

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DiIoz1dwiCymBJ2I1DU3O4UDdOCD1IYbLUI0voLUvMCBbKM/4INC61S/TdKSOoUevx63V7g+6/mZ
lHiHKW9CUA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o/flwcKffhg09UZzkz7gv/qZXGXaahpZlLeLvCPnGMHOV0tl8mkXW6lQBADTMwmBGUm7XZoObamg
kh0wsLz7sz0k84YCYY3YnDkU0s6XZ4yFdgj38M8k6+BTgeZETPuk8RfxBp2vQOv9zQhlLgklCWqU
H5aMJF7gqYDH9lzMxcc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3XDlc/RrM6J+fMEvhngyPf44nazd8NnlO+9fuAyN3g8+0X5quo1/68MLGc1czSBp+H9Wyu2aBKOJ
b7lFkbCJ13UBsZfTOKvBryDWOFa6KdkhYbTVSV9dfXRZ8PoouPNER1m+r+jF8e7EermzCIExWInF
5NIain6XV3z5eFAoF9+1wNHgh2DL91NQvcMqUhxodAC4EBuf80hcej88xks12032BecjB+B/gAMW
Fju2sqB0/mqHcdt7IfTqsGyFva1zLX5LMPhiF5YeiK1qj1zrDwFPgvhslJ9mmgozdcxNrfEp6yGo
skXdLgGuFnqjmzVIe1RLirf5OErXnL/7fcq65g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DYSqibotPAlt8I7+ZHxqG1W8t0MXnDrQyejnExd2/xGgdjHg+z1O251s8cO1MsyRynExFZebXN71
+rcOQqj1RiIoWzG/7+iJR/rcMh398jmqlJyWLU5IbIHCNoZyFsPrWxh/+WMiLYcvsaCPV1/bb8z+
2IY6rcDkaBrqk/EwYjE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
otEsDJz/b2bcmmVLOLfSwi5yawHEPe/YwdeYC6bj4QnDnh7iDtRlCB8Vxsd5V0BfHeL/WYjoeQM4
255fcpmsdbIm804UqNFTD5E3bD+pXsp5hjDUkd5BI6UEMxrdFYZ33Vo2q6da9Kuh+R1oMK735BRX
27ixqS9zhC9yoKM5h3EFDD4lGv1ah7oo8vFXQVvAoHLV46fz+yTbcdnzjY0CBY6ZcHBHkW/tXesi
gSqE+UJ05pdgmjP4NMP/1EbWm0c/tA0kZtZOMcSt52FHS77tvDYPPfsmt8s4x48hzc87BHtAtJLb
p2k4Bl3eRbmVYlntF4Wojcy6kk0ClpBDQDcHyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 32608)
`protect data_block
hrquASnzZlzqNWvQqD5qimjwmc6vQOv+I70IHdCWRQ/IaTWgK+4NRzhcWBhKbJWeJJxs88BHisKQ
tRlzzl/Ogz25s/U9xVrraPRVaDymgkFEXoDo+TVfpf+kztGBlrVpLsLs7TZh6vRpe13/RSBmuFbv
w2wnrVTnomYzXKOk2MewbmCR/DND1rwkfsA7DJ9h2QWvWgRpzzLnDVNexc3LnbV/yBQrnhKfwrPJ
cSkWwqdNccNmgVk5otiU3FeJ+TQr/bLXD3YwbGVMQqOnCPVm/05P8tz3D3HvkFYaIZIIBBg3H+51
1iDSiELzSxBfxZ+R/N5cLd0i1Iu1Urc5MUBiSir1/0t6FUY07Z87sRouel/XkEwzrhQn//UzUVKK
xVPdJHg3/1DWmaXImMvwPKP3L9+0Ev9bE+FwtQ5y8N6kEq6B8x0i83CoVlPUL+zoQ/TTgx5TJrGC
mJjGq+DyI1LcA74nzF18zi9W0+yFrWT4cuJS6+WqcrlRydcj3qJeawY4m7R2YGWEYO/A75UIS7J5
yNLLuUaX1c7+yyxnhH8C1Uxm5gMDc0dDpC+J8aV67JzStBI8fehMCNTuX6+tABVWTnoSE8cknehH
cOTOXATYpfqlLJa2NuK3hNS+83G4AA3EMbXgsbafBqtCjg/GqEAphKfPJgGD8RZL+vcEgWbghpf8
4yEQkzpg/2xoka1F916l1xztSMmM/a/uW9u1ciW0VjDNShxIUuLy4qWjMw4gLvRSToXu9Ve7GOIv
pa0VjXw2Ws8JmmjNpXuDxugkqbZanKE6MFU+LkMIH4pBxc9mYlq3aJDSCGj25gYth/lpUG5E9zJP
u4pkDo0KiTaRFd+r0WAZLfLOwp1VXqS4WMnAmyFL9duKNLLZESIppT0isF4oM/GFto/9lUCoz+Bu
ryJj+kzRDFMu7G08HfpWahyeGEXsbeDHD8qrs7abVgfatovk6oaj2rf9olNocX07QqZ48IZ6jow4
E5BDkb8bNOhA7fgMqMHyk59TyqP5TWMrmlY/oH4oLSMhWsSVC4bgPFT4Yhr+fIUK5mlsnS0ZobhT
xbD8dqvYFUN70XFn7xjGAQ3sTf9fuWZV6nQWPRUfdud602WiJGLx411AycZPVIgduhYr7nCKYj4U
e6fPTSUEA5WOttiTo3NiG0/z/sjRTmQgc8bbmP2Rnr1t5+NI21LdoG0VaT5iogfGksoeR47wZi8W
QmUNOJzTU6Uutz6TERhleL9/KwCge1laVAqSYxShegQMgvnk2TD+dBJNe8S5XDyQoPAEwdq6er3A
QwkI7+1yq1dVB1nTL50gRes9ywMYtvQ7j4lOitEDCfYhV8iR7AOyDS+XysYM8x7djwRqxUEfKhKt
hs6QyhKa5NMJBA+uMDnYcXgRoXeRpUaST8zZzWUF+/UiE+LnQjsIDFFUiAk7tdvlr6lnHYue+bDb
65ftpjipKLIf3kEl1EBkT8iwQYhwWfKFBSFsEUqGxflPMYmghNdVWpCQOdu+OrLI0suMS8I0Yltr
vX/bm9opBobEjIopACkAm0t53/uWB3KH9dcWPWneejgyJaO3vI3xnN7a6ppO7OtAkRXO5x29BMiL
H5ADXQELVnUABW6U4VJsj21x7nbdJUjCdq+HuBgsrKnTAYGtB9gWbVKUPahZOumNIMQdRq7VEQgV
w8dRwWX6OTJ50oG0fTlqj6mvtVroHZVg+U06SF0B3pM9TiC7OHz0ByMCxqRwvM2inEmZIpOp7vDj
++Z5DUMWowWV6wYvXCSkIBRQd/uKD/aZujI+hIj/DYboYQqXuigsnbtOU/cFwVzSL/o8BgJkulwi
CEMmKIdX7dji+hHnsd1ZUSvnV6EWTTEiKRMbCkfIKzrTN1uU6hqQsYKcrYEpd2yzOcDVe0wjtVyC
DAmGCuZmqsqjCFCXsLbtZmd2e/E532nve82hMDLIUN2np1JFid3Sexka8d7ln4qCASDBeF88NLCm
NSP2yUQW22wBoodMw2J0M9Hzw7x748UuBCFO99Yi07OOFO5n5hEi2HlXjLjq0ZPHEHToWCSQDakY
pwEtNEh8yLAFN7U0/5GIEoGqcfYl+EfZGZ8CcapyYIQH9dAxh6PkRK4FZMWvUeALJXqibJ7p05X0
YoursEEwB9nkpITbpxZ4tiiZmkv0gThZZJvYVf9XUtLKE5vinj+M9qq24qu1KPgzpWkgKTmEv75h
2Yg/tFUF7G5fJ3eBExG6GwCpdbwODb6bl+vbgjr1PK8m9IoVYP2jrLUjjcyTrsHREfGdjuUgUpI4
bT/1nRw0yj8BVRa9yIw6khN0pb18vDUUJvqeNG9U4gpVeLttpBQ7YT3/pNpz3Lj2ufh0aujaVuQy
OokVuwpzFe51hwo1c+7/I96YyMh9Bi7tPZFNCgF3O3mqy9/tokzTgpUEC2OyG8ln6lgKjOfAU3ZF
N8wrXbprDvf6u1zWZJfTHv8MYcj1LO/qoT6jeITS5JZ+ZGKBZFsBpEOc3DU+7NI80BritNW5g/sD
dOXVcNrtXG2n5N6FsOHjSsRDQKXelXwPsTRsqxsBgs1ObxDpCZzOw/Iozvlbyl/GeY6DfW/OxgAS
Bertzh2yRYtvxGciJQ8Q3BKuywE9GRt+xvzAGaiI/ru1Xgg0k+A49V3Y/WmoaOXI2x1+9yTgJmvg
yym0LM7waCC+bbDZDVYxcBk+PyJC+p9s3kgpgiLxaELTOwjEi+gsT6Y+FTfiFYMg7e15OjEacdwE
+W4Wk7rWqoxIK7zMZ565cxeocQjmYOpv1Xyy9vrTmqRumvbjCWHwIkN1e/FWaCFffbK2SO+NqM8c
7lBmzHC11WpWF/IthtGcn9Q7uGcqLKlJDMvLg7yJwQ1dhelTppfMh74E6vk7ch2+X/BiswKQ6sw5
ijiuCDxBpVUkIDTzDfiX56zOJ62xKJgcuZR++oLI1WEjyjmM4XRmjCUthgKJ0mDTexlTRT1RkB6r
KMfuS7S+DGPckvcLMFxHmvljOaALo8wCdv7/7nWDVtqqETpDO7li+0cg0GQG7OHrmXU0oQ4eXm9Z
H+CoqxtwGDNgqyGrf1/G6r05s/OnOhdEN4AtRSjmIlvPWWyX6+sqOSQIynrkFjtQa/h3wxhlH69n
Y6tucixoDmPtdq4FClB/3AXBQhKNVGnEJUnB7E8AnqFW8IR+yLP2GT4k+zEJsr9LB+lQJBrksxfW
aDNe7dNwdBZlb2moQzWTNEvFtrvnSD9fdtY1jOc6NjuZ53oBOAbtzzKpLEm5uD6BNnjFCiHWWjYz
Ly5GNc6UugSnhjbgGN0LthNrPcARrgQ//5gcSHMsx/9nDXWTbKTMFLL81IkeNKJo0siayTjSEGm9
yq61HIF1NkpjzGGbc32tvfi9uOn+qeuLOoljzTNpvajMnA4f/blvQuG+N5/TRM+8n3Yc0j/IOVsc
YZ2xIdt9sggDArwROyMOWVpZ0k1i5YCi4kpkBpQ80PrVhmreT1zd7chuXQow8B9JFd/x6WzuZOyM
XahdrX8YxKYkjRRUXT+Bu/9ZMEYFo5JF14kG7yPg/HlixU+mSKpiHapL3UW+UgzJNNlRbEc8mb9q
mmWOUttYFw7YjP8Qs6xT3mT/bfDskdeFlhHcHehKz26AYfF5k9Mm1hYc+S0RZIIv+D9S0vcC9v2U
cutZHX4eH+EAoJG8X2JWGfkjdIKBgFDkeiOtt299ZvN+x7B+goQm601oBqhuNWmvWC8si7+mVsVs
g4v3HNt3scceK10HZVXye1dkBWsQ8kMjUX0HB5u1imbDwCLAmGAdZfdU4Vzl34AgXg5rUHtFtmLr
CEP1mFI5cv1XdtX2QLroVp9J0CHKXoEFM6GfkKT6jNNKfvtlIzI6Bwm76cImBHpV73L/V8EstC/9
izf2HebjeqniotQitVi/6XUPD88H+OEingnmJVqjjKMDsRcDPPi7nzAB6IKF7iH4fsATXNPx8kRv
/Er/5116WlqW0KB4FUln6fFwmxp02S++BXtnXUPuKb5Ansv5CjxORNOU/GTf3AOl96R9z9B58btI
CMMuOM+tyO4zgH9jSluChFYfTPSaswY4tkuazgeSzpk5D6UeHiX30B2nLMUJuZ20DzvoPJUiIx2o
npye3J6xU9sBH95PaLyOirxWl9tld8TWGGXogi3QCVv4q2PWrV3UP/P3oq5ZtoxIlYWxN4iQa2j5
uh6XwSqSKlCmAyYIK79zKWEk1jXN1KpRsJbmQdPYzxLB2HPYyLtVXAeEDb94y7OAn9MklAp7OIVI
Y2TMbGC2t4NgeAqjSpIlMAVjU6t6W841ZgeWOD13Yc3V7Nl18YuEA1ZfyzsMqbBsydx8PEU8iav9
rEOuvVdqXntrbpO+5zLNjloRubMqMMJEfIMGUXl4MA9BVjEXHC0IX/T+7j5BFxYxOtOGfgwwK7om
sxUD7wZ25r9mltg+Qm0HMkRWCfuOQtyOC8Eup9GkScVfhQ5vCxOoDsqrWwJVRG/RQHfS9kpxDtYl
lw9o09+wHsI68iroJNapsdLwBv1ndKxN1LZoZ4IwuwW2Cz0rCd7xwJ5vBOPlqj/8DKgULfkv5Awc
2k/5QV8E0vi9ojzmoiQhRzENtrpamjBwglRuAfZWueE4ouYsqPyhXGJZlrqgfBSyYRRCrhlsfBJ7
YNMwg1HEBxn54p8vppqDYOKwd2CGM0BPDyyweG4tMvNAtsVlAQKvcFiX8kvGUEpn2vE4uPpxy080
b3arXafeY5n6VYGkilBHZWvHV9TbmyEDhnmYdGyK8B5KtWtl3SA7/dxWFAqe+MWpJi6hozqX75xN
ABONKkEfRkrpdODZtxLY5PWFXW5aiRwh0StvXvp5fiCHL0je7izmUnb1vjoHenD/ZFtaubqV/aEz
yvHfeUvZLhHHDauvwqdUMhYXBZE4qMaNJBOUDyGuXOccGyZLh19+D4/Ddvwr2Nap3fk/hVnq9qw8
LjnRmciB+bdUKcD9/AZ0jjxSflLiJTwcY+W9JnWFcPtEo+G4a4uclSvs/OTRxi2uCLm2lbqkmhO3
OMvSY++l8tEoMdvfJ1V+sSLcKGbCXwEypZOoIDmD/TPRAhNja19VBuAZFrPMG8irNmf0ROWiANvv
qk0syuXe+pFZIOe1Q1rrM8myBDwZW05IgSGwHpkLWlXJhfnNqIwOCC2dR/Qq9wwSJ3NlWDWuzSDw
UeZBAqyNkylfx2aXi6Dind1PXmcx5ZCrB7NsTmCxVQcFse3bsiLZyzlZHO8SxDRtNrEi/rI7r4Gk
xFnU/ujae/YuKPCoCLEyWoQobMddOeP48DbDoz4kY+ZKwaEfiiwWvoZw0tVj/OIWQlKXz5XdT0Aw
oEQ9RVn9I+j6l4nm6IE7WzuD0HWDFBKuEyxuZY9gj7PeWq0ijORGyhFKseDY8H84vUFE4wGKWuVC
Xpqe6rVLhELvwEa9jCEGxsq9yxy1UXR0vA/0p0JkT4rk7NY0qBuIKbZduPCsCanVtvm5GCCr9KSc
ertscg/KeUlHoOiMBMFjoWmQdPXMY6WSYX2WynqKt9LFhzGj3osEhWyPeIWiexVv+otkJhIuCl3q
0chg+emWsEFJvfR8QiTTACduSo6CO+uFIZ2svTy+M7tYcSzDMfzcK3KSvU1DDS+uibINUz/J0Vdl
YNIMTO2CFidn5+tXxZSt0mg/8vJkdAfxai4PPrcTTXsg3chCou3rBjj1yQNDTGmrveOWFc/m1qWk
hGE8JgoZ6gmHgq6fS1qG9dbXkfn1t3CNyGcGqzz7boxlesyd4GAKoY1oNQaKRlEc4InPvnwWjHy6
STgnUPSciM55BV8m5Ae4uSRvtDBn1kZHuEAIFZgSI+Of/8xodGjo6ogPj7TMc2cJ1uagwwRvAT8x
uO0yIKzlF93Fd2nspH5ouHn4uAo+zDX7DonQnll0LTAmZZoPQOr48GBa5Lyrm2muR1BPhdOptajh
bsryfjQRksOrWeGraxDcj8pWDn4nRCz40FXTrffp/3UfmS35WglI1Jy5ic8Po8NwCOD1vwLXjUDS
/CxCgSrmDf+YKOULWeJnEwEI3cDb4TsnZULU41dFh623Rv2XId0jFJ2VCaWXCBbyqIes3EW/frRO
1Ke6BTXr2DsUij0jWw4eKNhpnunfOqjJOA0EGX4e5cdyejIi7LlA5MotZuvIWWDuDHjZZ0UOQEoz
bZSXCZZZSFuLpfuQ3lk+vzuu3FmX7x8+Cg5BIyQXxR72d/dj+5f5RiMeZWoHgzy56muEtTSPxdSK
4uRXB3lk0PZtJ0K4oNgtPYd/epqSxuiLq8c7KZH/ZpfH5mkHf2/aHtn/NF5FUl4mXdEdMttD9Wt5
MZtIaw8ytWoweOU041YXbIeozXo29TI6v8rxpF5gvYbWMqGclwNzlEb51cOTf12UrMDOHHS6bqqq
3A+OdOWjIV0Ryp0vmcqNlUvgplWhx6QDorMiJwLCgtk2MWB9w/39A91JVMd1dlGEhHoZIDU5IpYi
v9ryuVNv69cnJ2PWVCl4mqrGfYCpXOBG/PRYOVGkf65S2Ao2xdZrweXskWwVwo2beCJvrec+TKHS
v7Pe0rHrwmJoLHDV8oruThQrzJflQ+YiWmCiMdun6SxtRpesBr+koUID3sZVMacx9j96GCwFwt36
PO/4OOL1MYzN4IMA+PcayAIhVa0vNyYzkZnaxnNCoc6HIcbKIpO56d2nmU90mBmcbeEV2JpKU4Rz
BuuKD6Pq+FE89g/8XsDm9pxMh7ahWagHWHK4pd0BqF3DdP1jpLHklJ7ae+nVyfblRteUk9qm+sTR
O266Swpkwhkhlpx05kBgQDKoHuAHMB3aajjI25ppB8HHiXQyLpPsdPe+0RfaByYWa4nKNTfqFJzU
0piqJkOq/lwbK7GVanu3TtcxbwHY0PTeKavnTrk47uSf/1BluAs1eHM/XW0pNRRgTbYw2b50gHrM
UB5Bc+CQIgUkpQ0u23+n98i50lNoihazOFNIkwDxBegDsYEf4uvNkl4xF/svoOkp5FTs8YiAoPMJ
Lq8xVG/vX511CmayiCXaxWeLvav0uakzFREEl+zOm/giSZNb1xspBAwRhy1NPUClXWfnmkIcJOJi
GdbJ/2oMbWkGhYd6PteKkyWeU6UanYFRUqMDcEWOiv6z7VEMgEL87iZidsx8SwDftc8QElUf57M8
A5kNqvEM4eF91YJVWP6/GCQAqns5scVhxgjVyy/pGlxiEN1j9XsUTT+umSmztUh2aZbvefpUzx27
2cWtPA7nDtu5pCLg1o+YK3+6EtZBguQiwEzc1gfcwfoM1qjj9h6ejh4wDLcdXozDasiHsFVncQzy
ve1Yr0GISDu6oMbFZ671vf0YcmYPZjpV3FwUALZS77v4jM6fkSsN5gPkTad6xiULgV/xVpzdmq1/
hxFIOIjl0JVW7iDKFetULFUUE5pKL/71sRZHnlvn0uOE2XpQrjNDspvWqstqcsnaxrclWBsEF9vv
mitHoeBXAze3dfipjUGdn0Cqkm9AnpXf1E6mYc8m32Dd3oNvvdkBWicgHKt1hOTLadYq7w2fYSJF
FcSFD9RhMl3vczyGLr7KLEAAoQ2oh6/dbWprTOBDAGLsdxE+ExHPkOs0Vq9DW7jPFmU/6ptfXF0+
/B9gjB9u+41am/4wTWX6344CKldrTyNw6P8CllukvmmQcgi9UOERm47uXvlUn3nuEPbFr3wFkhEf
hmgnDUAjxK8EyOier/GDqK8JzjRObD1D4cztWefum8rs3Lk39BaGX0b3eco/XmnJxBfN+TNtqUHD
mp9Ywk168aehiBhVv85+9VEOM0AXjl5B1tkRjtPDGqlIYkdowzPotDvfOKIEBovnGI2ymh+5Ji1I
frzaTagxxFqZe6b6EL/BNZa7XbFzAzdHALU6iZIzsAdEIc9ZGHUnBVQ+5FblsAJp2xLbzNcD6Mhz
qdXrudRP9COT5P3623exngoyw+2cG0TNLCxrvuueUMkzJ+g1hyx1tLN106cFYyK8HHQ+aN8DQQQh
Fm6gfdUszXgHt8w6gy87+p903AM/Jy0ouAPX9lZggN79zDpe7XBkta0WrlpNjvWf62KSRLVsINQn
VWeZKuW6L9pd641BkjMFhPma22VrhG14xQavIGdV1wVfs2hmDnsPECjYr0QrMoywrj1sDshSVOZr
Uq/wfV45z95u6hGxYfp2MZ31n4lEoHQwkR03hWQESR0AbP1F0uDqLMvBdWayuyv7NavXaxcCftsC
PdZHDF04RUbNMh0DHKBIvH7BXY+7HT3nD5EFITcfKmVbdbrFSLLNDQ+rxoMzYxTArgYQEmzt4jJ8
len/RuWWeNGhsRUopIJ1ek50+503/u6UQgo0nvDVyXUk2bLm/xhVonzYWIf5qIVcySwmfHfJyjMR
734TmbibLTGXTtgke1EqCT+IZ+OHfE8VZtj2Sfa2NyBIcNAP52jdsHlW3y+nPuDIG0mGHhi/OewP
NUJxfkYENSM3fjDhyZRtUhYM67XC4LQKiZ7E3arcntrEOf3Q9LiZKJ4O32ITEi7vVY9ViRDo9vvk
sE1zMXkxGJWdAUjINUXDBdU5YFIGIQJWfAZlAXiKpIw+EERLdaRuF1mi/G83nHTSHg3NzUPI7zaD
TksugDyhvZkZCrm9GnYUVcmESIg2MAe/AnAaehCLGiQf+sCrAL7VV+KjNTge71fVzKXTKYtQ04eZ
vv5slz8wfLxuqIhsUdkVwnLblPANqsWb3khXZyKogo0sJoOQb33houetduVLJdsCCKSm901Pg+nl
b4ipkHk7XPBetC/q/SRC2ldMxFNj1STtsZXMURGa8VZOl0imgIlyoQ4etOnxxOsz3vH485LFZUEM
3F/VLnOaHU12L6shln2GxNeYiAtXJgYmLwaQBGekvtnZDlXTg5Muqrs6Yls9tYP8UklJruVb1YXf
cX8Cwg8pK/I+OK3LI8TvEgPaz2aUxVx38XIINibpyLUr+hyAqFlAIYvNbI7yf2mDbbDjGOua5byH
mgx2/+WGPIziwI5QTYiXFDhem3xNdy9/aEoPh72/GfN3TAHv+aNEMFVEz0TlfPFIBxama7tuQKMv
hXQtmS7r2yox3MvdXUB9FAAwCg27lDyUtkgzUHxVIlsoiqY3O9pUsLZLd8aKoSzvT/Q0TTkNgYA/
N5QyUjRsqnpNvIMnjcuBwI+CBKxOmC0NvweSWVdyTVtM1cvSUEOMLc0VQTTZ1l2l41XXaFgyXQTU
DZ4+wWEZVtx3r0vXw2PdCN6sJ0FPUW0gks/+eOI3hgWy1613a86Hbio41+XKFJkfk0oktCGJ9Lw1
/lwt3FlzaKjaOEmCWAy/ZnwI6Gxj77A1grbDv08QSz90DqZBKvKCZNG7nRgQGSIx5d601+YQ+XpG
Cca+jvGfpEXL9z75YxX6yQ9lbQyy8E7wfm93KCZgetK6H2AUkWhusfj6mWID0v3NUF+1qhpU/0Ad
FAZRd2v1ZPvCu2QkBCHtMivwSlYwsFUMeitBqNkTCOTi+gARsCnp/vc9J6eFnInfhD6MNhMZmV+U
l4YA0gte/KtHBNjbultMMiy1uxRKCBp3rqp/luY+srq5rjt0eLXTytcsuVz5JUyIKoBebYon09wA
m0vRpn3Ko1tnTU9LH/C/ZnAqSyBn6IT4+nNeq9anFHO6TVKO7hx36wcX0y+vSZXXvxIyYLHfzBjS
jFpxXKHof03C+5o6a3FlscmVNo4Yn197VDihSq/9whgp5yYIIVAs5C4ia0LeM0e6slYBOWo5uKta
AQ1swEUn49Z5nSOeBM8Q7XQMKqcnsuEaBxlkLOcaAvMYRhDAJPiuLMy4VMH4o6HgGRp4zCFVS/sC
5DJ2SiJaRb69z1ZAVDshQdz9kpVKummvJbgJzE/pLWc9iYOZTc0aXYr4G+MrMqVf08KCmrvUGIZG
YcRp1oFzGTLZg/cQz19yxcqfeUANUuTbPBE6/aOws9Wv+Myf7/RjOGBlsOYdFy+7zX61HzFQBjQd
zpbRKwAJi0oc6WDW1T/FyZaONep0baKJuSr7GMh9wCtNcsCLGHO//uJW2/XEbLB1pZpzzppJh5C9
HGDy86+gUu1ZcAY2ynzbEWnqMQXruDTOcWCtar4NFOFNoQ42GCv+RS5sh5Ma4u4DEOFqaqEPNt8z
3dbGsCMVecYaA4lJDBhjsQgYjmZsfEyoEeJv1tDa+rY+5miXA7rOyjoSAueG1HJBx9ACno4/0Tb5
3W0wwsJo11hP1X9jVv7Mn8e+rBQlMyDlWkb+lR4JQeJDMqbelsbNLc0/zoq2ue7m+I15CFGH0VqX
YAcmHADlAoPbAREgolO1vzFICmQvXlyT5UuaQRT0+J2+OTJCc6W4py+WFsXpJbpPAr6Y0HfKCHzL
S1c4FipcbB1rRughw6qVmjhwN0es/Hjr6NghtO/8x8PqC7kWNilMiMEvevHPpa6IJEkWsvvP8Pyy
HoTL9mt20EN1OGwEIsQ0yzG6bWquvMz8hMG7FL51OyyIxH8kGecZjM+VaTWUrbKRPv+OW9Xh8NV6
Y33TiXJBzbWPddN5Z4D6Zv4g1AoCI01S76SbiM9eK5FJ2/UZQfqkwAYRCQe6JbL3OXpMzcTYf6lP
QVnX+9GijpScGE1jQ5GhIeXKl+X62xQjC4301xEESdxFO6Gdn5X3ZQJAjemKfDHLbbg1GA1Rztl1
Iay2CLU6v5cB3ajvbcNjCVZncpBITE/iLuLkbPY7cWGTvwpq+PunBg4VrOmd8Q9KRvOrgTv+Je2+
33o5n8CY86WeJm5xk1b23M/ZzWm85fZq1qIbguk/fgPwZ2YoG8FR7XdAWWdw1lKVkmHBKVs0lpIz
N9fKhiB68HSe+BUkClPfoBwH5CI5uV0gzITlWkzvzqpE34lyUxcxPCug2CvsEN5Obfl/BQ1Nfrqu
n7HsR7EtCvytV4xxZEOpGqNNlzXGuXbS6qbiO4VdSv+5cGETcmphlx94pc6uvpb6rN83/8EdY1my
KQGyTikSm7QZ/pTAtHj3GirRbDJ5vl0auiWHeS2QgOQiNakm4BbciXgezesz3qDIgmudkOdAAuYn
pb2dQVktsBKhOMMoqPLI5OGtSGFBB+O1GyNTRAW7lw2Z3nYfRGuctKVJSTHzROu/axr8vyHGpOA/
eGgTDpAHCcI4ApQ14OYgyNx5pqcURW2Yw7Sug3j36ARGIxawVZupjy970HLoWH3PMPHgli9XYTMF
kO/pR3asp11677IVQbAYTRhWYQlEIWU2DOQ0Sa+L//U7Qz8pZO7mSTJr7/fdnkDh+BZBZ/jUXeZt
n7sQ6a2poO4RUFc2KgCcwldzT5itPlxnOtyWMxVUnlh4DRzzIbcMV/VwXhd7HJ2Pc4fqkPrZlNRg
Hjk47+6VNVDGj8ydN7GgQj/C+Zf7y6Lv8x1mT9cjXy/bVWCgKCXmkaYPzSEqgTJtcYt4+PKMV+vQ
E8VLK+OslnD1G6un6kNkTWKushGdDxaR6RK0Uvww3XShFjuzOk9jO9ddyEN1hKDLZ7s29MP8Aluq
SLCsJZzGMWbZjU0Gx+az9VhmmfDMB5K/cwY9I6BWpM7ngLgurWlxJ0j7JAhjz8WxcZqJrjM69JcW
JRJRDg45EGRO9ECBWs6+wXhDWSHKlNPciTlsu50Qj9qxkDUdrRyOVJ/ykC1uUWrypk+e/BrMrt1d
tDaq/+jBgLaOD68Eqeyik7m2BzDvx81+NjFuHeKgq7flSHIsiy0cuo3xQIlEILq2tEQH6EoNGaW0
ouSS0k1OwRAB0y39sO3flseCgpp9FGLwzI1oP6hX9BTlnmT4gc+JOkXG7+dMWK22llZnmWWYdM8p
oBBK5v+HAokoubVYyOvkOkGj481HL1mCwFmXSJ1MvlKLdpKjUPYG+5+reFDFjCCLFip6mvZ0cjFB
IPKi4DSyAc3wEmrV/61kb5rVq4E27XdCdSSH1ibJisUpLakJhjEbJ0I6EZkpnYkkvtqUR3FGM8Wp
WhNrxRx3/Ctc3t9Kyn25rXPrL0qMskUCP7Ow9/PPDJk+XFiSJZE7/voWw8QjIvlKMbhMNtCiyyFx
8+NH4kI6tCAJK/DzLzPyEsV2DLRVgA8vGrqJ9G4y1FX5C7SCczMf7ijErzXbTJl9PWPXa4AqgYcI
Tmt0c14rz7NUFdnmkAUUO/TSj2I4wVLAAmvn+n+2aYKo+cHIaZqqTKgn3W/bL+rPcIOeZqMpDMtv
9MOckmsPGRWuF8IGe2J5vPxCes3WSHVCaB9fkwLjQF8RJSrUDp0gx18HNgeP0UntSIa/ICis5vuA
mKzvt2cNfgcZ4WeLZVuSIZl1wYCuxmY6aJh5kIym7ht8Q0sUGxFcbOlgQQ0PQ55WlxxcFP8nG35D
hnBmg0M7qxW1fcgKPiYHILRD9cSbzosAI7q1Z4srRyyZBuIpxQksfChITjT+Jmhd8UAlTxkc3L3H
DD/HCzRgn+oFwiCCoGpyaxWWs104UtqjRQkm1Tav9q9h2z06SyViscQ3FbmdyOS4J+xwG6Umacdv
Ufw5SiTIcDQeQA+7s2L4ek4hUSGCc3ygTnYH85bc3BSQeW7TkpSIh+HGAdCp2Gz3puqRJap4CbHl
d3gb36DGihokDMdDCYqFvzgm/OkiPARe60AJe1IaecWApHWWfYC620nq+T2yw9BgZrOOrGnI+v3K
XUjC37snI/Fd5Mmu3u1NGxPzJK2Q04W0TtDTNonaEDhHl3FZcNkotTXiVdAJ1TrdEHTLTDCl2cS5
OftS+LGWs/+EcyVnuv8ObSRZhZXEn+bh8d71nJIDlfHk2geP8zCy+b1Aff0Fypd3pNE0N9uia1Vv
HSANjQWB9rL4/oK3Ch/zfFBGqZzzKTFPAeCKCDGegPM0q2mIYKr5KnjzyoThj1bT12yXKYYoTCBy
ETYMJSW9VQ16mbzAWBTWuMZA8KtwgCD549f2Tvy6CXBKNeslSkhWRcAnhC99LtLl88mvI73/mm/X
T1kr5Pn8/E48ylvt4Ln6WWdDddx7UZ0qE93kN/HNvn0U+PSfkpRusTLQEVf1N2WsUsRZSfZ42M59
Uv9sXCkOHBpQ+mWJSSkeczyFoGzuwvaBeI37cpA3PkiY0viWSdYHUfKE/k0jFHEZpqThZsTCNlZO
3NOt9sYs8YdQNEB7rkR+FMfL6+csxDoQNQTCqXuhfNO0XqvpCRD+iit1rKMXnR7bBc2vUsXQlXOn
15rkxSv5e+vZwOiIrQ6wVh6XR4QniaBAF/ussPBG87sP/xyFpu1n7kE4T+4a7yNezQbbrC5SKs20
WZIR+K52X4I8JFiywy+AVmxpulfNpX5iamdz5T3dAj14g7hVTGQHVCsEFwbqIkLUAN7aNPdc1ur4
U600dOhf8c8HEge3K3Sbm+RCuyjgtdRSrwf0bU6ypzscjbWyIWeQIXXwp3qzavqvrYG8RGp8vxo7
eBbDwJTSMb8/sO4T6ptLlY8RoMkljETaitAK2+GxiLIY6GHT83Nv1OrvKhGT0/skcuetrP7vMrf+
gCc9B3jp9HK9dI7B0LjTbyP9DzRqq2Es0ISKxCdxZ0BxCypX+34Bmga8Kk76a4AjjXeNxcp8nblH
bpN9IDKAg3pY8OkzLQwNp9ZfkLTSZhJHOWb4j9Hqjc9sNqvDGc1240pmj7DfleRpi5BNlc0Ne9fF
rWu3G9guLRBseXbkbp295v6VjwGPkcxgYy3/q4s6ig9RS4b0T6dezWbGlE3xOC1EdrABBKXB6g6E
06jqV8npWJdOd1pkl5wlrC2OsKpN42C/LXJSxiKax+RoWYhTcjI/Y2aQr8Xvzp9bZbDyjHcZ8lXb
DjeMWYKwkLuhDt4jQmWmKTjwoYi0AwQCzfOmiFVJt9fKiaqrNQvF2yLcLc4dMUhP+PShmyoMDWqM
LErfg7tFraUG8Y05SPqeCxlsNRqpNROuY76YKCDZGA51osYgcgRx7aO04r6iR0HufF/X4dQd+IIe
JE0evWivOnFNN5II1JqPeDZzAA7GoG6D19Dm2wgTr1DjKLiOs1PeZIfFcKq5PodKoIZ6cVc7WQHN
42qaXfOsRYte3TQ6hIcBKiaI9gcpFaAoFnu1iAMD9y/03SGXiDsqXFBdqVDl09NytnGqxp4gu4W0
wvWZuFq+3+CXO6OpqSUoLioUXwjGqB3r20Jcip7aUZ2cW14VjRDaRPrYjNzZ6o2z028x3rXpGxHd
P/WeloOHkgUEBiFtRuLLuuUc2ROtuEvGSB9ACAzsKFPXVUbU9T9OQSXU72MK9ySBqdFtFCwCoJFK
9DMp23ewf3lR/zhJfGMJyoN4l6dAziZY8RXIytIab1doBB5E/U+VniSwj07iKwLQ5WKYlPAuYJKa
PZOGDrWHVN8UQ/v/WrrgHzY7xP3SVITRdJ2h9FGb48/ad0vRxx39vkD0VjQA0VXDL5tAP5TnNOEf
/69hhJ/XsQHl5a2rDQXbD5A7snCgMyJ+VIcyq8BPj1HSMS6KGIaCXOMLVyk9tgmc/09sXZ2COHY6
WwkesEC0l1PaA/GtKkhxBnFN+sxQuqeuLk4JOQVYejsKZ71tUxI/A80MUDMt3IaVYuFHeD4gnZel
ZlIZWgqyC0gEoip0UJw93+kkFc/k4V0oDAjJeI/fPGAhKOMophUiN0+jnp5eZTDY7lDJts5TyKGv
q0/NDgkeWDY1hzpucVPlnr9iejtsmRKmI/14MHIzvnEdipbg2WDgUF7GtkXS4FMOta/YlQ6dluxl
5NOGIuyhvTag09N3p3/CsVR8frSpV6i5mOGy6BgA4xBonFqkTTU2itXlihaNJc6wMonJyQEU2U/9
CJ/GoiZCkShVft+CLQViDzoh6a8ZnKxlRCZb69zNT19YzjoDb9jq3jgRnYuFz+xB3iW8pmTCJn4i
Kv+VahmTnlSaPh62NeaNBjyzX0+3cH/FO+A+m7aGUANnXS7Pu2azYe3KP1FAXUdtamdu5AibdyNP
qnRCkBh0deG0Xmw/b7dgBq/9xiSi+kZXbtQBdkkpFTbRhbPXRMPcnF17z4XzNZojMUDgoiGmKU96
nhAf3gy2ka+jSrp4N/x9OkieBXV0c6xL1n3tFySUUiVCJSzR+yUqpWjQ11kG9eON+ikma7dsS4qz
hZGQn4rPpyOBhGh5/KD0HuVE6LC64yNnCYBqiy/P0u+0B7MbbXySHYX9PP4Ef6OSK/J4yz0GZvtx
feRDZAAnZDfqp7CRR6USGjYhCq8OwEpGinMqe0fJRKdifFl7mMe4kKHqyjzC4HhZOZc3EnTFUBd5
F8f80vFBz3LQi5QfKu8kprzm/vpXb5RUAyIhQv3XuEAxPQ7poHuUVxVKSXQd9ftIZMAonUxTEMgt
hl0KOiVOwTiJIs2Bt1Z27XhigiKmVfMkHRPE+0YIT7wSu/UGSVOGBoamTX+CvArMNCq2Gq+n/jsr
wDwS2PFIb6ie77E2AWC7Zo0TfhFAarupOkEXY1ZKy47bo14wv489/U87/ukhyjGi3xqJ4o66wAd2
Bl2LAY5sl1iy5beCBWCAPV+IoI7kDJ1VT1weUgHS5X4+bg/GQerFWNTj7QyNUPtSrTovT2PIyvjR
b6lgIUdCe4nlmNQMfUh+e0nCX+F5mMcizYFmf5rjAw65ord6PAW9ldRywXyTfJgbNfVz1Hs1V5OB
mn//9r2wa2zmJg1x9iSUs8E+Zt45pnlHMx5oJopGeqrK9DrgLfHo3HOBNipj9uPkbZibgiCJRU4i
3WvcMQWV/TcwQaZP2zvcLsHwlyR7Iv5gYnWzaOFpSHJJN1bsKA/R+HLngxigtpkp+CEgGwWE7nSz
19WINb45IaV0pa1gkyNFDtrvFGNVxSL2XGKKSUW9TQquQyi4n96UjzjhnlhYvsM/5x0MABg8Ziwl
FRxBLE0hlDauSPHG+b4JIPqc4gEISxo61KiwJTGs1tmaMxiNJD24UYjROMzRL25MSPmrUSl449rQ
rBMEqpICuEQAJ3Yk9HZDVqcl/R5+98FhbHBiMOwnljIUZe2PwiNVOd51XH90xPMk3tg9qUGT/mGO
cW1MHmDTsgMHH67xrd7t4r7W8isrjF5IQKLmd5YB9J301/kdq/m2AnLMIzNRLcUo+qCYkLISiJgp
plpedtKWmbXRX6N5CZKok9YZ41zG4IhBnP4cyeM6KsIvCji9zwY4vlq1VUGcWtX2306UDrms33pT
aTApzBLuiJsCbsKB0qh9yoFLN1HJ2mvXLw9tuViBqEwCvYW5MGYuNmH2/yjE00cQoxsOVt5qHuiO
Eb9zPivKLg6hIcwdMCI/d38EAEXPdcLAGOrDArxnrFyW7StF/upS/bGKiI9WVlm0Ju7dCNFBgf6l
HhZoclhnHnPdBVDP0i8Mjgj+wqVdE1GQi9dtkDAi7ybnxYru5LiKOLADm8VgAcIw734WyNJFNzF9
EIU2YdPF1sjaiplLI2/paUslb6h7V8ypOry2lgz+TCAanmC1XnywODS7QTsxLSiaSbsbfRGr+iDP
+8M89fD0swnhdunFZqSjxQmSDucY1NPT9QwisFbtqWahQ655YqaiHUlc5oHcUCK0jA74vROlDSyq
oFN9ISJWVKIXiMD3sJoImINp/mSbXgjtHDisXSyM9NcC25xcsESja1l/1+JvsUkC2p9YLf6wGLlG
IKeiMJEjBHDMWJOTg363qJqQrM0FKk2Tsq4AOh7ujZ3PnVxGHfTPk1igbWlAcIb50XI6LXcg+fL+
AvQJdB3wz6gR59WlfXUMhr/8I/Ln/kQR6gsI7Wggj4gPxvcmqYO/j8ZhV46uwRA7Npq32+Nrwzcw
McdVzREc2rVhb9WFSJ3CIHSsWLCgSEuRJ+lLahhiWPl9tJIXsxuPq8mswcWkthWSCz5H5ZSBK/yP
/ixQLa9UUTVWK6vXwcs6L/qc68JypwM3jXQngCs11Z207eA2LBtDPxrPlxNgNp919N6LIJozc9j/
WhvfogsbSmChCqjqi2TxnCkShfu3tob8d/E6YibSVBB62oDp3yfgrlSfc3oi3ZYLtS8ohDRoU7P2
7L0mqxuqSZUWx3tu4xlZ2wxXe90QKXksR689hjRRLaxkyumj+C7UJEahvp4hFdT7FDox3aXXhUKz
9qUFifLI8nPHiu8Qh3yq91Mri+hgmyqvvylZc8mZI1IYIFaNO5U8mPidZkVHObyzoxDNaO2wYCQS
gDLrEAN+ZkltqW8izAIOiSnjIO8Zu5FrNDpRqRQ9YE9KCEC5L3PGpbs/sOYyPw79VEI0JmzqgRgd
4HTY3gm01i2dF83LA16N3KCDFFGZ2wSeT10dFtHUjiVPgN5HYE0FCZHBQ2y9PzsmEo2H24Jia/vO
OfhFSc3PnHXL4G/g+1O9NJijkZH8fnZGMDTOSsFur07hojovOKd4uCUHRr8lEuw696sWJqgSCiPL
ej69hxI5qibbBwK4TKv9aA0fRztNYEOupCXRa9MzLQhPCDFMoLGGrwaIwnStNsxNKWrCGsbMft2n
Ri5Am0wK71PopXIJGoXlD0FqTBAfLo/+mPjqhAUKE+yhdabrtzihb4uEswqycyjQ+s54H3GcRQh+
B39g18ov0IwlpCLzLAih4NMlIB4wkpQVEdEJar5Zg755vGBbRqtjlqsR6yevMhiaPoX556QgXl3y
4HdQgN6ST7dAq5Z3lpHHX49YP+2VyscQQdnEcHrMstC+5v2bZ9r7wjfZu49ggXgeOQcURjyCB6ui
2D9QiFwCKN5kT+akYCUH/KC0YuISbwDK0R4PheHrxpPh1kGhc7BU6ylJksw/N6dwy+yoPFESlpj9
mF/DqNBfbnRLJWBfLAFKXCzXmsmXad0hpQJxDluwUaLvdbjs+BtPY/NsNB3aPQvfvaVU1ssCEv1b
wkDhYoZWQq7zGQ+jZ2BytP7Ups20fcTvG44b1ceWNkziWOn95kPl3m/LOdXDz9m6zr+YhRnyvoWc
Y5Nz+J1TDezmQt9OMuMPm/2adti/gCz2RuJKfCEmquOKlF2H4IyFdIIJit9cWEwHkfXfXDjPmLUz
n98VTDMciSwFQsCACRc8Xv30mPATONo+3udf2oUSrGNasq5cC08LtCm381H6A2iADJomcbH0NdOQ
O1au7iOqtO1p7CZb9gUKd87BYBhkD03UfzCSWovUriJ/MDr/XdchDKFTeNX2M7kDWUXBtw6OAPpY
EeY8e66SE5OS3Y56NXwhTTQg5KHSjabL9UYq4f9UvSwESMujFcY2UfhyfyYdzoRQvJ6ePcrJHkex
IwALMhBg5Cr0YJw/wz1w1cTeg2IwqnE2iWpI3CYh/1umDjxyLsy5VKt+bJNIuByikXDXh/i9dZqz
ARAbFPS2QC+coIZxdD0ILjKxWSG0SXqqEQlSDWBgz2hYdgg2ZH8Rd6q+vsZfKCNV8PXFhddQ8qKm
nb4e2uPKRoPBTR1WF1xQvFKBQSHMZSmnexzMd152HpoiaCdVTgkizA4YWC3ZVDnrTpO0Im2Bv2sO
IfMxj4nNpo79y/1Sw8+w/0q0dj5lzXsy8ch/R3tJTGjo6vcFEx75BEWaoibwM9tVxFKmR++4AQ+a
TVxliNLkss/yOnsgpFbAYxROukuiocWZ1lp8+/pGoNYLpLy85jUV65TPJ9Pckme1snwooDs4X2mz
lhDNWkwRvF8zxqUDR4p/WWTMAARhQKmMaapCpJBkoSoAkgXav7yuZCw4AbB0MZRlaNPPy0i2ovpK
XKK44ASnL0oLLfOC47dCH4fLoUZB82HGijcBrvJB4DJwwKjiwPUe/U2DVsIUYTS1ujzXcdjYtU2b
MSuFLAEVffJbarcazy2yGur6TF3z8HzOtaRb3G1UKeWECiCUWPp0ht4AuZkQmneVRty3SBCIm0lD
On6f0cczaaNTT+qY66S6UtUzq4hxw7oY+Q9IkgACrAwhyI/DfIyRDN3CAglWfGMxQkNxpBbVezuO
GtDQle8XybarU/dBrzCuB+dWcpHhEJRwaPDoVChm3O0RnZv60PFCk7G08MejS67d/Bdyn/CgcyOX
+BvJptRotQztJ3ARkkP6imSxDNZiWOwTVEL2PXEcqtfBKjladPcZE6RNiRru7+p652IjHQ8Na1rO
hwt2n9cP4P3IlQoIZa75TwUtsFnf+OJBnnc9dy/syoyE4RsF0SxbXfW84HrV4tBMNSxzGnYsejnK
vvbIIOpwyVe0/mEJnRSvGmmn8qe0TF+gNKCO1VvQBmh9JMxVDqFMZc1WkSB4zQg5PdLZfE6jzx0e
BLtnLOshgOPlGt2NO28FRx7eqfeHVXakrMcGuDtk7fFQSteHzDiE1k29PYR4Bg1Yi2Bt5FPDlrew
eTz7LDgt8RfUhiu2Iduu99uErxiyEnVmfLp9ZqRfw/1rsJSlBPkby0guU3n+N+tsGeZDnQpCZtQK
8pf72NG8XCqyZ2+IOWnc7fqZLn+wDlNbM3d/ys/OjKz1DeZv0jnzSWJsAeyFzUQ7O21XkUW5O2Nq
C9ps3JJpwIUstSJ1Q2QGVJ9UMIbY33tC4TYH9DDYo4HEgxY0x/2AYTR+ECwneveqoB2Vlt42B3+v
hn//N6FwotIcuouOwCO3qXWhrX5NHaoqG+0Q9ILiSq23QcjKf9lKHMH62oRe3RsKVZS8tF3dT6bK
FuB3/wNh4WzOMWCuREdWv3Au+YpcrcBwFrvnMsKX6qqrcjoeDAI56YYx6/xn844KWAj9RK1Xpa5R
P5QM5ny3v6KLXEgesxteSKNHmCYp5VjdW4hcjFbymh13kt8YDPXuPEKZvsxqYBhii2Hu/rQEF4Py
bU3AzgAPJI4ZSgXMLfHJqtr9Pu6O4qsTbK/Zesb5MZMJWR8EZfu4XlsYNDfNlv3WtyH8i68qqHlY
SJTPM/Mc8Wtb0IYqnUa9E+pgy4OtIGIlSUD/5ZwLzOYirwzZAwPt65ObBZsN9gnGU6GXl35vcXAe
SzzYPl+7jjNoVzC/c+NdB8O/TRt+URKxfXYAC/wkwFkIm+avaT0GJ+a/UaJcu2PG3e3L9P+XXfby
4fUtDSWx7jsZMGX4qlJI0M00U7+xV0qcmSSbeog38dP6FV+/hVvB5mqzE64ErV5+sj5krWe+VJjs
SQ9JXRp/J1YkhhtOKdquzwjgfZC4LPBy3RmzGdbmcHYDK1Qj4yfYBn9C68oLeZcLrJIG/E50tKZ6
Or8krlMwIAFVfdvh3yfuTzODZKw/Us7Ykt9s84msQh/gnrdAH61Zlg7p7+F5cyAyZ8oPNYWasX/u
1dljNZ7bp51SvLvLE25+GxYK81qazXcbSpN+t78gCJHQup4FYrc3ElJLFf39E3YXcSqlvKkIRrlS
MthysJOAOVHsaJJFL33cVpWwp4L0vuW9zeoWsC9dEBcic8XKpXo1HeJPPcCZiWtSNblO+2MngVzP
dZy3qwiDWZEFFGChGSkk2ZyO06bbTQPwOJY0hS+0gCltjAioyN42SNC1pqI5seHIIAjOV5HAAcrm
8eR5vJBYIGUXvX6o+qmG4+SaMsS0WdZQp6SG4O++/HlKZ2EB9jT/gUPabyz2CUicawoJZ89eATgN
RJcI3fj9fZd4g9E6UreosJ1bqMC9zXEGa9LDLyRzO4njOfHJ0H4cKYwEZLgJH+y+8ffMmAVBjSzZ
i2NBV4np8EZ9Fg0aUnYERWDuivDOkc5ZJ7NH5IzYUYDRVHgFX+ECVcO2v0hZBDh8NjXmDXPsOPCh
+OWSO5/2dInRXbqunl0JDIWMuRMYQW1mEtVX8af6uKvU1RWFD52K6H7lWzesbVUx/vudw/xfUDH2
B3rEuJMOohXs399qCA7mkcTTkAXDxHVzh17mnZRrusV+pEfQc5jYnvhEvgWcUd1XSo8Dtmc4Evbj
5i1Jht7AswMpVSpY66gqeenvMudDUMx74jpXOo2rpM9xEpUwN146tSgATYe+Aq7nQiGHlsrAyCdt
DZBWjad8g+OGz/8NJ6jOoNONfRZYejGe7jtxJ2St3DvWUZjK5+AKIKZzXfw62E1Ibp3QNEa70T2R
cKMsaiNGb0smg8DsBK1e9Pz6DRKnmecHVVxKMTYcgvPb6c2epgYBc/I4TJNfgc516RDVQ3OAE9sH
X6fqYnWv1S7b59SuAcuVq7Sp+uydIdKMDilhNb6AipcKj1+IG1iyfTbfZgVyE8211WNV5/g5HGjY
9Awv1bR8IBNV22hNpllNkzdbA5OY+VbsdmCwDgcI4tZR7+LLk7m2f1Clb4Su4Xod92GoTlR895on
GB39QOlqLxwUk9lvny6iNsir0ccxi2QPmMV8ZHNx6lUDTkA4C8BMWm35AoAjIf58DeGdTaSglooA
fy+LQjbF1ZHi7WdVKOK4v+qbzLiKyD1wxZQZ2qhQ8WtnGiX3uJJklAAacGxOfFOlPJNnDjKd2EHQ
X/9U1v4lltXwiqoiyJTl+1WVzQd3riuUBRLT/HVxIldBQ6sXyUvsVNdlWkcUp+3vU0oxtOR01D5G
XbPqi6vGxWvdAufnjowzd2Y/+LoeHL0Q0r+R0u5nx2N3WAxkpgL69qkpuA/8oDN3JOatGMlWDtxr
tjJ2Kj01U6pKiOwtomLUtBgngaRCDmEWcjp2+euSQQavAaPcZHvO2GU2f4wFrDURF+pS8yhUr/Ca
dX28JQyunwwfeLqdsyvTrtW7YHzG6yRehqm3Lte6MxB+3zE1uTLZOXhLdKYKKwY3PdxoNAjZn3nl
8TIEyP5s2c4chGQn2Uc3v2qivspcnn+sSp5+9uTW7p48bLjmfzJRPtuw7hUTHapNN4Esvp2oNxuy
Ne4rRrgLqLhj4HVgF22J6lv13xalLtFap/tpXH1crYZIMwFKa3qumMxh3Ezq64SdqDwYqcj12PaH
IqQGH3LZujlhWA2+q9ae6EKGfQThU2wS/wwdK/cbCCyWKvRFY85XzmXcrStTFZ1iNm+PCvR4bj43
UX0wzeSu8cfb5SfsbBSOjdYZldQjxinmO4lVuRItRS6X7C0cF8+LKFGoVRkpQl3LTm+noE/BvMbx
720UpcXQnymubIyKG36tihlP3KmGzzuzRLs8jl22xt9muc6OHPCWLosSJbjR42wETrarbHEUZC+o
5E0xcSPhnLqXYlkXJnClZTqgG1tO65yHmFEeHTH2tuoT2aEwdUofH+d/7eH3FPabOQ/ra100f9fF
oRFSBxZD03VaWLX+uoC1VepexY1Ft3x70wf4E+aecP3i32RaEY8yJENuYwqV2hY6V6ecqJThY2VY
Ang/K4jLI29sAxw1U8FyStjHUDUZIkoroIvUeJapLYZ8IIfI9kru5gXP87THky6ucfqaC1gGmuAO
5imS2qjJmhElfoQAsyt6P87ncXvvxPDPGQEaZYv+2DD4wlV3fcUbQfisAK14ZydyfmPB6cqmGm4V
Aw7JXxdqnO5gZo7t6USB8cjWV7fIF8XhzaFgKlCwtp6Y8v4xiZil7Xh2iAdefUnbdXSN//Tm1L1C
Ko99VjJ6hW/qV1T6BXsnEBWNyLA26HsnofuN6IWHlosnAiqdeDNOHbwWc13TR0ww0qiysKu5dmRO
L3b/m9EppveT0V0Py6K2XBGi91vFQSVQ4tWG3HdPtdQkWDSyymUqntdBMCPDfyVIPW1MqTby2HH5
BDTCORYvGqsGa/Vc5E4FLm8iZdhF+xD99dXds+OuGBd8bhN0mzODmZ/1KZ7190i60sPjRe6FbG1P
RwFj/6ToCZ3Sjp9Yu5m5UyMi4rMgKaJPZJmwvAroKivb+fRgtcJ/8Yaif55aeiqQXdlLrtnp7jQl
FO9IFOAJr5kJggYjtwvl8GuN4oehLNi8ey7ea7BfNRUD7onDFR+55u9CBEptN5gsD12sAgY4bl1h
0HTF3ewFCEct0mp2u3AXr4Jzdk/TFUDEanx5SaYVLymCb2kKSpGxZCyZS0KxbJFQfSfL2y8Dj1mK
fjZ8TIfXZoZefhbKUXkyeL8Mk3xlgB1/uDwLr3k8nXPiiyvLMD7uGQhMNK419aJQQ6WEKA7K51c8
WHQtyvOt3gbazDWnO7HIBhDZ+6PcrC4DSbFwKgCekSIuiqc/GAhAQaX0u4AQJ88n9q91H7XA9pd7
tznRB8kTj542iI7cM3mCLKwnfd7OOvxvF88j2geKj++AeGANz06m807fxTi+iA8iEiLkeBj1KNrE
I6XrhxbgohjwUkrY/VHC+mceXlDEdlVJ/ttAuefyct77IHElNtHU3c8myPsNN1RqO0mpJ/UshojQ
1Hp5hnbPVSl9tDq+nT+Wb9zM+BCo4g143vw+ZVZ8nADmQJiKst02xPoCUaT9jGaX2yHYaUs3Pcyd
VDsawV4W54Lg9FNcGrQqokKctRs9TNEvY196uNkiBLCHPZzexoUdTbgAlx837ixMS0OO1p3QqUfN
gBFImME4GbeVM2V0XcWGRGNJC/aypYy/FvdrjM6TOR5ZfXuGHXNrnxzIOr4jTkgIOHKA4RfYGVWQ
tFBaxWP6TBbLbZ3agoZu5K1F53SsJF4prOQqZNktQFAr3TnEQCn9GegiLWC7V6tMvbOoFs1qqdMX
0Z3h17ll1hR25siAvSGFWqINh+JSETIzGz8tr7PkJeKBQ2+gEko/9cZVlMZBpWq2C/6J/I3e0MQS
eyz6QM9P93bWYM/b/tBQkRru+wfY5eRB+D/1GuBElMs4oeSDjrr/uB3Ad1P9LLEhXGlLmVX0xMhb
jAExii1jXjJUOrcR4Sebtw09LJbwwHB25ddUFsOW/34Wy8B5L8LUBWvXq1PJ/1yceZSrs1njKB8O
jM0XSdHHzOE1H2H/Q4UEkzApJvoz8hPYlzwX4jwTmFpNoim7IDTTJlZVjYXe4yEcJbynq/NrBxeT
2RMsgnTmsLiI+n38eh3Ci7/yxbTrYFUzh6qRwxwYY8xrPmJl8rtz/3P2AZhRq0mImsHxDjUuIkBr
hZylVYSIyqh/pSEFMEMOLHOjAGQSivTjQF/8j6Oe6X1NNcRP1QR+k31cBxzep4vpbj1T0pJXU296
Vp6HSmBATLu/v/rYftZI+/EIggaH2+rpEScgF2f6K2owwB7GvpHDRj0Pfyj8CLHBYowNo/mqilIY
q0p4xInYAjG7z3JORzuXZRzgAvkQLHds9CFUq9/v3FKl0LX3YtApoZRaoAcmWtxPym/6sIXxYU1d
WuHE0g7IEg4t82cg2PlsP4zsxvA4iWdqUE557dLwITZ3/8gGsey79yH0BO5Y04miLTfilLShsTLD
imUG8rU7jPt+E2WvISQRsIDnoCIak8pOFQZ2a4q5EjOZyyEXEoMyaN2HFwL0I/lMn4DsQ0smVXc0
fmT2iJ+eD03LBUjECk/Xft5VIQWVoiPr3QvGhzhvM9/8aSBh2xDA9iZ1rdwCagbqRnp/CYQficrj
X4MH6JtcWTQu3WH+V3/RLhn8Ayk+d60GYXF9h88BYZHifAQGAnmaMeuckpBKaisk5Y5K4ads9iqV
MtY1oAxGBFThDd3CoQunXSl4UY62K2XNFLs++tE+/rkDHq80oYz/ixm/fArde8s7RXVArLdNa/0b
Qdo9La+zdoJXsG0PY7vDVtIOlLww3mLsSX9NMlh+ikMt/IVCC6JdM4/d9GC6XcIKD/qcJu6UHlHL
yUAoMuYkbWQcEdGvpht1V5+KSBglHwRaYgUXx61581D8jignVAyRAT5mAVnv5R1T4aLwxVYau/og
Y31ftoXCAbpCqLsDCDivvklskb5UO6AUUOFSeqOAvFtq3S5Nun5zxHWhjpjS7YSbzL1mJAOgRwTy
JBBQ1oKX7h1AsCo0ZxinwV+oMwLcqowEU56kOd3QAdD9DnAcetFutO7LItqyOgaFAgB9YWnKlVlk
XuWK4RQqENmDijyp7Ck+5UJO60SOjTs30NtsAp3B+W/PXjuCtksn1LKzPLyhjn1r7MAetYSB1LAB
EDW0/QQC9cl/vOM8YnWmBAyMvGz2aPqYg36iCPRbO7NFPBBZgnDpTc50IWy/TU88STUUuyF25oLO
c3TQTZpuMeHRazaObaIsL/RPrCC7s6sJhNu1uPsrW6f8krs0fw01HRWgVa24zh+uqkPsB3So87f3
C+NGkTDJMxs/LJR9Gg8rsImn/sMthmQO7GduO23RLWfIBCzZvqQopdWHFOXRrGtfkfSaKPUaiChV
bb0G98wNf/OUv7WdOcr0KG3STBJOa69VFzRD7BPYN53kqTVHjDDZ3cIH071meeBtokEbxn3QCumf
NQkrfYA9rdNrBKhJe4ve5FXNVRvo/plVgrrIDfXlDY0o9a5/CZRfzqTlnrmT+/k/ulwvZEwoiRJX
Ec9hbkv+KXFQ5IP23TVIhPY/vwuvrlwAX20BUoHqrX2V/7R0V1lyCfmnqYWEOCrmhJLTiPz8GM47
EJwyM24RZMgm7RGPQWAlYN/JAMWxCC2i+GZZCVIaM4u81ARQCMhitUQigq2PdgP8oGA//lKvNSMw
BD/JPUug3+4A4F9Ils224Vm3BLylsGvOEqdhFctF8QNkT9scrYc3Jcx2/zlenjAcG7p3PmVvSa4h
aTL/dQFgi8P7QwGaausEzre0H81SRLtY0unKdoSix1C247Tm4GLekYsV6uBUu5MidwcUx7jkXirE
QZwv2TwwEWyCJ3gceOg9WPcDvaA27Z9y09woOTPvQuIL/JL+AHWEO76ob/J7GjIwWM+f5h56fVh/
O25avV3krHxRG8vMdQvLGIwZCTC1sZQzssdolNRLxcSxxHzBUBWkXcSJTCT8cLUxZxkpdu5jM4jM
X20bogi40dA/j+G5e6oXTbrhruNM5Fb/9d5xP0+xndq+9appnafViBMghVFYDceuwZy+Kvslj0Ya
VDYL1t/ZIKZx0AwcD9As+FUWP2jNZA3gcvw+S/cRb5dNPIBZcw76ntK8mInzXY0Bx1uXSNEnw6tD
EztprNrmLbyf+k7RvP7psoML95JbZZcEjcLNFlgfquDpgrYFhPJf8Wl/OThrgM4qL2Kp+DVDPxJ4
WFoISGZ0VW9jA3K/ikbpPI1fmvYgJGY7b5gk4zkUNpPovph9D1Cohoc45ISlXf8/lA7FCc5KsAsh
4ide8suius9F+GxoTiqI5NhVjNK4eOUwPo617H3DzNzvmB78DUCjzS4Bi0nlgeRDd5jV2YSSiFUm
LO4f5v3z/L2RhebQZYjG2hD+wz016de9lLsC113E0fmHmDZPFnFoKOUmQf+99JVc3oV+xJBlZRCy
lPzaQ8UgiEpjswlvpZG5bgHqR3V/jEr/G6CMTQU0+KDay2oP+78a6hiMoRKlHoqR1qbx5o5IGjoL
Edda23NIfD+XAlS4HW7g0KZO7+/RDFDdPfgAp5VuXS3ZT3ZljusadY1bfVJtXYZbDOku1HkM2t+g
TJw6vA7x+f+Y+QHN0UhCVXylUsRTO9q6flOqZa1oZQ4hr0U+RsbtGWTKWiRCE/+TQs4b/4nd2MGl
wHz7dowMhky0ieeq74jUX5S9y/lAOpBK6PYavzbaI1eyPYIsZbhqP6rXoBRIE1ht7ZgF5fFtGIrR
57Jkg5zNPhQd7g4I4ZDLePfEWX8p2OEXFkvmJFeIQSPU/CxBYiBmvG1kDyvAm51vJgGTfvYAUtgf
yi8C2jEDimBPzQagzSuIwqaFkzWmgfhGKXutOL2PhRXAQBkqFj5bH1Ip4JgcZ9UXqhl+GJgabqx7
+q5LwgfgvnoFTttIMSGyFgNb/Ut2AA9pA/TSpDXC+SSNucRr3tWm8NbNEnkHlCq/AFOh+rpDlSAN
makFShxIh+o5EZxEn8tb/VDJ5vFn2zh5n8z7f9uwOeBl133ogsm6tsqbFk83STMOXdzmq4fRhIoW
HGBmG0f5EyNf7H2aMP1Tt48kShrmp8Z/h9N8Bmx82r7jdG1wiSx4GP+Sv52jViS+qhEOaLVsAD/K
H5h1wunos0WV/rPW3BZ2wPXZoV8y0gtf1qsVaIAHgtk22P8sdkSHNT2zHFXQWjIgj2leIRnaia4e
EwED+rvyOCT+RJu0qXFZeWoxZ06yhn06ZmBY+dEaNzVW1kR3buTdqWzvSU1JwD1CQ3wjNK4V3l1W
J6AlW1XfCv7izyYXUaEGM4AqFUPbE0RwT54BBlI8Dnqlyy17dWFDN6muEfZi7yQI3F3MssVvaqMU
d47GflQ2E+7ibG5g/5E9+Xb2kAIbJg/gkaqgkpYoCX5cJhtoRVYj1cdrF5AtC/YugIFqkp9TRTGf
C9HcJbA7CLPLNKaI2gSYxRYcdk5XmK2jNcHk5D+FuxpBUQsOwNIhXunR8lHgfFu7f5b908ZMvPWv
jm8UVkgGRzbMWXP0gPr8rmgDfVphTxU2vOG5o1suyBfqLNLwE/GUPmxP9ECtCc+aqQJl4E9+Xx2j
bpOBgGXotp/JDRLM6feWMHUf9xPC4U01QE9cmN0aVEwGlhsKUL2sBt7MrDsssEnxfMTGIQBlW9Ab
a8tNxhfjkDnGzch5sTUd7dNMIit1ftqz5vWp3/ogGk1Ddoid1PrEc4G92IRp9Os5VuUSLkcQspZB
kHfnxYQnqgRCh8w87RMOKWBi5e7JOnLBH9z4GpnTZJ9K8OUehi52UWiLAtj/Wqpkb2kwrt3aWvmV
/5OiT7nb/6SL41qYeUg51WaLBrLcE3Yyxo8KgyvQk/dc64jYqNIblq3ElrjfYiPssNHtoyZ2kSFp
b1HoDy8fxBbQYoELfA/Y/DNosPKYXUiC+3ZkFsOOSiP/RTR3clR5vrULKAGdeiYVpgnOvJQWK12E
Xk84+oVdASF0Rrke4n57AF2TevMRAmwl8RwIAiFvwqFTf8EJe+p3JW7Rfb2olCES9MBNN3xSmwz5
fGHjaQryit+4B17a6k2vqBCkYW7yKrPpjgBp6Dz2qdj4oD9UpzXu/kdbhZyIpBZPJzYEC5OPeT1q
BIZGF7cRVH/VZYWG50tLcOMoc9081IAcwOqYMWgBgXq0c1KMn3T0IRTpqa3XWLz8KlvGJ7KQ3Ip0
wBjo3S+8yYAYLTJ2clKVU46JvW2ywvLO/8P1cC18H0M1cwjyts3KXbvAJCywhDDSdms/se1kFrOj
lrni386Lm2fBS3Ocw4MTBIMha1ImuO9wYHv3pjY91dLX9+Z5AriJmTgWncRERZPmiRSjrsTJK4JX
xVqJjKDc949ah2W7FdmIf7drdjy0r3km7JrMsIGlNfmw/+ArBl+tC3Nbz2htmfhQuwddBil3y1xu
B+4IQ0ZknBvTLD8fXykEVnr9cudA/VKLmtWMXFNwjynkyIaQ72si54OUOA5psbRm2VoWCSAIklwv
Tgj7owY2ObUEWDlNel1XNspoF5euoAPulLeQaXbkrAgnBapXtg01t5tbo0pIcj8xrxH/YDPngVBQ
2TwabO7/5gdLuzxzagJXimSVIh1sqrJ7DyokNwQy3XP7yqzya+QdHO5gCKcfGiZIvsC5fY118z/t
lWKiL/gxcEFpo3ATqBrxS/3oHg611lR2CfvtBFjHtv3Hr3ZvEpcTWQPSCMx4mUi6KfI4qeIyGKqv
6G96s15OqWsLeygxFd2wRKVEEUobOfMWniYKdLFTtSYXBjzMOB+oB9gvT+gFzzkUmBCPOcrUBvTD
WeC74jXPUZlgho93SRk6rfbQetPIa7RiAmdkBBw9xU+GMsmFe9prdO7pvLqOQESfmNLwYkz0AKoX
vvfixWQ/TNE7rMVq/wOmyrTRpmjUGvXb/vDinXt+EiXp5Zc/L0fYn7Qpp0DFSaWY20Zxv1S+GKc3
r1xnz0F4dxdm4YiFx4Z20+psELwBceUl3K150w+oRuLAhGfaFL9n4EFFsDz29kRvXYhPpcyCl8w9
9KG8v9440ej6jchz6CATldB7k8jFSrkH7k9eq19pNSJe6rwKhS+ptmra9QXH/SA7TAnYWUiR/YuO
IZP5QE6AWOdHh4iqrYPpaTJT5yKA+QLd3SIo1yJNkQ4h0CQXCzAntRTQ8E4ajoltm3IybJItaYbU
YQekKWQsQoxuJd2ZONvAEH0sbK87nXCMUqf6hg4rDT8Qv5eiY4Cf9qZGLkIRevykO3iRLqCF/5/o
eIwYkwwFyJ95nRhxXRB3SoM5s6XT3WmPHB02c1PCDYhvVwueJLbuAqaOmRSqlnRucXeWkA/FXKyU
krMK5hFYc4pckEurWG4be1HhPOG8gaJblQHzhN0fi187DxYBBspHBKMQMoZuN08o1iSN0bRmv4ZG
/ThRKny/DAIdE6UVmIh1YJLUpV/bdFav7au4CtvnZpa/y4wbUUR/MC8973GrInqyOrOmQZwwPlpj
iGiniidQ9IPJKA3KynNtnkRiUQox2zeh9jAgLBuIs4SXTJ5WHvjUb/4TnOqmg1gkSDTsvgtJ7NMf
YedV2I9y4sKroBX9ldj1TCsac7tWO8xseuRqXH/I8C88nsv/piJ/y+7s5gPK1yeXzec1/W9nYIJY
nSfqYptinOfXqEPafhxLU5PtwLGcfLrSjLY0gZGCdLXvi/bf67XF+GpqPsHuAUtmrfRHzzxeb1/y
rJ73ruwOAP3y3wPuNNdT81Aw20pmY1+MXsgNChfGPEGh798LhUmq0O0flX/AI9/LNl3pBqT+cmv6
9tfnnq8WYaAahnu4rbk5iyAOP75q7dFc0wdpCJtYrB0xcm4Axpbz7Q89WNcgkNX04hyyyD2Qn5Fx
2+H8DGAQF1RVhYM2L9c9Opv6YK4ZfNljdSKtn1+rJnHd98wO2z/8SWam0OCg6lrUp+vnAlytawjK
HqkHonwI3BzniQqwglRqf+idV5Rc7kGlWF9eCJFUGkfR4tyxQhcxu1L5otlLGmihm51VXcYXTTLX
Rodu9xDPhUlWfybExxnYAUJ3XEgKy4hHBlhmJCUagQKvmB5M05qQ4Y1Thg6TdNUCI79ZuHas7XVV
atQjg8vWqVh0WSNl1NoNEXWlSAJZil2LDjtHNBYbVNOO8xKAw9pMJUcwV/N3+dw27+79ty9RgiuC
sKw1ohz2+gt5lWUamwp2ofGEleTybJggXpZMwRaYqIcg5kUuAx+0VDw6SbzTOZ53IG27T/a1W4vO
NTdUMiTCm3IF8l/INl//UAWcYr/tnI5FdfqzXVfQ7CkdrKFdYv9/H/24Jh93lrLNMhI/wTTK5QM7
17mKBKoZuG6DVWT85fnTavLEY4FKGbc+l3ociaD0juICBbiwedOh2OmMW7PdC09nOeZmQyyoG5wZ
4a2W0BFE1QWyg/ZdavT0UqfsRENNqISathLHvGOvBo1ymPNobz3t5qD7byUQGrn+U8vG/A17Drmg
CqUmEuFoV1WNT+m47HYsV034qf7OkOGQ8ZUHOGCNSBobdM+sCRjUgLD+xXXcfKwqZwnX0hj6iOL5
me8w1iCvrkkxc+CF3q2H8O7kbLE+X1DoZZAn/FAgKXcaNHRx8fQtqovLo5OKxNSMOg9QpM6i2pbo
mIs+UYUT2xTmx5s4AKrc+RP7cYr7tYrEwQsACRHe9RONQsqmFlLwdPF/W/Gcek0VV87a9hDnC2ns
SoldooLiPZuTsyIoPobWo65oweOEb1qKoUFPymEKtnNRAASSSeEK3BZWvTJsA20zL7q7x6dw6HWj
Vm3XFP3dXhkukIjoSx5C+hrFTkkHfuhq/Fo3rz6E1c4dNtBPPA4jNmDxJIfheLeWkL207Rj6YvF2
ccl4i1uuygJmStUaashH1rvmTecYVcO0a6pJU4IeBEEou6eTMuIuQJ+UKSDPmimR4pKRNqem3Ds6
5YfDpKLxyun1xjNNnDQnm7tnxyx4v+fAfacr5iruVW491AT5hWEJxoA6taK0CGCKJ5LE0yiALtm3
gId92myCZu915KTp6pPGEIGL6mjCJDINxRr//kqVefXrnft42jH9KJZYVzTCTD24/rMOTDWU2Cb1
xAoTEYZq3cbDovwzKv6Q/sQ0zRTAJJQROf4jKhnks4FGMoLbZSFJaPNSP7ESARLvVs3LC11G2rS9
BvptGzaF5//TWf3QpaOP8/cqd2JzbxtJ0dF0f8Tx/sbyStwKCers8YOOB9oBB7aeoKlB3A3tKdDB
HqIvafG3kyY1dNI3bw6MXtmKsmib6bHMjINAe6YtQaywUERsa3n78yjnVPS4QUgYUJUcin+tYl8z
Xb82rGxUtT4xBkPpTD7zcvmS8Nq7fdAKDKkcMUq1oNBwwYb5MkxCc4vMBZgYMxBxJGA758A3n4PQ
wtDkJqhKDf/eM4XYUllSpvmlCYXYnzryfxvtUvJzl0QvhXwQD9/k2ZBeMMV0h4T+ibL8/PirQIZt
QN/hfCLITCVxitI3I8g9AEZNbPfGoelFc7dOAecC42F92E15sPN2BLa+WurhivYTNP7K0SI7HBbI
HAxNYgOPsO/TH3mHCmC70fLlfpduvIP18cVkCIpWQKOaz90S3r0Pd7n+MgoOiKZdfCezUGdzAJ3+
kv5qXbapMffI6MnNQmUk7M86GV5aUHZOntsWkG/jsPhPuLNDRw8vWb4zwXNDdE5Bk6nOQfgE+L87
kQBgQfQ6c63obRaWogwZjtqiYio8gCph8uDdvXDvePLBMKZIiZrz0Bibas1ReLwEGGK89Qx4O3qL
l0LYrhyOWie+a4gSpqzC4ufUJi6VXohdpvGiBCNKFoNPrIA7jkpbgenXAj9023DBYfOygQ5TdOrN
L8+1cw4/eQKP28n8SuO0mh53zI8DtrdZWnZvSAJ4KwL2/vORuKbJHP842P+BOj1URlxIThqHaoFy
KQWcDjuEQ1zGYThDDxcAqT3kmQ4/4wZ2wtTCHYwwzU5RE5KSw456zxeCvnaVXRvzQU5yW9FqOggL
kbG21PQMWJjioNfO4nRQfKovchF1rqgMC8L4oy6/ImYjFRSzzB2HrqOAcJXvAnYK8xn5GdV9NXSQ
Z8YGcIuhzmPOFhn6FDTtPFVuBzpPZ9Dm+Qg+xbcABdBDeIACYUu+AwLkfpGrCMDw1LByS1GncaVb
sZknzTWVXUNP05boqpV/DCpOjTz+WXUA0wPooB2IAOKy7CZDxYmnD1MPxz23y2BId1fI1nrdgNur
j2DTfzqyJCnyVNwazVlp8idm89gI1uz2Q6242uqkmwqfo4HLfqCVHrb9U4lcucEELBgd354/Ae5R
WXKHtK7uyX021iqzurNm6UwlglHBFkORqiTF7jzb8JL6hEBRcNdk5WFSREDOy3ZJJdwMMz26iXuk
eMcGCTz08YB63Pc9bz7bcSY+3vherDLDyalBHqqeeRn2rDVR51EObtasjWu+XeGYJ6WLtcXrbis4
ecG8tJRDOt/gGaG51hjghrOmiUHcwJPjHXepEnvuF5FWrlAMNgQnPyBPsw82gzf9APMFGtWWazFX
orhtKVluITSMwBbiVwMI/UypMMqbtMX1D2hN1XjgUQl0SFOqBkD5VpSa+Z+cdQXYY9vaL6Bu+nSK
8gsZxjmwnpuAWunnyHYkPI+q6OJqXQjhrI/OiTIusPJ5sEfzL2ePb0VocHi/8cGHBX/2qPEw4XVO
mGP1/QThILJg4GTRgCfgF+TRFKQmtpnVIma0G1aT19mKYtRi5FFlBwj0NI11/eT/LJB3FNeCK4+K
dFp7EGQif0qkeLhPKeSwHDEoEPbRXM+IwSzOJ35lhzrpEvx3B+ygY0a+DXM3t3dgE5mRQ5r7uSTJ
CT5FAJoLtjGFbhv+WYsVorMbRuwcnSr8LA+PQHAm8dGSIc13MwBUyMizf+KXev2UTFes/v316sgy
uFluAgIEuURsFTfVy4HrKFyiZBldJ8/nuJ1905OG+l3sDi2gtroUTFW8UeR4A7E0OBF6JSWoubI7
eMwYJ/FsTeMotoP95NPaJOJ3fTT52qh92Y7Wf0/du6m/LcblmIKhEsQuLTEpyAl61XBwJy4gQB8M
J4GEDQHyoZ++un0cIkm0xEJm26G8akGfeEhcF/EEYJ2Iwv3xJQj1lQT5FHdHw4bUZA6NmFyN74+H
olnuKd9/XvQKb7jqr20cD2lOQ6GmnAO8MiaY8MgqrXdZWEfUxzB8VzMKnBvWabITftHmYvhoXEdA
HqnZzaA4Uc2odCyjuMtkN/2E5QzGrpxNxU22x/kcMd3In+w/h7Lf5z1l30zxD1GQBblKm9nBWjqs
6/R7vv+1rlmjsGxjNb+NAJdf+zVe29Q1HoYxLQABbmHEzyrgGICCT/52AMwD8puY9nAIQvozjRGO
oCmMwKbasy3GPsFWtnLBBomJi00mIxrxnerPCal4vDBqcSaNAWXU41wNCNjnTzlf1hzPEpqFWME8
kyuKGvAR3LX4A+KpZwPXpBgLszlBb4jpg5DBqNbXdM6il/lYjlCJgzxEOO6OK2w8LsYQVzA8jyh7
s+n+tczEhlyol/NhHoiYxM7CZlKaQe57WqCY+ZgjSOj4lZdJ9r3QjtMkSnBggNN4S/cLTyyqlZlf
XrFPhQBt7vbDVdybJVE8q3QmdKdOmvmIA6n+8fOu1/vmk84FlME8Qfek5QF7+3sJacWoNALFzEQV
R9AAYqd2M8l5ah5ANFnzqwlK5fvGCjxkhomR448p8QJFYeoRyEsLLDyYbqEynF0KOpprGeGv1oAv
13/ztjB9Wcg7W91eUJqA/wYcxj4eAD41ZJmveRr8Zd0ab88bEs9A9tHJ8QH7Won7exv8MhR2h4nP
Fl/lDMcqVjtCKO7SEzBrfFcP25x/DIthurmyAs2yGR71fsYCfvbN6KKR9PnakJ65dznZsOErNRCY
5AWExKa7unGn2z0EHyN+yWIZTFxQmGbUEhWssp4W1AgSKKNNSKGcn9+KGaBQmdcfJcgaFpzOItvT
oz9M6YOVkdHhoahb3NZEEKt3es8jJUIp4RUc6MnuZmeKHvLe7NzKaUH4aVigqbUx2US5/7pC4vr/
49enOgXEuB3HGxL5dQkWK7gfh3cWrkvwYknxqx/Lu/coaPuSCX0ZNg6/5+Z3cGjlFQP8QnQrYEoi
AH5fybY4C6m264jo5h5I3khCbVuI1AyfaloNgSW9O5QgDGvVmYKVewR5zUQ/W5b6pvRJB6qvXcKC
5Ejbd2kE2Ia24XjUCpOBdLWojzpMsZcYMMN3C9SaSi897aaELqyy6aYB+UkGZ5zQ63DSivUZq7cO
ksnLIrcKkepWcE9ZeuNDsE1vwfN15+hVF5d0iUH9gERF3SWNFAVQhAd7p0KDrgSiL4kv0Yw9I68p
/+sjVSigw0OlIlxS3SDVC1JFy7LYCeeMNaU7Uz0gKe5UJzmJyj8Mu1C7W5DX/hEbFzg4uMwj4Hp9
lw3Vy4wvVelAU9pu6a2vq0LIWfM/0+Frog4cYTF5gx9BzX5fl3+BUQXXjeTeM92tN17AoaA07jlz
RTt5TZpy48iWHWi16hwseI2qSq+3+YckSx098ZhBgM87kXcRfkeAtA6hvH1GSrXMdFn/CQ0bQEiI
5FRrttu57gDcRGIDj2AwUSfO21exG65GQsIThxATyNu+QvyM+7M7x+sAfCAB9OjJzWorW0cQXl6f
DClYrI6Rv/bK4C3OEsv+c8CoikWTGYWyT7q2bLdSD3T0MA5mCpoMr0U5jBybFYwQg5eZLodNcF0u
bZsUNUzgRhtssqt9NXSRBJdY+QoV1+TKNG1h7wSPYgz1mkPamcwLL8u4tmeC96rwmKHuYJqzvo/A
s7kgzry9w3aGRD09FkbiGRHJTIlr9gIL3T588KmjZQmkKU9xE+ZzwOr6lZIZJiiIGF0GJyvHtaUm
RYL+6vHpxMOnUYN8+uVIuBDxgPDaTSDuB3EAJJp8RBsLikT9KrZEgCjX/oP6DYiu9q1PoAgixfdZ
RVDdW92hIP5Scc3Yl9EOwgCTFnS8wKyYOgUn/Nsb0uzq123u1HLgHXW3jInt3mKGUrXClsc3guWA
zm7QT2Sg4H6FmcXdFfAO5S5z6GeQgwhF3ltJZ0hWKmyqZzDBt9nBhIrAq98GU91Iv6q06ufbbLtx
3AwpwfcW8D5EuDjc5j1bW27lloD1kGwoIU+G6YFOg0XZm1bEGVv7ow7z7J5Jks4MWVr1h0U0gIq7
1cp8ZdJQr/YY0vGPOliSSUE2Pfx8FARxhnGKDVlgRjnu4n12vm2+geSBjrPJ/pvYvoChkPfYZ45p
BCI84cvfjKU15qm+LETOKacmXaxn3xaGFwAtCVim8/DyUmQtMKHO7naXvbDr2C1lb+b2isnmUJ3K
tUmZ3GnJcCc81/xFGNqptJoCg9o3865O6/WMjOfePnUz37gi+NamD7cwe3dNKOhJJqGrcVg+9RcO
qQQqTiT8/ikp5lzOg5WrHbroP4R917y26dzPe067kIepKcoxCJFjkAwqNPmGPuna5OTN5bRuenOB
wiX4fnVrtNd2HQVEPP9vwsh5vL348gth56PPL9VHhWhjaakPEoF8ZVFZFsOO9w32lhdFEeYarcEX
4AoPO+vNSkrkTRv/ED79tgE5aZ5VDkdGsMaKF8nUK3OZsP38uLMeC3sPjWqatOfDbs+3jWebmw3Q
9tA2+IiReaZh604Hbva+wVfeE/xZMBxxoR29sWAUysJDaAHyO+znxn4GEwiYMVqysbjV4t4p3F2M
q+scbiuulnaR4dszhi/GPWOw5/QxJlydNfVcOgWOdY9KT/Bkj2poYhg6Pk1731hnxxiWt/TxW1Ch
HmtZXEOdrRRABraj7ufEPfAiuT+iY85ElY0XDFM5kBSxfXJfeoOHhSdW3wlu5F2s/5B/gukJ1GnD
A2/9/4iAWjCpxFwB7DK89zTJ5o0zXVziF8MWgDRv3KDDXHzEpVd/GOdl/OK/+5/1Dt//5WN1bgjs
PkPnFnQZlb2MOOtpNNM8AmScwW8aTZFtahXKDH9yPSXS1N6HwL7oXnVXWpUlpbqCCrdaiEBdZ4OZ
CESVWApKE15j72RpOBWz/1iGTww8vgJR6tfi5kgVmR9mNJ9LpGKaJofpuS0fYnDdYn03C4CjENzP
nqu2Hr5726X38ZeZM0gMifaCsFWx5Wb7fn9fC2GcIkLtUQhWIKZxMWbNuSQLT4i0eVuGJDU4kkwV
Bfp198RhbhsJciET81Vykk2gTCAByw+eQ1We0TawRp0cTIBFGzwTJ5zH6mRuQzzh4IJ3RtR1dcya
gU0N6IrXqDT92elWHIvqd0xdHAyXtZtjTY2ywRrw96ZNOahnhWRy60uRbQGm7eRcN31Vb8cub/zA
DIyk4iRmWrnROPp/1dlOr5kh2u9lA1sTJbeyRwQRiQPOmfhpCusw2q8PzrzXE6n1wy/rK4XPZxzW
tltLbyXFbE842mUUcPVSF8n7L6FMatqRW3zsv+TllPXweX2/XOCHA2nP2TCdzX1UAknZUSgs5ige
Whr9tI8dHPtaVJcGZjwlElbnVYCEeeAZqzksy8uLzK1YR7mvQzlEj9c6+Kb6lvJfbYQDwEaL6kO/
SFFmlwK45PnHAX6XF9JB2GSXreIuLugRtLcFb5pBiFBYpWMrJpWHJZL7coPTcKcFo0vm7it+vTob
EZDNM0FmCSIpRmvXE1NOAXdAjbLg42v+MNThSNMwiLr4ngTTFX91R+Vzq58g+WNb0vCWdg5bm3+i
rGIBsbAmPc29KkmfIPlzYvj9+yVzquFpXVYWVoAeNrfS+dawuP3JRFy4T4QU/KKoV1+GPiIkSpfB
CDTNAdhu3Hc1Xnm4ePjgGSF3Jo3rNr4RD4hEeB1cuWvHEunCdQp3eM9z0w6e/9GgcaDgEP/jocMx
tDH0KsL/h7X6D9r9xvh4AARJ4aH5UfOO/MrCPnMmcHOTS3tz4kUUwTohrUDSEf75meNZkI56JnQg
+to0rX/pGbYA5PyXDgL9WMpcFSOw7HMW2CAl4NjK0san2P/OGd5/m5NCD3Wvm7qkTL0FBHNxMLOE
XCy3p4CUiVP4hcHdzP6pcc5erb/G5MsWgbGmtqd4DcMLltJirVxtZ4zbutc98yNKdwyMzs14c1AR
s+UDY6+S6L9QefGe9qFkJrs2IsVapaXfA9JCXPx8T0dJzOYY+B/DivFF7L3vgsK9xCrLRktqPZEX
F3w/m7/ds6CzpdS8jw7ob1xJYURPZxw7ooN9jYi2QKUZOytJfHruALNRptuVEgIbHdQzs5OHLE+F
nkLlD/9LMd4gCNB5ns42id0fXj0eRsldEElMo5X2C6zCCOrtaJxIh96yR3gfXy0dfJdKJI5LWpbn
VdlQMBHpQcm1eOfGuQKqj04VXWAWUgo1k+w4WZf1HAPxA0kpC7s7jRZW339eN+slPYHCahRzqFph
rS8H33WEWzfd4GyMuH4eseUDW5B4guTW2pPUXuvoVRymGthfoXZQFSUs3uy+2DNmrHsY7Xkd0FRH
H7NSYzRiSTo2TzecSSieAS9mMbRp5RWjQcDrrhrMFCr6LYdYgNLKq8nIBKeAytnLXTbLQRjj22lq
2zHBOVZv770gLSpT5HPAT4zXDRy2cq392zlyrQni6X8i2q+prjcXZaMVaTzwh9c4yUm4f6ldAOfg
9oJVlDWn+xV1Rr1/ah1St8tjzCAFI3wICZmXpnYhnHlDOV1yq5HNESChlwZ10OTlJJQvO8G82Ch7
jew2HkXlw4HpCQp8vEPHBvvQNXRTgKRpLCOCYNa6GbKmWg0JUUVnMKORB622z1NAdGlVxSBSs5Gc
3W+qXXEx8e14TAZGWqOVMleXZkBWgfNnP39mOch97ud+d1kEZH5rnEGHS0ywaz3SZrVgVBm3D/5B
khKMwNySo/OHzeuXpZJvCjhnx9uJiirZjHsjxGD1va5WDXjwFTDG3yu8PaFqRhaxEEtM9Hgb5+G5
8+JSYrdQvLpi0xhtdXIWUmZ/g8bLu1T55PBtP8QGYFhb7WQRdt0QMQGDK06e1ChU70J2Msa8w8na
VyPhIQ29xkJ64I76By0IYbbNed5J2ZQMmtNhPkjI+11sqQElVx+UHaTQdbPCQeQ2yf5y1LycGJu8
KqoCe3nMuSOnpLwiJonINmyragoFsF3Vuegzi6SfL2QjHhNwA3I9iIpxTDnwdtFvidGQWxtcZ2nj
iFcnIcYgrbaexOGBriKYeLY9bRKQix3PPN13DBa2WNWtBuPbuM3VeEVLIf681FXqbqrDxb2vXq1f
desdNGmUfcIzPLUTMKKbhi7YbNCt81c50rS/Xnnwk2r6a8Gk9lgLBJnqQfEsMUN5Wz/7JOEys4Cl
gm5mWIBnxO34Xg0hfTzyt8Du5UbpUZU68PGGtKxVYfH9KA6Jyby2Yu0aXBxH/sBFQPhQWYM3TcD+
IdvexYbkDEnHP180LlfzAXmqGCOhVFkH4tU/yGuO72j9fD6PZOM0igj/5P5YMpG2sir9fbDwFtyy
MFT3MkSKEm01Ksva54FmpFWTo5v0za4SBWhcfONZ1wo5mFeIClFS2hmIqMSh4JD6wDLy/2vGrAI2
8ofEera0CsJMen6W6pf8yGiwvGM9bH/Tliz9389nr3xZzy7wcomX9br4hn2ToC4anHV2mBkVb9YQ
db2rYoNSYDphw9dB+c+pVM6nBPlBwUpslQ13QuC0tzdQKlXDT71XHqxARqIF44aY3PdhudH2sKet
G7+XSOsgdX0fFFMzcZOChl8Lbe3Kg6o205VB3PUA8I/hIvW7sueFHC3lMctsIHQvQ+MxCZjfR/ZB
rtYaUXTfDILRB0ex/rRON5NQ0tHGzJIxnLJf20s3LilcvzKXXjTUjNf0zqKukSQbQPHOdIUKUwG+
Cl9asXwZFAOLF545CCHGE125SHJ7fnwrlSwkaXpNstevZtPlfSeIcRNplOcaGfeAecZdxTeqSICo
yFmKPIc4sRCvSImPeeog9/g7jEbO5t/XBlOzwL6FOEOJEJASuvU6+jsbdLX9/TVFWzskwtjAnCGr
hYijDriq10Hfi08BMD4GLsTRA6Q1QjwytPJIBMiDSiXBilNDOMIXAgpXxLbNo815l8S4JYu9WQHx
ukREdHFJq5oolyapxGpqBJYYLZeFWxX7yW+ITsLTkB45ebsJl8+zKgmaQdgjDePH1xdn1DHFZUC2
OEzE2jLzBRks1R1G0No3IEII7DAlPVnu4AzQHlR0jEcflt7+3NiIxHRtdd9JTMPbbX06Enl3rFnK
z0xjrJkEnb5f5Db7dGJ0gUixA5z+yEC+K+Y4RYpm8c9a9lydBVlARRF6zdLQLFPJY0fAlJfnYeqL
rzl6fzkxUDF44KUotFE0VZ5n7c4984jan2a+bGF/UO4Y/f0nExm7vlIrtRiXvwrFVAcZqYCp+tXI
iV/o9U0YUV5QAAQpNfTk+mspOil4YM6HXIR/nqQQiNNh2Cmpeqt31723+p56bRSc2+ZHDErOU2Cr
dCGZTqRCv/8lDadrlc1SXHEbcDwTBOTRbJJYCYum9VsPAYD6+vb3UZZA+0XCbSCE8Mi9gQ9iBT0H
BDg1nuo4J3qkoW20gMLmTTqzKMdv2e5F0iY7sUIYXyxDlwbCksnHYCMeBfxFezvy9xUYDFPJWrSo
YJzUl15t3TQQ1FomGUAMc+hzMamKHLOEmsqj/Tj1ueFpbVP/MrTuDoBn9c7/QccOflTWJe+sVgT8
NqF1eRrf9WgYUUxKUq8mBgesRMDWQeHVjuNy1CUqLWUtloIG8NYdwzBW/dE+tinqnOrct0/cdT4t
ofUzjUxf/C5Oa7xM2lgNozDcr9BxK47pZGsSVwWykftY5KPEHvjP4UQdUPFXv6nHYNufDsloJhmU
Y0R+dVW+bplpZ/q6cC3vZ6E2TZBU8PpQrgo/VscZInEVLkIqww/C0YAzct3duF3S2n+rlAR5ZPy1
xZbdFoAHI2I476hqOdl6KDum0bIp/RhXJlAy0ZFv1IxzAuNv2CcEyRSkIo7IW7WOGcSwPDdGLa6Q
PAqkfOMMgDgDQQ/biH4jvwNGm3a6f4c69NJQH8PgHgXSgbTo8bEONHj0BSSQPSngtV8DHSm+nPHj
xTiVQ2T700/huGp0j5wIkg73matfTWj9Dh0vE10JmiOGuIcoTkolOrFIUTDo7xsEH8CjQxIDV586
nZuAcJ38O8hq9RNDSXlR7bI9w/93C9uaCmxED+nQK8VposhTn0Ks3AZzf9XEpiZDoSrG5z4pPkI1
MkHMk2kzrOsn4lB7wL0GUjZ3ezSxyHLa2uOT3gDLEVT4mQpWGJdo8QQmCkQaUqMsGbNs8CSt20B9
yq0gKlnXzK1oeD44FAhWbHArWGaBK8RouAP1q+0rNG3mSNxtwpSJbc6GkNoG+EO7bfA2iykFIRVX
nBA5SjEaQy2H21Cxv4PgBBo+yyxy2k3wAhz3hOQLOQiakbMEh1dWGla0KI6PPwS58zIZcnESUiDv
NgwFpWBrrqjWBF1VDiuVDyDNvzBTW1h6XOIDzOGZuP4+MLsfine9KNe0GM4fkO/va5BsB57qKPjZ
wCbmjrbbLrNcuWtQR6rNROaTHBiTYf/F75Usg5oYGDOCxXwhqp7Ia6e49rKk6OasmbORn8gdsZ0/
0pkvJ6msAlnaFfr/S/yVRomwKhJw87Y5sW9yLvtkj0K31RGxP+UC9RYuQb2n9bbUhkWgVLOm6ru4
mm6kdW4moygaAey21a6f47NlmFpO4QcgEg4Zjg2sf5M4nU9+YdSO+SzGwsft1gWZCT39NO8h9H2J
NTYPgWrge01/D1RBBiIu2na8XwKeIJx5NtrQ58CWJUJ8xlgWBcpDarvTvIQjYTFtgEBtaV1gUyki
ImXuUVcpVQLb6g5DrVizm50N4pI0v9WYVmhjLpPPQItSmsxN3gAzOZbmYxjmBSt3ui+MsPQI4K26
Spgp/pPrQXbcDiS/mwV89/7HDGZ7ctLHSwFzGhBmcVAlJGdozqUoBGOFF492EHqYLrTvpgyGkunw
Su+tsCQChhHzo+o5lBvjTg+BI8f2vlpYazKw2PHAfXfuT9x2InZGIFka+MYFVzRJdCp2O8Vcm7ER
iLFPgz5R4o7ZLKaJmKa7492hYXxwp8rLqOdba5BIfnyKjZEf06twF/wtWjYwqpPAow4HgtIEnBTk
kpa0i05wBiXxNpk5P2Kkw2/Dk5MT5AF0TRkFHWvVs/Y2Nns83AdVIiIIK08eAvjkNfNt3hP3cWoB
OLa2s1vx7PYT3OpYphc8B8MuEVbsfthSxmS6+CMsRXfRkAY5++N7OCupIS3N/2ZG4XXpbPjwi3jD
YeyI7O7Qyr5ONsGhf2ZvD1Mu+RhDG8wb9co1OpAjCSABZh1l44JFC62U4W9SmyI14eZQQpnya/hs
4K2GaI0T1vOfFJRT5qxcg6M7qe0Y0reVwf3zNIDQoyy3spzU/m7qV2sZkL2BmM/xAYDjv+Dy5ENW
4TR/N6f/AONe+O2QOzpTSeHNN2SxG6lpV7g5tlI7i2vqKBOKO0sz+hEp2zCwX3prHdK57iH4wVzg
a8vsWpEtCxs0aIwFaQw6fR0OHyxlCekImjqWjFsDfp+p9HSKRI2y8mdwIw9XA19xPLTfWWiK/bbG
Tc1/7Sksm7e7k96nQLkZM5vmqi8rQdaJm9Kfc1RPkmkUKXN8WuW9sZ3Faib4V4z4ZQzEq66A5WKy
xqd5gYcEJ844DTHC8q/GlBESdkaFdLrUGdQlX2+821thavHRgFTIxL/sJ04dtpqE6SlcsAQzozcb
ljGBAZJYca+kJDdcoU4X6dJMuNXRzvQf9YKHCSL3YWM5SrshXLUPmm3qe1iKdIj8tTE5N/n4dteq
jOG7z4PXu/eSuVlsynRk9DJa+6w45C39QD2bC771SYABpG3iXnnNx6baKdB/NYN2hDnaaHdppDAt
zQS1DWxoAAFNjJp6uSKFnfKxcBO1T758CUem0tPyXFHLOhQ1LiH9y1+qnH/JBxiePmQxwqYx6Y8C
zvwaera35igaUkK6Ge3CugzCSKPcAToBQeuFEburcKbRoXYYpodKElIxXJd/+KnNQifCLSuFZdAD
K73JbgmUHfb7+L6rFtT0wVtfKA/lRMX6sDudeu0Ye/x3CmRWbSKmOCvoNXak23jMlKRUwj03am6h
atO3lsdUzgiMShncR0y80dIX6EZPyoyEpSZQ86oug1wuj1fBAjHxttMH5vgvXCQ/N88cTwsdGzxR
ZNSYsiTUARSiGSvg4sHLP2MuHmP5aYQnujb0/NVHBzlEzWjemc/bFOJ6JIztDp4neMvySQiSG8z6
BgZIKO02j/3CYv3cLViLuoMwPl2hyi9JFgYwWN5R24B3QRyvsUWK/21AWPWv46lNMfbvy5WdmtKh
Uqqk1YWf4ywsTYoNmk0s3OG+JhIxbvSHuvo3X5LYBk2nG8C6tOHAcajIG/uWJGc/DKLmCI3RjgLD
f9DarXPASzIeLsYLGeCs/GMU8SqMyDGXGm1XAD5BgOythwM1dVCdO/ry2t12hVlOpXAcPqpSvn1R
vrMWs6qmx/B0u7XgwF2rO9e+aOU0XGr/f5MdJ8PhokU5fGQv2wgK4t0DVZaErlGuf/p7CTWokR5c
vnG8v94/S6PfZwuuFT4DPrdXTpGKnLiZRzsiYJO6RIiiYSUkUaR5LwEDVMKrhoxcohcZ6/DGGSgO
TlbPgvy/bAsYB0wA2zUbtSRHWI8NV9OD9HLkmvW6wrvtvgTKZUXX9KWydvHMD+VL+2D0TGBHntn1
Eb0c7wYkrfxsXZ4XyO2regLqppVdXnmXE67ExuArkxuAcqFAN68q7Nju9WqPf9nxWGBv3/w7gRHM
N7I45eFFTVn45CBxIDVO9rVcKNXov6fZc1i7j0swHXnkE6sJ+M3gu0FFcxIkCo3uT/KQPR3FfHZs
aPJCCtJm9DT5LAXJGPuU8KUJLIz9Ys8iSXfVtkQ4uXJQ6Nf5hIUvy4yFnl5wqlF5TD6eamQtoeeX
ehylISi1Bmdl3NzTRGKAD0BtIyRUQTWjvGpoKusCWYgP2KSyCn4LLVmZ52XmrqqMofJKFS4ammLi
N69KqnL78sk7fxT6vzPVFDre28gi5mkfNRiZmnrHxzx6OTtGbJVm/HPg/etG/CZvvUjMfQwZ06PQ
0sKD9ReHCzpizFSgWEdqSwCqMpZhxsjmuM0J+rh373rivDVM/z0RRDgGd4gCBMnWsYhcM9r6edCk
xveUhPq4lI+7wDSM5TBbpGwZ2ihEb3sR50i+rURSqRzZlta8nm2FFs0GDH/VZNF5spuVDFxd7grR
8eRD+rtB00hYzyRJuGyoLhsYznKWD90YVUBrTI1G9gPgBwRDCcrZUISCQZ5LjOFhD3QfkPtlVsej
y3Vjb0OoDAIZZych61mC+y127fV82lfe+7yejH5nL5a7xd92lUuPDPsBjDpkfdY7Wo1DNCdJ6ons
xixxklRVhfLAwRbWqYeZMg4dmY+NPnDmtQV8nr1yaLiL0TNbfeWMWyUgwYrqnMX9PmIWP2tfB9JX
cH/B4AfqDyDGDD/XGOW+xPLFIPxfvCrEhg2YN4YnQQVNFLuhrNlkREYe5/QpoWKJWnYl3R+5iw65
TAqv7uRi3BmBUP2pcqRC4aW72E0NC23QqhK/siXWQBWP5NhFecjAhDDCYbbPqqVc1d0M7k4eP7J/
84T8nP335+ii2ZpO84B9S9ZoHmWxIs8pwcHZf9g44zlkblUS9TI4PemfMFvkJhm5Qv5J0t4wdzXM
TM7fbTVRM7dLJ8rgfI341+6JogDzCfy/puIrYa+8FBkLKETgNvNJdf6ZCCeuRaomq36JN6EDBeB+
4mycqgpoYc1c6DWBN1dHVRHUHoBeYv6fyzLY+qHnxencVdg6TohE5ZpKd71d29HnxMaHhCmlh3h9
LfzOqQ==
`protect end_protected

