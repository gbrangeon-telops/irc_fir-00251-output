

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XoDvqNcsUAMVrCepxGZ+692mBkX+rCE8HMYzKPm5R78cJ+RMc0dkNWWZsdClXOY6y1T5UuLnfOdJ
4pIk+MIfbA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GQd6VykDj7htiYnOl+4WVHQM4hKgz1J8Md5aI6kr8/Lamm+PnYCv/9ATHhzH1x3ZwU/+Hk75nShM
Z/fTah2o7SNlXBmxO/TZV+Cu1NdyZPM9aMjSfxhjbc4DdKhbt2eR/JXlXgPN+qqN+l8aDRz6dW1r
rhTiAjUos5V3YtoS0kE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1H8fvXKZG1QF+UJtGmRK0CnD8bm/+01l6RcgU14qYFFE8GVuJpGQyW5h972p3ANLjy1WRtjYQ4xM
/dkbNa4PXjLXaYaHj221vfSd3lB0MAvfi3uUVJSvclNp9cIhjsynHt6eX7sY3mGpxNDMKipfks7Y
7QsvE6SpbzMkIaxn/W/Og06vrJaRobnXPbk5O8bulSLgRIfqtOFawh2LDbI1+cySFds9EMjhPXGY
R3cSwZrw9voRIz0AJIAvvOBrLoxc5eVp/j0gskNHjRbPo5Gkm/B0oz1Ia6kiZiwtS5XXf5fYsvSq
8ip/JtlfeTs2FRpXweWaPr5rFOg0LxkGg0mLCA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7F7hPxr1ObCyOsY3iC3Phcz4OOcedLcCp9ggSn92l+/8vc/8WokvA1XgYsChaRHJl3lXf2X6jfk
OU2I7E3QgZVgyd5+syjWVqouw27C41FFBeCuGD1GtzyBYnFEqdtK4Wi9fPab76EJM+QSrUTFTxOM
vNsxaERzJOCdVgQoGH4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DAf8RFZxkL4Com/8UijiDJflLxIdfhDldD1zcH1XeixMo5g8/n+Yg5p6ecx6wthzScLrbvkfxjSo
INrqjZhuOy8JD1hgSySspkuAnlB/pYzsB41QYrTQXDdhODLQLAYA4QNlYnc0Hld5QRA0QsNa7b9I
jitn7EoP2gA5KtAm5w8Y3SJ5GziR/wWC7+Oq7vo7hHrOsipiX4kUa9vhXNaEzGvrcPOJN0YgaqRR
HJt/OxiJdqU+tEWkUefOFMVnQWevf91iZ/Fb0oG88z41wfeJt8eTwCR6ZrUTPInU5uj9Frdns/GT
RmMrsalABVuwLraRXdip/IKnMD1dw9K3eH9MHA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94464)
`protect data_block
+Bqc2FxN4HV0GKO/myF4lee9M8YOFpQpApZwXnmhUDOBLH3IG45lmVjItf8fl4smrPCn+u1eWNuJ
w70Mio0Rvp2nKnHPkwuOClMGWhbbgB38VO7bqQgJqWh+tarcgQtNz2yQyEwNmG/H2zrJLT/5iXQu
6iVbND79wK9LvE+mHBDsMwjJ6eHQrdfBE2O3hyzY8McuNYbsuhIk9AHf/y9s4ZGG+i0Qi0QM8Vlq
w7RXS+d3L9Df1bxFRG6LVBChAMUGpeQYohpB5Ylq0q3hxqsuZ1NAAr4DSp3Fffc/AJs2W8useXM8
yTq+mM/9CwVjNy+oh07zTHb99RA5WB3RvVV9nd+UPvsL2+0P3VpYhOlvUwDpCuP+ka2g/73VE7WL
C4UIJcVsxqSs/ijHhtMfKmJKALsNxsQIcf9DMBCG8uhFXA2dPHaD0loA2pEwFOfLxp73lfp0LJUE
ooaXFc5BX9nxv4AdXg1lW4Zk+AKyJJ10HdBSGtlSR5HyiVAU8aj2mEm0GcYehSsZPkGFoTAIV3Cj
XbnK/pGFDfnoqfEi9QCIG2H9eViWv6tXo8mwN5RA4YvJdTTNbkUVu2V01/39j4QmUalS48a1B5Cd
mmlPG9K7Ow6VgSvw+geMvXfcfj0Nv+4EUxpsAc/uVUx5hR958xbM89P5yd388vf4kSsJV4dVahs9
AA5OBEAy8KExUnpQ1cSg8xtK1F3uqOLnVfCoiuZwWu6AHFCOdPC/p6GJw9EHTWu0S1BOvqgq2tG3
QSvwVjClnM87RDbXzlpzzMtgq3usMM3WYJ8RnM7wuUBrZz0mnUAqvIzZymFbIrQPmd1+O5l2V1ot
bTshlhWsDq7c3PLOKbFcAx1icAZIy6Xzg0rPyZHkCW+GQqboCgp0d0n/RPspJ62bBAPpr6jXZ0aj
iUKDWTeFSyrXsjoGbZmavpYL4nwdGmrS2RSVLNqJhP2tHJS0X1j1jzTsDE3mPcgdnpfXLFQVSPBa
LJv586JrraQpKYoZkMgDZCxHUVCX2VG57ZNOkdlC7Y67vzWWMvBys3A96yV2oQJN3DBKJDKCpFwo
djV7S9WszXBDHb8Oe+SutCfN4wVixeOj9p4KJIxxOLrQmUwWqomAkdaxqsaxPh0jJWJUDn93T9f2
jYmgmxMIg+5nbgizhx7h2PBQuDh5qciaeJHQu9kBx7C7+VhNySBBqckeJaWfnip+n4ZLXU5jNio/
cgrfb0CEvcNpfQb7Ze4iD5hMfjx0ISc1iXI7OMAaCivw9gJt95CV3sytsotlaIYWnvCsqKG7R+lI
63dgf5Z9s9+66IFXBIZocCScjy7yL6G3AhrpdzQLXIshSEdC77GOCY5FRhHkIemqeykmyEMSezQv
xq3DuXPtIbVrcw/UXHPQbRKW18UZZ+pfXgiQVzMcITIdAezRCDXQjSKYmz+3z+QmamsG99wL/Q1Q
Sz0iIv/5E1Wgq6FxWZrbJUfQaAQS9b8nQfW813irt0qte1E7rKWVhkzQbAJ79siiOI/gJM1KBBJX
ORiYlBjBkeiWzHYnt26Xaxfg5+KYQ5pQVhIoVC+ZiQjm0MfkLkrMeNAVXaHNV21I5eg5G3iZxLGM
DTLDTSUYeGaUt6tkWP33PIDgpEBmqMGfJLXc4NmQskxn3z3hUgfi1uePzeXHttZ8VH39EidOfaAQ
24/T1p8Ye5qOTEEQ4f5ZpPoNEdY7hmiioFQ4seTT2Z5OTYnMhoSE0d635a1D4ZaPszcHn+Drr4vT
nW9Cn1p7fS0fIeJGjiLTqUijNU+XeBhrxbH/nSOeZz0y/G0zkfgDyrSTVzaTckafIlcYKxcc7XzV
Uxupjjc4izuzw/P6D+diaAhwmvYvfnCRLpIeS0BDeDhn6rE/mqwthfFMNLLkbIlg7JyGiT/eSUrQ
ymWsa4yKex9zg6z84C0ZPXgILEpGMGSohKdHOrJBKVQDhDMZKT9pmALTcFD4MSgUx8+Y3mdC4J2x
LhiDI9TiF/TCRQif3ehGXv7VQlndkkJVTjOZs2Nu0xqQqnng5fiMDhB9tJp5VM60cu3OJG6LoOPv
uvm5sNDzRvtLBrvxaMwaQ74gazGinfzo7VUab1k2WCtpz5YDHg/qjqxzYjDw6shM9mboxgCdxCX+
69rKZFMrgg5YCwrKgUeVAdhUTDons65jwmrZyWrUZ5FzkvT9WS27A5u7krCZAJ9qUhOYMKNOEsQ7
TQCLTNji+a2kMizkLAAH7P80ZCIIBV56Ur3g+T1ATwVw9fICuHgy93MRA3rE+O3ezJ5G9sbU2VLf
HjdLi4ZEDkxtFh2gssWoGTjjjX5pysDjm3eQ2RVuPOfcdV0Fcqn5+Rc7VR+gx4xqUk1k095MyhWp
XS1WB0Gkp+6NzmD31JEpCtj7jIt6Gsvwo8/dc2I3gIGB7dDTAgh/Nla0v+N3HAGOF5cH9fIkmzb6
U/cwZxnazz4upG8UQ0BGe7wtpcISJecexSK2FHFn6ezPkxA9srHBpN+n12QQWnCLaJJ+N8XxYtEL
ausDe24T83eywCnxapaEh9c8w4Ka4XUNz1K6gjKNcXQr9BE5+poBwaghDgpBlrg2ZlMVHDE3XitY
Mo03ESjvKxEe2BYZcp2txtcuhjayz1HsWDIeYV5MOtuYxghdXc99l8ZdLypTBIzecI9+HQQD8DFV
ZTNc/BkpG9FBUG3BnkY8OMmIz6rPB3mCqafGHtJ8tREWeogyHiE8Lk2hl55KjJNHeSm590X/ovo7
gsNFHnfaP9UohTg+Cj4R332mwJcg2vl+hVRu7vdDetuAxrDyFh7sprcD/hR84UjyKysH09hcUG86
a1rX2+ySNoGoKTXaxW+A8ZkSHxPTkhadIHjqc8AjEuETLtAylzSW0AOZtFxJRErOLAXT5p3S/n0E
IxOBH9nGu9PTsrYPqku0avuA8BujRTq16UodQiAvegFoaxa6u6B655r+X//QLmuwvFv1LpDyH9J4
ksy2ZpN0sXEmhmDDXH77XfszDsoNMrH2x1+sFGt9Mt37Nx7WZClInkVNtI3LFmhyzRjsszU7z1qd
OBTiI2oEAPPFxWSWpUVAwlzTszhbnm2REnKIFbPVI3ML1OtfBWcqCcPknWlHdkREYdeyk3wX7EjZ
hxAzyDp0BC/m4jf2oKa0JkunQ280gEwrmMhl+s9bCAcjNfj3CI0zGyocuvsj8+g/5Ojxc5/FonMN
e87QrldieWm9ph1eFAjiq5cNRsx+c94PPC8jeIXTplIdw4Zgd6rD3BVhh28AWZqOT9hlKMAVEvyj
FXuknGdkDl3AF1CvGnJ+R24EgzziXE4rfyZ1fFXFoypX4mUJDQehqYGdFifu/SWFOql9bw7IqML9
D6lseIMye/klcPxmDovxTm3T7rtqPYO4Gu9zX54ap380VQ/OhJCoDfGhChuVMW0+s4UU1G6EBvjh
Li2Ac9G104UFcMs8qBph4DyKeQVbTmBBiY3Y9ANC9yNT2kH/hxKrB/BCtYxzeRnwmE4EubdpMI56
A3eIDLvTSrQQPjGUjqU7Q71SFmjN3aO1lE572QvawIqWHfRuyN9HYV/mTFvqDcJXG9RJd/z4kIe8
zbd8COCmzA4DLspWZKtEA3EHFiNXgvJZmLouH6F09bA8DE7a2Pe6ZjLQbNwvCXCkzzQdnaCpWtRo
2Y3jdeEB7lXFIDwHWubb8K0UFzRLH295V9Aht6bX7Ci70EPmc/4uDhyIvD4pPYUvXnbZKK2QUax4
cePzz+ZliRSf5tpp79kc8HlGq1RPOeVCDn49icUvqH03QKMJKF9V3xgyXvu+zKUW6YTT3bUvkpYC
iMqz2ndFryUcRNF6ugLw9rmhVoYEPCQcLBudud8rvVRotN/ZOT/Es1WabD4ylZ5HATP+K6pfXuSo
AhMyGVlDyDS+qtG2E7JyQIKkLd3MbdDsbAzL/P153IyazTMKbJT7wfEuhcYRo9shjo0/V1IW0NFt
6eoIgqbyxQWsf3Mvzkm2mWtLNCh++yg/+GP870+v9M+ngnMPusHD4egCylRjZwPBF373ntLdOwQ/
HFegkA2+4TxcR/IQE8cOK06+P8RuSSdo5ajrT3MYV9EvEmPYBANJRE8NyIZOtlRgGLwiloMUrx/r
Xt6FdO79pB2sRYBIhTJBpyzJRynusnR3qFcVvivlTSOO8Jq6VRqIGn4VMU3qJ+YuV2BboNsS2bXS
VcJ9070qtcQKmM/7pC7VhRMOQZgynJQBzzEeN1IUD4e8jsBY+IvMZPbEa1B8l0VXXuvbAIQyD5rz
aHgKxuQvC6QRHBLpmYgQeRT4z7VGdcY2pywaiTZZt7Dw1hrIyFFOPXcMpz59GE/bZsgn8FTWXwmp
hE/s0j9U+mQshqFOFT7KrTH0/cDEJbMEiGIgfPzHkNd+B1xt3e6smCqhQoUMkwHpA+YD1fO68cUV
luuNo3W6hpIjqENoFR0CCXHEHskRJ7mrJE0DI25jFpeVn+HE+d2+ztE/IVOPB23B1akZxnLmbyqC
RBKlzUbQbKhFw/CK3MX/lXrKf+RR0nzWy0HPE1wsyu/6H/UoyCf7/+dMV1ME3lxYYxg3rHvmtMkF
hIjLOPYWuxkJxcPmY/NXV/GzoPqevH5oM1GQFSwgBXvatc5Us9gB+7DXdMAxhlvcj5MVe/+1ySM0
eB1v5Jt0HjJ1UUAkhP4ZMsrW3h38EoIPMqgFYfVXjSUVh81RJ0OZXuISHIZxayrHl9QzEyndiMkd
UWLYmjYNNuWe6UlrZu21JMb7zvW84EIdPOsnJdAl0FILY4+E9IcNOSD+4/9nf1WD8pGhBCSXiIEg
Z+Uf4hvtpNuibM4XZekz22vKHY8EXVcrLGRvICO1cU31mwgeARnYeTYSbF9k4/KL2q7uKtNl+9EX
76rDLUZeoXlYi5vPV1pYYTXe57v+7R69V+HroS5eJ580kCKOXIztT+xps3IF+ge+ewHj+xXGw2EF
wja1mYNNW9s0n1SeruLJIDifguBed0o1zsn9cugp1jUZSaokJXK+BFOLPCtAkRIM+aR8M7JcCACS
lfj01k41EonrYlk3mrB6rR7F2h6Rm/EBBNGk2BFnYNaC7v4XoQZfK3CXd48vuenvi955IgxAmifR
tcLbZgjNjrDLSA48ktAU5yEmmSwYn8k3P+rFLU3lUdy0lppApqJfr3MnaaPRcuKnGMkWA62a8rdu
fTKC2aYjPfnJ3qL+P/3hpgkjS746YjZPGM3B/e75sGt2R/M492e5yhKj1lZjupNamK19LFLv4KFl
ojCSqjnMYIGVfj1vflmjjlUbW0q4JmKipgxg3mpYsHK2tOHVwfUC3MROXAeIPzXFghVW0FuLaZlH
GcctM1zWDR+j1MsZeQikEP3TNICMYgiG1Pa0/JLLZDs39gbrAoL64J8wfjWPzNdSHCyFAKGaiEIR
q931gYiO2y0ZDZL7+jC70CnIK9lFh/8R8aFal5N1F5YBpZkHcX6se1F1XhwN0c+lwTkLNtjM/4zD
B0RHZzSK1BR/GL2e35J1DjFOB0L/R9zeCgOqwdHt6w9w+sOU4OFhneme+Rk34iob6D+XhDO8pwh4
fxGzieMNMOHESeD/8X3MN5H2nN3nIPGy7tVCkRvGj7r/Br+B0wbZyxtRh8eZ8broZgAG3Hq6+9dr
H+ULrAdr7cVJV+OBJ7K+/YgxIfwcFwAu98DD13vo7X92dMz4OWWSkqtwuybIiKSA5OYgfCzgFcP2
PW2cHOP5VmiYWLKlfluOaIIi5wk2uB0QAbC81MNorcIwyMxnAFx/O4TdnTVAnom3/htCTUywSOGF
9FwZIwcbxS8OxjbNxbC6K0QXyCVexlP9kU0kMLa6rYXQoxY20AH8idYf1yO96AnkKZarM933PoY2
V+SGao+KWML0AScNjlcmFNGP8wU6rxK9vix6sZgyPGHWM3p9Xt6N8JTGwTMj2A10dmVjgQu0axYi
PZuTbQFQcSoCO6vnxOiIwUimWtd4E3UqyXdWihpMr9A/WdrEvN64knptAjEFGX0bYaoGQZacRB4w
uROoTtrW1oLksZZA8JAUanGs164YlKilThrpPUaGUl3ipUypmEG6L+N8Q5rUe424DqQKzg7mpgY8
gGHzN1uslfanVBpq0kxXZu0tp2iL1nDW9KuhVZDV784Fygas1KEJan7rzz7VnPWS+ZUvc30L5BmC
ekm+AhJNhZc/sf+kvZP+ajIvTpB7fgk/y0C8ln4c7nZcsseFWL7GNcIYQElChsUGK9PKK3G5Z+X/
ji3HoOg7zgb9jT7T9bWVRSBcsrqeRPfyMJ3feT+xWum8rxGSSSxhvH3m1uYBytIIU1NuwiZOf+CL
aNEjN4BEJGYfEWVO8Obf0JWsY0sL1iQefXoktDRmjdcYkTeOiNjqhUhmgwt7gbUV0XE/zRrSpnPg
4kVt93QNvEAzy9bxSXYNl8baE0ifLf5iF3rhZTFt2+5sbmA4VbV7nfgarYisu5sAfQCyuZPMia+o
XjKXaJ+XIFP+e2tvpetew95gmoa5l2LhTxKRjUzMYEj5bPNTXGuiTQ5hox4Qi5ftGEdCF+kcUTXb
PZVzkq3I+TI57UZeVXI2SE68e8ZwyMrERLAxZg8UmNWp65DH/HSUTgvWoluHUsSmqLCj7z7MMj4u
7CXDAppQtNiOVrYqdU26vD7gCl80hm6AZBFb8T18RqRgdCtacTw9I4WaAaXnAC5mVRwcJFDvC/3q
nbvvmLFI00YGvB3FiA/WBzFT1KRW/eVpdRPUxzKwX+kfixkvyyl89D93fJ78XwHl2DGFW4hjdGLQ
CzFg0sHvRY05LkqRjaOE+DwkgvWy2JFjj34pfheLa+WayMw+lEJLIq9a5UR2CvZ26cYe89pqTLXE
hGq4BniW+f/+Re+cScZAlNRUSFPkwJy5V9uPD8iU/aK6gXaFRNU3UQrXg1bhhaHf/XhTD8MwoHNw
KB4fM4SridpjgvocElLUAFpMGVuWsvbtfVAl4rU2AjIX3ntZPYnq8gxkoQp+ZEqcjeGQwe2Hn59r
jnFMPnCfJVDhrPGTdu1GWdwwj04VNwZ55aqPgOCI2Mv1ghGi2k3ZpPMWYcIFcbftQj5oWE5TX7v5
NlOmUjr8Psoj3S8997bD85V+GjUKWj5bd16ZyFMKCJP+Nbz8Yy1mfxEDs52YnD7sA+vO9WqmJ2+J
IuL0SXJ+xus4WNoq8fA7NuHDBtQS1eFEhHWA5nK/zlIpVnL8J6Ux6X2W4hxkeRthW1hbC9TjgB+a
a1rdyirPOvJvL4CuyxeN8VegOPxM4Dpw1bcgs8dMFUM3yUuvM0soNYe1+S8q+diggMIQgfYdt8Bv
QA/OEuSsvlPHNdsywFh0unYvs2dc8e1ES4lA96WP4m/OrVKYwEP/to6sgTQ+rnN/6BkNucBo7D0w
3dtK37SE4KONXtX82Qhd2VL4JtItAipZORtlTL0v0b9XSS71xsClg6qy404HfP8Ezpl48VQWuPmR
KqSH/OqHPBzk75IF2FruzfpP0LD8d7v8M5PIvNFwAoklf0htsGBILpBTPgk6RqJlhSYLVIzTSrte
8/J1SRhy0Ss/ToIkAgyilKfkFfCkd5EN+4ypGE6I/7GKattdvAiblUU24XvIFo0OnpU4CPer/4SE
oh5hM6g5KA+lJeLm8RjWT+WzSwX48gl8VVRgZ/kd7VDeMYbIfjj1Gj2uQB0djrU4b3ttp4Ay3mov
3O1GWlYZTKzRRB6uTOXG+QJx99XK33qhSzz9SECgzi1EXXxS3HwhYY72UMlXmQNLZisg22fLpPEQ
yyBtAKpnFkPu38GBaPwRm+JNoWFQcDkrf9OiAxLxCWX16nH4W9DOyQ5/9Og+Ne9gfWtRjFLBYZ/6
atZoOqt+fE6awwpSKw+/yWL25vKTDf/mqiOZ8qI4JFaKN4iWXkWsKfy/nrAol+LCDdEs1jfeQ9D4
zYQSS/ghqo6E9G864aAZt/7Uvq9vPuGzTqsetQZ4Dpu+WR+fAuAu4y261aF/UqimyOM++o4LEWue
WXWW9CEtizrjfF8BFROEJEymBnHoUpaMXbAXjeksoN/i1qR67WglmBoWNUaf0pQu4XoDqUn6cU8E
KO56JYJYDGjUGTtFO0G6tMCOaArhf3DKFHs16i2bbK/1Cbrmkx+m0Z20+fz+7BJf4xlAa6/RxGem
Ru/lefEG6gUHR/+ftRXT1NVQMUX5EOO45bT3DznIYXwwlPkvd7kZQZMnbwca9GFC4EIUHTJ4y95F
Kcyn46N0OucpDHzKhl+KcBy5zh9h6Z3UDzQxx4/ftfgS7Pv8iBbZLCF2rq0eaM28u2hkyd83e8Ue
sG8fXiTySjw2oVkIztyzCwJ/kowSRT3tI3dmIRT3pvvWdbch4YrhdkCnMg/s5AQDQ7doqvHlzYt4
IqSppDZs3DyGMItLu0ZAz9g8C/0zZ971LnVT+jByyDTug9eFJxzUChcr0yOQm/GEB40k/Eru65hr
kngpDNx9JK5JhNwUbEgqytXqAY/2H2SKGgZMWoZTZ0yKvHvoOs4KoqgNyEtKWjwffLNJQl6QNtMg
IkqdcKoHaWw6KS1WsVj6U5vcElxfFBZa6znklB/ohWldatw2oQq69PEqsAAWM1b401z7OM6O1nB7
mtWejAvpb4vM2RpUkUSkGd3KcKGZoUV7qI9kFtGMc1tZU8z5YPhH+ba41WOdXnZ3gxXoWkedBrX1
ncj4n9eIVWVYWQGE191Kn/tT6IAvedLte56DwijZPPYIWtAP+qqiA3+n+RHnsvXf7N4nq4jHZnL9
+NCR0xjawhZBCvHpJx/Spty7dwpblwC1P5ic+bkx9MQkB8MU1Gla3nFhwNEYhYXIC0BQmCj7tFLH
/vTfi1u/E9Smg2cumL96n6AcxWRH9W2798D2vXRWmNnS20sXi7NaGz9GWukIRrkpCegI03ogP3J0
2xhtNQGwwlRhh897qQCb3vvRsdFaqNEVHTxGKkA3WvXohx3yhzRMezFO4iJGCEsQhXkx/4BengCY
a3oiWx6/zgmwZg6aDSLnjieefcVweNA3LO4gf40LqLQuXB++aWiysFRBMBLcn7XACRlurGMPmgId
1Y4Thq+f2o/pKzOgU4iaj9VpacaDOOlnSWVSX9JtvSoMgnIGUkSjiRJ7EdWJrCju7Kr5iHyGLeBV
S1VZ0ewBMA1qVMabkfOivz+NVi23eyq2YG9oz0VzPgVcuqiAwn2Fk6tqhEjbZSJAsiN/4HHEbhmv
vrBWopkmG0MHXt61XJkr1FlUQhh/WmAUtFCIWj8ICjSmVnKXfyTy2jMk0J1ta0Tntd0XYT4iyS9Q
GrcTVz7+d7gZ5BUWcc6GAEpqzLC21eTD4Zt7NXnfEGuTNCK7Brf5LvMfz88X48My6Mb+JNKg19+L
NUNLJj6q0/KmpE3g0uHYZ8Rd+bWCcrUDMg02prdhpDLoXD+cIe1PY7olJiIIO2xkiPvzQTRFjt2Q
v4Gwt5AERSoVKnwYLGXW09eqGav/HsjcMk3vRck1OY5feeghwbmxo+UumEYiZ8LbGgeQpBu+FORC
58Y0W9Pot/rfB+Sc5I4Ne34jdAMxBTtSLLkiKbeG3XkZmhR6oBf307H0RmepGkiyQCKEvmMTDPKf
BLXyabd9Ib9epn3twoRWZMhSleb8W9y1NjPsge+CPyg5GVg+LrB7+S9ZnXTpC528TYiFj7zJtQXa
1xRnCeQDvSDUpNf3cv1yV8/tC4Hy9p6Ae6ZvH5YRJ/iy4n6fcllFHDLPhiYMm0QBkwTGhW4iNzlU
pMqlI6eSg+02AZjwQWrLrajxX8AMGa/nSNJWcNIRqUK18NvQae7Pl6/UHDPKZPFXnynOsUXaKjMQ
NNPBdVy739XvRQd6ACpNlhn89jaQxfOetBpDsjDK1YKWvMLiPdrPCjZCPAgftEdv1BTUmK/9sVhC
O8B5n/rmYULf2jQSaat7Ym3MoP1QIGbgSyJbrhGH7h0rNcxQxNF3vF7LwH/CC3CqlkwWsUxRdelC
oTAS7MbF/x52WlObhGuRe0hHk27uTUPwCsOA0K3WUFjD9bFameI/6cqekBlvtuAKLAQKbcbmHep8
ufAvXWSicOJGIOux4Kt6EvEev3rVv8dIo+TJQd/tHuGFeLX3uZEdK7B2Pmyl0KlZYHbNszc/anfZ
NivpCCvp2pELVuh1ybCf6lDeoQVDIkyvranKER9vPbnqI5pHtzf2pisQOVMTTzfENNFb+emI71lN
B9o1wJjCAWT0yyG4FAEXpWZQhmZJ/DukruaKbEfmX0gmlgS5E1F1dhzjvfDd43e5C3nngcB5a4Ra
bf7Zuo+Foxlmvf4XfQNE2anYgGpjjUYhJsZWuCSNigNrT9s1O8Shic4CgFXiaB9JQ06HjSa2mdW+
QTVCLJ0fp9QN9kosuCQ6e4lRv2pKZlYZDM4L0uiqkdsQyEq4S/f7RIKWKQESCBV/z54gSVqbLtG1
sfk6WXL63AVSivZ2041uCmVWfdIJIVi36KKKpvVExSQZ9qnUkiYvtHV+/pXoeVXmKoGi1WpqhOQv
BUYKg8o8nxzJ/tJBv8OeQrNMjAuzP2RFCygmLNm67aVttHVUOwnK89nRiv/oADs2+2/viYeoSGrW
Twc2DcsqiDOA6FVIrvbS0EUM9Bx1ItkMOV2g5RgeIyIiv7QbYhvwz59NGOy/Ay9B5ttc1Hp078/n
QEOLlkzq41J71yO8xuaKH+7qhVURavpORYU3KbI0CPy5rO3F/aTW65m3F2DwrgxNPjs1PyYFlhKM
CPI13Zvvn7YM4VK9qd11P2D6+Xxu4gfympbvQxt3UGbHvJT6NzJPqd4jl8tDb9BBDBpB9Pvu+lK1
mnjoFSSw6rMNMlMolHY11S4f1009pEa+Jx1rlubPnJWZEuO0H0mZFYVT5EXe1dCbEQvRj+eApNtW
YV4De/w6vKmnSkNbIIorpwFwH51wXcpHMxkZZCmP/9ZVAsMBKixdoCGvztiPhGjoeCzhskjvG72U
aQRq8ai/vJDyAAd0r3m1+4IM3QafYHph51QU3j4ER7Z940cgH0vXc8IHodEPmNGOaeyt2z65oRxg
CcJhtzYoQcHAVNGUbAGSTEFUZ38feMnXKzifX8UKojxP1nZfTvbwBrzkOBePlF4sE+EtsdqxNOFs
PiqDhcJrnQ0idoi60NqHEkyk7/o9HgghjWX6bH4raOFdHIMDUKRs1lAHpSR/mEbUobdDGbhD0vh+
ctlvNk5/Q6p+Kz9/t65dK7CskLEpzT+sxU3jHfPE/9gsaJ/ATOnX5msTcX0kxsa1GqUIOtqNqy4S
P8v0ZLVjZiARxBQ56RhaBVcEmJCpiSCUunqCRopEyfPXxlzsWi2xcW2fCxFV12EZXCP4wWTwt0G9
YL9qVQNeNH8Uiil7/HUKKIYsd3Izzpy2fx3L5Vl+jp2hTU66MkbgB+PPQDFirc2Uo6N7lb2w5/QV
rHRQvBa0u54+4tTMAv9I3Q8ihxIYk0+fEDiMtYXnPcrbEcGKtc+ALVQTyGBuPsV/eHdOGT3iSSwm
7QGkuvNVRlz137aTxQ7f2x3Go62hHh2EIzhND8vCYHCnhD7O8+RJPSkRUCpFisjejL888DbW7qlR
OefSOL7HfHATHw4x1O10LaLU/T7BYX+ObMzbVIBfM5jNnuAY3pQ8RfGYrZHJMc4WSaMPPnAV82JZ
f86SNSOpw6v3J7TNmCLt+qzwc2uDHMR5mkvx+0B8KSuvmhKXc1uCN7TWwaKjES65SoukD2N2v4Mn
9XBNSN6/uhj9kvrVHoZ8ImDpLouAlFGeZW52cgbcjIaCOQS7f+EqWoKNeMIfOySODve0aqZB2v4V
dP0di7gIrlfP1byxHu8U00RE9ycTNy7yqWPTCy77+Nb+JDmWDvGMJ/dHf2mT/VO7GKHZ2L39DhqA
CePFGWi47lYDH+84rxmC0YlAZV9OtEohTK+MoiZiKWOwqQ45jV0HQVoH08/uO7laXWfIYJqm0PDB
r2JyYuHYeWFUNdiZe2kVB5Wl+ikEQa3dbDpx4hNDVj7RdG0j1qcwnPZWKs/bSQ2wmx6f2Sbbfm3r
4G3vTa/oMkonQwNw9fPDoQSwJvQLfKMkdjBQj0sZbbT5mYYAQY/jgK+zDICKUOTIG5uNU5LJ2SUn
1bZ00yqgeRVrKwm2xraqpMzEZBcbHmwm5n2G99h29dEyZmRCTKxzg1CiKSnJB04vrhllyBxTaKxj
b8WApDOyOZ3JMSIT/8LxXSq08qLuPQ5J3PHShi/DPLBCuByz3sVo+ezfdOSCtZaynQ8mj7+H3e+K
Wt6WIqZBslgt7M70U1fPCL+I+P00lZZ2m7r8IoxLFt9hoNkkWTM5NnJhw9xlimaJW9gThlshEz2z
wtfGcmDP0shxUswRdn893saLDtosxzA7cs7l+v76oR+iBM/Ib8TJjRjbkamFwQ/TwnMPLxdiyx6l
sB2HJlcCcbhCAjmNfXBKHPeJ8fHofLKZo9iX0U9h+MO5KM/DioO2ocILBZBhrewZVj1hloIuybTd
0HkSOWFOIhj3cR5GAA7sGP3XbM8M72EYdCJitJ9ovav0SCLLDQhkZ9tDB9qe3bF/V7luBooeUuKK
RI/LZCl/w5beOGjInbYWJy9HSbxn3dOwGCTBZ9r2Xi4SxtUyDEKwjKGZ8u7gQJxVtsvMNlVpAbPi
4/dCYfGSoi+qA7PdY1tXdQCGUPnMU2hOnK0dW2zgp8rLbMRYD8Zfkna8C1cKFFcbJzOHE2ItX/ka
HXlbjOSSg0O6DSJxxxBHoBeJBvFv0afprRRvmabd5kfBapKmL4loNXGE14L9HhmlRQiiFAva7t4V
fm8myphJU/qQw0PmqBcRElYA7VjH7hVZQuNUPZHauzs3RuPX4Sg+TdIHa2qEt4Z90Dy4kto0Nkd/
huCpxGhFOuUqVmplef0ydrfwnRvjmVuQOMLD9LtrtQQwvGfLI9fmev9tTNXQv8T/vRVuuU0487VJ
XgFUgf+DuJdnqZc/bGkqBQO1ecQ7EZbnR6aFNwgxRjGyVYxhY0r13blj2xn2YH81/6sufFTBngV7
MvqyeRTlGFS/oVQdtnnhOzwMxWf7AINgKdkegQEl4+wGcHG+QiLN7BOBqb9JHqcMAAvvCZZEeHn2
0EEhTxeke8BNz+hbsZB5IdWvEgQPp1Ahy2ceyYI2S2ngHgqNO4OlZ2XMrwY/yQuXvhvK5BGdIgSS
C9wFBnoUGQngwCN6ZvDuk6N/8i45zJmNQnK/Ze7aLA9gnOWTu5DaD4y1fmtPvgHW6ze+ImbV0Irs
MgrooRaUfPotbjgqyxZtiw98NgZd/kp+1Uk6f9ujP2/1O0MZmzYT8vJoDBPsC97drjNYObqArLFy
hHFcQ+wwl22R5bjS5o47AmCYhAe4p5K+QzG/o+vPbFe8SwB82OyNHZBdxSULsFMauunQd8Xpl9Jh
jcgjFsifc8zNPIr8qTHiF97tuoy4YZnHW57xMaZEWGUJmzZLNuWwuFd9c1uS+FEu/8B5TUiUKJz1
HuimzXQHpma4yq++6p4+AQfnYP0ffnlUvqPwgZdH0iAs5y7hKN/Fn0oPiLGkgCYjfcMpoTiJyi7G
SGDcnaoGb+Vwa3Y2aTDCtXGdE9fp/IxWoUJL9L8QC4fbvonYidHgjbxJA4FHTI/09iVYvUqG15uO
CxQk9MtpBYjYZVUxXmnFJ05+yJv/GLPHPacWbNfxK1qynRyIpehwmtSnxw/ojZpqLHj9qDKVaq4H
XOCLTpDNKwEC1xjC58vvhqPh5dU5WvL/sS7IhexuNpq3fyJ/M7+SX4xvWepQbDlqY0A8cwWv9wkV
DQTf7Rt8GgYZNusaWYh6pMkgvA4MHXQfhawDTCSZn1zAVjN88Ee7IuE4BvMelml6LKlzie/ZCIyp
NnEj6i5rHzUeVkDOlvNoeGcBG//K4aHW5fKV3cN3lizTOcDU4VhSUuYQ17Ln/NUFP/yAVtpQe78J
UtFgMJNiSn4XiILpCNlpEznd6e+mLXEKUODrEhjBzTtZRIiX4c6xnJA7SUa1ISOq7vwmopDTZM4e
3/uUG3BOBvE/25pUVH3Vk4E+ojJpsE/b8AaEuK5fzRxfR+Vp9SNtbw7oy6JV19eirUenVFtoj4lu
A/NBJGkwiqVAg6Kepy/GqJuM/eerqnmgcDpqdTHR1Ex/6njxq2S2p3qqFyjAdjy+pFRTwLE8Jhwx
gL4LBlQDs5ecUOs8Ex0U1Mwk2IdEZzVWRezTkKiMmdWzNsYuQDqHTLJRcSF/I9yN6bodLzAcyPIO
33gxcHwhfGp4/vumugqS8f8x6OlBnTDxXtnavjBI+57Db+3AqU/FIs2NQdD/EuBiRjFPCcuj41Rf
hjYJFoTZRiScqsIefFfWPvdwUAOYBfLBCx+wmCKTbr1333WedqZaBQarbHqdqkpmgW4OcFgVouGt
tzNcxYWZfcX3Nam6U0h0lGjFoiKOcUFYagNYNTq/R/0m0bWHKKF7ZIO279nKjlzgLDA0ypa7MM+X
ZO/D3h4L/LovN1d/IScyE43VYMPRGsAQiaOHR5//e3Bpuuk8K2B6YSFxnhqo1lOd3BuYIqU4UBlm
tAIUcXAnIu6f1DnJXUHOEX693XYrzG3w9l/rnwhTAn9umA2Y/2kVJtt4L1ZPCqH/Yqeego2EAPDN
XKTenkKNpTqfG7lpeSDFCWtDOiRLwkxoWWyLZTYBJ7f/DeFMWfb7axfmW6TR9mp5nHmA7j+Qy0A5
40ALPe8vz4FO9Qdg6MLthXsoSwDVM54Pz+FnH4b7Y9WKHhUrf30vRU3XvUn3n313yHtOev1Ch17e
uRWeeWLKgHjJ4g6srJQ6tNb393esrWHabpRBne9pPWZKXqu0fu8+RkblfJ/bjjtcmJowLp4ca9y1
6oWyqkNm8g/Ze0O/bqGKXy/84x3TBvKSAnmDzqGkQTHlRdmY12UdJRqd9DsqVcH6wOUMiA59+var
dd0FxWFqzmCB8ISnEei07U0Z5YUvJq6h7UGx7TK6tp0w+uw/xJFdWKKiJANfWIxsBl/242/g+ClM
lYQL9cEQpi8Oi8AD4EgcK4oaj8bOGx69vVw3ZNmv5T51homX/bpFS6BD1JZI81Lo6w+skCm+XNHi
sdopfW62G20/BoTBCWvJgwmolx8BBCW7/Fss5fkm9lnLBZQWMTW1xcS6gfoTljFVCpTFNio5IEvN
Fab97/AihMlKvUal+FAPLNUAh01DtkZl0bgGNsITWUqxvbgBC6Fa4+29lztNRSqSXL2L1CH9U5e+
Gq5Q9DGB5h96sN5lUdKHTvf5kv57OcltyWkOOthoSpgVEigy/jIim9wr1JR1t3ApF8FEVKgyTME+
s00T6ex6QZJVJnA4UEBomYgD0RDPCL/7kj7mr5gF5C4vRSKbFuNOzjqvYDnGxROzliGI6dzSKoPP
coCfNQs8bSM+Wr7lxAX0YB6808kk2md5G4Ubhht2RI4duhXi/rtjSYyFcaGsrSpNQ/9Lt/e54bdm
g7mGfCxZQKRFzBub2vNMJ9bT0beGwiv7iXclKq49nqAksYx8uEihjB7c16a0etAUNvE1wrLJnBlB
O4KHvX+jAWk6LYXp8qmhmxGJCcQqGadtf+rS8b9p5AFpNtWyX+3npah9erBgIPysFm/xE6Oy4+Co
walYJ/haFSozywZR86En0cQQodQZ8HfVUl4N0OdnpB2OL0z+2QlQY9bDLiyZSuh6Bjj5I0/gnn5E
LqWGCfg2WNgrQxFmdKfgopvs8IR/GMDZOtXsms+g/EyC1qchQAxbY1sJ/823MondjaYiyRUJt3+j
ylEp6yR/8akJ9m2oYAdBzgRidNgmmrpyacAHJKhK75AMevEq/SS1x3btfpY08iVyoOCtTqnRc58j
84k8TsJdb2lsY00nlsVFZk+ol9uKAmhKYq6H9Wh9vMHumtqx0Avi1tOK+ttOXn6WqedY2CXri0wK
bqWH5o4SCSiBkDQYZeptfw444hC1sRL5IpDnwWilwAHadGOwJfCHl9vdoc2TdOeJs7CImcYrb2r7
7xFJhjvN9X0mj5Y1ClH8uk9692mJkp6UJB0EInIUhS83KRyw6dPh1ZqqyCfd2Sf7WGWCKl/+cqoS
skVeFHvuWlA+xcZ7mIetDYCrCMd9fRSD5YrcNBx38veQWOYaT6TVEQGIf3zwH3XgNdLwR6DS+1Lf
RrxumZ4/RTulyhAUMmP5sha9VN/Sw4oVk0dPV6Q2mPyRRn6bepSuj7MBdJdWFNIazU4ffiTa8rP1
YyCjjkl/ldfMF6efUTOJL2QOcp6EAWuGr7iU8yeMNw3S0x1mhb+ZEyx1dxbzc2b01793bGV5oban
ZBs1gSEKbQArOW9tlJPo67WVcWMeswzx8I44XwDpIEvy4E0Ax5V1p+Iu7Gv8Ab2p+Rp9ULGxAdfH
PySZtLJaIFJnGSo3pR+lXBtYtalh8BwZL+3yfHDnt4yJSy4fwGooYec137rTOItpCB/Npr1hRMAN
Ny9k8TglMXBs/2DvTS7ogIEUARIyYt7TCB6RMSH/HefV3rgNY08DbDlnyila8VsE5lwAdIPeD5JQ
FGhCeoco2laXRuISKoWGQYlIcZ/oX+6qos6KTF20y2zzX/rOsgNNCPFssz10nPQRRq/raSKccJN7
62IVt+XAx2V0yemjUoEEXekavKQGlS4eK96F16jc1TDhag95RD/T/1YpwFvMA5GyMBwvmcjVbYKG
NW9ieFJHd6HrPYCZxbpGPqmiX+7dr8p0sJQlhnZ7OQDuatKtIWX5xcQ5n1LgsbWpcQcvrMk3Vnpu
+qLozZPbo3F0DaSkgX4+YCZb/H85hwjZx7k1s0H1HgvrW7uxrMl8Vksvg0cJj5zP2x4bzOLQ81Xf
A+oZOC8UffKULZY8cvDXTAsv20+A5tADvLgi0Ezsf2b7RgGHsT11+keosrBtzpd4Q6suriU9E6h0
moRdZTq3ghp5W9iOwa/yxp1gcpWr0TAIcIzI87Qw2gaDGyCoYtIupWPJcL44MxqK+XvZbILhSqJO
emXG1R9nxo+ixPzmt66x2J9CQjnDb6rzs1B9bm8EWSY7uL19iEAgmFWO0E3qASt4J0xelSqfhj8r
I1vuMe5Xk9TEhTppjD6lgoowoHvn0BIwCDijCWMOCbXc9oY866Z11vMIbFnVM0kVS+t/5LEFJfRM
oa2zDEl6YCh8BZcjnFm58KVjMSy/mOHQg3yu+GbZLsXdMBRjWqrlvn3jSg4Qs1IwBCU7hB3KUFhu
HQCE5MQ9mQ6wtu53IITBE1+RMAjfFnXCV4Ohn+5NBaBTS/akzGGrq/CCNssENsSUl4Xz5n7Z/V4q
2tfE0MVrxW1DTjbQnhwD2m06JJ0CXpo2Wyn9T/FNRUfak0fnX9ly/s2EB6ePOZHfveW96HBy/US5
cu+VALfhSkRI6lwgHqvYJvdDUBeg10aeztXHdhm/pLACuoyzJN3TZBd3dvU0STcDwENzW8GGKHm2
lth+nmkdbSshqKEyIvGWnIJzwZp/WHXko6sCrnCw5e4ohXkRYz6Cw56v+tpsrOVEzgS+C9s/H/Nv
E6/e81gWAhs0UJ7KI+Vup0tR9EWCWBeQhzBD+glVe1CMbTVaBy0crzb83NCVUNHcsJfdeVWcK12m
aNfR92otS/qXZtnX52l9VkuU0ALu/4NLUiS94mRkdxVkOzWzvkhTCQ/E6xJjn7AtVuFSr/1yV1h5
NzNU9P6wckIVLLaI9sM03mvG7JY+IKkDPMRO0GBrfa+lqM1NVoagbvsyyHPki5mpq2MIMPri4O51
lz4HJ+/DWZpTO2XzYGWotrITC9lsTtpAB1f7ZdeD3ULm2qrT6czrnH0d6zCE4gS7PbaEpViZpcmu
9Vy1UwTbNUBVQPhY77dVM6XpNVscp9ue4plQ9UuwAiCBsD1yHF63K4A28bgAkkGpMBiC1d6x5ysM
np/PjD46r9BBVs8nFlMcZ5o5p8a4p2qlhZyE3fE3+osZ8vo/xs9Xrvr7/WqYrkPpYfQ/erhzyYQS
jLw4Dz0igzcBSaUR8FYOaYGDYuX9ascHyjn7MfLHhOSrqzZAENF9Fxnqc9OLTpRTUdCRibJeAiai
TYfhpbCi1Fa4hI/1OUkKZx9HTmixLLirxzP2kFf8OiY9kSUaJgt0yrENjzvA6pTt63TbGixjJAAp
UQUHTvnLwYKKEbneqb2NVd6+qbNs1donmsWV28GP9Z1g0jvVzQlJEoqcHiClDpz+kCFET7LQCmQY
ElFIV1WfaSlhozWkWBCIoSbwqBc09/gF+f9zD28mfkfCXYUo8eK711yFd5RWnIU3WJYp9SENz2pj
4cRvUSHsYUo7Ei9TrsS1ykA67STWKbYYdHDrjgz1Xx6EzCAw+HOE2/Kf+0ISZKq/LKGyk4fTSw8H
fvuiYNzttLdXgTrn4IBX4diCuooUAWSlL2ilp0VGgyeIgQ9O3cyy/2MwyagbmtacTE+fwiaKpz99
JoxcS+lnO7j+UpTnCdd1YyUiLSlvK9SADjBXg7Bc/4j4PehZ9xVccRnb+tTqbOsnWdzCQMO70MVV
8tqX0HPO4Io/h9K2twkxnAVibJhX6ppsMXpHYEIFWmqe1pv+h29OWjyzV3qBqIFSXZWftiTCV28+
SPwZIo7z+1GuBPrOt6B5EgW9GrP3owTBSrMTpZknfyDG+G0FbusUEyww+bRhqITCqP0BUvCuRyKj
a3xsmEbnAlXaPBeLLlEAaiGhWTPI/kEVw/k6otSGJidaDA16Y5Ei2F7Pcwx4ysd/EvL4NykvQebH
UBvep9dsvy0YMJQkrcSHKyhbcYmbh+a4HuFErexpztxyadM+qcTOJnq0BsFdp7ix0Wwh1CZENkFQ
EetOgTK+I2Vih9zcQvIExnpT38hodzc2cZv7Ib09SgmwpoeTUXSLq/38BgCSOHC1K0kMogmK9EeB
6PaOXJ/BW96pcKVQYg3Xvn8fLyMFweJUFnLfNIvWqnWyMD13PWT3P2E0tzBC7f/OOpNKYBtPgypo
3+ZDKKA9Eqa2t0sbt6VjYzybFFfTNu/UKJOe273HpTXx6GE7DAyMGT/4S1Nfz1z9oE7wTedt6Vnj
BmiIqGXjWF4IMMVmoSZZF/L6P1LH/IxTGdGdudSyq8N4qLKcocqCe2mfvTMD+inPRXXgSkJsfzYq
XZ4MdQDSL59yjOBFtoAx7KVk81twp55elV4F/TJTL3a8/nFSmutV2YNH7+JeHnspRHsebI0+B1eD
rp/i2nPvLczwXVmPf8eoxUDdU7Vbeq8sS9e/nrePCPqaVCT4vT/NGhYGSQnWeM7IJ+543XSIpAZV
/7ODN1F5SIJ7MFAiII4pNxrac+aoWU43raVfb5Bab5TsErYv74ZjqNOr/o0dfNdF5rWphUlPjHwV
Vk9bvFivzXgJxaWHnlbdU585n61i9qP+L4Qv/UaMs47Y/322umiDIqeTwG7YvKcbkegfwWpTBNrb
T4daEYfAGp/l9g88DZ2983dCUMMW931ms5Io2DHnwsdif8PLGS0LvPeaJOnj/79VuoG3eKl3k0JX
iPJdWlXSMbhianii9rde1qI0EcaMhnXZNYRUi0Z+2gjf9JY3X2rFwjyypY/LzLRqKZ8yq5XGaIXE
TcRSh9qFNuRF2Lspr9L3zg+1CpMJr9hwBeTKXW/id+05RV1vI+viYA6At1H7fHoCagC8kErSp9e9
NIHuonzS6sQVysmVRfe4tV7FHxOb6tisWhEwskQuracQEN+vbYfAikCRQ+qqhuPyn3KgfMXfEYG2
JvGoJrUDHb8o8bbb6TrCKcRqSHYp9+An+UJoZ3P2vpcZoJ7549LM/gPKMkiwXSmjEAZ04gmGkMMy
/XmLzK81Ntp3cwW3jLDcJfGo748hmA8JkfZkov4wBrKmAMVrVSyZEkssYQ8TiVcF+/uckkkaXTSf
TKb8uhpYJk9FpROQ2Yu/MIjRP4Uc7bzqXjxZNMs92YY61gIDFaTbr8YaqjK6u/vqCglvMD/aMyPU
lcRNaPdJZQR6YOQ1y++yCADg5LUB8cElBCtgTKx8cCsQPAbUq6LqMtDmQiMDpZVASsjjOx5HJLKd
Vzw6tWvWEe+xa+QqGUEKmxWW4PazZbDDjtul8/dJtFIDHdxqExOTypi/lel1pUVY96kpwbyh823+
iD8O5bFc5ys01v0gF+vItX+socUwpy66rO6xsKb3AFn2Gx9rp9hgul+trGQvW9k1cX/oLrD9Lzz4
rIHB1ontdVV3Wlm0seOu25UwmX0I+zCrcEBKkgbROETcjI4ml6tEfr2M4n8sJlJCFQ/06MeGeQ1O
KK6YUuIvAkBVX58buJk2qVWzd5bzya9WG2J/mSoQTpsSBi2G3uRBEKIgI3pgDbgP5vY44YaSacn3
0PjNOwxoE66xQzsmaNwly1tKEZk5ms9Hx3R/798H5OS2vHPrDWpW0vGDUOPam2rXSqpuYRg9vF5P
iUN49I5viVazhmJhxoD3yl9r55uVGULo3Q+vZ6563Xo2UcT67eY/qlOJga/bhQwoAPSRgJX9DucG
YqclCOU8E8j5ro8Z11It9epQ4Dmw3KmexUnZX8rRaSvD5CgQpdSMZtCHipoXvOY0YnIeDeQOJ8/B
4RvCR1MLTwnNIfvE89IoMFevkDpN0v8hP82bOgA/HRXc/3wa1f+0UBOdbmNc4BIgXa2/rgo0lbY8
YG7AKg4683UUUntj4AFzWgZ5Z9TnRjBXI+ph4Jch8O0/wpDrH1mxC71HIPMHD395W9zcnQ+TffWq
HOL3pkaD4qG0BnbC6ticmhm7OGgwIJE76VTbUvDfbOsJJtozAJ9jL3AK5miD7ueaMP75WmzMz+P9
POT8Y0uswszjFhlGtosgH/RSg0+XyxTyEBPg3Kk4xNjUk2Ma2W7w5EV21oYGQ/B9CMrbfMdVyFXc
L/jSTQLweHK+f4nXhTzaoA83394kpQWp+OTfn8LgaRDrUYHdnsxz+1XJZIyu3jlLHnsH9sLwD5SF
SLeFDbsiWkbK9zP4tIwQqEtHVoAD2yx+8q9/VkVeOJvN3Qqb3KEYz23XcWEsvlK/RkFLhTesyn25
MUi8CmEa/ijKcGMO9u6/CpkRKZLBTSSuydvqy+hlsczqqEB51h9zjXrCDVC4ZmkvmKfkNAaILmKt
EGEQSeGxBLH/1nUrP9/cp01IXw580JjygQtD1/r8WZkVB9g1AQ5JqvGlqai6M/LKxrqWQUtG+kjb
1g2CuWx77hT3NzIynH9h2uZKtfaBDdRzMUvj4LsPrIaVqGuBlBJgjSY4iieFWxGsrK/8bfJInhKs
hj2/hmhVCWxuRZ0Ki//vWTf95yva9STHoSkw4ZPYUXj0IBHus4tgILBaNT1B2XhbsdBCOFCWra70
8ndkyvQ8v9OWH1ZATKiO/3mVl3FRd6tO6u82KWFfZjzbsxLpAEv6K17kLHCPa9yDmWxZ5bH96DcH
hJI2DM8Fv0b20FSIr7m0NvmZD2o92LrkOt1SlyC+upUaHZGWOpktB2Lsk12HNGSGABu7ILXRKhcE
gkqjMM5TRV4RVmIBca9G+dRKj7HFse0+m0igxV+3VZATxp2WYBMlD5E/xVpyo6ujKi0L0l6dBtW/
yZxSBxHUqh4NaMSuOOI73ycpHBKxarVbjsMOuejN4c8+TCtd5tl0GIssRR+7+eTYuy6dvuFiBgQf
/KUVEFX2ClbP1KmTdcUAT7ZRDQK77Jvt+1USyN/F+0T/ZrtG74KUhZ66cZrp935TxJefUHQdQNfD
YrRzxdq9jQy8MOo4CMFLhcJlGPy2liYfpUqxCeKCDWI4ZZkHgO3i8lOgITlBkhP3hSBuN9x/v8AU
cv1sf9d42beUhNGY3PrxfIoZ+h8dVERlXyVXELTUa7X+sfxUXJnKP3mQyGm5M6k3+rcE3V+vy6NN
3RAlkBjVdbFv//WbKqKH2EouHOVmgsqKKo0HXWn+k8tmKXGKlWQJ42TL2wJ89hMa+HsnemK1w8CK
QHKF+ENqyjttVPSKoeN8teyHQtZ80r845fqD//y4GTlZDnzcQcXcmW6fuhC0lpqzoa3VcBIkCpyi
FfB4Mysw2SXbEBQtRPDBD9ejv2L1ksAHMdT1kZKaqW5pBbh73oreNS8FM7qXaUU1wrgcxlM4Xjai
84Zu9w2jT3a6b93gKK2DLpnAaPiMIl1daxjUS8fb7mKQ2GzSca2v9WmQwgmg/0hcNeVljNAhSNYg
ymUHn/1JYZhhi6w2CYxhZnsO/g+aQxKptNw+OfBD/lSNcp2110rta/fCb+q19LLsCWxR2Fx84bIS
WuOX6w+PdcORN3nYHoh3OtgS8zZXDwvnjk+GEI+NzMwrCwSoYFb6SWO1D2BSwZcrHNfHTlJUH9QE
dVSu04v7lu30eIM2bWjebZlDMOueNON8oIha10VqUulnFR9m8xXpR0bDfL2tXMfG1+BMKCX80KMW
ccfEba8NEAiDZSe0RbdQjyTvbBwGpn/L6kxrAhtibqTDGP7mMCmnXZI1saR9BSH8X4+hjQkP0XVg
VvHAjZ/nMPgDlsGuRUQjtjshgg8Ihw+dbiCBPxIeL7/OFW2ONYjjf3z3+6/Xo8JUk5ZPDe25WjE3
eLBDz02BiaP+OYsefrInLDXPPWx3MBDOUZvdYw5D9Dwc1CyI7mCIi4padLdTTP8qKM3GOlQcNGnF
aF16FqiyH0ihnuC/tYQs/9RQKY8nyvrIMGulKnx3XYLNQxs0NxBtRBGkJewPFNnwoNSKJztuDAhr
MDODNoDgmADAvzD+5o9li+unzOF1usIk80cVlm+x6WmPptJyTNcVVRRQCy9/8n1yhxlhpYqO5hvI
TZinyqtT0xVQPDjg/W28jDLlldR86vk5Ggut0mgFZi0fhcNgcfGKGpqg9rCUsm8eyYvlRnroIzvc
O7dejft+f93t0LAkoBWEps+bvpGhZd507f7NUtE1NpVRnYZgGZJNqZ6JGxwb5jGjVTwkoq7m5MHZ
/ELwB1kz3mYumbCtdwm1HJQT2x0M4iP2Qy/PgxMsICQVoHTDB69xkNFcYk7DvPsgZUD1xtUsB4GW
JOoxQa9E4kDA1iJuLsfVaBPTM8PMg++lYWOtjjHEOaLGNNxMBjukEX2hlgZ75CfvnGJa5YA6FPyX
4MWRUDSJhCoB5c9q9XkeWpXO2Qg1Yus6+g3TnuYTZYROQwWbaCmBPOX/xt+GdG0SMcMhPzenX50u
7MAJ7xfzlJ85bcL6lqDdirz/DW+axcAVm6yEeAR/2vGCZdL7O3PfpkNd8Zn7cXq6sPVYRSD7ysqH
uBYEBLWJ68BOxzk1FvXQEHyUIUkdtd/JbMDL0IvfaUwZqeN+Ygk2qk3/pPzFYR8+Nm733lP1EgyF
8P81fc8nncgasG1Q2YllwkMOZjiOJjdMhSpQ/S7mg6SfOcljNknrS+bO5iPv5o0OIN4Tc9Wjamtt
yLjSxn7XS+BIGw3cd+TNwI49J7xiIhZCp/jRC5mfBgRIKsQjLNCIIeupGuc3azjjBmROYeijuix0
EL8UUPK7p4DMeWKiJXab0nt0N1JCjvSg3a/lMxFIwGVbp7xMJLXerEVJMyXSZcKGUtW3v2/8hZgA
ZEBHsf5AM/mepAMSDykLQDAO+TcYUyg5lQd6dGGBxHXm6P/BHD5wAgwwVQk/09I8x6bH/e8F2LjG
WLyHUv/w/WExZJw0gsDhahXta4cr8JIY/YiKg3BIv49IPxP0tbNP6HoOdFF6p+0JcA5gku7ozGQS
H7PkVZmYDXVr7Sqphz03IWaOc4PZ+wABEsRhKT44pLtzsRNHMMEgXB3nCaDmiOpO5bgTi2qDPsdE
3GcAvItbCMM8yfi1oC6z0vBIvxmocDRF5xJLa+vNstGXKNq0bf8ELUEIEuZs6zdqluFnOQpX/0e5
AQEJfJx/rrwwGOecDWtrzTbLzJXH3Nmgys9O4eEKxT+IhsRf88Tz5l5if16yFyW9mABLCTdttYuq
wYFSue8aT22qXP9RAd6VUuiuFv/8FwtOBm/cTh/xyscDOOW3oxwdN5OcUBjTJIRBokiR91AuWq5X
p+KOLl8QY9SREG/wxCDeenNALmrV00Y6vT7SHZuF7Z64mLQfkiydj4haTy2lhAb/wE5puEgy6yjB
fZphNzx/NStpR2uTXclEHBNQdn0zzI68wi6b7mtdP+9D71fYre8KgdkXbHXfW8iREEOGxLFByLbf
lq+Jzv1L4e5IEuQzYUYUolUJa2NB44ZDXgMKj7k9TrM3AXfvOaIy/XkWrbpNDn71qA0hWx//nJBV
j4sRG6LrnbTboD6CIec+Avfs4spz9uUur2ql4RP+FbVECGRsjXc9exJ4v5PqjpCdIXf0jxzR2LhZ
eHlMDiIOmfjZHVVsMLt7+hMcXXDgO1NPOcpbpww0FoEdekNrNGJOlDcXbTHNjrVRtBHD92FZS98o
ag9Cep3tKPYDu+B3p6A4sf3VZO8vDM+WyddfR3qo/8yNrTkmrRp4xrRViOaAM2WDfuBVvFTQdsTN
zHyAlLv/h0FZ7ca7f5Hia258G19OcZvaq/PIWt2T9Lx9mnhUwnkJfmYgnePtjHXukiQSWmhgXfmw
u69/U2EpaVszZpgLSdCPRRwAPL+m0DuxdmQgwiSHofvTVWYTX1p3TCLTMO2/1X85inmfhqEaQ+lF
Qcp3zjAiMOpVzGAH8m/JPuiO38MObRSLS8q/q6K18x2bn89HtBzcntFpflSx+Hnfge6NMgxz5Aht
DcfnrWSGzFCXskRpGXU64Zz7u+fosoyY1tZJz4NY37otByOB7XlNi9DCzIkOilu/PEmYrW9FDpdX
SILmUbYbFOEo1iytZcetrQ5yggMJDb9Pvl8qNHnVG0je6p49x1Vcx0MEigSdmy3nW9hfvUSX96A7
6yM0gvzYbcPQJ3V+YQvEQwxBx2gzXLuHFXR2zZ2KtlDxcdnqprr8SAdaECbC/9Qojlyy7GUKVUCE
qzKha3gZDx37Fgy388oPN1S4bPZ8LJ7vuNGGX2w3fntKWJIPkMvAzqEFT+U8BCGfe8nxib1gkSG0
2VQkb/JLC9MPUqa18RkXPxaE7kfMRF72b823R/qSLb+of9Qm9zGrFiZfdFfkee7VTJ0cffMqaAYW
ZgFOCck4wo9i3Akjo6aROKd12XXfCDkw1b0rclQ5Ohqh7YbQPzhnUm1RtqFcPDupOAn4uw3mrp55
p+S+2bWIRqDLZ7iZ3tlMqiW7HxAJkDPzlYoxXSaEZ+K5cYCXoducvnY+2QskCctCzkb3R6GUlyKw
DmYw0nUgaWm1v3wI2CssrSJRFM0XeGQL5el1R37yzVvhF0YMvp1scI82+QvVqfwQu0TDXo+UvEeW
2JkCOBzkk6pweVwm8+HZF19SB2FLD2EPtGbt+J2VcNDUZFcE2c9v7J7qoOWJ7bLY9INfNAEf1lvS
m5cJIocp1v+oJ4h0OgLkkt8WyBHgYQaVwzCnUKapjHoGdvZjoMYQu0i33m44bca9FzrTma9mAw3D
VGb8EP5fauQcPP2Kb+hTqtTy6P+kPBxB6nRboKtVOOf2BSIUYjgJcUZPKnzXtkYxE1hG6STu/9fn
Ld97tbhxYWGELdt8uLDR/8S47aOudQGpkqzQQGAhRXXXD9E5tNSBw5q7TzYbpxIBNaBJOCI23QFX
nc5KweJ2d2C54VZmEI2/kUQeb4KFVtzBieyI0ITXoaAkp9HBZTflu6SKt80t/r/qDW05zNjcF/hU
Iyv1YrWuwb/jtyXsilEnLDafvrqUR0rqdiiWbgvgV3aclt6HGlo1andyr3gV0dZkfTtjKUhXsFUE
wGpO9sUTdFCJaB3adp94sKusZb3WRGjOKLBhk74H6UN+2LRJ+rlhwQauBOhsQAcYrYULrk7tQQkp
C605Yyd/HMAcwA4+0QDeNzszyRT/y2qbDQodbpWLMTUpqiHOv3EXwQTaBiMRU9CrLxQ+3gsEGU2T
fOq3hKsX1J4NIOQaKX0RuMVAU5JG+0UGNPLJRzJfO99UsdiUjA2dSzsKpw29EYoOvFKL/Z4wQp9e
JnmKApRT2Kd6dRU4Qd0QB1Onoc1rz1ly8EXcteUzEdFwz772Am/rWQp0OR3CahjtwNgA9E84UC9v
s2U954xJveSqoEvaEFHDCRwxD/UbS7gpn1zCi6dbfag+95YN8ppaAnlJC627KpdM7JJBmc5IAHky
YIJBqdx+D338qHsevuuOzV+cNbhOLQ1LAUf1aWIfCW6bmDlnEONjJhVmUup0yGooBZcAs+k5QgCw
s6qkJA/iN3nlzhV1uZiT9ADOihTa27CXNvCHX7Rs+GAExa7aLHIlpZBRBMYhA2Hx3S9IzJTrAn4h
F3ITFjUvFl2fcLkL6pJeW09zLFnHaGREvYfv3sEqi4Y/PucUr1Bqdkgu4DniXmwi8oBt2LCyz+8C
vmm8cfD4M9foXhoMzOiz2sZGBF+MeReYbfWjOLUH2vTe1Y1uWZFkdUT5bgE4YTADbzpqF0o8ES87
xyO55dXnJrLz8254OfqZ5TlLDyu/hB16N3VOIINwWagnXs7JXZoj1GKeFo2oQhgTAcNOO27JGnYX
bD2ad+NVZIDVAdevEsbiUpl3jZ9bi0fDDEip+QbScrVWrJncF/qLQ1LhCmIh7YU0ff8vE4Q5Z3lB
/+cOOIKP3ebJkHleYENDlAnDToNy8VMp5AqPzme3kwIs15o/AQqqa3kWJ9TWttRXKu6T7TNOhtlZ
Q9AecqmWUJCuos1F2N0Df+p9XTg5P0cRkrEHZeh3Znd1UP/IaioivJh8c5D33F2QacYjmRdPkQ2L
Vrn3/Q+JJ0I4U99u65947iPJePc0ZYBbn4s76PTTLc85xXUg/JlKVBn06/PdFGvdwKa0zBKqki/Z
Lcvu34jOSCCu8HgGFBXK42CgalC2aXl9m90tfMRESHyDfq8wPBt88Mu3TitmCp7/+osiFIZnDxui
IJXEPMJg4gTracREp8w9pRi5hyCxts265U+hEfUmPLbrDjCw6RzWg7lRSLNxJty4Ar6ou13+CF33
zQQ6qWXBZ5sL9TWCMqpglT70cvqy3bQMfrEzM5FV8Gd6/H9u/MR0LRUnlmWmGlpAsnIICVNdiTnX
XPCKKX1VX3XA4ZtnWEd3jzdwHerqgjR21BkLUjjJ6zqtX6crvlajlYElBNO47nADwHv3XsLbg7so
/DwUet6W+ddFc0pdjH1c6Hb4126z52oG7tFwsm1FLXkiYDNwQvM3Bg7loFbOacmUobnCLZBVnvxt
IJCZDnO0zTthsE8lhAfWkGSp1jgWvJtO8oCKFpS5eC9xHy56tHPns/XtxJjeMNYZ0deaVX/9/O4C
XnKpwpngxOmynPPlavPkmYjFXuFmhAwYrYwvi1qTDr/6L5KvHO35ZfxsXola9r8ZNdKtx+XhcfGe
/h8E6uC7bdRl0kVMF6+R1uY3IcCbFggUauMrS6pJTRfamtwTtsiWYB41zESdjLH9hzyLP4gGwm5k
fPG71I04F9hoNhmhJ3+6wZjR0Rljeuc7PCcSbSeC+O+Qq+6NdI+/0kpfly6oexJ6h0nQ4m2MFH/0
zpgP0mM6fafpwul4BKGbjRiEze8yVwX6ZuYL6pr5T9lFXoUWnepbn5mDsuwqMlGaYv+QTIfLUWZg
UF6NJbEz5zJJXr3EdsnTJ/mR+b0X73u0Ymj7BeWVJHWj+2GfaowJ/G0YXnEgxYRMcy98c5g9xs8p
jrTmLJgCfaPWGqMhySLVt+oH75+icc0ETkSsu0TuK2Ff6Rqgc2O1uX/I3561bmS1KFa1jiEoWhPr
2k8n+DwYImC4OnP8cVaURICzFcm6j5uBcv9bxVFyCWosFREBIKvPl9MmWSzKosl8gKyqJInKCPt0
8NxDgkdHj1mhUQCnwTwDdHUBvUqe+jPZGjSHgnRqvB/3k1aMUM3e9iEG7RKtVgOH2bAe2gMrKvFa
P+ugKUex0cidcy3rSg3EoLHBETEJ4AFPd0FiXNK6Z2I8thYNLMahbwOLISpwKapZ2lCXpDf6WLbK
fbVon+d4vWElkrJqM6qjL7E8eknegk8dd1UNSFzqNeufd9TWi4EREQdtZ8qPn/xc8CjNnM8WZB7h
RaO2YL6kmWJS3bxesUVZ68an1CChGGvX2zjdUM+YE8mb+gTJK2Vub3yYVCiuIbDdbk2krdOfkkse
ZncUpGGr9dSdEIKjRlZKrSVNJki+0KC+KdllZF0hHJC2FEE7fpNglTj+QlN2rMVv+Ddo7TkN4bLZ
CMxdW4f+f/1Hr6oSHn0/ssXB13voapBSiPJRKDAT+Fg6SxaWoSEg4evqEJULkhr1D1rlIFZmaKtx
xwJyM5pi+bErcv35MIZg/kf8OXoCkgQyvoSmzr/UeQoYSg+ptyOcxM6oJEupg3cijcCvW4DrJzMc
MqGh/jJsERfBhnPxQb4yWe7px7Xyx+idkT/fxoEhe6H8IOUILQ8Ez0d0DgJEDAt//TFGjkRLCKAW
X0GGW5U4dW50Lt11fxnyHv/kW4exhlyWA+aXL44gtRBL2LINVTqIyYbPMt7uRiJ1z8oAnq9C2xbq
GMUtUq3a2I0vgHCZoBWunAj4gsdZCg8GqWP2Wu4ZaoYqNWlR9QB5kchAp+kke5/mM5TO7DxdEZp+
4zEExxmjIWTjVWx97S8sI5VHSabZd7gDeueNvBRdC3n949NAFDyrfZZn0x4iw1jco4bVAC6Tk0h4
LO9QOfrTVX9AqZgQ89UCC3+/xBuY/OCb8DOD3rXXs7bN90A99baRGECP849V+G8U9TLFiG7djxmS
D0FuDD1azML/GUwAM4VEwB569s+F3hp20Vp0/fIBqjZ96vzkddDPJcbsxKZyyBMNBVtEYAQCeNZM
F9RPg0oujaan5wfjHaqxfexMLSPW1nsgWDl86UIEQzAJZxrkQ7HeiQLhhOJq9ICKMcOxH6lasG23
lhQ8IYV/ARkpeflgedrD5OwAeSate77EwT9Um1Q+rUPikuzVa3umjaNhllmOQdj8PA3EOTsoxjSY
hBLfM4TVd7MJJewpQAqFNmYPh0HexRtcvPJCA4U2Jh5SuOJlHHvn1FpTpEp0xcqXJ/Xfq4EUigL8
RbWvEeT/GhpV6NGlAuMXyo+zOaScVFlq45IpchKc9jMug+c6w4TZeTorBy/0f8yoNHLKFZ0e5rdc
JZ0NZVaMTCJ3OEPrGAhXPB16RF9zxXf6X4K6nojpdH2fglGX+LTPEJvBxtS4jDfzV77yrwWh7n7g
eRIKQ6tQWSdeD8APYG/zakZ6datXcUAAGisW3rTEKVGqkc/MjlaPL3QCewg3qRBEqBmSSn42gTwS
sCcIfDkkDFdijabdq+XV82bDYqeeykpaoNmjtGzkCsxHXvOZn5pYTRoO+hQ37Xv04Bb/rxFTTKcz
xW4u2cnTiFPzAsgb6nUgGF9/tjnBk5xq5I7mDHeh44lEYMOmsV4YLyvzPDtYI2fhmmwgbbCOo7fr
j+Yi84VpvBZWDC1UOvtd7t0eBh/5EDOhkSby8ONvyFu0RwkA6AtLeZbEdV/DXoCC0IxwK2hjSSEt
eHDLPpvjk7ZI7JcFXSsnKp4W0SwdKsPZjfQY85JczIv0G/JEXBMUDrQDAu/7jEMHm0P2KxLVonY0
y98V19KqRRQposOckgLvWc4meL5ceZQq1XHZQkNxlaN9j5W3vtO/Zi6wD0oF8NfB4nYOISWZuc2S
ac2wRvfg2Zotb2BuOkCwsFbKwkH/ptymMFz7YZcBy5J+w/wGJpIU7hZuwoO8FxBA409e9zY6d/BQ
RWSmwMijPk0usb/vLrkzQV1F/k+JySr3X9lwVzaDbCSqZsoJ7H33FwEHdBPmMPjUbd4HtzC0gxeF
qbpdF4gGZXerotRTs+To0XrnWfBdT6QnLpy19yRthUHy4GOSNTnMA99yzeEsLFUFE+nbhEhD4Uw1
6HLDvQ9sG3TIvypqWWGYsfWsFVei26TaizuOJa4JhhGCt0AoXizHE4zC4HLk6FU7elq9rPzw/X8A
KA1KAd+RA3Q7TdXmqLGrTNjV3PDhRWJdiW3Q8zlVVL6mJgUrEHrKokoxqIrag0S+7iudbasomuzl
zDRAW9bmXbSBzczPdGfzMfaHqjSZB64LxtSfhIjg8Y1sXUNkbRPSgVOgTrvtosiSIyjRVMLIxNXJ
MuFkZK/a7PgxH8VqQLU0D7+5IK2s6NUSC/VXPinf4lxHn7jV6GY3/smPUmnr8CWEc6o3YI9iJxZh
l/FwtRTEcQY7YV/1yKfwHiwBgqz6PDCYT2o8VkKiaiDKhtanxVUwHbg3r3m1azK9ci/1AF8DfU+6
JSrlaJNGRskuwiBAaLdM+wNL7AxTry/7jZVScg5YYjiYKhaRgHRjSbVh1E7gFu9HeichRIEUhF2h
JUJBYpTGZ1CjMOWAsbgoOargX4X9ghFaEcacKnBjIRE8Y3wVkjddbkLw93vof30RXIanWZ2GOAhB
BA+GMLAsBHPl6pPuFIBAVte82stjtRmq/1uor77exypkuRMvp787oorE6mwKA+Vk8Bv3cHUEsX6i
/pq/coM5NtuANWs90iGMwfqQMuxPKqy78jBfRsGp4erywk0cFuusYUu2xuqbZY3l1MO71ZqM6TLh
pGn+3BcoBYSxahNU1uPfHltCE0PJAGTklfBZWOG46FOvXwSqt0ltismvfdjhVufMcfEz1nYdivSL
EzwKUhJpUGvc9RsH7Bn0QBVIKWCJYMkChQ1FG4ThvdPxO8arfZwW2XsW+2AO8NRlGPoKivJDabPg
8ZCUesIhn0YQv9pLxoXlqaVdnt2QPlVsMJicYEUjRlHY7WsLhgoBbltkOA76GmbiRDnzhrMQmF1y
vjJoPdPXAxtmXbbUAAjXnSE737IV2Fr4TnWkL2FRW0G0wCDFI+6Jo7fssv4LFU6i+gW5KJahZeO6
Y/tBdjgqd6gWl+f/5GDgDPek0vW7l+wLlB6Jn+ZHF+TQHD+XbJ6Pvm+SmZBG27DU+7OM3oZLOaXz
RlQei9XUrp+RiqAt7EjJMud8JgHj89q9X95/g7Wh5k6SgApSjvQprCKPWuQ0baeLM62Ni79nbgbY
Cd7WFRgftpiIEqv0vGiRE0ZcnvODTi/H2qP0AXYe+Dl2RzWIB2phznR6nJQVUpmJH1jQ975VSG9o
qCgXoM1/OVuq0baOWnN8IQIBgZPIbW056T12e6x0io7YHekf6aa+9bk3lmmIuDaoW8RSaz2aZuUm
yAK5oO9niIbak5OGyHFSIwSB6xJ5cWCeFmAu/IFwzTN0U7vLugjX1cL+H3NC5Dol0MColU6Q+G5w
87c8uYJzh5r4ntVge48xcwnZDy5VN7a58u8o5+7H//aBK2O1LfVI7DRpRRd5sWE2jwGQRWhP0OQ+
1l3UgGTKRwXjt0oTZTAh/uLSthtJFid753twW1WChZlqAOVxkyCBzoR98Zt+T1PQlL77RupFPhk3
8O7kcr18E8rUYgj2g4NY/+sxLyb+MWq4Ae6qNWGhdOPNNSba1RXeFaauyZ/ZNOA/hQUa1/TVwBQ6
gjDaD6gQt8kYQGsy34fij5TAQ/qJ4UR/TseN4xX8WL3pIdN+4mK0H1mCSntksXqED2RxEPnp0tSo
0xlc1H6O5cqrD+09puqL597ujXBfjaoDlJmiW8hKyaGElVQ5JpRsZVTVhrS255Dukm3e9h7KSBJN
Klr9utDEr6AruyNJw8juVsig9/M+2Jp1hsPdaR8jbMGqMDy1QKu5rfhRcsVAKdnIm9kXuhpy1EHS
OPGGIQKYMsgaOt89Fuh+py+09taDTpOgdQaAy/fXYgV9TaFgu8jUmhYg6vPpNN53b3IHya8BX+pV
PNbX2e/1GiCJwEm6GtWzrTESvy7YYz0RqvMYQOy5ocKg1iQPpHd+icjlzHZkzA0N3sMv9Nhbd+FP
b0vWZvobOpXBnqXKvZPUZ3ENlgTNBHCxLLPcZn1A8oniOej4dBIGr7oQflvGow39K7reOGY9FqoS
TDHGAP0RSXRMbj5TTSpJUo/9m+QzZ4V4SA6CeMxWZwtrPwpdw4/G6Mr+qNiXTCvvPqiwwNQbTjJx
BfE4iTbBDuTz5hbAoFYj5jxLVQ5bcLVhyWoHGbnKPUfsbWrCtQWRkddzV5CFY+h6fyAolaUm+EPg
XfFo7BHEV69MYoRK5A2qLd4lVWQh3hqcmc4YULOCgfYcXWPCxlIwGslUTIubbwuHgBdOdfkuGspL
A7+6nv842WMOJTxS1irvDP4ME6kcl7bCxcfY04RdmZ9tc17EiPD+kLqz7No+VsIN7IXhkE5Uubmf
ksgkAPn2QhCZ5bWDA+FNW5TOQ5g2EbspZaZngIyrXU1wCL8+uWQwKhtPNhXTD+QsfbIVQB1PYnIk
5OHqx4j8xF5iV51axuQmxqLYcBvZU3SzIZwPQm/7V+e38YyYFEtKDB1y+S6Px7ghJa51nefk3xtq
Huk8XN8G14p/3jit4DfosWwF+IdKQAwGeo0wzxgrtch/Wg7rDSmOBCip8fmR0ogA5JSSMqd6H9VP
0zK1ZOe3OUaHLjKgqwdxuIyhgEOCIr8HSWJTTyCvKYPJ2SHsPnVHFl/WOQQdUztptAtOLZghIWqH
cqC5T69W5BW68DgIqJq8gMul1poQU+l/R/NoaMuaIgnZ1nxRDaeZgQhzMP8T89It6RAygj3R3xwn
L56GCr6v6jwu0gPnmd8Rh5u22z5iuHLrUWiu6Wkbh+GSxWC9+L3BR7Zwm0HTd6Q7i0rs2lUd8bxe
1m6oK14tG/a4/c0GXQ3esDvRvFlt9HKiCYu1VK9UT9VxeJNsdV7M8gYvfvBmn70s1FAnitCuYAc8
QZcCxq3Hc20dVZe2SkmqHrRmM95tNTZtubHPXyvC90a0in10ME/GNutHXnK6ZPyZ012wZZiVSCaY
X2JW0cgPx52dcvnuqZcEYTvB1UHbJqrDMRZbWrqhwjgozz1Z5om1TYRK8DClvpU3J+RjHc2AfXt2
C9OhtMzrJaYiqVJVdibKVFs8jmhsiDu9Qu1NzLBoZgNvR7AfudoGoG71KCDobiOuAMNs6MR1gczY
f7x8enW1KSkslsE0yRjVlbFo7mtvRdH+27ZrpEKrHaoU2cpZri90a9UkcLzurCx9wJzLoQuRGCt5
LSGJ4NeqXMtRX9dU4kFAqdkUV6GZdzbHx+sM5Ygmtyjv/+rw7xyDHSPJ26Jr8WgE9gNemZixLfNH
Ed/rJB1afNhuzVkkkxOJydZRWMi8idLVXDS8txPpTy1i/KSlqBHlrLYiVqQBs67HB91dS00CMIsU
iFIdzeW2S5gtaL68zccg7jChqkUtfQsyybw4ioOu5zbisAp2iiUEfUVW8iNBLsPcMTLPqjBHfk/V
QwuPSyOw2/7IMpxCShLI1lZ9wR8K7G1ADx155KarVFkciDSpCXPYg9YhxCFdTLDeNdzGiEm0DZ/4
5wUapfuqfk1RMCbJoMEXJKhj9UJpDu3vkuRHsqJznbqM+WI1Iw2qqzygbNU3ZoJ7gaS84wW4muj7
M3cIv6iAS1W6BF5WafG86WqqGCYFRN6+bHHtPnqe0GbQjNnL+38hoJIs1q/EImlIK0qgLDZqFSe9
Em9H6v9RDsCIVn1hmrqClzhHq/bmRIcb2ZjtLeKTgbPG1YSgqS86ORx234uu+611CKuUPdFoCBiF
ljjRdBqpCCMUp6UxoK16Zcz/0oCkHIgrFX7jKXTV+/hO3h7B3LU+BYap4Y4ixWSkAwlnRpZW7nSs
CvrwuLkLSmWDcrHF8E87WUn8D+YoQnojOMdb22lctkiixUigNjJpuqKpYyPNbh5Av1loh55fkoeA
+acvR6YJ5PXrV4LqNpFu7LMiCbL4ft60PJqAPsZlKDSzZyMYnx83xt/6J68/QfvRg2W1US6rMqkR
QHmHxm7xmsLdPaqxsA/zT7n+Kso5kcURE6gcz5IpF9Y47cBifxtk147UNYLrj1lfbpp/e+CF5oO0
OjrGoLXF6t4U2XiVtpVLQafjvSXOP1qnkhU95UFom+RSvv4+7X4BjmjDzjzu2BBVXpuBq0ZtrbnQ
0u0csb2fcC/CST/Vi93+FZTCuqPvfNxkzuyRQOGlm0OdyAQoOLt3VaYRQCe3ahaLUqRU81PGRf1c
u45ULr2NuJJ40DupfDJRLJs3vOdce6zKMlYRJpwuCkuXMaPhxDr2FZdLfvdZmjuJZ/5h0cP90AfJ
dgucV3xU37/33Hc9b5YUvPUfNot2bj81YPuYo2WdjBfb0UkLU2x2KeO6+X/8+0l0CwQHiocZWzYB
QWUPU05rzBmN3uYb+RL8RjZZye/wwBsxK3s3Y7H3bZFb67ptl3lVGaAgv8sQQuBD8ofY7HUB0qay
LhIDahLllyaelGqVrWUTKL4Dz9qCeRK6Yd0kTylBBZE3l46onazozhfv+U7tj8zdcR7vxU/XguLY
9CUz1IxCQHbV8wZkMrT3u6vieKjc91J/oi+Oqf8alC63upSR6Wiw2rucLo0QSF9v+mx6vIAK3Aia
MHBfAFNCo1ApaJ5WPbw6uQhMJR2AhjPWvGQgfCRZ5UDJqn5iY8nK4/uIcMjyzOSb6+qin3zUcNqd
cUUKfYOa7NVXlvXoWiQV0Ez/fZTdHcB0QJoH7+ZhCRopaW7GZByZu598XbzNSReuUzdhbvW63i+A
pSqllW4zgZCEzRTuSMxeUrc8fDkT5uDEoPtal8oWn1i395Bg2YF4Trv3MKU7+MHAuKGJTg55zFpj
K85kiS0H9dPdpxDGWxrnnKXDj+zwP/XRiJiDbms0UFs3txjkcyHA2ALOaV0TAIXvxa28Aym/0CGg
QZyGojD6LJ4Ru4gsi65lwdqe7nAFBnUHU7diXGiXFihJ+2Jtof5j5XLExqnXrVdAgSoOfqXcCTTM
eH33+Mm9NxMsuIBrIFVHtIrMfk9ow0RQdlAzhihLS5IgbSC8gsV7X6zYeXfSMzIngOvK7f18MoB7
2PczN8+oYsI8J5OuTzCTMVnnShvgPOsawq/srNrHRAw/X8UuW+zW8omxhL9WFQM8KaqYpRbc/Mz3
V8tYdcczSA71HhjjzEPn9VOrKUKiohqWKGLuEXrDRprtJpk7vTM55FTCroRE67V9MVNrPHYxFWOt
ZhX9fyb0IlVNOKOrZEFk/9afNyygPJ6DHqEOyX0j4My5mfIVr3beBVwJFCezAxkAcTCtXO0mM/qi
OFzkNWs4DhR62CPboCXo+0as56oU0U8LKmg5sg+IEjHG121afZ/pmH6Oeq2987z0DQ+ZfvOJgNOt
5cniN23izjCAw55tgIAKQqmvE2XK4WVCbvGwIH77dJ3IV9XFd4NvDhcZxYrE3V5STX60gRXJovXR
2lObuiHM4RdZYXVb3cWiY1+Lymy55nVcmsh09et4S3dsOrCqeojI/q0W0+h/5JJ8oEyOTowlLAJ6
8gu0egKjctN5r1PX6T6YwDLK4wdNoEXzR9pVWxdPAZPNYPYl0HJ1UJi7MpbCMLMNx6LcYKMdp0ke
gK4MNct90/O8++pAw41bDYxCoW37fh6zk4+yi5uIPlxqJ+hEouCDY2cXSQOIvKbN6h88CVl75d1G
KKJmK0CcajxNE51QpY0wBn0GdZ6+tkehiYnojVOiOls5n/ec1RlVhpG+kLogPAndHOpvI9lJ5cf+
DRpbZ70nfHXCFvKbUSfyr6yVIW2H+k+lyknjHm/xfkrtmqp7ThS+KTiTxw5x+kGahaGGdRXE1T8p
iW942jp2tS+jRMSRO7kzbJG8UZ7x71pQ5Fqa7oTlyPUBtgYy5mzHMR6Akn4UDNxKP27rmMdzk0OC
LKQWPPRtgnpN891rra58iO70NVoqQ7+LLd+hrC6h7NV4/f0GDQVDJVwhBRZbHSE24oIDyiq3jcH+
193Kv1HJHTK+vo+rnCFy8nrG3ZOUidX+dFGDN06G2z4Wxf06fVhzpw1qkPtdWwZ1bv4O03bGXNXR
OBGUOEK1gGMtuYSac4f+0RbppxHBs/AD6K0qV85DssNNE9KC1c6YtbXJFULfUEIX+bEvDsJp9eiM
M2LYo5x8Xr4Bxfou7OVkXlFZ925TWIuUnDZW4n1iGU3Gt8ovW+4XM0JWkTlDU4Z5zy1b6gcwsypm
fchOCUSkk1oD+uDDp9Xbx0tdsPVYc+yqYZCNrumjxkrbieqIKI8pD7GHB/fxEILgh7M7A4sE6kgt
LnKfz8vdigyh3fTo7vudNvDACl/F7KjByD2Nu2tB4OZKqLWhFmWjl1FlKTfdy0J4XKdPqWPyqnzx
cfP3ZckfhaaiWuV7N5t8jYjG/B2DIUCC0GVZY1N5Aq3XgnbulLVMF4BtSfsTlHLgSiFJ/+B+mljA
ImIjBaKKeQFVBKHulrnoOhWb4f5sJ20QQQRCLiuVEcnCqW04ViB+FPvRI687php679aCvM+rpcbk
GnwISA+ZCJ/jNj75Lsmi7U4WUfy+MknqFbaap+BG5LG5XW0H4rWdHecpvL/2hsdlzBeguK9dnf7O
DCZ3suZb6cnaeAGGlsolA4oHyP+twOIFlimRxYlqYTjWZvjnCb8THRtzQzy7vsTqP3AolxS2xo/i
sYUy2sHT3fEhfJh87Ht0DM558awb7xCN0GiHeCwmKP1/YufAbOyHV2MYj1HLkzoOQUYaKumL0xPb
GeLH2uTF5hbOgcJKxE2f25tH4U5F0PK4+UE5kLS89fim2p6q9/y9FBLAeD6eAoxakcXJSlrarqf4
VZN+DGIqwii+LP1VKiyLPg8B7ktN12ePxQdsFEDyzHNIoZh3PQ/5765zAmn+snO1b+AWePWt4zE8
tJk1HBzzPXUBc1hBfCCQbuhT4EoQ/EQMgFYq9G3xMQb91Yk/pmrYJyHGtpcWlMoFDVopNGCAHHax
vcrGRpb/dTP0doSGQKuTuSClB5z0mZ7w5qEgfGycKmoYLEFY+R+Eq3F2WgLz1ItlekPIB5qlKRiY
I5uiVaEeYoRGB246UdUg3glmMVcwrOcBEmLeGHKqzgLfR1MC8h51DnsrQjx93DRUIuqiTQjaKslg
YRQOI6swi5AFP79ZQg9KvJccXlLjDklAOnD5OAApqg5rvJj6nVkWsAge5S8mYxLNXW8IX4hG64Oc
0GHitwlumaKCXcwvmQFX2v/7ez/r8Mvxw28zNx78lsL2SXef+cXx66997VEto/fST46rO5UzDv0w
Kqzb8Y4hRcnUoRZFylQN96Wt9CJgvxrUlxjRYm976jZyFUJCpgX5ERwPAQwkt7BEpmv7ocPyeO8W
jCAVaN9Eu7WuFHEb4dZAZQpILdOrFjYpp7NBs31WnY2Wq/YHNXiONi3ELUtgiM9M8qBw7pjLKw/C
BEuj58KLxA3TAqB/5yxhzR6g/FhGW0qQ2ges1qOw5SIINEEzX1GgccU2gErY51QITQabMrv4tYom
TBn4fU6wwnWeT6IZ2mGASF2Yp+cU9Da96y0vtmC20w3YgP8ei8zbHfkTPYXfy2rl49jaOd0Fy/H7
1yvpdDPjTCfoAg2k3TAB81qmS/0NOf+JS+aza+RFlkRAaT2UWRV5/MaDdhDt5ibqYngRIrnyjBD0
ypZTXLcVKp0a8PS8GwmK0dPttjhjTXvAxlPRzoVqaIHwKAGZtQ3ENkgdqHa/rDdcaZJF/ffzurpW
OywV0nDIl/UkaB8b9k7mHryjoaxywBpMI2595o0sd3Eux2sxfahKStBz5iyHenJHcUsYd2BI+MLd
1Ursq26qplcvBdr18+rOVLYUtpaVI+7YveHy+hjanlpU5RSA+dVs2inRhjdRcWwtfeHZH5TgpzK4
ib9xgA3pVkF/kjFpxKhipFCWI/OHcocuxY1M3C/r6MORXHz/E/LtGapKuaQem/v0itdJN+l0rKwr
U20Js3axr23S+Oz8rai5lpIr1xghf9uTOzKRXvzs/wiACbIn6+g8tEk0y1uuVIh1x13XlhJ3MJi4
pvMxriWLimFUTouuxk6lw/3Rsc8w37jFfo6O+coPFy3RRQQo7Lcd4U7DgkMy0uWUSbaf4sVShINb
DJL6Gsg26TcV47PNdaYVOVOywtbqAfj0C9aj85ox23pCE1RUlYNmx7Zgw/djXLcS0habWtcXrOxD
y1r950fWCmcpIuyvaEvdivaT3eJAP0E1Rw1N+cYuP3Ehd8XehGfZcH7ylWAwUQZ4dDUxo6nK7u6b
Q9i7WASiysr6wA9Rb4065N3P7xQsqNq46Z5A4AzilRyMcBv772qMMdJTjtMbCf6BeNCSLnH4W5e+
ML/OX8cc/34749n0s01fxMA8mo5pY2+OzQD8R+x+CYwf24NaHW6mDYsOUZVfadfT3KHVncl6l+tV
FiyMRTTO4QbMBjxRFppWB2w3gAT1QqdohViCZ+zADvd3BEaw0DEHgddECpU5jweVRv7t9e0KMIvk
AMB9bfYPJgasaVleSNGQpmEFlhYX8EsooIlSAsQlPDtmBt/dA53FyRp0VA1d66mj8i+6OXYWxAT5
LRjFByv2tL9DXVPaMZNvLxBgVyd9N4/bdfYHmtCnjKBTSO0UhoX9iWk3Iinno1eGuokmzLG+oOcR
/ci8oPOJk7EuexRKqe6dg24mJxWs+zGZEQWIL5sdkY5DyjnL7B52t8GO76LKfOJEuY3JljjrmY47
eEwAK9GWcOkXdqvLTQ2UkPm8jd/IpJNBis2OoRXG6jQRv+1QS6d/uVwxDtwXCOMuWCAxh9bGhRp2
0I1zLvpwhHflzMJOb9JtwMjbjnqKex0cz9msDQz9iwvpV8nhJn+qF7TALtYUXjDcB6rfdirKkTUW
dgKTE8qj8XsCNyFXp8lOnbHzfBUlX6J0CXEuDm85BIG/b52hYpG+zQd7lG/+uQZqg74mA9ptX2R3
UgIlLiMhE5CoFNsHranuhD+pUpB2/GahY1LOJlTOBsvM3vKLH7PbcAXJuKimQsGKnARt3EqfSvM6
+/eUy8D7zpYl0HlvaGYL51TFl2XYjXi7oQzRzYW0DFKZPNeM6nz61k1/tEqZR2kydtCfU18b1HLj
IoAT64iMkomjf8wq9xcKMEQH55lQ7Pv9lm5UiNPLYxt4mdATUS0OuhmXYnR5CApwI6dzDoD1GzZm
Xcet7bKkM6ex5ghNW5MAafQ5zPLVtdiFZGDl9eQT6emfo79UxI3WGd7pBdHuaZK0J9vbjeJXSrnd
eHlpJCQQd0r0E3tkKZ5cTkemvdjuekyUciKJCG+6nbVJKAxiL0g/ncMRaDOOWscr3OVqCCWRu7WD
a5+eNjALtziTFhPIMljLKicBVUITMcPBgx8nESaqTBKN+v/oJDT3F5b0/YtlQBjKKGbmnHXrQDHk
mCv3cn3S+V4FkJKg48yMm0z0NE37hAuw7bt9RxEW8YKfw5uTkr1JhhCxLtvOdnffkXykxiuxmG1l
q4SJVJRU5frCpLGq8Jc5FmFhYpgjgP3c3MCt5TmNhLkqGKZ8Wk22WE54f4+kNEs0vtsJA/g5bDtY
mq7gV06EyBMykWxX8DVij0/ChWOZgwpAyAAlNrPiO6hA8GrVF8ahQa2YuFOtoKCkc75pl9Qp6HSv
yi6BQ3ne1DY42QrLpz4yeCnZYdNVuuMFYx++FR4zVl6+w6Ag0XKJcuzt6b300NTllhoMyKBhQe5X
dcJPwRlAgOcitvCE/PrM2CZyMfKrLkiH+6drmxFV6h8jhUS2jIgF7mDAEgz0QFIhaaVhYQpg82py
zc4hHyINChHRDE63DGgSSASw5sRRIYra1t9ngae7atXUPk7sxb6KAxj5AMRiwAPI2iGRr4Drl8yj
T8kBydT4PCxCWk0JHjC1U4OCDkOYHyOYhXhPKqI65i41h9nx+pH0YVHCb1amySIc028YJjA6aA3P
Or1eJDOOARoQIXWKC4Fcy9hXtGHbpH9l2TYOZZVhWqhXVlvn30j6zp3Ghp61KP5ejgy1PtJR7JfX
nHGPpQ7atpCWO8oyJWKQA02JyngjQP5LztHpkXUMAJ6RgbG1J8Edn4erEqV790ugCLNKtnSAlzqJ
9D7Auo95X6Nt7ED6h2fJVLiHybJjoPUeyindF0tWni9OJbtLObEguPeDfArCLMPhLCmpP+jrbW6q
bUd8aCurJdcudMetderamvRayhXS7RxyzpFJFMKIL+L8iIFfAAowOzDeIWw2pCez9Tq9pD85281H
BlxOazJFuvJaadPSb8uO+W4Fyzcw2J1EUwsJiA8S4V8YL4x31O4CPHL07ft4o1D4EXd5vsMPprGg
sspmYpDRKbV/MxLkIjnRAtrH+QN8OfNkm1DWvpqW16HYs2suOm7Cgdz84QSCuITe7iFitjsXcfrf
eKjvfDu6331Zp8NG4enzSqJlSyj3yBGncWJ0rQFdoyDN6tI8op5qo7HMJCBqYAiJFRlIraOHJcqZ
gHvDhQ4mQMXcPs2g47ir9ovECt2CxqNPJXaIzBNUpSLgJoyDK9sxUyTRdZWWk4tQW2U59AsdC3M8
Yk3CSczNSU6s8T9LgZcS4hfjVD8LNUmpEgq37wHKuueE2TNVBdie1czBm6DrO+TrLMjX17TsZSne
EkLZjUy3jFeCALs5dBsR2NXiaJpdW/G5aH1q6nWCRLFqklgohxs4ejPMRG48PgSvCohGdrGdGSDz
WbVwS7yO74OFzyN2+k6BpB7je+Rj1PLroTJCJrdIw6G2Vpz7/46Tdibn9BbqOTXvQh3LhNQNK7wH
QtYIS51xl72ikCgrTLUjx8cruM8UG/wvBMyusk10MwJ5ZAOVUjXNP8Z1LEZaP0frIFDx/GgfQw+N
JY54fVy4zbyZwN6PvJjhlK7MxYJOABIX0n2ka3OBx7dfpEyo6LPSIwPhXuJT1A97iwQj0ueiI1nW
a14TJwHS3mu/3Zff4zkMajRoryNkbIjTAnu6qaVZYMX79bhPyaVfnWK8vkz+sQPL+yWBf5Spek/O
C1nL7yBK8+Immf/8nfaanFB2cvEUuqqvOsSnbM1U94NyUWXe6LBY3bAbnj4mr+6n9D3zgbjhDjSr
WG2mQvG5MzSHVbJE6B7LmbLKGOB50OikRfli4/LDu+ZWgq/NzHSP4CkK3Kn8fVUs3Iffd3eChPBe
CKaUBZWNFvfoOYewnAsEzHUxbKBl8NylXqt1DSg8UsiHY4F3jm696A36ZIrwaun+yM+6YTkyf/js
/PzGTO8PQ2d2sU1XYAdduwXJHewSHUt3VHkLxVKFKcp28pTtI6+uRiruD/0eCdqfr4RE7j9zseX6
EpzFZV0/Ls3RXgNuKDvHaq1kzwcIDXiGLdN/pHc/QB3xAqGccFBM50EVs2vQeQlwOvkXE6chRJVW
PX3i0hGOeAnClUPZCt0DV/Y/giucsbIMVMqyHK5j9q+LSXkpIKmPAnDGL9k569rti8lp5tLh08fR
SwPvqJtzwNa8aBr+hrh7NdgN2S/ohuUyoJ3aPCd+f3uW17/DHLXa70PQwKtcajmCIakMvxD0AF0s
N29HTnjS0+6YklkyUg0wJRYpGJ2Dcez/s6kH27qtjWr+Az5FUnljcyM4tYLaVAzBQXQFQRwcLdLc
5dghsXrf7aThjF1tD2XP8HRSmPWd0WDjrXJB/Eg8qPdPrq4TTV9HlinWesBZh38/dnza2IJn/U4X
84QI2KlXbDv9hfUAytH1hoU0wUv+jHDXXLL5eXHsi880w5KldA9QK6KnxBwGEoRbrXlgOUFhbven
IMOXhsP1xBjSa6XTUUSSmGqS2nhTlY2amMkrDHC2FFYhxi3NmNXsZuq83NG2eGCHPvPBmuQyCTYy
yMuG0vFjxuUY2gONr/6gAgI9igINDjLkEQvxF4aEeDFbxAwhbuQ9C94mtgS5lmqAba1aLGqe7+br
TgGbSWpKen/y3TLneWpM5a23NRYVFKT/UNgXPs5IgWJi10BzsRNIOuVYlamlglm25poAX1/j+gP8
LoFwck3TRPzae3inChrsTvssHv+GKKmT1OmchhsSnaPFcyeQs+80ylYKGeYlp2Bc4XG50BkyJw5S
4mBFL4V+Yr6ott63t1tQLTKOFziFSE1EVtxoIlnWSkKlzotrSs6U6+DdOFDB3BkMd56WXxtmgHWV
DQcXHNH/I5+I7IYvbZbLLEe5l3MtPqevTZS8KyZBE77toPkyW7yCGNoNMgeFBRx1l1MOyt2w+VD2
pnOs9XsyrX5oKuMh3KK5WwGYoV0KMGKzQRXwX0w1Z1ScVpmQXdXFa1j9mseyx6sDXlRTDWF/Qz02
3MgqWo6uG+/sVqQgbzWpHK9eqNRVhmOEtVX4PVomCY0ndDY7j/dWAfZwGcepXhPrkIb6Q3DGb60C
EWLVt72j6dYtgE8vqIHtJ1GWtWPOJpxU7mO1R0YiYKhvDdyw6+/gs1Aud1vb4FkNTXyvO6x2b0yI
UyPPMgfLIE+ri8xkQfTZmZb3m4poF7gnyyPXMgtkeU1DG7+0uoja15FSw12uo5CWLvEZVBiY+AeA
vIbf5y5fO2M7ZnQu0PcrfkPDzQDSuG1BKPHotogQ+CGiBT031bxhPJD6l0hoMpYy0H+vg4034Fte
zNWVQvgD+xizs6p3lNiK4lf36QEokbf3LnxcIDd0/SAGBewi66HLKyanh17+2tmBPLPTZAne/9C8
xN+Biuxs+bQ6I364ImvwI8dfMeUyM9CU9N1iZUUsEGc4Z3Yr7Eisnyp9zrf8g4XDf8xiJZ2a9wQA
jO3gbsZvgYwu7Znr2JvBYWDpr9KzXCqdBxr1eZrqm/lOPTpIUpgxxevgcJ5Sy4aKNHR6vgni0VMF
unJXFpOSiq4QBvAB+za7G9Tea1iCMWbzfyUqY805IxwtQc7+gZKUPPPDuSsnnpzaXqLV6gSrGZu1
lahMT2RV1Yva6HQS0lrsuiHIDCS9vyc263Pf5muBTORVXOQgrgapntCR3w0lIHnLYlVloCmfKZtg
Q2Nv+WdN/Ga8PFEIOkf0r5LnfGnRKINY469E22C4kCz2/40uBBMzBxpRCeOWIwUJoQioSBpzVExe
keddMwEGbbtbMzCvrYwGMjqb9vzOf6hFUgDbfeTvG5hKiupXCzSgzCLzJ3tiyke0WI+aGMx5SJ3j
ZSi94M96gekLk9707urzjI/acpvslVtBDv8+xI6plH245qjnB+hqrbIXUp3Mgpfi75v6BAjvG4y+
I4Wa6xSvy6Nh9wF5JEovSKH29CV8DbrrkBLSbfRc5qkfFr/FsdiyTQxkWckmc0xGulPWyB2DoR8H
DE2Xq0fk9t9QQqhYPeyl5aTNKB+Hzw47weixtX2P1cbn3AZ0pH8Zo59SQZ0M5IS8LYAhUqP/tuiJ
MeuBRXTt0B0wh4aXN8hk9S4aG+w/923hRgL9L1klyqaJU6WCNh6rkny46Wa4uDsjMfggHYW1WD1b
O2lPMc38Y6qPFR13mHSSAwE1G4NCgmn2MBI8EcBbcOoVeioYctXcpbSNMut5Kgay/i4D/LTRG7rs
hsAsCJ7RazA3J4dEOdLeg5Hm6wGUptsn/iqYD77zFRA4KUZ9fHnB6R7Hn1btqjVw3dnjlfgVo0M9
dWiv1HsBxyxbzvZGtyJtNzyEUCBcKnSueIaJDbKeyd+g/aIucsayWxwTJQ93kNGKc37eSwjPx4/s
hRBq8aVxYl9hV8tGtxIyYcnxIIVGtlpFpnD4SOCJaIF3g+PzECPu6BpzT9MeUTGu1r+nm4yVgIKu
u0Dwl1M8hEcveErmL75y88KZ4ff+vcQxMLaADDzyZx8hQPxTNqSR0K7Or+pEIQqvhruuyxgHCcur
dogtdPeyFGwWmBcamdFuKBDPgnD83Gt5DvQPjf+98LGvFjSMQoZyladqFlwB9DcaG0KZYt4KirHn
ELE4xJyHerhBBjb+Mdr+1QaaJvQ86B/+BobW0C/S5HwnZbPieAIFsJ0EzMdwaFFlha9QciWtVq5r
HLj2GXdvBWlVgn1kwEt3b0AXW5ylTa9T/6JawKI1gVwc3jKLj6UFag/zdRy+g7TOfpltxzbHvThD
gioOIvozhH4+H9sFAmctLSbVApBFyeW9hm/bYRUB6cbBZ5n7/2SCHKXLA/R9ADl5kUQ3q/tHR0Ip
Ia6WCtMKPOD0PKoscm6r+DwuSvWVeTQzTh/RCPi/OcCfH6FO4Ztj1H6oDDhyCxT9Qi+YR8JJDbna
8n0DG+6T489dhXdWKLYBTI62BMfYg3R5IZpV3KsnGt3MvDGdlT9eOIYTtMdmXHqyq8Yfbpq/IDOg
ea6JEv+EcZEFSz7akVTZXtY1xqJCYVUdMsfVH/CHHaNqZwgfjVi4sfDHlahvtCMuU1eevPgv3LHw
6xAB63WC3JiMT3A27pClJudBBg4AIZ0CqJgPbUHhYdRxm6hACIXmy70vwFxESEtRcTKDqVQf1c78
t5NzOY2rLEZOCdhGnaJbviGu32Fyf3MAzaPqxhJQFSJ7dByXj+OtTuXfJBaSUHDL39uv+9Xtp9zR
E8J8i6BLw0C2ZOqcwYALeX4GrBTvlpm4vTGaKgUH9pIrr0Zm9P3wSUCXHoc8mtCnjtfjSh4YPbGr
dvQj30PzQfUto5NWqWnD4zauB6S1Rj8DFlnANAwjO4Gs7q6rkYl8ZSG5QbpSzvFp5dO3I4q3Cr0m
8hWTWhCfPiXukARZKXOrPY8UA840YlsG6fe7ujCp+nSNmeEmEf4ALnCl9RNV4yZ6CLx71Q7Fb7F2
vrN6nvRjaKKcwNVdY/8YZvB/wID+dDko1/uiug1TRaIzRhTRL0KiicjuHl7XWSVVoPrRJay4Yvh0
LlUA7GXNPXB6hatsp4F9qZSgMK8fqlMq5tULOIYOgKhjsoTKqTjWcF2lt0Eqo2SJrx3dwEetRD2g
ncyz5M4QksxB20wLDSB7zTn/96oeT+XN/VJ+QLmoVZO0zvyb4Lsic++fM2lPr4anKUvPEczHKsCa
6mkn/+HTKTPfSYhUllYDWfxfi93zPCkkAqGhnSl11xX0QWlSD7wu8tnxIbsWQmHt0kW/R+HRl15V
JGObernKQn9weacdgagM6AR0+WaAlctyqjKjuAqtDcT9lq9ImBLrjQUxdaadUEt/DlyTIe7l0OsM
iN5w6XeQHQ8xZ46d6sttWCykmfLJJ2QGWbTDV327xki3ScsmjBgFZgGd3rw1u4oMss48zFeM5O9E
FfV60OpcDZpj56zlfrkNptYRYSwdPcIou3ebHw1l7S53tstXaKTG3yoywYITcT9z5kM0iZ23AgHv
wAaqUKQuLFrlVNrfYPAArYzUouY+o0Dutk2171KibDcEDGcqkdgK6hiW6153LkHTG8WvVY5oI4Hu
xM/Xt+xAgZ+XAsEiwz2Ko+BTgJOwpszR5FmhSceH6EtEut3Fc6EKrwEmyuf9D9tu3dAJyxacIfiI
E2Ld4/MKE//qUtAYv4H+YFehr/wYq/mnEjZ7Hx5mB3vMDxCwqCaPiLuGvl8BGjFX6bfIAskHwP2O
Odwnu1o48N3A7stYnmcMUG/ZmW1N4HBcsOKPoni05RKKkCtNABXPpEb8IrVcO7TtNr8UnsrcViSD
mEQ1i8pvIjV6g+K7r3L3Xt/T9z3K/pSZo56VLtI69MAiZUtIFMs3wTAuptUuYRUTFDR5h0BuywOm
0PEC5v7/jLx4/wYUOCU5knYEBIZwSk8uuF2yo39cUGmwAvZbsonDM5/XvgFq3YZanOcqv9G9Exy/
g00B7X84ul+vXhjAX9mc4qTeZKHTZJoxFTrJ6wy76BVOghGa+iMbk1DDDPv9ta4uHoRwxmhpVQmH
UnikJPq1Cg+QbKB+unTVon0yJ3lhVO26+1qX47HVfnu0Aci9YVjJYfIjexqqm/vJadog0huomuMV
Feh31FeCl/lXNcZJJ17q6duJitInA9/XqYA+709bskEz+ZjWkkotPpu57d56Hf5ZhPLCoD0tVs35
AZdmAQY0Db+iVla0D1JU3KzYpQRwyAgpkYPGcF6ekaVCldo6s94xcS3HUWSU3e4ykCeb+r0zIcxD
on3QEAtK0x5sRGP7gk4saWrlt9mz4ZsI5VbOStULclnJy5tnJshKCBRHPDfsBHF4+9xXkCL9Vg32
RhC/DdWQLnTdHqNZarL2JySqGC48v1MaIOVqDZ0TQcC/z6jIxjxxWbK5v3+QtEMMShEfETc/W6k/
xGv3qcgUNzhzGXQXTI2jzpmvW54sMwUD6jXnC3M2QJj00caV0Y4q07vgFI5Nb6obxmDi+boWXsD6
Hss2mw8mN/fx9IkIaiZYMxKy4tf+JVeaCCyBC+WUqcht49l9BHC64hCeLROgBJdn9KVoju/wwCzv
HDllqhUx9Q4N3wCdt9QZjHT1iMMdt5frKlqGdKvljKsUL3SBPpi5dNqYxTlekMP87I82Uk35jDVZ
9x0/D0tbP8qyTq8vhO8KdY9fg5Yx0LVK+9oBLtlF9rsnLrlJnCzaVfn4K2KwcrRk5rrsXudKFn4A
nbv9Ma6HOMI1CMmzDG2XgUIg0Ej8w+uQ7k4RbbkY0D/42jaGwv4sJ+Rm2n4AR6WQptsLdlEJnIoG
JV9hddd1x1ySeUjbsMfwLrV7ruxMOMeMPrzYDWlW88QrJtVMu6VDy+dSwWzR579xiCqnQXKvz3xc
WDp2e3FlkEnrnWp5pvWwCOiNSrG3tsbZ4VcioYgH72Y/RtHCOTorNl8ty2kAHFjVzRkt1m9cxPI7
LesPFRRinADiOg7blGo2A99yR28X+sC57prrNhF1GwwcakS276QDsKttH9TflMFZ5e2yXg2RZnyH
G9mK8K6tSiu0AX/qthMaqFIi8psXULRbeEDa+R5feXKn/M75swUdChg4HKJcgZmPImLQGBCbD7Od
fucKxz7k8+sG8um8cTSw5oMSEVSclhBAcpgG0Jdc7Hj3ErYwqqGlkzfPXQf37BvY+vZEJWZ3fJVx
bh8n+krKawGZ2JVVAcjVX9pgfsxYZ6SQJUpQgYzdQBnD1emvsqCTIMoQTYN9qbojA4lkmIlSBS5U
MpFsmNE/5eSU/31RUmXQ3TWhV+0Fx8Fnv+pZXHzM4hibH7jfjDSwebXl1MeWcJ5cHkhYvPjN6MUV
wvHefJ6Jq7HOF8gR2YnmXJeojMGIdagBe6f4HRokOgkCDAQK2S1lJ2MoIP49vh81aGU9PK9T58eM
FTqYg25DNBBC57OiLueNP/pLS3UvKll+yhxnsTtCJG+HHGVXhNNV+/bhLfVVs4bk4L4BCsCKmTnH
8uP/SPtYhpc7lh2fGB1OQh1IC8x3wh892zfl7VeXKXU0lZtds1Uy4pjR0nhY/wOmggwyFFphHzE9
L+Dm3vCoU2rPjMz/sKR88fqzlTq8Gy1Uv/swxY4dHIaLA9+VxtW5XUPVJv8sI5Sx2+ywtI7ULFPa
tOKJE1viN4KLwamz1PTqI7l3ujFrENZiqOlS84c67V3564yYdy6cuWFGsEyGKnzjgAZB0NOqgRdA
IwNRw9SaDkdJ8AcisVGcjCZV7quLSPIHB0TGi5YbaGUExserf7hNYixDhjz+eSExqM1rHQ69C5be
FzxLTQ/waOv7TeB8hX9mmMwhVXMzPlLOe9DngyEZHJQiF80wfEjjaz5cw/3KmtJ6CJeguKGt5kTv
5BEtxWf4ucF4jWHIXoXJinG0LP78jxhNL1UCn2G/BUh8ifhWHBOnemJHEXSDdGXWH24iHQoy3Ndh
XMzfLwMLiRQUQjjnsNlmfBuBh8f/kgHYFHVIe+nLlpY9t1KyZ3Y2GMq+f/owRO+a69sLRqaeWBZ5
O18NBooiimm5wQJq1267ALf2OBVoZXUWzd80J2Wq5fGCbVdIOjx9C5iErxXZXvfZBhliVnJn8M1f
J8BJdI1HN7DNTo2E3UOkXbopjv37+NOohfBX3Isk98zu3sz0ggwPDc3erXDbztId5b3CaIMNcCUg
VRwOsfSCO1+hwm/Olgw6DPLDAostJd15Z1b2FQQzSBcWXlbB6+/Qw0urAP4SXdhwNiS6tBNI0JP4
O/N8g4mUPIFv1Un3p1rRszFQIWbfCZnNUsr8W+rV39wHTs9+uW0+5IQov8yZv5kk5za7xxmjtPH8
adXyl12582ugKXSx94ZnfjcFsXI16cre/alLiTjDfHqvgeLG2UBVyWS+uaZkn4I8pURXVglsre6d
o4Vam5MuqWROcuPQ6pfaLgrphnxY9FagB+fnPnDPzPpLjnjnf4hhFFa9t2WmGuxecGYe/b27xxsA
lVplp+q9YeLIorqxyaF6ndtbJ0x+aCC5FiUpL/ibDd3D9p5xly7FSEVfZVF74ogsn79PoUbTDzKp
xvD08NMvDSX85ibgoKi/qk2mb/+gjXMAif7MuP9nVptY8Ai4XyHqa3fAjBWt8RqPg+qPKIFRQ77C
ApvxTic1mPV9UVtHWKrfDqlzgoKMj3m7/OQn4JFaNcukGFCUU/h9+IQ9CwR2DZyZeSikgYcKcgxj
0GjxxqNuky88SPokFnG5tGMUgBDHaJo/S2unEoz91rA97GyQe1PHpIIG5nAXCa6jJPRWnnrdUQwL
kUB2mU1SJ+m3HP/lykkxlcNm+9cwLMPQm4L5psn3rQMjQU8GaY9tMvVqjdhY0cgfT/Vv2ANM5VTl
SGCnRQT//6W+qk2hwfHRGa8LsWVjj7wQXddDZW6VIQrz4FCNEiW0rsjZrqEm/SOWPuX/wlSdWqbh
jRK6ZGh6PRqIfvYNuQI0JSRs0k3HWpFsww8hflA3sgcVbG0s6mKJ+bsKb/kfFVa5EkyMS/X8gZvG
K4X1I2lD45+qAVBqfyBLaBnG5Th2TXzTjzGT4lWaJ9ACjQeh6wFJNtE9TSiL1xzGrlULUtNtF8Mj
rFm8m1YB1Jp/d8+pUbDLLbbRdE561claVw+0pc/X1NPDW5tptOq8y+JoHTerNVJbYx6M7uyboUOi
IAykdJFAKSrNm+3pEwfhms+Au0guPGsxY57mMZDIZzbjdT1l1QZBP4V+M0HkF8q2dXNRRdVDgZiZ
EwMHPXj1jgMoDbn/3efj2QHhMlX3WbwLOKFRXv9GAddYqm8R7XrB1R0fgdRdcyfvw/jDGFg4JWLY
K15etKwOQ5euyIt/BhQHGF3IIU9grPDQmQV6uqb6QDo19fz9Wdsqti7ktlkNXoGQAlMzWrwEYleq
BOSFyMx1O/278tlkkLaKd6RJjLranW18I14AOF8d7qXs1JL47HlGNZKHml9j8mMLEgvCAm6CuNRC
MHq4zFLoszQEqa9fKUyssg92QRa9DRIB68cXIg8TKsHYKBHztzAbFbVCjyssRnWrR0GJu3pspaQw
yCrsUvE3LxjoAgQagMiqCWpbaVskwlpTU+78JFOJDagSejP2UD9ZqK/+0Y06Ueq9suo/oJoZuals
zm1hhnAVPcjAGLXX37UgT8S74isFzpKd7DgdbcKMVh+QttevFO7ITh+BRK7W5hz0FfgpHadR/61o
6Ghi4Iupnr5agJ6Cl8OFHaSJBQacwJ+lXsXYurQox6LUJ1iO0lYTDT1WQDMawv0cDBeOVkr1RohF
/t7Sfn1i0kPo/zitITprUqk4e0fXc4fViY+he2zIFdAbNJ/9vDLRmOHxM4qk7TXCBGN/e0zeYBka
ZyKx/LzFnfW4k8yV+slnW+hAeCbU37pRsbbnoKV/D0qg4h4ohZ3KRmC5n+LOKcjh40PKtqPinStR
ISx9eVv8Qv8riNLXb0+jJ4pn7I1TSpDfw5jRCKFipRxxXbjyVXivzkJXmDt9cJXQUV+xvMzczEPE
PGmBU0n1LphU1KsXxDuaeeBgEFUX/XUaRYDrQYW+V6EcJnBwDuOJQG7L+7iLTRszFGpWKu8kc6J8
JNdKNg45+iYjXIK+Kfra+KchriSGBfAdD8Up7v/SqDhKSPZQCPxYTUpGJZN80q8SJUwuXNTkuDY/
UzgNPjdKmatBEeF7erUErslYGwYoduiziXWx2ZB81gMDLTsLWHVdovW+bv14rf9ijOylm10HsGga
6JcU5kxfHct/pbFhoJWJiKbYb5WkVkEr6bSvLuAf9UHy6KX2XKzicU2zk8EDXtco85Iv1u+1Lmnz
qdTFigNLxLRpTZ+tuJIs+mSJ2iry0g7BlVrMOVyxlh1uzhChQG8U+3XDuDV3AWoEiQ/xmdb1Mx8L
eQ7jFXv4or+G3h04OUEH0XdeqG15ZnCPcScubH+d774Qx6B7G8qj6r+PrUSL4YaSOlANRFX2+ewa
gXKRUVrGxuesCn/CeHA18Cqx5SL8JgoSuHNIbJSb/lJoB4jDRxqhDHPMnlaGEd9tY0W+igs52yUs
0dLfsjuNPLk6bvzQhaCKfQYm0qULB0rPJk9B+CICxxLbD/QqFmUs9ycvaILUY+AVBNUYti6hVvGQ
MawD5iCBpl0rEnHrrvpSVNRnSxpggCZSNT1F65YrelhE8Wjc5PjEq/e4SHCNLQxfE1xaW+9LUQmx
g7t524QoH87wY40P3QsHvPJiK8mJQTzZNROlzhCNQYDwQqImVh5TT5gHJnJpm7SUTcgpZ8UqZmRm
5pZNrXGECsd/TeEWLrU7kp+3QJT0L+ZezFvKNtORFAEmN9jv5sp/I6avxfvlOemV5ZldDzNOFLsm
DSy6h1tCOK8kdsqkS25nRij4uyOt3XftQGY6xX6WEB17tbM81l767tv00fuZbT4k7561oP7CSOWh
ys0jAnU/HkWA9Cnl0fBN+64UXVpfPXzM7QPyvnka1doKES9vSHy7tfmK/411TSgMD3meWh3vBL7s
TEgX4vNhCL5JHQyQP4U65XJh/9D/yvn1xcEVz0IN1QhFrlcw1hJRGp0fR8DPlGsKV8s8XNdMTw1x
pGqB+VCa2nGNYdiKkzPjSMigV+iaEOtB8AkYXSfqEwYYNFJO2MpnOL/nD8SO/9q1hB0tYaXqajqv
op7nhG34MSSZdx2ihwpDR6rYCVwK+IZj/sQxgynMudyURHgixJs4ZBCoCcmcboUT+8c77h7sD9Wf
dSFGJnIqtlMg+8iIn+WvG+yHx2rP8AeFEgAbcGEYfwSNwYCqaKHA4sVLL7ZJRhK0w9O6ix86oj1+
jDMRvjpzrmsXHR3sV3Iqay/kjPwQ2xkheHCu7BxSpUSvTV1va1JdVXKmuIGqUex2ZU3XN9v47hNm
DPorFKc1k/CUxHFQtl9hrIhoFooTBi/vudyrPztMXtHx0dirvC6Ntr/sIkIWhCgd3uXqwFqG6BGv
EHQL3Z2hNfGA39R6EjNv+4dnBsCbO7GmyL0F8EkSWUb6KfmqVgBGF9xQZWD/IsAaeMWIM09jP0J0
hezEeZLINmeGEUSfqijy5bubAjY8NZcCiUVH25QthHO3sAQer69aZ45pSbTkJcGiSS/b7PqebnCD
P/++upXjx+Zki2AAx8Zmf6Pcg0vjwi6Zd8U5BTKMbK9EuRrtUO7GjdZLmJm5PbP32OGGKc2XANA5
VzgZ7Jlzhf2F0gi8l54dvZWz64ecfYyCzCoKe+JEt2cWrCY9H0y3R8zCUULUqGONG3bl2CYj1NDp
SJQjKucbLJ+gvSSYhh3m+xgMYw+e+YGuS+6Lj79XTs3PDXQzgShDBxiJbrROGUfNKkNDFgWagm/o
AVnm8wL4OnkhIBnKXcBfhn4DubKKNj2S6UzadTYsCX7RgSadqKKto551YW+5vhRiUq/QxyNYe1Ht
YOae/5Rjbb1PCmtEL5ONkSrYIUOh1kXgvxEB/XJlV4zb1rEPPTjvmWIduL4rUiX/eDXKhwkerKa+
sKxnRrv4j8jjwDwDfmA+tv2obanj74JKom0ZteOvE6GCjIxIGE3AfoeJnfhY/1wQdAmByJaUpYYv
uH7LsBM3CgQaPVA9Ep5IKa+H55V4F9XvAQy5c9hEDE3gY+w0A018TpHRBhq3pLjp+sFy2E/BWNNR
qU3JK3Vb9HzhjxHD6Mb78VPUhinDUD+hWkWzvXpfSdE4DfDw5txFYdi+kj3Npt+WXgLVaTV7czym
8hT3j/M8WI+OFFnMKLYG8nMGn29SF8UCtn6pf73+PCvE311rituX1fclF7+UuH+PgjQ4yg2M08sc
Rijz20Gdg6I9aaGcAa8DI8vuG2DodKRp7c+dnL48CmEw2qA7IhzB+wqHcwCtGpWFOgGxscRLpgqs
S+J6flmKPBSUOts1YAc9SWG5JgdUChdM7vShgzVR73uhABtYKj64hP6LVlqumL0msctu1uhEXRO9
11ILIfOlxoRRuvzP1hpAT7vGaheMNqTxF5IUws4b4tDgFjqkMzP9CdcCodNU2HWKAxmDb5WkFLCd
JwA9isZlovvdIWRKJ9+mLlgD3bGgv/mQnBY95RIzytg17ktOBzh09BgsCbjj6+UWOUQgMow4pfEi
zVeIzSHgg63wp/E5EY1LXElHTOJoYvnE9h67at3xkmuIF8F73uj37EDjnJIpolYoIta9o63yGAtp
MxNiV/OHZgMK+82Roegp4/Kzqqr5Qzy+vl4oICHFuNXK0fKLyvjvVP32GGvLpt8k7ElwtmT69fUJ
dZwQRrR03B3tMzYUh8H8hnKdGjkP3ddYAM7Eiu0lJlXPQbcH3R3xCLIz/jALF5WYZzCNebgyYbn7
iM9s+/KJg/U/+oeZG9vfaXeB2rfI+ob7RFEcPs7bpGHc+L3pI7y/gBw+pgPf211T+8m3f540Sz3w
b1l5r5ZtSyBZgJazf2ikZlcVEhM1rGS+k35EbMXImkupJ1FVt/aMIn2lC00cBjObF1yjcqrjp3Hs
ef7KeaKKq7Z4tbwGk3rcRFLNBQ1bCfE1l5O+DY+1ttBPDaf+SnoglDFxopreIw5vAzTyIbl7V6AX
ZBfvqFdckzqJpsDd5AILIO5/apWDkukCzcy7E3xaSEkfcCOLmCk4Tx5lQpn1Zg5NKd9iqZmPudNw
9WpnwsiddYcIYqmyuiTDMcsUs1u+gdSLKJ+QclXkuPPZXmVM0yFS5n1KbJ24KJXSvTdCNDeWxa6D
zrKgGTWJYdAETF7lfB8ToCccCegS8Bh/uQsRPjJjk+BtYZouoaVDV7egcLbthMLUXNmoPX5LbJHz
NcXSS3CsWUFmcGtlNqWIuScjo9wM0xHFLY933jtfc/dc7jmp8kEUTUgU9ckKhC1ChZtiMUIoY/Ud
TDWurFytq7a4sH5Wtx+m6iHpNNZ0LKrxMPk9QyPn/P3A74mvltJ6nu1ck9McuDkW6x7Ip9cQ2rzo
bSbYs+HVHnEttdN4AHCm4eEofl8r+stajNgCqXpWZbiMlJkazLFQlCroOSFdw8uWG6JrwTItziNj
CfDaiEPVIQ4yBo6YOjaktI+2yx+airhzoBEzsa1y5q8/oz3J1ESU3heHhs0SI7+Nf2UG8as5EN+G
oDr7SmNF5FZQYpzuu2jpbPwg8YCE7SY6zJmS4WLWvKiQ78TZkEvQAvHBClbWQxSFohn/MkVGk9FK
8/zKUViwHMli6UmC5By6ogFJKVM3CqAvCpp+/Yx12r+IhAdqQfTlsqqWeGVntNrMlvjhxPxnZMrs
Mac38/18ediyMoi1k9P3QYKR5JZRC1KnuQq+FVf/RILCQ1AWoQwVdqUPHlYYsJzAPI3BxUe3nHTy
sHkGHiN0aYDnfRaCEBCl+TTkNaoQ2FQ+YGli6+ZaC3TYPQo8FsN1BuV/Lfm/1Nqfu22kh30j/+xN
uSVGSxIpGkHHnOXoKPvnlyBQIukijJC5nMDYbRyzweqlF2LaZSAv2iDz7eUczsd+EgQc0D6BNtyx
8A9TANGl6BqbU3vFkcIO1WPy6T4QzVg4ywuIZvI7KTL/zHCWhFDGMZL4IP7HiEnhA/rwGhU9G35P
aph/Ezzt4x3lIcFS01sU/5znRUrCPUXw3hIqNH+mvbhF0Ff8j9b2Q1XLqBBJTT+5nQIhRZ88I16d
aTaGlTQ4ACcdypHFUgcnbwOTttLNcMgOZjWeJ+H1t8+YRjFrcgTEa1+JdOUcgZgoQAr99X4qrXuz
CqNX44F9GXzMKt/dN1fSii13hjUVNfx5e+RRSS98xISXUTlm7Wy1raPCccDTJILnupMddwD1AcIf
YvJNv1qByzNmncQhEvcFaAQaFVD8cBSU+CCYI4NSBS8EQZG4vVcoTvzj2GEpHpBKxs9mvjji0yJU
b7pQ1oO75HBwFjWgZQCYUzhg0NAoQPUpgshUDau2wtzzVUjXTwOAaDgPlQQ7DWDwfjlI7iXFMfi5
8rcURPrRyAJrU0xmKdUZ5wHD/E5NNULXMdT4a9+IlGjzr7UhRqtiSFZHKUpykVQchJKz/QFooxAJ
cPqhji2hBMBxSUrDkyakA/3qY/mJIvBxaASNDPNEGCVRFecx0HD2HS0Yyi2J9Nq5UDGJnl2OU01n
kiBGQJilfJFhkfDFzlEpj73bKDtinjgzcwqvynD81TuWWUmcPFguYM05ceK07fPJorEP65XPSZfc
+6zSBBERWtK1efHhMZ8aHP+E5MXyCkL6hRX9tGUawwMaITmml4J9Qxct8X3bTuqnbKYLKE4o7ChM
FUVPEIVcR5Q3cwQkk8+ierglEdMA/63HJWGIaqRR+oZlToyN/yJtamgDAgKF1IiKOOGTdcQATceB
eSFaoxQJxBbiCQV4bbSngwl6XfZZEytCeTPYemrWhxSIN2ZcXdzaBGfRZrv736U60MIQ0WwzSKnu
xmIYMbdQxSzGHE1x5tvgB+Uba2JuH3UNy5PTNMDGxYw+n+PaTMOCq8Q6uxypiRywE04Yi3LZZ3Gz
A9bfzql1xR2X57Pnd3shWcQaJ8Sl4498CctwzHdwInRFeGJT/9BfrWzXCok47GXLKDBJ/wDlIOGC
spOQlLfe7p0arM17vrn1XwW0cEYj7Ijp8Ysv+j/wDSxgj3aWRH/a48oH9Pg6b/YvCb5plgUGdvW3
9907vSktVOT7G76mja5BDWcC24SIArnQvr9aLGJaXhuxHHurnsk9Lln0H/JVK5xiIcS1jJerV2Ic
JE4COuO1wlrxCcatlaQzEbZoRXyRNsFaIJeQwifff5zfE+NXsqgSDc5L8CHj+juAIFez+Ls2NarS
vDtNxjFAF/rtIUN84U6XKKdhKFOFw/P0BK0xZfRhcV1o51MRIQ67l1VfjItS9yoHzHMOzB8I2VaC
MaCWMlaFSiON/XYFjN8c+ZD1poZyKNspMvFyGlxDU6/jC37mWxE+ojERpHypwfZroyy32Ey0yVdj
xpQ2i4X4NrWrlXvdrTXjPYgQ2LiOPwe0+O5vnX9sop9S6T2QHOHGLYeVPZak/Fij3y/OlGLLuJbf
fk8o1tcDquuS6zi7eBQCDkXlWxb/zMlPLxXkEy6D6XGtlYO6vT4BeZwpWmQFbQ2RXfoap7fEL0BQ
Wdfcg6SwEYjwN0ygK4wvs7IFrBayImNGwWKqouFOwiWRP2OVGEha/GDuUuIoVvGQRnBjsOXOftaC
r4j+mGbwl3JeEV3d5mqFZF47/WaEBwE0nU6+Qa+YRiQS3HZ63bBPLYzA5CBKY6EAAGsmG/m06eea
PABKljIPFJ1WSuUnN4wuVUFpIIAyrrtYLenFjI67aJZmPc6+j5TB5hgG82jrwUpVRozNqTofvpoN
V3SWZMe1I/c0VTW/MjbU7mprP6sZWKxWfx2awqFcy971+xxjKsbrAUMhGfX6O2kaB4Ia+TaiTGKv
ObEoU1md7bfEylzYRrOiU1yvauY7CsppdZoAwcMyx3NEKrqUDxbnfQ5JLYLW2kbbX98X2B1Q9YvK
jfE4a/JzsTv6nyyijIcnXMGiAgrwlSbEQw4xf/Dd3mWnnIifHkf+BW8P8u4aRUcIY9Y3JU8Y9jCn
UefmPNw3SQvd8yyWCMebuins5bhZ5XqxBTZTIsTS1Fn+in3qOtF/IGr9X86EdRHzASAeSggcyFPn
LIm3aU6wqlhUszKcZYQSzIb6DQvuIN+EPMilMKcSlQguzS3Jz1sD+8ggJeH4XNr0rYoe485pFyHm
8sUaib/5R08WYuHM2UEjluveTy4oB+ts1w0gND/eQ1pfacngf7Gj+6CXVa0jzdJi9gAD0oNsyWld
L6vsIeumwETIvP8uBe9nb36cVgAToowhixX5MKPeu2Lhwlh16FmOdmukfxP+v1U9NtkcVftghO6u
P8iIYykCNEQQbB5pmMm8xZ43HNePcRCjHpTyWFF9jwmqfRC9EzA8Hl5xwZOPCG34QowOK+Miyucu
saWcj5+fuSFQ4RkGCvpBzfsM8ZxF0AJabbKiyeewKD0E3qH6j6HxosnEEYWkY1IVh3EVGKWf7cWI
jL6Zj0T1tJZ2rME+/PCxO2bqIzrQ/4snKPZIvHUUIfyU3dJKU2FcH4paif2Z+Woe4boknADZCnSN
qSFALAm4Zp9S1Wh3ojy2TTfGcfyKVYgSfgi5Zl0Ax5oP+Ao8bB93R1mcFT3n4UWW4d7PgYXVZK9q
pIq2e32I9pAPdgEQfS3pVuVafXS0rsAMsTlZSQM/LJJ0p8Y9pXs1cO032+Hqbnr8JYlJ7lnEQ4FS
iBtGqVt6NwMtCONDNXHxAU5A2MNcbyDmGVoL6rBcUysvdEsux8ApcEEsDYKm783zwhhaCUBSt8Mn
1fcezsenvKvGQ73c0GwmH9/oK0nYU6wwLpXhDCVns8TiH092iaC/Qjj0j4GDPNxoF5iXMF+CEJ/1
baNJ3KcB7muSyrsDsJwSiGCpD4veEZDZxyayC8DjvfJa1accECafuh8pm8IGa7Efk/UxTOPAHfDK
b6WXkBx5mzqmQfjDz18S+2KGW6URtlkUTYWA90nYig7oFHRZJBqn4IxoMrHB8HLw9+ODMxzCkr/V
wXqgdytqVROT5BK2xVG1nhIFD28aJpvqGe44XryyJNsrQGypWkAY0KWItc6ALVePgMp6AO6Jje+8
996NBXnqdZa4H8XpqCe+Rdb1KFrkz1LQEmkzcWcnR9b37PkVGi7w5f8XhPSJENL0hvYB6stzjqup
/IcSAS+9mvupmhh/il+LkofZkFxdKKJ2n4i4cJeNuK6siBjv7jvpalwdYCoNJxI7o4xs4+rw7l+B
iezIUC22AcgIiaAy35DLxwSZc76u/hb6MBFBDvUNCJc4bOXtrPU64d9uDu4B7LGt5UkFpnm5WOuf
Dj3nItKeTc+h1yiOTO9p2BzgGPWORnAecuKiVtY2nIyYi0W/NN7p4r+8lKakx8UjeLYlQWQjJWrG
DY+PDFXu6yej07XGouO7k8YgkvOrMPv+D9ObbGfnWTL+b2sO56Cp061LnfXaDlsEDC9u8QgT38h3
4ItXc9Fbdp5yEwBx9nvjutqaB0kB+df707JHi+MNvdH5dOy5E/L0uJPtwHrcZfpbJehVofCRcgiP
vxwu40e3yZNJcMrRorM93CzmJlEpsu6DgC/2TB02DvfTD8AnSy0V/etKn4CfOJlu7dt0qnJtepF/
tGpnqS41fj0rnixvEZpN8+7ZSSyd9Y6pq5HHl8eKUVCULw6ZcR19ivlsep8NZhyolSw16kLQA8XG
HzLj+1oUzjgpxOaqYy8tvntxiqaLCRoBMxR8M+VvKtY6/UmAcpXKjNtwLkxlLaF/5GAfmYeDyOCq
jqtc2pqpw9GU+NMdj6SwzPbHL778jocKymEnpapvdgEz3R/1nZiuVjSUwMy3Wo5+su0/2XXX9Pxm
ov5bCTlegaW6O6khmNNGGK3lGcQxu2VakkSWzzYRpqcZLuzl+cYqHgIqL+wapnyxRoSeieiZ+bIG
ZCiWJwonL7wrYRAiCi1HJrOAxPvAz8Amk8IepEclYOjnWI2B6zJkUrOllkSm4nruBn08KYq5sFCs
P21H8LCivUtn6e66nEmXkXk+FtmsOl/t/yC4nPBJpluvLFp88WQqEQEPZFLOjUMPq3DnMcZvzl2C
Zg+J4eyC2GcrsJKoMxxB8wpHO8D4YIRibrX4Rm//9blF0Va9mNMOxLyrgqruGWWg3hZ51AVRmynR
eY4XpEfpzUBgSdVDNCjKopRaZQBVJl+4/pzWRmJn22xWI5MN69FOEytMHKhs3oVX3ffT5gnfvm3s
HJ27RqOyLzpl/lsbwZcmMRoLRPGqBwALmDCkSriu6CMQ6/AR7Kt1d1PzpXdDLi2+we71vUWYqawH
Sta4JKXgM9BioOiE0uCKaP4Gc5uxPG/SVBZERD8Wvc3Qt2TZoSOiS0VhW9neO3m4ZMUZjzui+71s
tUIUW0YVDaZf5FP4s/5XeKHnVHSpXBttS1DnFcxDeNqq+lnsDZlNUVUbIhwfj4vYCoqPyDBtCBHd
VOTtZyj4viODMz+12ibjRwZp5WEq2+mz/9ynzL1J2acpzrc2t81b3BSaL2JOQ7eKUkDR0yMvieJM
JJZ6y25ljjz4OaPnPiv4FD34dgHm3dVUD367kSrBKzrdgGEL4v2SFLn/ZkIqiHc554lrwCwUDb46
QRmua1oOF2ijFuVYecly6n4lnV6HWVZGknGYrfOrPDgA0TfBO0MxI48d75QYjcWCJn7bN22jymN6
X1b1OwR7Q3c5xJXuC7cEdht66MaabnR8FPa1gn6skydpOmQNAPEC4FYmbJhVxE+Og61JCWEmqSzU
kxjwyt2r9rLRtdEjoJVPNBZS9kNoCm3NCCrEgFALspEqioWNGclsNKtLZ2BVm94XOIy4pC1goNyF
PsalTShYde7EkL8HoLSOzaORqO4o3ofvt7nqPYQOnLcPd/wXFTlnqoXBTDJUDpEyQLxz8yvPuiWe
rIZpgP66V60T3RT1cOJL7OhJjH2T71iKQU2IYVkz3/N3nHJ6vX7tCrz0zjJI3gD97pcR/XYmiDW6
NH5GXiW/hlwLjklXztPTxqzLTdMK11taC3QPeXbROLC80noQhwJZqU3x53egHywrflaXyEuJFCF3
LP2+MRz6RJqWDTcCZJbAO6hzVGU3mYEq12GUR4hg9ctgheDFXD3dbL6CMIWk+rBFPsoe90Jf+AE9
SiKVYaVwKbS0IcSIIgXcsnnTr9rR4zaInZVHAHY+HQRyEODV+7jDWkyID7zqjGGDnnjfdarLNWdz
30joj3zQ5qIvIz8mp8kY9ccXmL0nH60zm7/6nohsuXdGAEf3DMQY4WIpxue9TRlTNSvYiUFlWbzH
oo7/mXQ5M+lTTw23dDy3IIcIkVkol03zPLOLgBiTzR/ggqrn66AhXlwxxcT3jERwjgMiDhq+p3t+
VbJTNlShDLuVNPCFTSffg+aEdNtDB9MKluM42cpy7HINPwM+OL9NFqn52mklu324/1nSo8SRuls1
FV2bRkgM+vPHHnS4PrGGXASQqcmt+UArADIsZRXOQDonK+tvY7/8FjpfChb8ZE6+ENBqzOD2I0XP
O6fEgd+qFPOBClwbnq/XapCrfPCfaFK0/RaOnNpJ7+yr/tE6sff1I697XK99pjgWhHZD6cSN+Rq4
j0SiZi5/vOY3LLh3SMZlMjb7oQB3CnsJ/SYFxPuiYpB7wg0JcAPTuHUT3UNp+W9nbHbtZYGVtkFn
MExvm44OWX9TPtuAen94Q8j10TRS/lx4Lbq2i4WvgXdK/S5NlC/TZPh9ROsae0biY3/R5+6g2xXM
fzZRIB7eRoT4l3sJ1fq+LbIpzAW9eR1VipCtUWYVdrW7ZkRRlc5rgL05jMoBxm6STFkczdOWBvad
mFvdBhDd6fCUr1zRLrJ3PcOqjrZeNxo2GtSqcMveMYyBz8ggXw8a1/LWaaFVrh87oZudIyqofH/l
qi5oWrWzrgAcEynVfU+LV18imIb/fdKwi5Jxs3nqACoa2HH34YFMXJ0nq3V/x0LeRAJ7RurHOCZC
wI3UCxUBrT9QhBiP2n811Ndwxs8udd2mUuaZzRDOuwzZMWTeuT4VtzPwyB008Dl6fMEi0n6Sp4Bh
LRiDy757P+EBp2++RuPTC9CqcJcnzPgfNpg7K9vHtmk1VFazcinliF9ZcWf6v2C5iw993/AW0pav
b2ExdiJRzRIQnJCBT1IqbZdDw9IelNDSl0oVrX5b2okfqn16YMJMXQqUxcruccerjhkqFFQF9QrT
zB5tzU/VFIL1lYJ/MRFBdrK9QG7pmjNqDoFOCLf/wfLRGa5XprO8reLwE1tLAA5+kqyCxjy9p6k7
lOcvKllUgnuabxs96yxgQFBsa87iK+NuWOjlUhAp7+F2LnZFD6+jw7UM9L8XkSAVKkjXdieVuF7V
eX1Tk1DjOYQ6YGv6V4ZnX6ixa1sMfHMBbc/+yeTzrj70adhs9Cy9j0sC2IXT91LQIhMNtnsFfIY/
U4OGBIQl/BAiHcLTp58MsGaOqnFtm6ST+tBGdiz3LZTvxhRg59laH/Z8ipeCXA+g7lT3XAo/ZSk/
69IwdzmZpuvefFOBBzZkg9vUZqTDQpSVliMKTLKJ4DyZN/djVf8oC7XOEE2mOQOEosLQ6iMhTMGE
nfv2Fwl+O+7ERPPbeKkhnHmuzHmvaFa/VatVZspE5EB/hsVN9yZQl1GJ8PlGrKwpTS61S4iRuArn
yKrDXOLDdlgbpy+bFqLea4ALob6IBAwxp703UdeDTUm2R9I/KMIeY/+aroxjJpusV6kI6n02Ka5Y
YwPcmn8kBNNf4EM3eU3L22QLa4a9P6A2Es9uLCU4/S71l8Vpj+1dHYSUNkkRL03U4x89knNUHM+h
SWpYCormgSRJTGlmKY9jBn9K3aymCXRJwIudRwc1QAvORLFXAl3kQ+4KJZgk4fsUp2Gdyv5O2u22
bbD+NdmCqyVs/gMy1j3xT9fnO5FChLltKwwSkAIRUyvh9hb15xbcW8zy017RwRmT6LmANKKO8XEJ
vbNAECvbuEflSMiIrIoZq11fLs2bw2YgG4ebBQV5r7x5Lr0EuH/wQ2ehvMrbXGYF++F6JgOP5XsG
vui38nR/80uVBUTpHlmdtIih2zEzAt9pCyoelKBlVUACn0/5eco6a2Y/Kpf6dtKX3yHG7QUi4+nS
AspJAsZLnWRRRMEdwHExrwmtjatJOelkPA8vKNTGv7xjdZL+M0QU8/DV0f0kEwRr0y/LajfRHy0G
NmRAFvoVnwYhDDgrclR5Y2VAv17bJBdrVKGNm+HD7ZKlQV5xK7xiIAjCRijFkfZqCY0Ey8xP8N4k
vPNsfr4pkOH7LKBpPFqG7HRSiixvRHk6nHwH105w9IXPbO/zhV5Yr+x3xZ2a/WY7n+RNpj3ADTo+
GlZ0IfgLv2IN8Wo8T2VUE5co2/zDt2Q311C+XwfwGLKWgsAiedfzuvKhpsDxjWFrBQjuicLoP07y
Pjr1W1hY6oCIwhGCJB2iR3+bencvBTrfcdpksnamxKI4ZzorycWDUXtSgd72xLvHaPekLvD7MyWl
zA+dvykhBmkoxcACjt758n3WdPsG2Tpqc+Ygckkfos30SCVSnF1LV/zq9AQ3p4jKhJf8UTcuyUCM
bdrHjF/kWxwguXxLJNhtNN6QhzOXPs8JIeRH5I/+JEgSNYvxlg5ilR4lHs57CHdcsGE7RoAzG7sY
8kc65VsFgAsJJVUhpjQWknUEdIc/i/Xi1DGuJxvDVfmmEl7twVtKuv3fLo6iU9xvmx4S4johdzWh
kTBclK5U2TLVGXgBHdjo0lZS1iDSTSZD0btG0CiC3u/dd+BobtQ9bOOozYiY15gk14sxEzDZA7Qa
qHl0znPjK/nwL96P6Wx050thzjUvqEO5vbmbsH11yGhQ1ylBwKZKeQIslQMicdGpHjDrYuEcFZ+i
+MfN2DXq0/VP/F30MmISr3Zmc8WpRGEKPJQlv/srtOpjii/Nbhx6St7j3ZJksmZVflgExE1WcxYH
uRaqtDB0QpMomXCYRq7v3SmTYSW8LuRwDgw0Jzu2/AYJL4O21XY4IPBESXtdwgfOjYg3kYm+Ek03
ce0XoAqwiuWN4nPbWk2zYpTrxzcl6HGAVrE88ccz9LvHfHA5dkcCTbai8g4DWbDLMyrCUN62p7zA
4nB3PVGOBtGwXHaCIkClyeNQkRwvTx6TD2YuqLEx4JCWMVo+FqpCKET8p0izKmRBfPfTdjT+2hPY
B8Fj/anBI63uaU2rHpiXcvHYoaKpnZzJA9J0j2Y6sdv+PnmQDBXmxndCB8gpCGXpo5clLVm2zvRM
zXEQpdhZp7w3A852rSA2UNeJ3huhsO5QDQHXmHro9bk7UrlooezfikKqxL1O8Nw31jiVTkr/77in
oXk8Xxbo9lvLP/TkIia9TnfIJb8EuhwqRmQdjtM/nds+Uz9zb8rAmSKFplrSI0Av4IqTf9WLhSKp
zqaL9KgWOo+uzEu+RRez9AwwrHnlXlWpNUEfl7lQI47qzNeYSZJN4lIx6ktTbWaiX95OEaaFLKcj
RAQ7nEoiIvT2eAsSXp5Oaxga43QpI6yPFZRpsk7vBU8XS8KBrBan4DgRBs9fak4vCtLBFlKJn77Q
6q/CtMEk5AYBIPYw5yCp6FM74v7dCN87dJ1+StuYKrur8K65JDWeP5CORmsrFeLFTyjeK/vH1Qz4
JsrfUVEiF2168bAQ9cvGYBRctlFZK7H7A8gy4yLRcEjBcwuFu/SBcGypIz4ggACzx8raILY9xvH1
xEscr0s9sCik6fECiq3t5Dm7BrWODxUe0j08dSlgwT/qFNImCfFUyP6oUw9eWmhvd0ZicrYNCmrG
/IlhwL85pIxAeku+vpfL5wyJ15pjApXiX9UitzO7w3cE6J2fcz9b6EJQIbGWJR9cCEB9F3GE6EPH
JTIckQzakRY4kHpzREt8cK2iCWpkZwIlf8ewKWhDkqmMopmAYR8RwrEaCtoqdnt7sT8mFA0vyZP/
S+Dwg2I6nkfUZjTGNsB/8BPAbDBazlPrRIwsbPQJGWn56Yc2aNb6KwQ85ZrcKzkB0YxCazYcqMD1
tRri2pdY+yBETPPPixXWqDqFKfCh99v1FPe2uXHz9Tn0lKaPNdKborBhVZBH0XqDdMD8k+lsfN3E
CWfKWhvW3A2kRniskZccbFf5b/1CG3vCaMjOIE7rwBvQ/W21FR/DNafKqSVHN4SxSXcrjXt8DIcO
SWhlVox0eqESxLBj1Tn6duKbo0zrEszWJ69enNphnUNf3cbxTk5XWG/b1pc+YHW6MjamobnK5SjG
vI+WO1mpAJIq1Z/K+UU1xQrH3W1w2VTMVYfns9D/jdTRzX4gn+FSeqtfe+rDJJz50z/HxGjxoYUP
ThOftjOTtkPBATMETmvbkOcx6kfuOStvr6IPAfLYzq3OZ62OvjmJGiXk3yBvlorXzVZx5nkigyqm
xAGTci5xFH5DsAIAXB9bdG/PyDbEQjecodiNBpLRJgCoc/3gbIEZMOuh9neAHqkyhEk8rxfukE2D
/WhJ+HUgqOqEuPKLzPXEfrI1HfhITdgmYGsGjdFwVSBOQrAQiNfd8JsgHjxC9teH3S0aaU1ksv6i
kV5mXvWHwDFBv0toSaKyFCJvQ6wrMEy8OhUmbECAIlU/p3/l0q+XzPDBkPz5vhDKr6KSsQG7FpaW
GBKuv/+cczpFY0m6guXA/xYO39+A5urctkmU106Q0YUSwTs7rK3NlcMhjC2fmUF1ddRgm+Snyg4y
oMntJTtobR42NLnXxw/3iP8Hd9PhyE1gerTeU5wpEFv3KDqVnBh1+XTjCaiE9SAfWqYZpv0DEabI
QuTHtuVpTesTN2KExPrMZET4lcxndndjE31zJLz+Yad2LGsjF33mWe57lHE2BCQFkxTz8CXYLtjF
3XXUpP2n5IiEQ7EZmMzQ4mxwndv87b5w9+gi5a39LoacUkPnkTyosOMqrZ9O+ZlIWOpBdtPR8UEu
rtvArIQlT8pDqn8lPtGBGDJxRr18zTdlMZ6TKZ0Nkkoc8yhxt4XfJKbG83FPgYRH8kgPOvtmzMcb
RF8POIYcZ9UD5qunz+8TAQaQ97n8zYvJKg8N6KB2D6oZodDZbunguAYxSt74daM+EnZ4+0nFhigU
ALuJRRioeIrJ1pUMxhRo4a1q2o6NQDYRnrdsB7wq1/ekQOT1DtjiCMm8Gu7Eo9cmNfl8zclZlfKB
I9GZgQQUZ2rl9GnwWSu08ZmCVHYExabYK7P/mMcTnZLK2uAv9gNb3BVeYkODLUpJpkBH+PS1NNOo
arOnHJazm1mLxsSGchEBVd+zbBtn/fH9P+jf2OHzNwKRV7OPmYvtOAUMv0KjDpkRRaWY8CnWrkve
V4BLiQfz1SBg2FjRMR/yFUnsIQ8wEkJQhfdBbtF8TKMPimJkiwUwMi3ptkRMxxsqwtFcwKqPLi2R
7LGLM9qCQ6ngbdmJS5Ytxc38fCrP39RJPwYIJHit19PUh0Z8/4eu7zhNG+Ap+kgD+gUfPefQDcz4
ktoAlpWExb88L1HbaX4Y0oQsQTQcww2z4bFqFN4We6Q92LyrB39QxSQCsdLS7hfCEttCMcRhgNwE
UfBracbOFlgK2+ASmhBfSTEL5JXjvXrn1ZMi8GbWTCqIkM7JfptXsEbNfFqTux6g4SSLbrpytsbF
uND9YYgGOnAkU2Ge6jwZRBDHA4yHvl8fmtfVfq1GK+9FsakljyQ2uecE7lZdYhLdiVjgf6ZHYHFJ
c2EMMJuk0wqRZRtnjxAyOcRLY/oh0vRY3YNrepzZepVy+MRXhHqoshEuYI3Dq+SJEO4ng1V/Xdkm
jNakvlBSIX3lpDGbMMzrThVMLprjCxl/EzD7fNIk6T1UmINsJaGfk+t9mfEokwYn+iSH+oQxHNmy
/sJRpw/5K0APQViK6AvXussrT3Uz2N3mxpJ4KiVMN/6E/zQOFqreXSiqpySK2Q7rc5YDDH2rFc54
zF7NFMd+qNlBDSQACE4JaGFyMyIZCnoKnN2Q9PEaGxsCWDZe6tuXZ6LFYivb1L/WE9wbWP3rJRWr
5BACuKMousU88OS77HXvcYJgA8w5ffH4OsMP8sq4Im0N9WbFWbsVdG1jLJcBlXOSKHFKlxqTNw1E
yAB1pgldJWHNXqDqZcnaHGhk0BiTJrg9F7jLAipBzBa4IfeKClqdgWMIf1/mLxrl0xWgnupW79WD
pdRsOJ2IBsCIbOxuMhA1e3U+hBRsJdemY+m1mR/PgyctFNsexttb0o1SuZcGJwejxzlK/9aw7AXA
Cc85KOo5DjNh4SZ91fjh50hDjBnwzrZhNzi0LlQ5+7G+ImYnIeQaJVJL+gu6EZFLZFRCPaGwFVsU
ocBCdnfI9PGWzV1BzbMCvl0zOeptPrF0q98Le7DMqEclZhQBfx+yAW6eLOaK27WKPh3UvDCdrGxJ
uegxFOp1SpZe89N7O9PQ1BzIDbFYJDg9HMvgt4fbTcSFFy8Qbx/ecudxnVbo2QZw7PKv5Ur2fF/I
h2G8XgvsfTmCP0B3Am43XlTek36Y/NuRaOdYKEMBn07ZQ1GCKe4F5onO/Cwtv9GTveonhVvUhjvp
eQJiBa6sYNsBljj7AuHa/de8WJjtBFF0b7D5UZVSM4Q3lr/rBDtsyIrrMwd0g4Ti2gIq/GCZREme
O2RqGpm8hRQ+B1W6JC/A7NVx1PpKEy+I7hBtCGksRZSuQiwjTBAJCMOGrGHZT77BPXbfvKSJky1c
s0PZBWKC/66C2N9cIRzbpRzNPtmVpOL+avxtIId2fS6C2tiVZWDjVhhTCMixJy3d4jw1YocJGFLP
k6hHl/v79I3CnNRU4oeiRl/ye/cyHJCNFZpSinMHXxWEKu481WFopFR4mxALxblYIT2cCOR/rh8G
S5TvNDurc3s7OP/DfYzWJahHDGPAiJT3dRh3fBV3PDsZJxcNwF5wa5167qIlHUpPGm9YbcSK1SRg
8yxKpgxxXByR21Y5n8YSRIRo0/twVZfJ5IUcee180YIeE+5uUvywCbk6OQ8xVyLCt27BvpWMneDe
67Kqs1OPSTQqq39OCaiHAm7zu9QPPZaCpOjvB+8w7CMctK8Rt7d/znlpmRvGz5OmD+9sDYAwsBss
d+vIRhuFYrnxmt9TwIK5KxvaadgON/hwY1hJsgtywCjf9g/ZhmRFKLg83EdvV3+A5l2Qkhl5GKvu
HXkVN4u4hMJStcbY3nY8G81I5aC9ZR/Avv4OQCGWINoU2x22OhfhLcvtXobEZ5TOSuh3JaF6QoEg
C92/urzLDFN8Bk/0XvvhFG31AfYokAig8Aqxl2JXFHTM8cgK46HO3m+WtD9TMxyM3ykjOOrxP2Pb
UXvlfegQSjNdIdvCOvv65fropDUlRGAxrXeq4EJMmjHJlouMQvx1D4EZYXZKuMSF/KjA1cID9dlx
48jyOw6mXl4pQUvgNXMfwzXSIWsxeMz7wUskalg2j2ikibh66HrzTmz60KLSrwWpRbhT/qSednoY
Tl3t6GyJhNvnBAshsY+J+Xh/QhGMzCa5Mzn4p4hUSILimzrqcFETiW+GKuSwUfv5tMNgG0GqGZnG
w9bRhAO9MCjSwE5/5sICikKjD8AAg6T5ax+HvM2XdeuIxlmdeaX7jrHSAH+Mp4bMYd1KgCLr3Ytq
icKk1nZdmAWvGdP+ZBe3PAwEYyTWPUn+Ta6bbAbfN5jsJH05GkrEXkGUFcfLVE5EI0K5DMt8yXbt
hfeK0au8/8t7NSZJCcVEl64Tpb4YuDuFn2kF+1V8dsDZJhhmpqqYQrE/TGnBoiN4ZbYoe6XgAjOb
Cv48oFh7jiEs567g6JDdVXxsfUWeg1tWzztw/tyqdCJmyjkR7RWeIJ2zB9mZcUpXv9IeMDcxim8Y
2ntHn7M4ITYblffst03ilE0FlAgomXIF3PXLJm2EOnzc3iYr9iGfz4NqODvrWex6ORCkpPsYJaJ2
8Idz/++UVFsyMYHUqCHlvzyOj6/YVj3MXaFkozJMdzvBB/+OI0rq/u9dAbDwyRs1+mJ4uarYKh60
3Qeq6BJ3gwSWxCK+m590/n9rFSeJP6LySXPwK8vOVJuPWncNQUkKxRlE66gHOQiMbmgIdTV6ttAg
bxBbA1yUolNd9UpG3W//B/4GnhkFkspaQpEvr6Iw5r8oqWkNHueo6+HPpyDy0LtIbLXIx77aRHXL
R+3zY8vzeKjM2gKoL2jlabBCDFakbk1NVF5CH1wKFeAsrRZAXQegmYAymfGQ4TrDX7sQxzEQXpz5
I5QxW3W4pUyMx8aT8n11eZWcG7BKciOeThJYFhKsmvzZ3hBTK3/CD2O9xTRcjCZfWrrnKw1k0EGL
2X7WVW8vlSx837ZFtER9mzR9ehFHM61rX0KrgKYBL+WBRepIy14/ZFnx7zlqzOTwAlgMkcyfGfIf
V0eJALL7aayLjP2B6+AX+g+HxXuAuJ4bjdDoZc981L77hOcCYcrzaoJR/jLJB5n5lDmG6vR7Cz3n
eT7x4DGEV3tp7gx5MX+HaLtVehsI2+C3bOTTSJ/P0u2yLkIFObyHCvnuT0AgCgU1TsdJzFVLEGEL
sQ3bHbcfqdxANtjDORGjWCeCwrHoANq7y48oO4lz6Gt4prga+WKaWCdIZ4WLXhhGl1jyy3D36r4L
nm4VCx+qxhxhKtWq7G+Nj9lCc7M3dRbTszc2yuGFt+osqHInwYKB2ujtqd1Wzhc7Mctl/HuuhD+C
Mv+UTTYeZNCAKQ1MctNStHGxE4gcHbgqg5pBt4Soy7EpgObETIqI14KySxhf/ohxjHaj5M5rrBXE
P1fU9O8nZhnD8KtBAtwLIhwcWe3xt0mXXCKIGeoIx1BQFOOh/H/94fGyODTfg0y7LxEpWSSOm7Rf
DWmqyfCyOi8IRI1bgjvHkJ7bfhnRK9ezXV2XUHMByM2rX2fj8RaTNcFgr0uB54aPcFSDCmVcIjS2
3GV1YcBGf5OdGj+Ol5dfvRkqj302RNBkFwwwmfv6J75/BEXN2Wf1q6ShSdv1cZqzFis+3Pto82ms
dneCzBPpO8jtDswafdf6uDUVPa6G+K/1M6BtVNmY955zW+IqV5slb8G65hWiWm+HRiVR6fH7tEEw
Ap5II1wJEdUPFAr46ZAUF4U0mqW7JRUIyrq/clNmVR3jGTpTmTVo3PbXM44xhcS91AeJQbcdtLKU
FXiNw8H7Ql3Vz8H4Znd4zsABfJo8T0CQADRA2jW8meCZQIazlWNFfeqDNC/Kvb8saM+flC/KFYFE
rzxrUM0H/ZBcRqih/S5/F1AmzefF0mzCAgoc7O/MiYttEYVvnhqOEswOspRjoJbDGI+zwCjsm1pQ
n6Asl5bRY2S3R3t5c1q7pc5kG7iVU61CW5ybN6Rk5Dqh0zYU8dhMlUWLfEIVQi/3XSMeVfMGN4mx
Oq8LOCWDdsm/3EiqLKIYMbayj2p46r9R7T0T1iLR9rIPPt6Bqz8MqbUCkuPK4mtDHgvGtnS7eKl1
xSs+Hc0S0xzgD/yF5u/pgr7s0m1mMdlIa3la7aLMwCfR6qQbLUPrgyvWfHLSiY0jreZFD1be57hQ
JZz6ugDpLHz02nRCwIYXS67gItl/PhLjXm9ZAT78TmXXg3PewRbHM1OjzSDHE6Nr1+Za9TIAvYxi
2Op7iwDq+M0kZIttOpXwfshvSmZHhkiTjwzGFi6ZeZPEBi7VFs2/o2hrcQNemeXV7nAHn+V7Hs4y
Vex3jx0d3UrwgzSjYf+Qo5wwCBCm2smbfvRNNMU2Odf1g/WuIlA2LsBWK3gOr+7T1bjCMy9xBmJb
UcsQACiAiEDKjD5eTAAuGG1IfADb1dGwuj+FRzgymGOimGOGZz/eIIAsccTaSUZEnexcfAIUrqcm
PgSP7CkyNVk7QQcVCI+QZvUnquLeBY/0WsNIEYAoGo4McuzBlQGtlrtS9yrH48VOyhBih+NqvExI
weyQPteV3k0duXuAUPPMIOX2aoxzrcyVtlGCUIU1VuMvi/mKcN4sPA63e2N0Fj/pNvcBVSfnkxAP
4OFwX5Cqh5G6wmkiKGXvuZDPVUzBJJzCtmCrLxfzkOus82/YG4PvSZkjXjry79poJ69Yp78yCnGc
QgYPSTR754+l+NvzrcDxX/d5o6YO0YxAPzaZoKEa1uyPaQq5eQ23co60M1eIXRiGIGtvqXrOaRHq
CLM1FZstDsmwlBMqROeXk0hoEbzVJxf58+F/S1gii4AH6HnkuMKlfRwrkXC5+MIW1dQCTzOqSVf2
1AMhhKhJSHq9Y3rsFhEIWfZ+2kZJX0R8i2RJnFd1vUTS81ZmGCStyXTX8S00TaWbeJvRZqD/bIHg
369o6Bc4nhb8Wh6v/drbkWXJDzZ9yVmPsXDGOVy5Dstk055NcaVgut3O19B+NFlF/P2Liw5W6SR/
cKIOeUTr513jRfCQdnIf6VfI5Yn3OtHLb8DmmrSoBbq5PGwjdJCvgNlMYaFRQ9S1J+Hoz50X8kcX
Mpb9WYQSLV2nmQEKXHYtpewhSJlqhblTOMpJxvEgF2CF2QtH4IhnkCHwnHYSqLfdEDfFer6LF8xz
387voPi9ZIxqwJqZC4HVCPw17Ss5tnBgTKDP/d3XI0iVH2h4qn1dLoEk90rtQawM8vD/MrjuBxvL
dthppFcUeOFmGheSDpM4JfvFfvsqlFolxmh8dkCLiDBGyjMtRZkPPp1bdlDVKT7pSE+gZMDHrPP9
Rz33s2bQR5pNOo9fUqb2cMQ23JR7WbwpI05OlND6FaBo94h5kqpen7sC1L23CrkbwI1hEs5y1gv8
s6v1E3y7Ur1Lss5GmV2rmmnjRrRcTOeLOx/5yTTu1hjVLtdU+O6hA5/43ZFOdFCv5HVO0PumXIDR
lBFwPcbvfxUPnwVZ8nemzyPsVRmQiY0NwLY+hv3AQaPpMmOYdRLp3g3/xkEFrFoR+PBsII8hjUin
U1BNvJ9RNa5u6l2eitRWoFw7/HTvboSghp0tk3zT2m05ery5Z9mmY+E78aUqCGHChd6uZeTjQ47J
RLihkb/Wzi2+T+ZxX8pbMpzTVivZKBHbpYkZXxDcv42ZhgG0Bam+ov5znQlpqBs2iAV2lAbVPVjk
KCdYwqTLHQ1uZPLJG153Qnpbp095jXdGsooG4FCNnNVA5CjhIOjvCV1aDytHXAurKwCyv0wb3SVO
9c0lg+87QVuGsHs5nMbZ3o6jiRpsPZi8fxDucWPlSJE/oevu8a29e4yIHWQlXLlvrijwwP/nvPvR
/6VxqkN51QO2OKbHRqEFl9VwztvyJzA4OP0V3IZEvkVoUa9Uw0dCMaD9cfSv9K7PeDjluh73jrPM
M6MlMckDDE3ziu+8HyhTTL4YyEmMqjGEwGqC1L9EpvPuvwXaeHRKokQyuJ+vbbv7qXLmbMPfLJch
4K5QaO4Ui91vl6mw9SmdwmwzWzIYBqcMNAR7VedmqfybVW9q8cmcesJ4svwL0MCfthSFhtYg+P8q
xY3NZpZqa0ZyW5Jhwo1aBglLYOXZcPdYOQ91/7FuplVPMqAzNm+9o39X+6RlGVyr5GXga7pu+LVi
/kuTO0M8PYGb7Q0x7Fnmd6d38/Xw0eltfIDIwi70qOpIEwx3jD/Q68v9gLjr68fzfCzW7mGVnpIH
328Lm81Boc8ufNv83Y8cbuNn0zb7G3DRryQSwtbrWxrpPJOoWel3rA04/tJoQqSalTj/gaMIILo6
ygjtSw9PXjxCsLwrOtJozw3emllDrzpmSXiY1BZ8LaAa/Rj/1zERsCHGf0VjuY0T8QJvswvoeLhD
HPVajbW/Ygyx8Ik/huBkOqdG2nWiypRnj0MIid9G+YKp8KXxHFM5DdtTS5RnCnpEdSO3/h8HtYEx
d8tQ8ZSv5LETncpmJjDLkvxdurgtfTFvjbknbRIj0EjKr8EFPk9dGO+YfJylhKV6E2xxy1HwrtEK
a2alh4kiAJK1jZSCHi50VmPswS92T7c3w7uqSnN6eiCw9l/84kyhRS1XCkitHUWuJ9DaGuKQvXuR
kSIgqIJ7Bt/+VVx/hQvhSq/+LkvSOs+Fav/CyND0rZLwk/4OVYoifo1gF7FRawE09J3L0Rn8l9EQ
+jMFHT0W9tXSjXXlgUwrGxQMZoCuS7h8kQWy7oQeFC67H/NuVHZCZxOd29/1jPINa0v5gkdlaUua
Nj8LYSBcdG71v5wKMqmEmu0W8D+8mkCQqKcdMFidh7dSYaKb/hcvfu3kW5DdlxJVCgT259slHeLn
FVG7Rv2m8vuJ7RpMcCEKo1ZuZyofw0rVrQxyr9pvqPmwe6+b5tZm+r7WqYzb65j/z67jp1EUcvrK
F1sw4RbI7G9MHV5HRRmXfIHCyoEhWoq1OOMz7ptwgldvQbFz2No9bgBKxIYyNFnBQtkLhp1syt5F
KsMDciaor+OflTKsminw4WtNA1qGrlPDspUykY0h4OeIZk509w5n3suTLVjvbrjsAtREW+IGzwUh
FXzj5o2iJGR03+CK9vmh3ldgo151ncnIcb1cj79VMGMGFlBM4W7+heR68jnURPy8FyAZUqCwld6V
wHn+CzXE8Bjgh0U8n1fn6vGtxrJkuCgnIKKxTbEbPScLzGGRssBumVDNHl4NE3mBRWtA76i3R+Av
cKgAcREOSc3lraht2mk4aHsPMmlgb7PX4udcup1EWUfbQwH9qFFLfZSs6ck+gpvjQViOk2KXd8gt
9fBXU34s2SiwYC+Id00/hUqkK/3gAf+GHwxHLyy/cg+UC9iBjg9aFqjoEwO3P1+znE3wb/gnnneU
CKSOpTvo3CEv4jF0ggdub5Cgohnh7HNkFVn39kUrF6PKQ19G5YuMvgNtq+zWFNeg5iKtz6Vm0/In
6peeGxPG/ncIBppbvUg/EIQ8ZOvt/lpGEIoWtjTiQ8ST8JS6UIZuo3v8Sn9jubMZOLiHZF7bgNHs
fAsajNZtR+zxya39cw3dIZ9lP7QSGg8leHj2n+WcQxcgkDuBTq6W2e4RGne6lxZipoYPU8HgXAk+
ADExY/rbH11v8j8JvF2HHKQfXwTKGSYaE3WPA9wyYB2yq9US7zIbr+Ng+lRgwOFZ22S43HX0zGpj
vN6Xb3Enxg+QIgat5P2KlurJ91cp8rxZb3k2TIcmszGtnDnPaIgRnWl/kjzw4r6Uz+qAVyH9uYjH
UwNZJhpOwCu4BUgPmaYm4xrmfgMeZOBj/Loc7Z19x+0jSOTHSlpVVSQ35mVW7YgOcOIunG7AGdt0
EO0+TMaPS0fxfwESL9q43HmABy1csGx/euXZLTPShQd6vmPiNEVk5FG3TJj1QlsYJ/XvkujX3ST1
e33kCrVeGv7sT+U0N5f7R81zVDeZpCH/AAF6QKKEGncIMcYQ8T9FwzrVLjBWoPSu3KWPAgFwMjKv
I3CE0sRYoIBkPqK9yhOEhnQ8iySwKA/spmy2z+NOAGAU9HUPhMIMAu9lPXjVGb1sfg+7FXHE3xOp
6r7U8K2rSSwJegIBJqtNDWv0ZWPWQaa/85tNfA4s8XlWQ6TUwb2xw+lRrBufyxugC4NACTfDeBez
eyletZA6/Xfc7/kV9IUSQplvF029A3oLAe38VQlzQnZq1H/LM5He0XzgIRd7A12HUmiI7c+uIV3O
o89rbnkbLUu0emgoLa/OPGGahIyzOaHJZI58o//tUGFQmEzg4TiaEeYB9SO6aPQBWkmfkbZuz0U3
d2tObLdbmK2W+2b7+zGUvQp/Y2Mp1j3NiQS93fZ5aEC3/VlPUwmEJSUKBi+nArpLzEJerMOeNkXs
3DTqmcgWi1Fw4G9NpnxJ/2AmPZNwLXOZt7vxpmiEeGDcs4+WjSc8KcqnmAaqB85ayOmbImv+961u
KUB+g2oGu3js0DzTfK7b7ZkA9Tf6Q3eAyOG0Xqk7jYSaa2m/eEJhpdA5W4Je6DPVo51QPr3B4pVw
cYseIIIHKXAoNwFpYqBGdUe0U9ypDHPTceVIk/ImTJVLZ6qcUE4jckcMLpVSOoHsHP9LyNGC5mgy
RcEHwqfGiCYP6AaBDGPD1fARTtBKydPD0kww5lazgefIbA6L31mT/wTqq7Yg0VU5CwDJjaWltu0G
DMGecgSWvi1Nd757m/YikrrV0HGoPdHWeGlQC5LwBg5dcDvG8o2CJ0T/tgEyFZWtPkLqLFzyKdyr
pH48eaHG3FrS/HR2PKb+Mhoad2a23B/dZuhAJAl+Tm+nO63CEmwhBddeslw+LvVSbagWoa1ADTiG
+Xx5dSaQK+DVW7AsjXKCmw6aonCX6f3CRD9e/mQ9KQlcWege70xMvmuFtNkTZSJ8YvLHswfrOEeq
Z77Lyh6BKHJTAIfhfENzty8bp8PXWiF+fDOqAbTJlqlIapQD3YILdf7uz3IDX3d3RZL9xU37b0BH
lG9Kf0EPQ9AEzWpm+7JOsrsFASxyo2CpDHZy49ldPVvvEH/NNPNLvGEiwCH2IkxniT3mOfNzQh7H
zxxZ3yDonq08WkQJAhh59jrdGMBOsPnQguu9b2tMKIx2EoE1TxEUh+FiyZbrFVVBZRRvLaKdbiFf
YGg7tDZTBMqqYb/iZ3dxIR3ZHZRVP/BVACbjY+7rM1rfLJWBskMaaiY+WLYBy04GBrimXHTXsH8t
mazVYT+ZkILTvVUejAy4fRNrkHOpWYyuMjHgvsikud16sB1ZMkPh43jMBlCWr4BBiCqCe8r0+xH9
NlGQaS4K0Dq6JmEsmZa/WHkyWt+an/FiEUCPRhZTe8YCvrxBoXuE+aMIS4vQoHJ7vYwKohXVRtWJ
lBUdbzKB6gklXZ5g8Kwe0mItw6N0KllGdsYLm/wC0MP/++B9wOTUUDYBcIS2mA0hfGNrvISKNate
zIBnGuYQuTXMzjLk1NiRxr2C/wSE+kqJhAEWY6Gln1mcxZyucW0bYNyJw++R7PSqjKb64NgzhkJI
74V89G2S+hPJHrUdmWGE0urxqpcW9m+CFeAar6CrHEo0CshEYAJB+dz15cYgmcurAYWGamVuKVZb
nZBvjWN4pTflzu3fNJ+rxu7P9QTDHGG3Yp9ybumNgo5KZkPcmHvg89Kv27NEMv8jUlLyPRnM1m2I
27htIeh6SQaLpApcNfrSv4B7scR+U75bzLAjFpTsMV3HDooSC2THbp4c9n/iiDi1cSa/T7CPhSvV
a88YQWC9Py6ydE2+gN/FGyY32dVHcsSV4wWF3TfDB2P+n4X7ZJEWOboVeUYNJazCoY0iLft/QuKq
2SIXxLfdF77iRyf3R3qRB/MqP2eyC0JCe9u2qdOqoCorrP5cgFvRCOF8PfmPvGnYgApvYSXYyQmK
FL2NgUxeNKenTL25opExmCtxn/C3rTJg9oTyLbYM9aodrplYfQZ06HTkUxlQzpDcUeB0cXZDgZpP
htleT68MYO5IvixwcfBqJq8UQJCD5XX3sx6un2DsXH+xRnOTrbrbKGsT3RjSI1Q+bYtsE7KZ2CUE
KuBCEPqiaBNSPco9pC816+9CqtyKBcRI8nSAakR2elCajMZE/L5u4qTYac04WR/A38IO8KShm30u
6GVSREGqqfYyQ+z/SywkMyqzfLDkVqoIqwT+BSleb5Y6Cyb69i0QdGC+7/Xvidr7IR4/ypQJJ68n
zBJLk+/5TB947b8g/EetC8U59kX0s9n4qEFNta2J2EJ00gYhxK+NX6iAxgHUkXf1fSN1W9DfYqt+
ea92ULUZjcjG1IuAVWcjN8uT6Tt4gtl4Iqg2eyTwvcOeic3fj6Pv+90KucoD1vMmKTqTxXDZaq75
3TQaUFBeRhOiQxL4wlIKEGHQuqm2aEUQ3zemtm8aVhhTy92m8vdaMDCpbWrfc6dPbRsT9y8q1BwQ
PTqocfE4m37myL9TG4Cq3dUk/yztj7lzjH80FxUCid143AipiEuytnFqDLnYaU8bNMiMA2Allu4m
nuC0yf0tv70aJXypQUXOgHRc1qeBARk1bW95uAc5LumI80vaqDOpb3NAz5QPEIJhTBA9hIzEpYzG
P+z/Tny3PQ87cD0uvdac+/AMrXSp6vjBPtrfRPmvsZiL7LTGerRFRDv+8OJj0n8U/9VAPFSohlis
Z9IGL/mTn4YGxYXUN3k0CDzo51WoncC7Ap2t1eVg0EcBxBlyEDatK6nWtDtKgF7nRVYExtNyhefX
WhXmKVbU7KIri6ppbx4mytigBel+o/+0GaKHKfvl/mzf8Oy5Ljyu6CyysFWs1iZZfp9Wb1/DuMTK
U41dtkwNPRLOvhN+u9msWxCs/swNcLPkwtYeRtnc/QJFqfB+31njBqds1dUnAYMgx2o5ZWN3tTpg
pdzAlHuSJg6AdXHkgQ5rgYOUkndgscNIlBCZ91F0WupiAiwzQ32bKq3mGItm3Jzrj+T4qr+vdJ4+
i0ECQ0QvVRR52B8q9Tyij6vGIsI4USJ0EK4SSE7UQCiZvandt6k6luddF3oRsYZPyu6sEksAkzBP
D7PqIb5E+i5/xDfq5p9hXGb0P5R4cBa4p4YVorNG/fWlxzEo16A+eX93vTIuG/B/l/CuGyC22vvb
aUO0V1ZOtUuVrXxy2rz8alNcl13Lh2pSPl31vaZbD9vwOW3Q5YGTx/52WChwqG/Jtpgj3UzcIf+U
KA8Kfg8uK6UHg7CnPG3VvLFrcLE0ugVG8ZZ5aS+NoOks8dnr/oZA/XLFTMZ46zZVosyLrSgUNZ0D
sIA1+4QQmLYezznriygSQ4WmXdbezjJg3OvC6LtLlIz5zkdDRrPnlYZ7wlsVooy9idq2kxk67tgh
MBLGwgvh3b5HB1f/9jW0tXoltAQ3dBQhPyjiBVGC3//rqLCMUuxtAgrIroliNaB5DhzijW3V9fDI
qUszpkE0rIYLWHgxCd9Pm/lcrTF3z83MgCLem/oNMMeOg50jKc/nrEKM948jHzJrkzopW1HTiXsn
de0hvZsF5P7pL8T6PBvjX99kiNZydwGIENNrGAcvob+/+Hk3fpCKGi9hMGSzAuXORdLiOBFo4W8a
p0Tjqeuf7hDVy5jehZnDw8reHs0udSOKyE0w61oLIEDNLSu/t13DVZWfYBeGhZ9QpYym2h4pmGES
ti5dg4BjjhBgdtC8IC89ATvEFjcXEafggJib24Zn8yNrBjpW3B3hcYEeBuGwk5stFLbZmxRKBF2P
QdHKJa78E4wxiBevHn2Gc9q/k5yM+CN5DMbrJ/mIINIhpfhH8kBFu42jovQXaUKX83+Rf1wFCdSq
tv+iLAAsjAn3E/srDMfCa/U6LkbOTq4yZLKU1en+QtgCHflAhcZyfyr+y6cqdKgE7T+iEW4gpiAS
FECerxdz3N6oF7MRP0FwrQwfDuZZPZ5lAjAmfk5HogETN5f7XVNi6QSrNjO9jMgvJJhflETXDSMQ
7odBN5nq++MY763ppb4VUXojRaeLQaLDUsuDLwR0oYnGd+ddBKNwx+mvfI86avFAseLfIRtU2WjQ
o4ALNVqJnE+aVl1CshxcLhYxM5eoca5HYGrx9kTJVA2FaN45fYpEZIqu1RJgGZfy4zIyrZiiZLV3
al2nqUH5C0dqWOxIXdp4/78XegO2EkiunKsRHhQpFZpwzXuWjNYe4VbrSnWOWq3uvB0OSPqm7L+q
YiydJVilFoMxSfWbmSY68ZMDLIKtzO6K08EVFteE1UlCSu+J3fZLMxiwpjKroLB2LOE8s0QgKOgM
QPyqJBYDlu4dVhw96svd52mlthjajbCjsllR4mduy6T6SezwDB09QA1OYcKI7/ELGID3oaaWZlIy
wJhgOWkNqjEfWXfr10wZK8S3NSt/OHqTUcXvjSTEZ9f/3B0pfyut20m8eD79AKeqhG7SLCWE06uf
W3arPgPFd1FjRsYku80/Q3xq5kHc1Q5ZQpHVx2PT8pWtjy2RE6MLRjQo/cPFFGOCxxEIdj8cElhU
yzKKe3YhGDI8RFBpEPc8k79ETZ2uWlN3RfvpgdlGiDy2u62Q1KIAXrRbOLaWc9aAqNOHNdUGMC5+
O2Au4tWRdASAJAMs18xM3ajJJ4YcFk/SxeSADk4XlTMNjdwJrhJne0U8uIiA+3Ea7N9iLWCNz+gB
mH6mgKR1QAdI2DdsBC2mFnbL715PAuyIDguSxpkA1so7nnleIL4Z6dCRwlrTh/yYWr6rVGPiVthM
aYZ3Vx3FWBxlKKjFMRivYClQq2emQ+wm6GuO9UtvcasFasShLCfS2WjaEJqgl4ArJp+IIs/BoG2O
OCQyDKf6AiWqM25NRA8JTFyHA52U4V0GIfwf5xeY08zQdNVfjSKFmALI9i8mZHIVAKXIPaegbLda
f6nk9+cAKytF/dKm/0oUNwRmG2LwLtzV97J6Y3COkRCResdIbQmdhlRw4JKbBrONpknE2iWK6JAf
zjLbSZk6S1gHrlYdN+L79brtkX2R6UBJHs7PyljhtBDJSGlGjwsBGgEnUQjcswHUfod3mw1BZXE7
xJLPzOiW0cb0wi+nN6trU/HoqwccHYYM1U10c/w9YkIxadvycbp3mIgpWTllqiaLvxyjTZkgwh0b
bZOdnH/hEfZtMnqSlbtDY6At5oNaK8cih9wxFZ8mHRcy/eONDB+1Ne6g1ylK9HTi0VNjCSiG2Vbr
GxMipa/QRwSvT+kmf9yaHKXshQOGRuNzujbUQhysVXQujqUqrQezDz8DokeKE/J1C5g9ZMQNJeLa
HcUFDxVvlInnhsQ7JzjRE/tfXiaXkS3EvF/kiK9J94T8h8iQAUHSKO9G35qKCZwDG+GU5jEQEGVJ
cT7xpRftLeq4wUiv4tYOZQAcvZ8TUU+lE+Gw0aNHVBb+pR83wMyDj8ckgGCBczyI+YMIAwL0Wgl4
veYcr1wjXWfZ1e80vvVtpDKOhM0iW4POvzjUrzE2gATid0d6EqlsQ6rVn1FI7PsXy1bBktsNuPxY
QrfX7eHzagl4xCyQn+zqjYK+OfyAxKazaZe1F1nQ7ASyvOIoxpXveS2pKHNWXsRZoHYnybQlJK0U
zAU9wQPpItBq9sUn8DE1dYB7vHQmP8JVowho/gJS+FLZ+/0buP8DbkRL4D42HfQYjRaQy7BAQiiO
iX8cgmBEY7Q5tqIhJ3ZrgF/FyAh2/Vg6Qm6PuZbMHzNWsDcgtWmjzxmo/MxIzOXHs7hzAjtqATqS
Er6tkYA2UQZjMwWzO6BBO24OLDwvYrmKhzREBwpxcOvzMPLe+84sCiOAyScu7AjbDUUrTnsynPHb
9MFiRy0QK8OV1cOnCTyv9SCDLWB0a6uqYTjfTEB10Sq2Z0AAKSTSK2rx8CpV1BW8RVAb5XqBW2Rn
sHlblPX3U4dGTLWLoNUd8t+Rr1WWq9IcbmRfZN14aBSPvmXNj3GlO1NkgbpnR3ayT4VBZI/7BuBX
9pD38PS92dpi9pXVMD4UNA75xApGj/jINkqPT6Otz2SzIRpXI8I03TGMZZtLSuFf6JEIE1PdzaVy
OQVEWIGZDc+i2K723hluK75H36ZXaBf8sNLJ2ivDSAXg/alK0LBHoRtDw5cHU0/YeAZf9MJlVldV
NXYflMPNLcGQ4Pj+hOrScysXjzHcbn7aVm9AKzfDemS/yk67s4ImfPghVK/fAFp8qtax453jRpGv
8Qjl8z2c8+U7aMyBuTo2mPwQbI5iCFiideELFZYLhGN9A/jTXvOyNLvaZP0jf2EMYwWbnfQtePkx
X766e1XdkM+NehyTzG6+euanSMjLuAKL5N1kNY0gp1eJMGs3NB3f3MQO0AStTQOB9UPG6Qi79fS/
PV/JSmDy5JnYWoVbjtYe2eX1b0eLS9rGE3TB/eMUjF8shKk/NWlaGLIf+nyavOARQgNxSekScf0v
ueV22ApG4Izx34yXlvLgAwbGhFKTYveGHL7EcrXMIdvUK4lAVPuD1SP3WUPCjbwFCFFQjkYHLZi0
0nDDOC/52zManR2X/Qfyso3tPp9L7RypGW5Nz/QtOH6zZL+SeHl+XHteBTsHoEzIaZvwFCjiJuOj
ZdDu0U4ED0rm92oMzffAizDqqQSsXuQT2x8BUFKUp/iCxma8Rh6ztiWBu3gsvfD20Xffn9plPu66
LhvkagHp6XmEEs57YHCEaqHpxNkPgcMYDQXoOtMNk1oRmqXroJNCHCPmDU4hyOfG3QKXLanhjlql
ZEsuApPvEQiM7/lfZUMlyDDgovFHrkkZEhR7byMuJDk3wpw4TsO5xxv0sakwWmROFbDIggtuFhXU
z3wmh9Gxs4bqEnMF8sHgFVIxm4EZv2q/zVrYmtkdOMvUDyeHwvsX1ve4M7CBVhgo8Q1hhZo4OHgs
HnYtAcxf949sy/6kwIucsn2oA2CzAsdoDLPlCnp44mCq97aNx2KSNFCE4N4qo8quLQUDEORHsscU
KDVQNUVIPNyhNso6+e+EuxvO32OC82JMxtmIVmiqDtWxmAPqHkob3tE6Tb/bSo53WC5IBqLaxku4
A3ArI5g8rTxkf0XLiauO7G5sOdVrCFjz4DknJ+QqxjA3o03Mv9vXL9IT5tsQ9jdr89pWCHG5li9S
b/3F307+e8Ztly12r05VxE2+ovcVgmvWwJ4ztho/v7E6ISwNziQdJPewwsfrTxScxxA/6LiGupzO
MZGCbvq1Sl+SPpm2Tr8gIEfqazGhMKEQ4/yo1w7H8WYGIFlYKpFZNOCCXego1BNBR3siBHYKyjjq
jTJXIbOApSK8YddTa4ldrNsfSu9aFYR/KRuDgn9sL8HYkSI1j98YHd075ux4eGz9AHHKywcvY5Ak
1+aPwwQ2Eia8w0WvaPjWG1JA6BeMtzzzqD4x73knhhc10iLIuGsH9VrtY7AWDPx15MolLQEHTHRY
mexUNE1mEprof3nDNyC5ObztlHqLPiS6nRkFJEawM0CWiy6HAjotxERkRu/Wxo9Aw5KA4Svjy13L
++6aF2DcW7oW9rSNRPFVI0uZ6GtDj3Yo5351cq0jtXHY6ijvQfRVelCsvhAbP3Kux/LgpcXlfYeJ
XurZp4ZaaPMVvdtpnc4/b00fzYYcx3TORbCGWt38HbjnU5wY7fiFA0fu0NPROqnj7prpPjRxtIM9
t/XNGNu6KRff/wgwhshwS1kAaHur5oHKzUx53FD5nQ1TcjsBjWMROGqT0Em1hCkrMQC8eVwZLxhy
ze7CZwRA4wlCN9fLQj5j+rwjg8KfUPetudtiEzznNRMPdr5dl9VSutA8OV2/R9vAuk51+4xJapOJ
fi0oBXZ6f8iARw7C/pnqn1azrkkvbSE+LVyKQVJ9JPxMAwR0206i0CZx57E35Bu1+OJz0FHpH2IO
71SL3X9NpyKyZ0pvzVkg8qaFeXHnIz+qgOlbBoHTVRzbE6CQos9EU5P1AHP9DpZcA8KuAb5tRgRV
yf1/sfpfc0cOESKGffna/QFxdijT8/lc/1TYedaW0Cs2FAymLkUwtPiA8zVKPTkg2jgt06bdt1ka
KtS2C0P+vj+8xbLfC++DSQ1JW5bLhxFS/JII9qUCcSNvwMk0Ja1icmeex7PJ2d77ZW0IHmQLdM3d
fOkZidOFTTDswK/BaZkptPImFPMIj2+NOzQRcwevlOMlHBWoIbm2pvcY8Q1ntMNSZwpRqz/8Y/PP
EIzvk/q7DH+49tgqpsF35TLHN5t+wvJfkOiCeJ9QJh0vVOY+VdKBIfY30YC7KvJxnznHuKuRNKGN
ljxes6ijP0r41x81uAQ43LUG4dLcJYGxPLj6xt1J/Aoh5D01n4/yRg3NDIduP5B7WNYJMDLFVCkN
wQtdBAmmpS7R1ViogZnF+g9KUtLF/3kACw0YzaonJOJ8VZhbeJfDH9P4BmTzuqCJ54rq5oUFkgBI
CcO5h3nn4M9+boKlbWbUzwU07OpofsnTksNohleeapaL/Fca9ZcNQxbz6Ix7j71M47zifzaaPrGU
qkvIa/JP2q7RgfDE7DP8cO4BeRv9cp56PcdfYvXaY0lbjuLKCDwjS0N3+k8AoFIVHM9Fkp8EOzT2
96eu0fklVODBZdl3kiTVRxH6dSHos+h9Or4j4XBcVRODQCsFs4uT9mD0T9mSJw0Ifqk3xAkS7zOz
m4rfSAbI6IvdoJUY8SFdbdlfAUcNZQZsaJbFeMbHjAqtVmgsa7t1TjX9u2OC0HhsQtI2UXZZlXui
UgMUqYbE/QmQjH7WSQzC4QIgnrU0Boo2/Iyv4Z0RRWugOOWWQds1ymOajzWZpn2XK6SH0sVcSZWU
58P+6wc2ajqLRDuickwAjOYASQMUpvUM77LwDOw+JF87Td4ACjpHavaNQNGSAZf4u3BkSxaIJeFQ
+AaDM0NpTL/6RUtRHKj4FV1V+vtS+PHOuxbtYKvMeriRvR5uk95k1iA+vcQHWjjSvBdjGwOCTBAI
cJy3XPPSvXu4+jzawIkHiz6FcTWizop+7F7Je0aKAUVbPIP/dvnTJn7FHoRaeHfK1MSRyFx0TXh8
7U745EqXBjg4iQBu2wPH+VU2U5oRS2QjGN0FuXYt2Id/+59lg2XggHeANObfqDRiZ9J97dyhJmDy
Db1EZu0HanGKDI1R3ZIJZ7AidJRUqn3xRXuO2lIH122lk+dQHB48RUAsOQjeo2s09/QZXues6GoD
7SNja00aG52YlU3SvQvFhRN06Tu1/I0tMTva1D3clr34l0ZN6BQQMXEzdahy7dtUpetiK8bXBBEQ
WAKQIWB400QPctWXRM8rI5RrZOixlXvqHfJR/nfyYIQmjVLj46ntWAMvzl4itIPVrhnVbHDNou8d
QIiCXjwJpyU3PHwQoeZ8N4X6lkn4g3TP1BJjHI7YhKfB/ffeXs5TOAun37BKQHDY2uJt9ECY+b0A
OxupGEyCQq1T/A17zO6BAqO5bVGGPvglHr17wn3VnjdzXbm1hYstoZMr5acM7EqoCJw5atbW15rl
Lw1dV8WUmTfN2yJ8IxHWfGkgEro+E0DgzL8bU+VbNpipBsiU+1SibB9BUkizMiFHML+CLI48Fv2y
wONFlgCYZ+mAH5OJT49qj4qE70WLZaFIrYLk69dGZKElniKsGaNotqEKSAfWqiap07yykIgRhVIx
no6WVSxS53N0uturIvXK9gfbvYvvDrsWjzFbFWmT2F6CcuKwxOzqFwpy5f4WA+520vxZsmxdtwfr
qOX7l4b293Vlg1oIbKmKgIzRVavbKXPam8JEdHWFkVlWR0668PApiQ7Q97VguuKdbmWO8tZaSjqv
OU+bum6D5wVaLjz8GRQOBPEAzwNybFXdOcSr/ooR6+E+XFP8ndlkmoPuylTUav5zUzXrqqi+O7Dp
4uE7phI20fNYoabE3BBo6GL/2KWeoYCDPAfboYDOkg8krowk1gWtWJdfLL7BdHAw0N+g0rPhBEQQ
rRIujFMZmMMTo655BEz31PIDw38GxIbdT3wkv3gNzNzoi5D1MLGQPjZbGBLhQV18xRA/ljr5X8RK
YeRt/VZJHXcsta6dJEc1/1e3P/FgHHYECLzE/3Mxnr4unJN9DrHHRIX4XFUKOkZJA7yCkNX5o18A
jNbP1lYVgBPMChEgDd1gDnHQxy9qHTpTKfJ/6GVl6VE89TpgN22jtzSz22YojWHT4fJQbDwiGedn
6gbVM8tIEsZvQMsOVfQdSB3eO6JkmiCglXqkH3buMi1Sh750LPjmaizdig5Wqds5RSm+2lHbYTB4
crAUJZ3K38B43Mxm/OhLHtAZMRBftne8TacF+uQKvl71a0mCqZiTeJgzhDFXysWudZ3iL/3VnuEe
itzqYHtJO/QyrxOTbdk1wQra2+o4WLw2HgPyuTvpjU2L+ppnKcD51gmpYxeCncDpwki2KS9/E6ST
s7Z56Ava4JQPu91WPrFq422J3daNGl7qDchKMBu9VvfRbX/Dy2CNOVRCrI4IM2B/2Gc/iNOqb8Pk
CkjHGcHqC3FLMeKQNg/HQG/XRayRAn+PfLlJSfR1e/HnvapsiwKOfRHPpWR8kcIrbPzvdREdLw+n
ffD5sbBfikjPz2Sgc+PsHtD1nopKB4OZCZj9FlQqIKff+gB9Iu42qMU7rb0KikfuSoBfyLjpQ8t4
PYZKR/K6dWimAQafhL2Yka9tJ6rBuLat9X/VtVyeoEpjNwxp68dxyDyPWwureU0AUXuG4yMIzL8r
zuW6dwFwEySafh19ym6OdlsxuafYbsxYGLOVEMYUwLO4lCRMKBJoyawVW/97uEBefWx/FrYzh0/j
O4lv6Kba7RNbjJ8zU96WGzkkBZZPF0bP/ajqbXFUQ1p+4XK4KLdF7pr85bhSf8Sqjl4TgMilySmQ
ylIbqqmnVjYDTbcTqT0JWC0KuZtpnuLjnk6EpnF6uUq9aj7+/2RHYVEXW7Vr89lMZg3xL6v3Axxw
QECEz+EH6UqsztQQRfzcWoo1v3LaWvUhjH7SN8KnltBUHqsJ7C74ozUmPL1dfWl7l9HSlDpSzRej
cbQXk6AXR5YkiQo1r+2r0G7JZXC4yo+9i9NAtAuhTIkqrzAYG3dnqdRY8K4CPH65PjL0wuVl9Qfa
YhwtiT8rarzDwwFBcUZrXgfu7KNGbfDFXPVMlUMTe5R72ypcW0tAQcYNeeuLlByC68TMT0rntnjG
I/Yob9vlZHNdUK2XtEdsT0snUryibp9ijl6tWjRGf9eZsfZT8CaPj6dsc4vm6tj4UoviXordIpif
2apYm1ho05ghyCyFRRSml6arW1w46khZ4PTPv55W7/AYbP6edlyZyn0IadiFvu3Gncq12lVN4Rdo
wgxn5iI6dcoHvB7UkOUmzWu2hr/OmLal9eiJNC1YrT6n6fSN/p5iD8iVhjv3ZNFKaCaY8T5wXi/m
FTUcHRpHVcXNpjXC/kl56cRwNcR5Uee/5/c/BDbosYR8ksxN3ZIDyZp7uF+l0y5YB6piMA9MoH5M
kBgtnoTabVbSpA9cIDkONIHcUCyG12Ay6e28QBAhqm9E+UJnwiQAtKyrKkwIViCaS61h+/4pAvsQ
WEYLnDa4t46SmZASwkKhyfB740eWMdXXtagSBrxYw0k7I8AOqKC+ITpxjn3TPVyzdOS9ywojErHa
Vntf88z6SnWB+iOb4S6Uo4xaD7GjmB/o0x7Gif9zOcWdh48zbt2TYnB+P6SMdhVbLJhkDmX5NhE0
Vr+uZ3ynNTO8tGbWrZn49zCOpFW1ST9Pnp9UJ09keM48LH6OCgPVhAKNC3H6AzrEC7rkhk0RoDxq
wr7w96vwhVKlv1QttlIB5UAEIJ5IiEHSWUYPjUP8qVTg5ORrwPric8DtDCvrnSNu4Mo/9ExmwrLB
dSuz/qXDMJFxLRxSYTjvMqn7IVviP3HURwUZ24HaWIPQNSvfn+yCyml/Ax4M9FFrERwWr+qlYSuW
jLBCCz5G5XKijfdJd05jFM7WMD6rzeoBBKNhG6ZMwNMBuVBwN3TKu0StUhY7CQqO5xePhfYvf8U1
vi2fxyb2BfQpUIQFIHArGqcl2hrqxVF+lshMTq7oBrm9FBHKqIkg7xKx93y+4cwa7Y2Mhwh3h1R1
5R+gcGoKC4w0+YbA/sZ8n5dbMaPkwulGK0Q72ZjAY0ubENc9bZJJ4ZkS6mZlbG4ye7/6xT/V/ng6
/n37BobBVQFuEfcXwZhTx5njdbMBPN10bx4UlV7V9xVJlwTUPffK98M79WDmfyPhKjACR0E5huJ3
xl+cvPK1jLfyIDUFV5M7DSoqm21hFN6kKIKAisM/WKhfKQKx3LKVFY0K5KEjvLnevmlBS6ZMthZK
pF3mNeWYcw2jXAzsirNpPrzyc00FJeUrYju0OcxXUPnZ/pn2iWuMTt0dR6EtB1vfUl6OGd+HMzs/
X+/DvKQkN2ii9FzxNV4a5qX+zSC4T/goU9z0k8yPS67UCeqAzb6ep3GJtxNQdQT8bC38HOkRr5v0
8a1vThEuAdHkcX3otOij5ehixefzQTDDoZQX2FeR6Jy43gYWwkKacuTQubDpv7qbW5N1XhK4Zrqb
mMgLwuTt9OD492yEGwwOQhGzDKmxOMzNpvZq5xvBxq6XZ+Ijv7AputK6Beq7bDWhs1MkW3V6gzYW
ZtaIM/ZLY8lva8d5uJ5DMmsQV6LKi2L+JmuGaGpBQ2f5eu5fG9MHm9QPw4yK2bPo8z++zuM/ynPj
la3PwDKAtIcVLKNfAmCU4Glt2IEZdrb2ozCQsoI6h+jFtIp0FEhRwbZd4wWhOXBFKJShoD8yZZ3Z
VRazDM1R7rRMoGO1QkUDh5Yn5k7vzTSOdm5D9OuiuL2QVni6isRPduS3gmVYD+rIKVibv+4kNyrF
Kyj7npUbRtiVDhgimrDnPPnspg9cms2z3UCuxCzuzKz7hJMmDZq9Xp0JI/+jHH/BO0nIwBvaX3wN
vf0a0IEnpdu23+A6c+py3+DYjk7O9LmwHVMFMZLyDYlD2BLYTEdvEeWWJZsl3xcPR0jhqR5seHCW
k8PkI6DtBoHDCkf5udC0kzrapTfhaJTQNy5Pmn8gGAm2XsR7p3TL06BzrlX1Fyj48rwX+dPOj7NR
1ElfqWkiV7AFb6c8Ig+P/F40xeGSDI3v1UdHYI4fRbVP9ub2/7R1XE3zaB9Idp2hYXqmQsGLlmzD
9lKlttfB6p/8cH9W3iXytqWA/FMcM0Ev1hXzpx82Dj3CVN5qe3HnbXv3CY2vD8Brj8u0bt8YzIND
kMBitPwbeDZaRudDUfdYrv23OgagCdj6IuGt/fvCr/eol8eFxQFrl2y/aAurQbyMi/PWzwjKzP4l
T7oSA0MvU6McgUyY9G49ENrgWKEgrUnig6PPT1AaPfbdGd/DHHtGE6SIavchzHQ+oMaRqivYSA43
LJlJa8WRUJ0M8N4+x9egK3sCe2JU2UjpEU7tx9ZyItsEd+810UgmtiB/Ok+XDTSaxg+TyDc4mWHd
BV+8yHD40QwveukVIf8Wjr5scYDhvBcXcAriFTRO/v+rYXqu5ghqg0YniipiQR7XbTzfy2aOraVR
9BoHfaIArOMlJZl82BvN5sghkMpduYuWLzEZ7+daoy5eLZeXkLIuKJOhR9HYCkKiyOGyDG2EhUEl
CmxzqNCfZc/9FXG0MshKNqHadFvBLl0Ymv0oPRRPQzq0c22rM1qPJ7kIjQzmQsWaLxxRvqVj0yKn
LKXBSEBqlKjOcRvhCtN1qoouFX2FOazvY6+e6ouluds3gN4s9nduiVZKrUmOs95r6Mi4BrlIuMXI
1/4bf/1tfNPx61FQbwEmkcS2wEZ/rnUPX1IXr7bafGZHKYjGujnudENdxxnIHGUMAj/qzNpUe5n/
HynuQyV7bAUD+rYCLQm6a/R1CmonYI+NCMQDLTFql1ysxaIaLOqF1p4+Ej13AhCwJttGinG0NUJ7
10tSvIg/3nP3wbB3bLHiyG2JOUFJVgTyclIq5OnM/RB/m06eeY7eEBvm4e0Y+BS+r2AZw4P32Lvp
MJ/74/eOzGCOEjSrwT4LrfzG/m/tEObtzHBrwmksvzPxnOd4M1HuFQ8c1FUneNAVl3G8A1z4Wk9A
Kj4aX3AVhd1+AsX+1LPP+IcFFhOynSNFvKi3MTSAvkj4jLuQRVtEZCpOjBUDTfAHBS7jLEf8dosw
r9sHPybt3C36LsZ7a++c3/HoT8MzTlsl5c3BauhZAVl8h5UhrcLug7iXf60m4QWqvzxFeHsj4amf
ny0gn0Ka3Op2UJLVWM2vh1+eudYQ5NXqHsgkDAzovfAWcZeeMa2M5t0RcEJH9WrVFT64DdDEHAQP
vrfQaN1TEzOJQReiwH13fSrpNyYiNfy+rTpcmruTwGWIxIo6lO1Ki5hxjVHByiaKH7e0XOSkhZ5q
2yD4UxcvTGmckpdjsybmtxuWrNcH5beBh+D6XBucvnwLqx/befs3BVOmKnGr8zYhvzJx7oebPyvG
CE9YpWsppIhMdaqsTs5cwDiXQOq2I1SEucb9Y/GBbMgTpoWPLJbF58X4UUvypIE/l1ROK27r1RKh
GxCcGpv9DB+9k35/2LywHElhBDzYG0PDI4mo8aPolZ8VnbJbsmtKb67TjYtG/ywLr9XYQWP9u3y1
AvloqGtikvR6/FKEf5XTbfXE/DDMzm8tez2mgekxTizAi3+BpIJj5YMAZT6v5KHIbQM0UsSQ3T9R
Ub/IUjYx3LbpDMWaRYMakF6bF8r86JDy7hY1MY/SjROtr917sw21mpi19oTAF9elE+Ead/0J2H45
KAej4ngxYaUUjkm37QgETL0rqAtOYoET10ZXcpyi4pwVSUhWH6PIBpQMC5glvzcDBGBSqGmSb5kp
Zmj8Sn2DCaGBDPCA/B5w14Qc+ERUHXMCVfPxYmpQCAVI8eN0UkeePDmCbNk1dme5ymtyGknZiItE
e3EtSbEMZu/pY5Y3+3cnTMKJUqc/6zVkCL7oCj/pUWPqt2U3GnIFa+89x+f7MGmxFXLP0+SAfxCX
MJ1nKPZq2XZqa2wMfjjhSPha1aADAuVz2OpjhQCjC80fH5j39B9GUE45Bv76d176sHt3oEHnBpuP
iNegWAAhXonHNpulfwxywC+cOGdbrznz2Qm3SeuZHbkAyYjtsWZ6VvxiGSyb0Tc3VWle6NPc9yDR
LOkSUsuJVcA9LW/KpNUO2spF7AmS5ogDzDb7TH9CDDQmfsJ+udXMekgEw4RM2fJwj3ALMaOYkTD1
bqIdRcaqZktGBr9v2bN87oLMFspKULpO6knCrC7MmO0W8urfs8ZKKZ0EFbJzSGmbswSrB6qZorP7
E73mX+8en7bLvFXC5e2k8b+udNg+fMPL4Zp23hR8zzJW+lUrgEYM6TRAHkapzLKtYcMElgiUKtH5
zTxCworpVHd/s3GQMfqZONKt0CACNpluALwCj+ZpT+CncB/VJl/LVqvvoHmMsqUbaTu97lAV5Sic
0jWHHk7JTmu+ppV+0NPfJpK86SQMKHMLmSQbLYSI0LPdPCCrywGzXx+FFWoF3n1xSb1tAWa8HpJH
KT/tg+1Me3+u2+v7HtVELqdaeS2xYuLibLaFBuv7KYpMgv9UA+8ToprE/z+JS92pFQU6XEWY0MCb
0Y4N+ewNSRLiLhREWBGNAqKbEPT2+r8D6ZhP/mqeJCrY96jJXySj+Jin5jhqjyvHZNsBSuNRvpXu
Qu7ud4xU6QMPRSysGasSU+cZVBKk+Orva3mwPJ1JReALEpY7JTEwdfxYnyVptqpGDYQOwJ1vCYYU
kM6Bm4tV0tY9PsV2xwUPjXUOJ2LCg/XwoiXeo18yTCyRFQ8rIx7TXZefAlRiqhMZSnbNUa2OLo9K
Agb2CTQ2UrScQcCNSLYVofVSKYF2kzezpEo+Hpap3caVaVSgnTt7fQh3PYQNXX4E5/v+AnFVTb3e
LmNj758HOLCgvSVPXJ6pfRa9dvBJkDXEVaPyG5M74rr51PYKUlC+uCmY4fS2DAoHCLI9gJJNN82K
QQ2GYAMu+Qk7spSjJ74Qkfq3H5z1KxfNhW682GCC9Vt0gkTxKICwUOlX0Hk66z3KIv2WbkQRTmYw
eib8Y1x6iUd6DWbAhh2pMALz/jlEmTdIo+TjAga8JF2nvjLeNPyp9sw3ml77qy2VAulgb9eHR4Ip
lENB5RY0Hn+f62Uu764D0lOVxI84DMZPe/FmuC8Yx1Vw72PmVuQhQx64se20NvnPXkmwbzZ1tcsD
wA/+si+SU8do+awwo2C5LQfA43uas0L9DlyyAe9pFTNXpFusLqsaRfdY6RwrGaVJgFJN5nrUsh1U
/dK6Vmn1TZb6/79Mxp8wupeJwPq6lKqaqqAJHETkZjGbkkAd+vLRXC7HOMi2vb9/Ric9jvrrmR4j
AtZz0vZpd2UBK52KF9q4KUJ2RuDOsskDeXO+VjkC0mKes6cNvNPsfikG1lAOrqmhFeC717B5Ak7B
3XwQ2xJ9o2YV4fsveHuzZZydeMSwbynrAb43BFV0CpmvXNYthJty2BEnOZ7kJoqWLZ8ZcVb27uqn
71yIBpYL4Y0b6Ck9MvNz8mqfB2DejhgffH/HR1XbyXob2jPeTBmSrXh1u2wR1DEZtb62TPUrYuT6
GgrSZVkzG5Lhh4ARcz+fD1A7qZC1IWZ7u8Uc/sqJpNx3GEj3qMdGi4wWn69j20ixXsqKPicOpZIv
FOmHeZWY9vTakK3ru3ytVl4D3s9TOdnEYPk4dvFwGaBWjmz0HXxOwacKDmLg4F+0NRps+h+xWnr3
8s46PhUtzU/LY79vwgblhMlATkdfFKZAeULNrbH0ImUZQ4heubmrEid+3oGFc8BIKMNAzsvBS0hj
lw5iQqm7gTT9eTY3rNkhpOEcOqEhin24kuaBQUFMo/wtnxX57vIuinPll8yrFbMkS8iDqCnNyMWK
A1sPTM1HfZz9fTxQe2ZS5q0KCkh5MrGn9xUy5el6GWC+snFbzlc65MgjdzF3bmzxumtd0W8cUmFE
1cznA0O2tNjIlbfG1g4DkYshn/k8T5cZmedrBn+PhDtcO5LoZmR6bR08bFaI/S9/fWAqm1rxgvqp
zL9VTXYvj1GFIfdPGk2Bv3eL/jVVvNJtI5vlYvv5AXJK7pbhHA1QeTbBnrI+tsUgLZ52wjzSA2bW
ObRRLO0Zo0OZhkyqGJo+XXATo0Y6kMllohG7j4XYQUwDBEJelLWkvlgtS0DWcq2qeXtY6ivuAxWh
xA8dsPxuth01k/io/zyRg/j+0PwAHTlfiVamx46DNoWkGoc8E1xjiSQQj5S0/JeXAy33fFwMpWDu
nApkmBXSEv6Va8RAEnAX7LioCjeyIYhao1nDINDXTCB3F0RW8yqIZHZawtlkHjS5moktwDfpbhHQ
M+e+MDl2OJeBBEevKhHAoB1BVwgvWnti0TMA3i+CLLA70hVzIdOt35B2gEd/IGoUeMaEwUnr0Gpn
SiVMd3c4iMQksAYMoS5bDf3iiBvIrBabSGllSDPHs8cvlmYfzOcZk5gq+B03uo7EJ2V4PuuwNgA7
HzeAcrAPosJ8sIir/fQzTftWxztSAGsTt/fq/ETAD5Qx5WMVa5xHgoeUMgq49HTOpLQWWFSKBXem
bf7LaHOnrT52AcS8XkB/cqKPANHnB2/FRkxd0BAyYmMb1OU7t/iJbKSDY2D5Ektgh0BsO+IY+FL0
HMUk3eHTbKknBG+tCZLF/b6yCtCxbt68v4/eqH0YTl1LU+K2//LNC2c1OiPdkRMZ1g/kgHs98YEw
36xnY6HrS5NMpcLJ6WSO6QIBuG98txytYXvZM6M1qMMgML6/WdsxZoBx2KYfYAOj2roTdB4tk9qf
4p2OS0ToN6uQV/tdctcH5bWgdyeM6Z4DytBOn02xce2c4Tu8NGckiOUW0lnEkQ7Gcc/jlNmKvuTs
S9IL0+SMP7j3nqcRSQCqjCLZBQaJeSiTX/c9igNlB8KvDGzH7Exlf28WeCeqeSoH1rckeQnmZdaI
No0h4z2T2ZdJyRFjYPYTjSmYU4u5JZuAaXdg85SfcLg46ogSVxO0GNJmJ4kEe0R34tcxqNsXnUYj
qgb+BQZ8Y+N/07JrNhcF97Q32DAAujU99EhH8Wr1EIymW9lOdQg/yLQO3WwMPNlXeYxF/H+X5PqN
8e6tbY7X+5APeto8LcuVHWHxVykul+XaFgfThdxQfE4/nN1ylUpKtYbVIsuH7/C/LGSXxRsc9NL2
37HkAr9r9R7uLMCp5XtqS6vRh+/d5T2HPqkewzuMLF3zFPRQRpmouHcS+EIhkQt9HaJ6ujlsB53d
I0z77heDUG7ZgFAWhJdurJCaSpz7JFGQnt1Ghmdiu//xsln8xokcD529vWNxVwK2bqMHMa6JBjE+
Wm6uYn/iFRAQK+k2agAPsMuk+erQpcVMDcCkZKru9VPAE0G/XYiQ2pa1CtBo9ir3GAN5FAj1M45W
x7aREB+V9oZgStEXorAGJqOzqyZ0/nVw1HoCPUF5Ia/62mM20lQ28eH5ZSrrNRqlObJGauLe7FvL
kny7FY7AFZlpOBOmRmF1TTrqoVmHWxCKDLn5SgJ2AKs5cyZgZa6U/ffEDlBDXrDRGQSrLxsz5msU
jf+79Zu8oXFT/9rT3NlMtJ3ifoLJw4jUp36etLJ3Dv18o0q6Nfdh0qc9V5nNQ1fPPS5o2g91u5xm
t52jutggOX8zvM7h5ulVgd4lARvg+2qfcJwpxs2iAoXNNwZdKl4vsWCBwk0ggFq7qcltEiMtJmNh
pNdH3sPaDS8TWlwqUrxeJDc5xXWyrK9H1oyW6yfU0Bv2Fx81Tz3nwis5XmKFe8iQ/I+bKLBbSQbR
CnmW004pf3P2l+P9FGVEg16J8qf+IBxhSAkyJ8g0G71jCFWmSSK3ZTp1CQ/ly7rr1tqXi4fuLQd6
5Mfa+B1kw2u/7FGcXYNAxIOMHOZkiXI7EYwqJuKiet3Y6BoQQIfY8b0ZYr5+gfJzGXt4t1yvTnGr
yWmr47NLANxSHI7SdbOHH4EnApuuE2tbPAMT1RTwbysihejquQ9RI58I+OEwQ1MaO8vLLV1BySlS
3HHOTjFkWtvEZPuTb7bAjMGywlwh0Qo/UNKhcoUuiGCdlYAHG/PeFFTHMGLu/aTet4LWqiYcvKL1
4uL1VIxx+x3xR4zvnD4lV12Yi4nhoCdeLVg5LDTfQceK5N5inWpXmoh5LjcVETUdi1aNqFQ/oQlT
/E+ZPXPjBA5Ed/i5owROQr/SngvvwGH0ii4fuByWN6HxHuZpjSVCwjBH83M0I16zDbRRKgNfQPIM
VOShmdpygG9wCyGnaQDNy2/YToK267ybaQhIJioi8a1YPVhaZGuLBJMuLUmtU6Cpa50jYWyaWUVI
7Vc/ZA3bz+iSDG4X6Xy+l6XJb68+eXxwLpyMYw76VJIG+UeIuAkP5kl7k8AZ2Z9B6kyWMGb+TrWu
hb9LLn8k0l8ONo4/OsR+CqO3llT6UawwjjgxVzn7JkctNYkWJIxNoZ4PfEagviY80J5ieeGOAwrj
TBA8UOKIhk9zNGpl2sCSz2zz3DyJL3ouZuJaY56ul4qwr0QZvNQL4YNRMCbo9Aryl5gDtzi4lBZF
SgN2kZIcDTSKU9uTSRNOoTj87ChxCn+rSMPkec8n7vJKRD4P9EEwyanKh6s/jx5Ny8eN98dlhO1v
MSgKx2rBp4f1+lxeewE1dfc7MGzhZoHFWV1Nubs3ptAjPYkiaGOKo9jEie35kNVun5/l1uL8Be8N
dXUKaYIz8jyeY3+QEFU+g/QDu6SHOHWBtgUe8UIYG3GlWsiEDe1eLxXkQ+mQPG/6PUv43CiC7IKR
EfpPxIUvlLttkZn/3B+4P+7rwCTp9n0FGfHaOknJo2XB/xlnphZScg/oCSEn/ogqGG/l4v6c/0MP
xxLOZdmXshiG1/kPMp+3qNJiDPqLkpGNRkGCu++og2qvkc4jTDUWGnNhAMocowEsi/6pBfgEePOb
c4nOlvrNmYC8FEcGBxKeir7H4D/ZD5F0v0BTa6Ai6ToLvNCoIrbhJr6dqJ9WGsVOwgUmZM1fgKo5
eV15GziBT4YN6g2TgA1PangSSyRMQKNo+h/2HFYZruo3P3nEFQE4BC+T6iGXz+n9LsKTFjaWnVKx
hAdVtR7unowwGy2UbYy7MLxU1oa0CZxjAyRZ2U7jrnPYIB4s7vvuVSjrYIPVpxrztd/rEaZmrODr
ZkAGC1dEFfsGMMmNblT6JNNe5Ftk0y5U2OBus+LAdumCwqvzlpjhNmFV1yvoGuES4brQStn3ox4Z
ILxRcaGuNeurY653Kd1kTmhA2GnvMCc6kzrzaSSaAuCDePqBizEnnJWa+PF9CYahJRDoW/VRabYl
c4Go6R4yn5yOoKPHMlS1W+10wLK9xA8t4xikpgMQVNdikeR5pLOtS5K7b5i4hq0fIY3vCNZhK5aY
gYRLovHD7zDMR9vFseQHfz61lNeD5mWhhnob5RSNf6/dj0jM4/THztwUixOsY7VVMwDaYhxfrJ7P
Zc0JFZJwGOLElvQLYjyfAhPduxCHS4StNU/hj93MnSm+M+9JV1+5d4dppjx3H3kGk6DObF368joK
P6l3xR8kFsSxAV4b+4aFh6OdGXc/hke5v+6AyKVdG6cbAwEOY2TO0k1lqKxmufnpUCDxr4v//cGr
OVzT66BuGMNGDbEd8NfbM6L1oAGI9vhgJMVyzTjtP+Kq+duYArIq6uJdj0+HSZeakr5L+Xlql787
n7iOoh9xv1PydtZkRPIKKtyI+NkdcPdgx6G9UZAwv5XaK1YC+TgOQeL+jZ9/uYyGS6xRM6GbFKnV
KkbQ8y1ltXMQRiJj7dLDqKgV4sZuna3pXrAefCKMzrassg7F2XwADEHqcvxCqXMYxnXfvD5lvmwr
qMVU9OyVr5jDv+mCYkrKA+1GRfWDLKI9rfK+uARHCr7qKoPxfNH9WuN3SsknKskh2tjgWDxWLnLz
dCF9t36H0AH7E/e7uw4M2onR+9nEQIgqSV1dOv9W8mCeaqkywEtw5B7IPdxya4YqedN+bnzwrS2y
LFFpQvU3Z2nYdZhguW1Mc2hZGM3IyMiwysys1ACRpohIJrOEI1l2hmlrmIK0SB1KsQPiWhPYVNsQ
4GdBJb+Ra9GyqjmR97JjxT3XqLsdwTmdQ6qY9uuF3QtyU2LS1mT4hwLIhuKfwvno/zPio/2ThRgR
axIUAFoQRxsxuoIiOa6pC6DHFFARERVaPC1ra19Qc3NvVdpVSfdKwC0GAoYZHZUagD0HdmxxkF49
kVi6IC44wbvtyzSA47RCkN0AXER8t4du5EEYgrK2I057znErJvx6uAtKLy6YMaaOg/LeAV77isJC
Jg/IkWrvktzYLJ5PVJ1wXi31OvMoiKceW/FvWKPVHiX79x8z6tkaKGEnQN0mqbQmxpHjNC5PiqUl
iu8XJkq7wl+Vux5hL2TicpjwYMUpgdxn56atdzYaWrXPkjPAaDHBSH7eoldGYMdp+xTnRm+ATSkG
qnypUDCGKaIJ+l+9Uu4zKUrJqDIa9L27NiRvzQzEDAko+ofPsjDLlWDod/9zbgeLCZGpURIaU/JG
z0bEzNwZX27nvYEj37L60UQ/+Y5GKzVokNFMBcUTybhDMMGb65Aq0gNAU47pGa0YCYRtrp71FrM0
25IT2GAxM2XcoIVRID99x6a9x/m3dOkmYa2IaPxrhus7NkQ6/FJZ7u3j6F3CrlguDrlUyQ/eGvDm
h3ekotQlKqms3OCuYXafM8fMTA5z/k89IzlRYJpedii/ObbzDXDUWGXBTpwgbzIUaf/aJRpiXUOM
xN7FA8M9wr7ahdwAd2+GXLt6MsPMTklL0XfuJKqtEzOJJBvnTpEPEliYkt5a92P4o8k5uLFRTuDt
FzmAu+eGprbS6Bm8yYwApn/fUqP/2GjYaRfks2hbsGalUEPHRjKvYt2m5PzbNyiQmA9Cesa5BlNZ
8vU+AvAeoHkjOOSuJlIHW5B2ftNofs6hXJNzltEF0FWd4S0fopmbrv5U3KNC4SF46QZ8PWAfF9AV
IiU+0RBXgK+WYUQrJdvZot5RHmxC5i593yKCtsHIc+3H+wKhvfaycZRxTh5qog2cntIYETDxeGiz
em4ts0MU27Y/7UTYNleYK10D7uqRRHX1tI/n/AdGavKLrtz0xqmM1E51XKRz2/P7EvqdxLVb566w
BNXJSkYIVH497FTTaKSqOmtcnUQ4rfa26KI2Hz3RruqL9fqWMjcBaGhSCEVLtT5RUeNtWh2khlDB
8Z2nm7l4XlSJbRAAbfKmMHOP8IdIytqKplrdgjHuALWJbr2S1yTdfnLIkigFcc7tdJYYu1CP/5RY
ZSKmSxmEea2dYLLg7tpIy9EP5O2+yTGEyQCGpMZTuCmIi/qEjruUC7ITCnqkEh+2fO7b4t/PZB4g
wiqOpWyxiJ+bbs2DwSAB80wUpgCXlbkn9HCvJ7QygvfH9I2cWBbO4TaJ/UMfDnmcup91Vhi/WdT0
oeYz+OUD+vy4/XU54XCCKCptENIecOKljwCqSNIhx3lhwhMTOors470gKTF7shnQCcqpqobA5cpN
nDfYqzlCI9aWlgL4W7IWSpM4ZvtmwLuHqI437f6EBFjj7cFvHw7ebBy8/c2aRY0B1+omf1bhsInh
z8oF6rR9/zQCy1yFqpJJpMO92ogFc2sc5KfqrkSoStk89Z+CtXh3lVShE8joO0UOEqGO2lLu5TbJ
1IQgWDMU94vEIjOcY71d0K3m94mrLVae+rvv2JRlFaqT9mwrqV9HdKjBvL+xCxDIrIqGDPgtA5V/
LIRigXqnGnWPFOl+L4X/m/7jknH5DJ58Sttl1rdqMnjOrbbuj3QoE/JC9IYojcOuuhN2sNXBrAiJ
gKnJti+d2d18e1GSE4zNScuymosGzBb51AsdRQDO8Van7SWcMATabNszeOGzuR93oYNl2NNsjb0O
FzkpYMrtGjKhu+fZkRhZsJpR4mZ4jBuPHQ/Sslb+oFooPR5HG+Ists36NmJT3/620tkmJeWScDx6
cYvsK+3gopJxT903goEk7AVePT5OC8L01xMoe4k4D3y88GkwZ4BOjKEjia8GJrpYNftl145J50+a
piTowqsGcOUFNM8B9m0pUgTja+s0JCisaiQy3aQu23NvidOP09iMRtE3hXgj3ue2AbBR2HG73WE9
G6t+9l/jtz6wwg0oK2w5w5XVQkJ3sYY9FdB04p+TTGfDMJWEi4yvSUM2ddBQuoz4kEI1wlTLwlib
1Id9JiljPkqYN++RBy8RXmJKr++CVqp+704G8nMytRaJ60IEvjzNiAWc4RXrXO7+YOTbEyqw2DhY
zOzNEREOdM9k+/twJGHgAOCD5dvcOq5vlRj+LFdYjEB2uDB+uZW2E2YbwMfGtW/fYT1cwMNP/mab
8EbU3AwLL9BnF3TJf4ahl23rISVdNh0dgEJUbY6SyaYf9SgFYg9OEisUOl+5eHNob47mtIQEI8K7
X/fKdYbdteLh6Xx+N8GCtaxpjRo1GJzetmGGkgv+Qzej/2oB7x459z2IYjTa/PcFBybpdHkDJdez
ao5KmJMhVtHKAdWMwmX8SbDI53LNjd/KMg+M+SI0pCYmAqDj6R+8YoeUBO1yDGmmgYXMyxS7waKr
tSE5eRGWRUs2heU0AaYqs02kQ9PqqCIY0hQwf5enq8T6rsS5nRzDU2AGi0Dv1+rBfa73ANKkKpN7
/G+Ctt9kqMVA0hRqelYbsZ86GJHU86pVSV08cLX1q5yKAHN7NT4cCesuZy16DD7WVXsJwgMqFWX+
9e004PX9uMdSryb7Tf8eszYiuAGF6/AqIJSQTxwmEGVx1WsZO6YUGKM0D41b55ktBBfIznsnHQcI
U2goIIwgTB2Quxr8PeEOFzVxQr8Nktxdy/wiBPmpKWPZqKBhm7W6QMnOoQI1JVTd/AlBy4lh5VaD
sNeI4wRZSFVo8vut7Y8jVpeWQlf80aT5lJZ0EktRitz9gQOl/NZR80Mg+t2KYc1lANCZ8E6UPpK9
MmStTwrXknDZHaLT5Qq7UGZLSquey7E01Ow+kN6QTNxTZlT4MV/8nHcTswpvRuiq1ynHhnMRuZKh
/9pnozGvheVo7PL47+0PaEMFR95I7BSpEWmy6HWhDSuoKeYj9t6Fd+5VPuqObBuvO2ObFLu+mmCx
fP0oK7MmtKwIzaX/zKOvvb3k2Bh6gBHZepTsWVVgNbSilQ3igOOPzLS7kVdDsX1bHPZ85BloHkt9
Q3LRN97a1dt9saY5Xx7bb1ioQ1hpTpo5Tx55UNtpYbS6t3eylPLi+LxKvpyRgfGaeEGbMb0zHXqx
pnauZWet0x8cNyrQYTUOdg0UU25Nd7pB1ymle9lZ/hhBvxjMKaRxDYjX2ME8zmYJSu6HmlLVVMeN
1KtZLZtp1irozbPxr+/o7l7znquNJEYZl4GK+l2ws6WFC/+LiGTJnXfCvVXkpbeE7Ep+VByhlPdk
sBhfKkTb2UzCAV8Qefe8HRrXFkQu3mUpad7Wcazqr1v/0a2uKA768gRQrGY2a7osiQyIvckvRSX/
R0PFLkikoSgrklsa1iw7u/qsgow3VEdhmRCp37RtWY1hjrWX+gfcMsw1mG5LqqHvQQgqqgkryzM+
o7llBEL5MQYhhi3YgkkDYPjJFzdCt1ZEj4kUQYMrz/zZLVq2yjx+156hZnl2qtUZyiImEc/uewfj
X3Ls4WGME3M/CVNgsr951dlYXxtAPkWuhmU+1fFWbOaY1FaFdIbMGJxuDiOjSimg+WQQTHg4em83
gAWa4B41dD/KpqflA5ZAihgwEiVrbIO17Ba3fl32JphZ946kNp/MTWLYGG43YGoQ/jsipUUo0aI6
EM+hk/g4F2SwV3e48IOyMFmMQhi/+Y1lPKhcDCGTZDI+skDvBDuJNq0rXa1hyp2OIji0+DLFTT8/
dHVVSZjTDdszBiEIAUUdetXNlrE6LAXPZMY1PHKp30E+B4/i/bDfRx+/+h6QFPzeUWSvyawYpEE0
/fqx/fOCBuU23FaQggSNkh88Mrp78XO5DMMzUqjCqiyJ0GzZrwA2414q5KEZYkCXeQhzoicLyrj+
Nx42mjq3rawrlQAW2hpg7reeK8shrR+cSQ68OM35i12WcLDVw0PIa5Dm1rCMbYdE2IzB3e4ToSJ4
kuOKI1cK+tlHZ5tPduvNPaTIeKF56j66XzgyiB7c81p1PApXPinocI2/ujNFhKMwYtM12SaFexs+
Gp2EV8lUnAbcZfYEVm6QjKR4ceqwmlTYZTbs3+krdgYg/QO4vwSNRiAq4qQuwpIHS+SEReFEZtNi
S+RR9cDPVEHg0iI+Ub9w+KI5rJ41hl7CbMC/iooLYNxbIeKeXg2jS32/aU9gFMqhMExZHIMXRMr1
OF8j3jjJXpcJEtc0HvQFRcq0vy9/dd+CUJMHxbdn8KFOK2qeMhn+v85m0Btcx7crbhX9uXhH8G94
W7psLeE2JGw5Ltatu2zUCDVAgnldmnJWe/gXRShx5h65ENDBkHeQzXw8W0rLjE7Bv2S627P09KLu
gNYND5CkoSBDobFvCt/Fw/9YVyqnVVE5dSZ4HLrh6K5MJ5UPRzoIMDPxMeLDWzC6iDBs7UIJEi6d
G8n58T127h/67lfUTZApdbtI6w024o1kt1YoGP92EJDtSbYoBcDSVgkXzNn8p3os7+rfDyI0Ws1z
bAmurCsR1IWoij8eK84TcC6j5irIK7TiTERZzjwp8k3+CgY2cRtuPlurpcpUZTKQf4RxEg452obd
1mDSAnuc1lqEWzruc2PVUJMgM3JCIQLk3XQ/joGqsMohU4rutGBaiJ8UwMFGpaeXVeVB1FaK28qo
JnzcrF3RKnZD9LlMBAqj2jE9arICFCxMWAF05m05thZkLxSJFRheUPcIMjq4uEzgX9FSBd8jHh8l
sFh+Ub5FE7j8Gw+zfXR/mRPeO6OileDV1K5FL+6/J6xzaM+19hokdJ3N+P+894EQ2YWGEHrihxMf
Gi7C5abtkYw9H/nMAIpcO9xJTQ7HYzZsN0WqG2OrfA3SgNj++IJAX6UHDPSKkPbBrNbuCqfugl6S
21+MNUJSEpB9GHu2igUBBiCyBW0aFWTeyNoBCUC9Z4pF/K7YN5fX3v3/aL6qfwwR/hMDy1nZ8Z5w
4kezdTmsreyKTgKOaCH/n75ct/LRVYiblMj5amm/H2eLvJpfpguY54da6n1XjdMnFN1HkDzd8oj7
wZ1eOSSmq4yESMvqaUrqkWOhzric0nj/uYE4NT2xcFnOI0FVIAKKXUQk4qiM34MztwTn6MWKewyb
txKrVHigG9NmcrWyqWADJ8ogmhPbL+nR89/H7YMtueIRQ0I/beBIWdjDg+YTvFJFaSVCukz3gEKj
TdENJVP5cKUDZ/UVE2WiBsCdIlVkYs0O9TsMxzGjCeZfJ3hagcBMD88blSv7+RU54rbcGrRc0+Ph
VUTOYG05+f2lsz4/RgR0RRWkzAWhI+9xGd0dbW+/VIWicIk8hxItEYp8Ca25G7SNFAT1GSk7PPfY
SEoVlPwDYKjcfcd2D+kARoAWKYi5ULSvmoDNSxmVlhxJNrWEyM9iZVvCbLr6t33x2qLlaxhfNlYC
BonFXzZ3sAEUiNI/wy702RWAjV/s7828MYPkPEi+vFxl3SxZy2t7VPO87sbgluGzo+2mcsIAmZjK
QHVjRmZP0LnNSg0yA4JPg2H96zg9VolXzXXbHUwYvFdMKzntcNvWx0bFzy8Z3Wp2WbolFPBM/tWQ
yCiBwsOLKQEz5Tkf/eqtFtKpU7myDVzC0UJ4w5QupO/FmqeUXKpjrilGeIUepPTsg/gh+ngUm/Hk
x78GBRuADzUvHZulfzNylCblB37lhPEOhMnq6sABvgagbeRtlMclDemBv611Vbx7GpAQcOVUUa2S
1fuXsLNfdfzz8j2MkcOyUsCJd+s5df0PnojTyQb1nSYHLWzB1qtpyPtnPozmaz1nSbI4dtQoH6h6
xLE/GnF1OsSVErWQSI+a1SWRQPAfKzwBRBqVGNSRKgtbYyq+LiLjCnfGeRjRtpFU32y+I896EfLf
xoWPg6jRuT1T2mvHb7v88F8/iBxpEcEBB7pDabEipw6yh5DlAlNWwBvpFELuf2l5mCdguPwOtlkA
hwVbE9emme2H9c/hTyEIPZdwsFDmn6raHtTPXs5otzKcg6bPumos3AA21IQqlhxOd9uoWou/8LGS
85hlTRD6G++nWOkIo3oN/YBRX5Xn0lfGRuujIGGVzJIocqsbUc31MK4OuKEaGmrnExdmYwZ0fFi3
Wzlo66cmrHXuO3NkiKu6UfLtuOshwyWKNY5wXh+wL1DjYdtT4nYhl4dPAyvRvUu0zPXJrhMN8ocK
4KsbCCTwCqagv1AdzqeUF6IX4bpuyLPVjXKXvP/OvNnpC6JWlbD8swBi6onQnPVL7ZkcGWHX78a9
97iOfW0QnCuElO2v1MnMDxBI5NWRMijNFWTgYb5GRtzVPuX3Cq+GJbLhGSIR+ZK2/6pWGNmKfL/M
mHoTtzbuRtsVJKT2pOkuw9e+JqtyCR/vQmlKrh0HWOXyj7CfxYD5untTOOiyiR37l9zugamfq7Dh
0yZIFpR3f/qOn8nfRygkWqt2oD7Uwa9ARRP2xtRV0T4PYLBNz1Ef4iIEl1symxVE+o8GGbvEDvHV
eZ6jA1e2CV+vKCC3gXum2jOSawhVWv2yAyfsrif39iJPKo1DqUMQfO4TBf7d9uXZ4ER66ojVbVvM
5dhRI4hPWDNUNZV0WWiCsT7xCUFOdT0zp8G4SELee5Mq+o2+6qX3lIu1dX/3GQ5mUgiaLF533eGS
LC1D+uE98ltW5eEnms45/RSmAz3wdQ6vnv+PlRFhDwGjC4vGQ43lrtAwhPc5Gb++igmV6QTVpJnC
Nfc8p6Wu7qYArAmwLEjxdXWUtOnnF09zSfJczFRQj+7Fcp3NsKfEmiDI//XZjR2FnmjfvlSHJ5yn
wntAtvyZgPRLrnrpU20SuCCIHHsMC+dpQQKqnbtdOi7omqqXc2zzrl7AKhDS7wzI+DH7FHdAFnlN
RwJpie999MQZ51EPO5zXJF9coz3SQOynXavygRLj7QxpTbL38plVoJ3erkJ3IID3IS8yPIr2mW2/
Svqf7+IoahP+vZuv9WgqqDTsxcKjyn/lOkAJdsk6EZ7GnibiP1+xTWim7DO+hWWpVyQD+xBVfq6z
3u2p0GZ3oZsThQ6U8zAr03kJXxlRhHQT7g3/a25RffghgjtGupZMpXUxfjy0gZb0p/KNqEPJHG+7
cv2YGegocUKP7k1AfVp/qa26fVRRhDHdu/OF06nRUo37mq9YRO2Na+UbohDQT7gDujbJ2wy49IAQ
BiqDp1gqWL7qRjj+Wh3MxcKQ09D4/jpehRhGuJchYKy2h7m9L+6q1+PI/NPf7AVgvLDiMuIix2C7
FZ84Rza8brZT1DFpop0Dg63+Gf472dDKXdjlo9wvaNtFtQrKZ35jNzOkAcK2rv7TSlvFKRqITeVH
a3NQbZaDVaPVBJxMUbemxvfuES67ugQPkX7F8IbMzR2IO+Rwm2LU+Ylzu4+QxLHdfJ9qziUpUN/g
Gnp3UopFq+gMEhmBV3ZE2bUbsWW4mehrSz89ch2oZMjUU55jZbJhDTYd+9z+RTjt1H/Ft5Ua69az
VN7rlwaxRQ9/RScOJRrv3s5GMo/ym7fkqDWCtN0YM8eM2T+zUl4R75Z4SauohXu/omza4VwVMgQa
JJzuMJTs+pV/WVps+A68iNctb+pI4WdWHXyMcNmQjAJCwb372zizMoNkj6O8MbbLV33mVh9rKyZK
wvhpxMtD+sLwN+pUcAQfJE8q4L66raRSDBGCAve1qNwxuRxQfBDWXOMjBDwOpONv4I2UqD6Y6UlH
XG149NaRKHcOB11QxVrL6bTBIbAGgQyV+ntcamOeP3PeSvXxcFbLbp1SuUHNgK+AwTj16j7Qfkf+
6KBv7wuR/6y605LIlu5iPg+RfNxWF0V6edub22Spjfbxy42dAsmKx1Xeou0AmyzdwwIkX2YbBz8o
odkU34Lv8iTdZ+4Rrfp5xFeujMrPTMCFpFzyOhw9uPRMGmnQL3Y/TIuz/0K+YMpqhZSdUsCHdrXI
Tsgi1hlGXwVXEWjQkPVlw2mv4K7/G1GsmMbNMtkr7Be9fd4vAXjhUkQUguaR2gmTECLQElTafb/W
bQMyx0K9IrLD2lvdRWIi9kMcqfavYSol1Qlh6yxXos27vy3kJww9DxSzXvVT8qcdSj/ro9yfNwl7
CkP+33CJkN4X+psUrWUyBxDFh0pS3HOgf4NEfQySJth84QlcxNKt5qC+GoejwBV5K5sSW7rmZmNS
Jw5ebF3sAeg3yK70CD0Bfg2LNVZOyw6UMYIfuvnDFjvjxoVi8h1fncIOpE5FEcBjH2hUCpm6Laft
TqmO80LQx1hX8V8ZDF9VkuqitW2u2Pb+wcVZm0iH1tAUS3c0ycjfhlZuxy8xDg3CAslLeBJMDn8n
uZohKSuQfCL56Zy/Q2xYcEcfOU4qH7BWDnBqOLDAYxNNuwYy8abPt9nbPv/w8sE11TcSu5DrfUvw
J5jXkALRPyiSh+lLJz/q9vIsbVpgrqOpvmB9jYGD+f0tp9XkVzuAtfai+R7l6avNi8W7EHQdwLeF
Tq1XwVYVpyyaxMf/nZL+QxkxGxqK5h9YWtxj4r6nAZfwABcAj6sZ0aJ7iFqJEp3Tc6garZOjFbjo
DnRwQsBLAYRtcFvjMG4gRwWHYq4UwfhA4CE+7QqY77CvJFSGTyqKIyLyo02gzLNNQO4WRazn9F9G
NAwcMfM1eNWTtzTwmwbdL19+7Y1rXYUkxW8VrF7vPtINwKbUW8SgWhJVU8rM5gjsQTK0xaVUoBfP
6Sy3Lil0iGZgP4m97meKPaCNlXAD81MyOLNNjTx17CH9kCtlFO182FnyLbJAqGQvtoZxAPKnsQz3
G9jb+AV3W5smm4Lcp743r77OVzc4Tvpfj4YPijIzxxVLb3nR2yuod6inoI6UTfTxjFxEfiJNzkB+
uPYlaYH7WfX4IaRER0uMGZW5Yxf5V0QMF7nPXSZUr8NkSsIn+Bq4CQJw4WgMUwguLQVi0hp6XsyN
z1j8lOc54WU2+xUBH9m7sxNPwppuc39lbot4ztUKQ0xBV+SruwF87WlECKFmL2Kz3q9Le/fTqfgs
F/sDtWq82R+4qNQub30oObN9ViGjK6RwoI7yln2rOyNYkkgSXtJVb/XK20Kb1/IVsQHozdVwntQh
YRirmDzcnqxmlSzleZCHW2JAa22TNay4Bs/TwQmky9booC7/Z5iotxzRvfp258tIDdG46cqcZEqT
5z7Ofq7LVYDAmQ7U6OXTG5BdeYNC10p72ytszDxJAkuShhJKkd/B75fLDYx6TuhWih1iw6kCPV1G
O+L9VlxUrrYcoSVHwIjlqL3Ad+Jo03yt4J/9A5JSi62D6HscVEufnQCo8XX/Yzllmfd9ouZDiKlq
wg+449zpzjcz8BI7obMBP8AG1ZJiJ/tY0M7T0VJLKdttjmg86LX7IfDGIADXtKz6eVj1/dD8hfVr
NbH6EIUezg1uAWam2A16RZclTJpTNLlCxS5hVBsxGIObk5zoDoJM8mo3DLuWT7x4c/NcJ3YF0wEs
i3fO6ln6AEftLsE0318E4Q1boLEL8LZosgg21buCnTjzJksKfifl6s1YFapoZUDxAvCTDKiolVSO
lJ0Bp/vWcS8Ieo2cD9bGOTS14H2gDLB37fLN5iU0Zzp523su9Rnw6HWc13b2Tx8YkLeiVXuAt9tt
jGPBkKXvfAKYM6pb/NBj7S5Aa55YV8VUoTofo93Ajavri4MnVmJb3TEfhq9r6M5WaZcmrxvKK9oF
PKR6Uo+ASEKK+giWK4zxPiC2wcp8N7/eMsDV0VsufJ80z2kVtHw2y1fEtOIF5Fyb4oXZ00spsVT1
B63RVI1brCIDpKiNUfA0RIRu/4kXxS8cx8rhjpP72iamT48GEyzXwf03v/KqQrTgn6tTfNg02/QR
9QnmoZlZowgVQxYwd6ozvHqvDASj3QuUUjYiDlSqqydW/HkIO5zF9YFh9lp2dFwtOCrz2FWt7H0S
RUHBU+xugnJsvNWgpWk8cx9Dz9hHQUyGLSF3qnkc4rDnp1YRMHzv4BUZw0CkygNVW2MKbje3G+Xm
58F18Fj4vUQW5vhkHx2ecpUcr5Bsmf+skkziVnkGYmMbOHDaWC37r6B5q2KLqG2YOhZ0I5CdHWPe
ucpS69GOLP6MXhhSNVznOxsABJM6MJaG0DRD/4WLgpwfPQGWl4U+OKcpZL5FZX8EHoVXCpz3SajC
/bz6rb6r8jSzIo1HzRnjlDh+hSnU/rTFmBLmp0l9Gb4q5IZcppw1OGafbYXliC5fza4FBJ6A+Wjg
96mgxD0ElfSFcqMkNlE7N2pp04H92w45S8XAUKwWcXif8bcoKtGiHcUolKW9AQA/iPrCiiFtrm9A
iGF96p8pMG7wSQ9s1f9q2dSKji90O2rJ87+hqQp4Ok8mQhpP07GyZ2rgo+UNws3I5aSVNdZVEZ6A
tFfZsTUXvrOP5Dpj/FpIsLn6xjwEAHBZkrMRtHi9TbKWhdlFEptRcCqLiVeEXVvrSutfhPIgq2Y6
oGmEP1yIlIlVwPnDcvBwJszrtcdMQet5n/OCpFVYXopUB+BJwcZeDa0am6XiFZbwAAyjQ/kOeW6y
YmsolAO4YWvnwGAeNBtF4F2wetMC4WbgY2qJr1LlezxWEcItLsXp7A+VvWcBf3e0JYvIxGFz+fKG
2THry6dwbzQGIOBC57kA81zIObSxJ0WMZreM+fxHwdXkCUQ7De2nVuRCwZ8OUfx/K1IIZA8qruwA
1htGBP91BLVOE05guv9N0V3l0eDyh6iRLRwSxCzQDAh0ddfJzEwrEDGn4lL3HnQ4CnXVtu2D9MTa
o924c1kGNp5z/6+lHepqKOMbpk/Gq7SLJQYGBrht8mEuC670qjtYsaRXmRxhvjZH/cL8CrJZyLp1
49m0faQqyWdyRd6flPD44actexO0QM92IvetUh00MHJkAc5wfgTRF6raP7k3CXxqIFrZaV9gp6uG
TT/8Y6fkuhEA2N6pyIw8vMpkNOljTIGOMlKCAlGU+e+BPnrHTNfOaz1bxgLGdiXKyms9C2zQCONz
yYMaaFQjUXdXwrZ9bNP5vIMuHVekcaruV3p46eYCAbYMZJCKe7wCx/HSzJJYzShW5Xhy4XBhbEGt
YJCGj45xTBd/qmeRTNGDb7dMEXU0SQb0ZVOpSv6uhjNqcaAG0S0VW62pTwEN/NlJu3KQFm58/hVk
DYrRXAx7GYTLtUtIglhz7tcW6ervzBCoOU+W0gpkTuFTIS9KRSwHhvozZllqPRSTErTqRYoOqiYe
BnZ2rWGgoGCa48cp+dkoiNOxHW9NRWzqtRT1fMmJwaVURTRQMNbEhVdxv827bZWe6uGtvOHqisW+
EwVYf4eePWRSaMKOA/w96NMXPlWyXLNP2zM7Emjx0fnNwOVH/0/bU3y4+eM7QenajXAVM/hfr2XS
R2PZezey/Nv+7dm9eRzTYMop+KgVhaE3GlX8DhF06V7yxNkYoivevLy7+8Yfps3QAxfWfe7GJgyK
9eWYX/UDCqfnChxQ8+cyxcctESFxIaEuGuvpdw+P7eQuB2CFF+8AprMcK1T/83OlzIq4d1kYE8H9
vE1LSxJ9b9XYzCFyQxUOZzzAZoWCT4RQZIK9Lu8SJD0x0vcczcw+pfYuLaHB57LIO8/w7pcFi5sL
YFWUvAfSKIGikCx1DQraor3061lVGgfCuFv/jPuS7bqQnjndJ65Xupl8rbAMjaQVAwiVf+BTt5l0
JEsPLRzp320jv8JR0Y0WAGVRhA90YIjDRYC6gW3L4kFDyFjYwUru6Opi0p9RH6+5S17+w3Y/0FwB
3NmEpgJFrgHoDJB7SvSBxLQW66XqS5aeh7FLvWLMd9UsiDVXx5uRQzljvqMPj6UrWKpdrm1ZEKiF
mCjSqmv7E014rxul873P1Jgt06UX8Gs/lViJcdXodMtJxhd5uZOzT1Zq5lwj+gwXpq7XqSJUhOSf
017KfX7+Gjih9DxK998LBuLUWAYVCXGtCWb6BgdtoAPJwHpEI/ECBBk3yztSG7vLjlkDwXbXf9t6
uZYBPMrW/5JWcAmxQfOvetrDI0OeD3k+OSEyn6U/e4VzI/VZvRbYb74oyPmAJoVNuNHByEr7A8Of
M1WSENPf0g6xygKRJZYQSxFUgEA0M+hdyUV/eXFkJExsvzyao4ZLD7Lfj1x8mCGEUsxq0s7YGHD7
8FUDc2klC+xfQ02frmI9hTVfsSkJ2yHwOPJwKLgrVnqNszLP4bP7T7OnieiwTyb7UJjhzYTZmcKv
G7gmWOIQenz9XlHmRyES4G7XZA40B3kZ/hKhc+Z9AJyYEs29NywF5vMRuXlLIWrbMOcudCpIm149
JJP/nqgtfZF9eCgVFgp7e6nQBQoPJYQLYUhtVWfDnUFbdSCkl7VuRSk+uqIjzKJ/2ZRCyLxDp0//
q2kUf+Fu4O+exlddnxy+coT3JsNPW+zjT98tTzGfLiEiXQjukodktAa07n4PDBKbv0UsPRmJVPqw
J3Yqhatu6oeDUiku3svpVNM/2hsM/6J+TETRIiidkU+gCKVFhxJEgCl6whfEYn2GCPOQTDRpUUN4
s5wPWEHS8XhzS/cdZrmv0dlVM1KRIKh5e8ZUXXpIS6r1Ae0ddOqgulTdVD8CNRbBooMdsVU5TGhk
3bDb22nX6SH+cF1GH6PGiV2OcI4ms4v6SJDGvMD2Z+kliGMwoMVjnw1IkN5UoPKEqLUMaAkoGYYH
u2qtTabViu/hBwgNJReONYw1qVb6MS/BprP1xdzF3FzgGzJRKPA1B54C2yDILehiM5+CAAWYOXCN
hyhjF+G2bRK3yNG19XI/88COpPP6zmEaN5fi82sFnGZ8nxA/HN7diTy8FZV3l6vd82hhQmNrzoyX
kNi/eG0qaNspcCdz6nQG8mvt4tG+Fy1HCfxabuhTwj09RYvLLngRwLuh1m9qmSOPkjfb1eJw+Auv
/0h+9Y2o3Phk26qvg4OnWM1lmGLLRKt0Qs4eSWQJpDV+Vwq5SdauIMa+NhmBhXGWLP9DX4MmP4SF
HpSbetA3CCrAOljY7xU1EZE/1jm2M6YkxpNpCWxI8ZZNszxLVuqkA5oIW5oghsZlx17r4rqJkSFh
Tu4YWDrKHJ3/F3oVQSa31tD1duMhshugWsvoMwAFiAShTdOAPZCvGzuEqmNnlgPFkG7b0m+fGuBY
V9FQohBUg178lz13vk4A6roijFXke35Jh/tM/7VWf5axv23vsxxSEG8VIf9TJoSckT6MaTlSK8Ym
qLHJ/puS3CLjUCSPI1fHpYeXf/7oFxagoirNDvdueMs5zTqMin+f5wzMRfRNQICeDVbAVAKaOI8w
/j+APfWlbHWEfg2uBk10NqQ65oWn09xC5imKGVBQPu9GNBWNo8SZxYWqivhtHuBVohouryfJI5J6
LQS9VaU6wZ4ThwvITX1LtIaAE8in1FKlbrXtgcROgS+inLdVYvBout76VF0D8EHM85FSfqIdXBMA
66qNTx2ZPJskleRZe6OWx2/LkTm/LOnvbCgVST07gXsQbHRZ/vu+hqBlqOHVvlsPDsf4DWpikZgz
mkSIDRKKn2ritl1AXwSeRfGqYmdZ83UILNbwX9tJTnhmhUcVncKSYK+XYQeiAHbEu/wTxbsAKoBV
/G+e5RSHfAz2EVT2MvTd2vow1O4Mbtl2mxIy9zj1iqG2QX4AzAvDgZQ6PXrtTf5FsHLS1Ix4avZL
DCw/6uSMd2PacV6muKpQFG9OQ7CxJTBxwry6nL8KAiTGmVYs2DWOFP4tzjxikpWGB1QKHqib/bL/
nbv8eKIp3gCLYWX5DzMpsgiFkUdYzXQiNXmIZ24Me3Wu+9qatb+Z+fXlk7JNuBYritVyUS/tq6bn
zmhV8vfVZDtPH5WnOKbuCXGIQS+cFCQu9DNT+VPlGEhHGPwmhfiy1T/eLqR9VetCcM5notyda3Ek
VP4a/14snKiwZ82/fOwSMm2ZnsxJYTE60kqr3YPq+vlGRdOct0zilmMhHbemtFRW8sNJ4YIKAY2n
maCE8avfsjuGoeXJMt4XUlY3Vsotgivj7JJhP3XMKBGOEMI4oQ0MBIBF2cW/WtbI3YKCSFHjPYKc
IJiOb9sqsAwykMDwN3chnQ4Q8o2eC3EXyTP8QtUy4je1ZnOCAmUJjXsmuiSD3N4A4RCunwivO7M2
CZjKUnPuDrDAqVHkWV0OMPTIYLy64B0748wW/Mc50LH/z7GkCp0efqa+NQ2HRyJyEqmBvaQPgE3M
iT6Med3Qq0dy1H7TSxhzw5UIn+qPN4Txh0rR2UC5kD1Kai0Hm+ZNQrhu6h0/B+Gz/F13TCeFoLdT
NtNkFym2gdeVDJ8/Ma6bHhEHtZpp7kFtERzYBGLaRrAW+0LWHn4arNz9CZmKFSVi7aHivgS82WyE
nFm7xObh/psPU6COUCMoXoUv2D7QgzH7R0SfTjoP/VTRigDPV3DT+JlTd4/2d++367NewzQ9Q10O
4Y0htkjENyczpxlJsvxJfyImONugzTkmoYk7nE10FRkArepAu+na782GYZQM+bLfmprxm4UjX9C/
XMY/KbZu/h9Lo+ZmbmXWpCBje/Bx9AT7Ej9LgHshsCNE9XFua/69fs7piStSkbrTdx6bDm39ZGg0
FqnAI2yV514bmYqW8Rj1vY3A7y7kj9q2/J8W4NVZXfwCZOXS2KeRB49lBxCkiL8wlJI+4n+jYzDm
Mfpm/7SrpfFb0a+RtNOcTizJ0gouEeUZ0Dl+Wc1wsFoxgSTjz7VdDI+xNK1N5O11m8uhtF2Q7TFv
DRnLz2Z+FCTsXY+bdMCnlPXa26b7ltwvGmccfccqK0pRwhJzqOjmQJ5VyVLJ7sJdDzIZsxvz6Efh
ykO87V1C1FMYiBNpInrFUnK5vJIcaeYJBy7zBKDFJmcw1/DwbQfNCc8bsqDxlAHDSXRfqoVNp/C8
SBdB1iB9Tl+7dGaTg96SbslJYq/u1HfW0hOiJAVLMqx7EaMS9i0ERBA+xhIZfR9pHymrBi4GAgcF
VxP+2SK/JiASJL0jWxEuxwCpJXT1zv8QqIlP7bIXhdME5amcUWbTDTIsGTAEQpVvr/j4AH4hG/Gp
3Sgq/8dpOymGLZuvbYWTRJ/szO2izENrDDjUm5BUBhCmAtYgThn8KVapgAASLI51KMdV6Ok/xUhp
KSO8keB7AqZ/ArcUlVvWayPN4HHLMunImVLUMQZ0lNGBQdvvRcmNVYfa28G9dTauqzchg85nFNix
7mK7y/9aGsloPyqnuHzzlIWDW2cFRHM0vMoNZRB+Yfci3KOH1o558LYl+Pi6Z/NLHaQE4COayt+n
koC7fImdGqiIYaiJjkg3YQUhbz72jaTsjabiwbeIi8+0gw3FbIn+VuUsvu5nKmLoQJZqEP5qim6A
HNMOZd1Uk27HEM6XkOs7dN12Mg/jk5ScczbKOdqJLT7YWGCEBfg2hjV1d+nWqKJ3OpGRP8ftCHjA
Q8JGHzfJ2oMxBUQ0gLWXMpwGmX99fr0ZgpC/3CvOyP7dkK0UJwtb+A9btKq9DqR5dR8JmaTqI0eg
deeHt8sh3Bn3By4yHqZmeLI0ttze9asMkUA238FVnImtHa+aT3P3w+14BsBgwyQYlip7UGycg+1L
7tu4cuvPu9FLVS+4fS860JxpH+O7d5CB/b7nkpcP7b4MffKoRZBnX4F23cQT4isevL+C5w5HYhk1
FN4TaGAqlsv9LZpJnE2sErhO/AiJUgho79sDYzXowL+NlzdS0SOTaCn4z6/gbvX0K0UefI4IBUdw
ZoAYu1Hn3oDbDHHfe03DN3EfE7LdsaLUb09i80wB3QzexyEAt/KY9345POjMYo0CsOiLHpIcBskY
7mI/ANRVjDZLq8/N3uoiZTUZGCK1Ts6feRwzra1qmgg1WrmJh0getab2LCCOVd30xr68mOku5yaM
HT76AIhYzTZ3vAJ+MGAJTxWPwRM/6A6q849L34nL+wOPmOb4BBqFcVd/MXNWYCMUAh54QOTWsGZY
0c+wgz1tkrFdZ/gILzSjv6sDxUXlhQI8pRZTTnoo++92J6a0ZCc9Fd05YyL8ucbdwhpI6KgS/jJ6
t49e87WpO96UqnhPjyZRx7MzMgFAExQ28UjfqEoNzXyL16hf/UT7fONgN4zzbsYRgjMIuUVAdhm0
rp/JtmKKaW9so20Hmi6fKDcx1QDuXJV6AIm1u3CLXiXLPlgB5vOuOSr0JIy492qieNINOI/W8c6r
iWseaeEVNH4KoYw5ryio3btNEPAtv73nbiIfVHOfxNMnvgYZX1JQfrZPee/UAHLjTlVD9EPDxA+q
YAWV925EsHGWO1DDCHP3WyAx0DwRRV2FWXLQGvd2WSXqgzptN6wyEoOcBPTcPAEyic5WzCd0z3fI
mlsEbP+3DQ33csMnQCX4IF95pLN2sRJ5U+bNoqFVSkJe5nJm3RA8fvEhUuXpc04cw7jid9PLJoXz
XjlY27RsNQgstdqDsHFL0oQzuy+UYJQMsst9Ri3dyf3vK39w8/jhO4keFIPy1x5sAAVPkRHE5p0V
bwODrS+pJWZOZTS1zLSkUzouDAEp9xNy4J7zbHLSz29+9Uw1XbVZ0zaEHSjw0QJoA6Q8idqs42k6
WWAlvrFY536BGQU/onWV6m4uHfIj4pXPFNbstfgUTWvR2ijAIzrnvgQESKaCCm6c2GQAoKVHPwdA
WWAP3YDN1oyE0+eksvuroudt9LAwrisR0YGhmeEIJhLFqjFKJJgZ6j37O/3O8iBbkeiP5J0DPylt
rc8r1upalcWevvMiDcJJElVrlSXHx2ZMUKJ2/2jQdFFxySwgZFCnqY+68ThH4Kwq84BnicUKx2g5
39Jnuu4aaLMh/WZp7KTYzuTUw9NjU/oIQhf51+DGgeTD5VDN42gzTwf2xfUpNGhTjVMgf5LAgpml
WVOrReayVG1gGzqLkxemiVpLybIBdXObUap+rLfPG0c6dZ+wbbqYyrHGSn6cElbDVEtSyBFi9RiO
SIzNG0JFjacS1u0VjbevxADr2ed75J2ZQotU/2rhnXBcnMl/Z/vMtQY5VAJNbJUj7ms7HlXV8WOp
cA3lI3tweTMzXiVG9xXp4txlSi1mWxQjPT+i9yko6URf07/FHPcsJCO1FauVK1PDodS0XxF2nysI
4aGYP7mTTSWRzg4FlCx5LNX5Jdl+xTpyotOLeTnLXKsTSWwSxbc1qmXg40aqj5RToZWjpDdxR6AB
glwgvJjDTY5xtISMjFP10aLn7ZHjBuKF3A8Cmbae/9HeQnd4EL3T31l/nAHkBCdoANEbxjgvS64e
WxyjYhrdzoYIGam7PdTSEvX+yqSr3EgaWo74DNc6rQuoEOzQvtHkss9Q3aFMoRLwRs/1DY/baqnw
LBD2d9XkNeQiURaDWL7xzXsxxoaPnwqT8ZsCVAlzCBL1esAqiGZSmjhKDadGB7mSF/EYK6CeSPoo
9UIVAQaB1ceUMc/ztAFyYhBPuc0CsjfKcrhZqZw3i9S1vFxzHaMlZ0QnxAR0lgf+ESzYfmNgUAJD
hKjeesJ362S3gJtxZ0g+8qVx85xdhoOdhGrutAzdjp+ENbt+HHz43QHHpRAAdGL9iTqzUKR2QJle
AvPfzxp4fPqR7sl3GAOQxu2XXlWMQE1rPWKDYqE84agk91MyXy807Sz6NGg0nyDY5fGuYRT41+G6
A3CRUS/tQPZ07QPl1qsgt/gICXZUAIk8gp8uj3tHCanX/H4kA9fzaQ3ZQyH6A8x8deRxlqlPH6d4
Ax26ZG1CNQC1ekmtq0CSOQMnL++DUK6MDIIG5c2M4MCfCL3M37cq4GgY1Nie8ztVcK6pPvk4bCAs
Nu+WV1ySOEox+6gBb0rdUOc+FnDqNJQ8SEDAZQFq7135O1mu1osN0+lN9v+v7v5WzA/kasDMwVwi
zKGqdmgRnU3BHzl85e6sT2VTC8ifLeXx8vQZd//pBhEGOsAW3FEQiHSFV5/xqs5PnYrhJ0dwmEVG
fwZ0Wc90vhDQQg9ZX4plr3a02DeVSd389K5M3j/hQNwyS0RrIimTZted3LH6qoPEHfSTaRfszy/1
Zu6YZoK8Fw4LNrEHbOsTArvEp83dlMYwHmnf12lRtovUt24FBeD8tEHPxVqcvf0bUwkDHFckVYDt
uiZsMimxINT5eiu4MG30XxNqo5tmSS6FOTG1Zqgfkh5u7wuBpoUJcfHcvMrsEV6fKzbAAZFs6n5h
bk40zB5dRWdbxkEoWp9H6b/c6JA03kD4QlLZyOCzF12FCQoi3DvCW7iwKDCI1aRn4iUsy4K7rpdq
2G4CZ0Ywuxkhjt76JSHEgn+KeFkbFEdWVvrEKmtrX+HMJwfZwGqgfdi8r71UPmIWU/b0D8H6eCYo
wtT2fASFKYUejDZTpIIRJtYgdfz/clO7gtR/dmzt+ZPsiTz1k/dkeCTrROgTYLLdXdOSiwL+hns9
KvWW/tw5K8cnzWXUQMxPF4PPvwKvPSu38CgZNiQXvXsTj9xGcbHlUY7y2nraFJz+NF9/P4bya2UB
KgHi59/j87ZzA3t/96BOsijeiW76fiq5mBDNuuxdfN0OaUIJt0XLW+FQZrgZJpfeHqkdMtoVVdYM
40zFJXSwo6ubrtryp0gmKDLydLSFXM6XjoGXzoWgSG+7753De3XR1qoCFRldZan2armiR3kWfD+c
u8WXCeyk82w7JpJDgGmppuwwrVrJtRuPWP5NI8q4bNt138MiOqqZYSw8rIw4F7U+Iqn0T1i+SB7r
d5CDKTKz/aOGr/DOO8eZMxs7gQQfmRSLjWDQLC3IjqWQfaZow/7UbJ8NQTmsI6JmRy4NPsS0MrXO
TGGA5y5NHzmpX+R5etkcIma73FShX6je/0aFgWrw8/3e15JwQDs7Xs7Exf7G8A3VO/g+ndG9sWfX
DdgijIcVzIVIsILQwEuKgNorBEM86hFzCWJe5tiiusMYJgcoUeaHGRlt6r+7MTXTa2i65Uisfkr6
X07hlgI/m4zJeZdnnQawACq1I2OKcUJ9y7DX/BIjk2HPEe1Nhpm/iNonkpqPZRKQiXjfvhemg+i4
jm5BGGiBzyz/PThtVdK1csL5yuNNsaYV8/5r9VrDDN7dzSLo2yJmT5frFTE0WpGkNO0Wg3WSPf/k
hol0JrBvhdv9nSz1BY+H31ps0OGvN8L3jUEUTGpeo0YZ9EnaWYirEsDkQ/M4pC4QqAAaCv54YGhU
EPJAMXOE9zv6zcQ7Vwtpb9SwRAI8RYqrkn/R0zp/IIAhwyEmTDOmj8+pJgQgn//VtqdFIa+UiKEd
0X1gb4n5lsfOi8zSpuzGWrK/TXW57qJwpDoDD6w7NIGkqWRG7bi6E/ScjBNmzbWob5RNVIHWoVsK
6T5o+Cjf7bmxEszMrMmMzIYn065p1wBgNQvKT80mGiV85z5SX5tZPMl7YGsfGn1RCjsKa8mUoC9j
DKH+T5DVt3PJyPzZ57JyxXCd5HLpkJxG+NgaAb5nGmDCkHv/Ly0ALxGP7ozZeQybHDQqtiWlW8Sr
qI6DFBH2wQ7cXbJukCHE0FcbMeoos/oVEw7BGL2x0fQykOqcQ0XNkE/K/rQSyuW+GJ/LG+o/OEQj
gZ6UMrRL/kBDZs/kZ83Ptg4d0c/lf2GHXo6ZKOfIiELbIqK7jEzXLVaSyfLI2ECfE/lzQc6+DVkl
KGuKydM7hsy4vzXwkCwJfCefgapAIW9QUfd2TAk7S2yITcR2NfiSUrEKKmhFEEQr/B1giobkkeex
um9z+ok4JvfwH7ORHxcgO5Ty07eknH1Z85rHLxhpXRvESeHHHBSBfaKxBc2fDwkfe2LSSkzDVt4g
OeNN9S0h5q1+FmX8hsDMjqm8xvJg9YwdClVwg8cjqUd0j2oLBiUN1UsEK8LzFyro8jtFdcHaFavv
rD+4dyN3Kk6b9Fke8lpR9GoCa/f5cxSg99jFzkoyEixok9mG0IFGcd0yUiQlADHS9CB/b85V+YDi
dWq7Iy2ZU2U805yD/loqSjz4JZC4Gfm12EofEoLVTbdqm5ufqPtzRn0DN612sQ00eLn1jnrKDPgv
0oOJHY4eOS1QMGRwfWSb5JEV1SyZ5vEN79EuuAKlJcbQfobLvdKNYSAK0smExe4nc2vt81TyqTo8
6ezRHHtRjYOsxJ9gbUpsSgcRRLp16RILDYwmDZn/m1fE01oVwLdKkSAo8DoJ3P2h8CtgEBUAIJ5+
FpQxQza71XRnER8gX8QqwjDRY7zDWcxVUn4anL6SbkCsce0Ge+82bl8z0KU37IS8TLb7DCRn6BeQ
FijwqiIA9umrr0uF8A9dQOjXEGl7SYGDzrNXs0z1QzP4nz5bfRVlOa60hsvslp8XM6LVO4Ydwbki
Ns6NusImza/0TEVaI94ZL/MFwr/bB9QvgiG5d3E1azWFA9aKje+RsDVLWC9q7xhYkPAXoXErrsEa
Yyi+hcxquLS+PLaf5FQHAw5m/qZyqW0VgwrPPJXmS5hqjlCq0DBdsaT4ny6UBdlqmUKq2lKivtDn
afnRJ+SiwlVZL6/hQq763vcVz89D+hHBUqmuroUpSMA3/mTutmRHfzjYtZmxmmvwqMq6x02wU6fO
voyQJ1oLpCuLYWd6BfWPAosyTb9LJ2SncMNvCVtx5AN5JeI7mVi9VzUYmjsHmL1fgaYA6yecBk0Z
z4wK5cIjrEoZns9/v7usqLSuzjWk4fcOOdmAhTerZ67fPRX0r8yT8PlBdH+ZoZLBl7so2YeAD6Ug
BIxDmISjdUsqQ1POoqYOH9dVxMX0NIsNakv7Sr//2up8bJ/KPPL8thv36IyK7bw3Jt9s8Gc75GGn
Jpxb1QuRJ2SEmiCc++Egry4Z/OGDTB5tAJyzVdEeYbMFKukCX1payhUj5xygK/7wyJx/a9c1me2h
990GX8BEKmy1Oa/vjXdZ4zhHLI76sjPt71GsDz20i/NhtdjNVvekotuED5BQWnSi1ulgP4gaCGQX
ucuWyWnqzlUpQiYhNAeY+4rn/nxIBBS7xXKPjeCur+RLOE6M1tsJzhWNrRwIolvNHkqeiEioLWf/
i0XUImM9sqFJRv/lpOB4jETRM3LFsiolSPZaZUmGcJKh/QT8ZDU/5xMuUeGLOn1u33QwNpc9W4DW
hRVVmlVrYJROJzm7M0JXltZXft/PF4B9ldtpbsEsQqcv7uTVsmw1oaVpMZhUITSEu/zw69Qa6CpC
RvYFioBOpDPjM9WrWvHsCmb0fndeSl1AkdUKawlMImY4aem0nJoxIqJpDptj9ga9hqMPlCij2dlC
EkgWIdcxBJ+FDG/ARjAUd9WZXVU4C4ixGTfmgKU0U32uuiOfuUU1123+y2QvlCQUFiwK7tR9YcuX
08RVnOyDpqh1AevW219z2Bh7uRPrry2aHAqLmS9HfZH9tFNJp5wRQ0L5qBm6sojMS/wFCO56fRCX
1A3VRM/IQBhvkNEtEjhRMWNX1vQ04EfW2YnpH+nsPjxZy/CwL5S8Vkfn7rEEtRZWD94GaeL0F1O7
jkTjNy1/Yq0jtWVzyPWc1xFeJmf15Ak93SlxaiJhGWQ/6FhTuJrrnB12j14cETeYKP1NAxIlw028
QyI8gLDNrpKeIt9rTfgEGOA61thdJFdtrAAf4L/q0R39SJ48xtnRIT/LAK3M0LMf+4VXQOFspGml
Z5/1cwH0uzYFy+h5Q6Pz16dQVHZ2RvOEKqTqk1aKgiTWb6r9LUW7ivlS7Ucziuo2OJJGD/J5Zkg5
bcjG74t2AlzYF03KMTnKiD24R8gmIicYsjAM2wqhrjuvOLo5TAYd3samI4TZVLqUgUGN+CglfLZe
KGKaO8DQDivbOR3Vn4PPPNt+8MckRYR7IuifPvNr6UHv5+Wc4eHU6snkscOvr4yn0mnly/sXXzGh
A/La/ktK+w8iWvVqh7FWPDDezujiR4eCPP/WU6NkXHIlKQ4EnB3tB2ACBR5EAY6qi+caAWBXy7gN
fL+1+RK/toJkNfk/qt8MlfaamcXPdHjifQix3bErHkDRKuo7b/zYVXFqBLL+ft9JRgeZoCYcDR/5
imbZG8FxYc9vMoqOdAxpYV3LQl75cuxEqI43mFPtmDuVbplf5zhnU+3EEK39qFAtj9Hfr/XggSQb
n5wllYpo4X/7UdTU9ND6FIe4M16YgupwL4ki2sBezHQr593p+4D17hRJHGpJRoifZWA3VAyVx/X+
VxoyeLjrBvlnyEGQCIP2ASA6REByq2nW1/BdsKwAEMAdq8YZvrKIiq/aFqcLAgDjGOB50teI1Uft
mpigbE3g883YKjXqfboW24chOgkIYsfTWKV4lOs50zqK/LKmMGo0VSy6lBu5LchlyyIEvuDmSn3V
AvYcKzNfn3ndc5Oxd6fzcZGsjnZCk3/110eJL8oIYZKXTcjMLtBRey3u9tQ1Tok3CdB4TOIroJf5
Z7vfzDnzE1hS4oh57JKJISocQqHFC29chazrxMYd/D/j6ht4do06JflMCVObhYuv1khFxaOFJT2Q
DXDH01mXuQLtOBtgT3um6PGpJ/kIT32ySUMWXApNhm7AGQSaPIfO5Rg8MWramWXX6TJ82Pq2Fhew
0xHixssJI1Yp9sY5B4S9SFWmRAdHf435OrzIMD/Q2NABHahMaqEGGLUTUFMRgavnQ38T5uQacoOf
uS1WGHOz7Sc1dwqT63TtrWAW/G759HaO5w6QPCiDXwE2WBrPi0HhK5hl1CvznwgwQfV2KT/5pR1Q
3QvvmYjvJmo8nS4zfNc/v6QwNHsZ6SocVjZ4bi6HRC96v2M8zpgULY2DyMn0CvyE7NpXuhIkAtrl
VSka3ynUUlFfrRJbzkDNVtxNOlZ256bDlyvY11qvMbYimz+QtZcwayk6Mv+b8FCXKpfX/0AddKxj
jkW9djHiM2jg1rMFk3l3C+UOlMQ7hHRpRpeb2UFIojU873eZ08c+o+TT6o6oD7qjj9rCAD05rW9p
orlArVxAH98ic4PUc7tVwB+vIteOdrmxzSijIGXo3p26I6s53qFhcn8rvehmFLXpg0MZagOFmR3T
TkeJqEBEYyujOyhknoJrNxT8k8Vc26o7t7P4U1a8f/yP9301Jk+whiaCd3bsiETXhRCReA7FqvXX
mqdNSi47eswMammVAczzsEoA56IJVhwdpb0T5YSICHKNNjkK59td8hExJ4djFyIYN9q0u+qrYJv2
d5yS6aQjaXrdTX8R9RB1p2Ax6/xU2fZtQjhxRxhz7/00U7WZ2KJwAfC8AyfU2APOe2OdMXxgXjFi
sSPvToYfzuCitfqBBUt/XG6zDaIV9LV+pJmLq6/hhNKYtYF7+6Yw03Qmzpu/UAsKbaOpZbtpXRBD
OtZAen5CKgXs4AwfoFMfYxexJoJerPfBCeXMtoAzcuwwiJ9LHar3YRxTfRWIwlWarMTzGetLICja
Isj9rowYlpoXoSlnA2oPis42Ds51HEeD05Fyapd5bh8Zwa0Ux+xhBzm7OYW/6af8QcKYrb4oHiKY
71VIJhBtJjhaJsEM8xjN2yCMx9CcaoD8UDbeuQQCxF+7SBg0yveAw/XYmHTGaOpm5INEa+Dlnp0s
W0ACe/fclqkr63CsSxtzqEkiuAaylrZxsYe19GCkuPFd2MriFFBV0LQjCFrGIfAOoRrXyn1KzXCz
XCYZWxss93YU5y2cFI5z8jBrVwTETX2M59JlwNRSU0FyPj8umssGNXavReB5PRqvSLyR4LmOIz7u
MtosnDTY+Mk2gUwbuJBNlqTj/pxgSOPIwuyGk1+VAZwiGqAiVKvMZReYNg4QCf1DG4vhvX1SECMj
klSJNCIiVlETjswSPgTD3fMtDYHL33u6uFx2CtQs+DoIRPiS85qdmd7V4UnNJhmed4Gwhx33n5OU
QYWG3DwIyaDtfHUKGCajUI8gkSz/WsI75agW0ibrautYADWR63aV8z9Z1z5CPjgcLZzpIe2Pa6ID
YxC+Xmv+yselgmWfZfNDwGCS51Di8wDDi9FTOVpO+Vha0K62ITdoTY4QIyylNr822BCVObAQANXC
6n5i1sghXCk8aHbsxKwtXwwYBfAxO0PQ7eDTM+wKCr49N7C9cncDeudaLQr7CaMt3rFwdVbqqx0+
AHze9SdBiOwB3bQvS53BDgQswOIv0i2M7boCrkRrHuwlJbVrvJ8yApZIg/w35czZMFT8lZk5JzuL
wzdrolIeeSN+xg0eBRxnxh+v17kkNfZZog4UR77YO4LtYKOjfzu+gR5u6senkA2rDCTBbbjJhAdS
8XHQz7sDHO8Po+KLCt/96JGQDloBO8+5ZfOHZoUQesGByXtj62wKwQ+sgBRESXX67ZKfXjYN5m1Y
4RGdM+gijbYqBtzcouFI4IEnsnak9xrPJxCO52CKjyMq6xPj0Mg/OZhdLkLUyAVoxcLT5Jop/oCh
E8onmzeFXFWMBPe24WmsxfNzYnz9lvQUkCoQUqFEE1YfuK1xQXtB6xsMbliGrjfP2qAwhERpPYa1
imW9jwBHaCnNTSTem7/a3vVcwricx2uAXQ4oNNGg7HIOKbqlgZGBB34sbETyndKngZywYcCv6lnU
iokOD3cvso2Y2eqpBAk7wFIW2Xh2bCNwWGxI2z93fJZBwC/vC5KauY3xjJM1uUDrLKCS9tZ3UOst
AgsBtkggmnyZQFsbs8Hx4EEE8buIFBhmLRP7bjN+gZ05Lbt68zKf633386t+sXggdP5cNCMBnan0
kfcXV8VjRm33jMpFCHBgyAnhkAfb41ZLGN6DBW+qiDPviy4gf9fWZ/F3qmzwC8/tmk3hUvJa6vsE
kTtqytUtbtXPQKuel3X9snk/gb6EtsOSNbvKgOtkIeXSIZo4VAWDp+/oT3a1Njasw2zpXnUM7suk
SKzj5Sl88RDu6GAyV4dc6lm4rsevTkSA66nlMmVxUqcaFvdNqzTenn8+ztUF/Wll214GJlm9O3NG
KYfflqmn/kfQKcUy4Eg5fhwZyHsrxWKwsJdeUj2IRrjWpq8kwF/hFLPt/6UKsD6jDqgQ5tIE4Gnz
lbPPWktXzCVmviA28/GHLcfec/+k4v+n0qhDgg1ispBojxMThz2aHHK1hbjbUK+YX5WRK/SlZAOk
ZtVtZK1RL6p3GwVxY/KOQrC65k7OXAEkHjvvO7LlrYPRtjwMjQZkjTrgl/IzH7LAswgTNGD8Ta1c
g7Jmoyi2tSjTRVtbI5YmW0lpsxk99c8+rCj0uQA3RKrzbA41y6rW0l/+F1AywTTTbuEJvIUo58ez
ksPyqBGjzHKqhl5mlcaymj9mqLgHNdh/cOk7yAjc0Id9OkqWNlG4M8wooV4nfv05KbDo6l/YaAMN
5VxmptEvc+cytypaiwtLtaSTockNb3hmKN4nj3It41cedKFO0C4MenKDaXDUz4MRw18izOLoW6XU
B+B3PcCQblCv0vyOoSeyyShH8k38O1zOZl8HOaj8SsQUDm9e6eMrlAYGvpjUSA3NxCv7OD0axG/c
S+DwR0XERCVIPTZ7wNDuyy3jng9i+ESZC1dwe5W9t88mO/4KQrkm2u5+Wn3YWDOqB7/OC47uCtRQ
pdYbwiDr6pnVcOEFKeJKe6FrYvPkK+YPEPl5fJtyjxb3cUUa6s/VCDT3cDAJODZnyAKJ0ouk9b3H
2SH9+MLVSzpIMimNQnhCgsIjRUQItbDjOFsqohpSDWujUJ+ZHS6YdswUoYc33T1GdhHXl4gje8ln
2WbN6pqyZ8/ZO6/6/XUqjZrMHKd5G7RYdZk+hUk5VZ0XaZmwULF6EiCwujAqdgHTRw49WroJjDdc
HCwOlI2fn+echIwmTO3qcqK1QxOz1J4ssADPcmKtOhStApnULyl0yt7325ERVFKYI8OYl6CvcwzO
T/zDVAyhtOqPM0Amrs0g/oYQZtufdOKEwTrHzEBsgaX5aY6Y4LIYRw3jtW7X3aHfC4/mLmjNaqfl
DEyDihfojTIa++ZSnrJkQjK6I5B7HCkQYqb1Lavlrgo6BbsfuRLkzio3iqsENBSD66+zUs8/52WM
JDi6rMAQOf1epQG8wltgoAokOpaPI81biTooO/PafYIqRzHAZgx0OFlv5nvlCd9NDKPdARUrY3xV
19T80RhSau76//z5qriRct0bVoLe4VVZ+e0EFA6dQ3fl440MHilq7zM62Nol3JFTNWxFsuFqLy5s
Kg6aAFLFrJ9bvGfHAjQVrYIEGw7CufQNlrDt57cwmMVbYJ9IqbIW2mxINpQxAfHtTbLNxkK0APug
v5RKUZqv/k7xsly9jyyRY2oOC3VG8gyMGhnS4lN4KbNH4BJ+T4eAJRdi3LCWl7O7+seRgSwEroAI
1/MiptX/BGHZ5SJS4mDsiNbfocc5xaEAZa3rmCn0L0mRBAAVNVpHTb81Ih5AY+EGJ/io4sjOEUuP
xlfdP/J9U7pUDXRgwqwCWkYsWrtDXakD7yt7HbpGj0sp+GIPkzDjiwuJLxAr44mwkZbR+cS39um5
wISEsZeU2vC2Gnu41HlxKldfIFsqVGMIe0n81w7JbA0yD58V4aWTFUhItDtBjAGK9xl0rY3FhKWM
5jkBEQk59c3Km92HRzB+Lke+IlxW6koAP8CIbGXju4BYt72aUuiLx8f0cRndBiu4KWZl5V15pCn5
GA68DMFirgni4ScuKpNaITNCZu4M5yRg4IwOid5whkHzTV+G8pN+TtJMFPk8QRL9KlhDPAgZizL9
9xT+NiISNQQ8J0oWhRvuv8nJd3aa0TOt+xlNHeHJvTvIQP1hXHLoLzIfyKbytjUAasdp99SvrOlP
CDhJAO5FoFYRL1waiCaSL0xIB4XJLPHEiik80Ymz8lEX/U03IIw+fJrounW1oK/RNs26w2uV7bMq
bmaUNqENNQ8zwyVSuOzHx2LwJh32hIuo9w924/stkiOOGh/cHPc6KnFdzVkny+O1U8Fn/VjiSxtz
NvR5bn606WRxxMrWip2xHC42woyEaJuVL9hNz1MWzpG/LYCdY+X2Xr/Ahva6wZ4fmZaG8E/of/uf
m7J44odg5Z3+/hTozB0quDA1JuQUWJUXa/vdQrA6s0Dyt7aLxJidaxoYCmEGsv7OOqtXCmXasV4U
SrqxflEaj+LpGhQE84bqd6vEGqy7dNgdvhDXFuLpfCEyNf/1vvlLjpFNws67xU1YcpP/N5ZFM2uE
8gRHyDFBIUk96mkxkUJumHfkMhq3Sbp1wGJJZTclMQydxgmieEKuNT4pg6n1I3Jir2tymr665HNX
k9Uh7SJid6N2LhdY++TxtoRIzEgEFszOs4wB0nDrs2YD3PQVbOoFaDMBw/TIjgtL6ZMOWs0nA1Jn
S0K7xOag1/oE4Y0Zk+YkW39quQntitTqJunDXODRhM0ju25zwjv0xu3HpYxl1zFBzTsRHaKPkXuu
kUxiyICJUYz2TydiW8JgHmHJ/HNgKLiXaxZLF+vCkRyPDJJWHUkMGLtdj65cGN0pCjOEzNHFIQI0
r39APNeEwAaSY4mbX6rQF+NXrK4eNQqePOMskOvLzGD5PDEvQWKjcY9KbhtmdPU3xkQqqLqd6j3g
CxKVvLWkU57Gab7oggF4zxD1qB+kRaKVTcjNHmEvOaRMvoJwYVlG5lbpYQHmnSlxDa/4kL9dKLnk
6CwFoWDH2tgFTXjhcFV1xcZV8mPQ25LxI9cFgLrko3Y/Ytu/Hv+KUuGSpRNN+vLLtArc+ExQ1yoB
m5ZcTiniuJB5328C9YOL3XhBlnuXdsfT6IUaP9sYwFnP+te7V311vIDs5YD3OSk12HqNoYucoPIb
bQ6Unb9/GmcdvAB5pabCwYpFbLFWp2xVayuXIpjqpgu46SpdL7TFZoBw8g2QRIjIggXn0i/F4VNO
zVDRf4WJnvUvn4jXsw+52NrVnSqDf2dHg7Vf3WPTzd1ZpgxuchmCsent56DmkMgXGs8Xr2/EPtTI
RQj6+mLqiGK8GCMSFQ+eag4HPxF+7nQhZVhe0WcuZQ4ivlvvuHWZFmYBR77lPJAEX5hPnUVyf0Vb
2nX3TAxdh3L2RQRP6wU2ynbR/KgoQ2/hW+j8gXTdrfZQsPxQrd6ddGohlzpHF9n9ReqCPbdxDpZF
aX3ry8DX6sOBbguePPx6M7KMmJsp3fW4RHUv6qQtR+Ac7XdaxWvjsk/ZhPJqsFwKoeJ+KN4kf9kK
JhPTXEc1wSgTlZmwS7hf34Wf4KrsKxjfOwcxah9JlwX1GfV8OdAr93Vvw5q/M4f8V4nRzeFOznkQ
47Lrl+0BLW+jsyLbCmhwtR2rEoD4APfA8PbVCC03Ud2rm6DH9HH586RXjS0mdZo4GVgIDmwkYQBp
7zTUJbszdbv4MROP1AQOnJBdo1xotkG3Sos2DPAdomP/FCS7HpH8dF3TyPlxr0Xt2GgQOhKvov8D
ajrrOirU0ibQWmb6c/VxcRGP/WC48/S6hdig0u4knNrirAWVaIWKrTiZeqoPVqzM0QE3iYy8kfa8
OknHn7j50F+nEeGJfalJwQvKoz64pdniFhkis9ctzZ0naiho/OKGjRsAcltbu/ANQxEroEnf8f4Q
T0oGS88IIonC+n4RO5fuMIInY7+VTMCcgwiB3Z2KPxn/1/dogeKiTkWtL27UupY8ek3E+5tlNi/l
fvtS5FFSpO9s9MwfGt7IHpsteaOX1Lgi7ekJ0UMTjrjxTsCEron1mNswxonhMA4UCKUXZia+ZRMA
TE84fN57fFIHrJ0LoBfrAPpm5e4IBumCtasblZESBtWu+ih36hynfQZGeBWskhxmYVJ4hlKdRXQn
+MKqEecHbdLWjqxzYNIBU0Y2wngTFr1lIWecguIO23cjndCLeW0Jp0gBxY0BIuB6IIvpnNoDBYPx
JOkxTTPK+5esbU/jA3X/UBCGvfJy/eSR79fc0F/AZAa+algHuKxRmuo5e2/Lv/wbtd3zjHrdc4WO
9MEdy7I5nC7OPnvr0CmFQsU9gUzFb7l8mfN+z99koN2LyQyylrqE08ZO2wQ7ASTDZGoHoKt0l5rK
M6vhwjDiu8YBohvBR8UynJFSElWWxiFeOCiQm2DNxLsMLcJUeCgFULZ6WlQX7twPwBmcXHFkWfKe
luLsLB2zkUh7rA6kLeTjpHioEqE78MaJw6G944mqApM32FpoWuRZCLj56LqB302NFrJ3CiX1Livi
BaVEGKvdukCMPTpPK5nDnOOjTLuug4FqiqbL5bwBz2HwCKmd8JgXti9r4pwLsVYGtr6ByROivuxx
MS1Yums40e5fWBxfSVf6JY7hn5CMnOKEchpe08+MjXBTOEdndvmjC7AFC+6KGju3Wa/6C9IQmSph
VzM2JzOMS21CPkYwPPjDmn2GRLfJs70qndIDh3OcU6jNCxEiNDBeYzijM5KIQRn/uJ3nusszD3AG
GpcHOP5Guusm1KNNajpAtiCtlhXtaZeuCmfqwHGM9d4tJ1OqIhny20OP7gDWcs8nwz+3I03gSV47
zj1MiNtZHLHS7aTMonjr0UFg5U0gbLaMFydNFQV4aQhhnGWwrLT402zZ/n/jzJcQz7UPj7+/z60n
DxfAaDnFH9EFFpSx6pF+jJeA1TePP53NkdYuXBQ+7RwqemrkMz6pQHAZqNjZiBW4f6xL5zDNNL7Z
/q+BbZMcN4nzC4RU245NV6Evehl8hv0FfSj7sI1RjPRRD7Vjjwl7H80u1B1RBPIvO3w4Yh8+mpLp
dichODmLT3KGE+DU/KENUoBRxwaCyEWlavhNXjffS92cERkT4Ezz2Ysj/QqTW586JoxB0FIeko3y
ul8P7EYvGxsqOP95CSEH98IstWHwRcpVr6KLS/U3+CWT+lU0FvvmpvTxflKCN1anhpzOnYTARdmQ
b4piZDmAxyMtBOekeHtr760s9Q/uAxYoOcgQEcmHpK46uNZ0S4Hd561rhbA63go2I/4mq9bbvwMM
KzkdcDnpzS0QhkckV2XIRWomJAnrf3Zqy0wqidp1aPOAOy2UeLf8B7VVWdMZgyOGSPAO1ydVSWwM
TElNl+Pbfsw3vGt/xMO6eAjqU2ujzVMBb5vVpOH9ugMYS6EpOigApBCIBbU1ENe8PQdU8kG+uLcI
IIXk0Nh2F6fgkm9sW6aQU1tYaQF5Uin7XpsV7jkTknl3LqThOFHdmXFgd1gbOzDoWsaqr05kqnS3
ZViFbTv5HzCRETZbIVvJXSgBW58o0JgHvoDLkny+qbfBh4cHI/4WoqMyvEFi8z/ODygUIw1pVDP/
fLPe+f9Ew2Gs/S2XbI3mWQPDjGozWha7/eKx74yU5BEDDLQWCsgBbTKtwB3EYTDpTS66bxjeS1BM
a8/aMPRzINDt2bpcnfAeGKRZ6xqgpGOUQikByseqvWK/9SxS437pVAXhlEAKW/xxWzT48Ygp0OkP
J5YfuR4q4inCsbCReVGIdkW0nHzcvVnxWy3tV1WmTNQ8wFC17ZY5Cn1D2emNEKFNWs5L7OwBJDTT
UT54feqdR0HOgRe8EOWUn8ZFgW7u5U+3RqNTU4jgwKKrJS/FXSuGzO4axlZ/5G5pDWlYxpwb0wMg
MG8lbUbvDMcLmVYldafEX5I4O//95EnVpYdqE1xwaR/t0RcSN1SxaRlMXhiTxQ1fCs4x0NtifAAq
JjGG7EfgNlpj4WJVVqiGkHEW7Tnj8qTtaHObnsdW5S0dZ1dsPJ4DKswQIib5g363Vn949p384K53
PeHAwVEVYRfXVIJ4SNwQNa+m8x4/TB4flak/cDFqBiixJsXjoi/upObRapb4/Z8dgwRWGNk6q/I2
UnRPLmeJdzQvIemgj+oEwT9N0iIz2j6NJdRf2qK7SIZuL+87xZxAV+zRjuXCIO5k+w5CfReQx2Ow
zONbWyvhR1DCquciz00TCEvjk0N5GpStMoYNOaGh+vI6R1k2jarWAIiwIhUUsZaibJ+9CZvjj8Ju
tt2pcCvM4swTDjvwMp3cX6eNIYSZ4EV26N59tQoKJPYgh2fjq1YBNYqBaLtv5KHrEINlfa7xS02L
HvCxzYko/KlGyhyIO88h42u6sCqbXo1ETbjAfQeQqsS6b/3b2k/zvWpJdL/XeSmv6TL2KDT0BCob
/TTBYu3POMLjPa9TvmISVXxAhBL7gEDSey5WfIffUOfC5kttoVDvmdCPSk1yDGx/17dH6brKaUdJ
k5IvbDzcuWFe+5ZowNPu4CZ6z5Fcu+RgQCJgWUNRITwL+lRmnZJ2rH9h0hRBpy23ERXp2jPbCpjK
VXDHhsnEgOKfVMgN/r+y3se5qkg1TDW5RxwfrWf2LNjNqlB+8YDnJkR4ZVEI9r9SpcihNlls8zu9
/3w6b0J2zz8f7ZCvFvrcL4GGZmx8BZAbDSujsveopBJ+BFOrLT3EfoxnBxpGkvWGr89786JI/tGD
HdGcTUtpVMGZIshOaSkgIC7mIcgSDfbd+p2gdB5etnlfl/lhg7MQhL3rzW/K1G/5XJgTByZn6554
yQMd3MDuiek6wzoMhsxB5kjmk9t8qxWMkakq1THLzQxE04wuGEpM/OKSC8YXtjGy6iGREzQyHYoA
VXQN4Z5qnCmquBpZrq4xOTjs2B5cEL6CRQj+zzPR1+xYIs78ZmpIbxgnVHNthhNeojIagiAAHK+o
rTH2m6V7OAkdCCnaMi82Mb6KzOnpMit2UgTUl8tzqq65hLZ2qg87tYX6TFpSuE5tG+GpYsBQu9te
v6OGGmgLmAeg2G9vTA3icQxZqBzat++DReUM1hV6hu1p76ZkTJVFuJ4UZ0fjL/lBLr7eeixDH+v7
uvdFP6As4lYYc7mFWONK8XR+c9sR8HqoeKEOa6UA6+Gk0AByH2EJnuIbt/Mat6rOut9cb/U4RMLq
wdLiua7RtsfZ8QldngDqLjnb91MxYaFlTD9y5SxprHdK/izptBsVHnmZsxeL4MIOpOrvDYSyuW0P
wTeZj886Eyl/bhIUuJZguK9LLu4SPdHy+3Tgg/6EndkSrk548YD2/P+tDDwc6sBj+7SfuYOYjKz2
WX8JnSA+p5g8QhSMnVgfKzTPuhX+sbsTUiVx5oS00QVq7Ahcy7UVFVmXJvtYGY/BoxAODUEZ+HXv
NZNgL2lSWfFVzmUbx7gpJFTjHYO9tDhGT9D6Lnj4gubQEcYHq9laBWThd4U2AnbLqiKr3UxWnC5E
FhOWLoARHY5Dp5fOaJC9HTCBra7jkKM7cGxFLTNSjjfTLLNa+cKpMaD8PYPaeAxYkvUTpZ1JARyQ
ByNNoZgzRqfNogj9MWZ91W8oWNibNH/5N/K0vcB66wPJNFTJb7w4+0wKU1qV6dUkKEpQPGzDS7u9
391q4Fm0O2BkoHvovNnLOr5ucQvcuLf7DXh3YctBRlwf9kaam2JsBKHizX+N/oTktDsDpdYICIPN
UYg9xBIWzRIX8HNYJzeVjeS/KK+vwJyQ5eDjXgiLacg5uoiWIoeilYsEo7cHdUI5C3krxGpV4BET
VJEO7eqrT6rqTkTJKIO4987xmoz0uIW3RecALOf+ItBsi/baBSo6va/EnT2Qlr6oru1QHLGQn+OU
0Y5kgyQ4RKtBNc6BOKP5aIQyRnLcaRwqPGHHqt5SH3YLdnJlXhTK804KZ+Bp9qfJTQz980si/BCk
OlZ5FeR3KP/S6VAJhL8TS/OlVvbGthVlbxs+wuHR+g6Qck+MLKPRGxttQ/ySRe4sgoYPoOorPtao
TCjFgSKF0sUY2Zhh5WKz2r4tuLZ18jboaecLznwyj+bOr/+hLHm2XUH3Ra73Sfs2vLvaKPaLLRPF
kCFX5TirBjw1dGHLhsGVRKjIJoc6i2M+aTrAxiicFRUuRtKBTNavRyqHWBixovLRhbfyM6u48Fr3
XpY1Xuxwhd+MZh/Uav0KLwIelJ4Dm/1D7YW3JV/LchSYBfhVjqOzv6mLjgJCO4aTYYyeT2DmR+z8
lXL6c6EaALf9BoTO1hGMTCXOnn2aJoQyAECBkEMfOFTTj/cFgX5KOWde1FEyVsl0x5WOJNQGhJlM
cv8bGT5MafAkcwzUaCFeVDqtfXuwORKq0G5tsHsYDwmsTSWPWtIwQikPLBITR5KQ0DyEKUCbCYDI
iRvPLFXb1qfB8pcDkuaCUade2In0vl1q1c9IiwkhgGUvZyGiVBcXUocOxCcaM9GrggqQlMaDetGy
BmEgC9UDp+nMc2LltP6n5hvPCs+N5AvkQmfD9K8EkUlUAc4oZ41ZmUFg+t7Tk4no+7/lg/c1D2l3
LMbkar30AOoAWu5yUAWs06tDS3Dsa5lEsU/tLLxG2suMZ0ch1ElqBGyIjSbCfremaXpUrQomgJcy
yz2PL7lHPmRO4MO4n+LPea9/+DSf00e2BnQJlRY5+hbWiI/3QFl6Z8pvPG/oE5l+HDo2IWpRmvsQ
A9CYxkmyBK3N+YcCGTsC
`protect end_protected

