

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MPaacDM0TWg8wcifAVW4jEGylx4PKrqc4CLboKEk0r6t7KyfUnirQwQAphZDsR83L059CNEzB4wD
M8AKmBfOkw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XUT3zAfEi3anHP5UZ9Q64SRw1RnMtcFX7nJsXqsc+jcNnlmbg5PdhmwV7UaFs/PrWKFdgim7UZCy
o9NtHbXd3iHyUEXXZiWfkC6NC5Dndoi/rfKSxw5AtxtcCSaJ3/cb/i40IG38fEOD0mldCmJ0WOZD
xOW9J2aHwV12uWmmUBs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5hB2z6qFvCHrfde+xOJHAAm9Y4Zd5X0rYu4ngUzTSYyHrr6WAc0PuLxe2Zog3gNAv7DFoV1y/Y4U
F6T4flnTjzAqIUvyAW8+maZzCAeWDi8VgmeKHRbLydt/JWB9Ri7GcOoofnS5/hxq8wRCMMkoHbQF
kNzxfXz2j2QXU8RR6+E7pvqcJkK5H/P2HIhS88SnGwppr+eD2lVT18h0s/QB43BH12kpY1JIkQU4
LOR3Ej9QoPTxmx24xAodMjc6qGME333306vLcWETw7evLQ7fHCoyGS8qVr9xvwEOuA+HtAnx7p26
Z/azE34tKzoImCmpb36r638Bv/NLBk+b7agF9w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n2iw7CqdgxuZ5kdEH+pm9NjU5keAcvOSKkOt8pim3KzIVtdYby3hWhnEsC/F1aUQ3kkgfoeHTv/o
nwfMP+AVXxDoH7hATDu0iX0A8s8avaGhFp6novk5xXzwMVnGP5Rbk3GwwADpRNWqzKN80je+JhyS
o3J4z9hQTmce/KBAfWo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sR/mTVuOveJs41YLuqwkxNe6mc/KV56Pt/6c0cIYmcRhmwLHOU3+/VfoPpEClea5ISswKcgmSmEA
91cZp5XMe9E1MxpJldN5YBxK+3XVJrpKIG8b4LM2yC+ZTp/81AZ6CpAKQXOcZAota3bpWOVB7WQt
kPn3pALJ48nc4gaIOk2j5GO0g6BLITkCLwe8Z4XOzYZAEaEB+5dJ58Q/7AbNKHr5UdGO2UVVG5Oo
7GIt9ETizL/sKscnCI3CshbxwDQPtnh9/CAQY2Ci2Oqc2ptOmylUrV0jpazJ/ulKvyLMe7D7sjb1
BOUUkYAI7NZU4AkYW+pW9jcllm96HEkuSjkTDQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50560)
`protect data_block
Jo3Fe6MnG4lufZqpjyVY+elXGrXJiuZpv1Gma1KEDdzoaQdpV+Rq0BNnHpbuq6PPrjpYGmHPBlkU
VrEc/Qfc2Ib2GnhAhRewHBKE8IRp5OkzHrdjHzIUaycoKgHIyVYmVT48vxkHwddg6l4pNDqERyDg
LqcQ503d++/vYkNZIi013w1r+U1kROmyYgJOHKb9L6Q40bvC5Vv9YT3yy/ducdrPgqu0PqTztnhK
NaVOu7ADeoiEXHRJMAaq/kVfzm0rA60YyChHu08qdTD3LKc2jhEZZYNjz1JGfKGYORK8+6Jah4o9
m/4VeHvCCTxsXGqmEkNQHzLKEY4S/FiDsJi21AoVxDxbTI8nqWi1WQ9pEZaJNDY6brX0QQuIR9cR
k/7jrBbOA9Qav1okntTfUaxgvW6e2MCCP9J7865beXV8wJRHPo9io8n9JvAfWvOhovcqngb/TOwC
L/LdaP21ionpsFm6Sp6h1F/HdgZDmhb2NKqNKS+uG3PDr/uuoQI3aQACQbyGIzcPHTGhtxTCytyV
peMB7QH7jDY1eICcP6Rop68HRBJFy+q/nEcWbKITh9ys5Qk5yp/CTeaNsYfsm8kDd0XNC8BdTmnV
uAWggx37fJAcFIoXJOuSdLP9+5L2Zb9seTXyc7Ty+jXIm/gsJeLi0jaiMoi8ENHqJlUOaG0jYI+m
YsKohpgHBnvxb1MobqgU2maW2bFAixfpxajL1ifch3zlAfeS70eXKaGpPcpGSgxDFCM1lA7t+7F1
tYO23FMgFsFs0715HmENRZaXA1T3pI113dkXI4WZm/Dke6wwKltfETlKd2Xp88sEE9+/U2RI8pmY
pfW3fGt4815hV+Snm6NzM0+13fPeEojHJ7jcvxcqFeDgsWN0UW0CsLfBglwPzCJ7jd0sr7QlnaoG
aVjTQRsY++PYx+xzJ/xTM0Nyi4DBK1joReMFlLxQwL+eCrnjbVEkPCQNrcS+KyZ1Obu3XrOCo0sv
1l7NYJlFhVdDYfLkKWTuIMAvK4GGsaTlCpuDksGxRgZYtKWTi2oOm6R4mm2NTukejnot2rc6XH1U
RUlO7TBg/tC+AwUAFMdIWIMIaxz9iNOeNIu83FuoBJ26BVy8HKFKQ+nvZZG+LF/FCV8OyBAIuHdy
9Ba2Aep+8s551J8iiiDa3PuO4t3NFmX4LXOnkYJe+wQVEAeUcFPTN8noFbzRU2siTsQHRPfg36bt
5fuq42ReWAIlG7PPBoz0zSSwfUyt+Duh4J4aC8Rkmc0gVsFpBLX1CgpIgWSGGFG9/xLvURcgPaOU
GA/mgBwsKjL6D3fylhHsC4erklr6/CL/HAj+TPojUoRcK2/Q2TgyPukZCpQ2vgmE0V+Zoc3CLEeN
Z6OapJ6LoGD+FtA8fcfc9u8p5PFes7zQjmvF9koAG/XBso5RvrZabCfXZfshsDugyfP9Dm3fCm2e
8hpZCxCw/gE1mk7jSzqjYvdtBJX+ebCchW2p1SZrS7/r/deh7u18bJGYwrBP0udYWnPFB+47lyVh
7jAqFi0xOKCs38yZNLQebT8z5dm9bqtXNQrGsVTwv6wnECh7QJjzhvHssa4Lnps0fjEGBdh7RVHj
mEPUFHtImIwdGilmtRZEnDwx/erZXza+0i/ghGrlGN0kLgtXMyiM7nsJeAH2O3APoPFPoFjMEEYe
olBdYt579KkKN+OK4swjNHx0Sy/VCaulTfYAYyMBtOMPKvguUgt9slvritsBYNebcCDUrN7zISE8
3cJj7Pfj1a09J9jSqimbi3hcLy41jcah/X2zodbGRetB323QEaMJ4Bjsheq9h6C1aZZzRT+nGxT2
gXha0rhwJEmewV4f4ouO0N2+wSjEl62QY7eT9DP+SObNmGH9i2v0UiA99PD9Xzi5i9N/GYmJjT9V
USOuulGizihH8v4DFKBQBcUDuJvUj7AKYFdmTzIitreZCO4WOHWmJHXATwyNUb7Ewi90lzUYWB8o
4omkqM7DgMaL48ucDjJuxsrvcKL1egtNfHN+mGRZoZ4DI6RQzZdz6gkcvnrIwlyXDYMykj4LCjni
ziMeDpm7NOVHe1b63Ozm3v8safamN8gu1vXGHCBx/QcTEIXWhIRA5bXR7jdbwJksDVGJhle4LUO2
o71D1H4RIc7TzkD1XDTnLHgVrb+Qd0TIn+o6WhmkW0TMzTPyTzLNin0VX9ZUAMS6MhI/P+4s/1wD
yTOZqi1YiUppQ3FI7MTBfOh8tw5WyklqVzwNT+khyyKgGUQ93lYVLqLohjlpFyyeZHIZPEieAbaV
cBBEupnRClZpMDlycMulodoj7c6GJ1IEAr/4eB0amxTKhdzYYRae09RmDLPtrkvs/JQT1btV5hu0
ORGUx2IctZMVcmN7sSyKs71zF61HflmnZOZ6NwPx+q8PxT0SngWPj68gqujmFmA4lDKcY5wq1CqF
17Zeajb7YsxQ9VvrwcNmz+KtTDHyqDtwmuYbje6cl0pIKIDYjg8Pi59H1OXt6mxvvg64WzoHPqAD
CWC4gdMR0YAfdMZzslL6FtyNjVIoKLDvN39BDND9MFt6IQtm2pi87H8BkhoXyzsshJgqcShRGzQ8
JbEWenBRhLlCLqvAve9YXgdUdwmJCz3eUQEtT9sRIAqUC2Ge2aVMk6/9ftZygy7JZ5XZ44wKSD49
WuFrfEzoDU422CrAz2fuWliqCyaMejJANSUQIwYDZawhuVaZnO+1RmCduWhlH3hFSlZyURjMh/lQ
PkDJSanuzYTOS5LMkKFW5bHZNOn/zAYakz9Tjj5Ad0Q4hLs1QQCXg6witAD+InT6bzGhh5UYc2D+
/Hh2kDRiJNOhr1APTfVROWnktgsQiJ78iZPf0pe8a053I5ZluL9lMg0XI05aDxrbJlvJtsTSP2B4
MFgK8EVyYtnASv39aUnxGCYLwKf9wk/kuFDAu8pb4Pwnu+PEvCz3sWefAB0SdOwaxZkkHDt5IJTy
Mjn1trR0zfjiHx9ORU/eviiQvhOqSmIQrYN7O/gFHIFrRqNnrpbTfc7CbWi2Ca4nibwjcT8P+dSW
pdegiE+RmAILtKNcwZk85BU3SdnPgdJpT7c+7K19/4M1iqHolFshdikJRSSgCi/mwAWYJtUhG055
a029BqpgdTlmAIpU/ZwbFFdtNf/BAdTqumUmbmR2OWCuPfOkjBmPe+0Og2OCvEIlV2ZAs1iQilu/
liNXxX6qAI89dhLLY43LJG9qDB/JTp8ElUJ2aToKL9/xGUznsV7kk7QpPhQ4pu+orVAL/Akyvs7f
xVhJ8lbFTaf0dnl/LcP7tUBnI68XMyVOpR2TDeCIcbU0ZjtpsTpEeZ/e/j/nz1dwzL4jArhEIPXg
3ud3Z4Xwsn9cvOdp3QHxYp+hpKaF9jK8KK2fkwRHrVXY4vJarzS4v7lnMP9N6L5KyfXh59RBlbnG
KBbrhcBAxF4Tv1LHutRGxxX/DHDxyYR5xHp/BiHGDZYc0QG/ren4tt3w8b2nYPqnDCjmtD3+A/ve
UU8Wjp6bylop4gOhnxnVCv2he0H2r09hz08MltfA9AoUzNMjlsiwoXsLhHCur0NofJCrm5VH2E7l
i/MalHLBLNaMlQ/pwVMEi75TPh0u8qRVksfYd3CX0X6JCgdU9+2ZzBdjP1Uw8oHBxva1me7xJ022
cKaMPZG946vZFGWAx0jEZIAwGGYguud9F7RMDj3QFyLoQsJREo2Y/GQCHdRjdjd0oyI8ivVlSHLm
86kXy2pRerfe+5c1xZjDPvTbm1X1J7KlXvZRlcGrKNWT2LCYqmRU29spOmsh2kki22N6GIe8IWiL
ZoofPNyfD4PLFpaPHnyvub0vtuKBxJRVpA89Y28vTCH7DxBqYTLRYAYCz3Pf6fTivcQyItWXIWuZ
r54p/MU3GASvc9IN+JikOTOASnQBO2xFvH8SehyQlqlHJEwzw9NTcmo+E0lpIuq3v1qb3xvQ5W2O
CRYJUKlqv0EHVrlBhAwEFApE+yGmkEOgV7vQOvO97UUa2mMkamnz6nYKRbjwte7w75xihNOeZqRM
VIlfyM7LdJx8J9V8MSERpKh78hyci/on4okUTFJibXNMxeFzNUgDi8PdgZwZDwKFXbbTLKbCncL4
CnAtuBwVngg7ezHHXGWAnpmzT55hKhl2hPQ+nPVx7OnA6WOK4LRhkhLY1i8BgKN/gCrY3ulBPAMu
ltewEkg2B/OTq0NvQxcToh0UkZJykHXTsrtseDWIDPfO1ZTHFwoyVO5rW2qcpflP7MRPwfD+Oeg/
mzwxDrrOgtWTUnmAqK4Q9IMp7thLLht4taV/CW3fdPqAmCCfPw5sfgw8VVV0rmqqrPOTXTzUV+Y/
ouvkfb8T5yUykyKEntRMKILEroFoUf0ZuiFg75z7OdlVbIEQ1A4M+pczt7zX+gzgbW8zUt10gXvg
Qd/K6Z0FVmDF7PrQD7Q7HaiYqLh6IHRYujplOzry9FNM56oDZjwBzGc3tTtQFyTi7VtB2ke+t+NY
drnWp/v/iDs2kW6r7ux6YJ5bqys9+iKDfw7DldFclLgS3autEvuYDSaR2mQ/udHpODmL1v5QNSil
2KCZglfN/+gh1XCY5BMr8PM9y4Cyp8VGT7qg7g69rVoWEsshnPEEy2G2h27ePlbJAfn1bf0tDUV3
nL0FrUSGiYVc652AD1ZyI0Siaw25mV9Nbdm8TN/gqJNe1QYPWh8Mi0x0ucdvK0tDO289NU6ociuk
TdmYvrrNlu3z8u5s7vvaZ7pWV/ZPPesbD4aoz71+UAJjF/OnBi3x6keZGk0sFsOsdEeJ60v75WcU
osQakdWO+aFG+t6VFAgtcLFbcaCAJYiPeKd3SO48mEh1t70EOIUcIzmDZfixyWCy5H0LqPE26i2w
IxaA/H67DfQAwn/Y4Gto5kn3YcyzlAETQ6YZSxZscBshifvppeek5l5QTioqXv761N2KjjdlHeUA
/QsXEWa7gI2c3E3IqOdOgeA7be8ikWIQLodnr40ZVI7/nkJtDj17mZ6mBOy5HfMXuYKgjOKukbOo
yg3oxLqIsAlJMEcYi4yXRiFVQQAIqqOwrdDd9vp1c/A7u2eXVH9dgY4t84X1CkLmQ2VJr5LxeX12
CKQjWXrcAr7qfdn9/c4W5AYfVEnjeYvL77x4qnM/n1ao13gSz1VBfehGYfF01FmQOyfazPbSqCsX
CSRMsGJN5HLd+BcLm3DiI4sJsTkZ4y7vs7Kwtszq+ri34Mmy2P/HwSPtBra8YGJUBcCH39fbXA9E
/mu36JhtKPJ2MQ955MhfRWYeznTFXHHXfgy90ICfcA/j9LdZy10mD68/dxa+YIVUf9vCmA5Jrba1
qwWEI2PpIAA8/pQeKTUE3RqSnmSU3zczDT0CTG8gvtpg8ca36UUcmnRj42yL1x0TJ7PtPWfZFuY+
JPWKbafy1oGXX/ye0Y1NMo/tK49hhjii3LrY2wwoFku3QUotC73q+/r3cdxaPtVoyOunRJV26maH
FBbZKfx58y2PAtk6N1Of7bDdwkdH3VmUYQZfAUe9oSjw/MkrZhRyaWFBAQsj6GwZbBp0kiFSQ9YM
5HoJdo2j/U1eet9UsNfSEro73AqN0sVR/UHYxD4o/P8mhLq/UICiFAE2N6jeEsJ4ewiFb5HIhNB5
QQBSh0daySe5NugdUmo+60RMcjVGczMQklyusbpg0AqgoLNZO8S6RtT2DKdMyGELuyLxWy8x8fwp
dPBcu9lFu7FLMEQ4tPEjXN8kkklnyuU2q6OVQvzr0H2rG9NVsJII5i0jRut3IS+KOD3BP8Gg+v6C
n9aZR6wR+QY1OrUopkoxfoa7DOslaylTsO62iTht6LY3ST1GJpaYqJUOqZQW4G30jCWK+0OkSTxQ
B3vYxLtU07EuL6Vt9wYl2kXfWfnzc16slByp3TikqZ1k36+5FZPVL+HpXwtqpFvTcIoklxwKfr0k
It/ERanDZ2R2DuXXN+eLLwqXtuLS1ItQVOeMC8FoG25FGOCr6m8heDvAjTb+vWavvYlCn2vr24gt
qfx7dTp3QMaCo5EIBYnMa/13OrL9NUY2anHbkXrVoufSdRJ7sopOzZYnTu4FFFFycWZMYQAa1vwC
mnF1/KGUNIF+deO0jGH8aFXG1kYmq86CTcIB4Y9peM3LgfEleflmlC2n++ZIUcqQ7/xW+Hwgivw7
cuIosA/tU5Gh9dhdESMGIioDNIl2ONFhnh+Y0plFdxiLgbGnj/3S9poyE/KgU4qRG07EFNe723e8
54Tlf6FDDFaBoDJvFhbsIqV/D5g/0rS2oJ9So0U4ixsTo7jjnp/AE3RvN8PesIeXSqV3j0ZcyViK
Hn42qFHyyxvQrHb0N/tOSsSfekLpW71sDWGNz5corB488S1xPTaHMA6Bp6gzs6G77uHVCvyJGHZL
PIA91yBT8vs+6y4nEhF5hhJQL5MEbcUw2UXp7K1blk301Dei1cu5V6EIemMWVP4sAFu+iIv2Aokr
YP7Y8Nqfx2A+priYXUUhcMmVG+aOb0i1e0zF/IiJ+vx69qiS482cnUuwXlGcBbaRaRka58w8PBaf
he5AFUXMAf7BpEBALoGQP54fvavjusc2JLylLDup+T2Etikrn7RU03+h4MhJ7viwkZ+bgu+VQ1oI
T/5ybY1GDa18z7DoZU089PPuYdI4HNoROM5CtKuhlF29UHFyvB4znCBGPw/w1haUnrC5njkb3ZVu
GAm46caq5iZrer/uWT5ws23zbvgNnOeeTj2oPKvTbKwDvioBZU894I+rT8nWPYp1Ni9fyHCmGzax
nGCYdcHEvqFXI5I+R/KD2m67TDfywNh+Jo7TSfL8BHlsN31Jjlqk7xxHns33D5n7ANolNpA/6PWT
oAg+qlH797GZRvPP/CtpfWEYMUxRXeIYMGxCEyacOHxQQcSDlnyqu8d+InQWN9YGKyiI7ikb5BBd
8o8u2YJz0g2RmSr2eULglEfac3N5fyG6DVG5LZf0kGl0b1TL7rPBfc8U7yDnnRuth2yYOcn/a3xo
UH5/9Ih2ZmwYqR+Cmt9Z2q2aQDr8Ypcr+rSAccB5TWh4D6O3JsjVJ1Kyc44QPJkWb78C+sE1GMjA
zkBF1nZ/kD5wQ12wN7mic0mQuePtHxA9eWu5Ck7WXp0pf9Hu53KgVQyrFDDKfVr+nAHgIwMSE99l
XWqIgr9r24Lli7EMJbwL1Ylx+PhhEfeYaMik6PLvdrVFW7AE8YRGk8KEkT8MErOAYHYRCMzoD/Ja
MabdpBuOiJ++ZniWmH0fPTOITpDoA9eyxCY16Y/ACbaa5k3z7lR8XZb23iyXj+qjrfCK1/3SIFtU
YRMwhaB17+YJbMZDTETi/n1zn2/NWS9TB/v8yxd16eIatvWslHxBlRfJeRmjjMEMio9ylcbX/r4E
zLkMqV/2DhgB/C7UD/UxofPVTjHOXWjyr10uxWZFadIfnH3NuWC/J4DFQRqcNlboTBBY19uazz7H
oFfIWe0vOYSgFXnwvj7XDO9gf62iVJBHHOm/Bo43aaOcaMnFxMUNnA+5T6KCAQ4x3eLJrVsfJPdI
YBZV0HtPCleDV0CQxsgNscyqqx58URKdXf0ny4q/fLt0ELTJcA7pZcrawC8ba5l4zFxOyD8Ri57m
DnaAE6m0ii2xCoRdUiFRSsVD0be99Wr47Rfwg1884y4f7ttMVEhltcFrQvdHu5hKO5uFMIFVTIsx
BnSNgC4Kfz82bX2WJMkaobFvrEJhr8ncDnhGjXajHHiWBxvX9IWwPaAm6kcgqWVIy5v9C70khlIb
3b8dQ5zIHPts9NyD77VYnWFBzPtWr1xVBztA273vvSG7yy8fadlbqb9OaHSANsB4ocHFbwcx3R6H
Hv6PNwWk2qaK/OdDqPe/+5rt7s10H2/EIzStxsBSxUzS0ENRbN5uAHEu5KP2scgHzILFQ6/pHzx4
jfZKT2DqDSmXGhbh30xxclmt/s2Ne78K5b3AoyR/b9IxEz3vbZUu73TA+lW3CuoRIYrGFJACtbjO
aqIHuCQ7+eiCC34S9A9NsqZVE1iOSR/CYNardyXEBVW4ekgERO/qtyGlS0/gDxKKWP3/+9gG76xy
/5TzjNGHTenZoXLotBbc4Uj5Y6es4vASW9+jE38hcP30k3jn5wx1IalCk5DZ3Z7lhNtO6nJfJILV
ilcUQN3iBiH/oqeVXwjwjxrtLSlJKBVBgvN7TUXOYhS684/ym/aFFDOdPUTNfwRY3PgICNaPL9/j
zrar4e691bW9J04WX4yYTVmNNTUobXseuG3J6KBofPRP+FF1oo9ZRpq2GFnzUy1ISz088VTpc6yb
hl0ypy3W5Ax62w2egHwcDYlc0m1wRjtV0rTt2PEsGdTxogTEL5jUJVcIf42erwgNvXtTfyv6IB9t
a7NbLkZQBkgB8vBZokUBhSr7Lc0jw91SJ7w92/ir75vDwzMVI1WZgsXEVFtpb/amqzZJpfc4OVaZ
5ayOp9iH0mvYyL6iTiTbHMgP8cuFslzvXYo2BuZbqS2R7flbqJkjYX5c0MIgm/BKKs4oSr6JAJuy
14D8qPRQaV7bnqwNcw2KYqGoH+ctoPdhDU+qr2iJOKNGmgmpVZeUGDawfghzOQaLYCl/SCR92YhZ
tOKzhRviItjiA+pL+6i8cBaR7WDdB8LFpA3WUz3Hd5x+crS6EQy7a1KH8T5AJaJPSiWNv+t7vbeh
mQV922tubCPgPuJIMLvwibZ7TTndETcH2VxwI3HT78bevSYTmfLXNj0GiAwWtMaSrVHEV50+ex0G
+W6NdILeLNH/wriZGqKg0wQi83cT/wBz8VraA4T+8wZfugjZ9g6GSRXOba88+DGqdwyel9vy19bh
hiSt6C3RRYqFbNS6CV7d/qvJsNLRqjIbcrpcvRq3i1lLbBKkq2gzkN2rWjm82ZdtsYVfSRAc9ABP
ny1i/2QBvRuNNl2hQhSWyilUy0eVKzhJwO94v2ytW23gt1YyXgPKIHdzYzpmCuvFg9+mzSwtJ2Bc
AQWhmeaWM/kKow8hzsthc04WVGceckh47Ox50MM2Rb7499MUbEaaVpo6D8k+BomkDCgFFz+4b5sG
HFS5w6ZsoUsMZa2EWrbxQzrlveZAyS1UfZwT3TO84OTdf/Fe/SOOmWFnpAwWWQ5x+3eypz0vM8rn
8yZZ64dr3VKPRzkgO80bTctxHHzYaSki9Gmvx2EeDLj/G/tH4F6XBJy7Q4BhTg7DXRgPWfEKemr0
mG0R5FBwlK4AQCgzXGcV0qdudfd2MYUj7V/g3NA7hjrjD6n9iqJU7GbRD+tcnnQaIilH6JnX/JHN
lFpLcCfICzViUfRPt9jC6hvM+oorg+iT4OLtd6vF+QI4ZaEOJC8Q4uV3ZVx9X54r2o1MJyCx6EMk
wm5DxUMCZs+m4T6VoSri7eDNjIiNjomwTAnxVN66qPJ46WxcW8UHpFRHnCHmJZo+UbK0Y+DWYum/
XFKyKoZY7uLeBiQFxgDp+uDiaT/TdLx/JCpnmdgV4cUKT9CSf/C60Ax2wIyQZ5F7EuHjSyJmamwM
1U4aUxQLs9Sa1GTna1RhDtoj93PNxNtiJilCPpitB+0I69Wsic1jXsV3q24jKvQcbI7Pwhb859Sa
8ySOFgD9YaPbCMj0JeHdvftQNl3PdwQGjnoYNek9OCDrm7m5wuc8Ya5BiJcdEJ352pHDoR7WxaYA
/VugJ44H+R2Rg0U3PAnxfBPYC7o/oKgoRfbzFo9uAG//3hSO05FQv8qqpFIGUieB4XRdNebb0GMp
c6L8L3UyoClDglMqWxCg6BdPhQSxmJG4pvMayvqQ6BhuNjE+1MgX09LcmOFm1FV+WqYAXy+vXvhh
74cX5mik2BfqIOtvguWXsKLJqVKlIMTG2ffB7bshG6qB9hGy4ZmUFrlBGYjHcQh/sfOFITgQB25j
7iqmwp9o/cdIK98OPUAHHq3TGodDR1AhEDBjL0dkoCK3onKOZ2gVvCcjPsGKSAlq1YQYZFus/uLs
DVIrD8gZYX7ez2NigLirW8N0yxqf3AFPAUeWbIwXfO5HMsVccr4MnHF+H+0ujz4lXRQZMD7oGfPn
Ta3sDPjLPbxK7Bttc1HLl2meuHGxN7LlYnWhhZSonho+ez1Nxd97agK2No795DUmejftLtEjS9jn
Nfv0O7R0DX716HVgBDVspKIdaA4F65N/bWx9Xr+/0raJwy9KOM2KsvCDwDiVSeDRr3ppvODmEFDi
4piaxD4/okRkoKDuRnG7cVCtqY/8XmDoISo97hGcoN9SDY5pW5S6kPFyiFCyhlbv0r9dhFShxcpF
i8KQ0jhPJ/zScb33oukX53jVA6v/YxjqnA5JzUi9oQoaO2yPA9cJILVGprQ38ulK0yINW9wxgGyK
wHm8jgBNIAZOnvC9nFZKGSQhETDev7YgqoTSfslUg9BtcJcf6rVynoKnENIl/M3yCD6kUespqTca
d9vWMp7do7tlsEZMQ17yCNl7cNZ12DrH9piZO+Ng48Pyp7da//q2aLsNTgKZqe1SmqGH5vv3r7LN
aPuH8i8gzCO/SVzneDJfH4SEhyjF9y8FhenZhtWBnAqYOxCb/qFEQe+JKCungDB5T801mGUoeT0Y
xxWFY4FFnu/vrF2GCOZPLFbU0BkrO4Nalq6XmzLG2nQeNG8dZTkfUyxvIveUL/FQfmvWt/QQNjBF
0z2nvelFjbYMqap6HhTSv1q4KVc+Fv6iKJGx5KwXhdyclQCax1E7sdgjhgsVX1Aem6SHgpiVfCru
l4VKGvN2uacIdivfS6KONgGXE76bHbxelNkSIL2bgGFlevv0QkoO1y4LwvGWgX+TZ7tvAWv1v/cE
6LTxz/edPyqGQEnn11JcO1ngv/hksKeD1oCvdoSTJgqvcbN38wCQmtLctNhIge3NsEa2NhQBB2hL
XSuQppTY9GmCvyfGV135KPV0tXozqHQ5yeUNaAKZZiWxR0cFHIJhuKVduzzkSGhbuXPFTxVEu3+b
K90YxhHOuQ7XoM8a+T0ByjRYGyjhIF5aKglwNBYGsaKPf3I2r2rePkrhF54WD0RLRs7GQE8xJB06
MVFfcC+Ri4YV7dOahG48FUNyQsJXtH1cFcuo01HJhXztLcQcFsQ3sCrycC7QJgEiZDhjRvmJn0RX
g38OFbfkSgDypvoQecLmAw1azhXUwhS7mxIh0pc0zw150OPYOZhHpdx1zxHlcwP66tDot84MfXyt
0UkQKtIFAQ4YQAMW1DhKUk2RFVNCa9QYKqzOjn2EBsgdQaolnclQyIsckW3GYUjvS8oDuXL8HT/B
D70WCJ0xjIwhWp0U8E5EpvEQCaQkYD5bByQy+p6DLNbXqylhg06ONk6phlhpY0L8B67YR1ENeriu
cithJbxTNdksTo8lH8tu/ay54e2aYmJo+QSFx701H0Clrv8WtQ9UJcFpMi4ykz98d8uAg2evjJEH
wi8QbR/NgxHHbCxeSkU2fPANkOaylkwXFv369v6HjSeRE3hKWi/XFIUbUi+MxW0eIactiS5ZBySi
QnFaQl7Qnw3az6KxjXQAtCLSObuBglUA+CAkM5jx+Qj9+gv+b+aHnon82CXCYLXVHV23maMEr3yS
YpbDAJYtfI5EW4fNeO5zK8VtZibBHC7gpjaphFC/CAIHnOH9GWDIpslCeMg7Wfa8RAGriEZUzQRU
OtMO/tgVVvy/uEYEr1YUU8pQ7VL2MDchDbIp0eOgPzvmslA4W2OoKGAX1MoGPq3ELzMA2Y6vNJEn
vJBZKQpfQdHGjCP5x5uqLRpDKCwh8LncJ98nDyXFj8SdCg+rCd8v7bhCnQnOx8Jusmfb69S5UJBp
Sd3d3UteUv8SVD9nc04yYdH7sj6oTcPbitwD8rEr3gTbPH7Kn2KGUwYl7P/j/FVUklzgbGCHUnes
KYSERJmn/XLvnty25jrj3T3CYtqlpraCtR+KjlocXYQPvYowcZdYzmTsD+QvlVyepVRUpnNrG/WB
tbrkYU9Fe7a9Al5FXekIRwHlgZJwUWZYBnzpWNZhBycTYCSEyg1H5ETTINA6/JoKMOz29pK7DpfT
Dzi5k2PDqK2VZLqMFU1ac+pAWVISrcoQ8kuiA+/2QGbjB8NEkIoaExdBjsofgufJMcUZ2K3F9IuX
6OsH1gNFrwgY1wLzeA7jRMP3CrGwx7HJQzgF3AnQ43skCIj4ijP0Iq40cVkeRwpUSbmwg5F1WA4K
4D4hQDbDNwUS8doHL/NE8DmN9Nni5JApDT7PUidFx/hqiHRIcHIkXkzZubsEF5LYKLlRlAg3ExPv
TXlt06qzMxACroRAybyIKIuN+a9uf2oTkukEGXB/z2wR6PTdNWz9vr/CSE9laFbGDVGpBaKqZWiS
KdByRqcsojPZl7E1X/PlR+FJsGkVU6ji4dcarlezJjrJz2nSH1t8VrtYMP/+KQA9/s8a0OTjB/s0
DzIH5SkUVDCEcd3bZIgmJp4Dibpa9wiwKP21tDRh6GjNYvY9idqFpLNJjGvnNdrzfHdZfroVEoa1
9LUf2wdadMYYj48e+6BBz1XeamGQj8iBwG7X+1LyXArOGw/QO236nlbcsRlQZos9WvkVQ2otIA9a
a6JBG4lLFHpvngyxxnOkTZV5oiWOg+1zYyOqoa47lcjSOGYPMnwoDbve+NE7A3I+aCaSmhepTeR3
0JDE17UpyG+hla+t8qAPk/1sJteklfkp3cXcbb2nyQRSomN+Xn4BVIwMAMs8dYGX4AcmBZYK2CXx
BAt0JbI/BYH4aDUv6tsvXTTvaDCGJQiVuki3S8VxM7wvF66A2ZnxQ4JG+N58UXWM/Va9P5Ru5gic
51N2Vji+bf4RtHDMWAixO7YhdQFUWhI5xYPXaVw5sB8g5QLtQvUDO0Hl6Q9YOEZHviR0Tf54kHM3
tPESXMowXjMFK5bZb5e64rgY8vovZUnltPeBCjgU4+3TgliJtEPzSAErNkuC6nkm3LWmbWwK/+Np
Mi3UGw3J9/nsVTijzkkIFdJEcnm3sEmpO7XvRlP7dTcR87CRPNGY69pSCtMarhXKmbu1PlI9EOC2
VSGhSIoQRGDCYrcrxpuFk7vrhgcjae4Eme1wj6ZLUFAp/FNeZ2nG9D2BKnYn9n4WiWY8FMDCRmTe
neGpzyAfFWrwg9rvb6CVNHZ2ix3VqxNUPI14LHRn/XuySatwZEjW5bnuWGpXoGIrryu+de3EH7rA
7WarGNQe4JwKTL7c0D6UmC0rC+FEBEUGxyAU3Bsop9lROZYKBn/l/j5Xt1rPOcUyKcD0vZz3v1YC
uZqp/dlTKu3K+jnMEVtvdKizafvLbSTByDACq/Y7YxljbGGz4JVgUhKQv0NbaUGxNUdJbeE+RxSd
Nz/8L2DotWCPATnddJHMJnJFaxVT7gfZuQv2VdGYQ19418eGNvR0gcSMBN7lhIEhdfup8IgT6sI0
euMR5NHcnNbiueJkszkTwU7pdKdPBK1a9uBEN/j4NeT0IOh2DXNIKGfx/OsSzNgS5I8pP04fRI7j
SBH5xa4Rt+SHsMIshOFB5hIELDHNibTGcAkbctLRqyfgOByw44aLz54/Ioj/N5tiVuqBBygM4Vlx
8KnRIi6MgPSl5EApP6pFoQ76jzgFm0Qr9oAhWYskQhIVqsxSjHBykNVirUSQFf1xw5mUwX2YT70Q
FRaL08V0kZpw1lgstYb+aEyfGgmBgCS1B4W4RWRdyvYbaEdPh5vGDS0GSIXuyM/58RwZBNd9XRA1
BOYKD+8aeoJ6pwTPF5Ou4Qqb+Kpfb+8X0sE/yK6MdYHP9BYvlqTCc7rZQyiLsr7JowtoJ6npvrJj
8GvZQLTrxinH6KeVuaI0ueVGsuodI1Yxs/I4YNqXIawydQ8Nd3Z/kB77bAHXHCQx0mMSV9QDjpCK
IBy3Z6iegHbf86bMA8gcwNaUS0B/B5o7VPvyoaDTaybT1Qdkc3C3+rxC9ekseJMnn7qGSUb8EgZv
gneYzMiVtvumDVwkcOcsFJ8ORz9sjnnwZJbdNwONHjERWHJLQQgec1S44Ey7zXtbK2jZ+KhrosC6
6+82xz2soc8Ud7wZgfpqu4MlIpom6FJevancQY3+iPuzXhJiyQdWuhOlqUJ70g9ONh4RaS9RLsME
w8IO72u96sR6QAr349udOUq6XbuOzEw2f+3tsHTxMKGnm/ch11dgjRCf+pDrZqcHsmk9fbGCyeN0
MwBaCGlvAfg6ZM5XmPkpvmxLGNvgY7YMrHPBL5iuB0V5J0Xb75UFY7Dv5kg1UC3J7sgJFrz+As8E
vbJW8YV1hqijXTsAfluQvugjg+sbrvzpIz78OrfUDdFiknmGsjfcrWeV83+iL+tEptOtxXSx3k7M
qBb/D4hswmoXV/vwAjbsUxwAUt4Upq6t16T6uK2YKhPZ3hK5IdM/yux/kZq/hWvLqZiWplbWhdbD
SPgvzk33e70tcnUGDjT2ph5TriZ/2EdLu8v6h/kOCR0q4y0zTMS5cmdiWAZBecJLx5rlSZ7q/0kH
6hD3qm5jlnyy1/IQzaGDExO0WsKQ5SCN0dhgkaFc0QUXZ5nHEtB3C4bYSTDNmzWanOAFIP/gEcYJ
vN5+Glt7ipuReGHIJXcT9IVOFBehU+EzdTu3NdkbeivaJoTEwYz9a33pt8/wopeCaef793KzgpYN
MdXs3B8C7VZxojmqQ8iuvw2wv4NamabU3fnjQ9m/vtX/QK6XRj3ANOVn+fwePVSitcviGx3yMvba
3/RP/+2IhalA1tDIfutdJq/VlG3TDOSa/THYJaCA0xWF6Tt26nsgWPeX+Os9jzi/UGqJwqKaU75P
x6DKDKfnKSuoNFk2cPnLhmVUD0ySGyDFwgq+xSXMxzke7CBMcVWSWrQVcXOcE8X9y3nDvhDCfiZ4
+qjw8bT0dDvUu4+R6kZzyv/8iAvv2T1YSis26zVfOCOo6cqevjiWjKjH78Z0ihwTJL7nn39viW5R
Z3QdHu/LDLb42hAjjNUTlOaWPDUOvNzRadbOyOJmF3nUnF43JyYkSheq4i7lOVqGHw+Shwv5cVO2
YsFDxi7DvFb8Dt3uUrhZrT2InF9PqSrEkN3aRa+yDUk/FG2Yi5bSKkx/kYk6MMtjoFapgIiZAVNb
+Ailx3kCvWHmJpjE6777uZbXLAkK3u/Whsneky8Za6RsndamhziwpV4ZN8BrDRy9EEzcSjqOS06Y
1k+MOgRQu8W3pOGGImAngpZCV+ySUEJGVI3GYPW53gWMdvWmR/GWOhdEBpBiJJq1jscyL5zXu7vL
kzr30rLOn8QRNolysVvsTp2oymdmo4QpB2Pw+nZiysBmrI408Zmyr8ZjLPwGfcr3iq0s7eNZHgzE
/N2weMQhJUi44xr4zEoTGl8nTxl4PffhDMy4IdMuwSZHbdAh80Xff1sbeqEomH0w2r7+oYmxjFD0
lcLO5kK3TWDsoTqotI30AwNugxOmtEhzZ7UfLIcR4wp0dh2rfc/u9S8SoyMF8sM7D2jpEmu4macT
Hc5gjCHvyOEP6SPdwXKw7vxSJigBhXZDu65tqQ/rxlZx4mhPRi9hal8ePvRNol6dR5ZY6sL4BWoL
O4NFoqFHR92HV8eFpHdVP5aet3UQe6rpO1og7KJqGBj+HAS24pdqApNZGouDfh7No7rNqqMX24Y/
ePEN7Zqj3Ttt+SGxw5XySGpdri+F/poVchF/kaAeYxWNoMSuXubX/ATZT7otA1ZOK/JaEDAOfuc9
cPVmT6FT55WG/EBOqdxHhSgM9TRNg98abw6TGFrfu6oxii2ZrOt28sL8px1WrH+6cgyL5uNWJ2e0
1hqswAPmBC94V2yuFUx2T/xvq1+A2dvzNBeW8IApiTR4LLUta+/izQWhfFnroeRKAvWlLI8y4XJF
q0/lF0zuaMmbHKt1DlG2egI0/7a2XC2j4HU+KT59qYBboBU4Q523SQSIlCMpkIl7WRVce6anAb3E
Abh1sXMcMcZZ9L2+jDHi+JpAiViVeIxbJLT7YQdR10Eih6/zTOcS00X/+vwpmEk+ArXIWC1sTpf+
L+iCj8763TlIWIwPAhT0NRfADYjsi20r/NTRcc8oIPgevgYbVDToYBxO03WvO/AdN5AnBqg3aAbb
2SOhMfxkA9KuMTuTwIEv7vgJ5XaA5O6CfY2UReMcN+/AI7YjlwHXsQbXMMzV44n0rtTfzI/UG0rw
T0vwGnUWR6AVX2MmoZZPAnFZO/3B+yVuib2PBYYTmJ3naHYnz6Sn7ckTdfmUeXnS3rgKcsT4GeIl
3WTWITe9XRSIzUCynn27Eh9EUFSsODSs//PMN0MxJtVuHzQsIOA3t9GuPlsRbndr7k/5ZEX0ZK3U
nm4jOiPPmBVp449xYqLhBMwfQ0A4dZUDy6mtSarFYqdKxpCtrmB2yu2ZQpk3Mxy81BV0+rjrmZMz
WQ4iPGjoE05l8gxdVUpHf+2PKjOXFNiquCwWie8ZuzEfZwcMhyjRN+wEnlDYyBk/P+eZ5kzKSe8s
XiEIqsF6Ppr3T8eS3aRCbI7P3LOehit4UX89snjfWh+eaeU2247hKXXteH6NXLrqZG46KCwri5UF
saHakkYVZeum5owqIs2AY0njOzyawbA72huNrlG1rPldGHOB3MzsOKp8oj1kGEBLyAkIPcTzZ+Ud
oTgxqHdysNghVIcnej8sRTmzJyceQeFs1doIMVyUT9FWoGONR6/j+cw/wNZLFY+tIFgyUiREpQWl
XEp0FGJ5wHD45GxlaINg5FhW7TbpRA3YExlr60T7L0EE88qPnXqmcTt4gj3PrvhuPyKk8E63DxXt
fSaoqcDUSxZQRhaTcwGJUXg1/LIr+Y93juYmuyrRtWMykhkMy3okqr1Yc0iMWHbEOy4f8xW3yNyU
O/TDaJ4uRZXEr47Dvm7olCl2ECJW0KWsYsPGQGogNctoKO016nNieM8fCqKrAZ6Ukvwkjtqaqvj5
WTQXJeVJTwoM2NGCpoG7Zhng6nQEh1roW8bh/JzdF4S56D7K+gTzurWfowOF0xC+cFlSrECDfzYA
5myR2ZAZLyM+iVZnm3vnr9nK3ctQ2sH0fy2pjsHN9+U8o0BcZ8VP1F3hTZFL3lNRGq/6GWh/JThU
LF7WcvFRe0UwsdfnuahovFgO4k5BKk+h663P1CvanccmMh10D9tjEEUF1KtSGujF54yZ1FtgKajH
SGTRjxd2rjmXJ9Uu+T6Ickj42wvqLwHAf1QrsxEw+4eOJjbuCm9o+KV3cYhxNaxuAe5n2ljKtd87
ZcJL4ElynNWqMEDD/4AS0mgYFQStjP0CoGnQVEak293zx77hFJZ+2X21QoVlfEbHnfo6G9bLZVZY
/w1gGgLXkKMkb5KA78kqs1CV1hFWnBU8qOlyAaP0CesNywhOKzpJ2aTIwkbeDcsJ3yGMpNxZJxW+
BduAtINYn+RO3M96N8fHhUkl7hgiPpioKfGbz+TBNl0sPjwxqTZbEwKGAXtoR732jcRSpvd9ZwD5
uYuPKfpiDSCXvf/YxNUARq0Mv9FWj+yd80jGIsanXj1g2SOYJI6nTyDzdQ/ESZyyyXoSLEItRIg5
NtoFPBM9RZ6CmpRpIeOD7WVJnFc8bxS+VwYeZOd+2lNAoNNyCYi8wG0TH4S1fg5S5lfEq7HV08cy
JPf5WgTzv9Y06zOXPgQj0tbkPwyf7ukX4YPYrNTOGcpVW4tH872pl9ll8zLlVQQVdgi0fzGqey3P
fpMuPhOGiX5RHfBzdaTYYHQkjQcCO9yPxYdJR0K1KvHo4lMMw7Hs42eFAjyY8vR2rA2I8eTFwHzw
m7HeYlyTk9O65N8MAB/hjKa2/DCE9vIHaGvxt75Wd0hXUnMbYSy4d1EwOUB9llcZE4VKjzefyE8q
A/1cIDK5uYiDQQwQ1wcvCoSkWxAo3CvxZ+RgEjrtxrj4O7Ldpve6oi6D0LkOmTm1VhejRRdP9xAa
WwUsbA45h9kSPvporXYzSD7BCqPYGdswlZRR2Ou49fGtY0ZCvyHtYeqpZV32p16I7YVoxY2gumIM
U1qCxwl6VGWhdhOJzBn0oxaCyfsebB2KcE1MO9QOuigilNOsCayWAVs0K06/1NCrlw1RIXFgGXKv
9rvHsR+kqmIhqKnFQC8rvcmu9q62UbQfrClhzgDSrT1cdgyecqvan9lhSXS4g0EJcKvEh/KSkYTp
WvT3hqvbZ+ZvXBQKs79vrcUda7g1ssOaOQC04mCdH0/ASPD5a+dfQDkQ4aNoNGYvTlWXJN+zhqj0
ZPRiHaECpv7Rv563jMhPKTssEK85XU4Sh49+jlwX4AGl7ZRWhBrF2EBJI3BX/II5cyHkKCaUsck3
V6PhOzsFj7JwxHRu4SEBoeVVMs+IbcJmjNCRJYzfFYWbjlcVB7kBFi3KJ92CKFj2w642givcvpAH
9iVWD6E3jRHSuNFfw0zkd6pTrXB2rhroUI3MhaRiva3/+ouIsMY1NDhQEVZfgSqPSXfr+vMyNMRO
wAlHY4IHlJII91LWtPJENeGSW6VAZcrWT1jQvNjWNX80Wt6RdKXGZabmgEt/BvTICYdOZ8bSum0e
DYGK9TwNzKD5SXxmWK3BtbjdjWF5tnA6VI4r941EuWD5FMD+mG6FjrS38J04WN2ytV5JrL/xoaKF
vR6B+Y6krHmkrwvofp9Fz+n/+cccWymJpTnfHDOjbCkB16YSbTK7gdGeQtLSec1kxnosZYky4gXZ
iV+VhShCSzhMNTRyb0qA6ITaXYYoIVSFF5niLL4LJbVn2ZkBIaVOZZSgDoYOowSP9wHCgB4lJqvB
hFXTQ/0O418Plcyip9Ajx3dpCiS+/DyUJQFf0TMTZ+U5O//MQEKEMCJGZ1+sQUKT4L1lFHnzNMPZ
PM+x/j6ceym5lWySRD7w7yzTC9nslb1WGaaj32reoizhcTqXB494lRpPlRCHm2lMxcV622x8WU7J
i8/9fCQtE9vDEXYyCDUVn3xWi/5u6/AKSkVQBjeXVSm0FwkukQHP26BoE9ucH3YFzoRMkFJ7+p+K
iiDrN9kZXoUvDzbtZjPXUy118l+kjmCXI4tKC9MyJ2BrllxkOp3Md19lAmBOVEOeONRZaak+K2eU
AJK9trE1Ig94oQJhM3myzLVmAqn2eM3EqLSNH3WqgGAk3DFOv7ykuYpJ4yqXgizcHHnuIjC56d57
o09pPER8lg3wwGPncYOoPeZWLhXrHHMUgjcbYn+0Dt7w5/9JjRVz30N64Fd2TaraR+F7Yhn67MRr
74cO1xlzhtcNa0HUPgehXrYkGnYnsNYUQ8/9cuuNR966PbZLgVaBWmktZDpcbEXviR44/CEGYmoW
7N1OukmP8pTEDJQYHgzE+1YfyRiLkSLPtnrhNp5WVl3OUakMZCKGuZvmml0TRF/CStIv85lK1IA7
uu1Eutkb6bmp/NtwY3vOJVaFjdYc0ISf/odp2aIoeBzzotXtyOyKCMV+n/dQN2JT9gzNJL+TZn1L
0ATR4S1rorgbKrTaDjoyWKzK/juyeG0Fzn+G8vLqFzXBSewHDM3yXmgeETX/Z33x2Awu/VHNTpi5
+F9YU2K1vek1Mz8DWQlKqxGGW6/DjTcI5MX8xXW13CrbFvyS5B9Ug6H4a2agxLbkaBKJu3vNuv8F
6+VkN9yf2UCsL2OAIe43OGYFCkAWM0AKgkT4c68wj5YUeoRpBjyO+pxMC3P32UUtwedqo0jdp7fa
4RZ/C0baspo4IzWk8hNymCfYOudv4qNq72nFw7zD+x6Ih0CfhK2/3Zx0qeiC+xHy5gR2jKCaQY9D
U4Va4qDKKqxNhY5+SqGCW6OG5zmQnAlWeIE0WbG8OCnYviak0GSV7ebHgi5xYw9lAbSjQOrqivfb
Q7sHREFz1cb5PIavMvFH8hS0k7yGb3tTojtn5/luDWWqQoh33NuVoSJyrLkRPxkEn1Km3YKLiOX+
ZBmyc2dy7s2Hpe4OfIFpKFHXva/XuOWp/qgjLpsz9pmhPiyRp+K2d4LVRcktusHuPuy8MtpZnDfy
fZYMZ+ySXjcveyj2vZplKR/6g4OcOrFqgrQSgijf9+mHnfIByPQruQtbBlHMarA6AvHPyWRXL5YX
mMech5HUvEJhWy/44PKkuiRl0K/jpxOBIksbCRkI/2tNuHTSoXYYiUhsrrp6Wkh8YuXDmI1zwOha
IRlW/gYfUTw2E8eibCgoOCBbYZG6HZ4PQ5QUL+dedcXBCfTiOUtv/UnbMqPesRhHvShsm5g1Ihii
QKhDGoLibGqk4U6ea7L+77bFR5vuuawOxLsogotRULObxAta6kd6gguj9+pnRy3uAZ8/6iqxOA5p
tn1d8QIZNZ5gmxGBQIkCxayJnvE7e27iZ1NcQGpfmG1h0HT9a3StWW1zUuv6/mh8qLwLA9OoY9i0
nao2q2xLoKvTDu5uMhn6uLsRiV0KmROYilWhuzPG52H1ApbCG1tqg3tSGVrWMf7i/mb/i3Zr9DfG
2i87N2/ikKrYSSLLe31RC1+FDb0vgBEaemh6nAZ5lwT2oc+U1w932VuOnFkTEOMlCFnmByS9akB0
zaBPNN0gnqEUBCsM+F+t0lE4oEiH6j17CVOk64tQPpDc78g2FD29X4O6Yi7fIIaMJxuyK9tSK7TI
Wi8j+2c806xMPG5AKTy5sZAtYFhBQW7npSTlcgUWGOb/hmQGSfpC0Rz0ST75EmS1ggqsekr8ADmP
Jnn55Aa6lA1LmF94uf9mYL9+LFrnGlY8t1XAd2W353PqKG/sFEL+EVwiknfEryico4NstCa4sn3s
/0xiH0Zf3bPaLSqFrX3CQW0olxEKZI48Sbei2JPhBZmj1UYKGJqlV/9kmtaWoVgnVBxXuB7T1mHh
Ea9J0v30o051k3SDIAeHfCH+9qC1deQ2oe05DEv/qeG2Y9UwDMrzpczTWU97t9YzEu97Xr4CCE8B
QXaL6fY1R0RCpgnpCfV7plw9rLZyKE5rbJyUPPqifOUVC8okSCWpCxkfyGqKcjMZeIVaqe1KPwC9
Hz6KWWE+YubdUIf0EvgTXIenLsPqmrmShkGmGXL3CgH4+bRSTCwZDvbPVpWqBmUSbsX3SRaO2rHm
l1P8OOPK7CJhFw0/SXIMcDP8YMEoEk+fYMwPHYAVQMDnPFjy4Zlpl3HQTywpNuzZoT/4uGdCW6Bw
TkpoZoLLuxkTMnpXyhCn4FHVMR/thGKkDofdeZBAW60b5msRcQVlTKzjdUrXDud81+7FWtJhc6h3
UGCw/xD2Ycn01e9pJzZQjTx9zCCH3uuLwGSyDsNJtOU5Oxm0pfbS08AQgNN+Hq686IiZE//aExMw
2KAChkEiiq9AqvrzD3sOOOxiq74JCcYwbloo+sPKGDF1NSRCqFR5CVxPXh1x56cWKC3yx+G/qnbh
Iy8t204jJa2Q/wY7Gkzm/wbzbeFfhh/xICVtiuGY5tU1QXQpdkgFypXNq0Z8jLyBO6zO8VFYjgs6
cJP7JdLMlvN6mHXLPlHM/6JYzpelL4d/xGCUr2WhxYtlFkWWBFTw2TF9zUKUlthv2VrkA4XJJ9Ic
KBB+iCEfbrIl+ND4wVE7vtPgDuMJmPBzDVbcMebdKVE181sbNLtNS3Gn0Q8QIL/u9NBfdlLFAU7i
64NLxiXvNQExwRr7QAzrbzEUas3TqsZW+Yjgb5ONEEdF0mwqsx2KTT64B4dU62T9bOUX6cO7HwjZ
8aNwtkkEic9YXJOvERPlEwuZaxiSW+cb7rPlbZnghJYYeiACvsYYQ1Y2g4WpksXQKFIXrMUfZvZb
UJTLhETlasPOQFa8IfCKUUjKs52NhbkJGgVEsljO/HhelYA3LAnv6eRYC2+RAbSf6Y9PC9wr0eSy
1BA6DlRMKbDXWwKB2rm+3hWqBa7+cCONdc7AQ5Hl7f8BygUUT8cFKKCrYxvtIgEM0a4BCt1gyhTo
mAmARYdu5fqeKNYjmr3Rm0WK+oq6zVXCdHKucLG2UglKgoeVNVUdwh/0RobzbPjbr4gGkrMHCTmz
r0EPINco++mxw9PqJ67ME0HyiVqBnAgBY2UVlmwajPw7dZD5OUCLHqHfyLQce0r7cBEG3WISqELa
9dB8Lh8Pis/fzkIGWlb10FZOI/GsxcPnmFKdUoIrzPnhBbuXeXAZMUdxwa6bpCat5/u2O7w1iJ3D
RgGVap7XVDqJFXO7B7WIozrfk/S1BTh8jemEA+NDddgy4cdDR3e/MYzNNaeV6pJqd52iVmiQCzlt
G7Wy9E7cCHtFkCLNcO9uig6j79su1C1M7skoltM90rpTaHJCkOltpZ4OiSNY/LvkyvpD19w4WLpy
WezTM1QkSq4WSvYJP/NIOXHfIiRFxdyTY//ek1pdofuqkj34aqZXhxfgyhGyBGaAdIvmxEl7DxZH
P99/2+wrAXhdIPpRSoEchyK5v3FXM/wfg5lggAg8Ep1Li4Tl+sVHo52lqSNVXP5DNmPiWo3eeYxa
lKH3K1UIwUMkPOzMXGQbI8wL/cu3A7OCxW7x0R1zz+DMl0HdbxTsPf5bJdmk/y/WxZt27VO8cbWM
YLBYFlQKidZ9hUX1UUUgyEaRJrX8cZxGxGdyrsRcOMdZZRAeBG6oudRUwD6K5ZSWqZTrQTjNQL0i
oPmgOX8LR6hzCEo/iwsNYV3C1P4hPlVsKMIKle7lCR8tQbE1/DUNQ/XDNMzBreWgbQ/3XZh2fX/8
ol3whYANmEgijx+7uNN/5rNHkGRCZ+eQbb1Kadc4G+6lWyxgNOafpE2m/diF7EoECwKaFCI8eGJm
4wGzoVCx5+tw9Tn36Y1figZwPKwxXfqZzaUQ3DgGvbBVMb1SEscCvndBY859C5Y3QXwxbasZBtCm
CutO58+IdPup0x1FCoitjEy8XqkMZ/eDlrm3udGZotwg/RIFF/u8vEHwkGp3DZbw7uzLsRoufhbD
QYVp4cMZAY4ee94YY0ZYLSKKzCvbu05BVzMdOppzUe8GblH6KQpepjjeRJDVlNDDBuA+uYyGWcQy
IEiBfb9hQerJbYyhtO+nlAs/jlOd+VmBrfZbdom9wwNzKR1qKbC/avA1GgfSQ9gbFKX86g6MlhDv
43ndEGEVNLxD2SyKm9K3y29lGu4+HRHAy34Q7NBUeIg1JKV5a+/EtBD/WgELyLlPC6bysZ1HeE0S
nxtQvyjnNYNl67fcuey2/w0Yl/TKlqlw9e5BszLgXsfnsJpJ6zY3Ek91+7mJuq0U7AwdxTv8hmIS
IWdmqBQRE2MRfYibOPsp022sEdSbgb1fA10qsX0Fzglf7yzYs24nADlv1e0bxo0oPQW5vS571RLD
srHGLJvSAD7LKY3jAneelNnANNy2OrnQ3EHrePU/TZ/Iz2Xa4ejZ6101dAbsI0yL1SHvRT50gZBj
IQeWGHVOW/h9D66kWsw4O8sSCPE9CwrmPKsKP4G2cqv1A/u5K0igP0oFi+sp+RkALZjfGMFii6s9
MMoYOlVEnY0Mf3hBhbRz4wwdtmSW9CFgQnnhV0DNuTNHVJKLdX1JHqLw7HVbj9E1cMbaApD6ssdq
hklc1Eh6KRWssAuTNV7obkAe/54vFqvbkz1IXxTJ6VtwMSeteV71DgcX52cDyd15RphKbZTdQ+h8
Nz5i0nMA8x5DaItxhRGDUw/vuSn1PPBI3D0oN6HshzX1QozWI4xlYJ5eGepPeyX7nG1unL4gvsQX
tZd3pWX91PIhwdoj7X7H8AJuyuVaaGWZ56JJbrb6VPLHJo3H2aYDtY6k2choze/JvmuzPVgdjdMB
5aWVHgCM8DfjZPBxStgzeuAaUoVtrf14wBY2m6XgVrIg4fyTUF5sw9qBBHwXirwgSJIwEWphJq5X
iZhtOBWVL469dNFr9PJMHKR4KrbNu5MuEJcOZN6TKObUUp+k8si4n2BUQ9ZUhq5mtQV7hEF7b2sl
ZW5Ibr1LO4IT8GoUlTxY/4rcl9U0tKP0DK/7kLv0csZnVAwer3O1QummheL89nxz9oAFwxqD5PqI
X29hj1C2P+wXAtLv9hoBnE9bMN6OXCQ+gy0UxrKVtxDFeNixfVIcFbB9GkVYTsMyHXLmja7aN6CS
g2Tugo9FAMgTDuE3DCVs3lGdvElUK/vLcsyIn47ke05FWsKI/DJr+QPNJjt3ZJhcQe2h0o2yQbqw
LksccN2iaW86twhPFAZukOD7QYp8Y0xTI1vqg2ncQD4bS3I7QZGrdm81QWDED8wnc/oFM/U5yJ5i
9DzFaE7NnJYv60Ipc4ioQSBOBsZJmqP+WJ73ZVmTAKi1/VVZ5gzSwH/Lb4SMDjWTMevYfYQr1BnD
UA0yBhtJRwiFmcCOd8nEIQ5ZqUYsZ/WFRt45kxItgYL9vy4uPG1fQLM7eJeLu/feICgy14CDTcbp
SOr5O1XPg2bG2r4zOJLb4slYT2eUoyShRnxkUsrTdNFReKARH3/9BQ09D7O12WzkFr5lPg6pih8G
PzDvdQcHyh/Bwx0frh3eLQodfgQl4dTS8ltg3lP45CoSavCgykbM8jRWrZVf9M3TQ/lfxyJtB9tQ
lnbJ6VBgQKK5JvGHtxFTCIEqqvtX8kTuorQkXqEx2w5YljWciKVORfhjU4aomXW9jHIiVXgGd4Kw
5B0sIVM2rCaj/2XZ3a1ohMM2HD5epOcL+dYr6zh8Z4FNW1VfQSBHDuB2gA/9wygnE5Ufgdl7NVip
QHNyxsFhwM2J98snfqCIy0va60sND89xviBl/d79YEW+lHlUh6+5d/QcU32MuWz1WFnXEoj2iTNa
HUhVixPoIam/e2pX2UYfYXL/JuWmtY02eWrhyVCaGWOvx5G8LjssFDNn4g3xt9u7jVNE3HTisf1V
+qopo2ejql30OQlTbvbvlimchf55RLelI/msxg7KaZHjgdQ3gmOD7XiF7Cd/iyT2NewmjDP6p8yK
aHS6/9JY8GaepfTb3MXP8RARaPNxRptaXlFFVFxrmgGE3yexzuNHKnmPrlpg7+o6g+u0CU0Sfw3r
CnNiPIY6fiH2H9wTnjnMd43+fgEIqnX76X8zvmWTd1A0CJ65KwQjZnCm1n+yNv6v0dlBtQMfduIM
nu1ddyiUcwMQ9mkoWbfr6JIkNpmuNdPQq3sUG07rnzTRS7sdWPavUtlfW1KoJTm3wPWqqLQ+RZ5i
NoUC7N838Ihn3SjaWg301C7zG9TFvsPWYwQzpq/yC45qQW70KhtOqdHcjlLH+ikyrLwsA/5R2IiT
ga99oKd83J0LJaB1lf20ayU1hnK/ijPnSHE+LnJIc6SlqN9/ISB0ObB65YdtZJ2ir/wLvgZyGGxN
ZuLWeujIp9gxmkcwQnxBVIlqdAj2WEhvXD5HrW04ADFpta/W8jqihhH9f398FTlgWkLCicp6vnUd
fODProaq49lB8SA4zS0RAO5oiO4pxvTPnIuuXbZBMcw6N0s1sUdmACEyI95GpRhLZTIDobEpuJhk
ybdFbnL9I34i6nlg/Bgq6eyOeHWZQFw6vE6+wBzdJ7CnLhrWEh9/QL8A40tAvn1oI5T87sL9BiLq
uJCYLRvP37+TxQtEBJ5ec4hhvkb496EtaP09VgJ5ItmPEl03NAsR8hX9ydrVqkbz8DKgdRuFJLQ/
ahw9K3z9gBpZKBH67rFB89eh5X/ce7zUh2V40/6usEYspyWeHizoEpKWJJrIPkEZ0iCqxvk0Amz6
L3Jd/mti8vbupKVrFk6kVRPGeFEtsWlmltwR6s7nwlG1iOV9/W/I9PfHvxjIP3IMzlfPwu5vFNwc
moZzaTeREvrUCVnX70PvhZnlc9dZbq0tl9qVp5rN7jEbdC3GGFPoYfKuqhPx2cSEuw5DRE4+rYqq
nRSQTvi6r/yU7J+D7icuJ3nHGE4QO0hCYvuSFfT30g1tskX6cwbU1njPBwxuNMUXtdFCiqy9cm52
p8vrlHsVJY1bEIG1z6weQzcJpmyAg7WxzvfmHUQmAfVrd4p+ol925CgJZbc7Hgy63o2qLp6OSfv0
6aF18cOBOxpvtFXsnRJxdpS+IZz7pWFOaXYwTEPoe4ZP1Q71AAvQZit1zBfjBhm1PiUln+Fh4Mf0
SJR9kq/uBKbdRE3oeu3hvXqA4CLSDkq+hQq9C+UTVkBIaVjBcZnsfK8RU/hN19vXZgra/8er63WL
KXyq6voBW5sXKcg9dUEOZQBrQmzJqQ78DMP+sE0Fm+zYK7CFzIq1RCdx/SMJTfytSdcgjr/ixEGz
3MO7LP/yfhbDR9ps6++ykDPXFoeYyx+9uSBaZF4ovQ5Hwk3jSbnizaHxHRQpMjoQSDmxwfYpL1gu
QlBzmf/NzOrNS1CB50EHBVGZuN0/9prEZNwAZu+PdOqs1+DH7QBnxuvV9sT2PfTDr4szfQ1VdTJb
90Fn4QLr6j+N2sA3khWruzvyGI4Bk1vK0BpO5+LzfJ5aQe0+BSvDidmMmEFi/hVfD92bF9F72Tis
+M4fDE/Hz7SvK3Q8MB4V6ixEo5s27d5uyVJJHKhHB2egnviTjs/T3MD69+T51rOnr6VUriWgwq+Q
xpEKz0OPa2erOCY39iP/KkXhf55SWhJFjoV93kbjFTgOj3fqsfc6IMFd9yEELfIQSBIO3ZaQXpCu
iOlFrIQHCf8io/AmuVsxKCTJvARdMjeF4uNFJlwz1+6JChJmlhFm+pnacF0GLr2btcDusF2yzJV4
D+IxH1J09sqNLlvUU9FDVcTUDIOAvuXHj9+cHAmGt+bAlLbv3ETDT54HjbqVJKuscz24dvFpfbTR
HDrL52LtBlDsmIBZ2cy9h8qiCHbbvWaM5fdh2jTxed+loMnoy4hjKj3tyv1jCFE6C3L8pwzMMm2N
fukI65NDkPy+9xVnTxJyPUlNq7TXuiTKjwVn5hCeKvmO5UztJbgFwrCBCNCCRu2eYdbJPHswDpPP
hTgkYswiLxD/EntlFaVprIYy08qZh46QI8G+M8X+qpyJiCrgeRSu9E7K8zJhJIkytu11yHt97wTy
Btw20/yLjuuy1PUgMr2Y37D0SGBmGPBU1vx0gs5OyXPT7ZzJDZuPGfi0i8LmU95Y/3SsJWyMRlan
cm3SoxKkVCtEHLO/TJyiE5v1jVoM9B+AYrYPYZ+EeOoXN4+T92VQsfhp8xL0BncveQz0JVQDMlRG
Sl/kFuQ2KA6Pi3GYzOr0PxsONN0eDOROQpcCoNTLhArxiHXm86mw9ih/K+LH6NvAIQ3W1vQWEgAQ
4PBwJtp/ugfU9+myoRcolT9w7EwdxvbuQ7rQ4Bh8mszPjpYox0lQ0oECSTU2PJjSlMebb68OdYuX
WOFh+XhhhXnZPyZ9TvVMpxJ2k9uulB4ZTL+0SHVOcfcNikzhdituw3PqtOD2edZOsADK2tIpf6rR
hhbl+6ApKVLwArm2H0Aj8JDtcVst31MjfiqXj3c1OIYHl7cLX/GRyufOJPawA4zLeFnEDJKSNcm3
S7YU8UrlG+2SVz64j2M+VSuaj/e9xe9isqN67OBKivxm0tc4OECJVdTAMVYhjg2A67T5p4RoZcvX
hwbBaOaOU5Ldextq1GL6QJ59ElM1YiZtAJD82PzyYeW7ph3XZ5gK71GZxOjIA8s/gRw/dR+YGr29
GhVfKT4HxaslEfeswAkXJul4W/8nVKcHTaf+XDIocOQhTadIM7Lmvl2kNYxavVDbwnPShcnbKD7j
Uez3pLn90VyYq4MYTso53x6zR6qsLm1jCaMnwRyF6cYWdXr9aVFFX/60gBW37H4oBgCPFJsndxmi
oqI4DTmAMUvxy4lbtOW2F5AjnGBmAKCPthD2Opv4/7ABAhAIRZfaF1I80fKrp9+XSEVF3VKssbp2
Ex7kSoq/nJRt5ex4DWT+j8BmcwaGC8ZCWrA3rzjkPSV6b2ozfnU9yxUtrAdFSJd3vPu13kLB/H7P
cJzrgHN2KG6rvTcAYCuuoBlzz5/hCjmZ9NMyccc8tAcRCJNePt5vaOjDN8nn29rR12/A0bCrZqwd
hf/Lyefb92CLx/EOdIJiY1yuESk5L7MTVEm05uJ+T6HHMA7ruO2sm7pFGlQVyqAqtsk8uoxfdatk
BogI8haN7ua4FAukRGBma2FgRcWuOUkOSzuo28ERhDYVmuxomdsg/cPag8++wzSW3vLo+tSFz5QY
9GXgp11I9z8mzwEid/9OcwTVKVtndWAAiHdT/DaccqhGLuI1Iz5InuaDy3ZJhiFxOjk76Qwn/tWJ
RpuFOv335dK6PO4Mk+fAQf85Vw4PXSrkXcMeYJCsFD5QT4eL9qCZ78yoNygiDcjWL+icnRbo/9WU
rIWj+C8OF2xwE1HVal8O1ia/3LCyar02UGqX7QV306ozDAXMiAnGyWwM7QB4oGdOi8KqNrIsKiK1
6YE5dt7mBev+mw4uaahlJ6x6Q3QhSCSMDIQvylOoEDWVltd7/cQZXOJEWMOMmODwEa5XoydxgxgH
qsETxD2dZVb3QxvQRSziUCc55Cqp/k8v5YMikTzsz1+gIPJYJ92lCKm/f8GXDcr6sGr+TSzgden1
P2C8Wfxv9UX6KYKNm7TtLhZvHQu0l6LOYLK7Mbet4wT7qvZAZDT0wl59A1K/398zyJsflia7MHuo
RBw7Qh61YN3XFV+eXbcdyLeqdVFEF9uxZgt39qfMIgxwedNWISNPCyzoU0BDJ2OR/SRtRLVA4xqt
GTfCHUjBFVNJHTPuO4KUxm8sCJQPCbzJ1omhY97SPXN9IbLl8UAsucT320yGemOUAapowmPJuDsy
lgidDnGggTH6Ambr6WB0+RIlZap+NzPM42By8e0C7131zeIt8tRlDNX4Ib2CQmqlIS4T0LgjaURM
pbDWIGoGCG29RL5YzdkiXlaAyQjLqUWG/nI5ocQVQ0GRavO5yn1O6Py22jKp7SSOJEfFbVm3IUnk
AZKB9dT7mdvM0k/qi2WjkQ+VxqMA2aGNbHoA7a5w287/+DeFuH/dg1rg7keLQPukwo79+GXAasLc
t3Y4gh+p/kanBoyHFanRqC1QS+pE/C6luebbydkZYibIh1QNxXi+qCfo+F/uoSgHaUFun8zOpNru
T3O/1jURuV6tumLA1sxZh49VfQ2qcFl21GbcyR/qr+aKWZNnWfCAGaUxH9Buwy+QYxxhv/CVMbyX
2TaEbeBoQLweF96WcQXq7KSLhbnEQHn95604RT6KC5XV0+2+zI6QyNI8GxwK5JWy2iyRklMA4lyc
Dqadl86d99vQs4zZwmz+kmzr2KTvY07LUh/ORN86jGE7ZldxmQjAv7vhkQlwhWghfiehjRJMJmZI
IuBYuWGcr02B02TF/gDXVK156EhAkWMZFMHqGDMA3hQKTSWv7WwYoYdwxPAS35nS5cfdxXppJtJ/
quwCPlTDHp3OT6WeyebntRCj39WPmOIOrwxYKP2edvpQJOuTWIV/ZX+/f0SmmQxU3srDaZnQZlsH
oS+FAwQl3rEvH0e2Nq3/uxZF8+fc6udJjLtgm/KQVPNAhlpqB/gLLm7y6SGVPwSHD/nFWynUshQt
gbTVwqCb5inPrB/RBhVrrpZVsA3SrtZqc+B/0b3Yk8xxLj1EvwXuybHAoyRJNFDEhdKriawHr0M/
lVYRQfPqet83wxgoGeXoaEHnOi/f7PX7aPEogJcf1CEERTwJfzQa6s8GJWiJ2vH+Fp3+vVZpBX8f
YLO7ISLq/jc7iZRESDzMJ9K2kKhKe3G78PE8q+cd2YBNKt+fr2rDc8TY1Wxp/2Lf9UP6VRL6ikvc
T5MAP0tULHabuFlReeUH3hW+QH3HLJmRy3hIlQEvBlyHTRQdIldSmmPwGHXs9Uy4EaYrjk/yrZue
ROeGMKsqO8yQNPPvzB6PE8TVLQzC9NAso7iqu9tTmUxElkeyhVA3P7vKqpDvu8KmIza7j7aYk1G1
lhZuVFJheSpaV6bPSXjFrhDr3IRzFmA7tiOOv1tuGXLYP6Denp3JqPPEjPqRMDjz43wk85z6Nx4q
yGm8HwpeojuIKUKqe9boyC0Rmn+SzEIFszy0Pw0ds6PbKToJeP23/pIO5oFyrZd2zItfTuZZBcTn
xr6Tw5F9A01DXnqG4h08dAb9qLzinXQ+kBCpT1nXspo4BCyDWSZ4AyfYy/h2NchtJ7RydIw60uaJ
1yzBW8MNgpG5jB+r1tRRdrOi/phEOC1n/wkvJLjlWI64MWpmUkD1hI/ZkcvDKWoifsQP2GCRaUmx
nAWeC3WVEcZp73maj58i1LCCS0XesW4okTBo5bV1Yd4xpXjzDPXJUh4VLjxuChkBmTSJdMFs6roG
mSd/OAhBtpMTFz90V6RYwH0JwSAW4nQ5n78k7P6562ibB0Lbb6BeZfNkr/x6JnxasAfhCU3O7l6j
di9OgGxrV0POyDFT5vJ6y2pAPEaPN9v1V3rtg6Wj7agsGGvqdQMidXNyR4j3sFJl1QB67CrXhO6C
LM/UuheKO0frwrp7kCuEORL26EXoem7quGKNlmBYrhCqB68btSqlyc8E118VATTxG92/msMNuJcv
BGJO5qMgLJyBqXw5c+6k+8CyRFlO+PwCzp2nxLUdQs1HctekMAunn+Xd8FNtulumX4/X6bkW51w3
ndOXGP3Wa44wzld5VrDRQx9BXnBE4z9mhCEBNpjMHKU61PNHBe8V6J7pyROy1922CwGCmc3eZ8hO
7ciBfHu5enN9sOqEPJaM1EUzg2dg2NKtzPTfNwI7AZacqBsY4AgJOyK+EQhE7417X3xCOSdfjQ+7
SYyDMgcL0XdSHmXoGurWaOPpsHKTSZRhNu89af1d1onJJQdCxLleCHJmHmhQbAsgGW+VxTCatd1q
NIt1UJF5U2DwqrSIq03BEyPiNuSvvCa9/OFSywtZsBgjSJE98YQLlI+AtfUtRR8Uent/iQGCdt+p
kEBXqm+T5zQsioJ2mLzSLGZfPz4VjYxn1Hv09EAV8Qbi7dyUCeJe1FP4we/cJZWw5BltjdleMGDn
Z3dNyR/dDaoopKJATM83SFOTqZ8Xy9m1ncbTt01z2OkRNmmWg+R4sOaVS7WLxBj9DglcNBFGexS7
otwJtziyb6XAMq62AlNVApDqcp94qPvFKJRSKD3G4h0/1Z0MYVqXp3Sce1NXzzler86V4RC4h3gU
q34KMmM6pNk/L/R16EacFY/clLEamadY5QJDK4DEu/KjJev6OCG++Qzt9a0oJ/+H1gidnCRa+7lN
TXQbXOzEEY8UcM/PZOQNBFRAMVkwUIsSVpbl6Pd9URYwOmxWbLRwciR0iUqkTDvuQ/+a0zoTtPvv
BN29HdaOtNeFuYvUa/KJ9UaV52rpM5hcZyOY7AmLg3X/2ZpX53o7WSXSzWUNT4y7DiS7Yi6gcASP
NhDcjqu88kiN15s/hTGvXgiycID1XjUhsEm1DvNG6i/hyfsQRI/gSgm28F3roUTWV+sY5IPmSKqT
FAFyviQY8ADqsGCre8qobL37nAXgDSP5lnJMUzsZ4C2rdJ0MvAoLWtVsNRxEAd/JrzuBO1zJWsXm
PU0XnXb7GUytmkoLGYrekv9oYas7EsMxEngOR92qOBUodSSVPMCu/V23FKvWnjhJXK4glN0oVFi5
Lpsw0Y+AVAlkA+3S5nF5R8PWn3Z84P+jBFn0PVhrI4H+KJ0u4B+Cab6Y4rZ+fjn/tYWNFwnnIf4P
LmUc4ENRvIKvrCWrSUnXgt4UV12bE6+CgneQn42a6q2dfBYvyRMrdl1vpyID/tkUio68mWnW/Hyn
VrmRi1yVrp9K3+8X3yUJyzZ5TB2J/ZQ37Ln+xLNTVyIvfSHAblU/3r9A49q9nhUfBcVicb/uBOaR
YhfXs7rKSEBKHlxQ8btRqtgEEwjKGe1YC8WwyNgV6yGa6IZRIoXKtT80K83rSnFw1lFCPqejH/BO
+5smh+5bveMMBJRiO0dOgGSwTA+XY3jT4oIk/5EKwl/jCqkwQLwKNOWG6Ro/h+XRZpEZ3lyv2tkC
y9O2Yed5BFiTMbrc7JYLVc009u3e/aqRrRUJMmJPVB5ig9O9J/T8mprwQiQsgPRqqt0tYx1O/mLZ
Cww/rTaXKtkiKXGF5QGBGtD7e3q7/6QunqpB8zIUySuKfYtDdhAVCBqZ4or3q9MYlof8tECDqEOg
89JSgwPdLz+Gg0+7A+HvQGkCn2+9HVYQEdRjC9GUh2SFqFwUc2nPSPMkDudqJDpVY8Sv4DCD65eS
mBsQdlmhzn/Dswx+/OkVN7XJxhTtmO7V7L8WsBW0pc+es0JS2GgMF5AKXYp5PTDfqw7BVbXPrwaA
sle/nOi8BhIY3ysBiaf1nx98W3u9gxPHUYdKI1s0Sb/qOQbwpK6VtM8GgQfujErOdYTwNnSlR0f9
9BQQhiDnXFJjn5W4HRMqzKHZzo2lq+M6xR8JjSi0wUu+20YMF6UaQXudoWkp+1Z8/rl8spe9m4s/
XY2+7D51NZD9EF/Dnzps3jI6MramVn5/N7xsRAVTaFyXMSe+97PJjPu93XeliljV6Uz1IZrBsZBe
2yxY2JYQ1Kc8oAhVq0tTZNLKSdxK862g3RosXROOzJa/MAuEnNSx9LirTL9GJXrfronIZY/ldFui
J3yvlSPB7ut/coc5jOQLNAqK5bi4lpe/s8fwodjK/Tvw9Am+xHrKUiDk7pxdf3Tg0h+BmOu3FjKE
n4ZP9/VD/P8W8jh7GuJ3S+R3PQu7Lv8+lGsj+V3MjveXfg64XDa2JATNAY2nn7FFFtTh3V8nVrUF
cR66ldmeLWhUYtvYqMkYyEFuCTj8PaXwQu0WHSbD64G2ej1cSHtcHKtStJQs3RY1BYuKevOaYrIW
MuKGq2B7xvX6BLI5lJn5He8EAqeDHzmsR8JSwKklpV+hi5qbBpEnVXHrEfnQWZQ2nY0LjJSEQFy6
kMdpUHUWts56IiA/M5LG1NT1f3jRo7GvHd9xGRabSHdERYWqOgANtSU36Z/smC86OlHrZyAYtrQE
E/RVaUVwDVjQAWO58PHyPRpHYMMOzhZ8gyQ0BYvD3nhWbzNsGRUbjWYVURBQTsI8smVscrZ5CZg3
KsbqxLLU73K8RigyHw9Hf5ogo7xwLjJ/TB+uiQKRMtDiliyrZZOCMlBj8JPjC50czYaFqzYrx5G1
n0NUYuvhuFdYVKwbFdMPDR0zigs7fQ/Y3qgL+xxUfroksD6ye7dExbDj9eIGhmLncmYgGr43NvPx
Jm14xaNAXiw2QO8Z0/22k8tkAgXn1VuGFL9CT/JDms9teof4Kd6IicSQavh1pCr5S8TXKkBWKPXh
HnU4n0cKmn0fp7a9N1jc+8vCOIJxjiUQjy1aTmzoT9//qvg0Ds/b8pIG/DUlsxJxjajtc2wCN9TK
90nLwQmUedhaYrXkBReExJvTO7NLub3wSWAbfkwMu+YebuJZp3bp6GPeL3bcnG/c0oH1U0TsmH2Y
fXXxP02CzHioY230ST5HjVwbUI6v6gmUA++Hyn9YgRn6Er42iE+oHCeY+4jJopgNhQoRFpw+8fbH
gW2h5Sq/cyHEO4H0p0KDgnKAn+2bpPLTlNv86s7y5xdqxZStvccZGSivHdQHGxi1wL7Rz2ZsguKW
t+0TtxO4SAFIp+48q3K8RqvSLuaFbPmSJM/06tmQJU4hgpNMX/bBSHSSm5KpwnEq29COsSOioz4D
plZW6CrNh6vzGQukJEi/rDCAT70wcm5zLIjbMVl590nUtyAZu1DeOA+6vY2VvYOXRWjE/93MtMbA
xZI86ISUn1594XpAJo1SuATeP3BfESVrBXL4Nxi56+Oc2/6yBEYBRJvIYYTrPkkDkXFXYm9PxlfT
msiTXSUqaP0wv8PF4/ejHHTBn3BtoMSw/g5qRfw+Af9fSZRyvA0r5F+bVvELH/KTpDNaLu3wNPvS
4stFSA5tHhuUROWOgk1TBBFv/Il5zqv4NOWV3G53o3FU8WAAv479f0qoYTpLkFHwCvntvDoXSRaJ
KGpC8/HutNOC3rSVtH55y43ZOMUQrw8izMWZtv4uWUZsZqHjw4zF8ArHPZ8Pd+rnRy+EckFw6E6b
4vxrVv7bJvmSnTticGVGO0h66SKUaJnZKOqaFZ2mIRQBoAKGJWZdI8phJ03ZhM4JdZOU6iId9pGe
vyzHMKlCbeCpAdwAOjZqSseOddmuws49pC1jkfGrWsgXAriuWUWd+7Wcad3O50ILlKvJDvZMjmEC
DkDVcR81Lx7C9V3Fx/Ip9Da/evCRy+PzkNm9AywLkZ42pG6eDDzldD7Ou27nSyzbWV6WzAtJzRE4
s+sa204Fa1MK6mATOHZRNL15WQAtHwqXRjGZXEKiODbcQcfc/LprJdzYoB+bSMbYjtYcrkfleeV/
Hpf823eNrdvZh3Tekblwix9o9I+Ovp3liaUMpi8jzBjV/6IeItGRD91u6IEvDBRfjIse8S9JRp9K
Pu5AaYB9Mn8tY9MvDXN76gGdTo211MayamXm/Jvr/Te98IUEsCJkFmpq5dYc8atEj1JjFsN26Ag7
840gskVQqnGTBp2wFZAjVRBJBtsPMTDeA+uXJLZgukCH91qww/UC1o0ktFfFhhdKG4tktZCmRyUd
PZfF+zorhy3Bb22wLfAVxsX8f4d6ruP35VJJHe3xBk0uSuBhru21wXWYHxc0wpsNljqv1BqsdiZy
p7sksCaQfOObs7jUMDKyEd8KQz5cMahpcYsEC8csl8g0P2s4VLd0PJKRWI9IvxvRQhc97jQjbKC+
48gjoq+65KnaPMvqv+WAfEn6d6C660Gz9N2jzo03tSrB8BQwHJamO/A78YW9qyHwLVSH5pUxGMn1
s/bqQHjzjsfR0Y3NCKGPqvSXx1X3BBkiNMm2Jty/w2P7xKjWPIwZjV7Gv1H5ynsKdQXRxR+2v57K
ukcRjB5WwwNB5ScfIOveU7m7MN8bt1k3u+E0zR/SNrVg/dtxYwf7zuMCyRHXEksy53JCI2pRXZGa
NfG50OpOwGwHG9PMJbp1s7WhOv27nAMvscg2sXjLinSgbdmC8sem9dXGEUteoWStY9AG0k8C7hI8
/pyFQjSZ86xlz6rGWZEb+fk514YKCajRZw36htSMw/fprsHCkjIB3frgh7oef8+IyAtzAgiCdORz
tNKqVTy2Q9lKvNJUMs8Ec5O9Uf5XmrUnCr2Ya2I3D7o08rZNHcEO3kSm+2k19sM/0MyoPB3Xkd0d
DLjsr2cZH7JGqFdvHwQzmw7/wEpVcJXv2bJpz01aghbLlkTD5YVhZjCDFk4GM8wLs7aGhi0tozzZ
YKbnZ90o9XLzd0tc5XHEE1edbYLSqDi69iT6+wPsZO8fwDC3YIh7tZzpwGJPZY89ZO8Hwt8+i3B/
6Cth1rjhYVLRHa8iXmlURo6K/2sbSOjM2b9+pDvD0UTRkxqhYyI22SpMKdRoiPhjPmpkK8+CayvD
PcV0w4OeMcGMjk5erdrCSNb/8IEUh5w0sPhhxQOYPcC8sQt2X2v7ERDXHMRtX5/dgLIO6fOgAo/P
vGMqwNHrrZwymD165MJNYIWfpiPggLqTw07b13bq9KewD5Eq9C1zG/HWkSzH9QAAgpMH/hoTc4hR
rTlfIIpAYi5GWWJnqTSEl9325tg11rFVZZlm1kLJ8afxO28ZucgEpFCGgZ6jIfhP121x+vzWhncu
wOjr4SyeEt66pryutxAJsJPRCg6fy5riJu9WLTM0g/5Cjy8IlX5T5wRgu73TsQkUDRkLd1Vty9G9
nvTn0DF/9oqdh+ZArOVX2V3M1N4CoK3+tbXlCvHvJW1oWLV6zYDh6Fr6oATLVR1THi3ICh0q8Hez
K4Q7o/HTi5YAOKKI5chCgxW2oEfZWqJYhBVuTF5dv3ybynOjyi8wNLm8Vr5ts4DPYlR5drWtEtBH
mAX9zlgOYvY0Ik04TYOV/hF6SpAeirWeVV1N4X7v9fXipl57uHZW5/bVT/JG7RlqcjxgzkrPTHLo
CR5Yenlqf5KhqcziH1fYa6iUuGP2WB881BtJx2dGmvRoRfB4Zyvdp5fdGe0EABRAe7oNLmRw6Zmo
TyPP6lSv/ApxcJpuN1NQEJCp3gcnYCpD/PZoXp03THqtQ+p8vT6dqpo8QD8RadxMnMj9JQrZ4/Sf
YtbsJovoOo+znngh0CLFoZLgIoMZStWD9UZNvvt6TTe1zbOOnWosmvGPscazGFrUkWW0L3lnbvKO
UHbjpn+B5F3EmO05CoV0j2MT8LEqIsloJmGx2v4/1S/czATfmR2qUCcxO56H+fhFi7a2go/kvcVn
Fu1oGWVDQdproyQfNnmU4AMF11z3UbNcz43amxY00qqHLOx4jL+mkBo7NvL13QgOvq6LX4tk+o8Q
LCfG6TphnvwLII1bknanv/4/1VwgsC4Mj2IX4Ueml7gsLNUC2mLQsjKn7AM5hK1ekZxn3csr41/K
1HyJWfKvZa9uRC1HJJemAjSF5L+C48kQWBcu5bMn2uVchJXa2sTUMIliy6JBsi9uFSVNbqjQ1dgf
oiPh5kcbH76gAD0kfN0EQrlXEE0YLIOOpUaZWH6UKawNocgoN1PXBE8nw/paskO40vW4viOCirDU
djafT11UlFA/m+PNXT+eXxa6s4l+tUzTP9lF1np+YZPpkZvkT1WieLKn2ZE9D2ytmN7X8ihIZGRk
nnu1xNuDZ4WiuUe9UvSz5Ui3ZQOf+a+1j0sPcxqO9RAunQYeDbZkVAGAry/gTb3qYgR04MP/4OA7
IrfhXV5usZAdDsh0s294lp9KfQwCR0Cc0Cs1kb2TmGxdkDfK0hqmZYbE3vKaRMCdDJSlfej7qFrU
yzMTrt4q98jDlJktqbw6UP/zZo1DIcXqEG7EIeex0tt+hqJ1tc+8GoW2EnBg+6+4YyFsgNUPvAdQ
OR+VEbiFiD+Ma9iWEWHJgPnl0i5AtyWY7SCfN+IwcbRnURPQQ8ZHQDiCyUua5KCXbLJKVCK4qp81
TtmLyiemiJJWT+Z/slbvJE8ydDEqjmO148RzfyFrQr2t3m6wnxDllXbYofCvy3dqden8mab4ySK+
XNN3XvZcGErMMLMWI2Sv3JUeKIwlNPTk3UcNdUWYL7KQVqu1/8JhZKrNYwGNoeMtZWhb3QOnUI91
Mxdil0gnV3lBiv7Qbxoug7Myq2JteTqClKgXkCPlF72f6QdQQyZW2UFBNNvhlw6M1AoSpjBzZLHD
HD2pQ8KW9u+hYDn5nptqE/vdG1u9Fmqw1nQY2Uswmr2IFuZbp8E3kkghDmCo7Kn2D+bY0ux8v08b
tG3O+xCEGrQYAe0zDvyRPh98VAuffhNOgCFE5L98XGydFarrRY+OYUf5mFnvdCn544Frl96J4pke
uV53Z/14mB3356NLb294sFkemm7MBmT18jmNsN+EasR/OtKIzXi8eEPS9v8RU2xb+sYnKjSbcIhe
3brYSbmyTGREMWfYja+yNJOVaRwgR42+ceiUsQ7ZHH/4mgTzC5a2NGg1oWf2kYAP6rPUNo86ZiSk
ku4kuNFWvxlMH/PcaXYaf4ngH3lc5EXZcQTxaDxwwr9/WAlPffgH2xxceJAqj6Q3J5HgEyQNDZ+X
yeKWoOZl7O/0JrPQi0b6JOQ5s/9Ap6fcMLlKQlWWduhSwqD4Lf/xcckDUf00jJEeXx+E4NAwMR/1
U56yoTeZc84aJ/nL8bAW+2xl1XR5/wuMtm8/W/ZVolRISUT7Jz7/f1kc1TxMNcfYOLu0SOVtxbuK
NOp1gOSv3U8A8uC9SXYLLeE8zCKSG3nlC7dz70SURCSTEEmKrXxg9P5jgAVgXjEqnIObxnEAoQGO
ebOZoyyg5/XEq8ih5vZVyaxd0q4G16jlJuDoDHyuIEqBL8tm0sidWhfOIGtt8LP3NIESITqMezCL
FfstKpZCfcPOWgM23+czWJFZJVyfJUk3GIWjCzEjwBvVl/a9a5pDZHcjp5AAeG45/yWkThqxvQnR
Icz2qbISUcznf6+sKiIlvueSWSoOfPbdNtckk59Iltjd6gtcCpZz7v2plLaxSAUF8ODX2TfMyMOJ
/9ScgjXBm+a9LKNa1iMNahPI5D0lIBk+DS2rfZ4Y1Jlb/HMhSZ85TgREof0Gv0TvVkJgTqLK7qV+
YEywkHPyA8f2nBtzrSaulw52bnlxTqwBa1lg5xN1DzP5bfloHsb14eEd6urzLJX9J+wPLh8cPjok
OasHAGso5un3c3nBO7hfkVv+MkRJyk0tIJhARmFjmYeAwBw8Pr6lnNkzlpYqGNSBZ7fVA8pi5krN
DvnLP0CnM1u6kxP8hN3CdLhL05zKzYPiVV8W8pFPf8hG5IDWJwX/VH1+Dws2TT9fKqsO9w/qLDKZ
oBQvl0E5umRPuJIsaHXveV6mt6FL/0cvGp1JF3qcZl8YM0n6OqwVsOfpNGKmex+sm6ybWKZ+r0LL
ychJAEZdX2JLj2y1Pq40VN2Lk/4zlyzsOINXMun07Nwurzx8Emf9CSDuqBoAFa2aPdoEPD7IYKkn
XTdUhep+oPbb+rsAT1clxsayN/Af1PSZjd//NRWDvqxTDEEdbaP30ePRyE6pg7Hd1RfryywgpEWP
hQzzE6SSz4KpYGPg2nU3HhDnO1uRiToPk1tU5iOYgzWc0iJHQ2xs7gLEl/5b6GrR4zBvlKmB3TM9
2ksS9TvQ5VRYTKsWdWwKXTl7jgqikc634TounPBdqv66thOFzOCV5xVGh5ymnCm+fSeKWWGqX4n1
DE2Nc4WXDbRy0mKOUa9Mjo6OY0svcJjzf0eN1gThxN2rfpHcXZNsWDh8Zc8HZsF90A+7wJ1AqzIZ
kIeC0hb+FOilByTwRRUyecSCO3JhU49q6kc62xmtti8lVxfEPPnmCjMvr2E42QxKJiZ5xCbM5fTe
4nDTwjbyod17BPz/f6pYKs2F+SqhOxfDPR/WNveq3Q+fs6HlyczNNurodQQOSbWr3qvzx4zggZvf
FqU1HPqSVSQId0UYWta4yDbEIh1W/JjypWgtW0v2nuw+GHAERFUE297fsHe7fQVGPUE6zDFe4+d7
OS/rYes9Fu7medInGfun1JmVUT1ZcvtKJLZ3sBncD+R/vfUgZC2bO5tdhg2+8514ztMzlq5C94sO
xZ3NmXEDbLrHXJhJBs1FIFWmUJZnLq497MSxAyr0Le1tZAFoWYVALxO9byfJVb4+M2fbY7Uh2ZQz
Png/bPIKQCEt24iWQZw/NZazc9wlt5CYELgZzKV7bJbLMUIq9jem/RIzjDyIVQT4emrcW3eSKkmJ
2J//sWg/CZ24Vc41yoRwUOa2XuYgxYLOXQx5+YvArLuxvdtA6cTCd33qMlDgk4r52J0qT8Jd4bkJ
zG02sEOu7eSvqmWj3aiXpny7jEAnACjBMk13V5Y9vvANHiGVrOaO0xPhpHIQ+hAxp3o6DzIsotni
GunZAr0vMttyCbrV47sHUso93KBBKbdsDgr5nLD5ecU3Cw2veg2UnxL8dw3Z9lPbkplhDvF+F2zY
NqBLqTonGb8jT4OImNLTCcv6ZDhtMNNaualKVdj+LNWievs2y4q6NPnw5HFaEYLIB2SnWqc5ya3w
3neMrBPaupAe8L4J9CcUwVSl7EGbW3Q8QXWtMXziRR6X3XsNp5CSWUHlI/QnFLSMxVYgdqWB1srg
GCpIHU53DEbpuXAmquJXNZhdpG7i2iZr1xoJArbJwUTfuva/jPDCe6E5+s9tmv2ch2DQkTvhoJbG
R5O8AFBZ5L9ax3ryddM8LgQ7fQmHjjJ8ubANs0wL/nCXGlfAGyXR/uvEnld9vFusMIn7tTekGujn
ipjZNYZcrAvEItlpZ7tGUpKO5XeP9MiIaAnd6cX7RPOS74NvAN0q4sfITGbgIhvs96G9lTXzT47G
++LIYkuvdZuTMmRMr3MVVorYUVeY2HU7WuUbv16eBhFv45CGSDta58GjIEvScR5M3UN1pz6Io85o
waJ6w3jm8LREXdvFys7Lh1QjFamvOWOArfw6WfUgV5AQfwXCAurLJOqXBlI6hAnYfa187Q7WjpNg
X7ZWvtk8WkBviNeK5FSJsGoquwxlQbpiM3Po+N0ePocgRzamXCLaZY3COi+1mIJ3Pl5EoP9Bcrzh
TQsmuYqAo5exyll5R4GCKUcP4PF0qnko3+9LhCOe03zkul4lvdlM5iG6OtIUroGEYEifTXhIvg53
W2kGzp6FX/jANYRf5M9KpkwWtY2+nvwfP78Z0ykK7izs+BUXUE552HqE+CG2qadgQ55vSvBpwLYf
fbo1jhhsvdQViZElpA3AUStw19aPn/cJWOHXssr82GQ6KqPf6UyPRpaUedb6H5cm57PTfJWmyliG
2g/cTFthoPN3phv5yiiXQcO40l807dPFSb5fLx9U/QYkHqA5btGmjXj2clda0UZSTgb/iYBTHTVK
uelc2UwPXPjcO96ifwRLAfJcs0eI0nxcGXXnlkFOOVHhoooA0OJxOkBZcP2StXUhIll2MJHZHEUE
EJmfYs4Pt+JecXKcOQbJNsDwzAlKWxyhrKPZUW8ItjnUBuokARESWdfA4XV5sdbJImUUbUj4xvaX
TkQtlebf/4wQWdfk3JCuIakbuUG3VpVDmWIUlXjOIdIir9Qo9qxR7bFu1zcFYwevcb1BI6YtQw8K
ABiu7esNijqObsDXBmafXViS7/vsqgkZuxM0PDwg74RfLHcGFPBTomd2KiAVnFoGb9zYNbYM6pq5
C+LJRrlFlFyB4XUbVTlfGqdadvCaacUx2fso3zSKAXN9y+X849AH6XAJfUZwaoJqQlXlEBe3ZpQ2
HZTknSkE2IO29C45UGBugsL/8PjJlu3TLBVL7SPddc6iLasec4m/7QSV43T0GwVE0SKZghYbxdSj
QscReA8hFQxaIBlaO30B1pAWIwbKZ6q8wTXSrfPX1e03mxSs8t0jJ/4n0S3zjl9UqIIQWPnQgZ0c
cBgtPL9qWXWEhnIq+AH/QmM+moGE1aAdJfZtt73/nIwxhGkyyq4et7IH+volSexqv8JDwPEfuRhG
AzWfmt0eyMZdsr+lYR04bdTaEcbWZfJRY23onTg5Z5hrF9dqkG3VUj7CbyhEU4zZbHNjwRJgfmCZ
HQC+0TxJd+jvHTT+R7vLJQpdz1Oyqn0Aq5CIen9hRBQLyB2e6fcWbLhffAfBYHFEDNfvEAxr4gon
oRyqq1b8lD79XXs8+tVAvCexa8FAybquNtGl1iO6w3VJYaK6Iju/htGRVq55a0VSzIlhWBqfJKib
CX1JhZoC0JcmWPIDWfMgSpNhaYmorISdGaTeF0dOfWFXf/9qeoxFHce3a4mxSWpLH1ypsb+r8eFx
798CtuaHoLaNdH0mJtm100nkt0RBQ9oHqBQ69XVz7irBwl7ZB7mZ0GLlyaYhj33niVgqoVhhWP89
agQa65e1xWjuHNaag78vMTBoRJNmiuBkBhvtdVMEZaVhu1MrkuRAe/nGPKRe81Gfk4nxWedK31hs
AkeRXOPkoZJAbMF7fIzUqVsnz5H9fbG6DCSwGNzqwreYfQykUyvroBzHZABYYMdDE1/AazcvEqUE
YvIGxAxL30rmu8nh0+FTGLDS4sdAwKqZ2ytTIkH0OWCULSGZOLdeHgeuSYqTr3toXN2CAl65AmCG
unXhKAWxso+EW11E2seHnbsCJO5WlBTrIcGhKCayXqc4v1lgh/19LvExpIw2EjNeMZntl8AAonI0
J2I5cnlL8pfComM3Su3Qv185YC11FdpnZ5qkf6Mwj9UVtd6RSaLjcfrMvCD7tJmnHoB8Ng/hP8dA
wTRnaTaelA3q9O+89EtOBxMBRxhcniACrn72gfSer4SKPP70HxxjYVTrkaerJRbMTAERkCQdiwMk
ugL1ZHd6oqpAkXE3/l1kmUn/RpMB4yE4AhVPhV45QQK6QdBO3iZzuntqewBjMytdg64zUSTPA/LB
uMKK9SWbf8qEwR5IF50LM8BxTS95y1UNZBE8QwXS5+3N5lktqt07T1Gr/kNc0YgyPFXyXWFTnD94
3BBwilaBANo6IVStHtUe7rg9U3U5sv686/kHjey3ZAR5lbBY7dC8yToB9mMFXpt2cJFaz162IIaD
vfXXfGYbpA0nrzLbibIq9SVHuVDrf2ip2LMjoRt3UT08SXp/B/I0X0UtXCQAMia+TuCJNdZVHGgs
kfW8wTCLxgjAN6vDNjaTZ7Vh5g/3N709VY/uD/JwTr7+wu1KO5XFVtTiDAx5Irj81lxhnluY6Be4
vZfDntxDP6/g7NdwqXC/CDfrMe3EFpDnl0V2qe7xnDC0pt+MTGJJ43Hr6VXLmCHFy5swtdEIwD1U
nN0mPDwpqZhk8tVwF4GxTFKc0Ebi0m0GvLsUazMFTrU5hlYn6r1u9HWge8UISIDQ5r1HUSTd3gsL
KiWJa1SsoLkx8DpvGExv4jdR3CSkdbaeaEGq3cF9ZiRV+fEbVJY4jiAxqXQ5HGmifJ3A8j9mcEkp
1i0AhudZgpre1mjiRSUuew67djWlwo9SI2MwB/07l4nbiluV+mP+UOLLUZ7la4TNMbQYit6am26T
7hpM2IhoE/7ycQYkrbDx8rggRnYKHkimHU1WvZIv/nDyvCt+q1n05YW+eZSiAut1kP/hWHIFPjD2
dN1pUdBVKVoGwpL/VaUSFg6gFpQaPDXHJjM1ISh7mooO7bGKq5f+CEF1VDV1YKCbfHT/54hn3uhC
RE+Q/xQSuW646FP9EroXwY4O+n9LNrriMwNF0JofT4pU7PQNrRdeOZuIm9X4pA6TELGAF3xsN5Bu
UseUYBSRI0UNKoMMKYYlbjNKitW4GBCi2n2XnhrQX+7mOPi5JTFLHHWGxNw2oOSccp6noGUFWyG6
tbPRAYgf7UJVQLaO0pOzwwSgtgbscm5k2wLcL4SrlLMgzPEMDWlNPUHmErfA0uCuOaPEmBNShoGv
9b21E+sBjVsYv33KO0IaAJ9ZiYNeCup6i1+rn+H6ahE88J39QoYD+yPvNsMT9G6jQZTsop5vmRS7
Wpd++ZLtTWTReuh3tMfBjzPt0LjfcAJpTnrM3duw63blS/BPABzslWKUV6Eno/RtWE07NacyFgqO
Hkp7wVOsklpOYbdjfn8FoWi/vx2hUuSmCkViAMaci08tXRzMS0k/C8bavbNyMRH3nQRl/y/NdG80
uAiAUA1lxl711ZpEz0hxrb1PY5Dr/MtW+3kb1pjRRzAEIQceswNySKry2gnb5KHNzrkM3JyZfpka
qcaJ606dATJea332nEzNCjK+k7QdbodVEHJ5gX4UR8KR0YFgJh32Z4PpwPgdfM9t0WiqgjgZlZ4j
juKVvHQeVAT4DGfMVtFekIE433+IBKPTbjvJCJcmTKkx5i62M8bxlgxeJDOod7/h5pJfjXSe5VSK
JZw8bzPfhlowZKNbqIQ/4fhkBx7Vw1qSRuznagRoxPYJC9KJF+OPcQG6FeN1yUpZjPyPmTeM6uk3
Wc5B6no/3w4EMHAwzPEnk/qf5KdlXVqcwbDb8rtEpeXXMErbpQSdo9ATO4d/eHtZkeo/nFdS6kCk
hSDQVf3F+SYYVzyvIYDa2hwrqZx6P+NlRImPEbA+iQH5sSQkU8yEVpJ4/Hof8MBsVR+/MLCEL/ji
Z8R/ylFB5VuN1mXoXmxYIOgwiOuvFugwJP5v0ljhU1D84t0VB9zGsD19Ulu55htM/Rga4gfuCeaf
DLdUqOby43Qp/Rl1pjCbDKa+uhfD/xCLMQOud53qVEr1ABXFCVlZCQv4Yg3z+8iQZb/OrpSjBeTh
13U7YaGPdXhOyE33lXfcn4i3mYUmcJ8emkG7TRcnHPu+66qcoWQLpkOPslQ0Sua5bvQX08XxcCam
TvxceQ0itAvMXDOfS6YkWsaFFdCKkuKDX6U8ON/ijIKIvwwIcvuNQGS4Wh2YMcqtepVzdfkibwUn
ZVTB3t5rzxdVWAB7Eca4kT2ViD7HKE+m9a7Sht9crwgy9W4vdwSp4HJhIGxHSIT9/to1HZMviR0T
TNKU1nXQyuTkMy5StwsORfqQC8lAfpRybByWSxLYgw1kIILUg9WwIUoHNo7ZF0MAylnntflxj99R
O8/hgbIM4wE4f6ApuoD1/dpDR5vYQC4txfdMHsM5WIdU+PL0VghZQVaTDJxP3XC5A8dnkAEyBVla
A7XhhWnXEP1I2Grr2aQKAo7XX0RtxwGVNWx1nN42m1zECqkeFxE8buENfggHjVLAC8x3q4znehBg
o/jX/FDQS5q7WPjOCbXrGM+c0948wD6d+hGoADBbpvgI5N0NfCELO/rSGCvmSjyUKmLcm1InUXZq
JtS+DXgrp2UdBpb0d40X0tK+Oc5haeMaR6OopmILChaL5muwOUntAcYYm/t7pi99TrwFFaTVhN5J
CZk9GtJP6eLFF/Ts42Zw/T95xm7RYPwex7/s4+EWooOnwmA/GWOXAlN1dIUbZbSC9NGcgduh9i/v
PnBF5TP1zZQCpFcqweLX+1gCpJw8EQZCMtbyVc5zMhDkGzi4RPYE4QzshKBu/5Bwl9iOktGAMj8W
/o7I3ERKx2vvX74wywcahLFywbMdpLmSmuOUbGZdCGjRQ30TCQJKG0ss7IJSDwaPZ8NDt/fLwQg9
x71RDWWhZEQSPkRs8vDex5lJVyUlaTQcBs5+GCdvrIO5PLhasNHOw/MEaH2kdg9wyfxYeruUpeSf
pTE51hKFZG1Giz5qNwBhrIMLI/PlHAz73QXsul3K8S/qjvotY+Buc3GiGoSQVQKnKqhdD2orRmw7
fQRkqK8GIYSIQ2WQE/Zv+/qsZGIL9RVyXiZNjl2xgsjfWurdVupVt09/N5omheAUnlGGzlPNlbXT
Nj3CS2sUgW0EEph7DUjIkkA/b5tMQ+odyrhUN5vx3g+R+6POAS9/IPGJhYHKSJQLTpWBIFqwkx1I
4wrBNpvZaFv1Y2KrwYEjTU6D6Tp3RzzHMJH+/IEDL1Nb0llXtRmxr9o3E5LLAzryMTPFBcvcg930
UlTg364d5oV5hg1xGhrMrfMqAvihcQk2uSsuL8E8KpwxXFOCJecqgwX6EZ3xI/HeX6lhG2ei24Tt
4WFW+XIN+BtD/PaG6wcpWtFDve9U+w/nDJ7uDO/JMCiJdchrqro+wYX2u6A9SrE/EJWPiaYgNn5r
RCc/rDMMLZLp3zQQakuTLEGBgLqFbQkRf5Xb0TjVtzIZuTpIqytWj23BWIwgUd3cs/3zfFX/0Drn
N63E7GWiQImS7AAllxrm3grQ2kkeTTSmCX8UToemrjK4N1tNWVzfd1CvosJPsQz+rnG6SWW057yK
aW+i++Jmrt3SdcLlqd+ClKvuQzrPM6SK+3Dk1Nvdm9aw/SsX9fzBsT5AwykPG2ydYNMvCjD8CvQK
JjdyhLQGxGD2h3+FXkXkuu0cqDmns70ZaTM03MID5mjqcVT9cah4Ep6GnJpray6vTdu3FYkKommw
s8hd4MkKwyKVwDMAXAPdH72Qbelqz80bVi2hIpxDLuQqCSjfvF4morBSS3KwygtjOtFIBjPo8W6p
O/sX8BxTXrI/pwf+CNmXpJSKE0G8pwX4MG6UKgF/w1bdoksYVQSvva9AaXn4aI/6ep/qBpKF7JAP
PS5m0si+QlG3LAgqnA4uuMDmFD8FMFOY+B2HHxW8ONN5gVbvu4l/yjHC6U7oKDzrbphrk86YwxYo
tgldJGBEsnwPcuW8XkS/+qdxQQK1c098qcYj2vqoloR035Ypp9SbNrnkniLdwjj1W3jPBmulo10x
h/u3WjhGwaOFNvWpO/0W7fZ61jekIMnZc8EirkMcsf2bWqg3jXvrU2ke9hQYfLbAeTCb8X7mxmKC
fzdD1T4a6AhD2WXg/bQc5ZFA9St0b92TLirXwLnBZTOEx11ApL4juS4VysbqWWGnf+KJSDQHdUPE
aOWy4tyHuqK2k/sgBc6kz/JqlEz2EUqNIc7BBJbk9TCNa44mo0HpvUeLHtyREq+SSBcVQBMfxqSa
Me7JTwVE1y3ieqSCimM0Uty1tlEtM7Js0S1B+L1R9BPK8t16BVntm5+buHVevUFOoF6PCY+0cHl7
Y/+DjglcIjZVsmFWW7LBUqSUGo7O7z4ZROunN5X8Vjn2akn32mSGeNVfe3wJP2FLG1hQku+Mg66I
9HbuGkO0VHvBERq2gJkSnT79JawZMNjwyuPS42HelVvuopeXaYuOOfuKa3nJ08eCxprDp6O4AGhT
LDyPh+9yPxDgoBL1lQ2qN3aAp8G4YdEXVxmJhiEopY3f4jXJfU0T8aCHHy283D8gZJLgp2n/cd+C
r78q6xRDHbWDX5rt60IRZleI23gbZFvJ5DWNezqs5deUbQbaJ6fs5rtS0rs2sVMJL+oNVE1iZ3iX
safuvpbtmd1/FjYQ1ncq6NLPN5Fvn/zzCrKqMTVZ8IYOild3ZSWNmCQbyUdAqYCyDot5lv/X5Yui
AyBsZ86+UHVtbYn9nzyIMMfdhPHKoIXxkQOm4+LvIPEjJ5IxQloq5+8QolfoxxqmQnL7F/7KvmCk
KF5v0xgdaI115ElNJytDG0+TXB8Cyq82newSDk0C9No07S4oYYOHzXy9YezBvGnOXlDiDs7gUUeZ
IFvedUuhFPvXEc36YZ3Hx4DBDCi6KMdFP1gExnTZrrhfkN0FRbv0B9hapmzZR4jwGq3YFPbx933w
6lVz6iYtszKTwiP5lN2jGvxx0LVmAKBmuhqbvyTqePNutpk+ITyEpAtLw93NIOjN3L7yF6ao+B64
sEvgDqCsRUhOojwO4TLRQ8s+ugJmIqgh3bRsBUCWlVsCsvuX6K1UNhtwnskwwO/MxX9XIsnCq40U
s/Qt6ARR4KrdO4YrZ/O5Q5eV9TvcdMahul/KrbxCks1lKZjuFeXUTtB1hXkPxqqWzcaPOfOn00r4
nfdMhV1Y3iyQKUPvsdJ5Kk1WqLDI2/zyX0Gz1RMI9E8L0VbXm1W8bJedDcjpkL28Ve9fIdHkralQ
yLB19yKxrHT3AzbEeuh1wCxarUWIiQ9xWdHVUO9wTRnkzvOHN8rIK3PVVwz1WuIaQOgQNqvfCHGJ
c5Txkh3vZSWDKbJX0BZqVJ9uQWztj1mkBVsFlmeID56OZPGxzlf4cMLmPCx0LPEhEDwFfQ+Vw/zH
Lre4E2rDuUs3rDS+jzNlItYRMOSiwo3YaE6wx+0FbP3NdZ/W93E29Ta5+S/H1+CoFLYI3IWQc5Yp
xWQLju/isBpFjhgAgKYe1bglWtEnGU8kfxf42UbVtNj+B3qhB9d2lJxnJLrEEm2nu3jEUAB5/rHy
6GqYIaMlAM1FZsGqTTHO2RJ8mHzITdaLvl8L66266FsEHXi8nPIfLnIoj5mOs2xjhvqz1uL4Pv++
gUVZcURi1I093sY/BgGIMbtteNsSrQv3jOl/m7wWUGQdNAByLxsVlgL7W5CVSXSiyJStmg1sthA+
g4uyFMH0n8JVJs2oMVo4LAns2RMm/FsCYrF7h+v2GR1PRcA5M2WgLsoPWaOGb5tSHhsEiyomz5yS
zfXMY4D55Rg/wJHnmpkd9AU/O35o7LZwUmu6ERbOZk6F3ZQYxhTtSHrsCWX3QlyY9cFuvTOe+mBS
QP4Ltwc9Y8KRRblox7qaag+ueUtawUBhAfW845YYiPFhlvrF5/MQVuX2hVPi9R/+t6H2y8A4/COh
3dn77SHGlaWY2nHmGT/U/vggTF7PShdfVnpahZCWoPTkfLic5RLlrqXghjYz27yUkWj1T7rvi8q+
hlCEIpo6w9v3IJtnTI9wpnhY6OBjOu5ADkJEHdTUk8fmlsUWndimlR4/JyuSHWpUUiw4x1PhPWWg
vFJqgmbwsijP4ENK8c4JfaqPaHERZk/WAVZfEPsvW0EDHz2G8cQlA+ahSg4e7m+1fPt36vthF3Gl
3eSjIgMhURbyBJ7hbLmPlCEoUzzukqvrv+RvqmssI1j1t5pNg/k1lY3ogn9CpxAbS0n/Z2LRTZ2/
VT2Rr1YlXGGNR+SGCLcqjUIOf57CaiIlzy04r/tA8mVMMXshZzDvzIOddF46/QPxO/zH2JxV7F8Z
+aegeWthcDur1ATqhDUX8CQes5VClG9bWrN9gdv9m+W03Z5heihrhex/UY28B8qgxAPtUInYB3ps
OP3gvYDPy0c2SXYrBSooldGeRw/e9xYo3YOshANf8u930zEW1TkNDn5CIryi1C+O+5qHK7eo27l1
YzZ7YcazcjShoxlMssLOtp7ppEwLtTnIejzGMEmyjXooe2uCg0YAqDv9WGHeGXU0HJWfRc4BOrmO
y4Ot1U4gT0yZp75tZ8/N5bPeW04V7FDG3A0cLOqY5kyfccm9uIGh2H2UmGvAi0+8S+4K98my+BSO
WjyTLb718ZTyhFcMxCuPXAdISThHlZ53rl45ifJjXHZi4KHSTL92sh2gJ7ymzlGSGYKHg7wA6Vz0
nGv8vXk8ETrQ60kL9W4TFUtkCCqzsld9PjyOg7OrqY+2L4dkd5oM2dKaWHcW73D0pUcQwRfU/HrK
tODPFSKEjCj+EAsMm6iukCmBUZxf0oTci7Ti96WPMlyvGi2tiAFlPq9rfHjlaQKq0myZDX9qWrJ2
QzYMvG30+WtVaPAUICcBOXlo9Kr5D8xB97CDRyPgGZEuO0rZPER5QWOierexEMuXtAnh4VXTcQ5S
o9DRbTuy4H1GcY8i9IK4llfc4dVislzkZcAdJjK230ybIDh6hqVILniaJrGcQBmeqaiDyqONkvKh
Hi2UHMRJv0y/g7CVzT76JC35WU/iU92MF1T7h+xiN1G1aTic9sZSVBrHwb28nnNyhfwOKsZGQawQ
i3oW/3BRgoparK6m3B4pdN/BNdr3AuRXdOe+TLFE1CIwI9uaDYHPhCiLhltFc0k0kFM7tpmPFsF9
lPHA8r7kzJtoAXg4Udpajm/GKd0Wni/OdhPi3Pqw/nSQubFiSc6YWCEmSN9unkOnJqArCK7KUy4l
S4zoOH0ZxYm3Uc6LucDitETNKLqBHwry5zh/O7C3Y28JvD0s8K/jYrxAQL+nz4qKHesNY9m2o+Nc
FakdH6Kq4SxGEIPtKIv3m+/PgkVtQfuX8igihdHOhN87b+ot6a4s4mblRH32B8jzhrsw2FNNjPg5
4GPvIWeeyzMAG5+Yr21Cs0ANCQCcVkzac8MsHoQgmzib6H4eM6cjnp0U24mMLKCSygleRLrZIVef
6uZM9scTeECCs4z6F8D0EovUZtLR2of/9ZhlknZlhsN33LbpHLYJtS3JkK3w8YQ6gxlRrO1dor6x
PcH5s8dtNVdQzRvNhYUTkMoITtEKVEMozfppXbPanJn3k/bjJ9Kj2bSs/KQo2P/BzzkXY2APJcfJ
wDhDcAPSUqXAAH4poTzAsIc9CNHphrI9xq1CuhM8NxMvATlcMAYSCt6R+H8ZMa4RA26vMUlSlsYn
IadrCPPvUA189vzd0pV7oUpthu4Igqa0tyOIy9mEiqaN71GDXUSSarlEQQnPQthqUSWETFQK6WfD
H+uk9UlrGawoZQC3/1G62YOspdCDLqrkTcLPftwhSsQ6dxxQ0La08GZi/a+4L7JmilkyrlXQwOLU
GI/zKwQJzQp89VmwRslAgXqouER56GTwhpbk54idnFmoDbLNFSj51HkeBbRRhEbI4Sfy0VOmjGwk
Bkz37rTB2FYuWLILcI+n8ngO7C5VH6CI1RkfGXl/tFRx2q1SV4H9GelhJCftSDfeVYcdCwWyjlMp
xQSGzvKKFTF7W7UPoJfBefLukcQk5JyS+WGemEK+c8B7lkGmbIQzsvTWlUTsthksqiN6yDXrJtZd
Rnv/K5ZUUsLrQn5Q4jDR2D0NEuvjTkK9hHpk7RMCEgfeVi5Wsg//uz5tUWdhSjAnWe/6UnWuRpD2
a0Ea8eGB+1pXZEKWeSSY78OX7F5DbzpX1XsYQUpDWRsPzZzSRVx5ZSMSjiGp2EWNarP1U4UPjUNc
kDZvgMFdgHejHajuWIWBWRqvnosHliPPon+1zSY1PyIT94AU3Xk/3uCsmIR8PwyBhCBgE2j51Bzv
b/gqhw953IGkbhopBJGvo5AU4hGFwbhUZ+yIijFOw1hjdl3AHxjEQxaK7KW6agh3JlkbfTyRALvl
9BlFPxkAhW1Z6CQtJqaIe3gpSkkjLKj6pK3tqmGRHCgFKD1Le4WmtNaVvKyDVu+eh64/ImQimGH/
EPWrzuOV1T/1FYbWjM91HFcSAXMWOk/vf8kdTCw3cMujquo7cnz7d3XxcSCbG5CZfzMdaYl/XXG6
tJWvTg0ixoVoyoUIN4xxhVMFdEPfo8XO+jj8TjVZeNK+n1tkPKOcTeezomobjZP2R2rKPGvA+Ldv
Iala17WKLYX0ve2vnnjOmxuc9Ti61gdyrC1yQwkjNHrOA1NpP+l0il3oS7ULsLItaMKzCzpuE/5W
i1vnw5njqCoBtpjhMhZdffq80KoANmWIp6qP3Qf3IVFo/Olx4O9F8HkWsm4dpIlxRa055lA28TTb
3SqnJ2D/cFMYoXLGIl6ahxKcn6GwEqgySs/r1WFjGDTsDX1RoiJT3TCQ50jNQAS4EMq1a6VVINLO
czj3Y7cH2O9siL6HKy+YQ9zpHUX8wwtUxacpjdeZeqNb+s3waX2HyLaIV7iauhgeAHyR4gYya7CA
3+iWIXQKxhRY1Tyip7XaAhxa5WI9baAPf6f48kGcf1lRzNF0i4Id3OtcwdjT1XULtP2qmyT7KFIO
Y3NIAf8d2vKF/kkOtcuORLROoYDrGTY+28FByUc1NKh2fyDOg2NJPt8zZgRNNOVCFiwK9oTTjoq5
RRHkPtGJi3IfBE61UBd7MubyEAaYI3/FQwEn87MRhxGV+ewuE/hTaiQeFD2ZtKYkqryOM0rKdirF
IFt5grclr/MGSyDSycNPAo1jT1frgmYiMzx7SiOFeWY6HqRnvsSpJiJgisxCdMC8awD89Z+gmy2n
7ZFxk5YoxsOqAOxmcYNJwcNl9whsflJ/xVnscibjaOGzByRsS0V7vVlntc2jgYSOz9/HHQBycqcI
rUJgTgfRW8/3mUsMpTf+pXWKP9FokBg74ScKPzAljZZaOVI8dxpiRIGpQQH1rxkZ58UymrHCE/lY
oM+nuyiux6KIX9kEkNVBPx/lJWEOu/ZQV5kBq0DTI6pOV2ac4UQ8LpAgvdxoQcH4JIvZtza05gHU
MTElb5LRFHpY9JKpgmHCZBh+KtMkX9rZKW9aLSgIvjsP6imr9Jnp2jFsN3eI2dTNnhS/jeHYHYhf
kk1qKCMJmmQCwYaLBNGgEN5YlxtCWvcAAo2Z2bNa7zAL19GW30JmR5OzY1eF2lJor3RmNcMszNdJ
0c/Q6A7FCuM282n4vG7tHGnmaXDjHpjNGs0Lq8JmTlop2qyrkjb47qRerUB43CElROwD3u99xclY
W6t8xp3GTG6bO9VLoBK34cZaYWDQlG7UMJX4KvROi2GkGmKMWwHuXSYYEu8bx+C1NiGr09uGxeUJ
UXNaZx2nTfXmVVJfSAPjyuc9vEXokFMDwReJVUYLMWF7HoalR0zx2Ecq3WUIPi8hVpZuIekE3IHd
ahYlWtMBgS/misctxJruZ3+m37J7CCI6+OMhY2ml8ujo/ptZUt1TN1BChnkKseZ1icfhzWDMWnnk
S9WseReaj+big4YVMxbXTjOPJzMbRUhSYlkN9/7drekvnmzGXSThOF56JYqJeSD98Of9WW/QsiEZ
S9kuF9UCWpdW8meV4jYXxgBeV6oHdSt2hCQfxEvwZSndOrPtud8gWOMeSTBkvQrvi9EwT9qvnjyY
OQ271xWurcvKFzvNgzL3M9FZ/fQYJtnvtJ1ThKFJyy48uG/Iaby0ZUv97oRnQ0pc82p2aE0ViNwP
b09hjp7kh7tNd/A0B5e/rNbaG7fm8W5PBiwTkL4pYoXEe3SNVDv7E5WOtd+FDUIVGV58NzHzPRFl
64AeYcEv4P9ckb+Jot5Q8WbPtFA6eLNJqz12CZs6+K+UrbSZ6/eSNBB8Iyn2R+/hIJ6lyFlUa8Qd
FZ8NVCOJ24bX6sTW6Q10NiAXFACpYEHy/pMH3nnWtFNXzFQdBSLHF4ITxDPnvTv4r7VXgLVyvhLw
02C5EIh7mqw/NFAUS6X9275py96BBPaSNn0KQHmoRfVtkfpobB8DWwYcKSVAyPlpTPZEyx74RA6j
mAI9D29lw793FfvIm3Ny/FBneL534igOjumQoXF4CxA2T8zQLObwZUGcLsH5x03hH9slRq+Hpyvw
WdtJ7Vqe1iE1kSN/eE10YFTmvXq5f2bg3CUugp0mykRoeoEr5DCdN91xGg4mDbDM1A02UosRxiSK
/yka/UmP/KiphIPZM9R3Z6dBumK3/eYXQIBnR/aogPA8TSzzx9W0LlKtUxnWD6bxOU5vsDh0MG0k
yE0i5ukUT/ABe4LGXdCY7ziLQNaTBreuqsVt454EzDlU1+HpDzLqRDI1vtdS+YdOmj979sNbJtTn
bYt/S4ZlGKabvK8p1v1yRgWHo1cLqhwaQkl8RXVNd5f30Kts0dg6iDCbctIe8sayFvbhmPfMB6+f
AaLg7UCGnbp0EOO684v3WCGPKmJZCNsYb8v/ZfZT7QAl5nLgKxFxcwIgtAVjvHQFeoUEN5IXPwDR
U9/5cr/HnBexZCP8wjdxm7C86cyLFWCjD2VMUK24zbUXAt1WOWF2i4OfpuR15WJPeyf1UbrguHaq
beZfmAYB3zGWlgzXUnHclM6m94X3qEPMgMH3kp9Ca4oDYFBDUl144LQR7kUS83W3jtTELTx6BNkO
EQqzGdaUxO0p8KNEbPEAOav5hsP+xIa/bE8P4k5RnyDWiiEtIfPAk1MPoqlbL6uUAYoXohxPFIPX
m7kT2E/heL/nxaA3onNCbOq8ASvv9m7onctfusDrHVImmoM3szc5GhiyzVFBca9BZCNivUgPzsDG
Ch6MZgJpq6RsytD46yxl2cYElshwtV5k2yyWUm7jpYBybqU2ZIkOQuKRL6Cz5BFoOEa9u40D5yIv
Al0qmqfjAX8ODUOvy5VWQXB+KduyN6csGmuxZCdRrU2KD4osJMdTVymMrlYb+8ePeresipmOKRQh
8G/dlmjhEEu8FYCmZ/Jn3lhXwgJw9YO1fa5RWAEOznJNyLxLBpsgDYMm8ewS4minRcWKJ1jiXJqs
/mZLmkwL/1fo0s3shYz1M7Fq5rXvo48p221dF1FNRfdcWL4uAXXZZZGeOLuOPGFe/HOPFX95DbyB
k7Seo00M2B1zkKYrbU0DOshzvD9QNWUcdjsr+b+Gg19cxQHuBHKqO+XAI5yeHqfIAiB2Y8C5NSa/
3IzgzhjbbGcqnL5jnUjBPqAHy+bZ/PSDZeiBez4Vt4SdPJ9gyUtwCdQ+MkoFA2J2XV0sBpBCxL0H
j0O8+greIG+7kn2l0ACRQeK56Lrm4nwtiq+qO/5spBtUBF5qlgaaMdyvAOXQnfoZ5MyiIJT5fkVi
MLa1NvPURJBqBb77C5pdIP8pQBXHyWiLIF5jODAhimS1gWjKIndXIHc2mglpeI7DhZc6EaNyBzVL
lEbTEJxQhKRhIylmO14m6W6Sb/KEIaYtu7xmDzWYvMjPDBbhxoupNDz/N/cgwfvEOiCD52BJwv3L
9A4gZBsdRnyCcENxvJCjDXTBEO1Var4qQqeNNaKvinaVir0JwsITkeuVJXBXUGRzH77WH/MTQulL
ZC2gcbVB2lEFS1+YGyvcOnSbK3M4gn2TjVERk+L51rcK/fRl2TRQcMjy1qKKJyFPKET2AZz9nGnn
/FqPXYLgYgcx0RuhZXRzcuUV8lpdFAYK/ALox1gzTBM2CdFUNezLUIXU7A+IRWyBzFS6ur5YPPpb
LSu/FWkHLgstAm43llOypOHq+octCwF/yjKfTbW0Ha6LUHEN+TNJoNYWMuawykke9nUhu6qvjxxw
L2zPlI1ABuG1jBYA0uxlgo1NWOSMNm/BXGFLiwf0hRJ/WLUFEAY1Omq7HtowSF6HK8VpO8FcA1w7
FxHenjvuLw8JVmOR3ZXA7qrPQyef4lHkundCpIHJqO6DR6YplFxnKGdTA5Zs/MaEmnLgWG6qQEK7
lTNlD83Ukt2qUBRn8QKco/e472UDt4xsF+y6imGAXoLdCXMw2bcC3CRmiu54YlB2iKvOgVZa25Cl
BhsEOviud415g5iNZIIL9ZVtXS06zBS0jkvmB8aQYNRpOzN8smOO03tPoNL75ZLKYzprnhmRP9yY
m3NWWcMzQMdO86t36tJx9b7Ra2nyDf6b0g0PDMvS3+V/4Z6XBP6JAYJ3mbHSx2pFdDl4RLYO9ah/
o/l/VlSU1fhKY0EpfAMf7mOrxvqJ+kn2Lsi5xzkiNcPn9QpGzqZwO6Db4Qhcxczq5e0tq6aZe8FE
KWbl82ZGMSVFj1I+0Hoygh8VoK58lTs+9+gATQ4UxB1QHMtgjgJbT9TWn0584R6+9ZV/THHljCk/
XyqlBblH4Wzbpo+XxBDBNwPiaBJPzvqcjTe9Kbi0AcvFDox3nwhqObdEaU0qjgJ6KuCdK5Wbuz4u
EuIcmdHmRe2NTJ9VlDr+Cg99IWY5tMdgo7ZWR0OsPMA1uuHDZQf5ZRQHF9wSnfZj0jegtOsaBmHK
cJ5k3fEpPaCsKNt5aB0VaD6ghSt4/FZzGIH9jUk5HSLqwSV7sTCyQmZ84ixQrLyXHh7dYPkU1u/e
c4VwLwtX0LPQSp0RfqEC0Tpbod37cKQ4de8HrF+SwxD+tDxqj27A08Jp4/O7IMfgCKsMwmMdFfVB
zwTSQ+zZf2G9rN4/D6GG+V/LuLhDnw5gavTk4dTo5JTToB0MJf28FroNiRKeLMaU4z5TQzgEj9yI
mIuaQ3aeW4v6KrdQyTFJJGOhMP5awbutuskxJuRFgP9CuSBqXOBA/i5gZYGWIbeNhFNQPkBWKLOO
XpQtn1uHUYY07jwlkwcH2872y8ct5gEowWF+SHIIUTkbeJ6wFNoqX3DmsBVBeuArDthtN13n8kBG
XUcFqvXNWGSXEoNnlnuYbkes8D7oKLHY/gmgKuyvO0c8B6KS8NQKOerHp1cWB9tLre5d8BmZHcHC
/AmMCg8FLS6JZTmqAy+ooRT3pRyFeH94/sdDp/XLUj4xhE7tfZYaBM+mQfs9i1cW+7St5V4j4uDT
G5dtxb+/cfryhm3eh0OzFmMc3xY69FDEPRzqew5PmDNP9sSJnjX3XDaC35Kk2gLEW6j256rNJjmJ
c5nuupjS6M6//L1FI9cH4pz6d1B+pIKfJ16XJhgftDtAEwOt85Oh3gRf/oYdpEE8xJuqMlUzbLEE
VsEQ2UWGQmAgkqorVcfASQ8GgpeYrht7AbrGcz4/SbcHpLcqv0/hsk4puh28gWDFqaiOacwdHo94
NeVlu9jg6Yb2KIZQfaAdzLXdNbueBaOtcjSH5J8RdMmcAbBzl0XGKbPK83LX2oCvOyCz0hNjpoA+
Yk/oy06oaEIMn63Rbpl5k3Fz73mz3HNylP/mGkwNvptX6uW+qZHbpdav3v+FSdP9XVz1w3+Reiwz
0hdv/skkyhAnD+AdmLMK2xR4iplMIRL0lN5TWhbOpKahv8j74yoaluAkP5ryFmH0Tn0xp2E5TiMy
eDP9f+aUHm7/fW6nUt6XB+AVhPvXr/b4NjVZSY6r7s81cjx6vsSxr2NxBxNt70Pj0lGM1ADLA9aF
GH/R3UFamV+x/8tOmPLSu4HZ4NC80JEnL6uzX4M0YZIWMfUn8CHO7T7dhx31SnpY5MWI+1mpeiP3
sU4QSl35qXFa/nFMNN4ry1zgeDuNsty8VDtRhDDtFlE4A3VMdFF5grbx+P0K8aSM8h/iCFx7sf3m
VAosT6uHGAnBgn4LkcNqVrqTQcklVUZMkg8fvolDG/EMbGNenirjS1w1n/Onzm28WV5kSukTvLez
m6xHYekzY0vMqeEdAkku9l/sdkzRaA3Zktfd7WYzVLLHuLTg0twYe9ueSQeIPAd35bShujhpZ4br
OFOzDIOdiOH1Ly1F4Z9NlxIaEILM8ODVx+/iOIj9KPjVIaJgcuU6UZtyAWJ5xwn00CqOxVMTua5e
PpN7NRwtEsZYYZlERwA7/RsMD2dXODU+1IZU+yhiLOI6fYgyN8cueI3v6EStsfJIyISMAvTrOPXy
dXwy3tFXXNaQSR4HqJcKdGVikfhVbeWmXHx7UicagdsfP+sYDz5kiS0Ob1eK1rDjGcXfw0eML559
jwjLezhIe0cFR4zAAKMth5iUvU/HHJa9gXM5zp44dhyeaHeORwE7hvtrM1UcIaVms/lvTAM0eaRL
6A5wFKf0MyWbTnadom5GbeboKHmZmdrXc7xkfqtoEVWsBZ8VccuJ6Fp/kITIQDGyyMzRWKJAANIh
VcINfMcd9QwAjdQalUZAU4hwICsCws6A/gPWg1WArmtTvMZyOHX2iKzNGdBtx7Bl1l3lvskFJFfw
9fJeWQzhsHWBz9eTjmVPbT7fa514i85+wrIVw6pcJ9Ed3tFCSdMmIx4Ue2rhGhON0MhYsy9hfEY3
hXiN/n7E/S/nUyadKGpHErObGh4Vt0uw0gsPamZnPcomlzZg7L/Ho8BXhW3LgGWovlmm/1XGxDF5
mZoITIDxT1yS1L8rzbyMStEuNytyVX7DvMLmnT3GBU+q4GVZIYNzrLv13Iu+Xe4yfL0MnWpyg+Mm
N9DYhxAWx3GOyHHVLzVEZzF5LybETlbXp3mZu09hhF2H7QWunTtfXShCZdgcCvZ9DOn/xstNDTJw
JeADUb6b6KqjYSHWWYwTbTNrCmLThcvAuW1lU3+8yA6gJV5G9a3JtTg5JrheSGcvtozfn7AblSLK
eDqHzjuO1cVXCqqJ8cPIBvdOY4oJ2ghb1dQKD2PuyLRh7SwI+WCL21xifkE7PpvZ4gIvSrhWqCWd
QcNWPI7ge1xXxyT+HPc+0VeBM6JtKDNVBNFn56mGxWJrMUwJPV1Pvq7iNcKf/va6goa25Kc1NJMr
O9dq46oXrbA/kPBmVrlW9hgSN8deHqy3975YwOt1i+wFvXTcsyHhMx+v5abk5Gt5Ohr0iI7zXrbk
7pbQVP7NfGh486g8dgokBRNr4qn8ciyHc9Qnfw/L5vq6vJmMGplwLZCrcbZb23x0rD2g1SjymB2R
tnmzdJRDB4zzM14Usu5B1FI8TmQnJUn7gJVyyDAD/yXfKIaqHQy8M1gPrHx5Jxq7+3lRbKhImOyp
FBJBgMVFcfkxSZVqObTB1zmWc8sPolRCXokEjqB0dDofmreW4UchPWttLPmaUvAcROVeZ7Jn0Xu/
ilbwkLRVKyV+dnWZhkzAdBqTcIHgsMrO2tdG0whSfm3IqfeEgerac4YP6DlKRVBJgysyiragI7QE
aYa4dq57fOr88qyE3YT/ip8qYwIGHUbTHcGWssLAm7qGIBpaCNSEgZOGAd4fPOv1pVIzvFkLGYxA
y30WgX/fBmLMe6t5RBR8m/WQs4M16pgczwW7yBFpMHp3HHEftJJEtgdxeN0/T06MCydKJ5n0uljd
DP7GI90EzbJcUXRwCEuwLP2yfPJ6HmQk7J//8rSc+UHNEmzLaCar4be/tUUY1r02+Vhk77TUc7i0
DPrgj6h4W63PO6jLtuKjWqJMlbePVbk7NKqtsTzfXbBlXz1L8F/1Pp3bCDkARAbRRXI6l6NGX8p6
D4n9ZMufgt1QJtpVcRQm0zckifI4SGl9GQY8+bt++HfnenmVsU5A5N+2dx03rEUCzLWPBOTgWFej
PieTCagOXbomxnUxf2ZWwVlgImc2Z9I3Mtb5O0ZAU4PCv/GUFOf//t+rAGbXunRBrKP3eSGzHg0G
t4hKbfMGW1V8AgGz4H5nYISU6jjEpWSzD2JwV+05vdbR9tNf1C1EY3kz8aCf8zl5xhqoKCWvjVHm
27MFgO/GahmjLMQmmc/6mbsSQnpyGgOAD1wHyVO9e9iTB69+FNhA9VatHW+VU0jIZJhXpZGVQV9F
2j1hYpXOYGR0zVCsNreA2QxZT+OW+johLBrkgDCF5rHBy7wFvFT0glzhxos5rX7vaHFmFtkuzIip
uJ8xeH3xXEm6OaB1qZ+gHECyDETY+VSn1o6JreQ3PfoJK03/K4Yo4AHehRW+Aw5HeLO8bLXHflK3
3ukSQADMD2ipY3rxDmQzxNSFqDYZblbBE4vbC8ZzxGYMep7wsIkUP+Xl9bUBZg8eU77cYDXdwoMG
6LMaainMmStE4NoHqKk6UXqKIH1EbwjWj5b694yYpR65o/+Astsxvcb4XXv8IV8YYCQWafGnTdML
KzlV4AGklGv1nwcuc2MOqYNh6ZQXRFkLmX6G/CAvnNgba9y/StC4GSFnMY60QtgffSY4PsIkcgAd
JlZwRGxpk6p2CMT+MvLC4YT9yT2qvOExR6rlkz93dIzDKEoYZDkSxXZ3ivJQkeO4tbGuBYV7rpzi
/z7LxVchWgQ7hvzfMun/pujzMHXyTZ+JtLga8TykFN2kRnzz8n75AYealj/8JE7/K85iQhwDUWnV
eNY1AfjmYzsC/5AzSC+ERPVvqaLkw1NOG3BGpE8FnHuu6zEHTBaDGCsuLnSWUjCOWXyeqh3UOFsP
B9lGTen3ZSgCEQvVvMURVCpgXQLz8iofsTvnByzLNZoCEOP4dEIeECsdwfCP76ieoDwwKXzrnOFZ
7dgigSlwFjnbhmf5vIbcTJeA3XPDfaMRHR7jbdYr66gh7KTwBkqvElJOOV4CMx/nTJ5+CMttZUge
L/GNfaQLmWQiK7EvEDNVohIWCul1FJ0UjYm+n2Q/4lxBv+1Vio0WarpeZW3eHDQvMUa1Gg7STNOz
4CWUI1MLDOjNmibbxhHVsMaqeCEKSoZYN5e/Qu9EFrSRPeuqX600cqMzclLZE22aoZ8R1FXf7qBt
8jUL9aNDHCPQajYFxV0WKRchcqwlDfphF0PuDElQrKiH7TmyQzCovBbMS2EsvD3lFuCBHQjjUWAz
Y+qW/yobOdDOkU/dlxi9Ra8B+rMHttMTIgJKYNBdB5Ft+r4vEd1n2p63+30VrbJwGC3Zh6lEtWGB
IQGjSc08BaO7ndkylMIRilEfBLCnKTNqG7wFCSvCtqfcF4eolx1Zy6nGmiR6qpVcu+sg+aH2bc2J
/gVJuczUU3NrRpqZgtthyGpWAWXLRh7/RLGtYbt5VypdGxgUvqhukvDuCXp9I3LMeHT/s+eNlNo5
D3RGbhSQ7fWvKtZ7njVijeBJi9OScsgrHst/j85I4+kvE5ROF9jgMQZO1/G+E+6B3rwkSTKKKroz
+6LoJ4XpJtnITVjkxw+mghcyj1Y6r5bjKQWzO7eOCsxkOvWfhThC1egmNE5cP/ec4vQPvBF8CqaE
MvRLsVgT8jzs/06jUTs1pOErFFLE0co/HoZfCQaaKFzIOwAAFdTF9/cv504WVaENfbNlRkCXDc6k
7awX0jh5kN5VvOsstIz1aFSMKKMuLdOOGciZjvWS0RoC21fLR4xe+k8gaDDDkxCjOljR5UzeMW2J
+lEFO0JLUXbysw27IzRnXf5uaK3Trk1R8YxEmwHxHhruNw8H2cdSTsxoI5yeNwNqJBQT6k4o+QVc
O4uQhe7OBI3q3zd0CxA8jVu17nw5CfQ3+vZ3bc8Q7PfTscTv+otutpERK064ThBIpaZlf8C6iQJ2
EjDVY7lii6zejvGfgZ2mPivI2uFPEUy/65jb5+EH6RGmhIh2WQnImMJng+Hy4/Wb3wVjQpMtjnUt
r59rqgSrCqaR41+YHKDX0Fje6HcZGmhW3HhjARlcQCJnc3yDIeE2rkPz+gIkGgle6WvlOUeLqtJU
iOpKASzfir5frYSgquOaTElmmY1TBqLpPYbl9DlZlI6rRYMvGWQryGWO3sFHa9okm86bRwB5LAC8
y/fpjjBxxaqs0s3NLOEu+dzzIVlfX7/53wS5LlV7XWDBgJVXkZ+S+4azVdMM/33WJJT/MhicL2Db
QuoelBsBgTuRnQp6eieYo11BE/fo95SoFqfDugggTHZ4rXWK2u8I0N/aP8ueBayMElUMYBaxIRTY
irmvtpUH/Hf25zEdxt2nqCebsPahFYzG8ye4xfAFqtDRmKBLW4BlVgitSR5XGJpgOnL5d1py/OSU
y8bXdDMh/6W5LRKGKv8gHpVRD9spvW1ym4SoR4s6g1Jq9B6vju3Ft41tlcwenrHX+a/I7G6B2a4N
XxQ51+SUNVSRutZrKCF750Q7UNWXxKlPWDvlmpppOFrQJkLzfioWkzRR/te91SjvekAh6Rrf7Hxo
5hbMOeWkgsM/oTLy/So5FixiJrvR/bbA0f0Yih3lixhbu+zGPw6IyeqYW7f1gCwLP7ix2y1/vyR2
p2IoTnTeqLGwdcQICIQO8F3j1yFNIt4BIS6dGr6F7FhphwnFeZEC/A8ovqDfuGSlViDG8seeiXrX
+13GNfwxaxRh06RKTjzSNy8FsWUoVK4oPEM2fxnc6jibAkQnmt0YanIloCkyWb/ouoD/UkdfI/zk
LyBhjtXJILQ1xQWeTTJMXe6v0sySuEbPvIxVfCg7ExIuJ5E5CmkpoI902I9cGjJ65F/P2hYqqwDw
lLDeRZnKND/fh7hGXMEiLFedkwK3ugtuQf3i5qNs/mI7c/zSJylW2SeWuEajFAd4TASkfADXecs0
jamM9hH1GBnWseZ9JucNgW7QRNEd4nNsmPX99lnDO2oxO9Gsa/PVoK2AyI1BNYuaLLOo4LILBFde
Ln9aa8MqBkdcCSfjyklNcd2tXBEcu8HJ4oCZ3zCQpGpoP2Qd6OZV18hIkJoCPruJsJXgifxayzj9
p8725Q7XzllScOFYbBSr8/sP87al78kMRDsKN+aDHKUrc8BjxSKh6zqOczPr8EcmEYyOLNUY3KjJ
SZdGBmESNf3Bg1PhRgWkcs9n3d6qXsviOs5wrjR/p13/Y53qMaxmOdLdMPaSsFaif41Z4mQKMVCJ
8dypKluVlkG9luTwEOjYZa/DhsbiHfm65gWxUn2ODV+dhOOoJkHhYP1Ms7rsJZwqFQW83tcrN7i6
SYE+Y185txCNxvHZJ4m7DX02310MeJj6Wfpi6R8HNmNDSW8dno5yAnLKxa8+hzY5N3+8p+1lUSpN
0BBBzoEFCz5HdjBL8YhngrotIkLl62+W9xnlrv2WQE0iNGpOF4OnyWOX6WdrpISKDmoAIVM54wX3
0ENaD8CR0a2uLWzZkg5ShoemnUhrkPcUeHXxNYcaJmKYO3vvmthgdGBi/2g2jM0axFrryFSLKwX1
1bBHTBWsFD9shmulHtEaD+MRk/V5EYlVZ3MtFwQmK3b9C4cBA4J0rgpdH1bSlN/RHhbCn+XONWMI
r9lKx0s7rnsaiKtpcrgY16KsikmLg+X1ZxDSfN7CtcYc9wNG1wrrZC2Ev8O8TLKlPtObscb5oGud
fSKIj4TYZRuzOxVpFZvCDZFQAykHc4pvAv0zhH8prNbqBFOF1p86F9JWSmJJbTFFJWkC/8BhxZXE
fKxNLQsbJNdRwzeiDVXIifKoaXJuD/3kXRR84tkssyGslujA1WSjuc9Fk83WsoCwHp4fEaf/Faak
ZStKwmB2+z8L8ZEWzAGbFlKcKsgDQOP35LiMdnKljMb3u1pePrKxm9FxTDMUOtHBFpYOWQPIWQtC
x/UL6cZn5m5EfZDmPEdJgznrSv4xx5NIxzMKrmednYxkSW2oPWD9zBw6d4SU5Bhvbx/Cw8rHFy2c
L/oLLgBagqR//5GF+x7Y0/ll3lVWKLp+a+U1Wrz1K6sbNmWavBhpgaJiiKxlJDmhiZbz6I+ajbSt
SYcdk2AVNSLibRAWyGRgn7nwKMwpono/PjPQoI26e8VBtfcl8opzymkKn6syotqWTVKUakMY8w8E
Bm29qKd16MkzFcYPxjhifBFtnYtJEex5u5N6jd40jilnWxZHLPUmCEPGFEHRRdKPaLAS7bnb0SKi
Ne2hml97NXCYqEL7zA7eIrZyeV4s7eefFuEPKbDjGumHtIotBcP/4h6X12Ah0uEa8ED7/Rrph/pI
0P7DA/No8EMZ2odkuGRAvLkyQpj1iodKQmR6aWiPuUqY8Ue49L9eKSsK18u/S/fWCqnsw+ez9889
5xnuSe2Rn+CUeqgP22+c0FVA/P24mCbvAEvZagT9CmYMWW0YUhuOMSNCGlYnd+yWH+uOPuGe/NIl
7y/MxVbImvA4uI9Y/3/OQlHnr6tDa3KipANqqRae7XYibypKCJb9vQGSZboPSCzqr9+5Nkdsji9m
VeDIi/IMVCocLZVPIVsvUBwG/6zRQbJikuw+tSgDbBqFqrpsY2aj3oacwwEM2Wozo+niH1WtO9el
wmzmyGLhQ7yMz3p5dz1vOTD/2Cj7IQe3AEeaMKBT4/FBp/ccIxdyDd61EeO9XJKAj6ORMMzDB0FI
oPxtelF+yG6P0topDR8Wcm6DXcFy64ymMrVDn5D31hXsdPc8X1R3BMeSDGVVSeTbsL0wY3bGPmH8
zS3hc1cNdNbr5DjXhgmBv0d0yU5VB4DpWeyBIkOZwmwT8Vqz+V4iNt4O7d5AT91OQShYISmOT9QB
3HEGk7DFw2XabFl59Wbrh/Dd7xbg1c+5k7k2YvRpGfjvAdWsgpEmPDfASELHffBfC9PrNTpg2XIT
GiQ/O48+mEAMFcF0+BYeuxMaBo48TDOQIEvXUKMaBx++7vDmbRZRzow8YLPG4ba68o9d/MqvsmiT
v/8BO61GEPiOIss4XdAZDL0Nxl00BtW3PCVTUIen4RmvU1q656yMyWTB5KzgOfhT6NbHzMU0wIzj
40SvUar6H/x1MwozQtcbfwTRasbWS/xilWnFddg7IUYFEhmdGtPV/es1/PNVlashyLpMkaP5ZLw2
eDmhuuAueralRyHhAcr7JmI9x6tEjRX80Yz18N1++UvgjWLbL65vCJEsHP7T1BtOIzPgvxz1QP5O
rLzvSFD/bmia67CRcW6cNQqqZJPYl6tqdl80WyEtOVMT8Jx/rB0mmZB7/4cvzzTtB+6N1EhohH6x
HJejnxVnIqeqMtSsTxN4jJZHkjvYwSDlILe2Jt+bur2voAeNJXruTKH5tTeNHucL/jZbmGWct8cL
3w0DcbarhDrycrquXghOFBIyNNVRrmUqZht8j6UFiaCm/CELypba/ifFgdjidjm4hmANlUfoJCRC
o43I9DuOnbmFPwk+YzflMvrc6DDDCu6jCZ6884RnF31hOlGDYiPUComSjneMdXIoC3+0QFEhoUEH
iUsFjPiWI4B8u269ZjwoHxcqsPfsLVxx0PptmyMms1MkVSr4GYAGz4a62ABf8qMH4nGQlkGSnlmm
FUs437n6Nar0uYv9Ooe89sCQDOlDoGxMuSPXKJaXFw7ahI23M825DYkXPEfchwgxrjpL5+MfQCca
E2mTaZGS97tfcdGsRE6zCU2iwIXDVRaGgLldq5uDCFc7PkwQnZcQs5OZwT/FA2EPrn8AqQ9+wffo
zOGIDL8BXM/3ed7l4ZlqUuoxrChEEVRvUOj2S22qsgGRZA9iRBRg8wVnXGRrNgtavRYKKusJtHgk
RN3L76JKBNlklQAN7pWwLjP4D65rFsmyEZEGHxepmQUZoKQpWTHqkOfI6bXn5YilTdK6nusAhHZU
6B33/pm+FS4xUW7ycPnpyYM7IWvkEEN/RBiYz/5eVISAFjsg8qpe+MjbmhfmUY6Y4eFGRunOP9eB
clHAvMQAxPRXiZsHfYSErAUhKOpaecNDWpI0Aj87xX9aH9rcWOB0p6ORlYzobbsqXiqcK37JAK2q
WIi9AqLJMk8N3tS547jz/eSEQzK5YuBxh+k0krtasTVsL+xC9w62ln2+kw7SRBaqU5hOhReJWHKt
FT73nfRW40qWnk7P/xi3y/10On3F9zZVwXth/v9yMcS/ctvgwbxp8oZJavjoxhy0Ah+qtfDj2qvX
CbguGzVnO6DYM+90MTbFsrswAb6tg5pLud/I44Vp1PmL0kbsK1Y3oZfaOuCi580t7q1v5F/3ztr0
mvwuCFph2DYX7iQOMW5eN8VIIwIjUYExwLz7QUfq1ryXiYQzTGCYkBp0FtYmIkEIhIqPnclrhszh
QiBM2DFAavU936KKZ4uvJLWKUT7xq0krf98D+n4P95oPOjDw4AfzgBYnHjXLkczDnU2We0bgytv/
vWA4f/h+Ue7o32WdhDm4WCWrp3flRS7Z4SAf9HTjC+hPlEiIWiBF/MFN0l2gvF7npoQ3da9GVlKh
HgIjVg9GvSydvCVmGr93yEj8id800AOmvJdTZEAoNcScMNM2tEbSfBK+X7RuUOEVAabk+c7E7mZ7
cIY5yferquSL8Qql7EuxOolKmv/mfEDbPvPoj21kn7Pn7weYP7VcTKQ9zKlSpVlcYZ0Kgaf0PwyL
PNFWHKBV5UqECSVIbi/QSqypuLAEKvjsoZQq5ylyjW8VdNhNd/BrDt4M8LxiaDoAT7v0M6Wb2Gmc
R2CWlVBHS5EBnjpYuE4Rb6gMi+AZxdhataiZ6hnzzeMQsCiCGMzWWhwi7qZ583HSbaTEsZ0KZHsX
fWkrU//JpQtsUL8b6apakIE5M70/nQmXr9vfkbsHTgDRdkkIVcoaeqWBzJxQKTFiwUEbjlo+cRUB
GoC25fKEt7GtzdV2/tniWCdFVWbw3RHWcoUDvKFZShBMBZpsASJQHkoyBoLLtbbcp5+zlQtQaKFa
p4tm4Jjuzq8L9ySEFiFWDzKkmU93OvC9lOssuQ6Nw8D66gdRa1og0/anVJjUlFVaIUM+Kr+TYwCz
2wEC0J3dPE35/Wmajg71VpCA9fpagmO0CpMbjBuZbjRv6hNXrxZP52bsJR9TiOSq6ZG8BWvQ2i/8
2OBcsODE7512JNo4OkwtMbIbe5y3r3DcYIDKjgaaomCTDVPbcq7+Cab2fjqvRQbbj0rFPIRro7V4
u4fBxEActjCzKoLdCWcLSfJBDnXNUWvl/oQqajVNR6ozb+0/X04q+n4NwT33A7zt+ic4pCJTQlm8
cylSC13TF//SV95qbBHNpUyIK/5IDOSzN1w9Jg9P23QK3dy9olz26SfFhz14+DjqDMuiltdN9Bh7
x/GjFwvWPHIdazIG5zWSgEEapTVtb6XWtZaAFuTU744ANxlKjsxwtWU7pk/eXY25NOlQkfK9r8Ax
2qJzvcRa9SvHHWssWf3Z2qWRiSV3rHrULqDaC9i5nx8ZfpH9tSxlPpRacC3kIXo9NY0dXzS0qr/Y
7wkJtSx2pEtXklJ0jYa0NXsX5bG1/JobRns9Hnl9oa0t2qap8qVY+Rm0u8rKMNtgrDoacNo9b5Dj
MECd0figp9Rw81wzcnuitHHycoPhMdkQ4OG/IT424IFQFwzXNQz+U13C3hIp7R5xzT8Oqv3oxd88
F4zOQoUnZ/NI6VNuV1/P0hTvnDyVS6eyd3yaGPxkTEvLN16OHRP36l4CUHQL7R9O8lm5EsIbYimy
1GkXjB08QVfq0u8F1FZfoZNZbpM5mAjiWzNlPE0J+quup5ya8zeyvDA1KSs5F3XJXTIlv8h3OC04
dl2uqgSYSb9gdcj+LfFb8ms73VGIdkQHuj6dg4ZkbWYs3aC9zNLacXLe/fKydiVqahE2z2aT//yI
JyV2MUtL4EF9fvv7ScvIcIb+8hCKSuoBX+MkdyhU7Enb0u2nV0odB/iV4g2/3BMJ6TmpDAe2fZAu
WmxTgds+r4/S/04g6ESLH1htJDve42fKYNcXMbAMq83zee1CqDDzGSgJmPy/07ZwWcDSToqapuyF
xqj6sZfMHhMDw2qQa5HkbE3ULfIHvdDu0KhcnsK1vIvJwdCNuE/26EhFM3p8LSo/gxXMjN8v639A
bWKyoxUPc1FtCIt80hkNihw2LwB7t883sDGzlX2xdjm2Hd8uzv6Hgb0RJfy6MxhU7ZFUiErLIq3M
XSNAEqbp4qFPJUie0eekctMJt3kD7Wl0rDI2h4VQX50EqKRRIrSzgt0kqZfUqDAykQbly1LBIkOA
2nbN729nszMoWuIH6exNZYGdAG5G9QRUbe0YbkuH1xGMI2za5Tpz0IfJIXs+p23cw/ErgqZbNhX9
tXD/KuV+bD4HExX9eHSIjeLst3vvFi9JBnjwYjBY57s6t/PYWxV7eNmdITmqYHBay7EJAJBObCHB
LUeFwW99Qsmy+PBMIOk4Uh3BUGYRMsiDjoPIdgvc4naL/KrK7yDwwcuQbZPNVPznGE+rIc8OxT3e
ydlm5xi881Ggw+2E3MYyjEusiiK7NoX/8w69jt6TXY2J98TaCiMNekolxTw7mY3UaZZJLD9kIDqH
pLsj94U+8CTSdbrGwqnJDjn+MrL+5XCcsdgVcIJjxGSsdZpuRPHGL5O80I+jtnfERElfCJbYRvip
Qrsgpg0blMGsgQB2f8yZAaJEMacdmmaly7sxxlxW/IvPIxWnbCF9mWWaCAbf85X8m5FYsSKEIlHA
FwBM29aTGnbzLH5g0NoBkwyEkJODaccG2bUE5gpYbhEZC33AqKnGHq6wgfcr1RS2C9Q6fAfreASK
yEHCCFSLSkaLiByyt/0xf3Fh59y9hBqwQ3E8spAYC1cBisQlTp+G9O3A/KkAGrVYmIMl+boLUm36
m+ECLVrKUk+aJX98ArfQ7g/VuzByLXNAMEX0laay7qLNCqv61Wnag9Rm0Hl6HLUEHhUSIG+P9qZ2
PHCBl65t+fIMJG4U+jwkZxGeUDLKrBv6E4aaYpTRnOAQtOaG7hw+KX37Vy10HZhdOtRHYJeFiw9f
y1vuMTiW6ZF8Rh0JQqBYFMuc0a9LjPHqtE9PCyjY3DGixQYESXZI5Ny9CsrTt9s/9nmALu7Yqdb3
q8bkgw+ow2qC3jYBBchcNPMVCcTAdEtvrgdypnPTPEJdvXkQ9qiqVoNMhEPS8kY64WEMNTS6+hQ8
tl/A+hgB+gujeyJKn9w+wGQqHthL7zRf0EBtB6Lk3xuzPXvlwxR0FpayK9vVT4LqmywbMpvmUrNb
QGA3Qv6J6WacVbSZ/5E3iBwcfWvIHf8Fa67G6nGg5K3gZbnZuIEbZqe1mvPO2f6h9EHdWEZnN7qC
3a3ylOFttPqXQPZBK0plFAy6ZpQtKh+XMwhcQPvraBlm0gdXUxBHSqFm/aM0lwUQGuYTc8oboxv0
9jCP39claiMY6Rjh7loH2ET2HIBeHbWpt2++87TZK6TuG6CWLsNJcImYA7kum7AVvXw7VlAFIBAf
Y4+M0hQWVcXEc6tG0aKpWioTnnJyLCJ4HsVXr7DWQF+/whhb3A5vGuzcnOJkjBxKEynWmmGbWVhp
h2E927y2fdvSdbQCOF+CBbyGskgjb5huaoxgJJQ2K2JZA91GSocytPTIX5FZ2+h+ZS4kOUe/c7QC
MfyZH4H8bBg8oui7GlDUcbqFfISqYm0yBe7qFbtD0tPCQg1gR/E8YD3HHpB5zegtZXJRTm5BgIgI
z1lQzrNJydV7KRxKRW0PbvtuockthjMpjOFKxaieXnneDwyICvLOJx6Lz6/JG03ajX7mfxveMdfR
KEmflBMqKitNGN0CfFOP1qjd2P5uIbNn48vQV2G6EXhT5z/1GeogAeuZ2C0YKfPD8VcfaiESZZX1
yUohK5rZb+gpSH/nyL18g9vaAutn04Rb49MXTxIq80bmqpQAakyki51y0uZpKMPzbiubgAJAzGEN
GvNW6CdNpqL3MFyaM8pOxc/5ZqQX559yX7zU+xzPs37y/T1wuxib2y7wQ89NaBkb4bG8NT5K4f0+
t8YPMxJQTAypz31Ty+HsQ97OaxaZKdi78x2OgzHGEHHO26+ZlzlRusbbsacoY/coTkdYXbCd24pv
mQ==
`protect end_protected

