

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cIiYfk3Xy6N5OP4pq3GmqGiiVNUZ6H5+UojetFJBvbKolIu21jc4BnJQVK6clVlXeOqxCwUuMeWy
2HOHrYFv+g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lIziGPDmnLk8lYYpZIaDaMbL8fBzq4Pr1Jhh0ulXet+pjCJLyV5jakxS1oSptZ+tHYCT5i9DwoXk
484l0YBwGxIV/F50kQ4mY5SmovR5v/32XWyGw8Sob1+z/rA/iYbfy53jpQjBFTMhONxMl2jPMKOr
8b4lWHN3CKPgzR7gpH0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
htRzDc7r6AHMWLJSZlCSE/9tAboPhTxPArTqmJzMnfBntgIxMOX2YAPT8iZ7gZlglNlT/Bmc3ZIa
nj4bYkmP/Ed/Ze8J5Af7OuS/hLPfbdPEIMVOJrAzPKtgRUGYzZFakpIpDVbTLnXVCXGbnWwhbHOl
N+MoLyC3ep/1xGkMFlPyLgKVegokAfOd/5ePZ6yal5L+KR1ET32v4t5eGaONowzpG0O9uY8LtLQU
iVJDGAf4BzpePmtzOyeo5v68FfUFTjm1d6csF3e9pbQ9fEwJazksjJfyX2XYuUZH1eu5bhyJMU/O
c9/o5sfORhKXoxNo0FDKepouEYzneEXI8uuD0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FHtFxX6m7YezwdeWAQ6jmWMHTTCQ3ATyb5990cCrfHVNkzUwGdq1shf9GRL+uR3C20sVQ7v4/+tb
aJQn0JjlSYvQTO2Q6FVyjXNHAr7wpM4t4p6I4KuMXkNXuNp6PVpERQgKViWQe974sEr/n8wacl6w
0ZeeyAlvAxPvOHeW8Sc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WrHRD4nLu8DRRwrUtiyMH2ZN6Vs3L2kgyFgp5P9DMlNKTdIDDQa1yTQPpciIt64OlniyoYCatBqg
Wt8N5KlawExwntwLmfujXap7EAFuw40uyJX+yki/gczIgekz/25Q1+NPVfIAzqSReCro4UUW45VQ
4oIxLBIF53PvEJm3CGD200yoSxIl9Szkkq1FCyNtIufy0im7xj9CnEg/iFEwxzn8s8Ge79lV+lhg
fO4H7eA/Qsx28fzoVv2RYnMwC/Ln7iTt2527VU0KjrPDX1WGbNCJ5ny6IM/daMbuTMvJb5fz48+S
KUNyOcNxuhu15WGxxGlN6mcj5zB0r8XxgsnOfQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25744)
`protect data_block
UaECO+Os7jgiGIhhGzxg8K28cPduFkNBrtCyQfTUjM6i53+vLn/MdGvhi8Q+weHmR7Z+wTI3pKLF
mmJD/Wx0JHjWUMUs2BoIvlZ5mCbod4mGiIadb+O+UZWmgSqDlocDisX7SBu+AVFa7spGT+gVxts6
tdLMfGrMl4fIjCyEaynfUmGI1tIF1s/UEmXzik/bQmTDu06qOlknH08w+2rNrnbBTJVjTFcKusuX
N5SWIePXulXA5Q9YHSmilvLukDd8O1S3r8OsmMEE6ycW2nlrlFbEhmmzaYZuMOvhCJ666HTSDGDl
z5emkyKobtiLgrkVsRgfMUsJL90P42i5gZEINM4iuwODvyO8Dlbvqm5zREgxDy63AZ6DEZX9BM67
wRY+AUvdLFSx0Vi5N1I4tQAC1AlHvtN1dsrekebhWfs8ciZKJHREshfV1pA7+ib211CaB/urnsra
orIHCOweSh+3EGq9MbPrVc4yLZzxW+LINE9JTZzHD2L4gOVgwLtsknmx/nT3RSgBsXxZsnuB06h1
uk6UBrMyrc7m1UTIZPToqMKzGSgf+LLRlmhNgQF9eFsm86JI6DII+6ZK0M0BuDxcsuUI3mfcerhK
rGD93Y/CtPSWIwobumoQIlFNfk+jR0snxg4qotRoVOAU4r8Go775aP6Npaf+xMA17U3tH07wn+XG
FM2nML8MVnXe+2bFJOsdDAZGkLCZR1Q8jSjHXWGACqq61Dr1i24k7Z+0fVOuhLnl+LjbPS0nlrCo
bvXvB8S+v4mq5zHakEumT699evMlrPyTCvhwuQlqBuqcgZPDQLMyK7co4KLKO6DO5+rItHRxY+0B
hXFDuspkpSSp3zqvd7IXTQgC+TDStewcwciHIVcj8ugu+nFthYVcvpM+i8Zom0QdIqENDDSTlk3P
eaCNf2cjVJNoblcj2Qgd9Dmh291t/sIwndN/11sFOX6d0+N5wdnrA/At4NEAijQR5mCjXHJIUDSf
zBZUCpt6WXmwdVzMxdds84oJZd37A75kQWgLaOntLQhMCqPRK2Dd6PTt+VDLVonYX1AAYBTshnjH
7xplXPd28Zwku7ai8R+QyLPfINhAs9hgLmeF5bOcWhwLEHpeWiyX0PWOoctz1KJN+AGE8uJEhL7V
A0Tr3d0KGDppZEDTfSSU2lrg5uZXQ7GuAVYRhoYp/O2CN57aPo8COnZ26tpQEj09H8nE3z4yH2hx
z2T+HXClUVcY/YaGU/1KxBWBkRwDyOT0yuhh5nuk4vFCm6SVOCPn1Rl/wKalA+0e+qwVs2ZtaPYD
SKynNBSlH8IUDh7p1ecGuHEWuTz1/2Z+8bQgX6rxP03G3BC4iHB2kYHiLvCM4ZKgU256I7WZ31Sk
As1NWO4Xh/QtbzaLlcs3GYZdhdxKp7nGBQhNy9zOGtz6IWEOGSGXiBlMd7neiZ7V7QQ3mu94SpYr
kiHdFgkjnwGtQVv9FhEnCBYPr4NW08yEzwNLAoCDc7opQz7mVsXw4tijw34EbtorwxAWenIQUEPR
YwdsUU9KTmgwlBY7M8kJnpdbrcSPk2yU4AvdwAzjP8EIGItxhnfvyxdwgCAxz7bnYjF82/GQ5lK5
5KGhHvHDDOkwht9AmUnoCavFgLye4/BpMAPpnnDeITFziIXUeBIVCWewHmCwJkUz9sbKkMnNGShy
zKv61y1scIewD8DwQnm38Znx2thHC291xWPcS7yBWM/cusBYrA6/AOdhHbnK9XbEeL//gr9ht+FY
TDNZR+It1RNRrJTdpXQdlu4vYvwNTDkkFXEbTmBtbkM5+ULATTB5n2iMmXPCVhy86L0+T3W+5n4e
dsUtBZIVUNly2OhvQhVvYFsw+d2d+gqjsIlc7oGv4U9oDrouwn7Cp6ISTU6Wu7RY9yO9HPz7E+1Y
+wp5HKaEAj2RZGH8iXOie24m6NBxkk3VUvUAFQuXXgKXpk5vf34w/Z5K1aCIn8hN3cCiFskg0cNm
UrCRlgKYweoPdH2M52ZOMqwaW+HlJ4pmRsJnRqAtYr/ZPeUl5kkxR/a7jiHP0m9HWq5xYAPUJmrD
mpDsOENVCxCXgVxGMn0EmrQXJaNaXq8CglULZHbN+C2tWkKThEiuuwxdob/aVoMqgW7fsPy6/Al7
7fM0F/UmqSWK9RcMEnVjqGU5ULnIZVst12Zt378Q6K+AHT64wVu+R5Z6i6fhbHZSQrkzwKItGUx4
jnj//i84i5SEGbh8lJCo4vM2L/1PEwStFyQlRP72BVVQicWHMunbrXZzHHmJoA1XEkh4ffZDfH4c
F0DqghsfwvG9MXg4C2NaEYacHyjDxEjed/+ESbo4F3z5ctQOOTS4GMCMtQWGnEuPademy0fvG3n2
gHWqEardNMGTz7Ubz2v4z7MU6PDU1oJ16RBwxftUXmwrUlJLqZWoaVeLyWr23uvH+KCNVGoupRTW
GBPtz400OmUhJCiRObWfoTT5WPz2kAnZloLd8ktEN+aV7fcPkWXN2sLkT3J4X0VqS3iyurlPHN+h
cinsDTkn9xXOnpX0KzL5wTqDNngpLV03lnPuEQb2HJXvIoUNG0o+wHtUC7K/flLntxOHt3xjTuH4
danWsUkatM0oC1m/r95wUKvEQKacr3OxaOQ4EoXKXcjjyzcik/EUnluH1nPQEmzQlQPB29Il7anA
957GVOlk0K4ueaC6sn8lk5n+pLjruyjtB890AXnnOYpJVz/gjGcXeER9/YLy7DE0j31n2wRH5KOE
UdKl2p9ZCDWknYYqbC0/fxAkeG1xZQny12Y7M5Upuho1JWCSBw11FnJxPuyNlXnn23rR2Kcrvq+Q
4JmDyAJm2EJnBEwflT3E5ZMMlLle39Em/1op/duEialWcGdRi3jNTLJTuOeppOVcjrcFOEhSOqPR
a2EG0dsYKfw4DujcF2ajzC3ss1vRTkOYB5+6BEf59KvuBF5yKqeBkEIc56v3MkahYpas4ceN4Z8a
62urUmc/jHlIucrVnvbCGMvU6a0E6x28RzUjUfh2xvkCNX0OlvhKz8NTV3Vl+i7WU7Q1DXtSvieF
R9ONYdgOjRMYhnr1/woluiroMqqMsMUKh4juvbe4DylzuyktvHFKX6/meBrpEBf+My0ZWJbn5AE/
zE3T7RPYM4iX7V1R6HVXws/rPT57uODY5UjuPi9XX8Vy1/D6j5mL6aV+obdDDNC3WdHshQgEhlA7
wSjDoT/BURAmIyG44u/8I30rmSUWgXiNzD3vVHZm3g29rk5YKKR4mAvniq3ck0yeRgPsW0R/6kvZ
0fujpf5UM/Z0W8zkg+5YVABB3qYtZAv35gAzwqiSiI7i3PBoUQ0kb4YhhZDrME0uqEDp0OxpvMdl
N/7tIPH3uyzpKP+yXyN4e4F2i87npIlafVHNrNI281dME5kQd8oSiZJi9bl+Er5RqhTLc32kieme
wcZKtF6UawoK32tSM7B2E2h33uC3Dh9q2FtQ34O9gaefqXYbiBTA7BsA5FGBNnKQ13aMBPVHqjbM
E8MQ6LRKyPoi3j9imcUHQTqqsB4ex+/UiSiVscbyRJwJbkEjVFliVIV0Iw7tWRv7ZM8FOhavH/no
ddo35NeyhEyoRMPLCd72UyRMMKcrN8x25TjtMG8xVM18jZ6QAWbVE6kyl2Pcg230W/2rIOzF/2Zr
tEayaWSKMOL+IPS/G+ANolRjCz09MHlkmVOf0Dzn51d+d/R9l/7AeiwTvLpi7lQt6H2iwIMizl+I
LhreCVZkxPzt2yedzwzelvzZ6hAOiBWRzNfWx2QTyTg3WFvnM2Voj7/I8upDKue9weYm40fWp9qO
sYFN1I5D+VvovCBWFWF9RDsc0ZhyG9M75lKYDAnop7gzk3075zDVNMzfuOXlymOXqCVdYWHtRP2T
vJ+tIznhzMfNFlQ/VNp0h2O183X5VmF4IG8vTSAtNrod5rzWYJ7pWMjix0yOric57Sr3l53uwI09
vyCw7ggTXgduuP50aoctDDHIyo1ap+RaiTJ1Uwp+CBJT6vmmFUKTfBCCDzQCMR49RrVcTl44zHRX
Z7JzAR4KS6O75N9ZuIMY5LzZJQ/RCqYL4ZBd79YxSOW7Avrn26wkHyBX/575GG2iljbzPVCjln0j
XM3v13FCy0X81VkanejZaPFFLrfxJXbxNCfoU1FYG/P2vBFHaWlbind8/2WcYTtXH513yXmuYhEj
qP3dK7TgNGf5KQA/tabUJBAXos7PRoTJFZTftapn/ZAPVjkysUHCon+crKG/ITbey1hXs/oEB8da
OMvhOkg9cyiTylJBde/5HGq3VRImJxrVZWKeqxRJOQ4aDgqu2LGNPJ9SfzE1OOiMvdq88JcFFQBT
cC3ZRK67ERhuSrYrmgF1+LBHsuj65MmFOl2wdheRAdIVNxPEzwfQUH9FV6H4BkMSAI406mqCO5+9
5YoHez8dIrRQdralEZPhpE4GfmzfmfRX1R4LxX+UcIO8hAfvy5oPaCyczEZi+d87f0zSMPqfQbLr
POJ3RA/EnVnyw7iETigPmt4/pN4wRdXrTUUS7mr0ZoLY7m2eoWXEyfNepjAoOv12EeS0uJlT1HiP
FJezLUtFr7ZOKQZc/QTshgDplu7udJoIo7gIT8w67rho/kDYXFz+/KdAFw8CkZb11z20+zLXCoK0
Kl21e3NLzIq0cUJn7VFH1LWAGhd60/9KhSpiuaYJdvjoYeoovqNnIWugzRmFAlm37mi30bKmGY4x
g5yzL9Ldi3pwFNLJ0bIVLW/31Pvxfe4y3x8IE1lhwQMpK6sOfhRxBFsRvfSsKu6HutUsx5Ajkk52
bHzsh/BpZTJo/lyg3oXAnkuTw7oRZefLsQ3B94xshypTcY/PpicZ5/N+PH5r816osPslABdLJmzz
8f4ZoAkga38GbJ8fh7XSnm0jCK9u0h8mND6Ew3B2UWiAxv20fZBvWKb+DJrNPNv5NKfrKzKUM70H
S6dcNH4t80oLEONpRr4xLtvJBEW2U+aci7t4mV2TDBDrV8ZppFbONGE4KBNl0/npNNqBTJkMZHLA
UtS6EA+AZsgj5ez4njB3PKFvMXnKZzReyLQhPF1QAIkDRoZfcfWCfOmiK7POht3IXmqQr30H/82F
6Se6teQ4bB44II9jei9K+R9oos//Vk+mBGT1BhkXmsO3MF+/XUEtiWYW8Kny/QNpmet3lUw6jxfC
YymM2Ome58kd1E078GMhz5l0uPLz8/4l/+nsS7Y/4yjlMQ9ehtjujJasWhQ5RTWGwKEdz+x8IKW/
KqYqqkf7TUabgIEwFlcf/ke4UszwX/YhHCxrUtrYUPwnnJP9feyKlGCMXg1zIK2e6AY5HLjfRaQY
T5cvf1H9FaxuXaGLWO+JwbAHB+mTnl8GygYSKED8LffTvREwrA2tJ/OaD9RxmKvEXdYAnnh/QyFW
1dyIeRITQonqy5rb4+gAUzw21xibrsMU3ACD3I3cTHuDfQx90H8Ft7rPjhpxrsQohSVDk3eNADWC
G3DqivyR6kBBWV3sycVJBlh9ECRxinb6fc6gJh3wULebXFzy5hy80HB1e+5+FiZC68egxxKioQrK
FLg3RIN4rdMNmEOk+Ikn/TLMrFD9DTFxDme4uslo/KrZe3dZ2tOCVe6/WPkkOQwt5perPZdYG9zV
pBaNaTdO6alr86H+yx/KmIm4ItB9UU5OTGK8TM0UHclFKo4EWaaRtQx06JFJjSgBzKV9R/PJy1kI
sV5Wsq//wo3CH3EVKhaQMPxWm3Nt3ACWiDDcS3x6EzI0gjBo5yjZJXf0XlX1nuSTbE8SVu5kx3+W
YF/3aTNlgrfpaldJKtdgg1+FC7VygkN8RYfQ6z4q+tLC4PLM0cuOqKv4X8sJkEA7FTgd63mo57W2
5U1ALW7Fclf2SlSgHiEMDXaou3vGbf7nHC7zn01wqo/NRYdNhjeY8XfijNW/QKM3HiMM82P9vJyC
+wGu0ZOg2azkhybm+8QC/jYWjmiLPzIH7bKpcsinPOWwuHuaJwa0oWViLplKEuQEvSmz5dH+tBtO
Ge+9CuPAxRNc2N6lqVwAniMlxP96zTYVFU0WqG8SUndUQaJNIPPm/HqQ1ECUcadbgflpUcsxB+NE
gmUJ6hyR2uK0lBFN/fjgxGHU4Ukn0nCV5L1SgBXkwuonWS/UnFo4h3MEJUSyXYNsHd8FItGG+Q9d
edQoU39i0M7+b5PUXXQ2ze1HnxHyGEK3kzN12w8yYio0JE8GtOwbB49EQ1IErW/DRd7uPU7vRbzS
vx4hyNTuBgOv/rvcaUpivPOSt9/AOb5prgfelL87SN2byGWweWfDE5O1L5gZ0uyuqnGw1pLBTXKb
N/HD0cz6W2cueAwm6RsJl8rM/Na30a77uJPfzsayISuLNEOpHlaflhO5vXt+bON2/PvXBpziXoTg
OMKYAPeHWeDR4/KEMt9zORZtpgVpkls9BANrcmPDztZr2La2r/rXK3Dprkdkf6OIzvlj9F1VnKpi
NocQaiJVR2dvI+s+qLb4+ZiQSWKkc2g2qapP4diZrrnMLcmwJlWyqmUZ8r9nhH/sw/VWVtQKPiUO
dz6aHaudFtYg09fvuThYu/5TadFUbVC0tunRhiJ77X1eSMs5bxPgwvB58a2IJcetjxT2Xn8Lql4N
caFptN36r7RRQWDru0ZUlTsxd6pYrVbEinCdplI7L4OKA2S4qIrlQPrNu3Y7mGIuBVBDeU5rSsrV
srOZVJrgRnO5Tjb5C1xMYvihML0cDAOhCsmMIpbIpsJjc6vLBq7AeRE0nkV65H4RKVgJtEk9DDNN
Nw2+moWKVTUDKI6VWWCUYPURfyVmm+k2Nugj6lf2+q7w7fazqWzoDyDnwo6LGn8KWSsgwpRBLefY
mvJHawtdXVTX98MqECw0c2BRT4T9hdGbSeFed0vLM42IWqzfgPwRuo9nsQxHIVk3RctCEDq2DVXM
naQ+5EE+UcwKOw6vOQstboM45N64rrl6cSX7tONq41iRoLNAHYEQpiNnihVEVci5QCWt5X8EeQtH
LBoYO1+x2/MsHrBcWVG44WXcSt0f5Xg6/eKFiuC08Xn+fEq1nhcOgsq/eZoRiYQj/xvjoN/AQDa+
3erlh8I9pVoDSA0AsPQomBLKX4zPYZo2Tn2i7Dr180onW0P+cqJwAf0Us2Hqk3Tf8Wd0MIUHH+4Y
YuYmffKj7o5fs5NqBcRR8jY8TbTFFtbAYd4jNXdvYFBc+a0pARcp8k2d6Z0mfX8yGDHyyuEkF2tx
sbLydnumH8m/EkrI/Rmu2z5vu5lnl6BF+eULP9NwoteC5eIQa7pdmZaOen0Fc4BIqb8Dahrk6sKq
KnDGzH6yu7upf+rCuy9uY34k6v6dAvOaEkRn2XNTuJJ5aVl0y2CEkvImuIGaf3aH2vbOVAM/d7FP
AbKgx7COigfDYoVEGPATl1hHzT4uRksc4Ef948n0DJiJcLerwv6p8IifLWg+5Fm3Wc4eilAfPgab
yqImL7Nc1hrzOHScrsKdX3FDbbfh0J+KGAE8e39woW/2FixWKrxJM8wpXmBuZQphLQhu7deKcFO3
/5hpyuRkhCdzPURzCgYXkspIW+DglqlqLLMUOeNbxDQdpbGCU8n+xWPF5z6cZRbFo48QmbEZpJRb
Uz3AKfYqzfPYgIyxufpoNvvG+QnCI18s6MHQafLU48POXS/bwvCc7gwBlBvgpHoAHsKTIMjpcVsL
6FZCALf7CnCaUIA2O3cY3Ba6urB0bfbrrDzeNZOE/OQz2poyuR8D/UmOxYsurt08M52UmB3yi5KR
Sh/35iOxbcvotZnONDSXfFqVaNIYeno6NdzU0ADyvBfBSnbvF6ksblhNODfRI7N1i2ss45k2VW8s
lHHp8QKnEXV85AfU2Mr34MWNZF57qgay4Q1v4Sm1tERhR6zbvlQa1FMIrdmXLGr3zFkJCO0+sWLX
7EeEPYbSfNu78poiUrAsFB0iz+7a/in9FM/1SitlddwkDYG8FR6X9PTCOzxXHRW5S+vkwSTu1IFa
woN4n5sKCtG7HGjsUxKPFyv6sBYQ2LBglMG9oT0HBZbZmCHExExuc9uz+oljQ1lfnnRHuTktVz8+
Owk4FL6Kcq7J8oWvxhGOc81dWx4fxchmTq1bYJ2T2b76gdW2jW5PRaxh9zZG60mvhmXYGatyZ+sC
8NImzQ5Pu9IEH/w00Jen5rnIv5M2/8kjwT/f+ny+dMV47XIvhMEmVghllOTFKogBpqML+nCFl3Vc
5/eTV5vMxMOtUCwf5Zhrxe6fYRLNVANyfn2YtnwXTppH3ZsiJfW3hkPtKlw2FcO5nYaNHwg/mK/S
NEiVO+ZuUzjAtI492bQJJchg/45+5Ugau0qU+j613FMypYrtyZrrCRcTNUulVHHEBHLdUvaNpVEv
aKHNNwA0/kw8/54vd+S9Czoe6CxRIkM6cfd40KRDDFbGhRbewkEXDkglxIaksurFQ2P9CbS7/odr
pKCJSdhubTrVh097ZsPqn648DmHjafvA7BNZvmOLTydgPTiH9SFXsctmKDaR0fIUEHoYZtZr4KW4
UfWn91npdcGdiVFKFzGFEiu4EG7WD4zynlkqRJJUV8iBOfeKSlAhame5j0leQuD5kxDZiX7gu46I
9gq4bzFAeENSKHuLLxgxyGTrzpFwNU2dc/ZM8C5YTn8ApBjcKrJlMQM0KSQpEvHLUWZbgSS0WE5I
QowvuLjtNoZgUggnkR7ld8DLhvLVQPEDCopDmT5ZW2hr0tL66+bVRc2xBjpLhDtcNRdYhZ1Y78/K
iske2MgdJjPo644pV0gGZBezEN1FcTwYcVj6NRRheUS1UpFBDZPkktTV9jGxFaOxMMdJEVh7HzJy
1foZbGZx6BcxEe2wwVEq3qQoLlJJA3h156Oh3qK85CaWHc/4Pi1idWcWN+HXmKI9QiPHT7Obhfnm
NOzjlWiKzUneFDZjG367LIByNhxGCiQgyBnGtc1e9dkGJBaJ0f7dZegcW2s0bCHjXM5qaThLhjn+
dNZ2Pp7MbyRxnBecVPhlZIqchdpkEGKxvDoY/H2OQUcdaNz449ZeKNbo8zo1qV0gRKD1l9Fv4SsN
kXjEp9pk0PBn2bMHxdMzHulHblazq+LY2Kq2YCADFXWYDAfbFI1C54cCK0Lv7ALzXD/sbmdN4iqD
o5uIIF0Z2/sBu9X5rIUB0VMTjTZk6SZW9OaAcps4/oBacdgXMJzD2qAV8JyUzrk24uBAiJXv3Kqe
qr3ozIY6bBM9ILuriAWcH2LmlUDCXZ8nmsRC45ET3Y3mqBuRlaT1WKMeMTsH4ckxP/2Tx/gRv8L7
3DOEVWw8ZQqBt/KHTawPdUTDkeDCEjU4aeaZSLyttvSv00yqzB+XOECg4C/SWG6LOloxKyri+19F
qSM+QN2K+kBiIChYMI7qWEtddOKAcF36KZrm/L9hWLQcePYzBzFzqPknmBdCP66UbY6osNkX4mvF
yja9Ai16j2J3hn/FGKXF2WwNcDs6ihmRDpSRYzol3iL4mt82K5n++fIjjpwLZFs0kTnHhG2Mrj32
QsxaDm3SYdfl2A8BdTCFUhRMMZimec8cSE9oWScXV9FsRyPwgixnXr8vzLo/k6ZyIx2sF6Yxu2He
WtONZtwpsWy+4rw8FLnc366exiozFlz3vL6+hlFHJvT2iPXmv3qcjsgCmKaIoOwbkIYiseKN3Vop
JogbNSP7VgKLp9eESL/M1pq1lPXjQAJIdGHrcXPS7NJ1GEZ1sOnpqHTMSqoAXOxFEpm9MgYljiHf
OlkQGj41F8UGg91Y9TBqxzZZ49IQNKX5OHNVNQ2UXUQsMiznqyKmrxMRPeSZTUSde2pRv1aXm/a/
BQcL+W14v7eaamVRvP2Pto1MYEncQNYHt/odkyKzETketjsdxkYvazJftp/M/u0aYVJve9YMaD7H
0hQjF41Mc/JUJUy6KXJmAVjrlEeCXIB0GGWcS6lDTIgFhbnwmBAa5rQ484iFipWKeKhJmghSv0OV
yvIFZasHTSLYZv4QM1d+DRegj3eEG3cNid/LZ8EF21669EO5qQsSG2RlnfA8DpOqD/4LQgJPrAMr
I+7MS8NEHPxFieSJPiYaKbsCEsyhGnnWcT04spP1s9wn6MUZ4tZ7R+k02/okLv2X/0y9ocrYPN3f
n85sQwT6IQ8/Gv99ZDYaMePaE+aLnyayS0CmzDVzdtsFRSUaxInKnxv8Vhye5oJGK0Oh8LJ9eMwu
M4uq1yKg6hcP5pQoDHoVJ+AQLWZDy4Q4KETgNozKlZti4lzGoPHgMzPxEzjGotJbqoLX8NfEB9Qk
TENUnkEbGNKqPNeaU3VcVLi+BicXrZrc5TVO6DtAK4aX87HpjSYZzPIUt8UMkgQO7bDAAoYYsm6W
Ryo/u6G/Bai2X6O/Eo2Ws8Jkw5bKhvp3OCgQvrVElGM7Vyy+clOKb/4aXVtij+8nn91GkQJvi3wW
awr0J4V5RgVPNgPdzZFnt3YHjpCIZxrI64A07bLLKKvvhXBYsMI9Phm4faykOmdbxGGjWw3k5kZ1
U9N1bH4/oSYC2fAYUSStmeLcISe7Z51Ie1Jhq5LqHZr8g4CfzRgbfkwy1yNrDPH6yb/+8SAocXKf
p3SOjfCVyY/laLnt4XGe7eovOJ3atU6tPSzCKlaKuE855Yv0XwDSO+xeXkEAjcCuR36jIr2Hpu0T
awxijG1ej9pZMP5cK8GFpvqtjyL8nP9nYf14rfvoF567/qQrn6ef6BWN5KkoJrE2wltHVcf6csL9
MUZhdT2tH1jHrl6SITf6sVxQYfV0QBrq+Tc5uff9mGsH5xtLqEWJfEJ6tebL0JYMpBS50Qtt7UKB
+4OWYksOsSUppYyg6+JdvHwlnCQc22Omrq1ZQPzaqUIpPEIWOMdc38OxM54kPELDaR9Nk6qKPSNk
2lHElX5bK5elcZY7aI2Qi1qvDC6CPEkUcctPLQycgaZ8vTnFdiQXf26mE3aMuORXd09+el0Mn9VH
Tab+SFDlTJZMFM3ck+Xmj6TqVlvWhGXT2j+obnOhk8WgPA0hGcQ026ZUFuMBotQkN9GAG07NMq7C
oP3u9196SD+yh2g617jTRUf51fQr5aQp2oJJ7d2jmqtRyWAyzWbdmuJzJxaYzFieYgQm1MJXaDHD
/vXcArrDTplCmGVZfN9sRUlctmAb7TaeBGKMIJjrJUW3dntX9M+J5LV6UU1ovLaM/J/frj9R16p8
46Lm02Il2zxYMzZkxHifAbR2ubaOuyuq00K7eIWXKoyVRqRoUTFA+V4RyTKb4nhYEgB1lCSTsJtL
l6YNpPXo5Daz60U6b++zM1fJ15Yb8NehpYHg/bI/3TlWm33R3gQJFCsrhJ/LNTpRYzV8aIHyTVgr
M2usDIN9kO1aJ5UBDYhoMN96y0ce+6WxsTiW9zL7B9onE/JRp5pTCWiWWN41NDnK8pxXkBjxthtW
NxTkKxVEL7SCC0IG+q/0bcPb6Y3hhyYPqM3h3CNg2P6U68lCGjHT8seMTKseV94We8X8sxIUvisT
zlhN8QPn9d+dwB5mfTzM+BP16byI1ajF5XnJcRqMEI9mtFbZiTglvFpjA/v0X2KMfIFjN1u+oN5n
YgkUPRTWhHhPPG5h9HknvbQibcvB0I05h4+i+wO5V4MtYCaqMg1MTe119bi/zrPALm7okE+lFQPz
1cdaNoIs9EhEEH1G2i0ZfB6yMGVp7ICCGTp+x+9hApgzFZaRzd9Xlrs57CwmnuJ+EVL4tSIDk8VJ
nDp7c8oeLv5LGbYqFSrSRfBN5mowGw/grPRCXca7jOu2JqzvY16dpIC7/NI2EvJ2YWkCyaOCt+uM
HGS3FVxe7a2F3FQKhDTc7C/EVqboUWZOZ+DhVxi1b5T4F7zhlHNoIO2h3t/BxGXEhEnkVZ4obUPJ
OSA8as2VJ03M/LhPNUdA2ZYpO1L701q/+tULW9aEnJwjdAckdDNZz/o+rEUmB2WjFdEF+gix9SyW
QUuFy7si5ktyO+fTT/2YfgFdQMZHH10vIdXbhG9IkgzQ3c6VSHQ9D3Laoi/55U5tve2n7VAth4eE
ftuhXbldwYCmorXW6y7qM1dcoR72VPZxNWso+6N3Ejs8YBW5p5ijBVz18R1HYV/X7jf7EFnBYWZu
/NOR3Kp6d7b6eI6jRczvc9GNPm18j+wXzAHK5Bluq3cet1d/BpZCH/jPU8CaELdAfI1cMlvezrO+
fSQs1DWYTXBHT2396GGmEvAH4BIzThSmmGSLMVxfHpd7ZmPrNFS2WfSKcegiXI5KyvNL4i5LpazK
XNA482hpoSHZd5mmnCI7E4BbCeOblHNTBGyOsB3AFwCQtMvQXxEy1yKnd1aSbvGvq7Xrq+s1zDTv
beoo6eopbGl3oPC/c7MqhPybY4B+HhlgiFsjwnaVcFRFH6k5qNs7fSOpXalllVlaRv+H+edLd0Xt
ugGZqgyBSdWZDyQ5tNv5jr888eAJjog9oz4cvic9yAtja6nb+Pbuapg711cE7regUwbVRqkbP177
23RqBCm56HiAATCb9HceE//8/VZHAMZsCdXK8s/Ex58f37GJmUTEQsrCugDQiZmMFdKv2Od3kbYQ
N+O7kNCpg7Xorq9LwdP/mlHvhKSZoxKFPha0TjiPrJST44eZLzgZECqfro6XxzB6RESOcgJVe4lO
lmnEKOxTcpzpU49GsrqsYWh7EviSM2/1EYQyHmOs1m7cY1YGB9qD8Ia3ccE8BXDj2Tn/UDm9dUYl
Z7IuLoownuYbqkfj+4mIhZTNxTpm7sDoWpKDLDs0aC1Rmsg4C9eZ1BV6BSwxxJPpnqRlteYM78pj
Glg7X5L054y06xqPCb5Ica23MdzpDP02z0LSRgSN729UXWM8ZTZZq+6wYcJ+o0OOpnbtoETzMmVQ
aLlaAfkoBE2olBNxrsQvQHB3iJzIYBHCWPMm3TYTd+LDxnlSCiakTA3WOTWBdA1EgXuAKZ27z9eu
957QwWHfld2+JZw7SQa7mJMlKM9uJrpNCXfj0Ezpq4LrQniCusIhdZSiNLgIcQxAlmLdd2Umyqn7
olwuVjR56oLWIVMbyFuuIwWrucU+TGYzibVBUnNPokalc49855DZN32x5gBuFyA5WCgOUAI+eS7p
uhLw3WKpSaZFu0Wo6Qqt/GBRKz5RJmNz+E64pKys5j7PQYG3g9nkhXQJH0gaeTn4XJZrsLKPg6tS
sdgBRF4TpkPx0NAujm6HEW4nVrKEIazGRnggtDsSdAY5b5vrgbi4qNOj+KJSBIlKKJUn5L3afx7A
JntKreRmTHMTL/lXpIUIK9BzWP1DxCp5EbxuYVuF92jTybnhVNvqHulxWh0y9RnZW6MJu/OSzeyq
V92/4LhVSCQpDb2t9oMg6dO3cRIJ6OhVqK8Ri+XtKQHZF3D6JnvQcPxJ3RuaJ8a0tMBbGbOWR5jj
fbL6Td20RSD/syPjV4otw2yAdyHmkI/EofnRR2K69q31o/aXZaQBn9Vs+8WkQxPS0yO/72HF8nei
XiZOdesAVRsiMqcoVDm1SBi/bMyWLynylLld7dokXSAlT1E/6eDqyrIvmAkvPGM1f3k9XrZ/eaDM
knLXVALoxor7i+yM7L7Hh/dWcJlbZAOtW3rJ6+RThX7xfFd6T7VRMJtuY6TW3sUh3/IyXLBiO2Et
XcdPKTj15d+gxpMl2ki5pBkT96NYnvOqz9qYyDvPVl/oewfbVxuI6fhVbS6Kq5yCcSBzDsbnQt+3
x5Heee5WR0SZGiW7MvJ23/WcVQDltIxam1sOLUMo6+b19p3yKlWz0eRFGtz/s63VC2+EWSDyak3a
SDBcuASK0bJdmCDlbIoFLLnRHIzRI8TWMuuOCzJ0m+FDW+BpCrbf688EX7Tyte+kQqG7PEhyfaLS
Sewz1ZtM+yCDCwtW1ZLq99sy+dZSPx8rQBO27Yvbq9diYrwbRKEkMYqWXTuXwHDeG071FSzuJKef
g5SKrsiRN5U+QZareAAIm3CKa6CeVJVvWmz8h8j0aRg6qvBkVorlZguDYTOG6yWJo8sHijFSO+Yg
hcHLQc5pPQ0c7/cQx5+2AXhvr0kqv915onVjV+Ue4vzRrL1u/PT6PxhXQA4YAs+EtNnJCGHdetcz
R8PXxeg3CI1HqcZUXMHY2RQn6ags9Px9C7pKk47zqp4GCYlgUdxy5vqZBhsqjfWHk+ONVs6wl3Pm
8OtW8mjBuLJ/KHpSYMXL8KTbgKPgXiyFqEFqhr1ZwZHFzSSf0JGtrJ4XltAyvGzz3+Jgzij0gx5h
A3SXNM1pv7l4l4ILS5+IvQ3qUD9NELnEa75jQaYe/zEMlC6c9UJvhNahSF1yZoAy0enS+fJV0fos
z+Mp5d2LZmsHVZnBdei4BGvtTyDzipM6cA1DGXHSF2vHeXTRWIvGX7/kFE1xSewsFt6RN6Ptnncv
0w1YLhqTuW1mJKsmBoSGLFnw4qO3XiF9mJf2l7SzntQJkPqUyZWTTHVGtOnS6kCV0CYF2ZlrXS+C
Vl9v3famzEQoTGXp+takHHEQi5Enl8XC8CVNp/GuTugxyZNtNIk7uSQLiNYDZFGNdyL+wn9jSbQu
7iofLGHROQgFx1oXJybRIkbWvfVbo7dJEAcYeabSOyKOmllISai9eELAX4aFCRSoa4jkoUTGmH84
Ea0dgTYT7bq47E42/gQ75ITiZGWqX2ztmau9HDn6Drg4rVnhTwVZoCt5D/B4xDE2pai5WBdukWme
FwVlmExBinwrefl9EZtCRMq3aWD5OV0Vz/41RRrDcOr4SnlpHNG4mlSrWqeHpxBwGJXbOig5f1jk
gXC9u7RMK6q5mWWSInbgZUNzaNoNoaXpq1b+hd5FkIZvZig79Aex6OLrMggqUwZc28bQGrxJOjTP
A4DiybqA0bEpgZwTrKNpX7SN6eHpsaLyHMOK9N6NYZSbKK0mH+mu+ecNT5TOvisq+nvtG7X5byj8
OYFZB94dAA+Td4MtUFApmyPd7miUKMcE9I6f4HUhOqsGwUA3ohuRIDT3boUx9gwOBhNbGuTRaZ2T
qpO83WTOw/oC9SWIQjO8z3lxAqLfr1+rrzwVdeH2XD4SJyds49COtZqUy2w3A0Ws/n6omjG9jB9d
4oct1iDcqRk+4EANwZL0RmygQmXJW6/ZfzczHJo9kdzhqM9yLZCZvE385dE0E2+abFduBvzKI8Wc
d3vTjhLbzMI24Ily81mDEwQDVOCEv0NJQ9XqLZOsQk81ycGB13KKIQ9eV+BOEUR6okt4tuKoHZid
tCZgGHEl8LAzVXJw/uL8/ODGdUKPhjeyvEEmAAIZyFLlAG3KiAz6C9s+vwABGGYn5+3I3QK9FXvp
IKC97BgcpTo5r9EGW1dNu2E4DniRuRHpv/w8QakmGOkYpyYl6y0dXYyMrMxdCVmPMDEfmRLZBNwS
I37BbjqHooJGF5WbzFWOY5d6Lv2V+F9sTip30xILEZE669J9JZ0RSyzLgHlCrVWvrgnIya5tVwLR
AF3pqJqqx8xA4XL3+B/COm/pBCX4vAoC5k4rw4pb1cPAF4bLb3kU2NgRgH4OnNiPqFkO9nyj+4Ed
RpRRUNYjvWatvHwrL1RmTGvsldOfi+gjGMbCjIgWtg0Wxs3Dn32q5RFDvigyOCJBif3+P/grLYJa
OvDH6biiavJAZWtUK4IXy/w+a+2FYr5IiUmKkeZet2wkJt5QbB9rl5YE0t23UtTktDCoOhYIjx+L
2khziR1rLkcEX1M9Ue69j9JUDjNvMH2/7b8U366HjqMtA6zSMzF3Ba4pe14ztxlXIoBtr1WjwM7g
89MT5Ztz1fre20QtbLirK16eimVpHduZ4DOERd17RjLRMAKSI6COQQVbSLugcR6Gob696xvgtUvv
s7JHPsvdA2QEq4CkgOCrU3QCRD7O39hmif8ECk5bl7+TlCbj4/cCOlbRIvT7LpYv5+p5NTH0eyal
t5sGvjOb6kz6+lGP5Q05Qt29lPlz7ioh5lWoozk8v0Yp0Rwt7GI7kqH/ySkOWz6eKEjMNPXIGWMa
iqZesD5paowuoJMZ3KY6EB30Te82hbJAPK7pK/RCpCV5NIoklGYrfU/du4iYi2X78rQFeczk8a1Y
S+lAsVgOSd5nYdQ0R5Qz1FfiugEcx5zp8uZ3LIVqgrBCCmCi2NZelLpRJDaM0FfnW0CiqOmC55wc
OquzQT1qs33rvhFtIIJWYvOQVkV99ojUKpU269uvMt8ogRfE1/pM3qCqWXIvWprZCCVWM9JQ6Deb
4iig7y2Nv8BHFh6anMKOrOb/tlgDvJwk6st8aeTe8+ajPBsVKVZrQqTHi/aAuznmnIJ+eGPIv576
zG+9TXnIMN8Ys8owtwaFMMMG9ygZpNqlaRCuuysMdZ0y9yRuC/2o/cUzuMwMGIo7ETV2D0x4fo+6
M5QFL9ftt87dCdZh7CTzwJ5v+3pwtKohdkuU61wJqm90knm77dLakcUCGruacm3A99VPmM73PIwi
TfLLQ+Lcjd/p3Sl7qC52ZkGjXFgfZ+V8MBWWGb78WsbYBaZxQwZzMUWcvnA5QvGSs/XjLXq6KYCZ
9vbzVj6Hcoqh/AIjaSOhkyCt1GI3eo10UzSt2bvahtDmD0kH9YmacWpGL5iYDWB/fqlqtFUHE/L+
b9KEdDaHrnSuyCRcYOTbmutyd7Ij28YPGUjVu/NjI/u4INZVv34T7zJ2Rdz4p8l+/0iniOAeViwS
PN9UyOdV6b+R4ST3hfES3r0f9ZXhfcci9IEo0/oDtCf5E5EU6z5hpnOpccUS52a2E+TBTmtFzuZL
8/syrI9wkJ4MyfWX/c+9Al0+60Z9B2W8syndxwTzmPSaeGl+cSpnxgEK6/45OheRDiwUWSxdf01V
ynuNXGez2eFK+OE2+EhYpZpz3gRCBx+/Zk/GJGjM8Xn7DjBn752NcK7wW5jvCs8GPoxdFIByEpvm
4NeaEUCPZy/ImUM07z1KPGAHbHvrHZ00aUx0Oc8hm9l+vjkSpkgLit6pzu3eBsZbW1RZ5k13ddpg
dHyyEX3Xypr5Vr4UJcZoIs+asRwixDxPdfbSTZgJYzVIAez6yF838Dx12w0eS6U5sy2mTiIQwrg/
awfLyfwZ2UexDY8hCw3jlTEtXmi2HOoF/dBNEHRGudhKlGbqXmDv6uwFG1f1NmABUcptetdqID+7
7ZYu/aTKgSYNR7LrmBp9oDaAQCEfI9E8vi7BdHD/OrffqEYXiiEEO8FKFRu0A5wgtcS7Gmo5Aqta
0WkxMK0P51D82o3gY1eeIbV7TRrvKu2I9y6d7C8SHIo2xGZNN/Tz/wrg+rQrPbWjAj0tD0RX/yJM
R+7BtNYipDTm/jNtJZ1SYUplena6b7yWW62fm+cHQqB/6QppxSF++Emow73agBBMISNfgUsqX5MB
oFN7YgqcB5HbTqCJYtng22EvklcHOUevu9p/ooZ3p60H21KNDAl1Ol49CL/CfHvdyNwLfOawm8jT
g2El7+1WZrabKUlxmyGpjF+u5VqWDiJpI5UvL/2GOepvFEqT3UWu1D4r4Z+O9Hc1pZJVxUpKIG13
Cl+XR4lYZdI3sW+CLp2LzF1jK9zEp1wXAmbKYzI+TWGfevXVMSLCJyjKmeF3Yux2KDbzU4Zd/9V6
JEGB3PDHvjZx1mtUM4rCCBtWdf1a2t3utnfUHm7zYawMaCAdtyUsqBYSH7U5to8ggHeztvT9Pl7b
xk7FREQHNcLjVuwesQF4oJqUUzZy2KY+CnqwR6UX7BBdLCE8+LQQtWREZTLMbPW9eOfc5PWj6soq
6zSrKSKhRwHz71NQQYnRFZxFpWhbIlS9PweeattM4fUnRbjnBqIsphTb0ZlxjlxCVPah9ERBPh8J
CzZTwdyXH9M/phkeJR/7xPtn4LtbI0jF1CnH1a+mFejsTnP2tvRL9vWT7pDXvuX2J7StIxQFNRFL
c5eQUQb4xnZTj0ys3izXWDHjaK6fAs4FOCt0NaOM6E7hcRycJhIh/Nwg6guArBx5jNuA3fshKDmz
BsIFTnfikBp9ccTPKyvlsUx1gLz1tfghIZUp6FQScTSglTdo984c73lroNZBiPJTsDqz75iz355D
dePMq0N2zJJZZRgyl+jsEpVPTP4QOZbYA2oHmbgr75TlKkNsf5BqEq/Oxi22WdBQ1HEqfGm/Mp4A
dSoy9UiTel1MlGKsZZ3LHfADDJjjHWN/cOyn3qN7Q4MVse2p/20WBSlM3dNKFhT1CMGsQhzuR9wi
j6sjwdR6Tr3Q7XKl2I9ZGZs7+8mqEFSKLZoQNAPATM/mwXE904Ad+GFDCLDiv7JnJySyOZBXRJhV
ttw/M/2h2hQZHKMqidq+Oi94NlUg8xbRjlkKVXpHSyZa22dlY9eeCfkkJBgsrU27GD/cWLcfnOge
5HMYJBBE+5NF3sRlU+fZXzwArNVALuF30IPZLN1VQUjqxayMAv4rr52c9aYodUYMiaOrXVTT6408
0TowceTABKiHEN6b0gTfCR4K+c7cwKijwIKV5ho9/+g9hxhI+bbMllYf9A7ZWBKpAgCYcK/gEtoz
NmVxRiENeDhJl48sWlpC2dzFkWHi6HPNlYQRApf0fbMKkPEWSWfiP+jTO+LTFybTb3mvQ8A8DI6b
pGDQOiy+x8FHyv6p1/AyYuyEjqSgLbfvYbAwOT5xbiji+wGJjZj9TwHG3i7CvcRKr6oHVchrjaRF
fFXBL+F15t6xYn1zlj0kfCsnZ6VrJNjFgmx+Nzy67Jb31Ofyp+o+c29tF8CW1lqzPmehZeZ8aLaj
tXGZRlLd0J6S66HD0xMDAfKHy4GTw8gJE/5XFbfDbVqwJ9zMBW9v0WvNt4yWSo0BRts2s+9ibM1y
8cuFlpJj1VRR5dyYXZTn/dH9XB7R+l1HzMahWW5J0x6Cb7453VBEslSHkRGbUvDYNZUlYiw9HoZe
z/Uc35QhrJ+7po/9MiTCQVvXRYJw0IySfLa+VBfEV5mRaqe6q9SBvGIYapWAVt+tm3+xKuk2jY0Y
tRmwsYZYfR/0T5c7XMtORJX31idKaei5xA5/sbSUE7c+3o2Z86ip/2M4HbtZCdyhQNb0bFN8bLik
st66SM+jPDb21qQ1piHz7CARix99/fGobFDKmPxYGH67AMtXutX6ryeOJeBFbpt3HfypM6SBimQ2
pZhEWzuNnFzmBZf8ByEOjUHn0mtHR8CAngoBEUQEuysOX1B8rI5jdewRabiQODcGHQY9ca8WpSFh
OkAhhHmOfo2NF3SiO+CNvPeL53z5NgHM6/7WCp4Dybv7EQ+NZdeBB0S7FFh6BM3v1/j4j1LvT183
OAkk41vfYuH5uoadmvUmtSjhipwe5q39lYzCnPWeGXn3fndMO87bhPBad9Xo67jDOIV6P1PpCIBi
whq++Pb+kp/GEN08Ox4D3Vq1VtSa+EHWt/GGtiZdgbk7FIKI04BUGUHH1LkWBUOZGZhHIGEspSj6
4LCmASz4x49UY1J2UNukNskW8YIY42oU+y11J5fMZuVnFfdB6QYQgh/c8IvDZ+EAZnz0VFvba1cS
OSN1TjDtDKc/N+brqUkJ8xVi4WyCwpvgqKXuZFndmz6bgUgXQO5afiLw3sHPMvRCbejUaoFmyqNu
48qDDk9xnadQ13dgzZkGspk+w4opPoJnvG1QxZbgHzx+H0adxkFygS2DZ1mPIfRK44DPOyNtxSfj
fDFK0LgYp+f2mhAJfU5UsiezpvFmbNeFKcQwAhZE6+44qjLPOM4GAZ3htEaZR366a4vMwLOaTUzg
oYDhA44/9rgMMUAroa6lZhHSK2x8B6wRrfZp4oOuQdPK9S/qGBrvJYoe95swSVyJyeT/oGo5Szl+
XcfqfhwLrAGz+MpN+WwwmFbHLiILozYOz7aKxsIzhDNxisZI4rNhfaFRz4Lv9Qe4MKkBUdnsILu5
dfuHO8kEF8QNF4taqabv/6491sOaSNJODPrdrOH5Vo6loIaO9ocYgKkUmWnvpY8g+1kJYbIw8QV4
pKmZj96ZqlmP4MpRciIRgeggD+XXYWW7/ew/qFlcyBpXCbir5Y3dPrn5hS6T1Ji2GrMPBOtXUcfZ
HiMRyqJDX8KWAIWlviRHqlPRlTjmYrdKriNPRRpxY2s1qQX9zdGR3RsPI5gg1QH0WgnP8UFY0MDG
4lSXNZjdw7O1bszWJrqHULHBOpC7HaXy6EH+t9l3DxwoCx84laFXgIHZXY7mi5bwm2/UvLusk31h
6dftyz6jlBJ8+nh2QJz6Hr2Be0uqLVm2nXZ49VcXmldd1IduBPGFKyjEyl4/+tBEJg15Y20VfSD2
RWb8vAS/XtymYApqPOwihMDlIKGP+aUUSYiEBtI/yOMzsTVzKlJZ7+6PxQS5kFy4PPE7mR7m6JU7
77vB8wsTyoCKWpqxzDrIyfugWsG4Jan8kJIuWabOvzPskiY8zFsgiOE50Pm8Ey5/HyxCcfnU8t15
dMM26QI4wQnLijiYv1v7aUDCuwk9M2D0g9V/j9LXe/2YT4ako89HoVbVlNpwVHxuNqPJdvt5cSdY
VBC8SxKDwBLK4CJptQ0mLe4c5cVr2gkOxROf5gHzfx1939j10veChpRDCxlzWWLOBLuCBod8Bz8B
TylZ0woXonHMzSbUX72RKkxOTnc5CsoBX4005WzJUGAn3KoZl2bn73oL1Z3MyvklTc+6c45Gj76w
eTKAskpyxeMHgJqlzjtZZgrvc5VH3B3XZVihazbN6kggyIdWoBFUHdxzUHiRYiEPJF7NBFQBuFiA
JeL3mqEFxCVZjSbGDw6gMC7GAG58N403k0h3DyIkfzg1rxoXltMvgNIPloK7gElMeV3THd9UPRUV
ANNgVVG7nooGpajIq3S97fDFVzVROl1U1jkUBRetcrqVrXYRsS+jihCAvCEK8ILwPmMweTep3fqR
Ifguz3a6Z/XRfxzpEz+S29pe3t+bnRAOeIHV0PQvfO7NIhovrnvjvIPCHPwbpXL7Mjx2gL891uns
sV4+FKXpxYneFV///jaA2iNkpWTueyrytZzgF3Bxb0XyMUmQWe9mhDkF5OhanDPxdsmpPX1h4Kys
b98MCY1foR3ExVGq3v+WQLHHwbFuq00vXvKFro5nJsnwfcvMyOkW7KoK4G0MreTfymHBQTPt1Vq+
5nzhc3P/QT4eDr0qjB8JqDH/WU1kdJlSFmxZ2VYT1CuczrZvy6Eas8RJveYMh4/aaC9yyF4m/xbY
1rs4uju2N8PLdBM20d/OZyxBNIXKiZYJoFbC8LXOg9xKJkfw41m40q2m80SCGLdOW2vpKutdMywI
1ofs8DgSupL63NI2qrkK6A8pEMQPM+KJhin46NCt0FYRt25J0m/BgtFVIPZdkxiDciHAKI5Py6/5
Ons77l4VTlwsut+QWuQYeql1r8gathYCKjgqRmosCa19alJ9r8aIPNGwwfsIGJTfZ4ILxtcuVQP3
yn1GHhP+MBIc1N0CZmppx4XKd0uGvotoai0oact8O//bwdoSYkH0b9A7WjkdiLM+9ZqBK8laaueb
B+LjwYZ0Z1m21VL3N+WCCkPNox5HhKyvMxbhK1jV7aQjYrdLARLhtGMiUDH1pukx3+QQ/KeVxQ6s
4UPsH99LGm0bBGpdPRyQvIvQFpAu+VOCTQ4MDkNdxpE0DWIImZdD6LJrBlgpW/fsyaTBQY7DmWme
HE0m7SClxUqqnlzNEZiLpI7LncB1QH/TZgiyaEIpDlC8JQlsrpDtWGALbewTLNjUTXdLvzaV6MWe
L2nxPrdGTli07A0+svrLMke/mWy07VfXyCKuScRGk0gjcLuZ+8+YEKWBmgiLVlvFzeNWj9zMgv1K
q5EAutTZjLshYkwrtXEx6sWB9zt3Ji5AlpB0Ojc3ba5HQBZemqBpWQgAzvV4mQGWzTR3cqcPYP4s
5Z2xmuHhT9HENlMrLXIWLmIVfy8g9mUG5B8pPZTBdtQp1MDSI3IqgwJQ1FbYrtFSmBzkJZOJVsDt
4MOTY05n70+XHsvDpYatYeDTT+Qt1KsE3/eDR0LWuFCyYh9zPrNegMBRY6vltiVjfdvAyNmGi7cG
I1fzNUDpw99VzwY9sJRyWbBfeQyjQxpiLep27yw7sxtFh5scGcEVP8PMIyygo/GeVxhE3f5VT/R4
w0iV6e0b1TX71sZWQdzdPNZL+CjC2VSYVhneu+z0iXxSW/QN9zV1F6ST4FDarkMZB9qwyT43SDKr
z090zKWa+4SVx4UGqnr04No5aWuVBCGkw5z4XKCJbDdMa74+hv933PoD0UxJ+r3L0bqaQCScZJwB
tEEHYldduU2avaVD6mBV4fd2vZ4Hy2PFu/l03dw2tRdi+1MKauC2xOR9BYSILN5Pol4r1ozyNXzl
OSIHg8sJOtiKA3UvWR/q5yFVSiuAXll3chVvWcffqJLDu8Wqoo7iDGSS/aJLrROkD1WjGUc9sWUU
SscWp6Sx8sBr0eFoL1Pl2t2Kgo1kT4i8bVUuqy+oC8MQXsv0ERXjUwGBa64w+/loE+ZEzrbpuICz
xydOK8xPnHs/zl5r/pFIw435owgDYDI2HXWTVm8r5OT+lES0lCaLBQfU2iHNCvX5FIaZk4uG/qr5
o13df5JQ7BYxYTo1g6qs5IvO45e9wkigvWAj9bwlnvuoq3vgLJ0bHaMpfTGs/W857DAytn9W9XmP
mKYTQA3KMM6YSmgHaYZS52xjk1c0O6CN3XGvum09xPExy7qLoRGGmCNdaYi0GNabK9X3ANvNKpEp
/1VYzX/zbICAkMu9Yjr8SiukTG0reMhorRyyQGVmHd16IwcMsycrjHBT9nTREpj8OX/it9xxaRjk
aU0cDwtiEF/fdLcRg+zoF9qoqtzoF9wC/EJaAHY5MFkssi5Zs08IuG0DdBEWfRzWheFjjpLf+Z5T
OBnnktUT4VBjtpQgEcHr9NSOQIgVXr4klPlC+AXdDipsuuVvbbhXqY91uJw8H+0cARImZvjwItJZ
/ptUkgk/pco4JkKaxaoDBYgEtx/Asd2y5rQ3pXHwPjF7vjbra+9JsLzZUTK8gy61QNEw30afkFRJ
zVd7lfmkGyMakJ/ZZOEB0QJX9EYXAouFqRjFtrQ39rIGywsvfOeoZ/nnNY9uvndLgiijhrUR3u9B
VM868XI3uzjUjzHZT9WaOlvc3H30VAyUXSCFG926o+1jlOtTfPotlDyCtQXpB8B+UN99L6R35Biy
k5Uf+JukMK9TTjbzxLqtV3Y9wuWRvNgfw4Sn15RPRLkIJfaw9g+rpTlarr8dEuLkhovMvMnh5HlT
HsVCmeRWEliJy+IajajUXUlx2fv0g5ed6k3DJNhpgodERYNkO6y8JZ0xsVvXAOAUzDoA3WFstsGJ
fy+ccRIE9byb7OjXiofIFdvLu5mP+kjIPH/klFcF/ULMVgrqB38fE/V9cTNKE9Pe3LEXl6ELDNuj
VmDLnrh9y30cCpMzWfsCq9owIYOqvSH6bJSey6TTCxNOLVZpzgAxUS8l39oO2uAZxj9KLQ/1zyc8
3tWG00hjXsnZ6C2DuyuSVAqqE0DeB2T0vvUwAdGRVylQDjTviW6DFDS/Y6wHxqDZBnKhbWdMJ8w6
WZw7UJIjSTFsVu85YaevhtHZEqs9i41cJSkPOfHLw8Yh8ZqK+3G+cRj8paBgAUsBAxZAgIgKzwWG
i0SBN7bzmY5vWWNeKyMHvOXkscDGjh1OHpB9lfVUec7dupO9JVYYE5vDHbHAApFHAMxFW52IZ/f0
zrysw3TVAvG2UKdy2ZIAEfpJHGHtM5X/asH5wCRjLZkpR0xBgI7jGKK/WBEqH5zjZBZcxat5uc3D
YrPNltr8XTtZx2t35PHYbGn3bY3t7P8aClclSrXPTueY0PxS5Fg1y9AD7AeyecEaKlsRvGQu3Ole
uPYlwpyWdTgyGmaca4h9Tkmpn92clg3P8C3yEiIaCXO3lkKfVSoq7qlpoiIX8ra7yU2g4iqtlxmy
B5owYEj/K2mqGeJAXEwJcJ+QukYN4S3nLW6YTvZ3SUm68aF+RzmbNICmIyB2up+wbXBfyDDVphCv
wyb1m+BGNW1BXVMpx+aSTWtsRz0XbgTfgLoXKt8XvUOKKSuPxUyZS6KnJ1RDX6cW5NYEtUtz/GU9
2VYnjgLkj3U0QI/DW4HZ1zKoNRGSvOcd5x3SpEntUiaKiH8dzNv+OK8C5bCBKNV+e3j++i6f6PYI
crqTel1PfA6YkBLZNVxWajp5D/69r+JfBve0lfOjSqCpgXduFYBWgEbgwKL1MGUpkfAJYqSMW+Y3
YKwx9tWITw+9tu+I2NZmeiQVQytJGO1A1znq0MSGMo+ugZ29MRtdqWWEo3cOBuISlDgXNGQQTEzB
6NSl62JJjyMmTc+DszJ2dzPfo5wvIJYDfurtJPMIa9gN1XGGG/sCJ39CFkWm+qciOoyMDQqFkxnT
hPICXWfllut3ddfuv1E6hMhv8owOf2kq1gNbdvSbktL/EBtFsF4hizV+pXWd9OzY0+X0GFDDGcWr
yU/xYQnwH64TLyoHgNFst8DRs16oeZYucLWPq/0NZkiCke6YoSkpTGJON4lfqEoUXOTpqHHTir6R
88YOZ3EplPT3YTSLP3YgJpNNna4+kTv0nCmuRkZiWpNzOdiK+8ADYLehBN988UgH1xwy+sNPdxIq
C3wrxW7nSdUgjsyxikPXWLljSGPm+M5mIGXHLZPry5dsHqzBnNv4bQoThWMLugm5a9np/1/OwbNH
gU5VChCSPgwN9XiD6TEkjuUSKRB8UmTFNn2KrtD6k29AmFuQ2E2TcClzKitqGwao61D7ux+F8bPZ
MTmUfTUQRhVmZEEghyv1TddQhCeNlLs1vRclpo1Z3qrXESvPcP4UI2+rWgChVCwZtp3El16Yeql2
IhTokf3Iu/0i9JEefzhGiUX86jIXYrBftGjVHp/tOt01Nx7mtqoNFmLiQZ7kZruvYNu+FsEJhuLO
zcclF/5uQElvHnxuyJ/MdVKLdYwE9gEKkTsq2WQP5g3G9pMAMV3niuhjVDWDP1fTSvIpPfOwLac9
DwebNW/eWskCRhyMvjJgfN33oBEiWg5UxwdQ1necmqq50lCf4KPPZhI5yxFiFSr+iqMi4OREGsJy
T5O2z7bdto0hNYL+3p9kRkoxWysKYO6sa3JEMy34h7n07FXtv+mGiYzEwizVvIXmpExYV+3B6TKL
6x2pWp5onU/Q50f9rev/KRTmSx/Q7qpCFhkqwwft75LOSYdJ0TrFgJjZojl99pHlgBCye0YV/y0I
XhHHSoPXXd5LVyAhUU2mxm0MIUL65GjZw8bJSDLC7Wzt/WmbXKD7NMjeajscELDZmD1DT7ab8gAC
gKTqd4IBxhhhKsE/aLTkyUUaUpDE+bDUtl1dprJ0bGhElbI8uUMDwzsXdsJrtvu4gO2MKfSjFhVr
Vp1afrYiS2eaS0OK0j5kD7WnmwPCx/ZqPjW88jZu6EtHgH7/ln2+p81prg6GOLyX9yaNwW2Vzkoi
LL8H+VFCB5r6RxFDcLsrN3BtDMeVfZb6lASD2xtKBVCDRxk7O3vPXOB8Auimfq2nrVdLDK05z26f
Mhm8SrvAH3c76Pt/b7gFeDyAfMnGnay/hAafuknERvEGyAx9c9X+2mJWZd9jiRVWQAHoyfBEOQxU
4nvOo9zCUnrnqkdiTsAZwv83B3FCxZZr6V1q7iaKlYYjgDHtljR9gcIgoOdc8/eTV1Ut2tOSrGAX
CqEGbZ3eprzT0H+y+dZctGXZJPanOIIpz3xvm8qCDzZB29uapqXxYypgfYRTJNPnB+rckLIWVjSx
AdZll2WeMkYBFFt+nskupB04pgc+5yYjQi1d837cE2C6Q6YBAabMbgqfIfNULi8pDFqpIeI/U8qv
ONlzihWM97c/2HCUYU+2dMQvEQDpbOS308BjwIpy2A37v/R+izsTDMqaublr7d91B55dUXefNn6o
BN94iABFl2vGZBsj9OEUkHKf70rukeAC/cwzSnv9a0NRi827fkOJsCP6JZJqeJOg0qonBr32Js1G
uSCOsVEgumMlNwdJ0DtcGyxt5aVvMY5RznM3J7uW/aZsxDLEqf2YQ/VxsgEzshuuPJ8mH0OZ+c+w
boF5tQaU3Mq7sSg3DvafHv4u/SoxXB19PfU3IH1nfRX3xiL583dFh+Z7rqjEKbSYIbrjn4mh7H6d
niHNAoCltA3gnEqmOTUryocfwZjrUPbSY05GBnUpcbqE2dE7gni7/Jz3jP+QDd7KgOuGVRCV+u4g
cinfs6paaqbLm93IusiqXkeLQFRnz5nkETZnozdMqHJOiCpobRCREbmj4bSuSxzZD5FYLMSI+Uqp
XUIgYwdY6zE6p4ZEsLmlQEQXedembmHzXQbYa4TtSpbQG7qmiAkled0amT/J89G8X9lS0+GhZoV/
/GqmKhMNvCAdkpSg5bnPcnLbbFsSgoQxBx9wyao3nm+Ncyr39rnhBd4M+6tixtk+AfAzPGNFImzZ
Uc2X26JzjbdOxd9CXW12vSCAPClStY4mWAbg9oQ+b0RNTuFZduj8UG9V2ZjvxDrCcDziZo+g6MJN
A2lQvfLTGfPwYDnafKNMo6T/s69kyTPRJKqh2ulBDcHhYR5m4NyJEJnfLlhrM6+Qbzkbe9cA4B/Y
3ykPUjRVWbpvN1INUC0zYz3wuw2eDYpYjxGfluSA1N+sdkZAMdfnN3eR46D2he8MLSyGHGKmBzZf
2BfZEK6kK7J4h9HBSxgbPB0Ysq+NP+9lno+Thja5d4UanyCi9ZE9J1s0tYBJT9/8Z02G7gs3F5wz
hxxkBd7Rprgoo/Xqm44JsTLBtHN1fVx464BWk/DQaznhTQP2QjpXh/O0iFGpJmz08MJkjToJEajt
ypBkH14CrNaomQHD+1TAKokT8BmhCvFZ+eb3NnQt2OgCJWwAB9NezMaFHqg5xJ/CIiQT8VQmqTGS
BT8GFh2VSJWOJIjXOvDB3v8EFSG/ryvlk5Q4gk2CoQ0ATbi5GdIk4zK5SZj5w77FS5we7a63YGF9
slJUEzLuW6elVHUQsLBpWQPoVetNFgIpqJMuk2xfmqtnAVbolUw3NgvCgD8zgEB34aew3Jez+kZq
mB1bhzxtB6XmOzcj0DVzE3eeg+N4puF7qtb7tb227NsA6qsBVUNdkquPMs7PpX/w2rQgiAyEBJcJ
jUFCvzMg2jzZFHJ9Bu2m5/cS955RZYBEUcey0625bCv3qPhLhME+eGxIRCdMatoGwIcotKNEzmFL
g/2pfBTq35MsmyfoxszBK8EoVm8klLpswc9m0Etg3VcDZ0A/B4XE39Vqg1KtWkZhRI8BWHw/nIHZ
0v+JJGYht/Hd5Gx08wLOxOLPWJ22irqvENLEfO6kfOxttvMko+MaN5piLs/03rp3dkfnYsX4fpD9
h7KL6u/9uQMJRchGhGv8mlf1S1DjjsmmrBgkJM+7aFZmaCoywKHNFUScXHbY73LA1oog+dgPCErY
cKHtaJql0uZoRjEPMDOKBQtRnA5Au7hA90fm1lhAENIO9yJE4s0JGKeL+ADdWfR0psL9E0ngiqYh
5AK9aheMNfho7MPqTXicetxm5QnVzH7R/Ri48uuQFeYslSj2pL+is2n3TzBpTM8NFAx5X4Dj/0ZO
EfQIuy5iEsSQCIT92E6Hx7qG8jibMf1M/f23U8T18Ymh4B/5tND7KKSNh1OxDsABVtXHgr8PBj0I
VsYAGziaQPvxAOrLebYneHB9e6Z9X09syMqSHEsBE2bNNADquCvoGnFscQZLF5LNCh9P7o6DXsWI
B9BS3M2n/rbv+gnZtuEpaswoivaYTLmBlajlQsi8TvuZg9jRGief1wyoixiZPGTuUUkGQlLi+QJn
MllSMlu5LShEyV9UK6DmGm6WzheTGQFn1ZhSUciH4dhB3m78M5hjrb4BNSFhpJPBFAQQ7BR6oHAw
0PMX7Egr7dbPEKfwKJ14NKYgpfS+TZhL47QNHOUNOTjcGeAGY/ZGZIcl0teCHIw791kHqLzlrWqe
dwWUjYkEPQ3TDrS3S+8XgDwo2eZdNq1w1fuCNrsZ6iTPHHdkP9UHeg1YNf5ybIgR/swB8mRzB70G
pf13MbzLrwNwU86jDkekQx/G9rUHN08RQGVt0akJfOLIYOsey4UHdHLF4Rge6VKWSmoh4Tp4+pDD
v3N9dRcqkrMLwrcaGTAeevbjCzJ246eSF29zRXeDMSduITIH3BNzW+/vkfAS32mc5E9TTO7vfz8z
pUxd42a0/aaydgOuII+nm1f9ikafOMUxReKo2APhMuQ1uhtgvHsg9XpfmPwXjEQkQ3Ff50RbqIlH
pO2PEKwctwpB2IkTfjKDRIzjRIbmRWWaQ/2ScJq9LE3MO2nhRhgmWtki5rvB/qwLjUNdb0hki8bQ
fHAEEzn7COiCvKN2wvuH1OlDqixzff7G3HA+R5KMmG/T7nWOTF3t/d2WYgjAE93qqTqVqaKMyHuD
vZCE/xulvWtxRyslPlXPwlXJP9yxq/XwjxXENsDsEDC0ryOBYoGCNLbO2QBX4hFjr9croXWNWhOS
Y4Thb2mFAWUr0V2r0YgRp0t3NEkeuseHF0STk3wdM8PqnLAzsyU04cWWuhPCtXhyHQa4FwmWTa6P
usynk/6BAnpVyIBBws71lSQt1+vqm6UOpY0htljggjqbdYPmGpG+hO6+1Dq3yJpGSJQz4k4l7B0k
hapjPh78I6fdtGAHfm9kTDU70/YQs9iAHm0qJpWcAclQlajB1K6qw6BJPQpz4DHRSTVBQLTMdn9y
UHA4odKoF0QjS+rOF6PhC4h2BwnSke/X1TWLSRe9uIHLMVzf9kW6fdKFNwLHL+BzjxaPLRWNJ51Q
u42opUjzjMFEerkKwOF5qTJOPBv7Z6gQWe7culOJLRujcZ4GKY5dnJ7+O89rw0tRrNhdMI5szGNT
Tpw9j1dcRRvxW5U3RpePJ2W9pHnZ0Qr+XmxoewAYIX8PjX4pGVTEpxrYpA0O8gHelIaP0IEX241Z
Qpx96aA/kL8wFc5tZ8DVZ87gKQioiywyaB+FX6RAV0O8xxu6g31/rvNaiPcr2q53fwDI78U1yH9Q
FBprsh1RZC014QXOwvOtCN2WN/nYSW9qFaWGU886iXqks1wPTrD91LDBMEgGXyK+j0j27J5sFEPL
pKxFBiOaZarcoenuCEUtvnLselsxKp50Zkyvg5jCdCcdf2kynZTt0T1hXQQvM/bXp0dcQdyW9epL
mzdOWa8OhLzb1QdeOcYgo0Hn15TKPuAYroVfvySjrevgik06DRgq77qMd2SVKYJNDJ20oisMpFc+
VJjuPmS+4lIbifRYm1L2gEzMayivIi07x+3obSJ/Lb3Aa4LR2oNDwR1G66oVB1EESKUwmd7TThEo
pjsPp0rSyKQoUmcf8IRkjLCO7TZbYwbZ7oKWfrvBY6XAHWjzokCEPcq/41tmhwt45og0ItOIOYMU
QucrO9NwrK6GtjG1HWXAeXox2uhupl7KMQFBEtIAOOgPTRknr195gS8fAMniHOHFoZXFTxDUiXCi
NVMqAP5izDS3IgiPbQsrYcENSM7Mud8HFYTOIO3axLNh2pQCrHgaylHntnUYOoO2AKsms36eVLzu
+vdGHy68KdQ4pMHwJIu7EtyYkAZwUxnwQ3yD9plHzeP7t+Jqj3kTecHT0Drd3qyaGAiXIp0fjNiA
YgXY2I3lHPuDT5jkAVlbhVq0T3JaJ2U41qVAvEqvIG1jVYRnmygnso2uU8anoDhsSNSEWozDYJfJ
HXUTfW+mV/7AzpHcr5+BTEqs7PyBLKO9w+YfEQMsSK0kgw3fQbY/f5Fa580DPianG3jRHtUHcs1S
dlPKKfhNk0Z+pVgBgGOlxPOt89ZQr1eB7zF+oCr4fhw7UL9KRFfAfU6ykX3v0UJeGhT/mqd2Yznc
GcU9COaniZdgyKZLoX1k0ui2TQNuF796vcCh1a0Tdromd3ae4D5WGVumvpu1LFct6KiiFb5+WJYu
AsKJtoW/ikRnEg4ZyW7rraoSRf34cZWjTvOW+ZoIjwAmfWGXhrd7mf7YzhFtDETxy2yL0iJjkHdf
+YYAWC+Qwq/vBiykrH0KxyXJc6awlnPQkluUd1uH72lb74Q7Zq+48FGMX089XJevBr+Q6g2P/L7y
uIZGkd1KJ777wcHhJ4WvM+VYT9PrwXMKxJ3kN+6PS57eDcBe30+XIUAroC6sbhp/959w1pzXTT46
CCop3on7bb5lNKjez8rSBORNWv2Ca45MERh/WkjF5S/fKDAdrn2uJLFrK7S2eXazc2uYLhZnzW5g
Eop49H9i/e75fJe/Nng06FIIjnYVbQ7yyiafzbU+qW8M3sO13GxniZRyO/Ko5QXqLmi+YDbyg4Wk
lbLRnGYD8qyfX0OtnhoL3aSFqU4yqlkCm6u2ZofAmstq++e3z/w3rvDUVuaFQT6+kXD1Q3kxPegx
n2W3si9/gHNs6dYiHs+J6OZERUP6BV6Up/ZyWg4QqaesctPGmFseqmcVmVypxCnxm5TsvSqXSQP+
M1l81+Bdk26RbYTztfmHeCVkZAQ7JZOXY0AbGjdsbmOJ297YECrfCMhtu2RAtFA1liDpKjrpor7W
J7Bsak7sACWn3lGkbTHlEiclfpOeHsDgn5nQnrfzWSQE4GDcps5JBzJbvX50wFKRf9zwpbenodJD
ZXQpzw8cTJnab5/nRCUyY7IRYi0eioI9rKJ2UU8jhwUlw/OG9vAUl9ygSPPjyO1dli2Ze0lBV9yG
b6MwcqyKnjCTwt7zX/VHzTjyoxxmvUD3tWjY+pC1kqUagv4Sc3qnaGPgN4giLUBNHcnhgO752s4E
Aa8e8kaMdRUuwtRIKQdVvNu+rM7gz6osmeeVvi+8CRMgGWVOQVqgLhWatDcJJ7idYWFU0Ow7Reex
de2p9NUs2FX2Vt89qF8QIiY4ha3nTb6IThnuL0OLtjF9STj8mPYQxtNStuZ1wR1OfgJx9cezc1gP
vbor/ZuWYMkEw6zV8N+hN3w5+Hp8F8QaZL1pXJNSbJkSfP1LyeiWP6Os6/J/T55z/NQy/qYsHHiI
RS0yVQv+GDSVad8/p6xjAVGwKyf2RhT8+VSkelVNwm+Yow4k951Xb849nWqzmCbU62gQCP9R7vgT
jHN1tpAW/Fn5YLwNk+MomjuGQer/KvR/t1ENJKhDh1rsDsttXrZZSJm+JXjEvKrqeXj+F1XINamw
lMSkaZ0d3gUt8Ch3qkIxIfmZiM0HO8GWjAFPjUhXWuZskdb1l6ijjHz634/lSBF5JkTBYexZA0pM
25JMs0wl+4rwGoEZKeMFpV+EBl2Kovlgojs38rISzRM0GBO4ZCss/yOQ+eY1qWsPjb6bY+Tym098
1e1ViEEZA4w7rsQXuz0N+ACrySUzQnQpb43VXDpTHcCfNxNTfI/axqVHi2ofgzms+ay14tySWUoV
qnnB25kzfaj8pft8ugEvth4W4M9risS34BsalglMG69SMLDHf7fuDXDN68Hhce+iWAsKQN+mKutW
Y4BumdSsQ0Lgi/chZ2GW9LxKxM1Cwplt+PBzuETBWXUYWrqvSQTz74lQtfaPoxJFNm3YiPWSM8zR
D+nuYh5nc4vH7mhxPk9DBGoz5fkRFjht0eyGw4cjFBbwXVuFEkR0gu0reY2mViCdWZAeoVJS7+3X
avj+UcPWaIh1laEpjqZ48MCCdbQldAUg1N/M140g5PpkDfjEa27T9dUj9+b3GWNDRDZAYzQwYjd/
v64KsThFYO1UrwhA39Tby/Gk0ttn43RxunTOe18gcKTUB5Mggb3W+5bjEbt51ijye9OxBevk2G04
1t6DHKFK2NBvV75ZkUyNcnVxm5nNRPzT4dBQ9+TFW531OALEyVZ+CnX4l0VBf16Ri+aD6itJEeT4
3904ykSEePcAlhjFTXV2WWJbuCVFOtfcSbPV4XxQXC4oJEdUtpcTbQjcjmYT6UTdRKbKCNtv0u2K
5eb0hZTgcUjx/g1i5bShlhgutkJLy8P6t6Eak2LxM11uSOfwWO56kj23Q1J+D0+6P2UkpkNCXu1F
pfjv0WvqfPv8EFajzCorfiX8bfuFB9BO7ZgGUjS5MwSwzj4oBdEY8HdINkTvt+qNIAwvK52ZbpOp
EOfnOd6LgO0x9TFp97ZWQai9HAOzIjOt7dnfXh4EAd+fkpm19/bw9nt3DBYmxc1dflIBuONp9iHF
DkFAmUYuJIJQ6RdoEPbHzXD2areT/2LNR+zvcqfaFoXw3dQd2+PkRp6iBhuy+m972ZmTuLi1SpH8
AiSsfs1CditWrzAcBFzHog3egwpDlyOsDTx5W6M8QflNAcPTxiNM2dGEDgiUVI9GQUuoGx+ZaqBU
7TkNLWzzG0BW5MR07vMsqZP18qgzW7OCRPSLPU6Lh2Z39CHx8BOYBe/kzy2W+ssFL6QopN6xznwb
QZF8T8PhWOIqkTZs/Ml4M7j7xR+wTJQV6NvCrBXijkB+cLlr649U0tNE7kZJAc9eQ3fDSlQ/6tzi
BKWAwgQIuYcjbVUaUl8GN7XydYn5IWVLJzf6rbrj+8We2G6Bgb0ehempVjcvxqq3DIf/BussgPt5
vyTUMvFheXHch1yluRMVRLy3Ea86Ys3NzcnAIY81aN0n/O3BRDEuqQKxIJZNmeQbb8K/6+XXU53o
QkSfpWHfi3RKR6hUjStr3KxC22/jRaJxPRwfcg2nNGkwF7Lv8D/QR7cj+7vErQMU2/CJz/nxIcZQ
0f7h43hFxAwpWpVYXzJXvhL1y8rbA4gns+xbVRhoAHp9qOgvwojRfQsUEvjv5HnbsK6jDHsHiIcQ
9XSPDSxCJGDLaGoFV4oOEPdy8l6d3cflfLCMzR7sKEmAXjCsvZiABCLWnYeOnebhSBRDW+2EeKH7
vqlY8VXJTQZHFnkU8W7fh+Y2a5yM5L03My3Bj6glyVy2PD4fOxjx6qhJm2mCGYhQcNAIMzjBGFoI
y0YDUbWl0uoVmcI4lD7jx3Ib1uXVEe/FBAiqBMj0Se31gjTFbOqMhDfsN7eb+OWNntZtdDhUV1XT
uwSOwnpMGAb4QtAUqbDzvgAPJX30vxUWdpj+AZHYOJ9jHo1vLwdZ+7EJuu15MQqYSvNis+e4U4x7
A2REqRVF7JY8wYUepxbgIZmsQzdDRDkAy9mPSz3aLkIlVaRNsWRp3deKNmind5zL/Ul2ly20G68/
kvjp+UFjUUL4tmL+G+o3uvLEp7VjBGFdZkaYcp0lYHaYl0X3KJuiAupbCJ14ZjR1ybmK0ua/UrNV
thvdhaWduHJZZ6GeLiDiuZvECAjjt94qZjphlVjkCi4I25zNLFG8jrJRzGV5KWmUhtLAGCcp+WAx
3+RHLfJoyEKLxXzQkkqHqR9KRKt18Auj8W25paCVp0Sz3fG7e94wUTY1A0qd6l3NgvMXz/Doj41G
amGeVaJgD6l9gi8GMZ7i6L64MCX6ThrPt5Lq6vtRmB84a9+0Dy+UeVDxz8Ff89v08q932N7fDeJ2
6glCg4GxZ8pLNhGR2LCSFkUpEtCPB0IqrI8Q1/ZmhzOiXrIoDfeajqJJ1MddRrU7VrGQRxq+sHp4
Q0sXYJO7/l3hhVjgArcO5GhN/0g/e9DHtfAGg1C+HOpxpnc4fa2CB6WgHInisnW+5rqmWAS5y0Vd
sSy9si0L07AsKzRGDN7gLlQkswvVMrzkwhga9RmCGm7QrcJk+JroxHBbg3BQkddBEx12kiJcN31k
9dYYkICgX/O+X20gTPPej5InXh6+XkMsO+C1iNfEo87UMD5WSvCpeQ0qoRD/MkDYPHtVfeiwvxgT
Mo7nzhqM3mefNbcSRXLwJRFYQDoL78RR+ZfX8O5hCIRmoN34TghBAmAbrGk57q+ig+EoOySVyo94
iYzbkReaX0vkbYyFGqkLB3JMcOAWZxF1eiScrluKUU9WbtS16XrlKjtYQ1aVeJT4DDnSgvIkf5KZ
m1X8rejDm5Gm0KleU5q3nyyBvBRbFsZBT/AuXvIY+eQqHniDLLPIZ0RRvggbA9wFMrs2s2sPTkcw
YEGzQ7SC6kNrQ0BTYQMw7FL4xqh5Xpfbeaiea9emJEvwdmKn7ScUeR2BUmazAbFqC1W/z7r7s+wq
B1w7kZeCOD8d+3bL+eAXdEKXhofxq/P1ipme3p88O2c0qinGN6//Xq/vSyzWmkL+gP+o7pwPcbbv
evnwn6qABrtj+Bw6Zyx1m40q/TCIZFjRxYch+zbfJlYguLA2a8azWGRLCg8iVGjSe+CVuS9q2piV
u6f1aweJwjcDzIkNjaPERoCOtBPDrkOu2GiSrvDnIJgp5Ly5Er3l98WlmHPLz6jy0u4estnRUgfA
PdwdyNAEB8cPWIDQNvn8iW1B+k1wUDRwPpVYT/qSN4sxofQy4UHf3YRMOx/NLMv/3DUjgTcxcXDf
Sk55IMpNLKQIrSZW2qMKutuFqcAbePZUt5XxnwK6Jcrg2ldHRQ==
`protect end_protected

