

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T6wVkTPpNtKFC5HWYRGz1pDJeqROUhDmQQB0XOtYU+hhB43DLNvsfjC5KYqU6Qt1lGAhH0laXWbY
sFGsB/1X/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Bo87Ik/z3ZMfvsxWdQ0fNuP7YOCyp4j/ygqxg4KH1VshQEFmP82QDe0umsG5l9IQ7WJ1x44Z7hUv
b2TxMUXo+JqxKnlgUE5S7j3ulzSH7GuiH1ZZMyENkBX9PvYGPAoxkfBZKwYBwge7dC+ekfgtgSTi
JmblFBaQfl2z3igDjdI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OS69EpuOCXkwKDIJ7c3PBFNFMJbX4CiEZKRiPCWgGoIatev0sXIZ8vRiD53mj0pSkbBqScW3T3bf
nStSylNR1BolV0YoJstQyT1+2pFYhZ1LLXaZugJ/oBE6vqGV5u6J3W5eW2CILy6xHulOJT7cesIj
cRuZgsZzN/xmRcR/wqC0vFpdgeypXB6mda8Kpubf32Dxwqfu3L7BPiBg+o1IuskbZi2Weoc3I0l0
OeBzQzAzru491AqXGKlZ7sf8bs7SXbbzXRpVODRt7n1NjaKD5f39RasUxEkDN/Mf2io8pxFG53sn
wj8Vha0LEKNulGqvG45lCg9sffq+6YoB/PA6pA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0V7+weIw8dZ+BPWec3DOIbteiwGwG6dN9psrs14jYpdIBALSrfKIpNuQOkhxmutTucD037ovCmPT
7tzlCJSh8b8Ydyh2TEeIpJfXn05PGHs6Bho7YXv+uAmzXPPeMsLwL0Zdj9PYL8wHeM9h3s3oFmE0
whlOV2wA/y6g8Y9g2X8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LrKyoRzDm4cxDmM9WZQaVOeA1DZCMC2sBI/JOp2hUeVDZFMUfjL+9ejUV+oaV3PC9kYwU9gS2N4x
T5QckNj/uBm/MDZii4ZX6FRa6E86JES6LqHqCKy4pn+VjDJ9xeobjj2ApHw2GympzRIfTHfg3BzS
Zkqs9Cmo3/2Uv3zdNyaGnk9f0Ojhxe+EEq2njDvi1AWk3nuKPvaX2PFiQqvWXWef/JYb4HJ0Tjlo
v5y52n4XeymzBXqfaj2Y0hccYVFZ6YVhMnGGV06K68vVbtdbUuaSPRKXNa9qJHwvtspPluLhH5Xd
ujRGgNTtTMlfDYr0Fh/3k9HYg9NPc+b+y85sOQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4096)
`protect data_block
yvjZdzWUZG7TslowT38oXK6XParirjiAGUQ3HAmuqFeWQqMZA96r/lLGRp+A4WebkBqrmB+mG6Uz
l1mO1oOdqFcnWGWHqdfTtM2QR3PaVeyIPgYEViBA5MZCib0tMXi+8llN92iUn4gLdgVSVRJ+tCVh
Mi/JnTe5Mew1ntcz6UFl5tjxy4VjlSotW925COtmwJ4I2ZoRdN5Y9gTEAjQL2VrjQ50Vu/GPCZQw
dXLWPbl53dQ9HCyVgw2tqQFUrabROErJWFFmu9AA65+SPH1IveA3gBEKiuf7mx3B/VaDYnqc0vOx
5CjC88oVzEn6BKjHriu8zq9Gr4OFilvAT3wwAcFLnB1IZlNx4umr2H5dbILAbe8eKRSzLBazfnVm
kKOUcOiD4KCsVOLbTo7/W5xZC1aBHzOxooQVTVWU9v8Svp9uv9vlPI92l51Vz4VVyoGiY+AhhheW
lWwQWyw/xlhUygXMqJssPkZORtb6uPN2d2+gE2sh8W/58tCW45BrWu/TiFlmS5LrnzDtMOXltYJI
No76QHRIxim9VAr5lm02N0xxnAltvnYPtbuGmE/baIxcaF3HEYyUpuCtPbAeDChZT25l3WIBalMm
FEGTuyVmn/3Op5Lks3leegqa9wtb0J2SE5L2FVXbA6hirBj2DEve2GAQTZ6ORneLqg8epOWap/Ea
fWas5U5N+Y2MoayYpe2V1lrSaqN4SlZ8MTuZRMrvj794m8pS+0LqI63uYPQmxcolL1I8hNg/kNnI
rAGSqW5czXZJA0aw/MAVoKjmDPHpdDNGNfeSbgo9O/cI4oqj68Sy5TMK9u87cZ9mub/7tgzW7ASZ
xUwr97kCvkcclZdJh2jTFGXL8teHCyzEUijII+WwsvTLPqyoBxVgYci+ID7J/8nKM6h91KNmB/NN
+zNCv25Fzd9HiJsZRWNWA7h5uslFAyjBfTLBDLHsU3j2IGbMV6APJDR7r6stINENfo37HX9zSvwA
sBY+yDZ511Esxp5iDmNV5y3v0gbA5c37bLi3eQ8EY3YxUV+v2gIRUBj0fiA8T0+NoY25WfmWqXd+
u7yyU+IsXcBxxtOQ7sihJo7MVkTXZRujCFdpAuYTxrelT374eV4LBtHlPNbDFo2RKpPfQVu6Do4J
uNLmZpE51j5L36ICAZ6ZV4AauJbWY0bYwYqpuCbHP4aF5oMAotMw4gWXTK7OGRwjNyZrgrZE+lZ9
JGWmn5f++gjTYHcVOT3d8NggtZJ9UZSP61py3CV5uA0W82nMcd1UFgo+b8cqHXrY/pOGqXMFdPqD
GDw/Bs4XmSkWS6ZPrILqGwW6O/AIRqjmSKkxRELE5DFnTXmD2QuTbQCRl53b1Ok5YdQwH/mzUcnC
sEs5JulPfZ5c3dNVSPM+5K+BUoBX2eBARJqlDiyEeL1tarXsj91TxdEkwvPiMYNAWrW46hpKijGS
9HIfc9odiPU2VEn751JYOduW7NSBI5LhLtnUdPdIffwc12+6N5rxrxEFFroSzr2eBV/7NboR81bv
vn9Bx2vchniB0AgJUsgJTD7Oq0Bca6SopTtsq/UmfMFhXy6fTx/VmBUSerKdwkLW4t+HmuJxfc0H
ibZOwTp5d7xL0BY4xgDMoiw1HYdleQ0gZOQaxrhTcyNQWpnq5wPgdJVYbVojwysrcfKwZtyzyRAJ
3noOByTXfEAY8atmCyvCnMtnfnjvaLvPolOeRLMXRdwDCirDrQXPNOOjk3p5OclQ9o0UyR/ca+cs
hDDjnFrPK1BlZOEqSuf6hqyQiujGQtnpW47JjqwGAYsAO2EznkZflPnL3WAu1tAOI1fLPuU1bbHs
yyxVKOahP9cgHLz26ShOJGVFZMH1TD2BrtjOtEzDjZhqOzotZWKgBoikNsV8KVTEKb74AN13I0sK
tYRvudj7c864bWvkJ7M0hS+SZ/wOE9vk0YcGrMSRC6ku+A7phvC/R3g1t2SKWUnFpZuI1BC0vAFl
rIbCufNMwcwgcDIQN3T5XwR3uFzsOUgy31YEWMv+jONKa6H4i+S1jXmu+yy0jigZ7/INYfCi7ano
EdTbzBxzcA03tVS2gOO2bCC8XAzAwpAcpXtGxrbq0zd5NzHHNsuLit1hEJVyRA1j0Mpcv/EVlRKS
pzTVWkiP3hsduwhZAYiEYDQ1XVY6cjdTmRqnIQrVV+elh1MA09I5HmkYgKImVQujgw6H/SpgTRv/
qW3iRR85vkUOjR0zqs7kBVQW4eTFJn65wU6lWiSVagStVQ3IuVxU8iTSVAjB5uX+r2xTdeJynrXM
MsDs7EAZkoBvVWCludLsBtNU3jr+69/l2waMuwkO6z5+zdf09Hh9OoODjTQG8W/e4uqH04YFovrp
+1BLhIriE853wI/pFV3+bM40smXX7Smx2waoc9H58gHljf16Q0nu55fLMwULkcSx42nQNm6xsBWU
o64NSX1UP2tCNqeS5I4UbIol1o2fx+WU+HiVaUVzE78EnMUn4Fn0B9NoDgzL0S/b//YO3cC2L7NJ
3PF8nwzxZ8k8QPAzsb13LQnt/mMgPoX2b3zZVbQcLb82N5SWZVw0Rf9PFXkUe70uo4MSOnEoJOqn
v1rcDGQXWEksCIEgl3vL+SzWyWeqihllQrPRxcluD+AiicWK1A8EsRFBflcNCGjILvq74RUtRbdG
k3cWUpKBFzZ0MaYwDSKPihBDaYrkp8P0rcZphpjGd8LiYwZGtfeExgRU1KFZsxN+Y3XhE8T/agGh
/x3fQmjiTFInedXIFNZYDMLyaVVDZQjGd6J0S2M3oO4zGIU967xmce9IhmhGhRoFSS4WOAlBoEy+
se/yWA1BStgxmxpKUgqLp2HopoZqhRnOsOVEvu5pVMuiMzi7dG0lMPfMdgaBJulOU7ryxyOOYjSA
w3s0wzy74ggt1CzzOqO/dFTt/cwSCFPWayNanKwRFRYlhTJQwFf5rXkx27EuRROOjRwD8HiNYFdz
1hQDI8n90zpxVGTP+sGc3u5PW/wKLBazjNY0ah5epgnnpSbXhexksB9mvM6+dsT3p3hRudJiepFJ
jXgdlGhNJVlRpMeXbWzMiJfedXj9qgEndyuRIO5DrMmRrDO6KWyHNuqKskwN7N38U/VoYFfQ94JK
3WVNHQtY9kxJGmflqnTVN9RR8fCdpLJm9s5F2MZ2LOzdcP042CssEU3LIKCWwmNNaaeTAY1zptx1
VvUxk9hO0qKfjh+t0VlZpYTuzC/kQ0PKAEEqslmkQi8FWQJajasA07Kn7f1Snou8kSyeM4Kq8ei9
fO4NCwnKrTjMJtNbnQY8N6wUcw5uSv5Hk+XgkavXDAWt7lADlQW5VPk8eopcym6sfVbYKqEAz3xi
XNfJEgrmBOX8rQMe7F0IWInp0SJjjmgs76teBhBoAWg+KlzYfl4Fp/K1pOlnzkuNceJEPoTeimB+
6XbGj+Sil14CJ9nFEujlCZWLhi5Y8AHU7g0Ag0mv+wCls/qvyTCgWbDVvVwpB3zkKl7m0cMyYDDA
E3ZsBGbpmSeWlYRQXOhRNzn8IvDUUvoErEE97auBRMmObw/lcYpD/WV3Dz/abNQMam3ss69G8fpH
T0PPoiLIF0kw0BXT+U5ophb6xqu7C6aC4eTdACsgk/X3dRs+hnOp4tWFreYXUY/O/i/XzVLAq5Y1
XjvBEFPSt37MBxLf2H9UwX6EO3m6Rap0vvV7MCCy/LaM/VdYt6XG4Xme5yT+xJZ5229k2ts2Ezx7
88rD4agxmf0H60hfkIfYhmIbJrSLXcnwtsNrGqCUgzCGkEGXZYdty4jD+BHAwz29dR7W9SmYs5Tu
vAKW4aA2u0XaxBAQCtq8UiuGN6QN5kRhFno1EbKM8dP2wU7+HpLGQ4u5BAJdKh26mZt+Z+HjBkG5
PuMUFgqen8uwNNe5hc5VtQck4CvQj/eIAlkTg2qZP+aF1iMO+r8XmYpNru7UzlgeAclCQNt+AiTq
C43n4H9ljLZ6caSLQLzV9OxmLQKbB1DEloC685T4q6heldOdJ/6wNz91FjLfkDAXG1ugt1xTFyPA
P/kkkAYdoy+VXEsZRD/GLCFM8oMC5+JgnWD0UtYsE3BHxcjg4OHIPNDIoB4fNkwh5TvEo4HjeSIR
sgK9TuroqEijae8uIYgJjHBlFodXQQiRIOUa0i7H9jTJsPhipN5LTGq4StX51Ff9l6YKOQU7TCuG
4I6v0D+8k+Ud3A1MZqPO8d4DIjG5z3rntam83ZkExlIzjDfFBu+Jws8QTAcim/vzwk7wltFwdX1i
AlOX6QZulLdAjpwLpsQ9s5Ioe91tmrya4EuKHki8WCvB56HIqFnZTnUD7nHhW0ive6hRAyL5XMa9
WBXoSkhIXyoAg+ywqh7EXNVBQVob2HaAHqlAvpUMTBiz4HKXjhWEWzC85LKfuucT9x1yxT9x7onZ
veiRHmN0VM9Tc46z5b1mWjOp3r88mTCDTg4o1jHRLxsTyPAoVUuGP8sJaLr1k8i+Hw4QGd6uRUHS
gWJEy9q1Ji4QAdMKtlR4A/YJ1YWNfqwbP43NLjPD3OZpIXny5TqPYH4JDNQJkEQFfYRxfh8+eH7G
iTcJLc049rWHQT+2cMLQcwetX7/oWwwHDjn/dpxzO0yfhZ45k8+te3qxlURADMPVhavV9lCnUlPB
h9s6N/aPNVTLi9Xwn0ujZ4nzMEkSfKu4NFHcGMT65IcafqL6Vmv8iaNgxPVjZF7UJaOGP/K1A2So
lfBNGXyOjHlxVB3c/oWsKyWY18FJ9waVBcTs9X0agF4DnExNW9L7s9F74DtzxcBKzSdFL5qS/YlX
xNDNRnlr+NM1yTIg1NQB1pZUBFBRKwa8X8A5JswmMoGYVGvDCVpaVebqdYFNBWN/c+BnqSlI+T1d
RwgqMPT4IFsVdAqTK2ZDSp/4kLj7boy2fMEi13/vqXPt6CxglaV7H4BOnGIISq+61J0lPqteYQBK
PsBiHi41hANGbausObTpshytiVbdXMky96IKVxOTObwuyxnjusDz9R0IC/6chaQgZEbe/GwWPHTt
/SMJQ1DfUvAiqJuHg1I3IBXhYL3INXq95yl881rfVLj1Nhja9jtPn7KA8F4q9YfMg+PnvUI+KYM1
Tpq0DScKjRSpwmxsutYjdaes0Xi+lE0mWTjib+TpxFCNoacBHur0nlt/NnDH19AbJegrGmqZslbf
CPbS4WeVhSA8DgkM5qyNz80KJi1/fF27AMGaW8GLY/2dIttNNLvsW1Ri23x7pYNy8Ez5/GqxQiLc
TunN+D7BKGmH1kVXs49Mm3BkpDuh2LEv0lz8fuDuyWKufgAAC9SS+ILiBFItUGbqVn86DS952Wo2
YGT9SUSI2ph0dxP3ByQ825unxAsjJ4MsURBGQc9prCLbp4Kl240xuz89K1wpodbiw0+lKn3YrHdN
FmlAlm6S5W0B58IlOBieMJ+8SynV/Xo8D8gUQSg33GkJ9zGP1Y9zH4EqT7MjDeU9Hg==
`protect end_protected

