

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IoOiz+BDpEiCAzehQDaKkNxXycZX6DxCheIbVmZVnOeE8xp7Q+9Cdt/GYV8eq/1L+MpdyADA71Q+
diEx2Z9pJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lwiDFOkaG5HcqeigSQ6a9WNJOSnncyPnebjhd+6IKLZk0I0Ny6LWNpdm2fV6AG4pFcvx58T5yWEl
Q+/SeuKD0HNAWdTl0b2fE07zxr+edW2hoGXyef1M8toS5SeJjbmVYB+jYYVGpq6G4uNelAjC+U6H
qvBM4HmLQCceNGUHSWE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UFVaQj8UYHzOV/s9ci9b6/M58BwxIhqPdXQ4yEijf72oAEn9ivW6AsDsNzmhpHIiBklSohpBNUDU
0Mva3SAcsX3+9Czy1ShJ5GBV/GrTCNonRWGYRXu6d9ADAsYZRaJCV+2s1kEifAqI6MJhteonJeVq
EumiTmv57LCQxMW5bGdt9ducpN0oI1Oavkx+FYROiHKMHPR5ux/CzqaZUlRJQvJOcmbQcmUZt3v1
KBK5x+Z9B/aBdtf5Z1OOegRTMkPGAdkXGlAX/Ax9OEiQYDv905iua1b8cAJu7PD39JX00W/YP189
CxrWyFNefwoc+rk+siGiD7Jjf0ooGeZDZmjyjg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HK3O5vzCNER9g8js4SKz6W+Zie9dlDlDlxGQF2WrvDyya1unL5bBpCJy1w0Xm1cUo/y5lNUI/ADI
uYqE7JGFvbSauhLZj4HImoydapRAa/ZLL9nSRfszIVrPI8v6qGNzlAIC3uzmQS48iAygYUrq9YT1
qPItKzIRjW+YafjsvhM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
haBqrpdC8sHCosML+5AEE8iaTVrDueP49m0Xd+C16lJUg1YPcQ6EHNHA456bk66+nGBPSp3B+PjS
04UE5wn9q/J8cGL4YbVE/GY5wVAtR6WtFplMeOXISx0KcrI3qk/KzRrP9Ji6/ivM1RBF/A3FJtrF
qq4E0RTyXYa205RDSyJAQ9RjkwZRwEtkcJ6VY2sYCysbDHMzh/lD130AUg9VBNSdV8LSRVpcwCzZ
sRog7YjwhxC0jQK02UyUpzfW4/xJ7RqEZDh6icr8dQvRuVfwm4y9IzcnYLipDLpn1iVw+wPGS0v6
ZJj/N7hNXBnHUH6mTiT5qnqc1qaRllFBLOzRgA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8144)
`protect data_block
8MtqhLQ3a8O7VxRSFdl6PPeWy0ica/WNd80GSP40HOjUtjbRhTXeJeySZlabSiwc/0WPSO1va41j
kPpFBZYCbwEhr23JVC1lnqfmf1VZhSbLraxnpPvUSx5FL/xv1OOTOFUKjBBJUd85F6e72zAyIKIK
Z12HVP7sBe8UI3i+GsAQjTwTPkr84gx1EjyXrJ5e3uSeHx5j5gNOPKCIrKXRfh5J53Ibi0ASFlnO
8mnN4m3pDxBIFx06zBldY1Lk2fWd7ZJfMrrWCW4QNaQN9L/z7o65kxgD+dFTfdwgTlHxkQlNCWb4
JLuVSdYERrd8JU2LSiHY+qOQnchXKemzlM29BjV0dXuWmBMl7cgM3zf0xQ7GrwGIUruftB/qjF+k
n/HAiW29i+uLTxcueUz5i2N5g7156o9jiL8fJ8b2pDIIIjnHIpUPKdb9sVQ4Zto0lQAAjCUoQUW4
mcdiRFmnD9kUoijN50mRp8f9CXT10cUBLPUqsRGjXnS745/Wf4WRJZn2NUs6tGHAiZdQZxBx8mXI
NBt7ATJ7vV1GPHpRLG36ATVJ0vpGF9ylr47z6w1seglERuiJx8H8FQEYnAoduSvwuv1lIRXuQrwl
FeF9/DT5IH0laf2CIArXBqrUvh1XmF8mMg7uHF4zv6023viSfpd1quP7d2kP8CkcYgiOffH/PTGb
vHShQO8B4bABcAIZaWaq7Xkx67LkftwQIIAVR46xoARUi3bakTJnvrG1h7+J76IZRBbQvWZlr5cU
eTY31RqA4r0PMWASTGvpXJGiouL+V5eHkhyxg6T7CFIZhld5fK+jnfTVWUv2hZgJhex95ISLVW/n
mGS7YJ+5KF0sz/WtY3tE+G6tVyHfZZ2mPOlDSDlIJl0Sps6R1jM6nXAQOpSuJ9Tt8spoC0xvTJVb
c8iEUEts4gynEX5AOMc64W8BIHsna1Z5N3BPIMlJktwwye/Vvo3vjz41NY+SZK5HeQ0s/QGnHRGg
hlRw3NpSHBfYVb3mewd2UZ3UJC0xXk1G1oV4ZS0ud+pG7zHcRge4kRrEJT3azurzV9E66gCzm53B
/4sGfye6/dKOskOQfbG2dkXA1B8Otf/L9K+DEsRoBKehl856tHbmOJoH9rqMW1JFpq3ld/TPSLqX
R8SXnyc8NpPpST290PXi4xGNfLcu2S9tgc6wUdWz7IDxbs9o1azPfYP58IBKFJHA/o9tpwYtUvSh
JkyW8/7UlRJEQYUlvPj1F1Rd05/cMc1hi4Xjw6qwp0D36TJYMksObkEVXFwNSAOCD83oA0Njv2t1
nulKBLKPgIKUl3EuvYZa3hsug4O8kjcqcOs9vRSjvczMDmKO8ejlJRW7I3yoS6L6alGPDxKxxb6D
K8aVxKl3AcTHTXMbVqkZMqJufD2Eg5ZyUAv7bg1y3Pn23HymAnEjScwbvGYRiRB7svwDtcr2UDR9
+TlAB1bPb7rkLOeI1Pcd1RciRIUSC87uF/qfiDJs9HUaBxtJF7Oy39fI/M9ij8vNDltSVU2yQDdF
Ak/kHPtmoK3QRKy7xrjRHxXWlmelwawTrTJALdwczqeJiXMqdl1zpmCDFezOAx4tzlVrsBw13Eh4
ynADGG73r9YM+kMi0n4JIQB07ASJ0CKkcANj3jW1ojmoSuBMVjeFzslj2GwIEtnt8qPJ+lzovfXN
OH2wFyqczRBILb+vSRDBocieGQ5r2Ehi8bcKS9y7hmc7ul1FX6FP2XTHcXAeI+IIEF1Bb2wZCVdA
qwVa9JfK5yW85FMC53KgxW4k6XMpiW2Noj0Az1/e1yg+GQlYl2n3MvDzBj4r9+9ustj0Zzjkpjx0
iwHb7Y4PFLaUUxUGij7vVodP+ce7o8pxQiB3SSW0rVqHg37Vi786vSOoOdKO/dzodDO2duhjY38j
9un1oQuACYEXxyqsee4uMuKYp25/jlsxmSXbUzLNcqtbLtUvBOwwR4SdkKLxLtBMvVfMMhawukwv
B0tWrt55AntgGtMK30PQ4QLLMxfrJp8BWNth1kbL/uQOATke5YQoZ4fDUdqw+FsHJ7TM0fpNSjq4
n+NHyK7m1zYXpEUGcF/DnsNyKGqa7lxb9+DcdkvlHwmFP51pWFcFbtDdD52RLVMT4gfxXtxTT2Fi
7DlPO1884yjA4cWwhkWoq3m7VwV0HLrzQLRa+MUcl3LrzYu6oxWQksorpiaUV6BOshRBwsiktAEr
/wK9iVDpY+cSm+HcLO78TeBGli7whF1W1ftX7Kt/4BThKsFYDczfcbGgMSzOiQLjRr1IG94VEsyD
49bwGl709Pdyutgoixgxv5s0wNxR5ASkwr6evgBQOoogr65wac4s+lMP3NTOBZswWbMlOROA4KV7
ymZEpqGkzaGm5b40pCwXpbtS1utlRz9JqBwGvo7XU00N59dMp3oQxHNNhzwMnZPGIVDdU4/c2uts
XgHUyS5dOrgvQVTAMKKxoVMACsXSpy+/o516xzt3+qoUrhML1gIADKvjBbcububnKTFwVk2ZKcwQ
1NFaFawIN4ksl0JQpFAX9vRMiV0C2ts3AJzOU5ObBFAhYkmrgcAGwE7sY/VRfL7vu5Au0Ok43Vsw
5ic7XtVt9bKQKFOya7swj690d+hDmkyY+rwOw/MHmHJ+Ip/swKOIGDHYWAWWL6IAEFo6SJ/t/L20
NDLw+cPx8sh2xOojawekmQopPYCIY13XvE6mEd33LfKkpD1zPEuJQIipEcrKJSk9cK+R7FEQemQY
zBn7T8bDAHG8NBwqI9FyLrdjGXSsa4HtCmCljbKR7G/2a/Z77i2Nzpn0Z1iOQ37Cddc2avijBrz1
lTxn1yUsTqFyDToRZbPlj3tkOjHZHgzkrsUqXmDjimazT9bcjZQYxaSukAOWPCC37XqMPc/M6Uqq
2NLTdQIoWArF3nhALPvALeDXWy3RBS18W3wyqgHwuED6TumF9IUUy8Z81xi0Aw45kxBSGQAEjVix
XcybHhA8FlTjriowdUOGmnOk4dP361NuQyiQWp45W9OMDKIyeZhIdREmHm7mlhrFoDHXvWtV1AaB
RAvYsHOcBAzzO0iolfxxhLZtSmMfOkE2YLrVszIbupG6B+SCaxWlE18cYFXAzZJsUEPAArvujL91
IQwcS2BaCbuKFmxYlQhSduJoX+RyMErDApFIg/7PdAs/Gm0iabmUZwRvTdWzE35IHRm8Jq0PC2D5
JX4Ll87jjwiuEBkYpI918PFaszaE2kuZetdD6REXkMitBBAAMcbnOLF8S2qiERYkqTcYhzYwY27l
kgAAmpadGX6W4MAkxNOzqbMjUMmCOPrAWuOVhvKWNL1IrqQOLp375CAKLLO/6t4qu9o1y3xZkafV
1XC3+noUsdSkXZBnVaJKibH2a+Aai1sBJujfwlDUwGs1w7ioliGlpa0x6ON3A03ZRJq5eGHmAvCC
15cxC1oGpBeV5pHtMgwIpisNpraN7Spzg5Mkkid68819LpgXOcbYaGUPwfo+UV8lqLhGioswL6YT
PgqQmN9x89kAneDLpACGIj0JGBlfegnEM6DhKuGwEXN+T9KdPZjuNwlnYTZW51xT9lruJhHEkAYs
JWKchLcc3DtLUlCt8NzRyvWeXWv2is/pxqV2gEtuw7Xq6w4JmzIfHoJ/yTFbox5FOU+uOPP74spF
P6WwvF7F8IcAHMoHzN0PmHLybDHtnXPfMMuumbwR3sChM034b6VGk/lGIA97aAE4Skg6GkShkJhG
7zHY49clsZIBskR4AAOAt1SMz5yJV9l//Os7qsmdaBBA4siD2x3GVERDYdWmLAHfvB2Y5gCv3JKm
9G/D1VArje8lXEs3UtShaOVmjVP8z3rNPA7nPgyGPx99Ez7wveXz7JFVSpHUF/1QXYdK+vX9zpau
z0IaU7dmrobzTZUJ4hAvL81QEULaXDOBig0RPWPGt/XgrAsWW7V49iCH0+VNRHNjcQ9AIpGaIfpt
pMt2QRVtJG+SdoIGQhfn7/NqjUCfaiCjw8oCJZt3WiTMBa0jm9+sDcizwQYgEonPNXPPRS45XTx8
eUQI4g/vTnZxPKFFBUifOzNNHMqMJDSxIAWsSoy5EB2J1j6zc+7DN3Wik8kwPaMXgmstCpwLXiYL
OPApwo9WZnn8zbJCR3WR/NTKWDlvQHbt+x1pAwE+fHnJMcjkJhP403TSEAWugMZPEmB0mGU95hxg
LXmmVSuoFbsKlzHHy3Qd5PvyY5tesm530czw9so3hcvBB1Fy6RTe6Gw5bXURiDOsWJ7dSDib/SAV
/+JCBA5pVav8oKpugO7IzjhwNsCv3QjcXtROXzMODpOT+gja1vjHCKcgUyPznsQ6FvQVmgYlnTRN
m4COaHBN+A5VWiCB+nDg6D4Rh1QfZXTQLNLCvAIhtfPeChs9bxiMZAJ8+wqIFVLyHdDe53wS2jcg
/jqDjBSpwQM+TaF7NogLTg2Bb3mP4+D4zOAOxOkDfEnPsSnzMaSJvA7LEbDKqn5KX3aAY3D1FNsq
4YW7yrKw//1pzR4U1MvvYpXsfsRQ3Bvx6ZEpASAolPy5aXW72Tx0LZARvmcT9t03dSoMvuXmDC8E
OZtKf2cN1XusW4/IfB8t63Fbaf3MAbYfX45ImesuQUga0RPlM4RRqh/O7xrTW+9YdETo+foBnGO3
JzezpvzDzf+/7goaZaN6P74fDACsJQj6NP67R5JE39ZH0clM8SZTRsyLlJQk9pMROtbEEnSbluH5
mez+Md3NgH3VJgAVXNSkZzjN6NZ6xiWNh5Eifqw5ezfd9v7Leegisc7SW4G5nchTBDzNVZFQoQMe
2W23uIaPImR/JP1dcUcIa1vNVN/E/7VhLCWXdYDdd43ekgKGI9v3cTcfClOUVjzPtcy3tXOwP4/y
7rV0f12FDeeaiXXIzdyWE6a72QaQn7nqC/NW/1Vg1lEOmS9xJIbaEx7Z4v0h6hkRahNofuTynWs2
NPpqiZclmdUVrzYTTzJ+6U40u+C4MIIN0fsCOFPIUBZm9oe0pZOmVeA1QjRNypZrdAsp8qGSM/dB
TqDkgcYwM7FEN1E21HdJqSW1qvBccYVJ+FuRCWkNgXLGapKarDfgmQzTP/NiHeZpKk36rweAm6Ka
8Zoj1y28kwu0eJgdmtDHzqjJL5u4nf44GpcIdpcrD1IbxrbfMOMgwHac6sPen4RSgnax+xPrMoKX
aRsUDMXYQPzx81bbix3cK+76YyaBVpEaytM5zk0fzGC+4LtqzSvTQ0YLXMea2jpDl8z8jeo2EYwj
xZ6B6FJzlespbEagADzDh5wMdqEWb4qHBTvu5UFf1LX1PmEmK45Ipn2M7vBrNxoMKL29AykNnxIv
JOWrBP5BhdLAsVW0t9qDugDwv3P3oQ664YLyZTwy5EEcSbJo0HrNY1tRkKz1snVZdPBj8Vsg5Ulx
5L8ZskHDnZGYCnaHY63LN8aD24BflBPfeIywHfoZSlB5VzKLgSb2r8U+/PcvKxMKeo5wtEArF0IZ
mB4SouXl/jqKiuu+HeQB2LEwT+XBafBQdcYXgqEEOz+oBpBhPWddIbXD1/ZrFR1Uc4JzYKSbSb9+
9K/zEBeomXkFXcbXsv3S+I/oniGtg0rYiFp+6vl/k6EQtqaYTrYXveImPyGthif+ff1vwAKcs5ez
4dAdBpOSkkt5ymlfMVrwILmDwJ2O4V7HI3mnBNtbjTVoyEG7+b+zSLxFQpSYIU3b5O8hMV1sih9d
Jj6T0tCPqXQqcXon0JxHDL01jktkNo8iU8+jlW/0/9tLljPb3rU8jkntzlGXAiOdZx/cpFGwAyYi
NPn1ArcmHxiokaMkQI8bhTTKOqwsje75q7t9zka1APa1yxgp/iKmfzuhSyHavDo3cdIAfBtonEZ/
sIfLMgAoamlbVm61IAE1otabMhpD/HEYSNzvQA5EehOTPNCG7FMC4GxqsbqygKrnr1LtJoJMO7E9
VOzHPOnEp3PohtmBSnawEK4MajP4TsqV7DpvgHDz90EpoL+TveijLyp7+Zat/uz5OuN4vsroQpBD
cdUUEV/DDTing/B84W/0om0RsJbXPWAMHB83WQ5NzGlJnCj1kv4mJr4aBoeeidBGhtAjsrOE39/l
sQzTbENVLZ5jcy+IRO/CD02Zxig4PeGsec+6GuVVEgC9xTdbMTMkYrJZhuA+XsoKH0PRl0dMh9bZ
Z0jCXo5nnNlQz9DuYYNASPu5koTbrgqL+F7x8X8cC0yUvbHCt8WR3elXPSrofwXsuXRWXEJE0r5i
AnAgIHgzAaJBk8bd7useE9whuNlT+Ji8r76TpsG86UufLqNjGfKI3gDUlfhTKx47YZpGp/1JcuzC
ofJtH8unnUUwhYfAfjsEqaDFK0uZVGF7kwUOap+rC428mmWRF6U4m8y+OSC9u6FPx5jIvS7jvPUs
kmFYAq9b4zVNwA3882FMJxTmwWYW5EJNIa3NRC68myKPp0j985Sf14TcnjjjpOrUnO+GRiWhM5y0
yDphOaT1X/3b/xXJSKadNuuK7g5q2MVtZkqYOQBZCRgRFVzEdpbdVtDFE4ZBGIYVbjtb58D5BzmR
Dz++SLbvuZ4102RDg6N6AE+EUYEfeAQ536X46PgOXlXlwWT3N22e2J++Qkt3gFdZKR24lrDyDdtK
269KTzMjJx4//pd8tgpLRjE5/9SLLHkTFv6Inan/H14PO2tOZIjW4VyOnou9mJ/6iWU7tFhJAHEW
wkB9Z9UhmOgaZw4SSJFLgfSgqHZdsnpdIGefx9E+BSK8tklAKbnDT5qlRDe5Nagqr/fSgOX2HL5i
p/5H7Af6pkDoM6GJzbU2D9F1nTFgnK68ipv7iMWD/yULv6dN9vtXzp9+pKuXKHXUb2NT0XFVfjjQ
ILlAwTt7fDYFBC8yzcsuHnVzbnqKIs2/B4lgmPGyLfilMl2kaMuWjTQxm0ZPa1+tBNxn8azs5Vcs
oDsiKz9OaUNsuvVpGC3X2QYInAorDF5h5WNapdd+ygocaDXyABv1WTQ4xMMgqymj9gzWMW60ViHF
Nw4sJucQzkZ7LNCzxNVAZFmupcFBAgLJzmBzyHMknKxjL1HSgs49zhW1y0ZE0yqZS68i2MeyaffE
5tQ+FWyNOB7L5mTbLL5+ZLY/3o/J31PLRJJfBLVczMccV22fo67ea3kXk4t3PCDIJ3OM+3Agb6/0
SqAK7venD1YmVOxKfOT2xr/35OirD/FmZgsMaZHuXi1EpAaMfkQRy+Xnc19fBWjKDVn5qeTKci2b
4/8YSur92959e3vRIkzjQ782/kvjagZV9xOZoT50LbNw43IPWHeFVPuwxzimmfkOrPuDCcawo/l4
Jy3LOmCtdMBuTbSG9xgb1IrmpgWUevqnRRkZq06RGeS477W9vYBHi3V3ukeOyq3d79iv92yNVCUY
Fhp10464jDyrOjs5rBOZtphm7/HefBHcRzhe8EcGBoBySh2//eX0wBKUZW/mkI4oSr2px1DlRvbA
fahUh8K5BbhdBY10qgRfVZnJ5UOa63nyhRkJm37tuVzaM5nN4OqLYtaNbQPzuvZsze7pTj0XnNgK
hd0r+jbEW2017uHrqpbPrVS8kME/FXevmo2wB4UuHfbUHrmhMhcUk1MS5ah3IdSu+e0vdRXhONWx
zZeKdnBJMZRaT3KbHVqyjk83ym8fDtBrkY3i9T/hu25jMPJT64fs8B4z3fycU4QoCl1+s/W255Cj
A8+JUzHuJSYbtfS0xhNrIDguAzQTh03U0JFsQNlBzj32t7v3AnL5yO9QHfiT2x5rOqdzC0/heRA1
OZaOqbh9DrI5msKmBFhwrlWq7SAdJEn3HOGe5AJcyBDVinObSmBP33uIeM32q/Thbf+8GB1gh0BI
72rMTTEEuDiiDqNt2kp6htABo8DIRjddivEIo/Eeij5jPCfjy1tcPlHKNXY7vtTCzDVtjHATLyO5
SuUHgqywxTgOfIV6cjSFeGLlNV/aky9e6jXWtNeMSwve+Z1xpnHc/TCCNDPCYALYKIFoVj3Zq47G
K1zhw+xWV4cAB1nlnwREaJvwLgslqGA9cjgQrCI8cuKJTLXquxJXuhIgCM07YqBDvcMlr+MDX/mF
+k1aJcLXVTdPjOuvObsN0vv1JOKEcucsLqYMBxC0uHyULeU1RkX774IWh+VNdkMOSbXpOjL6FAS5
DHOftohDd/l/glfWkENp42a5cVJoMMY/XCkOljEc5mSCmSZw2fp5iEdY1abaUM8tTT5qx+8TiF6u
dshvwwNipUl4y+bq9v2ti7nqFQu/TVoHhuj6uHzcqskn+K8wqlANoilqMiegWMOVFMgBdqPnTZ/f
PfHuQepPPZ4UpPCR+20wYyidGEckPcN5VGeHsmiNPgugXmYvnq3QPSoKvir3VVZdezGoMyFuaoBa
4mpSczmXzwRB5C95lcoQ/8SwKMTB6pmphHzGd5BXYnLvhC/MAhNxZtwYoUmcvxQ5OFYLOXHyrKs/
6Fy1/GUoFQCsSi989/noASrbfKIvA4vBoX9baCH8Mu4JKZA5ZY80i+tt0rlqfF1dcpMRkca+Kf9p
2Z5p2UV7bTZ8BJdp7uiDGqDHrq4xh3j+QJdxWi9CL4mNEtLl954W5btREM/7J03xZLZSWv6TfbLX
P13DqnXWoUsVnufxmLKTNUorY5EDX1FDdD2sTKFtXWmA4bEd+L9Ijrgj0xhKo8smSveYZT387O0H
G1TvS1TnNrNmkSWGgKq927Ed2ILd//SbO8uEr/+VXfmG9sOS/lCUsjIkm0ZROW2HvGlCEG8M3zNW
oNdYPTIhZGL+0CO9RcjrokLacJjbpwPWpdO6Naoya8ye11HpRWAjx4Ndre7X3b0F5YSCZ9Kx+9rf
bxz76VotcTIuk324aexEc5d9xLtpMv6VoBNjWFpPdbEHW+Oao3eh9s26ijgQGFlAcMmPxOt/4CJH
gYaSLv+OEyecnoH/JlPT9j/zbf0nlCZpb1yAP/in0pGLNa0SQ4OqKiSu81LW5DzXTaB0MIl+YO3q
JKLwbb94s3k9TPHrDjiDHB6QlHU8woxDg3xOcVwiVrrbkKpT19S7JI5LO7r3BGHaNTFyyMtzLsUZ
+zBAoREd/CffKccR2GHcmdIgZXISz9oIPz/7k7ccxsFjaZAe7WGvYJ6g48l/qK0a7PAjpkRsmqYf
cQ3SyBIz04Y2HChXFTU1UPyBj9GtLqGM4ucYxN9ib99kBGMPBK72IrMnYAxoz0WteE9jgDLveS5M
U6lW09h5vD8LfmyMnJ/10NJfc42Ye03i5vCaaihPnVGjO+7aCoSWCOEVFoCDJptQQlVVYdZa5dT0
dNIxnQ2B/Zf43w5KX12/3X3YChn/4cIDUbNcmCCDvxoZ7xqvbXoo28a3fa6VbqI2XkwJs5zr0/gS
EaAQsX3+n4q9Q0aGB/5fDRX/tzGZDiCedveYI4wx9tI65XrBk/BoENUCZwJCtSsmWoEPWH/qtMAG
03T65j9+ej2leCniLpGPfQOefaJ5du+jue/CmXWMT4ppBjKrVWhGxpcEQ1vGy5MKc6X4T0pkmATo
CJJhQ0wJ8aC2givr7Q97+JzOk8ybYwnj0KziKjpN0333WOEl11h0tFOJhWYzXMCpFoJnfdlzpSjj
RsDrP9tRZpVIpJnekst4QdgbQ9coCUt2C+nYKRiiEEaGQyKpUB2MkvOwJz4ZIDfFM9Mz9YuRotzt
fr/ikf4XOjV064fjF+pRgMyfmXN3FtHlep49gL2bqiysJy6BZ6xogbyN1yGrLyJhIO7UclEUgw40
iM7KNXOlUw1o5cZgnyh9nimxnXhGJ4UkpaV0rBaOZHNmRvIOE+N3LunkM1sXG5vwwRJ6YzwKRCAL
AX0HgVjQyd2ohXxYoyX8dXLECzdhwCjUctYrI4BuvgNDYKxNcue7/+4rIWzgP4YalkhugSux0cW5
9FftFz86GQW0b2KMGGJN99sidNmRat3EyCV/337tFne/JHGPXKUMCiwF7eMprfmcH6JO9WCy9DRq
tim1WYcnWjNJhMonLvMGg+qMEsc/aoJttEQNhXGo/Pvn7CDD6yOpqgWDDE3pzZ9kQB4zY/AwSlJ0
bdMUkGkrICE1wQpmOW9aqQ0/HBpzBb6S/GgF4/zhafJ4KkoRjvYGpFeDsn9x9MFOexqikZh+fzyH
0dz/PXSD8GSaDBVBwT2619ixVqPXZiHoAoYf9EKIH1fM+UoELFNrRCparh9WH20uOy6B0S+JxmY7
lVgsy0xb2UaUAXVYOPDf3ymczO7ONyIOWVhM8RbgjMeGE9qXVYtcGZ26CKXYY6KL3CIPL10urgcO
1BtfXMFyyJPBEG3Se0hKsXZFOvbLMUEhte1T722V+yO0LYA5hdCCk9EiF7WKo7CJ59qZUdUm1KOK
hONjz7NLPxQN2QG/2pPQlgwjl/9e0mBQN+P4ncWlWcFNjkOMJtxZf+gIbAd6gKGT42O79p6g0Btw
cU+OWc9Wqhuzf/Ie5qXDFE87mdRUrsJsMXA2CE0ZxQonzwGyD5Z4sGfL/Iln+YkdjYDIwgq49QXo
snLlW8xCoOJiJoLIKPA+WV6lGuTu+5s/zi83liQ90p2PeDGAu0gE0tg2qqwAq4922ZXCAUcrp/2u
fIIMGG7HgpjRa8064HWWNKyJttvgHewe5QiiFO9i4YjmUnWcaZsvCiuKiic83tGxjwl2NstN7/7l
hPuERPXJYuNqe1xzXEi9RJx3Z314R08G2abEYXHDkuY/KBB6NNvLxzjizUfHDJZHTZkEihMH8Glm
CsR61X1iGR0XKCPEXXfLQk/BixPEQoQWWjVcdjYEflAE65WGbdJMFK6N7q46V4YtsjRhBTgZpHj0
f+j77+f7H3moLS8ez4H5qA4RMTuglDbg3YukqpHnJKVOpM7jByrR64BgL7licPAv0jE=
`protect end_protected

