

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
q/LTCQu22IewzFL2xoALv0V8R0cS+n3ZGOXTlz6zO0tHpf0bhYU3nG7YhbNw5H8bMFnHmKPTo6eG
UeGsZXmzfA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RYLOlBm3BPRhwpOnNgJH4Vt0qZdXkt6+qKeUVOFaD4rlCQUegbI8dSeedwyfmRhRBYYfcasAbBQY
SHt4NDprJvJn/h7vAd6X1UjRiIi8OF1s+lR2yqR+Y5n/Ai+CRx+BajVy1wGHxdjiCnM87Cq2Hq6s
UytlPbN46pRkluJe6NI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5Onxh89dWZfdY8AMW/MOzaZUaP+doVdup9B0riUkkwljU4WHOna1/K734H9kkMqSDTQ9ivkZIsmH
DErXjPeoJcAWqHloB9UX56vG6J+JtHhxXpnFa4rDUsDzFadXGZZrXqt/NJt/7/nP2AP1p1qeKRkq
ksYRHunueBYG/B5LuPR00cTpoZaaCYuJroh/pzkerIy/CPNX1RAKt047HCKtvFBXH7wuqo/yaUyk
Xkrxw2AQ0ggYgz1hK0KOdWT2JckcbGgVwPsik+mchcvmPUBKx8qFAnef+ZSGsUTy+3gjDznrQOsF
sJM7rKdsAjU5OLq3k8BWR36ur9hbMdk+lvFEHA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fe81XuZ9RrG7wwwI46b8GZQ5C9RFsRlLr0EzhGvkV3ZMeUUoQPwYfJl6GHoj+GDA9GnY0KeJe84A
xt/fhvb4h1DNhpVnvsOo41gu13r2msE3kvHyK8en6IodL/Mdh8CmalY/a7ZhDb0W+KP7rEAgisED
MHKHkmm4OWbTY9lIJCQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JHuY2RJ1GBIZ6g9aWOE7BqrGN8uQypqLnY0uHGFvCX6msmuceGWWswz4xbJBwz2/gb4ZfVDTzfAB
RXiuZlDm1B8txxWQYaxO0lZYlxtzCU/lUn47fRBxEhyn9Yc5lQx2oW3B/G9c81S8zCONQlmapnrX
y4OR/jDZXLz2wxMs0tkWUSXHisAbuRctLOTsTUfqMDUsJS1g+TDQCDpUDXL43sWg1LCRd7wDn0um
3q29OwHxtysopGOz0DxmTcK07ZEEnSJS89piniLxLQC53j2zOhAk7sCb4iRKccCVkkeasTjlcMTi
rJCab5WZRXi1gu1yWZ5s8tCfrKbGVSZTS8p+pg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57216)
`protect data_block
O6Dkc6LbkrRfkJ1FecKV+cm/54EAyyH12FVG4kU1WsI4cjzMuIfEWK5v9A/JXYQP9mrh3CHW/i4I
asZJkAeeVn9b4CfjfxQ0FK88G7Sioq/Ns0VTn7Srw1IWu/0T6i455sM8MIu+5OrOtOBdHuZ5pOcE
fWiwzySI/6HEqkk/Vx8LtC//iv1EneDEuz+krQ7cm7V5GX3/hyUcXIj42U0evKgTlx0THxFdfijr
KmYjR7GEUHQgEQlXK0u8FkCA7A8mCR/YGkCzIl4JWfRullqCnuQlCwW94aaKleswGpMnetTm5t5M
DM2uqhYlGUArXQsFxOTpbXYFMW+gqW9Uwl9WV6l5/EXMzHfTz3jnN0VGpBbQ6i/u80r2oEz89plm
8N6FvFJRpmDYfq1h4t2zSdb7eg7yYFrNRaf9gBu8+G+Q51zi8uj5eu2TC9W34yXr2TgLP2iLzCU2
4isU0NRR12G4cZFHbQ/zCqC19/PF6ogejahtwGcd4YDHnOUaLD6rAgJa19DgYzNDcLcZdeVSERKG
Sdh5u6n9DkOessOK6dtFuszKLj+QjFWbYPveb8zmZlxd2GT8OhoeNoVfFx5+sKV+Ug8k7mts+lK8
Bkp0/S4k47gtzsmvwWHdj6csnyU271ECc8XY/xoh1S6HUEJBrnEjUr+3/I0fwlHEJmvPzJGzoI2d
tt+EQFfNHJYzBV44E8fAIfxj9RsrWYxC7xN8LfAqixmwaFGZIx+z42bq07y7fzG25cIY4HpOLgvQ
OAZErWEDncWkARooz0COQSRnwUclqLgDGjZn/ybEzfEWvN9D7BGGnrSgEWCcKaV6Kr7CNeY9f9rR
bVPNPfY52MU2kcuLddB23iWy9jWJKxRItlLKtsCpun4mO7hEMxFVVGzoKk2lbucGi0u13fn1RucR
olxqIZeBHveXyY41CooOdhXHXhU+NcaU55yhopnX9XUUjIfiokiZwYH5ZSkx9smmjz5eRjwR9Hmi
f8S+1++1jKr3DGuVPV0Lu3PH9ETqUao1fZmEKiC3hSmCcc/LcvDSSbY0r8gEMJz5oGplLnfFjJQI
pKmwOkyG+UMpOn6E/sOwSlSAzW06bg5HvsTIEbiKimzpc1i7spq1/A8IZgL/iFBgboM5fj9zsRfM
iCA41XjM2VLCGfx9aaUX20MdHuJMtWuZ3KLkHVsjEQK33W9vINeuHd8+M8hHe28kzQL68WIGczpV
FHLIsNPEgigW43cpom8/Tx6d6SeUFm1QX5GQPk+AhPpJCuWyGF5cWCW3F1v3uctvnxoI5sKLy0E7
HNxwhFgsa+jLRcq7QHWq+dBe7qcNGrKsPBqDRHp2FF2LGJVcm9+SrHMeKKlkRZtT8zyhwEDgfrgG
OpFqrONJO65u9DCES7yQGxxKAzlE/XD3GpFzC+nKYOzKrMwpuXTsHD9bwtoCLgc8NUj1BLc0dr5O
4zKyUIWBVFWTffxIp+nmpDxzOVt68qH4j8JQirrNEYx4n6WVjLvz2YG03qIADX1lzdgGWCP88Gq1
8MD5quQWvkIl/QjzmI+m6IrDP5ZX7gyVED7RAbLzFQ7w4wdV8m5h91xJSTiRWnxVDHH44BhBKXSZ
wQF+e8bI73K6l02PRoXS3bCEXX/sy5e8g2j2q3RelPF2EbztdgiQ2D6WwfFekHelBTJ1IE5inifh
3p5cuQ3QL8zLTXZ+rJR2nAFaMHalICS1QYS0o0Ghe8I1XPXU8Nk9wi1ARSAo6dE53VvzfwBKLXYq
hCZ11Kx1Adf/XNUdougR7TehGGh91CJc3oTrxJQR7ZiEM9vyFpgSI4aAGKTdwncc1HKpVbXIeFzR
SXZtpgj7eBVbvnYt4oNnlpWKq6bmxg7EL0uNMjegJ1fjn/8elPVrvXXBlWCfOamLiIV0yv0HzM83
tuQLy4HUaaBMnaXEKjiric54OXTKufgkUnEt3uEoUM7l3vpurfLQg4hYpO8SwbUAAc6oAZaHH2Ev
kCD6GWR582B8/SRncVFw/n84Nw2PvjZBUHTB/uzd4BWQfjZIFOA8n6FEE0SJB/2+92Z8TPrOQYbr
GXFx/96TlnqF+hCaBUXikI9URjjyoGzw3bfEbn0EbxzZCewCSqIS3TrhkUcUzB7giyF890+FXrFj
rY6sgQmoPVHmNCXywR5hJ+/QlMdInAHx8lN//Ga4WRvd6GaNfkQCgOZH5vs77M04nGRf1WaSxXud
+S9wzrWmFRuAa62K+dCUca2S2+Mu0VRiJFcsrg33AWJjD08x5E92GXDeLAoyhk4x0u2WPTcKwO2C
sjye8/fXo06DdO4jjBUoXctnXCpfM6ZAAqPhpQsFqZatgG1cS0FiiKyCGVcsnJsX9hAbS1TciQal
Pd7rxijAX1/hMEhUCWZJmpkXqm9GXaLDOi5/oEcsNOZmbsR9Jv0KTGqOZOdSUhinGRMhCZLSWEj2
7umlWCjFgCcPoaCdIY18EplxuM1sNQDsn3qyFi7311KqLlPUgqr3HkDqZOwTFbMHr2JzlLsacdmY
+SlhKbIHmKTc1vuMZpX9yOBxGpk/pMIKMrcXAY0PkDTrjEhU7zkRQpVNiEMGmy8o9GNhpuUAs6Ob
y9k7dorEM2LiwMQTbWuq7j//dDLlAWU+G+7XwEm0ddRAd/jkBlFnc2wIfcXsna7LNJckN+gjPQn3
Hcz9w8SeOLd/81lYvyGZkWr9cTEligUVkD58EqhMsg3F7DxzfKl4zEVWKZxiUSaVCmfHEEbQseom
2hTa7D0hkTC8fTEI44/KoYmBj6+3XAcYnIAmDQ2pOueSpiAr1H79WX1fiJ+6qPtonoITNJBoeyYL
aYgL/OD42V3HnCerbGruqjxQoAiXhoO12IA0mt44WT/Git+giqGQ3JIPWKzgeB7MPT3JoACPlb2v
iKa1AvCSIEagcYaaWoCApnvmVsl1JuM3zfd8/ruwdhYr0zut3c7U4OhB6tWzXw5qFEr2A62b9QqJ
xymzXEm43wvXSIbjY6lQg5N/qP8jNsEn62WNegaMkmP16Zq0Z1u7oLWBVi3d19Qf5k8TUSMXCeHN
t0biCccPpsOMsEEk9swYC87nL3ICVySCq/I7ni6qRNY4fY0yqIR4pnIqMGyBMkNPVe1Hk2HAanYY
OFshNdUV7LFEjKYpEUofepWXeBmZsajb2/FgxLwzwaXvbgwLYN7qHBoGYAOwQHopdV+fjB28GFcV
RQfzWKwo8tWuwj5pRJnSKuJmvxumXoNi2Hqt9vwUd8HMEaznUl7+BbH/f26VeHKDVjF2epM8oghJ
wpUtCtljsBxx2kqZ92rZNhKrbVK2fqwHA6dbPv05LCTUbOC9bXHWUaG467Kcpj5Shu+4gsHc101y
0rdcGlx+upmJexyHTUMDaElpOfPs1dLwBc9dBaYv39Y/gBOJXEqSH1wnTT29ZHxxTc+JDCMUQMTv
2GOq7q9p/as9ZDyK67UKZOt4veJXd1cCyybj4lLHRQpUgWjvz07W7totstuliZyoq9k58hTdTKqP
dL8fk8WB1D0uBlMdU7a+/NfMXIR2FF5P+EZMnnf7BlVsOs93ome2pi7yE0ZZhCtoMKC+VG0qHgVr
TysXymhCvRz+jYo0pUtGYiW+21YbXLCPcLo58v9i1obLDsujql/7+u1KObHSnuWxF8rEKUnzM9o1
wyhTvKktwPaJTDxUMtigrkEv0jtE2/QK9aUyJk4lQ2f8lnLDKXzqBGOVMUjOquK7dwHSb5ckTiVP
Pelo1CpibJB+mtnXxg/4UPrjXlRRW4ugvzOAywSJkPx+7WVZNLVYM2Qel4B0UiZ0RZpKuo9FdS2T
4CIHwbwEwG31ty5tbUB1hubejKLQz7o6Jro5p+9mIPhYsf5RJb7YG5vK4whXLiwlDCT+1Yd7fBOg
IwPOAVNW+LPnzrl/X51HR4UsrP1Lmotn9JvKJUVBFQwiUXLhiekRk54GDrZlepPJXH4m9ZuE0JKh
3lXDMaH/K66+rS2lZj/xK8+WSMjQJuumxnD4n+8c5m0FzzxXGnbQyzJFa5xmUcleVMFAg/G/cfaB
ywklwX5SOlbTeWACjY1LO/m0+sHGrLwUOXaWvPW3QwjoZXoqMnIx1nuy6CUOMQovSwMIc9iawH2e
djd1cjYsrac5x54KT9LHGoVS5QxfKks82ReowwQjhwsaPKwYMQzxHqCelPPbsf7lmu6CY+WKadHG
o0NVQ457C0XM3DrcNYEW+Mn7NFnnJDU23M5ygJmh2sR3i8hYXJqF8GH75SC6r1duOTLAAH9Q6TXm
JfGNtAiW4ShvfmfnfqXnAUpWUuMwnwRMLaEv2qP9vv58CiZofk1okoC49snlKNFq+6kpJ08j+8+g
1aeO3epjLlJVrBtgxl3fZNhkRiY6QuOP+/ax9r3vtsYeCmY6SSdYrozMOlrxqrQR8l5rRFN60Pu6
MOGTvHhDMG8hRrvEqWJ4J5vH5s6/ixI7SJuVsz+XlBnrJl9awSG0A7atWIdQgMVdN5UewvTlepWH
o8LsB0lAUcV9eNOvntdMN9r8DRdyCRTzZ3G5Pix56CSYf8CBmFiaUMuGsX1SpM5d4lOs7NDR/3jC
lI+GrkUk8+X/uD1GcpAMfpmGYhNGlg8J4rh7luwT8c3mIAnzUOFtmo75LEZ6nNZbewAwUe1f4G0N
IBlkz/0qfuZPMak52NLciFDW8+ozk+dltoXrQX6UhNdy3NLzGKtoOrQkMDokLTgHyPIQ8wLN8dIT
Z0mWtpFYnFTg1ee9Zt9nCbqsZF+cl4rH3HomF/dKqwIYNJty1hpoN1jzckMeFwKh0+dwbH8WXC1+
PS6xyLAPPBsQ/Bk4G2qynDgtlCUjgK41z47TLkYKCK2f+sVsEIbGULcFmY3MQyc32tBobwDozOJm
x8uElvpLntXHe4LxDRwmNJDMBxVD2N6kI0nPP7adkDZAwsM0Id3F8pDynT9/D+lXdGtO7u4cP5tF
avDoEsMYSFPtJ7R9WkkXjcU2svMWBZZHlj3rrt5+vFefJ4hYoSLxwNQKJC7dOWQRQZYcyyfyuXVQ
4w0hjmnUZdn9yd38GMrSZDusLMBBGm+CsBDWKM1vU/zvNdJqlQO5aAUBFzyKoxH0CXCxXPAZbMdr
8wNib0K17vECnElKgoUXLINoaebdNqui9IvOtm3IxFhWr5AAdJkQfUdmC24Rb30PahWdV0pqNwtv
qRL5RIIsXCMw8NBfHIXo2+bHM2nnYTxu33sjnaXsQkerY1RXnJKx4P79CAM4lce6YZrLipIpV6rr
vntPG54O3p3BPIByWlkhLY/nSLkzcwIcvbAZLg38GFnvXkResl2a3HNUdJyR0aYJXHBhwIJ6JiSm
n9CBU95nMvV4bio7nT16yU7rtgXD7o29hDRTANbB13efJUffIlPXlJS2pWqIN346q7ez2yP1JsJI
ghezSDsBGNivTPZtpjZ6Sa+twkbhcJ5KFZTVIJACFC0oNPz0aBvfxOGK6WyJEeyFgnfu03ohitai
vUfyLrJVc1tLaFNRcElFnv8WK7b+ySwCBqyM1fAw/KW0w6hhZFRsvaa8kUhGVdNFPOGCkl0433YY
D6Pp1hvoo/1XxHBJAJ86BqXeM88CWUwJ5tIPQrJ/JcOTNJlFIMR7Hua8e9tiE8Exl7sn9hs1FFXk
UlCz/ssZUvRzRAk6r2v2ND34RdxArRYoEBogGvAr/dhvnPj1Nutnp8eL7JA1OhN7jsrGzw8tpIRL
ga8DKY4FoZwPfZA/hjk/hL5mzGDK6ozhAYEwamWeVEncujj0lP17hHKivoI8B7NHqnDjzhI/SZ0U
0g9ui10aEsCIOTzRFY7oMdO46FWE9N8NU9e7MUQ9RF3S2gbIwf48op7oJww3QhRNMCM00OiUzpVI
SIw+Z91oFF6VIZPfewEE07K8q/klQ/vxJVQE32zVOeXEHGbNC5I3kTznAuOfxnDdm/lMt4FezXZP
+KJ8Hnq4cgFcVXmI6+qob0Aw2h/HGU8y1RAXhioYxp0HfRNXD0XeV2895+ER1lWwrOZGNi8gJT5J
awp21CngZUq816HEpZ+FYgz3ZGaEE3sIwEkuxy+Yo0KGajnmd/F38fuJYityJowgm+EO4MVVc5ZI
ZtMx3xlzOXfBddEAataPjThPETLKhhIK42xCIjYamHprps4eC6zhv9wU92oS0AneynqzymLy56Z1
WMlRP84OL9STFLvO242VIANiSM1nAyu2QETfMFIOIKNwbpQvVXSfbQ85jDZi1Ykc96OhzuBft6wo
agcSHKlFuntatAtsOXtBLJZsXSTDqwbCPWDIx+9aFXE00fEObxnu2JLzyFustmgmZUk8eNpXRNpH
ae27iq8YROIfrTmB6yxXHbfl1XmB8jSaiLszywTa1Md/gk3lm/0ClAxZ+5Nr3Q6RaTmGF2KQcm9S
68G6uWXGDo/B7xPteeLBLtbh4EVvPfm/hiBhvsJ0LaMkDIWBHa4X0NU1AlWU3SiILFYZ4GS0t1aA
OIAT8scwztQGTs/Uc+FoVaXo7u2A3r6wPfrXN9/pz+HBaPLRBiSe1d+S29mwGKLJhy90PUoCoPCv
wlqfxSm2EHUdnb+3L8Q4cqI+eC5Dy+hENXsyKnSRz+V8wyA16an9znT/VAyWu9aXirBvU7UUWfcL
3CY+mlHFQMtjPvt4fn4n27Wtrkw3hlYtL0KIZMzjymsVmOsU81vY/D4HdCYvyCe6nDBDSoRK4xYu
7hUS15oZJ+wsOkwBozu/50emfM5xf3MalJ2U1EYGw5UnAtuiAFTyOX0mtLUkhVHpYnY7IMRDNk8Y
a5pqq48QZiNVcVyPU3Hd8qRqGIoDDxXXqi7fLjuRsGWaY5tg7tbEzlbYp8tpkwhZFbHxRVKfZEB4
JdUVAZVGeP29tljVLKfdXM4QOnUehGCLagAmzUDFoDyOzpVqxXQbfUU2EZo55Y5UdCp6aAZG47ka
iW8HnfhNIqhX7Y/U9I3Qx6+81JulEMa02TiXRx6AKq7GDhNzhkaIIvhDLyqJX0BUH3YyPqOM57yh
LIHpc8fQzzbyZQYi3cVJj/Yi5JfFZwefYwFA+UCyv4BfzEy3ZZrR3qjWOFibRmb0ayM5zFZUXpGC
0DnoWssTM5IbCP62Hw9XpAg0NZJnpzHwri9n3ErT7Ok0V1dTRuoecJ2XjbQ0MJkTB8ICeiYt4+2h
PiV/5uwW0wGQ6c9YsFAMjVzYbNeeIQ/xqMwzFOJTopdTYxUYm0LDVIQnPmrkYRLvHWbvLWbVpUR/
hnMqGzuioQkPGsJEWm6vatqCfcc2Z3FBlPPfE5Dvd4n0Z+dPqroDXTlGyuaseP3jU0eZ4HnCRZuY
v0tov4ooXSD7MXtvRypQdaBnEjh/JN1pmUsRVbrOaL85mjzu/6QaLKglljyiEPrQsglGm1ze8uLn
l+XrCvWAmTqJSqvN1nyczh+y5EZ4tVNnLEw3Y1sH1d2q7FKEYksxo8LnGsx6sD/cB6eGLVxMqqtb
VmNsUl75x4+q6Qq42M0JtwjIDmxKy5q1ddqyx+fGIM0MKdtIz2NTOLX9SZp7G4Q8CLqQZr1Xg+wZ
ZgvBTSX8v3iEZJYAdDlMYlB3lz7x+e0w6yqeT9H8dNQHauUrPDdcYRgv6sFJ7iNDI3hlneBf9jMV
VrwYsknj9hQROJCA3LHL8I/GJ0B1bppnkQL4sp9aMiyTmpE7QNBctLhw4iFUkztmhk46o8MVoVDf
Sh3BRBzwdpOzBUOs0cMjSD21NT2sHAJ6+kw7g1kLqbVc1ESPowY7FwJZlNhLFDuqjHhiBWlGOeR/
luCd34tDf3jH/wBTd2kvYg4lP8Yca1/Dr+Puz/FSbfEAKGD3ZrD4TXJzgmOK+ne5/RX+iC5e61ZM
wN1cm3kKT02bCRIiJSu5dv0rA4XeglW4nDtDNuYrU+JBDVbmxiv3xqtmWxEZM8hXbUmZN2kzWSCe
1PLYF/gLcNaNZRFrnIDbKSYh8p7kqGexYiYzxn7ksYgZATgKiSrfuZmYJHemdE1wL3AVJFQ/ZBp1
ZUaXeynPERcvqvxZ56/Ysljen5KkGPHfRbVIXby2gkYEG3sIz+iYG6oO0VnodOakLw6EH7bMqif2
z4DA0ioarU1r7sSOpZj5Z1syPd6+c1fbT9I2Hp1sVYd6MVvXUN8p2rWAXJP2iUFzM860qMMmxNRY
oj5wlh7Tff9iqyF3bXr5+Z9Yy1Kk9fcaeswzPMGVvFt2DE3E3wmqbh7oeN9PpyJUvSBAmmoyYczM
imC1mMjPVZzas5/dgv/641kg92wYtuj6MtuqBccbi83yq1BAuHaoSHNDrSgCD/vgrsQrOab/Qlkq
+2Ozv9FaRQ1KSfMKl0tgz4p9nJqnUbjJgruH3iolQ+e8YNkA6QQB97ThkopBIhdUessmVDlcmhYz
0kVf++l0ezRIRXqqqeb/B712G8P/3Gxq2ZqBn89cbPTRl3piUbLrotlY8lLvBnKvmp+s8pzN+fRu
mGHXZifPip1jaluByPmP6Loi2EJsAjXJ2v2WTUAuKzwK2IIJ3OlhXGzApBucHGiCd1jHFxL5XIhT
V12BxJd8d+PL91EdvtXzHnuoCKSP/+/rhnNtM8YcKlJN3/ctKABPeM/2giD83fkLz+TW7RIcXClb
d2fxzmXYQCsVJ3VMgeNkMgdSfFJI6mP0RmGNJqXXQZNk8AMdF8nA/CiuGrlhCTbkfXLZGDkeOzJm
E5c+1Jdbz+LT20l0hueaNqo5/cQIm99sTtNNfXD+Z/txfDyWG40D0/68oAH2x28DFfRhX98T44I7
DVKhEMfCiQray7lMpDXN+UAYJIpI9AzmFxJ+cQzjCK3lQPhjn3/6Wt9d+MzIwrc1FeE4s/tIWhz5
4i++dFhyU4tfmeVsKMsE4BOTU7j4QxVEWLn5XcwIUzDRq1Z6P2f7XTOyqFKwkKNRr+17VyZaZDaW
pteRImLwV62tZtaMIRPVVMoQ8Pjw5qmU+eGz7/nmdAXwVQ9GF6NMdwxAOQ6gG9qwlpB47gBqv134
HtEdRZ3MOSMjBjymtPc39aKalUsgBj6LYLJil9Lakjc/pUNVGw20zGVKjkWZLSYH6Cj/UPTngCRH
4FaZnp1ygYJ++4FKY348kYgL/k7zPxk0KYT2jPtlJsYfL1RS2Ki3g3e8PpgKOLwkjpaLLEey++3m
I03QxpSMBX1waVA8VWSABQH8zmZUz/wQzy1Q16cR2MlgnVF50sF7HziGTYbtxSP+6TOhOyRd9Kkv
M95xJDITE2KxsnhA3JMRv6Cnh8AuR3K3MsvLaYE4gLsh7FIw4o72jIwOZDziySOF525zBJulP7rN
Ru1KSKE7S4QuAoRkh2S/tI8P0iBSzKqgNuXze2F+Ys+HUBPn4TinNeaXf/hgmPqfDCb8lI/YQHeF
9aBpF84wRtzHCaoJky7KEZZSeG5i54+3chVxhLRsRiiFXC1BlfXWi3rRnBongVvWBhc6hd90zUVZ
ipXTb071Eu5vLMdDmK+kv2oMF/Znj0tVvSxiz27xk/h9SqgT6Cu4jd7oY0B9pn2gA2Rbl1+WVIlX
HlBj6bpSgiDWJEQK9XuDW+zMZqjbqPHzYzf6YeO2dzOn7Fkp2zg9F7VzR0fPIiVJrpUe/m8eCr/1
cwb3KO7qGH/tuNYrIDPMeGqzQ+OPgsBN2gp+wUjcSzq1zx+mfDYEOOc/J3hp/jR2ir6isIYyPF83
zGXUTFQpC5UW3syC1g2jaa/U5jksK9sVvoWONIZyWFa7nweCJ8u2IS+CHeZplo2bRm6CSswy4uNn
bjCktMt/0SqoecJB53QPO3/R+ZCeZSpwRW8Eg2GScjrGVd6SalLQeMzHq7DnwwJgfrruTPND2hCt
ZI5/Vf80pyDYeO1A09e7RYu9Yxe/08oaiyXNG81bZPRH9V6wMleIRVkuAZnsBrQ/g1pnkMxNUz4+
i4pRP7ruap4Qqj6kqFzrzPJsuxiSl9/IOeBSCSQF0mmbI04wWR9wsriJpf9Gw5041DRF9OmcaA1k
zIquRNEQsB5WT2BDC9XD4JyvsivMT6xVdECfx68UG6LSMc+fe1I6SvBPs4TryNQKYc5g/0gfJNKl
SI95SVzaykKgjUXAOtw2y8/SwcApduh+IITBZ857jYUQphyabUQ2/S7EMJYNUQOmP/jaWaNdAmdl
zJsU1BTK8vknAvj8fHL6moP6KnRRvMmKsdftLLCpEcPW51y317l2ay6Rl61Q4SfeJmXYnHmZlOIh
IgwVbGdFBsfNOljNenDlnY7Mz8NTun/gwMoLw7FejXTA4JPTfOQG4Q+VpxgTf1R2Drrjmsw/BR+x
zypk7y2p8daiYJtlSlBMS8C1Moyd0cB16wj9HBu++GmHI+BkXWZgjRBp7ufDd/J/7dzAwkVkhNPI
gU7McYdyEWJZk6VPGV9xrGnccKnVkMM0XpmIwp+GXMp9eFqUrWgWtbvEgVy0eJ2SSDeoqgTyvIuX
M8cZH9mDYeiykAB4rl4q+v8wgElRPS5rjRQHmq9PxcTJy6w2YNAkg/9FbL2UN13RJn2nqKyNtdJT
Ijz9F3sY8UIyDq5tykoEg9YDtUDLOFm/SDgcsyRa9+ofA4wWMuZHMaXqLrmZjx2OBeVBLpNOsYz1
Zg9aS38DQOsZDcld7YjPdK4VAi7tZsOqP389lieFbtYL2NKY05oG1CG0LY6NYGhdxHWXRcTg9UU1
LJN7KFMvDVPw2JV5rJoszYuZVXRsGN+OETXpqGzuQx7lwjEztrX7O0OmV0ol15RMEviRf7iGuk5H
lFwJLTrVo/MS7/o3jM9jl573TnuX1qHp9+PuMDvrZaNzXaMhXqBJH6H1cINWKa0fiC5qE6E/hLlg
wrI0qLy3065wG3CPY8gzR6ZQqbl5vPhg5pLxRcKiyy/EATCbyfB/Um9QIfEDOXXqowbIe3G3inA0
ZZ7rz+BKekM7JTc0DyAoIM+SHOqf12slDIFQVq0x4lNLZsTpS68vmA8DAEcs1I1odVJpPiMGVYh5
JijzqN6qmzf9X0x0ZqwTT0yLsaQCSSCfpo8sVvqmODlPZcFMhF8fskqTUm6qXWlXIDU7W3cvUp6C
P6Fuv2xs08DuBwppaE5B2vuhsbEMA9Z996zQ9RMjoP/IK9dFIKX6oD4MgpkcNtI0tXVZ7eRqSMly
RpGf+tdJCVwK4iK/3u4XOFqhXAJfeGSx31Lc6NGIPc+MWAJbKG1ORL8zZLwoWK/b1gOxSgShCZIy
0n5jbaZoOH4uRi+ieOjJrr8AqfeKVTdqje8tpapFYeNATB9pd0IntFacYdLt/BvV/X7SXoFxdNUh
0nkLgM/Pwde/mIwq4linLewoNt7YYJzTmoh5N91WphZniTQtCN7BbUUZ0RGC8qVT3NAmUT4R+nUJ
XTF6U9jKfPTEcgYLNGYJ6/nOI9hWO8wNp0Tatj2xi3GlfaC3Ozq8KWm1lIJH//WOnBRQnq2060nR
lXNf80Fkg7XPAXQ04JPcZ6y2mljULQWrwh0RvdCc9d0T0EU2xcizafjPNTx/alkkO+JkI+vw6/fO
8zDOUFeTRRhSPeccVTEoJfAEgzBi/gabUdID/JUsrU53AiIXIOxm+IKdS7fogofbcZZ3qqTCEE1+
RP9dOobpqHKTnEOiyQV+WGqRCyUTrjb+LN+aJ38yxtmDJZNwnhi1xogcsx6Cg3qXdvYcFSn9u65S
ss22BqD95LSSBmT5xj+b1o7XAHO2uHfWJnOUEgE2StmIoEV+yflgDh4+acL846r2I5BDbisRIz8H
iQkCZBSKjInAOKDmgmAn8xxNvqNqysubx6tvngVC1OsBBOBULIzbkYhV1BIwaW46/zldjy3V5TL4
cWXmssDl7Ug7aYBibOOFz3LHGut4IAbbFE4l+u3nTX1xY2xzoWioUaYp6pLL3wekkDHlqBAsI9EL
U69Sss5C/Ela1pC3pjaza1Ve4LcXIFIlbthqxE8wBvjHwpxFksqcZjxSn6g8Zby+tNF6LNoxgBCM
XeleLy6XhlhfX9MRi8n9CttpZME/Q2Ag00Iqlgru9T8nchKcDTGB48pvpeYNhKSsRhRKA2n12gdE
tJAiogDr1RH2m+1fWp6jzElgtTyKlDCyY943f+E+I4Fjl09oyzi6tq8vsG94sqfufijNWR/0nsm6
ydPsQYyf745MvfXwDSty4DLN/FBON+L+OTynhw+bJP/vW+B6CVbWaX7x71RFzhn8kZGpOPTwgAMA
ElWhrg6FBnxhbi3+YAfTaYBTFW5zK7TjRBzZtBVghVyGb2IqSB2KSq9zAcXTu8GIQs2sKHzAsZo6
0whNnzOh28/Rhmdv/wK8c5xkOZZ2d4c3CUZ036U6gpaXyH2mAfBSWj6vBqx+HBHX7rqg2hHahIEX
u767T8o7YNI+pYSnd6ZQXad+99Vx+21ANmtErl7GWQxi2lajQM87M3Xdmu2v63IRmRVIzG1MtMe7
9Vy5ndtTUw234iWDWwPc8EzOCv0e2j7boCAeU88NqUWeb5IAEaO7/YNTuHEZETogYSQeBY3DC99Z
PxcOWZEbGDtdbc/V/Ylrz6irpXUQevwme2Rl1jMQ8tHmA2ujX85tjc3v4Ccz+7vehwPJDcIJs9az
Rkcn0nNrO83CEKLyl55S7tjWkgVsKdRVQvY9pxHRoV4aU0a+VOqQErv0UdNUuTivk0+M5HnRUa2O
jvyR/wDE7EiCyde8jKN9USJ4gaVR0s+uQ76GDFRI7otr8XTLpCG7K/MTD+Ua571LaSMN+CrBCUXX
Pd/xE+Y6V4GyBqWZorbLYQPU6ijVxI7ZS1PHOUfunK8R/+q06lbEEWU9U+BZqoSGYG7oayTbcKU0
YeuskDh4BaMW+wm9OROHooegSBcY0y0x4ja0poR5WAj9SnN8uwqupF+/EFR6hXmhUoUjDBE8mEqc
Hh/G7kc0DGGaB7wQm95oC05QyNyJdP7dYqa+ZFQQfqyS/OF+laL+x+BudT6zk9A1BxPWB8fd/WYD
mRc1p8dETMDkbULdnhRZZvEhoEtztbpKuJAQNmeGfIEb6inr11go5ru67/0Hjy3rZlwQwdGJlcKY
RxeZiiXxTO0bmEp1rHMvEft4fdiFiq1BQzWhMgmPhB2mO/mRQvDYsWiTVbDIKphokGw0kIhNh0+x
88CYMmbWs1bGW864GYe4VQPpgwkRFNY8Thw/9p2G/3GunbBdpPv6Ihr0wmbGizQg7/08nJly03XE
4eCo2qRILfvdFCeQPpsqY0gOBQYp8CuzI62YqA5EwXcQsICoIHHZiDlm5YO15F2nvBhw2LMejeMZ
iyixBiphHgEqCgXAhr8l+jUZcPknxzP7wgCWd+tydLaCrurHo4lSR7BznpH/J3o678KSftFiKrU2
E+rCoIod3zerldslb6Pgo0TYnz8djFYM7AoLZP0RMkfPq7TCR7BotByW2A68k5t0AW19OQznbnN7
o8B4+3RoHi6i/hVFj8u8ahyfqw/X1C4neAJBhfT2a6cuxZ9xgA/IHiHr+Y+orjigDoxgRM7rLmBd
7HDHcB4F2ZfhVUo/NNSQfRAwNlFyAtEEG59Iqvkdz4OQd1g0QHaxWup0Wquc7o45lRIOs6LntKFY
hvOz2LKeHgAgdL1egxtMbA62MEKGritla6c7rmszC9BFcxmWUDsAcs557tS0JMuVoKpjzJjaKk3g
lr9nwSuWmbVtRzGk6PoXbYPE87879+09Y9mWpeSMH3t0V1XZMQ401i3uUK2qDjPW6oDEKfbTiWtr
9rhgjzCDaZHfCn+etrZZiwU5ULZqdLJUpCLgT+4dsLGwnuDHh4zWTDU19fxkxrYmQQIMJ6aRGkip
0LXoBPnjaortKZD8kuN3s562hi9t+GV0njmCRXgr0n3AZW4w4CUMtGi7IfY7CP7wIjMcjHGgvakU
ttnnxRqbyKPdcCbiG9FNpFa+9AVkn2OKkhzVXYyyytAzwOK0J2tZRuEglWKX4SksGtJ2qe8mgMWp
uOqeNGCvpduRUTYJUekYku7c1at7Y+v+NReA+ruUm2Y0hfw1w0TB8ppl3r3tnjuPky5zJTdNTJKw
Z5fl7TIYSWJwMoxvca9wbYUEucPWNdBH8hbu/K2kJ/h23mbRTuueaBZ6iYWggUTGRWO/TML21h3u
EwYwBWh+azBEQfUO0g6adRtsgRyUYiHXxgmpGgjl1cXFd7qSQMlU2rVF79DT4vMpwc1tTVgdIcO/
iL8X7w5UmgwcSSlGkKdRAX0nnvi9nKinF48qdBR4eXWxn1hnv9xoFGUa7jwzefgLgiak0XBBq5NM
TWbf6GkcXoZcIlxdmytxeFQoObWgzahrUYWPcw+9ceIuAguRY84hH2DyFXclOcWM26ncnbShMlDg
o2RVV8BxEKPSOUUpG3yAXTVTiV0ovhLK/e9tNeTOvDPkNmhRgwrKSzRgE1nXANmE58YRfwk1LVt+
rLHBfvj1qo8dwG/JDXZh35VdwiVfDsv4ns1d4Svkn+BAxnUskMyFzHt6ddKlJBkVXVQArKi6YT4P
V/fiTUgbMtktA3G5XUYTKmU63j7u/JRD95bzQXBjfyyzR3vlGikdiJxPbxMylbneDCzhPQSj0Wpx
p5t/9DgzieNUJ5DTFOAgVZ5XfH5IVRa61r0ESwv4jAPih4MogdX5GCbC8dMKAVWHAdy/RbSfF7yl
N9WMyb3GkqtFSSE1aZDXadOK4IulCnvs+4OPk95+khSz8cGUFJf7XRbVLfqOmuWYrE+C2ioKjuz4
FyLUj2hITZYE6Ybw7h+jDfeIlO7RfIoAZ+5QQm/ahQHnmIetUREiYIBG1rl9cAS2M6gBT2ACMRG4
qbGKzePdWThhkMMRgA4Z3sCcTTdFlMTIDzrtcHMVMNS1iSnBGRCTllDhW84kngvqb3kD9YCiC+7O
Za4Nh++ybckb0GE88nzXgScAiHcArcn2VXI8JTvSWT5P/YIQ3tNIn7TO5xeg14qYL2DGdEwoPmXO
RGAwCK1+njIKU7u9WuKc6Nrjki8mcaaMePGagrMNXZTSBxKpnkBIUtUUR6FsegU9r9ssZlEzKw+l
aRQACRkF/CWgkbjfoqJxjsPG9pYOnNcm/ZZLYCB2eFWAzyajuYxz3ZGSuN8HA/0E8I3Fc/IjUF6c
ejLHKu/KSSE6Dv40DDsRusT0o8rL45OlNq5Hq7uUaQR1W2XbN/Cg+4fpzgvcJlY8hAToA/hyCnFm
p/8bgSpmMeiADxSDzWFMK9TKwSo53MYWu2QpD0y8WZ0owwwebCpq0SduaHF9/xF7aEK7gwXCS8ey
MYJVFhTbMFnVxID8RuOADbCGEpjSQ1Be09WisG1SIdxYZaRqYPzRWUa7KdIiIW2DWbuyvyl1oPbC
UcDZg6d+v68sY0ykZArzYr3SB3QSXG3l/dWqkjCxp4dIeQFwVzxw5ZlEjYhV8ayaTDXUKNM4hnm1
FHi5Hjuw/t4+oLWM1ZkdfJoY4qmzgVHrADEwnO12dfRlidZUZCqlYFK3W8vPgZRUsGXxgOSZCe9c
ZaRwtRQV57eqhnKu5zDTpVTebcLj5KGMCZm32WcsJDJvdEQyDvvqxHwzPfwwtOWVk62O7bqCQSwV
wRdAkKvNeWhw+G2zhsn/0IY/LGALkTe4iDOKWX2rP+kxFSpVaceAO8jrUhe9GvFnA2lrgo7RlDXO
+hNGeSRPkoG9y45U2iNb+3CgYOqNiKQlHItOE/cKO6We3KEHy9Tqtio1EFmQ7rkGQskx01XoSY1H
avWeNZiYbCnPJznOJMibx7viznY6fDN62v2+nI4TUhlLHqMb377WgwSxAAlFmHvEnF/qdPXqXGa4
UuLhs2HaYOmvs0vDqAQbSoM/TeGO4sShqR9rCOH88lD2KxKLtsGhTYIY9IRoPbhZ+w3eFksLVV2r
TCAztKnNH0th+7s4z8+BYxo5a2y2CBwT9ZJNNqskx/h7516LziaFWdOQKIUzAFWzL9Nv7uz/J17P
74xgZjELXHpazWoUUVIkNZI+tzS1dwSrojURvqZ0TDr8rJjZt7/MOVO9WfqPg853KxCzGsijfull
ELcMNoesJSPdL4v8GP6Hymdz0ZY3Ju9zDbtUCBDZzP5yzqheQRsRygzLfmkSwgRN1jmkmFJGBYZV
ZzVQNL93jw8EkeiQ0Qb1MEGIKhQoTYPhxQT0rlt13ZtqOCejyo6TgXpkuQkJcCT9yF+u7Wj99IbQ
0cCRXiRDe8Pru/6cNnBOF8zdELKV5rJAT8Tpx+Eo293pvuoMHXhxPU0GIX8GgdduokwdDwMIx70g
nFsag5CagsVJ92OqaW0MhwtmDyoN3XytIvhy1oNBGWN1hONdD7sWAK20HYceQNwAK4ye663SeeUs
1MK4IjcLpG/hPch9EJOINsdjySfb9QB0Ol+BiW2nbqhjNnttnPmLVaIcVj3OnDnkC1IEDnPziiYD
P3I0ysC7qtwb6AN960XpnMa1KMX/n4/IlN48aXHs/HaZs7eEL58KtoVXTETdnB4MBvziU8vxoCaA
9s9aXiWVZElD2w9PZbb/ByZ/8dXD7RlhvYBJfhoeswzeyu1UrP7boFDHiVEJhr5ioaKSpSe4BpLJ
prAxsyTfn1X87JyytI3Zc8JXXsNG0TTALrarCphPYFS3kiif5n4TAMG1eLwYl1vGP0T6fEfofxnv
Jsnkel0TR92Sif9JwYZ85vb/JaiUyI8o/F2eaxa7RxCSRfwsFjYUfZDn3Wd1kXq2qiaiHzQiZmoh
2N00hnDILftw1Wl5dO/I0ukYSBs6oAdhHLwK+E2fi1YPRrZ9tLGtFaqpuxcUdZ1ybFUe6hmdruLN
V29JiYSz4LpU93Xqp2+D2whk5/oaeBeH4HPgxipAzlPj+83cF3dVvL3SbUo1UgZ4uz5avocqn70x
RDrvIa1hQxjLF95kiFGrxZ9YCgRM44Q4nk/FyhLUKoTBir4+3gMknnwT3JarjsIxPS3Qm32u41Vo
W4rbcIqZkkALNh2mbRX3AP5g3N1ut3vS9z8LBCvv7W5HeDiqvfI8gUm7a7BQ1Ja7rlwMuUlfvcie
cRRXrQI8QfKitLPSVvMUclC17BcJBZsCh4Q0DME52Stn2TurqUVcPTO9KilfGGHGebsua3AxD3Y5
60ZGVOSbBGO2Od83dLuMrehX4M/pno68SnrINNxoJRW41nbqaN56VA+n6EmRzTvfK2XMsdnDF+ly
8Kqcv4N0E9b1gXZkCkRs7I1MGfHpURhEa0N+Xw8WGcf5RmERB7yz9hG9RIjE/BGUoaZy8O73UUav
Q3ay7MM3EUdC87gD8vlByLzInde2xHWX7LX9D5ljdsaCCIYLecULuK+stlbg7YDmnNXSOdTxnPhU
lMtCJGyej31OfhkMamvLlyW+fBPUuMeq5I4gpVHeCGNPHY7r+40G0ALPMGwRe/mSl34a3WKsOMXb
7UrdIl8Ix2eVLZO3XnQowEcKEu69VCwEntBEYqQWDPQvZ3HnEiACDYwDZH0WVJf2Cl22SQRdSFo5
/uAX3Iti8CKLAHOsnzFIft1LisnQGLKYSZJI+WMd7iUDBFaz5m2GOjsl/T2AEsV8sTbv3I70yGTK
NTtlHF68uJ0j4AiqgSQtU++Vmmgy7O+gBascSTe4DLEf/3osKZYr9A232yk0jV0jKUrNaz9IaeRL
K1u2hpoWw2J+C5mSDTCzAAY9YjjfVi64QFlT/dhltofo7jxpnNW9SAkflyFjwuk3PS1ecpXFWLh8
eXzFgdAihVpMzUOAMR9lpc8H+eaWQRfpZO8ToUqtzUsP5rURuGqvPEbmcV3KZonZZOS6yrWEhmgh
Pq3pq2xZjKvZjpNv+vJOccpy5hjpKP10wNwKGnRzNPxLKaKilUXR9AT8lZyE//vL8+5DYsJVC+Wf
DBHzFfpHtRfteJni8zsl6vMIAKqwhUMdzuLfV8/ynS3c9Kx2h55ZwdF7Si3mH/cjUj5nf3XAMb8P
h6hT1sHA6VjwJ/Ia4jyAEulIsZoWZL9treNFZwzcVbFqExJPfsfMXASYyrqJo/Q/TiZfQyoolD0R
/MJo2Em5IXbOD+5wk9ngi90Wk8OTHV+4AIf4MKCXiaJJYroTAfBeCb9NN8M+r8SBsNrkm9O3yVy/
X6PyLoEYf2MKkEcbeVzBL8d+ZpbOkpUWXGxu/EB44k6+jrSlOVOCS76s54Iwy5DPuExQMPOjY8xw
MvPFwfQ0FZ6uRqnWQEh/0L7ty737CoXbevFGpsCDtLlJp5qCqSn+8hrmWpmg99qjHQUUQlanEAR/
Eylfoq4z0YNPRy51evBd2S595tkX5Y/mavl+15YXyj+T2lb4nIDRL9rxOuMQ18XfsGfbRcqfvC8t
ZAX+nI3DWaZepvPIhnrD2dcYlIZeHs+Xx1DU6sEwQ4zhn2ce9Q+Lqkd+bjkha20PEzSnbZEM9ehP
j02zrDjEtMb1ItS+dEs3X1LQHVYqY0ZGbYyNFUhWb9w1WiRjffxi3MoHlOORSKn4GXx5NP1ch4eH
ZNdn8pY6Hj2GcDcCdc2yZejByso+uYQ+pNu2xYwOvEVlQpKcmeuEFXXzgR7DVujzx5zrwU6Q6+w7
tX/4sEz+Rn1eWoQx+jTj9d5N0G2iDmpSTrFwFHzfYm2Ik6k05IZVSwmPh9y/t8sAMZN/k20r/bJx
banLoN3mqPbb+vhz6QlvRMmD+uRKZUVGljQFOddqM5IiJqt1hsqi3/7aYzq4SCnZD8hDMjewwTuE
3p4sYmQK1SmJKImFjkGzF+RXRC+9d8+4oi1HOhxWtGwESB+P86LEU4D7wnhr5IT3Qq8ueJFYpOk3
ugZea9sBXR0KnV5QEff+MFU6J2963RCD6GVORbiUxjl9HE9OWe1I1eM52mbxQRTwK3VZr/E5CkEn
D7SeH4cUypD5RVrqTxJrj0WJkG8Fw9AJ2YgVW82z5R2Ul7IslPDX013A4xp2ONan2lUmA08FhmKV
syAWKUmL6skpxz2Fv4dCvxC4gXuWuG4mCtJmENFG6yaDYCaLiXkif3FbW3kfM+/hl8P3kIMYKNjE
wtpZv63Q/7zm+vkQvtOS4hni9q8e8XQjLn3dI3vSKtH5P2UEAzkxlJsJAfVbrr4IDtqqJqb7O6DR
dZOM47FrUTaLUp3yGcRCIB1GLW6N/8WeCTvWZlh9jnTrIhXZ7OqE1kNmyezOTrZ1J225QlDGWvLP
qZ/hnzlVQjcw5JtzNq51ViQoSBTOGi5X9pjHzbBJu0MXdKij7LIl97Pj7OGaBC/a97POz4iqC0xY
imyUJRiziQBV2NTS/zSEhNDH9eCL7d0OL1CDmhJCx/ZXCcyDE4/sKSaY/9J2Dfh03ckSJHMk9XRr
6km6Zqe3R8WM7gf1PlvkTY9Ie6DZWWQUkOR45+h35viynXe6g8uGTdo3s4tt5LqYLTKyNF0uah/D
tHFMm0aejTZyXQEDXiyOs8LltC6kHVdEfamgb7KQqnMCBacRZ8vYSJvS779izWR74X9iYoPwrGgq
s16Gbj+V2f9DUF/i4Corz69dkReuB8TcYeP5zAUkRlVrvdVlOqA5AZUPV4ZIjocmVb7WeOApYByK
nn+yRPj4jVUu5f9OdfxMRTLFKfDlgRNPOVkn+wv+GDtTkh3gPTT2Le1IUETv1Nb1TOnXNT3oLxGb
HbsMf2qjk9e0jbp3s0BxeJFNJ5AbvTdPSUZNLySqJ6Vtl+J2kqQWpjTng6CIGUa6/05lNErqPcyd
CTOHNEv5Ergz5nsi3PnHHKGHnVv0dacfu3RcKLsNcdcUW7WMF8teNqIkEzwuzd1AC8aY8Mhau11s
UABTfsnIW4CZSuOjhujA1lPsMywgPn1wiG+Hfmmr/YaK6zkGHD7bqNvBRiessvp9Zp51ifMlY7Jk
V5PdQP86SxEYGufldGDaZw7nbg/zUSXLA5Ff1flbIUnOKC3rg0QTQZwEd4rF0E/0ZuwznjGSuAwH
nMpSkAexWii/NQiMLgW2ylz2uLHkzEgQXYWhGXJUzYz9P296wnv6DoM3IpF/DHazOiZ8t065ChYp
/sKXYBQbXpuKiS+GdO3DwLmoBYtH8cbRDHSgs/iI6hxfgD0z+Ui6TgF49WG0kv4v6zzDbv//8OzE
jhjAjnJg8608gKIm0dSZ9EpOdYvZqd46xK5LTXhYWkozVPasMpxEVGhW0G5SrIQnY+XBNuiLSo0e
pGKwNKjWNic/siPkV9+4kE9pTeqtfw9EVssGpXB5GEt2LmLDDzZj7/plWT58yL54aKTsQdexGDOE
9PXLYBVsRfbQix6pyiy0eyXH7PxiOW+VxwHABaqtAgHpHVrJkoZJsby2Rjf+f7CLfOr2uEshtF83
v1YTiwNbz/bbixZ54YmA/UN2YV4+5cy7I+2QkThga1ijA0zLRJMulIovqVwKAZPe0R/ab2lyXkf1
Pz4MY1HAag/5rM8WVH8beAzrN8Niyk9dme2jZskxfd0xmYKdZ+RXEM4SIzoCh0hJx5kXC2NGs+6Y
cUhL9IoQdmZnyU7gUAjFhudAz7VyOGDGL5KEseoIII9pa2bc3f6jj2xQ2vAEFYhf497aclv9vpHW
K2yoEhsf6EFzz/ewXmGalXYDSQ8L88tamhBLVjCp6iCgfMVhuyszuqBs70tLNOfB9BGGH6XWPWI1
VrOLl/XMy51oQXkVVSYTqBHd//bs3arTJSFTHfZ5Vc5QhuRSWhjJ8ALjOHZmPUad4zV2IX5VXtzV
qMx0bdbqoa/tYAycc/wMMiW0YormzWLKdmBTG1f7lngNG+WsCDGoUhUC9WY6vnQPF7Slx+uXAIgJ
skKGbOlbbEEFJ++WH+OO0Wp4cMgPBZW6P6sxHD4XoqV1Xcb2yh/xsHrZEZkl6ecpOCwT+/qN3JD8
Dt8oon2cLVNA8ojW3gIlgBZvkRc30bn9kZBv+cQTFu6UacOrph719DC7QtgSGDcLfy1E700cWRWB
yzmMTEYzCf9bXJjyriEe2kpP9js4m7KM/m3zmVfSjPnaL8RNqytdWBoJBJEEN3f8oIU533huHznI
FK03v9c34gaOuf2sHrNgYQig3Rj8dGj1XhXIU4yX+XHnnnNJf3XjU5RVYI166LRykqX2HZoP6Bsw
BDB44AJa7RssAsu66x5+VbCVfCaj44HgTy4Ma+xGIblx2Hh6X9Asrj+pLkwYK7KtcFYkJd/ThezX
NHbYyGj+PwURbe8Z9X2Ddec3Q1AZIxTas4hUgP6M87jB/3XnX95IPEgc0TeEn+Y0AMfQ5DiK7Sjd
bvx1aqtWJ8qLupVkaj1Ky7rd4e3XQ02/x+MEE4SbcgCJG07No+JdF308t+f3jCloeDYxWediQkLt
xoGL/N6J4TPqLFIgJOJ9/XoKl3xdpgiGJBONmfEsDbHqhGocJMcFPk/oiiOi6bnH1UYtzjjFBBRm
eHr3HBY265Q0Tpbj65PMfSR7FgGL/v948gX+BwNXHa6n6e3PIZrlEnGD6f32dVuUsyqUqlwQZOP5
ty3WnMGYW/g1fm3BSA/0V+6WYqj71b5q3YXaj/bzxEPvZlktVkueNvfMqho+xcIdI9XapzIUhsNW
K21DPsq4kLxtezTve6P4kiUweV6BaY1pQ58tABdn2pi31Eml/lJyx2VUoULS0YI6R6nJM3o1w22w
mSC6FsazHdYl1PzXJy3CWGRrckHHDat6fUS7c818LAp16yu/Vch8pg1NvwluU6w9AijjDJBImuvL
eOpgz/UMHU5kD+Wbzwva7jLmbPspgXLNHwsZF0vbg9zsC0cKxk27HM2Iw2ZhT4KLQFLt09dil4H4
5x8FXtCeKaiG7et3EnTdyl09QZywlKUcoNyY+YNbzY3mDFthRTutu8IcqfmMq8WZnyq5Y5kifHkR
E4Ykr94Iej5TSxkTyHFi4NApmXPG4BMMAXmj6fPl353rS9g7bKVqddoT0rxA7P3/smigEKFfqgrB
rAG9RoGOBAxNnjotFAFzo8rbBetGkQ55/o8Dg974edHW4lPCkJPaNPXkBYG/Sd6rUAwLaisq4BAS
Cji2U5vEDF0JTUeVyNy2Bs0L5k/Z89RKT5lFRt3WlyNH8OKKlXLcCoL+VKsL+Y12P+UeEwE/PyPE
AbTe5wmQ84WFyKGiCdxHySCfVrRY8d/WyTeHP6WsBTi5pbD+6Aj6RRhMlEV13fayoiyc1SetzzxU
naP9cjbLQmhuLXlCpHQYsMir1rOMJE98PO6xzBk9EJEmmOnuKp3od6pxl0YT7o4hQN1TT2Tr0z3F
lLgPnEbbv4sPQoqUN8SSCCNdIdME+7/82MZjijax1hu23ERofrRe05E4+gf5ueYxPOvQValB4ykF
rfhdrlwLrWq62BLx9ZKl3/6kDv+JHFth0xZ3eSrzW7aWhVmEfP9/EZNg4YP2p9br5T6MwX5CxIH0
i84tcpVIgGJb4q54qelCuk45kI9euHjzr8kVAiPELZAmCqPRsa7dotBJbj8X6VptMTRDVxu7ffQk
+5CeiPVYladkC11onj4EN9cmGQ1tst3ovJWwyEJX7eakqS+gRnPqYa2byq+N5nNL42RDtIzQJbGD
ZnaN1rHi86S7bbIMP4Q8jifpN4jZbBvVAn4an94/K61gC4b0JpkVS50RFzx3wW0VxOF/PFztuQB3
J+GQa1eh4E2Ijkils0E1uRXgQmrYUXt4pxYFPxwtA/AknLBXcSiutfJrLOoVkRtYEckkjo2qyPy3
aJIT1liytm/bVhIZs7KCsxMLa1D/Vr5r0g7a8QK4ZsHkq0YGNJDpniiRoLB5TPI+2x+AaT+mF+3R
7PvHJQd7HF3+9cwLV66mrGyKd68kK3TqM2HZrdtKSeIa5po28JpE8gNbThR3KbwYAYwb32/utJvp
FleeC6HcMi5b8nEbLHbosshgR5ualQ4Jp5czWTIxWtR3qJOi4kT8KkX1ymzfdDPZjyCJyO3ZAmF8
8GY/15zY7oERpzWhyPHcK5gcvW32fIcRpySfThHdPXMx6dWiHQjZcir/3lExShBBbzGK+Wec3fVv
hdshB1fpJuman3mt1kzRySLCE7+5kB7tRL8mTkMiKY2BFvaNUP7g1LHDn/fdtNO4IsGRziPIkIt5
jdDwB0nzgwVfUKNax5ojN5dj/nfRFaEVRbKILU76Z1DI5NC6YC2U2JCA8ENqppgKgL8hvOZzP5j2
KtOBA2UbXgedpW9AvPnuTWOB5slfivaYD49fzvFXkNdLynOtoK+C8fptJ5XvvunOG23MHQxY3PRG
t95jE3jfoYCxbPukVwTKvZ5oRwX+IKkrDULi6BA4TTJsCG684QbpLzhi40kRO8w/Z+K3I5y3ZhKF
bX5y9Nr2oXSd3rQuEDnrQssr7EOkrSM0L/YXlHbGcnl5cL3+31tULJRpsE3Lt1T6XaGMBOj5r8RH
DuIfNpVpabifdlYz4j6S7p2bHRV6cj4L8yPwlcbeaUaAPfICNxPRwmG1yUeq0zME0pyhgb+5uVNk
W9CumRWGVS+mJeg42byzWtVB7eU5ICuKH8GIJ61mgFYwvw3yKIN9SG2DGCxYvShczITqE3cvMJpF
YX76vIQqNHeq9cOSY4pliRBYKXbnn8zgXQcmEIulma3zEZcfAnkngAhy3ayvH1Lzijh77A7W37Yk
0DNpl2MIBhjtF28xcfcvNs/alladZ+YkZpj6STqA8LqU7rN5szQkC9RnkFIxHcup79jpG5sbrGMC
g7daqkB1tpQmxJvtk9dkVM139F3zzUc2LRqr2AO0ird4fdYbfNOLR9octts6BbAm99D4Nf47G11S
hf50Bz9mzHmpMMjBILszFcU7FPGXXbh6P4cVHlsLDDiy6M8fAxXIqha3+MYbKb6arCfa58HZd3vz
6BlcB241aQX0J5x2omoTn4j2OKfLJy+LmEJ0vzixw6h5PDTi7sKEL5dZ6l/NiJ9OKxg2/vpZg54R
MDkb3Sk2/OMnWh4hydO68eqQcdw1cCHpSqvPe081YghCDYFuuyvtbF9RbVrmtAme+AV9nEsY71b2
djjARhIZQp6WJRdhHjJqEUczCW/sNsakfKmO3hXNszGszxu7x6/jJRQ3Z6WJSlZFH7mgY54iyd/J
eSm4Ec1qdg7nP8YX9QAzFz6HHkgisQkVxWyIUY6FqEJkBW8qRXofpoNupytFhTNTfe4144B+w/9/
268PxBntmfBriR8nxpLq+TOiKMmMxHRjSHeY5P0Vf9R9/awluHQ9VhbyxTsWrADFVEzZoGCzY2uE
o08urzU0ETHYaGKmogs42kwmvY7xdvLRnJgtmdKMopN+L77eZyk2vcEgvjCyW/CboZTB7Tdcds45
fGkSeaAy6jnbGCHThHmO7UhnTw8TeGoAopX6muKEg2zRCEmJjrBkrziUGCWWgPhFs8az5z/rl7qc
RN2/wXKsY9Uqdw1oX/33phJLuzZC5JQu8raKKukXDhSchF2YOr23LqEzJSBSC5Sf0B/umt4ZHQ9D
p9PfQhBBtMAsVJPZXjUivD/3n0HzXzbT5K+9vblk5a44EjE8oz2r9SkoQMggFSS/Y1AGgicbye87
f9msAaUJFOMtPDrqFpEIoqneSIK/7M6a2ZyE0AcsjEVu/VYgF9ds562B08m+9PrkyP/1l1rFcdE4
5Ql4KTGrZaB0dI4hpeDzg0h6JuEsrAJTYCFI++FB9mezSJwz47sAWGV7HfEhIRw2mi5bNtOhS9Ss
h5suRETGHk2gqA2q+IrSS+HZRdo3Wtbt7ejkBMff50zeoOE5S87mVysV3T71kCXBvIRob6LmALkx
3QY7OJED83Nn8C5cWMpzQJEiDK2Q0uR5Td4WRjbShZaHN2CxUB91xUKuH26Rfae0RdtjcqO0o+mR
jGQgSqkP2MDoHT28H9MEG+zdVNEC1eLfeT3/AiEiwa37yxwURtEbonRV62FiK6Vp6to92ZSE4ZPZ
B/Cde/PnErhO+u7GREf/Q3W7IaiTVnli8Qn1VUPOJtWiNMRPqwgqmCucZ3BPRU3OqFdyF6qJX9EK
ybySpVLSLFMbu5BdMKfW8mtewSvyGTa+sIuaz6dzUi1uTKzw9a/+IFllb6u1HPyvtnF4vlezYpco
g3LOo4dXWGOi/mWnYha8ZN7ktpz9vXNtKZBu2/YgrgT8X7V2OHpsyj8Gm6WqfdhRjP02vGBObPod
mSobwiJdgaVJ4NzNTvM6FsSjEXLcdjK2oHWaegKwwfCkDG11EGnoeONAVhN0u5Qd0KKvk7vZ4HeS
Fuk6Zf1MiC6fbm7dTqtE2XDZGgqf6V4Y7jZxLYL3Iz3bXdSIE8MxjcYDvCg1H3VPMz9zuKjBm/K9
W6lmNGfmRd+ExGWrI+E88NE8tcSJcn8Z6Zyaq4QfmUKaHZKSNVPK8QvuZKtDtJJBlcZx7OXRSsGk
hs5FkkIXMHVeveJfAhg98WpXejlUdj3QWdowO6e105E1QmuvjJ4URVsKzfS05DjpEF3W8wH6k1Vz
BnNHyK1GCIRduv+31hos3J6Xpw9dOjDlfCFBazVnZti9jCfz3SwpfVoAUWFm7M8dDVw7Y8AGReWd
53Q8NtXrMcSpd3pETcPv7oE4xNIP7cAuZUnwWJs19qqw7JXc+7EYsoiablH6i+dOVDsDJ7i+5Tsn
6HTWa0/wF6garR0r9MZkfJvgWWFE2QnbtUZ+veJUO3QXFhgyIMZ+0BcBLI3QAhOTRVGtRv/k6HoD
XOtHqu990hEz7TynQyr6zmkFci5FNP59rJkUQDup6Q+P76NKTcMimiOJRSGlouqJbqp3Jo00Ljzo
Etww6DPB67U4xj3RslJOfDs6FoYLPMcKtH9Y6xnw1VW3Mh7Q8k9wF2orSrekxaFOc1wvT+y0+OZs
6LkAdNGRBZazBJ70ulCHqAPutqR3hB70yTMo7M3xWUuOx1Ow4JDySBOJeDmVT4LCrNYILAqcRTdU
NAIlQCirjzWDwcS4aokz6blIhOgdT4tic75LWgKXdfF2e3BI8AzHjzYOKqQQ2lPabmJhwnnqlpPh
ok/3Tm+hS1HpQc2yRS54gbWcIYcD8bNql5AUrp8mTBj92eZTdMTyhxoO91lVy6vmqiExulyLZHqH
8KQU2iPWLgMmygzztV3so6Kt14yocJJQFPGcd19BTtQGZ9Hdzyvj3GUjK9pxNZmTFpsK1QgiMGsX
LUCHtm8lXxemfhXsXOqhmtBtY2hldguNTDXRvVuRbGVu/KUXeylFNtKbqgg2167cpBck57e2HiQv
nutfDNNAZnNLjBcVx4JUjIIa995xX0oJRy2Vgn5SPUbeI6EuRL2Fx1viT4HfygQZ59kccsRqNvOn
6q+z0H5yHaiR7936o41rPINWsRKDk/gr2ap3/3cWfJdc3euqA2wMYddYPJK7OHkmejT2wNLAVPA9
yA/4iv7Zh/QeBMN1ZMroINxUlE5OQEr+zRVAtLscy/+/zQOaf1x78VjzFzfvgllufBHqY3F1iWED
15A2AsGcaP96egD3O4thX1UT7g9NQ19f14oZwoe0uPFLREkeaRWwWTeA44KRtarOhM9LRTFXJXup
8yIOYHdY2v7h+aQteAMY5XxMLU5rDXZdwjKuMWfWgHb3+ogGcdGDIMbiGiMgw19IlxLzqIoe02Ql
tyAhyGyWs5g5cMBCKA23p4Eq/1Zuj3VWcW6/8WjLyf+S4MTjLVAe05+du8Pt67uYKOd68r2O9yfH
BPQLAOKchkZSF19Q5MLRUqt4t5jPQq/WjKF5dIpkC7gTlgMLiA3EZTlPqxzUKyQQOkaeTPazUkAZ
CHFbs6Q+hOscQ1t9OS8GhutAHzs594qIhNUPLUAHQCyffyOHe7/BIUvTEasHBVoUJ57u/5CyzTOI
lHhLjSddiIdRs3z+mKRIoJVq/M7gsBXgPIU8NuKd6Qtt4dd/e2ui5qe1CygEQoOjbvnoS6pnl98X
ws2RyX61yNrJj3mT7j8We6AAFgRnNzw6fMU1JRNJTcaUKrtBXuuhizZE80X5W5xuIQ5dlkIjki4F
RvLFTfj9wpfP/6mtj0I/2UP3c9JBYfGMF4ribHGKgsQCghSh7GJ1C09B9kWzHPt8g1+4dq0Sucus
BxNts1tLVzxJLpbs0N0+F/6sNgtMzRNXLfE3nY3bRvEgTnnn3/xHJCamfQfA8bzMtFYnRqMXOH/a
omTHvPpY9FuECk5ebGOC/1NIHUUyrSLZdRfFc9S/mAT6/HMPYCIG19yp3NgvxpkLS81hRfdAkjYf
gNSUK+YYEgL3vhtwS3qVk0f+XNTQp2Iv1I0qpXM0VrCsaIlyNHISOU+3/S7Huk/5Nqk4vWLpmh2Z
K1KEY/hPmhUTEFUWZwCwUTlqZv5ciLb68YpbDQXIEmH45JOZ/bHglBH0O6kvl7D1Tkk66sqq9t4L
qSsb9TXZaMvSo4nXXRdE0IaifOqaA9h9kOmjVb0oBmokOoo+mtEQptCgiv1Pam0NOQFsIx+RSzHx
rISpZkZezkJdKKZkOH8sV+PBHVs/tDLta0sXsh0KKxZetxwf/CIniMrC/cp2lmNztWBJrdQsfpnl
ZZp/HnSGY9lXQglgyjexpJmmdYhXX4JNvesv8OPLVhQfDTzLZdJNYj8rIuUtG5fE215f0n89WW3n
gIUQuFVgdTw1hsciL43vu9KJmiUV1uLjU6vnamlMVe8znSqNnrFSSjkxfpXEuMuALba50bOoJKnj
oGWULJ6/IIiEvuJhSZjH3IR45ixX2wVpd+hcwBdcKSn7kL/cqo7fDsZiBIQZxkMvUPmZhO6mE7G0
5d+/lhD7iGJIBe5V6cisKpKKTa1BL+kmr33ENoHLcIPIX7sSdoXkBLXDwZH2AHNRGnSDMJNS4Yu3
icjbr2BMivbpT2S2WiXB3SmjqEQQSaussoGWaUJFfa6E0A3aCUawvlA78WmssG/jhdsp96OFCJir
ZPJmZIFl1Qq9Yuh3TKdXWjyCJKCt90YaCi+2NNSEnNQMaa6s3dNviDB+hcC8TbhOjO4kh6skHnbu
pMLYacIV+5shKL7QT6r1CrPTHrcjjkZWOx/ZLKn9lqS967cOInsoUxfWnaXdsQnjSNHe0Boa3Cj/
MJNBadHIxCIHEUIkqS6ifUhAsdRoVT+yQ2xijQYBsjp2Y/E/z6wvxwLqX6LbTuux6BfTWMAHNzZw
GBGj8fQ+QeSazvFM1n36lttN9Erh+mqA0ulNYv5X5EnQwB5PaxS0/NETIQgKSHpo2fMOYygf6IxP
6mHlTS7kcYDPgdxM9EsFzYijILMQ4Aot6mxRZiBTBPmXCyZWfvdfofX/030sNWO99ZyxqnGxZ93N
tWAQ0rSoeS0gHVpe0IgMjTuNAJZJetGjIhIOTTcnW2wpcqttwTYghrcmMorSQ7SyfJ7giSWUke+V
x5R4dy8BCS77S8oaaUbRPJCONWC0U/w8Vv1POJfFr5P3lzDlxFVDbcmCW0b8CcbzlqazM+e8maeD
32KlgsriRg+I4jTTjxwMzc2aWuzrZ/RXpCskA4puysjo7URrSFJVcV9yBebaccbFQD9oPfWDj9mM
ISFLuml48ffIVtrl5ZogQhHf4DWBdRNaOG/+rU/dYKIGToHp927oDErHROOlE6D1toklrCynQEI2
tB7WKOOmYDx/bHLDK4DV/J/fRH1POoDka1aBvVrD57ZHTbKfl6lV2Uyb3ZNWEBg+iZR3dT5JzFnB
5ri7yVsZg6rS/dPR+cjBPMUpzctOharYH+WGQStWYRW+4TnhHa197gQ+fAJrRrAaHXgPmABHo7OX
KPx7x8sQcOoqHCC+VdhPual3M5JianE/3oZohrTZE2SzKE3KF15SNw4pa7TKGWQ0rDXgGQPNHyas
j+SfCTEMryJvoolQDR72O1tewkix7374CAn2IZ6cFxTnadSco1V/dXfG/jrD1ri0xCp7BY2mXPqc
X4potMSmCkeMeznE/8Rl9l1e5bzWD9aKzzgX0OZdQgl9Kj6Pi/EZ4ezi6TRVldJeCu/2UchYGbTY
/nUn8IpN53z6a5wHiD1oRBru//oXvsSM6MpdRqVmeJxVuiWQthdkDIKRWWIW4Y1xOMLs5+DnzwJb
2ixjqZl7MmvhKA2QMrFrFsdx/ESPsd79KGRadT9ZLxAQpD7jf5unesY1GOVH796ej1c/QwxkzDPG
yxwM7j+hYcBFeswxNbMEZZVU3kJw1G3F6TblAPmIju/vfjpdhDXzutwv6dVSfyzhMGW/9+mDOz30
KZb3JtizrAsDvr6oMTJrRAv+IIGdt0pchfBSiLh6s4NVXJgKY7wJEstHi54VpJZYB1+mjvzX4sW7
y3mHwXip84nmhuYQYZTGRc15PMQKY/QjBETv+hEKCE+xadR1gJcTn5/oSEeOKScIfdEptOqOTG+g
PuQrp977Ey3AxD2A1J2alLoImymbxSRsbOlGAf+zI/w0J9vEDPkdJgzcdVP9yQeSoWQgy6f8Dz++
ZXhNobnQYDbWS25HgyUXs22pS1iBNokc0DZR//LvLDp5SMVwQEGr7jub23HmlHKTgIHPT4gJ2F5x
FT0VizvsTLIHQe9lznxVm2qa4muo9ztQFKOaRs66lT9q8mGzq3CFmlwCqKdsgjI/q6lPrdp8atOt
731YSST1UaSBYA5+VB5FIv/JKiPZrIm2pY5QsU2hcw1wjLns/mzN2J+eyGVLZ4Jv7SJ1buL5y8Nr
ARkjRlhYVaV93ZLqU7hZgu4GGqTeG8GvAEyn+y2dAhNJSp5HPTDap6tRaPy4goO3MZXz3r4Sb8Mk
FqY5wnOW2luUS1fCNrgBnYTLCnKdugpuLTcRtYOXRNxFGfBhVUIp0aglom/I16IllujLK/kIjPbt
gOlqDtHP9a1WS/qtWgaAXfk+dJpknvOk9rNc37tlE52bK3bkphJ0VFHAcN1GDDI7/udz5OlGvXrQ
U9dGY7c/fnRRlH1yTZK1gGjLMYZ0qSlMWdDfF1hBU/bd93OyLMDqyRtK3aiPfPUrUVTRFOrLczBs
iJB8In7ORyoYmdkzqhUANE319ThSyJyRNoY9XHglvvAhLYC7eg+ErBms4tXq/j/eBQL2BiNxEE6J
MkXuCkLqx8GumN3QRiqUKH1uu2YEYrfs/nqwbbnK1yxC8uKGXrRnqibrgqspE/jZlr1BjOp2bwnO
kKr9uOYzwsAiA7p8eCfjywDCbmaIYqVowOJchqaswxqsNZOYMvdFdMFHky5AbHJvM0RY74GlFchk
JzQIZ75ZFDZV6D/zyD3Qo7FzxxlTsU0BPPi6JYiqW1CmfRkHD6oPzEmh1DokHjm/Fmw9PdV7dcHp
T47vULymjk/gQUZvLHsOyhTIJ9/IgEopydWdAQjKd30ySLZwg9BYiKTgSiFNKyuJxu81/ZVeBnKS
Ic2h3Ib+Z93ZE719Esc7h1ioB6eynm5ygYn+go/j8ApJKNgzCiHTKH7Kcx9ou7+FEVRYEwzvHfXP
CHYYBJ+KrjaoDxw2jikd67HHXvccBah9v1xA+DnlFbFJJGfyzU7A59eE/PNSxa2xya50JrLAYy+A
WZ7fKTk5nToDpXId5+i+u/Lipivb8h23FBHS15rjQ2uvYsuJ1v/xpZda4w1kfFiqz04qCqvbiYKK
ahPSt2zS4J8f1OssSIkrTKoDfmN3JwBWeOvrbIuwdBnjWolSkxKm/kfM6ueqCsn4c+E9QS2RhE3b
kn8FzJO+ebixkhbRJ1kY/oQuFSduHzIwfg/XmWoCl1QfmG4qNzwuiIP3Z7FoiCPN2Hp9beqGKz7w
0ckNxc+Oy79bsPeC2pSeX7WdqvCsTLK372EwX/3G8JURtVx/QkokZNJbUjviehOJZIYe5NGvv1Yz
MdU7IFWqJf/d5D4I3wOxW31pyxD1hObzrCrf2sBFqmtHzoAeFGk++NZOFjU3+SS0UASs3COBbkWr
V8JHZtI9SeZvQ32LrrVAm9x6m88BzN28q1opQXsljdM87caJV6sUXyuGh5suBfRbw56e0Wh9N85O
ZfdUC6ASp1cO4STaR/EKeYLAb5s+cksLLbbiMDXXPA4Khc7cmJdsoTdMIPem/iIp0XrgKcUJFXrH
xVacQImuSIhAT6mejG4g1QKdQWq9D1853EPaQUAUuZcc799oHg33QBICpZUdQrgycS+p0biJ6xLt
Ml9N5NAVIMH+CI55DIAwbNl9ZMz6n3nqTCjiKskBQRUBoc5rJ409rfRT97WxECGBR88XQh87wdb0
yY+ZlIC/l9cBV921Z+1anWi0+DqckQudo4M0UXvI/R9YF5Y0tz/QLMvtk8lC7HrvdfVTdl3xO9PU
jUOVjxhwlMrBV0uYWkBd8Q92O/unV9o95AhfknNabKZPCqhjAs9YvMgr8DzGj/yv9rpi7ERJqcHI
VfcjoQx3+F9AjvgYMlnZpuMIN5EbuQC/k1K7Wlxqdr9UaWOU1U3FEx/1chKhUcV2BmouvyQCK+zM
TCfOqh7wvoo5kKLZ508+gdLWKfxqsUKADcEV8pLl/AhPDLR7ZSOQe+HtKAzDn/mBdGfwkI/Yd6z5
/vcNrPrxlwyUTvEdwHgUrLPXplUO008oLKjjKXSvZRZdoyGuVS8LxlLTVPr3JhGTi3YIBbG/ZnX3
GiKw5tPEVn9oNlFoaWjxQY0yt2RL6kPH8ADnS53sRNK5zHqV73uBzV4XJsblHT6Ruz5MiRKTv9aZ
9oZgiFX9QZlOCfqBlsYFBqVnD5WEobJEiB+ai7rFb+wUMeA+8mSpweGTSwKCd3XKTNJqXZpVXVPV
wK5p7oKz/HBZAqMOxzTjGGTDaIk9ycOpbXtpxzQAd1a1G2I7of8Urfd3cvFrV3vOpWdhulYywXYJ
tTaDXyMwSbCk0E7Yt+ZD9xSzX25NwIVJdbU32UmYasGxEvaBIp4F/5njVJx8hfTzCnI1Y99RSSMu
rKP/9K4gp38QEzsLkB6L+EWHGOQkVsgDLGgYCqANMc7PJGdyrFq3sA89LgDyHW+vteTtioRgVQWy
0SxJGFT5qrAdKMZ1EA2Oqw1sU+JZcMbX7/WKQ+LxTGq+vXeofin1Gin714jHHsm1Sp7wrDFTAL2b
sj0gZRo1vL6eB9aTBKaXElWFSxsu8dso7aUJWhg/T03yJAqhAlvqwUKQae7Qsf5s3pH+52ZbK/WY
bOThB4ZEUY1krCtqrjd43wuxa6QEiqXkRPri0MIl0q3UHpmcERBFClIyBpdE99XHq/WAzqbttCNw
2OZne+zRnILRpRERHk63SHpD/17DE3G/DybmXSbM/KKHHhYUbV1NvhEJlAP2W/GqDdaZB1nccVNT
u6B/f5w1Cr5O4JBaPMOw0XbSiW2WoFfnhJOv50TXe2KJqgoqKNV9ewGofHhLB4wsRV7uYpi4RyOB
IQRlPobwUIFKnSRckuzB5qZqUIgB9MKWmmYCIXDbQ0gS2roUR/DrVyNZ93PaghVTXKnXAM5OJvC7
R8FE1rW8dvNXHkg9Kl/sZXv2Io0EX5tJwgbt2PWwJlUihHx/qASSPmg889BVNNhu0nDXUz6mVb/T
Z8AM0YJBA3o35ex/os9EeXZTjtCC88td44iTeDyf6gxlCE7aVwZ9ddFFlirlUzzkMnEOTxOMokU5
doZW1xakR4BEROfmfFyZiMtL2/dn1srdEV/BaTmgJTRpng3/hW1uAtckVv1k14eixr0wimST4TGE
yhBU9Qv78CRXEVa0clOMc5EyGxm/Wb3XQ9kPvHlkLDGauziOuiPluXX0TLaLeSBsW8++Z3DuUhXN
AcsRAIxBdQCwy4f3iG5HTsYf98ZH6E6c9bAyrHhL9XHbyrwfdFKXYs0UmEN2hTJQ/glVTAv/Xwsl
aQ9x/u56JKdiOh78aLKiJTPY+JAD2J6DLs2IOWfN5P76fKF4kzbQXuwoJ/pOv2d3EdMSH9yZM3J9
jQz3Pbiz/LKkq5qFbd4KaIcLdeTq2yiwq6lyeRRQv0oWG7U6vhE8Ok398YRVCiQHKaRSyWCiP3Y7
pQm2+BCkp/yes5khoVEb6t9WjloGiF0IE/tOer1CO2qg0HGpSrZ1spCbd6qM6LZwT0Ion2G0klly
6WMeCkPrHjQvKD3jjRPug3d9Lbo7e2VNcQM8mKSes5KttXsy1WHw2AT6C722JR/xecEp/5j4p+jN
nM7dYb6DSGx7O55BasFzTf9EHjHtozou8mUpOQp3Z32vrGU3rBQVAzgf1twshwciJ1e6q6u+5YCS
1js58JOCId3r3/wKWJ9SOuBFd1EFXSnmLlF6/mggYxYapHwo7s3FJSpjGYhXaXWyeJyiNlKpXyda
HR361KffCB1AC58j12MsO+dqY2YOOa+pbaD5JmRAT5fp7LlqosLIXMydmBw7vroJMmkyDLnIOZoC
TrbSuRuo8KmQPu0uPECZwy4bka9XfyUBXJsNBMpwAXhCRdVVZwxM6DWzWVMM4n23C/VJ6GMPLo8q
kInAE+2uExqKtyYYvtD9OGgxOvShPiCU7RSIEe1vtygRdetHjNWHUeTQDyNzH+OZpcd66jSxiA3e
CJazS0J3DM+tJBUwy1sdKkvphhuB6QiHTvCpkTEkr0EVoF2BmdiBwt+5Gxe4WLi78ukbzfuiMXVs
lOrp6VwU23ZtWDvGnfJ1UltzFCpRMb9S/oVCfeu4BW0WYN9iFW9CAVgWVW23t3kaUfL+GvS+w4Lf
hILDmr6WNGXTd/girF4Rr2vNW3Lr2vTTFPE5QReHMR0xFhvgUT7qfZICTiv24nz0/pqXmGh2XAnY
XSrd4yAnbQsP3E+C34HI98W1Za84vwgLjFwxsz2/8mywDuSPe9l5dwYvcZ1qNanRQxkIbiolO1y3
KVuRnMqUt6gA6kBajVpxFj0RRT+lO+AAQPKwUIorrxGGVxXHkFxFs1v68AQ6ZPsG5vLt7JbXBQCw
8/DkecoURIm40iEvn1UbdGlbXECB5aqLc/pjGTo1P8ptizg9h735WJu7pVpEOweGjid7ulkKEO0V
9ywHEN08NOOQPm24cAbba/K0QmrDEDCadFJm5hzHCBpXY7Os/1i6CqIS7tSB7GRL+J0cV4fd9tgH
AeEv26sQ/o2J3vr8olSNeUpe0KOxI8nU8S/1X4Mlda2wRluMTo8pGIxcHeU4fkNFn3/wl/AXQfIh
PiiL8fNkZFBnlDamKBp9rEg50cCvba+h27HjOKvyE2EXBql7QKTuPoUlFyT3sNCtedQMrlfTJzvS
TgRpjKCBLpjV7lxbE+qFvOiO8SgLzKg+319E//sUxRnu18pEWQmYWtdqT4BM03geuZCutRz814Pg
hqCFS+yceeyGYejl1EeplpsF+WbZISnlIDBvzXWY+daBoZGq8vADR2XZ06ymmwLN4xvGeNjGyKQg
83HorN+KKHz+3uZpT9jf2GdYc1BdYPFmAqzGhH1iyzhcutcfSS2r5ABu5X+0s5BMRjz/eLK5XQgX
B7n7aoqm1ydos6ub5qtrtDGRr9zq0XdYOugZ0i+QcCqejvf9cMq07AdcQOKkYZmpTza8eUdtPXUm
TFE3h+gLPvKhm8XKZRW47H2OiA70V7sHt7XiXqJYrUOUvIXSFOpEq4zzBF4GwoxEhS02DdGpGIRr
jxP2izgKMiMc1k8U0FVeTVWi/COw4fZ8l7m++ja22ORF34P0fAOOCSQeDszpx6HmKgc2Jo2zMjlV
HqdHmcsn4lu6bMbmAaoJQfO+DNeN0YBe01KqPu+6KOpRHDkpVd+3pqZ2OXXDvIj4ez8m7QXbKLHb
E4KnGBwprD0r1cF/9+nZq1E+7zGwE+7gCwOqcUA8NBTZCqSeZRm/25xS1WfvS+XS4Nciz39TmZHE
tTiSNqnqemP5xSZiv0NxdnDHAve3VeYfWAApiWZgEs6DRtbBZLPpMCk7q9jAF6KZysmY7PG1kyO1
aqzF88tn6BlikE6ZlU5UEPPBxWSlm9pbsN+ehMIEbaeHYX7aEC9TRThagTyxuwW92yk1tAKiimGI
4nLiIfLoTluygAjHXARvp2eWRd7IPSphcNxp33S4H8v0Eg5F08DjnBGhO47tM7FHe9V7x+og75y8
owGnQOiz9ppR35L/TG0AFaFTdLLcXIQUxx4x3uh6SecWPHHevGc5Ke7j7dqeuSzuLo0+srOjoXKP
4Wu0fkSEhqdHJlYgUPiREDnBUH1nP5oYQBvTrB4ftoVHb6nxMdx9Q/hUyvAOk3KyF0BJMMKlLAX8
fBGMmghMYry+eGtJyPv/IG/H6+oshcmEK1oNESmPcYns034iBlOGKULDanHw9NXambpRGojnyVWR
Za442Gq/3Xkjbhwgk2Ga4n+25zhMOnli1UokRcvL/JjpifZcsCx76sQPYEyRrFkOsXmIo9trsef1
4uiRjmaz0dz/cG92G7UQJg0mz3BSIdqFqcfTjcbsiOPljKoYQZ6NqTnJWv94gVAsTR4DMDchm7hz
bEnuzgB4NE4HWoHgVnKKIKCCR6UK1zq/JTACX4h81/RraeosBG1TI5K2J1fpNFIUecuI8zOmZJYz
8dLG0jRxd4t3NwlIyevjoEtvoT4FnnTx6iszhZhSRc0J1jrj0uyBzCWX+4a1bkERetUTe4G2QT4R
F3vp9goehg+BmNbt/s2nVHHYILkw9sjKj1ZSReIYVtdi81tgah5dWd6dSAXvhoqZ5hCQDlMYZ9YL
CzCWtZnBccT7r67048WOEo25mS8rx/yzOotmIdmeddbWCE9pgGZ52MshFOiZdR+Qxau4ne+hCzOr
/lGHsk8jTeFSi8uLEnw3OTYT/vsDEb/UHKHGx0n2bc3mstX2SR989aNvL3Tlx7ank6hmO5fnc9Ny
7u/XQe4mJaWzWXMFZKAyu57VB/jwMerNL4q6L1i2x4HqRchTUa98cMGq8kxg9X3a7nSJLAPzAXXH
9mJButsl9mEuDQdxApiaJaAeSlV4sCZLPYORe+Jszhh8tc4sjaMCsQsHMAbkwZAeViMVnpI5EePi
l+SDKoJObg6oVxFxFn3awxmD7O3E99o00HlsR8Eh+aISqEUBA6X4zVfma/IGKEjmdi47E0wUujs2
O4twbGqE7yNK4WEa1wz1VaQCa/INSfklz6QkEf0y+cDGlTHlMx0vlFC2GNvj4Ms3ehujxGfoVmaQ
Tr4nLMixUFZ4qe06Z2vi+OtYpieTHywxnzhksWyxgoYfPJEn5ZVPCinu89ecCRgJMZzVZ10Wa8kV
RzZ+CNSF10ud9WqVaQLiCBW19kV3F5YOTdFBxBHG6YELjsMqFKz51dvZEzTMDSPeY/FMn6bIx+Xv
uewCkgbBWY9/sbNIPuoE92PBrP1w7oRTSiPwMuloopSIdDDa9XrudJqG1D2wzaJUOr3YP2Vbe+oM
Ebxm3lR6EcntcwrWAwc+zyYkDNT51Id6kZDdT8AJQs2ZQEpp4HkYvE5DTH4o9iW7Cf40gHe2Lyat
TrGJeD0oJhhA341/vtq3CNup6x8H5Bc6s0PoPNcWAz8rhnKsf91K3XkQY34vNm2qZIo0nKX8e1zg
Xq1ydD32pS0dC2Zbm0Acw8WuppAw4GdN7OA2HVgA4z+9Vvp5dSMQ7IN/D/Lox/2LXqV+K/LJxkXH
fEO2yhX1bXJLm2HZe/tp28OJ6y8kKOZZOSNIx7vAbSapEX8zb5xZRl8kEplo7ntSm9qdQPoTzqly
Jb1cX5XSAYndo2wX39rMYGhxnkiubAiKja5n84/2jZA6fpY1six4uFb3TFqJpI2QjCHRjhlDRxSi
yUH9TcoMb6C+pSFDstMmn2CVSIvcQePUf0NiBM6UJxeIs+bn9eNTAdK70GM8q5GtadSl614RFKRJ
I7WkPkmucdH9VMhfi/AldIURhPeiDMS7UaIrU7vtqRzAv+8d9VsUiYVRPYAcFZQKs5eff9fMH+t2
07/yPIlQ8HYTSdug2AqaGTregeERCXj4IHyL9AQgRadb33bxNVCVLlarKEWUqtGM8fWxLQpyPMyN
0Uu3bTIlRTulqoAUPmSLn366XY9sBJDgHksSc9kvL9nPi3+3tnyoBuO2RmbSu7368DAbHTC4IbYV
R3yRNzBBg3UY8bCll2L8cs7cfzVrRv/NOBNg30dXq1ub0dp0kif+Ttuh+jwHX0+9fNPplnhKzna/
CvEDb3NM/10twnpXOr+v6HpdpUG2AU52WKXEptWsgCwXulqDmL05C+t5YPSnPiY+0WZ4pbg5FvvW
bbhkzZFvESrJZmXz2QM7abFkS2GR6/lhGEHZEwfX3KNgSd+8FioI6gaJhxuDpf1Jkn4S0WTFmbYU
cCP9C0FjHwt/0KPKqnMtK0SfFhLBbr+2hMAPXT5G18C7thVpf6nZfcDEAZmxnG+vDBCQoIqfRNnc
A0Ri62oVlKTqUZc+NmKF3HtBSIBe1DCtir28IQb3gVrYTldm93T1zh9U2kIkP+jj9QW9vBCq/cuS
tqaodbuEoBWIGYj17I/oHePj1YSH7fOz8v1ehrTlT4yovxu2n34WpODPpxH12FmN8+oAH+eo7ilM
NIh6B61SUo/RRC275gPA/pDshSFD+X3CipOv5WxzSBAshkYK8AQ+sKsGASgp6kKKSDlQ04HZCqOq
SCNeWOA/RaeD25wudq/rYUa5o6E0sJfUslMb8HOXlwjyHyKPWMKtsmelRTfmN11+PDBc3HPjrERN
pk6C+7L6w7MpTIdmiEf3dGrQ+TgFKQcMO7ja+Fsr9yQgeJ+sWXMSyDE46syq/OZ7EkXYtowUaA0L
sRVq4NUPWKXaVtlI5HU+ty0Uqt+XF3gu/H6OclO/DPoax3hk+FcyFwUg1MYrPdfZ5VBreOP6sfQX
6VZOPHniM/m+KmILkPtfJTELTEBndx0oMyaev1zowk0x63JHqCXEJiZHlEMsiNIbtQIM2G3zn2Ds
TktFoC3FzNPxQYLP52F5taFXWGHp2AKsbUumY8dkxtGQmlp6780VpqDD7koqjjzYIJY72lv7X3o4
yI2KVuUFEVVXIY2M3NMB5Y2FnHVZW6p5E6wDtvytpQU/FZBuGnOP9kQdNgxtI6lZs4Oy8iahjP7n
ZOmKj3uK7qP6PY/sGtb6Kunklahl7r3eC0qmQlqRpitdlHR3v6aVL5gm/46sGn0Z2CyHmpLJhugp
DXmWf33aGni8wM+++g9nmYlTha+iLrOrA1hvO0a1EnEU+iteRwdOQujpRSOF2Sd5Pjg8GYzaMq8u
Bj3dWdSgh0MrULOH/EulUzrhqiZ2fwgZMigZgV21bhNe0N8gkeTi4B0Hz+PvrzoqyVE0H0Z7KK2L
5fwwhNATYOy3bpplWsCk3fSTvdXzutseR8+ujPkUOV4KLDyy33IHQ6/QN0aZGUWUp4tuoVb0Geep
RNSgn4Z+oVHVEF+X2bo/gzq2vTanbqz1L5tMFFaEi8ce7CBwVmwTx1ly5FWJsw7rAWLN3OiH0zJG
motbXLvn0xjd4i6cKa/iwsZoihvGjX73Hedy48P/FXYYhYVUDcgzrOWJHLdh66SPlZG5ddNFw6VQ
FJ+x/xbYjT+ZKNgqNnAL7L/BFpzM3Z5OmttoB9l700SEGMQ6Rg5vbjfi506E/r3CcmK1SmtOc3rP
70LhcGoC6oeSVDXO3TGUwmHs2EdbX5APIp/eWoDfXqKFdOK9KJSai9Rd8KbU4Up8eVLYxOL+sGyL
vCEAWVn0BH91zQAeX7whwB25PX8ktYDyYSHKy8OhDc4Waw0fhJcEY2FnbRESQyKP+SCc/8jUYmxf
UTQPxgZVri+HTX3Vc7G1hGTl/HDP/ZFp/0aPpVDdpUHQhes3YYQi+xzgjqgaF4sw8jlKS2IiXUF+
91Y7kI4Zf+HSBPUSL5PKFh3lfCfuKFSN3MRV8v5IiUnZ1zNgo76YKrNF8qe7rVenycnEQosl3ibY
0ktexnY42deKTs/GnlPn3J0iBcrT2vhlep4zA3KUgPdXbOiaBvRnxFtVPHPMq+Dx3JDlTShbPVSP
nGGzIzdCrPvGlMe1ZbwgY+uA16mJ10Zw/HGu4Z2jQKAWdKMvEBxSR5P9TbFO0IVlDuYjBA/qHMXd
48nygCVE5jQGZ49/vozCX76BiaZdLh1iQkZjOtBDIcGaIfedoIbKY8IKYc0Hbt/Nh5UE5LMU+RI8
USPsWI1l76uO8jnDaeUL7nxS0nW4MfjuyOYclzqzpI2CfMXHjWN9o0fc5wrYBQxMYCln1FLA5NtU
gI5a8m+cl4nz19/WBZj5VexBCuSY/brxYvyhvpG6RX/Lx2ooV8hnAKXzzun4JY587JBPEnlYoKIl
z+huvXVgmiGqrvYTeW9dKfhXZCdTnjmmgRU8Hy1dcXdkUjbUlpgfiOE/UyIbi+9GC2p0pOYkeVGl
8y9ppE7em/Sdexk4Nwd1cPy47XCdy+SmLLP8uzQg3NtciJ0iZfpTnsGtJuGOIrlLzKUi3X496xws
n7tA4aQgCGfMn+WxPm35PKNeCXFBzqX8fits9QsPmdp3MBw7pEyw7fe5VSsavH6gA1TEdy568OHZ
t3cDjAQmADf/LxpBslUrHBYEQiXXQ3//qd89oC1AKFGTBtP6vSq8SSdAjVlPB9mrhCgYu7p4DyUE
g7wRUK16vDtsGQpDHCFK7jTmvj5+gSvdoUOBvxGM1HytTilXX2/88rN/FjAOcqd0T7MDJlz0QZR5
sTGSMdwW+/9sRlYMOngo9r3xVAEr2szZshHJOtJfS/I0zDeNoVaTmZIFCTy/eh43ALbkEXkAYYLL
moO/vT0hlCOf8qwKdAqMJs7aJ+10ki/TXMQRKY2XC++Iu/FJuOb4fJXEbG+hjjZYmL9luISm3iTv
xq0gEVd6O3YgTU7fVyaOSTBfwmqKEGUjicD/P6u5JHWP3QY30Tb8kKC/wsxJ3XHT6+19giQa86Is
kZkE9pYagXW/NhM+iw1N9UqVku5GgEqrDGmG7NEQraqg9YWEUF2CwFUFz9yt1KiapaKtKVn1s7nk
Fbxtdp8r3itbJAbPpfFCNuawZikFMvmfmpKTDgcAhNQtcXblTUGGcKM5L6x3FSBqJchcyLxeDlHS
kAoE93w3nLYW7zi3DngVyar057NMR1Wprd5xxk7FiYuowSEKUeq75/mOMW4P+ImMvQ6+3cmJi30X
G/C+ua8U4L2uhfGwCLN+zwc2vhp+R3gINxmiDkE9f+yipM7M7QIF/jMzvhtLuHbF946LhgfPAsjf
XymvKg3/20K6ctfif7WHv28mtqs0UQlEMr0kDnmO+m6gnVUrFwRtwa1GTXBI8kqrBhUx8dXLVBP8
o59dMeKboXsPpzKRVJ5yzhQm6s1v8uRrMwuoE+dDbLfDF/WtamYxu38k3ov9XIjrDZEt9xHEA8Ih
2zrbY9U+zVI+U3OjcP7iazIrv5Kov5pIkIpVdC7EnlKW1NjsPqY6zxYOpOoPSxqHcSVCuEKBkI1S
IX1eomJaV+rx9AQZBdiHF+walHeubmpcBKDuSeFSePZ4mK7eOJAXZAAujbBNRZ8NkTBh+3Y3BWGZ
sdUXHx0Be+prnUgPz9phfQR3G0Qyi1rDj0/hmSuGDe36+fRSw525yhAIdoL7Jb+OLiTVM1x6ears
qc1YiVtqg+a0qGp/M0DWVSk9MEa3HAjHdZ5eiSE2xdZweaXc2re0ffHf51HWcjr2bHdGSJ4BfTXI
gUcN5n0Ro/3Zhh3cVm89Yuk5y87ebQfsfpumCnTxdgO8Ypv7K2ILzk7sCqQcT0vx/FDcKwgSML01
Zu9KM7+KB/VykZM0Lu6vV2dNxAqoR0lzUpOF9onBOH4Bgcip8Ysg0t4cVN2+UxPm3fbzGNf06s8Z
l1omapL+vXlQGkuAlOCD6NPjtHLzRz7almWQ/K/52GT/XROUdQEgimud/mir5qyd/wG0OKqTu1Bc
cen89Sa+/ehOmk0zD6j9kUGzcAlskpi2JhlZSsIezx2sFk6/OsXllMW4CQc4VIsOGIq8XSnEsOGB
bhh2lyQG9t/FiJ6eL7BoKhQ6i+Fp2FdOV9QPVKyZ2p6fEyxjBClWtQFDkcOp1NSazK1VvRLLwiCo
2pAfwBCm37lOTguuNlhI3O4cAZzCJodJUyU23zR3JthuO2ZTLjxvg6pRT5PtMa9S94efq2w5WpLp
5nTIl/pu2Hpz+2iMM+DXAJEwLLnShoWjY12kxHiM/KHX1PbN4DWCVza+smlHFI6Ao543gJ0ycyPt
IgOVvMvy4j/1+oM9lotNGkSJBA2q4NUBGfoX6Rq3nwQCd7tiDh2wuiZ/IvroLW30LELZCjGswenu
RZDkT9omq+sXpQG/9bxPHGthmsEv/AOMQBReOHF7XwkGJKV7QJHFq0kJXxoBWb27hGnsyp283Yty
xX9icfnxP/GAn0zY/lSM05zk/jTgF9c7MBKGGzOlsMqLBiZr6mbW2WhZGazXgOLs6fvv6thaPQ5y
fZ9th8PyYJLre/hXJ3uGqn5GH7e2mVg4Id0PDAPkeGjlej1klWdgn3jhmj5BEf0H1K6Zu15YdrHs
Egz05DWYW9PXpOzXnbGcz+SlRKMVlR1PnT88kHaSoMswodcAc0TItMXCiVL9MFSf3YyFsHOEm8kc
YT3THXKanvGowRo2M6DbDzGuqL60JVPLR30qNaW6g8z1CvWAxF3dCGFlOO5666ZxEC9sDUr8L6J+
3ggR/HFRVmphyLzoLI87jaUa5JkhkO3DoUZBkU0IfrtNwA2/CCGUnlij+CDXFyVULdVH7mgvBU49
uAfIRYk00bIGd872eC82VZZT1UatWfWuxGsLTh87OW/sceKQLlZEHgiCaeVaguXxK86lbE4PMIqv
UjtZxZtPb6xnOqQ4w/IMMPFWjkQ3VB/AFxz+J5PImjMputxP2ms5NYqrxDSsZxvTqEEyRDCuIqqI
WaaKvRFe5mUs5crgYov5NnEkSOJteBk7KyOCsN9UISMkc0/26JFUt/Yek9+jJdL4aJF5w7XiJ2AF
l56ITRNUaOYqYug9C5TTDFlTTUaLWUkyVaFj1DBs5viRZSNDuZ8iFCb/iEGVJ5retdi62RTkF70m
nAppDM5s+b9EE8TvWUxb34+0UeXvMYMYqo7F2L4E922/C4zHn092TUQYpuvtFb0fO9ePjrZ7KOkd
oYWCWhgp4kco9uKnOL/vILRoe53X7IDjORwKrojwHSPu61QKG6k6JqsutZxzMT+nSQUpsJGZ14KF
OOV5EQOrq25x0N9VaeY5kWb0h4UOllDrEMy+gjgMp9qyqcHgQSWl+7y0rhPkj3GxSo5MEqBR2QzA
0nnLfff0cn/8FsfbMMQlRiOrdUlxsbWCnffLn/6O5mNbd6xlnI5Mpf7U2tU3GFYUnJ2Y0tr87SX8
tzobCIWDvr5AWwVGUPC7AeRDWVQjHllEowdQxxV/SqpBwGrELQUyMPFxi1oI3Qi764BfvGAJ8NTF
ptgSnWiS8DO5FlOwgC5r3xGAkw1TXeuWNxNWQuKrzFlvQgTMdObc2sOSksznYSqEmergGfkVlYil
nQjTA1LfxiHrxZI/tb2gJGtZ59IMoBg9qeGuVk26v96Gi9s8DjTpG6mJeEgu2QkSeQxzq5lKRVi6
wCTxkL0JHzkEblRy24TZ79dOFRSmzRZ4PmtrZksq/iuf3m1qmzvNZNWsCObi/xTFeEKpFlJsJ3Ko
Dd9iLBj91c4tEz97ZhgoV8YZWIONhMnTiVViO9BH9aSWWsGpdHtMzdG0qyrv7mGMeCiLqjNihBTW
EzsWfnpxO27M7gPm0SM4mPNEeIFVr5ZCG4UIaBN4PuEzmp5t0AlK6/7c6pPGFFdlEG5M9EcfW36T
74THpqrTjgk/i+VCJCtnNo/7X6kybWMoIP0hY/MRwSRrqopI2siU0sHrMi/spL4FL4ZUmXdLpPS/
2gJHlgcdTEFiFiu2mVUcTpIyYuKbpSMdzKkasmKM46wZpC1ZwIA2cO7xYbo16wUcZrZ5OuEFx1LQ
8ZWpvGr+Dy7WRF6kE03pcXBy8znC3Gpc5WZlv5t8c2StXPS38jmdWlvsmzBVmQ7IqNoy8aUwaSnY
21UPea2doPJiDIdKGVBMqj3+9FRVYqyl5g2Z8mgYgkdwGQadt/pge+mnQd3q/bW0W8oJj6eg6TJY
tlI3r9aU94F0047L02FdWrmjWGrxERWaMLBSutH4WEBaIO9lT5Fp/yvjh8+A7hEOLICKhUpEgoae
gHaZGWS44+9BC9+Y01VGYHkkldW3VAgCo6kaotVx6bl/Hz8d4L/wcEoFCR+jQF7QyIuuO/wY37E6
K7/ULjwCB2vS43Wo40qwfzs5ltIj1YkAYuh2g78VeUaLvvKB/v/zBklL5+zl6lvofMY40h2Ei4HH
593oDsXZ1MHTzxpTKjMixrDcnbeTUV0ZfmpdfU0trje8hda4PvUITlV2ITmYNW5pO0VBCWgsZslZ
kMWDRTF6PHbkHio5R/IcxPAoZGPd6Dv+wY3Hzdfv4hpHi1xuFcGrl2Vm/eLg1CqdEO7UEFTCy6Fz
J6pC4fsL0gwXcTREwLq8VGSd78kp+n1/y/hJeNd+Tiu66U+8fBgBSP3jTjbk6y6M59yxFph4qEZ+
Ay+bnKCboS/hmq61KFg9XDga30KIp2sPcvHHNafHWYVdol9FYtRI6aw6ruN1dr5M5bGCbOK0z8Km
A55c8CI65kibzk/gpVL1C51tqLSsLjJddtcjGRsrYSXSpu98m9O7o3Qg5JAt0z2jrQhIf9+xZwAA
fRncb7U/39K1u677Ghf1HjLIwY0iTrIktegz7Jzmk0V5dsHN1JsTlWO7DYYPSM/bN1ANu9iv7sw+
KqfCYTd5G5rKKimgs0himAqT6WkQUqSPPNZ68X85Zsgns9Zo2xGwrSlZYS+9NNllX7EM1ORsGBr6
cjIDR4pRBW9pvtiCoKOX/Xd6ZgHxQJ1zlyaWo1DKkwslWm7eeAENTdE78mcD0qE4JmtspVMB8uZz
8CA2Za8r22ZI8qdHnZx90XoajA9qBWiSuwjhTvwoAEj/F5Zz4qtTwkOUbpgM0gvgHPfnILkJD4Ws
CxcHF/x90Kh01F+VlJLEAAtgLJ25ETFfF1KeTmgFa0wutcKVi8TKp4rsKHwM+cV9bL9S136xolEg
fIWjTih4k1smVOy+nBci2nwRXdxiksj1xOdr6152FqxbT/0l+QCSjczTKtjfF73XoHryEFzIjmkx
ustSWd2oOV/M0Fe0MJ7GWHf/e/aG9ttetUsoYw/ixNaP62DR+urVFupNYJhM4Q4mT6TrdDRNmy8L
JQxAPfxXl4eN+sDFdrsp+mR3q9FwcqvPen9KcLNpLojXX8hSoyvxzGalBK+hx+nxkvgu4n6L0MvX
5MN3S9iq8RJ/Fsdi2NXYyaSCvFmoZR2FeJBnVtMBw+29/EBMoAiq4t78mhue9bnj5AiV36/PiJin
rPuFwBjdAO0miR9KAb9Iru2KGYuHsP0fyBaDL2J0tVIV1IR4mnlwfJWgfoaGnYiGTvpUajCBHDfr
VzfT2qzf2jsFYa6fFd+hakJi+FGFvvmenDc6/kJ2d4pgpTtEKwn/sdxjKdy/QhbtIZ//rMCr2oDR
yKWodJ70G3CZN00cv4W/xMtRRYjRMYQ98E51Zq9zLfL35IxI3lSeFrwa98GTGp0nRrRVpgcLEQcr
rjR7ld+V2O01XyxSJUzVrWW4ZguWi3WUaBZzn07zdfjUAQCShXLazW2HaFVm5AwV3yS7rGA0GtAy
OGuWMVAyulOjnUbJbNEHy1vuz36FS7xdczWXpsVBpeOevjBjDKcJRkukY3YXYXTRiUbvSir4IygI
GN9UDLgSYoryIpr1DWEoQ2tUr6oKoCFf+bhZUFkpFqioYlLO4mdpg2kX3FlAerQew06v1CmAaZRH
SKQIPunzX0ohGJTEJQ+ZWmlDX1LbxbW4DDLHaF/KDItis/RS/UyL4P0pKdetvhL63LS5J3GpnKLk
TSEoDH2muVCeohpGIPn6Aar4Iz7noXidhbJJtsJEFCJG/utpNrWl1MMvAJdtgJnasiY1FozAA34H
uc0dOa70tZrMsBVKygPI4eIy9Q0Cy6fYSv47XKDnAAdXXHW4pbuAwZiXlAR38rhHFvidnS2q/lAX
3TrMz+T3BT9Ki4eJcSINQybIYwsXcB90MwIqAk18xdlzSiohezt12wZxkLwfVyc3xYmMN3Df4b18
6dW+Qu0mPXHxn6zPrzVzp3dbtDMfzahsogJiphu7KtyURDoZpneivt1CymBEEpeftHfOyqx7ydws
N6jXWXlmRj4/lZ8XaklG9YE/KAjSbkehwlgC+RfZouCtcwWKmQTcOeTQLYrHbjZKe5dvVD/DlZke
sPTBxqidEQv0rEzVY6Rwq8ZLn50UXk5hzv1yb06IOmeHVDGeAXVxs2L0n8kdye3bNkm52nVUsDSD
t6ruNu1AldpZB7pu8eN5ZnBQkpmBhZWddeWFWGXFrIT34u8fLeIC49K4n3T8WuxBcQNtwmL+KrOS
qgmkTZH+qlrnyL096+Z30TerXfk6q+h/ggraxfRxAbhgTo2oc4W+jGpo0WRUgFplkGqTAVmaGVPG
8ukYFzClONFd14LN/HQnoLbu7VkciN/jYn+juce2VZ8G/SPaFUiRQ/2nPYNl7GKFxsAGB0BkfhTT
9tI1p9qzAfzFLK2rKztoNs81mFhQmVO3boTc569aOkz7exoX/FJ93RtszZ99xfL4YPONuEl7RGQY
x3GaYK+5d6rIgb6WzZlfmznSDT4aA8CFJE7J9T/A1xmBkWrsHvvB1Fxq5icbLoUPxxfaZuc0/qX+
thmVo2UQL9G0iHrfxVFS+xEfDbO63pnTC7T+cIGMn1ECWsCJhIMybBYOlw175zc2xbSMxEpZekgs
gV+lrIRpRN1D4lwvxTMo5bGQVC6+R5NFdy/bwJfpTO+pXMA+BtQlyeJ7kQwtUtFJ231pzYiKGZmW
eO97ZrOysEVDjvqwMTS2CD84bc1lKrVAayvKAfjz/iw9xNr1Hc4fY8JVRgDkB/0kDHSMAs3o9mcN
AhFBiPrieJd+LWdtFS8bbz48YC5XKbUeZXmlQxvwi2+g4Mg7/xbs9Azq5sIQKrbEaiuq5MwfoiL5
1aKtBoR8DBa2Jfp5+c9LG0DE5CoIoFVndatKa0EaEgmlmqiCZafKtNQ7EicQSLXOnVa8memjPsoC
NBFfLY6FtGdL+AFYKCcFG2yYfSRq9Wi8L1Lvcc0Yoi2oL56ArlZxlxtZT+z3HGX9B/Q0MA5TB8/d
1Wa/Wa3r6vJxzNEkduu+IQtchMEFoo/DxK/7HmUrdFW+twPCeQNU/6v2Z+2iEWTHNNdeRgNDu+gi
pV5tfHVAyIq6JhDlKK/MaZGz7TihdiB2nanYEr3QTFAam+qwgW3GLRR1HA8Pu+VDJhF8R1/42XKG
l4XbgeKN+3fkFdfv6T7hJpJJq1i5TZUEsMBkAwCVHZgWMI/ySSeDYG7VB90Ly38bofnmkdsQs2UZ
D+DkCvIaokx68S6aFXoN6alhWyY2wrfUNXtJeJMeOKe1fRQ1/ggPZh5up6McZg00vMJuTPKtOL2w
BcwIw13fxKjJPE4+zJM8XN/kd74hVtIwyiQZy1zggadS5z3ilOXXFbtuB69xYiXiasJtSGMxX1ge
o2sCIg6Dz5V77YVyHvTd4YSuPU8c4pX5pbhSEcJ2ThRg6ddQOTYFgvc7yxcC7+eXrTaxUuqvX/As
fxe1Zaz/3my7/RP6En1gDWQfOFHD/yUsRnILqYRLZC1G8K7NsKdZm/CqPoO+UMdqCHsotgqy/dSX
G2xYvVdAYZVE6GtRBzvR6nXkJv/R+ZAjjtH/fX5vVhf+ZVks/8//AubDUGpBmF8u9JrHcsUR1olH
QbaTGtoOnQsvXwCR+OzQdK+1+BVMPbzlziMsa5IhMXLQh6saWm7flZ+sw/wilK8gmnw/4rsu0+gV
AdNmheEIbOz70ZYEp9Mc+DarUhw9J9f57ofvkv6dl4qojv1eiQyP+wZRgGV7K3azB6hU1uqNLKHD
YNV89Fei8j2z9qs97D93M+sJScWmKmoI8nL7o2uCM00ZXmgwv4W9CuvPTMmTmDxHoeL5zmsqhwhS
bsu/pGM/BzQwrSVCX1Ne0K+HlNxAJeDO8/oDgLNKjBZZJ4tEvcPJlZpR0ZKKWXa5qmuHjmR1CmXU
syh8uEE2rJdU+jJKBmgQFeD0Rd1NBoE5dqefKn5KrDeI0V/Lc1/ZqAk6yvZI+gbaV/olUwWDJ2fx
aw92O4MGOUqfa3rtFfIxcCP7L0Ut7HONkJ57/jzC7xK0pfkuMaoqLft1W9DREnoNXBkfWypN8UBi
JOazV/w8gydWSWNVbrs+jQ0zWXdAbIr4hu5IOVY4VZK7jilxIuMIiZf8Mq5eMADGN04eae/Mql3H
xNTT6LHc69U6+pVS9P2L0gHlaayQLOu7fVr3hXtbUa8hi8DnbbIc+mzLGt/binoGZ4BeCXaxJgKt
OjuI3x/soGOor3Mpg6K2fhDaGZ0bNNdGFpU1Z+y4mOujI3tRRqQm9R+Cg/0zg31+7Fp96gU/N6jc
Hz9Feq6rfEz694AG0+tEMIgAqugcz7roTCe7dEdaYQEWEfMbdQ2qa9V/MeO878XsH0Y0G2wPJRnO
/MZbE7fueN9DdA9OEnNi7GC3L6se0AxI5jO2+lfEdK0zyL8wu29RV7cptb4XaRkJ8xgLMCUS5Qlt
fHBwt6Zx9yYm4ahjXo7XMPVUJm1YdTJcNlqQqJrroKjEKpxuYFFvJIRHfvn8Mcnv3OOnfgmj1u2B
sJydDQLyJ7/F18eztUilPeU02/1KyWSvvvaY15V1AHLHt+2tfbvUSXg2I/yqT5n9x2mNUcSY+ZCn
6RTzUNHImhZONBLmI8NF1UG/BYz4Qgcb995DPGgb7kUfIKa5ng4NbbY1Ih8Q4AISMD/vpVSv5zW4
KzCSX/yk0CTv8d94gLlxOAfG0vEf9Nvm7MbfpX5q373hf4vp1zxNYd86UsVK1c+P7rQWZADk5APy
wPXgV3ng3DCXl5jFXDlgSViW3TjlNW5Kf2BxuNSK/zMtTM5hfe7cpOziU3cdkVWRuMuzNjis64C5
g04eaL/e8RuYdE/f6CcYM0Nh7oxo3ITwXODE+94mjT2KvLpPiJV92kLroJYV1SjmEpSXJE80fOl7
wLx5oX6AgNdER898SjxMffgawKe8pJUnZqKp1SZM7dyThO3zU6Qun1LoGha8dwZVDnUsYcj4Nh0A
c3ol/IGp80z5aWAe6kJkepwOFAR56EwWWCl5/lyMc7YGK3PIuroSU/kKYS9ip/lfet7zVKwbFVLl
UjerQYCBonwy9oHf1pe+Yf3NNyeIQcqK35Cgo3tt8P+/ZwEFrWb/ATjZrP+W6onA4SX+tjmDHFp5
Ao9OKd7MfMJx0vJYFruHSVSpsGVy7eQ+qNHXYab3KCM3XW06OuerOnJ7JUGADHALg1Zc2RXLr3O1
B54Rwu0xCnn5K3sroVCD6sJCWKwIIDOb5KqrCZaZZx7jMgGjRpWIKOQFaZk2MB5/ljt02N16nHS5
kxTOpUIzb6rmi1rQoQA10czFmgErc8Tln8MnDdPI31x3u729oX2u8qjetbzzqrwdFOyNX54VmqR8
9WyL5bdbQDxrMgeq+FOXhDaXawN51SekEK7Khm8/0gKlWLALzzG2HoIyrRIsNtSN8m0mR6NAI0pH
apyRlbo0GXL4j/hfhTwt6vPk+lXGX2kxFiIL+pUk31qLl0wDXUXtzHbOoLRtap485PO3eSyj4i7Q
M4h4hprlLL6hGUGZjyYTJ9J957cvVYe4YszWmvl8K8HjpoRiern9NG+aFytkkbx1pqBATx8ZlqLV
iw2QxwLt1wKODVSMz12BfDoW6aUC+oc4OSOsgojUCOORSZjhg4rWszn0NargIJo7laIabCxxjjVr
A9AgEQC8Oo8YsRBhIw2ik2uoHOQLA9vS3htG9RSg9GwotbPA9bQyILIx5JOyTyOBIV2U8ywKhob6
0M5OXBEnZYvn3vzheiLEMG7W/tf4N4Wr5qdvzqe4o8KoVZbUlyfLeKX6f+AeiRiXeG/uQhtiKDrR
skHzofy7MyMOaCZBJXHrLlwfMrOCUv9Rl7JqDOH3ILBYs5U4fjB1lY0WWREerL40G2F17lHbcOXm
G6x4J1l/GUssQsKNBFhrHW4jAFUC0uAAJW5ev8NuGFLs4XCobs3f/drBNGadPUgFO/c/J5S+AHT4
zDjTxeG4EOWLdopGjitBVw8EAlr2QNRoDO+SPQDR7Gf+OeB+hQPsLSZuJOkl8LuuHZcY7Ta2WNOt
Z9XbLMJFBsZqtsBNbmdlIwHdD2DN3u9L/gZDsGly7Q/SEO58+1v/dzt15sMnMEAW5aSHaNHRyADt
v0fnCzw1DDaeuj9/ot5SCmskCT6uw/MnWqUFDuosKXU/cwTbI4XxAMIyQw6P869e89VbcZmOViJS
csyaypNzQ0YgVoVh0RoYPsbXrhTuU8z7v03nabQPWd2kToah2Y+q4huFkCDf9Hceb4pEnAjR71Nh
Us3yRm0WEahiSfjoOG9ZTx2EVdcE9v7+QF9LYvzfAfkMJz2BF7bukCdwcRvVpGG78Od9bDJCXakK
WHkRsWzJmLVf5CBYwpB7SVe3phfeMAOEFSypfqv9fKv/3Z9mghbDClZglDuEqnWiBCsYgqDgBl5w
2NG0YxUGzKHKRDj1GWylkdkI1J+x6FuDHkKFmM+PUj4DMau+kXM89svPsXVa9u8k9zn6QNqriS1b
F7LKwTIBa3WMkUSGrliHFVwQA+cT186FStbAs9VxhMGgd653sazyV/W1wGk3dJ6KO5qkQuZ9OC+U
PgBS9S6kXC39bOTnaE3cRj5tYp29xEAATxGNZ/yK5WzqlcjWnEWbVsMauoogSrBXWoafIl8138Qg
WwGwhBL6J8W87P35gy1zYt2bHxrHquE97s12xBqxB7wGX+qNSY9csdG0m1C7qwgbtWlq5chIw0Go
fYqnOocRPgFxTqX/Bgb/d88KnqoTU/TrZvadzlEby2ijlpUbtr8QTWIdNGGeakuOzAF4TjHItrwB
EXcYc2UgBJJXRCvgVH/znIAuijK+B4Ogb+WWCb9eY1xdQt5YuQs5yrDTg2323QQ1jF+ykWkIHm1G
f3tnDRQFSDJsXmOvA7M4F0b1PYrG9jSS3USICwKEFfkLbtxA8IH/1pNhSsOPygei/Tdhfno7wyVN
u1uPcqDkA/cSlQYHWPOlc5ToplR06S7Z7wAVYsdbD0UejH+Ioe+7GjWbBhcpsy9Lg67W0qERLj9W
sISUTYfsaLlAJuvbcT545sUofxbozjrsnhn4CWzZTJK3Qw/6+njEZsBYKVnJFPqlwbK/oHrvsrKV
pzD3yuI8lycFBTMQIEqBcpnhpx5lwtHoraBpHknclDjzGHkZ3haSdyB6bkjsfMWC9EVayN8qw3r7
Z2rJIP3K6WSQma9f0LRzblthoYh3D+rNzKAa+1ff+lMeMzyWqvxKrvPU5Cnm6Xu4I1UtXbQya5ky
MyZVrE+1dw7FdvDFnXZgFoXO/+wr9JTQNcp8lwsMq5XnqIqXUaT7WCDivCGVjjjS8xqNUIRELzGk
Heyp2OP/hU2auiD9hiV1qhrmsroejVVYEEX0f5fsXCaD+e12rpdECd1vWyNY1g8Vr40+Yaovf0VJ
BeQ892ilinGPEzam+v3VQsqtNMyhSb8jVu5j4zqKRWzumrZurvz4tfl/ERkzfgVsABgf+Qt1g+rZ
j50J3vDzfPtY1vDIbNf3vpIkskquR/7Atl2G/vreWhj5kdjENgwsZGjcPpzk4J9kk5RNtn3Mk9cR
3LHd2/1HWfu+ytE65Pp/mI2KEkdskNNbPk8xMnrVNIkNxhBVV08PJcxl4hPhgA3k03KQBm+CDBJK
5f6RXa1+/caLywtROL7ltzJRGLxfFVHJqq6HNw/Gy+IkXJYfKtUR7XkKwcUL6n810dEKXs4r1tFR
8qlC2QDsrdiui4uVTERehDCd70OpBxe0vmhONBpj8HYjFY8Pn6cSqNu4xHsJNtoVJAGRPSZDGc4Z
03PVy/8W6UtlyXqNSWfafZH71rQsW21Vkog/rYsJh9avO/WOArgcgECOiBrt3S1QzEnv7qOHSAOI
kv+ed1CJNlWQ6el6+uw28xE+Wb3n9JAsOAPKnIXFQHcITzFJ7++8dYxVFxGQUHxWIeUkXMV+8uaa
oxz+IUNikqKYefhNSmoh6dw28/9Q+cRsFWA7FZO5QJIk8c8bK7ZSMJUhcigb9cvttkE7mEn+4Slt
jNcqspMfbDPyueKZ1MH6hK6GJaCMNBthdsoQJ29uqbvxMWNu9lFJjxU8OnkWT0PHn5ZH6rNzdLyj
I3586KxwxAgY2e/+UrcEuJlnoh1rJL1kYHaT1aqF1ruz+L6gLdtPsm/rm0728vdsHjSd+807Hc3t
UJkyShyjnmWEr8+NWRA8NbQN8jr8w0MHl+gQoszBJg8jRLgXxk6f2Omx/YG+1IUOC3bm61ONVFst
pahbZqKRmnuslE4rW2pR7QznoAZzvs3SrKVdHYqoRLQS8EiVNRUIOwOXxIWcSYEwpPsb7kt2iSmw
HHetkes2xdS+B/WEGlUoElGtf/opxCTfJRHOETZGKqqd/6WeuC5EXNRwkCs9aBViIldwkG0Lvrad
avwIcXZPNlyIFz5ANJoTavEuYGsjVbMFSrt7DjTtiFYQFkFXrQZnb8yUnvBH2MrK13Rh7B5tAYkn
iQyOfun6T1SIfofJNUM49WMZ/KNrdfALAfzk4/aF8ZZ2uFip5g0uXNMxxj0Ji+W/exAV24fVugvG
UQlhJhnzriJDW4GbpQS5AxJi9w455ApQAm/HHZvIszs1LPt2RXX4tLpNVPVoc78xapSi06m+DMUb
WTD8TMbGCF7XoEIV/gdICmrLn6rLphwtMiBR2+DXeBOsPfuw8m/QGdz03wRLpCwcFdadP+B3mC1t
Yfb2Q9zsKym5EQx3eKryr5C9ZRZGeKM4+UvwERIztFVNqvFtxs5lR1zF1rcw/gz98OEEFYJkgeZK
tAl8PqNncxDb6gYz2TodQqr8gF9930FbbF0Xj5e1ESHiFxedNaVf50qGPA42hqJ6lIzF40cE50qz
nAiaXPrL8Fzm+AqZjiwbCOCqXY9m/xx/+WIV+OCxwjmKZtm5rw+Nq6rxYeX/A+doG9OicRmCm3AI
RchPhLQz4oyZyleT/syDFuGuil+cTd83VHNwiwTHspb5BlTwnYOmCdiY1VhPFGwOjptpHmmFYert
/+cUPMzgUHFW0y8fqI9LFNOcOPl4xtBpOq3IuGfn57gWUNI+cGL+3qJVLxvKQGFvNQHWcXq61yPU
JURXvkPu7PQaF6arvJ+Qwa1+GFuiQiyLzTDuyJpMX5uLnn9i8K88auh3656cL/K5JzRffxrKdH+t
OrhQDK4qFA1PSHbQTHzPnbbJG7nFgcLGPqBWUTnaNrEXjzChiQ802CJTes/kdQHGNvf5qoKcXm1B
brwy9VYDHReoqGqMJc157/qniPq7fIAjl0/QRGnhRWsBdyVlv85jIRvLbwXpUwqpOvq0QljYOHY7
UsZrU1dXEK5MYkcpi30ymBc+Q07DvQx0OekfacPig2Cng7zJakrgAkYD0LWiG2G0wmkoxvWJODuH
oj7yvjyGmpbErvuH2dyNEIjnWJvGjPJ0/vkadzlwHAu9BK37uP/aXD/7u9+nRjmpDPa+UzhFtOhH
+vQJxbIyN6Err1I7oCn9jn+AbBXLT6v1zZBYV2FNq589i2YYiqFUUyAU94FdkkOpVaoTfYdkgswg
LYVVWp6bfuYpZKel8w+YXXB5IRYn3mFIiq8uE2NmtABw64AcJtcOabiWEe6Ryku0+0+y9X3k6X7/
sP6DVw9gefKdREe2qxZuJrxVzK6eqOii+Cbs0u80+2a+hKK9c/N7Ym3sZzj/9pyR2jh0Cq18tZfl
0zGEkhn7nW4ICs1Li1/wEASWTwyOHkhFcZAnl+2wwi5MMfEOcDKw2FgARUY/7R88nY3LuqVPen9+
ZpjvOYwiMtdJY2d65VxQfGtitSWyYTSymPGpbhe5eZh+qSUMJrKHcDC8GphERJMqU5j+yE1yYee/
VkASfvhfyD8DuD4jHiJj4a7EVXYJvsJAVHJNrmh80L3gYW8NpEVSqnFzqqzczwghSNXX6S8FsPKa
Vwysz78y0+gR/CDBSWq4ukUuPSSD/Olb9u8mY1EUchisbiA8crV8bCbJnWFrFgpu9JMoy25NzbBx
R3rEDItho/vSidattXcQ4D2fwVWrbhh9bHF0+WwqlFtSp8+goLSItUkzV1cPb5rKLXyjh5PEuMwb
yp4Ns2A/JIcUnSMRq6jgRqbghUIGsjGsIyyyktC+tVJTFBRmw1w8x6zXeRgbAnlyhj/DfShw4rZ0
wbRWXVRO5ptxPeNOpVofePl7LSXWdOu4c7MP50ji7uVJtDewzOTjMcTNnr3lsFgLnAPU4TJRmzZi
nJHxZSvJqq3d88NFnQ4B+USEzFZ7tPu1GLIvmgQ/h/oaOzkmidide53ujgQ0OK30AH0dYYWJaFsk
0FFBdZrmD6FSx2l9Qf39NzdFH1jkQO3LSrGy/tDD/RERHGji0oPfMPg5Vjdsw7ELMc++a2kHdVQh
U0MUbzDBQnVZBueURGCFFSIxIVFXIC24oTo93uLiHUhAwNnTZFs2zUfGbABpV9PBYfa03zxUlCJO
uM7xP5zBbvW85c1KncPGFBPsp5kD3+RtgF3tRLMmBnnKCOBNFjePA7wPgL/2/n1RmUxpoVy6cYW3
Vaxfser72SxCKi9Y2FcAthzKuknxAmybRWn6s9Jp7mb75d83JbKY39MUjmUO4klxlOoBoxoUSvol
a+LDDZc24oFvKXRXQqohEs7Y1OhD9eUXPZVA3cEcRAqFTLyAiovk24+hyVo3vIcM6iUuQ5agguuV
AbECH1iw2Pt4eqVcq/8vXMtUOBiC0I4zOhqZU6Y4zg1UdQkgOEne7l6KcOsaQkgqQjlnJSXO+yF5
ksQXBNmBbJzRvc5ls/XcXyipN/JXAK6XtLsISl0/OIELAJJk459O/Y2Mcf0JPswRQseoVfSgMKCA
UrOxvDOOpr1uH250zZeH5c4FQTL73KVRqbkL/5PpGtzn+kKb1U8NkZ4m0hnMf8N4SPX4WVUQeAF0
/DgpsxVctardWlhOwetGzMXn6EIULYFe2X6nShjGp3aDBo+l+l/8iPyijjGFz/iRMRM006p1dGnZ
5A/qwqkBWVyBMzOIzlVbUHpqvl3QOeP+2UcS9EBUGGD2/pFGK/uGZa76JMkwZI5rIHMe5pWwNs4K
aPBLKRut62b8zhSAxITef6kGme9ax52qEpkI8aIaJavF4fSkwNLa5RlWFkEnq3CUfQF1mbaLYOFR
gp2bDsz1OwcLH7OehE7ZDWo8Z6lGqFa/NzCZEWPN9Jx5dwxd5oJZWoPv8bsIHW8Vxl3A8/IT6eBB
uWruzaVG4x+rQlPGhkDsSmQpx8sqZGII2TJaHB8mi+39+8F+TfIAapo0g9eUKyoDX6PSzyxyESc7
dPviwtO9ixRUD5uwH4yXzSdjzV5faBAJgBPf2n8AEcl8w5ZeurridNNu8XbdAGx3CFAbEcN04D8L
M0mn6ZKQsD3WXJyKseszSfzRR9GNgnFwBffDmySRKIXim1KUTcwM/1HGfISfFWnm0r6kp1lqDtIn
oNdFZ2gSVqq3krMZLqYy7ZNXiSyLpwgMQCJ8UUbt3kvLi0+O8h+G7aJZ9qyMtx63PluzHPsKiJYQ
+/bCt/qhmPP624rY6Nw33PQrO5BdbqSz6UQJPss/tabcjozxOfmIKamw8QVqxGvVm0fTHI3bRv/i
h/XW69R+I3W/ir5NpmjOnLBXdVergWfDDqoLLLVWeiU3QMtEysGh1FEW3eEYyeFYDHIDIK9MPw4u
K2WUwSIkIl2Dv39UIgpPsSVgLdYPqmbK9TIyn5TLWnIH4eLHB9DVdSPvVDYxs8dX0oTUhJOsSda8
dB+6AD6kyXdUq8szgG+n56fNg0xQ/RncHMwjQNZDkBEVKRYN8GxJVddjssGZipKRm6rLjsuRlyWW
rUi6M0WmzAU04IZSEpX3ScQGkhtmsMbM5HxFVvxUyqULIQq8/Y6JF6Q2fn2cwEccShWmeMNxAOmM
JcGwogTdmj5+jJLdaMGme3GywKXjnV8aHIHeTqIxYKYbqzqbHwWhs+oo4ovJh378isWQ12EMkn5N
+tTX0PIb2jW+LrzbszWoLR8qrEgUcCZ/ruzyfeKFnYFliPxw0i6qGmcVlTolBpMMBVEzV0g3LSEZ
Rbj7nEAZ9nKPAYRbGOWeLWnz+0O7mc28oks9cxeeuELtDFM+a35snOj16MP43H9UrAC3n44MY5oC
6Uqh0xKF+X2HLVAL2zHYtLXymhGXfoWP4sebYGHz9j9W25L+O65L+zG/s7gWoQgAH5Ez0EApgiTt
QvBAJALSt+Z0maHm1479LRiDnEvizQoble+7Z67uWawvUAugLv6X/Keb4U4JlMOqe/tBPB5vZRo/
d+s9AR0d+xqd22uBTlFEDZcqLwP6FSrpivX9bleCyhOkM9KpyLFOVTTEBc+7Y28YGS9gAHpxwQcz
LG2HOZ2cuexpnk1ZZWy4IEYq5piFjOYXCFzCuXBvOo/eHVAiLe8jOSI1Aq3VJmohajjeTExDUxzx
FZXWr+UI5Mv5aZDDerWSKxcnxfSy58lvfZQO3QgM7HkG2ffjq0uHWQA8IiCG7msfj8oujaAwg6VU
UOTnZcngEuxPwqBOIT+zT6wDeMd933djblFeWVaG5tDRqi9x4enF9qeFjX23sEcZ9Z2MlONZQ5+v
Sfm+jJvp/wJWHLKIg5Vbc2TeBw6l0HyV9eqQFD2ohksrnU/D3QqiD24SzUTNhSVgw9RLRYdDrgBb
aBQbmyoSZ9qDuilpSJCtTGRYEY+zpRTe12ah47aULN9xxgjQC6ZTXSnidE9fsyxG78JvExcNEV6v
i1/nyoWq8SlfBJP+68TQ273zDM/kwXYX//W0z0waH1Zil7HdJ7Dqn3hn7nn3qcrLf4L0W8645YFy
B1lNHmfyzgjjtCow004aocz7ufvZq+KC4AowiLI9qpTSzxTD0NyTRihIvkcMfCLMxXINiW9pKrmW
6Se05cd3R6zpGmL8tsmDwB94PNoiqRSYHnGHxkwEP1uwL1rHRbJOsRkkwiVDTUOdrZbdpfk+GBiA
sh3zjfx/ZT11K1w6hSIq3DRqjQlE8+L5VHMbBPjujo1ZpWc9LEePI1B9F0SHLnCi3PQ4JqHKyEG5
oi7MJOPaYU6wceSE/pbCYxTH/kPIZ4G9S2JSmg4uCNRdMtOQz/cC0DSbw1618HweLDXLkVqvgydI
Ubn+FGVKBwK7ouIxhNhmL8UeaxWXHlNlFcfN7ewiDzqiB8OrhLU4HGhRVMmTtGwHCJHvg5C8alnV
7uTffcC+EIo7iKFzwL/YSrkDENaIOY3TQR1Pj6whpAYPvvMO3znDCQXHrmooCvIQzGRfg1sF9Yyq
6Uz1XTCKASBGlACXSUxMr1UifnaNkj40lk218O6q5VMZkHfcrpVTnf5pq7zprc3A7SzoJkNew5cu
MlPbAPrE8fa/FmTk9KmmZvyRfGNVXM+0olO3Mr68jXvj1sRCIX55XKuf7fh7HEbfi6TMzV8FZKQe
GiD+rN3gGHj7mAWtNBIJ9zcuZuBafho7MAQzA8WVpp1euqj7vsBVhIdTGlB1wxvvG+ZJ3JpFMOt4
aK3aClXpd8ccuz90YN5PNWPf2eJALvm6rlM76JaU3u2AqFCKPSyWKoceabZT5VlUFRx1oTf+Fzlw
zjsEKvOpoHP5RdmyShoZb0uJE0qaFzCVmTorHQ4qYcJkACITl/lsG7RaI1uaV91DpRtsQfhM3egv
nvfz/7KVOBDVarN7j84b/yCioZ7OAhmfuH52FrFW3znLWY/9lyNq5ww5WfV62UpShgOKmqDwhJh8
eQbmFxMdYgMW2eIy9OAaOqjWm1SKiEJa4iPT1EKtG3AXuUPo7xSHfGE2rRCYMCzz3KJOYl5ePnPj
DO3JRI/1jf0uWUmdcL9Red8xWonsD/23/B0JPt4/WiyZ9PFvznViF7C7YkqDGkep9irdN5VFuHPv
92fh21Nrl0C0vDDSvFDl12OsXha9fOCNNzby1AxMOrAo+9UM7DL/CTydIpfeBGyikG7DoKIwhWse
TSZe7z5v4XplLttIEcwKWPK2RATtFDl3id5ZMsdEEnIDyQHCgpVUJYwWg1DNSv+pjCTBFxZyQ73u
n/9R507VzQAiH6rWg14eqEi+gOo+LIAHr5ti/XYi/5yfgcbE8d6nHWPAfvXdjsBTEumVy7QHoiou
UKaLA4SB51NjTwimO8kNTkOOjBHbAwqbF4wP1h8y9oqLXwV9f1VRM0dooLifaopbUU4CfHriw31D
3xxzuf3FfRkba/7KtuW5CkT/8NklqxrPJsv95d+oczyRLjVprFnjGNCg5p3FUuqnlQ/dp/pGyvJe
dMLEkMroYU5/8DPkaGrC8yXvR01SJaGHr/N6OXOQpN1i7JBEQ+8hLDUhMTTCMp1J54nDuOwttND3
RgQY2qPE+XRwlkkRlgC/OyoDHrx0YWcRPX/0T6N/Y++iMwxmsi+Kye7Z0uSDUL4IrFYJPwvSqzFr
nCo58kg+zoBJnxKwYrMB6AD7sv2cPYvwambyTXbZEuG1UUTS1S0cfErsxS2Nuv0o/LthvG38dNEM
4RJwq0vuNr9zpM+HS54UTBHQGdtrwKE52YJJSyAIgRy4AHxkpkW0J80Sq+z80NhRzYuu16pRNSbB
Zrcskerp4qSYi3Xr/Iw9CA+uw2degSVSkKS6fZK4dx4ELHVwYCRYnw+G7uW9IQJRfdfceuh9CDZT
zjOkpa208QTBluGwNrbK9brJkdGv/f7jfEVUDOyabGipGIl1tFioTmAwq0BPimJlJWMtITXmOjR8
q+KHWG5M8UvbmxjaUjcV9Mbcs6ok7mngfz0za4tV+Z8hRg2fiApmQeeidzTqG567P6lMcBF6TugU
fnYkNZqO33lJCF4/Ie6gXfPTg4lOforieN3W4OQmjwC1FcCPm/6uFrX4FIWHmI5ZlsTUrfiE8wA3
Hep9RKHX656T9BZfeib2GDbc36ZYISyLcaNCLm2qx/hIIQj9s8GOBhupfD2B2ojinD7rOpQchi6N
CTzBn6JaUlDGMFlkkDLBZ4pLpYdnhUDy/I/kANxjy5TNZNoBUZdKpjOeVyRFeVqW/Nvj6CEIIW7r
Pt85k3fEhmdmHkzsAFy9d9tIbWlcqkM48+m+43OSwwB8f5Zo3mE93PDun4mpvxcODrdNVESPHvLN
5C/E4A4YUtimkDF7pr1UH4FprASvXaLZgVq7I2wKwNguFIQa9sAgXcsaBDQuBEjGZmkUA8rTwV3D
5QUdxbfHpyQ+LZFaJgsSj+rIQjDEe3tgrg9GlZqZJnz0qJ1vyTlxd38Xx6oiv/zPdWxN7RzLdKpl
VQNzKlLucTOnKhLMNbRsp6/MaNLsOx+nPIZzJfXMF6sLqGtfyPtkcU87JnES/hAhJBSx4Gzh7uB1
iWMbR6ltSNjW8xU5rsjH7+o6J2QfN8T7CN1Spu68lHuEL65yZo7R26aUA3EUBdm8g/NhTKvRUjni
BxC7oyZikagH9MQfzWOHo0adFWCvQ7k1cTWQukkvFHGSG1g1d8WEAaeiOpcylMi4HIy3Rla3bYjA
LrMPpn/2vY4er1BO7xMhsFBTHlgLi5OlpKvkCGzzNv/HQDmWjx/WYVoeQI6hp7CZHJtlQAP4UEGU
jXCh36nxSefhaPjDXEQRygT4jn5SkH5cWUt9QVT/F1iR+kNSO+8OQDf3tbGEGhPD123ldzae+jxL
TovLY1RqfQ9uFiXEggR5GZOpzx3I0R8A0Nb2uZwRY7+p4WjvVQSr9q7OG4u/gQl6a6xnITnro0am
1uvAXGyb8gsHbjBbXKUgv2zK72l1exJQMsjqCi+CPD6j0VzHZ6H2GoImOmwIN83XcK1zYHHnTCnK
BuqpdrPxaNKX3flVYgnzuZvSZ/sB0+mnyiS6RBps8oypRK1DPisaJbrbjH6s1+yhtTLI3XP6mWQO
T5smJyCQ1B3SgnuSsPwQSFzGZrh9lGWcx5IvonIYzFdwDAJ5LevMex68p+P3ZbReLFM5SVIA7grS
Zx0RiIIvRndMSvOZ0P59tOKSR7wRFzqT6eoHkI6okKv9bcXcTxBOb1kmyT43899Jots6JNc+iF69
6JYcYfqam69exwCzy4iYvuxp+TUysGsMvUguKhHrB8e2IQH4qps0GodfvT2ehXKOfBi/hsShnKMf
Fh/b+CFx35byH50QC/AtdU3jEkh5JC/OgcKKBL9PFg/9kT1hH+6sk2vTQKFxoQppFl19LdomFXka
uAtzqjQFS9PFsla1H+pWGKzNpukfRvEFfm0T2pqndjFNEEDrvse+ln++dEnQHw3qnAIbC4DHfA9B
vYQEpaXpxGNGrIQyrpQFI1IwGx8NH+MTOFMYLgySM5kANMmdkTvc3Apcy8naRGRrXnNJyfabl1Np
M2qRGH6FDmZX4UMiNTRofZcdSsZa00mC+ktFaFcZy2pJNXwac9ilg9aLeq8KDgz07GNBBvrjRV/m
pkpIRqtpQy25hgaGB9hYTJHccoRAHBR3sq/Yy/oO7aJ7srg9OZoLpFK1Lu2Tou56RglfMTshfOpb
OAlGzmq2glfPtL44AFHYNYWb0QLPq985fiixWegN9iq4zM2Fw/JVu2BeKRF9HDlHPeShTguOoGkX
MOGjAZ9D64nw5OjH1J3bJNmxkWN+UJfrBWS+TV278m4/gpqODWMK7FVh4XzHp5R8RfG9BW3yBtev
laxsGK97JjKCWJC8ATKRiE8txhXyEdNOUi8/sTaCH9K57FEQe6Xd/MZ1AmQU9eWlllTmlAHQz+hf
TNZmdM5N4/B6jZ79UdZ9JvH20GVvu+g1tOPXjYnFwsKTSz3dEbqkCifMT6bqARID9wkjFWrjtjoj
ba2QRvfxWOv0Ae9kfNUesephdYq7MRfyTe1C3vkhLwdf2kYDWJd320ZFSn+wUUDT3B2mL2Yok4L6
Q5G139RnUBUNRloMHlvsuo4xHmo35kT2SUfGmIotrTYNgivh6Ma1SQSbodqNB2DVWWP1QFKg/6uI
Xyt9DlubC2TxJz2RY9pUR6KmjEXwPzKDjDqgCny76el59RYXrco8Oz/WoY8YbKdPPx1+FxSwrqIz
gyhWMShx7OHTJTnmNNLuBL8vVE/v0XZ2mIRio/Ey+f8R/DtxbHTezrw/69yazrdbzCoqwQjPHAvA
yRRQ2IDl2hlmCcj/jUpY3IpqPJ+Mjv0clp/8nnw+9bHmYg0uVMGz2NzcLFsYPzVNn1iob5NgSFQR
WPo2iB4FX3aTXXfw7JBdi5qA72ayAJzDXaW905DQUbbpDirZGzuKLAx4RKX1bUTxpYptzyhgy3aA
/FPdJpJ+JgaU595JI1zUNMfDMfI8gyzq0CjdRKj1x0ZB1vcQ88WtXtG1sC7ONfb/HwbiTcSD8N06
yO8s4clV5Pyl1IAtGES/VTXE9EQozJLm7FfIhfymZGfHPBV095UqESxvOZMFtuxWGkCxAskvafn9
L+MRNoM+wY2O3Ib5NaXXB4qx3LshcNiGFgGpHMovYb1l+bCUv9mvoCRLxw+GFacyaiKo9KJswixI
IvGGhYiRMLFu2gHZu41pUr2WWKKLYtgbzBwVO3uNYdLm8C/9nIktZcodNleYGvi4hdgFsyVQNo7m
6cZAiH0bAlU78M00N7BxwlZzNKfj44R904SwoM9fsAl0klxNO8EXM4P51b3Dz17NaR+C9DMfGoVy
tYh+4tpUwFA25piPeNDUnJN1yiKz0HXBULcGdlPiB0Bwkx7zkhK3gBYOrQdIQAyHJLDVAB/wtERE
fqiNz0r+58wLWnlgUsvUXTCdV+hYiWrTCY9t/Z3PrZSXtVpN2zoWkG57wraxBLYG9xciatHzHiPf
m47l6eN8pwwj82zHap6KrXaOoKIPgeqdpqoQxZ/2XxEZiZT5H1f6iocWZdcC9fzlhNeNU6rLpFy8
z5rnZxdEE5hh+JrAKBNhBg0ESMn6dIFg/zfsh608mB78qo+ejkVeyeTlAJ894EBvUdk5g3wOXH3q
0/R0qTTxWtUQrFJKwETg6U3heVGr0YdsTTIAT5Xs8WfE1k2egeJBl4N856DLb7nKAwvBFZNmGBTP
QZuACLBFHzYn2EXdSv3bBf+oKZM3nLA7iGIKXNNhNkN3Fd9WTUBdWRTvVpArW3g+uX8bxMW7NYU9
wN/kw8nR1ohjLNBaU3uxSj57PEPfAJlQS+bMDmN9bJ/beZeXFi3P4/TLPD37c8A1cPdAr5p7M7zp
fFCLRnf91W9sPR7aFMwiLA2dvOkMhN/fQnYYDWAZBK58jexJCaodTEy3GnY8QOnOp7CSf+UyAXZH
N6bSox5edLf2LbRLUeZaB1zNdL4b1X9BFbSviYn0L6v4eK1xjxpGSp1FyXv37XS7gSQUDlUS+LfY
jKaEctgURp8JwYPiPmUM/UEzxwLciJ4F7LWWGesVl+oMdvEzTa9QzyTzcYGb5wUjwOjSM/iXAeQk
05egJYzxwwTC0Paa1Xujh1aCJMg20AvX+DKbd2/C7bK04djCapp8uxoi91OhImq/UQlFwx1aE22I
vuqO+6YZk5SIs58ijyrOUU/7dT1IIj5mqM+aewXqpXbMtbhxRJ7/yS24KnXYZCwaN/L+p7pPqCpS
z+ECr+OpgiOxDh+LWA2D0hlFjAi+8bYN30VHeIr8H07Kdf/Lvgif0f9CjUs/VHc0FJXMeB2rqe5p
pjr9nEuejzVrtAIsdFYmRrL3+NDfHxDDNN1LFQwLDN4grgi+ooVKD0BP1VY0vcCH8RFAxT343UzP
NHjqLPj2et+ZLaQOFRrw9V5Pu3Gmf7a73qutL9KOUzpzN8YrrX3MInNC9pcqwcpWnI/NQAiycG9p
B1/EKkzlG2xcJjuJ2XcyQziTFRlDcMkDjS5/g5AflinYIWJIwCe/y/cB6FM3HeuSUn5Ky0IVRz/H
7nW04PAWm6RzPMdu9CjiF5imaAqUFga6UN2r9O3cRvb3jap6lQDyYJnH9j9ePsy0lpLRjsRoF6Kf
UwCtPmG4yUQGJJGM4tVJzm7tn/7bVKXT6P42mcmqyg1JPzysnb12j69GRTuE3mOCvDGlaKVEvDJL
AWzKpc7nAMcK+JCtWvP+cjlf+ps5HPBguUQ+RUF+dnekN+v+RkEuVZ5yUobxCd9FBZ3R934ShW+W
ePAHYiRxnj3Q8n6K9IWOkGbOBuL8ALt0CGs/cWqEufFdV0if0ZY+lgKpSG6JrmP3bEShwUQiBDGZ
ogJJDuUJeQJ1EX86VfwmxShtsgbWGlpKjKU5sjCuTH63bEdqFOWhDQhZRN2OOB7BhsNF/pPS3mv7
z1avb1bUcBVr150awxzaU1XyY+kmYh2VtFQt/VyU941Ji1LiaTQs3aNIDv3BF+UyHCWVnPpMpd/F
LKqkfBElkAyzrAhTO68dKAGPHbuzT9/DLLQAA9YpBPr5b/rEd7nAcJIS02QH8MR+SKNiQQsWegSt
e/uAfRanv6tnBiRRJ8P6w8WEqwiLhJjGxq4eSzy9uL1Wi6rujmKe0xD7bRAM6I4i+RmA5Z5ZJ0AA
oEeUDWqY38OyGdVY3UQGVkTMEns8hrCXXFzr32JpDftf6F26lUwC7r2K1546xWga0KoFG05niM7n
ficzvJV8nAPdjB+QB+ktx9VtKo9SEztLAv7etOb71Jj7bxFG3GOY1rooKB1MX8ydpWpEGQf3rZhq
zaZQk6cmzx6OpszksXYGGtjR34QOhgN+91fgG9NKLedvRPv92vezJAFu8iXx1VHzLv0zXP0f3e/b
WKCDGob+aKtz2ik5HRGxxJqCOJIsmlCVXRHZjBuECmXyGOavC+0e21xBGMePKYLlLA0M9TKRAvOc
vV8WUygDjMigTck1S+RS1yQkpR9owdbU7qR+dhagNsKWKnbRHphYGqi5JmwJXKqXuzO/giHf8heY
sLaG2Fo21UKoxh4l+MXPwfbYrJ7QJI1C1zEYEAGz8QcBoXq/Fbk8s1dUPQMs58p3dqvjw708Ymww
d5OlTGO5kxsOU/R4OPUlWRn0QypwUGJQn0SaW/U4f3dwAW7zsyFX2PGLXRmZ/TftPFL5jxrmmMUT
q1sxChN7drhWqD80f22NKdYvwi21EHPeuO5F8vgKjjmVWf6l7B4SPuinq4IrepQJfaXw69D9r27x
kggA08AsVB2C3lVWhcO9rNW4yQwMU6FZOgsvNBnLniBZaiJicIhTk0Sk02JozhZE0LFR/G4CtoFu
el9COy297Mh8RxX79kla0DOGEgf4Un5yMnK4BbMRphD/BBhmG6IbGfQSquQNO2RR/9W/eqxGbv70
ve2GgwjnrAqAyYAfhr3OMdvPz+pRZZIFMym0X3W+YzTBdyU0s7MjaR4BXUadnUxK+3X2YORTg4/7
FkmLXr4l1Xf/cUdwv+Q4Mj5OSuRMSjBi6Cq/srwRRugApvZ3Rw/qLKwA1u5Q5gdsKZOc8K6konQc
hAQj5tS16mbdoamBZAZ4h8Uh53huC5GudIZE2PrIepXd2uzHlkpt+OXNoy6V/l7xnmcXPuc1KYm8
2HXNyI0YhNraWNzVp7eHBmFxoi8x4GtUTnkwMd2rfh7xX3EFHOEkWPQlP1eVYIcLrEWRngfj52kM
dAe1YoC5tVRgb0j7dJsDJhTgP+R9gjnUWekXGrtnf59e3xdJmCThQhwQgjXCwCFuWaNs+msJEwnb
ZF5icgaHKnGxfQH2kjxoYWUeii30X1EwtgI9/Eob/M5ULrlgQn47mscHvvd78ObCZqxiWUyXN5oE
As/QsT6H7WLc7drstrJmO6b0EehX0Doy+6v5TbxtgbmNVPlPw3f8nXiy/S7eHrV68vTHSRJ0ahI0
jeLJJ2ndhS/GLmkvuWMmVt0JeZ3Pi7sR7B742JhfA2x1No6GvltD3AjQRbTyEhHWcRiZhIVBe0QY
ZVJqF/eDlPpXmB2mnw5ndR5FXV8zIKOmzzZuCuHt091G+U8qOB9MjwYn6Z9DURMwRAptxdNL6Tdi
dJ1pW2EoVblgg2I9KLIG+hxwFw7DnIeS8nCPQDFPiDTMAXArbYSQ9tFL1D02yB6tKjc2gP1kS+X1
R6G/aeR5gZm/DDtJ9DURL9wkZrn8dFSWlEZtIxSk3NJCMyd4Cu8s1wcDrmHUHlTOPib9gtwiVOHW
hCo3KnHclBYjE10gYvSa9zpM2FEeEa7GPgNtFwavODTThI4SIMGgEN82t6XypRByrXE/JPkalnze
pE0rubMACXUDiFl6d9LbRZQSHWVGzaYjn7zQXeqa0bGRBh8M2Zsi91GBegymmNZwCN03jHuppord
IVJGoD67eJwIvfcB83ebzhtcRiGqMKLxzO5BzqOivmT4ILBK3T3GMJzHBjPJWp/3eWzvEF4UVCC7
T3QaG6/OtS1VSTPnDWWIXB2q66gwCKrtofi9zZ295S+HkE4jQQbEvQ4esEAWSFv1YzaOjFeEC7G3
Wag8fwxnEWEPBzlBJ4WLsccXchzLZuiLih7VXiiA7kpJmMWM5P3R9hPGMq6cpqTxH3D6oWa8Aghy
7ymLXBqJQlSKBBR6d4tV0rcKHvp0hwsztPtgayKl0wamYymxcu8RxiE8Uf6xyOJrdaBUJo4jVFbP
whnhWkozuGg1hLK6mkC2FK+IVEntn4nBpJQ+CPlBjnhjjFPEA31xRIEOCF4V4MvGErDkyNl7c4wa
+jXejsZGmw703B0eqQLVdP8SNbec/RLVrb/DBspCdWDXinRq8vBSrxgtSfMWTSWbdoWBCUqD8Mcw
zuUaxSo7smv6XD8X4Pf+RovtmXa9locUkAmi/ITut3Wx7VTnp1+FvH/mATXquwOZXnob9k6JouzI
6SRg6YNWtNv5GHpwazLC5TKirYKalLjhhSgAwgBc9n6kH5XEX8nCl0bAA7U+zoqypBSC2CptA5no
93uJY0QeVDy5VmWli11UBYJF/BgiFxQDSCreQdD/BwA3oV+U7/DyuVDzUI6c1u3zljp8B9Wg1wJm
CgjQjdouss3aAQ9iPqrk9PYmXKIWB8ELjgTmZI2ZcAaOGInmbKmnerH9GwDfKSDjTatOE5dugFS4
hH+tZckNvzNdNZC8StvoV2W9ba1PBEz3rAfPlzPsdbVXBc5VfYol/j7fOd6ZT+eGsC1bEbKSEgio
3475Y0AP++nF/dKZNs8FbFP9DBIVgt5JxOTw8dopkB3SMEVZ48MhkotjxXR5eaBGuZGvCHYSWKZ4
KQmJNR5VcuYu3/bYUFTPT/SQE2BUFVs/A0Go2w+nJvG5fsw9y+Qfq0Ku5ZieVFAmmp7q6aV0IpaV
1HQpxOeUuPCbemNB+FRgD273twuTwuo6TlQ6es+kNdmZz1CLlCvtzsC5UW6wgc2RDHs1Mit6U+yR
rBsEvhI3g6hC5C0ykvQeJtj+QvEuYwodqknmW+lfsrfCIS5jJcOZ49sqtMd5LwxV+MDFvHcp/Ouw
MiIEB2WERRcyZg62yKTK36Cme1M3TV4mFssvKjcTyqk9jwK+lCwLf0GfakNSUHx6zkdugT8Su90l
NedmDDqZTNRUwdldznRciNTuddEYheSRIQFIZ0x0q6rBtFs2Wsk/2Hl0T4rQoKpeynsBJN/fLQ40
6Dj4uHKGfvUn0fGRCwwO+o3R/cNsjUE4Snf8QE+9yq8BI2dJ5uY5gqwpErUDFpDoSOCgYrNlyf+1
ZbrUmc7dhpQJLeA1o3hWuLNtTtguvGOR0nZhC5QU3FOlnHjt8Jlg+/BsjjZBG3TidvptsFVzuUXK
6qHrM+vDZeclrdncVLR9vp/G0xmNMWRin1fv8k6jf6zr5lEDbkKoaXEKHo/ZGZgtsRLGTnQqoT7A
5yoJnWAx+gFwm1hYJ2Uhtf5/MY+YGXHDlzeT2SFtzUpzheemdYmg4EsDLhPnyNGnXAa71Z+gfxad
V+KaOA4+l0kEUj4xIRoGluEeYFotLCdVzuPDvCtxI1/5z99ir62LnLvHO3CJzZnpMMzoDwN1mG5b
or0qDqn9KfAs4kdFTCETwwN6zktI1zc2jD91YSwr1G757VCgZzwX/+5swGE18+J41NxPcSEBME6W
OV4XDAjMZSQCwXA2/OwVEnd5X3fh6vRvUqfi7NFZ1DxmrByfhMxrZfklVk9v8b2RoZqyYsdDr7e1
Bs6ce3g3QD4wSeaOwsEb0agJB2VW7Nli5UBsG2Wb7bmWf8Wg+c25Mc0t+6JigbokWlDas4duMjvd
YCbtD5kGEmvg/u1L0uCU5smOaikAKdy2oZ+BTVCvZmqPiuZCLN1VzmbAU8VFHLVLJPRfXAj20cZU
abl1eW+dZtwvZMfYM8Luoub92dm3GdSSLwr5aUKQPcE4e11iA+FYHzJ+sye1BJW/DPxiC0/nH2JZ
gViGp9BqI7WeukON7WqPYnhOUkJZyPyir8XAFvJayV6o4sIs8KImzf7w70s1+uyqbRxrVL4Oypho
bHaawUciKdGIsqqP3cktxjMJQTcOJ9WIXO2OP/fGywrP8dQIe2oNznYW9Ysh09PtgwLpA/t4nrVA
gzKdL26lMWbsXbGD4/OW1GS5D6qBg0lTjiy7SM3fv5LlFyi8ca93SuBfpeL1jpeWGgiaW1gzvMuG
Owk2Mhun8ed/Xbnbx8tAsCbPcs2CuhqM6OeZIPMJr1XBHnRCoXa/QDldID6YCtHVVmg07krozE9H
xa60ABiV8H3VtJ3YXxHRTPtU9eJcHeCw0/bwKsIVvLgwOWk/vWZzPHNbW064PIa53aL35aiMdxJo
849VrhVNnju0uOkIHGLVJK10wv0u08a0ZxN9ufI6QaP2CJHwSowoxSHLPkNqstyjPZBReIPRZn8w
zV66nFdZMRHo2pMWRB81Fc04dwyCKz04l08Pf53upigqIX9tb7Ndy4FGC2vApDYyCu5Uv4ZwVm0E
gqgBKAgOlELjMRl74bevUgwxR3IC7kyDyf3SruO2hyb9MllAxLdTO4gQdU36TAcPI9ZdAXR31pIX
YNjN5CpzBH7XGSbF6ClnNDx+xI+c7CpnGE8LgY+ZBzFCInpScc1sGMm/dJxB8eX9dzQOoJkJvJU1
9bUownGJRhtvdQqqzk5XpmXHIbv0j6BHLkJ7SQxayzG3QUF2wlXO8DALteRrJFYGiO2dJ1TpCtFW
QbMin6AN5tAQYzVWHK91urarhCp07wgEoD27f5/+eybmEuETEh+3iqE/FiWe8zkbQTlQ+uVymtcD
SNiaUL0ex0W0TBUVuyVjIF0PqqefZsAM4Gl9bQM1Dshl8ccMQv+i/Gx2V98QXQ1UhRhIjXaIlNkM
UwzfJ7I11Wzaq0+hik9wFbPkdc5e0pO4I1FotOFMpYn2NYh0nWH0ge1oQKMHBtQOgWo78/shouYm
58r5ba4kA5pqAgehcBnpohGPo4+I1JlLllsFHH63xDFpYFUfYT4Cwg6EuxpeMxABTnk2zNKv4+cB
VfBTdcbiJMaUZ5ghaUM4eRo1hzi5oD+I0Jsm7kLhf2TeZZ8AL+WZbiJ5IQnMPig73nRKzCMqwcf9
wetEFgNH/en7QSabyVVg1448b2WMAlxBFb4QqfTkcssL9iZlAJ5zVWXb6uatGT0oT5K9D8IlW3jw
KgpmvbwyFqROQ2Ti54N3PcmAWWVisBoVupXZBp+0BiCOWQ3wW5FQRwsMWqZfT3i/RQZcA1DjGQfC
la0U0GTDRu23nt00XYFLDQEcx+rhATqgG68b/QFtWM0uCPXYhSYhwUSruwCvcX60PPKjlpVS3F5r
Rg7VIaC4KGmlQNFimQKIfJFdtkzvfSRMYwMzZkfDYJuEY+pQsHJVn3YTfvWx6Ynnn/WOXOIPpKK0
bNvmKNI1sC+tUbK/8Q+oKJWVyvvvtTfa+Zd7rYoFSksqNP0zqaBAAg8zfsIE3i46cUv8kML83Sxq
TvePfH45+nDhnE/E+h+JbznUFA4QNTl1lpB6PoS71Q9iXBGQmk0bbKdrSddc+TqDvaeBl9Y37VmI
4ux7epnml0/jJcAW/yfFa3/6cb0GkgtMLsjyEG74dclk9xLldhejlXnES66ImI6Br5OqzLhKeADm
Qb/NiB1rCVTfAFI7IIHmbxLTmQRqz/RmTiURqU8zI/17rpYacTk1J4Z0FffbiMj3fUwTpxxrDa8o
UBiIJnfurdOSywOjNeeRyah9tTarD77T9VygZycVpQYyi3+J4YyfdvwPqwblZWDdkkZ+2a+SIx/z
MWzaAYofm9v7TeB98ao9Qz7l27QnYmrB7wg7liFJxiwMWoRPZE0BXX6Utkx8rUcxV2W2Z3t29AVo
mTt2YUZbCCwyMIWxUa0sKEFZS9c6S+R7YRpfefos0DJ+j61SXzM1OZxOr/dVfYCPZAWpuv8jYz9B
u8uihEpXKMBpO7X56vv4FLT8hhgnM04itKZdv89EkP5QLtE5Wps0Ldoo8/bbnj0cFsk1LMHXhYZp
rqE3rYEjcRhXVNJecZNsYOpdKuJLKnWz0hLgj8WVo2N3nsdDw6cfphSqpxqMQd5MWAMAfqJnrSqQ
/MtTiFAub5oMURJANgzzmYEVBR99jV+ttQ7s/DGi/yM4595Gee9jQhRnAXiNYpgNTue2zSN773NV
o/DWbBMRYNWzBWNbsqFaOUe4X4tZlrQEgbs7F1hIsvnILrfRLBN4s+PzpGjVO4j+OEkqHQCj5Bu3
Wp/v+QNfHJi6bQ81dBsEF6aH2eTdsUCgB2oIuo5o3upApaF2GPc/N+KChxHKEes4JBScoZ9Ky62e
UNsMoMyxO3MsQKYPvaON8+fsuvXAJvRZkBNhUAbjI/53YzW4ZH4nbWp95S3xI05SaCKEfGUV9gEb
0O8HoXtRvIhZUW8nv0vWsCWcxnzq++8eLsFwD3ruOMQlit6dzt9KzLAnLYsz+1PsV6AxdFwHJ3tq
4GRKVPrVdhwEkvN5znWQujrixeOiolXAhrTS4rCwOQGFrLU8EqWV2j5SLjPk0FQV5uHnH1TFrRik
ZotMTgYvhhf5BUNtTLdYoxHKjfNrTSsqUweLIQ5N5jfdeR2EjKKYa+/zvJf9J3tERARLb0UC/fff
I9rb2rnKEDbHlpf6gXMkbDP/o9EJjGo1kA/o5SJyQt1okl2Gtkeg2vdgu3U4dsBJoLgyZbaBI7VI
hnAiIeS7o77EvuylXS9V5YtvEWiWqbcnNjhYPY+gI/OSDU8Rog9vA+M9rc4mN8q7bQBioniYBQPH
0o/XGZ/+ABQ+C+7K8IcVq5LnXdXTFDbeAXitrFag+7UsGCUzvdCX6SWexcxTKj/xkTU6x7wdEtlz
6NldehaR3HLHl0C5+txtQotb3UXwxJc990i4lsUs+6jKNljQpHyoHT0Y05tWAIXlOlPE1SEseHeh
az3JiixmufwvxmFSv0UMLC2oDES0TAIolBTfwjWCgS/+hC5obGAnk1fuFOO9YUkv7wNGSTp9atLq
P+5XyASnxoqQaVHSazVPrLENfIUduPRuEHCM6VlFyCKF/3UltxrA1e/3VMFB3p9TMV/YdhgRi7Og
eBWmFl1z+3auu8KhMKYaPgDYi/VzmDktzRt4NDYXBZ/hbNwMgsjkOthaIoCf8Ejz7OceR5m36T2p
zM/4VfKMTnATw/sCCPvU7FN+HPiVG5k/g0Y1G/EzGQogV7lYgXoMKtkqG3tZDQUuGcoVz2ujXiPp
CjKwGaF7q8Th85q23f382AHB9Kj7Dz3X0EOn3IFO+F/P3zjkG7YTgpKXSm2cDCVL7tkax/qyUHtN
zQhGWqGJqV+1wTJ0ZAxb30RoKJV0BTvKI1BNC4GZdOK9pEZZhmGuAaCSwh+FtmLSr5TeKjtAjeKD
FipC+p7PzLmPt/crAErnIGbs0FjUJDKA00CmfhaxJHy6Fbpk+2s3xh5Uu18MnLX853CDdvxc7P3x
2pKlr0V06P9fDF7Vsxs/1h68MCcD5BGEiM/gpFOVHYPgaJcPp6lRQg0sfmY9XXT9WLWpEhlYMmLG
TaR5L+M5TCyKaKeh4L5s7ITUHCb5Vx0iBzv0yBhHw0nF9ABgMn7+XiLBfqiHPqU2cte9nxNGEMH2
K3pV+3PhbknvyN9oL6dewV9QGFjPmEESRZqU6cf7srtBkqHWEiZNZB+SszJomD9ujkBFHlB173Lm
62bOkZ1InBAJaS1HDJDyU1JblqdFiK8rF1ic17y9I0oA4QzJH9IH+iNK4FxMUphbngZ5ptqeWnAu
NECxMZvX0ckS0x5nL1sHtet231o/tfOs58NfaPD++/wsXaxgaHD4/syNysSMJjlV4OeNBiYQRTYc
qVDTfScULAyPaIs2VpEtDbC9BzK4pirJf5ur7UD2IrEVfML9G+B6/y2P2p+1HMG7QwXcY7iadz+h
X6O3WjM00bddHC0zZa1oi1BxP8VUkKBAIvpiskrCezqzgWlKR9NnxKUU3M4NNvVkE3IR/3aJoqSv
LFj0lwbEkAMLijoTdv3YeMZ24VzJgKoMPOlIYkX/vc5gtTh26BxpbWTmeBT7Gj9+gX3fIBcx7AeG
J5O8KbUC0L+2otsmaWauwEUmIqlaDqe6mjaDNGkphtG6pGpCPpf0sMYhju/K4Heaf+rYU3g5YzQw
Jc+EQouFGEjY4l+xUJTZxrEn0B3q4m83EjItarUFCkaur7eCOhPPTykNx6mNaWdTDcbDsc61EH+V
J5wkkPEWrQwf6HdA2EAvMv8OD11t5XyGdRj8H3S9pqIAribOXlza1iovnEiRfR6uzou8g/rQdzaQ
0dUPw2ieWMcAli5hZIueiokG1gHtEH8xkLDKAcFdYBpwnNhTWQjiLJXc/sJ86FJzElPMGx1EoFTQ
SXbPG5WNsQkECripCcFzsqOF9y+N2QL9nrO3lWVZzgdN1miKTf6TE8lDYGENlSuH+iWFLB8nGFkJ
jBEa9D5ngHi8vmDHfFzz98aFEsVMzMEu8kaCBu0GMIkVmrkzIqAcKe1A2Yy+HJJ+gXSZvG86vCgI
kPLhy50sVcdHcWdcZ0QAL7RV3FLexzVTu7VBk2m+YnpAVJnqmkYcwYKx6ragU+QExf9p4SjZKNXQ
Q1xITozhnvK0DRtomvsYZ/KND6yq8ns6M08ptM3B+nuXKa/uEDnzB040eWAlS/KWKMKcbOMeFmUx
Fe7TucZJ+0bvrWqRR1RUVgs4UGJGpAGAXkinIQIAk5bb3GMg6/gV9sI9VsDvJqr74/H8t+cDnRi0
8IFtlGJWfER0bWergBPaJuBfrV2ff57s3AatKQBIYRttYXsnaRUBM8bkGN5gIDg4Nm+P18O8JSbM
Nsg3dQAVJzHVCxeRTHl2u6/qozSI1lN7RGMmYnrgy5Rl47QJKqez13VcAPIrZ2NiJCI/rjGddCI6
LLBaMTmCS975f8gevd5XuZp8hBltCkVcJb5EcCKCmaD6i+SLWcWe6cTylzvHy0IL4lzK1BZKSJdg
G7AZa4lrhwqViEZ2gke/OOHRphuAb/0Ht2mEPq4l14hhU81nLsj1KW/VZ1YEEj3t8zZM2OEDFrGm
0x24dDMfxwFy+sKhbGNat60as+Df454koO9nnez4bXlpsOk/6vTaIx6AmP+MUulOONcn5tWNoKPQ
i+K+aJSp2PAWYoI6nWyUFYRn2Pg19JV8iufvYlHYvNwapzb7BYq2DpJsU6cId5J6OZGk1ebQk6bq
yBaeeIfq4aYG2OpzIZ+4FSzAx/aPjZNctA+Y2aSq0bhMfsnMuCMFrmAawJKkZD3Z6Obmb5pxtb8F
i7wJXHO5bs9kJO8UgjOxue7/+ILYjlG56qm/pFbVy9XPO799hhpmcAxIKMBioWdLXuIcRwrCqH2C
VKLYEzD9nM/tX/Azx0llHw5SSygVr8ChT1OsmRX+K9e4X4qG4MiBYVXQMWSp2z/boNSYNANsyrRm
zsSB+dtmjDdwQofzUpmHtw7VJMj51/sQJAE0bN6cwHCBeBLbg5Vv3bTjZ91FlcwYkJtmEoiqH1cU
eoFlc606NOGaC3lP7levrFbmPa936/apX6+EVkXWiH20T3K1e3p20zf/BmCcCJWecugMUEbw/et4
eyRPD80O6oepFm4g17m7irO9zOlT2Hm9aMAOkpCOc7d0+NOuc0Vj9IXrYbtVxvtV51rifecGJ2ON
ugZCbl89+hm4k+3CcZp2CFUAgK8FYUqoPIN5BXHy/YVAUHgsBT8BJnH1G8CxQstfDou5yi/2GkBm
zBQcUbToPqz/tlo9RPBG0CzOljwe+6SR4CFPJflNmAraB7cdgvVSogv/NcZvXbUygBXBPG1P2pK3
f10GKDkYSmkIH8/QKdCwSfG72pSmJW8aifaRCKy9KXq08NfjlCADrO+yUPFrheKur0D3eQwI9e4q
VKIxwSzkGZb7/NT4L0yjWjWwZT6cDWyLlFViwVjeEML1VcatY2EbjQ+nUh9md1MqcG3/Vhu8BxIU
5B6uSEZ6d/cv2rouqmolIRGik14qEaLaj0qiGzPFB2ttNOFwuUVjNqvF4wCu4C1WQyMesEh8vS2Q
29QqPxpYpyBsgNG8vbZL0t80PNWEu6fpDSCo3b6kZCG7COdrtMhC7HPCJnjo8GKwL1/q9wHuUMAE
u0XC7Etb/q0tRlnLeGe9RL8AutAD+Bp4kUveySviTlMJBG5R61JiRnYT1VFzPWQA7GVI0I6ZxdGe
lxa57hASqe72UCX8A+y1BFJszy0qsBUSDyfZUWFrhV0j3oLaZJz+7uVWPa1YnQ8JX1Ba76L4a47q
7NBrle0fQltg0DwKdeioaq2EMmu4HOLd22a75uc7J6oYgrtAJ3bSGfq3f6DgL4FDbbDKfJ06eeaf
R5SphaGFLKQ4fhbLTMsSKJKd47CRI5YXp9r10PxqaYVDlvYzbOxjnWZEuE0PnDgLggjXc6o9SidB
wjMDVfjV19V4ZlNPITpKHZ71iMlZY3KtGS4dGIholQXK9fYlF8XOrouqlzaLvmJz+uOnoqRA2PIW
X6KTmirsU7DTTl/BxTUqrwl3yT3s2MSNM2oDGwbRAwF6e6a0oKTM6W414GT5WRYsM6V3Ye8aBngf
tI7ZXzQPVwXMu1k9QUbYtTCRC5NYfYfdqvCq6v0c87z+a0jvu7VkRuRVcdCTEVHWBHKbvV2pkauA
giei1u71hj3lB52S6iKo2YccY+sEs92ZoFIwPjdWgXS34iqdAk5jbxFDeuqo5ep2YA3ZeE9A6KSn
bKJr/aKloMDP+CxhGSd7nD3FMKKPhLlBzsTWBygXVeQzssVrpoQugeQv7Ck3CZ2/Q/um9wGeGufq
Y+KPjzc4KFzS7UgaakdGcLdz6PKys13D3rdkgKZizGqFCcAVcroHYgn3wnVUv7qr3Lo0mi91G55O
nU5lR6qXyEQbPVNszq9nbNGJ1nn5grwBC951tWKVemySziUcF5ucsKXkx/yvsbBOFKRCdIwcW/6f
TSrZHy6NPUVIxBF1NuvlFsdAonQmA8+JiJQNnyGF2dVdTbXnPFhTvkecxO1zDpy53+jf5IhmL3+B
hZmk0Sf6HTN4JaI/t6I8b8X0PTgOHrPNzcz1ky/tfVYrY8f3gLHElNabJMXRA2gMGaH3MDRSFgrl
TEqQqLy/nQaMIV7aV36eKFvSYgkjX+73pQC4BRH+FACGFprVd0MCKdtDffoxPN5BCk2xcuHx5m2m
jJZ9i5bolIgjmLxsXadWJQ6ITOMe6I2+nZY4/UpSQ82J5JItsfkEY+nmZQv5MADr0M1Caxv62Sgh
RpTvZhvwURHPF4Ubko3VPdmgZv9qkA4R6zVRl5NowH2IYdNujgAyOQVU9/LY6ocGK22wioWr1mZA
IBzhRIv6N2AFU0huWqtIwo9jMMfoSENWe+ibOURMuwtdXMCO7v4TlYw7QOm5P1f5CWS7decnYxv9
ePZt2RPamlSsKHigjVPOGnYz0b1X/fxbp9wd4z8DEOPX/XrVr0zJ5iaHhn3pjWdCwwNc9TuGwiTA
FWdwpWzXz/AdeuoVBmAE6SzlCjnZWLI5WBuiUfF8FFbojZmLm3K6gSVG6Bt2yvsZLL7nespcjNg+
Wt5kyO+cVPNQMW8ipkxGvy8/RGo1QNlX6iKGFlhsXmc3aLpZDfPB5Jy3EVeNS8OPRWuJSFcDXX7o
AKC7hNmc6Y8gLrxfzXT7el5xOmn+KbLrmEevyeXe+L4Tub7whDr2kLZAY7w3TqQKB2FZNSUdQRok
JhLozbJXBy0n2hu7qRF9a5iB+WwRkqMx7m3RWp4nzl0HtRUK1dms8MskUVxIQ0VmCFcrH0iuxn0U
Or/IcdlaS0v9QKU88B6mXbmOyZVVJtU2C6xbjeq1LicnC1Wbyw5luGZyQfyOL88OpETvURiirGzM
Yp4Pgzu7hii7mh/6dh0WLPAIX9HSiaK93Y/gzZjbYkVsJY+BAnR5F7SUG4wS+ZAPVzIOMvb4uZRz
EMr2Hfl0hiDaUIwKFP5dlcz+OW2IQEW5nfXq5MKkebok0My2GlW65/3mUB1kFyJyLMKHB/utDyf3
TzSANM6VgdbX2oZ3AqKOsvpC8QzCpCJTzL+YqCgRtvYlDT2WJIJpWOmBNbLw1GB7b+2epYDl6Eub
jIoC3tLHKbzOSPhoRTB1EiXTgF7rp/MD8b57EF7vMbz6+iCb+yghaoO7qjZ+PvgGW6fi6phg6E8K
Lp4fNTiFWaEnwFH6k38z5NgzQOw+PulhOYUYaLMIL5WFs3AfMTBdkrniC/QoKgxegj8/9Rc8Wbfh
nY9eood94aXXo+wH9x9JJLS9IMOLK7ri4+RZ5uQSgiw1hyGxszciqc/89gqM600XmOhieaL9EiSQ
igPizq2cElUFUrEwjyjYBi6bSsAifD5ML4m7bvNAKntx1jF57Q+Vcs1MvS06ti7pbG9wSSDJPCut
7hMDaK/gUhYB4/prr+DaREGiHoBR11LxFqJn5mwzGIgLldrStxTxL1wEU3xD4l3luCRjybX5wyYY
W6C9/enmQA3wgsbv0BZP3h49psav8G3lsP4W6P5aKNfA3miXBQnuvUyI0j0bINexGwdadt/yxPxY
OsaJuEGfrMwFQBqMU2JEB0lXwnmbnyH2S4a5uVjdfOAhGd5BjmscKnQkWlQ0+26hhQEF3KRidY8u
pPvbjNsnQRRuirIaS+2liedG/7uC7Mwluy45M8YFTXQcK/YLFy0cynw5PlI4O2SaKPp/ElGcBa0V
Edxl1lSzElF4iReEFCOTndfx5u7ayHk7muGMUKhxpXZBXEj54vk93ieW2kED+FEKfHBU4BILEtLu
tb1NgvrooUVydveCtIFAJF7P1iXueUT+wvJf/NiRHfcbGfVF42NCoXgkgWgVGiFyOVaxAIwGvMjV
NqH+39+7mo9TsjexGxUpwo2xFC4fwvcDq9EjQ8tPet8BtIbAlhU+hkrbLna+wIrMayqcWNdmLZNK
UsPL1/KKbbDf3clHg8vloUWE0JsUuM8yJRP//ujpj8w5DzBdhwu8mDi8IlWdpJNfMQjGLnMkub7B
DVtGytgQTr+0KyBphPvbt588Wc9C4L8re5tXWtMlexXA0ALCU12VapHjErJlQbLtZILdZwP/IvcD
5TMJ1PhIZj5d97FV0dNJ198/+oiWCUgC72W2jk42enqY1+FFZ7946VW6Mu8JlzDbaSjdXDgRddvW
jLE2APrJrZwDS3qL4TFMOumnSX7XSOKFru39tA4vdPM8KV2lCRLK419mXHl8xEs4M07tNkM6liCc
/tpKR1rkFxBoz2mOTF8kJxLS5vwu4ip+vgjf/pLM3HTisrcdmdP+JRNQKRzwgiSRkRWROgL4ckEd
iXFgeVtz2araPppxHNTOTQL5J2yM9q/UEGqS2qsW/+K2RErPhws+UHMOYzFshLGN3nAU8xDcmeUU
jPGNVg3Fdjiz59GZtM1srIGtos6GKh3+lCAD0us1uxqT49cmUJpWRlYUrMlLMOEWC8yyXGGWZG7n
jBi2LQ8f3HncaNDG3Cvi5ts6Z7QzqAUfJUJ1xYyYKHDpNqB7FvMAIHGQetLMn1dvfgw7MlSwEwrq
DHN7pQAt/VjLKKeSXxJdzK/AlT3Fh/++umpXE0dEmI/01smT7wIBeDRuOQ4Anh9c1eo3kLOGc8h9
PbAjxWfQkt/3iLpIRuUgO6irpQefMdyLp4gdigpXwt9OzNzbMT20ufjkSexJtUTDDXJ+AnsTSg7t
QDlRxnUb42kYNcuaVRcjcp10am/DIRX8hYSpJcZKBMI0e0wqgzE67nGFMnzmrUcHWy1dTafIJ36h
ZKTSRpRy0ZNNEZlauZ2gWWneNB3mspmNspQz9wSf36TuH3bNLlLB/eGCFcM1PpJDVP0BMEjtIjTk
UNIEdKmbIbsBNa1GU+D9SFS2I8sOhf2ebVKR4vySrodIuvSVfOXpzt4J9Ne7ZtWxZ2eUQNsZRlP2
RqfD2QzFUoq6+COvl9NyjyTzVitU+NKRGa8cduy12ecRcmv12TLrFJw/xWDfcR/tLtz+zAF9KNB2
pViA+PIhs9zqb348BDSujMFETeAn/kol6avxts6eBAHN7I12M9NyvcGmdmBOtwg5kOPFISAUWHO5
m1MVLt8f8Lwlt8ChDsk8+jEPrtZl5BXOMCazrzXwa0k5jnnEmdKhc9q2kVik
`protect end_protected

