

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SOOYAbmSVdMSmEhVcX6OANZAlRBhIeIgp+j8aWie5qMiZZfkKWRKGFlDj4dOK2MxGgpLi60kolAl
iwo8CvQQmg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XO8hvx7ayNrMYNs+QowHbS9oiS1GjnY7XWvxUBWvS8S0pBwgguPJgxI5Jawjx75IEBra9z6gur8D
+8bJ3wjB5uOzP0Op4TufbsYZTMy5/IRaR1m1haAiZDNWpnRaJY0iGIl1ZfXnFFB/FNm2d6rg/H7b
+K1wV2KmxNsYmhxGeUs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qrXPktUjITPZaeyYovMGSvjyrwEeWSEPCoXArB49zu0J+taotc50izauZkw4BvtuT10+TUqV3pWu
H2Y4+wBhbI0avNdhBTQ6WysNgxNkl4xSoIMSUDeWLPrThpvXqf5EM2xFWnYEsoSt1fOlTzsbNp4Z
xTF0/8eRzGcTqQK8goNirFS4li1yNxnvMyocM7UB0Hgwd4r1WhVfwqexmsE2F2aKD0WceDfUKvzW
BkaD/pggzoFKe9ZBj4krjm5QO6MJe6tmyETtklCe5Tp5KFVAoUG5SSUacYfOW5JRRQQN1B29KV6+
B/PXOjnEprmrDoW2/GvnZUOJ8iICUgvcDDx9Gw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RfdpJMuL5lneUspdc3THLHWNRfMy7ZKvo7MAlgXNSeMyJ16shj6csIbQx7zWlYY0s5cmQ5qBeuky
S0nRybRR8cWMHwN/9rEo4V+uesao4mJ5GbtqRFTH0pGXUIW0hSA/qLXBAZCtANiThLFmTTovXGQx
QWChhP7QcQZsZBRuEUY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KfAPtRUOpYg8KaNj0Wxd1r4Bcs5Lt64mregrxrObBeYBNNIje2iGcuv2d5+PQzzomKwP4NoGlbzx
CSYz6XLlhFat5X0Kad65Lvso8ilyZLrxVgz/cQQVMyGtqJsflyi+jbqMWdWQzDlLboEzDolIGqLM
T16l7bjdTv+UHoBJFQNNpgCUB8RCwZwGjuOrDkNOQRBxFbXP4ewZBD1TITGRJ+9yag2oeIszJxFS
OnxOibAvqbpn5K7zetHoNiQFD0HLxODP6ACT7OZWy2QVwDRr6smLhIBBF+7E8S7up2WgvZZ778OW
7Swo175PkHbmEfmpa+y5XkNQNOq7GC6XNCURkg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11344)
`protect data_block
466gnsh8j7oUBnaKygiRp76Q9MGYf6MUWY4rvwt9ng0HvW6rdE9ExABje0ZKVt/QvOFDL1SMeJNk
a7XBGeWeTXXRyUlUYB11lMifGP3GDQ5TJTXdv4fcQvQpcQLiRqLaVCUi7zALXgeAU39i6xnGdkTC
k7cmBViprf6ZpPRAjYRKHjWO1Qi53bwtpCUnaWWIrcCLuZbMWHu2nenknIhNzyR8QVaCuI0GoSLy
Ybv4aSZGOl4GvE+o+40RFtp7/nP7Bko07V2DTcpvSekdLxyMeOUdDWfvBKWf889bCCtcH2SQ8ouB
NEXm94Z9Kt0/nnTlNZJV8d2X+zRgGaDv8l7XgXzZ3el3y4Hbd/iQyGLY9quPwlkKBGbkT33mzzxo
GC3TqKrcRsweFyrnXkFCksxnB0+2uEcZAkeYOahU6UptMw5Mqf8lDKUCSZePLra+3GiFR8mAYsaR
R/15M/msx+u4Ddliti6LWeuy9wdcSxxeMui7i07ejV1WjSQdYJO8nIUkipR227aVZNjjqCN+ZRge
4ZOyKp7vKJprD9KMaecNT9P/FHIQ1kZkaFQm9/xCY5qHHMQS0zKteBzi9im1wIDvFb9Xwv0B+voP
Ynmnhksr38LPQUZf+uXfcuGTJzCOjSQpnlMRAvFBqBZiGa5rTGiGCL9D93WE2zbY7aTOwUee1Wfb
BvQ8jogKLu72pezF0N7gDgm15L4u0aqFB187fZj7Ek9DQ3GrB8ayAsXekeWig1K7LMcnHAGb5MtS
ktdVt699zx2VEEnCuL+UKAQdJyHRRkNfChYSwbvLXeiive1i2/fGtq6BWPLMxZLhPV8v2PfSnkLi
lUCBf8XK6FU9uPjZkn8Oi9Kp1V0ednfHkwU7g/1Xedk8WfB/YfiQpwC1rQLS9lNUS42gCVCjEe4P
RcKpzhNuTNJWRC6WzqAWFOIhrOit0rFEztzUeQTpROkv6Thmtj4bYFNM7eRD1DKztJQLcITn5eSD
IerIfmrhAXx3W7xG/MR0WO/gPzmURaDuBylwePQGGvYhE+kd7rgyt9NeVdFCR7TM0PCj5UNlzkI7
xWSUIQtcXvdanLm4KJO/oGW31bBeRccsoaIpEta6Dc0UOTmDp7XDAn1hTRRcIL2MfYMI+AUrfvGx
iB03HoDWKFRrORRHPJHWkNXxa2uE9nLvD97tU5bdiIXhul8iE9mVkBLEfB1+Xa2wkv/ePBbN2vJo
15WlD6XwVveNIZu03DYi5uDpVBF7Ol9K/y7uFNLvbYiqlgpkiuJvPP4j7+KTEs8etYRYkaiHv3iG
xqbxv6AImf+FFnH5FxOQhyedryZElb9pgL18R1bqDIyJjIoDfPV93vOIsJKRAfK/TaUGa4DEOO0Z
Gm4SB4+v9DV2h5NL1lyy4pvhfA9r5xH3E6erEgYl29ROg5qtqygvDuldYZsR26iDIF1Oo4WOkfNV
spOO4UpV0UcCkaPTEMStieI7exg4k3OoyYVgTTxVvCvtrGS97naIPX7V4icYvPp/tsYpiPyWmAZn
MdzjknuyhQgedGTm0viOmlTWAqa9dbcw+eVZGdesSaay/s0zA3nemWVf7yPp5itjEE/+0z1Xbv8Q
fqc7mBeMOkmnYq0jO2AbTSrhkBma/kyGKH4CzaZpK8qbQ5OpRk9x8jmzScHs44ONZ2mlPiGH5rTk
BYS88x7CbXHWAO/vRpeYN3RIRi3cM+EUxqoiCivGq4rhkU80ELC9zOnsQO+EJkP2wlZvGH3+Vovn
y08apQGWteFIkRC8pddu1thYg0ZSNHiYtO2WdIfmfrVYuwW0xXqpDEawLy0l/pSDcYcIzHG+jdUg
kjw3T6IsOMXDsBox2Pzzy4cG/3zRniO8znx1WB/EmxyphnWeZJDAULUz5wrGHPPG7ZQehc3tc27r
eZQ7AP0mdvJE3Xt/3TH8n3IONzDFI4ivzrAWTwPp6xfhGkkCkKNzM9mZYa1Dt3/UP/w4KP1EO9wg
trlqGGMnjf3i83rVEfCP9K5KagsWvRS6kdFiikI0RxVcbsRDk/qQrdaxzXm6Gfu+FdwWVhsz5Rid
zKmweD3thgTs+q9snzeU1dYErxTmyjPp0U9jwq5SYPzi61Ascx9DZoMLZL0nFp3RLLFZ0HQhk4de
eUJwmvgNNGOyCGxQgzdAyuNZv1YO9oIttK5IF1yjiWQElOw2DeoCT8xjv1LdBiH98QTktaYfEP+a
zYEa9bE8gBKSOnSwgXoJBA+bmWMjLz/swtuzlnrKEjRzISDj7QIS4s0KbDKbbAEBzDbfugkByJik
dv793fFEWdvWCsUTqFgzQH+hoUHYnXgH5HIjEfq7PTlUK/JYJ7lUVyJg+PEeZCAlwZlO6kxbabZX
/Fn9ZLnR0b611cg8IzvylXHSgVuX/2bGmW2ybkN81DXI6P7RxNEgKpMaO8lJ1DMOxy03iB8K30cx
VUgcqEFWhoww2eeUlDYuGcIzRM8hr/s1U8Gty6l3ZP6LAllViU8b9GghIql+afrDHgCC6JQDg0LT
uO1YcFlrh7InyVn0dTNm28O1xaOixBGC7+wrAWrtSwfKbZy7DqREkv8cW952jYCru44TlEEc8asU
2Am1RcQXFwxIkyPsZGg+eBAivKRLQ33I8gI+AawTXP2hj8YpJJW22/yEVkbkMvg0osTy4wrSmy06
y3MhYKiqMufiQaHFaLc7/rO4scUSPGSXYjoE6WjbM9GA5TO39qWioCzH1FKLp6Ecvf9BHQOSRrSo
awCXYfhLlgLjXi667zGiBESE4djLXdrUxWAIKH25lXCHXmAU3pzcgwUl5TT2LMwK58fCNsyw+hfe
AcZeT7anZjCzwXlQugq+WpP6NVsC/WI5U/ZTYWFbuVUJOO/ZKlx4V+ir6iGhsB5myBwmNH4DWVBX
L8DLege5RzGiJsu3XDuFspBoHpFzCmi75V2paOVfQQb27V3UYwE7VlNyH/AbpW6AQhgZUfUSef5N
MUq6R9ZLJixqzCXA6ynAhXKcnQdSIvRA4TLD54mcIGVO51xM9v8YZl0VVXcg9nhcX7LrAAck4/Ne
MdD0IMi7XYTLGLb9B1qKXLzaeONJtUmJSFpBZmyszwnDrVzEHE2+L8h6AqLSUsMS+xX+o6F0XaGZ
gofl+ns5uJg1ex7GBHGwg/dsJNInJPDG6S3cP3DI8bJyCEJgM9UBQqchma+hXdZkzuOYlFJhV74T
smD9+hPSU1Cnzb+IqPqqYifJgWMVDx29c3sd+XPzk4XZKBO/6epzwYY/UvlAeXY8+t9vALewS9UY
AsqunIGMrD6qktAd8wX+tIjpboHIDj9K9okygJkqlSV0VTKpUisg4cO7AE50Vph0ciy1E9fYezpa
1KIqYA/His6yg00ZGtTgHfuX4vbi0o5MGQgxodOfvdQRnM7+nVvufqrNDC0JKnWqCZDyhcpBIreI
IgJIlw2ssOQ6G74SHbvVhezg4y7/Qrx55h+OyvPumcNO0bwKu3E5mrWsGVunBm9qVJgQNjhIRQDC
1B5GoCJDvj7OxPHQbwjO0YNWnmosL8+dXVKMTArjJ+KhTIf01aY+ItsoAD9aj6J+bPYMWKtrjt0W
TQcisJsUKYdusyKGxyg9crYKKEqLePWKItBI4jJ+OEGSXHAzWYaSjAhTpD+PJZjz5lbEE+GcYeqm
Z0D+Qjdnpra1VigMn1HVOhWeFh4eAaazXy560Aycdmdl7ZDGkUu0WTBIFOpUpqVhIqrQeLcO8pd9
PqPVeBzYOMyA6RZMa2cre0ZXDAlJ6IDHcDEVMpmZo+ieFLyi85aFWJIBMEdwhBOccd39IzSDDJhy
WNLzJRL+AgjniiI0Eu3pmYo12z+0sdG2jUluwexbXYRj5mJ+o3RCpXa4ngjkqNAumlydMYw+/Cqp
231kYzZg7UajEg7Gpg2egikQD2r8n8Ar9CeR547lqApBHs7aW4PRLG533zyIC1rkLXTSQYhTnStz
Irlc4XgjEXaFjfrVrVS9bqANJWhzpm8WJBpvFyhcAk66F4yY9RFAw7x1h8giU+KUaAOHEw+Qs4tB
IPGDtzvxxosYBZTlgzpH9U2vYdnLjNgN1TLrmIyOhveVrGX1QxC0a90ZAyIDNyVgpCKRidbWBmy+
rjrl1u9BPvhcGUyI/O3zL0f8t5TJ/ecR/9N7aUHebRPz/e1P1wY826osts1hh6E0B2XRw6w0EuXT
n0FEoNoP7ha4eLkTXDueHaC5eFMVhJOOqNcZwG5IikL7h7KY13wPURb5Kcs+/jfyRZCBLoGA7yeh
EZMF4JLXSQzT9infHWoGgCgt/GL1GMR4/WcJ9plOVb6SdJKzBguDwCgAvGrFmD5s5QwuocJ4qWhi
4c/whY5uzfwHbMZB5XJQyKxOfebJBxNFPairGkNeIGhqQ2Tpxk6yUfmzgClbSmK/7fJV5/KW+D8c
ISEEFGQVDWdopKFxJ7WTDDUbOkW7I6LbYIjphgKPxYeSrKduCeUds+eHk/wAtWuzj8i22dv9WQG4
1cjM1RSGN6Y3CJrKXIL1k4Y23zPT7qLCW+oBgBdFGDXDu9CLSgaquLQwIL2T84HWgezIWzLNHlkF
mrmY/T6R+pihfKTwLelzk1kW1Osm0Ddmotj68ey7nu/7mPrR9bSXil3Z0ibx1KJeDybQlojTPY7Q
BRsKITi+IGjWkZC+67ApcCUlP9+JBe0fCIk2JMA5pYB+E2Iy3NMBHNDksTg4Nefrw60/11/P4RKh
qjPOHfoMfLbSnCUHBYU38aB9c1PqactvJhID79YOPLF8EWZJl2d36koIOIMnPS2WHsyznHS0AQN8
JTy/oGN91VuBkaBvJRLXnlvz2E1tta3pTeGF5l9oedx8J7XtEoYP6DPNaraQAyprenFKP6ievDOh
DgAFajbtnSUm/cC4jayhN1uPu4EhKoRhKVtYoVZf53rnXlEgetZyMgkvYOESrLKhYKrL6Zi0jWmg
zpNFRGjbFFwi2V4ojkg9oo0WUknuJ1JZM8gRghRV9LM5n7/r51GtZ+aSXixeOAebH9p77SWbxsxu
iEdLfdXVr32bEWXjiFv/viDXDraPvCpgW0m5n27+JiyJAixaHHt+xsjkf9/kUiQCgLU+x5YPH+0f
agD4RLAtf2ehEh7w61IPs7P1V183tE7QKKcj+ENaz8yg1VrDJt9+bxg1vkCBzeDfXpwJZ31yyvty
zti5nHhu0w+DuFNu4Z9XU4pIIcdnpZRIMnhrbNLpMLKGTtcVTtcpn1Lek1A6PEmj1EBrl4bP5uvD
emh++ujDQ/XbYs0LA7nuD/A9kPpcqQMFPbcRWuncDojvIlrcYtQ5EURqOlXEpuuBLJ8gAhur0CWv
yPyKe8Y1SWEqrVlbUAjiFXXEzI0IL9fFkfosJfVhROH4xLoxwipMHuQzXfbJ062UB+gQCJwU3uo3
IhAIdBzpKzwMDahycuG12JOsqhN3z6FK6SohVCVqc4ergBAXSaRMOOivT2rXjJtpoq6dNP2hK4WV
INhvad+oQheNduKsOvLLllgMAimJbZ+VHDFRH/wQRuik4y4exCXSq61LKUHNKd5ic5dZeQ7inXyw
/Qmz55GcWDsc+b/oxXYS+qlI/INHvXZBT92gGlWWHqdybXYMupkpiq7/0FLm+4L9yyMAvh60qzFj
wVFwa39wf6Irr7JwpNnC2G26HJe/kgQTSppsPHDObfhwqxUaoaKVUruJnTQYfX2friwxNAmB0WvM
QrcTEkuGik0St8UPORZIhjyZzgUxxUfZ9tl7qe5eOa2L6jx2JNMWXBcfHcSO6JKYmV+ORHY3n+US
ZdVDCYRmHEkKU0poeoH5YkEHqxggX9DqGvuUJZnlZTFtjngJO3WvwIPW+6EdzsX/WhbaOIdcbZ7W
20/4jO1BcohdyUJj58S3YRzJnG8+v9wbiDuR/WftA3cMYKYf3twu96jsiu0x/KyxbE+tyy3DyhOF
AAqE07DCfMXAFaaCunvbUUSwSoWYU5IpKEsEDcLSMoZG5JdUddQXhFzCNaUhRtfLweRr6LN8lKIl
j9Ry6fytpAH0JMUaAHDZu7Ngwy1E2jrhWoTDS4Zye+zDac1WwTZhlzcpMAbcyRaynvV9Rm+qzTkF
TdsJWhupNRJAegge1qr54dVjRMeYITcCMwvdbycSd+ePYgTaSNgEIvZ7lYUPsV6atHrKmealBVfp
tgHPT4c8p/8pIIYuDXskwbJXmV2LlTrRxvJX+2SDExN2SGZCONIeXHLxo27BHrabI0NUXT99y7k8
PNuaXv/q4rF+y/i1r5Eb7c9Ijlan4dAOBGhLOLw3fesXQkTOk9+dhqIJjWlbVLfn7wDJm5uOYvfW
fG2RNKc9c1AarX2F5IAG4Tz30CjUDn/57XJ8xsQYKvr+dLi1cc3kQ9ga3NXciJL444y8m/Evi99W
2pNYI1PoFa3BavYuAl4+GBgfzknJTv1ZPisq3vhYxDo9w26BsSGRCiucENYPWzvNcnM4rIp7FWvF
1WLvl+Fc+yqFruA1uFBEaebBpxGckprBKblWNUzNVs/P/CqJyMdqNEyGlGXqNKBVuF7CIuzZXlEw
PE0hKmfmih+BsHoPpwayCmZkSQxer2Hw+5wnIN0w4kvNwN4B9rBvRZKQvqVhzoiN00KJLgYjG7of
0wop+hIGnjN/2Bpd/g0UEBW4RSC+bbUfJXPsrBaejKozk6X496WsnhAcIh0fp+eEfbXyax2Tyu1M
tNeQXR3ejXIp53kvRvX+25MKKuGESpOiYputdotgClxq5hT998CXnXEjS66aaHPmrtQm8WB5T34F
D+6KNrl7A3hlbKYvOUuwr+CXi4pgIsnIGap+X4LQ8Nzm3x1OfZW/5mmjNvVK7Bz3hpmElWxRmn2d
PJ1mlkx8yeOHXdaILub2pTBcO6Xl6bQBnMEbXlwSmwSLtaG9/Ra7a40h0/gcpArXRT9gQtEp8OPe
B9AEXPG8Q2zbgIlUR+r4YugOLO3Nbs7tD2eFIrNBu7crloNliHKd26F6qnRpZ2GD3Z5+wXxdG6D8
hKTpV8w8qUtzDvaBfpi2BpYAmZtxXOV9w4Pk/AvycFQVkYN5zuqDqrOIqhrJ4l2JKbHx5QwYSx6A
OMSXhIiRAYin/G5J1EOZ7nmT22RqqoDQeOgiAXP8IdxEno74NxgXZbiq/YIbCE5fj3aDS1Z6kUlv
F5oa9fcUL9lKjRFT8sx4rTZl8nhWb2YmWKk2ZzbnhlTVRwE0VFmmj6jpyFZD/HpVUGcc2G5rWm7T
f35o1m5j0uQuaIMlFmpYQMDgrsHK8Myvj5E4uXuNvE/jFRBhYvHLDME7uU/VB9b0JqFwIS5brHj4
e7bmAgOadA9glc/o8MZUgwmUEfgJM1QXuEVDHtYJ+Qyws4mnbyEs2Z3UIvcW8cGM08PmSdp3wRMz
rfKh7hnr+3vWAmuQBbbeALTpnEaYFtuRcBTYr43IXeKjcMra7KHdF6VuRuO2Z6LZKn783VhNuYFo
/ivFxjzpVzIXY0nhNscHnJeBa8VrYeIS+ur6O08sAFLZgbz6zJAr1vNsohE+krgKbmS9eDZjEv/Z
7LGnSUrSqZzTjvdygqLWMgHN3+fB+VuAxAJIdSIOcVlsoEMdrmfV1l/6douDYAW7iMX43hH0GH6n
Yu0j8EHw7EAyy3LRDy+pKbwxQNrAQtCkIYwONhkAeNCU23kRTKI2IlDdFHVKL8WDJUacFimqenUu
Axk7Kl/PLI9feSQ9ETd0kXjiMYOGuOxbHEFdHK10VyuxLF1VozdxNlR29UPuaFNM1PepnYz9MpRk
7HKf4wZxBtOUVHITH8vOI7xO2C34pN3PtPf2G8fmrJo0p7kQY07/3syS9COFHa2m8YmkS1mF+2HN
TfREwitdogq/6wYbkacjpnxHjOnO/aUsXlVAd1twor1uAcOzH5XlaqRzlKEzH2AY4QqgyKfDOrl0
LE9wCvBuKk+6TWt8oZfKHbYm9Sci/AsOfMOVy9o3oO54e0hjDiJk/DO/lqZhdr85UtkMjI2w4cfM
0HHRXFpyPrwig41P2gbfES/n3iUHYhy6Jv6OPrh6NZeYjnIVVW/B4QVo0lF9NSHTSU//SbTNBzQq
UhJ3CnnsBE/FLPL5L1qLTLt67z7FDZ78ZB7cSt7P6HwYGTXmKWnmY7eRlSXL4DfwdeGE02THn8Q7
zBj7bYPd7ILfy0lfgs8D3TZtVxfc9fL3cfB7E9FACUaJRuUORCK5aGIEislbYcYGAUMhp7m4n1uz
So6/ESKmEqeyxH+7kLUofX1ZgYLNKLCqyBO6/KsEkx2rPDPTEv+rHwUq1E3fINE6p1KsJ4emtwBM
Svwk+2WnndN/UKJM41BXvjX1OCRwl86WY4EOOe44Bk3b7L9uNTVBDHvsLpbnFPQDE6GFjE7iyBFB
gM/uP0C2X1CIG7MeygNeKs6UznVUWMabYVVyY3j76NFRtg757pcpll0JBQHaN2/BDo7sedZWvmyl
kmQAI0Sm/RzLJojuPkaAZVG9X3a3tNV+EYQgIQGJo3f1b8aeFD4hVbInXydPT6UuFGsY6t79SChs
VXetP8csFcmiI+3qjORvSoWg3zlKTFKNflAeUewp8E5pZi6lWhIZtCv0oen4dwSPUbckHdyMtNRW
vUm3BOlHwJhXkC9IsczhrDWlqa1sO5SlADJZ5fwbEsM7DDjcJTx7gfirqumi2GB4JNlLegdoh4Hu
RrdEcZz3EMnIlGlwTlsIYvWDbFdfpM9r/kCQov/PQ72rA9vDEM+/Jf0oIB0rWzbXICsmnbNCXMdW
7VvyOsu6dw1auWkJ2J9WYHGhKfMXSx/6DMzGUMxEYod9VhkNxLPr6G2iK6/PvhHtvMY0Yw7osXSZ
hBdevkvGqP0peer3BwpX4wTpaFnjvLOAWFpYGn7AEepZmPa/kve5gwGLDt654RmOG/bCPn+MPHIn
m65iUe0PDgZRqHPYczcuHtcn67mLOxnDffnISYLQRbu3yciCGr7h06NWbdLuAYPeJqUJSKCyiDFU
Pnq8eqRFZutU0TgNIjRXwCkUiABXn47SCe0I0696ZUtN+LaFZf2xApV8aN3ZJ3VKW03b5Vmtxpkf
rZNbk1IOuFi9h5lrU4jz64CvGVWjBDbEJVKsn5eQxkAaDXgmq92kQ922Wvt6VrOqq0ldl710GAXX
a0T6EplnkbQfjymnSgoKdugpwuv9yVZzKtEJfc2Mpb7kqw+HeuJPVCDgl7izRtlbnDHMhhEgBtmr
dGg8Ah6ODoXzx2DwJXjnocrL6+xzFRYNmQCC2ne4TJVhS783BiH7a1GTJlWGAXN3U7kLjOfoWK1p
9raurrRJQ/vpvvx+nBCzA68EunPW0K+67V9bJ+PZEz0lOrMl1O0NMeBuFOdq7R8i1nfNpARsMc4d
h21RszDskg1IliERDWmo3o+ykVBZMQI2XJf+5nZl2Z+IVtrxOWmh123IidoTPT29yqO1fB8sxdN1
SJjFI4D+p37/J4GFTUBxVD/MKEWPBMIFOcJ5/PWjosPrQrH2cxXuVzyLqEgG8Moi7IFqhWKxt39h
S9r+rvBYwCJIo5Hbzp50k0QBVSiNxghf0x+7OU3c0+0klCkjCcUmZtytFnXbJg7paIijvL5E0igQ
2IDyFWE1PJ4/IVUxf3aWZf7hWzGA6lqt4R/Od+lvJ3EkxYDcPEC7/uAp9e+acB1MkIkRzYzd0Jke
T9RrdbaQdET4SoI1+34qQN+Z6ZxchTKNiFryGWDyUDIe9zfUQeCdsEdsgynJ8fdIXGSJtskomAtd
RUqR5Q3AJM1cL+d0fc8dUpPQJXAs1n0WSLYP682rVNkuDXSsfAjUaPwKVztNWR659gDlU6dSK63F
UKZb+l/ZHyxcSB8iaHbhNOmQgOOUKZ+3UdXbjFncTgVaFi8UpTX/zWmJYqKH+fHCL0rOx5H0foqN
zgHNBuslyg1GEAVMNv3wz5hTKohuoEcrDqVlACq+mNkNPDu9+cMCO8hNMWuSM1tsMg6O37he1yeZ
hnM9H86mvIKFgDkfnCOFyQBCyq2ODyptYYxJyV3SJlXoWxWGUg2lFgzAv4URqxSnbOeLl7h6Wz9Y
Bm1eWiGwFTkdjqFDqYiHyQSmCCK1FqN+I5aJ5wAt3cZfG5CHEPovFH8y9vVvnqoSM0/mlDWtAt0M
sBj/9Hzl0xeGWDggOcf/YVxcoAkbIjZa4767Dovo7RfNVW/Iee9ao6+wyCLtz9x14dWsNbSKRtN1
LQfUf7f+dE1zYPxKUEo+r5edVLqaOrCJ27jBoqyXEG7MjqpTL3dzwJ1tc3+oaTJPaMt+2pPVrxXp
seMGCWCMT3ABfVEt9eutacekZ58MFqkIdSxKI0KWN7GobF2ewn4ApBWm1aaNSRCKROE57fSrefm1
q9I6nYgQpKv7J2nMpVstZL/L+Qpm07GrQoEIvRLgF4+T/xYz5cS/TKP/dJkw+PqQ+8kASghHGIJu
R3E9iNN5csSz9P+VQMKXvO38bpYDVsh/LtPvVjKi237FSYHiqyPNvpnTSh9lu1090FyvxvkMU98T
2FeFhaQt90UjLq2fIE+vPIKKXvz+o6zziR0ntvTsCK/OtxTjejZ58BvNugk8hcV06APM0cOBsp6K
uzW4kzt9YMybNEHnqfabNhGRNvyCPoQIgtgmqA53bUGSwSOCoccU8RJlBQlEiugvccsMqoKE87qc
SMi5A/fLQD6f4uv1WvTcOTdJey05GeCDtMhIEQeiTsFJWRAf3CgQcBcIzDu+3hmnQVMQ2V6Bie0V
BS2RXbRAf2/DD7qjlGjid1nSrPBvKp1wGBRWjveOLJlm/t0Fv/4bIRxqrV4sQPgyGKYK4sqT/fPK
4jTogfLhjQtUcxfwtm/b8a2GhyW0NnovmplZeBsGHJSTY5pp1NN6MiwFyuGK5e5MxkwV7CgVUnRT
b0dMQ/cMNla3klbj00fQECwU1loVSTEB/fjZnj7VbzqVFmd5W6ancfa+0a1yLWrpnhjvMrvmoiBa
6JF5m2dlKQvPslg/Pm0dfRpR+aAmM8SJVc1izpGpSF6HCOrKtm68drzS4ZhlizyhVTnKW4EvWe2n
hPzwBfts5H5iTzQ2hl9XdY0W3yadpCRATpBjW5SB2CuyPRN6Zrj8SFSfsOab8ZdXoG6M3a2yQAhL
pffemBR/zy4wHS5zmgnwZ9jt3s+qv8/5QdSGY4XxTtZ9JImz1KYg9fRl5GaU8EFAlcGGsKYMGY9S
M/Hbv0X8D+vUq75LVO+bbwd+p8cI7GUD4+HQvgKOfc5CrLjJwD6JwZ0qJ01d9B6gESpaodJjK7bu
nu53A4VkmYs7rMKaRwJakbwX2wElESHo7NOPkmxe8YwNjIGQcW8VFtUCTpAOzljyIrTUxbbT22DR
1yaAECaaTvBr2XYR1+28JRXwSOxHUOudXFCnCaMrxrT+nU7m3izfoaunIL2aUTDafypRSR2Uvu/c
kSNs+pd2tY6SFetHHyFLwN94kFH45I1ca3WGGurNulFaQPcJc34i525wc4OF9DCPR1f8doZFK1+d
6JViakAmsaT9hMBWTdWOffJ7iETllwo5yyEXs2iJ/vTmh27hbUI1m3U7QOVdfw/R8Vc0HLMDUoE/
qjRn3GalRTYr4P3biM6lg9MJ8G0SbMKnno/0DoJnk5dKX9OqK/lDgA/M8qoYCLtfIYaFfkTOLjdU
tlIgVgV9g8zesBza7bzYMuUhAt2Ot1bBEY+M/GxHp1g4NiXnhDXqiXaIWwhzzKfN2FKJSFVKGDuV
hb/fts+BoI3gzamQV+8yKPWq2tKPVUan0klmyVjkE7isZ1FzWtnm7A8LSFdyvclo5zuI7NFHZm9e
HalhK6v5N28iXU1jqf2fm5CkIEToCyR74DVR2iAl9hW16HuDtGrETbceGR9nufny8EEsmEinb8jK
VW09AU43rRgA8iPSmWmO6OBfDwHsmNycUhfGOy87u4Z0RDvNzIyPF1s2dZI0WsGgV7/WxL1MtfCh
ObmbZOxBxf7qWgYFTNLyZX1irwS8f/JOWms4xF7rOIIWTbFKJ6l4eG8blyq2086uzSKX4aFvi1pi
SfZhGJvbgx9Enx4fYWFm/cAGcgy9Uxi6svXLrxkDTHgCOjI+2Ym6WgE7I27HZdmwvEoAtOuWTdZl
k17+nH4sIX95kEfBMQcQXwkefrLXyeQv3S87hwPCFaixaIqDs1qjnVLlrWBwIn4NkvIIEPHw3U8d
ljnwWlq4Pq1/qF6bZ5az0PBJoQS4xbh7ZFpGKLIcTYZg/3t6q8cFfrsz2rboyp8H+0C2lT7Ff+fg
xKbZe5VqO/4PQL3Q/36QcsiiYHXRBDikZO2fv3vx61eHsV+xq76aKxLBd3Jq4WIZpKQuMCYAO4mz
j31KaBoG5hj+7PtV1dW5SKz5RScH8LKIyTC8FXKLycqK4VMYIwXj80Q16aQR9YfKgYEKe3A3xjBP
VXOCTxp3F8fVtRyfeLAwMHsQQqtgaeNIh4DeWyrmR4sE2mGHWpyeD3McwrslL+7e2d5zgikWwkhC
JPAC5WPULTS67JtY5TqNyiZ26TfIsncoYYBxzqNNoDtWBEG3rcsgvraeOCPHZVHqJCPvznXNUa51
dfKeF7cEx8MPOCK6PcIWN6gD35FVKmUpxZTwTOYxnPgLSt0wwmITCFxJnA9J927C9NngjUE1lAVV
4Tzqnn0HMUZXvrNKayKbwkMYRpVBLqOXBUbwtaMjESrkaLTrMzPTvyT3gHD5nfwLWWoHsrfxFZKg
UkPNl7oYMkSJPoCa8/ugVSTIfIjwaGv2IwuGy2mpcFq9xGIc9fnHVRLWrYGTE0rAETlcZHzWQTRR
tlryqKcmk+ajFkV/Q6ji4tfrl8ahv/HoyTMJzdpmu1SDhQPGpxSpwaFFGn/tepvPOmVACq2SH9CJ
uc99tfsu5B5rQ1zeROTFKAWWkDsC+AC5DrxY2lArQaLlmihidRVK7MUUcL+OuIAihjwDlKXm9AB0
L/dMOP5PB0gWOmHk3bz2XHtDXc9ylgFiIF/YAIMAQeQPg8hekl6odRlZFwoShBNbLWUPTTW6N0dN
a2sUiv032yA0Q0QGOTzQRD+p/YLvPnMIa3CWk9qynzG4+IB853tmcMeMkw8hUmNjYz/AvI2rBP1f
g/C+tUEmTWA0BBi7v/yowrwcSc27QNtZpVDHktCJ4UBV81plrnBJSN1xJoupna5xp2peGUIadCpX
+SDD738SxQp63bmIuHUDXGkPnooKH6Fbbe+Y882Czqzbs+IsMUOZvHl9GrSIOQys2v7TRIr4fFrj
W1G6YJ7YdVok1Fokn5Ra5AO3yf0uJz9Xsn6yAsoYbgM5jaue2EE7rt/5hFtDZeko1oeL4RYlU3WJ
e1T6zdeO7x3aGWKTVcty8lfQbcKex+z0vFhWi33OP21HpxfWMDY3VC85xbf3DDfsTCx+7aEb9+TH
iY8DSSVBFV/xJWsR6vhJ235KtuhYejPr9cwaSQvsB9Y8K4m4DI6Y+xkYZgY0wDCnd7P7hbsv9ZlR
iexRMdhBdg1W/Xjrr6KxU06TYbKM6lumx4Y3HB+tLWWHlg6CfN2t1Iqi7kJU3zmXgR0uv8VXZnZS
lii8kuIWqovbbC1E/Q1g6ly83H54uDOx2ZBSwQZRgG4vQG18gYsMRQFVTaLmeOFk7KyKCnxXZ/Sr
0OjJSwqAL4TfuXYNMYqaOMAJ+BuH4W6ZSR7Wb9tFZRCdl4rh8HQ5tuhe2Lqh2/C1I5QzWAbbEyi2
AtvoGn5ziCosUCMbBDwfhs642ba4rTfVzdFSG2du5lDT/xA/pVyWWGa4d7+2Xx8od1TRRYyTDAxW
tDzK2kYz/i7JMNXaWD/CLjoNdBZbnKCbZeX/fYvDKI1c8cl2jANZTRaZawPDX93j8U7VXWjLiAAU
HerhCh9yZDhkQz6Sxb0MNuhJfhOrKt320zRl+EmidFvZ0mu4GyBtNoj5dktn+c+iRTmdtDoIOsMu
IxZx0+gEgdC33fEfLChM3jcGlHBseMiu8o5U7T2jNaqDLpmTCtTzdgNUp+Oye6t6Y1MHwQL5U1tE
cYHXeQtU33jKtJgkwvzgRORUi1XIhuhVmVf/xlibJMGbj9G66/zXxp2yhnQwHxU1qCIFEMJk3uEQ
N/xzkDnIxhlRIP5N2RlH2T83yFiczW52B58dL/q0Wik8TlX7mYbRTX/nIMedogJEUp0xol1VxZ+T
MuRAtTkkNL7AsXDcMhm0PFgaKYRB4wm659LXv6g7WQK3T3V9848z2CDL1XF1Ls8trUf4KltLo47p
vIjzgkrAVefwl6a0MoKGFc4rLozf6Xh46ejb/OdS0jdYrZ/Eyhe/MpdCHerMr+/bl20YLS9e3nzy
CbRbhKkOblfEYsDGxCLpVcS6IcAe/0RU+175pA5fJq0PVqL1lzjw1ObaWKjkfRUuKP9Rvk31fnFu
e4u99+9h0oUsU04Ql5yGmu1GdmXk2HbSzIyPmWvHHsGr+6iM73hJDWUud1n8JunMvqWW7+uWhqK6
0Cxg9va2FV2tgbOeYBkAyy12kuiLH5QUctQR8/lrhjtGxI8B7GI4klSjiGktsZPL40CJjL4nfcSz
htoIUkbUPfTxtvWhiFM5+1yF5kcT3x1AmK1UcqohE6qnG5itGh3+xE46JoSdSybJFjUorEB22pR3
8MrYRVcS/SlbECfbRaMp504Agih8fgAirlDZlXQDA9S5Zx3tFo1i9GDfxxcawvxVYoylPfEJ7zJ4
zEqOiY/sdSxsQ17aaj/NH1CI5UuiVNpUCF2NErJXsGCJPO1Xk2AbO7lglTJyCzKu/vDbMZRurWI/
JgnMPk4c4wHx3H1J08GSvpwj22OsgjewNrLbTKriQj9JF6s/eP9xu0Vi8xOdU2iTwh8IEi6KgNp5
w9gpHYr/ZbC+2npErKG6IZTq6F+unibR0uHeZ+Atk+NR55P07z3/3NwQxLFk7G2iHdOoIfVW10IX
f+kZFhz5IJCTMl5LMphuImKL2rCG3Ckn9eChy7XeIh+gEhFcccxusOukmGmhXXfSgw9nIRya7L3C
NYVbkTnEeI5Z9MCcG/XLJD0kBMXxlyLS5lMWFAmxdfls7X0sfg7nTtwIcDbZyE+V9716de52crhm
l/CGcRprZnTuNrG8H5tRfRDGhccwz7/sKqnPV8pk/yd19XBi24Wlpr1TTM+DNOoZyeazXES1UEvr
CA==
`protect end_protected

