

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XoDvqNcsUAMVrCepxGZ+692mBkX+rCE8HMYzKPm5R78cJ+RMc0dkNWWZsdClXOY6y1T5UuLnfOdJ
4pIk+MIfbA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GQd6VykDj7htiYnOl+4WVHQM4hKgz1J8Md5aI6kr8/Lamm+PnYCv/9ATHhzH1x3ZwU/+Hk75nShM
Z/fTah2o7SNlXBmxO/TZV+Cu1NdyZPM9aMjSfxhjbc4DdKhbt2eR/JXlXgPN+qqN+l8aDRz6dW1r
rhTiAjUos5V3YtoS0kE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1H8fvXKZG1QF+UJtGmRK0CnD8bm/+01l6RcgU14qYFFE8GVuJpGQyW5h972p3ANLjy1WRtjYQ4xM
/dkbNa4PXjLXaYaHj221vfSd3lB0MAvfi3uUVJSvclNp9cIhjsynHt6eX7sY3mGpxNDMKipfks7Y
7QsvE6SpbzMkIaxn/W/Og06vrJaRobnXPbk5O8bulSLgRIfqtOFawh2LDbI1+cySFds9EMjhPXGY
R3cSwZrw9voRIz0AJIAvvOBrLoxc5eVp/j0gskNHjRbPo5Gkm/B0oz1Ia6kiZiwtS5XXf5fYsvSq
8ip/JtlfeTs2FRpXweWaPr5rFOg0LxkGg0mLCA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7F7hPxr1ObCyOsY3iC3Phcz4OOcedLcCp9ggSn92l+/8vc/8WokvA1XgYsChaRHJl3lXf2X6jfk
OU2I7E3QgZVgyd5+syjWVqouw27C41FFBeCuGD1GtzyBYnFEqdtK4Wi9fPab76EJM+QSrUTFTxOM
vNsxaERzJOCdVgQoGH4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DAf8RFZxkL4Com/8UijiDJflLxIdfhDldD1zcH1XeixMo5g8/n+Yg5p6ecx6wthzScLrbvkfxjSo
INrqjZhuOy8JD1hgSySspkuAnlB/pYzsB41QYrTQXDdhODLQLAYA4QNlYnc0Hld5QRA0QsNa7b9I
jitn7EoP2gA5KtAm5w8Y3SJ5GziR/wWC7+Oq7vo7hHrOsipiX4kUa9vhXNaEzGvrcPOJN0YgaqRR
HJt/OxiJdqU+tEWkUefOFMVnQWevf91iZ/Fb0oG88z41wfeJt8eTwCR6ZrUTPInU5uj9Frdns/GT
RmMrsalABVuwLraRXdip/IKnMD1dw9K3eH9MHA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94464)
`protect data_block
HmbC93q4RDjfIINaCQRDMVLVTN5X0/BHcrd7DV1cG6Slcm/ChRPKvgsZNXJNR5ZAzBt3BMLR/lU7
89UrmJZSm2oDwornAZk96HotV8HOc+LPi7a9qg8ZEhMDlSRsVXIwTXLqJMW8rMq8BJ9LgyPDaKva
b0ONjdR59lCeGEln9J8iRuXh7qAXgOoDyUP844GPsA84Tssn1VqmY6wkcodXke4WnFOcEC6C1jB2
JnKhnBz4NtnU8jFP3sEHfQYkxTF1AvBGKdFSG5EO4vNwkFzkyKsSsj5k0qobzi8fMocTpdj5X1T7
4KZrn+YVdRaQB6b7LbS2pih7RYgwdeC/hVxqaldtkRF33eYH70kGXdhfoxYCvlMJrVFqsdtzrRH+
pelWhuGprEKIdB3hQPj0d4+IXPKQgN+xKKtZv8Wo6D4GbCW3euVj+8DLxGPRpMA9D8o/uHR5hUxc
r4QxoE9+FBvTC/z+aehoE8ypDmYx/8dyqEUryxOBQY1elTBFCF4OqsWgxaR1ttPowLLtchrV0sWq
H72F9ZQqlfZDvxSvETcl+2CLQMd/1gMnn0yULbn+UAeR/AN9/UmRjPC96+P4ibqjlaHqn5vay2Xe
Yb0lvwApEalg2rwx/OQNMXS6O6LudkiXi7PnXI0pnp3H3kVoiORScmRBWx8e2GgedRq+sMPii1+Q
BYYW3TNnO8Wp/2hti0jwpALugQHMWXHfWaHcoa5Mf04M8egsue2qqm+rJXhkAYl1QfWm6hvTMVSC
4Ud9wolHAQokZz2rYmakEa+7x4A4BZlxlugJniDvWH17yPJrb+fiG4P+H/A3UmuMTap2wqYBPe/l
33geCnbsi3wkvrBJuB6suJf5zol+rAOYNQNkGann7kQPkFaJsUQCiROASIKGkhwfv2z3usszS2So
fDHR8RGDKhekF4OTjea47l2JRWBKVIU6V4x5/vvcC5w2HJKISmjtkhlZJ4wcocxb2qPJxB2Tk/5i
i8zHqZr95dsZJY3VKxg2PZGrnXIAlapIUQ6KMq9veoIy5S2yiX/1c2lkAAfB3A234ceCrjTVCgxi
vKJpg2T7SAlsobSax0aRIX+akLX89x2+GGO+0a5tBLwsYr/LArZOcMEZuuJKcA4MqxnngSgWivE6
1E1Pk7Uj0blXCWsRjmc+9a9rK02QzeufFv3V/YZtx/5XiytJV/28EzwA7HgWsgf0kL4joAdFwgDA
xFC1sJ/L4dDsm5vEzrqLp8DKSLcDiB0uM9IKcFCsN79mTE1LFgBE+YK8siNUuVc3JZg4qzqv2xX0
Je9haUWdqZ62b0tN3VNeN60MynlY8YYGES1J9xUGc3kkbuis/aPY+p13Rg+quFZ2CJMMFi2eD5pF
U4/xL8tlXLQS6xdCFjmzX17gWwPMQoEd+kEFVYcVumrO+Sb1nAWqITqlHIo+tL8rnLJlEhQnh6Je
5FIokrxe7ECkbyiCqK1vtAlR6CNXuuv6bkHqpahykCULl9JfUdfcfyjDJI95ySpZGx2OBPz6Qri2
qQ+9xGrCcZOsPayP3rIyPoe9d4tzrvxNj9Hw/f8h5uoV+ieW3sAk4voW0EIToTZ78D2h1i9+r9Fc
z2q9hZh+R9Bw/AciUoy68ykmEA0Bkzhb3CDq4E1HikjxkJJqUlC2Az0vsoImHxRKwW3Q3HzP9363
dXQV8azZwY7M/YmDjRzqpfgt1e1Cn5T2Y36eKV6uQ+zlk+bvpZMeW1X8irGCSy5Wj70lmD3X4d79
OS9+5QnuIHXpFx6JKt64BwJrndDToYwtoUysOiMx241JB5dAvj8K03H8VIxQ0n1Kzmd0t9M1eMY+
jqBbtvOFULSXc1Bk5k6gTZ3ciMJsQaiPNfldLd0cmLm06FdRPDFKOLt4iRdtlw1VdQO7rBsyBKuJ
1HalCriYZkMcqhI7K/W2eVb+UymhefAFgA90G9ek4q78X8QCJUpVVf/YhSChzPNxbnbxO1wpkQWw
THGpQr762cC9SxmDsM48Bnzpis0fpBt8N1UGQDyKkRinE/CqFj8QGM5cp1b+Xo1lzf2txut88frn
bjdzgmvrLQH5AwDajjTn/AxFWen1luI8P0ar6ncPOSHEC9amH/3ZlhOTGRIrbtFKCJmZazGPIhs0
9bEkgS4FVP3hid1zUzpV09gbHUArUzm+QPyJG3vaFtAkCmiHnGUOSOlXUWU3VoMtcNRzUy0nMVof
AaFNLVw+K7/efCIAqjbmYA/WlfohEKmEG1zwEzl4IzktoStD2/Lh+UhKfRu69/4eCY6HRWknNjeO
BT/DyWJ7OMeZJTxTJ8SOCP8zQcLrqVoJjF23BeowJ+LwV9IJCZBnLp51p9DQNtW3FylYP5QVkWVg
EcPJ/K67ykw2D1RdkN0enlY1HzhEI1p4sODdLzI64M6jcj33oCrh1rV7MGigPbMMpgi4dKeE7Uqs
xsG7z6ZHT8IHJBW0bCJ6M9icY8HYwX36nNcGKo2rjCbmZeDvr+n/WunEIZYC/PhbmQp4m26H8atl
HmLJlWkTeQOb4UIXDNHZE13cqhu3DS8MtxYije2PwjcSf+8uV1Rp4qRipddjX7L5a9h8y3h2oHrB
kZv7zU4kvB4C8YfluGHIlJtvgiXCOhRr5rmcXcyz1YkQsxFLmEx1o3GgEcUa1RlX7GS3+8zoaLEJ
W9EOtuZICG9cHoEadXDE92qHenszcBC49GBhiEBfbzYZph5kuDy6vewJ+dMWiWkAqNtSE1qhmQtf
FEi6aGZE6HyRAK8298NyTphBCoZ0RdEueXG5JoyNfYYT2PbNathCs+qnoNTCR6IPsYWYpUgwa9Fx
FBIXr081BoNN4FdK83kM0+c/0ztzvJkLmsOynN3XO0d732lfRW0H+bq3EDvjDQMn1wU71u74tjTs
PfB0oqKUSoxzkWrVpU9r1qRghvFwIyTvXJ3LEUwxfikoZ3UUi8z/KHGdMTzj5M4IyEcmPp+CqIcO
X3z9S0RvHJgog8etHUI4P38d55jcglITjkyKISmC39cXbErbWvjzgz/clNYVm0C/5HSoBBUpnOIw
i2pc4++OqvGQrf0G4I8NSMdTv1bsuvBxltnCW5znjtUDbVzIbRCtGeBCRkT6MLbvUhcEbZdd87wR
AY6y5AV/UCQBXtayDQVWsoMIUnRSLjurXnORO49nHWnZA+Iwlx8MpGTfdxs9n6+u+3NvKMQZn/6z
WSPMdJ24CxkZpgNOKJ7C2iDghv+EbCYZ7Y9FAV/NCY8O4G4XbyTSA16zDTCPx8iiD9zrtAcIsxRN
ha+CKCz5vtI2tK6d56J6kwVjqmwffRbNUIius9X+P/0uroILQJiq1r5QuFrEvCF7u423/hKFBtSz
OMJmrxhhIcQ5+Eb9FWSD0Tf4l3CfnKdrY3RdMGSIHHOj33CqZAtPMmM21jOOwWojLEIzbOKm7lvE
l2uUCDsOxQ32dvGc3p80mEiFB5uNimNyl98hFGWACjRjiAZ9Eh1h0kIe4av5eFrxx/4Uarc0TZOT
biKpl2WKhgR6Aaow/dZOwAv4wnAXbnqn2y+jHZhPAJ7NqACUiBGJM+UNM2xC6r8OUD9k7LZ8Sgzv
ZdrDOA7hV0JXvcNcnLynnPkVUb/PLfRk2ryU8AZpY6kA+oCC5C0yKKBZkEWZDMha+d3fgyWBrEv8
r1A+ySwwIx9eZe8uYZbDlPpELpqKTfXOwkW+w/Yx9vxTK66Q7VbOjjP9BFHEaR5K/NiGAWSMqsaG
Rn130HKkgGp8KF/fGHNx6HGzSnDJ/TFlwLEhGA3bS/wDK+Er2bWdXJ1y6jL9Ah+dJNz55Zm54xgi
IxsmtjoQpDta7MFo6vtDxXjcbNsMmTSwY+2h2fNKeBG+TjY/YaOwyQAx0Cass2uYjs+AkVCDG7z3
y68YHv6cnHfcWpZxogmxXXgLMNmT78bVPoqyewFMNcNwB8kfn9WF+MXxvcb5HyqXh7mN4DCAQCDj
RqptzVwK5Yf+ngzP08symN40VQu1tP7xZDyzZyUhZiE1LA/Lt07gyIlg07rFufYLKs/I+jt66KtX
dMHx5upN7e6HdYGDrTXWR4CGfc+NuTteBAKPXjHodWgFLuKS2yIn5xToTkbTTl63o/urfvKfVLOr
PGa9Ypn8s0Ha0i6P2ZOSwJHR0EYwKFVNYqCWWRiGlhzKBN7aNH9gjGkALPGP2WzC1geYhhJk5rQY
afYjEWTwKav0VB/NGzDGwryupgIdz1Zxaw/PBuK1bO7qNrCQfLsNEVJmbG8dxTH+3C8LefjmWm+w
EtO+u6wpvzIQqEr7D7/2hrKe9txmXf3LJxxtVdWLNK/7np7Nz7tzXV42C/k6MFcd9Dp0r8Yrpm/O
D7baviLsCAQ3iQnSoZp43rzkw7kPGsNuJahscbgi93xpH+NpSrv/G8BML0FecwjGZjn74bhMJ8dp
dDH2tD6u/IieWcdVLsHSzoWiyxOiF9e0w25y5HtZkkzJVeoZylqC8JM0vPyo41ABIBsPLuk2Xtmp
V5Ms0WWx45mGhmS+cUMevsn3AiJMxYaoRBVt6U7jb2TIxXJIe/UVku7A/wV2awd2cFMDASS3IbCT
SMtpiUMyUQDKVDVWQX3YnfnKkYlQ/1wqqa3eCs5QVFSarNqHZFM9FXFjnpqkegKLoT3/D3BzO8VA
j/eKuFlBrKbmxcz9gBe4UAe+lyas+8XSXqFIOCUJFGiuYe1KadG9s4T1Vi6l+L76cRXJQJQnLlE2
2kTUVqP6UZHE2t92mA2Dx8cSZL0dqjbv/kN8kBGuwTVL/RTdN45ABk1JLP00Dv5GpQd0Q7YZFr+z
3GaM4PKgF3aP3tKdOZ2MNFmISl2GfbEmbTk3XBFwIgXTpPGXKv2YMByvQEcxspOGN5N18/JsS/W2
VZK0MmKZQWSRrOeJ4iTW1jbj0wBwKmQOY0pSRkoyXXuUah6XqCQz5LIJHwFZ6U5qg8KbJxsukNyz
6vkfp3oZwPu3RNp7RdezSH12cMa9QFJ+ZH4YMRf91N8anvs7S9uFlZGMJActszmapcKGvWE6aCka
cRSLsDKCKeSOnGaJTJC6jQRiFFxesa2C2JPmtm5e2BxyplqOFSk1zWSDKyMHkmsCnPtHpt3dvqOX
D+dwuSZhpTP6HG7f48nalgN2TqVpycoITXHETE88YyipNrFtpfaFj0dHWUCHcrCX8R4MquiGp3pY
Q5r8o70M2xxm6xV5kFZ7p5mlBmp8aMni2jaZO7L7InZYTKXcZHufLCD2DZtNqIh4ZtVW6cH+dv/Z
D+9pt58NQfP09Bx6LcvbaBDV0qSeySbnFyXcC8E5JsAumkOWw2/iAP4vOhZvh2H7UAkD07aluWh2
Em+IKtYUgkUo+F6QunXupEn6vbHs93v4v7HTJzajQRrg78S90HMMtzR26vM1fMaoRuit1M9/mIND
aqAlKLBEQTtMOnDkTmvv0bPcyPK1Fw9viVrxhP6SeCe671JVRK7HGRzCe0Qbe2qAmoPwoOPSHWin
2XWGdTmpfUMIJy9i0GJO7eE/x8UGrR3Hdw3TMldWDZkXvpbXbko+8QEqefrGrX3i7Os0IckLuDTp
kEQEXmsdcxvNjbb4pIzH5rLCrezGktdojkVtCWlFvEHIa1vgkC1TcHP4zBCRirGHUClm8sxSvhZH
ANI9tIH3S3iOBlx9gmkrbn5k3qN7KXjVbi+we2iY3Qpost7NJ9SnuZVR6OC7l+r6k2WmBTS1ACzw
Xg8PTxHPfkh6p6bfkapcyJTVZnmJHo0edWo8WnDt0qjxb0ltIo3g4miOtBVPJld/DgD/+Z2NVbFb
j70KfPkEPg15S0SrVq7NhptmnlBMozyLZar3PdLsCwQY2NEwXXvTMiAhjSS1Zv/my0kC39n0JdtP
ZTcmSFf/n3z9Xh22Uz3IStEo7JoU/glh8i9+V+rwhakByoV+BdcWm24xFFSoVu56B9pkErvN4k9q
gzpxa1uEqmgAX41vfLZdFM10aT4m25J5BvUIl1Qiib/BZJZnlGaj+3htdzIoxesFnPQKkQFnqrQw
Ajq4gUpsXWV0SgG2I2rRuHsrzKGPo6OH9BnwOLQika4ED0gMNArfo2UJRxZRh6zdvpNjQcxfoGBn
t03KuROQUMReJynHxxkHPnZViBEHb9cRFykxiJjYrdlTQqvRHpgjdD18nUXYt9zmup0r6CQ9LGYb
EcUMS+3KMPkEFwyw/yOW02F+Ah1Ck5tq0G8WTDfcHB7dUdxa6yYVPOkIQxDkM9LAfyKjLW5CFhH8
MIxoZjyzq5n7exwccpredptZXYgtPZj1dErmQXhZUBZ73aBntk9S89jixiSvPjXuKevgp8TntGSs
zzHHpnzcu93rjIoNYTtYSC/pt9YTx9kwkYbunI9Nl/rfTyeHVFqJ5787ptmalhk+pks5Z14Z217R
PMGUEYIkfkU5B8+6Zt8Wn7advfBKU7/iMPpGve++bEpOM9PlNKSCpXJGMdQjlrFGuEc629uIbZQQ
sxjHsNa8WzZmoigqAQDQKtsrswX2baXJ9hG35Tn46KjvowHVaLbfKjeo+M6dfGGrOdIyvRz9GUni
/7TdECbroP1mEa3UP855ZHa1yTmwScvT9df5YMBeSyKkFn/GK8NtZ0ZvC0Fhpp2lkVTC1/ryPY0z
Dz+m2QGCGTikPXbYekQZTLEiux88Dgybic1a2AZEEQWsCU+21fYcXvCQbgrjKR/HZIZIEv4KhpV/
hqojmIOSMFT3Oq7AVNLtaK4QqkVyJIMg28ECGzztjUDYgSjjeD1gPPLwPrLk2YViFapNzDlMrSOP
CkhGq/0+xyfoLojuyHlk3aFepU/juCUH8/kLtVxXvVIkVYXl7YEMQr5Wdf56g5S2amqxiW3olUkE
mSad5yOK65jiX1qOzDcJz/oiSVLP9DAgFRF84AN4NBn4G9WbrlCVrGlqMsGgt9C+hEMGgtzLQ8Z5
hwa5bFyGVCJHI3PAfkAWVs2RNz6vssrRJffEIomtArheXgyH6u9I3QYybC3s78SR0lHGIVqRAvaS
IJonzmRgIVnlarYNU5JjBezIkcmC4VkRlSeWLkmqfGhsNOTPXs22jDzqE578HAYkdjiADcYU/HoJ
m7AK9Y0HjaccAVqKKATKl827dHqmKEmw9st9lCZb4ZzXRDussXcut3Wga4Sb53UXlSTVWO0JeshZ
iPGfNcB8wgj7vSOs4RWHlPXEQDSnSgqaZkiYlzl8f3aKa9r7m9LTQLD5ymCKFGHZOOPuRrEBifB1
rfYqyR07t9nCF0RXQBUJW3n7SvYXISjzhnMopaqK8UGeyJtoczqbekn1eJ4GWa5Jgq/Qz9UPEwyC
39rXlGce4DaXaTnzEoe6WeDwuaNK/vTrNUkQgReLgGVj7IwRFcLBe9YhNGgnE9Jj55g2cqRPMKmT
UamI22HDsuA+hlr4cSsULjpCPY9ba1TcQ+oYPhoTRAeNvdUzK4TI4C0juekrQb3wJAsygLpHm44r
teUGvKqQDHRzVJOq29FdMc77A4wBMP3v1IEpDOO0SE7SdIxYXy5Ab2o7g5fc7pBmWgiLsJ90u7Hq
l1ocQFK4nFP1BITcEzRIge5S5yQo7ppfcXMVjYjWVha9zdjC4GrObBlU9IqxdKD0VGHQhkWv5EhH
N4U9AFNOc9ypcianF/7xyjnuG62Zt4vzqotJeiLUiQPGVMbqFtwMgEHEy3xMeDi4pCOSuP8kD88S
E1q2l5KTgL+7XlzU4j75lmH7y5w4subJ6CDb7ySeJ9V97cPvmRoAoKNNYZUDytJAbbN3KAecDdef
SD1rEUjv19Ac2G1mXSmgtyN43FUgMLu1ifw4GrQSHpHkGzKi4qMWmWFIvuHZTNKR91ZNSNBc+yuE
m0md4CetQwFcyUid7xsLclxSDJClRt8b165HUMYzBTA0hdLBue7b98PfnVTb9kFkb5UghMSQPKms
jZQGBtzbCrzUKQhK/DinmU6QwIV4h1LD3G4bSH5bZz53O2q+3uW+v53tqcJFUsmONXSmzWdal9Y1
K7xPubM7tpnbia3c9vlMKmKTsk81A/mvKHJXsPdNVFN7umI1XZlwNh/xxyI0qt5XFOcBhM4qx9sy
GEkBdplvmyM3JOUOmniF+nXepqRtwtreDXbNF3Vh8kf+zZNfY78iufcrE8UrkUVpsT/L41wkZNZv
/IRRy58HOgqegoNUq8IHVqR2nspbOJ5sHtkq1k7/kYaMID0KvTGDxfNGewgTDulDtH+JtbAG0XKW
pbuV/sSs4r41KaPQvFh1uHPi1tYZ3YZS70OzBJbkhz2KhPnX7O4iQRrzJYYLAP6LwJMTNaaiTXyF
MPYC1JrLOF/CqI4GruYEmMRgPYJCfrWLB7J94k37aLUITxLOxdZtb5eMml/+SXSFp667RiP46KdO
y/68ObT/ky+b0pMlgkSLExI+GmiSeaBnybJnpubYCg42jZra0HCYvdPSz0LW5A8IpCj0N0CP2nE4
9twU+5eO2lIhkAZQx9BrwFJ1xkjlaq1CfgHyEz+odFy/aD7sTvh3xmtd7OL1+AfCUfSD+PVY53xy
aMyRTNCo0/VmstjkbB9CKLfkcaPz/c/7FvEFrzPgdq5Jvb9Yonq0YBliGoeL6ABg5tvwtaiQKHE9
Lj7NPLYsrV2HCKC1Y9z7q7mT4UYBUtEtht3jp6705xP9WxSt2ZmKCRIxKe8dcLrFWN2I41zlvksw
UqLCjoZu7YsdaZucC14L3IUbiwz484vlDjoxWLTDmWeDq59Kt6Twr2SMGBgN44qMIf0pvAJyk49W
9bu7IFwfr2luNyIvYoMXriaZp8gTTYuj2KzWhap7N0Mm6Vcj26Vwd7leH929Yl1Cq8bDfnyaboI7
o7hNc0Cyl1J13DNAl0urBeNScKxrBc1fhpelp/veQr4DOgCUK1wfg/ESreMFwGlhe6uYj9cn2nIh
nv1NenAQqGPcFrpFLiKK5/90Ceg+p2YxL57iznOM/MK26C1VsFF5e93aWDquFpz/qIXbfrHocR8G
cLojOIeibFVvpZk2JFk9RJwBa/m20TAoF6oRX+eZ5ZKUTwzBD7xA97tE/K99Idc3YG3I+Br9sseK
BXzRNRzmdo3DMGO2h/SOdPV+N0ksThscUE2fD+piNNKh6k4heBHz43gSvZx68QxQYFJyO7yAxtrk
uywFX/zR8TKy1VCirOYn57KvJmtNNWphvTHTQ66buKDLo+C14h7yoX9juEknyh7IIIZisbVghdgK
Nbg597l6pgrf/GtFd11W6Xvztsa4jIBs36u1xQ3hlA01ik2Yfms6EJWTPMe2x01WNqn9MLmzWc6U
CLyYQ1sJiKOEB1KisFJ7hE0W7nBTnjXTUdWeq8KllWkzfi9oLBloNhWsrMuwN6nQgHGbWy1tYvwD
L6SFea+cNHlsum623cPUmXES9fq1IAUbYjgbRNLjedXIiR0yzdBnRa8R+5t555xp7ed+1IZdGVIz
eWuf9pIylMxf56WD7U3ZwZvp/r0ahVktT1Mu267fpKGkUXyeLo/ZwSZhpp7EllbcNaTdTmYcp66z
3OrWRCNZ84BvLrUa2xoNF2IJ5DzMe8TE3EZs7L+5SpN4xXUTLKh60mHsf0DCMjX6AySDTDX5BQZd
iXOqTvrNdJxJ+/WPlu0BvBtTxjoQWfCr/om0/f2TU8GuOVA7Zj3uMcwa/cScKYSQ1emgcxuqEBQ+
oeTrbENz6voyX+IsBwUprK9MoAqQFW20Bbi8FcdmiABklZcm3OBqoxpSkgkJhmxMdMfFFeTx0+H9
UGjwm8me4Ni9LPo2i3u0z9gqHF626HLZZzS3emDpLrn6S95Oa5X4Hjln18RY5NyTgAZOxZdvOaEZ
h3B80dIRpZPg7zq5g8nECBg1BsP8alyR0WSi1RAyPCUrQ8xaASeDrn+f3ZCoMl3+ko986c/hKBFy
XHmfP6WDd6LSNv0P7TDyPPci2NR2+g/7wZ6ERgi1wmCi1tYRAQ7n/+ijckzjNSfXBmsD/JZradFX
SBpMYDT70ZiXAbUmF3EhP31dP2xskAUfBhmwgYn/U/5BPjyPoR1/udkKVfRf/sEeMSy8s4BsDFkr
dFO6LHAejiGFcp2o25ywTIfJT7KmQAl/DusiH99ZBVoUsD1+3Rq6vcAq6zYRuELUmZJFcZYCqTPb
h94HRDhpMcwIAdPJ4+Z8TL7Pyvcgp5xgJlLvVDc+Llek5gdX+bncldkxg07onNdVTBJsQwIzB/i3
kzxluqf9sE98q4jbyu2xbFBNkWXbKZmK3Cv6Js4QpO3m7++AznynQ384p5yGNNW3f2RL9AZTKJQA
umRlnbBUPl0/M3gXyNt4nd0zPc/3G/pOU+AoaweCTSuwtIuzf3LUse12duorSNLo2vRZw1kWABT9
B2ooGVv1t/FgbfeyduPkO5tA4E8Q57fIsV23bVZWwKSOaBxyE975Ib930m9R2ScxBlREV/ae1Gl9
jdpMfzPDOTTntVh7GA6zc4zFFbjc9uFjPkDTTIfUegg/X6JaJoGN9F+siTgkxYdsdElFofzt0au8
knRjwUGzI5lXsYvV1UlE5MdM4Ncd/GTi0AqvGAutec7X8dylHLeKZf/Ede2hF/yK5GGphZi22Vsd
iAiX9ZxwONbFuq9F66PBEz+s3p8Dcw2AFmPzJ+zb8gHQrkCUg1JPa8o3jyT6qxZqzTXKoT7rQPCd
lyzMT04v+aBbc81CMHWr1PdSVA97BFIUcE+BtJ3AAPtR6pyyVrvldgkQHDJaKaXbFXfkE8FPj9/j
MKfV/LISV+BT6vWd0vK9oOZ6v5Zb/Ld2yyIZXJfJ2kY8KNjlJG0yfxUFh2EpA35Qrsd+sZUKGVzz
w3F7hS7XEGBTSZ6YvDj+NeZhQ31wLwprbdcNeZ7dZf6DIx1n8F57ipSGx5R2whTfKY2T3DKS+WT9
nfYgINupgaTygDT74uuaH1HFIf0oj8GQMc9H0XOWQ1WY3Fy0mUF45j8QuCTbVzAnDfd+uzZstjh5
1LRO/sDdhjuBSoE0XJXU8Bfkjl9a03JPtQuahRik4h/vvMcpwmzl9RrAwIQ3vLfKIGlZGxvBM1qW
s1iK+e/EQ+CsMjCPq/CGRjfTlhm3m4DXc5xJXjq5zlLjx0SALxOkP8olNFRIpuoT4z3Vse70suVI
d18VlXEGS1td9JQpdbwbrhFa9Og/ezncq11ReILFDZ5J/3DvCkrrUTnD6U2ahiewvbKu1Mcc4z05
KHKsZDpwD+QjFUfuXPdWjhcfzsEzqZJmV8rAVgzFRGunUcR9PedX9xHjxj9pK1YkO3Qnvz0bsPHd
xbTt7VsUoEYctKLaaBGAIDePpWCzNgyALzwdj7ttOM4RPomFOemQW9RcFmKdZD5uBe7EFNiEi5Lc
6QHpnPAmVF33rSO4geyk7JJVDELH6rKCVkZkfNNc52ZpUB7WBSyLX7AkqaK7orGifAezqE81AGQw
PY1Qly4KM9Ci2mIvHdl5vK2RTHYetF+6qE+4s9f43obxuI1sHKpOz7167LqaNyE+EzYE7oYzQg6t
HITJnUJK6re6dCGI3l9jQ/Vm0/uSgC0PV3m2x5qt0K8FJzNNgAxc+MBB91QuGB99OIebZjxV3o77
2/S/m7q9PG14qDoYmjhfZ6sOmGjJk2uTUa1pMnN8+CIdGQY7MsrEGeUjOq30n/wQql3oFf9sipaK
bEkJ+5jwggel8ozRjPF5LJoXjatX36+HQOCHpNphhx/gu0Kk2DwoPJUV3OcEfCk272DZ+f+nWIBZ
vjikp6HCOs12gDGyjTjVhSUjDuvd1C0K/5zfpIywYGAwgxrxjBZI8ElnfH/TSu0PQ+Ie0GGayXSY
ulM+diR5JVr7vQHT8+vgv01X0362ARapDrmOiYaz02KgvCAwayVr1FwGrmoENAXoQDf/DgJy33xj
Q7zPvKkidrEbI3ubIPmhVR0i1toiZrb6D9AfEk5mNaa/4hTYnUPg4Jr9RZTcJIfdv4qzVcxZOUvy
pQDdluOMl533NNnjA3gpCGCC5vuJU4rltxC/aMrg8Jho5mVWvHt7OeNdIIvikBOONK7jN4UFDdgy
pszzRBEV20UHUIbUOBKiAHOS5pKG1TwdCoIUs3NQsS6soW5M3/3MKoePvP6uwaARQBoq9N/YVKsz
FJYKI/ySw+kByxPSVP4pRIDWbHKu3Sj1hrho80HCzPudkee9WT/DagQ6PGR6uKg7hQpDWf0vEfLH
AxyJgcPZmw3JZh2i87wmdkjSjRkTgxwuO0uUQoh3ACdBvGBG3Uv36FJZgWe3SqXSNw0fyvMxerdx
MCz4+EBC7779ij6gMgIUc4AUeL84a3gFRLZOhl5Si/dOVyEW6lXOvNL0aJhNn7bhYKo1jCtiaCWU
VbSLVC5Sl3rwy/D70MgvPlpxR1y2JBXoYfZUshvKO4OlBy9EZuzmivEoueu7lPVnZMldY5OY8dtY
Cuz6ZOeEkU+XdKfLcd5hh2Ir7tfXraRuJO1tuYM3qwaJhdHHuUHfpl9QZLz8a5xPMHUf/XDlktxm
qbxRnY7rMiAEdUGVel0QKXJli1xPvD2xsOu2VMypwbvUdvHIxpMghEezfLIZ4gEpkS2b3srE7D5W
qh7K1ODZGqJdJoHjMPh+m3BNWrifJVSHNIaZBWxyMXhRZ4IP3k42d4jkhIlBEYMs8LEEoJ6Oi6WP
rO55y6IuFOY4RhcWZwrXGPctls+YRrQwOdkDSNRBvVX340nx4LU2oE9HrRounZ76LtQy3V3Nid/C
JnOsi+N09x9Z+dqYFet5z5nf0NwQraHGaPNzEBYyiccBhh09CFRqomRHno47pWTuwzNKWxOVsAYn
DGRIslZXpCDnGbaN9lkS6d5IxyluAw/lVz6bW+p1bIJqw6p5Hj+I4FOQFVbG1FlDBmF8D6+mlfkt
hNeHQqEae/4U79JEf1wtOTRI+ZzliiKxR236FD0eJ4SNENxGPYTF3fLt7WYtA63JzHKDf1LJQLrz
IVyYWu3WqcRJJqUKzvD5lq0+8f7fvnEiNC4bFdWN4kOj1aYA4DC9cbyQr6APqDh4UtSi59DNdgjX
z0wZfG1D1I3JkwO2JE0+kxYE90D59LSTqW2wA1JEUhMgOTprsFPdFTHvu/GmWSn+yYdhn/wxkwqH
8KVRBveewn8HXBJHoBS+e4VxiL2oZqVmiWfdA9cOUWX0R0anW/RfQODfM9JVrAlLYcNxtjxy+RFL
FiBs5fkzG9ypiydCNXW1GqqJDZGZg6fiTiIa6TimALDu+r5JXNDWcNHG6GwkXOVmHhQZHClme5Y8
ViTimLNwdJARIM3qYuCYA0lN7fSTyBMlvHrHhbiqMJZ/hhu3v9BM18gWRRJLMemt5IPBHbYe9xbs
aNQvV/pvvlfGJUHsjFgIExGMSPWYVpkrTKhxQX+36RQDaTGY/PM2rG0FW2IHLXHQAw7iiH2aMSYx
821XJbN00fW8+NR+haabslKGuXbdkZegvU1OiEFbE/wC1FHALgyjiw4q8piEDsd5tO1Vd4sfrZEn
alp9QrZmdusqZVxLDk8767udfxhdKOCiJfs6RD7wiMNFG64CCKuVGdMNCcrUf6SC4MetX9y79Uaf
68VnfOgIfzmaLJse9/j9nL16trJNK+SVc8oVmwsINJJDBBqfOyfvCQ8zT89l8XWo1TU0pPUJM4z9
0urb/LpEXwFDbgYeFxwsywu9OKFvPAWFEaVBqou8Cjb2KXxgoV0cZeauDDRIc61CyFDl0aIYPWYc
HlOMtolUCg0BeLoe0QJdlQ61FMlawCSEc9Y+GeuCHjRDdirEt3u+m9A5xUS3wHEx0fsz0W0r3lys
9eKPtLd7VW2lj3HGQjlXFH7waXoExd1t2BMMaH6fDTfZ5BMlshoz+xw5ZEfBJYuJalEWjfAP3uGa
ru8Ko2CrmtAvLjokEn5LfL/Bhe6W8sIAbnlFZigL7cNQNwgx12UVoOVQKabL4ouayvVzeKZCgnCB
5w/VJ/rQ7BUR55BKtfuIRsb3igNpM/AF6ltyLJFtactlECNqihsfWksFfJTPBsVzXidbXiS/LNwi
a90k4gxhr1Gmwu2jZkR3VClRvF0iB96Hu/3G7ZfFJ6LbHcxTdlRLeFxGZlYYbo0pnaxoZNL3+Dag
HBV2qbLExOzZ19pBz0Z/SztRfvZMvvRKjnZEipKwEhyfHN+3di50Q4VSTV4+5fdzIaVfCqMetehJ
OgUny3yjnH4gPu4DbR9q17bXVDT/I+xTuDVUdzFaRZiJxYEOZNsb+wU+Xr4Dsma+byjOnlZWs5aK
PwkU0fJEbs2Qx3TxBM0gUIPXxWT5K1clVdaFtEwaDD1wF5v4qEdcWPMSUlpZ+NYtQ51okVGbIrQO
n9J9cdvCCl7x+7s4lhPwX1LMYilhwYGjcQ2lErnYCupAXNkdsYxiXEroGcvbEtwVxBHaEBVeLL8J
2dxX10bbLCzsQiujjB9s/G5sUFSI4LmgWme4N8+KO692DiMZSu8UIZs0dNhyKVkvDDuZq+L1Cwat
QGgxGEY1Vamcps60eGSrhlKQIuS9mO0Jqz61xjOSeOBxh+jIHLgDgZXTkiu9llKz0Gt6q9GMmEP/
4nfD0BdrmPbmk//D16oc27gS+yFHEKF6skKJd9X1KMdS3y7sRKREjcbGgYFuhslKdQf3jQ3fEhl3
i8g8KdBOVIy0nEl8qRCEO5zaquPmeTu1O3T5bIa72j1mtP3rWKC8zO5G7FMefaBVAAP5ow+f3z0R
jHE0v4GyT2OEsLaOKRnR920gmrKIzBPIMhigm6MdRS/FPKwFxgygMdciWIjgtezICTBqP6zmNRu3
O19TXm/nvVz0HxR07k3gpM+CK+JVLjAHdGl5Q2mUP/ahWvKZ7nl1JjeHhDu8BaZyAAMWQssVhhn5
J/McwXIAgKW41hooqj0kyVDr3MFF9LnPpam+mee7CUrCvjb9FHc1iazZvMLsXoHYQ0vyPTp/jgVr
O+7iuK32cxrLGqtg6PSbeW2MLZLCvlxlZNulA4AlzHfkPFlYCUtre3+GpvIAEj9whQmpVWagQD/F
RyvsOYvOiqzdZpoTQl2/3DecyfTx8/FKGAR4IEirVH2KzsChKkuUN2/JwVvUG1xiM6Hv7clLZbJ0
iQ3b2dY0azb7pwwyumdpsu8qQufoh+HRq6ZNxp96ahjdC4sBVQqDTk4q0Wz2ZjC+d5sV1DjT+b1I
kuk42cv3gjRRGETxT9+NhErtBf0cE/zTP19/f2CmPEW9pKxDr1aebAiEr8tMgiBrC8KdKv8pWUpi
1g17Fuq+4Td7+ypQjAwGw1Chcm84u0tKuVyhHSYdhhUI/cy/6vea1Z3WOmEdU2gf7v7LIYzq8spV
DBiSyWW2CYAhbUFbumkzN/D5WlX3t+l/FDuam+1+IyNZGTEuoLy+XEh4bsd1Lv+Muvt9ei4i1L1Q
45Km5gZ2xs19lX5w+OuDL2XqgqZcZig37YJP9xTsfaGq7VxC7IhEAlyJf8ddsrHqby2KzxL80jCV
wc5bASiTATwY3xhAFdzvwSSz6YG40jUWsCkcMZtMOjNPpHBTM90l9NA95P2SUQmCnKXyeSu9J5Uh
o1lqvfl0bX95hJTjjezfmuUNdY4wHGRegH5RU/s3KSa8uJQBFIsTeU91KlwrxyyM1fqaWqWNecSD
BSVoEC1bnGYCify81LHu5PAsf2i1LefPTJZzWZE3ltV33dIkvcm+4hTNjiO0CaoTUQ9u6DoUxknb
fDwyHVFwHlaVx1iHD1rSq94YZfKTZdsMCxMOIe3f2/9qh71Dg6RYFrgZTpsAuov13coKyEghXhYK
eKSIVkOhklQa8Az59Q9yUlsREhZsisMjdQk1A9As2YZBzrnny1jau7CVMjirqYoXtMDfWlBrBSOC
KHseUGd52hvOWs+4zkJ2BjKFDH5b3M5cWzHjrVb26QijwHD+Ctv6NonfbbpzSKu8KYGMCqWbdmWq
lc3OaLX/maUyPu977MkJilxqKt7v71DCF8bc68CVqBM2FNaKA+WP4/AwMZh8yJRnTkEbQXGfmG+O
YbSmSvQkP4z0leefWtj0iAi/Q8n2d3x+cNQCC854mV+alc+MvguCuJMnrCtUg+RtOHPYQKghj2ak
i+/R24Y1vq1FgLhpRgtGHeBXGMuXrFUQYBGrlxEUQ4nxuWrDbSTWa6sCdHy88WteRXI4FuSn7oUJ
Faw8roEHSJSvg/RJR5f/veeYtnnCzpEpzwaTZg7Jl8ba+KyUibmBE3nY7D8Fa9BHCvgq0SGpFtF3
1EQSgzeesU24+Uhu3m4wM09lyp0e69aouKj9EJY0xJKsDzXbcKnS9zy45xwf8UzrjIFpvmu7xfQ1
rfhJVnaduqwh971onwARaKwSg9cgkPtKQtyCWUK183bfWsVOpln4eDUkf72JKFsJJGVWyxrDKgvr
pwW1DhEvjBpP29N/nXccnCAXLp3jWl1u4+xKn2i54UImJx5CRLihiLPOaEG5PM36JEdn96dOTZaP
pOBKnvJnRJMvjV0N1o2boz0383Aqbv3MbvPXG0ZG8k+EbOCsDCo3zaEBQJYfbTXaydg7V7ceoN/W
kyB/B6UqE5JHcOU+l8b0mfpLNT6vEEeLS8/sDR9qB0Rs7ixoPP4H+ii1EZH/MuNGwMC5xxPpm6yc
o/5EwQvac2fWLzjJBm17STfFBlFDKhkYZT6YOGcbvBcoi2o3x6B8Wd3/2ySzd7pfznwoZT+DKsYH
M8n3WpK/yhoAbassk+llPVeLO8SdkYnNLPDhVOeMYIhb8vum+YnINEywLJEb75G6CIIZ6iI0mnr2
tRVM+Hdn+fAPulQrsqK9Y7yHY6Kklsvh6+yXzA3DAecPGgnj/LFn1Ncv2qXJGPl1qL+bTXnNvcXw
bTtM0qvHTXTIvs1hYqmrLp9oC6oCLHzlOlSzxEYl40aTo/smpX8SAwhJ63ZFQ6o4tzGQCZJcJW1l
645dV2ZUBue3pMwXu9KZ/dSTdOfxg62AANMBLv3Bq1a95QDjKd0vjF/4uEoxaDl4yXqQy2bGoCaX
GGBPXQbjVBjeVOBpLRgK3owp25lgLbdSGkWhBabczhPzbCSCnQmJdzh6+dLxtJlVd2HTLDOKUSkm
Rf+vnm7/3PQnE7QJJ0vjJewe/4p9F2RRW1aWTNR/iQD/+xaHRHZN7s6+JM/KrKhhBt/1rtGkjxKE
962TG4+eAMZjKqLO8HzMDpz8nrIwcRNOaZRAfd3RZDz+jrwnmqgfBKQkX4SZqVMFol+QWSJZeg2n
7+nZxgioyRvDZWcvZHpY5/S9ZhfEaShMSjPC1jZ1+wN+p0lD+atAwIlnerc/umO5K2L11RXyvqy7
UFyZ+SRsXJO4rNirS8YlIgCYWYgfp2LZW6LLR8BZRwSEwE4QQXSlNm0WcB1Fd0eoDuDFMqDxPKli
jLTpiMrDq33iJDASZ1pS1TbMPneV9saAmKgO3+tP5ffGxR90NVXvzN+Hs/aU0PFOwhYZCNlA41JQ
op51bXi5oPtTpKNNcHEh46zFzgH/3sHPuxvB1a9qcoAiWLTy232i2k0A6QLtNBnak/cMOUsEpdGC
vsLMAWqyROr8smBNwlTnlOQ9e6Ey0Gzr0opF9mlFX19oiPhFLvr0FwH6jPNBUp8LtPweOvX1k8vp
8UmSJwnAONY2m3L3nrLFgs3mzH6WhaF1PS1ZrumQTxsEme95FiV7qcPG1/UT+Cpu3T+3w2Cxr9q6
kn3VYF330MakOK422WMvSmJz6xfbn60rO+TlEZocUXsR4oLbCCXCgV+ByYfjkT2pPaffvNDf6Hst
wtiJ96Q868UQpfnjfOkGkmXA0Cm6+n8dPRT9nh6QvZ9QWUVujT2vOi3hkql6D06oB37lPkZD+a0J
pWrAKP0NctXfScoIssBQx9wF/Xbnvi1hDqno+ue8mIWZ7ME1zzm7cXxvejCpGmiHVQDRjyjovI5k
D0llSYWSuygp1ruLo1Cfw00th4P/B7TfH/EIIIo21p0TcbCWyATryBUrq8iCRnvwHPS1OdriW4nS
edVABBqTWk1EC+7AtHFr5U/EBEALTQ9Ojlc2a+AhNZshi4W5Usbm7Vx4pfloZuDBYHGCcPiqFPtl
6T4ofc+Ajzb8yyLZohIEpCznV+iX8Jzlykyf+xJ3RBJxbBbIjZSaB6zuNqv/U5wdP+z6IJhQ4Iry
0p03zyg/S1P3RvALBref+VgbNWfApqTSdUrtawFlElGP80GSDiIZ+X5f4jKW4H9yDEyH1jcxrz9K
pYl6LvUytVf7+duvf+2Xh/CgVrsfsI10eiSt+jW1jzvQal5EeTtGyapNBW6FtKTuTnk5OAecsdsf
EkBT1PxrKPtnNsK+QTnGsSh6oGV0RZ2Zd/YwCBA08uUUhBDHzQSDkLyObd5XwAFY7WJhR3TpmlYK
IqGMwEC0ZraqYQ2sC8yt/kQYUfFF2QzdpyvgGWpejtKH/WA5cawpBEaUzDdRQZ8VOYgmGnrUoLNc
NAqppi+QldkWWZjRBolr4mrbJnG4Kke8UZjJQHbZSS7ejogNSswhoHW1NlzfPVq7rHPPIWbzV11T
s4NA9JnAyX1VgTB0mROo1BU7g/1qmvCDtvNQw2ih5PalaewZi/yk7wxtRccimVW4ulAr4HEyzCcp
WVzFJkG6YEFgogGz2ERk/upnRbq0LezTxnsC07LRJkpX8Y5c4BkZSsfv11Ew6G/yOzXVtkLIvDL5
EeVMtOcOQpl5uReumDe6vRyzYZvEpyUDolcmZxXP+Ons1Tn/DM7Nt9mbxas6OiRVsC2RVzoZnTPH
YEv6F1s7XeRCPODjMf4VrHB1kqT+o3CAu22lCutOfFgpUnJEfBUnr9ufiWkoboPZFLhdUpUFtPMz
BHe09aOAVdVKh41njpZzTZzJ0PRZ+z6/1UV634zOiVc9pm4L1scdpa4gGRExEEhoPx4FzcD0ZA5Y
FPuaaCKwgz+Jd5GdxaYnbbANLvZG647WiGdK5PDe46oDt36u9ytsWUip6UG5UejkYd+m0vvVK8gt
0plJkohq4/QWtPfDpnE0T3h1RKWXtN96UHADlziEEqDLIsP9JVwXOMwW/w7oIamg39ZYny20Vlia
CaKKUd9L1jVV1H7lbX83lPatKwERIBLWK1lxjytACW1M2ZJNvOjKl09EgXIVIht+IV5r3GN3mMHY
oP9x83Q/NmiZy84UttR7uaZwfdVzVnF7bygp8vt7yQLRBWNTF2Lo9HJX4oG3wELiDAYnCVM+BqZl
75lsUUhUYhNAo3qkMKZD2+ltPwhuFCP+dJHzkZvIJrAT9ZDz3EexLjVdajlDHMJ5D3ju2WKnWXzq
lral3pQYgxnfACrkQ+9GupEqn9Ku3dWAxoj2cnoRe2MzgjMNvdMtlMBMTmgvULmTr5hPnuMzhTUs
9flWmBpBjxZmkQx2mcVhSizwzxdIFY75FjVaIsuCB1qwZQaJv9DyIL1yoZrwNwAT1PiGtqA3EBZw
iOnMZwglY0a5aNl+EJqj0JgD5D7aqzUTa2botsbZnc2mpXA1AKBuchTieip+AN9JGhtMkUE9Es8m
ixpPmAH8TastvoW/jT9/+7qFmLajNjHEsVojpPAFo07/BpFvhI3EpkDkbZwMEzWECk/oF+LnXYLL
kFd/OweY8SbjVZAyTwqhB6Lh32SpFX7OenHHs6Brz0TX7tBmYhJxnri+X1rqMMDkuEkazy64b/LM
E6P/uynhkg0pVMzBJDXIbinL6dkSXZBEYmF+nDxdvkAobgBn9H01yjwKE4b9XpjKmFhMn/1KKMGn
ZYfEsAbWLTzP87VX1QNS1zHCKlWAu8kPJTK3DXQ0iksuu3VNPHkdFunejySZzJg4XoIqUTb/URtG
l2tEqOv3X4vyZwDMlyVpM6OHW6YSFzdHx+K0JnvPfR6tG4Kn3ho7quQA+v7wztK+GlQt9zE198jC
WBfiDUlE2Sks2v4gX9UmOIn7s08dskhu4YALTyrg0OLJL0UMAXYa7IqmolGKu4Gu3nMfQ5e14wZ1
3YwbyyfRrC9dW+ozWbhHTP31wsbi/7m6prxNiyc2v4WrUEx7LWM4fET2bhmd9fRrcHZtOetb0Gyp
Zw98e0rlVK5qJQ0bWInIZbOchZBJfnTrX5QQbuEGy+4hTeOP1UXxWJ9gWxU13ONeUyhlPvVP0C3+
md9nuijYuLtgNUnGFLa/Z8zHO5YVbqcKtkJw5uW2odwbpZ1DjTGLjjpQZR0lw89eUb6VzBrXODkP
rTDU8cV0jhQ4fzVa7mIglAJwdKXROa9g0dhcP5qiDzVIxVUZsbpLpsxYVvtWKCcChKPvY3NBSrKv
WU+6TUu5p75Icmi5A4lyEuKyyvcqK0dwNgV6owcby+NusCZKOBcHwhNYz/coBxj/rAHWxsommdSc
ZjkPAbiZHkyIc29/xdFrj/Dn527neu/kMoRtEsoSJ6WlB66yA7YHbfkGHZPX0Nkgni5DtwFpXTfa
1mNbcwbKdNQy3q3uV/nNM2aUsNisp+qfrribh9VnN2Re4pZwvWkgDWELeHBlH3hOHUiL+7hssKhh
mYWU3e7MP+TFdV4YiIK2zAq+Q9OdMNAHEacidGaFEQt+gUFCfntssyIDJhiqz1st86H8i2yVF335
1bQBco+yHDH6WQHnzE8+lPg2n9ZHE0MlRSlh6w7W21pY8bABELa6h9Dp2tT+d7rgYjNxt+92eNDS
IoeqklVCjmhBG7/Xzoak55/JE5ZK6PbMdg6NNJh3FyZvxSUuVm9+zjkA9MuCJybHWplU9yNA0Ck/
UjKQZGiS1roBJiAXamJ8eM6pdwWGPoq0iy0MQN9tMxzwf7BTZNnQR/Y7L7sGNqQDbjDhbuH/XjKY
X2LzH7rhTrjsKuIP5lHg0VP9MPQP4sS7M2WkjCZjMgcR1xmh62SYyLhFY86gCf4CUhyCSIaelQIf
CSfyNlG7O8e0XmoTeqlia2UmdZ2OnFB+i6P792IfbntUPbPkTKnXmeKFilmk6R21q0VhO4Q+o0qT
66B1S5eqIC3BRzItH6s6iGAC0J0q+b6FNVCBIDqN03qkvjSiVUpDbE7cryI7FeoIM2Z2f06ORK5e
baNlhwe8GlZVCfAQFdn3bg/++k5gaA9OvKTo7ZEsPLjWc49JADra42zoZFaGQBB3ntITbXvhrRZb
KvtSbQZCqlReFFAi25NUDPEKdpDf9peBMFY4nvzrUh2+diTfkTDrZPJgz9MtSjE2UC5jtUzi4mN0
rsS1+796pYulRzcUDFm/rsamD4vTh6PU3TceKQDJkMjPZVdq5/oxZeEB40EavV6jsJPWUP3pwSfB
YxPmERVJfBYfLUoEBxre/vHM3O2/OlNCiO9uk4c82/M91GJn+TLAvEDFZM7hbF1fNNHj32DA7g4q
KuZ1hmCXxBGZU2PuT9LOWE10TcOmqN0gSMq9Lp4GmwmnyUw2M+oBjIN12MAB0wpTMTIGx1fF2Nvu
MDZDPHPIZLlnXs/3fC65LyPHeHUGso+9Fl+dipc+wZgJUrHTD1J9eK5EuUYXN8sUoGQgAVvvQVRv
pHxK58V54L8iu9cl7NdU2h05UpXE4AcJ2nu8X5sbe+QmdcUN57H14BG4NxZBMb4H8XuW4uE4+bI/
6JSSN5dA06CXIR74RwaX0c81b5YdAeHceUzWpHVKmj+ZNNSIVqMYgjaifQNHWk+rqooUIjz/Ai3c
yOCZ2OzHuVKg/LQxKMo1VI8Dzafe3DcVgE01ldwwGaQZ+aTDOoUKftnahrP1yND8fHaA+e0pjXyT
z/6Y533/KUt//E+vLdA9IJpbbIWVlmdh5YoRfeo4lDLYZZrrK4hn+uCFOv4RS8j86ygW8enkoFi/
21/RwEgfy+KG4LuTOpGtiXmTc4ekVo36pSi+YAZNiYn+bVzcL8ugG+d9e8iFuI7qYVsPS2fQuEBr
SFzVe1B7Iy5pJbK0GpNBsM6JvgPo5eqWKcQ7MjQXRC1vx3Ycqb+cEPjsSCTUztcwg3WAC3oeai/j
v5hrrdQJmwTO5U9UIdEvCQ0DKZmUECEZIIfZuuNk2vhuOR/CExxqjQ00t24oupWxH8DeuUKbfDgG
/0jod+RAhGK1XkHT4NdPXF3uJJQ34I6OZkEM4NgTQ6Lsrez4JU46JrzN3dI99vVks7yMwPGHQB9X
0+AQhTidWIkgyKmD2E7cpwcvc7Rzs6+ujws/3zbyQ/N9vxN9bXUg0O7NdBYk00/cb8MplTA34riF
V2BeE6nARrAW8IxVmL9gzDQ5M6nfg6qXyF83Z6YNOeMHzkC0yKzYIRUCCIn2jMZl4i+nJOabl15b
MTTM7AjmclSWRMPSh40CgPBJxN7ifubSqaX5GKlyCi/ZPws4DqV9RwMFjS80v+G6B96Hew9ecHKn
ja0DcKqfmaIf6bcp0cgbDhVj4mcqK04gry6/VrguncPbwmkj3CoNcfT733SOW6awq7KTCtBdwkHy
SgI3ety2pmJVqsv9aykqTOmB90QIqakci9sJWV61AS9UkX3G3Z5WR4J9QcEMLhUjTBJ9wLwXykUw
28tf2GZuPKqgX/Foawdp2B8li16sYNGlfSza6W8cmzA2lPQ+ZPUvUoOj2MT3/FlrvPeW/BfTX2M/
n/4z7rB5ViV3yj0/0zCophZ1Y+m73z96qtKp52QMyxoB/Tkjh5TBTohPsuVhvOf0gwTf3BpgMrKA
foitOeY5LkpIHTSMBeaKir5LwCQShCfglP5cyGF8+iRFlMz3FR45pP/JmcO++isEn1t0bNHb3aZh
fpU8j4meHpnPnFTTjN02yOrXqR0RjnRe8s2Kj7WRkdOEE4DSBGcM8cm5ezvmP9U91QhXscTWqdBJ
Q/HPVD+bsTVSlDDfLP8cEJ0hJue8PoT3OiCQdI0nNP+9eXHR8qNLHzGSNdqHvnOtZKzx2Jjr//4X
9bNnn3LVf2/xeNqBqLIk+IieUF/NdTXgR9zr8nHi3CimnodyKe7AHuPFZHkNaOGEykSADpB+3z5J
wF/Aqd/r0xuO/mmvspkJLEJ4JslB3r+GS1Wvg+hlYrntIYsi0AYnlMxjX44b3++bNuIm9OkCWuWn
XeDODTzjB+KK1PIxLQEddYQyxLLtgO3GbazBEL5YfYZGrZZfc565oD9xUMwD4JFDYtLyoKoLm1Nf
IBd6+Ebeiv36J1KI+pwQw2UXn9B4BLgWrwdHmw7ZmY72w1Dc84lH+Wo37AoLjYbv2AALJ2U2tWbs
TfJ9LLcawh4aBHJc0dO7C7aDEv6FaB3L63uetQfyDV3nPVms3dZA1es4jSgsCe/LH2rjSthq5x6N
HZjcQ4Xpw7wdMWlvpnc9AbiU/13Ly0mTBYyJw+jXVu4FSt6WePuD0AUI8TtzNLeOnXwbMLqDgHpi
uL/9O0MqSwukEavJtQMlRdoE08xdLA+gdLe4u3DjZKf0WaqGOIbubu3X99GLqYZNUSBlYN3kzfs1
oQW7+4W4Fqkun0FuH3IXFRm2jLtxjY4M0a4GKbUNuOk3H1IsW+iaebPU9LbNi5ycyCI5JjHHLBXI
l4IcDN+7QJy0BTQUH7VBOaW+1lssxylwNKiD2bKHp6JO9FncOmalrPbWpKL8by5AnVcXq0vdDXIZ
a+7yUZY/OLjrAZEcvj35d5vKzZjeuSzq5t8t5NFu3ZxjK+X1IpbfbjWwFJJifPCWaGTWhHYCtPTI
dyPM+dYyB+cAUrrVCQFF+cLK1jetQD88rmziCTDbI7OMM4V2PhAoQmGSzcpzrgKRAnDJs73jZ2AC
YPberpkYh68kOiSn/1Ghf+PBw/CmwD/q26gpKu4bYJY/TnZcqiEAVfDqjhqyTP1Eu2+aIOHJ+plX
MDV7RVaCnt1kbdl8w9h1w8eLgWF4kM5iYvcFSgj9uUtuNzv1/BXSakMwhwESHGPWSZpxWGY6dGQZ
+kgS5BwIy9aIt5ab+hdXgeuMxN0pbARQe4ebP+iIlEjfs4vTGO5oyRL2clvvp6vAEZXei2sUdPUb
tF+FN60VA23XuNL0o6C/5GofkVhoiQ6+p1RtN4lBzxct1T7ErcbsTyxFRub04TXNWyYS+12CK5uX
5vg563elwVfjUxG+5q9cFFFZJyaOSbpXa8a16FP69gSCxcUPlbyDoAYyPIsUT58qdKAlA14dc3lx
Nru9QY+K8MpKqSlk+q2oLM1qsUJp2ZNehY8OMR+osh/ToRpYp54lpjjQlpkBiEgBPdxubTDYXcWl
sKPRunSjjmOiHsYuFf9o9Z8d4KS7OJqo4y8ZhqaZ0CVIOhDxxaxIeAFppvbYlQa/wR5lBo4ldG0g
29dwhe6P5ZOK64kfxXeS75iw+ioj/hk94lALlS8ZU0qpRPrRIgOxC1MS8Qgu+pqqYKzicPnByzcN
p7GMC4MNE+OWN16E1Z6tzXTB5VfvLcYZPVkn75ZOjsTKVA62fdovALecmBdW3FNhSYFaBMXNDPpc
V8W04Djsknl38UNPmWXSVsjUa2H4+H3fJRa/6O2gFNBotgnehPBgxNrNnXmdeJkCfYUXwLXheznf
su2Y4pkCk8hBvIjPFll+gleoszIOd1X6jZHkNEsTT7+SbhT50ucFxkQtZo+nRbvchYZeJy/7nMXU
04bZ3Bno7Ox17Vn8DXzPg4owEH0fKjHxlYhS9fa0V7KdmgYMbMrkX8ZFQ0C62/VzoIIhf8ruqOE6
8aEXKypHsV4Zt+ut6ft+eED9qFZLD7gvPJap6RPhMcm2yh2ioxgTbg2+3hzU8lmaQvpLtwy18vwb
1meCAOg6QwIbhwgx0HotNE059lAM8Hmc4EC5DTRPyskxMXcQOqh2UtO3R4XMB4rT/FHlCSU6HmqL
nKNExEJSLeUgsw+/IPTypaLVNHQjp+Npw9Uab/mvLm433sVV2IiE6FKF5LrZVlipK4dmLbrbGhtJ
cavyU2OZe2JqbDwfGC6aVnOI8Ob6mC5rTpT0jtvzVkoyOUpjcDC3OulDCU3vwU/D8BdX4qhmIHAm
aVU2ntzzF4Uib3m7GUPBl4zrjM+TuiF0UbJ0UZLX2Y0aS6fBuf2dgfGqSPsL32orZBljQiUPVtHO
aDIZcp5+Ztye2twFEimBKW2pxctR/hMTUnVajQbW3clhtxZyPIMzEd8mAkuI1oYuewxFIQBYRSGQ
0TUzCrulrI9k+x2c0q2Z3RCm8HEBWMVl/ZtAmSfWj/MkQjOiJnuqQ5O69w2LLgTrSprPO0c+a142
NwYSK3o0CufC2IHbiM9KSpP5RaueIWfmXos5LTyA4H7TYqZ/JSdIcn6IbXMn+JkVvgjmswU+/YvU
beBnyMpZ+/ICgS50njAMQo3UKDxp62sIjKNoD/kDlPjEUL+RmjYHcau8qJOdYAXFGpVQSNgDLC5r
sJJfaFmoVra3tS3P4K2wNjGuClTCmaN0ttr8MSZMKo2J34L5GQIU5gLa2vdiDyGnzdOTItTV1HGm
ETvBE+Q2inaznTRQybdgV9CjBCSoj4URVu/RbEUkjKsifOBiSL7QhcAIDQ9/XT+VoKe35SOXooD0
8NSOMJeOiYQdP7JOc4L9/xbO0gOo+RalQ0enW0y3CR80GRyesjocmZhMUtrlZ+wGpycaWB4l99RC
r38k5tDIvYYuaLD1sNZZsz0tvmZ64gk6Ya0UKw8j/PBI/n/xNQAaasvSXxtoVCbR9HW6BVDprS9c
YEtTFPXa4AG0t8gtGIYykXsXklC+V6F9CQt0P8xPp5Oc8IGrn7PMY+uz0Qvf2rKh2ejkknqFDB/W
J2iPbIduXH35yFFVZ1wCMElEm6uZ9UtGkgJYMUylUxIkr15SFBsnVuA3iD65LHcMjeYyRcltofWv
SunEMzUHZ4YFlBuZYPn7V93pYQVa8PQElyppiLfyqcaQmUUGq916AddqKVl4718jSc9lEzhGlwgX
Sk2SeeXZoI+wM05sVniBgz8Gr0a8HJt+Gm4s02iI45HmvEVdP3ebUcSHJ5tXZoaJgBrafyrWzN6c
/xnUpWeGKi+tgmBxAbzDLHBUwjFX2kJK6+Zc+Si5/zw9/Gea0YAp+ymjKOD6m3dqYTdDY6zVvnQP
WIjQJOZSYvMxH9T2BTArOADhmHXwfox/0uyWGqBmyG/FrMEgxgCj/UPJ77lU3bfCO0Ow60m00qhm
bq11mrxxf/FKbDBSNFJCOD9OJgssJSmbUM36QPvHUEXOS8S9wSxEF7qJsm5aqnj7j0L6cfP3jm8s
UYfwefhWLmyJFMlCrkIYUslXmppEvfAXvui5M2yIAhcHDrDlVfpIjvvUxQHKEE/+xrkbii9sMyYw
jpxe8SVoOhyRGj2+m87kv0gQNNkOc4HhXwN54cfw4CBfjILhGdKyp6C7nBaqQ8+Iu1nWYJkkBFwM
6HF7x5PQ5ooromz9eB+QsyK3aPIPZILEWdS9WbP0UGy/dIguE2QwOYcGjjmkaab91BddVdLzdd5e
reOSe8YiRIK8ick9vUxozVq2E2OZQgGz0cPLCfbS+rPNer7ZIQznDZxjNL1q9J9dOdtFtNVyhhft
Ie8QXnG2lFI21xxhHgVMwrpghlI4vbwDpGpUjTELdQnR2HjZQJ+jp+bh+vjMXkrh6T0MuCRR027F
wKtPk06fZsZqYXWvQLKslFIRjatUBZo9sIz60IRqSsbD0U3m4geG/MIVBV5eqkqZRVjFt/zfzN6Z
NtBshjwmNwtMKDtFVoZyH0YNYnJQhcQlA8PGHJ+aU4HFU8+LsAlHTEJpmPeOOltPBbmuLOOgyYPA
Tt6HQEeoFyVhqZ4qyesQz1RdFSr7uVSDb4/DWrBgyzzPrQRIxkrqYdDyv5226d1IHq7ccm3jGJX2
KoD5s3MJJ1lY/PgqSsFBOv9V7XWQJCP8ANWTdTLj7wy5KzA4Wv6v3yb2liV8W3bgJEdy+lnIbqfY
4SRqhEeKdld3Dk1G7NkgOSwgNOUbMzN5xSRc4K+WYQOSYWMZ6YuD4RuaZfuljD8B6oN3tNH+V7fA
LIXt2JcZpLSsXZfgPkDbF4zxx0Ie9SNRcUVNvtUNPa2umAasjr5QrSPdJoROiu8dUGi9ArareYoP
+sI67pAyaEL/TYU5AJkjLbnIUV8Ven7K/O5ynIgAXEtd4eoVhIn8DfhsYDO3u03IEVXG7dfhXn0K
6E9olkwxq1vA2EYMOx/ijtIrhQUhVLQn7vPRYlvREOEPZozfyjpacyxbxdNYNLMUBpGpyIa7yJLi
MLO+C/BNUJ42TsIG3RSYvzdM9PD1NyLcEnTfiDMBrV6fNQFNnEmTTsin1KmvU9uZ3lMsmgqyLV6X
epA3MDSgc6KSO0sqlyBPZwO5T2M0lyr5lHeoN4nfR4b+3hkfB4k4SraQ7tnKRGc9Y/C7H9gxrRfv
gKYECRmmrIYDgKF7BrroLZmk4W3XfLsLr1y6d1eQ6RwKfoL4M10LK5ttNooB7MoGn2wGDKP5AKKw
088DRcMLPSVfTxIJD/5JPMtXxzMGM6435heR9yUTgGun4GMG/5XGzx8uhFG4/O77eStfaS/np8Jc
G+PiGxs5WN+tN+TjMkxhYcu6TWhUzi7wzfQVs6O00EyDzBjenuHk4lxAA6T3D5Qz0Jw/A4aalD6A
eWGIVsBVZXzPDBnNiFbo8zHrxyHmxh1EIlBJDDCkJJI4zWdgpOShJB79gkAlmWSPTykcuKdjOFRD
WX3y80pGphYEtphV6rK5cPgzvG9X5G7CQfoOAzVFMaYz32VA67xfRg+U5rCVSmCi/j+fn51HUXe/
r5nzrGZBOrM+jnthpemulQeAl+vuN99qomvvQw2ivX6TY7FT2FEFgXSPxmydjybdDL7ekHDnPmRe
4/KcuyeQ5bqMEKsHAvPTMVWn8mJTVhcstoDVv9Wnseqh7i+ctnFmeS9qtBMBAQKM2Z33DJQhRsyB
xw41kjrfI75d8JI/TAsLSj1/c8omnjuZUcVJOIKIf+YkwcnqZPYDqAKeForBop2isPrB6sjrHMrA
Rmc3If1QK3KKadIar7B4bTMjU7ZyoT7+FxC7dH+jPx1LBT5J6dVPBWrW0WvVc91Hp7URxMH9UhLW
qJ04uLA3t7trqcUFjDUywSM+toh2XDyJXjBEafCNerh/BgkVeypwy9nab8VoSylejHN2UwL+lMZP
ntM2DqWd5y5ALPY1I845dL0akMDvoB732gjVe8VnrWO4GHybmVyNUprmKz1rDEGAt5wItEmsINlS
pk6qgfCzJdXpIKjjT7ySwZ3tgCYrd6YMNAOSkpx/I9sSINCOLyttM7OPSZVQo+VvG0iwBNk70TWR
OKFT2jpbCqlmSeV5mqLvnyfvX4CPrsNw14gCUZ7MFk4SjukmFWqDWRGutrur8t435Y1SNGF9Zy3S
PgGo8HJaV64lwafx8KhhKf2zCg1Blsjrq+Pplk7xS3abKtG6a8LwzLlPWAbm9UN8oK8etyFNY/wY
LHEq4oBRjGlIvi/sLlG4LvfAwej/3CzF1CO4GrBZPGBmE/k21FVpeYk6Jp5AdNObrXjbHO/HjrJ+
CMaY48efNpy0DJiheiNc3t5PdZvkL+mpgn4HTh0jPGYblnXzZiN7KuU+iSGhc/gO/gRq7fJpRgo7
W/NRtyu446uytVPKXKZQBy+A6b0Rng+3h324dyYpDeaiRvAOzEsEYjdauPvnL9xq01tx9177vt0a
GX6vTods+aFuz0fosJjvUpZHD1pCPBm3NP3mA6g8h4lJ/9brdTyG2kxKTRGmeTLBTVo//njt3ekY
cNAcHV4t5S+hXUcWpfk/X8zyjMOj0wzf9c4tSckSuqzs930xFHsjWch07hDclnSHFoyLe4KUkorA
+WIaxY9SXTokgMseBmHBbf4a1q3pJ7S01wHWheMfm1JBhBWw3f7b2zAU+Xuu8kh3UAuQqPWsJ1rH
w7YE6l5tjVEnMbTMAkWO6kWDWgj81KJPU8qDMMH07YzN4LjAjzYvn6kYPt33EZQU3c8YksxeRL0V
urHsxtC9AUYsM7L9UMpHJA8RlF6ek17zWyWUDHoyY4m3/SjatwFZ3Y8RFFsKAzFoowbuPu75HiU4
Sqq0c1ttXdrp7xfuKi9hl0aZe+K1Drji6bk4PHXTkTLjczoo5ajIrfxQAhBFYk1HYPsZSSnvVJ8w
cBR9XwN7153tNtx8P/uR5bfZZczfMKwCnNx8ipRYujuo86Yj0jadqHPTVGUabv0OS4/k8w+Cjh0j
cDqt3DvXxiMSJTiVeNAKisOdZsELL3fl1xIZNjJNg4yk6UhBy3C0DTJ/XmSBeVW4JVKoNLvppgjM
P/e6Op06KJLJjAsAQf3ihALCtjNIg9LgU/4CkunWlt1eKioQn0XSfWvFWMiAVyA37VrFo/KQfI7p
Pi/n5t0go7U90LF3oTZk1n0be84C32DhWxMKltMMpIeQZ2WvJSBrK0Iazz88rAgDkiR4jTnyuTU+
XShoVFmmjJq1+CLvk6A26bn/SvfRtQstIJKDE3zEJJjYwyqRnEHMVYJPASN0MQ8LJQLf3qp7kc3N
KkXJSGWDtQjOrS7GFfAcd46xOUBIOqwM33al6vRvb3593glQpWuK0bPv/L3d1OzQryUGMIefGH10
yeFPlYQXrpgKNw3RGkU0dU89z4h8hnfsLi2tsuGKL5pO9pJJUuFJMhWH407g8yZdTXF9xmSzkcmH
y5USlC3CMl9rmMRKfMrQuqHhVvcsFh12OEOg87a1vedBtp9IvZJImHVPnCiQPsSumEaU/YGI1CXN
A7/mZ429qJk2tU/pEF3szIkh2OEzVTxlPhWOhcVsrkv8HmlL10AGWbRSgjiTQqAeSInoMmEwdJnz
JlFi1AK7eFJU3ibJFDEJAtEZU4ao6JTwPelWtLVzKjj3DS2Any6kjzKCMQsCXDpn6K4HzJYRvD0V
Un3YK0UfCoZ5AOXVS5jvu/jFZuv+4GIjCUOQcEl+3i9TtGE73DIwNf65OZofN9Nvq3XICzTmZO0y
UI4cJqJdHK/YgegyyISNZga0QM6fxLS7bFzfN5nqDQ85DSqT7wa72mMYl5k1Js7lSBhmHBgnLt3x
TC4XFscUSp7GoFXrFxdGh3h3KM/8U3/oZzqvc3jus3LUDgbPI4bLvsLpZMC02U/96M9AeYNGxlem
FNkaQYUgWqpTpO9RmWitx3fLP/gzpg4trI6PC+uGH2O/RTrN0Iq9CLHjQAD0BMK3KGZZQbb22CPB
UmmSENL6yPcFE/qP6uthdi4dYjg1A5Wz4SMUB32KpCZxo/RuDshnOkKZt8TZZkDsHWCu1PZslzrx
lwBLXXn65vr4rZJTYCW225oEoxN8UDxm77+bMdYkOWvm3J7Db2o13X/lsJ4SZnxk9jEduwruuGTI
d9gX1l8kDYXdUbX3SbC1F95+r28XZGJDHFWPACh/FmDNfuwz4nLhxvrni/YyDnnOimhTDAUKcE82
NlUT9rb3Rq6eGCjR9QB1M5I7rfQ+qFKEmhbon+Hg4uQtjjNRdt3IR3IgepWB23FI/CHODIDpb7vY
bi30kGPez5BD9QsPnlJ+s3Pv/obfk3MmlV0iE0eW3cRfM97h9BiPa97HqtINVfD+Bnugia2pwwbk
JpvPL2MaklsEMc66EnxPkBJZ6ezI7e/JZrc1cSr7Iz4Uw0rMlhq7UAwGDwHyg6Ln0KmIpyPFlqVQ
zk9DyaCbPb3x76ly2qfiFnbTs1Q1cB1LTFhzsWwJ1kzbnnFt+xiqoiRqkhiIhGigXIaPu/xzKJcM
C0Asg2N6+GrBZrKRBHtwFJ74XjlsT/JUdGOKG/0h3Rkx1vDa2JHeVDT6fE8NAXKq1y70dYLpeZtJ
emzcn6cflzKaYBfmZTnibYBEqGgZjaerxeZDB0MCibhD5TvsExXJebB0un5V4N5xW6KOvw78rbGQ
tOKZlWMDNwNZBTpTB+A7BRgB3idTzaa8mciJgglEEFVS6JIAbIU0/Yh9vPQhdQJcfcDOoirHtal7
Ago2QmC1mz94QDFQ548ak+Xg/DdAfzQva1Y8ePKHyccLl8td9/3Ritz+zMosc8Dn0zHO9BjKux1A
XD9XV8WDMOMVwzmWiVBMjs7eTRHzDOhGFe4Q2ywSKbPJXszjSYivh9e8DX+pfjA7WBCVPX6Fs+IU
9eFwrVzV2NMlk91sR2uKnUschWQDfCyskeicxatPThBV6UjmCK3LCCrMYElYlxPR5D0i6IMDGILv
n0aX5ggqIhNakCJcYj2Tii6eTwKexzNoqQ4ckN6hl4VL1ylsZNwKrzPAkkAEiPtzrzuAtqWbbo2o
hvrdCHV/wixR037JY3yx+UMHkcBLJm3fCYAewZjAf7CKKbIH8VoqIMAitWEVz0K/7l5226sU0pyB
pT1kCkgVq90P5YTp1LG3fGvj+ROFa273XFLS9AgrkpwRrZfrlZLpFPWyv4iLrtxdt6k2OQy7GcB3
BdRxQSrXU+ye7gSi7bmoBhBS9+EnqOvjGqdblChOuYtCpGpodm/7YSBeujma011BsJY/mfa1Btv5
9o9A+LSK1bDjM1SxFJE+mBQFEz5KMFXIHQdDRYRLfuBqpVmesu1i1jFRUtXgQEqhgAvDf2Z1jTJI
ZIeXkCWOHNA1x3O74Al+lWosxDl1hRYXsJLWZZYbAnSkPNG8mVcBsXB2l6/CiD0fh9Hq0yIPNKKX
m2EOr3Mn6UKEihhDEN5njuulPaRs918fu7xCC+Dppybxm3hqBg5ad7XYlr3+xoVSLXXfry8mM6HU
eadC+Lyn+MNTFjU1yoNPufPCyM/pgYsjfDBb6ZWKqvyG2tLy0rAHjldyBzmrbDHbjhdRm1IdYYkg
c45damGjrmuoxU6hZG1FMRGZ1h+lvXWiVo4CyRYYpyT2f8j3qt12jN1/Mzcqn6crZ/uSW5HUzJZc
tUQV4RevTTxKpjXOw0sM8QH9NdDrcysDzBhccXCsBgdjOrnUCqOxBSJRihzH+iZkjQorHNVmnHt0
IqYQgqazF22wMTYfP5sAXstYdlb21yKZXn4Q9pKGG/lWDYTzVlPVqJs30Zxr2yAqQfKbJBVngqIT
Qn+e1g9khXGdVfPuRPlW/8GFemHCq8eTaH41v37agHmJfKHvD9SGud/pX26lHMy4nPnuL5NWHItC
7IdYy0STZRgTVHZ2AbhFB0J5I+16RxvF6u3jK7yFEyCU1Fc1HCQeEJbbthTrOeSqr5ct/gllSqcm
NbIv7FB0JE+kdmEkbX7LXaJ4l0RuRCrjH8P0l5uiyHpIm6R/sFkgAJPDPdJhgTh8XWRpqq1Y6m/2
6/AcgLweHl5bUeEvvsOQxqBrKwhsWyAm9mw7jXPQ1ZR4uSwsChM4SVsjBsPgJcKo5quBAwO+bL9R
PPS2lxP4CVYeU33ZqNgDxBCsrTOTH6FjgwP63NmUj+7lE1ADhVVzvDFWxaw62J4zK308bCQo2L20
EbQ7rXFD00vogDxS8WyvzHJlHC6qowv3PyX/xoVcrD+AowS+6apyTTnJ9o2ION+LMaUE0mL57hTA
cJor6NZIKCCkMD5a+8rWs5sr2kux/u1hZJr1Wy4DleWDpg4eICT3ylgT6VLQZxf8sxW9ExlNghva
IW4bt/YyL2Vrdlva0/6VCGpvGlkc2EjumX/uYVle/lC4J4ie5bJWGEbwEO2Ovo2frZyhbk4bSsdX
z2V4pdNW24iy1wAxXlGwdcZycGcy2gQDsPOwUrVNf+tR7uFQMqmWKTNzSw5LFoNv8y95pldFrKxH
ApGqbQDHENv01SWvEKo9emDgbyAVvosqdGNX00HWMgHEVn88LhxfZnS0K2apsCaMcn/Bl+kBRFI1
OvoPq0GJ/CUnV1njKsJsUPE5qPwb4V544dZxWDsIlJ/sSJCNTUKIeQKIk02BYqNNBEcKsEuJ+V0C
a+FPzKBzQSY0/OUlECw97ry0SB9zSQJqq9klovV+yHkNjV0U+ju2x5MtBqR5Kz8o6UISKAifwkZ6
5TQDcIVHloProAQlUD77SUuLWNT1wmU7K/oMGuzYO+80hUkH9vU51Euzw7iws69YySw2i6zIlTsV
313paaNBEoihETZgRJVVR/agKnzzZ5WEorlHLmAbWbeLQyhfOra7y+POT1qdwnw/AFiQiKM8tMZu
eKm2PpnEGCApLohF/aL5ZAoRgg5QFgjYfnnyO9UNIEqsM8v0nTJ5VQz/Ld5jC1dRNZYBKFyY5rjq
Zpq16VhMEW+2AeRhlGxSErUZ9p0MoO1Le0ZP0vlznF2/4+UIh/gRczBMB0ePIlbgV3Hvp08jpOr3
SvDZt4Vao198rqEDGCsedpqtquEaUlZqfiU3cTCOQ5a1XlXDKBkUxt9n25snbQpBmFu70/8Udm18
vPGNTgSUciP4krdNQhNRTccl+hW8GWIOtw4lkinVJ622iJjkR7bgQmCXCVJXrClEA7PUINABpx0l
J4Kv5xlpS4lUvJA7cSV7aRXiIMJVa+GgbFyT87sIGFgf7RFp3pUqEi3t/tAQjugS7zOb+39Qqrwp
QopS+R2s7SBXn6AtIG/YPx5WkO11FsmZfZmWBr2DWB1oEYZtwamKiv22mJzzOCR9PfSgdPkLDi2M
wR/Yi5KeUaK8XvssDnXwYXKkje0+nTO8kCDkcQ7TPia8sqP6ak4R1IAuXvwWLk62kMg28cobl9u4
KsVthYdceYw9UBVYa4kKO0fEdox/P9IVLJOpmpur6+TE2PVZT9ytpQC3C7Vs1pBMS7mfsth4SNpI
xztx17mYnkXDcdbPMFcLh3fxRYK6p31bYDWfPUMBKId3lT4hUF35mQmL+iMOliW72PW91O2cFDsX
e5U9WMAt0A9m8wewxrUNbgL8SR3YP91YkPxAw9BTt+gjxD/Anhlwf2W3PgXvaQWDNmh6D8vKRD8O
BxS+QrgRIA+bM7YxZQcBWUeZYmSf7NGNKpzJCRFayx1euyNPtYLz0fIVtoS5yxU6ZDpcDMzTTpW0
iHxc1jqJkdtfvpfUlzFR0eUM+D/jDC8UU8ih7Gfp+6rrhRQ/s4goF50hxUSx9yKNVSozetGLeSn5
8DR+43gYp8lODHLpxPLR2SwWuO65FKw+XuQ7E7/pRl+JAM4f8WrVQdfHv6xcpnRcV6Vmep6UtvXT
AnpWJHAmYgcsaD31McnPH3+Ng0rEsx77WjoG5QbYkJwLN/PBr/WoMCWXKIkg7ac4MRl/rcGW42UM
Uk8AxGB/Q8ZX8VQreQxH51A45hAsXZCzZmq1Zz8SUTc+M5dU4jO+IFvR7fE4bCOn59IMjVLlXpKJ
7WooUgeiKaUewbLug+NNPsxGx4UlCHemFAsSdjR8xSc1ubegtZdZ/djabpMMZzi1L+6+DJbQ1Bzu
gU2alJEMkwwkbqmq1G3ajtP89TM8MRkkvV98ZEguynHbVWSigWQZnTYHhCTXC5E3YbFdIua/X20w
WF/EmmFJ9CNAjNqM8SCfM2/SA6or/nVmfoYbjQdYHfVUBUco4N5y+SA3+bWKI0jUkmVmGzMhJppn
TtoBsAy0Ff1kGPwxxz1YHnZcxI/nTSFhxQjQRwqs2kbKNC2HUxkmmsRE+w0uDTU7z8RPzeBp6Qio
A1ybYbf4t/T07IDkJN7GmRsQQzhRjDJwJgscv9nps0UcVL/v2EeZwRb5X56GVZLdpbxmZlAfEaMi
4wnIz/S9W4NcgokSUdAMusb/7gx053aQ0plEOBjK1KC9MhQrjDRliR3MuYdCyULlc7VXdBz3iFVh
M8ESxjYgsSpOZK2CkbtXLwSKOb0AujRZ8AQDtuq+mVQtb263vLs5kUIE1Ltp8ywgdFetla3STx5M
IPm97GyOoYWnDMa4K+szOKsANdJSuMy0fc/6zTvn10qhKozfPdc6Tm4f6NOkWUeoHmEaBt2CPkvM
zlVQhuQYayyRFwGSREW5jf3RFVcptVTTJZvq3ZZE4G0scYITlMK3qkn+kM/p0hHL3qukjURXtfkv
T4ql1VfzrLEn57B+SQD3XiFUL3UwGwCL92qGryO7iEAcGGWNAJ+NgR13OZCTED0cKiJ90SRlitLz
0nGjwRe9dIeDFtCdnxyBgB4ZWMNvrhzZkP9yg49L8CXuRme169Kj/rj40MvkuIO3f2sQMJvwowWb
aHZ3iMmTfJIGpht/4t5Xj2cYxKRTrD0TgK8lTxbY0lkufvGKxnHlgIn+VfQmS70jZ19h2tVZlAxr
1GWCVtkNssafj8SfZJFcSEtL+ljlE5mEpQFGwtgRkEpv+u0t4r9UlkuOCZDJFCHV3mt7kfZsyaWy
H8HhsAVsXudHS9hqvDXdfi6LAiN4ekZfh8xkcCznxJkr1c6co9NC8JwSEm81c+BpjqbGZZAjC/aI
YHEZZK+VGAI/7EYekBacjp71hML0sR74rH+w7+WLYBBwB545SdvVjo5vxzp+tHS4+6I5PmeWXPhP
GQydbxqYgJlyJPXwuWPZr2v55m6xPGC5+ohLkrbytDTejPfBMp7j1WSKoHZlV3eeSOTl08Hzl0GK
mdaNwy/IMSbqP1Z7OFp4rtydT7ReQRYP7vUDLyIyvbf2qabnVOjAmP98OqcKPICmBiegj0ZJcl3Z
NYa0qMGkOEeuBJINrSQD2rGL3HofTd0kB4stWdekeVHZeQMEpKsC8ZyIiF/26KEloyRiql6Zs6VH
tRgXM0YO2Jk7XlNOT7iEjkOkkF/ti/Yk0xN6FnOIylFwmb8P0zqH9V6ieZMVlVuHoxoJi1QB+XZ0
c7FKWqR5+XGzjmt9axHKH6navvdnzLRL7dqUTJqgHKBgwdfaCiJMGLbmO0d2dDdz4TMgis8XbAcG
KOEv0ZUIWG0x0pSFYLTqzOrJfonA1YHdmJaQsx864ZrtRxeJbnsYkmoTAjFBfNURE4mpIYR6yK5+
QEG/SM3ss2oUgL4keQ5D5r3IEq/rbWtQ+V2QDRkmyrHTvoxkSt6eP+Z7o/1atiQ2HrwEic1msKOG
C/8L0acfkkSCmn3z86UWZaVrRBi891dhysJsk9aWrZnFCeYCQNKtQp75h5aSBmGAwr5v0zrm5nfa
oMzG80KFYhgxew25fkvkS0cY43wWW9pOVOLQV3z11qcbvpc8nD7pxfGYxgz6nFrgg5VIXN8Q8e+7
ukZGejkEEdja+XrRT6DXIxDsoEaIPlGIZBPR3UL/+YfxubIRF15GDhozpX39bL5UzD11+7ta9Cct
4DNu3vDaCfwsz2CvMnLRSBEmFW8hnfoQNDm46QEsAm9MhFfy1fo9QgI2u2+pGyndnati5dkiMsTW
Y7hjYndAyS+XBI98QgkuY+tRMm0JsjrS1eyQ8Z16+UFLEUU0GKPntEJI/PueRZ0I5LeF9vY10OuK
T/4N9+GD9BD9KRRZLI15zuMEkU4ujDXTHrL7s1vLkczfkqzU3dLLf+ifM28idKU/n/HTgSX6Yxcp
i1rpClH7TotdRJG+R1M/ewBOSKIfVKyWRcwbmJRwVkGY8epltp742iLWQtaFOlpHD2/YxGaHOttw
n5k81BMfha4yNA0+q8vJMRTR91Rw0uZqOxzTI73ZhDMUyLZjA7ifA9at4LSDdaqeVoBjwKn5LVOn
8miv0mY40GU1VCDqjdIudOHLcz8NaCxtXEt6oxJedbSnFrOj9ZlfxQIv/chih3cKZ7XjgC9Yna78
fVIR1BnIhRq2RoulOn10mdKyAuer06YoRCmc+0Adx4X612gc5Mvbch1S/rdJ5ST2CB6hB6mccXUR
8A6z2qQcVdBGQdBUGcBYtZeZa6RvaFlKeZsbUkseR2IwlNzQQU+h3x3yyq1iDXhDZNVLaa34IPpA
+imvlS3ys0U6NaV5ue49jvAezXewMc7UDeUZBaUeOIC9Yq03gd4aEHWUt4pFU+akI/2HvnNmqdGr
UATn4bGEbZPcylg++90zhD4QF+uAjYaWQj6wT4aaO32J48ss3Ud53gDFiS7HvlyowM/bLAEBsGiv
ifbpTWv2nV7j0usLqIUQSibNbqvfm90rnTIWtKonT9MP2+zZIEVIh3tJVhLMAgAP//CUJkQ6WZUC
ec2JfmWlIbsxYpnU7t9Igl0gDKCz5SxIaH1R/goOCpz01Q1kjnHMGpD/QHWXvaH8bBUf12MUZ2HY
GVwWjp0g1kJUahtg/tYN1UpFGb1mbqfseOwl11i8mvfu3eeLL8VdIEltyOB3dnNp6MAJej4YaDwK
kdk4qEtYZ/qYY+MQB4tqbu6E3kb9bXfFtDmbbQZbK6Glf1cNbGFXmZUdsXIZ1gEbKEIfDU5xkdXv
I4pQ2OGCkFMnsKoBwLPwOdnX98Mx8jTelqw2p/rh/eaS6qwd3pfRVowQwmnsHSDrru0qt5AZh+UC
FFlZrPM+F9jqbZjJgMt/dAhssn9gkTcV0Rjvov4WG9j/otfLQhJeSgQ03RqowVQa8o9EqKWIi5FE
iV/DLyTYOPw0jUreXcNaI8+mzZYcSvFwhBX01dcKJRJszv5mRyd+eUZ1AnU7AFf0esyFKc77/Sjx
tLvP0lLuRl5rnW6pQSf6R8H4oRJb3rkmqj/z/YTtSIlNAXkNgvWtkWwDX4a6Qv+9nDrHk2i2BWxY
nNGrdm8f48Lt5fLmhC94LFs2q3gxc6vHN7X1H66EUit7fjD0/axqtXBelQi1n2kPmNB2oNFUszBt
sN1xhwopb207oAxtIFR+AEym73QaFplacgesAhRBAUFzU6oFfmdTHWZFRqbWk7aPuOPfvIDlgOY+
+QZZOL8+aPsA4b/amXOeg1QgD56H+b0g96ZIFJXtx7atIN8fsnhR3aDWiuo2rokK7Q9eJdb0RKli
0QVcTNRoH5apfpT91TKfyS3WgNx+t6DMjmSA95RWmKD3PVQouJW/G/oMrB8ql9MV6VEFHfOIOofq
rt5TvW/ssf6oNW/4zMdOrc9SbLNmqG9qEX37tb6ea7qMUWAEEPDLtTutf+c4vW+iowSbjVZifIID
SynXpKyu8HjgRjqVNpuiAZ7b8OXj8ZHVS+HrHPhasOeipw5qCgiKIHNCrIvOJWMyBBnJVIZR4oC7
WfBs01iKKCQCsOIMddX0CUC7Eez8gTSIB8q8k8gD9anS5gPboVZeadK00Mjw1+LhzsudoKE9DTYR
mJ+DkB0vmv8kDjthXRDmAjh7zC20ACzKnfUBVA439Ov9KXoKpy/UkNgye/UfBSuzJgOY8r4qmTkA
zsCY5ZCEINBgs2oPeV4mMSyNwD4RA9Oc3nmz0RYh0G8fnEhKd1nFNPciTLrLxn5Au/jFw3xakY7X
4NE17b4zyssRpKr/EiHHKBP4AFViNcGVxQj4zQfNHhvd4oChqOQZ4H9VIKFWKx+GWhvdVq2sNAuO
85hbifHrIF0Q0uLFVX298qe8W29wHEtuCIN0Wkabmcwc3qXinKgMKCGLmDJ3hvPrMkdkamnZgE28
xklKTq+8L/+Szn1VqNPvT0U0Ns8+HsYQsNP/IifUi98ikQ15m9KONHpO4GlPm7w/d3DIfgsQYlGa
/F0j1BwoR2szswXQw75+WgD1OXDJbT3DKXU94yO3qrR4Ep5OGnZrrRo4i5iwT+4MlzORjNJMX71F
9m48AxL8IZfosL2bd6vpN9+TYJVb7WbzrbjgJeKAGvWaAlwBPmVzTIO+yxqX0WmqHKHNhXZudMCi
R8UV8SnyyNZ9RQ0YQkk/ZfR/nauNUIkqt5ePEhBNT9JvyVPRH2Mt9gLAYwKJp52rs3LvVby/bqPu
lY7s1SXl4NUu2pBDH8NfHHmxa7CKxcN9rN0sATZApGtfjeHdUT4c0cPdw7KAZZ9yzXvE3OT7geQB
3oviaEyAvM8Y+SMIakjsDtnN9PkrSTRKh6mzL1FwoNuO+i2zU7vK6Cn/LV3rEpO1DKjNB0WG1pY7
aRmfmAK4IawL36Wz5nK3W13QR0FIdOYuL7MEFX7ba4WlNtlEnUG6jlm2kXo2/KUegAEApSLPCjyZ
EbUi5wG0ZqF//2jveEVbaqBEOrckqmSFRsY5LhClYGJmGK/0zc4Qq07ivhcX18ha6zrEw/BoP+Ac
7rMYoRPZnKCDdqpEdZGeQgqOor4N2CAeT+Hs81role7zNlY3sQ8M/wdwYVsjmja/Ocwcg94/xJhr
zM4kpKF5lPcTf42+CXr4M/MJVGO6/qMkB/uMwbktzYKL5ENfEezecyj+7gWK50ijfJyeV37/pVjJ
9n4E83LeZK4I/zGr4RbzpT7/12pn5MKknbbR2Lr6S5h2ukk/2KagCXXOdhHwTShppSDlJTk11JSg
3USbSEZd6dOEPAVFwsyGj9A40Yjar7a8OWWXT9FCq8LvthQRrjb1363ddJU4AGHhGvu2HulRVily
P0UTepS+esuXkiMPzfhuX0/joAI8llG1D7daxeFxqwedQd71AySWkslesFY3yLSQ3Ynqx9M1f49L
vfQKdmloJ9eHGa4hc/LTF5ed+HMgy5iTMWL3H1GrI4RRl1XRHGqSDbuCSIZQJZSUxzTqAeauPY6L
icO5nbA117CawDEpCC9/sLZk0iTCuURN+Ow00oOdA9TGFUD4gNM4H8ChqErSvPcjvRltgDq56eRC
MifcS6Tsft+L5E0u2740nwrL+lzLinYIK2uhrgZ74vC9ht6yfOHqe0pOQwAgVAQ969SRPmA5pJIb
4klrdHI7D3FQ8BTr5Bb+4s3hbX6hWtzntDMW8Dq2KswXRK7f2SiLeQ1VZkeIlhpCsLZgXWxRfRAR
gwJFHepP2xXbEK9FcjjM0/0WVq5F8xg9RH3QNB0KG9qWPswnx8e6NvkQJ/V0DhMFghgjqUUCkkFZ
AIZU7bbkhIDYTUalJtsSr3eb3MVAnVVeLR+CvyrfRr41xUqLNUzURnGYrT2qneuHmlrAY1uOqsQf
igoEY+I/jPAfTZhqhNmbCchBcTHAqDhEBjNIFrC+XddJftzwO36InoqNYmJoKL9wHziGJS/xs2Gm
tga6JAQlURAYKFhTRVLMBCjQdluk9r5eOFp8OBmNIXx8FoFjc/tFJ1IGxIdccurV90xSFTTNdbfG
VZZwWxjvcoP/oiUior4wGMPzE+DvVksLqfAfXW+vDqQ5+WY0xXp7HArkS4LtejWHMT4Rzpwg0Yqc
WpSwd6o4C7O4pTEnk424XxFI9TWBdXLsC3j2+Efk2uWVn6ojcTOyux6rXMOx5rIKA5/1/5eisPgm
l2PU+Fcqf8f2h9yVIYJRucd0tRY5w5Dk/mydsiUixQjKlOtZKQh6R0gdJQXUx4jJEEPzUjzaBD7A
Qu6ACU8N+7+z0enb+uGlSEMkQl5T0uE5/nPpKusq2pYRMQozrStKEYfL2KHYN2Cy2mPQji5yJxPl
h9FdaIOz2bw1ehvSCDIxyYrBpTZJTsdWn+PUz349JE+r648tArO2kYINAsNjzG3Q+IXccN5gXZQF
fVpfsZC4umOqEukixWRg7+LLmJhpWtOxD7rPyK+IPvZDZmUCG61rBEAfyBHwQYufY2NS8eYZoPY1
8rtj/nEF3FS7uLPY5IndcrHupI/Ajc0bYPhpGmdVojbFxws7DCORWSfPGYTiDP+BmdkYDWJUtijT
OEaKIGq3AMbM5qk9bBQ5CC59SfA/y+dwIAwZ/16i/ji+fXMYuQuuEZ42yNbNHykh093uHnLoZHUh
0pDf6LQsHMdCIvOt33rVgI13POrM6r8Ueo0xXRsL15tFp4N3yybRCOURJvFz5Cuiph0mXZRk8Z9f
WxdLk0df4WEXIcJmaA5GZ0teKFKUzcCRf6VyS4Q+DPRqG38aa+1to9ECzDkhlrm13MM7zpVFHCs5
XWObETNwTzaYdqOZ749QHRstTHramBng60renDZQHnsOo3s9mrYhp8xxTwsmfiD/Y3uxb8T9DZQU
LN8j/c9aivGrH10Ek1eBr23R44/h+3SBRswcqmD22Sq2jeB7FZFq1/k7nmNIyzDJT4EqnAPB69/C
VgSAiv0PDfYLQ9K1tSR6jVHWWWVa8kJZ4N8KlzHOAZJZQw/8uwJu15kcic0IOKQenOaRIwNByAI6
0UEVvlk8m2d2g4Gu0fWVjuAHAw4pgF4tL80jLmDf7h2X6knxYl4/0oGPS9lhTiXJ5TITVPnxBUAm
VWbkYLGt+irMhrp+rO+EdmlZed2Gb+5wSKrWYhsA/utke2fhNsMfpKQEgOKDJk/kuzwB9cUG/WrJ
C+fhRue3vuvKDfKvKtv29CpOBXGA52JFBXW8GUDk9hgaTsZYWvku/WPF2lc0j/ef6r5/exiIo5f4
pyREYT0CPqVeaaZIAagAGQPZ8D1KN5ucmQ0BM4K2unOwW8g2xNA9jeL28dQXL+fBbhJNuXCg2fTw
PcmaX9tO6pSFXLKfbvQHxhby4DZ0k3G+rPni054ku8SB573E7RQd/wp7ICJkvUJoAIqudsTvOZ5z
cSe2dEHFhKaZquNZyZyFpJD+Ur8zohbVKuqkLSlLs58yYhMG4F4HIbD9KcP+QVmvdnno2YhWuw7D
0GgJYU++hpVuhgYh8cwfDvjUTcrGh8V/EDlXPnqKV7gF4VkhfpLTjJ4byQCjMcJH5IT9q2QfGd8B
EGpZIK30XcNZERoNr9CJTLgukfommhyLiniOleX7RkthqNd8r5VIkC1zAtzP5W3PMR34uJ8s1jP/
xN6Nn1ey2EoV+SaZC1YAfR14t+dBMOiwvN/Vg4hocZF5bAeWts5jA1ZzJ9i35NUFjR6+7uSRPmb9
+EVORC74hah7gfNMjlh2IJHc6RmjuwqSJXHYCumXr3x4hwKfZmW/vVkmzEbzbSN8X3Q2CAUL5eYZ
sAeVMe4a/m11CVnnrZARVsYRkeq+Q2Sax2ecFI6rzYkI1Hp16g6XFqkxViOHQMs4mbW9g98SDdZR
HXO46XoYj3p9ijf7IJz4Pp+88h3nxAaGB7tNU2xrZaYFmO2sU181oJt8ErJkZNNwjxV09jHV9JVB
b2WQB1Q5taZCQvS2+678GzTYdqXZjd/jUVT/zzyUfqf0XusGsqBBmgFy1n0n67R1HBAQIn4/DTRl
TeBOisUcAaA/ICuThHjkOGXQRvVlu5/7Vozq08iCzOCvBraumNie92j5mAckJMdGD7SBu3EaTV70
9u0nPl17y/k61Ctmtzluog6vM8EVuHfVAzaW8W5aqd2iMEyEENJntYvoNVXdECQs8Im3V/YSq7hj
+thqZpr+bq1quqAfEj32U/WPMg9IMonI4ZcudF+/19o8Wk3zTm7FjWO+5BeeeJJAj8jeFGMAMzXS
BxVsr3KIMqvYaXYycQF629g/jFtgSFrlyA9moCNCBcn0NIkCnLlxOnyplWf0sWErjFMgEhBDE561
yHTLguMbDuw/fnj+GNw9OZxImrK577oI/glm0h7Swdf57qup/z2Pt66HTONSS/dQn2eecJ4N6AM7
4Te9u8Fv1oXgE4GWAXKt3uvnXhBM1u2oUvpmH1u4x7Mxpjr+cUfrbJI8UwYGSetHQIWvADfwZEpB
M7fEaQvN1I9ICKPGkq9jiqHM+d/cwA+nSfQpOmXqjmUO64SHMj6Z2mo/pkBnjSPQyTHCrajU5qUF
kbMq/x3NpslCxbCRlWTB/X0CxQXC17aY3e/ZzPMTzJDTX70zHiWNIVJMrRBZMP1XmuUih7Wl2veP
jiPP9oO51Yll3udYUQVKpTl1r/+k+/tiW3EcvN+GPKtJXo5IWSDn6LQLyzcstMZVYSvJ5xYaTLxE
cR8N797aMe1rKOdi4K7+cf4U0uyuzPqvph6H/MDP8KWV9KWbec7Lv/1tF44Jk9TK2IeXL3jlrkHX
fFEBkU1gRavm0zXxmkiMg51OuPAQ6zrEK/hVcWpVW9O2b0aYr7JdI+CCLOnSaUbeRh2mUIpL4XID
HPSYJvLxJ6jOzJU7evHa/gP24+j+HJNQ0ZfayYys7UOxFJPXJZ+UKJf59MxyUy/+mab0Ho3I07FV
XWFaODUComc0gv5vc/CxrqfQh7yKfC6zuOK4ZWQR5taSe4g3D7Duopa1nUBEou08W/BydMleVDA1
p5jRIMegBsN+QMjihU2R9TeYtj1XtGilzPCAfdYESOFT/wpJx5kqQM+EAJ72RzozeyeQjusi2cAn
oK1AgeCk8sQToHuTFXD4m2e0VA4mOaho/YA8lZSxtPm/Fhg6hO7aU4p+C1JfjxdB51bcATQrq7Ap
1x03MvtLiVoN9bPDRTz+41wya8mLGqb8KN1oNToZ1Qzxi5nHcCmX0X6EYfynbcRxeQVIpr3rvzAX
nW4a7W6es6ftNN+hHFE6iHJp7j5BrrHT+o7x9pkYWt8NcfdPqG4R/mjRfkxX322Mv7qYpyncmqe2
3HfP+GU7QVANbho6W2OtaxO56mEegwuGKXir1vd783kSKXwVskEmjpM4o+i8ZEGVhLtNPnjeJlSx
lJTkoEnGlPTZmS1FBpUQaBtU+KhsbGVF5f4NLXpkkZC0JdCjd1BZbuCgxPb4AQxriG0gyCJaBHHK
c6fYhR054UowWZ0fu2dbUsT4JjKa2bJ0/P7W27DMkjTyS8ugTaDHuw2pvRsfpyB82h9nKx/u798j
hKZyjeBYzZJ5OHN1VmAOeLX+TTFNmq4Hg4T4e70OOm51j8/Sbjgm0uJ5Jh47CHmw9QrI1uigp4pP
m8XDz7uQ2j+D8J/yLJBfwxDDf/+/iWVo8Kgxu0BQxs23JFxRDpeJDtaifZoe5icnXRBhdv80gdA9
KWUXjRKKHy8jnxqFJOKHocVmtxuhrPxYNhrmMU9q6awImetmoNSdodcVnqMwb32zr122Vs3wG4oR
GG5D28qKSVr862oTvvCMdcUN8A/vjd1SWuqKMkjWXr0BnYRitrB6LVtWw5o9+k1m5aj9RjR9OKdP
UIPfH0b97USdz224cBtJESUciwZ1RwJE5l4bWhbi+9Tl4VKHKVZ9i1W+puPhNZrY83ch3R33Ti20
tFTo8v0l4ODR2DH+qKOnmKTmH0/xBlu+UY+QQlu+vqahQpMRDZlClfHfoq/fGeL7y1vRDRUM/u/i
WqO2GT7jG+auv0BMUw1vFOwsNOKAVXt8GdwQFR2X1LDIeNb/eDUdYqZBUcfFPekIGv6UsT959YJJ
kf9wPFmS8b6Jq3C3Dc3ZdLpcjoYkTYMPEMz5o8+z8OlxF00GGWIYuZJbErOiFw5phMElvTxzDE9h
44ZTCyYChfCKBQZLWvXGyhZ0YuYBPrNepKbg9UUicFAfnx4xslFEF5s7ABcZcuey+4Fql8zNZwCF
l+q+sBYYseUF+1i/eX1P73sfamzLaufeBpOKbKCYGK6EhQt4qP3qR0r9R6YJbmRK228GLXTYgp8J
WJuj+tBsnDCi5s9NEI2W1rFGayob/mFM87pK7aTK0JndbiyhFrFZ9gBhiklWsK+sqmXaUndwzCKN
5gAotw3poAu3h4EA5vMS5Hc0zBK+VmPFwGxqhHwq7C1tXUeoBamuMP9xq2mpR0mGkRcKkWcYgyNY
l3wEr+15oPdHI0jARgP4X/AzRk329nv80Xm0mW5Ef1sHA9MDIevitAhP1PHvoeTuUEPBmTbowrLB
AFMn3zOlxAlqi/toffU5Mxr33Ppw4Mm2Icre36yiDpdUh5xhflIo0oxq3jsFPswISC14o8OMuadC
uoTfZD9BJ1+jKiyCA7u4STb5aAckrJdgOA2jGgoiSF4WiGMkvCx3Eg45S6VESI4lIaZNuNI2+5CI
+hQpbSScNlGgYqEcHipclU6uRXJc5+yji0b7OpctpY32ozMx3+cA7iW+MpjhAVQ1/fLELNQyI2C2
G3/4LqGOYdoxTOCojUxwWEf/ZOIFvgSe72lqHMkL94oa7SeI0dZd3pUh20W/3/Up8j73pEONJllY
CsDrCxFhoVs56ofx9esu3AIf0zNKAX6Dlk1KdYaLarUSXPi7cAujNHEbmqnRs+JjJHswdVOckAf3
GON08nJPPuy3Un2J1bgq6OkYBFwU9rQWazFpfSGYBAzGbU6HjwPD3V/vDFUub+oJwzUNHrNW1hHH
qmNGJTlZo3X30yQ+rXGQPoey8n6B1v8oBjCy5wC5L0TY+btdRpSyGy9QVyyGtO6TTLqs1lxQaMUZ
NIOS5ECHaqvr7HJaXgD139lBJ5kQ22+GQtsuoM1ymhAVdiSv3tCnL+5gBE1v1QW+Q51rc3cBReGa
P2rdkedaFOCuNq9Tie3fQAOUWmjKQMlCYE9K/PU2QTIaZj5mKQoAot+aTPDjBabTFhBDHfQkZQ+p
2N0lKT2bghd2aSLWVR/jKAge2tOBnqnDCTvhv/SDE/82sm/QJkQSjVzXXkbTalEG24W8Y3i0341s
b6LWtKaYajvuyvoZWRqqwLUfIwOdSOOK7zAhsUNHxTSgcYInSAqAbNDnnXLz1vTflFtSm5Unxp4s
XTlq2YJ4cyHqGIayxg7unrsDrmrr/gmqIFdu8IHP7tA2ZM68Hu2Us2Ysyh6fbRRDb3CLKl71YjpO
Sv6Q4bLAsMsL3UG6d/7VqR71v1j1kNbgY+BVe9Az+xifb/QzBMu2pT03GWQWDGRzOmuFB7RfRO81
Lbi4E70YOm6tqmED4oVMbHCAdrzdfvrSA56/hmf0OrWq1jFYdVcUtIq/3KdjeHeqQhKd8n0tGNv8
v9+n6+BuP9sFWOi92feV+VDZhIbbWSbZH02seYZpgWqc/9MKJYmN6/JRlZVBx2fcS7axJumyEmAw
3dFgB0oVNrHpWG1jDJKkqSBX/cE4urqmYWM6VERVKATf/lvDkksnT6Ycuh6Gn04zniFcI1ICxZDR
5AEaO1SGwqdciVWpH3tLmzHKtYAIb3vNKZCp+TYLMnc2FozZ6Bs3f1zuzwabhRYP6otBU4OuIA3g
UAjAJfdmxYiZYtj1qR0I4ZN8n6EU2o9TsxWZMlQLSyIGKOHEBxHF2pVg5zmOoRSq3v+XSLBe4+o/
Er//9QuJpvx4hrCLm2XS3nyDQVl5iK7W827jMKizMII+fou5rDCKiB++rZ5rVI60Pl9qUK7s0qlc
2JLgRxFzhnQcx7iGycOIyiko9cjZt0r+BXhi1RhTzBaOsZ2cpmlxdEhzRllhfAawD+q5hFWfS9Qm
Zw/CC+2nGAn4R8krm28iQXOb5la65pdnG7d6JnGUP1YwQI79PIbC0TXqyEPtpFIZfsg4tNPyhV6q
05Thwkg1oiz05yTRwd1zwa9/tbi+wLsKwmGNAax0ji0hszAeRGgvoeZ4YZec2rod3h6Ux3iJvRSz
NI2bJv+LTq4IMgMcnGTwao2iYst7sCjCyQmkxEgdduWm9XoxlCfsR0ReeTZvZ//d9AmzEfbQAsv/
BHq/al4VHL1cXEf9ptwflCP5KzS2yKwwsvUgl1TaFW80o+yD+ksIArIFsrPdc2McW6uklQFT1sr9
QeAv+D0xEq4aMRG2x/tNWvI0FMtcKVFXWlr/SkGlQ3Qu1bgzPNbavA4M03Os66pp4B2MB7i0EyYN
gtz7mMETAdLtjXhhlEMvwOnSGenptkVVCMtYR3Dls/P5PAmjKlQAE/5QnATsRHpfD+04KzDFcHxy
FMCymYfbPuRfiAzTZpnDS6OmqtOSNiO6EfbUtDVoAHwU90SYIkxdtl1UkFLEHLJqMckVJ8CTKZmm
k/QbaUtciWJtjmuu6i9sAgczeoOfqXhm1g0OMT/p7YvYsDmqQCRHS295c4+L2w1g8e35t6tW2CuF
d1i/BTuY8r/uMnhdVyX+mZT+v1+dm8w4aB3mCUdfSGRXRFpmHiCzMFPtDqSp9bKE3Ri3BhI5tvCP
slbGyULgA5GV5o8k4JQenyETYstZgOqi/TUv/IeVLMYqI1+C7WoRokMH3+oL8235w5q4nqCdPvoY
gSGEcXyYi8XqI0sIH9F2KnRAOONgwS8KwBdd9IZa85pxcbwySaW8WHSnSVf96+ZrjA4YQ9unzo8u
0xCf3dHEAvdhAFpSWK53/cUkSgpn5Cf57CtTBk7jZD09r2g+DujQ3fAjEZjeX6U2ZqpwQ8FPoVPB
DMHSIWqdVszNPFr0KC6nrWPq93pOCjfhHFPSPAN3TvhVYZeeVM0+bRmpyoR8dRzTpo/od1kwN9Og
tWDMin/Vc8LKInzPol2h8x9/uvt5IY7nS90ycfrZD5bL2IDMwNl2wGg8nvYErm4c0l/yZ3LsjHmX
/lfkvSkGjOYjxeYn0cOTKbeviFMdlTGKAupORri85lADMVOTfrr1PUr2CMxAkgBgPv/oO+mtw9WO
4KfPfZIxc+GkKHJ0Yko06kpt6jHIYszEHJGzDv/VlUEmBE9KyhDWH+9v2Qys59a7uPPC1Cz1nnuH
Qbl7GbNEiPZOXfeo94N56doy+2MItWbpgQVgNyCn84eB89Rrvo00/Y3Kx/NX4nBxWximx9xIDuZD
sF0Moktr8zgoqKPt9gM7ZeL1P91jd89diBzwG77YFtMGBEwygkkz8QrPcJruEgVEWOZvFsfYm1lz
5RuhYj1DIxr9HlJfF0d9GPrvo2DeCHQIC4r2rPkVF8zxYGeT7qMYdkd60Iq/I9kzAxJMFEPLgzvF
1Rwiirmxi+0GhF422SLdsG8kb7peuby4Gr7tMLSC/bQbJS03sD2qfjZ0cMLhydtEmdP1zIdkLdz5
h8FuOTgu9xxQig/pk4iPAz1rFBk9ua9oXTPQL6TCADLmXIaM1Mcdy5YcNS2z/SoO5F+0KDRh2yef
hTXw4aDhrlFUkd8LjFkIMvRXgB3q7vxZ5PPrAE+r0S5FKmNYAMejUQimIgbkvsonRA46iLorKxnJ
s4ANDX2FWkpjHNCc8PX68eQ18Jt3gkUlU8jVpd3grl+O3Jqj07veRb4kmaCSbsv7QLthBMxRkmA6
ZntsLyDdO7VzZDFNP004zMZSZKp/p/GnXmRdnYILyrbyofcDHnaRI2QatPxFNMB1Mvilx18KRI50
NMwOpGE/HqSk0W+4IHbScmX6dP6p2HJhKLa7C9C8cm/cCS+DTKogmd/bP/uucY/r8qJlKrW80XKL
cUVdqkBjAyayqI86XRtj8SaGCPYqeqLYQBClt4mQYMeL4S1kc/nzxL+k8Q6ub7FHPrUzoBH9fQ/L
iexJX00Xh+meWCvsiMGecw2WbzMnTWiNxgyR17iPb5lG+p1ede7uq3tY/Zrup5u1MLQkkgF++LNU
zkUwlt8mo4weQ9OYt0h0VAjQd4/wj9LkxhgVOSt5ACYidl641eeg7ToD9tqGGhqT6d281nBRItD0
egLxCtHILgQJv3GwNRi/cAQlzJPEPNZdVk1wtgc11gUizcWJsQZFrkmOBDEq+tvL1DA9JdIiynXR
ZW7Hvr0v/EBwebuIVyhzWydsJwdCPZ414syY6z4H2ZKrX02FBOwN0G/IL/ptv8hBMBxHl3aorAQj
QX+322+icQ+jzM+baY3HtjO2nJGhocl/XFka2qQcNOkZ87sUV9F0D7tswlFW249Y76vLq1AzsX5h
n+zvMR5lYl0qI5pX0GoWqnnJIQwdK1HDNhtvLTQyyVaMFUbSgGPdiuRG8ivFSGZyUqmDPiGyzt3y
Ak0ixFkpoTbB349or3asFpP9fshRFWzoOZ7j1wGtlZZnaIit7fqrPA7cOv8TKkq4gyoG3tiCpx2c
34zrHkHq/1nVehi/YfjsuCwwFXKlcIybRir4KzyuSl/iOMbgIZr0wPDCy0WOP9rMRlEquCjjwI8g
jl3663fPK0GTeDtNEFDmGGRuPNnEGZFWiOt0IRRB62K17xFqbbaydQ0Y5OphHh8ZVHtWURb/ujtT
gT06N9vY5HQIAchp0AbQJwSpdGq59M1qDA5dZVPh/RTjj+jJr+9eB/XuD1G3140HAXcI2yWo90Hn
ISt4vR7pswuEtZq43ed31JyAoJL0GKZVo9V+rJRfxLczreXhStZY9wfEFYuqSc8K9xAum0rm4GVN
5guW+kCyBwPQ7V83y1w81vS6vZXrHvMWBLkzFUZ5rd6b6ev6K/WvVvz4YAN/WJmi+iiFcg57wyoy
nbF6/Qv90owpwFYNWEQXGJAl0hkL9WqGj/EjddvSUh2dcB1WxESfans9DI6tW+3higb+646sGvUC
KVfKBIwNTpccpJ3Mc29D9+pVznF6BCtHj0bh0fRUDWGLSU5BuXc3NDiAqQVlth6zDc5S2rHXrOZo
aBi+e88hgL603NaJZj1fa4u/AKl1qLcLYvn9Wkog7Jqd9OQhLH1cjGDwBspgcdXSvAuH9IaYmrmY
hZ++IYmF/8NtlxKnBXNvmBeYh3K6UWL9m37bbi76Ldqmcd9q5GPerGio4BRrZ2RjvXjAQzICfixX
9S97VCih+yvZK+w4VDbWZu5VYItqBC2Jq7Exas8dICIq646blZ9IHdWkcv1926BHHAL5ilLkatr9
4o8b1oTy6+DuhUfAi8vTf5F16fmSKd9vcgSt/poCL2JsgrlIeHzGJ3uE73XqjPz/4WQixHP7lEAF
4h1v6X8GDi0VLzDAfi6XrfQvbz/w34CliJa3yMN3IC79NivvfUdn2pFVRjf7tYgP4F0zkZeX1C7n
LahCkiCJRJKdsBoH7V80J5YKiMS48go8HD4nxnHtJtoflacJVo8K7fVzuJbkuyaXy1vr4i8i56US
9reIMWj9c3DPinQC+tWh4sRlfiKnlpCgDvQzUk/9T/PDyP7gYlQDCerfEPzosLbQoG3DC51rD+bf
L6rxJP+GZErYsXSmKEjAnvIyyTddQRZKBAN35C7W3DxKxDi6gpnFt59L0naCec6iwDhusnO1eXsi
TOmWzFOz0T9TJc5pL+Hrad6Cu7soeZ4nFFic+jD+CKoXzUFr1dPuqxMzRTYEYUk6xgeYfueJauDG
UKn4v/urhkZHHR50bd1l13uAcSoH02jQIHsNuIXF73cxX5xscF7OPz7ZMY4ojSTvmW8XmD9Ubo/O
LrCcPqBgMycbFl1fd8dHeAtVP8FoJUxaFA5g5n0PfOStqCE0DtQma4gJiBGhtmsrvPv6FpYkWTdQ
B2vejB/nBd5SdT0t8mUe0/f0xUqwtLzHixEZNzHge7MgAplLxMMvxu8odomzc/N1qJHqLw8Cv4CC
ywzRxSLGHVkBRDLl11GWAix2MSgpUiXLXmTTXpbsgKCU83KkjQP6DLGILDbV5ywb0Oj3tlNqobYr
tGiaOiqHHbrBd8+SiOh4AAgvZ3yVZzXSzUvUeNM8w6jMIgZl3WKjA4uSSmNA+6XW8YrhLtbUt+SW
Eb3kNFIM4kGvQGdOP5Y5XevGhrlyKZxGrvDw0jiulEOXt+ZAvVfaD0jFdwhbHD5OEGlcuesUJnWR
ygyLkl27wPMoE/qmwuMIvAhidCOQ0cfkSW8/AbagTcPv3zWJ0Iv3lZ/IfxzWi1kdoLmqQ+AM7wkT
+6ngv64VEj7B4avM9W897SQDfWDj46RvjnQqDZ/H7fivZN2Q5SYLB03cfx1GO2dKB6RldfAM9erf
3mhDcm9VYWtcwb2JGibqSdcQHRm4QFq1gwTYZMqthM9DHQHkDAcgIJgh15QXs6pybti7tKwAljW2
YrnhMVEYS1K+D9TIC+9/kxxFgU9bMgp59fNpOq2q8YEdLVT3cGPp2lKi2eKkLSUlriyibdph9Nli
ZF+eo/mJiXe8XZ+7ak3TB+iz6mwNthzOzB1NaT65A8B1Rj/4E5v/xD3HFNfssSTuOzJUHKBX5LhS
W10+9SA/icJd3Ep4RQ3IHbFqHAJWtqYuYEVOnQwTOytax06JL35quB6u/QmTA25tJmUpLwnEDpHO
WoFQFSgWeLizDwIXApTxuK7fMg/DINO/ysMqQUoQrtLTcv1ZGDTWqUdzVApve1+klJNJSZVKY9d3
YS7TT7KgiWSFmi+cokXzu1dLk+X4eL9O0ewwW1BfpsLM9dsfmOlYhfCfFUusb8UBTYWbu9GK1VP/
KEX+83y8lxBXOiHFmDGmeHEKYaFXRvAgW+uG8ET4RikEyWRo9PK3Hm4o2TQaQtDx8U/iAfPuhJiT
O5VFEN/L2WEufFS56ZA25+DBKqVElkvfh5LhiSKLEJ84gd3wHN8UECLY1UZIRT5l3FXXQjjI70Mk
Fd2Zp/4BogBjCrqgqsZWnc7JUgF6CWzoPZZUlHcMO6R8L40GLNMEO8vndihpNTpTIA7lG4Trslzy
7t4XOYkFHEaAhNnJoff7xnGaFt9N8KYzPPWwYtZkAWNXLi8+1YGSGZ7nxUpBcAMcxZBZt54wfxZc
WofJ5YGA/18bRknjsHZcJrJ8RFahGMNY5eBBKeroW9BlZFk4rf9hmQsF6Ifs3222VM8e3SasOu5B
Z6UXcIh0DoJVwRfMlZLU9yI9S6ky/F87oj7X9DFh0ZtYFk/4YcN3NTPbFeLeHEws97w9v0b2ajGX
WbNiwdhjFSuzfiF7DbIqp4HuwjfPc1vPkjDCNzTFev4pgQ6FYQ9RnqMELPZSAbsB1U8ZRpSdD5Rv
vV5E4QWdcmlzN5OO/vaKleURMVtQ7pDwCQU2EhXRarOr4ePzAFw0tpgJj9q4fQSZDPQ7YXGZfINN
NBpkarVMRV92otNJmGiWuJRRfq8FuUbvIlKrwXrIcxN0YlpwdlSIbOT1eUm7s8zyzGz0BC/JnEtB
PIs3G/p9hk5NbKrn7xtOblBOZwCAEii7TEpWofs3GhM+oci6tkJmT1e2A1zz4fcULo8rwYGuEsU1
xz9Zw4Fu4jXuXM8WUsSllqeya4EcQOwNYYtt6dqC+WE2NaVvCoL9YcWu0TYyJkeai3ZdyVG3xOvT
1VZcrbdhKeKj2TfdDARNxCZ5uhKanT9s4kF3MFa1kQwv3SVUdIyuk/fTjZhX8eMVAeRhdhcfvTDm
OfY4HzLXLTqTwdjjRz96LbHUFAKOns2cRxM5trTfws0yTv+zKl1sur25U3uQp94FAIMku8DG6x88
fEhloxTam0vhZflZXGo80pI/9/OJv53HPz8dC5kQIAsAIHZXt7wbyKc0xf8J0NC7BVXjHLMki5pX
lQ41KlogIZ2ndMHZNosc16FnymGEUTeq7sIiGl1OZAhk6T/5mZ7+E91yghqv1PbkEC2dEk2zuO+e
6WmzD/GpC24Bq3UJ/EaLW8twEeM2kxlOsVTnXiIGpzZxCyYIWOAACaAfnY7F0IHc33P+Er8FqjWS
oQ80cCqrUEA1F/Y7HOzwf9huchRVdDJoMpXNqxQe9zrcZt+FB3U8PVKFidrvEs6BtS3UP5h0TkK0
twgjKl1QEr/BuBQEl7B0ePALp6sUQS9cn3czLr/X9AjZ72e9s4mlG2jirBM4nqdXzBseVZL+m4oC
r6xMnz2DUFkGGNRQlwWyMQ8YZuwZCsGSVqL7tLVyPFzO/uc3QyZs1sRJ1YLd3NUTmz3Tc3r80wqe
7vTDal129fu+89y/J7edD0CX2Y0Lk3qZRh5QuZmLqvOF1+Q90Ygjfa5HhBFUWqoN+em0dyPmiYl8
eHYtgfpHTB9DvidxjT2kJPThEROd56fBRFe3qWrUPIKOybeE7sB689p3A6VjoYSgNvDPWz5j2D5T
ZrlWaaztW/2eP422XeMeW29ODPz8OUuScf9Os/Ehn6I/QKMIrUmCpYobfZHo9cXxZep6kSyGly8y
vm+6mLlhUNrmLgL4H7j6Qdc6MR7KzkFWZRcrOZKmRFX+foO4n4NXIMnIZtwRlzJ6zoaXsC0yeO/t
uMpgrVdOO47gNRLiyuRBrdPNgREuzN3fPKC8/HZ2EBWQN8HLgJ97RHIbZPU+Z/nDXj+lVdWlw8Z+
Sf2BUlSPR3AHgvo5xoZvCLVNuJnwlSp7dUcQyVsgadTA9IwDc4z18oqv8r1WgdwEUfRk9oMqGEYD
7hIhwqm3tPtCmy/xFjhQO67TEwJgeFuS5cI3EHlCfduW/lyeFE6+70ZBfdH/NtK67E+XNGLk2eZg
kk09dGocftQbTz+zFfD+kjIE/jHDFhgHy6dyIQXBCteQ0i53IRS6qsR0ujlFxMHTc9+51LS8hQCU
7j57JelGxlollxwL5j8VgXPZFjQCoHJMDK4PzCCib458oSyHlNka9lM4u+O+9P7cVmit5k58xCxw
/EC/LOoEWrNuuzyzyRWjoh6CxPqrrg5mxnYpF66GtDyQHiAzK108HvpHWua7rUogPD5Tict8Qeje
vB2OEolDqSyxDQQ3VvtS1AqaewTsgq/2bhDBGTQp+OSWE4xQO8TUr5zCiekdZ37/jkeaRcNcu0BT
qvtff61VLpESIBtQZ7Hcz0y3Qd24mPjByJFget48725QcKLpQpSaJe7TWoA9kvmjIZeLECl2BfMX
NCEosiY47ykPxA48+TL8C4bLM6UQQOE9Vs4NDoe/quWYeoNmgqtClBVO+hQtFMEXM55smS20xrDP
hBjCOOxccrNJo4K5oq4wdDLjrqFHwH/AshUyZh9RMENX6gaFokdoIY7sCBe6ICv7NBPhcl6mcQMX
3V40SaFrmJgidvdb8Zf3KuvvqFaPJiQWDgeEooE0E5xG+dv5opApngAvPV2F0uLxHXUWTYGcrR4m
jyP0ZY6b/RkyCvxOxVRb6Vy7OK6NVN0uCw68j/kEM6/TEj/NuqemOmSx6nQ5BQInNAgFYUL42Jx3
qjqzgGqKcpg6KCL/sswoOimVtMuiFt8nv+vpnuk1AVMjFmuTcPLlOhFHABwmsZX9SuJfNV+r6qM/
TKGXMnIec7UCIyqOkEwcrE/fZ/u38QIK91ogzoj2p6HbbJs7aGzbvzwiO/P2UAhWuHOggF3hToT6
qPGqbvzEKnshgJKquAqqhARBRzejNvFugb3TA7Zn/5mLiqTWsF/9kn6dig2zngMxsaIPzM2F/bpZ
t//KQZISprNvlioXhY3z7+pIUoVfeNbPRKXy6qt+roQvKQu9/Xs4oy7G8lTDEWoyiyXzpLPtov2t
5ydy3YXryVtQIQ3OAPMCULwt8JoE+yHBH+r1jHfXy5ELN0S1eOAB/xpyqdkuk989oglC6XjYhSXo
DbfYinA4SBPbdQesdv9vEctmGTgVCTxHgj+D+wZaqCoART4ayKlJ/muE6qEiiq9epQxCupdBQfGr
TjeV+p/xQmreZL7F7S9roheO1+pFCJaVac2TYxZV6b/jvFAnxuJv6BXDWlJBtqamLui3dRS1Sn7f
7SKqxsiexLJ/P5vj29Es9KnxKoWd+x+rK89SDwBGmhKxeCk+oPLqx6TK+2572t8BAFT/AAvpKEe1
NpGT5S77I5UnpngmPJEZ7GvTLJ0Zj+uHrwKKT4r2UkHIHMU5eJdXhVTx2FZyFi1nlQ6MEfyvkXpJ
2C/jh9oVASAGJeabYYQkdD/ZiVA2C2LNcTSZQvZTJht2xgWhiBpM2Sq4B6GcSbrif82sSmHywah8
Xxq1RC8sFRkCy5hzC8WffRmZ6lpcTMrBXoiFHG5CurcVCLkqwMwZbM1pr5nn3gQDRvdE7sUdOhuN
aH+YziGuFF3vnHPwkID4zkW7SrYG3KJGQ+B8Mq103kwBw/Q3NsovdEgZ5QJu/G4fWBuJ49fIbw38
17QpqdUXEOiRF7I+1Y8DziDskFxJm5a4hAP8NyrU+5x/wIWy7AdhU7JztjFpAJ/AkHHODcunLEZy
97iQOcZmL9n31ssL8wxo2GvHX6A3NbjcTbuKaTFETnr/AGf6M9sxZd8y3quE1mlAj9EMEDLwbU61
xLtw3b/5NHXN5w6vaIAwlG6W2FKNiZp1+iLWecxJrpZBeGhtYA1qLM0WFvL5Zc6WYfQ9qCZa5CNJ
Kxv3n1Eqob0+WJlgfxXH4xp7xPuUYcAntVv4oLR/moM3GE3ZcWlSMGdIORy4VnVjO+3CT79+PxuY
vghjlxzTuvs9tzjOXK98rhD/c2cklkb8b2hULD2GM6TVnhym8Q4lcL5S4ic/j+ylFc00FIbC6PEG
yDN8TwuDSSgzt7mA9tEeyNekNjWP7GHHasp/B/YMUzBgM0j42uupbGn95LmPQy/ER55xT5dGqx63
DeupZtUJpIbWSuG/48RN6r2mAGEP8nf2mAeCvt5XknAQdH1QSDmoJOxdvstZHk27RRCqeWlUa5hG
mvoTiEUmtBLLS1yahC/+VuIZ7gIijp/UKtk5++0MHJI3RQxcTPuVCM/elcVpJ4rWRpGXiNxgXCPD
ZtO5UC31oDWcnYDp3o/ae/GPOo7hU06fYk1uNyaW1N87GxN4sUzVi54oXSRXU50fzqCyT61+sNif
cEcVYn0/aXrpHPNS8MpAGZTqTNYRNhcnL5CuybwCGjwxGFajjV+W5CGq9+PwqJDw/WF2qHjW+PRg
hjUT1Ztyg0s6G2XI1u6eB16IWcx4TPJCFnKxcIB39c9BHUW2tKJsihPkNbHNfghsKVgD5uHHZkRP
qxKn6n7IZsxw+mnk0Of+0XwJjuIQWt8yqAt0yGpwk7RoTcovhGBqLTzjGHG05cBCv2xjMrHovLVp
Flc4MBdjafaNX+ThrLpPoGvoR75TitAg4J3FBBtj7v+T/wRNm3DM/lAbyHBmt3dlQECJo0T3hKFN
kxup7nHc9xl4fZniWtDpUsN6lsZTkbHSRwsOa9OWmLASeOYTJ6i+NVEG7XWhCsBIHSJQkddAUZO+
XwbExsS2D66haGV0In1WVMUDISBWQ17KoG6fX04QtSyzCxEdUtVJb5LMnPHZP0v0G8lsKwDCPqa3
NnouUTi1pgYlKXEcpxPV4zkOrDcuJTLqT1vb+ZaxUEIOyDn6Kr+LP51rGlXFouJxJDTjvDsouCji
6ZU3WdEwLxuykKQoaopQaemeHa8bLbIjvnXaYSJWhAJV68Vt81ZpUiEhV2rU6GjjVKoXWQ/UtGwY
AAJ5Y16jj4/FiH/IxnUiuGin4ICNs3ahlSZYIsA67hpGDMSWcMpSq+LyodLW3Tbi1yCS8gaUCwnp
W1CnnR4cieygbZOzRs5F6n7DYtSvqBkihzkIuiL1N2MQSZ2ZAzgrteacH4g80eu1O+ZFcSc8VFzQ
PE6RscNONgjw+ide/kIbI1Aws3wQ74GW543L/KhjRyGqxNVKXLFgzOInxLxgw6YbOZV/6CetK7Z1
B/A6HvO6ZnY/jtJ+AGPZ/iMTmy0becJ+a9kfUAvz0gmTc4DK5H3nNZGqH0T0RwQoowonrNEqVwSh
mru1riIi4WKASNyW2CC/TA/mDpgri2okp3U8Dl2k8IKic43Kj+BTm5z6zT/yAj1Kk52ejr59YWbm
VDNC4Wy7MJa6HCEUBondIgy3ok4srYQMsfOBToY3GQcBvHwWyWRtz95Bx+JJViNPIgoBxy4dYg4i
rDdKUNbhWCQAzLjZeySdoeaZ92SVaLw4RqCNnA8SyahnaxRk6/Y13db1NIyK22zP7BTFAsT9e1px
KkhjhMD38BhaeuL6ad7RxyFOAiZTNifVFE7P+pZB+0guaBowSv2XC805AVvLTcK7BBBHGbRuXtFE
SFQrSVXKAfq9JJZvaCCFgQ4lVRf6xBEZLPvBzTK3jnAaTT8d5SUTPYz6u2ikQeo+h+hQwAOrSHHQ
0ZgaYUjUaQwvuQ2d3FH2qLEn+b+VttzBo4MeZK1ftqSGhFzwZiRDBelJA42SogjxyJ92+11LXFuO
ErdVu2Wntird7RkNyQn8p9/ZrHUBeMJNqiU1dLMrLHr9yoZnM4ZxmHdiqNCPDpL6nVdJSd173179
buvtj6Gc9HkMpmTlgsd3oAvqdbFW64EeGVJJM4qIHyAWpTUvODPLgfM5VGKn2PwEpPGJdDAyQflo
Ga07YfGe/5pJwrl66CuyRuRBzI7QlUOnDmHM7euXf8qJMstkL9Dqi9yb7Ui2uNWMkyB+8gZMBR/7
Efarw3ivXJ0eTTlIYYNCVaBsxu1d+rrgxYASm5jQ6ZDAiSnU2BCyCLa2+CzaI5+LiMLuZ+o9L0vs
iah2a/lNLsVpCXNTKtW3eKRqH00UfJtZhNT16rhz5fYe97tO5JlqvhdevBwL/w44eqkzc7o7mpHC
R73hRR5m+9JSQ+yn4Ti3LsUizp6qWjROBcRIkXU9iX8CfmXO5av4sC5wuBxAQHTU9aYmG7Tdz4/y
N/c4xXkJS54K6vjpB+w2kqE4JyYUi1iP3RCPx82EW5aPdrlVbpbJntIuXQ1N3WkqoLUjZxnhVSRN
JOYVgBL3Rf0E3IJOs3HK8h8g4wvVtdB6Jv5fQYHO8SVWJ/judJookhX4MkxHmQ1F6H1ypqKpef0N
6rlZKg68I5zJXzNuvOl7URkvthyMC62COahd2MhIwAmNEkCcjEOhAsliVCq6cGJvAIQTisukegpK
hq6lRNgQMFoo3aL1KWHgPn0qRHIBhjy0qaTcptaTJHN6czv4wDKZg2uShUlRJS8kQKdOSz+Ht5Jb
4w+zauD9IF5lQVdWwr+k0C+xwFDQ9XPOGNsv7ADG4Ofe+Ov67PZ1C55/OZqThwTzpmrDkvPM6J6C
rBJBI632Boaru1MRbQyJz90s/FAVMMgSanNJillahC5yu/qWbsE1J0OltF3NghZnXT5p+JC+a2sf
kCUdUTXzfuCIPemweyXmmRVHUhcDQ/6xL3IgB2CKrQQyleURyhQK4Qu9tKcWAKPKGLmTRyqJC51n
Mtjv5QBjw22NQanNCZORUZvcb3pjEWTY3mH+WJTFRwCR+jw93wBPwwH4ifrsaSvVXMri1Xi5KvtG
Vn3yVvKJIP+zBynG68M5PVMMvt4vRP60dv9YN3807zfAe9H9NP6ffameRrWxcvCJBgZa0p1ckxMn
+4lizNkPleypXTJVz/iGboPeS5C6LkhXYeLsC5aLsiAFNSS/NccYQzS1u/MAv9tAC4ltPU6NH8b/
JDju+101Um5nWds7xjHLA59vgplE/Iqiu7U1YTrABpvdnSSCpOqOSwtWjF6o8/W5cTCp5bXp7IfR
hy+y89E5L6xuB1vU5FgOFRWFJwiFVITWa/kKT9wURZ+ZP42HuEPBdld/hPecgkDMM/WuDVp9ojdr
RetmBEZ4yp49Ln3WA+lTabObOfnm8yqYwHhb6bqsPcPT5pHZxvauxJvm0Gf3ukb3lcSi+NQgngZf
0cztQ20dq96BCBDyzTtxADPW8itgbLI33CueZCy8leJ2MxXyPQbT/THivm0rJoikU7L98QwV81nw
3/VsH/QXo9Tcglw5L+pTzL6dZ1gwUSHtDREeWd0mGEC//PFH67oQ6T+tp4bdOM+i9YC0q9eZBgGP
OO6MwTcuXOIq9T/CruH7LIrOmiY2SPDuRK3q5C/LyC11OFWf7zxdyvHUCoI0wlZKGklfyysY0l19
OGvfqdaf7Fj8sn+MfAmtuO+bpAv9hh5BiCloTildmVCcIUBq0MmgY3DtxjWpAd+HqCKfXsUDNLkZ
5Hd5M3aKn8wHRtcS9ZaQ/PJch66xj/MpYGjfhsPRefaxJjdi5wHp4/Jt6+WeuZGuqdPZoOA9DpL5
xif6ZcyI6EpBphu5BBkn9t8EVO4JaFUFitBOBPpdxXYr/PD6NVosNc9t1gTJdvLSMcEcTUmv+L4h
E1aEtMozEk7qBWcZthucthUL29PXHqMXeD/b9ZiAFEiyGxRFDasOhU+CKFrRnNZOApnw0eBhg6bK
cXygYbH47PZJL958cUbJIaWgRrEeGobf1EssQrXxSkLW0SJ66/Pd8izZTVnt5cHYqaACVxSwUQcr
eC/xjZ/BpcdYnb442AX8MGE9Liii40TtwDEljfNbzBguHcVf52etMoP2giLk8UjUOVwrAqCCeC6H
KeSx+72lMcBDHtZxT1BIpCQos0EqXSDBlqTKk3BQ9PL8cNjnmNJ6dx4qF871/vrNHDIw/OqzIDzd
O/litpZE1gaFbDk7T22GZ6lXPZvdKWEbuNSy8R007pR0VY6qTFo/6s2u3f0UoNfx5Yc+Ufwg7AS6
NIBI+siQs2aQKC97nXvpkJllgGG/6F5vo8baM3H3W3XnSB/uRItXNf+EIz8qOBj1tUWw8riOekRS
BqrIYjAKLor6o7HraJ5kzeYRV6T0yBaZN7hmfpz17mT23Xol4ePUVm4ZUoH21JdQMO9r58BWk+dY
7XR841Ht7162gMaq06C74fY4wVGlqT9dJ+CwonpoYMg8WVqkMAfsxxbHtdZkOkWJ+78W/AnW6Pze
U4N31eugtU4dnalMHkvHHKTn/5wkrD39pBQ1NA6SdkFvGKu9LpNTcEsFtFWTQbmAiCj4MoCnGTnN
u/C+VntEm5F6eGVPUHkMxF1yhf/IcutI9kZaBWbifS8kGMFXRWjZaJ4LtA8acQ9ne80aj/mJoslC
0TGgiCiDNpjosVg8OQIW4yLHBLL5VZF5nCgShQuX2nc563exqgZKtco/nLO/LHjONZY/9jPiPWkl
xHJTt6IUH5/NseLfdnl7/NS5n63nS+fyzpDGYZbIdSzQ1tyVVqiIo5AqjrSIM5QxIwyyiV/MGkyy
CwqnDToOgT3J09za2847ZVlSfwOoQWcM8LkRbWO5KQ0iZ2Yk2zoiS+1A7kfAT9FGFj0u5VDR7b/a
yuEEq4caUjgQjWe5AHvWdFm3UAQInT4rLb5AfeVVK6iy4aAIAaLe9csIRRotZZ4FaJIRG0dAygSW
0JoFcplJTggTK3W0TNuShM5eT43Btu6+iFt7icNr6f3mVqY77FppXfSg4FFFzwfvQnLuOsqjjhQ7
gVtzBuM+fFtTFO5RT0Bbk5QYcj8qau0SvNUonPsUNrsAW2vwzUNL8evhfdyJLcPuXSwN7GevjrEw
TJzSYiQKER/By0RA/IU1KcZ37bnOyxkXJDY4RdD8i+Q2DCNwlQm4UEsHE1pSMykGDgNmugSK8bhl
PNC/Csong/cBEga1dIjjdg7a2yx8gpRcL6gbB4pD2pXvcdLuKbKj8eADyco3BbtEE+mvBCFvaueG
ZGZE6rryl3L3PMd3GQPTwfmM1TCX3aNdMU1oQ080YYVkBGIyCXhfA9mJ8fG3scX4sGyM8JrP/Z69
3r3lfrLXNaKvXJGzuf+72kxBYaESPbSTYFAXVYlvvnkaXpGVCK20wjP1h6cLRRp0yXg+ZgUFOKSm
1459zZ4LpvYapRB7mDvMFX+q4gwrXp7YWdm1BkosyEiNrNq/VZ86AW1dJhhTS9UqEfo/A3KzoWGv
NHRSAMw2E1oTKGpobV9OKQyVw8AyU3q+9VkeN8ceRcreZS4EAPABhQXx3uzidh4PxH0oskJJJjxx
1TjhxiEKJ71JsQzSaGXifFPTlp13vlqwU0r5wlKpJA8PIIvXVk/rH5A6KNjjjlj4UDFfHNoott62
pjgMUdYYfm2b9v6K+XTKWOsIYtOzcMi8c6XDTM2VqCaz4A2GSDOp8f8VCImy7xGzRaQuflYbL64C
9w9Hdq3untoSL6Eg7PZlK50pKx6FCksyzB6i43vDp43QBwFvcN73y7KziTVAARNWsZC/kusDAHTx
BcqEWO28BNINKnS8ykaPd1/9uRn6xkqNg/PY11je7X4HTwaHNf1Lj/wfCNxlDNiGSkt89z4y2M5E
NXM8JPbutDMcknMmLMGJ+SlpCjnuY7jsq3vRLDziz0wiJf/i4kRzkg87JUwFC0y3VH7VtIvvUzpA
wykJADQsT6e2enZVN+bcKXs+VyJAqUEVrmFxJoZvxaTT6ILAn+ls1fVy4EFjlhcu+GvmX1auT4G/
AsOTBsIXIwXB76Y+uQTz9ZoeMNFxVF0WlRbEfZG9dzy1eySE2DbaFO6PQCsEPol79rhbN73t7adj
WkEfpij1IVzMva3d3RhpjukKi0Bwg7UCN2r/qMspFcx4Ti62QQaTeDDF8nSSxLsEdCpLobKgjf7v
TwZNaViUu2a65v8UO6a08XzG3cCCrBRyDRdFyKkQzaRDh0AntTbSj0PPD+vX5+kyaj5KEEHM+nLm
I58Fp/kbEkjfAyaCFFo9NC6YQp5MlMwe7UJLB8f9oubhTspJxBWU12KqQfJfO7n693ZXu9qrX5Pi
hIz5ZexZM8oDGPe1wwCU+FfYWv+Ia1qXMBPQhImqL+5KlUdnbSYaMhr77zVyd3vt5FP/ZANWkrhw
OXWY5vHK64pP7kgMc0+bl3+mQiw8KA3otOjJmJP04ld2NEUJoEbTfg9t3iQgM3ewI9TNecl4QVyW
UIveGsqHINPD7te4MxLYC+A6/QULy+hvGWrDZZAJ2x58H17bpadAG3RdFQv6Z+T9F0Cv3oCFiKwi
dmSeUhvLTB6fUn6tID1tOiIEk48mLoAlQn5qW/WD1VJMZK8CJtIbO8SmG/N6io1JRgmhjXrYizig
TvT35qI+0Fua396tZt2XOE8PCALainHZiRmqCHtfdilK7Uu6Lpcmti0qzkQ8LthMSzWdm5EUm24q
ctBaNKegLKSt6goTV47bWKON2qfmwpQhEIJr+myHWevN5Jb1sUWq5cYh6J3lP2z2N7WusI0kNJvz
WMKlMIMyFe57fb5e8YigDoOFW4JAk1pXZZ5j30tH45lzjpFj1pRAkO0j6HWpBybhAXf56G3ivvdx
35nvKMytOAMo1wUvS+Zn+Wi0692uTo31lncwdYEqVCu/RY/sg37RFZLHLau16egF8usi7jXg8l92
+W/KPJDYW3oo9A+5vziNmWGUJWN+S+1ogvbIBpHOkTgDYdE5ijHu8J3PNabdbx8ijEBEbYltr0jc
mC2FJh4PwJdbHdPmq1nH+1qC9bbmspePkvOp/PD6cRFQGgfZSr0rFUBPro2bFHXxFKgXcSx/+Fxq
r+ON0hK6qBhCCDuutVgmJCo14Q6hNGanDiTM8NnOiM/qpjti+H2ZBJQjr6eW9jIHv9Cp3+1YpTcs
h9cjuLga2h9N2MrEVI0icKX6hcNrwzg4q8uB9KdknxtJhvdWK3EmBdg+T3FQmdln+3Gc2RWQNb9d
uArUSHHciNMcQVlet7XNO5y1w+YYYZbAVKgzMqiwvQZuUtKTJDT6N4/b7YG9uh+Ks1ic3Micm49M
dq0zKXMs2Rs4WxWv44MJO4zpxqkdzFqgzGfOlSVq7EeLh0hgMx7jtz4XH+j+ZVpoGn9TP/rCXlHN
ocWq1Px5yal0XdeJj4sJJksQooHf13hj5ZqSaUod9ilDSEBhXm4mW+vCpzWzS7rMV0p7Doin5SDT
g+tnMoC+La5UUlCaKU1qyDD4hoihu7oRXq7UhlnHLUQXGB9ul7EeRMnXxQu/QjmW6N8xiksJfugt
TkTIkjjtkIfRVIX4lvryRE+WRmKfXldz9JMCsjw1LKuJ6Puf6UQjfS/RumOADDPmd3iMigxSugz/
PZApbjdRcI95aSvymN5qLFiSajY51O6sDG4VMWE5KxPzc+lkrIATTajTS8z74dZqkOv72DNeJYmk
ocpgdRN7+T1Iha8XtfRTKF44EKSGigCp9eHpP4g/dT4AY08WR1HKh5uIfB72LeeKFUOVrrY1nn/m
VU9TY9nYqizEteMcdc2kOVztxtOFWq73cb/fDivOsBWpD0SfvFfvhfF5OgaloHZvVapCjArc3BeS
uZhrA1edG45Zl6538BvIGQVzM/mzeSjO4DdCRP+qTsSNWAsoLGEXAqFiFBKMVoRf5fUgIil65+MA
EMTmkWTL+B95p/7O9rSEdHgbt1RPUWp0OH8FNnJRCZthkEVbQqKIPdtaa/PjV0vvFGmBqy/rib5S
ceny7ZzUNQ3/EPfrnubBf8SESkZQsEOPhmiwCebooMO58BsOA8DY0VvHLZUmHHzFQgz0Lli1MhxU
4F6f5WG5kYj6P3DRmHAlYYniKPycSnpUBTWP/QeEbz5lX050eYCxCZnI1lOEOSKmRb8O6emhFMXA
Hhs4C6GA9sNOovtemqt6VmX9TBalpo0GYEyZ8ASvCIhmqZOETjQPm29fN3gKGsZi66IeGGvHgT4q
rft0/5/EUM9Ow3cRdfTNBC6XAAcwyO9xsWMZA7SgMoxjwtrt3Kxzv2AvNgh3RwrdxSuP00+ohtC/
TkN5wUjBIeeVaKdnoO0CSvewmmf78wBI/4sRdH/5Pr+r4TU0BB3zNSq2OxA5EBCgtg7XJ0H7AAlk
5MmMxq3e6m6vzNBSfwGhxmtoiYSaQc19U2R37xT7L+2GmeYY6AIzHJEIU4+oMV7BnHNrJ5i66nw4
NthqHUo72xYrh0qyHjrQEW8MDy1rzyOD7wZa1GyrTxsLG/Mv7vPYHspFyYf9yo1eLGMLmnL62nrk
gRz2zna4ECB9h+cQtnjPHeOLxe9W/86BciBs2dXYooDGmle3q4pKqWOeDnL0TqN5dnHRik3KHj8h
XyNYktbUGPqEi9IWI/ipM9U+nx4rf44UxH4fB75UFwUZ6qfRm4VCBnM+PDKwJHnU+lTHvcuFtArE
38vgd5a7o7yJT0lrT90SX0qftC+e6QQpg8s4uypOC42xQpeAOzK0lpBaUwIpVYlKSmD9MSTBa6cu
FTnbCnl1n20BRAr9h6vnv9yO9q59j700br05G06QI3JXxS2BYUJl0oIHFnR4a4hb5zIaQSzavQuE
DRKTXKhe86kGxSRyLH7Cy5PrEwJje3KgsvyZglSyWWyw/5mE4JiWZ270/xVgaDfK9KNjhbss2dao
9eBJ7WgMoNZ80XrSsl3muFfsFRbkjwEy4BJGXVtyMH+C7d2OlVekSbecMM5jJZISpX3T5QqZ4Aw6
eVfkc6c00q0KJzenlXnLd/TgignIFggMQfCVu+bWRRBcMZbZEf90zFkcgZ8EpD/MwkkZY/bUoaOw
TPoClVIOTia3W7NIuQPknBHy9RfbQD9l4VgVv5O2sfUq0kNVTJRqLjEK/lc/e4VPLUufAQXlXYj6
y0q9l5f26FSi7fWa8pn3/VHqVH3fn+Zzi2f/Pmf1PYJx2UTRH9kRpDYYKOatS/jazXL85G1U6JDz
bY670Sbc0+cz951fEgfhqZ5H/4wHEoShpHS7r3u8VV0zK5TNLuUCRGgvGjuq+eGSX3XzyiMuNBbG
4HSdziAXkob4lZ80NF92EpbYbLobQkjk+SS50aRky4EpKid32yirAjYtf799QrI/ZZ396IwQNFO7
/s4xvBwRQQhwLY5xauQ3pwYNXkY2QHvNCTF6qKOmhhWFpsGbb+WMlj4qXUiCiplMSI7bdB0Xf+ZH
uto0FU+vCDy7Gv8tblv1+XqpjRD5+qQbAAvTHUHGhUA0cIRU63LbYKNQIpYjn618B5lnySz0t+V6
QCZExg3Vunq+B4EtibIQ1nMbbjb94w7CU3gKW3XyJ8cZroeyjzgyCTPiPP27FaK7nD52LSvt9dC7
OyIN5hyfi05pKfK7TAqtop2pMRgXNgoR8tWR5Dz9BrH5SRJ3aUVlmWlvtLBgOISgwcym9+tfFzxf
b/UVLB4rKkcciBFZIqTx8QOHJAWB4Fcg976juSDBol2OgKf3EYf21mupiN/8cDkFH/Pu0UXp2Tfw
05QUM7RQfBJGe6UQ0Il6kON4GQVLLH8tmba9J1UFOW5A99fMmfj7WzLjxSr77GkeLqjw8Z76fTpX
52+oV4SrJ/k1JfefUlyiVTA+tERBl1YyiWWZahr+h4mGfIbJTi+Sc3kEvThFCNFDLsCyZj0+aCGJ
u6QKjl3gRQVAK+dN8o3d1KyQnNZIFn6Qw2vXNb1dWkzk2DNJ3tkeEhLQ11GC6NtnijJhc6KmcLqJ
k3BhqUhz1ySV8wZRiB+XfhrRFUQJWnqKeg4xr/bXC0RMcpRoH9vj1pxNi0CyohELEI0+O3dABKVW
nHYn+Y8a02JqohD1FiBWqbC7Tynb4EB4w59aIq3J9whbPGZehe3AkmAqftvz/Yrw9ZKAih5eVffl
8xWuNmO/nxJ+9Q4W5zVYp0eIAWfXXTpVSn6O/XcxgBnIuvUsqF3k7jE+jeOG8dFENhltvsWQEt0N
yGGxO89DEl7XwEaojVBAqIaHONS8mwbRyD9fl2Hn5y0w8RqaZyW5vxmQlh3aMVkuMmbTJIkRFdJe
4cmjnompN0jvVMc5qK63z8H46CaaWscXGGlWvXnEfxmGxDqrng2E6xYWLdFdkrCiqj0FB5ChFH6h
GosdpX8mLnSbPvTnj+z5LU/F1z0NPZKjsUFk07yAjrVAJImbN4ryCvoiF+VbRsrVzGg9Ngs+YeNU
k7v3+iEvbE/VqjT48l0ZRGm9UhUOeaQVL7XAEWsZ21aWYDhkTccwnItFwXKbShz0ehp+kki3IEFR
5GlTQR0X3I1QuYxibmeFtwR32qE5+nmX0pY/cMZ1+UNoot7Udd8q6JCpb4fNJNUQIvXTL2pov+yO
YPJheI7tkO0F0wPXkCC4aOwsCduwGWIRLbORiX23tUGSKUfpxrThRhl05WlFBH8yD4X6ZBlEVzOu
w/omM/FkBGiu8NyAhjRE6iw2qcFYYwaVG22pdngjPHHn/9PuDk781aWa06SePwZYmbgUyU6g3Z/z
AOY1SL17C/vA9DUGIV6Nb7Fsz5TIDya6NVE+VbkeafuPW+NxS4wxDmWC09x6jSV0w0Zr12HXCdZl
Fcr4P5VoCwYGuAoKTFgcBhoBi5oY9ghkPPdG8hP8yC0fU80OJvSP6eF62y/TMfc8ZQIjoZzTmitQ
a/t+EnHdcibyhyyrTC4Mi8VmZ4+0bYHnovWVNyvOo+pjWwKR1nQi516pA0j+7sOUJ1p84wFNDep2
ItgmFix8u7By+wFKNHFq4Hgh+zYAyQBouQ+DxMBrp0XuTDv7z1jM4L97qMU/FNP3KsU+2WIGNLHi
CV5RNS90aeMLyzhrn0sxGsiHhVTnYZpD/whYjPVoTmoy4oIxG5XS7WmVGJPG058zSN82FueFE8PM
FpUCGMoT0PVUPRFH8DTr7UmwEnq3ytI1+z5Ge+Rst2pPJuLFN5i5G/LMTQ7AAc7sN7qjGmYAjXPt
xqpvkLrqRo9swva0DVHXFYsYxim156xLGSnQtBTxzoEAKf0umC7+IdQkgi/spga2cUK6Dq8SEZOs
48YH41oMG5+pLLuGEh0EhiRzEUWsiVSZhOhv7rJITQ/S8PHV1krOH/F+OJOxwtOySVihGmyY4fk0
oAenTQ6JSiDUTNAJZrt/pT5MiH0/f+y2cQEBlrJ7asAIkCj47zA1qGkb/kAS7S7dY8XXcVqPb/Ow
eCJM8MT22FNZp4KWwS60G/7n5DHySp4v7cLtUR2Z6Rj9uEl8KNJ9VZdm3FyoFfkbh2MoEmztYKtT
OSCPzEPKryNnYne5WI3KnEvPnyZurWIAxfmG9PoZnIvAofAb26IOqbxgryPdEiPdvC9DzXM5ycVI
D+t8bRuVDf0sa4AdgnZ6FB1qUd1VdZpGJ4qxvBX43kwDm2Gwchx1l337DklS6hMMHRw5lczaLXHa
2hCEKonbs0WF/fLVZjIgo7nQ+/k4be6W5E1zHXHzkrtnPs3g+yeABG9YJK6IbtxMDi79edY1uxB9
naTT5lfxthA1pQVciu8VT9vuSUZNCGdZ+INywRmC4tDnT8b3p3agE7dNK64/SdtOEl2R9eGQOxjU
9qQ5hi50EXdHrHnHr8KL7bI2JA6XupmLYeeuXlHrOXtJWj4EMEAo4AC1d0hp2PGnWOoh44di3hhA
ow2Zi1XD8hNUthDOroH7s7i+HZjBQLhMN61FobvLHyn3lxsUODA5aUXRPQIfS8LHZEURDdP+2OKy
PMgSDpuGoliopj7Bjt9FAa1MhIOLVUt71IN3ZQeLaj6S+Jts60JUdRWUL30usLiV/UpnIndqWao2
PAO6WUalFlCrFha4oLbv50ncJKdpeuQeNYbAfu4WUjTL8jmvIl1/NqQGMEUiAuoZDpYLrZMLq0UD
ZkuzMd5JbKUWe8zrDsI5c2ZapllHgeKb3/A+tZXGpYi/66EH5h1hEfdFaELzWR3bygJ4z1Agq94N
PI2zgTKnJxZrhh3hSAQpHD8F4atqHetX/Ldv6v39YcIsCOOAGnFDlF5Uuk68t72dn+BVavNzlcGw
shAHIBbi/hIioueGKYMxV+UE5H937buGetTtdgQaiML83gJwJ9SKAJydVemhE6r8Pdxi6uuXRljf
BASqfZlSjbkG7pvj3TgEO7XRoxGMD3B3oQxK0ZgWRjwIT4L1TGKXYC1UHN07pz3jGBlDJeGzFfha
IQnca01D0cnlFAidThbumwPQBckNlX5+hyWDZRao2GtMQNHsQYBkHtTFBJ4qSeSyY2K5LnIchrSu
uP6Ys5R2CWNwbNkxwhUFrCxY5Xs75y4nuCbzaca9TGs5Ipoq2zAQkKL0+Q9/AeQINjsRT4hTjYG+
GQMfjERuYGRfnnYcJdZiSR6puNbVkIRRjljKlD+YwqRfLWsujcJ17mGDFlbR1dEiopGcD0a210Qu
2QMmwDeO8S1PynNIROysG3yh+BH+ocpJUdgoo8qIE5c6ZHTXFmQFA3TscNX0hfq1zde5ORbhN2Qk
qagkd0pHgTQBp0Zx8Io4D29ll517l7pvK0BcGuBskhe3D49jC4b9MgJY7yK/t6ZgJX1k8eBAWj9l
B9A3pfkcLvd3ytmg5x7jxMdVf9QZhXMPqat4JUrtGrhl1OcGkK+tTQCsCoynJnUGGyBMvVL/brvO
UmbKbx6dwGxhhKKPJzbVBpo3SSRxm1+hKRMrwMlQOSgSnPB6QVpxnj9ymgt1EqhwDr6vOKiBMLu/
B/wBm3xcoEnvdieGSkTrpYJqXKcVtjDdohDY8QOggGcjzo/z4qI0xbyS9vm7iatbWMQ4RD9Tek2+
Q1sAYlUvxQq0/dp8HwIO4MWPNT+In2RRlifP6iJoGi9kSgKYVnzaH1NuqIvkP7OWoT0Wx7oMsizr
nf3xcJ1CwQyV9tddAnCoWghNIZgoztWmWat+S9PyETOqGJJ5nzUcfweqy2Rh+wPTCLWGzG/z2ho8
FTy4fAC/5ew9e6vZk7pPVONKtDYidc40RW5giqj5pLtnH6/LpH0QF5jHd3+lZUtRoNXOH8CtERjm
aDXY7UuBD0vBseGI1F1nK0Le4uxBz261bgvnDco7NbJG1nF5r+1m7JVyFai4EQplE9A8JRq1xpxC
k5DzxH8uNg7b4LHbWC7wSGnODEaguUIhYfQbdaxzQOt5lx3SCQ0eieoT1ZNu9pAPRS9bPSUsoGCj
YCXrc7HoYNnqtJGK7CFd9tG9ZY7JdH8GpGw4KDpyydZTsIsGWcd+lL2d1/JTqLKbLyZ0wjNA5wh/
XUonmwZRUig8UlEFYHQkWUGgLQxgiBwhOy4ZG+E39zEkhN4r/7uPRW24ZO90YmFE0224RzkdgCCH
F9NDLtQZPp7sm5SKAojcVdwdoFyBg2UPhr/W/gD9/cIzWK/zy9vIEEp0KzjN/GgokgOiiPPSy10u
SHgjb0C+IPIae7a1uQ1RTD2czAcw5PkWUxkTIi1Zijld3Z4X9j8n8i2Cldc/WYKzeogXRXm65KHQ
Vu6hLFB5zuSug+XpxdXYyuvjWx/gqFIDL1F/Tutf8gjLToV5qmWxHLIp2lCNUzgRbCN/bXnOpz2c
spyZt9piwCcziUOisEP1MsLL8feL1WStC5VpSoNbkYXOxxYNBMJ3gW1xGZOPvttXB5/0X+qAYCuo
P63D0TWPHZN8RN5LZ7nBSA8ta36Lj+1xzv7RzilJtGq7hXYLicdLMPBMFZzxv95UdlzfxfKzHkDI
5DcSGAKv9ayCubmYvjpbnthF4DVFuRnmd4Ny9CHH6+iZNh5Tj8DRLpSnxlwblCY9QSmTvYBW+xik
gU28s5Zaw5UxeCfZyDqEMKqDpTwgOp5zhVE6gg+vDCAtTmYP64OjhSz/Y/C+hCXlbLS4zzNA+rX0
50suE2cJ9o/RTrFRYFZgasQzQvmQxwdXTbOPWB0otFDOkqUZLpm5SMbrXYbzoJmz+OHgDyzcdeMk
Bn8/vL3sfIL0oH9DGKLg/KaSqWtmjKOoE5p6sp5ynj8TyQjvcpiIaifgjvYj2xHPNkQdXF7CCjN4
AvVVNOiyMzYWWSHfV5nRAkQUfKcSxhG6DcfJwNSXm1V8iDirHPC40BzTxsJRMiw8D08nhuvVX8fn
Y+tdA/6+/hn0pANCNGbJvng6ubpoYI4uszKH/j51DrHsJuq1E6lwOXMYtWbqXlPbUCukD5zc3QK0
i7vr2AM7zTFzJ8/G5ryRi1UCDiQ54iXBOR5QMrANdPWATnV7UkvRjIk72KjeCkm1dyGslZjgmFli
KogXS2dqvDaoxiJNB1mB6tau1TsDGEmApcXeyBDSzN5EANKoZsdkfEyPCw7TIaGtbgbDMuUIarWh
hmVKrhm+B0Vq5YWdArTAXvs5HTVsDzSuZIpLXJzNPeahz4XJe8HG9f92/s5X6DVJTPWBLxahH0t5
LHOqaivN3co4VHoclqZby1xUXdezivFJTjW6zCw2igZ0md5141AJbGrdL61vg2vfizWz0/IhiFhc
98sKR/eYfl+WjhuStmVjYKJtqbnnQX0M6Waazc3cjZ8R/ShA6CZRZ7sqd0S1Yd9aBOFpNIQc3wmV
udu04wWvMJ3UV1Z8+FFbyXPtR9Up4FtnHQo6KbF+qjWfRwfeb0cfWBIIpFPUb8SY1sGYGwm5vikc
+QOB43ErLVVkG6d8KaL7HWeWXEKz6A8FeiqEKz1ajGfVClwgbkZ40FtFQCRDCMhSvbz3DQAbfWmK
zpUo0qnKydk8zegfyWu/LrRZtvrl3Sg1iMFWloTPjE2CTSXPKIuHdfvDITa2V2LIEL75u9/lzE2K
ykddGfnpzYwrvGVBYOL0WtmsSL4KRggGonkXaDmYhnAn5HZuEVE+dmvRCMxyXccTyFh7H3pjGvBg
SGSgxARIp3ncMQTvpSZ+p0XpXvVUXtgql9cRf0GhgRRiOhPupIj3Tq/3DLY8v3YBM08UvT7Xf11r
GJlPXEewvGy8ldaSwWwZxnc/vX2DUa5Ggh0lzRCF2Hlu8ug8V8E5QbRt3wuVoc5m8KUitFej4MVf
lv3aoD0IM4Qsv1FYZcOJcBiWroHb2d6v9D5ywvhz9Vi8y8DiE5a44r+SDh7I8hAmW4fHKxgrZEVW
/CujrR4y4CRF6wp0qX5+20+9PD9kszBsRxNRtDw9XXI5TI0iaNrB85x3Y+tZY/thqWDTx62x0jns
onM/0lZqvgYL6NIEExbAik+r3tGFTO5BTrC+qzaneQAqQ99GCPZ5sspnPj3+XvRUNe9wIkLDTXBR
W04dcZ1vCTDLVYpcasUW5Ob7X+7jy0rP75Eu41jC3acdO3+wpMkr5MU/SZXaUC2aCzkTfXrCuo91
y2CyN80DQ/icHdsrSRaP8OE6VqcpMYn1/nbd36HSRrjZq08kBnZc+lkmlaP3Zo1YTAdrBaWDMyRl
MdaUb8dfu8hbak7TP47YKetB0E59Ztz0TK5j0Rai7Ax/rY83aBsmLh1umfr56BZ/QxbYIU/Y5tRl
85peV2qTJvBwJd2eMBpVKsvwQypFkK7jJCdl6J0OP0xajqxclCTFuC1+snVBhlnGZxhPiVFTTWoF
XEjT4HEgcv27IspC6ytHOrDjjWrEnqF9/zQxxY+Dg6zVTMvdwiizHi9ZHAPyji0Y46j1Rvlzf0nC
GoxOZm8Clgej3tygwFdwFo69SX7Ccq8l0+XpbwHIdMfuQ0dE5nVWNFP/3FX3A2txPRrFgQNkMiBM
vYH1mXQu3Rjjl46oGGHwMmLFskXBfd8Cs82QOkmwccX4c8YkOMuR/zqQiCdINPRgpG6sluD8Md1C
qZ2OuaemR/gJFsXRxA+TJX6u478s9mgaDj+BlJVfHg+RvRuE7JuiY2IrBtCDCjfnNmV6HlbIO8Ak
jueE+WiFIU109UCmWrGlM9cKg/En49eynOCc+jY9ZskoJgxGHS2lVxMiLrSgtwXBtTc0Ke7H/7Vv
lDb5+GDUZgZvrVFVHLT+Az6sjGrF+6Ej0d/o7ciMdsoTm5/YmOMQNclCKcm18JReEkiR9Owh2a7F
khxK36qfkYlN/ZWXX2uVB6KDW6e2OsDA+8I3lFhZu3tiqZF9dJLgCEnxEm4Fdlboe4ijTUCwBRBY
IofDDxMu4md182jUAnXsI3sITQYAYXEMGqcWN41Qx+uyG3EjfLhma0Ahi5O7U94E3pchu/S5gTHU
Qy3ha5BIH5hTXanuzYUisPpCvoMYbCalB+zsLIyEoHGpgcQhScSxWI7SkbVrWl+/tDi7yjPWtM7u
iP70sNAIeZj4XddUubFFkGEtzsN/5VgoCjTOKXmY0F66DkVi/LXnVC+qzXWO04rfHMy+uI1WzPij
fW543eCvI5u0Mog2WoL5ZA9rewat93zR5qgX1j9p4R0zZTEZNPtOsx3aj8rVaMDC5lES993v1AFc
k0sgFD91nI+AnSq39N1aNmz741YX1u3ajl41xeKaXxSdTDM4seQymLLaV4ogESMAZpxM4GN4hamW
xr01uauqKsrnQwPz1/vYcXssAI5Kd8bb7BqGoGWlT+4q8TyaDgHQb+wyBIXKT8V96dZvH/cZyJmm
+vaYoDGJ7VVNEgUNcr240C6cYNmK7pCS4qBAshh6NT4FEe0S1/kulvGVLTO6k4EaQVU/apdFdU91
OGQJNr7uNKgpbxdMwQeRLk6xmk4b4dvf6Xc2JINpkWrwfnhI3XYBwxh7hVkRYXBIf5bTYDjp6MLO
UR3wKioqeIJ1HcWRKSOIffoetNn5mnKckemnHuOUhlpyYBmla7QcDKuP7KDgQ9X7pYUdRs3BWA1O
oXTho7VTiBNSOsKgpruxQDhKCs0BRzHdQjkrVGdHdXYHUig/E4R0jM6hEwRxrlTqfIJrhGwJNg8I
7trTLlFyhQIhWBfzlLlgB0Z3fcdbeDaos+Dw4OD6599EmLB+2c+vVsh8e4ySciJxccKabtcAdd2d
tS4qB2x/LoD5RtjLZWR5PISMStPUxb3jePmdNoUwkta3NTxosyj/Zw+nkVFkyqwdiHl80Y2MbArP
zPOHqKdywynRalIu+SuRvBcuu+lkcEYQnncMf6GkyU2gkpommtXMSz2ZSZ60OTdzqK2DkiFbuvBq
EQoLShbthvXm0cVQOkvgGxTRxI0kKwmfEFTL7JT79RrSnfYM//30Fsei88Hjt9nYU7xMMBSilLwL
s2Qrfuy7yTY5tIdFy2oMWghQvlmxmaJ8HNOk3ip2C2P1UZtKwjDNo2XWP4jAsjsRieUF45XF0Qop
z4jz3WaRC0MvUiWtCozPQcoUenAFhOLFtu1JnC1FwA0G3wvpQqG0xiNjP7V0kQ2fx7An46bK/WQy
DZtp2qaNovh8lFvz97MUW+U2r9ncJLCOpK1pYfqCH04FBTdheyYUZdIyRBeOb3LjvVceCXwoV15H
h7u9/GhgeOlUC2pY7iqw3wG59ShncOwT+YOMsnGZINquxOEu+8eB4NAR3ZVkQeoiY6wzUzY/KkHX
o9309vpCaTx7kbK4FQ1u3zLKcm8QTK2Z2Kgrpsj3px+VtAjLf49qp+ZKO1zgDIdOQQ9IY/LUxUP0
559BbacfGB5tf5eNvRa9vnTBZaemfuvD/OqHtZ7UgMRiT4dSsafnlJymwg9hpith/J9rwSbwuhsP
DO43wINTNhw0ZA200vYDSRPZhi7C3oMDIEIB59hzeI/d+/aZp2hqtlmt9U9aWI/N7i9CtV0isQNh
bd69INSTuXwdX1PBHqJBQc47YE7leNqfXCtr5/8Djfl2VozNue70npFbKcuF0dx8m4pCjaPgV/RE
LsDvNUxdzf18nxVh5du/D5ykabPo8pVCKzQGuSVBWG3MubyPriEpUJ3ya3C7WD6APyxXTAYK71Bi
OH7h0i7WFZWxyppKx/Mqxa0QlSHc7neqQURc71IwBTzlBdaNj1aKcUZduIVJylt2t6Su1ItNlIqe
ntDyFtzsgg0/i7x1hLdh5nfM4NOu+zSGhcUePHo0iKtgGo54DiJJflMR4ahLuoCQytlt6HCnJEqj
zwcepD4sB6lhNRZjqRbMJw1I2QuIggn5pVMRxk62LAJR2hFR+zztdsvmqSIC7WIh0cycOG6x1bVh
tg5gCUG+TNB5sf0hMdufHCUp7wfEDqfzqLbzdP4ZZbNWdrg0AH6Oxga3HZMHBXv064wyugv+NqPs
tu0x1wRBhbmnWywz1Mjt9Iju524efs78DSLp8vKTqoWBQnTPNjALKDBqB0xVI+F4UIFM3OBCkfPR
UPhS8Jzob24+S5pWRDUIqx3RJocDqV2yPlROAgwsehMJQAT9i1K/HOdfGhj7R2w/V7RSKYVOkZN/
XcMjmUmBeJn8JLhnRJYtYbSoU4hh43y/JYZFPxRRQzhuhl7WXHTvys90iX4uG2urlsOcysew9cd6
A9So2ifvEADhrUeoTDCUvf21l3E4TI0oNvB3MQycjTeq6eMfq9zK7lh4/TUASeL/Ti2K0u9QAaKx
SaeQMsj37vA8AwV3e4iFaT96aIoRL/NmGCzIrJV/H6FY3/dFyQnG6Qu41u+a59sZ3htazpMGj/1X
y8ozXyYNpMBPqIhvmDh2LqGe/g8PC4CpQrI9XpUtWIVyGzQ9bZzXBaE6GTJ8x5QmaMKmGJ7za47I
sKWTSc5NEp5nMUa7m1PWLPA+zIXvOylxj2WV/aECTRr4AKc7viaH6m11QCvY3lTVdB3gxNUF01FM
tEDFUs03SDacZbpvuwwWIrw31ueLEM5sU0oxcAQ//C0ZtL6gUxkrzVFpOnwYRV2CmfgqojoRahom
Bx2qsra3rYSTxx/Ak1xlHN0jDSIYuwBuiURX98/wlkP4qBBAsP6rWVgLvVY8SlhE9ZtzIB3VNID1
T7KLfQGqkJQWutk+B6rzZrYcUBXzIV8Gn2HOjFFC7E52SRI6TbzOljpJQ7N8nTu5ONepdr73xe8K
plrdt3zgM+yWE0CcoHG6SbWzCAz9ktU8FnyolIVpTDZcFcpG32GlMU9AcQsHLvGI2PeLNJZPjBCz
82Y8lz0/BEiC3rcOdl+VZPUKOLYlnpzN/PcjDTyjrNWvrwND6shSOkbUJNh5scDr5eIDxy0IHwRX
yFSKLudrS6eoqYl8PDlqn+pmdCJBN3U1gjWbkhbTxF8aidY+x+pxWK6InWICB/70/RZkV4v0rtfh
j6IokHO73qJDOS+GmaPVLozq4GiSPtxQStMW+qek2EEOZ1Ox/0bzMBq/jLxycjF4k0vtLe73irRX
Y7RDdHnP9mRtTsrGvreIj9az6CXJSzwUs2x7jSz9RfkWX0KNVs3jCgx9q2BHkG7Eok697O1xCdzI
0Zp7cYHhIL7Th/vtYxMwfB90djCY1zmHa61PKZrBPTUg2DU/jmftIrNJp8PMhh/KSlQqO1yt4Dlm
zTYBrIIrfUqU0x7D3omSfFc/W+LaX3aozAmbhJlmTglCL30Oy91sqyYgKCZC4FoV8qQoZQ2wEz/N
RazuJDV8u2Ox2pQOljiRwTjxnZTBg/kp3eryoZPSvpu3rqLw4JNWEmXOWDkka1do2EwuEojrVYKq
k4e9Kk8T2gWdbnA+af8qtrds+mZRuydOnT9S6zimU3TLaB6wmUMupQHR7noiTZmhUlxBSSHzqV64
ef+mipUTBW1UZepUoOrwN9ozgV7g56QrE7oScns+OiLt7KSsqCHg6Hs7d6qgWnjwzgfBxrpMaf2l
dgghSMULVUC8UGjU9W1YnOLsl7v+iCMytADlPQxRHGILaqhZrNJfzjDVh/zAPLblZskL06SB+tm0
x87z6YbXWA60zqjAB/5B/NLLvJ1ceG1USeW6e9w8EQQAeNprlFhE5CxWCYxb51k3J2R0uRUMO6YS
rdtFWcwfhASs2Rw6c9jOsFFXkIjpkAiL/NRRCsTj1opTOAWg9eDRK2MLGbbGW4M6P/xTipaQiOZH
OKSU3Ze810FnQFBHQJN/OKzO7MEmNLgPLXrBa7/o/NsLscxQ3Mnwhvt/k+Jg/WPeDix097fk8vDN
JG0YjsN16J5cVkIqXmjnJvjReaZYnsK4BhMZWy38PolNmKjZmZ0AvBy4f+2Vr8cOHdUrz8ulZDDf
ZqO9X8VjwXUoG2Ly5MvhNwwz4rI3K7YJtk1C1TZGkKzC1sK+qfe3YBoH8vbRe/6LciiUQQ4TuUJQ
mQ90dPDa3FdVsS4HN8DViV0btEmmYv9l1sDS1/d6o95wXGPrvm70LKz178LHQ6Y2ad3wd41iRVxm
oT/BuYBdBGk8dF0ZVn2WJi5dZhyd09l/bq+zs9lpd7j7uCNyObjK0N3DKUTFhfYhjby/U9eXc0Uy
xLGRoEjdgxBHAau8TyT68i/mYQVy4qIsW0Qjk+cfUYLzBBIj616bU0xEjI51zhusFJIQN4EhmaqN
lIK1iJ/gSdO5wH042+RUQb7lIdCUqGW2AIOmP2Cc5A29urS7ohxPBrBzI22H483PCF2CEgDCQifa
j37ZPLFp0ac2dlyLYHVilWGSWPT+yEoH4nnfm5oG97G6mb5WhzXT9Xepp2As4FEEXhfnKyQiyig6
T3I4WBhQMZavnb7hmolC3kF4dJLpucwM/yIsFWUkaY8Kh/sbEX0lq6/0cD5Ofmjd4T2TQE8NBg97
XDFpk4gxdQb3+4ZA0ZgbQ7nxZQM+/PKacstmRiAcBGvNseZvpVbHWo34io3sHyHWqWy0WRnPQ1YY
R0PC54sVBTiINlQtEjYL9if8CHmyNgBq8UwkSXs7zeKQylA8fkHMaLSqq2onR2EWPPoP53S6EMjw
RiUBMrJMghntUEwkhIhJE0yBYVHzLeQXKdhmPcUom+zBExxokTcJKfSNZMKOxLCvwSO9fBDPWVgi
PLzdPQ+KYkQ/5Lv3XYGQ9FncsI/nMMeEFUnBBRQO6xHmTWsx6FxFds7wEJEmtTbWMFvxZnEic1cG
RkPFQcYRgnr4CZSmPN6j41wvdaz4p8FTddj9tn4iKO2k1Ktp9ZVHfiW+eb9RbqvpF7dAsfJjFtQy
oZLM6GZS2QS4lweKOKkgQqjgav9kMhurTgkaGo8gkStVikc6G/1gApTbLAGNfxay7UtUSxCHbT4i
cnhHokVB2uETVBmdBEogvAMqXMxEaS/CCwATz1y1zkX4JScp0SEJ0UQovCXPrSjaOIeKF81JXJ2u
cHTlf3xMecMZ3Pn0dxFTaH9DfmyGkCp9kH0QWVM9WwoKU9ddPOGuNEUQpa0DJ7scA3wCl3BD4liY
sphj3ES1fQD80ylwQFI9HF9k6QzrI2iqvfhMS+TTHgkp5UiP2vF+6oqvgX4tO58DCyMz+caHlVKL
g6giU9PN594hGSIph146S4xOMETEgJEzlPmYkiPURG8Mg/R7j3OVHgTw7zd3k+P9IaVFjpAkxuMd
aUNsNBW4U3aL9R9amCljHNh5SJsSAW7aBv/WhYtX3wFFHeOCuorQLiPAqBcB8rrnzwYfeVOpQ4Zi
TiB0jj/mjFqdw7WEWZmRqYL/a7xN+UnerbnCYDloyMZaT4WqM1qgObDAlqcyC6xC1nTCzXE2lgaZ
PYbA+Jw1JE5Em46VJwfCtBRweyyiTXtQqSVlL6qquf6OcNIk4mauGMppYZGkqwXq2sTu2iIZs5bh
NqPOwtokMzGnEQPFmT51LTFNi5f7r6Emw+KWLIXClEL/3x5pzFh9XtAPw+2gpgNqiqWM+vKLzRuG
p7Hgz1pdWmGCn1C/Ffo6efYpXMbeaPnx7+wKiz8Il8qjSjUgGBhTRMFDb8o29PtUVSbyuJGnumeG
TMpVqZEu/og9YM0bDZ295f91wn0iLeJljMqEIv4epp8zrkDr4+bB3W5NH1VYsiXjnSAoBtg1fqUO
5YpGSBG+IjpAOkXEgBlgbuH7PhVpi7gKj1ys5A5mU5KdR+IlbQeS4vHT1nb7BOG7HysqJHwjMMNU
4TwSL2wCCCwwpIwJdyZdLuNwnMa/YLCGvGhAA/tM5NAKD4aeQAwmBOrXczMfZW++DzoZPtSRW/FP
RLZAwz7gMDHitCRKsxGl+Ba7zdMzOpbbdiaL6vYKwckD8JLRYsUJUnJq+UrOdHz3rBCOtSPPXZxR
6HEQOwSg+7FzJf2BTH8S8e9uAUmNqnttcRUDujgmGtxV+U16j4/xnOYn/y5bbL1fTvGjmZzl/peH
ywc2L9GINVVQ40awIb6H/6q77gQRrbxBFt5wPBiBj1ZFT9OhvPRXNFeGsxq451s3OiGk9kzTZ5hW
s5UrETtLFP29IVhCr1YmSejkrhy6eQLMYwY4Il1t8lI6nsRv9woYdowfcSJJxo9bdvuDJ3p7u/xX
8GKOT4w8ku4w68ymqv5zJ0GXHoAIMY6gr6BRK/ZGU5ioU0GKhO85y1U+74ajsUT0/G1LEmBGAYk0
BY0eoSxfv/Y8eSKuLHsxa+clPDoGYJGehhLHRsFVzEb63rjkBafz9Fj5ZrPGs8O3BokbjlCjnkD3
wQDwLPnKJaRSOeIavsdEbeFNXfZzpfrbgdzV+OeJPSaEQ5ufyOGYu/UK1lwZ7NOm8D8T1tsNiFBd
Z6YMAOzdrpg7YjvVwECkmPW8CdX2UbZFb+H4UhPeow81GKII0+OUSoV33YNpg0qyVlaxDx9QqwM1
hMGK8F7uRsvG9fzpKpoNBPMjz5gm2GP0OryDnf5WjAbQcLqCW1wmiSOe7jtcsL76TKmhR1EYdQe7
QVie+JU2pKWTgS6AmWAcWMg0/eKDWyjGTnovMAiGKPVk4ZCbuzrBgpLyMDC6bMFlURBCQOdYSIwl
jiXtarMhhdgaZz1YEvTtZ8mAJcb1h753A1gC3xEuMlSQj3QpRdpp+7G20aYV2ZSUXOlC30IsAvVA
0Xq0szr08WBUvas/Q+wSHuxdtCZ7mS9yCO7aF8Wc2JY5OcSthpBD+B92szdUYgw7SDeuLEKJHAdz
4inEjZHJGhKLxcJoaz6ZWPaEQ2A8Dhn8pDj73THdtfsekVLGsyoWWHgxs6gTs7K/08AxjKGQHzqo
P3jZplMF/al0gU0FRkG0yvJ6a7iV1SR1suwptZTQ/0GNXrIBja8A0zZ94bFnGpIqeSHBaOfQJC97
FkRyTsNn2+Wo4kcB4/7bSwDKWFzY2c/uvVl0UHRnjRx5Sn/mCbgT1ebUD71ZArE/ARV3DC3KfQy2
NTHq92HdnmG3PueMw7tQNVmsY3vKtgKKkQgnyrEqzsaBm2k7ikJwfiLIYMf4OAFTig+DBNeLm4RQ
wbLQCgbllteaPaxCx1usINKdI9AhKdPW9V8BZ8TkDaNbPLnUOASvQx//wDm44JbNdkRoURjlKwc3
xZVnR0c+BR/lpQFdsGHEAAeSGizvxfIlC+FzL0wtwa1fHx+gQy7jMXpoefx7YLtFIWJDXq+h/Ss5
Fsqf7uDe+HlHumpORZLlP95Q1F0j5CBPyXsUTA3sN15yXJdFZWi89isnbKXwTHu0P5dDS8+WqmO3
jQicRa69mVcmHO1ClhCKaCtGODmxKLuRnALFjDLj4wSBERLbD9yXG6uQJZgnBIp3wiVL2xuD3C3y
TVn5HaKQ+AUajgZb12IMkAxvJvrtCfwvz6aC4WtFQfLccHNqzqAyx1oA6Gq//eyYtpWe+ga4zi8m
FlAkAiKAnaKRaNYExkUPoTrCctVyL77Vjfap5KzcEfP2frLmSLKs6NBYXwOaa1zpcLees8i5eNfq
YAXyFB+G9tD4PQNXhyAFNhF9AZ+9kbQuEdHYKmZTT7Oqfsx3Cvj5L+5Vfoum1JVvClri90qyPvqH
JdFxYuCwrbhjfZPydlT46vSTXsVcnvm9RDRY53QmbvUpPdajc0hJhu3QO16SbhH+FvOaA6cYtXHz
UM/wA3bJw0oVKqhXv2T1NERCWPGIMXmETwM0zOl1+kg458CmtwwHDiROPIkQwGtNgRJG3qUV5bxE
ME5LWKCxWxj6Ch0eZZLeuQbSveO5ZembCNqIthaaDK7UdxF3Hhi4tLoDQ6i53mFnl+k4hguURfoF
g502giCoHAfIYCrAWEbx4dxcA/2I32nkyMjD43n/Re89Qbm7rpjTM8SIwdywY0ZSHufGhBhtQPGe
AGUPSkP0y/RGEJC6xf2wACfvVxYg07XexgdmN+8Kf/Zng1hm1mJu5VbPuMDwBWi7kaHzQLC+Fhid
ygCKV+DacLMhqSYhxkZ3X4JMSvpUmaDzKE4LA9JmD3C4dqyCBqicyWhSPtv/6q67K/0yvz0GXT23
+BK8eMjMFYDhDMZ8szCU70CodhwZX+Motx2uaH0OJc+iGb54f1fgmkhjDi/6SIltsVZDZMsFbsFH
P918T+Dvem5xDu0pa7GGF1uSUFp/C8ddd2U8+yKJeErGVdZOF4dRWrQi8EgN0UgGEmjYg1HCUaD2
K4DtOvOQUhS7vwX7+kCJOAPRKhWITbc63OGcjfTLDcptY6txjivrVZW5zfVqEKtEn+OdeztMbhRH
9TIpCjsgOF6LSWe5Eb+us4jcWG/ZD4KXi7lUvbFzboW5xGpGeqbJ8cLyAXon2ZfhjaSH2rvycojt
6QWtsdogfHj85x80ptTro8UAFibOXZoQNVsTcw5xmpXF1NLk3Cvbhwr2348QgYKn8BlrqLp1ZMC8
fnnYJvC7bCgCyrt4H/QkZaI3DP3rEcVCxL8t0ETyN5ftO+vnKUoPLC4C5SHiBQNQW0ih2ZmOnLig
QWPLhgWeLKGPZPbQPn4hhg9GPyXgDqwizt7JbPz3IHwsWZdABc7vFo36wBX3b0C25yYdVeUsgf2o
B0km1r4h42s9MIFuCIVXosOhktowVYlIg3LrTJWw2wvLv+dY4bKrrKKI3yiWjjhEr0c0mfmceb1r
eBxjk2UaX6ZqnXGB4dsRS96P5oelzRrvs6pYohV4mZnzzFFEGyT8BTUKL+SBWTClTdvMrdhT7OPR
uqxusym9VQkofgi8npKSoR+qS61fR3teBtRhh4x3hq2csk/tdVi01KefvtB2D7AvJvH51M7qXfXW
H2YyGkxpfTV7BgU5VFX481mb7M4VsFdjyRU7c3vTJ1hyRILziFlA+/TNguQSj8DOXUe99PY+1HYc
17u+CuPKHrnCHe1HYGEh4wawzzEo2WGeF3ati1TyXbWIeNegWFORWnpAJAZbo+RyGXUfs+JJnUDv
4NYJrhh0o+vNcCW0Sou3uXnCnS52Ffxwy9ZxbC+XYErS6+RuuKDc9kwibeO0UT4ul4Vw/KfuK6He
7LWT9jMCZn26tqer8BsNkdmlCuPZ1B4D76lS9impoH6SV6UEusNONELAVHnXxRFPZo/SCEnRbyT2
GVy3mqcrIv8c1ccjdkxlmY3h6dcE8P0sxt+IQS5YREtpi5rFp7iIc/WJoj2A8Xgg5pqP//gBGLUX
KQgbhTp0VjG83i+5RN//+ZiyJvVcQnjxdwiJ+JArHtW8b6zIbM8LJYEY8IZwoWP6dj9C16QWxuIk
m+HrMr2t9+CBPJjHoFm5w2paVK4qXWeWfldLbNIknfo0U+oD1MPwNUqoS359O1mSE2qufHwWPoKZ
GD3L+MzIpZDljRiDzwYqgkGubWMNWRuDrRtOOr/WHnwL0iWzY4r4OWENZB9xtMTMijSqNch4D80+
xSrfJIpJ0+mPgoeBVavi/gfdVIUMVyDfH04IuyEFy169Stfv5rMeQJJBWQydDl/n+nr1PhfxFWbV
XkVdfB6g75+eMPKshMY/ETPz3PaF9xEtlK+YoK2jIiS+lg6OHy7r6B1rL60sUfsl7/IA6tbzibgd
IVLJnZDzcRRwJADAWlndyWklJ3zlLL+eVylVYZcdRWXFBZQOCbuo3Jf6fvAvR8F0pPPhpLfP/zj6
EOrIDce5RKbSUXcyxvbGmqWeXQKfm1hDSKIamkPrhTYWbPQcUdkXA0EwHpfOfkQr5+piJAViDchh
i1hzMaqxgRH9f/4cIzQYleYItnfVcrybFqO1qYIDbtfP8/dSJG2eX5FxEHcOzjH78qe8pwfkFVSX
rfmSbJLb6e+gw30QoCNeGzm6DmHJAZ6P7Wp3oobZ7b7IM7BknV2eVVil4rAqc2lGmrQuO+gM1FKV
hAKW82JCnk/nH5Ljl61TA2ErdpCWv9/yOma2jIChLXufySAnUv6QYpBdL3ObUXCPOzOo8zN0F6UZ
dRd7BS8La1safn7DKn37SKHKc9Uf35ALumAQok2Ncah/aB1kADEQn4PxVrDwWBTCE0M/4Rgb81iO
mDLTVG+xqMk4zYaKz6PpjaZc9ThKeCarbaIZqggFwaZLYT4igKcj2MOgvvQgehGEQO4JlNOLyNDR
3nbAJZsE0bsSh08R+2QIqJw8xLJzS7csEru2xHZ2HyqT20mGxlgG2smn7tAeluSVthMUZOREI+Em
bhRKB0cBK7j+UzZS0CpNG4rtKZYOtrFyYupUQDY1bGn7KuJ48J0tqOCDn4eNabTF6BxFWgM1ATIr
0J/EX0X17Y0JF7xu4GlgaQvD2GupoaF+FuP7OueJVyrdA5oUSqKVbeBrm/RlqgRoTuhkFokqF6Ap
hrw2EjN4Hx77fXQBxpJ6rbYQJNIpkSooh4yDImlUJhnj+r0+aJLpCLbPn8gnkiPLhtbGlLXzi44s
160YlXZbsCUcVSekflSclqYITOUR/BmNPTvB08Lzxt7RHpxZcBkvRMZHjhxjEVzPuilbhx6SPDnm
tPGwMBc0gUcTn1/zwm64z732gE3AFy/L1T7yp+r61yn04dWt7f35Y5THKZo/Fw3z759ezy+kbkR6
tMszc5HCafVwk+Oe1eH4XTEC7N7S6SI3JOBT76G7PYY/ttiNOdT37cSrfDO5cyIFlronBqzzChjg
G1OL2FRWIIQUnW+ZYP5yzdTyV90J4lD/eb4q+8A8H6hDma2rRuNpqe9onyZphd8Ka995xbxKqHuh
+gQXq45HncrfPMh5/25jEsNZkW6uRFrIsqfGxNAzhSDYswpmZ3IZ8WwnETRlIDQeNsjFnaO23k+I
o6XNqVt+WqpfOn/dwuN3oxDlhp+s3QH88DDvmkky8lrrOd1kEZFuE04JKGLhEJTxdlqZ5dXejyEP
b/HQHgVMs1PuqlFMLNtcJQTXNzxItNopIVK+gTlKqSTNo8YEgDoE5bH6KpORvUo7jaYdYMUsCWJV
w80Z414hknxlNAMcg7TX96VGfALkrYecDX1gXL6uhZd3JKK7KZs/a3O9pdor9NT7ymCG9ASjeDS3
ZKrDPloGX3sarBNyGVO3wH0hAcNZQFG3LzumsyzWWw8MlJFj+tCPdBh0QLtooxD483Qrb4Hoom9m
3RRDdBq08z1QEPR2PHmqz9bDfi56bEwyt79UOo5lKuURgLJdtEt/gwssNAXwY00mDKXeOVeNMpSh
IGzQTC/cS/nvWJBF9fAAQYZ4tRV5rxCAHAeqSxEyXbyBO7/Taru37iL/EB+co6FPw1UXKBGovflh
Yx1gS23JQPgiHxyZyGZL5H1ZUlYFaiTj7tuf1lV+6TkVAj5Rqu7pXHclNXWZtrOLu8egR8cQFqt/
HQDf2jAEsvh9CTfT+BTwz2eE9cw4vmzJVwbJ5XivoVONQtiySHFjyhd9CJGWJ+okoW5vxP0FVF7k
YZlE7W3ofmAODZ0IDfatg9TB9yMl++6NtnIt5Ucjxh/Mh+UwvhwK9YpUiQ1w5E1TqZYvqeCjci/V
Sy29AGG62GA9k1USAFxTLc587Cr8gqIlLaZpJ9EsfuQgGI6W4UGjRp7gLgnstV93LejHxnZsEYao
tZn47qksw+mLjJiy8/CrGbtkPuY+ZYuWOXzWraOVzzN6MzPiNZ88LloFPjzBKv575O4ACcAfPips
ZVpfODggQj8VQpv6zkCuaRa6f/2xqv8SLuv5gUxXidNMTYAiNcoHws31yBTYOhRI2+FHvCkwCeBf
DoBzAzSwY7yMs3Qqj32CT+pCqmH28ofqyHsHkn61W0FEaeR+HHEFQFNTEDmd72l2c0QU4hmIj6XH
HEA9EDrJltr/ClhpihnVh4EARsy3HTEhJD449N4AeEDx1YG6tg5wzMzG2otg+NM57N1GNIGb9jxR
aWA7twSxjoA2weKkokcdzlwDGHzDy4yDxakCSR84RPTTnZer3Ax9IKkpl17Ggkw/9p3u7uikt85t
0KS5A+ZFieFkjYOhltofiQIgrpfSzBYmgAdDCUaXLJ+dlu+6Iiiv/7468aJJ6r0R4WD0o9U/p987
Prlq0m7fDLjB8DYIm4I3kkW4x3NmaOcuLh62cU7OZT62jO9ckQrN3fSFLUUGG5Y6W6USz2vjFllh
TUmJs012uEsFbn+4XzqyTje9C72aygF032qACXy3eDp1Jobmz2onubSS8q2aMJMRTz94ullISZ6L
ydCf0To/DEjtgi5Q0lv00PtFigP7+UDEjbnToqOWZoKJtjSEq6Q1yKVgcemAtuvJXIVSg3feAJel
BhuZx+SzCgTszqhgI1rS6j9EAK0Q6RlKNQMe6VBXNeX0vdhh5FUfBEHH/iGF+KiNoqes8NdMHI3u
W7zVAXk7wpSZZ7wHiFPFBP2eJUkvE5JOACI6wEYjiwTbQuHrSVKFTpt+cf4rSOlJj/6Z5JljHg6J
4Fi5eoCslTY5hH5/ag28/YlC16io7iZb1NWpwoWK/kvUbwV9/9e8FtgCqlc4gVnry5/AUVbJiO19
AZ7Jpixr/Yy9PZZryA7BPFbVbh5RdHIZ2Rjz+/fX9M8fNmn2lY2Zg9U4XOGRzDoeYYbydXXUzIhl
comzegATL0mSOum+zBQrHDSdS0TEGrj10n54DeywqRqsxhsnXaatbFwFNE5LRlrUjo/2SdXhXK12
zfRSlb3J3Fd/NquDZ0fTD9l3kyiUuKr0/CaF+xemK5Y4FdYWbnfBSzl2SkFBNB7ZwmGCNnvwZbDu
iHain5QLfA8xsjRx8xxy3r1UpxGbn6DoIlWh3P6QC+Sb/1TrxF0tVMkbw58veSA1DxU7dNFE4rRd
OIcvaaziylmPWBt+ovKQRMktevIj+sZ6YInR3JSrCHauuB3G2SXQZ2mnKhwPE0szDC0YFoE5DTLC
eGpIY69aX8wGe4Q5HkZ8acplLXRL1G77h4XwbZ3CeRb8HkKrfH/RJfv32A3Yl3WY6ox5QKBrywhf
Wre/ItzeaijK3koYnrsQAr5D5tBIQNvI4kMkHK+dGgvAQ0D/ORV2UNpgyNaO2trEI4evLQeHp7A9
Bicmp43vQhKdH2mbOdj+QjI7xBjbtl5f1q3QhW1idbmJRWTFDeuBC3NrnC0N5PcGsr8RFXnbax4n
Ri11YxcbAzIceB4DqSP7qp48Ez2TpFh9YSyvT+hhfeqNfCEZZ+dewWcnJOg8zdVEv0UzECJGeTbW
8dDZ4b7Dooa3FliEJcdCwSkmlLWCpmStDKSgc9rp+zIDZ2gnVCYvi4T3cPVzrDIEPi0Cz0ERCiB9
VFU77abcS095UB0HFv+pQvzCqOxcvSdbknbgWgtkFIouKSbJbzXa6l1XyJLFRAvg0ON5VwCTedoa
921I3kGYyJ+iJaLmO69qaMk77tdesyhoGSiTytsBK9gVE+YgW/AemCRyohsY8g2qKZLIiw+FdLcw
cpxvn3RafrukWRlHqyLSlrxQ7k478DQxjPJJfT1O4BkDjc0QO0GDPMAIgVI68JMVOhwJrEovWDDA
kg3k2ym5Bq6Sbnke0FHWTo40zw97F6qltw7oLQbwoIvZDfTGJww9JTXAIhXv4i8VCfp5AipW6jps
eylw9uBiRKJ5gyr3py7GusbkvkXj+ZvxcsWG01kYhEQ6gxYWH/lTdTaKaU8O5q+YziuTW3SXGVD/
iWoG+ImrB/JXy+2EmcV8Lqpq81uzjaY1Fa/t9mHp85ufV6iXfC/UfZ8/U4PEPLoL7IgZDbxhKQJ3
ObdTNdFyRPOYe46I7FU5EECcJBbNhWJNuMrcTC5T/hsSGK3UewBRsz+Ns0LlaBBISB+zR3Nk02dX
s40MrZc77Mw/yisf85koi/U0QXXkgfv9eacTLDBnA75uNSkb7xdKpy/SLSA6ITejYr2HpMjhI2jW
SbPatrVFF/xi3NHifuRyGN2mnQBOQGZ2WOXvBxaAvM5Dk/8TR30wFzdNehKwZ3zcCgTMCeKDETdE
z8sqSTBVTkeXVr6ahPGSemmHwKxAf4FdLX6OCn4+3bRduGHXK3cyTXXBTiTiF+WeBEa/PQTdEMzt
McQAE6WeJ1F86RxPyNO58HNdhInYY2gQ7gITdubByLWYQTXrZEjlbvqjHcTHqkBPHBAGIInt5lHI
ihG+B3v+JAYpRomMkH5yiCFVM1Sed6rm+1ut+I8QfM59b4TvJnAWJaA3QJYA3J8KBinpRlx2TRGG
rzMjb+ESobh6jpwL/RjJkkYtNi3sRG+rGqRSmRQ4cyVXM1gCqpXOwck3tUWK8/CQcyiWyIxYNwK6
Vt8gn7b5lJ8wqWEjLqVVU0XSaCKkQpd+b+c93K5IYPlbnlttL3QXavniay1ip+z4slUTwZ3qYLpT
90mx/pbBmrTyV2AcEtUNVxw8y36KgJSiV0ik3JRmWbPPaUPY2qkP28DiDSJzlY0q8+F0ebFQBf+4
EuUdIKCPUDV4IPLQ1vlZ8E9EMzuPHCugol/ylHhp/rZk98lcyyCI5jZYcEUAqFc7CPStZko8SyfB
6UoCKE75xjy5EuLYli7f+x8ZaRhaboDcQjyf+BPbsA0B/mfgvb6asX+gCKptPYVceW5S/x7KlPZK
TXizhPp5gCrip1wbaXF4AgNx8qyMkaJuvGG0NW4VVJaOLU+JAz6m24dxD0j1qOgsxpwRUYcXh6cm
BAzkNpz4lynikYEpvLct3bX7Nh4qwjsQ42UmJ1o8lbfDbIl79qazOGWMbOZUE7dadZsawd05gfnE
bYf7KEduRHwthJBydk4dGZBHd5oyQ6+gG2DwtkyEZQJctjDyxVPX1XVZ8kpaOF10ujbhEnHNa3yd
G+BGA624TMSbuV7TNXix08CxVNZK9tawrj8Urnm75So+cOim5xCHM0soG4qEKrzqOJp1YD5ZdySD
9Fks2YWZbWPJVztQV6vIO+8t9Zp9iIbLOmo9dwnxpuiCiSzaLyMmrR8OdRP4P3YIS+6kmT5RTtGM
1AiuNWZ0IShEJHt+gpfWTxlIYq0ScmWFT2Grnamy6CmrW1J5ekdjIOq3vM/A8HXSuoWx0MxJYLn6
xqnadDiXssIcRV5P3sWs4/WD/JQAXxA7dvNKYcOHufEqc5H7CZhxE7H11jEK87LmrMTUEXM+ptqw
3xRDQlmEIYbEvG6WQHz7c3jwp/nzeA6TqhDebARv3IKJgKjuNvRjuLDZkxu2wHNv1G5mh/HMJ67k
AeGYdvfLb9ZxV6q+hJEl6VHvAf/RVXQt53JLs98AkH53OCgFKFxG7PbhQZ38qnrpVbY32/Hs8kQt
TAC/93qJrv1/yiWKaaDJh4m9cOHXSA69W1C2F754aQtEEETmkHBMebTcVtPsv2qcB4h0XGBfPXXj
504My9dlJRwqq/yk7vXkSsgIcYgOWApgcz/ISkiaqpoKAQjbXOBYoewP/HlLGC7D4QIo9FAFZUXP
6DDiKXcqHKSKjhjpiqZ/46ASkRhrVpO+uIJOP/QC7lNm7V7XlyJiKVJCh+KGQQ9KELFSysUfKRgL
GSHIuXcCFvibOgqz4DLQso20yXQgd91LfW9y7giYjBEnYf3zpx7Jz/thj2jA7XRmDj5fi0U9yi/V
DqIX0v8sZV4w8zMwytnmnVDSZ/kd/hLKD00J6rPyU14Kj4XjAmyXkKSWQ5ef+Kz7HPLShQqzXzTi
sE28+MC8IiS+a8AJ4oFQJzs+BuLFW4ptAzfz8fbnl593ynnfn/cfrohousHNHa+zIkOfG9dALwDU
T69oyXhZm+U7s/ShRfnvR0UVY8KgD0YrLlztl8pdSbaqHQJlOtF7d8aOqAALvUyP2dFkA7WXQJan
WPP34R84fKrLYKOFQHRLBhSxHqNhCkWAAUZXDHYDBnyIQEoGrzkpp2WgSROIXJZNrbfpqqRr68HR
OloZNTPwvbRd8PTyV2umEVD66DUwkJ71sXOqZOL4FqJdnUqJoj73gDaCq4PoYIpopsMpp9BsZ2FH
cBZYVgm1x0+5PxXbV7mUvQFNwUoe7arbMfVYxRo+KzURsqxcZE5KA3PwtL84oq3iGOcniCs8shlR
zqaKhvpz0DRFT1nrHY0FoHo4/ohQO4E6Kn6VLqaSegBx3JmkfNWrPAuhDpg/sVvmWnHWn10F+DLW
3O1orv3FcjfZaT/osTRC0TnS9Smaxnx8MRkoFVP14y6WMPI+F9FTSrfH793F0AYF8sEOV7ajSAQf
J2LKTOQyp+LsLXwMrFD6HKqnvbPHVBGljsBIntpQQ2Kngt75OXmjVvtUvoneN1YI0EvuF9qf9zMM
LPwJrukq8I5sQ4s/4wECYWUNEfqtiLRxuQK7AhrwM2PmbeN1u0RPgm8v0Rzy1kgJNOKO5aJ07oNp
9MrkGx/wkNfkjwCC7QwDZZ/AFQFTCFCHBKXMJC/OZX5Pqx3fYr46dtX8UEkp1NxZHqnsdzj0Q9yJ
M7KxxpdP2efDojQuL7WErzDk7ay3bcxFIvon3G5ZQOE9ZyMY8yp17kudl5CtAodY2iukeaxxheN7
H29FrAQQ9XAROVV5hHgnCGZSkBeMU5mrTPt1JHhdiKEqKZoWlx4MZGChYGOZ9j9n+PuP0xxP9IPt
P0/xsCOjl8hVQlW/qt+evUWgin10jha38hpQ5noU2W2P1Zm6IPHzx49cf6+OcfPE/0wNAk2ZRKAv
jTx/jOwGwcc2iFm0n13G06OAy+V61I8CJK/Y9yAdytKLYHjPbuvHSYXdS/fR2UwDk86wFX4aUqXK
QYKjejWtURB1WjSZwi3aIB+xFXHYKmVJ9O0o4uzBkUzMAzQV5JnIPkJ7Sh2nv0ItoSXg3MkrCaKQ
cTCfv3dOMgRdpLomUUHfcw6vupH75Y3k5HmNhW2fFwtzFWHOzgeuC/J1BLyj7Jktfi9wdJ8h6zBP
NbH/Ov5PCsG9N8ATy7XlY4qiGUXhMnkwXjv+xfYxeBt05MQvOeupy8lRs0S46Lxx3IhV1LPul/Xc
vklgJuGnqeS7cipJDjrzKCnl0+EvLNJY8AH2lQARw1xmxGCUKKMkKNH0dVLlUHA7eaH+QLj914zX
jYuCsxTorJWLWBKH15PH1i52OPrdXu2sCdEZIrlynO18Gm4c23VPhq3skCkvi3lEVsEqoezp69om
04huDQ+kszjpkNbHcH4/k8julng/Q7mUk0oBOeN2O5Dep0SbqK6HPcENj1tEVh5EFrHVRNcx3dl/
YtCbo7HVF+sBryoAqhwam7a/i4va2ynUxmEciub3Z11XOY85PVcngoN97tcKM/Mo3tMT8NbP6crj
zTz1/nuenXFF3AE4pl19XL9XjNssvlAflxit/DtayXvkWj1LwFd2UPOmvu6baMG4ByB7yJJLIfih
4Zz2o4tE7EXWJCU8mIoF54DyMW5+/WhOGxVUAviLwVn2wVXDCxPZliI+B1X1wsEnu5eTjJbg3OHM
kHdA/J0eapB8UbpQK9FT9OYITUe6P3EuNezJVbi5MR0nMi74CEYtaKaBsszdTdmIjuEHF1lt6oEO
Dui9v59tKvwn3vFd0DiN/ST5UAlJT87F/JYL09cJqJ901acVAXxcc3PYCA98qOBuCRWFUOp7R2Kc
2EQrdxh6l5t2gMNTW/ijlToVg9CCOFRjgq/cdLsRiZa4myz09eGPp7OINk9B8LTwNZ6si9ZCBxjC
5R3x46aiCFc/902oBmvkkJMSu3ZuPKgwDHxnIqgY7Q2rf65t+zQnXZV2PpwSFg0JU+Grrnr2hsjS
vhIubgxqOQUpbld3++sR3iEkDp1T53KM1vtsyz3yA48jst4Cl32zdQNemHUo6ibeJpPdbJd9ks9W
6Aji5Fk7BDNOeWW/olsB3eex/yHcGsjzwdWsRMqrU4iB8rKEG1j50kalzym3dd7cbGDRROYxFCa2
KjMaFpkx6xH8HD1iGdgSIkW/Lp7KZPn59tMA0JTEW5fwY0a5hWVHB9iIxIDu/4J7BKHjuqQ6p4mt
wDXy/Wi4lj9HrsiEBWzAROQQisiamtuGYjZ1KV7kjBlZa+D1gjxEA82gCbPL8xj1JZPTDx6yNZBm
CBVr1aD2Uco/AT+Dm+WCkVoKkTxJVOY3gcuHkZZuA90WMViSMKZdCQ3P/c2wgeyuAsXORHAqPizZ
xaP6pEFHYnf338XOYnabR+aMi1BiawV5e4P33vSjaLAgK1tBGqZABSpcYexbMHMox7D6hdBiToW8
pxC2UDzZ5F8njl0FVNeIdhox1ofkEBRKzzmSsyHdzG3pxzuSO+XzREEovffOUBNyd0P9i9l74vei
rEtvC9og7XfNdbSyVCx724T3/+X8T3XrycHPLh6DV8HhowO/I/WScQXVG8mcVnUy3RFHHoYKdMXe
HqJfw4pyrG5PI7xd2d+jDkxNuuPosz2BF90i/qbucSsmrT9Z7GGpl5GW35YhtdphTcAY7UbvvVAO
OcIXVAqTXz4g/Ce6IS5GlmxvpgXGbIf32/3tWxcLeuxDHHkKr03Y+ABHoBB4oOhj3cLTiDUHk0SU
STIx0amcAgRCBW2/9vi+4ZRLBHwmUb6ThqQURem7F+dl2xIJfAUYgvfdben/OJfrtOIQo0yC9Uvu
YkQ6I6xCH49rHlUWRMOLSGQDTH8bxqaVE3DrciFLQYyo9W8PG5TmcgcxZ860FoNO2fvAwc2loLAw
tUyLuL4+A5ONNwqOoiJuPqaQG4gAOJtJmlGZe3XOjEOpHfyOn8ofdYoKNMDFB5DwgtKHIyh5yZcy
s4E9v+V2syaKD8wSszZnPvUuHfUIbze3cBSSCZH/Bl9K5lwhbu2BCLVIsuQtMYfpDJ2+Qd23QlX3
Mu2C9C0g4Gb6/Et9K32a5DCbG/jXpXu/AqDiNemggIK3sz9t1yrzo36FOr7xSqufE8TvlxdygHdL
32OMRqN9p/XI/IOiSE0j6VBo0iWjivqryCVhbW5eAXDwrEvUzr1X64K2HVORPPNtbfPQlyJDG1L3
yZ/dXRD46FN9a6+psgTzLSF16uzP/XHTWYxtziYCSBv2o56h//DBoNvOUsJXCT3Bh7Z9LzOhyfRD
HlrG35Mx01uiEJHokKs09+zlhoHFuLlUwdUkMn1Wf64NxypFz+IgWPgtrQlJywkZ3Yna8+YJLuwD
tiHvX4X2S5kKKWPvKYu1Peb5zWcHAARfxWLRtl0Y204vG/fcNX7dybzqnxvhhGm5AraRHydnRUIJ
deWJeUGMEbY97VAkJML9HL5C0RowIRdW7ZjM9EHEaicmOxwTyLXvzqNQ6mDAZXvXMTI9aLPH8iTl
PmhXhsGjrSiErt5lOGXGSacYcQzMjXTpDwIY/+IL9UIlibImaEzXXQqHOKk8GkWA2m1bb9u/+Usv
1kebjI0TlweHD5TzlGXb9G0WC+WgEHu7AfdAfwM0VSTqj6LwZX9YfpKIRXQBQK16uw+523hkNly3
jYIyjMJ0uUa64HWv1kgBXHj1SVIoUROEDycNluA5SLU6QDXqH2WIz2DWsHh2jHfwgbQz7B1JkMNr
7rrBfXJ6x12LD7JaR+wBfpWEC2b0P/3q1mIuxZ7vG0tonuT8lbTITe7J1M1teB5htvPTAjQWMbQV
rSnBtJeqAEUv54nfP19KEThBxq1H7owKHXCZAsu1dVI2WlgsDO8giuP6g7Yi+/iT1ZWv331430SX
64wqzxJEutrfoNYtlBXwcTUvv0VMsi+E66SXptBShfRyK8pWnZVfKLk8PPmS92g7CIAJMOpNfqwR
Frn3BDloCsDAzEiiuLf64YsQ5W12ITZWfjGoPVavoE5aj86qVjt202qrP6Hlzi3xN+uLoPCWY2kq
cY8CTcwmiEMlWYqKPyvIwGElGa2EM1CLh8yHzZds49dTXZnrmWPXANPSOLJ1WUbKAmm/Z19y4HDe
J5iLSnUPbqK3ywDB+vZSi1rdxGMmgdjiYp/OmOGpQGEe9yOhc1wYbLvX3qccZZyH+VdzwBvF5r4K
va2Qiksq5DZyDfFQEfkKr2kHD+eJVTnWb5uPRU8+CzRr3wQ67RDtSC+mrvjltDbgKK7CQWhg/uzI
+e+zaSODDsOwgANSrMYsBg9bYqcCG0F1tpeip8n77Yprbcr9n5Ga5TyUZlOeCn1+V7upPKo/CdDo
332rqVpYOhpmYOTZA01AOvdMByTy3IpCJTW6sJ1PHCrRnTIQxwvoXZ4jdREmohXpn8jfOWxz+BYB
2Qbpwd6M9mU3jq3J2DRjDg+Vgf5SJUAkQnVyTqmygeY+d8UpHdY89BdVA7TOuxgVwE1PXz3nb7SE
yVR7oPATXIBPNHRtdegCmCZ6h+NxlsdurDP8yW2/ahwllW8pmgbI9QwzvYCiw/hLUWHZIr4K6SmC
WJ9l+7k2lEmcBRrhIH5SYI5q/enHQLVXG1T/oOjjaZSwuOCInnxrTl6cnB3eG+dU0TrY0mcMWvRQ
p9onBoISiT9stUKTifeLxLO8WN6iWcUxvVtrY/wR9kHMOTdxlY17ZOlofY5D4fCXr/17zAc4M5kL
ixRx0RC6pYxEnQ8ldYSTEOkcfjcq/gCKshMm/FotQF6rkq0r7lxuKe7rVfoEfnGEqS1rG64VLlLd
6DAW91qB2DAW3ZlcVwHrz7c4+rS03NzZ4l6I/8EQLZx+mQxof49OEMu6B+B/1Vj5HDGHEes3Amlm
cz9HY6ea1NL70InEAzalHVIUYp+AFWk3Iw+WxuAYZWSdicwapxnKSbSvymKDAsLRXt6MgFGG/Qfr
T6eOZMVxv7p9Q75qEQ+RQ66R3/+zk+SDFMd+ld9+t3Di6iDQqxhafP1j8d92ya5bXanykrqRaSp3
XFPphCXWN03y4pm+jfODm1fqBwwtMcSmJw0irBJQ37DKg+yBLZ9LGzZ3tRFxEPRdMzrQOiQbfKLj
+48JXEjXwhIcOIsBiL6xPYoql4XS25UQA57cefvssPUgf3QwYPi6V9PdOjQ6FBCKL2SElm8FQ3Np
1EF1eOxb0xsNLDr9layK16a4afIcFcCWdl47OU/SQQYwQXH7/4Ik+i0oLvNV2i3fa9MpSJI1+YPg
RYpjCZll3nLJ9siGC2uaqWMhVFJzVYTNJjzd+NdxGxrT/9IW1iq0aTIcmm7L9kovb/SgUQQSRt6i
submXQkddIcWfntiN0h7jVNsXqRFqNOXPC4PuM3y/rgfiudb7QYdBaRdO49kwQY24ipjeb89YYP9
CJJ+5Zq7ykD1T1dnDu3L7KwH+B46FRCsquGlqDWohUC7o23yCHyB/URZLnQrCQsxHWJinEZU0zvi
ePGMfZbGAUNNFMDcsQ3nCJRnzZegcxvbOtIrE8/F+S60BMJsG3gle0SIFA4m4RTWAjWdLwziSbEj
Z2+HUTLsG7+LCZFGov/zDskd+6K+eEnV+Sca2feY+1EVQBsNNdKYnyBcpz0UeMQrdrGV+njF3iU6
qQnp541IFUV3w/8Ef7kVgfUgYP+weHSji5T3sjOcw2hSMUy/B7UCPGlLauUuTyi8hTaz1aexKuAE
CPnpkgYveBu4PbO71NbroveaydggCU2BSb2qaaIrawPBthvKm6wPbJF67Byopm50DWUvz2Pw9F8v
/2bVgXis+0rZTBVjse3drpX5vipuEPaFdVjTU+h00tRdaBUzT/N/QInO+pfk1k8laS3DvYU8cMpL
VKvXDoAoTh3l0+iadpf+h2iKYS6jAnSeLPJg22PbVMHfkXNcj10aWCNja0HXU77ALiV8ftTTI9Ka
+Fg4gmN2D4ccGqtyZ7N92IE8eLJDWgiPDNUKrwPfkT1JYYH902E204GoA/gpau5HjWoJ2XP9RSD2
yVVsk5r8ePFEHG75jvfas32jYwsWISTZ3SBFESkVIeE57aZESQXeMhEoAv0VK+JBvZSidKJHkDTk
wWfa1dR0kiZyvgcjykp1zKEjqVNkM9pxGVk3CrO7pIOXj25Wpkh5XOqv6YPbNYED5ntxKC/pjNzr
QKiVN2TkTHuESp+kiXF8biiS8NiuaoL9Gn57D3G6VfWXepyFHU9r+ZxD9CFoAOvbLIINZ/dHIIj3
Xe3Mjjrs9FenQqibNSn54GcfKlFV+rhdWz7qltMnHaBu34NijYYarj5j/o2SOZAvBtIYLNgqlYXm
CyHi3lAo+bACD49Yr5Z+1WtgLuHI2KVo0oWNfw0+2nZ+3VoZUGORsP2GkT5cobn6HmqW0uTOwBNN
zDRjNgwPql6LhL/MiKmKrF61H3PheqPbgsfq4ZfgclW19IsNz5EyZ2IH8MoTz8vw/QoLR7/IOtzq
PmR7a59AxFEL6o/HWiKYNRdrmFWF1vRH8Hwfq0WXVYJzX5F+rr7kUniKOIctyB0zypWAJdPdIcJC
E7TiRfKcY+z/ed77HMzzQDht5LqTzSgYv/gYjMg5k74K7BIXH1VaBamPiRBiZltlvCX3WiGeACvk
0YhIGkMEpRnbj/9zmF4CoVXV3Ya26fJIyLhwQOB1Q7jVGBECcdxGp6cPrjDA+4eukncPotCEy4nC
Y26X4bLtRoD79NxoxWhVYSE/6PgEx6m1F6vM301w6OGFywtmcD3cCEiFF+mdkAV4hH1R84fY1BNE
p61XJBcWfS0ZVZPTcd3Va2uJJGXe9bm7s8hTk7zkGsSTFUXb0NN7UoebLOAc0Y26JdH1zU38V7O+
Zilm3TSnJ8+oa7kJdA0A420mxCOMz17DBru8fw7Vv8sOLpidQOzcL8eg9s+FA3jd/wPZdEhfTRpr
/tJnXDvUhV46wiMuJMxN1B8VdA+tnaj6fuy+19qdSzY+yU+GyMKsvJck3kj2J/tGPKByPkl/xRkH
ZN6SJQz0kp6v6mY8R+T6WARGob3RFGfBbaqQ9TjpZrbQfE2ILrzJt/TNAJ2bwHHNbT0Uhg6FHhIG
R531vkIBs3IOThH86HX/nrAIl0K/WhpOyxObU3ugHxrmDJA0q3+yAIiOZ2d58zgAr7vbVVOX6dEx
qkrzRmT+9roCgQlrO1YCoESvgzgilaYgVhSur++Gfxi8P+LroGSBSjny9jGGowsRKnxeJJvoZEc/
N3nJzWfK7Uq2wFBFEii7+TcNMLTXI9S3vOarLIwsXFjPQJCTP0NG2oXYZ2s39iWUIx6GDcXbkSjD
/gakbA6No9oXfiuUlD2dBSTLBk9Ys7g4hlIEr/1uZRe+hxwZnaRfqdvG1j/QSxx5cQSl4GK2OHEC
c/YKA8f97rnq4r+iVqNdKw552jexRgVRRizduMKm/kqhRxUcYGxiTnbMmaWNA5KRQWiluCCLtRGZ
LHmiKU/3oNRd3CU7qpTQTb94nuZq3CE6JxdXP3PT2VlMf7ZFzWWfdHi3PJSJSuh85cGxhqwYLSMs
4EM3uqnpgRNgCUnqnR+fpdI9jV17Waym+gF0dLREDGXsaJhsNQXToG0+GERBj9PaJrFUJ0rq3U6E
2zyg2Fz+wvzM9aHMeEZSk8X+yxHXBmdP9PG5GhiU5bkLIYRMG/1qGIPDO30pvrQomyBNCqgmSBSe
hqoWuaSv1nxQDlLEHmg8L/XUpdBCjwrmjJpjfXpmzuY0AI67FhrEOi2bAtkQcAdXE4zrvmRkFuEb
ZyT6wl+eIn+YSCr/mnHaqH90cuajdc/UbP1l6AKaEZpz5nnx3Yo05qFlaBCODHb8nKqHybhcRU9H
8Mf8gXeOg9Nv2mJqz1xuEUj0sd8oVL4Hi6OPEcptcatPNYoQ/RTqL8Zs83uRhsUGvUqxuUdE+q37
LJo1SAVr9YrP0aOUY5HqicUexra5tRmPizY8utOBn69baxzJ23Hi7K/zemYvy/U5TdeFtTpYUfN4
dw4Dk943kSgmvxYT5ZLu1uIYIZAuNdU2J08i0uZJi3fudP5E1XdvocMWfdEFAZHEptRdpfaSjhr3
8fZCNwY9YXznZGTb2/V9bOZpp57Bqadd6NWZ44FZSsK+IAbDU0sb1J0zDL5SawvwSifiDc8z+/Jn
H7KcsBVre7aXZPLRkHl8uCPttz5vPp5EwyvijqDWKHqSvVGyi60Po0vNdaeeQRk7TWK2pCe/4Jsp
QaT3fTCr3cq75vP2zlgffBQ6SnxNbeZckQWprnKK3gOneOpUAG+lT0SsMSUUcU+d52NYaciBVyP+
TKkS0bgS5E9cfQvx+aOi6+Lr9BbsWf5nyG7rup3RiUwscB86pzkppmYgu/AMVXfbbAs1tq/SnWZ7
9iczilIcv/Eh/s+gISkWyXSjmk2qSY4HynBK3sjZhltSjdjj02pzj8JyWY246qcC4lTJBtZ41F6O
u+bdoLTytwlt60OLeXHj52MqLH7/Q97Tff7cfsUeTNzpxhwldGZ4daksm5lQYXMCmAYQ8il/iZ4O
OjG6DO2K+wByTdC+HW6EgYzW39PW9Aq3TzOgwF4GUCPVMO2OULXK7OEhfzKCQL7f/Fao3abnk7/P
n8RJ3kAV2iPPJNqqkEReCRQXdGTaarRB1l+pBbLU9CXT475ZGf1PORR1Ljfa8bNx3UpJi+OQyfIu
HZwNpEu/MHs4OGeWjHIZDkyA6g/yl9UeQLwVcYe2cBqB2uKbWVQyoq7BjZSIhRf1jN9LgV2ZYpDs
RBonh+ke2n1ZsG5+RxIiyoPEBYWsDmIhGqbAbpIIDYfVcPM9dKd8hJG7aZu2v7ozk/59lCVuw0Ov
O3mFuKoQbCTcUh227JEiCY9d8/alvOQajr5AfNQWPy1ViMOZ4weO/lCNvx0kztoRBL2W58sr9xWu
ySBuNexI1JGrTHNb1BAsgR4sHF/xMGHW2tpRi2D+lW/H0yqu9X/44VmV1Y+HQF0Js6jbe+1n84aq
ISmuuKTi5mqM4rBkeNoUxtmhm5plApPFZqXhFYnrkrsv4Lt4WBIuT1q8HTLcR6Bjx0E0ve7XYC57
jsNcLlRoThrguzzyIWgiXn/gRExPIpoz0xyIHh1uvhNtnzEqVJ+7WIictFnbutZIqZrWFScwWhnv
YHzM0+kM+v4m3J3KWyfuJSAHKHsup+T50Xz2aaHAx8GtLhldKNhUDQoP07rxKoQunR366SLBZDAA
h4C+L8a6cli/qTnSnS7xgLve+dp2tMlnUfg2Wpk16pSTcffvy25W/MQnxDaJ9ClQ5qgqfJJ0sQsW
CYoP79aW32YT5J6UGbyl7PddIr5Sq46x8x8OEA0Yyo2AqgT4x5as6MM01OEpBsS4vi7yAlSEOtl7
mKrUD/xLFWVQLszhh9UpG1cuika35I0N7ZQOsNFooGgFKtUBA5Mb81XEHsCVc2mMYVlgjLZrZ+XJ
rf2lHhpsQEFTF8XmezHAPfnw97ABroe/pEU+li28I+dlu86cZYM88gd8Dw0vCbQzvRp6coBQpBtR
yUl3WWwjM4hr733Ee9+22BnCCRdswXvcbeTOgZ94MKQjWSDqLBek+sFDnvJWaiQ+tiK5W8XOE3XR
40woM9KSczFkQmEt+oCAlhnaI78yYkeCSv4YW+acvAlFDhF+V2uBkVNsre93RFReRgdxVNkGHpQe
d7H6pmMU7u2kwkYAKVy0Dgtd1WFx+DjyAbM8UAziR+VX6ChsGMQh5JNZvVR5mJmGlgSRrT6MCQdW
TUISP+E3I2AsOFyr3PjxYH27DcR+8aLz6yp8q/lVGJyFeM0xEpPJZD9Az2M31QHQcOIoDFpHkiTa
cop4+os06PKOuyVS0s4jdkth3w9OpS3eddsWqPxILcGmXewH1OFKoS8RTENsjDD0Nl/6cDcuD5et
gZa2PIsTv5DdDpVBvGKVfLkqF34R+dVdF/d8567dWWp1LzCMTXaH4FQT2Vxt7pm3bVHlUOAsHLj6
i8jGCvHoYe+ynlhtYE6PDqiQU5eJK4GKJQLZqHaMvtCvamr7Oa1w8EOEl60Qyocto9YZarf2RSWZ
z/UyZ9U5Fn3tThfJpE3bnXZskCmK1UbIZWTWbzIp0WfEjhaEhhfxs54gimavyziGNQk/xafam/Hv
zCdfMf1njvW5H1GPja3Yw9+IemEzcgL2j+SYDKmW0S/1/tk7FCpxsBYX47Vf86hWXwngoKHhhYeY
gcKdJCnmuUv7kUosJwnbW6xtViQb1uCte20wVmJVEle/hZtSeMUjRxpvRJY6zc6jOPm+bLgm079e
4Jn6GOzEE9n7Qd9gqVkbgVpqAiCAUdM9vroqmxinBoc293M6jPJwvw23o7l5MtFEo1JW4JzNPGUQ
dNvMer/gYoHAb8AkOAVu7R5t3SXpwmTe6ueoQzL2NPn0L2BVPiu32sHkExqcuvp4IvJMLVzzQTjZ
Q/vr8vBcPq4KEhXlB68iDAxHo9BRwxtYlRaZx9UAXdfSbXIiwHPr6vf0xa4PtMW+KdKfki4e5pU+
N3j+sn7m9UDIVSyhciiLKQ4ncUBNqEMLMmOmT1vfknPZN6nQY8bl7qFabvRJT3jgCxxpPoC23rsx
4jjcrWe0TYffJRJb35xLNYWJmrkGdsY57U50iu7LFO50eXmR2n2tNJoRT8LZxdE79KybXHEEEQUb
BW9mbR9HzbcDRj7cUEEVQ3THS4v11gs/i02Ca/q1TiamuCV4iRGp/rgCAEg5wfM2hYxD8+oLoYra
/xUBPaUZY3E65jup9R13jBi7LseuBjSL4GRNGaz0zwokyKRSQ7ZlHGZYg0ihTg7sZ+ds0nEqahBc
SSXpl143tMzuXR5PHV+dyDDwRVenGrJDkYmEe8eOjHmaf4Jh3TAh7y70gAyufOoCRIkyAfbz9hPK
BG4s7PmQa0xyfDt76/op+kFCUwzSYgy59B5I0630CnuLs2YOk2ETRObEGPsn3pne0A48UvdOPWni
3LPfYBC4IHSyzyv/qZZQOhdJlDuIAgUH43n7U886Xejm7qOZyjkJkv7g6t+ceCmFMXHL6J3CUpqb
1ZWI3G9W/4U3iueuFAbmz5fmkyXhQPFs1QX5+tFn43LArQxJ97cZ/EPEZOm1zmNRRjt4LXmaXA+d
/HVOJCDp4PsvG6tTLeLPzyAYi4r+GggEJfZZg3Tlv2TxbO+AC/TxahDh1G1Wd6f+X4ZYcx6dwHpA
3C1CrNbfk93Ic+ZTfoxKo58siBwwNbTrj6fPH83vGDXp9gpAXZ4WLNK+l1kV626p0qz2GOzc4A0s
pJ/1fZRq4ycBQIf8nhVDalbP1XK7pSAeaS2mJjJbj0SNDvEunw7N/2l9I0nrY85wvynQ1wl1n5zJ
8m6BgBQ5teALOfSvkrKAxxO6HaVT25WaqBr+/HJI/HAh2+WluTL13LkoBfHeJ1mfGXIUKvjVVmkb
Sl0v/lUPXHtRtG8PNIlS/0Ml7ZqSUSbnXD2ZRgSmoBuanN6FqippgjK/lPs+bhRNSwQFq3IwvKm8
C9eNXsXNP5yFjSw95uSFD42qFUJLSzXAbvgM5H96nACPNFbvchcDVkgDCl4JCm5KiN2giJmS3FO/
8/fbUphlwMRjAD/GlSJBtRvGvgNVvIDgaN/yzkjTFg42aeg7fLb/QMordh2HjdtPEN2MoMnu0FS3
z+l6qKBJZxrWNcLEjmEVOwz0hMAwJTYZuRu5pccCWPlGcBuaKTOuLw7fGS3Mg2J7G734HlKOH3AP
JBqr4inL7seVkflh/e2/ZB34th1lOcvzG6AkiiFzrjBEbWq2Ha8lIr+NDyUtxETNgLfpxm36SgL7
Tm2FxfsphEzZrvy2CWTokfqQRTKBvwg0APRyFjFKaXqRr24wmM8JLlEPhg6povdjrpEQsIFO9Zup
tnyJcrQpOLLVKPMU9/XaB8SY3uwetC/IkTTWJzhPWPM+lIlNnmEqIYrJLn0x9HK3b5oD6++fL+g3
SLOdxKkG0rkNKNZYPHD0dhHGzgzuUC5gyA6RL9UuLfV7AUdyQuUYNzK9xKS3rwjEWZPCVyDxysLc
csGkLMKq2KeE1bD5uFfEr6NdGGQ2pC+FgjMynTruoKt+JE78xJ9m/N59e/BNtInqI66CDjWN20dX
sfuhx0BdUqJurRJXEoLWOyY3+demyR/BbISVhltBYbZvfMMZDAXUVGlWmA/XVhACh7ca8bEJnE1s
vSCQ3IKI/9pa21iQQGelJdblTfrycpgx3YeGe7RX3vtpJzk/8QZWWzbL8jdBLT/KACyIr2Ar09uX
r6VRQ5QIFMyx3QYFVViAysmGdPOr8tnESZUojYtItQNsci2tTbc4q98fon9z0fOkzd1WQSjm8yJx
WqEKKdnc5qXRddoq9xJW8aokRYZiw0VuylXQ+edw5VJR9zlI+6ImL+DjAkhZvJlIUBOYxyrVrap5
A9QxylGhUu3XaHABmTIs9PeZFosdHSHcBXmWKZWzGOL5lwIsIS4jETEU3wmIXeheh3+fHxqKWkpl
S3GVR6NUwIOTsh29KteH3yu6aLdtyfjMZpXOotzTpmkKeBxBJusQ2SETdGORbpz5iAUjFldhcZj/
528HwveNldiZqiIsfMMhj0FrF/qgFalqZJigU2dZ7qL5VDMae8bnbNc5LeQB6fqawVkNokMg837i
HMfMjStBck3Xspai1nzCSOxEoNEHO2toF2vmyY/1ffJhAwlfxDYQl51vPtpBGfWa0MAS5Bwgcr2Z
dQJlOEl+zg3Y5Sbwxi/JABu4sgaLZkcUBH1ARFyA89Ixhsid/dTBtSb+IVUHb8jj8w3ZTzYMRABc
y2JOcH1adpbFasM3aV/Aoi8j4JxoFhbsswVTqlbbkv9zK7kuMODojJ/JiXr7yrease8Z18tMy6rE
8hScy8/7LoTBtIYb3X5Wdu9/j52IrSnyFcncyrr9wLoUr3f9MhlfSDbtYDDk9fcWvA1dPGaWCRN9
n/xESDJgTY8ncwmmaMzP+kHYdO8W8DrsMrx4Of3o84PMgUlHtxNqXrEQABrsf02vAo3t5Szwk4IY
jioYNgztYG0pJ8QN7DwDio11Bli8d9s5T3ww+WqYm8fHorBtTjCc/dIxU9JuYzsJZp3tK+704nS9
W9Muf09835HN+4feKQaMvNJpwVu85sN2PzJLTDZXwPEzBjhrXv5SSr91ahJfd++/OiZKq+i9xp1U
8DrOkFuEkfsUByAOQ+URDi/dYJrdF6T84EG7fls4c1ngCwnSNIJuNrjY4Dh3zpSMBIFSt6wxDpdD
ilvbCe4Vrl40vRsLwFe7EbaOTc+sWWamPTNmcLNLM8M2BSwrSXIyb9IzCqgMIk36IghHtQr982PI
BiEdYAtiuORjiTiMRhtgA4Tf0UQW9/LpwVD/uNPM8EdO6DyFP26KWglJBwFzp+RbwkHJQoIQIBKL
wpXIe0CpjetZzq996bY8hxUJAk/PftSoNL9xHjkrWOLMa9F0glpPgp7F7j4JKA3YgOoo/cZC2Cc/
N5tjsWO9MMwcdUAHxYrenToPXp7gkySu1BmU+hQrV8wvvd167v3O9Js/mn/KNzZ3Oq2N5YD6hT7+
mvcWdFqckxofs46NVZyQYpH0b76njEitNk2vRWym5R+zYr4Mobjiv2n0KLha/ALb5Lh8uGQA635w
YIxMt/nxGIsWj1xfshUL6xoFVDwjPJQCWt8l67l6V3+iouj6htH4UHJzCMqiatW7+8dJdbAaKv0E
pARm72rmv1SAawC8/OXKQGbJi2dSZLAhDXF7/AfhbuWDhIa6VSJdBSCp+ZlGIUG0eGnxXICzYjOu
kxBNM8QYtQRdJxqzZvahVs+UiYfOUv3boyWdbvu7NGgUWSsoZ8NV5CZnXMQlk2WfEQF3iY7YVahu
9cS1D3DdN1zKYQHeuG/fAfv9gVpLBgR/84rIORU51N7BszEC/GnS4XYGyUkhKyxCFjc45chuYdTB
XtBb9cGsFDtEmNBGCub9xZAFWwfQLTvVCYiGUdWun51Ez7mySXlOk9kdDzHyiK8o6SnhyuAD7Fl8
dSQA5Pwm5z94xdOTu6VU450Xy+H6Vx9cGXYA/8eJJJDIO1wezTPhKqBnDarZvnDaTangQA+rqASd
VYHxgSiwFvdfcKyI9KidbWVwKgDoR73MRZLA5a9KXJhXoBuLCjM8z7ta4AqtB6p9sO7vfjOB8hCy
M2bUGSNO5BnustbcPrfsldNImXTdY9nugfzLhg9Icxj8qjY8XSCO7o87hV9MG+Q3rrlEBXXS68Aj
XYFG5PGqOXmb4OSvZiCGd0y0FTwklpMwQHUSRJV16l5tNuGOYFrcasoJA44aqpKpPapr34pnMbL4
c66ILi/qAH62l37bHZK7pd3bTDzRN1ovc5n7vnuPK+kQL1zWrCmMAqZ1aDCofGRvfXZu3WxSzIOW
29ZhRbhymwYOX6BF06ntkLCqeXpLHxTMciGTr2CJNwcxKv5/Y6egRmkyJuFuAQ8TbfI3IPqQ7ebL
IMHefnXsBBKMR0/ioVT6An5bL3Pl3X8QDc+gOnQMsb979eYKdvusufEIgE86Kt8JwrfJeUbzqaYq
gHmI75r3JWWFkMXVv9TLWYE94TePID/8Bg/WCXYolDTZm3Z4XexGbvieNfatVK/Ywz4wOCE/qjX6
subeiAshOyb8Sz6RYemkK4ImjEddSFY9OCvIJLa8owR6xoGUocbPBD1ypIFEkOabBJ12aRcoMMps
ld2HdwsBqbRPGQZpkfXUf4V8xkb9ROHUdt15u+1EH/XzQw8GRh+nLDr8wSj/3QMSRXLcZOLClCvi
8z2Y4Ej4ZeyIxWwLfLm4FTibE0RspK3b9g+9GodjuFVXD2DyW0L8BLNo2WEx9ZQgh967xRR+0/1Y
MbBC/jmDpnn4Qa4Eo0w9mZXDZA0k15vEu23BILdNvo55iHqlaPsZSxZRUYXaE5aDOQManp10mILT
3ToHuvbaycItuVz3EKT0jA1ZeA5xoZIEpA/51JrQNg7w5pV9EaMKWTi5Wgvmwcwm8vB8uhn0JwLj
FAR5dPFXxJcdcxnedMuZwkU6a/1Xy46XS8ZUvOu2zOp7/wB2LvIKDo1vusY5gVgAhghQdG7NioKj
YmlyncJ1zzc/h8sUzl0ry9Y6eUTTWeyuZW+vqhJmbnldOBeZN2cNvPYbz2YHGFe12JFH0m4mB2p5
7K1ri7PFkqUsb3o6Za8+M7wuek433fM9xPgNWFumzJ3mFkK8bAvBow1pQ8HFZMs0oKuAN+nMu/E4
cbn/u/7VX9MxmCyaYu7goWhixdKIz9UuoOSGoL9oi80bb0HNZYGlrByF/rxVSLjN9aSIszwuk02y
umc9XJW6znjI1zn0SeO1Cl3Sme6ab77Vm4QgYSWR3N89dc8pCV1FtqDBOlkI5lJS0dRnmkkqTXIp
swe593YlZKI69joHWdbnV4sTz7EEz7YfgZCFwB4mJycl9EgnQUj9F3ekBsJ1T0dUs86OZBCil7/0
mQ6F2Ov3zaEwkXjo34TNMTVMQAj58nItdBz4k9Sdz8XMg4VUB3soABX1cyy/k6exzNGoMGzLoVAy
kHQ+ojkl3F/WZF5C7dQT+lL+8WByIZ5sF5k3PXbSYmWaNeugRZwGU5UsJzI7InHQIigYWqHqvZE9
DDENXPST1xuUuk4x52TGNfVRr5tf6sJSsGL+U5DubCUkI86coLWtJfEFqu5Km7kPGlk7nXIPpbhH
21v6x3Boi2c8d6V1KVZPexvb87tijL3jo2CB3Kgs5FaesIJnuODIUOkgVBhw04j9riyc4+0ek8Gt
Ok9oGJ7u1z7/iYHJhlLxcIHo7Uv/L6g1yRQKqYWR+2spGoAbSTnecNefHGA2r0A0mHBQa6aL5LxV
dSyVRJRVTG/Rsyt/kpQKlo/uc2oCtesGBGMRvk+hga8ZnrwOYVu7VuelcES5VUiT7Mm/C2N0paQY
4y8v/WRUTMfkXNy236OXO+58q3vFhkLO3+m7aqzWjWO9Xn7nwjlD9obppLOp/2CVMqh0izIOmYoJ
1RjDDUZLDuU2srgwcfCUBIDLf9JaLfqpWHLc+kj8n09c0Ce/3Rzrc4zyHOhTwqm6d9daHLVgRPb7
/yqmMXCobojgV13HkWBUQ1gaSAY5kYccgo2aWjh2bWv8K1QE5w6zZZ0R324yw+uXgthDk2CYEGd3
iTGD9MHyRk24Nq+V63flUYGYDDK/ByXX+yHvRJFeG9Cdm4c+a4NotU+BYWAqoiHGXUJDnai6LaA1
jCZYXsFB18GhwTpvre3JyCcAHzHej2E2LIjW1ZKWoHLprY0eMa6qwO9iA8eTzgyfuhi3ZZUJKFSj
Grm2ldXWoE2KWFM+q2HPRYMC7607BhpEuU//RR/N5mdlZn93Ig9g6nP+Xx3+Okr7QW4xQ4mfJ3nd
qqrmYo5EBKjkFG2an9ZGckd1P9VogvisAt1Q4Tt/KsB3EBiWsL/1wsLKSrGvrxgfDIxxvvk7EZH0
0FnBFW8XB9UM+ppkCzpSDmLFzMEmVoKzx8lDIOFESpqJD3hBPz3G+zVceKwBf4nF91xLiBAeZTuF
DyLGcbq6jtr/MWWraJoguyGjGZtscjxrQhJx6eRHWKnRsh634MXSPJlZ2zi9yZGfV0erB5nzt0YT
MUJiUWLxT0vrSTnOeUtJsoz3FmSaJiwHyep2TluLup3y8u0/36ToS94VbYwariACloseZR9CziSn
+g9o+dKI7R4v0r4/fJZxiasFcLXwio8ToLPumdYHo8yrLuyT//YMQpNwPvbx+ochPkw81lU872jN
qIlx2v1oJKVAwMnyQbnmQb5p1InOQqCCmIizBpj9jTJdQBkbtR5YkX4cr6TISWyjB7m4vUMgXtea
x260t5rNSk+/hMnBgZayqCFSNj60nJvde6JsqBhD4NPeyOQ8ERzlsdSI4IwGGgvTARRneYwmpwaI
MM11C82Du+3WBhSzrPpZEm8rY8OvnAF/9hg+o2QOJirxZAhQQmGwyzJcJj/1pVuwYBH1ZPuC7frC
RgFhoYtx0UodSKImAxIL71/IaGNZphfXrLJ69EfdliWYYP4dyNOulV/9hlSLkmlVJ4rhCMU194sr
84k64cWcdauWIJQ/74yx0EoyY0qP8wa0oXqG6ET0K9oj8c89VPz9WItPDVOhCjMxvIk3+Wtk0lZo
W5k4u8R7x5kF3qOZIhjhQ4D+8WDEf+YA2ovkp8DfyGPsK48FPAOaFQUXUWhDAaivTcAUGxvybWqd
xzzvhCnrPuoNimeErdvrieyeQ6QD1vKFgp5nbYX82BDWpMIIauAAMpp7Ytk+0rIiQUuULTUVypb4
Cr3AOpE4Mm/OS5qUEmKFBFmaw6iYwz9dMVo05W8kYeXRbnMksBNAcyl1q/tp+Dcn3TSsKz91XSNG
0GHGwLdc4Ti0o0iZdccL59y4S5FRKdsVk+DynqOXDqAuyLyUCelLmo0hznbrRRIngJbx5R8R2mmz
lYWB4U9I07ihn5xPr2hj+bvVP/KokevtKMvDuxJhEIBuFWkGq93oN85yxHXKD6ta1Q2H7BJcgJUK
loipT1qY9S4Cah2NrgIwNjCGjT0HGDzJNTS/IY/4M6VzwZrrRYcJN2fmUOMfdPaBVD/Drp0nL05C
1TVbi+yOVHBPinPzDBkSv6BmivoC3TL7H7a/eatmCkAx1MaY0bPOZOymEMhzwI0ySYzKqgM8YhBG
ocnOUOy3MDBLq1kSQsXbZVdxri0r+cyuQLJAyY+rXhlgJ1kwDut0bUB9w/2vLnv16SxLllJhvACR
u5pffA3NAlmripSHX+rNdqGzr1YU+H8yX5+6Eo55plJCYxjgjI9BSLWB9Z/Kq3dq95vNqeP3UeuG
AgBSHonKg1uZ6CPthxzXjaT6evD0F/RU2w7OtAKtj5YdUnH0H5uPQZxj+B6ZsI7c/LcRIaXh0/IE
ruJDFqj/onJuBHxOCJVjeqq8jPvdHz73QSkOGvJiSFShgWFAMpvz8ywqM8LMCUQS9hfd8rGNr4/2
51McSS2FefCiCJE4kpD3kJievoNMOzZh8gjqBC3Y/obTYTP+Id04WlBg36UTABWdMOTQtU+4g/AK
5eqCO3+uSBaNDdyy51qU9rGez1VNUOVcyrvQNRPX+R0hPJPSg3j21b3L8aH5QY10pPG+OAlOThgE
GJWe5NHv0g2M434oPpdIZ2VjU7t8Q6VUkmyaVMDG6Ig0/hAehqpqqE5GAandrksC2uQVxV8vx9cm
1wzmdXJGRuqB/z9sNKszwFRNGvkj2aSKR0/ityLjRH78UkbcnrPof9XG7o62qbPTpnRAFNqKIqmC
aplq6u5seTrOKve/2tri+DPH3+SWs3cQEzIE9XUcG+830hHqPNGV/eG7W1ChL1jb+e8LpwnhrPoj
tgahqiyepI20u9xxUwXb1V5F6KZVkUZn0Ygarg6vNwzsC4D7OXERa0bGp2uVFbiUFsr0LMjPmJtZ
evu+wgv9vkcp+KGVkzkIw777XWItJ8NycnE2ftqs/lOcrU8AFIUvoZtzqESCLjGF4YCvV4ziOGn5
2yyYxl3SfXGzbOw7RTsYZzA3vO3P2vKsA0hZx8OPfb8ClbSJSGN1596L62ZUGtrl2vHEaK54NMv+
J3ToOGSGbu9P6oe5KoNxxWljP+OWjqEu5OZrUuffjDTqe2UkBJPrd+iA2oWKz8zGXeKeoLuB/fVM
g/00Gb0INo8GPguOJp+D7/Qqh+f35DHNyISYCc081as4MghXKRP/EUvgG6f2X0YSmZEbZ+7e71gg
10vUb9GDjVhBv+6NXkKrZHBQsINQCF3Ohcqcn9hozSl8UTXU5zzvXnmXGZpNqreUtArN2fJMcF4F
AJfiHU0lVFGiRBJ90Y0IZO2uNONZMwc+ArGtPzU8vXwZpNFGAoJzfT985Hk42S7xt/kIOawJMlE+
wYUiXnXhRVmkfytAiDMDzSnBQGBSGzRpeKWZWCaOyxPv6Cebu1VwUwPap2DvOkXdDiaEvCOwdb5m
3mxd3t2j5AEarUUf9qmJ10ERW6R7UNCBXBSBiHFHfZu1nJ9xwHsBbNPzFnBz0q7I4HDK6z84eliL
pE7QnZo2pUrQ2wukZrivq46Kfsb8puZpETyHmbsa2Swz0FBq4SB2o/szgcmi0iL0k3eF0OPHtskF
Jzr760xjWqdNu0JGZtB+AS+nqL9OKOrpbWNT8DSSBYKC3gy7if0EbpMHkMvv5nOpDJWWhiLPQ9ey
9tyEDAwqPKOIgcVrkVRsLCqq8LvkYsFu9feCoMl0Lv87gT0g5o4/QHJo/agMeKtO4+AtTdxWM94q
O0KDeu2obJplcoi8bfnEkkoZcIayFAfhZzXUl6D5iHS7E6a0IE7RNo/lLk0sycKIvyNEYnsYES1/
wG/dG+mV88rgObBaG0amyc7WVHIBFoA/uNY5vChGUXSPcixu0/rS4O7QjbkqhLGWCT1xr6P503UE
PoMkk/NYCkZe5zBSKgGUxtUX4BkTYA8z8SCeTUMixTot+AagWrl9G5yF5HDZ1HLbJlkzlJzfp7aO
vdrgRj8HhJT/mq2LclOGd2IlmpqW6z9jBEDN5LBjrNBj/U+2z1Eh1pRlK3hUfUSU/V7neZLbOR+U
w/eXwglFqhGx6UvhoE00Cdwv++FKbXkf8gP1nbTHo2g1mNWplW4RNG03ecgv5LSCPXj5ELkcgOE5
7rXiXeaxSA/4WVfUjTFxVh2Gmect+X5Ib/gJW+t2m7X8kv2jeAeHm6nYzzlyoilponjNvVkCVeNc
T9LtT6Iyx3GnU91vwufqdP5kDqbePMkwGb3Jj/ERHEafdOm9lKo4GBfV2WO2ZCIRgcM5qsVpvAt1
SAE3qbyFgZvr83S2ADZ6Vzqabozymhkvm2hleqYY7+gY3K/YReRIpjMCtH04qj2wexegTmrKoXbx
9szyd1NQlyY9GR28KS45aU14fDuLH+g7uxpPCZEh5wQPdIn03xLr9zZp5QCQ+TcqR9aBZY/pDWzP
i+PTGZAz+w1lVSs8dnoKOZakWPgQnkZAWRdbK+G9aHf/e6zG5lBuvnwnTkyZ6XZ52bf5rvYUkd8m
I0V3yPso+ZFN43RMPZEr8T5lpOskJZSmz4OqWty+vkI5Wai8nwQ0oDyIl76KSKVP7Yl4y8Tk/sD4
9UXyfVlSoGhHO+61FK/0LhGK9pxj6RQdoC3utJFkmnWFOWzz0UXt3xkvF1tpl67m7p0WrAxno/Zj
gDLpafD6TSuXHH0/V4x2LU7XPo/cQYVrrHknG36MrsOVmOKpCYSubO2J/Un96FOWctkg6oZ0SYnz
31fbMpRyiJBt5WLsMUiNVEKSDa4zoHC2GRL10jBXe75qEZcz0xr5KxiyQdY4GsA6i8+e4gjRWxJT
3BuEX+n0KEY7YvrgMIuIdOV9yTQoLe8TspsUIwsOjFtKQgLYSq4ZxXoxYn4DOXn6sl8VhYCMgYeO
WQp0k+1jz/NExtSUr89sYQ1UERz2wq0ccgxJy6JbLOoBdOvCu362yv/abYBD625d92fjQ4yyjGES
WVfDz8i7JeFOnfHzLSx0z9Pm51p2EYy8BjQCIFixVX8lsypezATnaU9owwMU52SBLcohuxfuIEG/
8pFIqeyTI4En+YnYShnVTbuZwagDNDpdgRiPp0CcUXCyxuGQqfDGMsNMZOqtZFgEbf635x/l4OoP
ocuI8ToBxVhSjZVAE4VJ8dBJa3ftlCee/OvOQaxtpQqrfJSkSSYiCy88I718R1JnjMcONPgXXUU1
Q15D0iWoUAy5DNfU1sDphvI7f7T9/iHKct1OqkB8kSnkHPk/LZYv1TLPLNsB+uparf2DmG3sGXvT
tOSfPFKHFVfR5hlyODqklV3soEYc1Vv1ktW7onNY3hrWuE5DMnT5NMTBwlEb2rc6eOLa2458M3GY
28PgxmGZ7qz1msq/ZrdFcTSGXUNfWXdMizBCINNH+LDDUuA4+esA/zEXHqm+2FG+psiTnK8/TSyK
sQGcQdPoq58pumQi7YKS3dnAZY38y2fuMeiTZ1MW9ZchUXPigIa/FKkVt1sxGu1WN41RAXBwG8bT
FU+OYBjzeijRgEi9wl3eeuohpq6ZCEZ5FdNTKuDUZerDtj4jjQZ9/9x+lyOkhS+PRbQvEMdJhZeY
5z2x9DIG0PLeAoC4/SlfmTTJXjq3n16b+L1xUsGNE2Pc1TAyCZHJZh/+/tjnVbo5UoEE0S+nYYjN
0OsAuDYTjOsvd3aM/1vWG31t5uPyS5zGzrkfZ2/4DfbPNoefcI2da/NUY8u6naBOzpEXsv3NmLmS
gi806Es9pl3371VcBvisChLWs4I8LgEcHwtP8MYHyxqD7CoIBasJytPTtFu6QEgp4NTnBiZwS2ii
Y0cRb5RTSjaJEMxJzueSfNzCldeGHIj3yvHE60kPczRlxlVEY5asBUbxMBVo6L18d6soMX+560uI
q09dWDVi0UKb8vhpYoYWaRltkJDqea3eUdZ9SOehwN7MfVGxOF7L3MnDevvA8NnpzFayeUgVFE3v
jx0DmkLR+cMzaGh7Tk73SZTyprP8fJJ/xf0B7ucNeBJ/gKwgvieWl3OgUXM2yMbiKZVHruSBh/V0
fu7PRly8UvmixBPXur9ua8m/XKg4KFyQHbwi2/NcPJolatbm/YQerVDz2aOZ3qDCfCu9NkyM49/K
nGe+9sM1c/Ag6vCuL7fyZN0q8lCyFPnWUaOby2z/zxN5AufCAeRNNzoVRBSELqgwpiWWcs/rwoOX
ZDTSUfboW/01YU2RUckfL9HWVPbdzlIawr1IkSwN6HXD5dSvrcrCTs29bduD1UFSvPgZru6ShshE
fbij8YmgoMKbQuCYyF+ggyf9uk1OqfkV4heYZF7LgiEK9lr3XYU3Dsy1txs1neP5RADRkDCuxJLM
VPKLnFcZbkDmNpzVwYa9Ek/r9516RqQhm4qn9e6PXtFLyaD6yvZTw7XMlNVxlvw3pZddG8DA/vEf
xv4GclijQdtNFjzFzF8bMdHXt8gW8OC889ZFM4AmiFl4SOhViLrm/TJocFCOrjEwYdaxcgmh38Wf
Kxv7ZSixLBDlNdsTnK7KOaMYYBZo93PvVFv8xnhxAIYzkhrIntywnxS6p0hQrKKhXy5rAcnUbyi6
3aesduj0E2fny6Jb9a8wuH56Ztw5XX209p/c7TEmuUboI+K2wl3r2sTSHMBjxkZIIAcRvALzQh4W
DUI3SIrECCxJT2EuJPpXC5BUYBZ3aaSUmCtZtV70nRDZqp7hPJHYuiZL5HHaKzvdiv99yvusHMHX
xOanDiA2yUOgiPEvmG05dfvAK3LhpgF7EFPPyMFAk8tvMnJZVTqR8CTG52OohfrisZPaWOzRznr2
avRAFGnJfe59VvtQmLAzQxxAgvJOKOIQ/nSA1A9p0Sp1U5x+6wUTqNzzeoO1nRMfvBouuz9xQQ+0
DTJM+qxa2/R6bqx4J/xSrleEq2LfOybTtRN8shrHjunWw5YeXggjtdC6p9i+SdzUt4xz2FI3K20H
TGjTCXB/wa2njQkRYJDWzJ8LUq+sOpphH/TIFcl+0IdF6g7zq+ibPEm0SU0iMcvc2CeRHN65Kl9S
Pzxq41vK9XxQBGp6a5e4sYaB/noU4bcD/7sXc1eK8PDhE+CX1/23x+qlplx97n7Q9rzHcP6aq2+x
1DgncFo7ShrGObR48yi9NBPJF5+Ktpr0HsneQFK7v2BfZAHg+xKjIHDXJbOp3wa2+WSeJmoxiNW/
7EAtTfBYZmC8RgR9btS2X0xgI8UQbGulY8NAvWgFp0+Rag6F0p6eo3B8rYdEo94DOICo4pklTcBj
FKvLB25c7DDzL24XF8iVv9vvz8sOd+7YW6BvOloQ1pyuKyCgZRbhY4nB7bnh4yND2o0IlD5bdiy3
Dq1bBENheiRmd/uB9d1eKC0ZA2oyuoVVR0mefIe1CsBEWoskL1WTY+GYS+fIXWEwVVtJrrJYX7oV
+lukBwK2oeTMsz7AdL1wRbaoUS635gtYZr0Kd/qVQ4Jz2HmcaYuqMb/t0uCaSQ3dr5mAx3AuSBM9
T0m7/LIkFHENFZnEJ2AtO2CJbCUOSICfPO7uDPUNL7L5RjMMKvsNn+cJII3cgs/6oufMdisyF2DK
xKN/C5rdEjbZPuE+bneaO9gJeOOIN+PIoEve8z6rfm/f7os3oHYI7uL/Yn1Qr9maAFamnJyMPSgW
7jbVxO9H0bks2Po7sVZB8qc+EB0py2w1Cn1Y4+OtUvNqsbSNFIxn+Qc127sB/nTzbKpfv/1hiPZa
qHcenoiMvVQmHcs9sN2NqdKTcHAS6KuXz9n/06Lz0ofy5hF/zSWrz9XkyAN5ySC+SmVptBUMFmST
etRjjxRIO/ksy1OOurREEP8psAa4LOqJb90chbNe00c2VKUq4hCGk5+spRO+285Pf53Sbvcyyf6G
urCMIwh+Q51ZQYNLP8nEGS8Rhyb7TCPK8k+afkmM79V22LiXK2G66eUz10ix3f5QTI+kppnWdups
AXx4MYAM81hYQt1suOg0DYDXdMLrNqN/Hdju8GaHAEuHt3Ry9CW1DnFwKP1AbPak3u+vugWSQ3TJ
G9NZI7Q85Q0KkEwa+yWSoRpDhJxaiyZU6DUjpkLKUCFHyIR9cq/2v17ZpbDxRpnif1+lj8Pc03zI
7GqxVu2f/OGcjlu6/RZ6/oUD6LLC3p7wTv1Nvme2C2G/tKMHaaqIBxV1ek6vYnOYd/aUSY6FPOBI
TU3/xj4QqCa3/xt0L2ba3b4+wV6kEXcFe5WRzFZDFfh05nw2cVSkWNXUeCX6DdZw7fZBmjIcdU2c
EZf1gpMqHJ/VZcGza8U1DIe1Xo/GeyimchUgP0ztq3mK4CKBGUQgoxmedS11k5V3v1kmbiG7Wc8i
cJ4plYtPvZpHChq0YSZ+8C+tcEKXRE6g70lx1jDwZZGQ2yXqyzQJciP8+waRJM8eqIpLVPo9R24/
O9TE94BNkFHLvbR1f5ZOPMGmwYRitoaLcamUObRTTWldNXwrf8R5ogUkoR1Xao44VuTzt1I0+07x
w9ddWyFEr9GkHYzCXSc1rDT8gdhfwnGYWTc+2r3XRibO5cDZcJmB0y8h5/yl4I9rTGSs9kuINsVQ
Fi8MhnIi25b/NUscla8T5EOQ69GV9xkyT68yggihnksh0NRbVXmISYO+Iitv2K5bLTaRITH1sTPp
uIwOHpfku3wGV8sGfcEWeXO++jQF15NCA+IpX7TzjgAvS4zR1Ma8/qpVkSArxKpV3VCSFabFpXVk
e60iHcc5aszeX0DulT+DDvgeFVV3gOedRVIXZxA9uMDG/qjgfI6XXDgmuSzB+YiIL4CuVIJY7oEw
yJj7H9P24w5a+LxAEAFj3E63xNLOpjzMSO93fsPMyCUxkkUZgQhRN6h/HazAuCJoawfqkJejI40D
qSJ4nXFE7Q2Q2vAumOkAv2jbZF0gVTIGbc3iy5xPwADB97ELr2x/s5D42GiLkwVPBby7y5EI1y1u
HMgSAGLCE1is6mOccDEBAyVmBiDLczvcp+xzrdwze34dKUI75nlZIInKv5nivbFfhTObInWlNynJ
doIjccT41DVcLK4mVbSi0qUVajbprtYLroTNWIooExDJjynH2rFqSpv4hUP/m5+VI34vLz2GRelq
aSRhbpkoZXtX5fkdGKbpf+zuu+50iLqKHyioXQoCdeGDyIeRU7TxLKo+5Qm8FmW62S/z/N/GRfag
PKNHt+aYRl/hVrqb13NfaEpwpHp9XbEYLIW+VLgUMy2OGHBU+/ZnWHcb7uTBoDMl93gkM3Mm1hdX
wKXLixBlfXVn3MIU8pF6L/W6VtmC4Wll5x7kPovJ+spPg6dK7h8s9f0+NiRnb3NBLwiUm+e6r5hp
o46nZ9F8itevpIxsdq+7HeD6GPYIONhp6NXxlMAb9157aZQBrfHMZfUePnMA6B2A1WlMj2PHIQXK
YNCf7PTh49ybSH0iTWWGGAvJ2n8eX1WLpzvqf6KL0pwQmvT6VZBaVELTzsw0SDxMsqPEUx8KHzAY
ONlSs4wCn4vH8GI90a4WaISDJoLJDq6XvML7lTn0uyL/UmhSpwbTORL0JUKt/pSSm13+V2Qy/o1W
WREDxTxzU4ODCzynHSluuSZrTedHBrXwNjEsaxWTyjrXaB8RUWQ3j+Y70eovA1WhwDw4/ABEU6Nf
6T4TE+V07U4wYrYSONUeXjp8xveBPbn8dJr310phb03yO/cdLshNlWFElEdXijycGlvxwTwYl2+P
H9kcsJZsZJOrA5fJLc37OYi5IeqdgS4RZOcSUB9GhW+gdkR0LL1FiaWg6rPrzZXWFCtWM5t1SUXQ
OvBywnpbbOlvCCgx+mBOyNnJBhC7CBFzYuhcn967RUstuqFGaSgA5mDcOQgsc9BM430UmmVJOKTv
u8mOLFrqyJcGl1+YKt6eNC0sSNAaNffFOCWN7zyAmNEKU5chC0Yz0FNpowTtZICO8siDeXe4t6Nu
dQ1QS9xijip0t3DzrNPIMbZ0UZO+k3N90jr1oXoBmcyELTyOMGRt/PvZlRj9iTO41zQpC6vChoRc
ss+q4cj+uZTWvutP7gFGy7YJ47vkCik1AIYnZZ4rCi8VQjsN3RvonRZiswg8zW2BUKT/tPSgR+f+
DnUFE3AL1WVNmzKnnWP450UMT5X0t/snROHu6gE+1vQN02889uj2zsnZLpk89mxIf4hB4LcZsKdr
/LYRkh8AXqyk6DnyUPQKcn+gc1vh8mD11XYGAgp2dzjYDJEOdw2EDZYR3teXsGZ5tljn5CFkWKkM
+eGlYZ/GMErPm+EdCTd/vO0bylSkT/t6wXNNMnCUBE7E/wp93DynXU8IwiCCU/NoZMtj8fGjvIKD
IlQrk4uv8evV0mCzszKJeBFqMH8JhSz/jwaD4HpcCyaIZaewb3y8Rxf33K6XRrf96DDiBB+CRkr0
7Zpp9O8zSm9RGj/kG9Jjegk7ExEbHxy8siJOXaM8zfCCQy1f+v2mbs3C747OQeYPlgNnp88g1txQ
tsWE79GOmNLPHkMVKCpYbz3CFNCBnvQLCxLTPfQVZX3RzEIIsehrOWbf4K2UUn2t1FxNNgtvt9vX
tADWXNNpwCfc8+oboTUwtnZku/k+8wv6NqZ6hcc93eT16EDjmHfvvksYY6syTe8j4MpKZKTgmtNv
DKl1B/691POK749HXAMaKF0WOQEB1P+pm+jbzwjYqSHqrZC/iDiuQx6wwjBgMlEMVpX/Sq0Jd75a
Pkwc9eiS1DHYJkCoqq7JzWVLnO9eTeKT+TzrOZqHzxxWpe3YY+UVQgH9UXvVxQweIyWHSt0p3vdQ
CeLysQnnk1UpC7q6jkDy5s73DugKcbm3yHG7wSda/xW2Ll05+mD9j59TFuIXduSDUcZz4bBYMFqF
lNcmNHFEbX/NJhowhXK68QZNYV7LLRlwyeU0mHacYwJngeWkT8ajb9eUGZc4Cv17tDMx94ms9VQR
Dt4hJbAr/+Y+xxwMWPx7u58RizWM0RFJhk/3HdG1aNklUT2uD1JIhi0IrXznasoWzDSpw/27y4he
/+LIFQoJbXyIXTtBbPDoGJmC+JJEjBBwNcUCTsVzJEoqoh7PXLi7yt4jnSTBB9xN9wuGb9VW8PfL
ua/oWJve0a3YTo24Uq/V7pByag64xnCfUY57gDqWTIWTJ66sM8h7GdLuPaYgcRLuKH+dt1jdfV30
rhNROtKrX4k1DyGC/GcEC3L3fseqiOaVt+RMDRge9eSrS8nZAZVGAgK/rVGCh3MT2XN6qErELvGR
oWvvsMtiO8ZY1n6rpySG9YkQfbm4MvyW/KLf+W5WtGPI7yFAltOXUzgbnaq2jJ0wT1bARwIrRYHu
Z+FSbd02SM+4SaeyKH+5qcRjLK1BiK5zKbdGrdRkSyr4aDWzWb4Svh+wTnY/iYxoM3lj+Fi+vZ4j
S43mVoMtudlyGTIgcRLDqs/Cuu8QnxKf4tQx7RocRgxRrWZdKcxu+tzqRdu/+YtpA3VRsH1kUG9C
ZLbs5/hZTeeiVHatetdxILVEj35u8vuBn+VtcUUA96p0Ut6FDh+nyB8qHJTehu6FV5LTK2ywDCA7
/j5ZvKipaqhtqVwkGjuT0ELeEThLlka1bVeNHPISQ2+tQJzQ8vYxh/hLSW3X1Xt2NohrR4iQupsS
6ZSIvgU7/WcXlgquXxBtAm5KIXxN0PaGiuVz2ZnBkBx6Be0a/d0Eyjol9xmi/SReMUig9aVWXuOG
784KFXO/mp1GSCfDemUvpzlhB4Bi6+nX9TL21i93mhsJnV3J1Jf8YlpFv9+y7IWZTuaMJyNSPikd
OnUJFPq528cGJrBysUMA8n1kCASevqC/nAFhn1XkZtdqrmgAhM08RscseCl4XfWQDRqoYv2SrAYb
DtROZlrUrB0EvruEeA2OKkpWHVszIk96sVGyQmUFkJXG5Pa8whHf03/x5ICM1XzHLlUIpzjdcK1t
jwBIexndNSo61r92c1sQTJws2DWzgE+A5ZB/4WZ6hchhHQUUmT5VK/pTedIf7rEgMH+rka/ENEpm
hnkAiNkdmEsOdwTuwhYfnzrQHHdApX4HFWymO9GmMdNv1QiO2pasJ2wNMj1XCOQWZf52bch486ME
RxgJf43ZePPOIwa9CcYwVuP4Rfs7aXbGTITLx8I0h9KR15mCrWMJZ/Oym2LUg/5ZMt0hfakZB9wR
/F9dC2hYHTD6fIe7D2+VEu/Pl8IwO/RjD6JVK4jCzP4llZVp8HLainup6jV+sEaheRV8ORduO7qZ
ARujXr/0IsG+moCjksm/JT4FxCtJHCaRoFEhbwi5Dxh4YKRal6qjYAkf5TQNYGKnDN/cI7TNee3w
PotIKBDKjMJrmIVYDxyA4wc/9X9BYlqfDq1E1xOP+JLibvZaguPe9eO0c7JfIINOMR+gTiwSq15x
5zjuGqrpWBl0Kdfi+j4RvDu2eJzN773YUUh1LJjfzmu4Ox0fIRgIHf3NP+pVMyYWa8gPAHeJAI5b
aqIMPu1bo5yga5jv5yFJugdRZIzlNZtWjRlXFVv3+6K76XMRMhhGgMHbIJ9KS+KlDXSQ58/Ipe7F
G3ZcyhKYqidpA3X5iZy4F0iwJ9j1uEacsJTUaYAJJoFf8H9ky+fsNxBNDkubblXCLPB7fM+RDvb1
MI78kHyYGzMPHXG4QsEtDSR65c2tkiIhaIBSRi2ACETpsvE23BKqzf2yjR4obrcjaXU0/w65JLav
IofX2SMLyejr0wAK9ei1pgilFv2bZDufTgWrHEovuVUoGAHTZOAKwbcBV3YL3K4t1tbHEqO5t8+t
YNZV9QATfg6V1bwCtzOAfsZtE34f4ZpeGKSO/WR3VNDRKT0ApLTdUrVGZTaQSLUF1q623h5tl3VR
DEMHucNseP9Zndr8/9Csrrdkoglh8oXofHZZzLI8fPmdhDsIkBTN6xc4bTFBauNjqCXgVHQUWk3R
7tDzPT9tI/pA9F8ZMd1M3CIXBCZG46x/tAkyzcJkN/pQCmEjjzu0RdzDQK9pupPgN/M26epyMWQb
0mPK7CoMxEA8Y18GRozQxoGgDw/89Hf6/4UdeEO6FvU/ENFEcmhRxXAbqGqlaoQXCVEBysSDXY3K
FTmpsL5gU6PbPcQD5n9J0lcmyT8ZbcFvgfuPwzt5jDV1ruy8SD3SEvF5O8LoHWRWmCekNoGCdvIm
3mg1F95e0PLd+F9EeoG+B8UdD+c090bCOtjAM7vJZC2Kwqixd36f4zhavpoHptP2esnMwSK6BXh4
fI9Nb52kaGYUyr1doFp0Z75kx86ylCJvspTePKRMDRE7MNLtLiTpDqWvi5x9/brCy/El7ricXf04
b/aC6KgFWJvztg0bZZT0Sy6V9vDunmUtFRoCTQUMVEBF8h75K6LYIzDdGcP6bGmxbgWrlVQ8+xxw
T79w7tzWnfGcfO6RWzkLvLwNkS8BX3Jf+4WTl9f1i8ZTpnclQ1DjpA++bAq97e9N40UhBuHrMPf+
Bwa0wGfKefwvX7JvIPeVd/ynRjHf7dY/UIFjLfv2h6JNN8vkl4Rvx0K6oEkpZvUHPnnTg2z7B3xk
dQL4iNTRBzxHQxcBxKPLd/YtyxOOvv/hmWWoVu5XNJca3DlwKj1xeWje/Hw5efADXX957WTLKxEM
ZeF8h3ucRBkZ7zv9cygUlAWc8dDOJRfbE1RVR8QfAv1srN28P0CBCzLCGfVNo3+ld8NI9WhSx9zB
s7ZKyu54gEBXTi7b5zb708pPo3yNXbRsVnUaWvXaFtO5LHTxeWTX1KMPzs/t44U861wUbxSHmtLX
XyRfBGvZ4WsmRMkfsbzEqo6OPsweRlf90gwhwEg9dsxgpPP7u67l2cHdBPlbbRIoS+g4GBAqu6mp
vkP/tpHuuePu8TUGbNeKYPtpPHxmUKWL321MomycJ8CQzBoOlyOQimX0MxyQXsd12RLqps80S18S
e0cHo9hKApJWSNj497nUDnBMs2rgSmim6GIMA+2SW/xKKEAqVUrBsVuD7SPY1+C5xEGTWpJ7dkU3
vjFwAJP/AUWoU2wHkH9K9PPXe/rPK/Taw5jofMQeYkHLRTx1gZgKYvlgjeWWXeXZJ7nAS8PHkH0d
S38pn/7hbmm6lH7FhARQps/mUXBsDzmXh3kHJCB4G6eiFvhjkbAjuVeDTe8gfs8ONYIdLEVmZDYC
1vbZxf2RVVyo6XAbF/FC//hFDwahBLO7LG3sgE3wb6a9+OHPtLfkIWgK5Ui6JSwrPaSEjpfAstUa
WvnI3+qCETnMoINK5OV1Bi/kJeSOLu3RJDeqollXeXxu7iHbye1ezBqnf3MtmDIxakAi5+fps+4t
LiHaUUrHvt3RqY+Vgdc2SL31ouHqk8007bbSMFMBUSeLOYG7Zp4ejZICM3IaFwoVF+zzOVMW8XwA
1pZrVGw3CLq/b2f+n0sfSW9O68YBVy+q0OfJCIUP5A79MFbgUyulhms8zQnGMUVPzXIcNtMm2QBr
FCrIQ87nlLbTlBmuRS2+KL3u4MCPaiqhuVr2U7MvYiUO4+kMB/uA+djqLPuoFxFDC+5aHtMameRW
gCAs9UOz/ZO6sqLhTsF3gELC+YwB/oLaQ2ILwApN+nG+MF1keI6Hv6wSL7H110dkNff99SAxyM4U
YJq21i/fKOiDn4ZN4zSmgqrKods+jSutEj/BKBHZoTxH7ZxxujrpgyjlvObzIP7hWR/bFKok7Urm
B4cWJZNZv37JCzpR5CyhorVuovgWHxUdmJ+xcHR1C4tH+uXrCcnthbV+WqH85JoB03oA2KXRimE5
xIRUqODoLFQ8ermFfyL4Dv15XAdA27hr99Q1gkoDw7wU6DJnum1DIFPsu0q2VFmt+rwHi0cSHCH7
HI25xNxags7ihm5IZBNDh2SyVBvhd+drdKP2pe7YWfShytZyJ93fRsfAObw+f1aWwofDk9WinQOj
pE7LMfuIagpchvGGa+QfS7zMP9+YtJqkNR6ZbrOGMNQwERMurlA5mHv9vyKlzrMZoI5AJr1B/0Oz
EojiLGSais68bPRcp7n5K23NiIHZkCHuU/wO3qY668QMMa/L2tWkQ07R/yHNhzyykce3VpIw0yY7
s4jByHxAqa6/gJHji3Dol54GwgF9WmK/nGJG5rksQAScUIEq2647Z0++w4Djirq9pZfwEMzqxZOx
oSEZ0kfqAeqJrO09LH27WYMrb4C2vHfpvKuVchag3H1L13J0An4cETbFAhw1L4c0DDf/xSCCSUXq
5p9/ewa12LGdF9/KkkaabMg6+HvL3l24AgId8PNxGKYz0Smf17VGYHfFLNptBdfdGEVmIauGPqzk
6Ga3v4Gho2EZGKP4cyX+lvV4+buwYKuNlQ0CeGW8IpQApVQcqHSPS/d+l224hig7j/Uso7WuGUiM
fX0IV+n/jb6Tun74QiYzYHCAbXa+gtRQpW6RGNy8clWHlwc9slVRyBEkgnvX+cmPmmC+IZ3+vbXL
eJxxtMe6U9mN8J7n7MQSjB8H4j/zHT9vruy7m48hn8DY1xPCyLO1HgODfDz3gtpPCHr74fSuB7jn
7CwEmrgPUKFinGSkl/zeCvidVobTu73ZCLociVPDqP546uqqmSisMfszEMFrZAb0N3cBpixa0wsn
YWY0L7Rt2hdLV6M+m7C/2ji4+4gN7eIEZOBjGV/CLoWYihk1gn0M5v4eXPuqvEf8F61gysAbyuvc
tle+E08edXexNTGFF2Y1/XDbp3ddOZa84TWPRio5vsNlhwKtfZkyr98JL2GUxYirgFXqAzvrQnJY
u3vG+amFDR7yKxBM4UU1q3giGAqDLt0MW4SGoy9J83oLju8u5y95j8EEaWUzioUjBjLs9FxX/Su7
clD1SO6umC192NlcMt4JBvOQAzLnFLt0SsG+FAQSkIy3lVcHT9cxyTzXw9ysq1IYp20k2VPcRKgW
hSmur3ay//kM+MZgRn5mWAir+d0GYfVCFB1ALeUCsGBA2vukVTvhdDKmA/R2PFvfaazWtHaRnWsn
ze788XG1q/qJOFuHeQPt8bF8ZxRphU6C0GzLSx3bJUa583VvZ0fXbTzwXkOy2UDGONi+GRwC+7sz
jLCzvLHGhKMkjdATzGT+g9pMN/cMc6YUz7v/rAQvD5z++C+t31/Aw3TRNkxsPwWWtOqr32FZ7YhQ
Yrtf3KqfphSIsIA42zoZ7Ez9TzpIlbEOdcW2i2MnaSmdtvBzCEKFjUlrDZNJUdoiRz5a1ybu5rNJ
hzT8raQzs7vYfhSdm4IjaNN3wrVUlrqHDVoHyE5EPRr0gyAtkLgSTLMMd4RqY0x/LZXgb3jKjpmn
EKT/O5jY9XNpCer6OhH9DThl1iq/+HOIsGmDVi/ukSP/w3kGCq9IcHye8WHt26qoPaGrDQwwq0T9
ER3eWh6oIr7KBWlvoIKTpk1aTggzTSosQXd7TzLPQHrh63GC3QYJfrIxgxs2olbmGyKEBzXvSefZ
3Wxv8gCP5bVw7TvlnCqgPmIpzGUnEnh9djeyj7T6gQ+bvbhqJvELrVupIbybpYfydnPFpp8DRKco
WF7yBqJCH9PAZd33cWOiDMxIqJhusxvGgJjK/pwr7Szkq4TRf5lHDBEv7BQ4eCo0qvYXhfmuLIgS
AJfbhPxoxygyWseSsu1Nw3WEK9156USrNnnfJFZb8uQ3/aAWfzT77F07yiUeWhrXMAac4HQ+qRr9
uvZ8Fr5RwK/Ber7ogv+jObUXMUx295bB99yT2MMNznAnNLj3Mu7ILQbJ0RhMM1jgtfjjSoMVZD8m
JPjaJhcjnTTRLM0ALdHRk6z+0LdnJ5n57JOI7JeOab/qNuccrKfF+lMZnIpDBkGIxTbPYyoIFbGJ
k0fBX8T3Qqe4t7UnJqPRSsYgkKYV4hrSFPGfbHY17swXjKq2sVBOpw9TPVXMUIQ+dT/cXXOGXJbG
3AgRp6TorBYzNazi3W0Z6V5Ccx4sgCPU4fRzlWru3YNILAaFtmf8kU1Le1GdUg7koBPbQ6xZVweq
SoS5XOC4vmju0tUqZEaKVDIXvrkAiY5LvoL9R/Gil1kW3c7mXI3xZAcsDup4vkyRTk8yIxDcAINa
ehv3hpYMrWn9HdfdVsJ/SbFBi4oDANjBc8v2wXZ4UIBYr0FMz3L7Y2lQxqB830O9SajuPXjCnk53
/0cr/8cwTtloG29l4HLuR8TRXKiSsqukO03dkwih4yFVZjdkKagTLy5GUUf1RaISE443n/f06Hsb
NmXIK/Weproo0ipMfYudBMn+uZFuIsRUixk91JN3I1nf9xPixeTDMggty4nkhLoWS33uSoWNFNL2
5G0DRQ3q9UeWEaqTaCEdCdlUDbdKG5Y1WUzqkV3nNqKHzqRwz0T3EtRLfTL1MAhguJ/i7SxEpEUQ
95W1NLV5efht/CsUw/ToZxa351whwwbkET0jUcGySNnfL+MFqBflpr0KYIhNK9E/xF1KJXJlfFil
lM8PYPoyT2Qz1l68vpaK7h/L8HsTTCLoQsB56PI0bXKCscrEJIvb3lSNUkA8/thC27wBPctnuZkK
GgLbyKoV0k9lcGveaRBpah90UGcOvZFQJp2p3B6sTX3LQt9sMZ58BIAtG+eSefUn1QFtnZPcipGz
I7eMNMmmE2BWYMTmKsVOw8X4ZOTMlCstxgfSTtYag2fbkKrR8z4IDK8lbzBRDJPNQC1RwSUbyMZ9
a+aAuNzoRV+EJvanWZbyqwZkgi+3EU9qcUT0kp1ry7Opi4fVh5R++Evm73NllhvwMFzIK3DtM9dH
h/zDrFNYTOvSUTVXSfNvIuFPAsYrtnwl6jUlTSFbt44H1kfGPdU4MXkkoRxpl1YurK5hlSIrQPRM
AtNIc+PTjTX6Zq3S1Lm6N20STWprUZYeutbiZLLNrEI3Jakvn53DT5lxu6p43exs3cVYfruDrpZn
LgSNY+Xe7rVzRMG/ebmX/92/CHO6EZD82JvIuT/8fMpGKTL4lXb2oGBpswC6g6phrtJJ1eEBOnFQ
UAC3I9YQjJpon7TBystV4SWOgAik09x4ho8pDDuOsTG30xiNmDjIa+38uxszdbb45a0E/wMaZ59u
1Bg4IiY2cLMCdZu8BGbIInrSnoRYKDtz4wq7zZ4VyBRD5LcS15QwBYV3nkDsr2XSaoCtgNAhfVor
Jbd8XtfzfdJi/8Lp/uKNLviwbRaJAoWXae2ht0/mnv1+jo6DdlbaZp4Th6Iv8BLkvclFAgGVR6FW
LykYD7nfZYAdwVYNcRthRVLZIjGsLhigFe2ciIHF1GtOQmcFId2tRglduRibTW5qPU+Ufx82o+bi
rhJIYfR1F3W+mpsgsAYXxpGPm3CUVvZ9ZSD63xYxxLs0M99tu2IbiKZtlPlKEK5TZsNYtKQ/ilQ2
L0gEoCHOIR0j3rPfUFy1U8J7jMDGds4CtxW3H5naUQ2/TVB8+ab2nQYRvEyp5mvYH71DOv4CJK8j
H0AQuGX/mn+PFkvTcr+BP5WNhOR64nH1aTOeC0bSbRJt53VemP3YjpQqYSmxGzkRlDvzMfd64Qaf
oh3r59wjqxJ1QiSDaGVkIyOV7WRCQDFY1z2N84W92fpOpbZCOko+J+nzgSw4afTNBv2Bj3DleWwr
Rfl1iGwvHPsfRBQZonkztdEw2AhRm2mNrxq7eC1iBvAATWqM9IeiC0WikgmdeIRdU7NXXrSok/3s
mtngQGO1GB07WstLkZDjvu22eW/kQ4qfWjmWc7nhfiynzk99edvVwWQ7OLkBUG6OqptlLD5pUK/K
7SeDwr0lpxwwrAxTZvK5NvfeLs3fDBgkqvB61ff023eIoEar1qm17bZdHVNdrYtqBo+sHA2zKc9Z
XhdBaky9cj/15EWlDKIPnenPH+AtrwWH9rfX5W8yzot2F74LZ8+63FFnU4XhsB2cIrEZXLpQlgET
a2Vk6b42zk+LR1B9p5L/8oCOOcEyNOUuiqCDvAHw06hbQWaZbRe/sg0imQeGIbnAmzXXWypZZFLs
yTpqIu1+NyJEZ/0XiZc2QqlOxTSNJMwlf9sPCyxer2DXC6sFGCAixyTAzpcYatMj6umNjUyxNt4/
VpRChtUN5RWjuV+HZEIylDiR8f2mEG3d5wLztz3/QhdKm++M4n3WgZvxQR5LHTXM7ZaG61y4F44K
mGp0Mz544RjV4xAXRwceGUxzieRjxNYErveRTYlMybcENistEAQI2Tgre9sTwadiIQs5GwX0WLnv
f+GwBugi1rfBpc+4eOfMc8gRyT1vAMaWn1Dcaw63KbW98H0lN5ovLrNNptNY0z6tTMM6mKhwNS5N
K5JszY7wANPSJeFuso1cO6YFV1jT8i/KN8TblQMidiI9+VVgIS/rmxejLJTONfHQD5LXDM5JUz3G
d3sKqPCsfN7gHu648Zq4AEHcav5oNdwBes0fFv0bEFO2Gm/w4Kuvh26WsxgjeiDK+cp3odjqKtlt
ovg4NOYHY0NQvJOJPs+mN937IjOwL/tO7thdh0uHoWszWLGAOquagBG5zR8VVvJN7yvyEUMrEm0N
X1cJKySjpEnZNhBMrQijVw2BuxD1BnNI5Uc2d+3i4SdXofIdca6DIjR797hGgOx3q4ffYFL9Aipg
g4MBYxcJAJbXt0G9Q2I1zS1DSUdIjO2honKtM54fpkTYr5ENjNAG0+M+YJpbW3hx8YDeHkaIwvkd
wnJD7KGrpd/cjkji5RZwIW1vpWQj0pQEXSoSn1XJe/ut2pSvFf1Q+W/scC/Ztyyg2dZ5cL0RlsUX
GVf4nvfN6BDJNZackpDdBXhlBbj6jyliSRKInvdN2BiutdBRWUy1FI5TEkBzGgdD/B6XJD94obRs
QyWgyeH/nm7gQdP7ZfkI4NgxF5s+thRAvBHWRr7qGW+3enkj+YdDNLBeIH6nEys2xRh6jDCy5R+l
Mubdm/7QLa2Xs+gZloktO0Rbf7GCHg1bS4RpI+KtmHFJ8nyyNKgG/fk7QfK87BQf1LfaQClsoKuZ
8gAXQjmzIXE1WneGwSbxjZUWmJhoqpJxoAjHR/pOo16/U4F5MoRakdypXfC54YB6YPk6/dgF7frQ
CEMnPGri9UYzbPfLajzz4zJmmFiyVLGMDcEewpJABifK8XHubU0eQMom8U4ztuCIgDN+ezoG2xy0
tKZFZ/n88xBBZD+4fSz8x1zhLIHgbw3/46Z+yxPpTjSaXUDtPzcRkc4XCNi8Diw2x051ZnPP6kdv
2Z8hHqI0Q8bskfvWzZr+SxEcFNDh0Zp5mErucTxRJgzNyKlplQsPZn4ysMZ/qNPnZiEifPq1PSrl
oGRd+y6yHg8KIRhznbDhSy/Ru/5hrsBSJoZVd1TjU7goyjX1rJbgpm/uxbgAEwnYq6wMAPjvyYic
n3TMJ1E4pdkYtBFWswFLnocNMBiPbqNgn8m6G/Lw8HSMm2Oakum5RVdrSs7KWbLcec8wUIDmzVR8
GiJzgydPBGFlwAzhIOYyn2LxXRy4E1bARSbspFFG2QO6ljZcmbEeL7uDfsTcwwkyg5H10fgulizk
bBZbySKGE3OdfrgjKRHv7qXF0qbHlxRO2TYlUIlspl5U1SU0I3zS+9m+6S1vCt708nAgFxJNL/sy
Uolkzn3OKJrg97OectUQqbfwZod2WaHeMiAg4WiYd2icEmySZGQshdoeUQFhizWz0kCwQ3VB+KAy
CIyVR/aWmfpqfWnzXyzA3B2gGD1tb8v/bQewy9rm606cHqx8MGhUG8f64snX5vHS6aFjegZWRwLK
ZynOT5kpDruiq2Yi21i0IS7KS44QoyCO1ao0DNWllyNemoq72Op3BItsRfyq/sgQNIpk1ducLOTM
cxEbO6B/FGo2mOKgyyfgKS1pc6A31siuf1l5KGqo7d0xA0nqfA1KIsyXR6LVLAvseLTE1mkXB27t
QkGL+LE+939TLL36SqFSB+VBgrWszAKGZUUjNkGyZfe/qfqj7a2KZTl5/qovnV7T4F7nLY2wsT56
r90+NdeqD4To9xeMIgoVJ7PTxyHYPFnxxQlYRE6f3v/k/F39mZftaYQi7MxrkaDIJnpw1LOwTxYw
6kK0/OGFbMdi8nfLSrwGIwoONPVB4cWKCn756Gn6ch7qPAXL60Vmkqv/hCYopXxSl2U/IyKrhEtV
Jbj0yfAvnocF1NbvObYDWB0adRxNsLf4B+odM3GN6EVRUJd2d/BkWGy+t8i49xaD8albn36aFu+q
24ly25fEqe+iPri18yuvOMzBhunwPPzYw4UrnQCsc02sbHlztR1EbEd+CyYEakkH8on6AuoMWGvc
BHV7gVivMH3GRkUZj5J+NjnkrxxMTTn/5JAR4umjCzrsmPZDLBqb4BHAGs+cA6fuyfbkjDbHkFGO
72PlyA94Igf6wwCxcEqT7r5AicBymOMfs5uUaxL7rquGUozZTkL1ynFmu5mHLGPLYft9SYujQoJg
LsSr75wrdx4xNC9FhkgQqhKrpnlZbeJDp5zPHhe2Kbgz4XxGo03VzKY3TnGuJtB9Z808kSHwYatH
pjhCpamo3wvKXk68qGRLSz1WTY0RAQDiEQFQixj6ndikisoihYdEkHmZoN0C5tB8ScKEQqo/RvF+
gYV9DQaFwsi8ubIZ4pPlifa28auivuzF67I3wdDKJwtJx5oUnXmyw8RkevsN7nQa3V21lwHaxrzT
iQU096tJm7Ugwd55uKlZDLt/sLH2Y9m02Dhv4vg+XpmqZLR6viEJX6dPBYq6Ob4o6mgHGFUUo7fL
wq1d+3/8KqYlRdLkIAI0682WpMgC0qDLnxwg0a/ZoNrJB5dq4zkVxYd4NbxUAp0BDLtZll3/Chd3
4XLT2Ky115OfxCn8XVF9WT/mWZ6GQt5/9+i3juARfdoHxCngyFj3W3uWhx7iWEjQqeaoCNtklwrR
90MF+lAkU9GY3m3tc9LCxqzZ8FeX/V6qUcLs6L62AQr7ns65EUQhNfIkapwpJctVjZ8NkH/HZwNW
V8Ak6jkRpPQftigzkOcBAFncd/7g113EJ3HinK6y6L4Dd2tbPjAzT/58BTMlxBPUHR01hH8xEdV/
X0d1c11DujRQ/u3zxdnAX323BA/ePdcnQFxuQ/leSbvCZX0Ozc47O6nhSvG8k0H6uWYELEv+3po2
XMnOSRAw9fmFhf2woIRM69q5nPfo62yyswlttk/RgqR4Qi23WEffcD1vgw5xcmM7qSgkUpQrlnEp
e6SyrqNlMKSOnZUA+PAzVoFV6R341/QMnNB4Sy/9Kgcw2e1dLcnrG6Uj3KlsP9/RUKcJrVtuX+2R
KuhDSCcWdXpyapPs933doN9iNnKJ6RlA8anzXTXvN4cTEqehEFrPg3kkwd8hB66yzURXQV/h+2dz
530H6cPSWkNb6kfv2SsCK8GWm8XES6aVf6uNYMONYQ7niam2B8DI4v2z1nHNrjLX32hJ5MsvTgVl
yEDDoVe3k3ZCuSj0gnRXYOXd4QYQ7G/nXHGLz+TOMlaezcMlAjkphHLZBnWSE+kJosx7v73iPK8t
LoRqSlSZd2aZSDmsg5MZNe2/lEIScJQtnrOU8HGEBC60CpmgvRiJssRQIsMvfIwWaAw/REU+bxda
PliZ18gWOoNjnkiTmDUkqXdLfrpxiaInk8vKoMl3Zy8GVQ7k08xRb6hiR2YuWtekYOqyKwyJXdG2
AxwhMAr+dHuPe6wVablXMaI6X2shiooa/fhn2bfRKjS5DAAAzajdLYEEqbbh6tSW0VIpSdlwFw0b
dIpfHeL0hIQnk9BXpMg3R2JAElOC2TZsEl9IFDMTBZTYqhempBeTnVqG+Klt0UTxWRwq1eu7FWNg
7ymGMCsLiq8CJ5VoIwMrVAgwurjRuaumfNPV8XAOxUKiH9XNfh5jw5zNozczs0xVePVaxjiU5V3V
rYz9xTyU58ItcWbigDOgbQiwerCWsutrAdqU49k5J7IYg5h1Ysoy0LlFVptWq4IpZF2D49LJ0ARB
tYspAp3u1JBFo58lZbYEB9Lsl8fftaUzOYTFukV0OhHvccADixuTOG8/IKPjEMzfw7d4k0ahFbQf
2jtDNxcPpe9Yg6f4e7AsSFox06zk0kTSIxT9NVYrpAWyLa7qgThWX5oLqsZv0ZmTPMPMH8OLW6JW
wHYLKZnhGdtJS7rl7OgOWiAkxaygx9kMVshZRpc1/cPc2GbnflpeHY3+cznLECuKT5k10VMjYvBG
T/k3hHfzl+Znj6sr6c4i9JHrQGRY+gytAgWI94xL9iyLEoUIGXX0FQOdCjB20Dd+mvtNUvpJN6Pp
4JIoyUBGrzxKMq+EaBntAMmwRCO6Vv4OF+AZK3ZB/oKUWpz0T+STvaFB+o7wCYIBxQfneilBFjHD
rcmI4jtf7BIS5NCzDRkeChkR4tQ0xZSp58gcu0+UUZb4x830/OTK580ak+hLNPoik+LpAy+IE+fY
PUDhhrGJVA84VP6HlivlOskP+YBgS+yVqJV4O2bG8aewPPwBHYEZSCGy+fAm7ec7mXIDSC9sOhZF
/c7zq8cU3hCnHwPAuqZgTGMEKbZrbskXvtRDtIUlnnpdpj2LS0OYocTuL0PqDpcW42g1tTSzkDO9
whUnRGLpbCoKfzR82BG0/esK9SnaERvDr7Xw1s69fg8l+Wh9hJoXUyV3wrMh+/m9gOkVn41xooPr
xUBjftrI/QCK4Hb8V3RnY1jNYcHLpBIX2raF5D2VU8jbDBovUePA+xXrgXB1OWFABusk3mzzg4zR
17cIKIbGXqIPQizMIojj8aHU2Tvmyl7odHEfqJziKygO9YaHQS9KXdHUZeyhtuuv0J3uMCZ/SMGX
EO305kmYlenKqodln03r7pvffL7fIrql6K1V935mLC1QDCnt6AHvSqoFECJ/0bKoX/GpnQ4aF7x3
Nw2Ed9l7Lwvga1hAX2F8E420vQFyiLKl1DaN/3nMDj4Dl40bc25VJtF/09ZgXCZ78m5cKtUIdwHp
NEQ9/wxv8pv4bz8LkYC9K91ohbLErZU1mXGITWyRhD5+T9YLyRmNHdsAy31fJNvC7fqjGK+1MyO1
kEj/HZzg+c9eY1pviZs3BMTYjxDirumszRzr02e8vZhroioeuMxrVzVt9QlNNyQBH0T5cKA2L48Q
lzKR5tOWk8iRxX/O3VAKgj0IDdxwkjD8okCv4ly3HLLaY/SQtDczVKPopbd1O+g5M36ReGUVeCwm
RXG8NReNq979BRHgbAZJTgi2xCxaajdluhEOcw79ri0aF1NQ2dKYTMXtnRazgiQ9WWalYPLbbtL+
wHpe6E1ZAEWD+PUIZ3aH8HWu7EqCCulXL+wnVv9mMszx5TGOfU07dI3VVZ9xwVzmgWUZtTZDXa6Q
1qTyAOjxNws21oRytrswgVclgx0x6LXUQR/PvXeZTXF7pzS2f1FhPiYMbbcEJkfTeL2wlFZVkoNm
H4b4wBwCeZ5YY52tdWeq0Ic457ByldAnhazuTtU8zznN0b7Lv9nO+JTw42rSIKu6nds9erCmTPYj
vPzJgn+6vUu0Qsod/AAS
`protect end_protected

