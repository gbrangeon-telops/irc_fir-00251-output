-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.4
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : k7gtx_sdi_wrapper.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module k7gtx_sdi_wrapper (a GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity k7gtx_sdi_wrapper is
generic
(
    QPLL_FBDIV_TOP                 : integer  := 40;

    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP     : string     :=  "false";        -- Set to "true" to speed up sim reset
    RX_DFE_KL_CFG2_IN               : bit_vector :=  X"3010D90C";
    PMA_RSV_IN                      : bit_vector :=  x"00018480";
    SIM_VERSION                     : string     :=  "4.0";

	------------------------ TX Configurable Driver Ports ----------------------
    GT0_TXPOSTCURSOR_IN                     : std_logic_vector(4 downto 0) := "00000";
    GT0_TXPRECURSOR_IN                      : std_logic_vector(4 downto 0) := "00000"

);
port
(
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT0_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT0_CPLLLOCK_OUT                        : out  std_logic;
    GT0_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT0_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT0_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT0_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT0_DRPCLK_IN                           : in   std_logic;
    GT0_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT0_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT0_DRPEN_IN                            : in   std_logic;
    GT0_DRPRDY_OUT                          : out  std_logic;
    GT0_DRPWE_IN                            : in   std_logic;
    ------------------------------- Clocking Ports -----------------------------
    GT0_TXSYSCLKSEL_IN                      : in   std_logic_vector(1 downto 0);
    ----------------------------- PCI Express Ports ----------------------------
    GT0_RXRATE_IN                           : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT0_RXCDRHOLD_IN                        : in   std_logic;
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT0_RXDATA_OUT                          : out  std_logic_vector(19 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT0_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT0_GTXRXN_IN                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    GT0_RXBUFRESET_IN                       : in   std_logic;
    GT0_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    GT0_RXDFELPMRESET_IN                    : in   std_logic;
    --------------------- Receive Ports - RX Equilizer Ports -------------------
    GT0_RXLPMHFHOLD_IN                      : in   std_logic;
    GT0_RXLPMLFHOLD_IN                      : in   std_logic;
    ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
    GT0_RXRATEDONE_OUT                      : out  std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT0_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    GT0_RXPMARESET_IN                       : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT0_GTTXRESET_IN                        : in   std_logic;
    GT0_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT0_TXUSRCLK_IN                         : in   std_logic;
    GT0_TXUSRCLK2_IN                        : in   std_logic;
    --------------------- Transmit Ports - PCI Express Ports -------------------
    GT0_TXRATE_IN                           : in   std_logic_vector(2 downto 0);
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    GT0_TXBUFSTATUS_OUT                     : out  std_logic_vector(1 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    GT0_TXDIFFCTRL_IN                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT0_TXDATA_IN                           : in   std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT0_GTXTXN_OUT                          : out  std_logic;
    GT0_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT0_TXOUTCLK_OUT                        : out  std_logic;
    GT0_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT0_TXOUTCLKPCS_OUT                     : out  std_logic;
    GT0_TXRATEDONE_OUT                      : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT0_TXPCSRESET_IN                       : in   std_logic;
    GT0_TXPMARESET_IN                       : in   std_logic;
    GT0_TXRESETDONE_OUT                     : out  std_logic;

--    --GT1  (X0Y1)
--    --____________________________CHANNEL PORTS________________________________
--    --------------------------------- CPLL Ports -------------------------------
--    GT1_CPLLFBCLKLOST_OUT                   : out  std_logic;
--    GT1_CPLLLOCK_OUT                        : out  std_logic;
--    GT1_CPLLLOCKDETCLK_IN                   : in   std_logic;
--    GT1_CPLLREFCLKLOST_OUT                  : out  std_logic;
--    GT1_CPLLRESET_IN                        : in   std_logic;
--    -------------------------- Channel - Clocking Ports ------------------------
--    GT1_GTREFCLK0_IN                        : in   std_logic;
--    ---------------------------- Channel - DRP Ports  --------------------------
--    GT1_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
--    GT1_DRPCLK_IN                           : in   std_logic;
--    GT1_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
--    GT1_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
--    GT1_DRPEN_IN                            : in   std_logic;
--    GT1_DRPRDY_OUT                          : out  std_logic;
--    GT1_DRPWE_IN                            : in   std_logic;
--    ------------------------------- Clocking Ports -----------------------------
--    GT1_TXSYSCLKSEL_IN                      : in   std_logic_vector(1 downto 0);
--    ----------------------------- PCI Express Ports ----------------------------
--    GT1_RXRATE_IN                           : in   std_logic_vector(2 downto 0);
--    --------------------- RX Initialization and Reset Ports --------------------
--    GT1_RXUSERRDY_IN                        : in   std_logic;
--    -------------------------- RX Margin Analysis Ports ------------------------
--    GT1_EYESCANDATAERROR_OUT                : out  std_logic;
--    ------------------------- Receive Ports - CDR Ports ------------------------
--    GT1_RXCDRHOLD_IN                        : in   std_logic;
--    GT1_RXCDRLOCK_OUT                       : out  std_logic;
--    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--    GT1_RXUSRCLK_IN                         : in   std_logic;
--    GT1_RXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Receive Ports - FPGA RX interface Ports -----------------
--    GT1_RXDATA_OUT                          : out  std_logic_vector(19 downto 0);
--    --------------------------- Receive Ports - RX AFE -------------------------
--    GT1_GTXRXP_IN                           : in   std_logic;
--    ------------------------ Receive Ports - RX AFE Ports ----------------------
--    GT1_GTXRXN_IN                           : in   std_logic;
--    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--    GT1_RXBUFRESET_IN                       : in   std_logic;
--    GT1_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
--    --------------------- Receive Ports - RX Equalizer Ports -------------------
--    GT1_RXDFELPMRESET_IN                    : in   std_logic;
--    --------------------- Receive Ports - RX Equilizer Ports -------------------
--    GT1_RXLPMHFHOLD_IN                      : in   std_logic;
--    GT1_RXLPMLFHOLD_IN                      : in   std_logic;
--    ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
--    GT1_RXRATEDONE_OUT                      : out  std_logic;
--    --------------- Receive Ports - RX Fabric Output Control Ports -------------
--    GT1_RXOUTCLK_OUT                        : out  std_logic;
--    ------------- Receive Ports - RX Initialization and Reset Ports ------------
--    GT1_GTRXRESET_IN                        : in   std_logic;
--    GT1_RXPMARESET_IN                       : in   std_logic;
--    -------------- Receive Ports -RX Initialization and Reset Ports ------------
--    GT1_RXRESETDONE_OUT                     : out  std_logic;
--    ------------------------ TX Configurable Driver Ports ----------------------
--    GT1_TXPOSTCURSOR_IN                     : in   std_logic_vector(4 downto 0);
--    GT1_TXPRECURSOR_IN                      : in   std_logic_vector(4 downto 0);
--    --------------------- TX Initialization and Reset Ports --------------------
--    GT1_GTTXRESET_IN                        : in   std_logic;
--    GT1_TXUSERRDY_IN                        : in   std_logic;
--    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--    GT1_TXUSRCLK_IN                         : in   std_logic;
--    GT1_TXUSRCLK2_IN                        : in   std_logic;
--    --------------------- Transmit Ports - PCI Express Ports -------------------
--    GT1_TXRATE_IN                           : in   std_logic_vector(2 downto 0);
--    ---------------------- Transmit Ports - TX Buffer Ports --------------------
--    GT1_TXBUFSTATUS_OUT                     : out  std_logic_vector(1 downto 0);
--    --------------- Transmit Ports - TX Configurable Driver Ports --------------
--    GT1_TXDIFFCTRL_IN                       : in   std_logic_vector(3 downto 0);
--    ------------------ Transmit Ports - TX Data Path interface -----------------
--    GT1_TXDATA_IN                           : in   std_logic_vector(19 downto 0);
--    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--    GT1_GTXTXN_OUT                          : out  std_logic;
--    GT1_GTXTXP_OUT                          : out  std_logic;
--    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--    GT1_TXOUTCLK_OUT                        : out  std_logic;
--    GT1_TXOUTCLKFABRIC_OUT                  : out  std_logic;
--    GT1_TXOUTCLKPCS_OUT                     : out  std_logic;
--    GT1_TXRATEDONE_OUT                      : out  std_logic;
--    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--    GT1_TXPCSRESET_IN                       : in   std_logic;
--    GT1_TXPMARESET_IN                       : in   std_logic;
--    GT1_TXRESETDONE_OUT                     : out  std_logic;

--    --GT2  (X0Y2)
--    --____________________________CHANNEL PORTS________________________________
--    --------------------------------- CPLL Ports -------------------------------
--    GT2_CPLLFBCLKLOST_OUT                   : out  std_logic;
--    GT2_CPLLLOCK_OUT                        : out  std_logic;
--    GT2_CPLLLOCKDETCLK_IN                   : in   std_logic;
--    GT2_CPLLREFCLKLOST_OUT                  : out  std_logic;
--    GT2_CPLLRESET_IN                        : in   std_logic;
--    -------------------------- Channel - Clocking Ports ------------------------
--    GT2_GTREFCLK0_IN                        : in   std_logic;
--    ---------------------------- Channel - DRP Ports  --------------------------
--    GT2_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
--    GT2_DRPCLK_IN                           : in   std_logic;
--    GT2_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
--    GT2_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
--    GT2_DRPEN_IN                            : in   std_logic;
--    GT2_DRPRDY_OUT                          : out  std_logic;
--    GT2_DRPWE_IN                            : in   std_logic;
--    ------------------------------- Clocking Ports -----------------------------
--    GT2_TXSYSCLKSEL_IN                      : in   std_logic_vector(1 downto 0);
--    ----------------------------- PCI Express Ports ----------------------------
--    GT2_RXRATE_IN                           : in   std_logic_vector(2 downto 0);
--    --------------------- RX Initialization and Reset Ports --------------------
--    GT2_RXUSERRDY_IN                        : in   std_logic;
--    -------------------------- RX Margin Analysis Ports ------------------------
--    GT2_EYESCANDATAERROR_OUT                : out  std_logic;
--    ------------------------- Receive Ports - CDR Ports ------------------------
--    GT2_RXCDRHOLD_IN                        : in   std_logic;
--    GT2_RXCDRLOCK_OUT                       : out  std_logic;
--    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--    GT2_RXUSRCLK_IN                         : in   std_logic;
--    GT2_RXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Receive Ports - FPGA RX interface Ports -----------------
--    GT2_RXDATA_OUT                          : out  std_logic_vector(19 downto 0);
--    --------------------------- Receive Ports - RX AFE -------------------------
--    GT2_GTXRXP_IN                           : in   std_logic;
--    ------------------------ Receive Ports - RX AFE Ports ----------------------
--    GT2_GTXRXN_IN                           : in   std_logic;
--    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--    GT2_RXBUFRESET_IN                       : in   std_logic;
--    GT2_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
--    --------------------- Receive Ports - RX Equalizer Ports -------------------
--    GT2_RXDFELPMRESET_IN                    : in   std_logic;
--    --------------------- Receive Ports - RX Equilizer Ports -------------------
--    GT2_RXLPMHFHOLD_IN                      : in   std_logic;
--    GT2_RXLPMLFHOLD_IN                      : in   std_logic;
--    ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
--    GT2_RXRATEDONE_OUT                      : out  std_logic;
--    --------------- Receive Ports - RX Fabric Output Control Ports -------------
--    GT2_RXOUTCLK_OUT                        : out  std_logic;
--    ------------- Receive Ports - RX Initialization and Reset Ports ------------
--    GT2_GTRXRESET_IN                        : in   std_logic;
--    GT2_RXPMARESET_IN                       : in   std_logic;
--    -------------- Receive Ports -RX Initialization and Reset Ports ------------
--    GT2_RXRESETDONE_OUT                     : out  std_logic;
--    ------------------------ TX Configurable Driver Ports ----------------------
--    GT2_TXPOSTCURSOR_IN                     : in   std_logic_vector(4 downto 0);
--    GT2_TXPRECURSOR_IN                      : in   std_logic_vector(4 downto 0);
--    --------------------- TX Initialization and Reset Ports --------------------
--    GT2_GTTXRESET_IN                        : in   std_logic;
--    GT2_TXUSERRDY_IN                        : in   std_logic;
--    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--    GT2_TXUSRCLK_IN                         : in   std_logic;
--    GT2_TXUSRCLK2_IN                        : in   std_logic;
--    --------------------- Transmit Ports - PCI Express Ports -------------------
--    GT2_TXRATE_IN                           : in   std_logic_vector(2 downto 0);
--    ---------------------- Transmit Ports - TX Buffer Ports --------------------
--    GT2_TXBUFSTATUS_OUT                     : out  std_logic_vector(1 downto 0);
--    --------------- Transmit Ports - TX Configurable Driver Ports --------------
--    GT2_TXDIFFCTRL_IN                       : in   std_logic_vector(3 downto 0);
--    ------------------ Transmit Ports - TX Data Path interface -----------------
--    GT2_TXDATA_IN                           : in   std_logic_vector(19 downto 0);
--    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--    GT2_GTXTXN_OUT                          : out  std_logic;
--    GT2_GTXTXP_OUT                          : out  std_logic;
--    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--    GT2_TXOUTCLK_OUT                        : out  std_logic;
--    GT2_TXOUTCLKFABRIC_OUT                  : out  std_logic;
--    GT2_TXOUTCLKPCS_OUT                     : out  std_logic;
--    GT2_TXRATEDONE_OUT                      : out  std_logic;
--    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--    GT2_TXPCSRESET_IN                       : in   std_logic;
--    GT2_TXPMARESET_IN                       : in   std_logic;
--    GT2_TXRESETDONE_OUT                     : out  std_logic;

--    --GT3  (X0Y3)
--    --____________________________CHANNEL PORTS________________________________
--    --------------------------------- CPLL Ports -------------------------------
--    GT3_CPLLFBCLKLOST_OUT                   : out  std_logic;
--    GT3_CPLLLOCK_OUT                        : out  std_logic;
--    GT3_CPLLLOCKDETCLK_IN                   : in   std_logic;
--    GT3_CPLLREFCLKLOST_OUT                  : out  std_logic;
--    GT3_CPLLRESET_IN                        : in   std_logic;
--    -------------------------- Channel - Clocking Ports ------------------------
--    GT3_GTREFCLK0_IN                        : in   std_logic;
--    ---------------------------- Channel - DRP Ports  --------------------------
--    GT3_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
--    GT3_DRPCLK_IN                           : in   std_logic;
--    GT3_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
--    GT3_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
--    GT3_DRPEN_IN                            : in   std_logic;
--    GT3_DRPRDY_OUT                          : out  std_logic;
--    GT3_DRPWE_IN                            : in   std_logic;
--    ------------------------------- Clocking Ports -----------------------------
--    GT3_TXSYSCLKSEL_IN                      : in   std_logic_vector(1 downto 0);
--    ----------------------------- PCI Express Ports ----------------------------
--    GT3_RXRATE_IN                           : in   std_logic_vector(2 downto 0);
--    --------------------- RX Initialization and Reset Ports --------------------
--    GT3_RXUSERRDY_IN                        : in   std_logic;
--    -------------------------- RX Margin Analysis Ports ------------------------
--    GT3_EYESCANDATAERROR_OUT                : out  std_logic;
--    ------------------------- Receive Ports - CDR Ports ------------------------
--    GT3_RXCDRHOLD_IN                        : in   std_logic;
--    GT3_RXCDRLOCK_OUT                       : out  std_logic;
--    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--    GT3_RXUSRCLK_IN                         : in   std_logic;
--    GT3_RXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Receive Ports - FPGA RX interface Ports -----------------
--    GT3_RXDATA_OUT                          : out  std_logic_vector(19 downto 0);
--    --------------------------- Receive Ports - RX AFE -------------------------
--    GT3_GTXRXP_IN                           : in   std_logic;
--    ------------------------ Receive Ports - RX AFE Ports ----------------------
--    GT3_GTXRXN_IN                           : in   std_logic;
--    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--    GT3_RXBUFRESET_IN                       : in   std_logic;
--    GT3_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
--    --------------------- Receive Ports - RX Equalizer Ports -------------------
--    GT3_RXDFELPMRESET_IN                    : in   std_logic;
--    --------------------- Receive Ports - RX Equilizer Ports -------------------
--    GT3_RXLPMHFHOLD_IN                      : in   std_logic;
--    GT3_RXLPMLFHOLD_IN                      : in   std_logic;
--    ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
--    GT3_RXRATEDONE_OUT                      : out  std_logic;
--    --------------- Receive Ports - RX Fabric Output Control Ports -------------
--    GT3_RXOUTCLK_OUT                        : out  std_logic;
--    ------------- Receive Ports - RX Initialization and Reset Ports ------------
--    GT3_GTRXRESET_IN                        : in   std_logic;
--    GT3_RXPMARESET_IN                       : in   std_logic;
--    -------------- Receive Ports -RX Initialization and Reset Ports ------------
--    GT3_RXRESETDONE_OUT                     : out  std_logic;
--    ------------------------ TX Configurable Driver Ports ----------------------
--    GT3_TXPOSTCURSOR_IN                     : in   std_logic_vector(4 downto 0);
--    GT3_TXPRECURSOR_IN                      : in   std_logic_vector(4 downto 0);
--    --------------------- TX Initialization and Reset Ports --------------------
--    GT3_GTTXRESET_IN                        : in   std_logic;
--    GT3_TXUSERRDY_IN                        : in   std_logic;
--    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--    GT3_TXUSRCLK_IN                         : in   std_logic;
--    GT3_TXUSRCLK2_IN                        : in   std_logic;
--    --------------------- Transmit Ports - PCI Express Ports -------------------
--    GT3_TXRATE_IN                           : in   std_logic_vector(2 downto 0);
--    ---------------------- Transmit Ports - TX Buffer Ports --------------------
--    GT3_TXBUFSTATUS_OUT                     : out  std_logic_vector(1 downto 0);
--    --------------- Transmit Ports - TX Configurable Driver Ports --------------
--    GT3_TXDIFFCTRL_IN                       : in   std_logic_vector(3 downto 0);
--    ------------------ Transmit Ports - TX Data Path interface -----------------
--    GT3_TXDATA_IN                           : in   std_logic_vector(19 downto 0);
--    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--    GT3_GTXTXN_OUT                          : out  std_logic;
--    GT3_GTXTXP_OUT                          : out  std_logic;
--    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--    GT3_TXOUTCLK_OUT                        : out  std_logic;
--    GT3_TXOUTCLKFABRIC_OUT                  : out  std_logic;
--    GT3_TXOUTCLKPCS_OUT                     : out  std_logic;
--    GT3_TXRATEDONE_OUT                      : out  std_logic;
--    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--    GT3_TXPCSRESET_IN                       : in   std_logic;
--    GT3_TXPMARESET_IN                       : in   std_logic;
--    GT3_TXRESETDONE_OUT                     : out  std_logic;


    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    GT0_GTREFCLK0_COMMON_IN                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    GT0_QPLLLOCK_OUT                        : out  std_logic;
    GT0_QPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_QPLLREFCLKLOST_OUT                  : out  std_logic;
    GT0_QPLLRESET_IN                        : in   std_logic


);


end k7gtx_sdi_wrapper;
    
architecture RTL of k7gtx_sdi_wrapper is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "k7gtx_sdi_wrapper,gtwizard_v2_4,{protocol_file=hd_sdi}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;
    signal   gt0_qplloutclk_i         :   std_logic;
    signal   gt0_qplloutrefclk_i      :   std_logic;

  
    signal  gt0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt1_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt2_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt3_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
 
    signal   gt0_qpllclk_i            :   std_logic;
    signal   gt0_qpllrefclk_i         :   std_logic;
    signal   gt1_qpllclk_i            :   std_logic;
    signal   gt1_qpllrefclk_i         :   std_logic;
    signal   gt2_qpllclk_i            :   std_logic;
    signal   gt2_qpllrefclk_i         :   std_logic;
    signal   gt3_qpllclk_i            :   std_logic;
    signal   gt3_qpllrefclk_i         :   std_logic;


--*************************** Component Declarations **************************
component k7gtx_sdi_wrapper_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP       : string   := "false";
    RX_DFE_KL_CFG2_IN            : bit_vector :=   X"3010D90C";
    PMA_RSV_IN                   : bit_vector :=   X"00000000";
    PCS_RSVD_ATTR_IN             : bit_vector :=   X"000000000000";
    SIM_VERSION                  : string     := "4.0"
);
port 
(   
    --------------------------------- CPLL Ports -------------------------------
    CPLLFBCLKLOST_OUT                       : out  std_logic;
    CPLLLOCK_OUT                            : out  std_logic;
    CPLLLOCKDETCLK_IN                       : in   std_logic;
    CPLLREFCLKLOST_OUT                      : out  std_logic;
    CPLLRESET_IN                            : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GTREFCLK0_IN                            : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    DRPADDR_IN                              : in   std_logic_vector(8 downto 0);
    DRPCLK_IN                               : in   std_logic;
    DRPDI_IN                                : in   std_logic_vector(15 downto 0);
    DRPDO_OUT                               : out  std_logic_vector(15 downto 0);
    DRPEN_IN                                : in   std_logic;
    DRPRDY_OUT                              : out  std_logic;
    DRPWE_IN                                : in   std_logic;
    ------------------------------- Clocking Ports -----------------------------
    QPLLCLK_IN                              : in   std_logic;
    QPLLREFCLK_IN                           : in   std_logic;
    TXSYSCLKSEL_IN                          : in   std_logic_vector(1 downto 0);
    ----------------------------- PCI Express Ports ----------------------------
    RXRATE_IN                               : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    RXUSERRDY_IN                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    EYESCANDATAERROR_OUT                    : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    RXCDRHOLD_IN                            : in   std_logic;
    RXCDRLOCK_OUT                           : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    RXUSRCLK_IN                             : in   std_logic;
    RXUSRCLK2_IN                            : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    RXDATA_OUT                              : out  std_logic_vector(19 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GTXRXP_IN                               : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GTXRXN_IN                               : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    RXBUFRESET_IN                           : in   std_logic;
    RXBUFSTATUS_OUT                         : out  std_logic_vector(2 downto 0);
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    RXDFELPMRESET_IN                        : in   std_logic;
    --------------------- Receive Ports - RX Equilizer Ports -------------------
    RXLPMHFHOLD_IN                          : in   std_logic;
    RXLPMLFHOLD_IN                          : in   std_logic;
    ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
    RXRATEDONE_OUT                          : out  std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    RXOUTCLK_OUT                            : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GTRXRESET_IN                            : in   std_logic;
    RXPMARESET_IN                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    RXRESETDONE_OUT                         : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    TXPOSTCURSOR_IN                         : in   std_logic_vector(4 downto 0);
    TXPRECURSOR_IN                          : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    GTTXRESET_IN                            : in   std_logic;
    TXUSERRDY_IN                            : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    TXUSRCLK_IN                             : in   std_logic;
    TXUSRCLK2_IN                            : in   std_logic;
    --------------------- Transmit Ports - PCI Express Ports -------------------
    TXRATE_IN                               : in   std_logic_vector(2 downto 0);
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    TXBUFSTATUS_OUT                         : out  std_logic_vector(1 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    TXDIFFCTRL_IN                           : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TXDATA_IN                               : in   std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTXTXN_OUT                              : out  std_logic;
    GTXTXP_OUT                              : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    TXOUTCLK_OUT                            : out  std_logic;
    TXOUTCLKFABRIC_OUT                      : out  std_logic;
    TXOUTCLKPCS_OUT                         : out  std_logic;
    TXRATEDONE_OUT                          : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    TXPCSRESET_IN                           : in   std_logic;
    TXPMARESET_IN                           : in   std_logic;
    TXRESETDONE_OUT                         : out  std_logic


);
end component;



--*************************Logic to set Attribute QPLL_FB_DIV*****************************
    impure function conv_qpll_fbdiv_top (qpllfbdiv_top : in integer) return bit_vector is
    begin
       if (qpllfbdiv_top = 16) then
         return "0000100000";
       elsif (qpllfbdiv_top = 20) then
         return "0000110000" ;
       elsif (qpllfbdiv_top = 32) then
         return "0001100000" ;
       elsif (qpllfbdiv_top = 40) then
         return "0010000000" ;
       elsif (qpllfbdiv_top = 64) then
         return "0011100000" ;
       elsif (qpllfbdiv_top = 66) then
         return "0101000000" ;
       elsif (qpllfbdiv_top = 80) then
         return "0100100000" ;
       elsif (qpllfbdiv_top = 100) then
         return "0101110000" ;
       else 
         return "0000000000" ;
       end if;
    end function;

    impure function conv_qpll_fbdiv_ratio (qpllfbdiv_top : in integer) return bit is
    begin
       if (qpllfbdiv_top = 16) then
         return '1';
       elsif (qpllfbdiv_top = 20) then
         return '1' ;
       elsif (qpllfbdiv_top = 32) then
         return '1' ;
       elsif (qpllfbdiv_top = 40) then
         return '1' ;
       elsif (qpllfbdiv_top = 64) then
         return '1' ;
       elsif (qpllfbdiv_top = 66) then
         return '0' ;
       elsif (qpllfbdiv_top = 80) then
         return '1' ;
       elsif (qpllfbdiv_top = 100) then
         return '1' ;
       else 
         return '1' ;
       end if;
    end function;

    constant   QPLL_FBDIV_IN    :   bit_vector(9 downto 0) := conv_qpll_fbdiv_top(QPLL_FBDIV_TOP);
    constant   QPLL_FBDIV_RATIO :   bit := conv_qpll_fbdiv_ratio(QPLL_FBDIV_TOP);

--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
    gt0_qpllclk_i    <= gt0_qplloutclk_i;  
    gt0_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt1_qpllclk_i    <= gt0_qplloutclk_i;  
    gt1_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt2_qpllclk_i    <= gt0_qplloutclk_i;  
    gt2_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt3_qpllclk_i    <= gt0_qplloutclk_i;  
    gt3_qpllrefclk_i <= gt0_qplloutrefclk_i; 


 
    --------------------------- GT Instances  -------------------------------   

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)

    gt0_k7gtx_sdi_wrapper_i : k7gtx_sdi_wrapper_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000000",
        SIM_VERSION                   =>  SIM_VERSION    
    )
    port map
    (
        --------------------------------- CPLL Ports -------------------------------
        CPLLFBCLKLOST_OUT               =>      GT0_CPLLFBCLKLOST_OUT,
        CPLLLOCK_OUT                    =>      GT0_CPLLLOCK_OUT,
        CPLLLOCKDETCLK_IN               =>      GT0_CPLLLOCKDETCLK_IN,
        CPLLREFCLKLOST_OUT              =>      GT0_CPLLREFCLKLOST_OUT,
        CPLLRESET_IN                    =>      GT0_CPLLRESET_IN,
        -------------------------- Channel - Clocking Ports ------------------------
        GTREFCLK0_IN                    =>      GT0_GTREFCLK0_IN,
        ---------------------------- Channel - DRP Ports  --------------------------
        DRPADDR_IN                      =>      GT0_DRPADDR_IN,
        DRPCLK_IN                       =>      GT0_DRPCLK_IN,
        DRPDI_IN                        =>      GT0_DRPDI_IN,
        DRPDO_OUT                       =>      GT0_DRPDO_OUT,
        DRPEN_IN                        =>      GT0_DRPEN_IN,
        DRPRDY_OUT                      =>      GT0_DRPRDY_OUT,
        DRPWE_IN                        =>      GT0_DRPWE_IN,
        ------------------------------- Clocking Ports -----------------------------
        QPLLCLK_IN                      =>      gt0_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt0_qpllrefclk_i,
        TXSYSCLKSEL_IN                  =>      GT0_TXSYSCLKSEL_IN,
        ----------------------------- PCI Express Ports ----------------------------
        RXRATE_IN                       =>      GT0_RXRATE_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        RXUSERRDY_IN                    =>      GT0_RXUSERRDY_IN,
        -------------------------- RX Margin Analysis Ports ------------------------
        EYESCANDATAERROR_OUT            =>      GT0_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        RXCDRHOLD_IN                    =>      GT0_RXCDRHOLD_IN,
        RXCDRLOCK_OUT                   =>      GT0_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        RXUSRCLK_IN                     =>      GT0_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT0_RXUSRCLK2_IN,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        RXDATA_OUT                      =>      GT0_RXDATA_OUT,
        --------------------------- Receive Ports - RX AFE -------------------------
        GTXRXP_IN                       =>      GT0_GTXRXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GTXRXN_IN                       =>      GT0_GTXRXN_IN,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        RXBUFRESET_IN                   =>      GT0_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GT0_RXBUFSTATUS_OUT,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        RXDFELPMRESET_IN                =>      GT0_RXDFELPMRESET_IN,
        --------------------- Receive Ports - RX Equilizer Ports -------------------
        RXLPMHFHOLD_IN                  =>      GT0_RXLPMHFHOLD_IN,
        RXLPMLFHOLD_IN                  =>      GT0_RXLPMLFHOLD_IN,
        ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
        RXRATEDONE_OUT                  =>      GT0_RXRATEDONE_OUT,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        RXOUTCLK_OUT                    =>      GT0_RXOUTCLK_OUT,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GTRXRESET_IN                    =>      GT0_GTRXRESET_IN,
        RXPMARESET_IN                   =>      GT0_RXPMARESET_IN,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        RXRESETDONE_OUT                 =>      GT0_RXRESETDONE_OUT,
        ------------------------ TX Configurable Driver Ports ----------------------
        TXPOSTCURSOR_IN                 =>      GT0_TXPOSTCURSOR_IN,
        TXPRECURSOR_IN                  =>      GT0_TXPRECURSOR_IN,
        --------------------- TX Initialization and Reset Ports --------------------
        GTTXRESET_IN                    =>      GT0_GTTXRESET_IN,
        TXUSERRDY_IN                    =>      GT0_TXUSERRDY_IN,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        TXUSRCLK_IN                     =>      GT0_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT0_TXUSRCLK2_IN,
        --------------------- Transmit Ports - PCI Express Ports -------------------
        TXRATE_IN                       =>      GT0_TXRATE_IN,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        TXBUFSTATUS_OUT                 =>      GT0_TXBUFSTATUS_OUT,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        TXDIFFCTRL_IN                   =>      GT0_TXDIFFCTRL_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GT0_TXDATA_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT0_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT0_GTXTXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        TXOUTCLK_OUT                    =>      GT0_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT0_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT0_TXOUTCLKPCS_OUT,
        TXRATEDONE_OUT                  =>      GT0_TXRATEDONE_OUT,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        TXPCSRESET_IN                   =>      GT0_TXPCSRESET_IN,
        TXPMARESET_IN                   =>      GT0_TXPMARESET_IN,
        TXRESETDONE_OUT                 =>      GT0_TXRESETDONE_OUT

    );

--    --_________________________________________________________________________
--    --_________________________________________________________________________
--    --GT1  (X0Y1)

--    gt1_k7gtx_sdi_wrapper_i : k7gtx_sdi_wrapper_GT
--    generic map
--    (
--        -- Simulation attributes
--        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
--        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
--        PMA_RSV_IN                    =>  PMA_RSV_IN,
--        PCS_RSVD_ATTR_IN              =>  X"000000000000",
--        SIM_VERSION                   =>  SIM_VERSION    
--    )
--    port map
--    (
--        --------------------------------- CPLL Ports -------------------------------
--        CPLLFBCLKLOST_OUT               =>      GT1_CPLLFBCLKLOST_OUT,
--        CPLLLOCK_OUT                    =>      GT1_CPLLLOCK_OUT,
--        CPLLLOCKDETCLK_IN               =>      GT1_CPLLLOCKDETCLK_IN,
--        CPLLREFCLKLOST_OUT              =>      GT1_CPLLREFCLKLOST_OUT,
--        CPLLRESET_IN                    =>      GT1_CPLLRESET_IN,
--        -------------------------- Channel - Clocking Ports ------------------------
--        GTREFCLK0_IN                    =>      GT1_GTREFCLK0_IN,
--        ---------------------------- Channel - DRP Ports  --------------------------
--        DRPADDR_IN                      =>      GT1_DRPADDR_IN,
--        DRPCLK_IN                       =>      GT1_DRPCLK_IN,
--        DRPDI_IN                        =>      GT1_DRPDI_IN,
--        DRPDO_OUT                       =>      GT1_DRPDO_OUT,
--        DRPEN_IN                        =>      GT1_DRPEN_IN,
--        DRPRDY_OUT                      =>      GT1_DRPRDY_OUT,
--        DRPWE_IN                        =>      GT1_DRPWE_IN,
--        ------------------------------- Clocking Ports -----------------------------
--        QPLLCLK_IN                      =>      gt1_qpllclk_i,
--        QPLLREFCLK_IN                   =>      gt1_qpllrefclk_i,
--        TXSYSCLKSEL_IN                  =>      GT1_TXSYSCLKSEL_IN,
--        ----------------------------- PCI Express Ports ----------------------------
--        RXRATE_IN                       =>      GT1_RXRATE_IN,
--        --------------------- RX Initialization and Reset Ports --------------------
--        RXUSERRDY_IN                    =>      GT1_RXUSERRDY_IN,
--        -------------------------- RX Margin Analysis Ports ------------------------
--        EYESCANDATAERROR_OUT            =>      GT1_EYESCANDATAERROR_OUT,
--        ------------------------- Receive Ports - CDR Ports ------------------------
--        RXCDRHOLD_IN                    =>      GT1_RXCDRHOLD_IN,
--        RXCDRLOCK_OUT                   =>      GT1_RXCDRLOCK_OUT,
--        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--        RXUSRCLK_IN                     =>      GT1_RXUSRCLK_IN,
--        RXUSRCLK2_IN                    =>      GT1_RXUSRCLK2_IN,
--        ------------------ Receive Ports - FPGA RX interface Ports -----------------
--        RXDATA_OUT                      =>      GT1_RXDATA_OUT,
--        --------------------------- Receive Ports - RX AFE -------------------------
--        GTXRXP_IN                       =>      GT1_GTXRXP_IN,
--        ------------------------ Receive Ports - RX AFE Ports ----------------------
--        GTXRXN_IN                       =>      GT1_GTXRXN_IN,
--        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--        RXBUFRESET_IN                   =>      GT1_RXBUFRESET_IN,
--        RXBUFSTATUS_OUT                 =>      GT1_RXBUFSTATUS_OUT,
--        --------------------- Receive Ports - RX Equalizer Ports -------------------
--        RXDFELPMRESET_IN                =>      GT1_RXDFELPMRESET_IN,
--        --------------------- Receive Ports - RX Equilizer Ports -------------------
--        RXLPMHFHOLD_IN                  =>      GT1_RXLPMHFHOLD_IN,
--        RXLPMLFHOLD_IN                  =>      GT1_RXLPMLFHOLD_IN,
--        ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
--        RXRATEDONE_OUT                  =>      GT1_RXRATEDONE_OUT,
--        --------------- Receive Ports - RX Fabric Output Control Ports -------------
--        RXOUTCLK_OUT                    =>      GT1_RXOUTCLK_OUT,
--        ------------- Receive Ports - RX Initialization and Reset Ports ------------
--        GTRXRESET_IN                    =>      GT1_GTRXRESET_IN,
--        RXPMARESET_IN                   =>      GT1_RXPMARESET_IN,
--        -------------- Receive Ports -RX Initialization and Reset Ports ------------
--        RXRESETDONE_OUT                 =>      GT1_RXRESETDONE_OUT,
--        ------------------------ TX Configurable Driver Ports ----------------------
--        TXPOSTCURSOR_IN                 =>      GT1_TXPOSTCURSOR_IN,
--        TXPRECURSOR_IN                  =>      GT1_TXPRECURSOR_IN,
--        --------------------- TX Initialization and Reset Ports --------------------
--        GTTXRESET_IN                    =>      GT1_GTTXRESET_IN,
--        TXUSERRDY_IN                    =>      GT1_TXUSERRDY_IN,
--        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--        TXUSRCLK_IN                     =>      GT1_TXUSRCLK_IN,
--        TXUSRCLK2_IN                    =>      GT1_TXUSRCLK2_IN,
--        --------------------- Transmit Ports - PCI Express Ports -------------------
--        TXRATE_IN                       =>      GT1_TXRATE_IN,
--        ---------------------- Transmit Ports - TX Buffer Ports --------------------
--        TXBUFSTATUS_OUT                 =>      GT1_TXBUFSTATUS_OUT,
--        --------------- Transmit Ports - TX Configurable Driver Ports --------------
--        TXDIFFCTRL_IN                   =>      GT1_TXDIFFCTRL_IN,
--        ------------------ Transmit Ports - TX Data Path interface -----------------
--        TXDATA_IN                       =>      GT1_TXDATA_IN,
--        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--        GTXTXN_OUT                      =>      GT1_GTXTXN_OUT,
--        GTXTXP_OUT                      =>      GT1_GTXTXP_OUT,
--        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--        TXOUTCLK_OUT                    =>      GT1_TXOUTCLK_OUT,
--        TXOUTCLKFABRIC_OUT              =>      GT1_TXOUTCLKFABRIC_OUT,
--        TXOUTCLKPCS_OUT                 =>      GT1_TXOUTCLKPCS_OUT,
--        TXRATEDONE_OUT                  =>      GT1_TXRATEDONE_OUT,
--        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--        TXPCSRESET_IN                   =>      GT1_TXPCSRESET_IN,
--        TXPMARESET_IN                   =>      GT1_TXPMARESET_IN,
--        TXRESETDONE_OUT                 =>      GT1_TXRESETDONE_OUT

--    );

--    --_________________________________________________________________________
--    --_________________________________________________________________________
--    --GT2  (X0Y2)

--    gt2_k7gtx_sdi_wrapper_i : k7gtx_sdi_wrapper_GT
--    generic map
--    (
--        -- Simulation attributes
--        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
--        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
--        PMA_RSV_IN                    =>  PMA_RSV_IN,
--        PCS_RSVD_ATTR_IN              =>  X"000000000000",
--        SIM_VERSION                   =>  SIM_VERSION    
--    )
--    port map
--    (
--        --------------------------------- CPLL Ports -------------------------------
--        CPLLFBCLKLOST_OUT               =>      GT2_CPLLFBCLKLOST_OUT,
--        CPLLLOCK_OUT                    =>      GT2_CPLLLOCK_OUT,
--        CPLLLOCKDETCLK_IN               =>      GT2_CPLLLOCKDETCLK_IN,
--        CPLLREFCLKLOST_OUT              =>      GT2_CPLLREFCLKLOST_OUT,
--        CPLLRESET_IN                    =>      GT2_CPLLRESET_IN,
--        -------------------------- Channel - Clocking Ports ------------------------
--        GTREFCLK0_IN                    =>      GT2_GTREFCLK0_IN,
--        ---------------------------- Channel - DRP Ports  --------------------------
--        DRPADDR_IN                      =>      GT2_DRPADDR_IN,
--        DRPCLK_IN                       =>      GT2_DRPCLK_IN,
--        DRPDI_IN                        =>      GT2_DRPDI_IN,
--        DRPDO_OUT                       =>      GT2_DRPDO_OUT,
--        DRPEN_IN                        =>      GT2_DRPEN_IN,
--        DRPRDY_OUT                      =>      GT2_DRPRDY_OUT,
--        DRPWE_IN                        =>      GT2_DRPWE_IN,
--        ------------------------------- Clocking Ports -----------------------------
--        QPLLCLK_IN                      =>      gt2_qpllclk_i,
--        QPLLREFCLK_IN                   =>      gt2_qpllrefclk_i,
--        TXSYSCLKSEL_IN                  =>      GT2_TXSYSCLKSEL_IN,
--        ----------------------------- PCI Express Ports ----------------------------
--        RXRATE_IN                       =>      GT2_RXRATE_IN,
--        --------------------- RX Initialization and Reset Ports --------------------
--        RXUSERRDY_IN                    =>      GT2_RXUSERRDY_IN,
--        -------------------------- RX Margin Analysis Ports ------------------------
--        EYESCANDATAERROR_OUT            =>      GT2_EYESCANDATAERROR_OUT,
--        ------------------------- Receive Ports - CDR Ports ------------------------
--        RXCDRHOLD_IN                    =>      GT2_RXCDRHOLD_IN,
--        RXCDRLOCK_OUT                   =>      GT2_RXCDRLOCK_OUT,
--        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--        RXUSRCLK_IN                     =>      GT2_RXUSRCLK_IN,
--        RXUSRCLK2_IN                    =>      GT2_RXUSRCLK2_IN,
--        ------------------ Receive Ports - FPGA RX interface Ports -----------------
--        RXDATA_OUT                      =>      GT2_RXDATA_OUT,
--        --------------------------- Receive Ports - RX AFE -------------------------
--        GTXRXP_IN                       =>      GT2_GTXRXP_IN,
--        ------------------------ Receive Ports - RX AFE Ports ----------------------
--        GTXRXN_IN                       =>      GT2_GTXRXN_IN,
--        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--        RXBUFRESET_IN                   =>      GT2_RXBUFRESET_IN,
--        RXBUFSTATUS_OUT                 =>      GT2_RXBUFSTATUS_OUT,
--        --------------------- Receive Ports - RX Equalizer Ports -------------------
--        RXDFELPMRESET_IN                =>      GT2_RXDFELPMRESET_IN,
--        --------------------- Receive Ports - RX Equilizer Ports -------------------
--        RXLPMHFHOLD_IN                  =>      GT2_RXLPMHFHOLD_IN,
--        RXLPMLFHOLD_IN                  =>      GT2_RXLPMLFHOLD_IN,
--        ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
--        RXRATEDONE_OUT                  =>      GT2_RXRATEDONE_OUT,
--        --------------- Receive Ports - RX Fabric Output Control Ports -------------
--        RXOUTCLK_OUT                    =>      GT2_RXOUTCLK_OUT,
--        ------------- Receive Ports - RX Initialization and Reset Ports ------------
--        GTRXRESET_IN                    =>      GT2_GTRXRESET_IN,
--        RXPMARESET_IN                   =>      GT2_RXPMARESET_IN,
--        -------------- Receive Ports -RX Initialization and Reset Ports ------------
--        RXRESETDONE_OUT                 =>      GT2_RXRESETDONE_OUT,
--        ------------------------ TX Configurable Driver Ports ----------------------
--        TXPOSTCURSOR_IN                 =>      GT2_TXPOSTCURSOR_IN,
--        TXPRECURSOR_IN                  =>      GT2_TXPRECURSOR_IN,
--        --------------------- TX Initialization and Reset Ports --------------------
--        GTTXRESET_IN                    =>      GT2_GTTXRESET_IN,
--        TXUSERRDY_IN                    =>      GT2_TXUSERRDY_IN,
--        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--        TXUSRCLK_IN                     =>      GT2_TXUSRCLK_IN,
--        TXUSRCLK2_IN                    =>      GT2_TXUSRCLK2_IN,
--        --------------------- Transmit Ports - PCI Express Ports -------------------
--        TXRATE_IN                       =>      GT2_TXRATE_IN,
--        ---------------------- Transmit Ports - TX Buffer Ports --------------------
--        TXBUFSTATUS_OUT                 =>      GT2_TXBUFSTATUS_OUT,
--        --------------- Transmit Ports - TX Configurable Driver Ports --------------
--        TXDIFFCTRL_IN                   =>      GT2_TXDIFFCTRL_IN,
--        ------------------ Transmit Ports - TX Data Path interface -----------------
--        TXDATA_IN                       =>      GT2_TXDATA_IN,
--        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--        GTXTXN_OUT                      =>      GT2_GTXTXN_OUT,
--        GTXTXP_OUT                      =>      GT2_GTXTXP_OUT,
--        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--        TXOUTCLK_OUT                    =>      GT2_TXOUTCLK_OUT,
--        TXOUTCLKFABRIC_OUT              =>      GT2_TXOUTCLKFABRIC_OUT,
--        TXOUTCLKPCS_OUT                 =>      GT2_TXOUTCLKPCS_OUT,
--        TXRATEDONE_OUT                  =>      GT2_TXRATEDONE_OUT,
--        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--        TXPCSRESET_IN                   =>      GT2_TXPCSRESET_IN,
--        TXPMARESET_IN                   =>      GT2_TXPMARESET_IN,
--        TXRESETDONE_OUT                 =>      GT2_TXRESETDONE_OUT

--    );

--    --_________________________________________________________________________
--    --_________________________________________________________________________
--    --GT3  (X0Y3)

--    gt3_k7gtx_sdi_wrapper_i : k7gtx_sdi_wrapper_GT
--    generic map
--    (
--        -- Simulation attributes
--        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
--        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
--        PMA_RSV_IN                    =>  PMA_RSV_IN,
--        PCS_RSVD_ATTR_IN              =>  X"000000000000",
--        SIM_VERSION                   =>  SIM_VERSION    
--    )
--    port map
--    (
--        --------------------------------- CPLL Ports -------------------------------
--        CPLLFBCLKLOST_OUT               =>      GT3_CPLLFBCLKLOST_OUT,
--        CPLLLOCK_OUT                    =>      GT3_CPLLLOCK_OUT,
--        CPLLLOCKDETCLK_IN               =>      GT3_CPLLLOCKDETCLK_IN,
--        CPLLREFCLKLOST_OUT              =>      GT3_CPLLREFCLKLOST_OUT,
--        CPLLRESET_IN                    =>      GT3_CPLLRESET_IN,
--        -------------------------- Channel - Clocking Ports ------------------------
--        GTREFCLK0_IN                    =>      GT3_GTREFCLK0_IN,
--        ---------------------------- Channel - DRP Ports  --------------------------
--        DRPADDR_IN                      =>      GT3_DRPADDR_IN,
--        DRPCLK_IN                       =>      GT3_DRPCLK_IN,
--        DRPDI_IN                        =>      GT3_DRPDI_IN,
--        DRPDO_OUT                       =>      GT3_DRPDO_OUT,
--        DRPEN_IN                        =>      GT3_DRPEN_IN,
--        DRPRDY_OUT                      =>      GT3_DRPRDY_OUT,
--        DRPWE_IN                        =>      GT3_DRPWE_IN,
--        ------------------------------- Clocking Ports -----------------------------
--        QPLLCLK_IN                      =>      gt3_qpllclk_i,
--        QPLLREFCLK_IN                   =>      gt3_qpllrefclk_i,
--        TXSYSCLKSEL_IN                  =>      GT3_TXSYSCLKSEL_IN,
--        ----------------------------- PCI Express Ports ----------------------------
--        RXRATE_IN                       =>      GT3_RXRATE_IN,
--        --------------------- RX Initialization and Reset Ports --------------------
--        RXUSERRDY_IN                    =>      GT3_RXUSERRDY_IN,
--        -------------------------- RX Margin Analysis Ports ------------------------
--        EYESCANDATAERROR_OUT            =>      GT3_EYESCANDATAERROR_OUT,
--        ------------------------- Receive Ports - CDR Ports ------------------------
--        RXCDRHOLD_IN                    =>      GT3_RXCDRHOLD_IN,
--        RXCDRLOCK_OUT                   =>      GT3_RXCDRLOCK_OUT,
--        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--        RXUSRCLK_IN                     =>      GT3_RXUSRCLK_IN,
--        RXUSRCLK2_IN                    =>      GT3_RXUSRCLK2_IN,
--        ------------------ Receive Ports - FPGA RX interface Ports -----------------
--        RXDATA_OUT                      =>      GT3_RXDATA_OUT,
--        --------------------------- Receive Ports - RX AFE -------------------------
--        GTXRXP_IN                       =>      GT3_GTXRXP_IN,
--        ------------------------ Receive Ports - RX AFE Ports ----------------------
--        GTXRXN_IN                       =>      GT3_GTXRXN_IN,
--        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--        RXBUFRESET_IN                   =>      GT3_RXBUFRESET_IN,
--        RXBUFSTATUS_OUT                 =>      GT3_RXBUFSTATUS_OUT,
--        --------------------- Receive Ports - RX Equalizer Ports -------------------
--        RXDFELPMRESET_IN                =>      GT3_RXDFELPMRESET_IN,
--        --------------------- Receive Ports - RX Equilizer Ports -------------------
--        RXLPMHFHOLD_IN                  =>      GT3_RXLPMHFHOLD_IN,
--        RXLPMLFHOLD_IN                  =>      GT3_RXLPMLFHOLD_IN,
--        ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
--        RXRATEDONE_OUT                  =>      GT3_RXRATEDONE_OUT,
--        --------------- Receive Ports - RX Fabric Output Control Ports -------------
--        RXOUTCLK_OUT                    =>      GT3_RXOUTCLK_OUT,
--        ------------- Receive Ports - RX Initialization and Reset Ports ------------
--        GTRXRESET_IN                    =>      GT3_GTRXRESET_IN,
--        RXPMARESET_IN                   =>      GT3_RXPMARESET_IN,
--        -------------- Receive Ports -RX Initialization and Reset Ports ------------
--        RXRESETDONE_OUT                 =>      GT3_RXRESETDONE_OUT,
--        ------------------------ TX Configurable Driver Ports ----------------------
--        TXPOSTCURSOR_IN                 =>      GT3_TXPOSTCURSOR_IN,
--        TXPRECURSOR_IN                  =>      GT3_TXPRECURSOR_IN,
--        --------------------- TX Initialization and Reset Ports --------------------
--        GTTXRESET_IN                    =>      GT3_GTTXRESET_IN,
--        TXUSERRDY_IN                    =>      GT3_TXUSERRDY_IN,
--        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--        TXUSRCLK_IN                     =>      GT3_TXUSRCLK_IN,
--        TXUSRCLK2_IN                    =>      GT3_TXUSRCLK2_IN,
--        --------------------- Transmit Ports - PCI Express Ports -------------------
--        TXRATE_IN                       =>      GT3_TXRATE_IN,
--        ---------------------- Transmit Ports - TX Buffer Ports --------------------
--        TXBUFSTATUS_OUT                 =>      GT3_TXBUFSTATUS_OUT,
--        --------------- Transmit Ports - TX Configurable Driver Ports --------------
--        TXDIFFCTRL_IN                   =>      GT3_TXDIFFCTRL_IN,
--        ------------------ Transmit Ports - TX Data Path interface -----------------
--        TXDATA_IN                       =>      GT3_TXDATA_IN,
--        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--        GTXTXN_OUT                      =>      GT3_GTXTXN_OUT,
--        GTXTXP_OUT                      =>      GT3_GTXTXP_OUT,
--        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--        TXOUTCLK_OUT                    =>      GT3_TXOUTCLK_OUT,
--        TXOUTCLKFABRIC_OUT              =>      GT3_TXOUTCLKFABRIC_OUT,
--        TXOUTCLKPCS_OUT                 =>      GT3_TXOUTCLKPCS_OUT,
--        TXRATEDONE_OUT                  =>      GT3_TXRATEDONE_OUT,
--        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--        TXPCSRESET_IN                   =>      GT3_TXPCSRESET_IN,
--        TXPMARESET_IN                   =>      GT3_TXPMARESET_IN,
--        TXRESETDONE_OUT                 =>      GT3_TXRESETDONE_OUT

--    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --_________________________GTXE2_COMMON____________________________________

    gtxe2_common_0_i : GTXE2_COMMON
    generic map
    (
            -- Simulation attributes
            SIM_RESET_SPEEDUP    => WRAPPER_SIM_GTRESET_SPEEDUP,
            SIM_QPLLREFCLK_SEL   => ("001"),
            SIM_VERSION          => SIM_VERSION,


       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                                =>     (x"0000040000001000"),
        COMMON_CFG                              =>     (x"00000000"),
        QPLL_CFG                                =>     (x"06801C1"),
        QPLL_CLKOUT_CFG                         =>     ("0000"),
        QPLL_COARSE_FREQ_OVRD                   =>     ("010000"),
        QPLL_COARSE_FREQ_OVRD_EN                =>     ('0'),
        QPLL_CP                                 =>     ("0000011111"),
        QPLL_CP_MONITOR_EN                      =>     ('0'),
        QPLL_DMONITOR_SEL                       =>     ('0'),
        QPLL_FBDIV                              =>     (QPLL_FBDIV_IN),
        QPLL_FBDIV_MONITOR_EN                   =>     ('0'),
        QPLL_FBDIV_RATIO                        =>     (QPLL_FBDIV_RATIO),
        QPLL_INIT_CFG                           =>     (x"000006"),
        QPLL_LOCK_CFG                           =>     (x"21E8"),
        QPLL_LPF                                =>     ("1111"),
        QPLL_REFCLK_DIV                         =>     (1)

        
    )
    port map
    (
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      tied_to_ground_vec_i(7 downto 0),
        DRPCLK                          =>      tied_to_ground_i,
        DRPDI                           =>      tied_to_ground_vec_i(15 downto 0),
        DRPDO                           =>      open,
        DRPEN                           =>      tied_to_ground_i,
        DRPRDY                          =>      open,
        DRPWE                           =>      tied_to_ground_i,
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GTGREFCLK                       =>      tied_to_ground_i,
        GTNORTHREFCLK0                  =>      tied_to_ground_i,
        GTNORTHREFCLK1                  =>      tied_to_ground_i,
        GTREFCLK0                       =>      GT0_GTREFCLK0_COMMON_IN,
        GTREFCLK1                       =>      tied_to_ground_i,
        GTSOUTHREFCLK0                  =>      tied_to_ground_i,
        GTSOUTHREFCLK1                  =>      tied_to_ground_i,
        ------------------------- Common Block -  QPLL Ports -----------------------
        QPLLDMONITOR                    =>      open,
        ----------------------- Common Block - Clocking Ports ----------------------
        QPLLOUTCLK                      =>      gt0_qplloutclk_i,
        QPLLOUTREFCLK                   =>      gt0_qplloutrefclk_i,
        REFCLKOUTMONITOR                =>      open,
        ------------------------- Common Block - QPLL Ports ------------------------
        QPLLFBCLKLOST                   =>      open,
        QPLLLOCK                        =>      GT0_QPLLLOCK_OUT,
        QPLLLOCKDETCLK                  =>      GT0_QPLLLOCKDETCLK_IN,
        QPLLLOCKEN                      =>      tied_to_vcc_i,
        QPLLOUTRESET                    =>      tied_to_ground_i,
        QPLLPD                          =>      tied_to_ground_i,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_OUT,
        QPLLREFCLKSEL                   =>      "001",
        QPLLRESET                       =>      GT0_QPLLRESET_IN,
        QPLLRSVD1                       =>      "0000000000000000",
        QPLLRSVD2                       =>      "11111",
        --------------------------------- QPLL Ports -------------------------------
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "00000",
        PMARSVD                         =>      "00000000",
        RCALENB                         =>      tied_to_vcc_i

    );


     
end RTL;
