

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nnA1LvIFtXuhnEgnrDveU5DQhO4oCdS4/TzHWVjuSWRiJTWamPLe1zKRcIJ3OgsD949QJsbaygaN
jpuk7BYNZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cfy8I58fHjYLB4BFaw/VxzidETwabyuF6c2nxAde+hbLnyzOfkymKdOr4Pk5oDTY4htTgTDRWzMe
dytGdfmZXjp6SJIGysindi/Logxabu2rWzFmbsNC3Q0gro5se9+3qoriCL3M82gnhvX/joJNLiXg
rsFmmSylhS6v32W24xg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gu3bZVKL/oo3WMbeK5OSi9dLiGmyQy2yONRw6Nst9yei3DenlP6wnhfHYdkStFXi/uvWUBEeZ7hN
0Bmqlib8vQ0eJP09mki40prhGAwrKuqYt+2JunlvLYMjlmKGJOXPgQJfoYTNzbZDTWMAPlUaZkK1
oZkHNa3Wtk5m49sk7N6rE0lY6V2L8UfgTL/MmCwu7DKHNfTBd2W2KricGJ6ICGb/eh21T7mo+KTw
su5JPh2xN6VOnDqK2JFdz2Fe2UsNNdpq35qIZsc5dRna+xfhp64zhbzGUq3oNeTCYYFL7/rkWyjk
xMfq+Y7aGpW1qrNdKLCLUa3C0oRubzA+yEUHPg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CjIoJO7bPG0vgefcLg3HndCtGBfDCnGBCSVZItM/kv6K6ZpvJnvEpEF/v7GEKszxgiutC8bTrPRk
/jMI//klbN/ln/AMlW7lDqpJ5wXp83c77tloVq04bnPwc3DaApr08oK3Bf1H6JgBuFfaRFUfxoRB
6anIIq6YC6xrV65+910=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D/ZhWxzQ+2vaiYn3/fV/u9o/WEb/ogG/V9KccsPCOCWeaD6JXzbX1wTvk2mHL3gwIIjopxpeK8ct
Dd/kho1WYC462ZEZ1ijvlrdcQ6jRucbVeVK20vWFMC1CO9YW54zFCdUIFDYoBjMQnJ6IU90guAMg
K2P3LVnqKNh7XA5585Xm34QBVEtkbFVGa/nBjX2k27AaOcjv8CeFc7ihUp4B6D6YzM34GhHkOxNj
NyMvVJlZ5HBA7JHakPw8PSgdpMIr12xEOrEcLpR4AR6H6hPW9blh2XXVPneGey+XXrhV6WAB7P2G
TGbniILS+ojY57htkmkMwgWfAakIRm5HfiYkdw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4720)
`protect data_block
EoHqzELBBpmP28QHq22L1uH7AxrqOdUrA2DkW1GxGM4evWp/w9SLFa8oPR8QfYruWAbP6vAn+P+I
kSbpUbSHZc2DRewLf2tNcMR39Fw/tArQOwGwQ/3Jj2dkEU68OP/TRw4CuZUffWh9W1sRDeXmxlRl
s14zB5Qeeeh4f0w7NLw346lLZ4JQdLXQQK4a22+U/Wevh49tGew57GGYnD0+MzIbaScRJevX+yFP
qltq7Plo00ijo9NkDA6nOi+ZrxSDFhFwYqA+ipuFaU4DUoNUxjrsRZbC6LmecCqsvixnSjDUHCk9
QHjyuWU+COjus4+y2jqeiUkpMyXVFOmJwHTN0UlDhoBnHuYFqC2PkK54yp7wzIMIPIeRWJZ4KP+7
P0IO3u9oJF6WA7G8gGf3j2iySjHAI7KT5yLDH1KaW0h8Fv5lHPVbIoGx81kiu1nDFFU+GkuT9Wgj
y0z6Os7nr0ugxj7xPvCaQwslsz1Akp4XLMafrDFmx6/K/d/UieE3W9pjVDb7AxRCihc4stu0kDPs
vkHzQvlbfquEI+WVIOAih/UZWfLZqYCuI37Syr4Ng1C1nhJaBFK33H7nEdQIeYkiV0xTuoXU+CE0
bo0IX9tk3jBg4OEqo2hl25SswpHvpPc8JWsfFaQHwPk7OIyNly5mLsXoEtruwY7zU+FBuds8wyFf
J7+BhifkUCuY8Kib859jPM3wjNRxHtz+Chh169CXSDo+ZKCBE4L7Gdjn7EDKzBQ4Im1iF5fTkjnp
mqy+A/C1NlR1VdKK3ALHwUDItmQ3XLhWctf0JekclHCkYwkF5fog+lOsksnO4Q+G1l7EDpk9dAJv
/eJhxekL1CU60/fGecorycF6bBYS4DTvDhVpdgXk9qGElLzd/Mx+sRfcCFCFprysWUH4X2CjLU4j
M0kQTrPFgCwK/JJUwgEx0u2pJvDJa6T/4u1+UXI3FKBI6uhaBbxswIWEV6ZMFG3KWvlFgubQUQol
CqnfOKKG3aY7Ux12zneTi69eEP/Yy1ZytEqIfgG7FcAYKXbjbFqG80W/aMY7K8O+iLsyX4wh8Lex
ANNIlDyV2oDxVxb5Bsk3Y/fRExCuD017BTFitLLX4qJlEo1aGssGP33gvl0FjbnRrhF08m5EycE9
aJe5FGFaJnCc61MIueJZt2Vqk1qLo0p+kgm9UeM+VZHmwA9UXlNEXoxrHrYW2D6+31DzPtBzzr4/
e9izeWiYyBMAgDwJnyAGhGeRVzmjHnCl3xndktjThKO5IPXugQ819lFuMvgLuaRYCWEaJcE7eJNN
7OnIwNevUQmfZ8jpWU+Tkyp/4x4WuPL+BupAE0FZOsh9XeyLT9mZA4yPuJwwf6TLZ5vTpO9eah1F
S45U2gW0WMp1Pwafi0r3OZVrxQ/LQbaU7GlQzFBOr81jo8Ka0q3mpGhNyWGX/5pTrBdR4VILIpIL
IytjJ5ylSYrW29oSFdU0vkOZnLv/d+L7FT+ZB7RBlHedius1vgEXRSqBaFGcUYU+ldEdPjRUQV5K
uod1pGDbgCtCPeOP+/ckK5hpqVnKPN4BGau20lQ7l9YXm8o7lAN+au+fE3f5oTD5HwAl832HrsNj
gkqLY73Hb31fq5b7LvHZ3lZq4ZaKsKqiLT+tkLJh7bR+AU5epkrsLy99XT0TwnB4PdCZnySeLk24
nIP0I3lOuPvrBrMKNZn+24EcJlcWZDAYZwhHosHDwTLchwNyCU+5DYG3mP/GLdTF11AL1Vn/51XN
dEc9+eZPbyQBGbb8JuWmhgSb+1Bkg36WgejpZda3WDCQhMwbUGoALSBlnTqs4me5f6On1yrPzLKI
rI+7E1MJlXJcaErGIKuJBxbVDzW08/5ROP3ChO0+0CDoj8G57WmsUhaZz1g8p+SX5+bYT1XQIYa5
gbaT8x0N3dn5IN4RHmO2UTSeU/bIU7CKce/btyzNY898vbA/u6LoS+9hrwI0QniG3x5cMFsDJIvM
3+lhYonBuKkY1n2nFRr32emc8eOvCrqFl4dvh2+jp5hhSU9keGKfNuSOXZfo0uaTMtnSlUQ+G+YW
lI7jcKQYaSPI5/htY5BeQSayA+S9OrsgTWTcWjasUdtLL9+pqhzpx5+OV+UjlParOBtZ/v/qtS9l
A7bAwvsaIVZOwiJu4/f7m51ktQSS1+fRUJflbgydVA3N6OUYQOLG1mKbnHaMbNfA0OCU8oCrXjec
UJdf5yrJdoIUolXPFGOU2xW+D0BfuKfkv86dv62DKXwBo+0YaBsCDmzkLKSFBwQSsWwrqB3em7Cv
4OOsKKNW3iGIwjN03mDVuvpDGCPKWrfXTCvwxDL3lcbX+JcmUnxht2F/8k7SXPkRcEL30B3zXp/N
8BEaPUP4bscQVafGeYstEoOcrXz8HxRKEibQBiiDTKOg+iloZhASVPnCH29s/uK4t/u0MzowtP/H
bXHdOchfi2rN64zc/3umeyU3y/g4tQnxehdHt3uzI+kraKmjnih3VNItVckbq3jokNndXINrEWR8
Lh3T5iMEvwIqdbrqkcZ+cv54pBKUpPfewteXfZLYR3uSlWNdMhkCMtoHu93DPMpq/YA1KZLek5zO
5qINJrguWMVKI93MA/77w9TNlPFWOlUau94zbFQQlQmfmzi9WhBfTSOerIfAKUjA4irJv5/IkX8c
s7R1BOYH45NC1cdbdN3rBUM+st8mp3iadmssXpBrMazgImLupZ4o07QcDo3cZzty902Ghgl56bq+
agBcW++ou5/7SIlse+TfdxMNgUIrgqF731JoL+2IffXJ5RMR5cRHgnPXAO2LI920DwR9nK31KPs/
hiVTrjiO9/YPxRRoF+gFGDwYxGO+XOWNCNLn9SvzCr014CskapAxvylE2QHVAlur2fPSS2P8CE/R
rGXaSA/ujYRrRq5RnQdkXVc5RdBrdRzPHBk1trE+d7/COv+m+i/klgI+Csbcc7EtOwZOd1VUpyMI
32I3s6K0iHsQok/txd5Sr5Myj2we2kskat9TqRyL5Hx6MsR+FxNGqlqr1JnEPqkhXEwLErnybe+V
3rkV7yv5xsYIEkzdvtAwRPUDTITg+cIpoad5C7b+eR68jTvnR6W3I6lpASPSVk4KQt5lluyrYCyG
o/YcAZy2wyFz51DrC4qBuC+XXdwOny9h832lUO1x6IcFXCKo9V6qPcy8Na6hDYo9w2vVALKnqAiu
nEarX7ETo5DFgDtomuraTbbKJwNpusnrIILigt55Hgy8tTTJj2vFQMiIjdelef7HOytz6ECN95xz
J/jh1qOEEpg1lnp6zbi4mZ05n6TdCsA7NLfXv4fD6VP69JMSf+tghz/AngPDJ5PJRJjem+KoD5Yv
RU6FyGCc7i+gHjOM3IixK+bJ5QCOA6+GSLDB4UADIM/qXYWprOi04e/D0nfPukMl9ylXNtaYGiVS
P7DgIM+oqlWb/1Cc7M3mJnAMlCkUz4PWfJ1y28r9DSjxdz8I09veNi7n+mRYrmvgznv0MbjbD7Me
ytXY3bjrbkoBg+Ult1tAN8n8quNtcXPlnIaUfMxKSiOObCkYMCl372pFFwwTJ8oJ03tuQpGRnXZA
VNdsczT/TYgTFBzTfnstHg+obS0ILneaRqmdDWdzzioxSY4d4SaKLf85HHGwe2crlK/WJlN0y4Gl
i0qrx97auqDMFJbXJuFs8k4VgCwMMxi5WMfey7Evu7cRkmPtwHuhyokgwlWIiBJ0KCvLtdI73arh
bJP9ybKSIXdr+SVam7VR09GNlFUCggUnjHirmmJOA75qmsdyGWOFMmf9OHc4uDYdZThs6o9pPivo
UHs+H5x6E8TNffxLRYyFUv6Kb33XpJsOzLJ0VGhuZzNCGvkWHzWLc6gsWy2pVS8bjB7QwggO0fVQ
cy5WS+5R0XmehK300YMirQ5rEeNFPrK5jQ7KgSuFS96ojTvtpC33L9fq4aJFnV4ouRX1fXu5HI0p
zHUY7mXAFNbD85F6G/DmLd6FC4zdn636DtKj+54KSQtasNbyAbMS56bURAnLmn/JhCsB9HvPDk1L
+RovBm5Ie3coVFwT3fAm8cRi5FR+Pb/8VipWWKJHrXIkcaxFrSU5YsSNNcCe3PaqC5r0VqGuo5l1
+IsDzBz/lfHjmRE7R8RxTAAGx7oH8fU/jBKRi6RCE8IdHh4ij3xnZOSoPB5c4HBFxh5tZXy1GmDj
ixERMK1r3Q6fa1bFSEmgZwrbhGzKxh9SO0egyT+C0TlH2GMDgWEkiLXSc9TMrJd+DLqLqt8GobGr
lubzRLbO2rrPvxzGa0V/3lRjs5EzYLt4LUVQiQSp+jilSSvTsEpXDRl4hKU+1+TIncAhFTrCgNFY
RO6/GmTC4sAwaaols91aZxjZcu3jo9rBOW9pUqlAparHNKWE1vulBwcJr2zzBZ/AoL5I5nv4Ndkr
P+rQ5CTKWXW47tJzm2SZW+IupCmEPx72fKo2PWRgYYcLO+lWKKS7IWNASI5Yxo0Zo7d1hof/pM8d
t7b4QvohPL8WrsOHwJHkIngvXdKz7rZ+g//lKaA6kK3S/ai5hi+cVeNGDol0ORcuvU7AgmwRQ0kd
duP7Tc6q8ZGZyt+Blb+B4AcXYTKKKbM/A0hG5FqXtyKv6Tz26ekM8Sf57er8t4M1mEhfQAUFUBng
CxucIFY1Mx7lg9rqqQNLzho0NNZBA+8iz1cy+zdu0lf72YRSHs7XNqmrrcC+68NVOdQpOr0SGtkQ
6V2XWCOp14GhTibqD4ae0Ui/sCPCYBp1g+1RCT06jDiB51c3P3lUMRBsb9ZhgOpcdnqGwlERecM/
npArDtCNYPUBorm8KmP4sgSbbn56jj6BQq8hse9wroGSvKtXro54d9qmnsYBKczvBZQxYXHuvutd
HlS5L7tcPqkXyq83WfFWjJmWhzawiPbVgdXkwu00PMdUw+z1qK72hpMeH6wUQsU+1ijbZRdUmWKy
OnFV09IHiVYKh9faBELD3vIA+QBdovXyXO92BJEbDGTXBP4IQBcHvVprqQ6DP6CnD4JD/2y9gkVa
LQ8eLI6n0zRhah/HWysnGN/sUqjhDEnCmKzyHV3seU9jcuI4lXRQmk6sLOk94tXt99wMDieTZjUA
jfmyaLX3W5r/uqbutzz12L/GHhMUE1wZSw3qdvdVWWhYMdEJpvapLXxFGZ+PF1X7ElkDR21H5cc2
myo71HYGU+7PYkXIwRYg1HhPIPOL9hpkZJfawPerVEuMGHC7iqr53WKvx3ZwV54mN0FoXcCWFPT0
P/LkCxKqwaoLt0sKERSmxoY+kKCeiWqQyLxVK3nKx/k6i7NcSeyoVknv3k4638XOmK7AadOtNQgA
dlrhN7zTH+8AZ5296vD3N/v0qU7lmhvW4GDBtV2ffwF9gkrMlSrBjciw8oM5UNNnslY2erIJ9jZY
AFHiWf+L57agrfX8+GAtIzM2IE6on5zLNhEBEv2D/8SI14ESFhe7yvILZ150sQygmmjYtntmUX0g
EbRflykewyFkS1jUgbnu9YC6/Hr7PHIzQ2folprrIbti3Ro7D+KK9kWShDiT1h6gi+f5zAnbnIOo
7hHHCx4WYs+bfoLoHS1zrIwm+AlVh2dKjGbITARoSLety4RD1A3FmVLWFb9vjW4gWpm8015HqR4z
qHiEaWdlm3DnbUp5MOelYrukUjkI5X3m5jAHI0idgKDaIRa3oBEFPWPhJtUMn999WIBqsiGHd0xY
cn/3DJoEfKM2AHGdu+FlaMatrFsZVMoWxl0/6uymgR/cfzXVAKov0NxVL5zod577IJ6TnDZ2dDDp
N6HFMRTqehD/Fc2mj4tmjk9a0Imj0f+AYWIWGa4+QUslw2D5mWdTmBexEByQvyHPfSLCD6aQX/Hm
2i4c9SsNaPffVgTFn2vecP9IAaaAdG+LehY59sdUQgHYbGumBp4SKoc8S3AMRiKQnIrISyPuWTHM
mKrhU1A6WVItFO8b9lL/7g8RMqPtrdzuQW758wqa/5IKDdjewZDPBgQp+HmIMI4IhEGdnsfkrYTc
d3QL/nJ7k31rtjxlP4Gi+JUCli9m+Mw24gVsNk+J19N4GYhLcF5jOVn85frWmVOWnjCa0CdYptcj
fb3Q8AjqFbkPFdnvnS1zcnz7+JlwoOQsc7cr8sDUWWmV2ZjMt+AGCD+3Vf4tYb/YO+PhIjv/FAt1
I9pmKl8Md9jsqJ+ThhsHQGyHogikdVkNqSREtWrcnvJYBz0LC0HpDtjAYaxCVCDS8vs3XWSjEZGG
32nTtstYCOpuTG0as23kzAHsLTXjSrNzz5tSIwAhdpSr6/i3sAPJVrrGOzRkFA==
`protect end_protected

