

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SPpb0sHtYr+7D0Z/NdHkBGKHFj6bPnAk4zCT9Qd9jSi/NZdzqHWXjKwgFh3NrYG/AQMVJcT4R9KU
T1kWm6bsuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PM0w38wqoKZTqxD5ZMv+He7u+x4mAKOhS9vNWqYsLtlMu2ni98hkp4Js0D7iFCQdcFCu3Jaj2Vqe
E0m1H+UGB6We+zPa+TnTKUC9+mxtEW7xpi8i+GVKfIfe89n3euEibIBIS0WLtZypuPRjuzr2TWw/
TpBFYS1oUTQ1qwWguI8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OIEbVz6QJBHT228fhImFLc7Q94gbSg/QOSgeKpAp1zRCxot1azeNL0EHN3pwZU9Qs6kuTNEAn7+w
agqdilWN9rl3uQlRBfW5KbIj2khza90rK/4UYrbcPGQyMxF8l/LBS9RaSzH8pqlJgQ4YfgwGNaq6
EHHkNL7CBEprP8VBO3A9geAIYBWstNirz3P/01jzH8PT87csZHkt/KV+1ancvBdl8zy3Pi5RrOtK
WdR5qLkbXJ6m4DjaubrW8HdK/fqusuCVkVGxmajuQw899iRpx5AiTEwKYKOor3msJGxdK7STL4ZT
S1m+Ec1GdsxDwYBgiKT0A3c1/unIYBS6y17V2A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y9qoE+tEhAFEsAZgxeFxNUflksEoY80RYly6rjz4X/QwncMYkOdY5w8AxmW4IYZfWprQfyfkxMrN
8JuXogLHC84iIPhEFIhJ/+RivFHW4gCUIf9NTOGEkQza7hd31B0/7LZttbZHcfTR5stmYGMhB9xi
VCriwe4C9iR9zFvOJxk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eCcOM7HngIZB2JCDRQ//SPPOptJbtDQ6WJM03A6xR3t8OhM7+MFavTdB4aR11UrppwUsYiZCHTBc
4AdaSSNbTEcILhRaZMNZ85hgqiNgFb3YTJu8ZIWifM+Ad5U1zkzbH1xsVssRl/Sl+cf+TCDh9Psd
UOpjIzWfsyGgyfaSSbczC/DMklBqFcyspqzOP0YGdgI4It3e5xnwDvYeewRqIZggj0RyjkJH8PxJ
o1XlyTZFQZIIFN0x8sDbcPdsUekU3pOCvI9JK89jigNzKmLJRotLEgZQt0B8gMiz/gm5u0+k01OA
f/7Xo9TSexSaZ5evmswsNTBQhg4v8j39bgkh9Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7744)
`protect data_block
lqgIF1V9xnux2eUcAFOCjz1QTEmk+d8Z92QM/ZPJXkL7aKnSI8gWOsFBxlzxvWusrM7Ge+txARMk
UfpTQK7aP8V9iL/PPWxmnohj0hZhL5GW6XUYHNJ0HHkocYoRI5QQDYt3CnJNfgiJhBWdXP9kczHf
3Y7mSPxjyRtPuzjIRsYcgSszddNcduwiXy77a+/94SyZM9WDKM3OSzkxU1atjzrGIVQTfsJjNOVE
vLeXNR9s0yHbxP3538hqIaWqQB7X78c5ZAdOvAlRaMdmmd4vegf2XWHA7hzjf1xKTAhXza+azhRH
pMvnX0K7zHdD4a7CEh4WFcduUCZG4LI7mmvRmzS5a+bWo50MW+IpGExllIa5tGbpgsQCWNzbBAuV
M+UfuwsOlCHc6kJK6yqhwoFgbJnLQmd+ombyzH/QBn9/0qDcJlbxNjjairi6S7+dn50X7OnzUuXs
tkySTr4uBbYqzBeIAqhDuMKQXgzrOXIO5l0r7UOT/4rrPgsHtz0R11tDCxB4paxS5VLmM/169P0f
iBvEY/1QKxdBJ/QcpfJAng2GTCqGuDZqRhtC+jOAZ+NIgxAwFob20pLBa2DnEdMQAmO6mSy9OI6E
aXQ6jB0K7phWNtHBB6KV9sk9yqzPr2KV4HPnV988DNc4dRfsM0Rc2MhF4MJGdPvwzVaoS6WJtYCF
jWXHiu9pRCdxtDUXn5oimPKE58junJQHMp+5MEEMqVGzHUVXm3JGXFTYHbLpLqY1Aji1mXw5+YI9
ZBkzLhZe0NoRr9HW8+r9yCYOMDkIHpVWmYBizQWkXbtbwSqlWZZDvHBR8cic40QlHWleY35e4nPy
IX28xIA9JxWnFai7V5/x0z+D0XPlK2VR0WjR92UWSNeWVDPFgKn6Xscq8zgh7mxD0zWRdlglUd8U
hrNOPV1IBwphwd9nYHtf/SB7F18GYpbYF99QsTYtAWlP0bBD8CEP7poc3VWd0tzmFGQg2JrxinWU
61YI5PwoxpdU7lEJ5ef7qQxuWzzZSIX2EH0Ju2PwLJEwtNOJuvuiyitTBxrdV6T1ilsPZWQqpoK/
pO/go2EGb4H0hTluTN9hUYv5CBgyPdJ3bMSHsm4sK8Gc/lOr2+kC6wyaUszmE2y+ELi025h+HHko
yPEHutDo1tnWU9pDPYNER1JQ33BMIx5+yKz6iIJgfVWr+7KesUnus7pSyahrcTwsCBXy++epLkt6
eKe27Om7NUVVSgBfR1MLSngL40ynLOymxV6nPNzXG/g92IRBuTwdREWQ6jYJA+VJY8i19FG/P8TJ
PvxRnA1DuTVjCneI4Ly3pRMJmKwjrS81hGJAA0UnBR7yiqA6UHdJNkqkNOtzyMGYRnI0y7PdHLuV
iEdjz729IcYJqf2FjgV9zdAWnNHqPX24Y53T77CaW33hPn0ZhAR/zsD7zXzB+9wOXfLe4LMeOw9r
UjqmqkLiWY4C036Zpb2EhrOYgQWsooiuHXf75M3nTGNQBQR/X0xqpC3sVWWPVk5sJMQuFPko4XY0
W8qc4Mk0koLPi7v8eBxxQBCnRx+o+5qVvdaDfRZ8XHY43P0/ptwAsBONR6f4NELerpBbs3Anh40E
w9J3BDAwzH+NMMNHP0Ih2NjNgI9IX1Hg5X/7PjebPlVxqBcfP4MM7fmc+RSJTSP6cWtGoN99eAy7
e9xuIdwDC4azO1Zfx5He3UNnvFEreqVYJExc6SWxFu73mqYfSdfCqZQfB8H6e4N1yi+hzSj51tI9
Fhk3zZmoVA4ejMqDe34WljEHHDYGSl0cPMXc9cXgWGlbKwFbANK29JKrKUYw9frOVndSry11hmpQ
nMrSMuouhUXz/YI7/LYoHnxRwpi6ap7rmRmook1/xXTqoYUSjzgOptnfz2A078HWPLn8FCjmq6mw
V8lEslPJ+r6OcYHMv7W4qb8SNL6GKwqwJq44DBdgdbvL414JWbUMROZNSYV8QpHzm9x4NfZfgXZ7
ZScgAiyVx43gcm5g5Wus/bZ7Z/9FVDbNdnBjb6eazBnWht5EBCjJILEQDxMK+LklM3qiZ9e4dGBT
LBbFMxyQeFaaBuSNGFUJlFIrHahYg2e1cdgncgqBk7EqQd3ln8mf4jspnTODguxKY9jRXOkhM5nF
BOLh8rv31sPhGpfGsUIxWlAZpTgZzLPsM/7dE15pRAWymcVs3brkxhltUJnqSnaroytBX5D/xmzJ
9pN70HrEE2QPqCp51K1UPVOBe/sbESRZwAiN0lF7f/3I2NIbczbXrbs9grHjC+cCTs9eNEK5gDXf
O02azPpJ2spnqwmok2bQR3pzO4KL4N3NJ1PL5OZuIyLAC3Ti5kdgU5WhFP+KzfMScSWg94dn3TIK
5v/tlhpZCYCQ05P2HFMkiJKaYC3gN1x61PGahpAJWptysyrKlJ+qvzxBNl4CpAlSLZXHIEaKWfqU
mcLhH7a37zvkyyCN0KIXB1RJgdVRZVT78N0kGyP4zzYB31W76Wqac3YtksaSynSbraxadOMAxmZv
LFaxcZxlZnU8YRQySrtapLqUI6xIK++rYhR+4Gm9Dk31C4vu07oTnZd9yurXCujdaAwmn9dISMht
oFH1pI+XPAAo2Y1m4U1sjZGmGM+NCjPzpcFtDKu9dwZKlRt3kgKiPhAaiv7KSkqRpHW/iK+iIK0u
9DBnadpawXZ5uvKAUFCAsU5GFYtmAZMJZCGhDvyZo0hXrI5ndDpnwicOKLrMM/6nnArwNpeBdl/m
TLGEOe/pNqjlWBCNRpTN5JYKbUqe9g8nF/Z5OhgnSnNNLRShLLfz3+ILitGYrD9AzWrml705iMvZ
aGYO3XziM9uXTt2kGfJrkYZ53yL17xhoSgjg8cnt/4+AnsoB37iBI2DxmeKkCm8ceAzTexIfvWd+
MuG3lC1nL5I9AO6M7QLPY+RNFYCLF72yhWo6ZHvqKOT3ZleixqtYo9bgbWPJAObxqgdMEN2TNUEm
a1GVI6qcx56oduPA4N2DNmO99C4XUwdGDOntuETbnMdBXLrtJEIbhSOzOOvgUx1xpXJ2J1FDCiib
PY1We1Dw642nVfkVEdhvBcxXVE2VbueJ2S9wTP1XTAnQPADTAACyEN6tKEah+JatsdenU6zRTiIH
04dL3O2jy4G8smgjDwI16Pk9fxCRsH5amPY+GTK4c9/+lNcodn+mgzl992jTddvxSS0/lW/YZaPb
AcsJVRt00AfM1A9/jhoHRaVPV3zKFEzOostk4Y0aMttZszzAXUIpC3EkZEn4SAclboqNCk73hl8t
DUYK7FYGurruv/34RJVpb5PhPp8/cucZlGjBFQtdrq9OBGiyDQKTRwu8pIs4JlewRBzaWecVpyb/
ADDUao07MAEy5IysN/BA2vlU6Emhj5R53oCgs9Mrr2/2yUsixULOl4oj3eAyYQIt+dNdS5Fy3FWO
zeSf6dfHiwjU4jThKxQsHH7cZXC4gv8Sb5yLzr0g0KtbYecTTn0oaaNQNsLFwivppzMDL6gMsP54
OPAbo3E+RoTvBdm89qkfCpCk7eonD8LAAcfhYjdGm9v0pDjxl6NLMV6xMu5tNHsmjZdXgwLxTy/F
HZmYbztKjyaxdVUf3bLjIv5rpcJhYONlOPKDc1l5yaCoCOj/l0fNdkEDTY/LWdnDjUaKLk67s7bb
Nx3Apfgu4uZy7/lyrN3Lo9RyfLYXfnt1V2qK1qeVMiHh6G69aKBE7evA+KY4ZdznrxFbpuzYX0aC
cIwB2EH3pePgLkR9SXsqvT3QHkE+7PJzMbmfutStvwiX1bbql+NubW7eq/kcHK6WYkw5ejTDor/v
03Ub14lw9MIlLDP1vVktPpiARub/y+l2zEe5DdXv2GpluQYACvOcC79LaVMtYnlzZMKfEpESKc2n
aPDFr7Fzc0qA1sWBbVweZPeyPa3ZThgrGBsUOJw6DcvZX7movtk5GYA7Xo0uiBGE5IKx5FyjObm6
Vs/xEqegPRqD69/qNTjUCsJFV8T94AeREwCAh4eZJZv84HddFVRyjJ2hMnDB15DsTxezLy6rZmKZ
rT9u0hjB7cj0zqpWjp1F5t1LyihFBDBNFTHtpITBQma3wQm/1b2KtTlPU89aWsw02UCtMWJRy+Fh
we/9o4gXTkw4/HOByfyyXf1hq1Wld2fFvEed6a93oYoQ4HOh7Uso6636OgBi4KipfWNXJoKGJrs9
WEZ6ZcylTfKRiiqwN6hwg/qiIthweiwz2Ap4LfSep4bbORrm26kau4KFEOz7JRv1XN2UyRy558V7
eWVeFye5pYAEFb1FmcksDMVmPakO8uTt1exGRx9ReC9ONXaZevbi5/NP9mEBnaQxIZU8TtXd72eA
BMfU6m9Kmen/cwDJezHmUDMbrrtVfPl7ntvH++4K6BL6B68kpE+7zt10tov4slZl8v3qQuH8UkcA
CQN1JnE3D/CRNlxSeADJMU/mwIP6IKelXJ2i56qLrF/5EMOxzenG+CmQ8vHi3pBv33Zy9r0kIgEE
VDsTezdT4Sm9fQzUwgPN+W1ATILgs+qNiP4yWX/kruSzIrpyWmOURBk4d9YDv1Clhr9JlZjdoPvL
LkTNkw7hbCMkbbiXKyb477CPlc39Yiz6J8V+k773gis0fR7y8x3NEpOGsl9rMab6YSOMGZwrZgNC
MIydL4lmAnrK2GvQRs9kB+B4proYOMvZE7rHrIcoS7Jgm8PQxNYUe5DJZEC+vo7fKk+0NjDEWof0
srz/YkIxsYNqteERDUJxLA/3yuJtYPT192d9kEv/MuWrf02n3OCdLJKAcnaduTNkGXuoxBpHpUQQ
X9lbiSRbAwNUKZVNF5gRgsvBHUIkhqqJWU/9sojZ0AgsWuhta1K1J/DbEiXV1f08AVKF1YetjaP2
mbLdIInQv6Bjcf3Ab6Wa4PlhYaSbPwym62B9BWifG0XPl1+tkcw9OfvKqrBBC1GLu0zdnXOkA4De
mi1LIJ1lm5Ra9zui7lmQDiwRYIPwy4b1agc93MVkAJ+dYOAdiiu0batcFgg94Lspl3WQLukYnaAa
gM5W/IOMq6TipRKUEub1kcA4J/0ezL57BNaBGqNdHBVXA2knzJZd2r4akaVPyp7yx+XTlMN8ksER
PNn7cNEJ68lfIj4Ur2UNabQW3R48MC2EvbVpUfLQmTybi2tGIu408yQ383LmXEIQJwVmV0QSb4zK
1HLTfifYNBP/ZPiCwLXCjEblSNe8TmJKUWThhmk/Ua/89pkS4UgDr7n3tpn+un8WRtyeWCAsetEJ
2dXdcTqfVZuAEVNsiGEiCFD/lcEz0Q0OyD0fUilDuTxgRoB6QAgFXr3ppI2+Mw+HSwGt36vt1+NF
/uMp2oh4sB1pbCKtx/TfTEJZFuDy0zVGz7VSsXYP74wdUzgcpb/nV6QGf5fKUKefAkuBpWJPBatj
5sHWGpRPUHbRhoONsYCazIPX/s9dy9oCN3Er5XwoIj/dn/FjyAJIX+7I+VXvE13oVJQyxLOujW+b
zajbMgqEDFJENS9dBasc7S/T0bkoCpHdjX7FX7yaFMnFMxsAaKfQsgspWidyDiAxWI1Zod0/tdEf
0FGNlYiOYi3fUrAPrGScDFBcu3zozRpl7n3HO8Y8A3esMwKjOi3Y4ZD4Qfq5zn4ATT5LCtMCHD8b
OHcYzibL+YMe6yAgLmBmYMyGWK4n/Qq/Y6TMjtgIiFW2HCfqIXz3l5ExOCiczZlxZfo17mkZ3jEY
/oEuftvaFaHt5ZwvgZwcOrqB8tAcXfoPqqCJuVJrSU8cQnzletd5TgTxmsbQYroHmttglhbPsz6m
jNKcPaK042BGIQWyH8JKg5+cm3oS2bPSXh5Mvq2ZLHr5rjXxmzzznTecMdUMYaU1OdxUPGkFjbI7
P++PDYPbXPIWebid2LVtdH22OBSgULbPxUe6Hmi6vz7++oLU5US4z56d5Nd71Dsk1lyjLGeA38cu
bzgWYXPisGmmnyXNXHbeT5vWMeXmxvsf+MEaK6ibFQuIHXDRv4wchqjgH+SY8Y0WlXoblswaqL1Q
xH+ROZIW0z6HNYm2L1Ng/gfrv295m2KhNap0555aFgvLhOFUb12FdZsGjmZYySB8t2z2FvS5L2pT
P0+WapgBRQ0+3f2h4GQHNuKYJa9+1UXuiqVKlOO6P0rBjVBlaLM/vXtlAXNCoDX/e6MSPKPX4ST2
2Ti0PUBS/o23tZBnhqgsjNuRa24LeD0qgarkB1Xm0FMAQHJJ7qoqCGyOhem6S+nwjLD2vAMnOwNi
azzrKHSsIaIDM2pQ/Apy2Eqe0thEkSBTjaa2HkbcQLXqq7tjqizULoH2k16YaILCKVUGm80noP5j
RzhyXKIJWFibKlit0vj1wzKlvAr8z4xH0K0dBKZg9mVVJuZUVxBMzecvzHtpZ4/+QAV0ImtVoB0O
LODfp4NKH1SzkHR/WK1HOFLaHJSsk3FTbBFtouvNH1l/Pn4y8z7CnwnpOIojbOC3XfxesLLoA/X1
JI4dTQSuL2oWDHF6d0iKqtH9TkCOYSBiNvERSpvNH8ZKwHFOw0Uzj5jkMID+JnqW2h1rdop9BhxZ
ksByrp6kYANcJHxUjKF5yDqWWH0tcKUL7DpfTXIHe6piJbYf2L8aStzpZi6Pn14YGE4gaIQTUtjL
5tgcw0mZBTV5wfe86c8ptSy4UbLbijnyAdV5yn8haD5d7j7iFyniJQ49zshWhOD3JB11dV9nTvVI
G413a1FjMtovXYjE1wMOrOIEzr9KIENOk+NnTAHb8+JeWbs8S6e7Dbb+nBoQJL5IWiIPNjBym3Yw
8v7UPZqLNw56BeT6saKEgdC77LgKDpM4AhHLMyxmu84WzgptcXgDH71ICk58e1lbSJFxFQiUKhem
K5MlI9E41r+nbuv2mw/BfeV8d9xBd7rCP/6qRTdstlvGRKDMYRK2wrYngyuZh/kYqqiJ30vLR2oh
dpPVE4Azh2Un9c1UfrsN2gNZLre5s+hyM+RqU8GCtaMSXr8lxx13XNguI8PCmSeaVTbLcgTL1eqz
ltpFt2o0UP9/hehtDBtzQlIUZ+tA0oCwabkN89vywQVOsNPSGKRsWEoFARIoVcH0fed/9Et+tRZf
Udw569M2mrWJ86UHJRifsytdedXcNHY/X0S44RxwLDFlLFVWjh8ewOJgEcy2wa//5M11AA1lWSYO
LbE7eYUIk8FAntxyKg2aK2QUxccOOD1zMzomVd5SBmq/bswFdoE18emC2VeIUoX3Fnnk/f+rNGog
wKrC4QpnJyjgd97Q4J6iaHR1jZxHS1CEizcvANkMQct7hzf8Xxh+EbLi+cDwq48EGtN7FLSLr2rk
W9MUcgFK1pmgnOddohg7GrTWBE0eT79KNsH14EbSR30mVrJV0+LoMUFH6fKz9va/m7RkdAAuEHNS
nGFwgjpScz8zXHAY+pj2Gabn8CFnxGw4wr7NnHVnMbfpRHW2ECVtvG2I/Tjis3now3vDAA5KYi6B
FBTQ8nC85363lRpn1pJkMg/rGHUOYRbUhOpdbQ+MSTjzygmmuww2Huds6GHlPtFfbIeWx0wbpWAm
G6nKDrDFtW/lAtHvQGhZc9mjneSbZVU0sxbji7Qr1p/M+pEMS0sxV1KehqXnQ40eR4DMoLDvz4Gi
V2CrDNlkPM5SFOgCAztjpZSVXZiW9jvjSzQjYe1eRc06FPsy5Yaj1Jtfe/NJ3c3X1egcjwulwWwG
43K53nHVQjaJoOEQ0QW8XtGQUsKe03jiH5H+Qtt04/z++q1wv5wWjkToBPkSgDc7pVds9glpEIGt
QiRu5NjwI4eaYTvm4DsLwn1rZGXMr+x7/F8jz2kBmiAUL8kzcIz76rIE9Y5X6zcTqB8dO3kOv9p1
KhSC6tZ0H6iNml4FijUeJnERCQ4TLxYQjyxMTy6Yu74QRxWMfE1jXhbvFhAqqeyc7AxisqhfLYAo
M39CepuqIMm/yFuSWzS9PCIQYWYDJtBIInmlmjtH2A/fsdLOCWDhvVWS6ikcSo6nIigioZ0/cvuL
jj6aoGlEtYMsLtpBmY09b1ihH5AFQ8L6/ptStfBuKuttkiEC6zPClNaAHJyYgfwhmtUybgRh3M6t
/WHBudw1q8ELITwL+6FZSx9tB1M6AWuxZVOjiyfP5mBjnoaBcAkfKG4F3cOY++3nG+5ldxD1vrwz
MSmRoILNzeN8C86IvBDzvsk7o1kX46QTLVnrlOmAS5czKF8weKAFNH8ZOFQMGihf1X61zdFXTm9I
P4PmpYOFmy+avlLyesY1YiSBf6MUk17yBOBvnM7mygFyE/F3Ct/O9c5q1pZU1zGnfa7GoGgYk2Qe
IPnvxUk54P+2r+TBBYelXaKk+CyaeETts2QbaCsNmCzaFq0uIVuO52L7RQf4xn1CVpuhxbiu0N3M
m5qMV15r0D40heujIg75BmSNnoCpu3hvBn/D6Xb8ZZXDWdyqTSOqruRe03bk1UEpAkkuFJip8Sjb
wIu9JNZs918KmlG9amWTPpxF8l8KblVPX+6bx+p45FeFvzHOr4Z95BnR12EkrR+AmYOWEZG7zilq
ctY5Z6JHPr1g8eVhxRea9Fy2O9lkqp/9WVgRoxAYSenXtkqaFa2xi74kBwhx6aK4kKJg8zK8dLO5
5WRjJDZiPadn8Fm5ExQVe/wcmhIQSqbfs7btF+LGVX+ZuErOX80ucmi/+k/Rk/WORMFzfjUB4Ri8
84R0TDCoAkLfpOrfmwBwuXDytY0jWIwVohSKceqMYsSlgpVTRAxFgXt36GpDGc/JKsrFZ5KbD7I1
PlcuHPQLbF6q4hkAe6eIEU2M5KjB7D5jcQwDmraPB1GvZWqfv68UeUB0RXO4N45aXXGpXGmBoptb
aoYeuLUv3SjOaLfZuxoq/NdezSBh2XXq+i7k90N8U0y06ER3Ep+uNTJ4VzgrlZ/9Y7q2mX+JtVrz
sVNoC1H3AXaURGO3k5t5JUTUMEfGstfAUWjs0tYeU36q4U1BbnDnJx01OC0wkY/CxYhYZWmaU51z
rwXP+pYyNNF8JXeAP3vDO54B1eGwJ8GGx9ESsHNp+0X4RiI5rHa3hyeurwBW0L4pRt8QPobeZUc0
on8idKx4emxwVV9MdEPpiJ0wZwilRZCd2LyGDNVxmspMM+Avv27y6MlmhTseCPuHwN3Q6Nv8080h
xBHtv+qLX+t1Lz2Du+WRXzitZkWWym8slfQAOt7UO2aR8CM0ohhkRjTNy7G+6h5yPRPrPImTSKQD
ERx/boapvSAv/JvdIKlsGTbLJw7ig55+HhJ/c3Vy/gJzqgXVcs/H+wc8vx+os42xRIlH3bJ6+Fu5
6+jYTDfuH49Clo4VSHoawDVKVlev3tMS0+mGSF1l0cqzyGgXmQxz6yI1CFQ5JjjKmOWeqQZ6LaNN
wYOkh+d+IfYGh05gvZKIPKjwHbGNjyD4PMlrvqMpmU+LB7BclxROGx9iaSXKpoW/M6bKGGyQYF9E
iLZvpNnjT0KjoocLPe14liKbBlnzHECZ+0P1OZ/6rhpM9LKM9SRpZZiTJIDYse+yQ5xMGGXaJjuC
DnAB5UY/+zz4q3Z0UT2bvpvW606JBhW25uj7kY/HtPJNu61GllCTmYQ8JkinkqipKTSsS5NtXQgs
3Jb2bM1tp0U0SzLr47qKYEYqxXu60ayYyAPLACw8uUHFhPVgkKrVFKO9/GjIXKZejwCOxmjhI1Te
jK3DneiNbFrjgkq/n4YPC5SxDJv77LqSBDGmj0c15XpFN3Xi3TbmOxpW+GfZKfWt+NlEi744pVtD
N8SzQQKnK1VEGBVoP2I2NBnDpq/4BKavbR6ucH5vusZSxhngwoTIHGZoJY6kNWZiFZhja3ToYJ6d
SAWcsjhuOVgvBLMvVLS0ruKeGt4lBV3dnhk6+gBS82He2jy4lm2jmyPB97WlcJO/ikiOw3QAmG60
KMW/s4EWW3I+1h1nK/yKDXsDzhWGCvhKHq9izZWwUwxDSOT0P0CNKqSC8RV2tPRUitl38praiIR7
YgVnHxdI9p5DRkPBKDBiy+aOUavZsNMQUlpd8lylXxnBS1NBXpnYjOsdhd6Z2WvyTOcjoqQbrfTg
J3XFY52BJbVEumRKSlvxQFS/88hbq3AGEruX40kUUuKm26SkEQnLUM4KTTzTXck4qT/TrngZWWUx
0jbJPpfk0WsrGjWjo+lcgnE3QiKjAg/ZRFfLs0JkNA3PEdKfAEHAxySg2rK9xbFhOru+Xi39qTtP
uCRooNhpF+xw6V9gsFDBRxv4j2UjJ/3bw3hprgjxANYf50CefWw5E6nMTXArZiCajSr1dqN6JZd9
w8A6D1RqMa6xn01BBciktAIBFzSfAu4/bYkrWkq4Vn6Ka+ShZ9PFWQiXe3KaC6Shtw==
`protect end_protected

