

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jtXjITQ50a0ecf2Im0hc5gDMz+eLQYg/zzqRdEOtUonTsMauUR2I/zDZca/cFZRkz2Bn/e1TcNfn
wKr/p3+6Ew==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ANnTEQ5JJem4BDOpiZXGW1BGnlByArgufttfMLkwemXR407wjOM5c7+DduQ2B6Rws3h4VtvHo6rO
wrBVcL7VsvPq1+tV939t3BGzv7HmeOgz+bF6BolXyM301AxlRkWo/0oJhXt9sAWYr7zYDeoXtQZb
l76HOHad93vrCilEPkc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XmwNj23lI8XFGQYG7vF9oV5Kxca20ebqjV8UOZJpCCCr+xVAS7ag+llpfkHEOHuw9tSDfsd4Eagb
WTNoLsXhoBdOAYPEcNzU+W9qGu9/wjx0qrsJ9f6NyxsR8o/IzcMAojV3xWACKEn/35hhcf9UXdPw
jFtFMZBq82H3pspBY7rQB54QzJyh7kwXdtgWfJuR8vKgpz2Bgw+sWz2/D2DHqFf2M9nR9Jj5wsYi
jA2guHzbYFRqb3Hyb8w16e2ODRs1Chv6CQa8J/8jZZjpfNE9JYFfYFbj02jB3GIgpxkUh95YsKVS
nyG+AAIy66AvGO8wjxEaZssb0O8bFU7NUeHAaw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jhiEXYtW8X8urAKsC5DlhfR1BlhyMUwpr7b+LLkcXXJrwnqMhkaTCeeV/MLdD2fZlxbKcfLK7F9V
JGPVeMHqW/OgkDKoPYInFHgV4dQ8+vVlaEgOkFd21VNxhDMogpMeEu/OUw7EcrJ+uVFRL9Y4CZQe
7QVrICfnVX7/1Uf6PJs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fOUx+hBZ6Yu+THnpJi++K5FNQDW/3h2F0eesEGevzvwYAUzmUKIlynhcf5gdgPU7azk/daFeo+yk
Krq/01NBV0vQpvK8q0FHFH+ghuL05juk1koa24QZKqKLJESEoqe8+SMhcjfeA/1/cXTmsbZU0sOR
598davhiRIPeODK4SAJwb2vC+fldvr29ZQPfn7IqVQ1mWsnCoHzWBSYPyy4Xw+6asrFDW88G8kf8
wyRSd13FqmDW+hKwsLgtlOhvBagW21tHVBbEEW2kPEAMrlmNhaLMf5utkD/lTPuEPBItEC5xgDps
hn/cW4ZYOpIgB7hTnFioHxnAEnyoEZ+mfU5gPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23952)
`protect data_block
vd0xuXKupDyEHS7jedzu8iozMisjlpqBRH0MZFSpOw6KGOt4E3b85tjUsCWiv7cHtGmzSzDjc3LK
eT6OABdht1FxEeYrUSB3HC1fBDH2LnDElal1fShiFXbFAUSdIPoYuAcTY8BlhC8GY+Ojm9BKUbPk
xkhi3/yz8ORUuxt53ytCla3Ti91IkfLAV9SbTZ9d/o1RMUC0g/bhvBzobUYAK2ZfneKs5OUnbc8C
st9l9FMcHqjBkWpIELOXLn8DMESb7x4nIj4MuDZVyi5xhMjEVYwUvFE92XzZ5gRS/OlPIUOXpStf
0qelDiHOhof3eN8kJ2CxmoxjFdZyg4n1R7jccB8dMhDmEYlYzh6cdPLvtR30wvjwzbrd5DNMFG5K
ATIebK+7RtaiYv02CqEu3Q7StAKfDVYrAGRfAnA/RZZ/320Fw91nRd41O3m9FZ5qoLurvedf2Rr1
IRdITPl0QIDipRsLVGr0bfpKK6bY0Hv6AMmPuqc+9KzZjLm/F4kFk0YgGvOwe5/mPQEm29ky9Ps6
/qn8LoIaWV7bcLwcsNuezbgpKgyQXQs7qqZCd3zTp2hAk8T3aui7W3NCp/m5FsYkhT9+5JUOYjQ0
kc9shQz1h5ddFtMwwfLINHTeeAZZb6AWL1yMPP5k+8lXsU/q25KcTvW1h+DWk+83SDYSRbH8mmHr
8ji21CWffaRcJ2TWbmGuuYvs3cEmeHaaoYFe0lvCy4xbx0MVsktYFGUhvB+tcEA3f6tOjt/y0Sn5
W45heSVFZzuy1/EBQvXKyoEZhseEJFNDl+zRhmGjr36qMPYl1RePhk4Jk0L3ERr29SkEUPxQzc9U
73Fz+pX04ShcJSPcnTCcnf7l9O5+BmTS7vE+QIuBYIqbSXOgOxXidQEh6X9A+AQjITst0QJqQeGY
ryAa7QXl4p6VAmbRTeq0ODDMFv/bZ+4DtL1wlwwK6ZP6aGqhYcEr05orcm9lNV/+p+/cby++KWte
QuNdKIdCjXhgpNfsPQR1tY1jn7kab5IJXt15kfpFnT0ZJezdnQl0yTqyamwG0AO8uO8qriv6kOGg
MKdgq2iw4p/dPvt+BcbpT5L8J3AG0NlGWq3x8Z8lqIpIG8KjXkj5e2s4cFkZWlvl4f1MDZvD85wz
jz6cxlhoMxwjvkg2usSsQptPIBr35mPJrNkrEhw6aMU5sqqQg4f7ZA5+SnAgakSNbTHnPvjRw+C+
LRVzUcXgNxwV54H23UNc7GU1hjcPblHxhnr4elM6HBEor1PQEBHD9JfYw0x+vDHfjpxnXnKk189j
Kmdnftuoy1O9sE1qkKeJceevxnKIIRIHqcitcbW3mIAJRRcfBG/4nyKcxdpreed14QP8DntITpk1
Sv3pOmvaACzscA48M5X/CX8nikAPFyDAyVSPfEjptkFO4YMGOwb4pc/6t1Y2HnA/hTxUMSQIBImZ
6nnTClOH0DIO5AFW3hJSm9JR/QFhu2kHbRTybNVxtI8TJuSduBB70db8y3kjQ8YJ967mzF/RyVkf
vhRm8dZbXEGQ/USnWZILM6OaK25FOpWRL3BdJI6PhGnnoK0EULjYj8kAoqqAKbCg9OdDXqgHBWf+
cLGAUnpAayCP0w3MIvT9hv9W2ntQuMBPPIlQXbCkweP8MQuhsDnSi/n/9S2MOG2kaSuiHYhl75bi
feI56VgvpDTLTry1HGg9APIbFa3VF7RKY2DD/MVA1r96qfbrRt1KbNZ+cBk93loarla7LLKqn2M4
mSffmTtxxv1z86Lzj2QuFO8X3aQg1v4BHYKkBSyVG2JCcfDtVhThsewNcNnJKTV6+2MKOq7/D00D
0wHV9rwYsBd9LjPmz0gfRL8R9NUUTAIXU9geAyHWrjtiAzvUIhBjnUnL2lEDoKfAEAa+M046Y8J1
fSgmZnBlBjKB/8iRMyEpkKo1xSQQSruMfB8L3AHkATUpr4nA8e4ttbq2lrU8iAvwZrI/B55YiVqT
mp/y4Wnbt/6/vRMduxZ2Sge0UOtInqxXW1qDly0u5vdSuwFFuqkWcfvUTOpjjGUfvedjHZxSAFgu
lcK/8deJmeiwTk4FkFvdGsXPnmwbVooMazNxBUQORCFGUkUAuC2puBRXb/7hxSMVmRy6obVAx2G4
avdWp/vKQQNoWDgi2ULDE2zS43FHNmO1wqLFiYjfbpWaALDUfwLXOlhhw8SzFhKBw7UzYtP8ZBl6
vo+arTgYb0M3PhQZKDwXs/cXslKcCF2QfUM7zfXYAE4HAx7Jz1gUevOz6GlzR6Jlzt2qXlGIWr64
gXM3NP4uW8EslJw4Jiiw0YEPxyGlaJuxqvz1fJ3jl8wotft1ZuoA0nUHQBww3PiByRT2RdJAgHsK
QEpTIkI3WgLwH6ckTi4i2AhNh0XD0baroI/qy+IJAbAk761agAhj3PzJT/QKi41K1cM5Rpyo9cK4
JZHezQ3qIIq44yCLRsDJXf+YKsi749++96AZpVVdtK6hkv0/Fc2AJlCiriVTq/V90BvkNpTc6lFh
9sbmPZ40ouC+slonCvhHD33/amXZ9YdMTO2t8jVSpJccaW4EZ43oCUurctKZf5JjKXedz+mko+XY
8qBd0a5l4iCX/ImVCSbuVzREPTtW+bZmoUw4tmgC4dqLcIQJH4+yzH3U9aWghDq60//2Nm+wdhM/
ktPIZHMtiOMcm+mPYe//S3fD6PvpmkOL1hwa7sEUlnssU032EyyY0c5sbf3dwjU+lIpT4EtRWSPn
ii8KXfBGw3CKepq1LZmnXHe/yhsb7k3PZ2sx6VqqNFwH2y+ieV4eegdqiyXlabOL8cszJr3hCkEw
AppNwsuXobTBRWB8w64f8XyUQkzXjyj8tdBjvvdZLS1salDSiZcqZnm5wrY2sQUqeQGi1zmQe+U5
IYpgG4guV3R5SJVnYYbLcE177syPLMCT8T2MEcbTyzUQMhfg/XQfdION3hMOd6YAnhbhYh8BAaLE
e4wPVQtTfAwcBYTSxYWflzWiVGs6fmCQ31XQILy4FfmK5aVpGspirYZcbg4dkmi3RGF1Wd4sJOcI
xnCzIu1lUtN67dBq60xXX2MmuRox+MvEuiRwiOj+Zrvrpa6r9/I4TpmbqYB3MwbYKrcViBXGAeOV
2QY2gDB1tGB5h7Y0pPzh0lqVPwjWv1sdoVaYDEC0D6yApoBSYMmrlfG+5s8qPYI2VuSgIRlQUCcu
rq1QRBu49RRfL9RmMQ2/2KP4anlvODTPDlpLp4eur4Ak2yIDChwPaP6GJmDD3Np9sVWM3G7y3l6g
7gOVz5R5imJCcghbUuikfiXTsrAShQEmopW4x3YWnS0IaCPFRpEZeLRg8w6C/7nngrn8EdLnRAAG
ZJYeYnY2rtdAXFbGL11p1JcBCC+CGt4pouHOu67V3P9q8dgw117Qmajao9XAv+lOY+bYuq5BvGdP
uBVyWRM/xHqdJR2B00eoNB1HyfJoCQ22LgQBztX9/UTy4CtWi9U2J2Hha5aI/cz6bccWbX2Z+eSO
+ytqGFFkM0Y1fBVFloO4Kqy+xxQAjK9F7JeDjYOOz/4Uo47CRXqenk7aqXJOwAnOgrxaQU15yzFk
NRMEmaBIODVdW9HhhwDKduDilYp1TXu1OC6kCjiL+CZHGjsd7ErpX906uRJK3FOQBkVtu5bC8i0u
oorZDstHnjSW6h6MdFzElREdnkX21dQxca7XcaR6Gj93+ObeNtNQpLyFlXx9zJeDunHmX59cLCAR
BwAFI5S6vKdxToYeuv/P61iBJZcko1qvqAzT+A/BeJmyaXuKpD3G7w8C9IWZMX76n5lWgLuH5C9N
WvaHs+SxCbG/G1iQE/ZPZ7YxceRi/sdiwLHnTmAUXFr8m4JRG0QhBVM3r7e/2yBlan0McHfKFNoy
jQkFBrb6G4AbSDNki34+MoN7NDT6R9lpk0oGokDFHuRmcXE+lpD3sNMxferUgqfSQ8BtNoSQZHWJ
DbyFc+nZAPbExccsLN5L60nAY5oq3W3YbRSbvLVYHwc81EHIlLmS5A4EdmsaYj/Ky7PP7Zfyyz/H
dZDcuUm01pLsNN6DtLmSa8t2qQZqyNHWYDzwAi94sxsyn0yUo2NDKvsuSd2qDJl0PYzfa8kaZ+F7
0+ImYjTKoSda76vkUCbk3OovIhoeaumVMWXkWhsLqH97F6QINAlIqKK0wCFsFOgVgnIebdi/Ypdw
UeQJJFecH0Rhs+PF3ERNS4/FXgaI0R/i6dEh9SjagcUiS5l92ZpTKbYjG7NGMo+7mOiXBFA1a0H5
CBpcjbgvbs07XDnk/0DUjK/EFc9p/BmLGYnwk6PCoVxSe8kNOZhovyu2F17zMPceennSHFiPNiGh
5Lu7WSgvUNV6TXo6BLbylRe8UFRYuuDGSp9znvHkyHRwrh2VZjxAFSw+jha6ke7SxmgF0mzaR65K
PKPzquf0KMPM+h8QzHTIYABs1bTdHiYPoACDXRW3wgtktsIyDkNzPLD+v/1+hRJoAn+LDyD12PHK
czJmi7xSaooHDra7z3a7RfpogzqYyuOhVs3bpmV9AVCucHJ/J+4mzeSA89cGhvGz5oA9NnGNfDzA
9FExmUmRRrb1MLMAvF9oRBOZQimTu91E39BquptkM8a8di9t9m8wAUHatlXOljXdD8W6YJ15UxUF
a3RVcYUXBWWdHyybz79fTukCtnrbzf5h/8+nz9750JkPRPpDcwwly7jareoTtabcb3X6wQ1SiP4p
MRfxxQ6YU2QJJJ+2It8cUJ0YcBZWaNbzrdgem3p9b5VlPQSFlhNiegYp7/PLlQv3D+Do/Q98/qbB
06ptJL/C9d1A+kbcC9TsuC1PcrQxyc7QWSimNdFKCRBmUi1XJndEnkMbvxeLSQeQmZmpPEskDACM
+1Pw7UUtz837yANm4WQB78mgXIO4t0Yz6ts8SAxVp2oV1xqCC/4QtK2l96pVaF5q77b2pjOr/D+L
TgOsWmMYYZohN/hB4NlKLkiXUmfy4BLxtwVPNQiIHwFJdm6xJKJtfGv+9O7ZRJ3I4/VKX249JriL
4IYqym2tmczXmI54z1vW7ds9KVbthBFTBguASd81bxnpEC21goehJIWu86SNu/BRaz2ZH8a2gAXk
beZ2QZeDPGqfvFkfsTBEtVH4QVYSZd1Cy4/REBrYq6EFM72vRiCnl6Q/CZpydpgbfmKVBWwCPYS+
3zd00Bgarm0GMYQak84fEpqR90vEFUFFICGFjWc/otMaWu77qVYLTXtfGkp73poTnf2WfE3Tvbu2
c5JfW8tS+vf+nUgZq+w99i8rmnlEJylDR7QlVW4WlU0G4QR0MlgwZxj0QhIB8RhlWHuzxYKRzeXb
wUSnLRN0A3FqHbzPAMr99AgwHo3C8qwOpMmU8Of8AW6TTc/aazZX54GaZnA2T4pMxzs8YX75uIeX
J6PofuiqASbI4KiFCwOQNlbElHQboF1kWcjgFMYGWIpkXDfxRZ+I3nQq5Orjdfx8pP+su2lMCrO+
J4LQFtuHX0e6KO27470wx9kGTrwhf5O7j6OMcwhQeJLzNGq8UQsFTH2Ce3Cc/ZDI2quCpcsOQzHf
cVwdrxDWum2clg+X1Z27SxNktP4adln8CxNYwgPDD9LgVTzeK4A4t3fLawgdQdX+2ACGLle07VI5
ufpfFAtUd+EKm33Gu7os7SgNHzoO+fXR98TG3+0Y1pcIVWencn4p8oKPWieUK53mHZydpBSUGt+R
ygsgijmC7FAEfRHJvCcjTww+BE4E2bwciMVWFkkQEvBYklXS2l/wCf5cmQHhcgG8yNTYzGeEBtNi
nAt8a/pEGsxq4i7Ugkt5sw8RiC6Sv8Meb1xBQdUoKq7kURGzxO+S/KcSeMWId3jSsMfqJ1HcAVlp
4SgL0UMYUfAwAha8AOpKuIi9rO04J1OKF5GwUoyIT6UxRB7aWAWeLU2HPFwj5eW10RkcEEnsUJJB
LtwJShq2jlNqvoHiefmdnaDjirboUU4Rch7O5HTkeO+3jwrL5JnO4dMUG0dyKANXRyShWSMj+8fP
nnMT/YXYxBKO9xAS8GF3tcDEIYaxAOWDGlvGE/iBkmU/xWqegEo3O/aFiNdRmd00dHJuOrKsDAg4
fUK9MJov05zD4MDEkeYC4YsY0itdvyL8EyVi1vi9PBQOzhrKQDYb+DqgnHsZnQqWB+QgLeZUobxj
+IVLb7vJTpfbXPGC1lae9zUq+59ZlOC1PkqV9tyRCPemM0FOrhppzYd8zHAP/XYIHgfgO3qCmOSD
khsCBhPV8ad0DMnPdFdELIY3XpNALn6U8qB6Zx6iP51meAIbCQjfp3SNY7Qx6nrHhm69cPOvzV+a
UazU4E7taI6P8DPoske4TNMjRpXcVENNzJSv7BftubyRZVE6Lpat/WDTS0pZtbuoPqqFTI+sJ7Qt
YpIsRf4Z/xdRO2XcSAiPEkVVHU7957UABECJIpkgM0AceSamhkX6CquoBTmoOu9co3/LHPx8ZOBh
ujfW19KioyovB3/zMG1UMmhCQJQkQmsKmAtcos6YQ+mStsgGpuLT8C83ihfKTc+RASZb9c8SMd4W
AvlroJ7xihCw5O0EbpVv2wPSxk/348+omgtCJHYOY3RGFZKBFKL1wrFO4wXfTLCIyvLrdM3XUmEn
7bBzU21jif1C7gwzLSK7XDBXeEwpthIxCG0U/6a5jlbtLbJwQfJgpHbTML5elIwSesBZP0nimkLK
THUxKeBjuuuU9OXK7S1vKUcN9B6ysRNh22ZHdebbajbd3w5VgGOZxYI4Dj+gmJWQ4H8H/L6wOj0g
7KNoWI4vEwncFsV6BvJqvF/jJILUW2D+hhVh6+26QKTgmOJGjcM5TGrsC/KzI0wg5+M5kxyyvB/U
fmFRhwTSbMqV3yyuYpJYo8+p6VkqA4y1aFQr2woNJK9/JZEUmhaEw1gZoWPjWH1E07fpewRMOBOO
vKdqYMMPvq/JY6skGAoj3G14VMgd66tiiNi7Ilefl5QHA2WP3IzmbN8ur+OffBEZp77jYoG3JT35
/Y737ltrFEBlGpLTx7tHH+J3QFuFRbdjHCYh8FPXdi1bYhaeftVfq9j560ULSzd9x6u+CoULvUXX
Ks50B5Ug8zyzUOG+Qgzn+vTQBYu6KUmkde7aLv0CN9SdsE99vGrGCHGK/uZXDt62hckZwTAJEt/4
d43MLRUqJIEcJ/p7VOLIBOnLuwQoHpOok3AFf55R1/5nsuYj+o8bh7ln8VWsKPOV50FFnmJ193h+
x2li8C/TFArtTJB8ZZapzD7huxkm1jkfX2tKfhrHPFHV1tuUUfOGq2OnWqlkZJvzMsPM7kA4ejhQ
I0wTbSi00OwrGLNi9N4Iw3368of5UILXYi/Rufeq2sjSKt3QtzUWFYdKHA7NHPEKWbKNx3LCK0a/
InXDFeQAHtRKsNUDliLbfIke861/Z0k1Y9OjhJgJiYV7GVA8c/YDL/JCGA5cWPCtf5CA2CSB4vz1
1pJKLhIo7ExQsKAWK5y5BuaqOZbPSqMMHBylwZpUA4eMT85Hk0RiUX4KyYgQzOZtgtrPhEX92M9k
9k/2jEY02VBDbr5k2P6RBsHPN2oGoJKt5Ap+hqjUhHyhwMNaIVSaIVjfxiwYliM/c3tOU0b3/1+a
+0XxcodQGSZ8pMNQ2RNbk0tdujf4W6hYQzmsXs0+klqyzIkERqucTq0+AX+DpL4q04FhzuyU/B5M
SSdsRE/X5BeVk5nmzAT0lcReEZ2mozLL/Z/OnrIrMBRzbnxhDTijbIhBOZts0W6xEM17v+Q0PtUC
IvFZSo6uu8wAHaDQLze8TFUXeYQMkLnbclmvqIfZlcOgUxItgchlFd+HSjyXrWUltfozuQwH3TZ3
Aehxf4leH71oMNCw1W5lm3Bd/sesOF2iEJyqJU5Tpb9+PJT5bLnT/ar+BzQif2bJdtPr5X395+83
m00KDBk9tJYW+/qF58hSgSnobKm5mQ8csNQttSnFOVMvtvti8+DPtpfXxbP1fuHDhzXYG3d4nArV
LnIOhJ5E3rHOZ2MHWnWMpHCZx+7Sm1oSdDPS0fAunAcVnu69tRkkjB8r84M6faHrDMBZqNMuyb48
Xj0gXUbM/QVinyz0uIBV++hJtx12QHxieSZmOgfYOcADae1zXrEj8CJDLgHR5OAtg6HIO81VT29N
g7Nv1GE07Wjd+A21uQHKkDOdFHru1YAg24E/YAoGnVypdlUi1wOa8/i7FH8RpMZVQQ+aoEa5TX5z
bv36Ym575eblr61KkpwP0NjKE5S45Na7foz/U2AKQkpddowbUyn7IH/yjPWisZiwYwr8GTP2auxI
NhRb6TEniFlE2bCcxFu3HdUNN0pFD6YPQeQ1mmNDAQV4M7ivWZu3HC6Ty01eRQ8tuKRrJcIoinlC
sJcZ55cmPqlnONGefQ5z5aeCymhyarMnrYwwi1gWVT2MgNhycAmORyqsTLnPw4eK+k8Z7M+xaEGi
75cP5vlqZPtmBp0wBfGv1Wu6wF/oACol7MD3yaNhRv6iPZrwu0yg2634iRUBwXvx0GKyulVbGDkp
YmNnMI9KThRQRz1uXWjWY+qVn7ey3+w/jjfbfzw1hN8f6t/brJBZN9w3CL3T4RvcARUdinJ2r9zk
Z5TKwUwRFHzEqnYAHA3Y/GLrTQUInRlVB10GsYMtuPa6N6sbPkDDZXNBR1Idj5JidsHmbfcVhcLf
qa3fQlBHUOA9BXjN/UsJZPFZcLPPmd2noNMHlAWYJhU6tSIq9rUfH2SR5HlVNXVZ7otSGFD1Lzgw
bQ0d4RKWRlWV9ffmpJV2EIqgmJ8sCs5G64vFvgZSnF1NmKL5AnZXWkYnlkc0FMDcmRuu++j9NXQi
cs2UhaE4mTcvXjeIemKTAe6ZkzYzSpfgFfy5+4RjOb5YljvBUplhDQ7+kCvh2Lc9HVVzPTK0TWid
PRA2Dazo4ymuXjmQhfmdEEG2q+HEx8X2eknevIkoh4lcWCwOcAu+bhh9hasm0kw/2Qecuhr7+5Ep
yEg3F/UQsbT05bQbUG242OtmJQoXNEbQWTsL5ceH8TVo1Flp14tBIDYLuDGYoHL0ucxwphyymh3S
Q1uK82TbY5OkjQ1pydJOd1I9HimeMa9Qy6zOklPA/EOAq3goqPQduvHOMVZXIM78Px/UeI+ImS/H
x4levRLZl4El7fsnL3ib9XZINeimJ1ve2+5NJF6djLNGhASVHjpufKoQUpQVrXvHrZ0fXPI4Gkxj
ZzmVfFMhQJ5W0pQWsUG9tOiX3DKohL4uGTKDwte8eu6cUK9V7LSka5MK49qL2Ij4IhhL/edsjaK8
25TZtVobGJCgTVThZWSjKie01IipIWJN4EJ/SukT59Tmt7y4v0OmpCrw+vAWsfVs7ZtO5/R3q5/v
Ve4+WxYmMZtpBAP+pH5F7omg018allpplBJDchUHTTl+ASslY1ucxwPmp6vu6BTF9a6AFimgb/TA
UmO9IWHwudVmBsK1hJuwZXB5o4B/n71HKpyVWpPRroQrs5pxBbHPYDppMlTDlQ2zDbD6j64F/DMC
x8S01O/nFEKviyn5CqK+m3E7gqJQSRDmA0kpj9MDKWGjqmusIM+jw/7b77S9SfOKUchZV6WTZopb
SRIyi+ZnSJHy0V1i5lmQ/W+bbQ37LHsvCx9PSWBsnGbbcXsXfNVnDL/zTC0sYx9Dr1HuhdRVtIF4
5HKuwhm8j0a8W4CkHS7SWrjogUA6s5FgR/AX9fdPT+mXA1BL7zyh1QnVeS+uw33iG1hiosr5RiDP
H7AZTR/oGvfCff2HOyS/y9th+71QR1eGfXfhGpJ4RchizZzcK/LHJVzzawYRtmdu9q96t2TJkoYC
FEod3GrzHnANsPyvV5639v45vVHNW9ONY3WCX/1M/GS+R0M6VBWjX+rzpCbjULU/YR7AZm++/rB0
P23dnlYDGBLbcHu1gAGo7jKyavrKgfEoEB2AzNtKuWewGkKfS42b4vM/tV6EqPge7mMTN4nvtsxL
7Lh1zke4xtacqn+cPB7r4r3fgMw2SETNAl/r24AMGee5SaeqhCaDnPtZlqrvVZvMC9QK4wFaKFZO
eBDm1zCHHXkJO8VHf91GSKO8wXEU+pz9zQMAhnqrbDpSbQRtnY44KjnDJY3iLEpaU95COidcFEEB
HJJfzAYnYZZ5Tr9cd21fufFQswN1Qk84JkIPh10lJ14ULyz3Br/aJq/fHJ9JK+Ae698Y+vAYCXhM
G/+8LvayI80AA9vycrECsLTXK41O2CsaRlCM6GcGNKAPUbkg+9eiPejL5gKqOdUduAfm4VEX6Ti9
o6/6y4ZCT3e9tMgVCYgHdTC0plLVqbTsn+fYUe/Gedn69Vww61eJbuz7Dl9ENZisfWUvpnnir5qL
g21PWbdtRFzPIFrNchrt82dBRa7kDBe8uS8oaLqubvFPkiDBOcx/Vp2lQJhWt5oID9gOUy1BxcZC
Ovvmx3H9gS5MFl7JGCVUnr/OPRjpwRCNG8ZlogYopPy4J+rSUJe2ScoE5ei9KWDKJ5Qx7qcyWxib
VrzMMvG3uEsWPXmxsDJpY9LB3y6DFRcepmxVXEBSdnVJHz0hBPGiTLWsnaKiYAwlgQMMXCvlIcd4
FuqfRA2U2wEbVKqLzfmIrQCrX5EdPhIlAgAJBFEaxykFDF/4ms7fDEZc1DH8nJD5IrDMutRmCjug
B43iFWdyE8A/iV+A18yrrk3hWRLZzpKjCFBPHiEB2Mmtwj4apojRY5fPBdWgLmnd1/8nFEjO1Y/H
pf6uksg0uDLadaXYtonZuh/eJn6vP3CKjM58sJtEyjl167ZrpM/yXqo999RKroXf0yUVMKAuCcTQ
EBg7RobTolC4j4JaTOpdf1umoIBvhWDrysx/HR6mbcTKM9ZKgrsIGyCc2jVav9poAQncSUWOgeUi
qGdl2tgWBblaOegJMQd+xDa02t0xOH1Ux+8/reaFwiO+VNhmr3IsF+9tiG6N3twV2tt15DYH0n9w
OyOkgu5vf+ZyBt/xpnIGgP5PABSpFw+1w0hFvkFY0Tu5cuujQ87wdBYwEEzXLf14yN6fKA8l8y0k
eFdyV9T7uPvyqW2hBGzIQ5hTCAbhZXGDQ9OSi37B+ooJg8s59l2w4k3S8MXhKaCi++ymQjPttTO6
Yj4xtfmEkqjvpIaa3SWTn25wg0yarMRHWo5iMdmI4zCHSvjFIl5fyqoII+zOXOosNDjwM8ZwqrWV
Wg/oEn338C5byg1woLmFB7Y+9MBAfil01Xe1YyTMISB/FqpIL9FbxpUkoHNLe/YRpmArau5v6t95
sl4mbwTdsbt8kKJPSTfzXKtbVutyiAZgliKlYYsrlTG8Os5sE5sUYLmg11ZdT1IsyHxy3+odRRFW
+hmOHjtkoKu9iITnujyRPaTUa7Ps36Jnsbmc7CSo97mfrJsEWoCKuUPqGBGjtKMtAOQNvNAjLUAu
pUdAhWqCDAwYiQcEy3UalrnEf2Lo0q1PBMMgiin9l7Fmxlzz414mBQXrVXtbpkey3PzJ0EwbcfDS
LJ256fYE4cuMzZf0to0av67tHM2sS+Wsi1cLpNx0eITbV8pf3DafruQyl7HNTeop3KTZC7qCHbEP
goXu//5r0bmkdeoJDsBECLXhO86P5OIuAK8ArxwAWMCbGCITtt+Gi0Tcqb/VxUl838eeJ68nRa+s
InpMRrXc9WNAHkwMoWYortmRYS87irB8Z7vLPEHpkTUNg0Dx+qCOMQ0qkXAfCREjRhiGpkLYTu3i
+y8XSqisE0gfvSAbBzehN/hxKurlkHHLMFHekXHtJHXztesOCneqVdrtjHwg0CPNZ1Kv1DK1MFfD
GJk5S9YuMVUd7bJsoRtHmwuElBwhie5AKoeyKLCvAM1U7LafbLvDOTynPsqLcf0jm4gO0adhBlXg
sK9h8/KgAB0R9Wmr4GXO/5vrsgOUADAWXR4N3VZFg4XKDfk3xRQuwAW6t8FjKp2ecVaqYvcI/PbC
5m8//58FkbDjvCsrm7vH7MweG8k7ZfVIfK+jpvZxzqRmfyqQMf5BohGB/lW3oa60proQfv4icISu
p/onLvckIWYJsx1zaq0IaTOOT0ENxPh4bMM5uKp8ixRVmaQScUaWXJaZ/rz2zTIJhIgfYihjEz8M
igGINribRkuqUsPeHIZSi3Aeg8c2kkFjKRCH3xspz8QWhOvlWEty1jazmjJKV0I5kYBWgUcMZ7m9
IiUsTUp6pfgdWBUt8vR4t4KqYYqHeJCJ9wcgSnPPi/QfFDeA38kOMvGwo2F5JCMjRQTqEEKe3FUU
O7Y9J6uecYlrLPElscWgiUllDC8fqEcLp1SPlaRJ+gmh+LXbvuxUvB6nSfx9gupb6V982cFzPz0u
xBXvM2UUP4+rlALfocwT1yFpi88ZPUhD012vyEMwMOPJV/OrSWHrh3GZnHhU/Bkewp2HYgWazDOz
Eaa1Q1x2dfap8+t6LYi9r8ikCfXbvwMIJBCWXWUv/fz65oQQzKmxYAAyUHdLc+mHZN/eK9rkTrqe
e4IjyJ9zQZn2Ru+qbcIyx7A+kBXYog8T8AF98Gfu1toDqWG4xKTOgUQFtUG2Img5vZ3V093COTHR
fXUGS216UqYMkPb81MvsCbrTvSkCOfyVnOoKbALM2k81t7+cL+aNeTqRfy1b0UsgIRr0pQf75Q/I
m6bACBxmNkFXW7yXr9f0KJprQUlRWRPXq4aXwdnZ/rgriNP3P1d1zM7rtHlPKAqpp12DA5XYwexn
m4z2Zq4XvBFDlC5O2QQoWO1IBBxhs9r2ZdHOHVohwkq+uZOm7ntnaiDFSQT5PAmOxFhXQcGFMjvU
DFowJPRp2IEn77htv0PYIfwIEMXedurShwxkHwTO5rav4vHjW/Egya0Z6rKfvJPNQl7W1VFHL7QB
W+bCOF1J312m7VFwaEPMAeutjrIhhajSub3kMTa+PEQVXcGYHd0AjtVYA8SyrDeIUnTXGewMOqt2
0UFmHZMvi7MHOlQcwtTQiRo3kcmjgkIzEN8sibpnPbFw3BI5hxyKyFasZWSshbO2YJEKjHz5FO4X
h3kKfTHTBbdj5VzWwDEJRXLGgxjeQf8aWawX1wEMKwr0r2LIyIonmT4K5NNLIjt+aMUbzy/+4b4l
sYGQfhnOqP7fVWIg85XPHPzdQ3zCrk4mRu5W9JVqVOXWBvCp7d/ubZDRViO1/hW9Oij1yrBZTOCh
avQWIJIzoHzigtQP2SgA8YRSGoy7erbI1Rvuvt9csTFbbNpZJgQ/wGf6Su36RKYnEBRZhgmZJR8L
HE9anPmP28FpB9IZrdIYszpS1+2epCn3OfPmpT0pVP99Yg61dtfzlG30SEwYz4a09/AojsWBA7i/
7xFw2bc38+AflaK1nrFbcmRDuj8JhGRRZ0nxsHUyIZSKGf5t0NC1rblEMi+H4f2uKBkL4T8N3wBc
OQFyw8Ekj1o4P6WX1yLWi/RBohNoczEaH/uKtlWf7RemtxpFk5TyApkqe8j/3yXDQEcjCeZjd9qA
gysaO4FCHjs0xHv5ecZSTqUd+qLHn2wLg1hVU9CV/BBD9VH3Zw4tn+/Sijed1O5sVQIK89mLnp7S
UyCjJM0fjnaRwloojcyG7vdT/kgudq9tG7XwnGdgc3qWNkY1XxaXuDml7c/PqZs4Ao13xVUZ24kD
KKIa4h3H1ZrhbnS12Q5SdT43HmyxdJZ3ehhJ8MtK8dCtTVRHvdJ3j25Czwq1pTAFWH9TEglblJZI
dZdoEibfrX0SG9juzN3JR9ydC0Dcm9VkLV+Y74rkmaSGUyqXDWTNNJLE21K7sFdPpWgqUZmbsaGB
iUJfrhunCvN40ZH+LvQ8w+qj0IDQPZyKUwez+IWfd8lHts50lggvpfVfqDdOhT/L7wL0u1+FmE/2
pUK5pPXWOBbQvuS7uqJxz6hzg6tbbsSrPePLgulAaE4gyYmjxPGVWlgZApLWmF1LHrLFiJhmkd43
iQNQEIKyLvVZ4dKFopK16xhD6atHkH+F7/q0qfRzdZFAOJI5O93zLaH4WXnAEV7h3RTPy2BOXJ1f
AGzn2cLvZQH34Ur/ZhwcOcmHQ80FwL6bcUxFenIY5uZGE4Y/OKRtjmcCB17I7pN2BeaucOTDvMZ4
LPC6CJye5ea6UTJPG1hpQHA5JH5q2WpSHVRfv4a94CbOtYlQxCKSPAnCVlZFM6hCj6+0OUyKUMEp
A94qyC2VMv2M4H60cdWQDkL9XPlDXyPtYDdptVxaWP42ho6dfR3UR3QQijvO7bvsSgFLEcIe+DWi
gM98osKJkg2aVu00m3Ay77r/t/M8fpmfuHXGn9B1ER2n+dgCYNYx7gd7V0ZsGLuKuVmVjxeTSrFh
yrOD5fCDrWRjO+HYcUsHdqFA9eX9m+jXsDkPtGDox07RdkJ7HW8xxuwDU6+kQGzHE4QRtXB3VkpT
mAcmVGJktivvb6UnKOzCR/8jzBXeC7MBWHvsXTZY79k5QvfdF4vgNTJQsccfKafbuHPwmcYeX6wZ
Kqdpr6DIisSOfUktdxxh/wAaGV+iJeFuCvpG4/aAJhVOM3tf0Wu6tdRUoMxMp+TWKqaha0f9xYZn
/XMBHSKkbHy0VFHY/HCICiaTVzzGKrAKSmzCH3Kzmp8KewmdI5pcWWBK64RVrUZ5dSC177kDqmCT
Ir1eizeIWPcc55uLuzUk34NI+o9SUFqAGu6EajX4P4penTWCWDYSMwlyKGDPsKhbC5OspZqNKNVe
eSRA9fAOSDJdSo9OLoY+o5KeQ+y1eIaNMdXFZg9MCHfdpQ4Gl+yTwiIhfCPgWlTiZoXzoG5sZgq/
/zBaVimhUI4leyTWeGW42GnE3pbgxrB3Xg17NeBNanAy30RcB8z+UgPEbpl+LWH1oNtowjgoAFPp
IDrOd6qVVxgh6nv0cDj+qKjgiQAtkgqlLgM9G8oLoP13/zUwrYaKyc0xH+8mbk4W2GpTA7P0S5JJ
WFjxS7F3oZ2nE6dUc6eBDdbruw5DaU+z8uAtQ89vdL53+J+PwNZZJNXAkTNVxgY4FzfpJ0+Ch88S
UQDTxIGACFpaXhk/t5NqfCz6KniAiIkixtOQJnupqcQ0KjiZdI/RUe8SIIMt0v8/zVp2MqPC2TZf
6/jAWctFS7NNgW7neD79bdCmhWtHh89edJdb13jVtO+8tUoLhUd8ulxPkWfps8xp8v0UIftGPnCM
TXcSUUZ8ENJalgFI6eI9HLqo21jyQEpjGk+8RoMdOucPPnNQiqyWCutT/wKmWRgj4AeRoQrb3JR3
FGhvpcwYzL9v4wtXObtcFwu7D03DNeZVzPpPtIqA65o1v9LaNjvZosbivZw5a1X7UJPQ3XzhGcQP
5U7qA443KmpbJjT+/RDiNC/30LVUATba4QUvQANqUuVA26BR4dP+eBexbfklTPQ9VNjyQtPXkyVn
7qdEMJlrej+tk7UF/j2pxAXclMfyzr2Yz7jFN7pdd/UL/hChMn2pOfMRIeibXt7S6a9AJPzwdwV9
z3Dl7kVs9PXatTGBR0gl4PKmqXegf5sLd/XUY1ewntO5TxzG7Y0KNdsVtU6iQK0MGYFA9GFFAnQF
jvF+HaKYndavcqe2d+scLvi9QMZENd24JwikVgnEy+HEGFk4Z1NWcre6UJaWX2wBt4WXBjip18g1
sVtgILqwR+Gey61tJ8ITls29cIsYRnPvSrFsosw5ur9oLiUG4DVCfAh80vVqQUsQJzSOsa0cXOcm
BuTd8SI9vf4t4NzL/SSFvqiv2jI5o5MuSaOO5S6ZfWlaCGOjluwN3DwAVUbtkH0FcQGCIzpLr+xs
/HKSQx2Qk8GmTEk6y8hqetEZ8zWk3U6HAq2l41mtnQ/1FREwXrR6TOqF5nBFOLO0ITxHXpLmePVM
xk0V9M8WyRhOqqcuxUtVVaQPpGveVMFEc8H9+KIKusq68zaUBsiXZpjS8Abey81uPxHlGc4H9bQT
+D1E+PbmvhtlfLYWG8Tg9Yxgpyl9kTVFo+xQ3KGSmT5kC8+WR887SQf4kl/HsanOarNMTkAbCoRM
NP0YD51Ip4sOXZSY5XYtXuUW7AQfq8nEOG1maoPk5+kl8etxjAHOGmVeLsduPEDJUTm/eNd8LOc4
fKyqjS5JHTA04gP3mxnkPmX3oqz5aCR162+kpIwZPTN7zyDgVJbQKedlreyPibXFhmvh8GbiKM6E
//LPfVd1T+DGUpoYM9IDODDnIJNU3kxrY+MKEFjzIGJWpQxZtIjKQghNTyV01Z+vKp/nePTPYTcA
DAFu5bQokm0TSrlRIFxmpHXA1gBWRZrXMkSLgoNi1dz0dWz8NLOv2aQ16EpFbVuAaXJ0UpJQbqDZ
UfD+r5qL1xyy3k/Mj8BiEDhQyDMZWPunpt2UbxeykUDn5XlPHcKdyIYZeAOvq4c9XBRwvo37BLNo
TznByFfSKIEZLOdgzRtiymgNguxtR+5KJbX12OcT6fzn9Cefh43cHyO0fdv/oOOCIOzG1J5YlBdy
v9MFBrA2g1IfSom0Hup5ge3RwCCLom/KRRSH9D7PoWpljT0aU144s55uoVHFUX5eemUC+VuejjZh
0uIe5PBJd5yE2chSUJRBjgs9vhJ+U+iwV39mpa3eDfEWBhhaA6qUdgVecxFxEgetRnp91YQ7X89e
4l3FYQIsZJbDi1N5o3ZkI9QG94c5exifn0ue3AYEaZbxy+adSaw8xcXlo9XZgO6xRaYVICa12Zoy
Lp5nrjl0Lw6MEqXRU+UBLyTWIaSuia3XzfaH8KfnwIH7GYhQrhej0ml1jmRLjVPjnWp8QLss6U6E
g1j+uKiXEpvThi95+M3rh0L6QxykDGK0IVimaHeYH5OzP+qE5VZzXCw9WVjCCDpC1qKFGfv61pm5
Y44TvHm6W52PyPzOkApD0NzfIb3t8cEFZTWzv4LrTnvHlXHuAhz52aiJwDq/f3QtdpB4R6joRvRk
k5WlLh33KucuPSmMjQV4dViUA29E5Ecjwo4e0JfHtAthic3Om8X4lOCWyAuw7tbKNhUz+fmvRJ1Q
a+ti8oz6gL8tBfOHZmFI7IJvYUV1f4HJkwe8rLjBwszN8CRCNvvZ45nOXHKb11IKeWv/QQ2xdCXp
qRSoKsSWZuiefP7giGjZ0FqN889G9tu6OXv1tbihwQRYjE7qrmHsAL47HtEgUNrEcuOC1HIiwpcz
2dgVjnvnohZP1t6QVYBvVdirX1H5aITFWmslf/QTNBNRWro8XNWGMjdM7LJTjd8J9RKj67iNH2KH
cUZtXZ1v81SiNDNpCfbB2DmWTmSAiyg35KRfyBh9CzjYLhnrJvWcndvm85Hfk9k6fx0c8FWYvfnp
PUrnTKyHlVthDY0x4NRJXH7rj1BpDO8aSKiOeaU2L4tgFnxOs8G7PfoSpJt9DRyPSyQB+kneDxWq
pUpj4uoczJq5BfkDLm3k19jv0m0LCSj3lnBXtIC0UIeHyUdAWHz4czcB3hQvXPq+PRht4WkyeMh8
Zz88XqFw5/WYKSSmWnhOXKLpsmeoRKA0XqV5pGkJhQc+bGNBf1ZszNpTfNGlmMSrpnevdylmuMJW
Jbj8BbV/QPCNc0qjETHSbcdbF85XraOtBNyRJbW4JtoZswELcuXtHPnDF+TDInOatuZaEivkymSs
/R0mZQdQIbIgLz7p9SltlTGTG4flc+JCYZ18mpGcGMLGSWkK6uWVq0tryjcv+OZAlEpkTbSv5ARF
xIEhfbkFqfYtx5NmdBCQ2M6I2GCDvdeb4AxyHHVhmimsUCXEjTukVb4mUKIWO5dudBy4K2LBa+/V
uKl1CsIuKSVa7g3c3qUm/VCUo5X9yEuHeyD92ixFUvm9VxQ4s8MSIHsQm8+AG6CzbgOWLwYqurSD
T7bjt9v9/DMs+O5uSo6R4a7dBx3fbESng1DHwr3LoIywC3fZUZxPzVBOIxkJM8hbgiF5KpvtraaC
vuG7hRbUx8yE2bxUkeJcoeqn1BnLJZ8bF55gaBDW0eqsoegHU0BQFLiX28y/aXFGDPOehkuaJsG7
qIEK3pAWNetS3zDuwaormhq6F4p5iap8RCgBaJ729LwW00tKP/CzN2qwlEGApSjf/gnckzIhG97O
BN7lEU5okYDdK+yMNspQ9eMNxRYcLLyRZKk+hDMBkuxJcn22CxowrtA6itBdRfJDwmh0B+BzGlCa
0rUSks/fkmQiVJ3YCXAaBoQkchpljNMzCD8ltbyugsmtH0/nMOArLWqo+rtdUiWzPsfMIk545XmT
AlGhYu4YTbixOdWLaTC1ZMFOLQqp0nwO/2fp397ryqLhUd+zqiLdFucYUPgWAvN173h5YgStkQTI
4ZqRiDtXubMjh/77b9edFe4mwKBrbRe80VMaJlQqqvJsxyacxET0xiJIoEgt84uRu6NVDZi0vr0y
BBjY9F5hN6c2bDIedyaYF4G1GL9u6MqpGdJgNzQLVeyHoppGS0Iv2NV9xAHwSneRWmZlX3EROGii
nYWGzdRXXilP7ATFHYeGhuwl9C5pn/nuNHsn5/JiniFwCQ+O0zpGOhxA2yTty2R/7bRr6eprM4mY
o6RSqdoNgJQoxyRraVnO8a6d1v4dj1hwQNbO1PyrRto4UDHI1CCSK0/wDGTbPtspDU1JjJX95jm+
xxcg20YyyclZJBHXHoqrAExSRjUBmvXUUVfk7Lc6uL83Juztuc0XmFq8poVrJVxQ7vHmleOZMf2i
nFg9Qt5/4H+5b5vm7H6608zpKy8WemgFjWUrhPW1LPWcJmvQg8rkS5W22/OeG4HfXD3L4vBKHeFS
c+f5NTJICWRLELl1d8SzBGD+ClRqZKVtRsbNMqfOoTvAOjslpFC9mXH5yfoF8Rj9aOdYXpNAwbd+
hOimd0IXZ7uDQMqIH9SWWvpQhRPDAJvThD2EmdT8xqZp8vnapOcNz43ZvX3lUePOmc7OVYRf3Aqq
M7ajhkWMeLjus+vmGke7nSf2zunSNM08U57Lag5vb7ulu/eGYAVj3b+Mbc+naR8nNFLyJ++pbFRu
5140r1ks/rWfNml48iCCn/quVXwpA3PLfZZaV1IMjii6hqG7GrGSpdDsQyG8NzCsEeCjuVrGp42E
0+2it5YPH8mKSSKoqf9cgs9xQk7UYfEW8dhIEOSZgp1LZwUEoJiY8fhdHR4wc7vTfkrrlLw3+vdX
3za58j+erfIKD4g2w3IltdoCwOrz+ihiqGJZ/SYGYcKtGAOW1+QJwUpnzXBnsaA05SfKb+KFODQm
qNg6ZTuNwfCd+xiEksJ76jDodGI3m/yB6l/z0+gTpiEaG3Pah1NEHv06pHBTjTG6n4CcFdOM4/ZZ
KpQPYho2VGH618m87cRx5MhtgiBQUPHHd/NTbbHyZHOstBSJmZYPbFYq+vXOXOVwiAh9+Pl/ddzx
Fyr6azIlAlcqioYOaeunwiqzP7Bf28IEVraTeZ/2jSmHed/7ZSyskulotfYdL01Vt07OHldD3WIS
a8fbND5XTtqffIAfFhL/Cnf6wdh9tlfCbUZNAake4YrdKerniRoKByme8NzBIgF371FAUBldtiy4
t4u8WJy5vwO8ukOsa54yd9629lgDFspB6+Yzde2tXVi+AaMRd1su9X1YB97Fp/SnrrFOS4jcyoxW
syD3rXe1C6jRPZ0tKAKzcHn7BkJaReQMYJca8SPwM4u4crhCC8otexWv3eheDHGfIWep1yFY7oTK
rhHmUD7XvOdfgUU5i2JROFppqW7OTWSIxcdOs22C8TxwP3NOZup+4YEd1603nehs0LBYRM6KeEgU
xiFuG+NCmOI54q5AhpdNhO8xj4+AlFQs75xVcH1wrWd5JEgbqEH40VnKQEDFniyQbCjc6lUDhx3U
haWNRUPjcYrKdMyfpuAptjS1DnrRjKxml4vSju81SGh1dsm3eaKxhATo+Zuhm2yua5RU9dlY4+p+
1TO+fjc+f5pvbwGeeQF3rezXkkKx2u0nLKlEQ6jo3fuCknNt1hxWzgyf+/XLGv+NjW62SPU6IMFw
gkNw52lCcvtjMw2dkLYQYIR3BB41TYSH6o2ZoKY6NoGAqaRJKl5qoYOTTOuztHRJF7Q4cErSdlMJ
7PrAjEKxaXyNysd0ffp27kX/AQjEqHOb2OIHsEP7MZvtnU0FN/R+lSieD0aBt6AnpD5b7FLSFoAK
r5fyI9XrBm4uAQsnLbRDNraW1wKVj853jQKdv+fPrStwE7epqEjIck2/eutbBN/KApP5aurHMN1U
GrUORjm/0Pu3J6jbZNsEPIwJ54+3t2+cINDQm2sqEZ5N6RJRDQGJQWdC3zbbJ9aW+OwHSGHPnOVk
8qj4h0kCbLm5zEh5OoQcYZZdCyJLXTx8z7WqkQeODg5JXeP7wgYKA12USmoJubnfQQej40F0zthY
x2jY5tb1xdtUCSqnU49Bv3wyPCoothxLnI1nr8niivPgyRm3bmkbeiWOX/sA6e65qGLRUtxfx5Sa
/5HMNHoU562KwJgZqYPIt4SOosbrmX17/hci9mRCtP3t51aQumqySMbrPEUT+6fbcpLR2ngU1JqL
QVLBhpt5RG5kKKtZR6K0BrIEkEnDM6dAPe7wXjEQL1Aq6WlCPB7ONNfvfHFB3JLpkPfYg/3rGC15
HEvU4ipP9yUFgoEVOZWgZ952N0BlEARhUBa92+/FwKQsYY/4gFxzy8kTZpFCIpDM9v1ABKQi4XJv
HuQFSXhdggAB2M4O9jKmwnkuETVW4+FmoSC/4kpEhmGHGGO8fZpq/7AId0cz8BiPbO17r6NRKVQP
gcG6TS4G7hGyJTI2A6y3voxpzrYPT1lv4Rmcc0wLML82Q2GtqfX3JawK2xwMm7LqmfJJ+GrnJCZf
07PQQ1P65kfvRBLuN9J7iCbeTPQE8n0h6zQxpRZVwhmgJ0VDs7kGKnklz64Wm/1PWpeVrJzS4Ird
yrG2XdfgvP6x6QFe0d0COx/+JcXEfYELikgzW/niXz7XSEZEpXWZwQl190RyZGgqYrwFMgF7R/UV
/vhc5SxrNteiB77cqT0YSTR5bJUNzGiqUQXb5NNBz1O5L49PArGaW68TSKng3hxIE5X3N7mvxXbQ
EBrmHSePma2KwNAcNWrtXZPB5Grkjh9hqctZ4eBm0euACJSGwuz+hKMJfgOTOrPCEPtZDt3Z22qY
gcLYPs46uIPUhfxZWA0k+FlaKMXykxxsCY5dUdWHEOoFIk+DpkrEu3RfILQwCAajiNpLWi8JJOjm
LB0AcYWRPEvbHQIUo3V7OTDIgZ24dKwZXZ9/fM5hApaApr9lhdZsayV2QWKzZi/g25UNoAa1SIBo
QoX1XL/ihoMJhXZEP2VOIWsMoC1xUvFMWo2x3PpFe7gzTF7XLVErlzlMx/WNUgzNYolXJ1CM+IxC
h7dLg+3XL/u9JysMggwDGrna5kNxNemx/G/HAIMyVzURkW19oOezkK8i5XlpH+oAP3Lo45cEPZhe
WUVQ19DgUlqHwQKm25S7DiEc5kS96oheQ1svwDaCB0ucwkyDxWU+a0Oed1V3DcsCD9UtdwgDq1t0
2UqCTBDXS3g+wh6i4nXrF7bJIx4A5t+C0Q1FBB5H9zBBBmjRQ0ApBHkSXe8D1eoi14RFwcUX9b7v
Uox1ij3xevEKiZHKM8d7en4uwZbMdMHmVmhgPKv2axGJ/lBzY03MW76Ezogj61MUn6OGcby+p71c
/xeJOutrWHghiRhmXh/FW9+YiLKIfKTtDDNDhMfAEd5HhHL+55yrHzuc6Xe4PkaanJSXwbOi2tXR
J5RaqUgiYCF42XMDr06K87WecBSESHEXTn3dBcTlMVGNrvbX013yVmqYSiEwZNS/MdeX99xsEaLU
sb6p8lxj7EOveKGIC8UHnxCBzCI/YwZymx4ueQE2e9NVjlPaj41jpo8bXjZsAwP3zn/OnYZ2iUE/
/z0rDqPyfboFZXW7KQzBfEK6tg4mjOA0aLxKykGKVerm9CHXWnjjKjZewx+mB7I50LcSbnTL10WY
u6Ea9Xy6cwtLB1yGh0Lu0Q0BJsBsgd/FiFUauNI5HIbrGleMuQZ/RRdmsiTyYtFX1NdMzivcjUw2
MxazgWejgBtdAd24FKJup3KTObM3DorBWs8XdSRGrKCwyDWZHdZAJJLVKfYdQO58TkN1M/M2VjLc
dn1c+UHQcBM2QCXch/OJUkur64mzC4tFlms/NrpguV0PVwBbPBHmYUmHwowiOeDCHBUDWz9PUpPH
5pyz/NRfdQ7de4Qhu8hVkrNxRkVTKW84AqwyuCwd6QeuPTTXCePkY3Qb8PYCzSXL3hXwsI5g4KPf
Q7T3yjkpXRvGf/Iy+l/FlTDV6sA9ku8zn9xv9Nbc5V9S4CWMzJaPYbJNd0o6L8ztCYiwTxHe8d+1
p/JhRC4TrAAl793VHdP+/CL3n6xd7aLW0JAL0+Habmt6YwbCGsz3j0JoD+fpaMPmvtVMHENhUcie
qJg6AkM67vXSxx/54VA/+f2TJZKeAyE33whjpiOZpQad43NTfu16lq6BVmqgbAIt9Ruer3bM2K8x
z6pLjl3BsCddhpmJhzY67usb8eL2e3mPdHSxbnpHVdvitYeJi5BFThvqdqSx1N3rKWO48dhiFF9/
2S0b04EDtufO/DkiAKgUwJQl531X6FZ6TBlzU/4knEuFmpGmQz1R/rbhGk65LdIi9+P5IK4NoV/E
WnOHeIZb+uVQb/+rtNIgy5SpfSMZyfKxWLzgUem8/9IlDvqLYtq2DAvy7Mt344NARhehfmomkMGJ
+t4v8JSy7s7OqbsxRpsfiSXGDqPiE/noEHFMkOpGMpi6KfM3gYc+2NFy0hH4ToD+YPjo+Lu7D3Uc
uMGv3lEGU6k3DMdHqP+5NtUA52+k3Jo7vkjt755i+jWgllWYJgXTSV0WbiDdSGrOjCB5zuX7i0Sh
/V46wNZHpH0oTFyzkQGyN/yEKQph9c2wrsAg/0edxylwRCJhowvlmjjsmehr2q2rM6WQGx6Mzr/6
TJpgZsbarZLmZKLBH9T4E02WMcKxnHKo6jG67oIvZupEdAYe7jpf1Lri48yCxygCf7i+GyLZhKZR
ZO9BSgjZy9rJ9EiSC0ViKaESz0lZuIH/gMpe80wfMvTVL8Q0QdIsnP1NvccMOO20BaDR7aU2mbdm
/0Zq+rMqSEwUfzaE66UuhyQwxhAre/qbL3fnT+OSKF0JUsHXUeBRd/3g/LQq/IUfR2p5x7/OlLuM
rBN+4U0dqrgnZKAe0H8kouLMUf8SEgtrITg8QlaqOi35YfDPWxyq7A4PgjYwgm85rnH3heNkeooJ
f4fsADEm7y+qRnGjAaB/PCYniXUCzux/UuCmwK010QzsnhjWIQdQ5Xgkct8BEAXNf3XHIiKE6hrj
w5LHqDG+qOEDZO8Y/o3wqJAtqiVfMgyqkxR3AngmDzapIVOeQ9vl+B+/lrEE6Nn1J2gW12+DibpF
XFkfE02+/JTSRs08yb7cixGj5+LjfHiDddhmGAfEGTC9rYn+K93ZaKJGYAi7NI8GnyLksrEzIvm5
1Zm8gOk2XEzXYxaq0xwy/icn5nHX+r11zF/dQN8iZ+0GbI32D8odXbR0K3swzPmkPh8/AyxF1D5l
Ye57khZHQvDcoZqdDuXQv7o2PGVfscnm6FDf3YZFAGfKPBGG2ShCUd6gc6Fh0Gd0Sn+UCTKBGudP
wWyO1O24FD6AlkeyuSklbDI08HqvWU+MqTo9AAzZlaTOqPMs9XbgKmTXwQ/fz3MHrujV/OiPVgcz
/Oe1xoGT7Ftxw48O2SRrdDwvOUFZrTDksLXcJRx3WlnHCvYAreQqK4uObI0PQriB0Bvnc842jcUq
sWCwS3cCCwyS9QXXYlfMhR/nXFXqUrvWXfCuxR7O6KVAnOL3EMOuRGi17CN7ObQ5LY/DKu3HBGkA
auK2Noj4TS2Gg7/Rlt/StXg0Msl6EWyEzswGltE7EMM2tFUX5UxVEnq6a5+9xXgT+jLf3TAbu3qA
msx9ZuB/3l/igZ3gXw58ikZ8O+2gJKxHUhZutTHrzvA+EYp31rYUF8AXJCCYgzeiNZV4PuJrYDoa
0kNcXBAeQa/aCFa0qYpWjehLNkiK+JeihUR/iIbsAoStmC0WpKy+n2JMoU89EmMxYZ8zkLVPKKAR
OZvwEV4SvfgKEiDOxejPYQUdOsfH6Im7ecoh4B7Zx0LzVc7MPLpLf2jFq61nJeIiaBCcpFB9y+MP
4WB+KoONxfSTURVNhea1p5MO1lEIVYnT4/0sYJcyed9+fIks7tvbb/VGjgHhKv8YnNKMSS2XPlGc
fSoA2wJsQGR3YTBr21h1pPMk59/nXqx623zl+jHkcnRPYRzokpkpTqhYZ+n3LUbf3b5TMZE/QTcZ
EUoe421BJXQ65gN4DBuWYDdqNqaMJv3wMCGvfkpqT/KWZns0xxooKLQYUDbPzDLt5Lud9mVsHg91
UNQG8VoOR4SGrUfRvnXn/BTbcBEeImyqk4VIA1x1zWQ3BnUV40gOIJczLyJpn5Jpni6CdWGWUQCj
1j40mCaLXdRs8o0t/17z4FKk4+5t04w4ol3igKjRvYWYuzku91rMNa56aANIX4VNRPImCD4pU3B6
wRly5NvpVRMnlnWgIKjqLutJ1OmJjwYDxfpetuF7tVU+RISS9lYSeb60IfLVOVg5wfi/cYhC7lLz
eDMhta9odCSnBe7OJA9o3wqT6LLM63MIC8YEnvxeTTcBujIYZWzS5sMnYiiRY9/6AWEmS/6wcEB8
HDmZOg7wJzVHDqWRRFFc7sLUo8KakKfN5sdMm1hHaHpdbd7UNHCppxEhTthQNJqJq93UC4z71e7E
/NC6NzBrtwmKU314FI6uoKhJQ/vHxCXj0NrixAJ3lWINoSL4ns13LGPPBpPD8OE2Nqk//i9PIw7h
6G7nf1ZGZ9IEXCL1A7xUQQMohXa1SnGHeujQpuShqCMWoLUhOBoSuD5dm7Ri3o+AmXLUuzqeMNGg
9BytkZg73SnQU3hgf7TWH6T73s44uY9UtBh0/b5ZxoVBPHWftzPArRaJRJI+AERhe2w6OD6jDulb
F7B1XshkShfLb0gzU1+4Yxoqiqm9K5yDZOl3zjaEg2Vg/uiQrtvS8fl7JJslu0e4vqYR1q+8piD9
P77rK+t08QpCesgxx4x37ZmXCKfY3DhStgVDuUv/fH/753L8v/aJb2rvgCIlYcKmcPtBXU4qh6wA
90di63op06I22kkaLZFEWqCopQadcmJDQEET7PLEvVm8rxIBWyEcuJ1mAeRK20zKNuZyvuAwr7L1
lwcmv5RO7qhlGG6qdAqYB8V4k7cahhsYdMYCP++jXROHA9ccKRVCetmZLaI44IFxfizzSP+2qN1Z
bb3QdhriDOiHXf4Jc1fu0Yf5Bj0sFCLnG9RyLtmjoxprqKhVLiKwF3GRyeYZqlEiTYbXOYUjN1zs
ClDF3fJ0w5rWA6FD+kxUPvYewdt8o33gucBi5hT/ukWxXFKPRzRcD6k4syIQlSHJFMLqbA2O+zo7
UEGr5sGZ7syMMQ92Yw0J9mCTih3hwidZ9qe8HdqOApjkIbO36mckdb7rSZSMiKmL3q5ZmeOAGQdP
HkXocN2X2Y4FWzcv1IZpUutbPwBgc5tdeP6Q9p5OjxqcW1YN5c27sdfHZnVzvC7AtC/o7mZWcICS
6/wgQ9N0J2RKxKcu5QPRDMLevYekKnpYWBqnWg9FHGA0JfeXRN7WTjTEg+n8JpzmYwDt6WZ5ZiEG
GRqU+1ME1l1x/+8F5XF1pod7gjFInHJgA4v+K3+kijSXnok3dbQvlZ3wxbGI4Un94xSzrv2NJThP
zjI9hQITb0WsZAFgOLqbsQeyHzsqH05haCO9CexVTUV01mzqurM2SwvCsw5+4t2WpK18CcRkJ0HL
PlHp4vxIh2QDKXQqOTXjRF8jh/0WMkHbgO5aw3EOrIIJDghZlF4EFWDTRmJPKh9R0rrLaWLf4FU2
4KZfLsOn2lVxcxG9J1y6FePwX/Q74RvYukwXWsylESWLgGM1+c+KZO9ND73c5vfP5GpMSOnjmztf
EdWTdIgvK3dT7fZgyM+vILT95NSKP/FsCZ2hX/PWzQveC2v1IS9laFbTxqhVZSJMwvPY1t+yY4r7
fWqlzKlg9RatoiZJdjzRNQpGz+aqcuIGaApTMexNm5R2vf32pdGZD+cPjqEogjzfgnrxpbyX1Oj1
70BUxJIh4EJeE8hnU7Y8oTQ3UU6o3VDp/hNRBwCefVq9GsUNEv8B2efiW0ww2ZBo6mzOplRJbcOY
KI/GqTlbBKjVM8R17MGL1I/KfTIN89yxMUDDXZ2j92EWGVbIPKa0rKDHjU6kWlqVsjC5fBNmbRC7
Hp0VcxW2VUQQmDML9V+v+lhFVKLcvs7w2WJ2DsayyQFBcuMJluCGhICnXpA9koVx+3a0QGTHthz4
oOrkBRLNE+cJyZ0bPEgoaxXLqVuhLZ3UotqigEO1+giltVPIw4OaxbVaifQ/1lDWDh4eJiv03L3/
2e0XqLL6zQIxkvA607QNrDQoPtqOFEX7hn0PYbcSWiE/PAbojXI3LkcXFMwv+08Iiwq58oKrL7h+
33rZaq2dCWuxsZgNdqhG4mm/NH8YExYw9c0n3KpYFRxdnyMNl9j1klsykhbjDN10hGorFJM3U/q9
CHnReVcFJjuZQkjp82QIzUfATJeqFUe5rSRczEajfZyLPoO/BL06nz3Z6eJU2oRY1SNPnH+xjnSv
bsCOFv8UhCzpD7b243RaqJuyD8on97JYSkDjGtMfRFHS+2KbAa63B4iwv/bER7f4MxuajporJxwy
aM6hOH1b1kdQe/lnn//5wNvRY5EnzCu063oVN5aV2QSHhD1DMvLGDgfyFyxCFkSxHJ74XLn83zqZ
AHrYWfbvQ2/GaIwgajTc4tQ1O78SxRvdXMOzQj2aWkCvIx5O7upL+4GmE6lPYkPsebVPqOlyJvaU
0Bx/g3Wkx0SaGt4qL6kDMU9tSC8SDEC5CjnjRfBp/zBPDWKuQp9Zq2DU3RDyewWA0IX/cc/gOLUx
4N9YrICwfCNJuqINBNpnnfnfcbfkuDC9X+SPQG05fJTyYK8EFQV7P9z+8x8efCzRmRI+pqZ5MRmm
p5pTSjSfZZpJv3S7rq+11uEyImeTbKGztrWfCQqZ5Vm24sh+YCTfgZO7jcK82tQ2xSvpyQuK8TBH
PSAY5kCeA4Kr/H8VaYNHM5VQsF9zOdTO2WWUdlrM2c2T7rMZRV65wuz98K5bbzv8PhkEED7mE4jO
YySwOcq+p9wyFIHsqpRrVDqU/PPFxr1kbVDU4aTLIXMg7nvIQV7Xx/vQ10Ub6T7kHvmpB6mPlPT6
a3azQxJpraTMGh0kE/mG22lf80m89BoDtjgAGgOPfDPZBiurac4zFo8oUTFQWd3S9/j7rQo1mHpM
6jxAGbVrCFDT75yQpIXYbv23Bclwl0aBf66kuhxDGrkRXTWpZc5ygyCU1PzQ9wfBsAMvP0ESGuNm
pxzaCz4YfyQs9oRG6pIDpSEVbRDRk8fEq5HYe9ecbgeSMsW//TPm3f36cG3ZrcUFjx70+nkhcYNa
3kVB60mAItT5jZwOD0RVdH1bU9by3LjqwMO1KidXjOev1DcbqfLTXfdHmwSbKRrTg8c8iev8hFob
AtJ8jXfrLHGUXZ8UFzqhE1DgGIyJ/muBcfCZgFGIaxeMsKQnmu9qhxfSdtk+xV4D0OCT+RbVQpdF
RXLMKS3dL2e5qOi2Z8bA5AyfeWIpeoTkOaHH2aH0RVft+y7xEKLnP2nlQqXMTBZKq5PM3KlxNang
2qLUqEmq4askATyP4mQA3WxV01bqdxF9peW5CJIrEA/O1Z2S1MJ+mRyVEp2tOHDNrfRG1Y8l1FvN
YkCX38vw6LZFgL/8y534gtbxpIUO6LCXgKWsIyNA0OkHG7vJVZE8Ccghvo8UT0082/IWyUsUn5sg
nUEyOqUGj4dlXJ3MbjXZIPTmsaMSGxSMv4C1sGwGoI9peN5VByJ05rEjdKrtruafg4YE+tkMxiff
wF+QPcC0T84Q7bSuCBG3tdFXNKSUKY9FzKQvUeDGRfCYxk//59tIUMcPShdaP2jROAoIeRHTrpQl
9wSBZxsQNjTZdlZcRhaXNvyRRjVTbtCWLQ3XoZXHw0w+Yw0Q+YGaCywNPqvxmStMFKY3q1PXdrYa
A9FRzGJjTvqcBWRUJ5RDZR8UhMzqtnzV5USRL28aiGGSK50zxW97wlVSpdYPavqCk5OLyVkmQBYp
9nqVxhbD4lOlqbp8bYneBWy+5OWT85jg+6w9UbcLYtXw0qen/x8MjWF/l3BqQ8eEycN28KJSFCo2
2rnXCuKGJ81S/ejIThdph9IYRj4Y2Cr57P3dX7TBHaC4SPp44J1FmZWtUCzGdKyIhrNsi49aNp+/
PoWvmXWSpjWgm3CBIz0ekKdgbXTm1PTmuKGLHbdzLUnzRVVF2i7ReQRXc57tvf6VeYHKv/ueT2DA
GmDlCBLc+x13HZJhAuhg0eywPmw7/RpPzXFEdF2CQy092Oepn2xo3UFW0bdH9YnzbGLyGBthll1K
1ZiaPF7x6s2u62neDTqgBXwXC/Ne/ZHj75iFjkro9BnylKnaYzCSnU15Qdf3f2fg12GzKsA5MfAP
8KOtwgVxeVJCJChaiXltY7De1nOZvE4g10K3bwcE+eX0mTJTr5qHHtX5iVIww4JPdNLlBtszWGaH
DUs56f2+peM/TqrvRHcfr2fIkAAwrakLdzPFGZVG2g/nGCnb6bXqCv0j3mAWRdnp8UKLB7V3mrwW
Dg1+Im+o6tB5QjY3N01MA3uVRFFwfcXT/wBqQK94OmWqnBOW8B9RZEpAGoQJ3CteW9AOlwkQ54ox
FsysaqLr1UPL06dReXzF2dX51WxtFTVSga8ws9n0g2cQovMTQl5ae3KE20hP1zH8cwP4Fyc9k18+
tX0WRJuejY0tNczy/dOepp+1H5LXYqST1bG6n1rtUxrOIvJMlDZ+MreN+Ou7zJcnZSOh3IF1Pqi0
3pMZNaMgs3SwIM0j/Xhg5PLIcJKX0mEWFIjXGrRJa/eZzjn3J3ohiALBvpygM+PY5LajLehNElEN
7wBLzgEmwR4lPf4mx4HcezUmrCg3XoULPToGl1OPmjfUV2b7rdvj7NXf36qHUwGsqVuQNEHQQU/9
/U+wkhwHfBwTjRm3qJk6zWszouYzC6R1lxY+zPpHgqwqqbSIlm80r/IdUAG7pqCHVJKgeCWk5PCU
S+IZ5txRAUptY1N06Nouv2wjEEgc558geOIT3BbMhvWhX8AsU2O9uwfEL7/Fv8256l8OWj6o+ZDf
m32jh54JIU7m+M6LBO50ZhqzQpWqJ0wtn6Tt6sBATweCprCaU5gm2P1uylL+vncGtL/KeG9Ngnih
zYx8SUyFd1AqJ+iaoLlFSsUJlTLtVoAWqt99Rx/bSEMxnST+G1nnWTbtHfHiQs0i0463bgwNbI+0
KV5qW1CgESu9FZ7WYqTinQJB714da7Jc11S1W0Vj9o9DmQdQmvKjumXrVJ74k3B0W3B4S+vtQeSF
miPNKUlf8l6HYaoIcR695afjQ4dvcVb7UVkTVED8oJhO4WfGOM1yTg7MWDE83bZ0P8P/pXl4PDA7
tQnAdFTg2uVX1QL58ym4fHdFmh1c+rVT+nrLOrb83EBhKW0xAE4V4unvmGZ01VAbddO5Mi+H3NPe
1vr9c7xJhsqV+L859qZ/1ou0rZOs+57BfRPRbgflJNFTrtQjkd7w8TqD1pPYW09Bgo97xpU+ypqJ
elBw2I9leeFmFhTLSQPTtrccOSOHhr2iGku4UQBoP8kjE3/klHpDw00szkYOb7Z3nb9jlTIUMoSJ
FaUNCfgq1ktwLNPB/WsU1mWju3v55raRUF5KQ3XlsBKvgvTCTRh2RmX/fwwQwwahR3BNu0cUUlw5
fZKcRc0hXQ1WQENtdVaG790iGII+opCtafYvBSM/7Eu7ThJqdmKbnkGtjD71e/a4GnTBbqVUb7hD
8+vt+ZeK1YbAeGSMtU3JJM0BKZ2jRxmZThuMdgKJAEajVIr+INE7uYYp73qFTPEdKCCjLYFUWh5e
kcLtv6bByLLoUCGI+qMqSuq0h5CZE0fGkPZUB9wUhkP5K/X0U+OifF3o/XRbre938vtB1wbfor14
I8rjT+YMDKX/y9ldE7lofKOAuJ7veU4IEt0gTpyDPCmKKbKbRjojAt+jfCH1WiJ+3QfaemLGpVPO
4tdCEEpz38xK8Zyw+1cN8wKdUaiWD06yj/cjTKMRSm27/NLS5clGV2ExAeXJkXG2knXM6boIEepy
5QOptoFtKYD4YmqoBL21rdE1NJPVtr6hbRPAW8Vx74C6A1Pj+EQmDuCLWEOvv/kfE1MUekKEH5Pw
mOOav0QoGkafsbioJlKSs81p+8MvS5L98ciOC4c7nI23OoG2hNhQvedEovKSjOZWfYfoewr5n3EL
zyhtMre9IECyJdvcm5ZfzhD6tDSir/YbUK9ya73EsikOspHWD7PzeBL2p1KxvZF48nuA4ZQsAL1H
QxZnHdhifTEf/QSwJWFCtuSZb7Y/r7ClDXGspt71SEqngb+FnxX/7zwnwqZAJmQlWQxBkg7l7xMf
3hqZZglw8GK0TIWoGe7GEL6bmmfGZyHG3CxTgqJlTsKPF2qEIv2Ovv53HL8NGtypdwGPrRJ35i2m
BqSk5hWBilU6i/9pNLj/Cgi8u0afPpnP2Cs6AMdcBHjhuFzQesbnp0BtQnpJLZ2P2YOiYWfeTQ8g
cbgc/y8YpV117yGI0UzyvR/34AVZBrBP0oSDQU5hj8vjQZMxiTd/KZfjxo/wWKC4cqBN5M33qEVT
v+I9I7sPVJ4vRTTdQ1YtZIhrPd9CWpS4RLsBOec8ftMmrHCuRx0v7ZMpE1aqDZMpsbdykY9XQHRx
HFsgcMn7ThUl6s1RyoeRmkuYTW8kTK3GG3bfD1ti1mHKToEdBXo8WhNABwgb9+4bx2utLoTLc5mE
jsYol1+cl00b9dS/EjnVw/6k2pNG7EvvoFHiS4Lhl56VnbklN9sN7gyq25zA6QCHMT7JyZxl+89A
JGLhKPybPbTjoymXG1VfR/QWk+hVAXEwVycOqb7eSjbfgQQXaOr9J94eL1LoUU1jfA2P7VTC7O63
gvtpq6mReSkPPECnkg3ZMcDSA4P/NOQ0IXuwtjJBU3Rcq+UZESoMr8obmA+JZZ8CO2nUDEcUAQ4y
3Wexs04YNPn+/wbIfUY3UqSjJqOusnmY60KBWL7l5Jvy4HgNRp2zFZQQlrfQuHG5QxpSEIikODQ/
MWLR+1OkP8tWMM/44pzSrTsw9YaEA0LALb3SZMm6A8CZ2YFkuatxuiu/BR/JZg2hrBsV50uq/SMP
w3TKJP0NL81w1dYnvvJwHIMkgomy+Uo3MlGuFI1EdkJyX5cSQiVKXrMGvKMQ2GHyuEbHH40ULNFg
+1jqazMlXmoM2n31nc23cBZZYUKE2falLsUUScJ/IglN8cy9gYoYOqPREYd4rJXUF1g5dHQ4Egc6
egvNJzd1MObtB6zKRtCiQYZaWJKBFs2509EiJOPl2QSjTeo4R1TF9R1NN15rQhR3uhmAAI0icqoG
kyw7B68O9vyfZqqzB+xKQxHvLCXevVP4JbPikPm1RisvX4nzry4V23BzwRTZOMqFMNNXfbbpchVr
+e+b3eXMvoo40/VnjeFwt3eX8+yeropgaWk+yos6dxo6lYcdFRYMzpbP4lHM8afkaMvzFPtjZ8kb
l5ODCQC01XoBkdzWsO8ZEKpH13FD0lVW784ltHA20WgbhNmoEaM4Vxd7SoDjz24jhq8mg2KfYqi0
KCAo54kDYs1TDzuFVzQHRrfewc26giokEUTN92elvqtPKWQFZmW41UJlPO9xmH0EclrHcHqaBT7/
QHTdyPsQjGfltMO8YEDPjfo6OLHqMLi+1MF6Uf0zqyHzCvFKMgNQasygxbcFOgC/NjTecaDTDp8j
vAIoBNwK6cZllqDOI6heVv1vGSn/J0QkQL8H/uI/dgFhwClB9YcM3rXVE86XM4m3AaLpeqyXJ0i4
j3sPhK89KjF/bOIC
`protect end_protected

