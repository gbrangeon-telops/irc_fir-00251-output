

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Hz4PNZqDQYlRQ+ken68CUlKtwl5bD3KVcGYwK7pLDyYBwi6Th9L/PQr7ts5tJoXAIQRYcIzRxOvE
bOvIjO60PA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GP7r+Hw/Nq0CwA10fCvNkrkcgK45iHUPRmPqoCkPDKd3ozfduaGFS4NbQcQDFEPry0eRmQ2gSn3i
AGkmBiS/ZMkSitJxD/EIgYbO/fqPeNo/xyESKAW2O+T1ZwGwXyv6qMAp2gFqycRAbj6T5U/FUq52
EYpn3NB0sMc8yOEFyQo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
le8HFUmlytAxiraEF0H5rT3qqsng3b8xZZHcvlli3mx0SdV7s39NBBuklCsi2z+U5UKSzgnk8WIo
w7XOgbkBH4I5bMmtC280eEWQOIcj1GSezKn8Kq725OUTUl7WIOM9hdaAEgsyYV4aegR9ufM3pfv5
jM49vFUeG7XEd7xqdKUxYcrZmsZ8CqQuOZKMv7+xnku0k9eaKv42hAQ7cL1uIXuIFvzDlZHyC8MD
e2+jTkJtzyJMk7U2Hncf7jaM/O2gSIFGoRR2sNNwVB0ATLYzGBnoP+wY1MWKJdSoIbDQ5r0792eb
YO5yRbe6PhUe2+UdG6sNzgiR0viGJQ6R/9i02A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tSJEOPsqlnARL2Dz0wpm4XWyg0nGSs+Wnp+fpstkJG7juRdPH6snLi4H3YFLGcOIteaUd6+0+nV0
HNDEDrgudSIwom4ffSyyotXElk+U/5goIr091+0B19LyBlVHPMfovruJJsH5yPOjkIUbE3z//OG/
9D90RTj2hDW4+5DRikw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y2U+pnaPqDjEYN9Ag4nM7UfxJ44UWPvMFi6W/IpytPtcFc+Gta7bvyNellM8zINHBtaT4/XvwpGs
zz9LduYm/i37u/eaLh4notjKL1KlEzSl/RQQCOAWEkJvBF59EPqbeUalx4NMTEi6gApYczcwU5ry
jjndsvqks3Obkc3R6uXlQHIzKbPFQM2kj8SV74srGUscAjTY98txOVHFhIk/okWPW2x7ScPBZlnH
/p6enNTFgNVy7YICPLQQ9SjExe9hKly0/QrbtcXPdI2+m7HVD28iWrn6JNqPDPmkYTv4lqGhGruw
jT2AigpLW8vV0cP+HITHbLQV7l7eN+9WNmGRNA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 126368)
`protect data_block
glmcLJybTKQYw2NbsLWCBo9jY1hA365q2m3mPWaWe3buTyjER3nmaal33KnIcieCaigOuVJaaUIf
d5RxDGaA8BI11XbOYX1laetDlEGVUy8q2bC5MYmnJoMBts6SCvBch1I15X4WQbBnbeKGLUTY4Gx1
gTc9T537TK7znz36CSgzIj8r2OKKMSuFlXWUNkSSw66uMIn2N1076Zt+nSSn6xY7Afnu0f6kjPGj
HzW8KM2oknHGVcLCHvd9cCm1zEJfqbhLS+v5FYu7Dbb8W/wA5YpkSnRt9NXCXGfImfUqIcErNKgJ
YZQH1I17cvB3S1g3zrmJOGl6Bpsl2iDq/qh/o3QAtDuOtJEHnIHQqLDDLFx3AyKHQy1ecw0T2DOp
hHDAp3/YkeNo61aLUCCPNm4+tSg0/Dq4xZDDlWwTEjMF5dJ15JCgKkP7NJ+9hd+6XVFQ4QDECEDa
SaBmcxntBPVP+iDEE/O7T05Opcq9oz502YbvANomKsap2tx3iNt3CUe1osjFZKyXwtZuQwANzObo
P2C7vGn4oJP5DHjh6sB7Sz9SRtzqZPxQwODPxfip2Wz+MU3mAhueJUqWQ2LblekTBFe+sNH969SZ
AmK48XPXkSZIit3UMa5/gmNDtfjoyI1oZDHIw2qcjnnZNBtG9gGGrQ8VUx9Zkbxz5MIzfN6gqGY3
NIAt9koBCmtAAqF7Z/cVLpOVBe1n0VkmMPc/w3OwiT84ZcuROVQavfZL53lED0vXOUvRICrs1TQj
OxY2zQjAzoeyoIKZnor6xy0rBGsGToTtC4upxT2DKDMQenpBuVgvGcD2zNwRv2T/XU5ZRE1qPE8M
puKeJeUzyCdIdfpgxhl/PibyMiJgnqQlhqxq2IPpusEugaa7pt0troSiAqRkKPaFYNODswZOMBME
BsMUprFDqlD9zsIA1RAA0M4YjXOrzSFYAAg6htX2X6OlBl0Ums7fxyReLNfxObp3m1KardT4SCbG
mg/ssXSQV+65rqIu9NQch7fE0W7xESuK6Xu+wxDHFn14p9k+s4RPjtsD18ICWEwSsZGZye1adWj8
63ujwW/HMj+0BCitzj6fRu7SZ25hV6DwqVhUgIL8A1k817Md6Kr375jFa/5m42H+Te3/k5eAsqTn
GkPYQNvTE840ywiYFIO5nAC5qF+mVDVMGbgdu5EgH0k6OMISxcFPF6+jaqXi+1JAWvmJnQ48zZRw
4LstLuxve2axR5lEFZ2/VJAU9MXb9uNHEeRgwZwhPuAYN1mk/yBZZIf9IWqRs4z5Q26h4p6KdNFy
GJspDYBvxdrHjXE8YWDenP2cohJmgOGVLlG/L8dv3DYrBuj1+veWIypyzO6S7DDRyz3eAZY/I/It
nr5InnNzZqtwJtt7HsO65Gm2jtFvX3ONI2TGNuUftRQNF+ETxQ8Zs5hSaJk5E3CwcWoYOXOaD5IH
3Vf5pzaW3VHyXPbQTBPBLOp0ccd3M4OwVNt/t8eFY0ekxB5d6fF/Rssl9cx+B6Fgic8ejzF9McLK
1uPzj5CbxtL3dfU/mT5jZwT/jyJEKhoGF37M6fnybX3WEzJMQa6KIwOF63KHSMFYs3iSyBdLu42E
NTrQpH7g+NT+MVQov4gtUCSBFuZyWWIWrhbGL0c1syx9t1i/xfWk1v2YpYiU0uFaW6/LZCPxGgRL
xUeHn7QbR6hJZ+yymA/Xq5wquMu2Z1PuPv+clrhNAyT6NRZE/O34GS1i9Gc8n+nxA7AI5jGjtfPU
BF3N5TLKrAyIDaabkXeojkATpxIAgosf9g6Nj+I/+/VQq4wZvhMdgD61gDBNBVCqFlpNIFyZ60qF
+UdwNFYXnI5D6IfpSlCq6wwORS7JYhkDE2XuAAvUJLjfJcDToXvUVS3SsV80/NZM0s4Pv8nX/PvY
H0PPY0jv2wtuLQjP8KbokDZWt5K0zMRar2Um5VL7NRK7m7/0oB9n1+nG6kTaeHLpKpvtLH7n/HUd
RIUIBr43PrgCmsIasd1wNS2Q7O51C1+zL3cCFDoJTJrnY8P1GcfkMlncxjyGI6JGt5gtrVQr5mcB
/l1w3BzC6vH4jQ6LmncZxiUbV5IZHFo9r/zDuKkcTb2in1Qae9aiXhmnSykCrOWG8UeDjVCJh+iO
6TX24iGprOdlR/cqGtZTXJT6Pjlk1x6RaRBpXasLOiJYtdNoQQO2KOtBk5kw4NwZDrwzyMGGTqkH
/gokNzxfN2ynp8S/3tGE9qBjRD92p/68iMdLI2/5FMOkk5u1r1ObJAno924KRVQxAt1xMfKh1Kju
QqtVUQ1D42I1bbp3UEFg2TVbvJhoXe93pquvbGxb4saOcfkFdizVUmSRcA3Krb6cvdROuriXV1Ht
JE/tvle6Y5OMkQFOvZcr1EgXhz+MGxRrk7D8cdImT1ab0sak2jQYarwMPUTFhwfrM674CA7nSi4X
x5bjEwHFi4Hx7EINI2UbjmDdm1M1tRPa2VrdMGc/5Nh8DTDwwFwN7cqTWzHUfEB8YvVPak7g1VC+
g/jd2Mg6A/kPsok4Vz0C/IAcmLkT8GK0XNcrx6bxdP8twxt7o5r19D3CK5J+BNfnqYfai4+JlUV+
sl5saPqpCdpUU7TZWRPZ2zlALWxI+Kpev/+gKT54w3YVy6c66KVVOBeVO2ny9Rw08SiFMR5RO6Em
up1dONcQOlfpWYqRpJ35MSzzF2JKYX3iwCfl1IMiLgjIVP6kwKw0BbuH510dZC1lVVOBd0kUQNPE
lMFHIS/bCjlH4hxCCYBAtLvBX4U71VzjuEZAIoS5W/WzLUlMd73K83ofM2PVpsk6Ya+aki1dkJg2
zBDe0FNa8KdbZk29yGnGWFa2nZMLJSZAQn2aeXppj99wOnduxxuHjhoOToUFDaNPdoWmdso56U7g
z5wqRJie7pQHUrCpcwSviGfX0uIbZgXMvJDn/T8VcAA43+CG+woWfTM4ZDfl8jlmaJGOCVKEacLN
GJNd+famDmlBt18mBgZFDSnoPcPQmUq/76qpz3sIRA1jEe5ICQcdrLm52AKnJrfpo9v7E7vL5ltM
ZTzCGHPSRRgRpBkuimpgQACgiP05fLg+5JEK3FqrJBTU32ewTpqUCazqQhw7wveUhertaacNk5Q4
Eh6G4EoHnGBpsCRkIe4+1tTM44IpKQJijqkap3nFeZbP/ysZecikQ7wz3Tw6oqqlJaqXxSFZ+VJu
aynKHRPqYD7SfIAxQaLBjCBLR2bVmUcmyej6L/4QcqPDnpak66LrJZaUm9ZDfzgbq6ck7xa9TLlK
NTlPJekmmyLh74zIryJjGwlhgBRXQqnTPiC/VAPFwF6TLKM3P8bdCQFABw4Wt5N8gh6QIYK+37ce
Lr+BfETfAlFqWFHip7gN9YS6xmu5Xcpy9RMt2j5gpitRHHeUwRvoFNEpxnE3/NJnH1PZSfbIhhTh
GRX20zqmQ4wxeVb+zBurthfk0s655Y3CjNG6XuYwYHmW50potoPfxMZxYEdg9GWr7CCiaiPXaWqH
o6CCSlf0DsYyYo/BZ6Z99yHAmVJ2UmkoKq+qBuDlrCN0OKYF1ENARVvPWRiWGaBkeS91KrMQHqS0
2YoFCAMO/KfbNVhvA74FKZ8+PpY30M+SHkzCO8SywbTkG3VhzDQfjIv3jqefCnN7F0zRum9PWnEZ
VDZCq4PYoHYBYoMRLdru7jE/FlCHP53KlnEnnC6TKJ8XsIjS2Jw12wcM697VazKspm7/5spsMufY
12MNGRmCL/yJYcSpirl/SOgovZ/DKFITCYWDQxEEDbXXdcAEzogfFjgUQMKczf0OpNgTWjh0o/lG
4YDMAGUMcTslnKHhWHlh9JL83usJ28F9+viwqNcnrhc8T6H+VPojc1sXFoprp1dIshVQFXoY8UQo
4xbeKtZ9/ZIuFR6HZH/dB4Q6pXjVZCMzWWsa9KcCgyCafasQqkTCYxKl3hyOAZU2Xuz9S9C88PfH
l0+z4h225AalPevIxvDHYzNQUSwaz3IEHtmAe2OZzMDAvYeEOX6Jk+mVylalePDmMEPKyw3k2Afb
Fpq0XqQfBkw4zgijsE7/Nudx0Ia2jmOdJjHc48dCrb6SGRHFcvQJnbgDUXOSCzvrRezSvY2mflQE
SsI8HoOBTbhh7PN1AjDGkfIkRpXRAJ1OmjJsuwtWjA2+gGsSjH7xC9lykyAPANr4IAs4+rUDvcqm
81IW5bHr6fG60yqi+lRe3+1hKFAXTgo4bl4B409qQ6hL93wMDCBpc00c5rNUbYRumzAs3/Wgt0wA
LQN3s6VmNDZOWWfvvoIXKGNC+5kq+Gvqu+DBjVOCwCtcBbugTY/ssktqIAgMW4i/sB3gyOi714u2
JACxq7vyud0GvDJoqZr4rn9PEMTWxSn3vu1vhlEsmf31ftelxlJF+7Ft1W+ERHofOi2yBmY5nKqP
5qaheRz3dqRAFmgZ2kQEjjxnVLFn5e67wGwX+V8nw2wPvRtJkuV8sCSjYbrhYRYANJYB8Reia3lZ
2CINrf5ZFYcnWNr4EINYDjBwlXbKTjSmtcYrDpi+egOhXo2rv+zRd35cZqsXlu0s+UdzEi9opN6a
XssvPPbK2XmKcdOlBU+VI2cpwLsdtIN7aSkcHHNuKe+IEVl8qP3sUsNpOyyB0txL929+/Ds0p/X7
BOKDIlzKca4o1Wvc0bereiBZtSNX74N9s+HmXS2UtgmGb3RAUdtqFyma60nCfP3DnhwcOjD+xZCr
GnbAIjvHhYUyZRKarBknUXuU6y55CDMi03ghX9QIb7vqdzJWkxjsG0UzYYvdLRjQhjq07Daub43n
hj+K9T27fzFdRDup9QkKC8ao7t0iARMiv4UYLRFNvIV4TzeFWPDJRuCIfxsXUQHl5AYPyaLEKPEC
z+3oum4RbK+RdjKkxcungQNKhhG7ydIs0NieSC7hAavTi8vdYuoYrrgT1ISzw6Y5fmKpGpUKPFth
MNQy0h7tygsR0vmOg271qpoBRQVcJOGZ23Muc68/DPi5nev/B8yIic6RuQBFaZpm85QblHaWbXzw
SzUUPz9hnkw//EcClA1cWwizWRsy9yH7yctBR5sQvCvFPEZqMT2SJKwApbA8e/0YmY5cXxo4Hrke
T9bpDGr9ppiclIvDhYjPfHogzHoM4z/GMcKV2lnFiirMK7Cu/6SmHyz1SnxkiXTFYOZ1sVxhexK4
SsElbCQqvbLBNAHR57vdAdTHRh8/vUp/qXjOcBjI0uszxS2Ta2ZSRMjgtXF4pkomGOMQbZ8+i52x
2WVhqLmvwIj0qG8J7C/o6FD127tABNg1gP9YjHR0trRdFmcdGEhJGH1E9DwWW/PzQiKICh72Q/tC
rZPA3taOlq8jd7GmsD/Aqln1jthgu/4TE2SEJFVUil+muNTXjquQqWhi5E12HONfr1w4r/4eFBAH
isDmxNx4klAzx4Z+Ea8UUqmsgUlMevE8hQ4Bwrxy54YicwJPtEUeTYLe8r2BT0eQ6SA+osG/R7hy
UMD54fU/2620ugTGjnVtO7MOXCU4WYhp2ij6RNfBFXw8xwNJ7TKeSSHtZhMBJE1BpwfBtdsJWwnG
uzJ3qzJ+9zgOlX2Qap52nBgHDlmy4Ngg+JiRL1QWa0iUllqlDqk+2ALazx8wnh8Rlb6b5Qq1Z8xD
1IGlGWyqMbJ1P3R7Xuv2c+SLaTA/lIm1X2XrYKAInCM93WlL7jSBUDevJOIbrqhW2vfzw8SD6BjR
vzYkSmBpqmvy6HhEytAMOjQUeiAPoINvW8KTrlVfkRMDEnO6C7ctsMV9MVpmvGQi+XQcQAKuOkku
TIe+YQXKUZAjcvPN50DjNosbXHssbOKMNItiN8oBIXU4v81l3zc1KoOMMG6yR8Nu02ihAuWn5Ff4
WMnkt259w5/P3VEkjk3rU2+zgx4d82g5LiY86iP0dY8wJKsUwnZoIRtflUaKrUeA+dpKmuXx2tt8
j5gX7i5wwmNfW1YofliAQWMfb/JdzWtA+XTvzlAaT/kdxRJoux38o5DH4bvHP26d9BnppJOWMCC8
J9Bo0BzxT0D1ryHirmDxmJpjj8GJuLBVa7jGt8EpYMcLUPhRkLig4TiznHJM5nVO65XEwH68IN+g
3LVeMuNMdx598lv25RqnHV5zU0n+manIngAwB98skDp+AVoxLYWVcPVb6SfSyPZHv93XOCzYUfoY
ZRxqu8MqwE/FjWE0JUurzWCYEPZruWka8SCkmRwme31xCJSn12pOuGYm/sOBsZNexWBwcu+F/vMC
Z8ADs0RXv1eMmZSIZzWqTRgclK/jOEGXBuRyXgaNMnVOxWC6g9vU+DLycQS7P/HG5TH4znq/oXAL
3aT6WmEKLtuQNBs9AmTd3hdNlEekSUPKVFRlWoHfLAG40+oi0rsxwD3cILbcE1FyLy4H8WfplHz6
i1gY7wkHfUiw1OuBaXTctDFPvLmvX9hlnebGycv9lv2x4bbVL7lG0fB6a63pJ30Rz3y3RFjts5Cb
FLgamsONmdnKkHv5t9YAhp4SxEvGCuItMH+D64VXqEP2SStk+Utbxo+ZCvI2Yx9LypZnnpGG7EfH
Re2d3cOfiMeeIUeQB1Lo6wduwDh17xfFiNl1vqfkUhAeHN8w3wLYEbKruZRJ4X+Sdzc3rArITThU
O7gGHfG6N+6jHDVjP7tDCyq0uCdFXM4TC4WNwIhwEt+lxuai6wpjAX/X8f8pgvum47ZsmVwI/RHr
36TIwQc5dGyVXy9ZD/D+DfdL2EscWXKfOgjvXdqFNqW626uw1+5Y/e/ikCx3znPPz9u5jhN8M0lK
nvAHTu4L6JPOhLwv1/+S5SP61HCEfZQsn3JXp82iNr1n03tC84S8WFC8WvBODuPEr3HL1sF5qRtM
QiMg29fJNOXnxIbNwW1noYHsf9RwMEHlzNEKfZzHFmrghs6GvEWQ9oJpmlI4tXReQq+0Y0ANqaUt
AxNZZgtU+BtCu8bPQ3UAtMHOW6zK70lgZ1oCoIIiGbnk3jrGSbN702Os+PxsE2SUCXIos5WgSfrZ
kar8CU8i6um1pMzOkIWVPcIdM0WmTO0VMx5RKRt8gf3ktvSAyhv24sNDh+gD3D97Nc6MOioIQVn9
e4ZW0s0QnA4F3izhOTG1azrILvGYjqOjlh+cI2K20AJMU1FOBffHbVlOd7hPkZh5jYR4DxfDc5oP
4kgXS1T8wbN+UrlDnmtMyc4b1ed9ovkSM4zBZU8MU9YWRUrKpE+7hMO80L/stfDILcFfgXwuDQmW
/PysTkY3OV3FjRDE91A4e0V7K4C5YPynjrbNxccZYa4STdFijcd2BKGb6mTTJkFS2B4CUUiuvUNI
QNJpgV+4QhSeB4P59K3yajFvvTj/Rvh3phoDNnsSVvBAEAXwQJOY3i1J016HdVE+T+KBpYXty/zi
r61taAJM8hcj0OY7nKxJRB+QmaZk6Hp5AGeSeL8sc4wq8vfpnnqp7AwnZ26Rf8x0JRhydWJ1LeP1
nHOOifXU649JqSHfXyOm040TlWwdvqfo8NdmQSrV3NB6V18TMJB+O/nN+Sctoh9t7A6sKoqhAtpV
un6xsqQfS3/c9/j2LCjJaRh4csJMpwVItLoGQeBg9xTKDGxN4dDDgztCFFPN2xJLFWUJ09a76JtF
QTmmkRxNwgllLArdKQ29Bpevo5FeE0jjECZvtOmMQifb4LHz3GKjZWU4+ChaWmxJbkkUSHDUHvDG
us4DqHH18IUz1HiOKfoue/v5UfONF7F2f/K2WSF1MD2ELZ+OMICUSOtPnBolQ1Iv3NcOHIkV6v+3
+D7OFJYvtWbU+r4EzFfArJ5wXby8jo+yZeQo/1NP42U5uXuvIta4gqbgTA3qQRAoQlVn2V0naAfj
2DMqgMkTURrdl8h8jQkiixLFvyAxxsPbe/eq7npATD/YXYVvsqUWiJ3HI3zjCTnrVY9obTc9u2+l
PggyaFLpyeRSrA0KWLBr8rU+IpqaI9uuDiuXBLDPtmCredbT2F37mxgx749Ga7u09RA+V1Ly8Dsi
/Q8PuCjb2DmRsQ5r8blR4oifHzEFxNKXBVIa/uyV72kZ7PWcB62oxbnHhCz12uFP2u6/0sM3u2PS
NOtbiIDAy/Y/hVjAmqXHjZr0MApdJRuAO3i5dHEgE+Qn/iYMWKiKBNPRfgejY007byESfjvonRl8
t+46Mt/TiuCZZBCcec7t5y6qoh5UJ8Kkz+TINZWlCuTfWZ5QUV1F4zeCedo0mE9S67gNFJayHKYA
dytciYd0FcpdlBDVdRc+Sipsjf7Zyn4JfM1gima/R/AakUaOp1QKhHZDk/GpvO5w756f0FAqOszE
VITidr7Hs+yhj3DD9/eq+BNgpVAXWeCeAj9Tf7xaW3G5KpJ5Nt9ah5kbRlVNeg2WntaeqKPUCW3+
10X+C5ZzPXGkC8NMhzJQXplsf9IZdKikRZQaNkH0qEBQRd7PKPHPQ5Qc0b9dN0gCucMV9yzx6Z4+
alhXms6weKTWPiKhFcJBcxyzGLbSpe1yB/5l28lKIpH4EMOm7POHZ56qT25U70p8PhB0E3ecdyva
FhKlkj8Vy4LKq+Z/rKKBN9fYnTY0kYIMAUOgLI05rDGRMK2Yp4N2OFsnPIbfjHXuTk8zD2oTI6QL
pqFF6lLXxvXRNg0iSQJ8Ra2ZT1PrtvZLqhc0yhkhHc7Ay+1PnJn35W7ULGoj5QL8YjetdprnWLYF
+XIiB7x+eHaL8IofoAjACsXOwgyWnIBz4Se4W/m6/IXeYEdUYQkA+QnaJ757AJizw5v4zKKto7eP
SqJMqGOt91PEsJQpqrjitiVFIM/hXFa7lVGfsRSIQMcEi2BmyC6J+h7MMOe2tkXbEvH+aVKsL1mY
XtG8sm1D7FfZhkPgyLbM5fd8EeEIT+IjyO1EsDX0MuQTqXNAfduKNKrUQUB6hYC2A136CQTs4vwP
Q9E+NUZ0kQ6/oU8hsHJTyitNSyW7csqqhwGx3fm88neSoPPZ9HsXN8sdxznWCFvMjfDBZ0+RvsoO
lAufvj2h3Z3oF9ClKAdzXMqexK1R9p7o6Ead/yYGI8tLXSvwcsGdSvScYaPzohQ75gQr/7Es7W6B
vmdEmHLvsD/nHxpYseEoNBVqNVHG3GfkYqM6rk3DQNoejjzjx+47BpVdsUPsk/w+BFw11hJ8SvGY
FEJ2HUFqT3kmO7tvgT9YYBiQXsKGUR5P1/CjeN8O0tl5FmfqlB0g9802WiJsJ9Xb2ojspZGYafSU
4J+vFQdULI+DVu1er9/zjzqCmnBoEcmjY3GoDa4b5DUeueS+pAi2l7AIdWni+LaJFbyqNS2WV99f
oOr6cJl1mXHyiyib1agz4WAqyJ20IpHrc73sttPmnDdSOmBlrGj+6oB3mtqDs4oRJMsmKbj2j3XP
g+nwtlD0r2Y8Qy+Fz7c4bLA6+aQXjCmSqmCXUeGKFGbViVUNZPdFSMoRN4cfxILwy81snDCPN8OP
Rirrf0sZoE7AO0e+AspEcHszL1ZXi3joAUgv7tanteRSUQAi7Fn1kClxEvFQQTRpsa5EffZVlhRF
t4hv3S48Uv5EveksV3jR17sCyAMvw6BSbqdP8b/P9E92PfjD1YGOQt+MC4+asOP4PeIkUD32WuNw
OVyzMS+mdOq81IS6NHNPuqcJbmZhPqw9nEjSgMQj9f7Xq4GU3wVR8V1xhMYcSd2y+m/K9J482Tn6
M3li3CWIdTXGu6LVdt8knD+DWXKSMksorxo/aSHuB98otmexMT2FyuY0ALw/UelZDhRByNqyLgwL
XE9TNWBAhW7BtqPbBeSdGI4ptS7/rvd7aFjP/tIqMcxeOw3D0opOSbb+S7lxO9pU3kcZ9K5XPP0s
SjmMwxkn0Pl3DTq0ZPNcWb/ldJXxa+QPqYdCm/7Bt3iCNw+Gue6zujVf7OXb6iEP2QR3F0oaol7l
ozAnj8HRosTZnBMdPZVFTLMMp8tcfPbWae6bu1fa88vZEXKAAP8kc3oY1UU/OOhnNme/TT1pR/RN
dF8UrPYiMu46X5UZlQOENYddg3zXks2AdvKTT3H66mM+AfBTJD0qRS4wJ5/ZRXQNvhTlc3fC3n+N
Zur2EciwjDeusY1AyLEDRyh1tBtoavBjgMKm7Z94QyUL6cOV5bPsMiDMZ23ifuxRDVUcX0Z3Z7uo
w5J+ziFqkJ07dgh7wie3OGcgUt+W8tqaVtBlkGAY+u9VDvUJRKVLR0COglpxvOXRXg4BqncKtf3d
66F+C87m8rRJaWMjgGiJ/2cCUynohFfSjHT8qO39NcIsLr39SkAB9WmCyxerNAmpjmBaurZy3qy/
CP1NkYgtRVWDJc36awzHOOjFRdsZ3pbI8B8uK05BOUfspK8j4zMYUBazKFIX+7Yuk/NGse+foX/9
7NDK2NJasICiyvAjPmt1L2UmvaVqr3AjbRcc99b9OTVRi4A+Ch4mtr2Bc7mc3r/klLib4ChnjdxF
ZeMoZTpq4HqX+Tibm4Bc73ALb2pR6kh3W4fL9U1lHdVjTyppODx4u7xFbJM9PqslZZQwIwsOtBPx
46302GaER/T5gGh8oBuaqE4nVjRLhQ0V50fW9TAuAvDWbkHr7MAOU1cTU2uVc7JpEp3DtNFOTrLL
68Tp4LKbjmYDR8vVLvAF1WR6XvPNr++4LorlwEmfFaYuRr2ATPuwVMgtbl9U/vmZzwbbBdsQyeYk
ldZvjTr4mo48iTf7Of4GEpzHt22q+EZN+TD3Xdc7YTeC4XIf2zxSTSFkDXrgvLXwgA1Dg7XJaNhc
sfpIL3TgGRf5R0kYIeDN2mB5KWY9ubEHyfxrnL4yMjVjH9eVEWstXve2qE1cjuTXa3JCiD/AgLKP
6fW2VJEhlg1THgbTVuuM7+HgbF7uW/QEbL2wK7xq2rKigBmTtyhYmrbBoApLfhWvR+rwF6siLtSt
Of/HkG4Y32iwkah4W2lw+IIbw5NG+zs6TCvYSqzPuVeCUQRrE+FEByyzNDJCdASNvJSah90PxGwq
D8xxhf4EYrB1kIBbuiC/PTGg7WixVqzzFM2FrCchEmpdxVRKnUJlHQqQ8ZNv+UW3P2S2yUjstixN
1T41BQ/fqC6QBOD+4XSR8DkbokMF6QVWNtA1JJrdh33+yGJqrm6fqG3QFMDQLp0wzxgtt7gGNtas
PD8ZZdcC/8MrSquiOInjQFT7MOW6y8ZVXy11pAp31nPWbhTPmp2Al9nZwbfyElif5r6RwZeIQM/g
pK+0KMjYjhnsV7xDR4WylwViAJqZ5yp63IJ8ldN5T5EN+UE3DMy6SvUj3Dzrs6VOAOXAaCT509SK
aiTeyRF+UO7fIK4ZlyWIuT0bbdEgikT9glOdn8Eeh8+f9X/3KYohgqIgEztgKus3qzM6YBU3awnH
WJIDNeETWxo/uI4H5vcIumFiL8zik/VPTWYxEnw4IaxBRZNpRbXd5dcIiYjhvCf0nq9SLRbCndlp
UEc5bFJzd6c4nSZx0Qu9aTp4KxjqX75fWpjgP2/nxV2mBgIJ10FMaNk2E8s73N9+AqJ00CivjeEi
Dds04QNFrSG5gfBHzUsSULzE2U/hQV5ewoG67GMv0C5d6ZVe8dOLre4R73lD/W5N9tggMjXsycvZ
j0+lB+kLR6uJQ5/LZs0Pq9olFuB/EeJsSWsoGZkmrffDKyNYYWKlwHbwgjtjSBQc+Kkjh0/DOkd4
5VJYQjMkef3fHbKf/krV+Of2fIWez109f/lm6uEcFFC4uzu6/wc/L5ELoXn5LkVbbhwkVOZxvcfj
Sopfq7lGvlzsf6tt/642GkcCf+J0+Nl7vqJrs077WFee83EEnn66/SLLqTDyDAaE5IwZ9K4xydz6
B6uAmQ9+3BZdKzZiObjz0s5A3Yz3ImHVwy2Htg5aJtgA52/PYSo+s0Q21Zvdnk7bX5/2C/fXcIV4
J9iCdy0oPZkzoSFh3l9dCsrAPc6wXQB9oOoQ3k2mfXKsH8JGSJSJANukxUjwOLsEWH88Z8ZGKHR3
6ES2zmcjpYp5nWHvcJhrtPM94nmWFpmPQmzRjxpfCtqXWxiyYgoI/PFdTSoKvFZox1ReoX5zisMF
6Tpi1Rm8/ZglZBiBgNg9/3xZquix1Z9rqJ0bbWqWfXY03w+W2Et85tQznOUNs6iuROMHQaf65a62
tkJZvaL8doh1b0D8Q9ty6PI4QM7BScKqxfC94PESWFT11BJ8irSxQ5VqMKEIbt93L4IoTtDeoIzm
38EYFhskjOXqmuqgIFSOnqkHLXru+HT5Vkg4C4M0/ONAWqBhpn8z9IiTGgM/dKWq6DFGGo0EnYz5
GvrLC+GGYjVWLzwni407fB3wO8GGJlU/ZDpWwjTc+0NMz24daU6wi8Zdqp5Bor3YkZjn6OUtSt71
JI6FX49XG/DeGTqYasrdPm3pTAHNj/PIUgXPayoZfwV1awta1clHHkQGBzLdL4S9G5P1AspnxiLH
MYl1RRIxoVr+w9cFZiNEQiF/VS+uX1f3UAhBbQssSxXKY6/5yLBnCkqXI66DzvULCIDsjHd5kAM0
yWAO3UN1IjQgzrq8ev/eufxr/NInFfLzNFTec+a2veNXRtLFLIBNcrKFSUnmmM19TlyJs6YUf2Le
xez6zRIb7hBKLyVCnIsMGtonCXzt+h66NW0I01SAz6l/1/GIQXxyCqZWcIGo0jbobjbtrPMT2dxS
yKY2v1GK6StpTt2yS9ty93sSmQlD+8qACIPl0QrrYQKiA5kFsVdrlCy6I92qp8pWL8gnYjUaZDSM
kbYqmWGzUZr+JnYai6dSpJ4MVI3eRFaxTB7xicjXPKfdtahGl2bc16txTVZC1uiU4RWIXUEmhW1J
Xi2qQJwwIo+1RMTXwXCVfO/Dqespmjg+hPbYS96GoMfJ30QVDai4V/Z1ulwKLwvTKtaO+2rNPENV
zGSrb6K1KwxVgdSmM2/mAmGQqDJUdKVIELBxHLoVK/EwnqpypkYtpo5tkr5GEOEzha4I0HBrVLTM
lmMYFOeJq0lUK1gbc4Ztnsx6ysEONVPBGb7aoIE4r6caVeoqDyvtV9eKEXy7geihLzx/9YpaB1IY
nc5dFW5kqsFhB22JPwC/fCNTiYoHHJbP9rf38pzezAslFiM1yqO0R5jT1x2gFagXlIzHUwQSmpUv
I54GOIpLcFYlxTPwY+JN5bh6+ZxfrTNBhWd76GMnqbFQlOI06Vdu/C3cvlvDZgDgc3PhVEXYn6OG
KX8eLdo5RWlBSgkacsbPjy6gw49VohatYKl7K+3hxsehqzyczo6klajFQhn4igDsM3UNsCgFeo0s
o2MCvSgYLggkZbIPCV32fMHeHzxhVcrnTwopOahXV3mAS//Kozarszjs78Dcq2bjI2WZb3J/5YOY
xjwUqoFe0FCo6LRRUquzoOqBsIytjhdSijl9LLpxO7CJgdtEP13TmBQtTZMcsBzD4CEBySOfGw1f
ZmuF4sBuQMqTQvRyTahPYrcGAfQQr/qpPRXfEUwvOWgbzZOffUyvnVHkmmBmc603J4jWrT85nPpm
Vgr5I4lEmYHGG3AjZJM+SNfPokzlSwDgWHxndTF8DhJchKz98eIT85Q0TdIwVDqcrQVr8YiGjYcw
NIlruX7iKXLAOkA/+93z857Jy06pMvU0FNFvdCNdoYYhdbf6v+rLpUzpK+ZHqwBCVkPYKvYwm62T
UNSANvfZUIpAjSXP26cRaEtxhEMtxAlkF9yRO3NtWzts/zUDTmp2zULlNlywBotERYcdn/HMBC88
1DUmUr0BdrjAucZeVHpT4CC5nuWBKXWSHvUYuTzf5j0xO4E3YX3JuC4npscDJNp8R0LZtjD73+qj
CqdvrhwKO2xgVpkmoKALB0j/8YMZiH+ehVpxvNebF0Actq2uP6WCKpXyLCHhhwcIaxGdZi94ngXu
LfukEHaZCanqDLHMiROZvQ4cMkMG3ZdLU3sh2Q/JHdP7Gl+Tbos/ArsEDQTbadd73+ZLYVtbTxiO
PNuGGYIJyFuzH66nQqkhQpQst6SLAKAQ/oBFri8+cd7x1d/7huy843nFmL+lsxcQA6RHgKMyvDV8
yKRHZKYqHkD2s6SE6OVYwe/5JHaMxDOdhHCNvIVDLpzl0hIY5c67MQmJqEj15sV0JaHfYdv8OV7J
O7VNqUJc/ts1Rx7P+RDFHGvwhuAC6FzPCxxIdVKuW4HnzFNsy6Un0lD/JrwYKJ+MxsoHDwiyxHb+
dl9I2R/8ynVz8TQEeDKX8r4amE9KUwlH66AtOEJh/Bh7ItrYOM2j9gBhrxFaws9YUpOaWWatNgTf
l8wn32f3Wi/sj7mPspWAWb5GxDaTm6WqSoBsuun9pzGe8vfwlWUhU3EmyALBGqFWW+jmOc/liOln
1p/vtiVZh+wOCILV1xJh3YNDXkEfIoutesiiaEptpjPb6D6pN2aKh3QE0xSQmhx+tUN0HIut3eos
nEiH7c+X6jA8q1TLrFqcAfE1kWDtlCZK6anxipN3Dfc2btYvWYCs1p0iJfh2XdrqapUnz+oN6/OD
JjgVd7VUEmXOKMROZvaArS+pCSK8zmJRSmpEWp5sOYXZEC4vs5Lr0tJD0wI0CvNIqVr/tK43roo1
G3URW8paL0Z7BQ+3zzb7OomOgO0w3+0nWuZ9ghPuQdYFx8/eXCdHL2yL19PtnRSaI8L6bG8rSHPS
+oRPvVwhdsfQ02eRSpwYhFLRLV5jPJDYlJO8izsPNR5eWSZBKQ3Ve7jZztBTmRBHj6I+bdquXfLa
h6y2muilCKm38NPnHgu/VZ3QMECadsg2mIuyTmNAAVfncT1KsUpCO7KATCsGZlamUBOeRlG3A4OQ
mnq3fWJUEGAzm1lXoUYwG3Subn3h2bH+YaN0magudpNvslWz9E/kpjnJcNCTlUfki7ky75gV8bl9
MhBSqgKxi8nIlh8fi6MgzD+llX2AoP3DI8q3RFvXWcr96MfLgfspuc9K85SrkiOUpByFJptuhOPw
cexvNVQgTZhtplKQnVO8G0ZxRyjWrEzPLKR0Uc1id7W5l6o+dV9C3d4DZkoWEpPoyp0dbaPMRoq3
JYYImwa4MNepQ296PdRwrX197T4TPrWsr7rAoNeKIk42y/nKPhxE3u51k69G1umDC0NnsDyXAUsh
LJqm0KHRSv8v2UhpCd9+D7SngM7gJSh+W1of5U2blQfDnTSKDT0jcm0JJ93F/CSEJkE6U3B3S+hF
SF2l4o+WsijrQ3GbWAgFLMy2EyHn6DDv5gAjj4nzVuqI/iaF2OCqMSnOzpgDvoX4Ure/mrkAbvGS
GPye7Bt5mw+SpQnaGIpob8/3wdoks4Hoi3nFZuvkxBUwpJ6erYfA7KZmC5IrLx0DbuEEnK66Hpkr
sn+tWszXmkCMX8y40ANIehmYdTUFTI/4zOc+YhidLWnBd2zzjJoRM8sXcJw6zRGFzX9XNTi5rdQ8
hyUFtb/AAdkNZlgf5K+FBZwD1bvbwmfiY5o/uDfLRDhuwHpCwwYSBeNGSnYkLssW7csuhGRuZ0ii
4Mdg+WLTFo4kjbn5p4a8byNYX8AYGyhk/r10XVyOISjuPyTHEit3PE7ENDwZwdEK/K9xlAd1kW5d
asbhNCzp6mqsxwGh3fHDX4YMKcsL9XwYYRswwQ0r3ESStwCrKDmQP6RRimMLMmvHt1lnucqQyAxV
ZuZbm0C7eI335+t4VoVlWe3b1xPtRwZQ4Q6quRDh9ndkpKqWHg+hBhZ/Jo5btEMu4kippBzdjLdc
4IAk/gtEnuvTxu00Dr/JWHGw1YWWHv2TlQ2eiYHS6EmFDX/Sojx/GOtDML8rjHGZzR4mzWS+Omcj
oMH1yyRweU4Gt7b5Ep/CP0gvvkM0QkcwCdPmMcalhvUsGeM2k46aOoQj0RSRyqJaj83xaIsIQ8tS
8JGzPvDH6DOcP6IvgDGB3dBPo1m/Gnvr+3k84AyuevZVwc659OCuuflu0tTSLryvSvNoPdLv6UE/
j69VeQZWUa6na9CFYn74M1fsmS8zXCUZj/BVIridr8L/Dk0y6jWEYWJDrHUsJrzywXu6JyxUHdVe
AbPez7zdGDOueClJ/15Ih/wQoimAyd2UUpGUm2+4ANHuZocKnPsISq+gyQXL0YgKztrldoeTF56f
bXhCoX2gKwqFqHRwpDnsVrpcnCaOsz0vZEWaNWSD75NxyJDKBvXDNq7vaLtsU9I4Dy8ESceJZGbr
qgjMiqL0iYulgTAMkrD5EPioQKgWU58u/3bOCJLt0VNpL2QdTIia26x9kBhYzDMvh/lLFfngPESY
YOFeTWFYz71VminQRJVX1iZE5fON9uSX+KMfQ5z8dmju3gNwHNR4YmY5/dqf//bqjPMhdnaJ2srz
UlYyscm8MyvPzrIwdNPcZnafQ5WxGl4EhvKCCDa+Q9Y9svuNHat4w4h5dYq+AcEG5u7m08BajD+e
/EAb0htFia9WM0IgT75utpzWwGl+c2GOlFzMhxs+zerB4amsFNZsIqKHilR+xz/7kVXsccEFFzgb
OxdCCvEQEd5mzFci+C2bJJLiqSPdRwo/83OCcJj8rsxshmrZxVWzmayw3IO1QtpjJKh8R9ZPO34q
l6WRTWT86/zOPsu/PF1mmC1GxGeI7zTTe9n+URtDi/6fjlOXz6Q/0cw5Nosj2Iuz7FZGiYzx74HN
Bp6mmqXQyCBnq1bvtKnDA1NEdi2gVwpPMdASEfrZY/wgsPC6IJkR4BW4+Ju5Vk4JAmXGIdvKtUe7
54h3ilh3OtZPEBqolhJNdvb5J4NX1ynAdf3DWyyaBtDcZbVrOAV33eGnpisdUol5Z9ctIh//A7uD
5QXE6awAmkQQQjvJF+rvfdOZ+7ea37N1ymxItND0k6QaPv5HKYoW+RsPfXdVdVPq723XuGC2mE+9
bRM9aSFw+LSm+xTbcFl3Bm2LWVvLTax2XFjNxpjKOVJPAwOgzTEjqaa3OAniYlDtPGjr3lx9xWA8
AWyj+f8y2jSY5PE5m5DI2Wf7WZ67RKNVfqHqS8+wBEYh554TKQVx9E0pxPgitDytG5/e+2dt3q+T
wVGpKX9v96eHmA98C0Dtyx4XQrXcQv+yLFQ91EjDjakMlharLSVgtR77a8S79zvBTDzbnxpZpew7
nXRgkfKT0FBobZGqlP+Ie2Ydr3RBZk3QJvBJUQ++Q2VArtrwH7X3xvhvzOMJoN1nRSlhbiJSCb2H
DgaNfeeQmCyQGIuGWyTLNXJfjL89z+Ze+XvlTD8/vjykaw6TYEsMIcUPLE4vhKueP9Pj1Qo5Nm3+
HQB+/w1fQIUAKT5RDP9aq9I4rtJDMSv2XV3qpexjHBLRZR+hP8/51UL8oqYzrTCODnfSE24pvaKd
+Rpwo36sT+vrTX/qtPIsAtjWUZTTiZpoxZlVMkkdTFC93wZOZTgxu09UPaKfQF4Q5wq3bzHElfx9
+Z+XxzQUuK36tH7QpTrGQCZut4PcHispzrjsaqCfODOCgR1YdCEGvJPnBtgOBD5EZB0XiU2yCMo4
oMLPP78Yh82PiGmXFai3A4YtKOPR51I2uDhT1mk7/V1VjycjTs2tYPkMIlDJTbXwjZ9DOEMLry23
wlKEVzXJ39LAUjTPShtgtJxEUEwHMk8ULFwjeIi/9sNRgcnTrFXJaifJww5D4Zn12nsdG8LaIbLI
WQF5AGXgz//p20E4ejPOK42/rWh/FE8QQvdQRnhiZwz4SNvnh3VWV8WryPMK+6wM6vkDVXLkWSzv
JOR8YQ+5HA4ZbIJ8Ag1hJxRD9ThdpIS7hf32Ute/wUv0U4TVzZhDtGZBnWRdhXr3COJ741tm3weK
8RK7NVLYtHpvd/RePNDT4N2po+G6wGQ3mCSo/wKayUlEtw8T5iZ5DLvVMbU1RMbZ0WiPCPio0LpK
AkaqMIHaqixp2SyCjE+DsYFLDbRpAGxsi0r8eOhr7FggorMLiv+E/1Q/0yLsQwscUjCimDlIoem8
G1zQjmovY4ASeNmbh39dkGrSuulypOMPbVDuBf3RsasFitus0abyBcdQIomdHM8bmqA0hkUI3mI5
wwXLYblCWzUP7AdPVw8wMq8AfgD+U4eG4ZGJoRllHbToVFQU53EkJEARF+KeUT15D4CZg/+iVO+j
t3W7Tr+GFQPvPL7I4uvTCFoKou4eJUsQb+How10U2e2wjzsGDcLfMYFz9L84HFE8wqNWoUBgMHU+
UlsFolMg3nsttCOJtXITzVZlF6yQLAteHuE6b+knmwcffnNOwjz9jovPm3TUH3KqepjpHf5flNdb
8FHQObtjlbQHuiNS4M2EHzkPSqbpbt+RgBxCyT9PuwxXJnxALh/Po98CjPFMf0aNpyI94x4qcYUK
ptjVDtuQheWF/Hw2I1BTyMLHO/FrXtmDXJq1ypzJIXYDqyxdNJA6AGdGRp/+mAPpk9I1RYISbVgh
whmj9gMVXzoOBbi0S9s20VR76uOAZWThzEMQYG8p7GEozdBa29nYd3I9++oDcRUJ/MruP6qrY0xj
7jDO57uOdUVG57iXqzqPXJDMVl39AtPTGlSLpsQ4DGDLJ3THlHsErfzc+OY7T8Sc3bqhn8ERRk72
AL94mVT+C8FSc8uIw4VGE5ALJqB6yoSeaG1VeDY9mQ8zGi9Y3wGthB2IYkEK12jYZGunoDuMeZAW
DkOjlvkzwrFdipcr5J2CeIY7IoWjswv1JhGMY7PLT2XR4CFl9icZHartcGc40P0p0OtCE0nxxvnL
p8sgrFrHzQ0AuO9smLv1K96HvCPVASMH1GyWAHBa84LY+T0k/y80AHuxgfvhPmdSh1awGIV7z738
ukdoVG4Q7sx2JcM6PIwuD/pO79Sf/GPzeESZrjMJ+E0xQSzX3Jqxl+oGm2TqmgMBmaqip61+cV9O
VTiLfGlqHDwBQGqa0ukBkicOBB+EjNbV+wmajpf2qNxvknSS+Oxo6jJ57rJovDKey1sVVvTU7/cN
11pHOw3tkfdJ6tJ+DVujNS2PB34cOuutV25d7e9iDfJIA3gSHajChmjNaED4JuJecv8I4ubGHGL4
81BzGTCbcutN/QPgQ0bzxhg2x7X+cfnW6Knh/laiHpmyb8S+tB2RrcTU9Dex42HxYi4RABep2JM3
2V/WERYlwa6HUMcpbE09hQoH4Rk4YAa7uBLfbLacWU+ojUAG8ckGCtVBRMecPlDSzXQ3nMOoh1kO
+QOcsI9fXyWkL/GuGNxh0dLPL9w2zxG/tfjbW7jL4bprZevvKxncQp2BMsutjb/F/uGx9UNrBjnD
KxAvq9soRgFggYlfci+UQSD7+lezDOvcM3epNO/0fNtTAX3/eXYcNK5ff4q4TPA43HI6Sz6hPsf4
7PHO/mooy7jb0NspEzjrgm6Dqz7WK9ukd3RheP9d0nGy5Lu1SlgTtUU40MP/lpf9rcLwQAbLt4RA
aGNNOzmPoQBdq8zr420o6YFCxTQLlRRkb1MjCK2XmVw7ZEfRpIp/t06tdZnqsKJeVZlxATRGXhmS
KXukcG5ZmpxxH1An+YJcIy60lsB2mktPDOUzeJI/fB21GjkFFShVOuACuwaDrDmB/caKiEbHNbEM
l8E0+T2g/Za2SVC5o9QOmFnol+V9+P2r7zq6KG+BgQaokgt7wc/wdGF1BizfBMy3jJYGuBibqVt9
1Be4Q/MAYnK39JieGLwLZiIZogn9GmTT1deh5pinTS7xCQfCINLWrPWxmu7u8Wm43EY16HzikZ85
DH01eMap3dEPbzGmB+2LUNRxYN8zsSK3e7AkBpdN0BGaqr20heBQ8xAinrB1JhDLf3zlm+NkKF9U
GD1kiSURx5zitchGVlsGYRcJCNiQGJ6j8KsHw+ioFwlRK5nKY9eVDQIhuzhRlt5TrDsFibthWjfP
4wFmtCiLQbsWCgz/orP5x//5mJsl/p+WDlRs5UDZyg1rCSxJEjwR8PBFbj/WMuRZQxc4IE0v8Jgg
GwFDTZ00ZJvV6jrOJnR8LDUr5YxFAkXSndWMbHj/JTFsj6DQRihMPNTSmbGGexatTJDVdyvidXpO
YqPvmTeXwRWAeUqo7jTxm9zxIE9q9ReBWzZ6DCbDjv/UPXG3sOW3LXITC8bJsRjidgCM6Yqkj8po
EH2cViTaw2zgtOKKoqhMNH+D7h9RxzTDJD3Qb40u88VeaBgAQ/pFMRS+Si6X+QsZNeBxuJ6+UQmZ
EM/YysdpEn4VCeuJ/hD9iH4RVZzXn9pivuYHz2eviswNGsBBYaW9q1AVM7LbaOORV+xbyPcqyH7s
fXvN/fpu54Q5JgAiyRuLRKa5USr+ISqRZaHf+8UudsUArbPl2V0C9+j9ia4te4zPfW6nQlaueoPq
XPb8EjgjN1kPXZjWlXcTRjzQghVHFeYedpfRpsEV5MR6VcjjIbmXt4E7tVmGILQ9DxiNmAJSd1/X
ROKGAELH61w/7QwbTC7QAGTOuPifzDUro+CHc6flbIygtek8Fw1D9khC95GliHFNsOnjzlSJhvlB
6+VG7DNMUnlJZ3jGIOfSOQTiRT04Ak21jjnSuaIHhNewz7/VpjTWNPiz5LKjPMUjTLmu9JL8lPXu
mo4+6WovsIWwlSqllXkkW0s0mJgiMd/hbco3U3l3AUdU6Cd2l2FvesODquIXDbT+QZqp32+zHEGv
REurZugrWuL4OIKxT5q5Y0aDYOeoK+XpLo70gGBz8N33TVnd7V8KJac2XkG4hlyBkDhOnLAKszv7
kVruAGYZhXOVslmYY0k8A+HW7fbljBUyXo3ihRTIkxQyV3sCmbSJxY4bRBheIqucytpw/4rxac/p
+YijkBDbFRuNch9LH3sQ/t0THvDeaATr+lfkqkkLXn7pLdXhKL58HqJn6gjs07MpnNocUrjcPXOo
ibhoXLpczjzIbbSiYnQkg0kg0l/09VWQJry2YTTPFBqVfBjxjIdJg5uR9diakVw8bITKzwo5nekV
BJOfXw/jDYx8tdOfYvOTXVhbNuXOQk6NBPGGYkhCJXnElUjSVOEpx9kz7zTKCYlDo/zQe+SATEEb
23VD05sRUVX3VpQILHW+f9m4JOJ7A8sbOzM6ahPaWadn4njyn4Y/OTUZvZASPLVNBSCOKGUk39ES
CIoU8V0K89Rx3g5+mfkG/kqbVRSBCPwgI1Xrr71S75CODSoa1Lse8EkfdJRmkLX02LPV+YMYgN1b
yF/zYrnxoN2XB5FdYs7RSfL8t6gHBdRHEeURnvcTLyBKBeQZ02kHRsu8X7jG0C9c1wo+xo71puAo
7btiuRyjukfySH8d6VKRBGFUF2haXZRPFDQ3UxgvqDXwRSMQ02d2XsYVp10wOv68JUjBbEp3lm3F
mhLvGaakQK2ceMDrUH7wJscKnewoT2VWPPJMxJyqNQHbqD8NUbjJBbR8kT8bvIraH6HVbs2X1pXz
ShvUqe6ZGQZVB5tIqlniloQ8eRQvFDF9q6jSw9kMFlQV8wQWa4nl+pXx9y1EjT20hPg9Ug9IOoCh
mk9PH6HXdfo3Mh9q/83woGFKaw/oMUiD+SQmQ7p5QaIr3SAqFrpZsv3PJXNii6XsuyPaz9gtlpm3
0io6ba8/frbaHG6hQvT8seSZoL0n82PDcbFY4/Y8lcySt7gss/3UqK6yUcWa4kf6uQeG9fMwQt8q
E1BNM8IiDySOvwHkriA9B/eno/Bz0mGN6wi+sQ6uVIhYUl5epKQjTWE+nh1KZPFx989AwfdH9XTF
l9xQ8xd+ZRS1sL+Ku9xMbKIgWJ5U6ET8HCHkm0zoV462rGFBDauRnmgcg7O7fyBqopb4A1kyZ/j2
DCpErK9nyEwfIruklCyYCzFQx4vBrmYUOsAPWSvV4mQyAyl1H3NT1nTW5H06f6yqTKTF/Fzuw+nc
NEpeXxi5xOqE7Dmeo3hleZvT6ooj8Vv+oHWdl9AEJCg2Dj1kOJ6L4Y41nH7NdZCKJaVXYxm9ZhhF
uyBaNHoLongrOJM9iBdSluGr6sTZSjChIPIW1VvxrFoDK4/fsoiMln6wATFmqWyaEZ8nmfTVeTVq
9Nnowy3TPymozt561T1B6bbT8tLOSIXd832XLwOPHRAzbKWJ/DO1BW7qxtfGcHL6mPcIWT2S+zBO
lD6raFhbob4E/LXnT7/Qc1oBKHaqWlgxX+EBiN7WHCPF6Z6QW/TaBwqBlMQ8PbvH5FI68k3+rjIP
vUESSk3wKqI4U64V4e6OF9pDDGd5haTwv3GggG9ARCc/jeaV+cDqrIsMS2Nsme4/gy8HrMmpHWVc
JYVtI9NhPb+tOrLae57WQhgLkfZ87f3FwWMzmE7TnrEqFPynPQS1MjuehuDYL4uC1TBwJ9AvI3aW
1A61+rFIQwfJayiLtOLX1c0WZHzOV5ILsbtj3wu6MfZVcmXOQv1RfdJHQ9cp9BTaXuAzZLv2FjFE
AxhV0EBFUkb4J8i/mQcpDD9okfxtMnguz4ZTWoPFAxIN0rL8caAbrulH5eBAphd1YFPtdA1mjBTF
ucfy127OSDo9MRUJL6M2WxL+7aApeOzGOUeY5t9t6Few1n094gJRDPDPz+M1p0YWYKW5bSy1NLXZ
49PLq05DEEa71dWTvVDnvYlZhm2VTUvHWauO+WUTwAiMy2LdmRlZ8D5ZIrE4hIU3WeVJAn02NSol
hUICk9bcJCtHD9+8P/2e/ZNqdxOaY2OkdymreboARnOekVALUzOhQoCgyZARrAp1a4OnEDxDl6KR
Mlp/BVZV0aVJybVAmuBQErscIllbGjEoV1J+zYxnfkztLEtSxFmE8s3V8/APKiGk8Fm4tXeP4nAU
cMu+/0vyfxXqfrgp2fIIaPiDjyoBCar5cTn4sa5FmF2Vcmpzcj2XZ8NOMzQ7Ve+FuUVg2boG962d
831ARvd7dfZfCPLiHIE13L9DQAVaIr2Qcrl20OwhzLJF5SVBbSVAWmhWkJbb1r7Iajm+NKTx8sNY
UPwgK4jpGkowKRYCiYCUTLbj2PsCzbqOGxDiNWgw7DCKCAPMdKE+4gzlYZsebNGrY23mkFtkqZ19
ZVlrdqu2D3WE6a6vcRCvsgjg+lpHmythA/y0UAQSQY81QT8b75O4XpWTK97x+DY24NGimdvJIQlu
R8Y83kCaeCqe7gR6mUDJUtUfKPZ4aIhM3inEdRkLjURsa2LkbzQDhShAhLI0Pc9PxyzZ4sfanHPn
qccjA1APAAinkVWxGfk8ZNR2JAxYbZMKwRaBNp15V286a9k7Uz+fzXvcm/k7zjNjoyUUY+n8zcnX
UnrWxZR91+ADjboCJ82i2fEgJBZDkHoMZ6R/eC01BlYxcyko2U5uf0xEPLnwK8CRDooi+7C2eKRd
IV4xX2Ni9+wgBbGwUwnYGQ6bcdkYCLENKQeRiEYwPJdJdm2JlQlpHwKY/WvYZ1iVtB1L0fcEuObg
HQPoWolpVEpEZo/7jU6rq1nCERPGBxkenaMzzx8iPCUnmxCuseU863/UTHz1CT1Mvtg2W2aPArZi
1rrMU/uSZrawlnLAAZYiGsm4XSW2sucuNXGGvzPLyKxOPAUsJUDJP+ihcWHHX/EwMqV2youvde3H
iWLDdTxBTL1w0uIYETzJGOi74g4qMMc8nZKjVSGmXO1BmLKX2/Nqm9/VCUYPnQVAf6IJ/B5QWNO8
s2VotrjmuKqTGOSGEL+Sk5Y2DewFSFAltQctA5qeWybzEOKnpX5JKCKeoehh5W/A+92KZU2ytRmm
FlD7lkQK2C1FHPCyB7/WHm1nc1CMY+7ZCiZFU/O01sjLMezUxKjPzDU+jZKmGUdffOPfnx+IUjwz
wMJd3NxCOfhLzCg6/7jNLrNx4+zmHR3YLTlrpitx5911jF+eEEcASo6UbRaFABNCHWwX7EgXtzh8
C8P3N2iLuEcU7kJ2dkfmiCXqMn5EE6hKeI1OOuOam5L1jHH4E/RmTMEBcgSggTKi8VKaq9NACiax
4ei0dCRoZALOiFoTS/Z06JXp2gJDlyEBYVpSFYiDPII8bQPD9l0e95v+tk7hQnAaQJFtJcvYxHhO
9vyHHbDlOeAj3Af+ERNdNSXqICJsCkht0aGMpbJmhYz0aeQFUW/QoBH9M1dasZFoSoCjfl3wo0We
PgvtCxx55Kx+yPfmUmtuOI6+r6XkKeFFq/RqgcqoQNod+JNGUDzDy2d2GYLDAWwd4Fc42LmIo93S
Y+Ob/mOnCPVn/8ucy5EAMtgxdDd3sOez2ytocPaxNUaXdDv53nO6+sPc38aeNWFtdUKT0TvL2No8
t2mfAiabptVncgTY004lt+NKlFzjPgOw95l9qDmsgH4qHNHZwpnhpk0XdOtcj4Mwj+NbC+rP0V2L
m6rRL972fDcuZFChN1+nG1j6RfxO8W0j0k3Gnqcxy4m7P4UnPiApVnF1bDOZmuTS+FXm3Gq7pygr
AV/OC+3maMxCJiWZkIkzrL9AepT+CaCcDCdOKpX7glAsGhFFu+6AlUsNOlYIP+S7Xd7UTcvF1OJv
jtqxNyTLNLBgaON538En5Jl+GHZzJZU0ypptddQbjpKsZ7F+e/FSPJQvoC036eFBxV5/ZrotMVLP
r9NvSQq2VrwB/zVfEUvHo21GJ01iaCAL6HU5MlvnEdWCnBCensFzmoMrK3JR3Z/HSxWnV+6ZiHsC
KlbmhjIICQEXh/vg97RFRPBfR+mIh+n3pptd10rKX+bn5wxWCXS7LeTbKrhqFwIDRcaAkaDuoFDl
m/fpO7TxRKcF9OOUSTz9JWiCxsm7ab0ueyQOhHkbp8KOJKX+oyQIKNfT+bO8XaFu4lcUTSgzfROr
f/jPM85Q/NvRWzQPHuM52yKlQN4u7cZFc1x/1j+o0w7MdhFHZothNSD8rReid/FtF1YgcExUhU9e
6Q2egJ4JIMzteN/XPOQvESkNaPjXRQOTA59LHbOSSNflNZo4HFjPMumkcZ0KKYs5IQkOzeqd9Lep
oUqcHs8h5AqAbjq41+UwcxzBQ88wt4yhrUi4jfas4Kvq7ZdIFzD2A0e9Z/gvIJDxmpQwbUzszNgp
43rwvDmRG28Tz+17FXmj+XH3Gz7G2x8CgtsRVhd22rENkYvXHnhJKJZ0rspMolNu9sW/22EoGpIc
EaYwwZW8xRs2a/XNhkz7XyrZa9LEyY8i7qehBh2dGr1WJCmcntzgtwFvMQjx+idCKE/UtJMBbXMA
eB404HCkDjr1kGHvileeFUkSwf1LfFKZw5HTtKYEXKXo/ELaA79WAr7GlsGXjTv+kmZRhp7s19j4
6f+jgrSP79g4TYtZZohD/IHmAVFGZxNrs07J8cM29RtcridK5xk16w+lap3Zq9NKnKMo3NEipgMB
FEgwLEz00H2sIxzJBQWpWviSfDBA2lgJ/CMXWeFGnmJAzwsM4nEEWpu8cD19SzF0UIegg/U68CUq
9KTNQSzPj0RvFDliLCYy0PJ/wVPc7ga73OYEwn/5wb8OfI2U3K5WCPxQiRwnlCwRVtajrriwgX2Z
3SNg2LyDVKNc2qgH6/RUaWFmqtyCwByrKxP2FTtp9YBR6EpQFucw1HYv6WMM6AdgdQUk/Fvq9c7b
Q4509cQSv2AL5LypnYGfCAmTaReCdOqAm/OHOLJ7MF91b5wE/ggiDX3RvSrt+sRjKFBf7UP1T59I
SY3vFzQkyAJzcHNe/mo+qCo6yZJJ6MZnVBJh5f+XPQ0BTnpz/VoMAm/VTMXjsCgwb9yunjXnPWUP
tUSbPvv2Lq6QrYnaXl+QoCB/eUT2I/1Ku4BnWSSW86J9sfKhDnCQvyXI6DK0/5V2nd7mXZHeCeHj
yQKOhd2KI6c/Fr7Ob46ZJvsqBm9cTeOqyB8h5JV7FmONNsoVtk6jizcCqTtpBiDk4Svyz2F34/lQ
aprNLUvQ4exgWlhzcAho4oIpHiGMJGECOz2BlhsET+M1ABFS4hb9bURDQb0vxi8yiXZgwqDTSX3F
L37n+qt5/BHibKT48FB5VdcAc8QI/K6NkzBGC0lmFatczmLoKraLAWQjlmT9ZYS8P/ZRGu0ZGhpe
yp1PyQ4i5Bd5XS/5/G3GsXCssv2AcsxZ2k3ckF6CkvhQhNabo3OKMMycj+VJOE//M97+uxKaZ6UO
uOvjVTsYAwI+HRAgbaEsrhb1z9LNAhNmvxVFMP1ST8j/TTzF0dJ9yrndM1TgkfYKsKNkaT0DFlz6
Tqw/hLyK9h5ZZ+0u9DrTXww4ogYOQrrZag9EGkYf4D52iWUbIp9YK8ViTy9azuMQ/goQwhfihq/l
+gGxVpZAAnrQWq3+JpBNTN3LskKVvsf5g9vMmgbFcTUdk4oZm3tkZK1M+qLqlqppHqvzA7jK4jcR
LL4jwBW9L+lKa9utXSr8THMc3ryPasa0P21yo3eb3qD0uIQIwA1o39IlHUxge7SCua5CQryE52yi
01ON4yj3QGz54VidaXwpa5Tf+1VSJHGdJwqFEgHD7TUjL7Oog/bLAdHYi2ee9r2WiMPs0RWfhlww
iR7OkFHgsf+rrtKBlkltCT6vFGInUZJcMs3Y1hL4JqrpYbUHscKky4GsGewEZ/AOmKDiHuvAh1Yz
dCtZ0w+2D8E8tG+o21NvQxxl1qONBZXcqFDupJHDucBGOt1/VbfQ9JQaqlCBdIz4UsDb/Yv6ukRz
hJMInij+669UKhGJHUvIxnw9jtWhj/eYUOQh37ALQ9MNujidbYPKCxpj4qc641jwYr45mdUMZBWq
t8vUboe9k2eYo4PZ0AlkJJuH+0jSLHqm43EkqjsPxPhNOFnwcoY5n/MEQjOTENcWDbwxMG2uOCD7
rjFl2HYbkbbYjT+jYziKwysWpfiCREFL9hjooXRxouvGDROCBjuC2jwW53aarTJi35WZHSiLLj0b
1wD+iuu8KxOkbBCjJDo5G+Fsg9ui+1LjhdAKaBI9YUy88x6yf6dfqjmjQyVT5OoH0dAaCzcFkFEr
mx8CDGtpNR9i0d9qE4wq9lIypWlnlXR2Mx6BK2KTZVaq+qmX69G9isfHZmldPVeYy876iF8GzdN5
QxmGHmGFkY5gxRikLbpAKWAcjSUzcXdeJelpFZiXUjXg9Kj/swMdBtcD7VuThPo2K+ecTroSeN0b
6ntEbHbG3/AWOY0K1JIkNCXI3KGgmAzCZtYNKcGNJbu49m1Sdca0hd6/T7RcZ4bQSxmIOxghTvbC
hseFN8Kc4W7Gc0F+L5RaA4DwVaMt7nRqVWWSP8TZURzjDO3OJ1usHElhRfN+zYLOsxrNTVTvGMsm
u20Rb7PWaHiWJrqR1NHcXIFe2ffo5C/rDVEcAFTGXvr35tU6rbZcghSR4ezq38P2jB/RzunvRGIb
7sVsar80A1jZ3xiluOLntGQrcPSsFLGJuNjpr8nGysUjeehxJqR5dPawouV062uMZ1ELZK5TCMDj
blAzO7njPniyVHcxNYnlBK3pKGe51auz5VXAPjinT8nmeaXoLCPjdnMpIrUCw42AobH4cgUF4Aag
MpkB8g844XlNrn20Ex3Nw6RspxJH2vtZ7508jrlq7DeW3hj3WaX2iXSWzWhv1bd0RTAdXblH3iIr
ypL0FGpga63gBkLL3rSypZwiv097VRUc7cprNnwfd3H2KwSsaU7kO+4ggZYkzZJqYgUr7kuJuTYi
+Y7A1aDxgd9wkGop3FNe+L06T3etanBSddmJNCH7xk7vaOflT+Ep0VYMDsfL6v9+dy+nf6qcw09b
GBpo7d/pf4IPTxRWRCQ0kACiJDkGhXsBwCoQ0mkVPUnBsqgVuLMBTuNFPmMPdbimh1DfK+NVGSG3
uDt5nGa1azNxp1foqakSqG+PUA1Djoc2p7IhDfPc4SsT6lFMnz5DLQAjt8/rIkmyy48d7+ptcNCs
cdO+zMQqssjN5V0vzm0FuEY3IRjsJV55+387QQZegDYawz2nFlDQUAyzf94CE8EO9e6yNr+B7iir
AzjmVEb01L73yeMr40yTLeISVAuayiB1MGSOyfiUcu0gphylcF5rQ2P20oY20NGQ3qaFAYyWaL9O
ncnN1xDMSIKkHlmHXmiX25Q/LWFAzrouqviwEmzP/hgj4fiD/eoDHVt7NHWo4IZ1cO06frrtXLAl
iv/OD7AKCvPS4Q3PV71wwQ3fpypAroe5KAhaV+yUcCZ9N0lpxZs8Vgeu9GYBiPQIe/g1ou/QJlmi
UmP8LhHd3N74Gv4ahAwIsCDq4pytu5ElHRUzgIY/NAD6Y+ZcCXRfcFrM6oNtsIFOJrzBAI63zPEX
aUDLDE/Pa67KrvQ1lX60sTn0ccw/zpn7eHOl1X1z5aHndtp1pGN/eKxrNKDmUjDsUD9+qBF/u6ap
9Fg1NudDyOp0LO2112pKdwccIOQobsdxr14FWf9xWu+e+jaPYWBtLRl8isYQ5l4YOAGJtRU3lipf
dftBgIiVj31w0CXH/BdW3CZrLGxkRsNl1jkAGTTD1naCxwS3++Tx6kyrImdEiBZDg/0NYmA0oIja
fqA5YhTkXhtmtP66Zi8vxuwXNPFmB+KiV+1b0iKWhiTzDKtUYVDhbJUI9gwcx+W2ER3w3aVvDDnG
GQfwwxniusNDOcONbby2DFgCv/7ywoyH0TqfuQMZ+F5HLfV9XhKy4r3z2SbsocF7sQE0NKwpixbX
Mu8HzQAO/NZKYtT/wIG3gD7M/RHtYzR5/3/LCVsCM0cQwJ0RnoHvKIHMK947X6GYKQdj9R40Lt+F
XNjeoXA48rfQwsz4643O5kG5+5QosKS0bwxzuYVogGhVM/xq7yaWZWrpQ02ABijXuEf+v4RaT5R3
QohiugDMsH7MKApOnMn8bB7XTtTVyAmChcBD1tAQkIRG6B2TQyrq7KGEhWtEI6iKLXkqG3RwzcTh
JJJ++7WLPbBbCSSkmJ8B52zYlByIGk7PvvkV+HXEAmzburYsyPyaUGa2Ho+wj675oasfWLWtEPo+
MrHQkUlfhjmhP16EhKUBVYZM1ntrzOzYb9pvuSHLQ2m0zUG1eOwo8J1N/fIrLJ+DcyaUoBEc1hwg
x536y76HY5so9FR0iIChj3QBoe/pLaD9NUCxeop9kI9jhIwvmBiE7oD3fKRI/wbdR9zCM0Od4lSv
5H9hupxzwlQd+DVugbf6EkyxwuIAiGHYUdofc6nc0LZj0pVxxZYmjwMxlv9j7gDdTn6cr4I6jUzB
7cCOM4zq1URbd2DgC2DZ+jk9xPN4E7G32YablcvYmn3Yt3Tp9oVhF1WAp5wx+EfOBgXwph5gL/Yw
cvsnP2V/HQB/pnNTqlgyxFwTMS5AI07eAkR1jDnCBYXnMaCbLPnPoxQu95w/XJ5ORO4WHB19caWd
oGHHja2SV1MUhEVVhgUnBhLNz7RVFBOrQWua6CwblJW/YgKGRFZs2tfKcF3nWUVHCRODKSuyDKYX
7kV9OI0/sOqxveSHyeciRij++OajqpNPvRJDTxdJhG9Dc6Z3R4UiOe/RJdgdUV9D6/9J2CasJfxU
W1f73Yv3Vvphrv0oRmDAewFuAijsWJnB//6HnPVYzICq6dtghOa39iV4iCsGD7rOYszu7g+QPA2x
aGeT2kEtRtuSVXGnNQH4OL/AetI9n1CsKP4PEhEi0xMfBI5cSEn9ouaCh/sWumJly14QNC9TJ2vJ
Re5oCx3wQtnnRPyvYkhCQggE1OaWMw+D+b/PFaS7ePbM/UAogeORLUQ2a0zkUg3SAxmoeTltfEsV
etLNWvBZBXQn7Ut3GyUvqPWDclIX616RZ5hTWYnGx78FlqI7c3Ldsx/FMF8jZol7HwszHvMNeJWg
Bge2dpGuIzFKne6Q+ULuohAh+IWM01Mx2keCQx1t33f3zq5b7Ylo/MV1s/AUJa06ZFYcMDic047p
OYOjwhYB8RMaJV/fDIPSSsje5Yg/2ehHlJjjS48XVgbQirvmRHzo1ei8v5IY2ZylkpF3Q/dkNiw9
43k2Odf2GA9E5JJN3WikrgCQpf6fEGC2j05Fod0ZDQ1UwEWddYm8WyS+yN6H35KANA+WLA/O5Kpe
5H1/O9LSVM1oN7OAKZIsfGNHEVv7Vz4/XLeCySWVDOQ8rclbHIF13RYzdKwCvgxUzcYNIIbQSxux
zAW7ZEhtj1J7FAKdpr2Glv/4mtxUmT1YxXgxRFfBtVnQX88Xg0+FDgOW36iFFEQs/b6McFvfF1X/
kNuCCaBLmbQ9hN7oViroTg+s9M/iXw0t7cYMthhJJVkHmod5S34/MmvOUmOU03ggAQPSpnNhyyOL
IOp1oowChuSmcoTbM6NF4RYfxpbJFvOSkqXgoV3ZNk6LgJdyZbS4WcTs7NOb13mrhsTkj2FofY/F
9uVtcPHRyAnp7fYnaIlIUwxDIuhfS9O7YGtHEYC6kYvfMEnfR8s8Iap1bJjpg8jbehrBK0fElvNT
LtHnbawyDWKX1rWc8jo+sA0/DiBgrBH2kIadpjx4WlWz6sT5UoklAoS2CO4LeMn/r/z1rGcUmujL
EZEPr4syJY8et8GDo/FmwSw1qc4w8+ocIaD7rYhpnzoQjl9WHtci6BJey48GKMJvmxezWyKeR84a
7VU8SE4DXBL21cbgs4oWcuR3gICeB0CXhVhfXVaZqRNRx7EQjhTZepyXubQxb6ZgaJuZ4yqCMt/p
/7008YGrSh77UVCXY2OX30KofisPoekXhJH/zM8EVkRqFzZtmPIqLVqs+P1TzdWU32MWzSkGKQwB
5EhVnx3VY6hzQ43dGgd2QM8u540rZq1qTO4/+cwMGLiJQAlRgdPkFpvcL347q8kNtGFbjOOydIf0
mYmn6d07gLp22lga15HjKCMTozj/rcnLY4iLSnfka0GEZDBwBdwjMiHu856ojmCKaSK6OeO6u8fE
hntGEz6ozy1c0b7y5sNMxpUVAiQsN4YHIB3aFAd4A4RCV+NRmDYxw7R0435kJuMoVsJxqZS1dBF6
m3aYMCELI66bbauDbEwPM6IbQ2Q2XM/YIvyLHnsPD7PCwHxfCOyXgGeJKDAud3wit9Zkr47ibl7o
LnW6GDK2/kxuz+YnGGGvoXgw1FAva6fqpiK+37KdX9o8VjXqjVfGkap0AGT6C9MPiiwCdnB0kz8z
PGIXMAkyJEHPbD71r8H16ZEgmIlCV/sb4s86Z39frdY6l+fdqefNSr9jJr4c7+SI4BdptxaMlZOS
uyJdp5KmLoiLg2gzvu/vhCEjH/xwtKljOeD6VS+dbNwzfz2LbqJlBctVr8k6Nf/NaxIk0oyehi/U
whMh6OKAPSMOMqjHV2ZJyhs5C6Sc+We2yVtVWgwmR/JvB8gMh8r46CF/yUu3mSQ5Rlbm2QFMb33o
ocfhD8MlXBOyUgYFQPJRll6n36vn6kK2s2Rsx0emPZM4wNpjS4stk/xgIF0ywOWOuVIOi1hWR60P
UfGt9uEhmgh6oSrMnv++Y4jX84MEYDiKHw2q1pxiVA0RmZb5wiblJao+YJpIiT56janK4GR9A/mn
llC/2TTzEpNHyXFUDza1KWDKfs56u9JrP5ZS2OTcaJGfKyxn2FCtqjjJ+HqSic2xOz3utrcmCPFK
AZAlgULzIpbzLsLQU14HNixzQq3C0EDCZebF/UEAk/uR6HNYP/Bd4ugOQQhn2mBq4KDtXbzAeJfh
XET7MTbHuXMNP61a8EHs4716plC1HoOwCV9N5MeaXhYdoSavcprpPEkXcVIqXMoakMDeksvoq8VL
wDykLrwDAAtsaVpPNUo6jQZQMJeNirJ2KP4nbr4Hg+QKlNG7qhOT4qt8t84xNYSai6RJRM+jyWQU
wNK3W0Wo+dIY4jWcw6f64a352+oeeXLARMrMKRP/es9CkksZXxeOjPvkermTIg3MIs5jx2dbK55+
DbdGSOe97EmADSGLkM8ttmFo4LXBxEqjqG+DZjrEj4g2dNzuDGzcLuSgc9ZgmHlhH4qXWgssI4vB
zLuyH6nKeQpuozH6rwRm5Baw/posJ63LB+yT7LeABnYlSnHfDk7kpG50nPAOF7LmwSLaay6U+wAJ
10N37v31Ir+xV/gc5q7iTBy5+/zrXik75osRbyEf5qYNDRWBwYR7wTTgfgSESw+6RL7BXmuqpt//
j60ktOB7CYKcdFjazBnzy6iJtU+xoSacgbdtJevDEkdnyCYF5eMJG69CkBwKSH9FeC4zz5L9XoK+
YkCudkcaw1sNWwR1Sbm8ntKAJsmELizl+ArTo3mUy2b5CP1PCcHzs+btJzkjt1FEtzUm+DxlgXZP
ojyVHXUuGmCMvWzDpEC6X7wKdVYWDcHoSilW7m5zgKQA4pvWSvVwTZQTQIaQ7JpfjaxEqJrwPHWk
Y26fB/NOT4XayvLlHkNZqREBWDsTMFX3qfm6oCeUMFcBc4+9zdbEVmMoU8YT2Se39Z/4/NodT2r5
IhR+HWp5o4H5c6kw7dM0uWXr728X6yMn7mCJe8+8Vtl58J8RI39fkuX9hle68YRLRglA7a6MReK4
eYdLsyRdE86sU8VPafPzASAixebKxCLF8YHgZo4Dv1UOGcbd/NX8PthWdCtcE0Cculz3MSfnnjT8
2xan50l776AoQQ9XdG2DmlvJEoEGSE/lX74xxLf+n/pkI7PbbQ/9zw/CWCPcFJXkikRXEizsjAyL
y/45/p6d59f++PIv7UBdc881UwkKFBixXwsilaikNYzNFzkMcCWLyQT5vX/V5woxi/Qbz/BQn9ez
SykwKrvM6gStgc1lCWEuWwIncDpp4Q789+ArcOXtHABLq+oEUkxNeiG7fGa9C0UelFL4L5v3v+CC
snHB3WDNSFmKjNGl7VnKJzG2Xcx+iigircs+tA7uDx5YzVs5V10VUxkSbzAf6dC6pSahLEUfIDf3
h+E8dfRndIWG1gvircIMYMq4ZtiqTq8EQovYmff14FGCeRAw4Y2GaYDhImFg+suPs+ytaLx774nf
SiapT0lGZfNlw0GAzjJqlhbQ0XJC1WJllr++NnDkOPMN1eKI1IWh0T7mAs5BdllkKW4bcpybRR17
J8rh4PkE23SS4a5kcoDomEhxitys+4hxjEZA3vopWeVaE07huiSw+pDEH8ufr931csanqluY2t7e
QfmD7mPuErO7rI6sioLJuxt5xNz8+KTI5Oq1px25Pmzv+qmR69FgNCo4W6sskXbMQVod1va8eqEP
7OU4yjdJR1NbuRCF/kXGhH8cifDHQjVZIj/MbkPkMSeUlV9sn7DF0EosFQEHSuDKn8OU78+3iB9H
qyGQrZOibhV8ogcXexrARj1tIgLhmd44WLIHzrK2ZnLKLS5iT4gFSFbjvO+A7OrAZcqWkcJK0p08
stnWLxWLFIC686pHaqDotngKLE9RRuf+j4td6nOCRJ2myEgebfQd9fOWDIvdUDbX6PRDIQ+WMGty
DnES4NGguPNnHSzWf3uE8Q9SoSnLcrzkYF4aWwUnedaBg98FaHNo49A9F3mqNnEGRg2w89MdanLi
wYc2/NSEpQYQsmkX/1PFfc6qNQG4UExw2TFLHLHsW7ztmvaUYEtqMm1Owowd29eoznE8Ko5nJkLL
5I2ViYoOONYZim/d6OVg8JaUJ9dC6azF30DLArJoYxtCnDv6oDcEGqKKqJKgqgNDluZwFKG202pf
OdZVWpbubR3u3bIpI8eA9sXZL/M9jJvQ1/yKLPxcIzxFrIjMFYvCJMY4h0KwvsI7IaX6weEtaUco
hZ/A17izWKbewVmGoOhHo4PHBKmeEBgv+v0Na9sQ/VM2hPBureDqXkUoXzBc6ONclz4wwJnMluTI
Fw7A0lTzb3HvBjHRwgcrDz5yqBNb1Ta4N5INfu6PEzsS3l3p3c3bGRK20HJUsWWI2fwsZJDB22RP
H05G1lT4lSrMaQNPsHxEkI2Gw4H7Zb4m5agGn6prk63ROJeh7477FcISCBiTyGxehkt99LesU/zF
naEfjpcFdbYCHFn3beXzbSrPEFtiixlL7o2D9wsGxCeHVs7Hw7AihAtvvtiRYjVb2ON4oqZ8mvbA
ymwSjnucOBQFOl90amNmswNAWyNZn0BPuPCGR/VYz4tWioFsMrIpYxYQpn7ID3IoR06Uk2YPAsZf
Fa4KImHclo2abgKIHC1ZSfl5MyyoRmSkooEa10m8X/r8r2ROxpvIZ5KELbQY76EOuPeD6KBeaIE8
Ur5oxho016vSL+QUhK4+luE98txIqsuxCy1fZC5YzdP3kLoMiQWvtItkYVIAd7j3HebbfFohAvTY
fZlth9RAfQA1OdWdPrSVpWn+RdCQkw+rVbE7C6s7tGWysyxyOaYHjaYgYzZ9EtsY5Hllh2rWCyM/
x10zqBwPagvkWw4aDFe7NyDXJ2e3419gHW+2FpoP6Fk6uRgyGgWBwH8wPIhb1SxO1wWJufS84PIy
AfqwaQXJE3kjv6DRlObyPJiAs/psis9iQtC6Q736mfSvVSmSEB8PI03n5o/BUJtSpDtm0dJDP67h
HEVQyojY55zId0mjDCZg3n0prNttB+IRcoGfH+umK3FImiZyyo3bPhfWZNcuCpcoOO/SPVwSgyfv
Cy6x3OFwNmKbQjSL/cPjaU6K+ibG9ZVK0oiykAux5JbeeEW5C/DEAuAIwzsffZ1FtYiCiVoHdzZq
qiSYfJRgTxNOuf1PVyL6m6ogcQkeqIzARlJtr+7lBXI8pgHmXowBpO5IQgkLgvlBZ6jCeWt4nynz
TdDIZ4uw20EmaGOxDVfurpVo2ZxbxWVmH1S5JZHh8H+8oqH7KVniRTwhYvbi3hjqRb3ZzJbogwZ0
FbUhDpbaVeojJP09tyHpm5tX0WVwwhbBFqseXe9tHERVuJWdX6KQO/+mgtzNqUTCtcaRYIkQ6u8p
EtIsP+0MWfKmyGuS9bbYFICQa2ABXpWGwFg4bHm7DImqsq7S8N7X3e9C1KtSatJSpw9cZDWYO5cm
vusMohdszPkLxAW0KcK4Fcpn1auTiJE2TFP838JA3ex8Da8FkWeWUwHc8y0DqO5U1RdvXmdhF/Z+
WF4H+Kba8ZJtPGjtmBvz1XNBTwr0JoldtCuUuUeiV/0J+d0ezE20wFflizx3pn8Ewpq8RCSOMMQ+
iyjGXfM7ZnapYtFi9lzh4iniclLYuZDRaJ0YFO9cM+MSBsDUOWNeK0ODqnWq067KqE0yfqysWPj5
fkh19XsnAmYQdE29a74n4uGbgMw3p6c2BBSoLCGNuu2y+juryPuqRQLtK+O65oG5jWtCHjDy5MoT
vtdqol5vXN8t1Frpofq/Cg8eJRBEAIGQWbipPORdsAIS1uaqfX7g5DXG+qRf1WkoOGoXtlA8VAA8
lFvhiCxQVU791gFQBZO3jSOnESRpE7RppFSM4yWgxvs4EiYlFnqs2n32HDsB70KtYi/Zt2Wo785b
sLBnjPeHdfYiXGXaHqxtrRptu4ZYPOzhkJ0v5zL/F5aXFcT6EhwiBLyw4AQLJ0m1mZT2G+6k/zmA
y8vEBzIgmzK+LJt5vbUBH62mozX0elKm/bXsBpRKHonScuOQ8Rf6kWjPCj2fpL3/gBymLOV/r2Bj
xSaAS9FT+LQ4ZrPVG0NBS+thHTogYP9kGvMTJu+yYil4sopAgP2aFwTtY0ynyuI/sQu0uugXRyjm
mgsaeSHN7IFzO/ZnJTZ4dUWWy7WFM+QYAy2zf/8FeoBhGP4fulyvOM7yGws7OLtI5LNaLjeyjS7a
iMjk7Omg0V+uDkf6VAZiwxznQuZ/+YYqJJQ/MOnO1RNInGqyMLexa/z4iDrDwphYX6Lnbsnpd+m/
qRXOjorp91ZG/qjw+cs3L3UWdMxcbypqcA5THv8QqWLn6OjIZDia9XgHQdRO6Z2uIRNcP2jW86O1
+2NM03Vp7ayej0CI82JZds4LQc8/QB5XGh+grvBUSxgi86JdGIo+6Ie0uW2AIr9WRZ9NUQ7Bw9S2
U1Zgv8Tl4wfNPJZOBNJygK1z+tMF2oe17BhZA7ZhGubB8NkXUBAwhhRz8TlI1+GZFAGZRAtgTLIb
Xg4WfCfcOSGyWYVaBnyuwT0BKzJg759rOQ1QQwAKonsS+eBPRSqT9gBiphQyen3upYPtPjDcYSrp
SWGPo68vfj0oMrL/CmRqCCTdQXMF/97Ta7XPlHU/QLi0PXrLNa96SS6m9blYbvQKO+gcIJUe7jp1
ILyi/rjBOp7lmvFKoC+PhgsYKbqHqkAoLF6rOkxRaf9/wfmUFngb/I4ALfodbTWfDG7Sl7nLCLZh
SHMaFfjmOQmleJa4XuUsbWYz397Ann+tcS0Zk83mf770UfSBVU6l5Jj4fkeeOD4hyV5zPopIRcer
lMQ4vDMtBelLf95jKewPNJ+C6TXKXXrDUzD2fKuJhvmDboJNzCWD4CiXS+Spl7nCfUCa66EHvvJE
ng2ZQmpbReSgUppbqweyElP1ajwU99UsvpPqjqIJxL61fno7SA0l5dJPbgJBHJdjLzUX7WuaCbF6
5O7DbPcA+WScVwVmWa698NvBbew4X0hp9fO9+rMMMDj8Srcqmkrd8W9BJQksiDcXiucUtXnvAvTj
zwmoGeUrmuqfq8yBQ2YkraznpHEZMLZxAcOjWsIa3YOmFxG38Slp7AhTxHcpIhCALYN7EWaKX/XA
8tUzSY4f92oLst+dPSgQrjzWTNcs4a95IOBwYP1TavUpVx9wNdZOxoGaMx/WWygd449UQK76z1E1
jB6O2SAH5iNFcuHYj7FsnKITWfBwuxNSb8qy4lYRNs/SPCHPzDiacdYDmww079Qyer8VSndgJcuh
0XKsVmuVvTTqlu+ZHTuypQ0pEgUag0GFa1CjvcB39J8alTUml5Agm7wOenZDDKiacPahTon3N7RP
uXt6DkOqXYVa1fAHdQEug5K390yoAPHLJyCw+/jE51D6/OJqmvONtIHzlPDsCCUUj9YuLFennKmj
i4n55b8Jx8mnY/FvdHAxahWrSeS+I6ZCOLgWKb2OfQCN2qP73lMCLVTQ79iC5XcyjiYZTVqyHFmG
t1YFbLV1+EAz0iZm/4W+GZpALDlFjmY/PZLn81cQlt+ybt1CwB/iKXx1SuoKLFchVzjrWGWCjM0E
dXeJIGCKS+It8RRwiSuF19PE4uIJGfdZn5fYcKLMayCBix+EzLIPKId2DM/B3bJX8dIcufK0+z29
QOIjMTOpM120q7wdl1oGEWoyn9uMTI2FQaKaVlCnSrTLzN3/JCHzRbP20rGV19wcanxk3GsRK7Op
gfbQ+Xm5mQj0PKf39GvLrhADJICy8xLUJY3q2zbUZ7R1x+X5mt0ODKSiSm5YZzCTOByL8NKoDKDK
LoZN1DYTg6ovGkgI+IiyecpiiynXVV4hiuLCiuaok38RMTP8mfu0L5v+qn/HuW7R0RFOWfMQTpfN
hhJD8Ip7ndABwrIQgI1FCIJxKIjamDG3/Pw+5rCp1V24knZQFU96w23/XZWnaC+ZZPViruyGBira
j3KXMmZzJ0zpljckc1U5lqatDzu+GOqhdhVnIH3CK863k7YKKoWt8QfNiELmhtEkCrL6w0sXLDdr
E7VSIzOpEgXdxlB+oGq4MoHk/IV4OsiRei3BNWJkCIl8MgOrniPzOAjFVDll4x82x5SD55EdusaT
cbwHsfDKNCg+gxdAhjYNuA4kNTGP7KqLx4TnhtNygcWl0zSFE8RS11K860D8bH8xUlqxCRCsW7qA
uYB629gwRRGFFUehaa/FogIkfgtZq4XJC2PdjyrHMaj9rLZiv3rz2SeAKO3oc/tpNsiB63qK2Kki
avMCzQPZqx63cyD2PuyuMLCzN2X77qFNzRp3Ke4mZZZ9Y+4Iaz8gZ7HlPvnup2HDcO8lfQXetNbF
WTdKIgWGZJaDDMRoJG4Zox+acgcRgokMjmKzLGmMjrFTtOFCt0O48VBGPglKnE7XYZbHrTFm6s7j
6JAevF20Y6XZL5+Y2QQBbjwCSkSHrkCSEOkCoC9MfnUgtOr5WcBLuk5GKDpLOIzQHNJvZvBZ4i9F
pZulJtarDu48IJi6HpLyFfYT94l3CSYUqi72jQ8cu9yJBg1Psl0s2ATP5OXqorbrDFEprFCsojCI
krv2CuqbMwFqo4DnmEpELJ6d7aOUMG8gob3T6Un77YwDsQQWJxDyx8aBH8vWfQ1/Iz/1hyB3pXPw
Nrkl3zL0HWER0Ln5cDDBrYWxi0UHIICtBM5YCS/xbOz77ae3mTgmJLLOLnTd4fzIMvmLYQAqGXl4
5R+nP4O5BzUInsLkJGqfMFWKXoAblbhA1iiwa0Ps2ldhYaJ0924cwGipGlOcV4ZZ7o3sJHEyzY3W
w3gc9i4JWdWnX/MXS5v6U2+XEqhVfACu/nRkFmli8w+nFqc7rlfeF0G9UdhnOFhftt1Tdj3jZyv2
oz1El3mipxvE2P+3mM07UHo2Dr2VPtsul8zPE9ZZuy6JcqVpJNlunW9jutQkQyPMEx94i6dIDTnk
wVeSUQzxE85dfMzQBfZdFtGjUBy7heA4qdCmnNl3OnE8f6Q1O10PIKR8OITEWrshKVZuoNU1nnWZ
PKP8BTCuMpMVFyaA7qB/MmBsqkpcxvoHuTyUq4enribpK97s7MIz1SiHddJeR9vibjFeW+RFas61
h49iIiXa7YFOmRAYKLlO8Bm2vJGWPlyskBQazc50GViK82Fy2y39tHnjok4+TSX0Sr5t9QyMJcjB
xNtQDi2SzPD98INYDACPdQqG2JR2OhCViyoguUTMIaTKTtqEs0MzxA+YfpUwNRrSRtPkvOltUorf
JqFNlgiXEqeFzUfzs98gCbobXYf6OZkjaSQvmMwmnkdOEwxkYt+me8g5RR2uaJnwnV+EaRhtg7+X
ui21j8A95rpr0HSTdgofLPpEyc+/Hkt7NFTqpFn+1bPiJDSIklTRj2Esja0ol0SI3ad3yoMvvoED
YtHbtWd8Mj7McfwVo7tYPQchgZFD78iSrXHeHG1TxBFltCuMSyRXoUht2n86DZFajet4aRcK+f4n
W7M2FcT+nrJrApa9b0PsOZnpGvnjWXixcusXp8JduyBq7bV7adDsDHV9Mn9JPYF3SgsrVrdexBU+
bs0h+0Y0G3ma4iVtw2T1eIKSwB+OR7ohFlTYS3i6uKHkoL0P0/Wn9Q/NsW2bllWNnBxi9FVd0A+1
W0crL1OxHLSKoNxmDAfpJQQQxQ7DDBKDYmvYnCzhmEc84XvmADhKHYyeNX8kdBI3pG7025Xa6cdD
FY1A8cHk16vV6DfEoqz/K0ya2KQqBhKX6FrsSOEQLDXoDmsk4dRVhoyXLLuSjJHjz0RQKqL1rktd
kNRA4p+nbq5zuW5Hv1Y9vpY4a6xRw5Ej+UxncNQXaDcZsgAGucFZgaI0PY2IoimnA8ruVxKNs1p7
Z39eYXWl7xhf0o7RmCjvjfk9VfVH5KmNxDkymA19cGJUyuOf24XQwIXgJE5JiwOWlu3f1Isu8msw
fiwC3/UlO71+1M2c1+O3rQnVZPa55ztuozdfAOEJMNCzxVmoa/cgL+rAno/prdhfb/xZ3f9JADTQ
M0C77h5iD588+xqHPWrBqn0mEUlYzbC4vjaBGcdnFWU2pbjY8pN3fNwyC9HH24s7rNckaAWrJtPO
gg5mZ+G/5PQaNpyjMrzDq5E6brA8Ow2D7cOyTwaNdYBNLfLItuDzguSweaX9eZbvVlX124Pq3WOE
+8WaG0VmpECEk2xCsKbBoPzJyI6PsC7NzlhwhOu9j75KKJghBwGBOC8h6oUUvj1y4tn70AnDXfRp
ZMlITV7cYg/ssHFN50A4v8h9Et3SM+5uUz2Qoc77MAge1GYkFh4iKbO3R0//3ORiCOJIyw0gV9Q4
ds+vE4YksM8uevpAnmSi5FaJ3n3wtV2kUJYjqTbmBbvv188c/Ng3I4HyXO4FmmHLiFGKq8bO5Sv+
cZmIIemPUHAFjHCWf8CxEz1AJIudg+sN18m57uaV2aQKAAQhxFUZzl257OcwTgD3I8QQTziRuXMb
Ka5MTX4vVDkMpLNRAXI+R4P3Q1FL+Q6pkUP1p5kMaBttdXqiaZORxydCUQCdlGcSQEu3l2ZqrAvh
t5+D03qRElNTGcvJlKdHxgg5OUbfI+fqpjHcKBx6/y7Stp51JG1qk3+0aQKnPOBL9/LFbu5qt3/X
hpUfOvoHfU0S+IdpFiXbsyO5Rh6spv/vSmvrl4aSXQgGDRkoOI8EZDx5pyo+IOGHz7uFMpO3ZKiK
lRBV+zJr9kRjXzrJuZWEwtpLVaVjwQnuxDHOoWKrRV69I3gTYWIIVO6zBEkMjVPajcFHfax7JF/o
Ifh+N+wSaH55O3tkyJAVA2hKksn4y50EI29elatjB+xiwKBiiburmn9A/+osqkhtH2vChmJNv0SF
KTjK6fw9t4sCOlhVMgC0GyqeFR+OMaS1Hh1zTnAM9ZMW0VvVNfum6diLYW58vstFLf5kntuScAcw
PYB3aiDjCpY0rv75OFmT95Ovlk3oj1e47uhkE8kLebNb/3YA4bC1SJesHJuKWV1iflUUiwdDPHyq
JlkwNWG4X19kUlOs2G3roB7wUH27XiRexbEe/JU5mQ8aJMQhpec+Y4t2q6vvXtbCwcGQw0C0E6qQ
0zjG0pMo4y4zbZwZZQccl8e8lnyjq6gnS4ihjYHfQQqNt6h4iLd1QGAn4dRWtzpRBqrJ5P/B02ES
rdLUSuHyesppbhRXsAbCts9Ice7yBvQjo2wvXYYwJPwDfBEH4uKQbJOfy8zkjxbiLq+MANrdFDWF
AltwDpNhibiuFrRnt5P+uPq/ljSOAFjsEelIjFDues198DHi0EkQe+rZ2RzQDy6Ys2aNEwxNQYDl
jpeDC1SF0HDbAx/CgODhotHVMfXctky9a5a9XsCi6T6dEFgyexCrSkZhFwihSMaJklXX/aNLoWXh
5bUV+s4tdWMznEGK183rdqn7XJRXKvRSiUlXQ/A9nPLyHkLcXr+91e4DtGsEBSVueVEponpAyUeE
Fi331hlxhAL5kHBOASwfd7pmfrGxbVN/UhCOz5XSS0K8N1aM0LFK6o1j7WcL/1R8fDs81Ubla0hL
TzPBX4sMko6+nq+5wkR0Nk/pR5WOPFIwX83GfXpUufr5aWHUkig/ylCpjXpc7bEyTkl2DDE1NhWK
LUpOZ+zDLCUIbpS78vSFksLmvhtaN7W5Xt86pyLg/ynAurBnr5htLhBKk6FYnDQPNuZq/MJtUifV
MAl5KSRcYcbusQ22bJWdPhhBJexaukBlKKbJLZW2NuR325njhZl0pLQPjs08HMsxTO2TITi63GLy
C8zA0b2Q2W7Ochz0kGvDNYnXpAuuJgT4w7I53jhc+vRQgqPuPV7zYZ/loegJ9YgWyM9SAf27/TPZ
Pud7kVwD1w9Gc0Xpbf2jACoEZEfZMPM9hdckp7cGED8Y4/sg0t3FSkqcP6tU6Oys45A2olhS0rxd
2Sj6fW0oj4q2xMoOvIsCgbekNtawcA4sJhn5xinGAKYsUZeX76gXKvJQWZOjmqJBqlc3bkk9eOyd
pAzuPUpm0PW+aPGnzBcNFdD0RSoNTntPtyyez5zaXZgnQTMvSZSbZ4l+Kxi1tJfHU2WUBQwzXH9V
M01t6KEfg61khDF6zcC8dFCHHwzHq+7rq7auOh8eyjzHrxWbxW3b54A+tcZWIgeQtKAhuJKRvk5x
6xatD0gTVMq2uIjnU115mMeNAHcGjAJworABTQOi3j+APuCUxbqB2/6h2+0O+cqmOFRN5ZWuKZ3a
leYJEXq1KZma/HZv3VZdhfoDvETMCO1/ohGGPRTCOO+keNlZyQN1wgclB/XpO3S0CBChAQv0nm7G
HL7N+TEWjrCwo8S+QruULWUKpjGVGDgx6c2ekIXjAyxGetviYgq/kPchweeHzIN3LUXgp6NRItLS
ogaNOCBo8nZ157lnCnS51EcJvkB07jr1OzvSe+bBzxUBfzvGo1sa8jwuEayqXfiSF+Fj0OqAfg0b
RTP0ZQGwvsjd7nLtCnMRx0NQ5FF9L01q8Q9e7ItTaRh2JfxeFmuaIA62/aLLYwVki7PBKU5W6kno
59dsmnJjbB9PXkfuZaPXgWU9wvfRuoxR+XIoQfkYbG6ghNhyxvlKoxvHa+EgYZzMGSgclO8WkLbb
s3bVMxZ6G23IUQTzeUFmQd/za2ueyTP5j8LDu/uL8qdrwo+/FCubMNJXI5ALSCTPyKurYOWsSLvv
wkUwXDAC+HuM3s+uXDAW1N92bgkcT2H863vjBt05Mc4RgCHwtwRiS+2AhcOPA+KXkxnmZ2ZJlYr4
N+dBnAquVdaO2AdEYLF4Q8tgT58RjUQim5T5pqzAZ4hcZsxMQznxE0u6nvYHiOB/CHRyJV8HGT4n
YxXgteI847dMXTW6wBWKpofMhCZ6X/uFt79EppYuNcT3vrIzIpq6oMNJCjz30dWzv27WvguqUnRI
uwGlmHZIyeuNFU9YQOkzZ8hkckXRcjkoCJzdbIKRU1kKHG/XDI8cViAJQFjIamXVLfwcpRfhffyu
9B6N5ZaebPSXV8OA23k84Kb/ukjfKuYuvFAGJKBTAiF0TS3Ghhy4QnCUTBG0EwypRpmWJCZlT9wB
FY9D9XDZfQFG82FYl+T36E7dLjWEvH3i7ZLKMa2xeRmrlEKcTwAoHWkSFkm/xe2/BeGa8iTysLX4
PybsfoBPuMtrSfGjXAAsWMS5jYPV8m7wqExaAXBs7MC/nEVdvbJGk5ct0ndemSa15fMG1b2hMvCX
I0NED5fhVUAEcOYz3b59/04VCQeoK+mDN/4bX9ExXGhM0GPI0FB6fqqx/nAKxxaYzi1/P6QfUAR0
s6LalkZ51TMxv9RJiMpPrpA1MoaJIUeSqGU2Vhfevx7kJmVARmyonay1QnpFbO92x+xnek8fPAXK
4ITh7vqtLalUrzODpvbunIulMag7CN5Pva7jbglOBbRzVokF1NCzsV9R5ErGFsn8BimU/+VoXKNm
2zPUsLbqrKlIdOv5QijKN+WNMwECOH+s+V6Sdzu/33b1IwTFdXWNw4voBRw+aMAcNrXi0XW3WRT0
bq/zRHmxYBZ1Id1A2sLw/q1IYvZEran4zCoGA7Fy5ejMn0n2gtpeCFEKsL9bqvdfV8rT6mSapQoB
t25QnxBVK1B/lnePOumYdg4YxSU79B0bqH2SlDx8ymq46Xm/G+vlWAK2gYmMg7Y128J+BlwHgVxS
kN2rCZVOcV+irtwZE4US/Lv9NqSF3/zNdypa/uz1U9JnHrD4qMe2TFMsZwaVjCOAm7Gpz78BjuQl
fveFYyitox45WW2DGjqmfSgJ+7MvL2z6me9MYceXoLqN6RqsQidKuNbJoeJUtv2wO3SFpr3VeOd1
hXMeQFpwX8TPHKzLqmqykBre7fX/mfP8wZtowp4k721KyHoeHfkspe7iPEXtKlOpF5m0wJXZP4C6
XMlDYwE/Sm3X1dCULxwdndBvWbsN+UB2Q6RueVDKSoREdsQeiiO7UJSXbFI/3VyDW97q6CjodcMh
eb8trVTP+mCEREkL/tMxvyHXJktegdZ1is9rfYIU3a8vky0R0bCRPoICedokzGPNLg5gMZIrUmTZ
5Erp/3dVoRHyaHTBae0ssTBronfTEpey2OLm6ViQdyQzblEndVf0IU4IcccnsVENwfi038UYpyys
pOI46TefAb3LduaO7th0Gy2EZYhiiGKe3JaK5U9Nn126pg77kzkA2G+1oOrrOIgnIne4sI3J0Y11
Fis2oucdofuMS1gxmIi/+VxubSJ7yob4AHsIXxnGNXztvcwI9tGFSB++EfezBAPtc6iiueFmcyt+
FWT3yaWo80fh1dwLbHI+QScZaVaWMK5QWrHOGAZFuhvF+j9BO057KWHCqAOLxpWkUqG2WOfVuwHQ
IVve3ZP+7iXqtZkkB/JeEmedoYebx/jbMr5dhpZR3aK5NU+jR2P8c//E4vLejhZ62Aew7VgOLDyM
MZQB7xs+N13FVs3no07NSjg/xsJQ+YvtlAvmz3P84bRXyocGUTMcVi9WyDduu6Brju/IiiAs5oUk
awsX55kO8xH0585jS3TlNpzukkvr7AOqftTQnA3ad85suxo8w1WUXXfmcSyNYqj7sP6rZ47GDKpq
ylNjfrrdxee4SCurrnRbtqjg1xOY/Yk5z7wults9mwxOD3g8l8uepm2bY9nkT56ZrYr4hS1JDlq6
PffREC5vU97bl+HTaxi6dc0wNe/oYUoB9jDzSn/Z30ht2t0cbe6Nh2UDadA5eu7Tnldjz1ECpNXs
s5iWNbbd/A+9hAyNrZFq5ODwlV7oVjJNqtboGW7TVbWPWJae7YiYIRUOk9IUNRQZd25l8e/srmTO
ih3Lxm5AsyfVvUT9DLpiMTDadGp9pOy7B9sv1JK8ljZpyy+ESzCX6Z47XcjwcypwPZiB5//gURze
RrfQ97O0DTKK9z5aNJ3uhgzx1qOkbHdIgBuoDkPIlHJLE21zJvlnW7vH6z7tR9dQKB9Dkj1PgPkW
j0GsKZUrv1PisIqhF66atgNtG9HuYfcadVuMsGQyZbN+MV/6MU3xH3mPumiRQL8mPozrwT6dOtM7
sacIFPJGv6swpoRkUeOERiRjdORjRaHPC6IWTDoI/vcfFIxtRj4ZUsTi7FBpffOVnS2H+iLyM8BT
8uXVfiE/Wb57HsxDHjhxKjTcbQRuoWcwQhjXYPUruy9nqvQU/T53ADCcRhZDHYN6IAa+EIruJR7G
kP9yQj3GudGOenXyfgV9S0H/edPAg9MgoPcCPmGsd0EUVkXhrPY0Wse7eLXOwWe4eLs+kWLC0RRI
BVSatWGp0mtjii+NyWuIN3jr9nczosrshqUE6jdirTe3b4gepQlYnL8hbtzMOCovTIuOA3b3+VcA
uboBrS0wDNoK1x0FjQ3v5tTxxSJpg51GL3hoH4us0tH9bqTjEDD3JBDni0ca0lZERzHe+MBWbqfB
Exz8cUNsd6Bu8RTJ0lSt/7O8griQFUbtpWPinKMrkhMqKc9UHZP4eS0XlBo8C18iZnncSnfjLPKB
MgRC3rQxmhVmluNK6id5XDmg2U2pwEBC+/S5mMOllXivZRo3FTY3klpGneALsFU7Tj1j0PbzxL8J
cA6qLSCKGaa9i6RWiAzYMdyFCAKI7L2r2+2MfKHjYGfEtMJtNpeNWmqAl2Lbh0hnmej26jJn10pf
7GC1pwvVG1oObWzi5DyuHpJCohNWmRynL+4Ftp7tN0cT3ZiMDE32oyfHLGM2ZLVJLo0gnq2YYU4H
A9PRPdiHOS17imOhes1yU5Hg9nlNwXBVH3L0XWtuM7idBJVoMn2uZhJVGP3ZIeuIRGjH/d+wNmKr
FcHL7NROZmyH3ICtY4N2SqA6h8xQQchiSVXJWDg4ShiDFDFtdM3vvSQCFy4DAK2rulePVQA8ULzM
8yf+sXjfiodNBoWIDSt4XvumXUpGzEXEJlzg1MCKYAWh3d2C9ZsIdptpX3UIMqGN7derdsJrwU+o
WZvHLK6SuJBzwifMrO4IPnF2VZInfGQQcy2mXRI/wI4wtRkVxOHKbGHSoYPdD3BuxTnWBi1tHWMY
l9O/eYiQwF1VHZjKt08yrW3w9a2qjbDRChPskOI1FfYir5Y4j3lt/+gIkfp5z/eAU/AZqdmE/mKX
2Oi7Z9m7YfDb4xTQsPjCKaD5ayN1MhkLwk3+9PrALUN8pErhpRPpkES7+wxRjilOZSi4m81DoVra
9HMqEQHV+fq+7PSqDlYorxSzlj7RYY7RLSvj5LWd0K5opI6v2SiSDrjO3AFopDZ7Lm6SdXdZtJ7+
xz/6zQOUSH28yVRI5lElC7oXPGAOt/uFYer7sp+M5gVSK0RtaG9B9c4wnQ2ZS+RUS/iv3UnMtz2b
NCFNuL2r4BuDoaydTWcNVoNjBWYANu5UCPLuuENY+wkuDnO/aC6UxK2VzCy3hnLw8vok1BHaXtax
7NtXU9fBmHSep/iw8Ede++N3OnmKP3sc0Je6PHddeszXj67adQeIZOfGVu3MeA54/MV3BmEnsY5q
yhTsKhiGz1obVRMzbCBllHH3OasVQGE9QSX3AF8Ztz0F+TdT85B1TOmGNH+mhubEVUP0SNeDBoZT
Dz4Q8oqV2nhroV5QSiPSvKz8n7IIxVTFYvCN0BDikb3kJYZgzgMYtEN40GhIoqanHBKi6eLdxRVr
wzaRSc+BJ3VPmPqQsFnkWk831ibSFgfUpxRcghAH5PnjYTtTxloKWeire/nIPhGlnh60zkV7nwO7
erB5WAkp29wWvDyNjMCqsApxHYd6N7QhGRhW1BFNEMjCAMxcegwF3zyPtMnzmA8BSxxJ3wH8CtPp
eI3JwNY9zTYOJozAUZpS25TSaXoYiVY5V87ag1LB7tcqgiUAGa2DHtnk5Q2uiZgh9PuKedh16V6X
jmwQC7bw/x0j60SxWkan9JC6Zy+1YwhovuTOdzD6OlS+opCVl6Z88Zydobtq5l092ELVj4/SqK7l
njjMTUxDj4henEC5gudeAAAbZ99kmBy6fa+Bb5m3vjtusTdw0p1AWG1wf6YT3ZqmoWfdAXB9w5Zn
mjlm+XUh37cReZCv04O+LUdHIqiut17fN+3Ekm1vJ4ySK4fbfBz2dxwcl/lgVD/4UdzB4HleSQcj
s/jqkZcx8aMfdAf6RjPayzfzYRn4uW9sSpz0J7LwpSsrEYJ4NY3VxyUmsKWh5pR0wMe0lhCl91b+
bqJT9njeZ5QJ0kyYNknEAOrg7Mv0vpFRrjr/BYp8x76fhbRMay5IC88Ni+xiU9d5PQiQVHIzdXIs
B0rjTwOGaZLjiLCa9RG49gNsgh55C8mtpjCxMCROtkuKdnFKTxct5ilG06fRShZfxoclO7yivcE0
Esroy6+6fVMNJ659v8L/YW275cNlePxg2QFflZAW2oVpyz0M+KSg0LBg/Oe/anAraR2/FSOzxO+/
VynzBRhLV1j4XDQYvhqOmIPn9WW+OoRl2SAVOZ1A9TCc5SOgpAamWnYxubCrtF1JqIIWCybj8bpr
RdsysdzBOr8d/Zg1FDG13nw+BAak2KBBrQ6KQTvkMuiUPPWVptX+Fz07TdtcCUA0RM2E2AiCOhlf
uRESIWoTYVLajSLJTp7mlMOaG4mG7T/qMnr7mvpUKUqH01h/WtffVDxesBk35wRc4OzcBbyKg3ic
CBMbqJMfQ0HRMomqpc1Ctm10PqI+PJ3PbnSZju23r9TGMYJGDBKbqm4lWfnzUWeIQdkMhQZn0gAD
YBJxGq3xtJo5ltKx1pKYQ5tSNDvjrRxh+8KltWpuJGt5K+MsxKYRi/uCiqt0YeasjMIjrxl4oLkb
Ci4DbErhWY6zLJ0ZB2jZvvIdYTCrSxFdh9CcUeccLl7nyFZ0VF367AAB+QuQRJtVCP3TnScfSObv
dKXnNS+VEoUaZV0V1k0Xkl+fTjUaGbsS7+52UrUjE7LZe38tU2SpQo1XHHA0q1ir8O3SMn7fXRGL
XJGzFqVfSOSEoEwGh1mSLihc3TzeRGH/7Hg4+9kps2x3CA0iibzxpbh6Y0Nuikegkxi9dH9SGGxk
44486bWPpzO/2QW1IuTeX0/iNGZOQULaZOR0XZ5ZFk1ShOA4+/eLVfwhVwDYtcgK0cO2P2FpebJa
nVzD+HUdUBUPOZ0u8DzXT193bSmc1saZD+Vw3j5N3SoBRi4uDuzeHbNDZMyQ1XVBA0UTVKx2sKlf
rvpWiddsqHT6pBPvnvAPCNSNiafkZLaZ2p9ujLEjH16uQ5JQyGoLyCocdnMpPP+e6D0EmpSUhf8U
DZHM4LqxDE0lzT5XAGMJFlNtfxOKrVBKvQpu62OuTEXbD0MJ1PwJMskj71M4WuatlmpGJ08/de91
QogEjSQHKjzoijmvB8Ag80Pyh2MAmURcsF82yx2flMu5o7JUH/ZyGTL+AzpXFsx9cYFym5KtkGZs
S7Y2fQWAaq6+pQf2nc6nbC+MixrKnWIGQt0KW2GK3Nw3/Z1UbvBGQ0ON9ASLJkARk3ip6FHUoOzo
pVrOVZIFGFHFHEN6RDD6pUh3kTXYH/C8evdzRcHADexp4dneZ0tbSP6lQDM2QbbR14gubys6giKW
yt+2cQpzgJydIzSOqbnfmg18hnifKdZwEBafv2Nq5ifUR/8uxsF736oGS9itAsM+CGS/G4PzlSyn
QxAF0VnUScY6YgfT00iQimYKC3IYu+I0TccPjdGSrpz2nTI7A4fRCp8tikQvOYNy7G1l5lv8DnPJ
jm7m+BGYQx1nkQYmlvwayqspwPeGgJK3cAD1qM4GAukTD8UF3WdyXgHr2o8eKcqt4GP10pFbKEQt
vKtPYNRMmKEnVp22iDDiktkMJPhJrjWzmvYw51JSy0t6o3rZjnL1MqgIsKgYVh21mtTYfJqB17nv
eKhAbAEMgrpyrsWH0T53WuiHBYBKUDTkKF2gYSuZNGtW3Ig1oUfPMvzXzsVMoY6DJk135XKP+pPw
bbByvp4jsc9v0ZgemQcY9OEVs9xvnLfZnZB5mJvL6aOJgF1SXI+PLcrIkugltO29Z6RNPJFoJrOR
jmNAMcNaVI/BTSaviPilEBl3LeN4omqrB/JO514LIjkCyDeDhnreY+uY+hulqaB/AQcvH6EjDkHz
ArsvQtSI0yGc8DVIQKu/fquyuOfp6ATVWKHK/4iwsxAGoz1K6MbwzkOj5vLfabD9qcbZ29XnsYf6
8BxGeb7D6CoVFd5Zysu3XC8xqX97KSY0JYFk/iVs/2DawqDd/fwRf1WwA2GhhLFYXxVHT3cGV019
jM7wsPzjiPwxdGywYe0G0GR5BBpLwBFexWw49wN+1Nn9mlkhuvUyHryYh1j+gfzaAsmO7zxWbAWT
3msn8KUWh7ogSD/WbA1XX9cPsGThP2ArLh3sjzQbJ961zBve/Hf8z8sWQR6pAMb/1Mll0IxXTm2b
GmKGPjcK5SdjbOrvIZjoa928z6VdTge80AvcYQmmqslJm0U5uEGMaA5Zi6Fxj6gFgPscAUIWPSaW
PpXZVFmQyN0Tir3A++mbPly3nYma+Jl/V0qzNArn//gX63uWN9rf6KfGe3Wd0cdAOMOt9NMob6tJ
YV4yK5e9n5d/mytaV6TxsgVFWflhg6lWtUD4hYuKpGu52bvgdbxgSiet0ZQ0b2RHOkKlFncyvNZL
zWQpzlQc2QWA/wbvP3YILyhPa06Rl358iWjNgZhSsEyfkzAzykFx9XEehY9L2wq0yUxfHGdw4Y75
qdGZYEBlbloXjCH7cM3HJbOciim51+3L5NO0j9/KVUSBrDXGZzy9BkXMzfxAuuEqmzerN19J5FGK
j3smjgazHM+77MTanlYZA0HtpMScDw9sw8RgRWfBUoC5vgqsrQorHP8ku+8U1G9lYIHRF8bVNVtB
DxQFwO4z97FXvp/kUQL0KnkDwt5gR7zikSfWD58BEPZ4oOYK/EAJP+dCQsWaGRh9VUXQaOc8ZRt9
18QgKmQ1bgEAB5Nk2GuwAzo+92/NeywfnwakJIHw1azOYacjdmO5enoxYHz7PNh/wMLnDneQy1Wb
yvDClzo4/k+A62tr4hEYhr5WF3TA55wzQWE946wdPMZ0/3bfY29mgtqm/+5l8O6BioPJ73ZySLgQ
O6MjlKDvz94SEeUY0NXn9z2u/4HGIN7H3qfiQQveIEzBksAd26dZvI+xuxvt7wY9pjF5KMj1R68C
K6Rp+7dK7RTmQ5DknxJBWPMTDgINxbEBsKI8w1DcWvxU9G01ZVTGYBMsfOGjAtB3MYIV8ha58w1T
NVk9Dw5iOs4Jgq6jzyWw7ujmmjXIkA/Z2MGRoMRdf9GmUW63eRmyl9DzWifTytsV2Vv/sl6vSXDu
7h0DR1g5xX/8FRYftIWF5MaxydWlEpJHpCkx7cx24b1y1W4T86+nAuiWMxWp2F7ioN7IOHH2DtFh
bHVDEASWxgQ47SeLSgmGs5zb16xNHU2h/puhSqt43d54beqhIcprAXnIanPlk427T+01ImMr2vvI
j/N52ac9xTalFthOdKOF1KuDhwLloYoBGqiXdy9I+m6RggURD1vZRKOOIiKVc9zC4m/xSrkiVyvy
MfsfC6hk6xxC4Sm81COATzBB/y0/5jSEVUjLnX6Q8j41/xHcyu+9+AkVBNMQTJwQ7RJEVdINUUS8
fbZhQuf0vtDDL/RD7kLvryqNkX/56kc446DPThx92T3NUEIWLpPFo2sskpF6D6BW9hwB3XsP9UlL
7BWoubjxlEbOKQAtM5DC40Q/IJZ/XEnc606ZiHkexXKVos0Hc2I15x2sD42y6oAWTEUyN0xpnyIm
yHKWh1NL03iHsdHfbBCvyZvhBgL8601+76gOsUWEiUEoZrC61pQif0VWgAupbKaLhEwALOCzigJo
SZCl3HI34VZbheFqWE4Sf3i82JI3ld+ONVlBMpRSs1Ioe0URlJifQ2OsImmN1U4LxKl5wDy6YMOX
+91A4TAAW4bvig1l5Hclbe9Zg3Z/px2n5CWJfOqPJK+aApR83t9WsVAygjrkt/L0zmfEMTzqAqIk
Hqlsf1URHbPBHEk5fhg4AlRniudYrh/z+sBmttzdYtSwG3QnielDuujQCtzHP51dUO+Yo9eYZ0Ud
P6DCzIuozrUfNH2tmDIJQZWtWlmS76csPgENiPUG8ZY/rKjX6diS5I/O4R2XL/XtY9hv2MlmN0jh
UQ80Np0bverBNVS0fTG+ZFFV3PVhIzdH8ydqARhDsAV94cRt70BGMFZzTd3oNxg1IYD5dI3IuqbY
NztTfGzmdyhEEOIGqkSfrZGEIrfOUWcgl02vyDwwKqgwbOup837QVTfjqXT7HuVRiEkkhaTHOREW
3f863an5naXDXLqnbqGyglh27mC5d1mTmivr+xeonQ96erMOFxjQkg0jfT5TKVOoA4EzRciw3MdQ
0lYL/cKFqJh8Tx/4can1sJ1qRxNnXtYCV05TzLdPneAsZR1jCBRlbCf+q+E+NxjAkFjJJ+YM94ig
RLJMljMZggr6wgHaAD81Jf9XHUUOWNXiK0PSel0I8zgiXTHtqdk8zRI8aeEeDv6S8Fu1rsFXqgEl
o8AweHDTj/wIU5KNFxCNnvnjnajbeeTbH0zYc50Q0Dqk3PKQHJETBhkAysoKW6X7LjU7ghusoATL
JgXS2bpvWwcNGWcfamyjZN3wgpcegk1yk+0OAsC7SaWEEuKDnHEBB3SYIrV5drcNmNqo06bWTJae
meslHJvlcGcZuvFShLu4SVYc1FJj9bYRzO+5lZL36rNcFQsB6db55rgMyGjke0BTexVj/M+Pu75A
r+AeMaVIkYopalO7x/Z1n5I8udl5XdRlNOCf5lyv6HfmAl755eNcufdm/9Hjdx5GF93mLbTrTmXW
d71T4ZuBYuBQc4xIkLB2H9YBcyzP/h/AgGzRmFMjhGe8/PasrZVrIf+DyI0+w2AJXSAoH6NnXeeJ
/+nrEzBcaJm3JoYyienvOwrv8+R2WCHEpY5403xXIQ31OQopiN4bkPlOsSjbEFBlb+N2/crUn1s/
TU4o1EVKm50tfkdkUyuT8DCUEVUuxPmK1PTt4x0gg7P5BrzTCvMcZNNfqXg1C0FHJB29iXMKczit
2ZhjW9OvWh2mznsE5HMbUkNHevXorlirIrs93lyOjrTWmy684DJZ+RC7xzz/rpWc+qw3jUm1l7lK
fhH6nktCv9rup5r7OYSf7eCGRTOda4rm/K5a0FuSwe4COmvmj5ZU5XekKsofFCdPNsCXtCkfJyKY
hAMz9IoeX/SFfesntwAK3umhvP+zDmDEk8CsFIBm4XnQ77256BE38yPjtwzaDhbrqkw3N2pPIwCv
p1VZ0LgoMcxeaf3sGaHoqQIVs3lYkl0++1LSMy0XQs+PAUydl4TCoNmFtkvTeT5psK3oq8r54Djf
dtPDFa/HrCXyPy2BL0SlbUHKhY7X0bOixB1LrOWm2bGq6topXsx6Z/6c+WJ3MFBIniONmUs0EH7r
PBYueFjJdlunE+fNRrEMWQFsREKzdWdNJgAWRFOl6xFY6+BJ/Lz1V7RERw1vc4t3LfhXaOOrHW5Z
035yDb0DMJ0NuPdG7AQPlD/X0kX4DXjM5U63RO4uof6JkwD0bDLPXie2vSmq5KPFlXB41fyFPXgg
iWyuuKB5742K+8SSCsdsm36io80SO2Jssop9F1lQMSVP1UMm11eLkMv92RhFj69SbeH+LOJzGjEw
FlGu2cpu7eV63WVwANil8EYkTJodWpcnMquKM02mQ3X7l1Qbx3UoR/sXowX1T47aGhSvinMLw4r/
vNlZhKiPSAnZn8eAy/DGg8OpoU02YjQZ4Rm5nJ3xKuuoOh/EzXpHsGSqbcnTDUjJuaZ+IDv/KNYK
uWDaUDv9jps2efjcRX5n5K5KXOdoZB24pphbc8gIA+trCJu+EuX+K0UALTIXoXu7o0m2okI9hNBj
Qz/YqIdOvorY1W/vIhsXLreV6+gQQNfA+ymJAWzVJ/vRKJOwI2jx7oaRCas1kjURjK2IQfcjI3bD
kqr8j2Ubc95yqCKhPccwQsNNiFpIJUz5c58zImSVcAlouw/rkE0Zya3o7nzzKQ4iFS3Q2o6ihGs1
cwPJLnUMK0Oq9yR1so6H/T88wjEa6Z1FuUC7o4CALbNocRfEhxKiJR7mLWVJDBw3T5Vhr0MTY/CY
X+8wlrmEIK9z/SCsWXRWvj2SgiPR+KKPRJ90tHoWpvHFwueED/uKIHZNDZwqtlg5IcTcoEHyY5kw
zH/NANjvUAE1e3QhpaFwnkvzMGhpAnaEzwlwHyfPl4wka/RTOvx0lVugbKHx7jLL4V71DbqmcTVR
Q0/ntiq/kN37Pu0nxtDi/n7SztIiVrOmZaWW7AhGPn+5+0gBUACOrx8olnQw+RrL0Cu/+wPY3r4a
URD9QJzkIlZwA3wi++d2iqT7DOda40t0+6PSiaI1qHyQb5KTf6OKrBF0QqHm5RSZ1e6J1tNMO0V9
OsxHxqWzLgeMABT10hlIxNzmp6kS3ImkTws1eO0cd4heZ+uVmizUaJDTg7kxRjRK2vmxTvhgl5s2
yyHd9nnaprSvGBob9T8+juHdyL8I0Am0yM1Uw3GUXJ+/15Qw6XeomwM2PnhbuLHDqSPlvZVPEWLp
KNsAEokqSDthlQNzZvifbn7xjzmuImux5w+QK8z98ob2cJO4XGvQBl8hOcj0lzo0roQds3KjDfMU
sv3J1p1pziyXnu9eDnK0tzhwLrozKLB1GWnDUCSwdq3gjPeO01WhendEDwGdbCbVX+baPS7YZJ/z
SEcFlvu4SNDxbm1kMRwpkG0xeczvSu6lK5+f6ltAGecmCX0qhBEo9REzGTqGaWoRI8357A0eTjly
mNWahPFoA5NxUggTQSwnrSJ06XKbcyG5HO3DyfqocLDIMvAIYZLxuX9pXGdQ17nP9wRbdtA1dyek
zJfusUmAvYSi9Zzlo5HP1UhG8KBafOxHnh7GoHBN5dy028VJPEuHOwiQRmVizJ3qKCuuymSEy2mS
0DVWu9N5OEZzJBQB7ZWsfykn3GIwAKvWlKfL6VfRe5Gu0ASEXmPhRDMleiAQ7z4cQGBYgCuWcwfo
C651AgupuQ676UF/XuCiK7gQZ/oBzADaphu2t3gBQfhcWFF0B15GsLBNDwty55k52JO63OzgAyFU
fTwAbi6JIJz5xijVBK2XKrBLavjbRc2SQOotHo9WSSVXih8B0MHI7osTy730uCsHZjLfeXdJv016
SVY7Vekp2qZVg2uSAerqapRR4I/Sww/l44084oQ4BO2Ecz92T1b88tP/7tKHJcF68pY/CgxlS/9Z
vlzNiqyPatA0oO/ApG6r6g/PmVnzp+sTIfNxJjYCisPmOBE/Uv4dhL9sE37BGcW4OZQJ8PJmlxqB
j3KVftcWegA8X7cdhZNw4Zmpq6GejlaE2Q3I5zfKLFZHM5QY1TrRZ39R6DcmFC3cCRgtOBax8V3s
l6MW8+MDELIAdAW0UaEPhcFq3T1wB4J8UkYKPCOpfqt/MhwAA29Jr/Xm4z0Cl4UDtSOx9ERb32u3
wCal5EX96TZxWS7h5oFQ6g/an625tcugauTCKru0KCqneLrpS1qawOR+cEWmpztP4W2dnLMUI41g
svHS6TM9JUTltIdaSwlg9lYBkoyyw27S2t3MeVoyLcuqdvG1rqzNcUq+gshVPmuCFUlBN2yRgqOi
Zs/pU4orxSFvQrTObpcFiruOks9OLCCQeinX+UZt/IGdpEjWURJ64vtUs5eaO3GRIMV1pxbSZLg1
zVCQQ1AoSeFIb0JBRkC9tg9yyS0CB6SW1D1tyPuU8qDO3w8W5fGDJZ6Xt0FLo79tGVHxpCJrx0mc
VKMm/yMJ+opjjJjiiU1Qr8Jt05JqavVBIy13G6n2mqGQefYFp4tdF+zERsqwuRMhF7CIl5Qd5hep
J/N1O0IIOF4lEzxC0cGNbzwO9EjK/lDag/Ytok9Lgafl8wjTABE1XA9UZJXj80O+xExHovTzR2SF
+no5B12y+eDW9NNOpKW2+DFdSZN22uq4XLJ9dwLU8IFFe6ieGKIRyVHucqoo5YlpLyzjVAhBc7Db
j6p0O/v8BfSE4lVUFoAWrHV0fgewiVX/9AQIWGQ0vz5RR0+pDsvzdcvs0j5A4mRM/xxwdyDChiqn
IdrGDrzDgxcM4R0F2vJNAEVcO9q1GseWvtWw5dX52KjLzsiyR1uAPNVs+2zH+TKBdeTpDFK6bQBl
RQWZGP6iuPHChETpWVQxA7H2zEcsZmXrOMRhHD8kW6XtFYQ+5klTYQOPaGuDKDax6GzlT7fT95wi
h+GTIHVnsyTOv6uAfIcH/buuXhAZxk2hV7VFCQ0/fo+JtQs9xtALbiP+t91eOGruRYz6plyevniF
UBeRmnH1mADy0ePzECg1EXuRzDJIQFmsn4nvwrHUcf7tJZ4GI8CNxFGXKK0sSw8Icdkl8AuWEvIV
hNCpvzVX5CY0L9iBz5WWBumWvhejYqbb/pUHZ6QJ8bLdTAYq6PPhgUh0U28b0S4RZh+20opdxU8U
DDhyQDJ5PhQ8zQcwTCJiblNodRgInaMEC1U8QG+e7t67CZbcIYJKdagWahoHV4kSlhx8jd0oEuy4
65uyX4IZaTDf0vMw8E8DEHka4RLH7BaoHyN+qK098aatU8lOx9bqtmhhYHb0DSaD82t9jQPJUggP
g7YD5Ao/8l7/72N9vG9akiMmFVGrnUFwlo2X7MI9gdL/LVJfBsN2W7dyoxFZ2U4KTPR1v00FZCRU
Zcn7iKj7hW5SZt/sZxvhiQr/E9JfJUm1LeC0NX7MTQ1Bg/8sfB7eQUFU61l8+XKI1mMSuoZ8oxTr
ng0TZZkMpz5x1m4vWRu+H3YUl+v6kYY/fGSc5mG97V69qUQvKuAG1sxI3xkJHmlPhWe5r/9/S86w
fFmJTxnAm163BRVsSuUWNpRo30kyh5EkvAsflLHfvNwG1peVQQF+5UJTQmsCM6CZ+fiN5MdwEPty
TN6lzhTqg6yz93qDZJAlpeyUmJCg8IMLuXlXaepX14D1DODbXoEFi7+Nk1KVgAhmd+H6e9pHqdIA
m0+E8OdFRleEZfpWu2qoVh/v4GuGllkhRvUZflOajR9R4WGJ588teHHO4dd8Y3kKlCQKEYs7K6K2
3xNIYkada3fPMFKdg5BBGoW6ivOaNe3K34CuNvF/L2wHtnZRqaLOuNyIMbhO9864wW1oxhUflTUv
iA97pxweXpcuysLi/7HB37xZHU/eO1qZwabgWLz8B/14Yubun+M5z1H83cHcPQNQ5ZctPQqutprb
5cUF/2+6IB5mtRIAydxZQObkbZamUzbfUqsnlh0iNe3wmqbDlrdcZ65fRzTLiwlgXeYwEkTHdJT0
DhF+eLtFeeJZFGb0R1j8qHe1myRRfLPdavA4DlWkZh84vn9QHka1dYC798cPpYOMwWUj1itKnMK0
8lOsVbebDEx8O/2SfTHAvlngYd+NZjS0I3QmrdQkxy6dH1OsKHYXklUDm1NP3QC5vveJexGDpoZ4
vlOFwYy0zzR/pTOxbXcXf8InZyTbVpCOgaYx+AYzoAx7DTX+43iRBmWQgghFpD4FG+jmfkqr1PhV
r85ejBDse5PhqeR9k68Tn8tE+58xJCskdW8cnDtX4zZ12tVN82RwG76dAiQczOsolf52GalNnO6/
Kt9a0tCUyoJhLRgUxuYVhhXHz2G1u1O/Of0tO/zRw5KUkm6Pu2+w4bi8md95smOKiUp/N4lyK6Wm
NffKz4/kpzdNbcDNKCi7y3fux/gQAG0N5y2NL7xQ7d4uRghRJI8CkpYOS07+qSfgNQvongw81++M
dbEUDG1SAf8kjRUv0Xhvr+4+OybLWn0frX955JrHr6N89Gl6wtilbBd6oxOEWRH0jkU4Nn7nwPaD
4NLldRQO5ZY+42A4BLjX972sZ6N5eo66xjEDPSSHmp7bs4dS2sQhZuxf5k2eHZYKTc1DZwey2//C
5gkzfT88YB6Kr2Nsss7AQL15qJI3Pj21Sq2So4awpL4V5SDD8+zLqKkuyLe5deu4IjQCGR76q07s
KDxLqGunbMaFVLUJIjJQ1emLKL+0vtPOrhdGDURzYNX1ONt58nCqtA5hmb7ENwL4NFr/xdlKcNoV
87/WEC3qRhWpfGk/peMUv/V4Uzs6YwrtKWX4+vF/NKlasy/sy1M+UuLYZLyfDFuilx2CmquH5KbP
YxbBsbSHuj9wkf7npc6UVgZwEXayWnxsXEqNi5GEkuypI4zWYjVoD5awc2kU7uYroB13S1Z7dY52
fvNRnON9Emam2zuSWZ/dVLnEj/4D01HdGZ7JQLSResaVFhVO/jlcmxmwMHAUa0ZONDp+KiQA/ZxK
j+Jgms8AgMMvWC8NZ6IO2zDlQkV5QdUQJBpxIN2CXdtLg7LMP8NiaMM8yk6EKNpAJ9CJ56U+Hij4
8x+oz4ffl1sp+C/cgkcoU0gq6givyH65Ubnc3ifYK8KDEY75djZYcHimfmCTeHpMm4ltL4S1F/5W
McSJyxMrIdIEWIbQVWQW/SzzTxgz5TlqNcKyog1GJh4gZ+eWcQyWp8ugzc9yNXDiSUkLJY63e5r2
fDVQ68Ne8zf5b2edopCAH9rys+Y1MkNGHx0Xi3nbLUvUj7VzbqVc6EtSr23E8/g1KzFlUX9mh/7T
Otiqx8QbwqaNqxuenBE3r+HdHfTBXFa/BmlXUf22dWZJUBQxpA0mltMgkozwxTVZHMKhWWUKAwFe
dJHRjVJHkv1ms7vhDglrjYY3kJbHLncg2H+peCwE32UdGJuyIgLHZVJHlLrSEdfuDlI1t91JEzsS
XnxqJIlMH7urPrhXsxaaVrLUxxHLusmPclNYkC7iQFlqlBx9CzQWkiAzuFGUSCV+5/Udwq9yCFKr
HRWvdWjlW+yG6aF5OjsGd4Ykt/pxtJXOQA08tOIm3CkuJD4sw6P7vyLoJoCHB4Gk81MhTn1n0+UK
GWRMezJNH01pQAfFLIhLsGlQdBeUpE1R47y0nK93d0+f3IvhLSk6zc7QOTwfpMVS4guo9Wf5BnSS
S0mV4O9Y4olB8DnweLGhvpvb0uCbtgBBWY55SglUZcbWXErSDbWYlZouE1dK8aRtEauzDqEMWetT
XftUYZRl+0TXGA1oo+NmjigxXg0r8pdPpwt19jjcTRWn0b3cGrk1uNc9rWeQtZ6/HAQl7m+13HaJ
H69dbtY48LxZsD/BHf+djiOI6J1g5pGM/ztlmt6EpC8NgqF4RjYnIOMJEZRpvBTfu/HrwzK8iYuy
P6faGjE4kQGObAHomZDd9PUAtrCCFaoGpqXQvoJV9vDAH6WwcHZBj/aUtZ4dKQIYlmYfCtPo6A44
kWHzkSA0cQFtNdNlk4ZipAKmBN83vhTAtKGDTvJtQ8CVeCElcYZzhHfFNdzB991er4bRvFo5uEV8
U2sN6UWrzN88rI5zPkz4PPHSZ7/couT1uQg1h6bWR0cRV0c/TlNZWilRoGPwdGlOVMV0oBsuwPpU
NH++IdPUoLBXfAssPSdzcrpyo6lLuJQzT2wT0Wlx8QK4ZADr/BbRgvgmh9MZFq/tFvolDPVJTmcl
GCFHnQZjFPHz14iJGVOgSTbfYBBdLMRafi8oKeCQyhWIvBuwYLEhjzV+jejzfO0PhgIuLFbcYBjz
1/rR4YqNlv5nE/TdhFX6ZcoESwi2nI3QXobGTdND0gGfkWb3js8Dg0ckdBEwfRufFXmOzxdIjm74
qc6aWrUobRX4gXpFeasQTbsctviSXwoT/Yhtw3twFlxwWgubctfIJNvy8KVP2I8JApKFYCUSqcJt
VuDunJFnHdQeZnlndVJE6fsut8vUBXxOgwWagVy1qSXHln6oeqgN0BPZngj9NOgdoZnJcJ2Ooi2R
V6KCpWM9JFD4A56YVEI5sLHuEd9OnQDigH0lLoTlrsX9z+ep8V/HOTASuk+hevpt29tgB5Fr5h6H
TDJfLfMhcsf5IXlfRjwL6FajSstZkIFUrQOJ3+Plc4oVDda3IHiWiyGeaDcXwPaa9nAPWJ4okN1D
CmSL4uji9Mgbn65Q3kEC0TVUajzJjoBDCOrGSunADazQ2diSIGZ90FDXURFpxYlYdA+Ia2LIzo2W
MP4ACkb85R4lGTHyTD3gOAPVPZKhMn7APahGWsABqTnqzWXW4LgDADlSuavEMeaSkSV18jr++xHG
kEXFEJo7wcciUW3acOxovtXY+Jvca4G3XEr2CGQP+L5oN5+XTpf0IOAiCnxpuNLqR1ZV21exnXiI
yOTC7HT4jxdOCB3VPvgCEmlSPN6lPLFSBoRbIpL7VY/bT1wCSgeucMV96oh6zLU5VJvq2QHbxKQA
jrRAahU44t41MVHEZE1010Ar2zin8kyEjcXYTBdZsYT1zOq6Fi0I5qM8D533JknQUsH4RzwpYdjm
Utuuzy+vFKFvz8RFPwFZMFWBd1mbdsgFTcGpstvurJXTrVe3y/AVziR93FegEb8r7lnYYLDAC719
4KWg5ck7kPC5Jzj5UYtjc7Eq53PubLZTZW7nycvLxVGQX8938ZEd4Y9I/wd3dtm+6vRKtiAWaxA3
hk248zrJj04DvLY3xhdWOnS/AAnnuy55gez12uJcTsB9n6jukENMAwu4xYGkt9JvcYKfJqzVAKBr
M/5EnMAER3JKHo48G11MjmoLD0oj5f5UWjmvd85+VU9y5EOLU76zJBQgmredfQGXG4az3RwuwITV
mr+oOre9p4lf2/e8aQEn+3B9inPgNv+cdL9tBWI9wjnrTnz02L9UsCPrnwlFbVVknrUCTvUeiZgE
g1wetlac2AOEcsLtV7nuLWvge3HNf4pLBc3L5D760GDPMKAoCifeenvtkcVEPejTtzCuqE/Axi52
8omB7J+rmtrKzOHZpkqX5Xn2r6afRgzkShDzH5mYHodktdRpUnoHbYhqs1VFJHts39nk2gbGsnvS
7Vfbtvk2oQs2vYSpRVeDVhk8ocp48Qz5DVfDAJl5vMBbZYuSKcy9xdTLRdiAxRWOW4RX9NYuuARO
+wkEdBYCeT6Mv8F+HdoR564dVS/q8AWDx4ENgdt7BjceWrARvhp9MWSyCqvGToAkysxgVrwP0eMM
bmDAJ6IfnT3qh0ybZpvORFgtCn69bKNIefWgTxkXNQqLcwPO/Qg8okfk52T+oo2aG5fjr2+86bot
QPT4M52siICYdZ6KpVhyrxirCVbSU89f2FTnfJ4WSLAeNngjeBFVP6jf2V4gEIJiPaOfOnH3sCwm
C8EhPUjUJe7oI6gcGCEeZkm1xt/xdxx8UWOsZfxEKVAzJlHdrjm3iVu72CAdMcgKFD53t3DacbaR
mOa20U27VMU1RTUmP6aUgl5Wb0k++3afWo0BcGZpsc2aR6JAhbYnmrd8LQedBhJj4X7jJR3qbuyV
vw6fvk05MLwZ1iTEMfq+SH4bGwSiRz9z2kGJbTI9UGO+h8YzefAFXEqharDUJw1xeQ8cEUN4X3BH
v7Xf/R+OGlPG+PZhQMtFm6D4jca0Z+yMGs68FD+tf92JJmPf0Cdyq51Suovwsd/QZLLHjOh+6xlJ
hx4McFRM/sEaR8EHZMhiG0QufowxDPUTcVEep7tORkjBjLImI8KqtUxIfiu5wYGm3CFx7l50baNE
LbBxtiFcYMDJCvLEyRliwmpIt/OKqoZoPOGO4VArQ+we1RsLn6utbyXmGsEgsQQrvX/5UGXqNGFE
cY0XPfpUtFm5kbmNGcMUk//ZalXrbnyTdJmX1JdIzjjPgTe0OS0FUQuOK34g34mDg4Q2fcxV9JZE
Muevd1u4r/Z8wewuRfDum+oYRI/9gElWGNrTnkNU9p9TANEEGBA/DDGfk93BqD9RONsB3ISWAPg7
xAL5OwAqcskx25ZpX2xJTu34xbHZG55x1h+6njnVqEV+dphz0ZEN+Y3T6OOFLnISgjXwwUtKb+SS
EmFx5dO1tD45cUQIfP0pz1Sm9m7zvmyXoIFFHFiqweTnzLNZZR2lMjYSrGdtpR6j2YRppBU2D/o2
PT0+oJDBilnUC0RhWPO3OMPh1sSnNvtiZIGTg9pznkJErFlRysvqu5cNT6R00oSTKq9SHgY2mtY7
IuZ+aRb4yt4oTUJY2f78Se7wT5FKNCTQlESnJJsEItMPSSPAjxMSA+oPJ6XI7VWE7bVWjtcd9veu
k7LwP4VK6xTD+4H6PmkUPwFANpsO/yRl2E/UVxtqU9mUbekcoual9XLFxnbIiYN9OQlora5ncZNo
GDGLJcsa3Y9Vvi3GnlWewchh9Y8YeYoNSMPHfKsAuAXd9ZCGSGv1PcpXwTuHpngQvJVIYZfctlWx
AHRvVOlRcSdgPke29djMqldudgXwB7cZVxS/ckP7eNaEDlb2mTCaGoYZGfwlIZ1P1WaQ3t7lRFaA
EHHGM0cP4u+OCCJcaAL0aC0Drk+eLKHYxqvD7smg/8k/bupbRtTz6xXm9sBWS9e5aAWvsbzAtmwK
O6kRS4gc3rNKgYn9YuYiJyAo2FjHx0p9WeoQci0LIHBOpzoRBK6GfYH6frhAxM/IOnqsb6PO3EBV
/xYhTSENlCZ2BCqcbj5awslzgmpF6mFkws5Wcji02cGvMk3/NY7IUzrf97iWLmFhMu5Fx1kCpmRo
as1bfnX/5UWb5BdDHgQLE/vVnqWnvM1X0TMtVoAcWSTVeYHqPHaxwvQeZ6xTD6qqjDPvexHv3a/W
YOnf/8trOkaqmOXLYKKmw5/dxdGWZF6ZJyi+XaSOyVzlX5UeIuAn45dI5GMgopbeDjHxsOfkWnzY
sHYaN+c41mAbIvKUIN/mv75cunNPnSziEirZKtlvSgnVY6zbUcc32EQyBzokg2012WE1lNCzl9E8
C9ZvG7UOahQpO+rqkL1J0bBnoNhPpWbmRz9SRAj9ZdUxSKiXO5N2o9t4h5R8ewZs+LMNUwfutzG3
q3+P8rbPCQ2ZPohi+h6gS4SRafSqhaqg799OBPUkjt7+9vNcNvz/eG+9R2hBEIyeaz9xQPmXJIUd
TVcTlkn8xZpY5vzF4q4ES+ANxMiQt9XX3yFzvp7DKcrl3SfoDaqNiQik+K5z8eTX4DSx9tV+yP10
nfm9IBXoPKxAzA2xaKSdAnuyFWcO+jakyiUMKp5NFO77ktNCCJW4jodl7ZqbbFrvHxdpgcUzTnDJ
CrEBMOQtBdL769CAVhRnhD9jBSe1x40tWi69VClmPK5I3Ek+OivfwYGfZZipUFJncc1D24zH+4xI
LfXls4I28IwOPKeuDCxUqD+3Mth4CuVd3gMvTi+aS6znnLHw+i6ZaV6S0mF4rkQ6rdCQ2nJN6UOv
774j4VSLGh6q+HhkfudIAikIaum1bnozFDF4tBUhVJp5P2eFiOJhjygBPXQAmFxxbqHo7i04Pf4f
/YIheyPdQcP6siuBhozxdMidbXla+qjkcN7DkqLJ3I4T0+wi8ebn1jTIExQ/HeT6+rCJIZNHyi5L
ggeBEvya4J6kvo9jj/j7fqxjq65WJIe2UI9xu+y7h/eXTWqickuWTLyMf2av8bf7y2xuAlCD7UZQ
dhTYsB3heeNy5SEZ6mM6MIxAEETciNqQO8SpRAkOHYXkNNaZ8YjAIXmnRrC+s3upJP6/+YCRTdIY
eeuG2d/2q9Giv0qjOs44oGCIarewRMRF2xuCGxQ2Neqo2GzT9SUpyKCltwP4wzbKjWpWzJ7OE539
tgjSjX7FK9SFCTRGIYGEP8fjLVOOIkknRc6fBc5yDVvW5uYnVeyOBa6LAq5JCmG62RdxKk5VBwGD
2oWNU6z5MDuXGh7Ige7zObrVrG9iq4iL40MCl1fCq/k033BzlBldiv2nxgbdCi/3Z0c4HBGz/36d
yK77esqbeMHVsT/0uHGi2/yzYPsTQ0UR0QYdqVJCXZDfdyqTcZ13uUZ/mu72ZzAzDpI2rZQ6nX/5
9U3gVKRLXYkJYModafhuhGFiy4Ozgwc6XjCL0iSkuMoYpwx/SVEyD1PB6s13R3jkZvFnJwWBDWNZ
7q+Mpvh62G9KUkTl9v7MJqS26c/QrMIzVppy7RTdFmN74icLbAhUj8Uz9VL9OnUwM0ZUbV77VaYU
t6OdeAM5j1RgXD0pMC3ekdBsx+yN5fCkK7b9wV9DUtouGC/NKBavAa9JnWmoiVGr9wfyGLG2TMlX
ez336Rzs4acxEYIiAbi2ofB3OVMnbKMZmjm6IlyPvkvi2XTpQdoGdiNIB7LqAemTtRD2kvqFXbR+
WcsfoBzcLZmaNC5n61i1qeudpz0EzmYeFQU5PDbxKeQ9NVDHzp6IgeJ2QAcV7Z26HKPpnbft/yko
3wn9ZsQpul5hTaat+S39ufAxzJZgY/4p6cIaIrGPd9t6uLy8qjDpMPif867M55jppYRZLj6a+lTA
GshPSdo9ZEb25U6fHvY5C62WfG10UmMkipj2N0dJ/CA0n6CEf5kCj6DkbkMwyOcNrP4NuSmISyDC
zBP8y/oi3V2LOhNoIx1kW2+AKfgtEaYc0hw2k65SkrOjVmGS5jy783mirhC5w/bH+KDNYnYx27C6
pCFKZnQwzivKmxyQuWyyAZfY6/J2P9UoYeq6cQ0QHpiJkTODnmk0cWvyx5vFfv1riutDLYjEtW5f
0KyTjq0uzJx7/eEOV7NzJcgV3S10nQCc55KzGRcMv8xwzUXvpeI0VbLfaMr6OQfcUYzjLyddC+d8
/QlDZfUm9ath4wvPwRQzlnSrBmWmp6VpbwLHsrjL+ErQqATS2PoPrPbxIdXhAnRDtSUOklCFT0FX
cVOUQUSga1QmQWXGo3f9VNUTusTrTWZoQBATsck4vqoYpZrwxfRcTQ3QI+1UMnISmLGh/7JldkQ8
bWaYcqk9tO6UKGLnfcLAh//a0PWAnlksdw8v7Z23gsq0258gHbhstQZQ8YX8Fz9dXmn3nPr9j+Er
5AEx+e75848hxbSkPyH6uBJ2o6tL5PVTPslarX4lylEZwbG/3ZwQN4Z29f6zphx8id2sD0BWhPTQ
qv/YP74NKem+U10b9TIDAcT9TqPaaa/sw+uj1jdcdtqMZztUihhiGjs2LvFE8nxQQ2MSwhV+pwAi
zxTwjGAvGrn6aRJYLS2lkWpG1dUkgU0AQIHChxLc5MM373pxDKd/1YQ4wzVEiTu/w0pqvIKw3hnO
iv2uGjYbUHQfoTgbl7wkJTZje8S8PWNgMvEDGQNYaHJJuRYI7lbDn1hcpGRN8KQO6pnjNDLyCPp3
F4e3AoIaRL/Jv+nBTgu5JDlByvCd620eLTqtvkHzfWBKTgLjk255BLmR7wEuzjGCAhIqbOuv8ZCB
JkKbdz5LYHCn6k5NLDzmAJ2ik6qg6YbyaoT7YajTcJzpOqQjudb6VTDqNB0EDfDZCVpDLfwyaQpo
NiJK4I2DIOKjrURfx0WF6zh743qSqbA58VHltt+U33r/WIv4dXHx8V4+km/nhKZmqmJ2oo9pAeUx
LNAMiKRtvkVsjhZ7gWVKq9OyWivAVgYMYT3ioljocM277KYFyR01ItwBQ3qFeXWoh0cioEvIwEOQ
LOMr9uqHhbKEB/oDLsNOP9RzTPFla6ZiKKRyq33DTJYBLLA2G4tcserZbtk2CT6qkndSb9IcFro2
hrP9J0yvFpqru2xYHYVire8CiQrv20Z3Qc24T3QMet0BpxSS3WSux2W2JSkU5GgME71haA44r0g/
3lnFF97lk98tGe4M8y0XZTsqwwjBPvyIE4UveielgoJYbOwHcPNglAV3giQMjBG4CT3ThwAWX6dJ
cxEZkgWQufQPlIQP5m95121gYWxO162oVLAZzUbq1TZkQ4CSKONp1hxCHhptR2p5s7oV3v8p7TEO
LzFEn+XZVD0sxlcERbBjJ6f6GscdOEPalDV+VBlgnV8kGe92iYTsxpwymUfFGv0nqWR4OINXrmWZ
erOe+e+1UPDZn954tI5h2HjOEESz590dQ+y7mnhOLWLmLbU8bVymJaU28coaEEJIvcOuzN+VPkTq
ujmu6nkut8XyUyPlov9/Mr79oB3wJMKuY4MjPgG79clcg3Vr8nHZezfXXPtQ9nWEjz2u2RYyXSgc
AbkkQyDPC3RPoDVVYjMnpgQD5/ejKGAouwC3L8mjOTTaJBMsohvYXHz/MThKdpZoSXsQhcvsCQZ3
kCKA6GyHbr804DcwUsiQLtpiO33pPoMvVUf/CBXGAK3J6UhvQbuC9YI33fWPNfwkRpDqILXzWRRH
oeifLvz8DbrP/QuxC4oYpX1kE2kHQmyMNLoixofpsu4ItK6i2b8jTLsYa9ZTNxXMqjXNaiksbkmt
zgR9bzpIHbKien/UK50oURyiWDdJpUBtV0E+Nu5/LK1rhfTW+nXKX3tulfeMXi+WNZQuPQ70w/zK
QUOdA5S3TGkinFuvbzXjfDyhPnxd6eJSe11kVmKhXCu2XjsWM9Qkz9sjZIqcfcdwqepxjxBgymUd
01GVy02UDH+HBIaRnc4DJMmVejMicrXkwBp/0JTNHwxaDoR8ZOdxb+bh7F9erkAjIQlfZnu4GUn+
RAhGGSyheMfk0iucHMW3u8yt3Djb0B+4tdrmdOAp2JD2BTSFN0zWnOEP3NAQnWN8o5A9p9av7wVb
Ua8kljgInQ9Y2fkkSg7V7tbA4RHH0GzcJ9YTwFNmtZ4e0sK8ddpQIbeqmKS4Y7fQnRBckSX8J5Gj
AZPwlmP9jycokm41WknNQrxzQBKc3bn4SzXqmOLu2P1L+oEeb5vqeyuMqm/86bh29fXRriSI+EVn
0EK3GpQvhyDMvv8EG42jHfdB8w8r0xzYAxMWklsfDf1voAAnyRIz0dEt7saC3SzrI5JwlBdJgkDr
3OOsKEiBSF5D8CXvw6ptlSBGilmYpjhGxiDVuviqvY/b7rZy7i4/2nun7OQKLtJA0QvibH6+7/3E
mvAUNgggimabCQ4vZlETGi8BrXom+Fi/cUDDMc8ShZkLIFf0ND6Fm9+F9/lvRn4srfv47VveKoqo
mjAHQ2nDsslOi5r0oQfek92fZB0DwKAyP/lJtoMoPzy26igivo4V9GojjNE8T/B0RB0ctHxz53gw
g8RpHLUOaCbLSHP9djEN9RFRVc1eMF/8gk+Vt69F9NuNG59HBlvnyBCMN4++qGuY3UFYkmTB11g/
VFBrDRW1JOZMzkSXzLt43rZRBC5WZHzIXN7e3/x4QzP0HEhLVnz3Lzq+/T6H5Az8cEx3Y4zWx6yz
s/A+UgVfWWxLyAub6wDLCqQVThDfvtKThH/KvP9HWU1W4+wCdHar13PGrWeIKU+393bwmUfjFVjR
WOVCiGyo6MpVZwTHo3ssCeym/4wdqbDebd4jT4dA5ieI69XMF9VbZkYeLYnvjYLmsmVIUgi2zFsM
9LOhL8MJZ4rVpaiBujqQICCWljhwS8oNFPmeyJeCKsCLXPbjaYGEN/wUKvMZMTuVbq5H803R3af0
861tflskT10RvQYdPa0ynQIDfogXHdnWVHhd0clEj7DwHmjRX5XD5X5x90GVg061iNc8JH9hmrvg
MKIhZQjLjkPkDx9OPnA2DKhdP3c8Da5Jhlz4DfhlnUdRk0QZcu9DbwFsa+AXKQ7HOBqfaqfT3Wmj
XlVhDnh3bePi4RCfSxuvAphjnPwZWrM96v3G1Dn6nAQXrpE5F5gaKJKsle/M46XiQ27AwGE+zcBx
b1llcEIHEU+D2GQbY10HvP3jvg4bwlquPVfLF2irDoC8+AKnh4ThFD/CiW3yjb3OQKiSrCMR7KCu
QypPOr6MsPDt0e+OEVpf/+1Vjt8aijqJmuTV5iU+YrXdIB8DPhscmNhSpb9zfllqPvzTBdPMc+/5
1K1Hl32qNueODhNvSK9iSjx/wdLuKB0BijQtqzafzCD/8wMTq7KWFMDWsMtifNJSCYYf1DNeK4gI
RJdxDLr8AB7lfxqmyoGZA/bSX/uUlAt2ECuq/mKtRMZLB1WAhOEd/Ai4e7QjSyq8XaNyzscBShkK
Pl3hm06BOuZelq/ptNEezauVpNzMKIN7oRFxFA3zLt2E0a1YgXlZxDl9gg7NOUiQFKPZwvXE0sP5
Ab9ZriZVS1m8V7cil2amAsotInvHhNUNDZiaI2r4DlcTfcw8zKKBVhDJ+AmhWJc1w1uES797xM6k
cbmdVhDecqOu+/eYWKvO1lU2aAAnyZBZsw/7dxRHTt9yokEgd7B52PV29x+xkIYp1Sc5VE3UYLso
dDCkqrW5VBHYY1uE0TfBS9ck0xxV7FXfWST2CpWTKTKbxwy451v8aHf3RcXIJb2wG2rIuUobpLFn
EWd92P8XV5GnPEAFaBIIJQq+tIdbpKuRDmXlrA8rmHAGhN1I/cPz2ejphakDk0kM+h88VqopcHv9
Pl0EBPM8gG1CHai4lIJb3gw0+m0AV6z03qXVVo+WjWCOb57H9fNqzP+d9eSCUsIS6NpmWgFCgG04
cpUell3cQhjIIIt3Ym3Q82Yq9SxpIZW0OZcb5jjrr7H103nKjM2FjK/rdXEP/gpccnB8SnAzyhZo
0GS4SAG9mCRTd9ZwH26q47c3zkOeVJqwA389cbLzRqaxNd+v6QK18+Ifwd6GAVk2EFx9iwWCLuKS
pJ87OewWcanRCS56dotJ9Jh18OTCyqnIkSaIubPZEyfSOlqbT8LiFgGQdFm1ekNUsfMpZmnvxCfm
bV9DQNn5O/6fHkZyb/JRYnOu7cKfWuisVa2HZUxZTvTUkFvLmZ88ujgqvCgTm+hF123OJ2EDbciJ
FrikaLvuOVhQ+ynwtC8mimOcnfpfMr2sJsdHxVKdiqEJN2RlQZWKQg5x+JAWIQw4aNmAIVGWbTZR
RL+6Wy1r3AGTxr2166zh8YEyGaw6N4yC3JK52muDIR7Na6gzSw3tOSkfudxXsI094f0EznTHDpST
TcFJuBeasiumpdlLwu4caugpkmYIfzCceGrvJXce/02NXaQtyFY4Wcp0KqmdAlIHEae8crOi2kbp
u48cN3he+SThldcccGwlgMp5XhGwudrE3SNTAcp3E++K/Rekwwx2ShfYJr2LOeu7bJsW8K0JsK7b
gXJ5wQw9khlWj7oMT6yfn0I2TSLCkL9qSnXwwjFgytSCCruGZ1B4T9KP9OgySXb1RSrFhorQtCN/
/jK30g0eOM31jrcVsWcwtgujWpiFqoPayZ8TuMgzJ+bfLCF1WWE2ox9G5wCUPIhHjCSYR8utsXpa
YgFDhLEX8/79VS5zND4rl57rWuuQlXKdEjkfp6iVskP+Qm/70pwLc/8YSooLFQcrfwEJYhnTq6eQ
2aodu+wpS0T99wUdG7n6vv0+IHTSxFODwzILiA8gSP/V9IhU+sYDeegYVn27Culof6ys0IHg8l7N
lIn6YM4yvkBUXRBkZ0ovF6Rjn9mhON0q96WAI8f4ABBOpMT7FXjUSVGqDPOrTzkdp5ymJ3ROirDY
U27kt4T1JgCmSojvA1Vs9hM6vOzhbqazs7zyU3DUyubSG7o/NQZsiijEa0lsNjysDnjg0g9Q8az1
7zMYW/OisRLdk8yIspcEyn1pqDbOU9qtzM04ryCIkKuj/Sm1lkTikCTIqwoI//2outfZovbmFpwY
9XpXQ/NRTavXoRxH9X72VZw+jZbUUAR4WfbpyitIaCa5SsaEDmJPKWtScXgBnB4LViDpZNiO96UJ
DwqxyZujj/KT8Sz9jdbc+6rUzEMlgbxpNjKyaDZaWUCa7C6NB89YXMLANNVjPxUr6a+eZZ+jeCGk
KVGLgbZQecbql9XglgONhMWH8gwrznO2VGIP4lJPHcBlxS0CDBgPtisnmSq7bt+KV60JbrSeg2ag
q8iBsWQ1fHg245SMoHE89zdESE0RUiuq0oCNM+y7B3QIzTlRQFdO21lV7YavPeHRuIEk06hRDNz/
aUibmL/cgIwvllX+vYn6dPoYwfDxyjMCm/0ICEdZVjjqhFjTdzNaVyE4gqttzZ8pfT8wBlSyr0cg
9qdEq4QGEdZsRXBR0/ZYjrZ9tHXpxz9vY0fGxtPhhdaKApfqVRJHq2aWVNY+GbnhIMz5EwyY3Iaz
qAnSckG6FTdYXZncaHRV01JdWlGz9kIWs9fOjFx+VwOn+jk/3xadqUAW/ZWY4/zkXe3CMYJkxRPR
ufgfCCHx6C3xUDg5Pz2nyX6wycXhOAeik9sFjFz5ny22y5GTLo7lWQtUt6kMPPTpaDxlD1asQmjl
6Jprba3U2QLHnIeNBpRvaiEYw0Mv8843IwKmaLG5xbRGCsLetjAcmui5YuHAawNZhxhDQUYwpnEQ
yJzMN0enakRhmdYvlJjZ1LBtpw2alDatWNDQv5hr1zuoL3pVwr9w8N8skFSK/kcP3BW/182zYDs7
F8Sw6T+n2+HdWGn6Qigvg842IUE4reipCjo9GwaWq0tMaGJrF6SNusY4D0MKSHaJDumcxNoL68Bh
eiv6tKbQtmEVEMuG+TDj8zZSLptEFWzmeXcnf7ceFC1RGNDCiuFBZvs5TI0sqUbG01oG334YZTXY
KhSeb7EOGQQzmXV2HQqnjPjgCxusCCesg0SBhvS67KDcXUvkKer7gERNt5VgtWtcPyHFF6VcaWnN
lfn7q+PDE6SCQc7oOP0YYeNg3BwOUJVK9H93OMPLBFZKZeL0/dVSFByOWYZR0qXsjMie8B22J15U
a+LR9WONIptI5PCIxeMtQC/+T1uHU6aNcU0k6kAVIgWccoiDPvhGL2xP0KehWn7Y1HSJxQKWyvmx
OkCMwfjYsKTOCgmun1cHxzvf4rGRNg6CG0kN8GcR8PpanmnUCUklR7kYiOeqgCXFWs+x4T/ceAmT
DJFdhDl0B4PHff8pTV0oii9wtyWC3/0PQktxbMxU7wJhSttMXFQ3xv/qCENQ/vQIipbFGeQtByAx
i5tMmYDcsB6LuAubuNg1fSRnvYukN125jz9G5ZGCkYtmh/O++HvSS7LaEAHUd2vY7JuJTt81jQrx
yAV4xhrRGmYw8nb2ksdCuAciRVOm3QhRf2IPaU1OOAc/W1F3TW4BcHiahrRwNXMadHrNiP0KmYSl
SwC8EaiAcD7ZLEl0UZPdHJtAqwlvkRRH0r1Za8gQUCC7xBzArhycYHMlZzYqa6v8fg8yERAZCKDx
3xM4MvO1Q2aWln/2ipOTuDgYFREsE43x+SepGahQQTLqBulKLASNMnHGuWf9Z4EK5VLKNoRBfgjf
kISuADEb8ihg2BlAim4qtKErljvcrIZnOcxxlSrkkdg6yEZMgl46Hkd2kXOxj9riOZVQQGIkXmqA
UHPEngY9Nw+Vo+TRJnwoP7kSmCo0/gKmoiIgQYZ5Qrleao6ZOHu9QMm4G7nn16ZmUUdDVbAfAZLQ
506CvNS2ACicW+1FBKeduLmgfIazxmWN4nSrBXkNf3I4Wg76WK1ifm/xvyKt+44k8s48UiyLkkka
MVR+Cl0otXQEZqYcNYoeDCTV7j1Szp8vhGdbbeCvUlLLxhe4+eBKjKo/kRlyaG+jfFr0BpA2DX+0
7AExI+12owb1CbfDQ+4cCI8xHJR4Th6z6gc6xY7wRXrlet6h1wcDdKLlH3mFgMuVSuH+rbbo1zfY
C7SHCDAS8yRM1+YzPpOP5oBgJt2jzrP+TX42xponL+TmC7pdodoV91bJZenOAa1nG7V0FSeoTfiX
Ot+BGTZzeCBBvAhWBvEwYRsc6XUQ85wFdmufyiW8wt8chn2DQL0Z7QTWa6h3AHSaY5jGlGasZtXu
0/3F4X4BHjcC7SkBGFIfKvu6YDFr5Yo7llIIa2X0X4QE6bRVuGjtnkIL+3mbmVI0pPSF9GjsPbQJ
Ui0dEG6GstVsfCoxUzMBhds+zv3tkTlTRSXdEWT5HdhVMrwE1ZFF3gvd2iK4JmD5lGEJIJ5r0L/c
I3XKJXKOZTjBLQUdeDRk0PDfew66p4QOD+37sk7Yo4qJkUXV/kPpMM6en7kd5jaMROjF/aiYGGZU
UE3eAJ3+0tTaWZfFEI1S7c2g5mZ4yWDUkH7cbjuUMS+7T91W1YoMhCjashQXz17JcnXd3sMZmB+Z
su5hL7UxpGXHCBG8T18u2fjz/AsW+MTsoi+lRmjrOgp//hhPS2oGvm3b/HThOsKUbZscarugNDvB
T6vN+ME5RQuQZ8xU9CZQsicQ+Hl4CV5UMu+iTaWoTlPoUY35ityG4DTTPu47TQ23g7K7osBwUitU
PJnEFKptPOSdrAFLhYap/OyPs2D9/9nMMCeaLoiM/ZmW5s+UehUiZgfmEellJbuOXkm5TgS3xlth
qqAU57cIWYj8hzPFm0RFmBI+r8QWY1uDKFVCCxEllVyVfJ1G1k4RjBEs8lgLuV6uHX3NUS9ApXjf
mkxCCXIRON3i1bU5U3YewZULP0r9OWNNJdzKP7HNFbP9SEjJBekGTj4lSNhNlBjkHS9CUtC4Fkzl
4aMa6I9PsOAlIcJfxCH/3jRmXyFl40g3heQFoDfhh8pXVvXe6sNj0tkUnEZId8jcMsH3+tXR16/Z
U8NsfVfNLwMQUiadzeEDPBf8c6hbw6GwPCmB1nrmkv2FnV0kmTC8oHMLr7CmuVttZhAxT3lGutGH
Av4sCWPRW35c5my55hZ6zQvMOyIw3FvTlcSYjX2yiqXYX/Lh079/RFlroPIwi+eNV9jFc4h2/blG
zoQOkoDUUQUE2PynWXsrrs1pLVbcONHeb7cC4QdGlpQcuABSE6c/sQ9bJTue6ONVPlIawHUrj9En
vbyp+LsJYbGZh9cK80WMX9u62XhHyqR/g5ykOJU8nZLSN5EQOZKXAirXjUxLSIh1BCeOEE7IOZDW
Ml+2R18407yGnDvpB7PH+pymDFEoDBHe9p96/XSpUc1fR1ktLrSvGR1D3PS3EhJDC5KR5z7MHDf/
eKwvhrbPFqWCSOxgKGCosUh2lNs/xvm8KfdY0zl/GH2zOGHNG8609W7ZF8OffSORbaHHgWj9LyjF
T9BzqiOsA0j8Y90DHPUDwxO9M5HOalxhAmPlZWZ+01vwQQZoxn3UnTZvyESrHSb8xgR8xZpsdW8B
2aSx7OvQX7B9/X848RIgRVLrI3QURofxPyDz16LQrGp0DeSZW/m+rL8wQCTqVWeb3c7fMC4Vr+Tg
bbDrD+Vy7YR3gTOK4lNWo43RY3nfewbP/eI2coKLpoj37EJ56WzSbilBt/qUq9sOCjHGrh9u0XSX
tu30n1K1YmH9W8qvDpQl790ofpQb4PGZHD1UEVdILUwZ2scdoQf3wrwrODm573SgaLjn60dvW17X
/YXkG2w7YoHgyx2W91P6WXsv6/2Y0v+MMuyd3arhFDxwBAtcofQ10iMeM+wJJimSx9+z/k1UhRq+
VdoxQjTZjL/6UCwJTTlezJptpruHkgMhKfB+xMBp9P4NdJXD+2NyU+7hskmwg9A/3F0bYHSqphJl
4LKt24Mvi/lXHZkh+WhZMyA2rcjvRtA3fuVmyqd8Cn9383HlshEcCMAzgrEXEJ3a/voW1pmLvMAC
JUu5X5OuBmIfkpzFZzkRH2v3635tqP3Dp2yYKsN3NHMAG8J3ESkh22zvSLsIDn5VoJhyGOUhPv+c
XsFCXYctIEzW0Fl1hvtO2YwSYsYLS6bnCDfdklGaoS3BJzqzxqhGke1XtgtfhDYw5qyguDS930c1
+x2FiwvgsrNC3zSF8oOC1oiGA5iMHJapNdesSzwkHMe7E4+dVGwEBP6fZIvIutpw6veYOrfpPSXX
FS1g3X9Fe+yEeTTrYtsY/uWMJK/6rQpnxg7DT7xafIjFmFMrX2f7caxsehe/j/jPT6efXLK9jj2+
ameMjyl70muWcibdGMFgs27f74GkKpL+DMfmUviPk4Rym8VaDiTTocndo+rIxo1OwLR0GTwlqlHB
70GpmEQdARZL3lUfK7IDk8+z/6iCGlcqmVhksf4udCwAiPLwAHBo/d1h4ZxW4rK6B4B5vsFVfldh
vmNlCU7bPbCIEUuhbU9rWh1Takq3cDCAcdPBuM/oZwwx/KSfUBqq1kFVvZec7Klu0Mm49h2Ge6AM
+lYi8SDifpz/RVHLKXg3GWYT8Kp0nYyzUNCn+2R0qPJmLcxDphwXAFEqRQ+w5dC08sHh/AbiH+69
oebjdgo8kQgW+XeAlHpr8c4CxS8w2frJfVeLPANfsfSmvTTYNJ7fQpMtb5myzj+RyytkpqYLRXJu
9Tuzo5N5NKx2506YkMJauWB9S036glbWFMSqCgj9zplgJJ4ejOyXliYCIrYj09XnFktZFsNChueT
fNTE4ZKMiSjiWAHSD0he+Mw3x3iOytIvP18geh4Z4Y3wua5PLvZrz3QbsczezdSs7Arl+L5n9E3L
NUfJ93AXKXoTMRmA834dY/xfgsvWiiMhSdIXaYHV0hbNv9AxN+SeBXmDzEKVyJi2OBEz1tTIpBRw
NnP9FZpu+sboMpRE1rYeHTUx2xYa/nPOMl3vVaKaJYKVtkiyAUiFQW12XU87GUKQCf4n0mMSVT7u
5XC+/Af8ImQpyaFnbIzRX1gCeKPJdEjIqz17lJrUqN0H77W9Mt989iMtJ9HYMG0ye4EsrWkB0Mml
cfw1QGlqbx48gXuMPRghv8rPMAhZ03PULtZGnHGoUCnglYyZh8ufRAlL6VI/dlRa8n2rAeRNKbs3
JZPqsKa/oP+i+FgC784649KFySWnrgYF9qAufZOvhOvm5pTftD+wDOCIm00enU9vnDtBg6fxC7t4
iA410cLpOhPKcKuaV6xULjv2RKFkYpNQBvkOmnNnkvboYaGDceG/H2C1MQ5YOrmgdyo+0ntaVJM8
tOPxGf8RDO2hM/SYm7kOlm3L64dGRIUQJBN9fu6Nm3KF9CmyfihpKtuwVOFqztJAnxwnEAW9Ty4E
CBP112CFaKUEd4fxzpvungvJtwAJjQVF73F4b/jxYPr0daZu2Sf67vjDL7g1O7ETWvHNAdueuryM
WAAskQiuG99C7TlSI+T44VNsmmey6+eGbTBMI9WPXOnla+kdL9oymERWdisnB8OEyLpnaNB5JD/7
0YDya0RjZPTKsAwjzEUJPMVFjED45eeuLHlApiA+t3c1sjunAHnjyI2X/KqCM39QBEWwNIt9jOCL
QE2vaJDYpw8wLMe/cA8MxH2h+ETNC4i/tXSm9V40tmscIX1LwVUvbTnWgzm6IOJx+MgPNkDtP/Rk
buJVzrgiucoW+1sSncbK9vXIAm2LGgL8oTAVkYCAPawNs9/OKBxwvqR3AfZmPMkfussHLXfrmLkW
s2fCKHZ3WSEi9EwuUvlIfwxDW/6lmud7xTLsNar0QrZJVCwlB93W/+Y0YZx24ljfsAuZvPE0uTU7
6ivzqZLUnuHXTVR9Ac5dys7Toalrim5V4aKT77j6u7xJpINBbztRYFbSXxmK4DrHjogJ25eqie3D
tNkZfwqQRQDvXeIqjmpyLAhtt3rvNlzjPM7pUdCMI4ScVLIctsLTZZZSQ33SIQqr4jGO7jQgLc5n
7yCjLZcnU5FZ4qrPz72fpJkvF0bulAzthMOXC5iAilFHHALMEt6s/aRxHK3joJ3x83t8pmyuSC+5
29BVImFjRasfm3vZe5bZX5y1K6fy9LO3RDuCHdBxO+8a2/riF7VaVeTfGplhsi54z0bdBH9d+eYN
dWsm106qdYQg3sCl46aVR+cYQzppkcfi7tv3AktggsmPcKXw5MzFsUxOQwTcrPyRM9Sgk1mREEYF
GHXv57UZMIbVu/rpi4lGxpu2j+lDWDG3KLSzUyeySh23EMTbCogmJ1OYDGIPb8xrkH1Gxj3Eg0vl
sCzsdyqGaBS8at4XoZyHMiopspV8H2hX33CTG38q/GjN/+r1ceHURcdo2ij/5yvufS3IYQDy9x8X
GkcR7e48uYiagocamDl3jhdp2NdIK8UzFROmQfT6qnWw7HdNrNDoXA4JrxVB390My282lHQ912hM
NII6GxCYW8m3GEGn3rMevS9qNEL5BGE5DLabVL12iFRAwk4hANSYLSQB5zi55of2Z9LYY0lDEDOt
+iz8DKn9hwcBI2x1YD6ZOmwKyOdgz65EM9RTD2KgqfwqB3fq//5EBRQWtqgLpoL3/O+zPgqC17mG
Rw9e5n/x281oR60CoPOM5980YCPiDpDlwpURrEHCrFfbZBhUUb/Ziu69825sIDO/FrZ/a9ruzvoS
3+2zf5HId6uBzoIVJEhajOZpXbccVfVPgMCbrIG9I5coqOlDgHlJ0Ok64WLpepriTtVV+e8jdACs
vwOABrvPmK5Pidynf//Aaq31tNw1icXXI/2dlNCUcTkgzLDvlNGf04CL04/zopJOYXuXC/taR0n4
3peCIqM5GU8aYf6dC2dEdotUmHHUlNDqc/xt80WecELMOi5dVyDuxP6IPJJ/IoujjKTZo+NYVQjc
wLk4gU2BJ3A4WaNFXnJGxxBVkXMBzbNM7eKMlHVMmUJg0eSngNZmewxKfkLNK0GO3QxMhTwAnNEU
rcFtQWAXE7z2rYl4mRgWpa4N7QWtBCEyg4/O3vCpUgPWdseCeG1pTpb67+Au88Rh8ccsJYjBslXB
9gyNQ7kV0IxVUTZ9n/n/mGPfSsGEmPiYaO9oJtXH/EH/N4YJp93CfmEyZdpiuH4hDce9oMr0mfj+
o1nkKTTjY2/tX2JbHZX9s4Hpnh3oVVsk2O0MR0kCUxp8XKy4Ff77oMLizDXFhJ/UE4jwIE5c1EJV
y+CbFlTgKCx4tAzJsnOLBimO4NdffqOCniQc50zCj5hF232hrSG0+7BAnWE3qRvSAj/qm1dWFpC0
CDuFromERDMOhl8PfsKLS5B7M0g5wVT+zu6E3gNF2LRtYZtb9V2olE8qN0hVsnV08yKLo9a40UWF
Sl1H/h10D/BvUUfT1wNppbb7M/hOALcvT61ArC0vS5sMnBTB1ZxF4ZeZe8O3JeSVF1jyGfetCWcZ
QLVgZ3sh7v+jcUtJNqGrvTHC2ZGWs8CQH0ngywIbOgVgHVdnnVhPDZCDFzYZrjf0giQTRIZDSjzV
UMF/lk9DssMSqiV5rrOKsRs0tujdT1vBtZxYkMldQy0zUT+x/xfatlS7xnQjHegQT39RnclR3pXz
xx5KGPWbNyFbgtmfPGkYBBTOZ4As/j1GbMuetC11qWDRORTEoYNHZJLas+FNKcnYh2p4XPrvgurH
A+3qBiD+GCwwbto5GLXo/FYT2ZVI3zEAdhr+saxRScbPCHGbum6UM06gfdzZr6UY6g1BdNt1abXj
efVsav83FHy6WGsdkRSayiI8cC0Tqs4+wmJ/b08eWjB1xD4Ri2QsIR4QP3Wz/IS7AeXDGqAFW57/
3P5rPCTNT+haCBiGPHYsnmnbaOJVczQ3eBdeWCWnCh8LniBPOAJWTaK8RRH3xvxJf+0jFppQKIo9
iLvQlGLNfpK3/xxtTPmk/oMdfHzikTF5mzQLvrEkXGmJukhh6V5oqAnCsqNzuSiB0AO2NxZBuAXA
hcZBorUXxMA1M73ZT5x6MBT/65W++p7jbWVfURRIDNAhX/vCteHl3QQPTCJjWKS3Qv8y4qowlIrz
F2Qg1GwvkjQt0UkBgdpbbvkD9zGWdsm5oDCa8JmaedVztKTELPXOtxf4ojM+Co/MqctQxMpnBEuy
rVc6093HvsoPoxTCkJLYjlSw2P2q84LUmvXP8RrBSlD30Im+T4yLV5Vl7kZUBIJ7zLHtoQnSsWFO
LpTsQH+TVE97M0NKAYggUyiEDyM00YzUwlFrpmFkJYcXXaxc4H26NKjIkqDpTdAgx7+RXLpGokRs
Z/rTUL6AzHcJJrpN8xr3xdROr2DTWOeHXcPNA0gSKAaCXKASAdLiV6LAn/ptY6A63sFYgDbm5mqT
Ydc8Z+mdJuryhbL+RYlhu1ehEvqeBuaglXQgh9V/IFSSRDwV/RuCyhepL9pvoIzbOTGa41DPFSrU
KpvaBxMyFe1PiQejumQ3yA6bKlOh8L7rJ/zvoRH1N6zMgL+ykrEMJb6uzFw8jwDxV2motYmqc3rj
G05u6cBhzqVX7y1jl/IwzTj60mnGUgN773ifNyg3NPwOeu50reNf1g67JnF8Eg6SosELKMhLQzNC
UxqnYJMaZgiwZbxb863VXfzQq6z5U+q6GU3WOEuaVHFdU91jCK31fCFQL6/woGI3XOt5PBRLe0LC
lWVHY/3hPWvjUFcxRgi14NAozjEDukEfajP63+6iXC5WZqI2pHQgjSGwMGFb9aO+SaS3kijFE+VX
H7d0vuQQfFxCp/0w1lG2PnJwLguAhW4aXtQdJc/JlGCW7JTkk1bfrSIRZSJcB0YERnjE9A8egksU
PjNer2nWBKh+3cEootcjGqdMkVcOhac97Vbc1j9Qoga48dQHOPqQPZjG5w2AWStlrZVUzDjX9uf3
pkzj5ZAjZD9/hS2eXjI+phYbTRGJPPkRM8itXj/p+HzcJjhmN+ruFzVviQn+S+sUhh9RImyyNDKE
vJDfYjSZIVV/MGPnLik8yTyCv2cP2Z6JfLSrWpdEU8saJ6ZRKSGvIAol4p/bln6ai3ApYAbfNz8a
CKjr1lQoyoCy/my6fMQwQoVBHiKcMC2JTM0XEowjABUZxpzWdPSRQk35Cu7ic02Ut7JYtnu2yoHN
gIkGRIUDyPiaR8QYN8aoWnAc4rqCEPJVQOaMleUFA9B2/91RAmLGrYJH/10XsC7VyD2f5oqh7H/g
Rnc4sNUtOqZFcMKk7ZIv/JlZuJ4PQrbuKIcEET/MHxL8A2Yshj5N5pjHARELhG/lruESrDVbO4C5
tsSVds9hEa8T7YMqrIz81YJhXv6Z1+7RASo5jr//c7D1FwTCZ0saRSdFECKRD/4V6Pcv5S7a59+x
rYx8ShOajmaENlyipScEdt8kXqcFq9PVcvwoVjCSli8d2I/1+Gp+/U89NX31ZZosQ+4NtdZMkQmR
OqqyzRqYkxiUXG4NQ0ID1Ut8mA9FA8k0BJMjZQD4E78ylLfQ/d5zyFZ8Fwz3s69enu4f6P69swI9
rwecvAvtcefcOMBxYHEC77N8IWhl9xo8Kt7ZcO9aCZLl1/Sajnkhk2jRyQxehKUACwt8Hcop4+Dq
kMjEViVC0Fw38R4u8g52/tBMYU8ES2rHeJHqjgRDxdj33QIHoSSflORtEM4un/fom+C09NH3lkC/
ICROEFVISlk2/UC/n0EgwL699t9Nc6TUsbY5jJFCx+6WawZGG9wEnlEHG3QM4YGIKt5jblueSrqR
n7NiLd93gr9qFPE1f0BCMWtXsBij9x/dxwq8qV5cozuJY+NCnQ42rz5dg0pxZrxkfH1j6xBQff24
IrB9Ingwx1tREWwFeqN7ijeGb1JZHApqZFjmVyYwkqId5Yk0oIHUXIWk33NGqVViRBvQKZTUiCQK
KaizvMXXEEhgeNqZFXF4diAPfsDSTwJODIegfUHUpQjzBNiH1BOMMoZrwhIicOSJZAerBzmHJyLz
G/28pQwWrjEI4Vr44fPKMBc29OtoScyVL4th57g/DZGm1wkPyWwsZNfzSwIloEbB6Sfba4UEVE46
+FwYNj3T+A5aEad9SIaT3+s4sBu5tlCHR/5XUcdslx1XBfAjgAKeJvccJ+0jXggHUZe9LE73fs/z
E2uhQaSY+9B7YqW54M3SubQbzxvOQXfGotPO0PgC8idua9c+M2xdFbyCQiFqfG7auAL+ygMGcYrJ
8CnYZlf+SX7+Uqdu7FcEGdFsTvYRJZbAmkwjJ7YOGERDEdm2QYyNIdJX+4liyDaTSzsMOtvHtWmZ
dLdaljp/qvHQ/v+PZp49Z7UwZcqjJkkXkdQx5X4epOLnaM9+wlES0Ym2w70CS9+ednLREAnf4Lkq
No5EevvZpKu0UVVUKMjRw+tWw/6zbwiCdgRaZeBwIvTH2XknHHAJfZi2rBxEvUNthaGqtLtd7VFp
C8a6UDm8zTEwgyZbdvLyaDgshJGBe42gB3V1Adz/M6gdFKGkWlZpp41jd2Nyb5O6FqK7FORaSLiU
hqv7cAhNU6vQa65/+XZeu6h7mzlmuSoG7xDWeXgP+bXM1ZXQ6ELsTw1SPGawyhjBM1PsOnceO7/9
ZyEk82ep/LkHnp1/iqnDsPVdmSLgSLqRHCqPeFOS+BMwTCzvqCqFLyIfzhC/JeqrUUa2ENOWsVCc
a5++vQoJtzZI+ECZlA+LtynjfSpcAsbw8QWhXQB3LN7FliEKLqNtAx6G6AuA1JLIf2Xot9jfizAT
q3e9jKQv8XynaTSW3ttRtKuD7PnjCn+cg5o514MYsvX8C8Lk3j3wkXms0NtAlITkHv6SHn67J2rR
M7YG4cTSVuu32J2+nMl8EuS1ynkZ6FQ0++isEq52TJPTZoIJKrnWAtUfEjr1CAx5aKN18/IeXrWC
BzJytpaCVoYCDikqDvLxkdbhcvd5VfmHgMecbDmXJL9SvltAcT7I4kdHOHM+6u+iptxA/n16EF4h
BVdsH94Ome99DldzYJNbrMZFJtRq9J+mDcUtoa1DpasukBkpDnIl9gx4rmEGN1SokgJkSUKn4tNz
HErLt8l5mKqmluB1PHzf7jEGGzEsh5BiJb0eK3P/MUNH6kBb8kezTzozhRq44dqDL3mFGtj8tzaM
u8QJS9s1P9ewmhlyarLNRI4Mta4LdNqhWsydYeMYf9nhNPuwTy00Tg7tCsG9RZInUa8QcdRQijMT
z+/it5UQek6JajH57JVn3tXYhiU26mRlgPscjroxnh+VGWXd2Q27RxAqJApILLwn7RZUOfH3t4zC
KqfpLA1czg6BPR1ARpuH+LAhcOauuebmp/xUaC5qqNq9po2xkHfeJrpXxIVKv+LiEDMFL0cq0P/M
WlqcevhFhDXpRn6EzdwuHB/fruNt1gByuY/spVaT95oXh9R8eNWdD0iW/uh9+1REAiqIHc5LKJWF
w1KVxWGBMIdQkhwg6GKv0u0lJw2m9WmPHmJEoJPCqHhkrhBTOP9bAT7wcce7uvlzm8C9LtKgleSt
GbJY3ZwjYp7tUVv8WXd5e/iDp5hry1mnS/CUO3bEQFD3OqPMIH3yfJ8t+6XotlylrIqMXLwbWC8G
2zHLk19VjTYOm/Mo/VHvSfgOsAVqZ/Vp23jyXhq8InRHALX+Uh/6S+dHbcPrc8jvMAtfdmICpQm8
+MNCYdDmfFWb1sctmg7X4I0XVh0T2394wSZnbVsWdRmqWeTiu4czOUpGadvB5loOxS6WqM0KmWnt
rJEUnkfWTVcAwx/Tms30d0SawYFBUmm7bxxlM1zcyNyKf9EmHgBPdKxiou977zCbqcPdtXEYuhqd
YgszWx69inQwA2sx/ljkhpX4zA5fHlgxwaVj6ZUaHPhJzacMekHa9w4ia47EavFYihE7VuH5J5Pt
kspyfIfbC+jjhmpItknT0eGDS66iHZ7e7dPVZPRA6m/6sAMXHCKnndeNZ+pea4vlChiav1+ph8tp
TRxf7p4Rt/77tFu9M5dIwbKphxE080pBZ83pYTZkWkvyWt3cf/+/hzUThS/Jgrpsu/hYpna5QxdQ
p9hWuuR5WVBCObyGUJt92f4/oYrfh66gMmvW3Ft0dB5Woim+YyT1bqtvovc4iY3BPlsvlxZBXNB+
b9TVF5eGMFzVaWpbKFoiMjMNjPrcoI6mW5wu4sgcGsaR79cjjYc3oVF8I/QKnY1QrcGxCE+TET9r
YX32vKx0D41l1IaJiTwpDpi/cuIo9GT71ps/a9HIrGVMi7YoNcbQZa186DYshdjMwKKKhb9sUkBw
OC6kITl4rwl9AUssccDe3lk/tcEJICMGC+R2INMIn9qylZ+eTy9BGCo0MzHE/lQ5VD9OGQeCSpZr
sTf2U/m4zNK+fsQlSP5DHaNZtHodVXEOGGXf3Xq8i3zock3egGndB4qeHzWauyQ7/1p/RUhfF3VZ
QAbvt7fZpoqx3U7ZFuyGObM9f9P1+xD0zSOSGExUAScyl+jKdtW4N5Tn2TEc9DXrkJpg3R7HHg3d
zonomjZcT3xobwVNc/8r0smp7IB7RQlDW4EdSW4anIWswuqEz5rQGMT77mn4+LAGm+xnxvJmyb3Z
j3n9zghaAPJzuPc4BUU0DQMUBGDPms0OKvmUrRizmQasthQC+SDIVlS8ci6pEmFtu2jJQjj3kvqX
vTrWN/rTxkNEj1Co2jVm6BIKmtyi/gYUI0PAFS5CZzJzr6D2lsJ7sCeqY1McS3xuXCyuGt9MgVEl
+zWIFDq9RtC/kDXbT1sDneHm2M6j7OfRP3Bv8feqBqmzImivQKa8sHUjQ/VAjZ1V2y+gQ2EglCjH
lRCFItInvwkP4sdjdDfd3V8TUGRZ9RZN7obIuZEMKb2cKZ8Mj7gBLKBpg+2/m2Er1TeFKtY7zyyn
aZMztCTHVvYUEI+wZ9xfcR4ZR4vmJslrLWoReVo2LZSO61ouWm5TZsqBwSh5U/iK6OMlA1poQZAo
bvNRj6/b1KxmvuJyLl6YOkYiGsKml3TxzpUF8x8jnbMHTb39vHR3AeDqSt+AvP85AXjHsPpCrhPO
uqTD7nyP7xaJIJlHV1wF63+hWKAPPtOZUu24Kk/lOWjZD3lLgl+1oals1rJUAYdLsLpLOcKzJX7X
PiUOB+BihGjrhGbifvuly1Sl6UNKv61vVtl928owKwJyFpl7BiqizRIza+RXrs1S7pNxHp3jS6Ak
sF6yXhDxf15jq1Rnq/rZYvG/dWFDIsCMf4fENHYgVIQnUJJQxCHsyA7R+tA7R/lsEN+fsI2sWl2F
o2omasvKbTgp/R8Dzhk0ByLrMiMe1X6r4yX47OAuydGGA8FmbQ86C5l7y2hx16uT5uO8enVY3vz6
E07cxSOrgL1Zrp2LmlgIc5cfnmnCKTdG6WIak/E7zWRXekRAExWNIy4P/CtDor9tSJGdiOonQhh+
v+VpEZdXrJlyrg59DEBjiEDZZD/oJeu6TqlxUALZUcF6dMlP4yiryuS080ko5mtAXxFfhnsHSehY
i8Zsq3l0vL8crOUn0fO2HExQJcsXpiILq0EP8vomEHiCBO05FxwUBuSbyStIVyn+oCghqAs8Tkjn
y+4dI+xiPTM9MBexd95VRD7EViFzAcMlqt+AgpNs5pr2o245706BmG+myVKBKmQfEvA1JD3olpIn
CoEOD9lr4xPMXd4YtjJwsJoBr8ECRf90qed5/fVZqeED2kTywoJXQGrlIzdyYLVfDVFgQdHSX3N/
vAjmhABB/amH8tvWDBB8aMlfN1EztdimxJ6SMaQ0BNP1ZOaT3d+XCNZ7gK9HXGSE4sHBL/agikX8
9jiBy0enVrkNUc3tZuI+owqAynGoj4KtNxAR90aKQrkX3XpI7VI3S51G9TLrsV03JT8VsK+KtC+8
6cz7CFfr/2ZRCf37I/R+9zNa7k3MrOq9jZ0D56AQvABxFgp25J2qVKdid1NqmXWyAPrs3A4Gdjf5
aSZ74Cib4bCSCcHuCTCkzRbIC1EDp8QnNAHUWhroTnhl4iySKTl5+bNxxia/367IlhfRlB7IRuSe
jJlm9mxB76ZtVzbtI7VCLvFm/2w7JLS/NDmpiHLPiBta5sSVPzSc6LP0ropxUEk4HZyT2APGVsmz
qiqKUhSNa0T2vto+N+ZT7d8aiVeYR9mwSudtXB6xMbUWxap96B1Y3vdUJtP+HTgMAcV7PZMe7IHd
NxR0p/XoJXXDJJ5Zb76ggLjAWZAvIArmZm9MpioyarW9CG6whP72HPaiwRJUOziVJ48NPi0270w2
onXUVmliAMmrORMvYqII6fu84hmiNtTh8oZohJfY+omrgXa0a9tqeHMt/AY6xdDk8sZzVMMgU5o9
o0QjaLQkP+PRwrmV2vrOpfwwWUkhcw5WNu8YiCB7ZVuB1LpSdG/tPOdzSBD4Zk7QNVNOJNbfERp5
mk6s37ecDqjhzL6YArC0pM8aV3A/GAw4qflkUKRmhXkJ0wvjQr6WtWVqnZny11i1kvcK/UIkL6pZ
2e2TrWX8rmKZOUM/3beHjUq5CtXeBux1m2hy+5x7K4sOeSxWpQfXT/f9SNYglpxY6V8uvaKLOaC/
ZR70h+1zL5I8gMwYFJ337v/kCGmVHx+qY5gJVAbkKDxQPhGo4XaPI9iQDN/4Rxjg80Dk8mdmYXSz
Hobj9+DVOp5io62i8aiDodzbKR8VCI0FbzrEfVwBxOSrecw10uvEBWVYehykgS3rm2BA0F4r11OB
sopidS302g8iKgTBv2HnQAsIq7yK47TcKtorBNX0o7vErBmzMHC7kwOBCBAl9k0wAO5QQOxOF9kz
loDV/QKCN5dCazU0IpzASgQssNcPvxN/zOmkvLIBbJPyzMJKmow109Y2PRlYjFO+s/wCxnNDo3hj
Wk2GpvMHWCKYnAnjuUOXiRva9Rqy3no35FP2g9GwIBH/apedMHqV2MJ5M+2iREgrzYYWiTaBvu5i
dEaOTtnXvFQFzKk26A5GP3QD3F4XslpxDmbXEn3X/VQ+CMO2/D6FZij/mYXdcbRnKmcg8jSRWA/2
MVOtGPzy9fmLjebctIUtRI2FUz0jqOlD3xY61yujCg/CRitylJ3Ryp9w7FAF0bZ1w610OqIvQlay
dUz8IX/2/JaucJXy+FT7ZlKoQ8bJ1bV2/xkiaQkP5npssvAg1LTduuTuWxzbfkUc3Ge4K/nPJJYn
iVHZPrr10apUE65ncgnxf0GLH6TwHJ9WRPaUV2BWVGjcn7U6tjaAZz/ubvKJZx5CxRc6Y4DaeS7f
OURNJumcND03nBlsgMqQ89+GD93jAdKJT3E2A2MXKVNjbHXMu78AN/5cZ25G9IAKYHj3lHYqGYkj
hlRyJkpqZ4bpbMB7FyNHI0VerkuiEfZkEH79CAqLHhAEdAbYj9rsNTLzJP70n59CcpbZmv6oaDmp
fskDWfo9taMb3DbMm2mjVUwuIC9s46cC5OcWkrKds8p9S2qzsbQprUpJekQruM2BQjMg2l1i5Sa4
6wNH19ZE6Yl3TBEfgTidhk3K8Ef7/s7kwZtBUH5xV4nKhJINuwJTQaiXr3S/5czTB6Y8N9jk4xsZ
7BPpOY2HniFA1LDeYyNMO/2krmr3tXZq0g94h8XBrOciGeCcQ3PyJrdOo5ExY3XUi2jTIW62VI99
/FSe2th5Bc6p/qdp1+j8Yc9m39F5AvwjkCRDK2F99c56/nji5cTgaMbvEpE6W3HkOUw+WfpafRJF
T1EhVUl8UgRoeNCYWqhGOclHG6TsjdLWLV4iTY8IfIAUzntoYjpQ8TEV+0MtZ6m37tXn5VndR6DT
7b2xoHR9Dr1N0CocJ0Q1ZrHnxw00wHufWbzQjrrJSem7MFDmSwdOz/rCPrRkxwX/1Sv8PlTlcJrY
GjGXh44ygsVOqIaGkSpQjErVPaQFxeFg4sv525ltbIx1bffoLEfrBqgAHM7CDZreM5yQx6N+JGnn
oWBK9DvLJxzEc00PUQfPsXFPVnLfp9bveyzE8CViBww46kk8xlYJpxwYXXireMcdKb4NHBB9PUTD
8jPT8s+MFnUwk1VoYh90BogzOXuM7TuWy6jU56MnLJOrkdy7oR7czl/+KZtlmTpJqczFjOO9dpVO
AKqswqKQ+noHwW7uHpnKe5/3eTEMW2YFx5m25ekOpdpSuLfZBcJGzcZgn9C5NLGcoAYYHNyu5BL+
ZC0imSwQI9aWJ3H0JzTNctogE/APbaa2s7rHpJYDYIdgL4x+QEfjfO1RBW0CsljEoj3nt4CIxWGZ
tfpXr2s/tXSqfjKYRQd4ILXgUvc3FZ67Gya8ztwlbTtIm8CIW9W4AbA8R3q39koeRNhbL/STvvuG
dJBLewNFtRgY54nnIw55AjyFKF2Yw2aCTsl7Ba0wJwn1ZlMRYSedI2/G9UDiOCrYZhxlp5hFCNFX
vr7i64NKIG6QDrhkNTvhabn/RETGAruRIBqbX1CDjzKBPCWA4sw6nhWZESjFiX3+JriRAe1ub1SY
ejL2VhGbnlE1/DCs0drHSSNsTJkSDP0P+Y7ZqU3hDaxjF0MEnSO+s+kVq+16eWKMJLDHpUcl51Bk
jVMOMjzq02dzsbpynp6iDMLGg7FT827wNyy2oQlF8aYWJr0+ryj2t2XVUWCPTMAWmgThQdAJm4jn
qUVaWXYz8mG5a3gU/0dFGdzVSSCFeC7c2H5jNaroqEQ2xrR0z//LRlOrY0wek/Gu8SZSNIIwKMAc
7w1dtwHICt/1e2B/PeXaLpX8avgaxCIgghR+lx6E2rpCQRA1fH5HqkM899IXDBHphPoYsb4Rg2SZ
zOCt9gZfF47oTtTDqWirkomAAkU/QFwhCeSizlOdGI3zXzUB+/PFQBD0CSJpBvMnWOmoM/XQPdc0
Q+Dh+YFQs8F7tec8OYiNAkBQF34J6cOkO4hXPXHbog6WxmWXqZJR7RtjVJtzjbhFhv8f5uEn4huM
gGyWMbACcEJkr6BQnCpUdg5IJ2FPKIjMnjQ1F+xoFr++xAy4GsIfp7YDnnX1HKVlXlPAj2Yykged
LhKbmqyuL9j2TR42FKWlD6aMqUgUtFlRmw2jgq9dJ+8u+8homDE6s9gWhfIt9EIfHyzpF/PU0pk2
jtfntR3xnixwHHcHKUo6gtmf7VNcjJhwbsbznfvldU3ZM5zL72QO/vNiDpKm6/AsQ/uchtkL6gwd
XAp5KS/umWaZw7nAwhrxVC5O84e6vasoNkkrsnaUtilapHClXI6CQ8uvkg4YPTWo78RbeTJQxcSh
Myjrf0eBwnTv8Q1/HNgtewfc3Ey7Qdey1o82wAGCjgY3bUwkxbcEnORwD0+OcHCQHHmMD+9/UqpC
7kAzNNNChzdKLhCjfkWrXqd8EmjLQjA3+pFwKaWP6on7w5xoiLQQVElAEVWogEAdt0bb1LDAhFA2
oI8OWZR/duBFJW309myMDkWXkpy21rH4XpbaSOpdcSDd4WSTnlcxgCMrMbRgMS5y9UYPLrPLdbai
M1ZO8vFscs8i6Ptl454lrQEmhBjwXTr0e0ugLU9njaQq1cJk5H5B6L58bEMjrekmWYUJagBKhUSg
i0CoDFixxoxF1NJox4M9tJt8IN7iXMDak0NfFaIg2hNiYeWbxoWlAPyAULv3FgyoUnT0b3RrPrFi
2YrlXhLljdA7ISYSzRxm/pOaK/SFe7btZ28HKYGnHteSZMIUsLsi3oWE8Zl1gBvvSgqYy9f56tBK
Lh2S3vCIVIEVnH7DkCfQPeaFDthNs7MmJgh1B3YCeQDi3d7SySAN66vgfXIXAZH/qQxtsL0m6NIi
qjkE9KCTREXTKzxVd8eeUCHMrl2ZMhlFFZojjEbpymdtJzndlfIPLYboSn2biFv/IqGVqB2c6Awf
yvoPZgCyqo+WWTxs0LuFgWDryzeTBK1JwGdwelTuX3Ot4GWT3SvzvioD4RBfa0pU6A2vu/+0QYJc
cHcRwEY7cKpwj2rPmEm8hw749grWueKPFhJEeWpaTzYgMnDBdeyjEi6iY6KaRc3B5cMPIS4GpjX1
GT/0uQWnZWOGJvrmH3cTPNW2wRZpH4F25M/tba45C2nMgunlwO2TzVTws05IUvPQHMc6YEysU1K8
rjIe1iwd7yuYirxQHZe3iWho54AOH9Cr/v0OmAUzB5AYiAAUL3v+vaP9EPv6Rv85aEDUSctmuU78
JS1/3SuvpvWjwUtELpXOGqnpmxyKEI5R4OadvTweBMhNdDKRM5kI9rlo4tD/MWZ1rAvkxb31gq+b
f+GbUwDnQiHQr5Pfh8ez3ut97Z5IW8G3apyo0bCNQq8ZI476yTC4KbFRcucb4BlhEFD2qXv0znqe
f93GSV9ijcqyo56jDb/YK5XvYDlbRRzeuiDLVtsmUaih89uoqtj7IJnJ+kCTB8wiOA3pFKxLPboN
DmywnYL2iEKT/c2P80FmvfcB6VxiT9F5x5kNulmg9iIToDphTiHIIUoq2zDv9VQ9aZjkCeffByGt
yooZWkZqIebeUTEdTVoSk8B30zzUq70CyoZ0WzXqfjFwblUDisSR4lZpH7XCB50sVZRCTlhh4vJD
tklgqDXoNMb49iYI3nhJYa1KYMU4QemRAWMQOs2nX57q+Dpn6ytkof2yAVKEuU+/wkUlwOjz0XJS
plTIMRUFYta5HLoxLcT1BmZg5XqXR8nC8bGuAkxiE2uY8aEYdjuGRBFRusACiumM4qyZ8OZk7TuZ
gXbphUunnE8VKzkGysHPCLIXoMMenwwhmP7Y2XHfOOFC7b7LYwPl/HTWky1GsfBV76L8b0+3JdN1
eDzDwgF6/rti3TSy6m7pr2MTFE9apFF97IaANTyMP31zhRjssFwV7epxpoPu+G7enrR1zVzFLZMe
q/JN2xrZjsG4yVpD2u4hzB3hKIWc5Do2P1iTZYg1W0GonJLjv0yjDDCNAqz9EMEUqk1VJ5LYiGz3
pkAgAB23iea/K3MpLQ/D7b+CsGR7z31RFIdXvk/5KLsEOwGoNtdx2txq9KjU6DkmwpoUvFhapXy/
ZgAqj3RccaMLJwyvnZjvbBW+DpKzJCzDj9ExQGGcmVsntFQwgxjcLXgGocZ91wAEjeoCa1z8nHnP
1LUzX4pzK7yg+ZndbwFxE2/ZMhMv4IUAQMLuFI/7GWJoOkGCxc8Ri+GQ3CLNSdJ8gsH1yFZGqQQ2
udgcNigIddP7+yOrohzVwkPsx9IufnjNHXM6iNbYhAMmelcmabgHg0gk+KIom/4Mff56XjG7JSmh
E0NqF7pVYoZH8Mnv6/bSda4eB0TRR+aH+8AXI/ePZdL6r7OITiTnmxWfpwKVDmTvEkObrvSMVO+6
3VBX6sNmmcr7nEZlYdqbH8KL0kwvMcQh8vpTw3mChWx7/x5nRkrj8ibfB9C95UsCmomi5HRWso+u
dP0LskNFKSQMWpbZEBkd74vUXjqvL2MvZJVwjgyjUsSD70jEbcAsg1/6KcjDTbzBEWQek0HCXBe+
sG4SwIPP8j+hWVm64KwRkWY7wExAoxajTUEFmV4QGbLR1o6t+/TiF1/nzrBpJb/Lax0UtNlkRKu5
vFZ9qkag8zaKXMVdHjHBfmXkE6AN9ZUj23/cmWUxdzayI+6eocD17q9Lu+Hz3Nxv185aNjjGjzEu
llj6pTBxiPwlabtRHj1PsEW2FtqsVKY+D10OEusuatzzp7ge3QwzYbhk6PnwTm4lwxMZIAy54no7
gY9QHeVY/gzA5aW4DwHUXwcRZ2Tz/SamrXugaoxiavBzqezW6J+WTt3qn1bu5LXcLG1Z8XIyT2Rc
kIFs1y6Aq9WR/cXcF+SVIERdywECDOoheZ8oVqcmkNYjJthHQuPJ391Pqa5jFrIsPZVS/AO4Vq16
37hmDkbgSqMcVokHLXE+tvGHwrpYc4Hq5uGGgT32WU1u3oNK4alrYaRAeXOBwimDa7nWugc1fU1e
4e5XLJ2chBuAGUYh0CZdZKjOoffqGhTN3JWuV3AoiBwePKVdYelSSe9VXNRMWmaGWEgAXr/qw4GM
OwFylU3AuTMAJGMpThGUKQ4rIDK7IcxCpMcrW9lHkncXA5Ta/VeXgEo7AtyfIxt4NEjz4S5zb13p
IZxK+KBf/sgn+jGuVdXX7iQ0mVQIaHR+DMku2qs3w9EleK22Ykd5wfyEmIZEFc0dhXY0mM/2OH/b
wLv3GpCOkBYuaALkVsDB+SMO/rngJ7Y/sDk3sbs4kJ9u/D7i8K1BFSREy2BAbU1CO27XwSVQK+c/
BtZK2K0V2nH6jhPMIwa5FDv6GLJoKI7Sp0ycguteWey4KJTFZUZBEVk6GzvafUoTMkxin02ABVH+
O7g7zGmn4RnUB0oG6cEWUMcCY0w+UFKnOSJW+JF1IEqJR9YBpgRPYJj1xF7WNiKQq244DWAiCreJ
cYguO1NLMS8GP9Eplpc43aWdDFAcpAjytWJ7c5/++6BAH8njLw3MHPmPoPP+7gtnlT/8+XP1x3T0
HO1G4p9HW0FjfrXLnUQaMEIKauEF3LeaDGtgXUJWQunlRW1ZGoe3uPRtyZ4BsB7K+aoz9TbrNeTn
6ILjeANlT4ktP+4ky0pO2v2j9YnIjFFHAE0F+ageju+LsVPcDGT+yI2V3agY9dGy8Wl7LvjMuN1Y
zcDMZQH4IRKk+WmOroRL1pkIlmQSs7ex0Z2+P913IUGznRjRyRJzSmx34392KxRggiYMMtk31ZHR
zqlMf3q3l13tekRkPqcuVhj0RCE2TuYocnhkRLSmDoMKB5ZxlmrGTJhvufS+OXNaCi3NHGEFDry1
7D2eYNOO35nulUt8HLLz/pZhkwg0dnykHxvymk7A+Oin0dJG75sf5y+NlwSnmkPmJquFQyS0MaKD
9SBQ76Vixp7p+FnWulc9ysdgukatVidwvOQsUIUqi3lUC6gjgAotK8M3wR+d1pfnofSUTK0L4qHV
QSQCzYgL29J7QTyUSFnk7EHxXyKYkXBO0S8gIHjyeaIqssWPLkF4V9Kv6ewcZ9wybvBy6nKIeG0B
lLVYpviJRjENBC/iIWpqvH08sCKKS1gCvBbp9uvWajN8OZxoy0+FVYEhR0t5Cy+KtSr+WL8dhUQU
9CGWpaKlQlfJ/Fxn5U84jW60tpfJHITquR6/jR8DtHUtJ99ViBEt/AxictpQoTr1FBWugvQntoBv
qFGd0GzoEemE9xI6C6pVeYhHHc062HZODYZB1lxU2yC9ngyW2uMyy++z9CnIe2iBO8EKZaKQvu5V
7wKmlyqoU0ab99xzOOl13/DJ+fMT1nBbeSeNGBbGGRnghZyE/ia9Gz8SVYA/0cRAqt9uOBcDWotZ
MDYahhq8NfodZNGLJk2DTu4sOxeRTZ8DGrwBWWXtuyvEEwmDB1xyB95+1lD5wYq/A5ItB7lpR/Ga
xKT4jgZmBwqXeDM9b5iXixbTxaeNTAheh9xQzGQ6PgBHWJ93w4kPI2mYjdyhVR9+Ri4i7AmbQlgK
F9KzrrNkcE7oDl3w4smlBE3DefYPFeSGU6vG1Jt2IRFy0MglaPHnL9ZrMD+marki2LrRliGbcIy6
LwwSzomQmqldOtkk44LY69TRRpSy1JKslSr+3jIZzAgqo+gha5LRh9YbDuvUUD7udnOgYdosv0lO
vmWOwB3w21AqrbGKI639bES1gll50VzjRaxlFnFoDZxlfYrMDDBKCX54ebs/gOLTLjy6NjS84MiM
g8AEGsaO+l/J34HSPmYSfcfC5u0inIOCmQ1YVzE+Dc4wrg4TspwfdmsTVYaZMLQcT2FJQ5pHUoxz
R9B1gXRhU+KGxyN7I9fQ77/b00BZ85FgFHodZDdI33K9HelIeVls3tCKrnyuBOcnSkzYzWwL7c6j
RglA24RL4R+xjvZJp8QbMEjtsg4ts6zn/VJyfEAnAH7cJ1focwpIHnqD5m4PNeJDhdCQAkTHzVFD
Xn4pC+2A50VWfH9mQvMKn9wOxO5EOB4FJBxOQQ4dOaGrvaYPWg5VGKXAvDsHyXTK/ANDM6bbqDE7
05wEeCUtSXNJoCX+nc2cMWLEf2V8JRwnrhNocg0h6a5BT7ZEzF6cjxBnraUoWqD+MJqb/qymdXxx
bEMG2EUttkQ/Zort0EfxhjnAKRCU+VA8GHRjv2CQ8O4WPt7f+f/Zj+npxmwxNJam6sM2959SSVbP
kEkgxyH34nxx9O5RDMIhHwu83pI5FDkf5roadQK3J+lpM5Rh2BO1KrWiGv2YxDcG1luTcq8lbIn9
vjDGDjOq5imhCoi+0oj6ouuHNmsqowu/ij4NQU1hlN8srdErV8KlZ/IFb8KPKyhCi3jbYotH/ExB
hoXvD4FwjouKe3mmkTyhjfwT0uy3oy/hhCJQ2YSgS06mSUpUBDFri/cRWonBFEF1erxJ7+iFELgK
xCJUuQ5jEyaNhePOBvKmhCnUSykh2pop3oCzdbWyGOwBt1idaKvwTU46QxwDAvuRnkwcjk1mXwck
v52sRRVROUWs1vQuZtFTo6JQ2l5Cf4ui9X3BFlyornkNwL0EtHcNeRfVu66hPJTN/lUw1Xjdu0pn
FfdzsXl74Dl1rTDlRWH4acmhQPprsUS0LsXIBV6Bq4ad3lItEpPkfRwzn901LDqQdit1AqhRf5rb
jmF2jsU3GT3E+LZiuwV542BDNLDFZLqgg5nV8C3gk57UTeaHYzOablzyKtfSSXcEfCyhbozGD3jf
oPpqxH42dwzhqNv3EbdKkqGUZeE3dD/9wqKytQygSABTElETb+f61mgwjJPxarpfOAtZ8bhmKY4m
If2+fVBNKjWLQLMRcPLzjKW08345lKG6SGpi6+tiudHu7SMpOWSNGnalifmoWiQWf5q/E8KtciFk
PCUcAMZtMnqjf9inQVdFJZ74ZMIvwHkp95anFYB6qxIRR87l3UqVKg9a6EgzhT9lzDD3VAryxP8y
3VgeXLkyNC28Zd012a7/FW0S0Gbijl4ZzcRuX8KE/wMkJFp4NQuia8ik2v2FAqq2BjhPLrMOxvk3
FhpnZc0975KNe+TbuquLUeG+RHRqB4ZzhJR9O+lJGEYeRHI66UXeNyzSqn/cv/xWp3YaA8CMCOvF
Kth084Yxa8uoY6guqjECrMwXLMy0Syd0MP7HJm8JC2/v34UHRAg7q742mDVLWzYu8blilhmRidYL
Y4D9kJwY6XeG1+78J/YaJ1dClUhjSlCav1znUKweXzVRHrzg2I9HG2VXf8o9iAbRvTO+ae81wefm
Pxh5OfB5kowzDY1Y7JbYyaJpRLCwWU8Z+Vf+KOmiOrkJuwg1ta03ObLf5nCKSLJrXrzxj/BuI7I4
93/1uEdmWmcz97L1MHxE/OoLfEaL4WdHx4n9f4+vmEWA+meoXfxl8iii2sy7/vaTVvnlKZamgTnt
wm9N4FxWayDRMqGu2i1n88+KB7w36JfJA6v66ntNh111sLOzFuF0uZSYeWlOUmFN5ModlsuRV21+
OpMgQn4iBzlHfMKmeIN/B/0zQGIbOBHZEnc+YlTmIYeLrVipNdnFpkU4gFgn9O2eo+7lP64HWkxr
4Bd3dL9Ehjyf5q6AqgwxVsQQ+V2DGjs2i+a15nTXtzNHrZFhliY1u3VgnuTNTxrY2nn+GmnJ3k5r
FvbMcDjXeEfq7s+ILRRhMyaOuVAbM+4DH2imKuz28Uk99gyJiD5VzqA6zBWi8Usy+xtFSfOHXVZG
VNzWh7RF+Nd+hVpmcWrSplcEwLuiK+0+nKqC8MdSSeS9K6zHNqYeGMAFXsTWpJ3o+v+wVvx4B7kZ
46Z15HLGc+yiIB4Zob+lwyftKBTtZxtr1vkoiAweEDGWubBYODoOOOYM+v9Qf2TEsrXVkpHNTKYr
pORIxfse1cWV7pPD6b4GhGBGR36Ta42R3zlQqnTlPQX83BLjQ50u7x0Ge5Vl8QKhirLEmcN91Ulx
Y9y/fzrSfawcbdQL2fsKpFAiyncmN0Gej/2XT2Vx5zVrsSTVonHLK2ROTKlajIAGG2ZvKwHCbes6
8NhKET9U7h2YTRCDyFJfJdgaE2fUY8By5v5Nln3TZAYCxKrXyohN+71+L2NqgDpXbZiiAc2mJF4M
DrIE28+TcCzIUNC7hU88kZH4rCS0VGfS3Vv++nNNkaGBR3n0y8FnG4CpE0wCrJdBLC5l5Su3hizS
VVKc5oVpsEE3+mVRbRrdiHWoC2ScAb7grq1712iZvb61B4Bd74ERSrtjgtLQmSl0BF6S809RGKmB
XVlEdsFGaJBc43+medUEre/jZAOcly3wy/RMX7VHADJYq+Aoysm7Zm8OIb62ceCLRI7CxBKCO14R
n9Yq8PA62ELSZHHxZXy6II/OjUUfRQ/wCjz5uXIg2YrT4cy55tqwrYUAWvuB9unKaK8U9lUnpTq/
c6KpcjmIX3KRApEa1/JFlKknHYmNiLqZQ1lFFIXoELKTYhpi9+tI6+F5wr/e90AVRfyvgzgbB7ma
Kt/NdCMmAkicBdnWnQkmxdVIczseHW3qoJGOU4Fx24xVVoLH45yP8Cq0Cu+EXne9aAZGVTolvq2a
SB3irVGkh/AnOj3kejNz9bY51yS60e2gJgMNSfCSFECea1Je8/m/yCEJ/J3EPQAHrIFH3DFNWMZk
U4sapzCr45f/VfD29xFOXWRQFRHy0eoaOJAa3DxbF3g4hMetqPDC9STKoIe5uqWgokx/NJEwbJJg
RMy81mE0VmbcMarNvB1h6sJh2oN6nHXWQsudsEOEyL1GOSuF4AKAC1mMVbiGDh34WHgz+kNjHiBO
50859pURN9n9ndITtxYtWXkDvFtaEdHsDRELhwX9aGSF6E+PdeUmMiWm3O2mnQtxUVAS51AMx9Dm
e7TTBDHXibfNlBV+kgYwh8dq9gBQSGSxJWY/bQJjfkgIDWotEUiukE7onNomfUNbqH1PltydDESx
WZmcQiKXYt1zmLQqappl2k4mHHKbHvMUDkvOicRmyoPuwwsq9lYOdClc4USoIsYVxYkJlOUXHmws
s0ls2dpbFKxaKYTzYGp5QSdnL+uADdE0tIwxHIZsMmX7meErTTN3ZYuTgwF3ULm1FEInpUvAWti1
DNgtylqWhYPmkUb9zXVqN0hQQDj79pM/262/A6aCxCMUChJ94TjosI1rWhCy7J836A6b4ys7OZ1K
iXGbVI43+Pjn7Rk4sp8yw8VS3wrnM4A6yALTGp+gx4QfuDZkt4PXadk34BwPU/IJ45/wWtqe3OuJ
cPfQ6dtO/HBo80XAy/KV5ytnRuPRtIhZ1ekn8OKTfRGs9bQ4nR0ZbjIaXL05LxO34UuwIhBrEWei
oF2u9Q1tx6arVJsDWi6WuFXjMjf7braP6j8F2GX5+SosEbVM6pP4qT4Ss9CxLGYwGzOYiwAhJ4Pi
M9MovxvYMk/DYzgPx5ZP6ygGIq64ww199csjphzDYGOY2PDnjkQXD0nnJN0AAEkn32rBIqpE7zxb
K8EbtFLLXJbtZJa9xsmdOe0DSM6xfWTfAnWhU1HRvcmE6E4ekM+8MVrknPHWobROwXX+zBvYFU2c
J3WeR8gu51bE7/m6m2uxW4j4T2mMOqnzNoNAydNp8Zbo+5B61uMpncpX7ulXNhLkbMucx4yLnLOV
RjxIxpTcmAC7mpNBuXiuQ4kQnnAWNaLjceInI1dCPaJ5AmFFp7YQs9PXBy6QAeCi0vFp+eAqCRdD
amkCwNuWu2Oqx8qrKZy8AUewNt/MnjM91gC5JTbcvUMbAQTXLn0Aur7AqxGo6qgpI0FY2VhB3KIb
mMJ3MWs2YPLoKbLB+kN7uteyeHq9NDJ5mFNJm57vI1g0vek2/tbGwxFe556aFt1o5XTKH4WH2XJ4
5TMsTk7/473Jq43VpPByeMjlCdveEF4oHKI5BIXCcRR/J8auUIYWhVEVGScfp+azAh1uLUlbl3HI
eWjMTwm3+1Csd0Ao+gaWnQev3zAXYn6w0/QovPKGqjF54OJfg/tiH3ppUjH3zNXqZ9OVnYC6veZe
vg96WLU1US2LljjA21eDOOMSQf6AvqXxrK4tUrvib05QbtoSaAL+jt0T+Awc4SCSpcg43gbCEPS7
OagsmXg2X3n0bXT+r7U/19U51rYuF9QsvBncdchuv/ihlFXC64E3TEVErV0A6B4sGicjpjXtmvVm
wI5N0MpcldgyOAYle6vp3E0tLcf/xrwh7oowokezibkCigRRqh5P0+CgJgRU49sT0+kPDQc1mxVs
3JwkPsz4sOlLyAg5kw9QqMEEcXrq0PsiEFjBPMmmxg7Nbg9aDl32ch2RqizN+IJAlGwB3aTl3P0K
0eHeqYGzIodqk0CwAN7A1EC8+4Uh+3b2G4vs+24kyw0ADYMGfMXmfbbCgzwKKzc0CbDu+TFXlpVW
Oq1j0F8FAvgSrRc+9F+oLaigNn1hy1qqVKnNnvW+LYh2qGsf/HpxcWL0vEmKpjQxD5vqD/nIEBJW
FYK4GodXNwGQux5yHkgYd3Wb4eokEpLYpsoGy7pHrVc2Cq3qK2JPxY60YpcgNJ+UXyS9hf/JublH
cUkBequg2XhcNRkSvIX/aFgu3rCixL/Joi2gODJVm5jiszfDFKpRefGsbXvtx+ym1k8Y2fEH/Yu7
lXKf2sjozTVMCUxQvXwlLO93JaoYEklFvcIesZjHzU7cEVhTn/8gNGU8zMov+vGOQ++MSs9G6i3Y
2PAD9tDMuG5UmHOWQrWfGDi2+i3RUBW6o5dYjZfxXKkuEu5qP4G35RtTZNGpvbwkDfxyPLXBkfZ2
9WfCqCisgtGsHF/rLD7VtXp+/YShdFRMPMyvtCLsiIHDRzQD0i+wPNH4DfonggSvLnN6mAnjzXiP
Z6Y46Wb/QzcoNWf8WE/DMbGQnHVoCdDhneoP69BcWEf14FjdsFgATmJGAngBph+6HIbwGE2BOJLB
u5Xye75XTU3gMsoaOUXR7/D66Mf7C+o3K/Odc1j8/yn6aPcP3DWabKAoeSyuqEqqLN9yTWURFSWy
JuEtImrQt1Bz9v/UpGyHiXLOy3KUJ6V95exx/2iWEm1OzgD9md8iTdJnmLZM3WjydkhMKk28WqKC
Fbsx+FuQojsULvTra+9x7Alo5ol9sq/xrshC2Nu+R5S1o+TadFLVm0dbfKhMaYXeCznvCkSe1ixY
bkTymM6dpVpc84hUxA5dg0SE4sd84+s5prnYAYQVeV3MTewgKlJ1x51qSweReFDk07es0Yujlvp4
JpHY8oj0vZa7Q9ISa9caSsZ4uuPNbJqAVcDPf4T4KElvK7VlgnEkwGE+sd8KQZK9oqQrJjH6RDZg
cqZmFonOKX52i2PIQrRzKaoRu7XC3ZphlVy3IAS06ggoSwh3rf1gGonUceJLMU0fw5sAxfjcOF7e
CcgIpYOoTde97D3NtNPzNXMjwfumFDgn0mBCShjungdfagEgpcm1RqQy1urIf/HWoqmAC1RXPrVk
yUuraq/TBKgmGCrB7y0iSyPGHiYmglPpY9/F+zOPTutvFI8DOlUOsyQEpfB1bNaCnutZ0WVUiVIy
GndlKcGEFHEGOZTX1I2a497NukD4fKbR87HLbIJwNJ5z8zbY8sn/+JR1tCL0ZOglXz3m6kkMPGdW
ht6OMrb83uaw7/YwUXUWse0dNyNRxj/wkAIaC8kIHz7l6pmP2zMG3D8jh3JInU0gkV+rmN6OdNRN
DSNAtxhmeFrp7NxoRmPMy46gnau3GOvac3+QNg6HcTtcSkIRns6HVzw1l7Ry+LJi3X6qCtuo3K3g
/Df7+3E40EC9+7yt+8eKKK0IjyIaocnzIqHynp0Tdsbd6btfcrIaOqh7uB01hFJuLM5+8+oaxuaO
Urn7jg72prZ4qbp2WOFrxWe1X2RlRdadrdDRb4u0JEhyumOlIStyjAFlP47Lylw+cfZu7V5DXGO2
FCD/65PiowECy+1oZLygUXg8N3d94/f1Wzy0IxgTFhLzON+RMxGHAy1eZo7fj6E1uHLBoED8qZOQ
oiS3uc2pGtaibrJU2HVMBcb/j6RZ4RON2Ut6sLixGy9DgZdBmNYU28rVAAXBWEWXjQumqzOo8APp
utQQN9S1ObXNsDSU2PGsma+lcxs+T4dxZF76/leWjpbaFdlLH24SXrMsb124dGK/Y5fhvYpY9ML0
aFTEsbVgEHYAUiADKw41kkSx0zeh5ujGsjLlBsyUdCW9J0ejB/J/tjkjsqhwzMka6ajh4TTrU1Zj
p4Na19jK+wiBl7OsmymylHjaYjyQEegKsfXMuE0RlWIMJGxQ/o64dfYYN/+eNu5k9v3yzIVefYwt
teC9zo++DRA6GyGKNt68Nl6VHi/BMCFwdcA7xdTb+8OZPBDrkmN9oKJlRPObiUWYOi46vfrle6Sm
5S71MBmLjX8ERH4HO+fkZ2tUpYoEk5v70jHNCJ4dCeieDVbS1yigKhhs+391KchVHUWfFtQN1Zra
6KIP26p6Fc8BFzj1HjPYHTdljSsRA5Fs/y9ikfKlXpgcCoQsjHUb+2jjw4uW6G/lWhaHgkxjB3y9
WerrVE9HR7KscsavMAfzLaiIOFGLgsfrCB1JRVnbmpIta2vdbZnWanpe26wiN30wRaPSSG2EGCBi
wF2p1pEJVgXlK04aF39gpVwgkLn4Vdgz1qBV/tMGFD+gdCLWnN0af6HNgCnkjOn8gQgsqIWs6cEG
LuZSyf4wV5j3dssPfLVc2r61+GKF3jTPczPTC2zExrkuSipqXn8qsM9cUhDGR+2AgUlNnRHwAsiF
uxXi9ZMkS4W1QvQxi8yo70EBF125QU/L/jVYpquiBIMNotpWss3EKTac6CKa9QVu13ajxFO/Y9kO
OLJTx9RnJBh/blhBYEi/h6T1pf9+1H2P41yPi3pWVvo3uQaKs4GnQ0f+RKe+4Hx2jShowFSZt/Ig
ebZXm18x00qGnSUq9egu2GBs7YUX7iXppC4C8bJjcLV+yMqO4sIfrSKX+BG2dJhVN1xgHgIcJ5++
Zd6a3iz4BzPwkybhww2P+JkEcpEKV55SMdtDK8zBddnQhO7hEIhxSqdaUd5MKQ4NREVK/6BqYf/6
XoMX3dRABHguVoszTE+GJxaYpLAPlpVVRN6zOO0qXPAcea1MutU4P6dr+jZ9YIKUzBlsFXodCfRJ
xYh8yLewNHIdQaXYgCfnZD6cBaG15CbPwK7goE4lamhdy91cO7DWHDfNidHfVGHMFViIejJgr9K7
GSezZ6NzuxZ0bEZa6BWeX06vLtrNXbr5IPNUYNJu5JJCtYeoTKLT0QygIMJupCLMxefpdmbWfwAh
ZFlaFBsRA9TwKKzBTGYlDbT9NnUlfI2Jv8DIfXglbqDp4dvdXl32/sk9fSHW25fY2alsWGRmDQ6M
803BS/6wojRX6untF5234EVsSGvz8PFQMz2fSXqYQoVuPiaQ63n543I4EM0kSrDhBgtWKu6P24/d
zonANfFwqbar374xxOPWZWwlaz0d4MCVhHWs/dbV0pnqMfodpEDtIt33pGe41uIIkLfPTru5KrwV
pG+sFI1L4YeSRQ7mXAy4EFZ/sDVO/cjkwn0drkcGKbkEoQp2M7pObCnRw3vO11rwJH7Aqbitz6Qx
Xw/l5IR0k4fayZPHyY4Kp9EpEyXb2GOSAN9CM/5Ck6H/RFx45VyvmMwLNGuuS0Wy8FWrA2TlM5Zo
Gxw+NftMkO4lqWlEFme663GkIjBMYueSrAKrW6FMWyti0GQwxAAVqfGfl3+NYpscRMHzAD95Iloe
TpwAOWzohRxGpAPa3TAh6eobNnUsJ9yXwJIHbvStwq+BNVKNqiisZBjwTh7NBjIvpOtSeDOEi9aA
PrSSSP1sLOmTcZwLMaRN3Ex8cj5Z7Y7aYh5KiZ0UbR1s04Eds0cbO23W0m64K774IiWau9kOKQ3N
+nTcVyW8aUtiVscdlokJx1F7u9q7mBfNdzxsHSyAUwGDTKv2v+uXyyAZbNihVE/VgyTd/wI2BVsE
oJbpVvkCMK00673pahWcU+l2FbhPddqOZH9UrePN6a4+Ey3mI+ulLKV8UiAqysaccJ6AKS8y9Hul
SEXsRhYTpSjXf9BhPOkxF900dyaKtSykkpiIZpSY0VyLFilQrgdrpDwX6eeJh/UoXswWhs3ftlWa
Mk0N7OIOWSEgdR0NzKIQlMt4wGr+WFw+uhaL+ZObfPrxnSSqWdLvvWuIxiZGe6TO948K6V51sZOk
3wQb52hf6Ktc6FJb4Pc0H6vAat2Cw4JJwGGgku/9kXP6Mnk0jPvpwy0apPgRUrE200osHQldijVZ
mugax99mDrlQwoxpsP53wEqxvW5hHwHZ5LPp/ywb8RRUtIec7w3ypDEIc6SaxySZqeX+n+dCtxJT
fyGYnx8KU57ltcRhr0NcSdux+8ah0TYB0v4vRtXWHQUr+BKHFIPGyv2MHvsRKYgpTJC4F/W6MWxM
KOA4+miJLzEmiekzY4NpRJv5sd9xFX7K8/SZYs/t6rzkZP7lbAHZBrgCO4oAFtws6Dak5fKS8mZB
QG++q4awI/Vdw0ac0m98BxeSAtPly7MmtGKaIsG93xXGBbhpRrsu1Niyrc8my0RixkbStynmtsUG
Y6TOmgzsNZYbfhpbiawXw3+F7xsmq7YDyV1fWPVtTRfzOIASlcM8UXp0dGI9lS/xNWVkKnY4NE16
dizYWQ8rf7wr8vf7Mvb2yNafubQF8zDfJeqcb0j2yDb1/nCf+eoOI3bM2dD51ePQWnJu8qHrqXa2
32/08Tc3gWxWCrPSUBeEG42hn4pc2ipQKh8y5rdjoAX7CyHbJzauTpjng/ZzYLRsIU7QU1BUsfhv
Il1fkaBB2cDba42kOzGXZBccEveW/rZpwW7VildXzTUaZjcEdZrOC4QLbZ6EqAp9fruBr4cpIiFP
SwPvea08O7z6oM2NXiBY0X7dgC4nvv3PrmgmJ8NaupxLL04XKgJ5djcfABMq2VU4HaTrZoLWD3lI
tabVeEzgUcNAaL4ZsCyzQ/IsS1HtDLKfgGUOQjIbHcmLkKQQHgot3cR/Paja7dAlCYclItCz98TM
KORBzyn3ec10WwTxrFTDAJznE656iC0VKIltS6WjeK9b2xL1N76CsD6YkJ/jBoXzP01h8A5H5Y/l
P95ffLkQpQb1W5Yy8CxTTzmB0WdFW2AmVsgRZd9CFMBgeHWhaYPgrH9Dxm/VM15XcgwWwb4dAfGb
JHTZeOWg92NKEYAU4Yy5l3GIsoMb4s/gQYofDtU3bBIxpj5MgilXcerc2l6RbdoHg/kT2X5Qjpwi
S4N7QUGX62wHpM88VpMxqy1kyw4BOR9Bvxa2BQJlxM7atI23HpseRG+qocglvF8FG0QI7eBT990v
3sJ7pa72EPZ0v+8QWq9j8Ghb3igGMyP5S/dzyMDjWSSx8GPVo/f/RvlwG2rnX2RBl00VUwO0WjI+
hHA2C1DslR7p5qAoV+cJKIGicXlBRptXbqv9+gerGk6JEppvGFo0abYjLJkQu8BdBOsINKAZiN+/
zdSgR6E3IYkfsEHdf2RvFFQk02HB7VBXN5SPIibQ8Rp3LlUnrdqDqcJ4wabi3pHOL4IJee/ZUDtk
WnB9DMrT4C3+tl+dhelip8oOm2D8NSvDW0d46wm2lDoL4fkpmZ5sbA1/AvPxrmoxwrdvECFonSxl
bhujAW6RBETTHtBFrRjOmxjLU1zWbZzONKNSgtFIOB0n3WAvCVVUxGU6L/ncg2ZyZhuAreiMQ07C
bIwPOrGPv/4Is/G6vxoms6cJ0/1HDvKcSa4yHLOrCnZSgKRNiGphgiui/ZnnrZ8vwESMTXs3Y+a7
9bz+A1XtLfPMnRaJT9WFx7fz1Xyt+yHvaKGEQdyeY8R4D06MQfXjKfI/mTs70lcUr/d3rdKmvmoW
ZYOKm2NsPKBltvHxGTme5ZACHm2CNfCnUjhTapIEISBGTayMTuTHN+lEohcnH3Rm0ysiLuWeZvcd
5s9Ccaax5ytxTFmJw7P+jEiibeL/jMcyMmq00XjQMGA1ny/tgUAGxDqje65An8YQy0fXPlC1od2q
9XGNqNMJL+WO9UH+uvshR183fW6oSRwNH9EdmrnWxez3otOy3VnDXFWI1X8hv37YPkzEinr9IhEf
P5UE02MAfZQq7LQBj4BWAiOd3PVVcBQHVw54QcK3gN1HqnC2ctG9IM6dhyXuWWJ2uxrnXFp4qAyw
qQMx6cOHAQ6CMQCvF61ZIFswKFjPAmN/4m+iQCjdzTih2mYTnUiDRK7tVYnPVxEo9j2gtzlqDLpG
tLEUeF9pP32NFbSquDJg9VZ3ctfUGfFX4zAczCrnPjYG74OerUznRNvA5U9DrTs5llqADTn90RIn
uoHL9sR6j/gIvwhF0i4YH1eBxuEgmPZJNfqHVMvQRfcMQx39kPok9ipk6Fb8dFX0TCWx1rh4mN3H
LV5xoM9eH+OtIbdzWv34RV+sF0/GJEJN/7D9ZxxiX1j9I8nN9JZlZpH9VbzLguAoZ+flbkHj5s6R
p85/sDTcbSonTsJ7WoIuJeLRh2d1O/FZ6jiFUMEBBtCFBgJs+Zrk0uzuRvHCeMpTojVOyx1PprFh
hAJCTloF9/XAQSnJwPy5746xt4DSklHAbBJaqCw/qh0j03etidsorFqCTFHsweyU+zPuX3mpfBuV
wfedeZwPFNXks2LBZbbINmF7El+VbP10a6WYr1XAR5fzl7WKfJxcVf++o3nEaeo4vx9t2A9S3bby
KHeh34vCBW8FKZn23WmBHUZN2QDacZKipnlMMdeuI8SgeIGSXs3Cft2UgAp9nPvMb0eISDrla8hF
IvcX718gGutU2fy5/GlTxIMZw2rgW3Y8R7CRIat79rx6zbi7iBdX37EWDJ8dYpyhtllpbKRzDM5P
AnxB0TsWmgIEtc9xZZFCULzQJgtP6JrVsmkUkEW8PzIvI9qOicdaqr3U7BBlDof9wbKuHgGpChxV
c33Scon+R618kebPWEwx3pRfSJC1bra0XnVp1c9ErYHliVnlKyuRN0JSYkgiRMsK/fsOsbnZ3qXi
Rfv59s0x9lV29fHTB1iMrfyvzBqg9miXl2zrOuXSF4QuiXjJpOgNw/EstNxPRbHQ2aKRM5U20JCd
ncu7okeHJovDTxjyCKzQxKr1EiSmW092aFVxpPgdIbIGh2sbfE1joCKy6HXYW/wTlGYF8IRY+4eE
0eC8c51bkxlMpg4hMgy9G5f0v2y1HTEsllf8Oq2nI8bzDHWXJb68eDlFdD2kPCF7QKt8onEHxudz
ts/41qZtR4z0ifHSKxh1OSRLZyvdGoDH8C67Nt3pI32S9j5M8M/o35azUtSe21Q59Cyx/TwNn8aS
3ldWIfx9QxfN2z0CQm8PO3BqXS5bO3Sy2vMMk+xYgC7Cjz3j8qZCNFq/hh13WXCG01ludG2Iidnk
l2+HGW4c2siu6teZYDRD6dqdGnc0ZGuRzZTK2BboGYYo/HNOj4ATNJ10BNjWskHpp63NMysBQKZM
moEto0zDY3vypuXh8wRIaE5jgORbG8JOizYyMRSbfw75NIV7zIsiW7nz5OV1nfEJ7iwb1RgcnKWn
ZuN8ELaAzUksPt3bvTSBlKBzsZjxCXmaQ8CeRV5z3nl7IUGV6NfTB5jbLA3ZBBNgVj83fVw/Via+
NutIQdR6wUUaA3z/xU/5mmPtMu9k3ThqPg/87QAa8+eMbbhqGHQRTW2mNqa4Wkt14Ydvp6/McVyP
GFMlS1YCqNZ1UWN7A2hPEWchjW5orOolC3DloFDcVbbf4117CxTFAXlh6c0MPPtNQWfwTqwCLqtM
h4LqNWk8U8uyjrCt0rbB62MxtOaCpIRREUSYICxgV2t3hzee+27fEB51qkWS1FBw7oW01FnvoEMP
iV4RSSoWiq+dFeSEu6AVXVQls37DU9mxjoQ6MeY7gvHPMdzh0jBFFwBv4zP2o/cYY+pMLa2YSGOG
Tj8CNAydZS0xmzFMexOnc6iWEwg7GNbfxPVbYqzeQFa6/N1pPtYbpy0ULpUqEjlC7YCiVbKlqESc
l9MrcSjwFa5Tt1aeb3GqO4ayC8xcfFQKxe5Z74gOEj2QOgHfAr9pVwgjblTJrmdgil/EZm8IfAXR
Po5eSZEH8BTMtIw7331wU7Y40kv1cQBeqejgj2pIHARh/7ZnMaZvNCxZ7ZC03txT74fL/SaXIZAT
b0DxkEAzpVHczNWk8Wu+p+dWqneqPQHFMVkInGbB8KDiREHFQJl9RhUyHq7DmriCVCizkRgMFDiU
UNqz1dvjJU4nCTWFGF+rLX+MuPWYIpqjf4Sx3Z7wksaDZbw35ofvw2muNVJvmAeK1RzhqQYNlj59
hdCKvrCNCaRtYGL0EJuQ3Bz8roBfjurjuWkWqqRW3UL23cajaT5Lq5rjXvat+W9s8dMakcFyL3z8
F7/x+urj04aaTALeJct4Gkw3XvM31Fw6eV6JItnqxUe9fj1CNSmqqWxYs966RfshO8V4cscAzlDR
uXCJ8+EaG7INc2KRNxx5Sx5dulU9aICMmpTkmBTE45IHIoRyD1f6JHYTHCecDz1RprkXHZ/8OvKo
tZnuIHGFJXoBtB/hef146wq1//r8TU81Xr3Krs6w6HEPJvTcpvc3CFaxtQC1nJzj8t4u/7ZlyhdA
6sP+yg8y0XVgFW6BEgoZ6Dho2UwuUyBjcLbLuNl85wBIfMRhfT4RBxj1GUwkfMVDzKJIVc6QeQ5F
a/zuGNp+kZ6qDdascRYwkw+D/52aQ0IMtw/NCAHdkr4F7HCi2NiONtUk3O51FkrEiK6epH63CXKg
lmD82p0iorX+bjq+xtS03FdoAzhBLpH9WGfIgcnVELLKATe6yKFA3ZFgHb05IlC+uXalBUQ28xzl
KcXFBRBZ6dyMJrmlJnvXFFCVhepf/4QnlMCuVJGLG8hPnhvSAMSI2rU5Y1Xmbts0rVifKv98ZCeC
OFZts4N8fz30MXQEqwpjImExOXN6Ct2X1qDAqN9d773WZgF+BsmMCUnuQuEYBdHH28fFNB0EO0SJ
B6uR28HAK87bZcrV8qJ+/GtONiQ5QwODBSEAMBsPcvMHK4A1IeZNdAZAM4o2y2rtLiaUQmFMmBUR
V9w1s+EHahCEfYt6cn8nt2GP1H5jxJLD4Ji8Vwr2ahJUK3AXDL9sMi3ipeSVNMtwWF1RXUNLWUGe
wm7siAsTXUabVfQj5Ks+cLrItCytrrbj06joyoYyMIkDMuPQQqCR2vKZeEjQ2cXEYXaI5k7oizeT
rhTmjfb3WbFK1AYItk6EjQV8J5YArtjqUt6VwvCxHrhDxRRb31vIQ6KuXmcPqxSe30T3uKg0tMc1
NioCQMEeAEV0yGo7xovJy3VxUpIEQVMezXOGU2BT3TNm+IeSV2eH4lDfEvZkO5fGoqoV+nObQnbh
nmX6AcvJUU4wd1FRFE1m22n0GWN4lnof2Vf+lo/GjD1mog4MVfXQcLo9MSKP49/MiEsq78Ya0Z55
vAoidl0GjWE5jCL9bED32pkGACS/OgEuUvrsOSJOSMALVXGFp2cbSzLVEhrAR7MCLRLveKKFJIQy
F6BJpLP8JAAfAS9BCduGWb/cnuD8gB3ZOOCLiPQLKAzI13bLrjxERgnXb8ATOmy7SvWpuAX2yRU3
SzpQ0gDi55k0NnmlX2/mbv/+jhii9DsOPoSAk3zfUxSz83uP2sRtVV/ADkWx48qoTPOJKzdU21a0
FNy36WSoS+w5qPjkq3FWcLCGisypM6h7F9NAf0QThIFvmB0UwTP1cuGlh/+DIK9vyGYVbUbcRZx/
Nma1Z2Vs0uqJmsTyJpUvAKt/WwVuI8LvVu3lwSMkpElijc0lpzfKzj2u0Y9yUtkv+5fQyAXZL1OT
PWJrJzH7BjQ2vpKH1wQH5EODtfivJKjnrKPMD5bBAJdAyq7jFoSPziTmBZG/eM5/5pRTZrTE3li3
rl+d7Zv0fOVCcIR/+OrNyphmZVLkixjRBo3FOSH1nO8t+pItuoh08rJYBqU+NP7tkoERUTqfPr5L
+H6BR2cmR31a0QnORdCdBqGN9QML1siMADrWupQozksGLih7yR7EINVUHvKE+o30C0Ukn9vu8qn2
Wc8Xr/NaLp2UXC3ykXpYAand485PiA/mlOIsowjcbAGUd2whOxOh72AAXwcFtR5Glre8Ks221Wfk
ECZSgMf9jL5qJSxrqvuHOb6MAp3JzhRGjMbqEMqxeQt2IDhdG2cLdPc77IE45ps2jNxzE/IiOgja
Bs8gU2z/Su7fzM0q7xOUWiKqwzg4+2Xo3P2789fXO4BJJ+fj9IUGyB4XCyg1qFTVcbchiQfA4u76
BKLglQlR/AnRoEzgsAsg70YSCQk1OT0Nza/t5O8x7IQtDfBB1frs0L8nMoOppAi9zZzMREO29zrg
PNQUzYgU3e75hZJ1cWoDBQxG6WSHKubDpWzqprlVyDDfSpN9k0AOV9/Z1FmWqk8+V9O3TERg9jys
nMA2ux25DpSrDGyuq08ug4K0TMehTcJqJnzfzSvdKBWsy2BDv4Yzpwa20/td/AjSpTe7l+YjZauT
7SWJ7ekklRXHZlQT36QMk1hsCwozXwPA51W4D9tddjrmtCOVZwuyVw8WCR3geL7lQBhfA81nTDXK
u1FT8Iccppb+99L1S7ZkPKsLoU5da1t//2Z6yMvt7ToQQfyr74TiljUH/92RldAI9qva61qI50+b
PedpidDd55BVr5S5oiWZ7zzcRUFUy4viSLTl+jqi6y0ZKWHNTicIHFGj0ezIboynJ+9czmXdjfix
YPGIwSSGEC6aA1BGITnviWwc+701w5F69dQbfa1hG1Qc03AoS7kPjzh/EzYBwzSyzWFL6pfHCliU
76lTf+sCuVRZHIIkQz3HpLt+NfaxxkIQ8DPgb2SulXGH1BmwtJ6ldZgbOeA9GWB9gFCnWbN/2va2
qqR1hhtjWle0tgC4cVdzeIZdBCc+Zk3m4wgdybPWmyIRsWJjca7aXvq/ZO8Ja2tTmjGo6Q/gaEMu
9Oma1ZjEkpwqjfqe+H7tvLSdtLM4rvConEVsM7oO+5AI+8qmHi1Q2B/bWFr1hH447JxEnOo9mhol
j7caEGwd0uo+bIE/2RaOJn8zq5b5xE3ItCzi/viZZIpTR+MIj7ftokcD9SM7fVDaJml/VT1TNAWg
f5x38/dGqXTWCcChcTE09Kq8tcDAKe71krWHFBnt72Sn8My5uNTJmb4CX8wMqRx6rjuS93Q7UUxi
QoltGCiGvPQ8w1CedYFPBS0cWzQdeftSwYyEvx93fx/hWdvc96GlVbjcnPVNGVG+5FLowO4KuZ8i
0Z0RhdiOPS2Tg5j0pDg9/rdKe0qG+GG+CKL+ERuo86KR6cI3gAqGC4KHc0gSe/aWfo5MQfYdraVy
rSdesc9ayynHJK4fAFeRgfpkwOHGzZR1G0VgQZ5nDeNQR8wF7GihXbrH+Mez+khCtK4u0y8/xuPE
ENAc2pIjX7wh8Bc63S/UtvG1jqj1oLF/XO3FrmL5EUFtXCUjJ1orHd0K9bBSMKMqMQ8CkOAxDeZ7
jMepvsJ0rrPJ6r8E4EyzR84gWuFLz6r8t4NKMG2/2SFMWduIcwFm2qCG0dwgXjiNMBhbtJLSJgfL
3tACwksQLgL7w3P5bR+CUl/v2OwoNL1cyd59R69DDIO5oRmYEpQuUWYC67KYWoc2nyVbSRGgjxlO
4Iy6giLVdZIVccwkF1Ti2FIWTJHakZbifM7OdYo6Yb7X4Zidia7s0Vz8kZEyOZ820GrXopONv2kl
d8K4ouvkynjpEi5n6p3hs1BtBC9NIr7f5UWuyHWegCPtP9Nr6rTRfVz0H/JKh9x0GnABHVDTD1iD
B2cvdLbJjTZAq4Jq5C0NUkg10RJyTGviKkDV8VBtA3ImD69ONRt84QpBgHx377fVwVgJuSxcK5uB
JmfNUj8oknizNnjX7/mo/h6beQM+28+Za3pgJis4/3gFXfJgOaekllPxfNnmGczaRT3iwXhMYOHo
X2+tV13IsyxlkxOKe1VjncUchv3h5hUvU4PfBcX9aewTYvsH5o0rqdxr86nLvwGKJk8xp9x4UBwH
nIQ2pb15m21dvai6nF2DrfE1V3WZ0+WWY03Ghxm/kcUk/N+RKbo9os9J4pD1/QZc3PiTk81MC6IL
kX/aOror+nlMQH19zGpi41HX/KXTlsy/9T5YY40rUoENWFFPDQvsU4Gn3GIlD/17ezNfrbNYhpt7
cNyHDzseTKw1oLJ49zZmEBeYTXf1mU8DmFsTIPgO+e73TbItbtjqFjzKGoG1X7VZLslG73WTcYhp
ECsNpLukCfW5QlgT+3K88OaIdLICltMRFDy0gv+6eAwuB1shsQbcvFlsKStitgj8sLja0PYdRSlK
EI2Pgs9s8zlWs8rHXn+K6pDXG7mQ0pXr+/muIHY9ZPHwv566bHXra18TpFI4VSypQ5x9mDXlGDuW
tF3aLWvXu9EWtnoNNImTFcHdQPR5AnqO7tcW0z2xP2j3flxih2mCVZHtye72jee11/CfaVQF4jA6
vKbWPXH5agB/ISvm1Hw+m7Ds/0HoNkbh75g1gYL8tHsDGHdLRcUhk0sO/TKV22RyWpoe0PbKRxV9
rywFF2aPF5E8LkLeTC+CZx7WlaViGE7T+a0RJbxW5lcAAaSB0nqjv5RkYh9m1gqSf1fvydjIOI4j
/2NSB+De/RwRNj6GVE1RdA4Xneusc6aXs3Sg586JluLlyRaorPuVk+aC15HNHLeY99jqsVlEBlne
cr+bsFIIwYmbZRqrtPVee0HZPpaH+nfV1GzIoALlVzhuEWV1McO0+x1OMoBTJWh8qk4pXEv2Q+C3
TG4wDhT++vTTjADAbUl9z2ESmnHoypkxp61SGhUHOLfaGmZx5Fi3y3++mrXrEzE8sG8pV7o2OS42
75uAvYZ3Yw5toqXKyvryD/D2Cn1Iy59UDfQc44LQf7gsYThE2FFv9Si5kaT9Rj7G8O2vhfAJ2DuG
JnXJvo4i68QWy1GlIuz0WDMgIM/YwZh4PLwpyEH5FgSLE7xXP9tET4CdlJ5yVrNm4POk4V5+dJTD
/P1S670s4EpEbObo8vdPXqgUZf3IrfhdnLfU7zWvdB+Oe6tuxZvJ9xx4OOSnmve+CtCNpI34omU6
jiax6SDAhEjtnnsZ2Ydt9YR83KJ6TLXPuuzsFzUmBD8483gUvnd4j6Tq2LVk0ZtcWkVnYRDBlQy4
Y8jOQ0uRsmpGkZlIrMgT3OnQDTH3DxIBtQprx654IKcOQmdwMQ1iuTxUmEhos3c7T6H919Y9hUYD
M/odO4sZQwb4nZT4BvUu1ITJW4ybj0mYlCNXMAsoey4edJuU+Oq5O7d9N22rPrCzFX7CsyS34gxy
0GxtlNsPMHFE9DofbTldhJSo2eRz1CBLlkiYhHmrX5uquvJnZZMw3H0UB9BPW1CpbIJt7GahHWDz
I6Ek9hbRysFIMJ0w2S2kjllRQNxydE/2BW8myBMQZ7MHEXRIU8oKGB1CQvsgm7/g+I2ZauCXUwLG
KP1bUSjNoJeo415JHLaFJPsyQvosANH6LpyJ+bH+En1NfVqGJJcUabZi28Rd0oxM4yNlV0wi7tjj
B54akjoq1JriPjfSC41P4f/sWEwErbAmBUARFX53CwFYgOGm20eGuw5QaNhYInBCF0dMOrgH4iPp
PHEwCVhp9DC2h0eiECYuH567H9KJxcJzZaus6BmxfjxaMC3nFFOn045CcU4RZHrqBLyx8nYPvEnl
qJWnTJpihrk7/xAIpQcrd7laKwdBQP6SUOPaeoin49ESoYleAWhrxruKM4ej5owIChIYMmH8b2d4
9TWnRCDen2eddCHwL8CzY88SJ0Q/rRObPdwCU6SmML3Q+ly+MHj0/6fGN3GgDi8l7yhx8Trdj07T
uM7mnYVVhOA8VdyFnj80GUrdOJVL0cKAIeeiSJQj9RYwu86IpYGIIPJADg9xKnBj5tK4R3nfUCWN
XAFbUvJSzl6ktBc+6y5N3yPIdDwKJs2+iYSjp/tznpr3fMMBaEr5JOzltFG/NS+XXdlKdRgjybdW
BfcVlfn3gSNKGV6l7H5yrOxokt8jmiQTCcfNOUQ9dJwxOiOQpzjsoSzt56fPeoJuuqZXfxNIvW1Q
o/G1MujJeT2h0aafwNrmjx4YrmmoKQNcvD8JDj8rE23VcmbK11HfhnG+VPg+6YcmfV7foBumZt1I
G9LU2tDhrge0nmU3ly0IbmeAcEIHsdaqe73HudM2DMtbtxiU/y7YvfVA58AD7S8Uk0J5QerUXaEd
4C7LnPZVauPXvfbpgZc6WwKGzbSpOjFS2OaomxjjoSZYEdB5UgDDmlxzEacD86X/EcidKWSHf1cR
NdpD4/FxCsPcuHRX7674Py6vGKqq3SQGNgzRT8uq9fZA5D9MTini6uY5nblEDXiZ2Yj6svCul1o6
nOVqdIe48qnF6T2/k7aOdfN3soxohecOehuf5mODyJAOTw5N8Yjb2B0UX178MajGISo45H6Da83a
L69M38mllqsu58cdx2tP386p/UeS4iE45O4cU1UHMNBoJarTnS9CsqSmXwD8lxQ877lKbnqed5G6
XRk4IETGDW5V37KOrEUeJzJyUVxMj8cKbndvKGwI/Gxpl3UrweqUIX1AobaqrhYG02Iq1KysLzMu
t1riI/JyJWcuWgnEdtpfhnnFu4eIJFulOUScQ7E6PhDLjNkFmO9IbBIWPLjmP/e3PaQfrgsGvebY
3vPJOOFxPBF6d69HTHKW7HSUZReXCfmWIg5gks86RZn+QChnBof1HHV/3dNVnkQSsGZmVim14TH5
QB/3oWV+LLKjwPk54eE9zaKd70whC9il2BvmzKnZRHmK6Jl5qLOwzpBjqPeM09tkHPrsLc9e70cq
PLa9159gUlzfilNjn/+stBzpBK2gUEAnNKH343P0U30cQT0KDdWdv8O/4bxctrRYLa1ojGDDZRNT
YBkYyA1Z8ko43U2YO6WAzSyGTUfRL02h29MjzjdDLYj7E4a/vV9m9eV3twKfu7UeJjb77OQPoij4
yrDx1Gjql3qccgmgbwda2kWPdk9cJZs259i/HMcjsyIQPmB1bzZNVaD9sAw8Ow08Gdc43+4vrA2J
BCYgSN8WxXr2n3eIig+r5JxytynbhnxIxv9NJ8S/bZ9F5Aeulr+/ZiLP4d/P7O/A6JSM7CPNyxVt
iWKxfoSYmokLqc4W7sZF3DfyfEIQku4VlmotVstV4R9L8ve1UJmwrz0edc6LSyuGfavm+c+DmXBW
mcIpHSeL3I7trngT+rlQCRVMqqmH/hldmuXBVNwIO2f8dKcAeuuDy+YCvjOfilIHkk/E5W9P5RtS
p4kXnAfLwk7Jh2TuBjSk8JuAc1eJtNxqNrpIKhl4boNClt+t9zi6KywpLv5t0pK1s7U6KUK1vbG1
zCZNypVDA5aUg8AYUKAJmeDmfyLyxDJ9SVwNRI/ca0+86nTNDAIm80kjbJocMR2GrNox0Qi/py7L
NzXbsDcU52Ex2tc3DI484HLWiA9M+/sK559Ues11of/J6nm2KQxe6o+j5VT7m4Hm7A2uy47z87jO
6C2cCz6OkrMNTIjffXlzJfvEG6DA357nYbQFf8v7xhgqNRmKAfLQJPKo8dzOnQ0/lQ9WHMLRr3GO
nd5Bi5dVAm8xFOhwuvXNcUQ3ZcdhnD1PT1Of8r3vX8qe9JGqWL5gH2oHcL1dRs5ZxZroKEgH3Ay6
ELZKYfBZpI3khWyqw+qJt4Aw+cYgBYzyHgTs4XEajavNTo8GNJhhlYsLMhw4vISmGk0oVo+Swr9Q
Qdm/kl28MepQwv+zS4lsVldLkr7SON4a7FYe+HIRa57Z7Di9CB61CjOhN02YcqR79h5QNyS+vMS1
JuXxWMdle5jF/hh22e5xaBwYIrmIUH6or4q9M+VxEKf8nZ3je8VoPIfpaNGYRiD8OVl0iF03Pk++
H0LODSFkZni+yr5CQPA2Se94rJcHkp2iFKyr+PbGeMYvSB3x0tQj3KhqoRbBzzN5VvMFrYRELGKf
B4zySmtA0kndeOCOktK/7z3WhS51OkdcTHvjZ9yaaVFCmbnsAO+T8xcLcmoCSgbgXZ8dj5FPVayQ
s3Xl2A13YJrPUU3vT7makHFLaNO4EZ8V/PrONfGBTtQfyFleAQEujD0JO6Nj9a55oX4J9Y3MtBkt
R1Btosu1O/6X3bn2wtNLao+JR8+0pbyXbq/VEsSTuxOZ5WpzU0k0aRA03Bq+HWi87igqTPV4TqpX
jcOVtWqYcUgdkE9wWT1vK7Q2hnjva5CFeWQa4MQ9s1L91Jnljc7BYz98+nLHBbv46MBw+JRcS9Xp
vLiexCUvVdS76XoJd9nTi/Ca8CQskTUD8Q9fG3ufbg+o0LtZ5zmV5M+a1f82OGTK818vAXhpUVp4
prhRcTjBh6TbImjGY0pFbS3IAw7w/TqsH6wX8FbQiJMv1jIBjjJw5a9Awkux0JbipE5TCnqjvCbV
XiTDtdN/C0owtQ9IgR+TNpJIX3oaej1zJxpAhIMx02fSu+81O7Z3SdCT8GARrD4hKnTnlaU/Yd33
syiYQcvXyn/PNBWH80gsCzjrbpdjIPjkTLrG9zRUPvyaAMIZ5Q/bVmMnvG/L23P+w5Ad24cQPIl9
KhpdFYyGB1YgSVub4e3kNEBHgkqWr3/QTQyIjBdHutY6KnNvnfgZNonVAJErTg19mDyPbPS9mz9v
cW7916ictvWxN2CK6kgrS1DGoiYUqoDMs9YJobZuY8EumfWxRieLjRrXfpZI92+seMreFcs2aUc9
npvikcIh3o8nnwBXGEvP+hUqAob08Qq3UBVVSiYy/LecDPVqxdCQOuDnlpioAV733FriNs6Y2ZJd
9y3fez4CsTi0sPmGkodOQno6zNDJB3Tl8a08HHCOjFTeRgrLMHaq/KgeonRf7LqJIo0bFRgLP7HO
Zv0vB82GDZatPM4RaLfFfzlO+NT4X+yZLL4ryxUwHhRJB5XgiHJRJaMeQQPm13e2KPIt7CYHBaqL
7X0xJmNxYCqiclvYtXFJxq9NEZgk+NyO7j/G8wAUjt626VpfBmiaoOkJPoVX2ERq7BXJrLb6s/qo
7y2R4jrXSfRDeTh8wlwTKq5DEZcHzT1beNuReytdAv5hNxFiIXGtuzSuG2qsQ50lfbKq6IRz1RQH
AXDpocv1HCTl5GAgggwhYVJ26j/BuhYrhmEeFEJO0AFnhvV1F6CefbO1beC6Mcv/WkLaC4v5IpJW
hgnJEyxDt0eTN3jlBZKKKMfS3mrvNXReGMAanCP4D506Eo7DWSJd6f99YQpOn30YN/ikUdzns1sK
qn4YZ00SP/W8YfaPfweYhk5nQbqjiqsG4TQxBbpdAkC2HRFJLe1Q1PGG6z2VrJZynmP9aav3M3D1
5CompsZrn7/JJvnUhhqFRb87uPeaXO0Gv10WNpIrkcegtOjhN7jbTw3qJkM5W1TBIyQ6UW+UJcl2
whMPEOCYAcny5VQysEWSJORLvX8iURXObxhgDkDfH6Eze3Uhw05i0chcFYuOzboM6Z83XiOp62sv
1W0UlfEsiMTSXdA9fZVituIeK2amNh+Ms/lsEOC9k1ye52UoY1hmuOF8Sy2t6u7WubukviQh+aZW
Rrz6Y20nEB4pDix2rXVbx6XcAhZD8faudeYHo9JsO+woQ+2eao6QlpWS0n3Hr8+2tAJkC8hilt+k
EQyvpERPg7jprlNmRrqdFy6XVniI2q6VECosEGKbfVwX3aFL9QUWONS+pgCqg/03izrSGx/Nb9rU
8FSDvzLl7wqO46+MnK0fMSj4YZjPTF0/P7DIpJAp8KsjlDvF4wn58Hk55VFxKv42CBM0FfZjzY16
BEVeZsOlOD/PB3XsGB1AOtz7c2x9ThgkkwbHYvk8F9fBFFDORo3skjPdReUVzyffxo2I70bwJmk8
dW00B8azdVGu4f0rcDjD8uH7DKrexam3hPPN01fufWQb97M1cLy0wPXpiaKR+zA4cFQUC5PE+oRQ
pjmaiM6iizmYrD0fqLXICbryziS5rVp2CushS+ghDRmbJM5z4T7/Q4a6reQB+iRbBNEB4NaGmZTm
9KgzuGA+67WdTdZEku3NNyxfbRS5ONTW83DnQo1A70WXvO4W/iG8MSn71Glng2QlMMOEmWBvlWCu
TFwzM5DWiChei9G26007lAeA6OqVY5zQe6EDCiO7gcYRz1jSe2dvfmcbqvEEpwrS7bUCXsIY4CyP
IeKw4g9zuNDcScB+yV1qVW2AKPyxbzXDPzWXE7oJbQJ5Z86Fyox7z9qk/UthV8Y2/xvY/ucZxN0+
TYMaRsNy3eUDjtlTdZHR0wqx1duSD5Vxehr6LrJYZl6im775lQ8v/n9ZtXCQd0eTjJepLGVlraAH
3MxbBv51O0u9kKvF1nOuMoaoWzDlmpCqgF0xxcugWFOJP7coxBtWJqhx4GEiVUgKHhJeuIfP15Ew
tsrc6s737ESHBphNX+QJ1CDsk2P9VaesfiHHhA2AQKkPSAmmkylfAGgAeM3JpLzb/2W2b0aenw4I
xqYf9ftE0crigIbUFzCU5TSgjBYwcAsr6vv1ZxKDHLBPCmz9J4tLu6HcxDsf8oEl7Tn26Dnz9jpA
xJPy81LQKguLIDBz/jfp5QxeUnwobK389s4LBu5Ujg1QxN8lYw59V7i/AXr8RS/lM1Sa9l/13qhv
GgRSguRfUo4KQ3fFcLqS9DtBaBo9vI5/Tx2/krgZgnxXS3hGPz2v58TqRyIwWPLiAeU1Qe7+c5Eu
H6oiZEnc1/CLdR/VsomOzClUckG4NY9aQsHsQQAMoSHTjkfoiG9UqBuIP6SHRYoCSEs8y+g8DLN7
MwvGhXNNNC3w0ZCyhP/igmE11KFAkvvqkA1Frrb12ceVGVm4WgsUmUbTKXXoCiRFoqgf9yTXZn2t
2KS/rNJk5G0rSGRE/i18bXG9N6xJa1UvWel34BM2+crcEENM1SSzU91wv4Sa8E3HTdDE3JNym4ds
/EA4OYeQ8aoORsr/piP9ZLFw1nGVR7cBu123abJffvqWrYCutlsjCVnWbMyhhiI1APZC+v7hk/uW
ErBbsbCFNyoEu0w87cXkE3yu+L+PnIebKTTLBTWublWfXBOMtOqixtMUSGv26y/5bsk+FIVVR2Vp
ku1v0nKjCQ7bVtMgLmmQv1wfhRlhLuEumhJGJK30JaRo+dkTE8RgzI6TnIlzbUL1d5kXgDfSOF22
y67gvcq5rbkWjS5PGzLpV3pKcG1RKBHU+Pr4YhNSE5hyIqqoO7Y08EbNeYgxIzFAQVyOI9cKoS2O
xI0jVfmq5yqFsgQFZtytSwiKhbpKi3MCybyI/H/sGIncSK7rmiAHECA70RuS2zXk9tltvI4h4UKp
WVe2jDhFDT5AqFyxESEc+6aIS7nsY/Mox/NqKKFc7DC9Nf28q5+H/uWE3K1MLCepj9xpWsoUnSx6
kKmu8sMOEseukpHsZCzGSgyrhqxYjN2fv5yUqL90xbIi/rCZ26b2FzLXRtCbNudQ6uDgAtZq6Voc
pFDUn4+6iAcB0bEJSgk1mFtEJHyTpXcDd10X+ho6NlqsUVt9addnDrhsGS+twtsbibSP2G6QGOYA
1huTIFgAodoL6hURF0XxVngy2ygobPoZcuR1gp1Eq08yr4v1zhOAOGCariNnW79HLP7Iy2RcK63Z
A1K4skwNhCnozAItIzRPihZn/BM/OGFYMNqaq00cIq4Z2cgAxS65tjL6IYCqWxhsxNvtdUPPcxtl
4vWCjZPrX1/EFOWhFaTrxze10X/DLs+45q1247vWdNgVpV2/Len8RpUad33GoRqp5A2JppG7pjWS
TEtaG52pn1EbWeFeNX9iiqFxRnSwyNTqEWGBNsTJ5y1U+RLqpGqSe9U/AZYSIfKA2BX3x6a+GmkW
JaUjBHdw9VcrWEn8gFQOaDzgNazU7t4NCe+jHUB6RH46L06OZ4wVDrUuYnpuy2s6YaV4Adi6kncu
GHO8/a8nvrjM/KWCfQi1mRnQtNQW8ihM0ATtOXLv652b9PuqTgCBwR4cOD/NS+Nk6b39tUM5uWGq
9WVjmlvHRssnaUzeIk0sV935MAdp72VzgmJOWM75gMjfZGbDc0YNwSfnnT8mPLHKASx+P/ueFcfP
Wc0glXI3e4LtSxsJoFWrRtpcNDAZ0Jfs5CxFtzVTBxDmCYWClNRs+WAWWa5H0amFex6DzoIiRxne
c96ZvE83rU9Cq7vJ/6Gd3r/QVsx7Ag4B9hANOz8SASxwq/whhFgGc6qfecDUcdzECLRI/573k1tx
Xw57gYO3H4kVauL/GwRZkCOhXcT06/sDqtPak4jND80OQ0O3vObYu6EWF1sLSlIh14TYiM4hGrMk
FwZoD4njAhDWS5yQKO8Vgw1sBwuD1HQpv2cGLRIaFRrzh96c+BYdqbRoEUFngPd95HvitxCllxd2
LrhOYcR1bvI9kmKZeRTLIWcKQg/t2zDWpRPSGLdJBp09rrZphzpDQsEzI22ls+bePy2qgLdePkRi
NwbFFW+CN+3W91zmHyOjNkpAWB8rwtLmIV+IxBfehhAJIJMZVkEh1JvaYeHj6DU/Gwu3GdjjFBJq
niK9u1S3bSrwPMtmvLV5DNyO2NrA+vCdsqUr1B1Ob5kGaug9GikJZx2ALfpDmX4oPPbl552gufWD
69P+i2LJd+wyjU8thYaTmGPmDzWZ/SgvMTCw93n7ZjtUcgXQ/a6dASrGDufLSEf8DGEysV5+7bdc
QXS0pRREdq3r+cfQSBwW4DJ5PpmnM88xRX4+nmsf0aZLggpejhEE1YVsCh3fWWMX0L4TUDgQ3zaF
wP/EF/poT+Y1Dg3x6aW4AMphnc4GFgXJrBZwFHesRprztMLxmnqF4y6XjxdkBXv3uuUMKHVKD/W9
oDW3Lagw3L2H+zTjd7jOCjOezDn1PkTlLMjNetpMN6Hp7AxJGM359IegC9n6jG3wD+tNcoa//uSA
it81Ey9qMxKgPYdh7lOAHW7GtfNc2r3vFnLjF2qMvQVcJxppb8w80XfPP7kgLgi4UeI6mU+tCo+n
bfrZoiqArCvyZkeoTTgmJ1M9GvNp6RuNFGPFIXoJHIWAv8o6iBtgfPL516dgsltbZKW1ZFvFN8XO
X0SVbCjj7ue0j802eVaW0yWNee3vhhU7SqC3uMnc4EevMiKiBQf+BiUJjYrA3fluPfY5QnKUEeA6
XqPc1m9fvtK/sDD6EkTfc5PLnvoWmZMiehM7aBAHtrx+W7anNpYj7Jh+3iU+E7l+rAMwE7O7faE8
JQCG07a0Np3u0HSzOj5Eq2zq7NdAe5GGCcksvNAvEyauxRHEQF6zsiT+mmaJ1OW1QVMsCMlsgpnk
ipP5ZE4unWua146Em/Jf8yt3vquvtq1mjTrPNyMneXEX/U7+UgX7U0FsG8qXrze5vPk51Mg0eynf
3SV6+2ktcG6Wqg+6utc4oX81L6oZbfsr8BsGJOMY5DRrBag6Bjdsww1m9xEoALPaXc/IQ/Klo/NA
jbqMDTljDI0Ydf1mk1+4+3jmHFNEsdf4+2T6sSTTNtUcuXT2zFLnyk0bT/JEFCDAL/rtTuqcsYAG
gHigh60wRQaikyOiosZmEvJvBnlALZDJqxVQRHskdCcjVhDMrjA9RoTaFAvgpAHy+b7WafGi8MV+
j/syiZXRBzqKXYl/EbLAR1wfngDIqZCKlyodgob0QO+JM+RLL4u99mNl6guK9XSaxizqdy0IxvaU
jW8QxcdxrEW+3bGwGrE0te0YF9SsCTET0PyfU6LkBEszxJ6MUpM0wz5Ff0aS1UOL0dKETH7S3sGw
2RTkIfLkOotzYQctTQKTUvLD7KX+1EsYgzDwjId3GS5pQiN6x7bu2WvE8PduMw9KWw7O67LoS8LU
LCHRWjXyB8cnL3us9KV0Lpf6j30pPCv3NGZo3UsewfndmZ3M6wJoHYPFFYOZKHASM2XwnRIAQlRu
Jw2h6bEVx6FC8COAAj6a0f5jH1Aq73/WOeG3bksAspZGoUAMed938ulbM3asvHxZHN0XW7sNLrd3
SjLyzOD0/rPrg7SXtpSKv9Prrloiy+NxCKFYA0mvGTsbz40mkXgHj56/c1bSJyFgqPOAb8hoYfui
19b+yCdVylotPrgz0rqftZObHL7/3avFEojG/mraryGpHVBIzhEtA2Bo6RJeF+oCdZ6ennzKYE4k
GmJZDJ+jpaR47ZTQ8O3ef0HkvqFpQeec9vsf5UgET4gA0a4xR9OeqRHCON0zrnJ4jE3npJhKxrEL
whChWZXXs2910SDbrFE9B9+Q62ycNqIhYwPH6t4hg2JUyvIWXUrUhHSzbeY7ooMiSzi0nA98uhXE
+PCnsrbCK/XNcXOhecKrJQ9pjwJpDkMsu5yPGhkzwUn/1sXTkqbJ38xdp7MzOvOWyDDXPo180PI8
cSX81SH3EusxcLfunIFGfBg4boOsZuXVx5PPCFdIE1MZv8W+Mj3wrMkm27zOypI4TpHaziUjxFBq
alX3ClJExK1ijABAzXYU9YCNdd+c8mImLna4JD4mPvxMo58RnVEUW6EpTdfLzyggebf/lgWwt0HP
U7xbB4NH7xCXQxSpojOX8RokG+OCfAnhSbVL5PG3bwc8DFa957+mmkCcGV7wA9Hu8lb5m7fm265L
21gGHGbCNgDjwDyuhA0/Cqe55AdqrTC25XmGlUr7wpORYAni03yPN7VShvqKzxrEPZWc5TbqZ+sJ
1NZnnJmYTEyM3G0FMoiDBqkKaPN0Lk0tlFVez1FOxKnlsTPvEDrPXeKkhlaXCWaRL4kiF1STfdag
RmqhviwgyEKmAKN6hKFdkGNJbuji9nmXN1J1ofT44/eABoVX0Gl8liQrrtFC1sxKgUy9ANX1h1qI
RInNhlIgwrJOwuMY6nRYpyrfZgUcyBu0T1kYP9XPdxNv8Cw8kJBOjn0nKcnMIAsHKxwzcgtn1nJn
E7w9U14LPp3UV4OHa4KfhvPwTY56dybUa7m9ABYk1CzZ8pRDNNJl9hMFaETPn2gPf6QTp8ckQ7lx
3ctjPSnUDEAEV1IuE9hBbKcUhZeQ0s5EdraYptKGyoDoywOQqp7F0ILdiebQHljX0u1Xju6vrdLO
sk9STT6sXot+CpUQXz5Kjg9VWGW3YZ+ivTJELJnJRvpl7qs4UVaTjrPtSr/7f5V78qFOQkUk3dLa
azVHgRfDy3+B5Mge9An91Tx60el1xQSBw67f/OqhW+hG7UWCoEETEpHF3SxDvrqjrLMxcslTw9Oq
czzyFaF7V8q00U4eUhPu1oSKiR22L00XVyDgKlM0Vq46SCK7K2rrN/19kxzjyb2RqSPkGhlNq+Es
Vnx4W10LQHs0XjMwCm2j1Lo/CcZtGCtbkO8exHLcUGoISCjAWZPZQEsH9dKEx3dZW0vDzIRvzXyv
C5SCWFSfmi0CtRyNgyyBYE2d94Si5+SKfzeszlZMy3pN79NICdSDDzs+X9yAF/a3H4vjPK/vbBm/
p+T2iMcsSSIc7yD6ffgJQDqnK8VowiFug08utUoh4hGc31Liyzrt0fKE8hS7EELnpYdoZ2SCgeZ9
29ZfMEQ2yDTHeO5JOrEO4VZw5MOL85j9AsHNgTty4sgjuVFoF8V1FDGw7LkmMnE7TTzu3GLHG0bv
zo1y8f6als+0ZuokA0PP90lKcswXf8Hfbnlv8G2HqqQCNFGI1P1WPrkqxlGXHU3nWc4RjbrizJoz
5OHc+2TzIivddsXtt6ldPY+haTB7wP+EhxyX17XVqw339H4lUaXG80qz6ZAxe65IEZrbYELczzeO
UkLOyeoOxXKSAGMN1IpqqfBdFfj2QghbaHFfNryr2PF5wCAGFXqqDUUwMt7zRY9oC4yaPEnPglrC
NwPg2Qb2O2X9/96aURcDmD4OnVqq97yKYiLcEVZmMkspix0rMKLF/HtS3ijhRwVVYfK0cz8ZDDhd
Zf0PkHo6hUzMh92IFn8AcBJ+ouWxiv/bkEqYtz+V/RRuxFuv/xC/wIUfvweaYAHoRnxGzkDDOB8L
3kKhJKGLqa20XX3j+zmFa+Z8ifj4fl8BZcUFmkXZ3IhL3PgcO6sU48Fc/6H3My3cJYLU5uOzJSch
dBENpyDbPsWnX1vQBvkk4DG6z6hE/EvlZ8wNx2guMoBXyobDa3aI/ogZS9DTVGP3gfOTP1keprN7
Zixy/r7CXbxUKLqD9kHi0Twp5IR5T2S2xZD+cea94qxny1d5/nPdugE37GGJeU5vxUbcPZRaqiCa
LIwPFRfBmddmsQB3M8o5Xg+v41gpLFq70n9ipN+j4QvDTZwNKHZqbxAj0n/qEx0Jse/x9p2mnhrz
QXRPQTCDDmOlgtqlSFIs5+SpXD4SUKyBgO0CuElCrDrcJZcQ2lYgKzVwQGBZbL1J8jeDkrwFMnfW
I/Y3E0A4ef+O1bLAuTmpE7vukCN5GoDGqejgk/aoyx1ohgh7C+NGKw81fp/uVE4QeMD9btJJSgNw
twHlGgwx1y5M7pxdbz6SH6xgVKUfiGcqqBt2pSZvU9xS9c8hrvXD2Rs6q4fWIzVsDBdnP7ZKN1M9
/V/cpLXAnLFEpAPcueEZSa3HiOesYm/OQWSZh9/3k9tNoMYli7+A/xHi7JnuseFk52p2LK8YQy45
AyWjSLAyqzkjKOVbSV1T10/eSNRnfNwA9GeOp+M3nCXJ4l99UE/Qux9i3kvY9TbA/dizrW6lmlc0
C64W9NEyDP8DSGzrQBgag1ZXbnxbP5JqfvHn50LAKXCqnX9fw0RPtdBWM8BXkmzOfkujmg1+gDEt
hgxmRsv8CBvJaiCPGeyIWD1Fm5jRxlRGMQvmgd9t4BTMNxlV6X+7yE2YyoI57slvIH/n7YyVQMFg
UAtC6vhzEtiweJvXhq7XA8RzuzZqaEhg1wnnSS9vaA7bvObfEO/FS+JoPVv+I1lE+kQPIOiG9KD4
nQUzw8BWTxpIePFy+uoAzvDXhePF9fOgwz8Rkywr2j2yq71mCkeBohrbz77qLrq1h1s+GEyASrIH
UeMbe5dRaixrKfO3o1vgY6f3c+BDMUEqOO5XC1xqOErUqN8G90ia6zk11JkaYb9Ol9bmwVnLiCn0
l2pmGanbiR7Cu4MvIiijay2/WrB3EBZGiRflY+lAS8t41PnYg/ZO8iK7/oYNaTyRr2fDRrHRRrsW
y6eyBBBEzB4WrWCOETgcSBkBBM8FXhcI/P9jzx6eKPukqomxnLXGZl+LFSVFdGjoxQzX0A6BKEpj
69XvxxagWPAaG1ioIw1oVqQL3XGvtkgdGpoffLrggpyY4fJbKmpp6xHUlPJQThTGxrmYdLTSFRg4
xC4hqaVrY0qZVWs/qKac6p9+gQX1lIxs3PWpilxB1ouOs3oahNv3mNVIfO/zXma9J1fUWyjLwZeJ
vOL/AaE5hgdDH89NQyE7UAXngKE/XO5rhPyDXn8awQpcRoAaKe8ek2YjIFMq7knL5W1AZ7hIVMna
wDQZBWdydg+dDFR1lFu6jfDe1hPz+w1vAnCahAQqzcEJYYlbfhzM1YCRqdzQRByK4AXgVTPMlRE5
Aj/PAVw2DGwfo8ag6ozFqp2Sq4V0kbUHvKKx/DAAJZTHxhxMkzwNzv9iBtYMCm2gj2w3AdeYEJsV
MFdbyjgsHKo3ggqt0eGUcXNaSamV4pZezNsWnOVugJAdTzatDFRRTc0eeRG6hvYe5jM3ABNGan5v
GH4jZDFBQ5xPKMLrh5YaLy+M3DD3pNFr/2LYbLyJxFu19ynP58/gzqjMnRZDgOa4NdOY2bk3le53
pOy3oLFrOYCOOw7cQCMm9iX63HGjbUehfVLVNucZAkBDXoe0wvMkL2dBAtWcwomJmEm1lB1nIHEg
ZWI3wGDC773sgUFM0ljbqhmYckZVh0b5JZzApZgHAQQWVuvYYeFNWzfiMJYuxZJpXaOFJbU7zTRx
ch/8kzDqUl/I4JaT/c9gcdNjNjEIB2mgbDvgyQiJeM70FHb9VfB39eJ9/QRVRfVlQB1jTiqrRqE+
lEGmmK88JddbY1Cr76EArgSLhYObH9SOjpGSmFBqyIsAmF1Tcs8IpqAzPXavG5+KaTQFkdv4lGQM
0Vi3EkOYmyhzvVNyfTPzpAErByl7fbWw8u5hofltGnvV7FodhcSonyjdwIPf1cjwYY4dCPuQ+P6S
qEtfTz7g2Rcglpno/7vRK4VJ7xOVuMx4saOmxJWmtj0QTYkqkzroOptbIPl/uBeOy7F2VpqquKyE
cS+/QP6x6Ny8fEnkFCtl2tanJYZJYEA+M+7/27xqYxhKLk4tcAzLdO9NgKqiRKOAJGoVE+sWPoF+
wlPi3BOA7Et5S1dqO+bZBAPQK+WXsp9n40GwYkWgQthc/5QfCo2FmKbLkuTS4fRdQFheq5ljWUVb
frQ+A4cfTiamwv/VNKv8yShGkBRM4XTH8lM2KE8aiW/enG1RQI5GUkJJ8dg3NP6FzZXXLDy3mXLD
Nvy3DbjRpwfpjmBUz8xWz3DBvMhiVZeNQHlUC7W7w+gJHChVbX7MXbhw2jEZsJRbGj8bhmJWvcXf
3djzPo47fDiwDItLEAqdH7byfQJ8MTieCRwhU/mmHRqFTFQnw41kBH2725FBL95O5pryG5P0lJ6B
cm9y7zZvSvCCMknEt5tciru7mISKP0ussCQlVitDFwJQJ8yfkiKWIrRSHQ3VDsElkxTBYwKPQHKq
qZZFqidincPN/+oGtPbt2B0ILnACBrDctf0q8uN3Y/kuiSnqQgQMIWoMj8m6AJIcIkeB9caEku48
n2TyQdv6S8aLkRJ4Ki9kaI8VPkt5gtNa5HzT+FqueTw57ugmoRv1HTrrbHhhh3h37fywpKBmAe+X
QH7u3l0tcpUsPymFZ4SMith0W6+labvWBwz0ltPpaZOqn9BqJsxHhIwdiLb5YCpEO23ivuTRt0J6
WfIZuannGyf1fj3ms1IADhloeD9i/DfgsnQ7EHJgeYV2el41M8w13wJC0i3RxAUSEqcBBuwI1kPw
nGH3M7qfQziT3lEEocCw7+OWKgWc9NAkU2auYpkGYb5RKIM3yHae65hBkmHPWLXIYJud+L7fNoCE
ON11sMOXZm83MykeTMl/GKQmwBl8a6l34oMNekksPOPgO/E7PrAsFqtKSSaRQK8Yq4m7WBK4nTWV
vDH43LD4/tzcbpFTSMVvxyxrpPTPJttZZbjssq5pYanLHk7k4f1O4Z/0NmQx5kpwINXPXiz+QGfK
dkrM0bv+/N81Mazuun66NUcy5LWQfc4KY6pX2MVyL409mOi+2wkYxzRHHeGKI6kxcycCer5tLI1n
REQPxg6wQpAxBSwUtcXVD1bt8ReYMoZ92BLPTE27FYncL7CySnOuSUyIKwd8pwqt9tAJEWJh0q7d
u0PmpHRIgXi6/BP8bAK4LbD+QKmyIkpVaU5gWnio640j5SRt8N1tKbYAac/S/YSDK1GP7Qrj7DAR
SKz5ppPWSh1VcB9DUy0Sr/0n7LRBa1pzWdkLhcyqha0cfw97iSK70KOFi9j0ea0YjziiWIKvjD8g
6daZnELXVYOO4bpSAunylJ+f/LUMvmFo3PJ3Eaxdp9Tbh4bjZc9YzEPQ1oC0fSCB4IPlLs0Gaer6
4fF+04deHM2e6nZwwXAwUlP8lMEjSorbCxAOmg3klTzHoViWzuh+6cq8CUW0fMwq7Rq9d6uwT00j
XCrwzXGcoqKD88+f6Lw/+uCTfOly7aWXxBIUWJXkQNm+Rwyoy8JZzKVmxbhQIcIKgK89KyiidwIm
Lo4IPZ8WLHL/TFGOqbBRuf57QxqkaXZov0Q1QcmuGMyNYtAO9E6V99AJ1mm7CFbNCv4RuftTNPsb
OAm3REZkHV11c7cRnizC0lFMFmDDfblRwJkCOqFTI5tgb4UBKnUUVfhQLc9R59T7LTElcCY3en5L
MzJilIKS2VaxLY3T3jMV0uNnjgYDZHdUlH6yEK7IT1wHoC2xwQ6Wn4xuDzN+j6H9WsdyI5oKqq5c
R/1Kix0tOBZZEsDDXh1jK1RleujRLZxRmZXFnUmz1BMJ74fpBZ2+fRnmAdrR8e02BE02bWfLhrZr
KhGexVQYRW3AopLgjHMmAv6V8AC2ZDLUul3LkZddyqpo/7gvOriYvSGUaqg0SAN0K1AtAaXZI8W5
jLTc4qtUcvxJEyweKdhHFTOVRO9myApQFI2lk9Rb/4uI0tQa+Qlu3FDxRv7ktTPOzv/YqkNjPJCa
PzEQlGBoe4yx8gK4vwDowXYhYckVMpRcWGPWlC3bNYOgHhpFSXDfxeXmSfVeOWJOIFiwEDbFllHe
KjPqAlZBiZEHSHvfPZMUqpf26BfgdbveJXf/dUbi0C8LYitgaJiK2AmH6nAPMKOG/lQ+jrOHg68e
ckKg7v9jvVx27ZagLMr/RSLqrHo9xJr0OfIdkp2xuxmFE+VuE8kjotDtCd2wcodtmPqzc5NI7ha4
SPZT648OXn8suLNhp5qx2VQXGf6urGVGtMF6bjFaNezBmbOU5nmzdWWMfZAUG2dondsxtHx6W5iN
mypRT8+owItujjJJiIS6x8ZnHN6lNDH6deX+DG9wLVel1JiQZHtkeoVJnTS0lvHMnHEOY36UENZ3
gOStqbdhILP1mUX7737Sn+Dkq3SVMKxBQs06HMJAKzfCVHCDWnx9skaxTQv2lBKnaSHjDZVepPv/
e7j6Elacbj0uSUMcRHeHr3CL9EVWnu1hkByvVnaVkGqBAPn7XIQ8KzW5fbJqC4p2j85RifBDHPVu
jIELHQ7HHgcHW+CCzhsXQEqnL/i3N07Odza/8tmHlae49cq4WvSEluHnYoMVuzRRaXAJIOEtlgyG
daN4f0vMDfBBCNst9MaW3eMTpRrj0JcikBKrkWKOr4ba5i6Iclk6ywnO/mOPh4PfC2OIz/9RO3yk
7tAlFb9yk/bXYKUyv66gl0JpA1ADsMW6AJBfYsdiysf7t5o6W8wX8dJaVuGOc8ZB347X0JifADHg
oMuuk5aGp+Tdsmkr+qyI6qiCuPrtiJMeJRVoZ9HrSKk55y87OLNgt4DW2+ddLID9SmJ0r3n4hB8a
DJXWM3oarLmi4p4uVQTCXQbmfZB1hnMQEQdM1PSuDETDLTTDy5JMjA4Rc3V1Zo4+7W4paENdPqhz
NsNkYfLrDtZ7vj2OSueMYKcBcSdDxXsTAUuxdYSXENCcjUtshEUh8fxKCmW42vENCqpGP/DsxZL8
XuJzaVMxhH1PNZPF8dQu6HLgFkujI9ohh6L+QaIHt0Z6k3NACTeboqk3h8TYMrLrEta4uO5avD46
It3p5uwvT4Xg2a56Tn2urm+14EXDjJVtEmQMdQQnPKpk9pXA4o8AgqMCmS1LOjEEH+D2SiBSeSkA
I7pN1Dbqxjp3/Ac3XJQKwl8+It+kp7Teu2OYpZ/izZodCgXjgN0eX5G0hXf5n5rAitC4zscTyS2C
Y9J4fUZ0+wPR29XAVt17VzViTGUHSMnsgAwbId8GSf9cg0BDpFg6ErW74SVxseedZtRXkbSWS7LP
a8QG7Gl2Xkzf25+jt9SMW248PCSFwFZyMfoz//sX0ejyf+1DvMO7puT/71PudLTkXY9fXdzQQRqu
eOFUvh7VbzusD27HzMmaWoXvejtfsBQTcxCcEaRl32AAWi+aKuh9L7OBMDANG8hfAINzrHJdWqP0
wYurPP4HCADrvJF5EoHzdomHJgrx1mriM61/jOxWNbrQUuOqNOqvuioqgWjh4EyaXRcl421A82JJ
QPzEpJAoIRChEOuP+yaDohpa5kHILERsYHXCWx4dtiy/7tWzscRK6Xeo2+RqiVnxv+Fc6hX+nTPQ
LaduiY1iCly9b7ZNlHRlifxixY0UkuZM1RB3v6C31rFRvDl+egXavfjUtC9b8ngX60W++Ob0cW/x
EYI1jXXtxIQ5eMBwFUhXmstsRnooiNc6h7N+xiru7CWO19cYEMol9BWw4Q0EFheDo+OlIsTTfpY2
wBXBY0DPR+07rjE6S3aKO7XKH3TBM31OjHXSzRnPOOJ3KCYjKNttZdBLKfBOs208IDLgsqPKp5xr
8TAl4LMva1Gm/v3q6UYLbXRJPfC+12NooEh79bmJ4wurWQ7beuI/Frh4At7fmJ6Yz9ms3W+7JtWy
ZICcT2+lXvu+k/Qw+F9oWifM+pF+pAV8hEWCwPbG6B8RVxMKK2HLm/swpcOUgrlFau4Nyc1Oigyj
Hod+yTRAUnhaor80Ca+AEp5/t9R7lNlb+0BWtoda90REGYOPfaSEVphmlzgGqyPSVV0VJ0H2iG4w
yEQXj5g6n9Ob0mdOcPKL9HZhAarEXk3kgyaC83ALhWj4Og0Jmo6bGhkZRsn6mA/R1/L9G0I+AhH+
Ps741A6DDPRnVzSYnQKSp/CTaN93RJgGwXS6zk+ttI1fswibWHXgXvF4G1NKaHEt/bYBV8pd471L
PgogYUCP+HmhXOBLdgeWmvQMQu9WlEhI/Kj8YXggGMkJ7PF7NNhK4fugr2ET7qD8InKQoUSrxWt8
P4jLesGUa+W84Jd4sO3IHH0MVnAxzNOMrAqH5g28jPgNrE/nbOd4KDwXVag6OmdzCoLcy5YouSZb
2ZSY5d4AqRGtHOq3+RJ8fOd2oeY6Nh7uO50Hq2cdabD8NwpBAtPKIdUIhBcFVyE++TICmgecLhC4
1wpM4c+mqUv6QgjWmn7BbuHgHe68dzvhM95J6CD5pOphcBbnB8nUsGg7S7lycaV1GXbqo5wIlNtz
AaCvok3GeQHkCravvARxBQqbIVEAm/vT200FPD4+9a3n4s/FiOFUExljHUPg07DNo/59tXADsMF3
mzzh/QIA8KqI/jLE+cr7cJAtlg/vkUFioBVTfHjnZpbuVhaKXVW6QdpdQLnn3xBsc3Vj/7GOIojg
kOrNSFdmYIICPhdk39xUioo+VcTe3iXxvoSZEYbBVishtVjuHKHp3UwxsUX2jpb1R0UHOe5A1Hqn
iC7KQsBe+rDdP8mvYADIOkqzn5pChfakRpf3XOLH3jwaJr0AtWgqQIez8RtDhPdazVmjQAWRrEY5
VkznKmT6DkfTHf9am4Y6Kk85YHl9e2ccXG1cOwJz0YFkRwTFrx5UbawT316wWu9EqxS0GpdE1Ew8
pXlUAlONmnh+tINhE1j5sCx9dZ3eOU73yK53H9SGTS57e39e55FdQfwigSQWr5MtPYWGvKbMWeTb
wz0crAqo1qFN+PVRsqDkS6hsAWvF9tZIXkWvnIVANE4hKRY2ND0uQ2ZjRGlwF5vXI2ujiMIQ8asy
ivd0AnAcTgAS75liRLF1zZYwO8Np81ZEjkxkv54a5NM8kfp4pLGFa0Bl0d3oJO9FZEWASNCNw846
HhIw7ZEed5moVBnPz02HPgF0Uogf71+MdJ5voLjQw2HkyweArlJmR78Pdb/5WtHYYvWNuMSYLdqs
6Cre1aAoYPC0esNBpv18Jb3H38/gyQAbm9QD2YXdSFhkUVoHHRS9om+r9uGeNwJWRJ120JumdCcd
M7GqP4qC6+Obyq0JeMMRaVdsU2T7EBCAb/kS4amm3pex7QLVaCHfz9Rv0CYG+mzCkfYabNWoOkaS
+mmwgynXIKy+M1JQxPhmGLTlQ5phx8K4e4IgfiIca4ZYooTonCinSYUrGC9ovPOR2IESZrEldA5m
FeceI6PP/1uhJG+zljMJ+fp00kGJZhN0mDy0ESuPfwIN+L1IxVlXHz4L4fX5ysNJUz4FVWUhvUSz
LKv5Rl3EL0DTSsVoNv4oUwtgmt7E+VjIht8A1mn4kXeZqGQGajFhEo8f3TbNWCQLnrmR/fqnEXZg
8eCLuSZH68oAHS/EHBwsHCuleIlspn4d2F28q+YSzwOMVdxiQKBhCdLyl9pMIm97/KnhLf4UwvlT
8u51QdHd3qaYRPf2eMMpaiMWdXRqf0uRgCjZZpwzyTojmXQvfsT9mVTq7DEHKMnm4IAk266J/ZBW
sF1Llx1Ao4mMPMPARe76CxaAXh5eGH41wX0GBKofMDp2RhZ5Qx27zBJMsMITkaf5E2kEpxuTlISZ
n7iHjSfaqc1LlR+hs/+0ApXauHNQ9PlS5P/2mDx2ZUAcJJClWAT0EMqVEWgto3P3xrleqx3PJMCA
z+iSva6p7JiFRU26fZwgapsvCfYkBi8ntZQp8YDeCMd3EyXoaoSLg+MS8r3NEoS6LFBmCBJc8KGz
FwkCmjGZJDeKO6F89r/GHLic9yVaW7W6M0/s8CQBljFKLpNZTFcBOdpt0WnThQ/1dIcz7jWNa9Cx
Abq1RJeX3ZbuXxaLz+ezqOCq6uBzk8uRjiR8DgsLlMFJoJr95oR0ycGk9q9yeW4BrD3iwA0aF5hO
agIkVdeVhkuvY+xWq+nrNrj8fMbeF3id/FLPtjGrhEvEFY4dCXsWpUlFAKJWA3Ci3oYJOytMZU7p
JTfbddCIZXyXKeax9zwKfXEa5aQadxIJz7IWePBihA8O6cBoi6utqOC/XF5NUInxUXroT6tuUy9J
TI+Uk9yEANNEwRLFIjbdKQ+AjfnyxoiUIM8OYKaSwSOd/qzhQw5AQosVPnKyXcmZRm78eSeqX6dJ
mHBfBhrUEhtG8L7nYlMxAmrAyQjgUujMbAe9Xgq6xILBvtzYsyn8gcBvcGcthN93BMMKYNmXpLGJ
i/ZUk1w6OYHfnGX1RXbtxMecm2QSm79+8rrkYTpi2Mud6VylUDAoiWyDhaOoTVG4U1zgxllioyh+
NOdtP7RJ3pIy680dq3CNmkvJaPmJ9dHbWLi21ASa7VIzRl+RuF24DVUTfon2lceeUupluDSny9PR
hc6B9bmoqbyqN3GZCZK0JySt0JybgijpBdndr1UaNR6OLrEHHuL0Tj5xdotajUJadPfxlaeSGkE3
LGts3W7ZHAy0VsTonU/yqDL1uBpiT4x7EGeN2gJPd0ZwxRDEVW6Jc67GW6BXftJEND+NSE17rX7R
Wdt4KkC8oMlCrEpTDtAJFnVdjubdfh10asiHyXm9peiZqDDOFibJDM+PhFWUnNOin143iGQHlay1
GiDYwcCQ6UhwSbeMbsAmqezYEPEMIVHaIk4dcCpBtz+OZzcV7iCWMBz31yJetaj/iJSkLx+Uk/MH
t17o+GW/bldNlO5XKgPdLWHcpi+HKmU0i+weEYeqMPE3LDAF+KAPRj37jKVRLaW0ss0MhdDuw6OQ
2t9faaRvnjzoRiuak8Y3319R8eB7LbUi2IcGmAiJSSCfBLbkkCDkwHIZ2RCN8NKBu6jXKaJbIvjN
P8wFylAOPMMER04T6xEFKdW5h4JiOO3xj6Z/PDVMKuunx2XzmCyccFnSSHgx0iYQ3lr5YcxSJSr+
c+jdrii/aFHlBUuiPq5ERJYcMG7smYx+htFvdCEQ+frLPi3o7/x+KDSDqcBBuOGfTDY27htgvVed
zpzM1mcL+N1EXfd7RD0Dr2sKW2glQK0KLDGjFdnVNH6hywGGhrd3FtCtmHvMqYktfNHFuQmuIodF
hdVQFuwD3+vztt5FpIbmyKNwAhfNMgsuvS8oCgEyHCXIs5HuH3ml/BAPDdUdnv2cbyanAEKxIaNb
o89DiIkXznWiSMRSRlEYaP770N4/UnaXKApGB1amMK0efDXvWFJoOaeyngthg1O3t9pMZCUwbr73
5sCJexZb2Ugt0gVqKl4jWvja4cumUy0SRGDKs3y38Ws9x6KNpaIyBlu9nSdeHMtT8LGNIXwSYzP9
+0CwxDZ/ZKfVBfQL2cwNQKZvX+HK1j0M7jtwhKZ1TXOjOfmeh4vcTqfQ0ZxglvU+ZbktYGrSuTc1
LUYe43Lz9awPrfDDhlzGrk2PkHJZo3IY/xiJmScMZ7hhn4R93dRgonla8XDZjFR0yx7VIsGbUGnT
39elPRWO3Nl7NH/xJRGrpeGOd+hrPLoIvgdf8aazEFdE5gDGmEexSWUfAfE4kmoDsEW5KyejMpVk
aKPGxJXeCYCw+NL9QDEqJkKqDh9dKYa4SogYJ+gS4TpcHidFcHYq1lAijpMBPkCXXGOaqtdfFtTk
UFlZAT2fGGeEEv1ng9gWX9KDHdL0dj7c9PDVugxCJyObCFmlDImrQ+9v6yPW7C7OQrIT1f3oBoAH
792w/PLZI77Fm+HLIsPfmNGP3pfv79lEcEOFebo0dVu5D2WA6Y2zFTNk2/7dzjPA8upGP11lIJ1C
iiHx6IJ+YGUFFoJmJsHnEu22qQ8w84kHn+4Jbg9OHrdIO7cdO3TAG4zYPEHXLAushHuMDtRxk8ae
aePHzf/GHrZYXviEWRjvVBh02nXJQU9yuoxcPEY7IxRAGAMr476h3u3gHGnLpij6r3o0BGwMJFcM
6uqtDSA3g8sFPe4zHnqwaAo5W9Y9uGFp2lw0kOpvfLPCEzckXLJcIyzdtinrGX4qYACO+Wsrptt7
XTf2KEeIAAKywLhEfsTd7SS85zL63TbKGarRHW6FjqgADQL7dH/vOVUNrmivF2vALsAYItXnDQrV
QcSU/fC3I8cQnpdAH8sGbfVZv6LmodTXfCiU6uv2bzwb9dYfr0/bLrdgLpSj7BARHhCZMquK4/8M
IQSq+PCakzUQv+8C0OMJFoTYgPwqeb5YgIhUBH5BQHSVVRp+S65RS6RlbIf4py5BCBXu0VFTbUar
hnuxPqaQ5l9E4InKYoN92feppV9b17bTOofK7JXJaNOAXOuTEdw3z1sEW4dMpFSN5SD/BeAANRf7
D+cxaEMoZ7YFxr8YIzGPua1ssAJHzkT4PJF+4OFfnjzU7PhXTyqfa9pbdcP0ekx9T16mXcPlhiiR
VsLM4hOSH6+Eg30INuUKeeWVv9PqM2MkJOFiWqTugHHZoqw1LRD2T1L47iNBADroWfMTKTVpuHak
BXLvKsIAiFvLWFyRHR9zR4yuRHpMkExN/ygwdSO589rkA4d7hIwR+SyC0ctjMyFo58KoeiQHKiIy
mhYceH/q2J1KpkZvnt8IR6EQUf4Ymt7NU7CDSMKI8t+5wW4CoGIxG2V1IYwWBzBVmN0S09s48Ey4
Fzu8iahE/x7QVQB5pKcJVLTenuTf6HMr3J2pndIl+nukgV5ssLoDR54gXYJBeiEfQFkqCs0iSeiX
ZOI42nUp1ga1whqm57VKg1qnKJVkw1XF+ilBPpn46ETVUsovHCixsSecrzHRVXYa55Ib9kyd0Xn1
xGMKcwXJqwMJmfjTRmNnIdLQbgoxDo8OaCkanzvzQSY3ORRoPXXbz+8dKWI20M8fXfPRGmQmyJzq
FinGVk/WHGUYtSuddjvbs5eGr7+VYmO+4FNvvsgyDN5bkXEh8bwLHM64pAymQHW2JDh13mGYEIrr
hcPgdlGVnu4JofpzrQ5ffaBy6J1J6koXrIJGIWwl93pSqQrL1DvL6Oryh+5yfflsmG0E1qx8OPxP
tcWEasqESjjzssBscGZ6kKk88yn1wXVoRJ51U/ACV31+KAIqweadtMeNWV4XhTKyMWSg2i7aZJRf
ATNX98BIbHrSbk4dn8quyKcXFdT+RFcql8l6B9e7bYK8dAzPmgK8IpWudKAEzQNE7owUXgNwF/CN
TaB+XCAtE7e7KTQ+g8pOFAwMXX96OScRP5c0J9FY5WSSwyW7MkTMA467Q0J1nI2cBwc863+QF01c
WVjWa+ZZzmF+7i/Ngey5JnwheDISjLlbXthfpQZwWPkgkMmlj3bIhM4UUWOxJm6nQe6B1een7oXa
nrR6Xfk9mNneLIVc7OE0Sw7vz8oqiK9qGsR4VQc2ypfdVdlFJj9GAm2NVtcwqhabipD3ak5+4xEW
kttgPjLNrg2MgMj2+DEI8l2Pdqt5EoUCXIS2EwdlR4o3gn9VdcRFvLbhJ/M1tEea2yAbfV777c84
D+BDpLkp2X7wOBaWsEWagul4DpwzSCoeDSIzYfpzDACDemy4AHDrP496KVSLgFHzv6ZWXTecJT8P
5G3litGJefoGej/t6ZBk1kTZy6GUQqqiBvX7d50ssafJtWFY/1fGv/1bcNa/2+AQRL1Tcn5S/9bJ
0NcbId7Ikl8vmMrk8M2Uatv3jaqQrvAS0rHUOLT7uFrt5aKR+3TQI4w8iCjHg7EFN5Iw0BZ4NDJS
RM/8vOe6dWdO7PaH1g4qQI+5MIfBKv0hEb6vZdXytxSLAGRqegcNYZuk1d9eWuVMrgNtcIrv7phF
XCspAmHZPFckaBrxZawm99Np4ENslN5b6YL4OcjQHPrOhskf+Wma2pZCY0zDbhrcV6LPl0OBKlKq
cS9QXuisIAXiqkdSZxQaG5eVKBOb4lBH12o27Omv1n7UByZ4v+1mNfk33gSZ4AC0MHbTvl1mSAgd
79UVpUcS1xHzSpyATZg+f787QBWqI24LO0Uuf490xzF2PbJ/VXEHNr9h255bGYrx7RcPFekQmzwo
8lQTm5sdXYoCo7M8BTDjGjk7x9BRH3e5YunaREMDj6ZDU6WCd8HS99E0g4u9za/OnmLrTIUivwFd
YLavcie/I+m8nC2YBzq/yzPWY5NkcO3+UtGjl4jqVlXxDtySQ5vzaSVoau0xDe3nGLQpMtgVUAJj
tcnWg/vpbGF/qOlR5qY3btesvJSpc+D/JDCMQxPBHuyxjcOrD9eEtVGw+Nw+Ydp20j6MZ2tMjWH8
gcZH69l3eRHdcakHmm4rGt+MFMHzQW5M89y/ToQhtCSUn4LzigMM3K1YWkmhQQzsBBex2Mq717JV
OMxEQ7CgKc4zbyKx1CHIj+w979IIKXF1iPXqnKpm/mZE0h01yXEKVvlcGxHMmb0deLokbPPLE5I9
CAiPS3oRR7HAXl1YZmwKrU+2JvAfMe3eJWuRE6qum3Ji4wTG0YmMrAReHBCmJ42dt/vNgVApNLjJ
c7grgGJ47rv8Vd2SZDJME4N23cR4VGVD/3EF3yE0KVlgtg9C+v4UoBAJq18W+jYrCJZw9rfrJJ71
uR6hCAF/UcGibwUZQcW5s7BUAY1cUu7bAskC3fMlkeEkLItFHOvh1P40M6Kz3Us0cLBIOfRSXOUI
w98k83AY3xqJroG6szorG4QF5StqHiU5KWaZnUlLrKeky0NAEXscpQ21M4MivjH6jaAWoB0jM+Cs
N/WzgaRhRjaOKGLXSjnbX3rACTVmC+jHNZlHOW2x9pkmoH9z2fUHoIYfANgmVrjRbQva4vkVyBlG
ZgUGKlNwbhw2ipi9jBk6+If+6HjDiuQNuPA6bRWRXj8q6a2fZliMofgQ914TCx5dO5JhJMRwt7aj
2Gja/SYkt+3GRV170/UwSpuYelvVHCK+1k0IcJ/ev+nFEIO9vVO7D1vszX7iVPprg5x9Mw4Kjmj1
Vp2DQTKF8Pna055Vu+YHGjYQ/gkM/1jWdWb6Yq8WOnV3xy6nLsN5qFxYAw20W0zMifjRdbAbGiWp
FkeS/MjXMJKFRGKhu2ihIVIH213zTXClw2hFmz5wj9tkbxyP/BCbNjD4uTDjGIZDoO+u48aNjSVC
BTx+ydLH5Z9lPN21KMuqZr3qPmdHWq6I3CwaR+iOrUL3LX+eHUN0MEXksbWvEYualJKfOR17zU5K
0cEV7/WMCGx39JNw3N0hlvtMvxu689yNBN2wALg8joQxGGG7Ul5yG8lHWDDtwfdBRiQp07YAiyWz
etbm8Eh4C8JxnWZAGwc2MhMecEMAgmIWSkItip1gVcWdF5TvSaPX2Eb37s9xEII7z5gsH9w3vshL
uUCUwCwNLoAN877LXjeFaL3HLxv8Jmf/0IPI7AoK/NrWFKU8Klo6qqSoD/YUXB8wm4BTzL/AMijW
C4SxYuGCJzVE1Aawc/6K1KMqIb/eVzQRRkeSG27fse0bRbB/tnj7NIIZSS65V86w6ezzlFqq6wa0
S8V8Su6x2cqgY6FTZYamQ7ZRbw/p4dEN9Nro4+WuMa3CyCQUU8MA5crGMAgdhqWgiNfVjVMP5a89
+NqDck6Wsdl5KBMMjQbgXnLh8EGgIsRLhNTX0OL8pplDdCvXmPr9Vlq7J/EUAmfzm3J377ek6oyJ
mgqPs2RTWsJK6/L0MjINY78gdopCQrVZ3Xxna2vSQAoKkrMWnzAUkyir1kC1gQTjZM3tOdGoMRCO
xZ+qd3/lmBCWmuCbVYRaIuQkEzU2j/b3SsUwgiV3HZkuoFMuze7/FHWa7Q4/bVeA5m4gSS3ZZYre
31HifNq3Zg27Nj41liyv3WjoeARzcoVa03UJDJzdSaNBnWq3R3dKkXVmeeCVThpskOWq6dSbXzsg
OnVnArRJtz9HrWuFmPhIldbU0vyoiL9n7Hn0HhHuQc79sws9Lwss4hOWTxy62sVGvf/GhG7bdFAH
lmbG9snM/6XT0amo1sZCDZi7akU4225uwgNDExI9TJsyEDHcFxlhCbJYqiEjr7I7wrVZdSrh9X1T
VHiE7xPo/4wDRzRb4shH+HBWiXg+N8ueqMYQTf1AcsFbu8rNJpRu4wF9DoKRNdzjhrvbkY4KS8ak
LudVqz035SXprBf7ahil58ViEX8KdObiFNWO11CBTOWflokGbnhuHlCpOyPQvJN9N9IZSo+4sWoN
lf3ABW+EyWnV+A9s7tBWGHKieoLztOZaWglgTSMx4C2jdWhHdacVimnmkSRpV/SMNvECYUKI9GSJ
n0YF+vJAq4QWyQFYHes6YOTkaubjOtgDojF2eBTXVXd14hu+DQX4PwQ6nceIjsDJ3IID9ANRPcQt
ApHBmwRoNU6cyO7ihvXJIurkaTHZf3Ap4428QipJk96bH76hcC1PU/qe6nYF+yjIHJXyCAg3l2FR
YwNPPTaf61oyTZXWt3FOQkFc18KOuNaCNk4Hwcsec2FWlxlj4F/irA1GQqMelDHT8RZhFwD0kqjn
U+QcR1Sd7dNnkGFlF7X8ZeDfXCuQ2fx3RJUXCVYxjXkJd628VnKMg/rFX2jcJnSrDlC3t3/nGdTF
QaTjMgqcSD2GFKau0laLuAT9lcFlczSwJ7jfTDmyeFF5YBNf1fIJyDq+LViMPptinHq9MZ0/jH5N
6/wLu2VE7vZHwtMPEX3Olx61wsGigJ9TR2D+gVonEKFFHAuowrZv9iZCYwyMZTuUhI1CRF3sthXy
yXQ6HMsLpxqsLBgrA+gfKhfDasXP9NJQSnDCenT2FwpCxg+gB87i6BbwFsDBdMirOL2d0fIDpdON
P8h4Y19c3b7lzyPz80Cbb1mjcvwpbjlSHYxRRUhOZnXXVxhircj4bDpMTvTeKTuI1/lTIP/dYWI2
tZ4thFFUqLeBvMP8q58NG/exeHk82JZFpEdl0/vbXHQVUba8UI4fwwm+hz2Hb672UbT52t6BJ8HC
BR+3ABmmoJlmpAdQNZ9VuRHABxH7zMB70ls8LUWg1ooFI0DbuPFnBjiC5Pe319PKeiUGozT3FJDD
LBqxO2mkkg1qTOdOEJcTkNhjT1algY4SahkLPdzGeo5XW71mTWWX4orsupPsLjHEH+XE2wAbCLtl
94bofqagYTMqJLmmhperjPmSzGM28aUEJUUQxcNrPrXHh8sXlqxyGogl8LpYcjeZNR3wXxPZj9/J
e/XPqMqPhYnM4VBnAen12DWwJfBZKL1L+vQl5iWfOMtbM3bxSF1jFcAYmmAefjeCS+5+/r11Sl40
3okUsC6hGvMPV8wv4bXB5p+yFSzQ9q1KIy6Hyha3qt1YglqkGu/NsTJdheICC18noPSX1P6irN7M
COWF95RqhoH8b1MllMvp5egnLERti2BwWeDPDr5WKVUJZ1sFrf+EM2nH+GbDprUfo/sbHQuJPnyM
8XtH0e5eWzzwvjcYPrh0fQdEQid7ngeEVET9/KT/xYn9DvLRVR1fKIOAT1T+X8KEJftB39+IjRt3
u0nlCK0oYedo2QHrV/hfh9BQiOcNP/LOJGXGXhxqCQORzXhzyiMkpduPBz49DKb6Gu9+9bjDD0Ta
M6hNGnXtZXWnK0pmZjH1MajOJvXDJvQXpIY/eIxVQd9CrOyaOJQOEYY7VwWFDyY9oAU0BfgAzHqX
BI64XMKlzM2jtGUS1uoZ852UNE8/XoRDc1SOxkvdFRGwbiLYXBljB2Q2Mpyr3oK0krbEx3oFHHo6
v64IVEv5ouK1atenEcQWR+fIEvKo69a8ZLZQSXSaFbVdI7mSMsDhNec1wMGbMiZykwN7lNy5an/8
2d/uI2OquQh1IxeWmDq3YGP3BHdfKdXxITgE2Zxsdyn6nhZ0CIuZPZy9QudORw5SU1oK/7buorgc
xia970R4aVK3v/FsIxRZUmrtyW6uPTAb9TR83n2UnRD0wGkZ5fULuHMUgcuEnO5uoCh/lD3Gi25z
IiNKKsEVSFiFgwPcMoiQ4MUb3VruajC1aW7wFXg/3jXEJlWPq8CZWmInnPdwXTZBClkqbH8aEu6l
iym8ue918LauyqcVEMYAke9ijJRWFXzzGLKsIeB1O0VkkyOrinIey8U8Y5SINFklWllJ2/IQZQ2k
mmKKkaCag1g3LhJkgL44lCJVMQvLc9w23Ir2myYUWFxSpC/lwQFK4l0t15edgNIVkqYiFGbO6Lio
+VFAiATQqKEq0VE/ScuUgbgAlzmiLV9H22z8pSeQszFpQGSQukvanNU7KQ+PniVoq4hfa0kEaJ/8
OSOCCTtu3O6k+uOMp6cs6pZurSNCp+8U82FHIFY+SBWSe23sPficdc1pHKpsZylOoFUQlOcCG4WW
QL+95uqkrTkaT34P6BJ0iUL0gNfbKk3Ri3tS0vbtw3rMr6RNyk/TxhQkw+kON07TbEVlAX+JY/7u
CpJE/lXPbP4wcqbnf2a3jhAlJ4rzSZEK6yEg3dI3+dew/AsM0gDup3snEhtUeYR/GBE7sN2z/NBW
o+iN3EOSbQlJEXy8JFdkGDFNzIXZY8+KI8Rcfp6e9tUGKZjOUfeSuKOG5TXrYtCIZLgNDKPxqerd
/PsVA9S/Df2T8Dq5eCGDJ6FAr/hfnwQkUuRCgghPuSJx+uu/y/9nQ37871JpHDSHPSV3JnmoNrBl
yU1Uo+WmnJQ+1IzslmThUWglw29j/OcIA277kUBCEhJu3Xa5qR/FuQfs6sQeN8ZseEVYAzQVY2oz
A4GUxgThOc8e2XAqZ4Z0RyL8IhW8yX7rXjNWCMdNMuiga8mrQduhFHdEtIIxqqtqoNl7YWSaFyP8
Yf+MpRcw6Bre+4gljyMA36M5HwfNMxT7XUORfo7IN4Ttzf33fE8CCKFdsU3uoBF1IxYYFJFTHq5z
Bbn+gd2Du5xEySN/DZTpDUHYqMgKptbRBPn5ZuH3/bSe18RIG8Gce5Fbj49u0o3RsGP20IZHccnu
APdCTUBbNo5FOJ46xbC4ohUxyyr2h+fBu+u+iz1h5RYThcwGSpCIgRVJyU2J2E4dSTJd+qLQZhzC
ahlNIqDB9n7bJkQi+6Qbahhw9OSZYobBpvQCwMp4r5bun/OJkV+/3Dohk369/6b1/1xQgKFzKbpv
y7sfcS5FVYu6GJ/88v4SqBdws8dM0L96mp4rw49rwVXo1OT7s6NxZ+dErBG3P9lCwYxX/1PVP5cO
IGafNYjC5CxAOByE03EnBNHJTdg/7DkQr/Nmb2hGyin4KWzuDaj2zb5GOnGizs+SSw3QtoocRr+V
HncxyJzhYJIct92DHnAeX+nsxE8Pf4CPbd/gqhPHpKT9cQB0cHP7zEJ+5jq9wd3zFKBD7MwlMRbv
chb68GBilWzvlm3vSv8SpIy6j30Gp0KFS7Vh8HTgU5G+Pyky7t7Yye33KuubksnjPo7Fjdv5QxOU
ygKTkqyPU1rtzULoN6KHIbNH5fpFueh6bBULOgM8ytPBG5kDu5GyLaTU1S80NM43nwZBr8BJwp0S
y+RfAlVnYA10CwNpLRiOxZv4rSbyECvQNy/xh/9sXRQWx6gH6F20TwgdSTBXy2KAypAy1EbUbJea
cvOIfGQQrpKDA7NWIFZUW7DVDwgB1t0w0x0XAYmXsGfJ4bE1Mq2l0P/v2O0k4nUjGXxv1ATyxEu/
XUDepGpWjfSzIfzKRj537g7wkeZ6hpY+ukLqz2b/q4suZgR/jx71kMtj0CEVaYB1GTUB5eCo6bm6
QnQKvwwcjEi3gsu6EFFnYKOp35Yhug8mCRmeizmt7C7Xa7aDqi3f04sjZ1W35gokbA/pYUl/tq1c
F5b2HEtQ3I3KFaEtgTU3j430cPAcj42MCdScdyAAI8Q419W67mATZc1l+R7v7AedQT2pEveR3cMV
l31leWNAXeUcw3qM9HTmcHx+g6IrsR7a7qjjFKaYQM7v7vcAJk9c8o0Lsf7ieJDNFZ6htC+m2CF0
1d54NZHNMF0dY0U60LNcYGeRpNvcTywYjc5Q/HLFVAGMpgNNg253FHw+A1Mnra8zL4q947xAaCvX
wrgdTRWc43kJR+l2ULRijH/smYYVFLxz6quFV2gtGd9n7LO3LmHzEiOd+w09ZX3lyv0JFqtYtAbj
y96dPonu375MYu+gZj6Ufrbek6yvaGWIRjw7k82qoLkORPP/bsS08OpHFowmRkyaNvPgt7F+ANwg
/2bK8ZwtAEbH/+ACoZffSicoSI68l6ddBJmQa9H3OGDu0et1N7+5A0GGDQf4SBg0l1/kjCxCwzQq
eNRibyv5ABvY16UoOk5dCxyYQ6Oa6VGA221/k6dPtsjxer5jKI92D6UZrSASFULqe+NAEgeDlKYd
I7b1jIzhvmWeNzY+O0KoqUMCOeHtNkKLCOkiIu4aEACqfIXhgeU/1XfZaQP3B85DbEDP5GyXs34f
jipR5B+etsqUGtRqrb29tBqY6sU69tyvoNn27thJPOGGZwvJR6mq1ciUcw+kGWL2UGbVGGFETUYg
SC6pla+6KPTaFkW+AIRWajlBSGYimyZYHWaTYywSkXjWrk4DStu17+Wr3BKIkxUdPIzvCTB8yV7Q
Sbm+acohc+SjyQ2LZslSN2lKThvh+WG2ZFolxQ5yKWuyv/p+bUYahULw023T/WkBAJoeDPz4z7QL
hL7hJ4cuQZry6vPuqp+/MGkfBUS4GccRfAqRO/tYqE+uDxok+bDtUip6u1YdrhWBK0jaW43ONspq
g96kEq9rHBbvwfRkrUppCLf59gRihz0ybWT9D4VivfybpBfu6lOs18WzkSKu+XUU9gxOzVyp/APl
3nZTfP0MZatB0aguz0iK+5np9gH1S5fQ7fMhteXJmNIIizKp9r2tOkV1iuBdsPaYt2f/rVK3HGhK
tV060y/VfS83LoazaVBNMFnMhVtIoUmwhrlE6oPHIccZHbuewFGd4NNl0Y671uMSVo4KPcPJC++V
K6+I0/ndnW2AKESAkzyHo5S8poH6tGDpVRYegFZG+CqxYnjhexyPiGJ8Dh/qY2zr7+wHEKtEHygE
3aDA8Q2LbCK/13gjivFJQedNevXe/N6/bUgUgr077Cn1/zS6JW/wMq+2EB2MH/zCJz2NAQv1LydU
Byh+s2wNH7wNZP4pnmF9Es8s/LOHFY8w3Kz/0x4fJ2V13wIndm6ySdfbI8OzBQxxiSSzCEuwJ2SJ
5FxY8fYJlgMHwB6t2rymgmKduaDcXS5n90rvDe3KEmPTA/oKCg7CgbCic04kuHPwkmwxWzCrYvk6
dmNPwshMiajpSTomeble/tkKSKnNfMInaBWEWLoftHsKx6TqsqG/z8FnY0HJJuPQPvfei56bHJpK
XIpJlJu7rGKnT6zU2X2746XHKYhk/hb0VaqlgHr2pCnr9aSjFQMP0y1mYZr656biydlxiZzlOJwp
STEnFA65zYp3H1xpETX1LCk8WAkWcEAjivnan9nuIDos7MQtxmjHBT+JyWvCyMJjHvAwPVurs+j/
XzobjNlDgLd4HdtWHl8XSS9ENEHAz4SDTt5IlTDx0pXZZGVjcaFE0cZdvF7Ya7hgGwDeUVSqucvQ
QpT/Q2TfCit95BHOcxGIYizgxCHoNaNSRrGqmy7YBki0SK8e/GIFq2feVBTgW4HwIQR4RronAnxO
a2he+lfCp+0sPWumeWBl0u5o7YWcbCVuXB5u4tF5oXrAeKKZslOYGuMc/NMBeVMSlgkuLD7qEACZ
BgDQ/8oA6JXkVvPERHlu79MzR4Z1PI3lSXcxSQMHmht5Fhfe/yCCHEHZEWqsWjOyOwLhomk+G7f2
1KCEIhsGccaGrOIFnYnAgXFBhcRasQ+gG0NlpQiP8p61KhSzDd1KAsFWlOOf1Jiw9JGhYv8mWwdD
SqWAWPsbAwXMkSdwy13PlgYWLvX1FLeJ3OlPoEawYnhLYq1RpywsfB42yC5JqX4TN1uvo1vGjuHY
eiDiIXkOBtJs7UjDa5FpfqnGNhBCE/J0YLC7aJBxQwGQDCgEzXW3hpQFpuE6VFVTDn9V3P5LBj28
o6p64mbaK/mGL022XKheZMJJzFKH+REPzVmlkxMKyResqw27i11F5w+lVNY1A0uax8gKVewzqWLC
lc4U+Bg8xbbOKnPIJMK3qaU7kaDzzHhV/XGafz10SBivBQiUkIKIegg5OV/H0LCNlguPtYEAGO6d
CVV2HgwQ7fJMjamwhYT1oy3AmSAOlzoUBTBvz8T8k/2tnKe3atMIoNnSROrmMFJZDHpcMuNweEFp
5Zgs99/hqQ2flzKMfsisntBCRuz/7TUxoA2pw14ojjEWEVs/cL3A2szUhwOx2W+EcWsAKnNK4iqV
mnYsmvCpTxIO50WpFokAuD8jec2m/VM0bPXJZ0b9Skla+5ukZP+SlLp63QMJi7cCc2LDqZsNCXjA
ghGIIIVDSmoaSIbBpJtX+d/RNX4benHvzdwVMkU+lZYWU9d1sBZU2LN8Lbzh+tFA8g8Z30F38HcO
xSFFJSPyEWeY2Skn0QJcEu4JUQHyiVc+CaWzzyIYZB0YnLJo8OkM63hciCHtV4PQxIzzHrmRb+rv
2x99a1F3kojBrjkrPj2Ddg1J+PRKExHoyd4GuLWOLLa67tyLnvotMnO00VDkl/mHzEiN5R/5pc7t
u4ODjdAcbUe56vlUv5mqo4BTACKoS4AWu9Yfh2LvWimngmNbHV4YVZrP+esDJqumXqE1FpQ38Mmc
Y+zxL4bMfwq7pc7kFo5Iun8N6G07g9Rgak+GsMgnTL1py6/DrjxpjMXvZjcXnw3OSynxBbDb6s9W
UQnSYXn7MyUnVWq3GPRy1hALYp/6j+TvwirkFFF+/BIJy1hfTDaJsBlLCbnA4ZnUu700vg+KSgsO
7Hm3X78+kWDeXVK7ySqQEJZuahOVFrs0CG8dSlAsrRUo/N9eHr+9bFUuSe8eLbkH8mX1Genp5RPH
ar3qNDmbDYoiwf0IKNid+yxU4g75qc7EUR6pFWst7JzNy3azF4m0iVXO32TQpkFUn2LjMV4L2F0q
X3RHeQ9gGi3vVxRS1ZyzeMVvHZD1HTfyMyfOOhKhYdwQHdPlRthSO9+wbANIhcSvV+s/O/ch1z7W
TFzE4DjL5MUi2bjR0jfVPtgph8Hn+2dQ0xODSvDbf7pEDYOXXIRD1Abu6zCZX0ctw71jJg+BKN4Z
0eXKyYSNEyMJH4GZ/kbgKeht5JLXBRqXsfD+POh7FxrsI0K8Hn7CT6f3x3yaMscdX39cq6gdn0aJ
rT0ZycE2NK8YRrB74W1yc8HXMPvJ0a8P8Ap3zYGT/ppzqqEWEWk0V5zT1WS/VdOnXFHZGiT4wIci
AksWFuR0DQwCWvguokdwJ60KULeyraNDhlqgngkF23EACur6v5aiyyiVQnYFXzAL1bju+YahTtvw
NBMH4hSQL3J+xGmwWTfMrNUe2GIlMQbjkRA2ePS7p2tZMxqZ8MMpWouBBawAhHALx6Os/uBK7Qrn
fn9x0/X2H1JVH1qppvY1H31HnWzkbdyBWv6gDTLdDUy4pyMEebGgBEJOk2rVKzluyPlKHP2uglZR
/m0CwwH7irQJqrCW72m9x7CQ/pidbw7RXZWLhTG3pyYdqmgFQjH1tv/6PKB9T7jJS2KAepieikBP
gH/pBknxFFjXBzFPOXX+O16EgJiyDz9+1NVinm+wrXXDSzYLrXULG6xg/oK4/Jv81YPadkWWgbSv
LjASmKIsHtWyy8LmDqzFtV/6S4J0CFTPPnJkBLKZ7ISJOG2HzyGNZ4tt6iO03NHD2KWPmWdSm4y6
tSQSxq1KjwNLq3/hyaGl0HZ4BQKRMmvTvHxpzJFPWBBLfJmxfULtRCivLmRIGcGCvMB+t43BCOyX
jJeuf0CCCkXcOtwsjWkEIil+3BZzleMeth7wAkaGootGzJm35v8MYIHuSYfZLcJ1fQ2N6hTTEQZ0
K3eKDX8Dw1tZjziVF+EymU8zh2gtAw/9v8qh1OE5IsEv2HX8F5NsfJHrmRDl9AbD1a5Q+D/W9x9O
AAgjqugdvhDRZcQwiGyS6OiVNWITq4n57TJEQnAOUQfpfpkCaKMRYW/6cdGX9XHyFRUpmtdnm+PS
rY1adl5GON6m/cwbiahbX7XVpUKCiFoDS2kD4B4Cde9GT+wPpljD1fX2qrGoNq4y2lohtQu6pnsM
Fy9hKqwZxOLfWmdKDt0rezlCbFQfThSxjWR+FVAT4FSnaRY7WRrKjAgfFGiuo70gVrHXzqqGReKa
tKqB7TDQLCPwaY1NLhvosy3V+0iDHKU/fD7L1ikpWI5iVy1IOuyFmoROXxtysualxy2NZ1knFWKd
38YN/eqX9ZP8K0Xch/0S0ZBRyHXufggJfY9wCz45UMCOOFWv35SzXXZzYO4oEdu+Qz/xaaUmtWZ8
CdZ1G4QqQ2mOKNlI7XHqld1lNs523HFms6DKFYLl79trYKRrr/YxtXNcXCYALprIw2iYfQNrJamd
V5T6ZtVEi4yVLtEZm8hJX3zRQURd5OszOrOxId/8EwANBasUbnV373jbOHajbuyMl2hr/caDemRi
mzxFzCLjGJUMh5JxppPFinG3Af6van4pG9RjOSbwhOHwjwBi6ZS6JPqFkfA0vGTXIIYuQfWVL4Kg
RahTp1oGZHTqIIh+bRo/+pCRKa+yhnXmDWwRS/hOzFf3jGRQEb3zchB2hU7frsfjrWkni/uWR+35
3IstmbS1nImjcXNQO2f+lYKxs+TuhwzttdTZiHA/v7boCO8gYZJ+jwuya4AIUAwUDYnPELpeHfx6
M/FT+BcfZ8ybZp1CB1B8nzoT/3g2VuytfLnG1LjRGR9X69Q4X01ADO7iexcA3mBRYjeAxfdC2Zok
7sZaWAn7gty5zuI1h23dgehtFv5rHcodfjmTL36xSZhprCWvmC/xN9dXF4+b9X4HbiyJIGEFeu9o
3JM1KQOxocsYzviLcSrYSwpdKovDqCQRWRf9L28pc4A6D5l/y14XpO+5+76f/j2bw9OGvd6DbFHK
IEGbpuEj9VN8QANR9feU4oidT0g2Uddvo9olxqWCQZkF1duo/RPFy8lCQ4gyUC1YNfLhPHhp6jSS
nVUtEn7EXt0uy296XRR1nxht8ZqPLF68xBpkVG8YZHmwhuGHGduf5pZws0s5/io7NtKEXRLTsACb
t2+cCwfmE4VJt2PS8O+ew7bBQ/GQLsknY03TH1Y4r0AsCZUBKzLUoh79IfGEtIYMloJOLlv3Au/W
IkGYi/rgF5yUdHIhs0J6ZKMMEECsKrmv9VJiNMY44BDy/iJXCiYfd7453M6/vrvIjwnY59oaZ7Rk
DstqPxHc5Dr4GpOROhAjC4QZeU0PUk2HCmAtZ0oAw/g9+NmoUrLY0qTbc/GylGkNyaY0GbzKnzQN
jv5wAW3dUgY/PTTKsPp+qyFLXCjj64Dt3YyFhu/JXhB5vCYRAdKawmqgQmGS7lo1suLyB0bYo4sn
S+1hssRLvJ74j8ZXdfUtDaaPmjjCackQLXoi5+GSTgP0f3h6WGRjQIDA4DNBE0kPpF60ecbsVUf2
xZ/rWYl9jovPkzqrzwRD+Z18i7zP0vBiVx4+NiJjsd1owMDVfBoK7i6kisBWfmQciWuKx1UbF/15
bMqetrtaGn9dOXU71pD9MG0nTUO047AtMwxn0PGGCNHb/28p8qWL4Upu5Wu77Ug4yuN4u3WyQEp/
6Qo4epinVIh71kQpbd/g2F6vRBEVAL6zaIansfTbEcqzl6NtzJnfrKbDNXsAW/kcXBr6atOQ6dO1
Or1icJPRw+AubYkG4TKDuyiJ9kXMU+zm8OKz73gZBIS5YaQHFAQQewSn2c1lrvAVEVasEjABYufO
sLisCtlaFGK4lR+0Dzmg6ANHSYfiy8+8QKjosxxn3ZgIyHSwzEIK3oLdP5vthttJ4mMbzyCd4gfF
N4HPXdBvZSYbSkHM93NHvsph2UtNyyoCgbp9EFJjJkDMscVAIhN7IlvnW9QNTF338xP1uPbp9auo
4uXqXofD5H/IacucVaswoNRAZ8Ra/NXh67soVKjKD1hsVoLiEtSQzX7XUv/RscG6+WbnLXgRaWbX
/2K9bnQ2NQnEKnCUi0PSD7NLaAdhR4O7kgDIvD60Vdh9B1HR4ODF0wNMiSi1D3/tXG8fRmqsrkQU
3GZg4kgUM4FkSgdJpg31uMyQez1Z3WUjgaACyfvw4ZjOoVDJ8esCZgflHztyxkpUVtDzb60GII9s
W9yi+YFtL0ugSAQ1+aPygRifqwsAloYesFogI+NerEbayTFOqiwj2iO8VPSOThnopOiURUNLp1E+
powR01OsUfKCm+2Ul9a1DppRksYG+x1CzZHMpNd8aD3dVl3VgFeSajNOD+x5rdv9z712ICaVeqLg
9iF+OJeT9ezBiBIeRR+QTDPaN+RhgX0gOi1xgMpKHME384LB9vN9nSzMqlP25QMMOxqRCI/b6n3F
SE7kVahkczR9EXV8ch4jZviY3JwaeUf/RFOg+AO/qcEslFWW6kChK2NZBtzMdowGUxbbvVamez//
Fa4Ulhz18ZA9A3xVTkYMI7PHNlODqnDXr16fyjGhox46m1y42KkH5a7x+FhEcL/OsWkd3eV0p+2e
905oKbOwFTMKgNHtQmOMyBmvqnj02HRnz8s5cjTh4ZpTmjxpXxgulA0GFm0JYEA7jU+5Dys8Cfqc
8iZXE1FV29EBQhNyyhRjQf4gaiLHAdzpCGlv8aIH5S2ekPlyWlKtM9scqG4Pc4udhxHPUW3pxhy7
f/633YedCiY/MUaH6IH55QCi7id15e5BMN8oKgXgUzgXoBQ3UOAZr6VJeDZP/kCoWNOeNB2/ISn8
uTkKwB10mzRL/IIZmZILKEMczl1+oGLgPdHFMV9/mjJnv/AuvguXtQ3JLCzmBHKyWgXtqA3wT0D4
nCKCfaF73E4zYpJXF7qYccxctvP/sNR01qM1LCpcLNg2WEqBsoea2UctQdq14wZ36aOoXSC7JEPz
XAv+XsYrsz/XEnDhuWAKAi4XvYo5ieeyw3+e7m3R7PEEeIba94qTqM2znVAwtSFkMtj4kQmV4V29
vK1AvNZSmE79cq9RMO5KTtil5oafAJhs1zQQ+btS9jY/A5SCskpi3BODCBmfmgfbgTce/nB4Batr
AW+LRoWm89kZigI/siJrrB/NKK+HkAQzLbSyYU5PXmFbA3eKnt7xV9sFEGoNJjU+ZLx+6MVH7ijA
abgXDndi6r1DUxs4mbD8UnRF/2Q0vBGmwUyXM/q23zhoLQSXV/4PyW9m/Vmr02S1Eax0I6PTinxt
7yJMT9XoBMq7+Uo1kAv8LeV2Wp+tr/lfV0xbxSAsLUFuyTd/HXMqjLTpr1O3otv2s47nRNHsvmgO
W4Xp+HWP6lGRUHHygQ1ZajkiW4gCrrJSXThAGGnEY6sgOu3pfrDtpXkXJrPTpxmSkN+rM9zzoiJ9
toMB18F69MkQg2khXkLMxvbuIvoKAynS/nLlib4ToSW/B72K/Vqjcze8iPAg828atHOPmWgGkIuG
02ajo8hEl/425Lo/F1+QTHEd6u6eU8SsANpMyae+uAENrYRzLo6bJBT5Fb0U1ZMufvE3HXYzYQJJ
qp64FLlyS6UolkWc0aiBihjXKBz5xr1FGVPW2aAZv/RCtFUHdowISoTMH4zcPdVenILBXJC66cx9
EF+6HaC/r1iX2nqTnZv1tgL/hRVKcGJ/G6euTot8kSDTN3baz/9eYCrSLpw1NVC0ZmZ0OjzKECfk
FC6lAudJP13UUI5sL0SHiQ1q6DmZqqMKLxLKAPpIrzE8I5xv8g5WWkwES3899xDmnQ3Z4WMHJhfp
hB8lUY7kusv+ccyLUIGARqEE4EoryLBD3R6EeKhyvsQmRkdzOvq0xvc5su3u/6d3lQGcPiuhxMjm
ZYkViGefH8SLvt+Jh6eMeh04/ABjA+Tsq4UeINEVPZPiLajJhuBcaPDSP7+iIJOgd8Mqt89vnhjH
4v2DcnBCv+zsGjWfjq6bcy8748ByDM9y/R/egPpOCdFSPl5uS9qiOAcduBbi0n7gDcEOvR/tBGoJ
2MhWU/PjfaMxXryRMfIZcU2/E+Op8chIYGo4qzB8/obmP5NCEuJ4binvAGR7gQtramyNfhKOL3gg
jHGl+934yxYUhm1HIUsipNnYu2I2KE+qdvkvq5rkTw1AdAhdTyO+MAVa+69AshYccBxoInA9ZRv0
mhJ5gQPM5BSfg3qQnAh4ro/kfsgIKZk/cl2cxqIWMUOuzfpo009lZFeJ6K5wbKeLHcMUdhliGBEu
rIk9tQjyP97bRxDRreVLhKz8PCtvT7uKAS7UfoSJVP9zsbVrNHYPXQKYWIcBC/ampMfTjbEf4Eq4
tPTx75xg8JbAnfkhyfQ9wspXxM11rJzZ3xhXjTBuSi2B2Bryv2mwtBMyY6ONnaQAKCIl8B7Z7do3
HEBr7/m7ZDy5k31wiT7s3NYTWyBHnE6fUAWxsX87m1KlMrfy/fF/QzzOL/VuwjBWz3QIvqXfqHq0
mDWdYzhOo15wmV5uXT/XEWdJ4zpc41ZsdZX8PyOJKtkeCfG8Fm73IStsbjd5K/L2nhRXvcl+8MWh
ZVX9TscXkbPLUEPxCUhdeXV0aVW+1eUXreeIBl3r5bZiAndKzRbuJkPZn5UygO73ctKSTVAAI1Ca
f1jdfSuA8ueYcAOtWbEuay3G+Wm92uoytMllNfxLXWLy/pulyjnWzFT+cHsQsYaCvuLGjnt9Shlc
j9lHTtj/QguU18NBbHczZy6BZHPU/MCpB6H//3kNL76FHRB3cDpI4ULAo3DEih9Rxdo/jwpUGQgJ
Y07frVooXAnhnQjcPflhCh+riFZ07weiZTjOgsqcwJ+j8ZbkP79egA7baOFFf60hu2nsvDoZ6u+B
SKbVMT0gHXcWgonS8giWjKXLMCEQxPWTwQ7S7s8Z/nfVDtWftWS27Mm7lE92dUMNpMr5qQ46QyT9
kKWFG7fhuDv4g0oGOKZhNN+jN1KPID3kE5Ob2FwQ8Lzi3Uhgi+xz+QnzxjNU4bo24Ewf+JvbnBwR
kfKliWCehDCYCd2pKmkUQ7MHXdaL27Q9G9sVdhOwElt/Ig7lDririEL6JLL0Uf6/CeXBbcYLlSW/
8O/vmkievGHHxQ0hjzm3qbXp3p75vv2sCdAU/2YMi+YN2XXKkKJ8r7k1H2r1I1LW9DZhZhikmkbO
MJn5ZvAtt1Rn8SvETfCmaBsaS5UFlbct3toAHgPh35jwzjZXsCHiMso+SzYEBhvd/9aSw1D/tS/S
Mf5w43qdsjWCewApk9OEkSOtPjQAR3JGww+EvxeX/77kT/dmupyFj17jzle8VeA4KJjazNPmqrQX
w99UKHGpwTNVn+bhwpMqk6FusjWMUaIm68q5QdBdYPgjRBC+OXgEu1q/8pMN1JRtCqds7n0iCs4W
TXWvFund6dxjI9ajO7q8KJueSOXFjJyfHMQ4AEpSbgFieHa0QG9YM5WhYdvVUSPjrxJYtd9GM225
N9K/LPflfBTZdrnfU2pbVXSXtwK/R9cOPxtF3pK5m4Ry05/WQrEunW2bthy7HwR7+zplYrp8MX61
+HeHWYkZXOWPxv+34v7n07X+yy+5wWyQfAz7+e0wVwGP4Z1J6afz4+VfTxwV5ZVSCeAsWWfVTG4S
A8Ki3Y67hhs2uivN9ZGaK5X0aq9Ph+CFN1x/yNkSNKtYgHwfMjYisW1sW+BovnIbvmKRL07vJqi8
SPV0UvWHExtVVwBCfM2ooI5lM89tHzGmpzPEb9W9gwVqrDJ5g73o51bKv2HQbHWSBcnMZU4TIWa3
MiAicUI7bA24LeUi4HDJkZl9ypL7TJYQKnGRgiuHQu1ZmVseEhiQnD3TScsoUDcFMx902VqkZk5E
pEz1GbyDiophL4J7fv6ojytDcFl0o3/lRgK5ACjcaKSoUkMtsElLIjv+eCbEpltF/8DBQKaszkKb
TuahiXOdDdNxNMDGip8RjyJSr002UWhUx0MlWzbGVu1he/qVqGMQaQsegQUvdJbrdF7yjQCiz8FY
FXSMizy+VB5RdA7+mq5aV985hY3m7GGyo+ywqE7bE37mnPaBIf2pThpWdYp2QIXCn6yjMYODU62g
ugQkXJHuiJtAnBiggHujZBkctlVoWHylaO1jJlLNq5DF8qn5Fr3dHvryBjSyLWmnBTq8G6/KdVqw
NyqI/BmLbDjIRTbo0kWJO9VdtsxyT2nDU21a8Sm233Khaj63FQaQmeIBPUrPLpBnfCfAO5G8+ufu
/xs60EdpU7+dbO2WAl9DU+TCf9dVkX5/ctykTjSk0EF0gy+mvJqK2AnSaqCKSqg23gNPlGCkg8/j
4PDOf9fj/yGWbcHL2L+GeDPHWsXxRDzoqoawmbiCcI4g46GBtNxEfUN7bY0G4s+DVBNanNciSWME
DhrR6JMhTPy1JLZwbQBoN0l8gi9UJ72c5akwjZifORSpXZ5At6fzNKTAp750F+yX18YRMKHLwt45
Fi1J1Y95GtsCr+tQzPXbOO+39cToNC3dUuDJpWxpfxUhqnq2xsJMsGc9bUfixAm+2t3D7PYaVfeJ
CP4Rhi0nkiYeOO2ysRUxO7lT5LsW+KyUy7oge4jpaS1tIwfsO2c25lV/V5gFjNTkLiqpjJzsD/cs
mAFb22MmYSqSg2Dl92lKheDmP/C90SZ5SEHuCjMhng287JTylQxABk5QMNIEtFm3of3ivTQOdkI5
+Uvmqv4EwZMcxL7SEE5yhD2xKidT+OFftqeYxdICXPkrhGzZ57B5ZWQdq4EL72U8rezl7VbnZPSf
B/9roe/bpNsoeh6QUz3La+Q/Smck97J+wacSPn+Uq7KzaMrDQqho5DJJ2wvre3ave2+FP2IS7iq6
CiufWFIj0mYEZroDpp9BaAWWfqn42pgas50ZLDfZGSSPdHEZa2kAUH1k7mLqDS0upGO7QLFoGJXL
KPEWW4QRlUCkdPmo0zfoFD+smPmgFTpJ2fTYjJ0YQmswApowFX9WwY3jf1a7quIIolBteEXJlWZK
Iad51guHVH5vesTDJwmpfyy8/y3AwjgxM8+u0CQ7MDzNlNyy/zAXwF1gmWDSww7id0EMUYEOtg5F
QqAxYNqJL4GtsEcRTYmsTNBrVPeCrLVRGw+h6TMnhTl3/fcpCZjH/t3HBiEvchWVT58yKPVdpPLh
2XDcu96NfvGLefr4f4NfA00y2mdfgAJgz8mTRoXiIxUmGTcnojDosTrHaxBXd5TclCQ3W9KBBxU5
u4GnXEY/qacaSPTxbWbARHbZUtECzbqZQZCyH5E9Uly4h0iZHUuBBf3tM8aKafdZXIadbcAI/fxP
iw36QkZyeKAWpv4gPJk3VsV0qyngDbXRiWvwEacwOUQz2GBYhMBSQAxBi1PyX8JPgWws3oXdsM2p
3NgyuIIKrmO4Zdy8mlpICi/YaaPmS3DkfLT93o1Skfp9kLlfjOHRyJou1Mrf97T2uGkbLwaVcioL
Ha3fe/iCNOXcnD11UORXnZ42fcMNV/CIi2/IA0uj6EwsGCHta9jRvw+VVCQH+ej/pnpHtBJKdrpT
+IchT1CkOkbyq8KCH269MdY65c6B7ooCi7suI5xdD/drR9Ia1oAYNAx/L/2gymo2YWTNZJbyVEXI
Z17xDwx/23RDIgKnPi28YEfO8o8DwuRiuxymVoz5BRKEy/M6RMlKcDqVUo8uRC4JIEVlPXTHJ4/e
Jx1eWeG6lFs7O6YcJURFuByem60nGW0fbqmyfc48buSGBGLV80XDvrIaI+Vu+qs6+7HHFuf924Iz
TF5qQdS9uhyFZP3nOsDWioooeWenNAhaOr71fVC2hstaZjUOR7sUU9dYapS9PHay6fY4yc3yIxv1
604m8eH0n9WYgk8yF/z0p1VVvLQ5fj6CPycyTL4qU7sGwYIOyj+KMdfV/027fx0jSCHKFpAeCN7p
NrkJbukvmzBYmjvtj2q0ZMYi6NBz5maaGN5AX6Gb2Ke1kqZLhVZu7QlkVX9rlUfEz3R3qbWq5cZt
lOO5RURQLvL9B01n4aR9ZqQMUop2CAM2B/nq5VdiSAVyrUIIm8IWZ9pN7qfB+zWDAaeWtRvi9kEy
AmYgIEtxTk/Jtk2wZVA6KcOCOYtGah+0YmPJszkGPpAJF8f1P5/PLR7Gw2gMJQ84r7v8vld39m7t
PbbQlmVg2seoNZNaOKC6QzHn9GF5fEs+UhvE56/G38U7bBtLTJ1PR4PxxlDvONSgznNXl8SzprMn
zlDyJx5K3QWhlSqrkMkH/tyiGI3jy3TM+s24gAP712cRWGw7FWXgVRStre8eCOUEm7HLNyhxzHfW
grayhmjEI3AMTvW+ycyuf+mVEdWwK9iGiuTxVgbJwoJCNsRMp+itt7cTbJpUL31y343Rr2F3uxDu
yANHGsAQkudvAX18J654e3Lo69g4AOS3TKoatnweo6p8meJZjAFN5zn9CD3QrO8fNMNUy1Of0N+O
H820u6mmYYy8tbwZ7AwLEpFO3WQY+ZgFD0B/fbKlyVxql8zQAgFunXMYNmPmGLKZrH6WWktx8MlK
F9MGGi/CJfF+N4j9dmNBd09/lAp7zbsKDaD2LCDt3OTRqAXysBb+VAkUu7KhFZnqJhgiKZdGMu1a
z7H0/bB2+dxUdaZ5XRpswRCvOSa7tmnaTjGfPSxRQFDPOdScrrWXI6xb7IjirFZqKSipESQAVCI1
sA1Nkt/UB2SxIShZQCeAo3pWhvkgMNBn3vzuhB/MPQxbMFiZfNnD2wdCmx4ftRa9u7BTnG8BvlLe
gqudNJ54Us7/ezraTFaIgMw+r4+dQsEgiOU+21EDvvc+4mFwdRp1jhn0d88ffPnzK2ukGksSAPo5
tuB0lNCVaTd21VZ9iwXXxDamozIws1w+7ctDU4FjSF4PUmrua/Goj4qM1X/f7jsQAjC4hg+g7HOB
aP9zexjgq5UmcMpLRCcPVAdkp57rXY1ECjF9LDV7DLI6PIFcuuCWSxLuZcaETzukfTaEDadX8CJM
cqqsZfKesyzMQBOtRe1omHoehXJ2qihusn/bKXe3SpQkIdLMW0vuo8XFGnLaZllxlgEMW8N69jdr
c9iON0tisC2mwTFC9x0NSljDDLElCaMFf/0B03Y17Lmh3QBsOVtTROrglLbtnZaFUOEL+fNUADGG
vQrEQvIxYwmfa2huiI5cAUd/KmZkvOFILJIUo10Bw87seNHu6M18raaGw3uRDELN+qPc94nYm2kS
h7XGQy+N6g+uNKb8i5eKAFRNR/EYmnCz+ho3H8gR11K5BBKoT9jjd+SB5IePjMk9EqcIJZsZT3gq
w3eD+0Z7RhCOLQv4iLMcaEqIc4vt5m13dTfGGLQ/wYROPeTUkdGqE0JIdLovYZaVb6oq0q2leGY4
Haab+yFCkvJ63JciPdPUnT5l/zcDqaNeijrYUBa+8vMsQxsTcqEWruiDh6huPVV5gglr8qx9Cska
/YM3/pD/u8XaJX4Vfr93d89IVI8iysUvwuhQWaXBFkWE7AsrqZBkvj9Vp70wZmg6fz1olC2lpgJ5
arAr3TTAaVX8UMVL+4Ls5WsL8GRGuPKxpt6xvuh/UIstMW3axiWEMqmm2nNj9t9XWZhsl6ts1iYB
y94g2AtvZcyjnlegmxZUL9uSqi03/m1Yp1QnGTOHbgxyZ0KpRaigi9E/DDdvEQdMWyL2cNn35LE9
ZMy0xoZMA828OP/F8dkXGeWI57UAwvoeSD2r6vEXH5sHmc+rVBDhB8xDBJNe1XrnPzPq4DvteXPZ
O+UCQgc13bsM21L9NS6OzFDMnioDjWC5dh3VWjUEraO34PRQQxuM74mMMobQ4hLFfm0HfIArQRHx
K+1g7cTP/Fa5IPyJRDHgUuMl8FwuYckEE86FnleQ/pQdaRUvHQKi9PyoK+qpW9Sww/LOCB941MDA
glkKbWQAGz1uLfEmOI50VJ3q7/055mpjtbkCq/9yS01msgXkt0QeSYeMb9BsAULvd4FA5vC9T7lM
mojnd9bpOQPlTDOLROjeapQKKnE+0jJ19ySKsqmk6gyPqWIMG09dgoj6VwqdEXu7gW/SDOlYX1Or
IaX/Fg1YtBEFzEoWBR/wlQ9E1TvH6Wi6YIDNIoFw77KNhH2CJU3RFx8QnR+7+O3yZXZ5ZCP3sFrB
bE6pjLTJjtuB+40HN2RtaMSU9oUw1LpE7ZlRMHzLtweKMCs8cwU7MnXTHijsRFMjiZB5fbWs8M/f
x50o5N085fLlVY3SqBTcpwrV0zYIEeb1+nlJCseFu6HyDPCGiizXsQu6Yia19W05cdgdy8YkbIBf
ShhuKmcWEDYvTff+Y61eo91aBVtsYrWU95b7VTDDVRs39kR/8ll0zc/HkOloFbIboqonRVqdPoBp
MrxeNaDn/dlnjkdEw5nMqdTrlIdI2oi8kPcLVcq658PeUFhs85qFG6r9fp0rI3Jy4XZLAsbi5b1i
Ryq9VIo2nKd1qoTcD5wtaRgu8gwhvdqZPgpYOuWpMiA+NXnNd7h8jDmg7RlawHUEpGP1D3QPD2V0
W4zamaXDOaNr3rXKw63ITloRD+yaKpNRjCLT/aM+rEpJJYCJEb340l3PePGR+Lr+fHEiuxKZ4hMW
N9Or23VOYyXk6f7P0HR+QVj2+L9hlkg/07YjBvHAyZOV191c5e7UQ8EMyvrBVIhojMrWp8/3di1F
1bEjPfOKwqmlREPebYFwdSRHkA60zkzLImcjllHeLW86g+teagykJs49zhl5gQa6d//4XU5YhSn8
uxyHRiWlL/886UfqWuqKYqr5vTt0UwbhC0PllRN6OxrxkZSIFu3xf/Z2eTOhp7iVXaiTwHbWZwcE
vwEZpg83JP4ZeDwP3sOl+t1I+SxEEuSbZ3IckDYvyv0thHy39NgAugw5IAoDf6aavx8kcL2OKe3A
6F+VxdlwK2FxZiUM+WdiMZb0FPAVeWRb5zoPhrOyFd08uKy3MpCIH09G42vrSgrbrfI95VLx8Yqh
3dhK9cLmM9LPh0gXBJqAMTgLkprW/4/e90Py+pWUg5v2cxnKsSSwzkntXGVy0Z4J/+FeGjhljwU1
uIjb3ILyGCmq3vqJxor4bAxFbxJNl0Rr4byzjXcAUWuDe1P26aMwfO3SlGzS3X14jZ75s4b5RaHs
+mGp0Ss4aDTIkKkapY6A90rW9f1NHtfGEHdP2842NB9t+np8+2x0nTvWkOc9NiCFm/nMZaeHtn/X
FWo82RWDLxkNkIV6uOqmyfiVNmKMMX8Hq5c4I2PLCSF7/Rmmur1RNMVDbRVuCje0nnrUs2YxGw8r
MeaOtOAB2PDDmyzRwbTp8zIN8nqRz812MhLZzlZFueKJg6BUXvsTX4bsBnBrEp9b7e+MlLFHabc5
HK0P9WrRPV1TzDVXuzofMYAvKC7y54/c/mhYTkgERi+PVYvXS6XVscf1FXxN+3N2bM2Y1FNdnqKK
PX9WYhb1LV24GZFimW+yeFNvdlmpPZTwj2HV4npfsDpGFzaBrT63LUg3W9QV9l3x2/5w18fZ5qup
1hPAYV6CoCEAtvMlvFXYZsOlCpLilg5ZReZPiHiIXiWEXwDcYBRUcCR7x2WOsvVFU9meqF9InXov
FEbMcHFeaTA/esirId0KZH+HDscgXfAY+TroSo2OoSSbP96Eyp4K9+v6DCjoea4jPrG2qxjlyOo/
rTiVmFgr0cFygVvMI2EIyJLHkdq2jmW0oQ7CnPQP9mYqISeU9PMvWlCpNaYVFiAqNOgFVo5/MErL
E4+ppOdiwG648rLkbJkFvPjGAjRiudbYikA+KTe2bN9s73SAtGTqKPEVgyyQXU8LCpX1SgfaBe81
fXY0wMHyirTWuDE16M8UDhS/fYIX3oIIjYmL7qiSS/kE1Cnu1L9iyFtpFZ7PFTGWqZqvMFfRdPNB
PE6AVQ4qZ0G8wCJy42LfxgUlD3X+lLZe8Mmyw42WlIIfjhivjJlzQ32nKv/pCN1IqLG3S4PUq2x4
AsdF4/0jG0mnCWowxxJp8vmXVDclKsEvYuK+a+viNb8VyeeUzFrzygX2r6VEwcNZ3fdVGaMIhQWu
h90El9l7u/aBhAL7jxVqEr4i2m+eefslnY15EbOEPMRvpnpiL13lxf1Ftg9B/GIoYYRE1467OuT0
SE0asswfiupN7XtmlMRZMNyCylfqVKZGq1CaAgpNcGmRWfc7DawhyN1Cdax4Revqf9sfor2wyafg
wGIjNyyeGH0PTbOfrxv6KYdcoQQb5xP3DLp5s1APfmU3MnEsqkymhO8zOHzpZAn34+cXuhLCrYbm
AmhPQ7rkHza7/3YZF6l3iW8BmycRHRRuCsP4JQtPhmxAiicidkSm7Mys3KS99P7d9Gygp2UmSdiP
AwaBmdkcZ1mbqL+tiWcQEU0KuWH9hQodcu6LpTdC998lIet9zKSD+AsaLwosHbOvCKQqtAadf9NV
X2yp3M+FeEubLrnEbs+T8lorTFflMc6/GMn7cxVC0Sqp53Te/ZFHehFBDm3ZXiyN3ujSRKHhwkmI
e64GDPYC+hjy/0qItpPtGeGtKk9BAeJn50pQy9bihuerYdk/JtB+EW1xc1zAdQrwbTQvWMsRcpD5
XVJJiTWnHdpmC4Tu2WVZTqtInFdv/0SzMHDmMzHQaLEed7fEFGc6yo04IH270qBjEnuQIz6pxZVI
rcfspmYlqRDFZJ7/HtX7TA4n+eUPAu0npl4+bT5lGZ1EfZxVeT61P+dP5uQhSUD4m+BhZ+tctQij
Uqo1wVk02kjxOFbXe7GpcqwIDy1csw0DxtzcNXCvbKVDO1z8eupf7Qd00X5SiIqpgK6pnyjer9Tw
d3UOng997ndKzyqfqaQB6WvlJtRZlzAdZNydipsEDQE/Znq2iyvAlNPnkyN6tBbz07j/Z9ou0Eq3
lRwMPd60xQYIgJ3WjEmBCiuqBm9rp10LADhorp9l7+UoSrn/K+uwobNE6fEquKrKWt1mc43/l8B2
Nrkve2T4uXkXkC+23txnaqgqEThaNIGckpkzHnSrNWeruyNJ84tj5sBs24B1VYOp2iTNU3LPvjEi
0Wd+SSQJb3Fcn/nxfv0BaKRkRQwMTJkZkA7YZDBBzMts4WKQA3jzgCGRpYFOEOzq/gADbGONI1CZ
liGNGgGBlTHJPzW8Ono5RLFw6Wy7Js2M1BouV5CGPYefLX9H5mx7ffFV+3IvfkMUJo32UEA0JbXD
05/DlBGEcjkqZD5pUpf4lkrOVND+zVq5nsSgYqb6iWQDKff5/cpv9+8WYPsCR8CIVL4Wd2hNpRC7
d98Mmm5q8K3NhYZ/sGNtrZJC40tuFLSHfz6OqezjfkyeGIm1iYLMIY9z/1UsKmaXLeBxwAgDvyzl
lZJRazMP/Xq7bThSrWAgwfBkSySVlwClFSEqmPzJMucLRQYkz+atnNIp86d+Wmn61SgOffkuAKOi
jKcFRRYZhCJuu0f4FohMpWxjSXbMG1/JMKtZMYfJwnqk7l6VHaqZCTgfirp2XqWxhD4Vu2+c1HYD
RUe4zUpubXeIhRH/7TwmJg5e3MX38SOnYoaDjPlI5uorwbihGa7iJTVAv2SuLpIj3sRh+LVHTHbE
vpylJo1uawIP4F6jDx3h3X7mz8eYSigITW+VWLbaI0pGSU00vrWJ00smXALStA2pJJZJm1+IHSWz
z73W2ESmpur6+BuiWdr9nJ8uLhsTvz9ipYsFYLSlg9rE7z+7dFAVUhl2hfZ5W/NgsWNfmSa58eg4
i1zlnhR/OE5BXHPRGt+9hTl9X1XyzgkVGZVY02Tt79FZQsqc6ZGQTZMbBi6r4IKQer7ypEoLrul2
9CXnPIbZG5JxgKe98OcVNfhfsiUZUGoArg7zG17191fKIqQshUHfNeshIPmPdc3MCDY2eCjMDAxA
QFM+hYy2djl4CtXEpQu2kAEvoUCtfdk4zMN+ZX8Tq5t2wyqPcjCIIRcfxrgiSRJ7KoODwHpCA8qv
milgaj9zSuONtyx4Khl8B6wBps7p8q3u1mL2FczDxlkQXDtzGVTyDxDMH0Y2MgUu7XRyq0c87xOs
fwYwDQeLDzmY4ugrNzkkargOpLkN+DP6wp/ZMNGmYy3s6OiybgZebW1c9kmGsJCsvCKpVmDlbQ+O
kku9QWYdIneTfH+MK/apYzVu8m+s2zitQUtqmqNdLS559cwHAPqsJDdlGOHTC2RqnT0DVKfiwQDO
gL11eaDc4rUPLbMIQ80zZRA2yklbKAbsami/967aGt+6TCERfJB5BNUM9YhEF+LSUhjftHAfSNc+
WCp6jnJuYwWLkdd6mAI1MKWhQT9v279LcCOmRuA19e2hcMXNf+oxjRdMocxivPl+ipJEA0Z6bKW1
ltkdT2DGw+FwK64N5cT6FrpeIjtiZfBg/uMkKcZdNWX3/Ol+fRX6OYT8heDTs7yx3cZICQx9lFLl
fhfilMJqlY6oLHSqOnU0uRT9Rhbjy/K6p3l42zxpTB4kJLARGcYmPr1A1QRu/6nC9guspJh9b9mi
/yW6cGI1WGG2dnV4THY2bmcZTCzoAVqyk8L9V10Zd619T/q25Jm6IQpWT/Cb7DgKYJqEjJ9U842x
zIpHpzT2UO0ESZ4H7WBK037mZtJ9SafI6bEEjHX+MBpymKEzM04jyBvkvvFoRgkFkbVLOvDccZYe
2xU68Uqt+YqYRKF8C1X37K9FWDOTNfkoULQqTEoa6unM3f5jLREUSwegnl9YEBxsATlfAKT9Cwkf
LNL/z/f0lvVh3m0rsOrpvhAhJ6enJvKLP/4oSj44U2CeW+cd+lWa8uxvfH7HY8aoit1mQcdTxRsN
fHuxabyrppqOeVlb/ZXKbTIvuyPiyIZ9Kn7y2DwGWnlu5cx/63IDrVXIhltzFBt1nJgi/vA8LFGP
QvErRuARRDdfMUhnP238lOgGIFRNz4/TZIkoDa3sMeX4MoSbClSWh1Qx4kqmKDpDcNvMMEN8YjMo
yqfoQtUNOfpiIuCEawzwb74llKfD9kf8j/FeoLPTPn74tyM348NlfJcFpPeF7/vxpA/+44EHqHez
/R5xkdV24oKZjwX0vMRKnSsSXL50tOoCYJ1uJhv+67qa+l42FnwO4djObcuTn5Xat1zruj2DKKZ7
B/ND0X4yFBbrnOLgW07w04+53sa4lh8z8a4MKcGPqMXVntVyi3YpFFfPQgrMx3bP1dwoTFa0NvIk
FoQNfAGkZ0HJQtjrdgm6yeV/I7VsAyL7d0KOxXfy1rodsbC0HY8Qa6QShgTNvXNHIclOvBA5X/2h
4hg8P15wwR1Ce3WTK602d/qT/caeIKcmkuVMjiJ6h8fjKJ25arROZquqcSdOIQ0wz6mYkgaRexl2
gO0TiUuRPCFQfWKw00ZKLuS4wGYMnDO1Tgz9gjNYFzc9NyXCamazBd+mPJN1JMAxIFVnhr0Pudbo
Sm9I8+J+zU9bhV8TMVWQCacWWfAggvne1W3NWhxjoNp1ZDJOMixRDsQaiigNedTHQteC2ORTQp6Y
Lx0AtAFiPPUNncH9sjaFfqbefd2MKYSiXUStryTH0pWmOwBvTtieZXFn896x1jM5ka0DGs/9QPhr
XqVdWCm84kF8BTRqKfdnOenA7eOcI/dY87Pm8uVcNs+WCmwNilnOGWItg9nCc+gopd344Anx7eFs
AOcpVKetS8N/uuf/0agXmqa/FiatFkhPLDWR8myjOne4LTbOpfJNZK9LWZkxvOJNnU3jv+7xUsTq
himWHQrK0oIOPrIM5/XIxnOAT1IjZezVYt/ujxch3wSuFf4GXYqfbihRIg/qCw0nBQ+f24s7V4R6
59YsynSSmxpI1bJ3BQ6xe68cY+aHlsZrUqw1DUlCUO2PnukFY8jKNdyIWEK2v3AW9jjFs77PfaCH
tujXvKkJFFkh9AfjR18VSQePQ31Mjl8l7MhLOuDzAV91dvuhdpc8hqQX/mR2PGwem2H3K5xEFP9f
KV9301kl2cwd4jmBJ9ndgIfIw5s3OlU6gi2123zF+BxO2/e6cb8d3jY5dEeyvIML3qCu1t2Uwqxw
GUDTz/rClRXtnD+V8LVlfVbMuCxmqtjKWlMk8FmzY5aYFGb65GoKgw36tnjld1gxLI/Y088xPUl4
tHL2SuMNwVZbQtaYvlPVqa4bg3s2B7X3SganJOdDvNpPGWxyoBbp8iMUIgQWZ8YKNzXPM1DIu71X
GxFfaWioqXhWyyKEd3+pZ64epTW6Ng3LvanBmDR+aMwtX/h9YrrITN49kd7hMgbFi6hAJLNVLHw3
Iyzie0wsCGVpWF6mwQNOQzdeDvDeASYxQZuFDf9cXLLep7FvXo94pIQM7QzCejyI1V8GDuGjWT6G
AEnK+9wu/43vHls+7D2ILXL5KHpTixQHuL9VKtpK2kSLGlW7PfDo8IInLipXDcb7ParL3RfZ+H5S
2MLXtshUveo2PKceVI752Nxxu70S/Q6yknrdogizNh1In8+KatqaNaZC5TBatdjBkHyVeWC5ffh/
5x4TYLTOaUmkAarc/0GPYB6PcMv0zHLODk9lmVywJpkFKpjHDaE6YkdohKaxmqa/sbysWPVV1YWm
4z5W/49tcW3RvKkIIcQfqWkbdZwKccpPZ88pCqwikA95rQppq7ZGx/hGs1E4NUj0sBD/lFz5dJVx
d2ah18LAvXX1uIqZVpWbAh83BXinSwn0REUB0gg6hyMPskcEiPMruotEf6Pgbpr0hrMm/8Jgh+r+
KwwtEqDE9Nz42u3L0k3vf2b7YQH1OPw/3i4C3XndT9hYiDfe/87YuE68MtcFvynki4aT2eM4nF8a
tG4zihSKbqwjS/PZB1fPNLYdlBhbkHuS241pdvVPhLWE8CH3pkb1qcAR+nt1fnDCmPFAC4Taes6X
5wXFgilkXwpdDkCL4AAYw+4WlVQIKA/X/ayH/YDSSt4TBLM1aUw9KyGjdxQRICnlIDZF17Lmrwyz
yS8HoSfsG2QmKRbj6trkqVcIGB+KOrVpDqH5D259s03ir+AfxeOoYKqzHwWXzDS0bMmNuuiPyzWi
Okw+1PAVXz5Pg74hkBhkL6ffxSr8XYJU5vA7ddId3hukE3r2d34o/e9bSf6g6Voae61qAd/uU8GS
xl+H7q6Piojd0OcD/rZ+lvlVokZNBF3CsK12U/32E7D8eiGXdgP4lkYMDlAdPk+iITRoqR5XxwXb
FvL+DKywG3a8flrplUZOUW8ehdrFEFhlVNPg0TLrwBHAtNavcozVy78l/YzHTfCyV0Vc17RGrdim
oXNpH3+ynUlo8+FqGFP782+JzQHgybkOonsSRnc38/ZO57xfAYif2H5ZwtoxkbN/ooBrwfv9Zke5
p4KvZk5lNS+dD90+1EzfQ3p+3Zj90LiU+NUDUWMfPBBXp/PvlXQyv93fS+v5qqZfZwTlezjKoSq1
Lk0/v9R4rC6YT1gktaMH1T5OBVn4TvJ/anJyhQrduXLSqMu2+QfxPA+BvvPtq7YpUSuPN+YCfjWf
LHoKo3NhIqQQX5LcisMfrC3ae6/hJNedrO/GpQkdCavNGhgqUtgRItbQZ9hyAEz0+RuF/ANZrayx
40jW+q7jE1NOI9bFZMA1wKaTT0hT+zi+HF6sU4hjwXX5HS/OrqoypjQ1SQjzcYmvLbdldSjqTW1A
br35CHKshH9JM98GNaQEvTGmSa6+Z1if0aP/dyIM8hIuNVORzL7n5nT6pvDgAM4ELRsSoguiReqQ
gn8+HjoAqmAQC7pJMTSPqnLZ7InL30eZevZKNZl8ao6mRz71B0wPdwyH4Ftjg4IuM/YJHfyDj+0V
iJ170zvknbIqCwW/DJ9guycnD41a6JdwH1ADeSfXE8D9G5s/IqQ8izCg6IHpoDEk8RVnXzaI1K+U
m6HmKS+raZxYr1agPgk7BPYBeBeswlIW4HI+aR0FS21+9zRk78ALZCg3s+jRiujOnRyTNNzSjt/9
p8oIMKQmV4TtCmFLbWGUme/sgb3onIUNhFvi8PSzTgedbPxiiQwomGhj0ESKty+kT2TxZSNMPhGw
Ce/HxTXMyzNwshg005RT3IW2Gbwv7xLMO36BlANKXn0QKGq8lbLa3Ks+zPYpFOIHjp4XhRCzR2uf
YfbWHKuPeSbFN8cSk7CL/HRD16XuO/1mvkUNxs+wfqx7gs6Ts4SS+joptA8xfsv0+ek9ek4oXa79
0NhdQZbvxcUKrPoT1M+supi2OY8MUiO/03w/Ws93Gvud0OBDORTBcHtxFgdPc2iYTi4mP9VJ3AS3
YKHi3Xfi1bRynANuJeVuYskOSYW+QPsnGmOTuwlNeMaDcCvA+qqS8813mlxzew+5DTBU0KpQLM1h
9Jslj/Q7LcyJoP4SpWjlWSuoipcQFS20Mwhmymx/w2C2sSaJeshpTQtCE85AKPPwjufylXY3m9ZG
kWiNGk86qhmspKibaSlM1jFXXhajl9NcyH6niZd0aO/drcTgM3qXFGJxOKzvzRpRMKsnNAR0IB/z
QoSt//7THvoqkpjR6Q2WnMquJxqz9+ETNK8JS7s/CXcOfaIjpNdXR54tV1jJqC78jX5+D8vRpexO
IZjh/W7s88VEPyL/vS3fkD+R5foPH3rfNnSfa8zmlaQDJKU15UkbVwYm9fESKo+kLsQw++wfRPeV
oMAkEmJfejsR4J4SEl03WgNwxDEomjYH7z1/UwSnTfYp1Sjzd6JBfvDQ5MgZNuWvZNK4M4EQLSf3
m1uX3uHIfHjiDWcHEHgeRmRD9DSvWk4g3UB4M0Lso7UKZPVBrFJGjO6sAn/J803966AWEftiOoHr
Qs9NRPexdet6uw/G3ld9ntlkxa9gg+4Phe0klD2B7mxfZUblABjHxZLE1qnMrhWTWboESXuZVNIk
TJy6sQjQHgExgJ7paWLJmbAgki9WLQJhWVSnrRNn6LdLXzaWZdGmQudme6rgijZFxXeCy9neXpQt
XnghvaznxoeGRjsLFSk15bI/mi836LZ9ahvKUtiGZOg38a74LKPW42cQhP4cBmOUcFp13HzMFhQc
2b0eSsyMXUS046RRN6DCB86otA5Fcnn20tgURbaqzNLD9MXZTMQTNWRMMjnUG/nzZxeceF+KUoYc
Uzz4a5ZPsV6SSb4tJOrdq41qsXUi2sAnUjTPKV2y0U8HukYq0NY7av0HOITzq1Bg82V0zq+nUPA4
Y7KjAWIdrYIjqwD8dQLfRXQpv2EntIwoUgoJFekPgY69PpBeJq8OjeoFoIoCY52s/VbbhhQBtK3L
G1y31NtEIox0tkCRDLE5pPG4tYxAhvIrLlug5wasIwmh1tXyUQJYUwvZLsIM9JSa9gtulRtC0k3H
X1z5zvfVbhV0cuzWH4A6gJCUiaJ6htLAIsNOWsVGUSdUM/TMqxJefmj30ftt8l4GSAFxdoy2CBWo
XTxLTS2iXBJBpRTy6ZhjyDrv5F/wqUy8/c/OVMcoCWLSzy0EnZK3LkYue8ofJuCcYHsPmuZaBdiW
/SgKpiTdmS7dimzamu3Ypsj4i4gjqxkotvpzzUkZivVe65Ex9pWVCkifNBQrYdyeGv8fGXcxED+6
ZVlk6ezslDJZOlva+Mt2ASpxSmLCjUTiSuAVRuMimlng6eV241fh3aw/ekkNlCt4qr/NdHgcx6Lp
E91EWdgAgrim7Y3C6tpvqF86XLwwCx/RZjzUOctHWhDpy0jalxRdjbRLNuf2Jbx3uJvwBd2A0l/Y
YlIN+1qaviVR8LoFPa/hCUxInzJy4WpDyAAhOBU52oQmJpsdRL7EBAcgF9f1lz1Hm3Kx487j15LN
WFKzsU4un0iywiSycSVhV4FSFDNP5B/wwUK2dwG2I7Y0Tc/mV03xrmfbpGvwJVx/6xzqV4bAtQtP
yMSmCAN6anC4rcGAj46tQl/S7Zxa8X0BI0VGOAqgePWx1c9A8FQU6TZFYu2HXS4yHtaCUo1WMeN9
0aoPPW+0ZhHdEr4bLCX9xFN7nltuBB+DOg0kk7rhU2rs7awn7Lyw6HN3xB3IiL4sdlFD3wzIKrrz
GjPXFkPg5hwDH5Pj6D765UAItiK8G4L/DHCbiEQO0plwy6mv88SdafrvmVD7rYlaZsSggghEEm8O
JvCjpAA5Alqx43D30DNbmh9zSNlJK5yE3QG7FLezJPXZL+gXFLjL9eyw/423FzBMTxPn/aEaRxpv
7B+Nl5jaXJT5CG+L/E7djuEaFVkXHtjlGHvy6EqxVGDw3UJugx/5mlAcrdKAbMtazJqICuHreAtK
3J+QZO1acotV+w7KWXqbppGQvtXb4T9E9S6HQWVeSqst22HEp2Shu/0h+bl5crHIn5dyzT3+kvCC
IP20JA4tLYlUoDfZQPOUYYSaf1Y3h7WNcQrTGO9Nf71u8LwCU8j3I4S6dMzDaMFIYcs1NQgo5GPg
gy5zMncKd0rxAHmzi+DQitH4935ZiwnsTs8TgPK5Y5nVZsv55Xz4imSYGffCzqih3cuLqEnWc7v9
jbihwsp71kNfZn01095jjlFLnlGipo4azZm6lsifaAUOBIPlSK7dDxx88aQprHduiJcTKAILRGXF
omdSfefmV+iZjD7aVEFp920Ga9yANZyj2j4tQMIGzxYTYlXRF6s2frq4Q3W7LXkj1YHcMgRsNirt
bOUDt81nnz42+pWwYpIEEMvk3VtFZmi/IX2+oBX9c9D/hnkDEfaZoapTrN/8LBUJzvrW6X5l2Jog
eQmnzFZHHbqWxOfJE1542WPnxLbwjtxw4E5a2ZWhrMwQIc5tnP6VQbkxpeNj9g5bvbw/Zl0ujDJP
PnRsglDB7HmjG/53+Gj4wj9SO8l5SG7epVoc3QU08gLG/tvIJ6d1O5+NVvrCoNVLemIjBIkaSqJm
ThuAcwaRRfvga/zsGpDbz+7QfSYs2tgWeoe0KZaAoaSVA70UuPh+/wbSZYtuI23b5jTwe1+qHMLr
xA7fIRQymiHVe5T1tz/1PXkVrvERf6iJXu2pzsFxnD4lavP5M0qdoC0Bfn561W3j3mAqwSiGVbct
6wP1wPI3gFEA//2AWZca2yFVyDxbhhVVAbQLuwshL/qaBwaT0+T8CRgVSyJSLTLDJm/f4+pwAZDs
t9pILx3EzqdgI4/hGmTVaviEaAihysdBLSBEhI1OOG4zFFrUuqB4MW0EFQW/+D4MHK/7cW0QaAYh
Hn25vJqp7BWTk7z/5nyEjdY/PoAiP2P6+DDOFDzMS8gnzRxwEyEz8dcP866ceIraVQSi6bZeucTY
lywr+ioufWWWf+9cmA/30NkeAazU3onl7RQUftswAtBATGRH1gTbj5UVVl1u98c7hfH9Th0vI+wG
WTN9JTUiWwmd88fQqk75sp7QTbXdrpwPyPiWWQhY2qGCKQ3uwHdLR1OdXFdZBYoTzn5tH6RRaqoB
3i9bVd3SfCEUwQHS7rgi/U85TS3lBP8FFcYLoNcy6kVRj2k0zOhMUqcccKslJY43s/xVhzC+8ohw
sQrXpkhbQjmrENrxKeKVN1mDC+vW5twNo1rgh7wZ+k1Fn2YYZA2c9nL2cWfYDGSlvvaBSzS0OEHR
K7jXmQFpL8KzOyIVeYMjURyS27zv1PK68MQg7pt4BhMETEFPK4uQ+PIRaIaX2CYhvXOmNhuTRElC
bUimx7dd89r5J7v1k6C7F4jDkciw8ovpuxnsam/sbGmaU3dbca4e8GM1T5PhQL6EsnWgjmiTGVja
It8Dcy/4PWm+SPqyBqknkxCc0JsKogSLpMl67NGt35oUdSL+mWR+bTVy+AJE5lqM8giloGg+tlMM
D4OJDdBr9TuJwyJHh0uDdTXBn/wy2AcQHym1ilaAbQt4PDZ+G/BHlaTi4GK4MFlU4OP2husWZnxx
PmEMQbPCQMBX2r8BHnlwyh+RTgnFw1Na44NGFv9knaFJo1ucjwbYaJ4MTH8CSTeT/b/AaXqfEeiP
FO/Cm/IKwNj2O1j7dEFFCexyu+uxYnUUXsZ3TpGDjHV+uMEmqE8m6lz68bC9W44U9wL+lHr19wte
xGtd6T8UGqJnlGVOYyocougAMFhY5F1SBPcykA8dO9ZmI68XzVhIlptQoObXUdVWZ9Vk16Eetuoh
PvqCWkGdi82zbsxF6l8PIRIi1roMC4qoO/NrBckfh+RT+lCu67uk0EE8IR+EYoBep6XNTZxM9SUK
R0aKu10+P5e2eBnlAo3YBII5XE3X8WbknZQ2+BTYVABj9jboFfPiwujqgOOSf1qcVgP1VROC0Wla
9rcEbk4XFwKlVXSCvAbV8DVmiVir2CPSGlWE928Neojx92dKIzdbA16wq8i/0TiZQCK8yUBip+cf
YbDi64k0NSKGP+WmpleLLhvUEG9TIY9AnmfaMiXQTb9wsOQLqaIwFlQLtUHX7tZSPjJZeKvdWyXQ
EQKa+4CjE7u8eh2OKkhHBsWFQKq6RZVaabsfV9fCKkfQkU1UAbIjo4v9a98jgrLAidtvSQ/RcF22
Voxnwd8/BhMxVl6acj/k/LO8MxcsDhTJLCj41T0G3zOwaRKN5BXZUi93tew98hLu4WWzfscbTyLO
Hw/1ODfeVw3ijwVA850GzNbNWYcFUlEM/374fjIZNr6CdgG+7U+weKX4CnvTmQTKnHEdLEJGaYIM
uHpacQ99tEPo6r9EXNjkWlWV6m4YtDcEk6CSDmG7c678BcHIWjKqEx+DSw8uFDIC1qz2wVvNH+Nu
4ye0io10xn/R4WOj5kaNpXDgcKM6eKGZv84Dwe//SsazZL66/FZpLDjLTFU4KaiOW8qiq8khg3b6
66nbpUgC1L/Vupbxz2MuBSJrK02J1Qj288RNANyEhNMBzLOv+Lr77j+Up3BBTR4vxCdovyaLblou
772rnt7gLVfdCOJZjRLTooTjAq2GQ8G0demXS5G8l43OHagqn1qE8HqZCPyzVvTuzJnbGoaX5uwO
uut9oA+/o7jVdEKurMSHHakA3LEIYsmy25vfCpGD5zlv7OysnCK16H/XZnHmfAUiX9u+y3qVMaIV
DVcE5aZ+0FsX6OZQesebABGXO0c0u5eJRlpnR13ltumGYv8eYMAk4dJUjqtuopTkVCVbAC11hmAn
jMX5YfU9RSYarVZYkv0ymyx6QHcjIKvUPRfGDOlwRr2Qp3Py71DIsn14dpWeFgpS5CLEyHEpBWPy
0fAbqxqXfqLr4X095++KHdEcJKonA3dfSh4rtMzC5+rAcR2/pwgUeqSRq0UENWCUODHnfL3OcR7w
5JVXCDhODTgb1KNUog79VGhyTcTXBXXZkKbTGLVKGyztpSa1PCzDHsPfty2CufkcF8zzPRspD1CO
WioDKBPLON0UZ5gw+y4kFfEgIeoXqkXdgFSz8QtBayrGykWEeLZqsREnxLxvxFKgMMu0zlrrnYj2
DCKWLsxfY3JvgO4HPTlFWrKnSvuluszZCS/zYFlsmC7sQwDrcGuNXSWhEblkXAkbq4axYzunmELm
/GAWmx9nVMZiBlqQLk7BeU6YBqhmyyMhXeXlXCJJrsgyEsBAD+Alb7Qa2Ck2zy1+9BX+WLXQZQUQ
iIq+g2XtBQeExtqZvRlxQGH6i84lwzMl0CH8pTrPKRCDhiFougcfF7eac7dw512eA4obQcpyIvfO
n0/yZEqGkeT9sNfxSi42wlbXNhl9P1rcJLfQtpOkxrKiHg/NlG8T0tRMpSQowjRjgu+jt85dnou+
EpnM0ltqAF69Dqrh9zN6UjuMCcZkoIoP14hKXehgNnO/ItSehGDbGwJtWLHeGw7n3GKpZZwZOvl3
KeLeBIieJWM3VqN2SWXA0SRgDWVuTEgqI5ZyU1MODuB9UDTvJUz8RciqksHpODhmUvFkbLNWZkWt
qhtc2C9VfHOzErmTjY7Qs3NOR9AXZ1X8y+mQjv6cdN/PG8/MeqDGjE5iZBDJl7UB1kiDU9XKicnp
nZvPZ1L+JlW8kRoH8+gUeOlbw9VYlFoxi3IjFLcXbCFHqmNX7C4N4DVVLjnPVU4hUTik3jDLmhih
FpLVWSxk3gG7y30lPH4FA4Qp6IVipaIuG37euQXlVaEtTqQRyXiulokR1rpRw128cS/iFos+Wa3I
H5S4e6Y8+MIGkbUem+Eeea8duh4kKnufcP5Dc9P2Dbh5tL7NPTf3PGmPnKkInE8hh4BGdVvdDzsm
AkBJnchGFA/p+dqJdOZZAGSEsyA72lcoGQ+DVmXlDD+CWVl6atKmdb2ljVMqn1uE1nok4+CI7w/f
hw4BZotJJ1vzs0qaULG0mL40L6mKSGfS58hyAfyKi8R4Rz8mtClYcp0Kzca/R/WHvc4LMrp3/33L
6ojTu1tzYvx4AgrNsV/g3YcGynB+Brp2q2pWBQKlJpAL0PFdl3R896t7rZ7BdwxvDJs+lAjgUs+P
9KLAbq5fLzY6dxp5Ju8V0WUyzqOTdKwMghTl55/OOG9/tFVkImIM6JmqFvYaRUr2GIQ7lClgj70V
F7RsVBFI0KLXYk9UhouS5hp1qRRcof52lwKJqan3aaho459jUUUHnIKBnISytAzC4FmDVHiGo+v2
/1fSRmxliFV0tHKOQ46kwSffjAW+clzp4qIipd1ehaKR4/BtEae5eQNO1lfINO2y09fJMJR87Yg1
4ijRD1ILwryWy3CDSu2hL3vvDasAvdKnKj5cPqb3QX5IH2j7aAe23hAC5lz0d16U2kSqLi5UHJXW
iBwKnIv0KaE+DXneErEgpKRPoGevv5KWhoLvk8VNNWfdOQ/fICUszYtTkkXtklwCC/16m7n3jUSc
Vwsi3bGjnSLNag8Cv8n3oyrQD7q5CrkMlo7I008xQoxaKsp7ZzuuW9b/+Pm/pSmrLzDO01+KZ6zB
E2ZUqtcX2cwlk8W9cN606T2jKZJmaPF3VzAnd7p73WshFAl7V15cR0uQJjSn6wiyqn+Uxnz8Ctxx
U09fqf4Nqt4493AXbJ278zIplElbE0IAk6qHZXHm2u+wcfi/+w6FRMYuEqWonrErYVKaFiweHrg5
94tI4zlRmGnZZUeTgMxVQWFOdoNRcXsiTpfHn2z3x/P3dUZum+DtX51VMdOY+XrX+tGS7RVIAaQS
XcDymiWRioby1E4oaPtPH24feRxziEeAdxd6jPMOO/JuohDO6jqNFj5up5GlYB7c2/N02K5BdMdS
9qALtEzai1oTeIqUu1jDv1VpGtOfczwT6nX+72rdpgW/7DxaOtqxvCtSlTcESuXrq77Yc+mXymui
pU7cr6FxB5b4yPx3XHQwBgeY1+xvsx5W+DUCVBSlqo9njxzzkwQoAsUdNO8DEQDKTjUAFehxjCk0
QROuOgsgxxWDVT9HYCLDSW6j7ZBc/W5CqXU0e71gz/us0ggEVdnd5fTafa1RbfHQL6dDrPyvBzWD
BZ5WH2wi52GBOZjcwvzbUv8kztDafQcCMWhuZjfB+b0gHHC5FgRSEMQCDNAvqJYVd1JVPLup4yR8
zpxYb3hn5heixnFKzB0QSuKStAB7Dn4PvsWDAbSTdcVkUSPrNPwZQTnb9o34UZ/96RCllmOcLTv2
piSHKHLkyWWJt3DFuSwa8Zpq37vjkprPxZLUDEc0XqhZeGGQ+IxYKjO1QWJG5slrPbG8TDsrEmph
FabfUSw7iQ/PNoSkmMZaXW/2oCksyPQP1a7Lb72B8nXh2wSr6osOiqwJqkXsUbCZTwnA3RDwbTrJ
ucEpB74KN0gGCT1KWFExsIcxf7gRPb2fjR/bxgr0F9aLeLzyeSePS120HsSLe5h8pnkHzZSOlV69
1l4kTWJh8w00plONHY1Xgl/Y1HP+23Vj+vhNXZuTjw71NY7l1G54jnQvvhP6FD1Gg6vKHGDYqHIs
a0V/r81ElqfDtVi0I21jWDPEAz34k/tOlHVAE44BIXiwZL5oMwC1hN+ENZ99nsY8mX5CyeDtsXFl
6B6BnYgJAhkSlbQoWNb6dtpyipdpCTnT9mwg9pb3c/KJmR+q+txL7puHLZwqX6ThK70V1eP3Xnle
mKNcgG//RjV0Kxiqf918Ipkoae9K95zbSgKSgBHzsYMrJcJh/Ab7Bkbam/SCGq/eZim0A44+XwQk
fzLc+EoX378HAV2p2FV1XP11RXAln74ZHYxOHjvuhgBTXHlE0CXM+URX9hBkFPzK/soqtXGODFk/
5E3PqTgh5lwBh3TbMVp/blG69XHfAICXewTNNGSylHFIbYEJ3uTGyj2H3frN7nJOnJl3mKKwwUMS
3NfJN6KrmytystdBzeZd30EEe7jRhpdm71m043YRqL2c9R6D8EvOMUsX69s67JnebAYivKMHfCoe
1747UwVT1KSxz6PBN2sLnkn7YgPIxanMRJR6EnlJzDgsT0He8G1lBvS3Q6UjaPrJbaarCLUjti/N
seJO7eMTBokBBKSOqOYSaWN+RkuCY0kJNNJRrhfUef+X4LQbcloknh95J7Dygu57yfUS1aaI/kNS
suWNtAQr8cPBRF6wH2JEr/aqm4ctPg5GFnJNmLqsSXVumQhejX8BGcFSRr8hnYF1dNPUFlqYHMHo
LiUQbwB5RG/FejtoAc+A7TYuW/IUGmyHLSlPY3N4yCmNdR8yYs5p4cZQYzp7+UsJeAkO41wpUx9j
tUelwUYVCV2upuSdUYl/z/3HSsXL5wUhSGtpXyzvJCZNlI/LbT4bw2sQ3IMlV70jdW+CKEK4N2gf
wZxfr5Lk7bIxWIRg9JQUSFuBYEYM8ZR/uqbA6xF9lBWgM3v6+vYTBep3QkYxooj73WtE3jo2y/DB
coY3CGs0UeN6rWN+Hp7vha2v9kQBvV9CfR+vESJCYcPsLfPS2kzIGFw8s9f/Pyyo965csAuXJNTo
eUui8PCBy0GIpI6wvygNXJxH5iohRRW/sNdzWLF/QI+dXB6cx7Xk4MCdUyDlfakcHkQwG9iHEqLk
g+eDkUbbRXVsFT9vLwX4bsTuUB8qCP+OV/Uoil4dVuSUu0cdDw1WT73QvfKrLLYAgXHQv1ukaM5S
5Vu0INL8bJkkjKlItG2X6B2Gxmrh5AB10iCgAwZTixSTCSRRUs9O5rl9c7lUMLMpfldSVl6AyeXT
HrdzaVPdDzukimKrU405Bu7INGhvGFYvh6RltykkoS1mTp9aarWY2QxmWEbpzIlpjPs7rfacEtMQ
ZC480nds6iYco+vUJSRtSeOWu9qYIgoGvnM2UC1no+uHH8DE8FziMEEVdTzVxE9eJCVwsAaCfrSR
Z2oxEyVAREsZauAGEqySTfSRqEx7I7gL2ARtyAQe4xoh2eyzW7q9imiV+WeWlfBNb5ivZB3A66z2
PkxmF0clxYexfthcEM+H77Gy7MjjQJd1wcxffpRQUcE8YsQCHI/YKAn8IfSJQ4qgcgKBo3Wu8G4H
2YLR5aghvzrx0dTnYdzTsCC35Nh3S2lQNv+R62xAc08NrILN7CRKtM81pCDLUnO8dsHuDXvclTXr
cX+e97SsC0ycJiUJ7Zyt1vwL5hgr5Y0i3/Zz0B7w48X+XgG2BwIWUjh4mUkvmhve1wbpiXAiYyn6
QUf5IsngGGq+OPZ4X35JuiKEoraaJA9Po8CDdhBZRCue5MT9v0Z9aPiPG/UaVg56KlB/Xc9nYFvj
oknu3N4gnydifEZg1XbMnKPsRoPug86SzIJRaZpjfFo9IC/JUBrSBrIfX7wgC/T2bSCF7WMXH/Vf
GuoTZFY7bq8ag3IDBasBTbXshgMn7s/cBF8QvyvIxWxqVTtuIeaqNeriu9Esg6jYjub5CvV2CX0y
fBZLO2Qp1NGkOoMuJWum6TQ0eZtNcZBY7rq7OSYdVrhn/lXyqPoiMWyissHLR3RgSCHO3g3JIkyz
OQnyR6wHuhIA9dfQ1lY7yDj7tyGh9nOqUFKPQdh/S5rl+1/IClDDGZB96vGxHlmKa6VXCwMg3yUx
CTj6IUzQ/9mKzkmQ72R3bEw1F85+8YKqCsdVK//ztkVhO2LzOF/P5KvnjTMkYwHFgfh+HgfLKrWn
5bjxAgOV5HZlmbHHxJhR5fVNXonUV/HMRlkmHnbfM69T4q7e7bzm79OqlqUMuhZ3asAbyDcgz1sA
jdnWoLDJYRpwVyhLl7wrEkxINIBn6aAEQKSqtEn9LzmsyT2eqMptKEpWgQOq4eKHeeTGbIrFIWlG
nRlYcS+L15N2IY0AhoxbdiW8kWOi2PU7Qv0wRo3tRsvcvlQ9kAmZ22NMfGDc4FDhqnS5VGvQ7ZZH
udfi0wvW43vzCUS1HBnQ5yc0cqGbyvt+q1adjEfMiDgiS5hQbjM+3Oefx5efJES7/00Rz+llP32z
rXTv5qk1bagWnEbASJDA9A/Vfgaewjpd3ahvOkvwG8zb3ellwHLtiokMJMxXpQ0SSQIcPBhAk4Le
xpx+IGuLCQDbNKOAhC5sHtINMDRQAySSs4aH6r6znJaQ9QunP5UeUT/d4o2BvlV5fTxlv13tkci+
qd3U3p7n016hI5uxxfaO0MrfhyYjRFfXmZ6qKbDpiCBIz5+61w8BtrOChJq9KZp56vG/X9BK+8B1
dZRueJjez9ttToRQ2yCNVS5iq6tbhyW5jrAH2j+1u/h89NgUx1aK1rZjNJyBGW+JfSD7sgXqA2bq
4pENYGs6HFEBN+0fYIZ2Yf5mMFqKqreKlAHf093SjDoe/VcshML3iQFNecPSzpy3IwvSmTiIQ74B
dJRLb06l4llghv7QKrvx7Yvyj0SrMMM5FZ2iOkCnwydIdsWMLBtdEjDaKo4DiF16WH3aI8DqXKBE
xwe5/8zWpIjXWOf+Y2nsKGocIjcuLu5aVQvIXWTeUFfcbnRpHv1tOsC0EmyAApevCTfZNkoqrXnM
sAOM8tnfM45HngO8XuEX1xhLyX56k9j4bE2QDXqQMSZE/BqiAsPXlQbWrqb1dyn5+8Ug6GRQm1Im
dUdYhLdyxVLWea1Df57FoAWU9di+R3BO22Yo2v3B9Jk1TGmUswQLXBkuCD0IAt/KGawpFIYO/1HQ
9O9xJG1BCUOnXl0pPPS5kivsADQ1LVzaFiDCSgdzEK1+g7II+cm85ATHs/b5SHhC12GpK9dSnkK+
rZai4wKreGSh0JkV5K1NygRm4VZShdYL1S/v5yoYS+U+2RYtmnb6SkPlq/DLrX8O+scC3MCxccdZ
rUDJeK/GKUc7zSKvVIMK/lfpa/731zDe5kAu41KGxTiPwo7zcOPrwl6yMIs5W0t8Z/pr1G9ka9U=
`protect end_protected

