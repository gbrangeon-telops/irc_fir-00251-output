

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eddlQ1EVBhLWIw/V3Y4jUv/9vIqrPH4OG//oOzrJzxfxJoDe5AYwYtf4Sd3VIdakKHjGWL10tZxJ
4ECEoEAvaw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eigFAyj6GpLic/D0LIryLMG9xQfLbNW2aTMhx8nk48gxIwiUUV5O0RCi0c3WxlsD0Jm/PNvkmU9f
0bvLBoFrSTxK1CBf237YO6kwoV8FPGCIv6uN0rXS9lJQOPdNh2ZUFAvoavKMegwZ/325WocnFLGE
+YU4kz1iYX1mmK3UsWQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnusdFYP+cjTwVO+sX1Blw6b4HVRZgRv6yA9tZdzqDv0sG/5WALWkeGj2iueXjyR4cWjsJaH1ItC
lJVwVFFXjpYvHwJ5RnZSqxv5F4MQSqH8KyPuaWJ7fxXpna2BJOvJUmLpfNOHHcM9ZtydeUw0FeC9
iaG6qychgs0JvDwxBvcNWeI54FWlrduydqedwrfELAOgz2Hnkk/tLLl8ktgdmAuHiBSlaAN8i7/7
Tmw44CbQzhCNPl2j2hqobn0a27C2ELHJlqNJpm8TlXqvKo4J8RYyFeM9H9JreJ/8JZ5Gf1n3ys2S
lY+Rp2WYXmq0OKzkZyIfymRWl5zSUC9Q8owcqQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uySJstuqi1YIYxsMDiwNUjJcaDIhlVqhon/QnlfUo3RyDfx9K7bIKjrz+E5jMqOrIwDUZDswr81x
cRDaji9FXOgh4P4INZOlQhXe8T+6WB7arsOA8Ipz2w1V2sV1eY1zPj1AXh27lapbQpMmsim+eCnE
1jY1XASKE/xreD8Glkk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l0UqkRkbyGn9mj0GavEkdTUw/Zw8lL7XEPhtCkfsrXvwKb+1KR5+77+E7EhE93Pmbk2awJRlXYwm
D65p2I5aXxW9fMEUNE0pZrhuaqpOOrPdC2bw4gaCcKb2BQm2PHu1PwR+8skPqiaBAqZVoUwFCZE8
LkMHYL9PggokRGZn1pk2O/ghNvl2eJ30v5gmurH3kQ5VEWU71s2ecSWfrCtyS9G29Ke80rPgnbMP
zifmkvX8s5FcVU1LeIe337473lbGtzk/tTh1neIkyiQD0Lkip6Q3stpeftQqI/864FlzKS35OASQ
wgYvGQgHNq1FJbrpROfsgNyTrijicXvjvpG0Gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37152)
`protect data_block
kkk9fIKNxlFOhGpxsNTkUIg15CjYTZ9XAEayLhnhVZs7A125zWMVDdD5Hx+yZD9OPVism92fyVL2
h9rHiql94OshXnke4Iu4wSp/MIJDTGij2oiovgxIDbmNv98/3x3cGc42erpe7ozSPzfVfPKYt4fW
6Qhg0J+6WE9kV7g8D3ui3aELve/IXpVmkXzx7zhIyQE7K1n8AVV2QR6MKh5CRVA9DrlTyOjdgibp
/MCd+knE4L0tO0Awqs+7YWDunm0yJtUzeNPBEIVgsKd9CeN+GvRuHMHqJtlwrNrcp3VlaRVSqM2L
xQBO9EEqKRelzLmkpHZPH4jb6dUoqAA8n4Xpardf19x/pGsHHjt3CjpjWEerdWX0CqH+VH/Dp2ng
IZYyf5JoK4rSKn443ADxLpDoQ8PyiqucguhN+l3vp8UN36s3YBVlQQzzwHnDQ3cLvhVX1AM6Ct9V
7mJ9FUtGQfkR9GHdZVsmfov4oRPhxlkPxCy46qLyLvAer82kKDHiziez/ASyRstL1qyDiWcB6aAW
zdogaQER0QoviVwTjn9aW4FsBepB8B5Gj8MM7dQDHqctSNMH+twrvIr1i3QGIiH0dVg5QZ85wg5s
JgYE0F1BoIrK5EApRQ2m3+LjIFIgvYpu0QOASEap8jXQ+4OcEL5fWdPJV2tK7BLRanxyaJY1TSGb
ie1pY9uljqnkO5hWzGcQlYyYMcyBqe/hVJ0fReo0KAvyPsYX12UtJhDut3Itmm9TYh7e77xASDUE
xC2JAX+rrcdqPUzoh008yGATkDip98B21LXPsXR+sgL3TSokiYitrrhmE11DZpz7h5LmzY7C3CAM
p18uHAgkmBFQT0qDYFWJnwJQLT1G6rNpCnllGUzjHckwxcr83juEvqcoVPYOw0e5PG4HhjXzg79s
S5LqX6XSlgU6iHtSD/2Et9n759FhV9K4jt1/evVJ7NehmbsfveA2HF7u83kpb9ClluEIvAS7UjoM
G5tZ9RDMIv53QlVQT2YDdsR5gnLX+G1hK2tDbUVV1a0yb9UW+RRVo4qp8eDF3OrgNgGcXtYXVqYN
zYW9/7tv13BsI53HBFPLFgUw4XpI6lLu6zLoLHmoCz/zV5aGVos5G+HZMNGgHwl0ki3H6nQEMMIi
6v955MDn9zQDF76gtgNbL1d063UmKnlhiIHDBn99/6Sh3cXmLrRhhGh8pDlw8HzqyCOL1hJjHidQ
k6l9Y2Ajefyc+rUItCaS1olkVvyoXh5dupg/+ZE9B3fC6CxV5+p/1rhhnj2/jR86ZsTIKaNaq0MK
rrrJHOapJTtd2bbeNnRO/iZIqEFnjZwoZda+y2k3Ibc1vRFTrnjf4xiQYlPNDJdKafc8im00vKlp
pFxTkeRQC3MaoiehqOhtNouN+ORhUKouDNu/5ZUQ2GbEwLJFDEP1xvhhJ1QgW/4nSznQ5ZZNH1Vi
fcwh+HM+zRbaZYd8k3YkpwpkcIsdtr8wJHESsblnwXjIxdkGR1Ynh2XkZzEvRn+BAIgk+P+xo+hI
XQ3Uab2BMjTCtEDTNve7byAa/D0BGAJ+RvNGGOXkWHtBlVD4yfBXBEkwZ8CSSDhS6fW/K3yXV4b2
G0KrrClepbtBou+QlMdKcRYOJmvofcybqiy2CphTMUCDxHy7LRapSSGt0rbZIY5BsVVLNurviYOz
Gsl0morLuquUneBm4H4KKHEtBXeFR9dlpK7uNPaKJK7VaRt1sWcssUZm7++mFZt/sIhjkt/nMiUG
GBwaQAE9EIDkXza5qJpTeMHqjsSRZdDheDpg2IP0L7sfc6y8ddMXKZjuKj8YgC5XV5RzRgO6+6JE
lZxNyvuHyOA2OtDcCL4KH9qHYU8F/aVkUKVib0VIPKJF6nAZE60HLu1QliE+39C0oEbX/fpKf4PS
A+wHjHnS7WyfL+/Id/le0+3+oJHj0RUSGJzk/TtkvGLaUqYc4IRtL1mz88AD/kgwBRdvea0u+7kC
7hf4EsFkkag1KUVtJVVb1xAxoyfR0yGEXN/qTSsupTXbufDYYMAugOCD321WpPB7CFHxi3/OK3h6
0KPLvfuf2CzLOo2zZxogMocXO6xnhaCUa7yWQw8qipEzc9mI/JxzQ1jq2xS3f8Uhdmm3k4Daanla
mxMMsJsUuX4hW9/dPWnCq+BFaYwXot7BDvQTLpjM4Q5rwqKkLMqV8Xb3L/KtEo88rEnnWtgsSHoN
SNNpu8XKZOah7O0jnLlTtGfpYtup1hWWfLZ4G3VqEOyhz76w0jimGuPeswXWRZmYmnhZNbJENfqp
Un5d8TyPOQsLvFlqryCi+nwmvTwuuFJ2cfn9H/ntCy2yPSGicIL1aD0C5vtJHCh1sGVjoryMSITw
e0ZkSR9nDGv9MWwnSy5zUdNbOV1KJkrdobv6nMB1RzIGQfdc2IW7nmc1RRkfTXimO1W2gwU1lZBU
bK/9McQsgD5nkPRPqbW8/ruvgm9tDKaqkVsA+HGhYX/9cvhVXzwpT7VN1K8mpugAtIcQSYRpv9BE
hCWFxOba1I7heojoJagtA68x3YyiRhbTNlY/oV29lcfJdhPE1YcQaPX9L9cO1HfgEb3pnCzz+33C
L/rieaimP0tfzV2N30FIF2rpLncI0Qu0Jmcbs3ShvYLcbWRlVDbFs7wxk8IxbyVogSWXRRUAepwk
nUxY9CgK0H/RLpTk5CNpdaWuonoZe5/DYPayJjPvCgQDoh31TW7wEC1X5WLpYzw9C7XybVJb5WlW
oB68ieAWoXOGsREzTc/krNlZjlUze8XsHtWyXKgzWn8/9ybQ6+QKc3A1E8vPKTs2nxNfcIkVu24J
RllyX7qeSL2L3e3zNsWs1/GT6j8aMv7o5r2OwkgTlrLEd6FVt/ZlGmjThrLGzODrqkJIDQq/bOOu
TtYF0wh10BdEquIkaNcNyJ5SCwFJi1BukHmrqzJe3MeHLrhH2AbzE3BvmGwmlU16uJHGXaZBqJ6O
Wk/FdDfTFbSU1dMZYMWfP50BNq/pxmGkPeWVLMqPFkGeHYq9hzwCuzDg5lzIhtd2wX2s4QGDOppC
fLjFGGMOcPuMnnBMuFfAmyODE4IrrFZeUxi4Wz9+0FYum8W5OGCvgoyD+e+lfpHi+dB2nosLN44g
akw6DqYUyJCzYEFJoBmcF3EN/v9D5xagQRBbYz4Q7nnqiJ5npsV6qkZ24Kg5VyQWksuGUejw4iR7
IvgQyPSi4wwIU/lR+ClX6l/KJwtmjb0iluP3m6AlgfNmMAqaQc+gCVaobSM42oF2xk6XUoOXYvti
LPRdGCqy9ppZmblxBUF+Hs1oEYvX/5aZoUy9xfmjS7YEIdpKeKgH+IDp0suZGKMKykv4zH5Asbrl
gUZnaXm2sOEA6Vj3Sujn1P/fxOd+Gwk/XBhYwmWpo1Wo0mSxadzX9CXLIcQQGNYSmkYXHRev7jOA
i6lCo4tw34LTvAkhukWmhcfccgVkWIRzTxlg4WaA16WcmpHLE66ASCy6e1MTMeKrM+f7tS2CoU06
Ur/Kk7Nl/owCh90/1RQTjJx6t+QOPipa6fNxTXi1xOkj4kZAT2w3b07RCBGjWCT+4PLkAtj1e40r
WDIN766x/jZXWvsy5hHk6/PRQ8GFBewgXrgPSPS7sPqe51tRQnEtnuzgQM4UQDyqgmU7UTVj1Nsx
Sy0522+RYLxKTO66D6Lj96Ze8dy44LZBWo5fciuUY9swlJRjY8pokbouRxcR09wCdHwGWfu//nXU
IW4eUQJ0wOXuioJCa8MgipCgH4Wv+YxyLtr/T9+22iFoNXjJW6ofx0jHhWiJc2yuBncpEE7qph8l
cg7QhOd6C5fKp6S8I1qJOl63OXMJQOj8uHy4bNJ+1ziDkruZBXfWKy9TjG6Xs4Bq53D99HrOyqcY
xYMLWjhGkGKSBRYO6EQVTrhq5S4C+o2nqUbx0jwfSzKiN4QR6N0rJT9c1AkgO0yo3WwqHPih5hXr
lpdY7CLyNInOYQPy9FKYMqaPyq2CqS/WrmV3VOUMynZHOxtOKM4yq55NLi0BymKGQxwUCsHSWraM
RYU9b1g+7ZeC/gXPW1CPsm1K93retr0msxtrl/7TnC2scIhmrcdRgxNkCbOQJfWA9aIR0fTHYYpl
Nw6AasIf4fXdgvG26l7Bpdww7ZDdWN36kBSPmR+QDRl80Km3Gk5TYN7hntJDLUYAzw1RbbofRV4K
0/kv0O1kDx952v6LY2WdswR/qSD6Tb/6K/Vr28mDdxA6pEsR4w9UXBNwN0z2W7COHKe52gtRmsmC
GE760IZagx/UwsBWaAyU0s+a5CI5E3EVXtedb4qMgbWbS9wNJZYVFKVCCVnlUw7T11sDzcI0boko
JQtc1hyW8c0jqp4t9aEi5+V/S1q/iX03/HUFwt25+lq/5yef6ykZulzLtGUSUXw+uIIEUX+k3dmX
N2bryMDyPPbfsh5oq2kIn2z3Ms7RrtkDJs9wwBalypQfsSVJ3sQmpD5Auwj3d7o5pDBAXsIERnRO
jq2Np71CaHKDsgJY9yE0l1plM7sXKEz0V4i7kkTDgHtmY+hNe8eaUBNpig3HxzlEnuLhV0c/Utzi
oJzljnaaXU7gErTRCIQusk48J7BsCZcf4muOhxeK62aCCYeTHmCgtYqLCLYJhQZxS8u2C9fuRzQe
cS++ZHOQV444BPrnfXRBqZklI+6ulEelfj4uteFCCXv4SP0BrbVKC0HrfvKv9gS6Q+Km6Wnv9Arq
Y/plevfCwXqe1WDu36Hvg3WpjQ64yUhdPJpdSjbEnDHKREkoNlAxrPPq3kkQc/j/d1Wtgouwfm8w
bsWFPxL5iCComplTz4r6JRmIHFARUdUkhOG/xRzrfA5FSOAjxivji+RgJQwZfUClJOT0TgLqHcv7
mkkHwJiCmjWz+rR3Qr6DhV80coEX9ebT3U/VyuXfHnWrphVSgRQGbMBthBq4P4oD8Pdi+UY6D2gk
WI00h2+FYlFh3YlInvDZoypPoXNdjNznAQaq7JUflPeK5XOkKfv+QXLgaWB74xc06nKA14NIg+D6
IiwAO6PF4NHdTi1Q/52ni2cXitqPo7TXZnS67VxGXcCvgG3PUqc53p1yajCCHTwNDrM5n9k2tKE3
tnHevLaVpXT2mJYFdngAlq33vMlqR42i1ZR2WBx4WmPL/+XTV9K6K6lMDXLnbQDnd3Pos1DrP/Rf
yE6CrdcUa0NqQcm43KinKmM4OnE7/GaPd1WyZGNy9RKA7QK7WqYVNAyITbM034OxAb5D9M+0o5CC
VkGWGzOQR44aqvj2gyu0G3OrKre17MSYI2J5xIPoZ8kCJoqHAnXQKTeU8n0gECbb8L1IEY3BIsFK
q+kmvzgvBNMvsw4ukDePMYi/5CqiuPmXd3mE2a1JHEZDqlLkEcdJBg6ZAg+jBPGTHR+FaNqegxE4
QGfEm4e7wOjOC6bsUk48ejg5x2un7JO9xLg+e93pCQUO8NlTQRAirHFYmWgRi23FR5VOLLWKAqpw
rqxZvIbV8OwarkI2S8H5IJlQ4n4kHTHpDi67VlEXoOdCv53BM+amE9UqLM/UR2JL26b538JjuGiC
bJnY4mSqhapyQbUIKOBccY5Grlp/gZZTa3dgYGiXqaj8aajOdQYrgvP423hNoznA9XPBXY5M2tXh
PiYnBjCJXOHfY/H+PQ3tyS/fnHYMBg1KKy9K/nHX4KINz4671bdbzsj5OIdW4QKG8E8a2c3p09BR
8He5t7L4vqV/mEzjLS/W/g26tNvRN4hqm4AyPA0gAizRd9cJ0/LNde+gjPTcnbrm3sELctZqG9/J
R+pJMdBwBbGwxEmnjPM1F+0SJ3/5VqsPsncSPHu630sK/TMQyKnF25Wy9wwCxGaigclmw7wEl4sO
c/VFgCj/EB4iQ9xhx1bc5GlMHhsyaeeTARVtzHMvCJkovetN3hUjwX6x0cdEYQr/xKu58v1MqgGv
d5Ui2KKo4aK5mc7yNRM3mvQEryvi/UaXiDSpSPHQk0BLb1FtpzWpo+s3MfqzGHLXpmejEnmLlIzr
/UXZ24sh3ZlJwKhG4REtH0qgpq43ZvslrNBwVYt5HjjN7odLPMEw1LBPmAT2+5sBwLs2nyjRDIwn
37CppkB/8jqhQ1sVd+XsoA0IY24c8dHaCxP49dIfINVDHWKBBVOjspvaGr6g59au5aS4oYhd6mAe
w/fET3L1ComeMwBbg7OsgD/PZGlCz2bZnUctIvV+3FGpObkIvh86rZ8Nrpdh32iuu9ad47vrCNuX
51gVd0BsWix13j6xavqgZfugW+V5lVif/5/cCPzTPaMAYYZn4+J/2iPhxver/IjPt8wEAzrbExa4
XR1WlHqBDvgrsFTOAOgQT+pYsMFbfVodLgbGTOjrBkt/KJ7rVP03QOJqXV2JPdngJN0VwW2hd9M/
Lceac4eNoFB49NTVlOcV7d6x0lz7U9F7ghVyTRkE/TqU9NtZTBxpAowG/nPo351MSr2wMuVmNEHL
ErEbq/3W5vMVte1AeEMW80MY3Wk3XoYkCHbiRuhDsDcbreH7eEv5E/AIfXFZDOQqk/frkiZ+4d/F
KwyByDYLZ7uROaEFMp8xYRqg2VbdUfa2VVqDCrB9jX1TD2Vb6xCQfmYhFKxQi2KUxtruyNpJv0fw
68sYA/ySyFvRkZdyyY3BAmtY44zQo9Lx3grsJdFswxwr7VCLpDanE3pZ1gBYiwEmV/s4x0lTLeWb
x0PXdTyjKRkbkiMjE+3lKs47etOXFwkTL8Z7z9Ha6pKCJpyRS875lbY5N91YTBF4B5ZKTmY6EFEA
QUA+7EI6YfTgh1hO0ioxIEbMazbIfzMurK1CT0UFBo+NylttDy/COgUursNeRHsXzkhParmTFwOa
J0cEl3NHEtDc2wsgPLaTPSjbgxWRzsFvdc2OeeCV/ohxdxQIlEHvg1qIvgzPTFDVZ+qJ6W76rnrj
uWxgtR4hUcxhke4ILpzyxBI/ZFXMp0/inoQ5+d4uYakT823X5o9SD4TSxAJFXIArdvOZLeEhCKG+
ZJg3rgbgeZ/uGW8biszUKkrR9AStAnIkY77wDPK4MIG2AJjAZzIybMUqhQjslvrt32ZVtINhAifk
6SS+jycDK1Mhl0ki44x31MIVvF69Antl/eKEo+4GI7pd6F68LS45gueU2PDHLiVk9YLvKjXhcCPr
oDDdr4zVC8K02HnbbjOmGdLZJDL6bK6Ribeo0vI+ZGJQ+HOfR4bPA+PLaRkngsrSBHdzWHs4UMkR
+Tsxzk26QANM0zNcBIF582er4tVMRp+yKhsIFJefVEsvjMX1hGxRUCLZm9dcVmOo2vqMgDFVS2yJ
fUNr7mlkFpFgc1U97TsgvlyjXitHMmC7wM0AABD0GVys/BCEGQq+KtlXUEMfOFm+AiBnSuPhY5kH
QY/divfsv1Jkcwzlh8i/GngalNd49wWWO0Crmol5sD2OeKC6Ys336Fu1sJjVzImFLadJyi4GIylL
n8Dk11ah8lQ8w6CDMCqwrZqQQkfHHK6WSTMtL9pakAqs2+9JSILn7/s7bHSuzvCC00jFwErQhsV6
QboC/ZiXzu5G2reI08mQeePvP3JSq19J1S78yF5UEIqtcgWPM/Pro5eusrriUI54S4Ch7MMj9fro
b3q695yyPyEd3nuBSk0xUl+3mZFbP9T8m3M8EM6zxGVeNbDOinHvMy/1n1LmyAEeGfuTXKWgKUiO
30Cl86PU1Ys0c6uxjNTbanvGO/pHX3fI87AZxwNU/xEn3HVsULvsD8fl46T+w43sj3hlp4sJbj0J
IAPDOH9he4719Mt9ehRfvH+q2a5cydlood1/GEwWRhCg/PfhYhGFaj2dZ+/1xZVt8Phu+zMclS+Z
49C4u5U7vxSYm7qzOBBkacNlR544wQbbCatuQzJ9rimcBdnNGKUq865L0ay7mJdpMu2ri7uM1ZBn
5KN5vOyjrn9BupTQDhN7q+tZVtbQVUwDxoecoHd5EId+ONmk1hwDaqT/GSrBb2NQ7IZxlhZ2SRxF
uPgm8KeJZ8+mgejMEL+BmCxYlEihRrWl9f8w/Wujy8fR8041BUdwmDsiV4aj1paGP8EWigXj9VS6
XPEFom2im9TccX3jL/7n05ksQIYikjSym/qgatOpMhPopiGSR/5a1XxdNWv8CQAkSoF/XssHPjem
nNXBciQDq6KkKR47QvzjOM8EnJsMjlQ6mGo+Tk3G6oWY8IxQZYiwnxF59JMmoJ4GtsavC9KNVs7n
LfrKkkGwChgrPYJIT77Psg4PiPCme0JOyTwlZpGN0zLGz02lVbl8h59GiBNbeOBg+NbYjIvufTqY
C2yNSgFC4NrGPf15Q6GMK3oMouvpDbiRiFmDLfpWyWnufyIQawPtl0ZvfTSIHPGoIqUm8QG66olb
UMObIK7CPYkz/z93gtVeBS5EH+Q5tgUFNILjg6d5N4Ifzhvd9xrB0ghH4+zs3whNtzxC6dMslGKS
U4L7n3Zj3VGRkHHetW1D0DDWhI4U2TyacvGEXUMQHgk3VxZBPph2SEK1hT5QIaG8prVoyQQdCuBD
UP99nstSwtriZw+z77fjIlkPPSXY0DW55n6ih/qIT9vxkn2jFoRJskM0An6U8rP3cuJ+u/0cdFys
ovbZu36dkpxmP/ql9E3DduKfnXSizbOzDP5XHPsUstNHCPq9Lw3t7MF/mxxRhEWkca/v1UKBrKog
lMWvEiV4P9OdJP0l7iHePYzGYAaToJAzQltX2t1qedEqb10Is7TvHrQp8xCo/uc7h42nFW+KvRqI
cKQnP1Dl7WmhUff5Buccm2F/FDDdmgiP9xbROo6WZz9ZNiV8rCcArx7VTU9ez7s/jCeAukcUuADw
lUkQqzcBcQwX23nqgJvpyQFus3W/Lcf+85cFvYTwkNBEOHkRIFFifhTwukVNtIJgX1XPrRCkEjfB
MV8Tu6pMz2LNWuo2sSM9+VNH03vZNJEP+ofVIT2F1f9buNs496Cl6qrPoZVadmveRYAV41XCn/SS
/LsnylE2odAUoMSwExSibaA0pbyg3GxA+k1DTmgdQHCFb0ddPL6hs8n+lEJfI3OoPMYQYGI4a0+i
Rp2z7x123DAAgRx9zkYyR+CdLS2tgAEzmTwM8re/I5EvTLEw9cDFKw3vFgRs3Kdg/lZHmcpD+/UU
Yq+vcnOd5l0+7Bm7cNHoZO52Dh13fFNi2Pv/KlzTarqopMgxsU6GfuE+4anwBGPLyUfjZ7oZ21qo
ehwKueXyT6GSbntwVosyU4iQitSkh/tBmMC/XqtBoAaw4Zl43lqAgD55w9ECpd/ct6KiXdLVshI9
AEaLou/+FU7FIlo9tmrWYhH3XnhgxuW3ddh5DXxP0gnoS1HDPC1AAr2K2QGjbu0qKnn1iJ+Krqw1
5p6ATQnq2g8NMtvIqeF06SzGCqZkNRGItK1+Zvn/b3xUeC2YvT15NpSgZvvleK1lg67I2jOkG+Z3
cnnDYbDsmL8sXlndPcmTYp3e3Q256H2Kv0KR9E0zQdgYLcW69gz4r1NHZPBgu4OG2FYSnJoB9+Nx
mh8Q2VwgqpvflKk6yXr7zdCe2/KXUk20DoMY54vEXm9VQjKUMD7OcKbCYOnkjwebN+0bXM2GwVIF
MEJ/+zXS8epSlWnQV8sEiecBYi38UESMETau95l8KUyQyN23bySStYCImmf4nY2aKlcepq4w/G+O
R3K39YkEUZssdXLkPjqCmt2rt2dK4bFhcaEBSgJWTqpb6i+MbE4lTUp+wKqtZX3PWi8ckhRZUy6t
QG6y04YPZ5ibip16QScXQRmcSLbz/gmN6IkQqEKbfMM0Y9XpzpoZHJLwHTpHl1T3On+Dk8WvoCPU
Wc6DG6CyUzFv2V5vwTzmUmYoCekZ+o6yzoRsE6o1EkdAn9+rbm7/Z+xJ04x0InsHjewPBbRkdhDG
QH0h/DQuN998ZPIxeumK811UfKkSgN5F2Pwq2t2lWwjFWp3QNDNZF6GOiK5iuMto84CtyxXzMMYx
l8GjaoOiKSrAiblkGwEnvaqISiQYJs5TMS+SCWHrXwmnOD/jdAhtLr9Sm2scv+/2CK6G/H5dbGx1
kL80IlrSREhUnyLukpNKmomc7OWWJzh3LO7SUSf0QCiqiBwFPVnv4kGBRShTcTnVBZrRsYbDG/d7
4w6zeOvTqyoJF/SLMcvBUCUSWpEBbTHEt4XmMlNcjzykMqLM+amupGO3xQJVaQ2aC/EIRGRwmp2w
uUE0UIiEmDNrA2NL1i+rk7qJZKnqnk4SfN8moQBQ6ATQLfsI+MJbs2QvfrGRQd8XSCIPeYYaCUEy
1pvNe72rcSdTa4r1mx+h/Dl3S4PNtn0EFQx6fKmWSZ9O8RDyrmL8ZroB1tQVbaxuW1NDCBrv3mB6
mdPSGRvNnasvezRCIvc7q2VLitkaSRUwL2vK9rEihpWg9w/34cF8JbyHTFU3hx99VQ0EVqGFUVqb
Lhh1xqPJbIuFWi93V5y0dz3itQ9uwhD1ngB/gZYNeR76Ycfx5uKQ720YCpaHo22vilYqPspOJY/9
ILkKkK8Rym0Rc/9Vj5SsPgbafX5kzG49w9xD4w2s2p9L0b4/1TqQc0DHwKvKNmkfC4VKI7h66cyi
Gp8FKcUudBp5k1mGS51cNTKnVMuQ7JGkzLNYHskItedg171KyZsxbbLzCkRyVDp4KDX1ir0ANjkh
6wSsRkKtEh0JxkRbtso+ZNo9nLxiroWv4pQubYjxRtD/Gts4Ofs3ChBh5bgt6OY29F4DiQ+A6zh1
uLcIdSEf6Zmb1+WpleoERnaRqquitVEFni1ukq15K96qrFp/aRT8fJzfwtEQZnz2inRcGtvA+mTg
v6QPAM45oSOsH0juYDqP6v6Gc0uCj9yutCoWhAfjPWRVZ/Yp2BTIXYoDu6l2B4PbUtmTiuPedfxN
4LzX9Zfyud8FrZE6eFpO2trIJ2XPVKW/IRPs8oPgZeLBVmwv+dUcWM6xJ99rrWmoV5SDbhD6q2+N
6LkeTqvO1J0ViGCPpoAgIa+219W5RcPWbGMLEvR+NnjtQUdSjGaBonFpQiF3PJ0TMr4Vo7XX63mk
6QCEqKxYzcoHJtcqu47tqUG91E5UXI/q9Nooy6z9+BVgG1ZaM+B7TKkqIWMWeXv4AKpKEfSQHaJ4
bU2aUvQtJTHUpxi2mDHPPbQUVyIlLZ4kbydyP9SxHkwU7gOgTL9oCc7aOHwzfwA3OD0jNyl8sRia
+/FiuRVrcp6+9fUp/hm4W+LlUo/AjkGntSSkmt2PrYfIGM8EFdWghWM/6vY5zQx/ys0t6utICPXd
gn79r/95xNZGHu99FrxZ+fMt27+KRNvcDi9aPVsRwOdINCAziCiyPGeu0sGHLeY4UjnUkxoXKhwm
Wxk+9CxCaVFdujD6+92VCM8qqJThH1M4HbQDTmZWnu/UDMJn9m1h07kVjgtR7bkQcu2Vd8iSHUVi
rbbLcnjlcacyiAKKrs9gPfknfpuvCGBrkUTE72C1eG+h5OJSEHsWpXojUqbITAcEpKXRssBFG2t0
pPvLl8+HJPderLFNCNdrxhDz8WeAcgqZvU9tje5EGdQ48N+HB5Mqg7sDoNjkH5eRFag+anULnssk
VHmdn1geR69ZJS9f9rr6AGRUujQmUxWO0MPLBTAbk3yaHL7MIspcLBRQx59vBkwbj7/6rGks+nqr
FbYf76YFkBQG3KmIpjgC2F6Os9QBF+lEoMBEd2BjCK6xILmwBP+M7MYNjHDqrOkphM96DlLvDTDO
jRhILgOEO32TwdStOgP+z5W0NDOd0RCWsXQtRV4MmCdBguojeD4c9uTD/FnS/eRCr/7GaAebpy8v
Eh/Y/ZenT/4Rk4t42whr6z+E1Y71UqTCg0/YDQ4i+07cyAhcqSrWtfA63DjdAfq8x/sSxRhEIW4d
vbOPvrG6bd1hAYILzx8+1c548qjQN3tZQ8jZix3RRpWa1jox1pHJzutEtPZvyeelFrRB36uIVxZ/
xErJAV/2x9uzbN9CcTqpKJTpVAq8KtY12hWEu35kRy8qWCokAbZVGpaT+U6DdiBLDKpGg9/5rN8X
btrhow7pgp1gAQS1uUlTUVCOyGGg4B6H+Amje8C1RiVjrx2lptdsNUVxn2VRTi0Bl4c2j5PqBdn0
yNqspdZPFus7wO8wibEu1rqh1fjJjBWEQBGUYmX9KQIf5D0msRthLrW52VYu2o4OaLJs5cNhlG1R
I6/VLY/lUT2C/ZLDwNNhjBG+ckTeucCU3JzIJnRJRfvv/LJkVx4aoi2iskslvRjPiCrV+Viwmky4
X/NdtXjs0yzmzJBfYKEEpzXR8cIgXJLY9iFOnWkA8mlT07dM8gG+oQFlj5omlkuujv37xBzmuleC
G9g9nBntJ/wvgQV9gR1vcjP4nU+8lYufglLgsrH7qLzowgqV0DyqQJBpx95dgHDnr8S0XN2ncqBt
jPA3gbfBQ9aQsl3cFHJbxArHr7Skkih78Fg/VDJKYHHfdlrqwdOETDZtV/CDf6HS9wJWcK8ivQjZ
Q3GMvwCcC72lWeSaJspwFfZIQ7GttzI54j5zXGblDCUhUGKgRdWR/V3Lr/W1heTzOATnAJ7Rhr8v
vw76B7wFUa/dRQkgI1lMZCwB3oaeVlOlzNWHHjJ78nZmimfryx0WKMvKXh0/veU964qsliFRpVNQ
/btorp0Y2RrZZYu+f5uuduCmUjE+2FpiBHGkNNZMlk+Q4Wxs0N38xpN/F5NqP3k0ynyzPcdcWw90
tT3tGz9xtZ75WAjXbBaymjlntMAyOdg8MELhNo5WtihYR+eJK2T/ILIgKJ+kp36hjVwWmYYWymuV
NVif/iQWtlVrLbkPfPT8mzPRdZap+eMrTfQ1LhnMYFmKLQikT9T3C0kzjkOmm5S06S4/G5VIekXd
1C3cszYgNhRDA3d3rG4Q1uDn28X5ozza701gTnfMoCPjnmEaPuitCYGHrIJqOAiY94S0JTVF8hmq
dBj7MNANYsAYJND+JFYgFS+VfUTGrJzdqxQFnLGQR4JroDsq5/R/Hd02aFxSXP9VDU4nFkdIATUX
9U0HRI9fapmR+2bcf68E4nATwBcAvOEIYIQ2vHW1Zp74UtwMfr0e0k5sSpVL2FtxPGlGXr+YgSGC
WBBDyn0mpbibbKfC0MR1NIOU4JAeEA1q7FegT9d6dHZgDYgtS4gmji/adaKMtUocpIqb4woaP7gy
7QxbouOGb3fp5tyue6sHTQjqBqVdtG8vQvrogfvIcXY3Qn1kwbcLLkTaLj7+6lx4HXFMM0aXjIbm
aFtSeHkYKhfrj6bLsAkbMiraKzd6rSZ3b7R/f+MTg8cj1cOKMHHxq0dq2SV6ruTw7M+IwqSaWkp7
AACosxBWZ/RM0IV/6GaR/3KrXSoG3F3Tii9anG1rDDul5dkij/6eKNqXLkUySVRq90ucZOtw6oh1
uSP2PHGxxxyhaL+2ZP1GCfv5hd/hdR6ee9F+wnsWfjrsWerRcv/mZq4ykhQkqpgZpGlH5MOIIlt7
rVGk4Z3lhN4rtMm4hFWoEDLA1qsbKI+klDFi4oLI1ouHR0sSxbCETl82BvvRFUYgLQNEE86rIJNP
cQEEm08c9QIzLjZrb+palYhF9kn3djiEHVe7AG1BkBZsLc0taXAUjexUlLuaZTYqJmdx7FGpHyAg
DBJShvpYNeTYTXqo98cpFBpgNKuucK+bnN1ocvMUNQhCj5fabsPm+uTXkmvBGYkBROEIO10/aZuO
jLFNFhkcZPtXxet158vRjhkkXUXL1qbXnYBB0XAAJc+6Kqpb33T0EGQvY6RjsDHVUvvzeDhiYamW
u0/E/coaVwdfIZ4QVjFRYueqqxN0o3t3rhQ8TeXbldBe8cJXViCtvmqIJatl1eIwqhIHykMhpPtO
dkKypdSOnPbVB0rErz46Lifr2EGbEceCGtmvxsALa5gwvuLxUcEpzBCTZGkpY6kuGG7xWyrVfUaE
vLLtHlxxSAYkxLrN7663A9G4RzbhIkseMZZ5OIR8T/k0foz8OGJfE1ITF9re8MlC9lN/x/UGh1qG
jyEJikQWZZQZfn7EzM9rOFCopnWhW5TDd68pIYqe7pCdUgTMh1kQiIdqbL6QHUdOQ+WorcF3A7be
w4JfX6wyK48pW9doZEDXEfxcDkTGnI0rpMq3MVhdiIXejD7HkvA2g08xE1iXmmGXieTaNoMEQ/Ym
KanW0rAjJ8WiGhzVon7uBfCYwoH0KEItPaauJrb29u7y9hrdf4y1EgPj7V1xC1+wv9kbHgbUCbv/
xv0IHxxYMy8sCHm8Wd02sfYjlnKV5hY1uQhOSupbGWS4PlX93WlAPE91cM1RSvThhKwwYJPO+GfX
p1tK0ubA18YxYYnfuLd5hexSyPL3/0967nQYmOf/ABsIT0K1YzYX3QhAcDS2BRFI7qSbts8ht3e9
WrcgAyIFQjInzvHxTnELVyXuufkgwoiuAnzdDFcQZpT1jfYPZBR9DUl7hteMqJ6o9gVBdbaO1z5m
4kWrE12VcmpF1tSTRj2LOCOn5KFdGkVw7q6XYJPEDjUDt6/YAUx0mBAYeMitzc/7N0AkPlHhK4Yp
2NTZe3ugsMDnzVbL9eOzthPtiBbmJ5jl/knfXH2HL7FU7NA5z3e2YI4I6znPxxp7LI/Xy5piBRaJ
n5E6VBjPqOqQd29mnWI+s13kIqrITjWd/z2S2Onr5hodyfVIk93VqRTICyw8UCUG1sWoKz1EemG4
EXa6I2CEZvNCjTrHRLEZtJtHs5mcqFNrQCpPORwQlVucz0Hhrx+Gm/qU3gbIhV72UjdONFZwZWrC
rlfglZRoS0hF6eOep2E30BpF0Yn6cjQ6+QiVXGogPWmxJwvuILtEq+X+6ijXxe8ATrpp45g5ajL3
sOZ7omMRVGOIJTv9aIWuoDvxHSTphXqeTjnT0luivRygRBfnc8+h96eLU+lnEl4uwZv5Fibk9n60
dx5HuozLaOelIKUiNOFrPnYH+XI2ftIF4sn9K/RLOA4WxI9cxKbuj4SJkWSWwfqx6xLbpsBcEzUt
GI0cEzCyTc7VktDyJ+FKUrYndBcLzjpGi82RbetM7T2wR6Qkrm4McQbLO1yaZwW0dkEM/XZhEirA
C2CiZNTSOAMNEl2a59tzN/sKR3ceRTEJS+aeVWNsOguETV9hG94eLAIm03ukwXxtwjXCsOc/DO0e
J31bia2ZctLGD0NFrOA2tvugpXQs21xV4C+8ADTq8FU4J0mrEkmiOywb4wNKlSWlX1IehYwLQ0fJ
5DLupn6pOlyoeL8sDgvt8DyfiFiOx9fISdO4BBR7Bg/+bsxZ2REp5Qd9SK2d/G2eBMgaKHoX95dQ
165MI0O+CsnJbZVE6GS3HBeklispzKQwqB7tsmAsLvfP7tGymnY+cjqn2NLdJaTMFjyfXiLwlsCO
2RDeCh00nhWBjGl+2eAtwvO64cxYS/uigJFEkSfrFYEccU9GB0VhXftlpCTP6i+ZyZnUJMuvI1Qu
+w949Lzn2Mbe/Xp0PIEEmjpFXkzXvQ86L267G5Kc6M6E+cv1rxQ6l5Hr0O7M5WAYA17XZbJSi5f4
GebAz86KxWYWaVnVqA2bRFOknMrrOVLPe/XVx6C74ONnlbQvjAxATiaaAHQt+IE0bQp9G2xUn26j
yZQRyvOPSwPZImrxQOOPvfkL4LADPE3hvBjs39jYBRURrRMM/PR7Yj6tK/ICw7Ctfv7CciKXrufg
7UvwOUzWsYnGSE2zoJdFjTXQoHpYO4GsRg/qsGbrR5UVYt4tBI12IzHLvc+JLO7JnNPxO6pFxTuG
xTSnFzc9/e8JKsI8mg3ccQa060g1Q08Ooxshee2TfEHFWac3bdjWaXcV083a2ty8do4X8TPLZ+eh
8G3GAgu5g5RCCvdzeaXgfip9koRarbDVHdJN39z4mzO/06FGVyNYV2GSii3TDhhQhaXIgr2Y4cK4
Vkxtq5wdcq26QIoI1jMb2bEdiUUid7RBWoK0h1bzzEhp/SIhvOsQju6Rb4Qm0n8sRkte0L3Sd/Tl
TxgeWEcfGI5qESYg8E6Qua6zoBzIqtIfriBize7mDExi0urHDeWUxlogjISwq7u4ZkSB3ftU0ej3
TQ/tLHWR7rSmzQPE0xsxy7ISxte3OE3uM8msdpaGgxXmHeGiAHAdqC4n7AVr7/SCQx9vj4XTJ8lC
yRBfe043ba+Q8nLEVym06K/VtwZWbJgP+yh+zQsPnIbxr9FlEtQL9VOKztGo2suoda2cimBMQ6/h
QYOkJLdEOpss1fCjLVA8AkuuPBUe4INUdvFm6OfCaKF/wZetI4r5HRuwAGgr8RV61+rziur7e+WS
dkLDZm02IuBWnReIX2FAbz49OLncllvcW9x105uxT5B2/QZJjVHyphctavrUY9T9Wa0lhCVty83n
+E3dP5FTkrPo3rmpW9c4tnuB09HSAExnkMrF8t3EJCA3myr1+1YWCa4BpVeJl5lXY8Ury5O2qSMH
+q5X58Dcjn51ner+5q0+aU9zKJ9zYgFqcFS2R/GE+9vf0818xJA3iqyglAMKycIN3gdCRCBM2Myj
Hnf59lME7lyb+a649RpIpZDUQYQ23WZfoLQBzIhkprgieXtFD+VX6w4TK04mUeRNk9y7fHJ1CJbM
6i/lmMHTRHjUje8UcxOgYqZQBKUkAlU+i1PZrLfwgC79OFYa8hpAkM+PyBFebSNmkW86Wu1ceKpk
5hiqg2O+HnVaECmf3BFQmKY1QPuRrfngttxMjnUU2kB9Q1oIGpguSSqhfstkdMJTYaYL5wVy1SRz
rRpycF3Dy7RbLGT2NmaDf+d9JdWRGpkFXD9DjGRCnGhO5QwCf/oJQPwRXu/YH5aR9FMR5HT0hl0Y
eaPJ9bkOQedLsqqzw3VxhOQTt57KshOMNN0QdR/si6BC8JaX+munCfGKQB+y4ORgU4yuPaBZElDE
bj5roKX0yZbIlBOVTnuUBZPX4AR4nXxMtrDYZcleAJjhY2Oz7+3zASsfVf2uUhDwM+ODacjgEbG4
ZHZsyOEHUER0nLuG1BoHf3r5xbPqSlCcwixIDToj3ubfJwkEa7qll4n/5csxHSFB+iz1tT4BPZFe
vBoiAA8yDiPnWaoDrou70Jzn0XxAq7mf5pJIFhZe4pyq5ZDKL8xt6IYx3jCOMmjnJjTwvtPIztiP
wJ2anqvuf3FVwXn+tSEW/ft2+NyWmIR+5B+3o1SD2gsJF9uQhjZk01HoskySzgr6hoijFyyaGa6F
8z1K3zW/fdkVXMkxDhQG2jz7FBHBD2jJjR2DDxyMrIfn/7RV+Pw19uYeUTtS4QgiA9LrwCNTgL0j
4p1s1DRvqZZARYY/WWOt2T3g9F3A5a6mcYSgysm+eT04LwgrUnvERDCtRwKhaUCvHXs8gTFpGuDa
eVlDgNdvBvM2Z/Cp2wYNMpZ/VN/d0g9bXRzw+6ZpeV0jvLn+8GwoXodjVx4osF2GAKbmItJegWBn
leEwZUNX1/K5jwvpuNoNZUpFmXbXJGB+UG9+9BzHmMbop8nq0JUsPVZ0hNRuHDrf7JRTuqbU7tFI
44DjOd6CXJC83IwOP6N4QCTWfoFTHr9l+wkUttSDos7aQraRZNYy/VoUVZpD9nnhRthtVs/MbpZV
1m12/StRZOQzdcq46pb2fLv89QNWgsxrOc1xoTdv86ULNpFtRjT71399kOUopm/Et1kyg2qCTc+J
JWves9yCrgTaoLwffkaJ6g3JNinL/KJf9Iof6UGa7mOSXOzFMR09v3iUExg/dIKfwlEPEE/KIQ73
DR7l1U0t0tOYeGBUYh7d53rB5Oj5AUxqrYHHiov9sda9kqeEBNdES9ADoE76XRbO9k5yMPt10dVS
KVuAKx2Z254DJ3F5M+rb/2VVZC6ooUyMUc6b87ZEggBSCvxR5j9xWkxLDhkg66waGqsS1lZhmWGT
kyBkFy9kib1qMlbnYPHHaD3aQBXsanquc9Qae6EP1rFmtQ1iaPxtNGjh494jqsoL/wsu4K4UFWL3
l+En1eJ8Tkh/eLZ2ioS5jqOtGT75wgaHiNF/ZezBegw+c+3k45SyQMjN2ePUaMM4adstXtqA4Jkb
RMIPdaQ2iiiywW2Ifmf0hJXVi5NUsV+DdwJWLgL1AQjjgh53egqMm5N/Z8PmtwFDxvOVGtkbeLKP
sWD2n03Ywh1sh0ZovRTgILcinSM53V+0ZxhGr3sFbSUZdRG1qQYMmWmpdtfIhoHm6H6/sJ4P1Dgl
ge+4BhXIK7aAK/SNIlcGd7GBllSWQq9+PkbOCdJWqfdaYc5+ufC7BNdhClQFUX+qwETWdQq4z6Cj
NQ1X6dk+gGeE3rDjqIUSAv1lYtirPolUo7ZZPeB6iJXcuhFowHG6+lovSsoxiWjKdWfzElK/fIrW
/Yz5fgf42SoMGvqM4feTTYDfVxRkVyafFkghLsJ5o84lezQjZffzbjrUvatmS0Kd6P0hnuDznUNc
MfI1xPZTOwKg7KsIMpC5earkAWQgBOBsVPIVYWcaKsQbqKYJFH3x8qtGySM4i4nNs2iRByl2bttq
tlH7kgP+39vd3uDnFlJQoYUlDI3veIL1Arcn61ipK/HwC+WABYeeHYLg8UbKurupX1/2cjSX8C3G
TOvr5pZL4A5QLAtDvogoIjMJ+vhfivNqzivC4+bWmEB9PaQeV077i8XDe8sKyxfEXWUYXBSMNPIo
VF44ucQpQG4WJ5UuA176EyLb/pms4EC7KxmY4GiAFmO548KjwXRj+hI4InLXPZXO+CV2S3feulJz
zH0SCAf1D+86c/i+UwsuCJ5WfFrlKEvG2C/6yxFJY6u8Rci8jpLEihdHZn+f70uhR/jpyuBGaBbZ
PAEo061Rs7Ga/3RKBTMI4R/Vd6nwy+i+8aoi3o+LEM9PuBc6evJgB83YW7pyZlPD50QoD4WJOKZR
MEMrdtKAS53kCtE/m7ne+20WzwmgTj4nn2aAzb6o/ssXYHI/lYaG13jvXbsz3oDEFlAoZd7OpVTl
OoMTVaYcb/wkr1mYpxxgHxLavzKSeGgHTckJkDK0cf+CMvm1my6UmDlXF5iW4Co8dwXc8kgI3BMs
YQDe+tBl8rEGRUQrc9btzDLD/qufv/w3mD3NpBZ1Y2NZPnIMBmr6gVUE91lRvo/mN2s1ywkWHbd2
MiN1n0mLwYAoWm6inOskcT+CCQ2fyHzhuvNCMObgEDQf2Clpt5+O27rPNI/aifcgwhZduaCXeHqZ
2mLRN7k6VRVhuLUZUWeeYVKQCUuBAtLBpK+mpUb/YJi2lItxtkC/5q15veASi54epREifNtJvE6/
AGN3RakPnmzVieHdPCD8yjf7PjmtGVkqBVwlmkPuKBg9KkRkO5U6Ov44cTcTlPmgKeVTwOgvmsgc
3+DQg3w0uMnFJe+dT1vc5cFi1VjgmCdBbEjEBE4aWy9VhVFVFn96iwldfkxABHCzEBBYGGgATPZA
b6NE8Wedry377z56pFNB8sSk1zJ95OFWRAnc+V+NMc5YyonnKoQi48Sq0USXrpX7jIVm/AUaKO1b
VZ9iVhVcp2LHu2l/BWalD4zmgoEoufBr+0AmHZ17FURZpH0Jj3hOBojofgVvvmG+j5wix19GRgla
kyKge9iz2TxglIxwtdx8NOLBTrbn5NX/A20Cgh/fX1iAWJuTP5CUIQaLcyV1mBE6CsCgwSnAhcCt
uDgj6oZ0L1dAOVZgOBZs7jcFp0LHXbE1OOTACM3VgeWJuB48VdozLsIEzENXBYMZQTs1a9TrLuDk
a2nSV82k+AjW71HUA0n4pGYM3wwzDGIVHGfbIOR8kCQQwle6ruiF8AOoOEKBI8G5QN8Jovuze8RS
wY5nbXfxMZpOZqHMqQ237eubBJP3swcqKrQcUCR4Ly97qrVV/u+e30Ea9h5AgA8vo5PS7rhAEDrJ
gtqqnEeEuIE7RoTbSTupIu12jIFq+R9GKxfI22Dvj5cfDvVtApSf0hdB8LG2nkU4W/Y68CByIG1Q
BQfPBfYCJHdcVaA6IuVwBYaasWzfAViLX6QCFtH9kGiCcPL0EZvtSx63fmzMeHL3xiNx/gOgQ5JK
+Fxf1ccd97cmg1lL2MoCnpz9TUcOf4zlWNzSFsLLpi3BjOv1qN7/qLLOZDz/nJAM91H1SzhOeNxD
IEkOCmXmAw50LdE/2AbPRQsyH9tbSyof7Xv87JYqrenuA/mzgdA4IdIGFaesb3xwTE4teOHLaeCx
fvW8SaoHz99k2DisDSc/OEfgg9c/XdKMrWnMXllCHTzWqjaYsz6IkMTq7/QoDPcdPTH7B4qZaTjf
Y8mYA6kbfcKAwRV8ZqYRHxf2PRlulLuD6jWVG7PaA98L9fNDeZIqkPrlVy4XXO6snOpoIzuI2avy
O8uWURvgisiVeYevWNyDrLNgRsYb6QANNgEiJtcBk/2QRYbPVWJcI89ynUukkydcTl5i2ISdYVS+
1UscZFz/E9X8Pudqh1B/nhM/Y43BboRQJaapEuVrNzxMgvlP0WYLBb5707JgaFzpJfQZQ1lOOHGF
xUjRQtKzvsADUDcd3Dudqst7Lomo7sjFLFA08i7ta1lnE46V5+CtWgYUjUKqs3f75c9oJPnYCl8f
u7sbaG51+xP6Kwv8VtAnfTTXaY0wST6kxZElVaSIxci6k8sl5LWnVrHxF0a8CIFLFhgGh4EpCICg
nlXi+S+5Kt/ju9HQSMDdsfhQE0+TQKelOSEqWdZX/XH0q7TtMr6w92ca/nm9rFPq5pFeR+wp3nGE
LrG+FNCCIMjehg4d3WwhthuwygjDKhcHX7CWXloPZoDpRbQCfb0XKdC4FNRkkCAhtUARizgMFIr8
AkNZsMt+d9Ni0Oq56/TSrMmvoCmgKi3VW/ZmFiKGjRj9KzY0Hr9qXTKCTIfWP5yHf72rb0zvQsOS
Q1L+5QhHeOzOOOCzXs684IO0RmA3H+j7KBK3ISsG9eFAMmkzd1XIH8IPe5h4t+R2T3gmiPRagSvg
0kLXBVu+Vp33rDzh8IJwTEHJmrNf2WiVZEZpGVGPh3L19luAfX/gDiAJQkIyrhl0jycJ206m9/SK
oJw+AbRSBrgpB/1WlzkW3j7yMl2ej1hVI1UJPNW0H7MLCdB0sGe9+MQ5z1Txs93cyHLxBhafYEaS
wm6Yrh6blKCn0iZq4/E1Y82sjtAq3iALY/fijZLZGZgXfQZ9JARfSI7jdVW2ddXoKYYt89BQYXXL
dW8YD4nM/Mao0WpwQr6EhP+2m0/zJlrjgIm+vNTY5Xp7eex3HIF+HiJscbxopye46C/At7DnesRe
Uj7v4YPc5yI0PWC5qPAY1ac791XJV+QKL+TiALLzx3qBIExX9VOLhO63vw/k0a3OhdSxUMSqYNc1
9es/CFFHIaRl3GnMaYwUPz+GXh0+jrfpLvyvhD50TRqQ2n5TRPIsVmSNXlqZJemxp+gYDbaljPRT
O4o7At8nj//ADEsLdSYeZTpq5qxXplT/DVvIxxPl+/Vt/89KFQlFyiVpFc1O2nfd94wnZWAUepd+
rFNEBFcnuLV8u9qc2iotpygSOMbTGf6LACI0X39k6VAuDw7x+JQbCT+FMjZWAQo8sHDJtoqJ/c7W
5tbLpQbAbtdrN0T91s95neJCzRzx/+BWg3S9AA6C4b6XavxSkTAisZuHJuNJtAQ4nYAf/i1Q4ner
mEyb3nb8pmsL2Ur4g90L8Twc9JSZlLlb0YV953SpTnTO5DWt1o1jMBcpDUNMBPzyNyfbAQJrnHol
yg8BYHiJd2sfLFeDNzSXYSOV/l/vFf5m8aRX3mhVTc6riPmbMQzY+kVIwC/fuSuKPMhntV+LPrqj
y3oQzE93YP97O0UI/CEv2pnzhsXLy4cpvfrdwhiuYTX8o5dk/Xkrq9BFGsj+s4RO6zZiZ69nuchy
e4wE96lDZydBX8ZxTv/keXOFVjfhZCXFytXYj/uutTY9/JbM6kGl8kzsFMzHRX8l9Nzb4BNw6aD7
pLk6k7yqs9I9HENfwu0e3cmdJisHOQOBxbB8qUp7kaff3H9/Fex0Ah2SK75yH+h3Ei1/QoR57veL
YZ2029VVaqa2Tlt6XgZCvKY1HSqwpBqUfbBZhm0tkFwnNqHxGNqXyDE62L6JwUUDxACy/HQusWot
pMUmz7advxpMaMSxX8OGQa5Q6pCKfTGQZCcufAbFk+uvkds+LuNCdKhFy/tnjMGnoovv60n0SBgG
QxDfx62aW+7qU72FHqKU2mHeeZQ2aK67r6qKBYCAhSLKYW4iH167IqzEx8Ketf9bG+C5AmBzCK67
keUsT6WJi4MxBMx7sBCZVvmCq9qd1lSTXH96C+B6u9exW0SiXY5krhpatFyAhuFSF+nNiGZCGoKm
t2O4Ls7cvAUi8W5JJ8VPUf99yaEvhtob2r9bvvwk3LHBOy5VlCLI+h8ZKBO3q6/V3Tkdcxykj8f+
QFl22UL/qomxBLd1HwCAGL89raLiBvoAlzMCE39+F/3LDvscUVfWQ/6b0dc0oOvS75TXI2WEbJGT
Ju1s4o9/w0DZ8atXZ2XQoDLV3OKp5bQyiAOEXsJlZ8b1Cw1jXMrBnaQd3dBMHGBk/SdcK6OpROUq
/dNBRVde+YnS2F5P33jEIMv9jjfx2l6HN41KfcfbWETkinYbR9yrR0fMnGVC3DttotuR5f4ITfzY
ToYXJ+3J3lqHT1AMqYCURaZppsGlhgq3Uzs9+X8+3Pw+MUe4/XU02UaEMbcANwPwfX9oBPlslBNI
amXnmYWR6m4T+yVGZr1wAKx3KTTPeQvPqH+TDARSTaPdZNUDvgskTA+ysjtmuClQXGPOjL8863dp
1FaJ3b84k7hHRxYZyQnnnVNIS+WXbfohKtgDtWYSh/kYX7zo5SK2jt5xeXP0NbNzlYZmEY6D+Hht
A9XSNPK9sZibqv8QFbeCSX23xTQufFBSoQiUA3gvV83LxoSJLUowcYvwX/pll7zqdqvg+L/8rO7t
NZ29YwJtB8PAJRxW9VaY2qiGjw1ct/kmlZE1WjrnN3yB/63Mptq1cooH5WNin79X69bL4N/xzIZH
GnG+B0KUclaCzQEW7YqxKO0fB+5LIdr1Kd72cRIv45OPduYNrFOh3BqPUtMZWao6SoodiwSOHLm8
n+/Y9KPzCNoUMR4hvozh4SG1UJKyDx1w+Bi/JVk+T6NvNE8DoM9LdaGVrqccEt0Y9B64QDtQJBpv
ArW4WVGMIV1Resey49H4Ut48Dcutiy1TnONTonOSIacMgxjSM8MevcQtwxOYmMYwKwy9gwhnovuE
Naq8sQbZ37PPk4vO5rY/kllT+fjV4JyAy/pH/u8b2RBTG+7tTjs2Us281ngV5yqj46cVsI4iig2I
Faj5NHaLv08CnA2YpMPv8G6oOVVknNxzkWYQQFztpYIPuhpNxJHA1hJKg9ml55c+5S7OVH5Kp38h
0mVDgd3vnOExyktf1jadMPqAcmozb5WtRd9cIzyuR4tyPvS6FdrASFBg9DBzatHdXIcJGMkZj58B
3kWLf+SDMS2OUYMVIrP0Pn8kyIPD1L1Kl7iOBzmIvpFBfcp6qjIlCdw6xNBTzymyks3rVBgfCT3g
PJZvXecaxpH//MasZR+PvHRuvAAi2pzcpEzA9zDyD9wzqy/HWBn1mvCASFBX/lAMwQO9pvMhkrHO
mgJrlXqQWGEIUbd9Bx1RIESSaWugp6HCPnDYSbMc5oFk55kaQ4aOqI3NGBTLqgHznk84oDwoE66z
iQqcA0DzVAYfUoioRwmy2m08qkzjdNNvzg0nkFSLo1lZ2MYXkIaaRDDvNMs/YOdLNQMiL3bsvkXg
sZO1VkGT51CDwY0T0yIT5gCRJFJKTbusEZx4bEfFbhs0dq/mLKDPCuM3qAVKnFkIsOKbgIUyfH98
4BXPoSsf35Sd0p7PiOs0D4QUMhdySqMEecfl0CikR5Hu2vc69g45/FyNnRk6Ku2pXbZ9ZpICBPbm
F1OME9fea1HjFomhGmOroRFB96jNVravJ9uvq42Z5MvVgjb+9KM6/HUAx6ruIf0YYRAvh0mHeOpO
MlfHUZd+qoNOcpe74jSNJjg00zoH9xafCU6SJ1IUynyKm3mT8WZy6QzbXf0wdZfikK8eAM63Joad
Cm9dILWMdoCMehAHa+EsolEphYc5PPR7dF5RwIOWYwXIfHPhJretjbrZEJshbV/Ve1DRBQOqMmMV
FuC22VZLQ3R2FjAvrT6ck5EQTdEIMSXS1tsgOqDd1tgBwMmILDawdmNmsNpbFyQWCy/YBtvHymkk
iwNUTmvS3uwwQvrS3spEFASXocLOiWvs5AFklu9HapUhfLMHeh8RvsJwexWQsQMeVNrBc6gcmuLP
MQRinbPuOPwU3mqfBYJnC/9LoVBYsCDU68LMKHzSdazpZWKUuOWDG7ighp9z5o/0hn5Iu4ah6zKu
ycpSFt5VrlGUtiaHA24UaLAT1wdsIIq7tnzEP0RSymzxCHQsscW0C2VW6D1i0fc6/iO1mf9UNJw1
ZLVS8hO9m90eCNfdYYJwgiqDVBq0B7ysoGW9pqbRuDt4cX9hYcR/PF69p/WZqmvJ9OzBnX0EXt5N
+DEpEIQq6YycU2Y3Xfp0xDdTH6FY5NSuv8VKr6fmPgAnQ9Mp4ky9SIner6ZerlM9X8olZX6M2dol
65l/isK65nav3rL5g1FHgeP4GfRDPmGwtm5yA+G/0sGoLN+UqR9G0MCo5AzNMCCCBxCCZ7S9X6g8
Wv4iKdbYpSGrpEZqWncmHU4tuqy++EFw1p1KphVuZAr0LV/x6CG6gUV71yIuiLIA78MYryJ2Yevd
9x8TWP8WVzBrUX6bfFrMlBTDytFFzp+jIaYXJ1thRV3oogdM8ImFINIiASV1iVuBdJTPdZwZB//R
jv9bUbQ/um7Od6wA+RuJ3zwZoDlNQaAjYjrIPDzjdTiShaWAz9HxMGELYE+jb8xQ/QQ7dMv0zbFw
ltL/Y5Mv+VwkFbNLbzfb4xiGUIUhukrVJg6jOHddz3W6d6XmfUHOT2nB25+O0NwQ4S+C4d6weVYL
eBk2SjCCrWiaRWa6nU1Hirt/4MGlEUq/ShHW4R6ce01l7W5SpDEK9zxDDCAk3kHnL10fl0hbo1oi
KgyUErj3QtrLxpWcLx6EmjzBMTrRqlPQ0SwT5SKhcLOB35Gofpg4qUQhkZ3AGo/6qFnk8+EAk5kE
gPIgtUXBvlcjWfv6qKkzNDUuhAnb9Q9AMSwSfPNyAfdfXYnTE9JREh5LX/Bih7GL1H8/q6R8K4m5
gCpKl6448pZDls3JVpul1MpomEQlt89aFmHLAjCvXdkW9PJa5dCRDvbveCRmlPaI3vO+ShFWIZ2f
CAn/kyXhPdT7hDhMgrgDhKfqs6NX8riLhQOGb1sk/xs92K69g+RG5NYzM/wukcwGGIBbIfqbFMen
XA7d8uEeyjpxFLXtYjy0I80nDsFmhnD37r0/6s3KhCcQlavmMzu5f8UGbbApS0RsnsXbdkAhp8JA
ghklAc28MpTzzVOEwo1NoSNINC1MHKBJELHUq7i8myQNGAGGmf2QndECRLnET+vCBqToa0am6T+G
MGK2IKifY84QcJ1LQ7yGFzDnHWiMBt98r6YpYkqtoCxnkw9u/ZotAUMwWn1ZqQvTFFOIxfO7qYDz
CIUjzzZLRLPddExY/oZjlQhxGt+nOvlJzJ9lV1TYMTfIiQOhS+GBlZpY0k7pLosf/12gIvjbB0Nm
tMYvquqi2g0vIcpzNug1cj0ZZ3yd/iwdfzaHj4+9mqnE0RHZJOrhMNea+YVOPddzvLtvHLtykCUX
I883N5pLIJjpBGBrip21ebfbm+nVZyuFnxEdGFYJkP5M1LHmqxxSwmOm2Mbk51kb4icVjqZULI4k
jegSu3FGIXZx7fLtymPEm9CqNDZ4aDbey76cIMwtwg5VRv6FBvAvvHBtN2GtOcoHgMoSXHgq8hLq
C0jRwGUjymGKdKTKQ3AcHy7xg0j/vSO/Br0fU0tTTvJPKy0f4s8dWajWec12PmFLHx84JF6cfwps
TniQ7IWzFUJvRLQuPUHzdz5wbd0IV7rRT2M511uhdj0CJCsbZFrC+EBbszwIk1ITAcNpoQlE1qq+
VdU76YGb8sM70d3TI2VWP/8x/g2K91W8EGJ8s/vTLjJufZWhUJnJrEJFgorymIts+h9L3WQ7jrxN
7ZlitPtX4gWJ+tKRy88L3YYvX76uKql3MQZFuFGiuzxOieNHWJwmny5utFM1jAUiXOINL2zWQSIE
KTZlVorsLFDBwyFyc7p/oPRB4UWjQuSdMtPNfA7eRMRgJvd9Ts1wHFuuIKXWL/dT7YtoQo+TuKB3
r0cZ8l2Ukvx9dr5CT/NrPtgyrKcx7x6v13+FDxzGsyG6LDrY/pJfAc6pAorjihT4oHqhIsia3QuS
CIEMn1DSA9WC//yc82TdOwlVHPl7FRdeNey5Xofyvaqac0uMIpJTI1fDm/+0BJEpsCCdmBkniH3U
Kp2qZSA3aYkNYw3pIxiILlgcSx5tFB+/BBYxTB3jIgZpw3GeBrmJVVJ+pJT6olvcB5L9lwpqMnwi
PsjlGlrA5ur/fSmeXIjy9+hnGYl7uI+p9QR+okga4r9zX1k/w57nNPMaUiM4vNqiIxNWCI6G59Ox
j4kj8rAzfKb8hwpyNT5tn7iR7oXsMBigpqsZUYQ3q42DLyNoFnrJdOzyfosprFuAeRCnAiosoAvS
rxJyaGVP2oAlQ3E9GU8DdBWwNzKyKZS6K1S0nHH9XkRq9hkmoRvmZfx93U9iixt0hK2v90xLoWyj
MoXnBRVKFCWECM/iOrByVgyV6TFsTian1MIWBndM6FTKBajGsZ7OazYZ7M9//Vk5wW1QnoHrKn0J
iI2PgYhLIJ72AoknMxNIO+amamanv1DS7UOQ2lS3AOaBajYMemMEPBoJcyFRdyn/oCp01As6mjqx
zW8IAyP4xNo4SKqdpI1r6y6AoxHFY12ToHA+Bonn72I4ls85soJLXn7EZin0vf78512K4TvtSBx4
nJHGw8Y+OuqPTbzvy2v5x4PTslq12VtwieyhrN3E1cuEmuKMnEdMYcPDArAR7I+GFknttI7Poc9c
Eqr6HDrA9rv+ySM6Ninihxz15/TC2yzMWd+sEFir69RfR6hGtGcm4PEDmJAQ0kARfRKNMgchHyvX
5+Uk1etL3MYNKjIdugrEu4H4rcpxmAZSdzMl8GrOg3iJdwUcKZ/vzr1NOUHwkZA21vHpyBHnXGKc
3dDJYSzYjGagnvCc5xVBU5pENZNgEoqB1ix6oBkBI8/daz7dcgq3V08DwxoCcd71BxBtuEQwmZnj
0Qz8QJ9FuAtjagW0xSluMijB7Ynm0SNM5EaLN+20ILKku1229aI2R30da3YHrSLxTUwO001suXRu
9H2xUlnpcuHh+firaB3WTYAs0dx9yIOwqBblowY3XZ7jIroXGN+AOrIMDC0V9zDXbxnx7mmUQEPY
qYbepFQqztAc2KatAieXrfHcZZqrclK40O8sNvHodx2/+1jWLQ8bC5Xg5mxf+tvEoGU+NANO9+fl
NMSc32DhsIy0Mpmr80SW1SldHhPycUavtDm5sumqVN2ZOd/VZFpGtFZ/jCt5iT2QKfezt7bW2DsI
U6R7WC2Ew7RRA8T2y46IglGFvfktGMvuZMpt0kbeBBK9UU9MbLjXLpLg4YVY5r8CJuS/xKro6JbC
pa/snNFvH/ejnkvGwgVdUlX6cO6adG1pn77fieeJ8bzvJnYLzBbaGv/w9IbGyTydP+mRVFf8Jiwm
n9hn5L+ITMl8KEzBSjslyvCmn8+7/qfpW9a0coZovFpErhEfoesWpe7nBrRE8DdUzJJFWm0fAzDb
H6V1rgsvrB+SVFAPf95A2WlnlnyPkNQue14WdD6uGAxlPRiM0+MTiqqtoju8tVaSSaW/YFTRsgzy
EcmzraQR6XMgOTXoodqdqT1qHSGWQPLr2JE/PiMXwUIZRp7KfpGcZxdhroXxF/NHAlv5lZny4jr1
0e30S6Tu2TwhyVy4ggN/uGEcfjjo4/ifbmS/11Q7T905zPwU4gFR1emWAKq8L06YZaIcIsNa0Dk1
ZULSXjbWb3dYv4Qre+ECwdZFoYCmpLSHo3BsAIm2CFmv2QfykxBo/EDDfibPZ7gBiihWKG8xDCNs
SY9jl1Gnf1LZ2gm8K1+gHQ/RwftF9fItLs2Rkwx0m1njYYpWlUuEwboPUl6OphpT+8hCVeIu+rsI
dMc1U2VaNV55Jmza97RiFqertEMxNDS1DHGiCqaG+HtzsLLjfcUHWtOiz2SVrLQRPSkKcza0EkJo
xQnt21fVUXj9LtYCrnoc/xogBIPcj1bQw4J3gwKswmgnyq7J91n6UasdpLUTA4NvEg4GDyPncNP+
SjpN9jQAK2aO6dw/hx6Ef5PgBC8aL3jJEjfFbxQaGAYRqYQVmDbDw839Pj+/+aWZHI7OKGKuD1tl
hnJUcc+TcvXiUcUNkvQBXMXTeieX7uewgPReti9R538Wzf0LvpNqALG7pgLI59ZmrpaVNWdkjzvC
AWl12RhNup+aKDA3LHJnXHK5UGB6PxZ+j2xFxb64BcFHbQjZGhKk2osg7H2tJWNjS+x8tfiDdzB/
3Nrhrv8lp/5bGNeQtLC+ECyhPNKTrwXUPlxKPimvRuydhhEd3jAPjdZk443/lmHBOt1PyUo+e6Bp
AihNbOD1YpHxE8nvFsqTlL1Yx/AwshVHF9RGsQi98NcXv2zz4O048kN0un4hmewVSa2hJQXz+s0f
xU7PCZnIJjsHzfREcJZ5+Agb+D0d4EmeaZXQoQr2uaVjj5NmeJN2vaTuzBvlw6pXduFS6FnEyagP
uJRICF/ESMnrEOtd+z+Khw6qrSWHZwwFoKb/ngkMAQP/CvesYhjbIXVCVs7gyAY8MK4jr0vtt1fa
SZtb0VEcAjvWPzn37iQ88vp8/DG+m2R4i4sj3tWM2c2j6mUeu1XqDUhqvL8g+m/jPolU/ObTO0ld
WtiyGS7Fk1bEjja6RRUEThOc9UIdtJHYIKk3/CEX0/YNbosgYF/2i2JEMV5fUF0ajBeW7UUA9cCv
9nx1KSRydvisM/ne3WeCbSCU0/mXBzyWq4XbBX55X4qVk7UP8dkVnZ2XgpvgiZ5xZK6LTf6sge7w
PudJF2Je9v7ILGcWJYGnuSFMoXQaSNy6KDrjAzP1QCt4GQNeKmUiDLJwnVOrwZMVLx2ywUDl5yAU
9J3du0UO0YcZbpmkr6EEKlojGOwT5seaQEnEGyTpvtAEXn5lpFfZhAOOgT4EySPatGIZ/g7ikQEi
RAW5OHn92a18LtrEPeJhGm7yp9JNJVRuoGUF75bnozpLmDPl0A/+CPPisctz5JQR6dZShDyKgFfa
Tf5Bywa2jztQb+JYCHwmwLaFbwYcOnbv0KbGNsCx8LJEVOGItdNSNR57SpiP4d4IzcrnQTBvG8pm
Nzf95r2kxegrbjxD7zwH514gEgUyxT/BW2sEqwuwf0sOUzFrUqsY0KauFmVi2DnVYgOuWQ1xnZAe
H6Cyu9NALHu5fVlQMdKH9F3fXyre5sEY2Ry+TE8ARkrZzZwyKHjV1M2uB7nfcAyAJsnBHLWQe+z0
vUlwok1rVjw4YeoiKOTuN3alOcPQUtyQ/qf0SYEs4+Ec4Zmuv1NgqMI9IM5Q5WRq6PqcsEz0HiL1
ZCAgZV8e1zKjinir0qH/xigwJfSelfXNKc5u45mjCyQz36sZ7dGbsCh9TbPh/Enqgsi12O5VFwkA
8YrpaRl+SVnp7noHZnJDlcwjidsYs4jAFM7M50aMXj9kFHjKdqOswlk4kswaR30ksByUTrWlt7wq
ipJuuozymqqFnllWk0x0avcq0LfpIg0QIIa6IUQJmu+9AEwqU2ziuOnKMwv/MLimKR1BCP4Xce2a
INs4YG22rl0ofwLPdGIaxzHOktYdmfeWu/KWofVvIYKU7NYhJ39Pg4MpiIXgLX0VaqtxnnQwcTqb
gK//zfqUHp/+LP2BAoDIK9j8L2IYWPB9+SLlLLGguTQU1PGGUBQCEVDCi54mizr06jqmC2/oqGMd
8jlJ4XCoDLy9+muvd2X5yqrHeCeZURZ7kMyxfeMP28mxqQQJH0n8zO0QVxJ/eBd7z4OIwInlitrQ
9eydPcffwh0/Wl9KYQxYA8tVnQnw2kyPWBAKtRWv5OmEEnI/LObCAIFiFoKO1CrX252YwRf0uPQo
K3h6z7DVpZ325lSPOnIVpNb3BncKl7x1xKLQeqMKWY77BQH0NHH41GLWt/y3hU/G2RniFQ6AsSCp
EE2Khz05ItIJewu3T9sMug6gTz5D6RZdhoXe0CLUdDj/CUVG26DuCIYhZpKHtT+oLlqOp9rJLclP
QdGPyrRP8ao9uDVsMb20+RuR06dPatabO9/i6UZjJNdXB7eWJG/VDi1l8xp8/NUD1ty66XgQ4/qM
NOSPMi9HxyaDmKZSsMLkPSuJVHr2rBvO/YRGfvFipQo4t8ULfBZ15BsepdQJoqbrNfQil+DuxOAL
xhkgHlzmUbSMXaAddEMmdyffLq3Na14LbdM1Taw6jniJ9vfTHVSXqY7keXYa86rAIST11z4fDXbu
uMw4FqhxxTGonROa/j/p+NNjspAE7oa2um/cA6LUakmL2fLk/tA1HVc+mx4GT25+g0MftAEL0JUf
may4pA/6DMmMzyDUQIbtgZSecieI+G7C7q86XTGmu+pFkQiC7ZQ7R5KUexQfF2awChhUUekIp95h
011cpj+fAGd+NjPhSND6W3Vfv08jo7wBATqEf3M4kSou97/Nipg9coxh0r4Q4ZN9fZfb5hSeATe2
Cjic8Ef8y9YXOZcEKwfUcYWAwEYwHUKvWet3NMPiUTNHsZRzau0IAVxgn6gbo/sHYg9l1h2hzTq1
nkCgfGl/CR42WLn2yFN/Q4NQzTb+BjXapCKqGCAjuV9H7scXPDGGzww682oycTGEOwQ4IGyAqzvE
17Tq82GVnd161NsFQNhSCJiTu8tmHPNVRZYuasK4ZbRlydt0WJM8RqcPX3or3vvL5pZMONY0lUpD
UMf3z6WlKpflYrDvZ3KS5IwSrn4Z8EhkseL/LKuvlIoXPA3a9AkxpUpvNwgYiEOavIueTHDMIU8R
TSRQTiSP425UDNGHtniaF55+3cXYS24BUbJvTPk4IGJsxxC6N1fNdSD6CwmYPfH1znhiK/TM0kWM
Qpnuy6a/iCj8DxknLwL1Mqnnt3PT7/B2LwYKs/b4hX7I/Di9EP5hMFWGY6WyC+wh7bTlADscxJI/
QR2MdN5sqBFy7irOr4F4fEDwsO/VVtCzuoq+1TuKFyH73F7Jgv+kXXfdUlTCqNw3mXeQtS+yzFSQ
z0LbkI4PEOMSbo3Zw3KTs20oJa20hPnx4WJyvnQ5azt+mIhSpeKHE2rDw/BPsyRXN3I2DziQr6LS
W1qeMmmAB8w6zoMovJUzpzyfW2ofuSBduq1XXAH7p+Zzdc3RcxcjKj7pcZI/thMQ/VuVnuRMxO9J
XPiMW/MuJVAmBh9iY0XtNs6J2JP/YtRBIZrhhTeJmtQ85Lu1jpQEhKaYksG5Jp+j8twkbokq5NId
mTHYNpGzW5BNnDZutl+HosgI7/DWL+lUVriiXmvEhoNM7eD3E7bETXm0zx3wj0+LLPMwd61Dfxuh
eRvrTsogx1lsKVHmHfaDqzMsGHmb2ZfTf+u/sJHwNanzb44zW1NlmjS0DXifG5SBqdQQU0+bbp0E
0jIIVpS0bGNjiv4SR+kdNcmXDootyYTRR+9zvUidYhdtc+ZHyNhnmO6R7HY1zQnwUzHNuhFzQWUs
I7zIpra6MWtO1yD8zlFLU2c8Af/KeqSMY61776QwSxn6Xr7R8p/2lG2bgNTVi+LllKRnL6izPyEO
lJ0JU4EtFYoSorhXTl+mUSVvk700DawqpZ9V5Z/lzR7AaoJaJZ9LsrmoTxA2T2bB3oj60bhLEMe7
/b2xlgj2JtwX/JV+6KvtJTJJIHkvCWq13Wca+qauWRwtFmZ7LUxQSX0lokh4qKmt5l+de97o/VOH
50zoSI4QhAU94E4I3OE/f4n1QgAJyl9A3Xf1Pm7zFy2axNgSgrscrdAmtXmHi6RCctynhL3+Tw+2
EGvG3w+o4ULOBBzKez5oMN6zrQjSd07BjyCDCTi05tbFO6Gxu86ZwfmMl1wg2AktZHApneIZpLVG
ih6gxq8uxgtM80Nuxk8akBAE5VV7xDOIVTeos6PJpsjycsruZi5cudyh3S/X7eqOusSL3dQvvT5J
QW/xOnwZJ5ILZIqSv2yC36ps20rqGKwwXWPQq1nx0lheWPkgyc9d27uwZt58NsATnPSAwdSjvF5/
VS6Qzt6tuvw8FtIKMIn/iHXKGxnWkGXFJxiBvpBm1V+wuIpZ80d66r+frqkhWp+t845EVKWRNTM+
nq0/MaDfrSVZv0TJqi79mqHdJvRELk84VS56dPuYAkiZel2UqYmtMODZmcVlp6q9BjmDtmC5xXDZ
xwPW41mukutM854NtNtar5V0gbrBXq0Y7BaiVG4wYmUaawozQHEEjsYxmV5/T1V1t72j9s4o8WZC
LmLQB1qnboIk+KtmnKzwSTb6L2Sb4FjTYZqdWI+XTeKwDBQVa8C/RpkG1Yg9nZK0NBsykSNGA4FD
uo+LpXTX71x054RN0yKAYStHwsynJSuIr8oJSY14Noq6bQRdj/iLQYM4e9GvAReRxOEHI9qVWOCV
ka3kPc3an0jNHPODEsRYerQcR6bs0XWzis7qkOvwqSQmS4v4YmHEnD8XicyPleuBNIO2ePwsNRhP
LwdFkgjpo1UwuU/bV/TwoqX+zSuxdngBEAzBM4/2EIqkQyuP6rETZwsu8cVL7552cxAxBkT2T3Zk
l12lmjw3nLDBErlV3ydBeA2VrNYIJFfsp1kGpYPxjzoGIa10JwpSdY/uW6AbfBA6KoNH73f0/YA3
vd/svx9sCWUfB9dOXBo2mhAS7fBQ0JHeXyIV+FBT6P7/6g1JfzKp9xOLY+Y/5mUiZt+B7Q4AKHHR
eG2/9+8v62SuR72t+VApbQbW2c+spwwtjMmukFgU+UR6/KTL8dml3Y1MGxndhEi0rdZBsohW9tz6
GSHTGU8N6s7gllZXYuWYW3WnTAO/paDkrys8xjefxgvDOXqls095waiJQeIJ0XxirllY5MX3i3sN
yjq5NSQqqaXE7QQNaHjVSA0J1oePaPKeAVzcOXWi9cYujMEz4gQPx0yvjJ/9e2UrVfv9vOcz17AU
afUxHotHYg4HF5YFw1aSShCivO4IJItg3JyFCM2gDDh9uhfANhgvKi1UAQKrL6Q0F8HUNxRygLj+
4Ug7d5Jgd+wO+2wOfMacckbBQhSqJL2SN6j3W60xFLaMwQ4H/wj5DAqbTRdL6+mKCT9lONX/XsRJ
VU5jS3ephhYKA9ibc67T6cEe2fX8RHo5n7x3uxtKrtbBLNdXTNO0QOmoEzKafosPfoAJu4G0F3iA
5fsk4gO5fumiOAGsjoISeT+Ps4oJ1FCisJ9bC5b5RzRJp7dZVqwq/+3jNybXlFtaPPOm5EFRGxXs
T9SveXyqlOqAImjKrS/IVAzfIXKtrRbM2XKMiWMa5gUsSShfPnSQmNCqzKAMnnB3L1fE1JMaw87n
SpwmQIOCgj+tMq+gn4I45mcdSaqx/TUHac9Wl1yrqe+SNz870Sn9Py0tNEIRh3cFgakDEnLua/3V
EnZbOpksWFB0pGCrhSrn7/VvsMoMfee6ODtfDt7OhDGiIm62Sw21UFye5+njj5CPijYYlDHtqyJD
kJe9qylZ/jF91bQgWaVOWJpNLxAAs+0MheXjs7TWErnRuRBwc4Ws+kSlIgP4YcF/mcOO0jf21O+Z
ydNWSiAgf4f4Gc4vD16LL8jqSDuUirv/2HX1U27wrPdSs6Ao+7kk+gcCcnN10eDvDLG4+5tZscSd
EPnQ+hZM5jnPeXCpWjy0KYZB30nLpARqMvYoes75XUJENAPhzrd7ukA+H/K95QshlbDL7w4czfRk
imz3SoiA35FVIRfuGIHX9XiBXkKZ0B3G87Dz7LFB0x/6n+G+kEPSfplI1fcSKqLbOXvuSan+TMHS
VSE1atNszk/tGEcMfkd/X9b86F0GoDWE1hBgdEVHTkQCjU0OKwnDScIhG2yHZ5usQrQipVGOfgRn
Z0boPto6RO2g8dyi557P/aONjPa2VBpRcpsyA0l4NdwD3OrvTP5hxzSRliPCAwmRg3Q4x0PnSNHu
4dB4oEw4SAFH9lB1JYlzcvo9M2jQIyrLrpEmHxo0eBCpwrrN5dxfXR+/D0eBkuNjFEq5wAQtHrGk
zMXfvX4+7jJCG0hD/xB+s+Gg0ehvfWrki7vZnDNUdoMsy1AKvhDuYry33fqHOacPsqf9T0sofpva
FXVSvp9Kes+j1JzoH+4YgQ9KLau4zEYfLG9LBwjb7+mz75zoztYHJ1OWEKJsoaZq6Fc0c8wlPdTj
1vamJSxapFoX86VDi5kyIzRpJxMx+DXBDx9Vo67nzmOQ/R9V7Fq5kaJqofjeF/nbla+APbWvis30
gMXVMXA8ZoR3fAHhqoBU1sKbZF4+OCgk9/9AQZFTjNxBf+eaL5qAk4xJZqYIa3msZUAJBOY2AtAd
an+ryeeRQoSe0F/4j9r/XJFBtvB6931KKCdNCEBmYV33hTmun3Xgp++fLBcP7e1bM5JB8Gv5+OA2
yfHi68dtMLOxyY98ualwFGWDJSO/BN+wiSTeJT8oI5URo3ltWCG/P0ts6UX8/j5YXIKermdURX5Y
uCC78crdfKZLJu75Y8OwEH45/6+QDp+SAl2jkRy9a9RkUkG9cqEqa15Xl3er2a88JxPHYXrOmXSI
dX/d0vzx1CZCaYud82br5wMHEr2NBX1cpXwoyd/e5+Bk6ewBJfTaQ7ATng85JSKVtZ3AQ+fFRuWE
UHzaso+fCaZiK39XablWFplIlkX2bCoSBItPTnUxe3eU3rCshcLg/gmeQiBXDiykJafH+MPiDI44
QYdUTKv3KGcUAPo3ajWaIfDeNB3jZXRbHPVVvgD59so5GPw0g8EC/8DXAvwWJ42RHccfqsobX5vE
J+sC76Y5WKV5m0wcUaCVeiffMSFAx9qw/ndi1n0dPf7vjtoKeqUrUT83PUlG6wQJslDLfLylkzap
e+WWq5Acy4LPJWZKbO9hJ5hUn9hsCijvEumFEmPXBuB/nEEoIdPtKCIeKDKWR+PjKXTZ6SWm7INb
WcpGWSzi3V4qbE6OfoW+31BPmp4zI4ZYTPKaLubUdZ2soN63G8cX39RLLi/tyyU4hBhx+QpKf1EC
9m6yn5I+M/PcaoRVbNG+dLiawu3Klggh9THK/fzHMnP0JWI6dxttUyhoff67wJ4N2O4a/trdwRfT
n6IUNF17GFp/Q6BpdE09TX7QZZyf5h3MmE8kQOxmV9UXGq/whkuGgWntGyAT8ASnJ5phB3z+p2g3
N9PrOnqdccC/lCwKSe7cMk8+F5X0pvvAAMvQDlFmnZ+8wXl3wm1NrIoFqH88u0SKaEdHtRzBUIFS
T7eibCDIJ5F3EbjU+HbwSUduhYqqbwbYm/ThHbU5TjOemOwHOp2Y/qNij1MrfjvPWwSi+o+lXZzf
cHlZO6Yd4QP3J8Eof0cebQgWscx5t9GzgYsMk4IydpJ9fVlvqlq80PrfUV8o1uiFfYamvHLH94s2
CAvhK0vdYEsYeL6sZ0vkvAUJSSDETkmby3kEGZ909i6wTEFU71/tocO+Yke38M0nNYxzW1uNFs6x
qT6aFdEdwhcp2fyQnfhD20Hcb8IDvfSbFLHfjuhQ0HkYEqHAmteadGy4tQUkOTN9flIwA0YskMb7
MaVvGXsNk2LbJhtqld/9XVNnX43ylva7cub9JBj6XJrE1i3+daN8N9aP9FSK/SVJ2lI/Vz/MA46S
DaTQFLtTUyCfCcTnQdhsEUFwD8fDLmz/GKSkbgl0tLsBjH5Q2xkuvQ2f5FcH9opzr3PGabPXc6lj
p6PZtYB72LC5iBdSHCYBwuyI2rTwOHdTUa4+forbiUx/6okbeM6xBc79myQz878RWSx+U6ikLdI2
et37VfgpOmCSCiX9Ur56qv64gOIZWmeNqAmYbKU7UD2Fc7FxhxJ4damIPo3iobK0eT4EdpDfl/2q
u+FT9tBfTeYiIWz+VJ8G8ippyi5j9Qp1P3zZTQBLZPb1FUyNHB3ez+7XFpNWBAG/zET5cyCiFTSo
IC9Ci186HBPRqvb1WbckmPow9LYp/8PrX0MCtXifkN32+sOj/SPwlqf3bDfB3mFXKAbjKBT64Liz
OyRPuttyf2Zn19wBEdSEy5UUBhX6UPqPVzdnfS6u1zwNvQcGSwwZAv3V8gQKaFljsF5XjVdKPY0s
lnGxOa7Vfm2IKYDUnpdSAbB4NSyTphkeQsYk5AkSnu3FBV2rj2c6T7IkRDICdA4WPm/cWUgqg0sh
bPXXfikXIyPHwXPjs583FL8TbNKFL27XpGDEtftFea2QonboGdga6oIaQLtGMiUyci925pJIaxw9
UbjLmHMdRnvhRBf9vfGtdorT4g5RHCeXvb80f47dQEVQud2oTq2BSNoU/MduHH3Supwx4qjjQM3d
RsHA1jyf9Eq8xtOYViNIYPcqkZIV+yt1Tl7HJ60LnMI01/EBSIsRsi5/mJTrD3eJQY18miVM/R7T
aJmertC+p7ADfuf9XO+vTK2XNii4dcaURdw+0XxDfIdk9mG7xNArcS4KNVXUpnIYDg42vv+FA0q+
Ujt7ljdxTFS9Qs/SRNXmrb9cZBRXtOIeAUeATdByipM3Ue9Yv0Re22aPi32UWK9koSs/O9UQWoFR
LBGvJPs/gtNdvqUkGejfXOw1qZEkKw9iP/Jgg+CvBzxzPoapjJhv4GUMD3CSjhvfqcNJedFb8UML
gkDWuWkPLxbFHB8jFN4FnRhKVivatNVXqhc59ggQFbNSncZSV/4ag145fhqGclkXbmhng6hdjoH0
rKEcUbjTHKybxdndGWrWVIQgRGFJj706RuWK4Jivpbm5fIkINykNVQ9l+gnUGO1e3YoK3iIyEgB9
aR0D7hQYgzuJyAFgRLO2Dn1JmVIbdnLqRbyv5GiDysa3tcytg69Mu0qQo7inns5DrvBOOFFuTpZk
ZJQdqqUnc9TaK8exnAd6BEz/PwKmYGUMYaPaWm/4fZD3DJIixI/bK1RVP90GE6dC9o3/PU6sxYCM
fNOSZgl+Trn/1QH3vY6PkhuD9ciVze7gX7x1Ev8wvSBHLr8KcGCfri1DypSZkPpfcHFFXAf9+REl
IfFa4jdDJo0y1VgAnnDvBGaP+QJjk8FGXO7mwoneeUktsg/wTEsv9jr5LsvmZOqvz782cHyiasux
bB4anHCZJHPwRFONJ25ScgRZEYFJiNwkuJMryMGKRieWpE+ahscWboFP9m/W6OUAz6NhcrYyfeJz
hXeZ0YKgVbTBw1RVF4SgbkD5sJ9Wtk+9UHiqUcsa+2pukQ+BayeYIlKPBWIG+rAWNazBsksAXNAm
ynEsW640oYk4VEJIAv2K00RtoEfgOIxnvT7MZR/bTcRnLMtubWUV1+26hJfo7MCMzc/zRqaY1mPU
ZKxOPYAB/ubuxZX6+/Ex1vV7AXSCIIs3cxREzM3QAEiPNFoMlpoZikgS1z6+uLHZBs7B48z5Y9Px
rlqaFRoGSx0U9Zy6QzaBELqd+wZ2G3noCbePgLIlvgQopSCkr66C28SmfK2uy95u/x6DGIwpD0LB
JF0Phs3vWXyU/d2KGEkwdWwZLtp6Sv39fGiE9A+8bUxiwaOdNl2MGYE2nioCiZxrbmr6OJJ7mP2S
wS2IhxyBno+O7D3yc094wNTl00o6s/d5JdeKxhqssWEpMgdXWdqDSFZbfbOROIPju5i5Fl7WQk6s
cYnlChJZFplhgbboZm35CBkJxdjQVqeg3gTQM1oMXCD1zlP4fqm6I1DRTmgcgGtEVMBCJOeZ37Lm
Z+XneVTPTYGJ0g33J88wyneQSsiBRjSiqJynhcoT58Hd2678InyCeDmuXHUT3kN7hjQoNiDPkOKq
++gljRTZNVMiLHRX0Zu+aM6pwwWFj3dFqpDKlAOSQMd3wXUzEcZZS5tAv0UnUuxfvidH4W2Mcafk
cyHouI2ausj0mIFlecx57GjPZmyIzUwLF+m1RBD3jO4xa3MrD4YUqSAMX/y13vkabyjNbXbCEguw
a3SkYzPU42v6YT9ctjoCHkGZu/HxahIF0m8FSoUe/6GMFzPyDgO4z96ATBfCcS9qanslqHvqbe4U
1E0wMDiqWVZvrzapdVcc3ZmP2ien8RWxBVSugHEPnYqr11XEjV12uowLm2zLO23nmYjokoLjTOF7
Pvyf5ZlzL6yNPOzMl8Gf6lu4wksoLtvSZ8lFdRSbukTn4Isd3lYPJ2xxm3sRurGOCQNoxyY/2xDf
FdzDE56KsHfFHU2fnRF7iklYZWsm05ykxUwyr1Qm2gi+FeQ4z7koxkTpOzdmrkXiiD8Qy2dwYmO4
vlgyNJrxKteJSpCj8Al6gUTHj5Wct2yqBH/YrnAwkE+YaOjtpW6uc7JgwrZtVtvZ/fWmLktJSEUn
AvSNE+mJpLhbOxWHeY8V10YbdvaFMvhTaIhNyyG6HICVy7mo6iuWrGwOEG9KNCg5yNfPkxWSOFij
MwJ5glURqXK9JO01x9gKh43vtp+8j8jA4B3ZcVBzx3qO7gBfzuyxXYzn2sEe4TVCSPuIL76flpjf
DslDvweN+N4U8Idn0MeR9pyudk1TpDyu3iyHN++QYm6TARschCpgiS3BHl76InV5u3+70H/R3M7B
9fQRAIzLa3VZLiAXL16wAL5wqjptiQSDmDRXIaKtTnsNVanI2MRMVjwSOpdSiCatYU2nDyBxWytC
yq/XRPKetDXrm/hzE7Bb4kYdNNRhJKCp3UOjOdiyipmEB0XJ/WTaNGFiJH/AK/UEZufarfMECnlg
EgJzDIerOIfj1V4cG16J2XuUWKA9MeT+rM0EIh4Z+XObIwAoX4VD1bkyU1Zru4Hd+5xey9D6xQOA
WOKWFAuzo4vNadtM33sfyxO1+KJ4YClO6mNa31WwWW6ChO5RBx2nPvPFyRl93Cda7enMcrhYmd3l
P/t8g5YGrEiLQckCPoMMRVAYMDjc2hTZwnBb23myTr1jEfvykdCZRgdxgY5/k3AdX9FMJN41QaZW
HsgPujihbKpWwBjkqfGZrwI2A45hYAD78cZKB3Nz8cFjgb6vtG8gmOHfr8yDgihcNC2sXyRecokv
Ib5/LSMUT3fi9GcQt+5/EVzCaJiPt9oCAhi4NRGZQnNdAFqw5krlVPcNxVqpXyvuZipgEchzSUnP
vFiG9Lef8TheRRhVYCO8NAXN/ojNYznb+tIOH9lrJeAlz9+XH/2tT93TGPmPb4evIQ5uo14oLHOL
TO5eWILIsQM8qeMcK09c54qE/EHJ7XX708JJnxels6Dcrh6PRUsud2j4jDGysfdVzf7n8y6iMb6i
HQHOIC7uuV1hiazCPAAQMH5EtgyvtqjScP57r1DQxP6ogDw1Avp+kJO0zY/n2NeXKuvl+V8gRCe3
3PrJlcd0+x782Vw6loI2axN5s8bUQvP8LNU78Z2RFe13bQjw12WCuULcneS+yeWoqAChG5oy81At
HV0WtiGIrEtXF9UZuxqD00pvm7oozTTx51/nsI/l787DZ8f/+R+Nnzc/JR/iAKB4Hn12IOd7wjVp
GHAUOyorrF2k+vT3uE+Nse09MZmOkDZNLQpn//ansMJonma8PUSElNw0YA0kWM/0tFNgRc7g5N2N
V5TTe0TxofUtmf17/uMvxtr9FDG9dhvaAOUtHF5eBt9kNaZ3/HZFdF+WN00N+M6SEZ3FGiC4/oRy
uh7REfQYseOfrBLn86WMaOsIHHGfm5PqYhkHLQvmrljCvIRx/a13OORXoh+BRkjMwRf3SP3ZCsX9
rPuhB2fFVOc59xJkOHv3WDl2KHE7IFFiyouQWcGcbl03K4PG5qfuiexVdJWDbxUhZJyQ0BSQrp9c
jyJAU2/t5TM5HuNMfVzziFkPakCKejoorYzxmtHjZD/L/BV7zXhvPjTODKCH2T3bxWKeB0dXOa7R
ZVcJtc0l+Kpaz2eTrpZhxgyNxdJMSRIWljn6Ig9t6ZPvNc2Du9DutRVqWg8nC3Bih6jSPvfICB4c
VJ6evGXiIQM5GbHc3jxCDNtQxfj5Xu6YzJ9EYdgtCDTl+ZK8cWco5oOHSYTrt14ywfk9c22e6gjE
y/efP6Z4J4wqsgULnlbnYFlyDxvfyUcwIwq0GWnoGSM47bVYMA7y6fdWb6oVYHsecv10S/kUagzD
6pjleP6kTzQfUG7Cmmoy/OfTReIb7pEQUEsyJto7gRxao0raFnx8xb1b4GbuAIQef454pHBPGNI7
nESAlg+4M9i3dDk47YiaW3KPPzcyjMJKpwM9VMJLbmPxY+rnr8jfURcaC2M9osdNjfA84kf/v25q
On6KBk1pV6wypLqYZ3tfEGRtexFUz78J2MRWOdYlW0F8QFTo8vylLLzvUp5txmr32L0a1mnShXas
+iXxi9jLiHsfG1VLuKLtCq7k22T+tiU3526jCGG+v9ZfzOvLKQzONMMqSWm/m8Bb5iukI7rUgNfu
osumoRA8IXVli5OXRIEtn4HTyOJhn/5xh63+UvcY4eTjVZN+0AndIVm1J5OOyLYzhuuKOZRw561x
4N8Z+aoAQM6fnVyhYxBtv7FKZ2nTQ56Z2I4dpSRY2M2L+ksXcPauVXbeO48m+mxhTjMcsGBGGWZ8
jaJB4EtIvNRYttWk5F+BmA41JpxU1RAAm0SXlmeDNs6Q3+dcL1qK+zYXwQqXw+0OBvpo1Xb/YNl+
xenH6vI+Liq9z6jE9s8XKXhyyzvZ0+Yv11Es3ps9PkFAeSQLaDpwDp26XH57M7iSn2IYkqCa96Fn
s/qxBP8gimuAw4aNhcXpMYo/x/4HblgmVk44qydIjLoUgivNGqp+9eReoKJFf9teoTiNIPW+vXuE
3RQQC+YLJ1GI0fxllkNqVPOKCSe4oJXadOWmRaMUKs38ZR2rPky2RvAvBpZ5kOqw/xSqR3g6mQiy
+K8za1ZQomKJoU95aeHilkU795PdBCmrycB5emJBsOTKqtm5okEdOTCci6NO+CyB3RV7/0isfO4G
ds2JrsZt32ihSuZCnQShGyMTpcv4P/8+wXC41qk+1qvmsUWeC0M7v/XdgNtBRjcIAK2zYgTzny4C
xSmUWSI5nbhsL19Mnki45jXVtfkG2yOpekgnik8dTJbI/6qKX1sLpBKA/v3+BCJ2NTqyxxBHmvdj
Nd9qOcccKMEBseYdN9sjTy317/MmqaaV4SwhPo9MNn1eadkT9Qeu6M7YWz+DsIJmIEMrRyBochgW
/lbnegCPaHBPt6YMgTz8x6pZ9dODeqjGgPk+kquNkkFa5wnNO4CCfxu5lBsScYJ7pdgLKpoMGUzZ
oTQjkjWuJVunENToEGq2CUXrIC6t7Kbv0REsPoFWb+pbHzR1UFjCOZyS9gHZUnvbwMd47mumItNq
tn4zd2ANmkN2mqLq87q+BXQmqfGYRswoo/8D05nn4rHy063BuEPUfH6Z31Ox3dInM+2IEbs59p1j
s5KgNWKGNTH/BraPqxtoJ+0y0ZoDrRvHkrzJuVx2egquQ5ZTU7DpsPXhSmZoyx+en5t7WyT9mBv5
+BO0aIzzlVpbviErZnbRHXr0BYKfxDy9Fp1KnjPhRVs/OPy6InA/KxM988pljmidR+paqbDU9m/k
8+seYRiCN0ZU/Y00OeanYIhMa5QAHmwJ6yS0ECIfdoEf+4L4xVekQnnt7vw0ayOIaHOWS1eY2F6k
PaDq/EVX5FlurWrEh6qV/HQO8g7FlG2Dmjf7pj1c6gi8ZTJ6g/VHGn4i7eOM+loWIvBlWHg91X8+
RdoylxffzmcZHktq1DM9y9PDdIxbAVtz6OIRCVLjP6CpSCIID+NpexVne25AiMOIADXDPAXQ7aZB
ozd0eecAidaPah6Kwv80NqYGwoC8aDNl1LdDzTZoH2P0KujhCDDz18nDpkaGunVwwf8mDdDKKNd/
pfSbLAxL595W44pQQ7TON0cgCVLMF89w0u0WuJ703TR5Vt1JY0SnnDNgI+2uYhQvMfXLpeJlYnee
H1b9pZuJnfLNN8+6tIXf8pkCXpIPVMxRg/DotNACq4msRKtWFSn4amRmtzGsTf/8jEjbWa6GhYkZ
WX2Djzh6MRn4e5oDhZnHPw5NjMtlJ+Z+qi0Pekd3XWFcaM0sDyNJivIOhU/RGpwdQYvPSy0OTpIq
0E5XV9XJC2JJ8JvT1TJrgkOR7374NjnYlpQIbugr8bMzhlryClytDloUKDOsei3+HxdbGR7zNH/A
HbMDSFWxDFl2kBAfOn2AU5saA0GWZnTnZKUPZ/HooWSDDtGIjXLQ0b1dCdpof0j9bJrTDaGegcFM
Zs0eys2TpXeak63UMYwwsc07BIR7Za1wYY/nAcBoF6kHvo/sX6pVr/HrTGQXtu7/sGHJhjZU44p2
BnW/1cAPEiWgkxraoi/Z1jQb2+QYMxAlqtmzQJYZA5vLbaKj6M3Ij0ZACPuAGj//WGYOIIoraaGv
69354KcF399blsAhbjeB8ynYIPErCQ6hS/7aGJ4XOtqVq+r9jeHurUI014X6U2H7j5EsnV2pRQfp
QTXoUD6/APPrcreACThH1uSzFLW+2DzYekZrPhq/OWH2VRDPBO09x3C0Lk+aWENXWs2GiHXsnnP6
exbKy7cp7/yQamtvRckfKonAS1i04e8QTyVE2BI5+yDB2x3ELL77P24p1EzcN/aU5TAeqbCvzY+D
UwKTk0i0gFMY3wH6MqQ2M6ItsLljfQhMk/NYg2xYYmIPa2wz8BBc8y44VDJ+6PQRi1hcxPscrjBf
WKcJyeCjD03VRMXGPmViHhtPQO5lnXYv/EK6L5h1u4mawgC7D21ge9D/TQ/Ua0oz7vBg/gU3VW1K
b/o2GCTfXPLO0mSLpUH8vC2XQfvMv8EeNRFUMQqIHybfXEeVSIhM1dBsPXL2MAkyWWtcIVYH3DOt
rmHRcFU36TXHta35cCJ4JsNj1I+JV5Z35Kpa+GXu/diE8CJnFAa/eqjwiFkU6SQBvb/0Lp9JkxZX
BPWBrvzOdGgFesnDt3ktqea0RCflBg5UwHCEVakb8VO/67s+8MAfqCb1vTE/JcRpoPayzC0CSM3r
WDke1MDt1DyL26l3AoiIQFEpTWdj7md/ZpKmoIMpftJpWWo7tZvMFNsXQ05JTbTdi0dj91irI9iS
aKVwgXr61pEOWZ2sqjSUgIGr9f3zgTZ/AVkgdKiJCtxh30nJdgr74b1YZfXp378U2Z6k9biQ0yqn
7yoxCImFgCZ9rbo9+5fK/+WU0r/Rv2I+jIcqj3oSrT0OLno8MLh9rHmq1S9BetqUkn2Tx6aQN9Ng
YY/b0qEpf7o4Eb9fHElTL70SMS9z/URoRzvdahjSzIqBTCDQaJ5/bX8/QpbK6Sukv1+El+SU2Em8
qAOW7K6Vn8kvpR40Aw8sPALhJfWvPOhVS4yT8kI/YLcB5osCxoMTKNTpxS1mUQ9arm++TctADvbB
E8xs5RirJ8nC+yTK+hR0Ss9QpM6zFUywn6LB9h/WQPOWCeWDTo9d+2i2+sjOjyuS9Xf1shnb4xJl
lfawMoi3EMz32/KiCfdimyuWqC0hyNI72110M0leX9Lw/5irFvIIeHKeiJcmj3gR4O2wbGfTewY+
u/tp0cy6OnFHwE+IxRP1TuFc9+fYYooP+4uuLbm9g9BWul2lQda+xvIfnUL9vR+//bjm8Za1eMmy
9vW7Z3klQh1/1jngpHGaMSXcpvgGvnuyqglwN2q0ts+m/8MzgUM8C8m8Xyg+8e0Mhi/9ARgo/3zV
nH5Frw19tJ2KgOVfJR1vOYrspjo2j9+cA+xesxa6SkKAJ9+pAakcvVeL4WTuymectkJTryMIiPE8
4JEeZkntV5+PErIoHWlwjDWdlNr3EaJLgEuqZRM66FNPKE+/XboOhQ2Id3r7EjYOxY3jZbjika7A
5GuKFFWhd7onn8jT8Bl3ZAWuNmvw8xPeFYdDIxHXl12MSJZ/QYDZ0Sp89JvjQBXQX0mXiSimwDUP
h/ofjjGvyNYU1djcR8oQl+PFfPhhegBi5mN/ZrjH4u8BweGpOgVGROk4QwTnVZN4t38PkYSn0MFa
EOT2NVggQg7zcNjRyh2KwSqNOq0vodvdyhMyLXhlb4lchfp8U5jMNFJfSAbNyP/0RKaVxEitr2om
6HLugeN1zm+peupBCI/GGBlHJ1er25v2QNuoy+41WR2OQ0I/iUzq5OP9fdOXR25kFxGdO8YSBeKl
juohzGOnWIPZe1cBY1kWAu+7HkftKqDNrsMDZB5f8o/pD2y2bfovLI05jmqh4wbT08Zs7Ht9RVi6
RKGGaaLZTfSWIfBHYMRzoDEoaNLuZQHZYs2HEfpove8I9y8uqTIdi/sj3mbUgu8245qA/6sVzYQY
o9ELdpYiS3NjKGmLQ9xZ9rKRH7Yawo7iUNysgdiQIL01DIcdyjq+ufJirX/8/aNR+o8uosF9+WYa
+FiRDEZ+tJfsF3ijZogodUpnq1z7vtSm39b6f7hjYus+2iFuceUYLw9ERx5gSvrqEKlZl2V1xD2W
urjw8WCqnqC5I5rv/jWv6mjXoO5OOLDEvAXNKTiYe/q+dxJVIxOR+k1Z6y3Y3LqHklsx5SwUyJyS
+4gHHuGG9t4fTohoGDdFtsR5AF1F599N/rOMo2YETbjc3v4AelgqSF54vjIu4LYzHV6XJ6Vopqax
c6GmH0sF1CjqZUjdrX9SXWf6CBze+2VUenqPbAAzTwO01Rvxrp7uGGDN3eO5sIfbgIIhvZSpNW+b
oX61oKW+F0huXotY3k26wkBrxxAF9ONrdSQ0DAI9wzO9NMFow5JaoPaA5vnRMiTGmSLitXN6aJpr
s4h+w/HB29v2fwIm63T81qy6WU7WEhfEM91m9Q2MD3FRyBCgWL8IhqRKBmG5dUk4L4Re18Rs7EM2
1PKuDtPwkKPGct2spt3cJP/Zory/jYJSIjEN0KWi7fHsN5OKC0rMucxCmG6AQfnSqOqUJ+ffFuNN
08BDww4Z6cg81J6aNRpszhcREzLxOOVQ+qY9mM+VATfiGZ2s9R6A++q5/1EC/hMYuQNerbbyAjqX
8/Qf9g8MDlnfxnvcA2YyzQPj3aCSRd6uPVT+HeqjOjnZjaObgVHxdvdyTOL2EFkSZYopsZ2iN0nJ
fufZBQpIjEPp0y5I+3ru1n6kAnxQQq6O6ZvVt/i7k+fe07pR2dwP609g8GbJ2AzFYc8cUYKp3XRL
mYw7iYkHSKn9Z1nZAWXIhqohImP6+LiMWyW4xa2Zeo91f87+33oWiqaFd4aWlpFxL27kROe8OjMp
gWqEL3eDosUnqBX81/xLIcvAjcTumNgUX35pOzGQQWcF7vgcuHAUSYjV7EHJbSo8LHyjJq+RcoxP
90/zPIVupBI9+sg9knqKyoW6W5PRyPC4idENTPkLwql7KxBkjq4E8jm9/QRHyIXkVWXsyw6siO7A
cwBng2oW/B9II4i5ocRbOYwPxa1j3khNBVE5ZhOLQ4jvO+KMshTNhy1lliqoYzvg2UJk0RLs0jC2
9g954M2uVMAONEA9n0qWoR0zHoDALTAbGb4AIqDyOmB7s6U2Si+BU488ahx7B7GAQQcybq/F6a6r
3K3SXkiOYbSWlySgW/8AL/+DrXWzKEAtzhMmUJZYsdcqspu1g/GQiOomJC2TbEmo0RRmGRZv8AWq
8L/Q15VM46tO4nEdey6GMYPzfas5fzPaAw+0d2qjuWZLG/T48PVI4bl0UMzCSqfas11vs0WgnlMp
GesU9uI3LiQEp4RbSajaxySwpZ7oUSR7pjG6EuR9RrajHTyvhbudy0UzpcgJf4WXwvxKI2D6Lm0C
fMQCprHSlAduwXJ+TppUZnXs4LIieLZp0ZmBl/mBa1YPzZ9ABY7FuYP8IRtCiX49f8bEe0Yd9mOL
pVtNsbwNBCVGzrHCquIO4Yoyb04NMM50JJ5ZHdTB1Y6BhcnqZ+6itv4xCMpggQQ3AGfNTxalc9dq
vCJPAhfliNk1rySi0zClnTfz/3xMo1/2fThSUp8Uv+DKnfpjlYe+LOwlioNWsJXlY8D01cjyV7r7
fOYaGmNydbow1wtHFqtW23K8GYXsREcgEVlF11slIPefxW0YoqkZPoU2n08S7xas9GcGBU7rRTvH
stjDwaPX/HXyXDT8gqyiopQuj+G/vNn7aqace3ViMQWL5OZDrdKTQJZ1kvnop+lHY04Gy1pA2pEJ
87VzD/2zye+jVJsf4+br0y4hV8h2ty5bNT0OHEJUCi1dxmA/EhwkI6X8vkr//TdCaKKQ037iS0Ec
7CiZhAEE79H/ylVjfDTiNlP5H5EqHfFnKTYHYUweSUIOEn38CEGoA48pluVHhnUof6z5c1jlaQCE
XE85ccfNyXGywvT1xLq17nVMILn+69jB9bwF5KEvLPO6M3Tg/LXn1IxhC2Jekw4r7nzepkfqn6se
SHAhX8b5KCOvwF5p68jjGoxYc8pMk/X34UXiArApyBaI8yQ0xfXeSRwTRtSTCwMolVFC/EPQsuqF
tBgxa7BP5p59iwdDYpsz7uFO+id2AOnELyTkM0fRYoni7myFe4s+EjWxMrVV9c91z52D6AYWEXYZ
3eDl9l+cpXKto4vsvxbvQ+GyEySoQd+LTX8+rBmfGTr8lC/dZ/CuAiFz/9+bWcIoONCVL1i9fR/o
j4VFVpX4kRqS3inhtibobzvs2TYRPISLGvk+0PMkgte5fK2PpollnWsp6UnLVJmwiINA2VQlElCt
AO6bYGkWck56A6D/P3LoCVWCuq5CIMbHxX4URj/In4WERh7cTM/OTcmNgSo81Oys3suJEdNFdRXl
6HqR3JHQMXTUGBARkI7ewJ3wkEqsnO+dYMP4O7So+RCcCY354wAA77yNPLT+mhMXjpwsl7bbuTcC
XMKgkfRg1szUPb3uewF+nWrn6lVlYPsqTIV0FTVoj1i8bne3DK+rsgOhoFsJ3VxxvGQSEU6c3klO
5yyAYqc1RfQgLOJYCuuUz+OMuX6p0CS2nSbv9TnlsHCcKAhKpJ+NicUbr+IQuhliDPmFIcjyL7go
I59wLGGth0wgoQc4UBUJTLwCb5sVN9G0i2f5ODD8bwVBB1zf53lq0MMFKmQfbUsvVYP4JP/ISzL2
nYFJR1hSZArvzOgKs4wVrSYiXmg+hCZ+awLjFxH8NEBvWnzCJ6+GLRLBdo0cYTTGBwv2oVRjfnAG
sQ3nRRc7AbUxp7epXkbflwzuPGsAwo17ep+M2vx5h+ck0dpOEF8ttWzsx6OFQ9WWrFsiVLddUA03
imHD/ZyYhUC1GQvsm0CHVMA4na/f94IAMapORCg8da8+WCt7ykBk65UbTk3hexETdtxl2zT8K9j4
FIkAOUi7wZHUn3RmbSCzz6UIt6vnNZ5+wl4vZNQgBRT25t2YF3VqPW85J0wb74rEyvs1IlZC8EfU
D8lLrXZmZvX0hZnJy3+rKH706VL/4wkib/p+aKA/Ws0SNt6M2IsJYuoFKjQ2jAdi++jPV5yn45p7
C2hFuHTHqurDL3/khhnG8aNhaBmuy1rSj9P5upItdHcP+wg1h+/6KbBgQxJ3Pf/cH22QO7T7wo7l
OyG//gfZErQyPOlBTwG6qb3nOAhoS+57XaEWCjDq/rv2R9zysIvf3GXlF9/s8+DLIT0beCv+/ksJ
DtXhhM5d9aqECkU5n8UQGzvGVJZJuLPguViTSfDWizIXoSxfP/Xu0KLVghVL4JjFJ2l+OlLMKZ/N
xlt3bH6CdlYYKaW5zeo6Qdx02IpbJnOEcV4mjwRU/WyU7Xg+ivVT8m46J+BfB+7mRiTzBxUCL3pP
OXoGx+YRLYolxV2j0iaUt1sSNwn7dlU3A3ZPD8ydMBELf3y7DPtmnpf+YoLD2kioTGnfk++FMzQA
9pPEgjvseN5UgCZvjMpccb1WRmN8Fg/DpjxDwi3Rvp6NvWUzeIdBcjm7ok9ttx8o7j5JkfFSDEQT
8z1w/j6K3lx9EAhX1XV91zOP9zQ/4KlnVPoiC2g0KYTye0dOhR0+EYVN+HvXAIn+DXbL5WiycZtO
w5VUuT4Ovpb41qISl9cdPHur8jF3fwIhVJBtvagCG8td8IE6X8VyMp63X7x0DKTcDbkpzFQXtkfs
W+17EXCM0NeQzKkb0bAxAtCcZB2zX8QgedtAa9p6xJkChxvoQwPOaaCjzDnbmJI9SrXZ0FS+m+y+
3DvzQ2H2da8liTAgfbzUWF/pLuRR9mKTLXCUxBcBtx9IukkUMrrWRA//7tAcArIgUKLX0byvLNJF
FvblZyN6aSkiZ2TzQ70bDCEUWPde6RHo6jNj99YrN3fb50D1MDYyrEGyLZYXOEBHGfEN5HpxEheZ
DeKI1lyJc6e39JUYYb4ELbh4Gj8saU7y1yeve9oNj/SFu8R3XdOefQyLOauQ/GVuOAOfhD3jACu2
PcUr1Mhdfip/zXh3cWGj0PkM4mCUXEDlKtNhC2RczunIm89/dApfTGXKJ3eKoslpGxrOS402tTMI
W9A7hXHth6JPDcyMD4P4Ul1k1YQitmMoELigzxkw0HCS9m1fc7ws8yML3tYGso24ZG7ds1NwXy2O
bWNqHZ33O7zrCCbKMDLwJHwBf90BI4tvWUMpU+WLHTTSRDFv2KLmOawarhMcTIOLVI0b69rOqqMD
7quElAcDiiGO5q5bWLnj1QYA6fZ4hWScu9DNSu9IcMdh0dxSYC7BsYYReG/ul2l6JeS7XbV5GtQJ
GZdzfOnFXCkIz5e2LsNCJpkiu1PQqEUW+L2x9S7i/wNHV7Kt0q+1L/mHMRNCQ4r7kw/VL9q8DKs0
2+WN/Ir6tmHV3flEk8oTP3nPIJbUDHwLIoA8Rc/yrGMMUbf/7gnfQZZ/WXoUbN9gyRfSTngoTbcN
uUQlCQUJopcvAjoLS63SFqg4lmHhLpL1WkSFdbcfD05h0eHjM59Novr5wEye3D7/tqToDyOz76jK
tVvDnfld1qsAkD+zU9eRZx6h6VlEyImzgqD2+G7B/xkFt9BbmuOi8UK1h/N1E1Q+UtsDpyUtoylj
GZJB/7Smm+SolhUNWpSON4pIS4fRsxjl0gTOILvjQkzcmEKcPDVkCXLxUuK1DuwBJ68KzsRV1uUE
KPGaEECq38S1kD0mrJs2C1kQVIu7xCmF/yo7KaA0oywb+pX1HvjMAU0Da9CLFmbovSfj3IXwFL8t
BeitKctR8hFShOYMaAAjEyomMAUYtna4pRYT7tYvXfHKMBKB+ZpUUHB9N2mzeoBraZtVzoCoa7V/
nm3jLzdG3KCHMmIvWDY0sUk8sBnhS9on17gZH6UutF1IrcdUc+D3cGTDklvYh/3CH9xZTcU3LHiE
ZIHD9xh7nnYazyNAOUNw+NpJSDVEW9KLf51LYC0BiwFAlv5cjUVjfOVblyiqTBS07N16jCoz3ZtD
sV/wZksRtYPvU0wt0iZeC0iXJZo8KQ0nfNEY3tWgjtVEIcuQN/mCaUwAdCKMz0R/lN9XQ/NU8NrM
6dx2GY7HF+9EYoLnkqW/x9LQXRwT9Gmo72HeFnFm/tZo1olPxc8/+Tc16PLc
`protect end_protected

