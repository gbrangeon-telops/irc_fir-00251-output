

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SOOYAbmSVdMSmEhVcX6OANZAlRBhIeIgp+j8aWie5qMiZZfkKWRKGFlDj4dOK2MxGgpLi60kolAl
iwo8CvQQmg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XO8hvx7ayNrMYNs+QowHbS9oiS1GjnY7XWvxUBWvS8S0pBwgguPJgxI5Jawjx75IEBra9z6gur8D
+8bJ3wjB5uOzP0Op4TufbsYZTMy5/IRaR1m1haAiZDNWpnRaJY0iGIl1ZfXnFFB/FNm2d6rg/H7b
+K1wV2KmxNsYmhxGeUs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qrXPktUjITPZaeyYovMGSvjyrwEeWSEPCoXArB49zu0J+taotc50izauZkw4BvtuT10+TUqV3pWu
H2Y4+wBhbI0avNdhBTQ6WysNgxNkl4xSoIMSUDeWLPrThpvXqf5EM2xFWnYEsoSt1fOlTzsbNp4Z
xTF0/8eRzGcTqQK8goNirFS4li1yNxnvMyocM7UB0Hgwd4r1WhVfwqexmsE2F2aKD0WceDfUKvzW
BkaD/pggzoFKe9ZBj4krjm5QO6MJe6tmyETtklCe5Tp5KFVAoUG5SSUacYfOW5JRRQQN1B29KV6+
B/PXOjnEprmrDoW2/GvnZUOJ8iICUgvcDDx9Gw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RfdpJMuL5lneUspdc3THLHWNRfMy7ZKvo7MAlgXNSeMyJ16shj6csIbQx7zWlYY0s5cmQ5qBeuky
S0nRybRR8cWMHwN/9rEo4V+uesao4mJ5GbtqRFTH0pGXUIW0hSA/qLXBAZCtANiThLFmTTovXGQx
QWChhP7QcQZsZBRuEUY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KfAPtRUOpYg8KaNj0Wxd1r4Bcs5Lt64mregrxrObBeYBNNIje2iGcuv2d5+PQzzomKwP4NoGlbzx
CSYz6XLlhFat5X0Kad65Lvso8ilyZLrxVgz/cQQVMyGtqJsflyi+jbqMWdWQzDlLboEzDolIGqLM
T16l7bjdTv+UHoBJFQNNpgCUB8RCwZwGjuOrDkNOQRBxFbXP4ewZBD1TITGRJ+9yag2oeIszJxFS
OnxOibAvqbpn5K7zetHoNiQFD0HLxODP6ACT7OZWy2QVwDRr6smLhIBBF+7E8S7up2WgvZZ778OW
7Swo175PkHbmEfmpa+y5XkNQNOq7GC6XNCURkg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11344)
`protect data_block
8ouk4MdYXRg/vxxRsxM2cYoIDCY7jjSJo29PZKdlfJV5TsI2NakRhsnpFgyBtp+/LnBPa5ODomNS
LMK5LyIuudtprObbiZkFhrbqAXRVCMjtzBMEnSv61+0qHOnXOkUZC8shOr8Ika4TsnNs90wQZj55
8oc9lXhGXw6q5vzSoMNjBZkzXq0BSCD6NKWkwECwQhw+08uditCy76QeqyThtFcKOepN+JCKsB4i
EMgfB0xnAlJubuctAWmcWaIfj8BnED0Vc0bZuEhjMy8mCL8JjZ/TP4bDbSl4TuWdo2sJIGPLLM2c
mvH68TjUFCmOEz6FXOZ4Tw99nfRJfDrHOHcM6QlY7P+d8rCg6UapFng+BKGoqrQKSh2oCvn+0kSg
CceXky/LOSrTNFZmsJzzFJSkeRRECEfgdv9ZyM5P3JY2VYEHxBBKAAgXhrlW3b4TEn4OWyIIHxto
ui68Mb3LJPaQZADw0casHQC1elzuEaS/OoXSNxbn5EZNDokttxmZCet36a6XfY/zrioyueF9LW6R
1uHkKtDTTE5DbYOcLs1PmzeDvqGhBsgTQf/FT0+fifgWM4/s7YnQN8Nw1EvBsgjHtjuG+2/xbFfN
T+orEi1MY+C0h7oxTHDfxwqGb8x3I2alRKezDgIioOGWxnQJTyGDzh52aVZKU5PqpT2Y1AQxnXIm
DlCnf0a9nEfXUWVqeoDqY85KOr13SlcSckmVAxw7IJxrDRPtGkXFTiYKHScvNdcdPklDIZGgCo7Y
5fPWLkyssEuKXwEG0Q10IVPfG6QPCZNfYD7Jbezx8iQ/TdtHf140sOjmnMp1mtfEBOE7nwIpu2hZ
PmDicV2j0F82ZvDVZuJBpk4GMGRSr2TanL9YtJj8WBvYReabIGwD97/Rb1cQHwr5/smzX+pIpdrL
fvTRy06ERZadUgYpHiULmXbBUXwMYqur8LFKDsyC7HUSe4036Tb6GBgDK8lV9zf+MDn8Btlupddz
oB2wJpJV4pq7E/CUP69u/OEzKtmmrQszKikMv4EjOqPQ1+v+zeqisAlbqtOimBTywYz/Wfb3yT55
fFC6bwgigqXtl/pYitF8v9Kf0sTQGEM+b7b7M1YIKYM7pJFcTThFV7YO7a3POXeFQZnaXULmjibO
7s8U9dMgWP2B5wNZAyh16llz72U0T4d2FSUdjcXfj4XT9RDMV2IB4gIXYDkFsnKDEwlUULQdrMVX
uHlTTq56hR+IvIvu1OOR1AUiSVCgc4fLXm3Kk3tdWDPUjUt1kTjwWLPbrc94Oi9sshrkYs6vMSKE
0y27zOOlbL2RHejEyoIO42ZDRJhVFrAlk1HI+UrcbvxesxgxuzqRUmHQTw00amQq7OwJJbhcMTL7
HEyTsZYeAt1MoMCxGEbkSAPYU6www+HREE4ET+Mv7KNqB2wl7T6fKVW98rmywTjf1JLhgUzkW4m1
4Zm1P6/axLBlwRxPBDCVjjOIvjvNQ2aT6hZuuFUhVidC70TvI47FTWbSsbfV5QB2F6aahW1HSYK7
hwABlEGvm95WGb3mv7FPoaVHxvnYAgUD+7XNkP1WQYpigz6z7oHJL2JeGEL9d1DcSWQfrusdQgtR
nK/bMgP0CQbD9o9Yrn4spI1um0WDrWcF4zoL09/zuovrWGebsJ60qc3Tw8MCy5//n0SLR6xPNfm0
2IB9RD4l8t1VTmsQgW85132eXR/QUH4vAfnVGdoUOcjCRRnYPQy3VPX2ADJ1rJbMY2VN4fODZ5vQ
iBCFx1CxbPX4Yl3n6AFGr59Oa76fdM6UwP1qcWG3iEKtwW7Hs0IBGtPaE4Me+mYVxB3mUCcmAN9f
b3eAKUf7UzLLT46BKNR3JOqMveXV/urgC0U6wHLjkm8nw2/fW8sp1ZU9vKyGfTGbz1+ItdJ24n6H
0qSpJ8Dp0cdZOpbAL0ZOpFkkNnF6lp/gOjRRjxCJucLFh8NvMTNeei80vuTiZg0NQZNOecCgYqtY
X+Tdzmo58vWOileCo3J90vDHivlUnwca/fpxH39dUGQBkwDBbKMB/32yLG6eKlHKSjX64oNYp81C
Lexkuy9f3iCkci89skyUHaRVaHkCM/A+nhXZ6AeRcZd+HKHwNAAs/tSUjKhefbfOVvH+xvqwmGgu
2f272lOOA2LsCnQM9rXPfO+B0xAjit4TyVGCU+3TLfFUZA5E9DXL/X/VRQfERgZNfElHxR08p3Hh
WGFaqeY2llyaJP6qVvKpyd6w0tpuMR6byn2KO08pZH2RUP98ARMBkANLz1iw4MBa5oz6/z5LS5kj
Yril9pbJDD0hmIrjolY/WpyjrvRge7ntYPgr0aeHPXhs4duCRknDItHi8d+DqZibxGLxdHypp266
4uapWQo1bkpnUDHnrnkBObpHhQz1yHQl7XMy6x0+IOiCKiIlCVKn19+/mNcQh1SdMXddriQig09H
RkqlJhTxT+cWEqbt+tuu7/KKjuu5UAGUIISvvYtY6/ZeRly+BIJ8H3DBmZJlMzTUGROITeiN6cBg
jits/q6D1R6PNlm8cxOmXlzh2i9e3Y8qshX1bJ4aI1nTEhE+Ft2qnbyqlxD8BRj/olNvE+Vis+No
qnJMZuBjNWbZ4Y8UhlFouBGh0vYla3yteHPlCaUT5msDyzrprw71pxW1plktNnT5LiZVzKBXq8sN
FO7cZTo9FTQ9UalKEEYmkPWG/hVQhcvdrjsP66K5m0zJAwcGhlA8rV6ZtHfZN//c/NoH0DaDZGin
FNXm7mYcjR5CLs4zEYo86DgqlOhsL0aQ8P2PPof31wFtwyIWnKbRlV4X3vBLtHMWR9BsUpbJEUpp
ylusqZIJWwZxMNtD2eFzn+UDCeQdqnRAJs9tSKNl6tcvJPbsiibbSHPvhzyaMTeXUEgvv2amCtFN
zJ2qnLMAsZBjgbD279v2X7CLq7CW/3pRFBTU93xw9BuHtqJg0FJA0jeiUJSHWfX15fHr6GMRU9Na
O4kDauc784A6nA+PxnlXdPefUPWv70kaYBowIybgbIZjsofCsCCjLuEy9UR4O5W25fcgtgjMi9Ki
7ZifgojsHJaMDPwecfiV80PMFa/gEanPLS/tFQR1hfMX/ee7PC2QxnAyaXZoA56kPWwoDhr8fs+1
3ZjrKFbfSXpjbwVhsIzocaC5MFrMjs9BEav5MGWMcDGaDPACzAX1RznAmdPn+9qORqw6Z4HaQ78n
03WuS830cudFvEaDf54uiqN15WmSAW8zowhVCP6SubKZCid/fhEHw8cl+WURQjBW4yGPV/T5/S26
9eUyfmMIH1GMdYLphJS6WKU92FHsBtKqSHp0b9hPOHNM1gcED/AKfuaG+6HsGRD+cBf+XqtzH3rh
wzfbyGqYYFuXpTD//2n8wpdQYFQG+E+1vO3Qj8JSr6+PcY8CRJ8fSut2yobiwf4GwS31h7hFBtvt
g2S58CxGtjP6Faa/oLcF6D5MWSvQgk2JAOFoX6AYmxrXr3JkbKDyBJQFPAdyBc5tmL6j4OeviI9E
SdcumKct2mMXx2xzhmUtWZ+WdQjZNK1iGy0/eJY99P9WyFoNeUr6miOb1jSbhO3BU813T/nGxSHM
QE/cSWx8p01THDjx9nFZoKFsyim/6SvFiRse4wSVRWMLlnAXnls7TNZpX7dMt/2KoRlEkAwD4DG4
pX0lu5E9zweyplynlRoduPHMnV+wcMYbHi38UUc06Fpob7SeUcBfR6fwFRU2WylaD+OaQfCvpo9A
5ai/oXPE1vtxOuF3ddhP2mhgv/Sl8hnYuktI9msrbtI+TfELIbUoAPwBguVM4SAs4+n71saWOaLI
1oKUUP2nqUr2dnWWljGJ4J3Us5pj8FWPXWorQEp7aUSBWe/Bp2vJko+HZl6RRRrfZvrfSpxsKNBy
2rU7qm5szN+IofUtMnCDsxV6xXPLL7Te4MULM2JfSPkZ/uF6mzWviUl0v7d7NYgu8ukv1WsQQpKG
XlNLVsLaYlwZcMEMAF2c3QTpP81vKqWrnBLa72EeAZSMTyh9zcOWk9rR4NkXwNN2buRIqL9Xy/2X
i/vuIl9r7vU7/FKb/yWU72eR0bHLh+vYwj09xFpHhuICNcfqLDHqNUJ7RIZ8HBqjJcTSl3+kjPWF
wZdfDkBYoG9dO4mlGBt7oY9SsayT0mSPrPlv/Nq+wnEcaCad3KA2J9eH/fyZXvYC2xLcHS6cgZcI
bkBMr18iTtM6X/hmdXMVfQhZNVndrUip3bzLfU8PwynJ/MGZmIcIRDal3PkewUHIvQ1xw6gBEv9C
I4O7stqX+1BEx1/C+VxkhoLqjQnKiH0TbUE8T+Oj0/LKlOX2kFSylyJfBr9GCgIcNShVVBChFPvG
e8Ncv8cdzhNjsgax+C8cp5C6YsnTnfMdNEcsTYr05WEBii2BtC32OCo721/j6Uf0y80sKp80JOBK
ScPRuijl7Z12Z5lmu/qpKxC1GkihbtdAPhxZCvBums04HvzJTdFH4tPzUF89HDOGv3bbIRaYiacN
KJRKK9lQhEueFcncAN9stTSNA9O3xJxxeugP+nuK1HyEK8XGxM1rAJM4ugC8ax3+OLPm2TaLzzvv
8lwb+a2uIwvL1JYFRq1FqArl596rogEXeAdT5hEd+i+aiAQ2GJf5byWGXf5STX5MHAe2rQNi0rET
X58NOThK5BwBvk329SFRPG1/3yx0+aGeH/YF90SfFrRbqsUCkj4Aif39JlepBzwTQOoZ31jH/Uic
YRCCNAUGAlwNMj8Mk59KOMS2lZFmoZuDbWZVoEJuH8xGxvfUUy/Y3eyb/J4Pyn5cH+n6+Od1+li6
1Yoi0lD9yijFe8nvQn2+X912uJI0foRAjUlLQO+nSa54+3fWMtAup7QvrsMfHVPMCFvPsmOzH64w
FVXAO2WzOsDVjJ6zeiTOMq7bHFag3hFmpej2svMaBjh1nFoqOIJ7dS8WTlsY5vfE5UB29Lav/90S
3i5J7naBYrgo2vRPvuCM79qPQW439rHV+S9dOLRCDWS8paMtLmD7IUyS+6HEXdln+zU/BdOepNeR
7P+H/TfFiIFfcYLZOvFFJWta4rvV6k4h1r2f1zyEgFL7lFFc2GooNGZbIgvXLKX2yxwa2SWxXtuK
9DGJSKyagBXA62j7VKA9VE42/o3UNrjhQNCUFjNBq4WAEl+kCFiO7O7go+cF2K6cruFWDvgPc5Pe
7nRUrDYV8c6C7LGwtIAxP/RyKd7GLXf+DFEqa35/0lcA1J/zGGmOasOmtvQBC0K2BQxgWiG7PIKp
FHFP0VQuTS/TSGRj9xVMegKwqTo4PCPlf3EKHE2k0dGnpr4G64Wdmg2gXltRQvkgmMymPSOV/kyB
jYCGDbDocOUBIqSwGS7s46iJAe288AeSZAuzJ2L9NIZ2K1A4oWb5l9O+kpWUyN4sEzNAdclrvlZp
w2eHj1Haqn35x+mbA71tubrt3a95dRXAlaRLTC0MKbuh58hYDd+bBolEleV/JThjO/iYbLpp6t0Q
q/w22DevlsdsshbOtIqOHszuRvcA1WS5b3N4GWwKXLwo6i1hPSE1Ajx1OiKGdiwHCJMVtovY9PIt
DVQVcC5aIEWR2lxLH0//UQhiNlj8j06rAiFIWdvYnoY1O2ARbVlJ0HoVYMFeArNRfAkfTT8nBQ1s
O4O3iw4VlBjOkpniywLnfsHErxPLT5S4aFQdHBPAYeHA5yu804LNGDFYKbthHA/TqAZ7ZzGrh8LI
xjpGphq5YFJr2dbeNkXh4aQWOTGrmRZmSQZdFt270jSnaoYHlgDcu/O+4WiQYeyPtSc1ULjWiZsL
8pShtFadFjk4P3r1cNAvNnvFttI66fTXIZNj1jGPRP1xhht7CcQgkDoDh73TnFjNGIVh7y4PZbsj
miCJIkpqFJdvnywpDZof8cXFiudQaU09J0wlzDmnyNDzYykfLDlkE5H6npF7Hxeus5Ht3/t67kJQ
YyY7TPPbLkExei9buAgPwEW47H5wcCTFbSCXwcZ7u9+9UEG/vZ1rOaZea8VYfxv555a1Uyzf+E/Y
IX/3Nn6RK43Rrgb3n99KxHDR+DvCwoh7pB/FLVsBvsanfA/UrX6eNlxno7mT2ytzles35CaU539l
SA0V4Z4RUyvvnEaNeeSC006rxONJcVaybuJZHE1fjgjQQPa7TK1VxMtg4VQEFBK4A0QHHeYfJcN2
tu2hlPmU4r+RNElIYWmpw4n+BRp4ORnCgA1VpBW+IGe+NIrPBDo1U+I2nSppQnG0h9iZK8Zlfzr3
QVvXR10oq/84lcXlF5AJ24cdaXk/Ql1s/X+p4iHbFdnnqd8N2S5YwNcpUGNLgGsC+6BOhtCVcA1S
3u5kcMZ4k/cdVI2MU/X074kIOmbdOGUjFIdg5KUFKAsKnlBC1jqrF+sla3ls5/4eJN2CYbrKRMws
wyptYu1MtzI9VvNWHMvRCY0esCvTeO52JLsuoNsMygTaHavD5gnDCarhgo1ZPAGpXOxJIVWQo+PA
NMwIrRkZf9oMZVqT80T/D/1LUyyiro/DEqtf4KWhq2EFKUuQihmWy7Q77ME+6XLjAWxrPvr3Zu6A
e/IGJQ9nI5m2btblyy9vpOFmW9PaJBs2FLQDtXz22XYM96/wTytr1Kv/Y1r5qxdz5cdnc4OtG0YL
Zyo4qDZJqA4pxCHJt2XP510yd1gULZkHyNZpWQ/sUjsBfS44v5L4Vgp8IFabJ6FIZShNPol4HB+Q
CfwSd0bH6mIxF5CmjSS+EEAX7V0JxuHT5oyZT7vJx3SXs3bH1IF/czuhhKdAXAcCKI3dVGWRen8V
MH5eTeRl9TRCoVH/ZggRF5SIJmsbMxH2u9IH2DxkGXqrOphtu0wNXUqlrVtgmmKazBEgsSiv7XKA
+MMD4udNzJR8YYY7rSt2T8caMBczN9NEtvtGtPkDz998VNonh/Ar5aQunFY/2fyA7jfJW6NPTzsd
dVYv1AXEp3Xd+TGnIkeNYvdNWUdQa7/ojkeJXgp3Sq0svgKzVqADgXZY8OwqlhyVcSJno71Ws3cU
15eDQiNzID5JHHPISkk89vy6DeUlXh3WBc0ZZZtKYWsH5ySxWA73zL7Y6bpAT6nT04opfpQQtWDM
0oPIqyskBxJz+dagpy0j4Ih0cTaROF0lhPIKV/Tx7XmhsQzXJ09nx+BP9KGRhtkUmcgo/cw6gWW/
tkHpHEdK6q4k3vecia5QQruCr01QbMQwY0tYIteiLub8JIKvf6/hh9514tR1dEs+Fuakw8FnYgUY
jXC24msQs1enkD0JSNr5hvJNchexqcLFFTrD2u6snf+PQU9i1qAypPKZ99MXMMjuPvLbvnc8pBQC
y1sDonpf6OPkRzbSsp88Rh07A3iFNxsrZlnU+V3v87/5XNfJRI4GQTrE2DoLLehVVuiZQthqHuus
/hm1xp8Bd/AJ87goY8LjiJM8r9kkOZmhwBCiKSZSOZIa6P4+Q8yxcTkqsS0pbQXDwGed/u8WW9Nb
+tZTCII43h+zn/gBUpAIifp09vB6H+EaTnfc8pjjrzAIIzwu5+CW+qHmD6NOTVI9BZslWUjTdcFU
d/xxH2yyCVdaowxuGJFsjp7Fh/cNlhxzuj0rwkp81Niu1Qe0A7H4foQef4Ezz+hg0v4wK1D1c4UR
y7kKkbZXb5xgg56wOU2UTlOoxtD8C5WONQpprpHGcgJsLVhH49ZModWiaCOWaJPANv6WYQ3lpOSb
7bN3ggDRTJVsbVpZJX7Fxz7l7V64wY8ocIbdQpn3viMxgLZUA4FxdUfrx2FBD41T0QzmOEYmTX+I
naEnS/bDqZm7/A7xNC+jNYC/6eQAmnZrN7BpZInT1Nd1YSxwLssmAq39NaJGNiuKWZ3pF75/yQEu
iTQy6g7aIf2FLBLQ6A60jWphAJR92MDk/xXe5sazubfc8m3PEl3qstL3wiQGZ0dM8bIor+zzskKW
1ZO/SBiyrVpErMWrcxs+gwTrugGlyfFn1HUUXWHhU2pVTUwX/P5GW55Mu69vzA2tfjRDxgGmQonQ
8e7NIks1u5SocwNIv9qcNj623pH9+t7xTFSJQAnNuE5v+BPZ389bI2Xv1CxFZBIsf0tSTbcT5dvs
d478MVDVcVrnWj8ShX+AJAwiJIXFA6TWM9iZWbIcKl3SJL1HJkD4x2hzc8xaffiXDSu1p5v8DrEV
2xr/yVVNZ1wb0QPQ4Er0tpLILR5CSbGtggczTs5mNLW1KHrgAiZ1aqlGOvDQXWnBow6oV/mr53OS
Cu05gIhKtH2cn2eF1Jr98HNfdLA7Iol78/VHOTVaZ03D2nJkC3fWdhjcoq6IdKJ7Izr2YQGa/SXg
uy/Wn21ZdfwzO8b5OBJ2b4lBEFlKszdKUn23N7XOHuQ3iEkeqfpeGnEvG6IH8L1VwgPR+ea/zntp
OjDUGy05yxcdlHPewX9xRrqWIJ5WRHyH0mQlVfeD8px1/XHxC41obIjTmMLExcFgb00Pr4zRiEpX
1uujRnSms4JzjRuO41a5S2WrNkpvSyr+NTFX0AYHn3yk04Y3YXBXxBIxEALJcv4YSqT0xLLNNu78
hA6AzzpHg5dfLHzkcxOEg/q0dKSUc/EFiLhSXWhTGMrrq9lhdHVWSJpupc/aY2YujXzA55cIywJc
gOkkLphLnV8vS+B9oBOvconjU/f4+w69pLq0wQz14AhkOT4nDStfwgOc0ArXFEbDbZnTdVrWHkRy
RcZG2VivjoOrC3owtkKDdEYjlmJyFNWcth7C2WCJuWbU2oHtztMQlafmgm/3ki9Lv6MEoAMwQZlS
MNaEMaaLfh0kbqpXx4377s8MVL+3DaK6Yylz77rHVAh7rVnB1Fqx+aKYxr9LAPSSgtjmNx2r0syf
8hk6gJAGPHQ/3nnpZM3YO3rwXgeo7Rt0FuR5MrUWDQJQzom0D1FzADcLuaZd7d4LZ3b+vYRA0xJT
UVOjPS+g2RAlMZdRfDXHbvD41Wz0zb+pKgFqNT/+D4xxRTsaB/JIZTL9FhvYD6CUGg2T+7+MRZ11
/qzDsudvRuWFheo2yU407wk8MtjGnLEmsCJ9tEsgP9MSo/ghZ1qWnh/T5DNkR7pUv9OdjaVxS7Az
68hZ/CG+dOstszl3G4uPQI1dGTGURzHjpfk2qmp4yRVg4YWJO3aAbauNjmBvAmWS7hQJ3BRD4gIg
L547sQM7GEAijgAMMvRc57MmdpeMGk4eLZL05Y8jW6q6ZDbJ2sQa66HDKoUnQH+/7NAfoC0UszkD
3wgBtNptaXNBOM14P2xJpbVUURs2GYc8qqKHe9inHXeYYaErgKeVTHAmoHjhYfKktYQVkhpcXD1f
bcKRGLsVm34SZiCRJ5x/8FslZCuWWnxbIgBb2fuQPIpPYYSoyJNfN3GrU1Lmh/13t5f4CqERSdOu
XWOa1sDGtm7+K4kJ3Pf5nkEjLf7ayUNARhy3i3IFq2v2q7Z4NqP41xVwuNmQjoSFm4wz0Wo31Ugq
f+QCKF5pjIkk7kVxSO5N22OMBWR1E1NYAduhXEHYrg5hfsTDQic+QNunh0dlaX0p4YlbqQ+E00be
JLmG44pCQPAWNJgCyQXEJ70itW7XOrCnbcYflRN+QIUp1MM2ZlsewOiVdyL9uEUqfpBXKn9fySUU
yLVptJk7PwrxQ02i+4pQt24NXBre18960X+6uTydEBQWDk6Q6isoAb2Dmjj0xAB2XrmhDrkThhFv
dTNIKKrprlqe4Dqg9PSxq5vDDgy/VQgncLfkTmbOWdUe5xDrCNeV3Nu9BLCoRTXBS4nAcBJ/eOgy
jL71D6wXzad3MVZoINriLLARX9AwXU702j/1EKGZvAbDJkaxVV69AuGZWrNaZKjJmeZ7jFmNL1wP
yA+XfljWmLlJF0SFO8IrQFpp0d4/gsVg8aKQXTyiVR5PYtVkiendBcw6ckHP7xVmnjFIS5UiipNz
uAVRi/5iwNeUZswpNNKOm4zL9lfxS2uyRse+Pvsjda7OfVObo42+fMNcpe72SA4FlRCFMU+DMrAm
Nft5O4qOyOs3i7lvFtjl7cB8ghj4jIthgA9tAFimIEA+imTfk1hoioGqTRkAdCc1s+kM/6yNOw8V
7eaYpgP+usSo14IkVbGikBd8eVkn0BXxZYYNNHReqlD0TRREFyM/5xnG9JYbPJnhakpspsQwV345
1CnGBTOlcAJR19Bee2RevHlUrvPFUnsXUoZ+BhCTAF4FaGH31KjGRTDA6A96dS6Xb4sWraSDOYfV
DM48HckSDWvcaSHGcrM70J+XC+eqVmoUlALH80YMfshV9qV8pjjP5s29xZWZ315vbJ7A4CTZ1IOO
z7SJTLlPXvmgB4oDM3MpO5LMeU0z8T7PgTziSPeSVZ8vHE70euDoKiPmF3DZtMXA/Dq9ynRSw1+h
vWgv6kk4R6+PqbgW9jsKdEcq/euiEj+DrKqVgm0dX8JO1R3iKuISWEXJUTUPDmypmIHkyvYatD6s
htBkLyQ62owQitv1DdJE7ND4maoMLj8Sl1b60tbTePShNB9hhjk5DI9Fq9l2gPr6u3+5XQGcQm2Q
wu70sAiMlvddmqsTnexwXCL97YyS0EbhW9bcIXuDumHBv4ZgpUIyzECHASjkAHrQkRb9lGDGAUa7
KS6MoKqMFbKSpRk3dd+LGF4RsUsCVFcOzv3HC8HcwIgQRWK2zP2L4d7d6uIYniGeweg/wCP+/HlE
y3/GuOjLdHV1g86fob1PyXRPdlbbmDaaHa+39RoohzSwo5cI+Om4Nu7lzRwRArl9tGzo/ys20d6X
Iwv80XwmjylziUaxe8+5IJhqclwpCAuXvqEKHqtaS4lr2lt5hyl4mPsyxKktoWWHfB7anUS5JpIM
2cXtDqUb8QMoBRmpKxrbF1cTYeCD7H0K2XU2pYK2oQ0YynIRDJ1KXY7rlI9JDFqbYU91IBqdF0LA
gAfe6CuOatwW9tHIcurK8tNNL+Bz34w0/NoiF8PGih+y6poF0auAVKFRPu5D6CHP25ef/i8UDdXE
uf3vsbcwtDWa6/N8m168bID2WtfnlrnEmini20hPvle5T7+53lgP7NAfaASXfnzvBFihf6bzVY5N
y1gFjgZ3ge0OXOyucC2H5nQZTM+rzlz/TSU/q3cnUgAId0gt5TgYGcHFjO7O9tLUmGDkiI3EDdrt
Rrumkl/nkETqnGSZBDWBgVfSBBn5SS1QAtMpCy+g761ptWqD1pz1DkGqhkYXs3A4Et8AabDuLNJW
rf7rkfCnb+nlOiEHZzVN7YXa9sPHp4b10cB6uIsrGIeDDJSEfNzjoOG50DP4JOFu9+qMOuBoPG5Z
57ke7AVx7s1fiOSy/Q1Be2kLVD8cHxM/NUgOFnBUL2QZoxkw4ArSoXWldrzl33ztXTM33Poa8gLf
D4nADE1NPPzxqKBgKDuYZaIfDUhneBc8/K26iYIE6U2FaeOwrzdzAUhkyfNUh/We+yJbLMupFQIW
IpvGRM4oTzwJJq/DJqvrRR741l4WYYnPxE69AhRO3+X85C1DxZQePUHgGM/uLrjESrjhgOt0dGqR
aAsGmYwj7Fnnlx0+aHRiFUH4m11rOiOuU4VsrEjcwxx9t5CSiP/As0vn+T9/JL49bq0aE0180RX8
3t05q9hyZSDL0buoFN3l3soDEbcY+Tj2jMFtd3HSPeZDj0qTdCZU+5XYNGv21VK9JYpTiM6bdGZd
RX5GJ4ahdqvEY88RpurF/FvkaBs13zef3YHc9PYaaUFDqDCdUOHMtd1e+hiMCoMdbOVhZLq2BNBu
5I7OUiaL2otd5fHJQbETr57phgwp55y7XgzwQSI/6noONBmkI3w38Qq7xen4eHa7ZpMGeg/mU4RD
FfGS5rxinUJwe6o33VqNILRstrV6XFx8DF4JlyypTE4AuKKHUSI5h6tZNYBEqMPglvfVSdg/y84C
/XZ9QEcncIsupyBEgKXlAE/09+CxwtrJfyNuI4O25mqEV/ZcYXIgW/qtDv4+wBCmUmDs2PTYLc3m
PLB+tVy4+paYP9qv8TIREzUXWZV+dWNI2Ae7zIunTS61yLICs/Cl6UsnQDffWUH8PhGiqgNbh25G
pSOGDl7do6nO1iC8/uZuUE9mjmTAFA0Qt8cYzljCnWzt4VuosiqeiNDKgBCmI0HvyMos/4Kgkrpz
HTGJO9P68/lmG6SNljmyN44YSgTzPmZS9tI5hrJ4vqS2SBKbJdfX9vbd1T4OH+jDM/4Bx37r6lzO
3qIrkpzvC0Lxv4RE65Aq+tuDZTUMoefV7Y/A2Z0lO73QzzOwoW4eDun/w/A1MkwAql/H3zw0sPr0
/60zXo9+Ao4GUR+6hJqJSdqIkjyuh8JyzlLNIQNMnZi6KgdDqIzZfcUGo7yneZlvcRWhWGjnXHNd
0JOXeKYN/71DA1KD2PsRtum7o5VGQGvESEGQ12L8KwyPk4o3ik65yjNIwtbekPTF7ytnqFQxQ8wM
s9DK2M8W66jOCx+kOv+yvgpw+sLni69bZsc6faMXBBBI9wy/tUfWuoe1qnd06n1aYHYD/BRFfBqd
HeGQpCfiis2+42QUY+sggQ1+hgMzPQgp5RogZakFfP5PVQ2h56gZcraQvcrP9Tlmna8GNhTnZKir
Q/nja0qdZ7VIWXdBCdZsxq6XnNEYRCXUCJp4FipR6NF+D3P1LFWm0wSN6cVxs4ktTcIzzcGSWmc/
KGWvFI6ZAYEiubbAHycwoNiwmmSP2d4VTCpRKDkSpFf/eb49yE/rNH4o13HuGdBWSUyn4brakh0U
Ui50QIJW+POUx4RLaEEO/9vGQOuNpGLc8PtGCD3PPRxfRL7wgR5VeHbP6yRiGxMUjvdJQ31XfWOj
q4ufu9Wwjpp66osdzTzkuHvrwgcLmWkCqCp1chjjM3SpQv1FJ8BHnbJgJhuPGswsBANzQDME1uaG
DMeUNoIQeSLciouG0H2LPc6Oq4tJ+/GmP1A7v2x8SUJ2W1UNJnI87d1S2v4Mh3DOM1FaiuJmDeOS
XkyGiqCB4pAA0Ipf364+SjJGplj4mE9eyD+QqBpErtx91DfKxFB8hsa8gsZc9lx0p1gXpMVwdrB0
AiRZVPq+1dVC52S548ncYBEGQYBzh/losMqWRy3F24gqdUr5i4JJqSokRyMj2TB3wCx5b/3UeqVV
6tDWHwMQUzaNk50B32DklPi8fv5qr4oiyc+39gi6joTh4ppCL9w2auDjFssK5HjOnnXcDewonhii
PpHKUA2ykCefBKBixevGFmIvVTvSgR8hsyqOH7mKO/Lu+HTtRB5q5nxyBJ3xXxWeOfNtha9xjrw+
k6RnZSNNy/cSIRos+X/URFLpUrSfw1SS7QTA2nSaD2Ez6QHt40vWpzQn7nRsV5vsZAUBWbkf2OZn
07nSgGTelpsDZ3g5yNvMvNPr2EUHdyuTu+5mgkK85pFnj4iPIFzm97yjPbFQNU9vaNgUtLwmXmN7
OM0MIONJ+7j0i72ZT8sV8Dira1+CKU86PJSsfIB6b6wYLcLGOIsxvAqGwbVa824HT4MTyUtyOnCE
ip4pifnJqu22mjtYqJkvqm3DLwXRP4ByGWWYsyF5ewh0WSz/itR7wuendYJAH3HXjqEg9ttOjsGw
hI4qzaRH5KVuKftvEEr67eukw26uHl9u5VP2FzEzSjQMQkOaEsOyJvJ9nyLgWfvxU29WNnMqkbG4
A11omaUOEEHYc6T1FfoatZ2guJ/8Re1ariqTiDZ/+FDKwSKFnVze0bmQYzJT4FB3F8MTU040mhsW
z/tV1hAaP2DzMebPo8XF547RoNE+ShOBTJP3xIpEAQtVhOrXhkMWGKhxyPvGHttLUbRyp+dJbosC
rZQp80oU0qNzg73pS7iM9yEu03ApxcnP2Q6HiQSw1IhWot2iPzUw3tjVjHfwhxfWXthdKZ/BHzvj
QqEcLIKj9eejP8VazccFecVH+ROos3fUvjzEA6xfmrYqa0Pl4X5aD4kt8okGzWKRKofuuY7NTYlf
Eqh24JGm6swJWcnuDiSyDYtXFtIik1vPQJCbZBt/rgfqD6MSYrPg14YlKS/g/wuJZu5l8mSSNWqT
Obn1IF+pvaUaEFdTU+4YXu+9hdDEyZgZ48G7rYQsv4hp005OM+CBlpVmUtQVGAH93EwvrcGu7f0/
/Kl08Zix3rpoTHUVJ6+S6FZHXigYaFkLdL6BRT7JCInlMiGEfQqm+uSMKgGvIEURBx4wTDi1/5Hl
rv/Zq8bf2ecuvcT872chfT+jEF+G3TBU0hyfYrquasU988rtcxx1wayxSMOXoYndSUP8dz+8R6Ej
hIXG0OCvPw2e+dGQw11//ZwnDahg23mP3xtNYihLiGXKTNq0F2562G2CrveGki2Qlh+OxUkMwiPT
bKGV6kae4UHyIz1qW0PZ2cjlxoTCZ+XLwoSTjSPW7lB3SJV6WqHJPIHyxE2KmxWn0+F+PQMKcd1W
CJ9xO5/nUWyyHbLLyk72GOpGMqQl1N2wx2iYYbASDl4vjMjUK8feV56itD5xDO51Myubn7HeydfC
czDfUhTEJFO2C8Jm/ATZww1IebYNv0BsCoQn1WZRiirdxJgOPw/x8R8dY3+gIMNrIlm4n8grCItT
lePdF1p8mHozdRjpMPb/epa+UOsO7KYhRd54PgMwV6V5TdHYn0zN9Fb5BnATlaoAYFV5RKAIdKk6
VLiKngDTSyO/3nHkXqA+CtMFrdxEU9VbFz/4ZzaBVGnjvyy7Qpu2FdfTHsMB0hYyobeuuAlvo+hN
90iJMa3DSaV8WDQiCl4cLKSTAeYOUjFqT3EqfjhMOfGXhI//5wj1m6B/CpB41dRBvlTGV7LnoXPq
zQw6itLcUhyNNmD51xMa9NQQgBGXoLlPUpgRV9rswVJrogQLvxg47Qhrq4V692Ut5W9h1MKQ5ZmW
D+CYyOFrfYreeoJ8yDKZKC84fF88mnQX5aZYLxA+BM9pAufL672E6sF41kKzJ9oQ2AeIY/0oXoS0
XIIWKavbBF9IHXXfczDaGXBX2CnfYeKy3biMU0C7F8o7fTcxU2HqcK0Vsy2huPCUxtMM0Qi1lTOi
aesvxo/QeJsLhmxKYZDzSoJwP3PIRytXax3OZfPXpUzafRLZ/AppycDLdaV/qx4IzWz+iX7lHI59
EzOferq7grygXr5lMa1zwTqxJpWp8Sf/BdP+g0X5fckCnN/QxPV/qoxKtiN/3KK52cXG0N0RYNaU
qg==
`protect end_protected

