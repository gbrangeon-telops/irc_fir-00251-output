

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WH/1Hfau3yp/7ANrlzYJ6lp+xOi/gEnoXSHu7RquVCgxmSwM+u6NJ87pS5P1rM1REfM6bC/4VD/K
djLzpKr9YQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K9OQ7UQRJNNsqlJeKiLZja2cTpdn/7D08GuVLJ2Q7YwPyOa9sKS+3g/15LJ/yRa/zU+A98tod3ce
QlWEn4ue+HTvQflEH+MpavwOpNzd9uaRdRTecGrueadi0jZCWhKDECPBSOBftTcItmWjS+iuOrYA
UzNSV6gBgTESSUMmlbA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rfuGizF/z8gCeFD2+mr9MbjRWuTPDiFayAy9W9SH59KTv32ja3WRqyFVDNKefGFWmFgyXwscsdSc
S/STQk2WVtfaxUn47IIZV3HVYpgEROzZ8tdQyrDPMbi2HwmCfaz6YD5xdrfG9Tlx4ToidJJ8M9l4
XJdd32TWh7NYEzLxqVy6SlnR9JfF+0+Nf5C57mxaFcf8i5qJ+wGXhxEFyHFj5aPx81iijRBXdTZB
X7F/NtLKVCgLQvWL22LQZOJhyZVP7Cypy5OtaouwesfLnz7akydXxvJf1kqXrAdSNY4YWjxfZQKZ
dY2m3KiIO6F542kNq0ktevUOXRqWTgZJhPauRA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IUtntTnFOD14laEXhqBklNwiMVlWXctApP9259AAx8PFHjFAnJ8PvitVWk2w4ALBNs1tWO3QG+lc
7ANJMKcNRDw3DKgO31xMYxIed+W9fGmJO2Vhw+W2lfZUNPYCZDcGN5zCsW0hJkR6oPg9+0a7K7Sg
VTgdoWPi0vZlEf9gd0Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NobNPEAvOyayp1TtUWqLiTt1wnKf7VjSBi0esOl6kg2wXxaycO7UdL9j1KzK6yLaXpPqGWArWcdZ
OHZWjNgANQMvd87WyNjFR+DZMXSGqH3lTJ+rUOlsySu0gV6nE+CIBmIaadzXmtjlUXyV/oEoRCZr
rq22ZdRXEi/z57ExJp2QenIf48qX0mmYi5gFLdknqEc/38ewzEWm4uHsakTPzO6DKZ89VmneHDI0
7Rw0KBtgnhcNeggKkHBNrVAExbuEzB7b9xOHs8SicGFL9UTrJpF8NFV5zuKj6z6MHtvPDvJ2GC1W
BJO4/x680qEH+0G3sdhClIkA5Ln0j075tcfv5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73072)
`protect data_block
bP8tThTzcSaq5UPdwrv3i6hcfedmATTr4C5727PzN+MZCp3v01OZ4AbUfIg8RGlsEF2zxHCVMruZ
KuSXp00OE6bUCV/eiWsZmf3jtk3/+akG4vlyScT9rq27c+jB9muR42OGmUP3LDhvQUdqibiHBw8u
orEsikEweMDaywlg0yUb6vJ/vfqgpUnMHzXeNZUk58JHc296sAChegH5Tfg8fFQeqiV9HrVArFrn
zNrp93RF0vWOTcSvtqqXfJix+rWYpPzqgXN0YhMKcjREtKhtjJpCKiJcLXCkodoSmnsZmmlnt6N8
KHLWY5tVZy8gLanCxkwWYYcUIWgsk4rCbFpFFHopWUeqiakZz8MMfPZdDR10h9H4iRhvhJb+J/xc
Lk7sSIi/TMqf41O/b4A/CjeBQdCNi+0WBtCPBvCNQ/Ke9j8fygM89dmXsLvyxtIFl3IWVBYEA3rE
+7H99PFd4gi7FszG6GkSgBQMkTS9TG6kMHEEO+xR6b3lT4Zi7SP+4Zpzg+x4J+hnXgrvDFapuYfO
zeZ4GY7yrCZ7vn+nHpx7evC2vIZdq6BAoPYUsndpKnmK2ZJuA0x1mTShTLE9GjRH/iT4YpDUAUrv
zF9aajUyiBzwski5NYpwwDr8r1NHm92jwuBW+Ab5uWzkrxg7C0c1cZ/Pi/cpnx7lUCq06zp8WfpZ
AjmQsyZFuSlFvT2bKjDrYCVgQ//k5jfMgh4LouV/72+peOz0iO2ThKpB6exeWTN+tWvwlRZcuo3A
cbTa3c4mm0LXf1hd/LdacMGZQVYjE2cEUy9HGXW53Arj1kFy2V3xZ7o+Bo2m7vW2F4UElx5kUZTo
x7JS+ubmbUstgOPqVt/3xoDoo0nGI2Z02OJfX/UDbOR2iPg3KMU2L5h5L0l/o5oSU+r8uFZJ4oUX
jO4E96bzjRd0cModeA3EnpcO6F++hPsbr1QxxsFWth2S1HXr2hd28vlv5Z1oyimRMfyGh+c/SNAh
hwWvZudvVz4+t3wKLSeqXzLzbUIkFEoqTrkGgY70xMUH29yspWg/LG2qXGXd71SEJWiAqL4NKdol
GcSw3AUGvMbwViLkCPiz3salbyT8r2KsPyMPaBjh4Al/vhbfDpPQbtv+byE4LK9xlxlxau4xnW0r
duhrCJOsRNdE/tXzXFNyFDIN3wtC5YV9tUy8qVbXL/LhqDU6rbJz9IoiQVGPpUsCll7Sm7Xm1KQl
JSLs99pNLelvPyQGeesJm/x5da99+0uHCgakxvTtDRi7gK3J1vJMf+yZxYCVeDhqlR0FG6qdr43x
fufRwis2ZBUfPW8yUnVGKOABY9JBO6TmRIQSWLeh9UQ3Vxb+ghmKLWIPGlJw0Ox6+5U/Zheaxuyg
pY069HFRfqPTikGx/Wkb27TIR+nOP52sgp6F6zUkqEDytjGsSiFyxjxtErT/VzqKiVMUnBBjJr/H
v3l7VXrEZUBj4b4pIHXyxwIK5d1d7BcSSHXQkdD+itlQ0MLyuySgeycncVzc6t0lim2au0aUPEqg
OmihlsskXUwYeWzORbic2RZF4Ow8prM+fH3lpaZ5M1SbfDa00TI3zhQG75JKqyLP0q9c2Ph+vERI
YWNyiAqC/cIc3F2duOMPzYYXgzCqopD49/egyeBImYBPRlD3aeNX6jIsKlgQyrYOOAxXS7C37xBt
p6ECh/ghmJ5JdBQs1N6XHXPtJvwnkiznXo/hd8YRuqrBdhcbada8LcJgg/itiqz7AmWGZoo6w2EL
0icgqMcEffsM7jMSrUC2IPuwAFI8GdLgQsqvOINSx7xGMjuxoljKUTgD74yOMx48IkWpAvOii8Cz
+/o5+qlmwhDFdjAzqyX9vXosYkN+AdNdQL8SRC+0gHTxeYqi+NcBvR1vhlEF/Asq+MiuOISkdoKV
F96qDCrWAQQhndzN0VdluD53q99NVSAAG8jpuQE3mCOSpslTwC1z17IqzmQKCPuZ6PJEkNhXBEfa
4SPrtT9QJSVRnbufBU7NDajjSI1kYp3vopNcowKIjrrdYbskzuiy+danrlzzQHW3QVfejp7FxO0U
OWB10k0Xr7UnRr7GlwqwTKSgBPZO896galKJGhsQsToRny9RsDSq7C+hSxZ/VevDXJ1gupSm8Ek8
nQsMiFxzHk1BrRSMzsVZ+EpbU5FqYejYDOUTshV4UUf+e0V1O0vSyPy2aO7uifO6JrDtHPz4rU+R
tOah3qXNl0GVMsbOiIELZTGpCJ3LuWcVhZNsAYyrBOhEpS/pT/GbvO6WvYx1Dxeyx1298xf8QaqK
t1ItbB9Jop6hgMasf+b7swVlJQ106PYDp5nvUtjvj/RaU6BAbZzCm6f4UkmvgDFfrZhkWSmIeY/h
7S8heqs3SboXbFGYBPaNiXXSAF7sC8YvOMraBuvrkJI52iuaD2ri432lSuTofeIWPr09oGtdSruU
hUZwd6KDjOpkCy/1oekCBWYNJPulLEGGsh47t+K/VbUoQXbXZ4oQXOqx4RQ3W26jdjO7cgPbWJGz
V0OyEKnD66dRLe5Tyq49lyQqFe9+5awujw52sYAQrVGv3zfg6xUPk/ysBm4jQeg1Rsg3TipI2dhM
SR7uAez2cfQpwdTSdj6fgMRddwzrV+YVeP7bVjHJNH6aGs3UBEHaWocLEek55UAX9yM0xkET79Ln
0p/7G+v7IIIBktkB2w9VqADJbaA27TzIcMxyg3rQitsoAUw8aV5WUakllHdHKbXwErnpzP+M9kr+
mTMN66w9QkFsryVsKR/5JFFUC1JaTCLgLtXrMNKabbD6jtLeFkHmrAul8wJwoxMgEmqfXCpIpES1
2QbGGTv8Elw6DgvH+QfUC8pMa3TQ3lAmwuf8wOOwlMZjFqXfOknAe7jB2pxwYg+BNo07FgzLdO5P
ZHYkf9COcY9qOW7KivYtv3hxaEfTYWPTE7kAmx2zjD9Fc3wQZp7deM/MEObKWm9zROKjS6/0UCAD
dL3YdjvSHQ4mOORF1oTsUiDGURpgkxAxjEcu2Kb7TbFxpebQpoaL7m+IlGaV0V+EcUbYOBVP7u0d
wKZjteWd6RAlJxEpc2GRpFbGaVYJyz9TL030K0rXo3F5HpZlM4lSMpzdrsu2Ht9x4s/QzscII3jO
Pl5qK3ca2+G/0zGZbeNEL3MOWT8Mu8kLIezlh4IoprGuFkKLh7ByEU6MiiuM8r05355NhBoTRcv7
ZzhTyt7/g+wa6vkYWuSfjd1R+hTuP90waTPspRnESHGW5EczS/4cY4FvtE5fFgeJnTrQ0lYhhnVI
7JyjZjlK8oIsfPZE9rKspRm0xer6rXpqRX89b88fOZ0CHXHEt9TkDyoBrbYJFTEKxn5frdSfnRIG
0CrBGpWCQOOaQiDllBvxGt6L0g0Vby5stiAFm75AyouifwufP0SV/CJU68YbuQlhYbRYuinZH2K9
M4VoVXuY5L9ZJuwDRSzs7w/4lxFwJWOfrUTPs2oSojRFPjV0xoNtpDQ87+wKcDoUtritr3cEt+U+
1oEhaZS8BdDH6FiXmOv3DEIqfxwlVV+yrQxfiDMzZYZkGC+mvEmpqLof7Wp+p1Wl/3Q2lninaHjc
gThr04ZrFANvZpF5DAlUYz3AHN1QnmYHvXEt2nruRwcmYj9fC/d5rac2hG0ZyvueXmxR255mwNlz
uWy8HYRd02rh1qLrwZBq/vv5CIMj0k9apel0nfPopJfgH4UBccinkG7Jd8PVeV3RgL3M/TOFPsBY
W+z+hyy7dP6LnH1TpO+rUT9Z2QiDnXjRIpTiDePxoFp1uS4/zKpfqGL+sqvxeZ60a818oHPWOo1j
hBZk+2TB0UzjQcwlqiBlE3CX5BY9APAVeWeuDrq5u+J2pwbwE53pJ/YlvJjeUOw5aGwH7yz6tLu9
d0wqHTrTxdy9ntb6IcMVPK7RcsnMBJE5ITsYL/7n4i5ngsZ7/cEkhzfG9vpJMZrqw+S2EEslxdRo
dWzNuwbgq67LCozuiMUisMijWwiM+8RIFSn88mhQ3mEcg18YskxH08wzcPZTI1XvbrjgkZoMu1R3
WjF+1Ux4c+OPZ60g4SaWPZInFGbTkcRB1LUeS6MhbYWSSQJ+8HzFfW/Vc45MbSr3xXnYHr+U6pms
+hJ6EH/sc8DqOxTvaWt6aOFxxJFKXKFXIA26K5aQtTXEx+6RN+KTKcuFRhZZvXrRqTgM64HCTEY6
JzTbYwdwwhoskLmkXrsfo/YiPytdIWWHMiOIpF/Snm/fA4PwamVhMNU8AgUVeN0mxs2bqJXjXVzV
rehG4dYejoQEABYwZn7WjH2REEsS9C3y6523jjDPz4otx+/9Lz4j5TRed08p4ci04U5Q6AT+4Z+7
WMdD47EZ9aztrXq306JnkeZfDqe9hCe7u6DJYzXxaY8x12Bu5FOCcS4WFR7pruLW4EdvBan5Fcqt
cTBug+FGVUvsPnUqO8LEfJP+Z8IuRyqGf4YQOJLhkD1udM+LyyrO1OQjxkyFb+w92ZDY6WPXbhFx
d/PLAFDkb6pJVzq8KHtcdWjfwvuADWX8Xqm5bOBxC5m9SsCz84tDscBiN4N9+zNENhaAHTPITIcV
Lq0FYv2JQv+IAjXld9Ieap5mNE81DW4qCXYE9vdlbWL9T4Tj+VMUvxr7kb3lXRFgnMw+3o/zQgrQ
sT0AT8S3QcE0bxWg3TMdMfN7z4JjHR9I+kScTeu+esoIJbAT7OOwxJqjZ+il/PCmaSBlBjd2bVlw
lAOy6P5bM06Ny4EQneH4Wt5eqem8au1jNss/gWZ9JeIVr3fsrCi9NGLwHloOgPzveEWaPgjL3C3Y
4oOrz3uPVe74tt7vD+PNd/oXjhSjuBXy6iFjfV+ANqUeSEgDuD1i4n3dA6sRcjJHCFpEhfVKJ4eX
22GlSGOjW+YACi/brD3IC8HSRfm9B/XgMH96l/oydT7R/CfarHMN0XKmKcDjdkGsq8MH3BsA156U
6PZ/NRd3I9OcyktEZn3FDMIc35I6rvhTyaCJiQJtvKPPSXIzeiZr1cyZyBT7s2HuZcx+5N1brJkA
OkdCNyhbPWC18T7KolG5oPvUefCMsKc34s2jHJipSHHeex4xnRq5zva+KnUhk6lXx9s3swAv+SEt
d4uAv+eLuhP9Evf/THPHTPlOdBdC8CtaG/kUUXpd9ayIGey9cJLhJrIV9snVW8n1DmlRKbvazYbW
bU6Y7cDJAsiTwIpo0Xfm+hh7faFBpQxI2ecuXkkDXHOEwcWElY5Oa1m9MqEKHmErM+wSYaFjN/1D
2H8KwyupUK3rZ56FROi8/5mQyXPLQR7jjy0wahGW7E8xuSZXtjUkjUNAiIdA2QDgskONk8YwQNza
IQUxaxz3gF6Dk9SIwFV4Ewhwe6HiKrf9KKYrccK2A0BGD4n1wfTA/vZpBimOKy56cLqf1wEYGZAl
83xGYDSHIdZz58NlMzHMzCNlmqOlL4R9Q2DYGSOBDrXLQdK0tiLXBlPNHS12Pg2YpKABxF87V+EU
Lfk0HwYnS091znoJtlfp6sKj3DV4TvgcSy8OkicVdK6P6kifpv6/RUuPBxNlHfaajMD8KJEayKYz
YjgmrlgwFoj3iWVHxFTDQJbMwHCIGnbFwqEAPPk/PAJLDCUi9yz+kdmYY1mNZNJWfpjJ1E2vXnP7
oNzXCzSfctcdqKTrgr7ZHEKmsdOxsiXQ3MMYHbl5Z2aC/425d/0KwMNjS6Sg8xTtAZEQJhI/bmjg
hvgRviH/PZ1h894A9/S9rgrh0akJ+VIxxLhiBd7ss5UebQX0qEEc1F0VR46w43BTwva64PEjb9ti
uh8c5LFdLtd8GVM/F8sbMqHyM3Eci/1WghxDg1PKNxOa6gcz30RJY3UHVkLlh4vOr1U9R46BQvS1
rczy7NbX+G95qTPQmN5i9TTt+/iexd787VOz3sigaZc0//wEGNf6F458gF2Hewddtz2zvGbqNjBb
SxC4T7DNiJOkIJDEUPQNLOagFmG7aXoFKwDkM2VQmJwyEdGvhpJmsZGMwq1dny5ToPIgM7bAAD8o
2q6+s1mJrpIqBBrzfi3/KpibZwgzxgFRDNjlB+nsczGRElfgwvbwZUrdTwSREykxf2Idku1yXCBP
DQGINgLcQ4snCduSiT9RHJBIAmEGoBlWdmRAQD2rpCygdnBwL2HZx/W1iwlMdT0KXaaLK26th/wQ
ehip/qaeZNPbhQj7Agp+cUEbF/zmiOAQiOe11Lp/ZlQcxVX+paefrwW99r4bRu8ukzCErP7V8pvc
is+QlF0218L9ogr2GtXj6Lznfl0cT2KwEKgul2dkmcryL4TNRTu/I+8LOPgUbjASL6xMl19bWpcs
LglBpRnpxOoRpwnQFe3ZBRd/oCBr+dubEmRSZLFMKqTUGUWkGYtUm0sQP/EZIXkV5D8yS/y4lZDV
m7cWiJeI/vH1QntYHOOuBnddsYx2BhWlN+sngc43Ahy0XIhVLC2yIPb75doYfy+etBBq5jKc/Jbc
Hzd8RHbgs4Tj0Os+y2XipirMdywXLcj/IPge7ExFKkHi5Ghe8GIkzlBDiXe0wIopu7NQRGtq5uZV
tAYPoziBUzEXaLpIak79+4wPaiZEyBBYCqd3i2Gjg2KeAS2jn3t/FDRi4qPeslgyaLINColdpz5E
SVpV0+/vcSSXNEEPDpdA7+/jhKd74QL+0+XGwUgJWi6ttzpooiKGfLFznd1sVs9dA1P4xrOBxKxo
jH8B1nzZQwvq1ceFKNhJE91YA2N8whDc1V+4aC1Gy6bRC1ohWjKwrmfNvfo/weF+62jJG3DtAOuM
1zaV+cuzBA0QZEnPu/Zmwocpx7A4nE5hY82GNsV97HHUDemO5KhvYbJTRcTrX1h8616aI+Md88DP
Om/D7gSZvZbUO9Qlq4qIl6PSH3VHnA0G2dFrfg90odn94NFCvdFv1CfkhSw0VgSP9ZaNLQqsg/ur
6biO+Whb1INYJKZuNSRo4tWa9OHo6BTlpAvRCyivZ8S+75ck/Z+yapIJzRd8twK5nqMHV9FArup0
kbFs6lAlaudwN+ZcbM4rAijc3tiHw1jLnYuxJmk0iMZU4yl/XtK9ezHC0VJHPGCJ/tEG8MN83Wc+
lNdu1xrXPEHZKIVm1rjR7i/gQYIswWegyvG/wZSTOUlWHomiGjQYTEZWCE3dMnCPQxC6Q1TG4duw
4qSVqz63jCnccBmoL+sVo9otKtdc4qA1ZtYT/99o3qgOfNfPPuvFdwjzIfrg+3Xcq6iR3Tj40eft
Qb41NK+sDD65DGIvAKyr/4QB6FdihUXNAbJirNAAeIaGGOAkINoRYz5VQFJbK+9o2GKqtI7fUc/g
czgiqEeBvQsK6WDomRhaamcIOF2cGEky/6Nuo3PIyTUt5riu5IP7j4YxjS7nba9ZjqxkPV+X3Cys
aEBlPey886oJhPeWjIT1re4/edKY2U9/UXeV9u9PlRvO8A0Aac6CPfN3AF8UUl80JXzQ2T3Uqy0D
4EvsXKCYFbAFmPd+XNu1+W5f07YL+WnR2XaM3N+mGsOga6Da9ud6weqMiYKVLiXVLltQ5fcLzCYn
YdZzDK7/E+ANMZDkrU485mnhdVWaqW/wVSn+huoEdDM7vEPICV/KIw92RVpbGOttkbHC/n3SHKwW
lZMr/3/ducKDGq0dzueGHc32lqtHLV1fHitYmpGMRT8BuyNKHmxC/y/HcCu2Fx0+T+V1TpwE57hN
lt+JvQVr3yWvDbHSzkkxYKk8YotwMgCUvTtCBYLj5OTiAeoptXlbPMOZQBCl/WT5cKX7YgRNKmPQ
9IgxwWidINhzQ9MIQzuyW2r2gpQJNMeyf7MgSkzP9jasOKkEGP/HLAJXCf2D95FRXUm82hny+euM
k9ys9y//vlrFnsNPoDBhJThrxVi70ivHpRHG82l8ivScsmOvwEu7rUwcPC7hF4CcGKnGGRMNyXOt
YAM4aGMhOFmYTx/8I2FHewnby7kMlrq848KrgOhNy1uaM5Ssnqd3ucH774USbK2dGOfPS/6sIwo6
71KuVZlxW0acQGlErabtS8jmxV+yhUfLfsy+Mtq9K3Wp7NaSdXMwzEDD5WEXweerqKttk3EmY7G1
gVkPdZ6Ycv6QVNh8mSJ+CFnwGAkGj80dcuVAeMqHuTsnz0DXpJvgaA9Bpdxal0HG7pCXh6oIKHTh
TI8HHD/FpdtFJ16+SS5fepGCEuhH4fkMe+/PgN0IimZBQJ7Qiwe312hGFAIJ9fJJs6rXvigBkr0r
njt62dN0ncoXUR1vI29UkQtj3LEie2Bxv03kdRDf/BZJEtWYW+9GCJCbEQMEcyiFXUuqLZn9EVvT
6yObepyncu4uSiumhq96vbTe3fI7uLg81gBLHE8YYLPMIjEr7Dl4lvuEEmljZ+mAYy919W6j0ho8
Ck5u739VloDj7WgWrQwvdmLqxusoOgsysXZns8vwuaj7OKqwhDqPI5+HRRb5RgTqtmyJGO6qAlP/
Ge/fN3Xo7mFDaGMR/cgl5TgCDD9Xda33XGFyioilM29K97/ksUVShr+XUoF+If5l3cWs8Epdd7ig
Rrvrz7Rp3EWih7feCz2UJiFlEIKAHf2MaD8MVg6ccnF2p1i9B39sASX632utNiBO8ek2nXYi2uni
PwfZTiom0JPMvSYUZJzSNYLB7Bes4b4U/l1USLxAV7DlyocD1B5M8xvkPlwwUo1dZniYrW8rMf6S
E3oWJcnoWhFobbE6zlxm7qPC2vFgDzoMqB1XFWKvMoEYHNZbE/KdEDX2ouXvxNUL+CEQ3452XSS6
MNdStCuVswvRVqqfGFe+4kUdYcOWv8xGIVQbjl8qHA3JNzB71u+ned0aFVVbRnkEWWMaO2KAo3kF
oykDokjlGdPqZRRi1+WaO6+/MabbtBmP5kS5XzJUgH9fIZqqw/z1lmogjtyqKaQqa4O+YIJFPimC
SUNWO1vCdJDLlx4sB8EPu1hQGEbk7QaXnVtG3TtOmzocO6TE7cv+2/ZPwlc2xjM3JgvRjKXs4dcH
hsVilqYNSSuvgFUJEQOO6VMfPVw6jozvg2n2aBqGI+vFemQZxCtVG1XdUO4DGs1z/+PdfV11StJ9
YQoY0c913iRJK/jd68d29pbPC98V0Quzpn2c0Q4jHWbc/I0Pjw0uioyhsAnyuXhCOTJg02QRmX1D
iVnG9uacSD9YYKHCNiwBSlEh7Qr2U/BK8LvAImcyDW/HnxLT1aYDbzHJrrRbxlcDvD/HOKrCXvjG
qFJDXLO9JGcOYE+4Ys4Gs/aKjCeKREOua8yOoe+s6H0NNqPCDZ2bqZl9E0F5vimd5VnC9625dmk3
jqkFjow8igN4ifGN/RjDxKOiip7uY8yko6oDM42kmZFL3bJr6wGLBf414UDoMaUCPfuMQquy3+qr
0r1yMKfSdvWxzje+djUIgPaNw3ggWAwDJirBwZB8Loq4r4ROMKTo0J3gHdQlnhiTVP1qy1x3IyZI
QzfurFf2UBISRo8htuqClkvcJNVL4RJZqfdq5qpThQoNKx9P5Pm4n68DJbJyFj8W1iwekYNlfDKQ
C+wkoTE7V/3ZhtUMBXTy4/Qmrivsd19xo3O+UxFtP03k1elUxzMzX/3G3sGgYF1fr2zEtCXVJQlM
mSGU7JrgAnAjk3m3WhZiqeBlUxgiqZ6pfi3uymTtIGo4OaYhsye/grlgqYRfQem3B5+7imWmIuVF
nO+HCeAPABFy8jiBMEnQi5Io3gAZxiFMACJdibxHSjfeyb0hn26HL7z+g+jL/g9r/DfzQCDHi5Ku
fk4QTdSoMtWSgP3iB31lg+BttzkXukvfQI4h6iqjny2X0XHzja/cfg3HXqGEz4DuIUGuzzsJG8zc
g9bqV+QDDEKqwpygW88sV5DEX4tYlbH3tiAlBIg87zA6hnjJ0pt9ensU1TIIh9mwKyPzN64pumVV
OtSubaR0KW0/BWjnHYuBoB3PQN9VZrpIu5NMYFTpho5qmsuStyBXHD60p2mysfvuqUSFZS6B5w2g
sWhyE35IH88XbH0XjRYmjL8jtpnS97x4QyBEkNr8/e27PemjDEJG977nItgS2EHfdZ468PEROnfT
gFnaJwjrZzHJkiwqNJabX19YrYfWxEkF6rTzcytIRcqVEegHxQ93oO81D8Y+cYWREIUs73TmurLT
7M2oO31x0Ygf4gk+1nZyVsxJ6CDQUH93CWa9RldBofqjHah1z2dgGwD7OnCg6oXYkAp3IGBr5g4A
EgltcgASSWeoYv6LdjY4xDvmOo1kBF8NyoXwCV5WGfcJkotFfgq3U9ky6bFM7Fxp72rmNpz9kXmU
JtM06au/OS098hlzKTdKlyGO8csBXGUK9T03w4ByMw2hUF7UoQhOwYu10DMy7KZ7UzQlSbKqPwBZ
sPeRHHQ5ehcCpI1ymmahA8J0CBNoiSRKan4SnYHYxDlvKtw4En63iz281yHFaPGFAJOQAZowOwDD
/42Ag993ilNCiDxgYcY6/tXwcbpk3B2aEl6nTijsoXds2U5U1WSKi9UHf742eci+h7KREDnvvwty
6jiQnUqx1nhwrZ7/1fCDm5ykW9v0e1BkD5JlUzDmb+VDqR8SDJJmA/jKBDienO1YCf2yU8nc1v4D
PQxJJXa6q7SY+xyZA8qn0bVaBeS76JspVXeRS7n4veOnTNdMCfTlmxCUtsvK8Sv1d3Obw4jaiLv8
i00v269H3s5qxM2bI1EpY/RsW7EX/LpqDs0AVof5w9EbryvkPLQk+UOlCZZjBQiAxBza76pe07zz
3i+DOoT/w7Yx4iKTIjBhpx1H1YNR8q1rZC/N+D7Qy1XEiqRUDEbGICoCwk/16bg5snnGoAyMbmXX
pobpVgdS84MAIaCxTSF7gPK2QCkuepZ+XmadmnZyjBaCYuvBWz+4IaGpTHO3v+UFiGbNaf6faGPE
HS0Erbl8ZihWJWwamKEzOCTD0M7Jn8p+UiYtsk6LJzP7uQUdlLcJmaev29N5o5eS2EfOMbmTSeuK
e6NLbYTeoh+dIsZfmYFCFMMlft5dct3KyaQhRj5BIe6TuM6JOHfCENUsKI8iVLXz3iTpy7ejvAR4
m+TZ4scI3GZ7E6G/DMFoe6hB/XRpF+XYIC13Eeg7dVNEzgMmupfBF0CUZY6834PmRiwKz+9Z+1CK
V9yFTFqSvgLpKKzHPWnGyJoz8zTW4tqsCY+56fdGX6VHhIxCwXgp/8mnx+iKWZsFRAUEx6km/s4N
dPGZImGB3Co8DLEJ1KBvYeQGLQGFpiBXIqurs21Mci5k0IPH3kY5HbJN4VSzZbQj27Yx+ocgQpCQ
NJ6MujeysuZhhC9BDYyXaFlFsuGY+30f7pqsHJLNSBopXIg9NDwW+FHh+YmEF1pXFfTsK4+6xgc3
oZ7UrX+MaFxb+UVScmIztRPSnSfXNzSxALo0g0+Xk/eSM6bAsFrQFZHlnYQWOW2aOrhVtZDqt+ta
ozzYDpvnsnplBTdCQCK+PscZHlnZ2HzGaAaR6r9SYTrecPZG5EfFJkvbAFSygvJKRpah4MEbC44q
GN+NPvgfS+elevPYW8VZ7R9z2UlRbImDI39hqZohbdYjYhNU3e024CqtfIcq8zu3/TdjRaRXLPSd
L7sHRtjF+u8IDvcgHEvROJk+jS99oBoIeaL9Nda8NzpaQrRzzyNaUF5fDb1lTCgrdzuJCt/4UC8O
zlX5WbV0mZTfl4Z1rdE+vdoJgjlCn0HoI4ihZWDLLlT0fHq+Yfm2AM9mV8ohJesVtTnVIeZbBAmG
qqN1W/Y7CLz+5xGIyKlON3GZl1XhYc39Uz7Dw44hrJOwT23vIrNrznr2KQwyDeIvi4t/tqBTmXqj
3Ud+eFAYdNdCCnlI9Qo6xz+gQDcqHpcvJ4CFHBOBZPQaCMCY3eyNO0tsGXa0oIVvKpuAnoyKGWwn
LNm6WjJvVqKkYmAMvMvsGUGZu3u44+D6feQ9DzCG2NawNtQ5QDO8CMzvDNMocAcGZEhoJtKwqtfU
T8Fex30SX7xeW0JoV220czr2D+ot/C6rBvFhzTsxpld0CGyFm2sxr8v7NThPF0VQK7RpO02IsJMY
obFSbM+ljtgdCn4Pu77Qth/6rAs+8Ivh3G31NKKzP4MH6PqqjK08p4MOs0j3cCPYceguO9StMa71
oAVZUb6cmfxCb/SUiaLwBIlwsRqkG5de12C8kDNnAmiB5rnKSveuu2zZ0cWefHnr6dFTe7H7NlHp
BKTmgl+TKo5A0ZmolW6jVvhugO+SL/ech8ASyX7dW6s99IDOzQDukZtTR39IAcNJF0r9wsZOR9Ik
sjR0SmO8V5y/t/FpA8+8y45tByqOQvAgc4xBqZZ6smBvPGwGZCUUbMnnT7oELrw3WYuGrY4lDgBV
na2+eiIgeRztkg+iN33PqQEDvn2cBWMExfxm+mbCX4R5M1FWnKS02UBVOiADp+YmcnTJTD4jrT0j
FeYdlb3dnhi6foh53qGIGJpOh33dhks2NSdiLyThzwmA5SgI1FrjoBA1rpuQXqQss0f8nVsWpdIz
PST8eNfGRvJlNHM1qEz6aOYGgZALQtc3YqAImmL0fRhnOi9lOQ662xkdyPO2h94EHo7qtEYKafwI
Tr/BaH1W9EX00LRr+67PMsoQ4szn89l/7tHqyAhBm7+X3I3r1p0I4dsdxDflaWLpuaFuNf7kcXfN
5FDtWoaNjad8PQpbiXqNG5XoDtdjqqSuNGvqdz5XnE7Bl9vp56c75cV31M2wvVNNYkv+L5bbFE2F
bmVeoIVYSn9e+UCVdY4cijCJvWgvCGLYGOgjmg1PyHYVs2H6Oy2scrQBE6g/zt9rtelZrhuEzcBG
n2ZHs7JV5BXXIhg6DeY6y/Jlm5qNwxrId6MV+J4EtyMiJhaoYeMagIJ8QYX3B3qzoR+zFZnDzzeh
Uh0gp+VNuo3HDzJZd3GvZDyS1swmuVr2M2zQedaJQqoCYCCPzt+XiJum7xoO0Ob2/kO9uyLsKDD6
Y96jaW05W5AWQVO8KcbGUnPAup25lk6v//sngAq2CRMEq7kSOTupSy1niZUOqYx4hhQKuhFnrgJR
WQ4BhxNcL/DCoAXVoSn2Hnh+mp10827fu/AW9pzSc5m3oiGy2tEAn5kjGvZBQIkPqQdsPysO1q5S
FXixtuzTz0aiNU2B89jqKfzj27ZigJNWIt9P2v+GS//XIr7KU33V7iGiGZyzShFLlCzLnmfwtJWy
rpjIHp+LLuWtiqRLr/pKJqmnEF5S5J+QIQZCy+vyCX6QNL687nJ+mmCoUtHbmZ7r7ylFsE5FbmbG
8gUMmron7F6ri3yiXjXHGsvEpYFwdge2RHSSnCTHEebSeti9OyoS/Vzny7TUP4kpDjdptDkhB2ZQ
Io86FVjOT97FkImNT0An/hWo43mtsxnIaAwRH69Uznhej0zP2rv8h6ueLWu+HhJeHn0M+ScQm91h
e6t5GbQDLsFphYYp7U66FfAytAQqVD5Ymy+Nnyp+9+HpNHn0WYCS77WqzVK9FyyHV7l5bcQU1QYB
fb4mr9KMq/2z8lmeudOzW9IvCBoljmUU5YF6sUrTKdyieMD87cDWRdexI0TJSrkcJjfUPXhHPH4o
1UjwWd5UjhqBq0UyvOBm9Dq0J+jBuODmnDkx4GxG5H5moY2Kb25j6KS7HD+rlnMmceqVPRPEQq2R
IebJS2v8VD617NGhyt4Yf7FPnucSOGXe6g03kgJMUQ/oEHi/fP97ilaJt6Sh02f0r9/D3ybebjqW
OCUdBm0M2P548TRrtmgPDSXmN0qyvGnxIDT8Fd9qXSoWrbCb78fsvkhWJZVM9ylv+Wkg+nFPU7PB
sR4yjOis18mrG+54b60cD2aFod8y80OGO0L7p2fP9QavjfL5GMS/mMOdDQeUmpyTs9NxUnyd5Tlq
mmyjI4wkXE7Z0mdZTPFPi9UZXuoGiu3mHUSI/6YeXb0Ei5/eL1kz4N6JRAckK9sq5xaC3C4fbwKt
LKvI813ucHF8L3G2uMiN7tlvg+6gwLtq/tqxoEFjEWPXMV4PPUBdnQae55XTH8c4SraTEtLa2rst
O6PTAl6WnJR75nPYbPx3jGdwTYTigF8Wtz1ik7nezjVcngQg58K5F1AfqvmugB+iicg7JPKZR4p6
X9bN/023u/INu+US0oPdh/7p6P5pmBirC8RmWY89ORLP3K3QuMQiJYJ5Of15o3+/Ryr9k4V5y95v
Rzhimtm+d5w5pTXpbOXJtk04XNTuSQkkhgcm+exT5GhjTj//oN8q7QJHphMqpz68VPhorgsCy8j7
+yGkhLxBo8pv42k34dHaGruvqGjDbhf/h71UgW6bZS4oA0PXZAHEfFR5Lm93OES0wJsucTvqbOCe
331pC+maJv4LMtOFDC9kNWcj0QChm3eKGYzFgDziji1hUUKOvgW4O5bB5KQ6nVoZ6FQFLB7GhCFo
1UX6E2eGvL254djVBNZ/nYiTVkVy8H3JdCcL3JRSy5qyUEsJn1pheoV4dGqyzwn0teN2u8cx1EX9
FxdptGLtmYcnGOd56bR0LFEfpcMiZUWT84g5ixijhyouZ7e2LREQjUZpXSB97PJ1dw/GKhP7AFDh
kg9rAyxRUQQWWRmhp468jR+lij4Ze6W7X4ucPg0XjuU0xiS/6wB8t+aAUywy92HmubQqLRNTnZOe
8cHVUjC3lGe3k+lhrdJGhp/v3ross4DjKIGUGV/PVwB3eOiphuYxy0WNUqSC9y6zw/dbl2Ax+GiS
7653exE8R0/zqk7muZsb3zpJIwRY5p1FFLIqyyVtsI1LPtot1ULyCDgnZqBS+mOYguStBjZJ++lG
KoQxNEeMzo/e+g+/DwCbouo7rtd0TNp9Sv/fXInRb2ifi3/UCjKICDIL/eI1vUYSndqgYHmNjSK0
WV71q8g19my0eZaxcgKABajxCF1ujV6lzarlB7ZZaLwTJEFZL2uCuxtJVehHBm33XgMcP3uwcjPs
OihLf/CQQUvYcB1uBZEhCltlaXrsZlRQEZSPFJb0I09ma1IFU9xms+6XcCaX7glyoUlVRQ0vL7yF
ByNQ8Vv+TMLS+AK2yLgoeOmKNSmk2BcrrDHPupTHfyVVTV32qboxGQiYS0fvoBSdGHc7/IItacja
hqNQlGohcTQaEgiQAMFNxM11Kg2Am+VcevP7wRjbFyGLE1GzbPjXQY7DxhcdUQz7byVD1t+gsYj+
nlV/zLhCEpfhS//x+J704CWgDfVUgCVI7BGG53lcENXDSr0SJ3sFacX1bQXRaZ4s6D3MWc6RvQIE
a6UMWU4Qo5E50zsRjjhLdV/Nz3Jn5p3ICqB9f7sBAL/SWE0V6t104JEXZu/NJSfuKdH/sLJCuKYm
b8k4xXFAx8XA2Wr8GC8kcY56aGoAKKGYs7LEr47V2avKCo2f5bOyjqKqRpGGzjx4AV0T5/1tyHAZ
u15RBqa2zIDtCi6n95jMwSZpHe6uI884bUTii7HyLJi73+h3HHe8OA6GEXk5ZZVRdavlh7acOZmD
ODQxDVlGP8QuwNjIiMlWIcwfntUSfgvKmNLssT9tDhJ6g9OBS7FImdmiDd2JDPWMXaFTklkcOMsn
iLHJtM2WUnEauAdsD5ulpModbYyM1QkBnXkGWiJkhPXHrHiAm6VifKvXKcj6QPBPY45h7NqTtPxS
j9s45SbqAvzid6NFTokvieVnCSYHMnK2MoOAAR+RZYU4C3iEBJ8YSM2dX2WJLXiIbbYhu8zyo6Jq
brR2TfL3qo6joYLVdoyvVqWU+SP1Vzw1u6RZKNDNRi+XQV8grPIokqAXttjqjqaSB/dZhA/7mAzj
Gh+4AM8ExldaYiOkn/DBI3hJM5q6/vda3uMLo6pvTqKJZ6OoJ3tFHJIhdDXg/RykmyAiJkh8ssAz
d2S2qJYjp2kF7g/pzDoSntd9k0kVKDyJrLLP7+eOBPumRLafI4+CmdlbuSaVBy8ayQpfBk9VrxOB
8ddDujxtgtkc2/GmICiQh7XGwvww5SNlLHQ9v9bj8siKyz5ATaQA49tjQl3pyfWOohyo0TK1Diwt
8xGAfwEqoc41FB1/izH0j7HK6dWLB1cMpdJRc1Zkp3/xhtuCHVO/m53XeRIHWpMdficOGXYzEMEA
3mABKdghwZvpNYByKpg50PqjX1tqZyhUiQTAqiYDIy5SQx9VeDrnh9m18W2EhoKNROa/+9iflcg+
hRkmOd2NA+x+adGKbiHjKCk/4XliZGV/GfODhngQeYxFFjY079pafxMw5goUKn6chBp94hnBgKa7
SR7MgKQrj15sgWxMCrGxXXLjg02bolZkn4Dw7WFwque37UOzM5IJtmYepamH5AyyENwb215nDNsb
2bCKTrfGqhj46dFhKW6ztCjKP1VqoPvQQts9hqFzrsLjqshk2TIf19X2mUEh3OwbUkDCu6ob3UIu
yTEx1ZmOKlZXXWJeUCegQmGyxa6AnItWQ2jlrAZw46mZcgCL19zgvfobw0nmsoN3ELsN7ZYiIALK
uW2LJ32l1dJyYpewVu7i7YcXv+pQ4k9YSrQb7mS1/RkfLsU6XiGOE3jrS5WbQUnR5u7fgSB8kJUE
4NO/cwqWRcnLuPW5B0cstQeVT9gkyBbQX5pOFCwMu8BmpmCxgDNsTzoUM1/3AZ0q8SlZrXzsYoEf
uthbYXPyGCfyWfElZO3I53LfGJoy+snkvSQ3NU5GkvYFDxacU9jsTAIB6aJZtL93lMHPpw4eds//
xLsWDuxmaph9cHeWjb2sBZt44bbhtXBBimi4YgxJ3ACzIo286Rkeea8oeJBnPLpA7yye0dnvTQC/
4Ak3+HcQV6SUdxj9dIpudhNRpAJLfJY2ttcYdH2bY8Pbv6tiAx+vNr22YGxg9udEEnHfSx/LChtk
Gc891k5OJTX6XWPYxz/ba/DRcrz2POMMwzcH5qoUPgb4ibDOT0EYUNCC3U1RRbEUgbFi8A+GTiej
aIZE2OeqNnblQufF4vyGBuG2mtzM1vLN9uyGuTKy0MQsmXZftyWK8+ITn7NBTdCHu8VO1reVrts1
2/tUqdcSisENXuTcrMPkvFwWLkg44ZFbnyuAKj/DFkFWYD7+0/CySANEnyjkrHuAqahXlzcnLkVL
ApKLq07c3WkUTR1LNJIdXRvCSygNU5zlM3xU1tx8Sh9GAFkjn2Y2hLVjquGEdRb6kLG+3cRWsGII
JDViEZuuOaEFgJn6dvRD0qT1u4pbK0WAjqhSe3p5bnuaOCintQcYPyuOGhAJ2NVjMRU6L0Q+gxTs
9YnJuc4QOdEMJ5DhoxcktMhYkFfOQo1Oek6Bp8cnSquq0ihfoSm7G98fD8qyLOJFrcTMIrMY0m55
WRDtw7BO0NKjppJCLpjaCniWi4fk0Z9/7iVtZ+HG+eG/xO+q8NhITVpLkXqdbpFrVw5KFx6pRxPR
AhmrmHG2ThfwNeM11k0saWX+HEfmwHbLeTv9+mXPz9yzJ/hKqkWZk+PhX1VqDi1m8XOVXlqQJ48t
JbOSHpINCGQuj7quxoLNoywHLNRb5B2wdlDudfuWuK4StW7KLyaXYAQFv68uA/j1gxIX/ns33jT6
jOGLO09hNJJT38G0zOnks5Tu4jzwSqcIf5zJAyYU47M92ESL17+1dlS+CbzUCvQ9EQ1R1md3EhN+
zz6WDvpPvC1JNAn83gOrZejTgXYjFtpKzbHC9a4EJIA4T5UGxVbfK09vObLHJiKtUltyHd+8LQXm
PybqCeIejtm5AH9ZnQnx7LtplXqNA2vEZ38SnDuA+xSo9EiEF+w/u2Ud9o7JTLwG6svhvJLijFyZ
jTTiitNxOsO4anqVAPWTBJ1rDQLF3+HXZ6H125LE9iKJfyTUNdNvPGPbvel+p6a1pxP/2rDZ/V9w
zzFJ71h6gtGep6iiWrxCtQupLCXGCRxEc6WiQhkyJDy9gx5AMpP15aj0lMK9H5iT2NN3RRuWP0A7
QeIxrVt2buYAut4jiWco4H9yBX3u/JEf1KDnY5waPyzj8aKXg4OzgePjBFERNS3PXfq0kjyj/64I
TSrWEcWvvrqZagOJKnEJi9w9+Hc7LE/vtJzzISXL7vvUJIA+zXniv5yL2wIAMGd+Mi3XdYd59B4w
m8DcqROE+hEN/4OK8EhypGjqgoCz2DB9kUZVbtrFFbAjb2HvRXN+2nXhfDpvOeECaUoVLA87oMmi
N5ptJfMqKaYlsBj8R2lBp8m6ix7tPiuIT7dbMMAi+6OL/I6Rg2uocu5CCnDRvxIhgYThvngbQOQa
22EdL4dB6Vrf7Vo3rrGm6Zeac58HqriEhz5PLiRuPTksafdtHMPjPkSZVR9b/KPp+az70dSHPFJe
6oqFScaC1u5+Flr0sypF1+CBy1g7kp2w2+9YFlv8KgC1HGzC2oNB+TFuDAq8JYSKv2AUIdfuTYW2
BhHWKQ1we1qW8rNMFRvBeS+KkGJf0SJdcEN2rkdPEauw5MmJTuP4uo5fqhaDCR3+GW/QvlP9nYkA
hPPVLx9XekvMPXb3/bdvXMelnhYV9A7Nrdn2leNo91JaCVt/je2XMAzJ9zeXgNcjKpbJ/0LoXd6L
/S0X59R0zHtWPvdLH2rG6CbKD86yNdSR2jyckNkOpH5EwkPTc/SVaWBi2v3hI4YB2LuG2/ZYvyi/
mjyNXgVpI0ibSuppGXNyLE3uSNv2Qe93icoP3k/quOIsK3zrnPSAmCD96YR7lG0GwH2QrYSWBn60
VFeZft+0S2T5JBDq13lZdyKR47r8XVE1igyXZugkath/kA8XJuUVo6qPBaSPk+VkSQyQR/ClBmYC
fAbPtCV1llD5tWE46s5yWPBTD+tIclLR8c+AL+902AqfztuJ4Zor51UogNWyXz91dT6pRxYHbKuM
3cPsUTvdPakREgouNcjQa9VKjAuVMt/hIkWdCetIyesEIKhAuWp+FFRNtV0clJcB+u2YIDVNRZYg
Si9FSUpdHVdTSXGo7YwB5IZdr7rUmNIb7E7lkohIz9Aej0HiwEDtUOt7UmJHdvNdoMWcSbixaDdw
nbYiE1DUajGFMa18ITDjBw4n6Cb25a5ohTy/hi48VJidSZCdzyUPhOxkUi7gnWXIco2wqNvpALE1
TRr9IdoQXKxrc8PIo1F4+f9Mp0LQEU7ffgawNHgdHkBnhwSTOkWhlSFR/RYP9G3l6SLWkLH8rpQF
CmgIthGXfKf1M1cK/bqOPbRXJGUt2Q6IDivRXxPyk1k77pADCIDTQTm+Nwn3reDbjaVE6nfn74X5
5fHt+eGPojSJhjZr7SPxceUSyADpJQvIut5kCndJ+u7FOxVO7tzluaBtZjepNjOI3eJshmNuRBXg
3QsQ9ugiGm4aTLQhyPifb5A9w4DlP+PhGhX6sGnfkfC/2y7r9E4CFyrug5lX2xW8WGQDSu4GWQOY
f90PrvO6DNVOwifIwSwXZ5loQ5LnPFcb5SW44JQSm2P9Kos3239xa1WRnvi1sWDxWMIBFa9HUHIe
4pUlgkxpzat1nqjp5zmVKhQx+FugOsnP8AnopiEzTttRsEaWymAxwDXA+aVU610Sz64RzaJ84djd
rGJ8Rc+HaVonLddOZjrY/P9UL1zw1qZv7dNYx5R5ClXy6ZzgN2WOfT24VHCET13ao4GHlUwm63q+
GHmxAaptCSAKw15I1+UVZh2KM2LbNrUD71FHZdGTEC2Dc5I5GXNCKI3UoeX26N6sBIJMQA/7ZksF
i/lT9jNPdKyzthoaBi8BW38IDOdalL18RZSKD4DxRePvjfXw1FjMK6jBg/1Sa90L0sWc6kly14b7
ld6PG9Td9ZpY3NCV3hcgZd8vMqO8Gmtdrk/lPfidfsMSu6W2Bmfzw6gbiBn6FGMcWrIzVX2aB7CI
lq9/OMFxZcfn3syhhIQgxxDXGxEOyvLNCSB0Zk2XLeZjdo95VNH3JevN8M7+uMo+WAlUSm2zW0Kv
0NvF8D8LkPd2uvSlBYweHYHo+jLxldCHick3aSZDuvy/pqWQObk19fRy2bUrtH1oRUCS4eeEntaM
xQEWpJ7Or6a4B7dmKORMXjM1VH+w/kKa9LV3lS45Z+Q0YczpkR50IYjhBeh8GSC/lpcI+SYKaDjc
NRR2Tqtgb+E6U9Cs0hZnj+ITxmC7z5ptNNrBO07y92E1QgIE0fCjAiry2j/Jy7iy7RGe7pXkeByn
lFm3atXZCxRRbgLJi0VupKzmSp8+Ir6OJOqn9e3cRlC33UFJT0ld95JyNHIsPkO0G1C1TVLoax/0
qY2SNqPkZzzqcO/iWr6PQcvgzN7573tyNpAHr1oa05Gyuzm+eZw2MKk70tPxxpWQSp53UgOEdBrY
xlGQpS/tx3JxQ+UuDFBt3q6VkycmwbYDfdFwvJwPDEtoZe7mXMi4Ukvnt4T1YGLaN71xCHtmn+RB
iPTZ5yOEGijxOnRDkBFhK6XuzhzjW9/IwbU029P52N+gx184Hw8T3/DBIyoK0peketaW7iMUeksU
bQ2QrRUXrn9YfYvjP5umxqM8DDFI35lSF0TNMomOeZrSd7bU+fKvXKTcb9uOT+VJHPwiKwuxlZB/
pXnqr9iC2wJdqLtOXiAFMmPoQZtLps+Qezdmn3+a/FU7KLDRObBxalq7rQvJpU+7wRgfMUwGwVGD
wz9EP48/ET8bGO9YmTzVxexRr/9nHk3GnDMDGuRRc1ERPFfw7BOO1CJRLhVS2OjuR9TA7MfD4FcE
7n/qwzL/GsufdgBW1BqrSItHDy2Z1MCvM0xEky6nYodEa0+CVF/j7JDKSDGXj+/1b1GlF26iqBT7
0Px7MCwVSmYilGbdpuyUJ3kG2Xcy+U5hzJWqtrXupL0jujwzcuE0O8RYQmv+QQNVgZ5pNwsAT2El
A8Rzw7CL9JBzCUZlVSKDJD19h+JM2CwxYr8eue+PK1S0znCrE4eUtx91ZSk9t/hdx7QdSZVgm+DV
ugpFZYw6OidDHON4NKUXSp3D1xqp+fwPUAWo4xoNkajsXABNVIGAmQf2w6XGFP6CgMpBIDLrL8ru
mdlsC3og9TgbNG8gZeQdRGxD7YbtC2/fqzeZHKTahjmunr5UNT+1NtV5BCONlyejkmX6lt2GvOAv
vWQSl5AkE14LmV81nEAKkBUcHqXdoyjQrJDBrEw9j1upJ1GIJIAQ6a2qT+i5zXgpr75abozNfgAK
ktYShvX76pcYmLEcs9ENC41r27tMU63kofpEBm+kaLKKpE9WvrPWGYvqOpXJHCZvrVFrStlzODgk
KvpvP2sVuH/klMpcW1O3PlVhY/IOuWtST1NRA8dpfGz09WZJ1IXTpVC4lx5cfiOVvOiCT0R6o1Fe
T5T0bRzq+vq2zHV2B8rlsONKTxF5XLAMTFQ5tmFxAM3XpOeGWJs2I75GKIKPe2QwSctfjbOP0TqC
BntEsBRXRJlzr+COAvjC4zO22H7ZBwkUaMWbB5SlBUzTj5ICLSGkPXj6JkYiykhEtv/qzzlp9Mj2
gU/4hSie0s093Y0rMW1x1XGrkr5mG/eLuTB6ao+ZUXwLx+Dp8i82cC1g1ai4FTTK/kRaAVsJ0Gp1
DEQJOz3J6ir8Im8KKR+YUvIfz3kQOGKXrqwtcsKJjw+j+TD5I5bjdXetyi4cs0jHroB/EMJCDWyy
dc5sHDtzw7M6ashrwh+WF3uYXypMKjvY9xIRj8CL784Vm6c0EwUfAPF0CVnpWQgbAOh6eyehaFnL
cj95cQfxNFjK+/2vsMwuUlKKm6PfaU42lt0OkRG8O6k+obVAuQIYomMQG/VJgUEVonVIx3m39/nb
OdxTeY3y07++qv+XqJ6aK+eRQfuR3lYe3VtXJK6JmI7QpYhj+EPMSXGH2CwzoamPfBDnxp21qEC+
TjIiEyNbt7NaWb3bX4FoZf8FE3y7UyHaQJbWH9kThhSEQopAvB/ZJdJKgbRE2uGz5pEdCftOVin4
5OznDpW026ET6GVQlN7+agrkga3+3wBQUPhGT74slhenKuSKDPqn871QbY46XRaQs11BIl+c3f6B
Np5MPl4NhCW6Nz2wTzW20Hw+tBrqB1IekwNpUZTx/cNizLdxS0bPEJ4c0FByqnAFgdazVCclW89j
cf6Q5OSeJBGfFPI80Jk0lMFPm5QBhz0DIlMTVT7mXO1PncEdLVytrRXRGeuG0kDO3cMxHQZ7uPiC
LDD14sy1ntL0/ewvGSWbKBNWqrxnqbalufzFLQnpS5iVVoq8OQrwLkfoBaX04DwkI8bbZI0wd3OA
1w6sOXVEl2lHiAet9BTA3VgEgf2ca1Ia40jIEMamU5N+TIwxkpo3relGqmglCgCAOHzm1r1Wuw8J
l7JyxvFXV2ZqAuob2hUN65bDu7mAKHs2iDBW/B6t+9EUYQwa3puuaGwUOnCnXIZUAGHZtZoG3gdF
pbypIddK/4lvDqYYUz3Bm05pEKYnP2NjJ1vkQoLSTyPcth1o81CUR+Y9YfNsVDECDCl6lX5EFDn3
eTTT5K29uKADIK8NlVYUlbdka4q2vFY+wt0CjqYd9MXOaMJWg7MIdE0IGxYGm31hPL8P4flb9n8N
tRO2VhCt4E4UGoy4VEifI+i7SmMz0KT/9H6fedKrmBuOdENOLtGLU06rr/2kb+B1GN6ZI27/pfzQ
DjkwHhWxmq1p/akjYWZC6lPfAi7upVNOjOuzOlXmndaM1/qooH/auMlGrqfk7wfvp5f0HEn0rTME
JLWyCJZuHFID7C+TAhCFzoTa84DM7q08JWZhBDAKnjrZNrns9yW6axFfYSA8hfrc3DMaAg0Ebm0r
U5+6YzVd6KcevaU0HM0/VWnF1KiUEOxygY49jvY+yYDBXWVqv63XXstANHlpo4qLNUYCQFmW3lU8
aZKKuB/7FX6Xh8uEN+ifliEAc4lrBamQMJCyekoFG7ipftdVkap/TcsuGPrMy1ckm4LQM/TZtxfQ
KUB4Ui6rLL5xEsxSNavDlUwKqLWDhxetTRboWlybHor6PbSE0fPUmcUuli+3W5ltzrx6SozITtEc
Edldc0+bA7eI2SDdGV8hlvCkByS77kXfoizd4ZgrlX31kmafuWao/cVkaFLPJJRJW8ktCQ5fLY13
VDIW/KkkVIKm+DE776GjiOVyCHKHcj3b1AwYEwJhHl6bDIp/LwgKH4+lB9PfhdLIlnIeAAUpxOVv
5ZntQ4X9UaQAGYNbiNbM4BDCcH3sP5SD4HrwFJXazXvazMdsNLOTok8pvDqVH0IWSlOSp8UOxWdi
pop+VnOVhmIi0DePoO1Geu6QkN9jAcjaNFji1fZQcPci1ZFOYDtCT3WOQdegexsv3dR9XsgYBltZ
zsMAbu4mXDK+PPl+Qeoc7pRSzXeWObpoPhBKxILLeuwGvtx2OpN3B5n4oq3Ko3KWyHS8x1XsfAEt
iiv7r/nuzuePuKF89euiNfc4gUfznhVmBPhIKkHVxj28Y/UdPvv5Hr/PvDb/oEW806n2E6TerQeD
l2JnwrygQvELVvwBs7VlOAjQc3zq8ZRcbbYvCQWtvXB+6SiBpQPD6lvSv91dRd5mlEbTQVlLltfu
kSfmf9pcZSWHELk7HOaUUjgnGfPDTSoxNwe2Vs0uFyMPfnWLvIb7Qfomyu3uxzWweSHqLiqqUIkC
X5U9CwXAGZTzejslsUy4dOoVdeR3RUsVfBwYxHuGMcicxpbGwXKswrwMpyfl/wKywo637LlXJ/qx
//KT0QWV7MlqXwow4iLGUL9PLw3QHm62ISxtH//cUHk6uQTZsE+uzqay1B5avSoQfpGjdw5LHgJu
SgFX25TPBU4GRUM733F2P/qgFQbfaemA1+qoWYv3eV2tY93cvWGkgmq8rKD9qFSzWaUvgGR5Pei4
MtJ6cb/qf9pkJ32Dkf0RRuyS0/60nddonaJNcwGI0uhdJV+/i/bPyWEmd5KfrEFRqRlPbo7Ci0Cy
3iojMl3LN5VrhxWxDbGLDH18mSPd+fIsO3cHa9VZBB5dLMr0p5yTF6kgWDsvaRagVfsqGaSmW2Yf
SE1Nt2KVFO8+5PdpORZ+rq/G7qXdKEjziAbRkFIx2zZh03/kE6225hXcpQFQsus1lKgzuYLHk+R9
LryJ/kOmp/Ens5x6THjEBWp/cP14+ZweNh7ggAQAUPCrec1ky3VWdwdHGBy1Z+RKKiZar/rggroW
nrirJrjeHtj2dSndpy6hgG8qQ4MH2qS9ds6yMxWNf0Rcp/QSc88uLZOiygOVSpGWfRSFKRrfYJk8
0lgMr07pM+HXgJr4GPrGZvAhLbXZHDhSfV3sJUbLJrrRNKuvRGEbe7m5GCNwP90oYseZhf12b+0R
utqLFgVMlU2Cbz6UkHDBvuQM4EowaAhp/2yUhTxGZa4qnivTP5AdjGruwrElWWNbkgDjR3QAbcdc
5TkXHS1IH0MEsamzNano7FURocXFQnkiT6+1dW0B7PZ6SF1Zdf9vqFdH5RzvIFtYejtzMstg+EC3
M/B7Sb0elDzQzmH0gVh1VD6EE+AxE1FTItuAqajs8URrMV68iPfjhNilBo4yPlNuLjxi5SMfK0sD
yPxIs7AvK0x8DjqkK89CPGqqsPHNlKezzp/1l/K/gXfU+86tZcSOkkkySgKoNyiakNjJuq7cEJZz
QzUC7S2qECTIZFQkWVFyMLPRstLm2DmCl/5TWBWJ7pw4b6C7RlrTQ0S0P/0OOMs1JgN81hA0dU9X
ZNLncsJzkRmmYHvtC/zlScb2w6sZ4vBQ4mEQ8riCqwt4FNqxPXdQ7H8ZgAo4NeUK7K7fJ04OmlIx
hVYEprJ8el8Cr1g0mTbwZEY4F35vNK92AzGYuOZuaOTuIqf0Ti+AqQ7VuRonYwHxENGyjrbzomxO
RNC2QRbJIZLnd5xo4+5Lm75ZyfYSHo4nGUgnnjBHu9NIIjXcRF0dScn0fdhS4HyrbpzhHaw8ubOh
mRzr0vwLPDG18qsOgsRpSefeaEh375GjBP+mlfZoaXsf0ANuP4lRYNOCw/C6TL2LysDg5yyPOOOS
IkpgHI0Is842WDTIdiQeCBq8LZ+6BoqWHJ1nio4p4pg5LmDUDC5yJuXj/COtRXEYJ7f51VrPJ9DY
xPUnnRL7CcnTxUJpkGsMFSbXrwfkJsY3qIQv8RwflwwlfdCtw7pecgkhKJmn1/hAE4/KdV6dbMlO
3FNF3d7qZF1yQbfDIEWXCABz4j8+20ZLy2XJWcpoq6qPrexQljZsrKq24ZTB34lE8Eor4lBPUR23
W+vvfRHG86rGfF1TwCo69ywQ194jgqbuiJx4IAZLNonmAvRKqwmvDG1LDVmRR7IMnzz59/JEyXc+
72Q5iNmC5LtyKw7pbrIb18p5Sgx1rpz5kFrXSiOjryBW4oQh+AF2hy0XLcncNdrmrVH9JeV+RUUp
cVtZ6mXTgdY0VN4FSzYop/nu/PgtLErTTgA1OH0D5JDxoqe5koVLlEpo9lh3zxC8ynw6y/VWR24X
duWj1J8nbSEpeNdw9tap7Err/NtLgnSocbEQjSVFCLaj+KLQoxVCmDucl0nOe8K/nzHjmpHr3woR
JFys2jegC7PaSUhFB9tSdd4462e09Dw904thHhKxq6UpHXXA4IGWchXdARlshGFe/EGtKmMkvI1B
90Bm36lUCoxjOespH217gC/qL2l/2fzb1r7gA2f/Q2X9Q6xWioRMYmG9HE/QRMiInIra3XmfL2Um
fPKitII4D9JwMhU6pPWxqVghnYvdAXJ0xxP+V01JVf42ZBhC2NC32Xq77Iar1itSfi9hdEvmLADa
Vj1on3fWmDJ0hC93fcmNetFryZfZPorxUIgGD/qQNzZPZFFg/5jNpVfC9ED5yIAuWt50i0Kpspqd
5/6ygtXGaQez0ITznQnCSN/HjU64rjiXhxailsSgqjwSGC/acxxjZ+ksuuy+qCvAL83mZLKEs4Hh
JzQo+fvH83uFbk4kdvUOWBZpAr1qiSg4m4VAD1AGWJbCobIUxPWKM/6gXce1kFKuHzIzV0KDm3dq
MREuqCTVa/SaOsq4/Hd97CLlxkfTYKa/dqoA1yZiCqotfNh3tm69rQUkKXDX8nGhHObnJWKhJLd0
Pj6f4vou5fRWSvRGCV50buVJOPSWdqiUNN0kHcogKiS+SweFGZLaGn3fn0Lg/KhtZ2IU3apPjWX/
YrPop8vNv0KP3a/ljVSKxOx++E1YHOWFxe5NvHC/m6x1+k+jptyyxpaAZwy2ecbIcz0Lmq4io1Xf
75FY1cMI26G4txm1ZJ22o7PEg+lbeu8V+6o9YVA1Ict4S+hMqK9DXg80Lv5uaORpuYweWB1aLo1K
hlzpTSekoBaVd3DYzD11zmAN1aprvby+hSjoBt9FCKV+yLWCDUnZh0Dlu8JaOOGayd3mu5ekMkUK
rlbk9LjmXIjz5+VppKDvXKT06YF6FRt5XnWQyoMheuoyUnPzqXMPmuXwwhGojooNHGrnIm7TE0oA
CEqOy8ySKIJjjSW+S+GRgZOuKMtZOwxLfEUEJB/E2mk4UY/+ZA0eKVWESOa9R0PeqKusFMqm1hxU
XJE0oYa0lOJAOhQ8rQNTh14VVX6laK68+ahkEtvI2Bj+CMA4O88nRAVOIpfo5BAmqsktTrqcMPih
StCXzZ16KMh4ct3m3MqwWAfvyeIBD0nOF4xxuqI+zgjZeIe17fbL34oe9AM3dWSBLsjfGHuwf302
Jg/TrJvOJNQHebBPenTqH1He/y9s3UvC0pia68Uf/5gWQVj9OTvk4CkT44FangJJsbYg3NIwqzCx
l/oBYkmfv01hlPU76+nIxPDVEq6jJW42BmDjW/q46hnjvS94XQcphITVdTajhqvMRWBjHWNqWaDU
4U4Wsy4ZfOoGbhxJP94ZcL/1y9pygzyVuZ0hN7lueW9iFiB71dlmIHNelzaOYQjsX24rk9T2i990
WlV8W4zB22tIHISrbgKkfkXvJgJoPRoJ1QFDmGOOkAXFz3TDbJZNQHxWUrLUsYDve23n/N57RIGX
aMEz9YANjtSN9VZ2UyXUQM3QtJwmuCZtcJet+YyXBRuAJ66eGIH5aB0kVfPHpteu+qHp+0YdxKu/
uh2OapSZz1gItyrfEumML86Vz6WELLvLSFPyK77S+JbV1thxvXrVuubRlFeGv7+hfShTK7Ej2v/E
yhUN2ZW9W5zaxNPGE4X4veskrvZEIX5Okio4s7E2uX+UMr7SDSayv4FXbRNWFGxeIaYhUQvqtzHh
wjo7IqNJBP8N4s7axUSh2vzFUHHgwwYRJBmLqwnunwkzPLduDy0Qa24w8y038xejNenEQEtfYddw
Gi1FlGxKuGeSZsQ2FFaUzVeb83Y0vUMDL+7esAPo13DNuxsAEauuq/3vbGo8O01Wm7PYbeN/vNHj
a6QyCas7BL13C81LAR9QEHoTm0RHfvY0s87hrIPPfuePrw935+ONh9hcnCoUwdDB1RnRHlkjnzJg
dyyytwDzRxGouMg9O3MxUMwtwXS8BdEuqW0w9FxrmvtBFod031WnVRxE2fgF1JWwrhHbvVi+0CDd
WO7/EkrMIjDHGQHxOwpFCRYZxUpb+LCiv/E886s7ZeQC2ufCve6O2K89oO3z1SAc6m6SVgNiJfqd
nYpfGWlEZM8Wsw+QbPaNzVj/wiT8k8LCrz99dAJHhxp84HdK3PXl+FxNiLk5hJn0S31GKnCNZVUq
fpC2r/S2v4vK7AdCJNFoOtD8lC/uo2JLEkAaemb4KHqxprtunxtiwPqoTEQKqldO7qYWUrdTlCgV
cwLg386gHHlMtLN0Q5gU00tQ/do5N7VsganLpqn7/BcAU6GHbk0He3rLDjVHLbJwsDXfuDB2PGcC
fpV4Cdk7os9q5SRN7EgIkDNlikeJp5gS9n+I/i9/frT98BE5roXy5kSF3vGBDPcj8wkK6li5roTx
KaYXoAOEMTgtHG7q0g8ZNBhxDDzF20gS72aDKDLFex23C5it04E6zbWXibxhWqj82bvuBJCC+ayv
KMPvd/hmYr7dyOnKR6LjyTRh4g4Ur1uxqHcGbEp4VkDVb3YRQwtuMlZXvEgLTUY5FVlROkaDx6B7
LgdS8sprFOmxKFF7SCd5+9lAGsH3rSdRCAlQeGdLoXgZH6ROBrYSOByD77KoOWpiR3mbMEfdMPr7
mRrBz5/TAwQEb7+GrkEDbDOyjvw6oPqlg/F79b5h/hauqeqr5LnyMvZTx/TGlf0fJV0sRd6QN/Mf
9/+/Dr9DP8ebAKdtNipHJuWvLkABHRLkvRWaR0fjA+nu+dlkh8Y/EdZIeAsPnsd1fRjIaQV6jYgw
sQjQYdK4Q9JKoo12ualmHuxZEbwC8gN//xmMwRs7UdoHR5Lx7quMducWHmmBEANe1PFiHvMa/OQw
szFvFxcT/VjEyZHGYaANMhNVt8BjwQW6fHs/h/KWmoPW6IPQuFI289jg1RmD5VZaXmDGxmYjH6xI
unDsYRq4zbD98h+muEE0B5lJaqtCQTu9weFSUV8mMav4qSARyXNZlpQeXcefIUp0biSyW4WDohfa
+UkPG/NmD0T54445a6Uf8sF8l6BUd9YtcmHBagswjxqYNTJr7cwn4NsJPEANyALByvxrjiKt7pZP
gKy37nb54PYDlxOA/Lh82ySS6NdrCgUccZs0N+gLtEsgQp34c96LNnTFbBeHHA7Swl6YpNd7BDkX
7JbIiborz2rD2Yangdlq2tFF4yFZ5jpLFZnEfiWZNVXrU36nmsqPgd4+s1fUDx8b91+BgfXbH3Tz
Ip4o2scQVOKbVfwsIU52KjXIpHFI1UKvmLFH0AF9agxKsTiLxQq22V79Mr5svpUMZ+T8+Oh41xt+
DqmiDJy+0/Q5CMBd+FQFMiiM7nRu0r9XAkIEI92ItbJh3bS8C3FXibypp2vUAUiKGwqEYdsz99aL
1Pn831esT1XsNp9dkYiix3wVRoQpWCJ5bE7Yh44yRXJW/I08xSDAcIz+UhBYrLvKptcbdo/3jmYx
06tVlVCsfL79LvpcbooPc178rXk7CoQC0MpUHXIxaB4SGKuTkm7YQ7xN9gbwkooc6ssK0GssojrM
h12O/8aFjaQr3lBAqBTYQQifj1sAFBhJihzX/Ze/urjxwdqoVyGDsQElRTic6L5xkZ4dVBpAXkZS
9izqxpsPJmnlIZPeAtA6qSOloPD7dYQmQPY06A5Zv8hu06OCQylCd9Hnf3AlhNMqeeud1jl59Vpe
y7zJ7eZPR95I4GS5yusFgwe/ufae60q75dhvB3zN2lTIpJbd3LzmFIJWZ/+iWq07p0i0hMdV4lm6
oMt2GkZXXPa3ZLgY2y4zt2Zf6E3HzCPlgFeWLg2rnrPeLT8eaV03KzENbADMVbC4wKvRHCEy4Q6O
UOy4oDeN1hW6mgJENKm8NOHxLw5wX9+GMa5+m0g9q9cJDiQDJUhqqeSpatlACMaFw/So93HKfqf0
J2mILulI5Oooey7vRK2ifEmiUs2IMwOsGXcPChA8uQdMbQvK04aZqDVxWvgG1eTqg7Txq8dgEbAJ
zljky2L6yUXA8Ov0jTXrfxRW0PIA5xve7pYmIL6OirnLwLZFA1HJoyUUlrav0hYE2iUQQW9Uu/gn
VBRzD7RG1EnYlrWpozIkcQHrXtbTGmrSnlB2FO6WRDwnScwOPFOiYWJuMMcH0h2SClUaFaMN8tqj
XsRion2rf4JiP77SpXVMrxWtLOE4SJv6dDSA5nYRw1rjw+OAw6/d667e7cVI/C+Iw3dw99I6h+AQ
o7mLmTRqOvqnRZ2ZnkJBICh9FkjeEsI4CA1dHWmkkyxMoeG4FsmXK0sRO6X/+xKdWEPHmyN1Ijl4
HeTy9MdcdtRCP/zHP1WiNl39wWnTrZyky21W1ZDkKw1gn3iSf6V28dub+1lneViUrJGV/SPiVbdx
dr41//kAIYKI1OMLOK5Fr30r0PDhdu0g2iKVA2BOL+nR5HpAup9N5HiFdhyABjxIYJrr5aDTCVym
XS/EA4ropcZjl8SWw4L53T8JOAVlK4/0fzeDutF/NK3JzyxmmGpwMgau/mdNjO9AHR/gQgK5gNHF
g3FdfMAYsXzyB6Gr4y99igFz8Eqa9R1lzIEdh2JIboZCvGmdrl5PSKJx9UOnKarSKShxdnRXNdBy
vzll4m7agNXedKJXUqrUEDjyWoaAO5l5bgfbdgcnHpig9TbzrDAi8ZoUhKWRLZq9igQC2LEnnOYu
6X9TM4HJJrkjklO8coGkdR4CZqqXg40wYS3d0gL5GfNSV2EuCrNdaYA4EYjlyODLpo4xmQEhQOOo
xcN0payMASPR024IRD8nBoXtOPehIzdf09jfcLcwZjujXJj3ElwAqdbwd7QpG4CKJYMZthI0wqul
FySYY3+ipBPlelT8eHv1GLKf7RrHN6qPcd+aWbBKuGJbGuy4h+K5Yi1kLBjMZjkXxeiAj6XaUV2o
mgRTatebqzXp6m6A8n2Ryq7m2Llp9DpGO2vixNdbCQTO6xQ55ETOyLMF0XqN2MVaGjiu5fCVry2i
qx9R8AWH8+dvuauhUohA4Ohlp4/WNhKDdDx42CY21kTFBBCpLWaP5YklaiFhqbbgoafP2Q6aB6n+
/zGg0NgJ2Uv4/Vxzv+D5XwixiL2VLgQvH9A5ADZtPQvsUwt1MjulPwpHMRNztzdGFf4FNGocfcTA
yvbevM22BfVdUj4E3Fq9kWxy7GodXq+oHtgERQgMkLOSbKlFgDaEszPbVisjAQfLHQuPnS1KVLad
AlWV582Rm6IOdrpuODsvt4wc2qVPY4zeKEzcH++RRvSAHu0IgZyqek3U5FQZURMNjhB78GC4MjSY
XRT5gjx2Kr02Wld22F+LwRVw9KgDlb/vPOtRgvPy+k3O8WUPHXFgGlvIJ026G5PXoaSl/GGtXPvs
FEf7fx1gAdVZT2T5YiS90NJCUi+1F1v1/wK/wz+3WsvxWH9xwYiZuc759bdsBFVj0GWEQD7RsM9h
vXkRt0AAEz/EvZK394Wg1X5QBYLqdMTW1DesijbWjoWptKi9od3MEqhDK/6Z4PLAg1zHwf3UiPmq
z8Glc8C2fruedx23uog/q8ehqZkk4cI4NDfI8VcrsPdw8orlfsMZTFRStLTUqvHUvO4PZrP+qMU3
fvWS9AHtS9zCtJlu89vOkf5HbjZQ5eRQRG9wwN+1dlYFUiLm0V0jHjExMF6bdWjK5smyKAuraVvd
Rih0XxOyaNH468OvHuqGN+a1+KAbERKRIROsubTomntpnit7OEFIO7CoNRpuFifYBRXomVNoJ05b
LRuPR8H1OpkHTbJ4mTkfDAT4Zx8AGoxwzlxm1Y+UW0oMEUmrhLhKyggJK4fS7+08BMipuoepTJEC
/z6UJo8hh8Rwwm5vfS/P4idlNvcdJgW+cHfwV4pCLT4IMF4ZK8UIYHME3d7b92Rr5rF0hImrN2Ou
O5o8B/iW71cju5lp3NOnzRbyYlzBr0Bb2i4ETGDOJoePd8GrquA+r6naUdGI492yRurgy0VGgjTd
RW4wbr3xmEzq3MDriizrdTcigVojEVbbhWodSBkmxnOYQw2+GT0qn5uzWJxSvzZELTwfKbiOLPmp
I1mll5KIGdNQOtlyVmOyu1ZG9RETHPiTvKrIoI9PLuy16JBaN/cZoczP4XHAk9QsEXlNeTOdztsS
q8FDObqk/7GTCBjaejK00Fjyc79GEeqVdy0IFc1QdPXhk7crj795QO2IE5EfmmTgiNrqtHOfv/GW
jWe1Q9++PgXPPpCnMZVvw5qeAIuDj+Xovo4h0wEzSByAQwmrkwzb/F1exBTz04srrQW/0SDO7Mn1
F+idkOeKdHgLQe4d+cQQ+/rqJrz7vXMy5NwkypwbBUwmUxu11MTJtWFVEXkPqEPH7tJ4alqk8Auq
KgUFyprnEu1DgYPODPKKt/sZ8Ty4IjxwQf+6QdtDjhr3+DVRFYs3svBgKSj6UbnR5CF94A2gMWI7
rsUAh7S4rO/k0jR/EpemwTkE54Occ/y4T4ZLMIL5teRtwr+4OakJMBJg2pCM85Fiz8ljzHAueIWy
KG2EqMsK3hcrWNjnySPFwRNTwTtiycDXv8KztJ5hGyt+1h2eYFKpsmNwCkeEygEm6QYIATqpYS5M
V+yceLWGRVxDF4t9FS6R3eEeC1KoDBTqhyMivcEaX2pnqxTx/SKGxbSZyEEYS3vKBq49EeHQEsMG
JbVrBnkPgOrtd3lhhkTvi0OYkyLafpQkIV6PmXjCFqDuQPhxDZUqCR32Lsd78A56ecDAFlpQZQ0H
kx2e5/fZrq2YTYqH1IPpH2YP5ZzMXlaJIDvTggcFTV8Gk/ybbBDiNdGERFYH1lfQPxn0foEnapzG
JQFgOmdR8b2g5buWw1t1kUZ33HhGyjtC6FOn3pYWPR36Wf1tgdDOrBwzJskB2WMKdrjugSbhHwdJ
re3dUueMbQHRo+JSCX9nK7GFZ5ulTnCsw2ZE7o0zgCfQ9eelj6C6dkjlgq92bSydFkykLWeh1ScP
cfxTJuXh92fK4L9uARytzA6+6EyVJvXzBY+XzkaAEHu/wzZwMm7zCElAFxIq6MDh3ag4ZPU+Aucv
y8JSHVyQeidUQ1Ls8s6Btb0qXWY53qmwWgBzAQRKQ7t0Ibjud2aZBcvRionvrwdsvR9qQ0uuI337
FS5uLOEwbZIIkly5rnQHV4rQXsI3un0begrGLiMit1BsDZGxG5575180wWeChI+5lfkWoWF+tCzL
24vBtgJj1jGChEKH2Mvgv1BMPKqjh8emB7HseVZ1+ae9ErHUbmhN0bCD9HCmf6x1FNjaIqrxrwjX
rkaFhAr5ncJqipecU4XH+JFU5kkOoHqYxMm9P/Ri7nHu1p3wRm2rPOBIC/qJc8CO+Kx6lgVAsZjg
VOF9Hg/AW7wL4sY6AFSDjg+yD69F6foAnvH7qapo55UzrCnKe8qKoV90MS2611fEFjFeXTkoFJcn
7CK80pQN4K25EXectthHIuJw4KL6Mc0CHVHKjsCpMjNrQcZx7PWtGKvrHcNAKqIebqqtW6Usw2K0
AtVYhNJH/2mCEA8IVaky1p+av7xIZI7qfyIhfYARD+mqWs2rPlw6Ay1cEx44pDDfof+SogPlMaWf
P9IDKaRSJOGejFoqB41cZDoW1jqcz0m+hdXdjcUPqQh+C01p1oO6Yehso2NSEJk9D4gLJ1JoELrk
i1d0A23dai4/hSph7S/yaoVXdcWPtHlf0Eo42Ki+7toirB+Hxaz21RyYvC8Y+vuVJ6yVnZIK80ln
wSZotlQ0Du+BL+E51+X3cMHV0VVx7BsrJIyuzSSBafgudk2o8SsV/iR/sAMPqpz+/TO2qaAqMmBw
kAeIvQgfd6sXGQluQVonyBJxcfbPWRoXjWLki2PLtQuyvYhAScL6Sm3VK76hdwMFTCkJU7RH0eo2
HA9NfOiDBk6834Kr9NT1IqOxJmJ+m59eaKpHvSqd1lT20vHt8Qy7uO90dRK2s+f6fOhhIXNAgIHx
RKD9f5CP6MpRh5wK62dKj0+EmmKAADcBFKoSzmHPeNIP6fGOrcQb5CjE5iT8m7ObTyxy2l8sA6dB
oq7V07DeNnTQBQyQZsmIweKeF/7j+5+fTmhnVaYjHrXKPTTZHaJBpty104vmtApEkiB51/qDtVRX
4eOhW6x7dzmOxVohdFrXi6pBibEgVedRM5VOitwD2uPKF/pvVYmhFRz9gxR6U2grLD8Dq49gB6IQ
Uj11KlXZegcMjpZFzQeOmT3u5H0soH7a9CbHSbEFHgpQQKaPvdfneML/FfXHr0ACFIgsi1oP0hnI
f3n3mMoHmkBQGcMfrfJHdco85EEQoUXWuowxoBHswsxtun8+gRVfTzW8GDS3RrpQVcr8n/GH0tMw
zwhWPcIP1SLeynWUlqPyfZCkAxOGBil6AMiNOBswuxsbYe/HmlRUhbkCUmcD4skqImMhqaHDllFi
VdnakVAW9VD45Y+66bUQHGNoGUh3PTTih6lQtuT8hNHFsvee+9S4LoiqYVHazz8T03Yeffo26Zju
yg4m9QK8qH7W4PzpLPEcQ7qogGXNzv0E9hwLoFwPme+h3NrcfcbW0XWsHBDJ+98KWjjLcHJIYGI+
1AW/4aW/Ov9hF8gvHPSG/DpEZwtViCdwyMieydfOsmfSSwFyW6P/IjByPp3an0VXxcwHOdO5Z1GF
5e3/eb7NRJjFkZmwMQ5LuiV0uHIl8j7qL12chwDXqIFqRtNRhVYYIS8eVwL1xl68+1BOYCV6ynIZ
iyoaq5aEGj3TXCkPcVF9dhR09TI4Y6V/enbV1TMS6EFAOEmfZt+8BsQ8kYop9AGUyFPqU4xU1BRK
TWLnnI1KR0AtjC+5/7VoOCWWwmfPPpbANjzup6UAadH9O8s3nSyaJ4HZ7+lgWt+2EEo/U1e63eHn
hJJMU3BrtOvdGsIq1vOqY6V0g85rLCFsae/7jIzGlcttt8P6TsCzXOvkPkkNr7XCEfbZRT8Cwyg8
8az2EV0WwceMdVZR5eJ78otkZRx02JWaNUKfpMLp733PfIO6Y09fyWLgaUR76Y5ncmEYBH8usWGC
gcxFpihmA6WmAjoFDxwaxsjvRfetEtPI3XKIrxsINYrElbyzaajhFnS9mnpjOBK3zJcQPS7Seifi
CqQT6aYQmP9KZzdLuQuqnQYXMegUYVfM74ojGlEVuTBn9xI6nOywU5g/0Nht5NOxZuL/6j43ujLS
OzmodtHH3itIQIWochUqI4khVm91kWrDPHFPQdrARsq99a716DKVQTjYwajdmQUnxvIzewhsKpM+
eworDpNFXW59zZvEEv/WPqHrvNPfX57iuDtWJ/zkwTyE+wldq/0frAc0+8swQA/Uj84vY7dMjMGM
G5AtlKBEAU/GrrHJ3P2MUWjr6Ftp1SVT+5gnrjQvsjDPnuLdz4Hz7RUvlXC2p7ldA+AtuY5ecPo+
RTfBwqQLhWEaJBtkBIJSATQVmSjB3HL2B/4e6yiMjOXgTNP+qgidrmsQLgs7hOD3kyOzCJ1iXVAc
TJZE52FboW1eRtuZKNxAA42awNMub7g6xSoV0Vu5j1cBbxrocBLveu6RD5wDgKAA42k/ur08Vn1+
2ht771b4MH0mPbxY1Xx6gZRGMBLWzx6XZJb71ndjW8BMm9fFr4qWUUF5v+DUnSsyzyuAivyjS7PT
O+Z7pFFuHv/WJZU8mgo5h7e5RvcgSFQE4YiT1mGIjMM//UOttV4F32TfRFyNA3ySH0TMZAHzPjG4
GeuPnHklr5s6eCSFuNGsiWbhrl8fjjWbavot98fa5LpEZwPg2YCjC01p6+D5T9Hu0mtdb2NHu3EB
T2nhQRD/1DvdrBNpy1P9eSefNrIgenIVUkW+ScwbhGzjn1eGLn0vUixZXZBigT1QOdWPWVGdRp2+
k/yV38xQpzFV+sblJvHT/oU5tYi33VZlRQw3mWsYny8budN2lJpv/jU9g09Cwvr7Xwde8Rb8y4NF
QKRDc6gUscRBcaq8gQL9WFg2OqFHoPObdZJc2rm5lbtz0bL7nEA7HR7AiC+6udSaYGpDVK6PKOu1
njEIg/XlFnxbyYVL+Mnx924UGOFES+gh8EpdLdPWkGAWQxADFYYZO0FoHaNSAZVQDhj5QqcRRaAo
4WPyOUpI01auptsixAucWlw6tt4lFHW67BMUWc4wCmxUDptgOj3Ks4N//vVdLAufOwU6ctGo+PvB
orVh6P3yt4cRB+GVCNempkH46ioNowffouT4oKeLWoO8EjDrvE3MOAxHClBGn0TlVETPqsF1iorC
nYczRnvy0jJYk3t1PM66I7NIU4JZpiH0ms6xWh05WDCXwGFBOnpEZFJRVogNAqdLvzP/swwjxHn3
g29e1PJsKPBbNK6jeMJzSuYcUnNYUh1B239ZGZplbl6cbO81uXKkXKTpCrVyeUbHcoAc0rNOsUWg
uwop669ZDEaaRrpTpKbGNmQDLpCcfMNnUu2Ejizht8t98wqOO5zkSIrrQM53MvOQMMquoaYgnTY2
OSWP3SRwe/UcL6fpe8Ya4+uZE3jyyG9ynwCCuc93WIFPqksdj/egS7ik52iw0l9OQtTtasQzFmLe
gjOWOsGzaOL8LLxrFqC4saulS3PDBsid8o/3RT+AHth5N3c/dHfPi0CnvPxhJWWL85edue4aoxHG
MKJPduIVNv5T7BOViQnJCpo2EtxKjjQ36YLNJvNtoqcv5FjqPbMALvG+/+986HqvR52tAj8yi+o4
u7CLRjrr9rQEltybdwP+HZnNvQibfZ/OirjHnuZqZ+CobEI5jYNpJWN9fthXuimzmLOUphQC0vaY
wD9xfxXN0ICqfVXpeLiPYo4xvaJNJqwbWx2FR34HR9Jta+eE7Z49ufdWxjOEnnAHpPUn4cDxIzVw
xzI3EmsY9AdFXwvua4cGWuUU7tJkTpCtMlQzutR5HMD2QqFfHqS/FmHDcabxgJNUwA1YKKZMTVOB
119jG1ufBvdWc6BHuHUhacvkqQccXjHgs0XasD1hYS79CU1Yl0VXb1cK/GI8AzO5tBf+MGfQJWZl
RD0SH9t5GGhbOYNjzT8I+PCEnKSGwFzSFkX1X5iOC1F6TGPLSidyZOTd2nLHEinwOthTkGpPePXw
7XBgKOpKsM3JGKwm4oI7HTqYO4Mw0IvSsUd9q/PQxCNKOtbb7SGYVIG9XNLixcrg/QDaO9a3T/GT
jczDDBTzQfMVWxAEWz5IvJDigqo82nOf8dNNnyBLrLTzyfVzzepyVJmOV3VZ6PkerszEVeWRoy1r
bBSOAHN57X8hPo3gzFxyUPW0yBdd4tb3AFSiw6BOG4FXYiik2waebGqjjTL59BsNCugS/ITsWy/1
hSkBAW0MHZynz9ZIgGJ41ATukhTjtrOZE6s5Je63OZFm2DfQ3R4Knv7YfRdOsjtKkA+it0ghFo0p
hGPWQdEOifGz6uIEqD9q0yCsihVxHLPAeLu5D2BIbvuWC84bhDQ+TIBinvsiJWn4YecOOYDuPm99
t5Mc+iSgWVXbQneWUe37KOLeHuv4GHmnZBDcig73QI/7mKxTSB8d6bOFezvsPGj6u6QBxjzepfhW
UGoLr2vN8djuoPdgeHvu688uCAGelDPBFjxgQfbQmM97YxJQRQ25x9H9IrRULwHzXdxCRnLASe/S
DFWdYN7wKY38b7KdNClpdrwKn8kGnQNex7ROaKSU0OoIXzWwcqpCzc0glSr3uHXJY9aqv2N/Cvaw
yG7FRNHHPhrKjC5S6rlwGu7Gpz0Y6ieuizBt0CeCRLFkS+r88sPR2SEMRvg90j6XaFlGwpoe5SkQ
OSPBGv+Qi53V4jNbb8fApGW6BwjYSk0lrhjBShONIiEztl+Sv9DM7Q8PFzkSTegt44lg0zELyikG
XkwSuydKfacJwXy6iiGUtvaGXn4aS1tHcuSaLyAk5oejNJALz/qIk1IVZw04FTE0PsSIw+8bybyo
czxfyQgX3unbZDTBbW+RPtUlWLY7qCEoy8iAWQ2F6OsuAOC/de5fiEx3XV3kA7JjeDfEhesz/Ovb
5huo+sZY+F0fFMCCC/7FbGqEAx/c7gZ3JDLCVzE36VJJP5dILqnDow8sc1fwuBScBAPzCkAwIYWk
pxMu8hFgiOJpCaLABj9iuOfi4mrASpOV2H9vJpdYCu1lctTyGeB9+9cjlgTbuDM4jdKZJMNxZdfv
OGyFE02P7cgul8eNyT4wYe/uNsTa99M0W2URTybIA6qjRTkvTYesm019092xSeZYDgIO+qTyRc/7
hz5ixEx4iowtQ0G3As+Kj5YAjbmE5ZYtJleNmtgceofsKbfLqXDec5ZTBQSZ/UM4iOxKqJb/pvmP
LIsxVFgb8Kxuz7qV9jd5rdxBeXNisFumr5k6WXnkZe9PF4QpdTkzHASH8N5tZ8nqFDloDZaHMeMb
YyLk34b18l5UR9491paWPN0pNc72nNKe0hoGG8+dOHDOSJBmazNuSYQfxd0w4mHScVLbCqFpt7qn
8UT9uzgCI/gSqYjsZWFfftpLKFR9YMvGVHElwnVMq8ltRJeoK3jBbu0dRm08lLu2MH8Dx5Tds6yq
2pEML/QeA08YQlOvcf9rAfjHwB2QlPwQ5biWR6ZIYaZjUkNYVWtt1tN7EOPULb6QgAJ/bUWBQ64W
M7SVO/fpOPHYiyquOyWaUPgoCNAgSHGlGQRbjdPtmPtU4nwgEBx5wmeNHu/IToTXxLBDh4Trnn44
qaPDgL5Z1iIc3UER4ecvyJd30/ie/qH880rldluM2OQV8tTB7q5Bh2aA8IcIW2qdVH0cvI3VJh+Z
fw00s5OgCC3lOMO5D5RCLwiGNaMt0UJ2skg4x2LSXc7pMsLJ1tOBwQHLlBmn7X8CTpiknJj+4XDo
an9+X3mzQ7MZu2B6pLDoA1emBGgcM0XzUayqym40w/gmf1hAXH8SkAdYfS/EWnMjRv+PWPDMp3gF
oDSXhbSzHct7jkLKU2DGqkZjfhhI09sWDb3c5BFat4fjLFQdI6s1CfYUj+YHhPaynP8VtgRFIEfM
dCp5tHeFUn2+y4Xe54AQ9uKyrK+95ZLww+qPyiyJ7c/FyF/IhPQVRRt+bDjvSCiZliTaL2DNKeGk
7C4o2DnqUoi7jvPgnbXLjp9Aed8wsUQ86dxtw9R0JquiA8tomSskPvC3rcJD4/+5sAbtqhhjAI++
QPzESqns30Qw+qxJN3LhaoGiGRKMso6coLSSTqwTIOLxGggtiAf80LfurDoJSiil7RVHhK+LJf7Y
lmm+HMqwpdDsyDOGGM7Ex1YgU6dkkIZV3OVmn7+CPZKvANsASDar4/Kgeues334YMXdGp7cKRBgU
h4dwbR/v1p1A9OqvTm8GXxQFUJdQZ5ChSu94OAreRNgZMZkaagIhxwFLsxxiaEnS4M4QAJdq99n2
lKbofsnUaRRKo369R50gfIiJb0ajHpIRX0OdLGBCLrv+DYgVZqMRGmfsJKWUqGTxPUgi9L8taHgg
1PSdN/URzvJlQteRDbEPuLQeoEC+3Ap/k9doy0EG1yxblSb5OpLxj0/QPSWHe1IDKhfXScepbEKx
jiz1cKA0MkhJG5OS6JrTUlY/8kcOhB088T2qmdHHAakZyZyS9JEjO3NcvVfmrNKtizi9GQYUQxoN
ZRIJPzURbNokL9QJN0mEn1Oh9DHfPMMVeMqcZu/OBQ83FTd650hLrQHxDOTdnuyAKDJkaiVWB6sl
jx+i79TaGw2aAakAvDwIGsQ3+AeAQG9js0dtoXyYEti/Vw1uuvTFa7N0SL7ZuzbFgQJsWOdxM+S9
xfGKAgGpuwtZH/p0UwgCkAPrCAqlkRJ9TKeC2TXfuwDBnKftyFATyIV5q7f7gVamX9mJuZvRt1ob
112ok586eM6GeBLIg40v23NriY+WoDo5ghI8dHC4Udd40NMvqker5gWpsGB/sU0P/hNk5NQ1t1Bp
JM8LDnlseIdxU3k9qC2uF0eAnojAcBJWlapBCDOGGeRA6Zyv49WXYv3/j5Pypo1VNzT38DH/8px3
uMXRYQmVmxsotv7Y0K+sIbaxP8F/LMhn/AHJGYkACOED2Xg/w+t+e3nKSGsSrQbXnlNZYiYCTJTS
Yip74AAFdDeeZs1aPJHJMdFa4In1QUig1xW042qFLu1q8Qau9r64ynFCVhp2aIsXwqv588PX+tKL
m6AGKEInZRAF6Np3/JyJ7Ej33hQak3DEcS9iFiQEe3K6yW5Q5/4zzkuQH8FkJHztqM+dLVrRdH32
X/jxFmBBsv4357eT3hoQC4ts1HwDZP9lRdRk0Qn6ZWHZ3p6xSCUPhYLUyAK1ZlHI3nqNSd1G8jd1
OydrEEARNkr7KKKksOP8Pt9AgA4ALrBPEaPvwfuhBO+lwmKb6horE+uHuRlsY3Man8bz/6PGF0JA
9mMylTugVULGUMD9uO+ugnMbaoSQsPxwIrgR3dkDTAHiu8kb+dsCt+xeuggUw7+MWi9BoVBa9XQK
upxB9HpxHGaz+eTN6enqnl+2/UMzDDfXSTLL9prwev/071zNZ7BrrM98xgrPgo58sysBozvSGmVZ
0EybsLrvxe49mVylzjMEC1hnB4CX4J43e/knQSztmnO4FVNJEu6lBQ+jaOHqTPI0bfS3Ce/T1Mfy
ghq4SGbUQ/aA7wBUprDe7V1zG9QvP/Xj2TJc4VbMVZujQKv/RndDseWs/F8iXDV4LV4Dk+ZXIQXK
AQE1srJQYJA9qpXpNnFTFx1ozNX2V2N7013y6+qjNHldX85oSdiA4carJTi3A3EyM9EpMgSVGKyU
nshYnQPLa5CbUcp19kdci2PS89MJNGX0qB4LhnyAB7uRXxn/mZj6m+r8ysg4HsTv/AiGIB49z0IC
Le8t+gdR+DxyJrspHna0JgWmicXXKqvhVqcgGWizBzcIklbZDjMP2PUEoGutVl5keqC2/Koh/U/D
FPRB2NnFB4Y2A+jnhrio4h/cFKRSsjbTcwWecTsEYy0xlxEHUM9G4s5kZk8C0ZvYEDVVMr2+t+Y+
mBMoJK9sGAjW5DgpNret/As5uA+cTPt+mM/CU45PMbfRChP1ChiAuZokqNnmL2OeH361Rf4BkIeB
guhkEtGYpGe7+KBhwZG8UVgn6WZjMblZU1UPsuSY4QKKxRaI3I5FgqYUMdZcVVTLGWESVysxK6rr
HhDOjn8lJX72PVTmzguZGncf2KvX/h20WO5dKXvSOTIB7HrK6KYUrBmcukKIZGJMg28G+FgB6MMI
hfI/vhdCExGu30VpGU18zttS+kgAxWc6YaEQDSnn/3K16fyoez+a6jB6dZoId9h2L0k0//MsNbvo
prU3NjA5b9xdR+HTyFjNBch21Mgux0zCD0s/KkRpB61U1uBi14TAv8Dx8xBokSepnkF5Nxg2zfEC
W3C3RqNIXBmwpYYEyX0koPbrxb/9lRPAdko2D65DEYTN/hZegM02/l9v/GJiyc4hk66TDK8MKjkk
jiGEkRpeb5WTOUF3IMKqw7NylVo1RuXOAk2Bmh3aHmEaHy88fHItD2Mq8dbs+kY+glOqTUcy1MWN
CbjJn4BPyZlvCeP0KMYByot+vLIfMgdxp2cpujPe9CPpJO1U74T8FeFnI3IFnrx/pHbQLZp5Q+ef
o2Yz3c9rmZVOQ0SoFXbI3o5BT2Xwip/HRJ0UFHVvG0IhBNCSVrBGdQQRjFl3Io+lIzrszMJsBEW8
VHOvztI/ilvS9Wh+OlBDNRvSSqTQen4eaqE6+Y8QBC+yK4F4jDz0fP/bKaUsbkWqa0KMCMNaVngY
HWM5G5wyJrCrywBcSTnS8k5rjl4S5Tk56fxx5HojdrHG5r+TqQWhQ0MHNDndFWamL0yvTerrpJu7
nF0UgFZg+rPdgyvAGF3nYDrUh5r/2m+9AYz4/qSVRVWkhZXVZkP0kWhgpcKnuHjdGduiGKWxzQuG
Wzf5XTd1WRd0J/BGmB0HWw+hTJcVAKhaUOhoVed2xmdDXqdgFKRbj2K3hmyO/fCECfBLEzlxKtVd
JZRnVHAngKQNpQlNf6zNPq0OvjM+jsvbkxM3Z/04h2N822Ro8cShrnE3YSSQS6ZlrLbjcgUia4ZG
ch1Yk/PJ/6mgkZdP0IPq4jQfm3D3HFbsucRMHOSQx/TrwjyUfnuo1dZRokK2pP+feH1MpRbrU137
FQCQYuOGu6YItxaGPwfZuZKINhXeyMKe4rK5HNCRzeQQmSbk31GrtpLXBtlDNWn/JzGIEOu5TImT
e87BPzN02gKKpGLV9VAKoGSfubS/fNlSX68UlmSLcd9IkUo3c8n7opTtFSQbxK6qqr3wI+ik1Uyb
iNLpg2rIV6BTMC5LE6/lB4KCE02TRne8fDBjZN9bOdUHtSOYl73OcBw+R2mg4MhcFr5ZSHKadryH
+RwjArl8QtdW3tKVa/KjDoEkXyHyNN0ImHBmt1xAoyQ5gFZOXp1m+a+Mz041zP6aCBn8DZwoq1vU
LbX4EI4ma3MLk6dXNLmFW913Hx44UT07bU/U4Ar2leXmL4DelUhlYOgs+NDdIl6UhNjHovkc9C03
ciexeJCiIjXHVbL14+h+cFjhjNBI4xWRogySNcdvB7w5qMbpB2+oclr8aA9ecpJ8IoKTdZ09A20K
+lRIzoMXAnWhn1D4/k2P+gqyHoR+1hRex5U3M+wVH6vYqPFjvB4oMhH//a9qVZ+HqHtRcD6QG83Z
Ex2wwwDyHnBUxK9LzO2QZ+J0VSdq9r2vnbDxuE6BwotpiszDwYe++L/7H+8y1KmUlgRwiFNYPemu
g5jR4zlKBuTspIWulMLg5EQjB3WTir9f7pY9gx8mg7RHzy35y7a6lUbXANtayiXlix4cmIUEwmn/
QKzinWCiZL/lJEM3+kFiuzYgFREwaZ18Vs8shtUkkQIbhWRYz+jfK92ee4GMMOdsTRMwhiWKzZxm
SmXDyQcAxDcrU2eHhXMtKOlKU5SfX98IhO1c+5XshBpJARXIjQnmUQiZYFpr909lMy0zbJs3+7H/
M1dP2aPQolUxymcS5u3YElJv3v7x/7PoMFe06ggt6qWD8rVIYGN1cAjkaoxDcviacuvNwNhKapTW
/ul0OWhW6NpGPbevRbnszcYN1YUsCaaQOiI26FJXdWPXaewVZOyOKR/RGUf5xH/+QWCN7+LsQtDG
hFXH1C/5j+PcVBLQrhUjUm/1KBnzeiJUSgp1VhppbYcGdwpzzdy8UDdcT+HEnx9gOWNzSMl4Y5WE
QGgtJczn9LGl/riPtOe9CQJwUEysQKs2g6Q9icN7uckpMElERALLEI2TO4rJwz49ZlDAzSkh8r/h
HShhuDhOenG6EQb6aYSNjnOTu2LP5s52KDwjHZ6jhlIv0VlyZ326mmfaPL/1x5o6mw3sLxZ8LSe6
rJJEyDr6nBW6X+JfaS/oQ2hg2w1E9phXDlsjvZxhiVlKNea+22ahl+FJ63j9iwY9jP8VW+ExurF9
1FjIAXwuYkvGJdlrf+Iv8Y/svIDnK0o6KThc2mY6iLwg9oWxKfVtgm0CCb+/ygZ2vJHNgq3pkX05
8SdWXJ6aqOMuA0Up2HEINDu53QRfS3z2Aw3j16OEfOqZVfCy4hz1X1wl10SsJpkM1xUpdYkEosjd
a5xEoidefAS5AcEjH58AF8nogQWCw1KBtnxxnvSvdz7BIX3JCLucQfVpxIIipHKmNttb2q9QxGLq
Z4u/txyOdaEiGACVI4gAgQx8R1aWPZMriSL1JjF1lW135GlMo4UJ+hM2Le4IpzRrvi0kvJ1DD0CZ
kAv/XPsgpLZ4FF/52L6mkyjdfy+vLs6rYLjXu6lzN8pMK668zJQofpLb+Voe0hbu2f6BrKoU/oxh
WhiBcVpQywPq/6eilKgPCMcpucXDqq2GaGskMBL5wBUtI9UL2/j9SWb4Nhhxqr2toufo9D6agrC5
WVkLKxh4C3wPTY/dxHkbH9qO2mri1SglogQHKHMVMZIOtwAHXjF9Hlq3jBinTufmkkkRVYmPxpdy
nCSREMiEvLIIf6f/OiOlx6OnhZQueZsu3L18zd/rfa0UdwKYNzU0yp/n2dZWKPwc6Wubus6ksfR2
H1J3I5xnbRunPjBGPDIFNSRmsITIaikrvmv0FU/b9LZE5I5iov4Ikk14o7E6dxRdC8n6RGxAzqKX
Caakw3QRVxw7XTBi3oiChr38vtfG0rxfhuWXB29s+iUD78+787+tvoUUctiV55O/fMRwOlqmjR5S
myZNHNmp+cs27WeHXnd23MlIcY6paHU0yQuXvzNG61sNRfoe1p2Af9XZe+UGKVPxPWxwI4TvWtW6
zhqCIqxqrq9Kp8sXlgTBYCjIEFXFVBcUVQZRRt9NsiyXiDT2aKQ8k2+5IAbCkotnSz8W/2W4iC1J
Zyn5C+k9ABi6imH2NVLSQVrp3Dfw1jPlnGjZgK6LFQqWRtooKHPYBm6rqcfW+BP/rooeyFRCGgGK
37H8kuuExXfJiMe5GmPkTxpHFL6THlCItBqMnS09T68bM9uG1Aluyyz40mlY2Jsx1ayOoGEhUFh+
BeMXMV/OtJYgp2XG9W/dQ1wSbnrS42ojch/jmTebYqm+wu0mmK0IJ/O3GdmbNseedMyoc5MfSlb6
m9QYZr9QnZrJJh12okIKQZf2kUb5MUZMjej9i7WeOtIsZ0Lv681cRMjNaVklT2dDJ0hIePYygWKq
8YuR2qtx+cS867Vl+gUYgP3OiaqefD/InXY+01F25HvKI9u9riO6/dJ1NptsDrtk3gOqnRmLMgiR
9z3GZ9qmPDaCAeHnyOzO7VeVpOjt/YVzkW9Jk1uj80mcYSc+Xl2jVeYbyiPkLkFNqc1DOSxXFH6P
as3TxfM+EjPwTvm5OuIAGo+Z3znrHUpTdXu8/BxDD4fHHazag+rro4IWRv8hqYg9pP+aHmfmOZm6
2Qfki7fJGCQTC/zj+bapV3waRa2+a+4nzB3lo1KAvQdxK+WhYYq/uv557mG3Rnmx3J3j5v92e8yt
au2iYbMpks+0G2zSbefIMOKnzmjmF6T2wm5uNlY3EErRYHGuAUun/bfl66U1UwOe1CmUR7HH5tgp
TBxl0pRxM5m39ho0vhX4HIDYvAHXbFoW3DmmrEGzz5I8nGSEQWdLrgpbNXCUFqXYtkB3iOaaEsh4
AcmFw0JuArn8YkWKGWlx9uZVW97DF/Ln0gW/CNu7oEJbXMTKNN6GCJ1k46BEEXTKEzkydpgUcP7V
JUdmVkohcfQckb5ArNF37xZTK2fAZLLhyRkLfcblr+HuTVEUgs6k2J4bTN+iH+ldlTD28Wi6abDo
hbv4gn+xX5h+mMC0f74ayO1V00iHsBQG6g3E8PKJAIjSzdkbit7JpAGY2r5F8gpRJ87T0YSWBfUf
jN2cYWMjhta1//t4/bAaw0fzHMpMMdaipgPKJkzbYl3D816as0Mi1pnqrowHlbv+gm3no76pxr4G
BH6jMnSWQVDe+55Pw2FNw2vFtTRDTlNtiRZMiUlq7Hvbcm51TBgr+CpeHYN6xseOrLraOGyW0j1X
vGDNDd6XqOo5wm52O52jTu574z2R7BhTUeRc2DCfMbu5j0lOKAe6xSothBUJTzhoCkLWkdhX0jGd
M1B+ALnFKwSR6WDyo5G7M/dfLd90ijTtUmESLaOJ1c9ISVRhh1GSbFk7khT5aL3DFQT45Ppdtkoy
wh6+Ic7lsGZlEwgRC1X+pDPhBXiHwiUeU26tBXNguFBi8u8ULcqgU1RkLpaeM/Q3BuO2OVttPJrj
PypW/RI0u/2jJzKD2AD60uNddwQ0jKnf146gz5eNbDq/UBUAlFQDHu3PGc7Vg1ck53pLncw2Ofep
+j8cDtwVIJQrSBGBdVd5lMUH4sY9tLWr1nW24KatOqLRBWGE75Ms8UtAtJIMTkY7p+RK/2vQgW72
+b0LfpLPPQeUtApCRCM5DpQ5maoEMa4symjpvgaMKA9A601Gad6qYo6ogUyABF1W2hRRxi9ehrMK
r9c5X/6YsMf9VOJNUASjZYyCcK9yq0mN/nneEYqOKgjumab6Rs1M/FUkX+2/UeLm6HcYwXqjJjhi
jDq7ZvHczxdMJoL4Fu5TXZ4FpPIiv2CAGHRNQTVLGdQJWTNZrF31+SuEMCw8XGJFPI0hAWrBSMWk
t6BNaItLtfOasIwsJ+zxremNMem6aKfTdX/ga3DHmOOUegTjC2xaG0dKFlTV/1kdajkX/kWqbt/+
DvpZ2sce0vRAWpS9nQyvlCrkZzpX+oLrHP5Da93fEZRrVuOS+dkQdf6n31oWB1aAV+lzMMJ0Ct2C
4s1R2EMxSrCSY1iQiZxX/wsYI0EcH40ewS2kZ492D3htBuW2S2+0pXe2wMNMBb46sk9RXCuCGSNj
dhk47d+bfAR8LwWs6EjQKBrEF/NcuRGZNfUAQa7BqHHtLIav9QRBPp1rhTITiX76kfN6d5zKoAYM
Pt3xfgI+B64wk0+u+hNU3lrqilQHDJT8CY+5+5CVmRZHqbot80TT2a9iiON8R0zk/rvEjrQP5C2q
lHei+aQ9QPpp/T4w4kujHznWRRS4p6Kx9YfczCONT28bgbHuoMw0cJMtn/sMdoBQApAAClzwk8VY
go7Tu8OCMp8eZMciL8xaVr5/94WYlJW4U0uCibxFxw0dzoFGTfsHFX40/mxyYp2P2zPu4pAqwuDW
DxPQtBGvqpQ7S5mn3jEs/XTPjEddSAMbz7BhDW2VUW6U1ch9Hchs9Tcz9XcA1rYEcL0IIOiETGQk
qwzA9tbpl08RnKhY6eA4uN1AcepimBBv1kJyBEb1Yg3d0dFyvhujKA2HV6JFwh8ZochO5EUw8qB0
dsh4w4PE8L/tyKck6a4HXL8LEpu4eu9YmtxY+YvLDhw1yCeT+bwtFKDuaGYfvEDmgxED/+N/NZxr
zsVs2dk2NdSt3sjj4tbRf3Bp8uFEYwbjvst2MTvY7Gwyo+stpgG26mPP3UL6ouMs+UcXV65fwyXX
Sa4oMESf+RyZb6CwmVaa/EYB1EiBp0C6m/6CJUnYIeFNHxMghiUnn8Nuct0teTGSQRqNRBRqfLCC
qfKeRBRCb2nkjqei14FWJH4YF8EBfPggWHpq7aUdpkVDc9e5W3I+U0RSNrIR6JeBFgwLPgW8XyCg
EeO4pDnOnTXUktetMN0XjkVyp1a2Ql2EcnoHHu+LPzGM0HImgkyj+qDGdrM1YajgrBXCqeWvHzmu
zQAuAYFdxAUq9hdRbhacVee5IUemaqWJG7r87nFHqqBH+ZNhp4jQYZu3ZnnX53XioGugkyyrK3xB
vxyrtX4eZe5I1oocVAdqwCTOSlmK2THbHHJCMKRuLuTX1QuvkHov5YkZngAUrF93kG9TfPzq8PAB
rJqJcJ8kyNu+KK7fCJH3PEhqLWR/WWv5WX+fBs8RZRROJOMn12S05OBuxVjtjQp6x8dAWqCCLpdn
ueDtXwuaJL1pLCR9QcrWAh0bxyM6Cddi84Gxd8SOp7fGBTrYOnbUSOQx7IhkgTvcjLyHTicJ/Y+a
epoLRJswVFAqDSz/SQhB7EMswbVfOXY4BnuwS5g9bDD2yJxIAk2LGyRj28lEXfMJXgyWCIlX6aMQ
RZ59v6B2t0zGKGUukfV8cdlmK+VYN+gvuvBN2GFi29LUsqWYQi5S2D1WxPDeeWDCk7nc+W0L7403
2J7HDM82oMEseIyAySLVb3KUqK1vWF4NBNQXAFq0zVI/ZQ6LREhvYL3UesmXXvO7qzstKE0ElNA8
T5NN2v1YoSo2WJv5eJEwa9nlLx+EYhpwyLWbW3sC2OqrVqVdShY5mc+ZOb73HegPzZsUm4tZxywo
+CIS4VuBzQSPhrh3fz5pThiDdjr2m6afFUGCXpBQW/l4EW02UmAPD8EGw4QaOZpLJ34tWpHH/Tmr
okNNGLiQH63FGK/L8jwm4w4GytYhLq5yWivAivYWNIf/gFo8JCKWnXAab2Ld37byySL6lxfcV64c
P04/QhDnYa8X627NRVGwC2MDaYD+z7oNfdO8iSsohTMdSNP8EiUbvu0IPIsXxaNgYUdkLIC2SB0O
g/udcKN364hrzSaCiBNOCb/E4srWaBr/ULXPFO3qTCtZPbxDBRHzlaGGajgh+bdkjKG+VwnoaY5L
yVuDtpvsdrXse7TnaECh/xDJDLlUQUozOWai1IY1p1hiDXLgeE3aIaVm14+Jl57ll/fKepCMVG4U
mvRSjGxN+jmpuU5cXJG+WZ0D8eTmDi+sN/OjT7OhC9AEvP00PRUp8ToYMxuPPf+bXCY33F2v8xG4
uzuMhZ4cMX0SDA1JC76yAIyXzVy+5gCdrUHWfzF1DVp0iTgI6mNrZFSch5V57qSLO9oxIvggKeRR
SnJYD0RxJZaAEXSHPZz5pFcq9TJzf47JdOajcf9Kb5qykDucD/5i8Zmf9ak8uZKTZZVuOeTJ/2WI
HHqtxQ2R7mY1kOzNyMgWcE55PxZFUKwoxrH2WwzkhORVuunEnYph/n8wkflm5ayTj0WFUN0znKui
YtGY8G3dJmwkr++JqFWrzeqbjy/m+6PIk6J+unTk9LiinKNGK8wNgSdVDFG+lXzOGaao+w5vK90N
90zst+Jad4QFN6sA/iXEk8CYp4ErDEPq3anMClNl4/hNhmlkSFSdCxGcx86uz0v+5rG6EdusH1f5
Jl8RZo+drdDwlr4sT8ebDdpaEA55CaceA4vyRV6cYbnaYAIkYwcK7UgzeV2nNF7jtrmBhYZBAg2E
lusVQrFqpDac8Ftj12tzUl6eojWqtaA79ZUp+z0x/3/zxXeG9u6G/OVjoDB1iv0HV8v+pnsLAbzO
K0RZ1awr+OH+d0XfJ5SiJ/WA/1ZB6/vxlqYAD8z94Ixktq52xQKIHhtaFtx3jgC06UN0Czu/67Gz
XJ5AKqTeJuI5qlHyLeL2H8bKvaIXRb3pMoKuk5gx81+TVhf/tTPD7rF9Fax0/+Q1Th3c9/taS26o
dtnvw23cqrl7G1RR7vY5ETQnKZGUzZ0f1IpkKQAL9NZcQ9JqJ8ZGZS0PAjCDK1YV1iFuEmFSuGH2
dNYSjGUCR026eZznroMbM3AF+b0gnelpQwegw0eNessszoxc7zFD9aMDdX+mUIHt90FHSZejMEec
NDWAKAUX0poWcDJO6qRldCDOFXzJXd2AcfqDqIkuTv9UanWXYkuR1YYT81AbeHQ+UFRSxUVVPWmt
m1Uqg6eGgt6yLGA9ZeH0jCcB7HeizSZDE5kqezAiuIh24WlXQs/24IuRVnV90dwRy3gqrMTqydMj
nIwlUea0WUP31X4HMQsJeu04QQ7oCgEEjTAfJ/PhDhGfSoBN492Z2/f5SPYSntYDAuBhm2aUJD3q
CNM1Vma+hz455bOfF4NN5EoLmqu5mDymcETRT/wDzcVMOq5RCJa793L1H0r0gaz8wyrbSAuHJb+o
waHxbPOhCGyH4TNamubONaLoidW1MGhDY0vaZWMM/k5FBjhP1FnE+a0Vt33ajjKxzJXg2EAHzDZa
ADoCOgpKX2zq4LlPZKxAq38ucrgbwEZ/7FIu8zy4RR8xWkoam3hkUAQwt7ZoajIEzjZhZpkne8ml
cYMZPywKoJOxO7B8r8Mf88vfO9Qt/58TqDOcVz39ToPAMFnNfesd/etbPxeEFpa93tbqpVoIKZWK
kGKNiBT5jznV6cHR2wQPha8YMvIMDCuHuoJN5pkJ0dmzaGpaQSB0KbgxAkLV4XoWkPSdfP2YD5ol
SlLrEAslXr4Z3syQkIFzFRelQ11JNwQ3zQ9eeRh2uqasjLNgOBqCwliNivTQzT1+NBF/ocUDO032
s3mYeVehz9Pkz53UU/oFDLavvklHUAu2EPFqQ14bW7YfsQOBlN9dHijNIG+V+fa8yyzt5ceWp5g9
6mgIPP3K8gZ4lzK73KYb2YgI8FPCsNAnXsTzpTI6iVu+fTIJUudbYtdC6YlmGxGRE/UbY6JUKO7D
CH5uHoP7tdEz/inuC3STfn2B3npVbU9vFZ6m5cKcjqvsyeLzo5TZRgCLTER9cUkeB4BWeWyo+AO4
GavV8JOegOdRPBJdrYlyB652rZ3D/bGbYu8LWTTvVhy6+0agto4SCzWbVEE5DPLyW5qJ7o+6Xkrl
Bx267BKFDNwz0fy0Im/Tfm11owpgFC4lYU35tsCLHbmI0ufcOQ+Wyir2VtDGZqCFJC1MBUiwMtI6
aHju9g5Lr13rB2eM9gxV+QJaHtgfzIAAVKJhJCKZfGRrQIopEJj29+JeLJ6eqAMnc6+ieqnuOpVQ
ruKRBuYnFEZtumqohfYuSL7kc+d4JMHDyKNQ42l82tU23x8FsvpIJicEXGYVzDymi454J1j3E8m0
H0oY88Wbyr2vjDnKalwZugB0Wk8ULON+ootudv2xY4Gj8mIPjD48tymYjfkDBLkUr6iuUD5OM8Lg
enxKSrged2O3M2aC9en5JJqOStjqBxRFwdw0UbXwYOm898Rmb/11rVjYlFVltD35P4HETOPp5Kc6
55g2h5OdIDiIkvvcclaLoq2CBWsxf66OECn/cv1IsyPw6Nv1CcTtw4N5b4ACd7aUSpy+xnl1RGKB
anQTRieclUxMEO7JLXCSz5IRds8rHastcq9KTOH8ohIY17lhKV1Sdn3sk18gZ80lkGLGMR6WMHrI
/FfwtY8qvLJCv4J3Cx01cHc59TMta5ssUpd04B4EzKnE4+UHepis0hUcYdhhBq3ISPSiy3jwYm0s
tluKb1Vb3In2H5mU6Q1FlSmDzlnNwoamPnSR1WrvuGVZT2NzIMDpfmoL7rW8DBrZokfSoWWxtjK8
j0V+dLeRsUgVVuC4dvaSI9jDtaHpHgFyxL4ZwJ8w0/9wNAFW68b2OTu3PgPORWIWHCv27hTUqVGg
sp0eBliythQcKriw0WvT9FP/kYStyRh5BjjGf5wV5Di2DNLgRq7o+N8xMC6IwD7xl27Ea/UueoiK
kRGyFZ6Oz8XIlxuXCi9HU+6lsP+kFRhM3Jhs849aFqHvhq5fOjTDrOMLoNP9VqfB5Ghhgv8akGAi
n8WHN/bRC4WXjA8sKNUEWHM7nc+K6UcfHJ3mED7kx8wJbbMxZuQ9l1UEmCRKB8RWL+HZKviDwbvr
BoTJknJhMF7g/iGzfLGhzQeEuRyQ0HekJRyoN2rJrlYAuVU0SbRAUJvg9SIvUDuJ2QlSc8PyZt0g
eKNrCcLFLB7EeCHiQYxbI1j+D2jDDkm/Vjo29R+qawIsaI8EoTZhQ/60kQiprYKEPP38Q/whzKkk
4iSY0I7V9AuNkhyTnvVOJjMNYkoRQn9EpJUVMQHGrH24FK6VBz/u/0CBO4aUTbGbqGSJ2z6q62ul
+DscojspBwAI8831YDCOcDuTiKFIJd/AZNDdcqTVVDWPEsRAe9T5cUad7/sKOLl+wgw4G7r5z2b6
xpC8lnwtyonlMbIgbm/4gPFKaReMVEiHSzndvVssxiug22nhe16mDjhGBerba1bVn+U1wvr+JVoj
ACalccH2k9Q0jrQd4QC0lS+tMsHYA+zrYIS0XfkV3wkDjh76UpmrKx9W2u2Hy2UMy9hBmS0Y6luX
GL9RZ0HjIgPFx9J9te/CA5ir9Ih1r7oBcYFnDPIMUnLZNKdWY2q3qMsCRRRw5iIP1BF8kyBIIB+3
hsnu6CxnvJRBhDdl7o7wo+8ZkIouFqrzbXQVf8uxCxatR0hX+p84f0iJSWfPtoYOqPsmr91sIw2W
psC7mqYnoZt+YjNWDhHmF+9i7HcmEBSkWlk6Kfizzk0NFwaW9hfhkkyUNyjv8cTCvZEwrKNbZrmi
fyVt6aU7CcyN7kDyBHkdgjCHjOfwbHieDWoLLxnNgIySTNbPfNibRk93bpzlZkdbqMU7AplLMLT7
6MBShjRUQXAk9id7PS+AfzE3NJ24fcVzOu0hxmoYL4dxIxb07uwIjiKPSrfhUqeT8uZwgEVz2hJm
scat8YY1Hq4tfLqdd/1XpQ4+JSpWHAipXWnyUojj9KPkBP29/W4EqMvf44rxHomtupJJdfX2jsbc
di4i/6B9OUTUYyjj4/4GYiE7wDxIn5SumvVCMcZGUPZxSs9ZFLRRXMZhsMHICGaaHYwVqpNjhkDG
fmh2Api7P0ifHvPWujFDQ62/NVvrzFxXBzYVXwP1dJpOzZIYax8bZYPpqODOMMTvWqGyn8oBc5qJ
04DoYOjylrLWXlkjm/Ox5w+6SI/n/Xj7mrHS+qoCUOB7eBNwLXrUgQn9KhLCvhEv8OGmdxACBXRH
WFRAS8L29YRmJ2bP8CySXnQhbXXn2LvqozkwAV0+czTbVwdk1AGm9PROKeDbPM1zmcdMBFUEypWO
NFVPRtH1qTxiXU7sCaY4sFHimQCmavLqbOdmcmWdsJpGm+DaH6OUva/lXR9LlxzCTp54VjNXk5eL
3l69F5rNOte4O/26m6nGAp0n2uKRVMf0DCV5YTR//lquZo0utXl90OsVT73tN+5JAPO/yGxyC4ey
iOGAE3xWugPhRAQXXG2qJzIz4UhRuTJYPjJvrMBw+3hmjhDDtuIuNccN3OSauvnn+kKII8tnabbH
/q5BL+/Ns9msEhokd/nEl000mIWMzpEI7sA3vSz6t9zsikuBgUZ8WTSR9yrwoXH4JotxrE2F3eHC
H/BKqLS0YZbUoHjjN4EuZs68Q8zyc9yHGT050g3oCESqq99o28VLM3MfPtHYMDOgJN9aqdrfzxUV
A/OPH0xo8Il1M4iu5uJSBe5luCAn4ei4c4a7G+bAUWYubFHgu7c2A38SJ9R2CaFxyuKoYUxKoNFD
RDB2iAfzc8lmpRuPJMq5IVZFLlDlzZzpKZMQguexTtzGvYxg0hIgwVe+0uEyw6Fl28ZEfICJE9ZG
aQsl8hKPrqAtn4TvS2Rfhi8LJF5AlkjAA/sKaARzEq/4jfrfWGBnikTnXW9vW8W0TtMcPQrmZQD8
Y0adT1qqtpSRjLnTJ1crhFLRjZ6BSR6GAFwaHbS3lSJNcAGBWxiQVD1WjWfyxclX1328J5sHi9X9
P3qqi0GblE//0VQRQ5I7SFt5tLehqlaXFVu58gihT8P+iOMsJv/XKjzJ/VuavasShVtXZu4BCa9E
mcQOCKhsnP7CgLAUBcAvhttXPAE0G964TEPaJ+M2Y/O9Z5wJGG16CsOyj1mnlsByZ4piA6JQOfqZ
SMvQkp/t/CfUY4dZe2CCxXlweOHKbmQTJrPAfYJ6eWQI2dxos2DBgfTfm4LUablgWIdvIgfS508T
QCs7CYcTmRVFks95RqIyge3vrTHhWMpGkZFefVy828625R1p+vt7ZGsAWV6MEE73v8/fqL5Z4VbM
HPYQD/yqByeTH1QVJG0nh1Z4nGZFUcfjPo45O+Ze4y6wo+T67KJkPkExoKyCgtddmyN0lDU3DE8Y
/c1CLSLYLutaPdsRA7MgZELXoJ3qSMMspkCBzgBLrLo4tIL8EYQFWLII/qW0EVwkfaWMg48qU6xw
BdhV6MAVavnMcO+Ng81rGfU0wwZXgny2RCQsEfa+s8qxe1QHBMZJbsocC4FLAwhNBl9YlU2aY92e
sByJHYnFK8CVHVH/VQ2ybwqNR2PUzbX16pRREKjmRLNhrInLaXzc1WjQjgjEnXDF73xgfWu0Fnpk
P/V6ensXqXCpMlJ4QaQfCQ51IyfN/YhU4WmN8BPxn3lqeX57bau/7Qux0kxaF5kOCBzAiHURT2P7
j7fbPHKZ1vp8ryrmqBQ1c6FPgizT5zfRFEXvOh0395QotkMK4+g4r59fDdVcKfWhAWGkQ+/mOuG5
t0hnzSf3e7z2y0lT60gtS5Zbd9Q2nJGVaazpFEsRXxMQYE1yauiuWgRNzKz9wpLReGoTVbWJF7dc
g1F+HCXUgPEbO4Hw3/kLnPV/MfMfloG5ofhDOX/rUYSIGMdEVAzaNicVjhkPPxPautpLT6RVuSxH
4L/S0PQDHW9IuJ90ZMlhk4IMy6ukwtZjs0l0BqRZgpL+hfkPxHslb5m+ep3uiMTMSrBSiVXBsJi8
4NaiV0HyODOoInFLmgAVqBZ8q8BDTItPeHwK7WJ+adJeIygB+gxAAXmDjif4Gnqwzk/p/gYHiHMq
jil7pW5Nmi6NAK4oiSIY2Nx9QTJ6tKhCr3BkOJqtraJqSG1sd5b769vLY6pCzTi4Txr1xJVhcy6k
b9dmlIb8LnCweMTy6qmBweO3DEDw9XFttm7VGonz59uIa9R3pmVJK+/zQQi9AUuTaxJFxxEWUsLO
OIcxK+b8rKjN+0uA7As3S7fV7UJlWVmXhEexVFrFNOdOdlxdyTBYC+snltCranmAsX/1EzelNxDu
+2m7lQN0OLuuEzdyO0/1X6lb3E1umpYVSkYUyxCwdeO44/d6kNPirsRK+LFQVBahc1z108zruPWq
qjmxlLnKbZ2CthvgQqR13oDtQWC9aNeuTRtnCt6ApgKbV+krum9yPwakdZWQkV1zp1zcXYzkJgyj
FpmVX95hwbrrJjpVFANUFwoT+Ir6RbbWdquwSDxMqjHEZzAXsdFDlU8Gm+pJekwhOYaTgsC8KVug
9D3lyPeCdkE+5mj/FDaOXdeWKIpmG8TDAxoXJETy0TAGTl9x+jgApriv6NE2iEaFSmvPc3If+c4I
QKOba1mDx5jn0ITakwb0mcyz0wn5Mfoh/i0W63nTJbIqKNRCa+YEewz05zzG+wKtq/MApLbMxXzN
Y2Xz0QvSgexGfxsHpGpU5EIMJpOWIfraAAwraIpNGuVHslSL45QXedIxKQgYlh9zrv4VTc6BUlfs
/6oYYDtKNJn0nBzgvcUT603cbFRd2CDpt0cyDirWIZ3d8bkvXMcoVX83Nx1qXeCdLG2Ietme7bdw
7hUcW/GZXEQ7oQjhlLCAJqQaycoTp5s/STW1VYIHzOsbed72tH9S5VsJaZISagX3TqrZO8rRpqJi
jOGm/iFeDZ4pGKTtJcVcsrYZ4Iqinlpoz6yWZV63oseKeb12nQA8Sf03XPMrcKr4xlE00NAMZL/i
y2yiWjIws16zGLIIyvscNQGJv/NQxEKLdNrkPmbXNJiVQFfFXYxtPnW8kXlUeU8KwjbCAn+yAYLP
LWRLOB7T13/lpCwdTbBlZZUEMuEdUAcWJUDAcfQOXyOwYli14L2Dicl5YNIjLwmypLIVz/PWiOvO
OZMZz/2i77Zq2jn9vPdo5+ox2dugLUj8i/U3D9T5fB9HLZfPiRT679GLMJ86IQk0K+smtfuOInrr
E9iaisjkTgN2gxd2ddySTEGEhrrA/IMBrLqIjRo7KIWAyjLJeGyX8Vo9NDite7LmmeOqwMJFHdEH
bB0jbf4TC4E3OH9M+LP1pnSvEjHBof5bUmDPpN+nL9JqLI9HRAhbqi2LzgesLpBTrbZ9GZ6jU/bY
ihNETnMCfLHpyAn49sMH3OeoY8xGZMDIda4jFPeZF5BgvzacGlhORuK/24fD8pgSPvtf3O26a80j
USYlZSlKwdm2O3ljhWJtb/2jbXmCjOFgtVvSoCWvNnq7O0sAFBO0RE2CU0JQgrdmSvo3S6emx+9Q
TsqJweZqVLowWvU4shCbwFQ1YA/CLZXtJO6EzZg4A2wxOMXMe6fJTTvFZRfgRImv3QjaZI8EY2Qc
bqSMtaLeWaOiiPT4t+yg+yTykA6lPzz1ZSG5/4efZlitS0dTSNTjFJaeIk/uM8eniDkLSOgP9/EA
2UTP8hvhNbVGjNctFRhjQSY7LVE1/50PtgoAvrCF6p1P8A4dJGPyRATLi9FNOswmvDbpDzDh3lsj
Qd9j2o7KICulfyHroTD72CgJOrU2Tcu0wtjYzKAgfkq7IaOqASerfUVdPP3isWHAIquzOg0TgGM3
zRbGL1GbjzyLbjpKbEuNPzMoZ0pV4cWzS4SdVZnX+Ma3bbq/BNvjDfri7JAUO6wFoc6Jwb3QewuL
E6P8UqEREUdTuwyYbNfeVt9Gmu8E+K4Yc3co6+UnJPSePs7MvnUyJ+DNJ74lo2PhNpxjObDY52CP
0eFwpN8OCajWQOOEddhnsil0VdOG4pJ9H6cXYXdysaoYzBJMLYlE2WS1H2LxuO1DDXyPdJQjUq1E
uP8cg3azlanXhxspzXVAVEh8w1wjKx+b7+lrvkgVYDX87gO54bSXtyCWjYlnbf6cgxqgipAkUvCV
AukrjyENrMY8V6Rx8cMnmttMt6t+ObkazAUm9z9E2gDX0g5aVz0aWIwyhmjOK92tYPrcq941nKqD
GtKEuZE3AKsEDoAUtb0YZSLVyDyT6H7mXbIn0+wV5nIGw0YJ/tipjzZkb6gErp7wjIT99a0KP1Iv
9+wiWJnycTOKucN2V2o6Qke9SbSH/FEl+Y33khrvY2qWMOshhalCEvpG9kUwdstYOOGt+OORpQfT
XdarnEoK8ToAraZC7+u07Qk+ppoqByoDuFFNZRmRJFXzvPUH+2xRcWzW/8xZXnh/9xGTnYtKHF17
r2RKpUlW72iPMVjbP9XHLePJIEsRfIn84arT0l7oN9sWQGLxQpAVMTbR49dCHPWAntdKAzg2n3uJ
2QehJbNZ8GkY0QwuyJUmlyzHKo++yoydQHwC8FORB38wH4IVXfV3VypkAVda5Y6YzXPvaOERGIH0
WyzRFI+7FfR2/z4zN0hB5HFoZl028zS4571CB5fTVod9S0BDa7MffO+aNoYE5K1q8WZbuGjQOeIS
FPqY3Nh45MTU4lwO/QFvStBpQeiPMedn3LbbinqPd5Io7lMrJE8oQwj7WlV3SFg3CpwkfjGIXRRW
Uj5urSX3H2Fi/s65VClu5VGsqY31IYaEOssNgvqyxQg5proACWfQMWpu/Yy5O3pgjnkpojF+F91+
czTHwnqYybGggFIVkizmwx8GWdTFuI3tqa65v474AT8EUcUhlgGNSQZCvCHLvZ/RO+9uCwzdbGB9
zBoMfgKV849Oigyhqd87Ye9DJs5hJB9d+c+u93kH1u+MU36nN4j4yIcii2Bj//Yt2d49iY4xcVHw
EyWjU4A4zufWOn4q7wNHekyLm53T2nFmZbbwtm0i6R9hXN+vpMPG0XfWVj++6cG2h7wGPdes7ig/
hclfoEPH00U1NR0cftZTjV3wNRM8gZftT+PlwVSFLJVgs1rJOU7C6UAeQyqGz03K05pZdCQ57ILh
582/RSe9QSnxYXbVLKdnZ4X7Z6+EZsGTxozy+XnujQehf1Clu1mM4zWXNl0Mp6dK8iqxdQryOTlI
qFKM117ZO6OfXDpJcqVdjusrS1opyK/vlqE8mj2yuXHCafiP4bn7RWUzu0+YV6A4zCsow2RQ7SUr
kuLT97Fcxh3NPFlo669N3WjxpUXK4SWaoQ9eQJ9raY9rkedxqtimHJXKonq3DzMtBhfEWDEqF2KZ
VsF3a58J8/CnAWGZavvzxv+s5szlvbTWKweeP3l+8c0GuRdgxTqA8Y6B3T/DKvserXNrIMabeg4X
l4mm1uHNbOh4v0GtXiNQB7VQR6zAjJ29xU7G5KFvqp80hKSqktXsp7YQXcWiZCA2bNMe7Mz3XdCw
9JgcZBtFRG5J6tkHjaJ2B29X691AsmvRbHyq5NlCgJE6/6tv6EAHbRFcc+VhIa0tBO7TMafwyWFQ
waBr47SKcuE4p4j3SS7JeYfMi1NTOCoIP/h6KamdUrtzR09AIAKDaB8OwLMlxiMOqDZrliVUPLx1
yfB/4XVAhuvT7r4ZVdE5wc07gDgAulQpCJ9LHszggePuzfAzfXYJVzj9HoeeCF9KxUpps0wYnsb/
6yOtoq+iJI2VfOJ4Sp2LUCpb/e6mZCCnEoV+fFQj79wn1nswo7K8K4FtsKq5DHm1N7Iu2Tc1nFZX
Iocu1dnUYWeuvjowU55h449+/raes+qn90TBCTgILaxlrCi5LShDmz+c7MLnUYB3dSLcFhiES8MK
e/H1p3JjfpzrWshtTl+L/GHvJggHFay+nj4nSqMi7lgffNPpkb7vb7eQ0wMIyZkZO+2eK99t7Onm
DQPLw730u/0JOce4ZL6xBS8IKRnAEjwH8eauaq9dfLpz09viRmq7Ycqqrc8eMAU/4CPKZ4tHW7yy
tpRXRFVNBveG3y11suNV6b4KDdqdECrh+A8Wv/6JVA+aLhZBm+bHH+7oGDJuCI4OoggPKpOy6adK
khZPjbIob1UcXOhN29UpfQyBYDH3NO7BnllbEZaJGUW2FwFNTxm3YblluXlbiLw+bL1mVP0h7CAd
hqcTv/3/YjXCTrsfTw5q+1K5QySRk+apG/Aa5Oj95s731jcHP1ZO1lCLJoz2YuUlg+wRpE0aq3Cr
4h5KUQ8rs3O1u6P0PwPryAH9uM4iSxBmlm0n+COdDH48r6A1orbLf/0uXoSM/2An5Ic2MnSOp61D
T2GdBvWKgCsKWo2btiJ2G2Xmzm+T3f92o45WnghnmFc+TuXyREArF7edDi1eupASeMwbJbI08BsF
aTuDlkJl/z/YOMCB7DA02yJ4PuC2DQtErLS4bFXZkZyXiQe5SsIu3I+LWu3mbvsbc/4sEoLTYB/g
0h6cfCp79+S8CM0HdEbzr+rgZjU5V3bVEndbJRE9yrrE9XEtSHaMGf9rvxnMNA555inJ16KtpJee
MYFUUo+Pw9jzDYFWqGXzHz74gWjM0VdtCpayDbRzM1mr871rpc5WdVgQ7w4U0C5a9eeTepeCz6Qz
aKQPTatIRJJnxFDHr+anFVfDz6hmKZIAzMkpgJtNrkt8q8+KvnGO7pJmw1cIn02gl+M5n7KeMue4
4R+JR91S+jP0Axipzg3TKnehd2rfycMnronrooa5rqoaQBOfLhtgvJ0RwhVukGoZIfDUbPTuY2Xw
3me9xsxsg/XaE6pEtBTFj1Q+DmHnvDrgWvjyjlGuw/tvyb4Xp2Q9ZD15D8ozvv9oih6JHyvZ4aiS
M/UsBv6j+/p//sRVt1HdwybHTsbVZW4S7hkIai1D96g0GFMAdDO5FBBc/29/YZV9UUUaUQb2JOjc
0iBo2RUfyzPXFTPVOduqVr3dDQNhGyuj+dRZaHx2N7RSRl2SJS/FzLbErOfXwLRBs2TGCiy3SR3Y
n6xet0NPHb7UpK5gb8dsGnoD+m01Ok5Q1XReYRwBRZjCOYuGlP5Vym/pFWU94d+5uoviJG3TMd12
QFPgQHvOyL5Jm54Zng5nPGFjQuwZ5rx7O/CybcBQMs5Jzv4SYxgIwyF8v5R9chbWR8KS7pe0Cn8S
WsIRmkiKohg21ellQ6JeoF1g5dYj1q15G+FxPrKWum4wM83wrfB4stRSSzdAZQ1aFqJf7QFcNyRB
pv6zp1g0YMafSC7qwf9znFlHsLwC9kqpS9sn+3MQPyAkccZTZkdWlp89XbUhlFvPISQ8CnU0SS9E
jZQ8MWVudesD54Nm5l1W1ukdNwUbKMHt3aA1HkN3eqXIi1man6XFBSWtATpw0Qc7VFAUoNbrMx4z
jZtVzOtGTVCevzMV5qw63tV1xTs1E+mdTE59iscmR+21ZMaWWsJGu/Eb9Tmkp7JWqedNayZDKh/8
fcQ6KShxHLkMtimGLkivQXzFUWWPKavaLn83yeWDppyZhfPk7tpoToN3J1vqmq6noIerpF8jneN6
352Xu7QtHdq3w5uSkiVg447YXUWRKfx6YQWIZPz+Y7ECoRXl3JqYKIwyOpWGWZDcy8OA+2UZL5N2
R/SrYl14rvbD53TvRfoWoWHdE6IA8cko6q1lZZmBj8zg0cV4MwxAwBmG84OpIeHt/FfGFHjbRQzZ
yvxQgD0x1V/+1wpxttL8nRft6UiaIrYwcMAmQed3wOg0FAosc04wJH5hUBQgoyocDo6e2MskEtEk
cOwALtZlDAIEypI6kJJSufYGqWkKpo8o/f9ASETARfSHpgSC/3Yil2OSLGdDp6/jj+LMH8xUnnoj
JLGXURyvDHxdhlJ8m+p7ha4egG53uggW25l+ti7haJ///g9VTQV1pEa/zS7/8mpcQxl8slZ5F+bm
0032+5mlpupHoNifBSK/MfV7kKcR4Exw5Nq9r5QWpky7tMv9kK9A6UqzopiDJZYXQYfXTi1fugM4
A9SSVGnWe2vlB65ompfoZ7SzphkVkb3pcVNTpaBx0uYYPVMJ9v3RhrsrzaT+7SGK4xSevvXczsao
0uUEl+X+9e75eqKuSvOFQ6cMRR7rZ7qWYjo5g+T5xQEqZyW5vFLOIHSig/UMrxdCQX5N/wp6Kih2
lEx1Mjb1vcTiLLLV1ZSM0Y1RXOUS7Wb9zPCEKY8vCUp9C9LFzSlVPqw1KOgLVZRfYtagfF/rNRa/
uWkDnWaaHNrM1KVweReeJ0lmmrfYdORH5HSu/uqcd5UDqEak/xyhJ5mYC2adu7xcobUDdnZWiedp
z6czC8AQx4mJzqugTY0aMP7PQix4cbOMB2uPbvpJq5TsTmOOrhiY8ryY+O1ypEerIFy3GsMaSQ4R
eh1KGAli63qzWQqZewkqBPVJwjENLqOupp6IFjcUPJZVQd8Sof3RtMbX7wk3ryFxdAayrMdIXtEs
Y7Lwv7E7vFUZuOsluFMlysNngcXuxbH7TCV9NaEBl+vg1vXzASWwjSgh7siTPzvWgNx+gE3Iuu9m
izO6r7b2uQLAI/5jBVcAXlaloWD2FDawTle04eDYs0nM78VfPiQ3huTKmCffza82SmMS4EiXsUYu
ukMnVE/lbTPisVOFXiGY10up96aYHiDwuRbCzANOe0zAi++gOnAJfIVeGJqB5KrCVuhszxs6doWF
8CNIK8d+k5U4BpH6Y5si3l8jzO7en1fE/JtwoTAvWLdV1pXcFQOZjK/t9DRABcZ6RwaLZ7kybYtZ
97js+N+bIzaz6VQeLB+os+0CkeLjtTKBKhhDC1T+lUTm9EszzqhjylS/4ad5d0/D+OnZQQS98KjU
/O6UMOa5ozsMzYSyZWyW4+fkw/ETW8I7uY1f89latefoEouyXLHG54N7oH3m8S3FQ6tQR9J82BsA
Iu2Tz+uGRTyK/OaMpHMgvDNV0onBGT1WXcGtH83N+7By4gVTemx7E6/ZfDpKUvmIp0/DDVhXq3vF
8xmq5f7dky2b1GIqoxlfk8F21MgLHMJl0ZPz+0dK0X7sZ57dw8kk7e/QoA7wj0qm9yoJtjfXCmsw
RT7zgbowrYkmw7iJ2HJrD9P9dCX1HsflfE0o/REhc+DPf+xzDph8juNexuGgTSYOHupWZq7LbAyH
g/fSK4lMf7Hrttuj4O6gBrN288WzE4oXVo9WW3pz8qZ4axiDgXHQcbbI/+IuDOM8LAbrTSLzAfWV
fplK4Mv3nQd08pq7q/EB8GXZlTx+yN5W0wqQEnabvy8c8Wv5Nown57ZSDtOfOaFkfDIJxii9grbF
osES6tsuVvjwzpn4B2S0VrdLB6+jPTu8ICIrH1z98geIT3GH4GnKa32pptec5W6cQDqbHMNSc+Tw
Cjxi/lYkoclE+a8webzRMdmLYo0zd+pWothRiekGo4EZegJUm8w0QX0daLNqu+njsknAMtHq6n/Y
IepqRpUVcWL+tkoB5DlljoeakgJWDSmPC4PfQUyPnh6A262l6F0xmU1EFvEiA/iqvpZCQjLUinsq
WqO6wcb+8zvRexvqlxp0FsjOv8LvMz4qoMdtgP5kCsWRI8ObGSaCcaLXIIBb28eXdQ2K21dx+9kz
WVPkylu24Vdf7OQxG5TTd6iB+RPnmh1CN2DBHZ0ee1BeLzkIjsFothI5AQqVmj/96JcxgzyWo6On
J4wB7HMlR3xKfy+J6h0bui5mRgm/Dh8bS/CMDqUqVYXgvG2MPMMk9xRH4NeV4qKcYMlZshaZ3QiN
vcIpKhWrFkhY1MvknbAEaGtnMbTlh9NIaeboLVEZ6TxeeC5PKXFhqEsyZAQxEdoPnsryh6hBlF4t
W5B5mJb8uByAXFc/DTvhY3Zs7eUgbDg7FsHEs3COQp16EYdIHSf47S+KPzPSVG4fQA44A9FPTrkA
fDTdf5f2JB+50qAcflzYIfBCUz9uCsxef5PgZckPn38S2VlU0zKdGzL2GIR2Vl4xsFcsFcJjqBqV
z+i3hzrvf1QPBrHj97UMf6RPGvl0Auux3px+ytMtlmUi0vUWDiQy1k/gzl+uav1vcQRzM4O8R60/
1ULXAyi/cEK2EHvyJshEQ5lNULGXNs4EjE9OftkoOuOGCOjtoOuWLlgdeOGQP4lwY/52TbKUxO8i
fXAbJu7PYGMgRnNFHN3z+t89gl7DzcObGc4+T0vFGfNokzMh/b/wsLi2P9e0ay4hUzJyY3dpfX3D
VamkGjC70fXOm5i2ZLZvDDa2xOqL+wJUns/xQWnfRRYMbLsfkFVbsNe69UlJHjluYZ8acOyIZzZ7
NH9uzbqHBdzT64OKm35HbXOWYn1gVm58bMHD1axO/Xif7X2lQVc3bgyEoaAVQhcdjyewC2mq3pqX
yAytz/Sm0ysiBEinYFGcS0vpbkBv781VN1NrPwT2lTDK93i0IFpCX/rO6F8jkN7qhaLCwcA7caeX
YTAYF3pcPryA1/bLyEnPLR+oEL4hanYlhkIKMlpn6j/EgG3IbPPcRtLiCrjP0Gk2Sbzg9WMU5hzH
va6weM4MX4h+ma8PVYb1a7gHCC+fQFmyX2gJB7p1Xb5TjjS6xcxs9MQdQ0SrljoTrHiMu1BGqPT4
kaAzC48RK5/3CEpChYbQI/dv7/J5skAJrvPRbhuvZSdIe/TvCDO9Aafx9n26axzF0eb3zB+KSLzS
kXlqIBlzMtezc+jgJi6nfHTtLFrGdeylFKNwi+4nDNLBjtIrqZZ4L4PqY92vLqO1IuT/H/5PclE9
7LV+5d99k9hvLdA9zrImrZ8Ruvb0hO82JNfOS+XJYDKC/15WF7xPdFwdEun1+Y9O6WT+FrOHiswC
GhFjlhXgZlDJPFfpd4fwVV9g7cxFqGeQIzrMIw3FVWZqyS2lch4+46ioSCYlbux5VJ9gFKRziUR0
GXzp4hNCHr1p5IOny0i/lGyKjxrA0MkZCwDgewX0tSjjp+b8H/rtaVkZqwPUFVdESgUEuZmAMGLL
SOiZBnfQyfUceiwaQKEQlke6HMFxQ/B/06B/FR23fTz2Mn1FnDLjPxs3qeuPqRt0pF7pJf4Jypin
GvpA3XD7Fi2ulR1Lx36yoggt+mqjFGOoYZhRmw1j8c1IKl72flatwGarWChVKPA9dMh3A1ZvObKb
9WL4HowLvsNdPLQXE7zyatnBQ7Dp4+785o7dEa5yr0saXzysX8+AeTuFRzb/FXp5sEZA0SP+knbu
/NwItHaBJOmTJM6u3l5UyeWU8Fnrpq784gak7/JzsoZrL+z1uQW462MBfSz3qtLEM3KDDOjEO+7x
7uJ8esNz2r/BE/CKZR4kkFGgb3UCAcrWb+yGbYqXjqzd+5+OtWJpTR77aQViRFjZDTO0mwB2dgZ8
7ifIL2E+ZwvjkFtM7adiqhVHh90O/LcQRrpfEiFlF/pPjKCiPZG/4LBVFlmm0cxFQ/f/yK3YhHBy
wIeJs1RGvgIvrvEzdX5OcOM0YDkYKDKDEkBy+HiJ+Dng/UJLcteQMzwfF0jmaP0EeaROIApfyYve
8HMeWYMCIUUlJ1Y2MV7o1qT07v5YA6dJ6FG1Te3x6hsolDHx4j8jwev6lBuOIbB8hXNkEw1jhgJt
qo1Dd5ZGS0agOt+++TxRkAEqoCz6jYGQNd2ZQ8BQlTDvMfuAvattVM+n4Y8EAZyDaK3HI72rrro6
I8XMXwBFVUkriZLXdCEtK8KtN47dzni7gdf2ngd+W2m36+lmvZSkLhqyrmptropb1qCmOfYwSF1e
iUS9vaDaJhOIdwz/gaPpl5q/dSzpg7Edbw/NfNnvtW6/+9T53FXwAIRFhtz4fg9SbmH7KA2MYQtC
MTqKMc4ZgSxELEydwDvujegY+bB8x0kJW0l9lbvXAVw78WnQlXc+deguKrmLgSUupnAoc89G4R6p
10yBRUQLs53av8ODoTKTq3Slo8dXZ5GKmz7KsET6ybG6/LHJTylmDt38fbxJ5LdyHYP/j0XNqVLs
a0I70jXFTmZuciuEcb0es4JyDsTOIF2yOSLGuhT94mqJ5nBgUriVNhxBs1tT/o8RIqtcqFNat+FQ
mPAGa1dIvAc8Th7a/K35l4dYLFMxkmP9Ydjb7d3UGJh6G247MGpXJrRp7hv8hpwdlOxoHu3xFuZ7
qBdbe08pn48xystxxOUvdmi90ztut1ui3x7ZZvCxLj9Uhd0gt/Do+kxq3n1+/Ie5kUMkQab44/+o
1G30TxUjUxTCL7u9pjIlw+UY/aJ6f/PY/KaWMyJ/BBpWBJk/+YCsVnU+mWdLewG4PKIKEQwTv+KC
1tRlv1qBVl9dU3qflfpzcK7W4nZqICphZwMVtVWN2K4/dNJ8zZsonyZFWP3bXsoXuj8UcT6ai4XQ
5SF0EqyWFLH/R6eH1e0B6MODQBqvZmg9oaUu4/h8jv11YPSY32ATWGPiCLRIeT/JcTOf8BirFxtd
ZgF+/DA+hEnQzsIi38PJcNyiPNWNU1+DD+XUHnks5hbJ/AzByss2HSek8OqWcsmOBtdN4aKOMmnL
b0ITffyNcz7w2C5jY4wgsJe+Ryszf1lN2yEnzYf725aV4g2B0mEmIcAB3btxENtRPp0k6u48iTht
myN+H+jxqLNjUmmOoLY2Gsk5m/tPp4UdvEB0SH8iVw72i4y8FWO9trQ6/x56kC/kUeuiy+m3NV/5
4MIqKGlph/HcQR7BRsWlr6kbUq+HOBzYLMsFZ8G6pFB1r4CQjxdWWfZHGpbKBgn0ZM+CBRv3rYZk
AERUHPBHcqWXzapn6YGaX2SV+aPf+3G9BPsnHykQSZwAhHryTxNgZmirSHfPqQihevvhip5CkugF
xa3G/sFHZkGL5hWWBIf13Wsv51rCX9eMpoobqmfF//8pDmXLV4dR+9yzEY25Y2I2A1xIl708Z1a+
cLs6g4ex4jaO2ArkTnJXgW0GHheFHSZCtbEh0ixybHb+ulTa6TQ/WFKuO0ZtF+wqqFQPmssrhTEh
6ByCtXHH23ZJUrSqDhZOwjD5JUuYNwXPA2Z85Ft61l+cWNSasGvjdG9ks1eEACklc0Ki1mcmR2my
QF1iD+nEleIB1Zn+Ys64U+kBAJOQPjqPDkTfCj6VSdkcUJvCvM8L6+ivRILT2bcCXinXBYPF5DeT
RNy7DoU6jmpgIcfNKjaA3XonN8yXJAwsJu3dvTG9SAj75MWBly+IFMz0gw0MOggHRvKiZJ1K38XM
S+VQaQLRV2JUB+wvWL4HYCcdhK2YnI+UHvXlp9ksK7XTjQinTgfMjiUShweRGgtyRooGv3kD46bX
fDkjv6ao+eqfo9QHaInxKiY6LwK5FJ48LBWriZ/mi/00Ko4HIQRm8ZPFaqV29OPXS0jl9KjXdw4o
jaS59lnjOaK+y1Su27AqHX98fNOIK7LGs7QPVSUityi1GKLHpcnq+xrdCguwQkP+ykm4Po7hQ9MS
pngmJmghEFNV+IGSt4WCEv6L/OnpAsCnGs1lgQ4BkCJCsaCmDeH2uALzMyNPLxmAk4brtk3fYl/1
aK0ZusIR56luGTUx4TxmWmXVUWqm+SIsBzOtKMM++LOkPHn8c5PCZUph4tXQmhlMsZZTbnpXkwCO
b3C+M5QCzUgtWubyeQgvRwrtf7y/9TiBBogW4TTSZCL5ToyI4K6bctk6BAJXQwsxFirKimYBwVO+
IIT5WIM0Zou5H917sL1ECq8MK7XuT1KlSFfumVezboDUFDTeKqaZZWHGB/hdBiJqCEdSLABxo6HC
Uwi5Z6Bso8bwCIInqHIOGJGE22nRyj61sVbDjxroYh+sa15qZdl1hd3TMyty6IheNG9uukdm3y92
y8/bfH5icag3/hSdNU4cKMxUzAhKJhw2sjFRqJbOUtQUKsf3gB/YL+4Tk94xZU9s53/TyK4/5vCX
+cw7ajSUdGWqf5C1+Ph/htdflYJjyWu0ndwKPSxlXHZJ+iCaC81d48Vr00c+E6dEne7z7c8XK9WE
w3/02tfYARTPfKmzyHfQUFDUhMDM2OVtEfINMfGmk2rCHNfy4+loGqzsOViWIo4T+upWgtEGwefX
A3VCzBPohRPMmtUz4xcydMSGrIO3I2V2cuno6/gT8AcQYlJeKa5Zrg7mj3AdW5e6mxzPmjppCuXd
w8BIVWKt6Pb245JuVeH95DOHnWJBSGCpuBAvTViOfFPgkUvMHa+dOWGhSBoZnn0iE5n3APh/6sTY
SdzAqGWmSgAWsRxf+ZTpyVcCdNRIq5edRoZliJ2zicRBvvwldzETu0mwDGG06UAH05iHthJIEHUC
vePHju1flAMkqI/wEPZPGtEcdwEfafHx3GXFy5EdqFFgLNI3twJcQtFJAagEKRGt/WCOFAzu5Tct
NF43fC/clYlkJKfeyLjGa05DinBZjZv+pW6GGWxAAgWSMFVRGBgTyx5v4PAKr0iWNqFygyn+z6JI
OdYYZkr/csX/LS8nQmIS4eXv3Kd8UL19pAFt7imoEikjR0rMAMSou9MnrPEbLlofa6dbTxu0s8ig
zSVyryx69/ha7bdcMEBw6Qm0nNWtnJimZymRLRSLu4K4Xj9lOf3kpOaobUOFDRw9psGFPRf8c7GD
P3gdyeTSHIE+er4ppUqJazqjqmhHQ8Aqo4MPae3Y3f3FMAjFzcICAwglgkUtuki+1AaNAkR5duCl
5s5/WYry2nSMM6J1ORcld/Jh4Z0NDTkrxezfJqufiNfx8ncmZ5PYzhuMYT1SmEmVWgBFMaj8UQxK
epucoyaTanJgMKisdR5FCGVa1mUiGU/DaTxQ0qs1W6hW0vYvcSGXI46SomtpT+SnWhJSBEGzYM4C
BYcb4W77Me7ZliSHHjxp7jmVPBDw7cAZXXhw/FhGmxmq7h7DvyJ4O1B2/oEv8yQOXROWvLXemLgY
7ui92MRFEHfoZ6vXsSPKEM+UdYz8T98TlMfyBR1Bc2Mp3BYEpY73a5KW14barcR9dipnkanIaM31
NB8FadaQjpQVNfFVHmabNa7/96jHFmxDncGZBklQkBSaEu1YZVgExYAOgFal/6rzMm1aeWXOv1HA
cpuPZ1lrW3KpIEqHYKDpwSP5qj0M/Tbf8PgIttFs5YtQfrmB7pVQUFuwxaSN1w4SpaxRtvmK1K5z
50LSQXBp1Y8KdbAurMN8T3CTBZon27YwUM7QW346XpzlQ3zDGxoAT16xaBllkDFG52/AkoWqKaXP
w+965BtWr/7KCKkmupOUgH+Xn49CnYq3MATlVJbXyG3+gbLoFcSHo7ytmYQ8zNRRWuTZAsgF/KUO
ED7sZZGT2W90eeT1ErH6Mi4hClJqfSYBBBuh29mrXOR+x66+H/9liNVRmfS0oeOHXZk5pSRdi9p6
kwNMW/V+dvn2Vn8aXm3zTiNLrlmYkRqmUB1vaG6A3cwehVHpAKU3KYiMA9ybs7kVSv3+sqyAB0iV
GF9OQVq2oPCHXBGKK9sKZYz++D36uf4sb6CkXMQnWvCiPXH7ofADZ191wu4gEshUWDRL6wSt6OLG
D1glhKITsFECXsJbmqqqs702IMdTYI5YVj5VdVohIcm5g/t8CaSqTAKkPToj5NzAyjI3SvpavWhT
pT023tvOjY7UBv0hqph1dBu8m3NNytC8o7pZigoF+qcLq4+jDyvAkpeYPiUnl+n/paYti1YzGU58
XwJHa6AZYMc9imCAMYREVpyxtDfyST4nTvIDKVUnvUMISvcSioH+X6KEsI5JiliiU6Xke/IGmumf
7b4i4fWyhJrGGgmJjowgPrT9L1V5t+9IPYYSu42JRy+mHXE/blzwaik3ahMW5veGpd96IGvKvGTv
W6oBo8HmAXyh6V8sAvWc0R3hryIWrGjQRWRrCBlTZ0gRMTJqDY9px4shmz+jAOZlceUuMoI8gXij
TfFiWPLB57lg1/+WXv6MWq7Xe0LbcKyd2t8NPQiMLaNBbBtpbotCxXs9HR6X/iyEIEKt6NJr3aIQ
S70zIpJcDiasqwIR+ZK94izFbqTExLuL8/34s2qTpfpybJUA5P63vd10SFaq0yUtvDZi4hnccmZ3
7rLgq4sFVsK/UQ9l/3suyJvTvS1LbG/dT+nOL3Tly4Fji12LiuUcvTEI4WgBBI7lPyj8ER4BorsF
uBpRG8j3Q/b6FZL4gOQC22PE75OUBPiuSXaBDJgmyEQRaY192JuyCjCH8/NbCqTKG+3VZbxx7vco
i1LuVruzg/OVYQjmL5rKoUgciL12+wCnlsXx2UK4nlMSHuTyqt+K6GH7yh3IF74T2sIGZYeU46gB
uUxNXYeJw9QK96bQLlqJCtbsdZZ3SwtwYYzc2GQ0m27LJjflpv+JCSkM4WvdcWjSoJT/LfLtjtsv
qVMpj2rS7ce4OzqKgxhzS2YtmlYjTvIt7b4QtXs4lAtFq/C4OyCqqNZkbDqbpRpSzd3vGzgZQoam
l458I3smNIfdX22WHS9FWcopAq4ljhSSDAR5RSpGhCbnhRKdZWFeLjRr3iDpPw5ImLxv+L8os+Xd
FWxI8fQ+3eKoxiaiIFqzPbUn8DbkeImhqWTGR65aNR0t3q0k0JTLkOWH2AqztRdCPtdvUD+HD5do
0UpB6+CA7VyN3WDHi4jLj+RZLZk+NC+62xNPASOaQIL2JkjRuPewG0Tu13Qa22cWyZ87T8yKv4DX
+k1vCH2V4C64GHMT7SPUCBg/G4wrE6AIBJzI3a+L2xUa4zek6ZYQCaXDU5VU9AsLqF8khWGkuRzc
Zh23lTZPpGi2gVj37/suNyY9C6lC6Gs4d8oq/sLP+AvwD7cm1FIz8wLXZCDrfTHFEkOKxzky+LLX
eucBUSYUig1jB2lEMOz5x0RxxgLbAnVCS4jCO8y8HtrfdWlmleUUQAAaXoRLkdUW+KxTw/KlzFIv
pzKdQM2sVFcjloSG81gb1vwzeOmvk6999zSexzNdDErY47ohml/qHW9D1wl9QLUp21SmmIxpFXtS
aUCdytt7PsEBdOabFj1rMZ0LqKqVnqDwqLwptw2AvCKtEGeHel7b86CyMzuBVLkuAi7sP9LWCt0S
gH8GnCZRTBrh1RRBvsM4fHjBmyrimYfCinBC9XTo9rwBoyxQrEBg64eK6wR+0Ovat6GIWFbbS9Zk
YPRc/Jb72i++k6J1eGv0icqKYscrdLsWHgfxcizza2UhtVus/A3YDnlOVqtI0nLISHxZxp7kUEK2
3XHhw4EeDKbx7+7OPzwbOpmsX0YFooGCV4di4y8EPCpUGJCDpXisSJjUUUnLmSHUZSQW9F5Mctu6
4uqk+2XE2hUj032LMzCpwJvW89+5omeAViM/0Tm+iqXvP8VBInhBE1GtXt9EijBdKgikQULX7wJJ
/nHzcADhyXVgGGo2bG0I/JwWG1qsJqYWV7mfAaQ107R9PCrJRZaO+48RqdL6FdkvCDMqJYnEvhof
qGn5XuCHnhuxqN8SirrsMeOxxtB1cBTUjoOpuXijXXUONHrF5FpBrToV8nodiEHBQoAboWIbWHvz
Rw6Iavbg8yEoaijxcGqCspsnwby0S38SZTxOnx77yV9YgtTZB2c2rXMlxuV9ikYHDc+deYRfpOCu
nvNMva3/1pGFSs3mq7N9LukaN0tJP1RlMEeQaYVxtmk5V8QDuxyN3QgfEfgHrNpI/D8TfkadNQaW
i7vXJ4D4YM6zWNxXJbV9xpm3JuxRxeTCXjWOmWKG7Skw2C+CvuRnnvYuONHCDsvsfdsTmgM+YUlO
0ortCNBJvceiajPwtvErL6dxEz8w7azGRKvCI236AW2FhqdU3QyEjk9T3ovOYx77TH1W6JDsMVrV
Zspx7M+9A4dUjZ3jgd8rpegTnXj1/PZQKAOkkMWTpjz9+rPXb0nIcDwb9vAoj01fSuceNmri2M9I
nSIgv61SIrfF9Qos9lJMIeWDP6PwyvvBSTP5UBo0i3vux2ygVbeqxSLEnJYkVkvM9VoVQfqTvDD2
4p63b/+gwjQvbY40yxSgZ4STp29obw8FYmIbwlLrwRonZjn2qsBv3aMZK2BD/nTUnKC65TKGgXk7
6WNZYL5o0mfQglwYrsGYpfkmthqAnrO0Me30H1j+j/sU1n4Qft1Mk2qksDe5Gw4YntrhkDSb01Oc
vuai1ECR75dxBa2jHKpoRNZU3oXlnOhWhUhK+ztQLprae5eVVGGzMzOCTMwYYcm76L6SB6MvoWLn
pv4wYj1cukbzmKUkVZxktCj9cbQWjJXWP0/RuttTMihRaYtH91iweTigGRxs+E5qasTNIBtbCupS
AGqvjtE6IjOEwTXMWTIKH1b+x7QjRBaIDu7UUMqlJjBk7ikO0FuXqkxCx08dAKY5QXX8fi8Cupfa
HorDu2umsAMKerDcjCsfNvdTVSZ72uxUy1/pyGGDVk8+infF6LkI596och+bwkcPUU//r/kU2KQY
zM4WeN+bBvEXyxNJ10wuh7/biLFLqz681/gigw8R+7mDEpQcnD1oh7PS50qcI/WUJu3XSeUV0E5h
tySfqoJwJSi+gjoT/9McV0MePAy/oUm62EqZH5kR1i3c0AS5alerXqXQoCoeMzMOSsxPn+CpabuB
/QFNRrhJA8zejsBZOBmmfVJEKvKqfwD/Aby6W7SlBwbiIf7ygJM2rSVQoD/Q8nQEq3raj7RiaX/G
lb436zK3WhwnOlI1n7D/Ge42krtSRtI3/4SeXIQ28OUObz+0DUKxHMjCEn/IpB8/X81kAJL+zx0u
1L9BS+f3ta0cG52ibttR4F0eXwxPSWdpMyVETxYXS6vxE+ZCfjJxeyU/+wHT+9zV3NlrxsUBK2h9
/z3iRxZ4gbLqlrw/vyL2j3qRV54g9fmVKNBP8ZVWb6XKoI7LMUXGL9fZJjl7nPy4L2cShxpQ/rVF
gJ/8WpAguR3BYQuqJkPHrFs6HQ5yx8SqRmTy39OCdKLsdzHbe7u1FnWBrAHJGXF1wFaSTiB8kQYO
MRsx3U0QGPQKBn7L3Nhlrkg1Pzs80rx/yss3Ss0MOT+ZC5dy2gMIKVwXc5V4IwqA16g238KgANs1
xasu6PCTDrNJUDYaJxVWw3Md1jVQI2RlYOEB9bkjELsYdDGMgb38XZjyod/nZ/dwYqmcTAB+4Xec
Nvk1MwHs3hK2706a7wfn8I1HgEA424GU4VtYJe6pTSMZEC74Ri5gCBdjveaJ+xmsUBP+s1hw2gRP
3O+IshUfCGLP0QgvjaFx+ZaM2T4XOT2L532HJPQQmRpzUnGo4eSSRiXsg+dOSm5pxH4TvewhE9y+
XX6J7XC/DtRtQvQJaJDmKbg25hO8nd2DeU1NPz8SWpR6CUAU5Uf9twZVBOlpGEnPRFsiOxuCS/li
kHKu0EZ4qQPeg1jBdIWIejqgUjhstFWZ77IqcMizLXPsDRd8ku7ZXcZ8jKv3YbvtrevaDt7mMeWd
vk753RzmN6JwLW8RZ1SeMaEJU0Xzooh/gAEkE5brlHvvEZ/N70yl33LbXazaM4X6kOP2HWqzNmZl
dFPPAV6YRungtrgBs0EE3P5OgsVspe2Hyk7nji21giafL6L8uE4rkFU1xkfXKu5/ET/oPPPnr9nY
ZJVLLLb3+/1WWT9XTyLxA0lwqBcZc0JZ2ooizJ2ENLqqAGFTtKf073IvfKshLvLAqYD6XV3rDd98
LvgNHjoY5D0ytqOW2+6J3M7LnD0DXb1uHvN5O3ZRSP6lLpZE83YGtT8UG+SWPs6V2rIa0AjJb6nO
1WGhRHLkKH+0trnX4ZNkttn0JXwxcRwxLEJFJC8NtsqUx1/9JSpTZGXu06sEgFGmixZPOL3AuIl7
nIzf7FaC3ZzZRoTTQHj3XoGM0esGaO9apFNk/i4fdTUJzIgdDiW3m2ot59TH21d0SLhJATFqyMGT
S7GAEZyB010HPK/TeaL0u5lHpGqOx0W2EKQliagQWJZy8eNo3OeykYOAt/hchA0vq1i49h9nYnX+
7fqlsG/k/ydtEyMlytGCCyWAlJOLZa5oFzzOY8E02jgyYfONje/Ik796kdqdDmVDYgybhwD4F5NR
Sk9Ko1fTIExRe8pw0DJz7vcyNlPNzPLR8mIEdWRZSpAhy4YfY768CFMeNa3JbE4dRh7fsoMiASQD
Mo/dsXSqWQvvuNERyLsKQVvPyr5hAsUwo24zS29FNcpDyncz6UDgjmLzz2NJSwytwJEuUCSy5kyQ
3M+6H0uVmmF+4w2kePImmlVwQnfQguCeJ91xHg221ZlXSyJVDFCfkjaiEvA22rUiZcMapjq25kw+
z+mGL1sjy9yxIfoWENqcsxr/ma1rE7nCGZZ3fYD4aYE8FUtI81g/vXXkPdXXGeYg3dl5P2IEXmGA
WKSpQwZ80bq0djtz4Sw2WbrP+hCmAXWPwd3Yqe7kk4GVnNa/Z55n8hQD13MmpeYBcdaiStLONByZ
08Z5K5C1IgMAFxRm6H/OH0HVXQnkjIy2Y4A0mPUfzz3ivS7kWxZq6oV4UU5RpPWdRC1sQfvAoZad
+FRmMc1mEq1FneCbafZs9a78G5GM2gBTxZ6XVzjvZ2j+lqDusDzF+VuaSNveGtX+tJI7poXt8VOu
ee9aqy4FGB14TP8YkAZEniYwmbLimGi2+tFE5Q8H0KIf1gGaqrxJh7zdujmmtiTVsEjmTxzxGjwc
BUetJAqqSi/yxWc+AiBj3+Io/GQoVZjc9v9vnSu2BuRhR+0SZEn6gR+CTrLTu+Q4YwdRthpa+yWH
i8BuKYtTLMTKrQXt4PYPAO/TIIIO5YdHNlbZpUsUpiTl706W7yfdzumHvwyjSr4TxqbUCUvmv/06
ckzVB4UG4JoyfxGGIPCZS3YtXRbpb/2SVLtLWjon+HvW7qaIVLMdM8cnLPa2Wz6izFz81S2wC2Aq
mtazJoai2nhJbdu8Wvl84UvF21qEjFiTFVYA8/mju3vKBgqCD+YOCV0l3QtPhety3QYyCO/WKbjJ
2INWAQFEAkLxTYWGpqg9kTufTQQXw+/nxswwamZRbMhdAumXYW0BkYJy5KqFBCDUSx3kmOG3piFu
cpMhzjHuaHl+ObDVzi8GL2QQVn1+q/llXkPzgI3sJlGXZvkXCdDYVBNxDi2/V385tkn1K4wtpRhQ
jxdjQWdRoJICFPTvNaBnlNylpEpSL9i7AFCM6p4Tzcppj47hMiyT53QR9I0sPPNPV+4IVD0wevmH
rri/O6W5u5x3ayNwExGstXzSZSVFEhlJShsI2ZaAKQMqDGr1Ka90PxUmeUYOJZq8ombu7PQh/rZw
mzOmrK1FR6AoOb3nYHohFBUV/Wf4RaJzXuCUZYufu14Kn3HEYdFydLlJwCELitIcAhUkr8thY4zU
u2IR1kjWZB0nrM3UAV7lEdJmuf4D/STQ1A2Lx5TjHiXVLYDsAQHzNz1aksTFL+svc4FDf6B4Tqda
x1EqDarWz54Z5akxDTNlcQvnZEwDjuyIpv7D0ksmzGkssfClCmwMyzJHOfmKilTA8O8HpFOzkBcz
TLHQqHIiBBMcpnFSFpJozVsUFMPWONQAj8X0y0pqBx+6R05zaIRv4Yc4R4pi5gQsRs/SWh1EKk4+
NVmSeuMyFW1FZ95h31eNNnAyAaW9G3PbtHV6UkZI+InM8tDN9KTsWXDnWy2CD8cOIHalyRJhMA4a
kJuyL7k4h0K8VrG5b4j1ErmYmClmrHOjoENNIvh0Co1gqkdQNZ/SPPpnJ/tvdKHJxNL+YKK7wrWL
vHu5jeZ0xxmUUm93LlSuikGD9KtGRM9lY5COfY3eq34obiAUBqQqMfw19+aftcCMGaC8H+oELiSu
cajnNoL4UfqShflsYtzoc0m/GDM3lH48XZDw0VKYQf4ASeBNr4+OpNghI4osDNXvSB9ST64lugcm
PMgcDOHvi2VCKJLTIPZTbXdGSbh1nMTEBlWnAIZUIf5KT+yIcpVnCPcRADmEUyq6NchqID9sWDM7
+3Sw/N50vqqUgJXKEsGmILP2S5aSiAN2LHA7TIGPNHh3xyklCP1NkKDF31Q040WI8xDNj2kFYUhx
RUVKbImgnK4AnBetoUMF9iUrn6QCiI8Zr3bIwbrlec0he7+cgfsbXE7HbcsQI8GXM0J7UiZFmA5x
Wj9bKD8238W9EpEvQMJQAoqTsTtIu2566W23k34pzZzQ2xpWf09YHrKvJXUqbTAzVLqv/tMO7/1o
ut7UKvzxY5etarAwA+9W7vxlf2oQZlIIuxQQP26Y8KmrADEIK245LZf4eXHVbY1BhEhxR78xN4JN
Nf1KeQqc6pE6TnY4qZQpx2qPoAT45cUYZIlbTmT3hzF0yImuxS3wnoc9Q4aGhv6Yptju4OohX3eP
vqg0jPJ7mpTOqSHXLOp5NRBGcjenR2OI/gK/Gj+YLfUdaTxlyiGnfznUaSLTqxWHLEj+dML+Oih5
TYelPhZOYox2RTKqiFmugL1r1S0gYzSws792oy+76SKyQIWFrHq1Jmyx3nofm697H4NlBtcWg2eR
5jzVDpPZmna94uZeogEn6B76IRDy9sncdJ6DeAJqe4Qoj+jsx+mldH9fJLHOZwqEHQQisR4XUF9h
subzzYBPRVNRN2Qb49vKlLvF/UJrvhEO/czW96U1ZxDw+bDVwrDmE57jXTmcEjq1CQshLJcGbnGt
gpm/hnPT/CLj9kO85yzi++l2CY7kFd6TD5IcsKXjsaByepIUkf/+ZbVTb0KPA3rXCYxe62+8lI2X
3ol0fh2rxHjFaNjJDJCk/bnbbYe09j+Me8XnCo6FNb2fVVGw6Ls6sE726nTxRmYtzDHPDO5yDxxR
LbAD8N/wwck99pk3RdRIXkDMA/Pn+AZohi9Mqe9Tbw805SZkP227T4IzM7sr8x8GLzRTqXZhOHQD
+N7KMiqCLvkj/CRm0GSYb+BU7pk3vaXc1Q5QcTvwewRzI4PeX4K6ol9KaB9goz2R6s3EDcWEj8qB
Kawc0G8QPGvFMnfU3NCla93ZZ2FNzvS1oklUdSzpktYaOFc+FqxReOiDSjz8VCtn5aXYi10oQNgw
gDjpEoKubQ5/wnCXoM7nxkxpCkMOC88RcUGT5AQo3/qMXSHNYPcS5E5/jI+t21I9FunlqLgBVoUC
EgVomM2sD1haoN4i8+zooTeuy2BeeO8ZQUFRibGn6BohB1MWCjNxlrKLRF4kukhjEu5QxFZurSVv
iNG/SqG8u1tVO0houfxq4JCsCs0NzsSbgnArodicP+1hRAAp+Gp3+XprJDfNuP+B3kKnomtxg/6I
112RFka90thvGyJUoyANA++v2331ehrbjD7j8F3af8l4ZIYLpFh0yyJPxYq2IW237s1OP5O4OUVa
GfnQGXjWreeyefLLzye4HdfduNgE3uabCdrpATk7eDzxMQY78QPjhlYywulqrj1VYIjkCywyKKpY
DEmQsiLyFpH/pa8dYWxsQQZZ1K9snp6i2+HKdGd6i3bx3PKbUGh/2jkB9MxU8xXsw82ZbCxAyWD2
gfFoxyazzKAXVHEg+3G4zPSP2iXBE3iaxa/dgLNWiZP5EMqpdSfHi5JLAqhFNkH6I/8VKf5gs8cU
00uarEpU2CdrcI2EsoHuaKE/QHepHt4Mc/HJ/LiYxL4m+G0AvE+55r9xAg7DnHq70E3HRxH5KBm7
geJdIQcOOdRydrIdjxYsA5zHAlyfuPoHnF1qGYzpfzVkfus2TC6jD7yQFz0DAbZ0Wh/0V7xk9yRY
yFp91llLXZg7IurVUkVAFV0eUMUVo+Ox7wKvURT4clvtQ2cCP7jTSUH+On4Rv2WzdjFeP5cDYKlI
IERx2xaaUVC2jZXtuwJl1GpXpxaaUvL+ZP5sbB2hf+Quk606hy06f0GlTFVlfpkSmpynavYL5aV+
NsvO3ZsiHetNXTkAcD4LQiMn+RDzJWU0laDYKj23X+JtLoWvUsmCNIVH/HUxgselOiXCA7Srz7hH
pyWveKcGa9BQ/WTH1aeQwutH4vCLBVX2IgzNoCoSaZHu19uzES8gspY1bO0+SXwuipOPLUmgSYRA
mSd80eXntCTC4S5UhQ0D/Qdgg+0mLx3HZ+u63c4L+dL/cn3Mhl/SAvXjWZjc0q09cs0sBWbLNLni
nITFnqf7HNyyO3EcCfizuANupB1eWTdhGC0/jA4YRwZyjQjIfhu48YMmeTdK33eVy0CcZt/M/ja6
4A050lVqJdiVvvaLEYpbFpDzX2qdIltg31dqyHyIyEEwiXW76Tj7gklgJYHsbIpDc9fgGfd9KkpJ
sFGriAKYW+xZlKX+v0kGQpDzknsk7RW8jpPkqFCDF49IqzWvEC6CcGDyrj6QXD3tI9+t5xRTGkbC
vm0hIe2XypIKudD715Dqy03S0uXGFjlQU7wsX1YkMnIpBlwJwQi35GhcUiHN/6ajhn8AxSgcuLnf
/xhEnnZRjZj8cx+WZcHxjIRxpIgzayhRlAQsI9YalHsUQg8X6N+9WQX4Xd73TQaVCQNb1UpOEEgP
omOkPAZuYDZX4kIaVi1KsTc70ga/vJQiOVsVQH/2iNSaYwxKKfDkkMEo7i/3senrNXjOlH+0+zR6
oQEfRdLKlIeTSAaUzCjMF7pHWE+amzUFXPki7zTe0zsv7mWlzsBka/7LlaJs7NSdgE2j+0jsCctj
ltFhpZ3nK0GFdVTxrJ+42gGedTtqS6AZHPyhtvX16LgXLmfyJHUSdOt/T67UZvMIT5ayD6o1OdEm
bsm5FdZYdQ+K2fzZvNexcA/PbT/L2RGri3vhn9dDXbAKNUW/zz4hXRS8z5BhDn+hIfk28Tbmef3i
ZaToFNroLUo6U2X5u4jrIqIcz47MdEnXIhTnK3XkqlvMo0ZPFls3QoSgjxYX4CURsqiLoH4/sUe3
y8DLFs0sakLj19yJ7QMsSePxecntPDkvCshGZrLmyTg7pU6M612YuLv1ixxpTw1jzwvO2bwr/Kb+
mGEJjewR/9sKJxB1prmwa+6zyJKE6mstqMNhWSyiKL+qb4r8+s9+6sY5TRD19oE6qRA2INmPVrXI
RY36NA1ag3utvt2HfkavwfZiFioQ2Cpa77h03+95UVeA/E2GfBZXwcOHYHCEnLURhf3DA8QgKyLT
3V6LnNE+vrS8PGYIv/AGtsZCW/P5bHT6Mowa6fsazLYkRe2b2B3AOuCPIsfnBWXDsKV+x8qWffHd
e9mS+OJAf//uCIjVoIq0PfCWDwDV9Vhdct0A793YVej24CRPwQ77lzxthRxfnzoMyOAoGPAWtU5U
0LLrV4NfOq7edQIPhPBx/nohJ6yFradFcbR1B+WdKkJOTjWe0KsNQ+0yiV02LVIsTuB55t1KGGxO
OhNpDa44rfJNwuGJSE+1Z+h8evVnsTUSyOQjGf0kIVAI0k3Q23aJ6lwHxN91TGL/J1pyEki0KzQ1
WS4EeSXrE1ccinsP+h03OVQvr8KHTXkbl/84BXQ4q+NI9WUMiEwfnluF7T3ws363RvfbZYcowsRo
SEXsSv5H/W0dKr38RjGafKGg1V8zyEzaS3ZfT+TgEXixFgofMH7Ko/rE9n21fpJwDzHN5VW37uJu
fLDH3FkP6X//WsIFR0vvIrNHmNa7Wg70yDfhfQuesLu3tWvoGO//Yfs78OaQH5zl/esInop6NOBt
ZHmSl//8u6imPwPfQuA5Gs6MilNijop6at7ReYFdHqP0age0/RZmgVz+1vNKwq7xx9D+owkgSkmx
ScOSXaPcLhz0tA8WreLIM3s23zrrRIiUUhNhMYjjmyKM0QDrqbED6CXIKprUllBh+mvS/B3v4h3b
kgQjQN8C9b5KMshTZpMBjALGadOb4QN0JUF1RySZ8aPDxUPNbNs3Ma8qo3fgcg9uEDVJxvvJ/y+e
qXofZmqFNpwO+mahTKhJMzQhHE3/5v3ts8rqUZdwI5zhQZ9XDZyObkbeATCtXq6c0AYGtFgsgUIB
OaPTwX1EHvGkS70zTaYUpSv4Jmt97NdTkmX+dRDJ8HSzoVLWj/Xe9R4Kb4UE1jXpB07+rYz330DV
KcmEiMGSjsY3rrDEOhbYqL+1MrGXrDGDvhneC6FJm9FNsp0NJo3cOKzKJSqu/qAa0gzyB3F505GA
CtqdeRVWVb24wAx4CJgotMwxbZC/GMB0DEGWWuLo+soJEottonuab6L66oMZmXshpFaBJWLmCjzE
1/6KAYS2GR9I0JDVtnQUhJk532LnC3+6SDjJ1blRZ2ph2BN5PFAOpbkpzKM5/vyH3WE/9p2RC1RN
4JK5qjvs4sA8VI7DFWcH4Gmmc8KlBMrDn6xwdgCItYRKLwo473vgSoyfii0+OZc7sWy+7ZuydJ5x
er9k+EW9NR7KMaruRC9i/1/V0N6RpRf4q1D6EUSHCvJS/mBrfYHT9OGqCcQJqAq5i25VKooFKHkC
R3mzQ3E/wX5SCKY/rTgyLanpCqICQRWAApWxh1RkKCRSzMflAhcWtQzKsfKCpxk58NDegys6TVut
wsMP1R92JGlN2tWprH5GsDcYA+mcYCQn6jaUFZ30dicGZGdNR022e1Nq2KHyCXConTD9uuuhcr5U
ITQglqsVADAZkVkcN60DumilgkdkYiS8kd2trpfzVCyqBHSrHrGbNj6XamndKHoDUig3nH0q5Csx
z+/foJlB6PPuFAgD4UX530+hpMMAB8LU+ZZTdhYKsGINZFEGJPS3qZ+HDFd2iA73B97w3QgIeIUJ
jBDWbn1qhiJeuw8pXZfs2BlVCNotGbczGRWMyYGC13gqcdlh0rUkE2E6jVSI65STmNmacRhOV6Iz
l8GeoQfmJ7CD2NUwemmvppJtizP+Rp3ZhQS3/+8uVkjD8r5c6JTwhx/wkLZ2zYHeRcm9z02BTTBz
X8qZKjv6oAwqCxFba+NeiwjDV8IbdP4KRoLH/Rclb6HFveztP4sYmWzLbO/TxrWUL//T4g+gb6h/
yrrKc07K796v+yIE495f2S2OZmvr5KQ6cxOwt3FTVjmr/8O4fZ0BjtieXNbYS5u0gor2+UZtfgps
zZj97IaFllJSHIaPwXu8gfLfjqZ2Ch75T8/t9LlwHXqPAlxaZpZLh2n5uOTHwNMrufNhNSyWcQrQ
AEWJFAak0Yqu5Zg3pmL+8bnEaFUPOV5UoCoB7YzLcRWBelrVXSKywL4C7r1E1i6MvZiH9vExE8y6
JDbk5VDTEA8UBTO5Jmz1qslPslwazUltpcFCGSemZB7g0YCIW3Y92SQwvlMreoG23NTrjwCwDVn1
POmpl4mSrefyBut59w7zKmDCLBf3WAwWUssuSqUingFGgTfywXEht0Ze2Z+CoOv7jC5iUArKKajV
4OaK8SPYmGISEh+huqSwQ9GUTbjRQK8eL8/Dnz5lGo4kUFG6KttjRoN3visibpWFGBhMrY36WyhS
VMaohlUEL2ATXQTWxzYdzIIn5WP+yvjlqf+p+3MjjMNmvgm8Qe3X5+MxuTOsRVwj4RkdgJOGZEnN
UBeaipbeI53j+naP3Ae+Kacr7K+iorhSBWygN9ii3DSlwTD/4sGkMybeAkw68Y5Uw1f+GyMXHFqv
KLTlQABIMEUMC7E4XYsKLzyT2Q/bo4rEeUNS8UTs7Y1daNga+9LoI8Aal9C2c+WfAog2cNiegwi9
xMNOM7Jnj6xh0yoXVygB39rNbAUxnrEyyDTV1yEq0gdpgszZ2h0duFH2jyY6RKSBUyoAHMe4pABn
MDrfjWsSCRwOSpGd8/PS4dPddNzDunm853IqQkNoETiCYAkmoRQlhIwWHkHVwpQVkQGZ6rUSryVF
mQ0VyaJ2RSEaI72OLEJe9wZliNBVHC7J84TYvxbZ4ROBovFssUVJ6ff+iRqf35ahjIBAEgYRhj4J
njQAWaI2tm+v++RyE0UcOxbIqVN8MZA+gSHh8IZFlTxhbbUhA3cujDQgOeHscedkXy/7DR4QjiVL
YforOTG0xvVuRmcjfjAZhAHSoMeBsxUv8uVrWS/bNZLsdbXuY3vIbpFMyk+Ynkb+UvkZN/N5+TmE
o+t6QwWx8yaOeZhZln/5c39u4NuMq/AlxL2vnxf/oKA3Q7XC/rp77zw1bxrs6Z+MKHAQq32fnl/Z
9mqp9oRLYUskqhOHZbgwo9uXKUogBk6wr00F78NuQWUASeDD6OrZRHL5+NbYK9e63fG5NyJXJkKs
n8rY9C90Jtcn2xA7zCbVLxudQOwiqSTiuAXBrLyuvWT67kaOZm74fw0h4M4tzQ1Fn7OiHEr6eNcF
wQSlGsIsdDW3q1EYf0B/5wWJJ847GEE3l92Izg4k7LiDcrYSG9tMlkyzAt8Lg2O519Dri5hk0s+Y
8y2Wsfv6l1Cur0WrOiYsQy13Pkqy1P1WpLKlSDDGq93T8E9dWPEb+j6O1XgszL7xaJX4VBkClHF+
AN+2aqJLvhZdt+ayTwyAnOM9kkSaQ/tcO7V8aQ02ETAAno+OVZ1kiB7PioMklTSKHncIm5EtKdCA
rX3Hun3uA2cHciZAYnLmA0NgIESTakeatrQZDvXf2FNv/7K455l8ov7mV4EMO4EFWp4QZ2XsvfZi
bP6qmdtBywuNdeNKLyXV0pK5c/3d1EpdelQnbQao7eqQQDqrb4LpmKiPrt5c12I0YJDfylcbS2lW
BakD19UtsuU+qxeUB3WliGXCXpp9znpJzDy4tHe3Vhbsh+fcw5SeCPP5A+UPESLTjshbu+QOcizn
2/vK2rLiRd8bQsPilFaWWL/7Zl8EtnUnWOoT3l/0HcF/ckx/TqEiKIf9Z89V9e5QBj266kRKYHio
I/IbUXOBfGCwTseYjh5gCuDvoS+XHrsOoUoVooBgokMxti6T5I6eWMtpIbgDHKZp5PanTPBYHK8n
dRzkCCxBVJFRdKZP9zLf0K6ah58WdkLiehsnufmHlE6QhDwD48OzEVC2fc5J5KisEAteVk2o6JEO
NUqMLaIJz8sYQzwMLqyFjYung06QmLZXFZB0UFgH5w6/n1cOUKQS0YcNCbyoriZLWCpov4f7B9yK
VXEHfUsrNy2aVTecg9Ly60llg4B2xCa54ais+ljRfKx1214vwrK4UHPTvY+ist3HTrxW937O511e
W07VNDnqKO2Wc9wY4xW9/Yq0gOsLg3am01mMpS3dKlsfW7skq/eKFz9PVaXSN+VeSkX7k6bTEsvl
vc7AQWbhY8oNyNB0j2AvR+S6FySlzEQoSHuGqcylXzwVz7gZu1peMvALoLxzaNpeACXe48CnyCh7
MU436V1M1HsAAnM4CEjkfGJ95mhMh3lNPDv+hoIK2m3QzDI4ApUmYCiOAyfNmx8j8NWGK/jkCU6F
46sP+adJGyWl1euhfkBWxXYbjq5oXgunOnaZNLzcPN5sUBnbwwmlfuj6SuNN89UMeiczcQKf0AX8
TGyxySS/1gjuGeizxduRyjnqbnNPlHU5tNJrfRj+yipOt/IBQ6s7kgaHiM1euijgrJ9JFZHyWRpA
I0aDkMOxpZH54Yj4GURyB8VTpaHHkuUMX2vjNUv20m7LEwg6diZayIuaT4Swo0Fz5Ex5+iLS5h0O
zq9w7p2mDfbWQe3MxbrByVkRVnnXmARNOAsQZxRD5LvAFQWKudWduClF9FrnE9819I8rO53k1Lgr
4BcM9wVj4LwXVMZXorpbIFVtDQT8Ftj/EyvpDLxokSZ+TSYXf9E+I+rSzvKLN6AO+jx/b9zhnReF
bN2rGIs2ICMaZ/rnM6fp8n/KIK9XyUQ8dfYtePVGbmKbmIxd5Bc1u+fbLSK4fanmKT4Fd7ai8z3W
DnWjS1o4/t/N1kmQUL/jlre47yvjc6LrIWSqo+4Ct07g3B7HF9v+86JIz3QrAKVWl7TH4Q/y1ucl
YVhiZ96LjRBPLXjPNmLcse1TOsxzOKB1pFoBqNKOHShoP3W5rfE/c+43BuM9quHpkePEgZhdPOqj
KbrBKJnaCTnHfQHPjLwOpzZZ3mzqVN/2hPMPsTG4s/97Ohl0VPDgSkFzlDnF38qlpvVBjCmBvSZr
+h7wPKWNVug3PqeLzJ0OwSszXpu9A52aqFAbvo2iLjd3ZfhBfvP04cQXAU5Oijv9vAEK6JNqtkJ+
580cevHbGt1AA29yjm2b/ktlrFPfsc0OwTMvExNW2lSPVUCM/XU9i3S4+AtgteWkOnvaRsp7Hz0o
Zirda7nRYsiEnVBx7FVmq5llYkMuEX5cG5GyTaBCmTs0vHFYP8Fs87z5McgInD8kPvwsz/LX06Lc
r2v0atP3eBCmSEUaXOAgdIuf8y6/lFO9sfIiezT71C7IDmzyvCdtDi8CIBI4JYH/glOCqTXxmOAD
4Vgp0jTBmrOIUvh+9k39WEqq4EU0m3PNtrQnmai2Ej9Sjbrg7UnAeD4ds5MbfJJMI+q/CDV089+F
yZrtzRkIBcuSyJDC2rUQQYD6wWaEd8aTbj1KGYEvVl3avlmqimO+MnFgEsKrIGXCeF6nxlSpCuzz
t4Z7dkV66gBM8YRCk/N/tUXrh16mFIMWoFUq998meAqRSqW4XTu7WGoofo5DdiaNAO1i60wFw/qw
AxcfpbExevbifzRiUWdtXllBIEA7XrF1Nh6yY4ctBbRnQWRYv2+UlKCDipimlmElhPsV5OnczBVj
2194p/5/+uw2Yv3IpuW2sFq7mogFnikjxeZF38jI+huoe0I0w64Ak1TBdOA0Y8bTXNZf6GvRr6E1
4TFyBA45E5jbLsAlTnKclrFBaAqFL3mz5yzUPdmRz6JgvjVENXnapKp7DL2Q7P1CazyKMYAcFxBk
Wm/wVyFeUb0JcVoUZRmbFwC/uTIF1osEfRAl+eYAEX9reuL36EpTLSO35vMGLFhxfeoFEVYuslZ2
T7nzgE24UIfrvbFhYrLrzpUsTTHD+HTB+yJ77TkOj6s/IEIxcE4MACMx6d3ZWibpx6GF5DXk9F8l
UYShTs1idQyc52nG90hLBXXq/O4WolvfPsMgpTfmvfZdPG1JVxosf2U32/A8ShybIcwL+8nXF5Bw
xZ4W+KI4Xiu1G7Blq4OfJs9+fFOX25K5KgyhS59QWhM0kNZ+jlvzTpu72cceh0kNZs4b/k2f9Ljc
dvPcjLLvOmGgEzyibuT46E8do0wZEE54/pnQajl+zWoHSLZT/pzhNw+pcVCbTJIKbgsrRqX7mo/A
1cz3TcU/IuLXpOOhaqktQJ5xeguDyLLQRq82SlwIC4ASaCPGwwE1rHdFdnPuPiX4erT4tcu+3Onk
U86JmlUng0QiflTxEQsSiM85QvHXmrB4NSPscVs3T7ki8rIBKuibPRStf9VYPbKrI6VtHjw+9tt9
Zam2KCEl8rYoHYVrClOr0dvmby6dKt2AO3mye5YbCETp2fvtXtm8WnRBaefLhJnKjmMhcud9xlu1
OYy/HJKaX8jEC/+PjXVUrcLiXWIuzA0w9Ijciqg0eoToY7lR42HUR/ZktK0OFQ+ys24HdK04ykEo
joCVmC5ATjmSs8Ff2LhDnXA+Pv/TTRsg6HtiXMQvMXgFvIH/OVt3y+T3DTBjoSjByfgvVg3TMtII
c0x+7sbK+yd6T8+DkRxBFogQU3c8hH9XS1vK5W2VP22FNUXabMIVhpIiYHCWw/31wzEn8z1A1qbw
0pX64Xoh5hWdUgwJFIiwYdnO6zb65pJrcgi+Dpo/CAhfsbuRYHUpUYKsOvo4JlXedhBmCnTr2BOR
tQLocUcW23HsFLyLmq/glJGvmzo5lrmP+O5SyQJH/91OOjT2WUozHLbaWOF1fSM885lxvZWsZadN
YoAwIhsGrPGZVKAAJnA88FOQ+8Vk/agh2FAVCsnPQzj5PkzS1F0fdwFgsTBPmbI4p60lNEs3RGjy
87q31WslWn+3JeqfErLkIPAsh38eGE0mNAuAquCTcD45zZku3ye88SmkBG+0YI67x6wLiRQt5Dn8
NkJz+jJCpScAqYKQ+nDwpTsHlGHHg8FZLKN89ah/o0UfUmpWuyS6/EeqwkgQ/+I7tRx0rrQqBejZ
2t0225B5w4sHjbEBPiP0dkA6kxE4XMKeVU8Zg/P7dvtjZRfKqjCRH66MZx2Fsckqz1X/tN762sNM
KgD8j2dpp8Ar1rhVXLE8yev5M8wPlLmKqj17IHoKp5Xvh44Vc9ZLPqwUhMSZ3bDwP9hq9Z2GSJPn
tZiv4tVhptMXZyJC/qPHGe6GXaeAfvbOYzgsgH225CBg3bowll64n9OyyAPigI7JI3JwNLImI1LH
F8anjwHPO48LCCh4ccdbKBlwqcGwkpB8Zz6/8x2+1gP15mDEeA7F3ogFG7S4dv6uS2Uw8g0wmupi
sfvGQl4+SLqy9Z0Fm0p/wR/q/YTeexw7z3QS+nVTedUGVim+dIBthnmjh9ulr+jLaw2n8GUTztV1
PQSgmExLPL7uXH4dMzMjeyTLJ2LiCGWJE3SI6iFdU0C5Q/dVabgFGOJ1R0SbMVjdUDd+iISL8o1K
5D9EmF0Q4TfSyYsQX+7o3965EmVlJHYxsCNSVja8qb8vApZwe9xv1EDl2BllUmYOOj6VZWV+W3KM
VhrcQ01ZkQLhq9sDjq6QBSHFPDcPAxpUh5q7dtUFaRR40gmA1d1isa+SawdMmpFfSqwEjhPPwQwO
bv/HO43DciiOZidcH4pcgoNyzhj2QByUDQGHq3Ucri54gswwngyv1DFLLMc2VPFqFLFcbgrdXb8j
uV9Z54oU7IsjQAGyH+SE+fwTxopOM5uDIDccMRfjpeILwp/Hf/AWDj4V3D9K6T/Bo5ReNfz89Ota
SiDdDyXX9h0etw0jEuX9npOdaLzCwkdxxqYBWfx9dFyhndd3gcgsPTk2rvyPeNsEio3IOHqkkK2B
izR0n8eVC7/10OEII20J9W/HRctDFw4LCNS8PZOKfWHSGtR5Pf/pVloAuZ3fIf6vhf6B/r1E0gYY
XkI1BYMbLz5KNBpWRt3xiCAycv1X0dPC4pequUw1UjwmNB+NXJa4TGRP14g3phmgQBXUqV7+UqIt
QoyOuwe++LjKdgREK11KLxIAPcuJa4EF867SxxL/PfHlQdL8P/pktSwE9J/cSoa/hVhUsDHurRvP
HFdFCQVERto24z9s1iWzqOMGcg2Mka0YKDcckA3/erBSUqjLHRaZ5QTt0ovu70dr8QwrITqJIpml
ny8r4GpVe5zPXZRTkd5oriNnIhHy8SSWjbom90KAAgW+js+iuY0dLStiq5XyKcPcgcJrfoWE6Nsq
Dohwn9oxsI+gguKfdMneBdMWlD2Zh7PFvwqUsfGKtT9ob/Ikeb6l7H8WsMS/Qd4usAUJhy6hunhi
HFWU//F1kNjVz02jrPEZfjtWkzavUXSnLdnAeygmzbbjgWFoXyRV35tdsfq+SjEPry5/XGO4a2/j
jTzhNCDAdgifNXCZFI1KcyQnJscTddSMRV+h2MN42DCXwbejjxHwGYa9gZLNKwYt4tcoML9LjwcX
0Ra2LzPMqMk0T0KvWSaUiPaFkbyQMyHCdroQ1RDDu5vTUnWQPVL5As8y2Z83ipNbzFdKMSGcqB5F
6GGRVF8bzdfpJ1cVuzsAJisLGv+feqavgDUb+cxIh4QOQVPVkUgA3qqpbWv39HcU1GUt1qYMvVN1
wTLBTxFvuBsQt2DIF9zf9GfoqyYbA2glPSWdlenG3kzeA1HOQ1NvFlsQMmi3SCPUDVV3fLlBrdhN
yG6zD2yNyjE6ukhtaJIeZ0gf3nQL4spLr+pvhAFhIalHntEjnWUZisQM1y2z6D6IkNI/J/LVa5b7
wydsIZ0iIEQH++zn+EjGumQOUU+/gVkX2ls/YPrDIc8vGscCGQpvIQjGsoIf9xTroGDCHvDEqsoo
E5fJfKJiYU1IfUq6AiqG/xYk/nCnkdiek3uGVOUaxlHkaBlrsOWCH2O2+DVmhs/E3ocaMfcM80nq
Sb8YMVtl6I3X4oAr9x2qkcnnsgvB59XgWZLjkwxcibncM6kJy/WzP/xrO0rcP9b3Sa5skmtCcVMZ
eU0m4Rr2BcqdBP1wn/a3gm+psAKgRFJ670yF85KC2iLpBS9Ix/NkNx5TgtxIssUJudcQaihfFPuc
SC4ssSn5T8R/EcGzi2BJk+A5bLTkutdAvGrVdBjnZ0VrzmoW5ZCH/fra0asexpfNK8015XO3/o0m
Gy93zErUHIkLIEivD2OCdM7MgBwmZoc/NBaToPsBZM67eYB5hIQnePvt+VHAkMghQQ1Xrg1tlV3m
6SJ3cjjRo3PIJPIqEOIbfJXSji8igxQnI7u3OsI2rbnVguKmPHl38qz7Gyt/PQg3n3G/rFpl3xEq
MUbWuiCFjbhQBObvQyTJylpWuu/TOPqjHwD5H9WnTkQf1rZOG+0pDtTY68JFPL9Fm8Vt0aKZ0MJV
lEKpjABSVlExv+S0xShBHXUTsU6O2cu8tO9zcPJrTyUjuymt5TBJMiqnD5s/PqG2gS+qTFzMeM6/
lYXCdTkYmL3jE1WJzJF749BBjzqtfDLmcWekA3bmuSCer8u5aY4/yGVYViiGRU4iVxdXC07bVj+8
fdvq4tJALpb9HfPfhTlhxBFBZTD5Ps+OP+YkBixC0e/KA4RRzK/ArRkWf4/RZimJoBf+I000tZTO
GQv7V032HuIOHHrJje8zwBa4DkbjAW4/NiHLu61LwClHtqsgEuJ8nyNuc3r/5JaQ7Llg9qllysuq
uUDyVaAAfA7Gd7Hp2ZjU3rgAnZIYswNjhxkN2EhbYLn4YsglJ1wLb3nN1YOiNYpGbbRsC1rKtnf5
tlwqWydTTZ8UJR0ZDKWL8ybzA02lZNJC1l1LwDDVdmEkBDHO/ZEtLxwNsH0Cjnhc2muvqK0hwzWP
D3gJLNoWDylb5bGTM2Ws3Q+8O+gpUcuEIBzLV0x1FfrWCkYDBMcWNKb1FE2Sac4tBV2Gn8tl93NZ
jVH6n2Uqm7Mq/Itck1HUzkkQDwIz3K6O49Rxf6ENyT2JSLhvZzMaMnqsdjJvnpKai5QnpOyUvLkw
/pi9hKWZgomE0ctmrRJl4O4J+Zx0Aa4GYlj6JZQvlaIYddz9yjYL3MmxP8BbOr8MDK6+akKtIbNL
rNByuK7eo7YpJBQidy+R7GD4n1nR1bx9jrx5qOBLB5Jr73aVh4t0dDo7UqVcZRhKnXfJkSbNGFVu
96dTyawKHN3t+7GfVIj5Q1Q6hbBAvj+N8RUvWr2bR9jtXFijRywrGEh4dkeCP4m9QSgPPl1gpkPB
9I2xuqbi4k3bP5A50ZoXXurG/IxOFdpR9je3oa3rM94TZmKVEj2W6cXcF/euqDNXBalPNcxb/7sI
imnFS65Oym4NWIThkNicMOLHaKOv/ZErs5mzE01FDMRH3ZOTAj/y3y9EIgGZjuWIjYRqOkJKnpFm
gdK99MYwrhKWzIHf1ITTsT5Er6q12nemTyUihZJmAa8ktFdVH47UeQ6/oDkWsPUUBut/NE5YBLTR
L4xD/iZkOHNg+tWydQfWQMG+s6GbGRTSOOuz0KJMfyy2Tns6vQnpLKfBJw+bNOJ0/TB3RqfZBYyf
Q7GckKabVk79vXsS9E63a6FRnEHY+cde/SBHuHE3HJB9naLb/eGYTkNQW32032yml+xmfqVz+zeG
wyK6fBen79HaXSFSH4ZJ4gXPuGj5pNrJ0lYXtNS4DSO8buI4Yqq7+nunT0xte1OJAY/vmrv4hdS1
39caguuNUASG5E80JxqJ8Uh9IJ2Ut2u6JXO74AB+PKu2zjvky0MnsOr/eT38vv1qvnKjD5xABCJv
LjD4i3Az/f3A8HYS9cgL6G8nI6VR0vCrKS15MXfhke1sHZ2Jp2Fpif/gp+qXcEv0kriP7xsyZcW1
CTKmXs08ZdrE4cG1ufztSbcwkVBDoPWniDfcDVPnHgRWtaF6ltSR+1rbkhmlnD7DDmBz21T9aF5V
b69Ox7n3bbewQDvCrJuu1PcEVNbU6COue6LYxgLCu9BAXvIEElbvimfT259AEnWEH+05rJJA4/tH
17zaBMLFiqDDlwnWFJDp8tC/gUpbOCAAwFLqdSA41MMpqSCihz0BlxwI8wc0kvkvO9hB5LkYHFNo
mX9PWcjKqD1H8ZN+INC3yt97JUEmrRDyDHXfgptWsKa1IPla+7bnPPXRSqg9GxqGBSIy2+V8hnmS
KnhaZtYtlR8BTc7zhgeaio0XxurzeLiFtms1uJsTwKILnsK4d0KIc5Ebx8wWQQTR3dhcWy+Riu9m
kqI/6c4RDlhU1Qz93Ad7afdSRUJ0fSKUl5Zit1HSumy+tnpq/tXXtP/I/DFTzYLoKK7bNKXtXkzt
+3YryGnt5gLh/jD+kpqSc5Y4+0jSGQPb0Xea44ABOyUtq/8V5IKSQ+RGE4nxLl/cu6YPx22qoZXW
qV4b0Ce4iiDwapduGCjV+1ped0Hxp+jRYZtcELdvTqeG0U9PymHFsOROtMR3FyN/GXXx814GUHR7
/rZ/nXImIu+AzxCiLgVm1lS5VMifasLFdXLX4HlHnGvml4p5vdQzGotvrPjUlnn+S4rKrH0heUuH
eHWDAAjRi4jBJ6YJpnoWBwqn2Kdwbx5xJMg0KgOE/PEUvkSdglAdCgBqK8txauG93dfcxA+3QNIa
NyCta08C33zqxS87M2NBnU0yei64kebFWza0kxdzRZhTC13qvfrzGR5XmPL5phXDZbw4nMFLPcMj
aJtRbV1ynKxO7a0F4sFWXCRHnWM5Sit8eoXjW3stSLWDlKmbK0Gi3zoLzzK+NrRytcwMV3QjG7RQ
RPdmOnta+vCvyjlW1U/zLTAs7B4NjkV6t3mvyo8hg/WtgI+C5VZLqO+k5nsVuHsHiWpGzaJlc50S
jSU5AKdYSrln+Afrj+xL9HQ3Q4qdJE2FdQXSR20kZJiybFnUNhDFc2fSuORoyQrGONFxsEQyYwnd
a9AOGAAygQgcDjusf+eP65f26AwEw+oV1LJR8icImoP1VDMq25qP7sTNaB2UmoBY0LZWoSiUqg+T
dyTYl34VN2fum9pMfu06mpH4uZWYKOKmBKPmwGnuNORATDeCB+Iymuy812K2jHAwLLC5EPlJyZZc
dS7TBRtBW0KRk4ZixnHqcrC2i+O7o+Y04Mo5kkWiZ06DhEwo40r9HCKPJ6nbvwyKeRIeKZreSw0N
nVyRANtd1dpGDfKAQZiP7BQ7DoVH9v4UCtHl3WbOIPAtTJ7Tq9aV5Dr2O+pf9QEpr7xyfZC8t8R/
0zRiCjwqJr3Z/cVMJcWRPQe+pBj2GxKCLWUGDT62thO9AazN/4bcdE5BwdLUwhBJjbCjjO8Cum//
8dcj46NU4laTcvU/55bi8q07CU151MLLSwKBb4zK0JN+UddCPsIUHucUEvZdGAFrbwm+zbbVt8Mt
EeLLuNRcZ4qMg20a0o6cv2mgoKIZbv/etPUs3v43ZfUySo6FykTF1yTaN56gUaiK334uXEBah36r
NYrbmyhC8oM5sul26TRPyTyvzOP0/zarwVR991kWdnXgaZZpgqRD0JVTlK2n3/ukA6xOvpIHCx7S
tiP9KVijVTKj++GvQPgoDkn0iBjTJx0Yuw4eVe20zMDvZqcv1/ZKqKX61940BaVno7n1El+BFyQk
yRvz2kf5hWyGvpsHts0Uo2jh3ZSVkDXQsdW62aJMFEvIIpk676M57Ar2NH/6ha4QdFnUNtO4ZVSk
8gxxTd4sRHW+AjwkULwKjdhlIc+fJ/P3ZEYhjJzgMeb6e0sv4TpfePrTR5aURB2gT5H3AjvrE72N
wa4OdiOsze4ropGLV2Y4sVUGbbfI/UJuUW70g7cpzUZCHUk2tjeFvZzxYvtVx0LQQg3HwNFQ8du8
0so0NXVcn5L4J8Anl+uDKsB8zkx0bPNirZYnxUPL7McIZT/CBlbuVAJdkIJaygF3mLwYmxVKPtzm
xd48+1r/Q1R7j8byYqMaHmvzvwwWAeJR+5OfIpKydY5nAaQxfVUy4hSRMBqnIaTN1dGRg7yxGMyI
BjQCh80zKrfYdWZe8uVBU2+OAC1TkiOfU+q8fU2Rr5Bs1ohiQaLvEbmSaFddC8zQHvt/bmWio6Zy
AhkKsQXChQPYb5QsaNnjmofUEA40Xh2tPWLw+m3Ixa52qsWOa/eeyh3qy5dnn/eXcQ/xBlew6caZ
xxr2XwAV+QyJ5D3icaUlXO6lG2+jclWFOOPF9ueRoUtpbbNXV+OtrXm7n4j6CUsc99XWHGtdGna4
xQLs9qL+rdsKOzUkxcyy8LOmXcKA3iWCZwGdIPilHLlr5jmA5OTzgDGCp+Y04PfNPHxIFas++2cp
+lxQ7Jq8Lt+7imqp+fnJLiw3AI6JUY3kTq0ti/qlSuy1TMOE12CGrhc2AhkdHPEXyOUWP/ILx5AY
JlYB/KpjRYQUYgAqEo8U4EwGu/GQyXSFc8zXEgoZv4PUjSUV6ngLq12CqJ5X9qEEmrySMSyj/zo3
SjmHHcJ96tCRiOnuTJBEIbuprrpErzDB7Q8+x4gGG+/3dEV2PTtp6UBc32chm+wOgPV7btm1pFoJ
k8Wyj37ADQYwaz7Yp9NSt5knmld9+L3gVcsaGw54hxf+XW1O+gF58JW2IMN4C5K7YK89k9QQj5r1
PPpHCvE4HghLMsyFn5znO3UOZZ9o5Wz+gAmuK6m1/c62t8z2VYuf0bAORaq2aZ7ox2IivDApUL5T
p/+IXID6/VjbDu3rgqZJh3nvYVxXnT3w4lzuEkKHRnNZ7iVF2V858ZxFPiOLvUQJFhYVhPDLv1UA
zSBewKga1ZIxW0rEuH0NJFnAmqxx+ahUPFRky/Zg5JgHGTDP1iRkBq4iGE1rcOR/IE4xh/+SoH4f
ECWHSX/MTAA6ui0/UAhzSNvD0mlGGME/EhIqhamSzLpOmsPYiHqWUr9e5nkCisguV83KpY4HxMNz
+qY2zolZR6zAldQLrBmaJ+TAI2u0r+D4EtDS+Pbd2NTBvBqxAQR+18k/E12/3DKI8riWjOjEf1Y7
coPpRMhLYtzNju6hvVWg8o2i2zjqsJ5Ztkh4MvSvc8U6zTS/pVWADv7rkvHiVb4PykqW0lBblmpT
iGiQYPSMloMrPFXJWyw+cBo6Zi86NVSUeshjjp2k/NuXeJ8OhpZPVDUwt5+d3yPCvm7GzG4btR2X
VBIC2brrmvJdjoet2jn1rHQQCIN3lqoVJSqRP/68DjffAxzbWUrEMO7PtYD6pCy+99zxOSs1SUFa
Q0AeWMsis13PBViA7cFCPwzUlwNNGpdPgapuSrRta2AWyNap+NBIlVZaGKNEjwLZ+kP/rRueqrnM
cJ1H6xgGX3DyyjOK/v2qxGhbbsaMbtifioLQlkTykBTWkEnVNAOtcoV0S2WMOmMB/6WZU5HsbTz7
6LETyuunjqFBlCkBP6obVnA8D17NNxrbS+RiPvvCFu5t+kX29g2SmbtRAY+T3IwKSLffdI0eD7Cn
GjtVdeDesK9jQyaMJaQ1USpNcoyKWAMaNWtVhYhEmlg+yyUJoM+RFbU6EmDXd3LBksbpaBAdiDRQ
nhCfNQKfh4QlQ/jdvPxH3xhW2qnMOoVIfjT9HzyX60oSAYKOtZgsZLNktJIT4gvAGnmSg2wXv81h
c8QbZN3jn2evN3i4femx/U1IGRVh+FJZ77WxQJKeba3Q3mClPqrSGM+15ghIF2DWouz3PSyuIl9C
5hjt8agAC5uju8i1E00nKW4a7F88eg6Gt7AubCpWXviysTzy4rhl2bSf5PddH3ceVfdcQyMgS7Tf
Zy4jNrn1QPxqPDeCpYOKFbeG/PRTWJ8PCXg42zIfCev931QXuRL/kNHaLMkD2VJqHuWeWMH2KAmo
5nvIJnQpSaG84AopWimb2xttFMTKINpX7LzM+3tWAfEHyL3hwowML0dqH1ajOb0VLf/eBn/skzIU
MeT07hMIBNDm0CkC/J8APEBOBNzzDMrbtYTPjHClp+k6PE8WXem1H/BRQP75zgFf4nNDdUw1xmum
1O7Uy7W20Ctap6BL3XYvFJuub5hQIoQQQqibAQMdMJvwix8WHQpy1jekj2DN2X1cEkzWmvhYJdD0
hkfE4BJNhHJOm2PP+rV0YmTEjijWEBDck77WdSylMtFMaCvxyGYNCCcK744IMimPmkS2b26HL77N
lN9t8pgpm6nFCK/lZQn6AJWVo/jVLMOZjhbDhqCDPOaIBEl1IGiXdrZB6k/ga5ir/Aa5Tmdxj3C9
wLp6qYvY3Uddu4sJyHQEJ3DM8Ai5Wioj5AaRkKMFEUbbDF7z8ZvZSsbzkYSHwj/fKkWzkOdeM8vz
Fi8C/Bva8m2buEGTtd568slRlJKVtrzd/Ld0CKC//31++0k9xu4dGBkIZMBgo+Mqlencw2+eN6uO
xgiWhTp1xvgHfFGYG4YxbYactKdWQ8/bf/hAObXKbWQPdU9YD7C8ANJaZ4FFA27qJI4YTyGdCC8T
EzpgftJOgWMoSqLLPhU0kR9pslc7q2hpurHYBDfaWkhDGg08LmPsnZp5x8bUpL6GB0wPr94kSt/L
eUFw2PgCgtIPpMRrNkXPtsX4O+4mAqxQoMe1dz2Rq+TKyurwc8p69LWtM9KZmJb0Fo9TsKvY+8R4
6Vyl/G0VZMN0auc8s4tO5tTbhHIUS/ZBrp9uAyOH3LxDUjH2Aa0/xCtd1VkIbmcPFSnchXKQyxnT
9tv7hskyJRTtBVXFUqTkd+SVwrZlxpDuI+fQJaqdCP3VAmpylh/qDJj/TcA+Y+OTCg5PUOEFvV0o
VSvN1N3fYK/wBiYbQTzxgsS3ipJKX5oZZ/M4iMoLXEqW363x1PU7rbYqe7DNf7nFfRgL1XZQ6/CY
qOmShayIuEl5rZGljptfe/BNb8bLWm8ff0lrlYIBHynwyDq9jCVBAjfOz6dEyfBv6nppz2ibtLiW
hgWBO7X5wnGKyOJt1BGQuxhfvVSXiAtyv2OqjSTyyBQsCWZkVDc1qs6UKrqtDjuesvczFEZhz7sn
7LELxzIOl1OpymJRuQS5lk66znicIh+Gt1f80CGEgUX+jMAycNrdIOwlCtO+bh0AbQJU7pIKTCIg
ceg9YDLQcLiE53f0zJIGAM9z6p/gOJxKVwhGKUDzZlLA+X9DUvmwm9MYTd7grWNvG7mg8Rd+bh8W
oWAYfizDEk5q7ehYw+GesC8bHWZQ9TeItZ5zx2XByiC/xaSLt2TkSyeQv36KfZfUHfZw+Viya935
bAFmkNL6cIRS8Qa2ZNjCZNiy4M2+YCSUhxTtAqfzH/IGqk659irOOFx/WWIG9fUM37tuLdWY+6U1
Vx6Z9JDfp+1Vx+ty9hsFAoNiyJ1mtrqaIc+gurM+RiUUFDBIusCeDy4j1896fX8XiCDg0l9VjuSw
i8Xe8EoKVBHTxYDPZJGdvT85Ucm1m2X7vMDoWXD9Kf0CJbBrmegZYdc7yShyji5ovyYa4MZ8PhtS
fDszIjKVXbS325wyL5oo/nEwVvpWJ5Rd5cmz+MRNQ+iQfLisAwPuGaSmnisd4nYb3GxYAHwFqFo6
10x/eYjGtSOimTjqhThXmHDGSUiwrdLtQhZtwy7Z/q4UZzyMxkFKE35GAGsAcedHZvoLQTHjjMSk
jLjMPpN0rf2pmZF7BFP1D3CJVoDLiyCiqO+bJkIHm5F8ZyrvEoUc3mROS36H61yZaa22hhMZ2N/O
B2nh8E8BeIEPYNJVLyMm/vwoAUiFllnjcBfzmDxF3q491n07ArXLEcuF1eNVBIZAh6fhZTakdS1n
Z+w7F0hFFu0hwhEGRbrrXOJOAT1HonaY1t21Qm7O2WffzoLm+rEPOPhQEcW9W908J8dJOD5GfKT4
ACIajCjhDrMv9zPeTDEK94G9KG0aoli+yYy4JzqjRUbw4D5BngmXNvkwpw3N1MiXdA0Wnapq6Cwh
vc8qWC5v/MZaB4vjYJ6ZBDOwTFgm7+LWsutmDvMsG5Z70/b1Jxcf7knMsJgsdemvRmkP7muRf8Ds
6AmkQuMO14rlEvdU/uFAWGMIrdokNatQe+uM8o4tOwBOGG3FtCh/AFQq6nn2AATzo5HGEAimSX8+
pnFqMSD0Mo32n3Oj+jrHDFNuJEyjznh+CZsqR4Zdh/98pWkEpCwNjQaeEw5Ltg8vd8ycoWnssSJS
ECH0noE/Lv6VsbmtQGHToWLKYOu72x7+lKvEbMlZ7T+JUwBZ+E7eqzpPPKV4g3PwmfoueGG2rf01
DigPlN+/Cb5MfIhZXBUH7OUsgwgVwAlLgxgoP3jGY89Cm4/BlUq/bInIF8AuRDgqqdaRgUV0Kcxk
oe7dj+9to8DoEwSMCtqqmrXtnFz/zCov5/PSWrZXy/EonvzXNWC1z7wbWhXk+aRuYyBu++cSrjEf
6TQcHaZQpZ6gP+RBHAXc0GXEwqx7uMns1XEkhWgpIghsTtDnbOESzE9k9K3zmup66vDheaY3nag1
z2+fL7DOnXGSzIqO1Waz6sxHowLsl8asJfylHQsOoBy+qXXW4s1dRDkkgqOQp/tTuDiZN7fArRQj
twWP5aJzIkVILJdDLh1cDTrDQZdl6JXevxoca90/KGEFs8d2qdwTmCOXhcFcSWQ1384I+z0Ss0VC
FGG2OoYfYPDpBE5vmpbamwfWjrF0GR0PVblTFfQkAXKuyKhWmTNgB8sbvdUqreS4n2Nm/w7znD+y
CTBWs1y8jD4X78oL45kDY5fxNa8r5rlLl6ZziL8YrsUxSpynbwjVEqOdJIhsMubw7nIniBMfUE3K
wZp+3bNRqsVxqF4ZwskRIT0ebzBkY0kU7ONWAfHQavzwZx7UtcSbttz2ps1BrgpUy4IIRVP89Fmo
Ccdva1gD+PrrV8cT4KAe7fP0PpIC2oBZFoHO2klCMdkLztJfkFoBvCx6WzPPomTzuClcbEDWPv65
Hng4Lxa5TeKdDNgy5wWLahB/HP2NO7xoaghDPlknehcnoUbS0tHXfhDEPk88LUou+AQyOE8qiWju
FHClci3EOr24FESr3DNdbn6uwyzgueP1wKrZgVPw4fEpVZdbyZDjij6GKK09/2njhFIfr0Bnbze9
b1x4hPPy406y5kPmH4lxYd5+6RLqaisn8h8K33ajU2Ot/kkvP2M+2Z2ydS8A1XOgjnPe1dGSXsPw
KM/cd0rcjgX+QQUYvHoQsU0cxsEMdfw9Sb/8lOg8NHPqEbSeHPtVH7ZziIs2cw8QjFAvz1pNaOKI
3KgfyeIcmwmInbqvPz0Bpxive5rRdadfqT2dRdSzAmTdM7iYFZMgpNkmpM9xcXnD0KDQPJgpA03y
Y4J+ACibRj28UFeGXDaRJCSXXrGvvZNWcVwqINQ+cOhZXaLW6JLauyAQyUkp0fXjmA8PauUpDPAd
VisT1yFu3+IwCACQVhHqqbJBXrqunhBAkGdg8XSahRc7sTXPG7dRtbCxVorRAg1ZpoDt9wUAL6J1
je6fv32j7UH3qJnWuLlXj0q2w5DQY4wupQSKTlGPK1opDw8MME0FZjDENiRORtQ5rBDMMWvyMKUF
GXZTvQdjoHHHAFKjouBVyP2CmYhEPQlHSv2p52HELgZyJfKDDkZEJ9sqRHW8hZmOEM6sE4HqOTVd
xVDhgWVmXKa2k+c/Nf7R0JkU/LkPJBG0W7uXZwA+taWQEHEpDWD5z3NqKWQ6AhI0VLwn6CC0SrpJ
MFafqfuPqbzG9cad2MZcdLnoP1p7k3ebibXH2JRsqQ3nI35NMa6S7V5pXpxy0CPX9zpHeo+t14nT
fP4BH/ujL6LEyyyfGVzXTfvOd0SqADm2dQ5QXbRo0iv+I1y6+EuYOCyAHqFMpBKs8+oQhBfRU6fG
fqjo49J5dGoV/zRUrHfOVf7ueYKY9InMJcr2YLw2J8WGWV0/OrKArxP8glh4HKxO9Rp/WhLPuLHi
E2OB24famFo/ODXCJtz3TjC7sGZYHpzXU2udOkWD3BV85SKFtXufvI2bm9zy6DOwN0B8FIwdQsdU
WkEcdWL4uVMNTtMoK88j3zY7K+oboc9UAqPWWNMy4LhBJ8Nq71T+9sTVMzxXz7elBOQfIM4p4uB/
bEFqBcr0hDR+Elj++sBClZj1G+flWYGNuv3hCzpwUDjVD43PzndU+WpiJ9ezOwocSlsCmGfEhHWv
J3V5O2B+7ON+LYq2qpY3b4zgjARFz6rXx+d97M6XiAeGLv72WWQgPgtwFREeuid6Aq20HAFb9/qV
GK5XoHaJYmudA+OWS0Xg/VJ258Jk13bsnSN8Q5dos6uIm2RMKrMukitvGeDKFxU4pe3ZmNRtrEmZ
T3EE2iVj6qo5Q4u6lzpEfNXT13VUQ3sHF7adok9v1D97zejVFv34q6gM56WUAL79Z4mUoG1nhYP/
pdkw6f/5gR+d921ScgADkLuWnIXXqcpFLLgTrB7Cn2eH/c3FwoKe5Ij37wOK5bK2Pspv1zwIX1Ai
hQPLygD7Xfla2+7iAIoGFLnOrdJREBj7Ru8rHaaLKOFmPJJt76OlfG6tFL+ARvEstFNGTQWK/adB
o3Gm/phk2ecZLplY4cZLFLWt3K3LK5+XtWvyt9DrDdcN1ggXuVMruWpy5CwwOigUHQXfSbwmdG5d
NnqQJj7U/82OSAmpdH1UzD55mEp9dUYjABLhIyv4rtkMio4FrzAMUrgk6hkvGv2o63yy2tZGs4qn
Hkf/2fE8iURXMk+Yeh8AbgY/7lZFe2p5SfBN18ft+VBDOAFwWc3cGk8o1hkHmxg2jI03rgYIKFWE
Y989zu4kywGQsubL5HSdC66/55rL7d/yBDAIWGoQ99dx/mP9oPCBJLk8YRROr07CuXQKlUngrGvp
P9i/Fb3LHXJ7MhFpALE5o1enHNtgO80KsfYzJ3oaetr/9K4CXvQDnoIx2xafBUio/eku4RsIl7na
BXx0ymm4NIYFalFF39OKITSOGH63bF8KbC9LeV5TjhpPuLoAw5mrwTF27HOGiLjzlmbjRARxj0ou
rAbjwJTbOEyO45dfp19Hxo9zQx536ktOuo4znFB8+gTfqXxJBX0XCS9kh+KXJaGqPKGXKms+BEnO
ZyJg/IDbaCRk9YCml07kFqMowx8C8/psJsHlVuDAUkyHHqyT4nPnUXJMe+dOr2dzIeL+5oMKSjwi
zLfVHVKPvirTw2ZbElSOuOz3ZBSESWXTCB8gzf+NblQA6Iwd6la7cWycRLwlnWW6Lx/Vrr5Iw+Ws
La/me3Agoa2XVSTriO3vgqeI/7HHspyfhkt435FDMSkoSFn2ht5eZZBMhVn9bMKbNiyA5VlXhVD4
TA5iwJTBbM3T7qzWbZRpQY6gAgGcdzPzGgWqw1XSHCbxmhwFOEDlxIWZMYobrbxTL3Xb1AW4Pgc4
6LeqTSUS6FlaGInwfruzqvbn6g4hRTHmdx3IVwe9o36sjC1mifo7GyGmjev2h9abXzwZRhvSiSsw
u2UF0o8liDktocTNLfXDRX4lozjsDMZrYfteYA+Dwy2iE+tSGnN+bqsGG9BYVNWN1eoZbn9lM6pj
ix0mGaQZtnfUu+d9yKKS5NS/cRpnlr67ebxTqc8RyvBvoS/pxybmkFdtuJYUB1N8QUYudYUWhcHY
FVwmlTrPva37FhNcgoV/J+qokrd6HrHwyKmzlw+d5Y50VcJl+ZSM9lgdaXaGnpH4/EGNt7K5h1Ma
eqVmTpuQ2FHGOEVRhyQgMahyz0LdxPcsWP8GOgg38EcWddE4+HgMm7wwSC7pa08zHD1cGx0Rz9+Y
8/lV6wajMePMATVdZXtH/IuiXT7D7R2mtb5KaQ+xq+RxraIHpdjuje5Kf6zA/qop2XblXM2rk/ls
VbQJzZvfuvXBUKlMPEofgmpsO6dXwG2a545r5QSK66sho54MMzKiyyEaajiB4/eDt7QiwkTy27ON
cDGKq9HerODGZDaJPlOnR1ud8Ok1zNHozKhqavNCbGfYT2+aYGs49Q9NKCMH/aSGcNHlU+auFAHk
TO5Qp9mf1c74OcAy3UQoDz+kB+rA88RokVnsSs4/LUqvdIQaykx8mNJKFFgM7PiyKr4yr++fmv75
mDYyDRih0hRrS4SRoVhB+XybXUunVJTOk+8O2FDZfaLyXmQhIerCogZxDg5q/Um8z7X4BLHKgB2Y
5jB8sGv5cZ00TLlcupUjcUY9eYUrSspNinxxzfG4boVci+WnOZcyumSPXBG+NrkI5eoy/mHiIW5t
qCUN+5HpJRUal9AddYE3wMY7ULLW9+htOYVJ8//L9r/JaGWzGBS9WxXjFah+AZBBXL0b8h1uUZsd
tKlMKVnNYfrj8ohQjVq7NFzyKX2AUVSYpShkbeRkEIan8VpXNeqoFg08MevmJghXhtUHseopRl5h
khcqO968tzhrnRJQBhY/2NThF5G3IWi2mXWWF+yn76gSr3AxgKbCNYjYGoh6v+PiNbW5+OdbTk5v
xd2XkQTj61g09i9ObGQy8/CehZDMfTXOhtzJkKSWzRX9R1PYKc81Y+3zOZcYN5LGv43RxFygYeCv
q9TRkncUilMxGCezwr99DA8BxeUoYR6tRXi/CMStVqmO52+R6TUdfIOyvgqu9c8+/IO4zBRfVw==
`protect end_protected

