library IEEE; 
use IEEE.STD_LOGIC_1164.ALL;
library work;
use work.tel2000.all;

--ATTENTION awuser, aruser, awid, arid sont d�connecter

entity fb_axi_inter_wrap is
  port (
  --Clk and Reste
  inter_aclk : IN STD_LOGIC;
  s00_aclk : in STD_LOGIC;
  s01_aclk : in STD_LOGIC;
  m00_aclk : in STD_LOGIC;
  aresetn : in std_logic;
  
  s00_arestn_out : out STD_LOGIC;
  s01_arestn_out : out STD_LOGIC;
  m00_arestn_out : out STD_LOGIC;
  --s2mm port(S0)
  axi4_s2mm_mosi : in t_axi4_a32_d32_write_mosi;
  axi4_s2mm_miso : out t_axi4_a32_d32_write_miso;
  --mm2s port (S1)
   axi4_mm2s_mosi : in t_axi4_a32_d32_read_mosi;
   axi4_mm2s_miso : out t_axi4_a32_d32_read_miso;
  --MIG PORT (M0)
  axi4_mig_mosi : out t_axi4_a32_d128_mosi;
  axi4_mig_miso : in t_axi4_a32_d128_miso

  );
end fb_axi_inter_wrap;

architecture sim of fb_axi_inter_wrap is

COMPONENT axi_interconnect_0
  PORT (
    INTERCONNECT_ACLK : IN STD_LOGIC;
    INTERCONNECT_ARESETN : IN STD_LOGIC;
    S00_AXI_ARESET_OUT_N : OUT STD_LOGIC;
    S00_AXI_ACLK : IN STD_LOGIC;
    S00_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    S00_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    S00_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S00_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    S00_AXI_AWLOCK : IN STD_LOGIC;
    S00_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S00_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_AWVALID : IN STD_LOGIC;
    S00_AXI_AWREADY : OUT STD_LOGIC;
    S00_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_WLAST : IN STD_LOGIC;
    S00_AXI_WVALID : IN STD_LOGIC;
    S00_AXI_WREADY : OUT STD_LOGIC;
    S00_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    S00_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    S00_AXI_BVALID : OUT STD_LOGIC;
    S00_AXI_BREADY : IN STD_LOGIC;
    S00_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    S00_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    S00_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S00_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    S00_AXI_ARLOCK : IN STD_LOGIC;
    S00_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S00_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_ARVALID : IN STD_LOGIC;
    S00_AXI_ARREADY : OUT STD_LOGIC;
    S00_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    S00_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    S00_AXI_RLAST : OUT STD_LOGIC;
    S00_AXI_RVALID : OUT STD_LOGIC;
    S00_AXI_RREADY : IN STD_LOGIC;
    S01_AXI_ARESET_OUT_N : OUT STD_LOGIC;
    S01_AXI_ACLK : IN STD_LOGIC;
    S01_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    S01_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S01_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    S01_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S01_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    S01_AXI_AWLOCK : IN STD_LOGIC;
    S01_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S01_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S01_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S01_AXI_AWVALID : IN STD_LOGIC;
    S01_AXI_AWREADY : OUT STD_LOGIC;
    S01_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S01_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S01_AXI_WLAST : IN STD_LOGIC;
    S01_AXI_WVALID : IN STD_LOGIC;
    S01_AXI_WREADY : OUT STD_LOGIC;
    S01_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    S01_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    S01_AXI_BVALID : OUT STD_LOGIC;
    S01_AXI_BREADY : IN STD_LOGIC;
    S01_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    S01_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S01_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    S01_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S01_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    S01_AXI_ARLOCK : IN STD_LOGIC;
    S01_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S01_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S01_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S01_AXI_ARVALID : IN STD_LOGIC;
    S01_AXI_ARREADY : OUT STD_LOGIC;
    S01_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    S01_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    S01_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    S01_AXI_RLAST : OUT STD_LOGIC;
    S01_AXI_RVALID : OUT STD_LOGIC;
    S01_AXI_RREADY : IN STD_LOGIC;
    M00_AXI_ARESET_OUT_N : OUT STD_LOGIC;
    M00_AXI_ACLK : IN STD_LOGIC;
    M00_AXI_AWID : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_AWADDR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    M00_AXI_AWLEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    M00_AXI_AWSIZE : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    M00_AXI_AWBURST : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    M00_AXI_AWLOCK : OUT STD_LOGIC;
    M00_AXI_AWCACHE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_AWPROT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    M00_AXI_AWQOS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_AWVALID : OUT STD_LOGIC;
    M00_AXI_AWREADY : IN STD_LOGIC;
    M00_AXI_WDATA : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    M00_AXI_WSTRB : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    M00_AXI_WLAST : OUT STD_LOGIC;
    M00_AXI_WVALID : OUT STD_LOGIC;
    M00_AXI_WREADY : IN STD_LOGIC;
    M00_AXI_BID : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_BRESP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    M00_AXI_BVALID : IN STD_LOGIC;
    M00_AXI_BREADY : OUT STD_LOGIC;
    M00_AXI_ARID : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_ARADDR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    M00_AXI_ARLEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    M00_AXI_ARSIZE : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    M00_AXI_ARBURST : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    M00_AXI_ARLOCK : OUT STD_LOGIC;
    M00_AXI_ARCACHE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_ARPROT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    M00_AXI_ARQOS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_ARVALID : OUT STD_LOGIC;
    M00_AXI_ARREADY : IN STD_LOGIC;
    M00_AXI_RID : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_RDATA : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    M00_AXI_RRESP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    M00_AXI_RLAST : IN STD_LOGIC;
    M00_AXI_RVALID : IN STD_LOGIC;
    M00_AXI_RREADY : OUT STD_LOGIC
  );
END COMPONENT;
ATTRIBUTE SYN_BLACK_BOX : BOOLEAN;
ATTRIBUTE SYN_BLACK_BOX OF axi_interconnect_0 : COMPONENT IS TRUE;
ATTRIBUTE BLACK_BOX_PAD_PIN : STRING;
ATTRIBUTE BLACK_BOX_PAD_PIN OF axi_interconnect_0 : COMPONENT IS "INTERCONNECT_ACLK,INTERCONNECT_ARESETN,S00_AXI_ARESET_OUT_N,S00_AXI_ACLK,S00_AXI_AWID[0:0],S00_AXI_AWADDR[31:0],S00_AXI_AWLEN[7:0],S00_AXI_AWSIZE[2:0],S00_AXI_AWBURST[1:0],S00_AXI_AWLOCK,S00_AXI_AWCACHE[3:0],S00_AXI_AWPROT[2:0],S00_AXI_AWQOS[3:0],S00_AXI_AWVALID,S00_AXI_AWREADY,S00_AXI_WDATA[31:0],S00_AXI_WSTRB[3:0],S00_AXI_WLAST,S00_AXI_WVALID,S00_AXI_WREADY,S00_AXI_BID[0:0],S00_AXI_BRESP[1:0],S00_AXI_BVALID,S00_AXI_BREADY,S00_AXI_ARID[0:0],S00_AXI_ARADDR[31:0],S00_AXI_ARLEN[7:0],S00_AXI_ARSIZE[2:0],S00_AXI_ARBURST[1:0],S00_AXI_ARLOCK,S00_AXI_ARCACHE[3:0],S00_AXI_ARPROT[2:0],S00_AXI_ARQOS[3:0],S00_AXI_ARVALID,S00_AXI_ARREADY,S00_AXI_RID[0:0],S00_AXI_RDATA[31:0],S00_AXI_RRESP[1:0],S00_AXI_RLAST,S00_AXI_RVALID,S00_AXI_RREADY,S01_AXI_ARESET_OUT_N,S01_AXI_ACLK,S01_AXI_AWID[0:0],S01_AXI_AWADDR[31:0],S01_AXI_AWLEN[7:0],S01_AXI_AWSIZE[2:0],S01_AXI_AWBURST[1:0],S01_AXI_AWLOCK,S01_AXI_AWCACHE[3:0],S01_AXI_AWPROT[2:0],S01_AXI_AWQOS[3:0],S01_AXI_AWVALID,S01_AXI_AWREADY,S01_AXI_WDATA[31:0],S01_AXI_WSTRB[3:0],S01_AXI_WLAST,S01_AXI_WVALID,S01_AXI_WREADY,S01_AXI_BID[0:0],S01_AXI_BRESP[1:0],S01_AXI_BVALID,S01_AXI_BREADY,S01_AXI_ARID[0:0],S01_AXI_ARADDR[31:0],S01_AXI_ARLEN[7:0],S01_AXI_ARSIZE[2:0],S01_AXI_ARBURST[1:0],S01_AXI_ARLOCK,S01_AXI_ARCACHE[3:0],S01_AXI_ARPROT[2:0],S01_AXI_ARQOS[3:0],S01_AXI_ARVALID,S01_AXI_ARREADY,S01_AXI_RID[0:0],S01_AXI_RDATA[31:0],S01_AXI_RRESP[1:0],S01_AXI_RLAST,S01_AXI_RVALID,S01_AXI_RREADY,M00_AXI_ARESET_OUT_N,M00_AXI_ACLK,M00_AXI_AWID[3:0],M00_AXI_AWADDR[31:0],M00_AXI_AWLEN[7:0],M00_AXI_AWSIZE[2:0],M00_AXI_AWBURST[1:0],M00_AXI_AWLOCK,M00_AXI_AWCACHE[3:0],M00_AXI_AWPROT[2:0],M00_AXI_AWQOS[3:0],M00_AXI_AWVALID,M00_AXI_AWREADY,M00_AXI_WDATA[127:0],M00_AXI_WSTRB[15:0],M00_AXI_WLAST,M00_AXI_WVALID,M00_AXI_WREADY,M00_AXI_BID[3:0],M00_AXI_BRESP[1:0],M00_AXI_BVALID,M00_AXI_BREADY,M00_AXI_ARID[3:0],M00_AXI_ARADDR[31:0],M00_AXI_ARLEN[7:0],M00_AXI_ARSIZE[2:0],M00_AXI_ARBURST[1:0],M00_AXI_ARLOCK,M00_AXI_ARCACHE[3:0],M00_AXI_ARPROT[2:0],M00_AXI_ARQOS[3:0],M00_AXI_ARVALID,M00_AXI_ARREADY,M00_AXI_RID[3:0],M00_AXI_RDATA[127:0],M00_AXI_RRESP[1:0],M00_AXI_RLAST,M00_AXI_RVALID,M00_AXI_RREADY";

begin


interconnect : axi_interconnect_0
  PORT MAP (
    INTERCONNECT_ACLK => inter_aclk,
    INTERCONNECT_ARESETN => aresetn,
    S00_AXI_ARESET_OUT_N   => s00_arestn_out,
    S00_AXI_ACLK           => s00_aclk,
    S00_AXI_AWID           => axi4_s2mm_mosi.AWID(0 downto 0),
    S00_AXI_AWADDR         => axi4_s2mm_mosi.AWADDR,
    S00_AXI_AWLEN          => axi4_s2mm_mosi.AWLEN,
    S00_AXI_AWSIZE         => axi4_s2mm_mosi.AWSIZE,
    S00_AXI_AWBURST        => axi4_s2mm_mosi.AWBURST,
    S00_AXI_AWLOCK         => '0',
    S00_AXI_AWCACHE        => axi4_s2mm_mosi.AWCACHE,
    S00_AXI_AWPROT         => axi4_s2mm_mosi.AWPROT,
    S00_AXI_AWQOS          => (others => '0'),
    S00_AXI_AWVALID        => axi4_s2mm_mosi.AWVALID,
    S00_AXI_AWREADY        => axi4_s2mm_miso.AWREADY,
    S00_AXI_WDATA          => axi4_s2mm_mosi.WDATA,
    S00_AXI_WSTRB          => axi4_s2mm_mosi.WSTRB,
    S00_AXI_WLAST          => axi4_s2mm_mosi.WLAST,
    S00_AXI_WVALID         => axi4_s2mm_mosi.WVALID,
    S00_AXI_WREADY         => axi4_s2mm_miso.WREADY,
    S00_AXI_BID            => open,
    S00_AXI_BRESP          => axi4_s2mm_miso.BRESP,
    S00_AXI_BVALID         => axi4_s2mm_miso.BVALID,
    S00_AXI_BREADY         => axi4_s2mm_mosi.BREADY,
    S00_AXI_ARID           => (others => '0'),
    S00_AXI_ARADDR         => (others => '0'),
    S00_AXI_ARLEN          => (others => '0'),
    S00_AXI_ARSIZE         => (others => '0'),
    S00_AXI_ARBURST        => (others => '0'),
    S00_AXI_ARLOCK         => '0',
    S00_AXI_ARCACHE        => (others => '0'),
    S00_AXI_ARPROT         => (others => '0'),
    S00_AXI_ARQOS          => (others => '0'),
    S00_AXI_ARVALID        => '0',
    S00_AXI_ARREADY        => open,
    S00_AXI_RID            => open,
    S00_AXI_RDATA          => open,
    S00_AXI_RRESP          => open,
    S00_AXI_RLAST          => open,
    S00_AXI_RVALID         => open,
    S00_AXI_RREADY         => '0',
    
    S01_AXI_ARESET_OUT_N   => s01_arestn_out,
    S01_AXI_ACLK           => s01_aclk,
    S01_AXI_AWID           => (others => '0'),
    S01_AXI_AWADDR         => (others => '0'),
    S01_AXI_AWLEN          => (others => '0'),
    S01_AXI_AWSIZE         => (others => '0'),
    S01_AXI_AWBURST        => (others => '0'),
    S01_AXI_AWLOCK         => '0',
    S01_AXI_AWCACHE        => (others => '0'),
    S01_AXI_AWPROT         => (others => '0'),
    S01_AXI_AWQOS          => (others => '0'),
    S01_AXI_AWVALID        => '0',
    S01_AXI_AWREADY        => open,
    S01_AXI_WDATA          => (others => '0'),
    S01_AXI_WSTRB          => (others => '0'),
    S01_AXI_WLAST          => '0',
    S01_AXI_WVALID         => '0',
    S01_AXI_WREADY         => open,
    S01_AXI_BID            => open,
    S01_AXI_BRESP          => open,
    S01_AXI_BVALID         => open,
    S01_AXI_BREADY         => '0',
    S01_AXI_ARID           => axi4_mm2s_mosi.ARID(0 downto 0),
    S01_AXI_ARADDR         => axi4_mm2s_mosi.ARADDR,
    S01_AXI_ARLEN          => axi4_mm2s_mosi.ARLEN,
    S01_AXI_ARSIZE         => axi4_mm2s_mosi.ARSIZE,
    S01_AXI_ARBURST        => axi4_mm2s_mosi.ARBURST,
    S01_AXI_ARLOCK         => '0',
    S01_AXI_ARCACHE        => axi4_mm2s_mosi.ARCACHE,
    S01_AXI_ARPROT         => axi4_mm2s_mosi.ARPROT,
    S01_AXI_ARQOS          => (others => '0'),
    S01_AXI_ARVALID        => axi4_mm2s_mosi.ARVALID,
    S01_AXI_ARREADY        => axi4_mm2s_miso.ARREADY,
    S01_AXI_RID            => open,
    S01_AXI_RDATA          => axi4_mm2s_miso.RDATA,
    S01_AXI_RRESP          => axi4_mm2s_miso.RRESP,
    S01_AXI_RLAST          => axi4_mm2s_miso.RLAST,
    S01_AXI_RVALID         => axi4_mm2s_miso.RVALID,
    S01_AXI_RREADY         => axi4_mm2s_mosi.RREADY,
    
   
    M00_AXI_ARESET_OUT_N   => m00_arestn_out,
    M00_AXI_ACLK           => m00_aclk,
    M00_AXI_AWID           => axi4_mig_mosi.awid,
    M00_AXI_AWADDR         => axi4_mig_mosi.AWADDR,
    M00_AXI_AWLEN          => axi4_mig_mosi.AWLEN,
    M00_AXI_AWSIZE         => axi4_mig_mosi.AWSIZE,
    M00_AXI_AWBURST        => axi4_mig_mosi.AWBURST,
    M00_AXI_AWLOCK         => axi4_mig_mosi.AWLOCK(0),
    M00_AXI_AWCACHE        => axi4_mig_mosi.AWCACHE,
    M00_AXI_AWPROT         => axi4_mig_mosi.AWPROT,
    M00_AXI_AWQOS          => open,
    M00_AXI_AWVALID        => axi4_mig_mosi.AWVALID,
    M00_AXI_AWREADY        => axi4_mig_miso.AWREADY,
    M00_AXI_WDATA          => axi4_mig_mosi.WDATA,
    M00_AXI_WSTRB          => axi4_mig_mosi.WSTRB,
    M00_AXI_WLAST          => axi4_mig_mosi.WLAST,
    M00_AXI_WVALID         => axi4_mig_mosi.WVALID,
    M00_AXI_WREADY         => axi4_mig_miso.WREADY,
    M00_AXI_BID            => axi4_mig_miso.bid,
    M00_AXI_BRESP          => axi4_mig_miso.BRESP,
    M00_AXI_BVALID         => axi4_mig_miso.BVALID,
    M00_AXI_BREADY         => axi4_mig_mosi.BREADY,
    M00_AXI_ARID           => axi4_mig_mosi.arid,
    M00_AXI_ARADDR         => axi4_mig_mosi.ARADDR,
    M00_AXI_ARLEN          => axi4_mig_mosi.ARLEN,
    M00_AXI_ARSIZE         => axi4_mig_mosi.ARSIZE,
    M00_AXI_ARBURST        => axi4_mig_mosi.ARBURST,
    M00_AXI_ARLOCK         => axi4_mig_mosi.ARLOCK(0),
    M00_AXI_ARCACHE        => axi4_mig_mosi.ARCACHE,
    M00_AXI_ARPROT         => axi4_mig_mosi.ARPROT,
    M00_AXI_ARQOS          => open,
    M00_AXI_ARVALID        => axi4_mig_mosi.ARVALID,
    M00_AXI_ARREADY        => axi4_mig_miso.ARREADY,
    M00_AXI_RID            => axi4_mig_miso.rid,
    M00_AXI_RDATA          => axi4_mig_miso.RDATA,
    M00_AXI_RRESP          => axi4_mig_miso.RRESP,
    M00_AXI_RLAST          => axi4_mig_miso.RLAST,
    M00_AXI_RVALID         => axi4_mig_miso.RVALID,
    M00_AXI_RREADY         => axi4_mig_mosi.RREADY
  );
end sim;