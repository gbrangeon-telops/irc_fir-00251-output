

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YqipQWc4JFBZb16rc2dodhguFDkilKhXXsYOnDVSNRAjtkaR6AZEesZX9P31kdm98GkKMNT69IgM
oU3B8PoxIg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Th08Wi4CTujjzYeFPRrbrk96/H9lqJHT1fOXWDhDkZaqyMx5/LmUZnPHzc9Mi1qiTcgVKZeTpkDd
lm04xNkvaFBlZ5KAxEqjMNmhtMTNyj98wbYe1WGtUEppm4URdSaGhgzD2gvskrJEfU0HoVjNKsYv
Y8g1ek6gYioQSqVo4Vk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3ST6h9XhpdCHj0//nno4AUPlABBr9tQ0cisrrim6ayZf3P6t8TzMqSxgV/q0TD5pBIm//qvgm7Bo
W2S1EUuvf2WqWkW7p/E9CPizeTTEZkAYHckCfZTDk/HTJdolSIFeCHjfZiRizq3RlOIw44CUEMSg
PXhJE4sbT53L+d0eIaNmJBJnZPN29vIw8LbE7t+Y1oivoLSh1BhWy3+lZNV30PrceJFjB3Ylx53O
r9RULlN7k4FVXKoCkEg9NcpjWNJAX4azHw+uuE/ZZmEDfyzXMbaQPIzErM+LylAQ/PYfvIwSeBK1
4Z1Yudv71r62qTHPKAu2JCMEmzvKCe8RAmGoeg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iNgef8JJ0zz53Cg6UsIY3rdr+PhJG3ZSgPvV55cmHG2d6Sfxzk8LG8+nTrPNPEPV7qefhOfs2qwO
LV1XGy8/zcDatxxl7RZSBTwjwXvbpgbJIb3oKBLjSbNQOSIIh7oK15z/NbQ04jpEoFW8I8unz0Dr
X8lH8UO/ss4o3sjSRmY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gdQRq0TszGQ1sYR2djmFoWhyazt+0Tw2kvNbiTEjaM08h64rXWx+KrfH4Ux19p4jnBVjDnfhSE44
xN7ehFd8XzCnm6T9eZgkCDf8dP3IGf2Nl73ZHXLjDsXHqpK6BXZEG/Ko8+LkLz9nw7Snn2cWezi5
seVqFQ9T1Cl73kL7otmtLUuX7sR7LkwbgtAzFivUF8Ml8V/izjdNdzsqpzxjHY9vo/n9JWZSxDHg
dF+BgQSeU0ooY6vwulhfUyi8hYLdbvSFz9Xlr9vUXABI71kCIOeJMQA6BrcWbYjoGqM7KNL6TTGp
K4Gc5G7xM4ucj70Vz377eDl1W3KXvVQRmQSA0w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6928)
`protect data_block
4cwReeA+SZy9w93k0fVK15sWKuDg9Ux5eLzy2pS5TP3+mPgkqOMcVRXIEIReVtBPiIdiHLvUWJvt
eqP2Ixf6J7+aSywd0EDM78DXopMy3ySOLCiJD77mDfiHsmn+IJNYyBWpALKGrgUg+Uv3BMY1+bsz
Szce0BEU4+tOU6lt55QyESIK92J8wvZxXlrqznvOBvuEVB2GfXWNbwhpzSoHqlo3m5XwQuOEM6FD
xQlpAVfGlMr+TbDnyyYHCgWCSIKtcjUPIS9LwmaSMtNyt0WIzE89zbjOPWu2kVg/kqvWfD6FKycE
lpt01AF13uCpq97gvI57Ce2cLt+7K/C6oKW7IG5yGH8kLED9Kx4AZc+pHoWRHDc/5ROqlimnDGb+
4naKw2cWQT7IAhhgOEKWRGaIYDwA/7e/Z0UAEIqG2YEfeR4H/0YJ249Dlz63JH0/oiQmn7QlcZHQ
boq0chwY0a4/r33QHeUWvvT2FuIvDLgw9egux6iIWdUAtdkjnK12OaVb6s+TVpzn2v8vBwsjlQqS
QYvl2TL1gcpMop8jCluK0bSEnpqjmIMZB077fT1OPd9Mc9gsgujA3ox8DnWG1pJDvUkgtqRY3yna
Mdymushl5eeFpBouI9iGfCGJ1xFlXDl8WF05ScVr1tJrBoY5/m6nRYdF3RFaXkCHUF7UG2/k4TKk
+lzJ4k1jAl9nM+vDAPNKRPYOUZc3dhBH8QgRejt7QRiGe72gdBX2dUTZiYRur+QYcdM45jm5r4CF
/h5DY2OKZcVIheEQJsG6HlAKV75pDpFT9Z4R56/eBOWabu8MHpGfc2j1XltpfJ5Trl/2GjoyvEC6
Gsy78NP8Hzdg2alyN88TVfkHj5dkqiEa97VJkjDyap2BSdajdRH02tFMeyOzZjrA+p/BRFqZw+3g
ur1xq0FbWcD+d7u1lH4KdfED2vMmfEJCHfny+eE+b8xX5rdDmfa27/V2SXXUdkFvW3r611WRhmE1
sdpL5GJTqUsQGw/J1+/NuJy3O30HJFJaNSGbEN5wfTYdg9eV1GvNHlpRVf8hoGmcSPZDdQpi6aE1
XNlibiAOkaklG85Wy5FdRCd9e7Y6wQ/nfst9GqvBcgbniX1uMhyHFxPDqLBbvNAcGAANlHCojNoa
yzqpw5nowzAvW8Qe424H12rEZ0+0MuBJ/Y8mRftAPkeJ8AvM36soMphKibNx8e/5MN/yXYdXg3Ex
gvYA3GeG0UXczzQfkaeOgWEINeF2xsnk+fVz4cg2sifBaSBeBeUh/4L6UuVHH6ZHGlkwMoOagvlg
ruQXSy/GJiMRjMgBuA8mGDlKvi2BcaFwVSPt2G5RJBa6DeLki+uZRb6sg6RRoqqWbFGP9uVuobuH
VtsOOFpt1sp/vQcQfmcBiyHvseBxR9E3lUGvCPc4Jap24s4QhdCbf4BNmqVHEvNF115T4wR98RK6
qsC8K/wTAgBvDVtTC1Kx7NieXx19w9Kt9f3ZPe/ai8ZouwmsIZZNmGfUzGkL0uJj2D2nR4KclX5g
KMQTuGX8IFTKmL7++nZcDVpGNg/i7D66yG9mhzbROv4LI/pH/39ZCMspy9SCkR1Yvtv8E0Ilge0Z
9fdbZLByP+jYZXLvd0m6CfGry0VitFI3O4xOVkplv7HAm4MkLVQicaCgQQNpxJG5UhkugyxV+ee1
GqoA67ZpmFo+bgqmfaVgbKtZFCvZvq288tyd6SYuxKNnA/TOGsQrM6hVBzp32U3f2q9ntcXS7e3V
nCEnNAePysgVj64tXic4ORR63MWdjehvnYQAQvibjTudT4uzlzaMbGSWgMGZYs3PYfHP4DwnEN29
QHPL0FdJWSKEW+PpYEbE4asIA1nNRALf2AXTeuQC3ZT+ZOH+e2wggAzXdJju5AwtP49dPiB73zap
RHTbNBn+a1QsYqoyRrtBrazz+bZkwSq46kynuets5i5GKQ2IOyNalSiyS6BKmjVa+FtgxVB2Wj0p
QLEXO7rBEoMbyemcaI1bVTZ9gGZx/fIv7n3znd6KnK7UQpIpRKNjupYteY/kiTe/KBdLf4jznpmX
8ZWjAEGWtX+1I7Ks7UWDAPiCeGcVosSjep5glaVkP6+5aMn5QSEaiIM7+jQnD70MicTfp3Cf+any
aX8GSXTXtoTG2lWBywrYiqsvSeazAlHkCI4SHS6Wox8LOGz/vVsFBKMIxo5j1rnez2FWnXkqHWs6
1P+Mb2AYqBaCqCM5Ks1atVkhCffrsd804GhMAgXOGjPCjea0zJ+cwe/9/HMJms+vPi2yAq2EzKye
xEDTGDMjTpX3bQH/IJBk2AEYYnAnFccVhsOpq+aCedp9zEm+HCL4OvZsDm5c+V0LyJcPxVi1/TVh
piL60Z902Q1RPlnJNDDFwbu+7kKX9yJkXKVanrONPYd4xn1lR26jC+oEjBT29L/JKix1VH4jy7HC
lboRfJlG8pmCK7f0s9uhuyGbXBMvTyrLyuug8cVauu0ChRnmKfVW+EPlwJyjoJIKt1l7rXmIdLho
gLPfggU0lTeDMwonNyJowFA+rppBoxndgBsK75VcbvdTzhyynYABRohPcRDN25KoIIc3meNblXpo
9+t3W1/ZP50gpDlIFIELnHflc/9oS31iMD2C1mpoEn96V5G5yTJpo19Rnovkjsq13vEj+YvaPD7q
ce+FKq6wupzcVG4or0Upuv0/w4i5jT7UCJCoctblbQNXpcsxMUp+ttQquhkR+sgp5DI05Xrg9G9N
e0DY2NBgo8t5J29SNKTAFNoIAVDPxeyneOulFv5Zdh6xD3a0Tp3oYxeUEcDxiQ6VRrQRYk/2pEpR
9WH6UP2wU01JQZTES0/8rNj3rV68jtlfbDApueah0uq8QyeVt7C3qcuqh/MTn77rF2+hS6ZhQIsr
iYgS3EBoOpEgJkRoPyKaIhs0NZGUV3MoCPzxGGShE5qVBeUiir20kAs+UOtU7w+SVMJs5qTUsY0H
YElk5OnQpGRQKXeke94iCQqwcX+AE0t+RwHibPHmkPiqiHKrjMRgAPKUKlcdS7YBSBzBFylkDZqI
AKZqHM3NNmQwn9nnabhk3NxzY6N2Mp1118o/mx2n1xq4SciWH6SqizvP6HJqD5B1KV1hdR7JYo5A
S5FftWyJlR2ISmapdhJ7V8pyynHOGd1NvUt9PKFBFhhPLJWtIH9v6OEnrWHFZyRvBfyCQ+LtWiGD
QkbHjNpw3oK5YTYC5R2knejDCr9OYEWTmeE+uFPqTmvXr89HehTas5ahx3M7WE31LmY2H4msgd8y
pI98M2utJJ1RcHbWh8a8V47YmmnVPnPG0EXzN343tAtn1LX3LxsMTmUVAldhahYmL3AI3i7/MnCJ
NQSkoInGM60jXP1Onsw1l1dw1HKB5P37igSiCuAxlzn6ZiEQryDdjK/D01Vkviw8SAkzA9ykY9Iz
28Qs22NhWB/pO7TCbhqQCJX8uzSrBF45mnEefaJ67uvhbDURmE2g6ErAAcAD5hP3L+ModZ5WYhn0
7hGgWmtUlLM5qsw7p/NPKdQB8DQvWLmDy9+QTErhFBu29EWRvaVlGSuuJady+L3/rRSPQ4AcQi2R
sIx/znn8dcHFjyg2I3itqFxceCRrjDVfFk+7r9Um3jbBWNSpBDYQyhdUe0ArbyDHp8e07duenMSK
kECRnxZyiszsNwDS9aGpk/O+dmZ9Y+8Rr4fbqjKHiHG/qzZEBowwU65emtiMmKsLCUuSNaNRP4rg
wQheHLCbETcZSELy5uDEYJNvglgzj4fqgIRg0ybk/cO97QV6oUEPRP78Kw1P2Z/ldtzFKI+10ZTy
dAwLZH8Vv6LR+7OEfogQGFzyV3WeuOe1GnIDSseXdm1fSFJ6q3fbGD7TIzANOeVZGTTGoqGqglVT
0WNgOmk0i4GiutlgnZ2DQC3TsXED8DzP86NG+V2UcQyiRC0SpcymI1dU+QF+04lWMNDt0ZLf8+aR
+YVWGovYgNlj1sYm8Ex3Qa3EU9+Ddla9qKOvsU3L61TMg70c5Wa6Erp1lPQv4byAgDyE1/xnVNPn
OW9MsNw62oHDwwWQsdAlRm81/nu2Ubi/0ajcKLdyoqDtad869IKtXxL3GB7VMRtT4Xi6U/bAHGb9
cf0SfA28irNsCQLe9JCiImZ8J1FuIynX2AZje+5nIxoZG4HZE1QJDIDVf16G4pKyXZXjlHQb6Vlb
nTFTSp6Ofz6NpDrVs3QLfwb8fQQ56HvQjmzrZMielsdebyDz1mRLzT/UoEcv0fD5lb8TYBON4jUp
D8hJKvShImjyVQ3A7Ia40AHFb3FbTAKdQI1C3tCepRwtn/id5/5WVAW82Vy9BmV9SeG+JYKHvfWL
jg6MUvF+U3CqFxj9CZkpc4UrnwrA2MVfq0oClQqKsIpGdBF5uZq5bqVN5Xhu2siz9XC1ur7AfZQG
oktZH93LuzZkXJrzSRy/9AtvbqyTwvlwoGZAOufjzba3zwVjgMleC8t56dz2/1/cb9VK+5LN0bSp
jH256E4onByUiirB9b3Q+Gky9dw914FBoyg8N5mmHmRPykjXN+5UVwMAcKBaaQJ3qT0gWg3kRThi
1epa4e4tB7cwy/QQHeciH1K7g9vN872Ubx1iDPwJMZdVZPt2W2iN/AUIziPl4rGlZF10e0OKRzaz
Ud/zICha1YPOP0WSY7ZFW3TaiO8XhjUV7ktUj4HmLkqy9KDFf5JwDc1mPArIhD3z6QaWgbmjrbGT
bCCGDbIoxYxPi334FpqJZ+zGcE/ja8OntMJc8NiCNZa9QkEag2oUdShTgEMEWDAgoX1rZZtHslBA
H/v7n/6ZX7h61Nh/b9mr2i9lkSOitVy09PL40nNuYedEEPP4J6WkZ2AcyjROudgOH3u0A+wo+Dqp
3gFn4af0oh63xOxzCFfpvI9RE1AN/mMEBEefG+XAc9Rg1v0WNlzKXm29kyIk82q+pFeNn/0Lqzql
83D2kXidJ9bHvzFz7QwRF8IF+pEjPIdtUtOPfz1Ia+2HWcMgJqa1Sm3zJuCCYAVHwdXWzud+g9A/
9AuuSUf1pdQ4Q1+VSPxNATTb8PNqtCm+XqWSK4ctomuVJb7XF/5wslXowQ87UrE8JzXIEuNjXMqo
FIk95UAaBrwXozCqfQCR8qCaDEUd3FHrazvuZrQSPeRGta13srPl0pNvz8aU3naYOSmPdgd0mkVc
n0eqmOv293aawem6ExxRSQeXcBZr2q3fgjbgZ7SaCfBNWW191TR9+nqSMihMUTVJae0Sv85xBn5O
SMcWoLpKfZDaUatCqswbyEB6xae/7dlzdm4zZ9NafSTdz39otbW6HhhiuKE4NlRAdHSz8W+f/BLB
PR5d0iqhYyvlix5P0fgsIChp9Cmm4XCjSZAV9X9BeFdK5M5AttiuZM859pppAaXXMvVs+HM+sf6O
4KB7X/koOW64fpQUlQjRqiPHrs8xUiy5Mhw3KhiweuEnsv7DO+ZwDwvEpusdjxdnizenyMuUJ0wj
ySU/x9jHPLU5x4VIk60tnz2U04lTlp/RWr2GXliPq71rbYuXxTVIegJuVDBJEZwTQF5yMa5QDhlf
oK5PMjjCww/QAi4rFBZE+hKS6vcKft9k2/jspb+HTgToNnt4vnl7mJd84hhzvmg/Tj8VDu10eJRt
7FWuFsj+sh1gCwaMIEOYym47ijmu8NnwhUzWVU48J6m8u3mMlz955+Y60i3bguEx8Icbyb5uKLi0
xYMuzUays53n6WxReAVNIDeqsCPiWjunyDPyLb4+Eu96eLonjxTL2gtW4XKFrGCugsWT1KXEiOzV
CQZTl4t2cFwdDTr4xwXye8DtuCW1wmKcs5rqi5lpZi8M7PxLVDGcsJRdGbEsaxeN6UT6B8KMx0YA
sYNHTxHtgYRDMJ9IEjmXXhbt4oueVByh2u71r7zeHPqgJh2mPTMuPvO1OAvnLlLxfvnyEyivcbBV
CXRNJuJaW2EUo/y85uFtCTdLa0vZKx/eoT37d8af9Z51OosRdwFHKOUB3xT/Xm76sPoaGpmmnM/h
aeaZ6USvc7cCI2YtaexF+2dVOj1Edv3Y8KfegNQoatf83xOzJgvKL7lr7eJ3lh92uEpKlkGCjUNc
dhhkK+/qB3Q7f8bRkHsopQ/kj685FsGxNLV9biICH64eqLCmh38mugrQt1TUrSlrHjwKSELbSyFm
yce70wNs5mXljEZ0NTWu8kEIJJ0vGDCGHBdjk2GmfBJbtDaspmGQo5swCmLxKlaMQQP8rxnCFlhc
6fcf+cFm/Qubva5BrJoHZIpzARoWMuvzU/JB640jCVaq9j2HYLXJznA81S5noSVaeWHClp6e2Eg3
NWcjV47awN/8LkFWEBI0ooQPTHGMLkPENnSuafkFj4YNBKscwQliiEYWhqVUK8+ZZ5DvD4Oko4jg
W5W8rZoKUcVxUce/5Zy+7rxtZUuTBr0e7t4Vyifu+hCRPbGWGt8ClYQbaTmmfvBJqZIQBRQwuUKG
B1KMLcCNENl1QJoxscSWChDIOXC9xIiJNBPefBB0WkZCwcpy1N2f6BUPIefwkzIKQnpQelEXQO/w
kCoyewqUnE7IEo02166H/t9N2ESk97DuvMQe91smjFl3QatexPnOv+Kq2lRCKbmnzrCrQRg5ocqp
P+H7TEnh3Cit6Ev3p0DMtqgy1gW+AHTpYn6K4RJzQKA3RWG4EcRsKPtoA1iJwaJCLnmFWjgvL+RF
UVvdYq7fPVFTMCasVI00MUqjnXiudOGrf9qWbKtVuZhYePopR+Gttrbm2+QIWpUMtcFcz48z+xBM
0Eu89ak4pnE2VONIrTpLrzQP75LZzWgyVz3wzot8vr6EIZjiU5Q46OMF/K/EkVz2OacwvZaAEtWY
NUau2QazagMQkZVBMKs4mhcnLZnuEDQ6KHk3KWfZp8+9Vu7+3UyfCdXXudLHuCZ0C4+yyz6u/RkH
JyBwnN1w4wAIfuYD/S1jUO6qlqwd19R6GqsTLagI4i62XTIZbqqH1A7wWT3T7UM+M/TSNP/Q1jHw
KVa7wx3b86WaMJE3Ah2EqqHD7vFFxJAkZGVGCiRV4qyOhGzH/pwFr1G+wMSaoiYolmz9T/czDU9L
gD28UMcuDRkc+GDKop1O6vKyjrpeBfzVxAxejMv7SZBSrPL47h/kr7dgsf7DHkd6KtM6BGlGrHX0
UFlWDQbpjdmQvn+bVBLA5HyBuHfZ67PnCaWk2bYSSmjOJcVS0prDbFuUghEK0N3P+WcAw5bblcFX
ghOxMWl5ySkgCridC32wukHYY+fyjCp92DYCSsf5g5fNogPfE0qCj3e+wVZb7dGcJfRCLqVxDZCw
OseQeQtIVpGPuYW+2SnibiFhTHP/XN5Uj0SFjIW7EulwYeHnhKYPYKuYzIbPYCmCxcRc3DxiLikq
7AgLqpqAvMkjPgx6nDRTAG4ZCFtTKVYYoDhErdi06b2VHsTJpWoS7eUUD1ULilM/aNniiS+T6Kgf
6ij5qnOz4Syz7qrUMEqzvNaaWrf+ZCp04RbMVRC3OOfUuncJS7iqRT03THMxzw6MqZSE81MbuJKn
jP/FU9q75eRZDHZTEuMCdu+3uOAlfqvnQ6JbGHnMxaLSBu0b9PfvScERXjW21hK4+btfOReH90kq
26ereHlvsObI64kuj5zERS1FWTIQjs0JTXeWrPim+IrntulJJTEqxIg+OLCWEgQR+ARRUWfUVcUn
UO9ckLiuXngAukvUWW7N3n2Ehuo5Ht+Anrv9FXzYjAkOgHzFBhjQDsNvNRDJL+NXWZPYsc7EJdNZ
JUtRtoVCamTuPcpoz3dhmmkmpD1sjZnOzzA24rmW94fITmmI3CLYXBra/mTsJB3zVn5Hze27+Ia1
8O0DDrVb2PieRSsxyCoTVLJWKYNSy5UWFj+WGJ7OxIO1lPY+1Ta5q3CGbIHsmVrPi6wp4fLeZROn
hTiC5xMIJBnI998pZktbkiejVVw3BVTXficCBtYTIfJuiWM/nSnpjL+/KJZCZbc4xz6kCtCU97BZ
LbMW2nHZirX2pOU3JWhmGYClv82kBgyDS9kppGj2x69jrGtWQQnLe8jws0xtTBefnft8s0ZDJ1bb
O55NLlawH9onQawycUOsa3mqIuky92SB/MKhH6GFFMFVSk5Io/vQSlctY7e++3CChm541ga6svht
4LRNam8PdxWhL4xg84RkRvtiWGFIk02gyrLxfZNCXJMI26zo+bVijxYxEY8MJQ8If7uYlUpsjAvS
F3S75MwLMv60HydOhl/QrCxBuRuvD6FAglOVqornojX4ZXjJrKdnCvMLnCCpSYzhjPJCmoFXu4+Z
fXwS33uucIR8cjz75VtAXZ1DRgCb5tS3/cEZFVLbyYdcKNAFQIqasddFDYfe1nfT5gU5ZCpCWKs9
aFCWAf2CgMESUVmSJOI4OSazqwvSl4lNSLv+DfGeObav+NpCIn2b5wwgbroZX1mvFoRlQv3UtWUV
U5loMshFkvK4XwV/7m5B2UQI/sbP1w/OJ2nndMEp234S8PuCK+gBLs08WgJQbWf4UYEXa/yu4aXj
YaSV1sJZYRpSkoUocr4LxbBC5ixXfLYkfE270/bOfFJMfKbu4UjB8i74fm7MRYUpShJztF3EbKnE
c4Ld5szcjl5XbP28YNEtd/t7rwI9+1kcUOpoVDInh9uHce8ro7hVb0xPApC25FrPD3A54RG6tyS6
497AB3XowM2GjZUS7HINaq03MwKMSeBgv9aQ4XusbQW8tNBtWX8hISEqtdEI3LQ8tv8VuTRdIqNs
LLJhviKVbdkFslr/b+Wkw2HbpbSYXnwDrYOcOpNzspoGKh+pFOrD2sJ8b8CxDXGERslZPiHg6c6I
ylZE1sSPGupiM5G7DOjks18dWATm5AfBv4//dM+jvPQ9SIYdPcg59XdjklLjaKwklFF6IpnWbRsY
jG/DaktW0voTVtEUfhbm5Q6iDhImpypNGVsqBa/k+TcrBQt2OFzuLO0c6ex+BKzJuWffEwpN9d3I
Rfjef2gEz/GlQavnKaFrFyiqUX9xcD1ntFJ42pBcVxJ/NZVlWui0Obd5qwCgZC3jy11jJPe/ps5f
/SjYDQd1jTXjfr3BDeB9RYgytyh7N/Q8GJgKvJUcWBu9cdYJLbAdLEpPLl8FUP73322FWIJ5POPe
fovmm+j0dXpi2YXKwCdCSZoXf9TZXM3FDEnFZhgjA4d8cvqlBRAP+susin6uMW5r1YATIO4Dg/fE
9FNpiOLgcacqFQ9qQK6l00knPysdAHBVRrvLje6NBA==
`protect end_protected

