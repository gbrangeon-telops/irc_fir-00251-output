

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OHeaBmhw2WWXga/8pOVTMIzcYutI6Mhna2kzvZmeKvttg8GRcsMBDXpogvkdmdxp1KLLzWXMAKSV
fUAOBPVAvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ao3tKAmGrk9jDIJ5tmEl5p3MIRphIc7Vg/SqO4TER/rFDRMS3J83CwQ2b9YFrnde65FSvizCvsTV
0Knxkw8zoIma+TSgIxOnivhI3WBhgKeA2uGkUI4h7aI3JKyXt+ar8rATgfMIjtkwwZmXnAQdFAm/
DhnKD9KmESp1ihQZWxM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tIRCJBwrqw861TllYkYZisN+3Hf+P2JXRGH4rS3/mIyKaeRa8ciKvXh+DuDwE0CQ8FK1JKt0o7Wy
5niCab0pNdgMIWoeJTN4M3Yv3mIYHhxe/uhUY+qL9dbTdi1peu0ypGwB+pCVAaCMnYsMP87ovoxG
mFxz/aWHoq6z5hUiOqs/8QctFGTu5uGrqo/fDpwnQByfUDzc5kOGUXom+7Ix+u0CBnUzxUPMVE8H
FW15FWlEhZ2/WOv5odw8POvTaQir1St/I4TCBaM8Ne779Z1F4E4v1nyrImWHcYGt30Ex/kdASWup
x0rIb4g/F4zfpMwk2F9PI0IRzfsxsXBx1PSZmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vDR9iZfmcKoc03DxzsUkjAUcoXZpLGp+jz9oB+bhIzk9fA1B+YkBJ4B6wGhxOSVsIGzj0A/2+sve
cYv4/y/PnMWoVJu5GAXMXsNWS0+yhRlFm65eqZTnif9T4BQLUfDB3Poe8t8+8qJraoiNha1dShh9
FtnafnjfaWlgFCK4DSo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5OVsGiC3k02pbA8zjICborh5BXFBySD3cMhIIsNr8DZdx+UrjbiVbqZMU9Ry3hJ/1iX0Q8zDyFo
F6W3nmvV82n8xeQJN36fxUpz69izOLDYVC7B/XqC5I6fwrewIKThxTuK9lZtFdQHHrzj3T2ZDLDy
Z1+PK2wQ4cNjjft1DSS07aO+6gcWXb8X25cWmNGk/P6Hl0pzIcfFFHwO6Oq+bJ671kKmsX3jUKAg
DTTCgxx1Ex2XG0j8cWCnhZjmetyd9o4fKBdb10goxmIXB8/8Sn+4BcUJVLUQkMnRwy0YJGGtpiHs
ZxxUU5IU2sy5csUBb6rGbP4ap8jLGVFhtMQgiA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16944)
`protect data_block
ggCzI4dARKq5CbRn5oUhMybfQOSAA27V331WBo+FnK9/m98MJmw+ADQ4x7k0s+Hq/1ZbMRySJ4xP
dgmlYWGWABwbmxjISpvetmRIG1h1aEnbEB/jdM+n9bf6C6iDJsiOwuaV900S+jVp2dDrosLPGN/k
50Zd0ZC0f1CJ2FnqAKnvUiXQbTb44cuThCz6NOkw/onl/ibC1tqyitOeSgKKrxm5wXH3pcrtemHP
M3hPsCxVDAarzKi8FtdpgaLvxfSuUbY7AeICxWvEyeU3yGUF520lYriw87S0NiPTZNUl73+67DJT
qRE4hmIcM7IYIdDz7QaleCwp8E5w01CMkdL17/yz8OemVa6WSELaMGjT4i2u+1SBw1j4ZtjHG9OC
a1EA5YVi3c9RcAOWsuNNotIocYHy+lNkx+gsPbTiy9BBu1ByrXVHB6CYbeOjvbmhh+ov0R9EGnmr
pPgzQsk5xH2GcDNmx3SR3/2MIaJJHM9SUOz2knMNtXCThitYT5M7cq/YxAZ5t/FG6rTJct8+Honb
Oo2Ch5Ms7o3rdj5GWbSk/dDxcE81XiWVdLoZMnYexAHXaep044BNAxXHKZbw4Dftqp92t0wc8Sfm
b4Q4Zqoyy55EOZB3dIVyYx4bz/rZR9Eu5dSLV+OZproXzcl38l3f7Jo4GVFb3nrrSmoEtJi7xiLZ
vJwvvJrcHetNpg1wqe3nNW9A7CgyTcgxOsmTmVLwHckaycRJyo/YZDYBT5HfnbPZmckyEmqNhHI0
nyymujep2wczHqeYYGJieqz6UrASh6W2cStnyW2RfXKJO8/KeGvkSRofPwMgFw6wJF2BdFPxb0vH
Vmh6Y8vrg1DWOiO/wBg6SPJO42lxRTvnbRkk8ppQZy0mPjDwcrF1iHWo5FjZ9p4iS8ddFhJHgSHs
ku34IuV3arAvm3yhmlTwcoky+vq380gXzLK4ujqjf9ZifE5waYlIEVTR09ZwlKriry8T9Rio0AHZ
EZ8CMR4KGgS2VYp7EeIDccpJdmgZjz4AxhZ4XExZknLO1JSebaOuxNkRfOFDf4AdGYWOgQHEKVDC
MjmN8KVSsQUcjAjcITOVGqPm6wlCVpFZIGjquwPNi/J6Nw4Pue4EumEiXF455T3ojB5sMSiX+Age
uXYV41JTo/4wuCkQWS0G1ijWdYnQYzPU8I6YcekPox3ffaVZ0khs94zWft6ty8exlvLzX9ECITQs
dqbhApB+V5UO6ijpTeTwSACp24fT+7juznsyEZaA+H/JxsVxUseUCDZfSXbXf9IOuIITf41ULtJQ
obXxN6HvlUd1kVicMDSFWxfjYnS3H2y3xzCp4JYrCn8tjnNzfIgPd3u9IJLiTM4fw9bHJEV+iacB
gAw8A5FGJzvaoFSdZSAdFQLiV9cvHBAqm96RabYWz86VH9Ba00w8zLRc/iU81WNNNpkC3UvRg8wO
Cg/FncH3Kbqg4VmD0elqtkkSianqQRT/V5grTUaGn/ev50nATlB25/2H3+pK1LBtGjMarJKACfBG
X8kVf0lpdgZYheJgBsoYeGastgr8Bc1sPIoLLhC873V1l+Pc0aJbnIaHvMa/d17nfBDU1ECxTAhq
JiJMh1R6xaJT0HP5UtNpD/H4L3siKb3JZ3NbgdbDrJnA0cTRaXmuSqAqlumwRUM7h0HcvchhVeYr
so1vcu0bBf4tfk9/Utj5OBDVaMHmmK8iOm14lQbc0AsFdvWVnPG6huQsYxKfm9z/5QdnRrNdd73M
T9mma0rG4bEbR9AwkRVejE+dbVxIvAD+UA4oTp2IKyfwYIJxKCIzU6xzaL+N8REH3o+wLuvM3Z3q
RSyMsVXnwsxbXIbX3HroGXg3x3ztOkJwhL1FiLQJoJioUInRauGck1VZHmpoC10L9McpClIrZ3Lv
6AlVNZglSCUlEaJ976nnF8fjsrRqBbwUkoMxfhNzBIKKTxLUjFWrSq7Nu0uy6oshrBkvpL+fQYhP
B8yEqCeBdmmicXuFUmStfgGmcoWKFhF+MdlkyRV56aWT7/SdQPH6u1qtVgoIQgGi4n2LApKV8PRF
l3k+85XqFEPV19cebGUdWtI2xxnDQDiqXgHoVx+5D+wuZTFXJzpWo5WN1gpTghZC21wgVehmWNL/
GuCBi0eMX/6XSmkcFSwI1uUQ8ywikokWKwhugOKlHcVedKxbc7+i3ctDT/BPXaqpTW1zFJsVOaYA
vHlF1S7+IcIxQUpbPWhEiRkm5x+uqfCwY6pImVrXjjL+Ee0CDijEPZD5mGXIoY0EqxGFCN6kE5NK
HPPqRFcWziOVfviDUgvuxMPOWw6pXPgEzAe37ezf3dDY7DzCgd5dnt65KoFJ6PAitWgDeqH9JWZC
MsBFlhW/pPkjQGDyg3ovtzSRySrKUpCogRvmE8bNF7PSk9pojwHCONO61Nf4mNlal5vcDKvT7O/y
42vq8/iIWcqC1f7a+QYRdmk0SMyKLZZxlUf8bq09Q9THNqN+EqN299edhmvagXyfPZFtp9roLHoE
fuGL9NLvDyBUg8YY0pojXtFpfiBgIGhbjNfUwta7kPaLfU98rT+7+K/ujfugf16lT+N+yxoNLvDZ
7NLsnh8HAWNAvG817OO7a56vrprphQs0Hh1LPapkL/vGPWk7Za6FdurvBZzEY6dRWjyBeDft0wDX
5YdrAqi1TwrhUsi2lKDIoQszVdbWlg15SfrrG7+tzFP6d4cmdMf6yp7SfwERE5HFgOQu8Ul/Ctog
iCm91zPdxf8NJ2Eg5pRVMT9a/73N6L9fhhEAHcdHb6A9GJwlYRmMW3zPVPIRmGOEoP9lTGU8Co8i
/9n2lLzCshiLyEK9JeFP3mB+QiDg3DbVaBteBjmMUU2W5gzzc3VavVrvEzu3zwY9f+YOs6AIp4Dm
oXu1ma20b72XNJbjULb7N/NAyGIKnHNvWpG2lt6dOEEFqKgk7Tl/X87oHXz81j5sGcVKJ2ctVL0Y
kBJh+EkRT4+DSUlXRBo15AP3quAUccJWKJ04D2uFTt5Botluv+vLKa26hAskT5mEiTmBO1nlP/ME
pfF7pCaNXmsBmBpHhO5gEw0xmOihgNhXJxKpxrpWdsGGIZmjsfr+O+5t0Xut5H41rvXU6TN4vVL3
iBay+VC/KXJN9H9pOU4QRAAgE5508Ah3nXTmWgVlCkjAggnUhTyQ/YR2hJWiWDI/gRMYZGw0ir4j
G5ABFSe6ssP7w+KwuElr09YuBogqoKqqE+diG5QHkLJoEutte+pQ2ffylILD1sTlrvxrbwA0jQIz
lxbnJU0NFicZhyw1tWS8YtX3sbcI4Xz3aHequGDtp3ITaaLqrnFElaQ86pOvjRU1TLfr3fKHI/iT
K5uuZMtgGfige5PYmKZiweSIbJUbHYm7SG+ft3dhGyQbwbXSPMt9ZMslZi1VjW3rX97ef+jsVRLF
j/Ecd4cWFitIqF7S+1QJvu6/YU3Zgm+L6hgU5Sn3EIT3zCMzuLOsmNydLRFA3eg4CeAg6H+nHSgH
u9V9RJ5P5Ddmm+e2+cGvL07hY5nzQUSFXCOU0MFjkpq2l4qEskl7ODgQPa48fsV5uHJppSo9JUO+
1R8hXgktrNCqb/+EWcm7j1IlL1oC7buNJjh03GRrQb6YMhmvYs2UZWN9rYkBEr0tfk/B4y0oFbYN
jatZcSrskIj35cC3cgIHgl8XzEYK/XvXWMEgznWsxcnJtK34tmTg5kGA37dhkz38I47bMPCbF71+
b/ltOBSJEWAnKgkyDRQi7GILIFJCJGH6KWhuxV836gte4P04J1K8RTlSb7gaMvtHtciRmp6NRLes
aLFy2mx7UkIMHB5zWI6nhSXtE+cWM8emFfj5X/vlMswInwF9iUl9DrbmhTbYpPogMLZBTuKDZP+3
SESm+umXLC+etOLY1XD86jcjl2BOzwMSZUxBt5V2pKH52wFtRGvzMEzaTdxIw+8yncmNsBS5TAJc
vjzjqpfn5GPha5wQoJ5QWJixZkK4oECD/XhoZ9dBnqC7omX8rCSCMvjOjCcWlI/f+CK+Zj901q91
l55Cga6KmNyp5evhIYWtHuMwDmTA6JLGfTa/V8z7bGFlTh71DzHg3hlNxdUncF3Te9Zh80WTPPic
7CugtA5JjVxp3y5nCRnaphqPWmP0sdkxiT85E48aC2SWRywR5T6RCUWjN0f+/EmgdKs5KtNrR9AC
dxofGPgiMAu7ZvfH2P75LHq/l1zIdJpf69miuZdUUGcCYpWKQDaegvuwdzC5kn6BThDAxTRktX0t
dK9k4h3arxOiJxN3OxABapYIOmN+pRosPup9mqbIZMiPoNzU3Xpym1sO+B9eAm/Gtg8+CfbNaXnx
TN/ZQnN2l2hFbJ5+IaBMmjw00AKCEOOy/a2YQosUTIpv+zq3jIwpax2quBZrfctWMjQ/jn9mt59b
HopfHOO4KXVu4jYK9J8WIZWDiQtYaT5oZAuhWnE7+Mc+h8tPeedvx9toxC7oG0Chr40B/itOrAeP
31AoPrWJX3F23s7MpQZyyQV2dCLx/0ThrObHHh46bg7dYl45r4Z6WlWk1KjMZOmkTUoyoRF+/wYA
0+dMWACTSBj/hfNyLn2DQINJ2g2PwGtC7nAPezr5JS7WuNqiIu/xLBSB6gic9URe2Yl+yFDCYJMZ
NDFysoT9RjoO2fYf8Nqc6FzAMT9dOV6iGqz8i0JiFTdC44DUDQYVPdcUFKpxO8B04/lcvyminrFb
lsIMN4M231pKtGufbszi6UGg1l4dOeRmhM6UCuCgvuqqODmk0knG3jXGfGzqn9uAaZ4amXQ4IDmC
sQ3G6uvCIhQm47tyNAg6X/E5c1vQLVIA1UhLbl6X6AysYLwDbndn+/13+991Bhpj1t+uPXDTvdsJ
YNiTKUsHtz/x/jKMykWOeufCNsua7KfLpXnRChH9Dsl619tTTy5Ff5iBHQRP+ww1SF9lj94+XFv/
TN0IK4Zh+UBfjWkTjyzDKLnAM7Yf75a4K/B9SnCFKauedEffGKslaEOJhV4pTPnRymNvUQN6F4bQ
ikJe3cfVm3lL1cen8B35xQos8Yfv+N6s0UHYeXW9bzxstppU+Va/jn3pYu6lNNXdyLGGR3FsBWf1
ovgPqdg9BtrlFfLNg0gXlr1rJkeg9Ucd6LQWaZ2CE3HURrOK0oifW61e8NIuC/j2svcpeN945m8Y
7aD0h7/e36fJ2T4tAo3xzdRAsxtwTxx0r7UOsjNz9+MAFR17HLRulJLnk7ONhzM8cYsJNshS8e6o
UZATJb87WbscnZoyKWinn7UvQ/NuHohPY9H6h1k2RFve+5LrB52DzLAvcJqyVDeO2jgbF7SUM922
dltOE5Y7+bHYM/Ab0t0Iexmx0n3BhtLw+1UNEecCGKT3nCp/leKSd40tvmCvtElh2WNvRJeaLgW2
0TUn58WcI7N2xgZ8U45+xXEaMmJtFG+8zn7+s/PtEMiDXhxkvl/SBrrI1KnuXj1Ig+9tUlxG5k+P
GvkVaYIOlrRsqK9cjBS7CpzTKQD9tZyJ2t0H+wFPQeGpGsjGs32BN5r25u+rBkkeTIRE3mSDbcgs
AUuiZ/cmzQdmoSQ20SOfKrnABkMR4cwLgieCvK1vtKoTTmjzXOBbH1zkz8zqPGqcRpPDhyCXWpyl
c9jys68LKCATL/4+6ABJNaeptKk1CKaVHecfGdQE9Le1sCb54KDQhE8O6h90Rv2PCJff1OX0RTja
YfPubzihUZ7r7EQJuGmFWR5amFrDCzIvTBeljtWFp+V1b/7G3j5p3ayIKiYBjNCKiFMdgFQvbUa+
xGP+ssvnvcv8yHTVg8eOYosW8+P8+t2RcyeC1pJt/0aSkbM+vuV37BS2fncO7zQbtIEKfOrX/6z9
CFb+5O5/HZK8JcVDjSn+g7njH7nOgnEZj/a+F9F0/umRqSXp/4x83j5+iLDoS+T2DUbAa9NU5Vq7
lTvqQqOGLwCuaf/UBVoarBgnBb2ZiP+wXBX7XSRdq0vgITQ5nuYGSYzDJn8mKUIFxWZ9zUTyVWNF
F7Z5/QwWmnohG7trenYZ0nglzaB0SdKFW3BMFY1qWYD/RDrORVemfAXRFzBwEl0BPLdNICfBZi6G
o/rrbGkh0tt04DhiYXOUyn2oMOQ0NBSn5It2f1wq05DWFX829RvJl5tuZU3OjZgrz049jtZ3PxdQ
rGlJgburZ8g5LhdL80mY8bmUm+lwqBGJ1YBXNlNLUyJ5NqM6rvilD3B9OVzEaiqaU4rBNDkajapD
YQd2oHSL4pmxhRZid/xFs1E6ych28SZFZJ7gVJ4a4btJhU0HMX9l3NYHHdV07/zi7DYGCDYz17ct
d/N7H5lnY/WrO4VTLr4j3q7ta31QMmsEppqew/G50m99WqkdEPt3xToLKuCI5T0QRR6p8lvBJVS0
NhlHUhcYK3GnY5ea5P1X+1UKGTcW+PBTlYQLZTRHnsEAvaS/oF5sJLKxkUh7XEcwxTYDpPtoyZ/+
Bb+whFEZ6Zhz4RWd/lSsPG7KOc2cUKQrGv74hd8UHXQc/BXWMfOz92bIU5GPFgMpzt0BxPYqd8NP
BxVbdvq2e8aBsbGylXSSzOGlIbWkspmYaGj++Nwh0ZX9/Kds1jOawzEme4/ZbeSqEuCsipMohIHM
+0lXmsA790vYmSr9OFefNWZeu/LLJRGHcQrqx+xxt2SPswcHhSgZC2V4aKnQmQIzdFKmB62cibnp
37mTjhXwbTUSXj4idKqqnWEsrdz58zemrzqrxYeUYiuqW9PZ8E0hggHPKjiNgRkAErPDNgN1q3qk
GlbecFkSdY10H82CR5tUXSP5yQcgrbZ7H1lPe5DfExpVv3lJ2iy418d6xmCA8kWrnaLSF5hB16bO
PBdB0BPqVcx5dnYZKxxN27R1c+tkDyymIdgNI1TCzNmx/BiliTSCUMdDMIaoktMAPTAgeIF0vglD
vSdM9QaX5OcSaJM9yKkJ5DJfjufp4PBsFZhEYt+ezpMDVKwff7+h6pRpN3JtCDES5EXHCBvjHmao
gcifQSydV6hP7tDk/rbVSA6bAbdqI/A8aKzdoJ5c5wziqSBLdNd1/SPr7ixpH52kvGAEYvISanx/
B62PEDE1REAKGTCFy/vCwo4nyC0DotAKscDzAwJtANt0CLV/u7johLAo55IVp9D5zAPQ5cgU2dHN
CvA/XtVN5HOzlXdwRfqovSAN8/ygt0d9011v6xa13pa/GcuPeDPBVLCCnKnkhr2Gk2Nj2HTxuTub
FWch7qDmMdI2ZrszxxJBKdi3nXbXwgswUOw/2Bt17HAcKmD8NMLCzRXJV77Y6Wyqo3LYsMgdQyRO
2kT6rmi3Z5zdUxC3Ogd+fYXy9EecEplyX2zoCPYkzf0qLygnO3PpCQ7kvFCHHpcyfnExvPiE/tho
M1jQj+ROXg7DXaTBxpPv/2SO6LSFOwa51DoMifIsh7HI7kO2Ca9PS1vBEwDyYkYBsGlBKU5OMcUT
ZrXhXgja4scfwXFDYVGbdmCVbuN404ba0tcmDHeslQBHAMvk30e7Vh/Cn+g+EqhZEdvIJ1SIwQQ5
qP/m6wRS7QJk5yy2/F3AqoqDZ2iN0O4uNIxLIjPpuoi0lRzSwN0VMRsC7yUTXSos2O9QBd6m93rh
Oo83W8seoRPCM9IH6MLvJQs7csLarF2hy2VoL7idOOV7LZ+i6kCpfjw7UOueNizQ3APBEKRxSY6Z
07f9YF0e5iGB/dvY8gsgTiqwhK4CZkSYBaYe1SvGyMOp8QCQwL7cwzVwuS+Z7K8dk46RKOKCfmvc
h1XgcnTSOXcUJhibZibYWnyhNVuCZt5WzsBZKpCNQb6lwKmSTcSnfE5NL0TE/CHJSXcuFCjmSJX8
0juJeq7+JvHPH/IDXGEYIJBJHChNLQ+rn2hnegZlyyL6zBXSjnjtBcWMirfio8oDEQ4WbNLEzlZL
qurIZVg3gMnoGicHXF2ttnJcJiPUFAR5GssCJzcZVIlq0+E/JOTpgSLAKcsWuUfhaSGJu36qsCPg
D9wGLK/bqnl71GekTrTQ6+xZssmHV6SLbCdvDmHZU9HxDH789zEIFVEimkhTZzgJTg5mbHxTFZ1x
jbGiFvcfQYTBdrtMgSn8TPXQvbJw79mIUDN3HahZPlfDT6W/KW1+mgiCh5O0V+PG+nDHEkfx1MqC
8WoggOAD1VIji9whBsgym80Mpq+SxiCOfbPqXqf67cH0WfmEMM2VezHiOHPziHvsYbiTV1Jyhnu6
0avPK8OA/3qE9IpkydSV1FDlYMBE4OzLhnRyCYez9gGhxqXCogre3cr1zyF7RViig6YCTvWkLRXx
0YJv8yRBWth1g3JcfAngrqmNCsGmQHOPgslB3Q7gzv+IAcXs/E50J722tLVsSN82Sh3YgkNyR7cu
KGv6CqAs+iUZT6YByLntysSfRorL/fST2kbdYnUFM9k7BIWw9Mzx7ZGtNVioUoFOnSD3fdLqPgKa
fQZQpV+Riqx5jBv+PwsCKoc9b9EGspmf5h0mvI9Pjnzki6m7REsBuFh8b7LEoMN43OBnV2xZV2Dx
6/WFCtjDW4w5vkqyKRJCcnCLtxlAvplgI0aiFO44urs3npyFOsr6svQ4ySCYIYEPuW/I5YFtN0Fu
XSPdpIr83rQKAVMrTHvsjKk5fKfMH/hTeXREU6rRLK1DFjrKQiRIDxZQadkFwvqXXiiFbSR9WmkI
BZAO2KB5uF4AiEJDKfK0hsjRRHHIEX1E6qcmP11A5t+MSpWc0QFk9mNr3neONdeG/LH8VS0cUW+z
cc2lPS2RM6z0YjnynlUovYc4SKO+VIANR5BIpfEEQab27qmxv+gkeEHhxPprhffX69UhevJTFqi/
Au3YZqGUGpWuo8qBzRJ5W+osKJkAq9cz0ujN5ybRwSypa8AsYqOjVklEGt+GnhF/aF4Avc2cFRDt
kZb2DqjnwhFDNWinaDZltdq+GXP+PJB76IJiIVIaRWI3AA5QWO4z4aHbbOP12UnKVzD6IG582sS7
+ENUatLeaxv85tpJXJhQ/Lz8UVIQGL0cVGe3U0yCE6WsBZ+GWV36wV32/DSmpPG1OH9QfMc/CiCG
JhCxnb0dseUutUPOWN2B/bvBC7bZoZ8KDoBKVTUjw7qeiHQ3LJeiL48yHnDVDhXBNruK70jiFaFX
Q5F/t+AfDtd3hAL6jGaDrU8QSx8LYxJCe+iUqP9vij5eundZT3P1Ym2UdAm2PdnMjkPIWavu0nTh
kF0C4DlnNmbFUO1qWVMx/34nJJdLdFRv0t2uIe2Lqke/KL1Q+Y+5xybf/tY362cAvm5SrfQeefOi
T4RnsvkBjsA4GAkVrm+MtA8RuH6R4qQic4TKtayAqcYVJjgMI8Z/TPTXhkTZLmVg7KY7rI70fy9A
VecSid6zFDCWubiWh2MQvGcOoqQFfvCcZEwVVkKewU1MH/BaOHXQ6tEP3CBvnhVC4gvslFfkSKHL
4NKG0BuaZ8tNoqBzSW2iB0bn/LcJVzrNRHQlV7Qr5HXhjTp89qOx4d574pKwuPoxlDa0uQJzbv25
35VHxercSrf0D9JSOCJirlvYGY6nfvrlsTHDFLkeh74YcAv82ztKLnM/u6klwiS7UUSwHUg9y7Es
87mhiMM1Ez1XfXJthdvQY+fVrxfnDHqwgszHjIJXCW8ggChvj3XCR0AwvfJUcPaYHorrj1J1vrry
7n8A89KKhfx5ymWjWwQtWur4J73OGK/JjlrQke+Uoc5h8Hj29yBvqvzQHB+FiN9uHAV0zTDXmpgd
O93TrI5GYG2LCq83cdbh5HCxlh1VgSoYT2kXFWk0Y/orImb2xjnlHI+62Vrkh9K1zFn8DKzREnbw
1oLSamM7OGDJjKbDRoui+ocgDb+NW1th7DzbITs1aKImy998D3E3ART65vuCvASKcMaoIcoOuS04
mkPux0Kl1WkzVVL77AsIB70aCW3QAAEB6FifoSS5T4dhQwklaswfDV5qI7FWsLtX9+e7LTVXYTkc
YR22NWTST1QoLdYS3HbhVGjAEMIg3PbdHvY3/Oka7mE1xjWdasDFZW0HOnVevUvghl1WyDj4UNSq
Xd429zKrQVh289BKOdAurqBjVk8lA646/+d389WPgXkrZPr6RfJyudOTh7rk+a7moNblgphlzFDV
lKnv0v+Y0HUI8mWl9K87pwBSfGCdz1Vs68fmw6MSlSjs5lt0YrWcqaAMzP+dO0ttg1hzyIlwsy6c
4i/lEoPw5AEEPtxx5rX47CzJV8hXypPD4BfZdVlw81LTb6bETR0IE4DF84ii4JGiUcr3JJQTLsfq
JkeWyGhC6zjZaJFJg+aaoM2oUIOlXG2qBn003vvgZJdTAwWi/yjQRh13TK9Ib7R1Ncrk921wXTZv
hbuWVVVO+cIt9koogUEcVVER0BeNnK7dmFCGuLdx/EXc8/nQBQ/tVkmIIcTCG621VZfeqqyHFBrQ
E/oTYu44rnjBkhCYgln6Z3ACs/BKoGTFXlB4REr1SGvwGPYRbOvheOK6e01mcYxL7mS62oS6AGNi
cciHtzZhEBqYYNIiInTloJaTXS0BCMmu5X3odOy8LlZuwG+77Hf8o61dRpgTvmvMc9396SmNWyL7
1AXufBA5+Rnr/WvXJ8iwzapgxZuUv7UNb0Y+Bakgr/13ydmvlWekr7c6W59/yXJn2r5jlgggrI0T
Lc20k26zQdxqqEhBfUomfxwbXp5Hi/ZMoQ9LbUgrnUW9IKAX7vx0CI8pYKOWh9tasDQq9JHM2Qs3
bQ5zcYIvE8m8cfYby3/qJvXDye7IKLJ9MKbmgxdf79taH9G4RoP4qDH9bWXgNLlN//DXpV9Hewxv
j1N2DZTke1vQ+qBZJe5IsBL86rhVnpwhdSCWcUjHnF2kmh5SA/t/YxKWT5GSQdRWoe2Wk9OMj7EL
oJFveJ/CovNDZ7H4LLhT8ubl/C0FrRs2AcvjJxJG62jJSSIQvJVQxCZDuNp8HBEfdTWo5Zbq1Gwt
wymb5Eb+Yrfj7TsBHQi6OD2FXhaZTWvpqvkj7/O4vF5lIPZMK/tHyPAaaXgefQK9IaBRDMkztpGb
tShj/kWDmm918le1173XF2Jzx9ytqrgFNVe/iLbotDrS3HsxTXs2AfBT2Awvi4+chyV9oN+PDO+f
BMYv0MLqipQWrJq39dMngPAAVFI7i8cR3Z5d3qzIBhWoetAELse/xE6hxA/3j4Il/l+KcjwdcgyR
ANqpdkvnDbQWReiC9F1hhpkaO6xUx1E4n6OKJ5ScTDKpyKPACgqez6QzMGibvnAE/C+EP8kpuimV
4VRx/8f0AGkD7szdl3yM5rsFFWVlj+eYgQafk7EB3ZZP+r9yEWUF76sH34LKDSpfBPYcWj9/0TZG
T71EkhnKQecAtrTOyngIEJVFM5nLHJeBUKBv2rFKe/D2gqMJ2oo8JGNEL2xz6P1ez9mgO7iwXnjn
Tky1nyC3JqBpcdnKrS+ZydCkw3vzrTsI+i++fQS4PP8VdJ2ls4RRBwtcx2BuEjd1cLlkhxBiNxPL
s+3lt9nH7YOAkGwsdQmzlrBCsZgWZrIRYk5136Zda3UbdgjdSFZJCVLoD4YUsHaFrtU+MKqjXhuO
2ZWpfOwfw1SA9BitazakTB+pgtDvB5gG1axXKzIJQXwkCei9idppISx3CMd4kNSAY8BNN+vyVH2b
sI/Q/CQQ3ngT4MjPewIxSeLPZDz8tF36e2bWSt4gJAtnXXZIJQ+qvdp5J7fyhkUnLmV7KyMPQmHT
Xpoe7JCO+Y9tSznyYCthISW1MqJseNFC/mEe3Lfa/XfqGuQKJwzmevFIDT//NtSRR4kwx9fGrVUg
LDxeBZXvsCkowVWfKp3X7SzWtyWrM+R9xSpwqxoIEP4Zv9qtHUB3Du62SivKmTY9HhxsWMsgUcgw
AmhERcug8MC+xCYo+En7s59oSdHveaBIYSvHTAvW6OALi4+u4JQtLRXw7IHwyop64llC04azeYO9
Snm6jeZznZDXyQ5ddjnfRZ0aCHMzTUY8FdtBJTYF2cpfvWpGAyPPZl6TOkj3mzVk/ApEUGVnW50h
rDr22iaCeJXdYglu9HBYXgUgreOOhZJvWrrV5tr8GSF0p9/BopzWfXuOZYgthx+A93AN5+OplCbG
i9t5fGbmt3K4BEr2dI4+hlsYqax8tzhK6tKpXfidaGkg7Py9MO1uXoprHaP2mtR4uUESV5lBnBN4
c55NRlP7krUZaYHal8IgNyx6W8F+cqQC+SSwDOkWiTEI89tbCyz8nuFoNrl2eZ+a6+2uargOHTZ3
hYSh8Uj57q8od2z65CV2ZpHXB1BlaF76G6eJvdt2EkhGvocPjV7gmT1sL3xP2jolhG/Kr16wT3ui
RuZ5n3beE1ux0YauaArkE+4qsN9JSO3VXs0KIN1Tahe/CRQ5I72J9w8NvhI7wILka3fzO+41orp5
VdrOdYqFrCBpQbfelSRyLWQZQYzi2B1TVS3LW2lvyYo5mRUaSForqNmH1U1mLZrfJVsxrN9zGFYQ
VeA9rCyfa+IrtWw+p0fsJQsg4rHl6sSs1DtMt+uFVdLu+d7FaCTiySMc1NUSaY3x/7WiBnINsv8f
EvG82f3/FyzKXlo7CyRhFHo1QlH6E8M4LLhOBZGtO0fPOoFxUKNlxGfaE1KcCg7E7kJms/YOAmpL
qqMlRaR6dmlpOszmhN6dV7vhq34WzxjOVUUiYg65h0fJeQTa25kj9UDjLt50cq6tt//ZjvQPY0aU
Z0zeLnEgkWHy3LW6PWF1eePqa/egLGy/wgI5RvLnAfFYcqwI61FvvJT1HUrPyS3lrK2lDkusGmSz
mo4Smv2+iZL/L/g6GdMrGePAX9iG9e83ML4pTJW4yqhdwDdOaMI7HeVn8gT01PBMj1ZHPBQQaLwX
MOcqdHwBtmgRpuFNmgpwEPl2RTPMu7jXsHcnmFN7TMM8QaHvlf1EmvS/bowaJoRSpJeulLKsquv8
ykPHXB+XlfkOVXoHBIjQXf1bPu1sUQ4rJWJkB39Hh6Py0MzcTQCM/ZoHjmn5U6gEfzoIXbIxwuTf
CmwzLBvN5NJGDhz5DP3FD24yK+nJ4W9RUdODNFYZmJ+D0NmedZPiCFpXeE1RV1/XjYQ6eaz7AJO0
2jNPoPy4BM9Rx8UaPgEIPVGCAq5BbWi5JeWZUzq/WZ3z08vd9hsJ1HMrsU6N4s7RVJk/zy+C2kPL
acncz8K5h9HLlea3qMRLXIXqVyIAqo7XvlBvbHeAo5TOMqa/1VeOh2rNLf8BbVXMOnl/Wg8pIdaE
zA5JpTjU7JT1njj2JwFipUphKLRMhEkgmM4BuE1vBTL1UGe1OIvgS/TDRBdHqcRotRAQMRsXNwex
PCByBidlzqfUFQvOdd5L1XV5dg5dD40lwKM+WbCguYApEQzrK2WkfMoUz0eiprh6kQT6SDxeQ69l
seNK1s222szl5nZsJ5P6cy/E1NdUqYaUkqApwYA6v45hSgpCdDA4i9/I/RhWTiPMZmAl+z3cLsGA
JVSdecuWlq+Xaqq65TNGCtsWRReTjtaBwd6UdpuNvOQpEeEu5B7yszLy8+XFhPAl3hvxgS51EdC5
zBMO2CkRJPvdD2+0NNvRC7qT94yfSVxh4CMUreleePx6R1b4Q4scTY5059C4+oVAMzO43G0qo3OD
uBB0cJMgA9SYn1/HnsQSn0ru0Z9Vp3amUNdEIISPOPhapTYpRhYd5hfHToFSlP9luI4OeoZVkdyQ
aQQL6naMb2ET/GfBSdqJdRqHFm2JNpMXablouYSRXdsf/dkUB9dvHDnqvLykwnQDpx/S36WmceU2
uiqGUocYh315FIe5uU5xx72dhm4R1eTTgZDTcc6qOwEr6y6oTS4ULJiNWYICPjIVeI/TV2iukHjW
2wFXhVBil3jxvS30y031GxkXELmtKpixibampAi/lzkHwjoJ64s96SbT9RZV4imimSqcxhzPcDlk
pq1lAPmuRRwEvzhwbFARF3aRslrilH+8KxB+EQg8mHWGQ2+FU6mNzaDLh9RwK040fF+X5yY9CbbG
Gh5EjAlZU/NwLBb2lyi4LbO0e7JY0E5qZxZhLK3h3yNxFxKMtM70oX4Ror/bCP4FVUa5NRRhfX9L
+WOELkyV5T5rSLor3WVEvnC5h+SL6x7kvRaXuzHIGe/BcTGI1fWJSOzzHRAol2Ss8/KJ6O8+wt4B
BH8d13vio0vnKX1t2+IgWhubmdMUhJi+FCe5nIXr445x+aS4h8HXyxHuJhMb44hcGZYH11Z1FhsV
R+ju7ZlL2oiTuL/8oYcqMplAT1GWVN/9mFwm1Z0U7sFq+7K+zzDkF0WrIP+Pg1iKTAs9WuCE4zdh
MokIqZAA4FiphDFu/35u5suv9WoMNwkqS8qJn9XzxJN7QMVBwRDS7JcMfY9FpiTyWjShvv1cyBPX
1KXM++vg5f4rUYaaQYwKhOWTAVMIRvHInbAKbM8YvUeqYqKtEEjLJFc+uzmN265rgQ4ABsv0ENC0
Lwlc2FsSDNPS2YUyhUw71LbFJh3Iniu5n9Nrwz3UNBpws8DDFwQ0bTWWGRRLoA9ImObVD13ezHdf
2mo4IMFig5OVTNFcAoDa24ss92N7lAJExVGo4kaxBzrSnUdZkHOXmYHc9n1Ywkc2w/HuiDVk442K
1KgX7qkQRI+RnW4qxxKgkbrQ4PdKm7urKUUNZLq9CZn8WgtQ8F95hQ15MnCwWsVu5V+FtfTWFlvi
TOmufWt6FT9fVdh1HeCA/IhN5gTVWQq5Cg2hHPSPixGK/qfGfgDmtIW0z57dx5w0zletKVHNTxSM
ty5eF/XoWZsHPjqE/Fb9kpMv7HZC/Q+9bVzndVy2Dkzcci/Y9sGh0kPC0rOailx6N+E01R3Axm41
g2JkECVVMLWSLVZgYGFH1mnQId8xyL9dvMrCFDPFcV/qDustJDblguwj9Wy9LxlC/tmeVJr/SkAQ
KCAgByVsErOyQvDQPqXck8ZF1BseeGiEOg3Td3mwxOYMZduoL6RScnfrb4S3AeJrhxbirrcHUIHo
OH1v9FjNDCApamVgmaxtbHIfGr3mt4aSCq77O8B2rEd5LWaHEkzoBONPtbJt2Jertag2NgEt7cy6
THoJuG1kPRgrrvBJkqYf9hlAxrAeC93yz1jP7FPmpVD6Kn3w9hMFOaNGiwSTcaTjl+5azHqbeS/o
XMiKn34M1NZ6bPLUN0vXpaweBS2oZPHT0Qv9T3dOmHEE01qsxq7D7p9RC1vQvmrNuviS6PVz95eo
THUMnFky8L54/YrVAwJP80bw7q7Swoz09BY2G5/339L0jb19uYAKD5uod+Xb5mNUlibToSZ6jZUF
UojtTcgLPVc/sJGv6A7nJLQKA/8/dQEN6F09HkyyKvT+AUA8iFXidtAXHmeuBrew5y9aNA82UR3F
GoggjO93iogNGUFchiYsjxB7rinem57dM31T6gA96uJN+3Cs3/r5iZ/FfXeSf6d8uWPx9duQhyj1
Dvey7J8ONQOM1fZACE61p/FnnFHcp7208VVctnz60hOLod9FEoCIaMdBBXlCXpHcsx47YweJ3p3h
X5qqcL9NPphM0T6/U1G/RLd8rZAG3KbWfwFY+VGPGPInaIUAAvFC7ixRT955U/E6Y6PuKfUrgaH8
I9YZoBRgyOgnhrQArIJt1CCgaBc3OFGE4WYYn2/FJqnWxhW1p5OvqoqTvQaxkdo2EzRYCOwZ0bim
ofr/eWgUcfW5LENfeGxmI2cmlYB8yUPGcUXojiUaP5N86iziscrIvhOs5l6MNft/GgrTgTWih/Nf
4cbX01UHXnwD9h+YdiFmucFZgvmazpT6HjCQXu3FL+dSexkygJlNHrpPzPrXKrn07kt3tPv3Sa3z
zaRCvxnFhC0whEjR9xSQZX8XuY/fkbzzwh4iWTrXDg6hzvjYhBOYCejBjrKzOvYA2M62PuMk/bVK
73WZtucMCuY2AQ5nu+avYKw2rU5DM6ycPjDsuAAr0jhmgg2TsrACPGmp2rJiRDHwemSAjQDIyjFl
0yTPEHSw0iZ9Yj8xXXEJsOq0U8Vgb4JBXVo84YN4DJUhsqPjnjMJasCCEsUdo12B12E3LUib3eF0
x0I4yNrG7ybw8rKCFDqmJzQeg6V+jN0RC5XXqE3xcXfkjLoF1enbJYA9pNRKQKbW+yFXGSDegD1Q
ytmXfyEKYJuVxkzFk662wMmziO38C99GQ7NPVZ1jl9avRKK3lCJBriNz1Doi1A7ZmnVkConWpns6
6/ZJwKQvxNUm4jlo8okkXh9FZC+O/IBIIQ3iKexxZNbCuZarzy1aUfVDQPzdj5SZ+epplW1Y10tW
ckMgkzgQC64ow03PhgTW0KDR91OaZi0MsKS+voj+gVRAKv2TAJu1guo2vPN2FWKPcgLzMImqtWQp
QqtMSHlIbTGXA2NSvFfges3VMhWg3vJK7j2BG5Er7mR9zzcZEgMmgw5qya5B1SkSx3IAeHxLU/QS
ikxAEFpnd0gKDxkLCCMlwGrp0E/OAAx/xvvf0Ip++x60gx0RCRdJqL4b9Gd1WYXq+jIVA0X/H392
6P8wPawyA9n1MF7mfhnXCODc/SVcp+GY5Ya/JVW+sZHDFB/YFkN5cTgwuxrEAHgk4zWdGhICvLCf
fwVyLHwAbsNHJZ3WO0VukM820KAhcep8vR/F8jq2P3/xSJ05oFtbxuKRoy+7zBdoWORA2tanuG9N
G7WuQnSgws5AICxoQfd9XbNdtP+hpbb+mCwgcF/NjCHazLocPD0pH9P8VE7a10wF8eBwQzmaGRrC
4iyq74C7hM9s5TyiUupsW7a/0LadtmMlpIs42zqHFhqcvBv+WG42YEZ0wwZAF7n9KclYbzZ5e0CN
t+cyzX4beoxQM8cYDa8FiDHVU3S53UX4IKTNGS2X1W+THwgqsiQuPBjq9weIeyZlY8rrsXaBPV/v
KbB3I7pC4DQTuLup0tFnr//AJi8FqKhoayMgLmbiU6O9a4Kpue3UcmtKIcL9A5gGKvjg2f4Tl5BC
w3jctwm8q2h9VySytiihWM+xTlQ+gsrjUsgVSS7kZX5U6fKmwDn3tEDikTYVpNVZJ2HN5kFJ7obD
YQGzNQhhKxchCOewnO/Cg33z93JRcRMHbpsOFrgTcBItPlahoXmt5kRTTn2xNDshhjxCefXI+rvg
1SubXsZKz/htXeoEawaYpRirv6gx1j+gIPFtrVZfqhAMUx9o6JHsjAQu8uUSjl/VOa24UQKFMqHL
nD8Bi3iNz5bSAYXraSYIjJKnMXGvj56ZzAij/ufZGS32qut+aJDemqyYGzsZPOX5/pC2pZgs43pL
BGAfBEsw4wJeSfK0nBvWhlourWNjy9/fq8oonFbFVtMLOVhh/cGlrVwWZBEPqaqqbrWtnQ24dsmU
FTZOGRKtqD2xSQyh+kRXmxP7G/rbuwsivIzmtnemCnku2Ivbu6EVjOl6iX8b3HMbPi2l2j/bmHVg
ksb+VCHsIOGNFIQoYMYfTYjqDhOcDCPxXjWBqZ5RcU1htcB5JUrT42/8/nyQKydnqUa4+hn5H2nJ
xwVo12+ChVR5jiCy30b1iLV/ANbpcagzHEMQTWKswma99xBwXp/US2cLoTR59LXX7PcFT48lWf4a
iRacI93jEQ3+2BASq55CQP+LRkUThoV6U41wSW2OeyRviLHAqNPbD4mAx9M5hbtIbuqDZx6OH2vw
3o0HY5PE3x3MDVTcVVLtRRyHK0syRFIHwQDwqj3JmmpniSrMnQl1GMMsiGwCPH7vvtJT0ll4XIbM
gQ+eJmkTht4BUvfSDNBEDvXDQgaYcpjgvyKnfKz58LZgXcxgMAiZDsafjenvs4lADqxz1fMfE732
Pucb9xwAtfHxNmwDMrSBXMPRTWjMBqEcky+uR3duYBRDlcyfNUGwuDI2ds+T8TIOPLUI99hUbEhp
sjfRxin/96I3gWqfyO3qZUeVMsph6EfBArJHfeFu8UcApmHamW9mqRH7ebTe9hzg0slRoJTtzBL6
Wk6th4EFb8XuEcM6zw4R3qgM926dVmKdzNSAl8t+F663baFCh3DvXu/fnfEskvnPFe4ekWBap3/A
BZUlV6ttSqfyBjeYlU9iogGXPiyUndc4bYukqAn8mpMzoo+oqLmClnAZm7s0TUMNJ+34Nd3tdKZo
1NWEcghrhWQI57u8QBToCcoP2s6TGEq84lqSi2SKGNtLxKX2GlGfZLIs39brQWfTsLOuxTNfrePf
cannkYmVmCX8Pajx+5qH6o4LmBNdDGDrFGwR2NGhdDAF9CsTb8L1hjG4+YWYNBqrPgoLNS0eq28h
ISPEwIP3KevbZltxM5GCPAtKBkN91pRhXXWgM6+mgC9YNmUhPlH2sLVOw55mjIczQz701PQA3P6e
WzsYyWVYjpAJfr11yL6FfJPEI5VTbFAMg3WhntxVmnjAvFknL53yPFvnRk5MHQVvdQ1IB0WfavTv
31bEyzbai7LIf4Cqxle5vDlVGfj0/LgSplmadJqbCd39TfW1L+48pUG4iJE2cVYch5KZ2WZgl+we
uvEpQbiHDWvLRzdkk082RceaRFJxaXw+7hTyGyi8uXlUC+B2Rr5OYRPkU+lpnzTl0NKjfIe2rSmG
xfAfyEX/Gp7a2HdBY8Kq4foGY6qqmPcIia2lx7Vlol4ksIvugnqvGn6WYSQr6zhrjMZ/qZF13ZHx
44Z/eD7crddGJhTIzEJNwHGdnbvVmNNmxkBjTXv+olFAOHsq9qsbO9pcF3atWVmUpFs+KGsExIU2
KRmrhGtXBwtGThLooOoZKSbo76oG/PZiNv1z8jw48ZE9ggsovFi6sKQKLKGMTupdfR0PLfw26zb6
U329oQRUERJ3/VolGvx+a/mXlcyfw4Oyw5coxKkaOg2BCFPiKJc2nACgRbRydpNNv8eMt+R9Huo9
0FQeouyPr1eNqh3NJbRbjyC7JHxxy9XavvNp4pY/V8r5FEYyLoCOdtjifo+e4Icdc3jyKluoBYe0
9031hdpJOoRXvoznrWoZew5BGR8kOTNwlzoW1e3bsF3e/hsR5g5p/qflOnl7OwlKi2wRE/HqKA75
SY+RLjoJjdqBtmscko5/e2iuKvKqkRttU0bdPQvGuKpnHjxbu466DCX3wLrz2O59/bKO/e2nAGfw
KmUbmcjSgEdRJKX5OC0Aj4/APWVbQrRxiS5X94EgcYVew3XVGeVAIDBaTLPCxmHJ3XGOZ+NCmJYY
5wLq7ZEyBjKabe7ez/nZ+xpn+UfvouP9mrZ9g3U8d0qCExiGy0nsHmwpyvDEYJ5Yp7YrvFlN5Enf
k8fVLQbfhaycojWMvxdNuxHLZVkNfz1jXqcSA8K8Vs5PUABOA5vHVG7OsAaH5zq3JjAsSZGT+yGd
AdbiKFLDtWbNJ5iiOAsY+ygadvxfns5BfcqxY6yuv1rTHcpXZrEsh1oMHXv9ziJHJwY6n7Y56Fzq
0jB7I/6v4wHGWGjZZmi/5UDqfyjimxhUOiKHL9XTGfujiRSHSdV2k1t0vCOOVEspw12st1w+6iTO
3C5yjFZCio/uH7nb/ehpdqcb2oMWaNADfGBQIUKyzVMVe8DtcgBIhxuYRYzd3lQU91nFF4oqUIGM
c5sYZXBfmGMGkbUSULJB2DGgLoFBL54valAoV9/3RbAFUR2rXHzeuuQkodK7WUklbU7plqkNwO8s
TzVwnUkCKqw0WAV4S0VsdGu7qUwbH75FR2xm1ZXH2DK1cCuZEZIM2PeTNaLyPxHvnJGWIINaRUYp
ZIKw+HNOpnCdSqnxM4B5aplgjSXa29N2WAhv1JPilK/vm0sDV5dQOHYcuGeDQnB9Tl4V99pd8xI+
J+MVF1Iq3PIa8R2nXLrU1cfj3QRHUsoXaOQzhOvmWG/rp4y6obl2946ORj/1ntbvZNVlAqRBr9gq
/qmLoRTaFiulD3XP4lSlDClMoEO82QSEdBtJGSU/YC9F7MAjxTxm9h/oncSbY6u9oxdX4QPsHtAF
C8/3IN/cjO+vilBO7ind8l+U/qEjyh8GGenpcCy+IJnmQliq9LtJn5zWrYZIoeePTSD5G+AwiSSu
ucsZAb74bMTLvbPkf0JknbNF287+kv1Zmtv2mVSVuQ4cSRDEfamr2BPYo3Gdgh/6BkxfsUF0bISd
laj69djB9AQiFWb+CYLRz7Mwv6zcigQJlv2CnfQrzmbfSatXQ3ceHfe+km2u7SLT4+GRaQEOZTgq
p7yExJCC5DVpr+YKvRZ2LuKy20bLgWomNCFvCfUYdQhTLAJjHGXwkezCzGNTRNU6xTZX8kfoAcBo
fWdVWyxBTwa4wgDDBXUF1vJWFcAvWWyhM0kZs91FefEdK8QitnZPtwG3CtNT3OuNfZQnBkaRVHUh
4QaC9TJ32aIWWmHCNptul3T8XV0WbTFI/EE5K1h1C8IS3/V5ySAn9wqqK2OZ5Sry9FrT/JLAGouv
ph6V3DzidoRC9xaVnCxgkhrg0WAKYGq40RvakNv+MkhHjNJjbzKPpTDtBlweQ/m39YCsnuS5M8mW
kZInoEvgJQ/T4Ag5Yo2KuoXJAKJ3udDDMFFWgVQWrsDibQ/zBAuue9+FwaWsvR5a++TP97oB4e+u
Y2gk07TjqOJRRd+SaIFpb8SojidfS7SzcYCz0DW6IHDWOzRNYSJjhOdCJ6M6U13kBFQW6cYtBOLx
u9GWzyncxeU+DOAxcPO56HXFZNx7pNpT/LbusFLzoBId9Kp7mDdcEjlX7GotDVF7UjBx8NqeK7s4
gMuEaF2NuShUZAyQ/TTSsUlxOFb5xwTo7TNwfQRN4+/x4AVicAl8g1zzlB6dlTG1oHZTimZpIn1Q
45W08jp8Ikl/QRdN58zV6sTjlx+RCpn3/d2ehHlNFZIyqSQWy2QgU3pJpKJDngBDkYN9ggja984P
OTfAO+2iZPztHzBnBLkw3Rvg0rIKGdwFJ5Jrc4PZ3mBH5SGulFdCOt5U8xa1IiX3G9CxRbQYod0C
Lb5lJtScpsOPjdLUD1tbjDHZHZyjhqb7T59Sf+Mk/io8qs9F+fRz9VYac9Q22APaxhT5YEuIO2ZE
+D4pXxMjxl74M/3Jh03pxTkBBdoBqlWR/REs94zU4qh5DetpLj57xrCethKJbBfQdLpQ2zMkXeyO
+orJSpxiVJOM88pfIMUFgdJxdXjt4p0PCkM2A5BOVczKiyCc0Hnc4TIKOPg+jHGXDwxBVlmSgQHc
Cl6cFvNKyk4YtMm91j/eAQpVU3xUaz1M7SujANnti2jMrjfsNhm10aQpdJoAuWObK/IyREWVIBcg
zL89KEo18LkQx1JVweN8WUacuiYBwBkEwvaq+NDHcMyaMfOhSuMlrnq5KluMmfxrU+wQcmvpuZKo
wgm2QAJfeeUm/9jPjO1lnurdiOuhtvCmGWooXb6k1+cvWqWQ2QwqKXXOHPQ0dReh40coCx23kCPT
RszsIhEgU8lHtqxPDcEkOFd/Q7QcA41T1yBXULV+cHH2Rvo9B3nPci35uJNVcl3mvyPH0ZuSsu26
l8pyYGPsDDGVphBHWuMRktcChvmz8EqUgZmOVO66D78P2VU4cIUMj/+L9J0zaBTFMYV2Mq1i/zMX
aYE6bBysqHQKQdTAQOK/huD8xbJwG57CXM84xionH22AbFfiOrdytCvDU2UxLV0U5rRLPK68D9uU
mxDOOtX53CETS/bTLbnp4/0RQsiJ88nMHey1mJhS2cZ8iFdL0ejgpgygPbF1OV7rbWp+GII9oz56
MbDg455mlE5hnWa8tG3h+b/DFVn2Rx7RYj3msmkDD/TAGh1UGPc7iJ+eg+Cw+jRdzrLAt539PVDX
nOSbrysM2qlJC7t/itfoppXfovykJiFxxO8IRqE/vhsGxnz+Y3Lg/m88bRj8s20bFIenqBd6ob+s
N51ieZS2ocYQtOWqsJG0FA3BQaQ0WRuhQwg5DZ8E218QnQJNhUoBY5y3mWLPAPgDgdSecoG4gg3N
hUqlTFH0ktAvG9wtYHDhbnnT823Jpf404ttlsjsPFgkHq3WOa8mJ61rHX8DCPo3Ek+LZ/Bq4rKM5
rhvQBNwvxTNgLIP1yMh+0GnbyeOxMnhYG41B8IOcqPHktMHU2QjajmrqScHCGmtnU5ASpNc6Wk99
QBGFdMKI+8OPWIFP1JnI57mVJ2UlQjl9tEiPCnyFP8djI5djlO5fR4SMbcCnJvsWMXKa/UghUHCE
aoULub7E/yORubTaxBODu0sHGaf3DehZvKmcas8eFi3vdf3euvd+rt66dpegEoRpjGIvGlc03vv1
vvkiTKvVvcVvfjcIv1XJmcKPz50XhpYAVpy6OI7xsPp1FoiN9tHeMemlGIEviL1TLC+XeWyyx5wm
Bah/3YqzSAJ7vAQsoPBpeSBRg8J6WkWBjX9RTsGwwb5RkY6rzi16XQ2cjHwmACGVhtZ9wXy1plcB
yN/fYvdJini9WEF7grZ+TK4pDWoUgvQnl8F7ibEg39GhaPU52vJ8lkvOuQnwgOXf+fZwXvCkecoT
ORlBUQyhWB3TurqNQ73nvreJW6WoNdWLldDdGFuncKFd3u2FVjf7PS4ZCx1BVKr30P3/ExuIs2VL
v507MWoznACNLAmQg0QaBUVcZFk2KpSagVUleDH3yfZzVUBLiNdSBzOXip1p6LBMelw8rYPKFU7Q
vULL/cZemyU08dfP6iPB
`protect end_protected

