

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H5lQJsJvaeLLGFRhK1oe708p9zTtXNXItx2KAtknEaAF2yq8IXwKFiVPbPTO8aJ4G1wQZMrKgMvb
6zlyKbmneg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RUvUfs9jruf9OSb6utxk79ymugfgdQ2mgDnw22tbcF4+w9YY12PtlphQ3EwSjE1BR+YNcfcg2ppx
nVp8oQrlHaYHLiZdJQiFcET810isTDBwI9+sjn4Ry8+ftUrGRDkzGQghSG1UFCnSyA55dNVCduAa
//ZGtYPCXRggO0BwEzM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GRoj0md2TTeeyD4XkfgAjr1JI8z1r2plHgATS4H88EONpa3oaJwG10L5TE6c5MDXVxHb/m1WeMVh
VBt3w5S8h9pf8c485G3a+NVnNsA2vHPB4cEC1yhvDIpNkeqj7HvAUARW4zUkp2MDiimsNN00ZMVQ
inLzBlDW8A6T3Y2b3GmoYzUXaMQElMyS/PaVNF6Se8+PIRjTB8Dv5G+A8K7PF3j0h0gW5LdMZrCx
isigyN5NiqJ/3ZZGLkd5XiuLlr0DetrgHdwfifFeF2dmLtMjIx4kUkMG45tToYmkQS3jwm191cux
eXIUgmzmvPZHik85i0iZegdiOZ1LzY1yO5OyEQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UnEKB1f1t5V+eYV1nijBv/smbMsJH58WebxNSKYwmtj2m6R5AlGEZE0haiR3VYCxPRjmiopDDdr6
uBQOF41DIKvZSm6YCypTeVt9WvkLpXTJIiHnLWz3IV+uvKXohhIry2Pg30NMC2EWPfi43aTNvtNH
ROJrUVVcDZeGvVPmgRI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U8EV7GGC48XxGZ3G4wShg05dze1bZdqSUw7dITFWVJl+2U1VEqYTGCRl5zpa3cGdqM2+nFugC+BK
YIux1TwcaF2Ng1I+Bp1k4H3BhUPfmkZlNiGri0KnFOiDYzBROYyyiUUX4IECNCLZnG/OtNfakQoI
AjU6WqtEEQ5JSpZpL5mpGWt7jGfdl9gqPeY88IdcWnasDywKSPqo47azQ0KIzwP9UejnEHChmHgr
3Gpvmrmywo7/+/EQRujU1oGF+ysfAmqchOGtHLtDFJ1h2OjLVkv+puXArlpXpB9wZah1XCGw2FON
8d2jAO5M9wEJ2bQpFyxmedBeZ1Qj0cJQKZW3Gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51344)
`protect data_block
XhMeE+Tv8dsTX5NS2RvpxniqL264RRDiElowtz9gUu8rxGz5ZOeMsRJJFrIkZmOrgLmI37gUpmEy
1APsX+PZLM/HghSHtQVuP+ZLaLTgjoME7LOD7BT12xUxfUrSFYlXIHKm1HkcAOKvLnQkACFjJ0WW
PRg/oS00lp1ZtwPtsCN6LoJw/2eAYQKKRep+jNeuC7Dk5hVxEZLG1XXalIQ3DttPmOhHA9RfpAL7
KIBxR26EgNqaDLHH68CtZXbdiXWsdrTOTJTmEgHT8PhidkzOTvFc4FkNGlwqCYTFfpZoYkQGEITe
3KuEkllGrlQ23SLneCzq3Sqc698g5vhaf1H9y5Pcol+0nfrUsEC4snJaXn8LW5MPizXFLcBKiFoI
u+2H3n0ryixJx/eBF5juvlhjf4fv5Bfzr4Vkia3CKBAPj8696GeoV6Wl4gTj0QNxaLlrchW9lZhA
5BthHH3aLMksRLJnLnh/9iMFgKSOU8T7YFdn09Wb8WRt24BBuNLCeCyBqftFOCE7C/MLM0UvJrlB
4MlGiiL+z4ABjBiGuEIN5xPllAN3H3eW3PCPl3rJHGKKpkmlG8dNl/L78UQx5nYdpr7zdVKgF7NM
PQNEfqh1HERFmXglNPx+T+gRsbQyHJjSsN4R7D+CFBvAoBcLMIsbNEAqK+6JdCmAvGQ94l3YJO46
kSmXn4AiJKDvcWHCu2qlmCQQFHsv9azOw04LGCHtoDZyB6hNXXW0iCaz7WgHLCN35N0VJWEPyaXS
AGGWhRS7mjoNWedAHtPQpTSW2I3MLyByJHf1KGTTb9EU7+CG3g/6a+sQ7ZqRqqiHlwt2vIAonU7a
VzTkDkzR9hMa8fOqQgV9/NozFCZyhtUHTO8axia5MyQYSDGFUFxhStfejrOLqYa4Lhigv8yPR5AM
6bFFnMIl5odRc15XeYFFEmtDUFUBcStRt6s/BYbBL8nNVTioSA/H2LzmEAuDKaiIVakom3E5iPFw
EQdgValc5XvwgDA+A5hvsDfO5hSHJKf7Gn8fN7LGu7xz+NHAj0ipK6dDVYLUrBdptdcJEXcrXL4i
yvALEteSYniqTdNM+RSoSgllUxsRAmUnPakj0Ce2UyCZNdnJ7R2xVjUeFdQ9oYkce/AfEK1nBEdF
hnT9nxVN1Kho3eEbpBkit0gF+NCzTVYYxixwT7yAK5rNGkllWaSr/0w7MMVwyFQ7Ria9v0RPoMUs
EhXlVGGzLgersUYXMHvs/9AXZbhhSwEQ+xAuMrNPzaeGWl3nrgSGr2n8oqI0GI2LLVtl8hk3SyNk
UzIwfJriq089bqfDEjVNRb+0T13FdibnYJhRouE9iHsWpBLYreMYEPS0TWyuEhQqDhOh7AD2J3Sz
KO/Q0P47ZRM3ICKyzVJ6WNvna+TcNcqxoFUHzY9MAE6JE+iMXL94zmM6lCMRRkI2K33f1LiVBj6P
bZSAnotAWQ0a/feMv80dguYW/FmW2BYYn/zVA/s3FuGp1QMTFejJq8tonoQSx7+/B/JkjYArrtpM
bMeYMiOo3AUUwQNVpnyRA3bgL2Av32r3wmaFRr3rlfn12qEpi5ZuKYwfU08MdQTjkEaaaUX0t+lk
GDFnf9SW46g3Z7SeY1oDIpri0vjd6NYCppXg+ph2NHmi5MhVhQGuQ8NVd5XxpMC5HqjI85AxFqza
g1RlelO4AgoblzXRK44l9qg3s/Z9sTDIUU5kzvE+h6ucVd2DpQ86gsPheoiNxDU0Vg2tl8VyTT+r
MYsRD9EhisZPtGxk3Rw1h2ji7MemdP9mn5PXitOgKzYP8KBSdQcceww0KoDR/1Cf83a00lZUjPv7
DoGtOfcFHpKrBuTX7uMEAxBjG8OTIKh6ZQaAlHG3TfuKDeGvo8JYnInanOF+Q+YPZIJDd5lGnq20
eWBule9TWinic6Kvi7Eki9pIRDVLG8SCKxYsmRCylMSiHwvYal103ihSkLRCXkvpAKBdvhWr/k7w
2x8i/6swBJtj9n+V+UND3v3s7fppweghB5S0BSO8Yg3UB79pVuJqAGOFaZVMS4/Sfv7YpyQRhIGy
om7pDvhlu0z8XLalK64Mg6xbV0QkhknpIoEF6ErSbevkWvQH6/TJ00tSQwQaom946TbtPm8/1N9K
paWeGG0utDjRxMUs+sVGqYThcA0YCcdB+MuDm4Z5zcKlt2kxuV7pC+IiFjE2NIieDG5ceD/ljFph
v3nDJBpAU78mL+HGc5kTT4Iz8qRr7f62GSdy/jjMxiajTewBBzpxFEo6m0xIOWDDmqe6VchdnkRr
ITzwavXMQVkbIEbicVHycraItg+1vGlxwAnSyytxkxnq51aZDfRyiBQC0QS8lojKWBfhwNDfgYh9
ZjXld01u+zix469jB0DxenxXDe77W/ZqMME6PQHT5Wl30bkgx+yeRCo8w22ZBPWV8ZBBzE3MELsy
IzK35rxI5W77TE2yAp7ZkI+MQP3qA+PggPH6DZr9cTNmdgi6Wxij47GYIn9YU0H2PSscsmDVcTeK
QoW9CZoeO5X13SgBrCy9yMSXxZtelWTrLbAGJH8/DcGiU+Q3wfb12AbaQ6MBgCoKzn9V9tm0m7+K
fYNYsX3MDdsZMyl+rntMrbaLxTvH5mvC1M2pMlesjUhLmpfdXJpXjbaQG4Z3s+MP5me4aoeHAsqv
SPCPNMEqUiwxd7vMyP8sfP+hQiBdEjsUam6GDHCrBCADcmwQ2nQ2wMLKtN1DPwGLV6PXyM8QRA1L
mlG/a/OuIHEyJc7kbKrFayGwdRL+Zw48WAY1HAqgPZ8Nxx/HQs3nABJtzcnihv7bJppOnYgt9U8K
YSNcLpkUVRFhtCKCoW8IVOtj+GVK8kMHU9n7feodR2igtmjSavI4P+kXxgFwG8ZSw8dDFbzH6zQ2
zsrMfmm7oKQ5b2b2jfTnyaOSV4h9OvwrjyOIStT5SE0DOgqI4ldii5vKsPG0bFGDmKaCR2EHqTFm
hCtRGdrghyjVczd4TonLcXzGXy03Hf7ttCXpsgOl0VuMVOgwS5vz7sccLBzSCdOl3jjRXwQmP5VK
HyLfh8QmXVRR+fTXpg6eLI72WpdBUZVHgMR9owWA9A9HYbmXMnNZq2Y2Mb0efPcGb0LkO6CL+sOJ
d0VzZqntOopHWkcyYJOrSAGVry1mF4RArrExvZGncH4WK1wMOcXbcMY8rCxir1hkobtBxNF27xKx
OYjml3kxduNLC/ZBeWIFZcn1bBP3BayFn2aXKIH19TCbQXzfDwkI1A04f+unwE81l1dEB1DtyceL
8vQ6C+GHYqnlGYTxW8dCNVwhp7rf749a9NH8g4psFY4bO+dqyNUmOYpb+OXE/qen5Eq80+vnsftv
6tFOmxxTudqjDYbPpaGEbyfa8mDjb6NI3p2440lPz42eob+gB1zBWh8b5bHP9R2N0rNOJ3iHFvlH
HX+6Cw8h24Vfr+6XGV9yyi2VUce/dSvKtgTPxC052znqqrFxo9j8QCLnf8qRL5BvadulWXLpzEM0
5EHEF0R1giMuafW7Yv2+9lCVMHNV5m100xpVnuEd9qGJyxCXU0hqoNDaV9BosZ9c0Xk4YH3OMdWo
Pysd3tIjErJmLdYpS693O/NrKfEp2BMCruIoy58tAdvCi/l5ouNZa1oYGhAXIw989waQAOJb+ryv
B+gfQgTrmpjBul0MwTeGu34vDAptn40Ftbg5yvy/Rtl8h8D8Yy7NbFnn1OpmwMWx6CaGyaZknJe9
PERpsyKL61gucZ+qLGTRht787pgWtFXlQt6nNgr6NjS8hNHkz8voDWb4rF4pVQYdxy7rsBU0Zch0
E/MuTYrZnhJVIGDhYtOCmuiZNQWFi3ZsoZ4rFsfT9xl+hxy0RxkNBUtgfKz/Y9rJ1OzqdwnxQC57
CQImcBuHNTtszZphSyA0Xg+PwIPq25DBhKX2I+TqLR5jbSqP+wdEpU3TomYT4woGonJ3ro2IhHIZ
DQbdVmoWixpecTGUdS1kmhoM0J5kloTrhOZLj44rRNjZMrnPghSsmGEvA6c2ZDrtPYKNyz4afpjv
s5k2pAQ4yORjWmrLs2v2w2bmRKlUI4oA5CT/jTsLD16c6+/XnxBHAp3gp7+hAAYl5gDSCZ5RzOPX
uoWrQeTCRdQPc8GDoXjnyjZstB4juX8ePt32KOUBInNYol1fXs4SqYuxs4g7LCQ7uq3oKyH597gw
9AsNGoHUrs1ZCqLjtUmtoPznDCJjkzNQGHCyGyPb3J8xeEJ9/pXDwIegu7bfABc9TUGFIurwG6S+
8tS5HySfHNHHKLJNcw3Pal1AO/BYvj7M7NY1BUEKqtIst5VbJWAs1alebbG0p/VYtHolCjazUZOC
6tdVZJzNvuDO1+bdQbjHM6AWzbRdK7lwd5wNEh4ZnxYiPa660/2H8Xw9tKyAGfGexVEnOrinpYej
KIdVSgzEWcsNWOWPsuQoBJ4IBDrMhrmES4bGiXWEOLpc7RX7GbjTIk23Z0G3mpZqBunuLLFOqoSi
GSSRgB6DvxLYedFnULKGAP2LrVSQqNUmEEfjVC83nRK6mqVbrEiEGL/YEPcrg5wQBdaucEvELvX2
MD8jBQ+Vji61po51TTmQXww9fde+OJgTQQbGldLVttlgs5BXgbi/s8eUwh0s92BUqQz6RHkcJA+c
tjIxCyFQyJFSgrtTb9/2yC9w0On2tLmkbqOPeAENd3i+AqQh3n/Oqo/LrZBF4CSFrqDDIarqfBFY
9Ex3QzPQhtz82HUIchlQu5QVQBmoDvVqLGfnS1ilxnycEzn1xbSrxsjlmWwKZ+I/3n923yuBOTDQ
KeJkOdRpfueCJ+Ka/qHUuY22k1XHq0vNR3+DD9hsjfE2qzpGgrs5a+a+hvSq2JNgsha31xaCmHLF
XRcp8LKdsPso4FomORXjRXqsOXbiQa21pxGgSo5EUQWB9mJptynQ4GL7yJJBhAVqEWyBrLe/6KNh
fJdU8R4uP2Les4OCRYG+/G0HTIriMX+5t/qylnQSoj/jxAyq/6yONi0jjW/ajsVngm2cCU+ioHiU
K9ty8T//srGYJUEbz95UZwFk7htyubWHBNnVNynsR/2GVMNmRBZzbDAQ4loWJqroJs6E4pAqj7i5
2wxP7ZRmpuNam9y7MgUBRs+TPbG/g2VFkPsCWO1Wee+4lO1ENgKJgBLCHqQEXJsIwjoaybETagOP
ANpLa+pdLV0aeVkyQVCp3K4SGDbwG+aU/7m7u8YM7exVZEd4YtAzYsKGUXDD4z5k23KHZPkyFiDz
ebUg1IopnJ2aE+lUfXnheuSUW3zV7Pu6XsDdbaYw+x8F8hilROwCdKXy2M//tentpXl9YzqEqZj3
1MXX3swlORUmxan2euQPF0WTrGpv93/Uyj4qImPdDrM/EmSyBPyPLiaxx0I5NIbold1EMbkzMKo6
Zr/rl3Gu0brZUNlXOiMD5ti1KuOZWaNsATxQGPH9vb/6o5D2dbzHd2mWUquFqg3AR7xi2yyAPiMZ
mW+5Q2bRj0W+fYm6zlrxCpWpXjc9wr24t0Ug+BE9fXc+o6posPadnShxLDpMzSihBYVh6J4Biyqe
YH2F438HcYBqrPXPueMs3ZylzEkfj7SCyTBf8zQyJY4wMBI9HM377gmPaS8lqftwHjOe0oJybUKZ
fu4iOMqYPMM/kbkPkbQdqG7hHCE+PXlzpfyJymo0ETbMwGQUDO/8aQS00jw/bzzo6icDRtMhA1KR
hIBrI/mrLL+vkHvBcHQeJllwOdJwnhiuc4YSPbe9YzoVfJ1zmyogOtzcfyRtropoSX8xv4fE2vHu
tOP4SCoKp+Ooyw8bSccRRtq7OAR8xPCxLqrbp4/9oA79rPChQr9740WoTr8g+S88+hPvXRAvTMvw
xmery8qzPUaXt4EimSO/gb0SnPjACBC2p9t92fyc4hteZnthT6z1m9v5aW9vzIVhhrugh0IiJWrX
vuMAWtS0a5CSDEr7/OZABcb/+VVw4NzRHtFiAPr1mJBRXqekwA1Up+9ocS5RD4pdOGXK9M2u4LZ2
o+hGDhR1czQ8jcscnkFnfnvRnvKg5TGKzeJsSNuVqbztVYWIHMnMCFCn2bJ4wXxlW8bUcqHL96id
N7H3/713qi5wIeTuQoiErB2BoB+I5HWYph50EoSeUhwBe8rx+QHi5Fy0zDh8I7tEyrwxHuHVTRQ+
YIFMpU6tRUh+XipvYjgTTqOWHcBXW/tDaBd2eUDexV2FcwjeL7FZqJ+AG/gYQmMh6TckUe31T9XU
nQ7cCNRNBZKRleopWMBjlu9QOqAvOMMo3tAjlFCF6Q0IwOTwBPOWTkV2VyNw9JqA7OqgNJSj3MwF
CRpK6oqeVn63d6ZTr2kqgkbXPO/rlgukpgUkLDIreXORDiyjtYVEo1CjDxfkrbxOA+kAHMoCS4BX
QfWvKUxhpAexQVSUFzDQ+tgBB56KrqWQyB7Py4GmmHuP+OYlGnwPLAMyf6ie74HmQDdBUOILBgcX
OGt0xfK7/UgQdzieu6z31+5QBk73I/GiPg334MbYkYwyeBopaiYBxghFlR1vLNX4N33LbGQzWF2j
VBj/6Ye8WLSRqHwj/vXMAjp0JEOL0accsK3353Ig/YFbNCTp7iFNYlA9oj8eyWnOytAeycpID4tH
z3HHjrLNCrHzavBqbU5oLt1xJ4eVpFDjjvnCajsqLvjlQWND4dUfeLG/K+mUYEr8GpU/fxCHqRty
M3AL5eERHP+QxQFbtdHcmgpvXHn7oYctGkn/RkWGjZbS3RJU7RuEkY5OitMwI2gc6gXk4FreUgMN
cVo9hIXap+j8M0VTdQUP6w4n1TUMUKdn58na2jCn2G2eSOcG5DJfS6pO7bypZuchErk8ZNPfhG/4
rdbhTYvP0sMSJTBD+mvNzBWtwia95PfKnnqBHm3m+Mn7TumNcWvtMhWx0VLzbqTelvmaxbnys3hb
i7WYDWtWMJ1WAzl6Vq0P/egD7KOWVpjyokxYZDbR+0OXWxJVavTcIAL3Yr+DgAyIUDuYiOUDR6Tf
JxraOCwlXb5hnzgHZXIlHfm/LLbYbnVWjr1xFNfCxnwmYBCnuqIrEOwrrT43aHcsCvQrJnKz3gi/
vumGPOib9bTB1jkwSUbsDxFLn8lUA89pwKKjocnzWqJGcgItYqa2pAlDXnvYgMkIAkGgxLnzVqRg
0EF+vIkd3ev1k3UdVey4X3eYkTVzBAZ6/cTsXNCIcsi7xYxm4QhciitlsqmaSTHYlagTC4cx0pro
/obgoYsWz24QA01VSnzqm529gMH0pdd4/EB0CdwTmaVxFH3j9GbnF1aBSeJHOIU7wvkpppQRaA22
u2S2EW0uzYW/TCQSuCxHOrfOrYWlAWtlG72YHeCnrCX9CVzW6MMBw5VbGJTgQWwCgOMufDJHm5ip
+q1+XIRt+WMczm6f6sNqhcmLimxFCCp+rQBlqR/dcf5A9ASueHPnMjS05kl/qHFnBVD6UI4F9Xqy
IunkoOuM2TP7rcbE4oQ2HCsupiUFmzN1y4XBbDry52fIdOLTeBwKcQ2tON9U+7DXaQnC4EMBYYvc
Vqsc0vIP7oAApjsz7RXHd2bt58UEl6VF7dvlmnLaT1UVQfxx8eNnWyn5FzyCrPikYQmnV7gYJd3F
4pwnEV9o9p2ZkuOrCM+N/zpXdNd5mmGqOmyBLQUo/yVDSMoWi/73vo4ftgXuWcyBwdMAGgYwrDs9
Em1dAT8WrhPb9SCrFPjpuC+UVOU+Wz+RB2vZNmmliOu4o+SvbxSPTOvfzx+I4u1vAm1xPgOhzaCh
SPdp1LB0HN0Hp3/kJFzfyAwnYl0n564YFIIbprdQVSf9iny1Hmd9wq143Jxc3uidRxNrc4fa9lK6
76CIp+Erv3Iuzypjco9VPP1GAk/cKjWkqYDSwRIGeUcWV9p9bPARraiq4WLNZGMS/AkRXEHaDSrq
wmwjCLaGgJxfq8Wgj46MjLEHqW/mhKq5/s36KSPL8YLXoD6BL6raC19Iw+5GU9XQ35kMBaDdQI7Z
W3DMYMBY95hA1adBkt21rSUpMWVfwoT4OGCXj33Qoo0nHyF8kR5iiiivTWlkKxaJLo9xRLEKc3t9
cfjX2kU/b7ESXi645m9lj+SNPsqSM7x1j4uzB6azYM/dN4WttdwD+14zJl/XIVZzEdkvfprAGzZw
8/X/TyJhT4mGkiP/4walZfqZsUfcFb3tckjJbtcyJWt14/K6jDkqK0O13zHUYAT/XIpQuHqLXgdM
hknHgMfYIPsUbPx9ahZBY/cl/1EDjUWIKQwi1h6pBfkV3ktq07jlsM1glFZHOIGDgAlFq8nhZAHu
fyc5rpFppHJKMKsYpFZKgDBApNZ0yyyKn4mjSt35HUa6GfRucN+/5R6GcprcWdtQdS+o+3Cb+dnp
JWrTn16RiPGYT8O+1p+oOFBFMY6hSxikfYhbSZliePuPO92sAHD2N8K77z1AGJLWb7b0+XI7xxQe
mRjK22GqKzH/msSjEuMaGe8smZ2gb0KEPihf9nDV45Hy3m9zHICbAdDD4Cp60/BeLo3866bACfDb
14qDG9xtw80M8Qy66zNr0WNjdsCKwYbvoyAK1IMzDDJUnIPi1j6vac7YuoJL90EBYTFxAwkwk6DL
VXSvUwe2NIP5XAAQxJ3ccZYuBKIJOQphGV8twNb5IPE0vXW44hdb/qYiwqn7xjt8AxpabqIL1JLS
nZ/Mm669xwhN2car7IJgsTbcY7Um3bRbGk3zIdtVPpV+9h0T6hmX96hvSonFfd/n7BGOjJM/nKxj
QqyktJy13PaZG3qLGmCIwXUInlhiciEJrdX9cNwT0Tmkf5/J+mtRqsNSiygqh7mdAFGcSqWAOWQ6
3WhrpH0f75ap1Kl9iuegOgWdORRO2xQrDtTIFRgmjTKCpfkJBPsKDK3WIluklS424jBZ0F6awXma
W9M+tiKdiHVGrFS6fJydxzPOnYym/X11kh6l8kTeTnII1r3wyItTPKSfO+T5FlbJ/XHmLffxGnPo
BD5gwGy9OOCWpRoLipTb8KB9RsUXlkrBq1uiuqcOnimhn2CZhKlDTebotVSsL7p3GsQ6ghT0tRDC
SMWMnnCMF/+w4nAtMG9U35bmLmXkVx+hLIGnV6V1Sjxeu9mlR5XgWdTMPzwnbFsM2s7j5LHMzNHJ
y2WWzpyI6m7gifi82HG1X9ryYrn/P/ScUZidIie3rvyoYWSPD1Zi31DdWOYYKAHH50lMMp/D/X4r
Nd3ivTe2Dnw04Dc26y+f2wOyJTCnXfo7qZGA3Ix6BD7H9vQiWKZwE3Xg5KACvwF6KTlLEjRfosUF
+jNvoYsbBBh6CTWn+t+DqYDr7iXaQSeEi68+lHqP2IGZ/3GiF7elizcJAMvOcII82OlzXRqHKjt9
VPLXXMCPC8Nzz4Utk7+XG43S4sFv73nDypEI+U9ITHZRf7r3Efht9JGqH51pzuoqeX72pTizm0yj
HqjRHkMUJlGVXDCDmqJbexpctZsEFuTgOvu8UVdltEEnKiBo+FDruwKMBXigx8/HOZ6drq0Y2TBi
LTctN6PbaoCtyrV3MqXfaj/mcsYIVKyLZiLzYUbfytOPhE0CZ0V1UfoFNrvKYc9oiA/weDQswZws
rxqk7bNvXjazbph1nSWFopcYk9Jg5KOUysew2fONDf3yGwD/yI3KhrK29qtnEYh7TJRTCG8rGIus
i/ltsA0uI4Qa2bP++1nvP4cHt0bWlC/y1+69bCtweoAHLK6SsvEnWjp5oyZhBlHMdUbPcqoocg29
Z7uz+0rPmPkmINbGnWQxR2Do2xnjUcGik/T3EG1uvaqC0OXgk5aEPjSS5a+20XebDOPUGW+5qCiU
ZE7SLLtF6iayX7LFWXMW+5aDthh9mIViFbBba7qqJqObhoCQb5fzHRiEtpwMZZ6VrCqFUqJOysUT
L7762I9LW9a7V33EnjP1r1hda8VJFAeZbhKFhlCjr1GPA+wl7Emko0HPIH2GQNq3e6c4k7fO+4d3
RTpe5t+6YDAQdJgCraVIRHoL4sHd4gYQxHa0YMFZlYiZBh9sfxdHPjxUWOwdIgfQqmu1sNceLfsv
vMU3FMdcbagP8xCEuDrU8W/Y3XOiv5O7xM3LqGabZeZiufoNReKQOpHlaHfgt2uwvLPD3f2sa1Zs
jbjAoTGMcaTsl2/veLaAZbiCrGEJOeLP5Hn1lbDfLiG3FwrtZoLFoLc/KgONggPpAOw4qvNDLpNE
SVKsQ+H5o/dAnyWuOmzpuwunQD+ZvIb61B76BOSJq06wdHltkrqtyTXaGETlgFVMdWKtxc87f8IO
ccYP6KFvXBZsmmShVqn3w56FDs0N3lAbhr+qZA/gY0WmstFlQtVPiN75smaP6FDeSf1QABAqMBW9
l8vUBGCkiPnlHhxgR9APw0AzZSQ/MDz3JSO5rVyrJOg7I1yE/nV3mI7R4ma2td1fw7eDHBmz9FFg
htbV2F6u1hcHiYmX7eep9L368RZ9MJxub7NpRIKXyYzRmI2j8jwRk+qAZ01Ynf41R/Rn8+JtZURF
UDDhPyxaP6euh3vmqDyp9zQAqCKAtUgjMPSXu//p59VZ1joBKHss0Dat3wcUaXa7ibaiJVf+Mvht
88w7apewQABuEnd63uU+9EbjazrEAXejwJtoUB9ct6rRSpExpxajs9PpuB6ScF560inI0bOFvajV
7qr4akvq7MX2gas1dfYTOLERynbVUEzc96TvYFRlGH8V2UVAgOactrlpr1yUGEQc3llC1IwRvnT4
AB/dwiYXMtHIY+k6KVPwjWWsZaEAPedg2BQztPrREE2+2YQEsy5AX6yODhJSzbuMXIalUIYCNcs7
qs3qWw6hBZnvHnDuw+QpaDJzhkROaMTje5ji7bLQiHN8EjH4in+98UyiblXIoEUnxwhEhInOSQUe
RFiicKtTdttxmWZbCN2r++0+a5iRNts3PkYoCGpSNE9Pa/kLVaTevJ8TC3uHiWzG84vHbLddPctW
SvUWArz6GtMWXmCb1mkY9JK09Q4zHyAiYdCOqwNMBkuoT2RZnfHwHyJzegokW+TcHunTY5WOicTe
K7/M2B279Z9kuuf44MHA4oMn1PsAg8s4HC0V+vB6W3drINAuJi/xnNId6WYhfzI8rkIgwKKvOxIr
gnMDYKO83oqs2/RYWE/KNJiRlGOLZPtHiHczQ+nXGnKDPxWiOylRraklcXZK2+cZ4UZ8A9QgIZzw
qGMAS4A1Cz1Lrqr4GcdSJKGhlFoxHTV5uI8p/bdjaYdWJ2QIfI/f/Rw1C5kFncLaBfDuN52iav6R
HJKgQdlhadPfiaqJLwotxwyT2LY4zrv5oz54i10KK9dQ1eav8njn6XQt99/9aAkoCiwpv+C9H2fT
0Xn6WLpcYJx/fjzvFVvvThF2nqfVqUgA2FoRo8nqUaPXS19RSCKuHOKNrExpAWSNA0BkZR/19nfj
ahhyP+MAuRlJXG6NRcO9ciBZJjpbc3Y+ebNMxsfXRqqHI7eiQ/cN6sxZyinUFE3GCvXMehm9gMVC
kXonPrPyZ4aJd5o7HNCIwnlFnJOIL+60SzvRAf2nVUgdXe3moCBK4Ofa6HBrCb5e51q+Xn462GeM
XUTHdF/SU8S4KkKu3d7s7zeTYmzzYYA2NTyKVjngBmNGBxszT8PyZiXty3Gi+OvlMYOwDwryVgu3
DRfD5ARDuWX7y8oNHjnohyQCLO1jm8dick1e+HLdVXzy3uf1YHNw6nNhDw6C6ovGSDimKFIW3ZWU
p32HmaFpuMPtdgeqDOm9XSYPslUvLLzsV1ZuQY8aDKOnUaeAF0wRLgCjyU+Ys7oozXtKMVQaazas
lXLNkgyW1dqrR2c67M+A6ZjIH7fblOpnBLvBdV9Psi7wcRY/ne3NqgXnUpr+/usX/YY2GbTLrL1L
ECiPXGR1DubT1a3r/PZlRWPiLLgjdwzOKKKdnJ1rohpQ5xhFTZgfLMrolwMSWuxQipYpAy/dQSRN
iGZg7cn3E6y0wzr4QIjJRA+Qkjzez+I/Dg4Pam37DPVErvON1gEKlNpAts/WVdrpJ7/u4dyI7e30
ICWZltWsEyCzHGmtu48tar0vKehvOM7ggIZw6PbVZ8iD/Yzmh+v97CXEc0nOWSzdTNNjJuK3yf0F
ZZAbqkzVsBjpxAs7aPSCPU+EHuOkEpuIT/8PlVbcrru/3WLLYnPPLwy4zyej+WJ7kXX2k06xeH8F
V9LkgSNTWPfc6eSScdazv9gyLwOUT8RQmoKkkxOHDwozH19YjSgLdU6zNpx1oqxIXdeQnUYPZFQa
EYCwqws9ETeXr+B+vYZhcwZJ++YrP7ThyP2+V44iA2fvigEVgMquGEYrt36UQLexTPxFf+FxRQIF
WxcfiYsff9n/3U8BrTVL2SBzkQsOTO7kHx1EzTcoKojNuZgaZQB+WOEtzvFCrOia7S9iv++e1EFF
fxdF3UK1Iz+P7moJoA2ZC+08osmNFZ8AwS4fKm7kVeYmx2ipj4dF5YFK8Qf3Qzx43qyj+PX4mdwI
ssRziPLpBLpOdb5brF8cgqacgdjpXZ9HG3iC1K0QzEqUN6Ba7CbY1g5gOHbE8WD1RM/3yf3IP1Qf
zPc1qxDSZ4tZPSAwJvoqaGX1uneLVaf60W+lmcL0MBoGAiZZDWJ+8GN0Dtfg977DHiGj5CR78Teg
iW2KI8eB5Ip+exjZki9u+O6CQvEbPIXkR1S7a0H8AUfZAwvxvPBKPioAOnVUvTx9LLs0nZ8ScAGR
o2vIbXxip8muRu+l3q+4l+/mhHZFcWq7qasD+tTY1lZNE6X59X/GwsKjcHT/rQDMJpaQ/rEvgZla
44NGiI+lagaRhXDWetEMXFq7mh0W/cSO4LhS4ZFxBwDueGlID0AecM/YySASfwA+OTe1NnMVvtvP
55qQPFsFNAqMsOjRXa0zEkqcOpnhmXh/bwqCVuxAW1DLfW/vHO0bhks4d/baT4kjfl+68Cwdt77V
lJu2823C98jGnjvaclcVkUsgQb8PelJAQ3guiT9jSM5rh8IU7cQE2f0PoVcAd55i88vzb1Uaucpp
X/KgKuDAo48MCtKgKopISB3BgVFDVGksYZiz8fP1/Kts2LHxzxdDFpnppk4Up+3VrnwoHRwAzLSC
LG+xvGPBTTsUEKvMwsv8L4zFYNueewFGCuHrZp5kWuw0lN5XBDfLRUqn9ZsxOgT+daBA3UDJlL9S
aNu3wtdN519Qez1bWzsdyqcY4frcsrCEANlUk2zWOdBI4VMAu0GXF/KBVOB9ZBxqPpXWGCGWmyvl
a7PWqyeflEnevyEUZXmadgfRwjmAIzRPFKrI96T/LBl/JVi8ESmJ7PksJ7IJHAgg2WvpWYpJLZYT
xJrqHFDLNzw/kBFnMtdOJf91qVb7QnVlFTTif3q2l9rKgTTZGtaa+PWwBNw7UW8a4M9J+urm/sHE
tkt4C7qE2ZvHbdIKBRN3Y0mwdbiIzkIqs+1xJ8UE8B1E+3q8MunpSeEObP2Docm+PA7VzBCqEQ1e
2ywkRgzY2PPHulHYhiHdnhijJsk4KofN/lygVu+aQw0tlc5K/o3zvri7YatXYGM1IZjd7LT4l+J8
OPUWupXcpuVhGj3a5gNvKXhXvfL+bZGCpBqPk4uVcUcPHnZCvzJaPekeRVc6jpX3KIR0GAto5Zg5
OGiLOpe8dlRwQdBKIFciLvaUsqiS5aUoFrkNnthsXikEJJZXg573CstIcdKSSQuQP+gsRBDuKGR0
/9zqgNkFVcnfRorQ5aTZVpvbsIFDMZL32tZ9O0E+imy7WzbnCQUPPb9zNOdLIzb/wOrpUiux0mif
2pYBWAE8rXsvxa6JhgaI6xzn53fX2Us3FH4tr91RwN8yyzTcsWqmoZcIdev38FdUfnkMbVsFzLKp
/X4Y+9Spabdu/Y+5AGw6x44/xVGPIvCKQMCKABo9N+cTH+0YV2gx89IaVxKW6aNShrABnrBl16oQ
Y9WNHeUGqlY9sdqbq9Ii9r3m/iakTe3NmitT5D9HJ6w4G5OTjzqrpwh6nBC7WEWXoC4J5frG9fq+
TLgrec0TxIPyEw3fISYVtrvl0m8hpS+MzOdcy6PymgQXtciv89jysoRXCriSsnU85Iyr4mnWtiDs
CmJ3LWGTXRlir+Fcpl1wJznVvF0EWkyEsXqpnh1vkN/drbiA7d62CWmB5a/i75ggUa8NBAaDNM54
LgCvv5CwLxY3DRIkLMlRSAg2Aeij5c3JtBhG3fj1XB7qv22zlZ0VZrdRQ5Uas6Q79FWYQW+u7vpl
uQAMGOQdcmYb5P3cqPXIg0b1zXKWyeirkb6kXhWuT9sqYzp8NBxMT8yUrR7wWmhmLq9JsAtJOZwO
F6cM46mvXCqYW5cOTXil3nfDA8Qc+1n8t/zri85LQamJKviQl5sHEOsyuoBKgWd3Hy6BBWYwZIYo
asdxr4eDDQbvxUwpkKKYfrMTbaKlMjCY8Ex7veKpw7lx21rFZSpUyhBzohqPZRO82k/ktjadNit2
lxhs9hrBvWiF6hvZoKcLa5mIbJ9xlVBzwkX6kXTVlykVy6dU87KaD6GS0o5+iXmgWcP2MF2i6tlV
3HvLv/c0lB+IxQOd1+TB5gb+QmiQIIQeoBMlSPLE3gVFNhsWTvZufsqwpp56LBZ6YRYbOqUwyXbe
OiNXlfLTMfpyZUz1mHgrr242HTpfVWegniXvGia2GJH1JbP2m74xc3jwIx26adGgocVLiphCzI/K
qJ9BZBhvk0CC4XHN9jNmBImoCtNNORBZ9WrgdELqBo790s+gF/4OQg6S3Kr+WJYbwmjayA27Jizk
OkfU2YG4K/3RTKL9Njp0zDUDnf4147j884f8Ty7SWgqcQilFvvwEuU4lkv9kaVwd+e1xpcDayr2M
soExpQAX55CTFixtoA2MdM6MvR2bKoLe1WgY9ZhI7ERkm597J5rnrfH1Qx6c8vhjOltFJuiBBem9
uZzOnWvV7Qg2+OzgO68VmIA/WPROS+ZnOYGjg+Tf7tFFYcM1jhMeNkPYwjExVCqFzqrfY0Yc/rnG
TzmC7fWWim37q50F2g1+C5sH3wtZcTBx/LMe0+y5EwFuoYou6krK6JI8eqBJrfXMx/E1C3DMdXXG
fMgdTRtd0KyYE3SJBOMAUpqpTxlGkADKjxBlJmikPsxxFR+wKoqiEs+WJeaKtFzlg5lp6wfCpKug
KKBTJUbUm/ZhEipVRFM1TSfeVQU26NSbd4aA4urwijR67oEJ4XOhij3MLHbRWerRasw6gMq7J75q
LFeBztlyhqzpsBOhivufDvovM+KNg38S4wdMfIrCbe0Ng50Wsao4PLZGSsk6BR3B5Bn4i5JY2FEm
HIx4xTy9ZnnYZxpn0/UNyjflqn6ZD05H/K0hqP9S1vINA5DuHdMO9jBabPPuSjvAowZ6AOy/XZ1H
cCHUDIM36Fo3Ghor4kf1NmGmeQXhSPrX3RBLSoA+EXaqtzznJZUzfqWdb+NLi+dJIy+3NY8t9h/s
AiT6ADwJARq2CMuhitECIJoqtVEfCWy+pbb+gO+L4y4zJ0MT4md93e7Ye1QLL7M4bQW/gaZhwt2c
cSpY5y8quiR60TgiAlozfH9x2hLWO89HQLsuTDLYUYjgyuPyT8bfqKuDnf+xgajeBZMNtPZY4O6e
9rn7Cx9w5xFd9hCErhYe4GWgT0TCCTWJ6u5KNCGeAzNxrfDDnyjTjE47DVyQIos2j67K+EkpjLIu
b99MsTs2yCjSfs0QqCtdjN6fU3eC4su5zGvCCIeL8nM270B80HklKzLu3ePTXqNJtZEDLKyto67m
ctTG1oE3hHtvhnnv9S4IW3NPOEXrNGPAkNeJooWCnOEl5VmldOiPUGTLWF7H7KeFtaHvs2X87Gmg
r0bhA/t1mOCl18CbEEyw//U2SANV+URZonUEjneo6XxaDFevNcAS7TL88lP1sZGLPsX0hhT7iqYB
554FFH5pMjVe7fySGBB8Rhm53uKf7tjMskHSM462d7gml8X4Jovc0htIytq3J50vo5T+iW72uA9v
NEcwpOJAPhqOz4uqT7ezv/vqYaG0vpjvueH349Gz9gHy4lOK8VQ1R2MwS+pVOt5JmbnFh5s3NWSQ
5QlDnZOEW1thZEe+4LIdwAIMmbM3ThvJXeb/dALuWqyPb4dwz3x4ObFjonlz0jQyVU8waf3UGSfa
oKCiotZC3aO8prnBCO3y1ljhlZFWdxtb4r1U3p+JoZKTIwU28NEBEq4XJECK0ByowVW0IKI0uBdF
vcj+NQ/qnb6J5RB9WpHmWek5QekcqT219MeAsITUNkwCcwXKEo/myNTaw1lEjkE4FdIIf/slVjEC
+WwOInPobhpR5Gw+G976passbmcafywlpG//RLD3eg1quvelyCIaOIevv2y/pAUZFJWp4EBhQjY+
aZPRNLvbNKmW7TjE1Px/8SsgHgaAZvzi5Nb7TVrpq4Xc8Hdu6lxK1CnPHc+A7wTQqGLkaZOCyIYU
2SEv8j7vwhIa9VZcL5u7go/Xs3Wgln2FZUAAdDj/ohEBMS1lDY+T1U9Uoq2A13fW728/oV8ii7JW
MX0URs87ybugkmtgCnzGFmhQt1eEzaiov+E6TcxSAqI2scuXvNscsh9Qa8DfFqqjo3FHfVwd/h2W
/fJDBqxqXpndKHbr/QjXqiEaoT0VQL+hToNnNBmvv5pnd6CXsCedwQU0iaw6WpbUfqRQU37xvaB4
Fw8fXCnS8Ma2IgPeVkr8WnN7UNdopi0lhkGgZK7fQxb+uqQmjfAIcXiE0OdQESusm4+nEvMZOmXv
lMXgHTzhL907ShhPuRo2ZJKXwpqsvoRI1MfAx4dWhzER5MDjI93yWJ98wJc0/SzWS7nwKEJ++bxW
OMg9jTQ4sw6qgDC/LRSegfW3olN5SO/vo16CeovsXOzdJO2hQ2hk4QDuKYxXWi0rgjSqjKgH4pjS
JAxpgbBMSGoAsWnlbyYOzabOPmZRVswRSkw/dYSaTnNSaXdossy+8DRnFM76MZJCB296rHQ8OinO
ZYHPWFf/mg+WnOqfa7gS48BYlcnxoEWUx5b3rm23CLuQQQhchZC6xjo47LOF4nlb+jGJServwViJ
LoqSvSIvNPNq4HtgCaVEuMv84Toph+KLxgXHr3jeggHuB+mFjG9fEV19/SYubG331irEn1oG22GR
0eU9Z6Lq+Q2TR8y82p6Q66XvVhJ4El2tPHDzgNJP+wUifPeyNvrm8Ocv5hPl1wgcS0+szFnlk8tX
SVkC2kVYiqr4Q/tGc86eKO8IC0BfFMeS2I3vUDRRHUvBYDmsLmw3n38hCFAFgkOQ2pZoDrWAm14l
/IuuqdazdRKr9ZBP6PTTAaDTscfyylE3EEV1Bdys9+FSj6D+yECcTZZbn8mnN7tGTA6i5DR2a/PS
fCAPbZsY5r/KazIw0FxQe6WEtqBFwEFLt3jNVul1RaKkniT6+yCzFT1UfxkzOJ2ZM7wCz+yl8rO+
XUfXlllXG17RP22WPyF5byhWI5iQE0nMesxA8LTCPXRE3AR54ysgSQM6rzeJtREDAIcgOj3NdmPz
tfawg9Hr3KOKFrEHe4j/LQXIlFjKCZSC7A35ziWB20uOkJsfFrsIHExV179X0y91l3zHDtpO1I6R
yOmgD68mK45HNRFuMZl6VJ84mHIXnWJDGERiIZITSm2Qc0xlR2UOgqoIKtzTy3k3bwFqIrSjEevD
O+1Zh/vWYzjmyj+TCDqmy3TpOGRuZxbQjGLmmg7Rjb6zjq7HX0suHoYL0rl7tCFdeH00V1c1WC9g
IjfIs+/ZrZqjo/nx6Ct9/zfxFNgo7dbBnu2GLVE9+rWD5c5s0/3OMMT/uIhR+ooYYzunvhcWtggB
rCAQ6KYfioSn5BjHuiZe5Z4cktQ/IuBWnPdtklLwAo/W90ZSLgYdnksZxcRcahgk5sdvyfGsyR3M
YyagidJ2lS6pHkJKRb9DtYhoq4VTSOAmCnrsu2PrKvPrrqUpGGqyKMYQICDvUXdxV6Qr5BfsL764
pyCfUoZI/XnkQhoGM/YG9LYLO9AV3PQfBF80iBdpWEvZ0n2UFZARnPS5wxonTQvv7f24ucQ6bsZw
hVg4UoV1Zc0pZTbNC3WjJ0gMg1UHaO/PTqym1boN+Em7eFsz/SSJf1Ryf8xSNf3ekUEbAKqu8A8G
rvFVQFnkjq9CtAJqGF/JyQuh8/OdD/Pu8+5/ZdPAh32mezNOgvf07Yx5N/AaS98g+GofbtiYQV0p
TDTPeEClrvJvYCE/AILzHsatSvkLsb0c0JB8Xkb8bvX//LB5DhU825pGADLOX7AfdHvy1P1ONpnQ
vfb6ObPM32ZOtuM2xvhAA+0raCfT5zPmqQ8NZK8YXfCYG4iJtttDlrud+4thzS62cF5Z2ovSeyL+
42ATNtfb685N3AYNUHOmbOSxOTEd7DJz8sTBS+M9FoWxdQJFS8ogo0K9YWjndB9GtXhbJ2K6fxQ4
WuCfmeUh/o6LKUWKJ9U3RCPqOdvoMS2b/aFqsg7JSTCMFX/FawgJo1BxNDjtRVlXdAfF2zvMg9u9
/iauKIOTzYH4e1BcNIUB47sYXqR5Wo4Gh6z4KN4IrpBlp0eTY7eFmvA5dMeQ2hpIShF4WxqDF6lQ
oIJ+78FE34EdUDW+3yaTP+4huKADht07gGN9+XdE8l+vdVVYhQVhUo8amk+ULxlT5eBsWyJgjN97
5NY8a8dmJYvOJGWPUVHGMDjr8QvQQf2b2aFRu++6byAOrEIRKcNdwlgBTjVQhG3DMv2E7DwJUy5M
PUVNwpqfgmXJnkJEBrSxG9Z4J6Hs/iqDslFpiQiZnpzKPVMmebPDlSH1QX70GgdxbFPAkRc3fv63
Z9h2c/+appr4q2RnMLFb2lPlfwKktvhAQ2nlCovDPDdPDr3E/STjCe8TEAN8a4LaMEj7iDvEPSos
eoF/a3IzObOlvtFDV/5Sk5i3VEYJUDOyrzOZCjBerVf3zCHPxDxhgz4vt96/3j62qIdyzU6mKVNW
85W+cb96ItLucDakL5mVcVbtNrv8im4eua8O9hn3TVdbOiJDBEPp2zz5MeBEGcp4oBnzkJOR0YYE
h2RbyiLgx7jTsNAH5SnqK1wis0MJ7x4e9YoKwFv0N8fw9zyjUAoMHxUEadem2urfX+5WtJSF7htb
PwbAWeBAiFBE82JCfjWx7Qm9whv2XVXUTgyRM5RpcF1R+1TmRdVuxUvFwdC3GrOjVG2OwJ4KgBge
Q4AgSv0kEuEMu43iIxpk4shBn2C79b+GyXoBKry7qn4/Kv3yTCwS3VQHYfGrZW9vdes6hPVUZdyO
06TvDgr+zMcRruzPUAmLAsNfEHYs7Jw2Y7WAMXk46hilfBNK3YU5Pbj12Lbp6QJsJ+ALya+bokV0
JmRgZfArS/P5Y97/+0QMoAvPBwjNeP92K9u8iIXg2BqETGtICplKjw1N3GIU+ba+3dIT38Z7/wKa
6TUEDi2IUUai8XB7TUdDLkZmWRhMZnFjJpXcQ9EPrDZYBx+w4szgWky52dwyhLmRl+JZkvV2QwWA
tsfUzF1CQHlhUK6Opq5AdvHYvuzamG/j1BlbuD5SRVPkoSeho8lVK2DlRf8NF19MD3O2VGLpWOs4
PSp2pL0/bxnOl+8SC+ProAK6qQle1nyOCk/E3i70vVkvWX7R79s7d2YGxWUndsGgiUrb6MkUxevJ
M9r/MH67tPlwciqaQ6IMgZr1renHbtzcxC7Gmy0mGSI7eU6uulvjoNM3LkDjKEdr8NXXTenWoXAc
h0YKgv8OSHk1vageb6Fa2KIndvL2ewWkVQADw8y7eddYOD+CgHP/DrA7p/xmq/T7bdCrYH/DEeWX
8pzFbypDfLFeQ7CGlzNX4KI+Wm2Z2kvLCHIY5nHSLt0PJkJ/DKef0beoY300E43Wpx3fUdELyx5R
erkEvwdVqCBWqsff1o30QjEbcRE4tNL53J3A9fCCwmartb2jxtdAHQV1NKQVtg9ij518scL7/fii
Kk36kPA0NAlnl119LMkDj6ivsi81hhcNQC/oWYe+aBd1e4tKITHSEHVrCJROYQiN+VLmNrRzB+b9
CI0fx/q7IhLQA0PEwlM4FOO8mGwPtw36IKmIlDmmGUjp2WBtun0kC0pLRZ0iRmMrR+Senlihmb89
hfQuWT6j5BGPdGDoPdjZEVUcHNlt7U/OHVJNubxK5PSK1yFK4DMXnCSXjQaiuE/8q20yRkRYzlta
rIyf9/dy/WnpW+ovtv0wESXErXMKg+dp2lFqMS5MrQvX1/A6HQb+XL2mxQO8QHLzmxMN19Wwy4SO
K1sLmZTfTBp6pDtwpKpS0P4VnbVshRJv4gGJCuZ7deInb8zWBallpO8GywvJjJ6k8ffxrqwGA3ia
QNPrDAQko/zG8l7XP9n71tIcSSopU1uOZfwt3ivV9r4xAznxx48+R6AtjAYSSCCmZWNJ4SU1LNTk
D2owsMj86RzkNBSuVWo06JAXF2yppt2mTQ0FjwO83aWZXn9cdmYP9PzYbdBcvaHIKeZMwRlbfS5o
Z7qtvTdvj1fyww5ABdVjIyw202T2bs46hCDpv834afWmy1PPbtP7rLesdpewIziuh/wEzkgcew/s
55rK9e1Eszv+i3Wq4hjzylHFiwDNVJMt3IER9sVkMQJsqgMCkHKSUtjlUC/tdJnbKH2ArVTsmZ05
dGvpjO4k7wVNPcFfbqooJKA6v67kOiML0PZYI4URBb6T4NF9F0fKcn9Et0WUcMdGSQtMsSkRgmUn
z8JprqBLqMMJwN0GuIGXiWaEjKmcT+d+Ti60KtVG/VHUxine1Rgap/+uVxnqSFoNKATGsaRPKmXD
vNuFnfulJBPvUeNge+2u1iHv7XEuqr+KE7nr3bQX/PNfDjH8ONe2UpqT0mFcCF+q+jQUhy1rHGT+
Ap3EJJN6uvd8DJdXtVzmBOvI+UgYKD631mSH0sM4Q0/3+PpFRDQhos2WFVjt8bkiMX7fBWiZzd5m
8mIk+6U722j4UACKGPCBE7yuOs9+0P3H51iuCe+e8mTSr5aQ2W3jZp1FRtlyfJGsYGpTjeCxElR6
xN1lTUW2KGiIimPIoXrhzmW0lWpEfZfvbQdO0nioWzOIPr6RdMcfbaup4Oc3trIb83HftnZ4thZC
8X0VLdqBVFoZxXZ+8hPeb/Z/6qWlXo2WmpINKicjC5nWc0mI+kkadfhC5vFrEG64FOO6bKczedxX
mRaaRAhgmB3PpJxca4+Pgi9AI48XfkIQGIxt96OxbiHXk767ajvX0Kae/fyy8E1dOybiCNICfzW/
OFFju43Ucsh/FJPuKFw7//ZjbZ+mP9qMtBn7YIiSjvgPs6VH2r/Df6zhYKbFBchhow35iVf/8zq4
XrnNpgmSdaxF/x4+pl61U20dkJtZxNeeLVT4h26nsjsh2seojp8DgRsO2oiIYfW6+UMknDXgMy6W
/uar8pl9/m62cXN6/j6lUViQUPnehC3vMLa0icuGXbOTu7EtExXI6ZObE2USaQwA3c1Ha+zRwD1E
BxbFq4K6UTMUeTknNRwAj/dMcMP55ACTSnHrUc2edtGXe2o2ugyX16J254dMCYZ1J9DvCg3OzoQG
SpoViSde5qk4W6lrosVRpBXtWezkHTQPt9sslraGosqiU4dhd3fmBlBpxcPEMlnEAuiKN1aJUHDm
7l9NBbWB919NMa5NwLRTIsyHqgVzZN6IGRWOyQjE0Bfe8r60fVhsLew8ncqfnMyMGKxEvUehi2Ve
MKQQ4XMiP0LHBLSz+1WFnLRMgk04k0TKpO8QcOG4J8LLhchSHnGwgrsD6GlwAMhUbs49bNq46z2J
WzHvCyO6IvsTEjEuYfLvPOBi5LRaSG47X9yPgNwNZYKYXLt439quqWK9zV/HUvVq1LaFx6rqyx2K
fF6YlRgNYumXxqENkdNfhZAdtMV+N06UMGli+ryWpTVZ5R1NLDbLIOmVf+HaYZlR3WiFKeIhKfsw
mLaV3sAm3nLEuAQhK4EV84RpLsyD7SSJVdgOVbedMs30SyZJt7tmDraCEYDmETBk0vF6WVaO3OnA
RE+H+dLc0Q9YFFT54D9q+ISbHn6oFS9DfdT1rCj/bTj0zDQKBbLDi8i+xbRfk4V5wmdPJZ74Fg3r
KJMkesX2nvR7JPLUnaDcPIV1VuBochWPivvHoblIIdIUUFLjTcaV7ypD86UY1yPvndSzN2b7qjKG
qfVYkxbSzSdDh5Z13FlFSklrdHwXiTm8o2wwkuNnOdHJUOMl1AXUFPN2ZVYd8FeYaR2ZstMsGCfL
M1IJ9/oB13b/PdZzpvYcy1xjr0F7vaO+a/YUrKOjMQmjd0bfDAIVUYjAbombw4QWTwgy/xQx4EYM
H74/b77S70lVmt2ET0WbT+OvID8CmM5WcUGPvfBo1xuN1CZ4cSuSID6NZxXje/d+f4JeUeLOVHwl
9Qpbq8+k27Zb4my5qgfzWYI65KK65dEHb0+mUYMzj16Tz/bCWGSqm6K5AwdOMILiazVc2nD4G5x7
5IUG0CCCNGxl5Rbidb7BlhyA2w7EiJCdJ1lyoMl/myWoYHX6+szMCIW7VPqPa3hUqJEIQxZDUsLs
nftnjCrCxGKSxRJImc1ZagULy9Xkvp941nstrcCTL4gUx5znNvsjuXuZ/mnx6mQSzwE/f1DL9Y1i
swN6eb8OPnvRFqaY5qjN4Y3bG/pa+ooTgRdno4nzg9vGFqgeD/6FO6opO66Y27HBRwTs0LF4Rk+2
7m0Gosh8hcdn/+BTa/kZVkro6P+3AoKtd6KPCGYDdpG6veI4WmIS/6TA+uDydPvmKq4Xg7n+NVf5
my8jNw5rqHQVmlux5aWhZk71B/RyySKGDtMh7YfIXAsgqgl+LEaYyWgzbPY/A0SbWK835J5pTRAt
g/E9XJ3sIOa1dCADa+s9SjcxunuE/i5wrspW++eJWMFP+bY7wOhJi+wBzPXOGv1MkBKs7HLr8XzT
3+Wqj1Q9aLKJpW7MbTPFK3hqPfeg7eQepni5yB7x8ZozRyYxCPz3nmG0VSjDX+rEdXxnRy9a6+1B
/72PlgaV0dvuCD/WQceybM/IReexPMeuyKT2f++9migJi8M/lFyvPJEj3ncIRrBxmU7ylcRgpq1Z
sLKw2KRjmlvTkl1PB5q39ylhNWAeSPwH1+8GsH3fg3jONitTmCbyxSTny6VUYVw9319Rx9XiXgl5
SKxNf3g//cWPZTqMmwmrq6kxIGuAPc9XiFdFq3L6BBKs5jTyjTeeg3m+UJCVfjrt725xfc57nBx6
JwkzaaRaTyPDB3ns4XL7iT5oCyxwmmMzpgG3g3UnFrafJ8Bvr+d/eX3DFt9MB4dMAZX4WLK83A6V
Ce8DG1rE2N02CUu9DN3RnT6g9G3ZZOcqCVR+9AYnUBDAKyy48y4rgGuBfIv+zNK5x174Sk5ptiJZ
oFlZJaIbslxK6aM3t/WXv1Bo970hy+eCtrkNX2oJVTWHUgpOaX4ylP7WBYecx0lzWeV0SomJlGug
VL4pcWMgpE/UleWT9drhkRH9ZmahNex0OuSKkN7UG/x/HWun7/V/7EONhL34BPhmnYq1gekkN82x
Ggc8A4JeZ7uPThSzDOzH5OI1+3bIUK3uC7IBNsKPYGZg/nwkCnQPA15sQSfQoZNba5+X5pmXZF27
cWZr2oU4z5HIoZtRCuYjz5FMTvqxBagGs2jxjTN5E7hFjlRKNRP9/oOxDgGMHZOVkG1TG5dP+OlM
nNDrHhQ+ySxpkpX8U0fUi5BCKqcf71BQV84Dy6DUzSq5R02172Vl79ffUtrHyJGGlBzQx883VQr5
t+PZBUSeA9YQR44xv1ReIZz1DeALgklkqd/gwnr8ulwNEORp06WAavicYxmU2ONtEpBVSD1NHXlT
nOjYKLfebqUOXBFr2HTzrZMBnWxE+oh/IyJs9HFp6ETmQNN/Pb5wioovzI6TRowt/YmxUW6rRkfE
cTHU4O3ZtNVodoQAo6QP2czczLIT4Z1e/wTZ6VyPWBct8Ym0cSPlBghmjHyx/INP5v18MCljBLbg
H3DIgOrMKc58/Mhds/mpyk5QMJAjEVT2ZrQIeagLYMvV/YwLw/27WvLq8NF8hxh5s1IZnMZvPNVy
xmjtmbsIOB5cwM84ByugpIz+xQt9B84WB9F01zqtADSP8gJFAsUpFxrDL0YYP+BctDSLEzcWXeo9
zH5TJtjA87RmGfqTFcWlGKegtizcpeNOfkLC3yya5zDXU5XfaVcyTQmDgnFMhHacw4uyL69oFH08
ut5mlJT5MBHsf8an8Xrx9BTzyLgjesD707xNcjYB+UwPCjfmnO7IgIXUNJ2yfZEhkr7E+d0SYIz7
H66rGNetklzOPfAaNJXvK/AXOrndgSLRbpCp5tW9L7CvP2nvw1Dsvgv7E9QREjyOk6qz5M1/hmJ0
X2yb0l0U/LgDIwaqZQooandDcL5FZhMJteCylh83alTQOpHb7DL8CAIcFviFSzFPdlHFjbfw4Kl4
EBKS/nyrK6em9+STBWTkShF9bpQDL6uHsXKhEiGM6rUb/058cU+bwDa60mPBiNLG5oQ8rv8V4Qm0
fFY+hyn3VEU6xbrTeTrkrFiaxfSIP+GLHJdH9APuqUd9DxmoXMA6n0U6gGoaaKKJ5XnSqZciwqHX
hVY8flHvSX96AzPSRn+rW/e/zGQCaRYj6DxkuMm60Jx4dBLqdulgcmSJAd1/WvboVLrkgzP4H9jF
WpPXlomSOH9r6SXQ57yIWBwBdZTViv7h9tA8iZTzEHIUSluA0IPoyASGe2PUzzXVesL8bnFd4BSi
mK16K0Rff9Mp9iNA+HUBtxqiRaM2kdVYna9FMCgs61YWCMeqq3C6lELfzWifk2KffGwF4tB21KCR
6p4T4AuBAm+pRob4D0a9Alw3afOmjtIf5HDFTPZHv8S422m2fU74dup9H3C5E9awDm6WFqwid0as
E1kjCbXJhl0sPArMpuopcV+xrtrcadd88H2DD1GPeE9l1VmFRlu+K2XNMAMSDjKTpP1al6bHwRLL
QlnAI8uOF02sZpvjpuFkiG/py47DEoLo6KtSNcjeAZTY+Zt1FxhBhrZCjBXcrtRuVN6tNcqolRl0
f8Fsb7FIjSTKWV14+ljOmlzaFUqbfP0WVCGiSj9BHNxurn1o3n8/hcunuD5Vz8izbXKj4h7QKy8/
N4rfM8tvp1hF24dP8503x8iO1Q4YdAWSlz3QTgqxJVk+5xreK/gjycLTJUAm1JWlW9FoqMPZXMl6
GZff6PPmNt3K3VXzbxNB3wlEbkPBZb552TWy7uTdKmGqsPmrmwpNsaD5XiDS8WHPFzNsGkAGRjio
aUx845xEasEIXHebnrTZ9r/GHq5zIO9PIk8whzODL7zF4Frscu6bNkAyMOCNh9NsKygeiCRnUkNc
AcCj/Ttzccb+2CPz8oZtfmL+4CA9E8X6qPBEUR2ZrTp9SB8YBPO4mpzADPCd96bIGLM09yeN1FEP
1euRgqWcISpF3TOiviTD+Uf8+QPzoDRb62uyRwAKfh28Mg1MYuZoqC7oSNnOKQHxJ/WaPLI3upxw
wuheg/NiW8jexxVwushJXWukXC53y4/EI87ePW/c+/aomMAWYZEAe072uXMl4v5CBFLjKP13OhVH
l5Mr3PNHAwutx6gItZQ0USY+7WkUSvmQuC99WGJByn9tu9ALE0WAFq5ShNNEMEIfa3AFoZyy4Rfi
XxAmt3oMxEwYTL1e78D6fOZFKC360x82c23z+7bpMJtH6vXPO8n9n5QuU+nZGi0reGUBajtY/Tzo
XnQk6AHD4lKu/5Wuc9kSLDMLIa5eoZp80YZD55a2+nH+uThznEOwskgoLbGnpD+CaF58yEiGd6dT
bJSoKZoYZ8fmawESfysYcUQp6TL+3KpCg0PJ08MZ0ohVABmCdkBgD1IY5nRkkvF6haKamQVfhhEW
spOrmyfwnFCmLooyYsi+Q7f5J1w+ykto+YJeRmxP9l2RmpRNeshEtaY9587pnLcyYLnTBf9sUW1g
lPizOYRGr9hlfoQlXrI6r1qLEw5T03qX+MLi7q3yy9GWuTK2GSLf0PX+mjhhpM8yaPnavESN3qpU
ejVMZvw9qBRqrAIChde1LwARDBc8liYf+6shSX3z5g9+eyROlKSiFNlkiLLZt8SE+IMXP5i9SxtL
7BlvRSOn83VIzv74SbIM5ascXktpaHKMTqT2L0n6wObyx06Plq3Sk3wIFHjCH+BHGjUo71RRAnWL
rqonTb4LrywA51A86P7O++4wd3BHaxCUdIeCmqrDd7G+gaJm7QfnAuZk0sJrDNYmFIxyX817N7T+
+/7iYFgDiJipChx5XcBYSmPiYmFL74hi4JTboCqq+LV8neOAC4YYntPGn7w+B4tMNSqxiesyuUcN
YT+IxNyZd0sw+GEO1uycYSALzIigRZQ7wsVlKgx6/SXzQYzwFiD+uMKopLvcPxpl7y/9+dDJ/NBM
bPZidQVnrq99UmaCtNA4hxOFiGxKWwCo0vaGtJmUqQo0RHOLZOoYwt6COuSfSrB4TJo9jUfmslCI
IvI7pbuo8/Kxx43+mDVI7t7vdXgkajnV7gf6WnoIKXEY3kyOeDmoDLu3vhvI3YFSH+kqk6IXEjyg
k85BL6X366pbpEcZBcqSrs9QhaipnW/8qvJLFBi89F9wV28jNpDN32jotUG8OOxjOxsYMUPw6yKL
sC8656sVomJJAY2zt4cRUQ0PNQLJUn4JQK2YfiQB3cdhHWQt+7Y+o+37jXiAeBrl7WktAL1QaS35
NtudengGRyxCbb1rgNhrkYaxHx25wZzOyfA5/IPdjZeLZ55NGSth7caVDkNse6HCTxpHD1x0ZAUz
5sP48SRgMYMtDxq7/ePDVUwuxjNygnDce1j1VKmbQtX8YXWEsl0R5kqv8T6mGKyjxFNA/44ZD0Qy
W0oyDeTE4S+axzHC/ZkFn5Y+SgwFaWYyHg64KoI+mnJ4Z/oHjRk2H2UIs2OuBBoL/SwK6tZGnUJc
4b4Cqo4nsFqANkGJe1KSLTzOcNZEO1sNwPkO4in9d7+oL63Iny6t5wKD3TAufJHuToJFHHXETPzy
THCE0EIIz6K/3m2SdB9VWQUL9snYi1xuOJNtkuS103a+y0xi55pClneGV3/VOqhXE1BQC/JMkIVN
KXnRkjg+felSzJTR33Xx6gtTjmNG8DdFYj7ornNX+S0+Nr+n593nxmxwBfYyn6ebJq3F2zzGJG4z
4t03jO2hbSMFq8TX+oiYqth9ZQtGblPvfrsnp/yx5sqshRdPyCb9OyHzX5dO61XCICIKfCYF4hGX
XKszmg5UYnWb9GXF78LUklJcCn2ZOiAPYb/kNCApuF7C0xGvyju17m83YAPlWmhcG9ABtVfHQYeI
ulG5nwq3bb83qNEn5gvpOYEGxiVdzHT1HFdXZZVdfjTLRwzvlSThFBmSUxYXRGLA2jfuyPYMOtGI
GVDa0QOikKPS8zea7Pouj99l3ahIJ2Dmq1m30R93XyBifn3iAotQ9vBxCUPSyOjc5gILwQRX1Nh+
rgcVfrgz75xOmLzOhr95OQGshXlilDpinyJIP4LmKKgU8pdiZuRFCp8P/M4jeWAzKlXsIPC/tVME
boLwptdw2+wYEXsmGJnukOPiJBNFUMyvEapSTHx8GGp5ljbd6P+rn5aG0AMewhkNjRRcRQGwb0Kc
c74TgHh91LCwxNxcoKK79inlmicJbvAoBZXkgyOdpSbb7jXLaZjhdYpb/E/aeuMzMh9aUJox7S9f
lxAnVOAlhZv7O3OGl3KLqf1Rut57QjPT+lqrVutBsTHc2mniGiFNq0unsR8u3NbeJfaqCfZbzvaP
CFUvAE5tgXx2QKd0s+IcGGylK4p8PUzKgvt1iBxOP7owOKOMWGGm6GgsqTco/L0A5uCL4L9ADl1D
/HRIrYdc/bdQefNoBsPEyuTYFW7ChGJs36gz7V9rYQNwqxMMq1e0Hap/gTZ6JPvFX7s4RtCJSOYi
GzO994BVq/h+qVf6ofOKvtgE+4Tb3ojKnWQUNEIz1bADyJyRagpGZIbbjYMNBfIA3H/OWIVNh/hs
JX0woeY7saW+7ltvy7o1YKvXrV7Z2s18PWxWmCvuL63B6NytKBb9LRAEvL0+VHGotL2IUYFV37+o
j7gU/j4RKiOboXPiGmCUwOmAq19OdR29MeZDiF4UcdUgm234EOCWYfX4ecHthVmL21cLaDSrGdfD
ogKUEtR8679zW57n9VsoZfJAgeLqstb2dpZKDw9Oa2PBXC3l0Wkrr9Kg49XUiwZ1IcMvrAKstSDW
CCIHbtZWwsLkfdQYwVhfQchpa/IDikQVnMtxlrLSghyAzMwIOo4pWA1HXfjHFku6Kx0L9NO2EC6T
SiZdDKo8JCHC3F0DpBw9Dr79dEMQTtr7SL9CKzUdYNeY8zlZGwK65yT0t+p4I3nmqsY04mCtsSXN
XkPLAmz8o3rXniR2NhUU9Ky1aOOCd5HSojIiTazOh7mBFLuw0R6tbZ8rcI1MJsVkK7xTNSGXecAm
O0mwzkKuOSr2dZ+R73rer9lHyUTQp2vJMO/I3gja6+hmgAuz2dj0j6E9OqMcGWjvWM6O7GMlFbtN
8tGZBOPredzOfz0Jr2+iDRq4cLyVoCHjWECnX1T8VQ1dRFTKp4cZpg+kuMEFAqsM8q71eKwrlC3K
1eGp2gpfc9kYu2SoWRuaYt22oQDD+HfOefUohqOW6BvVLuthQL/RkwhgMYFgZ30yAZW0qQZAbk7v
zzX3t+Do+CX3zdiVqvNy+i/oG14P88l+ldpXB4gjhhqcUk7gWr53PWLcmhe0sitGTH5Vs9rvC5fj
rSYXvE5hTOrsJ4S/DmFbBykfEWCt+5DA0ye1K3xz5uWUlOWkhdHHah6FOE3V3VsLfbcW19aV8DfN
hXRO/PzaWPI2TEV7qgk1Sc4xPHbXpui9rpIzB3woFElmGcXyL6Q/icAhOn6ooLEuzeXmOfUZxKYR
olrVZNAwfwO6QFFHcKxn0gf24bEU9btJjrV7KSY4Tmq6soyM9ipEBs0i1D8AiVnHreJf0h2a2PuN
2kVuFFjCIxt/NoI0OGDVy8AhVxqxOvGaCcOkhnl+sFAkBOSjWdziDqGi7XLl6Y1lY3TV+fH68DN+
Itz5zSzyJvC2GDNnjzNEoq5Ez/6W+i61DPiMr7kRlH8au5mKmeJXWgY5wOTI2p1eK/JKP/FR3Gj8
xQChj/BU5HK9BazESjCUNULRyvDxCgLFG/XqGtiMnsE8CQGzI2YAhVuQpWxWRIx71s1/iyiPsjt3
UwMyyMX2Uy/7ARYQEnbaRA7wLz2zvb5+wOWgHj3CDdSod3rRl/k9Ph/EVgPaCI4LHuUo1+kqA6v4
hZmlcp56xoRYq09OfP2PO22DOcJcaX0GgKejFWFUnAlumbx3wwj71xEdVFJd+yKO3B7KKtu55Uq5
3YgTwW8sv92ZqElbFw2O7aqnL5kIYfN4VdLm4CrAXLlTr2iVNEPi1LnQPc8d0IUc7djOawpL/Ygj
KCDif3yPkVKRgcWFFm2metQANFq89oXQjcynzGedupRW+GMQdwN8FMavDpqBqpAjeYr/fRBiXPMY
6ePQ1HntxkhCT3EdO2IjJ5xt4izI/Lo4U9pN0zavHdwmqLDrxybQY91VvvjoGoNaIR1uEfiJFHaa
bAq4tp09gHfBPHCaChChSROb2gywSAYa0II70rCBeewIag0/uOPjYHkTDwOXjg3cdAs0j8IPmX80
p+Usa3Jr9zOJr1/xeJniyVA94+PjCoZEeJkBbiy8qHhyvt7jnmw2x2TBlAsSrHk5oPnIlT5lrsJI
4mX6DY51yFRf/rxqOxoNfX5HlioBDpmCXzK3NA0vupsUCs4Uz2T0/Ru60gnSbfhEwuheiol/Yr7H
hysCkE8Tg6j0Q6Z4OxF+Ra/VqFHAGNreiZIna5kI1MUb9FYguG24HuMDqSgH2w44e1PgeOehMTFr
0bsy7ZO0p3qlNJUjZMTwzjc0+3hVWc+w51eqXxzkVJ29gvG61sdvkZ7hnrP0AjAh3IqdzLfHH3IN
jHe7E3uG7mVSjEuXUceXtvusqzLzpdA9dLVwyl8cPFOTvR9amoQd4phmw+Jx8hEnItLgDPjtJD0O
b/62F9p+HVK9Z/4R2QBDEPQY6RG+RNujzvI80pfN78U3vE+/KJsLw4RCSfAYzLCUcsm59EC8lOA7
j3RLR2I9/U8onvMckhfVGQcKT36iLhXYgLFI/Qx9Pm/hPUBsBFpjNZxEcX3zpuJupe2OCHfPQTRw
OA9cApPPptK3l6cYNmBl4VsnoKmTJCn6Hc8CCCf4NQyW9Go99FfLBiT4057VGQJY/bKn/HtTzQQJ
u2WoIyvoLxZza17gpY4t4EYFFyFogTP27jFroN3+s76n2KH/9lUqqF5upNjTYpc5PtJT5RdEvsZ6
PG4U1c/q1wGZHLIj263c18I3Wf2aVPjLND7Xt+ZPwzt3ZzH3PTXF7qgi2D0R+AsH9OHDx4gGBCK4
IQSUU/UP+D+cBsVklKqjSiNFziu64t6SEl2RkLfviM/c9EdPIRS7Fto5UsMr+MaJoIcD/JAIyNOS
w6XkSz746oPJgpAUjXIaCs8o+WdBf3Q5bI7LApQUBv5lCR6OPD3BGz1acMoFojKXzIoW+t5K3fM8
ke+3YKg1KiGQN2XE4MvjsJCkP/IWmsS7jYAU6UPnyoMnl6kbqol6753UEzgfJQlSSeCRnspjXVkE
Y3xnGjiIcP2W4C8RG6sqJgPfznC3MKLS+OkTXBYman4Ufp2C5l0S42flukGh4jKlkExrliSJGv81
e8cIQyFp/KlZo3Wh8CWN2O9VTH5gpmJdG9unI47rZxyQQ4S5pwsknmVPY0uxZcliNhBfjIP/zrUo
24n00GPEwsut6s0tVUh+2pE+Tr0/3oLusP8EnC/EHq66uqz0GU3AxQDgMfdzH3xhw8StYSAq/w1C
S9BgwXIS6TEeqIei2TroxLA8lRZ8hCxlcFfbEc6jO71ApTnqjetUiVJK8lOXpFvS4gkhL6FpGiJS
bPcXXaEL78L34W6XILpOHneE/+0HiyBiglMrwgeH7w0IsCcAt9X2gqKV+Vx3zgFnaP8QcMZ04W4m
BWO+YENuKO7uwsb+c4rjDYDyPZprkm0SKJne80vxxuYhUNRQSqlsRjXuNyFlL4wdwVezZExm/fs7
7fYNq5+Jo+GVNDELIzrozOsTovM9ZXpMGxfBirQXYk6lLCNAw9xGw7zCP/ZWBJTNmuZJ71pAuGrT
rK+oQzyquVUrZnd3D3k5w4qJer6fj0+KYFyjXwc5w3s//IoyzDQ7YiZ0ora8kg8wX8SHV4prPXT0
h0zctaQ0ntPRAy5OY7eda7BGFP3qcGK4OzflGTPEHcRInkO4zqRnzlFxr0ebm0tVLhQMR42uFLyo
WIeVvhkkCh0KQaP0fESeXsfAR8cyoK8gXo6v4akAr6e4QI8t11nrvNNkiGEu//a53SovnCHY3kvS
cMPATyLC5Li+XWNZ4/87ItqX+NEa5F4BgoSgh/QdArs28oECGPizXhjYF0Ner1LYeHs4fVjk15Xv
SFzEarwjGXUsR4fQtNyzNoxfMF2sKYUBn0kVzaKsFWOexNbPHeTGCBeIfDMCbMNBYtJ9dtMyjA9g
uFGIjDQOA1KPcWPdvAW61q+Inimmtc//FOZaPAX3Nr0s9zqEwQ1e7F2Fxc2P0ceMHIHuZXxLxLFP
NRqKPiCh+WeoWvlpjmhywXXt8goXbFfD+mQVK8HLWBl60LIjidIMibYpQDpWhGiB5FlAUXlt+5MX
FMXFi8fLtkBtB4XqAaIZWhiZ9Wzm+JjkKw0Of+VCYeyOiSFK0ozaBAqinw54Etb532No9ttb+jvL
aEwQqzxwHnNmXJ0h8RSJ4JHUXjUh0XvUzBYnKKpvNJeQC9lshcNRkIgjYxmsXW3UYZRfISQ1ZWQe
SGnf0+jz8yDA1LzmsPmPstiHeG0faNJcQnOBShWwrENZGvMB21IrmBEiEflLPGV70zFjmRn2AsL4
pS9J1V/O+ZozQXe3hAGPFdgTP0PQdFWV6a1QjJbG+rf3Q6DtevZIpRCe0H/R+koSFZ6yJb/FckpD
bOQtxWIu7yYumlA2bsTEzvEFrI9eSYzDXUJofQUBGgyxn3CmWcD9F5/6QdMQr30aL214xM+BhNPI
jTc+Iq/t4EnZa/1pRGdzI2a6YAaPiWhBncCAt+UK8uEwElqJRo43ZXnqvykVb37UfuO0L9iRyLQ+
exZXjF8+QV2D/ya0uXMYdu4U0SwO3Mgc/bHkqGKVb8TuZhYhWOpNdm1X/OkBWmrRv1SDUxTb/KXm
X/ejIsQxtt1YY6VOkVwfk+DtkGw82vaU2UZAH4bZoc3GKb/LCclX+CQrOwXpr9LsVDNGBgNhDbO3
LxMDo5Kgf4DTadcvXuQMQO191b+Cgcj25kAl4ldqDRsy+xedKYslg+QZPClcyKkWf18+eKWqOf/a
R4w30AKHs4ggjUHie6ihTBsCEAbglE/q0+czTMRaEZjL1rQciU2GQzQXNsvl4ocDglAT3dEuv1HC
+EF1RR3pyflcP7PNwoELqV/ClYvIQiBDfED0weWiEd0eKbvGodCEKhGUI7ChNz6g66YQAFEedCwP
RCFb4poW6y3D7nLIxNGGlsDHTYPaiIucipFpfLXwqnmjV5uDnsDaNtHJd9WnRnATxPFBvSRJVXWI
GKYCcJCFHKqAHjE6VZKIIvu9m5g+2bWGLYl6JnftIq+iIsH7vOENdkJK6y0PxerdGTZLrSQ+Chxv
v1MB1Yr9fMvByKfbrP2sXRCIXpiC3x6NXTc4CN9QAD3wHym4mx31iGB3P6HYfvuFF2/QxxVZsZJl
ahJs+i3zDsCyaN801tEa5uKPVuniiSm6m8HtizDgYqj0d7vIVtbvhJqn8hM4UVV+Ryo+7ZsKCZhA
o5nWKYNRRcGXExMr5h0ItWpeTHkNQI6DfkvEqI5971rZ1M6YPjTB0Y5gSy0OoesM41C1A1so7j75
6/ik7BYYMCYlLN7UI0JzdEhP3+STzwukcHo2L+evo6YndkoZWPL4DhTnjl66yWCU14WwAzH+HZGu
AYNJXlGdr4bCnU0AN4jmdrlz+3l1l2ZW8v5i15gk8ZaHDbQqFCUo8vOraUksyWNlpiXLHNP6RPUS
Ky0nRZzhZhp2aB/9jf3NZtE25zslkrY7dD5wfa+8oYBbcviYp2VKsbED83zxa8zKSjUV5bZDZfqY
raGM2fUiPt7iRkwZZ7HmZjMdn9BFOe8qBdHqQ2z61BriZV3TFil93M7LYTkayVukO6xRR1k1c4v5
IBNVqhMWyJplyO5+RrWU9GxVLP6LV3Xd+ALWJ2ZpKgFS7VFgr7v6aXwRGXccELOIbAzGr2rc8Vfr
WonyA0YCEneYGbCAekM+GNRqa/oafyVyM/TEDgp3mrKTKcnaWN4c8tsIO/Eis89CgE/M3Q2CZM6B
1DxPx8lsSwVaZ/aI2NoCq41wxkXFOuoV/HztJdoBHEQjyd+/urvNsPeHi5acUpkIBxq70UQvXELz
A885EqfaJwz1Xyvu3AUWVFggXN9MNlRsRbOoukFVwb7NPNfJx8HzhbcQGN7rxvu28m0kQThc1HDj
lf0gO45SzMk1nyOQw1OlthglD7lkdQ+Fu8PxKyJsT1nmU5HV430z9PMgRSShGjFQB8rLC+tdOW6h
1Z9SIMETFgglY1CIVMLDleaFNkxVXWt9nHSq/Td5stn82BEiPFxGmx7Yb8w73ifUUi8w69QGUHq8
1JnHPGK83JQcHs7OYCOHKm3zjA6cYkiodKyQKKvk3MHiro6quqqvW4y1psHQgDmQYTtpnczmPMsl
YYfJ/qtkVwHiK7f8+OB0muRWT5P2e/XTQHgan+Fp81zKWk1d1gShgH4nIq1VKB84YJniivWlucls
upfFy7mtk9AsH9Po8IiEDS4SKPg+2ffv1hfn4sMwrTId2LjWplUqnnox5PSaKSJBVfIHOsj5aKPa
K4XAdO1B6w2PVZIChAcqirB3J7L1W8jkgzY8UfoT3Hz0olhOdYnxflV6lSEFTzv/UKDvv7CavDQO
wDeI6on2idHBDiKEMukEXUDPLWx2WwK16MaWA23O3rlhuQOVdYgiW/5vODyYz44n4dPSuLDp+lBu
1VmEYQlWdvZZ3eh9Fquj/8myZ1+7KGVMYC/b4R78DWXI1l2YTIBo6H8xyke2z5qJmGaGQRyvG4MW
ihzz24CXDhMrQ4PaBGj2m8mkumuFn4DvK38Z63v1kHAl6EYJXbLrHSNTAoLYPidnE0KgKysdM3PR
f6jAqbLuwywQUistTWEtC5seuJhzQDaPC9jgg5c8SdSZbYpr8KCmQm9QHg7WguSm2HjV6scR+dCe
dczZU0F50AaLuTy708Nk3rAlVWTXVDJ25thNVaVCs+I2/CYXZSzB0WrPGhKFFen0s3+GmTty1w1X
FJGYiPwdNeuR5S4G3rCbEPB8XxI4geBWXyP9EeTkiD3RJX32L2KCJoBBblPJvoTHim5AA73ssWu3
kkcbT3AmugkyOPVvDZs0ciatNWp++GqMRxwpjbppibu1ha9Ql47MEboJFIn4YeZu6qbkrBWBm3if
QprnMO1vpMROokru66Fj1MWDtmMlE4ijz6AP350suPbh+3MRqzS4Ri05nhjCn4aQZVEbn5XPB2BB
ppKcO8viXHmzCFQV87vMScUJD2Bnl4OAeR+M/qasb0p0pA0UXpKu2t1JZEaO7RayGUQjE4slO13B
4oAA+3Do5RbQJT4LcTOuwFrVCteMezEHArhwZ0s8szVPYvFQDDuOrHg/JFXtA87UKvZWACW6F2vD
dJfjRtq20AFHdOxLMTxXw+mdh06Tg3UROeEtwtmvGy3D/scueNFBtadrAoRrvsVQEvRJo0IGpB51
51XmQdHKcQ9+sWDFe+IEtTA/DljLAmM1bDbE+HUHJikrlyvC3pQOyjPBsE8sjSbDiJrQD4XjwMnx
OdFWS+8uAGDhKMTPbsi7wIRVpFh3ZecnExhQRz5FQfufoH7yyYegMkXgprRZLPs+LMn+OBnxoXye
oromFSBZpC39CT0DwTLDzv8HpAD2kXgGJbfLkzNj223hkKtr7YO/I6nWjWjJqMtAUgHLkfdbHVPN
nqclOIZzy7fFQY2c/zs4A7V5+lyGQQNMiz1/PGsFDtZ84RoLa1m6vZ4uP3N59YIIvrmkeRCShYgn
mrQ4J3X752LBkHnrnHpdo9ybPfR7R4vjxzwZ9R9ImvL/DZo6fwsVuOXJsQyRmWVncPvnW/j7x3O6
Taj+MlM9xK+vEPVuWghGn7lnV3e52zYo+a6WxWQX9U85x7xMfbJHNEBVR1f6JDbcMQcjYyN2gbSg
3TOkdkHlIJOY1uptk1H/Js2TDzZ+C7kYq1/bSphms86Y8kr0QaEhPRo6JFjnnJRvPYe0jG/uliE7
HpO0xoyXrFip/FJmuptXbS/J5BPhLuVc410Pm9/kwwiihis1LsVAZhY+Jeuzh3M/6xO2fb22NTUV
22EZKCH64PmZzYSO3YGppLGMAe6fa/2WFDFJrw1BcDkMeGUFGF2AQFLgkEy+hz5+45uCIBGrJgwe
X5W8xKorz8knqDy3xsegMBN/H2dVZDbncZZ56HlMtS/1pBCeJCqwMk5zNddJsgJwwjo177ONq/47
PV8fYrSap65FfANEyWn8EuHrXjAC4UVoprI9vvNWmQhw+UM0U0ct0wluPf5grcQ4AaAWSjHRkiOf
keisXVaIa4Fye2433uL6xxf52mNblJvYJItDbMriP+y1VRuhEc1JcP5vXDTM4dFMca9ldlAHxlVr
Hi1QzeFYq0f1PQIOavlEZq42dJg/ltrfZGGx562ka0VunjYXLOez3GjUjGhIKtsP3f/P3BQR3Ip9
PqmW2U56cq9MGShmD1d+4sAD5apdlzTw27wjfzzRvaWq+xcrkPbCAMzamIAdV0eO5c9rkRF2Vz7Z
+oJE0pPLfREkfBbiPbqfWlmsUBubMnzHp9IhEUBj4Q7qL8JHborrGxK1uSOei6pcCKbHfSNjzCl7
mNRZEOdcBlS1PfG5cNhPtvJxCtRwllIWO83lGA1AjGnOTi0amFwMtOpYN6Pby6fpje4yohAKrhNC
rtv8A6yhPY5G6r4lME7swcPzOp3JWKU1hMeA9LKU+BZpGOMl4Y/p+5mh1j3fpjioz8q5Gml/u/Wc
lGFIM2pGbnUiR66Q1b6F9GeYSEC/sPWentOZ2O10qojGoTW3biOMLCP/tgWo28O2E5k307+SyRK6
oyG7RANAph+Rq+INUPzhTCc57Hg2sCkBCxFpaEcYBhNFZF8ct+YMy98T8JFn3rQY8WQGw1IQWM60
UZA429AG2wW4nYzFuUMjPzao/U/ePhNTF8ubw1QBhYZ6Okv/XY1cJxNNuNV2BF3S+9+8WQDJKgaG
0nGeLBehHW5T/EDjrrpnNVsuRp5fc5iu+5WQ4Be1G5QaoVduxx2QHns5oeKPPQqypYr24Tmku3qs
haJ5DCBur2N08WtNt7DJ+kwgz1dBABW6xBFvnTslVucwWlWXL2IIJ9tTIX5S0yj5ODrxiCOThf2t
M/2M6k+h08xi/670ntZ7nJVAuXNATvqVA1bdJygl5/3vf681np1ys9P+KLTJorJxR69rxBTEBl7S
Vuf3RxpYzrK28BNFWYgs4bHnq97knyV6VZyGDjTl/WWN1oudgZ8fHyY/bj/xwcdpg464BvMN2fJg
Ra7naibs9dnSnBG/CQi67nv9dnO932CdyOQpyC1zcB2rVZAo6vuvKQS/QOHPI05x5QqXmqBpS3ct
3O2tTJ5lTG5qu08RYiCU58bMlztlIYkLq3RETy7wl85Fh5HE8VaxtDpqKkHIU5/Xb0rav09Alihr
QMOcZHhFnEh4cPwaXtp2ObEvs+/TBDOad/KNX+TWM1yIi6AUXZxa4FFMfKbO+zb4Jku3/ybWT4jW
gBW+M10mHMgvU8/b3Gr3r0yAkA9gTB3SEJ9oJoGcDCMfJGJLi1edbcm+12Ne2sCkzKb0tmRUxI3m
1/QIgMAFoIri98Oyv5cveyA0UAeqv8XuV/YTLpouEGHsX6ZqOdHKLMJBXvH8NmaKXPrSxnX/HbAW
7UZpW+ebnz6VGRKTKTvPB/SeAptW2OhGLDPicON69zMKucdWZ8ePirg5uZEA9xCQyz003wt69xqs
+57wdtRLigi6DnLOnmKqnaYNdJoeYbO1SrXibhgWDXHhvQhmrOxWK7CA/iCqiOEkksh5OPMbf7UN
DZhgNxyT+DE9cZwDdc23BRdScmtMj6QU0VequNPQK4fw1NBHxr5fo0LLcVTto082Vv95Liu5IYhf
AoXUrNWSW7C7+uXvqS9sv6foPtIBZfhaVJeJrc/nrIr0NxjHU8u0nh0FQVer3pLyuHwR9VogzFHy
VlVAeFUbq6C1Yh5cePdD8nC2fZSsYgjOht8J9+7HvIz1XBErUk/R3TP7qvvIP5q6cP7DJq6jA9K3
4nSHa+9Gd2nyl3u6rboUuADtNHKrpsRzzs/vW1Ev8m0N9uNGHEoVaLcjiXRIZM8SB4yi5WEdjFw0
2TCyP4UkPeyjkCVfxUswlc+R30K4IRzVnNJJOlezXpX+xvzsrEhY1CaJwmkESTCM2ze5EvhzbsSH
MV8ZBrXqeDtlmwdO8Jo9Y3iz+InduZsLZPF7zP26KAZ173G0Q2AnLJoJr3Q3W2fONj7yeHYwTHQV
s4ZNhus5+q2s3cGcMLXL6lGUNmzg7qVa8q76ThNBry6q1IWrDNbW41h95r0kiZlez5wa5c2wXnpj
ayNupasC3qEyOS1r6fawvqyoIpNfyyJHuphwgkThqwRs6TJhFzaC6huzD0wMDMv/bbv6fm4YvUUK
npVhwZpeGdc8DCZEV10LfOdxBBe0CanWjp3rk88ZmpDZuArFqMMNXVfqm2jDp6qRf0DHJcz53HTS
JDMHJtpFO94cykF5Z4wnmsPRt4loI3mVIVx5+BGilPYu5RN87hlER59lNjJ0kF3CuMJItK1TOPAB
G/VbIvLucmc2S+yLYNIOAnLxcW9fx61jsORM5soNZh90kQ3SymUSJcRopHlvVUjJRnTVfLFNTTfT
4OvoEfHy61Th7O9r15lzNmALdh/EOVvZQZ6mxnZoR6T4uafQamxlVJ3sQ8rLCUk6IIp5lRz2ItUw
S4/PcJSIgPEQ6sQKtk/SoBuWnhk6q5aFVVc284XiJdT2mvoBZOmyBWvh3ltCOkyoa2nd93bXLer9
s01BOMo7ridrz7Bo4j3l/18eZcZoDce4CAWV9WMqEY69dfiz1eG6LlccaYLQEWLHw9DNEeDBmQ04
GqLm0aqlUJJv/FKWISukxqhp6b8RBdYD5aTWHEAQBsny7N8BKO+WBFphstCrbZ+EZ+bCYI0obR0P
a6DB798BVR9jHl0aCe7tp6bbluNHn3PVpieWl0U95yWe1jYTIh+ZfTnp+4G1x2BvAP2fwYHjj5Ms
ttZJdNQVHc+nLdtnDszCDQ9YjRMp52vpsYx99yR8Cv0Fai5tWSZHDrDdjCiDHWX5N7nA61IS3pYq
+EluvdRycKiX3EcdzXMaZWue+ZpgGbGunWsEheYJKx1vCe6R802JGGL08isDXNC6kwCgoEpor5L5
LmmETYSaJ2Mp4YLSme8hWLznHOF1hrv6aF51HFphYZdgbZMd5migF8g2Oe4g2C/NVIe9e66xbdFd
X2XJtdMYzTSvpk8USuSGcwMa1LaeoLTVeuozyZvqG/HAimS6v3PQNsngkFRaj6peMKlS0PSHP4pO
co587+tUykP8L5h65o+L6gwIUwn3I/Hr2Ibdx2/vf3HCbwhUdzAChjiwR/eXJsbo+M6Bystn9KVV
fuduFa5kW91yv7Y0b2Ij8UKDjZTbs4EU8chGayIZHDybZ4Vbahrto02lXj60PxgOO3avZp8fwFm1
C0k+m5nOWYwXpebqV3nx2V6qO26jfJ7dAiMBMXvCsLD3lxtOvP/kSv5M+DYOKutgMlzqFUaKfKyM
jEqfFzWWePyzzpEfxUkPlM95Y0KGxDj77ZsoxrMoApByrt/trc11iUg5BBGic1I+tT9jKBIOPxTp
OGArdbF17aLYHvI3J5BQ/yAx6jJHITs/QhXu4XizmYbOaS57jkGNqhuFKETfT+YI40j7ULTgFZjr
uWCRI/zEP5IHfdCbCzJ2fsiYeWGHJq0eK1V3LtjvDF0EVcemNT+ge9xllhMyYCjmZBMqGWOQ2q1Q
chrfTEHYvS1cWQ+mG3jLQtwNo2kTtv3g4WaBreq7nH3FLJ/EEdmTZN1qwNo53E/PbD80PiC5wf9q
Csw50sPbm+hhOoNoKJLFzPZAqbT/LaAkv7hepnOWMt6/PXXUzwgOxphuaIR0O40JTcqRkD4A4Uh7
xf0kFY9f3Oj36wfCp/S3MYdwVgYLsI7UIXOnyrbAsfk7OKqpC7HkGuvExwDIfNph6aRvyLX9bBH1
0JX0XvCaFjvPwh/QYPvwFhhzEoGOAvcjZVqqzc+RS+wl1UC/QzL+xsm9jp2IFM41XCqD90Q2yA4c
2ezVWdJYC6uOB6yFfJX3jhZfDpSIkg1vQQtAaDJhLsor09dzHE+509LcAjnLpUiNPnyct6KGuock
UoVJeiEugVTcUkIvL2aMZGyBjCknq2GyNIcEVO7xztCzEFDR3kamHKlo8L1TNjsqnrDVcCKBudXy
YQv4Col1alkwmi6zRBgqUeH2PgjIHxDRa9djW+GnAoFh1P/pYPpdIeqp99AI6/9AoYmXLuKctDke
mbYwQkCYNTHvXczl4v/XELgt9M5b04j9bI/grTLVHn4276eIvod2D2PAwxnGOKRuvAt+RcS7EHgY
xtyR9eADoDidGv8fQ/Abwiz158OQGxpZ6e8RtDvG034MltmAgwqaPnoNeM4Vfb8apTJpo80/3GLM
HJuQYJxgVt4FApqDFsjhbCYVfeKTyStV568DF9/H8K/s9oLTu2jgWSSRIseKroIf1shACfgvRZDi
JcoeDyH/t9oVZ749z0WmntUcbW9vyA+bJ6ylYwZjFWdp8+G+G7g0rAjENZf7DkcfwYbvylGaXdAR
OE+eeUozgQgvd+zXH8j2Diu350wmjosscWFlxaUjvC9OqafozpGb9T2LYEHfXNJFFduJFAz0l+QG
W0gF4ZiGTPBgKRwVgffCvE8d96hv8z9vtrEEakULDwr+wU7PM4C9ljXU5aJiQgc7xxARcRBY2n8I
R63ZfsRnlQHMooocE7PsN92SxygbrCY82WOBLUKT4jItlfjoMvx7hcDrzF5ToUrIL0ss7Bb884zj
EZbZ611O0mPm6tfxqtcZFxFkSj2MkoMF1u5QO5Gv72KqaIOuPGcNfImg2Cw6W/oA1kxyAOQXoIX6
+i3KWtWfvXwHAHVrzov8d2mepPvE1enrehRFgKLBibqj+ljgUQdPH6H6WnB4QybnXVT6eii98jjD
ikMCVBHIIOUcNZbGI3oAgo1pHdPoBBdeTQqiSQKrmzj7xpE86eiEKNDbrzDvOM+HY2dzn4cj6C26
thZPpFqSUJ9w/1o4+vdROXSxU+LxPMmEsnL4EcMF4BtoW3vFYXTQd72BPBhqnF3PCd/MfSfBUjcf
Fz9ZYgNOitUu761CeDoxki1CuaciQjKiXKtwxT2fNTDR5HeaAxV4VJ6uK9Gg4Guq8Qfoblo3tzXe
DhQRyAx4V7cZ+m9kOrF1APJFdXY3B6ilRvUUOkZ/sCiOiddFX7p1LG7VANdSZ1f6fXBZD7tWY8H3
BIfo5ouHldORAMWJpV/PXHoLZdiP6ZNH7Yx/3/G1SU9htdj0j88QzOVRfEb9hyWCRK66f60NVv9x
JHZOZJkx7/lAMawOYNBOJpYdnAeNayxMaEfsztI+7dbRifhKOluneUjGaTFcvlpkfTNZ80HWxvTt
krs1pibqna9prWtV8AbbZZZ3t2H600Exc0BTyRVFZikaQeO2fpViqv9ENN9rwlV7OOy3TzHswqRl
byXkhui/NGZOXJbxZAhfUa0jn01dK2MIRUODCXkTnevyP57YrV5jafO2gtHITKESgaIFgEYF6alV
i1hVNPbITYz5zhmqKIAtPl/RjDxdS8kQDx6q92WlkwwOXEMOxeT9mb5MGk+14l75EiHtAfb9INiT
JBfGdiT3/+wxr1msOOtYCWTsjeoH9SZJkiMDb0Olq6br9/ooyHqh5UyEsiqKoE/jpd/bG+hMSs54
23jO+NwW/Z6dMOba2Izku6DnY8ZN8EDMtxBvhaofH5qV9OrktUjIxHm4QKtkKy5ea21iPH3xhUGP
nG3P4fRGY62xGxMJonFvnjfnVJgfJwR/M3ecKbG0NfFFtpfXwDxxO7OsFwqzlaTtfoDUdfcUQfkx
uJvMiTzJNBrdxDPY5gdedtDKRhFskmGB0NgCGFT/18bIM+n3/LQ9HO+Kfh3s9uxxHUW52OzJUeJ5
VhbAVMipMFQyZxEF8ZE4xiZN5xcS3V8cGcqUIn/ZrF6352UThcWg6stF4Ck7aXGUD3GQ/yefj4IP
nXkYGOxGkXmiTIS5JmMT2QUvvi1RPw9QJHjcpZ19hBmwq+ILgM96wR9/PhuDZ2QFqlBb01pDX8ot
vvrFnx8CU4skqWh5bqiYIpnyj0ZPgeg4+9QbSssx71fxqsFU+IIHZF9+zPMxMvnuOTRNDC8bMawq
7m6VqmmIFYA+6C+J4NZ07KA6PTUYjCrrbca5Yzsn71PoF+qUE+tf+11lvbYcda+DOo0BaSPJ34yI
9owJQmek8oha4aeStTyq+RfDJpNCyn0h49V8gV4gmPhc04+rBZfXfTOAXWVhxAWt0DFkcDFpucdL
7CJio1YPPlPiybJgZMS1uoTlIkDY/wIbsZ4ZiXHWP1iHU++8Ut3YoqsNPJn5I25ZjRHJB/A9/0nB
e9DJG4L3iyY/xVPnZMb4rpvRdwqZw9BWO0V/1LVw8Wx+5fuZzQ8eT2mle2WA7fu+YVDcKaVBOVsu
/Lnle/tLuzzaZ05nkxwaohFYPwedutiYDvwwgXPlGNZtkuo53tODN99oQQMfWJ0Z0545Ze07Hb0k
Wab/gxfTmau0h1SDiGpYMOXDg+0/3HlyrmWerSS9xpWrMlaplS6SHZLM3i7yERLR8P31aA3xIB2n
AFs58MIgsy1YiBvd3lWD6qRTx06bLfk7b/x68YNBMnwCcMdt2+xYuSU/iCpUxCdK5iSDRoxdNGV2
G6BOGRwAFwr/RvvGiiw0wIYhK1sJQIglExiXGYCdXNdqxUYfaRgbjVBm5UP8WDNsYGNOzNhy/1G+
SVg1B9lwbkh6MXE0EuxHbd2WuN3NWKrsGyjILQw+Ex8zcJAIXEoQzV5Ws2lnB7tGVEH/VvshCMKW
hT1VrxS+AxXeWAen+Xhgh7jp2YcJUK1xJ+ojdiNT80zEtxFIhtaSFwLCat2UHf66OODfVJBfnZys
k51qSBGH/Rs79stIye6inuiAn8RxFnKuJHzYw+Ztl3RYCvShkhAazKpNDu7cZ+1uwKYr0ol2AxDt
kHfviRF4FM2oizhJSxsjjGykJb+gwnvfextE0qebqIAdvUviF3QV5wZtiiALEsm9RjoIydip6tR8
QNRvYR0nDnhrxOtiM59J/b4C79ND++Hr84Zsw/pfjVjY8KkSo28STQxiZExlabuDaGr1xLNKLn+0
VR+qyGyBtLdEkNsVXp5bC/Rkgul2DyxBg8yguguQT6gLTRm+6N/3l5jkJ0eeNqrO73MRC/5LWgBM
IOLI6IqaDqOQ1kYRbU7fRmdnYUxFCKKaRNCnJqM47BWTqM64xCPAWhSa7+yFtg5rxH7DOnto1KdS
MuZSXdII1d6Wax7YR+EsQbApgJchpcYadfCWDqYWPBIGGTd3/lUBMOaBqDoumNOMXA3eiwnak2JN
Yd9TKW4lrsblcfiTByjX47DAfLe4JZic+SpSArVpHEcZZz8ot3MD3oVxKHLNXh+BN3GHJWdgxfMx
PiBly5Ur5TD0GiEPVnla9jIXAB0susFtqc6cQU2Rp6PATvMVk36w0uA6XBl4dEaFh7L8xaeG4Bt3
aePxR9rPjTC/x8OhwL/oqXVRv3OHk3PsAOyBAJ4pXDMxHZ966So5I813sJaSP7yqmAGP8LodMEBK
y82/uLlhHAlHDMgKf1pccx4gNyI0WUY/rVlk2kgXmTK9RygxFIxTCD8Z6WqBrckqHiuhyPHrIYYj
CUp84zbuxKpV49vKW0UD9cr39Cw06AIrmNuKDeWMw6fEauxc77C9e8kTdx4KVLzMzOX+b9rWhnzk
cTLsz4vtz2H5aqCjzWPQKFgcRT3p9ETXISBzWDEpnybVnHAUZiKGDDALMi8AeYfpFUyj0fAjJIDb
xCWa6P4JvLRRAz+nnbJYqQY8eaIs5DDx7yfzRbFzjTy/fqivNvXXyaw30T+E0cpZD3oa6wnFWnGh
FTbAbOXADEocgDRzEO8NqchrEEvPEJoe+9x72cXYXnqYGwfBTktGemUohHN1OnI9X0PxOXuzp1ZP
zH/7emXDVeO29f6by2fUubOMFUnHPvCj9YytTQJPAsHUBy9FV9gq9pba3NPGHFp3PRmZMBf82qGZ
HGvxNyLaEqbaQ8w0gBh19589xJVA/k/mUCFnwDJwzJMKXM9TXgHOF6PnI4TA2NjOixmmVsgx4TP8
QX8dkwmNwfIfkoi/pBYPhL4qu1Wog9ODmySBk76CxeSf/j8XO9oiemY6Bz+8BYVtdUcfWGvedRN5
L+0hLww3dMbWsucNCzU5MARWei1/D/aPjOlOC59qIDQtgKF87tbZko9+O6VVPp5vWdHciHs+d9Rq
9z0uulTOLlOilm3w9NM3q6GlX0u53O5GUeUmzai5CqB3zisfDCBYj4bjhDeY8QAT44jzXcbORgYO
mjNCK/PX7mpUposNY11uF74gUXfZY1dnyWRhsjZ3snDkz3V2Z71mQQCb8X2VdFOMUSfIHKAKfoFI
RBLgN9Vb4v1jHSXNxCZ+UJSDAwcjxdIP2x+0qGYrRTrT+tpE/r4gM+l5+t43zWSzQkh71S5SmgYe
j0WVYBG2vU3St2iGze2fznsFal3grGBer4YmgrdfJxFbP1N8tK54mb+G9xGAfJvC2HMTB/gLIwMC
ZuKE+hx5nMEJb+RCIF5VrJ5vqElxDh740L27MU+Uh/wTFo6aYYmCgTjW87ORG2y3l4zyC3rIPSTJ
EK77aSTbAfOHpEZc3yR4S3hmxF3ubiP94DMhgC1iZ2QkjPRO/9I86UjdBZvpZ2Qe4akGBmYMrJ9L
jbmur57wXNTAx9Uu3ClOGGbbnVKYWbIB57fGKOOF/hLufScI9JITK0QMw/WFg3mIIyis2UCKuusV
n4/WqQXsKIUHnkgfOiFpXm2ocrAFUFYzm5UoInAcZs6MyX60g1iP3/ign5jBtM+gxg6/2TRa/l7V
T7W7dbdbGzsCO16E8GpNddGPsmHU/i47KFg8QOwBb12CNmR7Q62TTg4mYaHfQK9afCYuM5DPHmM7
lWyC4uwbisJlOxA8pLlemTCUN8JS8gdvy4Ahj7YfO5mMR2Aji7UKF//uIYBRN2s2K9KgVlKpaCcU
lsoOGyG32dg+bGcMt4aCd2BWDlafeBijKfkq6JNuRlmtIiofmthL3iOio2s0BE7btJPeILOUn1Vg
qlmrsNSl4CMI0icRnzzNvOmeiykJAvrHvsy/Oo92iewH5aNYsLiEjsC6S09T609T6E9WTAmA1+F7
qQ0rOGyHj65BpsTAtPYNfGXeXjvVnHlimwRWTfcoBPmZTKygwGE7w3SQ+4Nvmc3CFlWFVfep4TRr
EfRJfi2Rspv8EjY1r3GSpZTgsxCSSo0bUtB/32qFrYiSBpAX3DE+ZHVUIv1NdAjhBv/qR55Rp4F0
ikm14JpVJmyEM5AYDnWyGrfxee2kxPFIuDoiIbX8P2XhIeXrJtvwyCJeR58nSMy1Inxv4sqw4FBf
Kos//7eOMuHVSOkse34YVumKaqmKkdmvxze/1ndFKTNb1gduVNDOKbn6m+nJtGWbz7ZgmUiALcJF
mpPV4IXRicgeCaKBJMEVLqI/kv121caFApVbRz1fhM6kb33dyi/WuW1lmH+Tu3urMVQ5XO6yuvpb
JUVIw3qZv265hkd5GZSnBAIId0x1UBNpzvHvyY3Lbp4tFCw9LHt+/mTy7S08Bqn4KEGdHMswTkFC
/Zsybjp61wPVzrOvksB7j2iQm+Djj/Ii4KMMeu2TeM88GoaVMY0TLIRXWhDSmcflKnkwhShP39mu
wxTjU5ak+Ri/beL/njqz3cIgf+inhdDCQl6Zqd5z7Ui0+ouhS/qmC30n3oClQiyZA6nr9maeNekI
FFpeAYgPkirIclz7ekreIuE3hyIyU0Hu8RZBlt5mWndhpU5VLQcJPJw8n+UMus6VQIFDWiQYy9en
Ns9L7PhtSYK4WIPcEsrN9YYiVZ4OvPLbwbWD8068MHDWlJ0Aby0MMQcb1Cj67oHSIpiagd8y3sJc
sO7u4BHTkC91Q1yNyxESsshrJ4olT4dM0J1vADnnhS9ojZ4W3WMWk3LCU4gH1dO+qykPvApPxMpp
csqUjhSgPq58ZAC+LM5v6zRAKYc+5S+du71IWt4x75S5phxtxIE2HrDhYdt0PUGBl323QlfvOHzK
BoB04l4MXFVgpC+4d775j5UkyoxKGcy4VI/Z144nQXi+vYePVGyc8rqfa0PaixJLD+AzecfJZZJj
JrQH1puEP9OPek3vHrAKVMap/J64F+/NVINwxngU6QVSG6wTWCsCUgyKklkXa1kwdJv37OGEMBBQ
xslGqJrGV1spJusXypb8YZIOx7ZvYf7e2Bf8y1+l/XhiDNEgY4xZ+ndAouSh+JXByAKnN2iFGgNI
MFdqU4GZh6wxfXbNFf32TWCFFfx3WYzPwIukUhqnmpFWOqrWQcKKAh2/AnL6WHxYPIRWNtPjb9ZI
iGNhrG8/H6rM+/6eWuKNGSPv8zRuG6WA10kN4Vfnwp+hDJJQ6VkytsjPUhOUrzbbanbf1Ow7X70T
scB1OR08JqEjrC/72wJmIp+hP/3eTzzwLHKyI1Jg4smAm+Osoc4xpBtAETwMz0q9uYexOmkHAIVm
jK+u4sflS1xltAMUwKY0zJkV5G329M4Za295y3dlbWPuRQrvcdh+hl0a4eb366UYjhbvGwLjLg4M
clyJKxuceosxcZ9w2fa43cUHKa1tJAuUj+bcopTnNQai1m9YGHi1OcHOtlzNWN48KqORrVP5Euh5
KvCCRcr8nDX35vQ8G11rEn+dZVvV14IVhdV5VIvQ0+hdKSa6IccjagR1xR0p+dSTtaxQaLY0LZ6k
LMI9zECTEPcSHMnI+6Hl3L/eoacPllJDQuM5QrJ6z8itqqe7dTN1SO6WBtXBapLM8iqPuzBHKSiV
txUbBrzB991bYObXQAHm5CoCwDVkHE8vvhaHDkgKU+asGRy9MwCqZ8BBqTp7qECjb+JVsHJpLNm1
Fwuol3eYZsnV5OXwUhByc3f5AZw/qJSJ0El7Kzpf5pu8scZnS5lO/ISc55pGQ46KQJhCLQYVAN+u
iD8zz93noM1F9YOF1M7U6LbpRXzwz3/KGPHgjcjuvIM6achFN1v0DTCNRbRN+ggCd3qKUBOjCpoh
P9QUmC+7nYZsrPZup8Pc5Uyeu93IYnooHWQZe1PHZuhkvQWBHEeTs2SIfgVJny2gWGc9ho2UnBFd
U56vLFkECNN+Sy9pVagFiZlUwkx6YpB6Zlit1DP/BBRhNaJAiMQwjmM2+KSrBWuSqyv1zvoDM/RT
dOEE53BeJEXk9eng62T1H6GcaGfdXqHZ29t4SI1mpOHxcgye1+xRcj5zhNjbAWHaxPOuZEO6DatD
Lytw0NHpk3A8QBG8yeWANxUptwDSedL3CHcuHLchmV547wyT+tl/Yv3QX73An/9pOi41lFyqYd8R
5MkCJH8LSlcnIS+Bei5cUIYOz6HK5z3tAKUvUKOmXlStcuiXYIcrOdnBqeeAmLZgROLkQQp+QQp/
UnRylfYeeRcKcNmYAdLDADfPq4LNK0tKwBFOH9uDLvKKs0LTohLeJParMme7oP0I7w8LrOtGSS74
MELOFtIf7yE+QppqNap2AjTYoARwFiuA96W+8TWKs7cNUtgOIwNepYggDEOl9GUpfubv7c3S0Oi9
rwmxtQDYR/thuG74XLesp5zb4xCSiZ+VAnOBSVXkX2QjLggmDdWpVI8rpnYfDuwlrFRhDWLOYrvG
xFh1j+FrVkcjDxOcYWfnCbMjsOZ4konaka73tJyYI/3v86sSxbY/+4cdvVMiTgVkbmpExKDYA0uE
M9Mn3JThFjpa8YfmKUX8uXUZCCiYiyq85G970EzfASXN77X44mAKAJV7gI0GQQmB82/9ODsHAFeH
pRIAkYAU0b1Oe/V4AEqg98oHwRRIE/GHX5CLnGuVBe5kUXKVRSHAz5otPLmIwJZfiM9gX+YBZPh/
a2UTPSh7Iu2swFbMHpCMZU942sfYr9R4/WLrjmIECNhYpudCcaWdUhlwIA1dH8MSE97lFeZGL0+v
nUJuOPnNwKbl90J20erU4/eUCdyYgq4EGGA17Uaqsdm9soxqoRcIUqhnZ3Ke6/XTy+UI+1rt+kTn
E9zVyH2W3Yzg3qAWoYD6NVMYG7XK014/3/Xhn+ARFdv1hXk44YQ+fok3X+r6Cka4Q7ul/N46jhNw
x78rKj/UdyWq4lp/QakLv6UDFaLC2g7M//7gi9cWzwad3sbsyyqo8Um7xcju1DJ5wsgLyxwYvlBm
vgVRbnYM8GdEG3/6IWxWf241qbrgCQtllSjOSIuHXOzldAjjqNWIky5bGXlCkiP6w+6vNAY5Q8bd
/yWfa8I0UdAKS9Mc19EjNEgnEM+uygMefYBjnEmxkcVFcKUfk7PVsKXOvD5QS8ma3o8oP0u3iuw+
TAnb3KgVVzCteQqLXV6hhTw+raZoHGWbDE7zYS/kzfAPPBJIxryg81UK4Xckw/WnMg3H6ViFIyF+
HWp07anx3TPfm/DfyIQ8Ult6ROKarYgMiLA7EcjULC+y4jitsozNDTvhYMEBZuezlsUepGloUvMG
YF/p1fjPpx7LQgsyT6kqchIq/9H4Dq5bQtbAvLKJWwGEHnaWtqLjXqJ4ftVA13WLmWdppcZS8fV+
NJdZqGlXF4TYUFiXkQjKJhyNbaJmlbhWlS8C4wfnh9Cu1tZHLeGetCb5WPBwmqhIOzU1mOT0uHMz
/f3tcBnX2OqgeZylBp3kP30LfM3mU5EwMlbyDXr8JjekPzYCU8o+peBAhYoEqfWh+R1vgHTcyDNK
DfbHKLhgCk7A0i6Fg/PEDmPxZHkqC4Rk0yt85dJdg77yWVzSP7HwSOvPigPdmkAuqN0zObgGd4IQ
URENsdVTMQg0B11iPf1XHGThAL79C1JwPr8o0u40gqBZxR/NVhaU+86CKaK3Txa4q94quUOmoP9K
UbvbvxMiF4bMHdi1mmE1U+XBc38+vE6HAFCHOwJNLarHuRF/iekHTMN/Dffya2SJQ+uxWxcLsQmN
Xpmv94VyOeATYCelL/KA/GMf61mdjYtCbiJkjDEVWirVL3OSJ3qmxsD59FU2nc3gbVnGJEaaipKu
PdGw+VlgOTmwChtGGUSYEDZLzJ+KAeMX9g45u7T/QR2h0lCSl/OFStGlAizJZ/DTNRIOJghrj6rg
PtIss+7y9CqiiJUwXj1jANf14fXkZHFUCCqiNhUrIFWfQ7ndrnpdc40Mptd0KvlHf5yW7GcSx8G+
tnNjheIz41fbE5EklBIPnyiB8os+P4QvJWvAEZvm9Yt1wyy1PfSYsQXe3WKz0hRWyMY76/7mcDHR
7DRs+OTWXPSg5HSYQ8LQJoqhxSzm50vXT3fXdZPfOsL2Kd35fLCQn20yV9K5VHuHmGzo6MKve3Mu
ZEYvmhPjB/KPG08SWYpktwl5Hc682L4gktb7c8T+4Eb4YK/96rX/LiwjlAAaHJCkZvwZXgY18Yys
yubv7nSsHrMvOP9xNLSqYA940dbF3zjvsT4uH2Q/5j7NuaDYcWL45PdNZK6tLghUGMT4cV299R89
QpMlj8smp15jUO/Pzv//tDHl22McLISlZ/Oq1LJp96qKKYWEZMiyTtSh3qgTxJBAcY2dBDEtXCeL
Mu9ucfXM9Nb6t6ce4MAQj6/5tZvLPzdxCt+RaFgIm911yxt5LOSFXDXGaFaYh5T5nQq7+73nsIu/
qSerGfIgjXfLZkcemU9bM6QoCL47nLOjyQD+zKau9MG7Rwxlxs1sOORMIua0RRxiCB75PGho7qJq
wWwPrbivufRgc7Mrb+932kDeJsZ6Rta2ZQlFHlQvFDKeW6K+BRlrKeKINrrSKAyexd04D8PxBPnU
gG87jrDNjeFYR9MRJovJtZ9kQghKe3iIi1/8dxGa1s/0qyjoRLRy1IukNKKLNS+uRc3/cW+C+AJQ
R2/pJA56Tr8tO5cjgQNBBwgk+zx9PiL5ZX4q4MGvH+65Upv5wNY4rPy1CmDo8g1hXAaATMfUAewB
xt/ZKyjfDMuhuqkRqiFl+HphNW8ctJKR+etar2kOP7ve/IhAoRdtegXeuKOyQNy3gGS54E4P6cBp
DjVB+8HrDWT5R6A41QyAWGQsLN2ByxFVXMx0+QkjhScygGz72Ln4SbVark54vVAuvDf0g5iTHrYm
6ahCoGCYWYewSSrg88tbdjvHAh07JlEltGvqi4ekMEKK5zLOXoSNxUBTVKfkXwCaexcjyFfAA1Vs
MoMYG+0Cft7yTcrwaGWi81pR0sv1GRKUEwQDmAwSSH2QGpv3pxGwGj71qwkMzgyypyT7sS86CZGI
dRxfwLlOTTs+qF1Ogtc4pyQoj/2iO62ymWcMZOTLQ6ZJDC9rxzIbQy2GxY+WRfyV8Mi7mKbztso+
b3UiyghNOHZ8NsmzyGL/TzLcLPlF7UxRWE7unbz9j1DyFpka5e7HCuXygOc3gv+7GxiMwwVaWYb4
+MW7i7GrzvnBHvk6dKV3TSdxE6lOsXV6Mq59yvva46k4VsBC525T9riAPu+ZI6fwmLEigHBYFHav
wzz58VR1lcfKAsIuMlF0yt7lr22hcaccU2nIgjpMWA3E8vnpfGLvPYfQLYEENHDtG+A+ObK/GC65
Nimp4j/Q5m98JIk9QmdlR7InAD5e0C4dElpTgqRCkZeKVkehCgSzIunwMYuccZQHtB0c9imIuIgZ
Skoqy0MjVjuYKkSzjbIIljqlLwUCj560Y5oTzpQ99+CfY80DCfpOgMLbFqxwUXVI0yvXV69ef6KE
O50xlQzHY6URbeOr9AaPATmIdm+HwQKYAb9L3FaiiGV+79yppfgqGuxopk8uzvl2w4wcPzCVeKc6
z5G5luDS3vEoOKAlzz3TBDfupwRkE0SzV9DReDn/nFkTLD7HYtoma35X1HswwojcVeAAwUApsN/A
SH39RQKBaHvoqcsMFUyz70AunB3TtyXesWngnal3aEc7wKuLBvrhwOnh/Ex2EOK0Biv+QyUs+bWi
hACvVPNd2jrLId0qKifs+wCWPGQIbsR+hY7xSpU/w41m8T0N5FH7TtpfgY+7TFve3guVIXOAXZnM
h3lf2OQb3BZHR55wdr2CsbsyYDUXRVx7A8J4jfLvfHkxQGw4IHX6cEc8GpuajrlAKzQ57IvTWWgW
FY5RL95ZVvmgz57b4HEYFPb0ax6gmYfzptfFYWNA07MaB7zZIaFIXLfYy3H5W/mzvC46ZobrQGsq
dpRK9+4ZvLexuedXSRvOzew5Eh8VIo0zCnbnE8gH7mSdm2X6ZsJWc1ooCpcTxRTa4/H5YogbHlps
zaH6dvpNR6QJnJC+qglJNBbTAZJ7cSYY54tWlF5NP1xOc97Gm2/P9oR22EqvjtZG9ejCukGWkZ02
mXeFMdbNAbHaFjbCf+3Wj8gnWKRLHu/OSrt7Kfde8/CGcd0uqLe6YTQq6tDSFORdraFB+y3LXsuH
+SQaosUtr46DqZUoAhAEhc0xOQpVJDyd7ZR3+Y35tKrOSn24V8Mpgc6ac0VMOgsfOWK6xQpUpcsj
av6tuIJXoH/UfMcpEZMeNJlijEKd0VdjwXthNj9VEQ1s9Jey/afIOaoTXuFb9nBZfsbJrGNOOGIi
avWyYVeSIqXWUvGie3GbjwyzLNU9KHTEdQRmh3trQYuLXwAmKmSZv4vwF6XWaaQTIZYUN5pbHc9Q
9M5uCm+2Hoxk0RfIpSthB2xqZ/54aw2mY5NrTNvP/2+5/ibJrDITZRz3Dh2CQ/2rSBCJ3HBZnCZQ
/g3mqnxaYcxzGnfxamDgTEkEEOiHtzfJV47YPcJVodWIy6lASd40JSSjvqSgZRpe7Ntdz8ZhfI7F
U4Vb/Ic2YxFMbGlEnr+V9l+3FfoPBYn+lOzBkGr0fr8fnKn0kYY9jaczO9Hb4/SVpTxtgPBZFS/C
XT7GunriW26CjcfmZIbqua7CJH/AFzjY0KvhBGzwi5dE7t914Yrgz7mxjJY4hs7Ngva5jUfF/WkN
yAsUQMxewq/KfHuREyCd9/hSam23mzv6VTPmwwgwFNw73e+dj7M3rFEm3OXb8uVTPipgxsENsDH1
FFeTYmaDQBuu496HyNwj9/NkpecPTLJNP0odmVfcE46n1SHZYmxAKrWG8/zRHsueDxZoeHvUsdWX
2bzNGt4RhVmEM+4RMR+v6GlY12RU6QByUnS7fikAniQFO7JPTFWGxLh3YXGnRyoQ9+iYwJ8APWD0
xX4ChkeJvJ+duxuqlxOfjjmN8uMJ1Ay/NFXBxSfBTXx/RQ0sXrR48L6iNR8Z2rw7MVoNOSTZt5Py
/yWExIHmXR1Y4osuGP8Pdi0gidc08/O73IC3tX5TF9aFcaUuoGS+jo3pLNcnQCzNIo9QE8NsihN9
LeyRnYV4KtxlqjLsNqymzAlV/Os5WPuQSY81zacohRQHAerboqDtjJPFLoYZNFqut3Dr+G0zJpH2
qDYnIiFmHhpRY8D1TltF5cgbt6LoUTTcXSLmNSmdFtoOTHmAnhbMXjmCXbVtZ0qd6oZ3I1k294zV
JPVkB7y8iGay9KDOy1T3zD0zW9qsoTYof+6Gv4G599HaWXjidVTYqZrk0xz0ATpoalg7JTsx4AFe
ZT+QxkU0PtYpiTD9a5D86CnXf0kvN/FqzjpxTX6hJ5YpEJ3bd+s/C1gDWUaIIRgCkPs6wMeNGFPz
ZpJDa59MPOZpy8umEbk3WhqP02usGxYySGByL4cRYw3ycl4ocMkQfV9ViGeR+Is5YNzU6IYQ95Fx
1eya6jWewQ0Fg86Eu96hq3o5FjlHgzO3uEZGElU2C1n2JgTgrkpVyYyNPgqbvhPU9TdluWEurYHR
ZSjefWFozVHMDQ7jSHJFcRGHQNpgCxKNJVhBx/X7f4nj9E2kjciX/WuwOdUzozlm9D5kYPB/es/P
4akl9P3ucFXW2KHtkDhF6554WkVCnr5mPidW+ylpYUJn1T5ZdZQw2EHslVhgxdEDY8m/X7sx9c2v
gZDrHVNHkYYNn07sz6ZsfZGwl5TdNoFrY5pOy8t9aGrS75WQjX/aeqaij8vWw4xwteC9i3uT+QQt
CYquTay0iCvDT6BNr5Z8MkWdVxtRUSc1feI2FY0CqZPtYsTENjLR2CqsTJTu+ALI8x6covg9XY4T
Rj+squMd+DAiOqU6239eYz3WjcrD+Nk0n+p9J9WP4m4yYuu0fmfLpqEe/9liL+SJ4O53BI4lnhnY
kybMHESRWVa4dweuyK5YTvxmI9M2hD9m3ONmdWff4629s0Lk9ZB8n3/2bnmYCXnoG76CgwpGCABT
iJGw1bchMU7ef7n5OWw3ttZWCrBo3xzpF3aBZhPuZlYglVF5beRc4V0y3W7q0kHJ38gNIY4/5JxR
lyFU5EQk8nf1KuHaUkOLxBR9SoSef2rdXHyS4vYETqUtPgAttNtRiDKW+/ZHiF/uCYeKSOSz6yL2
bgnzKmaMfQ3uVkp9cvRAK/EvFLQ0ApFY/hui0LxLsEdMfpM8e0SonAib6AnmOIDvEkK2qwIR3I8C
DnS1vA6mqI/6qBHJ9MbA1bH65DSyXgB6p3vD/qbio+K54ICdroXRScKnM5ccw4hlno/rzg5SmG5E
EJgrH80taRJwhj2EV8rGU5tCbtJvIyZtN1E4IHd9CdcVhOG1S1a49KOpe6C/vEmook7IY6cwHjNQ
ZL5LRblk3zsNb+xYUZ9iym4Q/Rd2WG8FS/1FrAhzz0asR4TkOrdj9pGDE6fHouTUMA8XIazNyboL
U0SlomEX96nLg+zRmC4FZeM5HDmmXBxawlICH7SWzM5Ln/ykNCOo2j4zlLgk+BBBvnJLtnmUyEI9
SghaJwYD5VNuuUWy65FRe9xDunrCSmFClcB6LxUqorKLPbqiyJ5yrgOw5fSv8O/eOyBhCQS2Z6KZ
Mnb3v4kX/QcGUALu/AiHe1y54q1Ko8rkj8Y2CbFmr+jpy69GB/uSzZUekKcUh12HI5ZxDZcGm2is
oFugFutkgUpQ/YgATTKYuu8Maa/j7YgqFWKzgBMQxmP+E6MeRtXJHvkCPQhjHgG8SW0IG175nBIk
Sl5CyqNKTOX+fX+GVA2+5WzDst/uiNG4GhqlYtjYyUY2wmyRr46zYw0dmfra2pZjWNuo18G9Yge8
yi1lgp3AzCrnaQLono2FEK7W8ojx+d7OVAPcGHATTdi2t39naOxY6KcDAMNDlEO14UbuobkzfYMq
QpQ+d70ARL39smzaTRJXvqiVQFC0RMvgUxvTiClBQzHW9SK9UEoeC4ozYJxyZGIqVHCA6A86tX5N
kG+JnYpxrHxDRnsfmbSF4dVgLb7lGw96fSjSW9SYI9JTuie9ouBEeIuX4v08gl9fNKt4KlB3i3BP
/k+C/0unKK5L4JLUIdnYSs6j+52DIfYJzvn2CelPwRQEcHX5r5re7ui1JSHRcUvdyFb5KvGjIMiZ
nvjlYd1s0ceP0LU24AFFG57wVZRuX8CIITi0UsN1rwLETl4BRwZVhdpR8zF4azKZY/9kJjW0wzGQ
5K+rOMGvH29VhkMtrWN9GYsmfPdI9N86NC4D4TXyyc0tkqyJPPtsFgv5T0jFwTADDnetm2qU2+/7
eGun1Q5xn4BflYvfdKETY4KDDnZc/aflRBoVI7z/5qnAnXJyup5RKh8ZT2wHVYMGZXV9Q96grpLD
l3H4PvRP2e64bWeqRTblydUqtABXggGy5lEBO0M4nT4KKtaKHByeUHSU2tVfBg6Z7busqv6J9BVE
7DIb+oN4eACRHi7uDmHjfx2neTfd81uT7KIb7HOqfA3aPbuBfKzbfXnn88GwhYphGtbW8kx0IAa2
uqRZmferwtsUwl355leUXUVzpx2WUsHbIzg/nD6zgePjWAbir4UPUphMrhl94jL9MExrHl8wPkwu
4HayIsjv9r+RqnugHFDt4H5gim+VXOYox57NuiIpMMqZJwSISRv32llQhKeAkzBLvouuRhCNQAta
V8xYxfnu5fCT1huqWwY89g+qQq2Dl1mFEqUul4QYsYDLLG0TpH/tTqBXP7T6oS5WtofWJktV/37s
YRj//2LcmFxDrCTWP5ADD27IX6HY1LWlbpMAYRiXq+kvbI2b6HTmvEZseHYTM60U8+pHjoJ2oLLW
NJ3CdqVxlIWTiWBDWNGkJ/JfCl65cWww8gk2fN+5IwVkdf//WSd6RRdT/oCFF7lANjNJOLIc2MNq
8AbvpQpcFkLl2hf6MYRLgmHWEhPsjxyHTwfkvAxZhsBIxp8sVc1HUQsLlMQUAtkM/GkdAnUNTVji
iA9SaUu2z30uZ7Ex0RpKQc9PXAtmoqc05+fw6YSZOJrHBQEhuYJnmbCGAisEraQKQ4uCfMnwm4nX
y1WZbtgzWrHkipUJgHE6UHqmd74gx/R2T2PwCGALN/06YUEQVjT7lBRWaOkuA9SCx4PAFxOi1kQS
Lr9sORO/+m63UnhoZYakJmqRbB0V1kRDF5DxL6pZXF2Uchi2DN9c2z89lColZWdQFHaxDVn35mUM
z3vWCTw4IORFqJEgyfxH3D8EFZKokE+ZMB1y53tk3Ae7mF5R2AgZGnOF8/hB7mA9CRsWUKfGj8uy
ZuJfYhaH8TLlShzhq8+SMRw1jan2MiaRF9ylS+cGmYhpgffCLmt/uaAk3rWmTUxpSfCv/LnOVx7S
DUYsjsHhC45JiqDYBccyMK0ZsVER4vLVztoLPRFGL+JbwJW0oc3eTldKaGRnJzFjGx7Lg6CUZJ66
pCyrPyPHgDUqDodAxxX5GtD4jNcKfds92qde7Se7Md0Cf72SYFDbT+p7WHRNRmIr9L89VvvZo0Go
6PbxeS8aR+zG2ZldN6eHufBKfl8RHtph/bDQlcCTbD8V5KSyDt49kDtkpyLZQ+/INjimHKCb2yVp
xrexQUwRVQuwWhRQhlhn7+IyUBdzxjq4KS9BxExDxgJaS5UHhXkfSOsojF05Dyw+MO6Ay/zWgnKh
i8OpKoMgWWzeALyDlkA17HKi1pPHr5ygXez/+Fsz8ZC+S9bJUMwOLOGu4E77W8Nt+RPj8aYXq7oJ
GlCqZuvsjH0lFhYHe6RbjfPu6FWt73dbPiwB6TLgKujRlBwIwVkWjJfk+sDq/R/tFXIdIc/r/XXx
/gW/Pt8ma0ffOXDuGd9JnI3VmgcBFlfF8/rL6gh852nHhw11h1rZ2ZwFI97ZoYGG9gzDtKmHh3yj
l4iEiPadwyP5sbSC5Y2BRqxIkYP8E2zdA+SNR1T978xYfmXh8PjnoCI23ut+e9KDUaRZ8vTg+6OT
2lbB0qI3CjQtH4yztM326VIZgGaTKZ2YR8cE2tomsZ7Kvseu+KVcupKd9lDXiwA77hhBOYbU0V/z
GulMQG0fCu1Lz/Wd1G399biq0cijjOx7DITjHd0rDp8mH2r0gAVf0mmFAqb30kK/g3gS/6Uue2/e
s38Qs0JDiKZ/MTy84HHZ05HnccHW1UJQbQdl8MIBv4uVmod3j6DxQk3m6t+w8mhjjwhCd4uewnCA
sv4jeOC+rgutQE9de2/yXwqCoQzN1m92HffpjwRK9rXUAyufJl/uCGQylry5W1i8maOTkL1AMbpH
8Gzz2OAnJ6MKc9p2jihYVSwVz7IObgPYNXf4hmpywbI1T5BNuhMpQzmRaeA1KFj2YOf9fdIvRbPz
7gmERBeskYnFkO6N8wZ6Jt+B0dxCQ6KXIkwbSq+Kwx7o5AehKmqlU77tLRfDywUxqtzeZShAFOyJ
wA63FlwW1ycXfy4LKyZ+U78UelqQ/W1awx/BBrsZP1YmTR8fcCXuq2TjB2ob5cE93CSHH4a4D6cB
RR5eBCr9ubMUprzunQpihw75d1bUFsuCrsSQEkWKLPdricYPeLEJ6gYJeSVV33uuRZCrc4Rd6XiS
Xv7SRguLwU3haFZNdze+oXKmuPYnng8yHRHHrUuvztNhKpaVIWVtJ0pi8NxarFiw7EudWd5QAN4F
hvV9aNPGoSaHdg5kAlXKZVAcnFOkx6ZHpLq4SnV+rVVVZTWsauRDGQuqWMM97+JvvV59PEkkKvng
c54xN3EQOQ9yT4POF6pJgeZBVSHoP4pAhx8YqALKjTnNH4Ypkhzs6cZrSwLJP8gwZc2Mqg1eH2c6
fIXefXuQr9V7yY32bvnuPfvJLh1k5FrX3IaDWujggG5d3DUbIWPM5k6v6kIhUJ6YgYODF2h/bCog
CUN5rS12NoO4PHshBblqraGKnYTuyZwMxpeqN1E8gLtc0jfO2WpvcZCCI33TDyn+qcnw5MZrkTn6
GipBrY0KWUp35ymQpojgMIP1GIrSigb+cyuY1tkENF5T/ti5xCCA3hPsV6EdVF2am9yR/omKmqjn
wsuGRj+7DABToVRQmCOeBmbzDRB/IVWO+LWJNBZjqB9ogiTbfuVrf2TKbkG0ckc9ynNR/+wdxg44
9IxFF0AgBehXQy/JpY2u99zyG/UebapPLthS1N8yiX8U/p9Yy0xz51Jk49Eo9g988wHoHUJELQ+4
UNdR5lfxJljoTKLTsdtm8fYpl371iYAH2I8nxDNb8uMgXZ5Ur+CQxsDn2IyVMQoMul6YNvjOc4e5
Lt7WcAY3LCQX8Py7O1VWDY439ygdxp6ebHCoInDm53qxB1r+mgfDdJPwoA84RhezGwQoVrvMGfDO
VZwkUvYkh0yPd2/NAEwBN2hIfF981L1qYbh/XfzxmEazNnS7isIGvJaS7bYaoqXQf8FAfRpzt6o2
10o8YWggriOIgUrxOcirKwWsqJi6fOYFTj8sAk+CwPcvGv+brWMIDZnJeBVpGUIAo1uIKrNC7EVQ
SPalKljPiI/eVOJkGb0/XbLlZGiMErjqnwSFrTol+IVRRzLUkE9m6FMtRZY9/vjIDDRY1Axd05kQ
15hLiVUzuhhDt+eluIGt16+/K0BOiPmxHG6BEoA1RpEDO+AS93HnxEbOnLuyB0vZe5GoKvZCnl94
+T5+1uN+cxHocPRTUg5I6cmDx0l4TsoiUdM8eUzjmd58kjwvC9W7q8oVDMe1lvFZzaKmX6houMYK
6JAIj3F9ofXGdtM89R7+c6ikowOpYkLk0deGXk9RMURC2PO0Y9PqqX31h9dhJdvBrjyXPaUw3QCg
EzONwNVJ591sGhdKy+W5k+0UX9mgzELdQmkJhQ9IEcLzUKbLiI0OoJyHY9EUGrNAI9aneGjXjjqI
RFQzeRKTsRNn77LI5pdp/ZDIr0iWSVZNsbKXRGuJc0YCjP0/Zq8Tn697vyQbdQVRThLzcBVaIste
HBNuE55Aqx01zIybEGjHJBbexwu4hH0mzkvmgwyxl3UJ/WRz/pHSKX+A2FKbg65LGM5nuQM0BO8A
6Gyx0CZQOEU5j124zpPnRhkiYVpUrjCovDjMOq9WMFj6gOjODsjIThf2H17ZlLNSX6cAK8qC1OaO
03sI/A/RGY85dub3k9K08TLt95zVLIUJPher8r2oI6V6wszzsEA5rrlvzK6Wrm7+5u7CByJbCyPv
lTKbEzE1ECOYyrrF2YhL65brYhRuPllq38HSY6AecnuLfqE5h/UyozD6kqNQiFMLpLS7ojqgUULs
W/m73FCNnGfEeKSxLNgQot26PKvZ5S1MrULdzgRKcbk6SXnPzNZDoqiIH0hJ8FZfahop+9FO6LqY
igsSTTxDOckDVOhT0KuUUK/FpXJ3zmvYCo05V8ZuGDqFrTL8mbuvA9nYHnfebC9v6GZDvini0kNa
ESEZ6ta85flZGYDfCeWGboSbbu6HUz84c5G4DRBBboyY383O5h1/rpZcQ4ZW0GTnZ7smMmVMiajW
m8I/O4jKZp9sDMQNgQJs3lbY9QlfMhUIdaRhSJJGfRywQrJ6AQz16mpZooaWCk7fQqZsHex1CHn7
pnUYXkv8vaZ/BJKuv6cf3d43X3iZbDjQf18XII/G2wNZ++7QD6Y4CQiEjAfVc8Y2/vyQCvvZCBi8
AMNcY5ghz8qyoRFHHf8SW1i4Gy6//mh5Lj3XHvAxXKS4ATr+mT76x6BHG7iuX/5ulj3jdiiqk0AF
MVih/4lzMDxxkondYQFaYYZiso92EXV6wRgEfSfY5ALCGwPxMb/ZgevPtHrj14yt9bxxP7ez3QgZ
tDOvRc3W1nbJXeks2tfDzn46GTFsA6tJOpOfsyoQh9djqXPOsNVWlfd5C7YAYsHImeAknYy1Zf5m
HEkVdwzid5FMqJBnYL0TN7PTser8uJNaOP5Db0fY6cRUdoy5hbWdYLlOgfD4ZXIZflSjz/GmWhKT
2OvqQhwAUthVsryVkuN4d8ykFZ5siS0/Mo/+74rrqlSghV7zqbqqvsXVf4W7ayOYZPAXVi13JbOY
jXrQtcSz21yexRiy92tTILq0jUKrqwFxRlsTGEGiXgxDpJ3whC5iJIZB7Jvxf8EJxn7pMzJ6BUmY
PAUINuVLhUDZda7ZSazuLj+y9VuJ1qoILavoJ5A7i/XcwNA5q1kDZro7u6BDgo/wDy0Y5aFBClCB
rQbPT1xjd4jty3t3e/+YDRlbbUxLcekboewiWKa9NzwltpxRGq5yjjlbiLpWzqKHCAlT6yW1atxu
C8MuIiY6+Wb7t0BiVylT9HDzqjFh6LI6543lzsLZhl+3rS//Gpn5VT1ldUFF5Twm1clCM83Zodbk
VkwTSsrXWYeLJsP+JcAghtoWoyX8usLjwwTZjcCKWXLlu3Kiy1UoyHjvLWmnWvdm/kd7+r47LwK8
rf6COc3EqeD1f87PpUZW+Xg6dXpfVQeQG/6jUvrNVOPh0zlB5F594wGkP4fIyB3dheYJ8UafMqjH
jYM3kAQ4Aa4p8kuFaCHLU4ez+DCbIbB8j2Xyv/E2yMmV4C1K7Or3yeYptELtNaeauBUmU98bH/3o
s0QjWbr2Shtoq0a5kT2ImodijcTZ5rhMYTM9v2uEmgow7/82FaQXhpE0+EL2PXwNaCtiS6JHUUBc
wJqyjN9t+Bip3U80m54vL9A0aY47Gws/1c0dVYzyZPjqbLvaWFnOBoda5pruIzt64OGIx955xQij
iUnQbGk5F/1fQdwV9wI8t5nQJg26tjlxmbDTgsvefl/HyFZyjxFumRirqtgz1vapvLe95TPUYFFl
2M9zkMu2FziUfuhojBnCUS2qeHpLV0mwczXAGoM04JYt1TXXRy5awytnrX/omL6xeLX3NdDSSnm8
8cOwTrToC29i4GjTp9+nqb3Ib/pTPTo7ypL/MTvXU35pAUidze4dUkSiqSLvyInDb52TbNDz4S0c
o7V6fH2IPX4UqQku8fKYCEbegukdCb9eRux+YmgzvIUwWwhLR96JKcEZufaqok70jvnlp7Gqsq9l
dvuMu6YVUVPhRHlDIWiA2K3jgCCPlBHYj1Tk4pWbBFB+6Z7aHC1YVQ+UWgvoO9Zc6Dx5tseeAcAv
krfLzc+jsfvsJDA/3hgm2kRX4yrqEwS9+l80//JDh3mOd7lXH3+ajoiYR+5h7mBN6heV1/ybADUB
uOKOk6o6qhz7qYPsA9mp81NXorjBTZ9SOyghedG3IsczgoOyLvVo7q++stTwaWHuh94RgN3fIU6/
yPzx32OEgQsRIN+F2PUqQgm9y5TTkhIDg0mFqUXvAvPxqgLaZFGEHUpimVHw0M8Lano5lBXgfWyP
abLmBrAjj2Zja7DIj7enMux54rblDydtBAMGBNJlpzl+UXSaunUwFtlog6cjm5UqcY+Wbu8zU3Mt
+QDel2shGoRfhOz0nw+7tkxf0Th1q68Dmdid2Bv9TunJAyK85yL6hfcAXms6sh2uUz29j0U43pqB
ZEQeg/8cD/cbA7vdNbrHAvfo+sdFPiRRktqoAkrq+Y2IxBq8UoQVbuqupA3rpc6UJhDkkPx9dmqT
pXR50aWgjzP/lsEANVfwdwR3JK/osfiHlVL1ID44TIKlLXMdM5E4LYxVYMI5kPy8PT0N+h9jlOJG
8tIWBmGzETIdIPn1cKyhFIENZ/X+KbAPBXIAXr1rqL3HIErWLvL/hOWL4IBJrtSZ1AMWceBuflGC
6Pr47Nme/8nvsnffdXz6NDkhu8bQzUQSNE7y97pbqUW2IiJfG3+iLtAuiWkV5shdNhqHmXHtpwLJ
z2+xA28fvO9kawOwQdMmLMRCme6tfPiCF59Nk2gta09foHflkrT6y56/MzgFNYzuAPANqLwPu6vs
/vneIbDr20xPCrtBczLJR+DfICsp5fTx+VvEjX0zbh5eIQUG7QSFMjVyEUb+n4gNh/zm0rn4MuyY
am1AsYuDfZ6R3EmSmJsNwOQe9BlqoOInRL2cpP48iiO9pJLhKy1h4JUA6qhert65x40fHNCmQGvx
+eN2vN/5ncYkOcQ6Xrq6UCxKo0O74b8G5WlMDDBOn+wA0cbufNqlAuKJQUvmOM8s43b/bW5kzef2
vI+sGywKg5afjVqimXQN/jEwVww1bsgYy5GMFtdNUOIAA6/7SmQl16qTqss/xLAfRK+ByrS97gvz
tMq3qWKZxqSvdsALHG0PcWlokjEeqEo638YEqcHzYT73RmbEVWKPvnU7+OefW8H/GR1LQ1enZtoJ
maTJcti+IzYkNGj/vnzDtdXdv7IrADJ2WIgOvSEqWHZ54yuFG4/E4tclmbd7kowkXE6ICyp7l9on
Dg/QqdDGTcgHlgG/9sFrU92ouRdUJgYpyUzfNjT7ddZhd7TdJhZTyNGUQWG600ah/7Qud0a3TM33
U/yAsKutC0fMMSwvMwbSyrEOVq4KaWP8sqlNlLyb1arjcuGaTORLycPdVg4UnqQBrl1eCKPyIntl
qCBbjFi1+/zZN34vuAFX7wjshEXWZwWX7LerQlcys1ICzBin9HIkcC7XD6UgrpHQXG7B+wp8x/sf
yDIvr2kRCh7FozqdQphruG/Ax6bwTtzWxMvbm69D92GgHmoiHT6qxPaN6Q0cTTpkywpzXUeuyANO
cHAdX0lY0TDsNp6tgp6c4IORjJYVQ3L/ITFei19begqJzEFVneDjQMkId1cCB9LGCpTbjwSQg6vM
n8gUDt/MN4C78qydAnAoAEpkKuM2MbXRb6MdZo824s4Ww+mx+4nvzSAsb+ufaN4ZStwYr0d8I755
jPeydWLSbtWU6YFfW2UXpo4fvPAyOxwUE6382Jq90s0GnEiiXcEbXFmXKvN/PlbfIdsuOHOeI4uX
/BLOixfLAwJhlNPPtm1rJmXHtV5eygWqI6tmyYoQIRn4jQ97YX6tIo5j2grNIw4zy1tUVloj4RdC
nvUXwYG3U27u6Uyr0+zY0kY0MRbMZssERoD3Ys9Eo300g3XTlyd+e3j8mkp0/P1Jnk5cUYfvqaat
fJMCEehALqnsgOi/54Dvr7FBTaBmNaNfdYAqjOQY/jkznM/o82Y5x/ivD0VZDt1EZmJqmDJAeCTC
q6WHJ+cfir+LUC8SptA1dZn8izC3lsiWi4GEUp/+IPve46dlKt33l67zsM0szGx32MRwKiwpnCp+
tb8EoFjzdC6c25IVdaQ6L6oulgdEh2XXUCKpnE0dYTH3BAQm+/xJI29f6+ovRi3y5DxVazSJugS8
YxEyzkE6cUfk3Z0F/W4SMvUc+2J+IQy5kpr4cNoVYvSUgF4sqqhJ1bgxlsqHnsGIp11rS1iIUQVb
cd16QUJZMFwhw5XQAawP/yH3yd+fifF5inhW1RbOAZR65C2sm20Rz2tBMWeGOmL4pF5UTA1NXW0O
AYWskAFMTw3AcgRXljrNZCTP36ckO6dnayYhpD7MELRnBE1IqWmlXLXyedEUH2AbZcMFsutAV/GM
i7oQxyG++pPqflLGHK+A17m9IKImqVwACz5iD+N/HMe6qOE78x/ZBsUkJfJMKxStdptsN5UmFLWW
yFSksf0XTf/MBZlHZjONMF0M4eQr2YV49RfjJvxNQKh3Pr7OcsNEKeN7FV+w8aUNKButKsCAC2Jx
UPNF5g5CwL/mqHfn9okOgNmK5dahCtenbFxzgXVfBonvHygfKU03yoVD4ToqQELzGvmAGbElmZSA
TYY2KcJMQq2Pb+fVZN/NPHzze+5pv50STsAebJz8EMw0Vn/fZTbktL9B1FikK4jHzEmaCpJUB9nz
8DHVwbBFBSCizDZXVx5XUVVUKECArj6TtRwYyeJHjjNVXNkxkz5v7q0ZYfZ2/J3cm2m5Sc0RQggZ
JyyuVvgAM1kdEOW8zkGSHHEmq51eMQv/gDgDfd29MFpYhlugGhZKpxFeRKxQSuXdJMbxTkUueenZ
yMGkBJDRoGMyDkBwzNpqme0nviAITxvH3jehsYXCBHQoQR1udwALrDmyde1YQvtUwun8GAOogeoy
nC4wQhZYBxx1GndRyIyC9fKt0AYg+pczggqJG/aG0rSsNg+zGeu+6aE3f9zj6l7g6dHZ4/dn8AEr
MMQT52BNU9ET4EPnk0INYdl6+bwi08hWQmRdSzvQ2Bh/CzgWV9uxI/X+UbhKPzDyKVV77ReVmGRe
LNJzBlLj64XvcYPfw0iQzPToatbSURNGDOJXWoySIl0PTfLZO++wrZrVvLLHHeyKxcDHL4/jK3Rw
4XnmgTJxeWLUfst/FG31YGn9Xapr1fhjf8Zr02CSSCA0vbtv2REtKYeDbR5Sp5/yasWKB1Ui4yCk
j5sop8vti/BZMbdkbr/8VfgxK2z59bKcwnx3dGdKQrqjhmJWJZkzEQZi9XCfjMRSdWU/jqEdTH0N
v3Iblv/PY8p7rlKlXH+KFE1HXVTpOr1la/EYM4UWariS3zzwuQilWbI9rjfmi4mNCJVA7g+HfiGp
OjFKG9oLeTiFKLwfvw2BVN53UsKOwRGdvoMRkU4Es70gSBaz0juZHgDwzPsXHF0tsmq4kAfPiyMJ
hqdNQjv8ZYRTdj3KRhr1cTTcF+CSluO0c5C85obDo0MzN2+IUxvUzEBrjO/Wy+ozR+Tj1sUlslFR
9xCvHbkgwjnT5c211eTgv3iaXZpa59kRlDIbGmmTDk1IYByi5NJbyWcwTMffza4AjibyNDRFpiDp
lUVoAgx3OQaZY+Kan3wofGm340A1He2ZS1b4j/nfGG1CbCNaHHruRIKaURe2ZI4XmM7EdbD/Rl8c
JilmcQAF6nGvAANyFkIlcn1s03GNJ12AFBJlWUID1eiZeAArcErjLOejavatkdMszXvhD+IvVr+u
QlcBAAI0acbLTol0n7xQWSOSQcYHs4xzBxLN5lkHCKmn7VlyOIFnR3C6Mm8csoAD0VExKb2gcUjq
mOgIQrYNs8hov8lThMbh3/POuveykE8iOKMHVJ6YINywmxA3fpifkmhUerpLa/N2VcNgKz0+H2s/
BvXme1st9701jbXO8DUV3wiD4zUa+3L7Zdz4X3mRXHu7FyTD63BzXi8dsgH5M9ZwLW8Tm/DoGsih
EeIjGON8bTUtPbWOge3u0YSBjATPP2AmyXtVn+CQ86mNQMdnOPbzBiAWnyYbASQ4wzhmY7f/HWQA
94ITFHraBWfOlST0DuicjnFAZ+KuNbUgH9EnlXObA/YwDbFBxq/E5r14PUugmJ1QE2XvQOdEFILq
+1gOYeMLwFUTmdhwFjPYMjG1ugfcQTt23sbt4tn15GM/KaRW31Qy8nRka9BOWCEwqXbmkoS6ea0c
6/bw60Sx8cr6OTwnp9+NMsHkiRrP4M0UXXGrkFSerPE1d4trMmbsPYXQ/vBOZTWkFQLwiZ7M7Lho
oe8Uhg4USwdshK2PlQ9s7wfLmqIrpXVcRL5DISHc09dUA0huCzYHlGM9T1S6q/o3URQ6K2r29cAk
Dez3kMpqmoT5TiFMSWMf8D7la+BtNbROhsEp19jBIdfHmvM4tfNWmXsWEYi2Su1R1r2YzrYildk4
Tp7UZJo5DNyoTn5jNXQXy3NpZTbwg2rJLOHiPMvpEFJrQAjYQMOVK4OTBDB5ctcCeYxvFXqdB0x+
lxPkM7H0Jf/24wu9MKeEl4g5hn/AEVpwiX6r7L6VWiLXig9Ah3D0oGMznD0zE7UdBmwY0d8UGJxT
9rkg8YKofLB8gUZICKwzm0XXiKuSKNXz0G1jJC/AZkvwAN+56tEWEwI2lS3TM55rZ/lcV/A0S/Vx
L8KoOa5z6CokvrfEeUnIzGo0YqwV9xKFLSwvIKXeD6uXzRw2GiuXaZQARkjo/f1VLZYqcdjSNcnX
XZ4O4gYv6JVtpdAoKAuagmUlZ49rmA1c7G8DRFFvcunOs+adw/afVFVNB1Dh9gZXI2YcZza5rW8k
sUQvR/AhrYc/5oY5rKO82KegKXA5O98pDOklzvC+96A3uEgns0KSvEMsmzsq79yB2LHZpdrCsvnH
RoTT2CR2ICmGNHelJF9iENP/neD83AK7YRGqYLswzxzTcfakYaIWvfBz8m0C89axDJO12+TVXTJk
aM7roh8V01R9c1HWMjFx3nuo/vjpq5hEOlNdz5mdlGE81MXTKhW86JZAiH7rUWNpOQ/xo2I37E1/
q0JpUWfcBnvYHg5y1S8qhBnbRmyNy9kej46R6Xux52DS1bvDzvaRtJJT6+S9ZToFZdNbnN9mn3Xz
2L3hAofhNiO+Q3HeBbhDx40EjELjxrY6ylByeyi0C/4AtnqsTOkhM2lH7YfrWTxwa/q2hB4L4dYy
9OB1KfPzxZxoE8w23l4gwG4bg7v0kKSSoEp6FeTa431kSqiQ0xsbMzP0DSQ4lxPRdQcDXwLKNeYq
KvF2gpEJIorgw66MqpISit17d0k65dddwela9tpxc9bOUt0mqTS+EUfiDFQ4RmJuXbsMh9MRHT7w
tgg3fKcc0SdOOpAaK05rPWKOoESI7/tmxJtdHpe9N0oluQ1o9XzZGXZhxStEAcdQYoV5CNEOA8iU
4nGyzMFfafu8Clxo6dOhuvJcJ8zm22WV71r9Ng1nQO5Ab0whXRn0JQEdq3gJlmfX4mMUu30rrXx4
SgOXVG62Xyd9YebOtz+WD/+LuAfo0r6aXOoxsCdoT94l+SsVJlxcISpEqrE6kbGD/W+Arb2ghnzT
QETz3cM5PusBX94DFq8KwJa6C4o9OXUUnHc/vLtHI84de29KTMcvP3+zuPBgaqjpg1DVbpT3tZTy
Hx2GF2wIWsJs5xVE6EFFt1xGsCbNCNQbcxUVo48+7qs7n0rSsXwey0fY2hN2cvgsF276WSjVxbv3
lbzopD8gSilgZbg6gBc4RDY9HInU41Q6nM2HG+6usCV7M55AFmKM6DnI3jr6FtsaMiW+g4lcD4PI
XbvyrEWwOvM2BGr6kCfewBlo1PjXUo6raetAwF2hmHNE0RMdwxSTpeb2bW8ttzTzQsJtjwTnTFAb
zEDtfo0qkkBYVoDHZolpACDniB2HLIUWTkcz0Rv6kct1msPubps7uglMxrTg5025D73kH2nB6rSU
CDD7iBkutMS4QyirFs83DgznztWs37cC3nQSeSqlqsyo+YjnxQGcO8IlkjavHz/mR3X7uoF3hUlg
QAVDOsRgUKAjsFhklgIEzHl2x0VnvswJht5JIvpUrKA7Yveikp7LvC5y0GZIHPZPZ04yBYWPRef8
htqBYGDgcmaqefJ9MCpqgh+9vnXio88eandUupzYHhrtMvDF7cd1dNHOFnoOLZMcXqQlCSTqwvep
PM4uO1qDRYayqTp58Hwa1G+c3AD64bt9qFgF/9WYc1fHt9k0LoEpf4KCPw8RHdH70RerpuYGwVI4
vvydOJfSyL1tCCSgy1Ipd3wqz4BnpER23HAOvxrtFdpNghMHeXU75bus3AAtxAp+Vza4R7irh6Kc
RrimUEbSIm0ZHGHc0c6lRIzMaQeKzKYtWjwII32aDxoa3ozIonfmRI0TV44WPzinm38ZDnxX4D7H
eNOmTTZNTUn1oalfLrJcnMGi118WX7S2YVL66UvKxW+kXwFmjiOya36f606X9pkd6oVv0uzpJYLb
zZ6Ra/JEWHxVqGVFi37vLUnhoUif45RbMbM23zX5cCFJbjn5YoIng8PaJkfvzon/ObY3vzOsjOKK
dZ8Rm29qzVxdwPUqievyyoaMljkImt0Q3aMCtTfwl9AwlC6StqgWtq1qP+BvzJwrW5xf4xjuZdD5
q7Yul8+f3Iu5VhbUzn3jSIBLQ2dGHsilKG3qrhMqO5JFpc7mJgRQwHGPkiK9Lb7d8LeVF6pAtXtH
oIS2JtK5RtV0n9EINnlsUMAdOa7YA8zxttck0+frXqmm5sXCuxBSH7sJ9xXABlnTIe+r9KJo4prH
BDNGyrKkA0eTfkLvyEO/YDtJ+Qd764Zwik3XSMBecM+oS/a4EFY5gJaL+2qRgiaG4CIbFLLNtXVu
T92Gf6O3tLdXFsXghfZUC39dMY+CsYMtD5EO4F31LCEPnV0V1GUyRhx/EUmcs5krC5lZgAePC+Ap
Z/PCcSn+aLLIWlayS47B6t8x5Xmh745k6Xj25LNgn029VVfDpN62Oot3w2nW0aq9j6QV6Go43KrZ
AO5qf8VfZPJIYYNNBy4/wbPDvKKpeBFnHavU+8ZN7U1uzraSYD4YDGbUheM5/AZnxXofJlGkn90k
CIkY1ndSpiZMbx11gu418MK63UlWMLKQwDwaSDqVFAGWJxefz7zCCg4b5erbnDnaFAEIdx+/H76Q
Qz2U3Mnazr3uGzu9mgOuuCEv8UbM+Dig7KMx6JP4ILbB6M86t8I9xZldYRTHxajrM06njIjxYVA8
qquegk6XbKMflupZ2ybCZOqv6fo603gu9gMiudNb9MSsn3eLUEUM+bugIG4dGL5uxhHcKlh63VG1
ZVusycZrwybhdWdfiAZIhs8iSv6Y7TJVxzVlC718Ve5LFwfrU5in2C+7be16chpyTYq0hkza0kHX
3jP4cTgHOGq76woszGFTBaMiUByZdYOd9LV2iM65IAj/3cGgJW17o8sOySLLRYrAYiNVuYA1wd/e
HZZK4SXNmYJN39U4kCWHFuFBC3pIm4ZrGhkzbgjp33KNfSUjO5KIgEOLAcStcokgG77f0J5DcT16
/ORiOKstI80nt3ketgOXh79/mcWvPAp6tnj5RhUdrSj36lisdtigONsjStF++aTJJ/PKp/ApG8dD
woDh0HXWUC5JVtJYUv5V9GA6IKg43qdD1gJ27p8JAnzf7HY8mvvRQHXg014m+ZrAkeCmDDuWNXF5
rCWI7PLpIeWJBuiEbtUVXoh5W5/wpv6QGvkbwg+K9OLMmPNeHfgq6+I4zKLqvEJD3cgAL5NdTPZd
ee+Rvk1Alt6a6tmxp9f4mGU+x4r+0cdeGPv6wrCp3r40zMRj+L3AKmxo42O/W9Ffx+Yrf9EwSFkT
W7s9/rREcYri2vavFNh8nn2o/JZSnXNXFLYwDHKbL2q5SaVZW4tSrKkrQSsJW+usIzAMF3P9/KaJ
Ge44PS5LzIew5byDBZvqZPGVoPU+yzK7DPyOeMEt1p3sxkNwEewSTEclmvGIx+OmJwZvlldcuYT+
NaA/HOY6p/Ap5U2wwv2VP39tTH2jRBR/aO7VKrifnnYwCnA6ULbfsMCBRg9Gx/QSdXIxQoGqzVpp
N6s9S10jhera4S9Ms6Cc4I09dTK6K3QLh0HjNfidpEumkrgjHJg/aIVsOm6WYoj+Vcv/uK2zVXzT
BwqLk22xRPUmPDiRKpKj757sD57OBPIYrkyu/pBQFIFS1h+dJYiAVpEd11Q4n9rmBBdD9/ApQg5n
j2DY9J3ylTxGSLAynoavRPKAArYyyh7MozsWE6YMRs8aM83WDbin28wGct+JobI2GjXff35LFYjK
uxuTGne6mEAPg3IwAGsBIKW+E1OfXTkv5r+o+JbqOhxg4w+voqx6jfFiUo/QG2t2vqIlGI3+VqaS
HwqcLg1QRqGy+MWmTiJYhNujOn1H1G1rlFIcPAkPY6nnj1VpOGqAe1kiCO4q+VOU4qWVPUAOKWy+
GVlmuN6bhCeSLXemyNoJhGzR5PjRvCzoU/Zigg1iT/l9D8BQ+r/0WN5eCIU+rR1l94Errbat3J4/
aQo3/jqc36ATcDUdNJFXkvDIGWhtSxmOX+vvcKvUHi25Wo8nLB33dkkDuNdCL9zaDQZFQmhoFHBr
xPXV9C/3vlJG4hh79RT1V/mnR+jWgSUcZSVKw35rxhDn2Tv8+4oPPuOgSEB0r8UhRXUeJFv+1tYV
oGYYbc5hdB3EveFabLcWi9qSFiW4CdUWIp5vcWP/2tb++BHMitE0AaFPong=
`protect end_protected

