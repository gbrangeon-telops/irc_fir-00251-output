

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IVTcVKz+qqR6KelbIxn6hKss0fyLwIejVgwej+TN1ST/vU6syUW6hxZyGugx/VRu65UT+0QU+88C
5SDN434/fA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W0uuDuJZlgdtFvYMz+doOP0vwnGc2SXfLiGH2a5FulZQF1GjNx3fjKnarWbbCm92Rksm2FFSGof4
SgtGKAeCq4Yz/Vqm5xuP6QHmdBwou49vkKDs52HUud9c3EaEYtdNlkb4+DCcueqZu76yWN8rf2DJ
ekmu+LGiL1dmyzv30tE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Da9hmR0COgf/nsNRjZU5mrjIzRjN0/ufJQ7crbPh82WrNgInUm192216ks1D/Quh1gQ5TieAOChY
26CHNdLfPPmjLAo5/cOIRsIuy2JD7JAEIDFhFO2BcC4GrUAhSArSC4/9FyqXrVJUKuDybwv0tWSf
qpHjmJw18CiVw84ne90mESBOJ0fW1ujayfbI70yaGaFjJM/DPm4Lq+TC+TFlaimxpTFNrAUzQNVF
VSkf44Zb11D7if2jaL6ua4hPGgYpPcisaJtcEYpURXS8Lw+NjmMExnMpUW39NqnMiTEPom3YBwag
JMKm6/EZOnBvVc8SljH7y69fXiGUXgw6Z6POkg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1/llP5a+sEX6Ky1I5ak8Fr3e35uMro1bXNqkrntPBRVTqUhQPFl7wfr/6Abnu74l73YggylsZJi1
1Erm6sC9oDhL9IE4pENErrDQRZHuFnl4+DlguLd11swTlNfBwauGoCBXbTtZ8+O70UI/sRzXqbZc
NDH1RywyQLhMRmSOjCU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OI4vyCtRzSCtjYNsCqL7rYkcvPw30aumOHoxNPQx0NU0Kc5/zvGo5pjE7sDqPsv0b00mAjKXUE8e
pVllo+uquegdt9Smrq3DaiQC/9hKGiZzOG1rJH9JbLcfPMXDGpwm1inP51BNgkQwocfUEAVndeWo
GE1Y28I9gt/5q5Fs/OUAX9cAh1VoS1OcnYX2wbgJSlzuLqnGWRIxOHl4+NkNkBq5Q3Xm589bPnnz
m+d2tBEPyqaCTvb13xXW7hqIf0ahuv0AQTuiClY+KmF0GjLdJTWJjDWPuRd9WYhybCp/lrgDnhAK
cnRXJnAOwP1Vgr7EPuoyVc3UkNsZTxEr3wrouw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11680)
`protect data_block
zIzwJGwpxU0+bFjoj+zv+bFCWQAMgsmzf87Jur1coCYOw4IbRuTiX//cttX03jhuMUyl8fa34ixW
lOEYiQzqa4XEAS+k2PkGW1R1Cy4s06NxaJ7ZsaTXjaKDDEuIE83xDnIIAckI+TS9F6Rul+Ox4gR5
rZ5f41m1CL36Tl8Hd1YKqNaix8TkwWOVRf6FAjZaLomelFRRGgm5IivxCFhPZuRqxmN6yUVHNHrX
h7nG4dO2oBvjpNCn+4LdYUkHXkkgabs2G/kTIh96yUOqiJPaU0L0lQP9EEThvfT1IUalAe6/FPpF
TY0AwO/R3NwFC+oT6bsdY2XtamrfFYxqDb9HsauYk8AGHihsWY5GnHCL+i49PlIK6sVsmzLJSzkZ
yLFAB+2I8cUuRvWR3F9ETgyEe/w2I8VPnGOvLftcaFcx4uBXhMzCV0Zdt9Q5iW+To9uGvugIO4AD
n4PPxpt/DVvGvSBDk7UqIGnC00cZ7s6u1ataBb4VF64qyX/bPhypRneH6qA/CGlfeBSimMpRIPvW
OIosIroDcdaztRaGUBcg+qCfFuShjA2/FHcuARqYM1mgHh4BSkNUxmfEWazxO1IkLtPkOi+lU68F
vr4SIjk9G7P0PRE4U36oEi/nhqUJVLBXcgtBr9NY0TmpYtEwZ4amQWV6nZfLuNVSOPCn/K5WyYJx
oeTto9iu7nztX+07ftsjarkv+mGceIR6muQ8ELewFoPS2v2SVbuB9TB78eNY4qcrEP8wk36FfIDU
pmsKUgw+sIjsJPENdFvIxclwNCp94pS1HnMQdjCelUrqrabwhtJcue1YW3gYaCFgDkxEX8Kewzq3
/j99+i679A5xP97BboK+90clA+cjCqNAr/VhY8egAsr1bcZvZ1ixgTX5SOtGdiHuUl0WbXXOVswa
NXolQPMMinmtM1gUVtZFLv3uQkE9eVQ4acbMSvGsJbFepgcr+Mi1AS4mwEvokFiYH2OnlPsSF3MV
piDcN0LECyPDFNLoJCiUBE8Ik8bBJ0OYTQ4wy5nE615IqNmDnlOKBSTFze2TfvYXBUt9jeJk06BH
Yx8g9HpM1fvaFwRzINDKsgqrjrO9vJIONWtoEZpEWH3GWTex0MU1/5XNx3aJxjOrmPBNngg0Mb6/
PSBIdqCZRlglSyoi3vTuULBBGlnVY/f2eB4v2VryclzYn2yEQUtb2eg6RSZ3AJWkzNRwqibdKJwy
YffaBhxUVENT/83JKemYsSUbMj2kQ5JampnQUyh4vTmUMQvRYbR0MO3xyQTAm5a21Zq+nvw/9RoF
RzsjjrizlNVoZ0gcZgCq7Mbc8FyuLjexZu2JEmiaFv3+ArYA5NNzZNCy6zb8fTqk8RSzjm8IQq06
+2xW7Bq1WVVDmYEXOAISOsbHt5nbBkQUk22jkMNM3l7und/T3+ERasyOZaXhClSW5tOxJF9Ojf9v
zqsKTqcEzdSdhKcDXra/Bi2x9vTpGDB1mYf2wfmrWs4YZZoh0UQTc65PmGwPzHd14RJGkfsKUcmA
HcYszLuHBzTesvW/6REaSUoW5Kn7NB096aipS5cOoGXpXpC4pBgEiI3dVLIkUZWtBol7/4uDubir
qblRo31aSQoh3x13uxRW1kfcsHuJLNgFfAX1ICipGi9r1MH11TVVvYPzdr/0u0ctf7ZjwHWODPpn
2pAUJEYOsgEovHKVp9vtnMkNjNukD/XzQPLe+qBwBTDQyV2Ze/TxjgqG701+pthYStaTirYlAcg1
qH6o34DG95X4rSLPJwxcr/e8k6ut0Y0gjr/m3qS1rZ4qdcB2nIQvXuArt6M6owEriAl9MKL5/VtM
v0mK57HuY3AbCJmscn9/+qEYzNGFiHBgPcd7bXYY1nB5/weTUIruIY7U8JUL+bgynVHWzL9ZyWc8
x6a4aQIWV8mqsps0JbpGxl8gy0UC5cN2UKi2IldK7XYvE7tdgXOfWFc8+Rmdvr69cZqVJ3y7NilS
seRUnfJRt8rCwhFCQEGuvJnCH94wXFYfWQODX+u5+WIlgoLixEKHWuIdsQ9mQvw1wGPG0CNpZ+5g
77H5/Isg7UG+iUMU290/deGI9h71BVLciHwPkdWXG03n/dEovkygDdQqlwhaRDJrprCJR9idFfvP
RMvxcITDFq1tGnYjD7K4LKaP25KHKkXPuT9sDhg2ky9a5WYUJ7a20QPu+3ZeD32PPrbUikkz/VL/
9W7UeMd8IlJdVkyZWclfH/IOPqeq8/tRKGy4UXpB5CDcDYNR7wO91Xe6bZaWUv/eOBxYRIyaLFM9
jZM3nBu4AN6fYOFuxI0lSKsUu8x0Ofc2flC1DdD70ttHm8MmJ6qgu3Ugp4/6CQUJjTVZnusi3249
0UnpqSYgsRXzinaLDdJEVg/Ja2iCeQmDvlobiQLBn2KpfStlegxGIOx8V4h8L8YNMRGk7/Ei4uhd
u7SECCFFo2hS4faSsCnxbHJBiUpozu8zvbqSEDU920CPcEPrenzFS9VZoAKaEJls4s1OVZiafnMf
qBjCyMIqiDoMaGoIIQnaVfK64qlHs5WTOIObCjoc35H2gI8A+enUMT9ZAuD2Qbt2MjyQCIMX7L+w
+PVXgf+oOkA+77DsrvOZzIjzCgH1nbxRtbKmaE9lemfhYRIPGyXYR2RVjiaICaFpqPslWrr9HFuR
bNohKDPZ9zuTOgsugwqrxQwXdvMTZOZYcXepHpCv/vpYV7Wr8aZT5KvL9d67JDICm8R7vLHnppuN
63l69zqwhVVK20V2psH+FNA4r6lCPQJkBuWxLhqjiZyz8q8WbwOwQpdg5g5W2exp2hI9auS9N8oO
2mh8QswMQmxGl5heIrlJ2wWgX9AdgofqhtHDIKp22Vy3DtCfA4eFmD91KjJ70a8dAlxHvgCjnG3B
UrjQlcpRPtjSR/F2rtr3qVPeO5RujAxC0oweEo/1IT88EZg2nZb8RBNdwzgzVTbtihaWcir89Z50
Lq3lWON80wqKEXcB3Kvuysnxzh/wUMPXY9k/BvvWonwkuVzsTondwQZI5Yd5Eg0iEt01wQQGT38O
RTCfYytC2AeoNaJZzZu/0KgEhD5wt9gWrOzE7Yw7B2hB7PznM+uBs1BLwB+V9qkvjmAnSBU/MqaC
y6zuSY2WYQ60/iAJbh7hV41gDdm/7PjyxCHKIGwW79Da1WY1fqHgns2+gP6LT9ypnt86f2zdvP6u
PXjab3w6h9s723HaLjfDs9XwYu5752sej3Vhb7Rve4bkklsLEi10XLDYbwOAGRtMRljWgadukpPQ
5HFDvqZwNx9iuHLKLlZZWHfORR7863l7xkIoQrdULrB1RC+thA2QtHaGzRHlcXU+++BkmfmYfID4
9lsNe+jEVt4f+n7G3cXswC5PYqb9dxpNFTLqw/zCwAQqcY3fH8+EZxZlSPQyops/sJYFelnBD8N9
xuaCzOxzDSq/u+WDSXYqZ2KHIQQoN1x8ZK7S9VRTVp9FauwkK9+qbwAZJNw0ckyWjhNNy3xf4phY
oshXir6N9M+vHLSLYzPTotPRpztyVQ2yR8WzyI+WrDg9S1LzKjr1f9d6M7iRFcLka4ZkPY4DiM5k
fDpZ0gNKc6cJzIi0yYxt1Qq7gLIx2Ar/Q3ob2URa6O/8BUWQDkH4aRfW6RxbOsr+sKOM0fXeHY5A
vAHUhI9caLzWGyNrymhe256CFpSl2NpMQ3z5WKWj+oPte08hj18pcIulMRmiSsd+QhMUmjZRnAGy
rnerHAisSnvBWy4ccvX/Rj++F4qne1uhwY56+2U50tknEFyU5jKsdoUtuSUAe7TmhAGCh3twCvVl
OSADX+aTKFClP4jk+YrCPzwxAYCEe7/7csjxRYemv5MgPq9SXuczfM4VMceL9gmYsxQHNMJ1h+YC
5QKXTUuVHBpi9HBNo9xzUrRkYIrsy15XeCY9SwOv7SBXNdlX7o39AWeuIXViav40HmjrofLCVO3z
P3Lcj5PMSY6TuSUBaO0n8YsjRlI3pYGEmpjYQbG0CmiVh6yeW0T9JlEk4rxKSLKX/gr3IoMdXRRa
k5qVc61Zsu++UiAsWP1euQnfNXb9INXAwMafoq61CALlH9y0HxFCI04K8sYEXjexc9mEFfSXqJzK
SJ8q3Sr5epkthrXwfhtD7thuQMUIAi8e9+/7VG0Q5z8q59CfEO4xBHmIXcoylVcKNfQ8d5SVs3fv
oo4Q7ppPQccTf7Vupi+XCZauXnOPShU1kjkYcuGt3UPGKvQWSDXbRg2nkVR91GH0gRQg6mwMUrZ2
42pTeRhshnlEKwVbdqASNDEtUnus90ONSaE3wZEWf2ZufoGVALXSXEf52ZVsJ+tDpruULENy15OX
IEakWkldP+eisfCGuzROmBkN45g+RhBRC9EBQKstaNrRuegjjAVfPz5xbqrknOooQcqT9CzZyQJ+
8llHnXmSk8igAvl4u9Xjyzn3RdF+62Zm5FDM/03sWQ2bPyLH6Ay7B+Hr3dc8UMF8CY9G9Uai2ID9
ComwKwyA25RrZtj8t/pHYdeEofaUwwRJNEPEpxKIYf3QDili1qnY0VYbV6uxYtvdHz7lL/K8dHK1
BzOHavh295MO9RO6cUBwKS46ZBRQt5Knpyiulge7UOZuiq9Fdv14LS0xw8+mppYBMtOlHyqvQDIj
tpldWZ2Vp3JbTYwUjKm5K1sjeNQoIvQXaaEk4+fBTaC1effc2AN6YeLco/kjAJ/B706BjlXNW6Rx
n63dPFo1eOocUGiEm+VscXV6AzSo28TO0UeMV0xdZ0PHXM52CTuPGyMDs9Qmvu/DYJSrPnq2nY7C
ikqS9XAoRhHaMigUsDRzmgVwVPZ3Brm6RDL78lrFMC4mUfqbUKVlE07BG1gx4RJhcu46P98NXSfY
MEppJFhKS3GzrRLOFaylvdnplMtyn6bn/rSVLbploGAVORc1RHoThrvPOhAUFJ+Re/SsvgWOrpvP
FnYLGAX4G2VuZCfxS0nrWU95ty7pa6CB9VaEa/3ZIYLupUV1XZqa+ybND7b5CJU9tDl87hp8LhoF
g+u/j/PqBurkP0D68DrHsBDl5/2nwcvHpEsV/Yz47SyvqonkLHQGv6ghJGq+0i5EB94TuenYYw/C
dISyRRzIIN1JpPvYP2pcYbg4GNnY/cN/yEm+wr06XCPGSCVSRGVM/UZb9cpR7N1DhT+EMAdJ8iyx
wWYEe8+xqOJMWLj84eqREEZWaZE+YDVzIZhr3ebGqok/xF7nCqQfbGe+QF3cnqxvdFaPvfAJVmWA
83OzZrIt3FiOUzPj4qePYXCNggT9z+GhsS8cVaBqb6/VBA9eAttp0/ZZ45B/aATxXnCXJkmb8txq
WAaSKTr9cNiVgy14nbJEYSjgIuMJCNNrEm1O2wSkyonwLUCwVkv8A30JCtpEE2xjrDYdhY+67AqP
OB99EFHhaUjI0He83uy75jSZtC49sNg87HrRhba3/glN2xx50QATK92lEu4Ga1Un30/3gOx5jZ/a
cPqUuv5qSQhvV9ZByGxTOEwyF0sl3AogzHMJfCvrUbDdadkhUbboOW6FQ9areKZuw7dQwKgDRDql
5ICHWZtp6ZF8xagp6VDbu+H4YoKGYrcepI1xJ2IhiH3ZuVnVWTxYeOUWQFS0fAl8w+Ax2btQwCII
y2qgF7HEjjP0wWmaf+9cUyIHnRp4EgQ5wJaucZHq1cWOG5cnJbnPhRO39AG86kgNT2DpDjGV6s3L
oj43czUSvwxg58agJsio10aKPF6LDgnsNHwaAKoMGH6hh/k4T8XlmFPXnETE2i3xkYLCSD6M4gRH
mD2iVYx+9mrzWog2yuXfJDlQU6hqeEAL/ouA08sbydTSgwRXeyZcWPg967T90DCz2czmmkfo2uWF
RAiTCpqeZj+Xcbr0kvRnkKduykT990gga8y2G92+taXxJvrHusFo9mg/INIox5k3ygim/yW/Z0k1
obeTpNCxTi8eImumsfNlS6m6pXeqK48EBy7mHUvYWB8VhZvmpuw9lU0v6hcGyTd6hzVPrTWYAiHp
7vtap0P7AoqRa7VWajlkdS8mWClxzURgEvU0mUAb0E53PsiYwmL9CaFcmV2sIcxmtjzWc2xNMx47
WzTIyw4G9SFsIN1pFvsp9SjwkCp3ug3rmBDNMgDiJzwOzXzJOXi0J23sz1HwWvg/h4DPzxThN4YF
iSqiSaqcryyhiigEKyvX0sfsZc2iUYOq+eOaTOdhead0EvxCJ2hRFVVXx2TZ7DbfVZF/Tg+KQm/2
mRw/Cn8SMKLfM8P2+YtYBkw+eiiZfSRSzjGkmx5yl69whJIuLBXSQCZnJng0tqEO4rSvs6k1JSnQ
1xbEc7Cw02knZ+m7WH5vPBNmzzuyr7jajEx08YTe4qnCClyu36V8vvMAMu8HxEK0gfbG3GDd11FD
WZgBhAsV7CxNFuPg5/4H360GrssGHTp6b+aoEgKmvRUyDup2eMDBJQrNYhhMokI6qy+ymGIcvRcu
u95+Ugw18S/F9LquGvO2OGEkP1ZtZ9IqfHruzvXKvStSd99g3jYowYMgNvMI8h1teiFAI5NHJcHC
FO//GMo/IA+xTLPL9FKkbiFhynCnrY1mMbaJuRdIxUIgyNaOfjjMUrXkcppV7RU1g7z0JcHqEjm5
Ueck0qoVgtQLi+Xp8f7Q+OXoxD6vAftasabkgVMu3R5TboqQ1Jk/rmtLp9uzqYp0AS65fdyt6fz0
Ht3h6tnuxEIHoJJSCWgXTpeGug9+4byJblE4BHmC/ZCDH2TNL6xC9STEjX701pCk9XM46gepYFi9
qiRKr9Va285RDFcqTPJOZgPFYGfKXx9HtVi/+xKaSY0sAYWgDmS4Bc8RRCoGMvVrgEan5RBVRZhP
M5JbrlpFk4e3iyLF1b4amhn58JPkqEumxkP3KuzTYgani1Y0/lmrd/9sYa8HfcWj+z+OTRLjLIFI
LHHRYr8Plk//Jz9D/oUp2G9wXgx5Mt64OT2esMiaRbM+SWEFA2lxPbDg5gLKgaRJKvP3nQbolvFl
OQApjWKv3gOd16oVYljdwgNkAUGH9WsB4ncZoAKmYE0Lm2+cXvMLeJivUR4fYLQI7BGyWqSUtVs9
NvtrOPwyP48tEGzn9bhXbw7P1ncNck87XT4MSAmijvTUgcNisFtsUIo+nuG7oqX2e8lfjvABC0D3
KWuNzJcpnBRxjwEh4sTGDvB+Zj8rxxtYPI8eWoFOInOTAHzoj9L2KVE+0d/0UMwHjKIOkdKRu7CJ
QOIMZwmjcJHk6c3VAbfBpPLIUN53t039kEqPY8xGtNLOnfTOY5YINWegA3D9j/U30hbJAbbz3npI
ps7mZ8Ld3fuBJwPsnhkB711Au/QuC4jDFFOBPE2Ofr3hrC7kS6SrLhm0YNMNHvCHq8FGwQRGyb3O
1Ytnj2Ci8ZCQqsEI9W/QY7uGcrbYRn/ebPu2Yg92nW/HtHBRUNhvuBC5kq4YUY8P9o9iRDPiTmuh
WnxfAEgBF0/3IbnjUVQgAcVeT4oEMA5Cm+H9pgvleM1oyXGltjQGx4eHVSy8uAIGTHcC1igBnxU0
9GV7r9WlGweXpdAk/Lntdow+NTgWIueMBLZsNbjnZ+C+S4MBpOmobFHOWK+lW5lWpFJaQyGwS3ny
SOvK0EPZrgBSigWiQfq+dlhgm42YGhc1+bcKlqApk6CE4k3qcBnzT308MS3T5DrdJGQlfAdJ/ZuA
MS7SkYNGHjtbBYcOb7lH98rgcexwDFr1fPk1wj2ndXGE3wnpcxVgIrY/gVpjmFjQs5/fHIdHxdBl
QYhETnUR4cSx2l4DMVHiGdTZVd5beuX+AgYXqeXKuaolTO2jzGisepVC6ldaazDmZoD6EHCNKUyY
34tgUJFlv8Kw4Js0JRwGviRO/7DxKCbgIlRZ29HniZ2AMFvwK2QNYlimaJwdVk8QEmLpP20OpXXi
bQzwVPm3VP2MgCGUf16bbLtfrXrYxIbQn8GIZGwVkk27y0NpUMShnmrXZ/uEInes+aTrMkGplYgJ
1O+bN98UeuMQsxtgdUDcw24QAxr99et2c08Sn8cJDfTXk7NFds3ZMNGfS80Q8J0Bw+nI9FEQ+VkI
U/QlSy/fjeukPexqIRNtYlfPNJHfTgnLmT/T4Lta6yJXjlYwBT2EHINSV2PLC2ws50VYDxLJ1X42
S9Psi3RGfZzqNLP0caVw0+GYlAeVCwowFeE42GLz4NtwtJUGFO2BdH3lFBwh9Iv9ISoW8PnZtTCd
MMI+jNdQ530b86YBniRbb1AvQwC8ZR7QNvnzbeFYJGw1tRtuX6PjMwo+ZOeBybb4dzTobhT+8A90
GQ8QKS595AnwAWyKNLlG61nbiUaajEpLt4MdRPqw9alM3amOmafofWauu/b74l0MSyBl126CbOMk
rj4xNR1OI89HRBP3rmGBSAHK03GoxyxDkRePDpc2R523r+VI6aWE57avK1FIoGdTaYspMcC5sWZW
pkRchvkuZslcKRPtxfTveaCCq/phaxgkyEeJY7EfX7M5OJJqEnfwP9K+Qd7CBM6jFlOFSFslQprF
oWOnUP6NGO2CgyRWm8NUt87jYWuxs/aOelyhKKjWadOemx4G5Y4CNNF1DYSpvpbdbIAFt7uPgfN2
nXEBFo5KjMuf5TWhf3KoKE+C58PAuMKv0IOQOsdODTNfKzr0cJTqA4aMTCM3rOFBnV+IrfFUIJPL
pQcb5+iC8RXPFLCN3R03qaq3Zd6efU81/sSN+IWy2gv4Tr2eGpNsy/PCb4yIQc0myIUGNet1HoUP
Zi7LDj0rwECiotMdtbgecHs5gZ4mi/Pu8D6EIG9D6QlhblXlp2JwXGg5Wvm3Z+xq94hrkwSM6Dwn
QqXhZp+y46iqzZt8xFoJL1Vfqx+5R6S/c7l6u7JcjSZ5CuSRmkxeiHwJ69Pkn1zK1qzRrQMqJiEz
jZRqyrQSe39atYP/LLmjaAKbwwR50RKvP2GQKDO1RpXC3H23oEqjwWwd6VHYOHZI3zIcxlz2xWB+
x21fFuZ8qOxwVUOGrywRZrg39FlZ2sAo+d9dXEukk7lpwjLzNKanU82nv9qDq4tOANnJIVz10zNS
fxUCFMXh6/2GsubX8gOwcbmbU/AekNH7NtexM7G8EB60rv45KGRRX0wCUekktSBttUsaypBj29ti
ximd3XRzwMuYxJcL9FvnIcxUcs7uLizxI83T0/Ysz6XryCXuM5rRwHaBBWN0GhbZKtE5RktEEX9/
yDHitq9oxPWwgqxYwwjry6kArd+tOzQoxIqyxqCqK97GJZ8DRr7osKyC2bA6II73qOnYCanIzy6w
diwrYiz/ssLm7kVGv0PzZm1g3/FFqWuC/xkb3yaV9NBl4eMqd5B6Uhp9FMZSVsB6aR0nnE41Ywgd
CmZ3Jj6SD4VTDW/IM9cTaQ3onwJsfSIuq1z8XPuyAkixA7/QVQKt00ME5aX/W6pQ2Ysy5pzitZqN
452Ih0bbIg49Pbc0Slp4UPujdjFB35RjPaWl6ma3AKLlSfvqp51JbxZesZv2Td4NBE+j7B9ZoZoN
lXBLiHboMcN2xlv3i91IiuMZ72SMmTEFYFAEKBxI4QRtgLARpvhPCT8YevIn+ZWWSZg+upoC8U4/
oE8GQvterJJD1l56edt81v0Ak9Y4UG3QKs8sylsQc/mgR5tOqf4lIL+ubmj52ykZvlpXLy/jS0bh
ZTXABiSzulDyMUTS8L7AQQUIe1dHpnqGx3843FEDrp95VZXD4OiBP+hlFFwLM8k7Gan9Z1IYUIw2
s9AdmKt944bxH/zc8qS35Nqbc7xeKVOIFqSKEOW6qkE8JJaVaYyjbmEyROnDSIrPzwSSQZ3aTPdj
Px8BlGr3qAALsXjVCSE1NsY954jbgUfKCV2J9aX1nDshcqcLrO42gPU+9GKGAksJv/ykkOhftu+d
oQMOLxOMK4rLIq9+BnoYYWwwAwB8QpqqwFuEtnM5Qa3KwAjeLWagCdAgE5+we1wEGjlS8bVUh73f
YG2EBtHkC9GyyIq6fcxdRt9B7ClIdEnc5J/vbfnCoUq1dpcUrncI2qF2J0b0ksvhitdTFU+43IcP
1TC6T7bKGUxt3R5BRRwOJDf68RPDCqPdejmu6fSPT0YRdJXpAXqPIH9xDNQvQJ3SP2n0FFgOm+Ma
LZQ/iIfi9I4RB8iK2957ePCoHWT6CNamqImGwFgvDe3+AsvHeln+p3fjyQmTp4isJBMAgX0k9Ap3
lpVk46a6LgoEzzdgV8u+mN9sRi3ZHF6Gdzyk4FtkTaUwhf+9qXbJcYzNlJ6u8aPvX1WxEW3QkdzW
5XQSMy6fo/mcuam3Yobb1bpf/Y1wAeoFQ7a+QhxPauabQaKqH4RsLXpBLMgky5vV6rKnB35Nv6xH
B48ARVkSEKws36jrXLc484lIlx5ddeyfyFRLWtgzPO8yKT0TpIkebMIb4d70MEuUNCxi3fm+RUBm
jTfWmsayIgUiLXE51rTX4T6+T2zNNTaGW9nRRpyZEBocz+2ZLoCCI+tkAmCiEnQqdk+mv+5ZXqnM
pn9sadJmth6tmqtWGC6+UAyjnwnvcNj8ch+RbYfI/Ic6QnkS2igOmsNEVYczTqHKnmLS9CWbRQQI
7s0xnCTpY+4bn4A9pcivuxELI2IF8p5Z1PTyvpI09+4SEPoUpsnST/STCVkUWNck/HMxAReo5VMc
qL+mFKar5MPSIRHnyN6IrbYOGY2q1vPQ76tTzJ3k1YHc2vbPb0I6tZIYHwnkmU05RoyzWKEBoFy6
itIYDUQqFdE781lVpjj/HG7YX0v+gsYfJatfkeUzlGdrAvA5nPzEUfnHelpYfgz0hyhPPOFDb2iO
B0UCkUy6CFb0WCW4HmnRX7WoGtQfmSGF/VaM+UdNbzLJMs2sbVoGd8xNiiDSMPBcPRGItbXnMSgA
o6SQVafM1rgemQlZbZLlibUoeU0MRJmu+YHhVMvH9gR0oc9kUqyJ0t+NWM3LOV9YAPcWvXm8dDyk
3nHb7zIBnS5grlhvX4Z30SSoPOWwy9TowwTfTtE1WDvC3d72Wkp7c+seYiyqhUHyCuav6ycEld5b
NcLQp7BOxcEBZPQGvx+RcGawmFJBDb+8sxCEynsa5zkHM+tiX8dGKrD3c412oy/zg/ofqTtssCvW
5iphQOlUh7lKislZTITqo0rAgEc5WpVxHdCBJRnCNv8gNsXKdUimrSIg3qK6QFU5F4A8kx57xZ/v
/povMO51FSVbRWif0MjKTYmZJe0dcTTXmdMfgKBOzIbXS3xvPpbODHV4OCzugiRw8U8Xw/lIHEs4
MApXiFfloX7oMG3fmGAfAvo0OQPPWELRytXq8gBiAoQOc89cRL7JJ6x4bhls/AAObSwdFhr2Ia+o
++5g0sswUhq7fAXqusrXXRaMPCpd89FVSzluUJtIkdchQxiINYTXphEjGj8XY/8bdB5wRPhMwPzD
hpUOq0ImVLvGWBVr3ioiRtwFVsnFS7IGpOSvO1FLtxwW6mLySnSZg3hd7FaKYcPmcJHV879OtzQF
u28cOU5Rn6CaYU2uSUC8jMXmiZrVw5dGae1+JdNXq64vBCc2mh2DwMJhlAZ1AxaEYLQW/yRRcH/v
s/KupwCDLqcAf7vujGathtr4ug0d8SovfMsApJJxOJkR71GKMQR6tK6zdRobrVBKUtY+RRRVcIbo
5cD3WoJxjOSBaRby7fkbHnjo0lJnh9DTe9/fKZkG6rS18Ya0b/v6goQSdWsD2KPj691JjJfAX1bl
hbWN3bcxdBsszXa74r3eQZbB20f76oa8ulfHOptNwW1SmoIlW6mXk6Bi4RD4UqlMgOS0mZMb2Tvv
PHt0Q+dL8x/2Z1QF2pxZyqXjeiz5+c5TaW4htPi+sFcr3rfdYlAiGzQ8yARq3zHP7HOPFUDV4Mo3
pbV6Vo0mxr4rdu97CGf9Rpe4wuKzZSSBp2e1R0thdO4jv+pOwccrabr4s8zF4+b7qkP2qUB3vAmX
XDt9frKh7lvOXtcM7nhEKlvwmSwhGufp7rAulDfAZwIODOW+O18Vl5QGHseqekkiX25j1Q+0RIYN
875+i9Ve6m8X1fKVUEVcO8qiWXV1i6ceqSIBMjurFwV3UPu+KaI452vxTt9MlJjnTp7dzDaOaxa0
H1zY7En494v5Tc89DeIAjm6LbsWQy57geWGdAG5qeQBanz/9ShzA0WNsUnkHYDLJGet1648HFAMi
CActJLh1U2AfnkIKDqE3285ujCY1F7QtAk+VG0C/rxJI0EqDe9IwybQ67X96OsrisjzAQ+30JKvZ
vnnCgTrWvgAeYznR1XdnEASvbyBSB3d3IkXGOzX+gsoFiQtXfaJHYrQfMZQse+GHxgB5eDFF04Wl
WHFJuNMX/WXWUMcdMtGrYlRMJO1UzN2Ongl+qZek9KbnK0sb6jUDV+rLBrmXKHlgmN9Mn7dv1gn8
8agfY781S+r9Zoxgo9FRM65fG5iryCtDUcZTWzfQXFi8a3lxx5NvAi3AFw/UbvUwYyNlVIz0Hq2P
Bbl4XYQp4zaTkQLxFfpWQGyF266uhNqnsZi3dJl/BeoFxhMj+JMB9nS/U5ldWTdmRthAsExfNUjw
uip+E1wQNdSaiOZxihLdHcGc1nrklDOYojafW7gKhC64OTzmPQR8wIh5cereirOCtUcxQix1xgdS
RocpTgp3qjNdlDeGhkL3cpjasYHS9tif10LpmIt3J6UfFiOkyO5LvwBT7Gx1w6CgMzM9aoQC94gZ
RLMUfi3VjufuXE+1Gx98TB0Q3FPN+WxBH7XZtM0btngbUB4UAg/fzHigCl48RYYXmKZQEMm6kC04
a99LlQf+mIGg8Y4x1rLn9KKU4eBKZXteeSFVCkgZau0mYI0GI6Y6x4mubyv6YUpn271zcnS/d7Uz
Eu4cLCb3J36KQjR4vzTPpbudlc4b79TvHTHaV3nCT2T4EDe51/QubQRJPTonv7X4SG77sQ24R0Q2
xKGTJzl32Q51yWWCRzHgcnMI8wCVC8HmlUI7wesIFK7pmpLQyKj2KQPuAmqQt7hRyPl3SM7B4DY1
z2CqG7WK12slkD6dVc3mpwZvvEnEOGW3/diM3jnrWzV+IzYxvrKdypEZJxT4y7PMMySWabHCwxXL
MmKNvweTFGyO32hir27JAdH+k+9hoxAET8YT4LEDU9AKJiNSaEqq297FeVwdIvHMtjvN51LQFLxp
7Wzl7OOxCNKVJeORTtjdknTAqYJou7LAFBihkdZR5WHCR5TpfrZVbpNKc+dCxgwbTTnth9A7sWFX
N7pVnfT6iI95w+nL05NTi8QOWYL+8YwBF9yoerLYS02nkx6DcVLhHl20PhlP5f5zxlZBAR6NvvAm
JWyaVvBJJKsGEXHzRg3V5CT/SwBPxjn25HPaoUsUrkaKkAEjSTo31/8agYkMfaO9LsYPXqMwFF4Z
FLJQBH/B1IiPyhFDRbjMaQnTIsjGamRw0mWRwovlPwUIxUt/uOzSp+KBUxcCfFcouDr4mlzpGsRk
NQ9CDQ8gdlHHlEp0b0hfJMU+7MkQ7kUN1xk780/hObnURctaoolwddtvsk15QFjPUpFLZ603rHCm
f6KzRXo1b3spf5l4v86p5rjn0vmZgZ9XGjxfSbK0BSUuhRZhWbjZcjc2KwkGZpv1o4xXAtnus/yp
DQSqVFCWSs4EMRSpi3EMmLFLe80ILImizwFL1l09IoRaN7Y1woUiNzB36dnN6074iVgG4YYNT8rg
e/sBGGbxMff79qn9c2+MhbjQEbljtPGR2q8gwedKFgJR6q6IQB3oNoDo/y/v731Ha4ZTMKQMMtY/
qpoenEl+cUZHY/fOOvvIqKNhHY1f6doNp2ta2H2wBOSAQ11nPsrLWkH6IWSU1P3o1W9piSi3uCnL
UN+hlhYudg4psP+PbYLS+ogyL/fnQNv8ftSA3q2WKHcv2nenSp0hCWq+LHq6xI2hwJ9Zhq9QWe2l
lnEKCKKrK1YUbyGNgncfYJKWYR8/87KXGvntrezEO9gnsZi+sqTU2pPR2rZSHfn5Me+Jg/0HoX+v
waS0Jdehc7d5DeLF2LYuO3wIpx1AMsdisVgUoqKnjUC0ftAl6KF2pDGlvSUdof+as30umstRTwk2
zjkmSm6m5hJOqDcdJSH61/lqKwELPu3BU3sVG1glk6wMxWPpj9aTkt+LZAT0cCICHsxqURD8fOci
6VNa1bUiZKjS2P62HWScz3tDEFa1uKZ4IqUNLtVq1PJesbC1tOh1OTnOa/XllYAzgbWre4ekfhsK
0OZZWTeDr++5uWCs1LPlfHIlDzwnTjhS/XjMs5b3yyX7KFhWmuDQM+2oH9RlxD63ClEsQO/kSjVz
KXUXLPTeatnxHBzDyr9hUZ853AGVjIaKwzQWleG+d7zfSzU8nvn7T0VrvDYbSchel0xA4kp2G3CD
RvIu8UedgBZdjwL0X8BA+RHtDvqWFTIBIRsOR9IfenwQqpbkwKqGW3f/Ssy2XfmjTetx6wQ4XZOj
CNORu7N3CEXNMLw++kkoVSAY6RurflmiT0OJr3wiI2bsZoX019P+rXIYLswE+PQ6VY/+ymXOXomW
vI6b4msR9hV7GkowXQ2Y5wjyWOKg42qxHYkwLI+c7CmptJI4vZfRI/yHoahZs/xUn+K+MqHrO7Nk
rcpz9M9qYibWqNydY8mj1ObRu2qZ78+5ZLhnFU6v5SOtVuREWUNDLKHWAnyuPvVL/YAkHJ8QUgKU
DOitJY7gBWNgnJ4Hn1qdCkC1NZjPyIGC9vHTH/I0L49yOgx+sNrCboD7M6IyDsSYxuZ7rmVE0tjq
gX7VmH8chSjJMKDaAAt7lg2jmZJjt+WFH5nogQTyu+UN3sqr1nxoMBPZmCN7ACz5mSPsn1V/NnNy
dr4t0SPYe96mObNnTIiXy9jK8JR6/36q8HiP5AcQFFI8wynEiS0GjB7ByeJZNqolJsgAa2IoakOU
q6j2tGhOTjis6RIlbuUlxnifyJyBvX3fckcz0LCc2v0hKS3UMs5Vpqwv4I7OgpIPRsUECB7z5Hp4
zxAmbZ5IgDMv7fJcE8oP6CdIPrHlFHs/bUtjIz+XYKMg8WI0IQocDC+Jb4z9PycJdsoOqkWsBx4l
TpWcwwCQ9pwvVmKDxLtnuUQYBPUpa11C36fXVAs6evi0nLMmxb2XwHSFlzT5wwDMP2QvIJ3GJzcF
XGczxTIf4CLiRUOmzGifb9b3OwCZDDwC99YPKRRmWb4LzUCMj09c1LwKA052eoVZnCtBEoNIrRhp
+3D7ZWdqrCwTxYY7Ajfj0r+fSomvElDiR5ZxYg9F/204Ly54H4zBKDjqzX5/iTlProKm3gcLubCN
ROXsv3BmuqPgG+4EMEPbHO81XbSDh+Urqon8qozJw4KaHVY8mP6hM4pHg5X65HFBcA8kC4A3Bjq8
jGLiNZ2VY7Y0MMt4StFCymoj1kT2g5JF3Pryfpes5V1BDrKW8hdPXwRO9hndNLKHa+LQcWGkWZij
9+bvEif2gZJptB6FUSru1nbjUSmZEBNlbHjtSTTRSPbCm+lGADjx5Ne5Ejn7TIr4NeG9YmSbV/8e
NI0a7+SLeVFy5CZfvilvD3ajb6M0tzZg05Fv+RNTsNfvaiIo4wt/hmYYtJjwwNUdIMyHiw==
`protect end_protected

