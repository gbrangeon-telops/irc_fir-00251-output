

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eddlQ1EVBhLWIw/V3Y4jUv/9vIqrPH4OG//oOzrJzxfxJoDe5AYwYtf4Sd3VIdakKHjGWL10tZxJ
4ECEoEAvaw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eigFAyj6GpLic/D0LIryLMG9xQfLbNW2aTMhx8nk48gxIwiUUV5O0RCi0c3WxlsD0Jm/PNvkmU9f
0bvLBoFrSTxK1CBf237YO6kwoV8FPGCIv6uN0rXS9lJQOPdNh2ZUFAvoavKMegwZ/325WocnFLGE
+YU4kz1iYX1mmK3UsWQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnusdFYP+cjTwVO+sX1Blw6b4HVRZgRv6yA9tZdzqDv0sG/5WALWkeGj2iueXjyR4cWjsJaH1ItC
lJVwVFFXjpYvHwJ5RnZSqxv5F4MQSqH8KyPuaWJ7fxXpna2BJOvJUmLpfNOHHcM9ZtydeUw0FeC9
iaG6qychgs0JvDwxBvcNWeI54FWlrduydqedwrfELAOgz2Hnkk/tLLl8ktgdmAuHiBSlaAN8i7/7
Tmw44CbQzhCNPl2j2hqobn0a27C2ELHJlqNJpm8TlXqvKo4J8RYyFeM9H9JreJ/8JZ5Gf1n3ys2S
lY+Rp2WYXmq0OKzkZyIfymRWl5zSUC9Q8owcqQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uySJstuqi1YIYxsMDiwNUjJcaDIhlVqhon/QnlfUo3RyDfx9K7bIKjrz+E5jMqOrIwDUZDswr81x
cRDaji9FXOgh4P4INZOlQhXe8T+6WB7arsOA8Ipz2w1V2sV1eY1zPj1AXh27lapbQpMmsim+eCnE
1jY1XASKE/xreD8Glkk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l0UqkRkbyGn9mj0GavEkdTUw/Zw8lL7XEPhtCkfsrXvwKb+1KR5+77+E7EhE93Pmbk2awJRlXYwm
D65p2I5aXxW9fMEUNE0pZrhuaqpOOrPdC2bw4gaCcKb2BQm2PHu1PwR+8skPqiaBAqZVoUwFCZE8
LkMHYL9PggokRGZn1pk2O/ghNvl2eJ30v5gmurH3kQ5VEWU71s2ecSWfrCtyS9G29Ke80rPgnbMP
zifmkvX8s5FcVU1LeIe337473lbGtzk/tTh1neIkyiQD0Lkip6Q3stpeftQqI/864FlzKS35OASQ
wgYvGQgHNq1FJbrpROfsgNyTrijicXvjvpG0Gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37152)
`protect data_block
QxwvvL1y+ev/P4jfTxHCgllW/iKg5XuwDGxaSWqkMolNipUysKcPxjcODZRwNNN4SZfXrPvkHZQ+
r7MCbiPWQmyx/I6k/x39v+eVdJlnWF15/NlUM91ZonmKlB2lVrKij4m3mK4QPrtf3w/WlsEoWkJs
okeWEXa6kZKsZUAkMmljmjtBzdx7Pd3tsCL3KQU1L8lKKFo5eT8pSTvMfMle5Tc/OvULsKyBzPyb
/HzYLSVew9I5mBXYHPyieWqzIjXs6EbYezwTphEGqo6WS37Ps8BLvrTvDUCow8ivjXPc5Cm6sA9m
RxL3B9xInXTKz5aHIETFnbTeA0MpHE0h/3tuNiucPyY5wAMJ4vLfM/oRjwHY7igj4/Zazk1AoJO3
wXWX9YUY12u1hmrP1W6ptKqO3dWYUIEztj1WzF/VifS7Rw8Y5K4a1MWmTGvn0Z3iBbSxDIYtH5eY
lmaUoMi/B0a/l9c2f6co1YznHxhNtMG3hTh7/0PO0NV22JsFNo8NyYU9XUwI42a80F1E4QZjdDzY
zmg6q384Sop0XFveEHZ42Qk6T/X8Mr6DT3W5Iwuah40etbN9pT4WQSNShElMBemqfVuiW4DzEp9L
Jk8ZTS05OSwOaaIWo5FBGsRSmwGeG75s3V+I/0gQ1umwQ1xVcKvQk5bmSSDsClaUQdz5/XMM0a3A
5CQJVU+MUYDqDs9Ep6MQVItiN2hfcs4q31eq+USsdDVTSNvYMeVadf0rCWlVSH7rLtkWl5saCHDV
sNXvhqpxYAy/7pgtLFse9UxVoNhbCxJFaeP9MLJvwnWcsL7/xT3/74ocOJEjlgprVefjzzcw7Hjj
nNBV4688wcoOEwWj7HBe2ZoPokF7QekAaMEOz4cRs1IBr4s2YMnhD6V8CMCa8h9Lbonn7Dmg7gjA
p+8JnuCRTA86JtkAPSr1DCsaIUXGpye6TdiPTIwTOG1Y4MLPkbPS2qjcwu6wMy9Fma2qW6/g4fQA
fxF6hpYHfq05dEvFaL1If/pYR6E/nQd6FLRwng4/bkwADQrWzb70BXt/BYyh287oE/GiO+8unkVE
TEPveOpfEGf27AdBGMaY6gv2E8VdInQ7fQHR+DtkfPvHLCHl40yqu5nr1IoD07vLx7nnp4+a0cNQ
W+S/+eFx/mo8TamkkiKbsygjHrf7VlJXdARvhqqvMOM1tY/RNbYbEAwhAc9hObL8yBtwvfOmy0vK
eZtXU+SCAhZduLM2CTf53NsTyEOPFsO2oKjZ8ada21plFQebxjniUGVTbfeGahCQuOLWsPavUGHa
96+NgqMqxZ4F37u8WeFfLZ/j4yAyO/CalORSv2RZBwiTEl9x7oKhIo7f8j1X+CA5rZLWiGX+StOe
SH0IWYa2yw11smjSYMite/eCYmlrIxd9qLrCOKk3EGLKgAsJT+kx+z+aGR+aJbf6r0WbZTch1N38
IDDvKptVEEgq+DFfd12Suu+lq31SFPYHQwJEHidqCcvtkQ/bFsAsOM7JLKGQseLleDu1EByUPCuv
As7I34XmYT9uy8l7FpRGYFkQXNYAwtxPkcBrYxIX+548T7/XZ29VOmRroyRl4zT3RjC+SNxQqmcA
haw/TiXagKSk56oSiGZffxUBskiouVEfeQNPI+cLtxFtfv5QzfpV4fsEHLKj/ZOzwDBZRqfNmzMg
4oEh9De2kGzjxxpEnPweyZFRw8PKig5/g8b0oGeK6izfAIi1LE7c08SQXPnZxygY9xOF+CrPuVQA
UfXAyzIVf5vqTMcw481N6wj0zhMwKLgDtkJdMPEwRrPsaeJFlpNNnsIqW8EDYkzZ/y571y48L5+v
Az8pysOjXnWYkmddk4+P0H1jHy2EeXTZvr7VSvKG2bvghbYcPVoVM2/Kns1evUH/mscUi++awC2x
WcGK4Lkgz396D7XSDGtjMfvn6Ovi9BwGkcZazb5jKai0UpWBBMw68WmUv4UEzYHnmJoaU8hcnhk5
wNTcSw9sPlp2MD+u1EVT8QOdWMqiSHDpYch2qQRmR6JGRcVFRQA3PFwdworu8nmymDMLENl+I4f4
llU1RHKCmKUCxXnxRePTePQapftJbqiHxHslCvtMPEz8dVPOpnHbrjUE/jgPxUSKy4m4jt1lH5Pb
OdmLgpxRbwQVfhcOtTHw1mp5m9N7Bl6ybW84sb8FJAewhojWTkzpAcbRVA+ePwQ5+Ezb1D3x4Yes
rp6yhGWTCYYJdtVigepdAvHAj8M6OP2xIAWe43VyRKjuWGlxysLwpn7aA0QKgG7yLKZxhQQBvFAA
02HWRaFQU6ONkd/nZDtxRCuPKNUdkbQPCVHB5sY4ZH1T91HFpFm/HuSBGAT1cPGViCwlIR8Vrydz
mxPRzJYQdDwUhTTBbuz/AcjEzISbuk4amHgIBm1oeEG2Me/iefB1cooAUMmLOfyG1f+gKq56cfka
r0QCLabqyfon3gAznrO++dAOrifaJrcDG6l5VJMWTHBbEr7guRDxuV4QAxP3ZOFtymfpixuXaBL9
fFtE3xbAxaB/vFc2oBcec4MUPNX1Y3AQQ39GvkjJRaTIdW8GXWNOK4EHKmKS+DDQj/Q1TqkZptgW
2kdKJlxZ+gtuv5+kkLWwhKyiYD0U2rPuKf5ZGdWAMWwos/SfbOIy9kJ2TtLSYpmpGWkz7EDiE829
RofR9N3vKhrdD8zzyHhsWf0pyAnwDnYCn4RKC+m8DHpf2CSLZRt6MBHGLzUcr7yRJXCECRDsAmz6
yZXKv5kc44OtOvFM7XhX2sFXTpg80ddBMgtaiGG/pEimAV1WmNdg+kEXuLuVEcS29bmSjjeyhXB6
YpU06gj6NVXZv7dF/XOYAUc+x91bAVjWGWEfU1MO8yBxewyDaXrDxcz12ajyatDEpMyaK2areVb8
EJHD6yv1KKBnm9drmivF5r6w99Dh6py5VnPlngHypjW7IJE9lmERhi8uBXbrZkbZzO57kjsAP0gQ
6e+D/HYm1WkdxCfndmqDSN2kzkT51z0f3JB/yZ0CBUmWCRUoHCA/RiNgiMtSR3eSox1w6qCqbmD9
jczUdAG1BhofM1SsQN6+cfyg6KMNoKpvv+ncpKUlY2+ukmqqy63xuPtcNoSOowfa3m+zkrHKCATY
/inaJ/DuAsBB7TYzExwPZc+pam3zxSEemhQs66xEyZDbZx3/kcgEXfVYOUQ+SU16PmHl+PBXCCz1
TyHxMTi89nvZC1LZ7v3S1+pXjDjN1t5U6BPIu7wv2CSjTLwaBRpvnPrnCO2TNc0qyfoJ1IMJx53q
qopQWHzK/tRcLFeOSvK+zb69WxFlwoXP4+Q6WyqvZUlMOmcMbSBDoBUG4uq/EaZgywdWTHeKbi0E
DSsm2A9ybTJ+Atnq57nY4286nJHFOGAx9CLQ1ZjwlD9LWsA3SStzpbxPHC+EAdhClXxQq6fqQnE1
/FQ4PPB7Ost++jQxnkRNYRwuBZDRYM64kckJU+B29BfIbC5kgvSuCU19eRLFkdIq/gv42q3eRi3G
SeheeTbNSqUU+l5GXcppTp3Dqe7UDj0/B4l4CuhwSnmFH77Bq6m4RwaNa396XD8ElZHK3eyK/szs
FsP2Zxr96bKoFBeg9IShnPWyNhC8neyelEaQ7toj9lGzb2nnuWY4Td4wPx3VMhz7AMgwgEmrts8t
hxsE4ocpPcxeTcPd14ZdFYxAkxd0CJU75hyAaiiMmIg5egxo7FXipaowjOdkNTt3E+1VfuGzQUc9
WOlpWj8eaNEL7kAAvBR+pj8hJhu9CDsLmkM0ELRp94LWF0mhmsvIkWHl6ZSRryre1tTfdJEH1sko
5LuB+6jYjjFyRssr0HKW/F+9/JTaCxuX0pt0Uci6PnOmLoPZexeTHD0+FXHIr+TJlzp/MaUEnTP6
G6madQNOKPAmCq5JvEXHkOqqV1ohUw/mr4Ao5MKt2cgK8C77Ho32xRvyQI5mCgKAH8tWrL5Zld5D
82wK/RylPG8QuUdY4G5TwrUPgc5tP4AjJCq5jmqgXGQ4ozRMAOqUb9aVHEO0nFm7VbnTMho9RQvh
knEGzomcHnUSgO5fV5AOmEo6WfH5tVrBIPFbsneVyaUe+JmsaDDbkcWU9EQllG6mIewp/sXlYl49
FuEE3lVK9TDwZ+133pgwd3WreKSYITOB5G6maxWdvTWk6/POMSpCtdKO7o0BLtJ6Mb+qI/LU+265
4mqPOAWg2iIGwHw3rZCFWjPfLK9/v4Tydi73wx/MBV3Vf/bH8KkdYq69qRfzUmthiLR+HJ41GdOe
uaZdCxcSTCm0ME0y2KtJ/H3zeNT69uQEYxQRBk1vgAuq6cLILTADtvZLBiuPAC7UI9lvqEFNU0kk
NbQ7uiMLpCv+Sut7x5mwkp9RUf7JTuzelgjhWeccjgFaSHxjElMGSfd72oc/AoS1OaCwToFDBw/o
J6lOhGEec2RoEgj04l7lQzMgqMnflt5AVM0G7IkD94g113HIPFWRAUbrWx76BbZpKbydLKX88yDj
UuB1QQXpcVOcIWFIk8ibgv5fomZ3DwKfa1UPj+kNg/pHHOh+CFIuHj1vF1jtcziVwWRXF8XVVHlR
Fap4wpl3Bpzk8Pkkg4/buvenN7zO8RBtDtX9CdnxxRkiX0sC/0JhCoPr/Qv3GL8qEQH/xMSDN2oB
6wz6bxcTfwGIPflxKE3bUM6svpNV+nrOWRwWklvbjRf6PXBk2+wGd8p2JC4+iLCcA6k2TnBIw4JI
nMsuMNaKO3sxGy/o8f+3ADpTHlenC9kgNnm5hsez1DIW1y6dZB02dZ6KwZN4M4oD6LeY2bqw+mEU
Q1+6cYU5dzBKl8pCKD8usPoE1Gti6vVRmdo8q1N+UGJMuizDclDufUbx/+Gqi+G+M8nqkp90hHM2
mbZXyrNVePrdDpfklGKI0HIiD6wet1Tqf8b6iWP7JrXhL//yF6+tz6Lnyfb+h8BRYcyT9uFlS1YB
3VF0bFO8aXC65Fi5jdNnneEIai8s8JbdJtAKnypCFIKfWceiGrf1c9yrkTizfNMXyP3Cg8K8m1L3
0KK/2sRHQh/RmMmzzWOLpzRmm+kbrtq9rdc5eGDgFSAFfRdF+oNQ0pd2q/ErC7UhbBrEsQA/g3Z5
ycwJpLVtzGcBJ8IBm2VmH2ElXvhKOCmdG+INpMARdYcl0E1mQwVwampID1kk2RPuLMHTypvut+X/
/xg2DFOzdBKsAsQVOjAQe0vuDUZtlQbXaJAdHeTPht5onr/bVLjUjzUOudHZ1/Rjcdsi+ND6Kq+k
LR/ipH2wsG2Rp0VdzIBa/Y4OBhcKg41oW/O9X5nZB1IfEWnGysfzGjVybHaXFzcJsOGVX3U+vEew
2U54EIcc3HdViNh2SltfMqq9Shma4nDl+Jt2zfo9HYB6MqtMi4+0JfHsP1ZQ0EBUwzQtAtGk7KZp
mcdqaKQ6kUaKU+FoYYKjIZpqsAnf8jNNMVislURGOZCBygmDY0qL+X5oIdKtHNqgdIEPxTWFTQ5D
l2t9wgsELKl5AHiGic2OShi91zMhEpCeqS3sPZSp4fNFphbiTqR6wGlP1rCDiwg0OEffuQlcd7IF
gPSmjSpQ6mjGkvgHtB5lW3EsRK1vHbOpEOZjc3AfHNSjTYMERz66ihEisa7Kg0Vc1ayOfXUYZmd6
yYn8kBqjGpHpYsvWYNpcXDRvjjP1hHcekrwNh7wLyvMhtjuBrrrHO3DJ/M3gGDry1MOPvrOkGUcU
GOV/mQG8arkqFgNVrQ5MXGiebF7oxha4fNyI67VSBeVxXCw7JKtBL0JHlA6yCrV7O7wBHvudKImK
ik8e5iRQKa0KaDQY7mmNz2ujMYm19IzYf5d4Q33PsoMn4an86qhXqABAMRtmY881UbcGAL4ebLQi
Lxn6m4bNhSt/7DmD1bX18Ep41Um8mPt53agZvj0yT0K3E+sWEw56P72OHDha+8cjjkfB5n3zIFn5
fP2vuCEMKeHq0wb+yLRinre9y0GcUIBExCOlfSR7qk1l95l4pGwCjOZVRRMg059pMLEaIpr4r1nJ
tACMKnC2O5snyY0nVAYNY8ElXKGI9lQqhm7Nc+YX67nVMF7kCHIWxrX1oEnOGDjNpQr6U62qDiQW
BtEWR4cY1e30x7j5Am8yfC/RYbhCtCl/XeOx0BLkyNuCMi752R1gKu/qU8c2fI3IHUcQ1abbWVPS
NH588Y46ps8WS1sIYOQgwXJpiXRcQmID7TvPhSlncfMu6rT15gCrelfWRUqICe7Dk0bsaQCA/zC6
qPxoE0vPww4jAdF+awk+jrDmX3iOguUArd0AvAgpYY6CtV+BH2xxA4DIrdPgoK2RU7kijj5341me
HYf3mPunUW/ZVpawz1cg8b6iw7bJI3oSFL93f9AhHTaKcneOw1N3+KgOU2FQZhVZw4Wr78BhMh3+
zBXlKMpP7N6aNcY1Xckju6wTOu20Ym2LqmXr+i1v6WhdGIeGNmvB3lxd4IOLCxKHggsfdA5iC5DX
3ujMAsxunaC+qFgVjWBcfTfDrgaR64rfObGyAv0lA2ZX9svUVqoPc4T7CfgAoFaIvhrdajypcKLx
yGMDkXm9cJvHfmBDUVq1CzAUNc11FBz1xGqypU1Td41trawC1LOKivl6FEdMvO7C4LLW9vqnJ25Q
kmY13Ue0f4d/XlAZjMtY3gojf38DXGPZsswQh/gXvYdHKuscLK6uyM8Dev/MDHBhGupEZeAZBlSo
YVyOytmOHW65T53D2YyJSuasAh8gaQ4r0ErtGFvWEN+Src7xUHojNjUqa6K7P45UERTVtRsHWblw
zUk/cY/Z46nw+JJ83Vqn9W/70AGeuPoHOxkX/Qjme1jigLirKiu4CsTL9ZEUmtxW8urSyqbeesiS
DkuKslsX95MYEogx8nP8TIeYZGf4cRvySt0MCVtevFg0n79H/9PaZ3wmJQdYfT68xgILlvEj0wZP
a6ix57vRZg6puFgomY1WDZKO0k6Yz1vW2pX6aXXK7X9ZoAXHpD9wjGMRnJGOsqhY50Ci/KjxdHdA
Eh15AlXYgK+N0geUy8clu+5et3U4sbE+8oyCODhHTYskqeqTkukJEwSCLtDCZ9f6CGNzlSDxpp9N
RPH9+JWSQjXifp/75PeahPti0IrkoRsXT2PQ4jOwqcDcF5aVXwq+A8MqYo/KpH9ESG5Bd3xHP885
4AyYEBcA6efqrzLjjP/CDuXFR9x0e1Y0yzelCZat8EozyG0RRe9t3zRS1PHWhKjDzqB4eWyYWB1D
p24sUAWe8309j4mUVBxYDeoVeBHo7zFE3mXOpr7uK5my8j7cf6flfwvnulQbRjtXD/RBSMoL8fK1
1tmzMQBV2j7vOoSnAMAb2xla3FCGxl0ZPd5dtTayIGtdux5S+UdKQ5Y2w7A8DZ6F2spb9jYRa6Wt
qUOU9nO3zZ9lXyVmB9CZVip7PDuRLdylBybiriLij7z3dJZFfhsD6yvrxidDg9FuDkWL6w/UFs9C
CHo0Vz0ddG/wiGv7vsvZyRN7Am9MDhcy1U4RDxA0/4duzg8rX6fMHsrYKDEylBJj912OtcwFzamR
XPEfNm6/57I3WYGgEqi9Y8xYN2HbAFYbhX6X2Q4HNv1m0PihRncQcmW/py3fmi+W7g2D/fKobtZJ
jBP3sAS9esQXeJGoG+1RPgVTWHb+sZfVWTfYF/w7hi09PG2Kkkn+aAD+32/0nnTKYCfP/7gJrpSS
RrUaWBVpNxxorb5bgsfoRXm3a0zaAbWNISrGo8m6zPGGgGROkP7HlTRLPSumneFMMAmhDzRjtCIa
xY6Amj3HS4qNtVddWwj2GmghNb4YzszLEbf2z//6Bn4dg1R2T+CBetxUW/+fOfcsG0xrgmx5E2QB
TTBe/48il01YhQkiRFHBlcMhlDXqzI4gnceR7IzYRDEQEVGzFiVm73KptRlZJcOd0FIR2gSAnRdU
dUwPBteD+vNx9yRzAcw4EmygZad+3ltoJWgh204TnR5pLwJWpH008/ueKu+kNZha3dn+CS6t4F/J
G2VR32Ge2LkQ0dsqyYYhP1M9F1EFZ1E0j9V5pKmeMCxOQvigGVTwnminXGmTkaE3LA1oGNg71sll
UjajP7t6vWwIg8+yoKKXPOPDKhVX8CZJNtW+ZvEnDqFlAasZUV3LX9XWJyc8gKhKsABlQe6NTxOy
hhGrIJfOlUNy535uF9KUX7P/PgeFsrF2j/Q71t3crK+31dxAYcPbxsMWTMWZH2J/9sreJ4e5QpsS
eYEVTjDP9aCHAhpXBwyCiUZXAAkge8PdAxYNQyvRTGg1Tu053rFFITj1qBnGwenU78qM9h3QbLks
GydI8Q8TJEMJ1qWLl/a8HVV9MBIWXZspSWXCWGmmfGSOolTKN3tdwOtL7/zL2UozOSUEqkoq52FV
ChTJvKoNm+3HFu6dOgNZnDn7/La1veIrGgvT9K5vXhEXloRCfMWxk2CVjnC6Di2vK+09t096fmBB
jKcyGfaxDdNQJmPV/2eb6wKdbYbchLoGqyoyOBhz2V5RYvl+O3GAEAW414YFWCegbwPLVMnAMTvv
ZZXGBVSM7TpsygsJ6I7kXafMdunF/0eWr0XijAfypMxLjHkmfILbxSnweC0Xga3/pfW+leIzkTN5
gpu2iZGttGefGvH3vGBlHc7FtjRAitxS/UUYM5eu3lUo0xxmQdy6VzFRP1SOfXwrSCF22cnTnp6H
001FlH4IkGNzpkf4UP7tLVkGL0CbGjZX8fZvb+yQxuf44MwH98yyuKDASVpms/A8WXVTmRK2bV0t
QPga9cWpGWPmt07ZaLT0ZPrJD4BEtGfYlukdTGNqqR7ify3oYtHFqPM3my/f0Pd2HBRZLO18LVaF
Kn2qNNff59abht5e58HdltyPM1b+/Xcq+RDoOHicmo+BOBOVhkGkOlhgY2L2BIdICJmebooPsh0j
uZWWw3fUhbtJNOR9lGB3I2Wp3cLvg9tBwV3sd/OSuhBvQCdauzwGlT65dVAX6ijLZ7iGJhvhroAp
mi2Q+/dFd0+nVnWvUD9mvpk5HdbXY4xXg+ReEQM1G0QbMebw0iZss3zdjqQyQEYFpBaHAFuzDB7h
g7pbhToeC2oxoKKv1ibkrBB9w3sgs5x78YLfOr7Jj48zpkmSKHHl2bllzlDaKv1LX6ug7uZ/PnQJ
Vhcz1MaTEE+CZE8y2dG4CDVMjUlDmT0aTS2lHbqxg2AoB8Jnuqg6G08w3un5PjwqywyF3Mw8MIt6
+q8o7Sv8wSA5Di2uy8/c+T+Wa879tNW1pNBdPNKqIEf3/5iuIoT1dSvTUl2rGpwPDmBFe93f/Vw+
cJeLJ76EfjcdijMJlWYeZwoTVOLZ4ldOhscsLdLpDrQEK6+zMMYLsst55t5xqKIRjxvvW5ebMbcD
BoeKbE0GnIDdwTZ7fIzHy+4SXv+mEtxEfX0hCnU9U5ALtcwNuFAa9KFIa1d3eNVwjrY1Qo6YTRee
QkadfA2hXG10r8m3ZgIKD11EsbCRabSCalhhOwFGLZYIJnRZ9nVscTKxLaQTqa6ibDzH9nn4Ktt3
L0OmkcyLumZSHGcAlnil31s0ZeZJaWAlHPx14C9my64MSdr78ZIUai5PXx9d4dl/eS4W8HxiB4O0
LU8fUIIf4uLf95qFSF2aqDtoJQutb+vCvYDPAuSQ2Gkbfek61VagZ8CIjOxoP4Fbkc4BIVsH4gOJ
yxpuyiqvIXEPYC41H4yz/48tBlskBazL8spbDIyDCobIgwI5keee/NAYymRXnVZf7ZoA50W7Kzc6
Ufhb+42OCUEvn/C6qA7+fXGCK0bSgZGPqvzXUKb3LE1IhyhLm3M2YWQOhxNP4Nb4nRuXRevf6PaW
w8tQzycxENxrkmLwzMfQdumIFK4EKf391Io8LOcPakZXze4BU13JDB09/PcdxYCQNVpEgMk8IYOA
8zploeWz28vKd4Yk51bUJWR+AL7eyP0kykdNuag+u8FjCoDYNbbH+zVGQPXmZAggqMA3cLdnpKIz
H739C30epwu5FiNfvCJoWhIHYU+zsYjUQzqOjE/x1oPWPCuPGaIp2VjXde7h9JXLxdDZ/VWvdbjB
KHGhY49AHujF4k30NOznNK6SFEh9qajyRZvYwIoerr5YklYiDaxC2qU7mbYo6ag60IduHgO+mNrz
5YWNmVUa+v2ohlPLDr9ZUNpM+2nzMk1ll2MKFMcfI7NkmkgHSsKjI8mHaYGKxvaB/FwEC76D/uPI
jFSsK4MJVss/QBRRw+QNLuJ9jDQbwhifzCaO5oWIxpFLlTGrXhdFUCj+5vkzS23fcVavMRezDqjB
QQwN5mzpvVwpY9Rd+zEGJCDeg90Uq9Hd5tZm1XXyVT3ygKUKPVjh4FLGR43a27dnVnB3H1K7Omb+
o8V3vqLHhgeKywmoYVRwwr5XmobSdhtzPWbAnHHjEEpW4ryaRZ0AHvpP4GBgoPdg9e+4TRbz6o6e
PYom9ephBf2Fda/jlPf0gYQ1tvSNYCm+7MG660cWJ+/ey+FZ2ayqsvm6gxE56gg1JR0bAGb0CvrA
3dHnxjBn8B9aRrKx4DubI+kjnki9tNaeTLDJDpdRKaijhvmlpzHFdmmtgJRYNTQz4LvXDJ4FAsVZ
Lh1S7bpOoeWhN3BsivK9xUPfUdfggIVaoZTA/yGCdV5JjmpqbzBA6T6vMMGTRD5nrfnFIGpPIgNc
Qo1+VR1FT6wv911w9dzT3ETHNqMODs39Bq2rWQUzYQsutH0eac6dCtbj+jPYprkg0qFpGDGP8T/V
9yCagIPUSpi3a91uBVqc3ZFQQI9MBtU4mmBCDD2h5bzF22uJG7fV7hPhPhiS29hGCIW3yIo/R9c6
MCI7qcnS8Oc0opxepbpCmh+CZ+/U7EapBlwBN00271ObCg5RWW8cHDHMv5ncdCIwKtyn9/+0/gqJ
IGPEmNVAtNa4Woc1NI5vkTP+A7VLwAYAteuMf+bdjcRaxgZQRT6K3uopjz0sFqPYi/0E8TVFQ7/e
Eff4ZOxvXqyHEvIzRdPRvLqK11iXqAYdsQWG3AJ9lkQSCqRpTYJWnxS4DB7+scOfHeD/dphXjBmZ
IL1dgtvDOsrrm4HPcZkpE7fHvPYedLgJmq/OCgisxT3gcbJoT0QNI2sWtL7zTHzl8Xxj77HZ+POp
ojk1B2DISb3UftApkKt6nFKddnoGJQvtad1aby51MVEptTJTnpy/J8RLnGmIk9KiIvBaXwGfDWBN
R3ozSg+YG/IHN9jvlpsnwec3dJ9nAtWYsgjIcVgWdriBwi0LRPT1pcg4V5sNo7sWNnScp9krJ7Rq
VLudoRWFiRuR9Yc0uVE0whOMCY35qCW/7cJXRgM+7DHhCjLSrE6yrvvLEcPeCvsTijf+nAzZV41F
kszxG5OQK21jRxR7ou1SczYw2slxQvJrZNTjiDjQepVA5TPeyE9UgR6rvKI4ceAFwMVog3tifpBb
lLz3WRxFZfQgb1VmjhEOoAVW+plwIdiCSFRWg10Pu70vBuRmNXfUoLwDsAQ/9Tj4SYlU+Q4ie9K8
M4DfePle1tqE+txXZOPFqHagQx8hGib9DsD8FxT8Ht2AoIbZMqnYdl0zZcXHeXyONrFmHhvaswu0
hga0IOu9f6AqZ4JfnG971+XoeJwx0O5VjDQjjmfFMG5BzuNKREZAukOMuYh+SDcAODwGKz7QPQYa
gx8i2hHAJHFvvGbCqzu5rcF11BD1gvVxGfSAvasCDCm3DovYXMZK9JkAFFsI+7oUIslepwE0BLaG
v28nCk21QMX90Hj88qp9py9/iAz2OhpkbZJeRqS3Vd9VUBODgKHIsdM/HeYuSnkoLjNPI95CXn/I
6DFT0ZBy8QN9h4xmvxGLiNYnDOAY8L3Ot9g9oCiLMKaGoaMuD0qdZ0rtoPgcbeW1WZbPuBeHuHkA
hAzh/qYz2u8qc4znFku5CGPwR23ZNSio0DJMS8WB5C4lK/5AhAmqxY72VgjEaSRpNtGLDlMjPNWK
lfPAgsvxLGJBfkoGsBmd8XlU9ZOSLRLnahV2cUQnLRw3W2cSD3TaX0mrYfIKhVMsAmYXHn1WbAMB
KetoJ7IhMvinSyL5guPKtbB76eAklpid5t7OlU9nup3VfwZPc/7OGboM6XMsBreQld8I8fKhXHY4
ckn9/BuIKw9h5VGAGqOW+h3Oa0XvgDolGG1TtYQQLq1LI2yL7Cdam61ffdoSF1/U3ewBeAlrfJ17
fPAmMvsX5+UOIwRCmcpTwmJQ/R//yAEq0YY/OIejvlxYohKtnCvOYyafN2DYd4piY7ymFNIVKPX2
y8VP+6HhyZ5Mj7AJVb/ROCwzo6svEc/b3MkEWEFunJ2mQhC0hpVqL30liMLBg97HfRQHRZxgFIXH
M3Z3lF2LD9IZFsA/eF2H9eIMZ3Lx35HhXKSAu9HqKCKyKySxvjRRd1bvqzjOhR3vQ09PX8Fa385O
yVFTyORc8J+Ngb7JPH6pa26Fy8Mn1i2DczDj5mYApDz/B/r8ECXVIty+q53zjjtX9igAIfe4WtA9
Z+CKPToXOloOSw2uPrRYOUgBSIbYybnZuUBgom4Xvo9WoJhHv5DSoJou6kJsrdTUax8kgaT7D7tx
lZTBQxChhoUKupEwwOlu0jodKhJdACy1Y4lYRDN8tN5Yn6B6+rud+0gbDAqERlFP/IHzMKZvT6qn
Fe9hxcY9ZTMWh+OtsRbPeVVRb5R9zlRUyhMbdASwjazD/hXvE99Hj9ekCe/rrtYD1EIPWOWmlvwA
qyZ5ePYYpGYVkydZovH+i/tud3HKKfU740qD74y3jxJPALsQjy4/c+uml0F3AoohEVbpPcB7W18Q
mNSZtc6MXYS9yHK1ctiUVmNW9l7ON2w/ynL8MlIVHV+zg2wFGpshpXWcvbMtm07f8OyfzGU26pm8
MSPg3yw4o7C3OPoyC43EeVbuxVeKTDPZ3WPeMg2YXY3D/pERxwU7Fajv7bVZDxvCsg06ghAdV3Bv
fhqIvsbkpdNFoC2qb9pAN2k6ahxj/JtdOuhfEosR3wnZRP6EqXGzZ3suaORSfPUcfZQOByEgOfTG
KH5boh0s2kr1CStM9zCHVdDCmcIqItCax3TR/wLTZt0aZEteF+pxx8dcFfO4QHfMTpYaOM0zFG/C
92ppZPmrIoXP4lppqOLiEN6YZm/SmYPg8EBuyfxTb3wj/P+0drsJIEAuCRiD1krzm51h/WVaM622
8gB5HaG68paSGgh1w9sPH3/RKErajH3lxEIxXNWZqAmxcPMzTF/LhOPrGm6lbC9TbNF5W/ov+Ze8
ou6xGJV4vif9Dl/sKHn6IVMCy1MhHiaaag5Sh0R9/UQZkSuRJVSYiDPP1Mmk7ou1YYJn7LIOhaRw
K6c83H1AWcitihNH3jcuWkVGFWRS239fRHerhYSUY1GOKIYu+5GmOYGB35aK/3DP5Y9yA6yz08m1
UXukRk+1vDAnoowNqNGftpNwFHslfM82o7vBGGozP7p6vKJAIYf5ZdmQYF8//nrbvIQqpGVcn6fO
6w52dCRCAX8bmXrPCiSungeIpkApQ+V65aNMSOAwaCeTyF3N4AlvTBfcIPBo2YiLKFBdWTxLttij
cUUNTcy41iHAiRrvHpbZu9xpwE6Iew1kFyOYm+ahDF080+nHVrlR13zxMwfR6cjTrJYVyahbvxDj
XzgqujOdVmLQNWC2jaDnr/Yz+dU/2ouJ4b5eNu22s6ZInr8PRXUA7KlEPCqjazLUNh2Oo37YJzDP
DzDHxHnmobAAgZQmXVraCvIeo5Hg0a7Ep+N8tOO3FT/InLn+Pez7CnMy1Ro14cuigCqXl64xmtFk
nTFtbE7GRZ09tYJD6xTU+/BRq/n8c2czBbEYvW0+P5BmF4voo9HJDQUZgdyDzTcD7ENkp3rXjU4o
NFwMsb0SLBUs94r4olJ9ew4rgo/0oveD3MNBFBp4T4u8NC4zDwB3/Rv9CMe5ncrUxT//CfLVr95S
ZpjWPWCNW33CaHrARKT+YVyyu2n1S8PTguKrABXyrpUlerfI8yzSWoWS7DOC5zwmeUGQt/jg8xXg
noqDwTjQFolfhjrOL+Xi+M5ahe509Rnt2gZHrUUwBsKgSd6b6VeICCXXpzFfORIrILkMy82cw2gc
BIFZ1GiGcuR7g2TDozxiKpG8zzE2KltE+crOeSHvKA/ZKTsNFbB6plzQOABSryVrxOQKvAWVoj1g
7RzhfnV3zNiEe7o5fBXMg85fE0QvoSWlBJfLbck0eRqMTP3K7zPbvqtzNM4P0jhxn2hqM478gICe
g1GsKfBEJ5x4IOP8CKwH8sQ9mWLsZs0YJQX+NeBd768R5ZboPzKc1h/yT8LBCHVeiqpoPu9cKlhx
Zi6PhWs+NxFEPv9++ccgwfmXgZbl0goDbuCI3ECvi0jd6MMurQA7wQkSNHIEe3uFKtjHFCP7JxHi
W+StvZ4syNbaSYbFMlwcKLBx4Fejije86wVYxMgelA74dF9PR6VLwtc/j6F2JD7HlX/X6GJMpPGK
arhot3VnOa+IDN1/2ghleUxW7AM3efZsvYAxCKXJTXQ17sTgrcwnExpHCCiksl+vTN6r2RiVJ4j5
pFOBkjBGLBr8CyZ8g1zmMDhR00JZasEp1eJVQUerZcSLdT1LFpU4p7Q23AlQBoqK8scc8ZaTKhHJ
xbyx5P0oOW7S6quXWqchx1RIX7Et0ZcjiGEeTbBTg49y32/1tJJIazg0HPdTLMgPmjeBDv6dP71T
Bb6VB1yabNEnSbqMWCnobZGh5xXyv+yWdtTKQLoswJUnZ1w96oH25LK0udTyYn1GELeexKLW2Z1q
jaJOKGovmA/mMkugQEf/ThwmoMpDeq9JgufWt31jb6ZjBBcdMBCPhXY1sbVbV5u3DwH7CdEVqPM/
jW0bpZGV3IPBhT2b2npQw8Y3wI+ttsEjTv+PGAb4KQMdS8otFFi8OXZyuDbjrfSqHVHWIXh+DNK2
GQDM3qDjcsY/AkIUH4nY2jJIow2rrfnmQMjbW1/T6YsyDFKWP3qMLnwONYnmr5GoL5lMqVXFNt+w
xaAumD8HXjbV9Uq4/P/pevQffvSGzEj0DjI2hnnGIdJiII3Kr2p/upPcdFE3Lh8CTRDmPZazPvry
0oQJzyHvr05BOMB7ZLffUhOb6JaCm7UDN9fGF2MfYgUAJXfueodQAQPAz2AtkYVrNZIsabrgB5G5
W2/H44rmkTatJrRtfPSdCjQJnovwklFY5ye/zYp2AT8y9VaeH5iL8eKAJrlv17hOk5MP9M0+tIff
wT5/zlDVyDmJHCv+AKPdrs30EJ7Ga5dWP6yNaB9j/hK85ar5h82/z8j9DQmzydNmw8vaazOioeBz
ruhckYXM6I+UtTtXH4vQIculz2PhbCkBYkTcplb9G7c9TfPtmXhC8UiYQqTejIDa/UFsGScKlJjK
VW/EmDik/r6kvYH5bw1RGofi5GfkefEv6TJwNkZmZ8BD2Ngu6T1z0vkB67WRPFmkXtAptNn+8LSy
Bhxi6JVCB1Xr3WAK/eGZoj89iEg4UUDSUBC/Fj67EyoqR8oIxhAt02yxB3bWEl109TFSGK5NepIg
r0yIxfcVYX5VDPbcNcH5pGFqDrF8cIFe+HxdpnNpIuvCeZEdyDjJ6Fgi8lKumYZHyc7vaM9HU8W0
DJSyXMD49yJsIG9+1QCEdA/XrWqnB4WZosFgu5gT03gNeNQPq8aG6qnn7sOM5CkukosRKrhw/JgL
vi9SIlX5br8KJYLCb3yhL9D9kKMnp2rkG0rEh12EysRFED3yV3cbG2cPwSRDmnsv6H4hlybLD/ip
jF2WE9+/iHOS7E5uiOXwCGvwJ8hyVPFvpQ9+5QWNVwCZ0NHirDqMuG/zzrrSpzEbLKEE+Db3PvGQ
pFnNctPzthbQq1WWCbw/mdDwqna4JHqthR8SY6S7Rn/yc1jkvtsNLT3Empq5Ga7bBd8HBp12MJ7A
DQLN/8zmd+JPYLxKJaHIXmL69Y0X5uxAUXlEyg8yEPi0U55myVHN1LJokOqvxiTCXwH4odiIq6ZR
0XOcV5DTMmXETfEKzZVvor7rkBIJn/W9lO+zN4IZFMX4A+GhhOc2bB9rl+BrrnQvxf2CChFfy9AZ
Fr7HAVa9CHsUomVOpiCftczJavnM9PEG0LmSEmxiNkddKrF9mFzMe4oATRU00UI6NdzMBM7uY7OO
8srI/0GY9PjR+VBaJSAhvYsdlJGIB0XGwF9q6IqaqOTUXX4Fz2Plu9x0KHBsYcf+5RLHXBQtQJdB
qCMzOzzVO/r4Jd8QSEYfxDkjKlv5agsip9bDqU5HxdKkdmlvgMjJvS7O/QHU3vdz6pyHrf/AGuMc
E1f6nRJnhiYbTH6yvSqwqC6okXgCwIDkcJreKbIs15VLPeKdsnbpgcL05FU84+DtLgWl5RSyv7Pz
wq3sEqwNrzlsDA2V2PETImtIOWiwOe4rourW5NsOx32YbTpKpAMbWBZfsdbGBVsWIhbhd2tW68Vv
h8iY5EBXgtgSP8Ee3y7XqJRXWOyXiMJFIQJq3KyQLpuEwYsOx3PxS1RrnrM+bW1m/ksLcZCW9sTZ
/hDaG39PEto4Jd9N7f0qVB/ZYAzs9KvUszRN7vAfnXf7d+eX+I0ytC1zVQTfpaRIKZXGbuxVqNnb
lZ6bXh/dvF/QEYQMdGXfkjoVy1Rw4z0oMRhL8NUczPNL56mwTJgjgg57M49+cPsGtXwUaDeuSQQY
5eYVveAs8BT2P32TAZ8zf9gzLKvLCM2oJQANkpeghlSvdz9Jh1g9ITW01kz2/c39IH0pPjl53cwh
U/Kbu/eJSbpIAYaJKQEN07vyR67Wxt5vG/iWkIz/VHo2MXX++n8MkrZRvhISJTIc6uN2ZKll8Qd5
UV/OnWlWVatJPwDgU8Gtl7LCpRuzaz/vZTOzwMRe+pBZS6i+afgcszC8x12V8nSNJR5G0mTqdQTy
xkKx8fJ9b5pSnxv5OFw6xx0yNhmsxYcIfT+UH7OJXK26bBCW2aRgU0hf6Ht6moFmr392zujF+/v8
vzjoCgVVl0D6nXKB8DiIP+xIcYTtUyJtvVp41y+b6DFBzhbBZ/y+2qc+Zz3QysDToR2Hrso8p5C6
NZrGEaMvvF6+a0tMfHADxa5tghWK235loJ/XHxK1DqejHE7o0+NQ+znG5861sBUlYYKANgfajNjk
Utxv2npBEBQxk757E80eUrTjsdyiTSk8acObLpVq4kf/CeXvDlWDl8y3D/nF7Pq1FImZhF/2XvFG
gnjPng6GvM68uFURapHac40zmu8J8tUXwPoPANwyoPJ5FBiUIV12DJo3fj+8qLh1y0jNEP9ZgMGP
k22zXkme85yFjgWqAUZm5bR3uRNSVHPfvwadbAge4hxI3OV218kSMOf8GzSw/yhVXMm5nRNphuKQ
dpLb9Yb6F5IywslxTXccHVia4hNOmDcp60FGeVgGBqJMABaKG/ecrDME2DbTmuyVpt1HDBmv8vmY
e6qsf8k0zU8f/xxanuOS529CftfVfkw8DaBccmYmBvY63xvHcQ5im8P6htlouQWWcFIFC7awfPdX
4EPIyuxPw5drVlEelVMF9t7oW95ajSD7izfMq64KZtBzcSL88QcIKzLcbrp1Cr2nymAFs9ATl+QG
k1I0jYcoD8OgYvKWT6iYEsqyP+807ivlSfIsiSFWYq0k92cBI2KAE7d2v5cVrJv5ime3Ely1uuPa
ymQdnxkWk5YIa098mdAROKuCd+vLaM9v6gM9T9CdIirZbPbsrMwGqEY28KYR7Hq0zjGNWM6hOXs8
AgTcDtUlB6p7pt/kzClojqWhMiewm+er5+nnmC2cc+68M5gbVhSdOj27g8DaXxatPvqQwCX6gk5/
l5Di30p8yFqVe7hbvxP7D1IaJ3c28bs1Y0sK+r9syHXqGDhbvAzfJqG8xeB11haywvY6iv1k6fW5
BBp0Mldes7cSXIGizB1arHHTVHBcgWo0z2y95zys3zhCJr2+86rmp0zdacXK+OR67NN37nv6yt94
cJ+Zo0MGE4UZDGwTHDy1LiFO2ni/7HqswuOM/Sqxbkfz94BVces+tTmwxgmOb+BgMhGM/BcjmjCf
Fv8cVWrJD4Zg1wqPTQRy4cHM3YrH1uwwXYF0At6rlLqmA5BX1AhxrdPZ0eCHCLR4lZI2stDERrUo
d4YWoCD8NJq5kzgeCGWtNcCt/2pgKeMxnmxTW8eHrUE13tbIbpJFoKMR/7QmzYct9HKx/vt/JUnQ
y6RMki/Oqw7XYPHhqSoNqyG+CKPQKCE48/qCA3thDPGRFk4wInBCvXsHTzQH1lytC91mOCl6iJLo
MqbZm4UpwkKoBYtyuSxqF/l7Uv6x1sxMdxEN4Jm1f12nTk3ZhswIgUkd2w5/vr/yUkdO8908gN6O
B2UrKAH2Nn4gGDP5i1dtIB2pCAvhlhPdJxTw8etlqIIwHrUBqVvXdFSalJTABhUPlBuOvhXISoGF
C3mMYshqg5gtPRT8dNEDIS8l0VaVndvklzXvSvMjKiX/ydj8LGyMAiYiVTFnNHd6yEPb/um9xxJR
IDNa12yKAfrH7ylAVlfPo7h1FZBcOfbSS1HvjISEu/fbZp1lfnMsE2nIImYN8yNGjk8tiM2oxGVs
L14V7RG2GPLl4Qk5IBCE/CRYYFuPS8grZUfiv9NevjK6a/6rKuDZZskWwZSE/ghnSQ7x/Z6V4ks/
04AaHPZL9QPFRos0iKUalGUy1jCKhBna5l27rS0IwC77iXDOSU5Aj6CpczjahPftHABK55JsDQFL
7LIszMfg7luxsfgUdc2iHb++kRQDv9941mf3fpBumeE8Age3DN5fKf2zpdH4mYryDlfyc7zWLSSh
DhL752kfHInjE+9NtC7cZ6CskfZpHfhf2tKQWK3LtE/UtpVnEIlWFC5K+haBNdrBxuX8BRUMmbqO
Peu9o4V5EXKSKQKOIoZh+800NHUZJtWothYv6NaByyvtmcSYxsSs6r35Ffovl2KuCuRnLiqs2KXH
70e+qCdo8suOKqy+2LfLheoZY3AFvaNK3cudaE+NpPzrRG8sp9FwHuuMSbzeptLXbDtATKQCrOs/
BpRJgpBxXaazHwS/k5Gjl/ScSGCkUZGECGuc8s2evMDaAvs2MAiHrlx8N3Q7YpExuAcxvo+ZDXOb
zYA/2N2ycz2YlUMtAJbKlfvkFRvPYvhokyxDPpQQZhmoqonlYTz4TgoO2itZy2Z5axvzFxNtI5dX
iZbKK1+XJyw2SIf84dWbe905BwCPS7OZuVRKYe9J5Zgqvx5/csd7Zw+L1swoqWI69Wg/E9DJdF4v
Th2JiGS4KXOp4TKdppJSuudQ/xRj80WbAI7mMrRv2RA9dVLo1xIKGILBz7sL1uKfDDzoem6ll9vA
BiUHgg45NjoyIvqmud4nqO5WiRIdq+DGAbPklOA3G0/lHn9Xu4zocKg6DkDMG40MfIZcv52TEJxo
oKmGc2b3h66muxOCeaKPRoOOqNE8S1S5PHIy6zH9H5NfaxUx/hziu3mL8Gx51CayQZVIkyqwpZU2
S4s7Kk7pokPxz1Mp7+iJCo59sc6pIwdjIOdoq6agIeBGVr76hShqckYVXp84DR/Tf5qyBomT3pzq
kLNynkcYi0SBt+VvNEzkemDnJn43/D/xRtl/rUKCdXLR0hWTmkPb4+o/YL3yQI6+S7Tt6y7cx9Kg
PVvxkojhqacRQslqyVnJpwfc6fCrGc9YfmPwYKf+FOCMkY8Ls0uGlYleTzGDLCSDcCYLu1L7coSv
ESMWWzWHtCa/uC5McUD7CD5j6ZhJhCCuspf3yh658F9pz7IZhBaGX5WL8MZw3zMdJGsKpqQBwBVo
c+SzDdC2UL+n7ezat2WnlWYwjIaJkzX++vIpXNGzSTcxQ/QZHHXUc4Hp/QvpvYZjOVNG+EuZGZjd
qNPckZzHKg8m++nSxnItqLlEOFjiibIi8rWe/HMLkGad5/lnobMxdAxNjiP9ww1HGXy1cln2+jIT
lVbLOukLvn15wPTuX2bKoksMCMm+J1tEk/5huY8v4ZpCtKlxckLT1W3vG0nZoOxbyEkcT+9QISlM
Go5uIWxwc0O4M5q6EfFU4uH87CkKMn9anQRJhCgv/5vfRtTAq8sPJa4mUX03Ld6veSGYzlHgXgio
/7HnKb0haBm306waZSyP08w6Mel8vtixlVZE7QxQgo2elEXScuHhWfhdfqAk42rjgKSb3cmPpIgC
NbMU9Z6bVBvGrHFWL0KXTHo+WEBTgJE7yqUcyJrH1zg3qJ4yapSZa0kZvGNrDAPsD6J7bLsUvIaj
FAFGRM9TkHuDKsbZsOariNIYhYGbBO39FIR5/S93KclEn42Df49xOlklHq/KL5gFs63BxExzowLu
AeooJVRybcG6eaqhRBBnW8MZGo/slXXERBXomEYUcxMWa7f0otmeVvkel/us/l5BsF4owTOeA2VU
dZM0bVSVnINzCpMh/oiJzhs5R9wotKvhclb349IbaBDBw+IlXJa63O+MAu/JGhXU5X0qKgD1g/ce
eRVQBo+0HkvNvXopkaMcMCVi6qEdptZdFHvsxJPbBttopAekbFy8bNUYaTASHQ3nv3plBL1MX3v9
VfVA9oqA6edbmX4JF7B8ukZsX6zdPTw9xYBD5XTTZDF/sSDJagFWRqe7dF1I+r/j9e89mIhmkriP
oui7IwbaBL5E4Ra6uDAK/ytcgo1994/HfealntVgCpKGXwYh9FMn1QMzmVK+I92RSalkKk0Ir+ZH
N4ANuSScBGqqZ57pRufcDGySaO5P5rVtg5d/XHzlDnf33+LVvZas62qBGcbZQjzNPv7s5KCscbth
IUU9KOZM+YnNMfxZXFcuormOlMwVdg+DG6lp/GWmhUFepZ6/yd9KxlPW6cQylKCd3WzON2Uyz0mn
a7/g9Q7nCwFEz0m22+ZUFfzFoaiHK/ccljxYXXztozfzo0WUEO/EQ35OqDIb9umZmAP/LKgzWFhQ
0rBFxksGyrWhiAAU691UhlMGLrHcJe1SQwM4mtcxkaRqTQV3grtXjLuR+tA49Aq1wy4HxXWwtVz2
KlMRpVC4ttys5xDLYnmM9rtrWdzhSzJibdpHWZ129SMK2z9QgJfsjTr7ov/CS5a48no7xZD4p9xo
FRwFNZuHcbqyhtrcnjjB0ER1w4boqHKfueoJNqR9Koc3qmQ846cVKvN/tSGNJUH5mMOy7Y7RPsQ+
661IPPUZTEM1au50ksvC3H8Fp0qq793ymM2aRhLGGnLdwgcrW/jO3Ld/1L4MJR/vkWz92iTF8gR6
wINdcy1PvO+7Z+ds7u925hcxbQ8Lq8DJBcTVIZGcOhLPG6Od39rCF+VNMGSkfDZcCIjyPCoNX409
S4DSyoSS9o9zwZsaPf4bf0LE7K3QwWld/hD0vjBqk2XLEzHqbnLSUtX+WIyx0xWVnNOMW5anSAMU
jIxrIJ342pS5bgUFdQi8aWavxzygPz0dpVpf2+EFy0gva/7jFckhKLyFCNW16dYWwehwqAzVRfDI
VJZM2Xt5sL0lbz5S8dae2yXXeg5CaOjWHVacHmGnlJIwudEN7deZRfTbFy+8p0FJiXJpZzPUPMLA
2LICH/uxLYzqhtmff389fZB7VF84RTl/MRLncR4SA6hwZiSu5N6ZeBJiJXn/jJy6w+KfG2SvPzvF
LyV0+C7ZCIzNSMC7Yr+vmvUdH4u0XGIlRBgb2MDyObKmpD74+H7/AdUhww6BomXWz0zy0NIJi8Bj
aATIhf3xdYUVpQdhG9dXEr+2VLaW4np1SLMsHPN7JrL1I+me+4Vps4GSWBRnSJYpjTVMN8vBe14W
7sDaFAxYNJv50Oae7pwLtgZJ06fklgzFYLCpfPHpoNz6U8S7D73z4Ot17VKw5c+LWL9CAsgka5Vk
dLvi42JDZgrFvJcZDTFUz/bgoA+2nQ9vq7pKGcRH3NeK3SSnolpV8v2UaXWpqp/UkyIPq/y3brHr
gyr5PZ1WLEtDozeeHIiYz/E6yAOefXuYDTzNYKaw4yzwpbjmYquVnznyIzI0Ch5r10jYUagqLClB
pfPpth3+np79VubRdBu3FCxG+QfHT1LE0BvKBS2Y8zM74ynB7UXBdefzrCsQys3MdXzsHITgLY9e
Tce5bOy5NtD+/NTcWC3kI3ZzS3mjbsECP2n29dOm2mGyGUXfdqrKEDuPTXytj4WK2GoGFEzRLHBq
3iwqdUCDSEpJj2QVDIQMEnLtnepzE6tWyt8+B/ooPOHde/hMn1ntJ8nsDSz/ERuMAG8JHq81HgQu
PHzYEYoCBbtrSelpRkQ92ttzyXz+DhsilFe12Hxw7lS1lY+AxPFaKAuEXStLWo+zmmYDA/dssVXl
BSRhirRFmM0RkGzc/IaZKkVhvfThTJkvArBMGgbYr7imrrIuvDI9EQ2t2aq9da8xoZNAp96v47jc
LDrkFSgAONclwPvSTs30PO56craY5kltr/OWJJZYdnAnkGfDPmpd57Deuo8lyNY0kIMw8D7lTLNj
u0GCZ5rWC0fmux6+WFaTRNYXPGZL76kID1QcqMP9Em+a7kQe5IbIKN4XzJohdO8azwEEAAfHk+AS
r4trvuvPBmBL8Ipz4aqH0kg3lYa1O9KtpwupviJPlE/3sLaXep8zJoQb2WkQi/pxuXykFXSuOWuO
3QcKsjHoOYzERURmDujLsaOePBgMttkEwZuzMJX6EDAw6guLY2zEV6crmNIv9QpGw2HEr9iJm6K/
Upk0s6dl3t00wkEGbkhvERoKtYV1wtNeI1qgM+VndCURaq3IcRSOWa47qMxAbJnNka2hrNLAAb5E
maMuyl8X+Ac5xP561m4snbNDk8NsmZ6C03C0dLIxXx3h7gRvOspolE6nw01N9eJuwZbpX0KBZJ6T
i81zlEALurd2b451ps2iktB8AsI7etfeHj/FLjSoy3ndeA0a1qdtWquwGszqRrkLP921A8grKTm0
A2YoVFmCCTbaPT/+uQ0innVQ+m0uueVkr9wIdA4sFcFLyNPtsgjrmLnGxb731iqF+U+EAGt1O+P4
XdWwt8Hzf1iIrD6OLjAj8mniViqgRYc7EAZmY70Koz+tolR6zPLKYqdi489uoNGW7y/DoH5sLj3L
61DznUgO3zjZmYf34TCJbdZeXlBZ9+SFlDHH8l2IMGUrwSB+aBhIz2G4NCtnXuq9WgmEa8XVCii0
WW+2Cv39vs04ow+btEcFAAbPFoi4HOc0JpEnrepku2n1xHX+PzC2+M7LLub6t4SWXD7dDhFBI5k5
w/m1YomazRWHYjQHOV/hsJGvEfti1UhM807L5BknmMWdk+HAg0hmjn2fTMm27gaitIlQgLKiOPK9
Tb8HCL7v9ImKpj/UEtpmucrpYa3LnaanxX/7f3DKpTHgTsMm7ZBxRT6SLw2MIGgem3OeR1Ij5BNT
5WZi2e3AoxZ3mIECYTaPjxMc9INC++feuDy4fvDE69M8DY4W5vFLwIEx/7KNfTqiqjvL2a/GWwnb
UGJJRNWxyONQw4YmyQ7Jv5SMrOPynRAC51ZTZNceDzIEkgawG6vTsZnRDgQx6UeNRdZioDXCZdGL
FNXZ9ckSZ1NhvlHVH/R4YNcBHIIlHggD4jLHfwsndJTFQo3qZ5r601IGdtXLglCXF4B2pXqII9i1
6oktaYk+Q1gQaF8/u0K4t9UmJprD3TAZpgo+1AKrZSxZKhT7voUC6SkMCWXPXBczIlkHCaz/hM1h
e62tktNOtSO2o6S5VeFlJWcDxlXG5gWQxsGue2/u3vracvNETtBce52aDyp1MeZZr/xrAts+WfCA
UFxH+Yrp51dDQoF4u6TUCsmLfif/qYFMXkm8SOCFUoe2xI2YAoIXArV1bAsYfPLfwNAJP8tU0ok+
/fGoE/PvU9O727LTrh+GfOOKoWn11YqeBe6WASdAdxPf3T0AkQoXIu8Htnvd6R8lgVL6TeOZtv61
OC8j6h6CV3cLGtqad1VtmbC1vw1+47q7CnwZ4g1XFrVRNNQ8kiGwBc0ZPGxCTerZ1T1dRjGAdTIw
Fk7B7coSrUGlJXSxbMNAzllZKvP8Jm81lB7mqjDWOJvOI+Mkp/ZdIGAfLq6h2weguoEu15Ib11F8
vkce0sJ58Eec2Qjw+CHmTqizdn06RGyiYAd6huu+fA3LEbwxXX+RDTAJEcndxhFOiEXWiAlFNcze
DCz59/j+hUjfEx9uIJq4mA6Yu8/nUh2lIkZmcz0oOkG2ad+VKwWBIhmN1uG/3WX54juhK6IBSjNA
nt+sSJUU4ZWpk3su+XQiXv4AR1AtgA694yaWXHyC/uHdXfpjCqH7lHkZs6PtISRB+6xIU9acfrTk
q4gEFANcCYy2W9S6zMZJ7HlGdIyKZ/1SYPdLn4Xy5JNHiAcVXLNtWNQ39JcQ/6wZAo29lnr0aLY5
LazaBGwMeH3KNZjKvVCVNb+2jTPGUZKD1Ipuq/Xq0ArkRkpPdcMOyqUDkLUHGnG/+4aS5eaHa2fy
sR5l3kIXqjKZGd7eipz+Q+1yYRybXvfjA5ihPhPkMnVo2g0GsXJRa/Tq8VpJx3IlCXiy4xX7RCdH
lUfOEHQp4FwkuIfD6m7oaARZuCplqLbb4wtHZvhszrywjtDB+LRxfPaQVvtQUYq7TuROzggxRYZf
lQbOjZkeG9LbzfALLC0L+TEPl5jx6wxCVjYrjn/Rn2YLTa9dOffzfg8i2NF3xx/IvhJE7Tt4QiNW
XAXk/Z0w9qFAx8QNuR26kvxLt3Ciqj5yp1sjXOHP3AqP12+Hio6PP1NyD/ibjDl0WEWEVribtl0X
lGsM87+3N9ztQ32ZcXvjU1VzDi60UFo/Je/iZHZ+6bCE5sP2+gjnms5GAR3YgGTmp1OfKfysIezw
dy5dLNlqi/G17begROmJ5Obt2I68mPgcBAY0rXwqYGdXmRkLoMDKIBS+WPop+ptGSKuq//i3382X
dmsv+yWkhklCfGRBLbJzGtQbUM9PYKZY8ti0usvrkkU4Ohrdjj2nSkFJmSi9li/hOH+U7S7vuYfp
JyyYvbWP4Dvo1l/sRNcw5zXakVdmTW6xaYoulcqi78WQ39TItvcUY+m4iuLMV6gV5lILNeMzvCm8
T8+yYuOnV6b8sNHBr+C68fsk3a3kUhi0Q3SwxC/4MNKU5grQglJsJXNeCAuYHV+Bt5X9S7Um4m2P
nldYreY9ABfzfn3Q8CPlzFLhgolWy7cd4uvhD8iRJO9qq5mTna84HTHEL12iuzFW4CIotSQJH1tq
HITkj+Adm73lWXjcSowhwjQf3PJFtsjNAa1Gb3kpkTZLwR5Z7hXRkzrBo99mP2gUIaWadP5QUh3U
OBlCbNaWn3ekkMkbveJ/77vhPm4zQm26roT/lN8C+rQz0RhW0kUaC90svwGw6XSUsZFCv4U7xc6k
jiE7wrge50Y19tDTFSNctzdwWFJuMewngqFOV6dPoa/PBp24Q0tDZIYYGeFbH7qpGdoFoQyj+dU/
Eg9EmKvgCmK5zfAET2cBaJzlwsjxnMzT5ecppMa3Rowb3x8NAxiUzB0X6yFflPJBr5RkDBck5AFD
0xrtLZqG+Sh93/eEHtYdxs6cefowDMgliivOJ+FUWOf5fe60bOTBizlwP8pTabTt2u8XcpuM3EAQ
/5MIsCx1b2yafhnkT/txbvDLXEUcSCPypmCipwV39WM7R0YOOXNaKsz8v9J8+AZuddeWcJhQtv2S
UqSeK39Xt6/QxsvcLevKXb4Y030Bu6e7unnK57MVFqD93cVPP11kOo16TZPNA1DQSbCKUfvJUaFM
Qf015X7MK1Gcu1a12jyLlYa2xrJ4OS5G2uzyqiT4KyMsEl1qZeCbT9WWI2qO/TsI3in4+viPpaBL
o2UXBTYutUBF36pUg/+lP3J/gY40hnXaFcGi95HCDbavQABrBwkapRSrnzzGbAvpB8FnjbEmg8Nv
xlFxIQOkmgKkFZUgoDnnffJf5OXCki404g0OM8NemaTXkw/Ih0BN68fvIvU2dlBpmUzzJ5pUyMqB
6vNAazNaWUieJVzi7zJC55k+MPrhdul+AyMCO3yBAIEEWp/jMma+7lZnSzlQMzuVgHNssYC1ihen
xlEt6s7+HW2xsROGADpX0TF3wd0/NsCtDQ9aXonAD0CuqJchxLn7n2aDSsGrej9H3/ZtulpWzUbm
HDZHb/Ly5d1v0+d+xqDq9cwiLnMU2Dw0kBiAlRjR+wVbeL7jtMNZLJ8lr67Lfic5x2SMtcqjvI2C
A8WnxsG8KUIgc3DJ34f1Fmnt8jqRNDHTD+gx8947rwXfShK36TyYj2NNrpsrpr9ejbPEi5nyhDIt
kQLQzU+y2/liBd4skPn9cOrftfFmk0SyLFg78qAakTtMltB5MCEK7h0KFLSYP6nAZObCdU1vA/nW
1wyRykoeOnMyTmmV6MuqDcBGyP6JVjPqH2ntX9qkhSwp/k7ra4KPiI1315qAO7AyZ1gIkAQtks8j
FP6ks8OU1Z6/O0PLVHOtBdwIOEvUtrsmrzZa5JiowjobfxONVyCO/xBvAa69zuzlXh47CY0NHL0T
hiUsPADg7+GVyXngwnd8HZX0uKwBwHgtV94mG/p7oDmokweCASx/hKb4I4QKrqksaVTefvTwW7HG
VUUZ75AfUPKhvlWzBKLq5d8KI5n6DIe4R3p8WxolgP+D/upQxX0GJ0MhrSRF3Ek+9qYMV34AHyom
gaZIFMSskTHarTFagwrJ3mjcpe/hDvikOZHMO703bT3iWgaGBqJvLNezaRZkyvEMYTPf7hRKFlQ5
aO33BpXiWn1mkImfESyejIaCp4u3XxXsQe+eq92JexrerAlCJxgvlp/8hnExo4sh03BHoegk1br1
U1Jipzo/r2qG+Jc5DMPX8mnOHPF1ENPJWuQppDbTmQgZ8nNZvk+V+wdz1BRKQ0y1Ez3f1alIIz9p
8+36TNm+uXQlgKCLj53LUr/8ZnCJdDu5r3WxDDXbSnw0rETNxXtGtO3/ZIa8s6VgnGhqaUfXgZP/
/LsYRhQrBEXmMgV+X2kNmzu8pB/4hxZ6+FoHZ5gp5OZ2gL7YrByWiv0XPPbH4JVAj/5CXzkwB7bT
wkIhSy4yOV7Na0FVit24usCTEO58kLlOAOqUqiboNGyY1ACPHCJDW+H01xEaEZOjWRmM8piPVw4L
bQ4mtFdvTG7BeSL/9q/Kk75ayAufH0y5WaDtz0cYbu0P8NXXOQ6Ka2dVqnBe34OjsfhjwcQO2E+G
Nik0dAeS/yv7Qq+vyS7NysRDaNGVG0B8TUyoKRulT5JAlmzOS4uVXrWuro28hPI5HKzqZevE6qxO
Xhqanqe1hQbJMk3YmFvGfSFL1/E51aYtZTINULCALfyFb1go6lJd7Kq2QBKLEsvNlNNi8Jl3JYtR
0BZIFjRiKA+EQVo2LBaoM1IerbnptcA5c5zNL+6ab6sJic/jUwoTt7L2ONSuJZGtARWCHFA/9KX+
/aBz8Y382Nw6v5MUNJckGvdME0FpWiZ+lmXNVSGeykelYMsNv8laAgN2J+z7AkRM6S2xQQanJsH+
gfyGvYiLiTDPMt6vw+y3c0bSq3XDdQSC5+ydchvkpUzI3Ynf9nZQDIksFzX6/he0lyCauKpTNIHM
WOLude7lkMPVjrPlYv6AGwIn+S4CdTIku4HERr7dW7CHpq+NkTN+UcLGKv6KBIvV9G/DVxPHZGVX
YaNKPUBOgugiVO4ml8N9mJrmUylLP9TGKC4hx6yv94tsQArIxxl7sDyEFc/dW/wTQ3K4sM8hoDyR
iKIDZTdDTxoCer27yq+ouTE4bBT/H2pn9IAstSKXP61nB997Koy+26Oap4hWA4MtUNTPW5a027qE
feVJNkM5/xo4WJQMJaDFSrBbxgCY4rdxbGm6Xy4O/fwDqSyXMiJ0V74OcHomA1dwg9FAwr8EmQ5j
t/t6REVynWMSvIkMj093IWOCwIrWFzcub5pXRZa1sH3YszXDOcKqIafI+8JrjAp8vE0AVb+Miltw
3qmSOW2U1poihScmfbST22u70uluIzOawtl6TmUgFZpdz7927+lxNcoUrvzeaW216pObDXA7lDZq
hUMZcx8BM3KmQ0HjEbcedmlwBn2av1Jvg0FRfMbOBrBlHFFC/UcpvRWWZw7W8g7T2opHsJ27WJIP
IYOX7dw2zqDRmIOCMfACpf0jfYOgaPOeREkt+C90QN1emcQ1UnbwFnhHlafClAgjfiMAv8Y5ih41
dJ4Zy9NF6lbPPUIxcJkL1E4U3/JrmtUSej8THvBRfu0IIYCWdo5rFcGYjl3BNPi2ZNx3fX9wUIty
vgiB766KGIurZx9dDUABQVObQMeNhNDciUGbaXTGVqw4xQXGoZKdzYLn4TutvkI9eVwPNKDrCX6f
JtFe7BK4j62QJ2UZf6TA+dCBKlBcgLVHJ9XnOK7uxaDx4ElJA7Z3C3cMJIhJ86EcSGrzDU8VjRxp
dTMAeHRZedUMf1YJBcfsn6defwYd4J0ZOTaoIL53UvKLh4aqg2cDzN+x/y4QPSCEBDUHZ7Fx6a/o
3rG1RlzhV5flOmcIFt52xWWNsMtAg1P/GTUqm2LKWRNuzjhoboikfQlOVZopC/fqYCoSoBw2IeB5
OFbcuTYrHCcbzlteC5OO8dZAK8ravDsztviQWA7Ddf6iVpydjMKZP99006+oeq21NlYG5Ug7ayzo
AYgahZmop+SpFaANDnh97tBoFVslcz4JXTlETf9pYJpXV4neosC39jwUzk/AQLY4BPFS+JofXtmd
JGy9AeabwRzyZbO3OhKrDRsJqDHLSsK7glgHmowQK+k8aM3Cr3naxVHwdU9fR3d1Wlph4QikDurx
SlJXWCWx6GUFLnzjHKTL/atDT4j9+b5A2+cn54MFhjJulpRLE98vvo0LFwDKlsfUDKUe5/tjUcAy
CryvHwISIhzHx8p2jfReXZ3xC7Mr2y6qOTbfYEk79cYYhEINRHSDCZzKwVlL3b9h5l+d7pRNnoFc
OhfJjDvbggkattlEBjkGR2n2UnRO6XQqbWeFVlZuhLOGJWRhKqKV2EAQ8+0xbtYAwoS90jIe/hcz
LnlKA8fCS5Hktwvyil74kbh1U+xVBcw2YCPhAMN8pwrrueCebjEtuPuOZGd44byMWVh0OojrkvP7
z3ae9vI2hAmn5isbJvPdFoitOha5BN0ciPNTdqwAOzN4MRRFHxG9A70V1x+IR4XSnSmIHokMNOy/
kUxhQBf+ya7lFa637fVrTawXAXRrnfaVKO0NhZiPEJhOQZBE8r2zzXRSRT6KcwDp1BNJMHDe1B+q
r6C9VYjs5vkKCv8/jGQ8lGdKVfzVFVX482DLptzCn+TzudlBrC9BB+7D8NdinXX5PGV/gaU/g/Ks
YEThJ401aOUTxwnHc/Yu3l4aCQ4fJq++PXf2taiDP3LJVWUy08/ItdGKskIIx2QmDcYLCIU/DxTD
Nk0o12ysdEwlvtQAl/qWMnQbMh/xUpzYAEb3P8ZDs0cTmgbqwkC9BFwKKMczQ5wkuC6j9URyu/T4
2V0x8Ezyrep3US5yD9R3aWIORRKtW6sh9U5EcsDE99ykcZZyp/O7aJnqAL5VHXsZraOajYPEyWak
E07HwqCo9WrcY9+k2ijjvOiRUZDHdJc3UzOl5gT0oIf7NggQn9qhJhNecEWilLe4LjDEKpbZaeTf
J60WtzU/UntVZIlfJ9q5RDHq1AFCJP6ZnY5ew5FKJyKcplPL3WUBuGOdG8rafZdVUgHJRVnTL1X8
9Jhpir2gcGPaJoAnaKrH7Zb6JHiJv/++/bStD9/wVmzKeOZ3H2pd8hXvTIbMWidNiQ2+zpVKP6wZ
SjwDUA1zfJb8ntHMQBFww4Uro421Crj6jN1+y7AqenSywv35UmMWwhzY9AdmXnV6j0u8p72AkDET
3DtmN4yEbXOhli0L1/jz8h7kzDk1hrqk9n4n+7mjMhWffQ9aYcxIy1PgvbJYNsIuRfGjL6NioseP
6lPXa02pMRK65Jftizh6HUck9OremPZJSCZQEy5VJjES/S0iSirm6gE53itorZPT2xyyb5cVf0NS
x/ch/WhzTX046LNHBDgkrheu7BKWDnNkID7IroKKVl+9BzyBSXW3VEKfIuQkYjyFXYTbbH7hgp17
ap9GRAnYe7v3iJC3yhoIcHD1SPheSwD7u+LuS7Zh8slhhEzlu5Bb68rJqQBe7/GkK3wYhzMzXMBB
1y5uTs52NORAgMg6quPzGTy5em6ZooMoJCbdTq3sWrkNT6l9jUKSOS1PNN2DqLv0zRo0cTivjtZx
Ml/HcCbmm0u3rteeYW+maVM30hSOX58yR11ziUhbewgX6rlRmvHbE1lqqWwHg3zMw3x8R5eQ9faT
2kK5udmJPq0TdDTE5KE+NuSCM1q8h8MLgHxfU8b/IVeLLVShqyhDO2gd6FFdocHKJXmnWkXqOeso
ji/z7pIZcItQV2Ej0xzalZbzrptDxu6c2bEPCEA4Asi46E2vOzs24qn59QbR6hjcuxRLZCR6lsPY
T3K+tyBpFaeD/ORB5C6yrY+eyVsc4J95wMJcYecbcqFAype0B5i2XsQ1jUQR2usLctUaMSun56Pj
VjDPuFH895bAxv78pcIy00k6Fz7NY0HMdTbBaXuUIHdmorCfc1hqfbWErgqRE4pwCTBsdYpAPcs9
hbzBNXhWECKVt5PrST7IhKXjAwGjAcrNNmOf91yzro93ulD17gY1ipQscxOPXakP1sxpXRXO48Nf
089ogSOD5CnoAxqSOvs0ovcBY8/fFS9wEcBT3zB/fFYkr67phURKBw/PbJKycPG+HjT+Kw3jGAZS
ZqNK9GbxpbmJHcG+BP/7JIuvR13eC39FiAzUQ0kw7PSV6T22nEQir9NEjvKOguDudqVvU90T0HeG
KtzSNHwSxlAO5ERNIlebMLMvLU1+6Pr5jyOi1MKE/p9a+tNCCNxA9J9HucYkfnhgLIfdQueXYR/3
VULUzE8N1hvJ3YdRb0K/pbk42VKdELw0WTichLLoFQVn99N+UqSDglkizeVfYr0il+iyO+w3Dg64
wwrj2/rqGAM2sFBAN3KuJZjHUSPQDIuc12lQrQI47ddSBQM3SqZxmhMdEwvVRfoW9nM5hVBZOMPb
XtjaJm2ApY1F1yCZU96F4cf3JKDIm6gXF54dIHadEQc/xCbuUyfJHp30hpylHlmAFPeWMrz8Ohmi
IiTmiUS1ZwDXrhxyw5mn20zXindOaDqbRze2rm6GhghlLJ3Mo/EEYoufQouRwnlsBoLKyStoo48b
aIaYQ8uKiXrcBWsBIxrQWO7gvrl5UF81Z6rU+GcU0F73J8rGjMd4lRy2OkeoeRzJie6A5Kz+4PK5
cm2Ad0IGGIENQkyyigcXFajxp/k54tq+GS9G0z6afyteUKGJ8E9+eYu1m93oouJNGjQDUOnJGDWB
fgaaJANBtWlftvMxNH2eEoFTAMMjA9686dL5UMHs2mNMJjBGo063vBOJ26UDDkEKsFo9u2fFDCBE
zqtWznFKZ9TIVRrTk6beJtDujqCRRa9UuoXm73jUhpYjGs/MsCFpz7fNa3JU09RFeVdBeLkIcFY8
e9dE2BuE/tnuNeR/yjEoMEiW+ooWT9dPNk5izhmycnxN7JQLL3QQNCxEgQp0WZP5IMZwKJfO8Ffd
iEUfdg2xbkmV40ucWztJ6HyezhCvstiZKY/Ica0YM4whPvr0uUodhEQkADsqpI94/gF1wPb1f38p
gb8y/5KAx1cc2Yu2+2hW8WKXTIWSMZd8Irm6iJ1GTuftfOtjZGLi90XB8V2mA7y1YcZDtbGmJ5YB
sxZwlyvHZ8+UlaVnaBGMiF0IIwWA54Me6VfHyUMHH+9J3qAI5XrHECnvmA1XO6xZGvoejbfjMahY
CarKKt/FLoqcw8X80WrgIhv8oDNVyKBxSjQ0qSFmQzIXE9pXeNLLESxH+x2QLH0W/mivDrRJQjun
D1t2GotCTO0ZNEirV5ucm0F3XlFgkzvjJXhr+r/KqZbiB51pl9qEmJY5X9ymFgeuuamcq+XIYHfz
Dpgwz1ycsC3ekd3sjh5m0HL+MLnq2nQ9WifKpIDGiYdW9NGx3x1wa94xNpuTyCKD8JHW7V1Selli
y1mjTIYBMSz33TBIbgpDEuPk0OYWwP2prF/LrhMiwTsz8WBHLwrmB7zqWSkQZyozcJRccovo6ElJ
28dSZyQu5j1J+95pjAndO20pHxQRHB90lPwC7ZZ4EkJN0Gskw+eZOUlWUxh1NKi6L+oMiQya3Twf
0J6VZT4YRhwM3mi+j/o3vLDgWXsay70lMtN18tEs+XrIA2wtwDsuUmzplYqV54M/3FYvnYuqaUzy
V2PAjB9RaVjbMqMYSBdRtHAYBSL2v+HOLBOhh63o3HMupaqKQpXDwvJ8lFeOE7VY7LIJeWEFyL8P
cz26urWF27dYNruz9J9h9Z8JgA/HFrRPig5CubM/HLi8TQQx51Pm9HASaLbPrpKJDK6mtYlQvR9g
/FggoQQzFj35yWTY0nDm4v8zuHqmtJUWqN6e5EVAnctXfA93lf0kY750rsUfp0iuVlgv4PDwkOHv
56HirdoopCzkfOFv26xNf+UVwi83NjuxBTwljgm9QQOBQS9QYC0L3ac0mN19d+atLx2BzHZSaiug
YzdNq+vLfntaNzpughBh+S7qCdpTSk9NlDAfUDG7LbH8ZpkjvQ9qJQ1Iu1WBA1PoFYSseyiQG74J
neS5zdpbsEireAF42FJzNpOl1bK3nSBU3bgbTp8CSWFRAm6q6uWFiPgy6ZxwCrBMQeY4mVWqYWSZ
DqOyAEaOYCTuwlL0/95sZI+jpNxjGmEMWhD4E/e5C8ANMv7nf8BNkterucHsL3BtUbV2lA29jOYl
lehNzJ+EcBcvenDxvClWIJ9hNb+IC+kgLZCbB4Kq0PeNNZCFTK32iXMsaN4VFuKXkhGEEdVpsEpf
XvEwRAvked5Xynblxd7Z0sfwPFpi2DC97RRWTHMcseYtavcvM6duDbq+GGCgf73Lx72mqcZIyrad
T4p0VP+zcMCJRthKM1esJYBP5Oo5U/IyUA+eF8KGOP55EdwFor4rR7800+kbIM1rmabMZb/Brgbv
TzGvqecKEBZOSFbPK4ZptLQV1qMB8S5F6Aya7DwLQauHGkaC5y3S/ZV/MtKCpwefe94kVk0Jtk3g
PFys6a90XyFeduHY6+jUX7h9hzZRk29WenlPs/7VcHX06TE1H348G3swrC0J7eUHxpo4wa+kea1E
3vkLLVlGHigQ1tGHAQhFcF4ISp5kJOg5BMK8CKrjkxVu7ZyoBXhakN9Q7BUuwGKBpbeOXUxgEsUl
ocxDXH0TZfSURlujLAmR2lbCSzxSHnCJC++jP1dPXwo7dshc+Gkz1Kg5ay41g3lnqjERJRTNiU9X
KjivRLY3SNp0Xt/K91QwiBteV38Cv8wJcZRqvRqOMEuH78OKpJA5CFNhBvbtn9jEYIPe8HEHDJvd
c6XtphCtCeWwBOmPUCYxM9n6y+gF/Y8WByLr6zPMQO580TQDmM+WxLgiHJ18Znk4DV4fd+MLMa0c
WykqX+F/C4z5INv0ZujOj8m9d4/OC3Q0i/5iyT8AyNQaX+KFaVZOQg5nlgMoZmN1BnA5lV3j48pD
x8MQjre6ednsBYshQr0ZpF9qZPuvc4F3BZYHf2dtZtoqXCBtOmGptFNJ7phK4Ha0LZrAgmvTy8n/
X5SVZ302cS/IZJZU4d+Deh/3QAGuqi00l3FWwBmnYaI8g/paz9F8jRpaiUdANKx59OfAHQdbkQta
Cdq85kZwKPKhyf61l2TqWnkE/Lf9NC/LZ8WtYwdM+ve/1cTKp29KB1FfKKwSMmWDX8dC0+lHRiBw
Z53uBabUaPedosTZjhyfDpErIDK6A9hDe5jbLzN2EaQ+zCWDFPG55lA22TrahXKcWP5oSOpvopSb
Uz4Zh0DUQVWV0VfIVM3KBKfTMkMJEb61J+9Lix2Uw/TPlQXoUVjYve9Iho6A7Ym4hD32AWFm8YX1
VUWLcOla2KlieQpimOdHIC/qEA25s7ajivkSmbP80AJYyyACvGPMvGpDxADjUzwPp3YGXoe9rMND
Hw7fVHH0aXiaOIGNwAf+gel9kBTREzXrGrLi5geIShGnc9Jya6lhPaiYO70r3YUS6YFqnX/AANGn
nY+OJ87dVYfolWV/o2oLUnhlyconoCDdIsfzvLP7pbVqvXk1L41PDagCfxQBaFhoLG1stKMvDCQU
ybLPkDFpVjaUbQKiVefm38r5Vsu/PvN9H8mX7aWQxB0V0u5Ew++KRkE39h6TfWjufmEt3IUmanwa
S80hqE4tOthuFiyyTNWX05Fo6OhUrsm0KBHqlsMzo0VNHFw9Y+xngzTbFUi/yn6XtBL9TKC1NHVC
cv6gsXJvHV5rbAxrtcyBYLhAiIqosx6IFBpPFsdiQ8Asu4Ae5j2QCx08EX2DINuVJnSM4/P4zg51
Zx7VNNHgBVXfpTFEpjn1DlHhOz3qc96kdRWWMuRqv/4WvVDeueWQNKLKXgnZHQXmKceK4M8EWXE2
dbvRl752ChY2ggeaGnBXMGhtdpV6ZZjjqFdNU03ItqAP5I0fJtIL8lqncpftFPu9XrDixINqZkMq
vbpz2UBH3zRzdQ79V1TGGix0gSWcDZyg0FTxqfEgIxUoM3zt6XXZKsl7V3QsOhoGtVUu7kCiJJje
phmC+B9Ojbe8kBarojQhQ3tz776MI5xZ21RXcnkvm8ns7akDexAtYUDAzcIKP/Cw/23KZ0uJ58+Q
Mks5fNJXo79C8BmiTYRNC/3eKylZyDod06urbVeOyzuRJQVs76a3Dpb6Tdl9IPUPoX5ykxZo88dq
pMgRnp0xzi0LKQ7GGqRbubJqVskb5f5ggiSrsIbbv1AixWUVCQYb+TvfbnmilgfmMgfhihDGjIfu
+h48WUIIsNvgWizjts9G3R2KKdeyBGB4TR0fo4L6RAVtmZcKTiVlwFK4U9bdgQiNaoxtIW09QOOC
rOwZy34SEwHJw8C9Mh47PuL3H+dzPtZxZZcnn+WCT2aoSpFKJy8wBYX/v0efOBYqjvBkiXDtSHZt
/aMfQv8pxeBZHBT9DmfpP/fm+wQjSt4dh9iMjV1QT31kfp9SZwrGWEFxDXiWkXkwm+TrNndRzAFr
3PYzZjYZvfOQpaJ6IIcqKKYbTL4R9GDCy1SJ1pw7t4Yopct3q2dpB3osSis0ZiTw0s0pAPafe9YW
yt3bSRGSJoxUlvYijK1tEZ9n1XEZ+Ne3jk1mCIljoTakdekHJnEiaXK7Dyof3n3WC+qsEM7nUEPc
l+sVhl/DfFDy+95skzGp/4pFYjyIFoq0aV6e+NTwkjZDdwFw//Eka+0WW4WTVqqZcjGcPH5qS5kk
akwLp090lOy2h6ItHUJtdyTxVBeF8VF6CjAI+DE4+DIBAWqfJRmzwYMWuITQrMWcD/cteRDHj2RC
23iA9iYYeE1FmzCmKVtAnpClLeVHU+1eyNM4BfH3B6mtHGPJ9WH/imtPIgXKoRmmzM3RCvAkUGim
50bk4VJ+G8uSPG+f6WBlWW0Bh/jmMDYLE51/XTCjsTJBzCn10FwUQ1/NGXugSkidaEOYEh/B/8fO
8XxJ3s84rpO0oWDQ1X4vY/PTOQnmIademdEp7yPlnigoljhCV8M5v4FdSRAHY5g5cC3UEiIXdy6+
sJ7RjD4WCx3G3a5fuYURn8QnzZ94xDyC5Eh+pdrooHDx4dU75CgcmqhEi0BGX6cbvxUhCw/gUJ5L
NtDA4jisB7d325JXr9DDXdoteyQg+Y35RMbizfg1cMldGCXyuDcvrvc1UqDivBc3bmkAfj3+5qOd
0xSjGMJF5MuUUw1cjVyJ6/F0LgO4fY+pdkZL6KbCpWBr3F7t/oOqjnwnW1VSFvx10DBMulwNXCjR
G2ocDI3RsxYcwSZvuRB8dwLfHOoLTmbKFlf8y4EJJCn952fxlkk3vvfgsuEUJKpiGucxqVngq5Zs
He21gu3IIOaFNRDIOryY/aflxZ/GrlPWdPS9ImRnXV8UCydsshlDn1M8D+IPwEtnxqg5aYXIIQan
g9PP40DI7PFih9nef0SiBO6f/KdIh/9qopJfgZoW8+uexnhWz+FmjC7L3kRHB4I5eMR6kMFla6WE
7CpEILfoHrw38fVsinUq8KoUq6mcnqgDdxuv3rVv/entfyXKAHAJQlqYe7J2zwBz4EdivztlOmf2
ll5BNJoRSW636vYSAOkpegrI6jPNAb3j6QihZe855RZMsNXs9QOkLdwoG4gZP1qegijCppqsrQ3x
ImJGEQGmPnRrFRVpns0M6qlO3gFkwcmW4UZiG/KQTXnA/S8xSG3qEEMt/Fk9oB+K3UESSYWsistf
Mjwm/lgGfPBZ5Cb9gOgC9BZmcU4OXZ+ahH9pGwsAheV+b6JMPsuw2BKe0cXbNaU7d9QkZ9bnnBPm
/fAYyolvWBCjXJ4YzSPRELWi301pfbY0Bge2YfiZOKm/ZbkgKNC3dw1VIchuRyR0TaKjpMekd4P4
vLIDKj6Wwgv38jLDyQpnXyhldI32p8tM68sRRUXAUayTrgj7mHQxkw3mBigPriERg5FKH+EWuUAX
1Xu1ZIb5LyIrrqNBiNT7FkpKy6vxEMJRl/LRcyLw6ql6dxissAAJha3jQU6QD19A06SPE44EzfNC
5+xte3ct+iNqU9KRymzzgBN1vWMXnhof3W6zymnhVVMpbh4aHmLK4VXk75QhzkOFRByVTSZhi9Jo
8ZvOV5eMRXbhwsYY3rDkcwWsaF6y3Wj0iSSxt/JfyZx0YIlK7LjHzW2h3Ik247EsCfBDdrWzxQCH
IW6tmXY/ieSBy9We/zs+B/jEYqducKRyxyrH94ln85rocDSWn3MdHk5rSf9ICSAAxFHd0qD3Itul
kQXZcOJkDmf4jZYUfnoqfAn7+EXUC11zBwE2PsuKdUDu8AqUrT9aQYeuSjU6N4gwJfmqHdU1u4fC
kqgQLpSjtZDhdnKHjWn+SQgKBfFhePu7R++u6mpBk6/Q6qpmF1KvBdpJDJ9hILmdDLPqEncFVv09
+EuG4zI5NPopJ1tHaS4GtbN9Bx59Yhs7aAVHE27g+WOwa38cGobqcDY4Fb+juy3jwRu+e9OEJJ6F
ibRPHaYm5khZRFPVzqAjrvgsSGS6jbn83H8cUwD0o2rPKmNnBD+58DfpVq+JPqyQ0QdEoahsZZCh
9sSb/CwQvksIsYn00SrWy2aVQUJLkF3AhlreqN88/+j8R7Kl5oVjuhXREkMzk8u9xaLOsQXDhtU5
VVlJlD5W09KM1XLU7gAsteYD4H0xPQGYO/250Mm/LRtYK0MDie+njMR+O5sN/e8LCrhZ34goqP/u
6fZVBgGZZ9Qd9mDYpNtQQrbtr0Qa0pweMul8klsn3zd9u57kj/DDjwBCSLuRRQtrtVEdiIF0rM43
yBfKdd87ikvKAaR0UwnXtRG/XCfBpX1fmotAenkFIii4tXElbpS2z5SDLDVg8sW8647Q9fSB7Nqw
V/bccZGlRKTkEqEzd16tCDQDpkCexF2i8bc4k/gi0/EXjYigrBNKbDOrYxtydJl/A+uy2vdxyEO1
qKSDP1M4F5BUYBQqxZqavfNk6mioVT2574lKNVd+E/D5h3rfg4uJEobYyuqCK06GxSwutcDw6X3g
N5P+YZvk4p+jz8GFgEgos8UN/lR8Oj57agNEPg3JIIgoz9+HOm3Htukv4/g94Kzdw7SVmV//WtfB
BNW1j7aLTvtl5Hyzll7WqTlekd+eIMza8MeOguFs5+EqknsTjcF+CBoJhDjB2TDG5impvo9zgbXi
JdZSk4yjNm6AHsCGrbR+GhWDeHX4AoglTVmZrJ4RnWRc47RHJUfP4wQdDkL1r0vI6P5xB8O36Ejw
gAPA2bYSLjy2Xogk2CCmYK5pTCmpUndCNpvYFynD3di00JdQp4UChK58CSpg419jx9St/lAM2Q/+
HMO8IPxHBsD3hGq4zh0Pz1yKl0/LIhQiG/8FuCyPrRtu5MnHaWym0+hlMJXWOIluHr65soIfFh0e
00hyHz+Y2nOLgKzBpSLSXl8gVNQi1xAewa8bAkIwCAuZ/hLX2oVDCVEKjycYTpCJ3E937qhK7Auq
8ksq0nuxALODc9tDQ6FoDVoMzpaAqoqB6DSNn/XuxhOZypM23OrpVc6Bj3hruvMPzi3KT9W8h+/F
sur2hat5WL24ac29azwdGLj8PX7rFEMzqNq1nfmcDUQnDgppX+ZyzXXbFCEnczc08anvWX6NQtL0
Bojlb7Wd72G7PCyzPyBivuSv8nFKZMW/+LGzlq18tC4M138eDMzQPLD6LhOdb3aFbdxFEAgjjFQz
uUPozn2GrjSfomvpNcHABqgE5JiYi31muSno3AqYV+LV8UQER124gdlu9KvGxqTpVm60Zqdc/ubR
uyNImoUHuf/p+wHQnmPUKkBMka5Ie4gColZ5HqDjgeVDZZw7EuDQRsG7s80I8xe97CG1vzMzBPFL
6NCnlV38UgHU0DXdKuOrVS6AG3fD7ztB7Zememar2qK7BPOXRLKlLHy5b3Swa47uQcv3KQiQj+vX
iXUdVmTiYzESIAEBcmY3Eyo6scKjnoyLcHdmsDamsOAmmMS+KfD3HBtWcJjzNW+3WD90t7+3lEUw
A1Iw2tYtQgPyyvOUGkDc1ALjc4Ghg+ZPP6AKaIHovNfv2mCaWqd920O5x44Z+yvpz/c8dKV9mHsd
l6ERh7FT7gL55hO2bYsMaIokL9d3u9Fk3qRrIpCs0wc/G1L0F6TA+S2dQESCvwRd/qdTe87zY5Y+
juLTV8vTwi9nnaHSunHBg8P6FAnMLYYj4bZ1Mzg/6Kl95YzKMHgkqCwlxF+GgQ5bpnJ0Rp76WC4c
NuLqmD2B/eQfEkNcqUxUEtKeDKgBcce6er2uAa/n3w557fvrSsLHm9gS1lXiEkWYRqKdRUz9lgdZ
+7DxuQ+xaS/5MSQz1jbnE7Ij1zBAZhms5Y47drh3uCBG5V2bhyINxvW/+FfSgx3AgslGNGncmeG8
xj0LCHIMoigp7lxkDzdJ3KRNEAornBmnwUrSf3Kb+H7yF3ZbSMna3XAta9ZWHKt2h4vzDT8440m2
LL5R9BE1ulAHNHlZFjqInMRRbXTk6fF1gbHuwkuUm+zUYw3rn/ETxkCD0l6Tc9Nkbh5/62yS8scN
Prk/lrKJU1BtuHOAxYDpLN/yXCmVZ3GUqfKQv3TsiMdDM1+XCdrZMrLT83LQzLiAX2QS/jqR9ZNB
T1aYTXiyVtcsJVwnz0Q3/xk6og9nBdiRvR5A9emoC2rvaTMrqqJC36SHxiBZBZA9moJg19uiTSmH
xm6golNXHjDIoMp8mDEexxmE+qIEJTLNo7icssAcH3dOKj8CwPcoEo/K2d622dXyN5hNJze/DAfv
8dp+33Y7qJOtFzMtCWbU1WN6FeAGu3K8fyw9Yn1XWMP/GHYLXW+u3dbOMol4BOWWTWqwQ98g5FnR
dFkY5vYp+qLGatzY6dWytc8hoCfhO5rAr8Bx5TKwhKlTvUy9pRHbWcYWAqK7KRFyd8HxJ3cwdA0G
ifhZq42B2IqLED8hTyhGZKJkmCmTZuWjmtJUl6T1tV42x5OE+tWrqeFeDjgtLbbnUmCng5SXDYn8
ihWqJKcXmAmlPvfBV49bE1omsta5ysNmoIy1WPv9Okh0ThH5/r/Tg7yzcsM+rQIPnwYaYZ+0tN9I
5Qe0gG/mzM6D398SlkMJVkdtU0UxfxQ943nbm8DVHQ2n/Q/S47hPWlvqpx8HZca2ksv24Ud52mAB
T54wRJdQA2cqq8XdTCEAkFqyJpoHg/KrOs/A2dGo3yD2Ae8+fXRSErBBl8LbKDCgkrd9I8fyf5VX
XiaOCmEKneKYGJAIKZ2VDmg4oPhN8L/hWrqgYdYu7Qu2/kk5Q/RhNRMY0uxX03TdATdEYvr9+S+u
8lGOXlBztMg4ptrAjWe+5Lyx8h6Qpv2py2AQgrTDOq389+YrVakY5Hn2XHW5KB0zwLciMEP8aho+
TF1uVCp5ZtS6Y5bEWKeAaQvCEyLJmxg02kQrvouPnvUTk3+Yl0508VxZA3qTnAAF3sIgAZOeFDUd
bOcFchXZ/G13oQIl9EMvOb08RP6MAxGpzt5dr+PDl15l7ba1KS82uuVJpz9XgEKQbue8/dn9coPr
269/dtSLkiQca5q1VeqCkc93P+Wo7wZkN9nhG5bBTz+/fOsQiCoZb4g648Qt5gry1Y7nnRmsUubs
3SwCsEa+6mA/pHgXb2lAUP1eo27PzV5+UxqbqvTVzQA9vHI5VLCT61/hM54QFJtZjBQ+FCF5fftU
YdcVmjHgh49tF4SRkYUYyioFI27BBNvyG3Ul58KdwfDWYQBjYLajbBSD/DWXe7sMBF+r8ovOUFo6
RxzY/3mw8XOY7Mb5JrcfWpyRKia4im+8H4xvmC3ZCvduws3c5+hOKrDPkoNWqdrhj6bDvxXnb260
lBhyHj4RMITVn2ULa6OIObH1VmWYY5mEJi/8VlYgnC74QiCGA1JQk4+jgdnz1zZQKXOhTAEpGeWt
3YHKLrIolf7N19Mm1b+4/XZVS4l5+NxXE/KBbQ6BRsjTZnGzEp4ybVQuQhSbjEGSDPS8+2uWzNqC
FpusoaehAWyrprritLJAMJQBM1hq//8v5qcmY2jAY7BDHpzSWraIcLwNqdsGBRdGhPTRnFrBx7Sx
RVOquURheSXjREKtTPcRaMMktchHSUuHRcaq/h9P/hfyVHSSNGUj6zTAuGiYP833Ldh+f20iKhHH
idacy663AGjP9dv1fmAAtE3SpJSs98r3VrTvRg9dNK5EHwZCvSPNu+BS5Zn495Ex3DTDS5ooFGPU
qGPXX2aOnoD990LYgy0cNoA3OW49q65bAerRCcMLaTMiu9iG03e9PCGAOEF8h7QI/b8ixKrHzjYQ
t9OoI9XNAfkYK/ALqTjx0bB13xPMJsYYELCeD8TXCPLnGEhf402vCcSjjEfZyjL4qG/ai3I1zQjZ
Q9g97eFxCsAIcRIQG7fONeXLuUD95H/Do8+vilOIe+RVA8b2EsCR5ujE+MJWhMEmBfMYOvNyUjxH
n+/8n6WHlmkpZm+8MjvVgnDDJy4PYtTcLK2kncrwtWy8vdEMWWI4xAobRcuBYTkLXpJtwI3C1h3P
PzEzLcbiI9zr8KXTeuyi6Po/7LDotx6fdlEM+xdZin6rmv8kPo4OvC27i0mMBGA+CKXNhN1q0ujN
FpreKGrGveqPfDkgyEi6XtsliNPVgcF5/9rvj37GjblhU9YjcaS688CU7yZ5PrfcwTyyeBje1v9e
WPGIF5ZKnP/1k+QIdG4E+CmjYK8tZN7m5nbpZKO3wS1utKOmFYs1HANinTLKORqlapnDYkJiH10s
3Suw9+Eqa/+NkpzTTYNj4YzCldTjERWzq+YQd4LrkRUeG1i4f/pvbPeizzgyRnQcbVFln9Vp82pm
MBV7xw/5XPYN3G7mUCR0Pz2djzY/IYKkovt/6Mf+mPstO2qPQ7BKi9ilrtm+/roXrbnqgwJDuYQC
FczkZh003zGpDcMGicrDTpBQD8bygt7zUJ1gCXjgOEGW9MzLckPuy+WiIgtjIgUFWPZCsGQsfp5t
2LiiyJ8JIOw5mM+JeT/YS2EbypOhPEtO0j3lPpIB6MsXDNUsaV+orMXL9UGNCoACJ8NovhGdf2yO
ZQHa3C0ZVy5TbYIykhzHgQobSDlx4wN1FrYKHw0S2vBoe3X/5/frCQFenyD2wXnYhe9DvwP57a5y
F9vFbNnWUaOLjxOAZRw44BRlNStfeDaLO2I0jAt1JVFIK9k3q9z1LuyHTjeSDjJUAI13RLPBePE5
B+yypPVuWQkTYa8PdkKmwjkKNYBLReIo/ZfhEhWpqRwFxkW1bs54luhapBVNQ38gRKpKr0H7oc9w
aWB0g7ZKn5RngoVEMD+G2EXhOYjEEADqV5V93gPF7c6bZBNA0XYLSi5DhiKnlN0Tavcrl42Lq+KM
p23qOHNzmWlHatAiECmnztIstilEZiMHP0SDvDUi87CJZnqN68DdWm6mfVEmjrsv+LWGcp+F1a/3
kQ4Y5XnEYnwq0vsq9yIi7Xe2fJcg+aUwyjNx1pBofW4E8w6w4+l6zVHtYi6/Vs7K05Rv2snxFA3n
4KAA14PS8z6rIToinvzwNM1EqJTxNgvrR0YEPPHM4PgDTnBlKUtT773pIyFXmfuX2Q44Z28HhltH
iZ48ZzGlTtP+ShQLiuT3bFajtXHAHt2XlmQi9mgbFYm3CxWX4DsMyatmVvOFN2sVGTUH9WgvpQrB
XbPTS+tNKuXWM/MiS642NRXEhTygpowH37BiEh5/60AP4B05D6G3Vl8Xo1ai+KV+lrUfsSKEI9PQ
sI6seShoXX/HjDSKT25qH/QqX8sZLvIy/CNkQ7Bix2I6oroDTOfm3QCm1aReiKP3OU/cY66ATC2d
ddBTwqTbztFtmH+WM/2Pb4iVHOJ45OIMcHJcZAR/LquUMZdEWtpqstu4tMM/R8AP054+FfAx0O6M
dohlG5Y4oBosuqK7Nn6euLf9hja8lA9bRJFlvBZNi5mcv+mVjJA+7TqveeOZNgy77mzj3+QRLPOx
ff98NM0Ywt9k6zTo/btovtQFXdps3pqr3KiWScF8JNQfzPloF/TS797aqe3cMFrEn0NCkZnZ+R7y
bT2Q/GE2Wwo7VWAASTdlOPKFlw3tnx8RRRddPmwVOcEUvXOJzD9Ociy+mcyrufxTyoL7X9UON8cA
t+fKZT8J3wExkBQVNcsm/CqXZxr3zPboDwtcyewzH/rA7CxawtMILO2Vb8nAf8sAd5aRCUmNwCX+
kQK2hbLHRli7PeDVETekNUpkgrVufifwXOuzoQ715OJksiY8gcOPanHWBBQ8ucBB/LD8vW12Fo+w
BxvL+kY3XPy/8F6jN1m9uYJzONFkR0wC0fa5C5nNcKSA2prDXvLZz1RBguKGBoqBs7W+dYOEk27t
4AAlfB5GnofAnmvgCrklE3OznwIkLJ+kjNdlhuHDZOapi36eyvGPETpDJIeGxvKdJB2Kf/uKt3at
kRr7mfnJv4Gy9BaBVUUs9Np0nxc8m8rySK3OKvabxQkOXf41Sb+6lbkcoftcLVykJeBQjgaiiAvD
pjkGv0VWDwyabY0/J9+yDMP81no2PQL9wbrKR5CxFNZjukHmSPUWrPt+VuAocleIaLMc/nYFrtWX
33hPEgcMhX+cCKG+Ar0yUg9kz9BF1TFaCtVIq0f/u3S9gtHStuHus2TWrzeLyEgjCxPCIaUFie6h
3ErBjhEva62kb2OIMHB6xVzgDmsVmdxE8izgT1UyHr+jb+gzU+IQ/wsDXPnJ+/vksZAuQUgMfuyH
IfNr/CX/YIVSFoyPfCZ+yhJgB3VwF1u6AnAJhkLnZnZ7BK0S7DWd8O8xpvy1NwOaRptEloQz/zey
WKfGOMkkJ4E6XhcyDg6ExLTqhJRtKNMM/Z7M2JfkBAiAFcyURJiNLeedSsblSExoyMfyR6rDD3T9
wepAPmAXxeZUQZtwniSdMHZLRzUxyjARABe7vWCr2Pza5ucWPCZbPUy0jRvV3hGAkNcCuTOP3j52
6SP1ttbkMuLu868xpeK637NN7pFBkeWCypKEuIkzBXO8TuKZk5O7t4jZRsxkQ6BqQR8c5z8WCC/6
xVt0Vy4AO6XA1j6pjPJPvDL97qZJg+t1LbJoOAjB4GTmw2Yf8Vdp9rlNz9LY8fM/S09gQ1yXWOuf
b1qcUVpKCBmIlSQ8SfMAJr4P1mLzaaI1F45ibXA7udPIoR+veGryUMbqOQ1PU2skzcYIkn6ttHrp
ADQA+lT/Vree1i+D51RfojwVYIeJsAozX2ewx0lWMMnAYzi8/VVsDQ47iJasas3MuWQhrQM/9ihk
0py/8eiP2hsGydJJi0fZRfrcABUSgjUPM1f6CKWcvwevFVKW+ZQdjxYbk3bCHRulEsS+aWEnTG0C
hz+FjSQPZKAP25P8OHogaQjE7NTOWviZBvMaR5hBMBxDV61/NsQuWzsSv7QVrWmkhribXqnBAMMf
0ybP1OTrrOpbifA7ek9iTbArQZFT7O3gIXENVi/MsgkfI3oc5hsxq9oP36SLdGvfamLfmTRXy3jb
7SJQeTcQbdW6N1S8vm5jPN4dMx/pWNNAtFeDTKXHcU7R9t/4QQrme00ynIlS3nYl2eav2Js+DfMC
mv8FtRYKlCS7cc6U13tKaeANOXTmaiBDvNN3dkN3R9dAI0mSScQfHMnQj0yiP7NGOvGlQQj2tZ1Y
NK5sboWcYsTVFFQle/tIJwOAUZAOV7RotOsvyPJVLJT4PnNJqj+sLCEa63O/1E57ZPk/aevPY1KS
kfFSsfbON+MVFuHUq1XB9Tx9/suPMia2K4uZaRfvb/03g+TuAbERbQ4eG9XPcLkEMBeFVnS92rLq
4KyMt/UMnT0IwS3S75WLRaiCJpaOl9r7ZbL3smW+fc0n9i0cgwh7UAnNAkuPp6Ji/q0LbhpL5E3R
VjzubeJR+WeM71T6qC+cWDgD8dL4fv/JBroOil4vMHB9ZBOzboJkIf7ViqxlblR0dYmrhIkzHESv
fli2E9TwsLzGC/GEMrpWyMKLXJCfQgmC50d3XgGfgpsYzE00UDPfSdFmrS5vM+D3zHxueYup3jMK
WwYnZnVUSSAZ9J7Yh0FwYIBBbH19Sy57T7ObMqc5Ow+4fpoJr6dJXBt2MiVkfh88TQ5a5WGa+W5w
bPq43iXKoqHln0TFKyietq/bSz+aLRKgNVg3lceXz5KhxG9feXQfnNaKFrq8Cqvi5nLOqXIEMoj/
MC8o15ABQjxS4Wzk4SrYCyV1SHLYmPcven1PqVtC36yRCXtD6B4GGDyqde7jBCFTb7MipJZu15cL
qSjaKuZPrKhgt4Bly1rN4Lo/7EhJL0x0WnHPbIR2/oZbkJbjJAV1lUK+zTV9jOf6TYKnEBwdZM+R
+d7Ioyk4Cyx0v/AEoGDXOhCcThXx9blgatUGWPgjl8bAfsh2rp7mLLYbbWC1vz/ip75FQe0R/Y+o
U1k4/n4Zi82XDh7pMzdYdwdmVFOqNx+EPQH0g93nkeJayZ37Ut66TMj6D7V80tK+O4pnn8vF4YRO
fXCenIeYvE1cSRK7lPtl0Y5hzyDbVFezGpXKpveYazdTqrAkutBfDYTD5BL3lynWkAsRfDzmdiq7
8aRWlzCC1wcTg4GXz8Loqj/g3J407aPKF2CDESH6tTz1MkgAWXGj/9SkIIOIssWCTyP+Z4S9MnpQ
/8QDr93mCzWFRrySS6WNOq/xyZoXa59KYQQiILVWygmyMwSuXyOxH9D/gnVK0viwBZSd56j3/kvI
/46QkhT0WB4GmrGU9NZoyoye/CUVcpcFH4w3Ge9a1s+Gm3KCa3B0AKqNGwBe8KzeZvakC1O+u4zs
D5vum6enMViwG53BKP9+wudFNHYA+31lO2VWrhRuKZzS6409SRnWYAdDsM3DcH/CBQRpBMtc11Et
8KC9yaus48fxAdUKftmGg1X90E57eyNZMw1888ct7Si7pHMF74MTOP4mWbDscUOUEu9i44v43P/d
FTJbC8NmWhTviqJhjwMpfDUvSChPbsCbPAptDKHWApvzlUr6Jg1vEDINDsccvxYmS66Prn/T8OFw
Xu1rahO7z1iJIGtwhVKIc1sfvsSY8XkaejP+vAMyRPT1pO6fyKiDH9cMsNw+C0O2ANpeLHUCNyEX
eptzCO9Ir9dr04p/DpATgY4+xYjvd8S/hQWHtYA6I8EYK60x4Ve3rv5Sg8VoJ9ELEPaVr0F0L9Dj
wnksQdplPSd1s4xR2xbgChnZYWK4/UM9NhqVPxPaJK7H9pmMIEXFmiPtuYPklOqoGIpvFzOQaH7b
QTSwsJ+BH3Z6snaniRG3Fcl95ook67pPMU1FBOX7DEn+k/6D8pQuz7yNHCoU4H7BF3Ri8W/gaUBh
ddP/0AbGqQqLo/ogE9nyxdeY84bqUfJvTPvBCyqPd8KUskh4Zc76CUqtzXq6Z82oiYA19I+7qj2I
HgNW+CTR3HWdfi3Bb3A7E8rQRkr2Ir93xpQy2fDjJXReBWnndUSWdZwDrICvvp/XF5ANtXL+McUm
2nH+iEhaxj1jBZCpy64gctkZ4By/b8TyDGTdXDud2i9lTV+b+3lNpr5A6FWLezOhqp4WkPFaMeCz
pp71jsjbbFjys6F4BybNW3Nj/4db5ZDMolvSdqoRqEu6ISTBRh5gdo3LYvrVenJQKmyc7WoPBAOz
46kY8YVSdxMaJAxiWgMdvs5QMV9/drpPHfVhMmc5weuiYqNhQVMuw+uPqTno5D2sre+S5tOkg7xs
9PgSzFBmZDaH+27sAPj+6YSSKR62DNKEs1sntdKkm1PqhVpKbSmFoq5ypdobbujz5PkzkKzw+cYh
HYjnyvXUA0fjgcW6QnRy1pVJuGpsxkJOuDvXVqE4YNA5botMvnlkj8RIkYUPHYOnkbn1QVnUQCGf
+uIoSv50btmLMzSTDEka5Ne7C0D96UnqEv4TFf0DzEQQKjz24fzVP9GAEahJaIi120zVA8eM7UBk
nZTIbm0LtQscmY8Gc5g4xnn87DCyKY9RRD2NdDnUCnJ+CJ1lMfUvEsymD4YWzC3yVwjFddAgYPXJ
/1mrMKWNsc26ZqBzLyk6yMQ3lbF/UlyCfcg1NqTtYQC3oGHvOkaZ/2Tatt0bb8fCYP8HYYa8toPe
YaN8pP4in7DKey1D/dIKosbRnoeNdi0Q+iWYY35AxcithSevAtzrPl+YYhSMyhVOq9chAUpPTgvP
vp2Vrfld1fhD886tdeBO/aZPo8VCJmXrO66F4GpUhT2+8BADEUHid2kde063d+g30msV5diCLb+z
FkpDV1skxZDpH3xzgKTs0I+eTP3wVbUmupYnFS8BBab46MmU5AktI8dd6WUhh4JlYwQ2xpRu2s/l
NzvWh5FcGvypGUuty9MkLRNBjhvNlVfYxlS75pMrWRkrZydm7QiObAB8ZT/DVFSOVwvmPxiiMhS3
xgXLoIcdDG6O0FzcVmgweoa5TMn/3Ojo8TBJ5ggBg3jsMfyrnsir0uGy2EpC0tsncEAHNyFcYLnp
10QfGKFHbYd6kU+w1TXHc2UywmWN2n4keFTxXNUiQOZGLYhzUBnQczILtezkcT52AaWaz0YH+0k1
jzZweDxDp8L0eG1Or3b1ce+wYW2zCwVgqyvKgAq8/rkSJkz0OfJhSIePt5R54yx3t8ca6Kdv4mQc
UAmaVsF01a6y/JDVTCteHJSfAj9mlxis/3DOk5T7x+K9CZHkduQjwf5FqgxHjkcR6c1DLb4obRrG
K+qQMqsREgOGjJlYMuGqj5lMx8BBP9R2jxAkUUV8BNTPc2gpb2ovrGN6sLxhLYxxDI+vOdPviF3F
3iYJ/OGmcMfrTgfMTw40Gsa6FVxwp/9wiZTXoS8KT/dbjrkr4XemtVDNwlK27gbhpLw0Sg7fvAG2
JPNMxkVQB9yZRDedakKEJvR0QnWAWhX7T5pp2acQ+IGHAw3NBydplCUOqT3/+HmqB/Tz2Py0SdYK
aNB3WQ1whMGP5HZuS60/JtSmr1EmVoDPEJK8rtEP3c9BUEy+c3+dObSJhZBUI64cvHpNThrDiNaj
5n7rYlbzlRQ9sgFE+xJybg0wR2aQLzaLYcJKtFa0MThkkfZHdAv3mPO66nwz5cMv5E9PrB477CQG
5n8atFbgxBDsUtcPEf7qPGijlifIS+aD6sBYIUcWhsBrxQQUMvkvbhClxk/MPnr18Wfy7wdvob2q
CIZSsoLQfqKg9LgbPv3pNYJSnd/xNG4PF9E0iPb0hg8Cceftopp2vWsQgUxWS53211tUdfvtddUG
n8J1+kYsQU6fVgELFA4Umgn+Ftzdb1PfcFjbMYFf8CV7cktqWZbp9A3QYAhjav91GBzJWkXBDBke
L90qCcwDVC2qmGpgyPLp1/YW3xEXMlCl1+GA5alDCxCv2SFYWW0eWGVRgg4OtsksCkdfqIs5T0AJ
Yo2r+bjVJ4xO00TwubhdHTGmhwLzmNxyQUdLjbk5agANgk56h1hGwDypHz+fuw5v/Q6uRRhwTYmw
tZErys6bXuSuMAJB+XzSfRcCK88KQYeZnE7mL7k5/81PccLwfscM6iDO8rUEd0hqISk9qKW8E3D3
cHSrVXNWt0DnI3kdu/wkN2KnwY2Rh8Kmob7wUt4YXnd2t87VcR9RuTRd7GjRPXwMIOhYk5E531Fw
Z0E3d8Qawlhm2hs1MUHbuVuWGwNMxsmIVRnk09UWSVeT9jXE57Grkq23pbLBBCYWyOn+920EEIAT
m3xZxye0BIE2tAS1P44RToZmAjtba4crePtqTghbr/5N/h9g2jNGUlS1Ax9HLPddRowK12xF+QOd
k2BUDxQduqCfImJqE625dRbSvdu70vNNslsGkO5XScHTUXUSZ3V6opWjDiWOp06qxwaxyrt8ab9B
ZbyOGyR1AnnPF6dO+YFK3+jhTBTx8AUuFwcK8Bs4cRg5yzmtTrmrK69gsArvEcU2T1h4XuIR6tpM
eLgXrzqbaa0PNSGs2fuHcyP4oTClafVDOc6c/2Z81Fg6aSVFabcFhPH8UxLevprAOv6v9zvF1hQQ
Gj8AR37bKVGiIr7Rs2KDZho1vbLGYATKY9qeNl4oITohaSTmvURLfKm+wVMmilq+EbHS1hPlYKQ4
nYmtkkFR8D08nYCs7Vj9iAhCO6ir3lseK+dwJk5+Zg8UkbIp0VZIAcCNwWCnIhad6ZwXCHjmiFin
3+u38RfABcANdpVYGMOrOmQr83N6/cMRdw8reozacLk2Ym/cSFuZ69n2RNFWI8ajq32oX/fkg9Xv
iestsea294XKZjiwwaUnwj4UuZzQdZ3phAxiw/UVh+LK5fDPfw2zeH8rlb5FflQYRjn9YJvIQ+84
Gsu5+X+2oJVjygThEXJK1UJlXTui1IxuK+mkN1sV0CXlqVx3kD/TFrGihJN0+pld1JoO4izRu3ZT
foPTlVlcz59b0QPo13wo3jvXv2h5qCtAu+w0OQophIHGcBJiKmksWl9u7aRipC+fThYf6ZXCheZ1
zSIQELy+vXq/FhrWQZSjXzwr0zmvVH6P6fw5nNEiTTdzmfvAMHFGDZJAFdAhX13qUgO7NeuezTxO
F3kSFlcOaOsvJoSHIQPqRpYST+2/Ul3ELomO0Bx8K8igDdHrh8DB+0PI9KPwRhTKVnDg/S9aGmC8
7rqOP6UZTQFRF2Pz6z+QCRkBpdfdUkE1Su3F5yPA7cW8phS+cWPkn4TsomIdpCBc0pdGgasvIT8M
bMSF2Iwl5smwtv0AkkzlI7Q1ZOnKK0SXmT/24tKRVm3Bj7RFm0+7+4QrkSW1XScc62U9mFNL8Ssu
UimEPy9gwZPQYDzh3s1qFzWVkKjrfMSYjs4XLlwsmalW0+UDRKASjohHFnmg/w+dMDH3/+Xp67fL
evl+kReMLtDv5xh80V27QfGusi+q6HUYdwG5OramZIKPKiRoOYDYewL191FP88ZHv0Bp13+EB6p4
jRgHWPoFpmqaPdg62R7vimEumA2jZ0VKaMLPej1O32z85WGYCEFhC2JJfLuoXPltzhaQEAZYc6kg
oTk5QHou7Gu/5+scmCC442SW91PxVHCbIjj0xA59l6ztQPJJ+hiyNuGFwfQh
`protect end_protected

