

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QA13xX+R/ACi8km79qumYiCoL95/JTNXmw/Mv/Sollu1nSewLnwk6qQvytLuy2zqP8g5ZHUfDkXy
dYJVTyRzKA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nii8tC6PWRY1wcl+Yj+dJQmorGaa82N6txtyUcQdtmyxn18ohe6n/SpcWdMXBCN1HiV+XVlZhDEw
KvXEmx5H6nBr5/f6eVRIc3k7vZjXpluRFM7lDsLgIpfE0fW00UnX/0rMYgmxn+5+4dG7smGpX72S
zm4Z5q7tYiBa+z76ex0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
yppU6wpcO6vEUEaOZTTT6jS7XbaY+e5Jeh6nknICBRlkmT5DzQmd7eWK0ShMWSlNt0Fv0kuxSdt3
PRQVKoJayZoHlh1UH0U//6ySDV8PrR8ZKYbnb5G7lC3+6hAsVS0WEHoXFsxe3QTXWezPX8OXISSE
YYTVzXqeBUtBDqueK1cvQyMM7IWnXgyQ/0dRh7UmnEpiOonlQALl1eEnWSxVZ0L5cd+jDbcSlWqj
VgoBh9A+IbjGjOjE8FOaFLUMzvKXmpjNiGzhwyN1qXczrRlE54AWkRUECVVEGR4zuEA7VTQH6H/B
e1HQhNsFNtK03nDJRyhoiacaeHGOBo4yneyZRQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xoEHrB3Q0Yfcf3MYYTBHkrbmS0WN00JVFDeAhGuvxPP5kv5812Q+oIM0e+z8RwGLEwQ4F0j3UPw9
LR04YDkbyd4XfjRJQED6GhUyhlVHkeZ0vYn6D/hB6y5zA45LPFz5aqbLudigfR6lDZgyof50XSaT
wkqaJ1dNbsbYXDGYiiI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SZoZou8zrLQYkyuoYxGz7q7TKCLXDf41gJHR/eNOYbjhVAUcJLojwHpmGq29Knnj056DtiEpAnUR
HkNwqIIUQ/PzBp2ZRgLcYUhgAGFauW9u5fA3Qe79SJmVAKU55R6eP+5h6YaMx1oo7Myp8ZHgv9LK
0atkww+rNUFhc/kS4ivaypKADJgY/Slv1X55We59ldg5OMI3+jFcKD4Ow4Gbs5tHnIUzKQ507yjR
1wg0oIoTMEm7GhN3wZnee1A7XeomsW7IrTE+3/M1cRWhdrj0rq5nqrI9yilbmzqQyqntfJK6N8Y0
QQNZFJ8oCjr3X+2kFBb+Pd3/scpZe1PtOU8TgQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20896)
`protect data_block
kVOlkw08YLkaFfn68kQrFCUDcgHAXpllfS5emIW++SPvNwi1+/9HeJbBH2toJxSoT+TgsSBHhmbD
2k1xA+rrT5L0kJXAdGtBLcQmXP5DX9P2jSYFytbjZNAaBxziIWZ9p5c45tR4rsBeCihWxXqxknOs
CEdOeYqJHa1U/lGCLblsc5ALxarF/fd2et3BJEkFgGEr4JwZXK2QcCMDQ8gl+80mPJULe8CVFXNB
ng5Zp6nEtuVqswEoxghLZAurftCtJhTpVEXSINZYS20xy0mnwVTKNQXWqPhiEEmxoPu/3BLCe6qo
7S79hYq9BP2CKIhjS4m4eyJtcFENfu4EC+sna3B8OwrmqYPSS15oSh15lPJTWEVBdpZ5StewxpgN
Qrb6ZLsGiEjFtAy61TSixQ+EtOOaCOunqUw1UwWMzoBb5QK02mnxhlFe07MywvvuQ5tVuyQEDBUR
Uc5btYIoRcgE39Wo8BiQbl7z/quRQBXUxlTl9VOJN2pD5VBTQJQVjLEq1l/ItdLtoFbPygMtTABh
uH36r++OsDLA+tqlZ4yBaOL0gji1oDKFiCaozCdIsJN5GmZBMGTFNOmq7SEeyIr3f62CzCfdBNyg
/j4cIpx0yRipm9cIliaXVf1VaTf8HPmxQR1xxO2uYH1xGAg/Ru4lLfq54SpQ7oC/XZQUS77ZqLOH
NeT3CGeVbRiS3/ukMTvOnmf3LW52vwA5Tl1Sp3yCAzziyt1w8MlUIitduVtax+ZqrxRzcnpiE0PY
bHJIKaOTQE4QBsKEcFI5KIxixZj/Aq/niYhZhG+5Jsd5aC2vk4psygN+vyfCQBpcHnHaEWyuAIlL
oQSmtdZ8rkUaNx+Vs/i88C7emuU7Sty5z1Kr0fOaEusr8FlA1w9qnSxJRV+pBllMT3BECWoqU8cr
gkABNVhZM6NqliX00Gl5LjvPOi7p7PL0qBXv0f8uXWQoltioOIub2OjQjH9EOZypPK+wc/FXSp1p
aNYBGSDErOeRZllWDj/ROwG7YQUPMyktqFbvwObCrPsWrkcpE6GvjsUagqoLfCpS/0+GzURx2GUF
RM9YAbpcg5joJsKmvbXS+vrqIOXkq3TI02qCa6U5mNkyJiBv3YNOfq3XliruImc5hnRaN7L9WG05
44DWsXgNpfrzbK+NqA82tm4sJA3p1A657FqssuXNpBKXlg09GMq/Sgd0laXG0UXPNzWjVkFYIM2X
ujK3siW0MEEXxDeFc/y54kWC6SjEeW5v1Fw9yXrP+2+nzDq4IFTT/TB3Sl2ZBePufaB8erMtnpR4
rOfAQUijX8E4xbGs1D1mvb4eoIHdA23ygVZEqBCpg/I3PaOs+6QjVox4WYs0GQVPhbmhNP4W9woS
RcWtXLgGTRvxRyQh6m84LhSzkzMHN40S9MUWerXpw6uqanEj44n5h9n/i9WtQXs2OqsJ9gHuYcsv
vLoi3hYzDvqF/puka5MODmpkYkCEs1jjTQ/MDFRWUzom/FEwV2Ni4ceJ1TNWUBzNUadXFIMPJF4S
/TfIQcgzfOSIj6I+EeFPxtPfftrlj9nBakpyXPQgnUHoGuOJKtc+o48Lje+Wxw6yPZmJchWQfueA
95/OslA+nMwfLS9YcP9BApt0fq4vm7U/8B3+/tUs7GKYrT4xniUtYiIATze2Lr4SxuwhfNbWG70Y
i8NqVuGNyp7Cx8l301AyF2VSPxIT8jNo6XKvV8p/CgmgQs0Vbg7Id4lmIv1jpbiSYJWoeP4V3C3f
wDTPOpQrM8rNHkcEUESrl+GQMZ4AOXY/cL5/vaa5DvX1OLAjxXLl7d1e16tmGcdPVeMaTK+o1uQZ
79Pmnboa90VmK2pVK45dMQ8LX1M5rql3D+tLDBAdJ6H4TeyLKbkXt99cQPQoi1gEHTJLQrgQw8se
9YWkfSPQd2SSRUwekg7V54bgWPIwOTl2S6DfaS799K/aLy6rv0W8RlQ2zOuxh8dckhmekkIMmZdj
qfUgQP3a4cUESv4615UiwnYnibpNjh1bJwsf7GKMSz622J6GbXpHdc9dyNqk2bdWqFXPHZEoe7G9
zwkiKwZfokLedw4jfb951xlIPZGg5SYRBxCjjHplB6rnJuM/ePwCWPZ85XUGdmjIu5nvrFrq30qV
VawRdLGIdrhq1pQljZNUrs2C9hMMjkkc5xD7Q0HFhx1swscQxTvpJrA5omuEc3PkIMqV+iV6XsoW
CcMTuORIytPFh8fbsKL0dWIMeQ1wP2s23XhuRzxT/gM5m+kn2w4jWh7fYLXmWzzX9l5iCP3lk8po
Anf7E5hhKCeQeDxiYvbwejB109MVgxtM+Hbvq/sGvHX1KMVSgywZsVGtv2B7Qjmdt9NsX1tqsMLr
ZoLUofL1i7LzbojEXUy19r8w9xOCCJI4y692Rl8uwBMUwwPpd5UmHSY7FM3J57M2zSl7qe3ixvr8
mLkOMXo9IPHvLRIGUpHyvSGsbrLLpj4evzERxdbNAzWese/s2Orf7C2KZlhNN1jA9leYXqkdOzid
xoLTUxYZttAcbadu/k2G3hFyz7Gst5dKl5qlDOu222m9iElSERMl71Te+VlvKZWQ0rrShrbtyFVP
931R9XhLRqkF7D1SI6Th2yC9JD1reU9xF9zCA+qR5YjtTKb5ftPlzNXQy9vjuJ36YBXhsCvTC5Ul
vqJkOe2T2XonlkDToxFZAm3uyVFM7WtaRMOrZPtCMtsMFmN5uP+1suDhuh3R5Fbye9hNxgaBV64s
jc69nR01xKP8XdrWuPgX2x8RzRvaA1ngDhW6Uy5DQhas1zKbVxLi2pt/vaOP48UlZ1KYjWMEgHs0
/plRphtiMAuRKHz8NnZiHjvsMwtyueGR8RJv53XHBVirbCZ8dMUcWTp/sJeJ2puEJHavwTskknl3
2k5H2JBXRsvJfW3tSO7lEUr3AGDgQFLuOs59w2ZtpvRVbzjf4qTytUGhkge2zqMxPHa5D7oeWjh5
x7dyf0tcZrDATcweSiwEFLQUFH0ai/UkUM3cqxIlS9AKNgSRYmVby7YnXHrAS6evF5iqJYA7CEmJ
1xyKb4rtP6zuIJaiKsN37WnTPLZOOGZAnAHoi2DZzMTWa+mrr1JwV6Kjf7pwJdQJG2CA83fUWYsV
4JnOpoh2mJHP/R55LjdrY8njn7fW/YvFvnOwHPv3PzPA7LOD+nI6Q3XqaendGbNge0xdJuatXBYk
b0eJS1pJrGViRMxE97GNQVHMjibelTBtcD19PHw+PoB7gwx4XPqD2uKgQZtU7klTheNzqIvOyXJi
ExWAe7uSbL5wU7xzYtomneI8UVo3hQf9mgvC9iIKo3uVrMDCQQ28XeQSd4LXG2c6KAaymQ9Fm4N8
tWvXmv5rEaBj8yXsiFUcdZJwQFmrcvR7QYRKPSyCsbLfFxJp9cz7X3b/qPda1zAFqlt/bRvHM5Tw
MYO1oU6K+TakSGDClyRV5V4KzuLXHMTYOgNX5Ex32GnaydeEg1ohtrKbG1nHiwZPABjbbTmcz16M
QCpMyLJlSMaKYDPlEoS/7iBWLToaNil0lt0rjBy1SOX0lhMdaeE+yJFzQ8lf68y0TWF7a2Sf3Mik
wCee4TlVINmIbXt9sdscJ58tMWQEgqx8Zc6g5VPmm3OjsL57Li7bWw/bEHBJzXJ6nQhgmZISP3/e
dcvqqHcFfHPE/EWYHArqZ8COCyU5H6o06P9WhhlpJzIToS+j4Tjjos0YREP1sRFdnZKJymc53o5D
mKaFLumoUg4cG8Mfo4yJ+y+EL75H/Dl6TJr37Kr0oVr+wotAfaULat+ry17mmVkiRBsZcqJEATOE
nNcjPyTrkeOyfZLZf5h2Ft5Cbi7NPRcaNq1m52EluwUiwp9Mg/umEbLUlu5UovWbe5KSOCIuXCl+
y+5jc4uTO+NJsNhO9CpMGYKaZqeWZMT4AFZ8yIayDHNDZE2wAQBIR5aU5hSj/h1PoHAXy6q+qNTJ
T4Fh3ACIbz8Cd24qtD119aJYmvUhVuJ/CtF5VtGKAhdzhTb2FVYWLj9XW3vvosdrzl/UVAjzQYB7
0HxyehaNyAHcNg4Us0ODv7e/kxgDQLWEM8VFUYfbkkXZAIK1SIi2VcgGFnV9AR6aTVpy6ghTq2YL
50cNQBV+VI2DhdKL3UNQIdvh34ClVIKUxLIgeqRpqKTf8YbHMJ5+W6tl3zPGbrLOjx5wiDta7kLh
u5hpvY7Cgs1j2rVbqhlLbV0JoW4CM6n0H0VKAih53mHyNsGoUJjna57FVKtC+72ZH3ry2A6nAfQB
y16OENYy9QnHfDTcVTIx7SfrxJiM0PWVPyklaba238pSv0oyw+jdcFlN0dUPSGjMtmvYzzWfgjwg
BvX4ztQhPEUuORlBuql8qgjxb9t+hHKXHf/fZD1FrvH4FXYpCCuq9WZKgEuEg9uFLcB58nZPERpJ
IhWkv+YzrX7n+gW4HWG69GA2PA/0FPmHXJ0sAyJJLO7l2WO7N1Npiic5Cz9uWLZg8A/TgMrq8df1
HeFcOnn/oVwncBmPnLBo6FWshGWnIslV9DKmfLs+NqDOaXS7TWdtfPSApwO1LLjYdiRM9dcHOtuf
ZCf9jpidI7xgaG9uuWSVmgjAhO/ZO/ezO59czwVW/iJwZrtXwf0E79FkGMPw5bXJSnM1E4Hcpytn
yvfDEKrBvF+6xwdzX4gS3OKu5F15Nc2KYcAk5E3i/XFO9VL5JXkTKFUCm6cYELzfgtUx/Jvfgu2l
6EeYPXF+elzpRFEqo8vs7/vpKaYDntWpP+U1eHnxvCVELSg15sZP+nRP37KIiB2rwfe7GZN1oNPc
45/Z4cxsn2FD+dC6d1lQxOzIu1PfKSPQYItPta5Tcql9AUjCMMTGnDHYV3mMVPkA7PdFQWKh2qTv
Ich9Ho6+vSiumOsv80ZoeyAeW5GkXk3u9m4VX2o1RsURvRZuBWnh0UXEh2MKLyR8noQjjDkVThK3
hEl7Ppnv3egSb1gNSduAgMVjylXQ4O6eyLrpbRwozFKomACV3RB/KdniLPZLDIDPVagpk+vnUgAI
Jp9PH+RWlIZ4wvarHv7jDWIoZdFYkvXW+lg++FxYtyphD2qX0hjhR8X9LH4qQcxD5CtjbRRY/eQ8
ikpbSgvLIl1mhcnuXWutMccdnA8xMFuQyh5GaLza7uWHoSTeknad/125+OAw9AskHcohZJVTBDbo
Otd7Ny89DRHdkg8YxIrAhiyxFN86E/BL7Gaurs+xDbTZS42fur7qDEC7p3EvKF0Gd6YUhrXYBIhU
2ic7vneV7iR+EEoUluWuIuUybiHb14A9NW7UsBGkV6X+xT579uufW0d1RppodNwLtzKlID2eo31u
+OHwvuAW6eZsc6MGpmXMCr/cQ/k9yLmLnzKuxcJvFhbNjAa06tq99IJsH2OA6mw7+k2gUlrrIWLE
gemeOVGCuqCT20r01BC4MHjWAUzm59ptihg0zbKYR+vyCaay+A0wuffu07YWWWoFa3NQ3MxALgvK
XcY12m3SKycy1xDqUFpZCPOxMOFHbb+G3rRBt4ro0Yo9Co6ztkYUCXm8xlUt9NQLl0xZOYNlDnj2
XR9yiugYbu1q86yjPUIefA4G2kCgdNBQZ5pplRQZyA8UE50VMJ20qqmvu6BZvIJYy74M2iYY6Qqa
7JeK9y2kqB5LLj50jdoPezXi6yUAR61d+Dtps5dkiLew1vEJohrxjJzWkeDXiA0Gt34bfsAp2Ry0
CAX/7iPdtTm3FsgAq7g32XmZF4+kl9w+W4sAuXaWVEO+6aS/sLqsXjOo05+zFaghVQ8HhZs5daf2
TJpCwmdzAD2cTq2rOHChTadxvNB1YQGX9TFvRFLG1axxqKSIMf6SU6NN5+yvWJdel6FP00F0aAoW
IIoDkp7zcbekwEn0yFWRhxXrL0G38kVbsKa/LZxrjopBgzKbczsC71XWHtXhWMeLH6cgpUJCBKUg
8gF2+1HCxsFSjyQ2aiRDT7Bm8hiOEYTIPGY2dh31gzOPyDDuQk39tmSdbIlM38rKju4ciwGzMyMc
jIEPs7YOd8+x4hG8f1VrNepPilU6Fh5+x/sKf0FMOwYkEzkIhGURnc+pBxv3yyhknlyMQD1DMerl
V86stk5i5jqLQhcLs3L7HiGVRfOfHzM5jHUMIij3PzaCFK9cvu+f+Z7Bbo0IC7IBoaaBPG0BDVhj
4v2sRdXQReWjozdR0ygdgDh7ByMg05B/j2ITrgw8GVFR1Yne3WPk1xsqGOpGahRqHLhoCt7UVsEr
HtDOUye0rXx6a4T/tzQ4g2D3BIVLXkweMh124fvrzssobeVFqLqkaTHO3X327Wn+RhSK6ZnuaLNj
dLa16pD2+wsBUNhQ/56OIipgyayIUi/+2j5pHmPJg4hf8EqRdu14T+iORaXrN2xPm4ddhecj005P
BOuxJWUxldIrGOUk+j7Zu3x31NuDSWcp5sBhL64H74ctWnlhP191zzkXY/pz4k+Pr4+4P/vKbHl/
JTIdp9vLzPDDA7Z7UYG4r14kN1AhyZ4UQdD+9IOz1FVXoTg6sjDBkWr/zKC/inrb9SqCgSOhhP13
nOU1AtJ5bL9F85TYfeiyuHIwk51XrZMW4oZ5jzNAa6l3h1b5XzWJjSGgPUvZfC3Au76Zij2VrZex
/xe5ynvrcqmmklmqHfoycOvVwm7wES4bG2iT3LCMyyw27IZT/+9DrsfsRyKVqM+CivCzlwpRL1R0
vqO17WS4aq6mkda2uHngfwpINov6eMTFOcRGiNXPk5squxhdBIL6TfgTZwEQNMRvVtGKDKZm9LX0
ucRF4bXXpploaYujs7bA0edQOo3YAvrXKhzx2rVUzQhWW7Exy80xhxbrGugUSXGMDX2uUzu70GfG
J03yLNGYAgqXVVHjTnkunxDacWK7ODjOtI3/tpI+NQYM/2b5AB3hRaMh0R9sWEA6c3V00pGYP/Ez
+h4Nt+Pq1UuXp3JdUkTONAcwNM9Ui8pI6CSxbBFVqzfQRKSLSZHfXb5aGjmSgJ8nQpWIqY8YYgSP
A8EpGGgLYH1KIV117lgrtyC6Z3w3FDs6d/srtDkbqtIVRgLo2p3X6Bvfu1ZsEyfuNfsAhU8bLBfC
6mgG3hVbGPKN5FopGzePyAZK9+YSNK00vcXj/F3FMPUHPGCkQJHLX0EneERG4smokyCD91MaUDzx
ielRWip0pws9z8OVyaNK0ok/p4ACDQ8om5wckzgWBASyiDt+uJso8V1Vsa8mI4tKKfd5vtMI+dk+
zzunj+gujS+DVcmn0Tj85fIRCvTpqiri/kV12w51J58mcHTg948X+bKUFHj1+RtKvyGnMQ/0tn79
r/I/rXKgaqqsAW7ge/Ly7FMDZz4lc2thZpTaCTgZsd1PGX46D2U3dlAUwt6CWbtzJEYlvSxXECAv
ck4cvJ8/Eb5pFt4/jATdc0TNHOi63ey52gzxrVM6V4J8a0tRvtTcCJHwWxmU4VbtvXP3vi6ds41A
zdPh8ac6dr4P2j0YoKEWHN+KCfXyAJhVWz5tkR1xISpw5zwNrg6JwjWXBAttqtGlP0lNNEzkA9JH
1PNlxESOLp12Lzwwd6H49olLf2ER00US3Nyuxcx66a/aRZb+n8cxniq0K/OPzRf9FFX4sfZ4Z9P1
LUA3khw80cV1wpghPhIoORGgfpk99bs6sYUgpKLV3Lsl6zNHl45XjjcOuPXMTtHD6e34RdSTuwqp
/J5myxDINK3xyqTy9Wt2lWr/vdXeD7oxBe8IUeX+i96uZBwzlUfrLBjLtBpxa1lfmlSg4CiprLa+
QmTJzJmZmv3fjbgQKS7KViIIPZDVxB8Wu6DCy8m+WVL7wR50Emab1A87WiVjFSCeq2BSBaGXzpoX
ugi04qqcqmgdoGw0vDZFOVlRD1lYvInsV7rxSACcVYzSSWep5k0arUIQnjXmvwUx9GHEFriGZUiz
qKcMMmJm9IO6N/BL30/kewQttKU+BTeDGrs1g/J6tx03hxsK0jA4Cljal9C9GpYZkNX8D8dOAAg6
ojQH8TfPLzD+18w3LktRhzZfyLNScdjNU0YDaW62AcLUaXrWqSOEJlKftm2gbzyluxgM4r3FnMAi
LDT9OG7neeIn5H+aXBf6WN+1B24VPpCMU0IHD8yi/knkWKru+fPAaDCjkini7+h5mt56IR1OVaAV
YoEcw3oRuc2aBvFdBpbC5fo8NGodO9nVIac84BhbttjsgiIQbkzSXz2t8MkhLB0NW9P7VtbpS89Z
EHri/Tk3ugzfvpNa2Fl7u5rkk/C+b5yXTQhrQ/jNhdwWshZE5/7gQmfHvSpoxJ6+PWJHNR+XG1Nj
HogpUSfLNZhLjud5dXKnJAKUxeZ1ED+vugKzcg/4NlufEiaaRSQB/Uz8JlJDkrLOhRaH7rZCJjbU
fN0NP62+u+Zzd5jugFbk2Z103hYkIiCgC3P6BXUW3kuYloMnBIaPvaGRrwXZhMGWxWJ6v/tPvx6y
EhYgKYqf44dFjoHOOCZLBzWMUhaiTpSu63PeUWmNOqXJ5HmDcdDIlE+F8yUs/Xo8b57uSuxsQadU
MMg902dx+ZIjKzjM6uyo4yEzH5BkkzehUqvqIFFckZOJvwdhi98qH3lVp+Wb/J12P2UOe9nuCURw
GComX++1A8E9tI2GWoTgkcOd8FR7Rc012xowkKtIJmKTtWUAEZlEZFdvznH5qtixASdKFhws45FV
BvAC/H5CuP1j0CoWUC4B+fskHT7TDR/DtuxkbcuDC0CqFjThjqAlOjxw00oyt7gR8eb9C28GStED
1TtAu+tBl4Yl+7jcZlAqk4hS2HyIWjR8109wyUH83OzQSW7wj9m82cfUwu+GP9GJUl5hRPkaPc1w
lylyYSwy4CF/H6PLERk4n2MPbU/ETE0Gr5l6Tjwqav4rCoOH5pls6iHPIsqDBkeiS+aq654LvxeU
rzhXoJVR3iDoKyEp+7P2qttDJn/jVFWRfWZEYqWuuC2CYOebGhVIUNOnlN0Wfp+cWIamkCa1sTX6
dTfjBPblyytBk5sUlHSsjB7mpZXPQQYCy7f1lFh5LxJ5p65lUE1OH6zduc5Aq4OXhn8bH0glcl36
uYCFTnEAMtC33/C9ftUtSl5Drt4A1wAGIV6WWKVvUEnWQDJjfiY0Sab39Y0BM9yIMhsyJuj110OP
learTG60tEMxTeub6Ylq0lMy7zS5Hm4elbSW4OEoUvTLVI4vKnV5KE8jZok1s5chepsJ5WQsg+GL
E67hHOONtnnQwfqsmumYTyh1GWXjbdAel7HpiOJn1IpYmQy+kqcGQjTj61kkumEh9OPQfBtthrTY
+4e06s30mkdfL083MSXa++HblV+U7HYLVPgKQEsuTNi2v87fLjVp3clw1go4SD6LNk+b6IWq3Xgt
Vw6gFWiSbxxu3+eMKJ5KqJgTDYCmYcrPUB4IvpvDhuDV9/oAdslMzAlwO34ODQD73rBA9UZlv/a9
rekKCxpFXEZ3XCJWMMHoF6df6U0TAztsqSuswRuWQJ6GeqemcmVrlLBLBdyPWn+w1onLF7+pnzJB
B4o9CvYbLe7qNMYemZaYaCMTA3iU38EDvT+I/znD3scCifZmj0aLFnZVTCQw6Yt1nl7W1tt8fl5y
6DCfveGJ3gSvcb3Td5g5gL72DJQCygHUcTfMppDvARcNl+/yhMl8sLxMi0rqsM0C7EA7Ygi8+PS8
7wXZUJi+h/kbNHvRgOSLWtekCiOHRTm1bEzIuDqZ9S4F1Y6gMGbfGnelPl4CRRPkUlAhRflk/Dsj
7VJDRcZ3FjTC7r7Muy3sT+duiOE57Ta3cdjA3OO53mHbhMpDq4BadIjJMIuNBoohpHKdixCf2+Au
EcTwgK2FqEj5TyWm2vHBOkwWOcD1mWLED0+iCWCAvQFNCyGhG1FdiQOQyoCVM+9CAkBcgaRVMSkR
mUuK0hDAByKi016nHJhot7XjciCf+ILJWidfeFG4u+usvv1lgA5HNxlWzHP42KmO+cIou4W4LlrF
PSQooxfW6DuYqOfyThohgU3fS4rnhPM490tXS9ldDgj3Dt5OOBZANPzoixpjCA8eMHKAKRrD8M+B
l/kdbm6g8uh2jkojrSgwMt031YAPc8Pt9CNvyoz14UYPtm4QlkSoP3/qCC05ty+mJgwy7VXXbzzd
d+evbs+9+qg/FmS2HurwntOw0ElYxMCFRpbUDWppFQdaZKQgpSd5l1VJ8vPxRAtbWb9BnVbTBsUR
mTmfgpVtBaxqvMquli3/Q+MRIy/FrLLG1VhjzsthV4v/tpQ5AmSDmT4TQQ8/BprL+Vm08BZb1Zqp
gtuLJ9qa7MW1NAJXl/EWNIuQDTPlceoL7kV+Vd9k5kJQRi1QN1kKft/9PohWD8JFjxhlq2IlAoRA
OJapA4SCCOZ8hQYhTh6AGkSsVqb1ZB+B6E4nu6JzhGyLeDXT+7BaUT4a7fnRXn1vE0nMw4Xd4wXT
WW8E5sVIN3YCPBrzDmwKLKNe0WHrDK9pEF1HxVp5vDaEFlcTPB6L+qB0PfkbkZMLDiHaUP6uCl99
GMS8kypZwwYC58BF39E8fZH7CC8W0wOrJdSwB9bA3TGG7wOupsUMfA39B1VcBnO1c2RUuVhlVRLH
fYRKnBLnb+/QbfMQo5iHhEd9EgC9PXEpRUqnSfvw5U13mwT4/4AANPw9U08q2rzPAj/k3Tz0RxJn
mvH+RVmbb54aKS/IQWXnlGcYj4ViuJxsd8E8TSmzynOcElNogsvEzlRv4ngpUL5EfDePvPDAEgyN
J2+WPmUtkQboQqZ7lPv5i2anPF0lMeT9anV1MM3vwGDdaiY1d5bgWiXTI7oJgj4Ft86eZlV/pwYK
14ASpZkxl6MKOwF44k2H5XzdCQSJxoptMwRBWlLnHri6zbDwdGyjITsrKOyMBwCCyVExhPr3HE3+
CPOeqWB6B9WgnHOGpYceIH99GVI0V7vcX8E/Vz2adEA7R5rNGWy96XbkrVAQYPQsmJCmdjS6xKjJ
QzDzdgwb5wmTQdLjmsoAGf0YCFrvbFuskh+F/TTWlw3iUCJSm/mMi+4IhlBtwn21/qr6wiCThf76
QDIHlxzOSAzlG/zJ4jaP1Tb97sTWG/98YyRiB1nfeGvGrS+mQ4RaniD8CNWwBjrKsvExa2f2eEeK
t3qlZ0BmzAQP6kwxRKYz9qnBUXfMEn+XXqTgRTjtLYqwqETQykKiCYU6H1KJ6Lwhhk0vU8bUrVXD
8DlLg2JL9EMRnVdkKJg/Rw2TxCFKawtxBHD8FHgvZR5TdA9kmXdmbCmSHo4S+VDcOYd6ahjLbYNq
+TylTSq3XaajFMteaVLKB1Bdor6EO7E2hAG6ATPp3GssROPkVA1Q2shoLZylcjFVrus3u6noHl/t
b7ko+TeZgqJSz0v2D1qq78H/5eWhHYTH2IUHlcW38Np31LHiXOGC+ny86HP1EHufWvDVNTz4Ld9M
V9sHbsFwPOz2nXcV2Q3Q6OJq0gjts8H+EZjr/zTOOablDjsWaYvDrMiFOKs6jchxscF8ID0rKT+p
dRWxgPaX5FDLqBrLl51721n8ag/kBXVdNlgYJr2fWJiukwXeewerqsWWEsBqw+sPf6pMOqdrtrNd
ArsVfkTw7oMPCyJzxS89utP6FuVXphpsQaQOnbhfE09RCiv06O53xsOeVDkbPRcMSIzD2Tviz2KP
K+T8Iy4fodCvYXdOVDn1j0Bs2LPKWhqFgJwrpXUNuUnhpxctew44V2ll7CrDV8Y7yMcItchT/iDC
7vUlb8oygrjq/hMeVBqiDYy/pDwKPW7W+p8yIuDUc5bnKtwUMxgpX6kNGdzD5ZNDZ8Wyi1tq4lNR
oargvzfbalGPFO124V4QSlIvHcCS2sfY5/KcIaPgssV1Bi1aDgUiTPEP5UAYmm/jz2IXT9kxJd5v
BY2h3gzmeUU8O1hijJ7facPP1nNvoTHWYNvuNJVt4SBcc8fz03Lr7MF4TsihmO574PETlFyE8Bon
V2MdXGvppHHdDL9nnx1I+RMEeM4wCuJ76oqW15xC3vls925toG5g8WDc1OqreojBSMb4hKFj63vu
ptovSxzP/mfH3xdA0d37KuIgBxKqNEGD/SCE5QRVl8763+1GvNZK1zQmQjthLcDaIXptkLtDfG3H
0NkApZ/YBc4sn/0jhqRb6qsL9+dTNkoNLkV9p/hnwfnEvSsrm7zwqBMZK2fsSVXAp/HBWJdblqR7
pKoO6AaCfdhzMtzG8k3f5el5rLYOtraDzUxy7Qmdcv/98WxrR8C6WLD4MDlxBiJflHTVgK2Vq4LT
X3r642u9xURuCFevE0FOyoJMO6iENFu9TlvPV/Jn9wcTlgmIfNdz82C8HuL3B5KtFVjb61cnpMqe
MrxzQCQpYIRcaY7zclLEZZrJYCuxxJ3t4IX71Tqrcfz1B6NMKx2oYNjTTgVmBSPOwZcTrfVZXpdO
pPyvihR1DoM18sixpcyeAbOAkfHayav+r9qQZ2sirZ3CMpBtOwh2cjMP0WTmyWk1rczjfOZiIr4P
tXJh1jJui65uASIJksip39ClEUP7UFXkQZIAWASnn9qiN5Nf5+gPHLaNh/HcV3QBLvJ/PgE5D9/a
30UJdC36M571c5WZ47/OortPO15EvrQLIVn6N/zXIAyvvtVqsiWCbn1SNMYBrdnKpY1Dk3TzMNBr
BCsUnxiPfTtR/0itkIHOg36iQa12R/AD5CGmmrVXqw51/Rsabjk/AOFyAselxnyK0TSS1L1tHafD
Gr3K9m73gSolRXY6SIIB69xte51DG8cXwMI5bUq94tDoVRprziUm9vs2SSaeh8OwK8gcjxk+8bnm
0nqQ3mW8QzfOgDOeSKSXBzVn70khjCe1yk7uSVsxcKokFTETUeiTBWqnx+IQodpDr2mFx3ZiWf60
2qZtzEB3lLscWN+LQ0bizR2fNcN+WQNGm3+IXrx/8/JczROEH0G6vOW9ZUsh8yX+JRiCdM1SlvIH
wAT5uLhG+pqTjYgkPe/7kuJ5Ptepce0ItGAdVKxpHSVydj91p0LkYRQ9EVU29n2OgUlSyWT3d4ui
wGApPoUDL6ldp2i+QQxhrzY+w1imQPTirzLJeM3Ko961P4U90oXjY+L/ILfVE0XjjdWJY3Mqhcq0
9jraZZ7TepmtkhYDBEc4BWUIxkpkTl3cmL/jKUGehA5A8OmGfAzZcEQ4JvBORV2ti+WEXg8EMakp
o6Y3jkk9vzRye0TtebNyCEjuyL1EA7zyhRRJq0L5tplwkm7w90DbLJHmBYs0YRd9855uU8Gv9sJM
oTrGPh5TCXE2JgOuM+IpWX06BLCZ/baYzxlAIznLEuMFVD913/Ko9Rs4GcX5d4pVSJM6MeZw+JfD
H5kZE31/T6TzxtrGFNwvVRUwFOxzUb/ymuM5PXjk/43KdTgHIAtPiG23phEsYFY2gGDkpKzLAMPy
v9Zb52RupIVeHg/KYgoSnShcijBpUbWads8R16eI9A2VIY2Hn8hsdzxtQjHwphSBVxu1pvBu5TPz
S2nobBE0t6OVwUxyS6qQP/w8M04RCvSEE71aPX2aIEB0h/g6wcOLWjUo3p8g16mI435YMxEjPWEa
bsJNlhUAvigVAJRxM2ZM+kpThcwT5uqIIhpAieW3zwtmA8zzO0jcAYx35gHJyobCXh7SnQ/aJrfu
9bOZ8laZXPXPxCuGNwM4BF38efTfntesgrBT02fnOidZh00v8gj6tDhdMRikpY7ohOnaVDmRrEAm
eYMTq0asY+gqOYTQt7g75dJ+ZzthlIFbWmszINnR8IhwN6QakAlP8NW7LmsrUi+eZ7nzvEr8tsUA
vvIVzHoW08jUKoIgP33BsfRuLULbrwZItUDJuvaBN7PhT8QXZCzfxObUd58NGsBQyhlP5rlqiRfz
essuZ87oajib+y7L+d+eejidTot1JWKTfGEmpFBtWIBegS/hp2yg3kh4AOqatUSyFOsP4t0CySVP
KatH22b4Wl4EpvfOkMu8Nm3pYotGZpZcWr03fLB05uwKTpi23BIFMJzriw6Ph0ZK7MAefaRngqDr
iceFLYhUvanIPPZpqJYuDkfad5jlt9Zj41nU6tDHxCd5iR0sjW/GMz017P6BdpktbV3UwYqDEwd/
wkQaBvlpayCxiI6xwwLPc1G67RxKfuFR/fHuTlluMOMjiQ8/6W5BBDNZQBAWpaJn+hqFZfdy6jwS
W+x/BUP/16ak6d8GvWwR1OZbRdV21fwXON45t0U19OL2/XKA+eJGbKPY9cewYb8zFxfJ4Ic2Vlzl
7O9K7TSvG9ksnjK64Wgy0MdyKz/qieOriK4WZKFgRjIzJ35M8iTDNuqyWEpx6cmSWLOO3kpTawpW
ZCl5HkAQvSFWf2lxxXgNtH4l09hW7SQqLWbyNFuBaumSowqxEWzUGuUdg8fdt9h3x8JIBc+jJFsm
4O8+cmkj0V5EQUC7CUwojoQ1EaS2SPZIeS1c9NJ8wtwhOdUSG+JKMU0xftbJX/qoOycUAfgoCZ4K
vPYjW+uCmkO2+ryMmGWsMgnF9rWtNusmS4MstEJIDG0Ewf3wUx3VTR3LDmkOZHWo7dF8P941z2ZC
0/uYGR1q31vfqoHBwMCpVaIh75/OOtzHMqJbTGPaGKPkTnrLB6/K8EfO10/WTA1DejLR1LZ9enQG
Ydn0Haspn6S38WOmWQsuJW1LQKic66kTWrmrXMfxqKtZ/eiPXSOTHjVinWHXQEdRv8YhEsqQATAy
8irML3JRRU0naCzoYgS1hrwVUk6m1DmlgejXgg8gvD0DVJB5YTsTY9hfhKDFHOrzvo3A0x/vWxpM
NpGnuic3OGzF9fRDC1+xrHsEys/RJbW5WXr060A67fAY8yDDxFT+YElx6gRBIyZlTW286jzTp7MI
mutBuriRTsKwSCvoCfJC00exRwx4fIajlZR3jl7kT4TMBwhKP9jcKplmpNnm4Gw8YhU6brZjstu+
pnlkRQ3WeXGz5Owdipnnnt671XHyeLQt1zWR/Cl0MFke21j9wudhJYlGTTrtG07K83LxTXjRPnkg
bl4N9ZYXipjXxepvVPt0GvQ8ArKof4iFrpXPCJEk8IvDDfpGWAlDnnZDK7nqx3K5PHEXcC48IYkG
C5V3vpiWLnOg+kiUaZLxAsciJu5TbIYIeNQ1uENrk65BtjuBwyCGX8Sx3YfRemwrZGCaxNMjcQGP
WQc23SN6Edd9J/8NWySXAsnLcnW6XAroEKBzgjORW6CliLtU1K//t9jk84Ck1ObGhn0KX+wslfql
e0uBSOOxLB2xyBiqErprUFIZWB/nwb3fAqEADRlgdgC9oO/5labN4bal3noh5gDrJWqTV6S5jiY4
WAJMyz1mNAZkj6q8xJ/TcU3hLQJG3O2K4EzIQio89yxbt6S/GU3As8BwJKc4QcFulr2iV8Ydoi3d
ZmA+IKRKA2jkjHLvdj54DLu55sFNagvG4RdCwMZcbgD2Rhq1IikQsprTI8xDkgfaTwHx+7ujgbgr
uDB57l6Z2sal6Q4k+SJcVFzGqVyxmYfSErbdtNS//CHqkOrcgysGC5LIQAidV+J+MZ9iZASWxQFX
Ow/ueT6Xi7lphoCZr9k0RqRWP/86s9d+TBq42aHqVvXzMG4CZ4U9EcOANcePE9yigG7q9J6/bH4N
ioiX63qI3PdGO9beT1+vUIP/0bTjGxnJly7qoi1gojl1yMasdQ4QEj7MdVGmCxorxZbmiUIDgSvz
qWUDKnITr8AzQLNY6tRjEwavhRymmfw9JpxKQWI44QndN7KEh4XCZ8IA2+RZpB+Vq7GWVOTejDdv
VChmDK/ZM4clavOX1huBC+8754vgnGf9uHbmZTcsaTfz8nBKzLdKvkYZfznkOwQO8ktXfwi8KK6b
s16bzVFOjGQL5QF+0zl/hy6e4/f9G0osOThQCrtdITqzAgMkS85jfnql9fLA3FxivfK10r+T5Bi7
fhDhLOFhLcQAFJlyjDejWA+Z+aIJ949IDHwp3rIfFNyuzzycG6Zj2alFx/Ta+q8Xdt0zOzCRo/TO
7tq0+lUWOf6RzZy99tPFOo7RLvxhIDGjUsvZTgK4gx0u0mw11zEEEwcVvxn6XpYXEzu8ulY/J7/D
ipjDuFdiHTAm4AD6cPRXUMlWz+DIe4vattXU8B8TAiUPbG10s2Y0BrPPZ63u1PoU9i3MiH7lXC88
GEysnvh8XAY+NhQNACkxP/+frMhiqNrkRBAfhv/c6JeAw7Z2Py3spOjQaDs2u4p8w7g+h/gZda5R
A5Si/JrGQKCxoiYbIGy/u9N7q7CdJYxqXvLQYijzoLh5s2UMk9ucDoV/B/SYvB5U16vnQz1q7sQX
R7DtHG+cUPcjSvlSexNS+qqzVNlNZpyQOSyuo4DVA1UH/eIXlW3NQ+VHODMOKUfWrfSEf7kqHaCT
bT9fOpvsEQTN59if8eGItgZY/ORS2bwKW43LGGIRDvG5E76XnJ/QmMC2BKe8fTfUgWCh+57uUsju
TofGwhc4ef8cvqVkuNvYkq7PKZWadCmoCbzquJ80Qb5gXiUDCqAcDWkefuwmBtlBU6Ra8LeKg5dN
Fz8fVxpG1l2TyriEBENdJm78PnifhaLnknwDGU+sd/BHkOaijBSyveXbdJxFNz8DMMbzefkcIZb2
YysKYOkwLLi70/ipsD53nuuQtp5fMv5MuieF2F9x00m4ZxLMxVdw8U3yC1SBEa9LWzlkmDZSxsw7
tUReZlMQl23pALk/aVeZOtcr4Yo3Qwg3rtIVqpWviuRLl2ilGootMJkL0ouHo9aWP2pkIsCvwbT1
4BpO5CQ9894+8yRti5uXp4gSEHhgVkzIQWGYTdO2M68V3Pa8+xoxrsLZeKIIFEqDzBszFpP/kGyw
yid4Ok1V/T2MImlra0IlgnBItgERD1she8+PK8kDVHZ64W25qRxkBBmEZbDVwPmyYNnfGCmTrsnA
An9nnztju4E1ef/UegvGyMQNePF3oOOxiZM/YyfAlCqkG+WfWnf5HXEY32Dz25heUJ7w/WVdB4t2
7uk/K3LnHhlKnu0PWw6CWeE7RuIjOOELPFS4/Pb/sjwU4jVAe6tCTf4kyT4+HfQ4ahl34M/mKFYp
dW/je5xWoWXPGCQQXegh6xfyv61w4nt5U+j9h6lgKwHmjbTBqqQoSNtPXDbEL0OqdJc/m9W0FgkT
esFHzq+mexNAIjHsr/BA8skLt1m3W03SexHwqy5DPbHOrAC9nJgZXVWw51rc6A0gIimsHFSXdjWE
T2Zh9VKmILq+drUmP+kXfvUHf4neFyT/vjk5DzIuyezw1OW4k5DTAe4dj8J4A06MshH//Q9EvNBV
41wp4Cixfqjpe5xmnpFWLhw2ZFWqO6Zrv2howjtu+lppJHtdc3N7qhy8qtC2HR7W/lWuc0EZz6Hx
KJrEd37+PBijuh83iCg0wTEivGDbfOgn9MspinTtDQxVI2QSNy594XBPi6XpVbTXH/rUMw4yafJX
c4Uep+YMjeUwQg60rzQXI/BY/K3+XJ/dqqVqHfkLl0RjvJn/bMKmswG4AoeG8O0hrqYKjfyoSMyf
+QfEh8xicjiBwWYMUAazXkeovVoazw8OQV6swbuylCsgzG+Ws4gtVNtiuq112wE9iBXAdav5rejL
PqLN6uzYVc1aOG4O7cizBj5rvoRBOmO92WdEpeTvYhdqGsSkrknGKEBgx8Swj0ffjUemVAGWa1/G
7OoYKI70g7OXMtv136AWS7e2J/qnIcq1jftzJAgxcfMIMTh5KiMTEj7aQRcGWqfmf33YJpabrstJ
40Ae1Pz+nE7LagkR8pvLtEgMiIe6yC5VlvJGHbazgjdQGEzh34OMUl+XvpY39+euFaicKlxKgDJc
dw39WJw97ugxr7A/PtWVGvL4wOExWpYklx3JKMeBxfypt9fdrGzASItzyTxNYYf1tF1Sma8vVKxZ
THLkAKJQtGPzYzSAh1iEy+hW1WqYK0hy6xYdIKaImvAM5myl78lfDMAv7oAj+C6w0LbYJMyPKiL1
00QnArEjPv2WvRGfWLu9mTGCxP/cYgD1lmNi6U7Ea73Q8ZH/D3ggIqR5LzPzhbFL8SDQzQqe/Cbl
l8Ak5Lrndn9c3lmZ1rg0XBEfM38jjcf6x5Mp80ll7o4AB+iNIuEKL+O+AKfFGw3dr1C/wkcgD6sO
zf+6sPMwAHZF4UlMJzuC+z6odkziWYNvWyjetVziGDpGmCMufWCMWyXw85j4NCitNM0ACW0hw6GH
zxSMn1jKVnJ3Bsuv7z9aWxi49kPgoljuNWmL63ODVr4vMgLaQYZMqvq25gCGCdHzC6wCIKHF7bsh
vSam3674M/sZXllG1TyxmPJ4Uws9RjWXShJWTNVyUrZXAi6qCDG9cTzBlquYeQKZ/jUsWgJ+eTcO
CxuSsNBPXKbYsDFSwzRmbZvfsKmEwlRKcx7T9CxJr9CFWe4v0LgMZP19RKEqlfTT3NhO9N8VX8p7
LrQ23o/AKZPpsBjClef2szhxhkl2YqIxVTOm4zq6KrLj4rtOuUjv6po/IHWO8bvSWYgw5DDBrsXg
lJHEE6KEbdDHvGaGHqskN/W/CexZWwriiym14E6NobAfeVZR6ofQw1jDp1mXOgTCDSuMgID2YK0G
CGBhwYqVcf4p1vTwiK8b4mwo4dvkdV99ynm2Ckz5EDwoRcVQLsW2kiq17KzCV3ZyR0pk2eIe0n/8
sJ3YvKo96QHbv9o6jtg6yTpIJ60PardrRmBWIcPxydpYkzkTC2sFYqgwmdSdRGVjMMkAd/cB61fn
vnZugv2gkd8HHwA3Y70rUC3qAgEmz7Bkqpvnb2bb8EZRJM7YzUpx/JJkKTqXKyQ7gxjVOlyJs7Mf
oUAXkDnQYt1+kfWARB8OinZItRh+Gi+Gs8BC/JP72ZpcNOeJtDksUjTiApm4eKNWxxMkKhX5KGS9
wmmDcLAcEwvHEJm4do5/VOGPa8EdHuEccRiKbqLCtvMKzPR0gs+Hq1a3VszPS3PRMPun4+bKIQ1v
rYGJqgD2353QgrruxGCQpUEOTtMwtsoEu7QbqfJx4UiDKr38f2m7MbevUYtWIK6Wf9XsQESPPtUf
NlNBWspIEA6n17aI5U1j+b0JYv3yM9KRx+/REpdcakiDBF9xYF7ECVghm62yGJDmh/89XzPAiS4r
oVUTxAtbuEpRgYInzlXcB4T3G2lTjR0eloTfPtFOQR+2upvTAc6KCnGXhHbPJworq719SU1deJFs
tup8kUSaT3o4OzIGZ7oUjlECnCAa5DqzmcWKakF0qBzDjLpFQOd/M7YjpfetciwAiG4n9xPLWAE8
D7TigOTClKbJuWW1dg73Ah+Qzua9w1wARzkwLtge4lL8lsGoInS5A9MNBB5oZ3v88yV6fHRckHy4
ZVzSvqR3/GOW6dyPnEbCg1xVrmOIv30xR9POX+ouP4aFmeNbeXjugyzW0Xtv1Yd3lbFcirVzBOJH
2caQ0xUSAjlkooRiB9elZVvkYlRfwuR+Ij0PUq4SfK26uOBNbaoCc0EnHfhXH6PQ4TdhPh4SZhZz
X8pn6hG75YYw7TwR6jgp38QJUDhiB2YSxlnJc2E8NKn9OppmaiF3CMszGLbQRxgKc8VOTR1WLNYi
HZLmkAZnVQyzLKd/Rr8uFqkiipypYMZk84zBKUxMP8dgwLO9qKQt8QPBkc4oMFGbl1r8gMwfU6Zg
iXHm83dpMYyetkSGnnOpMW4X6I/e3DFBF1ZoxamEhbjDTHQ0xj5Mvv3P/V4ifHhBS4HMTF9VndrC
B0LhiSj2/bYN3AAvIEFBn5qDA1mfC6S12pvIG6sW6uP6tMLiAaESIbX+3LXxuMXU1x1U2PdxfR6T
MrGVngDARcxs1Wft2yKCYdqwzDWEVJSSun9ntEcSOo0ZqZqsPBxvPT8UKneT0ovU4irL8obB5Jgw
rRXkZ3ZghlBHUvVqrxNidVJ3gdhe+rbk75mmJegsiuPryRIY2mj81qPo8vM31AJcu9aBgj8I/YhU
MGu648lVpsPTifXD4zLo4GgYDSpMCw+JZx/jhkMXd7DGk95mElEBo1MjefV+rpQyJkX3NwNEYIcr
gjSGYQBVtn7G+76Vdf6S93/e7rZa2C5Alm/njeA4OZ3QwrEzY++oOk7yWuczF5h9D0HupSi/rMgz
Ur5Ev2kQr9Lhc1x5TXZ6cPhvyegntEnwyk//yOS9fjmyB4QkeZfkrSaMjOFUsz6NV7n5yYx8RM38
NuM6eDXjsEIZlrpUt9nYCgOAfla3b1rPNaQcNeC5IpNwfxl3MtnmSu+9yUGBdeNDfS39Z8ANedT0
JyNiqWsuwn0Ir5iwMXdehbDTKsG5LoIrnCqlUQ+1AO0kMv4FCv9inKfHbJ7cSmArcNU8FWrDxvNA
nqNRESt4AfIlySEzxPuJ2y5/3+qfwX+Sv2DwsIFeiKXS3MEGYZRqvujBg5PzG6oDnDp+1id63W4P
gv2NTFBODxnozVEx+P/pTS+U+QUpW4p6dFiR4hVd9Wplo9xL88qDYs7RhbDhE271KOD5y+UuM4Yl
vu31kt0TYQadNo/uTwZTx6zjrReoMaj/n7EfMrruD2U+YAAP034xOOtw0f6nh6WQrW7ctV8I5dnl
t4+O9iSHGBmgrrceC52Asift5m0GS73gDrbtQTE8rchFlcgpCY0rf3WmDcZwp1hRt/wZMji05k3o
kdg2zFCDfvwX+/JBJ+lt88UvR/jSpU/qXhZuvlzDqfBWpgDITksNbDcSzD6XgmxWb3D9wTKQFavs
fFHLjy4L1RNDG0iksZW4SnujUCrhA9bgQRi20hsxyCyBq71lmJBrqCC7uHeYxLq9HBBQGs8Xseik
/Du5Gk9Ri6u/06uStx9ACVeTG7xTig63zgbSWIKeYKV8EnEyv9wubNwcL0sgEyJsRV6vomK0EIYd
q1gNYBxghNBLewCfP70C+70gh0gT9oNJiR4qAPW1rpgmwQsYWaSUaZxxA73YIVTdwoRQSjgy4xhp
nJUE7SqnmheMlNBJpmycVB7YEEy5EqDgVkfWiOnmgWQD+Tl2W5qNIf4fbZnYmMTP9s0vmRwxQQp/
ND/0BLezf1tCxDG1BqatrTYAvs+xff0xgoEFL5H9lQMgzuEhei2dpX7jPgAnizXyppJp439DmDmv
rs8kzOL/yJ7k2O25/hXYTlwtPbh0y3zBZ6vA3A6PS37o8z5Ur8gUfL2rVcSmn5WP8/exCniqvJjq
ZWrEHB8tdo30JPIZcZXfT4Pg5T4YwS6ARqY69fdex4u+eNUksPkDTFH2r1CJ87U8O06ahLNwLCGl
Q1YOpYrYtIURifk30pVGdDQRrA7kBffpoplzg9B4KGXnxHf7HVXtHYZM7Ix7L8GYD4XuRfkaH6a4
CF+GVVR+br1MOCD+rrKpClGLj0QJVL0VSDJn1/7Ke+LNR9HQapy7kdolr6LI/icI86tN9nYW/v5i
Niw8CCKvbJKT4+qyDz0wpxmkX40Lb/Jyu1XmEd9s8PrHQisEj81bKA8pLeQNDBKdCk8UR+aYCttp
eOxQHUzXx32lTp2vUpTonf9qBYx3dySIzYoa8+5qx4RV+bigwcuSo1Gdt62QWrOfG5Yg96Yfqz19
z9tho73pqugJ187LfY2TAxtTOw7lZeLmN0vvaUfkd69PhgHGHgb8kLM1SOLwqwM47u7NXer5MbSu
zlvZxs55bESxJYYgFFMod4ThcN1DQMPtpPbgUEdrscZSd0YCzXYlVmTkA4vqJhcjzGpSxhcEoEbM
5tSWa7ahTz2Sf2DbOaKKTEBu2f+rBXbnRvtTdeDScOvgSTwGvArbln8cvkV/KTzS9+54iiWjBH+l
HAnvbeQpnsK+VSZO/IFjsJmH2JMIHll51aKJPCSMkVWnvNTKNmRBqeu71kc2JvoHrKvTfc8jxmUl
ZNKMyx52v25PFXNUTzZ9j2WPevNnGu3/pjBFrmQUhNW3qeaRHmkkHZ4TTDXIjQra80RtJ4Fb8Jfh
sUr4+K63PNkA5N4B7zlShFrWRHOfjm1pReVmYeEGuBkCkuPDAHix9MwP16LH2YgVQm6nuTUTenxv
L8c50t5pPcxZ2dVKUt8Beya36OiQDchPCZkNmMKBTsMdlIt/Xe6FKyDnDpT//o/vdpd2ZEacse4w
S5XWrKZ0Lwa+sraoZm3wSh7Co+UViuuqlz7/J4kjCq3yT5NH/jIljK8Oe/ri9sSGSXdAcozxn+Ru
ifJTLr9Ntv/llLfM3a5q5t8XpN4jQ78AKtlBCx00+bRl3UEoec4KrRjY4Kwj2VwLWMVUYLeD5fr2
BkC9WstTVtZ6Sbb5TgIjcXmlLeLqW/x3s664SMtMdLSc2K7Qq3q1i00o8g9XDk5w/yQ3k0jcfNWj
OygdyswA+ACfUyEWixJz/8sCu1AmiykmHcL6gH74rKPLmOzThGPGPPXN8iwzbpNX8C0c0AnaSqAB
VUzw0WBobyfSpXiIMhoDJ+8eyqqsaYbQ+s16pFnRKdQBm4YWzH7sYbV0NCD91X3ZjEDHH1MKb9pO
DtHACvFR0jFPgnJ72xT38FXQCF/VI7Jv2Ezg8PoS9S2Rou09/YcrmmjzmOjLb4MOr1RpvRTJbQ/B
nAlD+pt8lAae8TaZaM34U+QpVSdlLalF6YhJLPDq0HVoikv4XpbMG8K7B9h8JbCLyZ6UUUlygJLZ
w4fkWWYbtJerMmBPZEEKJMJXi+a0u74JibA/uWW+Aj3ZT65Z9ZOv/r6xPDz05z38odY3i2sXvwBG
l7M2dz8Oovp68IzXIvV1wbkBEAkgIjV5La4X5i1Aq0M6JwitiBUT0iInwFeWOZw+9jWH+Y5LrNME
9rw3whdcvxOSVE7VClXBQuwWdpy9iv3Twfn1ArAhGba9lm3f4rElO/GDdxlXvFdcI+oHYNak6N/C
yHsP8zM6dHwyHZSU8V/h265sDP7qYj/faNEylT+ZozCfoBrq8LHQUz0H7ycbO7srTD4FWshtG5uM
9vVTjCfHWchf/L+W6hHTBO3qDtK/xJPglOuNvN+QbBHaVAZJtVqCWTihM+Cc9s7fW5nYl+Wsd9Va
L14kWbF1o5zS7b0VfBioqeyOoxJczrk2wwbJmEM+oVozOvneJaknieReaLgRwK/qYdIB01PO1MO9
XPb1/SUIxejKku3DPz2kGO1r5lkg6vjREpGl5A2cWqnO1rx/9+lth+2X/O5fz4kEtoUNzJ8r6QSN
dAi+QJo4gC+LHK+F4WphD3VmfnXZxmbZNWx2qHpFDdnddgapzOQ/Cx+uIip6pmKT284xE4i7qAQY
lb9xhwkjrsuH4Dy927MjwBtRHX8hzJIsOnx1P/DcUhsdYbGBd2LFyO3kj3/C4YWxdyZfdhhtw++n
wXvvAq4R5QD/J+jurttgp0BpfwuaLQFnZ4i9YlHBv09wSivRC0iLNAMBdvb+UzQ3LRiOx+HhZDro
y1bmnbOTsFE7TAL2jr9ckBx404V0RG/36g7+J6M3U1U/oHNlwAtKTAanyj8wTb2Az6EZC2fLQbVS
q13mQvyyO2tlbDZCEUQejst2hU7//XwzZaxuuNAWGhfDkTmdQK1TOZvi+gYHyoDjzzCjhYGjGXSp
V082QT8cQ8mcoBrT/KJltCY7UvuabiCPjblaTTTUujL3TLUyVq40K5hMdfyFxmyOLO+spXyL+OaW
7OJmkVaOe89Ou+5bUse0zmXcx7q1BGUZho5aSxci6DlrPuhnxYgX2WKNOijPQTgUacqrkdgAsRWk
62N2powQB641u1Dh8YyyepRlRuazJZkH5JM2yaHCRAcPRKJ5FESQOdWPo5V++AI3X5FZdMkUeaur
I2PQUidqLVMw3z2X/rlalWb5Z8cLBp7ijLCCrHrE9s2FADug+qXzj5eaMs1pQ0f3U4H2VTNymZYz
Elju9Zfxcty28qPuhvZ1D5HuWRpIhzmDu0dQdaQcgn5zr/1MioBv2wp9eZLXqNr1T73lPnzhykLB
7mcADtz+PeNi3pjtFnp074FemBUsSxUG7WD4JFChu53cDLZ1F/InGNexMU5nS4ssFp6o+HIOQEPT
igig28+XcoTt7MPwjo4W1B28P/JyZ+C4MoqBiVmuYRaFkmLXyuZVUIjFgx08tf0VBZgGXzjUB3Fk
n6UERKf2Qh0+wPmeBf7Q84zswpEERWIh1f0RAEtBZOo7dK7UilUDBQLDz5Wk94G/aB1RQyHYRvgc
TwbQ5suijX4dH9V4g4f/2XyRF0z+8POWwJHVZLCdaN3hnaTFE2rVbL3QUzfAJ8kamtodE64ixzM3
Jlxat44IzXQnRsiyE7H5qfFVgzN6eECIcv3ZsafmPzPpchZ8x/kSNIMKwyzUzQr2X6tjivLXfOsZ
6asobKLrNhR+2FtWyWXDn5bWp9rOrx00VIvOnMlPTNr97k4tkdhhmzTJiqwyXmhpDfCYPRfPimDm
Ds8JgBw+1ZsXdmB/SElSU+t9YGOvW0a5iYj2tQ86YtxZmFdI/ix/1XG3dEME25Gu0CDuPzeIQA1v
683q6Bcd14AF86iGNV3D5jHuTI0HB42o4ojJ6BxVrXeaz4weITr2Wq2/Vg2gGoUaJNml1a88j/mW
r7f6gjBLdDuIKwU2uIO0O8ZhnxqHadVOtjYAgkgUp3pxMfCtRtFy+p6tBTzNJHqWaa6mAWgMCNhv
naKm2igVR1R25SJSp1d69S7DyDWjVONoy2PHJnPnBVCWmEVJdZmNNVw8/2wl+Frxc5mq2nHG5Z8b
DvJdixvFubocFtg8icVfJH97tg4L5/C7o3alJgRRYDKsYgAct2XK3Pj7K6tcpBkrIRry5hqJB61D
VYBDNhxagyoCsnfX0hF9ro/WOw/9SGV5HgCUk1n1HfLQrIBEN7Nkoxsx1VQAuSNkTArIqPeCB87j
cRVtZtRndiUPeSFvLfqU1jeonKCbgj3WEh1OQw0X5wMlQ6AlMh6m9ZMPWwlGvU1R2EGDyeIRemxg
28KO6jiQYgbSvGl0CH8CkEBDbWg5s9ipdjErNIOZWedsuOgJb21qfPK1cw5ZnIQt4IoBrnPO15Gq
61p2lNt2myawLLHfpSOgfkQ0FbkEoJSdbhx5fryL1JjzcdLQlPd6Th70zo+PEpPUQyoTNcFKE2QU
GRojNuUtDrxzQVsV5IQmrgmLDYIEEKITl1ybcjU/F/n+h8/oMorS6LrJ9cgT9wrlpz/q61jrsRhi
Az1X7A0ColBMO9NWe82KGQB42uamuFFhbUoK5G1fQ/OLNzBo2Do5O72cBSkNAkhPZ0lidvtrLZBa
Gs89TBX6FU6Ayu51Al9vPABtat9w8gfAnGeeQtu3siNx9VqSc9s0YeUHf/MCYhTrO7eGGwVbeB7X
pYOuT48u8nEQOj8R2q7LZQDLop4gZLfYQE41x89it6cBvLdvBgRjbvaXAmHDOt7eoGrum81kLzRD
LNYTd7UzUIXmVuZNE1RKB9pzDpuy26gXlZSaxr/wEAaayLVmbnomTKbjZxZs5krOv7Hv8yQEAXxa
WURCAdZYEhGdMiWHs97/hWFryM6cf4raO1L/Mc2/akeMO//kzjmLrA5YJqFS8MzLuH6r9FsEf+3e
Ak5ZWuZcXvZLmeHQdQwcNNe2Y5PYA9Ma1tom915Bv1WOCVNvlWUNSSPVeMe7zq4Snm59Phl6DQVk
6HzC5gpbXnjzsAozl9Wdytchmpfk+0a+Anaoy0ps+ZhOEUA2d/Ne7p5707HsfNKZMIkXF8athg+t
lFbUmE/42ovS571nQLKOwMkM8iB5GfR+JPFc9bztVmE44O5/c3gCJaPU6iO/6bwDk1JOFIA9Uf1k
doMRBJcUFU1CaA4OotG4+NzLiz8EhXreuNKEuIhqhp3rMhpzEePUhXVWsNfCzXVhTZdOPSACf1Lb
KGbPDdLImPVQ6RKe7PQFa58ER8m+cG3NyH8wRK4mdKyVzJYd5L3geWIgw46kG4x+0YcSJeMwVqb/
3s8phr4cPeTjQ74zR4bmwmXLx70TZypFsguf49iLR1PIeVcAi58VWAoEhNRZ/C6uHKrL5KvpdPpw
O3oCOXRYaKRLqEdJQCow15i9It2zWpPwjCyKcfmiBYiufkE2UwkCk/DaaID6F0Dftt3FMQkIIKks
jxTxJJErovUxTorKihx4sdqZto+B5o64pxCwafi9Mb6394TDGYNCmJpnOTy560cCpXAMlUcT+DsG
4kHtiIO/qgIMm7l5CMSfSBhUpJ2v1S5wqapzT9R3p8HsbHnUiBJf2rC5SgMkPn+JPpuc0pMTCYNs
LpYsmS25fuIDW2ElyPhMvL5Rl4D2phFrpY90bN7mtxpm4ofsI+RpX7zS177WLcK3KIQ3nCAlYZa8
Pxqnub9oE0gib2Gn+Ns75VFTBcWg39uK+ztAqEQT6WUf2KTki5gsiMVD584l7gOM/YnkvkMBLL4R
pFfSo4LVuOPvMDhcowsEL1s/k71KdZG1oOl3hLSdgb88HfD4rE0+bU2trWvYLIKcf7wl8Ubki2JG
XnAy9et8At0+fR2xhur4qpwIKfM9l/i2ea8NSQqXfWXGjsWr32yTy1J0IaQo8YgaLbp/plAUK3pZ
YiEZYHSNHuLxiRywN29n2jebBGHn1L2v8XyVSNPwmcwLANV1tsOM0ONLytANoF01UXG5k+B9AE2p
WuG7JdYJR4xidvgIsDOMyt9CuSn5GZT9GequTqv9HW/jfWhBVmInon1qTyri4PEfIngaY/+LAAIx
8LL77LyOb/XJssXDyZT0OeCb52m4D/WgzLmSDjO7Iw5THSfi5XdTGBBwn/tt7dM38niUwA6QNsTL
pIMfsG/8n8YLjp4QPgqYALNajSDoxQmr2FnmHFnI153g+Nm7chv8yOrxw3DwfCTjuoqONJ4t+Ws3
ByDv2gTWVa/VxT/XtBiPrEYVlbjYUQLVNcbBMxDU7roTxhWhwGihGAXh4/MZO6AspVpdRQuL65F9
VGYVx53YHHChHHBobvHJn5hijpIpLv2RSkyBbNzm0sn/0/vDwVaUgqsv4QrPnsHjzp2JsG0EEP2z
izqbayuerTc2z52DsNDwLgu4stn+pp6ww+No0IslNAE/M+m08q5oJD4e9okS5zpFi66Ays9ZAVDO
wp9Bfnry6dhUVg+YVI2CtMqfCY6lapllQNkbKLXO9A1JT42dG3veYpM0X27tk1Rlv+nY62AaY/q/
JJbJ/0sdE6y2Egq7pSM2ye+BL6ZlDoIseXBrzWn1BkB1KufRRN9pflPX7X0GG/A50DvT2YpxSP2b
RYysWz/FGIRI0qhBBtflt6fu3LeKwEINL/DRape/zwBZrzHbdF/dePWmeXi69pKPqMholFKttU2n
Nu2rPkIpbY4qICJWQd2pGCBtcDes0g55VDwzf3Q6XXrFU8QqifNdEo2Z1Fq3LWdh3s0EnndxGEZL
+NzAWl9TNJN6OOReXYh8WVFulgdHaoMfUQfvmyNHQ7NlRwYwSHl/wxZGBawZxUmgKiMR/Aeg8CKS
lUQgr/EOQaYxNeZ+0nZnUxT7M7Mr55XcZmCQi2ImNSrgRfM4SwXD8juwSCHAoo0p/+UU2alVyhdm
UO9HUen4wmc0jBTdSJRX2mKaygCnXCmwkbBoC6r80p453FS23/V7djhI7AalQnlMHigynwjBcwZA
SQ3KcNijr0QpnggVE1yeFi105mqEtN/dHf3Wh3sFEpNkQFWMfo7LxSJsBtfXapRuhDNJevUgQl7I
wgzoWec2gX73A2+JyX8zbosNb67+l5/G0HrJDyRUm+QmQIf7FVfAIdCH/ebPyltH/KFe5VkbAhdb
yRWfd+Rk/cFjKDh4SabSZ5/Af+cK1WUCU64AI+4KZcQ+JHBPPlIfwd5fDlfZhn3cZ/YOej8bjqgA
mMhH8wnts7nmEmsti98U2VXEaDJyFFsOoY4HYzMibpySCkDCCCIawZMgLA7PPkIoQqRCB3db7btG
rqROqQKbDJxOg4uXc60l1tB1qarrIfG4L+++buDr0jvSiw==
`protect end_protected

