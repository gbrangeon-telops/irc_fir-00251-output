

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JtfK/+1JKYw3I976gLBlwV2xqGRbyVsJ3RDvlPNJRewqWZOfwn5MuTyc+U7c7Y8NUZJKZ6RY1Q/g
uXt328ut4g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SKJFICLwrmXfYqYNdiUThnnX5tJzUEdqxXF+PdKpwSGA61whpH8w+itTbLnn6xyBye2kcWPZGi5e
86BY4EjHm7kmXxm6GHfc5MWAMFduB72GxoAF5LRKlUMCOdVsZag78zFjXdMU64ClBQ4zjB8EgXvA
zXBqthWa876wjTEo86w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ho0WiFevcJjvoEEaYGtHkcW737RD7c5clzugQBBm9an3ZkyNmpivYZbh5x9redNVt0HOAIz4unf2
BSVy7qVCwKIsJQlB2q0JzVYTIfuco8FlNbrUR7/BeLSPV7XOk/MTxR/0Dg6meFJjnWuC3OrBGp8S
Ul4C2x7zg4t68SLTuFe/LzPmogzBzDfD3+nozb8sS3jX7ZaQAm/T/7eoy3grLVkFjUg9uj1IhVTP
59FDPnvyx1zZ/V9kzMjvM4XKEW4i0DGLbDEkqT5cZNTgcxi+sBHO7OnQuIvFzoIoNFONwh8iJ8xI
jfha3bFVgIjIJWFL/KzL8e9Uwq67H4YDz6GAsg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tPUgwDCRFsMzMdJqCXSx12cw+CNwvndABCoiKOSYIqrjgxTgSZ1CAyY61ekJUz6cu1q3fnTmoaAx
Nh8wOKV+UbnkqjbXLltbzNbjSEawEnAI8RSn8gStXvDoHe7R6pRqYg2wbvEPk6N6UhaMjVC8JxUE
Nl+LL/ApnNDqgvTWrcs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EyCeFS/0OQO1er1RAmOJ0VIpIQN1auXP1dzcGUAOeSe9eyc/jA1mhBpZ1JPfDCNxALRFgLLGYZec
wCmtwGwTJ9NXiyrouRmXyaKsTpp21jNq9KLTxpWtw00JZFdcekT3NPcfNHa7nkycvsM6yWSUR/cD
frws/8FBuaG+siAqTh5qClTqkxCmbJ08Qh/l3c/D5bCXbr8wXY+SVe6EK7TiYFpV2oOMuwWw5VVW
3m3/ZK4knJ1G5Nn68ZhcGx6rqQE9ZbHMigIgQyt/y7vXemBfmAZ3xkMsYj2X3k1fFfReGPYzTOCE
6J8z+FWVfzx6XMFACHDbKayB8gE3RAvjSqIISg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7056)
`protect data_block
JCi+P0MBUAH58FZo0lqvUF/FoUsKTOnQc691nCxKu0goAPHvXHFIDXXhkALsHs3HDzrlyoJH/Syz
lCXgXwIZKaSm2TnKVQCIRsCCqiUWH5zfPJ83r/q0YHNT3HPXuTQk00aJp8PhV96PP8q7Mv3Dl6k0
kve2S+f+m/SZPjcnHNPyNRxPkq7Ez21EsK376HDW2EzfawNDs1QXdUc9SAbeHexx7ONabqCWYtyL
I9Fm3kzYpI9cNI7woSZHk6Yho2eUfP4z3rdZ/cujs7K+zx35vxgSaR1mt6+6vFRsaGvsRLMAf6RE
qLk2wq5FTNDAwOLmtUdcKOYfDIxicy8+U2/gAczpV3ICeW+5VK2lxTEfAkvyjtXkml6Jy7Ccj1r6
BhHw3FH2fvssqNR6SPfTcyzEIDJYb+KtaVAESR3NP6MmH6On+NzluM1nuZILYGRaQbD32YgmkBzF
WcxACQPAIdePF0gBaZdkiufnBeyDqg9SqlDGhMaQl8xqiYMaj4dcMCdKNpDDsTWshJq1oQh2Cv2X
M+K8+eYrqhnhn79DrDO3KnspztMV2LZDSZO48DgnYQ2mf/d6MbX2I5wj7TVRWTKB5HsxIKnZta0F
aCHpLJGimOb50xkkw6PWteFYgyk9CZbnQnFnF8Np3+GHM3efBBbrVQvc3DmVAabdVB05fagI1m80
fDt92gtEGKh33QtZ7TcrdE4s1X91kVQj4scazEDPfb6O9BNgrmpyGE3jkyvpimNZkI30G2UgZZbr
63q/nen9py0m6MCwar6fzYJ+AT5RdcS5TngKzbjwHLqZQxohP2vnh7utSQL10oPkpzgebuvHiRhW
Lvkc6rk87PpoN9SuC7lOD8tnQhkP7g8GNFfs4ZVCpIFDX3kCjCClPzB4pfFgS5YWv1SrgP3UPTh5
c0dSveT4Rvm1rJVe6XwJAy5dkJDeD/oro9bGcVaM3gBTKOZNBbqqIHMQyDv1BY5Wzd+5/6+OPEyd
BZXOS6RS4uP2BEODHF6u+lZRvlNYfFa69xdOkkxuJfDv0ddv2h0Hr1QlHiescqr/TS+shDMvkhrZ
Ik17GJWvF3RzakM3M+tngy5POzGoyc3zusXgWFpR26vQI5t8fFnEGPPWFlk5kQw5zlWSp/Blru5p
2cyz9SpSopVXz21NY9yD/6td+BnX3+87fRKecvuy2YhkkN1ZLrsloucF5omxbbtjaUVt8cP73LWn
pvLVwk6MAbDxaaM1LkMSsSP+IEHh6VznXm9pDo/HbJ5nfbqxkxbZGhyXFmBPUMSCdTshGn41RBWd
D5KzyY90/idJMM6Xf+YZ9/8SmLJlVn8oRB7COvwt2NubiUCuSvVtlxVjo5or00bngjSFOgW/UV36
3F1P5lR7rCytZrch69RxkkvQgFX37Ac5Tz71qDld4BclHj04STo80fJpQEsxokIKt8rHWdTCSSpK
/CIkX1Zqa2yqB6U2ZJ6sex1AZMeXPNUCXJMyH8B9MSKujfB79SVK+0NEW5rkSaY3j6g9CmsnUrtK
SGcK6xUZemcPP6U8n94we/aXxDcmOb2GnKTNLtxRxeB4Jt9NoQGgnmKUCVx8PoKZk/X6F1qfojxQ
R43LtFlGPv3DDL03NTelxRS+nYEhu5OSJyubN1o2FQEcF4Si5gEPN6N4rU1I9CocASIVCpZm+rDO
V7Pqu0Q70wkaEamtQAi1TrpGoIt4RZ7s8bGRqh5WmZiOL4vUVfKQWuY5IWTGgdRydlx371F5TwGv
C7wQm9Pr2h+zVF0Na7OlIZdsWwvrIGbGagTM57m5KXGJA/hiie4sfwM4gcsbhitebMp4/EmaTu2I
O/GBJd5PlwkSRte9RDUmRe3PGZ1G4H86jDae+mClnW4Fr5iiCV0it/gLxc8slmJxoZvf6IH3Bgeb
e44Q7imXzSysHhc7stCDQzLp075PuoqwRGKPXdABUH3mYWNuQHWR0X7jALHJ865ILNoyhj43trlb
3SolPyNxtVsoslsF1lEsUrALY/pSGDu+dSpda0/MNs2uBt4EQ1jtu89hZmg7Kg1Pthfgu4UU75+M
I1yG36sY5whsbwnSNpr6WvDn5rEPHWFeqMNGb6XIYtdgocZFUXJjKsQlXug0hFyyJnEjLnMJwnTl
6L1S0dG+PClQQPmPHcqETwbpz9SnwsCecL/xdLyBTsuBBP3yzAiyeflrNI4x8aM7487scvu7DcOW
uCSIphbpJcHJZbIZFFoVAKenZ11XMaeAIx2W0FiScTu54VTafHWPE+xUf0NS7BZlNvqQHcRH+iNL
7uDneK0I7r5f0TF+KIF1bFO/m7pd3DXjyoC8WOZ20cOJ3lIw47/J0leFnNAXHZCD97kZlEeTXtLS
D91By5BAbqOa+gyq2dguRtb7mMwcw1O/zIrVqKor7Oh9p18X+MJ7zGK4aTSiXmuMhM70Uon1CLb9
4iYywWCCcv5ZQ39pmO/OyHjLRvEHqJ4suFAhbG51uKII49O8CW2QjeE/CbRRedDDzdpPL0HUCW8K
3LSLk6bnVLOLsikMkQg93L6uxLwnlunXW+QS8bnxqeeFnt6EsguuIVt+Lfp/EugS+r91nHl/YqFP
5pH+CJ+F8jHWVeX8yv04w9z/3TZRHWWW5s8z3LfOUeznoMpVGckUSB4G1/OT6+wmwv4M5vW/GRAw
nX64cM8T5ko7dzl/G3Q/TtzAiXYsnK+7Xw9o/pHo+DeOqz7x86YrHvpnUmSJcSGclPt+kZzuqzgp
JuqF/vXT2nYczJyMCxWjYmK4cNs7HtV7y1VcW0Mqf0JOFm7ho1ZpmpOAzmQMCWjRgwC/s8u3cgZE
OQ0zA/zd0FCmbRFIL+MGtxITyzMw0fNToMAXRAIAJaFED1Am42NHT5MXi+m3BW37b1UMiMmbL/Cf
jwKwXYg2RQr+NuQS4NOoVlsPb+a2jR0glwWH56n3nCH40E2lOqE2b0JpY9eKqJZnE997uEJcVmCb
7ZvzoGfw+GOUEkwnbA1xdeEnlPgG9kIfaxPC6JrsS6IqvVpxTUKpP8RybijwiCzw3NXskFCY0iev
pWzOEtfG6xpSiTPGVu/x5eGOi7YAmSTFH/I1ZnBqjYO0bs6ErBkn9Udc3i2VLEPBZcr+nlPffNmP
M4FFXAHaJlwEBY4wWvX4nT1I4IeBhlAfckNwxItsHO9R79Hk7HwXcO2zhf8wN0KiSwG/JUNS5FWb
HZApMxqnUQRf8bXj7zkwmlu44C6DKKRToeNEls+9LFITCPNO7pD2hEFVn2iWvUnbc/dU0LTLzkkb
bbOOFuxiIlvEN5cPOfp0ZvSQMat4YYCckejYqDr6FUtXwEPtfrBOnorhvknSTDqcwNfB/fF5cgVB
crhuL2onIrU/6WKn1rdEoBWk8hT8o1UGfk9w1S/hnzwHoRKj3NlyU+DdvOiQblsiriGbqTOL4ffh
e7+msqiQXppkvQeabxQYDtkxoQ5A8aR1UQ3qMVgiYd33e7hIzvcXfhRT8whbC65LINNVtwuTpfrN
X26/YYIRd7xHizxWZqJyMDG5hKrXZyxgHWZR9b0fAvI/v01Fxqua622BCd/U3iRuNQeLPAbVDZsD
tL6Lz46P0lxhjB9PKKIL5GptNZDJKd1HfVpEqG9bjTxZCiAfNqGTbPfD4EdSjmRQq9gEoTa8VnOt
/TNOBBZ2dg8c4g45+MkddZl1kqUI6W+xsGGfbNJVNEUYbjoU04sFTHCKWSF/qeQICeCSMOiLBW1U
8MgCzhExV8vj6B1LWDL6DYQPHFOJJOH/jiSK++CWbobbsfJjp03yD7E5bCefartK21J1QM42S4HZ
2S+vD26wabtfHLK4/WxUQo80lXmDIZ+T80OVZ8TD7DkkEHlZeRKooecoeqRL7M4k2zRAWB6gxKxr
F7dcRYDoeukELz72NLaorPZVHDs/JXbwyLNkWr1OTSsrMwDib2xgjvzcn2QXWSkJgb/ukeOyTpKl
j3erIOBS7QpStc4OoAo3/f861dhiqfT08TGUdnVaQa1vTEtixjVmAyXxV+vAjV4abesCDPV5x6GX
MMnKFBwaB6uco2lpjlzSgN8QPBl09FFBohVgrkzPtj3cAwLW7VrWwf/9t0g4NMuLdAzWYPt2haiy
f1gYoL7+zmAYMmQbtj1RwhH9pou3oGTC9vfmvimV/TticuMm1BfKSfI7p9UjnZs+YL0O8jr+QQEn
j49986zViQ4uen5uJnmtXoID9BmxcBuyAQe+31vB5s7EA/CYO7kFPd4XvCa0JqjI8zV3CH4hPVUa
qyXHo4N2A5bSL2FbCshlBmzgJIo6e3K93WNWeLWNbvn8AAdchytnJj6ucGCVXQ+NBZZp+FM5yAIa
OBOhTeHDX8qCI051dicOmx+0tmkAJK9lZKk/fkUQJMw77mTEDt5l5B0gq1H07g2SO/cep474k01U
NdhxvL8NjuQgvx5ygK2oZoB0ZRdUbNjHUfuEnHEXgeDr2X6BAx5fi33zfr/fHTURmJWf80rbXP93
Gqztu22t+1EDfJYjoZ0KqOhgVkETSz+BI8g7HllpENIUebcctBwBlPVIYmUmBc2CDU6QgL8uVhpe
8aPvHg+zv5cWExqWr7HfuakVk9zuSfgJ7P1Q2G6n7g5G4/I4sJIAOPcxpBQlCmvGni9Vtr9TP0qb
zNnLVZa3rUP9tPcIy74EwEiqHOqWESWG5u1BErOwYwhdjVnOUIwBIGgRNtfcTJ4T1bPIAIe5vbNf
zLf6W7albSFKQs1piwGw83E1VSBMFkNPOusbJ6121vn8fMYVphVpyI+2B/ikmngUxXUqqpF8oC6Q
NmsmxEw78JAgVtkoMtHF5E9ITZ9SFY52I/THLu0VS8MbqhjxzZemO3zSUPic3qwijCEtLouMFjqd
gLj4FPvqn9MXbJYUd/XXmpSDV1Fob//y1xjrXp4IQIE6yfyWyii5VqwwUnM4xNQ2FwK0wwbKzuMG
004Qy5Vc5ZQx8VBTStibgC0VeRnF0xL2mxm7N25RYEwgzRLnUA6zNcxp3+AYH3kz0pIh9/J7D7PW
YXdSf+ySdy/lasGk4u1MWLoIUny231T9ydP+yB1qZHpYY6Os2/JWhyyAto0uI+FqCRY3dvU1500n
URXrv2z4CejN5KNVict8o8pV9+QyrqatKJHixiYeepijeq1mN2mG47dAzMAPABNMzUyPZp9INIbs
h9EFQ6eovW1IS+IEJsFFxBGM/Oc23yOTsfFFs+suJDpbehY2DqaKBfivPw1qD63tTyAdYN2+S7qM
ysZyGQrvJZW3OWNco0u++Z143kQk+novH/MU3xDb5EliCtn2/iA7sshrXSVJrdoQO5qrNeMIE/cf
1HeqbA5LUoCknbQcE44hWkp0UNVxSrk2LnqRyK0s6Gbrr/Wh48IeLV3p5wZf03Vb+reKBpfdOxWh
G7q3hg2BYMqj1QfObjH9M/fvNA2VAEBZYmx6niSfoInixtvpLrrl7c1Y2xqexD32NTKo56OItqmq
HuqgTyLQu00v2aTVLeOV7w3KafRUYLz4aOQn6GGLZhesfAUovwoEcts8ayxB7a8aLTcMtHNgPrRh
VvtWQQbZrsL8+cRb1KYPcCPJVIemoGw6WaMuWQx7x4xzLSXlLFBXUaYy4VvF76BEk+0FWVjY4rub
A2YxXc38xWFkmFWfyTUDhCT1avx9l/blkFA++DC8BVzbWkAze7gnzDKshSwOlVs2VHPRctUAlDET
rH4hxssASs7tzvud2RW8BhHM4BFbxfepTUaI3DeMlcacZPeE9Ky7dPEBTU2dAHP+sPEi2UnD7q5w
IvnxNdC8JCzZD0RQawQIJuJbw3u3atKvd/9HKk+a5rZgHJteA9QxUO7+I/RcjEj23LqEs0XNWM5X
reEgmLfioIo1ys28YeocXf0gVf++G7+dLC0LPTDBylYFkcWd+I2jmUa860Bmq0aSsEa8vhTNE1PK
L5dZSOd7IIkOIybKctcRm3e80wuBJLx7DaEDdhcj5OOwjtnSXjNXpqLv2+4ZOrh9dWuM08lcNE1+
tF2PMO4d0+dlKKyHPdgTjyqcNG+FCU8xZe6JMsMkfJMzNRLEn2qpufgUEmdfvL8ZPOqW5r79bV7O
p3wtt/6XLbED41uwhVaACUJzJylCJK0KhgY1FVuONd9Dx6+y7PuczFCfVKuJKJ0awv/ITDflw8xg
HwGu4tpYTj/axDgHn0vST2CbXFGa2DLglgCQNkSujH3NcYUet8QMlannVy2MZtDVKPWYwh6XQB1R
n+YjcRjEEvu23jSuNrMQjlCx6ptfK/MI55+lr+nxxXWZgQnA0D53htZiu+MDeBEoki2nEoZXD22p
QPVofBSWc1pOYeABC4ae1eFpnEiBh9pjLHrTzxR9IGtGjn76V6rn8BB1T2OvYRil8pOqhX1o6eXN
MOS4U/I+2buDto95rG6R+836Kg4MY2G8R0MGu1jFvLHtEpAqunz1/7Mg/cA+yqsInN6AGoaKZk4g
SLaFyAl2wSM9gwlj7FJZ7UCRkgCAgDMsAi/4e0ZLohAK+G5+39h9+9mMmP/xph413d2wy/5mCB6y
m7ClWY+EEK1j/3g+fh2kN6yCi7f7UIWCb72MhnmT9moYNcUiWx9/W0LrkEj2XHzeL/b1c4CVyWvn
Pl18aG7dnGFoZOsIKUtshSZZwBgGDBH/sSZZOuBWEVEFJ+c4/zivbv7Cp89ImK09Uv3MwUqss6vY
K9GgvUWqAf21wYceC3bvTRLrotUZOydKUkk80zBugcXjHRDJKRspKI9uaRmA24jXeXNCVrpKHHm8
kgev9XpLA9pTZqHZBlHWCCu24XYxLGMB+Ql1x/1ZrsE8t6Bhby6U1vnLoRQY46+nV4pQKxIaHlBQ
Jk/Mm/rPOzzlxjjYovo/lTuLffYOzYTub6F2/1DB5rSxiCwGUIxopWPXu1M5Ha9XXT1GoSnwtQo+
hhj+vw5YgeO/kN0e8EAQ9q5JipWO0cAKCIj/qhR6BDq5o1Q/IiZsRzQhCWb2dCnoRX5uZhN/CNZE
W1/b795jVQVr0UleGp/qRbJL7QmVtFnQ7stDWh0IMhwnEP4SGJwPjietjT4HsVLQDfOzaBWdxBUa
RXgAchlC9tQ6xxv0E1KSkeJkdoZwdqyojgZJ0uk5EvQQWa6OJ/RNZgLbXn2EgennJD+4/eNrIiBg
SGA8HmE7RXWBcoyvCQIFE8pMnHUNuphwIgdANQgkxZincV0FpGx7xf95I5hvzmD1K5drjrpH5d/t
7p9mSKbaJHNy5dN+e1pHuVNl2kKVuNN5FM5NvSEuTraOR4dO/e1IT8uO+fHJCt/4iEHjFRN1kmTx
5d3XcQ9c084faiIgjOnTcLJZEB/O7qdZ/uniieFVAJiosBf6YSuUL8FcZjB64sAk5GLVEgnxrXe/
ZRVjFCnbmZ59x15+R2e3G6uKuQkHCEqzRAD/v+37GASLdket3+KacR0lnTSDpz14tRkJrqG5U3uq
vf6WZAgE6NYWwYtS6K05WrA52MDPssmbLRgCdbwcDnItkJcGNDU45nbxqDMWxLn9GoyqwE9GguUu
dbzC251wid6j1CoiG/KZz52ePVqNXtLruQxRmdM3pnkv53wih2SaNNG/nAPS3KS0EU1x/SanEYrK
8Rus5+qsLzccPGLzogUss3dvHZ+H5cisiX8AyF9Tdund91a+3uqDHOWdOTg1j35xI0MwQNfkMcoY
tFrgS2rwWjoFlb+m2Nhi/s/XFQiuhK+TSy0uoxYt4J2FUYjd7hvkUBmhWNEH8Lbqt7PzNJC+IuiA
mnH8w43jABJ7sVbL/X58wzy69d/sGALWQVBavQ5Hw7cV83Kn5Q80YSl7AwoKd23Rzm3dwoPhxLkt
jxJJnERaH8z9guF9ahgaxpViM8pFzxWeBzSuDKD/ca8a7MCJCu881mWSPxIQkPeR/3gBEDvDU/QD
vM0c2rEbH9fgvWfjg/bVKlrkyz9etl7C0bAACH0O2N/4xBByAHXwxMDK6gdGNs1nYAPSCsqihcBR
PlCeQl4Fmc/0kICksGhYKP/cSxHkJxpbo8GiwYQ4eY85ApH69V0VCCUOOIpcTO+63k2rOnwbeWSt
m4/aWlkXJtB1cNglYOceq5WyO5L040hcUYJmmk7OsqGR9zWAQokh6dosl2iFVD+p8WsmZF+/j0sq
Trvb9+AHxEz1B/eR9PtN+Ir4KF8GYEyw4ExRKDIyKwry1s0JYbx9aVrVzUN9LAUYwWZYS+NQqpqk
djHfVGpJZL1sNHt3e1fNe1/S/z8exTxcnzWllnWzjL65SQ9Y2S0YRJAFCLIRW4PuAGT6LdnDS4Cv
aVcnBt0qMWaV3WTNXjsRwVhakp6NRwIlt6leiDymVOFndFNHTgxbB//V2lN0muavYKo1K7I1KJ8a
4BrDtmAy6CzHI1XbAE3WwWdeu0K6IBnUNAFIeecsO3Z+8al/r+fRy/yeGEtIzeVbvvAI2SmbjJ4f
+1wzq0QtZUPEju5ulykAoVWkcsDsIHdfqYSGbj50tXn25mkqN/OkkQ7hLmVMu3Jy6Jv5NTVTj88e
WnTCaWBT37U3fejjXSoNzjb5akCbFM/1ooZVEWb5lSn7yXOD1XlfS4fsF/Py4icqmKr7ZIL/uCpK
7+7EbJfNud9uIyxr5CyB6MgL/shoYvXZepOqprOs7FIzx7BJf4HrDMu4S2/U3huStRChfJwBE70D
/y8sK5NS0r61CVHm7MDQKQoF+o5uf4r76eWUoh+jNmSqGH3gcP+mmiXb2hl4N+KEzTRMKLkbdI9g
O3YiOd3DY4jxZvF+zfQuHpoJis2iEr2ubOQYZeh36Q2mqd+psJW6iA0XF8mU748W+kasDMkCd9v0
+zo4mVsWq6A4NDKgLr8+OOESjhU68OKkHIEQMLfm2cLlTLNJ1E2R8cKenlrVbzmmMjeZwpfs1nNa
GzG3Hk/ZEntcXABwybFtCb6w62nQYIES6b1N8kyY9fVodVIKVp1loUfNxNXwulTxCcPsdBYmY3fP
K+xC8wvxo3RSGcBGg1bshSxVT247ciWN6nqNkwt+qJn2I9/gNytRsCWnj596KHZHmBqJUqaQRhak
kt/oqeghXRYCRH7b9MYyBALZzFtL0veysmbr/dW65BoG+qo0brnH4OEXVB8vdCmhdMdbufW2Ntzf
Ly0WGL7O3YVAJtI62S3UzRQMf4t1JkJmSaVefJ5vNa/1WkzL46oqCbUcszucOKndUrQNsyusC9dl
8keIgV+jCfVwIyrRCggLLRXRNjiqA5qh0jwpk7z08V+dsYJS4WPlCILdhNiBDDZRgA9xn81dWiKA
3I54PdfWrUkg0UtvWDxkjwexbuJ/RhZ16/znKuULjN8fLOzzC3l6sqzTP473/5JSmO92pIUOC+oQ
ld8zetBnNnk+1F3LBiODi4+pSK/VZY2dUtWLbwV428n6eZ9ctvvYwjYYF6KN
`protect end_protected

