

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VHfaMJ2jDU0R2eAkOntfC5B4/6MobpZ0NSnc7trviKzQU5KHakm896MNUQ/U/XUDUOQl1Ix9hEug
uFcdFGHOlA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jZ28dq+cqatvP/oWT0j+kbhevax+rcvgcOVET6FHORIxsClPAe5EiSXk6mDgtoieHOJgnr3iO4zI
pViSw9QXhHwC7nkjQzCL5GNnIAYREubhi50JKwxrsTofbyKzT/U5b+jDP0girnK+nPIjwrQv3vvD
PHropUlOeQU1eg5rEJo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wyTaR+5BBK3PMm+GuCvq0Bco7y5f/oiFqNMyoEJ+yA7qA21Rc24sV0Xv3v9W4doHSIdeeP0oUNh7
9I5Dbu7bsdY24p4a6rVQlpW5VOJjg7abnoTszev3jaBtBOpAM+FQDIkOj6hl9ZK+eUTOGH08ap1P
3rtu9S06fVXB15p5GUL4qJ+pbX9as7bXZJVw8JMDVFn1WsdJ/zMn5PNvL5qC5jZb/F7Sf9m7DkwY
x8I3vpZz7RsD6/RmMhT4lv1FkcH4MpJegB1J0hL5KoGG72FOKCqONCLsZdmnqz5BmJzgYmphlYZC
jJckdSX4yOLEg+jbosSObzMclIjrm9gORAOhKg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qekQcsRlt2+SE3/eW9XQwKmx/wWWvcG3c3jSLvuGiy4GIetXM6PaXqKAuGTMI8b+mux4A6dEdodI
mIX5ojnf5ZA1jyISA9q0jKtn/LDbiV/JtKzm0pK23fPqh9/IUaTz+oirXN82WQzZFKQ5TKpwrFn6
ZmImSJcOKVgUcM/iG2U=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tlEZl/v6lEdJp5aVMLYyANJmLh8DNrpNnDhyEkIUHbeTfiozIDqQ3eefGpJHd1yUjxDr+M7d69UI
c7u5loKJo9CP6qAEjMhB9NE50dWkO/cRVvdlBQSlpGD8Asrd28oTNAHTTge+6t1TRCmYfvMKOt+b
zBqmGPTyIDG3LI8DiLXNfUjWjl16n5IRikeD/e8FsFJjAF/a0Kjal/N8CzCmRiQPdsZhdMiruSdi
vpIRkNPRNpCK4J6asTfuTemt2JkEkG10IvEYhZ/qTCco9PECc5G9y0loOf9owc6R54o3iALi9D4Q
T0iTW1tROVF1jLbRTIe753z7r02QD4PyC+02yQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24176)
`protect data_block
U5y1kzlmlwv6QzwbC83yQhTr1UM2aqONE3fghqkDrFiTF5+t4Ey0AKjaAYC6R4JFoJOs3wuerLm3
tZJzp9KJypY3C7AphzI+pIT851StoRXztZ4UVUeY3hVt6F+F+hkvyGNxp3VRnf0Ximz4mOmRskbj
4d2YmtncCYdfqQk3prN7sBqyRZPoHLB+n/tBWEiwqM43OqSNdZZmp+9AnptnZOTxUkMJoVjpsm89
YdufVSCA47HqA+0UIMv7IA3usVR0Smul20BSAEt+i6xjpKt/PbHZRNIT3JxGNjzdsMv5/DgYiKYl
+zka29UUllgvGiSasH4nR06jb7Ce7BruOrhP8NL38mJHc71LG965M5R8UXpoUmIEcVWAuCmT4J/V
XTzzcicKkF3AYr0SXd3iAlTEdMHaIpTi3pKHPRKPd4JMAacrIq5SAYH49PEluGRL/nVoyF7h2VXD
hWotE4Zu6PfhE/fGeiiT6jFTdRMcCW9o8kCHumO+kZtv1D8N8ZM9oRxu6g1gXFNGDecG9LrVcrP4
+2eDxYwvuqZtpIMVmaFabAM+vqF+g+IN1qZZUOiBrfPpIM1Og9OGfnu86Qmv52RBvDHFB7o6pEKs
EBTK2ZlJHu9cZhpKDZsdgfJx8EAQzMNxoNclgsSslN0ncpzIlHFdPvLue9KcRHRaxQVAkLYF23wT
7ebZPQHNbXbd+erXxTuEdhWT3aleUq9GzHK75Tt8BynmW02t14/jDQJ5iaTlc5yzHEnaxwOVoz1J
8Od6j/KW1pmBXALKcO756VNj1lPphiOGo2OPu5q4AAy+d5JfRtV0+fDkDj5Pb9N3AV+yjGIlroJw
9rYiSij+x0Ka8eTLRpCNb8chmX2unkuyL6+CrxuuqaA7etPKaEHLeSL/GCxo0gy+6AHCeNvJzEim
1DLcFtPU/Ho80qMrOAUW8H3xaRqGvAEzTlond0NYa/+yGDVfgpfny2gHDniwoEp5st9hLXgE9nzH
fpcTXTJ6vqGSnQNnZ75qPBXFDTL4vaPCqYb9YqcqlNON11PULMR94TtHdtnKOZ5nuDSmI1ZdcOW8
mJ9lKsPiCoVMz+DiXCUU3bVPDQyOFQqMcPhDdCzqkpr5fR0nMXZSnH5mXdaruTdo8wWDFuVrjwMg
UwTEM26fjFUpaImfFMbt3NPoO0gcXeBmCFDhuZGEEqnuS6+JVgerMnxO9HfXju1qYgO1ge7OwXDD
37ouKBT44sII6kKqCU6bmtfowUlChBZuAJL8FB7160wVpRymeHTbtsV+Z7MZasb/UNcDyRL9uMKl
kWVngFCJLnIV+HCXEnIvGuZBBwuRuQg63lTKNtblguW9efzWPdUboI9JZyRFt9Es7x4cur4iu+VM
pQYAjAACSVaeeDPtvd7IwXIDD/mnwm1F+xbkMoFHdlCrqCZEKJspaymLaxwkwi8bc4I3ZQp2uZAz
lbAVilcQzpRQpb0DBnMGZVv2NYcaWWNMVRpNjK/MyEwvZBxYUg+Q3aemTlshcuYAM9XFgREq/elW
+jaJqc8WrJbTvuw8JD/1op0KxY1YnXm6RxLfw7f2LExSV2GHu3diesZASZyBwTJhZtH7CwDfy69N
XyfxA2ZlHXFEJ2JQ2jDUF9+UyGEWVB7QKgPdWCBw2Bnsku7BPwuHzJfXU8PPGPhAvQ0v/eSeWJvJ
zXWLw+zBIcwPaXptU8uWKaZQ+liEfWEaXKWo6IuHfml+vbhNK1Dhp21f8N0EhPz+08wfIq2Si5yo
3TeTew1lfpYzPrnYQV6j9a1YK5EhIKMjGGDlVCU/jlGS6nOHsh4EDwWdzPy58FNJqcvfTcp/VgpI
XYzOSIWw8AbnckNk6MpP+pO4tYF4nBnPD+ZiNs31tg3Lj8AsdAdMwfN6rfzW93vNloIJn5KmmlH3
DeNkwNPnROri9xa+aNKk3PyEtgtqgpUsd+2gAyOdjH8jhVQ/p+zWh7SD51MQfqJihvHZtaODXQAy
Z1foUlUvXg+KSHGTPloeaOz+RyRtvtM2Wrw0CyaPTCMv/JZaT+b+csasYmIqvz/8n0PAFcD89U8k
6i3JKhwUhxUArknuPaNgYFUEwUOQ8QVweXPT+O/16M9PzQ56UJ1NBXlt406dQyXF/LDiNWk+F87E
Jp8nzc76R3hPHqEXlLRLw9pl+iVr60cXcjn3jJV0YQnfCrimbA8psuwCJBNu0llxO5ktiBjIR3a4
kdbXAE0dppvZ5/7b5q7qv3cXPTt1kAXoqTwu0HnZPTlFBxvDP56JsHarV9tKw/eQgu0NOA6bZ3Zv
IE0u9qVPoIMoKkfQYbdbKiZHjHznBiD9cn0DPMUtDSdFxN0oZi6WuHZ59r/pgPhgHhs0v0oJFAWp
tO0vf3bgicQBysvi24XJmSYWSMkkVLgG36h4Qo42LTgyZtOrbzIr5quGi6Qb5/ZrWhKAKz3G5Wrn
fC1U1tLAZmotzzBJcKwd6qV7iqIqbZrE6p2xyzN75skUfW4kwJuWqzOuIw+LWLa+f76W1IjpiuDw
PDPBJ2KwrJeY5LhQk0wuDWR6OyRklu0E48oKWBzVtgYAGx9s0BdNDVEGAKuPozUez0+X1FO1bbo0
i5/PgNm9qGsZmFvB1hJYxy4u7wRVBeHDMXZg/JBRLlRvN6t+Z/75theN0gznsFvHS5is3LUMRFwO
qhDTDCB7Mye4QgUJqsXgl0iGTEXD2avN2+uK2cAluBvSWiJAriL39uplhBmR9/sxboy8SG+S+aZw
kNddsLsgwoqaCym1pDaURT2k3ts3POXJi8B6EXQv0VUYOoFcBFxXKYV0wwAdT6Sz9fSLWQDsTK4z
3DmD+sM+f7Pt69ZOZ1H3b6yfpdNBSSqzSaqPdqoyblY1OwtQYBtn6jc16biu00fpaNPhiPwAaBXl
q6snc0sQMWegpx3DEns5BUrRnAxvmk3H7vP8kb9nf0XndLzclZpnpNLctZ+SZy65dhdg9+7e4t8/
5jKeTQ1x3aq712gX954izy73MUyNL2ySd2Tv4cnlCooc1lxvUIXc2eaidsZroWD9d9QjLPIoxaeh
wZnvCjzt6woFMu3TDR/fggf9b8Y8gEkawKJFz8sVdiFOnXsAtleSM79Y13Z20nxJ2RfQ4ofrt1m8
jYwfHtGU/OtYoglqFX/rOfq1/Xspm+jnmTJVGgKQpWeIAu/hgUZp/AzDYpr+mW7MFApHo2WF/hfk
qOJNDaCUp1GVMNwxShXrvTZDWl/bxou2gGDQU4s0yZO9hJIHuSxxNt2as4vvUk/Gm9DqqdzS37Rg
J1QbU/BcpiwnAfHIqoq6LkRci8uxSNbT2rjzSpFXoR9rX6xTU+t5LQXmCAF05zY3wcYJmzJsbe5R
HXElqWzirxodFBYQRKn7+H0QimSqcFGTcpJ+o1D26WOzm8vyvdsmN8ffmltX3bPfc0u1pRWTuvnf
MJIJ9l4PurtAztYS57NktKnaZaIowbKW2uW71AffvOWfmlkysVSn52kQoKnSRzm5y7HuUGo7YOmf
p82rBED1LYOPMebhJXMRP2patnKLEnhMo3vPZQ2nD1v+eNDx6c3GeQy7nyxpFawr8dlvfyB/pHV9
5d6DJBfjVpL/l+SeXmrGFBIyKZw8kXr6JXI4AI/mq3Ur1GAmg+NZsA3QH08AxYfu0uFTpbl8DxTS
5NEa+K3wmhJ51+8S6oXRSbGlB71CbiKGgj0nP2ESQ0QddqBtumMZubk0jQ/INUq1pRnVDl5b1MgE
Y1c40jAXCRbExnk01wSwuEKBEjlietVpsM8hPiGFfgGuKAKZs720JiCkD0goA6tPQJ9NFdGm/fDQ
aY9G4FOqA6//xfKl2cH9aVSbHzry6vmCHUsiOgpdcgQErKf+CEdykosnIN5CtwKr4VCUPcXCvV/q
o/xELxVpDzq+UDfa2RtK/VCuZ3u48TTr20YI8f1m7i8+LOVFvZ7MZ2kPzD+3MsN3aJPeVsPjUdAi
q1CpaPN8VV5jKy9x5u3BREtioylQnFYoXHukdhvv2YEQtCLd7gYEljYWrz8lg7Feffc498m8Bkx6
f/fje4VhgmdU/ip8m80vm3qxsAsjfNEZcEqWKh9a3RB8M+GOTV9K06Z7F2Rzq8ZhAHJAaURqVhtC
ru0tcGAMCVNm9NVMYHBYIvy1zli7TCjYZIuJKcvnByUIL5A4CVD1nwaX8DCAbgOtbJNKR2yu7S+t
drz3r8qoS8F89GJAmUN+ZGTgNnEUmnDSfafhW+SfJehrSc8v2Pur/dgtttJNsaCSxekXkmDBI7/M
hW1sP5QdDQOQP8VFKvECEZPutGH0HaO+igOUwh2ZqIOKhcSH6jD56fGw+ULsVd1QhHzi3G4Q/s4H
o5OjtrYUMxjCHIuWaL17K4IvmXasuSo2z3BB80jL/HAMCxxxNLl1fZHGFx9NKSKaWK2NNgCXVg8O
Zf/BTUu0S4X0UkDdqK3OjRHzEbpUcurzbD3EDYVPN59vaxb8j84+2zrqSWfmblYR5G8jbZojCqfz
V3q0bWcgHNN02tnnK012uet1KjKTHXv6zQ+oNV6p/gdG0s2cUgEHufLrRDSLaCHH/wT7SnyImIKs
lC4kV7iQ0t5RbS+rLV4fJO3qTtKTKUhT+ayZKEuCaVHRX+kp6QSREr1LLqZxEuvog8f4N2i0ZbXy
2c6RWuM0v6HD7TE4VATHFMQRTcWMARHwSO7Lxp/AfTDyq/Dh2xBuFX9uMMwlorsrYc9XmoqlBoXS
ljIXh3nwrrWiDkPgF2vyxKvIjUF+zygLNW80JmkZBghoOGcDjTW6hZ7K4CtVyUOmP4xnfAp+CpCV
b/a1WP/0H95HxHNTlz2dgbKfaLBGFDhaqSgTjpPqC52oL14l03RzmYkHQZk+iXliDf4KbamcpOme
CZzMmEQ6zSWHNDP5IZR75MDEO2obtTZgoYJ7ut/DqLldnmPX201JwyjLqImc0V/QoNv3qeuKxcnD
SbLYmLfQeE48RhpKfobdkcto6OJFEZbga8nwh/bPbC++5ayDHpDtsq/kZaVNvFWyk7KDSI//kvBx
8qGCBPBQpSWbz6QDVe2PKGXK5COQ8KLTYFVGc3L9EDqFkh7Eul34iZ9tYwm0ut3vtX/Nw09Uj46k
ilBJbsqxviKcuQoGbkG3rzWRRVx5QAe/6iuw+2sKwNXhIF9L0Y7qy3clpSSG4kpTO8BTKQIM2Ucc
laK839PjlpYQYiHcextjzM2+ilpY1P1Gn/p6IJ8fpYXwz+Zkx4yEqK0cpSrlLMXLqmLI3jxRuoCM
I8N3YWKuX4hO844UK9/YVPBO6DrW69LXV4a7jPdqlcdh29YDmJznkxePmAFyZs1DFsKGDWKYIEXf
fuwuJobAAQ5jL8SsTVxW29vH6btQm9He6vTNAKbvZzuL1gou7PoXWmZmIVLye59qVGCKAlvqb1n6
wbn8xfkePPT9hKgBrMOhigU/d21DY6Z+I8LGTFo3jlm+8XnSuFZ+FXTVZQphqOsU5G+72v5sF9D9
etxoZ1CJjEz7v0BGoRjpc2HNRI9d0vdHzLy9g98NfezjCAYKuhxIWZ82bEDQqZyGyHXXPSc8uy/n
agrznjacgfP8GAb6aUitpS5zqRwLdXFVeIrICVKjF8h/uwyy0da7ArLZvipr+WqArhvekHncIYaT
4DXB2GoMvn0gkjz4itkHZm7vIQKAoftSA8SJCinkAY2UAMc/EgyGqmHDguATyAHjlg/r4uEFJo7j
gCWtHfbxACoQq+hcO80GrjSZowHAofva+SyoMv2KXE20e2OxUt91GmTo/ODxeAzjg9vdJZb1Lw16
W+9a/lNGzyBD24nBcUYO33NzN2xAHAkmQxgt4jdDXi3E8DRXTxCEJQjdrdYoDXEbW2Pac7ZCkA6n
udfRXs2bsl3HVoOZOa/UHtax0mUoH/G7xPEptGj5hWLfq7kyMbrGxiGNiudo4ziteCzGMjKyD3Sg
vvMhUZj387NDIGKeT8ytkYgH1ITQAzr4jQ1R9gUN+HMxquhKwrIFoANYsgeZG9Ax4q8536ainPN8
i4tOkzUJOaeC3KrTtVguGUUmCStG99v9q+tZvg3BMyB2b/h0sScVoztkXghbt5TsFKdxYA5pTubX
xyu4vZALrqz604ISfFgFsVpZdzI9ZcgKla/DVXGQlJ/7m3okLW955WIQJNn0vI879b4f/uTPWGlh
aOhkB9FfG5iD4QK8Eb9I5dckOZqTb2DkYx5zvJr538SMXlpRcsh23+vT26GPWZsnnSIvAXFF5Qrq
LYjG6oiY9fmMPy3jASGb1qnGT5ioJVsACpVpN/3yiMwTjZ3UV1vbRDYp3USO9jpZrKC7HBy6ReRO
J2VXXzZTRqdl0l3oFpX4z/rh8yWFeIysbdGGairLYZkDUAJ8GkAhr5bp03AweqDjnYcQj21R+Y8f
ZS4Enm4Nu91jSMypK9rYiwBgadpwK2agPikfqdyWMSyJwBl69W17QS8d7e4pugsFghdZL99w6oe/
fGKuM/sNsA+MeIEpDv+WSiyzEXTPad//XXVROHK3FP03XsH+W+x+BijHR0EejWG0RrORxSRM8tnb
kwjLEN6li4qLx6BTTHbZJpsm50+1BUsTZbXBR7zMny5kiohKo9Qi4YVQNsXy6EGDeR7XeRBVc/bs
aAD288n/nuBDkKjhCfw7RMbWi9MKb8/gh7ROLCoQxYuLnln14u7n/dDqkDsFgOROp679DJkpdWGB
3QeT7p32Iy2Q6SGN7aGj/ThuphYeyBR4iDHoExrSZxP1TVTNbLR9GGYNQTQkUW4vr2pizI6ziFo0
x515M+Oe8Rn7jEATZfEI/w3GNUqS9bDpM2KuSk9BAnFCw2Q15et6kuqkcHSP3PdydzFP3qaf0EGu
k6W9ysBCz9PX+ohUf/2N0MVpKXEcIb/VkjPizOtnpXBXycWRFDAn3Ne1skAFvjX8WJrzbb9NaIkY
sUWNCjHgzgoHCmXYl0rTN1uPqPC92dstL7uE82+MVxZ78PnOMAgcYxNYslbJQf+eSQkq9dBYtYGM
T77xgayd4jKC+8hjG4fSr5YymbnrkgTEPw/lDrRLf+wBr8SsM/MPPUbAvEqMnKy+tFw323FIDyDk
ft/mZWgkSmSCbzcTSNlbrhgwxd10/v03NZ2j+fl8KT6yOMjlKAKO2PpgEDllQLd2yIMDrahpxFM4
l1U1B5BLC4DB1sL5/d3XxnEK3yXFG9NRR3INx/BO9E8F15PYqtOdcMLmmEr6x8eyPuo1Dw/WJYye
Yp1xzpR140p3em9oudl8TZu8EHW+/RCz+kv35HEMly5VBnwt35CPk37DDaM3lXzn/ptlRTHlbiOK
MdrNuCxOwKwI9JTkD6ZhkhzVolHfSrB8Flv7Lv+WfkVqFzw8zpaX75wvYD1IFrBb9feHlhk/Vhvm
NI4YS5/Vbr8xNOIZOjjHuDXU3XZF/rAvNQ164if0Pelv8fBWSBJiFt0y/kI/Duzvz6izXxl9XuiE
uqZ70UMVUpRiZPVaGyPAXHh3IOZJtMHfin/JsC/rb3PtoWeUZ7aGtd2psv8zumYoWOD3P1Lbf/kN
NHSvwUTemTYEzbo73QYZjAYP1jPBmmXT9gRnDq24CPgBACYS5+FqZXiWjnkixtUQQ/A3/fDaI1h4
3N3rvIoU4b0s8Is1Fjd+zJzYQgzgTop5Be4EO9OFYCz8ADj6E5ihF9yvF8Gm0CCRkmmL7k8W/YZg
oljO9B1R8XdG2i6qP5grdKg0piIntklB6Udqk/vtNXG1FDX0MIl6U+qjfFzlP7sE7UWkqGGGzL67
y5wGTMjb4aVsuI4KNI3h/HgfwvPVpch9aRaLOPjoE4ZipiId8WDMWzk0mKnLtzezWdxmj7/39Tmk
a/CknTVWTmApTgwLqFPhOb8i5/4ofQJ6hxfKwiCMexMM4Efdfk80rchXjhRqijmwOKxw7rMRYKpF
FxPP/iiVf6478jgycptd4dNCvQg0HWu1RVsgnRzC59zPwq4K/1ERnkKYRqHb+U+rm0vI/6qrA66V
7GTGbXZFfHNwM4vZrLbI23rsFkta0YiWOsW16tJhOmAXBCmcN9u0me18qA3DfHf0lqdKkDNgOge9
sqUp01GKRp8m5DFmbk3LMKwnN5wjIwGZ0j8kcdrEQIBhjKn7K7qWjs7KmwYx7mdYb/XGqLxjQBVz
lxuGr6H9F7ke1r2hAney2qjTSGQm9c6zU7G/IEMCPXaiv23AteEspdfgAql8eT8+TppFFNpJ4p+8
J2/DCC9xn0kGwi21hFdjDnFtWCzWc0DqSL2x2RdpIo6wPNuog6+e6NljOsk7hQu26i3p+11y3Qow
ANe5pKKw+bHzSPorMIw0IAPY+d57iC6Vys526ibWvJDM3MGqxpK8ebKhUC5Y4PFaA/44JRGQucYr
KA91Zies0udxhSpQxomDt8+Sz8/yo3OKpownxABrJsko1t4P8tThG9jeiC1VWbDK875BLbLI6qWo
E05UEWg9piD02A5XFilTTKMfNV18AniAGSePwVs3zVdnw6xddWNrK79YwL2vem8XzRjgzmMfb9Yq
HKd04oZOOHLIm7tsLzGY//bvbk1li8MC3+/2/hIGyvt+n/3IxZkVNNy0kFO8Uul294taT7h5ZR2j
lX7o1d0b93yihbWajWRUxJE4PlxmrICul9txSVfn74uK49uVgTMYcoIQRn45NSDp6CnDRUNFLZ6g
MVPTvrx+lZeMkhrWEX5FXgdF6+yyfYKbfwGyrhXIEDotahZTyv06RvaWPOjjP4zGnj72WscCGIf9
1cjWdeV//c5V+7HcNxIlxQJNOqZhgTgOeL02oItuNA/KRc1m2efY5GDCyijezVja6T7m3VMwu3yg
pIXoMqifK5s+drW1xNynllB06V9cyPk5w/WXBxyfAhLkm9SUT1CNLIZxl/YyA20g040vyZV0QBJZ
VGMOtTUC9RJxdH97H47JfToEk2X0R94E/BzsPysp9b9tGdY4fXgiO3aqLgxjPx3ssOhRqBz19chH
JyBNRMHpN6EZvj2CC9xM0BKS3N3x4UdUZaqOO4w+/h2Kt4FL0RDZO6mNojbVJd2fYxd7U19oMd6X
CQOHc8qdU8d5duTuxMR+Pzb3hDqzAv0BrHlbF6rLk9xXF5p3INI6Nz3Kf6WC6rlGg+q3fw0GytMj
SfDKxRrcDmYFkreVzjLqmalK80Hm9A9qfM0hYUdkLCDxrkQeEuto5reZoGHNZxKrIwQG29YefGnw
mpz2lH9N6ghJI1wNt+nlVNPkFzeMKou8k293WvOAQiL/ktd6G8TWNRRogzkGQkCSD049PMCdsA9T
ydfjvvZW8qh1yriaGTwQt/q69iBeWeJvtOPyiJCkyg+8jimwEMLuEZ7r2N3eD0ykBs6u3rTzcu7R
ITYAoCRgTy58QEiuiFgcabaS/fZZry8EaTHXj4+F87bncqNYdol+ebYszITZN4uyPfJ9uG4TDSkr
vzoxXIWew+01ETQD9xfK94ZGdb0oowDVFp52RvU4BOjIXYdvb9tAmt+ailit6OinzDa7FsuijfhF
SEPaPkdJ8nKV7bAzJ1ysBJkk3mRUio0VuS1O9gX7OaRZUcG1UnwRTa2DdVz0HmSuADGsgolb/78D
zZkJO43QMXYCuEuNCP/YemFE5KGNNdWVFLwmK1yV1gO0Z9pB/nu+phIZGfxRdxc/3ClZHvZ0tR8o
gHwh29Zt81qrTWMjavPMXtqFiGSzPqE05kXkWlPXUU9DT045+OkBiUStfW0dwKwqm4MlKKUPpd25
Lw8JkyBA30OArzzN+9gj5IWBvwfqSgQ6Zz4iOkDliuQAbZzEiOsyI8sSTL+9HZW2PJu/lN05VYT2
dcW+HaRtNqOsWDQEtntmMaGmyZWMzNmYMXpwmZCWlj0S2ET7dt5zCGbkotV+S2oHxp+8CYTr6AIB
qqFkpv3LvduEKMrRfRd1Mdi5qwRnQ0+Buiq/PEtMAhYyZ8DbSd2FTyX4daKClL3FwSD800123LJu
IETw0yx+jXsn80XMI7VhFH1UdvIHp1tW1UEqh3igD+2gwKtRXoDNlPddFJr3tIK1skljx3u8DCE4
Xh1kYzSVfaNJjNFDB5o59KDAWlUF+ikPjB2OXIDRm0f/UuSdt1cCFKkNVEapBFHu4TWr5aqYyno7
uNDILDsK3NOISzYhRwmOoIcQptVe73DEfArk8FLJoSHjpTY5QBHV8802R5JGeEAb+bGu14T1Uvfy
JGkn6bMPbUHpUKRU/R1/1GJAvV0KuAqzQRrTYnKpmz7F30Q4KSTJyHnxwwZaAu7QDMD3Hjkb7erm
duEGJTHfRdxcTVkLgOqKJCxM9bNbV3eBlBV9ESNgnSli7B4jKUh12dXQJx13mq9zqTQVxgfDow/A
VP9uTYcioJIQfnA1opH+1U9lAXXbL6GserSHXDCFcS30ICi9mE/hBargKN2B85IJsj5wjSvYTeQj
edZejj1DtRdwtNz0LYU+S9iYRFN/g2xkCb80SHxjHj5c63GDUH91DYbtT2YMWrBgVnMHxYnjaiTx
wMjxdqr1SdwUKFYvrz76ZMjTa6Wnhuk4kr8o3VpqWPKwjTezCVCUMfy8Ry8IsEvLB7oLPuzQpKzD
PpGI7jCFOqfbKNepvNmF7/1DKTs9VkUhs+f/8f0VaTfh9j0b9ABtrgyysMroDnIWRKDl69/3WIvD
8yZ808po9Frsjcm9QUg1oTdCF5RMGQHvpuXKFPLO7WQSw6nqXUEvEfKhlPIIiLMmP5Dlm8tVCBaP
VFf6u1U17nGKy8v+3MrLvefYnkZF7DJOSSbuSDu0zBSCzmX6iT6ZQqIzKRupOVu9hsELhge+xAmo
JWrY8ZgaWIBLl/41nI+fhiFAb2E2sPJS1/rsw1k5YOaLnHREVk2CO2Zr4aVjSEIjYzz98noa4Dia
7FvtutVBqQElmBP7jdEamT5tw4DZubZA1IKeCkDDfwwAuZ+Yso9e/G8F/c603xMI/ueuakX7Q3wp
PHV7oFMVJML5eAKlvuReH5X3tX+cIV3K28T5HAwIyPZ9B+CeiRdDicCip8pkCHVTkqPqB2EzsEC9
cUQHlaGcmL47GuCp37uwN5Nkqy2E2rbkbLvpAMo9hw73jPIpz1F4fMI6f1lA4jNPOQacCGVJbuSo
ej2qDDfLThzttyFDI/wh+8uwaUTYBZcsWF/PxZ/j3BdJhFUwtDq+Z3UPz8zIPJbudI7kjeYTTmA3
sJUqu0drT6lrK6vM/1UdBSLTqwdSJ3/dKejcEc0wH5ltZG/ZFLC5BgIv5r6UubK+q+3+LSN3vBNl
dlHxLwMJkF2qiqe+C+oM5mnvk+3hi1PbXQ+towsd0UMqOB8i24QA1xuj4ITOd9LkmOTI89SmIE+T
e+FHEEUtkWgpdo2eNCwkSYN+xOr3QqYW6NwT3L7PsMwRrSX+h+uBnmSvFBTF/RKa0qfO6y2Iqxc9
vt3nHffFUz+OJVbz/7LAUDwxeoXGhBF4ryGegZTdRmZNm3BYonQyz07tTYnC+B/5kRXB7B69T42D
ztqudvT7xWfrq3bT+IW6rsZXh+3FEjP2URT/V/8+pSEB3rJrxR/d3FUwR4YkT2DJcH0SWsDOQkQ8
4r0yf07iQLNRC8DP0nZNu+QPS6XSrm90c7qRuoOn3RCPW+kG4uYz381O3guS64YrcogRVlHt988c
JXzZgWY/GYd82es1KAOIAGXdK2G1b3hiprMjpUg7Ol4W+lNnrj/+VdNzBDUUmXP7ckrgsM1LpgvE
n7XOhmOrKuOgFwY+4jPu4+CmqMqaTCmxWX9wRmTkNMH6rzmleZv/jr1Ckndokz8ITkHCcKKjzZxO
khUb2d0vIs09fbP1xlqwNykNhV4hlgd2ZBsKTUNnaZaNuHDBdcJW3NcwbyFyetbwphPLoCbM89rs
UVoK5t4CSkN9K0+9BO0Jjm/Yy3Lfb0K15D93PyaS1NyQzvbPcjsN55DqzgqA8irZhjQkB1bFoIQK
YMIURELV7FZLmr2m7T2PT3yyyC4ZziNEMW0XmZoxZRLTRTibadlhO5XI4oq8+SVB1MK76JRCJIQr
4s4bFKMxvP6/Ghugzz8kFMS3mXvUYrf61jKdX7Oeh8/l7qn5ItZbPKYl09s1Y0A6XP634574at5x
ASgCmCSggJX/Vmt3iIE7oABmkQnzrYMlu10lf4+Cu2bT23Ng5wP0m0+4bjvbOUIQIcbQzAr7Y0uQ
L441X1dKHJ1gTZnN+vE9NswlLa32qGsv/78AIlvEZZsCC9xnppR9Ajkgu0ZUTpBPMAmh5paMZuQb
vGWrNEeSvSGVcG92BMhmMhnVdEe2PZp7cWxIKa7u35mgKFzcHVc3zoVLsXmNWlpeArONDzxGGfmY
msBQjqXsEM1mz4G9xffL8mEyKRiLRXbMadePMCqsaRQb8tZ9Eht7yjz4g+xiG9hmM0D9od6nPX9V
R1phIMfEm518fhInXYaJ763pvlAf7f8A6cTSMLYJVodSAEs9hwwv19bcLAkhp9CEk/2KSlyKpc3u
UJTGj8RKiht3YW/kU3R2jbGHg/LR0kfAL4KKZQxIZSPnUZVOfskSS0edN6hl/1R/uSeFPT/jYh5D
0NCB5nv3HJuEIz660Emxp0M9wFPj33Ge0P0UXmOfs35SCU1e7pRxhxT2sEpbudaQmDjhNv+OwhyL
CVPf2bapXD37kvM4iRssQ6tMHh4wQWH+kP8izOOz+vv+hacCr1b/2GyDdWRaCwuc3vrRlgSHStCQ
zuaN2MBTp8pDRpSrvVJ4/ApySiGmLmh3GEZhfgeg4hZvZzU1zmh4Kh7pMNyHbWv/XeeJQxpWiVQc
ZF3SRESWuTciBYRbNr5gsnxvXRODKEDwRlIneTo4buos6hlAhan6O3MqSh/AmixgSQf8xVFLOe6W
80KcZ83qCZLx2dbpRp1khSda36jz8OcnkFzvibu2tCbaSTXXQvCr1FTI8iy6bt1ywyCr4WN36dK4
ogpUVWKme4E2AQpZSAZaQlBAvwbU3wTAO9Jg2xvMyJdnb+qVG7c/1vXjINoKqggz79noUtjA+Kq4
JR4+BAQ/EhQSwFV0VcP5ohWJaJliSxbuyTdVBum4QV5Gzr6VNEZr2JKxFXbsffed6FKW+vvaQGEV
e2p5xxavZbmvcUfwXZADyRSD9e9GPX47UTGHpNB8oHtdLEd9rKrIHBZFGggVxVGwiE2xK9quAcKL
Fk6h/9usT0nTXkc9VKcbBntijjYrK8tN3rzwVcmYb7gThzouJaJDR66HaG9Qi+tpdhgP8djSU4OW
beoHKLZ5NRcF9WKdJFuhtA3Rpyc8f/WPnA3NrQ3K4yqOJ3I/xOyfYeGwamlQPPrFEnfA16V0dBAA
M+WIDqg2lMMvMM1x+DOy3S7gxr//nqM3ZuLt5q1LaBjg5pU1fXbYNbMl4RvckBTbmN+vQ1Y9pKwd
XjmzAB1SKvz/EUlwDU9o3aidIkbKJdVMYC8+iPEy8cT+4PqLZyBP/NcX/I83Dp5qarLKUf119LXo
ggV524h8MNlwUrBclU67xqhMigsrjSrapKzxEp5j+7NaieVstzxCOOgtln7Ob0f9KgFXrET4M0Vi
YVJ88WIZJ+1Y8G/AfxTddrY6zL17joxaAm7fBGqa60puGWpq6KicWqorIUWSP+ncRdOWWlSmuuCV
2iZLMeoYuUeEoe/cAcml15A5FFcdqOcje/IwfdhtFLIaYKYcpFD7kpVzA+sGKNyLrqb4kpCtzlyQ
HwiBSn6FmfJa4m+QLnCwOYqVcFuSt6Jg3hmoMC1lHRjfwYSfi/HYce98JbGIEt5TSrLYhwyjz9Xv
ptG3BpJhzzZi1YXXwPoM3+pTAsCyjihGVrEYrGc5BXls6Rb1sOzNK3ow7BZrkuLDTfTfal57p2Eq
la0mnDm3giRBL4vHATmBL15XtyZMZNbEUf5AZaNDSr234hxCr4iNrzi4Du84/1wE36cdIbOnjgoE
xUs5R+U/ptf2YYgJluwt/IZvo7pWGIddOEesXJYxmHxxP9FUk+mzB0+divhjMz9WovjM5NlC+3YY
84imcr+eluEE0DFhMInPUiw+RxzS2QCd3jUPwmsORJCsjwCBpzmqu3sfjGJRuK3V3apUtJJmz2py
eO/pjM9PmVBf2DlmBNQGcmi5UWuRh76y6up9RSSQSTiBc0En9v//Gj5+VaspphH8fYzoayTxotf6
AWI1yEAyOMwQI117NQp1qcY25PLoCWK1Cn3zw/3Cx69oqUNa6ChWa6g//Pq1l9IVggto5BlQJj7X
3TBp2+FseY/mRx4tTjt4Q7h3uRFHQr1zPqyBRcAuDu+MsQKkvqcNriSzRx/IXBmjuUKcpRbdGgfs
Ov9r0alqp8gUxsskJWB4fG53XK5Jd6M2q3xqK9VErMp7LuzvryyedCLR9tbvMVkJHX13WfIaRjXq
HFj+5vqGVZUAQWYSqwURk9F4/dfccGntKmQhAtwDLMej1bHeS3hVX5Y3ow+1894b80eKIiSpJovY
Qyezz5TialWTPdg7bqFgO13lDWoBxwXM3vfReaI4925Go9qbJ3MmwLa9Nm2O+IPa8g6ZSjXIT1go
4PYbbiNEm4bUNAgCQPi25QyD1DJLAsBHOiPfiri7+T0T6NtxqPinYW0Yy54Msme546Pd3NbqnZ3P
D6DccSpT2GlGtIfRduDPUNZjhi/jzKXk58KN3kKt4BLZMmAMdSz4x2mVq7/KOsRxSr2EaGtNyUXO
XVcBNAQcJIAGYHbsLsjkX4+sHPK9+ZXCfsF7+Asela+7iPxokRegiMfG3eCIPqJHmlTukTVp17Wk
IU2lnIp2VFHe8b044qCYeujfHaJZVl/dxTimREsRLtedfmjD9rRBqS0XGhU6ow6/UCSlUL7fLIo6
99f2//xIW68+r2EiU/Ed+jAUVER2kXU1wlj713r8rGBQlF6C54tBUcesCf2j3zzB49xJPEujvGn5
gSKNEExfk2aolUWkCsDEyiWCDF9m5rjUg9dVqCxP+AgehfJ1JW8d3QubJt9tAACizjiygXCmkPjF
gleJxzq2UJTGsuiyVtyIKbKoTTJdCpOemyZGkwaCk31x3BncYu5y22eGCpuuFDKRJtGb0C+/njuc
cqUW5NbjbeDvJhnBYmrM02F/MCD/TpUel3zHbPfKI/oCMMSkwAZOP7E/tH4C4/5F2FkKXFSw18pn
i507S5Tk5OqyQDtvjpKiosheMjMaHyxjrU3n1JAFPubXMKgJJ+s+SRQXNqKEhFdj7qLECEejAALF
hcvJ83k/Zx/hBWRJydDLD0r4EnjlDjWBgOSOSHn4mvTomck7RdZXT3zUbv/0iTjTRF5thvMKnptp
Y4u2rkTuqAPzwtT8fWFMeyI09KJWax0V5Knu/PZVj7G16lKdbcrDC/W14SVlYs8w7naGO66jnNVT
YeDCUJrGGaU4Jaz41VrH8YKIVI6dFax9onVkh9DKdMmOIKuvoKGYwVIxhT0UhQWRXARH05LKrhXy
KpW6ysqc4SmMr82qsjNWEx6Sah/15yWbimw0bv9kQ339zlN3FGbLlsEUIaic0kK4rddtXunWPwE8
Um3rGEYqVTW2+4am0R8OLNrit5kYlovlCcT1aTGXpK8h2vOlBOIAf6iJmsjcDgBp01mADMeaY06o
RilBel8CIxf0VHecTrmadqeAGLwx4jclTfYCG2oMz9n6pjztHbcZpycjXdkDsR/VFb9fYKkvMDaF
p7aEmQBej/V1regUTsNV4R26nwc7tzlDxD57N5A5X5n9e+OzkLKXX97gJO00Upea7SWkRW1HcjLr
cNKyUE9wQTTC9BvhnRuSEXViy2zWwvggEFM53A2RtwGHQGmmRTxIEnKWAOxohFro/4afXtBV2rL0
LiJtOmpGGfW97lOH4iPaBS+f2xEa4kjAu2GFAJ1W3q153bvIJyrDRwDGvZX909dCcGugfc/CdQkm
sCg0V7/RRuwPsNopo4r8oFEHyNeZoUBxjKklv6dAh1WTRsqsOKkno+PCfK8Q/bnafqvK8fqL/Gvk
aYXUhKWE64gKBuUO8WhFPJA+pwQ5Wr1OrOkdwdnwTqqgLPPZ5N9ZoOmvYYiK6Kx4RA4FaidlePG2
m5uywGuXt4qSP2CD/YhMfJ3SZWZfxavF5oX1aUCjNQy3YE8oJiL7yIFi/4YYEMo5ENCY26aBpMrD
r43jU0uWHFAkO9mpw3G7BoPPEy/OhssGppyT4JjGlr59euuTA85P7ihxOa3I47QN6ajsxMjV8TRp
xjwUg3DxVe4GxyEU9JNithCqhrn91uRZSUzQsQ9qUHqUzoGetpoUfkevTtm1lXKLkKwlBg5N6XNf
42rEP4oLN349QjonHeDwS1OItzKJoUtW53Cl6WizwalQ5aYicH/H7gWKJPZirOBSYAWt/bEXip7U
7l/97FaKFNY8wck48CUGwIzckoN9GAeGk0Pc4dFDDiFqUSZLKsaFL5nyX+5UXB7VDw/Da8VSOgIO
B0YGv+k4LWW6jCdLj3Mfo+FrIDwddB0ESWuqDRyKrrviIzGh+Wyl3UVGwO7uq3/IWiIukt0BGJOM
Y5XF2q6q8O5Knkvymmi8KOYUbn0LgAJYu9y7jnBCwUVN5XHvDp+DUd2383qYzk0VEmSC/DW8oC8U
knDACJMx+/amMSX1ezT8scBrNjwwW9uoXBT55zAkXhjz1OrxJQpB4Eo0gcXVhvV4ftjFu0Hc4zF0
HQdPATckvLYM+xFVy1hx+ag61fy5IyjTJz9KtcJkL9iWaA67pTQrzAXtB3qFRnaPOfmNVrF+itMI
pDvZa6wZ2kfKY/+xTQb+7HdNlETeP34SackSErvyUyAt2SmUh0jHWCJ09OvrtwMYXhaF1NT6zpnF
qAQek1UOL1N6PiYHUE9hXg9PifDbYB+aTxeDAlliaAWqwzwrQxWweZbdnhbj3hRg8PxK/OC7aKiC
rxjRr3Ccat7/yD0fXDhe5nt6O//7Bn2L2FsqBOXi4PI4biq6aejep/dT7TwbnZt5/6tuN1YahWVk
iz2wS5bqgLy9qOIoRC+RXypK3OWjrbvg6hiVJ3/YDQC5h+0atNpycN279Fdrqf9iXjy8VP6EHpaM
GYLkEtN5FRhAa9k4729VcqCBm0++405dON5dgDbrwzuq73R3drag+hIKjHfQWe18q4loGBgbyrx+
Ef5Q5iRKNQ3w4VnUgZ8x7eQxbvcfE9n1xle2nm8HgN8oAJ9fETaX9kW8hQXOoi+BbB3o+gh2UG0z
TyJ7xuWu4f9FO74mPJp2pyEJxJxqpOHAbL8+xlRWi3ackkBvgSYrQbxTIr9HJXbkD8NlrFRU5bVx
TkGH/E5GS7iBKLAgozl4yi7ATFkLOEmuaGO/CTkFWwGEAow+r2yGwtpf4smJM+J8kRE6L2upKEj1
OBHeVk6j6KSdpiBgh6g6FH1iFdeAPVAq95aDCA5skVjrBbF5aTN5OUdZtqC5cK0FqP0gy6MazIwf
Vd5QJ7Mu8JGqHHSruRlFvI2k9LDUv7NX+fjnVjrK9rzT82t/TL7X46gaRoHL6zqAeB+nI32/P1eI
5KMq3r1ZGSqVdtBRihD3yqAtZoOqjcxret0zd9Z7MTNjEtzfw+VcDdTNNzpeXZ2VPuEtp/9BL85c
UrySoGvs0AoewMpLUuG99kPyVgbtkhLRcQD66A+kNtLnjIfulCHNRQQn7Wb8kVfgbr4HxjkEohha
Oa//Bmp/M6oI/H5ocsBfGOgeTJofwm3CbmWigiEPg3j9lM4YspErVKofipngI5DogrtWn+x9ZgyJ
PK8B6ok20rnDDStrrvb/WLoLOF34VRi/i2PhH0bAh/cVz0CZocyygEkMStufK6ak4OLRMfk99wsF
WSk06DneR0PwbmqGw1NZCK2lIr8D/Ss276MRiOpTUmPg8h92ZA7/nqR//hencxjszB852ZO8LetR
kvOkBdTKq7T/3s9iwspHtpqODq1IYBl0LE6SByfulb96yEfC3FBjgWaqRfPgPulVOvr7UMYBSJi/
LoR4kiPLEig1PagjTx02Z60Baf0YTAhcDUFEQKaLtYou1hoNTF7f+PKtnPQOjxZkQprMKfWZ+Ub6
t/wLhQ9ua+5TOkFHWjsyenl8PrOJ26bcaRHANi5wBmFHNMx1zE9BbI7Th2+wh0R24Vk9aJhMP04J
lgafTAtaYbMbH6efspN3WX3PLK/hspnqBmSnrrUYNbl6TpTTVSqOoWdDs4taE4xRrqSP7viT8esO
nWyV0foYeDBvqr3Ik9i/Mwk/YjMmjC3gx4YfA3qPZRg6soG+Io8IFFQ+6SxM8UNH6HZsG7X7YGNH
WzW5NgslSExFJVF2f3+J+VuQILmEg7TkRmEpR529BcR7Ula44mTAHxNDucN+eFBycPOw9oORVYoK
DKuJUASpnEvCfCV60Ap06qZS1wIKbCIIn6GsvwWQbxGBBcpO7Y/O/p4ysm183269C6GPGALXI1YM
beQd24fH1a5YwU7BS6y37KIQjay2l3M/zi3SfKnJCfsmlJuWx4SIkzbalxSeQy/ukhjRwAus3in/
WjfQu6E2ZFwLGqO+8NZOfRLJ0f1mUoa0SSj6gnRJzz13QNxocTtz3hIXcq4KyaIfuA5oqMnQph5J
/D5P1sep3d4XPCy7Yz69DJyQDRUjCVGCvzgGG67E17DL82T7BOWrjQFEbbab3+5bl68LqoGyy+Z9
OwW2PSW7n3bNjwhUBM6XC1d1TqvY9THmt59pBjhnsjcrkGtPvUr77J508eSv5R05T5RxSZnNnu1w
fXU9H8Ind09EeGRwBM4516+r6lLX+lgjHpjimoG4tJFwHigpCRY9DF4fwogZaImqywo+o0YBtF2p
soKV+pqwpRdvRLogiZ4/fXsLtP3avv5Xn36ordAtvGQ2OZYL1p9ehIKrRbE6ar5ZGjrJ84xiQ/Px
tSzlIdqiv6QxJ3CbJTirXrYNk4VilpM5N0r4+s1jB6s4zi/7GlXARfHrOc34naiGwq2GnfhCfaAq
CaFzwvV79wS1Dw6V7oNgdAQbDGDPZuesUFdRUGG1ph+kdbFLWZUoH5NirmFru65KH1irF3u5BeJK
dl9Jr+IpmKHU58rC16iu+QaFnN9jBoYNxLvWOfDG8jv72kYQg8p1Z4HC+8p78xUfUygYs7mhn3bH
HTVfHB3/tCArmZR/npwhE+kHT6/NOCsxHWnXR4wZdReMPcoSsg92gS7mLD7w3IpQJ/oH7OmnH1Yv
/HVHb12jcKTfEMOISRRbgxqJcDLbQ8GrHAS4KT+C5kq22FBc9SNF7545/O3CteJ2xzvRgruEVn/U
qK9YcBWUMRMCQVfn4I/snjCnfKhR6w/jLomkUexM5z/qytBsm/7PgiwtvFPh7dqy7un7F38Yt+nZ
BJiNnRRS1z0rD2IzV/nJJjFnIQvdsqhdRAz3c1+xdJumsC/WwsnZLaWJVa+pkCQXqjqowA4SDRz5
+Wlx/vTNtktLo7dq/orevqGf9MP02ZqzNdHFZX9eBBxXEsvoU79jqf/m5WMYFs/OU7nj7XFPgVf2
rjZqST+zFJpsQlokXBK7ikDrM45vMRUOd1kmEQC/vn72fHh2vB8MUMtowMXf5XzpRLxoTe3axVTp
RCyFkBByOibp9KJFuseVoiZV5RNntr+padrvUfv7xjV2V3IoXR646zoxJuox5fzFMUaYc5bvQrMJ
yEM02vj1wBqVFSWKsTx5csr65Wd6Q334VTnNJ9l+MtaDFobQFuCxq6nfoOjXSzpVX/+xS7v5xHYf
dRdHk+6Noncx4F0cvWEAUfAHf9etaB15MHw32qsra0uvSBeqMaO2D4NIyxeXYfvZ1cLqLgRSb5v7
uJqJK6tG7BmaFx1OUxfABvz6ehvXfW2BcQhEKs8atUcWqwKqm3LKQ0//oKjVuPo8JPZyBTH9KS66
GCUaf1aZIjgBIbGG+vifNkkz0siS8bQQbx40RsCdRcVCoQKt1mJSU/Y2LU8BTEB3YM3YuFPMrNAY
bVJ9lbdDLfvayIjhowWFmD60Whx7vYZIkSuWg1b6UTYk40UuDuHSR8CBTZPifs4zxd35UBOWI9j8
HG4Inu/hxUqWftxp/DaMwiobCwdaKojZp/bI7+WvATaflWl8fpxLfmU/n4sI1XFQGtC+zjBCYDil
5U+Ucf/Yki5v/EtTThsI8z5TYXCjDxwJJk+ylxrfK5V2mxFBHFsqo1KtZghe6rwyElZR8LOPPrGN
S3sfZ2JzBjN7YHVbMVrERQmvLEHELBkQRC16fsFWKvTp1NIylTD1UiiiLC5aZOITE8agw1g0usp9
UUpDKV+uuKO/haVzr9FZpjB8JUOXW4wAv5XRwEFW1isBx67QNMoosDUfx0WiN0GXq3ebcwuUjEky
ICnKlVBqKrhV4LYh0pplTYnaE2DvJhyCbcN5/3H1AZEoEgHH6y8wVY5xRcBrIyMl2WFMpJ041BPJ
xYEadvjd/1U+oWD/Chbhocgu2iPqemY3GC5Inx5WU1r1cdDyoTWAqHOFqWmlgTnNzg27rRicd48I
adpo59TdenOu2pneVf93TzBoqgqL4t+C0mdxTEWoONC4BI9bUnDCJD3jxHaN1I6eao2oPMAgK5le
xpUX3moKzP5WlWvvv6HZ8ugvcb47PupkA9zaEQkfi0yT2no5QX3XurDbTczKcCsxLNEHiJoUDs9X
sZGCTsB+Y76KY7vUt5oEajyqZ22xgdupqM+HEZIvPmImwKn8jeUhwwf1xChscmG1VNQ/wk3aJoZM
Y9y26Mm3TWu0CBOLJnk89knY9kkQ1sVP1UiNayv9MGw3E0lKWuW8zIobYFkvNfwranmHTLkAG23i
xDN19DFdCycFQ2t0rta4AH7Uc026EmJGgvVX1V3cIRFnkGgWGMASYDs0rLB/U9S5mmSjpNgQ6qOd
/TcQSdzDMiqsYkHKbTyc8uB0myWApDacgSruJ5BuZZa1n+5i/GpiPWjgkWNGxHclM+s9hzgPr+FQ
Q3oipjwl8oINJ7ko53UWmGMqp/Ztp6PZeBNN92/9tPjBxnFhhDEznsCubDngoW0hSIh16q/r8SAL
o0ZeOkAdM+pZuSXqWCPNMTPZeHnHlKNJ1eHS9Z3rRb8qIeJa6bJkwnSyxaoAzIHQFUNUl7DH93Ek
syhi4ZElryLm9oWyh44izrdP1GbAnhQtjvaBX1jGQ5J550OQrfAmZw/z4jA90jpxzndwlxkBkDhf
SLqYELX8836kIHdpRr61c2W4VCBaIgWSL2tSk0sbT6UFg6HJe7mqzP8fLnXeqwFBVrmGr/yAydKF
8dwL8vqvDMBbgzgintIyaTss3SQtdjpkS4RkOKXOEXHyxzwPyvkY/kUaJEz+bk3UBGQtoO8u5AOF
CB4KIuZxmKSM8PHcZP1xK5Mwy2NeF3gRnnBSLK095bwnFZ6xAfg/Jgk/6TMNjV/4b4F660GDSs7v
TbBPOLeln3Cmojxr3M6g5ctQnflD25hrTs7XR8VXdnfXPKPCPmglz48S4XeJtjiqKvyV1EK1bB/r
A3DavM8SfJMiGH8WuCikD95VnPiwQeiDMWry/LZF5IbfUHVmrRRJbvC+pW4+j3roCaY0wgB8lCJG
l9cSt1kDJ6dwWDRsS3zTcKU4ydrhsz/Hu3QixSw886zaJv7+ITQluyOGsJMnkCjFL50LZZCwx/fJ
N9ATovzmBdV8jAe2ZcgI/sGkNCADbN49V8SWkgYORsXahhNfFNK9eu0e2waYqZpxWuFCcvqJqMPQ
hL9XspbX2l8SbgRXKwbtClXOY0eNlmbvIyo6ypuRfosgICp9cwLd2m9d30tIoSXiieJNjH7+8jud
E/KSBMOYuSdHIDLKARsPsixIiXIqpzOG7MDj/DwZuUhv1aB5ndes5ImQ9fpFe10K7O3TdcxxMJHb
PmYERUqogj7l1LDHsDmSXfP8g/v4o99vWRTot4ykLVcU0lLedS5lH5RePydDeYkiWPg7LTSomI+E
nuaPjY98nf8dQSc4qmokha65ZJ5pohlWXvmY5hvwn0mBMHdMzf876rbDgwwXK3rRyWenhWO0b1M4
jKT8p4XchaWBE5MYxccdzFfbIaFMzGztVSuyLKyrQxE+8r8BDQoCNTHhkBvAstWcMT00cnf0PWQf
1o2oFyPkYTbJBFGQYbxzFyh4MXm9ELHsdZR3oS4IyGNqeqIGu232kTbN4UXv7KIwgmpUr45SDgZx
f1YAWDovi+4m/fojLn35rYt9qg0nJ15IK+U6VWU/mKqbo8eNIIqmtJ9e/HWfM3sp1Mgwu2tzYiYm
kmo1NaV0dS+e+fVn1o83jhc1K8kVWAtjRHZKNZ0JYW7IxHnVSjJz4Dnh8GMufJwOD/OiZmAsNjO4
cOdkjH35+1F4eKhBqtMW85WlimHSodmhd+/tSxklWXMHMfxHS0s3g9GYGApBhvuUfFo4LrmMRCJG
9OIAY/au/oMn9CKZp6Ek0D5kuZi0YxRvt6kBonlhwZ1Ve6NwsNb7S3xRVYmMY7sMIkWIpA302TcG
NYsMSvA5XHGw02jiAI168sP4GFK7fMejO1yAZKFGQdA/1Mo63TAHTKwc7obfuISVRSLabeHY1NM9
kg0Eq5KC+d8iQZkoIvdYVWoLHKcB+L8V5FN4v9yrmTqSsPDMwvB6uZuKbYj6wA9nbaJQ/RAKTxDw
jtukEYi8Qmxje+6hsuv8N45ntks0U6oR4pYsaAEVBJi8wZyEimwniaQx4jOh54yGjznYAPHNDDY0
VwkL2FPynz62E7bZDnaTevagwDNPxGnVwT9GMRBSq33N7s6gNzu4I8+wcaXHL5HVOLUXXjMxaZEx
FMYAj3XePXNbsFYHJAxqea8kzuOmiPvaiUVR4exp/YaxOMWObRhj4kf6qP5117sEnRBRvROYEc7u
T2AlpSYg9wr9a6A5lgNT+zSEHtKDaS6AR/rnW9TB8OgHOBmwFdiJgtxUf9D3AUMAztt7K4eRMusE
G5LpB5hl0tjKZIhLgINvBikj0HgCpTZN6YpRvEWXbOTUXj2eLDGT+EQC9WL7e4xgVBFij93wmOv4
U4c9Bjc7+DKLK9Mky7Es/1oywQbFiwrMbyYKdaNVfKbRQgtoF9vAYJq+9lVP5UWaloomHtpPKofQ
bDXf0HM1tnqLOLtkYMZf+9h6qVZHdPIfiFVeL5LRe2cV5QBa1+fpj9UvpPudIhj+91SwBmmSslZ1
PGefihr0t02Y6sCXh0Lf6ltq2wWxUFcyFkj8rYIaoHT8Xi5hMpGMqwUTO5BpcKocxNqGzTFT11kC
ZtO1V+2J7zivy8c1faEuF6ifdSWGkWADukvLNeqR48Y3maFPQGxFkC8hB1UYIrtBwNYRC+xPt38w
zx+MMhMiMZt/wcENQ1vmVIh4m0/24sQsLV7tTpXS8mlhumujDHXlX75wAGgMuX8HrSlvHrFqRXTK
QYUSYFBL+i5NMkvwCIVvebsX+cw9sOFuY1dggy3JzlKHTi5Z24Qvj/X0pJAbaCCsCCY7efmpI9so
26F5B21K4QAdTASYueO7vMDJB7srGS43VJ9dpSZIUMuBl4vcoaeCqlrOGQq3ZmsXYDTU7jmK1KAB
09sWr1T60dfIJIp95Zy6TLcZD1/vmDHY1HElgDyBogvzsot9PhliIA55Jmx6A+1F6LBX2mu9MDNQ
dkBnyYwGF/ksbAHVSK81B4ERK822UDsAfMLMwKRxCaQ2jOaUvkSZywy/pFHSJuTA4t1zuvchhxoj
AzcBtBNjyTSm1JewjbyTvkxWAzGThpyhEbpSuYa4biMAisek4nIOcljU8iBZWGxcLWLOS57bmSbx
G/Vzqkdog1nM2syh4+IaHsACp0l+eKLafH1iZuYHJ6ZfTY4A2pOOzEW8HVz35J2yMXI3K/VyqHXP
VLPkJDbJdOhZkSe+l5IpnQH4FeU8uILEs5fnSeMgT1LfR06oXRG7BilPcOeSC5EOOwxuZ61PITaM
hln+kmuDssO8cVbxugZfG1eFUUDLDpvEMtRyDBlgg7VkWwSNwdppPZA2ue9KW11UWFAmIHRPvayX
fnCBMZUsYY1vh/ax0rtYX9i3sJyuKilwagGTBYLkK6nSaNLPOYe8mfQ40oZIRYUNjcTKfBjNxLSl
38vpo1Jt0QhqMUVCRYiXpcgf3TJ0B3Dkrgc6PWwk+i9ulv/GMQwpkHGfS6/GWY+A1VhRQGVW+4EM
+TMPtop48pnza0fQEVvaCsUYjgVAx+7kuMugaI2ovBdY8UB+e2Rtr//qSpQG3MFBg+mFsaMcBYAl
/TQFtd6lf7YtPLzkwVeoAxHTbuHW8u+kMcSnNS4BloSr64F6kBIHRhowu8iabOhIfj4bmlhUZw3l
MRslkNWsvWxbPtFE3EP6ekRZUjIkuY0rzdmFhXQaptWryjXdacQEORAfed+29A36IjPIc9fA+NYq
kVj/lua6kl6sTEu98cC6lnq4sDDVWADQ08H3sHUB7n2hN6sSxAN7+Ey8lkilngjLpUvaBxy7rZlt
LjGD07d7U5rZbnUj7LvocdBkpepprQ4ljNw8fOfPgIt3ADNv+gDYHNzEsQXmf4yPKuAF2ZcWvYAh
7zMQ+kLxmYg6VblOv+43CBS/zIkpyVUS78VaLfJJRRCUVDBzDIstJoDamlfJXqFxkIB0jrWbQJoa
dTdpmLcPi797RfQOdc7UqbMlFcWiiSUvOUBNR+xxRlL6US/qwWM5YojJdsKcdXk2iI/79Ksl9JM6
G5BK74jYswNj+yeBpom5C1RYzw3PetI4eY6ypAPSF0w8y3hlbZo1tJ7iJmcEfbizAXt/G5Rw/ApN
yvwA/7aLGlc1in4D5fS9A09NgHW0DksiJUFOYPa+PZbHaR7AIxhz4jCpQNgqPCix6ekeg0vhQFRA
GkSp0BCmLePH2PHHNEs/oRvz+gtwFMvJHxXJFBnS38iEGzPk93REhdBToUlFGVK2ujj7vL07MDQl
Qd9fz+4c8E7WKwH5b5eLz2pQkqwnbHQ1bbXjnTD18sVuSa0Gdj19gw1lEG8WMSAEh2ZKwZojvMa/
3RfO06ttn2s4X0/8hmzOnUAOquReDcNkbAGq+7zHVT5nKuicIE0HJzATxNLQCTOFf226y3iN+ff7
Lhd4fwyDBHAvUEamuruYqgStWsg7UjCbUhrSx+xPmR/elXzBqPURo6826P9kvUdLpPInzvTdjnRg
KZUxuEQqrd2Oqv1Ct9u5G+s2fCeASrGqi6ZShKG01SRkklQUBBBtK6St77YHBdQLQeOcQySSNWun
bqiDEVnd/6tKOZ+X+yQgwtjONP4wDKXekqdO/6F6JBaEKyDwdnioSOmABDLMxpmTkltsPF/kHc5K
6utQxxSaCmya4CZEJUy10DZ4BIb5X7TWB2N10c8CyauyGEGiBbvc65+ONl0JnvCRO1gvBSgYKsqS
mIX57uWnt1S5kbc1MnSGBcqjnTZfWaPSk1FUshd9Y2hjkcVk6DBFWC/9MZUKFVKaqAscqIkCF8vQ
WelzApRG8c/bimjwLfxI3DDCT0Kjjp4f0gaPj88hN5vA/Jet+DzZIJ670QGNYpaSMv7j/GTtTL7d
gMr3AycZ1IBK6I+T7G41BpOOVSdOtBrOySZE+HwOVJEksCHzzlDBb9v9TxMQNwKn+AchDbZDgrcs
+ORx+ZZwgBzUJPv0SjKWH3aperlxASC9KvDDOYyCLqvhFMMqN0DHRSJZjZ6Ar+mUc5HVuRlVFs5N
V0blhb95wnVcULyq8fPbXnVy84m1LW5nGXq52+mIcea1ytahcC5yMD01819wxKK7P9H3K64Qu0Un
SF7ky0XRvHUDZc1QRf6gyB4QzALJgJK/gIFOqnTOVFj2+fbQpQV8TPqU9Pss3RMNO+1bu0laK/8a
vMuU2vPybILtyrDFbvh3k8hV6D30mfeFhWlQSDnNszjStRAIbEOMRstpxlJm+ex17MhnMlWHzcFB
Li+qUPEud94QkCbzsptO/1zW+TeYsJi/FmxZ6JJcvMsd9pRKglC+bHomD/a+r3LGy0rx/ZlnG3UI
MjUKpHN5CFVhG5BLgTKRy+yNw5OgBexeLhNawka5RFX3bNZRgeUDhE54/4Xmunt0AbxpX4OG+GRb
/M31l27nI6W9wSmaAKqZjh5Ge2YgyypX7QfbRYdb4TqZ3mdjLFECHDnz3HrVCoNtbLtiqJ3vE95H
CA31JJiRMV2PkzGuJ9Cy5OvokC+D3Rzb3EuUD/hqF91bmHQWqshypYeIYEbeY45UEc6sx7P2PIXt
CNPqho0V2hJHxp3PE6+ywXK03UVeoZj0FpyHjBfpB7Wjuyg5so+JcZmN1U4VmkpCbl1Xv72dYYZl
QLavoalUmGGOual4ZEk3VYHLuYt8Rb2uGOiaxM/Mu1wxKQ93jU9bqz0kqgj2QkjiLiZE90iaGzzb
2S1rxWQUCfK2cl9u3VDuN+BgYyjumIA3nMqUji4eJ1ME8v7sXsf8xGE0L4k0yC65JqeHWwE6dQFf
SWAEtkuNVgrdSu/93pidh99woEhfUIjOCs1OD81EUKohPF41m6OhKuGdOw0t6/TD0oFyRqQS0/j3
Ea4F/kCVXpmHIVgB/puXGgwyCKcxBlGGAn4UIE6inNqBlvQQsYSEGJ4C0T800OGrD85w1kTxG5Rj
lWnAsA/jxtCaD5B4s8cz+6Ni5oqQ5Z9+2OUx6qj7oSP+qJQZSOT72l3I/dxzpxoF/sZEiNCLkZzg
nptU3K4T6JsQJ40jhQRhodhztysgbmq3Bgus1mUvQ4A2YFNo7BloWiQeeJaH9eL9dfdILYxePiT/
6ISzQmKDKHBhtycxBam37DJdXqHHQCerrWEbkhQKawhTB9dOVRgCwY5tsAlnGR4eEdfoqTWixXft
77KLexKAIyqUpvBCAQXcvkquCtYnxb+SjVQeEil1hFDUMsT771ZFmHWEb7yId0FKg962D8VuG5db
uE8jLQdwmZ5T8p4a22k5jPSV86XeglD5tY5616Vpm40rUsHupaom0jaefOHS94gx7ze+QU6mIkg/
sDhQS7+aScpVlzcvRLkspDHWUR4vsTlMNdJ2nH4YQhbFPaNM6cIWM6CvD/MxBOXj6Sopt3sZaPE4
zOR1HLA2PU+h71s7ISoRvS8z8KHzn5mipTk6CHa0ZKLPbfbFtWNV3ya9bOXr+hnEFeqiwhMKQzla
TtP84pIRjNo/E22cCN4wyRIVU4a0ga4E6d+isJXg2Hai/wmlES4lPobQZohR0Mocv1C98fsq0fJi
7UM3ytiv6HgWRHN8m05T5G+gq/1uGJY71uAFD23EWRv0QFlTlZUk+7F1b42ZE9g4y06xFCKa8llS
L83HB6jJujLcAwObcKqq0xavoPNKB7eQgXw4i1Vgg2GrKf9JE0cJ4EMu/WY3RMmc3p137fz6m5Pf
yOlR9CzMA9kvBNrdWQQt7wJK0SSENnTEXkw9t+/V8ueEl3yFBMwwgeEU5KlF2uP4/r6xg+BV54Pj
zAI2uyfPzi8qAqttqtlpUoMWF4fVrsTTlcxh+FuBTMtuOuw3uYe5VjGmkpP73bvNvRPlG/r+nVNa
uaXHoGEB3J7kKYZo7qvavSZuvNQWBWuXjA7U7FYjNIEcmDUId0ZryYlpls74BvyTpSNtArrJR+bM
NtLOcO+09J3OaXS1BCahsGgQV6GQG8NSqmO4nOwVAmP0NRtYjLKyaur+jEuVv17IAAPP4GkBBVzR
3d9dyKhnGoYedr8bf4eyX6emMdCll2KpkG7bioAK588xV2+xiTYlK1xMF4/TCrmCcA4NaxIuuSs+
9JMYR7eJ81o5dUZdAFoICL5ly34sFzsSC9qKDgj9rTh2wNKE+ukbQDTAVYoyB1dRwm27A00dDzI9
WDR7PZn/4Je2cFZdU8c6Y45twpdvKTmUPZ/SC0Y/Hmb0Y486rWiGbOfZuhxKsgpVe/rddkB7vW7D
3FA+qnRhPb34uxP8DhmJe+q5q1sRVSwPSxR5/PLp0ZBJrSkVRtELBL8z6k1Tb46ez3qk7na99zck
CsDL9YbrUUFlo+rjpozM8OnVZa7GmDhV3OSLouxoL0onzyVz3o4iTe7piThBCzkDCf5EpCSLHdnt
3pDN6BSHWxFZ/FJlXG0K3qzY4DcNb5/amXZsuPYCK+acAT66Nk9DiYb0xc1Dnix9ssaKPNRFHzDk
FFsaJ1OzmpXbbPsoLBuq/RfFws60Ufeue74vX59yfRtPSuaCoo8AdgFUn5BLPicr6ReTpGRQoBCV
mGNgt+HVcgWMdqy4FuNrm+6DCRKJXNGMBWRVaqm4tcQ7yQFHtwLtHrYWDsyi0WFK7mhpqQ7OGjXx
+dy6K4Jwm2n5enjAuODY8ePYEd9yAd7boxQXC5sG0fpogUm9gnsEICvTfUeFLBMZuOIm6q78bQfP
UkrTzoKCVtEzWzik1a4J19Lkvu6rRchLk0ZyqqIRlUdGqD2PPBHaNMXmCh36+w/8kYQbLTplHM/L
zSqcnY4FMv2zETy5wAJtzhfHIbfUSp6ZFM1DckTvpSazqyqpGA5hza1vbM0crzVFUk3ZNiwmDT+C
cOzYYGOd/b/ENUS+UoU33EP2bdQ2qA2tcjZ0+gLuSvInhueYG/0TlnzzL+XV0QHLYe8EkxcWmHRH
jqNWIZWJh1LACWose4yn4CH+CMz6Fg270PhiECp5ARs7gJ6+5iN+1SItyiaDTBfYOOteRP5F+Auv
mbUWWYQ4zZpYyQoDeSeHzgESZOPV2t97f8EIaR/jGf9NbawruIsDZVhmoWIbU0BypylVOqwBo2b/
NS9SKzD74KPMAYMnkdrbt5q8D4p0EpZylDVZeQyp4oRwL9rjVwa8ksKUdlLUczyqdhgUvTT1Cpya
qBc8aDSosvYreHWTiNJ9jip/15uwIPYoGorG9LE1iAGNHFkkgKkZvNrfTujjPhwcbA8qaXwMdCAW
09wkLTCCl0ekRiwrfJrezIe9HFPp5kt6KHvaOLova15QiRjGKeSYvSJziAqvgLBN2NE8m5iBU6Gk
dwffuyPVC4L5/yn0AIYj78hS3E2hBm6q2PLef5w0pyE1ppztUtvwIMJHRpa+JVs2ZrT/oZzz+4ln
ZyjGS0pbI+m1CLP1o/MeDxdMShHNIhwG3PoGRvy2DNK8E40mQ8NrUeDi2iCjcJ+hUdCcLRzfp7lZ
SHcS2Shpu0hIQKVYlsDMTan80ms9spzbyKeamxoahJhMXhKN5MgH0AZNNLf4Ph+1pWyVgWbv+Q3Y
ymIVCWEDCUBkoKtKaRl9WRVky12YuMMzmxnbMnn+kq298TUSLPlYbVW07FCdPBwRYd1EKmo/mD8+
07dnWq00+2tXKQhafkIZldXdzDi02UpRLVurGeHc6Jd9au0KV4yII3Hx1T5OJohBanwMIg/rKMgU
HTow9Z1OSIPRjiZu9g5S1aX2sEBMmaVuBlXNk7TfsQlHOY7sTGhU5QSWH4j2KBqnk26VccY9Yr+h
yf9tkCiEsDTdk/SVe1GciH2pbsmWNu2dXKcuC+rHSKXy9jf06QMXIsWdVoqnVv0iMajtcXM3ZWsB
LVCu4//AJWA2f27jK3yXQGjAC8kU91NQqsFAHtB5Rxf3rlGrUI4k4uBFp7zgDavwg0J1LhPAbGCQ
HRSjLmNvm+YX4F//0VngfYLEIYyxQWI0Cf8NumiDz+2HVmpMNzBIXYXec8k8ttTOPRdg5P0QEk2g
f8lTmAhLgbrpO1J/pnOekG0bJ50lxGv3W/gUJhtOb5VGkEPoc9fsce/L0gO08g4UdDZyorL7DeEP
7UhYto1+/rXbiF5OLVN2Wi+2pzci93/+n21qBu40zkUBE8KvnqOKOf4MjZhkGf3UsdwkK2ZUWj12
ijNLShMhYYOzKdYgUrfVmG2N2xrywcGUfO9a9JqXqzMKOYkhTrsVbEgzL+u19Yzf5ngIO4AFwdiq
mFAqLeIHT+pY6Ke/nH9QKTYmylnTFAxsE4AKK9XFK6bV3Bdbq3vJoLq+zrhwhrarE3hVIQOIf2Vp
a1xIZH+aZZ+LTDlJFgVAXdeLKkizuDzBK1loM7XKfvN8j5fXIUBjPL+/G90pMP1lxdTqJ90fEwQU
hpxZbSauJa0W3HN3WhZNw73E3EaP6iURVEhL/Uy2o7jxP2Y7aL9k/TKFYxc2NNJFhFZRIy5IoryH
vuQVxmxyLX7P5zW7h9Sp2+b/T82/WPAowRqWjyt1FNrgFD5U5R31yMLp/RYSBOz1V7q21lvT4YNq
kOyum/K+SRoCXqSwXlIeAZ6AnTbP0q139YlANjBCUznkflDqQoGKu0ITZ0TeD8ByatZiN0Uo1ZUF
2nkGCQKH287EC6w26oM+Nl7Zn6BDJptyoCdH3eDp+SWJQbi2/VWeejsoMJMf4tKBH6toSACJkG5R
2ycVVMh6CzV/ZldTTHlw8s5RahUxDOQ1M9LFRFcau0vwOuZNAe83E2A56sSzIixMQCKwc++HhiDv
Wc6mW/U/ISe2n7kTvxLcWsXnktRnF5fELQs2TV0vFZzW/3bAFpCTlmpbZ8kkVeRUUVmotLMQ1R8f
leyrsw9bCbMh4sua9fvUE60glzhDzab5ub8os6xNx6XQUCv5+par5LAURDzLr2i2H7B1OgIPOEW/
ptEuw6yiFgxHh+wtdzJ0lo241YzgSYCE9cOtc/PYBvsl002Bbjc2msa/2Vh/TkjvyKfO2d/Fsz7f
0+fJxS2AdcMvKhxNSlicsNej/OfTwxFTccRSWM6zDJhg3FgWTLAxJQyxnM1qpKhL+wOfz4BNZIsf
HW7Awim8aWE4t63DOuzvxV7etB79dwTBLXRsVulEL+pKzoife+1t4e9TDX1igADEvsVg7wj3JqF2
1d2rL4Z5El93lwhgISZbr5m7Zplc2FAXa2b2o4x+BWsfcE66ZE5FkBuKTLAcy9orwWjS5ukmijNZ
mDZCG+N8I96bgfb/abxhaTxcsk9RN7caCPI3Mc1J8klVnClYpcEKNEV6qNoYTRZ0xviPRIdvNp+g
2qUQwBozUga31DLyxp73UzCUNXE0GzJxCZG/vbeI5HzE9yjjks8SczRjPOyFX0C3eyQcjyJFPeQS
q9CO26RP/SriXRtG7/Xcr7eBSmOtWTxuk+fJW3RxfBvV1j1hWNbBPm75GEdEn2kwRsFBY6Ftx/wv
iGscjAQ9dVAfMdVIdcvUGpWE/1xK/vldrmI0s7y302r8TN2+S1GgcBbSMnZFo94utwsY5VLG8cvr
sN+v5R4QhGF+oJk82rF5DsKFRokzKRkQ2IHCCJlTp3UX08FKEc8bEAzRgZgi4cbVklyOAYnt+Xz4
t7HmQWoCLyHDzIJKD5kJ82XZEjdWjxTJG8pVFtEaAwSH7WhZSv41gyOmIcTRTO23/1S5hGDEoNiq
ihL8rX4r6aIrXEhGyi3ZY37TzDzaR9jTLkqwoDEZDwPwArVPRGGYfospNDYuSKQcEK6sqXoElh8v
EjOEOZW74S2sXcXrzUWqzeVu85vNoPpDyuo4iuyegE7YLKI2EzC6snIjiSAEINTnkXA1SmSQTigJ
maDfSLpWPFbEUxNjyC7ZBcUDVfOyAKmWZQdPRAhpPX+AOLzUv/WHfOGos/0hP93u3Kh7W5p8GNtp
BxKgCCeyuEw5ap54Xk7g0bWUdjw5+LrpGDy4SL2/wCXNE8vV/vvuapBemb/ASFXF87QhAzwEkQzH
iY4D8ZJaqtJN4KqkgGRiY5/4D18Uk+K/0F3U3LROP7bHo+zqZZ92Vy9e7YYJlDBfBoqdgaG17J00
wmCEjHT7d5wa8kIV791qq809i/CoRzBVbeUUQv0rVY8NYXhIwowLCcy4YLOL72nepKoel2jmS3xk
wkvGQ2LcbdcW9Wmy8PBNreHq4mnDyf6OupUgpy/nEirOTnH2MMT7DpW79sVgX+WusaeTYsIOH/ML
2BZVkBVRZLdcmBfhr/lFbxnZzh+WQuymHEPr1GsnaAMWVPwigu9eQxFc302a8kBLfHKxF6/4X5gG
y+rK4izA5xz9jYzfWcpf6awaGlCjHS5uMooK4x6f4/EwCTUYHQG684wxPvgCVOuk/5MQSec0zJFz
IkoPT6+qgDLMS9QuHdy99V4MmcWklVghDW+h7TP4jeJh4t2Rf9z7yrLrpK/C1M5/DZTeLFBc8gKk
48r9JJRzpvI+hXe/+XJcUkFiwNoMwtw54guK+/eNGGsvzsWXgHmJ5JirpE0ez37DcI7XStNiYywk
dDOMEDL+3IiGNP1LrljrO+LvBbMe375SDER2cyADoH2s3Vr0Fmy9nFmomLDN+9HbNbdfFOveVoB1
0mKF02eobZpGPb8f66h+vdLDa5AIAhowapNaLMNiyQ07b5t9tUN6sACbcKWCeZ+ZX2+tm8e+RNKP
BAzTZ7r8BEw=
`protect end_protected

