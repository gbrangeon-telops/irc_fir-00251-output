

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n6SxQ4cZpYT/ILbURpz0n7m3/CtPg7Srwf+5G6B92ASMc93ahDGfXsRmbxfQ4itjqNp4bImRWGHp
TxDOCQa4ZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T+03ThTlMB5LbidY7dBVWlYp0mNjkvlbypoxh4ls7n36ZTLkklcCR9ZkGKPsYI13rJYYLwxb8HQ9
lAxKeG9QmQNzwwKufgYFwBDRimvj8pMxUUa5UvV+Um8vyzZZSQmIWtsYrZE6EEbBovwAJw8AOtaR
U6gMXGczY3zuLvGCvAw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xyeO5Evu10M+3X2Afou0ntsX5ZB/pwkUmxi6MkSVEZEp/q8vhRIBXtucD3zi9CwKskciGYDIN3V0
Echz03lkOALKA28V6TwxpTDjOCcWnPUs+SbNU9hrNos5LOcUeyT/Umkuwxvon+y1+GmmTNBs/HsN
LDp012R0drMTXSZtr1fQtCR1xHLj1REwEGmrPANPbJm5g9t7g3uQ7e+eNRUcylifmDkL5SHkZMiP
o5a6WQY9gEml+rOEV7XkaZKFEUQnZO3nxTVqbYgCz7Fr3B2jvSfBBfXQPG0AKW9Iz7aUGng8TS33
LFSc4gt02mCKBH1NOkwuxP/U3rpVs0fnK6xENA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UaJ6dwyNV7zPNxnKVFOwTBNM7GBgDixNLEFTEeGL4zxIus/wUjUkJRcBksOgUQrjesNLi9rSamfz
a+6oBrRU3NMz/a6LqvgLX0FtqLiIT69wj/tO+121sBluFxMRAbLYxwtNx0oswICZG6ot3kY7wUo8
MIP1BRyvBE7h7gUe8AY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iLkN9pn78C1qipOzfdJflxHJTY8JBXpf4rPYSCaQgqf5yt0IOulURCvwg0EGtXIXYL5OVuC8GGss
Cxal0AVlk6DQJUg5tnhgoani3XqnRusVYV7ivY3j4fNdUj8iyFUm29wArxnau/1wGXLQIbXlD+l5
Ze35HAoJRWjnvYyl2fMDrjYG0QtBEQHUh7moVIQ+kI8DwofjU8zFsu1KHGJsBje+80Fr1j2xEByY
nscMu+13hzF1cQaS+Ce+aroaWDuHJWx1kJ8/T+29qUQ8IgrJDtRVEWayMxcA9x6qrZ8JHoIeOcCa
xCl16mCCnpbqxuPBt6lvzV/n1cAzp3w9LmCffw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 87504)
`protect data_block
mKJYHd26GQhvizUABDHvIWqqy7dNjApyPJ6F09jDtff0Net5UYidX0QfkLs+OxUv6Q7Qrj4+6tPu
HuXE5mKpptEv9Iw9Pxl69j33V0xSH61nV1NrVXOJmkicWbMqHzJl9zcqouB31eqPwDgkiMeVbeQW
j/qBZn3bjLHNbFrktKxLr26gAYx12OPSVVhjT0jcp9Canp/Vz7HRgkUBFNcIGtrOgQja+1HDMcYV
2W6dh4BWNIiw+x6Hl2CJDCXNhmo8MSeXIoZbOOe2Qo5IYVXiX3x0W3UMLIegQd/JPDvtrZMpG4dP
/tE2EMfhXfHkrPAzK07vlpYIN4WW3chyzod8hI3JczCWNAl3S6a0b5o1djfCgnD7qtbgMnTSae3J
3Iw9v3/seHfq/o/vGpFRr6PrlM4d48np3HBRFq8yYpJ7NKI0E4L55IQhD9eNb6PzFGiZ8FGuwajy
Ts3byOoFdNT1FPHZX/Fv69uJhnDVOu8WmsXhNM1fwsSagntnLW0wctopOXyQI+cjJ76b90qExz8Q
a+ZSzuEo6dl63MLw20eQtV0tGN6plh22eLoY/tG92jUK+xpJv2HI/e7bfgEaWXQIj8GV7KDDy/sH
ns32XF3lvbtzJCWEddEvI+4lpmcv4mUF21T8Wb2oc+in+P9qX9iuNFH8SA98ZYJ6ipITqGMq1qwv
2OjwiLPKcLSfkxwxPZV5Wex/CBjaFyYXfzRzKHDJnrS1XtrmeWE00+l9wHzIZVQbgNMVKBbIYyYk
Q0Qcn7kMGdQWeEM+t2pmIaJVGfxn0gQtwMrNjrfgULMkDvPQfzM2stiio7b4zwcxLliWJoyZbvlX
TU+hDGsl7rRPOigvRlYG5KO+s7QNWcaDYE/1c9F/N7V+UlVc1gaTOr2DJAaBdjJfnY1FkgPieCH1
Rxu9Qfm2IQevmymScvg0781XayW7JFkFTbNZMrwxSRKIwuGtiZoiGlTW4ZSHsOGtYZ+fP29MjO0r
5jukN+61JRwHhF8yb3fKBaoJQbH+siwzd6T9nNIROukm+VRQ47RXXL712RLbMl9WARtm5RONIoGZ
bTA0Ge8dGj0W3EsRZAVPYYxDRZneXKn/iF+1daTvt3VhJTt7RHTOIYVV+arXdMbbJ8lr8oljbYyd
Jn7YmLZabbaemcWdt06pOhvhL9gBXIcK50UUR+CzYEG5O8stPdpM4rnwu+s52FJbSowIjMe68jUS
UT24Rc+VAqu+sKTkkPuCIGU4yc3did3UnM2SqbiMBglubZwB3xeUg+n6yKCZ7Gx7BpkEqhVXDyYp
ju/Lqd3W4Ncw7mgHg1qDwODEhbutWbjje/ik5x2G5HBZeG2p1lmUJutoFQo4tYf4nCFjF6EUC71v
0oqR7zRcraGdXNW4nLHoFJlfvrdB/bEZ5uu2TGGpW+Q09QxPyJk4hVJRXlfs6tHfquruFpKLdJ3m
3MZDqWx5+P0om1EG8/0S+SF/hJzZV1Tnebu52cr/LmZzf/lyeJABUZ6g2wX7REfXQSHnP9WrkiA0
VU8lVozNBkmMG3kmtV56M8JbT7dubyRZlUfC+FRtLHcOBrNWbh2wfCpyCguZeAlv0r58tyla7IG7
Wnxm6cOQrlhgz5B4/KtcNorA4JT9j0/Mi0AMRiy5bdrb28gwmjlfYrfqIRtNKHwYHa9XWhC/+fHA
wkqA2kLsFsDNMCPAUdhRSODl1WR4Iax0pyI5su372KJTkWuXOK4osbK9aN31I4XtcOz/VzHDLjDj
WWPR691mbC0FNpawLegnL7zEgB76sD8xRcSpMzh/HMnIdHt3JfAJuj1lgQ0ilyCnoEzXW4uVzTeq
NlZby7sgOzulYCF5B1MVBhCJnrc11seZTTonX5qQIphNQZtVzj37tAYwNEZ8lMqV1lq9oZ/pUo3q
032C6ofxbzj/5n7Wk9JcsBWQ2/ZXSE9g63RoSnWNm6WCotoB+16H8kuVUsXeymjuC7IIhUJC6+tL
JGg5rBI5yh+1Q9Fo+Opb+7Lrx0x5depRL7KLiCveoNMDLo4pFZ25xHbfLypwTpmDZWjSsWH8RNtj
+ADdmZQdcviOD9zqc04joDBiNsBUFFpQZb83ae8d9+NgfcqPN82pL0ld0/d/Za9I8nyXvG3KKYnl
B2muWUM9Ci0IaurgTcVzF2RBVpT4KfiXzf9NY99MzjUnQHuLjnSnPUaI3U4Lr97xqjqpqqFex/mo
lEKCLjCxMor5ggAAlwUirmPNJUmwKzoMaTY8z3InutOnjwSqmWtfWTIrOpJBHyz0KqlU/hJVRqUb
BzgZsNDkBJIQQKen7YOEJuK2QoDu8ZpD7ftlcIFAAowea4ZWSGoqe26cg7rxOgqKDUY0OaDRvGzi
QfRfd43Fi3NY4FcXGouY1LdiweKr6BdHPQWBcAZB43LOE/E4mrHQB8ijFBy6ILKYJ1dKtufKk2zP
yrnvAvmyjnMkEP7Q+nRrpypYkuUfSdizpH1PmDqEnn3JTXCcMJB+tQxv0HT1H3WPfiHW/0kFyakE
WXXWO5T474yyBZz4us+pUPP7r7I5cqBngsdIMKws/mIPXJpRPEdxscS5qlrC7zteH5uqQDX/1Dvj
+Lq3026nzgwU/KbQ6eRpTTJhPpRH4w3rEMHr8hj52EtlKO2yT2tbQFiopP8w24qn1DunTe6iEebW
OulsqDeEei6L6ONe+yhd3W5XGYhRiQQFfXjgWZTRV173tcbZWsfiWaMkFwElyRa+oOmgEZ0lSO5Y
FmDAy0IiRUgB5Td/m6DZrM5WWUl6eAptn0Hqu0bhaoBgAxmTSZ02L//8xftjLVOBbOKIRYhvN+tj
K3QvCKpP3hmtdj5TNMxDzJiaPOICQyeD3vOYtp+jkj/STM1q/pOcORYLl4IcZ5Lym9RvrfD553UE
Z7HugbUPorlkNpVAWBMPlJiw6ec/amIG68YDhFKjGIpBCY+w0MBK8wp+ByL6mncjWRixtlIdv1sf
oJNrxk5Q8MoZCo3cnHU3a8KsBUqtFdLBmpl+4KFJr9U01VRLRmGa1Q5YzZnDPMF5/Tk6EW5xb5Zb
OA7crFT91bdKh72KjX6Y7ifQoiP6zRvd9Bwko3ryVYfq+6bNobNdzknJJ+YSutPERj5gcTbop/dM
YE8ImXJcfLHnDeQhm/tKiIX0UUOcHbnBGXoFnhK3phscyZhqUoHcCZyFZbv8Xc7RLHQGISBJzg1t
63qiaUSttY+vecIsNvSDcup77Gxzd53L373HA2gr5p7p+DYdYUvr1ZSeH9eZUNLtn8rEfw3sbr+X
Y/S07zwEbaqj3D0m+JiRir0iYaEXPywhwokNIouoMgP2ACwiaHC4bAoyWMBonh5aWsyVBFik89hw
3k6kxw0kUy8sOZc/pKotg+gTl/2rVznpdEPI/sx63xYshe7/V+vtS9kevNKWaedjPEbIkmiRoQoW
yZnymhY+28IqBYygqqtUeAEuto4rfVHSu17GeMpHmIlTpUrvKaLuyLh138KLi8GHSG0BUMHxgzrZ
dSRzM2za+WpJbrO1u+GiE800iVIPQaCUxTGM7isFLiwyelIKnD3pioqalINAF8QbNOenTJeaR2Bc
4ibFZcMmcP82O8K2lRDwTCOmMUpT76vDR+8gfAYz01xR4OXU8P3zmq3CgJnxWHKYw5bAyCIZgU0f
ex5r7x3XVSyF+23t2lrwc5TbNYoZQAOSyDvyBh70ShrdJjPBnasva6hWQBqYHaOqiT9EmEqDVxjc
Pc8DCOAgjc/BuFlbYtEf38u5DlM4wfYdClZFwwA44IGhx7yYm8tTs8SBzA+k/GNcmoQ2YiBcIA9/
blT96wW3UrWGZ0W1U+38Zkk8vW75GV02Mm6nzSSEAQX4Onm2sOWUwdPetxHx2Cd1acKIgWaX5+LC
/SzWF8nVN+pP15Y7iMhwb0ek30/afW4EDEcuLvXuwtvhOTjtCvaVAautlB72nKrXrn3aJdZY4YJQ
dL3OS/gJFxbO47mT+qTB8povVJ2P1+q78lmr/Zjgxq6DoCowkeSGAReeIA4asq+DbkXzgSdYrPPC
Kht3z+z50naLNx4p9K+xpwE4eqZyPHqoA3an0UZY2phWnJZS8eDR/AWNQsVoG8hJLHm7rqFwihBa
tSWoaDgYi69+sLQePk7LIAlIlY16dU9jCxhACxbX2L3geVXXbkPboOFAGFDpGzFj+TIiT5BsvUBi
lvl5jPW84jYDkqH6k6zQZxsmA5YHl6SXUKB0PawDR5zFdCpuIaEMgnsrSR+xo6LnDkwCrCb3qgCU
5DLUk9BS3U+z9JG83U6v3Qph/nZUaSG32DrFrVliaguaBBxDYURTsd906fNBVNGBAcsaN2wjSjri
Lm8KyQPWbe3RUh418GtvxiQofeKYoeQmKM6F7bX5Objle4X/zBPDiWbsysPgT1IRZ41PNN0cYyYA
b5poCBaJr4rc2BT0/Jc19KP+9KSmFt1eHoIVUEC5uIBkHm/TVr1NO/P7YYn48Syl6l6HZAhT3tH2
1mr4xVknoywyWF3Wdfusat97ZGgh+1vsQnc42TiX6qBCzLYr4sLfLDYMWN5x/FHQZLE8l1Pwz9Fk
o7Tk6/4v+8KAj5vM5xWg7P6k7mkBXLF78jY7rmKW0rAWlQOIlqZx+Ii4vb6x4DRdzsHsblrK5u2k
5nr34eDNCoc33ihlS5dUPFzSQg/XpTajoD/XBpYk08af0M1e1mcdbjQ0EpeLKsyD3xBYywSZWQa2
i2e+EaSs+poAskgG2rOxhpL5qEdyNNeLo5ePlYCt4KYwqYjyVLCY5chvyZ/VIborE/2wcMldKxnH
I6MxDDSA7iR7ElRvrxjQnCQBmROAofT9r/8o7U0xUek1tn/ku3QdPvhuci0i+hyAZKZRBkjZXxwn
Tm22TBkMoO4rtjWxVfAPTjXVSeWaPs1/UTEUWSTzzFwXvkpvlMircwfGw8vMM6zFlO4VUZuFL+o+
aEkI1iXZurtOXwg9509Yv8tT1NYxG2b6QEagCMsYmTcOYBcXmBkrhvVzwo8Fs5GnrV6GcAvkwWRJ
b/iZ5thPbTKWwRWXMBuVikMBr5s+WxtvRgkO1ElfZLkj7WvCT5XBwwx5LYtcoN54/opHJ2WtvZgV
GI1NIdJ0De/xDgP/38t0IKl6vCxScU4+iCkXvWeh/DdjZNJ7bVTBUtFBljn8pT0K4brSRCcTlx6l
M0/PUXOZpZc3UdvzjW/ZmpOp5Zg59V8srXAKDt6Zc/eWEx2sV+JzmoMMaza9RQ+tizLdOJKbhxoK
cKOBSG1bj0pkmLW1yLNTOb6W5x0ZjlRJIBwYL8TR3UFU9VX7DjGExA2MXkc8NLtTQ2DnUF5+08xb
Zi+j7NYEyEAZdfp8qUOyzZ+SW5H8TZIOjeOp8LRw8XCT0X0OFi0k1Bad5pP76KatS2sAdDMG4Geg
oMpOK+hg8PEPqtLp25DkxgtbuO+gAfeey9cEjgOZBcaJPhcF62xdaVzyV4GeW+kjP7mspmM+pFaU
i7p9NwTQdv/zZ9VZwTMtiv87t75VfLoICPHnnoW0Zw4iHtMGUB3dWb9FpOFMVMRkLD3QMXWlXxtn
a2xC+x8M81aTjf9+WFWAZDBpZoAJr+Km+ywUREQuQURPh95xjxSexUX13BB19ZP2pfR6jPRbBw8K
oT1tHRn9ZjNNrkfVwwA5H6mY2DePIiKT2jduTMqaLAX4n6Mz4baD909Nmn9PHgOi34puojREwSA2
EUbSAaNaPJBHz6EFwmUis0Mtljtt0piEZEDr064JYFpAfTzg66YhjEtnQI8b2dmNhP5ZQ+Fe8p1C
6Y32kQwAqq2WpqOjhOVw/j8SxUDSyoneVkJZ+pXNUZrlvd5gkdTDXUFuvZqrEeatAYTDqz2mY0JV
U93VdUVeWQ1vyjs9aw93r33ZpU8Q6uODYcPK6aYbXofzfWpmC48a4UU+m0b5t3YiuAr7qx6vBRSM
Z9DAds58LGKSvCA/B/pPPmUAb+YjBr7E+oyRhHDhXHrwObVRibyAd8olUnYzc/YDQgTPtkf0BH+6
3uweBiv/balJsa5s9bxK3KqOXkg6lS0mNj2UJZ/sdxRheg/MsfD1IaRFFj5EOzqbx66ebLjlsCF/
JTRteeunA9aaW6E7zbvM4Z0tGXwWHvCMghSFGjT1q8lEu9b5ekZLK3xSmnhxzO2his4hpBLVuXgv
d/s2GoRgsKkBatH1kl2Gf6nEpU4snK+7wOhFKQOyR6sFx2lvX2faReppdoTFVFWFhIW0NUUshjzM
LlO7O5/aAzhzCVaN+YF/5rOy3b9/YZsrwTfcCld1cOH3hiOw0P3i3tvWCIiYHtU5mpj0/QDMZFFg
vFAgrQsKe/cH4bLkAqSSC/lV67fzqk87AWtx/qLkrrUESjNm1kN4RBjShxfrb6SHqyVBTXIvTWMw
SbJDWoLiCCHTyw6mYCKHg2NqpF3nmQSrP2yy3qPHbgBdXR0ppSdGI4w2Zx+x3SMnY3nrX6d+Q0uW
yIOu190fQdVC//glXayIJKXmy1wC0mCeP26r+lq469wQGLaMp/SgP7TwnHLYElZ2Rna2R8E/vZ0S
59eB5HxB5f7jYrEbmGGXFwioBf3a9aQb9F6VKiCAfCLLgGEivmRDOUvFEyEE0AJjZm70oRPGIX3n
wwhSwHiDCunlisqaMlgtXztzys+ObqUuNkU3LSu1XGMQNDmqpQvzWlqP2tPWOUlTve9KJGJXFi96
lC2bKKeEdVp46hH5eb85wpI1tKpXcZlu2WF8bnWNKU5lvTbO4J4LwMrVK4Vh9He4EBUDI7epkbs6
fRSi0BErfSnsZpwRVTOZRkALJgAgOfpM+3ZtednQb6AS6LHm6h/xRgXy/8iVS67NxLaL+pjGiCHH
VZX2sZHCgKjwg5i7JNnIcpSwZPaxYFegcObNtdI5ZebukDX/JEeRcpSNz0JFY0Odep0Y5iRHtWS/
X9JnzcWWzAw1oI0lZ26GcuqzTB02wytOBJxSG1s3CGAcQOvbbnd6GAd93Lpx1gKF+60SXLFISNYc
VYk4TCnbvGqy7ueuDfT9QWynj7wJviCjgHkBFj1VGO2cCcynz2amx1adGzlEhBYMGePKUnI6zOze
H/30UVWEvWZ4/b8GAgPHOdCgilfzd/BAPBjP254XxIgNaVFxThKp+ptmQqUQ1g6bK/o9ltJDe2Kl
GORD+yb24yYbzh4BHr8SNKJcMronKDNVcnpCoJ6bnEJBfevUa1LxI+pKMKcqb0QyE05CbunvYkjU
Ii//Q0KmPey3ltE5GZwc8Qg7rSrE5Cjk7r8XcYGnuKpXohzeDpsIAm6r/2OtL/hbjKGpj1KFKEiH
oD3/I5itLGMP+cvVUzgsiPNuNT7QOf+rJaK4s2qWu9wG1ArDn8AN0WQ5Ir+3zvpKke5mGqBn5b7D
1NMG44PSxHitp1WJXRGZMJeQTaOLUBmwcWxsdct2nUE40JhGqRAvPCb45QiZ43+DT/9HueMHf5R6
4TXjoZy7IjLa6z6CIK4g3+9XudPa0faVggCdWod1dIZhAdzEPgLyddSOc+Yl/AWaKyBp90QnXaY2
a+5FtyvENnZSK5ljb7bIg+P5mL8wsDJ9g3cZX1tetAjmhDFfpZCpsAzvRuLPah5AM476QmEvLS43
XuUApgP55iUxtBcETISydZ3D+eLoXzt8Z4SDAwPg4MWb0lXyFnr2ElKTk/Ns/aUpgSyBW9OKnRmM
FQV1/u/Ac2Gu469LSejl7ato1fNCMXAiSU9JsKmWhKsfoahuA74xsTcynkVxWmTCtWaS4D6cn24K
LC9CJJmT236WqQLFRROsJ0iS5sL2lep+u06dYegr7oHCODT2UlRJ7WkiaTZjaRD2yqFX0mcIUBYP
+O/EespPIJhyNfWg+eLXCewENa+ZkUwNAQ0L8zrieGvB6lPX8Wfaq8NoA/ag8rDOU5efy2MUTEyM
d84Q+mr1YENNP58KQ7qQv1rn1oNnym0RjBLkfMU0nf7q6acU87KdviWYyqOk71MPSLdQpeRN3HgY
S4rjfUfFdSx0bjEhWJT3fZufDJSY9FkYtkPTWKqzRk0Vtj9vWJmVnXyMUlI5bmF7WpOYRGjtO1n9
z+hLCO6Emb34FEAO73wXvHweiF8v2gXhVUjjIgSBUCuUhr3dhSAlVL0unWP8LaT3tNZxZkLu6oRe
KhcH2rezWHwLHQHDJUPLvxjtpQu964Ulyudx3xY8G5IhiqIzjK/1Gsa+6LPE7wbfkG0TvjgovWhw
vpBmIIvrYMndAIOFEPPjt6tcsLIFg82AOXWq14Eg2xxZprJfk/Emkd5sN5ejIaJmPn3WK6gZlhnq
ri0/G6TBFUSAMLt8mkOc2Osq1iDKOF73iiQfxEhvoG0QUaqHGE2RMbh7L+y8FM2tYnxHEG/HGVK/
XhbMEjs0w9y5B/udgSo+IyXiBmeP5fZfpMXXA0THViWMbKcnpZCdncGP7Y20fx8WTh5wvHM0dsaV
B0UnA3YdskJdKQkmx3TkOFVNJetGfT/1rhTF68TfOY0l7aei2hRO9ev60fsMw6NICkBAaHsEMWRb
c51MN+zxwhk5gkEf/5ntP7icQcLKeOwkdojaOKlx1YoPYsOc2GHuZPbNbjsr7VdueKi27aXWagGx
MAEVwKQ7YknCnk1B1ynUiU84Gk37Ty/1JqN8GLSCAz0Bo22wtYL2BaZ2vUd2IEACFldBJCgPl+53
HlmtBNsRppa9S1+QAlhcm5ZAbWZdWyQbdruAqXiG1nqcSEyJpQ6PJ/EaFy/slsbrDg2EYTkrn8Cr
mqKEJWEAvVc2yE1BK+EP9lBScLf4lZTbV06+vZoCt/jJ+07I/qL+C/jNNZl4xgQ3XvFT2VPjpa/R
8RNzc2ims+CoavEqJhbh/kU1X6kYK9nEiUZ0ELKZosAZashYhfO97suvrElZyihi36QhWQ1k8JUF
tOZAVxnyt8onnFNNKwvK9brx1JQSR5B0q8WgcDz58xfWsK/65PdI5kdJV5bAOstPKdYvjOsd/a37
YLxSMMyOximSDQEVVV4x1rD3smJVrvbYbpFIqymJ8nXS/xcZdVUOg6w9wRC1h+wsOKf1qLGcLsUG
xS0i3CwdjGbop8d/6THJT54MGNI7n1izDpFkYAAGZTeOTCvQTUKFFqfpO5z4qV1anIdCSnx7H3JL
4MXFl0TPfjbOzat+f+8V6ao3EQy+KTNAmDwOin36pb4I8cYTZtEmgQWICPk5kSk5+eQ2Lq9LCk13
k4MYPJOUp+a0rJMPNqgQ/JeXtoJECmDiFrqcQrO+XzMO8fs/LUbG+UFKy2SiauVFnVZfyZ9Xd53/
/bDgOhzeHDr3dHHci/20FJ9LM+4l/Htdj5uABZ+GFX6GiP8B9b4/wnHPCrrpcZnDjgb/2TcSPpx/
rtnzByDMcIlEEH3qtxXglffVpksQP1Vh6BPxrseFtwrF0zHDTtOIe1PS7kVnS4vPCsZNn6m6/Soh
+hL2Px6wig+r9wdzCT0zP7XNDYLPSqkxlhJ1+CB4yCH841xWe3FRnEv2lwQUv40RHhP/DwgQD38u
3/Kjs5PGrxZ7tdmbT0gYrVXMc5WsIscxs5q6ljF7McwKXGm2kmh4zytlvSo1QZX3hWRon7iRIC7D
ub0wwnnjnGTSIWJKLtpElOTcJQ0TSc2ilVcAbPGZBqJAiRHgPtrH3xbRBlzJ/qZ9RzxaA2X1FJLw
jj5wudbhZcJJuFqghMlmpWe/M0WZnrNNamnicUpm5pkiD0rV3Tuka/haqRLOgMojbeQ01Fqz54Il
cMHz4abOVjzqlioIkF98q8wP+Q5bZJ++8FxCAx+7zr/Wc6BpMmQ9UDpIal9LjBYsNojMQ8Sgbint
f7zQsNFauU+mW0srRLvjXzCKHQZYIv3GfePF8BnPNg3m8gdHlgSiy4a3uuG8ASNh3RIO/ttnJt8l
udySfhlcvIwxePymm7BYMH+QX9p/1dB9ov6mRL8MPNIHyXNx9BMQabyqLSTXbQOlZeNyDmElH9xH
ya9BMcazG4x5P4VIPkmKHW580/hHrCMT2mDU8Kv+D6iF/qrATWPTUCYaObjSLFkK21n9+rl8cCSS
uCd29udeGU097jYIhPx2pDdl8id9HYcjDG/moNyDTTf66bIafGq47c31RFvS2B7+eC49fts4BQUQ
98y8jDTGB1XRq9UfJDZ1CUCoMqfe765X+Gw9xgKkvy6kp1yx7vr0PJSm59gpYHUjNjPLUdMzX+C2
NAULPHKE2kktcdnncf1R5oE5ffa05gtkYjHX5KxXXbOHtG/9qbz4mjF9KhsXHuRHorB/YTEnxfqm
LRKYrDx24JghObszoryrYqs67g2CdSnEUAQ3dODHWRPp8B5QzeuV6EYDvchQddRpC6vlBTTyEV3w
bLn+bZgwQMjO8wjxhIsMcMZND76QwR+h7ygcXkEn33W1acNNF1m/umTT4HuGUOYZOBF55SCE9l4B
kZdw7h3ezOA2/2x7UHAc7kKssCbSUQyfLsGBeme5JJaUZZnPbB/E6FmxmJFkx+IRmcMAf6jrXhzs
DYyG9VlHdroOk3jt9+gtEgyPG9jjaImAxIukF1mzwqUP6KYmjzE7zn/3jp454MpmqCGG6S0T25sU
ezLSg1l4emfbIZMYufBi8TKT7sonXyQVlRv728PVB5jHmf/W9/E0LQHjuaLcsdhGVHsXlNzj3zFH
CoUuPxmbEc7ZYSA/HRqIPPLRe9R8aP14HClMtBH4Se06duVH9mJSk9ztOoQOBgOrI1RX4pZxnnFj
85IHILs1tiKCY99wDaPQfKAUFvpCkpTOC3Dnsvw+6bstmfzUuI+equsk78jfLMl7Gcqsq89Go96C
iLUOaN3puRdrQR5KL9LV6Wz79wrkbevywc9tD6SUaT9IxEEtP0kb/S4XD4WFFQpCraqen6fl5Wkw
efBLr8XKt9STm04B2CSvtF5yec3UgEr3h6CZzo30fPLvZf6lhvk0kRZSfjlsWtfyvAqV+NRlqqAH
MJTVg0QFsnurKexiW9QuI+N+KTf2HfDNUv6I4rYpOAOK8NDNwqkIdXEd9jDgkxNoIv/QMtZ0zahD
oLfIN/8Co9sEYTxB7rgvhLrSxrwFX52x21fsgluMfaM8WGU1mQVYI8584qNfEhCmKaQ11R/ujVPv
y/QS9AeH43vDsx+8PV8dRS+9VykL4EhXvV4EV9/47P0YOhXU+x0xkJCNZFK1XoH/Xh2wVFajqYOw
vR/BDVdKKu54rFO9roNzUr2vE8O0XFXA3kyrkf8AiKUjuQGHnTrYpqzb4OMF7G5hNARFw/k8MAyp
TcR7jXD/EM97gcalp3Ofhhh9yaHoMKGBVTP2VNtdyssxZWtCorg3nvhNksPRVRAUDnHMzNUmfYzE
KXRsdS6Jb025JskLodoTWCeeg42WWoMDztMtAWVBNBmGXcZniW0so5vBjuDq+cwtuF73Qs3VsKRa
krbIKDwdn6USFOA0fWxFbGoa8ugsnQm02ravi4k/oLhbbrnSz51L2f41SKKBUNV+gwwb3jxFfnpu
rhBK68Gje5HpJKCQotSUKr/4RuMQfKTqGTFFsrogHpKS0oqc4iX+w+2BX0S+W+8Ksui4JLdc5cR3
71XerPt9F6y+1vvTj6nxIHbO+Etlwqf4GD4fjkeawN62mKhrb7XlMOefLUdYujswH3DRgEq+vByX
Ei1QW8KPM6n1q1NvOFAzphtmcLmYH5o2a5iIdtqSHImgeDtmpa9GLCItkHixFuhj8ORwGnR/fnOU
D+B+J74ZRy3roWez82rzHOh2nEczGKgdzOzYaqdCzkYdQkCv4dRTTOzYux3i7L0CJt1Cmb1fhRbD
5H8UzOAkWM88OD7oRnwA66ov113DekyTsDblNs5cv93X4AQ42e3H3692GwbqVKfRzl25D9qY3DEX
MM7hmYXvg7JQDaAldB6+LSw7aXiSo2BzFH9NWRnZMrTEkdWEB8BmV062jtWBhLnNcvYhG4TW+wW5
lgE/S8VXaVJaakF2DpGbr2QwYcakO2jwX9P5eQr/NyUPO7cco8LFPylmV2w3XnV2FHDQU0RO/62Z
eGjJeTVpPPpOi0kyN0RPwJC6cG5ykD1TBiPOyuJhyUY2WqcxZ8IXfit21BUXEGjsCyM4Ds3FviZ/
2cSXe4ubrwswf8MEiZ53CVmpoWmHsktZ8tcC3E41r0xNUyZ3P49Uv3wWzI1+OU8ErDLUOzSZC5jU
qTqRm5u4F8xLoyov2GnVloMHHOplEHWXIk8xXl8pwfydnhAMwhuzrCJA7Or8LZpHy926C+TZuZYg
8G+hyfLBALWaB3Bj7EYBKjJJcqiGv+0sFJWrOBPdj+l+hJs8HypTI946P74+9hVw/s0wn/LARAI2
kSaIho2Tulpif/cJ1epxK5+cwEzMu0pFIULrPGv7yuKvn8LbQ88MA9rFbyAVSNsAhtt1c71he5A4
GYHlK2dRSoBfemncTV63GzlrUPuhtlb7dsvwSxpu5dl2wNloOrngIMuuLvj+CqPyjSyWVBQAovOP
Qisgn0B6Wkm6jAigIP22bfT4CaNGkGoTfRHMCHxHOrEp0CAV5rGcioKKcZ31a/povHixdY2yqQfm
IaD2ZZXFXgSnSfrEkPJV8HbQZqS2Nguw3Y2Ba1WZLI5YgG/g5xBn9bcFArl3W5YgDTWxj20Y5Wnh
lHvHUp9M6psREPAJRmI0yTHLsWgsRK3/ooUqdVjBNJYaZTL77nF9qFX52dOnFqHw2wVMag9d4Qa6
/GbfI5MZN9N0yYCyB5QeAFVd3IE7BQmLNOblkD8CFJ4tSomKZbZss35CWwlngVHTSoa3T6zQBenX
dC+Pf2zpbbnFWqdaqvAwVrpFnv+xulrdDP9UWZczgx1B8dF3yPRJFp14alqjui9npLxwB3KTBpaa
CevslVK+4Vm/c0Cv8Ip59pRXBzlh64oLeSpaPrZpxKP0RTgQO6PVeEXs6bBCKKE1Jo8DW3Vo9RQg
tb2wo2Rn3tLZgmhNSV2wR/+1MwQLtbzAaY2wTUsw2NiSaE6FzOUW4P0kbghgh80AFIb7CDma0054
1g8JNjLYhCN2h5BMHMzJO/eHb1DL3WxY4mvN/9N1WmiF90wPgFoquOx2NHNsRMoLxicZ8bwHlcFn
g2MY+dZVjqXqCoy9NfVqJHDQuf4//FsmPOrxuZnijPB8M/DKXuekGVu6uaTb2iGoYJ2Gj8bWVF4B
6Vah+Q++zPG3P1pKMhY5niqQ3QZmdEpxcwVPMGSJpl6bg01xR3gzqxXE5QTPYfMZDv2XadGo6btd
iAnpxZjHJz1IdfDwzYNkHLOfPRvFkiHsi3/r6rtgEOWwmqUx9NYCqQ/laLagO6Yc45UK0tiHrSed
G83MHHBzserNqyeU9OMnrvTSkTTobBJnFFKWuwlWSNzHWMcDyorUkZOy0yjw4HkDAkNLwPQxoIqj
YkTb9/8RlLR0hfhCQMpyVw5qICPG254NKX23z+Unyfph9jUfnOIBBu3n48QCrTqXomkXk2+iqdph
fSKhA/qOA+ytzS/rVCsqhL3v7nHUnTyP9ma5WS1u45dziYQcdFeEHpOpXxmur93jAIYIPiOY1GhC
bAILIy6WFnNsWxXYa3II33R5FIXsXohOfw2DoPvtLgQIB40f9S/97lTRmrvRJHdJmo948vp+uobk
n0SXaGH26P2TTQiaM5sqfNpRPiiE+aTDTMt514T8cNnyPh/YWk7jIMY/oy75Lf7mjzVo15yuCyII
VZ8pu87SZsPcHt0BoSIiM3o6heayE3rfaITJlkbJHlK1tHCMnXQGT/chzOvMhoEEw5A39+w0kSWS
8AbjEmMoxekOwN05k4WrZAFY8pme9QLgpc1NeBXtSOdWPi2G0J2RUdGMLBEMsf+Bc1iBLVv7eCBC
2wQaf1tWQs0endhX7EO9cMM+a2ryhSO11i9zOhX9nK//RX9H4tVK5g2yQPoxgacOhGmUI1dn+s/O
6Gdul6A16bHeaBQ0JtcnEtuFgf2Cfl65cKTXcxP9XHNEKkRYwFYAHYnHrPNnzBkStWvfY6lzL7c5
3YMHXBmtcLONpawOrYKeIwOYUShKLOKGcZQ4m2v+CtJzqi1ZJ2Xnpvm9aHPcFc3mlNYG1R47O514
ORUmhZ3GR9ElfpG2EnJMCxdv8xVzTDNSCa4yk2XxyhGWFotP49D6/ilr5ry7DILhlPht57N18+TD
tijmdKn6o7otDijnKzuzCJnSGgCpEyMIem3xXfflVJZCIl8aD1JjaAJBrkZVATM80gWx78xOxo+K
jdIVuNCUtrps/TDtrFS57tdz6VWr6rpZ+4BLyr/5eJ80eysNURJTyR++Hhigikk+2Bydg+xguBc+
4/cqturUY+S7hOmx3h5IG7MbccnxPGKjhl/mpuZysMat7ggL3SYGbyFvRxGs1w9UVZWw191JaQlT
+ieKLRyqMNL4S/I82fGe0pYwcqXkZfeoDH3Gfg2tvKVgEIAxtXYvWsvLq6W4qIn4Yry9mjDEq6sm
hyfpUb8/YI54GGpOSEbVnq+yDPIbVP7g7yXx5Do0UgyuBas2B/YOe4Kf87RLPObJJCYJlCgihoHN
bNX3XmcuRcCdBkyXzvicIOP6chNkhcvCIR4x6Ygn8yzF//fR5oMf2Oh2EErNplqLbG3tDDNWb8y+
jkE3oprBLtlEczRgingBelnE+T5PYrtpLnMK6KRzdntnRQhW/ndKx522sj/BmgewRydzbM12drG6
kLC/PG8CgJiPNwHqXqHSm56p7yvb12u5/hsePhM59zR7jyu+dVgl0rNIMh1zi0oKMv8AAGugCB2s
hYSILHkjCDKLxY3wkJEDx4hF6lcNdsCtdZqxDfWCZfRkXkeT//uyiRO2wTSmBf/QUudJHy2Ys10A
RVSGNbza0/xDo8iVilylrpKKo7lJvz91iuuBdtXYURcpwOddzBNkNpWw+u0+orZaEHKacboKd/gj
mALVR8vtXo+PnbPffYhnL60tPn8EFAWH/QZKc5juaEOgU6smAA7yfwe+Fg4ErhpYFbX67pbVdoJW
pPY+w5D6rU/d1ykcJdZw3OYkNFFz+aenZHED5+4pagTjqwn4YuLLUq8cfx6P8909zbzMaXAtWmWi
RRvdIqBCj66luBr6fRkH+ApwFq/hjC8Zv/AAUvyuEnc59wHiWnCjxMbEIeZRfB7oRtQyls9WiXb/
OwUDqf4helIcvA7gaMEP2FnWhhRIzL8I7NM1lPb993jYFTCCAg24DsqCOygFd0w7qaPyq76+c3zu
tKxYpmEa4VSkvt+bIyrwKamjfL9iupTwh1DGY4j18ZXhrioovlhvpbXo+PskzXbq7Pj42fzgEure
/RqySxFvw1155CzokmZoVQgtbXxnLjlO3mSQwt9qeFnn+ogDxrIWrdLC1vm8xabzOFthmmyLI5z4
ojXBS77IajlnjgoY5u4kH7EeMd3G94TqS+DlkNqXSQioRvVgNMqc22vS+T9ijhOE6nvJub0x6sr5
t3lSgB5oroMJARP4I5QRvOoBtImlzreQpILdPmRQEWzWsSlOML2YqmItJ5AkyIyYX3o1PMTxR96c
TyV3KNnuEV2ATG4GTRUVKlisXdJ+lamHLmFUoy5qHCbC/ALHTxMqx7mNHcnBlFXlKji2ylNPaUx2
d7DYzoZe46gPMZAgzzh4guIQn9DALYRKIKO38v+vOl9IsW8Bc5HQ3gI7HeiPoafZmvkKz64t7Ise
ktTUdhyXOaoEJnV7YpQ/bE6AegpZG8BUTW7Dcdehl2FtmaOcMlsv4t9i7sxNvudIGD47+A3+pkcx
mEil4ECskF4fWaWqbFqdjYdFiuxv/xezryA7a38b4UYm4LBSpPoO0uMOCf6ojM4IlzneG7g7VbXd
/4F2fGT3JmzNtjQLFIHySOW/VmF5aTL8BciwCC77/gMpTanCgWuP+d++KGbVf+NVglt+kwRBBS+d
GzojRrFJUm0Ch8985GyhUPcorM1uJY3ziFJfprtg/IBwJawXA1y6jH4jWUU3aGpMsgRDKHa/4liW
uEKQsniEnCgSleAalOUcuUbrZQGEMQGj6ncPjVl3ViA2czNb5Ii+xKFK3Z8JAWCAvay3DQv9GvV4
zj0nd921vi7FOORuOmwV5T56qS/tvHtA4FJDW1UfzvR15mjn1Ydo6L+xv58EHYu2Jxwjw5uluvxQ
+DPYY6SXSFhUO5ZlrbAgx2+su2saAV1BSvtmtXBLlf1aeYoekGa4xfczEgEfHz2aE0mdBzrosm6X
A9gfKWK14yN28LRel9r6Eh1A97NNcmqCJUoKKp/Ywiz/Eif4ImkfLSHuJF0pg56Sgh2l+ZLBK7j6
7KU/WV9W865z3H26agN4doroLVxIdvaCFyyWWxhdd0pJ6ZHqTMRkYGie1TrVcJhdeRNswVLSunOc
3JalW/pdoN+P7SZGJGsLPpmVU1Ngho6clXP6vcBdJh3eGzWEhc34+Z7MPoK+B0e0Mt3HYGSfk2BJ
mSia+rN7aYDoxq6Kij+O5cyoMTd7/3z56y5jn6iyunAQ7/MkGLKEWjyneEPJX3hN64l0PnYqezCr
tZ9qeKkQBJEh8EwXQb1utw67GLgygMYHjyBFj9oJVVhLckC5xhDflsU8ZwvEmf+17BIHzOw3ul9P
fAyGeDTIE2pW7+0Pvq3CH8qZHo2Sd2L0NC2NkWf+6j1ZQhkbUpUck8mqbQILT26zaXy9mo3I1+OM
a6c7m9qJwwypb417iYhlsas3Tiw/9kQLyTiNftp3YhhcQWQ86b52k5LwnB1L6k8UtPDn4KX31R44
PMi3alfI1RHkt1EtHm8S9aJGpyvHpk05K+/4RRcHv95VkGFsnhktOCEu8RVmTBJKXaFkEWgO5MqE
0nNLMX8pFuA6EcdwuI8WYjiY6folmssEWLeAZBois+28lB/KGdyhG5PfgNPkJW2HUsS8OvxoWM2V
DIRtK5yFFkSrFWNV7Uuh7U4jyYSIpNw4oxyex+mgrgPwkCVboP6kxd+Payc9M6cRJWSSn9FGFUU1
7oVQzfJBWIFSwaysC1sQUbV5f9T27r6Sw60d7nVy7ZwVaaCVyAaWNBTMSqaAJtl7H1Sx5RHpweY4
p6wVfTra+n9f62vgKZswTlycc3ZBZnWo4jeremd9r+E3H6Ueky/RiZAGMMZ0i1UNk2lK+5R4adBA
JR8vNka00tZin0lM81waRthvNxK3E712BswXeN7m3kW2fQBzVc0kSsRiWjB+vJsr5gsMXKPMtmJ0
ZnsWAD6BGIeqPCw3xxiFLXrpmbpQn3p+5wSQOsGmwx0IKHjcwWJsiGLApbnt08HcfYlKA71lEfbp
zQzaEUrwzSpajfP/adXK8gawQ9xuxaWagyJQUfPoq9gLd7B8N/S9jbguwlUdNfz/vCD32MD7CF3n
juWY3DgbAUSbdIZLjmz0Y+75RvXfBplzSYOv3hOd1EpTwN4KtIZGlUYjFff+QEM9sB7Zpm+Rw2PG
c/wfMxuEyHF4OSEDiYRRqjRFWF8O6sVhQaE8eJ/AeJ/pzje3XjAtu6fLk7y1l3N1aRTUvaYLyQdf
EzpaIC9ID7QGo4Zzxa0LnfmFvTFMwaOHJTJ6rJ1uE6E/w7eEB8R8aEehoyF6m52BjssDk/7qu/qg
eCe7kZpTo8Qz5BZZOPnFvtcvXKGwbpz8od7Qmt8CGGDQW3Dju+VxULUl42pjHVTW9+jwXM14GuW5
IxPMbE8zZQpW03jRVqZH+y4uU73dE54r3Wp6BlpYsobkxYfqc6O/eOv0+sPcM7H9Bw8iR/tGQicM
GdPuHSQk0I/uTsWFEHYZYon7e5MdJSgXwJW79U4B3l2QR/nr6l4zl+MPQa5XD2nt9l5wPNdvt42T
KU2HLn8VzLMCSxS8HSQlV4pudPdDWq/JYz6HkF2GdSIEj4WheFzkYz88RTVq0BNqK6Z2KiwEzJKP
uwDRJy9eYlHOA8LdhU8/8YmoSWTOMva7qww64OkcnOIQpDr76Ybhvk1ufLOwm4fhAvpsg4F2k2hY
5/Ffmc0rMuxT+X8TCuNVXp+RywKC14wIEp2h2hFyo8/t3NdIvJ6NTuS66FTqv9v2pqErSL0mqml3
kLU6mCYwpyjk/7ZmHWwgl9h8oUUi2bp4OFTraBUzS3auOGns/krKZCXZv6ylomlN4rhlj8SeK8qZ
F15n4Si09cgItkIqEYBuM9wvuggyb4HgxoEP87d7yMUMWScmojQ7pjwh605n88siBuCmdbyyJEWo
EDRQnLKrEi4UwRgdS8+ZGveHBhlauWqBDKZchRU7oiZ5cD6J2qxo26FGJR63PUA/QSuuwb8/OVJC
3ITHQJF/gGHsrrEm/0L6FhM4/IEH0lojtUrDdA5L13vB0fz0RNUvxfc21/vqAcC//oAG/9w/iddN
iziqmlC0dV7M64x6rwf9jj2spxmEQ/hwUrqU0uQsrgWS6zALrM9CfjxaCSRWnRKbTHjxHh9EvbNq
ufyRh6SLJjNG3yxwuqr9gs8PPnEFZuXMCcVfFRDyhEtOo2ZmiAsWHbzU/BGthf/dw0D+wIqx5W3i
SQJAA82NDy6+/IPfrbYMt1dipIZKkA6f6swp+xEXO2/xF/X4EAnglbrOx6ABoOS8VvHux063z/QS
QF0v51sh+5u2SmfwvT+1qUeZXFlJVa0PADRlBcHBBaMBEuq6ILxG/69uBdqoM7NyduyL+3i9wHH0
aBoPjFGLX83/ySSqWr3naTbLAt3YTSwiu38qro1XU/q2y7Ju/frBhriXq7hBZOPQdr9B9KpDrnOe
JTs6xxfZduNyStC/yRGijA4d8Uv77Aq7JFWcVJVIXCjOy2WPCxMJVc/LOCjj29Ob7CAsIPnH4MXo
QMHaUH9jr2dI/36ATySyaeFbsuMMHvtDe+iZ2uYu+jT+LMck0QDX3UZNZqOiu2d2R8R5D4cxKS+m
Vh6+D0NHU6KpvAQHFMVjuswINyyxpPgoVrF/CVysNm1WY+FdYD/HKcNxxIbUilPhPPHbOzaX4Fi6
MwV162qPFUi6CCDSYcJ/At+1P3HoxqN9HN8c09RRj3RFa6QmKeecjAMheSP/tNx4wayWKzS8cH+k
41zV5sMV4heFybkKBVBEpYGOx1J7UCQIeAM4UYnehDo3dLWnnetahhvh+BFWDxO5v8k31WBEBECk
sp6YZG9nHDsOMj5o1B2+IdjVY5YrlwfHOtWYML9+lcdRyYsuGIFpNk+n36cf3GlacNmJHU/xcBis
7KkhvqT5tfEAujoJQpuh3l5gTPMbTGnJ8e3zo1jf+bX9xFm55It7aGDw3dIYRZG2qmz7DiKa1VY6
eppAQ8Pq5q2/XS8yY7QvhOr5hX94pSbK7m701UHC8pzpt2pA8lGmpU7RVjAvdXmUn9RfIFvFrjgo
46Yf8W4WXoDy3ajrlZFdmZxwgQ44/4fJGVjkzEz40ofl7J9y/VdLlrfX5DfTdlVR0zP4tfem1G2b
MpAgUN/gQ92ASQZMdqxegyOnxs8vhbLDFm+wQP6sbCMnUXWRSHIoCFvrvAhSY7RYT/kaXYH0NUTq
t6c4NOjLX+KCcQLEqLmGPm7S3gyd6+dT/35JnX+Qilj5uJnAMSrMNiyP0QEmpzDpa6ihmRWCeRTV
Dm66x5tW6pjhEqkvw7p+C9gnzG2aBFMaU/Aue5UosYNEbU11LRpGSGJE64aLqYfE/ieEA505xa1S
ye8HfxooFBWTfyKdsUDo9JPAXlKJFV+LwaKaOmH7Mxj+amQhZqD+tNQzOEQF+YU+D0rxm/1GFv4N
6sjc0L1mr97s7gBMDZ546SDOjytmIWzIKq2ZiB4E3GrpLDIgY0hZpzc6JsCyoPSqzIjwnaL4lYlp
zypb2A9ILhE4ZnDsinoVe1Ycs0WN44tyFIV++4Ih6P53Eydbg3c1DGd4uRunKyzEYqz+4T7anIrz
Y095fsZ1nPbzwIEdD5Z9cNWebDu05DjURfGJy2N2dNUs4PJTj1P6IeSUwMxMFqJwq99P+6urOE2B
uWIlox5Vbwxg+anKj8VdQOG5IPBtu+dyhMm49feKexn0kEpRF7tKb6mQeliSFPzLsCeTpVy6YCse
VjUPnxFWJ83pt5E2AWdTlUAB4NlyiLrJmm+2mCxD56U6VYaQnYhI7GAwPCCPM3mlqAg3VGTYRBK+
8e7i8zDt8Tcl4IYV+WRcV9TULolk3g9kjxSer9jP9SzEZmanDJzYVMZUfxxHPgIsFYWw5Xsh/Jln
Tt5TP++6fe7ZtQQ7Y+g3gj2bcvNwCM/Ydme1O4BnpczHL4xyOVunJdqOqiz37YHJFZA+UPis2NhT
QTuFwPKrQ4Zh+NPU+a4LHuyVpp+x3yKD3dCsowo3MjCn/VzglWiA3TxxCIJnn4hlwLVGe3F7eCj2
0r/T9jdXP+5+kuTQ0lirOg8/EprYR5FYSgsp1Hz3cj28z+kV7D5NFRG3gbT0LKE1SPoNRWCLvkN8
veXgUYw48G6WXPBV6GIb97rlXUiZ+P5UoqjqsoE/dFxtNjrTaU2x8YsOy9TtoyVHe/05Fd6MLxJC
nt+BWw4o8jC+keqlzQkX6ZWyQq40lXT0j4ZAim3gc0YrYaK/4nbxkw8zCN0+Mh9s6PxuiSe6DHqG
FV/x8MzI96GV1Dj+tWqZr1PRb+nntnC+k4iQrGnpoUiGNJvWIJACCaqHZqIp8oSe9Erxe8MRveAU
N/t4qkR2d3aYuk/bdHVtD8oSd0DIwir7bV3at2Vf5LrRQLurYUij+UBei+ihLpm+8t0nvrKXIPWu
hXcTD+fr+CJ7YMKrEfQHjqgKHtVAYS4T2Zn6xCyPEfyByAm930YcCzocI5ypfmnr9xyOYuog2XzU
m9ArkxqPIboume7j1jKhbT+fXDrFLAUwijfn4p8srrJR6sGjuL5q3iWY8QOCjoPq9sFbnDp+gFHR
IOv4y8KfwJQ2w0TVMJsTZqLrTX80Xfv+jJxGqsGEOQyPP9GPgQav9LMy9Mn42N6Xb5ilEcn+Wne7
UMcGrm6nwGpPQXt9dWuFcmXuGRI/Ft5xxSmJwVxSkCuTo1ldKnrhOfiqIqUVLxL4RePxKwN7AzTW
98gOQhVKRk//9DZPGmMCpCe7eDchD/MLlKbx9mtR6aXS1leicn3TjJeGgfzqLvOi7EmNImagNxB+
DTIJ3V8AghuSiYmK8RI/X72ueDXs5xCmufM/iR0zj3DcGEtNIh6m9ku423SAjhQdh5XviE/1zEYM
fBZJDSNrb4/5Tq9n9In7s8WlCm1LIZN7FfSGVoNLUoF3AWT590703NscLFtqEcIFDGMPPAjMDT24
1gIUfbiJ6HFMy8Y5ChvLGfetudJNI4bR9Ov8cyUxLyDe6RM7LfWLu9v1XMz45dEsxayuFD5rMeCL
I9nmJjBpk9HPvND6Mcytzansj/l0yJMc9Y46dTix3mto3+yWZ+j6WDzdaxuOov3r1DgJ5k+duDIm
IGazA2iyVaT9mEfDgaANQo6oxzoTA6Vi4yzdI1NhxCMnunG7+IerTuQsKCoq11EA2QJqL4+3NSd1
nrvmxEBj/WDq/lYuD/QJW/Xjhc4qCis8QKKfa10VJXzSAnycWARLa4GujskikUfR3yHX+G44xs/G
t2qcrpdOPNND/Ljb6tDgyAGCV7ia61xadqGVHHkdqPjKCZaEOqIXqDlTU5MgkGCwnzj2zH2rJwpk
TPhWbePuI8ZKMVjJ+yNlGQzZpjNth3tWUOb+WFbSp/AZ5Lyfz975ttcX8BOic8XAhfILUpkQf3Ni
Ekq6daaudvouhk1wisC+tMXvJWV+q28gSz/cwtFx/+IjnCh0irtqofNmbF4UQVMueId0M4fRthzI
sXRPJ36VDk1fBte4j6FmERrYR4eENrVyhKC/ihOdukwRS8iPl7QHOLwy5uJkRcW5jz6U+eVXlRCg
RbOQPUDZZJkfrz1ibPK1dCeODbYIMzX9onA0TeqvzhRBd0QtE2tpdrHQ/fu/HmSgfcxsFyrO7MAY
+QYggcWREfHSek1WMJtTDoaTd7jViJX1oaB86DXIJ6Nx/osc366wdia6Wqt4uqyCFX4pwqz536DD
4mlpjMf6Y1xTm7as5nAbpYwVoZbq9Gb/N9OsrXRuie1FbLS484cmdzmm/6V3J5e8IAMLbNDUbhU5
X/p/Pd2dCUeft4Ldr1OW1SqXjU7UCIN1QONcZ7YChBXM7I0cFuI/4R5gkL36YtdFyNWmalOjkDxm
U4gZ96K8ZxyfQ9oKI316ruqZNT5LWHvHzh5b3ljIUQndIpkHLMKN+C6kmjtaxNJHzEUqbGmUDn/f
3SWVP9+S/p/6QIu+xBvkQNleJ6OSiIeGozT5B4dFC/xaIf+Ud3t6qup7bvQiTnxoXOiM6eV/rnt2
DIh/i9rBGri6d8w5zFIcu/lOX9El1VSa+HVssm+58MpyxaN/a7wJcE1dIUrvWNewCor9esvvmTUC
IE+vQNhTNsK5dartMVVJf3KV+J/1XEcnrtJj0ZnXblJU9cHeqUWb6+suWktINoer4SxNVaVtgjp7
/U4GEI+XM6W9HLHYVekNE0DQ56Uei6RbBvXv+5JwvAMAU5AqZty3Wvn0hBoWr6L0utQR4Y5Jca8i
CQV66L3knmoJ5SqgMG7E9HYpIt9a/H8QPk9nZQf7I1swARl6f7t56V6cacTY3GSQNNIafQZl1CgE
e2dYZ/9JIT7QN44sLQ/RTy5J7ZePzczxM2++Csm90b6CjMu1/F1SqXeQHt4Ks/ouJQ7MD/naHA0G
2rHyjymM26Bd9r7z9jirJn3sjkuNzzsgte+qx6MYb2Br7evjktjEaVfRTQHgGPLYiSFjkkkLQ5Ff
l9Qwm7KbrMfKfUOAZlwTP1emU097ooVghBxTtxPKMjtc+HAyMkaOtftpNm0EYd15AznHnvfT7/4v
gvSq7A6NlXUwXv8IDHMokOI2DuTLtyN1ooXXPyNfnZ1ASf4nFcZHq0vQlg3b8Ht/FcfN1lRD5GrR
HbqMJlWs6xvn0cvi+NiOOEXma5KNZ5uMoLCsf24z5KWX5+KKUpoetwFEgQ8+FmL3Vd5bX6PlcpCD
jDx2m8G2l+e1mBAYGA69YSAIGv+Z89gdaRhbQFYR+XfvcHZjmqatGhf6xLpqp/UpDP70m/MDziKn
cQVftVykTbcL8wNag9AC+vl+fSaZwfJ1cIIAHHBp/8gz/1PrSQDv2xEHP/hFF+ZxKSlA3IcoeZdF
L6WBQV5Ftn/kZX22w3WB4pejy5pn8c3WfloVoBdLr7SEOJV5WcOqg+lgb/Qck8qcwAMtXnG8A1VV
W96XPiid565HHlLhgOEHny4JEotWxCdqPDUg3qMqkW5zShZR7wN99BtJUfEFoOcG5wkdZ7yulaIX
EDsZhlk7U4rSWZqFrEFPWOg+NqcVOHjKDHonXhuCXby+OehHUGBmmxgG49WTyrO8criAP3WtjY8z
dPidB1LDqQLv0qHJdnKopZ7qhPOfWP7h7m0WpCmjWM5qGiN0LAu9x8ddcwgRAcyqI8OJC1aqu3g3
4unzrLtkXRk8NV55dqjIoZzsjOoz+KOnaEsPu5jAadq2uzv20qXMXIGXI4cm8wU8ZIW/0EJ4Wfsh
LVDH3U1pmYKR0RSltdU46sBP0VVt2PPmU+HLrJlXhcx0BA/4zxeB6748iS7KEVOyiOQictChDTpo
Sanr2dPAbS+4wOjyyfZgJA3MqHjMf9IdCCpdpKeyeAG7PnS3fmR588WcaiVEGgnK1+HdvzNemZ2Q
lvGGSdlhU7BufJr+S/oheINTQCL4sI/mQbAl6NjH+mU3igKm7f10iqHt7Vk1gG0XJyFwIK9K127u
gZ/goGMX/LSZm+ZubrvjcC3X+UnlCSGvvdzuZabNOQ3TQfXGAf2CW13I3+BMsUz84/mx12tFqAea
Bam9OIcwRmgecls8ywXIM9FB9UEqD4suJqnaLTkLvNRHfm97VJKsVI6AV9z4uJ/QViCLzGlyyMU7
er1gYZoMAmNJywHrEjSwYQL8lfvwkFek7m5LrR3LyuFkJophkqYIgSEyejH268LXredVgiX2o/e3
jITs/MxP6bGq2kqA8LTfLW/pkS+LGC6nmhdhnfKN9NCvaWKBE0IAiyVk2LxbtFtFzbBsuVzGDlnF
EQxQ828G5qwGAWLxC6JfDsluvdWTiSqm9HeffThuYyPgOnveZpFt9/j4gDqweRuLvwgKo9CcVw0K
Se7q+kel4WFfwRwK2kBNCPc5v9Cuu3poZ3+Z5GVIJE8CF8yvL2NUtsUkqCwYTwRt6LkhJcM7l2C3
Fy40F98LVtV9vQ+DMPMDY17alnTWRr6mOKsu4gvno4jhWXx/pALN7LRKbO6RViec46Mjd62JWiSz
AjdwUn5Jmh7KCS/Oz6CR4krsdpBMrKEm0wnzEkLHSptrT+QBus0sgR/pwIxZuMLSjskGuk0YmLOd
kXDPv2l1B9W4yW2GVEBvRy0Zv+yuEk8ruPFKgsJ2uJR1yYdkazqm4/S/AzO1fgeTHC9nAbmp5eqL
30rGM5fgZjGLXtnhQyc6RqEeZ7scM7ITC+pe1aDquOGIePeuKsbUpeurEdF7Qw03Vlxrq818wt6y
v/3KawDbWezj0i+doHYllXV647vnjxYy2j/ZqrQA15yiJN2m97c9zqWoH6c6eXCKr2qrzBAl7pQy
Gs45DFchyKGaPTPvipHoqa68U0RfY7Kmr+ojzOM2P8p2rczmLIeH0sFuF5c489azA8CZrfeJNX1H
sbB6toFOAU6zjYAlhqfEm3ShJlmhkym1kDuSBFOWKLm/Ijy6msHKdjpTtwCamKfvJCmK46jL3r/7
nxGwtsIi4j5kAuGrwEUHJAd/kr1FT5oZcsLIzlGeOXV+4NhQ7+MejTdDNtgLKMhbtNCXNEfv6ptV
+JUfgHV2ALhTwQHxsmDjB2elTxHySPWGf8TFR56AzHaU31WfmFcwcj0I5m55Rl2an23QHhs9Rqh6
RDPTfLSaVPADD7rNkED6lBSs0/2txdtrVed4qgoMr9duHkPrB9sM4syIv7fQ07wVtpXSV4MWfsJb
TGza0OQxC/iQo/3Fju8H+aaqyaJEeWwqy5dfRq5ozHUOVc5tDyJao7BBJURu5faiw/qejeEh87jG
W1FlxPzPwuM4nhaSnQSyWbdt9SDh0ae5p67X/UItQs9oSpbGEkMPmuqk59xETP7y8EKfL38ZlvHU
HSLS5hqSNd9V9AZq0ISyBvKjWSllTrlYk7tjWk5GTZjcU4p3hUrIUtpAxsn/OI+QFodjCTm9+IJK
qfPBZaYI/N6pH0sSpfrZ5ofWoWLOhXaCxAQZkdwepBFP4SCemN2htRdoK5yqE2HAJl0T1VXfSyf0
vt7QrB7z+N/XGVHkGi2Ss+wXay1Mye+bzb2hOQgGO3JdSGl/4WNFpfycJghhnKnoyh8fFd2FDF6n
SMpVJhIbtNgX8fIVEvlU2wOnaY8SEqYYum5Ye588SqlXMyjyKu21jQCrSu5taMoECYc9OQErdEFz
Or3YacRREM2n4o8a/pNhJw2Ut4bpfqmfrlcFzOFqSL1++u31Xt1JTNXo0OV908x/Jic+/8oSxxKC
zEnNqtzqotc5iZyOy2KcuB/jUR/ah1FMECLrYUUO4DPjAsUsrvMiMI139zTg6NOXh4W/3PjlCjIy
YReLKPOTQp86wnNnCGVkarPhG4lmuQH/iiyRivaiQXotrQzX/8JGd9M37V9BVnO9ZWrDGszWUiZM
8pxvf1G9RJQt8NzM0I1CnHIJB7eiiAk1wkM8y6iHz4qQtpK45vbmUIXnkV62pQPvSk7G1RewLpJ7
DWrzQbX88ZuOfkNYS94BZM5TIgxL7Cd+HuRdSVjAKNdHEYsQcARIXuXtoE/CgJvMwbzOuBs4nDhj
pUy/MHQ+zTTzO40QFBzQlenrDcLa0y5FV1lIQckv5h1z6d5ZFfLhYtJpUT7BG/MAJ2jfmHUtAwGS
PzrQTjRdFkxZwj+0go1iJik6n1fkLuC+CPFneEPfUHYcWk28L7HEbxaNuaTZFQGmcCU+PScoW0Of
ewlIsc1b3iCTUjOjEY4+h7gllaheke9l9E7jO14dm4r8VCbpAkh8R3b+SpTDg0B4nMZTag2Cr0FE
FaZVHiW8EosJI8d9hkGUc+FaygkKtD0k2Rf59h2Ow6e6GQFVBjOPHkPNnJTtv/3A7QVg4DTd3uqs
FzgoZFpO63oWir/vmBwoW8PXBqEokya3TlB4bHld6VR91hnFE+j7vW556X/KQfjbFGdCzqsPO6Dr
IGZiP5nYqYFsIuQ9mRRxqZeGT0WwXRH+vDljjUTR9aGFkvXN6j0P7CsfnWpG6OLAoLqH6sFlEIis
3LDlJ4h17sjiRQrnmCjmDmwOuF4PzAWLSlQtxBANAJ7uPikdgn+HIr/Y6V66vnRlQsGS2oVtBtt2
AVdg3rFb/yIHgQBez6KAE7+l/HTIc61yI5B43NWb6c3ocvDL0qFcLbje0YdDeyYhEC7+CsAlW+PF
9w1TfPwxRBUwVtWnAhTxLLAatWG2n9hQnQTFi1mHB4avQIR0q99J7IT4wXVyJ7BVpaV0lUjFxtaQ
vlfU8ETHraKwCPVpKwYZ/vZLXiShBezlAwSutob2t6+ufxK1mQvJwvFCUROKfcyRWLPiliv/LmFp
9snuNA+98nNBUEnrHAvRj8Iykwq07BsbebYBBl6U/Cl5SeSGeVw1d3kom1cfprZCTpxTDzt82IfA
HtY0c8GpEXfFvsks1mjVD/cI8T+COyJE769tnsoMcbsSzv42sHslN5uqvaoEh8m3oXnfaxG3owBm
MR+oGtQmh4AZcans7m6wFykenRrAodxqnil60a1i7HfKOOZj4nmIvgRi4uxP62J+D0bb56t2dqZ3
+fXMFscND4ZgMYRDhtUFqfgoXIZQjK2obje2Agaa5VhdKJ1CI/xfHvdvA7JKmTm/Y59aPlKE6WKo
I+V7YyBsAyX4z5tH0jGSqHSe6/5zqZZxZfXVzRsVNscith3VJHptUR/m7qVr4bx2hCkPfnWuaTU4
o9WXaihzBt4NFsSBI6wRfpBugO2hE/EcEcnCbZUoxxhbL839GshVyDGEId7W/7i61oiv893l9J7y
bKbDbkHZIo7OKoj85vKpQ/jcD2uokA7bsBYFlX56OAaQJQndD0BsPZru7PrTTRCxv8DTzd//rRF7
KoxL9qrstS7K9kYVSIG/xoIyb+yIVCWQDcuzCet0TwhzaF/pOUNX7oqye44n6GX1n3b3ucdWKM6c
BGQjkUbfkN3LzdTpMwNfCyPpX0ANxYkm7nyQz4CXqDbXp9n3aSRNRPh97iuYV6R2IVvpkzcSfOyC
fozw+Z9QXnxl4+ig7VMxv3XhP0tRcgyuNV05gHYJX9f1AR5E4XXrkfc0k4WNYfA9hoQ2edPfcVRc
q6akWr4X6ZE8nlQ/QYXvD0AmkUIzWjAZGadjf0sONRkeKo5h70UkP3AgVS6QsWUr9X+LPaCpg/yb
hkuu9SltDLSDoh2rmOurEmKTWB+8tW8tzK1cbd+0tBrp2RqCPWxnyyBg1I+EAdyZUlWmpBg9b2Vv
zL+00rrf3ec59KO94sADx7lTKtFMeVE1PWHEr50gW5VYCpuoKVyLNr2WxB5APp+c63lFrUZDFw+U
vPCp37N+Pm+rT94ahTuyGhHX/uqMoMHwWXx8uJgJqnNthnB1IUQmpMaWu5pvAMnNfdYdWHEUax2c
3qS3MiDzmYUxS/NI4/UTXWMTHnj37FFUMpPejt1mQrANImK1SjWcTcNx20EvOq3y4xi9PLlAU3zk
Z2tVsn6hnLu1haIV4QXzJRj+CiH1iBiVHhlbXLDOH1dI48NzS8zoWjgjaV+Oqr1kZenmqLwRQrt4
FWACrnjpf6oWPNRwS/sKy6/3tjtq+gISOxFPp/Dg0Xw+QysEVmsy4cNN4wq4Ue4Am+Z3f1zRZOGr
QMbSJd8w3ak6S12pBzI2Ax9JWF/aTB7w2MQFYYo8XFBDB7opx6algRZpVRVAtma1sVU0WMV0LPtP
Bblsm62mGkNXRSMNAACzhFMejRuqAJa0OczwiQCARhOJHGkpSlKemV7hIlSxt9EYS/K7f+uNXI8g
GtsaYNx34PqHvnM29DQv4kZ/fDLmFPkQuMUi0hWmRlFzGgoCeN78YM2YBl4X7584EITOpQkK1u/d
jclqyAnYynWTHlTW2mcIt6Z8Np1TLv0sgmrOnjAzvZmZ4jopPaxVWO/N617yvjxgmmKCNVtmu30K
Ihn4yCSqciPiliCtjevUG9bnp5wGHzNtPyFKJZcpMg3Z5BM4AS1icNmn9Kkh9EDQ11UdyzXtLqkn
0gwGnLqoTkWbWOkqND2j3jY7lU/ov6RNV/yEvodb8hAronRtG+k6xjyuu/aLJO6TQv2iRDyTwI2c
4mdrxZimKUygpMzx3jSCgkR8qAQk3B6hfi99AkCAzzLLaCvsPeC+mtSgj/vZ/b0RqVoqPVp72ycV
BdbKfVZdZoweJqzXixDkQ0nZtuW7nmae49qE0EofRmlqEkIyc/G09IWaDPwsypq+oShWCj6fWDj2
kIOr0ATtnGyERYf5/8J+Ttf7Y5JQZgIUh4n/Zvf+9rIznii3QFMl4VzI2Q3PLW+3wIOZ6ydblVm6
1phtZNwlraOsBZVJCFKxiFaF6tB/tNwAxAIMR0ASSFAOi4q/WQje14pXQ/StrO1arPhgjpZYAG77
51KePivNWOqFagN7Z8gG9zvTNOYfqDYTF5Pza05orC9xUYhauC/r7c1AgKTO1dZv1YKbg6zlJo/G
YqHZvu54t8B25ag+A8qsujvNlF2YS96GXA9kfX/Q4n8swaqd4UNB16hlJQrBGAcygdGE0tXopHG9
g1ZTv51QVXkqjOjqhDjceH/rerHt3I1SFmc8tsaaap6ZF6xqsnViP4JXoEDfwcO3iG+VWPPxzZ2S
Hcw7F0PMGtHNHW/V1OiK5jae28+Fu7gBX1qsvs4B88kD53c1QUFYHRyZIxXkwO4wcU0yzBRL8MOR
GxeyTMIsxEMrYE/bJVEIiherMLSgJjMBGHLr1EmaM+kl/xgRd40GzEgOzMz0BHKw5ve9lSXY8LO3
YPicvOxeVMTdVE0KuJY9aK+vSePftrhG7qTzDQBODz2qvAsXcmOrg4nYsgsKX5mCBJHuoznx0Wtu
CdSTZVn7jLgn6YNrQ1dHtrWqIncZwqJ04l+IDJiM4pHHzLTT46vGYzpUsKAOOzUVvnq4SgZu5dyR
aQQMiFuZ5Sd3VmeUKVAu17XHh9X4NHGLzj6zxHi1SJmAUQVJ2+eHnQf05KgzkGhSxz6bkGlXhrfv
lTep7z+nrvdZUuVJJCXwlrouvfAmW6RGCBdyU1gk2f8UaPjbgy1E8uINIvycZCLGl9wMeGkbO6Bz
ftObX3gHelz1cORXnuAK5WpJca+rtgwGMdsY3MFHFWv5k4YJJ3s/AHBU1l/IGn978tMEKxKwYPJW
988sHpFzCDE6l6DSYb/TDo7NUPjoYLoCSbuPPV/o1q0eIlNHaqTLdripGIrWpKVouaHPNRBeYZW8
aZ2IVYVLUthpevf1bIA5H9zvZlEZ0m9nV0Uzz6DDDkExgcvukLoxoUOaHyNjzODyJLv+eNtopVaJ
AiHyJdIR4vKWR2WG3jL/Re5MUoRimbbdsHRlPS+beN1D/+Lfn7VcdsmSVsaVLMlzGzGxVQjsbNcI
PLA9o1lj9iSLUUUrwo5huGYN9+Sk783o7TBCKhMTNwm512dCpiUQ3ekTfEzMlVcwt/KPsxWXLf1a
1oNybGqW+KlocG89gg/aY4g+JEPltLYWU6ULVExaowySgO8aitY4O4gfRs1DwhAR+8LD2LcmrBxx
kRWZBVSzd9f8nM4UhL9K9Bm/hx/SpFt6N5fRmWx/YZ6esC5TDINMraItO99Z6bCpDpYIufYu0bxE
qlnqkyjIN5iNxgF7uYPL5139qMMqDjUnkW5hfLD+Rvz6Ct350gjMNvv4Vip7is3mXwayTUC+N5mW
ZENtcQZG19gHAWxy8k0WaXblXmGs5l4ZVkCJUSKSQ61mP50Ro/YayURWTd00ix3CkbjRDhb7ADec
Fd/YMJtVxbhZs4mzR1EJmrrSI3Q+RnyZE0BxruxzYxWakK+hVCNUHDLesdd6grzOZ4rUt/gUh+Sz
WNUmoTxMSzuE6S0VsfL7ULc4Af02nmILpM48fAWAQFbfhdJRH3pG81r503p9n4gtJArtIw18S/Y3
DiEwcpE+rxOWh/W/QhTdfVEnb64YgQBzkxfehjqlFGJGfHlyMLltHYAnM/XF/lhDNUq5akBM0p6z
J3nQQpksIiK1RLtE+qTXmRBns+YwKQEfCkx7MioZ+1xXCQ3svx4+Bx+0QASl5P9iBXHDdC2vLrZl
301y0VB6VIJVdAxtla7982sD53KnahChMXtooeeAIcr4RvIg/Ekjj0ge+eTUj+GtTdiQruGb01T5
3e4y8Sxh6TFakLA6FMDMVoDnidtHrBk/bDSmvSJ/cybQxOlO9NNlTEB75E4aZI6MQfKOHhDes4CD
PGTZO04+CchxiyoyePLweC/7QY92igT/8a2xVewvY/PCcrBsbPr1WzbPfg2aJRhoTdiSitVrxmBq
5xO7t3GxCjLHzdEcFC5PG+DQZAR4U+KwkikIaWY3NxWTRO2Wn7R3GMNDQcJ7IOLYy1+NOuJYmIQc
Shbyh2aitjBWhgSO2Bupqbi7N6LvPsLCJXRM5BzZHr+n+l1srM+NSjs+UtKPgz9LaQm7LVpoYF4T
WbEd9qy8cPl4OdLnLrTkYAMaSn9C9HKffURaHwQW0p8FspHjDgMUpsKX1G7OvE7LXokbkv6JuyZx
8sLYsxJjEFTVEkMsJ5t+r8yH2zc7Gt6iddKnBrfe/0YxAWZg+bdMrCS6/1/y4VzftDVRBWikgKMO
yt4rgECcIwhy9Oqu3w0ad5I8AmB+kOaH4/5Ej8eVFFPqynWigVoVLu0CzNfftj57u6aC69MahyDj
gq0qCQN0mgt9+lpCemWjcZkb0tShJ/HR5vrFFd7oZWcJkg/AYQ/5lxS9lNCld/FQJ/bkVWe890nC
Y/9Nn+xJcOIEB/EXboYH5sp/K60OAZkRMQZq4KjkIregCMXrLhhtlcu5OVOYUGEpo5Z9lJ4UTwro
NKoBO8yIhDtpyLRMZs5U1HtdHQ8HT1x1xtK1+94RgEqkNFK+AouosiGYlDS0P1ll0y9shKPNXKSF
hyZlyBM+O3bym7ZuhilFjcF4h1uhNxY1hTQwotWCAzKo8XLUvQKEH1xBAn3qye2I8dxksHQRLIYz
nVcdx8BvSrH5cV+hEz5Lf3M+aZKmk8dPpU0IAPKyc0BUppQYxCdFT9YSGZb8QIjtyNr4bsQ/kl68
DiwRmgXT2O3EKGJ1wwi3AmJ0UtcXa1hMQzZniEq5KCk/8lY33vr0UtjCTfuxrhZfGgcuiE3P9GOP
lniad2LTDBmG0m1IJ4fvGrO+PH2m9NPti7mmFAvSFaGEdXAWRwcFdQG4S1R3fOZkfSQXOlUyiT52
zXMR69+wKApv4a+y+q+ppiMr1a6KG9Zoa4OFThkOxqExn6kj2lMEr2i7V62QOmQY2k4UyxUvNuSB
J9DmUdLIu+P0ZFzgAVn1W1dvGatBCZzJJF9qCDcicFKnV/SqlFMNQelKyLdqVlWgJvmbeZLIdU4E
mKwPG2PFzF58OQzpaG0B+XUrn35lQRli4sA/dz0cRjE3h3TAe0pv5dcEOpGH/QbeyfQ4d0Yq26iV
l0ahm02NTl+pfQwIV4GkgI3C4XRxm9ATDAKcIFz4HGBKOxNHn0S90yq6SLcxcGt+XwdIVVFM35XL
sHNLzkHc8ESRzh0W7tkDNuxqtrFtNDv6wLmwHWv/js29Hc+OYEGjsUqQJ0wbP2CN4QrXmb91KymC
mj64TQ4YV1rJW12y75oMAYtmwLUNPc02Sv905XmBSh00TGpeZ5RlLfe5lseEm2/QbTC6JA77Hfbg
VCHVLwB8Au3pZb1DxQfICFe706RvUE0PC8V70g1llCeXYGps/GHSXArvhNjrZF6Y5KYsI75fhhGn
kKn0y0BhmJ1/jfnmYZVz11yZhVhryNh8EGiou6PEGGIq6Mu/AvkvSGU244JR+7nf++ivF5tDjr+z
Fvy9/7a3ARZiWBNCw+NgCv0GByoFpVnXrApC2+hGB81LFvR8uzB1wjKGALUzTobncaqNrkUUJJLG
bnBU3rZ1eXgouPalTfh0JCknGw2xvnSkiJM6A8fnzO9OBjEYqeItOG5dEV3A6lb7rIa1j6zDZ0Dk
nIv/s8xufSInMTKVcZ/BlAo+FkIENbiKPCSBKjilkTvriIcXWsDM/Bd/jbhm6lVo6N5iULv5Lrpz
OL6yyBJoGhTFk1ILoEr03GVAG+FfgKIWQ/EKrJ4M90sngj2JU+rFPJIYpnslfER5w6F5Q9h2G3oe
p0TbgtxRQQcY/9mwShpW+wNwG9y5xwxVSeFbgIk2iZBpKAzBM5mnTlsxTgjroy/AxSZYlGmGTxPx
jPXbhMEAd4OiWRvyklJ4VP/0Is6sjEE/5q+sh3TYwiQ2tEELS1o32A8VEHalZZ2sIamYMq+ZWuCr
w+DZ2lAV0nuhhQzm7UUKu0F6huSKfIW/87wUfJtayErLoZMdFoFN11HH5Qs7pzjyUiobs0U0N0WR
MO1FvLnYlVsDmAy9Q4xt8RDtaCEbQ3OWze5N59yDYWzmh32Pk6oxlDLdF8BdJTpO2R1iodBXI6Sc
g9Q1JHN4x7s81V3NmvXUs3JjJqM9ILn3eyTDxGevwrXI+Kyp7qIAv84gccCf05Z/jm0h3u6D7Bei
rpIeCPtchZM8hBJr+iHwsZ+IYjysFOEhJAY0pieM+bLfB3zueLAqPtnvjRQAJSbdUCzAeaPVyyYE
0m15ZLFwMCySboQIcbpM9GS6Ob/yxAKn9FdRZaWzIdJ2xdBvvfBe8pVB5b9FvPYQhHzjXtp/fPB8
ugxk96BHIKxhXYJkcNVh8zyR7i/jebwgak7vcxZPV0z7ga+GNent2FLoQho+rDt1mpC1JT0inRaC
KYuXGTDX/Rlo+V6vu0j/3AUQWMsInJBeHA6ZsJZ9IMFtCzsrEoXA6d1ARFXVg8w3Rj2b5SKccdI7
o4xdlbWPSZ3wj1AAsFjkWgHDR+Ft94PpHdtBzCTagSoMm9za63x4F4N5C2INMJfIOPNIqmSdzNKJ
a9jQc5WqIr3TV1cnmcgKAAOPGE+EJg5+lSRZRU4XXf3aLM8/WY5In/5/JgH81i0YuIxMErMvr8yb
Px264SKeFxJ7aZcvvDpsJ9WvTbAtKXGjCtNXJ7Wl4aD926vcfX94JqWq+C1ZyWQWDQJ8NauuVHBQ
wZ00RCgb5YKz+Wpkcm+hcttVrsl7FolWiPkCE6V9r//IWyy2zPJaPLOq3BIushOlAkrzeF+TTR3K
LhdbATZfE03LKlqg1nXlf6ym36JycfazrAOJkMWQR3NNWzeqnXjKowv4WlAZ6QYoMxk2ZFpbQYag
YPFgduqRah5Q8EEfCq2/ojv0cnjX2sRBV96Nec3Q0kOE0rRTVnsS0JgoFSe979MjVyow2dLslqIj
h9SY8OcmSb2OPJVuzUT/mo7aiArZnKROSM2OeCIo7/+U+IlYILf6yjQlqs9ObbA6eTmI5fhbRvU2
UuZ6vhbNwOXpQKfFV0F3QzswHHS3kYD9c2LkNyL4iBBAKFBTo+FdtcknoGPfehmzN02uYu3uak+V
86OfIBh8AqdYrbrDKeMSThgxD9J/rGTxZ0Y+dkQDrv1OXq7mJs4cG9sYF4BusUF0uEwoLQqdJlny
tP7TKTsU7RSXoORx35ZAixzp+Fhw/a/attcD2fTQpe7/Iz2Ks0hwzTdcOdyQANiRBPEr1mZBlFze
SV3QFJrdoRp0i/A5puhK/X52LnUJJQMSdaHiM7H5+MQ+9H04/otPgaHuyHVn4jSCHcRTWgSzICQ5
8UvFSEdjcT9Yp5TPGySVG6TGihBnhE4USWOxiegryqHox7WclQEuNW3ezs+ImXtcGpxMP91jtbqg
J3/ktOkjOhV339g4vVEG11xiHSFe5RtECi6hU7P+Ai8l8zdKF9jUqW1LjHt4d/o3hIEtxfm5btt7
2jCHab4p2306XaKFD03NsMwr81cLsKFMPODSs6uggA3SSZ0/5ki7iyMXVCS9oN0GTiFiueXykxrl
wwnKRFYAl/lOJi9np7kfTuwm5EZI4b+8qKkF3pyFGH+G9G0JRpu6NlALVBJpkW87GtlfVRXoPh5h
ieZG0HJ/z8GvosvmP+e/ZxCwQ3Z0ipkOmmvQIokRhtc9AhdHwoiQBcvmY1AsHlfSYDghSqODftyy
3dWtLHShMQjaFYSMtPfCIqzn6li52LPV8/c9pppmrtRoMhh4ZH9/O4d8yrIZC1xSrChwxKBwfjAf
t9QfX966TMU6jF4/KkfOg0aIh2nyHstX+vmTLZcuLdFjErV12H/G69CiJjiFanUlx+hBgQVFmAiR
SEILN+OyuAiMKQFX8wNoSwXjK2WjTREJ25duDR5tCHaX3RyFQ1Ua39cNDhClCykjkPnjXpQDzP/o
hHrQCDU0FSmyHIz/9Mmx0uIWyOCQ3kmmkVPkGHbq7SpHecG9auUPfgSco/rI3BAr8PpB2TE60OU2
m7a0YWCCBOrRX8rXtQKz5rOmOjCgNJ27NoyeznPDk284/D+ThEESJgpVRGzSbDCR1p8jR1yG877V
lZetpfJ/o/pPq26lgO2lH+v6HPdI6LzDx/K2+s7YWmhxldhAIdu+ZJxX2OuaxyD1B4XID0W7YrX5
zdw4xQvvopI3+9uCsGZeBuQFAl2p6N0qeMJd1XzCaQ8l2YBSk43/GNihbuxvLe5m7rgpyJJZx6su
Wz1uz+J+RnHcra1N2aQPeYEuxG7YoV02FF4PdXTwSu7kQJVpTMBs2LHs7ARVujh1bTko04RNl3JH
PlTfuGi/yR+x3/EqmdUtTnLoxBYkVwHvKAIuEQE4bPszxCm2CNrtySU+qxs5oeGxPeh2FT8CdHnS
6wy2UD+FmRkkOrQxXz4KT0ZezwwobRDjVA2SO0Vd6C3wm7/RcvnPUJJ5Um5bq+zIlBvMDeLV/sSn
GW/lWo9GbZbo1Ec2FYdnamhsQP2YMsVRavQ0q46hC8ZhUJBfkz931t/CUFTR9VY7ek/fmu1D93H5
9Bws9QD/Pgl0qi7M8CrAwNzTEXjcBEiDNTdHXOxJhEO61dU8VYjrGCqmFJ88F4oE9HBW6hnVY1jv
VbVNLo1F7qWGeyLw1DfMvJsdhrP/UmrESesDCA2Z4Q6Ftd94jz2REUP4Pxc82mlppm+EiRrloPl4
rGDr3B+IqCIoHt40aq2cM4on0B5gpzRzdUQCia5TVKJckQ04HoBGsTyzXkYre+YUfJrsLdGFpdJ0
CP41gGTkFUB0V33zGG4YgQmYj3nojz+5AuMQORFwUVdsgWmxHc/cEKwYkocvzuKotXNNOxquhVIw
QtdqI6J2V0JMK3oBOTM/8t1GxwyQ+fZ+xaJ18SVvnHVvyYS1gY0RJ/KMErrn5byq0dhzvRMZ/B8R
SvaG+7A1f19XBRYbZNLp2LiPOELolSST8ZRfDval9BWPks5dcbTv7oyY9/lkVe3TYhUQFWpfVicy
v5YH257lwz+HENSvq0WFsNv4PMvdBnIo1mcKyuY3EYGtpo7rv6MSchrgTJwLgY1stbSC0Wt7VCNw
nktXlwUYkjqBTuGjO7hb7FEdWD6yz1iHIHJHfVifkX768RJdqw2jqq4iWjKmUJhNrnbkulw6ww5q
nrT3AcHJ0j4NsyFGO042Oxn4JuU9GonT4tDH79X9cJZ//3xu7l9DLv2gTzcxPsKo7FypFBpEdaXK
QMuz6mRCGQ4V9ZpzjfxGONby4lK3olDt87bUoMTJGonm6KyvqnnHkf0YvETbB5Vq9ZFUc/rBLGN1
UD3+8r4O6myTeNWIsVn1sf3CvTNIJaaEFELkr2QyElxXbqvzmS2WTHUzmlYEWphR86r68x2MsdGV
HCcI2YtYgXBShmp4AhXsfE3OBypsDEGXHCbIlagRx89fgKOLIJ/f7R6fmOt70kIubeCOpZ0R/oZB
eoAViKvcgZV+PcynFa4+vrRX/hO08/a/udvnfG9oPtskxpc8VS4av9KROEQFqtJ5cpVwrzR3AiuH
qNRZl/NGlYrIzyy64AdnVtx52/D0uFVZ6ThsO6l3JeU0VFd18v43Cj98bVwuPLlDtwWLCs+FXVR4
wbqR/9pO/qSv8H9VmgYRndixV1ht7p3WiZ/XRqaSVjJ0gF4RI8IHdX1gCD+fnuc2NOAF/9wXIyGY
Hu7BYNbq4qxIiQdLlw+glSAewCfYTum8fhPtBn8s+fEw3Ln7+FvUtoPBFXmCMhd1KCi8O5YJ3eq5
RAoHxypRKv9H8lfcAYCghkABgBGz2+skkt3tVQYeK1x5omHukGHMyaMmO2+P/zpYwNZlBfxSe5HL
mR5tDoZAx8mgSqgA0TlkjGew2lXA/ldsyF1aePy4I+CZdHSj7dP+xvr40LjEfWswpDakPZ4miMo2
n+YUVm1k/r1xyVhQxn0B8149ALluG6hQAVlwsZaaV3AjV9b6VcicgZoPIh3Zc2j/oJSofq9zj+v7
bpDUofPv6oHpmj0bjc73NiuZOeoTe52sb/XN8dyWDi321NGe1XwUl0q/sUz0iiAVuYi55tvydp6i
i0laBZsVA47luLOzdoc67MjPiO/+NAjjiApOPdWY/FpQGgRWM+RFkGIwkV5Sgt9cui/VFb8e6tt9
5VY3K/5IwFP+iNOwfwR9x+d9z7s3JeY4/O4uGEZfIqq/JCciXVdaYi0XpvjXzfPMP+6D7XrEFfvF
ooVxwH513HUgGookJDLOZNvsr4cDOWjepvNvNxGbIlgwxnhLNjzeS0HqApBhdD0QgG5qyvmOENJf
wR5sjOOoVE58Zo+iHu1FEdQdAIwTM83BGy8FgnDQG2PcfPBq9QsfReipXMoFtc0tPzVVmHRxnPCS
V6oG5qmVd+gmUP7xaeG8/3wbf0qGJ1HmVVOkC3GYKL2cGCH5iKiNRFZx271tokkWyNe9+lyokzrK
ZZXXVYgyEP0EGOi8qVEU24BXF5yiBzlfEHCTFlXLKRI9RZH7C5BC5ST7/hu3zmYN9wAXN+5g9dBg
bJcbWdG9mJqT7dWmrW/raKsFNDJM4LinTm88TtqB3+My/fUUmkE4FxdGa+vszOjqhnz0SGvCXXo8
kAsSU8ORWw7B/Z4ec1akwgJA4MQEsm62ktoKr7+BWh22kgtkKJl23N9LEt/JfzT7/TZCJM2wa42y
/OTmAVTIR0/n9w8zfEK0714St1Dp9CeckhUGI7lOzR/kcM92ng6bNuRWhVQjgO2J+5iMaoWAq5zz
Xmj7CySfh9Bn3RrYMDAgJPHfqB+7Y28mVw5pBcVTMj/PueNfHBpYSacNmwx+vyDeJL1Jc7JLh0yr
n3U3p96l5xmluthR1V5XG30ZJjWA8A/XJluQW3JqSrAfaIOrzbI1Stw+kpQsFIjXc1cnzlKS8nXb
pm/ROaTuCg0kWEPoi4YxVGK4BfzWZIwuij41NklUyme4I+2H8sAn5dwNDGzQGLiCpXAo5eyJ3Uy5
m07QX0amqUsozKgeNmqQC04b4/2DYxiAGkzJW8bCB7DFkWNqX12/Ffje2ylRgDZzKqRx1hYQY9f/
zZiQjNvOgbKSkKPuf3+BTm7NdnPM9wXqD2r49yJvBml/IeG68uCq8Y535FUJVndhCYBRntWcPFRH
1OjBAHD1BTWHA1ktu4Un51uqbsC4OYbFvfevfP/ufGYaBB+qumnKxM0pIOCmCcYPuEQZOIuazjnU
r9fWw1dnAxUdhf+t/oh4ym7eYUEY3fad3B2xKqy/fDrMx5oImG3F9A8yGOv6f4oimbT3jnN2SsMG
K5h8VH1EdcbcIsZf7muStnu8hPMvfFMWZF2AUwjIdCUuGgw4X7XaPqgUpoROvWeRnotqQOc+DIpm
TUmwyObWCFhyTYQwN+WXFnShOCYjZtnjpkH/JPg0HuRY2mcjuSS+zIKCKHcw4aPeAFoLw5TQ7cjx
QrjIA7gzI3Z/stQe8mTQrqSNi0i6+jSGZRinKvaor5BP4Xpcxf+3pOVGYAeYB034uox2FUySNiFQ
G5bYvVNgPld9ywNyTi7as+DFGX38hT+Sa52aVh9A+6pC8tVFYUxfwJFhzcQkygeXzn7aftGQaJZU
rO2Vb/gCsCJvTcROq/Xxuajga9+m8XDCUOYHANBJHUnQ9/snV9pUXgPTiBCAcNstMFiF/efmUAoo
c7npS7I8t/KSOmI1LH+ZnzNtFsfRoMQRDPtTyZdBGX2T65TSMsrUG9vAMQzsoh8NCTsYWZyGFtg3
Ql5s9ddNkZ95ji7QMGJuPTH/MlsktUJihrsbvvbLVPGgp+MA3Y96mIlzwWf3c5Mh6VwSRFv8Y8cY
Q151v2EwjXGysci85qJ7/dM5pVjBIkmIqpDUkzKj7nLXSOyhAMZpQCuOPY6sB+q8+iG1DDqASluZ
SuDmsYZn/6QBiSmGLlisXdZz8XToR5KJeE1SoRbMMLUkJ0ws9HFdGkwhju4S+/QYWZzQUnO8eQzy
6XAOjz/CFvL93a4T6kM5V+SOd2CVa+0jeGerUKLNvIlDRqMMxjsEDHmvUd25aePd3DfOumf/p8iA
ZC1Ko/SpfoO20Rp+06n5VXAq2HBaKXZDvfzLD6BXzlHX/pyWNwtTn+T6aLeVvr/7tlktUBid/r2Z
g6UKEOvu54jpo9Bxxzc6xaE0gxGgKVQQv8VB1VuJ8BNvh+c5tZZBGa6AO4Miw9lWUo4aSqMhB9in
fFACdTaXEJG6Ldwykg/yqIZ7EGTKVWVBWweA50sP0v+Mb0c4n/OR/pM/fQVcLHU45MBZZXqmQQci
1R/3+ui+RX9+wiIsVLO7mmvExe7KsPMc+9g4oXe17KbrB2Zak0UdbQW2AwfMq4SmKTcQ0L0VG4Y7
PC8RzUSWEhZL0FAGKgyHeQlDaok4IS2MKx7XCQHgIC+KlsQYJ3JkjXgXS81tFFoHKAANja5HHQOH
IvO4vudChVMBg+GINZS6SZPv2YOZR5ShvwPgoxpg2Es86u7jmU2q3PhM2/Rs0dZxqknBDhgZzs5Z
g4VMocBv6VJGaK1TKRfTmyw6gmBjBwEQMnn6IdJW2osAD8XB1CHDuGQO/WXhNwcNzkzmDrHVB9Xo
idtKGktNWuEQbYCs18gGMQVZAwduUprs+FIbdRj27LC4TOcg24Vu1yYGTfDWE3hjefoW0PUXu7JF
Tp1cNIncqdGU1oxwZOoNxDWk1hgEbAjlp5YdKRKayNDQ252km8Q+MQgCUfo2H/dpKDDTLGUaZCer
qQFskS6dx6IykFGP+kuR9M5EBXnnVz6qEZTRCpbAwr6G8bckC/Gu0TIrTcvV6P5o08ZRHfchlkAx
FM7l2n8eDymQy+PP0tv//qUiiTYQ4ePyFoYifJerVzJVycSBIMJeH3HF+NAYehD4NsXu637OJXFn
VLdFiVEv1wUMexXmB1bfTk2ZfQMWNQQ9LjwSEN9n4WJnczc32KNZ1jWcsH0jWXRzpqRAM3oTQx1h
SxSuL790GbDEdkRa1dQl7UknFRJ0yK3zrZa9mXLBngPZvkEFo+WN+mkp7uTvRHFHoQJiOFWZXCzN
VRj4Ezb8WwC6pqqlK3Hn2E1Fwf/9iZrmVKjashrxIK5/FCRbqL3GVNw3Hm1i2mG+4uRo5x10+Z45
c1MX3AU+ejw2nfGaSEtC/McaxvA3IeQR0hzqY0UUpy6yHprTLIKB9i1+hJcx+IDaazQvvFzGGagp
M8/I89noDZCQ9/qcR4juH3JZIBpQT4PZFmm8uupuu8tKWEa5sZALmdN6Rc+QhDfdOh0Mn7kDaxs5
Bv48cxvF6N+pzVBZ9tZNRJjO4i2pQF5SqZ8J1NvCU+sIPIowvKSkyXckn1z7m6HojUOt1pNDQBxK
1GAl5LRYqX56HZT8UEZaNkiqdtU14qAYe6AGmZCJ8obI4MAoyzVhUVsrGZk4kr0tdRgZJHLoth4i
b8vGVo5OPgSaCjWpvNFdGj3j3w9FuGx46bTRzPXfTR+DSNlWH0w0b56uAjtE+PfnojRrxio43Hxs
40HIyMZq3uptnPvAEIHR4tuYXpo009GEY1eo3n8CCNgxj+YdsP2y+6zTjL4TK9MQAlvKfu4/fAw/
74BmD7C4sgm5QBLvQKVPAS6ItSl1A07cD+CFPU3AYLgyONX3hblFRgbZU3mMCeojQCLKN6YyrZfA
d1x5QMwZBVWRtF5N0DtIwcssz+Vwf+jT65fsc8xb6KJ7OyUcD0hBIB1C9go2CPNOCpu4aK5NbjiO
f6dHgmkucUVpZF6P8fkdMmVBgkGYbkL6PFonqJT41Fs2o/jagPONCzaubIiWLrMx1bxjNRPD9p5I
FdRkLn291RejySvnFgqBIk6LFCdt7NvHNgsr/AwSXyuY0zWkNhUBCi8iaYfvdmPGAhvQJeRdrrr4
Si1ulnuoUesl2hlrF/vI3Ili4gv5Zmc8FC4Dz/SaKy4u/15sxccakjaPgIQVYyJmIMi4gJrVFSuL
/TuMUIChbMyljrir36GYjAYJaWCz0X5+p6LYkxLNuhUZb3aYqOcFTC0+O80+lxh1Kt+bZO7BlBmP
PcWLlstFL/8Pb/q+c2HlhOoH//0hqNeILQU46cuAkJexCU3B+lFgrlCc1icSlSxkyZ8RCVP40wnl
+OsT3Lex/C6Z4AsYHrcr4/RLDl84JnMjWrwTqaHME//X4VY0hxHJTP1g8ZXfSC9/fxeaKCSihjYU
PEqF0PM8zZXm5w4v59UyadcnnWVP7eu+vnOYSNypl2dx/wAiWdBUoPQWxSGEE3Jkm4nrMTkhDJDu
O/ApXeoNJiZJMevm9TC4/ZbxhDvu9HfZZXWrjLfnMonEZGrTj5T8YUUHZ4dQqvPsblIgDfchOL+Y
5y9vKutLu5QlwVfTTXhkvUZYBGs3ZHky+KYlmjRAeYyEY0S7ngds4qXaANw4dP1UyMbEfT12NVHS
6fzQiL/F5V/16bCjxRzyczuDOB9FbOogEC9VSoMbGSb7VZraY4rR0PgfDZ4A3S2gKbqVgwvv1I0N
DZL0emHHe0OmpKmMBtwJa0g2+aFwdQ+bb4FBcwG6sxH5kRruiJVktxtbPER0ktMIZrg9VBQ36t7q
fkKwHgZN7fJVLSse9+HTKvtZf5Y4+kpAgnE7W7ztGFyYzk3UbM1BDLNNPyfZxyo7mRtaNbpbNzZ8
ErXbfl2aFbDH2TVYeTiluYAgCyZtC58hEvUDBPbc32PXQR5nhfEiZyYW+KTWzT5pf6qJ/WjtPUtv
lZtCR/5BEXX7LahlVx/1yE+HwlWw5qfD2+p2g2aV1cd1lmXelWo+ZP3/s9ES51qNieJag2lcwIJj
0K+GZeDlhZV18B5JHEBQb2b/vcvUN1uEPfBjColLt71Ot1vnhP6ugSBbJOS5QsiIWY0AK9KM3mBx
7KAXaZcMIYOLj41Gpv6/i2YJKKdFL4TIEmm+OiMXZNnk7nN8Gs2FzDE/2nzuiKwAEBkTeOCPqYH0
Jpinh6QcBRIuUauEfPhPbv8h3qAKgcqNeyMCwgcA7TakpzLmF5flNi8kpEyOi2sl+9j5gU/wYXKk
A2VqTdH2tP7aBsbqoBquBN0M8FcjsKzdE7/ILz1CN+y637QptTFoC+LwXlxEuLPPmMq8YweNTnzB
MG1bZtahaJilwvmQmYZnWDKAGUNZqO+7HuX1eP3S+PrY2nLJDtROf6PmR3SXIJAal5rrJUR5SPdr
4wLDvGhjtWEZ5w9rF1RMCEBcdcsBUl0x1fwYEWYmD5GK/R/VyeT64FArbRI/sL35NvyB9lWCSmYK
uPDGZTrT/En0HBhJ7ewDbr/bPjFCt++JZNRDtNKBfs/nYJK4z8qVQ5ndTzwwDz6VXCPrT0fQ+cKu
PC3gC4moCaJVA6hSMa1bLWE6q3pkCeRanEKmk5Bh8P/DXDlBxQpP7ot2/bLAsLPx3TeEp7loZQR5
Ch978wqZl3ChSwKzVzNK+/m1Br1tjY6UHLv25rQU2eMPcWZCfF2+Eef46Jh7iWyQisD9Yx33L6tf
W025kTgzPsdbYBayoVSST8d/Rsu6ckFTKQDLbL6XL243Cq7B8qS6hyIc2N1xAe4YFDoOO2EC5Xax
lKQ6XCTCx62apvs8JDCRPCthTQlP3zpuitZhtAGimHyebw2czwV92gT56LwOrQjmdE9ReeYyLvL+
3uG/YuWEf4OG5Dh0cHgqelAvZsGzSYNpPFxqMh7GsFQy2D9mA1oZiKo6TOp/H6YF+ibi3XNWlV9k
hxCRk7G0y8heckdb7kHJoJP9pnE5yZQ76BFkmQSmnxwgOKdcaZDopKpU22svzVIR94ToMZUZOpKx
BZF6gTUkoEWy0D3N51+iPSLZayYdZdcMlu/E79bIZVXqDggtZkj6UDsqcpBUoGcWk+Y9+BJHNG5+
AWfzws8WoxCAhvnxHWM3je2mlRcsTjN7YHEmJGXAJDF2f20z9xTKHRpqtDngd+hud9B1lv8Svd1e
0MYuUWfdkV1sbCeg/hPaJV+Niw43qrebZHnpXMXS/JfyuhedyBlXxQzQFo5yWHwdwi6YCzA+SPpV
kTJnQM0kjC/79m86zrKFeh5cfJRYL1xKrE6MgKRXJv4SkhLrG/4+9lmhgNslTRQlDEGLOIyNlq1p
r22LmJR0OYY2B0w6X2b7laYcRNJf0ZsW2JvZQ5y0SPVoZ25MESbarerPj00/rRQRLMSFOFZ1L6eg
miw+UH0X+tjxPKKIppE30zj1CCuEExildpQmkmNndHJxaMIbqnxjuSDVCWdFABmRVhkhsK8wO4YM
42V655EhGOCBIZvR5kqqDUtcfHuDiaetLMerddnArLWZJuQkFFQ8T4AEqsOOkvgnCfKrQOArsffu
EEjxIm92KAcSGMShg2Oq/QWu6lydql4HneqZLuFcJF0l+qNRAvV+yTDoDZXfEYjZhTfnzrMk7/Gx
Csfw1OUJpXc8XwU38GIUr+VdxE3NPTEmTLOqpgKb8vz1Yzg1kTdcsg+iJQax+yDHSeDILUV58l5T
4V4+fEY8zxQPHm2CfqmNGvulW8PtkFZvLJJZH5mTU5odl0Hi3829cGZqwdKKrATY9E4Q88+3fnj5
aWU+4HdEWp8+QxNZ/aVQ1AiQWzQAycjCWhDwv4oefFgyopyO+oCeiB0WX0K1VY/+MDYpouPgzX1r
WvYgi96ykV51x9SGMWGMa96G7rrpdXwTfXwIytDCEfaqrCDCBVaFvbmYN8mAxdsXj1dgKPGeibIr
n/Iv8G5junFmA4F3HEOc+yuevv4fM2Qwhs41jnAziSAuGGk376mQBbsZqTgULRjmgzFaQ6ujX0Iy
HL4qrWNR01DFoq54/oo1wAVEB8PqHQq4l+6aZKp8DwX6cLaRRlSBRhJtNeYGLBsSAHtDNa2lZg1x
2LfAmPyDwBmXmgjoSPVp6F1ZkWiq1ZMN7zQRE5jf1ej6Omw+ruZ0V02uUnISDxIeDKWC8Gp7JeMt
IUuwJMcyj+FtClG7b1psa5hI4z7bGmerUG8FfJp9eoBGbzY1QX9XK46sXuwAw16N9EP5fcLoujLj
gnwabh35Ao64tpfhcOkSuRkAqemaVcht0zFN0DQHTrIX2GCtJ/d24i5HTA8o1CqrIpUWBSEJDR4t
gBUMlKPeWMMx3aTiSQv5Y1U09Oynxwapeo97eLkaDZq1f8Gim20k/V9KUzhtrXnwBzJnOe8vz3HD
/FgndKhVEnwNzJuk1kZi3XUbV1fMS1jPTkhfxbR9uaeV8WNIpACu7w5XEKofrCBHfcRXS70rGkiv
hV6hsONbbibiRQebYsQPWoA0HcXe+BWfKsjlGIonBdU2i1oNj2MwTA0rF2pnT9pmEZDzxJRER/b4
LbUnC90DTwW7dVegbVipaA6xGTzPyBmqhW2Nax/gWFagbmYibD92WqQW1YhO6axmlpw7LWw4+3KD
jPJO3e0O84P4cJlhpj1pd6+39cB4jmgtrAznWyVE3dsKdGH8B3M/jY647cpZmQyIqV4wPSvDztBo
sa5l60bmae5bICV0kKWUNJFa5w2yqJ169PvM6/LPpu17pjZdAAgxQpM8XWyKTJ5OK91M0dLfde6p
Xx64zhVn8tFnxNiPgKEj+pgAQh8HhuDyVsikf0SHupDwlMAHZZgvfQzxx50m7ytTB0e5hBaz8aDy
3f9aZOHVAGX8qeApuzLnfXCc9lP8qavPiV2s0QPsLmKW386/Fg2GNFrB5FA+YBMZLR6L+MxC3jMJ
3aOs3cG/INrgKsC2inximsehDUVWqraZMcRNA/5X0P/XH2N5G7tnpuNn8/Jhss8fLSQ4ImHMtIvl
YDZ4TCxGY9aL47RvFPy5pzQAR4QPbAP9Gmvm4JzKRB1ygbwxhOPCTwzmLlNc1m7aS6nf3+TE1hUi
PH47fY7cBgfiQTCBA4H7BThILTIE7uR5Z3OI8XLhlq4oUb7EgNXZl3T/WsVaKF72e8UAX6mQPoQC
4SeUTUc6G/FSKz7otgN8DuLho8LjyTKvnEc7A8sFML0pcljkspkE5y2OHRaNITk83EDdPztj1zn1
ilbQrYjyMpeAs4ZJFVeYRtJNitaFGwQd0m605v5pzDzoWRqiJO6NClkWQ2pyi2JaQhm0nwARoMnB
0HjwkPSZxGsv/90oYvHgLIZ7AUQdRYSxTBBmcjpCny6SqUzy83WcIuZ2pH/WSIItmMF1tEbjqXHv
O1BEwxiZlbrj+/Ro549WpffjAzLMkBe5/A9QFzbU68aGLJ+yucQrkzhnkn2QNBEEynXjj7dmXzV/
00ZRvxuDjjGkSuVYmAuYYzi4FIdmIJA+6+jPHwwgjt7uwRMeEExu/8ZO4p4OJvmVrYViTTJlohIk
r4W0bS2wmUs9XejDx+DxGQ0SSBSkC0lxdKESsO+HqzTc8mkjPmGFZo8rCQq6lzgaSlErCp7R6948
P1t+OIZHHCAmFRkuHs+Jf8uorFwPHzrOdIgnlkyC6MF9VvipN+aOzqMAkYs3uEuBzAycwwwbSKYn
Oi3SBT8MwMoNVIGD0oN4EryP5oQD3nmvo9+Zyk8M7GyI4fixr/47TVmj/LqGvnk3d8XtFYKBvkFw
yUOePe0+To3X4Jqa04g3jTF8RuxdUoYPPV8Ydo1N0xjZE6cHeO+oSSnMoCWfv7IHlHmL7BDPuyna
Ohmg5vGXVcH7IxkR0YzP1kqYKLeZW13Iq+/pp1esbvulYFMMDJfemoS23/zF9KOC0tB2BYALlS7D
UKpQjNE/L++wRYUcG8EXhhnIvn4TnQAQoFb8+k/Ca1ZG/VruZSgiO7yt3CzyKZhknbBY+/miaeu5
cyLLUpn0qfcwZMdQQ5z8mbuZhlE2XpN5W/i/9TxjBheKIQZ+49A0bPMn/3S0SOqvaqtq3A7w/NJu
LGCKXmdHaQ3bntKVwUotItm10hd5kmF47qEM4BBw8tI5reVHEOvM/jnMfeQHy9RozqY3HX1rAYu7
dbziUnzICBX9mntpTCQf9H6IXSzrruVGzWucZL0JYvijf1fjABsH8lM/eYTttl3QmgJ0lFAGoXf6
NlgCo3nEh/Jam9yY6rqggyQy/mNwU7LHC8IbSCnh/UHRTBhCyjs3lkyh8upFu3Uwi2PjjbCBHQ3O
lsCc7wsZCn/cgJ0JOEoy1q0A52jZErwYvSEUi8pvo1Mz5BjsvYYX4mSYMXLhSBt5ZpW5cE3HVPNw
K40Ee7a2v1bHLxmwMjX8CLZgUI0xoq6wIKpuZ/P953hfohNhTIEd/M0Fb7WYCn3tvDRBKI1Wj4sq
sPAkVy5iDpbWbkxJR4TM9mw1IoVmdPIvtOVKqUsjAol4gl3ECayG7IvWM4gJNkn3wUuv4Bl27EPv
u3wq32KqUucvrGYRJ2a60iMYWnGT3Jl7rVacJhxxElAMHjQHZebZNwpiumOmjA+msNnzqwlRVTZY
VCT7DDm3Vl4Pr5YrWv6d0eEEseLQ6+aohhEv/e0J7WW4+0nXYjdAr6xFFU0g9iOho65nvQwmnRBr
cWizeYA3xOYI2AHBI4qffA3BEVqd+rPZecDrGm4Dx7ev6D++eh6FWCA/qS3QxMg9SYZ0O0OYymiT
X77tO7jaT13SMSFJ+BK7GpXWOtqKXcUp6ZE/stP41XldAbj06Vk9M+OYgeIoDpbDFoubNAYUsfSH
Xc0HPTdoFsAxsBQ+bekTzV5n8UG2UahYcWSu0cD3Q/mh9h3m8uZrrGqkft5HIzrDFhaPxiYUcCId
MwuDZ16G1L8blxRcvFnyg0a5X4xjtp6h7pPU5sIAmbbOt5bI0VMu73Dq7Aa0z+PPJ8VbfO6WjqaQ
TdnRKWUzC5OmbMuES3GSpjfDLW72MiNn6WWuD304G7cXPmOrKCWnhZ7dIWLZv0XMw4n2rSDzBY0I
aIgp4SeIix93ket6gnWG0pDMTJGN8BlmXQ/LZjEdcLmLNCR/aZESoeraelqQE2df45kDR4xcgkQ4
HO69rgaS13lUGWxyQpVrBwTqCS1AE0+xZY55CywjzDsQiXHqvmH2o6+O9OkkIsJ/fqnSszxamh/L
VAfp9Do+BYioQU+G58gmELJw0ZUkeZht4g/qhJAhj7cN+gkRTws4TzqGW1oQZHM8A1Ql/qFOti7i
o0ZOcuJRo//9VeoTnE+LAYdBbryjRbcJHJklYvZfo9iUJ6nN1mqy3QOqkOyX+Bexn4FHIC7iz9yG
ro+ltJAsY6n7ydKfM2BEK1u2R4mCdCnOhVuNxtlcmsKab4HM3K6ylm5L6wk0Ud2AZLv0kgEtyul8
J/EZLtpM+2/Xu8W0R1KajdbtH9fldtLKtQtcNxMzrlWNaq8LMT4L/C+oGyJadaD2X6bm43IJuopp
CR+NU5JhGlJ0cvIVU68OBwb+7/Yt3qBJwPAH6jl3IJTH/CEw6xal5VvQHOUyLHSgOmVkpr2yj9+F
IKsD2b9Mry/p0GWzu1S8FOGdvSxaOD+TUuMYeTvR2uGJR95NSOPnOaOTJtIA9LA0+jJpSlf57BxY
w2grUQwrDqvbfH1CHK9OT9PfKLETqWHkiiPSmBiSCdAWtQgWLkM+ikI7FpbaaHygD3OL2UWZvmI4
1wpNkqImlaXBuxa0m5bnt6JVEF5DoutMRAzaMEb8lL06v5L626dLqVZ0by66FOy5MEUFe3EGEpuH
5/A4a/I4pjEX+vFWySVitXIXcw5SGpw/hXPj55fQbuvTx+gCyMDd+7WPYQ+85we1jBNMDndsQkoY
flZ9rHLJnITKBh/wH4QCx3H0BTjdJ0BJgBcr/edQnfR+04FqcDK2Oo3fc2O4MT1SKNOzpUvz/9Dq
ZvzU8G2P6uL5itM0lnP0HUprkcNQwnipNqfJk/W8t4BYfCNc1urTc3mpVa3DTyHhf5YQB6T5G84R
/OHEoL0u23ii0+GyTj/rYqHOM0wyiYMggoa3hTDYs1KlFrlzuQzFy4aOdLDbi2n3l2YKMOvJ3Gq6
Iies7lQ9XnjPGVH6Y8hzHThlanOU5GZhnZ6DWsA2MlGTv8u4rObdCl685zWU/uk8+DoJ4He5X7ID
pRGxSRLBR5eK40wvAAOkMaCvn6g6s5TjiDP3eM3X1OwLm6SVjMlAIKSLrrSLWgiJ3SOpog8ObJH5
dvLmVLNGjUITiS2L7ovppPuEfAM7kOHlby0w4IWIRlgDEjIG9Y7F5opxJ/XyLiHun0xUtVQBb07Q
yGVbA9hh5hbaFUKwy2SNcMEQuRFNVVfbU4upp5QZsRt5RrmmNUEeyhMK2IOQqGztpn16trlSBTWZ
UyCHaIU2BhEOC//iBgZ/6OSEQ0mEgH8dzjZVaHsoOY1yQ5/T8WRslu6g7VcsybV2Ckpi1v1KghRp
GcKCqJyL+qaEVy8k+VXFnc4oSPLxraLGErUOliAeqE4Xrwodf0kxRPxGukHp/XEZDDB2lvliMK7X
smW92+GD3s1GGwUBIDVAh7Ldd6G3wWqky8eU54N6pyF4NQHs6nSm9pqX9FAbyb2f7VJNBnNLpfx9
U6kO6wuC6YrjyV9mxMRM7bOQyq+lqqOAvmQnKXqEDDRwSCdesD5EtaaLzqXYxNJFZss2kMGCo3kl
fyM5TjMYQyRs917AIrBEHLKKpKJpBGOnidr1iH33NLeIGtIX7W+Y2Bu2DsN5N/0aP1DjtjxzVnzT
ur6BGZ1VqNqTdWsUCZO0R6ItQvJUM3K+JenuOElEFqQHERNlhALDzitUqRmzdhhIq4k4hQZNBFQ/
T8IFVNiv9fBkItoZN26ZycTcoOLHnim1BmTUAjc8gApnlZL7cWTA53xgFRXvhe+Eeo3a7w1yGSDr
vx5d3TL1xkeDOvBKL97CeQTDrlqmT8wdlKoriz65pdo7bphjk9lGwxx/xCmCDE+C2sRlSXzvIrbv
P7ZJZmzVBI+XhTNuyCf+oqWRW1BQuICHStz2OxhtVx9S0hs6AqBBIJanJQ1UybRT9Snb5NY8susP
Dw4ge4ioqRGJ1OCcyHR2Okej2fv3wqGJpuEF1o/B9RDzA6HfCbUbsv9H5xv8OdHzMHOgHEMp9CHR
CtcGVFUF/Z99+4jIrYqGKJ6HIUSMwEL8/tas0acOhdji70CF7NAbDv7Y2itJgZVFFeSX6lKfP7pv
r+0Em62gX2cT94iaOQp2LH9Lph/05WVh9R30fWzy4ffqblMDPTMvY6Ie23XK79+RJQeBHrdjanx3
evDqVjGDBo+wMxpXYyYQAewpnA9YdS7XQZot+pAnFSD0te36z3+W++v53RBFgjUVlowF9tdljjzY
aRo11xfUeg7k7WZlO4Ysgy5uDlh4KhqfWU0fAOH7+3kHjg9SysYJDZxPwyvmHBTxbJ3yX+jNxn02
5x5sul00bCBpPFqqO/TSyt3W+o3X2cHLOhGpVfGG5uHTplIRh85EeaMaOqEwOgIxfyk5R3yHC2Ov
GiObkUNgs4gszOT9t4dtEGP+8vMbjICv0sSCbwvfHSsBAaS8gojUM9nXwkIlB/5k45Q0hM0Tsgk9
P9kVrZ9uspDKsiSCxUILvw5BOInyO3T1f0IHFg9uoicrwGwrEmHYfMl+CS2g0m0RxVn7OFPkqmcl
nu2NslNU1gdH1PCXZcRefyQlFxKmYQipx/IeHbJmH+8f5o9MUyznWgbUuyDaly5liOgIpsla8msb
PJehymKgDdFhlRn7BiLudIyjSI1CM2c5U4m8ATia7EWKYZ0p5BppXd+X9oyeBdhGtNLeR9HFmF4h
8nSCna2JIoIz5swYCJM9dsh3tUf0g3qZ+XjlCs7cpXzKVRO/WLmH0e7a32y4sE+hmUAZDb698OAO
l+TG5t9lbXpetOj6ZqKpP/rg68/FPtIf1mqskK0w44ClHLeVjo6jlchQ0gNzi83xCTOI3MnSvdgf
NiEdnKZNuFy+yC/k9kOaJPLTWhUGfnw/0KMXdoSIQeCqSFHUNGwAqBsbYxUNQTDexJCI93fgWlcf
nRWNRquGkKus8mLMUy5d+6MXFUDNNH7sAJXuCQQod+yXflbhucgvwGbGCIgdwj/Xu/P09/MAIMxb
GDvJYFET2rSTh+h3MV+16Y4FCbL0Zax0dIYO+ouWj3NFMISdZUFxKX+09b3jBm9LHcL1gDU+/PQ3
YWUbL/EIxdbpar9fHEiG7/NQdPX4yxaTLpxEZxQelWAB/sgeEPZBT0tRexx8a0YEgB8k12DViZy3
Cut1FL66zzxoNRvAmlU2ZvGuQbEmoCCOrLqBSmHryUUbHvW2x6YeeBbMvK22pIy06+iWdaBNZWu3
gpSDPx4QJJWF+Rjj98SQeS2CxdKLFRGP3jsQtoeOVxBFiSXajAzimb8JWST/eD6WSTxIIDpl+kVM
bZO76HozHsjzPel4ccRd8tH1SySQk2ENbcUwBe8e9xSWIIAetB1l6vy4fuUw/xKYhC7oeeaXuBwC
+Qu5+gy6z5tMXOZFNF1y8sdMSJyZBEXreFe15Lrn2EUt/YgV+oIXGa3FcYe9PGT4pCr4Bt08AJKP
12crE7RI24RPDMr3yF4J/cKFXtb1l94MlapK4CS9Dojk2MlanZj2zK27hqALKqXNoZmVRH3B8IF9
Q0f1kF4q33R/SzpxJK+Vbc6d6p+ctFn+QE4p09Y46fXeeOtOKSIYfmXiY+seXqdsBcdq3i4TASnj
IrlduN8rJSjuUqGJhYjCn3gdB7rVIe6Ps7XkXoVzu7aDumKrDi7v8CJKXlIM8yXJVuQZXEW9miwC
5wJh+3BImYny0ObwOoscSYziTk8MLVeKG2wa+GTlS5048jcNz/qGZJe/zRtyyZj9Z2YQE9vOR6k3
7ITTDkP+SqSW7FJq8BH00q17PgOs62KZ+SdGTI9OE3+jMUtimORhtXV9JmBZjC+quR53gyjbQjL2
bhlcK+mTE/2g0VYxFItNfhQsRUeMGHrMmmONL4Glmgy2vKEPn0seg+0iG2oiM3gYnT/LCOHEwHSQ
KkA8ptgjUUduTsQlwFoClzEImAfbJ6hufo5V0cAuuZ2YKLPUDsSEjB5UHOqlrfhNUhzogCCaCoM9
Rtx7KHUEUeTcS/SXCB1egsKUpTfKrRxL4qS0kYHJBBxSOrVg/VSj8SS75dgbkviIPvdrm9ig7HsJ
Hi0o3TidvshZ1PMKwSLJhTwhsjIYXBWjElZCZLOE+WJBoKS/juK6geCbo/JEesrPf8XxmGKEfEez
slY3uKI+CmeoI68mxEAV9L8H0qRvsJuwAr58c8hLYdpo2H6xTcCA1XDked3KGI4ROTxWvtavEvsi
BcpKJ/R/6Ve1TKdzlt74u3kKRkQi0+w026v7P9QxASvGO9vCSlV05O6YyATlCsJ3qXXgYdFqNbsX
fwEeVK7PSg4iVsj5QjbXLtr/eBytmJHz6rVjeo+nJkCZKcMBVEv/AgjyhY+ZU9faz/fACn9YLczF
moWMN54pJs8Us1rwERNK3+69FEUq9/M105do0T5b4vS06ckzo6b3vhKbRPgqxjT6NDe0O8KlKza5
KlJ5L+6BFBFcEv/V67e8iNtzWrX0lxIEmU+21768+GlRe18hFtRcisjd/isb/BJ84yR95Hd2UYom
XFqooXJPZn8T9o6WIsSg7el70ZsJGJCjGALQkyXuCQLmR4VTA81GWl+z5wUi9ixQqLMiDk/M8Dbf
Cr1cS5KYD242RjKs3dKn+fKzdPyoApKICybMmeRi2JP0Zf/Ye609qwGpr93iGTApjm9lHyfaJ3oX
jmo0OR2vz884ZXsqYXU4NYjBPpNlvoSzLjn8UmS0FCglgl9ugBk8KwwLTxjVJcl/CL4E49E/qePL
L0quMaee6LAs0YY6/yL7V5s/TMwmdZj+/1nVlxc4bAuhlSvQArm4N0KjgVyEvBZzgUPFWnZRmjRL
akinsvy7bcW4yZdslIPCBbuICaEedsVpVC6fRxy8QhWyoxrA5UL2yKbkeEe1A/ciguCEoFZooHw1
LdMqyTqpZpxI7ylGgwAueHXwbSg1OxwYSD3zTz6vKvklbBBjw/N65PZqL0EA+X14ZkTRkxTm2LGr
/+4A+vkwJ+jaX9Fmsrewf6iuMahRn1xOWTE4S2iLIjmxV7cCglqAlKxb17V050E+PRPpIooDYKmy
RtoTg5x3GxqSeK6+JiO50X2LXahYAYm8BepCfcnXprjbYbOlvUQduG6+AgiVWEc0D5Kxo2OOVSpy
4MysoV1KFtBVN4yEd8ljuALEF8l+Y/Hr3gDEieQGYxYNGi2qQ001c2ziTVnrgfAThN0A3TIZ9xdr
ApFWra78K4rFVg54clj3v8TBlXfMRsA+xgFzgeqG2fAFBrsQX4e0BsLpYIkQN0EysiDXP2BTOA+y
olhQ7gtewYSnJuQdZlRUekPEwcNZ/awG/+gsc5Vtt0Ljg0vayCct012QM/llyJOXVxUA4C2WrgOS
uCEjY+yHRELihpQAaE9AQpk4jcFj9YlHx9UCS5rKrjG1AhStVUELCRt+boZh1MQmEgXad6djn+sa
jgaJOU7+6fux3/C5GDLxiPMWAuu9gtXR5zcrM5ASPJEJCzSW9OzzG4eBot317k/whdIR5kAQ3Qr5
oCdWWXUOa+SaCn1KUZR7S384AlnrskOKyIrTBhuGTlfhcV6ubeFPLY64zTb4ThQT0Pq3asrXJkno
rD2gOXLHeshR3nAYHmKKe7XUwaCPG1DunfrGvQBxw8VjtYMs9X1jwgoxyShCicn9vAdPMtJrjtyy
MkzFGcwWgto2uOhKq3HLgzuCqChoPhhfVpR1xyLuCes5IZsw8nkPndyMqvGkGbuoSzc0hP5E4mD5
QMhAFMYkd/cfb0IKFli8pPRwRR8+ZTdLy+TfBIDMdtyEIjmE4PyC1Y+1Ouo2sIrmlBS8hWOaGJUE
pjuFxjeou8rbCvOOo6i9M8FikMv76pF+pIx4I1OcdZo+K59Z6FFI2OgYHWjQLAbQQ/7AHCSyHEHl
e1Q0D2/UEZCkp46wAcVP6YJ7ysFh6ORFkQHCcSxLWPBHkAImeXFreZC1Un6h8pMxkrsXwLQ7xGSE
D0uWK6+U3FZ0v6W5meXzDXADZ8QE2+JaOpyxIkB9hp76OMahLLFdbv/Xl2v8Yalco69sZvEoQi9k
YMIBd7AZS8MQd1hKdsKNOLW3qP7fzOCHnRA/pOiOVgSMsC95YTHQ2E7/luiYCtnECpOMV3Ak3YqI
XdAYV3lb4YLbP5kIMBAEWICKjq6iL7CYsKAKuSimg6TwPH/6V36pQx4opAbT5aj89heQ/Hxyldk/
oh0vV94S2ffrPuWTYDAI5H63z7CVI9wPaIzr02hoImRLCZSq/CbNuCh4sxevjXacMJ3FiEWv9PbC
Ml724ZO1KxcqyOCBflh7hcBbGPBXMvz361EupOvvrwxjN3tlYj5EYEIH3MobmZXjW2amo4fDz4Qu
Wd9XQ4ys5SkrPqBojtMnjdt5bgTVVYsCnOvP5nBq2ewin7FmwnQB0XIsnjvk68/zLt1Q5EEuUoiA
vP09GL6f+TH/jS454/7GLbTMLMkThMGhYb3g6fUFTVfRPpKh2tIvNEaZNdu3JM0eglZux8Mr72bE
qOEbC9fszrRD4kWOrAMMuCXhOEgXYj8yC2WBw/2cLFNu790x34Bj+0d7XySRR79LdMWDGrcpHRCu
rhOkGA+0uPUzRuIZrfW8nz6iGybeYMiCsiUFX8VFjRoxw9+GHF7Zuilron8DCpBF/wG60IbRJEEb
eywLQC54+BRogMbJfQZYYrxULmyxJuTFWLwHuNnXkORCcbn19UHvBjmRQALomwCayeT+lcBWnS8r
qWbyrPfZ+sXkDjq438u2AmF5rDFV0flkr32yxSAlRrpSkajvL0Cbx965kXg/BfqY6BSzGzq08UVE
VHtELVW6Is+ZEOcfj1bt8ePnRmRjjbO7viLILqfI2eth+pwlHuwpmQCaJfy7GeRlWxiduYEuAWzO
5bhgbSb+aaCNYIEiW0aOPU0JGP9fItjjhch0o70O0wU46GjI35/jyoxi1Go5m7aMdAGSo2/h7kWB
QZa7Al5PBjRGA8ntZZMRklthC6kl/RSNt6W+7Ddp59R+jIq1uI16ciA5Gc7lAwdWdWCOGKcpRBT8
kJ1dXOfvbE5vU/EJacgV+vFSvqzX1QyB93HwQErefFeq0u+iooyxAPnAnt4svTqK2NGusR3B+MN+
Dh/u11epVyxuaNFSDthhvn1xEiQ3dUOxCsHFuu1G/LTVSh2FQ+3GUkPSFQnRfWSIqDDTiJ7MnHqW
qRq1IhfrCfl+0cG+e7/i/Q9Umg+r5uh9Gytk4QOfxHT/RQKktD9NcoQmvKpo5/2OHx9b27SCOCb9
QKmLXRy3LYGeVX0fv3Wg0jKr6x2HmNMqNegxRSU6O1DCNELc1TWrfK8ud0aWQVaFNnsqkni9iADi
MKg2942BWzmTXfmBa+yuaEe4oYITehdykLNTPTc3hhtUVqWlrB5SwkMOZfaR3GkrHc1BupOQ/loR
mWGYQYM1C/GpXhr8RYSyT9f/wjKEUqZdU6LYQJNxg3dg+eHJQ0/0uYeB3qvSSsWp/kmDXsYtzfj8
RekpZORRzZlQBaIk061dku0LMJM93frOclvN2akn9jVaqLlWXETEFoUhGRoMWmxYYkgtyteteJyA
QcU8wS9FklFagqzxLI7n733I/mdb0Zd5781KCmu2NX769y6q9hNkUh1tNBeByw7Vh93++AyYy5eN
r/ExzaHJgX6IxuA7subpqII43VkqSxUDUmcbFK94VVcLgOSdx4DkQq0GxE0yRkjTLMGCnswl7nRe
hMFsWPZFOijwCYeq90uAemWcd6y9sxbu8tMw/vayyCJyQ1oS9Ud4VBPxw+bhkKLv8AcUJoHqbWZD
fTG8gAtYwOmG9Swlt3qMVq3jvCLPVuL4AElkTvGO5s9ZElXGrvHaUPvhhx0hIrbzoS2r5Li3doRo
aTUTcXrUZk3QCJDnOKgljHc2+5HN2EEJz2qqW0xU/hrfb9rtc6nK9KifYxbyjpFPxVjj13sCtsLW
qEY0ASYAkRLZZkBFNR8Xml4fp34IqsGMlavuAJibObeMD6LzUQlzUkYbZP1BrmWEroGEkC2Ff45w
aodgbDdg/N7rB2B2KhfIUVsSenc75kGDYcozKkmNbkz/xusFVV6bXZS+pFaHfHgoIJSEFHxUv631
PxvskpafGB9GZ9bLQtWaB8puCfjM8Smy17dPF1qHwcqbqrOlM0yajBOctekNUg3cEIm/RZUwAhHZ
G1PBLFAqSwhLcx8yR2ga//iIAtB+MPEabcOEkw0X6hr4NQt9/pHd+NGxtqeAKT7tcD1UfZsOB3W9
sWImjcwk+DZ8k+RCA51vnM9ta6zcnX6AKMTG5eUPcrHzLa1yOOFSl/ZZk/k7cs2ypSH+8XncpaC9
1OSi2AIF1vwYaQepKHNFK1DO05eOavdO2YX8ZpWSAhMiMVeNzUC45VnJUrSgpbluv/CJ7TblBGbq
sItFWlQLRFBgVISLa6NBxcc90bK5DMlPyrBpn/axmSDD/2lf1GstsjXebbkeH+r9//eP7avOz2AG
C8f+8HRcpRjoLOUAv8oQhYxVLQwPZpyaqov0td6FdBGWEFk5WTEdB+67fqdZku+RVGlwKFy/2omF
dQb2wAb2Osjh2hGURfBNB8dPEMxyMyPjludq0t2ycEhLuzshdsgeU4tyvpv1dCcwsVbWoDdmiTaJ
4XFZQkzS8s83OvPacsFtHzVD5RUXCcNnHf0t4SoA4WS6rcasLiOEjNx72TrhDImNoBuusd4Ule8G
945DBtEgNgspDtk5A5ADR9rpWjWDiDkB7RBnzc5Hv6ovD0xJPcizWINedfcdrgm7QmZL+dP4a9fu
UMVzc1Jd/godYF2Z9Gr37YvHvHNN6mbIe8h0kDEWRSP6dNuRMFD0TA2FYj71RNiyg37HQsTzPWR3
L/frab1hyTdfJcWDlRBi46+w9TC2D9/06xuxWaOI6jWN0LLSdthFUS3wALjxs5dZd6HOs8OmNMTP
6L9ETQd6nxp0/F9Hi9Keop3QpgMajgpG6PzEtsMbhaWoHhiIazS5BOMbAmEpP1hj5SmjTBsbxsAZ
0wn2hUBOf5Qc80KyqOTtv/Ogv0n3EKuFbZaA3K20csW7d6ynlCB63mCODccQAlerUAhteSxbfff6
u6CThCwg1aCQrYUD1wChzBwkCf9vbwZaAZXDKY3FID1UFRctos/EkVQgF8VFOtxZeP04jYaoHYIL
ubQ9Kz6Dvj1A3CYRJ8Doa3BP/ys2Tqiks5+b7s1PG2EISqLvmfaU1OcLAVaJHF07P/VoVrq39IQs
cmbggMhsZYJk4utBW3dY1UHWe38Pd7mGE/52i4DboukgwzkaknEY1wahrVDiDIlYHPxUkYPDqIhM
MaBDpem1E0SnHhjQthub8T7IMhum8epkfiaHz0/9S3OxhJvgTb9r/YPB2Avj2Xhl7RVVoPhlIsk8
KDVsLE3jWrOIk6HXpab2LBp4Stp7kSXVFdXTUysF0z+Wj9ejDDtOHudPrj9hdtTN78iTMIX/uhI0
JrRxXVcitDEjcJkTNY4dGQIp7eyJCcK+SnNIhlzK5JZa6bP/vibjFQa8/hHMnbgGhc9/LUL4I/UB
vozxcsV2dIDap4RMiT24f+ay3OfDKHWyPTxjwcW6UOFLeF7P68OLK6pgXOK6gFmRCMMQsn9niomi
azaLqvGWeEoh3rSF0pppwxOEWXwKK0YkNvX2GtfQHVILPjFqVm6+QJmDIQhgRzSMi1UPd3jL5vsf
+GqASkoghlzsN+T/GlYA41P+GsFDyfUFHTHCo3r1jXylOFrHFZvIZ5Hds4VmZZHH7qXi25MDzpWH
P/iI8UCIpN1pNO2NlQsgvouLOY8c0Vu8RyIh2S2Knf7mplr23E9geilwLShCKqQhWAdsBA6e5lGK
c3UoxObIzgqyVA0Z1VkK3txMBLJEy+fj8+0Y0mYe7hSljFOejY/cpvq9uFm8jWd2zqTuhhJCtyHH
i1PlYUeb1FAfxuehMG0ms8PWLoBh1Hwddr4sK5nxHy7BL/xfBwA3U6BYO33vUbXSHK0Lt6mx7Jaw
KpFSobh9wnSlS2zNpppiLSAia0xYrrwdieeVMQ7ksQ1J7bJo9ZYTQmovIWN+ig6fh94ugxeUJ+xp
iOBuK4JRHW941JaN4SDl6GqU5cwm8zqepTUitlwe+nUlV6gxkpsm2dUJy+dzZEoCuYyl0gS3obAj
OY6/ePkGSK1RvzpjJG2iS9hsn3ty/NmNOCUWn/DCZ3iK9Ger2HmK13YY+RhmJtpfP7Jw+UtxMQeK
xneVtY+V1KPrM0WrvAA6tQmzDDjSOFLcShYNoH7qIRDjPRCpEQD4lvxmXax8rP8+Dy5WGfsu0CYr
UnyAD5T1zYwFJFu7JCx8iW5CxKF+mZcMixKeJlYqsGs0ufaxoSr6SuIBAOrbp0V6cz5Hg84DdTCc
qGDfmD9oYn7K0vVjtMzsYV+So1YVxslkMO1sjZn+lHubg/g1GNYP7x8jr5mD1/oCFrb55Muy/75w
5S1NGZtGPQSVbyUBNi8jElZOwCYbS/Fyvpsca8jqRrRBkiTPItMtftNMjoAez2wAMLTnBPRILcsM
xDm55TCXQifm8JYTYRp8xqf3kixjiYPGyE7e4yMtWu5ijZZiB/017d6f58AxOvCzVJcR7Me1f7+B
MgfxTNMByqsrWDwScS4WXSAAVGu4gBNfQF2ojzzQ91a1FIbsK+LeuxgN4bbl4OFoE2SzzYZP3XUy
maTHgeGTi4qLSGSAAdPnWIedOjHVMqyM0uB5Tds34vUTTLDgoZW8YK4ry70BfxKdsI9aiDBcaDcv
Yw5+S7ZyAcSa/+MbWBhXyTUhTx7t4vlU8vS9Xa9iG63gluzmdAxAjBeswkB1GN9GnrnL9REXZ+6E
XuN4ML4v52EtzSJ4AMKXm/n2eEQL/Xz3NyKMT+5BO/EBbCAVLmnkT0g6Od1VgSbrJFXYr7TQN8Vt
HPabySH/h5NFNVMaDLyuHe1BiOkS567R7CbfS2CLkBiuTaDiV9ncw1XYmMDL1Pq2M68WVEFKgBzH
cT6dYbywP0/9D3TOTyK2HhOZw/HnmCfmPjZU3dL9632Ks2Yph8vNQQeWIMhK6+nwkhaxStD6K1CW
ic5IsdaRJgv0bDf53whoMHPwYrwQurQjbzYosvr+ZDM6tHeZ6ve0x+ufdElI/wjmArMqn4LSk26p
KF/Rt70R1bwjx3EevFyi9s/4CZskbQU/f26vvC4GQCi70Lf/EvC3qz3ROMzkctisV3ejFEALsCaC
FIteo4iL9GVXxZ5eaJzpFGumkbBWEr3+ARkv3UpMImjD81MP6Xg46A/6DYwfCK07Or+we7QUBGMz
NwMLh8CRmVuU3dLYELlJ45z5ZWcfVvYWHi7zK10MVTtc1DGyP16zPszAQEcZAU5wjtrSqJ5cqT+8
91xrgQAT5x1Y1cWrVjPfKs0XLOCJBKePjeTQaJDg7CsDwf5AeZsoL2wEpp2x+4whWgRuenCxoDI2
lLEPTR6RNVGERAF4TpoBlB/xG9cgyld0E/PukfYMwevPipizYyu6nvnoNOLNgbsaCtKDq+30i6FH
5BVmZ3tEnjM8kK2XHwmsM2S3eMPV95THzFMJKMUeiMZSXfMgDXCkx19xINqcngGZ1IbXoDSPuWDL
4aOVgzq1UrwzGVyB6k0yTaqY/gsoALS8UfWsXrZcezXzM6ISWZAxFeAySvzVB/1FXEcq1+JoaL8x
ACJaNqzaP2xSKzLSv4qOShpjq+P2PrfOmUcck65sIEpWlHssWCPUKwTY2VZ3p2QnGPLnv9ZzNntv
3ee4WyVTG9+pXe/ihDuzCutb55JrMoCRK5bv5wko8IxubykFaJvZWakExMiqxpN7Q8gLvyWTOBE6
iMA1FnoBbvtg5Ybv6LpM35NYsZEGSB0Piik/qRZhxBrB7Qarj9m+pDMhT/yGZZzWwT323D/E2bds
uyaZU2609LNH206t45mNgOFErSmURano1CZdw30GoxKCJ5xp3WYhbFKk4oeWTZeSYtnoJn5oXckv
Q6j/JR0zf1Z3/JZxTPWn7CFS6CGWqaHP3Hkume0txGYJ9miuMMyrd3DgqbTdqEGoWSGo08me9ell
8l38dsIS4e071Q1Fc8uyj9icf3KoUFsG02EruAQ7oqULsq1DXmM5Xew5c5AVSTErOs3igrCg+gh1
WT5VJeYfPNCxeZ4yo3vjh8YZaI11WnP+9nYdcqaa6nrg5TF4OFJGUwmuKE3ePhTxrjeJhPKR51dC
Tbg4XDMlYMntIzT0YPJl4u2bUNw6e9E+gy0hUvWVlG34Nl7k1dnzWV9mOefB6cJXr6VeVRaFF/Lq
HDF3/Hq+SnzBrU3Ewdb54MRF+QrAO0cnYwAwF2AE4ZM89UANjg6WEwxm/wGK06OiD46ke6dZRGpo
rxglW37iKraHGEtzdyyquw8gmbVeRTO8XbJPrwAnRb0D1gUhSG0Ij7E8AvPReq+mHH1STIgDBQkz
s36TYCcNXAdPQ+Dp6r4f4jWcZ66cPknvdm3/eNap7rc7So8mqPdkIS/HQQHbfqwaclOJWNjVRgBI
CwuXPY2RijvxyAE5TXIvHslwx/NpIKBLFHTjdBo+jtNHOOf6T1y94SBBwzih/cs2RP3tMxCOQevN
hV3wBYYTK3Yo6dqS/cwHOKiu8BFEE1C/IOuZ2QR+ku/7rR0H2qLSRZtYVxkLbs5UAZS1YlRPyooT
eRYK7O4t7FTk3cSSawp3pZ6yvsCZNGFDjWxhTQFxVMs0fMvlLrhMLhBdlAjHJ5mnw3K7zoSCU55Q
2y31nn7GIODiQyLix5wSyl662RecMdPCefnZYL5HeNM7g8P7k784/0s/k5+bkdK04LZDcT040baM
jsALCEvEQLpKzWiiC3CeCXAclcFR55419ZOBZwsBvMWzNnEnzOsGRG29pm8g6S2oat3+w0NoIl+S
iGVXpIAxxoUETDxOkNNNZxPFkT3sj9p8fa5XFGXWKkaXiM4KT+nkB0AW9+wAQCMwitMs2MYZUL2D
ejCUUHZXGA4dIvKvKnLqN+diz2SOIpcDA4BaJCPiNf3s64+Kqq5DiJXtO+WGQ0aYydH1mVX0GuLe
lEotQwwitMOUcsZ8skxN8jjYnIcxebVxX014LNZyWtKnDDclCLDCazMqlKYclma4fRsEyymV23cN
3mL18uh9772kYzWNIFppEiIE3OpWlDQzslRPKNc4fkd7+DZlAY8B6BZjGu/Uc8zl+dps9I3JQ7Lv
JPBTwT+HWHi5HSUoF1NiQSImsFaJ8hc3yXhO5WoLzwE+jr90QZmm2bXE+XHmvCdUvir+X8cMSYYO
JRnu+0NVdqW756JYN8fr+CwdO5llQIJnzBAj/IyyRa1rDQ4/Xlaias6lKVO3l7E7f89zr7MQ5jJI
oEqTtufebBhWkVDrwRzgc4FomEe34jzAn/bLqEeDcffDwxUBPJMQ2NO09t7p8kXWIvoS9+RCFdkw
mQDTfjOeGw3K7ZV4pyyjfs8fBYE28e3OMYnLH58Pwmku0I5exGfkPK7JfZ1Nu2xHsN2elnX9rAhl
4282X+T/PhQIIdMu2Egk843FoCfubufNBjocP393rJlto417Gv0n+N/Vwzc2f1ar9JiLQBSsMKQT
CPzIRYNTxjxa4WbChuq704wjvhlvTo5JLsaz0gljDGBUOOMYExzczaWSMGwmA3tUlJxsdDgHIMLD
VM3EA/KjU8TwKrlGiJrDG/Va9hEUc5Ud/wEWN1s+7R1OW4Ng7/tjiFWwKA4NOtk/xP4jRxp9R+kw
sSKdwhy4y1v4rUMbinMNKSgX2JJHFdeg3QYSxAf5FeVWHDK+0PldsaIJKY8RW6/ytpuKXKeDiWEW
jFhZ2kVaGoA+31Pq8VYlDZhxSgVkgW/I6YLTfNDzhQXXWuVNX3vt35eiJadW6/xuBJSwSieTehB2
gwo4f8hI9MUr9XT1TWcfzhFDTu+Fq6xEr7+rBp8u/n/4om8WU7r49Hw7/OfLY8MeklP+NVtzZXve
22JUldxkm3U/bXVEWYrq2BurnoUcSdp1psVYAP1chbJjXC+TB8SvDAyldkL1GH76QRuS0eBzisF1
I1nFXsE0nTsoFJwMbJYmDkBnpJiFNtGmEPU7WFIUjpRyn486PYnNfWys5Uo4SLaRpjTzRqDiaGI0
DAc1FB+kdbjhqfFt3o0olplqwMbAFCEzjWm4PdoO1w3C6zGPmI+dZHnothaJPsSgZg9NzbHPhC59
b8elwbjmcnTcYaX+jx7fnQZPiRA2hlvRLDNqF6FwTx1w2ZU6Xg1ejwKnHaN8wLTVHm1lKzdAuFZC
uw65KKp64Zs38A0JfLhAGu9CmYY0HyRc8yrR50+jJ4rmlD1bBTyhmfpwxRlaCRXXqtWClrafLNLm
2twlFa1Byh+sjYcQvjxFM4fMgzApeuNP5x8Y/y3yLcwfR2ZpfhUhDFhWKxoqwJW7jYEApD2ynoX2
FxowH8wnwyPYADbYJeVoP41eZlQKORp8R+z1NSZ3wSfqRNp1KvTl8zRBBKicA9Y6+zYrUU8qROSk
b75GHd4AQrb2cUpVLXWJHbt7JmSQE3VnJXx+kOV4W8Hf6Xo83TBN2YFg0QsVmpTtTbEIBDRP2eiW
qAJhEGWD+x5DARbwQnbqXoxrZs3jQ2FLUsd4NqL64oFou0fwExZldICE1GkKVGhs88hhNGoBGPZ2
XKw1C9GVfadxHP8iIFySicWm4evktfMFVfs9jNvFCzixUGI8hH/PnXuMEhbzvTRS9g1Tyi6OU6Ul
MG9FUplGHN+3e/hZYm1dDxSqhYe/ySB/BXlqM3A+F4QCESq110nNuWeAmOsu6Zop+dg3WHFXexXW
9uAFU0p2XnA1RvZL0FA/d0ohhQNNc3hooEF3XzsMWRVlU4GiCLlcCRGrY9S8T3VxMA7saDd6Yx71
gZ7P2fQRzq1RTTPr1+UrMO+EM3olwgiVthKfNZ3DDHbSJZz/zh0vFXfFyxaBZDEsUs870uTYJK2q
nBhTxDeFYF4P9IyFljCxrEUGoNgYJHsuFkHnNJuH0HsbMmSDLyqR3OWhbAOJpzb2hI7dF9+1hdMA
AJhNJoDYnl1FLnwxGDx/bWcKjIjCqX8P10l7dLGqruCc1HQKPrMDK5/q+GMv7BB8ypSbfwsidKpS
/o1hifguVFv6q1Pcsx11bo8OSh5TEGrUXwpaW2W+A4qjyfT3FuzfN/km+RuOZpj99Dm0u8QqPkzT
hXBQbJrioOLVLWeobyGdF6bblcDeGNyeuEacAU280KIVNJ9mIB9Kzpdw3JeS5cFN2oQ2zQy/HBG/
1YVUC631W34oH5nFpYvTORe9cDf8SFXM46nYYDzLyIkTKRbcajfBREh7zhKH9fRjsgtspKrpMNQb
abOC6KtbIvUYZ88d+efarvmeT1Wfl1/mU83WTsOc/FclmpCWvUhAxV8dUApQHD7nxm7mdbMcidEW
vGr2S4UPM4NdAmo/TbP4T0atVIydIqbMHEGEhrXbCVitC+uP6qefLOJZplFo/3UppS+g30uZVu+s
BKv3rcOdgj+KyW002ci0PSwLnuAjtF6r78dS8ASJWRTId6f87H7oLknXuDf5mP7C3YPaw4jR7ER/
wV0zbkoj4TVDSHyRmaGS9T8sLyR39EhyoOTriqgqju2nfxDXXUHZ88vzpDoM4ufwIAT3XPJPzD+d
0qZ+W6h76LH6WnikAwIzFpVehRR4GlBxoItQYzAignn0EPE7yMi90iR+Fduk1T3apbYjmvYKBL1X
YhnErVpA2dN3Ag1iu0Yn/f3DzCSZL+pI5bMiHX1x890kmOsZSbMzBifCs0/ME9C72ouqt5u1xzPx
/migiEDGcG0gaXzP1ac3g3jz+Cv/LRTLhekEReDM45CwprRLlJiVdKT9HzlCxhMP+RfUttNJjSTK
/imYhAXQzkkYq2o18giJ0syUi27bcV4FeD0833JdHebRp9QjDJ25QXPWat10YPleHUXH7Ytz7Ep4
whwG7GyfQCSbY4LBuzTs130DLTVaZD0AQEJ4aee+P0Xd6w6Drkhai6m2DRn+9ctZksnjT1ZezEyz
1/l/gw6XdzQ0Oimg562pQkkoN5yEUm6xy9j/ZTK3hDKrDREHU6B9O1UJa0G4HiFNzSRpy00VXu9T
Gc8vGjviJLcQJscT4WuaYaQSlf9l4UhVHOogavott4Uo/MS0ojHqBxfQhwz6QdPKBXAGqzMFEDVz
qCxHlsdkpbwFel7IPdk50kT66P8cwUZeFka0VIwKf1Qs9ZpFvKqljOA/wtqKw8L/xu6Qsv7dI/rb
5iGpilodW1anuguATcltP2sg+1kf2MhRh1UyXot0gRzr4fuIQZZvjmq/wrNtymjXwOU3XXo4OzsD
Ct0h8jbv350tq4cyEJrdq6VTw3dXyFXfcXTFOfR71vtPi0gAxEEMN5d1j/ytbdYkwonl6OUwcyX0
83/hVijl8e5HTOSFC9VWx2AgWrKz4mc1CjVQR6ucavKwbG5+jfFt6RsGsm64x2GFfZrYrWiNu94r
kLX4aw3FGHcq3E3tkjF9cwlHKTFX9fz220r3JK/LJH2WyigjuOHwPw11VObgCcobE+rLYzburnhk
QusA4zhFMXtlMKCp35GAhnjpEyq4vcG1hRo5o1z0qyiM90Z83efwcGjleaXzmvEUABQgM6PfV2Ry
MdGNTcPq0509xMQSbPBVDihA/rlNJZ1Zqes5GFwTO7OM0b5+d5xMxDhWUcsNFs5N6yVQlVxnrwZw
6QscHDXLdbgwgAIFMlh/FhQDHJ6YhtnCRo7EHP8SIpcCgCUoHmJ5Ix8bhJA9XHZS3IfjmbLTcsNQ
NTAXe6V8t5qtlVQdvalK2S4qcWCacVeOXapjP38bHB0WK2mMrwBaEWQBfpgjqFrdRpxwPQ3l5gjS
0glh2eTUnaiJKnvcD0AuJSXvH8kfuRcGl2AI7kCLMk7rNwY2w9ybzdhgviAGptBdT6CmjRrMIMvF
NtUn0v2XXoo2zePHEUDCOiMavsDAteDly8qlNlR5BsWH0KdnyEw99GTv/5cwfa9Z7nyEIx5CVomq
8SCFIqgMNt/6F/oLmeaupwXn0H7yJmkfeMDVCncj3+qroOffvjrpW0wPZXuFRZfcEwEBHcsml/1I
56VmbjXu586skgOUe8llaTT74eAmSuSBdN7MS7mrRNXbUnquW6LHk4KETyBkjKUqPAuFKMZtGUoa
/qZXmg2zTD0aeRIEFd1bQhak7vQy16QvaLgeQybGWSVKdWPdC1K0ocDwhWAV4RD3rWBtXmreyApG
cEcz0Jfoto5x75jav8tcSB1rAC2SAoF35JWKYCvUUvAbrZN2dJ5DObUaD1rkGJlTsQtW1XRBNYNi
ZOdjYwRr7Chxee7HR2S8SKql0ncxcS+aAfrvEES82mrNsreAWtZukuwo07U/otudfIfXy8UIKbRf
olDsVpgD2I2LICrVCLbkOh9td3g649rxDw6pki7sKUoropXNUnaJq78aS+/3NVohFCDG6svn3aYy
vWxOkfXZb57ENPrgfWhiFhMyq3RiX5Wq1w9ZPEVMbqQxEbS3VK7KAyouVPd2c0PcpzU+DJzPUCb/
Fops23kd311ujqxNJvum1G7rKu1HTOLTkD0Y+kaXcqKY5QCOoElI1mmXFmQomSReFUvRfAxx0n3W
ueYWoj/GwTibPxaLyRpveHUURW7abuUQ3Y0xl9hln+CiAcYpDZVLooOqQEUEy6GGvJ6BaIpo+6oa
+ZdRwIavFl8Lv6KJoQVPYo4LCHeVWXFuocfECygetW+by2xeJNYVLlV8Mg5b8pa/a5oRBMNVCVX6
nrn1fIT4w40qA6NQEKNcuribXpPX5YBFQqHE/bjWv1T+5584G4TtCDaF7ord61RgzvbOK+oiRHP1
kLg0MqCWmFB6VnkiQgjcQWEg32eA8JbGMCAuzqWDnnhH/DK2cHlOEntWeP0FKQB6vycJpj++OFl2
AaGJKhcklucY9c4ftjmWwm/73wcvAEsfLr9pvu7c8A6Qe67s1PAIA0FSSTdvoyoU+BBUkaGYAgPF
fNJpMja4fCDESSqrAVUs70S8dqPYz0D8F6957gAzHviDzi+Br5388YoBbMX2XX0Y20GjHkRpbI/Y
0lz1fARhTiHFVYf94beu3y5e+TLmx7cCWtjW9Y7m5F4UI2R4SPUmLewri08ZVdFUA7mnJ1tA93tW
IQeQV8VjRvrpfpq41MMC9Y/V+8Dtsx2YNQQ5OnJljegb7kRswVuGFWQ5zGiSNZQpynZ8YMD7qCCE
VuJekrzkBouTg1+ezAhAfvZ9SOUbnmfNg6rt38ec1t4iA+9+5UeV8Ir+U0KILOdWSXGnw/Q/9Ahk
wlvMEY9qCApuEiH9p3RkyQHayXy6QOlnW0IVpelAAy317qC3zsukallS2rqpQdj2jKTZyFZ6Lc8k
ykt4akUumCPLoLeWwXRx8itKUFEMZJUSDIICuUqwu9WhspZ9k2AYgKSUnz+IIz1w7GeiUFHIt+xE
lIKgv5iqA0DLrv/RB5wdkqT4MBhJ6gnL7ML56BzX0sIPMOFbZI2UOwl7FV1/PZ9KXiAZJjTdKfbZ
lXSNHyK5IcvlQUmw6UKRtw5tLJe3ViyXtH+FWTPI4Jp+pkbWJ0fGnWkTuxk29jPHAeR0yn/M/gBp
rzDIWKpoJjOglT0X6iOSg1HSIBceyp4jMScpWtDhfTA9cfsEQPHxBCzmtVZmf5NDCysPTzLsWn/n
brQ9VrL6xckj9mwRwS5g/Gt7S2r576UVW2dDW7NIYu3+BcppoFFvV41qwJYNPQ5+d/cs2BzE0lxy
asO2mIOy4mWDIvZZQz5iCN0NWUlqMgIjfDaPz8DKD00qZNpGFeE/49rODE8cJC5CeK26v+SljY3l
XKW4ArIQPrOJRwY/+0dutJama4qtNIZx+fOzmvPTRqjvOoJivTLatIRhOWquJFdRlOorcSV/wdd7
OELNc2LeVq/xS34gaGpo6miaogOtqUmg/35EGiauEyi+EAx0YNiwH63oPYOY0bNYTSXQq601TxHL
6BdBPYCcdTm7UzfPsDeWzugb4X9nI2bqWO9PvFVg/h/W2MNDrnkzDeHZpAO6qgEnO7kNBkH/j3pH
PNw33otM33FjG/DZIuq6yMHVOx+FnPRFtTm8SiRDuF0Nztc/2dYY8Lh6Yssp/ui+G6hAcorO8MP1
zXodb+bpad6ehN2/bSx0oyo3QDhDSR5vkJ6q7+H/1IOm31mOqjOCxI0h1+eeUBKINwSIMt00Rhog
OLRfop4J7V3LdLSBcjTy3Uk38GAJRoRp3V3kpYlxEgLvDCMtJ9/jGh8GKF/ZokjiDayf+oDa8lGJ
8nk+2+Za1vXMnjm6Lc7He7F87imVkxDSyrdptSmX0xAIqN3Hz7xElL7hjVutwMJK9yk1xchwrtKs
iZoq7kCJ4YxexhHd+xXn036rllF36iCBxryXLveymyeACDNMTklsA1tMCDhj4HegouWpNuQ+SOLX
5hb7DN8/SQ9LQaTvZOcZeJyXueATaFBijrOVcB4xzJ7u+KgXxoe5OvzGDkls97BiaJMT+yeUzysx
cXr81A82KP/Y51ZbPwb2LNkOgQKKacfuolfkupEM+T3dSyRhYxJ1RwAe9IBAqCQ5GKCZgZN2blQt
l40ZeMd2tR8NJ0zxJKBpWA30JkAbqbs6rczUEA6S43EqZBh1UqyUQ/Sw7SWX3hLzHR43i5JOBWxC
pwA9L4E35aN9hxoCK3flGm0A9g5M7ug506ggXZa+P18Hkaet1Z0HXzYxdhE3FNUKIe7Ny/mPU4K+
3iAZRqq3wlr1AHzBYzva+luZf8xfGs7d7QlAoz/d8dhY/Zk8hk8JZPedC0X3J3wfoJBkOeQQmmhv
M0KpHwOTo/xJp/mwS1jt36Ih6xBM7M6Klg+nw5y/15crr3a3CALYuQPNAtF3Xy4kV3OWJ45z2VbR
TcmNba2yNOs8bOOWbnZIQIZ6xqpVbD4aXh3VrnqBBq5YunoA9mIP58TYlOClIsY/l5IBz/wK+bGx
t1vibYT0PaF0F15PCz8VKtlq/4YqtE/6SaLBipMUCI+ce4VHM7tkq1j6+QPodPwZiClt1+ruaBu6
bSgg13EJitUXWXAc1LqLzHhhdXtTsEsQphlqqKbwA/l9KI07gq5QynRlsdTms/VFTBWShTpYIPro
tPwWUZPH6eIa2lW4uV4AqUmS/79rB3v84/whq7Zyx//FVv4uz7anK7itFDrP3HWGnoO94FEaxM1l
qKRyy1P7sur4lFmd+Cxx/fw1IQ9woP3pI2aRlbQjXL4dBOHBfnP1syVyuV0zbR5Qdc/yWeoGBT/k
lyjJwYVgqrsSY97b+VxFVrOJa4BxzEhFEDqUyvsKO4nh3fz+wZjUcsdg8/yl3vj6G54eGIX+L1o5
qsHGUI9IcVTRPMeoTL5Rphzq5QaUt3VQtDjTJJ9L1JsN+Wg4kD417Ej0e47sdpLYijmo5/0UImCw
FFtRrxhvcIWws3PbeD6+NUOcyx6BoWqYlpNKsmleu4G0Y8xUP4bTGEWzba0cUXvehDs5CPuAH0aZ
/ih3scIMYkbKtMiFm/aMtKFr99YNGEBm4UD9YFh5QHsW5d0WNaExhp6Adm2PYLDdeaNG5C66LhzC
45ulI1ZRye3osnduraEv73d9z8/OvOJfcy1MVIwcEy1tY8A6xOFBLMzSTaeUfoNijQ6snSEA2ZA3
cN54dKSiwo8pVPiPAgJkiPsNuEIEnkkPXNjtT8i8gcqPpS+wm7+1jGzCF4TePtmJVombXG9MyNBz
J7A0xH5eQi+MnVcMCLCEba6AF42QnYdxboIZAfVOtqiT6t7OHKNPwKXkXFnSfjQhA8RkqiGnG/cr
603sjzIejGlwnm2QDqRsZIAhWRikhtAhmcZACd71zr14Cmx8/EG44fcUR7f2SRkJsrgZlvghAKqE
VqMGOe4gwwloec4tr9dTMsqhg4cBRrYZbZfdC0MAIbTteeglqfHzgqUAaKM6L3M4qKvVFr79v8Vy
t2wlOEhcarrl+AbAIuk6tMo7N77wKV6Qd2jpD1CRPkJK08dj9gnLwQMitsfrVvRKS0DhOzH2zzrL
+g9hgI8iH4i5euMhADHqCFUg59xS1sicNIRX69nbgY7bVO7V7wjOhnRHWfGdZhcLvqsHBO1FQexK
vkuUp+Onre+9TbR7D4219EkvAU24ty9epiymP8SLFjwwlESQ6cLycs6yRgGJ6beAiPyQ2owuSXEh
BAxCXZJnKUs4aDseM9LOssWaoEqU9w5oFwN+p3paWPHVUOmIL0kUaND0PV2uY9v1cR5V9DmM1OsT
U+2dVhmeXPUAWRli0cf0bi8k6tCwrNyTVPntrq4aPAbBYMeAhZ3fmS0gOOXs/0q0MfIQpZQBQFsk
QDvibDgm5P6bH3AA4L2t7wObI2vuL+je8HOW2zLL7uQoGKdT7l5DTyGFpLZAPoL1ANRgoiNeXQ//
LBgeVYPYpxVoxZqo5InAss49AmPPojp9D5fbimqr0hmHQPDAeJmiB2sxm5QMoWurgULo7ajaSrez
PHcdYNz4Jahh405jOxFZ49LAkwhzBNXsaX7uDkD1lDuo1D3S3JQq/c5+7XXL4tzH6NLujYGKJUfn
HZjHYZEPf6QR5iYzSsywneKE8gSFK2Df9ZOcKbGZ/RgK/sP84EVphzKA2xZLKgiEsWRP7TV/P9Xh
hMIO2QGsWEcW4OphP8auRGLKdjbnGRguNPhNjhtXpfij1QGg3tiLbFT3KyQpqIIyKZDIl6wgs9mk
M9MQLw8nBQB1hcwqk2b4QShfKjatS4mck3677mE9yWVkUGRFp0h3R6Bd9dv8DHzyAoWD73fq6fCj
g73UJmNqotSTFWDvFDQHTu3F0BKInR3Mm+kUKRuOOtXSoe8d/v+dPs0QCaGC2O0fl3e86dId2+Tl
soEx26pNo103YHVO1M53W/Dz5mhhq8MiUvJkQjzxN4vJXKD/ks8YibMQ5Udgq9XOHR8lW8Y12YNT
cu2V/cJwBfU/o+plgL8yut9wLgyFkoEwZqHp//IsTNxEeWzb1s1vDvjmhAijrfM+Jvfabwbv4gIz
pyV2RR799Rfv4rEI/viu5qJXMCj6lgDZojmM2tmE3w2cbojci3zvEQ/579n2UBPt7tWHyobJvxjQ
lbi6egUBsjPt1raDcBcrfE/1e1Quu0OH/qrWxvXnws/ZB2J0p6dnV2VOFBnSpqTh62VUXvc1bK4x
9d5Cljov/lGYVFPpBp4Y/CWAfrH4rKftVO/80s08JuLDw25MVTUMo5LLEfFA5X8mmTeVWF57E1ua
AhDejnN47lEoFxmKqSZ+WD+0hJOD15H78on7OHWT/vQATEpVbTPXKZNgq0oQ8OUXllJGFRkkBepz
rdb9Haf+PezePJ68sytRyI9nXSsc1WRMA8yDVcBQkHCvlXVM2rNdp0gzjrUsaHieN7wVY8Y0LloD
7CvmTg+Ou0mCpYyFeyTiIHNCUvOEiB+UuL199Rthrlt4adZRX3JVoUyd8dC/6wWWW/SqBW/KPpY/
nAnGxL1he5M1Gr/06yxZLv/bRiDrmHHgCE2HpRHvRlfdxR6g+CGecUv2wVRDroRmlq0EnbgyZxiZ
D7kc2T2IeuAxLvQVGaZqPQw5asOeqpdFDuoc5sSTUWhzhjrcaUzP0ChTRSMsBujl21GSxlccFjPo
UxwY5CvYtJXjfBzchEtMr/XNaBH7edIWyeZhhXgCNvdm3kn3xlIX3qj0iZOHSilraQULBeQYzKPF
MfPCOxCog57JjzlDlclV/Kj3nLeJW7lJe7z5ZeVSHCkohLz6lO/eTdlfpKANCWxfp47VSp/r6doD
iLMduTrNyU+0ELVUHXkgrOWUaXzgl/kJHlEKrYuSpFl6PVSN+DFie6/QjsHOBnW+mdpSk8FzoDhW
BM9wxUKV2gL6CoKPbbKzeCE9wzr8Rr40MhSF5iVrjuqiSLtu4JrEiD++HPqqxDITxVnoulIkzPBE
La4mp9iZPdr/y/WjN4fhsjLKwyjL5o/wP4MXn3+T2ePzBLa12HkpAcmDOwOvH6GohmW44dI3fveJ
zAHqUIMozfVs69HX4YRUHN72TDxKsvgGTwawSpdfMtPtWRWjzZR9UOxZgB5GZAxGO7dCUyxHxx5Q
JCyqSRflrdYTWbQW7MQZ00ZTOvNhhyNVC1Y3AIG0Sx6IiXuUXs7Wsm5Qlk10RSaaEdKmlY/vAWxK
RRRJVLuifyrm0HrERUuDXGbCxxrZy0YMwJgKnddejPuof0/lHM9YX0IFPmtoLCpplBmsQ0FdB+1+
4e7uzZW8ksvbIkV5d9IdOdk6cLBv9UEXn7BJMP9Dgj5hIeEaK/lISRZxn5F2L/5/9G8Cod6xAOlT
h8CS4hiUDI31Lc1hUuteUks5lIxd2gAUTC5CVeQOn56bl+5lR1EYGn9cvvAFHcFEbOyMrr9wqq5f
nsBzEOoqvJEi9TYj4aIihyP4X5AVd5ckGIwl9FONSMPL6X7TCNWpqRXA0TcRoRsfVf9KMGjQc8Ck
zIzCOuFfEJsJExSl7Y4Tb+DEkyAHySiD5F5IYvPjYedag7QO6isENRRCNw7CUiJzs837CAR8n5Po
hhVp7LxuAtM0Xefx2jELIrlSK4lQ0cVAT2MYuwmJ9ton2Jf9oNSi20KJvq8mPk5hTp/SC27vWbdI
/Rdq0F+eQeFSsknL9YoicU9CQFvvtpuyxHdddf9KgIRsi9ABVf8NS9Kk3f/li5cfz5WUP02Fd6qu
vidmwJa9EeEV4/+TEVq12MJ1C5TgfFABUoI85uQ2NKYkqBPxS6Di21UW6ysB9OwE4lazDe3canFb
NfQhJwhT4gcvVwfsFm4az+u0zSLUAZx+jDx6z0Ms7UNQJQFm91xNMlkdQfTkUbdXP8+EhuKuL1nU
EIfPfSdtsVV/ANEDzV/rJlXihn7Zoqs64haTvuyJL+UAtG2ltcuRuEQxQ2RLwntBOgyGTjNlS216
TxmtTZG6KHHK709EHcVExPUs6XBgrM71fbJdhMqPQT+AHhRQWsSZFDwmG9DQYbxVPAFP0jhQNGPB
f1MAcxEwsVFGVAbU2quir8j3uoRd2CYevm3YG3pQAgioCnHpZ2Xnwext2NOZxO1kjIHY4Ooa7Or8
qM1eFyMmD6QTOI/wZZByh1nLVmNsX+EWs/EJlYp0t6j1u22+DlXFmlyWZF4/HkXiIQxC6sNY53zA
qiIsFyiMvGq+akLvcc9dMyyR2tmbcWpPCTNLUN31NiyXEUpgDKARf7f66rFgk4UK48aEtmnC91C/
7w1bOky7fp0IDxDRlTP9caLLD8+QvR+QZOqDV7BH5QzCMZjpCaulZaEEB9R4TKpnJTDX2LgQnXRn
ueTixcRkNY61JBAFLb9SfVGWoT/dAdY3m5xIlYR4+sOHyfswZnqC0Ak2o65MzREbf7rcNM312FqN
sjkWQDCx7M0tr6eis+FPsRWhV3fskixTc1aMrXb5tahffCZekZcAhUyfVR+WnRUPEbbzJ0v2gnIR
phEfIr4eINAG21a2/psztOgC1BYs3QEo5V3SK1ibifoSRguu0nd7cyfoBVWMsYgU5ioOd22gAf1u
F4pPSRHJLDC3PqCta7LvhJpXbxayBJKrSOxl7yT+/8YFxHfYnE85mY3+kclwJvdFHTRCm7rn4+As
uay3tE44Uhj1Zs8kYJXe8qGAKOPnFJ7RRRYLl9mxt3JKROVqGnbltghKpqMJlwdXYcchPCUzhcdT
G+HCUynGGB407MXX3QZ50gbDINYMv6XFlGbL2SYMWqHLs6buagK9LL0BGSI+gfWptPqoUL2XBHIa
d1p0lSNeI+ozZ+PRZxi8ab40PiGEUqdWVuVGsb770dK/QW2LkM9p+EjojIFDnmRoOYk6jo+jeECw
ZLk+muznZ44OZNryNyA4Ebq13gBeLSIpdOqo3wI44nWyPh8vgCEiBHdJZh8VzAKcODY5Ta6454FS
XCZlBA60yQTFMKPAHc+9vBIKs5L0q9JvY5Pgp56x3e99nzvs18CnZRda8LlHEiBrUtuQhacyTkAk
oT22tv34rbTWBXBp8IOPYr1un6FOuzAqgF5HAFY+raopWKAzSd9Z0ELyYehUoRfiXfDhI+zKG2V6
SYLq7JaHjv/Doag1RSMhpga3/qQnxOIj/EsO3Bp2qH3vvt5eFpG6+UGAAim6ela49n1ldnGqHPVF
Q8qGszdNLhD3fpvzPMY54Rmp8fSNaTzTy/3vqY1MdAJCkDgcAE0qRbsqC99u49LzbR0i0bUEqSOR
r9LGwq0xRJb5DlWDVNcaMOFLJDJYVG1jcw7VD9dYclbi/11P7RTatp3NtP0I4S6onaCA30DOrv20
hjwpEnEU1G5gnOCigzIdBzjZW38YcPo5/N0M0yYbsSodgyG6RgPNUAVOf4hDUbhcxl9tSgzhu9Ij
0nlZ6rjg16trpdccTUxvBMo9eHWHClUWJFvDINDOcpEBaBh2AxV2yTHvc4n51RXzrxHy6qqKPvAn
Lj2M3i6Z75fYov4RnmVmVms/kNnDmow4OfBunGU0812YH1SxgTdOxcMGNWNG68Q5mrzrKJD3RnnO
EZqsm9Sw/fU5QM7/+J6kJvjbUucY9PNDF4GJHclwMqTRD6zomCwYSLKZtHlx3F6DH4x6p33dl3hs
Pn8hSQm7VR2yXXdhpfIZxGYjt3q1e8U49MaAhv9Zd71WnpSfOr53g/hTfB1gGD0aPEAlfMl0filh
S+JkEB9XHRp6KfZ2rPeetOscjcAB/wfh5IF9tz9gxtv7U/z6JHiMKHbrfgTPmJZgurx1nJM1S0Ta
QmSrvKli1RjLbXmaHyiNOP2IRsneUsvT0YkUX+nWmWiEPdSLaK3iOE+PVjNUTgiyHaXfQohlau/r
U0NlKsom3XwjSBPRN5a36mh8VavwazgENLGIxI2GisvK3YJ5vKaoBzEdC5xa8zsmR7NFBVq58sIb
lixQB/lvfsiENN6BEKItmHHzQOaoPXik1jWNn4c54Sd2zD/ElQ1JZo9hRjxgLCJbS0t+V2WwFS0i
9/jpwA90bAP4WOZp1Xhb8jgL/scsOjLE0QJv8mRFUvVErfE2D9yXVEGUa5NbgVG/OvrqRPprV1EM
1MVXM4hLCA/SvQlocfBZNM2VNKHF8E9c0KBbAM7AEK8egD0GmIzFujZZtSYDVc7SUNL6vwUzSc+7
4QdJAvnsbWR7gFI8j+ymKNiw+yPSoMc/+oklD5jnrONZfBQBoeQKnnaUjZuzXLDfRqGg7Rn+tY14
1LOe9OC5AGNCRYl2dPHlopRbyf2uf4ugNSkskRAo47g13BQeU9DfyIl9cdRHyOzfVhQhjdqTJ8+n
Y6yXzbGDPezyJXVPgFSBPq9Y5xqs6fmMuFAQOtqC6QUaBhj7HyUuJ21W4fVUZZoJsz45KyfD6siM
/BZ5VpTpX+rrrmraxIJ1S9Ufmm9zaZSgKmAamEJFzef/58dpIqcWJbv/tLGZCyCT2uqOnRNVOXaN
NxBjAl80qddbhk0x+VS4XEznoY3cWFWusXWGaKHpgrmNDSuYV6daHuKAcMgSM08dUiBgW7kcRAjs
UrTMdmpNR9LFlmelGYiQaB4GNRMokVjgvMM5BxPuq/JO9j9fifwvSrLuAUG7TazBPT/ROmAZNX0g
rFm/qCuG0izCE4cJg6ko+RRedJq2IbHCKS/BUGFxEY5g+LrVyU++NKJ70CcK08hIjDb3lBwpA0CI
qHB3q+RKNwY31I/dffN9kG9BZTuiX7tLtOBFiA+MftunGxGnQNq/8Kpstz/3fyzuoyIQK6tMzo0M
PfO9ujTiER7zBiR0O9R/iW072nfwxB6sy+L8fUx5LJSzUNkAxRo/uJBPHqmaa1E1bAduJHlt9Tg0
cnEpBMK9pxS4RFMKgWwohLvD5VN1RjztnivLycx1psGm3QN3uwifjrLZGiWavGGBt9YtTeucQknB
H853Cw3lgNYnQSOCf7zrtRV+mYHr8zIAm4q773Vj5XUwxnd7GS8/a4xgk2GnWHH24j+seWjnsCgQ
AY/IyGfSg4XhV7YOuDO/AP/zxyPvduD04zTU9rX3PynrS4p7OaVc5dJbciF1yX4HCOSyBfWGUy+i
4Zevvn6AtcXToEtzgfFLNJlozq8LxGRjTM9UM3JOmChZTNJDThjIySD9falFw3K/qrdlGidkxhrE
Nmp7xwLQXy0AUrmnEk45aCSR0B/PHgY9G0jJ58vt7lmBzC2xEFbHNTz4w+rPxUFUkRyyrU0j5uhD
cYlNCGj7g5LwejPm1SeHPdY7x5tl3CGrHtIlCn/kHF2/pKG0jD1V/odoghEHMc5gnb7aRTHlCIAF
+DPYgC86gET4Y4zTiCOC2fE1qQR9Tx3/T8HJLAqNYLScJcKQfYKHRVIG/ZLYRgWgsyWOWAraPMix
qKF9I3Ehk89qNzSR9Dy1K63cB/rTdJLovjbKts78DBAgssf8axqAmc47yV1hgutYhjuGlaW5QaZ+
6LWP1hbUkGKRRm+F9apDcK9f8vcEqu+6gO92QSUnCNCns/YRkpVHj3nsC3jAIagqVIBlf5Tzb4e+
HWTMnbBRcM0+ZjCGR0qrnqvVk5PK7NKKBlQKwOMc0lcDGXWuPUPE9Oeo0ZaOc7id9d/O5qJq6M20
xrWxHHRhWw2hiC5gWwMih4j8W2lsW9zYparzG40+WbR3f0xSW8bJqQ3tw7rvvXLHd7sDKI8xggrx
OQaCccR1uctv3U2WsWXFI9QQhVEiVO5hkwBK64/amx4Gk6A7k7krxQkmoGk0fr8hKxaFfJdqptUm
WLbibrPI5Z4DSEDKNxnusvMslcdh4ag/4hQ9p4uxFcHWGApxhV2gfVvDi/JhLDfCZS0I13fnse/w
If04Qo74Xd8W7i0dzkKwScOQm4As9Jn7R0s/CpfEL8vTfetH3kW2TSv2Ao69gXzIOYxWQ9GRBzvF
YRql0FSgZz0nn2c/irt68K/fblMaCI1MRt4HoMGa4lMP4w3T+OEdrbjNc70E1G9Er09FzdUvDjkV
ZRNGCxX8iK+BJ95l+GbYDjLwJNfmhLSxgKWLGTaVXPNwAcr4IZR7grP9XDAdLoOc58Peuch0TKco
U2GcFayUoM+kAwGslC/b2J8fgqx3YqsiUjPNfXez/+49Om80cpcyG4h7m16+JSqTnPh11Vh+UJqf
vtXl4TjoeULjOkKcZuEDKec/LB840cLvL8so3n+m9Ef50ecd8CK6VEmEA/IfMTSENB6IF/QhvRif
zg+O6PygCCrq/ZiKAw9u7sTSM7uaQgL7tcYCODgw28e/7v2S8aFhwhLejpGyQcy8jF7mbIGPI1Uw
ZvQlEgLw4E3lJpRSIN9sHfLdx6F5oOcbInaBBD8nj/Kl7yywG8Tc1AIkHoptPBxIno4pSoB5eQ7a
PH+rQja4P6WkUDJNz3h/JpZNfzjzBSKgJst9dHd5qJHkv+vY9vLm2uZmGE8U4yLkLSRCwApnW4zR
SfwrbF2gUuQskSKAwzT3b/6dp59pkHYOZrxPns5t0zj92JGeTIf1zz4bHZGgiMBCbS+MMCQDx6lZ
mUHOc3R038AIxiDLRitYPnxgfWGtG65eWUcEtF0UX1eldSqGdbQMqNmTvCgNy0Su7dEbt4s6jl5H
HIcpCnOPp1d+QEOEm0rLq12X9ENfkKUb5UvCheWMuFObEt16E2ylou50rv9NOhcNNSPTpb5Gut9f
aLy5QpYXv7yM4GNH10ugU9nQVlu3iVxBuG21LJ//B6YwJVDNynWMYt5P1E3TDLs/xqV3gi/+tOqP
LwzgtDmkHbk5SOXZjG5FolDsJIwmpR6uxTFCZt9SWYLZV0e1GfHHpA05JLmjfGy13JJ5UBmlvMt6
V7cflMS7tZZd7vU/a/VWPi9auH2Pr1BRBfvp/zPwSQeCirnSXEwBC89OYmlxjYwC7d7IFRl0SBEn
oWlVGmiQBJ8XYHcg0HkiqZIYXtGsiINzml+QS6KxaSEBPy967qworRJ7Buzpe/GNhe/arYGuGuQr
M22IM6bNXuDvZE0t4I5WAcogkf9RAPZ6cY9rk5kFpjUOCpNSXUjVoOtAY+gClnLbxrjlWhReiItx
eE/32hCLcaXVu4DDPWnshta7VQrevyK0odyHfkHWrdYwtXj6cQ8wOkuIFVZ72eyFQ5kdvWJFW0O/
camlQou5zpVTNfwzJ/vZdP13GxPaRSmFI6L8V59wKqm5htXs0YbcBNaWKlJD7B+ZeCmg6hGHP6RN
3qcIMa/3AlEQDyHtLOnhqhEYN9hsklni6D3ntZ7CQehuomFjwrKzAv7hMtwa2KIDiZIgPk8d5TG9
w62h6obbVO8Ak9Pzh/yve1zXu8i0A+9gEvj/I6isXfZonqUz2y1Lh+88LpeRvvyV9qYTd+sjp5mP
WKht9GQzrUWlj8dHsLVBl4D79WBNOqkecqcZ9Ha6f1D/R77Nghc+Efat22RywqLOtgIM2gw0DT7P
k83VFKP47rZBKRzilXi0zu3inH+3911DsrOSL5om6dzMG7MB1PRlz0a8Gn8hgHkxJJr5VUZzrFS8
SaALabuiZca+porPCd1Y4tNyUxySa9ka0KcX9vYvFA3MGgH+0SRojsNcbnj5RNjNdLTmISEaFRdp
12BGOkTfATKRUQG2DhFpeAHiKpQ+YUXoMeS4yGnsA3z2B3n4f1ZCEU9VTNAebhCuHo8FaM2oxmrP
CoIGdmszWGILnP37jBlQBf9DShKd5Roi79nCfMPI3D9UmQJ1s+BL5qqR4aIxxOsbcGSzy6N5spqa
QB3Ss10JSH4/5Ky3HPE9VVHKsUfy4ONtyNKPhsjt5OaE2m0CpI6ZoLGDvD+d+cVm89Vthc52R4XL
IJ4r8mlTUYgXdK2rxY6RgkZlicV3qZOmhf6rdu7eV5uf6jM96OUH06mb+H7fWA9Cx95kqKmrEemJ
wYqbNjPyEiExIYzmiAzgndKwP58qlZ0EAHS8itaN4kmF4WU1JpiWWoCd2Fc3JtqT5utebvc4BGM5
2V7djSyNanlcVcrT5e9Of6TAIRK2evbeNC8zgqHogJVvry9oHe3F5KcoPvovX2y+ibI7A/s2LNSt
/8zQBBZVHStNZCpvjOQegsN14i1+QbXANHDYyA020afYyod/UkgpGd34ndpEpQMRpkrF8SVbSwHG
Bc2xMUuas2cgEFwnAu+pJJ3/hezHlNI2PK1tGAjPUUG48ApmxQPzbpl2bXL975RXjjPFLZgUDm7V
aIkkHlNvWgELayPDwXptXXogPy/rgvgXrBECQgdSgAQ/iZRjgL5Qd0ci5+DqfKg3N2IYsb7d8szb
9taxW2H9ikLGliB1A8p17U29qEI28ZmckAlm60BhcNjXEtQhkY0vyJaDihJZuHUHcdTvsg7KhH0r
Uce4IDl49M0YSjHcKBLC0BQcgmPZQKbQE7bwi8AxoPQUrz/oPcStCAlQu3p50xiRfXxRe9LDXHv5
IBbq9Z7oJOlU4NvJOnYAUJZEpkITCF3uN5INXHnY25x7GkJ2txKWP7WjPvBjjOK+Q/COvokdRcEV
DMYF4eRNCyPuHBRFtLqYhv8tXroZWB5jqzWMHacLB2ILiAAhuSdrcXvw1oqAT1SVdz38tByxs88I
u0pfCBEIC6+L0Ge/UgJqnCOBRHMo2woCLLy3D31mq9auRfbQRdyOYdMvmFGKdUhzau9tBXcid32A
wPriA2dkpatd2Cx0VDHf6PzbgUIK29BAYIWG8XZbB9JbEWWO2cl+IwDjWqMwXQ2BlnsKkJLJf6Fd
ye85FsTDwnViy4m1LXWUT1v5NUhFJ5iRnq6mEmADNvp5gB9weYf5SzF0Xazhg6iPYblpJJody/e+
KqNY7AmL8EoQaLi2UlP8IDbzpdUFCMt3VnYmm2B4U1330uFTetbCgZ8XkRtBMyH4jEsmqAi0JNhL
j718jSV2Gx0ry6lDo5t1FAxN8+IBWoV5KH4v2QlLpzGxgKeLSPkA9sqPUe/5rhG0VwGCm6GBw1H3
t3OW4HMIerPUEMknjg1ZSfxr4Qllpr+7NhJa/IoxJNzQM0iTKei88QlqRgotE70AOvIO5xcEUQOU
8Ed8qaLtuzj7mAKd6jDtj8D6fBQUIvAjrb96VX3P2u4Zt4YS43pFquAY5eIPqkRtbM50cyJrrYnx
gl1s8sxk4rzH53li0ViWXHj+ZpA4CMQNYcZN4GgxXLdoPchDlUbSq9Chn5jubfBRjCuNm2sqlrYu
VHDnrAwizlzavM2K1w6lUtbgPcgg9TtKGANBv/YiXug0oUC8736jbW+gy1Ds0PbdkDnSBq0PGmBg
wodReV+qQgCxb9rQuTxtMcaaXYJd6oyDqDiwJOLjEZ9uTHjalNjdcxxFCfEIld1cDmVzl8cM4kR4
BK+BM3p7Gdl8r5mZqdFdTxrJkMSOd1iuaGxkQtIvLrBuX3BjLs/mVALlt0aKyg4hKP7RnCnGs0og
NXYu7BVTh11Sz34EqaM2PvL0XrA8tad+hlK4tkiP37sTsobLiHsCSY8h3wkMhCSk0vvSHNYDaaA1
X2SfFjHzupsdqwOBakRKqFWThpViP3tF6AArxOMYDUvA+MCoEieWYajrOleVR6O/LUYPX36LGeU8
sCZr07WRQs8YJtmLDYatq4+q5UJSzxBiFTaGDo7SuywgxKvviqifqLMIqHZYIgnMR9AcBepmB92B
l96WJUKKYwXZ/tpbvWGG2LQ+pswEv0GcRKzOqeGR7/8qkCHMJ9nOM6Rk5KdnFBJlmqd4kBD7BoXC
kllrlco07+hx+wornQUE/C8zZDzDxQsYdjXlAj8lkIucrIFtC7kH0TYK4I///6wlTtwPdQLoWQWq
lPtO+YSuGDJIyWfI1YqOgMsgNKvlY74TqaruiITbMNo0uM6SgtJ0BmVDUC62c1DQrMwJndsbMlhT
Vzv3ULT/BfUbEbZmen4mPkYhc+9OvQOoTh4LgPABIv/b3slXWQgx74wmyk8pmUZmGtgHoCiOy6pQ
Wa9ALKwhlPRH6paet3tmNjIB5gH0QLO7SbbHzKqX9WXfZdw5EJvTyEt0YPRSnmHiFXmzoPVXqFca
JvPAcb307ktkc9Nq/Rs1Jm0EF+//BMV7QkPbzinDaxFbWNqd9cAj3miSnMdIktf4SRvbZYsHCdB4
tlKY8rufWlkWXuBSVUohT771sEzkxDPscdS5gzwM94fTIA0odgm1HW+49yMWZNc4naFp5viuD3tU
kr/24WyxdV/HfWx2PrETwnmQ+0QMI1tObaw8rg7YpMVJpb6GP6Q+WWIkNYxRN+CKIQmTeE2UI/LJ
/iuUIRUthVPmt5P7s+m6ZI06hLd9Ydju8NIrm8HdsnJ+RvSlp8Ro4dAUTDEbQ8KNipZuWyx7t5WB
bSVfjwykDkyVncdJjHGOspeBH//cUwTOTZ1ABUGI0I87cvbR40lk2fdjVyhqIrVihzrk0ukO7PHf
hWlOYWah7WIB08QkC9fQnYCsdx1e9ihT71Q5Q2eb5D8yNx3rvRVNmMCNq1PRCNzyyESnigoReVc/
+0EXE2jqGWNLxMq6HUHllcXH9w7pX32kwFXUXs8v6LlAosL7MSNCncPcuORx+GCWoaqXCSpRt4VR
9Ulu5sXqLnPEVMXXmaL/pasXt32TfCgI46m4ilDO7zEMv16BHV6G6YB9/R79QnWPQ7nCfLuV+Eg5
/mIV5bYmougvntVFkhP/C9vdEKeBebAEqvqkpfEC6fF0QZgSBUwa2tkQbIVw1F3VRKAWufB/B4n4
q2sR19k3e6D8syvWNu4FTU31y7h7Az8Glp4kmzUDIeOse7/yKAF04GYHxbpUmV4uvP+SbikaOPEC
XshMy7+qivOZ9RYeUh8H992ixfaHwCc7EafbggOw+PJKXrJGHf4W8poqD8Fg2vo3sww23wRNuYg1
fI9OcdYBZ7fL07BdStU3xigEmbNfphw57XCxFfIH8i7ZNESJ7OUgRpQ5uom0iRwEh7B5ylYCYpbg
M5LasiPFyUa6iM3Iixir7HooVCI59aUUvTHqiPIsGy9CntqK3E7S0gpVTP+aLIV9tipDVvy2ndjo
8szcNno68t2cB2C0jm4KoKzTxtM0pU7S7Hw1kq8bvi9XVHihMKieSa4KtDlkdwM6kLw6waNwvhXY
nfOBhAzf3wnT4q0492tGD8BtbS5bF/Lk8r3U5w7F+soTxF5FnedyaaJ/W4tVOv905FCYiXuYvcOq
+h64KBq5q7QlZ1EVyYNFHu6vc8p4O+lEXGWsTMSwEKUhfpzFE25XIjOwa6NRHyEYVGcuP+19UMFL
B6c6BxrSmMJZ080gdvtyjMFTuJWqrVI0hoDgrGf+i+kPcysu1uJtvvOd1EvVdeLsfLeDgpeKj8im
sqEf/WV+UKhQQYDj98O96sI/HUG9D0neqmdmAn9tDC/M2kBZV0cpJt4XTE+kcDhPJ1loMo6EQLWg
f/f2ZAfczqRbwU5iItd8P4v9+HZZO3hYBPy8+NW80+lYW+DBq7Vo8iLKLH+owsTLKTq2B68W4YhQ
iPtyeVi0w2rsPQ14CXGhAEnIxhGIbEqdJJFa2ttuKDgeQiiNlZyzJ3acpg2uL+dFegKKXETthO6i
wDYSoKdbnE61BSivsZYPj2YCykN5XJ1YchZv4p5h4wG7C9nbO0cUKy86Gw5LxC1+eig+4TwRI30M
Ga224Kt36mfpUigALT/E5P7lIdUbnLbi+rA96ivpYYY/yzMVuZ6HCVeSAW/LOZI2n4xAOgonfxAn
96NYGdEKX0jool6jpHflRX0FQoRfG+D9Jr1qy088ZPzxUlqAySoTso71KBKSkMe4CLg1RS/+D+12
nrAgujEVZ7PJN8aQImewqTd3Y1DDZKJ/Sl8AXPb7/qo5c22PGP3gKZXu9kJ6L7Tfg7Nymnr1YKPk
hZtQ0dYrl12/NkFsgfofZdXqdu1QORLw5ZNwk26hjf06KHSPmUlgFoPHwGpL4dIM7leHl6Kzrr6r
V7tiF2i9YNUh2Doa7VMJhuXSYYbMr5JOw4oMrLY9k1etV//4ZLCLvM7z6lSLby65xvUNrM54aU7x
oTj6rrYGzhPv5yyi3rEJAGccE5k/64EXLQyDlIaPQgDFMnevfSrnp/W8GgeaVFoLjX37uRE5L0vg
XkahCaGGSa5YYs5Gtbv959ujEKySXf0KGWUcWbjTlKwobvpsdHP3qD8DQs2yV7Vi7jYVDSnmGVjt
DHsoDsdIFYPoBA3aJ56rsIfKJtDooPx0Nf1PcNPmpiXK7izarhTlL7qPTTwS3zlJxY+0G6BKlZpr
JpQjrVglh+LhebyRjgf7GbEE1OiuxnlI/uYEqs7mSfa5PTI3DrbrvEj1Q8X39YrhSf+vKI3n/WEh
SzWn5WkuxtjJ189vbwA+H8p7q5OwSIz2wdTub5u2B12dfLF+qSuXaJkDbzvswjBHxiCYROqpATMV
9qKB3CAJL6pZfJLM/FloCkuVKbJ8T7UcnvLMKyKxPCWd6BsPEvUiVzyKo3B6JRut2bq0qyq7Vb3g
5vaywBgtGa/lejsLZEUnbFZCFOGDyv8zm04RRm2dBRPjtTeboqvRJ7/Anfl7sVr+rTCAGRAvqOBM
lQIKaJgTSK1RnJHXRgGoq3bELt5DphyWPlEGxqU/2s8nrR2zp1Kls/Fiwd/iywUTA3zzxvo7ABYA
SNDhMCr7EeuJgLEWxSsBgveIvYoMQnk8VgEk/yjZ6JfLn6rrQRptQ34r6/a2LsQoU6wGrsP471V3
FkYrjVh0mEKA/880D1yeud+wITWUrRbniczNT+t7mjj+U4ZBvwtD2i9ixW9CcnkIJoSjZksSf8pn
jRSSQc9TuudPhDm8p7JEjCx72yG4rQb2o6J0/G+mCf6AFT/xaHMHKHCh+Ph9yrjSsMTK+mGuyco7
Z9bMQ7UoSMgGmbP1gAvdNYPgNgbTfQfZkDuqUrRFqgcmiqGrBGo1ByNYP/ht5Oq+pGWIqRt023Mj
op4x2yDsWZQTSJcZM+zjl7t30pomQ1PD3T5RudBe7yanxi+SyGu3zTN1cB3/bAxpsoL3akzPqNbR
wcTg6s/XCZmwhPc6uyUPKJIgSnjQMwVhNFz8UJ8hbPLk/O+G5WX5ju99P3I1x3G8JOl+CD+MnYsS
gqZTK4ZamkN+COGx0RIpxOp19JjeRC7VAeSzZqrBVjePr3UjbisqhpK65McYgPtMUshd523Gj8AR
iar/6Oa6lW+6hfNRmd3s648XRku5nMnYGfo5ia2kzVH16SPKh3uamOW5Lw5/FYLE+b0BgqYCdYOh
HGJLfF2p8KRdQxfyygmYWUnLWGIsYFuuGduXFSpSzkGkK+dDNiBap6JtusTikke3YR1qL+/QaTHy
OQoWBmLfG9hA2x3cFyrJlm01z+fJTfisHG5A9iQ43RK3ZKZhyvVky/xarNf0YLXbd/+r14ZQCm39
bdgps6/qilC4XctoldLz3xFs9X/sl0uEWiTxHvTArl7d/tVZneYXNIzxr6qOt31dCitA6S18m/Tz
k5ntvQ1oGL43QMgp82FmT8D7dyUyO0jYNNx8aNm+phwpwJP0GOIqdBCyq03XTOhy9MH/9xAr3ol6
Tybxi68JqgP6tKkZy1Im5jU5gYJ9I2EOKn0w6zL10Pnpe40YVGeHTQQns4+IHbvmwvvsETbJVJwb
ITtdmqPt6naVAWi0kRfTTkz81n85dYv1AyDYoJ3YLHcnpzW+WzVDSM8dvU8nU57WGZNWvw2WEqQ/
LPuKA4MssaEw+vZJ87pS1IsAiSfYw/6xeRA1J8Gpumy/0YoKaJZYBju4sK50EPUeHazrvQjDE08G
ZZKGtON3XOcNFwAYPnpA5FuwMEzLAyguqWIRSG6SOWYFnL4MO4sS7Yk3G8PgJ/CHKMl/Sz6jvjH0
ACQdd7pKpqzxGQQDstcjpqd5JaNWHo32h/JSy/SS5NjQVK04DqbdpzesLGqJ318SnL5FOzR3fxTL
UZ8NHozkdT0TenpBNEGTCgmJVVCd7vpMuoanikK8W6I8HpO/FLqFeFVtU4h4fgxw65OyyRuAlt7W
YkxkZks5Wcihq0K71xC1cv00fptqy3+BoUIPIj9tjq70PFCff+yLBVuyZgR74qTDCHb+EygTLihC
MKwVO/a3sZV2pL6hDDIxcMeyDb/KUe9J1TQcqPvpQVjEnMjrCKE9Xdo/tCSNoa0OOozMTF/n4qnM
GDOfhGUbRiYtoOV2fSRYclzh+5REu+g62QFNOUpxjJa7Wjc+NZxT2vDgPU3g/SxN3bP950R9z3fl
iPiK4FZ/OMp13gdl8TN9hNoimP6b7eykDxzmdcDvbNTuKglAYjPR2SdV04zVMsTtIQZGF4Ap7M7F
HSfT5JpubMQlFmy34/4DQTpnnUTlwAn2a2gNcqG4lIcUltBqaEWwtip2F41eYPC8rNfbNylk1ehe
VYs0nYRbEwUNufBD7NGAcAJ1+NTmqMcL8WVoH2rx4TMU/y8lndH1gobdE2JTQIO9nyxhOgYb6KNU
5kOZZWdjmQ4i2Y2NrDy/1xU0kpZlNVqOLZe4pWFn9gVgYgcVBYfw7fhtYTqZiWi0mwztpklj+qZM
c6O1ngh1drKv0pPLREnCO4IVfvVdFyRez1e9zX1zXgXN2vDSkETXXxcXYJ064T/t70kWFOvLjUmu
ZQTywejS4VYhlHWbaTrz+sOC2MqVfAmbKf8WGrPfuJaMnPInqKYfW7tOQSeBQJaccEcd5heqqPKb
NV9hUOLikUKNxxw0xOM4nsD3DtgJyxSAtJCLwQFhwgqazoXbov6USJR8kAVuXCsKC+YUGWz3Bj+W
hXILz3TQvAIFK+UHEZy0uUF0ipHiW8h4KCZ8fetIsS+C3c+F+fD/bsGoeXm1WuDc6CrNq2dpdmHP
chCCHpbBl4WUxe6rJqwJGO8vrAax1fiMwwyCLTREzDkOWLtlre2f7IH5GB2L6cFc1NFvbZy33iT8
2usm6CnveIAOpqe6kLcVDSttkGZf5MwV5wpJLa1GXCDA0fas63Dy+vMZTGeeRcCOq3kMbsHkt8aj
+53vP7jOKV0nFdKaCkHuPm86mouj7OaFPLwMojk7/k6vbECpKwFEgp7yPchNbF+BiDV0gynwHvlO
3r0i4S+FEQLL8I01rfSM6I92cTO5v9xSPVMJ3AJvVk2COCZNvszVPcG4QJRQ/VS0nMHA6PRzK14F
AH+XOP8gDVjHa+F6Xz+iw4hVaY5XbDE6OUkuruoz8408I2zidmjmqyoyGV7X2d6Oz4HeVIoKztwm
Apj//Le6ELHaIY3NwVD6nqZ+IR+TNumLvtlZSDWpikm3jXzXbQCg0NJVsjX2eVfJ8GI6m0r9ESmO
ZiF35GNeuiYxc+pEmPrJS7iwRxTp54eS36sSg8ajV05rpOMFC79QuO5/YzK0S/Bf/m3IwzEVqkEQ
KXgia8QtXDlYxYQiFUDxhNaeoLmMQcJPP0MrRcxFhT48BRX5kPepxZRB+PKldVxH7OR28EU9E/ch
MbfKN0aVglYl4T/fxD10iX3TIU3i+hSpDeHCGQQuO1JM9q/QtoqcHmu0AvCBIyJ1+pAqrgIwOpfK
6ZsgxJ9DGYSlImMlf/DNchBu6Owalw6HegGgagJG2iuh0++7rK/dtZRx9zeuSoObbdJ+CMKLH43U
AxBJQrPTdxdUfKMwua9mcjX7U3KOENjTIHfRJIQX1PJ84Lgssu3RfM3UZ0lzIyS37pahgtiNJDmd
Y53vTJwsSnTTWvokhTU70B/bAtxoc3TthRGMUzCU0sW1Wa50coqyLWYKRtptpDhgV0mvZW11AA1e
eQqQVBUbSdPOwsBl45TZ8+CIbH1hYCW2azOYJWki5jdZNYh4fbpJrQWn3SYNMq4DDheg0U90feaP
6QYnL4K8Pe3vPGsmvXJeKKacitUa+ALH3a0onreUIGzehYxQaW28YLnlf3EnjMRN4UI+nTskkdco
qq+hyV6hZffCufKjHL0pfmlRPnveV37wJde0hLxVPplUhJxNjkuguFQQKm//zHRRi1+utpayW2j6
6zCmT2CP1bhCF5YgVXylONMOcuDL7J3AL4Mfk+w49KDnc7grma72VD1BjSrPwm62buOmXklwLoxQ
pS760N33QXZ447v0ZbbZYSSFXRWa9566gcbgqE0G9vmApfuXRVlGJGSQI1NgUne0g7lgUlSFvXK0
ZDKVOfmDM3oLOJHho4xMvPHGLnqMalmweZK8g787FrEiRE5lY+pvFsOkSs2wfWg6+rbKasCu1yDL
BkYVj2gq0K/XnfSlIxT3m7EjV3IK0gwIpKOZJ1iJfL4vsuw8DRQ8USymy7KW0VjNbHOGB9/ZMsvP
CPrcyQBBiit/N/joh0b0qUSkrqo825kQczC0o0Ho4tWJG/lZYhzCLY6LDmhamXH+l2KndzVisOTc
NLzwZlTs0Qw2aQByWf4Lh1ruW1OSD28wUFT9aXnR1IJFs5pdO4pMg06m6yW1VPGXjv8mIKV/HKg+
0vGRN8s23Uk0M1AKcWOsDXU6U1QMECjH2bnDq6mx/emJcJQjLq77RMwQBiLLbEAbzFP5Pib/nfpQ
0Gci3AhzUJ0o+mEyNli5cIzBhWcPPZsuqAEAM/Rp9TJrbqFtXGM4+pwmW5nQhaBhMZsTntcpwblB
Y5tkMQlmmWBFIBoFgFLXM0qnH5x+ZL1+k5QgsvN8v8Kcpb4FyOuOE9sJE1AwNQsU+IjaynIOLJEI
mVxSVX+xrmLC/bsj8HhthHdO9guvyKtlryQ/ASPds5mHd5X2gZjThZjzb8L5nxYmibH7pOmjAhc4
d3vE66TqGAkGUATeqhDjA0aMdIdvLnl8jpcBS1vZKOuvmo1YGSuM1nZ1r9a2bsH54r2OEgtcn3yj
sDJJ1+7Ns8DXD7HllFnsK8SiB6hKPJji3E14p3ZIQ0qXn2Iw0QedHmIkhnXG+IUPT2fJlr8ELa4y
2RRxPYadza67MXLSr/EZ0A6kAMH3w9sqhpxLXBLkw5UGPtva7dYY4rQ3xZWJ0uyglR+W9v+gSrDO
baXu3BWi+sIdywzTmV6DweNY3CnUQ1kDJfShtfx/AWb81foVf8rYq+tv1ZMOId2yaAwhpy6v7q1W
e47Nzj62ZithC5D9+lJBTPt3df1GG4AB2XiP0qiGnnY6LPQ7st2+wYgXH2iJTBa4sRgJhjiPlOKT
UUQo21v9iJFskDRK95T2jg+maORVqJStph20KjrbGud6R78ikYh5/F1oCVN+bMgUqofkxCKuF6rr
M/YvJoL+GEIQQrmlxp27rm8Yd5QscTky14PoGAobXdVej+z2nUZs8y//M+oYrWeaObUhPOv2TFu3
blLlCaotvCmm+RvtXJ3nQOluQTVqVlsdSInEX0Xu9cyEF7f0zCCaz8IQEJ0GTprLgOJ/vBS6Hpzn
0I9BwVsenUYTl3h7z+Qme8uJ45vf5l2RBjMs7FzsyLpS9RWWwqhBK/ylY6OPMBbBhSHzota5AcmR
pVj4rAeEFBfTEqGfR94djopy5NXXd5vpJUWIZ3Ww9xAL9sap+DlAU4wRHzpg1EeeyMQi9btKNkHv
qtLWhFNZHGyjED9DO35mMcRTmLom7pgSj+UwLX6R6Ybkudk0duFY0/SWhbKkMQoURYWGu7OPFQ0d
cxzrSmSQKD4zVrB1GKkbotVhzoHxUW7I6TFai9ylnNaw/2dmkdfZo4iEsGLiBCQieYShh5SCvORb
R3il93c0xp96Je0156kNyVcEHUuV0T3dmFRW6xrcZznC8Bb7TCTXNFTSQZ4z7enPH0B2G/h8lQVR
YruICurR6FF7mLB9dBDqQIPJATmJkrHscFmMYE6fXf46rzcUyYwQy5upHrKCQ7lHvkMZHrJy4/6t
gGEO5uWYpnFMzOE+EwmYAZhZahXMGW4BmnEMz7B+HvYbvGCTrT4PeqsAcQKDVEX80tb4o8dWteUD
O11NDwYG/LyFeIbwHDm2F5na0rULdBw+V6zMYmk2MFClYG2MlK1dU0S9Y8eVv4yDIua8Qn4I5d7A
k4dD4GLe3jROE5gHpVPdw3Th/l3bYegeHl29jWT43fjtbOfUTrdRGQgq2Wa5BL5/XBr+eD64h9DQ
7mXyDCvlwYA4Ncoo/edgSLoJBWBCKLwgryKgzkQdv07Ghc+aBOaD7eBOWg6xiALw9ecdPmC3Jw7b
xBv/lyi+e6W/Cy/DFSnD9wM3jqumzzFmxKOBFTZpfhhemlBVewOEQe80ZEjT3/RCoNrbRZz1LGhe
h9+UC5riqaeSGqfNAOiuJ4tLjAifP6q/3QtlpQjQNuOkRj5j/gF8JNR/RsTyFD/fsyPWTOaOXF9g
ZWcEOIEVKvW2FP6lH70zXEja44IIBrAmoRWMWzOFuOLkfxX66yCq6TCyQUkxY3PxwXIGqUx6CuJD
YlBTZG8t+Rc4VOwWzfz4m7GRyKYVtvpfL8fjuldmHEGDk5GwId5QXlOqnTwyZCGMP8d/CdJkAHP1
FBjV0FFq7aNj45iO/JLsd959ytsp7dllEJ4HQ2sD+IWXXDQWHjbPJa2cMNbxrJ4yPCPXWKVF3HBb
+LuTk9P7jjSpEyCiwlWXBXvxt7reGv1iDBJPTrGXpgPkRNn30tvAfMMjyfC0Sxycz82UzLT14b50
aVCpRWuYf10s2YqrmF9xa9ylWG009ds73/HWzdvlsk+OuWn3zOtaMQA/6UvZRKB5PlkWFLQXbAAg
BWkHyTZwcT+qPs1YZEfrOCRPX8lYiQYAW4S2d8HM/JbSr3vQc5ksytOluihy+GlmwseDvxTPrUOJ
OuJi8KJ6taSeCHMwFBzsiOPlCIxj6A4uATImf2x0IpwoZ85zaruou69NUuFxaFagRTMgd1b+MEYd
N9F/5se05X/wq1i7Tbf4IP57F84/53DsBGUzAMoPdE1DnnG9pffJLakAAIBx5UkYoLj4OANDlVgW
9INfTrfVV9xW0j7ueym2Z0FyvF+OsGcqS5CV1Lo5x2uv1SkN31lEbzsd0mZm/OoQCdWIoDgmsxex
kErqq04wbczaRHHDDCB1S6NhyBXgWEdV1NHScu+3t5W1trOolVasMZEGiIB5PH+qqCcrii53Mp5U
KOpNpnJuCoDlUcOtVNgZFIhNfEtcMDRl6iZo1DFhtFA5ZyDyLPfImdXJmysC7dL5VXb7+a6yxx4F
/zNHRnos1UgX2gEhnkQ8RaRVJ03S2J6c48J6OTkdK+c/B2pINKVHkQ1WmxrU2P03BTVZQS4So5s2
auMPUastHIreLK4hVR0xfS5w8aPTfRcegt58RzppboeCwnn+LqeFBvxH5MOG1WsnXRcwOqWvsfhD
QiMVHt9z7LaBSLgHeiTh8P4vIWOvq7ebJJuirm6XJ5Zm5BZS8vge0hvlVlbQkwdiDTcOeUcuTIRP
4jXLNPtDVvZ9fDkarvUdM/pXYQyHbYWZTX4MhmZXeOh0HB9PRlJC1I5fhALIbrGYgSI5n51K25Qg
Q9YNNJgbNZpTYcI/keiJ2u22Uk9s4xDOxHOIaMzexTQIiwJ4507/lA/5dWJ86rCMu4hat8u9/N3b
MGWBsLCA+FwATnWhwH8CWQkFSjK87+oYLRIxlyslTwIH9++iFKhR5F32sy49Yg1p6uCvHOmjSp5W
LS6aVPVS4iC1LS7OWLKtZyubbIK/CjcNrhcds8D4I+ZyJKYZ6uDdmgiXGnH5mOBdHVJn8WHL+AiL
RtoNPySjeLHRb9qG59FHxm5cfrIwv58enTGya8SqWoTEjnJz2+QB3FbC+O7FHdLWpgdQq9gD0ieS
BuE7cYpnJks9/AfHVwAySPaSGUKZm72rGpq3q/URALTkf8nU/h8/lHZpUtg3y1TS5lpIkbJt8gEE
ErscsSuLQPYBYHo9yd6DjejhfedU4XU5ZmWuO9ZQscHTp53CK8zVn+4rMyuB8P2R8+YSHqHZ8Gaf
5pkns5LX3gS0ivnXKQDfJZ0itHmWjPCulK1kPOpiK2Q4aMKKyU3Yco/mPCl6BuKZs4BQuzmXpYFw
XToKjCtT6hKOiNLDGjJenmAXZJmro/mR0dlXGN2tz2lDqQkSB0sJUD68cI3rRt2RLhgK6U4Jn8zL
6cabwdWM1OpiFoO8MK81nZFb7mcbHoWKVRU3mhqYq7nDs2OaiGMVmVlk6FlTYTnSHzKV7mq31u4q
rl3IKF/qwSz9HBPOnbnLP1ZWtqDvyEo/44h5IHuTD0sRZ7XA7P1QFwzNWP5aMj/7zbE6kwG29P98
3noLO6ODFcqaZI0AiifcB+cBBJG8nw+jJRO6eF8ILjxzdZDH/3+497lqYzBrAKWTCqIJfBhndRSU
59TqfX06gJGfkf+LwgqBW/tsWKeqhZHGZLvdTm0bi8CDRxBgcwnMClOw5kmfScEcEDmJKzS73b3H
XdJx5bkFBd6IlI5egfWbW1kVSJa4ijcAVbbYLLcOhz70hiGTwaFuLTbA0kPEFs+FNbovF7xcNOJh
K9eP5joHF6/ZXJ6AgyZJlh0iV+7WUf0iZbErw5cvJ3IA18dI1hmPbpruxN5sTE5P8EGlJ0nzcepS
lDfYNeqovXNhIBvALFGyQPJ6zAHBGUhMxDnuVvSLLZD+OIf5P+AO3QFmsh6da9INbmEP0xL+mwfI
HsMCOkx0SGsWU+M6S7aYFESaUj/Gh3dpYanwvCPjvJ0ouHqokY2ugxB3eR2jHimNyHt84N/XHES/
fqgLGLm79dNUDuw4FNRMv++4HLPWnFkb7u0HNcs9wJ6DWq6WCmoKQB692SedN9BnxMGW4EN0r15r
FMMx8ajqTtt7pLHctPYhHT9B7T87awHYWuajcKqQSKINSD0tuMRTcLl77IYHuvtll7q//ct+yIkp
PUnuxgPKEuwZyhKnjdc21GgDAaub44TW2GeKk2tLg1mmC7DoErg7saCWpr8ALVuzOgcA4ESTVG58
P1F/aloO8LmNlJv4JQNVSWl+B6dwJiLC5JbVYYD4lm1X8cWQ4hkBHGlLU1QcL0iz9Fp0iLvBPuom
xioe9Xg6Far3AmUcB3euc9UFg8Xd54wJamG+1MEscoczA067ifuo+QHJyrEDgR4ymZ3N/ARnBJ0o
qnAj8c3GUwdfWuOvvMPvM7mx5H9riQWOGg35ftIXz3V7IyiVYvm2o2CMwEpc6EH3yB0pD+pXFzVe
LnIcPmJFdyjVT6ozwxph61T8bocM4wkfKJEgpboOhIFEcDu9w9gSPcB0G0/oFZ+WakPDklxTDcKR
vU0/fUxVRineUGlATTLUILV3TsNeGlfwVJ+XVYKFyp8RKU5+Y8S7BhDvpB7/A46pAPu9I+0K5aNE
f92Eee9euO8M2W7/pU1SrEm/YoCBeOC7g5NITNTwHW6vAmkvqD3UhcsGQlSy/ibfap1sCO1oU1CU
3GDvOXPcNx4N6sxcx7Yuur0GJnzpErf9Q1c0SczJf/ITiMB7uBN2zfJ7MD5PEjwNMfBm3uewN6e4
ilAxno6CuR1UilNx31LAt2ZyO8yY0qMmtvL4kdecKuDhplxnlBIu9eBCrMjfX1FbEhL4m/jzsaeh
eort1bIpP4ylQGTtaa3kuGjJJN2j1k5vMrzpCsgCDBM19GKWkp/OkFsQ1VMYslPeVLYdJtU8wGwI
8rXbySPPLSjv8xFKaZsX4ICpQUXm3K2cuxEeuNw4gKuTTDhPPWmZejkZZls2aOk+DsgN0LN8vjiy
ZjTlU+hX57nWWTuTY3fPtp9E1b7Hw9TON/NYQfeCH9MkCZYjOG64Rde9jHF/HOz+Fy+xbaRVBPgJ
IeDPbC3IEISkgj8RUzzofEZFYuewi4rf3SzRBN7IJSvcr9i3MocGS1JtEoLN8qC4pvVsBkYXaQWP
zYQeyBEgt2shlTD5yp5soHPE5wkRSDWI1JmHboRTK3muaa3OLeV7Kro8w2hJbWJ79uMZ16GTNfWo
2p7FWV0sQ+wFJ9bqx7o8bh30MUqM6H+/seJ4MYLsIQJS00SsGh3hYd8rH3i+kGBZU3HGpSIICf/G
odENiv6G+i4WlgmJAWErfSKVQccnvkm/uv9cYDn6EtidGTa69HgrBhjatN1glTdWn21NorQgeJ1s
Kmxx4XZ+s59pyt30xFfeHpsZjcuMDcT4vt5PvcpBdLmrBALH++Au9cWhG4TIFx2EbI2wUcvy61XE
LmkE1tVZOk2IzxQv749dWXQR0PsQVg5/MuQ0EG49JnNzf56yoIb0PoIqnUlr+RweUSkm9pEqu8a+
auplVhFruUYiIMe6Us4rPIfpWNsDpO+vUwkz5NEDvLApCqGYwsGIrLrZZA0Z8LBOR98aeMJNlRb4
VEbNixMTsWghEC+f5SityrF0lIC+D8+eQO9GS276zRqiq+0+J2CiuxjUhbrftIqWBnyeIcZUHjkV
uoi/S4k3vgo6erqJFjNRypbrImCPD7PWxhvSi91TZmLCrEAF7uFxT5dzbCTlbZFoh5vva6+kPikO
cfDPp4RrArusfpIznfxJmriZxzoRAvQGRu8i4J2GczuhOnqOwVNqGdX893RK13ZRRq4c7n8Y7+fh
byheHJRuhYLMYLVJzDcp0xC5EDQ86nsy9k7W7QAF3ZjNAAAQsnD0XjcI5Fw72/90QMV9AMBnY6JS
XvpyU0ExYdEsUgAufccUlFhcrf3OWpsYBukSRh4RROMy5q2HAkHSx5FmGtdQAn/5Uy7AoGGC/2Ag
3754myJuSFKOfzG5OWYwFcsqWap1lgidXu0NNvIM/WnuqSloFoodip0d04W+IcnSRKZ5a982Ihqp
YdgMbaXCQD9Pc7sVXtKTI2tNr5yQuaoknsxijK6FK1Re4a3BoNES3pNopWnWP7F2GklHCMQHp9RF
dqxoGdQHPH/7nbpLEv5jWh9jtKo/j+V2Nv2/cKDJjHNJ/02zfXITbcxkhMIoZPMTl0bhdJPCyzQU
K3fFskdPCD1Ko3O6P2EhhnkZ58yNh/yWWei4Q0z1ggEO4H+fbewq4D9bSOVVG+ykfzLdtIdNrde9
n6OFZZDe2sGWyFdfD9cAj/TmzFStnxuElUOQ/PlPfbBvpJ1OOHtduQUtq8FqOX/PUM96iKvYrPvM
sA3Xq5yC2+fruofp3D67hMsXzC8oUIP+R2C4EW1jc/N/IZsh88/matNZ9DmQaAuT6xIwf5g8dKad
cihoC1Yi/CqF+SdlUnwGSKrPrzOjgZ3X7OFCXpP9tPGAyJuDg5KB4uGvQ2OD5LVPQ+g6EO9PjqNL
OPsTYsgeVIyhrMrxUpPsdUsJS6+XHWHUGuzcSxUED28X3t3koecs7PVtIO+fOWNKSPRZrp12prs4
HNbhLtZtSrn7PeFGpsPydaDcht1LAnFaF9y0cUpsZYsg/7kkzJXxQ4gET1+nyq+TQUTrPeA9xPDF
jsuB0TI2NTXU5MswuEHMaR8ZKIb7+yH/xlZ2Fr9q90yyA7dgqTPB1DgVso+1JX1UO3K8ZECVMlbP
amttzjE5+Z5JYOrVMxCnuoRPdQqpV2QBGzMs80UUlbpcHu26X8AAEGWDcjsrgKrG0WxH3IaVeZ5n
f41KyjEMlTE4xhEMJRnVdQtf42ZI2O7yHO4JsGgt8Rclu5iYHwq3BsGE4YKM9qoYK6EfhKjxLOv4
y6YjsANvoZSOTqqJ3pvTscmU6gFKjRQX+cHWcaEM5WCAVKx3yuai1SgrBN1/77TPhvOkwQx66+8q
pY3dfsIg19pE9uPx67fK52Gp7w5OMhDJTdgigB4KRKL32dE5LcpBQa+k7QsgkwE2Jx9Jx4e2jNzk
cV+R8XC6dSaG2eMNyOxORjEaPzcusKuszYYEocc1Fe/KBAN47MwnmwqTcTVTA2YpKLDBI2TM3P7l
RvK1l6z93JIkWh4sw4yG5eZ19QQYdYVPESp0KMmnq/sarXltTnlciBIVJWwNKjHjxGz12wvJCmRF
M4Nka21NDTfOK7z4mrSpmHRtJZUP2HQXVYR2SaqxBsc1yunYDfd8mjppt95kaQQa0dRBsfg0nVHu
uhM1SEzslEnShN8WNhQyjTa6PYrytppcIWVo1DQnzcHmIOTESuB4TTQlB3Cfzw6Ts7ioLCO322E6
DgwYlB/OvrODB5DWaVGQ/eCQD6C17xSlgF+U9xkYX8ImdN1Z1mN9wn1ao208iYKpMphmjEbcqI9r
v2r1OCR0YixcGVWF+XQbvOV22ighDBmdoLSVvw/gqLrNkqqZ9qgBEwoxLnvOdc2ESBmeWm7M9D7p
lTkB46wSMb/TwHAK5MI80tqwZ9jFSrQZl4pDNmQQrfD8aiMIH7iID2dpMA/LpSgP44PAPafJT/uf
Gn7Cum4XJk8ZpvZTN06nskxqUdcoKQGY5vqNx4NkU8vKP9IOXnlNOkGFNqvz4VxL6eDp8RcmzmS5
tK9i1e9H+LKPnJ1Hb/EgHBmfwrDZUB0Hth+5x/kaQU6EoKO/H336604roSGldPMegAdSXDjFUI7m
/3YhtPJKcff6DDKcjwWeIHjmXHma4Y7oDEptEDS6VsJUrTuDZ1JbEjyOfFAyq/aFGxaIyni4+gP4
TW5fKQPP4U/JeuOfALrmoKnFUAQ9vP/Rs4qtJL6UgpQGqbta62RF5SHcC1ZgwQ6apM9JoClMYTTH
zv5ZN7UdDCcudxFUkz1rGNin3ufJF+2kpNZxMFZTmivcLwXSoVGod6tCoekiRStXI9+Yz5stsNyk
zsu0etX6yLx534gV5nPLQJafIqgjswPSj3HCXjatVrMK3ND2yfiaSMhIyytOBwizmyRcCEj1u0V1
jUOGomW8wEvkPYeBbhHq439B2MeKSlFuIioMwtvNMfBvwmsDbfJtwKoLgWfPHPsDBdop76VjBpdv
YLQZ2FrihIPCDH0n1fkswCa5qY+5BWyp+0uaMSkWKqFEaPFVHblZa9o49U17r9os5vd5hqe9sAAL
7b934lXevXKjrvHPXLlfcwsF5NelZIzL1P+47D3Ysh8jcnU2FvWJeQteFOeFs3d29p0PXzMGYaXv
UZE9uk71sYBHvc/VXMnlASa7i/IhvLeSeb64BeFwk5WEtQzjWjZw0dGbG9bmVXyyVTmS66S4Hkma
Kx0OeXSw1rD5QIWi7vCcS0arXMus8wWugOYvkxFQVind+id8hTfW5Sx/EC3fV7uv/zQViJA7Mvj9
P+JJp2vkH8IqY0fAujlQfQNJ7V/W40wC0bzH2fCwozttqJpoPKPulMf8/vZp/mE7B6DHcECX79Xx
q8jiKHknaZp9MWlihKisnQq65mrta5uAI8csmekJmYepjmLaYIlki2DfNMy891Uu5D99IhQFqcaq
4niWdI+JAxPRnUWZZ4eH0GH2u4nY95Dc79P2jRYcUMj0ibnMXskWzu9TmIHJhc1sn1o7/G9habK3
KT9D82AixRYqyYixKMcfyAH4U9RujG/rE2mjqp9VWWA4e1+kP/aH9glSiNi5HnPM/2Lo1eovH0nl
WiUWnYYxlTTB7ux9Ib8eBws1KBxLyTdKZWVjQhLuYEzm7jVFn+GZ85AxS7wpKhH8wgNOkc3pQVuX
nm9KzB6rcNebWjTru1NrWz+w3htjra/xjjRqf6L/zI+ZVsdtYXAo8+jYMTZMfiWDK2CezobSa+NR
cobVwJ9b0YooMesosyAXKqwNW6NjSOXpOkXJln331gB1KZPfYswRkBt3LFDk+vm0jsmF+0aCq/S4
lUjI+t2vtBJvMf80JUgm+P8O13gbw8WGCFWm88zFakBVoSlDsTCFPywj1V8m8S3P083Emw7oo5jv
FQCUYu1Zg3vWEHgegj3yxGrAzLfsKdpdZYyl5waozVs458W+Hlf1U/TGgVwA9ruTjAymDUCzlEGU
nHfrjJMkSFikPkpuAGLBvNpaQmCudXkG6I8zPkiZxXfKSm6FVyyc/oGTGrAltOitgR4CyfQmC9BC
7i6UfMbxudaNdGQfEdEtrH2gU45cRZR7scx9y33U/6JSqSf7mGesVHNr1y+pL3gWlyTXtgqmvc2K
VLbtALKm6rX42XiJDwRe/mreRvoAkoTN3K8p3A5UKn5sTbSoNwmK5BpET8Q0YgZe1OJ9wncJuurP
dBeOFXE2z1l3NcJTPF1evzfeC6GKkojUAyfPMQLipzcv80XhM1FYCZFU6I83kDmUCf3RT3kP4eGo
gvdzfgqZOR4oyKVBtneTCUbzL9OxnNJEtpQ8yYh8clsqFhRA1mfxxlmmcxUuDgvSWhu58kbUJqNX
bxYMFvMhyniy2LS1loRhz2NiXJZekA+3J+LwJrf7rWc4Y77RWTPPIZv7kEyLNz5WXVsmRydCLwAm
pAlUGC4sDc6anrd3DLsYJPyf5eHK1HFzMDmK1KJGVqKu4dltlthEwNGFDOzUPGOrHZUAz/2/9bfk
hnGmEpfVqE9I2xenM5OO39KTkRopADBO1iD1KoxMI8B/jANyB3yv2RKDeC2Jy4HZ6LeweC9nxV6G
MvUmpd+L0awfrqmOECTqyLF7h4EXv2WRSfm0a7thZZqjfmty6HVNkev67pP8zt0fb+EeUa776tTG
Lam7WOceuwvYB5RVImZcE3MHkXz7gmveiSDdckGdStZOyyNewANRClqopLxIj3dTnug2CvryO6SB
kkY6ENyNtI1cu7Jpx9ZFhe1gLot0fXzSOoyG8Nqdau6IwJUP0vVGswS+eeOFIZhoIWhoY3LuoUGR
KArot9CVz5jdJqnwrWsq563Ef7JzcY5g9ergS4H3RNzHgY6f0HjUDMZQBBNDh7sX5xanlfVqCuqx
M2usKc3AC5ON7a+t/MgtstL29GadEMyCnM2ONHPHuOmy8urT0Iwzo9mITlxRbVo6Fdmo3XagCc5a
aWKQeG+/wlFGXAQz4oZ/Ht5nkxKZRO61x/OE6sk0vVCnelArGW9Y3CmToSQPzZXhYkP++e8DmB1n
PgBK0+l0tU/3LxkavvbzyH12XoOC+qGbeCn/vGMpVHdg+YlglqViUKI9ufljMKbR5yErM7SdiBZm
akiG3a9JBAedp85B7UFsNsiHUktcElBlvtQx27x1ogOi5OmzBTc8rb6zeUH6iWu16lZTWZK0sEm7
aRD4gmHlWMyZ7JcF6gnztNLHd7Y/udpU2Yl5+tvrAQYLifZxqXC9kSyvWzTad3gLqQmAF8CKK80W
vWvRjuRa3erWcZzuFjFab9uiTTHPxrb/TpR6ze9fileFuSZVqFJyzGE2TaNOt2EL6Ll/8VKXSdiB
tmWxGE8MCm5K74bHRIic6xuXGwfbFM0g79EsXYIj1scpW2pAnAn+vrYUXKLvg83kEjHnwhCVSt1A
RIf5+T5tYyv4+Mg02HH1S2gPUvaVrcYRrQ+7CvpnglrHy+gXP7S/HShxss0Yqskx7Sul/9I95MPW
Cs4jbvmygulHxyW+tWxxL9tEGYd9C4jGU6ge5m37T+njwMIf2x9uy3M1OcAD0yLFnniHmH64GxEL
QnLAsj0ZgCgXL7yCHR+tDgiTBE5VccdfwVkUjfoC0ZBL2MAKEpZZQHmi5CJ/bB4W/LBK8AmsktHW
CykZYVtWApK0Wfw/6tCB/xruMrFcx7G1FqAsttjjYH/6sU1lzMmoIOslNUA/cTcht+4IzjlCKe83
J8m81Jp8uUCMcc+GDPm826WyhM/cnKp2pg6SREN3GgtU/LGPN5muzXbI+zYlOHblyUJQAk1vormF
ZTfbaASdJrUv8hFIAQKsI5haBdK97FTKXzuF8LhAKV4Es5cl15B22koiwZxLZGEEpcLFGWbYfaIx
UPKC58sl1QEiot3Hb85wGdN+CFlNsDzTJzWljjsqv40N72R2cXG7VJoHGcr7lJDdJdTXXZbncqF/
RqWHacjxRHMB6cl6OwXCNNcovuHdzxpDiJimL3F93BrZMbM0X5vpXZfEd5m4fsg6AmV/WPxV3Czw
WhfDkDBZth27WhFkfMfcXb+RqwQmtlw2o5d1uN83rya281ODqLrjY2AER67ahtwxrskDK7cEnyWI
0k8Q8Hvx1tV0cSOXDz1mBOdtZcMPmO5k78mT5JyNHikS2nTdGiQMama09ChuGaeLYtNVSzNL7mZ+
oXaPG2QjQ9DqhN7Gl9k8ywBGrxEnrWtBF7tyuxA87q3jCjKo0ihwKQR+LErOVhAc2bDuWoDj+mkr
cK0Rd8HrbbOALlFg1OOAL/RaE7dyShG/GDr3PyyAaQsdS3c2NfbS+QYV0Du2E+PVV29jmdQZMVvU
j6LR8PHJMoE4rje6QOo3UN8giX0bG7iy6131c7lOHDUuGB8h46H+PzDpRJeDsO27RkEKiuVi7CLv
Kh6Nz77F2b7jSPVRxR42tDekfzBj62aI1plxeqXNSPUEX6uos5Krg0ITaetaPfWfC/ShrIZ30rNh
hwL6I2iiHUTBiHP15IWK7S3lur7MCk2VzxiZvhpmSpFKnewFq1cLdSDNuA2L92xFMbU6NVQJSCPd
jdJrPagtR0eM4EY5wmLsx3v6o9LNm1qe6y0h/AZr4qDqOzmQNPUPAcoHXF5M+qrOu6/P6emF8Xb1
QOpuaODRBCoizmKWkMpLb5HF9/3VGl4YzO4aCKW4g4pCYCb0OW7wL2gzfT3rKjif1HHTx2n9zyEs
ZaVWaeTjfq2jMftxUCsqucg5UI9WTbFLuWR0SpHI+bxvrA/tbaysmAdTsmJ0mIFiFRu/lXdrdQIt
xaSoVIinh+odOYEK0taYl8AN809d8/n4a89tym+r9R7gUeXvBJBPGLA6rM+gpl4I5jPF7IsfbmEL
3o/N+ruCODRvZQFiHrhWkZCohYbGzRwHwCWI4Q+6qYJFRIRRIkuOi35P2AeepwB3ONZ6GNi0PdBq
aZVz5CA/GTYCFIkdmU8PGgQeIC5qcT0O3En+7jaQhzy7lpngm5nciA/oXPA3vxWlkJurQ2piGQex
L0ER654VzayOXV2DQMWZiUe+0C1A8JSWcqfdPTlC+xMeqZyJ5pOhI5Z9Ad3mAmnW+YqA3q/vWXmc
zAGc45HYBm210XkFaiFNPOR21eLrm9tBVASlefERjKD7kIXyY9sEDqbCuHkMDSn4goe5GpeYdf9r
GU/VA+76q09tKjB+r90yq387B2sGUXhfVTByB7b5CmhYHPxRf/pS4rIyw8mo1344OI0xTwKc5Rwp
kaokifl9zpfU2CvD4/MJiXmdFBdFArT7KZNu7rt62IHVhSbIjA6ToPANjuzsbSWevXchFKEae/0G
1m0Y+097X/5qhyeMf8FITLNR0o7vWm/f7jYirVHdCoeSgj0C4C6FTtMe8EqurYT3HG/XY4LyavyK
HW7/UYTiaF1/7NIqDfvKNBfANQNaV6fBuuVJ7uE367K6MXpun0puug310ICFfZUaAvc49a0AOaJt
PBFP1DktnmBjVq3ySVWK16VrdD9gwYwVmEnWXkbCRkBKNnxrsmEtV0a14rVPkmIbTVrtAJmOhn4z
IRoVibbMGr1s5rBkRwhRuKJs1rULv0esLw4fHThz4okJxD8X2ypI8VeTwwsDwAPNshJNOOjUn8da
ZXEi1rsX3DciCMWbE6aKn4/2DxhMKcEZy20tgTHjD0/ghQJIFe1IxI7anpmK92JYdDwYnewZ2OZI
e//H4BXVgPyT68QT6TBTnio2s2tYjpGoBHbxWyA1t7pgSTlHDrpvHRH9dJ/KvFI1k78mdWAYHXSu
0DCiibcX8/5n4KQGtoph5GDArGqVl4PxjdvKYfpqXetkTNjxs3dhPc6k9RKpGBIGhSpp+ppQzohp
2yAov+e54eo+JbNxryVJMSAymnaEd3xJKkvfdOvyDoV26PW+9kcoB/GUwdZaTbBkj1NwjP6lhK2p
GykivAomBvHJATo7vo1WPADIOQ2lX9RLZAdpdYOks8dlkJ9JQgj9Px9O3ku6Qkny4OQYrWjjTgPx
126G/d9wq7xCJzsxhLU3OFxo9hR3TlTBwKmMN8KFbgEsom8N2Be0XIkTeV3ixdKJxDoJQ1sJNKQ4
n3EY37whAhW35v5EepCbki9LCrMTAbtPP93OR+CfsVwxwXXo5HnrcQXUOspvS8VAcB8uSmnzx3eL
8kVFWwFe83o3Fo68K5LI2hp22rShWrd0Xb7s8oH5s1giBQ6fDSUgJ4tWzu5elLHi7JreZrofphh7
7A8GOYMIxddS/sOyY9/dsiT+f16BfR8QmUuHdvslYXTA29ypn0lkZsz0y31QlW89I/DoFhLTlAIT
P4wKR3vZdFeu4NDxRBasCN9J2aB3lOh3FQX76nQKSfCe4F5+Lc9HbYXrrTFjkQVDq2qYn0jhf10+
GEGI4EtZQxf77jdHrE/giM7pkiebcDoBzq1uHPgRvaCWlUmyYlPrLP561PWkoyM6wUOLxf9tnPt4
a36X2wuDRdeZ5/0qrkWiEjJKdV4D8Y0cfIPt1+K1ndMlCy6Y8dCsExTOfjmH57FmKHOI4g0ntAP/
AwXlAy7jvQt6DuuH1qhlL8ZFAFS0u0N4OD7bY2WgZsy2c4CI5StRiKxMn6K3+Ika45jcDW57OFI3
+TUekGJ3kpwJy0Pl4hlRWvaavhnMgwAqESHUdx3VkR6umnsCFjm5eAHz+FAaacl1Gc/HPWa8sRIk
Fcv/ew3tTyKwlz+OX5rVE/fCy0xtNKvIDR4Ef+S71ljHyUcuvFM70A1jU/ELj/m9KHqsAgMU/x+h
vtcjl8alrRRYBH1CtCFGbDKNvL0dcLkBll4I25+P2SSeOiyFR5nf+6WCgm5xBUoSi2oQTohmHd8M
ZwIlHitGNgQSXDrfrYxMDRacqkgbbSzG1Q2pphzeqH9a8OpZ/CCQC7PG2NicPUEdWxKeQNOv24XY
2Gzo2e3XerUMIwxwOV25PkE9ElclYPDIO2zhiB4tZGuIlR/qwWwZrDEmgyJ0KlZx1/Hep5nQWOlP
/aGXNT0YhOQuGd5pzKKTiZWjntIiI2n0WjnFfM1SNRr9y4fd7OrOp3ryrVayeiBYRts18/Hy+Z5d
ZcdeXgGhvWhSifCRRDDveg9WSkyyWbaxE3nLKv0z9r4I7VqbaNZvuyVmLwrPrNXknuUQT8VgUE+y
q5wv3T3DPlP1IGGa8janGdTOWsPZ9FicKxGafJ01DxILQ4iXk3K0vL6bsvho6Jm3l40fJYMszeTC
UoaXSg32HAg8YomXbgySx1+MwirI62N6hvMpDng1yFpsxaPaICEg3PkeynVwwoFgfci2Oauk7Xj1
EARfZxBXAmFIZ7qCnOKFDpvaTvG4u6+gK98qrTlaKQaP9t7IPbq/cDuz42CHWzkF5O8dQZlOK3nR
waB1zCUdIXLAiGphIb6RjVLmsHV70jf0VUovkXJTeqRrbUrVer2VY0N5DXQdZA/wSLF09fdftvL7
Wj/AIdF6HuDSYZmuTWc/ac6/jpb0h70LxWlBK4s1yKCkWz2lfD88xr46BlxBBnMSLqTCfKlPT1cw
QM4TraAoL8NU3ghRW8mNrOSaFGzDIBlXrbDk5Ezjy1zqFzjG19SDVTKZ9i4t27mbJ7wetuxeRAH7
OT39vDHZub93DDNlAQ/om1CXJ/fG8U3BPf1qHWRwLlMQWdTRxrGk3OVHwMPN2tQuKaOFHTLr9TEs
BIJbEhXSbn9w+Q4vAoCqClG/E12qp13xRuzfyF3UYxw94w1zWK60Kkbd7ScIMGgapMCnv310/IEA
6N+fSeuRenseu87Zl8YRG9T5gK+akjEgJ36Lr6i+x5YNz0yi/igTk8aD+81gjCcuFAMiRFO6Z7v5
l4xQRnYstdpsXSXCKZSFtrojNcQLhPmhy9U3Rri3O2V5fo2aLRiHDMsa3MbIndGYFzWpzVfXotmj
5Ooo/nwKp1f4tqiAfar3IIt/0Pgq5XZuc2zgoE68G7IF2y4sLuI1KmU3iTNSuj3XU0ObCj/EKoZS
8KLNaxqTM3kJs1cecgw0oSWwnffKBpcGcFsKQ8W1Mp52qiZxAzUITGRIhzvUE+VZXn0TAbN1B2AH
1f+zkRpA+OXCW3pCorq/Zby8qrml3o0cOA8Z7CbrOKzErZv+T5l4gFC/YKPeiK4gmRoA/U+eUph2
9Cx69H5joiOQWbn+HcQgq4URbxmjk7PAHoBM/ekV1B6fhpzl2X2FXoJU2M5VFDIv8XKWchksNlQp
53IKojho3nN6gtIb3qi01aLBk/95QYVrntBKPErEOtmIvyFOs0M3pXIr1jJQ9X8ML9y91+wzMQr9
1QDiCnG9XTttjAIgQpcea9WVwk5A1lzR8NudbF7ut+N+VVGRPERVbsstFSpZazYAl9dmYANrdZtJ
0R2eMDsinSwzx+IA1S334HyWdqBEyRG/iQ1rJ8aovCY8gQZEq5StcttbOri0JClGwJUZ5GFDP0j3
RqIIl40jpYrjsnyFx1N+FKm2XkD+TBiWs0RK09if3eE1kw/vKQiVykb24o5ljjgkGGfMUHrMntBd
XMj0e7PU/D3xrldoRSWq2IhTyry+Wr5mrAFrtpXx7OWnfUTSTOxcX8OX4qWCjpSRKjcd2STzlECZ
fq4gXEUnc514sYhtBvMGhNhmkMhbObu1uCZQL+u+2DiQeFR3l1I7TX74PBIl2or9l7ndRISVb3v3
iHT07degBt4rQYJSpGgBqqxCx88/XTUxDr4tF24PSU+dd7nI/C5jyA7h3tbaLsTPOPHqkclNkBXz
hqksJZHwOJ53nGf4CbEmqCsFzyY4s/5W2oyK0cEvEReAQG/3yrkgaRW4WBGJdZMftsOR+EYpvuJC
uReKjGPAQ9vH4RhaXaUPSbSCrsqdoGaw8qR2sAhehQBQEWOq0sWwNMfnP2khuoI8GJZ6N0xHlDvY
Z/ogWIf/SVq9ZiNrja0vW+w49N+vwBMe8zmFaZv9XCHFQHAKtxyt7FmVf2lAANUoD5owORc8zQfT
ELKSi1oqQBaaYMbYi8TblqOFQfB4RKTLEmpH5jagzWUKoM+tUhcWdoySvVE91Pqp/2E7ophN7/mU
5X9GwFll0DQPQd+XZCptXU4JJmXrFVIlu34RlfvZxLhsTMqB+FH+3Sky9e4DFNkJqcc1yFtsIgaw
2XBweGKfe8l3V2hXC6B+7pPZ3TnCkmE/DESroFyyWElim+bfeJssHFnRkD7iQsq7GhU96G2jnIWo
qTrU4NH/06Y90KrLBxms///A42VuhO1E8cXoFrf7Jc1/6GBms1EgVQy9lduGB2uZpK13fxUBw7xc
FSu8PWMLqbfoZisGnuaRmTCj+3HKn4Zi2lLToBKDUaz34E43+r3SERQqdpRSBD+NKJfqqidZT9cZ
YVV0g1zFTqDKbieMogYY0yDAeXBBy5JAHS9GdvAh1t/v3gEW840xHct80lpuUOFs0CP6irNVur0/
2tbz12qI/1Cu+VThRqA8Xy01zYu3tGp6+nmYedBSCULNA3WsnN0xA5MYTL27XRRoO/RuEA7nGVJj
znQXxej5PXMVfew95Zzfo6NoskjMK77vz+JoQlEoPO07WriA4W3DhijgJb/kAZGDQfAltpFIU7Fn
V25ZA3sWTfzyUnkclHKp+AoiI7Y2Y6xl17xfVjT9WV3M64UA6AUHoGZBNBXgvnrt+afkJxq+2zYu
pe49Tz9+MDd0SjVV6SSlow5IUo7oa/PUdTb7IXru/L+0AQaU4fr51ip+v3jlQkXVpzLsi12ACrYm
+vGAG1Q53fcXVJX+WgZbKElk6a8PXj3GGxiuC4rOFvF/bQQo0Avz7rbCoPZeaDKsIAFQCYEWzysx
/JpFUH0Yi0Hl9gP9CgxBRSysDG4kr614rSJb/priwOu53cF6PPMzPsy8/6MzW6hq0/yqZP3AE3p1
P7Z8MpkprJqawzQsMJ/PpLVw0mwGSNXDitIa7EKhfj4HboLScG4yaItqMEYAvoKKKP3ksVsN6e1Y
pHlPCVB203eGErdY/q7GblDva09nTsfmzA0QvNGsmfNyWfN1kOAKXyF3nmfcpv3gRHLtcgT02B4c
28dZCrNDqQOmE/Gbfs5zm1KxL8WhqJq0a8IJ9khpH+V7CYFaomYB6GRgro48xXlRma8Dl4MqxNoR
ClkRCdHtGfgKDx2KS3uwzOCFxGCmf7j0SXHOtBhDcnTxXIAFDlHuVXWJakHEgYRK58uHS/Rm58K+
n5V7YkJk+7oTVtRstzmKCQnkl0C2lnjpd0EXtrQwwgt+pyUDkQlruqKbmh4E1aQMqYsvaeG6iAbS
MqKDUotXX3qJMigCC7ICzVPzyi/TYnFRhUgNv4kVUWmLJd7U+5MOEOy2sPJQW/BZoYXWao4bCUTC
4M70zHwUvrTur2FEXfeJYDQ/wjTz7cy5zGSrU/KnrFS2bxZDvSio9BC+91sEqizFsKViuBP9AIkG
6EtiUs1ZOxkFHxuDeLBhQdIi9//1dOTxwA1nJYyQhJY/fWd3qvhonfef7tagJhBezI2a/yH5J42k
xopG9WKTAhmq02r5OT5SRHfspBpkh84Zmc87YJimMt0yi4t5KXK8S4B4UGCIQkt0DtrBffzBiImg
wSJ16D3CuonKt4rZc2SLFjYKb+90Vdylm67GTWLeIXXsaLwcjRur2GTG6gEwBjNkjzye58KaSZI4
hq/mVaL3MNfK+U8BIsLY84QnEBvtICCWWYYvBeBx/aJJiWuNmy5iggjKj7i5xZrNYf+igDeZwVYH
lJwswH9H6DTdoSwWAqCxxGiva+1brkx4TI6DkAGPn0+QiMR0RyfNNIpGwnX6OtGxCr82UxfYrJS3
o1O/A1byHuTesAlm5t2qKFJOjHNjE/pmj6zuC7bR1TZ5XQxRGuAQlHlQ6fTapV2FjtRWGpGCm2Oz
i0GT/Bhe3Gafp5fFzXnEzP7TLy3dVjcoCfaZpwP8n2L08St71bWxPXP0NrHzv2ww5VPwgiy9BBDw
RmHln/bMtKk/1rY0HFqhD7JX3XQmo4gYddkVaGmKyuiKBGGSuJaHxjFCkgndAgaEbA5/nV2NAh/K
FHi08HUGHDc0WXf6t9LbXxWxxKoSvf1f1HAgBuMHGxSDMMR/NDQWhPJs6fzMdazoELmssYNgrhcp
YJeCVjEz5V6OeroGsUvQ431AkwaYisVF+QNT8qBsVIlLU0oo74UyI9mDfjFw3lYfoqxPx28LhdGG
LG7jfMfaHHzzigl2NtPl2McDp+qX00hSHq0ZqmiuzxcbzJfiCo1wpyHDBoBITKExbXEjFSs3kM7a
1GFT+I/HjG2CGTBQ+NY8vZBh9qCqit/0/53DgQpx/GHbwZy78eNUXZ6RaKG6mTtdVZ1jRNj57m7a
gcoPw5zVXdSUcUSRA0ElFlcuojLybeZQh+o+wIY8zAQf1RqwVy8PHFnsU7soFQRAlDELbqQKdAWO
uTmy4L8hw0rlUiAHIyvy1NnOubkymAn71k5mOH2s/zRBrkNOq41Pem41RMmc/iAaTZMSRYLFuJUo
QgxIxj6y3e1D/2uS3CCRDLBab7vEBxxjJk3h6icFXAz7HBvXJLUYjPXkEZqjVXdpSbB7hsxuigS5
9NtpLQCY8lFrD2fqKjFETIzRLOm0nt1hkZBEaAOpioTA9/Kxdlid00Hhrn6exxQG0zsTdoxHyYjV
J0wFVs7O+YJ6euwhBm5oxgyaAqcbWNc6CU0YGTPE+xPz7haHsFrbwQ+8yTYWuJ/ZqRQxdcBfRu3o
5TW2KnUGw8Z2lwmun33AerEninMZz+qqoREF4oE7aoa21fYj/1KAmT/ZMZuCb09qWQNm0djhUpYc
dY8M4avEvSNxbcCFdGrmHKtUFsCuDLNjDCotCZwWVjcYAWFAz+Y4agPN0v1KtJCwDUpCOdNQfget
YnrkaVDxtehe3ztrcfZKEc929wdvgXIvfLl4/+4xVAfiw3xNcvKhlMnls6JIOZKc7oX5Bh2s0Hhn
MD2vX7BbplzOEqvzLaCoF67shlQc2V0L96GVCSfUVjgzWRbfvLXlu3ohgvzhOAamjJhLsi0Eyv0h
7bJQBOApKJ/IbjTbESZaYXRVCPAwFiiYOWI3Qkxj12OsMdOLFNCnRcxynJMIIyQo52j41EjHGHg/
Im2qUCsRa+Fqch8LJsoghj2y5slilAW1LC6xi3NG6iMVOVnirSxTc3KjhJi40FR9OMqP80TLoCr7
3OGqo25Ln3hGUOX5gnm0e0dTUtUz9z8429BrpSZ5V48MDAXjtm4h44dY163PQ1l30G3QyS9lo58G
3dk1m1zvtQh5d42pSIU6ReRXdJOKrti8TGCtRaR8pxIBw64qt+WnN2+nvcJiU/Yc0BiDDJNJqXLw
Kz2gJlJ7z/LcK3aH8lVJzTYIfk+TiQRV9ItfrG7NFeZUgECBg29wlOcY1MRlGve+FMTLoU9T2PwS
bmy1exVnFl00zF50YRBs/088oYbreVjKq9J7MNivjs789425nqLKKorPMN0oyKeN9KUb7DDweQS0
ma8KxjGaJb+XuONW1dtc5d8FUnnwB2PtgOrY39r9a4k8JRgvu8fw/1F383nHuLDrxd5LpFWVwDpo
VlQH90rK1Yga7omxTOOT2UjLnB/Q6y3OiSNCgxtJY6NXKwi9LgmF8prLsc46HJpW/xHrkY0EreMB
KIft+1kGt/Z8UwYLFE34V6tMgqRQ2K+BJ4KVc5H7xP2nIZ4KRLo9sQ1SZP0ozXCtV/8oa7QQsLRc
EVyKcY59K9u+cxdYBGFDcV3sa/lMJT2Y+u0N4jD4qDy05aZ3joMAOm/LRb+heYY/cuXjvZ4op4ti
hTM5K2hXvequ2fMrKkJfWSF/x1Va/qilcpYDhyEVIIursX0owC96WIZTReGwcFixOweQBqZunS/G
xbmcbd58Nh7ZQnooMUsqo5MvRfI6bBJkZntBTt8QYgFTcbHzvWLUr/n0oA6vBdLERa87Y5JtZbtS
iBbuj0QPWYiMJTWI/3LHHuubYlUEotda/xuvMO9OX4v7hnP3/WeZneMUFZGyON67/jbW1q8luxl1
DCGs24oCQoFpScMFOfFEa1zWq5zGGx0IBGw1poh0S/EzndHYXxItx85R0Cp5LnOSrQKB7geIgGuu
Hqqrl4koXVfUgv+JbOYz60Tzyi4X8JCpvYb/Zh4UWB0RGItypu3JDDoiowRMxoi1cvdAISJLCeA5
GfN2MM3hXIc4YlVV7c+XNLBDtIRVU5qPxPjUBchdta+YoVf3qzHcNtmbt1HCwHvDy74C27YSLXu6
5V2NUuiCyLWcBeyGZygTRsNidC7T3Iuit+vIp3ED7GXF4FZUiBertwRqAu25PMf2b8tNnIZfR+vB
AgmFkQrqQtc3JEyq0BcmgibBJZc+z2pbVhtExoPVqcXEjH6xTWs6dm1bp60nyD7UdtQuKUG8YM2C
uyxM3X43pR09yJMOnoSWXLV2aXIs3lgOnlmCL+POEj6XQY7BWIDEJPlpY5fj0ut6DDZdX6T5H8K6
qy8DDdrJOB2p2Xpu2bgqVZTfMpiES9z2Qix2LKXA1lVxVt3NWThYefLN34lkv1HUNtXhbuKN0cAU
5ocxMISa97IrNRLzkSpuBun7DzSbJzpdlXGlXW5nLx7K1kS6Jlay0Kjs1OqGfjV1ftcmThrSQ4Xj
7FxkQQrmyEZ95V4MQl7oCwVxCXQyeY/vbp3JMvpUB1zsX1994EbhUVKLtN5qh8lCmEcn+0InCyGC
8+y22AFJ6b4eOCBTSXkKiDaiQqkgLN7K5XS/qK5vKxtz/bJatUbmZy9OXEWdXWpLdrGAQARRtEjs
cJvDlWv7sVNNfABraYvvqmyu9HZeBx+bYJrr498dCM8nH+QwmLMVVnjswEP9iN2TQt8aIWzMef5P
8wuOF3PvLEugfxlfwVC1b58GPjfcwo3IUcq7m5DXaE/AmkWPdmjJSQ9RCVrNAWhoL5cNPH23bEQx
5rHl2WlwWBz9V+ahHqSgAbVXAJ7sjSxs361FNkwMocEnoi2ZPG4hyC43HgTwYWES1y2UizbTnOVr
tvaI9/tn7PTFn7utcfcnMgSzb/RmceuIzPYmpeHDObmPL+u33q9+UugGpZdZFsqMEdvUm0G/8my1
ujeT76XXhc40sq+G9ciIiqM9fBuLNsTWvIqhBNBB7ineqc8QjWwho+hPOco1t5XqzuGpBiWg+Fio
aMrFO6JIBgILvRH7mX6nvuFpW63k7k/9xtHm/66+m62uDWU8BA1WcnQhcVVgdjdBWHxliIN1BZAh
Jt57hcDl7+SJJs3WjSnB6bizua73Y5PdWkqHOchm5mqPzb0K4+UdDNdBuj+VUdbfWfEEQSVIxE4I
djHXnJfgSGrU/Ee53/pRlg+Z+R+lDyfpFFyf8WGohcUgBxZoFiNmp/o62kprPqyLDIHuX9LTQ9yn
BA+jY08H6Shb+yVtrnkVqQQYMeY62PWOq98FBtwbpZjIJNi5Vjut7aUbo4vp5kwJLybegOiyJsju
B2nlh407m+9l10EBK0Zn+bB85hRPQ9S9niVouDiaghhDovWeLFLVHLuk1HWhDKLV4M4FnyWIYc+O
20oGuot0LP671RmPnYeK2IKLRCBG6/RGM5dCQ+W4oERVMv/GnW8jwqrMShfZhBU6VdZc7VFKn58q
ojgWhumnxkr+CXR+/ddSA3CXi6wvXTMdxih1WrZX2uTrYsdmQrITuJq0kQypPYdOTOm4oVEOKptp
rakrNWxjp1t6a8X5Vk2vElKMfML/PPtBJQyivLXsSG0XPgPzlofpn0lux/zxEGIiPfbWz+P4Fo9/
YS8s4rqqWF7HdRM9mN+7o70xVAs63Ei1ptdamtqiVPGeP1m6Wx2c5Am634AsDuMvfqLmRD8kcE0u
BvWQESNzRLw2aCsApCw8Uqdqy3gSJiuthAeFikvc6gCuxyE6Lmv/2qrnURAnrHjfMHGHQLTnq2ku
0TxGafLN93LtuvcyLSQMQkogRBt7lvwmBP7cPBC20ZALLvkVqV4zhl+PmOO4rpc0Tre7idihFIDD
8SFAG0IIpvp+D8CXEAHeWfMXTJzAgRsGVsanNnbLLQqnIcOlytGvUhvmbRlup39Jv1TfQ6VMbP5S
ZzWlx4dzy6G0pBfmknwyM/00+fZs4iGausaSt5r6lq8piDcjO1trfMdsWqbWykdThLwBU/op0rTx
ZXo9OEs63aTku8dMZifEm8ausUlcWyz9ua5gjMBDfFuf7cPb8uKZkupSrE9WEfypDXzP/6svyDhg
ueHhwKwwgO65/oJ2NYxHcDspnkmRRdh/HND5z7oY2ewkR49DL2/wikzcPMOuha/UREZ/s/ZchnEV
SL/xvwgn/L8y+NTE8TQrL3V1DY9tU7KPf79iB004KPteld+5WAsMO7YjNWBxsaHMzGmPcxRXKLC/
/OuQub8DQYfiSt5/Knc3bKTrTsUB/lECxNdeVR2mRW+xUvF4DxLgQ1vX9VtVUdREPF0db0LMZMr3
riFsev2rC+xmcB31AdGL5oW397XgErsNzTPe859++t9fSv6VAVzTqFTTiP6fUJ9kevIiY9CZYRnx
qxAdYnhomEL95Ha1Xise9ctTC6UpCrA+tslfw8sfte6WNHhmi7zeNDTOZazQs2/g+JdVhigOkuV7
WK957s+pkqpTRiUXEfSWF6bGKHSyHGWZjxsaAvdlcz3hVQBkgTIO3WbFAUgJHxVhvfBGAC8XF+S0
3/dEognPCRlEp28JFUQk09RYmWiuPA/NhvAxDwkwcKkPBYmt0Fn+YszuNoSiEJWukLEgu1WQyvfc
CjO4rxx1jFFXATwLUVWPuuqOj2wD35W/sWeBqvoDyJuqSsXhZBzBjh5DWtcY8AokJkqthW0gCGOo
tbW2UIvPoRpbjZtIzz3mrZMNPNRWe/XgTU6CnQRtJwonDNvVj1CvJABgQ6v0N0r2fM1gdLG6Ce4B
AjlfnrCa3H80nE+KXsk+QrDIqu6pV+119yxI3oMme+fDU5nuJxqP50ZuNmFKrZrpaGcpDDk0Edvz
QcWIwEJfygaaNCEjfBhpmZedbodmpobFQ/K9+gAyVhS24b/fVnOUIWnMKBQv2KNgh5vGKFPRs3Nc
2pbyZBkKcNcLpLcBTW/0PeZGAFw46m0a9ueVNjUppDRkg4UDU7HMZvtO+aI8yjZtNiBKSGduV0fl
Xdkj8tE2236zyBkl4rV9qK1jZ+bKPWjxTy0EzJ3DlVrWj+3lvcfmRBo7PnHqlv1lJRCa/4Y9QY/J
a0HH0y/ThLRyxzpks5e4q+wzeXT6TxkrPq7cn3TnTH2ayEBkOBiRBiXGVrJKTMB7L8IeZXdY0OkU
3R8t6h2D+mz6oGAgJT0gOoe758wN9nSxh3qG42ZnJ+KiqDfz1Gmn6v+OoqzMdZ7eLKAD0KWpDROk
4KmQGB1MXBt2pfNGXpHjb9kDSz/eP304sFdF/FmuT8luVzbSqOHDDVoFKdp58z0+1fiU9oRIk3zf
BwMR4smue9jnplu0nljHu5e1YA3ScUNaCA8qbgBeFv/iBuVbXHamtQuml7ys2IW5HXl1+vmZI8Mg
ShqkCyZpv4Xqd/q6f+11Uxr9l/aNJg98D8EJkSSaESWL5p23ceK2k6rzH9YrbHDP/HzK+8pKdnV6
BsRoGADFBstV+Cq/cwX+umTP1eH5snNXaGwEXYM9C5tc7a8hXTmYqzbMJ6voZnBnVOI9LMwYa9Ch
QqHsOwQh74neszNUv1A6yiu/SjpzUHqinXT3LBC5eE0zYT4ADrLWyjDb3d/4I1pSaot90pRCsBsT
lymAUBtzj2fyP1K8/CgE4FDJnOsCorO87seG58tDPWjLgYt0zsNRMiK6OpFxULA+cdXsuL88bCf3
78b1Bkdn0F5epW+ajJEU1A/TKHuKp6o3qYpncu908wVgX2Mslw4Oh83Z8RP4a7qrt/paqVy71CsE
EbqCEslpEqNuv2vv34adt0jtV72AbFbQ9dKiBiY8zuVw+YlAqwxbvpl4CTRdEVBrzLZanK/GakoY
I9ok1pdN6FUvtHPUvKgW5l5nJ7+r7aiTxG5ofmEzmeXtAcMXPy7ZhW97Imh7gyGYcpyFukbKrmPB
+a3AUlG71lSVuLG7wcVnP+OqAspD0PMyL8n7z76gSiD/hNJ3NsTAntpT+pKFYEQW79SW/Ssw3DmO
zZntat86hjgsCgMWJSpTtGtAOr/+13802OeYjJS60m+XtilBODqYazN+ZKMBFguQzkiSXQkEQ50p
r0UFw33emTXcxdU+metSaRaltW1RfX7Gk0DIS9V8sDECBpTewcBcWvDVmmR4Cru5pkhIH2iT0moZ
D8Q0kH7ERxcngNTQX7h5rcqQWXqV6NUYB+lAGdEuF24c+rFVsqFi73Ptj5uC/zQR0NlyuzkmTesq
0SuivRyIbS/oZG6UJjNMhKvrkobUyNOey5Xro/jfunmT7muDTVJqXSrVuRa4v/DxLbOedQYg4aw5
sUlm0F/WaPP+Ui+t4D0ZXSFDNvXjjAaLCiSIQ8bT2OG96YgB5xtLaGi30XOR301d21z7+he3Hm8b
5E/xjR70JbFv35sYfFv5jR8KxflQ3vfEfHhDcSTz2kjJeVEe3WpAldXgs8ZuEMHl4kmA7kP9nZiJ
fwcpLgPDfvcoFqx1wAoC+itJ/PcEMo+72BTNYPK6m712+5CCTBrTaGP9ZAApGD/AE8GY0y0P6toT
tsmvv2nmnQXu9EW7ULqtOhMPnIdasranxN0V0xmYkG7PkQTpoKxGmry7YQgvbm2AbSYlesQHmPjE
pjg0mkCrSyk71YNDnIXbuZEtcZ4JUKxK/aluctryo1p0YQ9oeQ8r5V9C1SwUTGBoOvE+qFLa1MBx
jpvJkpchH6DI58ElCpP87uiTQHQ4ET5C34TGk8kZT/zUZo5Tzb8E80dXIudwrOhQzvrXzKNtdwUX
3JPadTPpbQ0Mto/t9ZHlRAzjkUu69hDMAYRzxgbWWWrw/sI1epuAfcgan3Am31cVcnydCakR9zPT
faCbZRLCIELodK2dSrFPLvwYFUMdmBTnxKA2V3C0r8I3ez8W5D35k+YHoFsoUONTp6HPy+wbOF95
YXRFjpO8Pl8qWzbmwebWK/pQ97mOVincL7l7u/cKhEIoD3DVZQFLR9U71XdWfp3dv5H4oIMzKGst
tJFQEGfvym+IHz/Wrie9JNSUONMzEndQF0S4Lwxr/8Su8HL5LLhjX44Oqti/vS5w8WzfuGMY/b7/
05XQ3J5bp6mdwZ00BjDdHI9pFEqQbjOLmC+XsXJwoOlu9vK1Z3qkhGCGkhXbfZf8zEB50LX9WgvY
MIdyXFvNpCN8weRvY1000DxT7tZ+XxKqaCk8nQNtYXnQYIyH0gMrGlPh3+LcwGPkQgSZA/QRloRi
cfD+L1nZuzNTgwq3cZIn/dWab8ETuiiiIVYcHDqm4IziFQTXGBfLOsH6a6KolmHGaOiTUlQxst/s
im0cEzyIsqZC8PJu+LEG0VsFlpAJuLL4RGDIXtTTB8MUmmID2Wq91zMxMO6dCfOTy4cimIbuno0G
S0UlTOzWcTPJKtrvhOCXdGHA9fRPy3fuHetTwOCpsDs3Lv/mRJwZyBmA2T4HAHBB9O/rv1g8cKw3
unopseDztwAhYUuBjxb7A+HU2gdfMx/rkqBKwS/oOCBN/JFwVzGYFlo6QvBxn7rxnIZUXho3Lepp
oLpDSL9OgBEvkQNMV8SQhPpNLnEV0T3Hma9yOcm+p+rXfVwD4L8gD9kXxq17MpqKCm+iqjcNVu2/
0oMwsUvT1jdldsZEhOOAo93I6wLYjTWWXONvxdA7126rlqwD3sT9dfZftVZ+xybITtOJ3PKehszu
fT/wbpmfRuO5nC1HnKtfuErBxotmDCq/6REL2FT9sETpPEPE9VPxKU8tpJ0JlwJnFUt7fCuYSz8v
Nbrmjk3cgL5FyOwJDz15OA9K9JGi7Kpaqc0MAOI1YqYFxAD+YNyBGBVQfeqER0rbUZ+O6UXYYD5H
HLBQFKmCi5B4+8TNk2vf5N//Z/5801WnMsh3vIQ/ADtFI4yByPRpYahlDD3Fb0/RqNL3hOctqHHR
Ur3ypdCey6GgG4T+GifY7EULJ+XIVli1KCeqBkgfLbDE16CFrmgSqxh+QhtN+MOfjstiYQsOuufB
lXvnEJGJKNypZXCbP1u2T+Owgv8grtQsRpW2CxRk+ryJj6BVlf1p2Vr0W0pnSTqgwf1ax1qbOoXu
Y7fR2++GztS5VRlNDBb69twI/rqDeeXD/yDNWtc7ys3tKUt4kGIeptxKHKQzFJfVcyOO1TF+N0ox
hYXF/osI8LnDCSLv6ihtsiUQTBUGnqqZtq+k6TedUQhGFDS7kWY7Bglp7+2L+aeVBG9vQfA6+bih
b6OIiQiOBZVzWJvPkQ70jU7/tT0PQ9yxKeUth+r2tnbB0Dcadwhcl6vgWTVZhQaULBLy495rCera
xs5bUsmeYUP6d8qzEImeQYNNaMA2MhLDi/qw/I/ssq50m8uzrw0Kg9MwfHkdEHSxjM1ldFInjm74
UHok0p9/gQHQyCe79wrpjLsZ01VfmleE0qlUO89JKOYi2zyWVhrEeTo6CW4NVeH9f8IAURmWrupC
rPzNkgkPQ1IrU5IY+qgyP/ijIFG17QdVK3S0sjiBUAeVjgT9lll12+y8/HL+beN5AE+IbNNQk8HR
CGSRyjYAlBR9vQp5nTMFuunVdeMbagWvoKSxjsIYgCnd3zCAhuICX2h2boT2i03ysjZ9M+IBFShQ
ZYjORiisLzw3hlG2yxkKvFX/ozUu9tkHbaamNbQANUlP7kYhh9l27DfGXD+bSgFw7dQ6qWC6gikY
4m+Bk+GR5ppD8mEXAqAGoWXJ/yMZp7i65IT4nv65b6jQb3gpk3Ye4nothSaS5F90DuxRGM/4S5VS
oVeFJa05KGfttUjiK1XIpgSoYNbiYNlRTWT6VRzGN9ey7JADmRgXPC5PeTghVH38PxN7xZEGt05U
5nysR+UcxpZmvCpfOVaf/MBXg0wl7i7x3jUzr/GbEManMlWKrlrZuhJcoziSwnxyx3sCQT1Mjk5w
CSpXWmg/FzHIxZjIfFrDPBLXw+jlHvxLGVrMEene3btehNquIsYA3pjizcKt/0Cx1VMjWtnixvrq
VQmGCwoSKi8kYi5cS3uWKO9+hHUfxGYIz5aNreuI//g8MvqWLwMpKqCg0pTryM3/vQ7al8+PdiCJ
aW8SXSjeUQx356JEMuaancuzdJwWeIwuWl3OCm5zU1z3Wquizdmh4uQ4uHo7y434d3ZVVCRoU45i
I1JGGRoyBESVh9vJ1dq51RToCf2JVUKK8rW53lA0RlzEZcmAHZm4Ta0KzAvB09KpOhVqK0RYtEwS
wR32WxsfNLpPTtZt/SR774rjJYD+YwBirAmkSViu177W6L90HFxM0nAOo9l/xB/GUlAB1Wbv3DTv
JZscfPnsMdwtviW6FoISHF7IsFIQIQ7lgJEKL4iUbWQA+LDa9mbbtt3B7mqbO//x4J+wz7PNRCpl
y2twqi4Gs11J1LlXdvV/+1T/t+5ynBYslheXsjSbxXnxHOPERNZYyCog9ZBZYQBQ7QrzuFGisld1
07cR2IRp5L/rZyU8KqJEfWfxt7AYIFeS2dh5qEwLXFNfFSt3SlMZ0ewGMCIORtjDPIBCwfSD8PBs
5iS66sNPrcrrcLlMuyiNGzDMmof68+9MoBuQT+bELx80P3cM4BiemaLtpm8IVJMHKNM82NhdOCRI
j5mLE5FqH6MdjgS9wL+Fb9WJhUm1MmL4eFUsas/WNDOBMXHClSG+M9acndriptBx+wNzJMLQ+Puz
Tg/iIe8iMUJI63aOGBeb+cH/IW9C5Vh3ormOxHoPq5bFpG7Trf1rohdq8B03ChcwGDO0y79J+Y8r
gOh1SNYxUT/zFzzZ2EHDGMnLUHMDuTW453TuKb0zI/j+xfp8Oyr3jH+wgrAXSboid7FvQGPrS82d
ykqSInMdMhuVqY46saZ7kOYN64dws65KCO2TREVQrbPeT4mX/iJRfhWqLJeH4UrAkO7UrszSwuK4
ttzXsGmsS2izFCDjvYGC1BA3pprJSDAftARsIW0Noak2XqLU5FygEEY1hbG5GsI+f7z+3FTVdTmI
ecpqd/9uPuisUBgdezRSy3HqRSlAih2+COlO0UuP4HbwzplXuWC/SKZnKlTbhKTa1/8SZuUG0sdw
2iU0XoqN2xY7PWlryjQOY0VrjY023llCpyK/Kk6fEC79st2XlyKLhLitO0p3WFiJVe3W3cAVax2E
FcYCf3FhsF31Bxh/uzowONF6g1wLpMjl//dAHSKRkMJUwJFj0toj28V/5aMdpg6JEK9OlNvIXqcY
b4i4HufH1XhUL/00oW7kEC8GL+yVWwnp960U64+CushC71m7+8rtahWQzsdEQaMoUQv9liKH2lK9
dnlhgPEoRQkD/3o1IlXJPH9Q4WHAQXZ5erxW1/gQbAKoYsxzplxYzW6Ug5DnE5ibdvdcQ6i61vaG
o15Ts/0RA9Q2o4r9s1KQct4psgPjX8BObVEVinkOFDmdtI8GSauUrjLzDsrtwX0yAEvFi81tGnb+
Baw+1m+YHsZ5tMzn1FKH9LN7iUaWHZhAu1PpfiIwIesieVQasKLEyocQ4o0YvM+ppeslyu2bp0gt
zLzmt/O1uQ/s7B1gL1V4EqzOWSJOLfVFjKoxK6E2nKRmTIEY1cV34Pm86TwzSUUtB2a7VW6mX1G7
ydKDB6VV/BgZox7HhAqofsIXsNOAOnmwQxXjlQIxwtvYt98vXbaXNYTocm4NkRa0E7KCkdz38RpV
LNgsitxhwkBAdi1AFxPgQETr99LnXE8/J9hFatjQ6dz3/0lL33S2yzyRXCfPOrtrfupnhv9KKbOr
K3AK650M47P+rdVUcPyYh3QARbtG0VdUl/SrvvoW8L1+E97zb0Ul+hCJXTVIv9wVGP3wzSgqur5V
xXIzMeKFE8Andr9iMpxrp8nr0q20duTSRXkZoN7jWv13V8sukZ5+HOmCHeJbPy7mAUaCT35M/rNx
cwSw4iEcFEHnw3poKKnQ8ACCDiWFMibHxgl3j5rIxKmiskZ0gZsC0ayFhIHKzvYMxgnd8n4QvDRQ
WKIwQYVeLAEk66Z/gOd8TdP0j3czG2AGu8bAh9IL2qUI5ZrNkTdZAO5kCDa4lKy8SG2GkRIlh3qu
Pqs9fiJC02GjbIcfxu4SDgSf0xPKnX189OSUEs2jUiZr5LDYZ6ZyjD3fDv6aSHolVIk21d8UoQAA
uOutfH0TNTht7PggS5pZFdr/w/GDEVwhOtoOCrV6LjJZgv71/iyj5MvNR3MlAB5T0e78pCW43YwE
4SI2yI++YPIAv610m10xsfSZz+dd9yVAF2pnMGs4CBcQV6CujLJuqkSj+i7932VbRaWtsDgBUc2+
QvgY3bwXmOCu3lJxIJsagVCC2heduYnx+aEu+xdkqdbgDY8nOkqKVXV5RNRhxVF3/JcHpK8IfsX/
G/vbJqa3Wo4CEF4je/a9l9fK6r+XjTKRCDaYtwalGQHv5P84lnefDmN2618fLjbUsSAXgo2QeMuy
rBu83XzKpOzsbyMJewB+G1Cjs1JUyo0jWdF47f/oEyJknelc3+2L+MbtUbBGkqP2QcnDYW4zvB3b
6bPcWnOKrhBHrLC+ePHOFhKG+NpYemQ+wSCdcWlRHgLGnzj02WdtRnBQVR+q+gA5vPzzl4i4siHL
XqzrzBoRAQulnzgIZPddQB2MPCeLkAeYBEUTXffhOcwpLDlp1ly6QOxDZq1VpMSy4PcrSBoh8oVq
zWdPEY4w5Mvqeuh2tStrLacasKxiAEqNRxMZZD7sR76GdAT2yke5TPes407nKo8lG7XBzrlUwiRT
xwoO17lo8qKPGn2hPwWwTQcsVE1X5BjYOc9CukuSKFVf8uhZevt4GADlPDbgOgBGAwL52g1xzECy
gRptzY0Fj+MezlruZJqrWbGtdYjxr+pSgycPS/vCZ8JMmYmUHzyYIHj4rSvgaq9bCxHJVa8A3v/M
y7bHZpD8oOsv13xPeaL/TewTapf5qlm5T6HjOQ5j92Coc8MINsDvkJGq2QgfNXwQM7jpACvqXjFV
RyrKrIyVFkx/Ac8BO8JTy+w5TCKqkKuqX9hUjVVwSuX/JOWWEd8VFs0wrepLrD2zy9QL3831XB64
ODF/j0SB367LPFYPnpkbBXH1ch5UrfKMelJj9T6pqPLGJGmdAjPWCaoX0vj3SaMtf4uG+jABi/5J
LgjMjo2Kv45eLvxLxABkkX5wSdnAdUEYogZAVQemdL3SIiUZ4JlwykOmgdns3Mha8h/QVAr2bJxh
QMaPnWj95V65qEhiMWVePdjgcRwsorqzFF6e+AkOaeP9N4Zxo6kWn7tjWsJh3Xb1kRkqoOW42gFR
XAc2jiyVFTuoNJEwM8dV4aDp0QrZCcjxOzI1nYrTDnIKoXVdgXjtCokZO2aM7zbrPsEBpoEZD3+q
P54B1gmEkyTLwKpxKGLM/PIjhCA05unNDjopOh/pztmIvx3KPb3QSTt0dJRWkkKizCg8PP3uYO/K
YMUxSAwzACin1COv7bGwIxGZS0mnV59ojfgH+a+JBdDb8EVT+xj9QRnXqOuUjr0Rneg+Rudcsc1D
JCetSfknYzYzpXYznagXEtye2iPtUee9GKiElYo+4+cpihAggW1aeHGwHMZwYioE7SVl0HudR7mO
lJ8xNLGULTjRXrqTP6uv2S0dbWarRE8phjdohCV+YJTuI82yK0bkVbnUNV13xHfpO2yT4Wk7HAZR
urfZha0pq/ufq4CuiJKrb4nVQajVsgCrcguZmbDismc+8oLCGev7AFbcWBg+KfQ2VbPRX2as1ZqK
zqBXZGFURayIlzzCysckqJC5ffZhzIUp7JUpvlQn+V0q3x7SprJhKeiZYipZ9LE6bP/Ah9hDZm+G
7SMyGc+kQottnTSV+tViRdN74JT9v7W4unRnc7a/0Ha2ON0SVY7AI+aSmdo1jcDGG3T0dNtAFKKL
JeEdhN2Bpx2B0314Af4vCe96YmuRKbKc9lJUBauKdE0BBrh2jgGQOyHMvxgsrCzK8SIgdP3ARzFj
v9TuM5SboQrRfgtWVmtG8VNkJ4LnWgJuIGqDHJfSdiTIDvrbCa295aasTVO9+4EI0gvfvXsQLxP/
Ig+etpfWdY5YKAkcNRHwuicV4ITQVnI2iFLyYS11xpAvLF4fblPdHHKm8/HB2QBNFEpAA/rihccz
gR6ovmn5AlB9WZ9WP9pXGiV8QkwRDkT98pjHZQh/5hRded8HH/WihXLp84VladwibTPGqA59wl00
IAew7SWbqobvmbj8J/C4aA91GT2gpePP4ilISrbCU2/WUxwvJH430PIrrR3GMimUUU7VKwTt9Yf9
4DEoMMs9j5b1otJwoFXb9saGnQO6DDyq3Wp2hSvMXgKXwxANkqV92MBD390xMMJEUZZrOjkYvZQb
faAjP0mRJ2gWv1JYn35rTQPVNdzNohVPn+YFq39NMpTXFvr/LNmFoVXl9V+fbHgroB5bqyqB51Re
+dpD/egi6D9pE0dAb/pGZ34jNX3kt/6YqFr2cbHfrm8/EwJAH/pioSJ+X1yRb/Wv02tYBeW7XzSp
MyjIC1xRjCZI3HS0E+4D7zX6xiXhcJMp+yGaA8R1OY0jGp+cVsY5QCDGq/wDgFaO6THqfcRXVRSj
Suo07aMG5cm6
`protect end_protected

