

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gQ4CxdvWgnieRLRQ2AMwpJaA+X4QUP23A7mcpTzLH1nina2JWDwyro/SbR0koY81VxQ8tVNBYSg8
3s+EjSEjvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gPnHmBrjBHDleV2Jfu7AAgNyinLiMa4GswbueiHBD8y67DvELbF4ryETXsYzyyRC60JDgiQTY9xS
mNBL0n+tguqX8nripcl2WvUcK2rEIU4vEmrY5Xa0k52V9uCE29ruqODz0JXngqZvaosAn7R3hB73
7cI2IgLWPL6sayUHq1M=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bim7wErRMWV5FSeSCuJLdGVUUYEH+U9HzwEGlgElmMU1LE1rxBL3MWBw6E1Qg5kGmxPZcrNQKg7b
PLZUD5Dv3VyvXW/HR3jI7P5DnwdmPcuCjrrkZwCh4jjzor7rIj0AM8ubprUHwkpicj6rKGNYRGRi
+lmT6hjwlretXlYwE1YClKFDSDei0UBfS9a5tRfCcNpmoCaImXf0uTOJ8unbujREQZSIp1snYBqM
Q6qvNMpDqcLoVSU7OrgHQdnonXWYqY/ILDCjdL1o02B+xcnkuGf+oGCDs8KSCPuzYvirbLqI8N91
feufkvRKEcc9+CQ7U9kVuEQ2Z+MB8XwJtiWwVA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HhRynIQ+TRImN/1ISEgCruTQGOfZ7yQ0AeSPRr1UgeSXeBV4/j+sqUVwy6KpjxjyOB8/Up1pUaXk
C62p4kvtT61bX2llnNuuYjikfaIxGUWJ2S1a+GpileS7Ui7iwtZy8qreshTy7qb9L+4SycH2S0Vs
ofqZzZCA27OgdUdAA0M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RhnO7aE6HcfX9+ngWNOvpaRDGHOLotkXich9kwwYcDEBAwcff538vS/s9YC3iM7OnnDBzfIjK9PG
hZTnV6Wbh+heW3iD6MhhmPxC3a+3h3Xr7G6V/gV+8tP3qbjwLdyiI3Y3Tl9GXzeddtSNdvaD6764
1AS1CtRtG1cyGvfnXyGxmyDzJ91rqIOqSJbBOVjL0a+NolFyEU0BYVthKlZ39r7JI1kVtcM5XAND
LnFrRp5p6iEzVZDFdricPTs3V2FwNDnZSvZ0QADHlENUl1ofRaFRtXOEIahTDRwJJzBMRTba/K/s
3AtKBuzpWzTyvSqo+1PWwgrrClt60fAvHko0Yg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12608)
`protect data_block
eYCSxuM+PKCTUWRlqOqgPw9S5qcPctlJFUSMiepZtjTUpF79q+gbUTjK8cDOqnYX7xxDyISIwVON
wpWOqYzFDLKefSVi7a2OweWhnqyxXS+NjOR9in/3wpV2lgsZGeRBu2DlZyKGxiQlfOytcRsIQsCz
woSTLU3sQxQkuN4pHHK8nz0dp6JT8G4MwgQ6kItAHowdua1QTz20RnTP/8k5vNipgQ+31EeZ6lBZ
rF3tzzaObSG8m8Qnr/LeO8KzsJ+tF5cwMuckynjAmxRzbIQ+mglUvUVESgA804zYZQMq58qXvZrL
/TJqqVcg3OoNGUle+qrMvdcqPbScGr3TyyLRxT3FPFe70qt0prXRRm7FzCNe+TnMo4LIgRmqKsG0
bRh2XnfcU+091cBwRUCjU13DIv7srIGgLh9TDP3DFZSyD+z2LGI+Odt6tDWkf01D/TLve8/zIQoj
hAEOHVd7m8Qd0qX+2cRrqQeVjByVHFenqN7kmJgWRa34dAJ5BznEhr6XUZO1ALx7VLrhv8bFdKWq
rDIZR0p9Bm0XYojRSKkrfxzL0sDqOJSRlQuP152FP02oEVYATsyx5vmdofELW/eX7VRO2X7O+rdl
MabN2VmK6aNt9SEJyWyauVM+Z3y0p7PEUP2LJqOuG6Y7X4spMYDw1g9v7or89P79mRisbneWFzZd
PJAhcg1gMZMrhbIPCUdPcwpbpvxUHdy5n+kj+pQ1C48U0tjWMKQHHkLkeSc/mlfXDR7SgkXGxwxD
6xnha3Pz9Xm/C/OeQRWyWEAWRNFC/af+saZgutKfz99phYqLBDReUf3wPiqFy5QSGTi8+OEYOFLL
u7bQVl/B7intNuM/t5samDYX9knWJFMXFwmInssuOVq00DSdEz/PJpswueykmuqQHyoKRu3lizPg
+5jtV4phd/L1IECyzF+uri6kcxXRCPshDUpip/wJMfoA2YNHeFNQfYZ0/TtLcm2aFykNpANfFfYx
s0LUMlCKd/l6qszsMwiPfGVB6Hk6CPaxj+moXYa+8OnAjujbl0NI1btaa3OaV8hr9wtfdZeyjEHp
+CZ06zGNwZyqz14u6Am6ZI1ODE+PBrZzy2xDelbWodKqUmGMnZsfjU6LUGn5g/PHA5IbwP5NTHuo
enWNZzh4FTtBdxlKbEIfUsi2FnOESV6aOWlQelVlsq3a3AKeMPMevoCVcBxoqunoPKa4O0/AbDmq
qT+gZ5nRKv3sO2wF2B2w+/UHTF5AqURnY7Krt9tSbHiFiPLPGl/4FJ+7AE1o0o9TZ2v+rEHodUsC
C2WZz6NGn7sLj8xHnk2BnXwvbaKte63M6u9evtXV37bFGjfAoV1CsomCrijwsBWvKE9PAM5BmPoW
JiwiyxKX7owIGuXz7PRWVPMBimo8Tj0517QviTqeix/2yBzb0nnmxu9ALszm9OSfwJj1ak4nm5Sd
xIU9pSRKjYc27Zyu9FkO7S8wMK56bdn+wrcoSR4Cf64O9zxVgqGYpmzoSfBvRpQdLLjvneNs4tk2
3mCxbDYmbHrr/Wo7GOPeMtAHgNAbAuKX7XNUj+szhcxTFR+PTg8A1f/vraUUNOAaknt/OrgZopH1
yyyMtRDlBVw1ZfMRVy3O0ZHIdsns9xnpkX3GIUNfXTEby8slLD3AhwFHU2zPqWHrRd2ZRH9DKEdU
FYwsvEyIKvEueKCN80PR4VBS9VVi9iUXs44I76HtHq7FJ22kNTIDLsqftMjdVmXK7KsFvSKhabOS
h0r3ixwNJNOx+NlpZBQyNl9Q+rRAVJeF6QRvgyv0fzdPUk6XJuDwNoPrh+u0Umjj96ajFuDWwmGR
HosBbgm1uQDvk0QB9tyjSPXU1caecgts0m6CfDD04BhqFBP3fOf+FARHlIR7VpYoiR/GQwYApq0I
dsFZ9RnlGepguhqyXwdz8bNJTUZprWYh8ylPGr2YCMNQ9jl2A5ff4EpS0Z5e9LH7vGGiqkaUCcq2
G7WBbqG3thGefTBWHC56wVvo4N1bnFx10dGgDOYrYqqjnsi95UObN5xi9yYTIuZGUThbilCJuFkU
88N9VEGHbL+G/P6SadxqVFR9n6BYmUBzM1IeOBxze1hY+fgPZAsL+1UhE+Bjk736eUbhN8fQGymN
Z/UkD1mqPVM157/D9ONblpN4X4bspwjvw2/8qvPjNQXdgd/tevrIwCtSH3Hl9Da1NBuCTDF5Xhgq
IykkL7BhZhutMuzIUCAPe5wSNrIrUCPpX2jRm2DNt5AP5pnYTlwv23nQUcKYJZgnBcTh3ayb/4P+
piG3RFBKwOqOZhfWaGcPpU8BoOzUzdJUDC+TU1/xPCsGJGyroIvhVId4EolNS2shiGjY55ypiPIS
q1o6eU3bS4Had8QVIjtqrX+eVlzrvfCCfONyUcUYEtwyyXSRGC1ww8q2N+v5MfTdToCp3aw7tVGI
HoiHyN3wQmYaSCRaFEbtWCTnv6OmHgktCKMtdtwggSX0HUi/Alwi2V38A48C9T/hppyyofIk6jxw
T4K5fGarqhoMvBcz1YYqRxbULrOaREqQa1FBINEs2VGjgdD3Bj94SOLEQdDfzFO9mazZI5VRYdw4
na2aSzMQVz7vQgg00KcCT7vjECaQAGLTuJnU6TS+t7RLSN9l9SHjSBoxmW/IYH/I+En6Rm1RmBHx
FdWktygmu27kx95qhocIdTICY0riYgA4VdqmGb/Lw4MjtErfZhbVIp+c5gN4GYK79OVvXLhYnVsd
1FteN3Sd10Ft62vHH3DUA23rhxFmcp3qxE29UGnkcurwF8mOsf7HwBLhVBuiMAvqbn+W6oNFfAPS
MDZlS7WkgNX/0HRL/O2dAFjTdqbOfhLBCTqfC9NuqxNVNUZOiN4n+10E20isO8VNGMZ+5ll4jVLv
P/ZcmXagrUQLHL3XsWNp+hP2uDQyY2iTQQ6ZFEr7gE04kUGPqcEZvFwUMuCk50ouvqhe2cBfbbzT
cIOVnm7C91VV6JHPuHSTUcbk9d+B1BivCn/cIY9q7gZ0M/764N65PzNucB4ht6kB42LkWeC7/9lx
fc0DCXfrdystI2Pr05yPIje/F+vtW+xJZJBSr7XPurDQTbWnd0IJlhVn4GM+QVgdVfkTq4MTRQC0
EBeawQxq6XdQOobbscWfeDaq8Zh8vyUIfMm05AY5XAWQNsRBi3kxDtR99674rkqdhnLukT0A+4qT
rZp/5Fy3vEdeZ3f7pjP246BHL3YtTJB5IvlvPaSEBT1x87+JyzXQoVscNP+fQdrilMSZ1gpYG0sZ
GS3R/WHTOnSLvc9zRzsPcUQXnRnVa/KP71NOlTr9CPV9frMGLMTVC/0YxHaGiwR8fZXPhsxAKaZS
JIUwrKcJuk+UIeNIbljGYtdb4+L5Sd+2VXu3wuxv7ct6qjpp/i1G0Z4CuqiLeNmV7dSVDpTRIqF3
ggCv/XKvdE4L2fayaVTeF0lZ/C5tpdHbdiHC9gzpgYjwTONFqTxxq5033S/yO9I7dnwP1b6MVrPs
R7433oXsfSFwZwpOEfa/FHqo3Kw9S9pUaFP7s+CPB1Fs61+01Lm1g/ML4u7rNoHV2KiM/dNQpDrb
0wToie957xWLMOS0t/xtkpFttiMHtu/OpE8AvIhyEGvfpbb4epuSuvmj98+v+txJfHqJMJmO4KOR
ZZKgy6tUqQebUBkHxbRxb2ucmUfG+mIh+l1bbriqMfI2uV8AQSje5lScDfB4isO4FmwB5g2jqIgC
Z+70MtGuRYxw0pRK12A9XbFGc6lHf7f9YGuts8KeNBaDSni1JfPr6R5MtAM3Tumq37CkAvGTvlU0
yIE7oPqYHNL965vYPnt3icf6kfBZdaEfLrn4MqLqhafC+GWH/w+Bu3+8EZ5tnArwcPVXYiZkQt+c
0JgS/TOGwW3DSAPW3f4zbbPsd3n9HQ4z3Cnc8LCgCtGO6EVJJTZVvYdbFK98ixBOVtcTPJANM5Gx
2r4Y/7TEe4taewtdwbXda6VtrzSNI3aEafRzLADihuP0GpxLRSY1l+d72Qu+4psF/W0o+OW5OffX
U6EAK2vz13j2UPMxrdFcE4p31iyN/NnJKduYAGNpd/N7jqnLyQwTPIPXUPEYiX/dDclnBptxYpVC
v6syO+zAOn176lrgnwlDiTdRqnufPZShmOYD5vkcT8aWvTE65XHM4a1fGIPs5sOr5KTYtgtGYyRK
SBrW8vjKQCtVsBuags4kOw0hPHDql5BTEQcfdQVfNMrEGNDQp0+cCpmSrrdsIlvD4uyapLQ1eQUP
X3wm8yrc8X1Kyz4+ZcforywCunMu48JpXqRxFtGEguYHezSSbGmeUZ48BnACKxfTLShO6i3bKlyW
Li/J2JZC7ljN3zX6+5vRTJVZmJoUKxBRgh1bupgL3LdopZTiMzzYfwsrZROjqOKClG1SMhWLoJhX
NTkBhpy4u+0TwsMfij3HQw8W80x/aXEY+ARYGuG1wW7L2SinJiHIsfOkEixk4SNl7LakjfZmDTXv
n7ywnEYOc0hrf1Kly2H9sHrhnDlAyddH3CiNoqrfjpLQEIOJaE1H3yFapz1YoSOkO6Wn0UkuVvwV
uloaOzMe2U/NTnrhHWhO8lpoTKib1kNOxzgOTmFPZXp5OI++/CkKMndNDO5rR2LpRSMCPQVTKNNZ
zNeKojgZnt6cJGYCh+B188/9/xm+i+SNkWJH8IJ+M5WWO/gFTKa4+leb9p2fZjJvmCSCjf1AorbG
N3HCL0bRJZfP29YVrej0xAyiBUYDLvOJ5vZ+CliyZ5CNRnNdcPBs5zoDvdt+SzEhP23T8R4z75Kg
jRgKz0j+3YtQ94qKVbHUZrCe5m+X1DAxdZuwbWZOPJvnu0I7sMCBaz0d3CnGuZ4uI7AmTADJ+uYS
gOFI+HoICLkmZA5WuLq1mC1eva2gRsNiEAtPVWCg8hosU9AhxNXy7zL73AD6ZNvb36euuoCPTVKs
2VpG+qscaeTI+Nk0AUPX/wAsJJh/0blTW8e6zOWL0gY8z+5pYzKGvBFw1WxloB88dLt5zAvHnjB4
s2UUGZFkAd6nHCoJp7R2jNy+NnkKzUccsBsNm30ig3XZRbmXIbVP56PAeZQHFEVcRdMYpJD5qTvH
QwLFMvcmHpucCLVnADC6Fe3p8z0Gkt4lZm2xOI/lDHeD/6VOI1ahXsorY/C2axzfRpIBCOdpoc5M
kp2KF3QJGhl2rpnf4v1ONgZ4Yo4jczVshneHNS/GKN/fs65UWXDdp+lxNG5yY9emVLK2vRf7+LCb
s2DIJDdTYYKyM2qx26OyImnylbDHQjxNUQ4/TcrDnvdEtcxHbF3fdFWGCnSwaAXB6UivqfHPCGVZ
qCHh7R132yPZx5ITvEFkMlw20K6BUR7zXFVsYnp42RpnBCyO7W+xBF2M9yxiSV2l+zr0glrET2y4
3S1fdBGt+cSFqUv53qo0NBfejP8M1KVq3km+nJEYfxVfMmY8P7izr8nAc7Y4eVfqswwVsUNiKhGx
R47yAWYOsAV6b1diY5WJoCL+CEQtCBlhwfhWDUhl//sbrDxUmAAlxiKl+PMm9lAwofbcC7+jDiTp
vdDRUs2xmNomHjVEpuSHn4hGpzi6MYNCJ5MytXK/WM/lgU+vQvBj8Mm+YH6wrqdhOMA026O0mqca
bHbRbTPkwonTpy+k/nWTMrEYWeCnTlQaDfypT75CkLYkw7Ywz9XzdEwXxYoRl32kjXyPNuJ81YKV
a4ezHjeJY3xA8we/z9w8GCWU1p3kvOdf/+qxv7SiCpV/WZ+ftn5251+CK+6Ymn8V6Wueo/3EEJ/f
/kjuncgS8Vv75mxCF6BI99DOJ+vSA6mR7o+9mO2DgiTVd44A9yqMSs/WlATT8ffC2xqU6H8Y8U8J
N89fHRTFCV7DwaAbebcGTtmizZkSbZuCPM33Z7qK20rgKLBaUzgFpjvAWs/NssG6FuA5+3yiLrQ5
UeLhnRmFwFxH33MgmWzjR7Rk4aTibFJEoUAL5bKu4CjYKFoXQCOzjMNpjPUT4HBkrt6NXDYkLZmv
sIva21w7oRuTTeeP7W0qVJXof25iKESCZb6rLwxrqCHwmvSI4hLMlXziyhY4MbgU36grt9PRlSaB
PZy8LsajP+ElIpIS0LgeozBd2fGZ5NwtEE30xlUoTvllmWiQAmDRzDB9jF6lTVDf7baJFulPvxEl
sHuy659y8oafSvhb6jctXqPnyhkxyiicd0PpffR872uS27Qyv0AcHBo1bHvTL/kmxBM4wy3FKB02
Hk2DI23TBuiCUkgPGwq3mnKs3chWWkV0ydu6pamCZXtwkJEeddlxW48jGZ0/gjePhbk6ZhOll9My
oecieIbWizyCV2T74bRfqtEVDXr8wODzE17eCstG5rIoqHS0BenoaLRrH0c6A3yjZlkAT33P/x4v
qYZaguX33H/gvbYPB0zx2N2ppmqUaR0QoLA1bwZ1V+mvfX3ToRhfusQaIHu6rFIXjypmZV+dVs1b
NYVTY9kt4jQjOYesBG1FcWeoR0mEwyRJtA0APr+HaGCHRA7LL8n2mN448uGfS5XVBcGoZNeT3/aY
VzgPHoIrGHNjPmsfm8U3d+Slbszz8wOIM+LhllAeYdzLLYvKDDYX5Yq7M2pVUc/ioGe1eoN5gDI9
/gC6G5dnK8pzKP6nsqn+mAns2RtDJBf4yxNqo069rr6uiSIz5ngFooucHltvbEKaEp/ohum/2LKy
hrNCuNqppba95BJBdznivXuGCpvPZc65JTucaN9O0bfipE0XHguLcET7ETNH7c2VS25Gbk6oqzRp
lC5uyG67KC+N1Ubk3Ug6gOn+f28TPhQIdYm0s82eti+uwMYNhRaG2JHVVy1Qpr50agcfkcSOUGWN
mehoZ6YwXeAO5buND9heAmoGzflUIdICUJjVcf/pI9YJd5Y70LUto2IgXB1f/cSxGnySbngwG+cB
jalGjSiGdQRkhqVGNGjdW9GV7vtv/aEb+gnZpozxomNxFadfqnYAIs0NEEosTtVID8YMY0UY+C+e
oFfNJvlM2rviRKe1Gf6m87Ayz/T/WB0QsED6gKoR+56NfX2dv2G4zXwb8lUqk9L5H+JleMCu6gqD
yjyAn1oJ3f+KBvv3oVKnrVfhJbcvpRdc6jmkEulKGYCmEghoeuVuINIDbfssJFFSkbOng5P/5StU
AyF+tvcjGeqjYS61ie4n+j6VljRgrpD3NmFmAAQzZOEFvQ5V1npzDGLK1BytiRUdJqRFYkbsUNDm
ZoLwkRfAjN65kNdIgjfiEnGScLJVx5WJbXYKO4iQghpvuP/KaBGSXx+HaXdMwYcMHk1T8CTIBT1l
uXDGfNbp91bUNlv5uW/R+7eomr5B+1yEYWUAfl+zwbj+FGB81xa4EBl6NWwfTQDKnLHex9rDj/Eq
TWnQc3LZ4AB9v0EYgMahaSpzz9AnaiOOiZy5kbd+LQh30tIbz8tEm7YOKcXhJD1iJaxiWDtXShkn
LjUTeZ2yPWH/+9FoflZJwvWWWaJu89PvaY2jAhiF7X50YCw+Cf+VvS/P5+Rp+S5swibBuDTKVX3B
juvwh15dkA/RSvzSY9x9DbA3TVPb1iIK8JazpU1nN3A0XGImloh2vRYcWeXwc2q5O1A0mKrFlJTo
WT7pNPAv6kRdb98/uc/BY0pYLCgEPRAshq8gZ7xyogIQvcjHrmk6ucTD5L5VZTCzl2utV/yM41Fx
QawDe299MbfWktAbqGUXupijkrBqBMjS3Apjr86v6lG4GVYfgUdoGIwVZkIgp4PLe+da+QwltSWY
trilcgVox+z+zHGkOqrPQ1pcjw0vIvQtcBx2Mk9kFD6c+3hdZcRFcihZzWM6xzIg78LPl/3EKxTz
bjxn8Sjf4GYtyz5KQqAMB0dUJBNEP5S9mLkB/+BOE0fEmIa1PjkK/bqlwfvsXrS7D3Jer9lGvq4o
XAOFGJyPRR4w07ktnDoHDprL23R60BIjKxKLitGYOP0yyPjWDxhmtuRSo4JVYYbERz4UKZqMpM5n
QjewJw1QKV942MMlDE4fBAkjBor7EADtVYibAWQMaNZ1d/ZZJYQ/zAcCgKsmp8qNVrzICjEVr2rh
0KN2u6yDvwvHrunYImL1sC8W+rWxYw3ewxwq/2gAHYlmIqlZCOsceRHAw4xxVJl+5DBQhSnrDIHJ
evhH7BLPgMxQbwhqFVZ31LuG0YMGQ4r8jjz0wI0UQ3woTvcZZP57LWl/1ciN+cCs1oaK+fvOHYLq
8hMUf4c6zCaqAKg345lt+1G7P93QY5laNwSex33+1nSm+9ONdjy3xkxtQ0zGX47MATBNVtJmqxl4
LsJTC0K7FAQOc4EY/ADLMJ3qS0AwoH3Hc0Mr8PfrWu1PF5mi3LdS5KqanmQv6HhJ6XxMAwCCefRo
bV7fj+YGctb9aEDKmrGCHoohMMiIL7jyOqNkmxLq60qqZFxhMdEVKr40fBBzQkyYwx+dcR7h/Rfm
JFb9jyGs9ttOQzsz2HfnoMS4hUyzEI+ZVFmdav7WFMmXa6ap1hFwIWf8LKVgrLZ4kVc8KD3A1wMs
3gpERLJA3caCgD+CIZCCHef7E9rOr5X3yMt75NUoSMlG/iKO8r8+LQVU1s0ZyRZISCFqXWsRzhby
KiKE8rk10iisHCoS65Olp5/7pdsmFxT72xWwZfNBblsomQPf9NUWtRkG3pQK2J2ITBmJoPFmw6Ur
oscdi9GE0O0EXgWDkXxkaCgOdIf93C7kRy7IzMSIPzYDW59xLkoC+nP9jEnRvA/F9bv3bSxs0uYx
67G0MkyezBJ2hlss2GGi0azFBO9td7ZoeIvLvy9VMSWbn93lVVHfhoJwpEo0U71f0P5tkLcmRXL0
sGCFZx6Eosi2g2BQeN4WaB5psFrB7++c2z1RxahlMaopNFtyoJAOqX2c8Z04HPwpdt/vKFwRJbE8
qM9u/89MclXAn0p4lh8LTfbCOEgRDPDDIpsIUs0xVg+Tgwp4LVyw0ymTioetbRkmpkkyO+yIg+qP
adRjr8brM3V6lqYz/PjXoNmxZzWldSzmVn8AfNNzdPVBLGwvyuzk9zIsnP4Hp1EmSvcHI8MSRRFb
m2HDPQnwqE02RrU8Elv9lgcNNQKG/aNdbagBNr28U+4Bc70Xns0PF1ApbmQUwiZCAyHtAHWLYViG
uFPm36dbETU0ZGRNp+t5/JXzqsvXFxbK4LqmVxCZfUHxJ8B20qNZxaXJ4YyYqsg9RCsq727CDiY9
e7LdrG64n21lNYStpnG+eVpjzNB7xzz4dUsnSKZdAN3zKeyUe+HeEovg61g6H5/Bpj0iXGhIB2T2
5boFQTj+ilT2T7T50p3VKEY7X43tcR0YePiOztHDLgNMHbVdQMXY9rs3LdLY0vQ0zZDyazZZ28Eb
tQymxuMLExfipLDgI7PIDM3qVO1i7Pz/LmTsPxFOwTYg8AUSHnCO8QXbB4RJdnt7dPE5zd+QKuXJ
LqUZE+3HDN0Rktkxg9W7yMAlzP+OZTaRXun4Lcz3TENCnRAuhZEPvmTnOuXjg7ZlD+5PYC6/gKIu
s/h4H5tQwjoHBWPR/veunGQwc3K+q2INMDOuF9XKF0w1URQZX5A0aOWI6qAdH8B0zDwA3ZL2rR2x
5reXwycXB2j9BS1PL3feFfkjTrRbLTFLUTAlCQoly9ldt8U4CdkVa2l37LcaT1avRBOlFlA9dSta
JpXiBlHR7/aPWY8FgSCZUT3YSV19Xc2MLk8wriGj1wnaqc+6F5AJ2Xoih8xo3tRnHRu/0gcDKFZZ
2pIVFkuAHt5SlXAUats06e0SEDiaxS5Qkip21luAwWbOAJFTAdJDCronpaTg052RCrBiQu1LD8vj
rm9WxuiYr/14jNNQY/R7ITb6VSvd3ADry5qelV72HHb0rI3S9uss0fu9mzfFISOLEiR1Az4a9jGB
4rVVp+fLqy8wCWYTpM+yApn+DtuZIOZRdJQPBDwIuwJ7W042IXu0MvL0+TPJVI8YR/7yGAZf+8nm
JhnMr3qhh6f/Rl7x0ADGObHont3oEwyfGDeedroIaB+uXlv2t1CSzsXvJCShO3T8dkOTZ5i46iNh
CK/NHg1yRRfyqI8cuR6pEOD0JrSOSVbHYlW/8jwkapvCHp2JlYHMMa1eXcXjYH1nKSNMermBal50
u0LFkQLDaTBQTyvH+KagZST86mlRKWHBO6P1IJdcd+Gwzlar0mo0Mjt2udKYLsf9Vol71YqGWa+I
SBPyQzIW2WUvHCPNgSIdT174iNNP2uVVgph1CEmg8wRzHmXSULbnonLvkwzeeoulMMkvGO9TNu8q
hAWE+q/wXhouwhCWqXT6mYcJe3/wACv4b9HzxnLfKe+x2mkZGXO+V4wZE5jvUlfzAY9UxS1gSUIH
3DpXAsM5rvs/Ppk9oeX6W/6payz8YGrnbiorQt80D7fTk1Ww7rAj3I7zYxrbEvMHHOnu6U9+WEr/
vnZk2Lxz3lhKwoUVDxqzPeSPEiCFn+eApqY6Si1JdKREcAunVN8qmRqGTuvqwlHF3JX47M9MtLYR
LYXNdOCW13gEnYDDpTtzXMO/9B0qOBMetJYotY0oaInXSJcT9F/tGg63/dY2WXo/58ynyW7Ld+rL
ECJqV5xFNJLeQcxRQcD3vS1AhqmTg6DDMt1eVvj07WgZDARtSfs/4veoPtyehLJvs/z2pt+1gwZp
TyA90k8oN9rZhgrKsV4OZz3H4VaHFV5a0QfDHnYBkI9EbD/cPzvzfjG7R204ptyWoGdzqibNA4i3
TCxf5cHjWifBb4fDdshZYamFQdBRAZsmCVZQn3DBa1RxXZWdMD60luWydBPALg+Fw+Fk/W0V7T98
bP15GExqR6Lvy0K2kRXvavlJUYW0zBckfzSoF8/+0JocyQd9804d9yyv51/CAUoWjC0aDFS5efzF
lPCnoVdPOrSxayIrR/zW5IFx/MKtfFwpnhtyFHNRZNTfpwpQSUkquxlXZroCC1KnAvp9u8uxvwoZ
9M4MDrNKy56Ve5ZBidLpk6IdxJq7xEbye33VLw0d/x2A4NXumuhb4ZyFvfVIsTRPnQRhe+lpg1xM
1gz+19t6aFz1ExRD2ekTwHUwMaQ5ZUfOGewgA3ZW0+F0kA1vct8jgJwzlZohaOIjdBTp6aznZA66
OFE0Vf18nZArH5MiX8BQg2+WEbiLmNRYmJVCtNdycaYSopPLxywFhBW2g88UF2fh8iFMm5wubVZx
ubWLhMoJ1CJHfBT7zrOaTP7R73l7eT9VtNp0LPmX+xZZ8PWUmCqiDGVu+9ChrzCIIQN3ZkbPfF2T
9wptBD+nm/0vLc05sz40Yotmak8S5dCVga1EkY8ur61Gga7XYU5reIXnRp8K0jjOkCwulZZ0Wg7K
BYtp2WkGyHZuUZlx3iYiJKPnkjPHWSt8yx1klefzl8lRUIqiqzkCywKvEzaBGZ95U+K0Ncqmpaml
NDbKWRwmMsEjGqbeGCCIb2gMwr1Pd/0omobUPPJuQGB8ko4fjCcaUKnVHD5emvOK0VydEWbjzyC6
787Crw64dOd9dEJr7BFXVJMpMorwmYrKxVmQt/xgm63ffowe3yDVuS34yLEaEBAFVu6v3HU5mrK8
zYQf4Jl2wZHORfTc4opnm61IVLXLCA4lefUakPb5ee2aYEfQH/7HRzkp8JmX7uB3SLUDEuCSBNfu
5R1pacKdJ7QqY5x3tkejVOD6yPf5sdTgWUxnqA5FZH+XXPDMPyuqaS0JxIWytvAaP8ZLLxhfgDtD
YVgoFCyE4AmxT70PcCipWqp+2eEa3pKM9SPwb7hgED9EkI5h+ru/26y/AbQlYakocQuXkhS5F5v8
sO1iij49pHxT7q7k7Sra2b++4wVoSuhu/knwm1v6p8m+iIJPIHm2602PteaiG6SefpY0wpNpEw2Y
CrTaG6Jpw6HxqfzuXjOpjH8Pd94vGxb/XNtOUOmAbJtY4kBwBSkzjpU+M/vrz0HgKbxE4KOLHQvW
Dwg0PN8/rbQtJxG5LaMp9aytDRtMxvVThVouSc9fV7DGJjftyxPVpTHho2ucTukDGAmNv8ZqigP3
JFHx5EKuig4KtHHPeH977UIBuy7vHpZTZJdZiMXuNr2G0qlPj0jOD6NC/enSD/zm2uqvXZME336Z
YHR3IKoWN+zbVQny8m8Sf9T6k2X0oSgdu1esvZ8RdUBiDXhEC23MnllkiLtwP8UnVyWXmULM+lek
cvQ03ZP27P+dTbmYt0NeLqALxxAC/ncDPydnzHdpERU+Z4ca5374YHPHlxNFzZWQnz3rVEj6/tWS
a2KRm7yRVNJ5k4fhqJ6sEGTVxhpPQH1JMzjD4bZUmjnnqJEPalNSBUiZPgIgz00+a1D9a9oxj7Ee
SNyfOYXY5rqCfzT1EXpUZklU/Dy2EMB8AkV+tVluJ4FYd6Hv+MPzxpITCfIHBNSS8uLOQH8xlEuX
Fcwv4EK0F76dMrMrI9P/4FIYBpbg6fHt+vW+U95aisWj/bciZbLovPv/IFE1fz6EkrsTOFaF3/C6
ihwASQoCfBGGZXrFBuITvePL8/AfPOz3Rri3c3Nb8pYLf2kuEIyQfjwwNKiQXNbSwJVM+abxIuku
++GaumPLPFNHQT6OLlnqeFZDWe2e/znXIUNSmq8HTSKRIJLqxCbYbvXfckZEBie0jtIvoRPV4K3x
5AfW6+Cb37duE9DvB2heh1AiqBz0CCjAMeurvDtg5iBQ/YJA/7ZMs9xk/lF51s/15Aw3H7t09txC
pHj3SjK/v1eHC3HFSnDsBLfp8THayvAbA3uUWCr/3Jj5fKPTKA6PSET1zgCtHWRtaqn6EfuL1nqn
j3UyG5Z/F+1UeoeREHM/qVMewtSTWTptVZ9Yaz8KqKeK5Zh/RsFzYbFwIV3No3FFcR/8R7m+4q9l
VrKeUKDO8afbK/ysVk5mFSeWLLatNzHcNuIhcpwqPRFldQCR8kc74Fr1UIgSGJseG2IJLVw0r6YL
lBcnt2k2qZvAzZIXwfdXpWaVAEulXYS1sZrAQXvLyZetwwa5xbdkHdQJvdyMa7pZkvWUh64+S6SS
NLbZyqXq1EaZaU+zWZ/RW9zy0kEOmJ0QdwEixTZLAMhUjHhf0Qfy/sfXBwkdIyAGlIgBmnYYAjNq
6JVjTUM6vSMiTzM88oZ15+y9b8JwPnBJYE8tS+kXEGuUmCIWavQhmlS7lbXcM75M3qFBQSyYx24y
Ecq/pnf3kMou6FLuH2DQbg4+dohCxGeVaFwsSS3aMnX02AxTJmWGnnshLseLa6pD27yd30iSDyYc
LIfBiTsaXSt5LOkgxrW14IwMNM7cPCNCanzpP2SwoDwFpZs/SgEzc28gVZNYv/1nDta4Nq68cC96
Ytyr7OnN9gSilFLSXJanqjv5BMlnbwk1mdBSnoEs82zbGyrYoq3d/Yd2YgUvj3I2RNmyLvgbRnqq
wEypC4XK0s18z5jh2J7b/anOrGsPOAwT35Bej3btOgvV3qnUp0IhL1H3E3bfzB/8kIxlI0RrA8kY
2bOvTGDc0+90Trlj5o2YSSht0a5NVK5CyGllHRWgrDC/whZymyl1yh17vZV+T9H4cjaLzUI/O8S2
naR6a/qzc9gcHBvq0rkTZ635TAbafTn240xp2atJyVKHTM2GoBJ1kCHDFupS3Gq1z2rmUSlCyIqT
AkyMa1NtBK439P27Wx/qqxZqnfs5TX7EKiREBYiomAC/knm9OSQtqDRES2F+aYV3RsD2YuZ1M1D9
sD44VaA6DnpgV4pUVjFByI3g8xXYjd32gyuyvoJPLkmvRX3kdaN+E1a2hDljj6Oka7DzxF1bisat
QUFgiey9KYa39lQfgYwBinzTqlyckCB27pQUotUNVig17awl8/77yTm2Gt2r6vW1f+x6Adk1St9D
St3+AvFHzl5/25EX+o1rZFP/t+9+OW57pVKiZ/spracnYVL5ppxLKsMR6JJ9bhpChbTp2C1ja4QW
VaFpb+fQrm8iAE+8E/fA//auOHvQAsG34Fhc3oVqUt+n91yu4mf/6GOaS3YuhZRd3xcdy5/i942P
OUqVyr55mNuqEGUm4T0GryJXdjfbBPAYNqHofEbtzLurgwqHdCnl6dBZou8EyQUBi98IYnvk6toX
hNiIEDTcNaik9hsNPhqdhvoRXEtOMskCsDK/Du2B0LMfd4Cj4fDa05lX8fTlVbwndc5eIV0kbBpZ
OkJLmOenk69rTFgs+PWwQzN3RBJ9LSl8/AwtEF0CwoJYiEHZ0w7pA2IoO2g9MhZafRXl8S+TW+7y
FLplHuK4nGLHZcWlkC6tZ6WR+jKNVNi32rUQyHKYbo+xOFwHfTSWCcVE5E0t3RdFyUUa63dE1Dwq
9L9d4tbmc53MxawA2A8iuq+U3Ymyl8PoEeaS7jXQYVWXON6JAB46ayzoGSHXKYcxuhbbTuvEodTG
8byftmKqSq+ng42V7IoEtpYWzGoO6DOf8BVHKqhaW2PwZsW2EOxJKToqVUWSo4mZjcW7gTWIFpS6
VaD0R3FoQHynkCU8vtoOAOBWQTh/H4k1obeNoOrgYPZb3cXKix2DqRpD3bu6tkir1pxBlSi+FlCm
NhjESrU3dCuDU+ftnywJ9XJ1ruNmFpV7qeg+LbdgdVNVLosirYxoiXbeA7C4//ITlRwQ5jJhCYYL
sIuQMJDVGRiuyRhXT957ksnFKrbgTcesE6YrMKYEB3cJSm2vf5jyIy4mGRMRu3f+eBnu85B7td15
R4AcTEZxDE3cKHWlJ2CtV1dzG+r0V4R/9ETV5sGa/ZHT5wz/VqRzQao+WNqGBgiOXZUyFpQeNqAj
l5axXgJORSUe/Icwo0pD5yep065KCslocVHh/zqhv8FWyuXzcAvfYBvhxWIAj9m0xKVZKyKHNET7
UrndlRCh753J2m3iwCQSRU1Fz9o6tqjnqyEv47I9YFVZHvAnjRzwIR8YAtRVaWDFBqMw5uJUKQzj
HwN5D34hXr6E24hmdeFo7crco9m4TC2NKP+s1XEUbsM1ZM69RT4HLL8H/uXHwa9gqf/ccVumnesU
shUq1wf5HtaB13eahc2bfcQxw60qw/ZfTCE9qSThYl6vWYDkMbcLz6hrug8hb6QMjzfrdkyz61gX
YdjMsQ6uTJaQnZA85cKEydC1WcjIZdJXhEbUxI+d2rlUQM4srqpKIG8aFAg8uABEcqhPYCouHQDd
bhgLgSsc2yBolxKxOQY0Xb3kYknITQG10aJPGMLSROtYoMu+OzfUPVRF5Mji2ULGvDixiNT1BlCi
2UIzbCPqbdD8HRnCkFM2P2XKyGY77IFoKclqw+BDfWQuqWC808ZnkTAZAJEQ9QOE8MuQyd0ZVdqG
5cWul4XVu/ZbmFwx3VcQwAZC4sync5qMlV6lVVRT8Mr9JfQ/H2bM35WS6dpYF+L0X2yJ/uoGiYxJ
6dzQnnyWU3nYR1tt1WOg80bN2fHx0B6Cn1AtkUvCm7M/a7NW+3jqAMGulz2R4NtSIyJTaBhRRWqz
QIw5KaZtj1Y6xncLmQkuuo7knqKUv+hhE/eYsCgZ4qGE+FpnvxL/7/Rnmmeq9YQ+W+QISevVr2EZ
LYF3gP7sfxgwzt/3LUfh7V7PA3ylIJOS6OlxUtC7DKAuQUxcz5M4kP69sO1y3wUTzdCqvK9SzPZe
kBFTHL3Axok5giLaVoAvN3f/raIfJ+3iUT/bSkv5ejaWS2KFjiyf/Rcqrd17WDxibaOYgZ/DwLO3
uVXlG1HdPfQ3R/7E/+9N2lj7W46+2UZ9+DTI25kP+BCv4j5DxIZP1N35s5I5/EqmUDAtUtKmVOst
kygnHMXKN8jLZo5Qzh1DVylCPpU7sYO0T0oFPIX1Q+VSsjNXjJsqTFRvdcUi8huLANkOjU5vqRys
xzlB/2GpqVgyVg5ITJ4QVNpzhGRIBViWgKVFQqi5m5+NSienxQXLxsqNdxGFyOwtespTOqLWHFPP
Tc8wOlSixtTxfoRiIKdrPrD/cVa/sY4YZPQYtTzlKNzo3UJ8jgvddARfWMWspgSHyC0jV4xCxNl9
zcZDDrAkXXqXODVp3LbU7JMdHBUDGmyCRp/U5HEXte0kVm0MICtrq/V0IpFboGrDh6bMbz3jtlav
NZ+Z/cAA2UVHEsPESH9+zOyyFDD6RfbvovPh6MsoWIKA+RQ38rqLVepH6neuNbmit1Rzh/BefVqO
/3AkvorDNbSLoeTH5A+bhDcDDNt7LzyItGL1dfD1rVRwX+8ylou7TLwpR/L1p2auyleNMLEHpNQ6
UHrKLYevdHhLbJ/zXVLgp65qPFxe8vIPAIltMivgPfLtUmwHzlHmocoUeDhaTrOOoiujz6OZ1Cn+
rBgwauP1MutGq8rrZq7J0ATPjFO6AEGHfiGVCbaRnHWWjqk59Dmj6qfSfFACTVv56NBj1rSMZrev
DgfZSiQVoIS+w6/4sMcKv8McciuyRV/70uBGw0ij1MvOwnefVPlZWHULZLp5LRhrQQ1rBpuB+cDq
MQk8c+CaeC/XhPJPWBdEpn5Wp5HDUSfnkKhxoQ/fG7uZMa8o1QhCM2McENGWDqV/Eb2oRZyAHc4A
kZi5rBCEuVD/luri2zF3n72Booh8Q/Yc6QGQDlvN+kQnwdoqO77h3ZG0eil0+c6jl9wf9do1cDYG
RM7O8eB8Ec6pL1RLnHfOAg4UPz8HmEfaU0huqfPJB5ilxb0DKpY9qHogEDXbfHp6gyCSPAAXG7kg
vCD52JJr6HfdcyMQ8tnOV9KN38Gh/fyVPE3+uCqg34ueBTsOMVRwhd8l6PkKsmUHg9sLvE3zMpd8
RcZJhZI/5LFVqdd3lj2n7L1RPSbCIDqGxzChPTt7nkpn4E7gpjpEx8jRneOzpT8zf9AfxIyPoCGp
+jdIZg1d/LixQJA=
`protect end_protected

