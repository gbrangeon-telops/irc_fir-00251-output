

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dKfOe1Fgzj6faSFeL/IK/IGbXRIzt9OQ8DZnq2KAQwbAq1xs/txiDbhMB5jT5GTGOpfv1lX7K9mJ
mDVaIsrDmA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cmnaZ+nYMcuVxuKDdMnuchBB9inZOxPR3/E/irYVdWCPhl0UM4JuWPFoKMQnAcsoQ3vgnwO/qltn
0x8JvlvddPokOTwabXK7+R741NBmTaawP5Y3zobRhI33jusePpwNTanCHaHjalZxzALXRseOguzG
AwGiKgpBkrzwT+frUqs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sUxQSwzYYe52m4+VJThnA3rSxL81p7y01A34NmBjYzEeDRUnhBCVE2EYcZxUZHf3SzWeAqe17qZn
+OUEYPsHFdXLy5QnKWkfeT6eelEedeGrqLjWta/XE+CwvggarDRC3yCpKHD1RObvSaidPkoLOQaz
Mr6i41kRIdL7xQbC4uLsdgEZKWh/fWAVQ0EsVnkKqE8EuxaCZ+UTjEptEyr1FyibFlRQuCcRV1zc
KGcqqHxwzSvE0/TqNDvaxlN4HZAny51ra9dxL1achi8jzJgZlO8wt9Agqbh7GQueaCXon2S1zoWz
ehgKeTmxlL7ytzeVDSpaRq2XKBPlYb/82fe70w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nlRZm6Q4mAeDfFS8oXcdcSIf6QMcM0qJWL/GpoNfKsPw7GwRrG7w5Fv9DZ3ev8dGDXi3ZhhDXcQa
Irin1hT7IkRZSupkXr6uysVtJeCdG/feYDkdTZzOR87EjbK5yer40aqraNg1lVIuObcgZ8AniYE5
0hMf7gQTkG+H4+tX0yk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HiHN8/USAozrVtx8xCHzL7SU/8fs0dpiHUe+Pxq1X1HHq6PWwlbojxR2di+cVlcr3m6I0F2zjyVW
WLu1kh2il765GldD+RCzgw8JhGbJOXcaDKXvV9p6bqICOBy5WCTf6gQ/vOVRu1kKDvf68tu0aJcM
5GW26Rwq/4L2jSNVHzuzVdgC87Mdq7eVgLL1qlhKwYslU6Eg0eOYTUfGfgCo2Z6Lcfi0atBesKpT
DSbchvClt7fyjz3I+qeNhclJOyfOLBdaqFIyBSFk+zxyw4U3h7toqFVwQu8Fc+NwLgyBezl0ZUBN
S4Kep7fupBYYGAqkU2vi+UvgcgkZQxj4+5jXGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14000)
`protect data_block
DSbg0HbvWYNvOMEBsyEABfgVsdjkr3B6NzrXHddj3Db7nG/zctJzPv95tB0evll6Yvf3w3rbQRs7
g9/vVhvjkr7dkQ/TteyuKVE6NMKy+imBWP6Z1ZjUEQpRv+x5hvYFOxegPa5ZHqr8kGv8xat7jvBi
LCwcdE080MWZbOUHSJcQjOFbGM7B24pSr9iyAZy2AzubVFCUdH1aaPl4xMCmGXkhEzuSMuoTWB/l
qyp7HZml8ewO8cstcf5JjQGVc5PTsjYE848pBkvdyR7VFR9aIOoeUCgP4SG/Rntbqdprh5NwrHqQ
pbkRUpk1ygaIie2DTdjWNvesztnssL4XdEn39bCfcSwtaz+J/gtfiV3xbo/usQ40MWRL7NcPZJ/h
SQ5h+WdYlRA4gu4SyqrgzifTZ5uZWZdSz/I7DHIEqqbJJwJZGZRf4ud9PseohWwUr1jdrTRFxTcD
7FvZetuu30O5F/92pJiivGkqHSF5/Rqbc2G8/Hw9P6PbCIacwDE/BTaMi+Fet77PD9HyFPTr3BgP
sEvZvKEvMtHL0GaisW0+SmdBbCoonFCY32f3JQcvbUml1/7vNfQzoA/AYrxj35wY3BPK06flNpSE
uiXguee1bHbigvX44K/cC9Z4u770Lxls8mFrF2d+pci1Pv0aAqkyb1CAbrSGm3mtaTHeLvmzPVvp
J5d461uyszWzbbUITmgijbU4u6fF/dL8wmWh3DeudF7ADMALGwYGsI6h/qwNph32K+W34n0/yvFT
bg7CifZWiv0eaKaLKxVn+RfHgocFcFgp9QJQ0Rt2ZK+i06ui2NwWDfPQcpONiWq+QPGKERujJKni
ti+dbYqequSuTVe2GmgIS4QsjEOkge+Nci9s3+CtgwmfKFQJwi8unWCrKOCTAS4PxxiCMYXvXc74
6U7XW5fV0BWTEq8eK/K+Fa8IMgwYDW3mI0CSJZkxriPOmxN+9SGSG7dw6HWVAvQyVzZQP8KsafjW
JoN52mmpY8Rof0YWdszE/2+hqP2LPp7iAfYJ2xWIhdt41RR30clHn319fpC8xwGsLbAC2+4n1wxV
IGE/qpMMczMtBSMVE8p+KlXRyEoiHP8s7IAULtZY48FHKL72/YIiRZ08eD6UjkBbFwYyy8rqWuj6
zBHMKPIT+R+2iVwJbB3x9dQYXj9YLq6qdf0eequKqRdoLV3EfURtsgKKrJvdQrB9D2ojvMQo5KU6
Q763hu2PptKKX4p+cj8bWyMVaZC7A/1/j7MgQNwjxhpVVeDHeqAMrkNWNu44T3IMeiju4NXpDEHP
u7c4igKIUr+8Rz4Ee8pEakPK5Izmh1FwS2MVWw9X8/l1TBdPq6kptpjN3TT/HGNNNsgJ9Z6OqYek
Ub3WfbFOx0riOxhj3rojj7hLBYGX8M7lgNdyjGu5XP2IR4v3D69Wojsv83NQkn1eicNVjK7uXFdI
u5pCUCHDuX0vNTHKPhDTCJpqrfIyTuLbgaDNxeBCaIrmK4oktVWXLt+XBa2utI9UMAXQnanNguc2
ietQ5dQH3D1L1HZoyz7hSSoJFQe8dljs8BSkP01OkOT8bDfXXRZUtTi56eRzsw5xzv3bZXIZVjqy
HJgkHqPxl80DHkANwZs0RZ5t9i+EQGVT4LDaNTaIP5h11jSCV2Xx1+iMpVDRA/eRsS9WHIjJMozy
fWphlKQhgexXdleTHlxN23WOSIDaq3hTs+DotJ3n8QLuqpfUtUSKWtSixtaVe6e4BQW7/Jl9TYLP
pm7LbG2kDiTUpR9obFreg0N2Lxxi/K0AwGwYxN1zeoPyD3U+uvz/Aj7RQbYq+6frDr7Lfs2wm8+R
KXlkXr8+6ynoy/HQIFkLxytGdxLxoksSU3FZaBmSTVMdbbOoU7RKXwJWI6aCHXe6OrWhW4Kva9YK
Pv+gfitilaTjR8Q9IVTp5Ir1Y8DhEdnrtTWT5s2aEdL0kDA9TXDn77MjeY5EWxDkTApY4i7AINnz
Xeo/YemYJvdlWCTFJ2kMZPxbzq7EFyfjokTmEpSPtYTU2QxTi6jGaZCPytHl5HFXxHWUBiiY1GgE
Md7VxgV9KhCk+I0e2CV0h5A2Bd04YujHl8vKWzNY4d2Z+sGvQSgx899QQG+UoA2vCe4fOdlMUWwR
CoWX2sY7ExhsmakU2MNTJ8/T4ocJCLrcq4GQDQJRd90R9PsuqGbBWXK93sMs22V0FUIrqV4dGjt6
JiAa85vRUApuWEVStH5BfI7we6Lmzyl+39Up9KpnvxXDbuX3h8nKpq3SG5s5mT9BYgQmoAZbzGZ+
R9XMdPrYLl8QBk/y/ExJo7DsjpBtAuTgmmgBgEyzFTxAqKID8zYJ13PQ3dEJ9BjEPAh475lUV2Hr
P1dkzjvUwnHEacT6bv6geWQ/Xsl1jO21FxWnK8xybB1RChBV8yqZtlnAmpfR8Pqv1uAvFn/aSCXT
c+WnWgzHuWGYcynWsLX4W+39DgAYb0HPRLcV90pYFsUeXULhlX4ZAtgNkZbY5rHZRAjl0VVnnSdx
mVd14+q2jkQ1m6hh9KvDQlxtxEEWKq30M2SwdiO10NIMspxqq2D9TDUdUmaoItVmdGPNEx3ug5F3
FmXwO2Im2UIeXLUk3+BrvJnPpWhHbegFQnvTtiGX5ygDNJ/lVt3tBjft7Eh0U4TnWw3U/3UoYAp3
Hufev/1I96dHBmrZgTflq4HZb5JwB+kpVNLz5XxodujxM0ehutMSI2se5O3voCf+XK+FC8l8qtX5
5/GtAkjxgD6mR+PCKCp5TsdCoqfW0fOCT9VoJp76tDFMrDwOR8zLCpELqfqp6lHIs+J8V3kg6jJr
EcdqBKAsur7HBXwqSCpH2Txhcp1j7Jg4Y6JrCK0qMQFazaIbtuf6uHHVef4w6G1jLMrVDdSMb/C7
GdKrsnnGfsme+MOG5pDa63OU5OJB+m2BEAYqKXicAWCX7WsH+gde/VeT6C5C1mHHSrRykqG8qloj
BCrBrrdmVby2xseZHsClFMtqc5dnkdldmBCdsZrD4giEOjNX8uIj3g8jV0PB9f8HY3a9XAeNKAsm
12fMF+1Sx5kOBEAqnqTgJ/pbbWdFsu/pkKcRVRfNKoN5qgh1guctIMZYPBkRLzMzCc/Hav4BZryz
Zh751zjY4i/m5KL+uwoNOFsRFZNl5ETpHOjDzqFZ7dibsrNLVZqi8JamqrtVeWx9HTOAag+h2zA9
Ej2g/oLpDI7KpBzhxw9guIVOLz0FY4drqrKf6ah0Utsnd2+TobS3YTZNLG5f/9I/iZGdddArbNFm
Q6nAGD/O72EpUqx/v06wnRld6PJoif2Y/mRChBc09vG9hXJdSMw00Wc8GMZQ/AvBAF7lTECH6y/W
Jy7fCs2bE6rSMfbxJMCYiBUh8DzHQXBz8QoPW/F/tfNYBP02o9s60ZO3L4+mZVzsKIpJLfky2k5H
ahu6oxuXmG3/TAMksijfUvAfQFpi1RSJlcp8QuwPtaVQ7T/PC9KQAXz8ETPVNBSn023O8JB5+063
ygl/K9IGcD5GU5VpdQMhd3cRbhsMDlRKdJs3seuvGdPn3CXavCocUDyRc5UYUyWL8ZEgKYYFKwTz
bcuwGGweQVX7g5whw9hD0pKNS+h3ispfV3mJ/gYPuTNv1F3RIl9k5BsQ5dsHnwP9e12g0CY191qq
ERTEvr2YlgiAMIlgJSXeQ8XpkMXJ8FSLljtKMOpxEKe78sHF4Lfg2nDAj3HC2VhShTha3YaLtcHF
KHHCcHK37Q1sDohsC6Owh6tOmnfa1LDDSoh7tIlNyJkB6pe/sfLPMzVYhfGKtFHwnVvfqc91xvVT
OvGC+4THd8vxe4duBfFsZWLqBA4fLQ4LPiNJ7z3zFdlAowjCrmnMmyh23/Meh3BxBToZx9zuTAte
kNzgNE7eGJ6UPSeAlIs60jsAgTQW9xccYfJ7Kc5CiH6zKSpGTpUemzigjEQOtskJ3tpxTZwuafOC
YbdU4L3y/NY/N5EsqAIE5gLDqaH4YYSQISL9iLTNp/3Qd6NUD+kf81o+g9RiRYvjltnwN1/xy1tR
EweSTV0PI44h3YS9ZzwKNhQqjGu/+/EhXRRPIMi2GpOWysDgFaCVfGshyiCx+plxXJuI8bv8KDem
mw2i8w/Q9Yl4WBdBSRKiTJ/Cvf13oDZClIb1t6cWpcyppFZQWTDwyu53ADps20FLx+i8pyL4QRAi
Gbk6HvxL/EuDF5rAJZkp0dheQmn5IKdxyYp45/EvH41MNPlEr/djFpFqnuNxcLWBRaQuFNC/igKM
J39MZZ6wb/MZWL7EGdrGYsU9eG08zSpe6R0nTIVRus8Dx6/gHxk5z7cCvkZYwNvQK/XFPs1voCOf
sy8OPxGSlfzy0U6YsRbMF0ZcJ8ycLsVmJGUy9Cpk3+OYjiNpgvZTpGGZ69rUToFJuhRPtuujewuK
0NiLp7wXUxgQwjhwkYyYoR771zJlCFCeeXgzgTbUQlu8pFGgdiYiYcyBwJylgcH90Jv5NzGkdt2J
yzouPluomZMVVFagRGdWioO1PnCpHmUAOBdJsMLQ57Q+eCzMRMzjCEM+DYFsY/0jdtyEed7zWRhP
AkeWd1j9O23ZLs3idVq0BDsMFEOoj4n+qSXdPXYehMYfVV9PBKTK0q1ywbUu4wtiTaO/sGldLZDC
MtT3Tt7hNjbuEdp3odU03a439V6dzNtCrR/dPgZRyX7c5ubYTC5tqqwKyyBBcxtxO+eWyOM0Ozf8
nuHJ4E1QlDQDr3Gaw69cktAXlNWkdWrAZH28ECvN2z89k7np3W3eTQ66P3TNE0IDqwDZca18l8eS
c4BmkFlTVVfqLiQ+Af4lmODeUUXkCkE5adUReOiQI4FKJChGjZf95S7xoW/r0tV9WwQDlgwsaBY+
Tn+cpmEWPj8EQrw4+JpXVZOjSB8qmdJcKbbf7ZKOMDzI/lAGTEEXE42CGFRTM+rVQ1qqs8uwiekw
/6Oj3N9Ch+TiKb8/1eW3PNUwLLCQCtRe2aIw/12+gOkQrC5FfXrBsjuxExU2qF3E2qQEHliplmJY
O3L4rWtNPS5kreTxCb1IJaTwphe4YoyBAE5IHHbUCXuXRGjQ6nMAjSDBhnw+r/vwWGHzpy01o/Nb
eeBFVhbIOmO+NVtEjQB4sT0mUenRX9q6cO50WZtMTp6fwVnFh0jQ6J/1c1f7Iz0miKO6ylCVCJHF
HQ/21EOCVts+52v3lSf0s9McHZUFE02fnHblOdJSZOKUKfcIazSPbBkiotlp6siIJAALWo1GysMY
R7NXsmXppOQn/qJVcl6DuRhEgeShjgDgGO3rrEHK9pFUBK2FCC96VBKdGdvXpeRHtIONlbjU05Sf
5cPOAHcvbDA12L4zEZGEuQTGhTVHM4gVeC7xIK4QHXmR4VSSnFSsuAwdwenHLv1lMHYIolUIgOES
bYv+Jl3lGg2oUfEQKU4SIOeHE99oLRVrlCHVRdnwjzaDWZ4EYRtcnUSWFCBsF0wpKvgJMmqidMID
IZ0hP+vj+B55TI74FfHybdA6hz0Z0iJxH4CD/ZIe5yiXxxMoSbCSFS5FquiGrS1Q/sBHEw+iRQxi
H4gnGUZBA91+bOm/VHmGGhTaCiOCZ382d4TLttMwwSIwtj8yA9esIyYaEyGaiIEozwClvrLtkUjw
XVO2a4Rda9w33OEINcCm/iKtUmbSqZdsCK7+zKFV+6rVp/JJgN2R/mNOE9D0YcDlPsmChA4aFueb
uwW6Lj0GuqEYiNWCoxzXE1rm/ndoWoIcmJl3SqTsSvxHER3bEABiQSfZ3WNgIVgGn7zUhj98ncVW
M0z3cX1jBlaVHtU9YobGjlDsy73xKr0m7j2t6ji5dWMMtI1H+EBOcPH04orRSz3nq8EHxtdPxW/k
ROzB7Tr5jS7i6zdLukm8mQsNKynmdoq8POJm/CsTTgdm+5lu2Lxx0PmF1gM3vS/3V+kjHrD7TR2i
bXrB3C4xzMdKR6C5DcI0+cub3crOq/a0DHHziHNoeXE8+r8h1MUy2vWlmrFeA+IRb8ow+dc1gigR
N8h0VCn3NLZMDvTriZgGgjAGf1YR26EELLQiya2ZdxlantJC8wh0Y2SD3MiNOyivNu3gWvgjLc+0
MzzI0jCTfhmP4Xl7XU9dPYSObD3n+xxTZs8D3wJkhQSbFdATGhOBMMCVM6GfGaoYZN6PD6dfL28U
UHhfWSqii79x5G0SalQ9FcqWtW4J5P/ngTLVlcWhPZGMEnnLdTjB/G3Jtp1DXHkzgBAmHoEN6lsy
dpWlWVeHir3B1JFyBbCx7QLOdnIsdx2VsuxJYbeKWpq/AoOHr7+6jdasyxNbKQEDNTIqSZnrqhvG
BZDnn0TDkximdJmq4739Epb4Uhswq8UTRz/RWS0P/55Hk3SGB0UpFpSJlaBwvXWo9v84IUdlw/zo
qT6+wC43xIbpPiOQFgbh7QxQ623TtmU/TMuK/+8HksayH4CX/VWrm+eYXKA/MIhNNGRuyOT1UTsP
4sflOOkm2TDs6WnHk2O6KFav9sdEV0nf9MSgVsqI0QP05dR37e53ziga7938pdcPqqHuG1eHNzVs
b+zp1Q7eUlXUrNieXlHw1m4a8948ovr8HqWYYYbQaZkg8g5QhpHPkg6pgM4qF1TbpoKG9z0mA53i
diUY4OBk3qUgHVm6zmBkLXI/vVNoWS7WCAy94po6jcl0i9YNlf0+CNbh6miJEXQw3YC/kUmXS+v6
RrNaHQBNNGVpKNmC3MnBRxLVPQDTPdlSPoFX283FsCkNQ29N9ZP5z+wa66nW4uTtKV+HHs2FKgy3
zRazl3+O+eeQHFBnZLrU7ZOi+edbGhREf7JQnWUJr43et7cWA8lOdC7D1i+CbowIGgroviX3CJEr
FPuvDeSwD+OfvmfB81F5KlBpqqROUkza7GYEv+LJq0FqE9eojwcjYl6sGmeavUxJS4lqV9cWvkEj
FjEGLhX9rJT2FxJ99vEl8CAMwD8yXu0opQ7i5XqKn2n8aRu6RHSfwmyJBesfBceHgG3IoxTkVuzc
IL819X1ICyqHoxdPoq0AJ33lfmjn4mhAJCbrba6bjH5vrJlCM6fqwafT8OMI/3o10EOVRbmWQ2UX
+hfd3pyn8NjF88yvXr5Zm1FJuPizKYe9/IbjxW5nPzayKD9QqLoBGAUKpj0xET7/f1WUusc2Hitx
8C9wlbIQf43t7Y1oVCI08ygiHw+0GvYAkkoqERhtDg0nSaPfrDzgN7X/SfKBTNNmXB4f3fWqkAzR
3zSZNk5IvBa0e5qXgifZV+YE8mafJ8kBX0YyGGV91PY1bZvY/M7UlM20Dx1A4vsK1nEwsUlgtA6L
LEX8wzCcKANWJFOafmumniP8ulvx3jBrAC/d60AOwxzcHeNTdhHM/V5AIfFv29t1QBWf7DtwPytb
YbMtW/z75O4zKvkx9JO7ozvDU9SMxC2tQ5KCUxo8IeLV5DJ7oyO8EXpNXUJT4nJZKM/LpKUhQSZY
2f9Y7Xb8bnnnd81WL2Tty3SrzanfGsACNWTkds2peOjLc9EvMBzH68MYR1FTte9VdyJMrndJ03d2
ACwfeSicgJSSTZzGxTOXtksjUqIDvm0qpNGQjOvujH/5IZ900qQb36ho2oTZGfDbJx59dAVWRfGW
0eBGq3dhajv7kzmTR2NV1LLsA5/Pv7U/IRsBsMrFs5gzj+pjl3Nb2Szqkfb2OXklv7TJ0kSyjt3O
hlmXBBhIYD5GV/eHgX2+HNRsrz+wE7Syeoi+zuXzRvHWJy2DkfeO+Q3yeiGCjMWQZAZr+7HT3DnR
FPKUvseyr/GBy2FIOfIx3TIuSE+DQQ7c/4VeqkAatL5M3vaS7oS4G7GopGs23ZiyzQ0/4bspv4xq
2gsVb3H9LVhkYnW278H2/QauuB8Hzx7/nL7sENuOQ4E+GkbTECsQVnh4zi8CBHdJKPYO9lvvEytI
/AQqRSp6NCstRX+IUL3pBRxLX+xCFkoAxY/e4I2ea3ZjWn63hKsB0MPcfjwAU2NDs+QToBlW1YXj
9tAGXcaAY3AMAjQUYR5sA15txvM+au11PK6fnGrijnHKr0G2kXpFar5oCsU298aP09YWdL1uJSzU
/yKS5WjN6kevc/44t5Q5nDI5zKBcUfRq6DIY7vyyWEEn9wdtPQs9nt3szvBGFxLoblv9esjuwN+Y
7WrhYr7O+iYTnuXctIkcuXKtyBB/9TiIb9bSaNirWLD6cVKzrGoBaNkSMXfKl9cpwQq2m/JP04Gr
RcVOWuvVEm7+WDWjgQIRL0pltj5Jwc9lJHXGBu1TG2WwEql3j2X0Q9e3uShCNToG5+y1+McYmi2y
nn2eONygy1XOVo8bymZLL2MwWMIufkaimVZhX3f+lscIvXK+sAnAP7NAZU6YMHA773xSAUM80G0N
CQztWZFTuXbjlVZWJfhZNpHGwyyrkvjKxrkBEQCYHHJ0tTGyZJsxZwSHgOH0neJeIoJsfu3lJ0Ki
utx413o1oonJvQm1T/LLQALybaFNXJlct6nqQav7oGkj18CZhLgVNZMbOPE6wflcLa4PEtknN1QJ
E2kXgz5JbC040Y4fkBETPM23LTlFdAne2XFPQdiRsosE+teH6noATm3iDB/zURLybNxGTFDj/da9
BYOAL4tNketppi0croYejC2kUFco/VEmN38L+uGTyKzlVCkMnpv5SJskg14HKV7SPfhSFwHqITea
/d+gPW4zN6hPZBM/rtCSsEEqOrRq2v6WETF5f5Gf54R0A4luGdZfJquStFCeAurW5pLuOBo/qeF2
vmU3kl31INN5lMYWzVNsUowfk12ElJy0Gmhy1FW/5DPfK0F6fkijAhKMjO8igEn1g1E5bjfOs4m0
ykJbuAsvovsJWOKI43lnF2vBAUF3nYABdfnhN8R50Menog4Z5Lwes22YksXs3ZPgi727XzrYQDY3
nvS7isu4QYWgX4A/VWl5/MeVRj/3rXny8K6jGMqsjv9UQ5GmI7L5+KdyTvw0AhfaSiopbojlOoD3
lqfhl4suFpYcSR1M2gRbTSEXvSOKWyYBX4d6zF/hQe3O1wmIGPHUTDWE1qL7qWPFikOh8jv0VCAJ
d0DYQ4fnLgzZS8F+Gc2vBLwScopqHU9VRGnKNHYg2Mn/cJs2iilAJ87U6EuyBVWkzE5GOSjBWYG7
zPIJjVzSqNr7ENJdn3XFC7eJ4Rkmwp8z1sv+pHP7EnR9/6rVoSED1SGXke/JyVdrkkjxcv8fzu/6
JjWb5MMgb8GFVqoAISRpOjz6uAYKxbXgHZKcoEaYHTBF2N0Lw9MHe810tzjVGOFgTbs4DBvgxRh/
ySGQXmN5xuhK+TZt3pl5SUporCj8zNjPfHf0fa7A11iXPR5MAW+JEJ9FVU73Fo5N7k9B1vGMjvdI
ZrWgZqlszcXPQ68dNkNfofjj2dudRjHmWhSM8zu7RAD0d65H3uFz8TPkrLE49bxAADVW5PhLLA3v
sX0T/Nwo3AyaLmX8BbFZuuovPmm77efZeOr85bKibFkwQCdFb9e8WveoWKIZskxYvLul/0sqqhM2
T6gRD6wpN0YdrN+3zhOjnCkwYt+0RvOdPL2Z29uDSi0xM/zngWWE5CNx2dv8/Le1rCslFs7fRQ0F
u405Tl+KIY+AOqDiLVXCYKRWHBdq/Ue/t7j+wMlV1VrwGkc/fHxRoC1WUh/33+xgXrV4aVW+2Ir+
yDsbqa4Wh5L8Xi4Z0Q6kAVt4+KBLNKHX1qKNXvAXMdrXw5oEZKw/L96Wzyu0iukontMiPMtXpyp6
Fam2hguWBau5e5lJoq84g0IDiLx9VOtTlTVEXN4r5qbnwvE7ShLRdh7uCeCKBJR7qWR08KXazRJ7
+nhid7m5Cw7VmuaxckZnAMfdlddQazqqmtdzZg84BB6IRdbozdJVH44wBCXOsF4+mzmfXVi/vsYO
USRzi8zUenT03EH2uK4n57D5alwqtuxLczLZ/8unQl0Fy3hpSQ5mwVOr7rGaxQawJ7YKnYQK9jiE
Hj68EGcdYy1/l/sojbiYbcMyVO3BUAM3BkxTaGvjlpx71m6EEk1vbTdO3tvV2Vy3aOV5DONJ7jPP
10bMTdVgBeRDbzeF5vavSlfwuAKpg0C0pUcuqGgYnWmWLgzFro0tmDommZ7wmtF8I4Zrf0SxoPry
xyfycxvemyvFel4bSCJAUT0EymQRW7P/K5RABMtuPSXHLAxek1kRkl17MoD6vcHe//7es2TC6msq
gb2uKOxLol3VX9dS4p7Sx5UcLJXPj4mwrWETQbaHRrgAGeaE/Q2A/qy03ulrNLw4qRSuWwu3TUgg
UaEtWpL7nAjO1NTLvTmIFh75ZCIHpWxElH3S//8iTVZUobd0ETqswPODvJz9ehIPRuz26f2LcTmt
Ay8fVHUZ14XlYZGL9dBRD9XfRldUJI5Vob+yCjMQ6TxJQZECJCRbCTyEd6hEhF9cW8ONq1+ezC7y
0fYJqw8cG3a3guSQyPlSQl0RUCFYaDx8Jx9iv8k7N9TLpAobQ8kqoGXpkfGoJXM8nqvi4PIiIvBg
Xy/6uJCGbT3HaORPyq04DRW2mQ1m0EWdWk/omxr9SZCDMP+9A5kuDXdZ+8pr4kBS2AWxPTY/WJdC
ZGLDt5fwXIWmvNipqCQlnIewkdn3AHjlpcg3qPNGkRKLDB18eHKPBH7kKFW8lGWxweHtPm+JVzXI
7Ro6B6efHNrIWfFNMwXtsGMK2wuFYSPy0z/G/kZ/YVj68H/xcit870Y/tMtxA3Z1GSkzKCBPjA1Q
lPPEMjxDWIoEgH5fqxPaAkP97dUgU/Dm6o4X9L7m49W+aK3NSIvFsVoF1Oip+l2KJZ3sTLNaCtOg
0hRqOrTk0LSxbsu3yoaPgrMoUjBNrtxVhn4c7FsLOFvm5bVzZmeRyu7rIonShbgZmZ4cDJOnCpic
ShstRUPdGfA2UcKnk8k1n7nQW/pQJlupWmUnnrzIJ/ht/oXkDyimnAyMOkcKG9lvbqT0lEfc5UuA
16KOGh3HlMqvBGEzaCG6RdOHXZdn/JtXVpR+OSd55Y9wDr65Lji6M2+a76lbMJWFeC9XgXW86ttS
5v3bOaGWU3rEl7U6JxzohwcNk/btwwHjqEhQ/IiJ7ORRnuM2coxhcINvTko9jagJLDdAVQyTDPLq
2I8EnitHghbgDUGS750Rb88EFYKmKKPV/lOFDrkF4S93TFCFsAoSndZZB2nttszvIah3dhwH86ur
6UXvCLYojVbJw1b3cPSbuaTyvk0W45nEUCf5I43MQJuKzwz0G5a1GQXG17f7aQhPXAlkdRbFYN35
PbZxx9drJFWkIv/A/0/llGbJyz7kyBSqhPqaVc47TuEgVXcKM50AhAYSzX0/DBlInFQnhnxRVhHW
mlSSmfjJVjcBQa+h0LZifZNM33ayLot4aOQDwcYSSXLMmF0rXZBfQjihzGdCuDHGc5bRbgtnEJeR
V/hfZgALY8RWF8FUoKVKhys+Mdn0pDYt5F7Stu3Mk+1AJi/SoqoDvFFyz5bIE66lIiZXLidpHaBv
27n7nelWm4n6ljJaWN4I0QAxQ7LKdlARtkeVrFxeddvLlFcv+mXvoOAUrp1ZxY/pla2lhYj2psWF
5iLfjfW7/o6/xOsB81Bg/RDKd9OoCBCpZ7AO6c2Epwv7OwuHWtNjm0hLD4ebSsThkWsfdmb8dLkE
5aUyfZq4zdsKQgSgnYIYmOzasmJXiAKsnjEBmOcZQtyX2+GrQOi7D+4hlFKHdCI1ex1uueM/fLt+
OsrDEfs5hFP5Sgw2Xd/Ue1F2TMTXUO5ZqXCwPhZET5YsQZ2aio3KXBZ9JQ9NyvFBaMk8b3fdQICg
mANytf2G7niK0I61mRzpgILzwfQrT/PRKQM31sx+rMePTRT2krPGbl/8OOndQEPi2fkzPrqDM9GR
K2KRepzByBNH4E46Z2oq0yYRQTigYwvH1RFY6ISJEHUa5NGjNyyJh9wXVWzjH8RquVEFs2d+PqGm
pTi+35shp6VuaxBa8mUI2LbF2r/+ZJ3iD50y1GT5+0/2PP2uJ4x3tfYquw002KU470uWVDsnRjqm
5futIDQxAlg1UZv/re0YIzlki4pj0jnaX1gSTa77g4hfEKPy5IwDLmfHoBE4EX27LsdY1cXQedtM
BJF7q+7HMwh6ZPRcVu4jrD27dEepMkwGVXy2iLlXwuUA9zNfqsJTsqIRVp91InUkDLkFQswCKi9B
5igcUxxagoz6nn+f4zKmudrklllab4YpHlED8FM/3XHroq5j1yGjHeZA1aA/mu4ZRWBuLx5LBJOb
fgMEye8+JLlfRhy+xPyiiEuq6A76IcZfsDk+rxwgpaUo3b+g0jJwG/OJbqcUqkjmLhSt+pE/72PE
pLPBOl8zBBfvFl9Dtj0Hlm5BjF2IdbpFHIHb36ToBfEURv+yT0bvm5c386M7YP6/TT7gN2hwBeri
5H4vh76rDJMk9nwRmsfpAtQn1t/QN4qKKpPmQj/nvvX0mod8yj5qwrhD6vmEEI8fgnJHsD2MNfJy
2PkaygKpb2pm5uZ6XepGZrgQJjNLcvpE/5dDGgJ4uAccntw3zfENABbkl04vI+eJHxh5f5DGemck
0uXuDSJRLvbzoOh1kvsTCu+rqC6dmXMQVgI/ViTcrXyegJicCtMfUVx22MEIogJHqyoAoKHT3LHP
wAqwCSJff3NqoYHHJGkUAUf94B6bccOWodBA2FmEbKKFvC2sYQqzUmyL2Oj2D71G05smvg04UzmF
YqHLRrRGc/SaVlL8sv8BUZ/RnPzoe4av7zKUMrYpbejaZ/HraD0sokM4UzczqQR4N2bFLyyTDY6z
YWRAgqelPbjbOFpqfCGOfMdxgrk7/mJVVo77ZS1nhBCCDmzREbW5FVOpseuK0986E5cN6SWT0vtT
pQp3eXkB7mklxhScIvo5ZdZqpczEFQbEj1EtKyvzhXRGlwHtAGdH3QJyHIp4Y3pXIkLqC9tUYgYq
bFBpZeFcSSRCCPbHn40ww1f246iK3Bp25nWS2d29c7Yx9QV7d/6jX8oCvGJkbYKo2oW6WjkHk9sc
l6rsrRI+M0L2w6Z3jMvGGLvXr0oLh2mUZ/O5Nvrt9jlxv7i2Xe41KPogJle+udi8a0EGZl/KxVsA
BL2nvhHFPRroZqLItJDBXOKp2uy4C82177Td8QdlijiHxHG+DyAPrv8RGfZUIDII4Qm93h61vVL3
AQYo0I4LlFiEZ8e/CAsIYeC80Rf5SF5toTakFPmPMh/SJuZhV2ybPBhMksIaGW+IDFii0KCEJdql
ixstEeLJEAJssHMICmKipKr9ofVylSsVX8zdxXpBCMypu8sNpB32mVU/SYpDxxYVdCDG431myRlG
Z/TAHc7KOheXYkspASCqCbToy2FrtAzTtUY0ku/ju4dWmpSUSHjiiQ3Dx1jVt8wgHlmeIoNJ/XF+
SwVuCK+HQcrwmG6oh7BzMoXhJ3rW1k8EnPs1OY31BgdnwBqc//8KwktYIWvPrwiYjabiZi6n80vJ
z7RcL+K3ZATEyDYG1FF2E1VujqW2WTbRonFTjMV0DGY8qUNbTIJU3oeo6ETXOXvy7Da+DLnLCqAV
Dw23NrDvqkCE/IRaa2NG5vSS9V0v233qG0ah5/R9g5VuRCNbojRPM/bqfMj6oELLPveHlWlkQ+d5
fMV7U99GVkz4kyjqbyaydo+zs1UqSRn4c1qTCGfKWA4+P8/I4rm5AdzwOsjuc/9QHQUsr7KYotHK
khrCs/kLZ+w99VvGKhzek4LsQNloL4NcgUaexfe5GzBSBpSsUMMJHxJIuh8gFvz0qrqFZSOfrDWJ
K+5ef7gQ3f3hRNogUdKLWERhgRdyB6mGj0e9GWxUtH/rAbl4CXHXmvVusNztBZJOcoJL8vHVTP70
0Ze2konIVBqvjxPsobGE8UjbEdOlCkUh5jRcuiGNdQJAUYxelo9j0k/bmgIJ48g+O5MJCFjIwilj
JU4af6uDNacuuh6mKLIFIt5E23iUvx6qlc14/YqdbsapB9HpMIBUfH+VudKSfOKxdx2Prd63lu01
8V+X+/96OINYZXu8L9hNPBmAHQOpVcHsBgNNP4UE1Bwob93zuR3qxH3NuDUP4pyVLMXC8j5hn8sE
3U0m504SbLZJgJYQurd102vIOaQFpiJ9CdFXIA9ebPalG8c1nqOFK6ccmkPOMzr3yTr/UBdbccXn
tJQL1zvPZHMiusg3KipLlk2Y/MmpYb9XPXUfi8VSFhznfyGmI85cJD0FLTtTFCxubOhEyHuvXUUP
mm7K/1R27xHZrP/2rZmhzwe0somxeL8M2n4FDeNEhvCKd2H74fwS2BsZ0lIuOvieTIjZXs2nT8OS
uTSecVYRZ9rZCIPit+QJliJud4ymR55nly/v93FC4s7XkooAyFNDul5OUP/CuP9zSmuy7GkUls8G
b5OZBJoFbbX4ccFNZL/EAKoi0KA7y6HEtaQ8sRA6DFdBAd/dbDpEVU8F0TS5eoC2zQhbUwjz9+C1
kg3sW5g1/GOrTf5P092lIbCJI30sQdchsEElKM+QnPPzsiagQOPVodjrW+Nc3rEMAxM+rHTFl+K1
c/pmW2Uym4MKtIshiHk19jsCdslAyWT2a146nFx+S8vy+9BYA9vUxMO+o1fHy/wpS5JSurcJO7X8
pE33S+VwAjLmOWLA5FkHdFJTNhlot0VvXl8ssX1UKzuBf2zuTTCDjHph/TtxqgEkxFVCUI6ABzhP
atTkn5ADpkw88H7zYfUJ7jgsJQQz0Q6+0wMdrbSh6af7t0oHnzu1RZlHZjjPtiqYbbQ+BYwv/Aza
LWC4QQg+dx9d3/ibIczLVuGxzdQwbfo4DNDmk1/v019IiAzDv/qp9l82x7ZkhXUZDuXBcTMgx92U
Cq5twLqfx8Hs7Y48TPZ6EFnLifwFTYjOsrtynciJJEC/mVtRWr9PRnOlx1vTCpljUgFjqBD9Bju+
iDGEjNQ8ECvzMrnw780ss6cNIWMMBDtMNS989ZH4fEywrTUh50jvgEOUw3fEG/farNyBPE//7Bho
asoq4Drcp21F3aBfnAl8O372E8pha7ULHLK0935lDpq3wHOiv+Mcwl5Xv0yF/ihx9ac70Aqc+Ua6
HoG0vikbBJ4zLNwmLFcD+8HB3cwS3BTRqvvxUq3VvASYT7oght1cKUlU+3JVNt3uTUGbiu3szpBT
/aYR3OeJtCfTcx4H9qyawt6xLcMI31yhec8I3znp5KApe+I2nwJZFHaM+GzjgxqXkWGE+VJqZd1y
hmWu0YdxCBK0U5U9gbng80GzDWgfoBay0j3ba3rT4xUKs3C4aymuJdf4MfPpTTxnx3xRITzPeBwF
PszLLNi7YaaHh04azCHwmCFIBG6PK5KJdNE5zNwM81ycp3QLw60B9KClcve/WpNxNjJXunuGmopL
ocu3Ou5OzZFfAaWmkTQg1vrQ8Wy/w21I1rmasF8CF496gpXTbR3mXU1oZAZV1uaUPFjJR0IdlbnK
G3qvcXYcPuQnsAhhvJOui3NtgFjx/6LeSRPoBhucCKkTw/tEVc7C+FRcxyYv6+UVIE2dFlQcLfEm
mc9tX3hZnftv//9EAMsfMubrBfFZJyITEoq+PB7PLWo3XoWmBYrKro5oFLDCtN2pgQZNpHnkYxhx
Xd6yJzKuAtFK6ThqzPNp36CBwO+tBWehLDAAFDiGz8Buf7BMK0H24NVyuPN6FDt9jBTl3TEFnOeQ
Pa0Mx92DAHxRfRHXeixeY7XwdajJsQ0rF5tR1QFyslEB0FSn5KtpvD5DQUYtP5ykw2/4oN1L5h2f
RT2wrN8oRozfSypWVvQuT9UdWCMm69lZjdpoSevv3eYIRU06ZojAIfIqyshWHt7+ZLTEW8KxY6WE
/86bFngsyHz2wNghMRAYioDHFgt7afbmElfpPF1UEoElqaq+qMlJ1Z3z5uTLV5WsNYu7fv7d9vsp
HoRVSbJdXtpRsaahCVbVDyWclBXvTpcgfuDQEL1nT5j6i3vqYYCp7m3AurUVxEQrQ4MzNK4a0hMx
Tf114PWLskNBu+YjTRasp/pR6HxCHEyoFXp6PtsJSCAJ50lnhUPl8XBKXzAbgmNtO1O6Z2wCm0/T
xFO+wS1HOlyC9WzbdGM6AoVE2MQ4aKOUdt3Uk7ZJgVZK95/CDh0sS+ah3f+5CWfphcauM9pRmhXD
XOD/OvjhYU6MNkYW3XKKF096E+mCTg8RXdFqG0O2J1hFZ41yOHAXw0CxApyOSjZPOIJvp0Kkw3RD
hXiO0d3Wegi7Nb7nx74AnbE5S9XXowcUc6ICXQK+EeU+8HhKuU+SS3f4OKMCyjMvzXfF8OT3xpYW
unC+i/0mPkOZjwLxF7yNe3UDfx2rc6Ui5LDqyyo+LwwHJEdUBtpMNWDsMp+6rhRV9yLiY2ngukzD
PemYiDb6VFSZw2i5jhtzqBX24BIRsYwKuzE9cUhQOUNheYCBbq3ciBSJCTOcPskOEyGNjzFpvtC0
v/zS3S5/5Zh0ljK2xYtTBtke18ZySPDGSP8kKfcSWulH+6ZGYxio8atEjAuqs6ZnL9JbM6xPv3r0
Dx46vekfYnsj6lN9KHiumCAalHDF3SiaAnf1YypwHothcFqsU3+xVViBq3WNGGDSidztIf/07Jlt
zjMJyBwbyiwojbDvOPP/qDohZSl9WFKz8HWMDnEzv3N9Pjurw7HFt9CxjQVpR8AO+oOC4Rjr7yyx
J9uogFteE6Jo6Dj8QXD4F52XO+ArnkYV8fcYLJwrTXFrpg7wfqDvztofm0imFfLnI8DyP2zlLKnf
FGCNBiCfOy+/2sGBV3SO4NcAHdCvn5UHcuYKmC55B/wgQBshWOFZP7mVB3u2avhlOGlUtg6faHa6
d/7rEZiQdd+R5PHta/Bq1aWnhzjSMzil89sBB85TWGixjJgDze3Zwbub3+vID5H+GA78Xhag8Pfh
unKtZRSEKK/oqytvQ/jQVEDmFdpL1VHv7iy7VFj//0+14PdzKAgbmNvjnV49u1JaRcyVYK0h2DMo
+8Ik6gefPcV8iwFBYjK6Pu7D3sePJplfQlKWyE48wV3Qs1BxtNw758CMOy6fJPKecl8Z3UlMHBiM
Ei/zsdujIc+rFNk6o9GI+7GUN4VHJlI3JTuJFQaubnl2iRrAvBEamBAKMyFCCxsCKjv9/6pt0Hrb
nDO1GhBP2fq5j0FCl56TH9nd1Swj1gnQhFYqKfChWUb56A4od2mm/As0dmgjpfjiysGQAnJ+8PuG
PBAtuB7rBkNxciT9E+Qv8arutWTRUuViLcNJpG2KzoTMmTxMuYK3xxz9aFynu3fSmHECOPu84FFM
Wrivny7sZ1doaxW4ImaxmDlRWuGCu3d0aq1xxU7ATS/wyx5X35BfOmUA23Y1hWeV7DSLVsCZezU7
EeGp22AXFg659Illt/vKk1ilTlDk2deKw6b6Qosig7ug13TMvFhkcrBUZo+OAd/yB6xnh7zZstnn
RB5h6+kES4XeT2ksoWD8jqyBKD8/diwYJcHUOmZozDeCVTTa8AeSMUt9kOiLu4ews5ItGZ4SCAb8
XsI1GYu2M3Yk+VIH8hSg09k5Ex10knoioGh+mW76iOoYSlkYvVLTmPjTKcGiHnKE1QkLe5AWM88a
+LePaXeKwpMqWumMqA90jydFCqtu1bnixbbbEpxuaH8gkK4EzJfmD1woJJEaTmj1DXL9Hf2TDFMH
htJ8pk0Isb4TSWXHhlGs0JxrOc2RBuUiFVnO1K+1UfwgvY865mfQxTkfMFfUqSDhWaWy35wRCNax
d6TSKhnSqQhQ43jT7A5SA0NrXArUwJkfRt5NpuyJr+M6VcdmntveUPz7x4Y/p8Go3/RbmBFr1CFA
93dIbvg8a+Sey07WbgzK5GdUap+WUtB+AjbGYL3yImqE/GazI7WpAZR/Vv2o6As0HPqRk/mG8wLb
UumC4ctKn2NMon6XP0WIaBOuGYBddLqrrqOUKB4ZWt/MBc/SmuMKs37Ccsyd/3DATcJ3IsmXNLNe
/u3XWFlSCusRAh376C3At/b3ooknvp+3uBxuUoT0NXAGuBJTPbWoYT7Qg+qAbKu84k3d4UNVPqum
Z+mV/CvSM7janHxLydiZUfuxHufAMs2fV1bOPPvl9bWbG1j69dhnMFDBrS7LWqjBK3Csf5uryXGo
tNtKPmwmBovBhxmXm+2AAen8kXlGPzb/DCLsug6OD00sZ48iqXrudnKh5DqvJ0I9R/lfLnoiDL9O
4J+HYc83Mo4KILyzNU/jrgRERaYCsdpiwQcwfxC/0VrFsn4/aHW1MJAq5I58NqtN0q8I2yEoaBoV
KJ1TTjsPqCItIyHOkKjYFWJC/QoFX7QPVylZfhx4QipWbxUUyQ1uVVYQXNIMXHmTLsrKeLkSIa1W
C+/j+i76RF8XGzx9xhc199S6zsr8CkJ8TorEttu/kNSMn8zi4W/A19GO/42wR+FWwJvfSl2htaRy
J2ZoderZ8ZCLC1l8khkBkBBZuDDf0TXapXURwevCbiNRH92G1PjF7HlZR18dVFpc28H9exoDgXW2
P7+epWznKQwDNOXpy3QI4C/usesi38ry3sTC5kSGbHFN8qqqv3Ao1xx7H6P+KDix5xd+K3N+RDsd
6TIrDW1H87KJ5R37OiJcE34aW95fk1VPhqLwPoC5346N/HWvnx7RRuYqKwbNWHazpk9V9uJQZKXA
4epJmQckLTBTjA3JU9KJbOott9kN+2n5Am8bj823pFgNb7o=
`protect end_protected

