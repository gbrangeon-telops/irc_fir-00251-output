

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CmScm1EG7+yOvSHJHM5cOhdqnLzZOcepWxY9DkMOyN4kLbgbdLuAH/l5P4gSPyg81gBN3kT+DB4u
PBXNo4263w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fwqNpFcMm3h5oYp0iLLBA7jw3Gfbtf9OYXqaNYQK5M/u6ozJ7zqm8z/7Gi9eaTLXS/9fpHpwK0LS
QxC2diEfybnFW6aKTP/iU4AM0T8Jfwg1fYYXa19VRgeHNuXnOnQbGrbwOzyL+M1AE6VgNshYAcke
HFUgdv42HBSaLBuVCGQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D3xIUFHSYN/tuU6xykyZi+w6uytCi8PG1RRIohuMCP7mdmezS82HpITZGe26wOIBAYGliyfJF+bm
//Xu42+HAg7awD4lB8/Gfse7Vws0SwmUepHhRYxtuQx+Hau6aq1uL1eE+GMEUXgxZ2vOXH0ipYrS
hLEg3TtjTbccTVimoRhbMQB8xVTXKgd1xaluMo7+0fNF3EBfFdhrX7VNbbmxpV636ALP/wC6VRmP
XNe5xXQjiv3FP3uE/Bt2VYm+z78C9QX2joRNZHnjI1wlv+JUs+OBnQx0uieg97dZpGTJDWS/ROJD
yUMDQnx8oeo5Aftp86QvBAbfaqE5X6J2q/lamw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WD1VRz/pLvBXDYk7fWsqqk9E+EKCxbcP63KaJV1ph2old7nkwo7SBQkXHtT+4KqXUeTJT6DxPa8j
tS5RCAcDnWldx37xHa9SUujjT7DruuKAJejsjhxtSfv6A/nEW4C6nOkCH10rAuqtBTv7SUZEElTR
EXiyr/yJfBZig+juuEc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TO3nxTWXykAydBE8oLE1lWHpTk01Db/e9HeGVQPfEOiTpRxWensjccZLTO1P6wLTocrobkWdnzeG
BxBt7prIiPwnDDfhHMe/xea/ckp4CqeBr0GVOckjbocHEF60X3dEzewbdNfFWYT0uATcWRkKB+5o
X3VNEsL1+rzFW3yXd3oxwxLZl2hrAEzHGv2AAZZgDP43u0eLOoQsuloFBUh5XzvTCc38IZkfTB7l
fBrAnLiMxoJyYNeps3ny9evx3MIX3RbK+6dmn9Aviq++SNxcoN8Y4/1btHsL6F9ez079jTeANSEU
ZvBBfKlGq2n/FXU3NGHAnGxirPn//Y4kyfC2Kg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10960)
`protect data_block
/4IlhF42XiO1NEwbmk8ZtKQ57ykOhO3Jjv/6peCmi/KlbUsmhseI7C5ivERF1BfY+mhohBVcOKdX
bJo7oXDldLaUGJXpaNzhcLzZIjPfH3masl+/OnsWeRoJvjZIGseFfEAgKSmdMWmnYI9x3kU+ntBY
TidqpxBKf+uZiDPecIa8+1KsqwffPgqmmzq5PSgZVhcoGpS/1nhw6qVEO9WyWbJYRwJu/jEo0xy/
t/PWZNZEctnwk3ppDRZGmoiZ4Yxt9ZIMaD+cDKoK8VgM4pkPs0EA8r/mTnhMue7e4Javen5gPByX
bGFzOHdan/fRsJSeDVaCsgoy0z6hslKlzAVB8KTHVmJjSgKmq5DSIrI5HXKXZBC+Uxbdi1Qi6rJS
fmz2AJSCy/X+BJcLy8jTIeiqYvC8c9s0SbhV+fa17jK13UYvdyqZOVHUOi1qM1uN2ya70GHqs9wO
4dtRFINVceBCvtYsPrsGPZWVGD5eswi7Hssw19og/3nPpZqrYdsWDVr3ZQU20u5s99jSQbdyuOUE
KJqVSmFjlIqqMCISoApOWsJk89tWItTSWFr4ms2Kb1XQf0WyJlMuUtw1O8ygPCIf/Be4bnO8pZPO
fJ3zDntT/npV9Y3XmuL9eRc1B5hHxa60j5vP7/Gla60ygU4pcUbrsyS/zfZghiJrYkPUdif+yFEB
n9xNTWQXNEwWq2LWm5mWmFzVgqntuBTf+frpFcEvchSudYdIH5KCT2W3LASAyckO5BDB4wEAne/i
HJIvAricB8w2LVOPwRytS/A0yaR/PqLuYo8NzydIugyBgzFLu0C9GqapKu8b4mIQMrfvFWGCsBDR
KOwCaG4/iQmjniVhYZwUKyOl9eA5gXcGSYDafqq2OKQWzuxRPPyv5Iy687lMV9VUuIeu2Kjw44Ve
IfvRB/uw6gQyn5bqnoO+923MHblLRq3bR1NQtioldwdi0acDRvUWFevxB6IYPzXK3J2lMXmQgycI
1+dmiLCbycGCdve3/O8igZJHi2+rRBTo3PKxc3i1vBB4/UlYDq6qAZ7/ZgWfarWLVBq8vnvO4lhI
mg1LchXIE2AJTw7P89EqjcBUjmGMX0+m/WF8/CFRtZ49WBvioLxwCJdX2SXjaE0EbE8FiA+yDS76
7oY8siEhSsfaA9HLvQaC2NkkFRVa46tub+ir9oNmUMduMeWn0HZ9L20C9o9iVrYPtuHg3ZvP15QD
1b5zIU6JasRTLfk95YmM08RnaSHOX+oLPFRDusgnE4V30M7Pqo8PQuu6JErlZttBnUiGmbgb3ozq
QPP/7iCk3AKQMbAJG6djJynLmpoCN15rP0Q89V61Fu5LIDgCXNVDbw1o8SLQoPEVd8rS5q4NU95q
mtq5OGwIUu03+bmruab7/Bs6uiPWyAfij91Me1UeN4Fc+Wkw9yCKcjdaZ8u5QGyHjnDdfu/zbKhG
a6MhqIek1dWfAx/wvhCPsRhC35fQTM6I/gMVBUB64zw2k5nmSrD3/E1vwZ71MezTFMKP45RU6VdK
QRaAKyJCIbXbfv42HPVDpFHQZL0YTKwxV3cNNYDQt/QeSStSSeec00wZR1WWoeCWTcUrZSh5uUeH
YHXQ/D6FXl4n8ktfeaGwjbWccV9afDGgxlhzTIDqQarxSxNXPWu4s9vhIfLna6ii+eo6smzRMHTU
DGCbJYDnVUfmreq2eqTC042cobNZh/VTJArYUcKgvV0zv17x4sEj2P3Wny5HvmVN3sps2Sk81JX0
TsldbqtKNshFaJNl4+twuvvzSUvno/DyTNLy3AKhio9vDarhOyXUYFBkl4IHrXWiKDQ9lLGihKBv
rcIGjbNO1vU7dJcshO7a9BTQAnhkgF7i/zr/oQCn4BPaAIjC/axdFZdHjC9J0qAdgomvHrquf81P
lDTNKih2PefEw38Kuc3w5nvf78/wZYLHiAS4P/VxpcbnwyS5giyhMpAcJ3RgbVVSzFYyeniz/cy1
0iQPR5TcfShq1fPFXCbugVrzfrtJ7Ur+C9rfex7yld90znbRJ4jMwRQlkihK4QfgDBl7Mm1IRzUB
tD95Ulw8yh6rVO43jnN6qTlVLRKoNH7k6B4Cvfj3TiTcEdYfezmvHCqG4dHfx+woYuryijVMfPBS
D5OmW9+rOp4P2exmjBuZNQzMTsZI0Q91cxKM8oP3NT+rr1AV2kk/3Mgd1vOtih/qeVPqELboauvn
mjFhjb2r9+KCkTHvHMCMFqu6gC27MyfHsBNzma+pO0tOUOfxW7E04hg6ihFGgDp08BcCAYQwRQ+P
IargenJvZE8a8kJAeLjaW0Qts44+IqF0ChnLHPJWBmiSKrXtToSpqLYxcdpzgEFL7EkYhDXu27Pb
kACYYh2D3QN6mRzQSZD/V/foIp1AK090sbm31OpHAW0iGWX+CYCaAGfrC61aqF4sysLW9OZC4EsO
hjPSIfKQeJEL6gSzKloY/RiME+jl4ra39tGxnZUIuJo9zcvMzac1ttxfVW8GDpJIxdU9ZUeFlZY0
eiRkuRyZlbK+l87JRVu5sTlLzVP7sOJ3bCmfeuwPaC3NAYjgILYkr6+XYgUtzLqKGyaCBoxeAc6s
fzZgPeAj2oES5cNWeo/g4xbVEacXTIuHA5BdIor60MUFgvelNIsEu/dEiv2L/5eaWwR9wFtL7evk
KPLVg4P+2eVp4DZD6z6EYJJiQ3KXIr7c8VJUMS4BK6YM0n9s29OBvGD4tKnoaPxaPUcpRLYt2blu
+OeLVNhjSdXKH04ChpSbAjwDIh1bBkg1xbiEjNWiz3tEkomSiS/F600qTa5sOlKTTkYUhwkzVPRe
UnaEKXICjTYr9hBVETGAbK4UbEFuUNheqq0tWkWjnUNQjhnJ/sl6GvTNq5ZTa5oz1PTtUUGal5dt
E65jYAS8XMXnS/pDP83XPI+GJpt43dsgdpnIbGLy+zQAwCee0cfVFD14Ec0iSCXuxhGB1S/dbAvi
buptbmRHm+Hnzv55/ZdbSDl18zoqZPSIKWxAdDgBzB6Bu5djpDWWcqrGuKYn8RhHZz7/7+XH6Py6
kqM2HAjWpEui8fb6j+gO2ZdZe55EsEDTvyXFdQnCmmOYMXLJ6vSV4SnTIiXovWDYljfL56xT+e/O
jy6eqdqKl8IvmFpA0CJ2a6RJc1uX5MGT93yYtURmqxQL+Fr2pKE8R1RzzuqgH329zc62aMhQLpaj
k6X4PGTCBs/2RtDo6WZWN2X+jpqSD8yCcKX8h6tUnDHWo3kCU6SJT8fpN0tzMi7/de3/ibMgAzzH
jnaa7Il2Fk2S0vqUM8QGiqkiE8fhbPtOhSB7XrhaZ7lm/4xukpSbWDmMPrKqeD2JqDgEmv0DERka
TkRvRYuEMk/18wZ9AYCYtM/bveK6TRcUA6im70KoHT+nLud0De9gxGEFQjcxRP40w0kVWBFpim4T
XKaSl38O1HJscoz2pxWGs8KOMy3bSyFeW1gCyugljrqXR2jspSCrXyKzrvOZyu8sh2CxFyKGnvET
XpK0mP6/bbEyAgueqvEw+CJCPQew+gPm/1iHPWZTzon5lBJTNPIGQFridok2g3rfE6x6AWgSqQXE
9WBscg7lJ8hsbeMKIea92IcxzzE6hVhTYxhPOkIT+OLw48BjGWi7Ve+UjHEjQOJTxCNyO/YoBMVx
ZktGF4+66uUdEA4Gfh9SLMbkR9nXNU0mikgVlxhdwAxLK/Z2eoHhpU6xr93KycGHhE5LYkt7cd0A
9BkMQNp3myQoWaLgNjQ2pbE4zUINAhdrRUrcaJisgutkGRm3lOqqfAf9EWBXkQ2CiGcBh7FXZA0H
rbPGfqx1zWQiiU1NGS6/IUmiyaGIDQY2NPUeeTIO4YfgqUK/9JYCfCTfN18XgLz2I945HgxIIzs9
tP0GrDxGTUZ5wtPTK1Ct193AIBOf74Oji+Zb+leiYiE7elrNqZ0qDqoCuIo1uqT3XUGMUJlzGWwQ
qYM50NNKhx38G7+c3SjTjPmytfMU4hm+55Exs+c0qr1qEy0HdvVk72W3DWC5s7yuoLL1kOUSRhIh
erYrM+6vAcm2+MvbuPfvWBtfvY5wHCoZ9AgIuiwSxRYIzRLZ0b46C0PLIDz8T0IhHz/5RORpaUDm
WPjkJ941TQ8dS4gDJiHt00z6R9Tf2IFjBgWRJavYTByzTL5F53TIhuAjygMtuXPn1AGm7Eig91lz
dZYOl310zZp/+K/yNl5Q2VTjKrW4pJ14KtSeo56eA7+qGk0p+c9jODLGcj07EOUQ23bt4c9tVKKV
GGJNhyyQcpxFvaVq01HHSA43Zjb9mW2DQoF7mH2SZuOUD11nIls5Gs0mUp+FnfCvBbB7kcQS7vcF
cvptTcDXPrBZoQqZh6Ik08kgdfWSXApxuqOSUXceuL72BRoQF42dgcSoyfCv/o9hic6wC728XQW3
3mQXskC7/5YXu3sXAO8Di9T9838xlj7r0uDQivX5Cow0L4zZpv3AuACb7SBgbASmNGtaDDLfNApL
yySgxgCXMNQhBRRc8K7DYVXDnoMS6WzrTrfxcqK6GBqiB74ZJbOUd3B/bS53Cnkg0DmLW6dTYCPH
/Bo8uQUIkYeOuXgNLophkZ+kFOeiMw8QBVBON50QcWQYPskGDmVm9LEg0BVpky/4jh1lNHZRwVN4
Kj0vB0foBo//Lr5RnhBDJjp5JFpRdcmgcxDoGg1vUHlaFKOG/OF6XHMUOSq1X9igM+1ZlcpFRyYQ
sr8kASall+b0HUZeOnxC/ptXZ/TwmViURnxNmweGgiNfOmZAzaObBz5s8OalWFNSVr5ALO1aivUu
BNhMyQ4X38J6sOCKhj4q/BMjjxIGpNJQRrsig2kuhL/vw7X1XcuFDS3oarAUDPJK5JWfl8wIed6n
VrCdhYn62VpJ5p5DSqa3/SDbV3YksdZH4nWgLxdyuDauZ9RJRUTSyhHIvyyWGma26OssRp3qtuHT
uU+/UC84qc5yjMAkVIhiIKm5XF1BTYIEUSPitM7zh1Anl6Ew7LYV1+ZEAg9Q399HErwIveUHerPd
6gpAtA2dcYklOnElFZwiGvULthnYQh8XMmkD503Urg7h7uBW+b1IFdBCmzny2BYhi4zkXKRAVJ0w
yFepvI5w9Njux2K7C0Z8/dvSicCP8TlWYpTOs8/Eh5/NqdFdlw4hYnREWizCV2QBIpBJs2aOaeg2
lg4VF+jFhPKoaFqCbyIgeAqOmVmH4zvJknRs3DmEjurEGFa+sNSS9mhSR3u8q/j5pcuz6mTrFS69
XGF6bEhuwhdAWCXKRDekkJy2BA/ZWvYjIyD1zEF3pgtud2rwNQaxychQt48RYpzKqCEDSS1VgUNC
nIE3nFK5FV5Ddrt4OisfgkyTnIxwixEFcDDCYDiLI2kSZSK6d+1CYr1s7c+tf+hdfXxz0ctsCivs
FSC0cB/fiF/MRfSNq61NJIPDfAhi6Fg70NjG5vIJBkcLE3LoTdFrH3IEA6WpmgY6zVeCxZIin44D
bSJvdZrA1EqtzLfC9Y4qN9KJiEHvJFDGUi7YF2mlRfnI0X4H+GCCNvHeVukwQHE/OTPlxSXnxNh6
QOIZHBHrlc6dawOEt6D/EioEGRS7N8A5A0UB6LyrHQKW9LblrIHLVFCd5MQ6F4ugJ68mpKrfcAlE
+b1XaEnmjuTdnLR+ZP13ULltTuCtInDeG6WenbKU1KRPLV9OhJPeI5FQsu5EhQh5/jVuhNqc/PRB
NI4oVL6ig1tQodWIFZlM8/DdwMDoWxGw/r60cBp2vC6OaYoFjoKuXg5H6y4A8GKTsEpUIBgHrVbK
ZHXsl13VnW2gCoZKRn28xPQbtgSOKFW3o7kY7POU03/jIHjUSMuUunKVmZUi+O4Bhsm2kDL2vAQf
ZbKrqoD09qTIhCtR/3UWIrmfVAcbFjZ3XgBPVq5kUKeEUv5hxgKf9NzotX93WJ7HOl5mfzKoa5/B
P5iMQ9lOzzwfkDPXFgJAlIlmp+gMHdODLL50sS1D8prmDxckNlXFXhs+2Wcb9BCsxJgXQkat8OWs
jq7ZFgsp0MPBYolVwL6TMk6UWtELJ5R0CWTaLyYriXWIfPr8m2H3d2F8Jxxrixq1LcyzXERlfMii
Hivq/SfXJLnHETO35UVSFNyZTDnA7iDkyKzNL14CGKOuxJKJEFIep3fPGuFvqYR9X7gXFo1NJhKe
nVsQyoWOIadHCmMEt3BrwigdXDUBKa+I4jquNyDq8rRHhyJEiVYcVI1hSWDudQSyU1hoaT5miTcj
IPyn+ZyhJ7pPPIIMRGuZ/R1T4BFrUG4dhyqfGeUY00clY1STj1UXjCQc9xL3N/XmaCArxKutBCYY
iVtR8jc7ypn+UHt4mz1JofVwyELXDqg/ElWLXVez3VkjbgPg+8VPHwBKX1ka0PoQlBLW8aQ0cqiI
4VZF/QnNn6RdzZPwMZXpc9E4jCQwtMxIvhSqTNTvHXNR+HqMe2CDr5GDfsffuloceQRK5UMy72Ct
9l2dvy2y/vqb9zeanzyMefZ/DVV+h6M7JaetH5+OM4hogbAyKwMQx5cVmcjk4HeoXXCI+bI26icP
9ktBvmNOUuN1sYeSmhERlFfoG4//BIfRuATE4cwheWXWpbkdYpS38RYmG9GpTLkyNcrKnU522ryD
635hoKl/S6bhaWRsPb804NoQkFgLUxkkIAXv202a5M4N784fjMKauPMP+BAD2+hdxs0sQIg6Vmo+
ZRmumeDfrujwjbsbE3rL7yiRBHuO8NozaQxpPwmKYV3Ic85l2odxSQ0t7Sbd+Rawss995/zXm9DZ
dwqhfGb9c16VNERa7rGytrrz86+OUyfqwqdI1W8hW8iGApsA8yI2VRYX2d5J+Fzk5rYhJ1bQOtIV
4YCAvF7puCppswXrreysnxh6mn9MTMQB8w0xgSUGvXTmjpAMPIr3bTtPCLD9fycXpvv9SwlQMB8r
SKeoctX6rvK3cK5/05AOUjodWabBAEfNHIBnC7tHI3PBo9ekxJ3R1dWdzpcJGZezMMuzfqemwDGL
8/uFfQI4zFM6FVm2yBT/nRaYsNf9He0kvZeS3ZoZCstbmMFEo8w2Iv6ypIGrP1DYt+sHd9UsRatE
c9Mg57jMaYQhMftBW9vmgLRC7XEm3UBYQt05Qy80yz+5m9heA0fYSkdyusI59l4Ok9PCZ0yD/6a5
uE7mHMOwTFxoqolceggfRb7WKXYWx1Q24cDOvMh5he7Bo+aPW8C/gDmow1HtAIQnbdMa/UEOkJ3t
mnUGiypC8MkHgt3zBGXuNM9UvYg4kvbFqctWu/fjgCJy5FV+UKeqNN7WRGHQnGrdUlsWWY7OFHlx
qP5BNNdS/rhcpai/OpV5WUHZ6R4aHrwX/AtJVmnk2SwnlllrwcP0+Qjsfyblvk0InvDQzDcLMlh9
aumXTLtiXJavghJJaRIDsk7olg5qOYiTeFw7LX9fIlRPBl+Uhi0aDnvijXPbOBqMtbK4RNgiycT7
CYLVxwZFNsmfSGH+jbdcVsfFPfY2MOb04DVx86UXvN3D/956AF5alNgZkdLcJ6Fk/QUWVJS01o4D
ilQM/ZCfJqz5SFv/1sloN5+6QlnGlYfpMP3w3QbuoSSTtmUxKNs2XwvrZTh+isWFBIW5XW+jIW6i
KvS4/DSnEa92PuXpuS7I90Er3QuRSnuvzwYq9UR33df0gCibN2lcqMatLO6lqvNqPxiIDBL2wtOa
neQI2Ag6T5x+necr0zXqS3l2s7PPFTZCLctXGXdnHZs7gDPAGDWXbK+kXqeppX6bUztDgB/fJ5bZ
e1QU+ClJbf4ks2A74/ZsifZm4jkfLz7Rok42TvXI9j1DhgfaK5vWhjA2UYUc/z7gdAX8poe1Nl0h
ENfVCnn+aQPwoZXm3e7UsEeVAhTJBNOh4Og9PJOl/gnTBT7xx+8UWPs5BoqH02O8Qn9G5L3fKApl
iPzeLOIfbBJHa1roeNaoqYPwnBp2LWM9UzfejJxVATkILU6ElT28m6kg6fgKhpcReA4kFZlJRijL
qM2Jv4AO8FQB1A/Rc7HkgClBdVzYpTTsrwUtUVgpKM/4P1GzT+HAQpVOsfYL+oopAdGhCK4xIy2R
5I3QkiW3k1fiMDRFKUFGSIS4mFK+Uz2xJ2mCJohP9AoqI5uTP/k4Ng6Py6s4H5owndn0U25ReAgW
SXN3YmXHtXw9NE68RZ/SMqU0Pb/VlvqRgOxwALKO+mJfqRVxHHQpHzLCHPtOK8eyDW6rhGEe8tYq
xE0Yl6jXKjlvDpG5emrwa8wfpWwR0SUJ4gE+uwvQ2WUNGlkEP4iBWHvvHv/9/Z8d1Mvyk5377fAE
5ZUIsvNePiiqNlXHXlTl6vsg2435aO8qC5zM6UzhhEXOCn2CqWiHaUmjZrFAF1cXWoJ3cduzTP6F
5x53Z2Jv6458H0lzjNtSYTM/n2YT0FK3TJ03OMazALEH/OCxSVs3j+G/AzwoQ5TS632wlroKOMhb
nfKbCW52QBAfjxbBdhvhCiR/rGwOUnPCTaJP59uFkE4RuKVrOdEfMtPLltn/8JQ2SMN4SpArYv7v
ee7Q+cPx9TmmQxQc94zI4nbktlN1svNQ1Bga3q10nIVLVgT7XPL4FKdA8gApvlpFv5sMNlGUysk1
a2L/H40axmbr7OElqSZo7P00DA3uOX8Eyw+SdUfHebqFlv6v14KpvCQhPHr1jDDbKWxkGDQEiynW
GWJl9emZShF9o6GqISaLjUrQ0IPAvGGZZIPy3LwEEBDYpF+E2hl0pIaqTqkuYUkbNZ7Ztekk/2Dj
FIyYu9hWxNhvQVlamj+JOUxZWvlMm/pE3Yd4QshNuenQJzqkIyvlLaYekGue9BxO2D/dSsTeXGFe
/LWuINogVO3a0RDHcnjppJyrhxtR/72WKjKUrRMtQESdhqyW9aK0vobTRA3oOHq3mkRU9SYpnlBY
pAXZbFuYoe1vTL7WoEynzIQCaiyPSTc9owHuK2/AuMwBhz3asVmrz0qwo8Vz077c2b2Eur7VEAhU
zKjnrktg+tzNJZ/5y2OhuUS4Q44wue2Sqh8dq1slk4dKFer1tk/ffg9ItaGGoQZheWDNr5RSrvw8
kp+nMfnh3+mdrjAwDKtS8+Gg+MzDaAf1nHiTKrbgb4Jss0fI51hB/i0tCsesAcgswjcvgMVKit8L
8hPWLFcod9mf4O/OI7THzl5ZJyy49VtWNIJXJvTsSaZ3Znb6gvhHaQmcuzmCIqjCubspztpoq/Gr
G2CDNtQGE4cQJJW6K3EbIp0tgkerj0CAr0s3Up2o4ex5nYcDnv/K1prOZZ+FgPF3fG23TY+cuXkx
NIj7XIt+/CfZ6ys6602QdkT0fTJAUUZyEmzat8IiT7R4kORcvl2LTWnnYWMlrWHwDNQdS8HvPREm
pjz5ICg9w2hWuCq5fIwYYJ2bvvez3OFZJkiwf2P7wpAMFvCvlha9QY+QDFgFby3PiNsTcAl12cKM
cHcj9aiawtP6GGZ2FraeAs4nKoSoDaSf2SVQEg8KpU0OPqvO7DNAy4urY5OtdAWeNircivWfAFgs
FftSbVBlzw1rd8Ln5bYwpykOOOSmoGdjBFiQFuf8MLoVRpdfVwQCPo8gL8H+f/UpIk8iMahP1m9I
fFQkwu/n9G1/kBXibrO3RLy4bIkXiPXDlssCW/ANeSgNiBl80hHWF48L8lmqQZIIWONXiqh0MTx3
qQwpXsQ62yRMHZmshos0P/qmdpLfiZf1GOjMMmvU0yNsM2C4I2eoLL2THzHiIZjne8udFu5J7OXH
Vh4CZK7QDYT1wkvaFR6BpIKS5dDohX2kag5qtcXcJyBCEBu5Hpa0GnGcVPnuUbneC8ikTm/FykaR
2su1i9ABuVfXQEbmmOlTZsDB7jLcnELJxrSQN3wnhuF4+cb3/GSEFMtw/ZNRy/6TDo1M+V41zgqe
tSJDlOUyIzLGk9B9JyDXwEnaimK46NEJUuwcH38WTh26FTf84VSNo0MKKBiV7ITinrA1/tgKnd9u
WmTH5my9Ms9X89DaOIZvMx5eQs6SzGzdqoBvlJq0HAdVrAHouEQLHZzPW4iSGR2SDmRVwqGCTc7n
82zGVHID2cTaz3jLOycsaSzVgG84x8b4rfzmhWNPnJ78+AP9gbulbl18Y04Dh1l4JihWcdfeRsv9
YeltVMbzl2O01DOrjig/R9SmHjr/mZr7E+47VuBm9ypxvOv6Y+ing+0WL35ctsGj+Yk3LbQd+4lv
tLJyre7perDLyRut6XbG+O+xpDCPlbuyuIi9qkVxsrO2WDkv+682LsQAR2O6sJ1AOc6xAVUKjCJH
S9DP/NP6RXcDLGGinTs9U2fVH8tpqiYx3lrfx/rADRW7E6LKc5mGjm1iDeroACerYEh2XMOgVRqc
8MOn7HaYC1BB7F6sMXlFoXCD6vn0yKQrXjvjaaUvfw1d7TI2jW6WavONj7jav5Iw4sHoriPVBZiU
PyCUcTsSzzqsBY1DjGiRzgWMX3QP6SSPkULQmECb+QkM94tJFMbpm6B5Y/XH9+5rNEDOTQO+ChSD
EW2FZVDGckMVss/+TsqxuPKldixdEkX4mKbOypvjnT2w+uvcQUMiSmJB0nd8R3GzS6xHqVWI6PC0
RSZWgFljBPGgDCWRjIEskd7/mL4s7JHDA1ETvGb0TZf0WGnK7GxPYYChoH0tNqvs01vdXaXiRj5C
Iz9SCaMZwH6Zg2RkCmht/GGdYhorPkqbUTofzk/jjsCL+U/43b7hZIM96GmLgrUM79CuvT+P9G7u
4gLt55gKNHN+gW7/Sm3wq2kE31enSSh8zrv9XWDWnSBygHN41lWsrM0yykvSpv6v/Bl+3zYzZZW9
hZOkwW3CYLvDzVWGqAc5V2OADZZQZnQ8463FyUlRm34s3yOCVVvJxhQefs8yUzhd6vIasPnpisNr
AS0HDl69ev59FlugLouwkl/yhXdYp7yt39BHahKf/rRx7mpQstH/6MWZ5wn23iLxQfjSynRgdTdW
iGYt9yFbhBF5HhUDJM73Z2DMhsN88t3k3Pd45wAtJRZ1vP4H6lgEW3pGjhHzSXlnXfy/sXo9LitJ
81twonKMqSL4o5MWRHh9hligN0Nwa0dLIRyePqefzs1+BCQFsK/9sHRmEvXf1Y3f8vvgGCH/J09Z
AEdCrsTLoyxaJRcUOr4Qiq9OPK5Fr5kr8YTD/uf/CWOQsXDtS9VXsePtEYoj6FJl3SkZuUZBC7hZ
s7CkspPddONacBNGQIFUDUWhH7NfaguO3vo26gbLGyQOqPLoUVxAkoE9AGtrOgw9Zl3+qcrAP2gV
l2Ub6e9JOjEsqQcTNibybl7/MnVWrn5z2JVYP2eaC5wtKUBMgpGXm8/pPcexwUnvffKBx95gg52V
M1FSk31MYVrcRMTbD7xraEUschWIZWR7F2meOc1k9g/xfCl5+qpemmRgG813Gd1+YD/EAQUJ82zV
Zi2LhuT/gWulBvRt35HHapSngSFl0aDQFY7ecrQTXAj5C9IJzLGgi9IyzAVMgNriHF9qYl1dXcnG
Xumgqly+Oobfs5vsxkx9zWJIP7y+sCCKUnavUvd9HI8OVzWPTjOwIRz95kpLyPaARFcUWS3HeK2d
dxtGxzKeCIWzyOWJkZ5za3wL3kD663ngncG2PgdDocZHF3toph713bbrB9qFl7HNXpXe0NCU2ORU
2/Dkbu6Bgt75kpafLW8rq7ddjrOvlT9KS2maxtTvvj3xd2SvTvMgc8Z07qI6F/OwspYrZyBmZCYt
JORuPvRi8Z5hoAvGiy8vNlCWI5csVUY2d2m88KiBLz0NwynsrdQdEwxAnM5bAUFWB3BIA109bBcg
qbmoMCxTdbtmv3SLvYY1H2sDrGmzVTMqS4+uWmY8GvqM6yKxdnL6SyyRpkIfRqRwig/231b2tp1Q
DgPqMzvv8jVTRIbw/nLVHaF/tQsKW3xFCg48SGoZLfjs7yYyUOnPE00uINPYAdpyj6nwhFVhYA7n
HFXgM1Y45cUHO1ewymebWkxumm0QFCAtTR/xTL0GW9X17+fMzv7XaR5kVrmH6d+skxs81TusE58d
RwBYeMaAmxrfmAfV6X/TU7Bk2nt0Zy45qZKUIilefXPUWgcuMFdhkVPqmIRFpfOsB8Ksh2hWxl5T
+sLc3f4DJIrJtD+J8LPKc5zvBZRBxecFPWmtBRcyzYbdoClHlndAQAl547t1KQOFeQ8QdwH98Yrv
R6aZnNSUFSxeg0YZa2XnzJ/gJ2/Wv3LDz0AHGKkZxtxgMSV4Bm4Mk3QMpBAm5DRy+vcz6Dg65bMH
Nb5nHHAt71DY6kSu4M/BZi45HVehXw2pDpjrl8hR0fFtep8GdZ1cEJo+PP4yw+8Kb2Eo8egTVnng
4Pg7Gk2lStyzT0EXkW3tVwuRkVONHPysEV2jq/zovF8TUmocKQB/pThk3XKVtVowGhASFGSVDGWd
1mrpWKEIvmMLTuICneZLmbn2M42wXv4bFZ89e6p5s5FWr6j13BvGWPj7GkUzRl9T6P7xoGmQvR1N
RMwnU9dFGpf83FSbsD/liCCtEOwJC7n02J07Salio3jkgV3C/YNeh1pcgxFv37W2GncYU0LZm87R
08nk1Gyh2sJiVAQ0ler6/YcqsJRWv8dL3Ro2ZnRf/jBRJZVGxnQnavqTxp7Sz2TA6+nTQaC6aJMT
5a0VH5//+sMHWvRQ6EJe0AX0cV6vhZ/87nx1aKQw1SzbNhkttIhWPO6suYxeYp+UsD+fILfwrzRJ
k/j25N+QGLkGgoI3LIdoW3hyba5E7Ru3u6AmgRsjufHjNul5e/MB8a0fNf9kaRsf++WJvxAsQPqE
CCxV3ULcvPQiD32AAnwMFfQrtuk9HVvq8f6ugZhEYPIfYdlFbh0wB/ZCy8QA/PQydIC6bcHuWjTL
8SSLDcm1VpEc5MzlBYG8cm68nT/CtTyck2iKxwtsv7dzwgbFZz64iWr6IrUXnNwkh3kTRK8ATST8
E+IZn172wcqlNPmwlacNBxivm9d54rC9KMgjCmqFV68h5JltF5LEhQMe9VtGmdeNZ6cbmG2STEDi
EgyepTz2Kal/kmo4gmOIQ9igZsgZRY+OUO7Q2jKE2RFLccIi3sWrC334qcI306hAUm4ho0HNhC4s
KmCIbM7mDLMaR7f5WWd1viDyKGrtJs7FlT9ftK/gyNfJ2eQp4Em7CtgNlkMLBPTKfrbiEWxvu301
jGUXVDDgRpJ6L9PzGNeIsIHqkhU0NzDtccBE3hPeYQ9/g5dS57haOmdNge1GSBxcnQoXYbxqRYXn
iIsZer2SUEX98w210VDUne/KA0qkaw2e1tbKc5gIyqUa1SWhRmWUB7IAk1OIa9Wxd8tW+A8ZammU
S7M4SSncHV4QXM9zXOyaHSpPiXzsdjC4jSBQQFvQhSk7P05lzj54vznWuougPQfZCbIZJYDKTdAl
wRZvU+ecdY2p7Y26bEFFMSVwQqUdpCe/V03rwQruRVSvnuhlwwbd5K3EY+xZc7tIq1dyPPd3t/9g
X+lWPfT5GFaW8y0BWeJnjy4EiQpgpc3YOBMNF2hPtvxp/Xdt9isvPU0aOVDaGCqu9e69BXwHriUW
/YM6Fb+Lpf2jyBXvfRyKsJkxzEYj+rsORsS3i5BTUhhd0YxRcNK6ebOGn2edTahiQGmcqor1Aesu
/4M5SnURnKFsy2VR6eMudqmZ1Li6NQWIXSNsOiwCtyvOS3HpbE4B+5E5S6cltvz9BthsuvotsIyq
jveU8+dggRulhiTLLtxu7qfx2FdFshNXvphEJYefPbS0tvY1QY9N4jVwue8iVuHFSh2126bOyLBJ
XiA41d3s/VBfv6rMpWLPDaaT+s8YedXASt/at4dEM9m+q2PcGKT8x2KwysYGumbkcuJj3ki6XN0L
K931LypfptDjNfFMu9I8N4s28JxS7+joDseXHqBCs7/VJ2X0gFZ4V7luHv1iUeZA5efGJVQt7dzh
v6vEOBRPt65WWhEf3FHJ5wl2iyBfAu3+xqbBINlAcIW3kUeujSFvojBvptR7jAQhh6uCCvBwLnvB
GyQGK+i0HV/uVcGo46CNHWBHXRbS4u58hHR6HwWuT0Q6P41VjLHKu1Io6Xhpq4L9Uml4O33pvVIO
Nubj5V8x9juNTvPxB++JeSQZOvNJo+lhmunG/p49PdqFP76dSaRa62+32tZxFCZbGM/gJOgpoWhl
5ZGu6wmsCLXrYozHwJAM59XwReV8vIBQuljGiS40/MU3EqbsICQp61sFquPynDCv+W2AQtkMWFSq
xUztC/+jU6DdebYAhB7kODR31dfZb0qjQdMZEJfnZEWLALt5ReKqEXbqd3dby8vON+lifzvNpwVH
5cMhkYJuWTurCrS6VzxeqFRe8bezVTaTMWxv2m5RVSXO3A73gOqk7XU/J76HikkrwFEb/lDodpdE
SYwCUM6w0N4XsDSAf7n3aJyrVLuLv2gqBVl/jJ9m6fW5oaESDHvU2502sGBpgAZH2khTy9Zz+EPP
59n9Rvisn0x7n8aJa2+RLXYMyRsKHyzu3YpS30m+2psOsWOhFZDzxwvWgJBbch2C/Uq3YimyqdTw
jrt0mIRDu5usIUFE8Vwdiww7jTXBCuX7UDHdeFYuvsWRhJ4SV5TRr8v4TNZ25di7e0Q2Dxagxcc1
e5bPxnDkpvWrVatrPT1YSQ==
`protect end_protected

