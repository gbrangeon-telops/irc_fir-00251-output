

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hezhI5arYh5Ll2LsYr9SKRVb8M09iAN2m4JSbciXeqmprOA6kAYKyNVYZrZl+7uJ9rCbSy2t8SS7
C18wuehlMQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iG3qoWxeKUs22C9+IygRgNw/Ob9GNJdHtLxrQAtYdMzP86eceFi53EP4Epvud6QFqZ+YCcJAJz6X
BiP6+zFZ6SCjFFuXw9pefFKNSIH8+q7UF5dPb1d06lbHzIZD+3mRDkhnSZjrqT/zLAUZb/IQ1Lbm
Z5oVMb2d2CoW5etMngE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lCcH3M3hshWBn3vT8V7Ds2ckpLb00IXg/NREvwDTgQ0x1n/TYrAfJvH7lJwH3QNYGbvde2S4oTtp
dxVz5eb3NKybz4CG1wYBC2N8cyfQblBGlezgCm3PFTB/fb7+0CJP6o+JNkedc2s49uA9zPZB2axM
QOZ+WiL1UDOqHRt1CYUPiwYxRC9z2R+kY3HwbNnbrtScHXOfjyqwc/ifFZR8DvMU1CEJYRjuFvoW
cH+V2gM6YyOHMcuZuaYjA16MxseT+50plqCZJKvjkYTDhSYcuZeDAun28dPbdfRu3AO52/Kq9gTu
MLy1G+7O2B+746vqe0NC8W62Tyb+rHxVnOWRgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NvvNy4fG+VCfM9NYumsm2clZ8IZDrJQ3Wi+cnwU6WbSkr/joDlB0ZRXsdo0mhVbkhlHdY0OhRpkR
3RYDWBuljULA6BTyF1sag+KB46HFjV7grhZmVLUbBkCWRKYz0xq7bDcNxf7s4evpI4rWpbAGWyJ9
TlfOT5npzM2PM090g2k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KN7EzciqITw/PNwj48fL1Z5o1AjZa3hMKXx25N37JjIMxkR/++b3PX0LoYvLH1v4MmFRO2F2HE6o
+A9StU1NJwej2oLxLD63NMJa+VjJBFCfkNayO25s8BHSFsZkhjc8mIC5S+PHU5t+p8zDOXzJvXOx
j/qM+zNzxFnZOpagckJWraMSJbbFjRIGq2RuUI6DTykdz7949XyxajpE+pE2TrgIaNudJhMJkV8s
PmKxeai9osJTVlAQyTdS+HOwcKIcXexlGTP+JSkiagntbBuHEhDR83LTtvkaJx0GY9b8oHB0RXsI
Jp2E0CkC4MgVpkaduxkwBZ7NjlyO6dFeIGiehA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35376)
`protect data_block
W1UDJwQjrfzo4Xsd2fxXVGU4CQC+uQddqtK6s5kSm7RIpCiPgIgW19xyKx8WN01XOHcT7cGdz1lq
ZFmFXG6lj8WTBP0v0p485MhsIs20+Ypcy/lhtRMak2nZ/swh7gGBpYayTrfc7vh4SnTxzor7CrRn
HZhdSG+IMpPTNW4Yp0MONqLo0ixNkHs9u6/EZbfHV2m3ysfP7fgvbC4ldYcZxs5Cbx+qzMcd1Vhy
5VF8AFU+8ly5niVdV0UcySOQiQyKZxuUTl1f3t5YO0SkT1m6Wv3iZuRvT/IWjL+jjVUx8ZrPQGqW
EgT20SK1/LeiTRVfGEp3i4QYm4gMulSWl65yVYKt8nmowMR8eiiUM5gjFEtFkxgWhOS0qn0Y7d7G
nTSteXiEzpPUBgJ4x8srkP1+1lYDgsbJkEf7FXOxyYNpBsM/dksdgLHJGx+VrOIupj6AZ/4jRUJF
ttNKTP3B68tJwmBxUhU9n29CK2T03xIvejGpCWWx+MgMWofEU0z79Zkyg51TsnHJpfnLl40vV/GF
1W52mgBwHHb1nPkzA6ZoeK9JfL81PZKYJcpmE6b2G2QnChmXkQZZry/KcB6HGZ10jmJTj0+hmKcl
TbVcNIgX4SMZxXTYJorgNVuNbTTIN2IFqV7MqhPVjxGNuF2XIEUooXe+vVU1j7WxxdiV/MS9eTNS
23sdDhsX8zbxTo7Hx6Ic2HXc2fIrv4GabqtccoaWUaTOcLBNIIQbpk2VHFOxHKlRwbBfHgqJRmpy
wKt90qoTomcjE+GeY5aMx8lOgMI7mfcUbEEnuv4kq/JYzhjXRxG3jXjZW5O8yn+aUuPMhQK2qKmM
9HgDvVnRqDEPVVQTZ9Wy++0OvHVXxrOC8yFyA5HGLYccVho7tKH+rC47s18TvMGaIuenfCmiUrs8
CQsj1M7gvYU7txiaNWzQEZMISIiiKn8SDh/zbh/eI61Ienm9Z1EXKbjThz8DwMg084bdSsE1wrEE
OVuONxGisb07teRLT/WD2sD1S4pFLZsBe1SAdpWTJX9DpjgDvB419i5pPkobNka+zoB49jXMGujM
cMrWZ3saWEOvFNVduy2Ec6fB3+BtsUPyuG5EccVUy+3/ivjOKHSyIe7/FjZ7b5LNjNjTckkeMQJ9
sSelhw3SjMGmh+oX/kRMzvfE/ovGeK+anQafSuTPCHk9vuo3V/wP9jgRjTp8rWwVVj195EUju4f0
ZmWg0xyWyrJjW955MKQuh8eRyka0fpkIad87Wx9stv32vszLgLatTZk0no2g4FTy9i7qEV0ZThQN
Un1fdsxi5SHE+jDnP7gyrArG88RypD8FUoGwtw0ljjsWPJeALQlZ8TZs2wboJBPI1C1Tos0liQow
iDBok4WyqX3w1MgjxQq/o/M0m6hXFAN8bZ0vAmlXA/fV9tBP0c3+STaLBV+NwOjQFNwHFGHVKptp
zihF3NWyitBQzZ+zpYZcicoAileWu2AOz95uFMvCNya2ZHqoTvZzXU5fZmhR2nVPxwN8ycM+CV3B
FqBILZfvJBHE7vqEY50hvp4U9SGJ9xqs4L1ubJLn0HZwoWKs1pBAzX7YqFPYkuwi3VImA5Dio6X+
dXMppsjwH0ObhPvHn9QsqncxL41ULT4oRA26Ha3okwG7Z0ywZ9zfEx7LgMH0DX+KvBcBhXxzmUq/
Tj+TpQe1sEqIinx1T/9Cg7c3clzXWcPisLy7ONAeSsYKFTfaS0EkwFMd/PUywg2ls7xYQbvth+c/
M3ZCpH/YttPp1JvX93DDDIDgOpRRzTKaGUEZUkHFpDNQtWYEQoYwLDfVV4RCGX1S/SxwYgt2yJ0E
on/6PjPD/B4ZjaPCoHnZEOt1G8IH8kqtTvugzYwxBBBAQ+8QrubI0DciKPrDoh8+LS0CQM8ixaU3
BsfwKkTcVpBqGA72IbJvrRe7tefAiirW236dmm70++qPUTtuvSBj5sTDsC/mKB+0rutDW91mRBHe
GQpZZ+sTYpuJRtIWiTK8Ntpk4RHdjkAAwR2072fCxo+VS/Hx7dASzVVCjFaH2we7R9HX9P4z+vqU
dhA/NyILfN35jObNBA5SiHfwrI2ujYTxDnscmbQ7+wFvaO+myO03ykR3tj+3bswgCIHeIR5y+uy6
R41bE7pTTirOmaD8G6kBkjdi5o7+c+9zfNHCzlYv+DrjtgfVp+anrGzMNYAEYdispESMO/vZAE2Q
x8Tud9RZxllcfWGHhVl/z+XCLakoq/qRGCeWk9WEBtgmemL8+ilrsWW8p93JzpS9YQQIIVgjueX/
CtJY69MCU3uOmjTLiJCtdDGmqrxmSjBEfm9v+a8BSBnnvqBj9X8AC3l+m5ytGY++Sb+K4xzXEN07
B1X9Zdt3hH0QwqA2F0RogcTUe4dd/J/ii9T0Qbb2k6+H2BqrFTcmN1VqgylWuMvVQ5LX/9fBGGTD
J9XyQdYi41DhKxmqdw8E6gvosuFl/Pv1VUhpyH/znubQo43ersYI4DdeN1TxFGDH5INFwzG6qkKe
FpKx87kP/0tfTmY3/tpN4tJHSAQCIdIY5Yrn+PbHZ5UlC++cUEyXRj0Z50AGBcSmxUa25VvfQY6t
NfU2xniFNhcBXH1+Uha52YfxNY8GQyTQx/yXZIVGY5h+92ASnXjGiL95ZfHkb7It6Xt59rWJvq7A
VZAmPEux/y0+grBEA7zyIg57Z+wXpbfYKe2o6G5hIBF7edBmnU4+7G8a+dptpJFY/ghMKGXcpEZY
Z0CJAq9ErtgLc1lA7Y2DoFMZh99MqVO7Ip7uClgGZIkAp+v0uCUqGFxW7HvpTmJP9uGiGFIsA3w2
d+1BnNpYSSwf8yNk/IXr2fwQ4HbOND4T2rXtfaC0As7rh/FDAi5t5CreF/HWdH61/OfBOnxppRZE
6Uo3PW1ki6GbcOvYwYwl0OcPkv2oRZ8Fx37XLbbNraWffFiOhRbkb5oJ5ViLvvVUSgRBunffWNfw
PY3mQaRprK0PwYKhgClkgkgxZP01i3KQYdpsihL8b10v1rNU+pD9YhnTngyzoo7BrzYPPc5zXq9/
4pSYOkrWzuc/ywgg2sYTrmBuGGrxWvmTg02edqdVDH2QK2uovOEf9IG0EKvnOoI7Y9GWnwBs/t7+
64KBqLmMEikjsIfSVCU4T/kXLeDnmDCnBVWc1PPK+K2y18dRmy4uzquqCXVLNzhThczs6PJWXPPw
yjV2IYA2dvOocf3NXqOgrYwXHEx8wrs9f79RfWK+DGXiEHMJAIUyU92PUJQwjbL9N/eeWe3eGS64
Ker8T8RiyzLrewfubnl4CYvhr37MIIdmfslGrUiUYaghNvFEI33f1wc4PuwcZv0Y+5+YBefzhl9P
D6ZBSQb0My3hLSYC0PR3FnxbIqyq0WdJ+YkSNANpsVngNvblxZJ7mIAapXP+KGV/XFRBj7T2xQBO
+In1DqE87LpcIJoq8s9KX6MvYEGOOoAC6iTjsAJnUY+JiATgqdha7F3AO2Gk9ezG6O9CfcqqruE5
OOZceibVezNiekg3U6KAhWQ+YqYrSe+Gu//L+gZCVOPPc9WiP+xNYgYIYk1AvrI/rumyBWkN21CL
RzMzRjAOxg31Rry+SM9yFwp3NBdQDPIBTc98aamsmYMcHnauGJNfE2PXgaBWkW/FDm+uMcbF1cx0
UdBlDoZ8PvEVWipdovfQbbwa7BcDerNTf3daTRXTITW/GWAfNiFdSQzvACR2PxwbYs4JBn0zSuTo
nnPuh4+EjAMPteeanGDkg3h24OjyHZwJ4z6VojbgR+85jfSCGrwhFU0YvH0YcWGiqJMVm0nMa13C
wFekErgW0hEHylm7r131AWm9PyO3vSbyocHCvS75jqoa1rsz2PnNWjq2VGqTMoQqlVap9G8QT1dd
7j8r4VRH7M1uaNeFRzLkFkwylH0W9wb3MMF7/SAhyts8cqkr++hj18j2qZGibB6XDrpoMoiwrJO4
AJHNTMhoIiJCXTi6Pvqoy0+N2r7UPYfYxYKvLaDkMzrSe983FgE8vYQPmWqVrVu/P+GVJDI7dnbu
U+d+jaC2IVE60GQ+cHzxVZcn9dXA2D/aa3nR3ESks04EbfTDVF5K3YdoxN7ErekHpCuDn9jU3Tw9
w37KCHRdlxeeEMK0j0zuQ+a9N3NXDLczxINBGQDCmiiV/2dXUQEvVAGgli3SCx9MLP+7VxTED2uI
NdwnDPHNCK13y+uNp3lr/JF5voGu8Ue+zOg7Gz4mxZy8Y6oUD38y0dBBlCF8K8VYqZ8KVnQUcbJs
OCrvqx0JcQqNaM8OV9qk8ArAIEy44Gzw4LPpIZ1E/lqcXFnVbMJGbVagsJDYx8tOgyYfvIGakWA9
uG30SfNadNhl/D958NlPpxO9PzpUrIjwKBXz1ASO9gt23uas/I2rPqpjB5XAttbJyM9jW3H7qsS7
1WynXfqy/kOPLPU7SeSMj0C092AKBhzKkKKLkA+OxMj7SRsRb7bySpHkdPrwthGMl85+azb+EywI
6IpiOLy6Ati/BIXLI3l+pAYLMlXqrYwhmfu+8q/rrgCylFQSTGKBnGgB4UUcSHV0amKxOy3I0SfR
5Ak3aq7zHYkHyDymIFTZPkQbBXYKW1L57FwsmmvygJgJh7HFeg+9joL8QKgdghMvXX8ZoeLZEkI6
c8uLnrNkDv7X6LHJuTOqmWmY9qPcT0/qLqYzi/8j0Cb4EIPD6YlVIknjfGRvXaYL5NFu/8OFRZGd
y+DC1JU61jcSinYB3TsoZPSuUWMAvRqjzlqSUPPh/IXcx5SMLCY5nKlMoaMFrDJNIROUfjHbEDf8
XRGlikV6wbsNiGLZhEHvXE3Ha1dqVZ16EUTyPIv61c5zKrdefLTzZLQQ1vAnuToiR4C7f8yWmIeX
IqRdxxkGpHKARehBSNQoo+KbymR65du4/hc3tRTeS87tDhL6XNUMMhaVBS443ofO4m33N3sYb4Je
CtKT4+6l0ebtTVNYsfx6w5tcovQobywtluQq4KWMYpH76LY4/nytwYt2OrUSvrOLVFHavmTVpk5l
RvW5Zkc9ZYvEc3j20fTC9Esuo6P2kRWqGaSTrWvo7MSKSYrvG5cqBibyRSaOFYgG176Uw7GGAHpR
8E4TPVE1Bspdt6cxnJKVwgJiUnYAD9JB7w6HhAXECRVa+yiMH8pvJd60APQg9uT/O4/G0DUrZ/Qe
86tASz6bG9hRG4rID0zFuAtfwnxTo/Fe33SrtfqfC4+7j0FXo/XhTlhpfmqMaoQRB/Bhpp+rVsyY
btQc8MM3fOWqjssvS0z6Rc0ElGZ1segmRV3PuENMu5Ezdt57hlyPi4ulScm0PbBKbdP3GLNOjo6U
SDaBl9DA0a+qe9NGYmSimXchG/P2KBPJKvoxFyNopdW7eWBOOhPbyfvZazQvPnrv7mHkVGGlIKYR
unJv+DZ1DP8MRap/ClOujy0ck4aRjrNSa2yW6ghmxuJI03VSKFQPiIIda5qRuuMvDx/DJudS7L4M
IoCAH253EAtqPaHUni7G2MI0HMDNrfpqB+8FFJ2h7E/RsojHuuZ5St/BqHxYhqHab2VhfBAyFGQR
PI5BaqdyNgLSHA5mHm5y3Mivm1oHkLJbFdruTTnPpzVhdV3YqNmktLHuOVu+S/fPbb4wK5/tnEzD
/PHSu/DhVaVKOpvBZHcuMGl6+xa4qvandJrHTldt6feqggb9U8hYxwIJl0KshE8qZ9Rp9+VEzf0X
isuPuwno2XuyinQG4yjnlQ5B4LPhm8Q7NbLKeMz12HfUr+M9JafQ2y7X4tIT9jKQO4u9aKUiKr9F
N8ls1XUPP9grulkIqglJWit+HfloS2pNkBiuNaMKzHrg1/oDTQ1Yy6fIEOlHh0yL5UdlX5FaMBsu
HzQUuAc71u/cPY7eVwVAHTwgSGfSZShW/E5QKWBpbMTZmq8JobL9oQweQjlWpJfs19sS3h6eksog
g7p2jUo4ClxgR3oHk9oeQvssnE+jgVs/7+7uihCoYiqk/6phTWs2sp5a6KHMqWE6NaTEiAMZilma
hx6R/phyq0nLpl9aNjz+SBB0Zv1U7uz4t2NpcPIMp/ukil3ybH9zcjQ6NDP73iKopT/vtLsgVj1g
eIH0tJsYSJDijm36JHYYmfjtKEsXS0+z19Y74j9zJCkszMOGjtQ6HDUt4crikdCH30hM3NvVAeN0
TiQlrNNP6hjqTqRLx/CUjMFVP0QXHxQZ7kjPKWz3Oa+QczIT9Jz8b+tXH8meoUZTg5rndrHD2Gh4
DdfFYs6nQ9s0qmeLkr/OGJJ1kSoMmtTMYgQLGRBUiHMVZ6AnB4BGI4acZXB8rDth5QYJbaZVeYum
PkbAWMeqLtwivlTVesZnp7j9Evh4zzx9ss3yBpXAkDDyK+xzH4LgYpSpNKyKr2l53XhTC+PIAIBj
WWY1UZeFOBt1YPMKR1hlZmjWxnTIMLTxZmg6EfQ7k4+ZKMBvkK6rh4+qPZGVtSQ7oHUq7qD3Ngmi
RzjtMA+tVirx7f1qxXDWU30mCyy4P5JQeP03gJ8mMzQsXHIp8C3vaixZNl0UPRWeEYgbxPU8W0nz
V0fdrXQIP/Tw/VU6f+RZiiybJ3PbUmeGO0JceUPZaieV12gEpVxiz1IXAF+g/BeLz9zICBBK/izY
NAwl8+ahkMAsGlmFuPbTzcA5w8CgpCMQGt9Ciqas/tInKyqqZnW+5icMDersrXT+lMElr/ErNvO4
qUes+Wc0Ky5fdJSfpjl13HAkcw6JT9P/s27cN2tvkkEUo0GYSQAkEvOD6VEKzCn4H0rSRkR/DfWF
/YfrXhQ3+G8yWsKdop0+k1dRIoutiXQH2twKehOhtOowIiB70R80bfrvsgNpYhPQK5g+a623VwMb
OFhpga6iC0LR1ojxYE6Ez2sHDbgh3qrpFXFgSAxOaEo9iboGP+WPg9ivIy5+ufQconrqJrVAQwS+
sRtq9BQynVJtTgsuRqQDEwl/O36w4PFOtfat0Wvu/EcpbfOXBaYmfxttpCGNBPBdSf/NU6kQas6p
DBdA+KnZHny03QC7OwfS9Km8hNjcVQhr4rWnyik0j8CpfPzbKrS+/Q/uNLuDwI0v62YelmGItEHJ
MNLir/QOwmp8ejUr3vBgl4dEcgmN97UX21xooZsc4nsCX6o8/XgyC98M0tPvBfJEgkllSPd2oqyr
gGC9QXXEIWdaT4eWuHbNgzSqTrlM0qrLXB6O2Vk4yPrO/iqK+SGNR3qDSte4aWlR2+oCuPDGTW6b
ZBLtiQDIZJd7ePQ2stIqy4T4Xn3Z8J5rlQnkO0DR6Ydm4V4En9PFnGFn+t6m7qk/UaC7xSkb/tmM
vSTRG8vcQjG0VR3/ErSBiVDe/Vym1YnVe1V4zVTV7eySXuwhxD2e1cKNE+/j3MqQKT9pfc4/0EJu
Y9teiZdXqBIltUnJQ6eYmwNjj0ezeXJQ2Xns9GZYreAEUEdXKVfu0E0yxCrEEB1dmxQZD8hAaR3e
fnhpdNNOZ5ZfNYzQlxXPGi+6nq8YMaAntHx45tHBYZIHNAWLvKQN4FgYliuH/E4wvGPOqaz40rip
LSpf21k28yduYB4wQm4hllYxoQEnWf7mlnSnR5Ri+h07uKRXur/L7ZEPAdtjmdFBQH6/I3uD2CKO
pOayvFw33WteHy2Sx8g4d1GvS3yvH/9aYvoAo8oVj/yW1xkPS/uu1U38VJvyxReOz/gXI64QRvur
jm6xmN/43n+zuj9VUtL4qdMsxbtke2KQ2ygQFbgraHJ2bjuUg4b2GxgmtMUaN4O1LLcBNyulBa+8
zNLpiYS8+iWpEuKnSTMRevHOwKgT/JJYsA9qR33JOE34BL58+dzQVEGnLm/KD0GKPYoVxOSwoeNR
lrCqr04lnSB296l3BtFYva7drmYFJuFIb4BhRpB59WMkmXEAltT5/3uso379C6KYKiTt8aO8bbej
kJq92eYy7THbeS3mpewxmAuh5BhAfGBG2VyyGBuHpRvagBDT7KinrmDSeYMf5sqhB1ZaMTi5WZ1Y
e9aCFo4I7p9Z5LVtaQTfwsRWB83OfqD9c+iRrNXHebeIdIBH5E+F1XrN+usiUm98NlWMU4Q3GnB+
24paoV4bPIxWwWvsWBYvolCPx8TEDN1MnuNM1iC8Lw7xVHsAchmpiuP9++9lzfKY8EGFiv83ui0G
BRwiWXTpZGGYDstfa9Q8vPEBBDBNDynrHaX1OSrsRWfPegiy6g4Hu16WUfUA/kE0tn11w+H0hCXw
m0OWpI0VQrddEUphlDKDtzRCBo6XFqsLdWkxwnUjrzXvcxNnHJwfZJ1SXaUicejt3kWj3VY4X0uQ
EsdkUdRAKd1J+NFgWsolXXEdMKlsIY3vYzP/Xhc03mpLioDerUgUyAySNyxXnV4qTmhgSy/+OmMP
lq+Fn5kKQu7yseoqh35n8+WVzxCcyObnSv+U4GXgsD83X4/P/bZ5BR/iHMY89Gkp9UyBZuDirmpR
nMX0LaNqHphS7WTSiraMxBPQqonSYOOMLnBT+7G85Dn1fefS2yu4M39VHEedPiFsX1oYW2eV4MyX
eI/vHbe26zm824IaS/GsdVieBNQIUVwI5J4lzdyLt9lxQy+mUr4RpxVe3Hz7942UEXXLHFm3zyef
AIV1FLO4H404tmdxLS5c4zBmrv8nuxKxmQv7KW9GNSjHY1dUGk+3+Op9ybmv5tCiwr1XkFW7kM/z
lgpUP/mc6KjTjo6n4JV3EQPzoBRAXPPwi+0iP14PI9tsFcO1prwlT/PyYfc2O9X+D2NAbfq5bDiY
zo7W9ctEokhts9dIg7QXJ4/BOIqWfA+meGU6oAtXmTG7D+LkT2bqDXzGbTcoPYsUpGUr0W6I7Djg
QS8lmv7LZoHB1+AGXgbXupPQ7p675ggVUDWI1/5GuTNJF68QBh0Dy3nTXEVjxGleSeQGISnHaWBX
pOcL1DuWXwYTu8stljw3zau1aBMMAaji5b5qL4/meT6Qh7IcWA8j6zF03Lf98Kakyb03FWrPl5Ci
Kul5/y9NZF99PHzM+K+dlTfa/F8wINmZlUHUKU/HMuL8IkMdTz4UUh0+FSusQEb4l8ihfBSQydpH
lZlfwHw4rc+tGxnpsBjdeZJfnTz9Q4IUdw9kTX/8s4ZPbrqx/5uYjhLKNWOlEAZG8tM0xSZw+ss/
FY4NHMijZi027SjQsnDFDYt+b2hD9l866ZceIzYKM5oVDY5aRyEX2carGV50MamYaQk5UtNzg4Z1
oMClPdfnap4yO3ittrbOqkYUNum1m3pbycXrwyJNY8uGN/gVNY+XZYLldszSUrknT/uQACEY0X22
1d8hZu2rHPIqs1rnsaxMwOosZ8RzqJ4QfLRqSGDLW0D2Rggq79KnNnOBxQ45lrKJDRm/P59oEyxx
1J3ux4z3r7RlNZYIY5FHEIoaIp5qnaEpyeikA+mtAIVVNK8oabYMr1/18tiIoJToLYCfX0GjjS5+
fnsSgMhLnxRUAeYC2hqLd1uv0GLpo89p4nAgkjc6kxHxapNzyXa5a3zsmhhR4dIeLJVBhGUDa6Ty
VrwtJkN8zbXrKFNWQXDtyJo1X+hF2y1kmt8GtkuQYfE6zXYM8gT4wtHwwTBQd1Y3HWXyIRO1P9Lz
mrXjPwGBZvc6eX329TqS4JKZqc+DgmJ5l88vyp//zf14qYUPPo1Ch1+1u623wyGdscnXWCZBHFzc
mHe28bRk77/0uPBP8iamJD1GU5g8jucbqJxi2H8TwrHLj4RBI0NEk4uE9vGfVUF8PceSVNE1+u7V
/YIFuVSMecwtHMGIJ8KKKXCw3UQD2io+HGnpVRSJomOGIG8ZABf304ISNSIFX8LuCuXjGVIssU2b
+fZJHC7UK0itVHqm7OzNoSdNi+0P9lop23GJq3lR7JIIp+lLwISEYkIUK4vsnYnaPxxAQJDw03ld
eFfTRDJIltDozb0tHuVNfVipd4Af2g6u3ROtPAFkcYlUJYfw+LgVxgpcObSGCbdHVLldJ9xvJJzK
JrG1WigegSnTbR0aPyZGHqMz26PH1regOF0Sf3PvmMsoax7UlXtMzC99D+qtMJlXfmFvBjv2C6Lo
X/++QuBBfjeqWZafaqX7yxUGIsm5oaPrRiS0mTAjBWt9WTCqinlqu4DVjCkpKmMJY+QCjhf9ZIvT
fwExu6IbrxtHDgjHblHN0IMd6Gdh+SftYTFaMP/latCWsW6UHi+jgF9Sv7HX10MvncORgm0th99d
WzrYGJIQ7famCsQ9BOpliYmmIVTJp5okQtN8MfhXy+Ho01SKus+HYQKLrzZIJaoVHNViLOqqAlzY
Ry3SjXyQzJej6MY/V9Cr2hKu9rZZwq64jjh/Uqi5p1R7pAxIltilKOn8EPeQmwfzjMlKpo9WLZsN
QjnZFaM7wf/sLwuj1TWQGpuclcdrd0lAcgVY5x+ee/vFqLYkuzcj9UXPsSOGvR4rF+mE679kmKfn
6DX2jeLXxHLLTU8Jzp/GO0AQ5UBVr8dMcqDrhTQyJAbQ56FYbcdUYnUO0B8WGfSqqvVdFOKAwNcQ
dqLKJjLdkwKMdfarePqROlQnsUZKx5ixNs/U8dMDpISppWt3ZrXciCDl3KxQuGsQW7SgrCbeL576
fvjDaugHjH2J3R+OyJ4vZbb54fvdTr8agS7c6Yo0xB28SuzkKzpRt/9RCuLSOUBSaVOZV8dFW5tD
d/1Wa9iP8Pmk1yHySfJjjTz0X7bXi+sd4oZzRJooPFwAGucMOd9pySQ2mVoLzd0YO4bsx9S0HeNQ
bOESz4CNOrtMfsuLYpnl0sI6iKuFqc5+D4sALF/LDF8eto7Yi+6Fj5m17fgjlVAdX+rf2TqWDOX8
VEUPodAfRu/VRlTKrid3fYhiR9J7GN+OtdOtc2DpCWgPtHMRD3vyzQwsAEFERF6n2iM8Wxnu/U/5
mC5ckq3q8Ld4+qkVc3lEOGrvBio1DCRiG7r68SUt5WiaeMq6Tshxzb3P8pSESBi14SailTLOXnta
GEh3l3TAgJ3hbIAtriCp9AXIwDCukX2yNOcSTeljUi8RTJPYnVY38bp57Tv0ewzkliXM6xAnXa7s
Exd6czW+HRSo6i1KVPv/b6waeEFCibeLETW9OD4p7c1E1EuQgo/mfMS4llETi9nz8NyMTMDzm3o+
OqRupw434Epc4HHjkEQ0/JtsnkhXwIgFzxXjzss9Qu9xp8D3mO2dBazJPvuRW7TAcyJgEL/o4lnm
YUMrYtHGiulBSOo9xn4PaPffN/X+c4YUdOoZAXuLotXJBhCU0dWekKFVFB3di/O0bznJakt/Hcpt
yLdbq/vZrvtdP29TfcVjvSwTj+R+Q7t1bZQdb7dMsz/gb8dEt7lJJAI/PHFXhu90pCdCa+QOrl8u
9PBdBclt08zKE4E8QAxfHQTr/PE0hPkduS0Q0a5rXcucbLet3MzSbgEROuKjX0zy08V6n4LTn811
OIM8HveGJ76qCCDKbkrBx8yQ0i6uyZSArHSDNHHX3m8IduRpvy0QzDCgzeXf4AHCEQtvA5VeLau3
AExwJH6AvKMcLvBKyOX2L/qry+nvkfzI581ChAvmqYYgmsGooEc9fcUYHRi39JkP+RZVPF1mU4CO
sho1M5I5wwyszkmOyITdWYNj8RQS4c2gffRn0DfWSNCCbcR2Icsw6A0jcVihJiE/8QqOdPtpNTqM
za1q529bgzA8Oyp4EFqRsbbf33n/MBn9WEBcMaLWYM+L7Lntse62dokjKjzIocfRXUQrnek45UfW
qAOCtIoBbKC9h+q2vm+PPCrKO+03zaEK3t7Eq0JCdsrIAQ8CGPhTRk80rilPqPs4xlgPLbNuKwGb
Ken3ySiSu9VFNcaw+IsQRnN8vN/AN10R3KhOSe4I0PM2QloKrzqjp2F+QKEHwB74LFzo0AEJ2OV/
T5V7GCqi+O3ZPXuqSn3SBTyZqLrJ8Nzu+2AlgUSgCQ2zQ3C9W2zDBNIPz8vnzKJWQjsys0uN4K8E
Dj2WDGir7GF54FSHWq+Sio68NRyLwYfw18b38JhVufCf02ppa89ZtTUIUd3IAIMcp3+WHVWIDsBx
nVDtu9kcIdHY8ZLGXVjZIYnaW4hUdtXoyBtp6rOI5wvbNHseqefeYiCV7kBWr+1K+Um1OlARX4ov
NyEwBT3Y+DWbvNHgig0vyInzG4xEXCX0e1+56wdD5VFHEIlVzqPEK9UWukWCeVO7sY4jCY4OqIld
3J8jDWM/ShkH05Cbi/VV9PNovC3Z0qmdfXQz9QwofQI6nI9IcblbdeQlqH4naj6Is4763cnCYVAJ
n4zRlwqfOGTIp2HLn0oTMkhrakuQkWGhBs1+XqHpx1oxrsH4nYGGPKk0uBL9m2l8Q2g8QBTbKMI0
GidQskeKnRLZKSE1qfwjiBK8T70tLEi6X4c+nTVsCaKRRKgfoEEvPUY9qmpQ9Ov5+rbT1eDf09BN
miuiWkyLTM4WGtWkbezqCb1o7of3qBo3eoWImm5hVlHXvQstV1l43PhZNPolsXAu17OfWovnlsc9
4R1yfrwGIVLQo2U8P/msetscC41HlUx94QIDTyUSqnQuLFNyrozozWbMg6cinFV/6jbyeSNkJPzE
TySPotPWajWPNjoFJcKgcUt/aef821YjYC6rj9DDIaLFBD/WBkj63Uwr2fMg6+pV1xGyymPYKpH7
ReWJL+ykAY7Y45Yz1uL2d/w3TE2hdusKaeCPBMmxV6pqV87rNFt1q1XiaLxbV6CXreSosJy92eoi
hTRcCnsaT57RC/SQvyskLBP9Q6ZC4Yi2qHOTjWjkAS0F5RZff4bd4RlrZ+gzJ37S8Own0yt3yKHI
6ScpDkopgsIF4kL49sWLuesj/5lmfQmjBG1/PywpH17NX1OZAQ/2X7J3MetoNCY7AHrVTu6KqHzu
b8JVFIHKFL2xEoTUcKuaBeGI1jGorSiA3hyU+xSZmHYkc2EaTRygawIqYZlHFiW5q9Fa9TNykJO3
ie+Iz6t5TuxzVvDLNmsexR10jmgnI5PPqr/mKgxLE+m7ZRHLV+YXhG0BnfYITxzDDrmi3pyEe04q
3unouxKK2GOKg9LkLyEpgGbg4JSQCzH+tvwzvd6oagg83VBm/R8pCKN16eWCWWIn7FOgy4HCK7Ut
b3IwQWTc7TIgyuYBv8MkqA5N5y3dPf6qk/US3U/8JUoEpKZckgSulB3u3ZvVstRyR8q1JeKV7NyZ
101xw7ZmcPjX8SB8OHx7zWzWlPQF4pTOmsAKKlKaShfOl/sgo2znzKCCPUmEvEDVSqgT9W6PfBr5
RT4tQl85v18QE52j3g7PH1okdqmUrt+4gULjRWmRH73eLwBfbrdikcA1n+23mfjZTf6PTe61RSlu
7jxthR1tQ8Uozty1YElBVAtOvq6wCIJ2vNBcpnVJ46Ekr2yUT3v/tQsDDo5KcxXaDXsrvTa/YDGI
Ca1EDaluHz5eguoYGgu9bqxOJmBNf4vAJf8dmXJCInS3I4XI6HOTAuPmOZTv4OeKtdkiZ+XqiJGd
LENwPGGYGQpAXL4x1IEYQgKzkvsqCQW+1ynSVlPMvpfKFjK6uHUcU+YCms/3eCI7r5TRT9GWJ94J
WO0K08ZbrXObfP9f/5rd0VBVkkZsHkNMHSOUxbaOQmzdXajtIqGVjbLXX2okpe3u126V5lFYoa2Y
5n+kmMM1IZFEZCDN8YXUwVXk25c77ps762D4bAuB+JFHIVi/jDs1lF1tO0irJiNvkil9ZyW7RrZx
i68SXFLcTjomDk6G/OZifw2EvMuap1IzXBWjOWqizbDRPFDMqtlDBXnzIryfK9zYdI5CA57lb+lp
tXp4njGsqaZ5Rit9kCzZwNpn5jdG+ApOjFx2CSNwFtnYHd/SqnlqS9jaMly7WJuJo1mFG+Kc/Syf
xqeN+s6Wl7V3WWnWYXHsKdSTgLyQd+2jCfrp+Mf5c82tTpEFakOxRxscfc4lF3RqlgwVU/in9TTH
qs+WzDVRpRfQhrFmOjI5g2jUj7uJllZ6pdVg3MuUUOQ80h+5f9WEGydhLrVPW2GPiS3hoqjR/5vy
M1z7pftoYo21dU+M7L3h8XPFKnz2YnKrnBy5/EOQzzHyv33RbfeXGLk7i8dVvpxAZ+LgKgAtPzyX
5mr4zv4RCtRbGpKXMSAYJ+mRSOjm7VtXb5zPvLyCRIPfE1LsAvX+kvVSN1y0eWxHXHEwmhzB/mzu
Jr15Nw29fzew3XLLpHAV9+hwMcuatmVIheZZ+RNWPA8ZffYVvoIqsOvr1YcuDIzcic7iQ5W80ef2
2OZ7mi808aKT2dD1Gsern3GGkBUztF/ZVOlv7Aey08d9x9f/YFGenfeUCTjuFuxFhfFCFCHR/6zv
Qwi31uggCn02/Sb3gqVC/jOJEmxwnadxaPRMHrCIJv/MpkYK0palcczHzvSunF7bYxGAFMQHP053
Jiq0O1NfudYhCxXsO9TfXfmUtrbZdECWjp8hJoFsDv2Qxsqm8VTdzhzq1Ewb3gIqBxEUuaiyGIFa
8d36Jpxxtx43OpSjHNM6rkeiajce/iavOq76SgfyPWFD+peLHK2/f8j6Y5IrHJZIghEEfjwRs+oh
iuR2EKcOZcYBzxnlrbLn6T5NL2lgz3Cnw3+1Hhw5I1mSP170yEXhMzozeprITttL5Trti1x9bY/E
2YAgETEJR4o8D7Sdds1jtdcpMV4mb/wG+xX+QkZv0+8gmRYXcVrODn9BjXDEkSYIpk8SWoS8UPGX
FjTIlh1eSj+msnVtAy3Lc4BcQ6sjwHY7IaJ/uRoVB02Wuo4i/JzCzwN3bEVgkcV+YOlaYiVO9HyZ
OGBGbwNpqR2makoU3xNCg8nEwO57XSCrAin7XNRDg7ozfR+yiy5GBvfMLa6VmbXtCsFQTH33B/W5
OMj3jrKDOdxG61t4I+5MuzzoIaGca/WuCsPHsLiQ4U8Y77CiWJHWsRTMc/ng/pMvbDlxIFHXcYPd
8vzZ9vwAnX1fyZYEKm1A8doTBg2K5Gd+F0pBxAjAD2rHG+vkQHTSAXxEaFClD60uEGXlrKwEspgc
aG+VlRpSKxCdnxkg3KaIwqihhh8v2Cb+cdiQuvIcwGA+7Px81W3WxSwa0FngnT0KTlD9FjMhN9D6
YEogysz2m9MhKNH8TeJm4JxIwYxPgKOzZugaI53drhf4+E3b8UViLPW37wHlif1gujrR0mjZQH6G
Xp8xkMlMd6NGHLg0k5PcBuQPN5obI5xSV38wQXFqKzB0fvFjGY1qj4X5Qzef12SmASBQzcSIGetD
orxAZDkIeymISrnmACRkgincSrZC3iiCZhxUe+feyVbXRYB3hqaQz8Q4xQjDBAuT9x/GPnYQMzq5
toomzgLZs8JgKB6IIm+OmLePdfnfjCbEnsyS786+SZviJT2rx8w2Rx1Tw9lbCRfqIo4pNEvS5P1C
AHvxsW9iVx4fjUozuODoju37d8Pkyp16V8XlGx1A0Zmh8Ib+LyV+7smHJHRDId3sJI8IRDfxSonV
WPlT3lgyPg3srcXPZKG6tQwAjvOb6BFNxyxuD0al0mphZb90rfbZzUI5w4Jv3IRjgC4Ev8amoltC
jTxJRMkg2rx+ndDBASG35qnc0zhj34G7CudZV+sMnCer0TOmGC4cc/KVU5aNptVj0bxDqjBpCTrb
q0mH4B2X3hMnYrhlCOk3Nt8NawXG6+rBkLw0IdLrF4NVhXWE2ZQdcr7LJCfwx+J1CuYNW7tHZJFY
VkerlB1jVWeO9at6FyywnPKtVH5H3vmT6TyNnBnCiG4W90L0lTBImc0hSEYyiLxMXPfLLrOjKlnH
wScVpL/MyLF7wgjY25xAI8w5duIEl6WLCx1FRxglKiqfJo+vc4oD/eUE1wuegI0s72bzIiT5aJmh
/Kml+7a2m237Nxp20ZTqAT+GWaKB8P3CJztoEwrXbn1fslKjbrkE7VMcxgptZmrmgCCQYDYDzP5F
1hVjHm76wKUbCNFxy982Fv6Dl+7ieCHYCqBZWn2n2P/be8GeUu0kYQYTd1tg8hBT/HyhdTcyDumC
R56CsW/TvIqz+WNYq4L01YQrxH4VypOqgPYnG07mH5FR53Wy4Cx6t2uxY4YGdeNO8s0XT7UXEzpJ
OmpcIE9KNFpKsckQGJkgLqDpkxxV6Am2ZrF9JIKnqnmK2EPEjAnYvLMcSA0SU0oqUpRJgR6jS3SB
HDa+heBqquwmDD5Z+Jweq5QMdTqxeOSduVFaROWyr0VSrSfVgyU6uXpH4aeH6K3oKIBZJX961zhw
sNepxbDdVFpQRRoLf7P+hyveVl3tL0oSDtOcNXTpc1Ufzj0V0TSMiYKkEhKfFmq+r0fnPrSVSzEK
4qc1TAkisVz8UdZk36t+2AXjg4uEMtKdmh7FPqeo8leDZjVNHX4GevDkIUI6F7VoH6HtMz+v4GUi
ad/MA3zwijCeVe2KXpMbBS2gC6odqPHTbrDe/TAIxRyd+AIwSSWYcNsLtYSq+OJptlcdGj77pkdm
S1B2M6uYh5FxlyxP8TPNb2jMXCKBRDE7HkAslhboRGTLgoNmQMTIK6Hi4Qff+pqPQEgj3JdaXShN
bCe2+/NsxatlVrlZUUybuxwZo/lZPXiMcQi/7s5xf2PdRdR6OgsvJK6XkiUJSWpWtamGE6HfTSe9
zksEoI2udO24vI3fqOzlpYjUZnCDoLzkW32g3AoLK4CqEOJPrmF8rH2WOoWdrFoTiKn90tnk13sA
NIrT0riyXLQ9piw+jOrLBQiLqzjQ2eJll86ENLMpUxmap6zyLsRF0AeJe2dExdb5eIC5Ts1mMxXe
U0p98oflYVR6g+qkdfAmz886INAW4zO4dsCehqSt4PuQD3s8qzzmg59cNWLraC6QiTgZzQKqddCd
6YutqUgSwGnlFrBHRGjzxjOc2fgej/iR11LHOAE0Jq8D7E/mtpyAlLD/LUUjoGr1/G0GKS0q27ME
sAAZOmF/QXIN0YNOuk1xg4h8736b1b7SG6vYTcHUKsAHmDxZpDtjO61vOZ4FtyLXdkDBQ1hXN7Ox
vaTAxY4Kr7XcQKw05RsHteYaTG7HSuaAuomeo7EEVzVqNuO1Ee9IhM2Bhx5ViPshewCZ8bVAVrYA
Afk9ZQxcV3ygDvBuTFE1JCGQDMdrlFnn5YsbO2jIJLdFhzU9kfvIL9DWA0o3/CrfgiZc2kRchZOh
KaIFC3Aa3elHtKGIkpbdNigfrjX467q/goQbnEt2/txixxO/oECUgzMLqS61BB2NPVfIFR6RrNx9
OdiuBKlt1dA5qPJ1iuNMechy7IHZuaqGBWYpttYo7sFQUkVrrDQBB4GcdI3O2nBLE0cVVPvmEVSX
o2oi/E9rM/VVl3YzZYe1D/yrJ1p31xaXh8oTeU9xoUXY5XpjZPPB/dx1HPJuqsSJARDSsZy+2po4
PCZCq0NC7dLfLbTltDtH/9DmxitaywdL1TUdGTxgZSj4XjpMqCBjjGM/kdnuf71MTFpbqmkNfOwX
kCYmIzfVbiMr2Z/Dq6FQw/5udJc4n5BGp24uEEao4Eav2VAgkYB4B+Q14HpOsm2veQRDbvph1Buk
4GT9HeTKQkL+zyfFyXlBk2obAMMvkSBG3Rw6qjhMMZMkAgMmIoKoLgsyeewS+jbXfl6zy5c3WfvN
GQEVhhx9SiroLyrTDwNtzXjgk9KKEnWitmcdIGa814jO4GtcqdulNf25Guu9sEao1Fa0JPyBHHd+
OQ3nw87JkKszPyOoTd5omOpdx4iqP6rVLnEQx+sMFD8gLgG7E5TH/9lSXHt3pMecsKCplWSvE+wc
GuNyb+T1LTOFsp7Li3ALei5BCOGFsFG03e2HhyHXh9AAAu7zjgCZQ4Ze30yeiBFUrmOBiMs/eQ2d
2Rk+4oudAmzsh61AGvWZVH5dP6PPEAY1t8FKQhihitdPPNZghq6KSICEb0QEj/u4g2CJVUaaDZnB
U/3+lt9fBnlADacsp5QQlZu4Y25kcXL4rF21mSChn03QL078wS3xG5R5m1hp6XDYO+Ne8cH6zsQv
5QwfM5IdNZ9p6nI9OsXJYkTHEPhLIK/4YfT93mHLT5Xd6ZNOnGpWrz+DTw2elt8fW0i9yhMQn5ac
QAAwBxvEtQBhO9IuVIPdBfyoO1LSTf8ppZYM6flLECwxjE+tQDmrhduiXLxY7b9D4/ehuVnMw4II
AvMNXLDd4C3odJMvHZugkt1vOvJYlCV1qq00ByBLcknNk7rkS9tH0PeR5e8MH2msMO2scGbYOXMb
j7Fe3Fb5ocABl/B7DuyIzIOUq38afvjjKkq44uJ4MWubkNCC5uiiDfuoC5Kv3lWBEe8+yM4raP5b
OgJMCM1U/W8VxTdq7KWQU9qMev+AF0lm8mtWSxhll7dk/+nOQijgVoC31vk5ix9yEd6w7yaLAEOS
K7vasWexz1lAf6DUOIXWpU5gy0R1tyErobnahSIlWXt3ya9za5LFJ/obNru7kbym6Vo57Dsm4jrd
4zMKNZYbKfkQJHKv2g/6TrAiJddPV0V6QuadtOeZaMoQZJC4D+1R/SnV1AEfqV5p0IJMKBU5vzBv
suHITHomMtMWXuF+TdLfHU1t5bpXTNZJ8PPWSBFr6SibQI7RVPg/w0/E9WM60+/1ECdpZ8QdthW6
0kAndGnZGamLYY9gLPiOhwly8dWac7/8+8CzCYEukF5vmaclxrMeOXd0xJ+qCSE5/v19E+8L1jBB
GtdqrjtiyUoCaDai5Mj7mdMnS4xef52CuxzMA0dpL5+sC7NbvC2/b5d1NYe4cKeERWLSBSwcOIuq
OygOBQEKOLslPO+kklZSOCnDnw9zdeWgi89fHvuiSpeI2IelhHnvjpdjApKLX7Ip6d9rocKMkywq
9pDs/HBOrn8B++7zZ5X57xwc2ONeDDjv4JcrvSTFd/SkygtrowLM9Hjcyqxg8IfnDoIf+r9HDBgY
KadUFhsoV859VjMnUccJWvoKP83psVGkHc5fpvCu6ABfu5iNasgUw+cdXQjOaajObHKWzcKutHKO
UnyAtG9n5fYwKD/zeSAAf1tjs5xIKGyjHsfk8xU3mzryO2LJRdTftlw1E4UFY70Kem111cHcXD97
Ri7+LNgvMTUtuBr59GIH6WhxSC4AFH9csx+uLw+abeq83Jfyz9h0tWs1W55lgtaXepFoNRtxViqv
eHPROnE330yFXbpnpgudGFPF92i6b0WNyn26hCcyWevcV8Ke/udV6JP7b/qUoTMwFlFLYXL1pvSX
m3QFUGEGHWsZk8Pb9L25lk7lmPSxWLd5mgO5JP6A3QVHvD9SJYhuseMLR34quC2DCoinXvIZrNc4
2QTWpfhFmvFzY0Aus/37fSi+hC7IxkKEGxv7eISaJRMr/8ZtiIqaHws4yEgxV13ngiza6Ywa/aqp
VxliVaUVMCQI6uor5fUYqHcdHKIM5M4UzIkdS0gWG8yglZEQlYzo2A3X9HR+TpZ0XdPPXlypo3jh
LwgdFv9G+cYnpcnZ8ggAig3wTy59jd70K82OS2q40j6J99SPMd37sT5RqaSSnf8p7T6luh+dw9Ko
ivBtPtEEWcb22Q+33CgXnXXltgbYzIRfQPQ65K0fD30qWbRmHQe4CPPqAFyE0EtcCdrO3v0ak6kI
dvImvn9UBGkh/UTBuTailvtpVFvr58Whm/aJ2QNaZ2CFhW9JHXDxNTPXUqU/hFk+uhiZ4RUdb8el
OoVVHQHy0dB7ij2YPgmQPVsXf6jwcgQChEQRtrx82+ANPP/6DO7EXjtqioDGCMPfWTi0QGRPe4aQ
RchUvpW+dr04ZUTo1UDlnxpxNahPN4i0pdQVXpJPa6U07spasCljj+0VTlV47w4b8RNT6WCMg1DE
15hPU53nioZANhELl/IzJweJnElpK/ArIFRTqpG+MzTNOX4zp8XGT3Om7BwCq5k0yZ+cWI5dLWBF
1rb5Q0aXS1vY3fOnvlOYR8ruhCTIPHFbBnzSeJYoiQ4vZ7RvyRMrxXz+U/Hk+UnZp/WcK/SMLM9Y
dbBwuouS32Zor8tVDXWOgHZof2AGMavsfJdt3D68G8l3zZJn34roOy+tapWoJfBuWnpubaxbumk3
MWHqDmFGEY7SgQi0+xWxgcPnVgnsA0YDnjSX7E6iM5b327P6YKKYOKEQMwl/DW5GaMGrkPS1Ee9m
PqgvCFSJoDh04tAOKiunaakT1KgjhWcNEKIfreSuXZFMZT1vBFW80xFA8hI3CZsyZl45tIeKl2ip
4xtCVHi5PZmHEQmhST6O/pzu68fn6P0SYmO0Sys2o2gTgf7NeGFF5vTr7knOI/jrh+m/Muytwe/R
mncdSlQ2zZb6Sz6DgVUZcfkPzvpyEO4CpwsKnjYDFf+bhxEpjuF2DQJv/s5fnF03AY/H3zdfnIt5
axxXzvzSC4I9jr7hSK4w3zRaEhy15OufOe8lzK5jx0eSd+j6+go9Pvc9WMcZk6flNPR676phpPxJ
SpK1wYU9hgk8pYUaccWQxge198oUIJ1hQ6pr0PtUoBWONtbNFZUqDDnPmAJW9pCXrlbSQZtaQRmf
ZJM8kHW3lrGt21ED41ktVgfdMjzPSp6ews1uMwZSElbcKGNFWKdooZQ7zqA3sCNsyj+cVhxiu2rT
wfCBC+BOqPLg2vGDw1Mtb2o0MweuUGw0v61cOsp9EQ1UrEHpm6noGTO9WLm6vje2xD0LLqOBwQCi
X+d7HV+anBUhk0WRCj7jWMQW97j3X6Ix87NfpjnmnochVrAvAhHwi+0XXI4Vsn8+qZRCh7K664f7
+oGQQ3HUG79OE9bSYtec0DM/xaZ7fcuAcLl3PqduuRZ/6vrtFDKD4Vi+blX4mBb6oZtwBlpRUCra
UedCPIe8do1sDjaTY8QPcXFM9Pqp/N3OLM+v01VfzY48GEysFKBGHMZpaGlhR2NBS1Jqf36TW2qT
lHTa0LoZgZdvUg5knaLulQ0MuhpL9ZYH7EdxbaX0Qy0fbidMHk5YfsePem3FKvoku7tTp3ilynEY
a4JcklvSPHgIelFwGVgse4pH1/VaxBaFlU849EMwdKqfc7N+pnmOSzb1NzFpNXg8cJQNyp12mDgL
YfUyX5tnGCPwgSLWzQCtvOVMXbzR4ttXkNco3dFcszZ7/j+7Q03YI5dylv/iebjiioRRKd/PMpH3
cS99zIe8otr+ui9zRVfZuQSioG6MCtHblv1gpeXWNMwfv2OqMIv6aLj05GxG/KErnzIlNwlta25s
YKO1gtxsYM38jjY2n4kjtXONUXmlNMrn5bDFx1BVhX9eYXzWwz+tMXIc2i+FzSv6IUJtqlGrdPiv
cb9qzT9JDNXH2yiF7o7Jg3Uhouu/RD2Hrkm7kWceDGYxRnsL9eL5mnAE5JcneLHI4+rM+CmXjPoD
Bxh4KjUAFUgonN69Tq80hdfwQhlPVcGTWr/LPL4UkPS1l7+ln6OOANGlt7721zMEkIQv1YcbyIlT
DTz0BpNzbRCVSjePZWoVE6HwQf9gtUYU2UQY2mpF1gz0us5uc/wnr9Iu+QvMqnV29faoXN0q5M7g
puaB8n/RWOlDrR2GFSl/QBIUw8tPlSCc/yrSY8KPx1GGKt+gYZi52KdeUK4IUE+pL/ExBODcgMSx
/fjA7pO6eHU2cmxA3z8DVaD+mwZ7ffIdEF0sYqst/FfSu/GIcpZZokAmk48S9bP/at/awQ51orFk
pWDxyWcalP2OEiKbWzeIFIPiM2BnHnCXsgCNYoBiD9g5JW7noznq6rF+iXsktdtoH4oIAtBb3QCH
KhGlrOapflILUG6APYUx/MjOvVFBsC8iMEHYO17hpLKMs678rIV1N62Rzjrc3VluJlpx62HsxpOT
MK4WLejdj6djfw0usSrXXZ3B8pDFkSrgU3/Z1EscqKBAK8wPueTUid+zOu54mL1v0JXu4SSvYqlP
hAlHFGXNHfUoWIFJQIIbjZPyZXJFyksZy5wUe3S5azgP8M6c2zKDXf/1YzF720/iLeO8dfw2tkSu
Ta2G+eR5tkygkcDx1nRJYP3/rmqC9OXNIGJTQjyHAlakBeoHpeE3aDsNNs2D4UGaBQccDKurd1eb
kOQTZomlQGKRL5Dp+WWxBiQf7A7aJM5nSV/nJgUtPV6T2H2BatDTYdRf/vY3XObFJu1R/wqJKEKJ
5E9BqwwmnI5QJYTd6rPKuYoXuy9Xg5I7CtcTI+V87GKxwjqnsTzPLtjCfZN5VBqrpPz+LxAfHl0R
klZIZSBn0OzIUdMby9qxypYbY276NDzLwbbQgcte6mpbzds7iBoC1bnKcfwP8Ib87ye1YntjLWth
wy74eSaYevDBSGXhlv59h2oJP3VrnRaUA9j1xiQOfG1ytcsNpeao1XJ6w3JTGl8RllXRAVbSAfOG
5B5QnZmhE4CWVT2ekCHRomfc1Vop14pjU0loDw91SC7E3pwP35QQek8/jo3xqfLWcMACyleG0RD2
ix/6ObN+9ZGOweJM2TZGL+cSxDx1AwwTHf2Q7oT1GdHtuiBo73BnrjW89dKSmzmmWyuHmEmLmIVz
ud2jeORPHMxhtdp8Xesm+5g28v5889RkaOkvQK3E7aom+zpCOo2ZfRLt0437TJksBJ6hSK3qCrZH
2wF6aWxyPTrEejKsd7j+qjWwqK9xOvZYS0Q4jjWTJmVS2TIsT3oIQm+cL+eSAGYnAC6ZLhvjR9HD
OXjVMnoibGvNCdhqndfbIIdLwQPU4c4gijxH8DlNk7sXVjKmiHhLpAmBwMknohYR+7DMykuSHH4u
xOxOcDkna+YRGTOho3m+gB+D99f1s7isJD1eyIqQS47KqSq2gqDfjIrxzcu1nKAF/2dPMhYubUU1
Xvm0NrWmlGDLGnLxBVe22ULJ7nVPKOFUDnxIs0RdevlmDl8jk6aGGlcYcMXirGp9pLcIuoegrReK
Eq5xBnRTvUY65E4vnysE7N38lois7aTgwzPT9dVNgiYO/JKv//mLSf8PL0IWt4pOJiIV1NkEbKt8
kyvCaCp+purMT7b6h0HXYFWwvH4ZKJ5eIT2DFOVrpCUPxS9VwxmAUu2Y3c0RVRtgIDozeXOpQTq4
/iaKXejyTq+kNph/6ocKbdzjsKljWxMTEmPj4vO1xL6qf1gl52m+lwuLFLlQA548hpjc3kkTaoLR
TLPkHlgJoP5SC/o0K0gnsm+/nKs6b83WrEVI3UpP6+5ORZ4OVGew5bWsRGd7LCFtY9lg8Dn8zL0K
1lQgjWeDEEHQsNQq2DdliAnmNYKU69N+ykfEsGdBvmRvrWXTPtaxo+3dY42QWUjydHymeihk8nwY
O4pQmmelm5rsI7qph5vz7LVpsDhkLpJm0KxomWDOf1Wh3woHLz8tarKv57asIfPo3pfFmH6m1xej
hIwCc6bmUq3GoIGYE0q1M5rPYy0GAmuwO3JY5n/WvedLAECuf5aD+eGZFGtEu3lzteIXdq9fv+gt
9yflE9xxhvARNmGIVGN42uYvLuy5e2eMIpFuReRDw/oLOwfKhwRqk/8S5RLqr6fea68Fn6uYhNg4
v8RUEt7fxQFFxNpRU60ilb8CYvRShPoglc4DzoF88BhgPbzZMuOc+mt77Subyr92Sm0u5Ix3H5SK
KHbe1yRaary407xCW+uXseC6E4tHSAfZahWqBGRn9k/KwCMvbWDqNbSX2RwgOzGkdAuogRjG30rv
ofg8HZeS/2uBjZnUmnoWxvyDzWJya1SSgHg+YimOT1olPi9A/UU5jplTbQYI8r5mPWXpmSyI/gNz
LYpiSLOHQ0/a1AempJiaLVT9ZboYluCOZ/jdJQs1M7r/kazqQ0Rp5vF/zTvxnnk6kJWfBxlnil5I
gLZVelZinwMeBZosILs1uhzyQZr8jDeH7z8ccyfwDLHb5L1ClxruWkblx849hx7ceUMG8AODBaBx
cpaayP7URZxY/i13bR2jGSNEw7Vfl5i8ag2ZYZ64rH8gz7peGX6Ldg/QeA1zjgtqv8LAdtl9xggH
LM/VGEkr9qs0sRmdwmvLwdsGZlG24WS7gAANBOJh6fO7jLPKTwD9VRbnuE5sGmCgnIMmAv1FqgQt
kZaezkIsiJK9XQy5ZSF5XaR/VwB55tIhe4VdrfIULhOFbZSB2TbbaPta0KM3vAQz/RpQVJoUa2k4
wyutkfKHy8CcNiCNAdVECY4GtDoIvQniYnD0NqnOvONxVFrpi6b3qsirUhaqDF5YvQqoU++ZDP59
bsOu0gwEdRvz3VSvHOvn0w6zc+H0vPCvbZ4oOrFD0ti4p33hbgvjkzEe2htm6oopQws7Psl4v6Ra
XXdmuFURazI0OgMoyuT/4aNzQgXDxFctzxa3fV7iCIZJevgY/Rh94i8a88WnPkPZQyo38KpAhySt
6FUcuj7X7ARJaqjiOlWhFvhSO2BpB9IoEoIgr5FdapfV/qGbaKuMlV4PWIAAtXATboLB4G4uPdzG
V345oTuXhi3h+8soMbnngvl8n9QG1cNV4sacHqWHlFPVDAtiQ2T+Vcr6jbtIRIzCzIEsXFX8tThx
W2DwCro+Yzi147c9S3zOoWoQaU6tqxDPMYqHDMj/7Tx+fYS33QYns3i06T9B2zMXjp674FoSaHxO
cJiDeCwukhlLJ5xS2mzfOthJi/qk9yNPRP+tKCEB2/OksWWRqLWwtPt/QxidVq0qLtuxA2Hsxo4V
GVugSEhbFrN2QTwe+UdrlyD2Wk8QO0mfkvyry6L3ypXdlrGZvbtUmu3S7huoGT0HPqTtm67udxsU
qL2N5QgzInBntBXVrA2ri2OaINsY06Om+/0/GX19fNeBoBfMcCWKg/uvGuJH+tIyPN0aZOibKQal
Xr2Doe/FYpvtSD8JvaTxcP1/GbxkkwSDbneqdrwIXTEr5Evr8dJE1He3QeRcJj/JxXFKOB4Wjcau
ranmwQm2fb6vewwtn1w0VVZpOgSQIixMIdhJyqa6hXZsVFKuxXrySreDfPFaYbPy81BraMcOEtf2
vjVO6FD5zGI1cJY9nhA7vYKm1ZNGZ/W8MLf7lTiu/3cDKd4q4yKTM/tMdn00pvfP5FTEW6exG5yG
x8Y6fLbVrqNE8gRUM8ZLi8D8FCVFezwSql1X8Cs5feF9Fdb8jzCmVC8S7pMq5MMx4+Z+PNBwrFus
34gLU3ndonmZLl2WsMioqQ0THhmkf2Qma9Pv2WNUSBSfQ9v1AamITqxCJI/6+LufH6OurapZSqn9
7cAV5FT5yMKeJQiPzjahBUuq8JZL+8d3r9eftCMmVODV/9MPoQAUA8UNkUncl53c4XKaLBy6kLcm
CkHPkX0Gzerd1BqXphAflRlZ7H7R29VysNj+sjGfNQEwCWhkb+BMjjfpwcIsaWd5SV5pLjU1mJZj
6Kihm9HUfYctSiI19hEkpDqlPhFnE1KCVC5ko6ag4GUqJXmj4KWSrYlgudB2U2AaEGrHnZot1cdm
OrPBUM0T6ZJsizE41r+w/w63lcnIABbHtThuvYge3sCZUWg8IZcvbCs6G9qKuB0/WTqN6bdgIuhe
7y55cVwTja0YW1nnHC0ggS+P12wTCJxKAK6Fo8zAYCPO0pWIPcvHWdZgKzp3K/wQ8l/OUuiFaLWW
UBhnda4RWu8LrkCTOJKmQw3P9UzsOg8hfjdLK7rP569RhduRjxDP+GoDygOLysKc/YzwnOJc+FE4
1hOWcEA3aAZt/4mt6KJs/8IO55NyWUZI4vFjwY2nftc3m6NQl8W35osb3gqP74D7A2NhsFOACs89
HACRS0+FdsLBfyhDZqeAUJcINZ/+2RB1MKSktISWS7+V594PmVe49Ch+xg6dkuAxGSCfVv3tT2W7
2eLAKuWRjPA8FyIUlM5ugbdmcF5vd9qMManuwkrjQo2d9A/FZD/KlpIeLIP/fPwXiIXfXW/Lyw88
xcdBgYGXuhjPB1FrJWNaczZ5f/ULoiGmnZ7hspfmy0Z8HZ38kam13sOJ3bXuAUB6VFwnNcQDFGE/
T/hmAwddpusky8HSy/6qWbIQt1obWTER3QTnfw5QX6kZRaXbQJl/9DFxl82Na+YiLQ5cnMeWLuQ1
rMBSkqaYYYCiHOUtTBQTqoONPvXIoga9Et9qkXKMnatNjH02nxCmmrFKHdcF1yhuPXXVa2ua+V6H
HRCqFfQKINetovPkeklOpnsfVMSxOo3a6+mCoxiOzQYhCp7CjkVpHWYLlcE7sXbQCaVSBFjsnomd
3faQGTtR0+MepHuG8FT3tS8SYu1CVU12BXjon4E8SPqmAjr1PUz6rEfC+WGawoMVFPgGCI2EUA6B
PbQK3QQtKLDaVKr8x2jeId8lF4lTV3nkpzxnr3M5nRoF118qw8wmbGvi258MdjT3Trtvf/7bqHUO
qcMvDo9Hc2w3OCnG1iBQdtgEVI3rq3ZjmNYhtEDL977ElifxG57ePauDgeD9PTZXi57KUlKMuLh7
/8obYo3AreYLLy5vx/Izx8eyOITaI8qoA+pANqBXy4hfFkeUwdIi33IjkhgT2UX6TB+x7qJduL4m
pqmUx0ammHjOr1fBKvFFWaNhrtHpamjHUYVSYnJXJfCOjZW0jNbMjD2U6o49la3Gtkavm5wEAC/A
h7gT0h1nNc35iOahDgrD105vQ+T+6JWAR0Zwc1sXABm8aKo9jzymPlbltTNNog28jd5QjJGEQ3LQ
lNHX1CShHkxFr1KYub0L3n7JXBwJqibeWly/wPZIAloGDkhYA3/8RsU3QIG6ji3hAPKPrloLtcn4
m1dNkpv8RTtkgIzjB/Dx+iRCS6t0eHwT2DHE9vdWwCJ14d28wkDh8DjR4BCzyfdW2ba9mpGb/USm
JfM3ubwGDi7F/CH3haEgGRutKSurvdfQeDBstZTBIBRKjG7QI7Yy0g7s4uumXeVNt4Sxsd8JOO3s
38bLPY9yWs+O2nctQ6Z5RmiDKnZPkdj5kMLZg5WEkPLy3eguYK5aK3LtpvtmlkJZeUQynhao37Lj
2t4C2HN4hK2UVy5VcA0CuK1sgHzwhjQq18qoPFPIyMNKbJueTDzhyCHmEU8jTEcn09gLFUPQ3etd
3Y54MA3dG6UfLpDi4idflWdhMPEGKAr+9AS9LVtITnSqsviaHfQHAdCD9TsT3CO708F8ptZoAny5
V/JbeeBQIY0qC2HMUHmcSY8B4FNMqwaEFx6C3W85vj6qzMR8b0MUT8GVYr6PV6SrxqUZkVpFQiT9
cIlWyReQfzAgDWb8YUxBAKOCF/csLks3Cc7DoxtuwPT16Bl/7Oxr+3Hus/WM7kAFN+ur2MIbpmkL
iE38M8/psmjGX5KmZu7hv8cFPpAa86uddz7Lu3luksbBxc3WlXTuNAWoEgiJhg5c5FIuJ+/sfnZ7
D6OoysMo5NT4FJyG8UWmXBr5xqhT+X+VchbDWfWGs4NCZh95SV+Pm6yJwCzzupVnt4G1SMySf69Z
dRwx4EL+f2mfkLlT+DAqJY2i2BqZAynG3NTeJ/M0loDWl7FGCcJ3pHkGbKPOU8SNl9Zn9Ter5y5q
rP8YzLQWf49iZy8qljnX3LJbkQxylphlh31cvGLUIDvIhoG1llywdQdv4rSS1JYRPuYpmKUbwD10
/nrfj5ZgquF3NITC2JlgbankehMXKTglqqIP+Zft7ccnG3JWNroYNZsYSKLw+D/h9cgS0Atr6jCO
Z3rO0zXKYSKXnhRZGI5bAn+A8x0Al9EPk9NfwuNIDdswsPVBeT26oOm1wLr5BIjqJDpaAUv8p+ws
Zzf6bjdpuSqH2ADaKeOhNR1xkD2v3ekA5CZwC8GMVl6CZVedR2L4M+6W8Nrdcv2AFpe/5Mcxt9kp
xGj5KgWMAJGw57ZfMehhR3e1QKM4PYmZneh2D84NYaVcKBufRgbAkn7FXck8vhgyhTTEmAvnXk1Q
SIYhpA1Ucg+p1nPAR+K35/JE+i2e0a8mYs67uyvG0NDlpS5pcgCsFsGpVk3iCtQ5v5tIts2B6724
eqDwDyTsqTNZ2YPPogIvUJAYBOxKP+Q2HwKmWGc8gL2oOlmwTvi9E5Yj+zf8VX3N7kUl+TJJfqsh
VkHTnYplkPT7oB7fYFEIQY5yD2az8OpS6jKY6MTdKjQrGY6y0P56Zkg8z7Zd7OMCjbKUhmlBYd/t
98z9ytbyvf5I31eP7crdBtqi2gcqQzfzB4EL36cvOZ8Z8AsBwcRg2Pt28BfC8hNiBofxMN3gzGZr
GFjdfo0nbfO04bCaXTPrzBuKh4JFpFZDf4vQNuqdOgCtUCbOBj5QwRq3pEo3qI6BIGIa05StJR+a
VsaUIF32TtDIozsUTEhwAXbhPXTXkYCwJxWS50kVdHK2rDA8Nx0ROjGlgQ6tiVUx5urCLGQD66xz
m87QvIYLiIul1rSCaiANICVqkJ2jHcn9u+T5nLNddI3ARqRnzxUmagupOsu51SN/ZSpFQDnMxG77
oC7ia/S1QPbvjv1egEORMMp05+daZxTKKGK3BuV0OXNSA3mZo4LzdGflx/9L7t9G750VOuyATcg5
bu7nfZ4hnb02Wz0fWNKybfFDHYYQlIKdvZ8UC86+asiCOZQcQHOXzLZGwtgnqd1i8XjIfYRZMwBV
rIt3f3ifdgsXGxjbHPYv1PqMaO9O72+WQEuKX7e6z5fF8FjJSZwxb15j6RftXYcadokRij/lL5dr
1lWc8Jo8TSLvH6rdO7XT6YSJlZtRXSO5d31t2H9pDCHHiQ08F/YzITqWDMym53DGUdf5eCCRGFQR
EKhoxJixImcEbZH+b1tHlD0F6ySR/M5HvXfsaZtw8SDHW+2lFuh/WzzAkzSq6Eqzv8dGFT4IlfqA
VyPYOdfNXhTBvHvF23/pooqfXdLt8QJtFicQHScR4MPjsJToco8BeAni3hVFhVKF3PNmiMLc+7dy
COzyXm0t8ZXKEoB9EOQQ5mn7dKyR4mqNutJlWftRkhNATzFAskpUS7gERcPPFiW6mno6/z4qx0pM
3c/0DUVwv2CEW78BBguwP4XIWa5O1ZhZBkrbccU2IW+Uemhze+H1pA/+yPZHjRskckqKJqZoIugf
F5NldxtRLD9G4qOjZGDuDNjufS/R0f+0sEbgrR0bLIuVqMFVW5zvBvve3dpVIBwJWODjaHTd6caP
oDb2CKRlFHW8UYNzlCNjmVCFhElT+LUa2KBjIEynk+DYHxVSiWuAKRcpx2/3LktqOBWwjVVECQHm
2Yi+EREX5gP9WS3txkVs/6q08mUTsmIjpYp0SyUmy4k8eEN1+n35Ol3LZbnMFHaH0JB/3U6tjzC+
OnohGv2IkvDZbdzRSSi1J8lWhBBszJW/cPd9kSs34vn4lm3jHs5zTXioPD2b5LpzpaVVCJr7qd4t
0FzMXVxSrBH+Jvoo+uJBOjQX0axvpHijzEHAYXVlkA8SK6+P8LEOWvWwLj/iDJFciS5OhFNd9jeM
75DIwDXSp98PhswMe+JWX/e8AlUD6WlK5DQGKzyPfVWskacK00iwjSdl4iLVrKIu1a5YXVw5Sx5d
rpanT384qGxiFMoxmmoY0mqpIVJrFxzoLo+INmkRW+M9xBBHb/OTLvJHK1nTD1WzS9lXISoNEY3i
2eqkSVcEAtgi8MfsbAsKJM8XIk2bFGouDxA6OqFYnXV8K0N+ePyDEDxEnMtHmUlu5q7H7jl+p/Ip
vuduuhFCGVjyFo8jaM7zJ9PfZdvztta28ndzhlvYWDcgan4fqFqOo0K9ANnkqP6OlWX3V+bIBHxC
v1iO9bRYePaFbP4KsNDsO/d8H2a2QXKSlLJvqZS5NaJfmAV293EsDAmTAPW4Kr4WK/e0CTSBmZcL
zdSD8PIgaVHd6XBOJRJ4Z+otLCjjIxCeFIhrLJK7z8hmG7k6+HQoG4ls/LoAca3fI/j89sczjx6u
FRbcaAZRsb+c8KGPdmRNtOvq/p1RAxZkwKOIKCALWDHdUepkjTPktPeqoQBjTIqj/CMw+JBteYrl
UhAECyDketAPPlPp5JP9UJJEJT182gf0z/D717sH/r5i6uXMksQEPx/q5N3S6QFQplcW5kbQjw1V
zlPlSuO7GqCSCv/Xo3acyBKR8NLX2QcqmpWYenEzC0vC8BJvtElp3gOcQHegUipv1aBdAnhfsvVs
a4UqlGguVePDlQDd58gf2AD2SRnUKS6H69tRpFGvHlnevtM9d7eyIefP57xrYjBInyHxBtVESPAn
pY9mdfDO1bGsYWHS3sU7QxffTQXTHnw6iS+QUrVNG2mmu8qGxXJtHgrDeRuRD8t2zaGR01pW5d4Q
hoiUKd3Yh9M95g5GOXgNECAmg6+E5y3NWswh+GjWFnCiDlhS1fSFZwBIkD0R3vy48axWzM6ZJeZQ
BqyAUCaEuXW8q77TkQYfMl/ith5xS5tqy0cTcSj/sePbefOZ9ZKb+/eA04TsqqFO/M6BmEXbDrWP
z4lyj22aDZbamU9L5bxrFKut1D/7Y/ahppqr1AiSF/9K9+g6NzNQAHmulJNTfsmOm0XcCtyPjbsO
7QQVtgCbNkl3JSnqEshf0Bt30vVgUsm4ybBeMm0st9Y4fWvXQCh8i+KXVLRg8ANlqBswyqL1QRI9
nNsWaZaozcJ2HXB8aZveE++E1iOThOlpKOr965UE3MPeneuBWy+4YlHAMumkU44oFXi4beO5rUJC
BwqkvdMTO/iYYlI3zxwnT4iPE6NaM59L+6i5Md12qyiSwEIK3492CqMPXuEkHgnTLHdYiqfzmYIl
ZIFxK2tMeub0P66XCH6cmfpSXV2qRf0DypFUtGPWB9q/yotPcy8vaXnetU1K3494Ef2WLTq071Aj
I8WdNid1GqWnUAXuq4noGGu/u/UxL3gYHggBil2cIxipyTiFr0J+6pegq8vBMWuRx6nmZqlttaws
L3pv9nJes2MtJMVvMt+Wz3QckVsbPts3ENI5FywIdKpjcBnTfaZsm5WsMtWssyY6L1fd5MbFys/G
9HUezIDSo8lQKZ0F/1W+ZLdSQZQjx/kHcu6zikbW1IZz0Jo2VZb4r+7/djaeDZbGv8MLf5APVHQV
ZistJaxZO6AYuq+D7IU/skqqrT5rDIyjZPBYRckWZhjaQ2tAGg8cSncIonIKMZtO1ysPNu+ddofZ
6EZIVvGkdd/dElp9F5E98not+AoM0NG1w4hM4iukjn2Dr5DX+O6Z8Qs0HcV/altd4ysKH+/d3+RZ
I4rC4LywyPsLDeRdMLa64r8xi9smnVP6SgZRjksALf4Fds8HhgI3q3UFP++l9rJpB88wq1RJ5f90
xYXOauytalbuQfy2b2+HHQNFcm+wx6y7ADaQ53Cc1XwfthK2+9ELFkd1jCHU6y6PjPOgGqKlossG
RdtKGRQuJoYPD29rhHQblqP5gXFMhjVIr3UHGIsoyDxijucz4NDKY2xc5GY7gvIsTH7FcFF/qMMt
atfr3rFzu6Lw6VrIaNSU+SH3DtlLz33vTOaCwLqzAHBAvap1ZMwOaRMu+KTxTo1L3XuTu32EdYKq
13NHpSzWVxCBzWsaXOjv18sDyNXgTqo0Zj7WO3rl1QqJqfWhmmmFAsp/GZD7WYNnIFRkg2zJItAJ
p1y10WoIQmpKydR+1IUmFl5PetSKz6Q8Ejpq7CPkqfd9GmC1pVKR/yxJiKPG0KNPEX+rwP91SWHf
8+qHYu+Mh+6Xi2L2hnJWgnYgQRPEYNKu1c7lGtVeGhvQ5sJ2le38BLt5ukrRsimEmeUQEyWg2gH2
aQsM9S1Fvb65By9n2LQIuo7K61W+R/VDGy/nK67tWQbKctjx2J4pnUvtZH8zaijSy3CWCUib7l7x
CldOmnffoWBmvMZkt0idHU/teIMWrV19C+u5nxyPiku7gWoe98u2z+iac5cSghJiKRptxAaA+jG0
bjjOy9wtxlRH7ak9y/h0GFToj4FIUVUIOhPqUjSSSSyUaVvqUvxjRrv/14O//cHSM8iQ57KG3gHA
z2yFm/JaJCmyNNUUvelpvbsZmp7jiKlDjkUpBbM6hBPVQknk9ExWVfJrk4I+QUPDf4+U5oGlL2uN
3WbVGak6unY0i+WmNwbfkNChaW3HJIwfTJ+u/9UJJFmE3rNznewJjSYxH7nB/4z8WhpXlPEtpaCo
Drm3IqMlrJzNrTysl5wlTmufAksSMpR6GZnz6JI39t/pHBXO92thRnHK3t2DoU0DSvegvl4/GAJK
Zsht5ffp7J+e3N+MmbV2FAPT+FI6QuvRy5BhdMcpVxNUZjJ6lg9j9GxAwneKCaIRiwMrcw1a8OTq
TmYUBmi8sZRPMK3EHGuXq6ALB5U9cpQ/EqfpWXpHpWzpQJQtm4zC0IEr9ce9ivntth/pw0O1iOwg
VID9wlGLoQ7aBZtG3RIggqVuBo3JbSRVO/VGHBCTRJpSnHXbjMZMhPlJ0pHbosOIGxg8UTf+BSMp
aVRjXO31VhNGekrZU0QCfKbbm7JqKBzXkqJ9FclWkuwPQ1xj/Z+v+B8RXSfKvMCTxiWsE5mgKU5V
kIQh8P9KAgjCS8vYJ31bd5oSq5WkFWROuMs1ioU9aGdYdfl3ggGbX4GlTB6LKoDDISo2MlRXAv3J
5L2lYfkqIxtHqk2Qu2NpeKxq511OXc8/oH0k/C3ufx8VN4DpNM5PDgeajGGK4JLCEbou5g+8//Py
Ek1wDhUUmrIsa2Gufx2mEHs+qg3w/XRpxFn7bjQjFNCffs4Uk8AWoEu4o1Cew09hD5OmAwG2FQgs
Ih9k8FXVifOQPQFLl//mHvQvmPSakaC4n0mgEHAvlvgiurUlmjwsW9i/HkgA2iMI2oZozneHYvjW
JlZETlJF+QtIc5WWNWxDdzq+omBhuxKzpVuG1lGdRgLdioLjP3aYuhC0Y9S+t2Q2wFYPbVPsYkn6
3E0b1Ued31IeARuzH4v9ctWYw/jG40+qesLmlAFPNFVbC/oWXZMkUIs+vTOoANE7gfXXdwEEXrmW
NpIdeo6KgljEzW2Qq4fe7obbqUHFx7P83VUON3fvRjjJX4NBCrPXEpJyNrWntaM1smmuVYiRklUO
EI7CI4eF3LHOZme8G9jw+tworRgCGs8/Qxi0jJdx53kyQDZP7dbOOsxe3UafOVHW4JRn1Hg9hIHI
SPiBtg/OkyjisCYs2HV6UmhHgpS8+RMUc5O5k59Q4JdSj/OIn3MusYh8QUtVZ56P6ubsL8yx1la+
pzCnQSQovlGbxRedd7yAl32mSGqFVdTZ1VdEU1hK1xolzNEEruKpL1VcIZ+hEihsm+0cEcuZLUU6
Q0Kys+YifY0WdLbO7cDD6u6lGwUdIC+O6VR255cUUEeZdEVFMzFJD4I86S/zNgEe1SEq5cL0hX0W
z2XLU6F+k+2D9f9DvqGK9HbtujbVfc2QLfxdxX6KprYe1QQD6J7TNfJbeqxbcWQLCFXEfo7rjMle
mZmTHycolGfw0UT5wyMtvxeAmBBtdNk8U98jV4P2rKpGKmiM9YDBqjw5iD7yooIihAG533nI11A2
E8YsIFZakNqMKnFvFMVdj/PKz5LDfTc0TAaMl3dYV6kbVA18TN9q9jcOj7wOf8pDAZZubC3IDFz3
wVU7qvRCE7r3K3yijqXsih/7mlQn0IvQhuZ2wXBdwTYhYQ63+a9M5P8obJO1fMtpvsU5mt4SlzCJ
fkLEKxwh1u8lLs1C/34tNOSTrR8epS5IuTWIwVVamOGy4aqCH6aVvuPsazbo9suzA57U6eoSZIK1
CtC7XESKNA5T258VM/vjjg/F+1df9Ysk8lWu0wMwua1QRMjeQg+cY0E+7Dw1JLGwbrXsiSZfoKUO
JUczpQNFjKFjRY9hr8KadUd8kGgmB1OrFIDqfBSn4w7qxMJnMZ158I9OK23z9DamqpeR0KJ55vTO
vk02uQBPTw5o9XKuFkVInN2sxE1fVzc4CoZ4Ga0SerM8bLmYQnatjWYTyx78FgOWM+CPXVfZ65cw
3+gCR3jAo0zpn0oN7F9Xy/08rMAK89+kpG+hI/Qpwqg89TwBxgrmx7NEFJQzhOuHu2SYda46wN6n
1EXwwRR8/Tp2jdY8fB8UKprCrLrpDjzyO1pGuIjHs03UC7qfWOycPPKD/YNzVHfJWmj09LU+yick
AsOnNMzDa75Kip4nSpt8ANhUqQFG+KlrC7BqZoT6GdKCfGEjy0qxQ7rHzfi3fahxdamKnb349CX8
u51fbXzvM4slvmF+vWwZ/B1pU9cgrC0iBCR5k1knr82bHI6P8+b/BQv+Qed7VRL1dMm22pwKlAYP
oLCexGSPgRwicVuO7yKJ6hcttCLi8LSD3e4MdZwzKy0gJ7hLG3PeaKjbX0p78AOQQIzhOtjqWMf8
jH8W4uKnIG8w0jpvJ5WUzJCMdqiOoA3zstk9uP2rIi0fpW12CUbXklEF5Ph8C/TrMCXzUM+n/VGu
GHmOKD8KPnOeagOMmiaAzjbKBoiBkyxuIqKGRO6NUNKh3v9Dj9808nqL4esF8uMDzfsLEznWFtRk
9kdCTxEPuqSPiJJ/ShzoLWS+n7lpKE3eiwJLfE1RNjdLWMVv41wsRSZF1dQ88oYHzXcZK5JCeGkI
VFHyjlqGZqk+QvEMehiZNPJA0kWcmYMi73yH5MD87TQ0JD18xoIdacY486HfVH2jbtYVQ/R0tLvF
MNj0Fnak9gz1TrAnO2K26O5zBSL6np4CbezpG+d0xBdg+dNKvAh23gCLCVxsaZ0jpBPa8x6GoXFS
QlB4PuIIKCgaWG86IpUWq92t4WkWETzoCNaPJQj79Eoaabv2QCgW7n558dXuxaksjTE9ZTryRBa9
K4ReFKZzRed14cGYdyWwSFbl6vZ9uOLiao66jYhVtfPp34LtWSaWc3BnptiCwjaMLEQMQuN2Rpjr
dfTa4AK/ucmWGORogtF3MDazffoJdYfARBJlsBajDtnTwee/0EkAdn6VVRexbxZbEH+BqQ3sQaps
Aecc3c3JFFJorkZfK14YojySpCph0IOHYbUChbFYj8R8EwF8Ie9RlGJb71gvwEPhuoE40Hvk9fGe
Oq73KPcyYHSqn589/yXuNkX+JLjgYL/otkvtZ9GX6h81vuSX0ByHd6C7ha20IGyv5fnGFHwBcyYG
GKE6Ghm1WupDkCgrPwJPtDsXDS9+bDYM/HL+b+uml/otW0jZZLO3B/pL6FhL57ImQ0n+AuAsmbmG
OtcUnqlxvPGNsHvhVGy8vqOSdqhqqRtwqwiXJIsoQufNan6lAu2ZNm3L7+knAyWtFchcI13FaoWr
0550yx035LAwcgNCihOzpWlnGMi2GIub4+tzrK60vmlLao6ftqupXqP8YZXVo9MgvzUJ41Ta3xsh
r8nikzG+O4JQpPGn6/iHh9kyt25X3r5dwd4TKDVehmFyT+52t9buDxebJbIaQB1lcDB0dj1VHsl4
kNHp/XFAJ9shIr/mzAHHFyBEzA3RH3WWKsRyXDa7kT+8Y1HmLoTiLYRlh02L51rEwCJ3/FJ+zpPK
LcjeYc0/SwhLEPA+tj+lsKwQ0Zc0uwbiJu0Bv+GP62H9MFudHxHXyziKrExNvIjZXN6cBZwv2spC
0SIXjekEyVS+mwX8wEn/E+AhI6/rGHzkuW7VgnRNcysvuKlW0/WTXtX5YEGFbECO3tU9PLQYQ/Ia
XqJiDLXdOb56SV/1i7pPYOSk9A/kGW3MnxoaDHr2bfPFk9CW9FDSA4j7daFAednrTukvPlHQcGFa
NT2NCsmdX0ETWz8Z/65RcfWNo+Br5C7kUG/yFxsA2s8hLl2E2bh38sKKEIhh0YT5yFIiTOd1YPH8
wus/NycIyB2CEgawJeIsHO+6uB9MzADK6lmdl0c9qMN1dAeKLFeogsSD6x1CMKRt5dhBXJrAp38Q
RtO8uec/nJCIoDbq0B4IRUK6qGg4z9k6teyooqdh3UeDB0BLLZ5jWN3vOcajTSQP80Agb+e7FKgC
tuMqs4qbrYgEOjPg+WQMsZsi64Ecl6r7gkY9zbzGiUKs0hunKHDHtXxooK9N+F9QaL1c2MpzXCDZ
8UldRNPmcOQlgFPkuln/Vgblz5YQPYjqKArn5dJ0YC+Gp2nHfhor+OH0nM4pyB0f1+U6fB8b8MUV
awE9SWgT7neuSolpjsczO8DjpHxEFa3ecXPZ8N1WZR0mEaIrCqLEPyYXUhSoegwGGf5nbGeqn873
xyQtL4z8urmahRcuq4j58npUGPH7ePRsN/UBW/GuF/0hOdqA6Zsj1SUI8IhfFdOxJ8uQnnosMUij
D5mVN8IgxDjjUW4Suru/0FHo2mnr2zpA6XkOz1kvY57enZjzbBhRkn14vevo3gzeEX/Ercyo/9t2
RTPEdsSgmZhAKaDaxfWxE26j1PNwbSFLU23whAgHbQHVToE05suQBgBb6FRsIZHCuVkbKTAI2C9t
MnLTccdalT3eoeycbTzsUMq/j6v/IKWoOPlY2TPVKYVxdbxz8crCpyFBI5GR6bQBNOmfYGMNdX5A
/OoUP2XkdF6/RdZnlolQN/KQ9gBARE2Ye/xr5bZdoPWuzxinPWGd+bE3HyIE/7PIwYXBA3C+fGdy
wf9hrfrFFDCxh2Q+c4WACKBSNCqLhORmQmURThZ5mt5yYDQTNaH9KSEXSLSJ+J69ZCYKhqf5Jl6Q
m2LNxU7paX5V2AyNxSFgnCegeWZcN1PU4cSgBLRdwGSLGm8/ldNHpBxfgzxw5aIYlfgKiUgAbd8T
Ak3LY1ixbH0ed1zazI6a4o8Jwz7aVJQPAl+bG0R4imZrZltsb1mDPVG1Xedd07l1Us0r0PWWVK2N
2XJ4arM7siYytM1t6DhPCokQjJu2a4A2vmPn/pcK6+q18AuNvRf8AfTKHhS1iYJV4OFuCqLRKQfX
MIWVO7Pz29K2tnskY0HWGoZ0AUnJjCs/JNhjQoGN8GR/sKg9sD/cNKadqfeLS9AVtkDvyOawR5Re
Rpni7Xm3AY7qRgWDGpt01dnKgrpT+VVe0x5/18fusFC1bRe4CczZxUkVvIb3dP1ly9r5FI31kqi6
5Xvy/EynFV+nc7fN5aPRqU/rpiYT8i1bS/shCGhIWhby69bha7n+1g+drhafaXqzNkvT+MqgJbpx
LrJSZKrAFatm9lQEog31QKrobPcoIYcRVIoMmvg8nSIlfCW3h5xQW5Yx/lv7etdz0UNWH++rxt0J
b+E16dOOhPmfa8sAxFci75b6lyhDqel/rctgGn1ggOf4vaOjbNwZU0wowvQrM67LUEczz2s0uCKM
fER7GYGPEJR5cxoGoVX23pi6FNjEKMJObMRULDMvfumC26i/aozEjQSoPeoppt+Bym49PzfRlWD/
jdoCluAOrjxdtcfklGZajbjM630BQoSS6zgwRd+gwfLB51Y2+o3KoE+3ZIpq4jjEr0IxNnqW/SRt
aMa3WiSwVFBHOZ1AJSQ0sHI3FPoJJVPi2sg6vwjP3zMgxNOuVEHr1UbtuT4y7Tgv71icj0gyNuqr
HfA6c23KGwr56R9jdHrl+u+KrzhQgldvqMWjOpSB1DKPPc2HFe5hCEGk/4LwGYB+fkxsC8qApt+F
47dM+hh6/NXEVyqz5D/eGdwrwIIHrJ+YNPZ7QdxcBUigPWPJGtuAUGcw8wpQzkAZzl71UOh6ocig
wf6R22vtfx2OtjUQnSQjHdiIHkirG9r26sRGK/LyZKUJ6O+r59dZMP3siWYOJzID/26Mv/9glA51
HIuKkSWPWx6VAl6iuSdOg1/NTvzkI9maF00oSF/ByYfSfyRFcJHCLuzxRIZw0CgmVWF+baZqOS2U
6/VDiSuzdEKxo8JkYBzacdlzelOnYPlIkajaSjcP8r9JliKXoiD0JSg/0oBrJvQtwSeLGy2BMSrv
K9fN5orZSLyHvdgtY9rMEbutsGKbGqm3qgqBfQM8hY0roH3G/8JKtvsc5GciaS1h0X/RMRGv99p2
SJce/WCvtEycyZKsM982kj/xNvxriQLIm3VE0H+gEPNSk0X0izpU+jbdij26q0yZ97BR+Mu44l4q
RGaIUqJk+t/A865pPneaHHsuHIAJzIHDe1c//p0fQJAX6ODJh5NsaVnLPptXHE/NBKrLwJhMNvTs
uHFKxmD3mMVucryOOhzecgRNEhlh9BYOBV0BVVjOfDrHWyAY2hujemWbPvow8h2cDrdlgn/yV4wV
i/qhXSa+vWJ2sStwjX0krTo4j71Swg4JFvK8yYcAFzw9zVDWtiLs+Mgndmcqdw53bt9/NxUkd+t2
uCV2pH7tJBJZswBuGIfqjefDWyKCAvEuKKBLNcvwLSpz5iJmTZyjDdVXcxk71uIUTAWKDGflvCN1
zYu/I0KMDhBNKU+Ipai8WEWI0KFydFB9OdML1XnbQdjPrLhUlqj1Y/pxIY9fjJKjQpWCQQ67wU4m
Utsi8osnjudJI7QwEt/Np4HE3VApeZ9B6np6LbsmDV5Yj1s98DrFUv/GDTyOj5g5LLIr7sxHdZEy
oeKhfQIiwc0Zc4xZesfX0rYHhwkNo+/rKcviy/mbuSqEofuWbrDSGJbOvYwgLd5Dza+46QhFZKn4
aFtwkctkL1BHZYbgl8eboq8bePDkInMObttOiqtwaXKLcE1amPFUrsUmDFycJLGAUNtCWFROR51u
nh/hJz+2auql1xrhUBxwZ24MXnzbYw5R6GCjIxUe7UFImG4Kya5gnYBgJH+dMuIL4wMdzEnT5ZMe
00XXWoWd2NvUxfsswFQr6lg6WbM1t4og7HF1jJByQJyGldWclONZyvkTIBBtNpX2PnekipGh4OM4
kxWByBxaMCvCHk0kfux6yuAwUPkmrnctIxDeu3rw3zJ694VWrmo7DcCv469S2hSxR17KnUDTEZY8
0OsnK21YJ+OFYKFigPXLGlZAULiOim0nPlYlzR6MleJ4FxYi/4xblTYqQ1n2mt2JZB2dS6zwsYhs
I5M0ogzR7UX77s19mCdYO1mV7icMNeKlYNH9o9ytWSB6WhB4t+aKKJ1/zwzvoArD0T3pQElhRLVd
BxcABkLOK9Asn62ZDypK+8jYlEYkjREZKSeRgFH/vErPI6T9hNsEmNiEu3lzZS22vQ0yDY3SLpGG
JJRBhnT5vRzCmuo0msaF+ApK8tozY+W37b9E32k7UNWsyf0zj9N9LDwCaa7vNrMEEwoOkPZgwTiD
UeEsY/YJ/sTsmooX3FYjaub1jG4x0GRK1MUtXfZTPGJu0NMi3MIO1lD1v3SiRI9RTJeBsWZBhJdf
O8UKlkBbkszYUUed+pODvvVXHFbL6lxAPTtx4rj2vIYTEklf0DCpz+aauvExSQ+AJ+G4/TshpbAQ
rwqmGpUgZqVXvmjV1qwRL3WIccGOb1hDS+iwaH4TMKfrzjQV6Rkflc+hKpy1a+W7RBQMVHE2KlHv
V+BtD+antlm9FAbZnm5swzbnMydMGL4mw6LxFhLVm+ZNJZ6MVRrXeA6u0Nk0a9i+wsh5llJyCE3k
vpUuw7REvxwxz6ihZj0A3ESld8q+8ZNAZyasTirZOPihhp7IW0UfSQfake2xIjeB6dnVxD/OB0VC
jjyjXAPs+A14iw58Zdja7WLW+h7748H//aufUBw77IA4JKfyTQtX38oYF81zGf9GRfIO8TtR/EYs
fdeLdyYNz+1xVTyKT/nggX1T4NC3dRL2yLEpAlxGmzFUfWDP9ywYdYwFMiVV+8Lz95SYvYPxGU4z
OtaA8g2A1KNa1PBquqKmlQuXVhiGTTqZMhtu+U90MZQy0rXaEz/60sjhLCuyp0wpTNMfeH2abfkt
aGx5C5A/I1y2FxZJNltYlN8LT61SC+IoXrwl8pd6MkEcc5oPLVd2naayftuxavB2Jm6vxNXd7Xc5
QZvvTWC/izm0jUEe9lbpZBV7DJHgM7vXzIHxxBOFHDy/A6vqeSSpewcEWoAhtTZa9gI5sEVhUrI1
MxVpqL+nmb39UqTB45Uh79A7+clYOvsfMT8uDxaaG04jhF6ztZTfRG5J1WNh0dRQ75JvDZJotwCM
Crpao2vuJ8Bxro2HUD7ehMbuhntKpn1yrHy2dVWvxVKMmA6rt6Q7v4L+sQORl0wtWq0S/WOm9E+T
sd6mTBSOdt25az3ogJ7GvFgla1bAqFSJK9Peq1FuNju80qgfly6ssar9GWB2r5aLy+4VeDRuZYDm
EK7U0UYe6YtgAXno9bj6mh2BH1swyvpcSPUfrjqfJvnvDGZXfjKb3cIqRKg39VCDcZ4MlFy9bLtF
DkV2YH7vNQBzFQgwShTsUW6Xv+6SjnetPKlqSKeQ9aCS6SJVrauDnKJFSzpxBoVJdMYW2pzZLDUt
333yRHz4yUVp4NFGkcIOvu3jTN/NrnF3lzYEIJRVZT+WYkTFpxHeZM1lP0pJ5UFzBbLP5KDGoiIs
5HUZVSvdYiJhDG4/l8ZW3mPpRT/drcBdVxjZAXzuvk8Bx5PqSW59q85xUCTmvVHUlTLfNVFxj2F6
iQCOhFa2Lh/2eztsqbp1jSmCDSL356TDlTWXsD7NMI718BexibJQK1KTwCGaNotkUIXKU9AYp9Ep
Kksof9bY5V206rCPQ+s2FmAEaVpNKXRqgeHmf8UQ4jSCEc/SPURSYmjP1ocibtlABQ/75gQJcnty
jZaR2CaN2qWUjSXiFQG39gFoFrLMyWDb6W9uhJXieqPIdVNf2YQPF4eI5avYIadE0JQQg4B5jjRZ
ptd8dXGFRGTZHToaZjdCUgz2ehCngA/3ahuXcrnUgIrNeQYVdyVu68ApAGJBdCvoThf1us2tQaBp
5iBpwAKj28EiDh1/KMahkW6NnzwtojFVCBMUzMPa34ft927+858FLIUvKFosULsH5vjC6y108HZC
Aw/LLY/fNx+i4RlbMp4WNDFsdiosRn80NmafjxR/QdmURKjtZTf/v9LLZ3qpX0Z2CcWuZk3eVryK
TawCCqQ0e81Ci7quc6XA8N6lBoiL8MLAaS8xrSiB4jwNvsCCFavV8dmWbMzrLo7LJhpTSYVUChWc
JC93MR3da6PocKahtu5pnuUjAqUYxY88yzZMzpNAHMU6M8WF0gIMJjHmeuhx8jWcPeaeHETBahLs
SQ2VTEJjyf0/d53XdWYurg+W4FlkKi0uLGvLOT+rWaAogH5bSk5FTwgOG1nU3efcAmjM6LCC8DHe
ri8fq+3Rnb3U+iF7Rr/CVpjRUbm+3r9E1JJeVR5TenQbBCROQqG/3ddDehgcGop+ICzsN7wyFvWP
wdekW4dcZ6MIYc2UcTgMw9kwvWKNgLx8bMTSwwWYZbwLwlE7OgP//6OcUdbuLUCvJp+feety5+Dl
wPfmjsoXomI8pNaKm8xXgx+I//DQ2XiNilxlpcUGJj0fh0SbTKcAVu+fbDSwZoFSaT2J3weeirad
beUcuIsupcuMXeGt9tEkIIDdv/yLshpIa4OPEkfWFw81e6X5fWiCsDNxm0yh4eyXAs6xOg9Q1HGB
NFReb2VcLJpE320uxzUDrq3QPBsVnj/KULU9LJ1Qc0uEgFVLanDUFCCTieNniQcNLo2103pteoTp
23dSrg3AkcasOEbhjfH1P2RDNt/EtmPY/9HxjUS1U7RCfNj+X4cSb9w5AbKVWrhngm3lmY86cSr9
OA8t6+FsU3StIuQ0supN8c93O/jUulEdPRMmezub/jkjsuAN8lJZbw/bdWbJzDL7tqbC0hbRMvp5
iwGNC4+iszAz3TCyCZWhKM13o9+ZJDhgEA6/tCl7faX8nFZ1fvXjB57RhPJ2RgmuTQAIDStv1Rt9
/YXwG70VvYJk9XEeK+twED89bqEEo9vbzGs2TvgLrGSRMnOn2PVHyhn0CH17GdSnAEklx8/VlNM5
Dh74hNDV8VVp1k/dAMb6b9YeWQ1WgquI379gPYc64Svd7bWFJUbt9UjGB6nNwb0Jmchn0NLF+OL1
DKTEZzNs0sQnLDonM+ryink6LJ3funuwjWhrsn7RUAzjXrKFGgb2O34lQ6Uxid+SpdXQrX/BNBab
a2GkXs7FF/0fMybq5VRoAa2t4B8jUx6ZllJf8dB1AMG7UMEirOhEhKDueQziEjAU4yhG4sc3TEWC
PO/yh5M7QYOzbWdFDpa6xOSwZB20mmpyVaXbsp1WyZ7tVisH+QnOv5LDNGiL7FAB8nX9UVtSZXch
7+Ee08RhsCqKAqdg87FEfCSbaGfWD6uXvafgIE+uNuLJfZ8R26wAl2iujRd0SNh+8q0RCrXxUhWd
OtQ+DjhSMe0xUlivFHe4zDYqHspxXvMeJR+TbMb6ykrvi2V2YQhhMzo6rQcOLqDxuKRnvtFqOXs3
AFQcFcvgEncZ+okzzOoXiDsyiHdA90ElBOT8Ypmg3GT5ABMsYVQpYkd6lko/DyULwRKcewGQez8m
f3rtostxDUPU0RMBSZ7qO4eXfGbPT7I4JQq5RtYXyJGMAQZ+JKF+b/Ho7w+6c7sSVA2NByD21/C8
yWSmo1z6MdOKO9U26ciN/3D1ab+08x2fMYHmkkE8SnS3e+hfC89V3Yo0KYyEgwkO/W2cSap4mxKa
w0+iO8xE5kHxaNu7zoyv27IQWYMAkptrUhkioY6tHUuLPUz1Me49hSG12mvqc0mZ+bC+20OF7R6n
qlZh88XN3uS0X4IlMrlfddPjDf+ztcc1AGvFPlQJSplwkVClKI8BnvCRLYNwO64kTG+qWcdQRFp6
q5q5Tth4a5eflU57JwgVKBHnCVjoaz8kB1jICqY3T0tLdctKO4XJunCDOWltTuT/AnL/DrUvmCgX
NDDLkDnvf7St+mLE7ioV6XBSTBO9FeFKChcQOeQ3l+T/nbd/XySKdzB2CWnDMwqT9jw0LFnz8G2C
RRwLdpsbvgXIfXneS772F4OVSMqpgl4lkskYQd8TxhrxfRAg7LASb2ZSCoFDRfTeFI9ej3kZuvaw
3C5P6NN5ZIh9+79+XtvMSLA9dXfbr510BMe3YiKLktDvDQPlMVf4icb0R+B88wo+9a53GpqxpymS
VTDVGrh2lzQTgrPoZN55UP+Du4e+7nv6IHYgJOJCeV+sqilWf4orCrjY4ALZL7tVqYI1U+CtO2m2
Ifj1tCLFF18W/yyPEMUraVGQ2NwhJlJgylI0CsXrjIhR3s/nPqlAVbZcpMQurSZA8Lc3d9OEa4jn
wmKdsxtR6iHtzHGKOkz1qkZTKMRSUw7VW98REeCAmJ6xV9vg3DOqIbCiC/zxbmPnkh/U0PRrlNTU
FaD3cAIZbDUfip+HflLB/vXuUkaXFsBarcqRSSgiMBIiPqiDkeM32UhvEoNuEsSjHZ/h7VcFpdX6
8Sx4s7neij2AEdnCmR7AiDpBAO7txVflAwdBN3jJPocto4YxlNyhA/1mr5samsuPkQHbEyBaklKx
St1lY3aayvu6NrdA1LAm2dxApzgGLRDmXfLAH9S8HwrfFxoNgVOKLDu/mGs0ns789kEy9r0vIBEf
PADwtwSH4NyEyTzCeOauGuMaOpHNEXg2MQPFcc1SUIHI6ONs6GDuY+w/j1xHr8/XcxqX6mK/RZlv
zAjqd/R1kENYSwHEORxXz8v/wVNvfyuNj8rKHVEm36i6x6zATqKMn+BIeOt8svNPs4oBUy2RulSF
0uR4bQ0Akk8EtvLdutSG1TqnWmIYVMdaAe6fprD87axI7CY6Dj52ETzEmPqSRu6iY3/o/XzeujYR
QU+q6dOgN0LxClxjDsTuu0JBpZSUGli88SwlunwtciaRp2xtQXs+t2jtKrNRqWqS51bZBhdRHV2T
hiVBr+xgXdOdOx7RLpd1P8UXdgf6wmVrpxe6NqebBp3vGvA31noQ5r5+AvID9sVq0sD5KHoy3XzI
ufLGjhv+BCD/bVjrS8jc8NNerEO6Cd7Ktb1DGgSl3/6jzSqcqamniA84145YPa7Q4QJo6OqujK/t
GJAUOWqmJDQDFy3Mk/8GgOI2pcb6HTx1i8hX+DUkH+hYtQncAWmO0kjSmNS2jg1emUJll2OxWVTN
78n8vl68nNlnAdW2FIlkqq98osr7IGfS+qJ48XFZ3F4BnvMTKxrygGKdzDBQ1gQZ9qU0ik2huN+E
VZu6TuZD0t1hJMZkXDr0rl4TwwDcHMxmWrfsrSOZy9BQiR9lCi9sA17ivQPW9ULP8nPMfF/xF5+J
qJoNqJ4sVun8CAJqfz8E0C8i9wQYKCRVKzjg2gFkYMxNdp6Aslg0TDDmXpNX+LuU8Hfj/0z3JsU+
z6Sfc53rU3579fc3FeKiDMpBQttHwF6X9j8ncUnuXM3AG0AiKysvp1RmhItQnYWpVezKejU773tt
10CIvM9V7AgCm+frR2OKQHIaChH4vCTvie7v/jWmmPF39UlWIeLhJRAJHvu+Fb4cax498kY0/Bbz
RcsNQFpmKRHDYeBYun36cAHszfTye7Af1JqDk2CaoLrbxjcm7C3tYP7fCOuse7wS1AnXMbVeYNkw
D7CcsvDKX/lJOSlrIcAOkuRAQkB59o3V+yb8YJTpxxhCxgRNKppFXVDsRKr3ZUeYX+eLOgkQquwT
kd/ePhMNsKlGKINKXpJolok69yWJpHOUL+n1b1gHy7XnPIsaJpS+qSqApGdWdTKVvHdzJOofcjrv
QP3d+RijIVPYhHJ2mGPJObj+ja9grTDOC9BbA6S+L6zsfKynr0gwvlNdvLWWP3zCJpO1yhq4hf3Y
Plrqfj+Eb12hhYbHsbkt3ew/Cn9CKKJM4iMgt3yr7QmsMFXfozF8mJE6/YOpo/GT2jTY7pLkR4mk
mpvqvrUlndX4VWHX70kmVEPEi0lNHwVLFG5zb56Xb1LRARA3TKUKu/yneEgPDjfSuOqqAdkjCDEh
tCzkhSYMOV+XlBQApRsae4bJkE5C69NXGNtpUoogXzVpqf5tl8wheX2193ixaVru8rLTN0OVi9tM
s1qAbtVzYxJ4qoam5G8RmkDy7usATTrgSHUdpuXj7cVphpLwhEfT1mjtrSF8KhBcOpnU1FxMQg8Q
h/Ifjh734uGMktJgxaUHb7jAqNfd0GA7vneZG5krMfVzv9fVZboNgPk9w/T9PJNzw4Ar9l7nAz4C
Pk1iF9bf1pu38HoarCQYk8fp/jLT1zRlnQwVKYhhMTzdCEDEEtHXYdlLi+vlzVugRtTlFpcWxEvY
dFpBI31viIy9Ith8kEVwSgrhoxdldK7N7h8Icgi2bxP2MFSfuft7Hq6h9G0waWqRcp8K+4roZX1D
XZL/gNp6Km7Gl8HXA+nbRN4+fnjeGlr+EG46DaRRavgb5fKMyXRqmkpw4F79cpkG2doO3FND0cFQ
ksAW/BHEUVo2VHRCkoOziGc5XESJKLhj55DXqCH4kiMp7lkI+mI6SJ2cdlzkoUIJNvCCH3JXbcCY
UwYw3DzzblWsB9zpmBx6pXqEIY8AW8JQ4LGRs/eLWjzsRBksil94zZl6HUE2WDxZvypY7UxNelZ2
lsuyJi4BvOH7pZ1DrfOcZAnilqBJASEBy22kqSvaUkBx3Db94RDPIr0X3HUiUdBdoTkm3oHH6MhX
JvtG6ZjoxtvFtBiCHLwRG9VGWnjssNAcXek4/xM9LjvypsRpUaQn1muQUrWSuF+W3wI/cJmhZFOp
C4XSWcLb9f5Op1hjWvlFLXjrVitX2rmJVwE4J49+4Bn8MKCtJ6gqjmQ7XwBcrLbp0fKB4v44pOqU
Uw7uBdLerni6qtkJjkc+JTSTuONtTrFPnT3Vzot/z0X5WFAIEEju+n5gIo+OoGMUxF7UUe4KP5L9
M3c4zGmh9+pNNgZRddohhLHRiE94DJIy0ewto505fhEPOspP0MSmzqUhN9jO1KLkurOdRHh37PU+
aqVQ36MFSsgb0cm73Vg1UcXSs8ag9AWhA0QGlYIvqIYHtvgzk3WcNZ4h9yK/N69IT32rTjKNJodX
UW0AXKOpdGrFJ5gRl5ROXss9ZnrKw/G30gy9wzdXr2XXvTlfpPqijA/FDmBhMxG8QGHgwqtlgRYt
pP3jT3Ki3nwzR/TJZ77ZQ9Pc4UxuiGZ7UOkgsM804UkpTalzcr+0NR8wJ0+i0VNkUS1w8hpx0Qzz
9jzhzMcoXa1xwaSnnoQgh54DndJ6LieIS7hmZ0t3xeeXqWKPLdvJk0gAiqggodRh1M0kptyi/irg
uoUNcT03KJGx6HztrzvPP03KNFQK6nedAz+AHeNDnsWDfAl0Mc7CO88bgY0ydKw6zqBSYC2eV/UF
q6QUyVJ2gsKQPeUN/397Ptp6ADryiy6linC1bot+gxvIzpNL/QOvlRg9eZYO/fWc4UFkYDyJeZqQ
tWxDGm60y+lEJNEyuBRxZFajJvNOygOAtkcOWv0b++LdvB30bLlXlQROKGbLch61C2j5Ssqmsmmf
j7y2pms41dFjPwKXg2o/MdoWw6XEK9C5sk7t93PXqcw3K2dpL2naZMpMUf1ypH4+/uQw3OlHNSo2
Cplm4ak+leEIrVyeFJoW+rAn2loqp52rNDZndFlf4YBHlm3VTiPQ6n4OV70oZnqz00SM/I6BbDJO
oP6buEmXr45Eu1snaMw9j51W6LYJtR71pg/UXjSos0gdWHVL0nXneQGnCFk1B/+0Wu0faaKldKr+
Mh8E16y0w6xWLP5WpiQVr/rcxMJtwzN7mOpotgen1G5FVbDwOs4f81+HV98M761OYdO8dr+fuKX+
1u6CwpohySHMY64VRXTo+nfnjxrazBzB1n3JWhpxKWYTPoWxlhi01ATfC2dLuvEVzGguDFhJ7x1f
xFqTCTdODDEuHMXRjJNEsr8mG+4MkjakxiqL6KVmk2QDqoax4STxiE5zv+PkCxacEJT3JxPKeZwc
096/SGmCq/1qmrDWEQxqpVyPsFkKvKNtnAuuApRUU+em/vD1whu0ffzwbqZRzD6HxfLJzhdTF92o
jhP/kzIVfM8jw0nWdQ0hxEWMpTkNVsyiSKFvMQqbPolhzO2KZLkz6iUTRtH76OfYQ2G0RVrOnjSU
duWe5C/FMkatQP81RLWqNNw4pXbbEY4jFjsYu59SQ3PWr/NjUTs5DzVNtQC14VcZvlWYEzgyBAZs
YJRmQSmfLUZOEA1DgbZCGOqvzuGD02L5+vTC+oOj1anmRl+H5eknwOaLcKf3DSo0m01+D0KgjnBM
QIgwU2XxwTzUMY2JkkTF0UDqzo2/sE1FcJ6VHzq87jLGETZaZHFJiPLJcZ2yszm8GPKVPL6HdrX9
hWQATuGZZx4kcYCt6bRH1Qj4byTdPeoe+HAboXRP0z6j577PbRzB4BqAh4vQuzcPPa9pCYWGjJJ9
UDKpE8NUrSSkEaq8NqYPKiSDgE40+kir0XaAjUuZUAl4T3uZXp0c3eqXpxWz9Nv0HJUDoZ9HF75S
NBNoKhC/doPx/T5cF960Yml+VJ+isZdM48Z5zFOv8MiOTWBQQdU4lzJemigF5gw07wJWUBEnsjDc
oTuXTu7IoelsBmpkBxORgtfo+97DZvZE4eX7b+I0HtHE62BH
`protect end_protected

