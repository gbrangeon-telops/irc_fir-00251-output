

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
E82wkdGPZb/+6GZoDi5HpckkoDtuL8TGRb/JCIEDYKunG0ehlHY7rWSAl7AxBVkDytYXn4VY0NY3
tD816aZ/Tg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aN+8nTYiRF19Ga2xgugxmmkjykOIKDSAJe8CuGlE1RsIGMA/TeZJn/LIOmkC0L4RXBBy5zkZr6mC
39gWvg+KhH324/pLiKCLqvJkIObctxdk1QghQFlwGyR5AgwumO5V8XR0wkFrGx5lcmF5I1Ic7QCL
4FCmeVtU3m0TggWFC7E=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aDXP5DZMSmAZ37R6bG0c2an3UXXBQ9f2UcCbZO9jybJiEbg3jaEsz9OP8BILMEuM2Gg6zqGospJo
IL0GjwnUkhmqiXNrUyuU2ZA9j5Qfpqi0cT39WDwUPJ8gireHKMW3Lk2XSOOhzAT2gL6kjlBz97a9
e5WZk5XJ4JpzHsyykVOoT9yBzVvTvBYrbMxRFsaT4GZ3NCp2/bL7FcAdHRGbG5cNEc+P//C3rwO8
4GNkm0wKVMVQq/2HclGOKJAykNBN7fGuG7zIF27nKqnI3IBVFzw28uEsxwVFMpLMQ1Amv9lQcw/X
S+F0+1sbjSvaH4de4WOv3cOUzYKQ/wzN6fSahQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c+SPO+b2cpVqItr9nAdAKH8LRjqZZjyv88QHjXDKD8kCd5SL0IXE6XqQ/EIjme3B6XJax0d6vBvr
92G/L1QzXOo8P82zgbpcUFM1hqtYFVROwwLTcIHV5QmMcqgWTv/CxjwYFY9l1w/ADUzzHakm7vO5
G+sQHpPE4aud4403sjY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T8GeY0or01NdwqMo6UKJMUTsmtP7APuN0oCIY7KzFu+PsK+FyNTk9rSPzJS4j6dAZuNV0qTymCiX
Xbb3asOZtqkbmx9Ts0TBudlU37PFSlhj9aboLv0+uBJsltC8lWgypATvI3dldUNiHT8HwKeBDDaM
ge1f8g9YSSRm9Jao06pgbL/b6i2WQcOEh+n+/rJDy+mhlYh4b7sJni6U+KkkIH+Nz+FTmo2KpEia
kiQmZaPY0KLlWtwgAmS9D9WXDnBy7lDRle2NygR7a23rjPwxBp5MqpWylPuquQQaCFWvB6BJrqSH
TxLzvd+PYmz3XQMRs1MJrzzaNEb2P8EXhMkKPA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12384)
`protect data_block
TmVFpU1c6A1zFYroIRwkju+CZze8NmR2WcmnksxUBxTly7wtY1si8qv7MY0PvRRYYdpWSQ5JQ9Yf
yMPXhnV0UzE0fBMeaYCHJcOtbwmUW+UKh7toPye+cr/M+GEddRViDejY1UG9old8J9nWhxRVSPLb
vzwtMV4ayhcG8Cclr1sYzFnwZYtc1yMPtlwi5LXZo6Nbh5qb2Vz2LLmqNobn1mlUkhcc1DaBvDSO
sJl/hkNH90NBtR48OWPg/YTk3y02UEcdy/ciNntQzLELsSaSjSdWQftjKxLzVlbZX56GYIvZOj6+
SUnOcl1oqr87Sy1ASmuAWgG+XBdoK7FDiKZLOaiygoCQdrkIQsZTY8/C6yzMa86nsua0NuZycdRM
s46xRz2ROZJNEvWMW43G0Yjmpa5sga+sn6QL75YrjClVV5ynOaNLjZTsnJn7iE3Lu1Ep7w0awjIA
u2TiZz8guWd1cLYoKpGrM77Zf8GotjI6V8pdJxfvMa2KFbK7HosE9g5Bagk/NGLOwbsuQ2ZACNfI
+ghtMLhGy9vnos+iNGOfVTt2ChezsIJruzpPQvUFqorr2zYkIx4fRJM/8HJqrVUOgGF4pYY8XtCR
s84bA3jRHsk8RO9czGJBqwAFds/xo4EtVN/NPi6v1JcfMJSzTJBbIE/U0wjdmy7b6QKy9iRNUgBd
ExOlgAc7kFRHGeSq+R5SAeiFq89ckQhLknwJHlgJYbqfhpKfxW9VMB+Yq7YFferiTW++KnXZS6Jx
Ite9hc7FBL1IctiGlQ+L3PG1Fb/VyA98y/QScIr1//AY79KQWPy11JjBnYoZoWlPAYV5dNp7lIP5
mZE95Qk9GnJkwuPVcIzn7Zer5fzhkoAmLQR1oxFZZhRppPIxF2s5VqrH665G18TwCmlxftZiRD56
eNMRHvr+IfPEGQF67Gpyi7GgLVy0FxtjxrpOFECMRUNcTl9sABzcQQLKVXkP5A900cIi7IdNPtl0
orcaYB6YLJzpOK/p5fUGqNoybfdkULfaeZLRQlZRJBmeDEBlGrty3H20o2hsL36JyiB7V3Wtx5Fq
a2B1/LrNeDAn4XX98w3MnBVUxy4HwrSfQ/ytJDlXR8+r0B3DEnXYzLYK4lNrABYusDVYCbtIWGli
DbQIAlcD0FtFtIEf0seVkxyjC2dqPBMjLEjucs2OQHimkYKnatTAszR2jq7LoMf4ABZMI97RSt6L
kZn0UrfgYLIpVsXob3c/r5g49nZn8/WCYCNhvniPJYwsPItKrGsyb+1DcZPypPdcv5zEMt8TLAUd
DpEkRi3E+Z1r8uUft9+57iVCMZPRHIFAupgs4kDuQJjY6mTonalJ/aq6sLziGkXWOy3komMaLKcz
R+PJNq4l24x7KXYPX+Yn+QuiNd8uU5hdwH5CetENq027OSdY4BgQZIiTQqyE5cww2m/Lj9sanWaT
j6SXwbMDDvOXS2XqQfyQWuh9F3WWoaX4EdPMGXVkdnKs2A08oS92itqHnLPzDI66IMQswauBRkLS
2ZuDyg7XKAr66uPYPgkYsTSkKTGZ6KH++O0LpWIHKVN/3pZTB5QHkMd/q5e8hl52S0+0IBTN5Iij
BuVamlPdyIIABCcikRtxszoN3+aHC23tbLYAM0/yqOl4y14v2vaR6g/P3U8H7v0eU6Jn+uNVqyEl
izIJrlG8HVUz7ogJtATcfgJXSJO7WTLjTHjgcq/fNrrXJyeCyVgScZ6ORvuiAUMCYfdfMGsHJ+g+
F+pdFbmhpvN2HQE8zUMtLF3ybnrvKV77Y5/+aue9l+UTFztRDYVChPYL+kSn7VChPlV/Peb/+n5z
ohp7LMRa4dTZO5L9l9NiU9+eav7+CA1ncDgPNjfe7D4L5RfvEWW2lVIs9JR1wtddv6jmmaCxVXcv
u9+9xmVLa7k5GXoHSXc3B9qA2yVblRjZEW5s6GO/qQG4qP/mc1xEufLNyhPXbxXieTESjpYdaUAt
aq58Ps1VdKq1mzeH5XgIreakLi9tduh6NlN19WMUo+CmWBFLZ2K2fePd7+hAJwgE+fYy1q2W+3ts
kLYjwyTDFkWBuGhd33mp0JXwHd3z5n/JQl1mcHtqyW0TFtsyEfabXwu3+Xzc7ppMyjfXQZpeiNLT
TI2lWxZGvWdBKDdfjTHwOyeXCee5FIItmlIN+OhjlU4orHR5G9wWgIBP6/1m+TpXMO7WEdZO1Dm6
XAEpKqs4Dk6BXzWqtOUQjr18ks6ucNkTI1FdcAd4eOuMHw5uFxT8dVYrU5jntIb4JjUI0HVutkbq
+okfjvbeArFzIVANfaAzp4fZLGFbXotibCE/0nn4QLSc3kJAYAq/M8VUGpP3xsB2iR0UdW5fB25D
Vw8wp2UX+mbDrIG5Qmv2l10pgiWFSS/nKrB/0IB1KrWPyhtORhC/kPO/FlMy+yRGnAmpOJyQ/zC+
MpR7cVQGXxsfjVLQRSBytSB0McXl5hykytr1GFndQrQz1FQXwkq/uYMeiCJgFsH5UJ5LWUEzfrJ+
kRT8urg+2fsDp00LGlqU7aSiBz05Ss4ubl4nEUhuyAYOvt57ExeW61alYeTqDi5moj31Ap7DbHuz
z1jclBMHXNytWr6Ix3HTpYdJg8GinEbnvxVTdc9swuRUj7yqo+rstWe65+6ZyF0rSWYeZiIft6TL
1U8r9Gye2rFlgjwOzLEWh+GXAGS42vOIybnXHgVBNH6TMHQQGANPg4njYeonaqDL4+4speXyNcVu
SCC3Ooea8ImIk93rVb/I3aXIBZyvFnRVojHvM6nPVqIks4Wd6IqzKT8Gs5YMAoA96rW7XiIzxpcq
A2Igr8hszIvflS6C4ZvYhk5v/kcD9+HYf6jYQgv8Rto0fQjDYXwVukveb5eNwDHJRGACdDITNqCZ
g5GnyzjLSo9JNFXPK+i1BwpqSh0w46d14YFhF+ug/MMYoGdx5LZ1QOItB7z673n/+FdL1c0w25P7
R3y7mqyP/PBkbpO1OZp7r2MxXZ8cinXnbgJGW/Qup2FIHv5SvRODp8cWZLoaI2ij8CWhbz7spQ2P
LfR0Hf9gxKCrQt6qgGR6TasrzjUkvAzaPXHi1YH1pFj65sHhxh44cSfBRIR1ESzFeNDbV0ZI4VbN
DlNGhqsVFZLdujElS2B0V5uHfE1ijgkooLLjJf4YRl1+g8Py9u9K0eSjATJj7PXlT8wFr4YsmcBA
/BDs7XPN8z/si0J4mOaySptQFHoVbek9GMsDTV77OD3S4xspgx6l+RI0u6GK6ewwUV7o7CDzcRXL
CCDb1Dg1GjXJ7i5EyYN3kYBsCuVw1LMf6M/C8wW9LUafbE44aM4YA/edVVI4FvVnbDSYqspfXulI
SXz3sPRXzfnLFyuOYHbICC6JV8iMsTXRWbbwU5gz/2PAStc1g+SUhFzKkZzSC/CRzQW7VEtPL/Im
tNUN3rbmpnrMUZtJWcn0MozQ0PSkTIP4MCaTXb1G8nHlSDyK68R4OflOjhOctj2GwH62HjK3ww81
vqnHvHz4oKydsSjisnuFCXd+7+0+SZneoZ89w5hhOkAEscpsRatvrpZXzv1QPbF00oelttVrrS24
58wnL4RyTfLteASm+Jt1ox1CjIxJvRl3WGj1fTid9JHwtvKBHYwF9kE2VyKk+2VGRsyE3C9ZLCTA
9KM7uFnovbF0O+3gpFQ+Arnxiyfc3h63CIIagN799WizA+nBdwYIFaPD3ShMWwithaUmrw2P3K0b
eTPA0/2C/G3wJg0bIDRYatlsTnWtxF38+wb8Ow5YtxzZH63qJhZYUGPi0eDC/EkQzpXYQjmXUQe1
BobHzefRVBAKutem5HaL9f776GOL+3DKN4h5qg4U35PcbxkeuJ6eSqMCYkInwZhqZB+xm8WryWhd
g7/h6P8SIqLgYZqLVaExVZ4fQuHzXW1PIxj9IrH9rgj8N/4PHPiupRSboa/WVLRVKWFxjGilUMhj
0fUdOiwsNoXSxb4lJjlfPNJ8juq6Mn8GuXSNdnfssKNd+Q9lZvYLJ33Ep0N/QCpys8Db1k5lkESa
VTSaUzUzRZb6h5JDtdAXfCEjF0I8CgqDkVsqQHwmqxrAXA68JlR5+A7+xaEsoyyENT3VhhryEr4N
hoAOjDQLHSCaorYWuiu/xkgcx1nQ8cznMIqbnFdJC+ThAPEOfV8U+TDAn4Acn4sx4nfhbSzK/3Bs
WG5togV2HWAg1QqN6yGPHE/vGoLLV8bzwuu5fCX3kZt609A7eragHBr8VvGzhz78XTNzh7Px+1cb
h6Y4FDEebJRe6cSaa6FVEByUjq+No8jeZFc7vqaVCJ5zR9wda5lMZuJ4yBqZAeCMv3fgDuXmqCqs
Z+jy2EBY6sprjg50UjM1PXY1uzXSuvK4/Xy3Fwc5dedkmCloktS8yxLRqhn9geecQvQ9u8fiT1eL
QN4cd5Wq9OiCtXhzQqmZBQjJL9UBcrpQIKgNB0In/32UqHeOhRifwWvSASbCIUunXUUfnBJ0qLCa
hDtXKEh1T36laNkde9J2bwkWBZbiEmMQxF54V6lGa2lzqjBUFzdLUNhlWvjAAesfko6/HyMAt9na
T7IcPvPVrZ3EN6TMmkFEe/FAIqXJZfM2hcMX4X1wFgbZMX+A0XGj6H/t3Y40Wg+fOZeVzUC3bgI9
jG935pKA0KDsTk9hxkORZszzDhV/dtjcXAwtJXYCdJxqSKZlTi1QeUY82RAlA70U/Z1ZTIYz6rO2
8mrDxYa556lGYooofRylf9pan9CbJL1RELUeExrd7bECT0bQ2Bo2D3RMrJSOK85jVhcwfEWeulfS
ork96Pjqh7+yiAVfa6vrYEPKbdup62aaa4WG5fCJOne20wbDpNVbUXSpD4hy1jp9T/fHrTEqFzZI
9779FAN1+82trYR9nDBIrQ0nEeoEF82wJwQIMA/ma9hn6jPUi+Ad2C3fOCR26cp8Ne1rLEJc9n+5
4dfl2x30DH/F/euYpab+NU+L54A/HNfV5/x+NR/ac4DrFVFrDdlnHUl6JYick8oZR94douYs0KhT
lHYFlJy683PHkCsljHTPGyeKJmm97Hu3qmtSUodnvLSt6WqnWst2wbocQbE0dPqpbhPtjEUtUSVp
ZNSOA0inMyD7zzcgVbkiihOgQUk/sod+oapDv6Gd2WmjRI7Q3/wEwpE1MqO5zTPPA8+sdzRUams+
HDCEHPv60+JyK75XOhO8aGICGlKCutXo0JLBO3QKgIb9T0DOfwVf0llcHbPCMS6ky4VOSiiwOF9Z
vS7t6PhXjdIG6T2Q1WLF9YGe4kinITWrF/iJEXmZ3DM1qJIH8b4eeFTudnV1frydOCLdhk0+k0e0
11LJ/jxvoEUd5yIKLvEllmf7X/rgGLdihzjZ3PzaslOVGOdmBB4fx1R/T+92ibgDJVEblvciFo/9
7WBAYsNqyDKLJLy3MCBgp1ZzpGv7zqLnttji7cckL6SFxptenomuZuDTyXri+XWDu9OP86qRzsIB
O9KmNB8dt1h1eL1yG/dPQh3AANTWTKN7ZR+k4BZ2DPyYX2pkHWMX4LgRHCFZmKjZJbRImtRaZvN+
AcbioBfwY6NLdQSkqeFqBLRFV5liIn7Mfwf+H06CJlafqlkUYmt7Zv5k49FHTai7MaSYG6sOoTpB
H3TVfGe/MFN93MsSdf67pVnV1Jdozhxz1pW31yZqKs3WBXcwqGYEWSGn5eKuBd9PFyTGgIlFrF6j
ppuVcb/Ggck8qzooxQG5Fqha7cdwObV8IcjFWcprkYs9jqiwYj48WNpAiBGWTWmrYqBQ95LwhkzR
nNBf5QU3SL5IR/6JGs3BrjhsQ5SeQikkaKHYut2WAHSNxqaNRIVhu+HPTqbxAquLHNBs/PwFc2i3
ah/gv5cxDYptImvq5fYXBMgv3jEdQ1wgB8/ro7fgcRs5toxUgpkwd3QA4LBSlxmAZxFlRXBYQBf8
FQjXhcUc6cSOZrUqyIhRW5HhmTcOcU7CGlEsU7yXkWSrzuf8mlxWHatqUmX9OEXCwGq3JGnjuche
H8pBIyAumfkY7t16IU5Vgt6p0FAKNm265ktHqE1blkM55mveyGyX3OvKfsm7c1Sx6Gzg/NhZITUG
6w4qcAqZpWsTPCn07mBwLUbdB/H+tqLbzVNAxAHxbV0YXwdsv08sEnImqj2KVWlZ/7MQCwAiUrSt
dxfZPBu7mRVd2jGoH7nZlelNd2MHoOuPipX0YMLULiwCQ1K5GHqjVKos9KUHf7lc3RHIn7JB19uR
IiixcaYOG1U6fcSe/Ab11l03XkeEwvYFcUnJdbUJkOUjgPSAR0oQYE8JjBUYuwHM1eZdxA9FJUNH
qAHHg76kdLi19aTTmvoatWWb+nBuVVli6fNiihC0bBD25s7TnPtB2uGkEcqXb8HVJAdGCQuj1ote
FRe7tl8LEmnnQnrJjd+WtJ1qUgaqeehZdXYjRM9aP6hFm5+B4z1Hg1lvPwfRfapdGAqJbwyd+epY
LSeHYUqNTaR1zHDPNXW/iSfKI5JsDWWQ6gKajm4GEJbQMXgsWw7tGrYK7d0y9QrPc+BjXCGn0w1+
k/hRXRPOeIJ19V4/C+P7TUaLNJYSs2mDQaiA0B1b0ZFJ+OWUh8a8NasWWQzvpGgndzH5FMM2tVpZ
bpjYAfhgxBy/iekcsHreNH3ZbA5xnVaJ7DKxS4UdH9ilhnpAtJbefSilVSeTDl0VgmqmPhYa/rmC
LEx5AdwXWMa013l5QniZxn9NHwZanWwlmbtI+0gpMpMT0Jh0buiHRu3oMWq2DEwQjQKc8WSkac5E
hCik2dXLdSzXaPRGjUVnQqzwr/tsPVAAps9HTuQa8x5Q37+AY/Gxi0WQidfsWHRT468VEQwTtJiy
bP95VFXrq3J1qBC5m3XV4bZxMfYQMVYIdJ2BLKVP1fhfpS0PGP6mZ3AWUbg0J0+ia38LCGuIecgT
WCnJdL+OmZtQxT+r//k7AYtyjkx8RFhqXfQuGHcbKjwj+QKTQPsvjjphhzktURmjzDWRln5w0r9C
dADvV9jtvM1wusmcastceCjKSlphwiL171iYkWEr96Ijn+tCtkSS6CUyr9wzpIlblWl+WSlXaGgx
6bKbctr0IYELhowr8GY6blgSyPlrLtA5d7klEbvDr2C5Elz6keK1Bgn7k/pPG78Ytax0j4tZtl9i
tQCCdTSQ+as+eZozi0TvAB1SOZoLFjgOBUc9PGV6dYWbuZaV94BsC0z0mGUXZBRMXuYkIyJd+YAJ
LIFdVWFoinRlyIBeFwiQVsVpsLBgO1fRjmM4exQb6b4+lgoQwtbMBgdYHXuAp3LeRcV+NqNmw9O7
Wgc1R4B1OFJzRytelz3pDYmpm9M875fXMtyl3Zfc9Ou2rF9aOuStRz69gyE7Z+O4umUixvKlSnvt
OD2r0cdXdGl5mcW85f5THPKPv/wSLN3+JEmRMbJ84DV8a463eGkJ7JKr3we8rxdDREFvmzOWaHFT
rB8hVrhVITsshfsnvpMJcs9iRP8Nnq/JB9vTppRdYE6AqY8JxVe6cuDS0wM1ZduQPLjuBHA1V+6T
U1XXjbv4W+yQIlKp98NpNtV3+ipVRZOgCdPJAQn5khBq5DbQE91Q45DV5K9/SbMUptjQbE21M0e4
K+srFkWNoWTITqvk+eeqdbizmqLUdnDLz52EUUDQP/vGrAffosiTI6lPUyrio+EUx53Gwqa9cFEx
aZ/tjUPkXATunfHZkQonD4mWwfFNqgW5pYnQQfd9ZGyXP+rZuxFyLAqKppBhcdOJ2hZUlgLo1klF
sFAemRAotqxRq/2Yj9gHuV1ivKBdeeUyAQ7zabJkjFLB/ijgrAW2QwfJgkFneDoiVBBLrrkTDq/7
pmS8aXimYbDx5Of253E2q/TFhAcz+rU1J+4LWx78dqx8libm3NoVPHTU52mjiUaDN1HNX5Acu1sk
MnXmgD2Q8iuKucFuEHu3p4KnS22O2Q1pxba1BYnSc2/0CP8k3K/UQY/k4O16Iv7pwxpQyDkZhji1
FhhKgKnafhxBX5MHnaPZ7rp9kRplMte7U07Xqp9d+qH8KKPUqQ9dzih1iHRVHjNNjnHnhJIwLzqw
IbihBjl26k5YDZqSLU/irJYqIlsbSWYadUIcOHfaJkXn94qkgBdVQ/cPp0zbjZyII74rdoABd7ik
q6/YPno+yXwAQ+QCkHeskN8AnafeMmnJW8cdeOYj39ykacG1WmKjU4Dr0AIzIpxVSwKZ825PJpEN
3aCEf+WrzXwvRuOiHkOdvj+9nWmBN9lBJMM9JAGNfPU5Q9R83z9rM+rloXsqN77MX/N91UjHf5T7
1TDPvP/4PCLND60Qy+FN8bIUJYlPCV5uiMJa6lN5JqXmGD0RKuYpHHvw8q7J0ngWMthjLl0+Kr7h
cw1zB/WdpB7+Ib0A5ByqI218KEYm5RgGWzxP54wOWonThWNMwYtbend2aZpqJX0McDmLSio6SGLu
TPTVq+5+rFKmjf/iY4maORiHa2E0puIzZ/lNcGJQ+d/RY4SKzXVabqyLBTUlYG/C/4APhUdPJTQc
I24o9px0/SxQlZH1qSzum0Pa74nBWXVeXGp0bv4Sf3Ux/Zz2u8AHa9BbEq50inHVqkpWkiVIinuq
R/21PtIZHIDUtBeRckmIDI4R3DyAr5ZhTqcmStnkS48frBi/JKf6aIpRc2rZwW7+vcsUIkijuBw5
GmWPt1OZgRLjRqrKRtt2D+VvRnLR4s91etJbC3gfURD8osW8z4DJJwgdeOR2RhQ23wKo6Ii560As
TL7HHLV0APjlQk6lgJBu4EkxYTYaDsBmu9XymRjdbNjKCCZufDY+u+juk4dtsA1LX7UQehaQNfFG
6vgRRnItxUi3JDLsXvOGMpblGnmMXr79zmPqZ6yMrTA/Eom31ujnusJazM7RGYglm2jZ6djfYA29
QRyHmwgccEyCKhtlIisoAcaSv9sbWNJr7lwusWJAae3cjM1PvJrFD2jFhT1eM8B51fuZmklH3l3y
NyZNxVf1wS3osuUvEohC5q1P+0VHM1tLU0Sk/t5vBjf1toozu3p5o9mp8BX5MFZ8LjvV8QAjIb/t
uOcMUAbkhGibiJ049s+B9/f0Nr8/6rRJoXQPFQaWA4qS774coxIeO4jxQorg/Az7dR/rzYOn+saC
E3tmEvhqD7HrTB9Il2Gk2KIm1TCZiZnGq6+5eaPQ8mQdvVFk7XIt0ixvnB4ODEjKPAsAyQem09ga
6TI79fi5MfqjKbgBb7zpY7pJGUgunvkWKW7H7nhgAsmxT4mzavMmN2Z2n3/yjpnrBjAEPPfs+vA3
nPZb5Av40xtYKS9ENBF1oQnjxav8A3FBnA2NLsR81lC/NmU4EEYnaMt3kqkXxXtRCAW5ULkNjVR0
kO4ml6zETPqFj2SfoknnOmaMMufuOpAIYC29p4fy9g8+X2RRNf0fK/WTw71H/7FJTY7+7IjLzkkP
pIy2OrXESQyqVc6hrvsiYjOxUPdV3e0kfcCUpIgwHePSW1ogW2LLyPv0FgfHEC8NVNLSwip2YHsq
S/+iqfSFKRJYAJB7CXPjqINKRq7h8/ydE3Hdl5qOM+nTsNMqqIDF5Nw1GPDuNqTMbPLAM+33GyXQ
GAwqW5eTEsto1YORqFb5PZXDlgwVZpKVlLhfaxkQCK4ouNwjZzYgDVUw010QzkZsKio4ng5rdEF9
oDrXsln0HFJermWEVWHgBHk49oOY9T1gYlFT19kHfJqqH53gO8dWZR+FK8ouzt0r5oAPZqqcRzsu
weiArlLR2e8h20i4ce1gsHOrNp/q3suw2L6vtvzW0IGZunhA02JwAMnaaqy72pOK03gCRtbhK1LP
5pvp4Ova8jQ6DcjzFtc/JJx73/qx9xlw1qH1qmhhzBvNUXUx6rTDIPbLLjLVHG9/juwW60s5DLMn
EzScN1EM3J6Q60y4YikdBRDQqSteVElZfy1fBdzhv7Z/6R9ClrpMCUdGCnqPOzB1pwZ0P10VKB2l
eoACPlJD2XC6+fGNEmrZ1VcjFKNADRAaEG0vO49T62BBsBNFAtO5Y4/u39kK1Wu69fsvx01sW7mr
6MCEW6Pg2aI+C8KGvDF9YWJPYs9dc7MFKN40gtYJgj5GUCE7P91ly7xklhQeOM7ludnAlv1FUo2L
sq3XeWTCyfm2pzHTLKTWkGRDOV+cu1pUSNVeSaJ0zmibLkZeSGfoXAkwXVyEpY29zUgdamJvrEmb
jSdW6tIaJ+2RvshRGcemrfZpAL1Weov7+CWdQkMfdSJkgVLI2Dbq/GCoWzGGGi1mqo5IOL50omfv
7FrBQRCsFWIl5aju/8R8cfZ//EGqKvmPuprZO/xD/HyeZJ+MJBTo16M3lSxe8Bua+O/mTc7tvqNc
RhagBrZaDrx6LQYt99gfD2Mcyp72HH/RoB6F8C/ouCOtENy/iZFQm66tmHoey6XuNu5bzFHeSBM1
NGMQ1pTdZf4eZJATZd9NQhTmfbwb/z8KglEa5HwFF0SDcXmaJ4Z/pMP0kipUPhVYR2xg6ayh4bFA
jCHC4WvhIvFEvExAdCr9UkbeHezqaT9bWlko+7Laid8/iDkykST8xCJXxQprxunhq3PWlkE5rqPl
7GX4O1CYhgClZROx4CcKyOqVHQ3v2AyV3YyxXiQVedW/5Sjz7yaGXeJRGSVxOqE8bliwFT+VEEgm
4Cq7X4jGZDZeYhTuUKncurOKyFruAsqXxXzhm1w/9lGztRIfGFB8rU9ZBZ/bu6q0APtj3wM2ZCKK
cGK/6L4Mt+qR1UQjjcqdLpOkwg6m/acGfyCw7lvF5kkcSrlS+SIxJBsflWGTciogGnpVC1fNAdHr
4pcTUuNIzBkbP1SqjhPgj8XrYVuHZwsdRlRTMFV845evPtZWX9kNuplT4FcFy7RR9a8Xn7dtThAf
B103KCs/035m63my2J+BzRwjuEEhHh4McCwc9bHSa6HQj2ojV/NhUn9AEEue7DPCG96ETWoECsBR
DGFlteevG/bf1arhD8fXzF8t+OXzwZBGnEwyXxfRKicTy64HnM7FOqoy63jR2OWhCl27P35nGrns
oPHng8HcO1I7xWhuWClGLwnK7voSO9+cen7ZH0XKTMQKggGCGWMqhmhakF3sJbKrRLlzQjyRVHE4
xXM/rC7UycS9wHyZzfrBXt/ksCyiKf/nCD+pnKhTM42zFtDbhO9h06QzV5gWgS4+561xAPrFrBJV
adaFv4of5lwNA8TcgCcpIGKC9oNuN4MG403xDdjNiG5jiNSJeAxkiVzUPsJM8Kf5zurBmfjItRba
vFpujZVzw4FY/Px9Bk6HtvTAvOov8EBepqkb1RFghLW//6k1pyl+Qhxzv3zwx+fBskGUVaTg8SNi
KNAIDiFqaFFUF0LIRiZVAgm8jP9ROrCXeGnyfTaHx+S2v3V7Xgn5Yx4MH80q1pa0FTLp6uunB6Jb
p+n91BxVlAa1ETel15kZ/3TNtCfXAN7twVA7XO6k7Zw5PjRnqEopZ6vbgO/VO1lpMwwYJe51PfTF
Do3NkClJAgrTLcjD4usnOEZM2mxaIlT0S9zhTyqxx0b/H5P6IPOoiZuywbVBJDf8o84w2vI3/URW
81J1SU3hRu1IC7b3YNo+72eGvuBCHdW7tkbt6IQD6MLqfM/vWJkm6xcm+2pHV9XvfggY48Bfdhea
AbhtMXNBfbZo21gYxQ2h6Lm3dDC7iMdN3xEDgiMDrIJk+gjuEo3a0p85RnBTqE/LDsOC/PXwGoG0
tv6F421CVqK01r9uT/lWCTFOecFwT7vrsfgf+rG7f9OcRlt8+l46URmBzDs4zIomfu6f4IhKw/Mj
eY/C7wZ9VGZG5PAqcFyDatTAJqyzxRZvM+flR7oAq1yoINBNJuIcaqxghuJYs3tv7gZvrXxgUaF2
qyjBzR7cdZSDIiAS815U4Zogv6wIhk2rudVQe0GgOHh7oh7aE1AkwuRuSO1KrsEfV1yGOmznj+GP
/rENlV/0OUcCUip9YXwjHOFr/Z71fgSk7fSI0APWF0lJS4PxBkWgXl9WQAHQMPNDfEoy5Ygd7DZ2
of1slvejg3oiRxaRa7d6ugDcPbCtBppBLlbU7h0gv4puiQVbzOa3oF4DXvv6p9PTrda7DLgwJBR5
WfyMHr/nqSCS/Jt1OvDYvicY4B4O2H1jacBWkjjnExwg1LLjY17M5rfYsah616TQIGN5TEuHclKY
nue3YMlKvD7psIVNBMZ9keaKRbTpfhSXb3HlQrd5bp1JynFbX99fin0LhDuedYmzJWuKXOXE0shT
B43X4Pqksirue1Xt0Zt3Zw2aoqe7OUrycv/jMkNo0CE/Lq76dOzkD8JmrRR2BtPQPt7azCQ02VAO
P6c3AepBY778HFZKz7+UF8GtJpTAfWyjvsJuuzHfjGexpbbIgrRr+nolbLocggnt3VdWvb3ZO1M2
4D6P4aMj/MmnjTTDsTNpVsnWP0NjxcP/+cE0QlNJVUxIJr8dEAADYbFslokLc8V5DURW99QBSNex
gJ7YDPUQ9lng7eSCs21+9kRAqir7Wt/mLJdp/comJKXTDyBcZMioxCQO4DVB3z1mTYG0cpoqZa7O
t5P5PG+EiapGa64BYSgVsx8aUDeU0yo5QdHrHk54OTjus/LWVSqH8OG7IwFx+MSTY6cz/AxcIS+c
TrfZiQ4f19MV5rdl/pGB7C9BrQQQrASj1PnthVuDwwR7KR5pQOqxFF+0HAkyBQTb1RtroHUGkaRB
N6LWQq9vyGpSn/EbRpdz4nLVe1GVW8RoS2mhbE97ePkfrJF8rbQoJ+QiiVc1gsJf46sa/uHaRKj6
sfsW3dLRrkO17NVmj2yEh7cckqALCviTaqE5EG7rbr5i0xgo3ik63CG3grTPw9KVuH51xNYysJpV
rtzv6OEHuM3G/hd833njaDWbtjwgZhwU0nLvVP3UV/ziw5kAr256zQy4ua7khEV+n0dQjwM2ESop
ITgyt37tkTZ8wVIf989BQlPDHyDpnVbGkAcSACCoPpX/56zI9wCnPlv8SbBrBD5mtxdZrMLhZcCG
GfBD9ZUpLQ5wi8i3hGnafRhiNJeyICB9ipV5aqwyt3nqH54uPVGI2EqZtcqwZDhmzzXZoXajFCH8
zUcrbYKCI2DvxApzzM3Qm42y5QyCaUyi6fFff4tUVv2aOddq1E/Jk8aIPehIzr3vGbbNvA5Jj9EI
ZFtnOP0HDNajil1qNlGv+lcqb6SPqWyJfEE70Kat+FQTbDMt0VRyRjcMkZGjOHaQBCSKNCRX3jGj
l7p7QlGz63R7EAnTsFXnWoFQOwjY76mAwooTO07xrxLaI9GoLKmpg/iVjsQgnf9OmAR+3OK3G+U+
YJ63WuNnc09ikjqO3yb5vLCNDHqd/rYMMUClG5P3ujHslbpOTYuEPbvCTEnGo/xNsEiA491xYiOD
QKrrndnd7thD33MmnrFuCaFJNTOmhbwbQvWWZFfF51Dbaoapkrqi52akSbxKy3OYW8cy/ab8tjqY
qNDexM3KhwCDnVQ1+gPZxAhjQI3pyGomydeGrvy3RTfwutgC4jpXWtRj9+uPDhggcnLIYhOqD2t3
drmtJYurSNuo8dtwh9X5FtiPTl7XFR3sB4JQTYM1c15vycpq0S7XTL/04FMEvKEhqdaF8ZdFkkqg
vHerSJmME5o0SomFg1PMkS31ouBGxz6j/0ZI4MJeISgrhSnx4I4DwvpHKVme5IxoJbvBlBfHW02X
e263HhonL9FhS+NCQUkANdWYnw7RLwxOmXU8b82qpFBbACXJst6eP/GSoGkHdTLvsecI7bnhIqg5
TCZ2wAHjbg2aeLE9Th/i0W2Jyy41OVTPJPYtRmratmPH7LX4b1aY0XzCJmdJ9nO5T3+7Ju7SnAht
FLU+SKPtDLXdHEWrWfayD76nHBC2fNR2h12p5VtZOdOa2SGH+D9WDGCAEa9v/696DiOq2YvThiKP
xv6H77aH2QvO9vb8Bts/FjjRknUeuLdwHiQ4xz635dQR4K00Pvax9cCAA8aV+dITmB40qi8O7XC2
UIESKaskU0wYq001/BqT9YSvQRDtCOx7aJAugEg/ud4mmJfF2Real1r6tDNIrARsZuvOPBgj8PXV
aiGJQKsSRwcj5f4GiqyTip9fd94a568wJgWr9HMgtbjlJLr7DV1yUPNe9fqka1y/KEoUBpAOOAuZ
h8MUEzy0z8BFLzOLhISGLcG5PCd2J66vqF5E8OJ1F29uiUzVdUDHeiBs8/Q2lRW7FSKoChV6p6pp
6cvkMimoEjx36SNFplkmST9+O4tiuLqIzGLQGe7+wKH98QwEor/34Q1olg3UgjcDMg6CehxMg2f/
NwlpSdwjFiX/CKvFtIhrJnLy44w1/ODqyMyTyKHQEYjXAKxC7OZjOaZVEnFRn2SpjIfMOJQ4M96l
uWL9IUlguBjGEF3PSav9GuTHasUQlzQMIq/8qnzhhGlPGURJKMVWHqhN8fJJNiADNXwAA2Wu0Wf2
vfpF1m2iu3S4TamOA5g3tGYpz/9DXkSRaiZ0W39KT+/ZkE9hcvfUFJG8oAUS+KQSsd/QxAP9GfQF
Xn27+b3uAYsvVR1cQB6tg0zg59cBznZsIvJJ6Fq5zqV5gGtYu5JYYzbBN1Fn4Bw7PXKx5yDBpyNW
DckiNAYLGEZJ/unJ7Cfa4tEym4IhqldorFxdRlOUVP+EOj5JRdmQADYmLu8PJ2JCyBN0KTbd/m9x
xRNwlK7Tb97pXI24o1x6GIv4udkXqT4BoQNVieXwBU1z8HMHbh++CUjYVeIWFGoagxN1QKK6WXWY
A+6symglj523sUpH8y33E4YhSoUIFN1emI9Yw7RPiuLf/NVu952u6FaoOdjIAoBfToKWud4yGCO8
bVhWXkQFqu6iuYh/gKauhHSadslSKZxP8b4p19R0AZmQo2pnbIe/N2DC5dYfPU3dfWJ3SehGgatH
oI3si6WxK64zL8Ch0EU2hEPogL9+mzOOAZ5nHihNROg6YcGFhHtU2dNntsGMnYHdXbbwqNth5Wsc
RTdT+Z8xRqUkH+mPZLrdxt1gV74d7IWf1RS4E7fuISdoLi+R5fEnQBHwNv/o/iLhA7VVVSmU8JYk
1s3OnZfQQCzciIxadqlQk/tUhrToUBY8xZNsXhpTbqarzgkFctupEzVYEDCAyumZn9yfn+0AWtnt
3AilaXeGRvIJTd9NP4LFlXBYm/IKDUc8qnXFC+zjqLc9rTWi4enLfmFjKCoZxtTBjAtL/gFxFyW4
YZuAZ5YMRsssAIWvgd/mSQpuF6g/YvAgpvuLDjpnLbiaFRgC+/dN1+LEcq7oDRmS+aH5hld5Jf+/
k9vVOmAAKBLZBjC2ZwWKJh6Q/Po94CqoHvrMjNTWExJvejfT5mVv3YRQ+gE7ewm07sTjbZ+Xa4hg
hk3AMthCVlr5xIsvdJO6SK+RK1tE83Le9iwq+IMUvA9WXFwi8qpYzWUYY/b4cOxs7upufEStBr6s
WLIFS9iM1IxAqydW9uchhCGeRHP7ZgrQ8wE6Th6x8HAe80bx1vh7/v+wuL0dWhjNCXC1fkxlrQGh
5Y2jfL67j65ctdp4j38lzWv7Zz33f27vJ1l7rkxySwHElK6tYrvEBrVV/rhcmUVQ8rJxjHYK05i9
pb2u+Fw6BAHRdNScPaDYNeCQ0TxDNywmVZW+wtTkI5dw47z+L+kh/pl+rwd/D31OKR/v/eGf6CuE
cqHlJeDbkhV0R4ThK87pevBni5KwNCrEFgmsn5gSu7Ys7Z0NRGf9l0kfV0VJtSSGdwiQCQdAmHpG
kvNfrOYtMgCt5ehMCOV1MXetBo6mqlE9IgFBpBsXzilvUHISE+E/0E6xQhux+9eP0fGyiAzFZaGl
Qt+/PB52UYD9hYR29xksSJwqs3hfbEkU59aWZ0ficwsFwKMJ0ISKx7+Ym6SEHarer7rg3RbAPD56
DHvKhs8Aa0ok5fI9jR8Pn/T1sxV4gdAx8HUQHWzQ6gp/giYb/lIHKBIXeYwbJBpdUgn4sg98nYO8
PpZJnF5k2YN+3cLW8+63tVlyAT/h1gWMqLgs0BlpSHbY0tNLfjGaFHqnrxbgOY+MepFYWBJM3i9T
dBAReimIwajwXb/CKzbSSdm+tbgT1LHp4XJMVWuUm0cEMuppYPqtOxdlYlMmjZHkfN40mMsK+bG4
FDHj6HkB9Jk/NiJNasSOK84RCnmexeUvCfnA4JQz0a45cfSzGZ6n5+ZPKcZDHiyFH/uqgm+BCD2G
mliSidxdFxXN338/WAdpZSFmi1hf7vBkHtQqrh9R/L98X6gzNC4WhMWiKzlh3Zj405lg+7rX8Aof
QgzimRFUolT5aGay/O9ppegWUcZ0RdGY7QN0Rh+Qfw8MSzjtlkxtBlocY7lF/5+vpFiDHN9W6eI/
h2zUNb3jS/QptkpnQEpE7HILDfG0umz4pCNrQNPt9/Ekl3y8FyBfl3HWcOdV+CvVzox7RlSVnnaQ
dNy2msbMzki/yXVkT3OWotWlW9Xguxii4yjyvZl3sHdRo8qlO1sWJ7x4m5N9czP7qm/I4gOadFxW
O2mbXMmxkWMFuPg+Pnu8
`protect end_protected

