

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PFFltKdLY0A82yxFqahMaWdN+zxj5kThYAcsDyz3A2vhpKKQpGJvV8/AkpYYPyltKlIzJB6Md9uF
AN2ca05J0g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
obdm7XtHPDQGZMrK3kNZKnRt8ypfk4aZ9VtSDpnSwNdbgwrFg4uylDkc4YjBW8BFR32vEdXmCKFe
3L1bSMhXRkPXZ88hMJlBty0IcmSYNatn3RV9VG9yYtXM73zMkJ4NIx7KoDtvOCnGQpHNAJTknAv6
BNEUXajqHzh/vB/QNBQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nx2eU410BtrBCSzpvDl9pNpIplyp0nHGgzB9LvwnXgdhN5HNF/YNjnH8WXRfWZhIT380E9zFeNz1
cIYhUxogcuyFP2sgar0PDv645GG14wyLd7prd/d1E3Ur29iNukQkz59OjXTEIN/U9Gy3hPt+oLVA
TwpP0P8RgeQqCkJY93IlvPGfZ/yeDQHrxDZUMFMxHHI51HM/LG6Y5RjcVEJMkX5GTsC4gSd5fEHc
DWDREOSmqmG5Gmciy22xZEiB1SI044vcLqlJadcUhINRbAw0576LfZrf0pjCGq0s1+nEKeJm9MeA
baA5VHd6hhXLwLD9jRkKDvFp76mdZ8cpvFpcXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
my8iGpxybuJuMik3+8MRqWVv3aAmCE4oY3Ij0YIUQTpme5jJv8e5DOlNoLmgXWhUlepBCUyZ1Ysj
JGlFKQ8MBs9R5aa1TLi8cCVfI579Nm4AO6VpackDfb6c5/BXCbiBb8XeC9Q6z0hKyH6xYDDC0Z7w
m1jdROr8ONcmGBJr57g=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pEGUMbCVqav8XqUNf0y2o1L56804gb2pssAnfqbrEzVo5CXZ9MmyISfyPG7HY7huXkJ9tWIeWtYt
bUG1XTbOUAj3uDqhigkZ4KnTE/68izmD5rgLlGDQ1sI7w5GLUgtjCBINeZsiQZ8IbdNK2b2sCu2x
1k1tcyPPvRv3myvuFaOhmiYYyCNc8F9T3cW6mq34yHrMb8GcN1rGLFkL16mdIcoRSSN9znhYYcLe
21llq9uuuR5MD7mOGEYx4bKUQGVdPOHLC411Ms5bCd0IbhTC0qWispRkmO0D1uXT6TguY5Z6gKTw
vMvXdJYpwStmSqzikX3kYI1zljpfWHQ7HMzzTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 66352)
`protect data_block
1qTTaSbOXmFqMDJE07F2qoQaoRnrs0o8ZGK0BRAnBEUWNDpcnQe5gb2JywmfAuao6cHUMB5sH8nM
GKR44hLdu7Yg/bVS2p0Peavenhq5zRUpUcFgYkdW0cr7hX3j6c+lJ4h7kDtNFpQei7Neoi+q4flp
T07oYwK3GzN205B61zlYKrdzxLnLIzduS8f4+6KIie2poCmOo3hEpmvVTHhoj+prQ0ukeHaPu7Qq
JxTuPmHcCfnzWaXkybe9aFg32TY4wMAVv/qB8UQHyqwiJonW7YWiVh+/XNaKhWH7ds5Jqqz3pnr0
yFxTXz8Z1Ky+4mEfiA+HDe/DqVjiEm56n/KBIFH6pr5W6KRY6RnxhQVnWPYGzM2Y2izZ54p2Zqml
stHWknFQrUySWoqCHA/tq/JHTCjV658HnX8jrSIaIrYt1exV9RPsqufnjlIDR57a3sP9P4XDe89I
FP0O79woSMMYIoaW3j7n+7P/Vx9t345dJK2ymBZkY6nyZhmqbWO5RU9vq5wZ+9Ev1+b/59un9rZM
TSzlk5ModbczWpnwiR4Tzf6j0S2qAFDREWwF2gxeQyMquULDN3Je8yLPrtMCdMP6xkA1KnK28fMR
empEOOCU99Y7VqGlobtZQN8vTKr7DDutzVOxKWWnLMK9+z02PgKM/QRsjVw8Z37row42dZ3qtK0n
OUVuUV9NSEvwIgoA+UJNfmMRI0PqI9bg5XC8KFHvDRf2iTW3N8RbYpaSynqlMeMyIqhmpPjj5n7Q
K6AomFCWB9xQLX/qS+Eb79GqDCH2Pud7PdBygrVothdplqfzLwZzMHR6aqZUnQ2PaOb60BlbzSq+
UVSCjZehFk3QeQkTmCQTMi8Vf11LNVgH6YPyhnWfD282v9IoCPs0UD078a6ceugkwnCKrmuQIje7
/6xqFq4W86rGZyLIUck/Aqu2VXkJCInihFjrtEsh0+IGwM/rz1BaBhTUN9FPf77dv7OWUwtujOmu
4XBxLxn+KLs+2ToejjBfE4xnz8Y6ReAdCtKJNxmFAGj0/u+TAF7jBjsmtglZsm3igMrTMmuiCcOV
jen5X1jNFshL3IyegsNvtmihZ8AogxMu+L02nqF25T3SBZ+E38hqeJgC0vrPTEWVhQD0WS2a7cRv
ruUf0SKWBNoQkXgnAGCyjUn+AsZaCm3lvzjGNcXDuBUQO4OPZDXCDWo4RssJ+S6ku1Fm09B4wpK/
cP2ojuWOYx9qYpZN3hTV/jpEG6xRvlKe/hVDde7pSYMpiUzFZEM+SMZpqmdRTCfBXo8Bo5fxERZJ
S97FuSvrm+oJ4rS6F0FsKGrGshO4f6qBIciKSQAKugZHYOJ3p/om4yD9xEkciUKcXjHFfx/Enr/w
mhqJ4oRHiohhctlGWItULV4mN4/f3EtKWS9tBQ3o/7KRJ3pezD+8hyHbPtuSZhkFG4Yl7PuMsao6
a3jeuJT4AcrD02Koc3BAjj7rdi/MZEiBUmFNGha+o/j2jcs15wsa07hu1WdtCYtwtm4UH7qGogUU
+VBAIonX4qS8B5yfBSrtxbU2ZQWi3mpiIjQNWSIAj2Vw7X9YtxqvyZv0v1jBpuBIFcs8XARQfvhj
XBmEKStr80o/CDvyuCzxiTUrv+aG0ln+hC9lUpegXJN/yhSnmLSBWtzOxO8DFmtGZl6QItB36Ao2
Kq+O4Ca2pWMrqOgYNvjjv45CfMWruvWWo5hBaAszG1zsJFgtGt9ZhU9djqSW6NArIrj6Irm3fWox
SnMudtQRO1v1kKRg8QTOGjbJCX3ehRisfPrNw6vPq/yjAhTVnJ7q4Wx1XA6cb/37cbSO7TIUOw8g
BFqvezCVU+0ye92vMuHIRTtLwU2tHirH29p5+Nbf4RjiVEBadG1Plb7aA5d+OWMnRb+rY1p7Z42g
XbujzOIKycm08KE1/mJzWdDjYRX2/HVFcJ1OxFpgUGLMyiXtR5Tbye4JHtXIN89FqAS6rN77jJSy
cCASushGR4UMWgIWNy/0fPkBSI8ZchQj2lR3+ZpnX5O5/+du3neVhnreEAgW1hE283KFVufc0EZQ
VK/HGTIbSSB65MkMylkoOGDQ904LSPybLUGrNmcjmf7aEmr2QjCtKXd1rByc12hqLMT8gcTDv74r
LMg9Vda5SVl7h7uhbmfmZAA+Wlx1PQrt487IolF1R28h8mX95PfaHaF96XrKT1A0SZ0QRP3znPbN
r3C2TMnsfBtUXqDn5FERvkr02HCFiaey7EB1p2XFeTs4yy20BQS4YJxLOLxhkOb6w371B6S7E0RS
tqkyqdAC5boMR77gs+EuBCPx5EkYP7LrlP6qH4IK183KA+XVmRUQbbjvVSStFsvmxw2L3v+6ikxb
4FGz1umKGtde7G/4OHAU3bzZ4vogqQgUdsfnQFQVvAiR9SHV9vKOsiVT+fpiLIAIHXdoagevHB2R
/GWvF0hhiACQ4yeZTzd79PFD+o/+mvFi4TgxJk9LyNu510WIEcvbfU1hUXkgyWiB4QNePdFNMpQ7
KytnjZppcLf0Nmtzt75OBxbe+3T7dlaiLZ/NKhWJUZOqdAS5UoGoeObWSkQANXdYsndBN6yMQqRE
JMJ7IqGrIjPxGhv4VY4KPWrl3t5UTsEQsoQEfbfh9/Lw2Nc1oZA9vYqMyXF4xmjSIDx3eO6wNNrE
0GTDNkb3SBW2lxdHRdcCtlbF6/S1JMdMIDLsQu8FxMKFy3kPJjOqbPo8thUOgmv7RIqOx2EBf5da
0wuYaCoaeSCY0T86h9k6L/mLiOx3LHno7LLVv1RtOKQfs4eMrZlUSw7CqdVnUthgOz//fFdQdyi7
Dv+q3qZ0pcccEoC4yo2cKqmEc1hpo+eMwJkUBq/+IUVxpt8chiJOcffQSbnmVidzfIZBxPxR1pTk
bSLHy1FPM8dM0V15T9hb/E6dpuJt/OAgR/aiZslYRBHOm5IjqZnXg8gRsOrI/TEoCeBnOuQ/0V9o
AiPdzAAGDaDgBwMaDvhjeoU5Vj99yafI+VQ7TWHe52hbryNU6iUZZwiQY7vlxqLfI9MkZlOeZJcj
IBI7iJiFRiE1AemSUWpKBkqyQqxghJsiZSL05ZquwK535wi2+HwKmTti2dsetFxWC0stS5C0Y9CE
n5W3DuQVtvssD6txmuIUG17EGr5hicj8KvbFe1wOjBhHWn+WHeDcU4NfDtscx6m29j3OX7Qcyt5r
JCsc7eqWw9+YVND/95CCK40hXwm+7lx3osN5h3SGWcMzM0KhYc8LZdwXx+40qb+mDMqSg3rLZ2Uy
xfwjDn0NggZEDhlrmfb5ICw4MceYaQ1A7HdvR4jCz/PUbbghIT92bOAn/+Ot0WRq7ICCEGVEOAYy
0KSUR1MqHBiJwR/2ZrRidAz3Af5Ikn4s9xxKp32EEt2pnbX56BA5+kFj0FTvSPTHautFUWXyLXN2
nk8AqiejyOW/3JNvWvEFLCeWLFG+oO3bVPNqWDBKdtkYsslmM366xPtmqJoqTqpkQPmNhgjXuADh
zpwTbv7yB01hRlHkW96n2GkJZvdpDVFNuqn7mkEuPPgThFNc6bR6np1Gj1QoahtWu7c8Xmcm2GPd
qya9ScfWsjscoA0ctBr/IincCZPwAkJiSFyiHd2bb0sTIGJS8wezMMBHCvr+6Z0azHaN1UF6yi5S
8X8HbJX2WrufwTzkibDlM9b+i31PC4ElGzjH9/uoOV512HKNc40QN7ZZ97zbJq/rs2jWsfEZkjsT
wagIBWbOmy3pc70rvru4r33l0a+t63o6Jc5IXNTNqJnPaYih0Pc8y9Ntgj8UuLP+aRJWu43HOvkY
Qq7XPZOMq3oktCTf4D00IxdaOkU591ZBNqOZRBjRIOw4zttaT2oACGMW1YXMbgswNG6J/ZFTuRUX
iZl/KEF9X1ZTD54daeZ/j0mwAzqBO+H2gTQIExNbONkb49+D6aTBD49Clt0Duxlrqpj6IfPbArPG
0es1VmZKrQ08slVzzOSpKwHGDAlTKPy26UUgIBj6LdmKkB7KB3LC4JNAkCplHC2w/3Ptk+vNpo/G
i2eg7dzyBxFiNLFmVKx5+O0HYc9rIxelHs6LuByu6rzo/Pq9lBI5CXLGXiGm1O4RAgqLNcOAJp3p
xh6hZqiKastyfKRsiWqO3ACJecv8fIIpZ+ixVoqfL7sJ7X2GW/DD0c9i7S09pwoVZhmGl6w2PALo
t+7QIJ1o68BRrHm60FQPjMRH7tm7XeRnAw18IoRhKUznhHcY0uHdt7Xa0EWdezQbm1g2m642BFan
dPnvW0QowpSSf3As+vxpUHDJFXic4a9mEDgSNGWLRaujO/W+WzOG56ufJzeMLYCbpljwPm+AcDe3
dHEYeQu+f58BLESFKJgcNWW+JeYs7vdCMK9OVEkIDu/Tln13mj2X7H4rSx93/EQoyKTfFYxzo2Dg
j0oFBSWqtnK6tvv+sEC6DXyM/JymisVy0fvKNOZoNEsxH02mcfG1JW9Yyv9d0MplhobiwOomUPfD
Ys6EKlc5/nzPdsHWorvsq5uhqgj5w+fpp13QcVbfOVqbXqd2Gtj0Shfwk1Qrjv1SlQBiohLSHYNz
BXASTXM4gcDFPlsHvkntj/od3EBx/VABG0N1U0MJUOYkBzRxXFwSsp1bLmDtShi9hYU5b3c00i9o
pSzRQBaq/ZQ4qeLW+9RKk0ClbzTxGz59iGa+GaMgr9xOSucJgFRowdVn31P/ZK+Y3TeW79gimK1Q
PFuCqMXFV3hPVzKuMYUmfx0UxmAH1bTEUQfQ3TX4gPMnqJcg3/c3MiLTXtKg5Syg5DT4mMeY/8xs
SP4AtU3hg2msQBch+CutjAM55ZtoNaWhs0nEI3OQW+0ICxAuTV7bsP7ReD2H4Rbe7nmojkzdBH11
iR4gogLo6G/kSdaKroAGykWd904BXSiGuAXwg7jRNiHGtm5ZBzmzTc3ELF7/03Xpv0RgQ5nNDc+I
Pfm64pdogzzOIHaM3AuwpYjWfR1luAkdQ1q5RxlXz0wD5dPUuMnHfaV+VI9EhF1leo669ewCbglG
wZ7vSr8JC1nS5J3LTBzx2FzOz7VBHCIVYj4Ot+GJ3ZR88hZQHX6358jfESFVQw/CXCQbv1SfUGXY
vSu46sVVbwAq2aCY/WSEfiQesyZr5u6vK+xZSiH1BySPeas3Nekhg+aBCj/4IOcI508I/KS9rPkA
u0imsjiPb06pBKutiox+95MuDRjVUCtHlZtLn6QseUda3WK3KaT86dIuLz+PcB/vGsqZmGlYHRSZ
JnQPyFe0qidn6ZU34PqlxcGF+0zMwCFT6+rUeuaGbUekHiw41voRNU1+Kmtpvb4s/s5NDA7rsH1O
OSR5nQvKoA4S6neAguUZ4PrJwv9/YouBVHNReHUm71jYRnUJSeGyr3l59RlZ9oiNsfy40XJKoB7T
0krffNyCdtMILO5kdUvYdYqXauJtUPYFALFyiiWy1iEmRoR6FF4w9jNYa/5RCzEBUsAfKbSA6DtF
TZUEMcBkPrnMo4KLGFWHXusQLnWVuzKoD1BiL6kz7NZXm9ul+sN6MFRK4wdSIfsXrjLQYYlFd2fg
P4Hfy7Y0g5DFw3bg238CdoG4S/vHZrWV4i0yBFKbrFWbXyHhJZRSUSu1VIfUsdbHsK625GnSHfAg
g2mN5Pjruq7EAoI3NR82Z1BOOO2SyRx3PghDKJv6uhM5bH3ELaAUybiVqcZyL4uRLDlrblQu5qZ6
5J3VBAawR79U+HTZazC1WrHazSM6QpMwE18Oyj40SCeBLwZecqdUUqQDs8hwi7Mcrltj5JEUiM+z
V9h4BvnefRtWbEU08+TNvZujCXJhqb0OkeRaoxTNffArEas73zP8QxMIaSUXMRG5Zc7yof+L2ors
AnW1pg5egUSC4zX8pav+egvp63wemqv4PtbDs4PR49V5m6QRx3KRJ8bSdYfa5b2A+bT99/O+v7yU
a253woUcaCIhwnJ/PDa64KK+zL0RqO3p7YqOZViN0LPcqX/SfXfmrGDEtgqTVbxU1OwlrBPizvZ4
/4nVNVhC4w7ynAmh/RvjLIPsICaEzD1QKfZgoFQIts05wvqbYOc9G0jmGuM7U911akgh7BndhVjx
NFW7qQlwXtg2zbDQgsJgRYc+HiNQ3nNc3cHnLa98ZsA0j2OwEnPnsBzgsY10NVCMgoMexl663/lO
DGIaseoAzAbAmTSkjooUOkqtjDOOFXp3uSmR2ldB8gAvxabGjDpqIEJP9Kk0dbXODqQVFvdWzpiy
DyMOSJDHKomHUWtGak1m2L2uQmDhpW0Mh55TntgTzhvMI0PVoF5WyJXKA4K+J/DAbkc0z8u7/0qg
PMXW4B471CpXnnMVGp/+ke2ka7iWgnFFziEwh//+wkgfJDCjzgBVKZViiaFfyQYWoSh1qzmDinNp
cJo7XWBykIbmcx3prtkbE/UmPkUG+IH6QFB60tPicZElgCIGdRtJoWowyd1SgN3VCVuHNm0lwFkr
hnYVBdDoPrn1je6pH70TJGINN5eIRQrMYEIRN5GYV0N0sn5SrPuMFuVjRVYXjYNbOtFfbLSKIgRK
uebtgJodqrQv/pQ+/tNP5EBAA/9ZLM+YZONOcqFG9rDmG8ygSoGSGMts98yZ/s8tvQcgI6iZkJ5M
4O++j631l5eGMmknr7gUiZ7onU5tXCxM0ady8qst8wZYT4e7EyQ4+5yoekkOKwdWuQriG2lV+cDN
FvjehB56+xPgesBpcGchUcABoBvTHc9TjHdSQCnaEd84gvWsAc51W+G0x+SiDbl46n2Y7QlqAKRl
xSj/3kLx9UGizeACYcD7JXZdSeQWH22eVIWvbCdb7lZVoRUHsSqFQ8yB6elxTT5HEsg93pmTHFZw
cZ0RFFD7CVJG3ULffaWa58JseeUawOYKBKMovTSrg3JEj6Pi7Xel4KcQxGKOuaAcXK1qLwqSVNJB
QCkT3j5fE+XaWBZT46QIt4fuExPf46TgdchSTxZ9Z3ZUEUI6W9oQirEhOVXMH1rh1e7FLDHc+tpv
rENRO++Slvtc7AJF8xqVFwRoX4ThZwEtZoOwYqVqQzqBahwz9dsvp/qhdXNMDUn/vB3AViLvtvAU
FqT5Ak1GOyVWWIU6v7M7+qDaBfKx5vHgrW+02zwjCpbhKzbZ5KQXWK6kn6/yMciDR/uQIdUvQLxb
lQPIyrK1SkzBpr1WAYNeUmlN7AgXjc9zQVZHZM+3lohiVc3u3IYGZznEqBLDghTSZgw52OehMNea
roMKCJemAMkPD8TSGOkCfmS5S9EAxrttMHTvNq+vTfRqwRgoNEhpQN/pyDtzwboR1s5/BEhzxaKS
jKhr5USa39emVkObLS5KMxMsJBw7cY2E035X/T+xnKITAryJ4cU7+2knHPI2xaBSB6Vdo92LJdNL
CHYFEzMdYq1Xt6iWdDzEqTfL8z7HEUlgUT0PVcPaWe25LQBSqY22Nrs6NVnEzvwpa6VXpoCHmobP
FqT744gaYBYaa8SPEY7pVuZROQZmLXr6+5Jt62TvzrTTcM1jR4/Pqvi7Oq5/h49Vv0E6CNdiniRn
CT/oSIxK0uX9ZsYJ++GKu0yq7SV8c1czfTd/A9qDDUCN5JkjNJlue6cqz2L3/Z2qhaeaOqODRspq
X2qj7NfvuoFkzwUEnpr9PG2oVjWkV+y6i1yZn9Uxavh56/A4r0MvE8oM+JOGE83wsLzyJrgFudo+
M+BRcTKdsdCfEnGfkgV6cK+v82tS3owI5QoVIlB35xPRd+HfJkBTm8K+Iw3XX2pap8o1aXtDyMov
TjS3GFbHAtdUaBlFyGHhc2RxTPW8HFw5WM/Wj3diyZ5uYFHEeuVdVkA8i5XNaDoRAp7Uo07xT0O8
jCcmlnON8D5D9JGU/ZIpUCTdOiE9EvOdhebFSCJ66GDUNAfOfMANweN2jw0e0CmqaE8L4VLCmuaU
UshwXgJz+EMJUlwi0tfqGKQBVoUOORTqXwV63cgUiYcgdG9mi4mUBh2VHgcjDpxsFqaR0cY12dJz
O83DnMYCb4RjFOqSuO5c/0AvOszEJL2FvGOREqhz8p7FpOR1gmngX/Y3hjDghGrQgZpWNrL62DRJ
vhix1+WkivkNmQlaMFZoJ3mw2hpXnvbbbHSlQfarnyUAkxJpOV3xHRjbDV4hi1DjwEOkyOHvbKVd
LFIikPgEJFih+OIGcJF7r21FVHZmRI29xrHSoep0kXNYr38+vaQgETIAc+WyaIO3UH29QzzZ5sZG
OlbVjWe0SeAu/87XkrWZq/RH/CSBPupBaOQmddx1CwZsZDy8D9qzRJsnn8NOpNeP9AOL1X+wI05N
oTU638aIsNWp/f6bLsTmmPSBPoU2hfiPIbAkVSE9hfkXr16bK5FfN7kBOoWSw8+hDrEFWsZCiDWZ
RTY+eW6a8CDYVQRNlZLj1sOScR43WQvmZm4yrEqEMT9/MbmPzWDfr+ZFy72VRhl5oJNmxyo3dN8d
3NSu1NwMlHv5RbDhXfVjhL3/IKHKV3PEt5Jxditnxz8aVdCjlL2WsBGBuT0Xsd0UCfocHzneYcNc
3a1QD42cePGZQ/TrzUBQJmDP7CzBo366UdjoPGNz7PuLSTLdoDRWdQg8u8YyUMdVA2/6R8PpvoG7
UltGzLAjUwRtbu+FN5AR+R3FSAOP8wjwU/vkCzxAuMeMKJgcakFkqD/H7JzL1w3yNOyQFX9QrgfM
xT+Grhd104linJaXeCpQHcH/mMLw1l3ZUc3rXXouBY0WXhAI60iCcW4PUP6JDKcPZ2NV7/5RcB88
hYDUcSynX17vwp5DjWnBrV+EtFVEn5CFlhdP+vmK4ZghNkqh3b9KQb4+be0tJMv3q8KkcLwucQpv
X5TwpjE4wXbB0ShKWL68cwdLAgoLIZ8rTTfKXlbrk8aGxjm0WauYgDkh1sZi17X2hDl47HixNHlO
AADYEFjsKskGGkHWPjlVtgk5vRjfMHJMsIgc+QgsWYAK1PytQWWtigQO9hpMkYVadH2v1NLtgn4j
JFogxjeuLMtc/laAeKM2hzpo8eeJ0g6+Pjmm0LJ4gGYlHeVQlSayw58QLKZcxM+kapjlukcYXgJX
s2wSCVrZUl8BkvRwUHie270i0wZyxnpWL8UdIxZunMIkkFe/3+OV2/M3/KT7OYNjHB4toAEkeSsd
eCZDwD41uB7Bg/SO++zm07UpkOibrupmhHUSmM+j//y5WWosSVi0YjNoOpq+6DB44VwFjFPRI1OR
I3Dr8qr0LrwB22UJzAZxavdBubjkL6MGSWTdMvtpiTmzqQi4q4ZM8TeV84fV5DwX6xPGQsnwxMGu
RP+ZAw7hgtjapXbmyUOB8rm7f7aN84lV5X3EU49tOAuhBe8flBXNQqqOj1TJjOz/YDg9u9D48EWl
C7qjMjAOiDNb+Xo6u376uM0rLDsJNxV6sule+NZjd80RlkRf6vTo9RWM391PUNqU/NM3MnOlhAhF
2Zg79Y3wYiYF7fMoisjMuxb3EQpDyY3VZfEVUGp4SNwqsendgL5UEk2Sxe5rJyFQogUJQjNm0iRw
9JT+5M1HIn3VUX/Ag1jd97v0kaNcKJmfUfe55Y+ij4zNwVv9HHVbDtQLibmCt9cjwJekbmEV12dN
FZ/MuNpLHf5eEFeOX/PH3pEKKy+1yVtk6VGgbedxcenZDsAxgjWYs83q+0rDRuARBRROEbkesqKp
EQ3UTZvn2TehF5y7UfRQY9MuKOT2Jn/c0uFtGc0ZTELVc8zKGsHP3Yt2g/B9hNjFg0Nyqr4GnZDz
AbylwtSBHhM1Ynsrr/7GuEp/vNpFJqdyx2EhTGHaBFEg+yLZPFNnAg2DoeZEMfJllujXNhGSQlTm
nNc86pHyBFwhBC6LM73AfjUGOPskcQszEwq/Xky0C6QInOiw7sqJLGZy/U8AyCd15Etcejuaev4v
DtfQHsz/mqqNVxDjxyj7d7opWpyoKlLHNCgyvM+1ftD1P2s0wJPeNvxOlLUx46cvCd0A8vEpFV0J
SNJaVrmY3wIBqGZnjLu3AKcI9nN+24lYTAjFXQfTo2ub8DmtQU+eQcXJ6xoJ+R/qIsvJnrVik1LR
Ovp/QuwbMX7WD4I3WZMKyJCuf5cjDBmm9+qt70AFEx7iRwDU70kXemcSkC4sZhjn4f4iaaALVT65
cm1r6aiTtJQxKUpBLMcAXcvlcuOostCSjha6Xa+cWLTTRrgvskCM5Rabk6gqE1t/L0/Sh4ZbL1AK
DMKl1JApsWCh0biJ6Z7XPRPw7RmVUgeizbgD9koWnWjRWGvfOQIh+P4xtJbljPEhTnc2LmPe5QXC
OIg4xzUYVqs0WgAATacjFIvGxokhks++FhfzhfAB5X/KlUsiB/znadKSC5YWNxYR627+YvzlGg+y
y4d02AnT4Sqq5NgWN09ZSeoFbK6VGLUCMVacHzwMxRewTCH3lhVnTH/SOjLq06+XHHFORexqgJQ0
9N+5JKSPcYLLY4UaSkdNUdbYCefTCOx14URM9J2IS2cQWCfYOM59tgvYatpTh1gnNfDiHQ4sE/1b
obf0kLMHBroBT1mPdnzEhOcp38XYbphn1gV41AQE8f7clAvEpWs5oRJROpEU+vBybgM6aRqPrlkJ
GFMA30IFumO//VS/7sfd8qitlbBOUrOSLd1imXGCi4AtKZ67EAiNXfc1uofoT6EVCbOa6WNNFdKO
kSYXSnaD8BNvaN/FFtYp3gb4uZfV3udXBocBVipXDAWuDTY2GRt48OfzrS5fpRKo3SVOT+zx3e+O
90h13rFOMidEjyj/n/lvxn/wIrsxZTj3hf2ftAR9qod9V3+SxrCPGhLKIxwfYD4BHuVdVcOGuk6H
TmHl0/te4+DV4fMysNg+XsRgokgcR58T6BM+pTh/fL8bPlpvWCtN5JYJE8pLxgrsIL3FCmHR64xl
jWdk5C7ePbqb+gODadcfbYHns9KyP/uj5CE1V0yL6ROm7aKmayK4NGClXBwX8msshEFRVgvtgHiE
PSnZeroXKfs41O8Gkq/1obEEtpFGBEwlv9a9io1d5nxzZzGyzjFh11VH2wu9Q12S202JipVImQfB
WUqi7OB3bLxgYX2iaHn92/ibHlt6NER7LrgbY53ijWeh+S2UcoUQcRW+1t/834p14dhL9IMQkm2/
ozGkTLWedJBLVuyPm0U2sErmIt8O/ip3QOQDlaqikGwfCMmywpmtdVBnDMLl8VCZDh8/XHpJyQFW
atpIxobAwHgv7L1rGEAcSTJ9v95HsQQGQYCRGhKoA4vd8izHZTafd7d/XSdj60z7zpprZeiqe6/n
BFA3QiFInDSJM+J0qDzgviZU8kXoPM956xRwtD4yahfxGGoM3O9hxQqRQkq1E7q2BaNJLhM1O4pe
urRrJqKxTBNCkW5LHJNDyPEtPhgr3+kCM8kfgGp+pz57l0Wz+pwMKkrKp75RF96sp6GZacCI9Ceg
Lycb55jfJq1j/aso4cWpbudAbm4SrRIDYLl0mCSeSgRbrz57/VlNPETfwHMi/2nGq373OcUsjSz+
skaYgGxTszPnz3D3h70gqpHyWEpFeSb8e36s0iQOyA4dgG9A0nwaw9iM9KOqQ6z63fP1hRuK3wfC
y4q9pPJ+Spx1e1fevDldyRucoXEEs2iMjtXtM6ADW8RIX6EJ229fIBAFqIkXKSqo0OCiDo60JN9/
H1XszfdhE3ml9BwF02L+2tYkLnYcBFy6bmHyksFeB460vNyMVgM0id9FhtBSLazz+QuhTEjhF5Mj
aAqMurRZQoUBxgBR+r+4wqfZmCXUK0vXLxFzdj3Lvsi8a7hnCWP9EYeMGrJQUtf+tJxhjh7OGFyW
/8YXcpA0lx0MKQE9aj+lRoi5aTwxo8Gr5eq+v3ae3vLW8Y98z6hb2UCPSMeZ+nbSBEloEX7GT29G
r8j8I98TriFx1RiMNKQz0697gspISrrXIuPRunEyMSPkkm6b3qfXCRz7Fref9C4HRG1qMkoJF9Y1
MQGZvD3xnlbj8kur2qmzLDD/zM10k2pduVoE9D8k4jiPtFxk3hVgsba6MZ51DxD7qbU58TG8Wsa3
7zClFS5fYvOY8MsBkcGJ0Am5bvMKJnMWLMKS3xbheZUPlT/roFj+erQfrbmcVK4oA0O2JTXot6OK
XGe5zxAdc04rKLY1CJE4tgxK3cE+HbU6ZPpwVTEeftMpMmXz/hpk8+FgeWdUdyPP+Jz7G3qgb764
gVDdw2a/yu6e/9qfsHYzLdGWFpVQBJNLW97zWVqGQXwN6xNawoI2Rvxd5UIAct5w86OwRcPKXJZK
N0Zi/JQXoD+5TVE7NmzL1pg5KpHNYu6GYE2SrNMoQ+TK0QXBadwWq+t4XAbyB2caa+wosLf6lX9K
ChFa2y0wJP+3+L77KxWpuYhr6h27bZC53vhzNZkVsEzInC/F7ccpN5t9Hh0fPazxCd3fHzS7KZ99
wvzaGa1O2vs1IWQ9RFd33nRBdaHNEHHeXmpFeH9cz+4mE586ipNeschMLA/opdz6C6ug+cgFvWPa
BCm1ZiVwLXUc5AyDOTDe5rcr/sp/pcInKD/iNledj49fyIF7CeDHgTicTBzOrfHNQWm9PNAmvIZ+
Js5AZaGwYqSDkjByu8RyTBTbikRQops8/tIoVmVo1v1mGVuDHxsv3IZepjp+cvo9qErio4tjY5tc
igaoAkPrjTA5zAymxmFIRszqH61x8zcXQBRE8TjmkdiCe2AxKeoRV4V/A93ayq5sIWnAyDdTPOC4
HPIKTa7cdaJch3txn7UCdppoxfGwUlWNrIlBTrQB8VMG+kRYm6IvNU25gOyZ1KuLuNXkfXfwg6zD
v0ArXDxgmQ2VoQoUHxXJcjNqlz1ZZBkwRtZ8xNWqdwa4FUuuaghi4wJUCUv1M5QiftlIV6J/piJ3
uFLZ/dBOhbn3cZfPDaHXGLzi7GmETG5uCmfmM3i0DbdcemYPZ0Y71lCZyoMHitTAyuqDt/oX/hV7
42s7g+GNLZ25Ar8IRjh/13dcaaSC2PFWyDNpzsbILYuxVgZ8m4QliInovPAYT46AbS1R337x0F8F
VS74J+KNaOoi85OlgJR6cuRhDf0Ssid2FBo7StlPjPlrAQwnlKner9xy9u5N0OY3sgl33ler0ZDp
Fq2mcqpX4Ad5GLUXRW5vtByK195nJUuut1z92LwXrKDV1EYauY7Hjg+DdnaeCvVdLUvjH0/70exl
6LE+1KaLmQPJX5HgiX0aCKTxAO/cMOcKhxnF2EbPM6OYZCBWUW2XrOIrr2Wh6fSJRmB4bXjT+eAt
bkhq6QG+1sDhdvf2vs/nhmEdpOdO52GlAXgQcueQry5zNdMp0mS8krG5WjLlZkJU7guoKH2SLZJ8
W+QZSwMLMZTVNPj0HuhxlL7jh61F9T5E4wDYcv0vcjo9s0FqfLYDyVEhJh/pB0fOOElqo3YQJGph
akqYgixDNydEL2D1MCgbvLIy2hPUJD8OYrZcq38K80CqkNknJfqzK2u0stORl+gm4VgomdtuaJgo
SpdoZhcNyClK5tt4dlUirFcncOF+astf/gl6ki/57KB5x2dQG5Kv1SLo9vXm/3VV/MNVgWO0jq04
9V7CXzt7eca3Ja8JY8wkolPYdE0IU87aYpJ9nm/YXFQ7FHEU3NxCkmnPhrJitqX+er5+mvUyYNUi
2EkEDnB2/uFyawg6OYrBNxllpuDZv0oZWHTuam7BiXMsLK/D/3Fqi7oVWdB1//IGSoYIdcfiEtqM
KlvQZ5jL08us4KFv9YtX4orsF6L+krjuUSo6GZJMY2tdJI4PXRj4sU9O8OxWT1o7O2zN4UQY0vb/
tszP2KkRjSMYpHhvgSD39wLmMHgv3L9IDnG0VbUtLmMcD4lc3K2mh67Cn7SVDXGAcrG7m0QeeCKy
DZ6bsOi2F8Pz6ZWaE3TMyKAIAf9y8hOBktiz41JfttE8Z4JpL3t2Sh5u19++bOEuReVTNC/me6zx
wM3/mV3bUcloxSz86XiuRSXrgwzCo10dTRTLamfgxiOisAjChF9j6iu0hGeON311UN+BbKx1Fy4L
w6T5uUxH+SBRczeIBz9BQCajLWWReG7Y1TaT6v6X1av4iaA1XVyRNfRrL2A/nc5oeQAFM4zLc7/W
i3ZPQMffTmgHta36lnaELqMlUgrOFnxHbLt5cuFww1ztCLczaSCX9654fe0VMNvan5CkWCechIXU
JMZ1JVInIe7gaqITSXyZxHYXGyjtT7ZrR2fFvjSuk1RoSHZfNL+WJuxkN1xMLfI00etB56e1IoIe
RXUYt0uJrU7Em/dHduVQnxSmvdPUh0fOC1t62J6o3aDS5pyT1EbW2sAfK4AV1rPrXIvbIPccu6Pz
wnE+89nGh3FJtU7xEjQ4OHLegSKV7ct6GMq4ujS9lOnlAnnvGFvHsN40QcqcbTAe8uaT+QTB3Rbr
+B9meoiEqS3vdDR16ANCLENNaNJZ1Qu6SXlg8rfIqJR4wuqdE6gNzZFWY/yOLl2TwXmrcNUFU4hv
RcPnJIMfz+WARJ6hzy50dUfPJ4DCG44P4H0UslMsKBNGxxnnkCa3DOKsJ24060sg74JTo4Ih1P78
5MfrgVZrtD17vLRjLNOV6ZIUtWngvay7oqILPKi+Fivi1yswaD8pH3IK4IB29XDK/ptU8XaLSY6p
cyLUxx1Y12xM3Oiqa/r8yLgk1wT7FNF1o9KmApeSSJE5D/SfmkRDNA1FZUF3oAPb1zJWLnogVX2P
2pb3o1Azy8hGgKS0xTULrnUeoJ0l3zwwioUmg1IY8sPWHUTxrBzzXCD3K07KHWFrXDBOsq3XHGZY
HcMLfC9LJzOAeDl8zx6p6w83HbsoH2z2W6+5J8k9c9rwjxR43RCHsOUXWrMza8juAEjp+5s2DCbG
eGfSfmVTWlceCfhDgSBy56f24BPxR6+RsQoI2PzwdmsKQdBS42/PirNjMGlDewagxMqT6PLazvz5
pfr8WlHLGRzZISyjDD7ovpijlawGKB/54FE9KR3XT6hdSdq5nmqBaaJircgFe9tWTbaHQvghAKlr
TIvHtkk4nZlBqx4YHOQslW3UjvAqCQx/Ypeo1UO8Kvr+zVbxl1ohSphE5jxhPSY4xjfnQb9DDhQo
s/u+4BlW2TNE5o5/blk7dzRKF0BAdBMK08hwMzuLPu5whg8SOhQZMGTlABIqxtzzhhpVK8P8Shva
9m6RX/0TSOLMMSlsJRrKMgzSwuUxV+fd1ws58LixztXFcjou/RCGEiMUyUpoXXRzMfVfK5ln49JK
4RHXLEeVj0tIX0b+9zOADbrqBVUKu3qPjXTPqV/j9r9HpnpEj+9HSdpTTqN0R5lUmAtrRwhxfTzu
Z7YsKUEMUCzUkP2mRaKHYiliN2oaFoTXhdSn0nCwDMV9C30YVxfgO2DqKEM2qN2d1CezQegRIKHJ
5ZvDHlhHPxOWg3CtRGmho8hNEp+HNx1zp82fXtfqQzCfDL0reYR4wnNiyEX4icLL3Ddz1KQZAHUX
dSXHNTRW9v+H4kLUdX9VKupBjrOQrawVG2wsUBqNYdDogpJWfIE43uKQX6nwsNRdTIMMhKKcQNbb
K+9MMLJH/+6ntcgB6Skg2/CQlEGBWdHa/uTb1oiv1AQbDA2mUX22UzX9xmtpigXvhMZfogXT6FMh
HbwA+QiJBc1XdJSD3wzP4ya0aAWVDHKRZpIqexU6celAqSgb6THJRWD5dGd175jRIAn1XAoK5MTE
5dnHF10fvspaqCq62tqWstcd3Vh6NqF4JmPSVa+9oZjFMyB6yoSTnAeAS7usvOZCumd48S+zxO7D
z8W90QMyOeb2oRXSx+KBFCp1c3KZ/ImSzgolcGz39f2yHMi17juj7d/AelUdcAd3C0EqcF+csv6x
UgaGU6ksP6g2mmGKd6v0JjWVL0EoTgaAEk3H12pGkUe3TfPoymT6KoA/l6CddBCubCKZ8an07FFz
V1LuMvzy9CjVOTRgxO0oJuWh4hnUTlrSSdu/j+KUjAk3yAjPXSJCuhPnOMv9zWCkgPi+LTBHA2nx
aJc29THLzjoLZUZWZJJPro/2X/L9gvoj2solbWwnWjOSvDObZzPUwCyCOwpRTEZcU2pTR1SoRHkk
OV+FnI0mPnZz1wjWltsZK9IaQ5B0JksD0UrD5xbMHQ/KtpGA4Eu4h8GA2UhMZlxcxgwI/Ient+uu
LRy4zRxFa6069XABpc+JfkQ1hu6YnHWCp9ebzH//XtOVQrNDLh+odI6Kfeg7bWDbghi1vYQinDC2
/vxvRBHVt0f4SFDep54lJ3Kka5ffYlNpLAoE5zVeX6jAUckHDA8Gpzt1d16rexZ9ptqOkCmO0pGY
UGTTAj1rUbQp2Hea50rP5et0RT9cr5vwfIUscglrMNzwEwU87nZZLzJj6w80utHmoX4ketNcxc65
bqU2JKPZIpHhJ5k1IQkztxTqeT0M318L5n2nnebH7140CU8dDVmj0EGiq8gBZBXqVKhxX6Wu2T9l
gflrh0KHKxr1LuHDqvUeNWf35LU0hXgBktrNWARpMEuJfY2K/m/k5+nkJwpC1GaOaUaIgI9e/SZx
6ltWr+ibs5gFbfhsSggg69z1j0mqehQKL9YO03NFGnFceRhC3vQ/oYSgay4Z1DKhYDkO1NM9m64q
Jpb8eGs2L4bQaD0qTsgwMYCi3c3jO8OmQR7Sb5wpzPnwIfEJ/Ygyo56glnhkygscTPEk9CB4JYnV
c5ErXwSSBagZ+H+60KfLjAkQNZrUnBpoDfM5ItwYgkbxFsELzWVZ0/vN0kDw+GtXeReuktgijsnK
IZ56sKZSpD+FcfMItFEA3GySkT4V8Z+pujtgWXUzVq0fvhDln6zPGD48qJNi+I7D4bJAAs3qXNwZ
I/YfuuN3Or9ym17dJWC2e3xWvw4HCgVI5lWpyrX+bH2K3vx7vTp2KNsr7I8yY5JFFE5+8Rkbu3AA
7ya4UIxwOe08a+3tKoKw2Sj1vz0WlXlsY3lnlFJ0PaD53sJ//OR+6FqCUxlQ1bxJKcezrdFPzxAH
uTGTa6W1DzZsqqsAyW+S9bYMbCi0UkUpBEzdcJqb/0e5O9g1+s37XBHWRQ3HHMJ5f26I6vuDjrh0
9MsUuc0jHTpxPfm9eZ6k38MEERTKWAEnGoojLzEmr2A7bDYM6CyAQvuxOckKyJh5Y9hqtcu2u2HJ
hmnXcjSwDyELR4zMOYpl4kvvxuUu63jqZnhTsYVPbWJX9Uy1QRWbbzRTBR2GRFs3zzt8T9e1VaXh
/TcJ4skQ3+tVaojYeffnzKzN5vksOmGAuR8x/K41S2wnsLXdA6HcxCfKZYcdEBeBBmVjTYURzFv6
NJCKZP53xcjmBmTbizRvQR/Hm2KBce+z2iaTU6Efwrb4lt2z+EtRRVDoEo7X4bpgeB+7MIzOtNH7
B696qU/Zn58ENR8Y/qUzxRVkIcjQt2A616+hEwrJPETX22gaNmjbajDzZFYr1wGL6m2BsCoDvgoU
2x7N/F51nu8Cu9eROwYY5RoqdywlNiHHNyEwdjlw6BKSR4PIwP+coNmlqh2ISN2eMsYvwtCn209G
di3ZP/2O5zWBUkIpTSlmo7Z/2jPLWisNP3xbPQ0km8eazFyKwjNpcK0/rccab/0Fx9wrRgss5zPW
YtpsIfVHkHkCo2J/Lfo/n35+gyt607sUMRTpOeCHtfOHoC9r7TpeTpLKiIHkcAxcabYOZLxJb/k6
9FJVfYZpj7YyeHddPC9JIbo28fJu4Qa+kFiDvBS5jn1yEPFMEpOwYVbM2sJLsh76OZ7RcQ0+sTSO
8i9m6HyyqkeoKLAGBtDK9xAFNlX4uxvQGWszIN7h/kd3RFRzGPXxZIe2yOhoAbkzdTyLzTgiOGgv
/SDU6Vreu/wf9dp8+u30H8iEWhurneanRsRK496b3YqDdQp1njqrFBrC/PN/Bnw2oa8Av37/Dfx5
7vL85PZrbGlWZhUZFtJ9jjgnsLWbTuybUnCi1PO72FhDv+awjmAdz8WjuBuoOfDhTceyuaw712Ou
tNqyH7BRWW5bJ7TnEwOVZCZZ2LBWJJGE6L3XS5KINMIRx5p4WSZMkYPvmPX0rBqIN0hXt6WbspvH
v9alSsLX9fy1abGbGzf/wUaFFDSwSwFpO00CuRPM3Wa1eVrqpxnPW9KgNN57g5bvS/5543My0KT3
cpkjSrb2u3Rkfz1DaXNbC4TyI7DuS32uKe/BBBf+a54XaRxYWjG0cqg2fOvzbiG1YlB5g3bGNgtI
dV0RJCH0023FsCLUZaO6VOKW6BhlHSzTSKepDDalABUzCxat8EMQ8UK/qTYRyrEMMPm7XOqos2c7
W5AcmTtV0HfiIyZH01J+04MJWxJ4WQmxwdS4a8LN1lJUF7YV1BHrChNK4wgI2UChAtLf4Ess51i7
KGXBTqdog3JIYtxJ6WNKgFONOdFwVxDVOoRXpieYf0Oeg3BI7OyRPIgf86+d87eaFXf8jrhhz9Aw
qVE4D8aNFfNTk6iu1AW5ozW47RPWM2/TzRMj8S9KHmaEzLDfb1Ev14p30JJprSJmLhtDQQH+ynWP
ySKrAoXys+zdrpqMBUS7eomv5NReHs3cgJU95JVSAPh7MQlVLutMSmWwM0+bObHUsd30IHQd08+F
f4sWjSdXFjvfkKC68yhG86dyiK7yunUlM0mmLPddES8nx15EVPNwB6fv9b/vPWm6dzuUg1bsxfMc
qvGLCXmJRI5eteQgyOozELC2IRUcKiKArgsT2tzNxbPZyp2rNPCiCj30WjGUwYqTFVt8jNtQxU2k
VY2Mx+HBsI1aQjGMfa2mKXYIoPs+j6Nro72/SsBFwI2usSnbNpbdZ6IyGkpoX/JuTbK4OizMrpmR
Sfg4Qi1Vt083v4dkj40f+dl2jpuMBpK9rPIf0XZ7KaXJf3UYjFONb8QwA/8zXLhzJYfNttiyZFhM
J46XfecX7/Tl+BPRbIzwFFBdC0p1KmJqCvZWqJCNa83E1TDD85vosaQXV33iJnjYfGsa9rGKOlzY
B49BYBBoGQ0U3uSsY2Y4b/zYfdwKqyg4QKnX6GRbeb1Z+RiERMSQUx8KFQ5CKW3hOjh5pgSjVed4
ERz0XilnL7vve8S7wgUZPSA8BkjuH6FfP7YB36aaEqnw4MBUuKXRYbNfTZaEqTPf7TeqnZ8YOsMK
D6B6+93lIE1s5Ir6iWPWpc358tGAA/OHkIYpaeKI8M7UiAyGrtmcuK1Cvrc+8Jo08w3V8YKSyekq
LMhKDgtb18cxvjM0aJVpZXTjVpFT1/lIuXsFl/QwuXeB0zZ8+k79Kbm+XVZ6sOBGiDAXLwILCF97
Qq1fHKAgcwoB1bJJCNAnilwAkcKs9L+cg0jxKSvQCBSOnkKYumW1Kapx38ckV41WXSV8JhhmWArp
u8zxADRmurKnazEuHJ70fPxqTW1LtGfVGnVXaX+DXlQQl6WGSYMojXhxY7zggZjyWlhkcLq/wi+Y
dBmH5D525oW3SHkOaOpgN7ng11xjLcuQXAfRz1/lJycwsjIYCtNikUaP394Dpfwubf5fRG1cY5BV
Dxdmb97E1kyyM1Ujb6eBPbZOAf0NJuzfBKbH2vutZjcVRBDoHBrdjXXDxYa42+ZeTJ0YBpY6a9lA
zimgjQ7ktzdxsmWGXIuyPll7ZllucIUn/kSU6h5S8y0CTOQXUeOwMfCt0L7b1TemI82SJ+aqQvar
BR2k+WC3w4WGvxqH27k57ch33KymiPySfLo620gEYspT4jzjSofw/xnm8oaRvHga/kuyCn2/yK6/
dpGoh9p9+zQiENTZt0Vdm934+JQ7z2JOF19vUQC3ad05JL1KzvX0EScVEZtpIujRN813F0zo6anu
042f6vRtWVT1Pdgf+WdoFHA4RZfQI/Od+6aNYoS5AuQUy2mnADO3xUatAJxqscCTkpbk6vFkrLq0
gu0OiZTsFGLZ830bRGQWcWi6xup3hbBbfqGL5eFjG8ZVa/cwr9908SyJmi4jwmrxumc9sWe1l7Rl
EYj6BQ4zJipbYvCAQCNT3n6evQQcBw3ggsd6BcmmZNHZbIzUjXYoDsIzRuros7HdFRcKCtrr2Aww
m51Hu+L87yQen5Sj+1dQN7O0SjNcrSazSI7W+YVp3MbDm4dD5B8fnx8W/LVnDEYevfmV20Y/EAoz
7krdrClGrEfWClSvuQ9UpIaRdcsRnNYdSvseBCPN5ZHnzLVNBaKNUS/pwwK76yIZUySeZOBZ7I9d
EcEcUHw9g4/yw8thauXkggxv7rQVuZrMZJh+rneIff1NRB1EniWrZfwm9k1OIGxNGp2Er0oT274X
pWuSSNqjWqAzMxFoRgBeKe74N5mOty79CjKN37RfXpblrNgB1wihTlQ5GWh1XCglZuaqPoe1S+jI
2L1qi68weGIqhE7haX7dKdetPZDQ05RZHBnqmB5GARYucZ5FcEX0i1uafEkgK8JKkemFEawPCNp3
5YigHF4G68h6YMctTyot6rm11+L8n2zUUo1SEt0jLhz8ohSUxPdq3apwSH57HqBMddCcmnDl43WN
J6Pv8EOGCgP3j/Q5rZ6lB4cnhxafo9hlHNKlUSpMox7V508QgmlCE9d3Rj5/BTi3oCt7EOSh59bQ
OBrV/HVvLHqGrMUFzFokjwFfXH/JsF1/VY/UIEab+V1+xVhDIZNJb0d/MOhHS8oeVEexsklrRU44
pGF7nw2ugmr8RUzcU/VPVNXa9YLy7W58e8d0J04dDarknDbg9JKGxch12UQGM+szKn8oxSop6U8g
WmmG7JjMu4ZbArzZtn0I21S6mV5978fqW60PVL2xhdccuKQxwCdpHWcuaWdwGqODDMzsDnsSBlT3
UKaPwSoQ0hRoWaFzm73dH7Ue4Hs8aeLoTS2m9JTQzl/JV9Q43ut3rEUmrHRw7MkKUqBxALPasl3g
A8p5gPmVCOVBSge2YFX3Tr6GiBminN7D0wk/6k0X48LLpMn+BHmg92/8G46bkVrff3ioSA5GWUBs
D/s7R+hs5bJMXdZTQu9gEjPRwD6AsQSTKHTGAVABTfmdHnY/p6GKcxPVirhoHMoZfUIRS1MBnfYK
4AQR0/piE7qvkV+JnQph5I3ZZKvap3FME5hWWSkmSmZJ6Tehse2V9iqT62hXav9BjsOc5Zrmxo/U
TMXa93r9qUo505XtU+LKf12MSH69HiPhnkbi4WgWgF/t2/F7pbTNY9YldVbmkwFd6Al/Nu2kCye4
vSYEsUSqgGCRLWN5ZO5coOCEhED5YmMNNGVHhk9jWWG9w2dODkwJlJAKR9cQBibtgi/toakHYWnS
kIGH7BhuJs2QTkh1bo7fnBXpJLI7IXQ9amQrlBCdVBPMlm2JZ8pFuhGyZwNOshZxYfZRvoViVUYX
QMsbP+Wje+9uE5OAjSJDC6U7ZDq4KysbjzahbswSYY+AK5D4rl3hIWMUzgU46gzIbuxIoe2Mio5S
zjJDOp0oggu9cM/xCarqZLgH0LeQwaqGmVwIG/R+4ChbV4g1MTlW0Iheef1KvFnS9ls1xknFD1I4
NCiah+7iIDGwGFQu5/OY8UjAmzq1zVd1l6pB+XqX8vWcSkygTLiy8LonPQkl8pPKNWGpCZnVLVox
/4T7Vi3eMp4E1xExi2CiryqION84ubjMvYd+S7Any0dSMD85YKvD36QaQnLaoqt3n0+aEn3JX2ec
LzWcIUAWJCpGJSo26UQYX9qYFt5x4p4t/ljx3zBDxkEt4Qv9D+qyYpvau2uF4uumEd/iCqVAvsjL
vtVN5UhEm5Y/TagUlpV6gSKVijAenoV33ncjJYCugdEZ9lbd3t3uoHGUSwRuaEZVJMwWBf/5tp2v
D1CKfXz4NTN4j5pJwU+pYEAz9L3CDQjTyOpn4bya0HyUChaFxstqSJsLDvTqBt4J1pyYD5CUqtV3
GY5IrM1bbdH0hECBr6oIW/q9Mvq8sANddrs4BhYbDFsZsxDmrGLgy92AWr1Kh0NmOYHXcevw70e3
5FxUY9zoZdlsELaiKSaKGaO+8v4p5zixQE27PY7gIaVaHPU1tNtvyfvI/HUxjPrRT2DAO7vwpl6e
pe1o7h3Q3RhUyZMwYKiUYvrSjfHAdAGpTtFPeWjmLPKcoSzt71ZaEgXSi0smccGffEOyt9CiMDer
MeWaOS0Nk3DchppOUs2JL863mLApWDwMm8Snz9w5X97jMlCS/dBn9cBqC6yhqJD7KDPga1tdqyeM
4v3bH3gwVwjIAaRNlX/S3I++TUId+oZieiqERHwRyH1rGEe+C6GpmS/Tpced8iKTisLMx7FY4B0O
JUcUx0ZANOFssC3QZXf82WNqwMhgotVZTiesL3aMyxXFYf9+FsHQPv8Ia6l8FcSLh3RujjXdODYd
voU1PrJZkR9GjQW6RymQk48LVhuH4+4aiib8NJfclHq5JQPdk+8dQluC558VA9UYBQRqrdVvbGUa
C7iQjSFjuLFDSlh1iiqoUxc7yUrNcu8z1MMrAbR9RqCg/Tl+EBeItjhKnYXP/vCnjMd5hVXnDmy7
BEDDxVWb61S+6OkWlzNZSbKia7QZbNa3FttZDxsJn6nudWUkVAAHRtYpnUNMH9HlVpkJbKWywAiy
Rp3ysCJObVHqT/ZTTa0ViVCcqgHZa4rESf9JEVH6eN0VAyz8joOQZvtWTvje/B9mEc0ovgQASoVx
IHym8vowQwRbd4qh/VBDdb906p+sVVRyBU8bWNF87JHP9ewTrsies8YbxSruF/uuk6GAJ6Fh0A5z
/88NZFipCMD6Zk+uyTR6nKLfJGX+3bCmyiVZ6AvDPpW/nHf62QPayc2ZKXezvpyXYjLHFdbHSraZ
iw9wqI2U/ai1O28xRdYP+z4ykj+LBBP//QI6EC6Tl0+954UHAIL+k72Yym0BVcnKkdwPBuwiKzez
FLfmNrMknox+BDu9ii1XpszG4K0ik9ABoA6bp5mH4X0lr5GEA4VEOnt7SsxS/uLZGIJbAvrhNiSd
9idERFA1sNRZICl1V4QFiIgnvw816viCn0MoiMRSvRq/RiyYsR8k/nZliEsmDmuClBtZLoJWm54I
Et1XLnp62PNEuwsb+8ZKXEaoDvYgiTBTlcInjqM9WVFxaZ8YxmSo/C6K78mSl7n++lVe6xGcBp9C
w1MpgXjNtM76vMj9OxsI0iWZlHFKOsUVbTVwGf6LxSpQs/WlvG72fI9fF4HJJ7j6EPXpCYlR8xmX
55hF4Gae76OVhvYbMj+OWrUfbEqOnl8AeTAVZsBAPpCJPi4BNdA6e/eD+YRgjGFHEbk3JE6F2s63
Bra+VDekfgMGwpQZaKWRqurC+d8/La9TilKnA9gjnZ9V6MKdeJ4wFqfNqsQgyzXUec+2DDzYpsa0
1fNZDC8+xxPGk6m/TGrTSuSCGAgQBrDr/6NRRNOkx3um58czrxjx0P2DpaI8/5DH7pMZD1Spa1Er
HnwwyusSYKLQVc1IEM4SQjf2PjcRTM8o5e0pypUqUjSrj3DMeMUDn0uWYtU9boxZnhdORg05SyDl
vFXZJTLbrMpGvDtXs1pjZjdqnzQR5Q7GRRy3DsNxlgPkvK40fgqw3QD2KQ1398EPo4h+RBnDyuTn
Wm/ANIPVb3DjGcEaD1BMHjGELKbnLROgzQ26Kk7bDZPeN2cR45O4V/ZXqncA7/mxIKnNfrsaLMKr
kYuDpzuGPHyqs/QpLZ9iboIg3xMLNqcrSxG990fQvQPoeOSeUx0+GDN9HQCHBkTwBrWwU4ULm3YR
li7/dYdAsIba3mmZZyOp8g4UFPJ/DWzpIqSDUnmqAQSB7etAA9hx6iW6/0rysZ7U4eBhIcTQqJ7c
6BdjaDVhkHENrZKFMRGcFCMTh8VySE2VeidgZhVLWY23qSOAnVIVYwTXH1e9X1eco7Uxe7EaKqTn
kLmQ9GzFda8X36OWO+CJhMiWe1QPbNDB9ro449c5KJ8Z9u73Znox2cX7A0+bBDX1bkgTYe3sA5M2
4CGqH7tp17tP+G4nCgbFh+cjbSM4YFL+wx649lI/M/SczNXYn/wimjYIlatoEOMqvqtbs/jLkMdl
Ip/pTXlHsnedDOBA6xmtvTcPJZnpCcRRj1rgHCsxAkAAiccdtcOqOiRj0EBR5UnOaJA7oAsBQnGR
K9vTikVQsSEdNOZ4HSk81NvrA8MFYXmc8GKleAbUTj5bepiqDhYWRlG9CvcwkZ0yMVuVoU4H9QM5
nYMMYhtTZhdNybzvx+NHpc0ThfJKP0hjyw/B7YrtbBgu0K87pmkJfvI5BQvGq2AWMmx+hIEcrtyK
f6INPtE2fH+yYGykvujWrUl0rR8MN8bCcVu3utTB6S2u3LYqDByqjZemxEmqgvChx6NZecOfwqAD
aRjch2F2gmZKB2zn8tDjEpSobCBVDlY4hmQovoFco8nQPZZ2rLeK4qLEV/wGqaARUr6rWLTySCv5
H8Jyv7gzeyd+ceDU5cdFccDJpDV+n0cB7O+k/GnuMiSslBb9V7s6yKgLl/08CwzkWJeZ0D5tL9uv
VM0fmT4djZc2ZvCqcL/a/zhbR9ERWUKKErJrktLQG4kWpuc/l02+e+VzZhtbVLM58ph50Eens4HU
9Hfg2GbQyz0LcFBYl4rBe6VBwpitYBUVd6PkXeaTCF6cARIonc1GgYrsL/L8ya8uB7+xqQpGnWUO
Yg9jCRgFU44CWvM+uAAiA89g0fH9fzF28I0J4mhp7b+43Ljj0leraAk6gothBGa/Afm7heH2x6Fx
7gNGu1CUWs+pVlXp1epKhE4XTtbe9ZCbpWtt25vDS6MFHZHbHjhEYA7JhAhVGjv10pq2lm2xYT+W
3ArwtjGpQLWNlcudFL19PIIRKSZM5opFbD+rc71u3GDO6XdPeaoS2eYjwgvQ/+9zDQTtXdMhfPyu
PBTrfwQZhL7um0e3XE9228+WybqPcrVxgfbYS9AI3pcIMIhs7qFvuaUqv+DTIMwBKTyh3jeXhZWG
HxmrrnA42z2062k8kDvtbGNXQnhdoxp5sDb3FEBcD/0UIIDdhaD+hRD2J3fH5SX2gMar1hPx2cOE
lXHxOApfIuXnGLfEhhs32MqmS+Eybxo7ARuKCmB8Wo6KNXoKPMaLYBTqKWkXcP1PXvadwRq5COhZ
hjyytFFRtSIVz4diyLqjA3UvP12J4vUUVkg3iMEBA/iiK02B7VY/ZY2wLpFVkWK2KTl5pDbQ6mEO
cOC2yDDCRMgy79ZyDAY9GPiQVlHoucx+IO4CE81FY1K4VFoLOJ1jDi6rwTKUxMtKHVrdrIOnkG/6
wgxHor+0YYfqp8PMeWwkbgs72epph23NEk/mIw1bcaF/XvEjj/9qVDClvrmBTX8kVVO62FqDuCtg
kB0z++YisEet4zCYtofpjKE66U3RetISus9cTGP42x58MA6hA+tLZmfudsI7IFUoMyoKw1E9JhKA
3RwyOnqU3HIwviDGlX8kwDYFtNqCCLGas6xDy4c7CsSmXskdrmxp+U8kP3rKzlzIYgCrIppJ2ZyK
LaE0tq8KcoWioGdvV97N9GyO27nDSS0Y/kpm27YDTK5YzmLkrGlbvQKQCSifBkeks76OxBP5MbHu
DF4sismIm8OcdWyzelzhO74NWnovKTTp5io/nYlI+2WEf5cKFwlxqAba1WF+nxxq2ZcW5UsXepRQ
xLHNEpT5ll1YYZQ+vQF/PyjCAf6gnCOUsmt1Pb1tfOWKWZ7MrlnrhJogBqaq2V5lskplq1/rY4JL
i3AHx1RGN5VIBwzd0f0lZMjFJB975PZQhdKBcQ6YofYXlixDFvut0EYkMW7ATbXxmdNtTpLRA3N9
dRU15i54GWpi47JUH44DQNzjlJTsVlbvKxRo6ycw26E3cmSyXmQOxlH+YHjyOwXianCQ2LWpxJm5
PLIlDiGWdDM2kaV3efY2PozXfH4IMZ9aQfvj8XXxdei9iq2aD1hoN/YyCy/HRbsmUc90bBHnSpWm
94cqlgA0/St5BuCilBfGZwYD/P2EAkHOF5Z8O7iyE3FtzDSyfWA5BrIUxzfVCccoLRw5LvISOyTs
tLO3Gh4+GUPO3jHyr+cHD8W3ek3Mu3ub3NBWm85zFRmoSF41R2hh9KxOKUgADqG5+2iKCRSlc2n0
TvCvwz1oUGi2Jg5qqMPV7q6rM4rqJ/uKsre6DJveut9fBtse36M2pC5cF9HjPPcBXmwyhh7yKq69
/rqiF4JZ6wmzsDfKE6ls4An6Z3O26L0tbRoWQcEe5agJGdMPZFVGokGVKWM4VjEI1ailQiVa5U3f
Pi2b+U/ZnNfZdr0Fk3/vwJK+2+RiPHFCwPuDhxp6XYbt4TsmpkDVDHn8TPSvmx6r+18eFgbrJoYk
4cM6B9xQXzeIl/StqzT+vGSMUf/LZdBWeMv4mccUgbEqUZXF4da2POEJXMWxtgXRxrPKYBniIuBA
EOLWt1K0NL5sSEIyEd9ZuBHgDd9TfUWPfLrtsw+hny84AiaJp8G87wuAmGuIuv+sIKcNrzD4bFvK
7UPIOAjXrMIpiYyqO47lyjE8b5oBarrsdHsHZV1o8wvokd7CMmeeM9UEFMRwifq9NGz68oNCxeNF
NlrcJiNiAwG/WcTeyaNMRJvdL+VpgeOx/FmRJO7NdtFY85ThYHFszvMs6sXAxdxFX1YV/FY50V7V
fUDIIEfqDmz+xkyHDJUL2fHHNqbR/TC6c91bLR5SG4dzdnmqYv+wfDyTYpP3CFyDbzud/5n9Fwb6
FJhy5t4wa58TrliFOn048DbG1DTaoTiAxl6fBGrVw+iN9gpAR++g+w48bbblHG7/0GiUHuakSTso
J0pabkGhz4ajxFS++6SRn/9onRE/fWROHRR0tNrw3QmAdWnWQtuT/r2IHWicqFviGo/xnrGcgKBj
duU6LcweHD9DfIDLMT2zdppq8z75IgjoGyjoEDVyqqwWcbuXXAqvDbz06lRAJLS+abvc4HcRZ5+V
MqtgC9MZGfhj/WJ4fEvXycnYskbH5mfWoTvpujakqySTAa78x2Y6jYd4mcYZqBHvZLcCXIDeXsfz
FvfWj9/GPsdNUKJXDy7jCdsd8F2Q8fuu/fBYRORzVzvkm9RrLWlbcelYrMV+FK0yyPy2AoKS/SSH
LAAWgbWz2Jfbp6DcvBgNioHyJKlf+1VADjUMRlbj8nLT9qZeGGRMkxq+1Trj6HCusrKXUGhj/bHY
cIN/ygzAlJWY1Mym63Lp//yfH5Tr/Xj57bz6m6eE1p2FYzicSaGW8MSoKxPuxMMuweTTrbeqCKmC
rdx8GvHueFvwkoBmjPE5vkiX+t/y1Do3nkOWznRNtNsWFQexN9vDEnd/KElf6jUJPi5SN4ZS6tVH
fKtOHCY8SLv01BI+KQI10htU48ghQ+s0H176pzlDpy5Kwl4RJWevGxCWmWiF/NSY8b8fXh07CQZg
9A7DAI0J2ze6Xw6zHyz/Et20IMjhDOPUc90Rd+Ll7NOomFjoF+1CDnZE414TvaBhzMDJgEctyYnp
sbNrlqxNcXjFdMKRA8cuas8T/abPJINsHZS08qZxgTGslk08/m3L4CS1rbZx/X81oIe3yKD3gVIR
ryjRMv2giZ/fHTb2XlrqTjavse59EX5XwrFzoQqvmcpDvVGMsOKkucbarUHz8BVxnUYRlN1xOTfp
N+Q9HH80UBkLXztvVcx4wkPWBcPGpaGBuPE1N5EFN9rl/HZjXZdoAlnp8kXb0SHhlINvqJbCHbHN
nU/THtqKHF8blBjz8HPRC5zBy9J/I0GYKxqaEtQQkTy7mY5HPI6o5DYrPE/dgH8TA3Vu+avfUc0h
9JFKFQUjLdNr61jC6UNGmDzbWnBu6rrdgcSJon/8rZxkk8pp6rT0LjKas1CC9Y9ov1vq/JTJfl2p
8+JkzUxOs8G1nUxkmSOVbaQIHOsj1J9r8lQMxzmoaZ4ghiO6o0W/9YSIK2TL7nHs/EZSx7/AokQt
0URJi7kwcOYG8MNQwpmqgNdzLkLwB1mjV1BxdvTVP5CyfpEjsgB09owgpWcKEi5baUUZBYRtpmlJ
O1dLcJpn3iSqY0Uz0zIVBg+3OhXviQep4PyIy+WgD02XGdXTkaGEUN1mhRTJTF4HB+uBTxEKW1DF
on8kmo48Nb8/d4Kq6+2jZSA4rrFWcSGb+k13Z8cW5RvqQdTKJ9c9dxKBu8svOZsDTQZ1Qzhhd/eJ
2F7XAR9DyKsHeH3gSOlwSh6vOWJ69uRFB5P9298SutfRQURqcEx4h8iAIGIvsk5Bx74leJgNDA1N
KhKdZ8tUtvfUkF7qiLRigc070LdZ1uyXkV7MZ2oJybc4a/C3XbrqS84OFc4PWweRabCAQDNrUCLC
4D+wdxnw+lScH+NUN6oRWDWwpYd+k5IFSqcDiOFm0MxIPL/dgzcWVqdK5v3TGTdfjl71hbijnWB3
horMlqhXkx8EcvJQV2/tquTKxRr/iq1FkxLwAAdmSysZaGTpH/43btkLkfb1pylKdROAqoF7pZ9D
z8H0K/ccaUkFoRuClR5WxC1XHia8Oc1saBTz2EHlDL6d0gh8XLxjkfZChEOXNmqRJOhdISLlj0oC
S7fSm1bYt+ZNVzH2N2rVZGzGFoLioGCli/RnDLpshC3Kv2+4DJuCE0ltaRdEYhwJuyzvGsc0yxRV
VBOgiFzXXT5s++ReQ2GIBiB5T/zaAhbFLiBhLDldqi1/6NGNXQGfC7LPxYX2sBl6yQ/tCvUhbXED
f2FthGnBZMH4MoWAXgLgirsTQPlvvO/2k96/p0OLneCbfAR63ZLPYMy+B08/8FXDQHl2dVfrDopN
6PIOCWasXEu9BJqihEP9+ulmzFJe2CwQRBmuLYuJ9ZMfLtQ5Rt/QXWgd12xT5Hb11yrpQX0wxnz2
pbr9eCQnqap/Sc7cWcSKh6ZhjfXsGRh2pJS6TZbdo7ZU7vGT4t6wEiohnNyA6Uwvs6iCWx0aZOfJ
cYLH9MiOLGrqG58VPRcIP/tj9TjB7FlTizlYtf79hdwQG4F4cgEjMwq57PHus888gCLu3m/+eZu/
uwklQ+Uc72+R2nxQq81PHupYJdcUWbhdrVt82e08UsvduB1fOKDxAZoiCHlaWs/Q8wuvuKKULjfK
LBfordHrDFBPwV768M/nsKFOwK8k2GcMIxb5tjDbjFLK91GUZtDwLTfGGyJk74GFUcAux6xCuAok
m7RhWmKu/+BGlTVDc5sCtCbt+NMLLWFe687LPnb2tZLkEZwFfSQIkxI3p1ZQ8znPd8gRB4CsQtCy
b3VFhQNUYGA2o7WJHQhAgHAChX0hgv1tDFNMiJk1Qwws34HnXF6+zvGxhSYAjm2LNVPI5iZfpuGZ
C4DoH22zm5YrPdUdTXvXfibruFZsE1FWSmpH2msW3yDpAigFAJMWl7uqB6C8LadrmWUHE6VaEld2
pH3qNISxP9/Eh/3pdKC8hAD2c+jOpCxZcHlvqx5toCvK3EydaWoOEpvxO++5u7J0v7AtYsiLgMPE
FehjBRtMqFl4hB1ZXtk6kS4dGBL9rwN3z6vU5icLxPQaAZ6+JEX6zgHw4y60j6zrMujZTiy4065w
LwR3OLbZ348nxH29u7mLYb0qmet8sgrJaVMjbAvHATYtmR7sdeCbZkEtcJe9S7U7uv4uHq2ifdzk
19irMyzHV/UGAoX4UNfY3WSZ8B+1PpTivjtpUYGj+WEZPDyMn9OQ6MDu7e03NqyArXibC4IiSjuW
dFYK/DCMwPPYl5EEWMychPZZIVo4gkLxyYNTbuJpFB0uzEc/OA2o/DjvkBv33DwfO4j+2YRM9qO0
YrZep2sVRDLogIjvBvPKHU4oIg4XVaiBaMner7rxgtttPuaFA/7Uo/cAgFGmOXWl6Ov1m1z6QSLF
FJZXEFyR55iWb6p132d70+4E5I4E9GbkK7Tzdx0IbPVNPpHI2SA+U0WSlRqxwIOB5BB7VC1BK9o4
L4C1u5GT37q6SiNJWMK6ZaTP6EhDq3xlbMczPyFjPyfEIhhvOLCn2vgm7UINBj3Ncj1AJeiGXrGy
ORhyKDX7nXfirvlUhUkbu85QsqmoU5nS7AbJl58tJ3Xuwl6qmdXQEqOOKEjwFAufw825O26RWOVY
deN/EU0CNnZ8PY62hT896CDnqGwDnZTHUhOGoNRLHi35REqVra4Zf/FAlJKY3dq6SrEHyBzZr3f9
DBKKXaGmEDSG3Mqg+eJE12X1PenO8oj2UhG4PrzhNiH/UwCw/8LQEDDZuXyXPqZuMZPyy8uso1NC
Y2AUqgIF/tfz/zn1FJ3vOX5YZHWTiXiPJ/RaA+NXfbp6B0oVaaLGzWy052iWvLP07hF7ueJ9Lb/F
2pOYKGwlS4Gwqvd6h42rpuN2Xr4/dzuNG0Ql62Rh4I1kFBJ/IJ2M8X/HuStll6LtS/CqBqRjx3qz
IXuQ+E9HxnClaWOvYw/C8HuJbwTq1tsdrgFPOMa7SKd/5WqHG5m8Xn5o6LpGRmkykI+F0jDqnY5b
qIChmM6cuuDIM2Zq7ZfRfy/sM6vlDwVmL08eWQ2ygAvftrj1dubKO0Nyk7Nr2/YuDxR8rUvLLoTI
Xjlm3D5yRDcf08fVNE6txjGjPzsNBynMegUydYwg9paByFjTtSrdCVmyMB3dh6j3zx/dnhprDUQm
ky0HqOf5on698dLr3uMxu7Dj3MLyxbtbKHFoj9BtuP/f777Jp3NXJh1zkDUau35kiVLAYVpQYXFy
ExbX8fVdgCfoN651xFNlWn5NXEfitwpYe9h9Z/vpmQ4blKON25CSSzCSsqIyOT85jtRoBWZlmH6r
+16iKA7HuXIhDzAIVodHwgg9pwTF6gBVc4Cq4EeeMWHA23IO1twmSChLvDpzgdrQdTsgCBQbjsBB
S4C01CO/UKcphGVuB+oLzWop5eYR2gSMObH4+XiOZmXvlR/eqllsdb3WvA2FXJIsvaDfJRkxeboS
ACdrbxkFe+cU5JNJSzsG3et/stZ4W/Vw8y2zofMpFbnKGQ+nNbZBsDcyZe5mPJam39OnUUlTrUrW
62Lg27iXVk4wYzBBxokFB4EtRpbW08A8yRk7DTKzguxhQoNMkA3EociT+YH2u0qpiAc8eq7KbE+g
PbLO1vDp/Z/WxIGopMpDjIon1/AaDsLkUfaxZJ67njb5fjLmifjnmjz5Y95wc1kKhxTUdBwApjRK
EzGmK8Sri++IniWwZSPlOD+LUfY9TQCc34rfNptQau9BdSQEQMaIHxPakZ+25o1r4pbD2smihB6s
HesZFna3XidZ5/dd4HPjXOYeM/KILYAPC3+681GAc7YM3kaD+nSrogM+GyfPy6P1LKfo6UwsvAOX
Le7CekbTz7xhaWhE1brFPLFIouMHWgsZznTyIqIBSQOc+kSDcrzoVKv7eropAZ5pWctOOVRTo7sj
rl6bcUJXk/17SU9Bmfvt/+NFBdCsyiPQPJnCayL1ijTbO4Ye+u4R3u414/Tnh8EJiyRVqhobDXrb
f+kBprl8nj4yjGed4wSnT23UG0Mytuz75AoZcasmTEXX5V9Vgnm5vSkFhi71ItyH1EH/Pu7FHrCv
gao9ABgYLADjMRwaChtvgcoRb9hgYHz+fPQA80+J/vnGY5UC5edSxJpMT6dflr68HcZm3XR4j3N2
jWL2fKufUGMspOZRPtuYAkBMMoAVTATaBXRl8YfD2B2NI8MxLy8pUqk85aoKNAG91tI+OqBjbJCQ
5/6dPgSQFfMRXKAAvfmZafEm+dZI8vfgMCqGY2NokMH27NvgqDlqb4vJptKbaYSjsB1lbsikgAl2
VIHtg0vFsRAqcR6DGdsxc7Vm2A4bUULLwf3KMUS9XpH4tmuVyX3OtgHYynE+SqWAOu/4WxjL+0Ht
VLFr0WTOXNVQYOPhhFR0M/lpaAy1eZwTMJKS6PxsV/D1qLj9N0a5KDjO/AKvdAb9O65A4zGGosKM
qf1v7O99WaGX0sFjdMrTvTvWTB8f3yQ6sVgP1NeG4qkzhdP/SURl/C1slsUAwUJ78w5wGziPHjdr
X2QyGwhelARSXcynU6Vm0tdkN4IdpHhFZYSIW2/DiSPNEyKZDuvqfzohWrJTf+oayKHxNo7eEXO1
hlmj/jpnjxZW7nSdnx/QI8xVWqCShAsq2paA7DmelC1C3xwaano5agRiBb9pky5cdJtYEID4PFxV
YKZiPyyZXGEMHQJdyBP4PVNcqf3ODfg+Xtp2sJxfNG+yevEGPlxnwrrcGZJJNWgaiR6qzi0tu31e
7VBggQZsCTuqZqrxHxuji4nqim25H5Ozi1ZH9ZzssbUH/eV8zjgymrceRRQe9auBIfrBe/oxXKB5
HLUfm4X3Tp8qnjC1kgEhw7ayqjTltTEcBASgo9sNep7/qFHosfPOoKjiuhtpC6cjSPex46oG6iPb
NC7B8oESLGzuAo8DHnrHcUAc6yzWsi1O6bxcejuYbVLxwFKo7aKieugzQU6EX5ou6bTMdr/U47i5
QpI8AzochbVfUoGEYx9QP0+86wr+VEjWbTjmVRk8+OLh90HFWKmBNEC1NkebRWjZ14fzL6N0iIdM
FfB+GRbpsQkucPKQSHtwqsL0iy7BcoU5crACC6ODVKXnC4dY+XVHK6yUpkrfY7eb4NN8Z147DJ+U
z7OAKBwfdqYQXXZAKvA7wjG2mH8bqw9vI0OAYZ2on6RHHpO6ZSx8hHKEYVGPOsx5psURBq4PUZwd
9bJ1qJmPLY35BCNokep3gsgFRqsltUFymU2T1neXz6Q/rtqbviTGjB9KFiYzXAhjV1E6YjQTMfUk
VVSvkrrn8vg09T7kBgimB4XT6G5vZyG2Fixz9bvbIqVoH8+Bl1K3EIuaFOyB6nTpqzJNXu0u4oJz
DSdlYS6x5f6LohgMv6VOnIlGnLBkcjAAbqF+nBZq263PnMmxH9FSuS2zqg0EjEoWW+qD+Ullbw9h
cGvgjAoGgUfSzUof8EREmHZsHboYaiaOHRY+7ekx1GZV7rvXFcM4u8jr4DFZ5Rv7B7hwrqjmUsjK
t2SFxlwV+E9qTbkfVl9R5BlxQ4uyxtA+L2puF0lXm444zNeztkadbSxcx+AnMO6538fXpvHSuidN
yLxYUany0HcAQO0esEla3KTjmWpgyWdC17WS/wZ6+6fbaKJH/ZJKYHzXCbdXHy80Ouaw0/v8JQ6y
3QYE6TuK4SWRNRwLbUzuUDdiN9bd+ylN6lzph7REwGaXrVsFJcjafvywHNy0Q3QcFu77/BUc2r6i
JBdu8x7ku8FmNSTNdFoVn5Z5PoG9Fs/gyz3bTFl7ObtQKxGOMP6OyjjiaTNxugGKsIMDLLpwqCxV
Smd0DPdx0VfKwl7rz2y5Bu67gbmXq45NuymvU8gQBatYo4gMrPuCuRlDW73t3aELBrWUWMlGZxzw
12R9I5Kmde2irGK6qoh0Y90jF7dfyXNdLptHgnd7k+Kvt3UHtplyZXgG2XPRv5OJy5qRLDgXf9ZG
wlX2h7oF0Y7FUbJWiC2gYTxeXHjij9xZcBGbHB6QC2GcOjZy/vaDa/HrVwyrWNBBnTqCJV4+SYiw
LSqokatd/kbVfmA5fH6wa9EQr6j2oJdd2mWqg4AkfQNrg8TpU00LAdhu11McpqRhuYOpVkfFQn3I
H1VSzOft99JeH3rlod0ftra8mSzfqblW//+faBu3+mkC7ZyvZsP2kv5/l+Op/4vA91F9lKlTKANQ
9nZkL2iaiB6hdZUhwmDgO9uKujiUan9aVt+eWlqUT2wCrCoJZhGECV59WmaHywXjlAJC4i4CgZMf
Gq7ZySr4cGMq2iM0K4FYr55NbTlt8haGG/9ljsyVhd9YxT1Gswg2RNAj/kmgtc0S2lnnw6W1lKRs
DM21y8pXXMmY0Xg73uZlby93oR9jjivUjNtdIj8By6T77XaNNVW7SgyfJEUz+z1iAyFxgDe0ZsBX
6klxOw2/hBZyiY5nRjq52Gl3Nwde+l2RvGI5/RXN1l9/WsO+2jSDurB9yVkvjNQIlYHelbE6V4vM
YTfwEYQDBQPDzcmpZ7obfBDUfvUR3gO0OVc4HxLtoZhud/33ujxbTY1SYM98383baJtWuMPqB1lk
jXv4Ng8T4aa9D6zT+0Jtue5lEBEjRNDnZ6wHdMSGNrlIgUdnreBMrn3U6dS/1/vaDQ6OcYVuMs+u
HUOR3Y65Kd6teIQkydQTJe5n06ILYm5QkqQrwDq7jmgGCXja+2/ophPo8NM31cj4KiTtSq6bijC/
BIhRJUvqnvCe/w9inq5vulbjDyLDdnxpX2R5i/sCqpzZIwYZG9H6V3BHa4F11X2ufKzuUTNeQfAm
mercKN3pfAYHPXRsmSh6/qMnYak6qSq/VYiyFvdS7lCRvSdY4qChXh4xBR1G3Js3ARXuAGuAizes
6a7QPEp0Ygf+3d4vWrLglT01fdR17pqVDUqjFz/io8e458YQ1RyDwhJ5ZhJERocY+zu46ckt+6yI
9xqrSFAsRJVffbU0tyzZenbOvMwh7Ch3s4PdR9dzQP5tZcocMRNlurRVf9IQ9NjK2kzndOz+WjPS
UNtBTIFAFbDiyJHR4lQ94OZ484xM/QWPMwqCqwx/ACXIIXMMxQE91XpTyLb/LZy7lvYG1dwveNYJ
cJc6Oi75OU3QkF+DAzgWQvvwN9z4ffLsckPthrdxL/adbJmsOBhBUin/50B4/JAb2HWnXFgUUfCC
vvKaT8hROdzZSbEmMmyWAvlU6JiWVHa9GoLuRFCDnykoJ1d4KnL5+PTUggiVONu9Lu/74+r8PjQ3
7U9YBi4GAmhfnE9/Jt+xYq6Wk5Mg7D4zfDIZkTtz4KCIvFOT5TpGaNByfdJtm+9xrNyNp2cxJdaj
V2TRl2HiQm+j25g0G66W9Uo8zUVlRiN5QcHGDlAlGtnVYh57WNv37JVdUYaLLbSnr1JJ2bsAszmp
O6PPnGHwdedt3Zj//jzW0c0ppaNdSgwnrcnIdthyOOvBBCEu7Tpp5Mf/7KYp3er0hr7r6pHF0vDs
ZXAl1VtJmJylSj8ad7HNHNkb9eben7xpm21r4V8CHrAjrJbpeVaypi0ggsIICXckmI6sjPVIsNAh
BDqq0QA7kWza2CELddpTX3DD2UiuTE9X7u8XoDf/QQeW3SYaIT5UlomG+mGXvq/PorMFZBcQiZIO
+g4V05tZkt8hrP4goxlwDHAfwvXVFFc+ZSFDG1fiKlohVETlQ0AXx94rKKffKOqwMhw/8pFLL3oT
tYmtcby4nCwpRslXHGWLrRppoTfcvwHBEaUV7GplTFoi0e54JQWSx+Zw4yoo8EDHz6nNNrQLxkWm
UEm2xbQ8MjVekp4vuMBID1FTkeG0XMtEpN/9XhYOHqdFQsMvmX1OEtZH9Dw1L7lbbomUHn870AyC
Usn5T9/3jw0h/dzsDa1VwUhNKW280dzWz8zXGMqQvFf60p5L+y6CS8sb47ktNSd1xH86U3y4W9bu
70CF9JimzcoV2Tsk4Q3FmKMooZyjuxqUSdyYuVtSkRSYsXTJ+XW3G9YZEKXEm7OrWfPXeHM/6/vh
L3DMMnzEIHRbqTD3TKQcJ4plkLY0Hhb8yFRSyns1wEp9VIyfdFMAdwwNcOnTZnb9PIU5jbvxq4zS
nM87IJnfvJY+KPKI3pPGkgax9d5P6rA0zBKEZYv5rkVRCjbsSACJTcjp2s98Utp94QPfOb0eBk2H
N9AL4gruL1Df3Ycckroi1U+c+DpYD9zfkBzujk74K+wesw91Babwu7fLspVckaYOMZ65NjvF611j
cL1tTbnvZb3RGcmzkfx/ndZ1loqzYDRFhJAQqB1E11KrEo8kP4z5mIEmlKB0JMSr8bHe+YrHqiaG
U97i5bZ5q7AWkWURPUr9c1A1kga6LOkRYAekH5XaPR7a6tgiBMNEX0REtPrINFBlvt74CiSC5D88
cor0bXCEKxYRFleFvAbVbFSavR1SMDGStBfqbcCJaL21Owd1toURC5E8LjZUrPuFnUQigS6pbjdb
auw5FOK1HEyJsu7FQNa6NQFwSyjAP9dXFEe/oHsqRtGTD7hc5iRaGwvYe9J7/Cb3XZDJhCThhdbg
eFSFKPA6RWP34qFSxvA7WuM3NyEfG6cNvkykaGACibASDd7gueULLfHPQDjXDpCKi4Ma9S7GfBEk
F5KbG+rjiBP9CJpyBLtUXPwg6Dvwj960HFQzjaLZZx0cqijpJKjA1yDKV+BCfekEUKiVxbMuRtU6
wDcZ88FM/4czuTmB8EgMbmUdxeRfH6kCtAczbRAmBMZOB6TfvcRSM2Xy4VH1/YOzOjvfnw9vCvwd
aZ/eTjJgjj3izBKa+vqFNrY1X0dFvnSVl5U39H75S+En9yAH4g1Ccq06JQplXH+rIy/errs9+qxM
9xoeWQztOh7/iPXlySy2773R4qFCAjJqtuVU1It2zJ7qs3gCfyARsRdqoglmOTtLkEWBEEMy8fT8
5U220wYPaUVcDohHOOFf/J0EpF8uxwFmwMBNfISKRpg/JW4+M7yA9Xl/zzQGo1QeyR4k9XmKbhjP
wt6BaTlcrP0nu2fzeG9MZ13eJshLtVRDUlCQ2NQdTh9yThjIDRFUUiFSZulva5F6OZDXIIl1bxBc
ac/CFYIhMSpuB0pEmf+0Mpf/9Rvuw6EKF+qsLDr6tHL18h3M9CNdiS4/oNnUCTY5TDk9n3S46we0
i2XwyQGs+Odf6/jM4VZqfNkxDVuCYIGu907e0Q5GHq45gxqaTTg6DKPepVSDYOS7wt0ZccEBICC8
zGzIU8HZRIe31u7yXP6HjE6/IO+S5Qoiou0tXxWs46D2V4crGKUB2PSLi2gy/alXxIEIMxtG9S78
ZJkyL5IqSS8qKh106rwylDXMPGY0qN/Hzxuw6S25++86FDkimXkQ3dPeY8WLwBqK6rpkHHNngZFv
k81zUKXYV4BQCQV65fenEZZcqHIv0C2k2g1E9EavXv5lwtP0WPVWAkvg864H3wG8w8O8M+dCAynF
U+pa9gweazob+JL7p9Ryf0sctYEI41+UAktlvBuE3mxWWmSePK7lIYVz3BdJI8Bm3yw2SWyGF8Sj
iGt9KDaGes/x40HJ/BPOGeYEQ03IBKzXIPAi39TFD0sA9azkFAgtLjde8W1jLvwuPrg/gSa9gbR3
N4iufsgTCTuiC+LQeMVcXOC6P+rxFdRlr1ra73giYXVuPpQFMBx/2MWMs/6WvHFIEMtrAsZO0LOz
YnA5iEC+wyiBfkks8tHkU87wf6NfTz2Q/EqXvje0FFIz8o6GZ30ABOYm3Po0+4n4UflJ1mga5QnQ
8ZuMRU/hea9GihsSSWxNT7ljNtjGzxd4Xw6pwPHspb6Rad3j/SM7MBAVQ1H+zrTsik45Yin9bEFD
vyX5FuwIc6+91Eln63BoQXlwt5gzBIrY8mTU2JLppMxkyDqw/T9h7pfmsO7ZYN0cCY8zXjpfoml1
wbEEqTI1XFlqNTJwgq4RmTfqqii3F4jNSRiBX61heES3u3TX69HVmvlvRTYBYtBdS6uLRFytS5Pm
8+PzOByLSciA1XnCwCfHXxWEUpkRtassif49CvFa/hRgBKWADAw3jP6i9yCZCB+1n21/+/rlv0pT
76XYiXB4DpPQ7skQJeKIO2WEQz/f0oHQ6GeAxkSmI9sZ7fDEmcziKt4Zzmq6xxiafJMTiqSXlrr6
tKElfXvHnlyM9TUk7DE5TBOnjh/5uJ8zFDhvsNwaG7hYMFtU2eRgvggdkk7rEfDlg3cpRmpvjAON
uSlQ2Tvekfm+V11QQsL7fsFRSwT/MTXWKUBwTtSCRyysoY+Mvvs0o1bpSZzeoZcC2GOzijNo89AQ
fQBN2air/TprSW0xFEvHkfa7VRoPgAqG2241PjuY9FkCd2x0FNtzay60yldJehkAOqHAzxOAHDDx
GWhXRO7fOU/4y8zjXn3Es6OE6qCI+AveR0Rm4Vn+8lxWri2ThRQhgOj6R0wAfWWWBljp/+D9fnhb
DrajeGDJ+WfkAYOMDELUsV/isWNBxdfcxhHpKW3UY4kdXaO5BnPaeJrMndBDlSaUxseQk8895QTd
Z/WqJjUGPOw6xmGRLNSDFbQA2GQMRFL/67ZFVMHvb9oGsdiVNPdCUtVfjFkknEMjUetnxBJ4UiXI
nLyckhMKLF2RIHsPNBoZHGaAQVdpX8SuHtdifWgytsqlSdHgzTwx7HAwUVmTW5yZYClMgRzhKokJ
cxd6qAYdAMzzySKfaXvaPLq0a5tyuD1ii1u6gh1TyNKAabbdn3mD+G5FC6TD6Y0/7IrwV0F2tcyA
sxqm+rU9XBpz1Wrk6vWfS+ZGngLo1jVsrxxjwwe4owC0jjwnwhkxMR3B+vvW3BQppKKYLNCCTMd1
8MHXSG2cv3Iez5Scv3FRnMBQocoLqr4stprznufAbzDBegM6qbVCx5fkrMByFwLdeoCrRveA/V6I
EfdxYJcnlDKw/bugVC/+yvuxh1jpIL13R9RwIqsBN0rJeXG2T7NiTA2kwuJQw3Xb+AryxkX6U5Gz
ut69K7AmLXh6CsoE0CDly6nTNmG07AHM/5CujjE2MVxtEY3Rwzy6iDneF9QtEIM5q8A/zdU2MXA4
opZG15T1YYjY9QPv6scBZMqGgJ2RuhjByoLPA+OshHWYK2e8sQHRIekYE+OZJCFi4HASwIcStQYs
s33rKZQl4zITpNMV+gqSRgj8jG0ECbBPtsYiwW2uo98xqza6YTmfyJDidKARPFENhp5O0ok0IAwA
VsZtTJ4Eq8eSK46bf2OEm9jwwsO2L3r0/IQ3NyGLd4okc7qBtI3IE/0P+HhLsy4N/5aj69Z5W9b7
t60REQkGALzWYvRuygIBANcNhnYKgqix0nehEjylJvll4T6KBrpxemsWKeHJ2GELg5w5YZfGyVTQ
j0pPlsz/qFaLLX6I2iNOdGWUuLE2ow4cZgtQdDFMQx4ZlJVcpNpUhP3N73KJVCxvhStDJx/CerDw
3yVrVoaDhBP6efTS6lK3aHwRmE9QG9POJbJaD3kCYFp3GgKlwPVhaPt16e3Dd9F0fpGgSkK8v2ie
dD9CSO4N+JO1a0iU/MRY84hSwNVZEVVdGnlchEhMfF/jxsvwv4pGFOnotP9fjhDjiEE/+3MHdC70
gj4mIxM73kplpnsJwyTjKxA55gWhDWtvNoUT8dPLAmLkdYfst4Nj2ZZKD9+OmsulFEI2ZSCdXzwC
+5dj8JdrSmX1o+oLD4VTqOlBHH71KrEyQ+0wprr/utPOOROt4c4j8N0uk/ZzxoCK40XQT2UuO6Bh
v5bY3CkzhdO+H1PaNLkxKRXBnsYFFMM1oz1gOwyN0BVMqBofpTB/YYxZgH2GVPHDqH3quPZfXgfy
IDaLV/uXEw2OKubdqfL3/0tK6MCgCBt56QHwfxnP1+yZqy+NsmA+/XV01H8IlouR29DilxXmENS5
KHg/Lmrc4oa6Hog4apmYForVvZh3vk5nP2f5iWco2e5mmxC+SIxzENrrsgc4bASblQNdAQXBKYbY
0F2jWCakvwaSwRt36QjxEnjOPQeEjG1cIzBD4DYQgyS8FsNm9tdxUIxhSN3ZRZSNomKd0ne3lnXy
+KH+rJtqsBAM/DjxHzi9fDWjJLx5g2ih2kc/juQOWktRQhDtB9PThqenjlevtp0aOCrO7nFMWC2U
lrnEqaxPAFGK9kjDxXcGcarfwIwGFbdg2ENMfyKtlJay67gthL/YduXLtzNFlW77+WdxK/rvuHr9
HQUC6frj2El5VZMyPDD16WCW6uc0l/3ovMURblqnEt4J0pJClXPv/vfvltyvawgn8C/n8zvjU3hq
wNahyXa8hPK2IcokmalD5NklmwIR4RxRld68VbuTmhyDKOq9vrc+ZN4xkYyqM1Vo4eWxLpuXiFJS
oJscVa31EqudTsgR1RT0g87dprh9KCBlK7u3TJ/7Wpcn5EWjbJiNZxbp4AB+rfb35DU7eSB0CtAS
hTQ9ENIoRUhmjRbLgiqvAFkw+FSETlY5B0zE8oifEu5L+C+IzL19zdW0rMGnQycXw426FDvpe8FE
Z8GZeVlj73yDuyF4iujeOs538CBDe5alCxQ2k1hYrc2SvN/5g7TDMWxKWctt1zqEMZB1PPF1j1BE
ZVSBRJ3R37YJr+TVUiPjUzw0KbAqZLNgtql+aPk/mG1sfhLWSNPYlc3i+sVZdKUUbHdoNOLENCqv
AxMXRyO6IVDseYJbbyvip/sO/mFljrLLrrM0vK4FH979us8Y5gG2oo/0zEAMJYUsSEhRlroR7MD+
dhjieRTiZqkrGK33ZHTLlmiZ5o2dCd2cU2MvzE+dHPZMEeSaS35KRPSE9CPVc4Rh8tA90TZzWVxr
/0u9TfouK90xZ8ymHAJg1Zso9piBMJmdNIAqShdBNB51HbFDm6OnLfBA4dZkNyjwe4SZSRb5NrTP
GROlq1rtinzhdbagZoPQNMUN8ShKdfSRPXD0XdaZ8iHITgw5KTRlS+vO7r637OolcaVl7tWgTgQI
1Vs4V6EQqpd3Oc5Qo3yxw0QrP+VU0zygAuYmC1M6wAbh6csR3RABQ+rxaODnBokSND1fqt1B9V4D
oYRUeHferq+opeZs3s3wFpoOIZz+GdwVYh4sUw4sTOnx5CkCtT5XhPIpDaNXCCTqd/rrIPEC/VYz
CK+Zg1GJDREW5vmJgePkXm/gzGJojuCrkl8EUENsMvfPdQsqwDSRWLU7ZMeJFOOqCsESlC6TwYyA
rkBfHkfsWsno5zzjY0+mIVayQZWP3hV/A4g6XhxNhmwSnzwYFGRanPkicxXAQ6U8n/lB51AaTBTe
G5nmljBIazcb8ozKB+zz/LYcM7AAh7VIRTmZL3ODs4oK6Peg8NWhKUcwCELm1t1pUCR2JeHuVraO
zDeyCSorFA0FcjeJhO8VOgHR4dzdBY+x0FaqShO2xg8QK8/drcb+fUuZPeul3yGi/iW3SJM/Xffx
tyP662DczvN/oyyVUeL6MPhondy6AP+9ZAoWV7DrrL0B202eui1e8t6lZC5PwEk77veP+QJUaeZS
W0L2Atsqlpf0jDtNuZHZaPkmCdGg7YKGNa+CAQIrdvhcbY12iJX9s6kxoqHZhmRm5VjAQZr3KYr+
3BktN/a6XMevZ6TnY2dZezTWxoQFfm3Kv8lvH3leGRwnKU2Fk+ldDDnKQfh14G80wMVs1Wh8LCNK
MWq24lvDSYrSAWMHWEXlXbCpUv6uBnLnvjsFVkv930ZSnW1kdWO3iyQzBWp0xngczO5V6+31sN22
nZo6ZsUD6nCdjS9iK8ZcFbQ2+jymdL14ExZR/ys7Ycqz2HOXcrv4KtBMGq9/dN7fndoBa394c7Gp
DsqKUCxMA6gbddO9fo+vnL8MNDx/Av1c81F5an/mrZGc3GTa+sx4MvIOB3DejpD4CQ/CY3eXOdk5
LcET7k0tcpQYDuAAU0utxhp40Th1PZj0KeV8K0WDVi6eEWaN8AWskfSJ1rh2bS5v7ReNs0QsLujH
g40S9vQiOySZhK1/EvN7CQf9GUbE9CjKjOK5wd6AQdOhsup36Y+ngbHZSi3l4eZwLhQDygRsYOnU
fCXfS91GgjEMM9wEwKzJ/MAY/8fC35XVgwqzo0SW99EZyCwAF6cfbzJL9QuqyjDOEFcFJFbefm7n
ylOZ1XfgbmvH14nLJg0S6KEHdB4O/u54lnh+CqaDYRQm+62ksL9H/5OrgvD8Ejn3nyOSYAET3FLY
/tl51Rd/67ejkEaGG7bW5MsWkMsZC5Ue5M856VPCC87/BrF4ARbO7mj78OuTnSUFdMp/jH7D3JS3
OQoX94kPcZVM0bqFZUGLZZ1bM02lS+CicF+1PsEXVYaAtRH+j7Hw7f/1bio1x5f1QanptKh6uQts
UDwjip2QUxF1bqjXdjA8KyhvVRKyDUikUsKpU/BwpzuYDuYJOOYIFg+U3nY711qgbWc+AOMQoj8H
B6yjHpX+u9qUnv2iYekSCYQNrf/O574ubKlZizfgtrOrWWridCFSV7ogViojYn8J3rsiCYxRm44H
9HBZgU9O6No5dYNjwCbyQ0RVx//Xat5C8UIdwRh+E+rQBSRUnDsd0mWFb4db3U1P1ADYR3buH9wW
QFhsNwklUruBv82d1N1RTG3d+uh8oEuUU7NIXdMqROsk+TaQ5Hr0iCgfARcdon3ckud+4/kcGCoO
5BOK0V7Pr5Rpn0iiZCKnsupYVcRmRP4EtuVgZ76gsdD5XenlSxo1IyfsnwCZQzC9rQG91z6EKIr0
IhAQtaExExUxjylaMosfI2RsjSvkt7S0A3NbNbvt3LeyYkn0bfjXMv0c8kLwFMBikc0mz1kQF4++
6RXEYA6o42oOfiSyW3TvK7O9Wdcec4B1Dxs/Zr+pkQlfdqTbGPFTikp+UvcwNgPiMKO9CAXIrYi8
/eluYIpdEfyICzpbrmQ3/vSZVizZVMH6XHZSZR9PFHyELO6qY9bJdwYmHlsi9/NKFfQP/wW83gjx
o4YbZLEuodog4ytpYttWqDZNHmjUJEWk8d1HtLw+vDO9TsXvmJHrPNvnQtp3qPwVoSTw9JTek+Rm
/UmpOhAy5EIIoyXHELp4Fiewc+UCgpWQuzMC1Tip2tFN+wqReZWZkmTZhoiXYaS85j79DeGbxhce
EVUVl9PuoViJ2GTn5+v1xpcUcPK54uRNlfa7nRlYyb3OE71YBwotCxve2yJBrdOSPcDGzvW2uk9T
KB/NRUTlHVLHCcTzOtQQjaAWBypfLAiq8y4g2riYDVfU+eE0WICnnRdZCi6+Jz+/nt5QegDjUxiS
o6c1Zb+bqgvCbvzWB8J3qZkicqoSa1iUL52nfvEacUEyKSDQTQ2fKD99CtOrNsW2urJmxsashIYX
wHn8QQDqaJfD31P6WLmFEZEaQqi7SonCEcxgZIvZp6jwz+0j0Y1FEFJjfTocwb18BQl7ejA6GFsn
eOmBCKDIXctRV/4b0P+Q0S6EeuNw8G6hTxcSID0YR/hmcffRvPihIfRkQJBrJ34FE6ely55Tvkv7
t/nv/q+dAs3zuLYliYc3Gb5UwlccH1L3PZ7L1HtdBC18bYi0yxz7potTD/ChHyHc/ijAnZkgSR+b
7IyRAR3yVPFE4o0w+pMIr8TQfxca6k82Np95dAYb2DfOqVtFOTgM8bGVqXD/CWuIdPKJU4Fsobl5
RYBxTSbGmjegzLZuFj/N8bXXQEH+/OfMt0StK29Iy8sZ3lNZJKYaX2a4/iXJubjB9wYJzI7WyZVB
4thw/0lwjDSpJnijUo8zbrAq2h7ilk1sDaCam2UcjK9bCpjK5Rv+L017fZAIdpNHtEdwVgLeNUFX
j8r6rk+ZbDrcBtfJ7WVyZv8YeM7JObvRWQQf7YZdnVUtlPvdNbpT5lkfdfAHkqJqh92UgQVz+5mr
ew0e6gO6en7u0xWdlk+FTtlO5WuDZDSIorthquBIS0FpVCfeah0B1CjJ8bCdz5jwi3L4zqFrcox2
vH5tfAbhTWTcd7rAOfHyzAd6g+8Z/VGzFUySTwJ3rS4ZKD1Knr2klhblBuyQngaiwTN/cRIbe+OS
FAWa6WmFyqZxfsbR/Vqm+jT9Wh3CB2iUXtdcQbvGBwamIX58u9zauGI0qnCgkiD8xsB5SQhx9OOl
pFzwtR79E/YNs78KMSPPBy+jYL6As45HGDw95NuCYT/K8qFAetpedn2pKBiUslPVSzgPpuHLUpPh
lI2a7pDjgSirJkm+F9coHDrSQhUb3/Mba7f6gVpexyxkB/oldY/Vz8zmGIlDNCO0Z2NFOWPH8cqz
amguyrF/mDPD8+60p7DjJA6QrC2UDpysSpu3S7smjyc9Ned9kbgTGkRkdCEoGOK6mmKpc9GHv98/
EfICUYSTAmQsONNttojKd/QO+jVN0K8CAQGBxacmqAw5bSCCxu6dNOZjzo9Pcv8phXKjPuH0IhuV
lIBsTf/rA+ONF1uU3RfM8xDUGktaKo+3q3q60jxmAMKEHT5KC6T7XEmYYK1cAl0aka2BhG5SObm8
VoOI6qNVE3hSUXMOWJp6KOFOg0Qva1CF7Rnb8FzmKX/qttjeTxvA3VOhaouX4OKk9+86FrkBZYHe
JotlBlXFzqyTGIrv5C9RifmeXfhO2G+REmXLsn4mHyLo9FTsHxrhSCeXTAjVTH4NdO7iorfq0fC1
qh8BunZ7f8MDGePi3Z7jBiEWmaXFtfekCKwbrLrQ9kvIoGe1aGotTS6hrHFAKIjCoaDc0shqWHIU
dgM3QdPFTJydsqDy+oSABhQnT6TeSAeC3YvW129wBcmtmrV0ooFkuo16SITrauQ8lMsQPb8iVgn2
R4LlYekeCmhsXmb6Ngzl4REGCUr3HqCx3g/J+Vg291KNPPSZYQBBloplKXzGdI4X4I+Cy3ZG/4mU
cPo5QFuXRwNoFrq1VFkztH17cvYubkNzSOgI9a1OU4KYwZMiRjIit/QYhs0dyXFccoz1TzYb+XxZ
XnTEKbQ6r7WMGQdXs/7WEng91ubRbFa7/j+/MSspNMLi958WU7V/APMihhYQZLKQ2sMsp2xN/k02
r9KsSO7Rk4dib3Jv8i9pmmdvU5yLHvvBlBynQHJUDvUwAtrKTiy9mWR02g1PTkf3Up8qwdN3/y/u
fz5wYOqViCFXOu2cdm3aNGavt+jaxcCZca+MMQMwsApTWt3QqAAKEfhZiJme1J0C6Bj40SqP7cBD
b9FldXr1m44pqgw9BsUvV48vKskdzii/hUT0OKEbTCfRuqRp+xnxKq2jhyrroo5DhJzGzIUIZOcd
LjkRNw2vrUgCoZcHKW6V3mxE6Qiub1jMU8GY84I/c/0g6naEWDxB4VXy3I2YvGFsUG5BO0c0/L00
pyxJDAxfNIYBvNt9AATFD3PkYZEKFgg5PSwNraS2j6Q62mi+94nIgwYTpbcJPBMBTK99P2IUEJKR
CIuHRMnpGAKuTqYnitPV6wxTzUyv7ls+FshtvUFz0b4Fo4w1bkeQN890OwmYaH+clAhE5wvFLKub
jL/G7tYHVhQJ+66JYaMX0niF1DUAm4dXR3nvbqwA4HTOgxxOPn+v9hVpOelc+lP6xV7kF3DncQlY
ykCM6Ml7lwOCBj7t8RneFY+5aQseEZEmqkm/iS8310ClORUhCWk2eEDke53rmjvi7lasu+VgMevm
KiC6qFM1BHeSgP46nJb17/3F++ZaRs8bp4mdZ8sRyFuyETs2GvJbxaO9LL8kXY/gH3fOMsYAU9Kx
edIjMDNP6g8aC4TElTIWIKJ+psCJyzLeA3QY6fWVmEZeA7Zi/KnJMg6iEyFChl+EIhQyzJvPY54e
lntSLsTutihpM0h61CW7a9o89iYyaMl91JWW46t9pBSMOS5FXBkSaYqV+LjJY/RhLTWjriit9XwH
0+BrRia25HtVTFoaXmHqunhmTzI3TGGXZBFrx6459cyTc7zXx/52SyJCZqli7Ymkwg7bSWkpape2
bMMEOTD07CA3Rdr+MtIV9z7If3Rt/S984xe0IH+gkXI54oVb3/jN17b+N0Jrpp5wh1a59RcIiDJv
Qnu+q6O57HDGckwPjuqh3rtPx8Rt49JKmX+yA8kPjurrpJ+XCEoG4erqA7uCwC0LJw38VG5+Sagg
GhocU45P28q7TH6Rv9kx5c/p533eFb+/T5czOtpjyLezL5wmdEVX+f1rJ3V/zbAyE9RoGII7Ie0K
Sargq3Z1l/KEUTwpdZvdJsyj6aEhqUAzWHmB2jEL4mxwIQ0nL45kV9ZDwbk5y5Bieaqaaq8ox23r
rgUG9jCl4Jg657DxP4GRgwgNYD16ISb7WVcxIpxV6PksIMGNU633UCghkDrIKPcx090fDZvzBORp
DF5xwrC38NK0v3GTPglIDUrLxRWme4E0XEBVLf14iwLig5+Pt76y1fVseRefCdP068cAF/PYOuz3
z4247+AwomOf08bkRd35Z7IXeZQIUwY/jEsGUpRVbw+RL8Nm7XrYgWhjkFIO5bgVMjO/wWQrX4Vs
fP91mBE2j8tA7Y+OreILKNrlsma9mmGqiD0Yc7kW6VaiAm5FEXEnrwKNRH4ZAjGH5OhysNywQCTv
Fzl/xNIMMHYnaFA6Jl2/M7PBGqEhPSIrMT+ZaxZkkbN4hvU7Fbrt7IGdr3ZwJpZgIKvRVLY+/oL7
ik9mwf1GJbqnqBzUPTC9EA+C0Hp5TRBXclsn+mvELeEcxSybbIksp5LC4xrq9Ee5yCkZvjfrbrDX
T8tjqI/vk5X2PTJut4eH9yFiv/xVxWs6GIR+3OzhnslLJSGu0/Sv2ErBjHCOKUp6O8ULXbnu6h7o
M8yePRcjTciebjayazQX1743X1owP5cQhgg9rN3I3ir2T5UvuGNO6tr32LwWxs/+bPJcch0qAndM
qwtnPdpX3nb4iSHKfgYVinz6IuCGxPachDBw7tGVKRz5bjCfN08Ga/eQB9ITqimYhOFkbEMEvQ0I
EN/djMncYgB2moPVrVaKHDS1oDYf+MhJxAEszwY1fNd8VB8oKlB7IFKRvmuFx6lo4E8+ytl0fn9Y
EZQU4D7DTrXSbZuJmHWYdetNBDyk80hTu9uNCF/s8uQoH9vjHMGNCUOfUEEgMsP5sR3TER9GXx/6
FWhcI0vSOHuNAWLTDSb9SofTP8DgpcALNoQdGaDaojNQUVl7+SgVC7Tu2yHBmCtm/jYMbqnYdujT
K4+qIcYrV5PNqTNbbSdAxLf/nTQ/ClAa++8qHercB0eLt/LAiE+FQggZNGT6g6xEi2Yygtv7AgqM
rrHDCI0fhGrt6LzQ2mq5ZPusH7BHK70Wt7qd0GCmBm5acRh8rfL8IR59EmRMvZOCL0iuD8g0737D
urrY90nAF/5X8n5psBq5+nNdJeIajCULoauMsL8BlF8FoddknVxI1ql2PJlxY2fp3CO+i2/L89p8
SnxMIaMjVNxhyXl7aEdSP/9TQqQ6H3vpITOc58LLS2UJr9Q/auG4ZxQl0BdrzLzLxudS5EEzNNb2
2WLrvVjr7M1F5BmhXHCCuQsToyhFnolRDcU5+6j1Dleg1VDPJJUaHNS+TKTXrTqv9dihrCRhknad
ZWCpB2xoh6xHa+G0dIXa7QJrJJOGrbvdMmeV/JvZzu+Gwg2uyL+hUh5xMKX0SDMu+hAhoIWs0Sc+
RGfroxTjhKf5UVr6d7TczKD1lOiaK7oDw3XvC5f1FxUXrONoof166C8cai3ocb00cIpe+NFyHooN
L7omPiMhaCa0Ug9FWjeMEGGG5NdHENRdZIibwQ26c4eUHWRvo5h0Tv4uGAGRoFVjNqNw8u+OLFQl
K1ajyqUt3W1dnF3GkR0zwThCv4BDi9bRuqUNIclOinQ+avMVplnsua+sqBA4TIKPFNaaxGEKTNYn
15jcX5bX6bfDJfflz3x/RlkNAYYbqG+1rJInKo8fE6eO0/EI6gVM5ToLFXzSrp/Ijy22te8T4KHS
WSzmBjHMHvTQwY5urA53JpXRAibp66DbiT3Gqfvu6yH+bO66q8eDFAmPcFwDiPV1/3xCPfo5d9YE
7AbPv2PA4P9VQMyT3WAWGQLNDqzQ1cYhruzSa98iHyqW8LYInU6HFpUhmEWDvXAbfp2oil3BQkeV
COfZSf5s6ldYDnDJGfBenvB28CKCcIDgNRUp9xpRMagXBjZc7REoVKUf4Q6VopLbq3OpM4yQahFA
DXugkpJ+x0M65Ms1ATzycsYgUndki6Sac1u/XyjEWCb0NN1n16mcoWV+++CDfZ9tdvec65fF/jNd
/NaGkNPFDKKa7MGtAp933B6D7XC9Bta7/TUgnA3rJ5c1bgTFt9FjN20XUXs+easq1bdAYPqifu1h
qDGXtEF3snNC5N1yt3bDOfQOIBIpZikPhSjZHgb35b9OePBSaVp62hYfkfV7I4dzPo6+vt+3zhnq
kP2W7EhcfclO/proiy239h9zOJRElttkKqAefEu/ITq0kyaHzO496jXmwVbfZLq3nycbS7TG8+ND
5wj4I0MkFVkrSc6vlQdBIyUJEv9kBD7Xcj7zbKM9DdenDy3pScCPogevR9AWpYiyuE0NbbOK5wAu
MfWd0VilOwBo+gF0O3zo9ufyNmh/ACOho6UVfsi3XVh+omc27GtEw78vQTe05pKYHqJPcOEbmsEy
DZfE4aHHyEC8CqjllG617vjXIhqSUS8JuwFIpyqHpyb88EkRuRpEq7Ulu7qQd2Y1gD+aiRT98If/
rZCq/eXmNoyBFoHbxmBPbCyWMh2CDnTLg7ioMcjbp3yvenxmSt5j49oByl8GfDwVy7c+b8p6yYoh
kTo4gRwFNAJyLgnJEYSPDX9RyAKqGz5EC+w5B+xgj11DYl7hsmaxXV4Dvx8694O83aDxscroAPGz
CaqBqv8obKP86qcQvh5gX/I5nGnv7PY9oYenSQODxWFr73/8GTVyiexDBmNBDpyvEdqKu3Nfgf8C
KKE+YLG1ZfyZMT3desOQ6P01+62Wi2dk++f4rS07MMQeSJq+vRbnbIX3mI9WPUdMHJNKu2Ozzrbi
w4LGYYSJyYW20+L2O2WW36ZYVpIdy5M047hZ+VyY+3GPiXxx+62kYtaMfeyzZUXhc7To81HZZRcf
gRkNJRqhIVUI7rBl6l5VTQRNdOvi/STDYsTgTYnXXCSVFY5C19AtTF5ESdZMGli2MkgEhbz6FOuX
j7X/tmhVKqPC35ETy5FJIZCJX7IahQPVrwbApl9u86Q50AUJvfwEhpe7yZ1ysvVdci/Elon2xkWm
LrNZYCLdrR0Dg8mAZznCrswTtDrhpbCd16MS2MwmkgmD3buGpAYkGMHpCRjph+XL3ibO5xGp2kgs
miywO/fQXb/YZPOxfXe7DnblyLcnwHTsXAx95EW7EEH2VNoUQzsAtrhE7azNnEJHhRspl7OMSdLZ
Qubw9qK89WcoNNR1gHx2iS9YnjYUvDKnGsn3n+QemCucLgrX/LbH7/hPcTX/XeVTPvrWvoWD7tEy
rBIkpwlpYjLKEOk5YdZKXJxlkO+YywX1soI1iJTzh1IXYkHvAitYQ3zxVApFdRvBCaCO4j6lb3QS
dykJrA5Y0xlvYP//ZyI8vZ//xhczsdJGvg4Tl9qDX4FNBtAKGRsk/HICOG3/kk/60TQ4DtPGOoPD
cRvMlNh5ZJhqJtlr5DQExH3h1rI7+b/jgSna1nCvEwk3i+dpsu+D9PaD2XKKs/OShYeouEchxoRB
Gd0MNT5DhouX0JYrv6KiwInR/W5J+TsM0Hws49flxfphgu4MM6FnwMbscHo4Z0P3Gjz02Wahm5wL
ls1N2kg6jDPi5htdXEdz+HPlE4MFmhcoDlZgShkPKU8CXVzpXsUPmHrTRVmFg+vG0opdc0jorPQZ
6CQQGAWeBEl+YQoq9MshHTxcrmJmk5KM18vrnV7T2KevjN9Zq0U/SALUBGok1dFTtCQLxpSw922Y
3tzDQ1RsU9sPfYtI5zjb5J2zYMtfodnUa8r1Ar6We+Z7Ckw5YbV1qznrik+wsQcZ0tY8W1bR3oIH
2LJNxFclGuegF5f5C9gESnPK+n1BRK/AJLLfPlu186a9hAsVoOGM8Fv/1xJvVsqeQ3bNnm6ZTn8M
E8mYs4tEe2l7h65oismrPhaG3MmBGCNlm1kJneceiRph+lwIzzQhD8ihRXLzaqK3D9Y3wfNLzRAh
u37ukliiSunDtrXAexh+I/3BiIfeLr6P3ooGG4tPwcra9t+tTtzW890vFb7iREmx049gZgn6PlLM
xyONWLqi7MP38vFfVWr4Ozzqz790+d3y5ZaTFkCTHy0pWnoCjaaEzF9Hv4fVXl+L0YvCAhnb4Gqw
bgbcPUtK9IB4koH18EvEqEZF+J9JQWEgsYbtp9lLPlJkI19jmn9Ms5+IUTbA+xxW9aQWmqMBPQAN
s8niTSLzlQqdqaOALlZFG8893gQpTYbaPdKNJnG9q8YU/HGDl44e6vodPz2MscLB308trn+3RrBT
AqOngPKm2OPL/oFicbFmE6JrgcTCUARVd0WWBO+CPURJR98AdbZELMt5J7cqDTYMM4mhtMUUp8PG
kzmp+3AanQhxn/ZKDQy7Z0DuxnL0HdcvCouFqezWIdmWU5dnDJQAV/fyx5xwrFxgqn2QrQTm2XMx
hnF68jwol5JpvKZXwu9chC3Q9b/T9HO9Qq/+EHXIqODblXINSL3KzlIlIbJpr7qYj8q/HvfTuUzz
XWUuQJp9lniQzp8xU/g2k5t0h2dWjDY9dea7/866MbPCnH2b9aw/BKWpUEZ7AAErI/rKNBXaZVAb
u3ean/o6t3NOZxMGriBRg/mukWYln0jhWs6FpIERWn8JQf67vbKmhAGgn/yDKa89Txi98txlT1+d
qWF8AnSWQI0dnnQ/VQhLxaPJDI6OvpxuMqr7f9Zdlc29XHEAd88NWvogw7xa7Sp/QkPC6T+ZOAFm
mFZajVpWmYzQZUaLEmp1/mXtx4pRCV1gPWfMjsXJwop0HwUk40V4fxYU618RPBLp4MZe7+qagMOQ
HoD/h+NUTXTG+AIA2g3IYLbQGNfBcaegDkZhLsGoRS8f4cjf7Dpf+1Nd+/0dYA87SASA0ln2s2WH
dSCypK8PlpYSGv2/z3DZICmFHztWcOkdDlnC4RQRTPgo8OE4iZBn9Z6YhUDmCGtZiGCvvemu7XI6
gd/pzyOlOlZ9dtYcnLwiv3mDuRgF0bCH9O7p2mZfL/z4z/QPSGwYvEXk5BPkCXi9hlc9QzsR2rzQ
2PIQXg2IHR+yDqmGWT2fjez0TIJAa/5LBGZouCXW8qchn3afgtISu6S3kDYrIfsp29HIYM7TVWhc
OKW6R1XyQVG9COqIzayHxJROfH8/bGjxDyY0Mck3iJr7R5my3zi0f3/m0Y5GM4WOdM/Xtu7vSWzL
0AqOROciylYzG7wbCmWjaHv8xh0MOHrUw4KPiXeOBUrki6C2DfUvYb22jxhMu4iRrg6Th0NkljJI
bWZALFQd9tBtJVIrJ/EGThOsD8c8HjkuoSYMJxCeZmwguULT7dRNyvcO5iB1NyiGAk8e+ktXqsGS
zCd/RAfQnn43GC8UXUEI6jiw0bKEoM38uiRvLR+iJu1lLvNwaY5v0Nj40uJcrQsCyoJgxqimtauk
kBX6ivZENZVk0uUiQ+pJPLx6yz/bAJm+5SuYNE5DFBx6HgjkPDNG3efvNpKpBduj3VO7xQYQD1/j
8r36pF520X1/Ay6fORQmJ4qjaaARVUgY7piTOIU/YFVPtQGVa4JjkwdT5Rb5My4397+zvOZg7S0Q
u5vxXdvc9lRc8tD7rM9CuLA72Lm2fpAJjcZvfuYsZdYBQPWnwqr+NlhCpFVHz/Y7V6pRmjp6R3iu
Kc5XtYB2tt4+h3vTkOj4OP6+qk4AkLy0zMj+nMbJ4keE49SxTboqzH9FHIcGowUHKQWnrS7DDJsl
KJUaw+tdhzmeleovxszwnZ2Cr2p022EEC+194Bzy2xSE8YwHB8WCRePDMk9PYjubeMK7CK6+8p2J
2PGJ9bKLkQNym4OvctLp1gOOpG+f1f1wmSEqvlUPb1Y4pT4sPoqtjulXKI0/jMjyUvTNzoa3Dp63
3IsiwXuW+ngd9ql5CccL2gkL7Cv0ZVlGio/2Dk2gRHp4kgodn/o4CIfbowFIBPDAuADeJfhWmn6a
/59THjcUMlKzVLL/cfrBgqAWhEvhQqnHfi5nkilJAFft0r47PfMCIGji/GDmtP9PZ6Re5ThWVJPJ
moLaJWGtldFjV63njsYFbbyGT6oE1GkmZmNLUCnaSpjYJKuAYH+Mbr4WWCI27F79X5Q7PxGR0mqr
jfUQ0yFYNyAnnA4mCR76R8sJkh9jbyWhJS3A1k5Y7Tf1Zf6nZpPYyzSQ6VAAWkFD8gM2lY62A69q
jzlqAkQbsEEY7VbbPi1eall5GUvljapKR/B9V3DTxYCvIcTzxnj79Zlg4dDvO8yd2PIQWfVU3XtQ
UguC52IjoLsXCpMVMjBTkBOHcDS6ztGvx754rBXHJMeAyLL0VhbMvVKDo9h3kdob+tbFLDUaG/Cp
2eTNhYS3CsZKN3efWgHcj5vL+2WXGxKrr6IqT4H8TemvHiaJEnCnl7cL0uZd5mjIqac9oUBeYe04
injdCmlBCac280d/qXn5vkynMAgOMUOU6q0Cuul0/DgngM6dULmLbKWgquJ6z9tCGW+ErocZcTf3
F3jtih7m7iGJBIcfTDBB0YJSlfCeSkRQVG+rhK8bvEWCaBRObcAHE5BKhU8DW19Y678rD5nnst3R
0EcH2AzT4vJzjGlkAFAcm2nRG06McUYgKIK4bSOusbRMnIbAimqGKDOQfDp5n+B019ZWZ6qIqT37
tpaaoTgCl+C0WVmaDRFflgSrZN5xvI14r7DAV6kdm7yYhK9n1tdI3FdNo6AiBrvKgZ6YsjHOSeaX
F8FcURvLHrfzdjMNaf1hdZ5vzm/08b9yrEpEVsob94ZchQOaiU8FIGgR38N6jRH0qXFEZCUzHjGC
iTWnwmxMBjGID64RvdAdwFL2tw5u2YsolB1YCAY8Elea47tS8ajlXyonF/0tU56dHKxvLiw5ctWu
AC9TjQl9/h8N/QlFu592MOG3DneJE3/00cl7/mNG70RmfVDyJnDBGeQLrzafRS7MWJpf3pnVmw4e
mh6i4t9HCa+3w/vIjHK4UcWvkXq5p2BfJEGxPDQG+2lXoNbeLFtf6VMkT+xvrSfJx3+XPj/rYiE2
KM5K2U1L8Ch1OFU8prlpEGUTsRvIHYUfX2m+StZro1v51qrLh8ifAoTECgYCyWOdvwT7jnusZQdy
F3xrxrgzC0ZaER3AEy/b3EwvFWHDpAkp9Qh5JKEA1YIT7RA6E8S2YtaFlldsQNFeja59zTjWKQzS
WYO6MrWzRCtZou6wljlZyZ+ovGdzFYW6I5VE8y7C+US0lgo/8RubQbXZdRxlrBTnIfliWXJJbtce
QFpIIENt17YRRr+kNdDch4V4Osoxul/0bO96DeoPZYHnha6QHQHX9vGBVuY49mVWO9TiU7Ne0XQ9
MXolAActnwpsvIvM0CxUA1bdLUttHDQa4+ieHul96o0NkDUS5uEanYfPBK79MM++u6JbNe6b7vUm
e6ViTS+LkBPQpiycDMtAvWLpRBrVTJgrIdNakbsR/7MgP8HlobeOf5Mt6PGFzz/uy94j950yTPis
ziBsISJVtfn66WfVmLlu7sY2+lK/kK81MqcCLkoRXO/3FwXyu9c+J51bbrExGoHdgVV4I40PnQlq
PBeOr1P9XfZTgq5Mq4vdMVVid2ugDEM72nOa30iGWw3qkK2DdtYPXUa/OjQ8yGNDiZrd19ALkd9x
yvCOtbE33PrD6C82NU9/YWKiXOZkh4BIKCiY0M4DzsAU6vg190hjL4qwhli1Ulr3QdgSD+3rDup8
dz6fywL07tC8lAsVO86IqCu/bvFyE3TDCCg2o+LS9Mesg9DiCGUDRVItbSCayd2yNE4Zri+QY/86
/r4Lwkaj4vRdTSM7DbB4COfpQ+HO4cliy/C53Tw5JWLvHzxBUTARhCAB532iu/mQBWmNHPFy1N8/
bwYJlYTzDlXcCClFROjv/bCFqYpDiTPzFCBwCfBkuS63a2nb0jEITPkw2pz/YnZLnTccXzLxZCUA
dAYk8Bm+jxzkBf3N97nO6REhtYwH6p5dRkI4yt23An1oLpUb3DqBCbhwDf2wGadFPH2MBRkBtagM
ldFlgBOs5W19o4MsWuUFaiGWWLPKOxRSHC2TF0IgQpQiTdVJVgmCAy6HPru9nlf1l3QTfETpbR7m
wWUYP79WQJAkg9Lsefjd65UEI1Naj8X4xJkvY99IVUqGcz26S9t9BXIy3/O4sjNvXS7XAYNeSGAU
0C09+P+RGPhXTne08SsoG9LEFdcKpsW85ptXwTXBy73/j7EzSXqaVLyfApUMzSGm6JD8pOm3FeHa
yjPJ3EoGRmhC+oSfg9K1+JAnkbF668C3zmf6NqzgnyMvFkemTlYEAbBE8vSUufkftD+4T9jLm2Lf
OnVa+DvcjDWtu6dGTvKsCxb4N/7PxK5bST/r5lGcRGOltkIMzEj5W76VB/yZ8QbYy4Iv7TTI765R
uAvRFQBVObuh0PvScjrjQqoPIMrwJkSp35sD5D6S5dbUPBL6RWK6kYT/iUTvcbvPLCZeTLV9eLzf
U8acZCkHiHxmCMAUo6UKilkewC8d4ukURCCYnlgD4DdlrAi4hkgrFiUnRm5oWBk2xtd99qwi/RPf
hX2V6uD5VolqEcuZkdZlFQZRam9+5iJhqgxhRGULtitDniR/C8QwaPgWR0V+dYcNE97YYzxrGaHo
okG1jGlXcNEEJd1Ul6c3yLf41P/GzeEvOoIEuekiWmm2IabxxNSCAHdrTOnSu5n+fVAxuL2pRK7B
TMGkeVc9HH7QNhYyQaCRTMQLUgjSMSEX/k+DMzTksi1AWx4BIlgeQSZfvbqV8uoP34vzVaD2kFtU
0gUqrYqG2mqk+csyDSeInbXnnjCsp++wjhtzas4xnXxMy5afBFhvj4ykctPo+/UqdG82zH/Remg3
5nlKwkQbQBEDJOkLealCxCTUME0V5kUBCCPhZGd57qSHvEXBIKvHBCPzJ2ZcuK0aJ+MWB5raqp41
IMoqz4NiQKPkqIpMDGriFFgCfMGPXF263Z18+3e1l05jYqjiuAVduFSf35d5cBAaLBliLVoR8HhL
+NFM33p9v7L+NEiNzmwR9+SfB4WVlAcZDozomFX2bkmUolSk+LCAXgsBcsvgvuH3ETElpHehh527
q4ZlPFmsNFpr8jmHIM4G/SJ3BpcPgkkDcycYslbxWkshmu2iv0lwwFWFD79pWAMQzcMlkBOZo7so
45AHkhVwf12qRjhLf+UXLrurJzMJuhC+gjKQH/g2VvBjV+e103aMifPvlbEkfk4YeJwHd85kA4qR
AjsO1V0XOYCQ5lIQWm8eNFb+HxTPHNoqNOUZSnijjhKQD9/hoI+a3QKvc1Z5UCJrMIMSILUzQuic
uMTi8Rcq5ziQl2KRDPi6fFQK6KgZQBuU3k40KORFhfYpgzQLKJ/PXUJ39Rl48/7EGl+IpI+/Tx8n
Qc4o1VCcg11QnIFZDUzshvIoRWEwR5m8YyK1X8PC74JPZEbVU0ABBGbx1ftNyRomLr9TAT8WkN3u
niQS6qmIzPpkfEr6nAllro9kRkvsi4pIjydLCKG+o7SkQwrrvVJuufDuGYS8GnO4NtQxzs6exJhf
c43KVqT0FtNldEdZAOeOYTxv6UWC+jOCi39BXkFpDIuGE71Te0ptQ4TFsEbVE0oS8Re6F9nN697i
8Bxn4dXIz1hxieLtGEmL2rzolcohL0kTlU2wBSEobhlLZiElM4CZjpg9buFy1N5a/nhoF1dAmCjm
jG1Zd0BvwKaY9IRMXGLdZnmRBPiSk3S0qrFZgZmT8nQ8I5CmZf4vgVf4iIaXlQ91MNJUQERcq7TV
30lCytA6TKRN3msb9yAZUnHI5LaDs41cd5i2Wfq5sq9fYkZKPcHjdEgAqEedyOL50dVNi9F78tVW
xVObmTewtolEo1snZQWmg5eCjr+zRdHm4V5hI2EYRM/5EXEAClhFwOqcJqlbsUEOrbCTbS23XXtL
eNit5KId1iOAGjXjvOI9LJ9iOaHyBMXngyR/3HvFPpGJHRoqbknjgeWKZck/+puiojnocJQ+NqVg
oxQ3fPgTZy6S4hMSIFVrYsaJWwG2/ABHcqfDQ5yPXHoCCGAcPnrtYQ+IlPdmwu3T8aYr7/RZNF2V
5+p1j2y6BiDZSZa0iXFepr7W35zNMuwGKanPYIsJEOm9DTLhvzFl3s9KYDPSXcaA1CSGVcsPS7zl
UZX+1HpqOeKnvaaLcGXEJNf8tr68Ahbm/c4ZTOSwEO1zg4CWBUcSg/tkC4mwG3d8gLkEVopfMrWZ
ffl5XCjmxY1zo3PK2BNc57wBe3g+fZZF3UoX+64pfIG+S6iQ4Y0wjWg2dmKk31BdvXlkQGdw49UI
LeM5R5PVF/JmE+1h75wFEOz+3niVeOn8rfA4xuhqbrRy8M6MOxf4WjH8XfcS/5n6lfmAvUlJAQzh
hZdajFKkKBfOgzNngJYVi48yeRHQFgPIge57/FFmBkMp5H5+pwwhFAMiXnMHGMUZOMj8VHuho3RQ
jrqyCf/GBMf1cOPXQTiYMEFnufo6c4zbgX4144ohpiBYiyYChqfYGyM4JGwydmLUMaDnHJXBdwCb
hKPsAAntswdIsa3jvnNR1AS6cdL0dx6Xf1oJdGOx44UiiIjcymXzD2y0JS3CHv4v1z+hE/TXXjx5
112QTo/LwEZgkRz+3a4MwXvA9Vgl7HmH+opXiYrtAv4YvefhMWs40CyZ5NpHgLpAKeloS2YbmG13
TkqNuX0v22btRUR3n41mnwDmCOv7ZuZevvI7qcSRTxcIlvxCu7goHI3+DbR/aQUyy5047qHY1g5x
wTYNKFIbCD+xMR/AzyKJZ/3lepip3AYUNNpyDV4Sv/t21fsNPhQ/mnHK99y3qZ3EjU7OusCvhcXG
PkiZCkXZZSCdzKmQvmahWfSqVdsYGFH+GhuKIzSC4xUv6cDlOY9tMyvFrcobAYAYZ4q4Lpe7FLJn
T4NkpmKDE8RyYX+e+9uteMPGKHqSXJVyZy0JZQ7cDMPGoZ8AOOyjm1vCXxXpUtyfB702mflcB+Tl
CsfaOGNX0bWSj+SoDOW1R2TaJi8yvqiC8OYW2eemxpuVNHqolqbVw4o/cbeaG+rDrtARyLnQ68Yn
pI/I32amK+5NmYRYsXA23nv3rV66oHKnDy1dHye6fG5+6aBdkEv5usBXAoGyo3Dyr753pgE2Sc4x
T1pbt+h4imJTLX/n1VdMLn8TgUxPUExsibYMX5fPiynv2Ww02zHYjYj8EkXOgM/XJfdXSNfVo0w2
PzbF7SUy4qMBysnCnoLRqY7e9SW/SMeCB2z5K+2+GyoYIv1DROHM6aPbGslqpB57KsWmvtomPJWF
LDnTULN7+eNxt4ZS51qkVI14kaVokt9EfmAs/Z2NQTxGnk6T3jr3WSoStaGv0on6Q1gCffK1SlXK
rWifM/vpG8Pdlp9bFzRmWgAPoEM79qmrWn3RRSVOcZ8G8RwmZGbvLSfbWVGKvt6ZthOb3VTC+6Dt
hFh5y3ksnsoQfTx3kbrLhqOXGPlbdaycAIinwSCPuQukvK8WLhQ7SpIVEL8jf3WcGE8ClnkwIoun
/hVKua0Ruuu9ZqtiPRfGpQWy9xJ2NNJkiYLDLWfISOXP4HfhWiI1EZqlzaDIuBrmQY6iQBvKQDme
cBUaql+N0V5R8A0JhjTsHRShNZjboK2e1g/nLEFQWMKubCyOf6c1FA+46QejSV1rLsPmjIcQ6Isw
UOU3AlglZQiaotNnnIH9L2Mcs3vgsBb+GeFnCVO7xhEao4nHCxgV7Y2I3tWUPuNLsuvFQfs/ee5+
HyPptAp7e33mKHwjpZDr27C77uUl8CYMHmTtlzdIQBcHIlu0+jrpXCDOlDb0gFdB5AAyCal40VmC
aQ7mhygzm36cpVVkLdMMnOf06loq2punyykTu48yo+PPi1FUkpzzf4Dt63Bj65z75TB8qu232On7
TrfpLae/akr08syhJcaJaGsMuVW6h8/w1DGLpiqFlOPkjva+Pq0dIa0X58cddJAskSmE+hgODd1G
AiaGRyglFYhEoNhflcAxdrUrZOvyrs3HPQ1Z2g60AADrv9llTXn0LWOomlb9oUcPzSH+9M0sJxfZ
HUMvSsA+HIp0Dy8dpaanXL/uWtSDcbUk5a+XyPfI7SZSMoZBK3HkilNIah8Ht6jz6iYYeXPbYetJ
zBcIwzGOqKReyiREUcibDS4OURQEyXbGDb9aQ4ThG/8fyZhMv+7e17HrC/GlrqGl3IJ8Ow2ovYeN
ffB61N0zITpBGTAV5H1TGECF54eyrFDZ+9wic4rJJTmBIisRiQK3EM5WZRYHgTfrogGbgI+3AW7B
mwlV0ec3n68vr9Z2+0mxd0Le0EskgTc+oaosnyJSZUCxE+cZaQrsNygBdMggnHFAl4/Vm+ipg2sO
joJxFhdUltdSRo9AHevIP1Mmr7MQ+wu1r104K4Esx007kCx3pR2LBhd/SjYYWR2PnPv8meRg/Onc
k88hP+w5c49WbJE1xJgMYBKwVIxJxJXEoYdDebOZvVQ3pJsNW+WwZH30KynwjlQoQTseImwohkox
gpbqL76cPyk9VVvTNh7OzXkRJ35PnsWBS4D6SlqQW3KlMzaYbDvKw+QXt6TWNKvNcQJCUKX+jAF3
dHxdQ8TcBlXLK9N3AWyNVqZQra1MCtD53575r1IPBtrSO1Nf1Ea0nDK1JyEtX79firsi3cVS1MxN
qthapWwwBcYwgJIP5u40qoLHL0e5oLclz1Uf0x+dSmNaPw5zIHg2jxxaeTMDkaLiU3D7iCVfotsW
1TCD4CjEdr/heeGG+gO2+mnvi6vkYASiWazOsfQO/AibQj5+mlGwgEC6FJvjHgl7rv5egRyI7CXJ
OiDwi4Nn7784f5+F/v2jXMwqbbxa/OEIuqb9nKASKpGdeZU6+eqmzW1S4WcsC7+QHkVLhV69izZC
RjKDFKZ4SFpW7xMiyRBag20nd8XSofPxITD8+Z6u2h/7vF8szdVDAAgSJckpFPquj45CWgcRZZbg
CZF+LKmSWFIaH61SP4vv6+RHyJLzcZVswSPKXZuRPEQKTbqTT/2QVi84fSi6uDCns4mHsysfV6VB
RuCWDcK5FkVdmxSB2+iEtfR3FxaDMI8fZ869hNKAJ0fAr+VuTyCX9dlJQXPAUQg+jnlno6C3Ee4T
ZsnzpqQlPw3dMB67qjl6B/2ge0wswcdEoKSNYHEFg7a64gfvN5B6/+lRMonuJTBJOtn32C4kuCUo
K6RiUpns1g/DXqH9fR9i5REgAeeTmReM4mBeg2ev2SSt1B+crTtF8F5AftKFc9LhUdmF9Txqy9SC
FgwScjnDKaLuhtoZYPpGwbuCrIP8jdO3lRZiSlrZnfuaEOzgiZZsIGJPo13C642YbHE7T5U5nNZB
ixFjNPipCJj1fqqmAy35eJD8zY/pJZYzxWGbIoekbraQhkCvg/tE/ZSWz0rj3okTjLUCPYRQHNKk
Rb4yz+wkIeAnYTFTjOvj0kC3ulSQdEh+Wx6YQqji24JpKfJMVHg3CSbj4Jyly97QN+UauDf/Q8D+
uFBIgXfWkcUIs0nfpMQJ0ZaygEIIrEnl9aW4heiImnszd7ewsPCF70Ca2qHe/1aZ1bCmAmskxTH+
sm4rsABNwj2PbbLM8zCMFbxhfHvQt75rZ9vbB+iVq2ESjlCbFO7Sf6aO9huJoTKjlumoLvhybxwy
gmU0YE4iW0OaBLQl+RHNQTZ9vbi0qGZhMD8lCyJEVD1tsFJ2iVFkYyM7rdmj3rG7CUgj5TEnuYoo
QtfIaUDNfy7kPWHlQ47uOJb+wT9Pt2/8vb/5u90KX8JPcnJmKpH3gAiLz1qLk1QDaoO+YmrIBSmC
0DEvoDXcmJkTItzP285FOQR6jRY2TgxvZx/7/o13R42FolDP3weBeo49p5SZoyuavaaYYMZfxnvY
dbGzthSAwvbFvvbybb1zOH9T6UOPBE97f9Nto09nAdcOba3kVtdCz12box2RAF19xw4sjLc1unBx
TSw0x99n7gw3p4dNF/XyMPEapmraVbRZHFKs/JDs+PKvpEEe2VI1pz9Oyn6yh5VSh2FsMIHMexuz
kR5+QLmvYOEOdWprmQHOsNuj450xknjSQsnqVJXEF6UpWVScQSF9g9EBeMWL9HKMhHfw6+hWgqiT
LfpvgGxLV/aXqZhZgkX5NAKsJxQz5XZesb0ZZ73vNb232FMSfMlOSe8E41JbnJEM6ANdfJuCErj4
m4pN6/fsUC5aL059leAjsncSJNDRu/N/oiRGeyquONPzrRFM8Ci85m82G67s79T7aEdKO4pOcd8E
00J276uSP1gi5A0fXfwdFWTYNG3uxZQFNcrqQgIhHOQ2gFvNY7MwEHbNDOCz8Hr/WkALxD/YsAcS
+O27Oc5NlrNcEVdFCMbVjG5N3HE4BjQAwRgcKaBB+ysrS60abKVM92CPArsdRO2IQlMKaYcVxmwB
aT4gtx7wRA7LNh/CLXprZRM+DAGxiwaZ4ZQgVR04zJLXNnC3XM+lDNzxDXqWi0GccYsl1A2YzPqJ
+CCMReeDXS+gLTxoI7YgkgwM0OUdmTjKD49MuA8jKzbgcCZ13W5RXa6LguDjY+MyiW/1snTuxs7R
sq/KfV/fJUKjtwLfS6b9i6FTW7aKgCYLdISazUZkJNB2GSoqUmpduYGpqv06E45zF4bqquilS3E/
aOO19jBFIklRJKQrILn1wIzFhuYfmrioYRVU3etTEHKYP5UBKKeV88/HBGs4lx29RM7O7ysnMp8c
yHrMk5jpLeqVO9Mrh9zmZBRxQGUQDO7vhAJqTomzyKkRsQICWFHkm1pqlnUidDA6mGRIoHbt9/Fo
J75az7BAC9OiE065lAnv3KDLi0Yq6QHFRi++gLg67FEHR415fizOe89mdCuV4D6BVh4wFLF6wdum
K8d7tM2Kd3rCQKfNAPzu6CXcgDEbp7aPQincPeuns2JkhekqEQYXMiEkkfwrNse6Rh8hdZ35ZCR+
1Gl1J7oOZg/iYsmjWbyul5rfLjEoZASHd8qpNWsOFaos+LoSVAjrWhroJaJV08N+OcMbB1Sof/fC
XFjVZBF/hH+xOJElAaMUCpNvJ4teLtkXBXCQQm5Uwscs6Zi+LqJ951oBE1/1ke8FNvwg8W0wv9sl
6+JWUsLyctuZEuNww448VYKJ76VV0Tf3t9qNlcyppo7VtNhERMPzAOpdRB1CPT3yKPZvuGjII2oT
NZDQYPcy6haygzzCp3qAr2CYTccesW50qQFo3glYDbFqxgqLN0VBxEDQLo3Ah7uzoEJC7NYnKKzI
NVtxwqMOpNFzFy/0j2YKc+wsUWkQQKZEUYQaNBKFQc8+rLYZCyGqG/tjWkm8mf1SeHcHeHMRPvnw
Ld5ZbyQA3wNVv0cQt1ka+P2+7swjwrcgq48Nm77YbPEc6plNhfIF6HZQXeg9f35lc7oPZfJTqnVL
T4KQRgLX7dsGJ07xs42MD+beezs5iJtPmRnKlMeATpfPGW+dq2mIaz5kLgXxP/gzfBawSJc5uJ9v
Ic2me4z4JUYddOqoYQC/aaFXT3nSHddzhgMPOnUw4YQ07ALXpJeFiv1itJlBuRLciIjpZIPV9csJ
skjPMIjJ73yByTZpqSQxYagJc8LPM9QMmmqhdHimPkLblSO+PwgdtIeKVCTyPpaotUA8VzW0Znly
N8biKdSyE/vfyELaTDo+ygzSJwQdZ2aiZhl+bn0+BjszZcQtTRHh58rN+MlK+Yr7RA8xCaT6LAes
nE8Yxao3TL6wmYvY/glAynIUEQGQoVKKkMcFbbM5bzjsXfKd1ijLnzGWRZa13DMS+BWQzdHm0m6u
nCGjcUb2tJR+yQ9VgRosuns3vHFDyl+qAAWAcTpFAlUYta4cRinbdiA8QoQiO0avciNDqmECM4Za
12jDbEC2c1jupeC0DV1MylhVk4Nc052c/2tlpu4Qy2CYGxilhMjdA3S9A13lpnIe+54Z47IjLwwO
LtQzctn1W7EubFu5XU06xVeGDwMNuenxRR/5xwi23ThZf1JhyDDHK/r4GeAfTxwY7uSNyTKRwYV0
F2jQ5nsWBHGXsaOfnpB+II1xKDvO5b3wU9u9ks7t5PO7X+WiUvA1uJ9MLfKR5MW3kqQMXsCZdPKE
8a6sNE5x3L70ZBsbxkTO9xI1RNQwP5dPM1IwMzjcDzt3ovnB2aGWWUGh9cN9XrBff3T/eTcA+taR
79IbG313xw3g3Fbea2DF9bOQt0S8jWYwpfVT3wcqj391NAMYnV8ibwfDvC6W2WF65MSE6ZUhu44k
8A7eAez7AAz+iaoz8TwqLaSXpdT57Jnih6U7VA9cQzRtyE+PPRKehrd3jW503SOw3hHxDew5sOCx
7byg+bBUtJ6oKR1BHADhizwJc1zNOShownVnOUrL3kPIoSiq8VFrz48vmfYYD3d+f3kDCVqr1wQO
r6ITFsShJNvC0qjqdGhj0F9RT5l/w4dcephPYR68S84Lqz9529lmneaPvYrwQZaogdmJP4V4lCOE
JvtcX+xTEm/tGg5h9SHgeCp0XUOkpk84Qyw395+q71BlN2QHh6Y+y+zB6bEsFde0jpqdONIUrQbo
R1TpWwJr/u1YSP+/KSDMW6FWjj9+1SuMob49Uw/EojGho/0JFJ1tDDQ5xMpIfbXoBC2oMlJFEPQr
CdbMG0xlmaQ4X5abmD2l3R3ETzyEW0pAvwb2jPgPn38kLTe3iEmfpazcHn3qRviIA99mjTDkLKxY
zJZdogMQA28wOwknLymXpgqyfcClmjMmcZ+qeUEOIFpbne3ZMOdi8wYjBfKarTuI1QKRfbfLWUJs
L98j00xdUkZqaitpaTDysenym1DVq0a9uk6PeA/2YuOel+Tl14jST3GC/WUZo0PHIzyPcp7cLx7N
Lie06X9fwi6WFbPR5L5/jJPoUuwpQibziNLPhKfxcEdYRFV2p/eK9FD/ElZJnS41ZVkAjLQ0Tx1h
1QgvldmvnAcwD259R8W8r4pgb/83mEyZL4j+U92pPeZHw6Mb7Rpv+wb/qfAG3HEqlSO2dMKPzN6p
NW8ZNbLUTvIjDiS01+rsgmB32MfWDkS7dw9DX8BNxxSzPzl3fURRpka4DdZpWtClRJU8qemo0EJO
8hx/vW5iWV6sCiaVxzj6H19a/hqlYGalgmRfw7kO+evFQQKOKdaTG3MY+9mH02Kp18omoozP3yvt
RxCcdZsrhKqkzWpOnhtIxYflcUOZpmB4uv3ypWq3ejXNw/nPQUCjsa9qsFT0wagIFhLTR8Ko40D1
1ywU/mTIAkQlVEGBXCES3m4SoBsW4Qqw8u6QSL5shTg4RSpkLyWYQPeSayCc71XsD+Nr8kIFUhuB
Q6xYDKI0VRz+8cgT+ZVm9P2KaH6LnZLZDkB4bmyUDBU0T+gu3wcOmkMXeF2fgh1ivygxQyL4orp3
ZFY1hRbcXNUygf4wUWkPHb+JwH36JUrSsWBjaT3De+a5akOdZlfcfN+/FVI1baR7je1hTWnuq0pw
Qie1IJqllMw6P4xf+hupseOh6ui8xDzxmj+3zXpcMATR205f1KZ5MvA26L70wJ5KhM0XKTTglaOo
P3VZT7mo4g8/Jlj5AmQN9ENIHuj6FpdO1sCMxEi4c9g8oY/lBmrmslHTaUYupvwfLL9wejxxODrt
SrCPKKbvahy4z+2GDlKP7v8pQIS6a+/Bu5oxjXo6M8akNtGgYaufxFhYWN6HL/OuBPHK19ySXYoj
Dce+7N5vdwTsMcY7WY1ab7ywlFq/eYamEzClbQCii3h64I2XS36dRYN7CLFVGsr8iZA4StpnY3W6
DErT5/sOg+EniyOFa5KvBSsupiU57lY9r76jUYPEx7/YfQR4CbPcEAVVebpwQyHqz9FpYQlU/kvE
vWuGDt2sgw6PDOOllydddg8tl8DA2O5wDChH1PowGLig2o5Z9zADRSip0zSfvmwD9omBiBhOrMWH
p58ini0JpMp/UDGzKL1MqSH1AVElMU2zJJle3m5hopcV3lx0izu4kscZiueqHX9KGaQrjvp5NuIM
w99tXQD2iZhM07L7d19JRlmkK1WgNzE3NHkRuTOc+rT2Y6AXxLzLTd7at6gf22KtltAkgClIewDQ
xhRyGS7miwEWNWQ8LSFARzMStsyFCMffi0NLwCCoLPXZ/JqmGbcA/7a8YoSj8XI1+phM4w2w4fd9
JJtiwjD0io80LQXoEOPBm4LPZJ1Ix7tAvivvt4TJQ73fvIO08zL/mC/sEYsliy66Y9c3fDGJDltT
+yg7IYS7wwL/SN5pjhhBIy/quyTV7DZD8vlT4wrtFPTnCJ3dib46qELFk7QnKBLw7OrfN9IwrfnN
T6xi/TNWlqosu/GCIuSFigMBsjzwuuBh3dP1Ic3NFPhcAIrKZimobGszB5LLojQoax1W2kwIiQ/S
021gGKI8il5Hj9XRhqMEsnx2sopJbUL/JSbKMua/HBh97AOTM5duzokqILrTPkQneg2QUsJVSzyE
JBERVofgKfCRf67Mgtuu+Uelbk94uXtG/6sSj9x/l3jzfWzeaTRUcyegOxMVtaAmEY9KZvbudL5A
U+DQmdbqV4A57tuqPIA3ffTrjzCLE5Jlkc/fGrs5bnD/LifLmN8E0I/Zu8Q1QNrP07zKeFZnfbw+
lrMA+I0sXMWq3zj9sZnNjCZOnxfwKTTNQl8902boEif6p++pV6aDqOrtm2Z2VWdrFvqSdjn5IYgY
ilVXMQ0d1t8ix4AJa7sU6EDe6a06FRdXKiJTKpGNHyY03BKp5lY+64lrxfz0/TEV5Y1WGT1jEByg
+EmhUmoaNtdbC4N1FsNOH/Vd70ReXffJg7RS1DgPN7f9iNIW+Ovcla1itj6qZd+066BrKFcXDpNp
Tf3VcJ2YuNWd09xZWZsifAg9usetMzEFz3RReI0xgKv0Fr+e7O1AlHUu5aFqqLwLQdvVnR9qKucA
wdbzc4GarKnqq26Ly8/QrEwpSPj5Se7/d5BzR0WCzhFi+ZfyAMRKCM4KZW+4Nl13R4MbcN/4IkG5
Be6yPRw2uzMtMdzK3B9byIXrFGQHvrwRG6mCXFJ3Iht+vbfe+9ezC+mG/YhpK/5S3S+/FfJRHNvh
9pQigy0vu0E95PFlhQhP9RWaIgwULe6f95/p0DO7B2doUtX5Ggu60/CHBuQKdO0sA3kDGaRp29nG
uhL3oIusMIiy4UgvPF0n0/5CFBDuiWApyc0Uqgb2JjqqGX8eWsTu/jIErWCADaD4fsxdZKtj2Pik
DNGe8/fg3Hwe8EiYXDDmjtPnpkmajvCYE0islR8pzK//s6RfQ1r9ty7pOXoAZYXezX88yY9r9nZC
GG7WxmoK7jwH1Jgo7GvszkMxnm/IH6IDft+g5N5hdOdhkZLm878ZC/H/BN93Thqc5ZVCrqLIYpLs
XhMgj/KZr0bLowvZ0b3ooFgkYUFmwdWF1zuL3N8OG2XSrYghrW+qPPBA1SiaYBlRU5we3vhZtkXP
Fto8pQ1872zN1KsWX72maR6/aYhIS2f4AJ1q9Zg/Fdy/jEYg7LMjimo68H9uZqsMuUQ7p9n9B1UQ
rew77Fd8it9Br5KICb/sqdg6NRoorIMc8HYqwkP4dkHSnd/fTmxJ4FlS2/HWrPGsQpHNuL39Rq2b
GQ+Og8JCkwXNZybrIf1GScCA58qagwp/2egr8rK7xUHlksSxUv4Spb0VgJs4uJTo5I7OanXruD64
SHIrZluZ61hn1926PDec9wf0KqaSNhMBeuBsfO790HcQn/R2u1DDCGMKXWoPHA6N94Up7CBs5KO0
d04Plk4fIHLevhH6fEOK/jJaeYHoOSoLWdqyig+sw0dUAy10UyMCv5gZfmN2D+H1jVuJkVyO+fU9
ng922pn0aGJDfrXxu/G1hTzR7vXRKqrEiCPF+kut0+Ku2h7w+vgQxrCD95pw5fJvmnbFrQJd/Ruy
SfZY3iSNlefOhNoqj48DUw5E96MUnQx2RUoV+bAYVDNQZzBqzusETYju16D7Hlx3jRDuMSs9j8H1
GS2YQn/RIZYaHBXIB7KkQrPInXnGlLKwTZpK/dUZIUmb4gz6C4egzWWvC7XiWvaivStRLA207/EY
A2ZdwsYNAo5N4RycSue99FDxjayNc1zQujs1siTvBCYD3d6vkZr3UGWJKQS/Smow6dUlNBZvo+EC
lshjY5WuIWkDRmxsVits4qxdPBRHwOt9+qlPOcVJY0IWnuCnp1YLaINxxWYcdoxqyam1czU7aoZc
LxC71FWluyFR5nHrWWrP1DbLMMImElYvpcTZO47d3esY9K72GnzZktRXGJKDPIoBfbNUSPVTDIU2
78Q79xDdGreJ1W2UyKca6ekeNZ0fiKGIAv1ylD88HI+Rw1xQsVD3PHhIzGAhnLOH+w5IkbNgVacF
scloPO4m4BqWokJN0uX6y9js64BRkYmSzpvMr4Xlq7zpSJ6MSvv5k/JdJGokLLSp2RSxX27mYUy7
dTRG808AaKJLV5mRyxaKAhsDpG/quJRgLaYgiH0RDgEbjbVeRlUltd4J00o4iN7q6pMDzyzNOOet
G/bQdgFM6gZl3O6rCB/vlSeGUzQxZLka8nvN3eeqVUVYbqOFqy/0R78VTRAGSNHBcoOsuu4ejYZ3
d0lvPrWiK6nv9s9/Rz2YaAZIOj2a6rFXGi0roRw7mNls08JbxkD7ougFha1/dCjYVvbEitkPamNv
7+8xupFiRmPxTi2RGG/xILa8wNwlN5MGeMRdwGVHxaqB4ocU1FT3Yjv3rX9ooRs4O7mADXH+0goG
Bb6Y6JGySYYWADMbzlns4IgV9W0ELNjEutMuTl9iV/8CRxzaxW/uP0GrubQ2SBr1roIglT9/KdSC
FR46MBucpTaRAybAQK46FdTvKF0fcca4mr3yKNQF0oEnRK0/5qUfAzCWfAi2Dh22KM8uUYwLBZAT
5cu4unapJ+oq5PT7OHs+mS7PZ2U56B92AhflqfXPyc4g0xdwMiCi+fsyY+cFYowhDuj7GgLbtbkg
GYA7qgls59udrf19esOE3Qd9vMBhWiB06QyJI+/Pq+KkUydqn2XiliF92gWJwqEQ8ouLgPBT+o+x
eBW6uu6+1Dpe8nnpLPoM9juasRfGupS2tgIBpNTh6IfVJdED3q2dVbxhafGxv5RoVjwW6fXpvr7E
5anMxscT3nVfmH/uQ5AbodNepZVpt0xjnVVztX7wOl3bY8Q4hgVlVZYiTZoBWexTzrmGQUe6cCek
5mfu1Irml4cO9AnP/oTSntE8mQxONz8kosQNraqVkaf0IBjjyvRcWAavJiyl3xjaJOAZl1Yff5el
6/0VujpVhdvFtqkyNutG++46ZYIZcFWWRArt7B6FatZxS7HaCJjKc925d4YMSgF2REGLlTz0aQSX
J3mHKg1xFbU7WIOBuV2dF4I6Hxf6ZzH8ygYiWWhl7Lo623M/lE8LkPZugnjJ2aTeTlJkX3o61jwA
CRgfs2IEXkgdSqSOFxsoW3I8BGI3uD4tCZpHkiT4aji32nbsaLufKZTn2Yoi3hjJuCNVXZ/zX6J9
8DRCEyezkf64IyWfxewOsRUaYdfSF0L6iU9LF0UeGUTJpqYaltThM8UjeIPQCoXJmymCQyGBiude
6rQfrxhgrJ3d/lz/38NGTIYHiPx23PQTmCZ26NZ/0s3gM12ZtCfjMe7tBFJ57KY8HF+vHzazRWoe
lNb9aU8Ew61IO+ejsaR4X9QfOhVmvJ3paQG3UQ8reViX0ReODX+B1yW38txtVx9L716NdPT1QD0n
1OkJEGUG4ukQKuTtcal1qLhxzSAdZI7A1/P8uWESe6WEic30uZw7X+zEylAZUbccPrWStcc8EI46
Y9NTpYHw12mVm4g8W4ek/BJj5i5wJLXHnK06zYIfNOI4GkAjS1pI0mjm+I44eiK6W/cjApM8QI6n
55jPFjHLSi+QHXj6DzUCZyT/gMI4PHTB7ewLIiG/Y5uYkjrfeUeNoYcoAsbDdPyaCQ3tPXF+kCyi
fWy8a4/dgfalKnzbvHjKBbrg3xt3KD9HHl4RvxbXLW9IgxzpqXfwNBk0xJRJ9/KIZBxjFIek1J1T
7BYVvW9A5VbtmgIVuoFvG7UHI+Nd2pH+KNnqDTjYAZfBOM25Xh3IWqKilv4pmKEcAVkp7wKg30GQ
tiHHG3YmSsYpAhqmN1MB7NmoZoxcam3/YYat+SNxInX2zJ5eDp1/AlTK3gkSFuX5o0WnsSp4rG5I
gvXF7Al7SQPzNPCh2BDsxs0rRmpermyjbSUeVK2Uf74XR3U7tUq1MXqYmUo+gT6RCT/VLNAF0ITb
OvCK8aFRcDkTomFYcLZxG36H+30N+ul66a6Z6Ef814ERq/PxNUwYeJI5V3QFE05XzDR+gULKpNLU
wth2ARX3Sby5DoWlk40dglF1Za0xam2vp9otndEMs4P2dJA7wHVFhJNnNJMO8ydh3rXr/Zq/TuTp
AAwPETb/n4PhgTsqDzzCbG9l0g/+QMgIlRliClT39labnEQmPLsSzFR6hDlHwZu0rByqAeD2wdYG
7caMlpVNsaNKsvxy3f9m6XIILh6fjAdg/enKh0DLuOTTRH6lbEpx580FIUyzmDMb1s0U+PIrKtYU
VJlbFhcE+CjLBQFUmz14Zr6s07C/JkCLEl8fRgVFMXHBO7/3OVkm31u/CuMafZ3WyrLaF6XBHCot
gxzYh1DxfF1m90mPobIajjcCOhDBx0XeMolc5JliOxpmb+z8v+Qq8Wfdz3ytluPjys4sGXihWtBe
m7URgmfoUXulx8jzsCuZTJKOJhk/VW8BPx4kBwj4sWnfCs8VlzTGlVhmmVLEcnK3et3uSrjHZem1
WGvkWM996PyFesdvFotJ9/CLAnNrMYZKSn2amEbdbemmgfadTNBHwNY3yXBDHynFkoI0ju7iooUS
1USJ9/KCRt5ATNtr9BG9MIwyunKgFPvo6WGMG5pMVcdDCtGIh3a+Q7lQSb+Gu37N788PuQlq140X
VgrkwUa5z36WSGkLnaZTlGbiZ4UMkzDpmMEv7GRqxNN29CmUPwpLBy3oX90sXc+yluHUaMyM3RKp
ajh/lNdNJMAz8BDNpNtE0iQug2v2myYoeDdL44SkHjBocqcP1GA0m4AG8G34pTffO9IwRF7Z/CDr
15JCjbS8/w391se4hbqBiWpsTRfyK9yywdMQ6f/y1qW6aG1UFeppuYn3uOpRX/BRWcYm+QJYPBeC
Vkolkao1HUQovLpGe//+FnTqk10j3J10yNUnDzL+lKgcEWGD2fAxX4Ye052bljETQK4ZmjVl84Mg
raNpzJGfdi0me6TEXeZCVP0sFQw+0NZTNwBHqwOAKquenDSWW1vFWq/SNdSQYEo1vc6sw8Hukjcc
x8P5iiTPW8CTBfyzs6mFnKoUNiapxsQ/o8Za07eUpsrOyCDMTkmbm3T1u/BvmH76qXNlN6/ENvna
DyNIZwPDCPY95jlQbvDhfvc1LKaYTMtH+dYNm6UAIIoOUBN/uk37Tr3LlXMjlkAUmtw56HhP32xN
g08j0JOwnPJlkM1FH0tLEBykr2jrecMXtMgqPWcchHwIOd4K5qhNYdJkrMdfc4yxEbpQx4aT/axd
P/x8MvACDdhwd79VuhrAHB0GbabtRVXh8RvSH5B1fhyPnBEvLiY7lavERtUapgixvAQ0tbK+KWjI
qqbR32a5q0lBDoZBZHRYO7zDlEDte9Ep9I4TQ3AwQ8sutrmtxMFeEg88QnuPhwoTRZTs9oZxZzvO
G+e0r38wiE/O7HgtDXM4LqGviBzUI7mhLSAaWn7er3pqmoWxOvFYpZoMDu2j6uAWs4v1JZMTOIH4
/+LdRKTG9vIYTHO4/fINNWkmutL8YY3P2QEwFSFyjd5YajZovcDEvG19q2R8yIaXnyQ1rD3r3j/+
qyx5zfhfNI2p0jjQAp0g7j6VxcWwFOX0wP6ZWrUe0TZE5UiHD2nOZO1MFaqPRptTa6vH4W0yCYO1
7LjblEuCLXjpNRpfr2sQbUrr+QXl1rz6HoM33h7AQ+Qx+8Ar122YG1+myz/ROHeVpEe2DSdLUeo/
3+VpnbBhmf2oUiw+LifEw4wism8P5BlmC318xF2tyGEodY5B1taYgeEigjPDSOURY3gjtADh8DaZ
9lNmWKXDQmRdnL17tlSmq1f+VXuG/ZC3UipRBu9p9FcF3TwvZlYOEQ0+DsyiL1b083c7KgGGrNGn
5xfrwN1TzZ5CwR5vD23mEOYcpD1uH0bm0VbgWyDAGldsaXa79uR+I/t7qpvq8aLNYHToeMXc+BBZ
OeYmdeCPAT6y0XzntyymJCz0/7vTPTDL/9F5Yf751ZYY2Ya4WmBYKVBSRYutq/i0mjaPm6HklRG+
MTVm8eTGKXLcriR68hEzQe/4hDC6LByPTynGJ/rnV7/esSEntNcsAVwgqiDyGG5EGb49HxkWQLIy
H1NWv86Ebbb8nHpgl787HB8OOwz1flP+e1u8shy0H4NTKk4KMd2V+ir7am1i3mAfPRb8RwiZkIeD
VUDVY1m5rUke7lfJ0yZeBGOe35zwONGwu30EcFE17R62EuR56JYSre5bQbaFkaSHUeh8XndeQUik
IHILjqlKKiWpxiHtOoQUIiGcWewVr1fFe4VunwIRtJWUILPJIFN6lCH4L7uPIri7ySJz/W/MnDLz
534w88sBuIz3wCOonFGSLdJMq3g625m8SqzIOD3izCW2+R+tAgcX0Jn6YfUb7I/6gBHx0mYuSN+4
4T763ogcYmxnTbg6I3DdWu60zyRg/tzb80Qg2wxSkAXt0QMQfSzf1JXSI4Eo+AOk0zh07EHV2GjQ
f5k2BfdkvAhFyN7nLwBUAuRCLMU0gOzbk7Iu00yYi3viFnMxImR0CQGL428PMy58zGAtD12mfqmt
kOkNpb42HzdqgNowYwiaQ3tGwLnZXSwrmiC55KcF1+d+CZGIneBfvG5WKd8EWCnss2rZq5cAeK9M
a6AYEOatQLjJq4O2g3KiXqPlmt0BjDY2qUBn8WTOHwS2EjhmKS1NjC2UEWTITPotImS2GyPg4i0Y
XBFxayjdAQMzYU6iLO0NrXENIV7mixU/VEczjxI8s40Y1Frhtbter4G+WaxZ3u5fV7yQrYOq2oCt
XQnMZSIB207zhwsJoGSk9ecDwfsbqcMiWxC4KkEen3/NosNu6aRaDbulojFeu9+a1dfner/GSEuJ
syJxfmvU/8Xws4spDE2Ans7Oe7HLtAQTOHdc9G/sDvHbI93p+jV6zi+Q3Md92FzCOWzKuTR62b0L
qLrNHCIvjMoJfK1Ke/SLiFK0FMTh2eKyxQNzUmbdK09CyziiAqK/YVL7dFjSBfa6UIhYuQk/SCsp
hkrB+KjynZesb7RMF9Zc6gtVJEvvvwdEgxE3FhUK3RARGjwGiPy0TFXpLx9+GpwohtBy7vCMDF/E
8TQgvv+oXnNLjxc7K1feBURmaWrzHM2awgohCNwfGEKejuIftYfANlgUKDGE3D2CQbW0hbaCnYvL
+s2eN85q5xgujs0z7TU8i2UxudNUXcDZW8E3KflgoOztd+/hUrKn+z6k6PPmri7yJlaJTSFkcb06
9ok8Rzc4hJfwCEFz3vOQbw5OlE+PppUPB6dq3fl9z1L9D44R9Pp+BZe1Nn1Dp2W5nV2S7cIe7c5C
Yb2XwpogMNk73URqgrc/5CS9VHPprWkliDjgbTj201cZQMQaF93n7YJZPHNXWK8xOWnBZkdjlf9p
IdYQoGGVBw6sYKMMomI3h57i5o40WaQqKBDhBi3idL99SK/bfoODrS/VonXwFmbQHdXp1EGS+/xM
dmBdJbAJtCXv8GZIxjc6/uEVxF8GmV3ttw/5NTvZ30SYLgMPvbVz3OuwiPW8KNMQzjIxjZIIZ4RU
f00ce7pSlzonO5WmGo4Uoby9tm5rSSVK0RutwKbZqKzlFkHHPSstNvk7Q3A+sxerFdCmq1S0S4Rm
f6/conxfDDHtGyongNjhbnJJwG3Qept9g4Uelayp7jJjCTUK1Vya5K3zwcmhzrLOgggaPKgqtZtu
DOVVBI96Kpqy718UDAK1T/ZNbBCQn9jFfTBXGvlD4K1YFHAEkNKu6r+Ob7iuTURMe7JXIryFTWSL
HE34H6T9n81Qrm3/czDh3Iv2dspcJQLh8RQadi5qMqsrMuqw6x5w00bknxAyIvalTjorE5o2yU06
LjNeGcm1LP1km9sdJE7y5yjsBNG/5smQfDQXukGWIZODmn9DXpsqF51rh1ZEtYG5q7jUw7kZVekh
lc+Zb1ycE6QuS74gxkjl1yIdpzOYTHHamhZHlURPTu7qV+fKWeL6WiU87BqPzlHgUsje8ztJreLl
IjYtkycgLASsFi3cwwLb4A8BPBUYbtK32cwvjToxifNB00CHCSDyowJvWE1GMJBoKTqybVpgQhz0
9gKvuOCUiqj+Ofjr+CqzGVKDXyiJXbf8RAlYMVDXSwmtDzrt8+rDASuY/bxk4SIC+kod6fJb2hYw
f9I8e6nVojf1bnnjGEwot/QLRpcK1o0Q9vGfxAErAi+9+YwQYj5BxVdyQLhL7AmqyMYqFi44ZQsz
m2DagYgcObCHVwNYCu6X3k/QtB95SXpYnr+Co/D6O28lRAQY4/uuurlgzl6LjZTLrjvK8idfk4C0
ZOEJdzQgHEr2exbwuXpUEmvIu7M81BkYRHH12Sjoxrzuc1QF7yHMXdI15saulh1QxS3ZOv9mk3Sb
mbe8iFRsYYBmLqhSHEmWawY08Vx+tgv35XWTDkaWaRjIjhp+ZUnMTdafvYWm8sB+qeiF7MFk6nVX
jGoVU6YoJN3cJTG0woBo3DgnOhuUJNY3CW6nlOYJpG2FFpn72NH0IMy32nsVN3v03GuG9oqcjdW2
NyMugJAem23I+hG3Dy9esDh1zHJpxY0hll557ucF+wPkp1LZUH6oFEFP3UKFsI/tFNNGgj1wXEWg
ji0zv/pY/zMp+7fjpXvaN4vdFJycOAgP0dAfDrDi6QiYJ+GfZWlO1qnNhqh2ZRlUOfp38ju8dDib
tyhLl2LDI5IZV5ui8VkItFiuImGRAQO4pmwl9U7R5YySuAM05jc0xhPnhPVxhjbXKVYWyabuESAR
Cu2YIlDzuG61PLcRnwnNYUl5ob8GhV0yfygIJDN32CyCa+JvGGaeay1VDCO6tstXE/YcVDemYbbA
xQg9jBQMeYbFbdBbMoXKjRJ2hXuD8HsT55lo2jU9ikplSk3rNaFh9rVHIGx7kIGsEJGIBhx54ATt
2kjyiHYzxK1Y83ILJk/g/LJvUoFnsNQijcMblkOqecR2zGlQCfT0V6mU/fJYf5EaJ8Vi3qolZRNK
IBMYxXfbyvfI7pbfkychIe8i8lhbvBlPLjua688t6q2jiABjeLKHCWxamSezBuBB2tIvmCTjoJOj
MhlboCnOW4osLoX1byg2FyIAE94/pTLqqHPim3a1W29xDG+0Rn5pPiMsPM0327cr1mdBuFTBqqDo
iqpaJUZ/2jCBrOw8e2Bo5kdEhppzT7V8zdhGultuR3Vg4pryjWMvmjI3lAiL2AeFnSe7Qm9Xzyj4
kAxdu2IKV0t+94aoKEZia/Gljy7E+Nb7w75YfCk1GMqrvPvEOeJw515R7HuLukOVDE0FjhBPwQin
U2Es3enDfXkFOHY0CeO4HmGfwFHepbmrElgN4aMfx6lb/+ntdA0ABX+AINop5FG/hpXkbt91dXHj
FH7+TWwKNDxyPyYS6xNe5AGsRsBygaQ1QP+x0JNJUAA1aPUTEHcZ5ZhhULajFe1Z+3CeM/524zkg
Tx2w2g3WYNRTaMlYMkunb5WacVvks5wxM/b4UcB7cqTUHG+qPa9/syyVC65BNclJAsYuuoQcVLl0
wvU42db6HOxOoBvJcyZvKxvT4G6MKtsFqLAInmGQXszKFZm5UthMTq9Jv8viRWpdav7E+XaCran2
fq+PK7L84yly4p8Sk2+MTPP9DVW11p81G65Hg9Ee6DA7ZAUL1P71wGYqUyvNYf9scAm5/qjHLafQ
KTHR9DWNkEZWiR1f8WxTJkGUJ9MO2wA54G9Nl5miCPyhXCMKijMg5miwguBdvopYH0NE+bCIhORd
Ijb4nseWgrXeYaa4EWrwbFVLhSxpzATPF5RqUWIgWI/gdVb4M57dH8fuBPE9tGepPb+up1quzpuR
6VvJitWtXZl2ziEwjA82OppUgGykSKzZMGUfGJ+IzoNhxc8NN6zFcUil8qh+mqtpzWhAKVmJA6rt
yCW/dhajc0GlWXNBGeV0cSuJrXfSneuPCYodh40zvBMOUP7j/RhIHPvAF+QNLgabPkQSBiaL8rOF
fINJbylGSzk18QwKt29firQSF5iXYz67jdCH30ROilR4k9BI+VDOvBl/459sJYnUuFmkNQtKJIBn
ZlHCxKB9H4VGJ0nsuQJilNb9ZYMMpjeKO/9o7CA8puvujpGi7Xx1x8+Q+tTQ+Aykv1y9JsywEfYC
ctuHykFs60xbiYyPpnb86Enphh6B8tviqtdcXYFl1kO9/zK4NC034q0/muIRJ+4xnYHkK9SrukD5
zmf/QT83pP8MM9WkjrFsZ6xOv0kOGu+FhxaN1kca3zfRsH6H7rUzPaF+rlGUOWFZyKkMkopA281j
H21nSaaxEGzWI5L6TfA4FfuFEhEhN0ktmueyO9MpVCqIytKFMh0xrKpI80YRU6aTTEQd4X92Iw/G
T1Xyj+EEsAUGc/RD6siKmx6PTP7oJCWANJDqS25VbfPrwT8KfrWfdL9hssWzE2tSDOAL7JRWMRGm
a9MLuYXCZOXy8mckie8CoOYqduTNDa5nAROtqqt9iQUSSul+5zU27Q+wfl7kpkElgZ+4UC/uBU6g
6xfTb/1Kys/Rg3dOXNZTmMPYh8fLR8SLLVN4B1m3uwZsRmZO6EzSiq98iWGkc37zHI9ZNUppOpQk
Bvbuga2EC0zykelmq6wSxAp30oP6thJKVSHYoGLX8+6nmB2JBcdqel7d34xcTaY7LDZ4RjjYIHLp
0J5uY5c6rrZkAz6QqEEo0SSvmik+7BWilhEPijD1uTN0qjciRhPJ8Nf0cCROpFqbChmlG1CCOnxO
VHBldxFTBZQfrXpCEWOt0pYSxEZmVukhz4wIVB/ffKW7oE6vKEXogmvCP51OalKJN9zlpafjC++x
HfDl5M7QfMevX5xo1sbNFxEzroz0S21YoFblj/miqmByLQ/Pr5/7MeZRv3BBnek3kVlvR+zCjZmD
FuaS5gDWlY2Cq7ArW/dZD3mX9agRSHmMbcpR/0jL7/Kq+i8qBW/m80q5/XasHS5g4j407sYag+EZ
tGEiTFG1mPnuoNxWjYqFZLeNB+k9KbV9bZ9Zj0lgdB/uk23dHjDvU+6gAD1CDuqzyM/K84uNs6P4
cWv7Zmag8rHtrefE+wez4SVA4x5+u1KvR3lbIIRZt5LIryv30rZIUVYyIYaZdINyZWPFRfu58eu9
VMeBUl+MEadole2OlA+6DYw2lO8tr7P9idHT6xT04hTxH1S7a6maZmuTOY63wLsaB9FrWNfc9n7T
rU/jKZw9EEBeWZVKpf5kI5/2F8klrKrZXe0HY0l5Knxh42jpG35a9eOJkSJYn4zfiZSi1915gdYW
iHtcxG8+zwuS31LHacByWaDhaG8rdxxjE5Qq0KhdKgGBkC/n2ZvbSf9p/5gTFryhriLFzG8o7qdy
nu5jVrru3fX3O6hMjUCBLg1qGRukSA8xVw1xzkViCtHc2N6Q66GfGV48HotkqIIMr7eo6hCwSZ9W
I5sWTOKIM6IJn4WNjO2yksmtCJym6r80nwomNbWjic5BifnrTAzu8AvsBiAHYXtU6H6WqiIbUjTW
AwhlX7TMTTXVWhvKLcjAG6RWh2LwyFIHfVic5ktlsNMqnv9QC2bM69ggBh8TcyIcLdQluvqfLgO/
oWrAf37NP8HwORI+2WiDUqnIL0l1pfUfgRWoyVGhwZusolqL237GPbZnh2h6K5YiNpYvnC0bSltJ
Ay9tnvg2dw/ey+q3OfYYCSui7w74aWMIxEZqMYIoogL0OKmN9UPZX9eG6cYL/GtFpuxYuzoqgptq
tPO6GGrG/uTc3UbgnjqK/NHyqkS6d0t2eqgFoDwkkGJihrxntXuF9dz2K8tKm6ybj8/BmzxJrUZs
UUr7Qlpz+Q6VaZgXffaJvoZu5xEODbKBv+nDRHlX+Bjp0Cg7Q7hPTBNdYyv9GVCiVEmii0moWx8e
4SYv1VX280/sjh45omqzgzf2Z9GpvNyWQumh95pt2grsVHSvZfT89ROlBBEyAg+A4/PRVbnO6Jei
u5CFTEYb0+P7x01sD4JjgHNy7GNvvXnfje0H0rLScJE859axr4p71Lzf7Fuh9ZEVuruiput8TuwB
1xOHi3imjTc1IbMZWrBILGn7PZoeUWhhmyn9CKCzTNB2al+HU+dVSgO7aD/ncHNOYH/A1u8cXCMx
t4v4yjk3sitSxVVXE6vlN8CWHWsY5KI9tr0GDN4YbLqFCLMCQZaTNaVVxRUdgFR0OOIw2bbJ+2bQ
//4xP+w+OLe/TEvBs/EZxUwPZNPRPTT8DAzf9BnkbP+xZnhsBwUaz4J1PumnvD6IiyYRupptuD/J
wCF3ufqJ64TgIQ6klExwHKcifZlBFmz1mkp2OFVhKxAhpehSdbicA5WxI8ftwul8Nqppqa4k9TC7
8xjCYMd20Q0iAX0AN17XwnNc/85fXMKLHCI6zSeYvujqiFwzq9WSSz3X6GjKjW7JoE8xV0X/wggV
zQ0fzza1RleqjUJnWWrNR+2bHowRhHnP8vpgFrNSYojjXkh10IMj9nTfAeMYydk6xfYlDUclF4X5
UBJj0cgUHA4rbdmdYKqpCiNEiwRso4nwbxgIs/v7wHFxkk45URPlDvJiWkRzGyn9LwoKKe8tw/qo
9YGyXx5kriDreC7Z2QbP8mLIgfg3OLg6CveXvRcYzuHdiM1dBEqyBn7qFunmdah+Xd52eBN6+i4w
c58KVsWX+0Km1Xk5SewshsD4uLt+Bgw5YcHFre7yfCD1Y4+5yJK/PbNUlTinySwJRS85uSlQHY3C
8WVjI0z648QvjS7cMa1KosYuwjgEn4ppxIMwWiRRBpYUuEbTANiI02DkyQ02lJ/Wr7Qo4h2uvAHA
98nmJqXC+BlgNbzoW4pPQLp36uP/KKQH8JKgPug+TqZedhh5YYZKE1aH4S4kAdQCuuArFBBPTXQ7
0zjrgubxrKCW+cglcuKH+n1SE0ZGN4yVb66r9A21erjga0vtB/mCPQDyoH+vaIPcNWSCRgV8y22V
+vGyk8ZooFr66NZAsB2ld5p+z13jUDpMTBkEDCdByrafO0d6el6bOitU/Q9GMr2QVK1wuoRNDOrT
4Tv5t3Ga1Z7Wo2UiwHZ+l1Ycmt07ho5ZoKQXyv1N914k1clrFznH2SA7VSL9b3BjXH8+htJhjQ8P
C+J1HtG7FQhkIZOrVA6hoMtosQ/jAdCBK5ZTWvWuiX1mKM734N3BU++Lugx0sQk3UtipI53hLjhk
v03AGEXGDyGgT1bTbN+WLMTG73h1kX1mfKB3FI03Uyva/jq+5YAws9IjCUFYhoTS5vXSvnTCcCsV
4WzpDxO0J66tfoHgCPyGbeJD7wlo8D0Q/oPUvW6YVR5fcihCQGiRJ2QydS9E4nr6IU+YKT2Xtk59
wGNyb+hCEzNlP7+88dxe3Sp+LlUc+C2TBnzcTXhnLVz4QB1/QsXkNzzyBkBgu+VEYiJ9o5GVy2b0
ukIOS2yZPeQN/gBDwOoQyAuvbXl+lp5PFWlsp/FVs+QNF9qy1LAcCUGSe6Og32mtZhOAXC4xt83B
A/sPpbAbcwrLQoIrBnvAMLhrMjx1UHLHuM4SR/vjhfifLGC+1JGid1f3BhNUz2rNVGG3tF/HU5XW
fsYcge6jksHDSKNKfuD/1WocP1SXRFKbNZgvWD73ZOH6xSHC1ZAwhsq4Tk3MSKzZWX3ygNOkQyRr
Wxs9GeNOGe1IAXqtijYC8VZPzzoXYRWAeJy65N0ZqDq7IYGo7F+IHKYXnxsK84Q9idZqiIF+vGXP
jF7CgoxffbDbJwvsCdBRyZHQ34lEtJ4pwN6awWBs+5/s5bmQoQEj2mZrIVMEXKEDexqfIS1EiZKR
BnMirYuPmqfFcEWJ/xQEKWwAO4S4lquElhF12moTwsVYJZ01NY1aTFiYSflThCyanibqEac83Y0S
SWezMycY45iOgtZtfOX7CFPJJlzEKhbNBzX7tbAj3wvjvF2ZsRUyr7hj5w99ALIaluTKibhxIlX3
WgJRIYdqnQ9DQWRt/fdlHcY1dZ1HP/seQpsTfjpLIbuiYYqnT/gG7BudJpJhzER+Udg+iOKFOK7b
3NLLb8CfhqJqomYxovZOCWyQoZtHxaspA2KIecpqmt2OMDfZXEgnIwaImbrLLZ9XbNsMxGcsBWIK
MbQI6NNs+wiClo7wLqI42kJ+AzuLiV3iGxaT/qLMHd/AtcYshxQ16s1ekXRR8BPmRk5SAtVF0LaW
Z1NQnyyLGyrlyzSGBlq5FALIoZdRjJeDf/RQFDn06r9fRs46EaQbWJ5jrWrMZTbMUXv2PC5pFE3C
ZB6llgSYCs6gaMI62Sct1ZtjqPn/2zYizPBhBokno82EnFoQuHzXKxjQTaQO1zEOM4/XdJzuWmCJ
mVSHOvOgTo7b4AmCdIQxdCiZXtiRuSeOqU4/JFTal6ruuGVRT75bMLYONj3r5xY20TWyLx57ptpk
CCsXQXiLrZif98IUTYAOSFAaN/64ptG0RPB0f30EX4X2HpDFZwNpni5Wlh4bwng19Rpx2XL2ykvS
nuFdi9BeisYlr9Sp5+P2rXklCcu6mX4RRDz3hG+qwhahP/SAuhtKejEe9iXMUHgGRUpLykBtTeZ2
jDaSKE9MTNhBgtsfm2JjA2fUEwb1Hh5lOYTFdalSXNQoemRoy4Lxxa7C+uP8LzjhK5dhwW8m14c2
sce7gCaNtonHoT9wdcbR8NpYqtl2Veh8NnoK7ZlpSH99shb7f/ChfX/XokDdgHfRhMf8lJsXFt6c
RQx7CfoJPYX5ZfEhKlmQfA9y+oHKXNGa+UEe6ozikNCzF4o/YH41occI16vyVB+uKapX64ULBPQf
TrKRv6OSU5nUSo+dE5P8Nsx0mARhVcZWvwfDSUxc+dfqwC0KJxLfEKW7rAA0/J0l77ore2XnaxBJ
kULmsvCErkipX1dnxyvRGQGQzF+xUANUqezDBHMoJ7PW9n0Lghnq+GLjlAULw5d7hWir6IjEDHhz
Z0SQabKe9ZF64MUUJC1bbeNaLsGpiMnm234mDlJ21YVUwWp0GLjg0ZQIcv1NpPFhVfX35VkfvHp1
nX8D2bGu+3aTzCvbZh3d2qhw73mbIYt/0Qabfp7fjVN+qbjSmPE9bp+PbmF0xDUaWejLt/xaVPtd
kt1C9diuNQlEX/cdIhtI3GgsuG7n6vIWvtVJSNNCYsYo6qsM4GjESjSP5TOPAWPh/GTIFaCbMqrq
+Njq+pomVEiKeBIWZSlbm5wTWp1WDhvP5tSuD9sXghQPuAaRmfbLxXgf13cf/WcjvkPdzCOzcdx3
d30x3McQZGfvqR2GkASFV76OMBxlBlO0tVEvc3slvVWXCqLjVg+V1G074884zR0DztvWBV74tmpT
aRvBVQE2GJk3LPlZXqqIXKvlzNcadTOJxBitSVMQYvgpbNjU+RWY0PHtLR/c3TsLFFDHqf4s3JpH
xV9mZ58Ape+b5xn2IoN22u765EOS4BIP+RhT2ve1QbYIco/cPDVCk+cNpHzBtt/fzZt9G9FtSZ3x
S9NqMCq4yfQ3hvxdKFYGMXzAY/U5k3jeKG7rnFnm9nqRXT23UryRKfdR6cT6BErXgWXPrYKV2m1Z
0LQxd0ZBYog68Pmi5h01rn8jua/oLlpjIivNtV8GwNkPcYpZ9TFrSc8nt1ZSc/yS/OMNYK4liqIc
Ieu/68mx0fcjYVNbjZ2VkAjj2o/INIpZ5dBtcoDl5UkMZWCbqawHs6vkEyk2UTiwrN55ghvZyYW6
vhTDIg05Co04LKFTt0z88PJMwjU/avI+zsx2chzn323aB7QLJGhL/+84EWhsFsBI8d9z4GnGdKTb
ais7FQsTUsEWrsj/jvhg2qjpmyO5l/39BVRv37GJLpNDuU4twFavBqqJYp0i9zy+oZd9JQkPuPNx
ehwjZrgzBJ5FMgCrXaVSz1iFQGFODH/S8/dAHqXpNpzcbIZ9T1S8ANFMqcjjwUZwTciVNkW/djbn
The0hWsR2KdM9iCrobZFWiXMzuKGvV8ZfIij3s9W3xT3DTwmNFggpIxP4x0sLGQ7SgNLnZR5Jx4r
c+oViNY2YXZMSRqe+BvWJK1ZLkTQPdWs9ObwNr/28XIPGhHIZUcztCOQ3kP+On2SjxM4rb3Tn/8/
uw6+3Ec3E9Mi3q7S4prVKy6FQl3M4qcOsP+Hp08va4KgOw5p7Zc1HcRkmhkVfA9mK0R7vpSplkWf
4859umeI8t+S/I1DwfOo/xNlSowvMzfEnD/XyHn46ZdEvLE/fo9mZ9J1yZ8Prt/AeE5jcA9puQdC
pHICc0gKhDkrCxY0veCz0HPIFlxq2SIBaVa0zSSx9pUi1y0yZopHaUA1dzcPUQgf+NQZl6B/Dxkm
SlmNL0tBvXd5Ncbieq74EWD3MLNmsZ2CG2DdlCPgv6q441OWEPnySBYIO5v6cQ55cGXlWA3IXB0D
d6BsHAYoMb0JsVkVwwTYunjgJesvcRPGpHQe3evzwQBOvJwZIwqtPSy8TmMa4QxYLS0O0PK0nyuo
zXTwNKKkGutjTGTeGJGjGTALlFThJnn4111OwyhRZQOIdyKieQmKR13AZIebFZUJP7J+6eXramYr
1MjUJp1MMhG234AcEiFO/2Is12Kpj23DXPWcp7Ej3QFkvF4iHGaDruGniCu2Z9av6rEt/Ub2bSzH
yvDQycHevokicCzTGWc/T5tiXDaP9KXPKX3mu7Mqh4jCC506/nE+Ln6jd5zACbYWe+YRAcOeB26t
bRLFXj7XB383CNLjCPlFwIU+mqKu3zcusVhQIHyBE6qvtiveZ+TjJa4v3eomotjnANdmHNsRFjOG
SsIkYt2H4UehSNa/EB9BMJBheTokG10rdf2oKP9QREUWOhrZNQvkpF9jFPlkLx02735cfwvKDc+7
xe5Nug6H3wiKCt7kPyLB23rFg/eZR0VkHaXbD1bCZVWREegXyK2UJkqiZtRBS1xcqdBP0RzsVF0y
N8sI8tpPA0kqemj+IJ294LnS0SPEmDZo3UnJo+3dTWf2B8tAxd3Cbm7SEpEEMYt4xZXHTw9LaTPz
5iskIm2/qnHZY4dkAd9D1geXpt8ZDg3E+Jx+RK1UfgL5zBxqJgv8QrSNKGam7TdQnjj/C4povdT2
IC5enjF1qXaCl4+R37kGYjlpLMsBkTYyP3Pcy4kvFPLyZyd8G19ksDvTnRr3+vabTBu3y+E/Z8oH
qJm9NY6zSscE1PkBKMUi3SuGW35AiflRgU/MdVaz0yZVuIxKIE9KY83NrSO16GW4XAYmJFwVVnNE
cBsdLZFhqMZEoGuiVEovPfknYyQ6WNL4mMt+9cD3XZ3lUoyzPjALNoJMUNTwqlJnR3wvi1IrRAy9
VcT3DTljUVEMMdI3m8z4dLkvMxZF7mZkeTfpJlIhLQIw4XSYN4h20A3QvTBoRJP9rKlaFx747JZL
fCeg+uKKR7sRAaXtwIlcSj+YCP7VH7v+JL+FBj+0tqt79UAxGJMg211CKvRHKkU5YzZvmYXYXBaL
gb8U5admtRsjb3Og6jxXZdhOARm5HFKf9POlCkohOp4yrF0Oe8Nh91UjZL1GFRr7F1lgUtb4vHiM
ACZtzgo5fdzeT9TC1VliPBO/RNwtny0zdLLy0xBo91wkEXkgSUvuciRzKHiZZHN8y57cpby66JrZ
ZwivLvwgKiC5Gmgo5q+Mbm7j5JdVNC4/O8di/MpzQZoMfvnMLB5yEQtLtbFcPiwO4eCMO8lb2iLy
ky42nzIlMrOyU+CEHXQuKXySGS4Q0OM48/zGIbp+ETH8h53W2kOcysC7pQuiA1b/AHZT6ucnsAK6
sNlxCLIRC1J3Dl2BI7Ls67qfKmy3aJZHC4cRaRTTIYqFB6r7ybezdP6rlBOFcHiSU0JYyoKz+BYb
YFb/gc5HrIf2x4mUhl8PLty0kZ5l9Gk55KYFaN/nwmdbpIB4vm9qCksvO626HZYJOXuZxz8QQRCy
ig6M61nxJcuXI4x3WpgngYfgZ1LladQCK+4de2eX2acoHtS8KUz7ZSNDMCuOaYvMxR24Iro3RGvY
5nfDBkR+Z/TcR8IYpfNQz9TKEvHjN9RP1YmjN4h3LR9+mtT6MhK5fKsHYavYxuTLA45n6ZYoxZTa
nbYGZLbIAIbeVzDgLUWWuLNNpyS+KDGU/miHIP6V2cOF3qk7sYkzv6gJhqRX/8RnMC7skq3zYp+F
Wt1VkN5WXrnO9mzJ6AARrv5pvtxcNn6Gr54b6sPVeM9u4J1eCCeXOBL/Q1IcPJ+uOutZW8RlIWYD
55y5pmnY19FqK+4Yj9ItNUozArjrPDLQR6RNcj/eI/wV9q6rWNYS/6rOr6QUB8DcF+Ms5vxuEcww
8lk2k4CC14fhwrqZfv047u73/fV9R0YicetoEqgDHYP+bRkPym/MTMFyRVDnfJaLr+E52dY7HAx7
wpcU1dZCr61QFthMilxPI1iLC2hd6ZIGA0WZF4Ot3cfMNOARLfuPpbNZ8Gzo0dq6gk2O9eb+4Eed
tyq/u3wOIQjr7evGjVtdVOvWhEzKcq7AYwe7PJEewQ+YQ+gLFZcN6nmxm3QhtKu/jcA5Y+8rwduM
YddgNhmMpLV6v59I5wSTESCQHhnPPoTM4ICoc0prh847sL9arXrnTmthb5B08CfBugDi1litDXI0
X28Z3FRDgIUaH8iPlhjFaOEe4FzyeYjedBT+AQRw3XsitSVDSZ80Dxdqemxk8EjEfGWTCVhBwpqx
t2hHCCaa0autCsbzA88fOcBErF/3zQZI6ngN1NadZxWwH6TBIac1L81SCyYSCOxuPOckAChLmDa+
Amo+w/1oU4Fh1txtT9Bq4rHXcxeTMr1JxIb5SJp2yufZVKIteZ9sHrD7lhmOtaVd/KITzs82EVv0
UhZ93mcBdx0Du/4wR+I53KrHAOYztKTA73GprbrZ8gGZPqeGLfxC4rlrfykVihkz9OdAZD9S5DJZ
dd55T6Yxq9PZNz6768gRZ4Cs3OIvLONG7eShcPKFIqxtt7FaN3zBsZzSpAJ6+OTKfHguAuJgHR3p
+XdwNZ4QvNmRuVTkLOmVRVMNaoGx+2gzaih0/RlA01Go+3DDi1rewGOugFV6NA+ZANCg36E5zsPg
PgYLk+if4w2Tbdy51UkAs8Uz2S0gL6vNmhhb1JLadEM5aGyLgjsIJ1vJeDWIb3CYNiCyPuyD0fHM
pLJuTQ5Sp3WPjcCFhXBwl3R04ZCVW1vrDgQKmHbosNgw0SfpM2weZ0ClVXxiAQgxcvcjMiq6nMmH
dfAYLq6l+0dlNraYl5xzpDwBe+wfMdv+NTMiLA8oz/S+bmSrbWeG0FgbQNVhWLuPWb5PqI2hPQxN
T2MhiLE6/9uBmyGVyzO0sbXOkB3Y24yKP4Ep9If/nRq9+CUxuAKa2vKqcyLUltyCdSfkGdWDWt/Y
xzGhryA7gu6S5LFGoux9d6cOy+WZKHTbK8mIO0RDgILUDLYmxsgRI+zgIyJxGXL1o67An3MyKm5y
idBswx5djISSWMGmwvnQUJzc5PKon540tmiMUeFElF9J7cKpGlvyAwoVNY0EQhZn0ceORz1ltdm1
nK9IeCklkucuJsZlOwQitee4YJQ75M94+rJFKrqpTttx7ZE81WBmQ+o9iJ6QKSOjwZfE7QUhRXun
BVZTXbJ1ZoYYiGvcZwmW1ab5zynqy/sSf53Q/b2MRI6TO6DaD+gGPZkSi9CzncflfnWj8bKIybCC
kD2PoL6bfPqkqHKfld1NXGxATdq66iZf7mayNdT4e9xNU7tV4aXD/e7/lzBJYx07vsIGschF3HQc
RE/teRKvW5EdnXM2OgLmZM/5f8DbhAH66hQ7EMmo5ExHduTFqcDBgv/k3xe7ssfv60+cgKa6viee
m5Xg5mNY1qhCV1NxyOFbh8LQ644kZwg+UVCrcD7PzJIx8DpIsU2FhmZXm4aa5sCHF7v7mwPPWF7T
iQdwFt6x7Y9MkrMe7yigIZXgqYzqYwfIRlskjou7awS/zgPzddGfN7IAcPVdkMu/tR5uTBwxQeEs
MHWvKx0C2IKtUKu2ntfLumEyYxdomsYX0OUp0ssO4vC5Chy4xdXVouFGokHHDnz3jHk9Fe3VOcTc
qAl9J4vua331Qo12fWsMsakqsXVK4wGuLFtEdNGHRmZA8mVJejQJQtLhgERV2h5DsYOz1FO/lWKL
TntnfhF7TSE0mgyq+ZbSxxtxdxFOd0358RL2z2n5n+7IYpgdn+VgXOpHY30ZZeI4pqBtwrmGwmmB
LsxAadl6pqgkXRpg5l9FXXMQNS2FgbR1SQHrXejGhDAzNARZZXFFfPtpYfh6lGI9OBJQ65fgfO58
tTOyxSLkFmB2VZPHTsSBF4BqsLK5KQEkWfE1uY8t0iMEl3v/tSUYQJyDoETQT75gx1/swQ4XnxrK
jez1RJRauItniTVBY6YZnnnK6c2OhJ2uKtfeASzJDY+3TPDEz/ys72p0IYL4B0VlTbLfjUhbgHUh
i06koR62hSVjGC0eDFbNuFCPCrNuJe6ymmB8X8zQvpl6vtruzSJWi32AXz7TZxZhQ3MBZO4vlkTR
1TTxZ5wN8BzU51Yq4q3PagitQQ1rAUZUMapRSCjMSK6xCvRZO0209Eff7vE4C6UT/RQbZ7sn3KH4
R/0Z8aVMDdZyk/NeXPnUmC8Sn5q/NjuOay1/IuA24dVqWv1D4CqSzVwukAoBqhOKwd9Q0ogTPry7
BK7w+oMIotbdV+/mZbiuEOsVlIz956Pxgy612/lR+Y/bqz2yXawuD9EG0SZNC53HLOKiiB9YsYJ0
TwiNGGGBmOCcbkz56V4lKi3vFjOUJdVHHzY0rclaYIVeTusoAfrxNxoZXFG/h1GSPYZ8GATDPlOY
nPs2li0f+lJkCIqFKdGk07U/GkoRbdvyHnLzV0kamGpL68F84nnNnuWY/dHlO9zZHiZwTMpR4P7f
OQamY6iodBXKNGZuLaSXEZxM8UWtgzaX4+ZbWVD+h3XWi3mbCZIAh9UfJarup/1bWulxMh9pKA1g
E63OhV7AVcPDt/8GvFddHsfJVthc//FdciRORyjNVR/r4MGi+pxRATRlbwAxmINyA7olkMjCcfV1
aehiKjx8Dqi3pyy2Wrt9TQyv6doDe7xL8EQN57pYn0Jnd6wwJicHLMfNnCXxhYB5JVf0J1kURClh
+HXkaxFl94kpHC3Wg8Eg4chCmRFCI0WrGjrmEj0m2gmw+OB48TENFMuLIqUxdLWeTX+AoPevrQx7
TkitO4UGVx0Pq8mODXOMaAXB7e/U0U7VUYTxmcKIFmZGdQwhterA963bBBmK/jujafa/mXk4f6RE
0eUfnfrUfNhgo9aRq+UyDc70nq9T0a0H8TjJnfnDzNgj1vVhdKUYo1Wcmh1NeRkDoaV7se6Siu/+
TAwF3SPAjrGl0f7tltpvwzi6dMQJ7wNSFqtnusBnPzfN80fJuECKtNZT2tIk4jfnZLxLGa9wmVc6
ECTOSVIle3dVHEawkm2W5LzRT57adqK8dr49az6L28xu5itV9fZLwiejyJRkhlCvSN5GV56VCOeE
xGxayf7+/OhkYFdru17fLtUuQSzBim3XrkcW8oeDfxf25BP/Uh8tuuMgbJbkDGCkebxJAqsm+ez9
bcXonCfRf78lhixfEp3y4wsNH120Sw+wnBmdMYApSzGRpu/DxRzmF+LHsRth4dsFo+s1YyWg/2Wx
eGU9Hwgu+jMBReszSvKu61n8GjvGoIOHxDjnGYjXgWwdoBU4M3TcHdpT9ytkRElHioCQUv4SFEF5
lkyWuQdMbwiyQ+ug3qTLz6Rm0Vccka2pjHX8ZalG4HP54+cvU2ostSA9AnqGS9verexXeWPqjEK8
L/Hy8w4SdGj6E+BGpUF5W2rzyFhN2JKgeeTO6eNefVI7UNXH0kRrOcc4hEy8lKd1/hvj1aKMmJJ+
HgEUYcwE/ex71Iq8DAW+BSABzvi16RmhslnVY89XnR5NIlfs+Lm7x5AWmbZZpBE+5cAdLBAFblmL
9yI8rR8cz9JORpwzcTicUa2IDX1S5zf8ZtrNlqf3o3xGS3fwYolyVqvFDcJTEeFx5umbHazLVaXX
v+ocZB7OY/QNEiKe6HWTq6ZOSGCOw4mDQoVi/jjvsypW50ZyLwiOu1oIMB/BtpShJHn8miZkx0/O
JlQ8WloC1E8QWRB3VmbWWpnrLb3AW4TxPlr4C87B8XycwVWap0yMMyxjP/D8ivu19vKyTZbakLaK
2mir57974idTA3cZzYKpU+doDt9lO8TpUSUnjPbSkRFe37NdWeY0aNGuur1TNKapmMpn/SuZiBQ4
HAUOBIWo9ePulyH2AtxBr5Jz2XVhzamD2oQOIdjgxu3pgeK+qdi27l6f95m9YDYdsQxW4bgWFkar
PXPkYTUN6/WBZIhmxXZurY0X/7nkfr/eKZJ6+ZsJYhklHx/sZu5ahxwB3OJwcv/7F2Y0droinRG0
KmmvZT1tqWPqdCeE0ZYlk7UdYXXU0CJiLOY2v51iDuptC/Ps7BbOR5YZ3/NFJenroOWDyO7u4YZK
AfUqXk6RdAui2KbHa3DiXt87xEDraMkdy4z5OQLWpHYF2sgH9F7TY7vWh7sQea/QMLO3/kdDoHse
pVecY11gni04qOV5ohmNKMjXYUGedUiEEAXK/YXRlR5keepU7sh2aFDRSpHJ08bJ6aXhA+p3cld8
u9OcNLCdsWgHi88Px3tPAccShpyPWJueL5uhFptFtVxldrha0m94gRhzk98TtFFfNE2PSZ4qECmP
nYmARoz4iEPiw87HyJ/GWk7gPU1wO3CkTjPGF8rBhQF8DpRAETvKSl+p6EuJVnClUHsHmdpKGeD6
jKiSHNEQ+VHO7wdi+J8/58q6N7b88nFiIf9RcsUGOLFtduLIR6c5eJlhDbHKvMDbn+t5o5C8ihYc
hWTlBEYsu1Q20wZXBbFnrs7XasZ4S9MXIKpU2mapvnWCfazxgZs+6FQknE41te0vuGyBidP+YqTd
doSQLj6IuyaPcinIEBPkIzbjlKNudF+GoVcbf9QvtjFvt4NcX3E6lHr69+VTq2VC+WoFz0K7D1Kq
pHi+YM24lVYrYk3p6iraP86FZaLYu8i8OrweJHau3kj3pawNEJXcGeMrilg97gjNa6tqpQzpPusv
QEUSOmkh/C9ZILk2F+3UmQLdspNm7bH8BPF2tVCJRF5eoToS1EQW41WKfObIvSiZ41WwkhVC/hF5
hD5p15FHGsbAxKM8mNz+YD/IIKlViethF9T7YW9hLipPBdZIyqsBmHQdIijJaUQpO+ZmhRNxjTa5
ioygYfYMH7Ave/TYc+i5FVrga1lqL/7hVtlVJ7XempBcpFvC17GLi/BUTTTyPlKRznuHBWr0+sdq
oxrZG/g4IK46cX6CSfhF1kJanumj2/1J8jIfZJ0l8Kv2sCf2JW40D5ptKivZKLR4EZxEzy2pwBGM
ACNp/AAyL04s2+DZ7c5eN2YZCWCiKxybZhlLpbz8NrrsgNo7YTcwmlBckc1Zg8C2ivvjBNdJ3u8R
sUYea8a3asyGLHwiX3Me2Wi0XYSqWILamvzsZLwZlM5SLD985k4lCsozy3wxjTyUkuO+ulKJ3TJ1
89SAWk51kex1/5WXTH4idSw907r6IosaMd2w4sSgbcMJyuD3Pw0FEJeDKX4IF6hTZu9Ic2imyuMW
7ZWcCz5OgJGBQZkSRSWa9KtVBBwQz9Z8yHDEaDOtVOIx4Q7gFTSqWJJjTPg9Qcd54ENve9Oo1MFR
PsF8qZVekH2XYRLFYns79/gkrwpQgBPMZNo5f/mWgVyfCJ3tv32xu6s2MlKZoW3I3zvBAnY4l/fl
XYEx3iWgxinV6KJ3++9jjMjbq413xA7GUErmpsx1jJl3N59R6yKuYmP8fgkEqPCkXU0YzVbxOxUo
n5XFcs2QfIbvcHJFiTH5s1ZhoRWYrWpqMMp3tDG1Ge/F+NnqD6zdYud9CIcK8vocVH65IV00/6MS
0irIBPdSC/MpA/CM93kTQVvIe6DSX+urC3fw2MQRUq4qzHAWBbSuK3Lpvpl8disAiZxosjTbfM+k
up2w1KFUJvlFalcQvKDH89QHA/fMGVycj7g2X0CYeRDDcigypyTKPQQ9d0AMcqNz+4qW0GW0v8mo
kIROCQDGNxKvKNjCNQJ0z7/BTQnSYH5N2L8MY/Sv+t/8Z9ii8h9gf+fsbCrORn76T9L3LXyGKdXf
KZ7CcQ8Zf0kexbU9U12dMYL2c+GIhYNNTLuJKY7HcINbMZcKrRb9DgH2V4sf+LOAv3hDifnJKtmn
r9nwHORDyYmKpqLG3HDEOdkJQtC4rwK/lVSGj8KSRfzlstYtCidBLJHSbr8kArn+r5ZWv94XLWEa
D0OPpebKSiKdte15D4Bl0Wa23fqfu23nhtxwCrDm75LWOSZx2X19kdT6/6PCzNo8sgUX79qHyp9D
LCI2ijG50anH85xADFlxZqyacI/C7BJE+qdnFv8jVUTq4Eh+5BAy/RuKKK7OUaagCCNPYNtkDnV/
qRy5HxYsejxJUy4dkD9jWqdkB3r1xNUTiUUY15GhDiPJvHQ86aCOtJctmSuEXLKHy06kzmdiugsT
OUmuCrBwbErcEO79E6wbdf3UAd+OiNtxJ66JsmKuuZPNueFQK5soKvaigpYQb41yWsgMLfPJ9yJh
DVxXgKsUL0bFKuif/cyT4156FJz5bTlJriHmg+PLGaJgdq7jBgic2mxX/UmA+ZJv98iNogGUMNx0
U7lE6GIyhAvIq8V+hTgYe/KvKpjonCpjnI+HyJ5ye85lpT8e1+Y0AlEJOx+kdsNECh9Jq+NCQP0j
adW7DlU++5T7Q694vAByenLA+EPb6CwVCNGvXh0pBetncKCf6v8vKbZfGHsDBULoVydCJF8coUBG
1psTCg==
`protect end_protected

