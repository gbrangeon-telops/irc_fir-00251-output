

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cPZ8vU4rKWICMycnP8ASghxteX0KiiSQpWJpCIK7voNSpkWhaLkY+/QNXKrCWexA6C73eW4MlVqP
U/aYYyUL6A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LGoeeEeMUHkj3xBumwl7JSHXwdKJWR3APWiWCdcCy3wVC6g0GScQrp7fjvXp784YBiHqjtsyG69d
mOZ3fy7Gj87kc/h2xvc4Kp6GM/IiHJc0mbPVp01AJelfAExlIEaVGoQkcAXR2aVikeaMxuRKkb9m
THdehu5n5eHx4/tJQjQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aia+xx8RLMhA3IF4tHoW0Vw6LtYVDVgU/c3FBWk9RJ/SaLw9lkXng6eXJGNs7uUJXmkzrbSEXjkp
9p7xWJMhovE7nwsp+7RydSgRQ0ttqPUbPZE1eqSc4iNU9Q/KQ7cPFMFwb6o48JfKidjAmSeXX5a7
n8A9TbJ98klc/V+a8Nj+tTPfVP1QI9dRmdzaW2w+actp2BkWAgSALKaGkzvCVGa/MpfN/fdLNjxo
VsiL86HW3arw5N+Ra4HD3GVUtLt9RoCCVRrMaYywuIwp2m+MgGVDwi2f2wZCZ3t03UamXKangjoy
PBei/XvAf3p1OvrOrKNUCVdwEg17DQWfBwZyYg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iSq3so3iXhp8LA8lrAo4ElVWkZ4sJhg+rWrioZWefLcgVs70gDbHsh3ghf5w2wiNXalSfMYzUoxO
skfS1+28WFbvBvygndpiSNMXeXmzWGrwBeHtNO1nR5azyndKvNsun44/B61XF3kTINCJNR54A+3f
0Ezm1jX/FmstQisPDpo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fHCdwSqtdLKfkpdCYo92uS5kFXmPpII38bIISEYuCqZyK6/BVCrCUL1HNVeJEgqGnb0uRqkye2CI
eX2LoUaDxy6iVejnRrRRAgNtgrlZcFVc3u1KxZQXk/12l8pxvVZj8jnWgIvX3TEsZsoZ6w/D41BC
6xhd1LtUfJeg6bsnb+yBYV5+H8NnHOqkZuFtJBsUzS1+4qFALyFqcNVJhhbdB0k2hn6z9cG6wZBI
hB8OJAFj6xON517ug+qP1OJf6uK1rHsG0pxYXoT6xch+UowAmLY8V/4+ShcI8rx6DLYpPvJVhEGV
fj/RQD4+HY8CEDIrJcGjF+Rpk986lOFjZ/hvRA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
KQihGqtzFgiKpEZe/QoXAE2kM6WkK7Z6Hsvp7hhWXab4M0UF20AKQgvN1NJamXmsKDRF1MPVFpx8
WnUl1iI11vY53S7EaGHX1nP2k9FQ8OQ1VDuDYqBjerJzixuoAPmqYIOuoSONgkMGFH5QORi6AnFj
qUN3Djjtg8gUUfh3B/yx3fSDzmakoXIi5DPljJnVB+2o8PyaQx1UwO1mR5VdMlHjkXYfMlGYsBwg
VKe3jeIRnC5uESbbT8+FQtwC+YoXK5ROOD1lMFNHLoBdE5dftvoNgqRvH11WZGWBuQCQenRSIkeG
5jaQ8ibS0yKcqJDDkzmcc9AJRKmCofSzMv0AQDsiqs/U0V4l6mVl2SIqtYz5kmIhzLsmBZE6qV4z
IlZjvDzln+dr6PWy/gFJkc6mmkQ/aYNNdlw0JIeK3py/gnIoYY5lNu3VdjaLFMK8EF5otYvM+p97
vYuDaNGTzW2V7j8Y+Xpheg93avQKqNepmXuQT2ouU9+lDRBaDX9mDAFSRTygxpXyfIO5v0on68DV
J3bVdG2b8wyrVABJ/fgb9sRdypl8ZOXggecDQeDZsBw0Q6GgkMmJj5m/jb8auv7XjuzoHczS4kY1
UrxJrvuw4PXsSFp46uUWCFeF+50X7IEcovIFH2tCJVom/mb9GQs+jHKjlk6VDLd/Oxlxpp8OOR2Q
10D4ALzIQp6pwHfXp4Xyagm7zkkmclYoo0bPqAJJzG2LQI2BtrUyiuUlZhe5EaoTY3+8SjfsjaLd
i97hs7R28g/78BpRr+V69EDqeH8oA94dd2u1gxvA2+el5ptZ4mOGDHX0G3DgVryZ/wBlOp0i+HAQ
Lj8zXOyfDkiw1vTUWzwPB5nECCwqre83m9ECEogSsnucQ5R0sUqE4KIHWS8wmicYouCzQYrFPfSt
5zFuZC1gDUl5Cd9dInM/nGwy7cH6GO+EImCrfLE3Y0J4hdrmNKbIztbewRhGjP9e5UiRH2wPMymN
3qN1NdZIpdJjnTOwXywCrB7hcu86G9Kq2HKR+nu+e/UWuw31pvJhOpruQCp85VvYwEM1dKZPIh+c
ENSVbyH2czY8753u2xhApjOAzL0HP+ychIPA8t/DyWe7YpIP1o7PqJTnHEnc9UzAMNff8xRWOSez
G9oVxQz745LEe2llSeJ+LPLsLx44RzpZjSOrxGwZhLo4M/tWWx80HFCjCJDbCrEif7fE/+debKQw
NRTK/J6AOe3PWDfSETjtkJG3NRFDhOIRI7hGYR8fchCDCkETWY4JXuQX/24d2Zji0k6Tq9L+WRPH
swb2QyFE8tL3BWmSH/2cnHKRFbxajJ3CQqwFa7v8m7h67zu9QkFfGnfXTG84qlqgUjobe7jGuNT7
NoHJH6dCEVGJ8W4u9HRLL32qu7miipX23N5W51Bprz3XelXEIjx9rqhAcZuP0aHopEZcY/pk4fq9
cyz+149S3X5OfqO3+/e/uZmEfMNKXXPkCvhcgIXluZWxVKB1iJC4VByURNdBlOBaR60ZRtZiwHPP
F/xKhuxliGOZQuNq/u5RacymhrMa6m1a+d1mjObnDiELHlvugn+FTPV8hIcjKyq5K+Q3/L21x0iP
ttP2U6kR29qiP0dGsOr0+kVPziAME/ZS4zI49MTKnxztNWJ9W2qT/UCmbUGgukOYiP0Kp/mkV3Ro
lQ//NWcm/neyI2PNacDhOt/APfVgp1BNpPDgkSz/lAOKrSaye2S5Z4qphiyn4L3tz7fr29Z0cxSv
aa/zR6UXU4R38t+9TLMKlQn3Q47vidkegzUN4rmWoNO6VtYhaIkdqhRwq8E0Bf7tz8E+sXY4TVUf
eiaOPvgeoW36UrbE+gV2zSY9RlE3UrQuiEeyot2RvnSgQjgMEOJ7pD2XvTTuKSE2GHvVVClzVFEA
wEh2mVb39VhZBEQo32Mhoqsr+Uktc3q6ZxYJ0hMNGreuIt9/RzVbPiSR38H1lEHnuzh+dNBlNwEa
g54QeEbedAv0gi/ahJySdr498mFsNZ8JhmEEa3TteROVevsZ/pPboXZPEOkc3xHvqqgU7X6i+UUM
lqZQyFnKOZ4V8qh9uuTz7Bi3gyW/WslNd9HtzWVduHWa3S4b58jOSSw8fdK6Q+00UT5IVKfOAGbj
zmyMVlMw9G2OJ+oWz7SqZmkxb5OdUVKrDKXe2WSNghwXu4b5nrkTFyL72rW/MDfR9/bD0CAS0TXd
9emLmCG8yvK3tatbNnB6IeBZzgiDTG4ak/zaTk4d/ydkWH1O8lKWbSfuQ+wmXDUp5eQgT7hVF0Qq
QMulC5hyE3u+gUM6t//ATGwKPGnqaKpdL/MLCj0dGiRpCaxWwh//9tIgm3Y23wv9TyZdbCtMGzCo
oNauQCIvHVrVQ1tlWY0cPcm0XmMOv57t8u3DHMg7iYaOcHpzGMP/NoNoQuICutY8SyNGhmvx5EG/
+cdDFNrcsia/GW8hP121erwHpgUh0Zdt4FMrYSVxE80L9y6Pimpd0tDTp1XLfuViHLeUEwjmnP+v
HaBACWx1c3vhJdjVdp4rWvmTQQeH9q4bu6fcXv/O0JykPDXi1fpsNWvkscX0kdh/IUXfv/9xWKkq
RX7c0KkFnv4yRvFdjC9dv/win7NVKeAMK+C5pZzt1aLVKVRZi3mPIrfQVSKekqmrR+BY+yvUTLJL
mDcvNGqn53K8fAz5MUAJxE/seUqb3oYU7+MkoR6O5aOJjuGzzc2iKEtmhbOmRN7ZPDHdJLyXITlu
hHHDDj+BM75jrt4kfj8ICFkMmxUz3wIXp128oSZMTIT+v1vpFH6FMzq9sg266Fs6OI2CwYH9uZ2v
dMaD64kSFk12rZr0zLWnx1RlILeCFhDF7P7Voqo0sdKxfrKbV9qccWModeyGA8Vyzi1bVczXPGUc
L3CS6PVHTqMp1iYIS2xWtdKa9gEY9QzbJ2fYmbtNXFKQ1Zyt7QxuTdnsQig1Mkj6CDFpI4lpNftC
r46qBgWkTvjidCC6zFbaS453f2hIO8iQXqQ+0W9THffvgP5G4ufGIqfZ5R0PBufOyBb8WQ/agxP9
VU8JLlfBmwtJAeur8eWnOBfZx0XYW05rObkfYHccPFscRgrNg65+z2lIpNphMLXkk6xik6ISahp8
CVM1ZqCzq7U7CwV2PJEWPBHNXjI/fg34fOEbwm7x50Zjrs0upSrWb8z0w15X0ShFtgrIV1d/po3z
R/15stBCeDO/bgbu7xj3cTsPR/UXEyb1j47SA9jQYBSGnv/TOVcZEb2PDtqwcgvA6z5ulQ9cnxYi
DFkKk2WefpdH8dmgJsbXqJM3utbPR7WrGISLzztK8Wade34RQhiAyYaD99/ZAFDcyd04siv8HrnT
hQa6dyk0cOIpHb+fKspGX+pLkQBAkHkkiqoMUGYWgWRUWH1vmMaSQmta4qHBJ23PFHywF2DzKbo9
dWssSbIh/OA6HR9Fe53gxRQNCBCBYlDkOPEuxlf48pwG8ay7imFHztZJ9J363YtkiBnn8H/BFpHx
y31fnyBgCsIhKBWfoA0VXrgbT76c6HPMkZf15HiIGweYBAgfbMWSR9PVW/dVrwDwxJP/qYfsOS+z
a2kRtHBtXmaRQjbGkZbIJBj/58xsvA7OrViGPRv5+YtR+Y26PQ9kNMzQr8zDbTS7y7Oi1HA+h4CT
enAaJ1MgCM5XTXf7BvKeCU3LoykjEjgApTL4Tt/nPjENILvCglK78mm6s4qvKEctGsmt555VtHYo
9pHZohP/jL74+ruQjEoNJartT3uIfl95ovT4zRCk0EyPoI352z2JB554KLdD7wnyOOJni8ovxOB1
j1yqt+cd09jsS8O27JC+UUmP566VkXIuXJ532KfzqMuQjut6B5RqMJbWnhdv0qTptoTnCyl0W0Wv
bbz3WKCpUlM3YDyY/OLHYCTXUuCWXIGV/9I77e2pd869Kdh9pRHe5EZB0W8XN/UXCsTfoNh5cIKA
44VgqVgnBPxDG6PckJ8VgUAeKiYk/72ntvnt8QsKO42brswtmQr/X+Gd8LfVBJjtkB+Vmkd0m/eD
FohssTmNo6TARc01Hxl8pqaQGv4VxVYwtlnq1lMB/wZ6POGWoQcpoxJagGZAEQvD/Sw428/inBiV
e9hshAw+IvonBEwOKBbjuh0WJnyH9qpxReI8nDxuzrmQDK6/nkV5ieKMPJWwyoGT8TZeN4DMHkFO
sK6dansQ1p+sOTVkEVqTG9ic/zxlA8tb3XEX/rKjjLxBAvdYVGeQxclpEHtbU9DWAa1AyWgmq27f
evEZYhlzlv1OTiPitB8aUuER4aAiYQuQhKc2V5UEOlkZTOPzznnBGqSaPOdWBZxwKlM5ZxlfwMzZ
XhwTEOvbfy86xBMQzOaciYx32QUU2gLHoZyNxVxGYsJ9vpz7fHjQs3obEjm5yu0a6v5SsInadlKD
LQjP/PZRMvNPp18pQVdxi7pkGwOfSdvfpe5aRlGiojFf/HzTx81dgK+qebkx0ltTct60GtRjv9kC
eMZIAG4fBQQgtDj66VL0cvSAxhwK3nHgRGZY24woziQ61wc29MkACAOJzVa/0TxlvThn3JwikbUO
9lYUdgmg+3NfZsVEHHoX8JWcSg8xaR3sNi0xxOFCXacj2XFZsp+TZyonUJzCnbbdrHVx6sad3Vbd
SaqNHzBm9BzlNkD40fgo6r7dvRWVZIVoJHJklihaFBeyiURael+Z3HX7jq9JYgaVxEdKmfw3msSn
W5PjGACiX1TNwGjimiBJBrhniu/B3XvB8SItr1RPtfUo06yQq/sqwBjrq2VoN4gCgVC3z/v+huZx
EwxfLC33zg4AWtKCb1a8DWF9DSTPatVCfY8bqupknRfcc2RZasnFZ7S/81yBiNy0vWEKAMFt8RVq
TKrUz7nhd32hn4Z2NaZk5g9UgCNoqfv/BOMr9RtFMl1N1tbGp2EfnvwbReWPHAWWeQfvBk2gE9Wz
LZBYK1oOrrFrtIpv1BtoZyZHZWZe0oqbJpbsQSBsPUmxeHToU9BIzKzhKk7Zy+B6UdAuwwgJ+2Qn
VqkOhxGm14/NEpVd7TQ/JMjE8gMI0dusCwS0ygGZfHt3amIySlkZkQR3gG6VJp4+BObJSzwsWRcP
IRasELI7bja3w7h4xbIwNOdPh66zvrxL3/+3ggNb8KUT0/k+HRGdvCcwunobjuBdye2xXz8A3SEf
mXpEWF+/NSEdXg29QUY2Dac6wk7VC4SIdVcvXeen23OxfGoZVXJkvRQC+F1bWjYXPP7O9aHwSe+6
6RiSj3EbMiDM1tmhch/pDB4NtN03Kk176vcBpf70fRnQtuQwK3hNJaH2/758Nm5FaRRM2OdZw0RG
53aW6K82OxVCfzeMxB2hs6roeI7cw0mmt2E+/vn4JyBh9HwybY1Xlzk8jk7e6uVAfX6gcpt0U6RQ
SvOqk3p0Ik9TJSTawSs8Pqm9wDnOvKTmldFu0vkqHHQZaESf2KMm4eEVMXhrFYpsnhr6rPXK20vF
8rQiXGcN+wieB1uH1E49vXwZ21U2sl/41ZFI9ViebHLEDRfmkE28L3yQpk1DNT+qIVw+HQdwdCWg
LM0LKL5yS/PooWj+euC0jlSIU/alXcbM+AqUzCPD3v81auUrac7GS/P5UgFL2udxSHo08XOkPOUm
BZgH42skQWtckGZA4S0wKRPx7la/k73fbfTOMAquNvN53+XK4DcK+PA8eugIn0tQTTyClilBLfdW
fkIiTmdpeABzmM9siqZ1KeEf7lJ749DmFXQYQpZXMdNFkbpqwR2j4NwYIZvz23yb/0FcXDkOS0CT
oAmckuGoAhN2O4JKGEDoi74cLt5mKiUwP9zoE16JuzmNcPFW8AkUtQ/j2SlWkqmhMhlLZMC2z9xG
Zk1DK3qnlqrhvq+/vG53qqCPzuA0Fn2jCmLf3Lxvem8ORFavtnFMzqxUD+iXLrQJ+JcSRijTe+rk
SbxOAEESJHQwEMlBszKgtjw6i2Uyo612bAAl7FMoqvll/MbeRCFxeQINjtaDbjwnZCboOEN5DXGG
tSdISx3c/40+Cv2FUfOGYuiHlUtCTvwk/PgSKyNcIRqdweIFWylGcW7a727y6MsmiKS1/36LVI1a
hg2IQxj1VFKjGGsc3moQfatFTjrLmE1HJt13oHP2OjtZJJNelXD8uqsvejJn4NBxHHGL0HlKHJYA
E+q8nA9BsuHEVce3S08TSX1MeIqtmmOW3h7ps24CeD5Cdp/KsMg3Rv3LxXl3F08TSH3JVVC0WKBl
qWDoFLWJeVlJ29ovuB9kwAInNBU4m30q3ceylGXm7Z95i0K3t0kmIzjNbUJz6pWaDftSJUqsZpyM
yuljk0CVUb0N/th+hmn4tAgXBGLhRdNS6ypW99n+IPScN5L+Cb++nFnVhOMCw8qg8/UsSbXbGIVO
1lYx3rnJb4bkntcLo1B38AikNmiRL0a42a/OIwNiQYJuU/FOtoX4C8nyk17w97XF5eSds3+6lcGR
xOlo5JPBHDKqWeXO4g29KDKRKou3w4L/FaWa7fBAnVFDAk1FgDw8B60IyFtyApwtaPyW9Q5IwpnD
lemHvCafVe1Leezoyo7Mi+65qH11Fjvl/ZK2RFvPbw7VlZmHQVGnQAtf6ZkIrOsPQPDPGMM1Zk6n
z2ZeUjXz5JiXPjD88tGUZ1Noi2FDnGiBTyMHYVLvkLooGSNavLkPEe93DaI/JnqI+DFh1gkf234R
1KX0kG8gUdq70IyUVJRDax+3ZVK9qkLNHpOycExVzsRfl17TC1tf2I6/wnr/A5DSEv2f5zbEakCd
2sn45WV3gsfwqNDSa7rUNHbUzG0+sEi/v1N87S40G0XIs2iRVEmZXnjhFXfUG4isE+Nip/sOFMmB
XvjPBaNGm0C+3hALeRi+Gl8pmJabIcckxNp729mp5R9nFe5NtYG8T0sTkSI/Xy4vHtLBCMoYY3OK
ulFp6ESkYb/6bWRv/9UDdGX8qv+m6C/3ZnP5JaSZjLhoiLxfiqL/Xv9w8b0sSDCxlNTAqH1lqOR6
8HNAG0MrLfFo/4JQLGKpcck03Efw8796k7qExlmUh+zFdSFS6Ez+M5gIL+Z+CPec4BiKrWOy09lV
q75rAM7YjXNa9KidhLMh7jcHZhqdLSy+D9C+owEgiv9JjIH7bplCJm+Ug9IeDsqv32qsRVIJZxtZ
2k0GiLtgQVSxSqkROuoE5r1f5uKAXQlw+SqXR53VcFWwmwWJLfrVNqX8Ek03Umcohb5JpfUeukUp
pJ1ZvwG6pNXcfClE/x4IhDm0x8Ytd8uY21EQcTG4QUSbo7nMo2olGQMUOboOsCUIhBYvFC0IoPwc
aMkSht+Fuz+nieCC5lT/StMKdybSdUrXg5fypeDG7f96fwrt/yUWNHSXGjQrM8lqxWSbQhLSYAq/
xxDL4imT/uFinFItFuYnhEAQiyA8++rFixYoZ1ng45TUVVtagMy9KZQ0rzItcYQV09VlVJne6DdU
iRU3ZItqhFFQ9UZ9Xbs7OospLtK0t4ZbbP0cMVtrPAtozteexd4pqIhyZbuGgxzHfXfTHWJU7+I6
KcTV4QQxx9XzF6u81Jt7NnG+voWIJW9navwQDA8lGxB2Y6DGkf308PYQNXt3F4pHxXvhKSEH3Y5O
pxCQ7h/yF6NW+DMxVkTreF2NNjZwCzYWf5yanzJNZ9poeeYxd/PSNC/nPa51NR1gC5aVoiB6H4Yn
JXCcKzYSOF3goTNKWhNplDnKUBCD/N+RYTWnraBas+wgEhDLinvfDaFC0Zjz5MI2iCRQhLwMSDPW
vXYkGjF4XW1OmDh5d2VoPJAIQ6mwRoIYIVADV7cry8BBGIIkPviGylpj+KpIKgVALmNx61C4zcjR
2igWublOVPjukI7BksIJ7E7R1ZqxrCCR4F/qUVFouArRCCGO3g7li8CV9VDX9swc++Nxq6LIb5bf
BvYlFx3d7BZr3ZwXi0TZRSxE6w9NThx/dMIFoSxqriXbegsgICpa/MAs5XOWUoecNtfJTw0gJU82
QaxYIQN1pmXAatUkTyL6SOnxv0SAqr9yR1/TAr7eq+TJHHqV6j4KE/7WnPzbv1oB0H0NKRf4kVC0
RkvuLZJ+0uM8iV/h/RmJaMqxWoECEexLfc0TGrMOYpxQZrECpz/FUQpr3W3XoS5c+6zbNfhcE7bn
C8TD7aGYD3zQs2FlGCcDHPLVI6Xqba3QRvUluBcd6SeF/6hFl+Zg6d39tv3NFwKwRDbkqXiJj/OL
A/UqIa0rI3SYZWTZF0uO5mxKXhG0k918UwmNQK62q+7TGshEbBkJ0LhG5ME1RcOxwulOx0ZS7Qhh
19y/D3l8jsEU5IRneHMP3M3YgCp5gQimxxLk8Xtlr1LlQkFMSzyiMOfTrbszXrfwiv+Oh+XZP4El
aNhbOEEpDaqIktw1Ng/Iwoa3acXAMMC6GeinhOU3YBlmNf5DOGGvMqDbNfpeHUn6VeG0JncbNgCg
kCZkwW22Tq4fKb9rSeErT87wvvj+vtO56bqMPy3AEeQps9FfuhnRr5p+ctqL3JZRtXJgDfh31Tq8
Pof0WBUm+ngP2n4+32FSsHcov5WY6Rbff5KVgEbgDS9hYIdvlNae8e1xr8m8vk3wfFa5fOJuyUb/
ZxSQZQvfKHwfaR96/GjyYpJJyDebnvehqT3ZI8buVPcY9aKa2fkndy8EPHhayt1dbXaiytIEZHl3
QHL0rN/C2jopsYPjNDN/indI/eQJdgAH3njBDkx9VwOv5iDLBokK4Z5RtlG7ecN9CucOV/S62RLd
Uph68Oa+GOxJG+cfVtt0jwfmzpvtwpOs3ygc7HMxdCH4ynSdQlJDE5feNsuBR4SgdhbhTaChXSCl
jVOPC2pf0XC1eV8QkDLgsZKXr32VZdaYKFEjb7lE8NNTa65JyFoMUY0DPMBBzxKc31Brf3bHisEl
abd9hEIoxwECxBoM16kG9NNl/7ARruL69R4z4Urb6dqYMaYxBx7DY+whuJ6Mgtac5tdavQ0QB6aq
8MNGFDLL/k+917aYRZTTONYWsPxjY78nZ04B51+AnOsc0S/rrANFQvF6XNmTe0rN3ek4q5cb4Gb/
VhCbBXgDqLBVsBPP0Sc4wh8wO/8VoGti2CPDuyb2CMgIti9LHbtrMe4p65sL1bpzC4bkiuw5WwmB
f0V6tKrWPNmC8sbLrfhztfZAWI+QW6WCqPHMQ+hEJXyzTYZS+Jn+B9fEyYaTYH0epGdQ+EwaxP0+
TXvQ3z/g7vwBAkn2I8C7uCfHQClhI4hHT47ml78hNI+nSY8ppx8AfFZ4uyohUfRObjrKgQDFFDXO
tZjqCzyQGqGWbaN8OncKXA5dfMxn5QF68M9LnzTSVJa5T01Zg2jIupCqw1mJX7h46e0H0DgNeCIv
ywZtSa3KVBI240oKCQpF/Euk82B4UgDrLPG2M+B0x2xQWsGeF8CgsMqoxcchUVp8V8YXmVZiWiIV
gOxyhpQZimqlfRwGAaz0wrztTmoE4AjQiwfNv1/bG/Cl40eNLBAjTcyp7zhBSGQdHtyqD/qDZE/o
C0k09BeggGGvGLG7sXppKie/hWfQHe7Xrqhb4zaz9/rx50u2AM7eAKjy/fV1Fjr3NdJag4XLEr0Y
wy8gI3q2g5FA91vOtahxAF29BzA55NvkEFTyg3VF5Y0QJMBU7Wi3LTIOyyuJLZuUtC9qO/JgeQMM
ZAvuGz332K/uXJObIQb2g6VKVl+ent/epKyrbtDV7a+2WqoLaqZNuyaUuP/DIOn+yz58aTJ6VKJQ
oMsIsk60LBMgFUpynWWAedb+AfJoWNILcIcconDpwyHI+UQBNb9xr0wM2TZo7dbengksJDMfxCCZ
BvLXZFl4i7P3ESFPd+SyaysOJHvaE5hsXyHgqX8egOlN1DVGsz3Fc1Z41EfGb2xQ/9QdiQLHKGZ5
eoCQxvwmGNn7mRomqnCkyLrHzzppGb7EWZSruP6Qs9/SSUfhoECiLYi7UEbauNJG+AC+bGQbYK9k
RdYaYPL58q6HC1ZeUlVc50+TwZXkCY395k7VDxWISY0XOCeJ/8MsK9fdVcYbuyUNqFs32Lx9JCAw
GCPtxUR1k1CVxH+Bj6dMm8vTaMXSJ+LiUOAzLKiE8Q5OmI8DucXcrWbCOmNDbaP0FniNEy3azx8k
/aiB35DKXjgwMNyRf5GI/ar8JNEMeFo8uZEEcYMr8z9Jbt3OCAxdWVluOlI9qKBY6QMHtEGbnVDO
2Bsp4xE4mi+Y6RDUk5yCXnSjNeudKZDLh9juNhYk+gw4TO0Ans5dRl15Xh6bTI3g1RdmUdPL8WkC
8b+Zc3Obu/oaV+B4BDsi7SnXGjkPyXvykMR4rMJkRYTis3PTixkMrE7WTU04EwuZ4GUGFdB0dX/K
hzoGrHqPhQqW58mJrD34N9SjKkJu5B97xOc8YsSqOtY9zigjvGD8VRhf14POW7RDkgyb3V4Xh0Ii
Af4t6g+49thJtf/5qXLPLziftWm9yWKJSDNxxy+GYn2a/gC0dUCxneOKMyCsRHBZSSJJIOHfZLhZ
TNhK51zBRt7TBn+Dl+BCE2BO/xnaW40lVLGg37pma9VCg7oGEChfVRQ/fEDEi+ejJ1TiOA6YD26H
N5Qh3QRKjUjJxgtlwdoFGS638RUshLAq4F0GgEDgIuetA/IV0iccsTmeoF8wpuSchOpcYAU141lx
hQ3XO2H0yQp2IXK4iZdBy+NofdjIAvSuEP/rz531e0rDiwMUCwT0iaPuLiXgF6SYwt3fFxAvahJB
vwKiqi4tMPbCZrXPDcoNeJCC3vZSpGOXvxlRZCmPnnXutkTGn6/bq0R3Zkh0UUs1VduajgzljPcP
RAx5pN97ZTvo3igI9RekauE3G2jFWC71dxdV6VXNNJPPlmgkcMtg+7jDcQpLyj8UzlZqlJFJA9F3
dmLVtkxA+UyOx7EZnOHuMaUiK6rHiN0Xgzz9Akckg42tYKBtndPGVDM1fd4jIxrjf1FfakO02ZQy
jf3vftg3CU1ZwzEhZ0BUodaNTrcFtQuvMUjkFiaeWZSPaQ3ojEloTK761mx3sXWwRkOcEjf4a03C
MwyhHbwRITWeVdZLrdLsLT/g6QoVfOXE0sfFOVJ/gBjDGBvF6AoVK+c9JsoUlkSJB+6MoaK9kkv7
j4KwiqvfViJmfQsUlBvlVcwJFsynfjj0iTT+5S3hLw/Lsn5IurZy6xd9znl4wOt52+o62tsbWNqf
Ebhf1DwX7+0SfgksWmiyg91hj9I9p8dUdWMdj/diU6chyq8LBU0/e/2KB6xZ0pUF7ARoQ51oLIN9
D+Hn0JF3q6W3QJk2t0cYOyugh6EIKMM1hwUcIvlVazgXF0jYnOmg3K+EZmHYNk0rA7mpUO+FpMJm
N8V0UCZQZjYVjI5R6dIfL4QbunOGUGJKcDcuAqi6na5BPOyNu6udYpHk4HYweQTUoVr4lBlkUYeP
v1IlMt+vmHKA7pmWS+VVhExU6cFyN1N5tj4Hx3wSLuChZw4qrGYPmTJ3Eu52YeXeajnswJ7+zxsK
D/+nbZoLa1OgUrmCJeGd3kn7f30O1IVH19FFiLuAACBqIv7xhXVnJgOuf8sR08XBq22xxQs0c3G1
2WAIoUiBhxbR5Ehsmbu6dvS2nhjAzMIi6zYuHlkNbk3kvbGf/VZh6xKlvSDLuAi0oSBd5j8co3PU
UMVaT/8pZui7n2lkPxpGyW6IrEl+Ce1YJ2rpbMMZutTzWULCWkpHhlR/uRBzkkOxriE48SbRFa8M
g6qzesVLj4WjzUlJjEaa75S0qEWUnBUzKZuIZhH+TMk6yLFTWUMKJQoCYjoIZ3Jkt9QnUsV1f7k+
8m0MmMbhZKND/PwinoUnDbbEmLACs5TYWwIifHeTFm0lnxgct/W0MeFQZFGJw40fIByWbFKKp/dJ
+R9C7Kt+AWDDArQx3QTiznnNSo8vd52sChftHfI/IxG79wViK/i8ZapgW1fJDsmhZPl5LSi2RtSd
UDCnmAAj5N8F3JvLFZF+pmxhzo+/zqB8PB4/uQKQGy7FkQ4DLosgimsQC+My0hh0PQZUnwO2kJZa
aNs06PcoswvX8Av3s9vKmSdT6HavB6id1AtBrIZk2v6B7Q+pMoA5oFYbvov0JEHqVanICjp3FvQ6
nfIVz402bH7Sbhzs69oV/hZFh7uHNvzhOQVCToZqmqdl3XwIuhX0WygV8RPoSwbjfSKL5qjbRVDG
DbU3M/fVdTc8Pcj7toe1miMgGRJnquopCl+586YkHmdhvzOWvDhyUdR78JflhgE5MdwK7j33RGZy
Dk3i0Fqr3J/tjkZ9zk0gexSyYPVlVGHkFaAYPk7m/XIAQ1G1teIoT1LcvqGTODaZycme9lOxEYcJ
ivhYDZ9AAvaYZL0lO9BnM0WbDCmmvUBFZEnlsXcliq0Nx5KuqDNuDa5ymT8wTmWvhILSnxGKgYik
dMNTdJp3VKt/yQO0kCqxhrOn/MDsT3CPlMqXLlvXloAAJ2Tf2CPcr0oom9EmRg/68/iUFsjXlGoa
gOd+1YY78HMNOHlR84eERpFPXIgym294LEHoEfhoIX5RH2UlMkHucC+5x/FNOy76DCkhGnK2f0r4
F1qoCbGvnG0IwrB+SlL/jVvbms5NXZG/GYU57Sa2RJKlYSkE+cAn2R9l2xoc53DnsHyerA+kWqJK
z55LHtVsOLyBdfSgmOSeye7lczixUOIhSQXf276Vfd05OIGjabi1W8X/UaBXcTuSzfsODgWYy7NO
39Ybri9qjUs2qfu+HfXUlBNShR2DWl5Dh1Dfvzxe6Yc36ZpK5Jn+rwXtfE7mQS+FRWiSR9h0FX7v
3W782KRI3Bhlxddy600oMZD1wh+DggrVAPiWliUtelFzPfittAUuOYRMVGoOLUUj7yPEgyqwDKHd
85boeGhVIxypO2Aq1xCvJ2aFqoa7ruge404UGJG2GCEMfckzJJh00N+rVA0YmBakq2ft26k/eVIA
y8Z9XVPM67/nFGtWOwkpNz72rS+68Sff2yKfQHDECJck/N+52s6RHh4+KN9B4zDWQlk2SAs4bwUZ
y+ZqSPrXbqOZ6VBuGoPLUD5w5Uo8IzWrRQPNqq5eL0VD3MpRSTdAc3vmc1TiXB+hq62Zy28QJ2Qp
CqvfdhBc83pF14WtybJN+xa7KrKTWbLSJGB6eed1+5U6Uir+xpIVywDn5Qh3Fr4QPMcX1h50CBhl
ikslOY872Ce0g7x5z0PFHmpOXIkMy7nM+hntOuh3LEcEFJCzxdb58ma9hvUS7AERniOLzx9+lTj1
PQXeiWSX0Nk/6eNQSE+uWojUf1oJa/BVJQRfy2q8G0Qo240g5ob/K4WezMIOz2+XXoKYXcVdhPE+
nZTjQiTf0Vo422SX6HdqKbMw0JsHU9MeYt2VBbcKhVp5OkkKpGsHlwqHPgSyFFoYoVIzIdLVRgEI
H8KGaPTayj2t3Hasb/PkPxi6n0PepeSg2ryAEXrOoT6ElzOYj2FZ8BPxFolOTLu8bj7F+Me37UZz
MMM9T4MI6QQMwo5vD1YxKkQCLP/6WPGbT0P1NzP40e4ez1TgnZ6PDMk1veHziaJWBDRByqLXGu8f
r+xTX3Njy7Tf1zuvccHlv8N3Jcl1VAuCl2MYE0hlFl5vxBsQlQg8KHdY1AE5UyUreh3So8G1/uzN
NS7+iTlulXkfD+NFo5wygUCdbJs+HUT3tXZpobLTlJHtHU5CqV6b1f1EnWHvzZXPyh9/OjIZZWpw
d4tjK3wdaLMMsA42nPWkIfr+gCEJMFOMBijrATFBJLAny5xz/dCaRYr7UEf1SbqNRWziQu/S/zbp
Qs4uEPTksoxmGjSy6zcxmGvP7zzV1T9YISnjbARHNYQzPkl0bZk4g14NpNw8b9UotNjR7jNO5cHI
9wHPeoq5G0A+QcsYrkAAIYjHJ2J1FyPZ6Aq/HZfcMfnXOZ3b6emGY7GJCg+z4PMlOxkWDDXh19Pe
wRx/tyxPfS47hDfI1wQbRWLo70wmns1Oz5Wv+1VYCdSWwoyJxkvHHuf1dZinWO/hwLguZSO1eKQJ
RGcP6kW5m8ZKZBntN8jd+Jfv4M9CB5h8oNEv6ZaDaz+vzsDtQw5lI6ZUp3eADFiAxiaGNqSOlo3j
dg1TQEBVMhL1QdqeN7WRtJWegvuQNDTFZ0wJnFhDsjtEryy/HFMv5XdpH509lIzV4QGkTKULmutt
dleQcQsgFMI0Krcg7ITy+yZYSs4t0Sx0r0kJWRYiQnHQUFWk1TGCaBBRZnzKskD1dBxoPThecC39
JJHyg8nyyJLo3y0EjglNF4bpNHoBJG0Powh3u2SYToA9GPt+Uvw4oT3N+VNPuIPjBLA3cB69y5MF
mDQKJzQAroDs0MWBUG1Sodrdz5XWE4Vus7eqCmDr88eL5Z2YFKfCCybPyEXxoMAa8tZiJzAI6+oE
f1D65mUEehcVY5lc7hZwH1+371/xhb9n9Mgp8x2FSE7xdp9q/QoNHtjkXvdwsFTZacUvkuUuwIKV
gZotbtODe+frvesAO3rzbd46qglkXHGKXj+UnyU5CHVQrDXg6gO/1afUIzEz+GvWjEUwTCPr0ddI
VSMGz3PdA6rhoxAelr2lt6ofsdmjQJmG9EyMDn7mLjIdj5etaI6rdYem5Tpmi3vHVGhWMIP0AzKw
Q78lVWaVDs2trSsTM0uET1ajiKoAZLDiI492LFkdcpyM1qh/R5Vu2MNWifDbyeycJwRwatGpULuT
tR1hAr9CFLBq06pcZw/JtVDARBvFzhpz0EjZ479AdrgHz/4gE00B0OzsVLX/OYsJWPq3JZ6ETeGR
PD5n88OZ3LsBI1lgExGb2jOigbj51bmS1XNKp4D7PQTFWVfgJ5UczQjxiiSP+MAbUFMUywjDRaLW
OQTplwiQnUvClTZzz/VoiFcoCyGxO+ZGUKelmE7IWEgef22lm/xHY1PuLFdMGBuQtJCNKOH2hl/w
GnzuGFjmyvDFon0bVMC2yRE4/4XUyteoasNX50fypElHlYhzcFUxQ5MpCUup1utMD4V08EUDWKWj
3/kgNpCWVL7UFpAm3Z0poYhDRSzHPoR2ogeFph8HUnu6/N5Bg+5Bf5vuv7E6sgy79zpwLgCEj/s7
wiRfggxILB/XDaKsoGjGDhjDgftwzUhHBvwhi13yo0m7kJ8bjGROlebGdLMhjw33VtgEY0DT2Xup
E4yKPEkbkPWzByxOPj7+bY/4QxE+GHYzuiDaL9Sq5Q+J3UeKgfs8SYO4RxAKdPZgsBKq4sRCpiqz
wc5PFEY0uFeyvgt6wKseJwexOYxR5yqTMvZxEG/KhyRozDI0lPRMCxYaFBf/2ZM7PE2pgXwr17yK
MLDB0CACrW1y2mt3Aqxnmuc9Fe7kJrSBmQEJ/PHzEw2d+HV89xb1vbeFMZmoqIe7yfOXhW2dRwrW
HCxwgnGoU7kD51cyK/0JYslEiM3bDpZwYfX8msKvzynGv5EZHth2nJOvNzl1rvXx7HJAkepbh1Zk
4mBDcfSlCU/P80o4SN5leCR8O+x3agsI1mEi5LLrrHFVLzqaERCftAJ1nhJm+CSSZzZ7GCDtkh2Q
sEr/3/HkqJ9jUGYDiFDdWArVy/BMNMSB1O3U5puzmu+3YuDLEYqSSEVYDCGPX2gdZJhUtwhmFqTt
OZa4aFZrDQdWNhZ7oh2zkc88dfzg0Cb9x4BahRgejlVzerI9TubJv2olxeGu5CCMmpSf7zea5OOT
Jg+jjFwmJONdQGV+tmbKMvehNNyNNMdrcYkSl3HkUaCob9D/iInBulZoasd3EiKeCDIuYpWPZU73
ec44ORCkRM+Lj6OMaxMH9O0SViNjkD8Q27BcH08dxoUHj2Dg/jXWHEcmWqe9YrYE3PddU22XugW0
ySmoFHRy1B4gx2KphBpPEvmmjTz8wijEU43GqHxHmQg=
`protect end_protected

