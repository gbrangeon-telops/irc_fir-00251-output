

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e5HXux03McEJscFg80ZeuZznrIJptNO1SFQrz1pWkRP7P3QoqpS2mJZRj5k487CXMg1LSvaDqmT2
OL7PFCCTiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hgCd2yd1Ey3kW4Xi8EYui71ziVJlfu+yPA/iSZYYtw01d1xCQQbb29qdxk14t+CL2ulbT/AG/Tph
KVRTNfPiGK79TWiKACghNYtvZsEbOSiWp2tzfhZzsTJKt6Q/Tnk5KS0q9lShCg5S46ZxNmKbnoII
YTwtWH6VQAWKrWw0gQI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tPm67AAwZoJgqE6aGdH3UBgFSYY0hEjWFTT4t/9DwITm8ODgcytWQbTKxugKHOWkwgxnsfouuhwt
QO5L1ilTy6LqSek7CTlbPwPy4k6tJZltW8YhAKZe6X8IJvIcPyG5jVx+6vlxM+WibCk/roITcPkm
9mxr1ZYPG61/YergLsZha0lMNqW4wq3ID24jQg1utjPuifsU4f5hPPbAaCmkiuYhwkMNuj6VHmIU
m/hi3cIAvUetwb+LazrLlZHRjTpygeOmt1PlMgoOOBXow6h7AJvjUUWQmikWL+0eXLxGX1SKnX5+
Op5qf6RZYmh6jR7nN97PHzmxB7CCeLZXWlS7Bw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
as6iakL3FcmLsNV7kgkV+92olQIBIL1+cbziWnl5Jjo3DH55nMZNZI73AcIS3DfwFYnxJCqB2SLa
SuhR2kAcUXkLjAVN6C44hN7PokTEYbZ0O/DrWDwmWxnool0q47JMJkAhu6l9w278iR2KPAv+EoYt
+JQKH1y1F/+RNrZ1eYU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BFKuZqEfqjecGcxpRGmpCDvmWO5m86XHlx1Avi4sYpYvtXIvQdg65YGdV1jpIV3rjwKZHTLGWY/h
WohbbV2nhc+5Ruu6dAeqtH04PeCXz8zphv8vhckLjpwnJT0GWHiaXAcncvq/6wuXR25ASAvhi3Ai
lvDf+vNs8eunn+yE9uSpqndZXDEQrdOREqbbPaHrHScG2A0wHmKCr+QTb2IHKcEfLgWtjt/VCXIv
5krerkdmS143EXlDVZB7mfDSlR6bwswWViVYnH2kDpeepoBCAgyzi+PoFfcxhkn8DGVtdsW89QDd
rLaMLCCjYMVnBfrYxBWw0Bz0mfZcivLyxd+wbg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18544)
`protect data_block
y11IlABj8nIf8zkMHiVxtZfat/jnw+JAL0olRgVyZjPaIoTiNb6cVSPQjBqSlJGLWTwMh5DohjeX
6U7h3+G75T1lWTXE5ppTyOZ64HpmPPvHyjcM2JKGhJ0nO1+2qEF4rkTaV9a9TZM+476yDfRmDl+r
sFdR7YRBqr4BQv5GtkoP6QfasxyaWdlTd0niBCQLLKWfrlY0b4uvXGz2Umh/AIO6e/vt11ecSTxW
fJefDqterS98yAn/xy7Eer6qapdpXd8j6X1q96Qytt70T5wRxmo6W3ZtYicQWO5IHmOBXgkHlo2d
WBM+79u1YuTf50yJ41v716Isg48Ii+2hBL0nh0WoVVaW/b6qLbAU456VIa9oWrNqjulLEWD77N2q
o8bf3oQJVhU8ABrjSvKPB5NcvAt0T+6ZvJCpXZO2/bsCH8R+ISHZ05+KWTWlGVazFJLzYBKZjxH9
6YO1BrVHIxIgSiWtke6jrv3GODKk8/wMFFnB1nzyz+JXswfcflOZoP/hR6GA0zbu55Dw0bY2/q8r
Fo+T43VQ2P3hzuGXTFJWEqyhCOZ+s+jSnOEhlVFtkFEhC1YdGiyIb427PkgbMGNmJoiyCSIXzgOK
vWY39Q584HCiNMWy2Of3QHR5tIH/lZMDnjsZQmniBQ7MkHNM0zwl5CXV6vSHW+RGzGNTrRnZq9yI
DLhgY+o8b9cGiiWr+ExrQfwDOzYM1fu3eswMiSXHIKhsPmfbuH1wLudGyEGuxB2TdCpCVO8iQ2GM
XsJiNiraiU9FX/UVqXaUUlVZjO29rGnATq9NK0+CV453eivDwhEPCvQ3QuvcyPwimRLEDqR6P/Xr
8t69p35tZAZC+0OtWL91dpdwD2gHW0XVJVUacnoyzfiz4ou2aNrQtIhhDqejTlF7JM3kIeigkj/T
WxjChWsPRipHKdA7BX9afNuKL4Hp1FGtvc38yED2bw+8Y4iooPr3h9abidwkRaTAYiZhSmisJlh+
bUlBIPgD0wcgGE7WeJZDvYKG+2w2lH4wWGU5slDLKZcmsB4MjGJT1V1gJrI6haMGzE10QE1eiBJB
BcEwTAKbJ8hWkYhMciyL5P8CLXeNBrhYbZK4ux3CGAv/TPsaoFw1XVugrijOtj9OTUJO81W0iDcC
3uqPW+Zse8Fcf33n8QggHiO0jFLNFI8Kdsyu+h2tTdW57gYEViWv17FQVtB9iaQIkaPzi0P+/cdY
7nNQZTHLkcmCn5HHjFGqj9mGlWqPYjya5kzln5X2BFWneQWPuhxxrRg/rSb5akgs5K0vAbuhVIEf
ACGYABF5/kzyWkBmgCqkUYFjHXM2wWdW6vmloGHBZgPd1OfRkZ6Dsb5cS5RgFlvzIr+pKVptbB0A
WCo3/cbK0P/E03yVgwNVcxwn9egRFRCzOy32eMDmaWLnC30dgi7oUpXUdL/B27lxZHSXg/xXw7j4
/qu6YOdtNxxGJfztUr6K3/bq2nHCRVOW35hfVcc7UPg0v1whZdccY6oB7eTNZ5b2rhr2QAPLz7O4
e+SGqEW72gMqAkx7zG3iOzvyX3Q2B2tu2IdZw13JIzwZbIxfcCyvUGu5tR3v785wb7dVq9usmem5
RrdX1WM5uTm5BUw5n6vz2AOaVDWAeZfvgl4/wDfCxMhkXEZgthJVQonXzZ/fo5eZskKeqot8ODOL
HI9V2n4KY+a2xkzrmP6suASLBjJSgag0uSc+4zokf0s76x7opgRqvsg2RFY/cTbhSt3kggXB2QcX
f3pM8UHLKFIEQsXo6x442iVujkbi4MySeQNs0CbFlukGdrgZuExyzzq5rZD6V7TbbSsILBZoIylM
b5zNwWVg0kSXEiA9K1a1VXaC8pfUWbHheo1Xr57wdhxKaw1Dg5VzZj3WfGGPV//YENzENlTP1J0v
xha4K3PO36GKgJAQ4BAP9ncO57fNbjPz4Za12drutqjGjIZw355aZqK3sr5Wrdcv4SoPcsvfJXBz
Oge0WJvJ1Yyli886AKJcVEbLqFLHMDRa1ilIjbtqdXxyxDe293JXiHToG1BezQhZo+Uy61+tVhxZ
epUKGfDWyRT8zg1KFZ95e6EeySYpIbK8v9fTHhHyz5Wtk4CERFiscnvmW7Vq7vEDzAmjpJAoNEey
GEb63dAHf9C0CT4D/lPCLlWu8rp7oNprN1o1F0kJsdVfnqGgBRMDnpmDsjg3m3KvhVt4Xovun8xS
QjT0HJKw8S86NDLfJYDCLu//qfu1DMWRZJjRzLQwk0/DGutg/G8YEaD6qxRxk/Wcr5ZlgdfpJP+f
mlpVBo75xyPYl9ehhj6OLQgAzzsb3d8MoFNvFoIouXzt2vTVPU/OrB0W7Ln5xjHiqprcPvQvJ23I
pHuhxBV76HL8yde52ns/LsJspRcM6GpXUJIzt3X7OySmCC41Xu1X684W0XfiVH5xzUH/dRQVouvU
qq3IEexHKHv7WidIoAJtuutJXA+m+IlUf/IfrzTxhb7iCMwq9XT3MCizMgUE6wu5RXXb7mTiCrRC
nu/RnxVJaL2cxKwDxcpMCIAPBwcAT/T9wcbXiAr7Jy3J1Brtu/euiJz52CxF4iZHtN9VsHeDGRnW
H9+61XOeSJKLzLSa8CDrjxpm+GAehGyOcj7mYs9B7+9fbw7RWJ6SI+jF8Jh9wibrFWtSPQ7RY/MY
6FHVDe61ZuOW0NwUgtnhSXrTLMJ/VYDC4D1T3yDP4qrWLQdMnRFDtOkdeS0K8zOQ4jKWKpZMcoJx
vzFsEURKlFLYF2ky7PLeZpzgVgtEByQECfhH4+TqduuCZjHoqOCGyoqCnn+n0ffxqcrQ/4x/CRhb
+T9Sp/0nnzYI47zmnXTX4Nnk2BItHni1XJpbAtLTWz0bG9UmGUZoIGfWvn50B9vUdM31lbJWVcmP
ZVCmxNfjYfXXo9LfJRX/ZD31Sqhs+qIVKjW06r9b35dgH8A75osUprGBTBYbJPebaRuPLZIb2zK9
qYpRD+IiKg6FpYrxAE/HbZOq+67JjKd38ABe/LNQx3GP0xb3qW5l/mXDXm5V5zbxO9/VEO9NlK93
rvLwfd35aT5A1O5sd3eT0EQD8J/mFTFoqM39mcNE3/n4Csz+YST5mnyTR3vmJ2CUX6YBLqFbfjH+
HnH/cdIC7uarWtQ8lD9hakwDv9O1tiPmhSeHJPr5kQ86KyN1M9mXjKGvrvZMxAUHPQOpFvQ8D7Hh
WHN4BYP/ZA6o3Z9N3S67EqngG2KphQx93ytDq8C77yZXrvyAkkxBkW6fHEEmH8a6h9Mu8yPohMvN
Etck5K00ffKLdOziNfvbFEZa/wKGKD7cZoymCXRx5kpryEyrcCkY+prEiLy0yuIjj95/0ff5KE5V
R8TE5B2C62oOxKV9SNSNY3VjJJvVjakkOFGWkBffS2RJW8VTiQzjajuvpCaFMCeuFm0MTyg5lRoh
ktzeFvlPF27E1x2tktjffN3YlKFmMR6U+1ddV5DZJgCVlm78NBwDbOf22evHl6vL/iQQthyWNr43
enpVTXbCJsPJ/nBVOWq1b5F+4NM+B0YXUj6DBIf248iktJkKqwZbkmwKGsogfe/YadEi9oczDGsS
akMRer1ywhPXzQ2wexsxxftHOExe21DJJpqQlgu7MNFP/JaL+sJcKfYPUxrMnaObUz1GEXNpKGdL
ncLqHjgflU6n1/Yzpcffjh3lzS+foh27Ih0m+L4mzsUbc8h8DB6CLT7YuDU2/IHtXX/0DM1EHtlX
gPvTxTOV3g5A8X1tI6vF6lv+XGFlZhGIjZFKvqzizswp3QSPa6gozbvMIMi5E9PNwsfl7kvBpHtk
il4R2yLr4oEWAe1T+P9bi7SJemrcqq2viPrxyV5rhGlc7V3AXaWosf1lRvxdFbPyHg8a+I4PRgld
cQvKsJZ2xBP68krbs7WplGXYKtWqCsuiB1ivhNgJbsM3by9P5E7rbOIr/8AUacGvQuasL+BQ0GjA
5YuiqIRZjNIgGeBkQh7JoDCd+DFHq4AYsTFhHL6Y3+ZFwlSmjfIyF6G/o5QC1f8FTSTAXnq7Q2al
YvjXSzy6upBoRixBGi3dU4jcRmotO8I1I7zm6rV2HbWEYQWZKLM8OdGkwPPnNx4158y+q7UWh4Dl
YQvKZOmecM06ywLyQ9l6teFMngQ+ra2z0KjYK8eqva1G9CEt3N0qfAb1gpCS3O9OwHIY7qEGzDcK
OocsAAU48v9n7GRdvtDQcvggjB9GIBQvwJT7B1Ok5mfWutXeSg54vnuTpSTumMc62GVgnPacvqI9
HEkq+HOu2OjsEiEJ+sa/WdJ1O5nCg0+7oHjTTNikTW7ok4fUCRvSPq7YJoL1nQBAZtJ334HzHubo
WHFWiVIBxDuO4dnhcu4LNYaunezclnAPmnZjWw48ViMVAkln9ASCt+/6+hsWqpwq3468sku75EGU
VyQSUqMZZistCiE6SSwP/o5A/N7P2d4kKXLAJn2UAQzGB/Xw3CrXltAXlfJp9TugjmIqjGKLrZIw
7ogIYUNMbLqLmcCDq1+2U6IhhFoMwmkIAs9qAehRRdCZdONinkZ6+5ap8astMOmX32Qnl/751AGL
qBrkwsUqzLFQUVdWoRJz4kiePGYdlfJdzr+KdowajqjvKoBJ4g4EahawI4XPQJ2tggArRwgeFc9U
Q5GKKglR5p6K3aJNxGWmpt/iKA1vk23INbmSD9Buyk6ugEnJa91XVBVV+/l/RBsnBood94d2yUMi
4yAlDeiQOfDSwhUnOn4toELY1ecpfMRWRa2eBsdp78Pdo4/xF228y4+x3/EM38BG1R+o7xN/8O17
guYUTA+oAMJsInVVJF87Nj7Vs7QqSRDLVwomt17dy/Oa9Ssyrjxkm2r0Io6dOqtVKIhIIhUf4vKH
fEx0bublMc1SiTCYg3pLuTh8mm+t7bFStldbxLlza+ujm0zhYu2p4W+cHGJbo7D19oT5wnLhrqld
xXNcOB0w+7dqxtXKKIjNTuxF+7l57Ye1Vi/qVnk546d2MlSg5pO0x4zvYTyg0iPpuPicKgYedtXA
VdrbmUzraC21+lVooGSHkxCSNZfqPfiu/O4+3yWX1R1/K2c3rFOCUsgjEhY+fzfCxAm7SynE0EUW
XRYkybYs63ixYXQNnDhP78/VUz0Oo70wf94vuLo08bznHyWZ3X7AntfKQ8aar1eg7QMIqQj9msK1
TISMT13MX6L+OQ/YL5VvjSzUoblUWDGGSE2QYzcyk4org1igYjEpWmf+UvTyMTTBngZUeVBCSUvZ
R0XAt0fw+9Xc1UBjhkJxj9Nj8r6KLSmof+hgyhjBcEauvwn1QV5qUda0AokMmzxofTvjZS3MUWiC
0w61nMBVVcdPsFVBfeZWPxhl9nPb+ddfYqsa01EMlD1oe1zVHdR7ps6LP6Ad7mMJVSsYza0rLYD2
kXelfLLatXNmDBJ6FB4Wu4ZqbmhxHf9hCwO/7OWs+uYAUIilc8gmsavhSjAoGGDzUgqjZAcxKsnF
+L0mECTDybDV1KxFQm5GWFudrqrR39nKkJN1HSvvv35UVtDHzp+NU/O8JQwHjwdRzezOwBozLAu+
Z3aiHiT6hoRrEEm8gK0EpLvrL3zFhaq0Pa0+/ABpPEzYVdar3+WAw9Jbnmmsq8cRNXRcpF7YuFFZ
YWQpVX/onKaJVGpDHjVqIZIJ2TZJqTWbTyR6Bvw13+4JSP9qrWChuzf5qef2aOJ9F4kwdbSzu5Gi
sRyX1CIjtvb2BTn09zDQHwixBeIjZ5FCae0gSaEmFJYicl3FWEfSCp9l5V610cASMjFbOtBY+REJ
s4ckQFoYqLQo6iWLvw7/pG/XuCaf4pZTQDbtq0jJkXHkVXHphEkkBJJBh4EbnCH8LtRkgJQXF1yp
vOuaCnlpEVJ2Y4WA9uQd0cEiG08QGz7/mRiXEMBcZe26YIJwTlspty06+lmrKR0bU8LtlPcoHKlb
qnFkJ/dmRm8SXibs9Z6YJc+ijJQcasBvavks00pLIYfMTLqFIwpR9Le655NPrwvsEagUczoOEdq7
A7Mxd5IynIKqr2or2Km/0bjsoQ83TQhlEKpYukvzrHcJEeDu7RQoY/uQ5kjVP6QNk9FQKvzDEDzC
kX7x7QUKpTsgH8Sa4SAVUPweaUI858jBm286XDdmi6Bo1hj1GDm1T6sH+9LmNzbdRhWoLvMvJ+/m
xJW/QOcZUDQsXOMX1f1rIRqWBIGeSjZN9C8anz6nJQRTFH1v+j9O25WaI9MFs0hvOeQ+q3lUjufh
1SsEmvXt9czhTOZPTKca13KZ5Nq3GcZM4RV1nhsyjBfMuWhvf7ZJOa6qZ+8juiLFnJB9Kx8WZ2ux
SQxt/bIKhFNRQ8vuomcQuq678Pr6mIYo0imTNFuQ6V76FgA8VfVM/amKenJbCclRy2cPjnSryYJX
QW1iZF7Q7IVnaR0AIOcej1+Y2lBVQ8sOz8GHqUG4HReLUx53kk0f5kecxLdMqDt61JyV9A1rRLkP
rzOMRMjlQ+CiBIhPKhmU6Ouu/fDE1B3ZlxFCOcx+zl8M6ZusxcSV67kG4Znm5rITmlkpGqtQydwW
ev3iIYOO6irFe0oWc7hqMmex2f6AsdDTl9CB9NdMHwDcjmIluqlwuqxRTRiwSE2sqXQzJvtsFR7Q
MelbljQr8B/Kbw2f6qe9QpE4cCdds7Cg/+Uk6oZR5twTRYs+JMmv6xCw2cqglzWSEDm01tqL4LCI
ACgDbw/mK4fM7ae1t5lWn9VjZ7d9gHtmtjTSW0ayLVltcwviNGM3inBIInzYPv2Feqxl0RYG4oUl
da5uUXPicOGA+6vKPgZvRFt9TbkS12kN/ncSkcK4Cqej2JorGZBkaCIqBQWpVLhyBFf7buLTVysN
0rbk7oL3nguM1N9Kbwi8ccOsmrSlcARu9rDrNaeb9H4ik5WajzTliOzlJUpSyO++Ne/qYRpf5Gcy
jIF4zyUbIUDGE1P4BjcCokoiL2TFRm1wGL5sT8oEMHdpLXv2x1wrSobL3B8pL+IlVii87m8Mi3un
onO2kU89SG6rKdp9ZajDBVhzbuCc4xZBMiT2P0vs5eH+Rr+QHu85lW002n3fdmClvg3iKz46Ho5S
rYX3hSbjoFV8cTqWdYyYnyWeyXsZyo4qaPJa172g0jq/BIoJuVXVKvnLiteYn+5vlXsYRyX1XB5l
r2t4bq/wZGI4heAhry0lH7BqU71mcY3Eolh+ntbgvB48iUTZTxj+n8TdenvqC8zZ4qpFY2uGmqNB
4COGZ+u+gyn/tEUPrTq+RlZ0LPVuUbWsqEn2Byk0IiNDKX/r0sF1UjG1oJQyyiRvvJIf2vaRF+1Q
bE7302BoVicywblRPPjVfpPX3d88pzeL4jIopDk7UdhRqQQTZh7+ab+ClHKWCvE6Z6idHaVWu8pE
3VFMEn5UDevdwF9MPbCCohf1PCRuT+6+3LD3MmDzqjoLuyHYdR2St0Bg0SrFtrwfgxcf8Jm65lwp
iFmhxn0gUY9oUb0V0nxnt9IlTuXw/LAiPwcIkuGVH0RfrcDbRRqEGVeoEbjCpC8QrLS7fFJUCWXA
G9eEr9k6G/+eMOLC3ydFFhJTTO4FSIJzjWg0VlS32AjN6bQ42HUpj0zyRl/BftYgQ7H7N3SQH+gs
4g56ki6GZQ8/tfUIJLhA0GUKPT/GfSErf2yo7btheWrZmpY1Bi3tk+TKx+4npH1x3ryvBaAfX7Ha
6ZDx4NvgB3AxSYlOuSWmqHIPx0AcuvVVYJ6QMIGiprMmEGUE1j2BEYAAzv51fYgMBSbOuVkqqvMj
O8Dyikp+Amlqj5ZpDPE3TUHURevz4vdHeSIDl8rVi7T9S47o2MyP70XLr3suCcaKgFqJjygSCM72
Nwz3ji/uw9B2puF59ov9iaExx1mC6ZKuGItU2xbGJesRS3S33kuddtGA+Xxjc4gWj++dlOm8fjB3
W+UXinMN/c/F7cP7PKTnCZvOs7HO1hmKhiCAmEcXtOwhBV30yoFlUdDmdyCrxQDyHwzBpBJY8pNA
Mqvxrt4wT8hIaj0O7n/hJIhutXx+wJYkRjYSsFDAIZv89PsL2Cg9jXcU7GeeaxgQNJr5WUvn1MvN
wv3PHAtHZUXGr7+Zby7Z/2LfcQbsdRVGVKzYKY+pf61onw3etfS2471CpVMlZaTiODVzF6BhDlYw
4Ey6br5J4uo2t0HaZmwj8qG9v3WDrr5cnip3tbf/aXKhnpbd9vLUV0CfI40p19io2+leCu7di745
y6Cxrl+6Y5iJTrtimSFl9z9yFNOlMDannDtzYueUAfbfinrUz/IPXnkY64EZpeIOaVajJaE3IL73
+NcjGSO92ACxNPNvC/KWg44NbBwceVieuCeYZSGioafY/IWUTe+PYkdGbVOu1kXMU9bgV5VrgJ0S
jcaTkCecm4GSHogXLZ+KLuUup6noYy6lKhHfZOrUPaakyBQLUmZqNB6lZrahECkuKb3rE5lABf6o
nzB6n6TcMPtGRaXOzGHayI4/FMFy5fNbEDRkoqc9+3TNDTpjbf4EW8ifuKBf9HN3IcHmd3XHxyFW
QB6Ajfkwx8w/rRk/Mte9on0QGgePUUAIm9z8QHvl7ZPV09MIK5GR03l8AHUHcyBrE+KYY4Pyx6K2
HAxLYm9QDY7/+S8U+9zijpufgV7CtMeA5XErVZfbMUK7yzVaxE5gfMP755DJ2kqEgT3AL7srkXQk
AYInoWzxSRHXmqD5KUnxzIaqPg1FdysRglW8hZf9GcimRlQsrYCvZhXT4GNsH5yqnMubxdBnQpxk
PZN8TJJc4o6hOVVsGtC98P/oMDLzC6WzBWzHNSz6kH5OxthuTtrgwz9rqaOIDNWm5hAlZ0v1Rrut
6xWKwjAsCT/37/iAq6hgsxYgo2tRKDKMOaO4+Nmax95/MAdHWn69G1iyZUZ6/3wf8/shaapr09WF
7JvFaj7SzmbCupBcyz29Ic5W16ufgIzLRmYoZuGqhgToPrPeCDNYnzGNxEDwFpZKjmEYLTRlaH8w
9FICasxmk1sWw/Z5xJpUJuBPLQNmczF9s1i4i8mPEL23vzYSYeqgFIOodG9TkxyAcvNrXZ0IDlMI
9zOxUIbO0NLd4uQexEkEdGMHrKYDClYm1UwSBWhR61lAhX0zX1k56lWl2jwPYqQb4YXWJY20pBnf
1Pnq0bRuUDjA6bAJCD0+HMXjNSzlRvXktOcs4ktqwXWbH7C/67CtUtKVAMQZlZ8Qm5IwmD8QKDhk
CShZgvixs9Czh02bAf8Ed56rnRydrJDpbd5ylnbyuIfxRivXJjpyPYAAm+IwuBPEXYB0CXTNeVy1
p/koAT3by+bK7jIL1+LwYO5BbM7J227T5e0F1lOJ0fHUo8hwVUl43nCaKJxXIK/PoTRY+wxj6Tgl
snHTQFkrH2cerlheLHnT94x5dLZsamNlZdLciXHTJkZesFuOdETKnzGK0zBM56QcKhiL6AnNxeSI
ip5EaktTZD/V/XlWtsiUxsKg3A614V6U8c/9k38DsU2K9q+CmxQYvCVk2tQpoyaHKo0aUDL5VUh2
gohJvYaDFygO5H3fCcfBHHqgU0EGP6CDdEA3dfIW/Hk1Ie84ycTH+hAUXmPhOQZn6/nLtL67C9eO
WoOVetpK3QVak+uS3/EuelgF/TFKPxzAdaMCvNgWFiew/27lHEpznMnLkOxlyWoRG89DjKDCIjfY
/B8DCU4ia+tPQxHzvOa8l/vgHBkjaR4q3qaOcw6U4u8KWrbNl5DLt0ynzpH3Gn5d1bLChXLqf4uz
mV6RL072wHf1NE9kBMzagME0hjh85nWokwzieMFfeedZA6wdr6Fnaf27kdEOEe4enhkOoQxzTSEA
X9M23eBCZXZCkbLyN5qqhpPvPxyzDLoecbrS4MT4tZ+V/nQ3JqA2gxwqLHX8ZKnjRrf15vr5uPiE
isCyq9ZDEs0wD1GBBNJ52kktlb0yFMPvjeAaKMwXLBzV2NKtlPCswEjBGchvnX3W4SmnK+682sfq
4ijvrQsfVPfpD+fcxm4VZYk1ga+9uwur1QY4NpeulR+SQ/7UQ3QEswTIKrh1wkOE2d8yOcmFH7nn
/4dTQsLJXR07F9v+7a6gMEJev/MRugV9hhdxqjHnGiFlnUEWPfSSXbWDIaKS+PtN2r9/SRTWyOWn
3CrGY0KwqS8Sp/piE0W6jaH2KVQuhUWSS4U50xTc3W+4b67eh0KKiWJ7NMXTzZHfvfvTamCy1z9U
1LAgkhlFfc0fZz6sq3iBtfTGCZ1wl4q+VsVka8hpyhd0jDzUNVfOitJ1PpkI4ceVBwU8HAaOtj5y
9kyTQygVoHHwkbvPq/DFiJKSL137oLv8bAyGpjpmbNhnLqWo3aWAmsSrCKUyiKhRnf9vrDrtxV7x
BdxZrJuPkCWDS7A+0PzMkW6pqOmguDDwZSN8DugR9FeK8DDsvbImZvRZA3aj66NCR4Nw5Al3x1c7
zNbhupdLIWO0KOFfQC74w5ANvuWNNFhxkI+r1aLThGv8LMtA+G7LvLLNUo56rObzHaPtlfV8X6oR
4jpWgIOum/nloWlX0grW8hboAINI4DqUnxCqS2pJBg5yHCTXAH3JS6ulGTbVZPfmxb5vVmBJQD7K
AL9Mri5uhLgtpggDmcCphgGroJKIPyJzcKDvTNmzZXp+2R3JKiFqJWqI0LLyMWKw+vzMRGG378Dj
53JKzthe2sXW2tKOA2+lY4S0RauJq/+LcAMgDfqb0f2ngy/bWY9gEstNUaMmpZsVD6jDQzcGEnjY
ySM/aF+j6BmFp4UB6/fqfjh/Um6/f+8Sjhxjw5oJJxIACMiqdhWUI0Ore9+yTfAPU+sDDnK7eEN1
O6EDjGSk+lZvkd6t7vkqFq+e+TePPl8Gu82BV33YNWW71v8B7CNWaEQaWVstdeqZ31+og7pV/wE3
wMG/iuhOQEEFCPzczYG5VrC+C4Il+mdNu8BtogVJ0NtrX3Z10ppP0gkKav1WpaaZoi2N1N4BoFiV
XwwNxAkxqBPqCUWh16/Q08JtycLeyhF+G94m7Iq4prXQyyBdDacmnBrbxZa8C0Jv+kLW7N+2GD4I
vZkWdcF6Nl+u9DKFOYIDBneLpFQr6u3QV8yYLno9slxVr9ydqGkjOBbLL3KJK3fOuaoy3AYYdIjw
AYa8lB5ipXPiQ8dmA8oeS7AUxUD99SxEibwSYzTqSw5n+jpMFoAvwTRjes3zWbzrcvDD+6JLbsbj
eLx3oo593hJqBXbV/l5UnVDCIawYOiTaYdmKubnZnufruGUTSGcNklFBu2smfV/cUIy8BQRBtPJL
0E05wMOTswv1V+dV4H6o6nYPgGFMkMjk/MuF+vXOaxhfkvH46lxPd/e3s9aeQXUDCr33duA4ains
XHCNxehF/iFzWcQDF4u1xv62eYJo1bhzheHKrIblnypyqMSwFRQ+pRBbxGfa+1s5UUAU9NMYSJbX
S60Z6ylVDKIVKotKo+NaWFG7pbA84OtTtwsOKZhNea5eg5OmBs2WnDY0zWBoo8l0kkh852FuhaVK
mlGj4FxFltvME7z1VFzRjEBoj6rIgBFgp5vYXLX97J0MFVRreb88AUhzg9VZxo/x0m2W+q1AgCE+
Ywzcj8ectiIvQePCUMNcP3O+LP1MlQaFab+lHD6248XIu+0bbt68pVltTNojhbwaUYBh8WQlC4uj
BhUcg8ArXA0+yVYlOghwu/WmJQDMO1GShX16R6X91LDMOpFgRjzIOUXxilCmmAqTj5K+woQFTTE0
jC/f5H2LcXFcZWFEv1fdnn1XowcO3R1+QfoA9iIBsXzSarVjv6tYzOsqRfuCwy1XDBRHTYL5+jUb
pmaa6RTtKtZ8lYXcu7ZRDMXglnBTrzyZipBfUk0XaNDsys+dexKKrstJ+7gUoNM/lRhy162bruZG
ALiRDDrrPKCwk3aKTY1mUVveAYKSZCM6vMh+NXUIGXLEjeec3joqlY6oQu972Vt0op+FR4kLrrP2
rzm/qQxz0K/SA6lKmTdmkWa2IuUutaN1mhX8nWZ23zRZKzkWwHughMjx51ZzZiGqDECOraQ3VX5K
Nr2xr1q3ijKL4ttj2j4+2b1dlJIf6rE1dvCYwy4qlPPlELjUib6jeN4tAUKgyT8Xp2PZhrfKamuI
ui2xw9Tqg0GcINqu4aCKKLF81ofXs/3Foz4ZzLafnX9KrLz2fJWDijNi/TZbCG3GWHj+PbupbQMZ
7Gu9YEpYubzcI2vtut9UyNTnuyZN4LZv7px75nDSPyLyaOf7a6iSkgxxunPjPX3EdStvkW6ke1IJ
iX/y0b7amqPUhuGFuDSQCttHHGYSR+GX8ZHGVSXrUv/l8GpNe4vjay3HDt2ehGzuWEgEjVGGrOe8
FdPOxI2s8YpAlAbVPJPdLV1y4zjDchaenZUQ/8qxusgxyIEyG8pWPIFzSY5/HCgFBMMvydEixzf1
hvXM/geqxjmg2zoRpouHJAACbV0sHjCRwzO8aVfD3CntX/rcV5FAeh71MpW8f1WLISiUf4KyL/Oo
zCoJwff6/NprwSJxz92ovt7bMoDu+sdV6Evb5LYV6Y9fiOpoQ+g0XSMX8gerlyOcnTyu1iKbt/5x
wLpmGLft/cS9RifR1n6oWcwvNqUg2BAhbbrwQzVGYlOH4cDWL57NIN5e6jCqObThBuMDDILdaaOt
3J3efUxu+gv9/Y5bK9NyNEEGl9sWvCtl1WRzspPYCC3IS2Dl/eNfZ8cAgY9Dm4d0NYqJSfEzZULV
fP+/1VcYkbvhIZHdFOT/e9yqZPXlelaqTCwgtY6AFkYQS1lSixEM0pua5P8DSRJzmoUPTmejRw34
ItyT+vGxkpswBbYOZVyLpr38QNCAeOGgmNXHpQ3bymbZndowty4A5nSnImogJSIF7vYD4mvYM4Sg
y42OdHLP6U+k4dITIir7F4qSNomuAGVCOK3DP8fvld2TFh3jkIvtMhBY6WV3nHMmvYFEDHfNay4u
D+cPWUFiiWLZOhHeGHrOH01d5WYYOLiiywDKhEquKfl33w7fPTvA1LsKTIlHaphd4A5z5uzk2lgz
yDBplBoP4VyyC1STQ+BM0+bDnf09D+IOpeMtH10DXTzIxlwzDHx0vcq46AiNdc0A1Jz67ZJYONA4
SOYJk+R6RJT4BSGFqGemv8eHmQk5YCrS6xuUCe4SUefmcKGSVKBt4tl5DaXDcvdn2DdvXEa+L8NI
b8cvcm9zWLugm9oWvLuGS6kLvPpuptJcCt6ZT1F5xn+8UxLZXf3etXs4b+6ZOcD3ml9ayckgFHte
qiHsoWFzmaAVfBHJl9I4lDDoKjp19TjoJbVJe/zHqbG8UZIsQUj2nVX/QkX+4dpFxQuncgN7ablC
CfvxOySsjq2zXVGzgKkBlxsJyJXvM30qwyFRyZ7nB3b5BtEGVIBaYUwS7TnX5hSF2xX7UjnbT4K9
FxWtL7fq4CGj90GNgj+/q/hnzuYOGHqkqwUIzkMhqHlYwmIhWycZFNBKri8PzGRh7O+umKBKI+iu
bR0aMEaDoL6oh6LnzJD5ue32knngdwMQ3uAggP9IhEbJesljBQfzApfJazBTEx8wMGiPLpsjVMkI
tGJMqHhjI3PFlhXa8VibZU9sm9EGnWtY5Ttf5BsXBoGcZA94mZ99C96q294tHe7KWadDCwxrqtdQ
i/4acN5K6F3B+yzXbnPmyv3URYAtTKOVmzY8uj0HOLugGACB/VUy+PL0HklF7Oh1lpK5JAJyviKb
oZDDmGKJm56SArmio+Iw8ST3xDyrsh//Ro4cXPOx9ssDkK1/rMErfhfR92tVveqMVpvRCVtIkTBP
v1WpyfefjmWu4mHPvzm3vqis4vyl42GgwU+4quUrg/L6MtYuGwdzjGyh3ZdjJmYLP5SRsmP/gxfW
dQSn3hH5uLP7B4EWcVFvyns7SxbEFF8/5jVijSHBW0nUEXfFN8NVj07+mKScLJUW2pc+Q6e87dHB
qRcHU+63bWZ5MRjVNbNIEBGEcj3t5u7cvQXj6yCgxVKRB6TrZ8+mi0UwnFNkZQF+auzM8UhiRz2Z
oOXJY8RuSCHMcc4j9RJVOAXBbqkr+fak/6fUwmhltZlZWpe4pnsdZ5xrQ3Cxahq2tvzD5lT9+trO
02o8rQUcDA09u5ACTDpTCXrVpZyCSplvEWoPXvoLWjM13ydpwDG5Aayfqkr1wAswvr+H2R8NoRfK
EjomjxUXOH59OSxYXowT+lRxh3hCBF3UNQKez8N+60Br+UAHYofPdEWe48+/KspUyK//kYL9ocGp
qDrlwxfbl7J3CGR4Dh7r/mT0vsVwjOJMnLKvoodGUAfRe/dG5Fuuyqk6IEXC9/QyUOlLrelH9gdM
P38yj6Coeyt9IHShVR1Cpdvi/jV0fioxRvd13ZAn+sNgoJ5+8CMV1llBZbudzp7VlpOTDdmEZg4W
py3o/ZPpM5jNlbsVR52exDBEuRUDLBpUk5EzLoBAHgSzBkhJeLqzts+WZCfraI8l5kT7eh4WA3dK
gIrx3/ICJrf0l+WW6MWmHKb5df4daEBTevMamyiuNowFRW5M9JwhuoP17x3KOm2DnlPAem/AS4GU
Vjs1kUCpRJszDT0GMW8KB7mQ8nheOLGsL65lh7T9TXxL2GYX9NCXT5YpI0QzrZtsYQqloOmDznZE
xvh+74u9YHhoKjwCP5Nrex1CutuSARq3gcJWRhzZjlQAwRsutmo40pyGSwi8IP0ROk67rqWruTT7
4gSTsxoLyYNY7YvngxLT8/zDcIjeFyr3NDFj75GAtAPJvHOUnlRulNqpXXVUz4vyLPLTFjxedJo9
4o77EEa41CmEJi47s+Flflw6hQbcDphM/9RMFiBqiqeJ1GJGwTaBpP3XM8RAW+Sn0tl5TPyOr8Qw
L3+4BvXSshqO2PMFbVWs3lyNL9yoQQffyrnqcxdvykk/EzYpRoVzWjqtGVJBYMBXho7C66AxBkmh
fRIAiP0JzyDIj/9jies6hHwr5B0t4Zz9sCN6f4RnFisKCv8JX91YpcjYyuDsbm89wQrhOnun6Reo
gzQp8XSikLzdbGrIt0uzoP5o4dRT+tQoJUgvjhMQByS6nKVstfenMo+urwlFNWZ2N+EGB7zVr7sv
a0xiK4bUPEDltMGNR6A2t1Fd9jsbIvFuQ5AJrI/sYBCCuSNauzB9fgKVwaKivOsEnn9JkL/vkYy0
CC1/gBfugXPiPYe4fC653kD6UXL5I/fFV6zxRjwBptmYj/+/MwoI1CGD7k9HDbrmgQonOz4qIWhU
nNP0oABikyTOZ1/uxmbS+Z+ciiqN3WzttcutloPn31HQZ1xFRzYcmUOfTmOAdMj4n65RL0NEJWjc
YElczMq6s52THvXH4vMzjBd1/RaT5pYHcd/N0A1yInoEot8EOsb4fRkkJrz7Opqgzy4dEGjrPgXI
VIxWG14MhvYPoVtwvHT2ybh4yVHpWAvl8d6AyBput6IN9c/N3AwdxKFv/dEfBdZt2/YdESwZA6Wd
+C0MkdevxwNwEHAGYkCxcEJS3zz267ZYhmDG5Rf1WxCQXmS61GdvO+kzofRVc5OyYMeTxx5NyPFC
yy5fnrfjM0iWBfikHwF6Luow87fDdC8PFoeZZAZTRJlxRpH854SyjJUXbCj+h8nZIkeaIpbHiAxT
HewtiU93DuIz/Cso3Pjgshl/1SExNdgI3fHaV0ck0dckRXEoDpU3UOkWwIx8L849RcHiwwts/Oxz
46Okn+kyVQOOIATAoo/uR9iyL0zGh/5KIeT+5mKlcglZ2492R0Knqq+0isUmrsfp+4UsH5BLdhRb
HL9EAKo1WY3g5b7eAkDRI/FYwzWmB8Yfm9rmdlQRX3IZUniSkSvahnHueY6E0NzQgN1wsvnItG2o
NrDmMH+mvQelehcT8dbM0TIoyNUlpxeT78EHpycl5cdKlMDIDclAk+xkjlQBiwSBYoVNWYIEPGFT
RjNVUWvRDqzwIiUX3V5eMAspZPSlzhRar74jsM4TKLNSCicJGGYtv5x37mpb+bCnwiQP4R/fkqP6
NcA/XVy7r7WsBC3MbLcRaCJQoLwCDGe41ZE0BVayP2YOWBEn/q34KFxrtFvVFBs7GGxLCYwpx3jv
Fn4nnQIf/A6yvv9PYsgtkJ2fIn5KLc/fxtvkIbrlNV7zLUvWILc1nHP2IOHxRY64Yr/VZ+Imi1sF
MxQ66WvSbA9sfzh+LXs22dS9lITIzTEUTDfCM4yJMt4EPknfZO2G4/LUROiBoCsQ1voqab3uxrdp
xhiUR/zZM+LjKoqV9haGE3DoWc4Kwm4nKMQJI7KrA7g0+/9iCmx7Hy8ajUnahqiSX0jSmXwz8Fp9
ByKZ33hh+yUpUBf2ISIVP7p97yHi/U3Gf3tbSNcUxKcRPW6csKJSdMKtzlfeXajjOADjQ9o8YKjo
MFww7tFduQwZtN2m0wAP03ynWZSCxN+Ua0RgCQnhtiJ7YfAceAl+zI/WL2cVcVvehwXncOa/uUlX
D6zeXrOg+EBITbH7QWSbfckB9mTQW/H14+fUI8oQxoM1goB7VYBOFIy+yClur2I5iSxOxAj/uLWM
U0uz/E4vnF0kxdqEHFn2nK9hoHMm/6IiAI9MUBdVVTdcbjR52EgnbllcfmumvRtMawGpueeDaY1b
en01QNOeZmNbzlkuFLdhaZXpjaFXORPf8qsbaEKUnsDTgzKtMKcJSjfdSJhMRYRI0tLxZUDHJoXu
sekozigc8Y5IanCr+hl8zu8txKbMXckmtisGOQHaKweZOfA1nDT/MZtALSL+0YrEPIHKHIbe4W9U
8DdNQmQNC79lwwKWWYpAtOznqGU6jOeDvppf+q0dSrbDS2pYv7lmD/L1qKYzrmwQOfHW4j6aC6CG
dfMUvcYbqS/IZB2Qohbq7qOr94BwXETnuTJuILjbDUMMRbZNp0l5QF6A5AyocK3iDKFL5OQyiyHj
To/WTvf1rPrKB4/JpxL3jENrIwo13YtTJ/ifuO1Nz3e3ummHUUUnDgRl+cF2+LiUS6VDEJW1TQDM
9WfLpDXbbt7ujvAhlHCXyc18L9mwJP8Pjby6bjTpH+qfd2/whVya2vQFucu/vnPSJ5kOa4DpGiQK
+PdGjOfF6IJHLN7xmC/jwvnjElmmjypRJwaTJLnCo6WOrPryRMCLiGacQFTi+4JZndie7DAlO8fu
thcN/+R1ko4XkY+C4My+vWz4FxBOB6cPzj32m1754v0XgpKmwL443Uf1qd7i/hMS52M3gLJKUrEe
frS+zeSfe2ILa7ehpwpW8XI2/GNDYfEYBhzy8sb6n1RebcmNGczKlTwfNbDOaiT/iOpSMpGt451g
tXyZxveOONtsOjBdYdxjO9N3NtToiUYJZ2hqhoZMriVVIdlXovnUwPMVDFKhCEFRmx1MHahrITgH
DYIAl3IOVi1MaQ76A/zKzZaGOkXlWGeQo+if1XoVF8YDeCYzUSvJa35jBKfi1yUh1mlX8jpeRL0I
22LT4Kl1SFvbyTltFmrAsnsCdA+vDI6ImHCukTIk/YjHAGMzztOvRAjMNB39k/O4KUe6tBaZvDU/
vSgmNXFFluCMgK0NZia3qAqcY5nbedPXtSQOm2x1blWvNz9p/hOnhBn4ly6nDwEOA8HSxbVljslW
uDLP/Bo+Hg5FXmty9vDX05Q1MeHaXL0sW6/fy5HgOkMCGxCC0feS8Xe/R6n3lTGa3ncp0XCwU/4a
tZS3mMd7UB0mRlquDHB4lC3U5ZQKvn6Ij6/4r/ygxU5g9zC3dyCif/Df2s6mrMGaMOVBAKL+kzvx
cuEAYunNdreSG3huPPQEYarDQI+M4iSYKDWS+pj12R/6xrH1X2cRw80UV/4+9tMXcoXEWuk2yrBZ
T5RZZPtDBOw+bSeSvl0pgx92sn0m+yLWUcDaTmfaePl5FOHTEvN7JMQofFJTmoo1bA/wDFDdfRxq
JU8n/GZG1pVPB41ORU/k+GX3Fz1tG1nhNmOG3AHm0Wjm2dTpd5FMl1JX9/JWuYQjJGTkVO/yw/7w
Sa8doB0FdikpkRtaIscbGGpVbRxG8gGLPOc/GEhPqh4EX4jlGMPHZkPeX7qY7ma95jlYnd/jXcTA
Pp+hX5ChNUjmfcjxb1GHlUhb7vY5o6dIcJPQEdEwkMjed3yzIEjhu7AQgpOO7dn5KKLmdlOY0EMX
1zDfyioPxVn5Zl0R1wfjEF1NBFgftrE0OoXSfVg0tIOUq+KeF/4KUGif7+srZzpnggQF+G8N+YqC
xsqZASv9QRlkxsv/X+/U9QcPrCnHlz984ILWcgv1d/8xZ0RJx0uIrnfrorvgdww8rrvzKNxNrrOT
pQxI5Xyhq+3qqVADxnZ5rCyJIdSu7utikblMsHTeuH5WlXmmkk+IOK6oZZRZpQl5uTf49ndiJTf8
77Gud3JoG61RASFayDimoJyYP0B+VOoqUNCQQ0b/iJX9ZUR+tZaSK1B03Ox/Ve21xIGAd/DTqhON
/PGf6aZf4tSkyUeZmygG0hFGTuiOvws4rMWvuYtCkgX5s2Q/dCp6P3lL0TXq6wzhIxANLpubNQgy
ZHhkITV/ntPVJYuhwNXU4v/FYA872yMWJWHnoiv9IBEV72vXMLSEn1GK2JgGqfiTZL0+IpcWn064
+JmowswP+kmYK4HExw+gd4KPktq1dc5Ur0NnrvUSu4J4s8jGNESpUeEWtC/iSxPI+4wkf9HvzM5g
uXGl3hm4mgEKlibOpJC4M3CvWuKnrbgfnszYcMKwaPC9LfPfCMOFdrDx8mFE7m5EbWd/5ZJZv+Ic
eJzcOmIfUmaN1iBEofgRSgwjo8/eOeQ3r8pdgBvBFx+VQzlZSJvsCiyalLC1kixDPlpj5SzG0jS7
3IldoYKYgrphh3QhjlFd7E2H8vOMYKrLpYosOExp/kGfuzDAJonjr1K1+1mG+0o6wnVgjsjvPCpO
cjm4YUWw9HGFUydNHD1okei/CfiEuvwojGLxNgFmkTXtAh6+2vGDBr8dFR6IyEfvN+ErBRkGsDH4
lx8IPtno9uPIpjz74VduzLS+HL6c+52e/nkuXsBWHUUcF1hUUfge0Hll3O7XdP511UwRwH8xubNL
NZxkczuuFMjtx1MpRBcGyegjXcYmpwz3JcCqikKvMLC6qGUowTuJjK+beY8LfPci6hlzwHZIA878
kPZDp5WCkyi+//2k5z5Qyt+ZzErwozKyaGDAqwUftJEWUh2tUM3kqYxT3BESPrLKpeJkfxySz9aJ
kDb785rMlgVEJyPdKf5PUDsQj/UiEj3Rbc9bBUHl5x3Grpvp80gxs+NgzGBzvx00j9YzDho11wZ5
1y6j+903O2M95tQXDsdygMFlBsnAGJZfmuACeCEez1EWcFiGDIyGXc0qFQ6OM0qGgDXi4yqkJ+RN
ytHb9+hXLciRMgQiHZby3Phn2HA8thmYdN5HVBIKOGKjLYndUnnO5DKH8gfSEcM4AvVEjmu7DnUH
GMFgk0B8IeJMamvSpFdwUZyh2WEiOv9Fe0TN8Rx9zdKG2qROWNZJ2wjs3fY1wEcDtD5F4UsGM2n1
EdjyyaU30Ci6cIbs7vsmWMOeCLpCSWh+MAUqHF7B3FFXKGQvyAaFIxuqtQdS5/SVUY2HNHkLiiog
XWqHPTSKFPUuGiiwKsM3oPtVIkJLQFILINNCzDBbzl4dLjKlFACwmj8nmVxHj+y37vGWayq261l4
Vrl38CnBTVIpO/jb3Mj/BsRZ4qSjI5aE/Gub2xkrRQvNPKOVv3IQcAV565hqFY3PtNlFrzC3BSJS
Hfc9Jx4pcWptSJuXrIRDKpB3LBcan5EjvgwpqPcZ3ky55l6kUZOY8jY/zcLyzchzxCoEFIfHcdqI
qZlOedXvtxW46OYRgZKBqpGFt2dvd30EzEUM9bAR+aC9WlBZhjb7iqP7TG+RNosL3C4RdcKIQf9+
j8ugGLYIKLJn4GjFgEUUHlfRLZnHcnnds3QlzOzHBKufQ9hPYXY9Ao6kS8lVKfZNgVexJenF/U7D
QtFjL/Q8qsmCmSNtODFXpMBG/SbeeeTxXwqZsr8Ofer8d2aaql1pKKMJ4qZLB61shgapKaHXRSkD
FC6MQaqHV0cB1es1VtHxYVzIbiaO56hBPUdeugI3KqrOHR8G7iZh1gKeW7J6YNA7IWOAkvDWWc+6
DuVA17ME1NxX8TnVb+vrX12qQe7qsUOVGQ3PxlP7gFkJUTpKa1eT8Lx+fmGovvtFXIAvA+HdhAHM
A0WrVcttXMFMkIxVeeRXhmtKLiW+gAoCJ8jA3AVDuQ55YzF7ZLU3O4i4qXwpma8YEuoTJ+z8hMH6
6kQIlUtsP6bmjTcytKZJlG+JdlIRaNqhBvEAcXEkdSvWCfxaLObGGFkbnQCsPvBtk/ff4LPG5a9l
eEPqm+7RFTMfTA+d26EDv1+XmLPDJTpLFQkvzVsrFH3D4Ej68IZ4jCgbq6HG3m/9IVtgef+bLxgw
lOWFLRsTWjS9LyKnNeDRriDB1C6HfTuXwjI7KQO7MTCI7eWRoiYgUxdS/SHuouxr6sJpR6oXRiRG
0DMwu7m5XTt4ThSxv7NualPV+pHUupCsaZPceq2nOg+Kl1C5e5VyhSEZMM/smIZUNLzeweL8cxWG
ttsnwgn0L5NWqYddvdkeAKsp+EoWXGWqXIemjKt3CkH//QdAIZ5RhB40yjWNJfimmr1//JQfuK3w
Knwy+nOP/yHxYaLDoYE0Gf75WxVT8LvsYwoQMDYiy5FQjVWZD76lYhtn6XO0zWtq+xNy4GXyzx5m
Wr0InOyXbaRm4WJqw84x3EY+MgB3xP3uyT/8YUWe02tZnddDwWHf9KbnB76NVp53RmctgrVBqTsx
Kgg3ib/3dOa9mXdW/lNNPUWPCIko1xsEy5KRmes6hHzEuIxgr7hFSV7rG0fkmbedHinnNIYDiJdo
TeRaFouc1ardH5+kAau5urpZamz0nUMIsOTmPFkREXeXGFx1/1BrsFZJgE0HaMVeyunx8yie0GFK
CQ7qiBiHrhklqI7dBxnteOAVj3it40z2dO34qahSbW2HdhApjEmWZHAviqjlFTzcwhxapye7jssZ
CMMdzSq34vJS1FDHlBjaGMT1KBJDL7qsKS1LNCBPKKiIFcmTgglOv4ym+aqJ67tIC/+CqZsXWZ55
Z2NeFCagN6PCsoC46+FvokGbkHvnRm3PklGf8b4sTt+JBjuooyiRq1XZUWPuqZig0mQ+DcOsqQoo
pjyH558IQ62g82BSnAzWRX+RznUx++RvrraMWCdi7JROezLgy2PzS9dEWFql94q2DUy4QOHSsILO
/wNDrUP2ZXgJ8f8sOJbnUhHiWLwMaOtc0X1RaRVGbKagAXmlvo4ImWxujP12zDH8vN2iYy0S8ud7
HSCQApkBQip79j9xRi71JWpZJMSQ0vYBXsF5BOdjTg2r/MD2HAINoIA83CibpLOKmwA3zb2N4gRF
JZDzymzmB1DnlptFbT0iKSdwxqFnE2Wx1nC5Q8qGmxrcqr0GOEDTsUTduhVIpC9gvogPivAKFzDJ
Ekv6C7qtwmM02T5M4hgMrOrXZfp8/vMmlY/qgu0DVHQ2n3EjsEl3eDfbVL1s8RrX9aUR0YZDfoHS
ScmblbuJjO5VTBjTpJBSV1kopvMURJEMjDcAbGfkCt4gFSlqLMIDacjIHGcmJW/0NqQd/2QwacFC
z9jlR2GtRRUN2t/N17o/6zbu7/z9F96D7Pd44FB6DzyYzX9bzSAPzsiPsIHPR4l3zrRVtYpykO7F
hVDRp1hpwfiKsJaAZz5SURZie8nkNLKZgJlJWKjVWmWklM6IiwABpf+zeh6uzFHAyOC16bSPNOJo
35O3vs7KYqgwytDzvS+UbsQ70ipMglKR6naG9nNbhfwCPUcOWPzTbiXA/6BIaVpLh+ZbJIyKJ1Db
Qw4igU41p0Ud5plpHnrZ+qcYOx212b+IbrNYiX2wWIij64WsNxKUHSdsX4GiUV9pCvIEdHE85RLl
4jgAxvxepWL7HvHvw8enEyn47yz89xZRILGAl+Mi2VMJcaGDjliL6x1ScKhUdv22hNZ8/+5f4HkO
ZuFJWE1y0oy8Tvfg1D5WEMkE1D9g2LmNghQJijNpm4x/TEuz1lWASDTbuyDt7A8z/YZ7H9alTIOn
Sy/t7J9S8CSJ+PoQcGC2U6kvwmgDxJOrPeYKDmNWF+if5os8FDWeXV7X0035gts47eQg7m8SPUOt
5DwcAvRCf4dvN/8SPZu+brkVu53EcgxjEe3tzCiBTq/OLORpHHBjPhyaNcypNUr+AD5/6PsI1fkl
OwBIfXArQKslNovF9aYPqxQXd2T8+TWbqpI5BmGImSsuLHNZgQwxWqN9tUuI5Hyq0Vcl7CYkfW+Z
sez8iEyNJrdthewY0/9Et/kti7dHGnS/TeJgZVM0GKfFlkAl4QgkpxHYKlvY7FApwqpCSMlEXSy2
ObtwPuna1Kiv5nAW89ywTIv/qlFSzergyfPax1slHYFQ2y/bseMFSzIDe7xf4M8LQyjde7ed193x
ZHFnwL/mOf/Kb2Zr6u/IEpGsYpDX1XH9TKFShECVQABHoDg97OlXysm6fy9ltNzpPIj3HM7FqgxF
6jcnzcpqO5lSX06LVBlWlPOLwy61usyerrdWZaUpzw+/C9B8Kvrs9virxx9AUT4x/VlclDNi7VC9
/dCjtcIE1N5SdCg/AK1jiamZt6P1KiTo2opiKsYdS9PX/CTLQcRCyL2Zf8a52bAYwXZ84xekdQPj
gkEZe5Jhuajm5Uv63QcilY9P9XBB6lMFfKzjAONZi2JhRjP4T5HTc6kXwsY6uw22MS9GhwgzpEIk
RWfZ/DCV4QO8ZdX+fY9xUiufzEGfEwrScPzWcKd4d62ETldFQd8YYeNbMCnR/eDzUrdMaF1M0KIW
7cmi38woO4VwIGUpdvsjWfSHm7bGfeYiYX3SVWS6f/yaTYJLnU4UtpjSYnjqLQbYAtZoO/hr6YBK
IZKR9eMJHcYArboq2Ciux3VSGyXV7PO7nzDAvP0qYLebHPQZI3PlHHg5sEYRE3Z3oELbKBvbuiOO
4OcThWNMhADWzwpgAafGrs45RlDjyo2WWwuEyUwv31fK31R1TRHfL9cvDPsd8WQ6I77RmIwl4x/m
MG5vNJO7qo/YrnbrFgvzLjxlc+BXYTvtbJTv7ARlOrBGOLACh2ONJSi0QXFvYYL/DZvd+PlT3y7j
gPyRaDFztwgZEcaLYeaKFGl1M5Wq0dl6mUXQjBCkWpmesW0Iqc3tVCzNwsdQWySpvG7AsntYC+/p
JG8Yw+fGMzpiX7dVSmai582/MuwYNd7Pm3WtOC6AAXj2blPcHqSBiFn/3BD3Rm4e7Js5Xgmi4xN4
2uW2y+Q2uayAOgiXp4mCrp3ilUes2J2L7PILBMeTLEqsm8fM9rVBqIe0R3TtnkwDGOIdkVtBmB55
TaCjrVoT/Iyk2HO11RqpLDE2lLcekWc631LeWtkhBopY0nCP7cVwvcj/RzH6crQKTZAY+63mwJaT
qPaH8PB2mtzInV3OZ4e0Y9nvGICdC9mFw/cElZ8nBzR2ZrRkIdK5TXzVEx0gbEyEsRyZ0n1j/tMv
FJWrq78R29rTf5xMm/Ly6EQWLzCjER0dtTcI/+nGB8MG6ythfdcI/3UoHzqizhrVnEEZc+KNgU24
xDJdfUuVPVSjO/aVWMuhu06HlZJ20c56x3CcHZJhsE8WVM1eDVOOMOFq9tyN0wGfjgTM8EDB3r6L
g7zaxxTW5oTGiG6DJYrjZxjAUdqg/VCBgS3ZEpawtXCQhppQj9Ta1ZaIey4hEk4beo0hAfdIeJWR
yWobj6/FXwGilcNP06giZm0jZ3B8ejo/Kp/22jiID/qco67coNN1GG3BqXvLnq973KtQAYg7SiC1
9ZXzb7WDmj3+KOB2FJxiQYoIt4Bs+3DYK+YewG3MB2eUCuZ6eHPY2FRm/JDqelG+GM7NAiufoZ19
LzH1FN4Y47ykITgfvOuxLcLOeSvVDRBXb7Fq786TM4EWmDxyd41cs5IVd3C22GeFLcECiPt29BF3
ODaor+/eC85pypPnPbqniyf8n7CSa3xhtRFrkZiX0ycKhf0mIzo0v6k9pAHO1pLYqOQ1+fQLUWCh
/uy9s07Qled3TekmlzAOpM1PV0+RYdYWEiRB2Ixne3vtY7Fl0Ej3EO77KLSs1AA5qpyaEgvIcwM3
Kp2yyyNVEe4ZJsuZ1yLdWg7cfHpMI57tpMf5G2/awgSF2XJJELUOC3UL49tqSdYmA60WuIfYtvnf
IUcJAIqHRqYrLL6LSPWJBBFQ+mv++Pjf2ZR/7cG+YB14TRk2AnT4SinKsbIHTfKVeNjLavg20FE7
S1zA56J7kmvMePh3h9cIGOOLNmGl0Vke9enXlnPQ/cBBRLYu6A2RI64QKYT6qRJEum6sEQ8miRJr
YffyTA0j2kcl367T7PbFZRkY/M7h7uZrbgIDcx7EuLqQKIPXvSVIyvtpXfA0u8yVhyGemU2tthee
aPt1wUBYFjPK9INnPEvWZ7+nEjBXgR7hBbsUZZhgb7tcSWBQw64NKiFbzGpUZbCKTyEnSTIdo0IF
Zdd9zblWhaoWEEi4TCUa4tbpQxHulpMSKTOqzTfTcA+YFL/DtAVhpNq76JzIdP7uR2rbyPRUpGZ8
hNmV/jZX7oMKsQocewIeXJ81dtGo87mu8Csj8DxepoArfwWtTYudz6FhJAcq/K/TXZWhVh5MRuhL
WgSmdzPxctk6i0kk/CSCUQmIVsDon088tgm147FN6mql3VMMsBUWhxoaP/iJx2p9Xd3CSB8Q/zHM
qE3dvok8TQowaiiPo+flxhrOpA==
`protect end_protected

