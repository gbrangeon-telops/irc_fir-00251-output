

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e5HXux03McEJscFg80ZeuZznrIJptNO1SFQrz1pWkRP7P3QoqpS2mJZRj5k487CXMg1LSvaDqmT2
OL7PFCCTiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hgCd2yd1Ey3kW4Xi8EYui71ziVJlfu+yPA/iSZYYtw01d1xCQQbb29qdxk14t+CL2ulbT/AG/Tph
KVRTNfPiGK79TWiKACghNYtvZsEbOSiWp2tzfhZzsTJKt6Q/Tnk5KS0q9lShCg5S46ZxNmKbnoII
YTwtWH6VQAWKrWw0gQI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tPm67AAwZoJgqE6aGdH3UBgFSYY0hEjWFTT4t/9DwITm8ODgcytWQbTKxugKHOWkwgxnsfouuhwt
QO5L1ilTy6LqSek7CTlbPwPy4k6tJZltW8YhAKZe6X8IJvIcPyG5jVx+6vlxM+WibCk/roITcPkm
9mxr1ZYPG61/YergLsZha0lMNqW4wq3ID24jQg1utjPuifsU4f5hPPbAaCmkiuYhwkMNuj6VHmIU
m/hi3cIAvUetwb+LazrLlZHRjTpygeOmt1PlMgoOOBXow6h7AJvjUUWQmikWL+0eXLxGX1SKnX5+
Op5qf6RZYmh6jR7nN97PHzmxB7CCeLZXWlS7Bw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
as6iakL3FcmLsNV7kgkV+92olQIBIL1+cbziWnl5Jjo3DH55nMZNZI73AcIS3DfwFYnxJCqB2SLa
SuhR2kAcUXkLjAVN6C44hN7PokTEYbZ0O/DrWDwmWxnool0q47JMJkAhu6l9w278iR2KPAv+EoYt
+JQKH1y1F/+RNrZ1eYU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BFKuZqEfqjecGcxpRGmpCDvmWO5m86XHlx1Avi4sYpYvtXIvQdg65YGdV1jpIV3rjwKZHTLGWY/h
WohbbV2nhc+5Ruu6dAeqtH04PeCXz8zphv8vhckLjpwnJT0GWHiaXAcncvq/6wuXR25ASAvhi3Ai
lvDf+vNs8eunn+yE9uSpqndZXDEQrdOREqbbPaHrHScG2A0wHmKCr+QTb2IHKcEfLgWtjt/VCXIv
5krerkdmS143EXlDVZB7mfDSlR6bwswWViVYnH2kDpeepoBCAgyzi+PoFfcxhkn8DGVtdsW89QDd
rLaMLCCjYMVnBfrYxBWw0Bz0mfZcivLyxd+wbg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18544)
`protect data_block
qWgnwEzx6WhSwmURuYm31oNGhuaFLMwqPArHk3Cv5B9TSjF66I6raNOO3a4t5u2+HoK55O/KKXFv
+LTHVaO0w8t5q+sJKAh34rPbr3iMeH/CTgLoMJ7a14fjf8zVkYz+/u+NryDzRsTr8ZJrgyxMgE1w
pFM/oiS6Tw4r6zd8YR0kEPxWQVWVs7AhHmUoJwVoHRhYWjQdoR3IxI+CICL5JxfXQO8MZtE6Tq0O
tHmW+1SyicMWciKEgyW7uQ+uHj+LgHj65mO7ENuhV+6rNl0Q2ZoNxln8GkHE/Q94KlCuLN1f+Tw0
IqV7f3OvEtunQDdrXhbiJ3/mDYC3YJ6S5JNr/9m9DL5FqZfQuWgV6XIa1j5kYg5UIRtGotCXhiOQ
Qw75AjmzfEvNWwnSwuk2mOlVFRj/UmcjKbsO2++0vR0nh1WqJ8ic0fdevwvw5LzYjzGxs4ijrdvi
lSVN5cQwqiyupNx9FOfVWhAa/Utif8M0/nHAtSVTkCeMHMvV0gQiWcpPt1/KQEd+6sxny7v2MuhL
KllsQNQdGb9u8xBuj2lcPfrcbQwY0yzFSs9UHm08BLzzQ5XyxdeSz/iGLy0Er2ujJXi7cwEshb88
8mjq7qi8MFx1UcLK/gNYE1TJRubQybL9C+zjrUQ/mjd/oXM9dPjuwtU4MHfOLBgAfc3xol/miu8q
196jjYUOqQ4Psi0JN8IENgKN1q7nDBS27o2xcHHa67qBkICNrYGDPhidlKv5X2Gf5IS5VszF11RU
kK2yhr8jAWye9OSvMVx/C9ZzY9RhFwaNGLiJeewswWG/4lkMVjWytQ7JIh/vRTrIxZ2AYnDRyZXS
IxpVAmi0Z4S6b/3QDqgsYbVnExAsxc81NJMEh4k7Qm1spS2dcBy2NlLsJ7r5kPJrYPl0qpHFgh7s
EATW3il8Qb8BnUuL0D9OPzxen8+q0E0axa+t12aGRWAaannval1LigbqGD8XbqEEbt8cDLoWJzj0
ZdLa72yWf60YSktqxCjU8XQqhdJN532uTKFmvkXVVuyCnCkU7EUNt/4jPcUFsZhmSLx+EzzezRbY
rBw1yfGCiPHdSOHRT+iY5Zx5dE2mo7hNbJDHIhaSa9Nv1v0JFrD7bOjIftp9fhCd0YEjXjp9C2OV
1BQnZfpY24Hd10DDAFIMks58+ejB4QpOkxhv7P9XQ13F3qCJoKQk6voRcKP6vALUFG0WNG8mVAOS
d9p2upia4m1LQbqM+NWGc+bonp9Jwg3tkHgFU87pnrkmEyrIt0RUsc4BQt/97DNvukWc8BYJ83bd
Hpio25xjrw1yx0Ol15wBWwt9Yg/GYlrBjPEkiT+dK1OgiwbR1U2ErUo5IP/IcqEHoaPvq8BW3yrc
OrL04C4SSzGyolvtT7yvBAZUSTYmmmm6KEamUyZBwuQlPKJ6RxKR/OidsPnzLf/OOP7u3l18RbOI
UhgpplhWdqSQ8meBqJTY3U4rsfRLGLBt0DiiSIPNTx2u+rZZ6EJUWqcrtlI7slFVUUdTcIYtXKaK
KWmeOXnnSuejFq3M1LJVWiv5qy3MjdmyHIl22jHVftB5GycQ0DPozTqPYRuuxEhZs0QNzoSDb1BG
j5hR8AgMvqDc3j/CgMkx2rwS4BOiWaSxrYeywuQK4t2kl15ZChHwV9KC2ngnp24In4xgBl4eQmYH
IGGGXw+UwyKwDUlNVcTI/nKB4HiUfRQU3B/0FbRviVEWP626e1FsjvERDqoHcsnCBNJIDgpFQxiD
kDbDllt95i3118Bb0QDhjCyc2eTBu4gwGqqM1Nnc+YaJeeVhN+epACg1MWA+RlJNDhROwjfgZtwe
IlV2b/80GcZ6VEIunPgWHIKKsE9v3Y66bDjBz+JbUcG3lQ5CsoEqQXkvfsz38dIaR+I51q0Sd8DZ
WutN60d3cgSmkAH6musd5WHMBJ8VFxNcyUOYkgclfBEji1MCy3yhXQw8hm9nCOkVNqsg4AAPTH5c
j6puC+e1rs2XhlV4DuzyE6iBol3cpa3hON8XMMnaROKHgSjg//+5uLpHNlEsTei028XQk+LeM4SF
ykapNE3u4cO8V3OcwR0UUuWljXwY0v/uFi0ieGI+6fTljrZXzkiDtB1+WDjV4PJE8pWuMJZ/MYWB
p4Lw0pBx2DAn62xGcaYT3uIwBP8hrseVe+KFY1Q8c+CkHitFHa/3+mszoD9Lmw/sdasoIUn2WuwZ
y/lpO2Ad2GLFz4PjscwttHwA2hfhbD3KVsgfvXDl7fNV8nkE6d5xvVBdEZ6kwVU4fre8MUeGME2u
ciJBv1YmFeFHKLJy2bkV25IFVkz/gRCO7NQOmLiLGP+l1sejPn6jBzsS2iexuYV4HbWQanvoAyPm
lIif2rTz6LwseAhBfkpI5oasg6dq1Vu7IX+cBarYkT2P4cJKcDnWfsVnhny1X3Rkf0CY9fJPbxol
1z0/ds44/+CjGnCVGqKzAYVBylu9jR6By6rE1eFguncJiJWe6tQ25Hjh3mOCgl2Dt0+QEoSZul8H
FPygRhQv2VB6kxSi8xnUGIKmfRQT54XqUZ2hGmpsTx9jptZZups5rhj+/qQuhWH/txFmt0dt4Dbj
qNgd9UsFiWMHU5Y57aKBIMDFT5MAM1epNUD+Km9joz8N0oWECvo37fUthfUI73eDoXUL7DJpIRIr
cueJIH7B2AHAWnPcx/iPT6aaVJHIIu+HkenUuuTfFCvNdmlFfW+rNla+CwMXqZ+O69VPG72fOoKO
DQWYiIAuJ+r6eRe2kN+RmF7G4YteOvVkFem11qzD6fshbfWZ7cgy+6av0o8rE3gZsepmJgNkpw2+
55+vqAhyDwzOUJH1lVYH3R/59E2ytATz5IUHhJ2y2OmMLNH5WDH0vY7bSgjPvEd70wbMD5nX4Wp5
Ke1O4u0WizhrHD9IFiWqnEK+8+7amGNzfmQGDTP9onb5anKEkok6NHeOmU+A36xxUATMHpaPKpjc
Tt9GNzqX/G0boOxQLr4iWcFOf0zmn7tx+zy3f4ci0uXytr/TsGrAFRR9Iuk9x55xdij7WEi97kOO
UJfvRWYzJ5kETnrAGPqbGqV0UYBa4eIdy9BFM1EQsLIeIszXlz75xu5w3fbEox5NNnlw10ocISkl
146ZO6n36vaKAqqU9no4paLdISglCqKeeKD2+8cm+HsEsCvOJyVeAuZ+V87Y/+NzVtNszvlPC+X0
3MEghfj6uZ2v+QdWg50Gc81jM/uf5DZiYv3yWGfwV6hL65wEMVVJxY3op5POxNfmIryhqCoQ7zGu
jkluoXojc2IZucPjKS2oHRQ+UGlZsXamFEBPktwseDV6a9aklCFmaGgpEHec3pHGE0y8NLa0tbWl
2hQmDdWjxbhDrXrF+fUFm+hVIvX0BwIsnnfFggrIpXYLBpDrO+7sMyTZvGrJEGjnqFw9KFZ9MUAz
lXAtijKsU9bLgGeLsbiYPhQsiMA03zE6NbaRUbyKAmm2oKTN9JYGFjSqSycTe2WJI4+rJQI3NhX1
Z20m3ql36bdEcAO+POTSGo4ioM1tz3AxdyuEcQ+IfHpwSvAFFTSyn+V6jEW85G6X8XuWjpxiDcLS
zJ6FkrxW9YDzN3EwDsT6wWAu4pKQT50E/1Fk0iDxAqT9nZho6zrtuW4sQR46kWt4r2K49DGFQv5l
aGlsw8toOE4b9K34aVQPWiIqf6mfllG1oT/kftFFJGmzoqW5RFqWjmYco0nthfSQj6oxizvHXX85
4snD4OrdggzDoRZSyPEay1bshLDACw4P9USO2XS6c3Oz/D8uH1QCOMZmkEOQHo/UzWinl2O6TbS3
umaeFnE/PGgu+GSkQ77D65lpn3cjVSfCgFFwIl1FGs4rJEHvo4srlapBgp0OiVlBaSbSUyN9uEzA
wqUEPODMRNGRpWNFpFXQt9iotln6t7MLBvHx81Tb4W3T5fRee8nuD6lua0DSRbTPxXtgzcwFg9+l
L/vV6jsQqiUNWiTi14svxBCvrDKABevrAaMRJKX3povUt7cWo4vf1FMSMfzzDnzTxD6LWXr7Z4zu
lw7QQPDFcxbR8G3i1WZum7t0dagKPs+RfKFn8Vsvj1BINURW2Tq7hGCZiLVVTdF2x+opbH6RrXme
/qswnn/e/ZRKJ0q8hfhPSMwngmnc66aG5qXUPP06XHDyVfeW+ZGnxgXXDsNTplysbhC1Np5x8lkc
0HCmqmXmzqz+BGTvYxSIDJR58CuQLLeNknm3LyOVGcmQQmILPp0e1Qx/PO1+KH34Lxaj8+5qtZpC
Rajn5MYI2Vnq2uXnz76tnnMGlIfGQTaVXf6lB33GSpohwnrdacqDL4FnnDy1cRGVoWu4ffs0Oy9K
0qso2h7ctdRwMAHZbpFhoZjaeabMaLIvfDQl6jwj2C7kLwcmvvxQ70y9UfwfSwy1AXDSvCp8kTBs
NL+OXvup5d1WaBNCjM/G4wWU944Qk97MWvTM3SPyiGxJCK2hH+XIoC2hRQVNJDgcv9+S70OMU78G
N1T+FrSLs7LRG54q4qQ7Ki7bZIv/3HSgz5lNaImRxHneNPX+U2nTg5dNiuBVQDrJr05cZ3GmznDf
pvs4Zo57louP23eGQrRup3aq7FIk8myFnKqLun2QS2aFbHsS/UqCiwileJsMmRQ/D1s6SpwU8LYO
iPHSh+L2fkB3W1Nn8edMydvant4wRjRYxwWgHUhNuigAvYNksCGZpIZP5uu/5ycXy/rwpBQHob1n
5nxhPLOhcrpebTzlexNiTgNoWYoNs/LEeRHFg9OrsjujI2AdE/QF0CJOv6RW+9jOXXP/2gL/7QC0
xdFdL6lyX9V//wdphTr7UF9cBbZAGNrGb6aE94R6DREM/PTJ74bKgnnG7gjuga5QhvxPQjgJFf41
WDIbTobsJeRckhfnQlVaQpM0MeeebYbMgBJQLWbLy2sufcXxYDPIEg5Zy5dS66FrLbGniEkdPalh
k2PvlzoQyfpYcv9p7if4Z33WIJK1Gpv9JVl/BJB6M2L5CtiLjWehwXZTggZtKjy8m8YygnTMmnNL
+Y594i7t091c8x5YQknWiYqmiFdfoCh2sbEw9aFO1MWxT8RFhbFWOWrrYBy0Qlqa3fMPDBq0fYIT
KKH6ZiH1vLsk6+jyP+CIwF/nhqcSXn+3xN/6Nzpn14IyXUI3/oEFfGERyu7UyhtZxvNEWjQz2xNw
qjJzPCGxyIUaEjV6G3GLjoJ2V9eoZw+Rz1Oo5I/6j7NjQmZxEhzMy7h8WgJjgAyI7G65kN+JBwWO
jjc6SnW2SSSxpOtdj5w9VOm3rjR0LNkJbTWQGD12WpsJEqRXkep3gezYOzXTUKYdigzgf39tTzVs
ziCpt+DRS1f3ufLtA+SuYkgWNf638R7IuSS+mZ/FCM7HhspLW1oDbchRtOoG43hnvTM8rQRvbx5m
JUyMb3yRX7JbWaK/amcuMLtYM7c1Qbhcx/IozU/dy8ysROrRFIlEIXRgq+rucsbGvKFXE5ybWdoM
cZX62rKCKziFMpEFGnOCye198u2or2TbuKy3D/Vy6njuYODpYeyy5myQBEzVhN/cEVO0olqwKK/p
to7RWpzgWJ+FOto4d1DUUzUYsE0OntgdjWufFbL9En0VmpQJd9Z1wFStwEci/CyDftdu4k+7iXL9
pX7zAoxDd50Rv1PfP5kP1I8yHYfr82WnBDnwcq4isqyW+7bg4neU3H9R1ZWgJJMGY8qAwGaGUm9X
9sTeVkXlY+3j2OdxG0fts4w9F2yOpS0M7eeKgAoAhhGaxsf2kFbOZPeIW5K8mfoK//i0oJJPBb+W
n5sAG3gnxQDMvVas7C7dbJ9UaIy9uAj+KiZriq+DBGq6Y60qu5pFNVg46w/5f3w6lLmZ9n4/aK59
vKYYMBtC2Au8k7D0oPCn4BN7rAluOCHr14d8huJmLW8KQxI319EVpHswdLECapCqCqUqEKAmzn64
qX1gECTxqKxuZfAVnjeHr+a10xNJ/qy7+dgW4o+SnpvjSPdPPmSmSC81cmfykm0Gyfk2e0FCMvlt
hpZ7hHQlnwSS+YdprdavkP4LTEv//nK2ccip+dkS4oOf3rEZHNQgKckupQ4nRNKf12s1rP5jYy+h
gIldqh07BD8CrdmqSX1EDTebVh9k4vYgwdtGw4ssC1L8OcVNukA/CA3TmhYjqibFo06rc48RynaT
pNoDYxhby1ao3cQM2JkGDG1DxUmMhC75msiWbrB5udyLgVz4CSP92Z+bxB2ITvUCHq4OOhlxoGuG
kAfA9CvP2x0xx0anV+UosThq35KAK2hzqPM62pane5RCK3ZP+ELzsDvOXG9SawUlFwhbTzsXuJzZ
Kkrf/rpp47FtRO0VlX1IiE7pRbFuFG5CDOUvsKqgCIKR2tLVusYlIsW74KP8ZnMmsL0ejGLuDjjz
JMusYBdL+cjXzJ2v9K35xVvYdre0iSILoW7hAzPZoVbXXDm89umUyX/pcZhhKY8SY64ZKgw2wZ9o
4jF68e7/wrP5nBVc/dYMb70ZEkOfKF2MpRMAuZoWdH1+K6c5iRb1pVlqOq96Lz1bRQItihxvAO4l
r9SkEcG8xwHuokc/Su3tkWWI+fwoLESndOHeqCeGpGPzh5H+7yqpeAuC9Gd5DST0eKePanSNfnIz
h4B3aTReZPllSxojgtp5RonSI0wry8cnanQFIDtiY/fqbQm9RcM/DS60Ki2sMMXMTOBu15ik7Uyy
9ns8umLFfOkL5noDoYcNKZH9IUjxMz1eruT/gfgVezfaUZo6WApAf2qcxa4vW5aXjGI2MwjLTMZH
3Y4JecggEPbMouRqTvGVMKQw7gq86EXC3DgldTlZeB2LCqHAaGaD9K2UCHMm5MiaKkZBwEuFB0RT
G2DXEUf6RTm2vECw1Jf6XSzIxMTvecCxjig2wUCl4zRqPhQFvgpr4s8Id8ia0B6id/pCg1GXrKpD
fXbyIH/TRUzplTvQ104SgP574TN4oiqJrD8r6IdcldeX0LvPWITnZovka6E/Ft0bTn+vg0KPNVR4
B0wGQy1d6MjQ0YhrsjbqfPDDbuDoeH/e+XH03hiDLcq4UeHsPqthlkh7LsVas0eMbZIUqD/komM/
EEYPW9jmg/261y4JlYHxfyFJUXroHmD/kdxVg8krcI3srFNES1H7WexkFBj6KomAQFjq/UhXD0ez
maWjoYHMahwZTbx5cgH9xPMlUrftIgBqJuL1XQi+m1oYJB18NngW91zLGhxPzBuPJmEOEwWkwwjF
QiTjCAnZD5LYogVZ1gQJvloggFyjeu75H7vgtuRzBT0dZWJgazyaMiJ5inu4EmSqufpttezj5X+M
GRPVG40l6vs/G2qVFOuot813NdaOvo7JbX/vWmqTkznLhPJE0JaLhItQdVSIlug7JHnzZNpHzUGG
o+T36SnZwhc2Q0cqJ22ULCn4JvlOwnYKMs92krjR3+hLtSJfUzItnoFkhQmGyDxTNnZXOKT+InwH
J04BThYz4ig5qzAtudwyaFvqYGI1+cbXIcOHAXIJ7fNpL9FX0vxT+RDcD04eTboxxKfErcfKQIYz
PS586FaxtUQb7GgWzPn1fqiy95Q3JKqvjXaACS5NNRxGQJIrQtqGFuJKXMXt3uCI1Qm1kzwlvEsa
uBF+je7+CVTaaV32HTJhuYHMpojwX7kWDt6rkWh/e2Nn2OWy29edq2Xxaf4v3Sz/0SQBm2Q+G/Bg
vSqTVo7gw4URst4Z9S9eINpcQ+xZODWfyDr5Gfnar+09GIUIbWw3jW4r/Q66/3gQEILpKtj5o/aQ
kIiJYk6+1ZMKrG9ocGWtPAxKqA5eixhp7mU1XJIz0EKgYLkfwgEiInyKwlRGoxdjTbp6H8bH3iiy
pV9QbQr93qUr8qSqEzA8Ku7JD4wyJvSACel0MrB+Eg/XE0liWzfs2sej6xRExwRVpyaYizk3/JqO
4p9oBAx2IcD4t6xrFHpiJolM0vfotc5i2/mF15WpYYAQ79Y8diS1XhlgYH+TgTW63TOPuW37CIsy
VgEBuYAPqKhpY1PQ45eHPrB+vu4cPHzn+yp3d16vYCO/juyhQ2phMcjqwuHGvtYYQ1MJSDj42IUR
TcijCrhTugIyHXwe6oLhSyqRfyBSq+CIfN6kZJAdARG19mXpkkKrpKPJQFbBeaaXrDKgW9cXefRu
KzkVsLaCw6q/BdGs5ILPDP3PvtJfV3Oz5go9hnxFWftjmq0161Yaoy78xclJaZzzbirTttum1xeB
R+1Pmu7PvV0V1FmEAVTL1jcnNHgQR+vHvqQAcaF+ZGtnTEmKkQrDIiVSY2acsDnjR2emwIBaXII2
8IdsaHldWTbLHt5rVAp7/hQTG6m5DYJyJajCpv8diAN/CGOHttnVtLOA70uPh1EWDFkIXepYvzpc
vl0Cl3g3NVcZV/JMD0TS1DjGQt/8Cusl87ItrktAqbbkH9hmNL2e4qWfXa6IMfmFMP7RFWO+HXWr
qlNheUItEuQOL/DJf5UkedUVt/C5Z4iU9t5C2fdjCBs5Pjjt4m8JnHiXukuWITdTSF/Eg8KU1QJr
e7fTlq+VlZwjA35ldL693HaUl/LUl0kCejlw9VmkKC83uk/eWi9Ppb6lGrQPaiWiWlNps9DMt7n3
L5wDKmy5olZBLCQL2SjlMqduU7jDmVK8OJ6hQS7l8NUJf93ORF7KmFyz/NG0zxA1bgp1tYEq1DC1
SYBAEsUQHZZXYMqymCAySAsNEae7VhZdUsSCXvyJ3aZNssnjU1MGHq6whOUqccHJXdBLDLJQDzQU
GuvvvPkK7F3brM88+QMRK9KrXnLRZos9PnVkVZumgU/ordz69/Xa9/wHTdJyuCDUL48WH9DczWzF
qJJczsauR6CdvekhQbJUaLR3yyuLn/1tq4EWiCt42/emmzenU62ENzRc9RhMdnZ4LwpdhdntQ/T0
SwOO/JGtM//KJXYhJbLa0OIZcZlw0h52iR51jk6Z0rwkhtJWKPL5UYXtVvxrcEQt1f+5wG/iv0ey
vLOCpYytC4CjN4QKNtixwe/vfoqVcEsNWOOI6P/09D0UTrk1Rl+GMW2Xu1hODXCd2Hxego3n7E/R
mzdHQ1JAGIvGawDH+zIvKkIga+D3exSt/cZkLwzPV3Y1YlDw0kYJGlYoDX3YHLH7LUWcP8luss6y
JyMssjX5i69KukJ4fN5PGWMAP8Vhp2mSWCBOK46spWA2qCEJ+S1FK+5u54QKEBBM2FGLsYEuBf1Y
pO7dW7L7z+EtIfO1+3bmkAdFcdqC9YOVnUn3ZBKURlDAPGFR1n0O9jtjhiVwSjC4aHu2fG2sXKen
/i53e7suz/wbYSPmmzKv9l7K/TEI4UuWKr05A1pf3i6KEKi9AIx+Ng89oioZb4P0IuJnPO17y/F8
CisiuBUJaHSoiSMM97pFNqO0dWKFXsQdNtq4EIj/bGepnCwJq7mtfmu6xN0NoYC1nPGEcgHin7p8
vMWUwyKN4CrFIYVAhoxq1HHPIZ2+4fMp35BElGHs4L43ENVgTEVbolDvv+ur0TEvQhjNHT0k3YDm
mOhmy7m0i03gpjk/JxytQ/CIdgKDUPvUGoQc9BjHyDk5UjO6rp3w5W6YNhzO71xX6XeCpV5SQA2o
dRjzdMYVU0YFjlBa9xQQ1NJEodLKk7qeYl0gzfWtBqMVlD+ZjXOHgzizVCM7Hc+G6r+7JV+Imllz
46KOd9642NhCFyZzkAIsWQGapHjUwiCSPceDDX7TRycDtjz2L8w8gudpNR6RQRmNp6v6JUtAZUj9
IvDOxgv6cSwXGiptAXGMVQG7ZSnlyMH6C3N4f8mbstwIVnwdZ9L9At7ZHzGQl0dchwIHWcrq4j2Y
cxJXFLA/G940yTXXORactilJL5qmBO66IljxV9qQIFlvHn2dje/h9Tma7rWmGfVuU9HFMJn4c5zp
XpoK9tTdotTef+ixM1EP+HFAEIJAbYhuEBA/ASFkvUsB0wi1YJg+gSb+/q+t5QiR67ZzFYe+YJZp
tKKawdIVDv6cUvLrQbDGiRGcJzRqm5Lfs7QF931OeMeg5SSmDi77xCac+ljotowayZ170OLLqGj1
t+P98J8xpnJ1HoSM4lsl8W80jCOXbFMuzmvl5vlr67uHIUsNybwTQz/HQFxCKmr3bPCvjWRvLA4u
+kRkyX8i0LqmWPMuXwCxAadujXgEw0VMVW12+dx6xQYdz/fcxGX8+WlH8LCIY6XfkFivluUTfEb6
QlV3kqbtliz3ENT2bf/829bHGH3xcmLURNoh+VYErOszl8kj68nGdDZg8e5V6wlkmGCmTSnN9V5r
MYcJJnkQFO/kVkBMX/E58bv1FZrtlV2ZIVeugHIaCCWmKgRdLxVg+g8bsDHPDCQZFIaxdfK0CZWQ
4fxhKThgvsF0B88XxPWNgB3fIr4MgSiGBShGbWy3aZsHgg1RrLiCiJfTSXDTcCxYZ3asdzQpYnhK
127J3mMxxic+RvLIQHFk9M7s8E1lP8mU5WQPQbdOUhC5RiUANBoUNqkr9V8TPzK82V/7KxlW1OnB
TiQBsw9aIvUlpklGKEhQUPldh6eEUG6J3lEhy3iAXYXdIuyC4O1TOf5tLUaZucMDZ6JH4/RWOIt5
I51ikR7xsH3rkrEipPhDk5y/65DlBkDlm/rAj3nAe+4W7nOFcXI1de6s8tS5+F844qnCUNXvlKUf
0ElAy1qdQT01hSz6KvzltmzSU0ynlhmUzAoCR8RHZll6/ahsTQlksPE+fi0N/iBkelGyqNAGSFHN
uLRB9bc/RopSQ863eWMnxyLxMjOe6oZKEQDJsXgp7m5q9Ydp2DsOfjjY+WyP8eKl58U/Ul+W7ztC
AXI9lnUWX9QL7OO64b/cMSud54IpdcZSeCI6edhvh7tnz5nh7CUfdJnPwr87ybtzVUzE4oOVBQCS
qDcM9ywIqZR+CNJ+l05ieyPXO8I9O058/CVL0RylFHe1rNBfILoM6i8+SS6zD6Dknfh27qDv8/ry
o3Dl94GtApukbuT61HBMNHPJuBMfFDVZoWYptn8LwNbW6U3qA7T/TGwCG6OEtX1AZuHE7zOufPm/
pvncL2sdv9RALHojgFgjcspa6VJq1UPM75PGbMiFOgYN3BqihKL2uPb/R5eenmoT+7/8YeHRC6+I
KPCGNFO3Km6jh480MkEw3scymPoUWNtDuAtlIeE9HQ3zhnN/O7x59RUQPdVbHsjre05dS9xhUBAC
SY1DGWwICa974wFvaNiwsNEMTPCM4YT8n30pv1TGgEC/sKe+tp6CVcpaZzX69UqhaHZXOeM3Bq9d
rwiuQqaFg8boOAeuh7gSi/ojh6oXz+t6z8rEVoZhLT6U9Nlciti35JybXy75i4Q2aLON64qBDtta
OAw/rLjhPHjlbOI5YtM7cH4Zea4y7Pj1xKJ7XdDZGYudJUSsb5WsS+6UKO8enCDuaozK4Ap9JVye
UKIGwSNk7XGx2fuWIy2gn24Zkmd7A4JpSvzG79MIkNi/tfjJF/lBfeKuUJFUrHujHA7QOn2glmTa
h2+/XwGRW3nzfwyBztxqmW9IrYbsKWT8dXM65hy896HFr6jBLrqLN35Lkync69mRcil1hiUg7WnD
12puj4B4el5/nWIGJiyNEnT8kUdd2xxr8iCHcQSMoaG/XCiY31kCnMh6QHNZEctUo2ZzYRzjwHDC
Ktl+2vP7+RsNeVs4Ld/zVtpErwSGLWOmEnQ0Ute6GoCX/J4TifRzYsIf09EEIjz26y6xLKDYN8ul
0MZEdCxll9crkBaMED+54guAJnmrNukjQhQdoHPt/O8AiJjheQKUPWX7b1QFjw9appKDJFJAtHW8
NUSJOz7HpBoIbF3AioKs1G+zIUg1PzbhRdJlSLoPImXjvBCMtwLfF6JGGPr9BIxvwhWCgPJ7j7C7
4Ps0XZObVDES8b++sJzHa2UxiNoL4aln0J8A4qhtnjzK+9Zo045BfRcT1UzHnQ28yiUZuoRIs5Gn
DMhphIaxkFD7tEFmvTPbm4Qo1/4Ki0CLl2jzfSU0k5H7MGca1JILoLMVRRkFuSOtlFaPGROoMcUH
moCjxr++buAso0yXmJtom6m8EigGJKDe0h9s9iCW0fwwktiqWjgE2s/kiPlKRuzVIxtA/l5zT9oO
uaLmTt6IVUvXqvR9sSbdnMqCW9kB9/kforQuHjy/tHzHopkmRKGxJYvWP2zznd8n6a+WHhiNtDhF
hbShZPxzHwZbv0CN/cORwvk3jxXpdHx45kCHPz8mq0rTrzvZF12BlY7GkZBwSaFCaXYPZ5DtG9Qy
syR5ycbAzjZ679VmzOjuVg3RzmS/4Uo3FSRu+Kyy4ZeUT2ZZ0SkSmZAWv376YMJEZ+Jtk7jaPi24
bDP1bqc1k5+oWXpS+gURw0QOd3B59s4qufh2NyNZlImrUNc9B3pMSS2/StslfvNPZR5hSFOSBXvW
p03S2aoxHkmku7rvsYndu4Dh+1v48zvx6u3peenzs2/HTRnFc7cu1CtuVOS45ES0rYeByO2JLBsC
5H3U2SlvycKV3OjLBLt2xgt8vu1QKmMDi4K+wBKPnWgjZLSNpvUA1r1+WqwnGiXnq0JUDxcn0auG
wrsyJxLuo7G85mx88mmFy2s8Vnf/r+f3ICKmYgrfDL1jKN/PwT1n0kjzEFwNBlyBeNpjNc5SnPQa
D3MW32H3lgupyXyNeytkH1L0cP/BEzkRyxGx5JulXKW8FNxIw2pJ2sc7NCPHjCvXznSqYJETq+KM
pHSrWJr3pumfvztUIo+E4uOa9pabeAzYR8vmFKtiDEWDlxYY9bAw16ACnaMmu5VNrAtkzS+oDoP5
LQ7EYeNxNRxdNyTzJ489gR7CkhKCrSHK+X0VTKQoG/KozeIPmPTBhBfYSLEutndL1do1OdG6SrHU
syIZkAM0HzE/L4taf1nIyn83mPWlCEB+meGc5WtGuy9//9pohMsMtjuBOpcI8zDQ4IBnXxzchTHr
4kst/pCj7z172KyBzP7f6JCN/lo2qgNDlkiB1bFxVYWDVH+8rrnCTLvyS9srdObo5qcm1zku83dk
qUQ3VmEvwZuJZrEgow6yZwO4P6UhDQ/+wEgGIvqRSXd9VJ8qtV+vIjx4OamPqZblGol6Das5KTYD
gvHbAIBNpiuzafeqcNOOIlUgZkMgIs/FRiM0Nj+kNawXd2Cnu8YtgtHSdkSLdwuh2giiIjrPkRH7
Wr5yrTk+k73xRRmNyF2FYXRk5mHr4Xcbn8muoFdY414EAFKupGD9omgCeIC8wggUOtEJRUykmkdr
K4xBmm8rencixgJhZJt0s2vA9EVGg+ToWy2KSBje2YMAfEZk2IHIyphjf7Wcy5LSdkFk7M0Y1gxs
l0hCiiAVUIFv1tWHQH/1LsWvjojYWohmSC7dgtjnIXqu1RN8zooVp2MHdzjRFSjTh1yvQp4vAk3a
qzHlOI5TTINsCE53VOHiiOPctcL8R6R7HLeyzwnhuBqa722v5fYngMbiZ45dSaiqR+ylXkunz8xy
fYDyPEsE5nzE4Oyvh0U0zs9MA+jNPoV6HoRKs9jZrSNa2nTUKwGQ7abewQIyJx4lf+4gE9zfFqeX
4jE9A//77dr8dVzCbCchDVTWhZswPf3zS6F0rA1xZ/Sx9ohlMdQQAWuxO32u05BxnMnZiK7S7n5b
KwUnxn9X8ZsbfIyBSVVOMtnR0kwZIMRT+kec0IVJMWCMRbXOCL0rK1ynkLTWz6sR1CnRcX8PYlBK
CEfCQ/KpibEJtVQ5mXb9oxGmrJ3YjHjTsvhqMrOhHK89Zq2mxjUB9t0F54lQZv+kKx93SRbudfa5
ph1UbaZOfBMx2+GnHCdotanmp76FG6H3QiABImcnfXfk0SbkXIyZnO5fu5WxGDbSsxkWAYKBHISG
jQad0YWg1aqALyQXjmjvSEQAqv7+BMEeteN6YLMP2GNfge5DxBcgHtZBJ2IKbu4D/bHIcLaqHaD0
qNscn4VuG+ygkBYxpIHzGx6xnSBS1fYe9kkz0/y1/+Fp8vViOus5K53GUdWdE8MJ9xcNu7nzIoUx
dFXYMWFIg4HzNN0wCuUVlJN9N6AlM3yZGBsHcpgQL2P1BBV9jRuET0jQKwAey1h3U9iEgTdWQnRe
USP00TKmYaIgd/jWhvnyoyHvhrfzp6Lvq7RQqtrjfIiFvRK2xWy3JCmn6iF+Ih/cykpAyKQ6rs+E
Y5yWC/n8JBJ8yFPSki7uiEucUP+JWMmzpQ3SLoWaFNV6wZ9lPYoH5HvNSjrLwtap9KwQndM8/ZpC
/yc/r7KhvmSLQOca3kCwXrVQvBcugXcJuhzByEpgbLlC/nBu75k73PQBGCyMX/TY/DjsmZOv5m3q
CwxIlR+Fxa5H+gjFFYiVzCKHe9bu67VnSAsWJNqpu1hy1/Pajkab7MFizgKhk5rVaISvcJ3YeL18
vRhx0Ca6z0CfBea97dE0iD12HiRgoUUNdy8nJrImO/jZcIU0N0qvyVhuAGGLW2uly9qUKOxpKMk+
W5WmSp7WJWz2zu8T+dwPPD+cXG6I3f+WE3AoLzoSKGcBMOLj5yNfhcuXDgT3HYJMxZYsuFQbPdwV
b6dhRnQ181pBCkJazk18hBpHz0cexSM4K8of15npOftNtPfcus4SjU0mVvsGAkLa0oFMZ80D+n+v
AScWOQWS38Rv+cJRdlFrywt9dlg0Lq8AXlUnPQVutNEV5QgRzEVMKZ6QOzj34Ks24Ajfo00XewbT
sVM3fioiqHiyZSGw+U6Q2d1mivXkqRSQcrpVhMob7kd4H/3gVBUinpDzZo8lYSneI2CP6cFkb7pJ
rDS7Q32Jc6ia6rnIFA0q56Nem+gbmH6gh0C/5twlhmfqN/NtToBHozhKpjF8KhK4QsAHCOarYxH+
h4MRuaMKmDEbDv2T5jY9KPrDU4iAeShbDO5go2CZK+nX2C3Ybbi+37Z4n1yHnRB3Z+3RumDit30y
bg0Cs71jmnaUblvKB+b5O9XgjMzdQflCMbqda7qiHZhjuyvcpAHIjlOtt/pNekLb2gFYOjpZ2Ott
RdCjDey/HOV34LC+BgaYdBeArAvz359qJLyJfsaa0qnvdxad1P4zL92rMtYb3ni/z9QXo/l9KajQ
JlQtsStp+nJIRvv8X4C7ueOTKPfTEhpX1llOyUeOO3RGt3X0szmLOsdjAnBSSuqUFtr0vrTzzXme
gFGyG12aelVF6/ZNLok+lBWf3QB9nti5JCsJYbra5nJ4tnT8r9LdbEBkE1C31KvHj66UvmokvQ6+
jUaPdEj7nnGWP2EpyRwC5fB/saFMHo9slwd1SFnMHvMa5SEyFAETyfQroCjx4lIaKfYR5/vPuWvZ
WHoiaN4halr97kotm3AYoUJ2nW0D3WgdK/RtUh6/XHx0NFr5xoY36iEtvm0G0rFm1zwmvwN4DyJU
Sdij2FQBDVtKxhm1DEaG1voyoRgoGVAZIWH+GRuzHubfaK3/vZx4lncyLGYI/DVurVV29GAsg+4Q
57PvtAr9MsE+Atihhm7SfKJuDmszlBcd0OmzqnJKuPMt/rUzXI6nDG8ojGg5akCBxJ3qFrOwu5AG
Z8zFccV5tgLawx4TewgjDlTG/+9m/2DqtdcWNqFREl9ZhHt1JBEzXqLYOQLQC7EPrgn4wgwzS9yR
iTSWQTej4nBw6g317YmFUR6fvmNf/vRAs5OsVYMvUdb86sYkSWscOcC/ljELgBSkd5nyUY87uGWB
KAMCE2si1XrswygRUt/1xm++F6Vb5WSQ9btPOIswP4jn81cfzoZluZdEz8aQGwVdYpBhw+/GUlGZ
xHP/mxZWi3TKEbNvYI6VdUcAV/FIMd4yF3xs1L8Bk+nSoLCBmlY9uqxng7aTx69+ur9ccWAjuu0m
gQ1LGoomcjZllpbYoY7o34GHKCcG8NUp8i31y4Cw88khNsw6nGyy+Or6yZermYgz+uAMPXDdUll8
KvIEZ4yy66ZGOSbFPXJW0SWhLc0ABkvy0XB4KpMTFQX4mjpuJ/qnZkl1031fIGNs9q7tPIgWS48l
oDTeJRedri42+NW7/3EBBOVoG3TBx5VJFxS7+nUC87iYDtsA9rpRQMnpvvRM3oOF8/BqXCIreEs8
6jTZXE9jG9qg0kic3o/PHF/5qaiilumX5EjFfoBFz1ujjXK4MYkLUWX8oG4Ad0NImBcCPDpIBLis
ymZxI/OFvd/1sh7H7EHOOvXa4gMYd6dCtG4HRHpNfHg3pF9eUq3g1eF5Wmrlrnlm4BiQY4lDYSVw
w52lkEsQwaIqkd/SOmA2VSt6SOd8ptSoSv/Lv9QyqCp02B65H96aio8idaNskrOkorWZNZVBUp6U
bhvn05l1QRzNbuTZqZQ56hTmKEzX8fAIK27gtlOe73fvyAJ8X0YImgYEkbVyPtO/ZinVdf+Ol8pT
WOJ4fMKS/2cihlFh97v58ekF6lu3whncqyrERrA38eacrz34OjVkn2QwDWups5/PJnHqV2XaW7u6
GhMJQpABSitIOqWvhw4E49zDMeENntrGp6KgFb6owiFoSo8SN+aJObmYTtry3p33C07Ul7Dcy8zL
wHdWI7iL5oOi66cCn+5XHMGbOcpO210mG3as1tBFSKRz6HSgwg/7nborUuPAUFSBlY+XLVw///UD
mimlg9O7MPmgaVCgGhrwEUJUv8CIpTHpXh5vkdUkjgdPDNsMRuE6mbBFeRnypJRmqknVeHtnolnp
YzpiJHCa/Yr40F595PPj5vfl47AW+6JwIr4PTvAOkkB8U7dZN2LSDPGqZxm3W+GvBCPlJH/9ttOv
hFQ+6rHbBUrXdiMLXgugzFmCwEeogWedqZx+BuLqwZ+7IbNGIFoosDRK1y5N1l64YKanYFWTQPkq
dd2XgVrm9L365NeoiD1QvU2zYhrPzpL/Am3o6bhrFV01wm1TQhVnV+XOpiIvDb0um3A+oDFP4QWm
Vs18LD2XlYBJF7bNXY8TTsOhqx9DbCEIC7DT4nYZuYQ/V0TuSdcjQywlFOtIDxwX9cQLpCiSlg2f
GRy2rsg4P6F45sDqrbGVfBRLrChi54J0YDuY3/Cs1FchKYSLfaFdTWrBQOmJbYl1jN70M3He1CPD
SPqbK4tCtMN85e44MyqQ9VdL0+gd9z42X1Qki365YwpHHmOTnGl3kmfFd/AS7aIYoRs1fvs2+yKe
c01tn2N0CEqkgCkDEPdSLKvvjZ+GRt6IFEEmjo2MC88l/YXcsP870gG/bU3gmHHgX2MxVx8GRJLK
YbsXjCFhJCb+hd3rbe8KxdEXyTMYRqmvj7BsutVvT0NH0hbRU+QnJZrKGZe7gjfWgUnCc5FMtGFQ
rDc4nukkeRLz9Rzgfyt0PGUrJxttAh2dS5A3/pT7pHtEht0/9N9YEW2Qbkf7mLl6UsuiAHUTcWEU
qBSFqCNOWNgROoSaiJFbzdW21a7qjw5EYSKIbPBbMrOo7geZkk1Cvk+NF0fcstIUkc7ycLn8d53w
iKcrEJF8QYBra6pBlU5GE06KOSAOWOAW8VoN5ZfqS5HeHojwqXUltvebKGHeBKjPIkyxVScHwycE
hGbyTnUcM2d1EYx5D7v+7Nqc/Y1/cXVFVX2hdiVtZMsWWrymy3rMWDWFD+pAIS56C5smJywFDLUw
z5HQ0sUJLKIliA1vhkTmzZ9FJKeQeNCCRkjngVlVy39fdszor2Ef0OJAmzNWFxKcYG36nAR8F93c
dOqSDL3YsE9Ukavfzu1wYcqTuf3xn0/9VcVr1lWfW/oOxXRtY8aeHwMDVj/HI8hOgT/eZEWbs3Ee
eEAdrBlte9P6BkmSFBTR9ZYzYdvNi9Ux8sHpSPtq6jtYOyEc5UQIEIHcLb1GikiVnUIjpNCp2of0
vvQow4PHYR/iGADxFl03AsDxOGwtRJEPlw5LEu5wIWJlAIViDD+cleGoNkUE+939OoYB3J5XrkT0
zK4QiUMKN1D0cBKmBAs7OZAq4DnNiZH/K8yZJxILU/z31jukEK/CqK4/WyI0aTCylzI8THDJ8Vqc
QVhyv5m5xaj7J4DD822e1blEZnkDlP7YKTKigdVxzAc9QgiNiNmG+ChPJnDewGjxcGxPowETN26d
yE0jaDzcGnJ7plj1xWyjQEufSeWVHC6epeArBrFYJ7Pt74eeqvJphT633UW0Oz+D5XPp5PN8/1Hz
9W9FQtzujxmSrbXDgVVsloeJQcf0Cr2IBmUbQCrw4PScCoDbTUsULQ2kn3UCV25ii6QtVpAgGKze
hd1j6uLPKx6LWPXKVOt6oxMa0Db+Y6If0zdUVy3i/6AUFATGYg5lQlaCktHUremxjZob8hb/hZkx
yuQ3LIgVrgMXRu98w2kJqo7GDDtrpYc5tMr2Jv6S/trrxlAE8J+sVLaoL4vAj2OXIg1vYO30KAWp
6EHpcvxrGa0I6MzCs+64O5dlYW9v7IJAGldoA/ohMv2+nUaakd9fJdfZ0kVjAxkkHFNJwBPjNEAF
2rEnKFqxwzidUrXE/9EC6JHrhYmFYym0WxUvIQkb5uLTMCmrZOwZ2L6XRnrsFTTNYU03oHsIJ0MH
36KF+OT8qEaS1wqKWX2dFhh5Njap2tCLpKQ1rvIZoo4bw+UYtzfC071SebA8XkpWQ2j1jasNMug1
9fB+NOuyLVP7+ZL3q2EZ4r3FBJVPjdDiI1BMXEDJiqicoVzqU9eWBGuYCScua8OC+pL7y5t9p3Fu
9YjP/CO1qeEfUMlDqd3THY5nPwXtrvpj0Hk1imWG5lUi676Z26ptDF8hQIYwVQ8MTUPvcq9aJsVT
j58IVwYhnN4fCXdz2wFNJMBYHolgoyq7PVUlbb5aPgyDATzsTFCex0q5j8soAIWZbMlCp9GfrdDQ
X/jJ0UgobMoA0AYjV5eo8OnOHVSygs4Q2MK2Zrx+4ExRu+5rSWpWL1DOT69lZwL6JABgorl3yiYt
ORP4eBJfBR8HxHMS21aeFS9kRimM1ypOGlN/0yGuOu+mzsZEHf8hMYjau4uTXu9hleavBKXb1jVp
qmH0IKuw8RHpc2DkKh+UCG891en7oHbQVeFZKBVRHnz0xYbWiojmXCk7IHUCQmc0FJBOJxqDnpW6
LllasntcoPUM9ViMf96VNaHSmhktqkY5UON6yoQzeDM7520wZ4+ToWgpizDSzhZHaGxdnNcEVjVt
S/m7KD14YSuzLc7vk9pM8I1tmIgLQmzYTBK5lXelI0DgQ98WI/ONc/jnTlf1OWZtQJqYvDbp0be7
gnGxTN1vliCoHTdfq35afLYtXoerqljFFkSjmreGXKXzQxY3E1wAnOkIjnPmwnJ0A4Ie0zOjzKRc
oA3gYoEro98QaTjrFIGrVywgbfieIzB2KViEfcR7t6RMmcK/MQKG1o2vxuX7s5+7X3IPhu9z3tBy
lUAZvsrQTS4hUlsj4hYy/Nn/RQwvKvgyuEMFbOgZiVPU4WVLQmgUdTRoDgEkuGX2741N4cFCGf23
xHz0pBy1EF+WqTkcvl60rV9eQWjGv0PxJTtTATqnc5koADHziUVkrH0ea3z/SCHDVVll1Y7RpU9c
4P11xtRtWknqbwkhfglC7Ga6hv77DGxHOGU6Fy0WOHVj/hk5r+/khOKqqF0+fS+uYgBxtYq3cvo8
VA2zHmSiTCccWfrqnnYgBxMfL3jxq2UAciex90YgRVl+MqQRKQAphMHVrClQyvEQimqaQ+6AwpIF
MzsJKcHrMaSEXvmFmr2raPMqvEACeuDMiIwn9Grg8IrRsW/YMZHMnLmCFm2YlCbAoaMa8gF3R39n
Cf6vY8fNjesoAG0WSmoP4dPTxrR6bXGUGhW0MLGqYkrxEiLa/plrbSLUFDJwgiYeWUcefOdz5qVa
Du8prjuhUrPUAYkgLVFOnP/0YplBRQoJlgro2o5z0xMGVY97hNzJWgs/eIRFHPJgbWEKLGkSNHty
tNvXAx6ITOkXSSiFQGIAt4sS3oB0oYTmKtpYpPT5WEwfruknkUI0Ve4UwhlVubifN3HyggN19uxK
LEd4ZgFRkkSBNsqWnt1zahVb2FNIL4uPVEN8eyYcjb9WQcdsrCJtwZQwoTlqzLYL5FBvF6PlVHkl
WoIBylXZwbBstK/PzPoVN8Hh/tXuzuoGMTcnm7hMisERxoXbkEp5R0TIjpPfiTyEhwF/E3ro9au+
bCV0r+7C4moxoXFoMTm12o2R1sgjYSPioiN6lcuy342i8XvfvlgNQdvRTwMcs3fRDCmjh2LA8lAt
mJD5qB8oi/tw9fCzBLwDvrlbkCaQs9sMUhwVvjNRemoCz2EiRtHhNHy8z0I/XE9gOcqhsx7O1Bca
jxt4rNhnmngodQR2xzRkVa3wy7vq68P6zA4kD2ALxzl5zt1M+cTfr4WpvvR+Js/Pp8aJjzCfTWag
gilBHLrqc42PSlzCwFs1G/MC9BMMDH8k/kgM0MQ3dW/Ys+GIGXZeHD75Fwa2OxF8/lHbIjc66WZ6
BLuvCgQv6b1E2U2H0j/H5MNrKMrCDNTC6wwk9Zr3FWW+s1NhXaiWFX1TU3z/+bJzTeV4QFDz12Wy
157XJ04zYRYUMRxhxpNtjiHDON4xcDJo4GcB5ShRyHqkRbtJA1Zn9q1HzKW4GtpCRkKUoyiZJ7TD
XSU6ypXxR6wLCNO9TpGyBVcwTBPGZgWw5CEUISLnYLKLEsHhAqXe5ydDWvVybJpMXL1Gb6YUqWhw
mdYs75g00aiaLi58MsMhG0VVb7XrZk25cr0cvn81JZpb6pOuGI1UmJlcdOKyazH971Gp1ftLAT/L
BexkeKhUaRGRxz0GmvtF4MvRVKQh3CBAM4fdb/uEqdxXIbkTf1EfFYuZwVuLxdTeNiSof9/NvFa+
rHjxuIqY6T0I8ZIJ29jEw2VVQ7jWkbh3WNXvtRFOzZt/lUrDq7BgpfbQ6SN24kgzFDLXPJdd3qp3
bkqw5JCovlWHG/PnJprSTtzju75VtoHzGuuj2aJJ2A7Z3VunA1bnITEqLE+9pN0yQjOCbFp9uSEC
lMVfmenOHQ1fhDBwhxHE1Il0RJcGohXtUbrNIYsjNDrfHDsV87qFlPLpLuKM1U+gQxVSnWRFPIxb
Jb6xp6pR/fSqyjVigHfuzr+hCPq93AZLK92HuHhAO4aKsDA2QYhOycn1UPt8/evF95y1rClQU0c9
qZaYnzEnnU3JB1XyydBF5ORVQzc+djhnPlEPdoNErlIh6ROC7C6WTwYao/X3Ss1uoD2N0JlJ/CUl
nO/CYyV61HqI11SP1n1f0b2K6fv+qK3vIZ+Omqm/SvWqfZRQU/+GrSGXXyVSphzixjrScRiIMFHG
HzuDFVnYRqT6dBRsbMc5ZJUQA/XAtoaQeRLYcM4oSeWaHTpqIfzc7JObUJ3N5eSZJg0EPY6waK/9
m2et6ist2yl3lsNpSsyQqi9tofS0D/Us+x47tkXWNQFVPL+e+/9jQp3JeOJs4NYXgqKQYEvZ+jCf
UlEimW0phbCM/UYBCxCFFoBSniSTtMooof0VG8fVIckbTITr6JdiYgGNRNqNMq/QB9y0xD9mhldK
QyglVr8rHbkaMXsVjUdrJzwhhKl4vo0S5KRMVINx9B4iAqB/Bg+me67SfsK26D516PPQQU8g0UfX
DH8z23S6Yx1jV4JAVNGWOK4fNXYUIApFGK33PpCgZvXVe43CUix/00snwvuEJYOKF6vg88QkuYy6
TQpV11qTMHLqW6eBpUlIlNDKwnrA0IIn0xPlHZOmXLnkYD7l5y/PI+gQVOmb52rGiuqO7Totpmji
xjCqy0gLQ9W+/VWtPCxxaE7rjt7TCzhtPtO+8zG06y1/VtJcOL3PycZhdS7a+CYYV9t2KdqPoMDP
hB54dWIcmKVbk73yeodsIv9iNVoQ50z7fgZH5EOafg+EhTwr4MQAEojYLuxdQlAUtn2t4pKATw2D
fB2g44O2ps7zjecH0hnvQHEkxU2UPgytkgoXEwmmVEVBHGrFdeXMNHtJaNlWLHNzafHES1Cn0yyL
cE1JCI+2Eoh6Pt9s3CQN0t8VE62zBgIkjZ9JdJPGE3wsgf4E8hfOQKOFxXegFcOR0ojVj0w0MnIT
pOrzfQ9uEJTkQ0mAdLT3i9ucWca+VI7SyxbwEBJHaOQUEf2vUs+AUkEp3FKdcT1cSpzA3AUJsVFZ
eb9l9MWaSaIFQbbEDGStKISW3Sm5Kzg7CkAx2NVtYaBgzxB8Oe6exkytOxhXJsXZauvqJAKEYR/n
qW9nauGjIoQqqDuwTgyi1DZgY3wIXtpouAUqRjgJu243OcW0g4l7fkmMnZW9M/RrDVAh81poK/mJ
fhtTnkdnOKk8np7UQmaOA0RijKPyxs9WfLnhBzfTeD0qsuUvWd59GtnmrccdpdApupGjivm1+BOZ
VfXY2/9rjTg7oBWWzsMcbCapTHcGhG6P3Fd3K+MnTHMEittz5LBiUUchv/67gQx2oU0WfVv6NboL
uZ0FI/rDyZD6XxmI3BfA26a5z3SAq9LUC7mygUJ/vim/I6xtP/6VHTHDpWEQIMv0C4mdKlseBr6t
eC9csPeuJ33WaDSKcK5ZDqkCJJc+wtkiYuM6/h+N/qLl3luTlxxRcBC8xb9zOaD2UHDYuu0VHicd
G/GQcrfxd69VKjEQujoApWJpoTkqELyzxWtQuusB6ZQ+WsXE7+Qo5fx5DuZuz6eJraoUvxPJPSvf
lh1Zit966B5OAotwmlO19iBnHjWA1TwT/aoQvVEILnmDUpDFdXYIFRt81MWCgJEnj0UTS2zcLOsA
3J+dTIgaBfQ7xlERV5q5CdumZMlDef3jSmbuKQvE9j4Cpr9ZKb51vbPSbsfp7bM/sdVW6oORuQ9n
is1tQHExzH2u9K4nSSt4h6BnW2MqKBQpaifxpIsEG9VOFeuVruDBT6ND9YEKbcXPcX2VEiQABs8C
k7DIY1lLa9mqfeHCSoopvWWxXF2pOqQFG7h9kuNdS1WyN+LoId6ojyZnRwGQJGfCtPIoqUu6yo3Y
up+v02wqWZgMf8XjmB0mN0JpVet5l12JKbMqWAFXZnimmf4JmC9rXgPljYCLyjK0Jmb2bN8qAD6l
GOOjYnTAeyZhWvbiPEVGRRDBkGxOJZzOTywBTjLf8oNDrYdWYtQxc9bOKcnz1A7LnSk1R/vqUhYm
hbj4Ha7WW9gOORu4vMubho05gD63PSAVyIjrj/FqZGQWnCfNe1SpvEXDPLgDqchyU2N8KUGkPcMO
X4HHCauG0gH5u+6GiQcnZEMP6Bg/ktX+lQS+LsfPH77CCaFtCq86YzTQcZ/pH29i5mAuc+NysK/d
bo+shSowKFOL/RBz/hBmYhIu6CJQzP+fcF1BcrVuHVsF626X6bg0J0HRFkU01TBQ6hbB3o3U+pBi
NNK5sNU90y64l/0JKq5rr1J1Eo9ZFaEcicR37CSKGgbOvLux1ewFCY/AOqiHYW76HYKyGOR/NZ40
ssod+8TVEr/U6E8vk6XWT7Lh6zOREoxZxH0SmozaCmO4Lw15uBprj1rsB+5enOBnNWZka3bg998R
KuRDDHP+jfG/WR8oRFnCzxpqzsmCedQtD+FCqLYoOm0/9tROsKV0/75BeHVArQVGcBLQnZuRZdyR
JYlHGHmKnKrZ86W3+RLhiDFn+ChmM1yDMVVRs0kD0eboloadATt8myB7H+jkGdnjh12wPgY5T98n
BOQawjEjqwHsHSMlF/sheMMi8w0wK6uaq/yQ5sh6HCmCmJ1ljV1vnTK9fCpde+2n49BeldtyFrCa
IhRRYd6B8F2hXIcRy8EK3G0KOUO6wfqWr2gSY1RVDLevAGyHa10MojleaSUdPggD5BucR2lRsMHJ
raeJ73U6zz52GGHwM02zXNzUhn0Nzgzo1L2ZGaEWmiTVmUxNZ1lQt9ycUyp2tYb3f2h+hby+soBe
pskMoAqG/du5p/DwmW57YwxE5EdOwe0yzmVN/HHLc+MtNhuV/ZPZ1gZMRB5hwLrBEfvRc3eGWxPN
LmWjWjSPcynXSE8SwL+oYTTNrphMb5OIcwAl0/MKyEkHVAcEVw6C7PejDC5TaT1gYC3nwDTpM20O
py578nJaUuawNiud81YXXYG89Nd4LOpY1f9NiME7t1siv1tqX7Z7fYk42I1ZQ4XLpjIDE1+Mw7jo
TK8gm5fDLdxPqepfpUbhMiChuF2UiX9ZqHemWxCpAFL2VvW2+DDQ+B4EAb+G73heKamdQ2T0b4nn
vOAMuRz0S8p1qW2KLfaL8UA+NyB2hZkGgfmdJAoIFEq8gV71voavokD7Mou/KVlS/gzM5CcjIGE+
XU66fbLvhUFt2u/TNMM9kWgwLU3etYvWhriLDgJ6JeAVxGocz75IzSertUwdYaWB97P2u8gunu/+
p9DC1qgbmEPV6eTcZXAMtjaZJGzILUCvKTOknOiPeCeu2NIPCJIal5Ap2Z/seIIoUpw67vPWyjDR
GOY1z7Ym7gp359ENyd112Rm0uB0tD/4AKYqGAmDgsD69XXUxLCYnB1pwQm4EQh5S7cQWoEnLzcOz
yQjs2TRa5XmRZs+Hyarpv01+pP1T4VtZAa6pyKIEmZbNjDKHY4S1invL/azMLxoHzq/A31lhPcrh
T7k10AKhhdAfRWmS9m8CdZ5u6aQGWMEYVqQq+HlO07ZJjsUlXXHTs0xp4AnDYN9HA86bhhYAaUSJ
mI5SDNai24NyQPZlQDp2SVaYUYL6px+F5PeeGtANG72Zb8Nin3zth3SjI2lA/0AqYdUU9ofUAayb
WMSCkcahEzCyEbG9OVIXgXBMrh6PqzyUar7Vg64KKTSxE4jNvGt8E9i5KCJHQUmQhYtvcb7FrHph
PLsaqsbbPHvsYsyT50YpnHa9rQ==
`protect end_protected

