

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ccZ+VLNSpHtEulGuEKVDJLwcsmbh6zDXYYsSS4iGpirAhbXM3BP50jl4c3979n2YR8HDHLXE3QbX
SjQosk5Agw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b11dY0owYoWaWqrEwg1RlK8C89M14CAO8cS5xZSZiTQ60prhJpRDDBFmDC0asd3vpmdy6xip59nG
z+R5fGAzPFXPwL2mdZ9u5u2h5M7NuqWsd4/PSQwIb2Zc37lWRpOZZLKl9FzYzSgF2YNv5/jfYnLz
E/n1SJLECqBWTvKh2d4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NDjOIJz/ezAa2sanfwA4cBF4MUjfAWwRdI3fhKW6WomA0dTdlLUaUk3d7HHvjRwYAFZbgsshlvRP
BFUgnI13aIFlirt9v75NS6zbC9iHo4+u43o4DjI7erTR/V7n1KuL02bh7njjYqFW2TM9DCTV7yyk
HpE/bHTEqhTIUHhN3s21EIF7fvF256QO+AgjOS/tV7UeysPdiXp6gUoJ4fZfor+WTfQVkJeKE9LJ
0zpHP6pDYIRgknpLIxX5LP5O6x+a+epaip1DIHLGwD6CJeBzPxV1RVmuuHt0FXHAwR75O/YbsdQ3
OLvEz7nBONr7GpqlRI7TlZBuj6FdMW9zmU7ONA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
23D8eH9xZzeJ+Ojv/tdSxXVchNNJmk24MJAcRI99YbyO8+bv8JOBxvZhz4Qlt9qTY0ExdOGGGFmU
aQ35HO0+71woQEgUY5FOSxt7Z+X3DhAwHoCaoUzrhIzpo/Vibci8Aq5CktZeDbbFyKqw4AG3L+HI
gLdEde8Lyo1jpmEidTc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MgM0EI48WvFKRy0diETe4cjudrS6vIt7158toM9vdseTaMD0TZIog1UmAGNvdE72kJ9RDo475e8B
1F5FJia14jZNw9OSBZ6rrUB6Tjk4EmqoYQgrN7x0TfSl9ybfwnnJEUbiXZrL/obnsUVUxuBuPHw9
KwRIU7YdWp4ONQdRCD9vZVkexu3R144yonCk7ZQbQol5voGa98xXkFS5wJ9AioaVUGfDCcHlVgYv
dd/x2xkSx6aLm3qbkMFW3ZMl2N86VVdkP+mRZE7JGaPyJ93l/kjtm21dSkDxSaPAALmdawaPAmzL
9Uhkk9hs8yLNZbslAd/6iUfM8JK7nIIDO1E/WQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20464)
`protect data_block
MgkGPvqC16YDzQ4m7+IVxo0+R0Cec3k6Yc3ROrp4tbVpGOVZBHEaEjo97JiMh5s/HafQiBeQt1Ur
JFynQIRy9pxnRay8jzuaWpOr2KTIj8xcR0pvkvzcckK12bo7AjPaXf2S6fyFN/02wAA8f5KDQkHd
xLtkOCX5STy1nRvyGe8SHlTUr77w7AhHAncL4bQQygRDAbW0SMEUDjOvUaUE/UB3qIbwRmRiyRdN
/b/6R+hQS5Ine5lu82w9Z4YSDIHb5erOn+w5chJpfQ5k4nB448ySaW4/RF0Jds+W4fy80n+finNi
MHRjM2lwCZunRQGZayJL/Hvr8984Z4O51xv5jrH1pZOHpHV6s/jPHfhOSX9VxkxHFiRJiDrfdYqZ
pn3DexjkfLEdft5sfTlgJm1uHnJFIeSZ3fADNvXR02xNIGShr3TYXRxBJbAIElH+Tm052DpmXT+T
nT0OgzKKN+TabxoqJUb7/az+CoVyajeUbWfPmTGA//zvlEpxet9hSPMoueXigEP+f0KqQ6RD8gRG
p9cRpWeVShdmT9zxfH2drk+NtbyZ+x56+zcr8KNhUDItuAG3J1KVvDbJ285Qp/YrBSZ/W/4ta6vk
DbkJnRa/KoSLPFb1IvPQMmvUyNomhmHI2t04XmUlQSJjP/bh/lxc0xoVQ9FDv5Hkreg6iLcE27dJ
5k69WW9BgRcy5fbIyT3LxnN5CvvvH7y0LM67pj+wfJ4kIiUASbFiShn0VSUyuKroaJ/dafyIYRZA
NVcSvZ+hAn92xonru1JmQjTpZgUp0eYMDr9YRL5YcMJZzhJJUVRVvjn6APtvAIqoOWTEUGAqdROc
aOuU+Zq4+GcMgDSe1+P5Iw5i2rE8dcp6LM4mwyR/jfxR8IHZsANyJyB+F8dZ5C8DtpYTsG43ReLm
I6iqKpeKy2IaFL4acfcPkyR+WiEHAo2cKzB0VOaJI6kwpSllMT5VkBmzWBamtbDi+ryOV+qm3uXx
VI9pKYW6ZZ5rLUsEs9tQJ45tDMppQ/apCjKR20KlSI+PX+uvsEDe3vkcjRoqHGB2PU16OBR8dT9L
24p7ZdQQDAEzMhxUYt/uv2TXTeEqES8EsneOKsPzGIeizRLGWRJRSBUDnNUlPPf+BpWpWiU5AkOd
ijuX64qo4FJeyMczRNRAb4wfWnPjNO4p45PPDJoR3/HvWNv8QkH1ALPC5LRj+101NGV2koRCjPgy
+m0Nwic07PvBnlaGgdytcFmrd/jXm9fdUXuxZXmuYFozxRRdCYTPmZyODrM6zBQdsf/y4k+CNX+z
6Vi09DNOyRNzRV4UuFWMNQ0Lmsr1YjMMXkSZUF475uLghc4mQS+9zO/RYsQw4XAEgjSG84+5XKTK
eLAgUgZfbHcTP96t+UdKlLdZMrR4Gcne6wH7Fbrob0TNhwurK5bfGuHTKorhG66dEAz6LZEy8WVA
CCjJEnla55f1Chjzm6BWlAL30k2/LAK4R1tNxRdZ4Di450I2rMU5Rdyb0+SE9bvjXWETM3UPLUzR
LmkwxP9z9vSsQMGVy0K2SQKzuvsi6qI/SfLEKww34FDVoYq0E6MODn6ZNzLVb3thpdix8HKMC5y9
O+q5C7YPYOjxI2eutq4f/NTPghE16WvDj0RtqTCnMYn4kDFcLKlzMw1fqd1arXDInkginxl2HkK9
jN8dmwbctEWKz50QzYKHXpJppqalPh6eRIGucBKntG82rJvEb24l9tsOOGkqpf4XZpktfcXzmzbC
qZLiMIhvNJreIPCRqwVNvWfcm49XNK2WWWzd22rrjINALFMQZFQakDEwh9QYrv+a4vv2nGjlv+EW
Lc5W60fkk3UykEw9y8AB/jx+vZjPwIf1yghCd0A4KeOtlaiIOqbMGHOcLYagi3V1HD6ozrstANov
3jiWYyhEU3ACG8x3oEy56WOcVj+vqxuScNvhZUsWkTvVgXzzoo78iIk0t4zoS+O24O0mnQO2Vh/n
hp4HQapYBuGDrq0SQe1AuUVZPi9xXa67YWPyIQ8aFrqh2xzIOqBebfgPdZM5gKx/d5v22oRZnlCg
cwcuBDrxYnDF/gKchpTmbr8rFkEzas3/J8ZHHKXQNE/N5u2QTuji3mjjG0m/jTWVQ33SDM46lYbw
NfcF1XgBy0sbuv05shPo6+GBBamVbAqC2YdzSK6CBTe3r7I/D01U7JIu6tJWdaE0MQVZ9CS5V3U2
/JM5Fv4kZoghN5EU0LPH2MISUeS/DKF+e/sBVPVpgXd/EJDvXNay3hP0dXlKt0lPQkQCkUviIjM2
ZB6RC6ivQ0/lJrdlnOyFKK7s7sbhLHog/wM1bUBbeqYxCxbMaZuZBnSwgyWmvzcHyrgN4XMWCyQ0
SaB3PDNXxLSPyrnviw2R4TYXz2QcVs3sD9j0okV0wctFS+YJZ79zyM1imrbntnVLG8G6JGlbR39y
4mhSktGfel6VaC57xcmHyoIBKStXnPycBHo6KXeUmgM1egsYYMlWE9uILqzTfV7adKFEqKVti8D/
SUTIpXzQYi+NKzbpdNJ90f7dkNeud8pg1DRfHvj/vqHgOZGcmvHxLbIAw0TucYBiHzypguEj28nx
qsZcKTzwvKeKcD8j7HbLl75iabNYw2ynw8GVm7u5JaWmFX1IzBwqx9TdE+bVmt82bzrMxRIVORhp
cpxvP3IAJsQ5RquYuQ/fscL56ADGE5DQyvhcblL+64RfRGNzmKi67gucI24UFoRNcQ1FWqDQZqml
UCXiWi0p9mk4xgWhDkTFRT402qWJ7D1kB7/dVWT7B8UsZmaY1YfynDj/GzOaPFnMtGyrck0bqoT7
gIpmOOLrDZsUGzaenYf9WlUCKvm2Eu1sCmnydka1BEteJqWKtv0G0g+0pxa8PgQXHkTCq0A/O9y3
Dv904ONqSbiDTQ/sPojnJzPPRrIu3A5scMIts/efK6xRHFWIq1aNLabz3fKPicqCTvEMksV2mmwM
VpXUcESy/JV1NvUJyjfb1ORCRUcmQl/dORyEQnMCMg7E+4CHCAgBxc0kbiyhnpmZL5NzNnV9/QdP
NHw5ALW7dF9ocN95v9kRdhDl45SSJIHKbbr2Vz5CGR3Tf5Ld6F+vr2b5XjmbrWbKmnfUK2FswgtR
qPDVJLH4xDhaeCtPF6vTl0S5yG8AIJOecjazfEmrecqHjjUkA0Nbxf5yIyVcMD/w7SKKdwabVwYs
aEKrGXZCQarz223Z9nTH7sXiskOuWGlttDiGHa4K1fdQ0gJhGejZlOL/MRSzttdfR4xomIje1x7k
S8l+dMkE0Rc2+ZaRSDk+YwhN+s3MEu5a98FVNE0AQl3aWGMz19t6AbgUvGj88MkFgHi7ZVf7zcTO
8rIkliFm/5fxTKMhaS6JnqZ+WBWV5Ry2geO+rC23rRAyXHlp3cMRc5C57GWLpl8bduWGZ5G/SI2b
XXMGpuLB9zBkg/w4b+cqtvjapz645NEphmBDjgIJiMvpFd96dxiedxHuog0gFglevHMPz5jSi07Y
lgbVVuPuKAAO36u5YY63D3gJA0rPXhiDZMsIwn2gCLXB74wPYN1CPo64tZcEyAnfboQUQ+JFsuvO
uhOWZ8sXhW882Q0raBWEjgRASdBGq1fWhlh8bqL3wjPOk7cI8O4FfL/h8GdY+Yh8+M5rX96m2XfM
Nth9Lb3PSv1ob8spbXsXlYHNlATmCVUJEFV9r/7RpJYgRZMU9Gbjelc4g4oKrqTm9kfUXLQXCqZ8
98U8lVLRwmU0T1AIcO1bCBroqmNDtcoI1pS9NkKEvKmO+BGkSSRn1pLvZttfka0Wb0LrB41N5VWH
dLAughi/jGn87kMh3LGbHwQCxbuiokIddW2fAayzX//Kfe8SOh08Et/leZ42lGZq8hSZ40DhStNY
7NII+fuo86M1W2OSJo1pJSBBzQVLDeaMwUtv8hVtySWmysSL5QKrlgCPPOj2UeIM84t/vMtylThv
yiJHb/Pk62RgxdWKGhvEou2jA84/xGQNV9UqdbtXV3nnyW6m6cYai9NJ5NVuNKBvGZR71ApecpZz
NzAliT/CsOSCfPnXJgsIaem1mwT1PGJKrgvOy073bfAxZUW8G71LluNzu9Y1ICIWXnkLCAoUUdPh
CeIP86sQirWX1lZdQ6IhjWHBD/EwccNBdWUGDDlA2hnDJ/EpnPwg2cwqnbQMI/EHgkcpJEYNAxTg
ncb4Y6keKi7F2GOupFUfoJGCZj5xPvLcK/VJqp2gyKgdbWE0WmXwPXS/93eDH4tUtxKBX/t6s7Pb
O5BFJGXZbEzvLRccelnjZP+xWwrsxxNixk9apmZb1J5OJFrgxRaBemGJxBB+ok3ryTqMhjErZRSV
SqChbSvLQYkA6D5xRCSVjOWwcjCWdZDxOmei9BRo2Ew6EC3PhEbngR84FjxTgiCYROGqM1IepLen
9BwBGCSCgqf3JE7PHeiqiWQHwiCKQV+bv1iPC+lUyhaxuDoSl+DUqy1aAnHkUElwX3nH+vhruJQS
Eaw0Wcz6AgjPDeDzYhNkZdl8jCc9nz6AofWhlRCeyakiJykNqwgzb2YbEYd5dFVJDYygujuztlUQ
78jJhEuDcbOgq1Jabva0SduKy3XSzflkTAUmyHh9L4mJkFMIDfg3xqR2xey6WUXuIWnP9IG6ZZjR
s2MjjQguGpk39RExKEhuxudPC7ksQA+QcnX7LhINJq+B1E/1g4qVHENmEB/Vryq+39ALg41/HUEp
YUZjdZ3swRaNZIy9BJxwAPZG+HYFY4gSGMShcV2ujnQctOGU8cmmCvR2drwgSEwKJ/RB9CO+jNLS
OXgq1wq+3zIcqcEQx6fcldnqVDoQs47Ca64MlNagWWQnD5wr/gOyIcnqE52OK2YuoBtO61GXocxI
wHcUDve6R9vpGpnFkIsh3tUo1Bx+NVgBSGzb+Pjiov9GAkTFIfhHIR3SVq3xFmqa6sW0HiWTguL0
kFHr5cKV2chwHKyBNLCcNH45M1AJhhT40Iu6V7XWdvhEsP5f3XtYGPljY1KuuIwqJp3qqKh5XlP9
PNEL60Nr38fsDcCnR94u7eT5h5H9+MT7N8mpvNQWHVFHHebZohs+a6TFDvx5DfGEuzUtBfFUjVcF
2c6PHImRFdITX8Hu+XL+3IcAlsYrerbY7G+F5qN3dICrNhEXIePViiMEuKTAGyOUxwoxojVlujck
yEGdTOHA8km1GtKFZSU1EY/27E0Vl/2Z+sjLMOhhMMP2cQwr04GT7W4xF+YwpfuAdaOf2xh9pRsR
AiQzXKHSIhCofCPg6Ey3DCtQgA90s0pPSgbvZDwB01fkk1DaP5vw95ebIXlPd5UOQWyMPEplB81F
49kXNrjTxfemOHjZGOmlrRSosdmHBR4CTwHTCUlDiNMKbNJ0GMFo93xaYIGZykTYodTBnrGCpmgI
1iuJV3wtNsi1OO3M137Vo12C1V9FynVlrD5iWxlwRdgP6PYC1rAKCEMxxcJb8+z5CsIk/WNJ53uH
kIXBwuZC7V/FlNEMKY0gstPYG1UB5kpohzK81VaAfD3PUhlupc0EUzBuCWH/Llh+tphkQVb+UoMJ
sbOAg567+LyNJV7hUOJ2dRHZc7wUor1uvV/4jnrY3hkfIEx7/xe401v3gZAoyydfGvQOisbKu7Oz
FabWFVbl5i6qFzmABBP0DgXESLsvxy8ESiCw3WgMiHzZe8TBom7Ao1sh8eyKj4NBJysaqqLTDyoX
izwHuTV8b0lsFVvBXESc4+zF72XDYZPl/N6ObBHzTieucM/VZphdSOMvRONBEL6zLgaaNEXs4UuF
KMlvLV/KIunqBS3acBMUWcTg6v2XzBjHXR/paxo3ixrVkVeGli9xoO6fX3d9PnSXvkJGJJMYcCzw
ccpCnV8HHZy6zyibl8BnzYDPaC3/JejH6yo+mgPx2s+1cG6VUIAZXFGwfqRZImCumco2DFjT9t3O
MqC/CfyK3/vwkuYiPhz9dIB/JfV3nwDXSY8bcUIxQdHcbmKO3VrlLA8OnW31kVKf7elyNPZd6se5
ELW3wBg+0LtmClup2qNbxxDFqyMNsF49hmXHqH1gL4QUCGisbWaqDZbe8HtBoJACyukgjXE3s+DV
V+HrhqbU3Q6m9X4EKWso9rt/gbNuk+SuG/otuQNykWVUGmHURumXwobWIWv6fWaLgCjOVc5xcIFX
OmGTQfdEgajy6S91QB71oroa39MVF25s1CO5CsbBGWtFKB2ocMWV0z5iz+9qUJBStzrJ+mMpuJ17
0zz+NowSeBAPFLQ7fjysQd4iVVR2eyVleQs6btr1fbScd956NY47PX34Qc/yeCtF3aHJwHkPYQDn
srFtwlo3B8bM3F//ZR49S/v/YfdqUjS14TNGVFhfyR/RAkBmQMGFZwI9HnyXRuFQYZUxMFx5BT4X
TMgP3qxlWY16IeGFTszlO9AVJqYP102xe2StQ8ZyM1Ln/a9cUmfAuviEOcC/d/Bn1kIwJHz7CZSA
w50n6CH71STkZLcjuB2pj/slfWCnTR+INw2YP9ugMYAeRa+PGqpAu+opvvnQtgfknuuw0MS5Jnyz
mV/k3gb7aVCNwMZni8C/638R4O112B2Cs1AOHLHJ6poMr5wLNBK9xiFBuwQWoFOv6/HlIcpXb1yI
61XpocwmJGxQSYUGgg6NV4GpZ5gADfrC3SWKVsaGhR3KOoczPRZ9gTdVC3VEqQ1G8U2QUlLCDhS7
SOFb90PvrCXug55GyPPFikENPA98wO6IhfeeAPhsoVVlN65Nfn5sLvqU1CWhxaHyrqFOMk/ZBlm/
G5GW9TP7oO4opI1D8rHx2Upc1vyIWuEXAWbRmKGl63CG+1wubMAqq9z+Z006Pyn1kWlhny/LvtcS
Gv8AAajvp/V1SWD5Whm5g51saylPM7jlNpCqmdeberKUxX9scjQNNFtj0RN2lXdLOsZDcZLg8xG/
8UeW/7SDTiDf4UW4mEh4DID6zCowiANKtQ5bRFZgGAXlaUqln+uIThZXy/5DQ04FP2eadVbd8Ywf
HYcsCCtKt81TplCaLrOmpuo2A8JeWihbOkWt75kgSuqtZNlYcg+ktyb3FV/XB+3mU6xA9HkakyrV
tfxe2RZHo68CRhF1XhSVw0mj8H9xm758i246Tbk8cW8fUVhNm5dA6lnbswRub10pzSLqKKsCyblz
mOiDRHg2b99WsaH44xism/DSVPTRz2mYKJK+YgTeURa6h6MYiBdp7bzW+LKFzgMOSNdW/BroQZ3N
CrZJfFOSRsQs0fMQOqwHzhFkT0qQTna73IJv0QKdGmAwcUgZCGGXqhtcaRqmFHcO6T9iPTXb7nt/
DMcnElPht69gY/oq7IAPubhlnl4zgocvFlF+k3hy6eNwlwE/AUqopBfVcZTkIFtqWZyJRhJEVaw3
8WV+hVB01G2qj05QVeR1CY5el2GGj/LeG7AOxWw0BBcwmyyl/3CsuxHRNQtQ4Q0OOzXkbrBrRHnb
WLv6sYnNbuyGdveSEvxw9iT9wstQwRZA43TPMUw4l5Ph9r3/k/VSsRHgPF9HrNcnfxEinaCC9l2w
MOe0JFdKZucfTS9GjLW96NBG4trd74+uq0DIROe/P/kqAsne3BJ41XpYs67Yl0WuNAd2rcj+dsiF
hKcNpm8ItppnrQslA6DWMDhDVFkEqbYae8NOK/LXtsIBqzSZDhr+EadIcfc29Gurtwi20yqACwQ7
se+q5PDbLn8VdlZgRdF9gVHr0b9zazoSNfRbT29Xi2b7LMhOMX2GncW4aFJe3AHQ2Q6QBimgAKwA
HGoF6vgiGOtT0OltRIXDFmAa4dLfAuPKKgHYRlprf+jsxDT7vtf77cq4nlRDWSWO9mp4rGKk/ZZt
hKRklLPgBILz3Y8ngZr8vxeneXjxH1O+Tcrg8F05wVjpxBv4DT/ZpaunPDOXrQanVF/lcAB0kKpZ
iSKp5qk4sLNK2eFMTJ+fnstmMn0mYcvtEuIqnNJqxhGbbO9XuScGUfdMiYcvOe34Ra1mgGmxds1K
Tb1UrnNNSp1x4QJZRJqUYQ8tf2H9dHEwFurw6ixeVp+trAPhIMF6ruRo0eLdU3lTfPGdHpLGrECv
/ok9buF106n4plVN3uX18Tt4HLM5E3OKN+ybdSjlMcESxGFAkNLfX2ey6aa3D/bHgbiHz/5WCdEP
qoLAdR5uI4pxn4Fw20upCh5p5EaJnfXtcTFpS1FQWIdDImNRQYhUPsUxylCWtLSSWm7Qy3qKupb+
07GSFu84gGKJQTBUZDptLXElIfeeBOcrI0isgBb8/lrUau1/mm9RsUMKPpy8OJHlQt/a/TrnH4q+
HY0Vp8QedCB/RT9gbquOha1sG8Xs6iYL479N05EzwPI0+I8lW30OeAF9eSdQQum7cWLqQpyAtUys
yp9giaZyw+mMtoc6GAFxDr0Zis3KpTu8qdGD978e4xI9KFRxklbdCu3197MwVGjWwuvrdD+RTNXE
qW7lPcRIldKrL3539Ej1EyQbz0OIGATpdmUXbVDQhjqBt7iuX5aXh/5MN1b0bNGyvIaPsF5IKCcL
X9Tk8J5BUN/igCNu6GTkJmajlkz9KxKnIm2rjAvsdPf43e8dLOJOD4k35LurFOG/C2X9oJUhiUVu
yL2+MorArrDIrb1hShXdP+DNavhTCZj9tShfqngm9GdP40wckz/MEOkpsDRL5XwsU8PqPR60a9NL
ODoDy18bBByuvCWttK9AE/3O/ytOWBF7paZeOXeA9m7Ubzb7ZG1X+p/3NikGc58eJZ6lkty2VQk+
zTTBepQQz30nV19cKRwBYQZsJi1cYC+zGWRRuGApjv2ihFbqw7KiAJKVr9rciGTRZSubMqk5nms6
R7IalGE2O7yy4eJJXTw/oTJk6ytrTXeKL1Rh1WizCwDHavGRniVq5VDx89XdUwafNlRuH0pIHV37
1ynxh80j1CIF6Q2T0zm1YjsTmBHdVDnPi2TCqR7YdB0W4KIOtz4Q6JT6lZiBMy03JQ99SUCxxrH5
E6yQKCqWny7QmKuC89UHO3eerlgeiMRgklrMvq1LeJA4C/Gi/YhHBgoFl3GlbTIq3td3pWQ9VmD8
oKvXr66uO0PBn5Kkv936VPT2yxv4P1MBn/8U/ZhUjrMKgTh++jRZEgUi92FckJ6xGG1D6eWs2kQ9
KoFKfm2a1TFhtubTZDpGR8LRem29ViMtHd/WiYHd86TcjUctAw8AYeMhSFyt81FvFrADrnwvI0mp
mlG9AILkjyj8Muv5IKoEMd2+B99ycOCRRmCLU9kH2qO5/d732IMZJCIhM+IJs7iYWeE7df/BQgkX
KXxDyyvxm5VedIx/cf4jiDAtbeVjsCkWcsThKFnkNMICT+IRqOsqV3osEO5EAVDl+eTIsjZBUUdt
gHeyOTNWM6Ju7LztCGCHBqJQaiC499OAhCmR3TlvVpXsAPiOyft5CF0T4UYyLfwbmulXLuwjTWTQ
kDvVm8HYutlnM0LuQMmge0RGQzENtTivii5pGp4kMLk8aNzw8a2SdgjbIVAPOBd9e9VxV+IlHVpT
EyLQ0O95lT6Ae9aUmNKVfuTdf6MjJ8zG+lRyBS+lrYZHGZgczuVI+l0Udvch3OWWAY/kUtaELA4G
PYzJ2jRWPLrjEUsBnZ3U1JHLyqBY4Yy957XEdcF6xn9m1HOG6Dpe2cdUG570QvW2hWhBs9fNBQ8N
DxPpy0hoC6Y7f34dIhwaso9PITlKXnvF+eitz5KprCTie/hxk0oBQYUWXZR2zgsvjVhlSalwiRkI
FNU5EjR3cEWwT/0vcnONqFz3HTRLww5UCZK+NmNxaLL+tfhu+KsXlMUqBFyHx8m2ijwh9ri4eRQu
VGCyqQk2crNDO0kJR7BrNOmsQrWgAGCn9EWByy30a0AOOc+aDZGrMLUH5eG0yPnp8MzZXYDuT0Eq
/MUH6jxommvCqRBtl6DtcN6CJAJXSlmF+jw2tHWoiqO7KRrk92CrAzi5gt5oNeAfpEasCu4YMHzx
R80JJN8CAjH9ZDBfHsaKPrZdn+gPBKOSFR078v1G3/5CvFEZAv/GYqrNFy487oeMnH9Rcf0rSqvH
pFYxFertlhnCD8EcFZdRx06LQEFtDVhh6JU4lBPpizgCHktbtiY4EdfGJnudBebaPleH0hIfaPIO
/MazzkUHne9MIa208aedhiRn2V+6q6aIuXfBAhAHJEmKL7mKvxphkgudlHCSrhPcn8xMfWfq35bV
kT7M7aWFZgamEf7QhDl0NAncLjzxNyGMGw/bQIzYgBOP3BE1Cn4EyaiMbbH/3o3dEArGUk12JwW3
qvaGrZaOItjwY73D7C6VHBbT7D6SjAOW2ByPJ4rspShySkQ0wRy8RWx4opyqBYZONahttEV3LflY
UOWflfCNTz1oS2ZLTCUR+JnJZG1mfP29Q31xOgaSAYJC6hyU+ehLp4yPlJXycOyzxM9vfS+g/teR
HNScJiOk3E6cW5ChC7y0Jg9qJC09x8Tggq1lEw7GQ24OpA+r75k27TyQ1IHHAZb0l7T23fEA3G6o
bTcRMhkNcSUz9hY12lh5xbF9n3kmT4E8nhML0m3Pd3iJsvRt7DkC6elhPTIIBabCXRKT4U1hDeLR
T9aN04w1QqdbcqsC+D7deJ10JD32kM9e3SSMrhuhangvNLn/NbbGM6jPPF9qb/RTMOZstGKUsP6/
6/pgmnKs6lh9UpB4EM1E7NNKHouGeVwRECU828tXaZCgcK7myoYWf214KTnGw+5Pc/UE/Z3j1yDM
xOaYcnZ6WCBtkLMfzgQAfCbRk4b0qINcnWyngDwIDuGwlLu9dquVu3ISecIl7+d62F/r+FykSz5p
jpPWGk+GvGBCI0GNFlyaNWteAnfbDl0CtblqwVklpnWQLk9YdQIgQHWU7U97e7hsG8TlxjDPP2p4
6W84Ti/9DxOEmtu+gDH4HOw0gxpdH6zIx5LEQZTniJANBTJPkR2sOuyeEt6jqvAUjmn/jooePI1F
v1SaT9yvdYMuyZs/zT/652HkluPnNuupOShb9CTQdJVIDAEDG0+BRH7XfF7HYwH+f4Y5ykK61DxI
eOBtvzHRMEv8JX20IOG/4KfF2vOwXB1HwgxbCxiGaCwxzzxWiknFfjw9LNMcRNI1BDWyOrABLRhv
3OUGbSGfpg3u0hzsj9bJb3Xt4LI8S0CDjrshljB9wOOVaIJh6tJ3589Ozx8MCW4BySmiInGVkR7/
82h/Ax7Rtc8QKh9pCb3Sh5NuxSQYpzDyBQnUIYZT35dPPGW+LjdYiDbdrYmDAUd0eV2ILjCszccX
b0LcHG6LsBa1+DLhlC84gi5krtDsxDAUEpH14XssjVNTgOEvL6O5StpC54qE/hcrVhrdWzGkgEzb
NXMdt1qQ3npaN+gYIMfukfcmZ5eLq2X3T60y+Cj5C7QSPb3xk7T3BM9Ba5wA0AC3ZvbQWOgX2Dqz
zJpLKxcmiqYOdMW8se7nuA83XQuQEneK8hzKJvOQxMXhPj0ggv+2uJ1SKAbJi8kXFhlwhkwd8kWG
K91rF2ssaxzWKzaYsejHNtXRBBg8NhexQhxTRMyKIN9V7TN1icraZeVpG5LIAO5uKznwii2CcYt2
Nk1i3OdUlw0D+P3IbSgQMkaKewV1xKwORb2tWvKIByD5FCU3+E4tEuV9Slqu+SXUKFRYMMP+fc2l
p/S4UV/++fd/yxczQECdd/3/GlnQNCT7s/+1Uggr23DEcapTvl6qYhgQEnGcsIBDhQx1sCmbfuKd
aLTr9ZPKf8ZP/N7YMAFRssFjJ9bSNSEjk1aXmmp/YC0l1mV1r7uk6y8gwVEtV2OOWoQ/NUOqhHYW
BWBVJ9k5cfnSpyI6rXVlUQdYwlAcQo3da/bt1/qJ3wVXBF9PMZlnBAcYiTAboKKv1DBIgO7l7d+a
o7rz49Yp+Mzw+eL3Jq0P4cGqY2YHl58c5qIrt5KPNnK2T3tAq9Hw+1OGLrfAhm11bZFtqVwfVBdv
dXh7YNETN2v3UaA+BFW+Y/JZ2GYE27V2WuLJvYauc79oFQg6LD4Ub7FRR8vhwCwWyXbvyioALNvz
liTww6ecQF6rLCAK7XuPS/D4tF2KOeDdxEom2CQnCML7MXuFsj+knoeqIl4UNgeHZf54T8Jcg9lV
uR1P4kOL/++UHJsHBXVy39rSdsj+cHPrwA24Rq8SxUTy5kNQPp7xLXLgkcYodFdBj2YvNRsOUzCU
28SpHYa8EF8M2Ux+DOjJPs5H6M9Vj/IDejk8n0PiD7qE1BQ+4qZgXL/55lLcKHWTOqG3+FMiJau7
syYOXB8LWRVrbi/KCX0F2LaxifvHYfc2oalaNt2uc5iseF+AH3A+eSkAr9R2DbvCAmaIPL/LBC4B
ClcuO0CZMZNbRx9EfKtNXxTaojsEV4gszJqfKjCzhMaJjPwlPY8Zmm5O8FLX7292+tInLt/zdpdz
8Q+/8A2M/xB66iHFiLsFSBNDDgNkfgr407nOyqVl8X8OpO6+f1sYiTvAfXejYdhizT75R5UQv7xZ
QEbFZnO2b8Spsez0vKt6SBPGG73AQGP5fqHwmW9zY8rXXt57HX+MKO0jHRA+2e8zLmPMLCBB06mU
5OqwQt06Ie4UOW3ee8bD+jhxTytVgoHNP43/RSYzlHCZ33X/ADlrcUHxPnBbkwXE6m+5X9wlRS6i
b9ssYETdNGaZrl6E60fFr1hPtoOwv1hckjDlWajU3yTwvH4RknUwCr8Dmxjkq8st7SWOYOzG7HeC
nuIfZD44eLO6MDdkgiekYnwXFNwXz7ZTge9WkjHC7vEOhPv6iHcUeSoF6VZG8r2eluyB1yzSOUEi
2XNF9iNhKpnTNuMOWhJ9B5RR2hwidR/O+xAzlq+NiEFc5wi5EcpvIy7qWSfslKCvGz91Hr6KvYNW
KxB8T5UO3bT8+0h9Mg1dO0Tuk0AxGSeE3zZkKQE4azwOlp82IoW6EuKc+wfXHvfgyBfs8BZkAgdX
4F28IbDNwflATze/UYLdS44QDWxkqWpLVS6g/YmV62MLn6FoBLKy5hhtTnp62i37xQUcipIQHFZy
8wLAv9i9Eb9VwRtmZHR1dhfauwkvC/HJIVZxZftYLqrsFsieUPxFoRmW0QULiyTBl3l+dfc9buO+
WNxUF1S0GH3Q9XpEfv3ntH7pbnVE67092SNFKx/Z0vqg/LV/sEqL+6Vui3heeo+c+RuR27FvNCzp
l5eTNolC12DvGjDmSV4BWt3HKiquURosXMofTrZYy8jQA6+8Pu74JvdpuI9pQyRgsuyWNMsxpr3z
i1WMZ0qcOUIu/Ag+G/+8l1fBeqfcQdOOrZAzFEUgo3fzpnBGhLEu6RbKGqU7xKNk/cmz49czGJUF
k+RX0pVgybhH2fDmuH2AEzsrCcj2APnDiQCZAkL3SMpm4YiEoWlaUD/uE4wNnHXk9DOaxkoMWsc+
cPRrka0K40TYR3r57Pm2pQr/+5WSCoJyHj1cIJraAD5EYurVKq0yIEl2Wd5NRjT675G6Hg+hD+Ms
V1vr/gk8/bVm8CMwVpVgGBld5r2jtzwJzFBD10UP0qdZXLXxOcptBlng1Z0V/WCpx49kwGWWVP3E
esEUcK1eKddfLTgNkK6HX6KIt+Ukwxt++sQ4f0CkYO92Y+VGWnKddRikkFd5rqPVAx8EqkM55kEM
RJ/FXrdtACQh/HqVMIUwMuonFoGekxQ/ej2BstDzhN9x3/aKUyqJyyjKjs75SY4bNgtY8dGauzVS
CUNwEM6vRbi/5ULeZ0CCqLqJ5MU2B/3uEUx2iiIzfnbvEVrtIaQsPbxVmr0i7RuF5kpQkFNmmX6D
A0ezSHubWzdayxFDh7HwxWik6Ewh7xo+rjDDSHMl2MyC3oZPMoM7ud/+9YMklxf7zCR8CMk2ni9x
BIDl3FDWkKVdSAi3lbMNAUzk9YEfijDB+W8T1tXPiZIoJi5563a1wYMVbthvg8nMiuHa07R4SLqu
aBDju650gDqk2iM9OlRYyGKP5tHz1fCcJWIt7jlti871l4OT8ma8Em/gIHIvPkI3ZRvVN6nnLpri
FRS5OzbAfgWfQIyH27NbYPJ7utTGJwn1PrECXilOCQ/yZftK8SWw8YuPtKP7TlTj83puhMMh81op
W1DcAH/RP2nth+LT87HQRI8h5KOh9CSdJUrBeaI5Ikna7P6jYIWvZttr645tMvWEJMzSueI8HlOu
Ghg/AaIMgdC51IAVAFl9+u7OmlhiyOCLD0+WzMN7aeH7v7KR67+nivS40zAonn7QdWRpWUsDonAt
v40j93F2YpCbyACpzTeWZge+0p6mbqSivviJYaPdG1elxfywG4jgJzc7/k5cot4XbeyzCLShPxB4
UWsCKxuj8xVatsjqss8HxcDoG7K4LUe8t5as2nXbTa8DOKceSAQ8AUjNf657zfiSTf8Hr+ETCmnt
LBtrF3RB6/HR8L0E1ibbta4ak9Fw12zdTB2sU2FoWKe/qR994q9x6PmXYiijQqTBA+aM4b53iM3l
5TeElzU/djHTUX8nttwzT26DQL99GmEm96Fy+BE3dYb5f2APeLiSSS1MYzsTm5CY2XYLRzU1t5Op
tft1RrgBCdukPmmnMGvgGvupYuDOxZtxb9OVB5n8nHK9qz3NThaJfcbmKYzGmeeRtwnFTNnYnzhZ
RdekD0Ig6lH7fOCAFrCdgTXmnkC8jG12MbiXYRG1CAVh/skZnPQojW6ExMXiRkiuHbcx/SoPDmN6
5uAdOCVR0rc9BtaLcMrwELvhhJqopohUgIn8ghTJ9bYv0U4re9Kc0Wwa/J6KOJCz6GDQLs93Tb3J
/Cc4pFUenwtp6P/Kly97rdx0xpp7+AZop+ZbM0tl1pTkqWXksRE102CcL1XzWe71sijU/rBASjIK
14OjqMycjw0NtAm1WSa0meuXqEOQv4zssiSLtvCVQdLtMdqlAvSnTES0mbvSq2Ueq/EUansCdWkv
yAT7PWpOoPSYRrzqCzSCGyPlE3tWxpQAA3nFH7qu/c4D5nsaFxk1sKJ+iHc0LraGYssSG5ifuxZn
c2mEl+hlNRqdyYlPyuZi7CGYEtX1xk2A2TVe4DYZIoHnYF9E6QBSTGvAFrQiZiDYkvkZvcmrLrvx
PlCE1FQ653Mj0kKp+FLYWMf4JB29a/ncH2c0PJUO98bjx1qFa5qiUev25tPUYUclgElXNqvWyy/m
VjWcjPix/ZatqSJigp3Ms1bw9+1K/1ZCSI/tPshBspr+Bxc0wqayahUxE5j67X5K+Lf9LDX/GaXM
oP7JQWUmJgPGKLhNC1aJw9ctzdFQ6bR3GITXYP8Ujz7+6uUVvO08XbGxg6jVv89/Qf9GveMlpc7i
3a6PYSP1QkwnjDtcjZ3THxeoLdX2HaZ0rdgMh9ZJj+XnaKhJshUHLo8CuTHRkXtWTFkexfMTgYBd
Eut0ogu8w9gyiKR36BWpmKInHOMbuGhOROj8pqsPq0OdAsP7yHmGyd70Dexy3PSliBEqNJqonKcw
w7DAtXCV/q4KdBIqz3pV4zWwW3Y+VJe1YKUnSQdlyijlY4+dxaIRlJSVjBGYKt+XiDgnWv0hLGNx
JcIkY3Ce3hwSccUGElXf7Ki4RfYzBGOzDTsElx7XQkyZMnb+y1ZZkOyG3xMZeHmQvCfZ9WkvvL4H
jDog82OvxTpHhVOgCOXDlZMW/fv7BBqYLTt2AGAbocRLz74VDBkzKDPfB1WFAP+M2cg/kZt1CCGX
vbn9edXy3N/8Nbj/MapWy8zUGgSvZoi1nj9FlNKm3QrENrN5eV7M9Lk+zHYrVvboHxDEHzXnSYzv
TACkh0isUP9YnKVvnuiUCvE1Wp7axskkWJdWd34LgtzXECuGLfb9HZoUeWy99W/+O4dVTeJ66xZU
du6yItltezxYkIrbmxwxSsUvTXXsQB5Z6k+rHCuRG+pF58stuXE9aJJ+Zwn357Tz7GJaF1G4Eij3
Okw0sIPMwGpUtJn+02q8GrfRc+pKx6V0m1RkAoGlSyB3K3yqWYNXnwwRPIAKnj5j+daF+StyFlCa
0H2RPaKHjmoM6zAuhIPKhvwTZi5lvP3W+IXe+8Blgu3FGNQcPNXnUCj/imfT+wZ3G2tEQklwUghU
rkM3TVmpbWs99GXpSdFpN6uX/8HFrSjsqYV+W3OYiW4xNOgojp8pAa14YKkWanUKsz96Cs6GcZqW
U5Vk6VfbtfymnHRus8eREHUZzjVNYAGEBpxB3xRuw7KZJ6Q0QyhHb+r47ptBEJkLHtzik20InYGg
2YWWeIUJP8PFGTj/tsueXE8JQVAW/Sn0R0s2+g4hhLpNKOq5qdK2REUbu8XY4EjxZg4CsdqlML5T
TxsnWjvVLmks3IxucOScg+WVXos9PahJSU6UMyztudIYlvQYidwIwqlQJa70V0wwNtYgfPQ85Y2z
ObrXB2jXf15CilNLkuk7tvKgcNPdKNk74a2K89T9cGl4z6EoAUd5UtNbIuAdsS7T0mJ0CSWe0oef
6npuRf0FlwIlSDabZnsb7fByqQhBaqs9VOGeVCFOnniESUzVfQ7mqJ9RgOZP21L83tqyqojJkN0g
KyPqhZOGW7yaFvTinwfsMvnIwu/g57kAagu5RsgalAUOcoTrJtgNEwZZuByQE/J5Q+M7ULrPv8lD
7/gMQG6fTCSpScfdT70jizc2E9n8kDqPKFnAD5NecfJUQftTryf0n13IqAwRK53745U2Z4ZloRpV
WyCazzeD0VHBm7HpNw9N2uy7kKLx0ZBNarT6lik40mlIZsPAbAwyo1RtMaLOsvA+fWAjxEULibPB
BECqRW2vokNOSnlRfRAOOs2nCDvo4ext0KFfTlO8gWaE/Qiub1NyYQhLwoK8blg677Sus2lMyXAR
4ZaqJAZugMQBez8BRAKfawNF8ae49beXmNM7qxLKvck2g5lox40nl8VecoJVS6gC6IjjY9qSl2lm
hlRUbYGCt5NCYDeSFT1/xCsheBOAaeT7eqjSu/2LS2Fc1LJUzP2VlusH0A+YNgzVlRAn+iRuKpE0
VkK7jRN3+/nWiDt3AhCyBzSBm9uf880SDeVLl7lqXoH8r9Q5xm7ivJflTa4Wp7GcEr00Br5Fjylu
7rSXicqV61408cN/eydYDrJvRbouZJjiFVfO8YSkhfojbFx0U91W5ttDZ76FcH0wD53TQ75S3xTN
7ow3MDnHH98UeOJwfNoHwqkwYMK2qjPSnMY+QFfwp4+351Ej1fhOQK5i6qPxDVA+tgedzeVBq2Jn
NnSFDxCfkTJZ2gVmLN2YBJ5Jjfowcm6Lh4nSbxbW9Wf7IzjrNJ78GkTHN/Nt+ddHp3aQyH+CpCR2
VlUofy2BvBizsmJMsPq9KJMRcv4HbK+u3MpOQs98vXpvGqMRC0K4N2mjUZTuFkUddgOoGYe1YCWw
4gd1trSrWP2Gljf5GJmP94ArUTHT8LcX1Qabx9sZGgfys3xYmrSKaALKzTX8gu5YVnegbFwfn2X4
GPf4BM4Y7qwhUEVlcZNG9e+lYn+2ES+s7/oKCrCbBGc7SSrXm/17ox9hAl7/2o9bA5WJHNg6igaW
FlWc4Zrj3zfTJFPBAP8rPBFXCcOebV0Z4WPJz3a84Mx2NaMSyAyzgC/nDc0pS0gLTEUYn4f0nTde
u3knqkKj9zfYM85schUX+85O9MhsCgVzvFH9S+j2W/NlEV0Qqn0XOuvvsohPNkhdgJ82Sf3mh/lg
Ci2SQSbB5nRiecFtIBHhZsen/uXzmMjZvYUpUC47wtuxCIby+JD8KIAWunGYyfmFOesE6lc6Ziy5
cbF+HSLb1YBbERazSBhSPVrD+lc6dLVK75bGXX+JqyCY/SQJraY3uKcFwOgM8hrbLrxMnrzdsgbk
WbAOVQaGGfqRJxOxASXbd8GiskLOxPoXF/TIhJM6pmNWwUjdf4TuCw37UWYHK7t7O7QP0/bSDdoO
OfF6wO7O4PWGEyaLNO54fZHiO4JkDbige4LzoOGRC9rG2cELUTK3hv4mhl5Hvg0d4Gb+1+Q5Xffd
Bi2v2ZDpfexxbtieYxVn2Eq/9ue4Kls8iXib9QHV0/dwiJonc8zJdePBD1rNvDDI0AWCOMTOXfDV
u0CmxVweJ0SHTOrAifJdTHfEwALO5Q1LPtp5j6mPym85wQ/fJpmgrGccPA74n+syGKZXad+wTdU4
GM8F1PbsWj4LfZ/EIfnJzm33FPK9FPFkx7tnmeHwlo05jh1z6UA2sSpei86jWLA7+ZTVHNVOO08c
xI2Of/A7hqLg9Wb6d1Vrf/vwYfhncgxghSg6C5VLjEoZPI65z2EuVS8sWttUam184tRmcp8O8BRY
VDXcJ2SfRQGOtaL/Y6BZFs2l520d8mB824BlqxNXH2NK9p/HbaeFSBZp/3F6oZghFic0J10nLpA5
MP9ho8RBMwCCSOdNTpZyg+FIamR162Qy7ZkD+qemNx2YreWeyQC+4zx8X3yGGsEq9yl3aa/Jv/7J
aflbQFElYRS7080+d6GtTatHrEL7U/46dB4HuKf+g7SkRDXoaqHoDq5c8kYaik78fN0Sq5N18pX/
segmslVNTYIsGIEIncs/zxOL6jAWZUjpGOJ3jdyIGSfTvxkIpJFPbYOvwrceZEY0c8HURmxELwND
0f+McTK5XVej6ncskuceURm++QhstxfHTV8Gum89DJlulTk2OGU5xp2CKHW4bsHA8cQVgyF5WZ26
BkFOy2ITrl1yzwGo50fm2wTHNsWYXlo6H99Jd9nzDCd1zkpKEGjWJCPVatKRXdSHNog3Gd/qzsm2
LKcNY2D8NrCsGcPKUWNG4uTApExIdiL3YbzS7JuEpA8bK+ziIyISt7gn+RR2ZBfp7XRWNjBUpGWG
vP4c77LVpHMtYBiefLyIACxbxBpK1NwE2fbcX+ZiOoIaDscyFeJ2iTye0Nq+2TwtAsoKtVCWOctm
Jors2mYdYDjIGCxr+xGIh103FjbT40BjnM765hsHO70S4KWLI9ErFFPk7jszPIHuIofZRueLEdcM
ir7cdln91htVpSuip2hDiC+rQKPO947gzC+IoH11jc9VwsiDc1oXT1KnbiVDhIW0to5vgseS/5tE
XRC8HGY0n4JYMmE3cfPPGHVpfjBe2PrA/VJzQ/4KFpfAQbPVcXT3SIEeiQtDcysbXousAdR9RIby
G4QeF6Ykh31JLoTaBO2SbJSCSdxOkk9yoUhJtniHanYGY52pZmbLXn8qWwxLwn7dP3jyf8IVN7rM
nIyg//70e5RuVJKzQDJ5wJ+rhDBEG5+bStqmAYzPVf5vO7IwW0Id9JgU5D3tw3WzG4nxV6SeIvds
+zeocuYCW3zZ5iOo+HxZNM9OjI2ugB6MeXQzGmHbmrqj3IMSsDBj1ZSF0W3fo7jnOvI8Cqm9sJPB
+Ck+04pmkz9xHJWfmyczNYlKqQucn2hhyxol3ZnQez+6YNnUtC3rQKBBHypCr8xjB+pByzNy4gLv
wv/rfp6xif1Rds+CmCw5YUSyHPAEk6QcWGWCJnqpXzhFFNFHiVGKzwU6P+GLs3j8Z1d4rs07kS64
vou20U2/amNcoifQFcYoPknAQlf+uutVV0fO8qYn5MLhDiU2CJemm81NRhnMmARx4Xz/7kKDKPpk
FdVNnfUVOTY7fp5XpTQSsb+b4e0nwymS1KNzwsKFChW4dkzG8RXnGkQhgkt2isWa1UvlBqNfOduy
pvCfGqb/Jz28M1q6ozZqxaLcfSthjfLWvSoQYQnUUJJN/fOcdb8GoW6XU2gYUGbEnV4Ua20n3CQO
xn1fnm34XFfx0tw+oOJi0WhKgllcWjcWxB1FlpNaYS7h8JqBqPw0MjdccGXxKHhKWyh/6gRrB74P
ozsALNianMM6mf4rjI/ShurQBT09UAgc/xHp/KLwK5LKAnVdShU5c7EElxrc9P/jhnDSgSNz3vyM
KR6Ovnq6M/nYT8vY6zq4KuO4BguHXpACa+HJQWXnnLpJkliSaXBWYOoorazMWdsu7C5wWofoGMkn
n194RXHk2+M8GKTdW0RZv2PUZ1Eo4SHlUebGA2HKlYmWTWQHdae02l1M/HTIRcTZrw07sMZ5ioQg
UJ18CbBaBCTBwnNe4WRIhvBbV9Bq5/fXasaO0gqPGevj1gIXTVhB63zHVOuUi7D0Fh6mwO+kSuW6
Ji3BcZ3BC+DrHlEpJTMsU0U4Hcey9mEf7jgQRn47QnYoR/YmBxzd1L2Hzku4/3uYF4rnxKtLbuf3
2OZy+N0YuMguP6vbkGlRxwn/FLMSWbByK3scOZGeQsay+7wAJZKK3bZHEFSaI/1KjTbIj27Hm9qH
lqMVDUMqiljVmyA3fscEMp8xxCQr7ozlnG0yhxOUxVIERlrIvkTL4qGlc9Iy+sR0b3/+nXrdlT6d
6tHTHaSU9UzZoIXSnRy7aIPl6hCExeQeGfPIHpFar1p7opmrMI/xSArS+YUVpUcs9IgxJZTOlrUl
SfnzzieC3cGtXPPFvbSKQ8Cb0Eo1r2j2d5FZa9+s35VCU5crVRs0LlsY8AHMdew7kxFyMrYycSbD
L5iKUEUjhO/c65BkeSJxneN5mU3O0cHyiDBZnEVUMqvcgGu9RlE8WWQRMPqJEoerYnJ/jwhmMMen
nftMihGWgW/vwsQAOMv00G6hhKyUt0LfKka7nWFdw0ws6GRDYxtkwhBXQOOXfcBa158KieI7eaUk
ydKKrhS71O/l99y6FBo/WAQSrQ8EJ0SAIBZZxZZ6b9A8B6PIjrpyjPXQVk/c1bbU0NLdtJ2VlT0I
Omtg8+1eKQYqBVuthycDD7qbW0cXoi9pd8rzxAu4zkWY26PfmtjkzhOHEJkf2K1zcZlZBMI4LjUK
LoN8rZMQELqgglk1+SM2LPcntqf+owqAC5reP4awpfHhJY2fLJFE7jVaaJk2cbnSwYR/h7vHMoXn
h8UPjmgz3WU9Ff+qmyfkypNlcC43Gv4E4A32DdgVx5/XXGVGSnhi++cy9sXqv9rGIggwtXJGrrjO
E8M3RbEf1caYFX+IqUjNxbd1cS2u69O3cGsrUebA2TlvFbqlQfTqZr0p0zRC8I8/Iyj9rK6MUSa0
GpqJmneHJBubRV80KCRCa6Y6EiKXjmVUWrlZcJu7KMXRBTCJ6xwSz3PNodsMEw1MHJZcIkW6x1bC
ySEriLRtq84bogUM0RH5Q7FvHqfm1fuk+WMs2LG6I4Tft03vtKeqybLa/rAHVCayKmNq3RU3/dGq
eUbCeYONhzfmlpsV/sPaTW1Bq+RrgbiAAgAdVLXCCauHESLA5HTKiIwSM1EmGRAh04Q1eEz4XsZJ
cAd7U8tJVvx0vFdcHKLXNkkBBgqR4F6afcHdYLcOCeeB9Flrx+v1/gAUTTbfYouxJTYlWe1tZtOf
UXDEuUGdWq2dA0e9U3v75z1njIVdJ3EAdRRsuTiVu0NpVZ+KBS8Dd19YXsPDqjoEd4Ccj4oRfl7e
KGTO0dTzZrhQVMlzd7aGv+TNVbHExP13bx29fmZSOtPiHlalDbgp+bWJ8qo8cK9dZD/ByY7vAhBq
4G8p6hIfRxfTkWi0F2dGjqYLlEBQsM5gqRsZWYSVGf46LNVrC+WyhOkfVQhyxXpjDYbQLRu2O6iv
HW10scRj4G56DC6qTalV4B6aOMATa33WH5KyWXCifa0noixAHPLFXZS5Oj7bEGAN1h6AP/g9tum+
73JJsEKSZV7R+Wy9WKjxyfJEGHOG830xQvxL2TTugTvniDkr9tJsI8WCxDE1nQ0DZ2bpxNPEElX4
nQQgGG9VfwWXxuMgv8ELPpOiZbltrsgHuZNSwd7E2XXcT12oCk3zV4L2e6HdG3NDnERfJZrwxCwn
s99YIyjWaZu0t/qCaarJk92N7CIRz2AI+7clhez+0ozaya7GWnMli+HWmfQtO3L0rjT7A7G7Y9KA
xqAq205rs4DRQyudFvD6urVjJ8BN/u1fQxNyjOivnhgM8TU2X93h7F1wk57fIWnraRBGNB0IHNRG
UR2R6Kq10xoBEc2URy4bhbCyrYZDhAzVAp0YLgUClcU1tGB2xfMmVXwJg4Sj/lPD1IdoaDymrbDC
L06YBdh/Ipkb7cT0L/+3ePh3i2l3+G8esvPVPnzkwhTUYnPZfYeP+6awdZFEDnF3vPKlnz6Gd6VJ
uu7SM+/8SL2aTnQgBBaWqQtjAKfI0SxUGZjfIkL4bOhoTIl0AwwZP7TqEtx+Eh5Ayv2Zy+cqEQAs
mJ0h8j14boxzuMkU4DXJfYUyRWfcsPXQh24HwekjpmWO1WHzQ22uIAEOMH9aOxVY+O1H0ZSeqOQe
aeOFST42QO7NA4pxqK4n3bFafE5wlA8ringsBfNfw1WvHgfNwQLAPBnu0j2FiS1yVakmoJdS8kJC
7o5IVoSXHYCv2GfD/jtIxF5Dor9+j20iEhmEfjRqY8zKApeQ4IP7qGvEAoB1uDmhLaFDMPKVZATy
twKd/QW5F8Nno6rVW4EAb/qWZrJJy6OOa4lwqQjzAIzPw3oagBcJAJdcR/yjC5qE9wciXNzTv08E
IqT5c7bH/BDH/TYsKSy0PaJbUrkTrYeg7xMCR/WSfF+KKCFEVDEaSAlQhqeZwbJIJQS69Vjxg0mr
FHW5YOa1aVaU6TcewLRiWLVqr0lrgJqL4DCeXKN7FGHA9PVdl6bRujAea/yRAlbu9JRBZJAuN72a
gd4BFuKuVDiySJeSIqCvQsGROYWGLuaj4ooyuyM68esD76qJI7NaJuqH4QgbDHLrg2/XDmNJp+Yb
Wn8f366IA7ehH+YbBSrf3n1johAlEH8lhI2ij9kE4k+c/hRGCOyhyn2egy3bioajpEZyZjv04yy2
3ibdOmMWUttZegJ7iGyxALZ+iOQrTkYMQ3y4gABJJdWiVJvPCP9SXOVUydB+uW8z4B9M+33n9aSA
7uFl11uMz5TXiWzew/K+3Veb5da0a4qzNL1rpQUl3My+SEEIGLKr1CqzgB3Art+t02PKZ5RUHytg
0lVi8mG8TDaARR9cqTc0fv8RnwQwhIjenUattQOK5aKAtfU8eG1x3bwya11itzitRoX1gBe6xqAM
fTEqdkRNPU2qSb+21kAvazMJiO2C/E9tNgf8u40Z6yk7VyiVQOixR2EZ1+6txwZ+uiNAx/zDEZpp
bCztmpGvlTOZLy+DUdk+XOJs2FEG/A5aQ59dBHEDnvr1zZC34ZXY6qaldN43rfP55p5/LI5/9E26
YOzNUUF4hv660GN3POKXmgV0Wcz54Ji/MeQPuCiNFLpgcc91Z/IwwRP7ZJaRAV124yW59+uBD9wA
c4x2sZPxgMiVa6R+zn/OpoAsFNHzE8B2VGVyvrDZMVSRwoPMKmzYgZtwrUXx31XA9tkAI62MeXnW
VOdVYAaH/ESsP5BXlefK/C0pS4DqmHTi2W81L3+oFHWTtl7n+W3Yk4enJKN8f+9D9+jwaTycNzTA
sjN1R4ZRTYa2b8lZSV8VPYx3Mr7z2RevhtDOIu79fcEEaHOAss8SGzOs1/SQCvi8Ukg2g/ALF6il
4iSFo2/ROEhXFWenqOWJtm2Ucx7KoP3ELKs56HGS8MClTHTxtqE8nxJW8XN4GANaaWlRQyt5dCE1
RK+cIlrkFsowD6dFua2rKOmJMAanm2JngdZqFi4f48X2TGoeY2Wm9jXW8AW+EimXzVsCfAblMJDN
7WyYbVo61LaFrVNi8RvkHiGt/4mN2GvCoZyEO6K4mTC5jjj3gMUjP8whmhoFS0EA45oRDkIbDwiL
7woPsko41nJkf/dxZgSZQBOATujRjDRBIBXU+gRiVdmGoUlPyGe7LSFTB192BSkxWgKJI2+aBlW+
HRcmv8e+lH87/9u2xvzn2BfCih4X2cbIlgEdlUtDl6RKOdSguzDdgozqJMDNVC25S6JJxNegQ9Uv
lpHZstyqmxMxUJVHkuVJw4elSZQMzIPdffoE65qy7/Nadu+yTWooRVsXEifi+Wz8a0ujArmxI1oH
C26kA/XoJXbwLLIWeDLR5W4Apmjhg1M7ehCXv6OiNGCgZG5rLaGpNBlOG/ldHi264mXYY0aT5y77
5wQSgIGSn6rFmJjXwvTN3SKHA5GegsJYH5fXGYqxND40WqJict1jBTpOrzpzZgKG/oXBtaHqZlF1
r0KjDdGa6AYATom2OPFD6jehXYeFzgff/CK5O0/27RUiCqGazV9PA3Xc36Sb87b3/5pX4AP1UvBl
BblMs/hZwfHT7OfkYLog4EC3A3HkpxyBkSDM/Gu1etSR9jrGz6NCzrgDR4mzisYquMARR2HXlVWo
h5I/m38mkE6jFyQDdtwNYqTstL+OcTsIb6/90AHLRSPsR5WPuqVsN6SAcBphNiQyRIL0lXpTGrgf
+XvYhjuESqg5zxk9OU/NJzuv4dRLDPxAgriJWTYUDJUf5h3MASoNgv7iDMx5yP077NwuWmrzFM5M
qoRD63pA+JYPCdOThBK5WDfJbJ4YZyg5JyI+4JXAkHamRv5Ht/mcCc8NuQUx+wj8aDVulDUy6Kw8
f02hFUCZ6ycZfjUs7MUGfCiFsf/8AfQmi4sPliK2edp03UgN54++gMpEPhOQQ6Txfk/iUUmnTYnm
nbeLq4kCg+LQPpxTvCwHAU+JLQ5k8BhjkEksvrQS3YMksfZkgyqKkNxjbHrVHVfJOoXW9L2D91Tq
aYqRvrfo/jYuB4KjqBlPO/oEp3oVL/OlS/aQO1ay4yOkW+KlCwnMWNtVgl7hEReoRB0t5+A398r/
MxAGwNfD6Sgl6oxmviaNDhAzb+n5ezc6FFhMrTvegXSxlPBbKqdmjVkcv80SU7yVegSZ56NVTg64
Bz4Bs/OurpduC3hWhgZqTTApvNupbKSaR5609o7H8pojo0oyY0SIQRzwRFTwbxLyCCKMWumaePU7
GHiKS2FDwYtiJ0RVLzGHCXhX+G0o22nYvFRkfOqS+GX/QeLF0Sn2qOnsjNtXwozYhuSEzoqIjMm4
cDRUsnsO7WgvJ5qQUhrgR0cU1xuUKLMgR/b74e+PIzPTL8kJbvracBhUUggdeN+00KuYiKnLjHja
Jp7A86jt5YSrFttNwdl7YsDxGFgsvc1+l+bHaq1MHx47ZI/7v2KJNencA7Dsz3G9GDZNlHFwN1Qg
4uRYE1xQpwZyckdpABYISNM3YUjxaIcoqvlq7iuc5PI7R7OSn6AiPLS/ATGwn81umaLvA0WIGyMb
sg1N2tM2ICny8XDh7zukE9Q0A54UHlQoXW2mz+9rB4ZfNo6Nnv3vAhbEhLmEJu0xGVyVeexH9PEr
kFLBvpjxL5COcW06WWJQjm/Ij6i9FyKqcKBpUkZvadknL2rs9s7OrvUtqO/tUUmAncuEDXyy36Yp
tPCemmsnJEI22AebjY+59NYuKE5SFxa8MJQng8NO5vhGbnNtzxyMd0PM2xI2soz8NFOZZwHdSPw0
e+jS+DHF5qwQkw3YDO7kNxjCbQUm6I9tz92Az+k1u42SV61goYYOFxHJm8aKBQXzc3AeGdp77ivV
j9EYlxaeWggQQdqKQ2/WBE1z/lBKgSTv9H7aZS4po8Tl3vJq7CWc/0eCf6MIajjYmzRY0NW7CcXI
AkSmtPFsNeHSvoVmMR3G5LI682iBoRMOG2OmguSfxcqYOFHl6Ft8Mc0O9XOVPMjcygTTne5tTs9O
xWOVhvBJpRhjQOeWAapjSu6WLdRCZISphLbOQlM2MToEojIg5afVRErKRyhMWlZjY5wulQRlxtBa
kLqr4L+BN9S+/x7P0Zr3HMvwwJEet88Lv94VvAWojTixALcK/Wqf8Gts34NI6XmrIQG0SUD7ZoJ6
OFTlbTyWd7ELM7e+oIi0RBAPRIeA44wHqPwmt0Z/wK+aw0hEdPtMr1L/jI/AFEsp2wnQE/b0JuOw
qGUGFho8zMAYV9ozo157cHEJyTwYSoYaYDfnzyAxWpic7Kyn2zhl3k2hSuQbXDYerHzlZON4taf8
Ldzb1v8A6qFgwDg+NjMzJ75F/mFsCZPPd4PFMKjsySwHxqUMFF5npfpGKSKN5W4/ChiJph36tFHP
7dt/jRcfWp3IrTXfskCHQWytdHyGuSplC0gsuwnOBmbkr6MKem0gS4L4FYvBFCgLOzuYfDqx5G2u
5OOnhXsXPKCldNCSgIFqfg0T8c5iR+5aPoUbwGDcb6fXh8t+WhDDhOTSolu06YZCi+1Nv/pNfetq
rK7li8hQFdHktGxnYx//wziFDC1vmyQnH352J6GFlZRfv1AkdXRZ/FCVMHIuvXQ3bswU91n0dS1k
VdBlO0QJP1esv4MDBUHqHkoH4XKe+t5BzmwQoWWbcg1iZCO9Dwj+aroVCpevjcd1kMyv3z7oojh/
waQrVz/YI6RQXGyOfupWLvINGL5F7mOWeKeBE/M7XabkhdJbwq41N7e/JJPwzPTRf2MTEuGA9PSi
flsCBrfN2mXPbmAinkLb32jqG/hzuaXAuk2d3/yQ5NczxCdbIR2MQkJvdgDDSl/RMrklafD8UlbS
5XI1lLDINFMF+KjnBzw1O30jkOA0IO97nInfBXdQNTuqfoLK1WeH3GyEE8Q38iPb/zimrOq4QD63
80Qoi8udDLZybG/rrpKGKRU0kTxpeUSjRUSi2RnzPvTXHpqR1lKi0qjfDSN8pxnPLT7QJEl+poKS
oKHjmE4MKL8KVL0wBQSQ9pSLu+OuqKhA61a/NhvGdwX+m+SE7YXKIRnHXVjOIZZNl/D/loLDJ3/S
Yn9i3fVIQPRxhy9BwwuddONgRZNK+bhVyoljQugFBn3knFi4z/BKbwMQTFEHIn8igZ1fTdSf+2N9
qviJXVEFS7xWGNfhuAFMqG9H2ZhA209PmGduHZel9t3+yLpbY/Wi+YkfRw2UHKwqk5e7n74byB8v
ljr1Xc9C6EcQ4VmxCqAWiHBBz+RxhUclnCFvlldwWZLDk9ta1SxgSsqrobK7LrXX6yRcWnA7VhjT
leKptVxc6H3D0mwiT4S5veAJw7ZjUZKWdZGZX8eQw+FOaNWEML04Nkb1rXgEnb7gr2ioq8cgBqiX
IL/WBzJZCNnN2BUzcV5NlcLZdgUmcyBzjXw9gmCwKuBAPrfVdNA0hX8VEN+QshX6TNI3JAB8FrR7
DZCA7pwviyrrDdAw9bVn8ZEVOWD8MI6x3x8x56oBIt1gUoycZ1Ty8UWqtc4LDmIG1tEpDpZFcYOf
m96v6DLR6Oa2NBi3vfMzLIExzKfUgfyCayvSo+Ph0InGCGgEIL8yYUkjBnKu6/JuvbAJ4ATsNsc2
4UGRwONo4v0TItju/uYbMZtCi0rYK//zI67QZUIxX6K48x0BgeSzo8BOZnRIi6eTSqJvoxYn501m
tPS3XYFvzNyKJPjTagHXuAqSoe/exYV27tzX4lqmVxkuulBWpEVmQ4q4tzRnu3qiWrJVDTbu76Ch
Nw==
`protect end_protected

