

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YeJs3h9nPnCnr3aRxIBZUXmhDS7WeTgKjgxxU15evXAwgLO5UoYuCJb2fGld8H5MyDQGWc8UFp3Q
QS1bcwQeLw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QMDnsLueMbfhPqb347LcBnHgrgkl6fbZ0QORe+igLd+Fn4pMYglXhNwzAsr45PWnZnHEuCtMe3Am
9p5sJ/ms8icpsPjNhMihj0/+LhkVUeJEYGJR6AGOi4DauCIoKWFsirWy53ZScEPa2MEe+a32HUq7
sCpglfzmrbsWEab4EEg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F3FpAl1oCeVkGEm2PKCJ71S6Z3CGasBF9SuzLFWQnXwmvUuKd7HyekhOce1QfyX+pLQcgfmP3XmZ
qpZIDWOrbZbtPCk3pZcRYdM0rjk3gWPTq89GN09GyodyzYH5nERal74RXFzqDSlXYzgzDvsSzAku
WQ8fc8R6wi9d8ZzaPtv7Mn3RMOg32FvlzTpy40zwgHFS17RZjspNh23gqb62COtY3bIw5wgzOnnc
pwYSu+4rxmNM105eSJdh2TJiSEN9+pTEYMITQ2PUZ0OLL5Qstj3GHFD8/78u9ynXfzh4PnzFHX+c
DtImYoh20HOPJeCFpBeWPHfekXHEPhbC52n0dQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lq9ua7Pc8cPhzNKkRvioUx2DGTzaswIzLnIP4rJJ3cLZM5wsk5kiUTKl9rdBpb7G3yE/zCnmkGDT
ZEvIhQ4CGdpOb9ZjoYg0BIc1GhYnGIexWpvkFarqP15NwctZCibdBpj579M1D8fvQ9Xw1j6ILLQ5
gUYJd4OzxaJCHTNx0vw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qzr81pSyvLThhRepJmzjPLJdFa8x8hA7KFKfUSPL+CaCFf8sC6XyXYts+1DRzPvdthUp8ISKrFAv
jy1EBIdnZB3D8J/YmjzA1s/E0S3V/3tyfjjyCDrQgRkpjqKN1zwlXCzBMyGSBWpl8ENwa6XmbY6s
fYy2IxFIrKpit7mWPaxU1OjywKhHRwk63dw93KzE2hJmtDZhJmXSPJNkgusdN/mkZzbIYUj8bMZ1
mRTDgqzRIp9L2zyHSB7GfUn9cIiKtJb71ztIZtRMoFGfKpLMWPUiRhyoCIz55vgxKfE+F3ghCh2A
ig+nnH/YWVIR6bKztafV39mEL7utiMvwk79iag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8592)
`protect data_block
KnZUzGlZlfg5Hcfx2yJVD0W/ZYB+0L7+uBf+eeoJvS1QNDCgLet13DSLUtMcV/6/GElJO3lP2KKa
rz5OFjBTRJRH7n2RWg1kqhV2HhpC98aWNAKZMuRDauQB/v35/fu8unOpwMPdgWpm7s7U4Xva6irw
8swvJ+YTu/ZpwFgLcn0mDOxiUHjsXkj0Bwr3YB3z3QFfvEQn559Cq8OvZ2xycHbDwQ9Gw2lY2Bjc
tJyCDkgYXGbeSD+QNlzlpE+DqsQf2rJqUZFMM0kmeChozIQ/luXPScdbUXnka/quX6miyzCI6xng
MHoUsQ2Nf/NcnRadGMsGPfxz12U72I+XmevqRjpjwUpWDQIKmIfZf1hCB6/IKftujci3bIKGLDGo
Md5YunHd0V3stB3QjFH/c1Uf5K59/pYOj6L0sWvj9RoN5g+8fUWUGVwrs3j+B8In9wYrOfZhzxDG
ov3jDhe9ZutyvEbIWVoR8zozq/2uUkBgTFFpFLvReOod+rys+NKBfgfLL3hDp0PBz6D/wTKK9+nl
qfWj/43d090vvw65zC8/qSNcKg6b38I5xrsDALBt7UbW/Gl5+h167qTZ9J44fRl2RqeuUolrHuWE
IWuADyy0jEttvI4yYEyFRJrv0doVm/3k8v6nXl5Ml4l8JnBuVycq+WXt8wefbS8gewG8ujdfmMu4
inR8ntGuC0Nual1mdcwQozKkQ+12uv7jz0bITevl03JulK93AAhnnKZln9DeBRWUf/8RHg3T9n9C
ecH6ZD/e6iO01BlFnjURMjFCQf8UsEk2nsy3fmyBWz56xKVKRCs4yqX+DJx3VXIFiGWnsPeNaN7I
TfeLPUdgAjXZ2eTfpiLg22bt1sXWQwsrVzVjo57fg4OzKLLWjdEjAYP14wiqUt4Pv02ebl3uO0m1
LkCl7jnBEXSWGYloYkEvU8jLR+woYRVxamoK14YSa7FdqgsDk1OzfdlWcnREMdrKJnb9WYUrKHGJ
iH1DbWMkUz0VNkyujcLjNbsetBsSgE8I8gWPCa3hYJYxGUQgSqjMQc5cTEWoXeGwc8mHfh5s9FLz
2sAKgReTnt+XZ84COZzv9QYl2pLp1Zh8dtNUCZ7c22VuA+GpS9Jku5+xuQS3s8QQOuQbnSHP5Azy
BHnXW1uA0s4Uan3+CUIHIignsxSX2MNXtV/zidBv7gOvfBvuLIVAQa0eESJyVj0/fozEiG9X6z2B
ACTGCpymTRQCP+r3/jk0qClfzf6qUa+Yt5+QEkNEHPankQxeZ86/WK9LyaARfU3M3+Je/zD4/PVK
SToeA54ZiHhCU8mRs/mF2w8yUkvK34gjRKGneDZs1dV8q0YcmSkmO9OuD9XEkie2N6VY5YRcS/dS
py6lGK2kZx4NwdhJeHBOHHFez5+uosqqTfEcgegMN1HJccjz4B/tHb16HTEofk2QZYTYcCgVt9eY
ROWQgco63TQD0OnBEDSoX0ocezLxgCqwcDJAwHkMka9up9fv9RyUvexV2tWmeOvBzaodsPPyv3jc
7REo6GbCGDlxfopI4GG3IV7Q2YqVpSKck0UudjfbhaCmce4dR7kDPRNJIyMKuNbTTc3wARnGZc+X
hZYcVS5zT2pa5VofVmjuF7e1X/qVvx++fSmFBbK/uEMWeJvAGSB4xIdpaA/mwg5fZsm/j+1HcPUz
HJrL2J9q1LeIoG7gDYeewoS1ul5zehnihDsKeOMBDD4FOx0SB45yQC8QLnMD2U/qt9cEdfo37nel
UcMiUUVK379v2+BPX78t6mFAdDWYqQuF3MfcwbDSaWUIVrlY4KbJJgg2g58PJXU8dL9TRztgUmUN
QivOT7kAyxJSaLlcskFOijpFr1lBxsBPvSJaiLYqMKegnw1p8LOUG07Ulr0KW8DVCFauUJW6hP+X
kMuqtp5STaWdLydKspO455sBTsOAJ6hvvQNbs00k/qnIDuXEjqACLcanLapJrAvpec66A8C6Z80O
e2d2THty34GTuyapIzn2LmibVCreLa8h9hOokCiPNXJqygMUgiZcSTs5rbTwJa7FB4EU6lp+kM9N
LvaApvUSm/OYBnjNVvLxV967N1QBBGbM0bAyAfgd9c+aZVj4EGukdT1HlpIT9KerP7ey4MW0YaeR
7UxtYbgfUNLlOGyCwUaCpk2ycoDwlIIT7iKt9TLRrBSICILPsQuA4kMlTXVBFmvMSQ7c7pXrTX4G
wqYoKduvON/8L+khNSDGbqMVaBOcpv83f16ZTnQ+Iu5k63nlmlvB36VklMp2SZc2am9nNyZ75VZS
Vui8mVYFlsu913z5pIWfJEchPeYvzG5psMnwWuQmDcUQMR+xloDIY5Y8WQ4SwpClwC3NfMxFJBX9
3rFvyYAJnBTu4GnXs9bmJ3rXWtrmRnZj9QkT6Y8p2f0PKsKzna5XobA7G5z1fZmtlfHtolBLTvTy
dBv+ZHGyqGwJTRL7JS1eDparQ2w0pmdV80eFmvJ1Tcw4Qpn9NVaEVg8TK5qwA2+bzTJB+7UTcf3D
rSm2GSJ+SkZt6jvvScIivb2pJcK7B8fa+HmBRjk2e3x7zIAWKPFvB0oNbgdvFk+DSXuZgUACBQbI
kEOrxZzl83iJzKeS8tPP37/swc8rTtLDR2P6yFqyVEd3xuuy44kqF5/wrTx1ycRCHNhiJS3Uyv5N
jw5NVpI9R9gXOWaSMjxT1Gye1nO3bdbNHixoqyKpfcXbhjRYRFWPBbu2Kt+VmUis8D8xNJscJQkA
7xI983xylWWex0gjQwfWbYOfd6LcBwuMEKlYTSeLc2JFC/kVTolm5sBjvo0NSVptN2RCYYYFC5N2
FRI21uhL9q4Sybp0AciENYtUw242grhEhASz4cs/wmh6ojIPij8iBxCJchgT2C6DLFG3oaIbI+PI
OsqxAnizII/ZnsPyzYPIclufjBpeJNcqy5LNjtzQ6L468bxvL69BeMjx5uVA38K/ZSrEYd4gpE8u
nUPeQm9IYZtVlrRc2BDB17TBwSxqu28Iv5FnCFTYMQkstgwgd/zZ4/HOnZFi9EMxpAKDe5sdSD3U
Tf4MyuzQ3S8t2EIqE//Lh35PToLB0n1Lv73li9BBnWAPaEB89o43dS4UpRKrKm5dmh3RUFBI/nMP
Dibon+wnm72DzJcFM2ogr+duor8NGZTMM9aV/dOv7R79LyUZPxmfMQUxeEznjMwmCWF+6bkLu5Ev
i9LH1gxL97JxtYgkMrARFJELgYxDuvSY0zSvTJPbU98mdpMsCBb/+lzEPZowBQXtqLDnbQXDXRtH
cCPAbsIq7uZy7bpwNNDIRPJB3y0tvmLoQzQqtc12s4lKJHYwF0AYqCoJecL2U9Omyk5UD+Se5LJT
0wVYaB2NdgaHAz/APNbjN5aL2m2AhGGC6H9ut8R2K82eRUyhhhECAUUgmLWK6fB5PbYpkVdovQVd
l3tpXwUqhfLvw031yztk8MzHeN6oM6UORytOFF0T92moVrEPw6zSMB8Z5pL1JrZYS68p4J+aqCsl
B45nu8J1WKbP2sPvwr0J2toDqW+BerSBJwIr+3HCNfAvUO+L+Fn4sMqd72iioUYnDxrk3s6BH9q9
PXs18qluTV2GVplabG0vy8dYDVa1VNla5+GohB3F8xWR8Bx2/ZAfV3czTDtYaCySHjZD366BveOG
586I72ywqWyZG3jH82FO9T2+zbJpyUnXUWv2JTiL3CEJthEJqY+vZ1O9DN+TGVcurRuD/kq0+B3z
hlVLRoRIyXEfRImMH6L11pEhYAe2lFKiq/iRLB2dKiVPFUkvVo6oYZb7Ne9p32gIF0421riUmOjp
SxayxF6ad9g85fqaxY4n7xf4CnbrVfJibj5BFhOYje4p74/xDFauQRJZjOiilbgGU0JjrGcZrHxF
BjanuJN/iwKXKdzLDFgH/mDBUSDMa8PqTSrZIDTy9LWePCu4CGuZYYdvGLZBcGCfyKVce95104b+
si1sk8QgRg/TR5Wl++OVayraCnx/NCKoTSxnDopNJsk6tyZKqDXlIZcWinfsi4FEA9k3Xog8CdMs
MdfB134uT2yYar6xSb+xLnrYDAbF4tJxPuc4BXL64OxQ0ddbzhSyqFNhFV1H0lqGbyV72fT6s8L7
EojONq15bvbVFcikGHs2Xt48MH+sfxcUqB4srKWRK9GqngU1jQ8Q5HgSRgvfzCpnfR4wsNkcL21p
Q0VZ8iXdrDxxqJFycsizcnxBmPaBn/r22nJPq9gPZONsg8sPL6nmTJ0kis37ostrSTQ2wWO/yCri
Gbq4bUs+YunugM+MtQqgO6TM2Tcid9OAD/3WYkjMmdG017pnNfnQpsTfp4/38ELT5EkrV7PUwJHL
2qnd7OCPoVXvMQjAOYXgRnbxbXwXLu9okPnudFV0+BNCf2sZfeW4C4GzlezHBMCfUizDqftk7wwW
MpxAxfxbeR4057MUPTtrNsaECl+Ctsah5DMx7FEE6X7WAEwS44BhiqCsyn6C/NIosMBPfUp+VGXy
+d0up044IkRlhV7qWnXHY4ctKzhSJKKvR881TmUf9FVkowPOTgGZ/8n2qBf29Mltn4IonGX10RCj
Ezw9O4eQWk0oKOqJXBxpVDuzRbfIejcJ36BB4fXGdKbuiS28XbpngbDJnJRk+OzczNyrHZjhn7Mc
SFqWqJRdV3Po1W+Oe1ajKTwt7pAGQz2SIe8aKsZ6mHSpWauMqPj8v1yYA9pe+a7eAkvc/8dUvoPF
gEys72tHb7nTIkh6MX7GSs6MyBPJe/y39J5hLLEUP2fw6pKmmLLmSYALlzqNz4XVmCbz61GjaqM9
8eJ7VBuQo1ls92qAhuxMZyJmkEarDF7BD1dJboI9TghUsc3YQ2QHU3eNElBlC8LF+K01cepnj19x
+2czjGecKuMLEdb9JEsShdkZnn4vBq4xufKsOAvb5F2dLL9fCGMrp037hHuw9yBhsRwKzE7XELUj
U5XWyjIbDSYTiu51FCgvL8Zp89CiA1ZgCyPC+IdpN75Yi/9c29engSCzK7XlTa0wGyoB+5G4TZ4q
ehwus9mhl+kwTOCZOHUUip4yVtGp3SZoW7Zsvv2YNbaVWSj/hBlszJ716C02u8TjuBlnDo+Vr4bC
MeK+q/hJ/D7yLbxHSyTSZ3KmyQ040Wpa1jDxT8DD0UbOeYs0N72AEBSIWx9A8y234zX/I+cAQK3t
MPt8Fsd8XZhL7kiKLCQCcG6bC7mfsl8SwAe7MubmcHufVXr80Q1CvJgA/jng5Ga1XbOHfF05Qcz0
3mBwcMYA3QdmdFtETvwLbTQu1rzqjbnP4bmtqRLgKq3NZ0CG4Uzm4+rvx0EHP08Jkneee5xpzyLK
cSpIO8ebp74KgaHfG+DVMCrLPzD+35LnF3hGr67IiSthSDIK8bghJh55pQlpviEO7YB3aXpS6RvF
IOYbAmoJM+1ji8w4jcq5Kh8QktLZcBoy4oByd36+wgJaZLjnUCBeAPE2s3twYnMgOcXv60qdN/1A
46JCszvtGAssdvZKFPXVbffPogikqF0q82Ujl62VGzwVd4G3CrJ9I+4cjnfdeblsTcZQbyZdKEUX
D/nGhFh/gy8qs2NcQIBYqh2k30rbSok5uRp0DI0V3S/eA2iZlsd2gCMeTz+KqpMHPot62UKdnjcv
R8mzGpvdrg7xLWTLGY2zPGlZhGoWzDWUSHm3u2FW15Zg1AWw5edwkoG2xdl8+4FYckDYqF1+VUU4
HHzGk5zz7QNcdo+0sc3YFb+/pf/d9D0Ts9gkVA5BpLJD8vRTMnfnjiGH5IrOhh3fjolNeW20cz6n
auBdXZlM3i3YOhHhmueDSaFRct9HN6830xHk5WJbvkuqfGLVgfk8mLjempJKX3HmLai+XyD2MZFZ
TQlrkvRn7mu2vnezpDVv4LzpLt5wJSlN+l1nMF6QcFV0a/WGxi84TXRyg2il/nMFtEtYgbINxQdF
YTLagJjCc6ePslNa09hy42VernlzbsK8474s4fWJqfOirWM9wxuBc90uwFwkTy7AzXqTVMf7my4C
c8zK0GI8QBytWcmTJcVrQAhG1cZP967JvFX2AhrZTG9KLwvQ/1I3ioFdicT72kg7URNe/a9OTYYk
FyMBqc7/2LZZfWoLbdIf/FNUnM6dDMrg5riLdhYgxBsrI3hhtJjGrwzavc/G0KlMYSonSfMXAU8N
B9vJh4o06++Ycuo48sKvDTz5VFg7UMiY95kEplGMdv5SEVgZld4xZbyBw3d0R8LnZe1F8B8KvitQ
ikc6WYG3dY9E5lqHSNfM4eLToarakIzUmLsPgv7A/aBJDq4T5qNr6ssCWSjtY2ZfmAqN6Rdek010
5z9WMLGzjoMvc6nAnvGlEkeF2RAnVg7pAbfYVCdQpDOjEwu94V2lFktU4tw+YEnXc2nzT/pA88Cf
QRuUl/2CmiNc/wBN5cBi2eY9/zl3QFfeJKOyHbBe7HGEMwaXeXj/OLv79mJY1rtR2ALWE5JiaAoj
x7vOU3Rw3La9Asc2OiQC2Mv01KervoaKV8r3OL52B2Um1nkroce2oqEHsZNOvsq1XrG9NCQrpjgm
g490uG+Lkle608mf9xItpcrUUJYEdHPafVcPXCB5Cbrb4234ptPr+zM45tBvkpzXRjSWFdympJ7S
jsXdiWhSgPz/lONToahCSOKva71F/ay9ZQk6oBcLWGtZ5ZrYFgjX9uzIvWjoVumFKR1+NJ/E83bl
5JHgJA/AUx99DP1qtaYb4Ql43GP5L7JqO8eS7g6Fe7oyliVMoi3T6kjTDE674iL9wwdSHvbOv2FQ
7n9+MLA2lqaryKmBgMqpX1f534zSFGvDPvSl3QITOCx4S212cHB/qGJ4mnatLZXp+eH891KtsUeQ
/aaEGO9pVbG4yZcgTX0gGgRoYIwAPu8w/uxcvlaKVG7IEU1uGME6QeUaiEqQbMYovVBSGVosJgb5
yoGrBNxYzSmkzpM/Gc3Nc2STJGDRtSi6hF6sjeNXWKfp0hQP7heCXVEIaQyAYjJdadSGg3qMsy4S
j8zYEZnK97mtiim1H3bblczbywgk4CA0ysAakJmd0f5yL0FpEZkmRyzU+sin6SlXQVNjy5J8kQRY
Z5nL5P9A4L+5PjU5/+PPBuYtkJp9aMqSu1U5BsROLuWqEFVejoDUs08xO39u2nn5HVMD0ueL49q+
4N6PlHhXU1qKoJ/EuAwNouNMnxzTiuTLOSGlI6svgaPMxs3c7n3BJKpP7iNsKyH+wnO3Ikf/7Q7D
fR7EkqHLbIig5j2ugVQa/uXS3up5j8sEKc+QaiVUkZhYOTFGjT9+gvLCXBwSVcID9/O1v4KMI9SD
471T+/g/z6wCd35ym4cgFe7c0LVWdrJ7gQnIF+rmerOYuYKJv5xj4LpepPTgNwCwX5yIwmJDQXdg
Y1tEoj4r/XCmZGHdGkXAso4CCmhhwsfevsELZ0Kus11S/2HYpmy34nE//LhI2iMZUoLk1p38PTW9
jKOKR1eJVYKRJ/dkeOtvRVDDq83lsNmVhSC5DvbW/7wuPx+eG6+FW1rPc+XX/ZlxsS6QStIW/Lan
s5QlVUmSq8uAs0bwAZZDcYL8MV6Ve75saqi8Hzpwq5+BDKl9fWEpay8GKB1dyZILmscfjQYpNTg3
qEI3hQgNBY56sh1TwykcHYgJ8ZpALD+zrAL1tizLKf353N5mjUrZuvUSg3MGewjshQwfOpwnbFwh
HmMaZajLmI/wP0OKZ/kRNpJ5pnQ4cuWDJvZmfVI4h7nh9Ur3FtFClzTpzjfb9rKRz5DC5WsnXKeO
IF9bI9sokaAmXiGrDHzT4JBQXrdxcVgfanpjEFJ2YjqVe7E3NbS3oo9UPE3+MCEPpz0cpv16nrD+
izy79HHEEXjScjmlogTqB0jS+k5PI0TUXCnna80wqffL1YEU7aaolkPIZc15YAZqMUxS6Y65OVfW
HukzpV5BuBSNhurIiaOINRJrYzf5MA5HDYObztEaTt+J+/mpMKph473zzBzpav1fVgOirI2NuKBn
zKvy1+t7XnGAVZ4/6IsjfcLtznrPmoWtuyE4/4mTXlr5GJ0IIog0hnfETN2U49ZxsM9FGGgzbcBg
R4fq0ELGrtcAsoy97TEhTQXPzgtIrQ+6E14FtnBHweWsB1r8Iy3ghNLXh1DYjcA1egYl2UbByCbg
KOVNyEf9Rf4nRMg5Soq0UrfGXguWsi0IxuGlYORzJsXSTuurwJyDluAlaaDAoPNto1lQVBEsUAh9
IDBrq8NOoG/chiFabrOjZkeD6eMe4YSUW72ka8NaclOExKHw9JIrhKBqRYoHKm55nC2P6qTFnaHi
Qw5vHXlERtg+UmJERTWRMhfZFlnGtCOtaLZKRQn0vJ+PKrnMQor0NpImwwU7qa3te2n9v7fkhp2C
zyTMY5o+igQaDsjXY5pRrbmhlzXPetT1pPAX4Xl0PPpWHKUoEaruURTUBWxPyisiHjp3O6qqtvm1
hDhTEd+sn+lONKekw8a4IFYTFM54ec20TO6oP9Kii/kXiRbPlRUyugjJID0Bn8IOz29eONEvUNBV
cqfISeVNqQQL8KLwstOEqPsqT1U7BvgOn4Xs+QGglW8wO7NA/SjwnJxgkJ6vvciSQ86rpKwPliW7
KwQRSMUzZIJkqp4HybHDR8Dx4hWKW6XKhE9/S5Du3PaWZY2FPr/oNTxnU4WffendrSTjr9NKdrEG
12jy/9n4SUXV87OqztF5HsMbF17YcsP8hIPNp56h+PrRglleMkqo7cgQDOiC8BAUMp1AysFiSChS
UlAWB9owrnYliTo57XlfViPjsQdPqy77LlDUmKTDn2FJQPy5Sq3ICA3/fwq68NxD7azhdrtqj9wL
SsBtUBqHFYMuO2nPXkf2x1ibN9gPs2QT1PRDyGIHB/XNVfxOP0nDbauWhS8LSHII0//B4Pzkqu+e
ir6GNMO9/Xq3uhns8Vs/NfmjoNBAXVQ9P0gPr3AC0r/bkkC0F4NKxY6IRfhtGgq8kLyDJLdeKIVv
jhN3jfhUjw0QZPvfnumqf8tuxTrumYqmobW+cnKnt8qvjSA6MWyNnaPRSO1QggC3KzGn051PIF20
I8muAsQAJWTQpsiDbaT26n2BS85lls+yKvOIlCLiVpx953+R/5GLEt5bgjy4QYYf5UC/P9q1Hr2s
zX2gI5zlFz1R3fFmpAwmNGUrU44maD2cYMnwN2AkM5IZRjFGWYjGB96bn7UuvCVuD90wHfeJt8PK
eLsOl9L2lxXz/jpesN6LgqBlZE9xfrfJtg5gowaNOBYoWqJG5uHLf1osPPRL786tNXuaZMQrhaCC
ZmI0Dp/974Uipb9HKke+1xMheNEaLgqwAvOQUJnb0IIzA7fiw6npnGjvV3lbZsr+xTD9dVEZvY1+
tV76BaDasyotKmN11LasN/abuSmUYk1KEwypm6nRkwZBYis+rjLion7ef1lGt4FSvqi1tV9+Ps1x
+bDPQif3dAjb0LqonXVDUScX+Surr8hOxYtAaig4Pd0pBSUehmqGsHyxxabs1UJwLQu3KbnFr1ej
smWX/0/g1Y2oahMrLcNIghn1EVH2cq4QFQ20ZAUQaFHllHlMW0pA88fmYvhOe56AM1wmJKRALyf2
Z8O4Y/OJO/TraZB9kVs2WOrz7hC5KMj4dg1oFHpsV1Qrt8kkqhrJczH+NeuIuAIee821wAOX4GoA
vWeUtwLlVoagajG2jlLHCrtnyAq7AlIaejU6syuLKGkl3Dv70wk+/PZGBrKfLD2ZuR+I4wXQfAgL
MMjozNxdJttqhlF742MbOOblcmUpX7PqnHAGbaWhKJS018G9yGrgt8MiHhk8aartC3J7yrDtpQnf
pTUr73A6ykvoYMkKRnLR89ilfXSPIcr8tjBkxRg75cRD8MN016dCKSfUHipN/Eyhj1hL5AJWUiIH
BKDzdGm+XEKjMH9ztxYgls2CKpu8JJPUcjToOPfqBY4zCgfCw54CZhRuV/g7Dha3hZXNu145KdD/
48wNJfnq7xDsyLqGwKs7A5Zf+xFLj2pLV6oqUJX+vz1JCpsQDi3hAb8eYtVpSxLEbbNaWBA0n4Z7
Zfh6Nc5r4JG8QdXG4UGT5wsADpG55rxSHyAiDMGFt+qIgbeJZFwbjipf3wBaB3MOUv8LzikT+fMa
486T3o4fJqR8MWd4vMN2nDgy4jMqkwVFRGn3G+JiC7P3QVHNDKj8dN2ffF1Pgn3z5k/oiGBqtuWP
8Vb3UZ1+zCGF4ikObtI0zl/SYtG1gH8YnxXWelWRc3a/KbATtN950zkCvT2pBr/2AxcBYxhQpK6z
Epa+TsHQQN0dhNDX2yoDoWg26e7mtQneGr/Xegz7O/QS0OhzKzxB+1TLEjPOH+ncKSHvc7kVHNYC
jxoZ3h79MgCqhn5Z3PkO0cmRaCgQEEcm4YNuYYGg+tIEn61rxmDBUTIeapzu3yzhn68fyQU8UsyC
OHr1FW4yA0h+X/ivAX0mN9NuKb13sKQinBD6FmgvDSx/vzy2AkrO3iL2xlKxd3vYJ3swCTTMi7fe
dJuStGvv78dNbSNUBuJw0XpUi691SbAS0hFCuiB21HCDwelc4AdpAzGlrccyyXxrxECkC3kS/rEf
pSiRCPJRDppZmLaIqJgOSB0louSeeTJgfSV8ZuofMF5DSR4ZuPv1wRGHmlNhkVT9Yv1m3IL/HaJf
R2PMg4G/Zvb6kuD06hICm9yYv/LnJ6q6mIfJs+lTlLrRAJJk1Ry/zmMXeN4pcSssiIuX4JjlFa6F
z0V3ZAykPrmIP09aQ9U4fqAZNm2+eAgJqvpqbZ1te8rfQUijnLIFzI0qw9WQyqluggO5+4kpT29W
WyZOO4iZorPWseu+g6EfMYlIoAtD3a9qsKTcQRyv7oJFl22PwlewSh2Gx+49e3j7lcVoNlIMZDG2
sLffRYroTShV76xhz0d3tgNCUVZToQtwVyP2DYRXH4NREYb1o2BAh1o2QnmAYa63BeMSr8I1MIFX
hDRFtiYoekVLllqFS4h5dSzEzY6a75jsJ+mR/mbiMS+yQwTiSaHQu3oF97AqTyaA2tS+FmP3mJ46
H32iCtJUhMivtjFs6rAOpUA79DuWIGPn3tK9wj44iLqoo5Akr6kUIZUjU50Bbry1bgyYg1y9mfc6
tXSKek79/nzPmvIq9e7Xmqc+abWYWqZQA36nHrmth7PTGqzREozv03Rcywlj66gYWk5PBG9N/nFC
FSI/ZvY7HRSW0xSdsbvxiqEjFQXd6RV9LZkW1SK8ykd4e9sv3a/BwBou49UGSW1OEehYUtlmHXXh
8LBHlNVv0pP2eT+aXt8B1/9eMYg1yovipXml9PNjTnmUeS1DyNHjz14tAmUI7zvH14kymWKVrNUU
5yB0BCngHMJAMBQyeBmMfSVjAoSTbBW7yCYWcS1J6lrMAXCOlAGfJnNvSy6JBLiRjE9i4SFVrF9C
KxJXBya/ncAnV9IicwnJHLO2SVPEF0Uz9elNb0B+rTKUe6l2eLs8JGZi
`protect end_protected

