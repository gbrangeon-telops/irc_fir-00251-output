

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cIiYfk3Xy6N5OP4pq3GmqGiiVNUZ6H5+UojetFJBvbKolIu21jc4BnJQVK6clVlXeOqxCwUuMeWy
2HOHrYFv+g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lIziGPDmnLk8lYYpZIaDaMbL8fBzq4Pr1Jhh0ulXet+pjCJLyV5jakxS1oSptZ+tHYCT5i9DwoXk
484l0YBwGxIV/F50kQ4mY5SmovR5v/32XWyGw8Sob1+z/rA/iYbfy53jpQjBFTMhONxMl2jPMKOr
8b4lWHN3CKPgzR7gpH0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
htRzDc7r6AHMWLJSZlCSE/9tAboPhTxPArTqmJzMnfBntgIxMOX2YAPT8iZ7gZlglNlT/Bmc3ZIa
nj4bYkmP/Ed/Ze8J5Af7OuS/hLPfbdPEIMVOJrAzPKtgRUGYzZFakpIpDVbTLnXVCXGbnWwhbHOl
N+MoLyC3ep/1xGkMFlPyLgKVegokAfOd/5ePZ6yal5L+KR1ET32v4t5eGaONowzpG0O9uY8LtLQU
iVJDGAf4BzpePmtzOyeo5v68FfUFTjm1d6csF3e9pbQ9fEwJazksjJfyX2XYuUZH1eu5bhyJMU/O
c9/o5sfORhKXoxNo0FDKepouEYzneEXI8uuD0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FHtFxX6m7YezwdeWAQ6jmWMHTTCQ3ATyb5990cCrfHVNkzUwGdq1shf9GRL+uR3C20sVQ7v4/+tb
aJQn0JjlSYvQTO2Q6FVyjXNHAr7wpM4t4p6I4KuMXkNXuNp6PVpERQgKViWQe974sEr/n8wacl6w
0ZeeyAlvAxPvOHeW8Sc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WrHRD4nLu8DRRwrUtiyMH2ZN6Vs3L2kgyFgp5P9DMlNKTdIDDQa1yTQPpciIt64OlniyoYCatBqg
Wt8N5KlawExwntwLmfujXap7EAFuw40uyJX+yki/gczIgekz/25Q1+NPVfIAzqSReCro4UUW45VQ
4oIxLBIF53PvEJm3CGD200yoSxIl9Szkkq1FCyNtIufy0im7xj9CnEg/iFEwxzn8s8Ge79lV+lhg
fO4H7eA/Qsx28fzoVv2RYnMwC/Ln7iTt2527VU0KjrPDX1WGbNCJ5ny6IM/daMbuTMvJb5fz48+S
KUNyOcNxuhu15WGxxGlN6mcj5zB0r8XxgsnOfQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25744)
`protect data_block
TwWhg/Kjsye+XcWSSNfvVydjrRxUioZdbZV5UxK2kbF918GkoQZ7aDEbL72okx6b02rQT2gMjxTu
eXt+37ll9r340RopF5+y8wdkJz6MWJ8AW+q9I4ttySPM32Is4H3enYO4fj7ezVOR+by8tvF6WPSa
oVbqThQuvP/BwvbG47DzSgB06xvcZiaNHsm6v1rvg5LGg7edECkLqEvXSm15fqypcvBF084U4eTO
pGdfwih9Fm9yjuOeXt9t6CjKaiJS5DQ3xJZw/wdGGmtLjMxTZlQnW2w6zWQRv94i2z7/oU9BphIa
7DJQa0DBMqJeusT9BB0zdPuf8ofwIc+IigSmHJiO29dS/Oirn/mVsG9EUIbNRY+Jsgkyrhjavuzx
tLQ3uoBXWfvhTCKyXvgvNZPywtYvOq+EHzJoCcDgtI4WWRMhqtTdPJwH/cs4gI2n+sv5IOeBJMSO
m26+U7wXXhIt/dF6cD3rHHMg7uxhKih7AC8aRYX1rCtvtfj02a5/EEClmX6HrCx2H+ZA74q78Ffi
6fNcdwllI2tU0OA2iNtxnL4Rc0MlAuNYW9AF5CZoDiOcK+veCxI1X3zxNGKpHnKJb2BOmhXLkBZO
nDENIZDdIX+lh45NgCmbtIwN2TW6CWdcMTQUDo9JbIKibW82B0xERA4gtivmBoXuQ02ST1WomgLX
2wknSZ3H6hUamHW1p+AULrOSqlJP4oODbu5ely8ScDIlOFSGGZ+GSI0ycabLwz+XeRhGTz38fnmC
ljMRspjeeubgev1UmVNThxZGACJTzY39VF3t24SP1Toaq8bdnbKJPHLtdtHtBne6ebawNovJnTuW
/fsAopdIk/d3Pqpvg5Joh2+j+pk9zRa3qmlN03pVK0mbnVg0+1RI54LpfIdsthdZHReYbkCeWve6
xLEQmuG4NGEPyMyEfcW7DGzUcIZB3r0Qomt2sJaScFOvXIb0dx3a9DQPcM/nQr1vk7QStJQ53d8b
5mvYvh4r9ruaX+BZN0ZrsAzUTIbn3Gbo4vPXCPdJ90XYv5IOpka6B9DxuQctrJYLiO1sWnGfyE/F
8gFoGkpHqU1xmJ9/RUee0KUr2rWFPS/ORrVruzOlWojCS/tfEIJGBghFNy26p8kcDsnZQiltbqiw
foSm/bIu9J8ygfISCSGkHerWF4DzH4EjZQUHMPRicp4H0g5qAzdsKrtc5Cq9UP6C0Yq1L3Dlrgq0
pOhBaF2tWTgx0iVhot+yTGHr5ZeBZeVVlOuQNSnj3exhQMparhjRAfTd+6ChrEvtKvmPPIYoAl3u
T4N5hqkFzkRJU+mDqUi8+aXl+KlC651D3SJePyUxFw54VKkE7TitmyrapaY1ObKlfLkAzDsnK86N
J+ohkRKfP9NqAw8mUd0Cdg8wCSfmDXoG3rr6fnJtKgY2fnNS76SQ8jKWu/vW/TItQLW75mz2OA5N
EeP7ciEqa2N3Zw/Ni3m68gyrmRs/qAs0ubiLgtQJTtLV3aC73zOB9N1eX1xlFzOvT0yRirI32lJs
yN49/bAxIvV74s7RYwDZXd1WFTKu6atUKuFu35tIS3JKPNbt5gIT4+PM4JZF5nHOzJ6k7KAK9q+M
ofHGMn2XWuUzRq1D8k9M4J93YZSsEUyW58CNK5lFTTghNfNUBKwiMSvQOmafzJO8w6dgRcQK0Fp/
pKVhI8b6K8HEb4BFGiSc4jc7AKQnps8XV0P8EM8DK56RSlkjiCu0oFOIspUZArvYZM48Jx1AF7eU
G3ufkoriwBRWxBV7vi8HRsbdyh2OWRWN5Z4A0whLBUmORpGugvOmMUSGEKia82uRzaUQHMJY8Cja
M8kuzhXGqolwVU/sMxxFLl5fbCZU9n4Dbttdrwhlk/1RyOmCqwhm6T9D+cGIgDNu8qT2MtG74uAX
LB6GSYdca3FNZ6g5nbuWKp+7LGZZnkNN6OcdLrsbZr6FB5FnPyVUw62YVWAP40kJbeVFphbXcEpP
x2N1Aklq1wRFradISB3FkKpLf5mF+5u4Tnj3/uzQ/DeLZFMcj0Pm12yEM5m/LWbAINEIJB2t7lcu
eivmadE1OYbav11ABZ2eCrkPzHUuJh/pnvkIVkTLaaq0hcorGgMKMRTx0NBut1d7EHAXB4Z6h9Ub
43w3xReDBlRFBwPF+bPr2gPkXSIJo917U6ozWQRdrEkJxQbBASmY3R3OlNeXKTJq+FIdZoHdPIdD
SZpdGRDywrhiwxAt6GSQEYcv5rBf8ukenxc5bU/O9PJnUeDaHPXlyBFvVBBCKq8SjyrI7G3M6Bgy
Jawq9V9bROtps+NjwpU7UdLpQKjgOQ4tqB/WYUJikaVpEh2Hfc6YiMRl5n0qyR7M6a5UKBH0ik3l
yfk5ce8qwfT+e4fy1kEZ3bRlJHwNZD5EVboA6scKcCfWNUrVyLkW9IYf/YUqyw5UTTLQvwOSBivg
w+sYdz9hkFI6LI5NW5I+IKGzpHBpNqnjNdsTEtq1HGEkR7wOpABg5SsLxpZa3bzv/csfAGhu24Nq
nUqlM0pGVSeO5tlAgQOIUNsPX3Crmo0jsucFnctmiZa3J60S2xW8kjtf6rTQikXvhcKEiqhcdgDR
k76zemKxcHdGG8YMuyr8Mv0oxI2adtBRDtoTtwVlnOmbk/h9K1tAoaIBJO4UH+gl1r465vj9vwj3
SefwzBduaY8dpNT0Y8BETUPZvb/86ep77rwBzuQlEGn2pT+22Ph3/qqCSB8ztRqVEbRGK4pGTG5A
beB7cSVW3BzaehwtqGBFJaDc09TAnTmVTlc2eXebiJVBxDlAWnZSaJDrqdkVwSKkwHEnV/MwWBvo
+GklKpYqqJ2kkEChvHTHJ7qxFFIFf8+MrK4+nQJ1fX68O+6I+4bca1xIo5B69CTEdhOEoQmrtMeF
o5IstpC9uiWKZ/6nKterV9/WXgaSXoWzJDCW56wak4IugOYNZDU1LawhANDyYxF7K6c+h2UiTmfi
rG1Bf1TL64CgBjNzSlYtQj5hIVAtiMKESX3L9dqLLIp1CEjQcNaZvvJ1Nw0GU7SwExTsV+214cLH
9MFioHko8Yq/pIqB4YLY+QuKYCdohtgloWN2+qIqAaZ8RR+u/dpGb4ib9SH1YkKAWmavBYnrVAA/
yfVL/c2ysRYnSnxXGp9oFOO59Jdz6M1zKKKi7iCJp76rs+XtSGU3Yd9yDfuIgTUuVnxdzpO0An5g
k2+9wSQ87yuyxLN5Bi0jMFL//VonbmxIPXah6/UKNG2aoNqmEFzGJCOrEp7kzuh6Erx3+3MJLDYI
zf22WVm3c9LCP4Lgt0uGGv7w4YtO7cKJZ5x+aPITjp04ctua0kmVQzsz1vN4iPZWqIA5qb29TwWr
eaJQr1sweRkA6PKaU25oRvVkGQI95I3nZidl5TDQuEl81dwwBHzMygzq+abKJeEiUEt0RL3jgqff
5jyeWQt5scCh2O05mfQWqP8wfGJTgwZEW0Mns0aFO6DFwKtd4eX0InhPhmCwffiI+hxSkISJDP00
jBrhjeS2wdRBWgObGjWYfW94OBMb8jcWMS6LMZA4h+ypvTNHVf/lmMuI9v8BcE/bZe0NvOl93vFN
8dGVQ3i0tz9v6C09AZTGolwd6kQSfG5St0lNY53IoeIjLOVTKfoU0VE/9zhuIfVQgG2JbDlROd0e
nxc66i8UF/8uagSObybWdHKXr4IsCLzGk0LuWLghPN2cFWqXWKO3mA3u2a3zbVTBGKsiSInB9pCM
xf1aoSh16w4cJSxx9JqdEjmE9ga3F8dKNxez36b+yJph6X7GHuSuG4rT9xKqrzf9Ra9EAy9LsbwN
DapJ1shHIeuFR93dJvkgzCqqmkJ5enAmTfzxqAnC6Y/ovmJBn/HBQq0t9tKc01o/DNxxOH0gM0lu
2VGmX/ulyUNanCp6EXj3iMnC22u2MbKmFbCU0LKyIXM1zPEK7fVAG32RiOjag+DX3lWRz+4WvZ+n
aCao58SXw/lfIGYbu9Z42rrAJqB4vyTIIrkezYlDlMWqMPiIVKLNDLSVRQH76T+VhYcTvWIP3VfO
fMaa9hj/eJNKVLEvmp5kVbyzRRx5fKKR5V9H+LBjxXgpnYKAdi0+MSiAoEK8pzBLvqB9s9GXIjgb
H8wgonJwxFu5uvZ9nNG+ZsVfsb55fyNO230mCr2Ha3noWpXrET9U81MiCuWJxBzbubmyXb39S2B2
r9Mf5EoGnu1XeYEG6Mamk+605/XRRIuWPaVaSZAUAB8KQUJHxZYXZXTE4AH/Q3AZugTj3NAnEvi5
3QhZ8haISnHkVVQTEzI19CAlh3W967mHv77lP8viBgVerY9aBqtRqtfo+f6VWPd0Oxo1oZTIHlf+
eiRTpCZ/iZh/WEG6N7aLwZusRDd89Rd+bSUR0nVP5CTeblH65S9lSNlFhSCqkfyoATuI0C3Bq6nJ
wS+jRVgds4ENJR5THgFkZZQq116PzakdWYfgR/v3XX7+UbkMuEXYPTIuNAmQq1Hb0axRONNMEbQ2
NKkHtzuOHWYGufKaU/9XTTjQ0qod7ueCW0zK6Hb95EeXCc7boC5ziqo4b+4czMkRXUCT/SFnPPr5
xo9K0f0GHgkrjlKRstlGWhaTqj8cL1j8WPQH29+g5wd1Rsw3aXEdfcMZEXT1HxlTaCDsFGXEcSB5
ZjE6Amfjrbmx0Zu16SUq6KpolWjMzsQiwIs+l9fSU0TB39/g+NFOwAMQkqItqZBhnZz2xjGvtRDi
qwCnOtx0+c5bMoH7Nanqi3ehWvr7Wj+/QwUsSkW8iBocbfvsopRdaYzJa6ijjdYUigg3GX9S/HLl
GZnHcT+aQAoZGiqCPIZm5PRtAK6CB4qY2Hz4QsPi0p/MWDOlQobC7A7w/m7ouLr7F2m5lM31TPBu
Lh6NkVFTf+jrZYUGVCbdrfpP2wSYDThjp3CLsP4zKkhTjte9QS2CGX1m5MEYAGFw/Oj1PxOzcdVm
fatI7ipxdjcqeMldvROo6HR5GUGdT9dwgq+yOAyenMd1kzXnJF0G1bgSEq8h/R/pTgHkwe4g5ck5
LSLSglQy45UNATyQEKZ4aR81767RvPLTkdO5waULGCIPB/Yq3s65/M+cCUaK2xE4R1JbBhCRWNRM
4UusvqfsqYKJ81sguvYso7V3kIZ7pxNZef/to6xSXmGq+Mj8U8fjzGk/xfCRqMUY1cTt4oRmP9h8
s8Dd2kXhbgHIiBVJ+HX54cmBgONgMtLnJImrM55d97cjvPFJLpJZEQA176UPF6R45lkPA0IjPaBh
rw5rG0Mx12cYSs4cgFxAPHP7YzjGUiVgKj9t21T2Sn+OoNLM2CDqqQCqMLcLeGQv8jQQOLCBrDZK
IF2ypbjOZtIRcWtKo7oplDJ1ybNBx1kdfHKUW+pqC/mZJRP002HCQ5z1+OGnmMB9ThBBQPh5xXMd
wsHn9AdPKOTFd9V5yUeeWX5oH3N70ClBRHn6bzF7lg6ORFNYFhNn0HIunsXHsyS5Q0SNsVdsDlqy
oh3SvLLPptp9tmkzl5L/xfK6g37UJChbQV4ACfdWDb7I5x2vk/3diiTqJvAaK5A6byZMb8u2LhUD
WIayrJtJ7oiR6XqwQxyxh8Bsd+uVATsLbaaPP+0SXiG/E7OyFO4hkt5f4RK0d3WbChyR8FlvSrUh
F+iNrexCd2R1v1T3/Y8ZWkHmg4UC1vsAft9iaLSCqF4eBTwQh3tOna7MZQ5u5DExgJ/sMWp51gZL
DWnfT6jP+rlEPNq9yYtsCaURdmTjCWQn5K/Cl/Jvcdr4F34wI32BDLoRx6XV3qBpY7yXEp3GyUfB
ntHZK9Ba2Tq7JY1dpYwyxUKwmZHGowjuUpfLy3Z4EEOhCoScM9r5+V3qRgfL9sB6AfhbNDDTxIH/
an2oZ/NBQLElFTDeoHzd1BgOhEhiJe28uB5uLxUcYsmVWd85p+TavDBqGAAUpAN2HoAooYf6m1UI
gBHVhUhpGttAOYb6UGZVdka37GtVPPneuBlWldwd0Ly3RLpOasNwkmjmNgIHdcl1+oLPRLl6b5d2
fmtBO8nRVHBfJTecLRKcpkhiueLaxzmuuwGXDwyozBidzobkaXrVqOm3mKb7pXzcadixQ2b2h478
ohnPchkJGSuV7gHCTtleJ6NpmPjnzSBcWYBDjMhilMqGVRsOTXQcUYUBbRO4kxWXwALBrToseTXj
FVVqJ04hJSUmcPHNcv0yykHrlm+LqOUtkbCK4slPp6FIlnngQa17r0XxyKVZczwq85Xvm5cuNHzN
YFtG0yS6Cn1JMeh48JCvKDmhudn3+j/rJu7VXHPd9e4gVrccC6LxBdMEOoTHUVrSDbgE59TLWSQr
7Wf9lBvcxd4WbLXygOU2jLeqB0Ogjk2b8BsyF1Ds0bWnUbuaJsCAijBd8gznaqDFmuGChv6pgBHw
COF8NLThGrbUHwcyzV08ivzSUfMUzAXkWKs7bRKLhW0FYDm0ISDn7Enk0K9Ts3PWglor8EqfVgOi
r4o1tJ6Tw3BsBEjz4g/D8m5fyu8s2etfMqyzA3Dh++af28AJhRmDQINOXS7TkhPQI6MPCibozsgV
aggDS/x5h+XEIksm8G+7G2T1zSiTaJec/eseJmMXwRavkhJBgnLqHBDcxjloaEKZ6kKTezxeXn+g
mqTGWpKVtMowoX2C2jtOIkAxlgu42lF1hxRyKawhJLE0EaIOduN/JXZPtMIDzWs4E5Cm8xatQXS5
0hFgMeWBLnumlTl7v+fxxDhoYpnHepQENxVqQCLR+Jmx6gR4YGxd3b93+mVBKc87ppgN9vs++Jr9
lJSFsyCSrZNiAA8IibxBujbpR9+gOoWitVDRlYGmxj5un/JZRljvOrGT2pXSgcujKszUdQ80K6we
583kyyOiX/TuFLywdMcCqmG7UCep1FpqURuZEQe67QoSRk/xiUCsHlgQLimZ5Rsdgx8t9VWFE1U8
kv1LRdbjuA8V7xWWKWz66BtSSGyV4MWMHn8mGl90WBL32EPtzJtz9JQXUoPeyLPEPNEKnLkAT9H2
WdVDrVvk24MTBArx1GeaiKjBWT1G9jP12sQ1AhwTb1XU31B+Ifq7kvdC8E0CxLPe6csyO/imzlXO
PxtxeWZFrZMZB/0ff3UFLKqHkTtZSNwpLcCYZiWSnd4BYNCZ+F+8kwQJk+lGTDEb1zmu1pdlBix4
nCRXwKgpgAv5Tq7rAh7wukmAP/cUGb6ju2IKXpQwRBJvei7mkVUHy1TtClUSimGfVqZKWFWkvnzO
JAfOdcNW3TfDsf46VAenXIIqiKoqhtr3ayONVksu9EIlf7e/L11qyrEgUqajnKLGbD/VU6f5wt2s
jcvaugn7A+TBVhDuCvraKfio7aemuwH+nw1z96yWKyuqeGPmdCvzf4qvKSFJLt3vzkXPaiPBlR+Z
kKfKHQRbUjvZgWqlKbJcwR7vHLo2yZLBh/mEjdQmY5WPsi3UmzrJiWqUIyh0q709tRw9fLsht0E8
KjKR4eETg0XLCGVqGqLG0+VFsAvqv0Q93B1pLEaRFN/YZ/+2dtHRjOec1+5tgZlrm4sypwR5dl8s
Bt8wE2Xj0x7F6UnPCr3fwY++lifdxZIhJEDe22KYQ0nyP16+ygdcKh42qFRLqGjh3AWCVo8el+qU
cY2ZbJdtI6s3Fn/PN00NBrSrtfHMY4kFYezBAT3XDXvz6z5xHfIrCC9gtrJxqCRBcy16N03och7R
2FXEkkFaCQzwXCdZA1H1G75jwbMUwMQqeaMw6YL8N7SbSktt3rBJH+rT0ZhS98zit95IgvR++i8t
nHOuDdCOUn70qb/zTsJ7Fa4WVLGuCnOawu78CrXsiIbueYYzeVGqBEmivZiUiXhrrVYca4+00K9Z
mVwPhi6SwMURY9h3umbgZEEGH9R69P+foSYYIw55Ry55Y9MwORZiun4fpA0PLSkHZv4vhO3RKMce
ymvw2WX83ldzPoHORhDpB3R6mRxAJim5SDcuv7OdEJ1BRij4AWddJwbH69/GphvfCvBZ4jTJOdPV
cy1L3jQ0SpIchTeHU25jLyye8IrpJ55q5i1lLiX4sQVMQFHecDKJryfR52a0sVRR5AWR2KQAT38F
SFzKgH/f7+nHgU4e09My5Mz1JshRkAPnr6mw09SVruHmCqRkCp7yMm/2sXNYd3BR6F+V+lMtAozQ
9XqZg67q551g3kSYkTca4EzmAm2m1MEc8vFjlXG7PrRbYsZuxQYkDtee1yELDzqjLfVCK3sGbeeH
+tgPFtI0bVGqg+fbesm4DYcFEWr744NI5PtUP5t2K8ASGyp9l+azbPW2fBhAIKgOrGE4T4o3Cs0O
9ggkVs7Vox3yRxuOoYPYZLyJtuTKxJ9D3AUTGH111SQQOlEDLzQq3Pda2KJA3xfCv19pVn6dMXwT
gSNgwKYMJg1bpUAlxQN8tUbfDAIgHzmyF8Y7WYrWyh65LTfMxAtAX+dEOh+dx4L6KgL6ve98KVdX
WyB5KBb37PG/oMso4caa0h+cGUSziF8u8gsEt+kImTBAeNJ7nwzrDgCJKeKdibibrE6iYhnZUfuP
eSYVrw1/jQ2nzu+ogdfEHECPLJum74cUoi5f2BuUeT/1jke9LG01gAHLFHJYdNm1vlaGqUImpuI+
SVgDpoPVIJYt+wP0L2eWX0Um6azfZsYAZEfMK/TbvFE559cVrKY8Ou/pu7LuGTnxPIUUGmtjDjwd
PCS/r3baQDZiKRtrdTK8nrcrVV+oa8Krn09HhY3Y/pl2r8d+0qtYdLlK2+3VcYH9YDksog+aDZyu
zs4GmQUxKAouiMhkf545ccQLHqU5YWC/SjVoVUjpCwAY6UmZCx+uGqE0B2idn776W3KIjp4YqyAF
05caQQxwZXeekCOvvkgXgjPn86B5C5Lk/cbwcmCtvyY+5ZGLMpILbundRrOSitNS1Nv4lRyl+OWi
N9/QjQmCxWar5OXYnkSirL1ZbeGG3UrM2nVe8yWnzvOMOtSadN0kZ+EIGmcEC0N6cZ/UjoxUom/N
1KMqb/L5yTQDoX0ujCRMHiGUhETYM+04E6Yl6JQ0Q+Y2FMf45sRVBCnQFLNHKG0rvDW7uGxvBe4k
nd4ITX2rwEyFxNGhAFgueuPRZcbNR8TZQMa9j6vDuJAZIBx8bcj0fiip6YRAKE+nvRUqx8rUK4M/
7JMz1dE3VyqLPJbLSs2Q9H7vO6lsi1ZZI192+joRJs94UvDAOSMdCwHI8sG9UBxfoOTPE4WT+DDb
hX8soWug+cy4zZAhR5Zh3Qr7QeGIvlqorJBJDtf+haHC6Dis+XTUAcumPU+G45Gx0EkakfzPiWUP
nZovMq/6KuS9nNBWfv0RkDuOe8z8Ya3+ICxItRFHLg7qCTtGTMTaIoi8AemalRenimQX0E8jIz4K
jRl9PAVpQxd3hRvKsFER1qEczpVBG4r1q98y/ArTPtY+Q6oPZYKtOFtJEbITxx3twvI4vE0R1M97
A7uxKMluV66a90ounWEXTw4zikvCUHMiBQh8zTaQqc11BK22dAOcNRha1iceAQR5PzONji8w0Usf
QcSwu6TrmU0VXev8tdGNKjRdp8I9nLR4S9j5Jv+5JlnNg4Qf3JBRj07LTgeTFvAx68U7JrZOzYys
C2fP5WG6XFcJldBDAJgxQ+R4BD6kFIG4F0KAt9suXj3jGUzG+A3Y107wAc3ZRbn/xaQzIu/rO36P
cltGeyyMV30OK4aM76E8W+5pr5IMGsauLNY0hDWQ+9mRNKQXdOF18Vn7LuNp5ax2pZX7URH8kKGr
9NsnB+uBXY8Q+mpiiFwlRZ1CBll2EseBM0cy1jG+Sr0UAbpT7JJbEW7RYxOClDAEl4YfqfN4dEZT
sqktHG3/E79wp+FYYZxppy5ItYIZuiyirUcUSenJzxBgLAYKCinFYdX2jkHUkfuba4U3TCS7fU+K
SiRD0cKt9N+3gGS2d6eObfUdV4yRXzJbBzBrepSA+gHNehnT55e1CB3eu0QxRI8zDMJkbNOFp6ot
wX8nH7g6n6jeMWnVncm/OfK/bruI4ZAtai18cbKcRc7tU0ck8ThHGiWOWy50pWKy1YyP1D7CXTUf
29MaVxMUnQEYqnyLOnd/9V5cgoYoUuGQ4S4ZZ2M9MQsbX01MwEGeiu1uca9Bq72YYD2E11efBZeN
izvVn+aC3SCT+I8dgsdIi0RNFwfDoAQPcvlKvXddteSzC1ickGxV/1qZJk8PVMxpdnJsK4TfvWZQ
w/vmbbbjHOKhEnN73hqdt3npX5tjpU5TFu501+pxXXpIUz6uRdquEwJfW0KSzwx8jzEWnMP4b1wa
hw3aEsCsv+5n+fFHCPLKmoOumITdJtmX4m8elGyhHvcn4tbX+H3J6TX2HtWtGl9USkPkghW+AoZJ
1KaWN7698r8vReQgVQaCzvkl3PM+8lz160vSCIVLKAbCZyned8BLiHBx2eM4v/Egi8wgY6KiuYdA
AM8o9p3el6M9lacl1+qO9oT0RmQGBD62OCWncrP75tlmfK/ocOWHn3Gf5ZnsuPLiiDS0f/DGa0d8
l7GhljT8vUG7NKhTfPadxyuaISEmGuQLzpeGgDh/jTFfesS/A91Z/XPfa/Kmu7sjEikCcf4aE2go
G57GGXaW8inVbJB3WgWPCByJAOzC0FhVxZ7IeYU8mqZmHKE+HwCz5EDePyzdHIz5bkJmUkrZMIQ4
DmEbroV3H+/IHs3TDytobNV2neoh6kiR9xFnr8oP8d2LgX1XZH4seMjCzIMQzSmH7EmlHtUvOnOj
HsP67uXKV4EMi7FoRVFEqmN5LMjc2QyQGvOV10w8TJN67vXftDCICjeUr7Bo0BrSrahG78f8zeia
orySf8pua0GML9ti9p9QA0qouBvr9bQM0xspOZLyTafIAhmjzIssnMXCs2SyLoJnfaGxCkOBvsm5
fPtjvyDwNJjlGN4lZ678Mpo6W2TEIvKQqjoDaTcuVQTMHZNC9hgHZ2tDg8OTPNxW/Vpi/EMAI5ks
STp44ROHJ/tBjMOaU65rnEGGZoZ4x7R12Od9OX0tXA9SVPCxMjGzYQwzzZRYQzs6ubYYuPDq77Kt
P8eu2jtn5NpYIuzq+yOT0VfS7LZ63gEs2ylJv78e25zYVZ6zbIZl+oZo6vpNK9q38DS/kdcZW9IG
6P4NdJOeqohMDEzxJJoZKs0FZyrtUV/zIJtfkBphuK9hbXk6J1f/EBvSaslhXK45XUjH52zF3YoO
O9NXTO8VKbl9paKlcEhhK4QUZzrEyHFsWAA/AFEqbo+zqNJzteYy5L3e6nU8pAue+y52ufXdPAly
pD8JlQm3dZtZNKg2WJOOW5ajW38BkFUDhSIoBt/bmKe4dM4FzoD8PGnJ5DR2uP452/liSdb7k35e
IQRiy9rJH3tLsM1tC1rRjP3SLEZspHRi4+TBa4vNmk8u1udo1h5+NI1hNgDiqjyXy03cOczR2GdR
r62PMioXI0n7Fq797bn+51XPBlcMNtC9ImFfwavkkyyYpufdWQ+001xvT9ure3NZEYbGXs0QRnMl
KV47wq8o/lZz4Zsd8mtGtWPiDjUyAhEFJWBtXhYKp/OKDH1bb8W3/bYfe3YkcnoltlAt2VLKvibi
PjAAtMNv+GWS4oMXx25Is2iSKwa2XIGJon8t7xw2F3HNytFZ7zqC/K4MDDfuJqc+TQVSX6OTvMFf
XC1oWCVGKaZMknqUuLDtb2EeGkTtJW8VzCGXIKDheQifEZtdbDcnoPhJlKCb2q00QGlX0wTUfDyl
dmD+0TWij969UuiabJTTRnCXFszB+vvcaAXg86oJMXyKgIJWBGGiSzA7sW2B0N5diiiZjDHpcgDn
JtE9MQvL/OHU3kG/1n0FhQZBnE3hGAgwy/o23Pc8gkyE7VXVOBoXQN6MyG3it4CDpl5AfnZykXk6
5O6peesH9k/TOueACXG6xkOCpi9Hs4kpv3RzKvtucSwmJStrF3u8Rk734xwE57eDyZF9QTttY4lX
PBCWLGy0Ez6IKVS8sXeoh7sfp8zgN4BLdHBX/eldv/Q1RQ3EiZu9g1tRYk0mJmtPiZngUZb/hWOr
8kjgCwmQdip3jbN5bfPCZRjddJ82g7bvc97wXcxaVAALBWbea3smdtkWwel+46YQCrx06mckXLsH
HkU0BBCLuVYVjDw4mnzs/kLqrjVYHyl7Ct0rktPdCjQJvFE/r7NxDN7CbQba+qECCc0uaJ17Z13r
iWa4mU+dycrGu+NqO/F6dasXMBTIYvKtfj3SPwieadP5AC73s8mW42dQbdHqPpEnyCF7q0VH/vJ2
efvHspF/gRUmOi14YJXZQZgYllb6JrNvLHB4cnSi2DV3CkeYVRM0mxhi0vVEl3cPffBYgkT2UmsB
2DkkKAxz/CssF7WnHt38SoE+TRSbp7WtIL9E4vM3mawK+/ioAH8AbvwdwfpLrEQC/I0He8C781bq
/yTBdHi+LI4CxdDAkcnFf/ExdUU4+Djg7bDUubB0jijK14uOOXXQe/Keq6V4tqXyum3zTFfk14C9
YWsRY+Gwxtbcu4I6lQ+q9zUMNs4CfRDQmjElaOzZ9UdWso0VjS+x5EDalhstYan7JwNBQvEvgfni
EhRhx7VIkhuVj7qe6XNieZtgV8pD8z+yb4uvdU4HBqNyQ+SR8YlTFAhrrZ7QKQ5vFEFIsjfKkhsv
RtFEc+d1Vxm9dR1jRD45oBQLNEWJDBzGePzxMseRM+4lS5egi5XSNUVZF8VnCohBNKLfWl36zLsW
SLgZZ/3BM5N+XokzExq2yCP7BUNEChPM+vCFgXzaWCSFDLZD85TGKyqsapJTW26G6zVMQjt7hpki
MXkU3BqZ4K4VE0mzIh9spbfIxzeEajatmfjEB5Rx87whzXtw9WJmtmnJWMUSWIyh7BUPu1egMfc6
brpPv5Ds5t0GTaq4xvBKl5RGzCXoa6llHDk7TLwlk/znba5QAxUX5vL6fo9Db945VpEH8V7BrYCI
xyg7C3aAnybsoU/jNZP+8FZc9H5LHk0J5T/5Oso0SFe2ONL/4xad36kcOmt4hIShjTfNBn+tKx4/
DZIvPc1CDxY9/F7rEW8yI1eciCGOkCAQqT4xsBRLl84cuY3FpJ137TjeKDxlAlBi97vjGlpDTa/c
SrPt307jDD8XT8kXsqAbMYsUscFownZagcvN0Fr58VwyzGUabQOxvjoCSpFdpsnQ1RxXGax9pPcZ
j/hpr0Oz4NwJZ0o4LZ68MP/6HenWqAafdU8EeuJlq1q/m+ypUCTz/5zX4RPo3dn24dXUeDMW1O02
CvSMZu4ahKK24sWWVXoOynv9r3orwpOL7ZUZy8cipry4xW8RMO+VDtoDhQQnUed3BNx3OmTYpbqy
vicfoiMciihYULHIEBV8ykBD2n67TtbNy2x46eunQj7S97LNOz3IgpA8DcUspHNTB+2wLZJhZvBW
CMiiJPOXstxpRPVYYMOiKZO1wCEVOb8d5OUlsG9GCfmfe8zS1TerMW0dgo3gXWiLIKeRMxTDtb2v
kB8Nkj7LdtOZQFdV5/XVArHQvgAwUeEnkc/gL5GWmd/7ki9F7EtPnfzR2a4Lha+B3BvkAiV1B1tm
R8i2t7XJx04xC2uiFSEt22Y4pRsKPYQ4ZE6MBWgIyd8faMxpBoT49ym+SPrrN5sQL8NEAPy856Ou
ce6eheLd5jH2OPNprerDGX2smOk1Jhq6RsK9eEUnzHSn4me/SWjy9J0cokKwO1Pu+0tqFqprNp2V
CQeU9Y14JhZBvfGdmJld//6kT60MgSS3ouo4JCZy6vO85rJ2kJYfbrj7Ofcz+0QFqvSPqsliw+2H
F7GubUaYwu5ba61oC6hK9YeQYRz5NXjHGCx8EypyxTlEJyTGLl7gQmV8TQqgnOSXSNubVbKdJvD/
CHzcJJu4P1SagmKMTaEM/iz7LOpotFO0/99959Q8YtaWupk1zJFONLbAKTyyBG1DZ83Fi/GwHYa+
VBCf2CbmpYEo9sNUHpQgeKqU9SQG3lEyqr1rPuE7h0AkuGxKCQwqbQfezChLz4Yh+7H6g8sb1b9b
NOYwrzBonA0XNlIEVd+7u6sfc4HD/hybfB+P6hxNy7j2r4XadcGJyT30iQiMGGVZEA0hCcTq+Wp3
fgspwQ4J4GVB/2p3KMvhoYapTTkq4LrMoS0Vl0jSdyuzXOLi3DdAXWcl6Yd+RVwy7K2O81UnO4Tp
JhkaHJOa+dvTL/QsjSI3GbJmuJhs+AKuuVPC2BFOoS14VbDzaYEF8+phnqBh386ZtPr3Um200Tp4
S7U38aJY8TvW3RdeH+sP73hU9oDh2nnpC51wn09qU8UhSJNfwkkPzTsHICUTOirg6iJAj+jRUxtA
UutmH9j3Ww6s455f179gyFZ26vtxe3VBQepR4GB+2u+1/4fiwnJHGR07rEQ5vQOmkweVbH2iMx8e
0SXE2HCqKMPNYw8ysXIWjLjqFPuJ1dZ6hdibDid/V+X7xLMF7G65M2jUXHKgXFeeQcrOsLnUh3zD
uzz1NmgPwLUx+9ZiH7E/tmRlFIJIoc7SWRonKM23/m+hojThMBTXo7ZHwDm4OvSmHnxta/1GVWjn
pOKgHRVyWRQIBqLlRz6EzCVZb6FWXN3bNUf8nXvJRO3Q8zQ7V0QuQ02SBA+6JQhfmW9m6fYAzFro
2878OtyOL6SkYf5c/Hhyim7ou5jyMlKo76pr1qaeXo0u5TxKzK5x6YdoLpl7Sh4cbBw+HAvrDk5k
oXExWwm74K6chY+lbzVT0obYlaQBMXjZRBMdIWKVDgEoIYnLufKydhExgjUY4jAdmeeJn5Xco6gN
d3lNYSn8pRSQdPlV/2eBmWir8FiDZxPKJj9euXiYlSWxWKdLZgp+Go34fSHWHZll3Tp3PaLr6Cyn
Qh2G/T+QfxAPeLjIK1uAci/Vw2cPMyoE7DYSGjAHNmv4zQAq7trxxGa+1VytINGlC3IxwS47WKv4
aeLZ1BQ3YZ8cqWC2W72sdLk8d9cmaP8r8oHCrqdDJslM++djsI/AdRpQyziIloMiTXXcRarfBSnw
gwJ5qdamsQB4BblvpL5NEvaBoADrjTaBfPMOQOoNa56qbNH6bR7i04PEbFeNH3FnZY0kZ49KI0vF
K+ewkt/Y8BBrfkwVM99w6N6JU4Iqu2iBITQAvNobu29Cxwwt66AEXNz6C7DH/8CKUpgeAZ4pjvx4
il1iovAoblCofZKMxfyKC8UWbwF9yuF/Zjmky+1xwFK6fkQVY062wC85MCgomzgek5On3Xs2IiPN
AQgzEouAciCqouYTB5gacRw07OqMaDK92sDQgWZ1sxMPfiz4ls59gqqCfFuFOmYPB6pEqjI+jRXa
OxjEI19/u1Pm47KBoKL2TofCg2yCguOIIk0CWao3L3x/L/Azn1GMIA2gdXSTJF2A60c15i0Waluq
ZZwhYq3HSm+i388nShb64/CQpl69ZMVqORjQk7dBfWYvmyp6UlZrf6QQ2aedlmRTM6tmfAvJWSfn
h6T/S/0ROObJN0h4tLlMu0A/LDl8lxgetkPo5w87vrw87b3aWZ+Tv2TkC90v2RCHXXF0SzqoNjob
ZREYxirNFTmB9JB5ygFIzADE0rsWhIBb35pR/rTraCupL5IgNTsj717rRgzO1ua6hjDDh7jq+/tN
yPLTmZhz9eOsPAi23iNlDycOO+puiGZOReyc11TmMt5QKYT6dUsn3AHr1ZiUublpJBvjqcpvYDua
tpfsd1kYjlSK2LgxS+bKzqA8n+VSh5hj8IvCTmg0FuuBB2HOItxk3/PF/F8YFPRS9z2eEi5K9A/y
BR28fMkV23R7IRRsk2mK11M6jnIQtSKmQSio4L465J0m0BNVcCBX76toBQPQuW0U577grrRloz/h
Shfz/FUvkZS3rSsqaXOz6Slmxfh3G7USWTI5mKrde1tXjRbsRCo7oxybGnscxeBKHJlKptz9jHfx
WdXwC3qJyY3lgI4FKR8UP+gCL1vkGzuOiFePe+4e79xtpFsPbCayqe8XsouHLayIGXiVgUaf3WlR
dbwzTHOwz6g88snJDIZO7ICUE8i5oMOwarRtHuBClHnUUL9kVZjUODIAWJzaqtbAFKneaPgVf+5M
Ue2cLaVnbDrWEnPEnVcKeTDYwjos0MEk8qf49S+Ek9g4GeSvem7mYY6hc+7wN4T6gtELYa82uhW0
13OHUhftOHnWsx8xkbG8LfTNZ9L56/VtWge3hC2yhZODMkr+47sKkONnLCjKYvOGdE8Es1cuqYhb
QdW+dadWQCDn5jCoQYAbvsZ1zPvjCLqQF+MojNSrAmNoEGv9bxm2T/rqCruu6LXp4C9bjkk+hX3W
uBmZl1lRK+RwtDNXwFMby2YHOpfOHhKkE29arBwTSkRWX7ELoYdgj+qyYN2q6HlamQBAXx5zBY5Z
Mmzk6x2TMqP8Z6RZvqxdeifwfZ1U81JLxnxfYaHKw+eiocLJ6nnJdrKQBbUX5IZozvMuw1IXEw6r
HowQmviAUXEtlNGaZIj597YFAr3e4vVlBWMWGIv1HGDJ9HZF+DW5ZtvhkwU72L07ehEFvcJ7+zZ3
eShrhPNojwYenRhemXsMzc86oY8yXu7XZhZIs2ecp1LGWmCzVTX66A1GJgCo6SVp+i5yFexeUC4T
5ipYwGIFD+tlemKN3B5fU2Dj8nWufF1N56yllXeChqvqZXIHiwfI9aR+RECyZVlQHqEjgzYE4zNS
33rYKhjnAqNKZVbyTnLAJyYntu/MHUBmTO9z8ZKcFRRuXfYLLPww/InmTjKKI0KAtnkAHtq2LMRL
UZGzckM7dqRfvJc7pG47BKfrLyBhL3neabDRiKTDlsut84/5L+0Bv7YLXQrXXEuFbslAxzY1sdCZ
Iin2lkkCk+9Ke0aPnRIjqE4dhubFsMPwX7NJWaJLAgf1SH4LXjhNmFrEYMLCp+aisUhMXWnJ/+m+
4AqH/G3UnzY32IDKA24jY3k7XKNH5tmosMXEn69hbvTag8Kmsq73NVTxlcPz4Mx01c92iNaEY9fb
I1sqorYqqkBcnZQJ6TIgPRHpPmQMi54wziXsA9hNY5SaQTHyZxNcWCMyGHHqT3FSnBRIv6byf539
4vi1m5hHw1bLyVvshFUnKThqA25yjG+DxvIDqGpnPE3yHBuPPxuD4ra2t741wWTnTnEfZbeMTNIa
HXySFVY+c4nyTW7GOoAAEjlELJmmzBZE/pCUzMMSmmIBpFdXhwJw7kS/RtCWiuDcDIVm2wgWHoG4
57KweQzKc1BWRhbWYpxn56d9hNcRRUOyxBXLuiOx8a7AZAGzc2LtAVmspnKhd6KY6SE0qOX9GV6A
zzfduWopAts/lBL+U0zyz4YV+z7deqgZJ3mfoym6GcgvrG9roiIL7uyWM+6iQLmiz5LWNVc2FAIQ
LkrLsA5eTw8F3WJuvLI9TY8cZkXFWTMgzTyhk2hUcskfO7etId+GhHPDezALxyNLrM6Ykg2BHFp4
jGNlSudxcKWVrEMwhx+Au410MWEW/f1iEWcnr8tsrAmoMBEUOxZHJT4l5PeJTCTkXsTa8Cx5p24G
6zF2/kSuksqyggQdt4RmtiKb2bfO0X8nV4N5pklW2XKtv1jrdvSx32ps4Mjy2fTMBXF35Q5xzJfS
mO9rnm9PFSNJ9QNrr0lhkJp+pMBCxuQ/QlHGnn96eaYTjnvmRmewlCAd/erfrQpyKYRoRoWom7TL
wgtf+/nv8Q1aVj/O+xQ9hFb4ck6OagWUGQ+I6EyJTodxTI0A/mCLAH9Pk1sGB2qKsUESp99lCsZ4
kg8tgV2r5F6uCId291eY4dBJirRXATxaEFwpSVBjyy0irjp05L82IYLAZG2k2AQfSAlkCtxpjzMn
Jb9Zb+PlECy4h0k4mzvFyVKhNz8ksHIQqLbw8ck2NBVpK+jSSvZjUItGWiDgp7kylVTgorZZ7lSz
buRX9vSBR/RV47kJcyrQUzzsRF0/98Mh0Qhx1tyXcqrTq/6cBUJhy548j59a/jTYJbbgjvV6jE+U
efehVkNvzC1tWvbblpLFRnm2zVWp8KQM9R0Gor2VueyIJ+m9pGj4Cqva9LzufVBbcaYrVXL3oQ2g
W9smyYRnj8lucc/WMS12xkTVnim/0fBS0e8qJnhcxeI2LsCpFmmSVThArrcNZlTnrQC4Z/kzxUK3
02oyHBaTc0t0h3k2HKPvx5yRHlyRtX44qNRNsKW5bnVl9T/ZTw/giPf4ENxvSKswVbfHXizcxJCC
pHGrk6cxy1BAQ7yqFNHRhSe2Aczp+JPLEsxTFfnPOpJFtyDLRFrhy53Fsk1l0JIhq6NwX95P8kic
WBwomu9KDRRoC5nrs7/DZ9FY7watxBiFziOQ+swPmP26z7U/76GVJl4Y00UrP9KeqVGlGUBIQQzG
uF5ovvyU0UhpofKiSqCGss76Y7gBdQWC7v6uLHYR7BYz0T01/yBrMDQkc33N+4wcfPFpwvL4mOvT
/VgU1SqJjvW0kdEtCSjb79PrBBOUI2F9nrUGQ+N5YuzN4daROBPIBM1l2qVDUOFb+z1YIaZgiKGZ
Sk/ERuBGfJT2OPXx8UZBR7J5dUASPOEd1gM9IvrKg/9hP3QluTwpKGZ4xEFMfLIyQ5aqZaJ9T1/X
LoY8z/ccal943w95l7qI7X9MR4fih38KuVWpgDSVGLY4gmdKYfHq7YWGoLc554F9snLQsySsPll3
dz2Pz3krr4pJb/k2vj2gTG5iVpiVjiGvtif3cVeZqo7WxGpTePdoIggkg7W6MDWNiRvMQVajBAyJ
eLmgI6qHnJqVQTJiNfp7VP+3yOBfyj2HqqpkPHrfa3glosfLir2TCIIpE2BWos+D1DFRoIJ5mHoN
pxhT32SLBm2hk4qeh2ggJkhWU3njJuXNelRG0qilcLjDDt8Roio4Ig5wrwmvbz6krGI1qHxvQF/J
YVHUdo98wV2Q3n28ye7aZsgawyoyaBfGdnvtNMNHy9fvdmEGzoB339LSP8qcyRNSbraK+2z9aoa0
mVoHWdhs4ZXXQ5XeE46TSC+E/GgduXGO72WsohhBlYWzqZs27v1qR/SVZMm6sT5h/WNSYJFhL+h4
r1pSq7qg+1lgUOCB70y7hSer/dAeSVXBrT1NYz5WDAgydqCco8bqNn4v0f26h3SvQYEW/N2ni4xA
kFh7FvoLANSUyeUXkQCg7PXL64UJaVzC2wxo3OhqaXLAzIW+OFPMV6Lzx2qdJ6KbwT0bqzjyWZzM
tu+xxZtqYfrRru2Cqm2yhtxg0zjcokNTZC5fFxRzLublvPwTTro+VsDrOW9MRvr2Im0KjFuBIJD1
AJRbhpF/wnt7B+XsbDW14+5KOefKeYmVRvDUkOUWbTpDNa5y9JVCRVMIihLdyw5sqbPQuQpNcLtr
yIkbRxmeydDGvx+ALwxA9JBpdMr8stJTfKua074X3nj7p3AEvUE1jXQnsejVcoYnluLAu/qrdQUc
3jeVTaF8juea/K3G+CokG3RhD8WcA6eamDfv5t5WQjGM/B5GKBjEJd9GRTypcWUNWnBMs18rKkWb
/Ny/OoTyJoQfXyoug8xcKYbp2uSGFNH+MUCYqKmGghNiKiGuz6RyJUsKEUZ+flA6TbkMUpgRc7Yx
Fid2nYJ4QQPB3nAguaWjwh7X9MGM1wtkSxvRe1K0Es6mJUJxh6gEL3rgR+e/w4dFqxZwQvKH83WF
abRLJgJAPfPHuhGBxzRiqdOAZFpeI3qyr+A2+SOJIRJ2i7fy7J4JTBagfsnFUFodFQZjYyJBZfKo
/DS8wmTe5tPVUmP7FbVNIbGG93qqES9o0e3XCbo+Voo7ZBe32we/YOgWo6vjdGH+fx1zR88tQLBr
82842eNpvN3v7rBrzImQiID0c3A4ZQIWEfgnSNW1xaaqmclYMI4h7Lc7BE3qmEEMvZAoaFNYInbj
bhKZEGGSROqRt637OT4RPsT2FHTMK80G7dgu3gAi27VJbkGQfMHCscXLBVTB0siR7JtKBNjjaHrZ
gYI+/HOtz6EDfzb4rw2TXnfNWmuZqOPxEqS+ulEZe/zMox8cjFsGJFCbjsTXpXbn6Srr6e5dAqjt
0iyGogGZcwtT/sXaJu/eab22oxizdDVftH9qzHmnucFkweFdTegK2/qyJJ9NhxzhlYW790nwIcbp
RgaBhSf771ipPcPZ+3fHFTDUjLjCeGrQYk06ywYA0mutubJb7hqTW3zz5LZaRaNfRqlYxwMk9bmJ
AOVAjFcu1wDkDCJ7mQeiMSGEPnxCLWklc4Pk8qKKEDYokaw+vJ7mcOfEGppVHToUYhF58EnTVbLK
Xu+uYDAShiaMGWhmT8kQCcSq0vI52T5R+1HTe1rVLzx6P0NpExAn0t/sxFq2b5XVUbTnatPCgmEr
FU2HvhmI/yMGyfIBGqTnNBiJANrSx1m5s8aeK09y/sYNQWCCAONUwWIMUbsYunW/GE99f9pDRfIK
EuVwYnzX4mjAYKogrppMcTgLyyYNJ/XIDNJn3PYMrDNgSmSpinETZx/E9qqIrgHiEo6ep+VDG9DE
RKWQli2OfGdGZFkHoO0iqGaBpLetP5sGCctd7whTWHBX4VjTrsuLlzaU3VFBIpBy4KCiKOBkYB28
CAFY1o4spVpMudCro2ikMEgahoLPNxcJv7S8BzTofUvten6oDxGCm2zfvUy/vPXg1wDD+ZdI5dVz
A5nSGreg6Xn7p6610BEnEa5MM5KUNfdJ6O+hDD+W+lSzQ0AFrfwN9TKCr0vHBlfCEBY3KZgQvgVd
jZb98dej90bw2Mj4SV/lO5QmnmMYi2Z5Z+mXxFSzI1m70o7Sm13hoNjjJf3DNhiLSqTqJm0X/jY8
NJKxZRijqVljKbS9Qi4HgxNO9Y6SH+FFBlW7YisOmXTsYqqL2AQp2DxlDvMfmr/4V/XsWSNSlSfd
Gw/Np1sHqJjEl3UqPvWXbGMfxcD56bRG99q/8abHbkfeEolH+/5gwN2pUQlJDG2c1js+jymA2tAq
lSJ8Aax+uF5IaKkqYTC3mnPnIa/gaAClc4REN4t/FWX/9lQI3hNQ6x6ScLnG3P/HbPmfAVv11EZi
XnJD2mkeX+eppi0Fkif4L0IdQH/8cYbU2pcR6Ff7sppHcMkGwi7FBDfSc1DD2PStIW8+wg3nJvRF
art7TU8czCawNHuPVMfDNP0zz6/9XiseN5x8ffptElxhPSTQd3kgYsj3kHhqxelBNAst8E9iQKgz
pMRBeIp+DC7aU26UgDCOZieSOoowKK0lYiYuO/s+cjkzxIQQULjVt62SJ1tku4pcfRQhCc/+P8Y+
Nb1SP40sJxqa4vqmxj+MK8Sw7MGL86e/i1SBV35f/p0rqzlCQSgGvg129QfmygtEUJ9eXeIgStSr
wYnTk1vlWcpxztAfVGQlv7EX/QcNkraYsyvbN513LtUOoPZrsW29ocD6O9rzDoP1zqrZCxrLm/iF
Ud9kNEGev+PUkrYoGUnUOQfTcC/qzt9TFVhw/uGysm9i0Iw3LDv2Fdav2MrdW8IL7N7c58nRYfcv
4zFJjHSHer5vSg5wDGSOEa7SgvfzUqvbqLsukhC2L0EXf4UfFcQmdMrW6iDc7ZR/RiobfFxdiule
r4fx5psaKXZCN5+9SvJtBdOg+R25CuHRl2qt7Gho0NHLuA9kA0uLYWteI4nguxm6rqYrgrpHy5i+
ScYBQiQLLITa9ekhfC6q8+SYWblrou0mueusavr/A+xb1s16m4OY8JGw+gliU/jVHY9PRjfd8VYg
zH4yHt+KwYJauROXFFZlwCvMa3LXChZemY1OP94QfDRiL8bG59NKqnX0KJhqE/+qq6e99t1jRsVT
d3i3UMiPx80Fu4BfVcUpOat8M459nEYyTE7lcEaIc8cE/Zt7hLU5QQgYluKkpF+SbwXRlX6NhuYd
RZ+NpnDLRPu4UfhweN0/CIWx2enQwk8fviUhJryojm3nyPK18/5JZUiDcNTvPjvQhLIDhd56WC6K
MR/H7mDt+68p5bY9uHihdLFE/uAUKUtJjE6KaEZGAaPZEuWUS6me6NmzIrpEdWkh7mkx2a1W69Kb
DDF3zv52RM36P24wpd1eBpNSi7KL4CBjbTG305SKiYOgEd+cFyfRuU97pwbG1Vgo8/QT8V+epyIl
21OW0gcKdlcJZ45+ZexXpHiiQWpzXFbCw8/0y8TVSfw8E+vT9etPNfAkN9NzkuSri6tkRVvcrErS
2wCrZEypwYQJhW9yptYrN0YPRnN+wJhOen8cxN8q6zBEK24Qsfra7rHJ24f9Qfbv5JTdILxIQjfX
jQrtNKPga9GMp891s19Z7Ls33waAONOJtuJjPrr366f9IzpyLoU4+wjq0t1Hvq2KPo4+3SMgM31e
cVDsB7P1LmP+g2RNCSfVCCzP1WBx3dFRUVnC1vqeuG3xkQJ9OYA93xUdwG25REO6vXycZBr8PBHA
KOE9m3hzIKtAIs5C2z+84YpvK+bOaJ7+Q2rWfFpjZMHceGFPG1/Snyg9mObHu+rSEizcfRg4jKXl
NlP9AlCljluuhaQKT3Hn+m6tNWdYIeKxK3GGePjvywz0IU1066I59/D/BttVuU+MEsNufdY5sJ7x
sBzBdaQ1dVlFk9QoH6P7AYlmBAdoJcMa/J1l9TQt+Cy3xBtqvvKRb2iuVFq6HCZvu3v53qQJzkr0
PXsPwjSLxqrnoGMsCbH5yfR6Y2zO3QshqhOe7LsbD8+TARp8gR0KhAFrp7iFFBgs8Tndfsx0WTb0
Am7TkUCMxlQeFBjU36dstPhrzv7aUEJbGG5+OThMMTi/SesBcw+XfjHeKgFHekOIIWNTMTsLk3Gt
IfBO3VBoOwaBfQYrwh4tFHzenY+zYu1XVLsn0Nmk/SiGOhKCvA5SrylchCofV7HCYAXaSPXFD/75
vbgY16/P2BRa3XrmUyoZIWXShQ5BwqRbhQZq5u1yPdyKta8hFRBUM/5lAqe2gJ+SepwnObBt8W3a
Vl0ZyIL56J8HQ+6Qq1X50hm0t+7CWCUtvi0noe3pmpTcL6ME2Y3E85y5RqRKlBYZYkjrN3l86PlO
vCiqQ1zfXJ994MZoQaPVf2opmcZgeVGHxy2QQve3Flt1E4uLkgB/6pC/dF7h+2LFAo/NXs1pwX9n
ZLZMEmSF8CT+wt31dF0jWBSa1+nnoWps4bmmCMddjtKjgJTpupRzO8EwrJ27UoUa7IoHeVHTNsyE
Byqyu1ujVn+5ISI1cneuuvQriqfMCoZpu+rOO3fq5Tt3TZ/tK+hMbBMs31YsYHmujfseM+Wzu8zZ
wN0B03/jzQe+7voABN7W2uaPjQLXfaLq90tIzTBPBtsdJfsyJsC3QdDGkSHJ/UeaPM71r51e7S+F
ofpW7sI9TkjxvY4PrHrbI1r7jb3wx1FTE05XfA8Dfx9MkN0K9IxQVrr8X6YSjTT5XWN+f0kVm18p
gvbhCkZ9L17rMki/rFIGSpAkPk+OBxMfb4/LHl+DObTjH/E0hws+bmNu6pVssqik9X4jUDMPkWBv
RLJyHugHpIj1OJJPZJEs+Uboic98S+s3dPS2SCENcbK5gHvEQMSijko3LrjTNb+8IcEXJMbbeSet
by7puRDydiXTVRGpMwDXiKHqucZjZTAb+4HUlzQeMw74Lc2zLFBdLFQT/9WXfADJZUn3rCznE/AY
R4cLSBgKB9T68pGNrQ5FpN4+Y5noUpvpVt7Ex87MfOk26a+w/R3zalztC5y2jvDDvtD2HAelOQJJ
9Ykn94APZmk2SIrOBacLHbdnx/GEHndQXgAUUoxVhCXvlejxV1Vj96zNvDZLH9ruu0z7reJ50ioS
9dwanTMOYRFkAk5eU48kL/mtsDzfiYK68DcHDZIefqavyIxdD2qSC48cPS8u760pVwj82tUlzLfB
s/E5x+hYx8mxKyYgP0k8jw2DUQt7Eta9fEe7dYVq3cm/LpgwuoH0iLnw1iFKx4e0Lf+iodSXfSAe
dcyEicibN7J3lqratmP8PpqfZIzMvOsxZmbtWV2dGXMYz2dM3G0kI8cg3D1HaPjigzXI/H0isk5k
GVK0cYvYylQQZmqhpbim5s3PpkenAgg7XMrhHY/3MIOZsM8gdyNbR8sqI2dswlUqxdvI0+h+QuCu
Rsw/tQ+f7GUlAHRuJzZbvAxBw2Bux/+hyTOO6CH2x/u0xgLg3HF1sjWGaRcSH43XkDs7TV+5BkBU
pWV/9cViUC/e3rVt9TbaTH+xGtCHSeMqPjIzdSV04agpnppUZOZxFj5SEVK+CaTuF/t9bXDzuSft
wCqfQhtSnmyNSgRJjxE3RnGUJqg9xFQNifgqwPli0SMpf64U69jnEh+c/b/L37pxCm6G43e9UnA8
9JSZ/s9ZJOzR4rx3LuwSmHWzEJ3xL0T2sgsfaR5NCYfHHNXYmUGEX+7SthI2hCMzv0Ck2+/Th33t
qTqmMZBXWTASpvTGPDEUlFdLkgZlFoXWDchbb8VTXrbjTCubKXgz/ZXQr33fQFVqRRlc0Xn6JsUv
dRCX3mFhlQUC1Yby09sZMFeWjsofBoBJIyvbezGOsbocsqBSB6/LINcP1Zjok4KG2NCOsfiTynoa
6n9TWqVv1YMKP+IVwRBkU/xXjy9bSggru9YUEooI73BByIlTASmDKJ6IrIfT9iACpG9GWbuImcPd
dt1INywr6bIWj57UqYfnSQ1ZXXf1L+2O+Vh3E7SKzZWMDjGCnLOsvSN4jX+1twoQe4S3AyTEWH7b
lYomodFk+ruvLzF6KlA1qDw9oPnqz/1e4oilcDlSsGZ4OK9/xbYr3OHY2k33825s2fcdphM/WGOq
PmKcda3WwA0AWuHbuay8MTk67tNp7bO1VGySkaH7FimnZfWuWMImd10yjdtX5sUZoCs6jC/mEbRJ
6q+caeiMB/bYWs8/kz2BbpV/TrPn+2jM/qsYlGhnOqPJXrNq5nsX7a44nBk4yo+ddXBYyGv0Zvr/
NNENFVT7vG9lbQx6TgJvUul3GmcTHBMHBEz8TfudMLxQtz3c9BJX0LQvzJqEClbkTY4WQZ6zMQYN
Hu4zuOMh75j1ODiaV+h2vMgRK/H0uYfw7jTRGh4xjlqoIVO/PgpXK9QxMmI7iciZTHdWfaRNAfaB
ROyO178LX0gGGOHCkeaPf64DizlaaNheS9SUp6OYZjVlCHE8K1u4Wv2Wbi//7kgfGdmNerW9uGTc
1ALfj3uxMaOVC5WDqPf8Y7Yc4CbrdwyPCcfBM/VIU1EBR3ELVrzbvDS5AnvYjDQrLKhG2EjBEOUt
zS84WCHSGENB0YS7O6ntrqKjYblKlMiBG813zpE1B3KMIIgwQFXQMfqr3JHB/rk7M/8cNmTfh0GS
kQmKMoN4ukPqW/XgjK0KO2j1YwHd6MlxI03vUZRD35vGcfU+BellAHfii2mzyU/qD63ckG58D1Zr
VD7m+te4Kz9XGWHkcrAeIXBMqH5DR6KRkkCXmBuBwOGh1YG4XwFpuVJnyqagn+r3EOdUyfJL8BAX
4BbBQAmwBPk8rTLXBe4tX/zgimOdUmAUees9Bdc6QXNzevAUlOq4cT3FAio7+s5Mqb+8/kGHPXIe
ob5cZsDFDU7QgdJf0OOy5GQYdbvkzb1gkZPUiekki1SPcXvpzyCRO8rCVgLi++0vNMX8FB3egUTw
c1ww1bU1LmaKQS0olBmDX3zl/REZvu27r2lrqQxe71NT4PffLRwpOWrvoJN3eSYYLrXMsc8vq/w1
46XcZCFK5jSExaf5Y54eZAthDyAGaKsvNVpDZMgnLVSSz8HTYvgDYSwY+yvftFHLmO64vGUe0JOZ
e6xhp6NsaS+QWv/UdyuoxyuxGoLNwLl2W1AItur2y/3NihixfuQ7TdKGqEyxjN9bod2+cF98YjKx
Z6JaVeIf4qU7ih1ekTFw90PpJccPzEtrMV07XMY7bsEIU3LsVEX7be0X3h9XHS2sjbeoPjKfswSD
vhMLYQXDwH78qq3nX9MQrNoChmETXBiLsRDRDpa6o8kf/l9Ay3Cb4UBizQ1yiq3hsmR5DIoD0y60
05u2C3Z4ceChwi1zzIDJWMTipMwgV+nr98SqCOOhYQdsnI9jwZFLnZZ+5xDDNu/miSFXFZdYoCH7
EHbN5UAlYznxjjkTcKLbYYHMeLVgO6c/Bu5LFrbRpSLiivTQFe796DIT8MoXtXdLzRXrxfLwlJ1u
88/JVytW6M2fhFqQQPW3+ojfyIIhP+RIlq/bgWs5naVehvkfZGCYg2PEyeHF2RFqjCvKlMmbWvw2
5FbFvgmiT5ewt2Xfyvm7e9f/gLHPlaGfcxogHAcJBkzSRAs2lbDkpJf+H/THf9b+Zyq/tWpPJqde
7obSOaz0iuCelNlsfpnlbAblfrzNmbKbYLb8zi6a5QmxcEVToZBrt/+MVZgx0BWni4nlY16pMdXV
OTQTJzPXd62RpmFmr4tvZaTsSdZIhCeiSma5CoZWxDiT85O19n1ZomKt1A89bBfzWAMPnj9CbqSO
eZROjKbQ38k693AVbXbT72Ed56p5OaWffIMTBAuDa/EO7Wpd2Bu8AbC3EyyiTzIs7onGC586WwnL
Vb6qwIVGjRJrd71Op2MnoCm5jqHdxpA6dFMetc9uVpkor0KNUluurtlLiDTId7xI3k2wn8WkwpJ1
ga9n2rRiMIs658vPmIwwUOvyR3K6YUd7uTr67nmCqltqQpSsJ6MzDiJvGbKROeXYpKbBP24ZozZx
4ugLWfVl2s+U0JBGhQlB5J2+aeYKYqmcNMYSS+SBIu3sdK2541twNks3moGTo5+usgc4svM7zgvK
/YD6Y2rocwOASJDQgzOisxqZn2IFayqY9VU2qLesLwS2XyabX091uV5MF9mycFEPbE7CMksykmrj
A6EigwUG+i7qD3eOgbGloQqe9gT7Lbf6FxxEtlZTldcmbQt1qcjSwoqAJ/UGVA9QDosAE61K+EOa
+ww5UKkyVO/aUa7JojdlMroWyNLFCX0fjuk4y01lAlr8/Uxur2gW/eUhFfmjRAx5iUb0bujmLOYh
QlufMBMxu46OWhyoo90Wb8G0sfu73AsUcKB5Yd4MkyvnvLT9U8U2FjQKSvz/jHsywglBeqmME7IJ
l/Hp2dp+ToBcmbJabzQVy7+icyWYdOiDx5c+lxjHIyrlc3VvTlH+LmGGj++ruW7RuAkrsTZR7mIl
zVwqASNb6KX0EQ1exK9kVCYsOQfmiUvCLuDNvhWDiyGOtsEGb4ojqbB1GokUqSjTDgJ12nMmY5hC
93KtWvDFCCUp0iT8fetVGKQ4jc/WBlSQNneqZIMRuKGAm2TxLd6RPQOEYBQUlpib3G9d/Df7eHva
MzoqWFBvVdQuMI4LUyJM2KZ7cDUSmwl7ozxgD+cgV/xBZ8lNg4dxAG8Ny+N1Jvm946WA+gR2AFGR
fAclKB8FG7LNWqyqmFGXPVPANpsEIhRoJMeYwnnZTUjRdNG5y0Z3qVW+eOHi63rSHKQ5Nc11kX3G
3Wunw7ZNW/VErWOArXms4JZNFpuq1qUAdO7rxOaiHOI8+nzjtsBoPXakvfO4kIT6bXeyKi4Vpbt6
bdT2EAX2ZmazcXzWXabUgn+vusUMomaSrZjqhSPPUys1KCrdTfUMUAbqhJ4bP6KdzZmUQxdYaWho
S2F4XlyvdDVpVbmKT/qrJFoP8+2lvLS1gpUkmL0rJ2MIhXUsQc7t8bbeT4VkyksH+3YDWWTUxpW3
ZrJf4yVFzdKCWMOG+QU27K7A2upyxawgUNr8KX1F3eUfaoS7tRWMQNPz2QfK6Wo0JHAtmVYZMOjN
gUNNu+C1+hylpAhlB8ESxFsoUn2wyGeQ1oPbK7k13EZojGtqguWx9HwHMwfuInKd/YHTuohf65/6
+ZCRnQ2VgZm6LDgCIi94733GqlmbD1dKgaJAIrgFQ9brXW/iNiyTWVDB79xZJxnI6z3lP3MltGb1
lk3Nuum/iAVqmXmcJ5zSvIMVvMhFjkwLJ8dLCwUTD4Qig+CmfwBWvUYKRJS3mYe0b+WyRc1Ww9zs
4UcQveaij2MEwCtG5PiT5fl3aqSLUcqvAWhxPUO438vi0DcPEOln7JTdgFxQzA+ftlqp08KMQEsL
aH5vXI7z/LmQ9gRhOirLa9ewUxG+uFYzbh1xJ9c3U7brJtCUyeZ2crP3+cTbE9SP08mj+Z1XJtVp
UxAZ5CQLT73eqyhnQB/ChjCuWkC8Erml8V9eMrE9wEvL6TRqtDHUDYkYuJMWwC2njME0woM62fzg
ThD5MFWVs2Vt89wRiTJZ6olnoyVnKcd/Z7swwtFU1XC5+0Pezn40nI6chnmGLqPSYDDKHsEdv3sH
I1fQ2D3ofV+SkGlPzBtgR91w+YM4Wizju3kVVVF4749Jm4//tx7tmPt+J4+oQIHU1+AKC4VJ32pW
1I0khcPNCwJ9shij+e96dsi50HDiVRUOX9pd+5PC4X8UHsCJYV1yrG7ENSnZGJ7s0h1KlzuSqG5T
NHmuPki88yj8wJrq5JAQNXMkn/z/0AEKAb8RIEi1WiRYCDCcH9YDay4VXKoz04tNoqRk/VORsy1L
cqgwatq2k1KIHlMqtCsx3rFA0hc+R6x5JWQxynocQbu2E8XcmlOgpnnZdgge5JiyLkKTruitrxtB
JUmUaYokLnmP6f2Y3AXDm9sydBGeyW3ihWHUwMVtHqrqYu1RvTBlxTJl2lCl6OzkdPyVBmahiJvF
0Or+LjwO5XKwOS0L3qJiAEcYsCp8Grh6qb79947NXdXAisOICT/H7r7GGqTn2B50DkHo72gfrTV+
ppL2MvI7PaHjKeDzVHxtc9P+B3ay6vJBvsPw3FRsO4H9BP23As7g1YjRnLpco+klJdl7wafQSxap
YlpcPV0Mm/PvI1HbZCUiD61DqpNTZZaoeGObMvZ5Uzg1MhIZFducSRlAD4Ywp0x784f36dY4Yr37
uToJBBNEov8OqpXXZYnXPdyiSNlszki+uSXz3qOZugZvr+M4bmFNpxbFz57IfYSseYGUWUkJ/Llo
x9dqI9Z0GoKELtjL1kasAQKG1b0rQY3D6IxA4a51sxgkI159+b6AGlr0M0c6SgZIszbN7IA7PxuN
D92bbwYaCg4QiHh0lsRqcpAOw7l74mVJdlM4wF5XmNccBffBOHfm9xIoFqPdhxf2LWiYDpl3yEwY
W4HzpqdXnY/4QJ/nrl2kDr264X5v1DzDg1Y0oztroC28oePJBocNFctJXPxCnygTZe0GZbKFYEy7
MPdugUf0Nl0+aWNHzz3d3lfKO5seCBAkls+hzQeoPUIrckSqCmLic0/FPL3YNpXDoS0sfZsXxcFt
E7MNFkALstWSWK0pma3YBXBGCB7nwu7m/U3b4hu690mGvwqjfn7+HN7JET7ECUiE4IhQI1JLBoIx
afisasPs0BOm4rwBq4hlbdEIXRNKhCQWtdvV3lxBOgNjts48b1zNl+k78ZkMuiwXfuN4rjUyhPkb
wWbmIbUhP4CxvIaWawf2TldcEis7ckM5pFGxLtcEWukOvETctAFGiyzo2D+5ECZJHaw456TAe5DH
nIqrepUyQ+Anhm8jT/dn3f/AlJ8auyG2XudYB/XwuHAkoOZiQkZdL6PJFI29OQFJR0E4XblX2O4q
RLfopB7gV/Gyw4os2D3PZG3OdX+EMF7Nxg+x7gkSAGg0rYKY58gJT8LNgXukr0ueCBbCK41FJteQ
onMAHC8mbHm16I8gBw2nyoXAFRr7iCwiCUUGVnMzpbHdAu9eKcDbJ+A5updPUg0SpwVoN5tnBdY/
MSlCPbXKwbpu1mZpfmm93pTw+wUIe32WeI/2H96EeSAipcp4yC2bvFc97V90fg/ogDt6Pv9jL00i
AmkSMXWHnhwS34FfYL0okxYqi4GYuZYxHFDcZVSyJHYyVkOmI8bQSsRmz57jJEfoWGU5Nxy0n32v
WlTPccS/PR9pTa/daYfyojZsjQNxvrKFwwJ40FpXmnRyShskqPq35YIFUUwCB7MKmID2QRo7ltNw
fOXfeCqfcq+ngJY0zy+1bQLnDG+XxtIEsA1l9CEI7o0oAXYq0+krJtOhjBF69bzDcGoNu8kIcWOa
zCsCjiZgj0dEgGMFneSbgzFJKRWKWwlbI13nuzIdQGk2NUZc5IXa+cdaTFdjgv2hulbqg8YMoqdk
8AFCETKONXdlmMlDzah0mPr6Pbr+pks8ihycBK3w0mhM5mtyEnuayPguJ7Wh6cqXjSyiRuJ6lHTy
CUqZEL4ORV6qw6wPv2T+f+3/Scm+fcXZKDD01KVHqkCVgyOE5ejUM49IgyZClJAhvEgsAIV7UjvN
Wr6E6uqfcAfUjEvubZHBtGDXliUnIn2hQjWOfF5taMPfHwf3jtp/GKYLZLYBUos/IAL12DAw1Lqq
i2Dw1Y6qYgpmYTv8sT2dshVlDfQyBk3oL605qYKYD4/YC/XsJvXKtrUW6FDpOrDNNeO58/W2F2Do
72U5rYOsWmwBnmOSCpKzt+V0UPBfXCNYX2ZlwuecPWLPCou3nmoG38SZqrdbg1nUmHk9mUTWmlot
qhiOBO+UPpqBaBEWHxvZz39OrajiIWwVv0FlbSDYyCdduKMnwsbtkeNj82oPLvIFtYu+/n55cQ5o
i1Sy1dG79ASfSi+V3xBh9b6UK2D5B/ECnNy0Y8PTZ93XVLCkMMOZgrgE/6hRsIqC5Cv45vgz/7mi
FsEpY9oyjWibyVy+Aa6jYqeetubWRtQ5HHwft+3KXI8NEV/5tpcZD+YFpcJx/6OBk55WLncbG1R0
7P91zk8URLSH3eZXW3qtADekrJ4jzUKLntpVDGNyI/DbprtN/WwjPgceS++BB8AR9f5S7ByOA/Lm
+B/Jjaez7sxkFVfCZadFX0BDdhZGzXX6uTbgEE3u8FHpPuSRbyPl5/LmQxVKAG8c3eqPpNpUE5Qt
I19CHYbSn4q6QDA3iszJ3UndoYEclbkMZEix26oXkRkd1zTDcMDYu1TaE81HWzQVJW9KeP2DN0Mu
/ouWtwM+P3/PDbyZ5zsMaBRsW/IzD31mF+rBoQInlOmwz2yBooFGgTVpaiO5NWZaVqc/9M8yN47M
QBMHMSAD6RO5WKJ6311jl9bptcieY/Fts7DocTS4suEmAkBOY7OjCnUzvWF5aHpaTjjZRRFHgqMt
N+uSpbXQMyOganpqzXUN1zhaULToumUtBDt+Zo7fjVSgCEz0TRw6xV3mzDAAos/6OXlkpxfSCvGX
wmHFocW8hRu2abWK3ZJp0VqkmnWlZqZ/d2JHluhl6BclG617BsHjivDN8z5O+WUkr/cPCfnU5oB0
e0XM8YapxGSbLsLCa8YEy8/yla52gyv3RTg4RmsJER4P79XkU3YiAg6Sss0JgIdNb9QLcAvUe3W5
CTsceP71aKOhhkZtn5zioYcMqwX0YYfJxxJDW0pXwpFcJlC+g4ZcX18gd+5yP+W2dUN8ZI1qoZ6A
AOGn9TcJKulmNU5PRVqc6lYFnN/xBbn+No/NujNPtz7WtI+ZkTT5NIP5orlK6UBytf8CvooGJMl3
TOrmuKt/OJF+LBm8LfPTsfF1jRVot67QSQyAjHGXOXq9ZJSNtefFWvCMnyCsOXfrM0+AZ2kbPVMH
sJUIQ21rfRo0RhimV/iTGacxHumNIcd05HFxOvnfmhVGZY4lIdy3yqO+Im4A3ibx6HAIMSOfNFro
uHvW98q4YholM9KdRibb/Dr5iUlzy4LYpY2h+1+XB2hvXpJRJc79jNR2RZDaT6mMQUS40aSCtHo7
rnWEh6YszlVfIInJIrf/924Lwa1ysO9o6r/lMHbPS11q6ACgKtHVpNGOIsDV9FvdGf+bYqasSZ14
Px7qqzoC+PCeVM1lriufmTl5Pi4VE4rWc6dFcDrYpAGtHjEpMqSX9v2J6AcwZ4zdwrVCj/dIspd+
cY0Zu1o738AUgl4rpl3lRnIUgkcc0kAD1VVr2faxG4my9ATmuYNupDEhMqR9b/m/hiNc/o3yRieH
N6bnzaC+R+zp+zU5QGalUn47uPdgj+2NyTeYN5e8gwWoliSjwnRaDvmz36Udb2YORDufT7CRai3S
pSZa3ZKcy6g261i8Oydq3gaveJC129+2JZMifooNHmdncvMTVQExxRVV7WCyEeWNk/qSLJbm709+
OSUGE3I/tCTdPDivlFCaIQPtO5PORhB1FN6x3XvbV9ScWhpyrwYnXW8F22o39u06RSfDdROZ2/+j
9yu+fG41VNT+VAQy/dcgB8hpnEt/FsuFrh9yh2B1ovbfTzUcNhvuZHBkcIaTCp2/RBnQYpZGZ5nt
iVlg+XE6xO3wchAGVAmhivixUpTBjK4jACp1URl6tcP50pMMXVCbiJvFA/EFpyUmqBe9ZqKqtZoI
vsD6tlRJDxX1w4QL1A3Czodajs4IZ4SLDOTYoB4J3kwp2TAslaVPrgG2CC4adday9XXQPHoLMMl5
A5rzLzqtyl6VpfAfQ7HvvvEL0gsTVqiCwsmvxLAcEW2MWdhm/jmkkokZbEOAeH3uTbEvQ5sCFrNR
1b/8WN0w+DuIWQVq/w+JA/6RPQyqCaSwUpWxPnXBT6kWJ0yGJAZsLDnBuPpU+T7R5NnmzYRco+p8
2T1D9qj4DdQet/uG/UzqyGYAuFAQjS6OJ2MO3rm+8RKlh97+pQzi+S7k1AFnvzG7Imln5CSD4zMZ
xIFDCLbR3ZCpWmAgAlYxcNKhJzoNYGVSL3XqWy+/Z94S4hHHIZuaTwlDCHUOWH4/L5nvWdEWj9xA
SDJS1dgzyPNFwplVnzF6P0Nph6wb1A5jfqVqfXti6BAfVCUrJlxkpwQ+urFMIDWxozPLtaKNOhdE
yaYq5SPR11D0uH+HGOePm+o/47xl8VjHCiHtcpqCn18hvNhIovXdy3HP1aRhsRDpsU7fr2SXXUZS
Z3cISO4WmXdjbURnD5jz3kQFtjjzFGQdmPMBhab2+wMkkyDhTGIY+2h53ycp0cQkzTkPeDujQvqL
tVbgghAmeqH7i/eVQ/K7ETsKeza0SZ2MyAWNlrDk74B82VqMewe70qBu7BcnPVFmTphbqbuQhhBb
QROkSfEnKxJ+glAA3fo4OfOsBFCpPnIrT9ebo69qiHW7BNrLq7Kxr1/Rw6YxF9OxfALAho2MwFvV
Q13KDA4uzUjMdQR2LU4HemVa40ReW2sonHM7tmoXXZt6VmAC9Nd/KxaqEEXPLh1HTRA8nU9X+9xT
bu9RGJhq4uIo88Wt9V1uQ7+j9G9qZq4SgYfhRJKTBCt0g8hEYwzbyiqORgRyM9QJjk2rOUgIeOcd
1IZ2z5TGPz+xGNHlXdzw631wM05GaTJo7XwGuMOSJx4BSEW1tqXsFf60E2tok/jh6FCP8VD4h11r
yDJPq4J8NqTgh4YgDW/BXgPbfwgxRI+6SvsuiQYSIvameFWLDuEGpu/LTlVT0Adyjzgr/5s82sTh
5yv1us1m2r677BR1HZ6syoEPevbogrS1PNWf33l2PEv8X3mFlpYSAIe9A95+jsXUjl+G1qMvPpZn
T+pk1gbAEZ8LkAMU/IlouMZSDNkpz+nIlfiRIswVQz3WKMb2gKEeITe/CIED6gjIMndjI4Kwx435
LuxdpF52RolKr+HU9Sv+b3n6UWwoaXDIAApeAPzXDXYYuXbJLDZ+JztqWKFG75ijWDzmcW/vAjUP
DT+AYbDXb+gU8MzvsiQvZ2FTKafu7se9FEnewfSvvlNApiYflHX8o2JTubPXtvwgasUv07AN5r4x
VXI7BY6QbBV948uO6wGz5rlphCgcLgnJjP2sma1Pj0PDxu5knKIx3F7cg9TzoNUjl432VI3Mmw4A
P2YxxZp5Tlm13Qrz0lb3Q3QJlmnReiF16/R+7aC704cxCId5DKz/vWxtj+s8xcGb15r5lE4dLgSo
ik7YPJzLs+pa0EfdztwdvFGJkao2haNH96m07ru46zPUjJCrHdQK+wqJC4GdHNRrD5f4vcHeAMvc
++7lWPk/z31G+ObeQhbTISFI6U7Fc3iBKlOi7HID+o9ovd7wG5DkhztpbsVZlahNnKw/oGNqMDjM
xnAbMBduTaUjV52yQCE8eAdZHFcl0V9jQ+6+XB/kgy67Il+u6FozKzjxhLnrat1ZtYjXDBrmZA6e
7Fni0AvY3NYZ69tVguU7iTf6+RS9FjDGrqPJ4jMw/fL2W9vetphHrBVjM32QOmPim1FPtcCe1xgt
t4jSsaIxdj9z0Idsc23dCubUMSqQznaqf9oDaYRr5VCYEMVffgnmPDxPt1MUOMqtKdO4DxGuGuu5
TWKjjp9YD3ja3onijLgkL+oMngiAokLQKGVE8bOKRKEjfLzZT6OBevkKz7+SlGOyI0wTlduzPD6V
2OLMsSxgkejyFYCn0zw4O54QJtgZUAFbaF/lrWeJKdm4BhM87zlmMtZTF7zzuxJez5OLpARovH3a
tLBO8uXqYoFaaSFIcYAtf0bbreYisjqqjxAdhNZWYE/cZYv+IQ==
`protect end_protected

