

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MpZqUX7RHqqBov6r9sp19cCgAmwWMQKz/kilwg6KfQHVNd7thNhiMjNr9jWB5lhCnXS2Dmq96KWe
V2+V1FG8hw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eHZEt9aF2k9bUkzJgCuA+q4yfEhMdqCEDNKyWFDaQseZ/ofqbFQAQc2uVVXTRkEXQs+GrviVm+j7
2wxr0JrS1Xw60RqMKKhLpfqRVe2BmFAKgU2BRL0PnA5WtTOSGCOmSJGfPa08juK1otVgwc2Gzis9
06D0/bVknfjjRpJI8Po=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s0TU3tsqHiK9WgquIx4poaAXQ17I+2l5Vqn12DnbEwMyPpn0YeINJkDaKFxRf41aPK1Wkun6v9Z/
YYZDqYBgVO9Z0NMkbD4LC5C9cZSBdk4ezqdUWACnMS4IR+6qI0nvPM6pNZernzgmYtMGFsG0h7AO
2CLMNIzANr+bYhHkAqpdx/KPtV7Deh8xOAkQeNSD+8rjhU0z6Gg+2FjdPjkTgWwsP8xrTSENuxiw
xPh+QM3dvd2tDQbC1sSMu3CzeLQh9mMzJ/R1uFQDv4VC1TFFFPI7VMPMlrl3y0ondyZNERO3SeHy
Mn6aVbKjlR68QJuFwdsz80LSh3ZTJ+foTk16ug==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIfIqnJL93Nk48nDUNvQ46MGSw+0jZe8QEp6D5vC3ytHCm6yvGspxOPTR0O/6R1kGtbYGX5AVD6b
KvoAJRDP7Wr2E6PTOWfFxWtEHCKiApDz7UksHM1gqF0d7SCMfsYR0KKn9LnLJiQxmEJD5y64ve5y
9s0qEeMi9k4HxMVPc9k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XH+fS8ngHwfDFxF50DT7MdOHeXbY/uKmg7Eva1j7eQ+2X+a34Rn17d34wKLf1Z56AIT4ksXzo17E
WT5KT9rKAQNao71yUm+YQAunOwqKEPRyxOz3bb+3Zvx3y9p+F7xTeZFLan3KtqwByX5rGkNJtGjN
oI8H+T5FEpTIirQ9oxghooMSVVhKX8RsayssyrgajR3SSX0Q0ggoCOy3XtjsFKfrcDNlt7iEsMAt
+8vV+volJUxGGSYbt9ATDx7fk+pYKVnFR1jV5fEpxyqiZQoGjkjsnbN29jqgiZBfhyEe2uAb7sF2
RnfrEGY96pFoR0k3gse3XEc9radVftI75N7ROg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5808)
`protect data_block
9uumo2yHNCHpsaHIkOIV0iZ8o079rfH3hyuylZcFvf+jgK/R+7SThESj26Nh8KDiUinA0jFf2xSm
5bb5sjffikBu78Jc83oMxBqK6LDjhKOoUu/7Sa2SVB7edh6wj5Hk8KTyeckXCJlZzPvdIV6cBnUV
K1NIxDgWW0fZpclVY0N6GKI3L5oHgg46LJljps+osn97XdvU4LotCf2c2FBlEoNmvqGGKspeWPof
d2nKDfswSV85rR5J7RZVArIc+AyLjDp7FDLfcUfgn/WpmgsQb/JQJn1ZuBw4r39xQ5i8Zjn47vg4
3FZca4g9WdD1YKQ0RBWIDcCVIFm4cSVRpDdHKokG3HTkPcfm0SNgwvHD64y9XtyIBudpDXiHMEts
8zXUMk5m4WOy+Ca2YFd4oW4nk1rJ2EAbfl6MsARk5egrvO4Mg2YL4rVP6Urltmc7FKZh7SKPwsyS
uXSnoR4Lz3KqFjlCbmElV4SKgn0UxNStX/hZVRhkGD8av9LQCwenINBO0TSn57mi4HJ+tyQETt9M
DOlbjI8ZbHLzQsDQoY4+Ry+AnbGYI7TV64n+NfObaDoVjSuEuKsxMOctXx+yUXjxQZgiTX1uPSo0
TL6WFf/6sVksQv9EyF4qE153p6pkeKMoI9Xw0NFtZ2da+KAFIA7dEckvTpsa7zdMl2U4jnBYiGFO
LW8PImkbni2YJ71rSTuT3u8grYdgy9pr0XsmuBq4kPdBPx2uOOy544A9fbGdYMKciv7THzgCophN
9lQLjcC7Dm4n7p3xRFAHhof6vZqTOaX2mpBy/7fmO514Sts4Cnm0djYkuV8hrVWRjKb+3YkJAHpj
r4bnE/5tgK/cZ8jqGk+hX7C/CuLS5UPbiVKOxZJGzKJsp+Kllz0eARJ0LuOYnjZoxGl7OyTZnokV
LyPgh0zUnHqfU5xCWMRH2X3MIHySEjMFp54+LOZVkMsJMrwKAjjB45yehfsdayt9SctrzIo3rF1D
Gx62NU0H8s8Xm5v/yV9dvpKqu/UiN3P2/drkgYf+mRTINRG04q5TvjOzB7QM/B4zXGeh1UsxMEOf
L+dXUnzejAhAb5U/TVpoD8uNZC8NMUaUIVN/BBffSh+9taYQZY2qrDgrnjNM1rYto/iUT1OfqmWn
D4TxIidsWmi+M0hMTbKJlHluyBrEF9lqzNJR0LDDDHMcEfh4+VCPLGgZbhN3rYpwEMvAHUgJCmkd
LmH3wbXpHGHVhR33Gdmh7GHCzkde/B5ZgPYlgGcuHEyb35TENfufa8iIIZkkjENLhekvcfixY6cZ
Y+5oRMSnICN2+jxdKudhTo8WEIy5TnYlbHBWsXwd0n/F/Or5iufTbxvEKvKhnL6BpLCVXSbJ8Dje
EJEcMCIpweAb9sdHdRAkw3QtfFysoQngBpVteX3sw7HgXBqtnDUGUkMHRBKc8999hgOwdc9ViFtO
o2Py6/oG4UMrchjFF2T01F5EM1Jh7ucAChKJwDart1LHjVdBk30gjz7zu2iiThwiQVainRk3W8wF
sSaEmo1heql5HuWxo14RYxBlubu0jYPxG+3RyJcfKJ1LX/8d0e101+is+haerYX7zuR8qwDE9bl1
1y6MYcP9AZJX0ghQ3CQYa/4uNcF4SWw1GvQicd1dPW7trRVXY8NuVcaWX8ZnfumV12MHmATqO4/I
r3ERmail2UVRmwK3jvGLcNO01F8LPsAl5rhKri07A3iDNVdcFqk56/hlitU1yKLhSX+tiI4wD7jv
ueP9ahWcpPW4P/naRZCQQx152WdPZuu4+odHc567BNebmx2QkXrqlMxpdYlRsCtSWYz0uBwP1e4K
lDXFDygM9iAbLCb2OPvIO16BqrTQGEtxIbRgHolcGs+I+enzJkFU2vabZc7OZLUXrLboLCUbPDpX
GXDxLybQ3pZ8SNjRoZiPKzpKtZWjaDN5y4uu6BXocIxv/H0gpWYwwcAmaNp3zcxr2/sMSGJLV6lw
bLbhRzygbBsy5icFQiLuQsOEK6bil30gYT3Yw7HDMrByuRFzpKWPLoREI1qxuB7qjv+apIdI5Jrs
WlO5ebiMruifZ30cXcarYu+3UX2Fjh58RWhGyIiknPvHwAJ5/sBBqPzPCmUEeuPEMqH3dq83lK+w
VhGHjbR0/TCXCGdirf/GRBvCdg/G1d26fjIEcFgK6aPXBn2OlnWtl++m+nBH7UEc3cRcMzADfFr1
koGpQAmu7BtFzAlc5tNWnXv+bShegvPnju34x9T59Exx4fe59hCyHMyj9pldRkMGPZtZQgf6CKT/
c87+rxky2Zdgma+OGOP5Tc/8mJDkLD9whwuHez84hLIh38CRqxbUqcNPlmUVfC49K0smfaI/MrHe
hJ2BshxInj6AFPf3fTC37c/FdD10Q/46h5at7/slN/464CaK0uoagjG1a2MipCqOasL4GI7GYZbL
DBzequ/Bx1oJFMA75h00e/6aYat5CWFPPydee7zp2EFSPNH/YvQif7zEZ+zqdlMeyZd55MjzhrjG
lR4oae/PlAtIFhqwPLQFxtADMKAh19rj0G4G1ez7dvj1cLvkqHLgvvxSo6C065iUkJfFLHKPEaiH
hBxIb/Hdm09WKF3jvHFXIaLFaMeF0219iwshtw4R/xxwXo0zjDlTVgi3DP325/MwtwZO/T2zxoZR
NR4Gn+FUpLVNJnEcxHwK6GeXIhamupmZPdZw7Y7PfTUutKYKzPwpTJWf1OqnPyLj//YXJhR83fPp
xo0XS0zLFH4qSAPrpNUZsF92zVJoDS3TVud9MSrOXGhdMTRzbcpSV5gkkvIBxGH7pOsnZ8R5gFx/
3yNqFeMJO4t92wRTR9tCZ4g7zHq9ii4IWgL7eFpcdjhZffneSjNFAeJAVrA3qc9gzjOStp483M2r
5iGvN/hN/wymzXMRC9+nKieNmg0SzdaPiJueAn8v9pb40FfWYMT7o1bdSyzAwjY04aIhJE203ZA7
huVeYjXmD4OdcUAjFr7s9s939nU3fx3Onxlb9Be+46rdrn6zo8RxaOE3fa7uHdKXU4CcBerRh3fD
JYKp+wHDft5OOLhcYWFlz6WepysKquD/+kqFd34LdwioP/nmS4v03StXBjP26RjFcbaLiYEysMOw
wV9qAfb/hrM0cal+AuGRZnb6NnlWkNeb01eKxoRgA/KItnZDh7Ps1QzO1oVI7QISrZx3GOv3LQUC
39P3I91121SiEQi3XMEGaJ2nXGY+fUrG9S/7K1UfHNlwy3RDmx8nHW/hISJLQ5QxqHQVC+wEZtuF
CZFVAeh26qyCJS8NsCDlL3E+5tmaJ0OOM4vxAJOteomAuEiyCPDKAMTG7ROARy3AVwxx0UjupdEJ
E6JejQjXESsGZ6lRmQr60xBq/MeJ9zgCyuaUjhp9MkYILeNgsJQOp6OkF617zu2WMjNahzHaLfPw
nZmX3kE0u7NK5ACrG4MKB0Blrc9EUhC2fniCkBu7aSUgLJ5kURkiV3LPyPKGvkwfMXU12/q8tJXI
zwM44Y+aIKmrSuZs57Z4n78ofeC8MK+KDIxrtrb2AEJNO3868eGAWDTNpieux1vYQi6TeowCV6IO
pUGi4QFVg9H1K6GuImleq5llaWedXUFbNZ8pQoGI1iHvUrv+f+joJcm6oa6dyvChpBGklv0E1nb4
hzHh0AkttOxPVTxkB01fI2p2AF0FOeY6oZD5HkhYmtJccNrEl3vRhorDQFJ6rnrzMjBImbf2K5DB
YkVboBaC5kqAAt5TwX/XSrweY+rY65NPmoDWaF+nyGVJ6gN9KhW7awrJN9/sN2f/b15fjq/934T0
hN1lxA+7+3pMdNJa+89lSpg9cnCqzj+j+7c3kGN70qzLRex+akrHqbZfoMxp9R0UkURtqrvq5lRW
KXKWTwtsy9UCqLV+0rsvruG8axHE5n8NlOkr9oHJjBFSA0Qlm7jSdq9mg7tzrDKpWPthpJq7sV96
zMECU/QuuqkFtYH8ISIIvyJqr9H7HWNFGgSx7T5jNwgyGH7RmpUi7rlU8sqWKNl0qJeaLf403chO
qAwElHGtOJvEfIYME1Xsq7KDAE1htu4tTuuU18whfGjAeL7CDSjzcrZ4fxhU+RuOZDYBGAtHIDSe
un/mQB/R3AelsRT3rZ9AAUGJN2Bucfv70aZCrnSQYE2qZ7nCvwMbBdluDzVF4FFLm9ljqTVaLuhe
fB05jkxc3roSR3O9OtP8JcF7CIJF/UAX7QDI7lpHL+b69BAF2ta4emuxMOyWwZY4mxeMwix+BlBO
/QfWMGxGeDDjAKg45O5JxTynVydnQpdoZ74uhIupyH2g+mo6kUFIkquLftTr2hx0bLIFJT4ffXkh
1Hv3h79AHRFroXv/sjPK5zRxpQCkyHv3LH6iJNQY2+Kk2rQGJnTA19OUqOrhnIXvyl+nVeGhxrTz
yUQgOV3G4/5XeJwrjbV9WUi2Zd6QKcPAteA4KBC3DUlSluBKfrtzvoYkqc4ipnL9GExzImRJ6PNk
BPCC0kGQYXbd3ddxCYBatJY1QpHUWTRYHBmDrqIkT/Jxmq/lZg7/JzVSfNH5fsVJmJeesEk/SAgP
KXwjXnRYx3u7pNln+47HSgL67kWQLtaIJ7eEtehORzvotQ5HGCKJpbCcxo4Q41wULOul424dPx2t
r2XdDdHBOWty7LGNrm3QNWbbdWSg0atyt5QcpqYR/2UknK6fyEbr6kTlI+LXHR7he+CKjC6TO5m9
MIvd7R57xD379P7zvt4skgauh5YI8mBCraPZsDu3qGvr9a2bXuD+yQIwF5YidSonSJRLpqnbv5lU
sMTlkDbCfKp6dL4NLKgtlThW1oZOXO00eK+jFlynNEK8GD8wTMYqeMYPSJjQ5LQfjHP6Bw9mS/xb
v4L60dw8OvIrB+psPTLOT0RmgLGDWrRItuQD6Ndl1O217vuaK8yMjBHVTHIMHxoy0/plcmReLBxH
UbKEd0YPbouLBNRgMDwNECArh22KrW6mnilutI2rxE4buAyTFlWakRa7ulqUOCauuT0sTgAWHys7
nN2jUqTn/t/Ip+Jx8PEnL+rsLadQlQgyLO4b7ibexGzn6V2t8ghGKpsXQOQjAK1q12JKg6m+9coQ
GFDFO5uB24oMeDM01ZtohrKCD8Fpxzi9eXCt9GpYPJ10tzYK2p8/UbE/alBj8bwOmJ3q0BCGHBUQ
KfJyScBT+XUcDX0M5qutKyDD8841xd4Qsv8dL5Y/aN974AYL8zB4/YQZH5e2IB5K8eCK4zRaTGi9
xmTm6cWHO9nyiq/fW0ztJC1N2CEw/LAXy4hZpO/SRjDXLh7fm8UvzBG3ho6bal76/m0uOTZ4LR8F
C3hJ6+1v1m90jnrMby/szVUjDeHoUX94KAg6ZQaGZfi8OIW5zvvHp/X85wYreP2Wfy81qW+DSSAV
r6kxgdxr3t10mRs2p3z3V6PhHG3KEcq72J8+hW5Hgofm509DYGtfB0Zf5Jr4nGnaM2Z0/1wdBmY3
xZLwB9nl8Ov7erZEujj7BuSILyvcnCteCpTx42fZ/TnMdpSGw/DiN1janQID/ntAFjV/NxnXbfDo
vSnFtgdtnBjQYstGOl/IUslLuDpL48XWgJKAu1umcKPmz8ddcUpa4Ot1C//C4nojs8VC5VsTb/Jq
ztwBCIk0WwFCMZbaaQe1AVeev4SM1knKRPXUjjgmEsYbZEgLizZAhNCxpR+CukHYjGgVJZ7YCv0f
HiljWscnpaBWF6aCKJbPpWWPFoo3Kq8X22o5cTVT1H7keXnfgORvYeusR7/jzrFCYj+i9a/cys4A
wkoLgudIxEKDS2xGzJtRkgtP7/miPbq0gXNm4+OoetIpdmJLfoNwj71LZQRbunux0lSDtrFjxf/e
KYrHWptZ+gG62MOrZ2zA9k1IoLctHP8r/KntBVndDlNBkdXB3Om4/d3FoFPrzo9FX0U6PZA5vqT+
OPWkIWjUU0EbRr8bLPB4+LMO3xscfN62vIb3loRnjnP10woXOXfWlfeNVI1bq7RwUQsQkahZQSeq
zgB0YmpMbQ0ASDc83lWGp1Vrvfn/Y/yOk5fue+uC1WPXGajiBM6gAJf2cVc5qe3WG+Fogd08Rh5/
WTPwQVOM2Zo405G6NXi/YXechwt9nU58yubCM+nN+M631hyhAr9fd0ttfS2PIuwfSR9iBkxbt8QX
hnnkBx0BSbQMmh63zXWESVIL7malh92sBfqzeDXNfbOPrmwvXFLTkpH89W/ZXcmxhX4ynr4+NPXK
GGB1AyR9O9dwJwj2YeRBGplokfLXXM6QUHESPyDJqwfUP+c1b+S6vq7egUnBIfyVso+TAU6bWKPK
k8GHSgxv/FzuehuXiuk0ncPaxxVb3V6N8Kcvth6DEmum2wq3TqGmOlOyRJ0Am27+d5ZFjTEj/iiC
vLIVMKpvLXz7zH77MwS8iEASbaj7q9p5Sq+yAlaWeVvyzpbyxYw1rX/jF/fGFd8UAjgTaXxYPK50
1w3xYO0rYJxi/XXrnFmy6e/hpVeO+DcNVEla+m3DeEFvy6PWm9GIMVmz/qmmGsCsOMpC6P2tajjo
FVuvkhKau5JDEIZHrfyjnY1r2Q3T8v5LF4Q8INaPlVc/gtnl9IQ68nopx0p/XQDO2nbdVEVJ6c5i
1HGR453boAjCuas2JmmH8qSM8Ie+GHSBgBfaD4NbQba3scv+G8ln6jRKJTCdgchQltggeXX8Igz5
+hLvizcwb/L5NjSJ5PFeajNzcEfhZKPYW1Zpa21qdMvtTv9ycwfBf8wlXvIFffEJ28zGhkJUAWFD
gQKIwY8sFV2JFTGhEOOnSjP9jHBizb6Cd+CMhFkWoaq01L0Gh44L8Y+WObCG7R7gRf7yDQCn46cg
DocvEn1AYJig/8EArSIyRxaJ27ZYf7muD2hl40HMM1+oGus6qr/xy7B/tGozk5HFhjVtziXw/bbn
r3WK7Emgf2cveRuLVCB5gk3BsuHdcgBd3H3rZ0OF9GwZ5QWUqLu2szXz7XMlwSwdMPD4fBEZkEBe
CgoaoNqUGJCUTkEFsfGnE9MMipLauBVDY5njUxRefNT4F7nwNS0RaweijvlZNi1bNktPPSYRV9xY
9iVc4KvqAnSR+1TSU5izPlM6LFPbghBEhw6RaPChiG7K7KkEglCf56P4RGknlcxnRyNAfJL6FPMs
5MM3gYJHhN5RMeGZVN7EKSZI5hwGRO1XH7nyo+oZ1GcghsUgHlttYRQfwfx09gDDBeLlcLYyY8A0
aLhlwjjVMmdE0OkRYzxSFyjQEThP22Gxq/jaCq0rBz/DPrySp+WT7/BF7fuAKvtNZ0+Jn+Zy4NYS
1FvjrRzUfEPT8lqBQs+Kw5Aftd8jyXhMFbKk7+j5m01ewlakG9lHByqb0LW8xIVv07OiVmQ40exH
NLvaCc/deMWZs4NKTc5VS0FKQ8BivHhekIsChxMjnPeQ+OAVYXcbYG9M5d3l1CbERRkpwL5502Ds
UA+hSgQF7V4eDxlmVwi2oiQjAtoKBArMcyT1hOtqJXpccOuqsB6P5O5JLuw9H0AXCwGTFjgiIU/b
+nCSC2LWHTwPZp5N9iEHmv9DYS0v3fEOvatt8MUqk7cbmx/2XXhu9SY5hCcBPP1LSh4Bb7mGc8cy
ZATgxKIinJSLuxT8ibE3+BbcyWjn6P/XsW47cZAHBH4Gz+EeWmYxmOnXTws0yC2jg/RYu9ake2rM
crcFKVIhPmYMO2I7g2AdiqAVwpjXESjy9feLCOFNjdI/yGv/XQBkQRL/zrgpXYBf+zQf
`protect end_protected

