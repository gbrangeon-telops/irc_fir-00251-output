

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VHfaMJ2jDU0R2eAkOntfC5B4/6MobpZ0NSnc7trviKzQU5KHakm896MNUQ/U/XUDUOQl1Ix9hEug
uFcdFGHOlA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jZ28dq+cqatvP/oWT0j+kbhevax+rcvgcOVET6FHORIxsClPAe5EiSXk6mDgtoieHOJgnr3iO4zI
pViSw9QXhHwC7nkjQzCL5GNnIAYREubhi50JKwxrsTofbyKzT/U5b+jDP0girnK+nPIjwrQv3vvD
PHropUlOeQU1eg5rEJo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wyTaR+5BBK3PMm+GuCvq0Bco7y5f/oiFqNMyoEJ+yA7qA21Rc24sV0Xv3v9W4doHSIdeeP0oUNh7
9I5Dbu7bsdY24p4a6rVQlpW5VOJjg7abnoTszev3jaBtBOpAM+FQDIkOj6hl9ZK+eUTOGH08ap1P
3rtu9S06fVXB15p5GUL4qJ+pbX9as7bXZJVw8JMDVFn1WsdJ/zMn5PNvL5qC5jZb/F7Sf9m7DkwY
x8I3vpZz7RsD6/RmMhT4lv1FkcH4MpJegB1J0hL5KoGG72FOKCqONCLsZdmnqz5BmJzgYmphlYZC
jJckdSX4yOLEg+jbosSObzMclIjrm9gORAOhKg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qekQcsRlt2+SE3/eW9XQwKmx/wWWvcG3c3jSLvuGiy4GIetXM6PaXqKAuGTMI8b+mux4A6dEdodI
mIX5ojnf5ZA1jyISA9q0jKtn/LDbiV/JtKzm0pK23fPqh9/IUaTz+oirXN82WQzZFKQ5TKpwrFn6
ZmImSJcOKVgUcM/iG2U=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tlEZl/v6lEdJp5aVMLYyANJmLh8DNrpNnDhyEkIUHbeTfiozIDqQ3eefGpJHd1yUjxDr+M7d69UI
c7u5loKJo9CP6qAEjMhB9NE50dWkO/cRVvdlBQSlpGD8Asrd28oTNAHTTge+6t1TRCmYfvMKOt+b
zBqmGPTyIDG3LI8DiLXNfUjWjl16n5IRikeD/e8FsFJjAF/a0Kjal/N8CzCmRiQPdsZhdMiruSdi
vpIRkNPRNpCK4J6asTfuTemt2JkEkG10IvEYhZ/qTCco9PECc5G9y0loOf9owc6R54o3iALi9D4Q
T0iTW1tROVF1jLbRTIe753z7r02QD4PyC+02yQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24176)
`protect data_block
QWKolhBabcc7fFcq3o6DUmwOMSCvFYC9A7uSOELR/1vmsCX7K8Wv4EImo0bDK0WzyR1BRuAsPx1g
jqlgOSYF5N51itAhBYz8GhR7kpo+iYg/vDmJTBs3P2yRtpnkXFXP37EA8egzeuj53uzrbSj2+GNs
YJS4xvehMuhfg1C5CTT7xhFoDZL3Eghnf4xNB4OsViZsqorGda9jjGLeNFKCK5VNKIiYQkQwpvdM
Jo3WEM0SGgZaBj+fl7R+C3NhXeqL9Nxjkt1XtdBLBHE8e0r90fcqqyZxwv5JRRnw1s96aCOQH7cK
XVdAPHaOLpD6v+/2PPzx0OHlHA8i9SPz42GbCr8q70MOp4wF7OUyYlWFNZ0iKCA5s5qv1l97GIqE
4uaneWK9ht7dH8Rv03yE+2nHTF5Ox5wVcUQ2B/Z02xmsWM+I4cLFIOCUa5V0mAnSH+5WYrnOym+b
+Vx1mm7IeRk0ZqMZ5H+lHu1QfdYOAYaFROvg9zrl9Z5jpYNrlLtlZ9m+1dTwFp7IK+wruTlh85oK
jlQvRYYwwdyIP+XPZMU/2wzhoI6M6ZJs2A9gL43jplnOduIjNli9R+pg6VNsaq/QkwreOQAIr+hB
o/6v63TsQ98IRO+OzrB4P6D8y8PD74waOCueEg3nKfEH467LS1fyrFINOPHPPc6dgOTOp32ZIvOh
pr0Ysy5aBVEv+D0No21jkXvotkARDxpCRHH1mCK5g8rPPhkgs61HUqZ3mi0WRuLtOl2O3fwqYpYs
cghDXE2TL8Ouwlab4jkM6FYtD2wMgE88GZ8h/3v04MwxpDGdKvrd65AmaUlaJ1whbX4pAmaEuyfv
4KsSh9/euDEBvK6GUrfMjBPs4T1mDENqCcQcacBE5j0HvqgwPxONv7vjLiwxuaOQjOroVKOTeUki
uwijfu3s2/k2IijHtx/jkD83qfStS0CfH+PBgDAKqe0dfnV7+xS14ix3rvlRcrU6f1MM7FK/SvOs
KmfcMgh9xWwOfy6C9eqsX/iCJbl8YEcqKrEqXRPAnA24pUUK4yQeweB3xq9QALrPALVM3cPgMKCj
Uy9hh97s1w8ryWz4iLuH1Nyh/qRcwcHYiPIchuxQ9yRrLXbOh4/LuoxT6rCNYdNU9KxPYXHC+arK
eVOwLVVBO4d11nGt4EU7d8edqTvHaHAHg9oGOCqYHZlVdHroZk3nNekQJquEYsODFkN+MzChXEuG
QCRyk8DbcE4FOg9n1NqYoSnbyRnc7bHkYbv9WkDDbYinWFc2T/NQ68rg2MWxVVTHt7oay24sjE5X
w71UAZ4pDRARVBWkMD05Zvr4ztGp4GVX7aaa0s1Oiyc0bBvxkF21UHmqlpKUOXgQ9dpkTQMIF1f+
EgIqEL52LV/psDKtdfrlX6tAAJakIQ3M0Mcr1oj620lwC385PpVkALjGo2z2kFymjjsMCy/IXsVa
ANJJHE/grm/ko9Pr4N9r8zvciEPnp26WcF5mUHmL4wZZyjoJ96Gf2c8Vn/O6Hrxu/RRDRKTVINcF
MQxbUKuuldhToqrrdg9ik12g/RNZDW20vknpTjQHDasornAv4pO7SZnTdGjbKmC4Mjo8CPhPrnRT
O2bTzlrFcPhMxu9uJKs2zL+MXBQ8I+YKsD1NXKSUBM/ODaIqUIN5aSNN2NyRPaZkWpeRhhaHsj4z
hxcG6r0QtopKfqfpms5MN0UbkkdxbQlXMHJgfbYVXNOuX1WtwWWg7ohvNPyxZe40mGlSg8QBqxbJ
CEDMbnBuE7eiFf9nwIHR50ehksPNXAztF2QUl0A4aRkAD7CdjN0xbSJehkmL5UmmOf9BG+oobvLm
IxHNSFp/lt/BbiepOQCSzqLsU7w1/stJ0B0/4pKyIcANecJyQ4njReVg5S+LnQZTxa0fkdZxb1cd
KXgELq48LOkuTvJoRGQPFR1iSQtcBIP35Ia3HhZLJEDXi6tcxXG+TZFq9KnUW2w5zsu54sRtSd9h
mmRYQ6lSxEx3WWjJNSnGNzEZlOCjwjEXJmvKAwuZan7zeqi1CsV6HYW7h5cD9hOl97nPgtJUIjaV
yWPwLubEAd7iCD0+u9W/hTbY84QeGKwGUaZRgtlX8wFWFd5wTjK6SzpY8zPDruTDEIHBAHU8TrxS
0q6j2GOg5lIZmtUHirtMODtu+mbb/mzQT1EIkkdtsziHMU9PoUHV2xLa0zMhs8FWnei6pLhKjpIs
fnRQGFGjUvoxSwReAFPARQZ6QhqBOTgrYV4U5rObakG5LwdzH8gI1VyErRsiJXGeNK7MsWzewLzZ
EBLkyEyS74M0WI2kywRsLMe9TW5gZk5nR2BNl8V/PgRn3mp7zDGG44fz1/fBp2VHI/qdA6UFiQM9
qHbUWoenGBS3ax7GVonrM1BPIfuBZ9KA37+nB0c7fcu6pulqHmMD7I6ia9Eh1r1T+QZbKWLSqsE/
rtr05p9/WTWXEJQ7zgQRcJ2WZOBvGnl3k4IAbGfvWx89ydC33yz80s3ujiZEaiVvoESSg4+o7q3m
pNMyyWxcNm2KhJL41c475nDZqVRshhKNgJXrCwbLNL2hWw1ei9XpyDi+xXiLdmYh9dJMZGTH+fZW
NgixCw1phz/nVuml0+tP32MzqRWLGjQicL80d3FIjxVD1GmAgstKI9AseK48xiE7BxnGF7ozQGOW
mDPY7nwnzqsVeTjc06KKR0xqq3r5YUc/cSpIIs3bK32gV3JCuN8S3ibyeFdhhshC3ebnXKZCsLKA
wn7/rCYtJBlkBIiptlRKwFrvpt1Y+7eZ3uuw1pQyPCGAWqVG/9kEcDHLxE9srW+lbdhhvsVeV6xd
wx4UXVntagFUsieDK3JTyJ3xrBKfRUgkzfKsNo1Em3CO6e86VDhbjFb1swAqt7aGw1E7HDhzb1/X
PQT5aeQecwkrKZFxnnn+Kf7LJV5XKe7GVFUDdt+IAL00zuk7BcirwiTxX8/2OyoGuv/fq3IDaIHl
YFWTOAk7FxhZ5p+DGBoXPIIevO4LQ8dUXdCfizak3oQY3t7xjZpcZc6nBxkSuelha8U+vfWDmnnb
4qfpvpk8UVkpXdDE8SmdF3khs+Yfjl4luXiQwWCbE72GtMqkS07/04f+AaUVmfBym3LKePjCVbm1
cd/4tcCLDM4XpWkbTojtc/+4yheFFTC/bhTe3SN2NS8AQqGn3AACSaYhE7yD9rYMbCnNWPss6GR7
yCCMY3mqdfx/k21+mxo//xy4IaMIzKpNSOwjuqVmbHrZ46HC1EOIbtL+n9rvC580Zfh0rLsyQa5a
JhCzKrMKjnMA+6FFODZDBR53HBdfyCsjjAAE8c8+7mGlWv17YAq79u9E4TUQHpLbD1MkneaYOHfk
n7rV+bBlEcTBsQWqadcZbdMSN4Tzfw6c8ci3YbHeggAhMQqld9b3+UmYgXF7QIxe1cjpiQpJT7In
19wqU2kCsaqEErt/uBZ9BB+RJdsZBiLD3CGUj/m+dIqn6V3NqqNePRV2QAb6T4AgbkvSU7nLqh74
azo3h7w62y/GzVxIa/7UwSY+idiB/HQT1nk4U13zK2tZ9nj3ivw8ZuFWg97tgN0XOaeU2v7TIS3r
nDmNVpTYa6Wq44a8ESEQWO4+F5fOPrDkr7oLpQbXisQx43FMCf0n7oZ779PnqloksMbd2LqLJhTg
2ad792wMiNczNeaE0aqDv0oIZL/yb4hF2PZ1fMjat/Pt9Hqp5EE1vCc2jOBzIr/eRLXJsemksGts
9dno61uxDignMgO8mh4hmXLiGFb71xpiVDp7xLmY6h3hqUspEiTNRReJS1ClCffjMvte8Q7cMyOE
bnf7Zuk0885XvTJeWf45+9r3MbaGRGnKBRM6zu3SEucHYpeJBAS8CUSWwPxh47tWhOpBnicvfuYD
V6ONKPuJSIF9YG9dudnqOm4bD6qGA4oq7Wr7bPBXTtvawqfu/wBQajcDQnrOcxCZoRAMFvhovIpW
0tFiTTKVbxayA9qARUuTKvLsiQlIjeU89dlLW5UZsZAlBu7dLbk+gP1rf4IzObLojAPjquqd99fv
yEVNedWZa66HWXWCyQP8tDdLoYvtZDq/1HRxab0Z6yFOZZjiEgGbOqUkeCOyCOQ2Nkoguyb8tFnI
5EpcwUW3oa1J+4CJYEy5JozXSG8b36qgBx2iK4q3OmUUXDC7qfLXmwN5k4gFifektb68SsrjOhWK
ySTZgDSCGqaqxLiFLepSwbknbWMCepL+agVSUxDw1Rh2PQF6vo5P88KkzBzGD8HMcVrcQEBzz/KO
luN5UxoNPr6oKDbEUmMJh6DKy0ITP3HdM/e8wwCIhW0mqjF1KMKc8g3ulJWq4kW192W4dYl76qm/
oQx3cjp4FlIMjUDC61KAgzGl/wa3V8kCygfbWzy1799MF9/VXgQ6k1Q/aFkdNfE9MjS2W0r7C4iy
Vt/WlN//kONqqSYPXW4t/qchDA6YXr0JnHt8v9Z+76NZuKh3VmQtJmP2Zg6/m5OxH1tf6F2QPexs
7O+0tECjDc2B8zeILDoUUqew7/0LvE49i1tJzP8F1nuf5MVJi9/wG058MBUlClc/IamlXzJz4WPE
rfXFmg/a86/y+2ASFxZsQauNUhQWmfuF0tIZ8II+3nk1qtPkUwEciTvF0MVjg2Yzf3RycYHRVXp6
c4FakdOHYaLBdT/rtDxM8eTyTGmSSuKZgPin3wWoTxg3ksOv8CZaKvOrQ3QSJj66q+oUbGDjuGxo
f70SC3AItqk3s/Ec4ym3bwE72R7q21dfaNCqasEQM1am1zXU9NZJ8olA3i5LmDgxrJoaGPDXFEqZ
IxtHcXuClHRiDQeMd2tN7F8pNVs6y17XskOrPtJfZ6vYI1VLjTJHI23qL2RCPq9juT6BpwFj+4LI
QCiO0nbcAKj1JfzJNIEPjWbp6zTWBTAGXSJBgHokikrIddWb9MEJ8LK2Tsn2Q6+wa/bZWGjw8QMl
l7GsrT7norooXDwUYoIpvggcwKFhFPOOWIe2LAj11D3u2zannXuNVlYxiNSEXes4r+ctaURSMLD4
3Fgl9oJZ5j/gKO9yiP3VfEb+JpE4eyv3Kzv80z/Oz8zEtGN2aUo5E3QKhcVIqY693D0DmCAKYYz5
E0pP2xQaiRRwmwMpKgbty3vY8wgOPt6JYwtaYChvshO9LUceTdN3t5JfKGL4daUZ52F/Nt/lImfX
b30TRbdQrVv/Hob5Z+RQMr/9bGwgzcALNeGzIkR5M6z5zUj8gwyaEwSmgcOrl5Azujlx7M1G+StV
Arcf9YCMU1Y0R6aTP165JmNup1DFHuJ0IgXHlkh34AV5IfJpklNNvxwV6RZn/zDRzXqc9w50yAyB
Ql3GWMWilDpdpTTJUtk8HXV9sHIHV2FMMvtc3gbC6Ype4L5ORr5k3QuW6K9qiBpHyqtemPO6Dxmo
S32QdlO80chPr81VHukW9zAa0qsi61cCFlfa3owC42lqhZyU87KLrwFTUsnIe71f0na7yK5lGMB+
hEBKU2JD1XhCTNBe2HIoHPfNaq4xyR2mO+/9n4kXIb2O8JhNQDfz6GUnPTMuqEJxokKfbF6nuChh
5hfuM0PH4l64Cygmy41Y7HdBHVjc8GV4DREbE+cCrc79/9Gm9dgVBzcZS0v4xchWyj+ckjh7e/qv
H6tTcn2kzijGi8PxTELB2gyn3NUCCaRkgbLgSrwNusS8b8159Ylo9qbYLpRhfI5VNZA+5+/disTH
4UTKnXAczbBRzwXnazZ2qTeuKHmIVvI165gT1ipO4qTJt8U4R7EaKAvejSwTAwpFOZEirDhQ+GL+
B6/c2LLLTQWe6EUJJCuFwdmqC8A52w7ZN/Er87HWfdzlqr1iZuM6FVbZqQh/pE78VCDpN+1EH6+l
Mdw7qlhiA3kwzJSD/3gy1lsKOAxGqRISZuL85LxsinpnysQd+sGdLAhOlpeDsUzDYmdElRhR7Opu
8qymIBPS14foODq3Fs0weGEs5+kQWXU6rqfnEXGOa+6s7MGMUoUhqL1PDEUzdyFrUirjZB3Wjob3
rxN+qHkynwxJz3NP8ggctKDaQo2Zd859gMKaLVIC/VRQYMwXPKW2itwaJ7GcEcjkLYWT6zD+KOQD
Ya/BUa48x1CVt0D7PSipegZ+twc3aI8kCK0365yixbWCyqazuYhipF4LF3ZlYa3kYYAQOsZrcBxo
oelNjJxouvZPtGn3ibkTTRPHYW0+B6VxZuMq59ygNdC/IjyJI/8XGzn8U4ASxCDoY5C5C3GR1oWZ
U7OpX1T1EqJKrERHKIpuc/xJcuTSkeTY6IJJvMTZ6oDcYxirI3nuZkyqZIIuOZqPVReBL+obab8j
nUFlaeSAZyF3HklWrs8L+Fgbz6Oi3vhvBf0unwyMvwt5AkZ/TMkPkcfuX9c5tO2SNfUDBmPV+4/x
TKymdXEnJSnm3OGkX43o5pxJuPSWlWuaDChiqM+04UC7TLPaTe/u+ghRRtjE4aD4hAYRZeubaie1
hx83o9w2x0kylXW7zUxWWuPXCK0cd18fc51ez06JJj002eZtyz9d9BwWiaJItVuz6UBVR+eJtx0E
vpfmMOACV7Y7lcFKwAkd2L3HEu3Bh7aTqDV2773LUojNdK45i6/GyUyx6QSJkPlU3e6IPYrSw6zt
7m/t+O2OUkxUYW+QStWfKzSCZVU7L2QiY+2xYEXdWQOy+fWi/XHio26NwkQwuKebH2BKkoTOQDZv
+ObFe2HVQCJNQcxeLjAVcRS/7ZbLezmBTUwT6A14LdjjYHNEpSS7gwmL7lEbwY5zMFff6M6oMm64
uEid7Yhxh39MoOhXuhhgPg7tbztsC/iI5wWcQXoRJSVZq3k4aVmjkNrKOjbgf2PbcnoT2izegw6q
ZrLc2hkg10jUr9XZxxT/VRA8ZcCSI26xXRSg2GmXD+SEMgHO+x/0xrPfgDOjAPKUCeFiS1QC78H6
saEnjRa8AqZRrfzkimyMnkaJZgAbaW5HMXAlP05eN4LUSYeUEM0xpOxpprEi3XXPD/YQN8wxnVtY
1xIC/wI0ZllZuZCTtYjEdcnyHSzZEFw2ct46qlYgoN0wqfXFUec1VgUGH+h5TwAvkryGcnK9qcyh
tE+RiaKnAAIuYYEs3zH0PCxVlTtA6lwHy60+R7FTOztLEmF3yHXcdpmwAVjGyljyv3NEvuxEjDx6
yBz6eiqa0J/AxOAsdsfdlB8CxK7WVOifXAUWRaWp0gYonqXqBWuY8OyaAq9npHb+YfGPX4cb38UX
Z+SEvw6AC0e9NHAatUegIqOFXiPgZ7WG4H1tAP/VirXyaV6cNmdzKyAzZR1OGoaTW1fYTGPIQenE
hPuahRcMwT8U99d+jlJ1SmQqenaFQqcN1c3sNUkzS/nM1UsZfrjnmV+qxFkUYwj3QDzomWivBAwq
wA5GqjpqEMgZDzTZa4xLaqvMNt9qvfSqHjtwuJ2IxVyUthjhTck96Q1RR9wH1zsGorA5vrLUKhEO
D/hf5ygNccZDs1/A/Ut3K3170oGIY9Jlca/e5IspAU89IrybGuZXyWrO1dl466/p345/bQ5VGaZt
jIDNkRk4fDpF8ow1sIBTgIDrIhESEzj4sRvzpsCteem6qI9chN19bc0O+2BqyW4as+xg5TtYUoBD
rlShizyHUxLHdrOIXwMJha33R+RNkoPVS1bkmpQaNfUK35b+uSCB3HcmA1pY+M8o7hdKNnWKpe/6
5cp8DYhOutqGFKx9qUGyA2FoY+0ccABxYAu4JBzB9OZ5F+3wpOwqFQcGTDF7LvGD0ANeRL491fwd
RnHGQsEJk6HoXcNMJv9hePWIUDh/mwm/JrciUvXHoo9k/RLzUlcJ2hZBpuXTDmu+/OpE1G6z/HU9
hKmjT7h/MNfiN8UUktbQx8XgnRSsTA4ISxYGEiFI5sueK5EJ8iKD35GFeVrZcW9ey8Tk58Ryru8n
tKzJy78u9QvIFzBwekx2hGjaiW8pXz4IM1yGgXcluUvyfrhAjQCbHljdacKFYh2UDhk9QpLYRyOQ
sAgKqxVQIL7/kgipPlP6yaARQhf7zjYBS1yhMP02gtGAr9qPMKbNk4FqQKV3NABx6atefpqkVQpO
6LqavhVzatiRvDNgXq+tSjw58On9RQYycVZOJr90HJMU5+IXzGn538h6uCbOixMGttp/7FnwrF2k
UHZMqUP+GGDbSPshz/ADGL9uPIyqYzViNbzxzWLTitruyj3r/ZpLNKhcLvLrvl7sSmlBiM/j//9a
kBnZM940GoYpzQsSF1sgxx7dRatlYpZFsrBH1khiEHqBu5zZezFS2d+xFc0Dbe8VLq8kkW/i0QX+
PWPRBuxj072ygG1CNEsfI/lGWRRjJbexmteNXWXelpg4sdpZGCi1GALPtJaTP5g3+0cfYZKDhvGB
+r/m41F9pGVjUijPpOOlaVJhQQ9iJVG+3EkzwMjf6tmNn1IDSUsnhb4pFMpN3k5dbIvR5wCTWFp7
IQ3ZCTJSIA1/5aFRjKhU8a9I2J3dixieqDu64EbzkvEJ4n3RpaCsQzntqMGzfxBlvzOt2kwLBsfL
cBf56lq+q45IVNazZjb1E7pnidiprGtcbNbR55L9XCmM2HBkKFwXs5oGqvqGiRCVCe3S37py2abC
pn5UCitcyji0b5zub4LhE77OLdWAfQY1Am2xdS7cd7MkdfRoTWdHikjyH5ywFVbcvEq2m9Sg+ieZ
mN5PHy/ecakntwtzfmajOQL/IS7YlOMrrQRShSHS5MNPIJYc9zgywtDgWNEq3+Ua9lamy/DSWUzk
EEEYgghjHdNyFCEpFzcCHbKQNIZImnD6SKTekXoPjL9UL3SbiFICnF93soiMgXknKlxDc3fSjqKY
0WlckFRzHdnmCaH1wsjGmFrG9zLz1F3v2rEb/lXWWT+UZLwSZTI7TVLZ20VOqf0Ot4zw0fyLle2+
mKwfy1fzx6nz8FOcThMVIUHbt+gqgYBnb5ScFnMLhlQ25As8N/YwTcyOwJO6t+ZnfRaBR3K6+Boh
d7fClQPHUWQDFErSTu0rNwKDdZ2psb+ovBS41RmhDNkmofz1IkW3pieLcX+Jm0hkhpfxShBPB/30
zuKtPWCsXoonbYayeBElPOTE59u+4ED+mAKMRsKrT636esfGgqglUBExJ6rp836f/qbyXMVbT1xE
L/qPfeboYbSZDSWzqtCKjKeBHHSh0lu6At9dh8lmcJFJcxhadkvwdRLy+r3FcN2bJsiZwl4RPKCl
Tn0Ej4ZJRZT+R8plxZbXahrlpcPUjFlUcDHIM4sgNhUgNgiU/iGCNoAydHCabmpEkLsUyaGgU56j
JqVKjb+ZnD5UVyUxfgPyDEw6rRd/Zm0b/09n3AlGVXu3zWcIutKkgOjr29yvwBUc3BcanwDsu8g5
oMH15nDyFC0YYr9wHQsxfXPK9ZHxysk7TjRBh2H3MtP0Y5HEsyhmXcvkJ6yXiIA2m4H9QLCwaz0Y
q99abTTk3RQfhfLZIDLZ6WgfJvLIfggJreThUE/XtnORXUsRQgBiM4axL7alaghEMO/fnHNaRBat
A5i3+/dOM1gcNx0bzQZuU3kdOnKW2PoyokfbW3DVPSjgErwV/UxpB6JEYEy5xnvA3rWXq/R7TZ8C
SDAhJnDmh1ktSGD7zm6npwwI1GKZIpRXaILv+RlFMg+fOYlxk6fx7dLs705kQNOLYmimlZiRtq4I
2tSKJdA4ahc+NPqk/Il0ON+hpMbWeOHBSJ9JqrODfXhImqs/Fgp2pAqNSl0mAS3KLgJhsieBlqer
uehk1L/h4q92zJHrtvKcFI8ofOKvIXRw8uF57PaQz748LjYbN34DTp2p0XBBqhnREHSm+4mHngRb
s8yyaEE0tJJ1/wTf1ZveTmmf44Qb/z4d5zK831nOc+a2QfBwfhWm9M1PcsgrKZFUiNlQ6/B1Kia4
LZUE78YcHG0ivLs5GnbRJqSIxfRkUVb4p6oefJSjK2r4JVNVM5ci7YhvFows+cD3JOSg+fwFtzFT
j62Lb9nWx22zxu51hT5thmR8Rz2Db3XIMTIOfj3vlvo9rxpjpmxSy6QzkSG7z1C74u8n5ySHQ8sD
07EFzAKHnXGgLy7x6JsCD6BEIjQzFaXI6TZ4jRFX30BmbYUR4g9ZTvPiOGwhTMxyOTkFuOBg2g/A
pwvxtA9qmaRg5Gh7sTWPLLUUDgqcS66ii5B465/hzph62rcSzo5Mgr40+iDXpnMuSwurVYM0cPrQ
1iqJyyzKggZs9CU4IDJP3NwUdViMKwcQglcB1ylflVcoPrKKavkHvVU9LYQPIPPz6OGzliqgV1BM
O/pBIJvtoBD8Jly+KB/tmJJqAEstDTZXwZi7TBdOPh8XL0+it9kUy7pHwJS74YTNE4x66bPA/o93
FbHdWRFCmGRnO2+rX3Wun988nZXlD68qmtyk2D03lw6aeGDBal/Ff8Tr3uceoIbH0FbmgrllIpf8
mMDqHWs5ne53+xIqnm4c+TlyefTi1Sw8PhpgUzVs8vT6cobhaDMhEbvQDWJ4wtqDXcCAQhOqpNGZ
aKNgT35WGfqF4W3qqagoKUbO06GxXJQ2HQaUfyxVZPkixWkbGcrAwx0lWaqXqiWpoD4w1XdndOWI
O6TXjkDLyrBIDurvziiWQVexbBeuE60IoFjKm7LS6lMZ+oHR88kzsQ8JRb/xi0TvmDvUcp7es1+I
cFpIK/pfporLjOBREXc+gv23y7ZNOjW5uhFCs69nWSHd9HRf3ezfIRkJsFfMcKnunlR6VXFDEcQ3
DqUrUY/Bhmg/F171KXav3/MCr0gEhvcnTDy5+/f3Z4jLehqILBbZIEykFjeUSA6dcLMn0G812Aok
telIz5IBQ/jAaic3iRysnFs40vFoz6glF/E03+GARSpro7cEkR5NW7IwXWDCRf4Hl5/k3xPfLGMv
8uoyQITwFTPbkGzibes4IA1PZuRz3RODlI1P3vnWNzBkKqi2SEKFeN+xMUSrpSPPQyz7qefhkBlA
seyfrMCTOidnaPDZTQoBxmyzeAUw/dbwHSDqgRH3T2pdFsSdzWmk3yzB4LjOJhs128QfFyxBo3w8
lE0pVg4m5J5jGuMHAATU3gWG1wxsNAolGr66522IkyyZ8rcHTWmUBkkbtgyNjjyMKM/tWdifMlSu
6G3NYuANm3ykxD00/xZJnaT9XvICjidthjtRBC4xPOog7PsvaZ2Am+RMry7jm0YOgSNcDrgiYkwu
Hz4Q21aAbfQH5Q8FNkMuP6G62sWtKUyJLkCh6W5x9DFKoCb03FsLFQM/5/svdqJm3rtfVV2fETgM
FugI+dCmE8u9KB+Knx7/5MrcPCrlQAO+/HkaqHotv9GnAt8p3NKAynnSiAqTDAP0kmNVy4LuLpKP
PrJ1OXl9siLr+W9Z8/GPQadhLt1atxUsNEUYcYO+1RUdVEC/mmGq9RtBwu1kVU4kO7ZZZ7YzERhL
isQM7KgryoDKGQ6CUBsqptOZcCLclalmmEfq/MLDRfKGC+obZnG74yixqcNY02t3yTOJEotxz2T0
Jkt95TO4wOFycX0ftdBKxdEZtMwAwyoF8L6OTwjio2iQnqSGbjVaV0T6VddvOSirSNb/B77b+Dqc
EYhZ79UeqrHBATD67OYeK7qNTBgfJFHIUvHsBk0KpMy7ZqJgEZ/1GQrfYoBKkv30XoAqDM3gG8A2
MAkfgdPM1p8Xm+BYQJf7ctTGzUKrVJlooaio9E2hCfrHGIAj26YWau00TFlwgIN5ZE+r1VxU3GwP
Vb/3lrvQT76Wyw7UdGFC3/h3GNWHMLDWYDGdD4NYN6hfWmCHwMXDj4VJogupZsl4C9+fWtnQtfGC
jD1c6URycS4y8sooNomEzeENYoO1ANNIgeinFF8/Ot4gTVMBe9Qzoi0LxHQN/ySm9bS6qWSGTz5C
bgtSFBoFAcUIkQmxTOPJNgl09lZ1iU6lXUtn2rpNWGjJMXkmDPJQ0feuwZw5Ak4EytIAgm3Mfm9E
WOhNp6oKupbThEKEBgGf13fXqlMYWb7JSKjaYOUAxyf5m6G0wwdYa0lBEg+lVPKx42R+8NjOFaYC
PjXCv7w4Ocx8JuYyqV8K14ulWEoOoqulpLXoArcH/s+Cmn7Iw5KR5EJ1gQkCDvyYnoTi6ijlfJ/Q
G9Pd8xXN+hDFQ61+0s5ok3bt4YqskXVhTter2wyTtulbIDV09pzrZ5b5me/Fwnp7/uLxSFzn4O+j
ZpaZ+3c6vKzM7ONi038w3eamDXjU/FRdDVMqT5g2lIXfZRpkW97MovbpZYAN93ti396ZxRHjFl9+
BcW87FkKd/XXnlpCddnOX0qQbAg21exFD0eVylMvADC/PopJu6dos/L7ZgKcO5hmacxM7IpK6GkT
ScPPR5Nf6Pw7ZM+ORChMLxC2HzZvGky+WZPgze+PGpukR0Wop/WUqBsES/WExYfXUIINu9MqDXQN
bcYBIss787M9wCkVdNBpLnETKb68l/QWcZBmRtgbnskSmvnbw0NRkQiKs9q3Xxfrkezb/EygG5CJ
z2kAssBgN4Ern7Qb5+AaSCyG6Ry8NKGvVExuV4GI+zZ7lYHPnckLgrXESsLd7PP1avWKQAWRKef8
WRCtsznd/zIAVGcEtsq9nE5TjNMFpgsfM1TuBXg9pYhb7wiXBobbP7Bb/THd7JN05UfSSRn5ClXb
oZB685/lYkk5J/r3AQ0JrNxB220EYHyNV6f8n6Z9fZKnXWebHmsSPdO9i9+nkJL92U+zkjvkf2+t
ywboIV4mvkmtzNEG73rgfs2tVTACLBfeLT2CC3o9IegkwJkFTpU3lTdduP8Mt0KWQOn2zACn2U/e
tfUTBDvajRgA5XefSx6o/i0BPjujQL/ygDWvkad8+4b+S5S4lSq5XskKkTLQmJXuh5NXLGZqkEhQ
pPTCckBS/Hq4NITi9Ct7D9lRwHeI6MfNyzJV+309c4grSc3xqSV/CBQFB1bNbOCjGvX8Ome3orjS
xNDejr1AE+0aa6cgoMAQvfkK8X6+DsawOPjr65t+I4vdkaKJ/lCNkIOXLSZwxeb4rU8nbSLZ3GXF
mPCXVSPt+k37hM3f4uAfEljjKyHZntSk/k+UFhkbqs7DdI0BN9qw2QoPSr2YXp5NHFqE+XjCIA3B
aCMs3gX64/nCO36SrWVxFzVG347UV5I4ieueM0y4aAgsmU+AiDUDJlIBd+orqgELefzqi7D2BMam
EQ1WwvsLxAt1BjARQISX3JBWyvtfOnqIap5JtuZRlx6hNVg9+P3cuByJr9EPiFZonDVTvocf8n5v
t6v7EiZZSBf5wGdwNyu0wrY8iXNyBvcdlcC0VOx7VJTY8ncD8T71oL8rxsXgStPBPhpitEQfnYrQ
sSlJ1LgSG+1AB13osnoVEdjOY9yPYq90i6P1CuYe4k3ARpP8Up/BzeaWk2OQWhckPNTUOgA73rcD
DDD3Y0QLYsqN856k6svr6Le/ONXLCHFGYpv6crAUsvXQ/2qkUbQeP8nt0hR7HNrZXhx/E5xJo06c
CY3UVYQ7ZnvVfASXeBzx4zv7xeasjrrDaSaCW+seEns202N//J9QaNyxTHXWCdl6G3jjOxtxnWBi
wyL/6laOqqPCo5P5N+UNGTDvCqGm/XUz+G4bM9owZ4pSIVZFgHRjulPeB1tXbPSGyNR4zUzHF7Kj
GTnGV2/H0optYnjRp+pR4i9kzgWP5579WPM7May5efxrVprlu3RbrIbf9WlDC7z595Qbem6lhn3u
404dbeCtNMo2YWt9STlqNKHbFbQaxVKtoi1hVVcoaQdLy0fXIIsFck4w5Cg5WUkgWYoRby0Y+p5c
DZ3Ik3QYY9bChK47Z6oVdkWyd5lYBMcQ9uCgnlsVOAIm7aVJozViLrxUJQHemfvb+lJtOxqKRz6t
L5UH1yTPZPZpe5aAkGZ1Jynp6FYlX9SJIIyE4bOr+b3mDhiXK9jCiPsgFLnmOwS/MPlAiEjV5/Vi
sA8NPs0GvorNpN5Ys6swDepBZEKY2189wpb9Lhs1P+t2NOyosxONRmnlIvm2Jd/dIKoCGgpnTo8m
vkdYmsTSf00/lP/6P5wCMH757RhmBsc+NhgJ1CLL6X27FQXH4HD3epXAYTZLreuEv300wIbeeQz9
1sLMayv3c3/bb9AjSr9ufAVtoR9r34tKtokuZClNSM6NgRL+LeEiqfwIMb4UEXgz80ptE8NC9MlH
aPuVb/EiQxHWAEi9eVBrxxgb0/UdS910JH0AV5Wzou+yqzbvBBX2sI7sfh8uykijRe/9n9mEqoDU
wTcOquu4/qgfVVlx43TDM3kt9Q4PFe8de2LnZAvZflzGwWCAFUTGttsoDP1HMC9Yln+KlnD6BQrt
weKR4pw2LNR67Nt4Qm6kA4JiClMwjKh7yWk4amITMjPmyDcVmHrKi0ZDQq/5WQh1MWRFsJ45WqfA
7eJfmLnXswNJBZVXhlkKYw4GF8bchL/xscI4zlRq3pQSqox65w/gh2DlvLN8fLC0rvhuAG3EV0uM
ASl0HdoTzLj9Ds31ckVhmE2s60Dq78635wXeTsfFUYH6P1QlBZUBJfkgXUv6xkva/qVcglzi3fWj
ViaLAWzUgH2UnyS72A6peCZYskMTGavhJaQBKTfIWWjHzjHELVQ5dnIWlyQU619SSAYZtNpHbvzj
/d5KXClePiUCLKRo5qSJ7l0ffxaVt1WE6CwPa6/zM2Qy2yPfA616VFOl6NhK80Fi7/4tGCEjNM17
l7jzr/ENyJZpa1QBEa4+KjvVSa4wKp7BMW82OxWxjfu5HBP1L/8z9TRZ020YxM6dPk1Yy4/X9qTk
CwG0Zbgeyf25YfBw8NftBiA16D30h5w1OSU3h0Nsgwoefj7v8nS4l4feW81hDVSYr/kN5ZOMgDYl
Bo5aYu+BX7S/qudkdhrBePlcmEQwpVaQyaApkRsFr7D+xGJyaeXHiyxYoQwf5AGieXcZTsSTXpTj
/FMu3I/ptt1gblAZGrLDLLqy5ufhYeuD29JcrQWxNqZc3WP9FMua5RJgMzYVv2Esg3jGhyz+V/FJ
C6dfl0Mi4xQCdNYkE9erR5pp6ChNpUJ5fqlf2mTfs//eCB51EHENHcPov7Jmg6NJRwksr9RHG+mE
BTdRT4dbalxpO1LdN4NGKlKIpH2+vMa5QGTogjJ0p02N1/xnfRg07S5qVsQLtcNpf/aexOnLk5hq
vBvFHiKokAz9m05NTeqydc38fS1QfSvJz+GVyovVpUFQkND2qOuIPNerS9ujYO4EwZPpp9gDUr7p
V8mR/AUQX6xYEkRFvAGs9pRmHwHI+o7o/MvKg2hZ6gTx628U4mfXUhuyjO+TeDvCJPjicDgjdUcV
HK2hMGtGpbZmFQvaMCLqx/UG72y/rJKHHnGTkj2qlBDvoWEo9Ppth+gvO9aFpBX5IRImMKDQVCsQ
JpmU3CZ/zNc1ZogVvKm+kbvBn+R/f5lgr8jp7h5zBu3qX1D9nQRSkfiMQgszi1XgXYXNnixCxZD0
eyky6PzcwzgTLZ0StDuGAx9rTbpZfRPRW8r66ssWT2GQyJEBWwEBn5HcUg6RXpzM1xm2dh8/P5EM
251gtaw0qXIt4iqCD1gZ02wGmUXxILhmDjSzHTpkzZ9Ldm6UKeXntfEp2EgfpeXLkEr/FlDS7G+W
5jQjD6stF0em86t+kozpi4cPCp/+eLc7fjsr+zVXU/EJ76IVU2oij+s/pLvq+BO8lD/spnTzWN56
KN+ik8oEaJrF5OzXoNMAshnJr94Q1gf23nHjDm7E4UdXgLX8X9dpqxbscvNDXjqyk40hWhGDry3d
0AyCe3ph6eBpTp1OmRwsQlGOmsirT75njv7hXdNGBiheV7hSndTvlcyQhihhFXbtRP6jSPVXW41Z
tCKys/qvQlvkcLsXJEi9K9UFKEAQu1M1CrH5nUpU4ZTpVyHueDI7tlIcfXAxvGHwiu16k43kwvGm
p5IRLsV9/R697+VehJQNQCCWWhiLm5Va53zYm8Fk681utsPqGUFx/B9yr63zaN3aS1LQF+14BraL
XMriAr6nzU0eoIFTJ8Uwdd5cH5mJNuB8Vl5P2rRcrBbp5T4JuYDc6rBntq1m+Lpz9PtfMyGNakA2
2u7pQ94Vf+xsZw1fOG8KLriG+h91oKo0SPYui9OT54gnclNX/2Iz4ySnRdIdyK+dMzdohBcoMh2B
+AdQCYD2eJiHhwjIEo17X8XWMZikvlC29Jl/rX3chOgLUiZfpq598CZHOO3vhNUTLFp2dfUKuIqd
OpxbBZlPWNsMlJKMjEis25I+p3h6bXB3I8WyOgamMRzGNUF1d2wScJAmYqeeOQAktP9bgZlvqvLw
7xUTFP4dV/OlCrebogMJX64KNo1CmH5k6dLZJW59MicKVNp2nqOQ3KVDEnv0XHHs5RIMlDAEnX2t
vlhQZdJZPlcFUgqVClN+Aa00sC9jgxKyD3KfoFOvixHvK+F6HBHYQl5eXUVMFvNxSVJqVphIhTve
Vtg8dyysCFflyXVWrMVUwntW9gGg9sMbI5apyXngJhJZPsFSoTGk3hCIpyqlELM0gZkjkQkOosEz
WlsCKBN1EQJSJUH6zKb1BVcucfJvdgnB6YVzvi3rL0OKklnVMrvkLy/L4da87SULM2Yem/gZXDhj
QX6Szz2x949s2r3UA1Mdrhc+s4YByikIiA75snBaOFTpKZ+BwoQNrSPIrefGTwZF8RMw6iRkcwKV
0JOFVmL9qcg75pMu8YVXmpianw6sueSpb0Re+mbkxH8G3tOS4xIhnkO6hnfvCHzBsICfvWVysr+8
KF/AyjOP2ZfwkBeYBjHBKyEnrK1ByBuvIgnxieh4+Lm+6HRdt3t+OWuWO8qjXp1U/KC8J+13raEL
YwzO1Lh8HSHZgPGv4Sh3A2EUqY0ZkfZNfdILgU5ONAUGB5YtQjtlqcNxWVpDzm1nEK9GPj2FwtxY
EZehi3pErM88LoBLRhbodPz193v5z3vIORzUBXr6ofdIUzycHvqKhMeWl6V3aSwLnNLZ7n4lRAUw
++pJ+gMknn8v9TetbLiEuELDnB1PQV3Ad9GUdNtThrQYSTu/g5fsX1DOSmYaPzR8KBKdnR+TzMbZ
y4rHAPrfTQp7mde7jvF1WbvmmnpacylBtJVqy5wWqZiIgRBKwJpaVqVUpbKxv3XQVMWSjA/Ci1EZ
DZtUUleFq3fLpcloaZ+pQq3SKO1vERPT6hUOzSco5BaN6OGviHL+q9LLOsm8eG3y5AMabKK7sznX
uDIeVnnuaYsbXSVfzfMJxbfxz2qsTG5JOXrdqQ7BXGHx7eCuNu1StIGRFMr9uGR21qLr63nj+6Vi
0VzL5M67u/xACsee1S33Am+7uJZTGqajYW9lPYZSDCmRDeyaVB1JIV3AS/dcmoDUJBHHl7iMJSaC
dTWW5RX3aoIttnSiipcKS47SY+X8HLDaLQ9FNOb2OeyMwgk7/UzDSRLP9CjxI94cagLy6kYPZ6d0
O244rJYka4MBwSTpD0M68Qrggzoio5WRnBhOmR9BMkC2/i/luKgPYYBPd1cZQBpNVwnSjZhqNLGK
0gqbIQp/w5sf/RO3jYUgisfjpLGU/waR0dD4tZ/L/EJjWQ5EE8WWYgSI0G3tq2IY3gY+MBNQHXmU
9hmvm+9qFMOs2ZCtQ1AmNTgxybaGSb30qVlEUqBt5Ym/42QrZPy4mDCbm5u0Ju6RLTLv1sL4AbPQ
cJOTuQUYaXL7Dqlcpl293SORm/fKB+2qKa1zQ3l1256OC9n9cafoLyX/8cT4jcWCt3XW9zP+p6AL
L0GkupsEO2CKJJ1dudaSi9oaTu/9mdJ/n2PXruDo9xlsEUcns8LYuzkCi/12N/cq29pKr5UvHjBt
PHR6q5ORib0OATXAnzzb/d0gIk4Red4jXhW4IjasY2gN6RSNL9g/NY9uMVNKfGdVfeix1D1H4S0b
OmoH/kC1WXMotrYMaOjTkYCHyHOXb3D3vNU6kZhkmwBChmJsP90Jsjyi19P009YknI5/k3OUc2Cx
bIgtJ0CTK1IbDRpmSbmROxVtg55VLGoxrEnt3vFgqvoEJX6KEtIWp8zBhDqIoa/lJxfPL3njpPPF
9eGWzqMkmveMpi92yqz4gNAUYIkz4Rzc5USGz4xdkeJuLoc6WBHlMC/V+wyCIrLENv6A149zzOk5
4Qj9pcvmUdTPNyCaBB2V47jlBHhqfnFIg+oPIBbHkI2IGTDrfjD22CViwmyvRv/ZOCUonxdbbxUq
d45C2rO5bi+OSoyt5MKsQ/iPp21yoAW0m+1VAnKjiOvuSRwWg4XVS83iB2GM2CGcHVrV6qCXwOtQ
9XollOE62bfHy1j/RWSFFqZvJtonmeBimcbyb3t0VAOUhdwC/diIi1x6zbD7cpU8WAnQkBd5Ma5A
WO/+IZbduv8japnhlAXYGHvsdasmLFs7b/ew+2I5mbioIgcav2E34oYs9wFRWYh83GFZzOgjbHLZ
hmJibwPmAOTeJ/HPVSmjvlNRn1UGesu6cMLg4X+vS0vzjXEKxWpyFAwpELs4xBKiSdyG0GE75pst
bJROFYDQQMdHwGqpAsXSAlYf2ZAwepqV/Y17icSfdWxOPKmbnu4GhXSivUJekOOFQmdpowP7VHhP
2Y1GLnNtvhhkFK+u8K/jCDoaj8rnTINKuZyCwzXgMKbKi+55jvlpsH1q8S2iPnvyWMnx3yX4m1Vi
Vf2WOCZEhkUJhwuj3i1xUBV2bhpS5M8ppSSI+qQ1FxMgRuDYMihXg/0XlXkUGkTnAm91pv1sJvZm
2hFnJG4tJzR/QopR9yT7pBpQKyc/35GxBczKN1YEI/fE7awy2n8pSHSovQGNMhZv0FQQvMWdsr5t
ORSiylCcMYG+lxrjFG6xKUJrSLqAH7NifMSdl77+jkiM83MWbh+8Rwr/X0F8TmSG86VzWiFQXf2o
eNs0AUCvT4rbyQ3uQojVap17ikwqQwaKzRBcnBVdc4AOvU4kct7QORQbLIftMs9lHTdKS8hkbmJT
cPFL9sVCICOcq8juFR8FAaeP+UHN4qdyZYLS5AOpBwJVUv6omj158QLExBuVGI4/j5iJbphbBAeF
mKUrkSzgxEShqGJZr0J/QjFWJRG+Fr5+tNTUTCNiI0txGkoV1stkJZR6kGrvL4Atog2VFPXdVRrp
IaZr1zWmuLYM4yTb6LfdKyh8IaFAQgph+ObUYD3n6XGonlNm07+AFO9QqddvfSlXfP5wspLpQLti
Z5DYDpwu6Vpr9fBEz7fb5zO/4GUwXM3dDgjrSjW1F0x36jscGKNr1gnacfvoOPsAaIS86gtCHe1p
+1VevD9XwxiaNIzI2lBgDwsO4MKG3z2UMyPCZ1eY1GcaDbmtSSYMWZVkEHI7q7o1EcsnmMpy1rEs
xG88QECN+cHY28z8K4hnTXeLeQAnp1cXbKexp9dLS3taOQhPdyhn3NVHUgr3Uo1LfiCZp4wbRy5f
gDBei53F7tg3jX1HDiOtBBALMRCXIq95jeJ62g1A1Yr9xWDTSb1qUFtfqyWj9evwKuzlEfFXhfMK
Zel3/T4CpxzDhcFyJaC+OtiLfYwikE8A3971FhFbqu4HXBVYbo6nC4/tlR50aXcpIyoQNK0tLeEa
DZPpZF8U8XGkFqdqmYy+CQIq88uB9kzyVuyRuiRNcC6lRpql9tTSdUdf4qnQfOnV2n2tjcqqw/FC
UJBkouHepFUOhTztUjrg/6ecqPKvt33EeshY5FjJyKqYDvgDfJxlIJ6YzGgmu/I9a2zUMU/RxEna
w8tFJm4ERw7xX371ByX2yrwfbQcmdIuIZL+Tv8ukwCV5LPtScsBHkpQOt8dB2mzKFDQxUv4IUio2
Ey3Cm/A93bj/GyEOJwO+0kxFcH87A39AHkhIj5iuRNvDAPu+Nq7VbpbOAHysTw5KHKsdNAcxuCUv
vQfVyfPr6+e25V0WcK3sK7X7d5g4/N7EgA0X/J+0EyCoBe/mwzvoAHCXc+OliCLs5g/pUIqnfEbk
4YWwqJeMg9fMPRHEmUq+jJTNRF6c5KEIzu+TLvBWQfXA38eAU4ihydf/LFCNhCKUXrzcnogCwebk
hONTYHSPVcdvmXdA2FrGzVKPkTOsCw1Z7KGmQ/CmtY5A9D8ArG5SwBnK4nI0183cq06x/uqmLHxE
KYpJZnXAsMASFUUv0nk4GC9P9sEwVjhC+ByaloB4NG6WCCfy34eALU5SWRbywQi0moAquT9IThgj
Ocia5mPT8id7ojoSfTUan14djPJbI/idY9gPaa/UZH3LfZuq/4KwqvcN6EywTh0gX8PyaKKFQFtF
dyl9KZpm+zAHwiOrf787tTx+on8oQwttRE1r/vzqeXxZvDwpQ0g3chTeYwJ/cjoviD1gIFHu5aAE
VZgMi9yyf/E29HJhGGMEESJw6MqqCKwf8yn+kbJRwJei9SNRtSZiaFEpWWfLAjG17J33eGdc98+h
H77zfOvDi52xHIDQ52s4DFr6rc/0Ew/rK8k/aKOWTmbaO9Sir8Pkfvotd5DOx+U3E3fb+iQFFk+D
ZgaE5lhXeHwnHZy4xVCCEsAaOn+PMWQ3/1PFEiazFlDBCs1pmlp6SY/7H0lKKoHGO7puGTfeNcBF
iqRPe2sonWVmjPYHEhEp/kXfpC1xKtQPD0rrNu6akrWe04V2Km7zRKnsTanMPmRXVRLesmokYxe+
TdTP8y46GIXIZCyc+lfRCVfBlwNQCUqEnn1I8hvxwXyq6zySqS6Li7IoDqwJ8MPfhiltVJoFJgPF
SmlMedamiUkCv+xxZ63niAqn8UTVyLj4snHb6x512l6OQmHp0p0bKX4El6M628ElijsgewzFO366
Qgrrt9zaiTlqpYw2arSOK8FxFAZp37jgQtA0c/qySLP6lxjZV2TWJjkANnvjFG+lviYx6ET6CyF5
0KUsz2hR6gi7JbHEB/8cyg1OxV0RztzlgC5LumSZXE1/T0ap9cr3AcZax5RRUerax7s/UGi3EKhG
h4KjvZrkNrsK2AWQRo/NC9Wv1MkvMtlOC08oUZFL644oZytq5kWSXVqvbQ8ktyAU2FuugYFLHkQp
kIWD5qozs4XhQLXAlQGsHaVdRWNAnhwAMCqNlTjvxB1htZWSLkEzTaxsdVmOYLpFFasq72IZJtml
0uwBRLEFikekusOhjbkn18llLECPFaZWihF1lx/dO3u1SY4KU0kSLtmbp44shZbZxzXzNV0jpTgZ
hogRH9J4lJYeIwGCnpPRJtmZ0r9ELF2N0TQkKjcmF++JXj/c/p6um0GroWqGk9EVeQYvUbC51zam
h/CHrBTui+NJNHICWV5poi0NtVJLU97w+s4z6XO+ecYZ/udOVmUwucECAr7XUv6IbCtW+CAQwuvW
jtV9PVrv4ktgN1290VwFuTJKZwNxVgj9TMjCzhouTVnIl76dDp1gsGlM9Nb2HoAPYY6EbZMnFjku
e9yRZKg5ENHQ/rRNQ2STFNKzOseqVBrQ7mMvkmaU27ut0E3lJcyX7Uq5CTCcetQEXC8aeUEdXtA6
AzJh2NS9/C2AILDwPkexUjeRmOaHaQ+beQChEAEO9nAyqKmDKG02VS4VQd8mT1KNn3yX7oJL6Kcv
yuD+hqy+J8qf6ciw8gBlDjHBvJG3yb1g5rNdaFRDMjHHfbGnOWGo1gq9fcTe6joqxh/DUJzUhMll
wSJfcdK9fYr11X5Ukniy+hcRuilQVJREbUI2enbQnL3/UrXO2AWrTdi/S47SiPNpVPavwOPp37Vo
7PtoVjWPdenYMr0V177jMAVyI5JSiUw4VwkPDwz6SSC0MZYBo5z1+l9LXHOkXgsHLP8Cd7xmkyTL
Kiw0Qc1mW+v5sU9owaZziB8fpZfaNWjYiCN+3ocW1wUWnPmie0ui8GyR+EJKd7pHJ762kF9yRieB
a9H0yLIbijbCLFWzS3+T4nnOIt1n5STgdFvSvgBoqHTe0DQ36W/cleXJW5swJfJlopYs77EXxNqW
t1j+I3d1ODTgX1UEgCwQ6Y3JZrVZvF7iD47pPgXoPVBN2Rrd9vwqDZJ3FisdxOk5a61R4WUtxMWC
1qwFUVTuq5b78V8lzgdjQSkKXfvQVthU1Nk6dgLHv3v7H7d57NypJhDHFZOAWgWuDP5It3v3s+x1
0CDwj33hyBdjm/VyHAMB/fjbwqY/ehdzYvljdOWiYCV3x3ZoAFETbX5KoQqzkG25AxT1dXFfylci
xwIu48Xs1MqXW1GyrOGhYW+UJOeVQkVGmjHN4hO8vpOyFVMF2t9yUnD0Z7dwVUP5JIOobbOA9RFk
wpv7RJqHJ3IEY0tFqOHcYS/oEuQXujXOY5iEFO0xMhG7P6LjuFxoiTnlC9gkN92TdIvXZ6AXSZsA
vc9mNLDNlZ7dkDtd80DL+HcHFrsZNZz4D19IPyrrXmb60rYrzx2Ld6SXBNkjV/Vf2VgkNJyjwypK
eR8U1+szyQML+DZcO8AnAi+CFGNlH8/hanOFAuW7YYbuXg9kjYSnOIhTKOVB+sqtPwkcNQK9Fqwy
xdzKgS7FIbx7iAQYaChHWzyR9oZ/4OOvFvxa/ccfAj328iEyV93HCidaqH5QV1zMbn8uktUvN9QX
31CXzAfCYNuMhN7D9njBz00YIw+KtXAtn4vYk4ajNmfbbLkJh/dkxNumbJm3CwICSIcuocgx/avV
fQxxz/lZ79HhMs8esZX3sBXjYW0MhsGiT1pWNjrAeM5ZJ+HS3DEcBAKyUvkMBi5LPBNHzfGRPKIU
FJZeauAFvcJDg2vkOX4xFDx24rydnUioY2cerb3FMdAYkyNHT+yjJdc7S0BEJuwhEHTRu/2Bu5jk
q2Vz0dSZsTXgaCiMSSOC5q0JmdN4MzyAPZumXlSY3wlQFWCytims7VOiTcVfx+2TCxk6/9e2Pq1e
Njjv6O04C9+Fze8wKQZxxV9f1lQfufcG5HBt6F+gHJC1nNU/oOutRFO98OdjgkJzzh/uiNupXTcI
dMMUY2N5WPCYQvrmQT3ZZPGZEz2mrbaa6mifBhpta0L6KQ6iYPxGSfESPPSMdo+xI46dDiVPMJUe
M0noYvvF9FNT2J1U9VFaZ6dcIoT68NI2ObF5yGBpoWVCUyRzhWTsAaANNYzCuvIW0jCqgvKNgMx3
LlKyBPhnQq22OmRFtS2CdeCHra0Og8nY4VuE+2YNzkibD0GQl2siIN87SXBV78rz1OiirMDOn6gw
9co1WdxO8ivoH6Z90Ebo6qMOSxz67+vd/cI5ivVtB5E2lh/+qA5hVAlM9VhLwXtGxR5FzIoxqp1b
00TDhtPn3FdXtNCpViaITGVuQOt0SbTsMx87AKonqWOdqWavSWzsDNjSb30IbQtSU67T5QS8G8ND
UQbwdFmqzkJUOEnxVMdLl69pAVIzHs2grIsaiaJjzXEWbPby43SErThekZRJYTSXe/PcyDzhlt4t
iOJ8wGLeNvq7GYUPecYcG4CCjX7NrUGvABWafj3vBONLoye2k7YTAh3wjmX8TtygbDnCXG1XwA7Z
DOmwtr0s+hkhikBP31kBb5kwtpp1p9Z10IOVM9fMCm0eDmh8QuQTjmm+Cho+GcnnfOotOz9fRhKQ
ZIfSaPrrs7E5m3p55+F2ypd30A+2s/Sg+Cw1+irv9SQ/5fqoKXSWZVx2KkaVN3fl40dtqkZn3iYw
qw6FFAbe83F2RyrQfQvnoQoFczQj+J1TkYWbM0Rx+c41HHNSxAPrtJgZdtHJsA9T62bjEeV9bcO+
n6Op2c6lBTkQgLNJQwo1C+3ekyQcwzw+fxJSYVLdmIgYmtPdlV9K704Gmmuyxx6ba94VUWkBtPXo
aqwt3QCI+PGwROM6z3IHgMQly1/Lb918xZ1KXmZLuOYak/H+YjrmdT/3lIGXvTw8EDPmCXoHVou6
hELg1htJKK8B7ZQlQ14m6OGUs0JJ87RgI1gQf82kQECWmpJmnpu1Bt17VeUlrz7rtenBk0+aevU9
g9lrxyCnBlpCKEySCyZzS3+FZ74zs+Snmj2TSmphk3IMpDKnSxnIMxsYNaGjzhZlzB4cxQNxksYe
udPZ4LtBTH77EYtQj42FLB6xNM9UPbbWlC8BGffpOOuHbOUli/RrJ9ptmpQsiIQxRFwpYTUYIET7
nJyzehuJfstxQCWPtCl1BlRT6BPuAJFs6FCKf12W/qLeZ/qEWh4Th5QkVxa2UjmlqOoZf1z2nPzD
zf950ksL8qkPosfuCzpCFCCnzWLrpO0sxGCh66pNyF6P7Fu/pE5bH/zALlAdCCuJL8pfm++Pvob9
ZC89XIcFxMJd+7cfHduVxJsS/ta0K0zWUjc1bVqa3l2E3GnfliEBx/6vIsuKTn+FRCQWeNwZ7kD6
e19H/vIdnmL+C5k8KW/JLl0XeFs1m8JgGHQlvj+I8zccrzCLgsxnVNo7M1zyJ+xB/Wk1Fkz69Q5M
IPJAY8qkNgeyWzZzSzgP+Get6QwWjLHH2riwtc1bCyTmQuKAPjYlZC7X5jv53kDO9UqEQPH5WsHq
7ujYR8EAc0v+N7KnRscAMojkhOsyWqtDP+IEZ6iemq743+wNWIpDkzOCtWOKO08fmDRTkCxeHy6/
XlQNBegvZc56ledsZyPfIkm9O3whIUOoGJzYwYrgyB67N6w8czvTrabdosAOgAtdimWV6F8j3gAh
y1ura1WguZVDNx6gkiv4XntKjOAxMtJCndKc5aGa44RQsg2wrcoIVB0GNn0p+bwuVdogJhlfTjI6
B0V/cezjAZqZ4JBpKskQh7xSS5bj7G3/suK4sXJ6Jl/pGDOsNZs8/T35Yv5N/stY9v24S2xHdKrg
sjWXRfnX3JzJc6R1uhYKEfifN5F4fkRTTO5CvTpmnwWqN/IkXPx4erLZtQYP7G7pxMbofBQUqxJT
jQexmsQitDO7F5i6xKbDdEWUaj6xAtcdZ6icObZihIVubxqAI20uUSjtN+P0aVoztP+5ctiXzDRj
9hPkiqoTfyev7MDOHA/PvZQu/MBYtMQLgR3XFD4QnUOk5fTTlF4zXXAzmix1E0VxmultSBYVE1OJ
tuQL4HY4RcAtmzDwE2sTbQSbGROVJNPY91kUqNiL6jl1t3dPRX8yfx+RI2ux4jWRGYdiz0kJTCI3
LeWj+C8hjImM9ZrIfmJIrbxet2Zgz+ncsBLfZ/CgC2SgaO3/cbwJSsIQU6BEEXT/Pv2tgZPmwKs8
08tCdX68uIEoLjsEHbfMsevO5ABJrpN/0jphTD4ukMA08tXxDhmmY1t60TTGPilXR3vbGeXOtZJx
rTp1FJk7X++3ICAKmiZejfjjPesmqDFdGb1hSgQy2Dud3YFDDpHsudzJaanmBe8YJD3s+ZHjpKG1
ibMNyVjRvD+6sV/tbc9rxfRA3m3Kb+AHyoaaMsv5SdC2+gh8L7ojg+MDP5VaTmHnmMhvlvP8G0K5
YiG0afKvGl/9bXnGQMfI0WJ1jdQANBW8OzG3hqtCfYskoGSx3486Ft1NOOiT+/7kyhot37Ji97Xj
2+nWeVI5EkbqER0UmJBUbjyGYhvYmfy7YRl/X7jKQetbdfXRxYne6ZGxkO4PEDUpn97xRtVNYYR0
OD2en8XMgy372XtwYG5Ou+lMFCI1+/y1palyUhEdJc3Ab0AXVBDUdkqqTEzHfHJ4+/I8yLFVpVNd
vozwusaFabJ2yuClS6+eeSqIewpXJNQGe79q2UJp+gFjdbb2IK4yV8aO8/UypXNcz4nExuKaSPJQ
z5bZiduuziraS0H5bAdVN+/K8dn9u1mmmqxVkQa7IZ27I4fDLfQMxO0u2CVD+dJB9fYI4PuUk1IJ
+G5UK7AGrqysllbaSfQ1mgDyWiQzi4dSfg16RoH7vVuQsEywpCAqm7Vl6VVJs32r6J4BV+3Dr5Hz
5GuAMBv7vN/umDRKDA4I4XNAak24KRrBanYVrSfdmrUDf9txI3VEY4wHPYXZO2R5dr40+L3jiYbO
6SIOJ0JuIHhC9b4aw+ct+1PO39rbOWgsZa7JI75FI6vRUrjgfmH8/A2v4f3goehiBwkrd4Q4NWBt
nFg8Ef0QIw5fe4GBmGx61rzYpNfzW9ZE9bi3exnlLneLP5d3H3dKw7r8UTfKJf+2i/COgulLUVOo
kk4rP5DcVoKlNChUTGRoSMOmIyPsv7r7pc4RHJzj3NwbjNcQWJEiQtAt9ZGvi7x3WVkTOx0o+mk8
dHNdsadM4iSCVg4GtiGCVBUSd8NW32aO3fqqxfWFkD5gT+pm1V3KCXAiFmrgzthJG0KJ53eXtV3K
ZR+KXmlLx3yL1QpUS7kCsCtr+L7WyBuyGsAZfH113D5L+387pe1Ujh8C7vrbD1JqxYmlGl6MJeTh
xhY/ErPl6+OpXEqwVdwMNcoFwge2dwGU5q/DYyMha4mBeuVjwOzQ2pB5CpFXEq6/0mGeWeqAZoW/
+pkiVSRHqWDvCBjyZwukz2Jzb3zCYrCdqniannPY5vGOp3qD42UoRj7F/+lReLOJ2lT/ElQ4kFvM
Ad1IbmA1aC/vPqLoj4/2k86SfXdcYSqrwicXFzHOeS1i9HeXhBh0qNAgasmFqlLTly7bGa+BFO1P
SJ535psh4EKeXj/E71o+NFHElai6gLtZNKLpYl3/v3i9nbbZI0t4pMmQWeQGjaot5UdPrORBUvh7
/IQlcIjvuoOb/WPNvdY7kX8+iZVLtRaZGUkTQiRjYy0f2HDLUZ3pnc5hht7q67lmcT6Ip+rUgOpi
5gcHuvCWmOEA+PACeJ5QV4uxI9TPthtL+0ba9uCy5ALaj2NNB2gCmcHuufvbraslXdADuW0lhAMi
RVdejFleyPDmzlUMhuHepbVg0DzqgMvhA4PqpndoxYkHmtV1iu4eNac8k1IiD+XzBaVCZ92eaknJ
T++JS+nbGEzraq2ntAp23MJpsgkeaq9kO+LyWRo7a54/VYPynh9khjZ4PshrldgdVR84KPehPxGc
BqSPvvg2tc0eEVaW7PhUGhxOcQHph0UYqxsWV37lLHSxyQZ3kb2bQW6VJ39L0f1L00Fz75tQhQsf
rBw5cW7ma23Afr6rTVUuNDm8MGoXEZCIAgSISJkoC5ddLArQfYskywIvubwekXhLBhPFJ8sdL2C5
yS1Wa5SR+xY2SQE0gGazVLKbQFCiwpVdjuBykQrYg/5/OKkE+Uc4Uc324FbD00B0zjivq5y3o4rN
IDHR8EP569gcNzcnhbzTtg4Go3XW9s06tnmH5s08d9rBECMQDFs2CceVNqpBbvJXRhx48LQyoYcR
i5dM/Don6A6qVNIY+i3FM+qymtP6phTdHugg3L+6hJfkdkUa4QgztMKRLenM46tdtV9Qulmg/B/J
ednYw8XdMbKZZYRileVlMdzYdX33Us69VweMMp0LivzmMeT/KnbWkH+GIJfIqSw1HJfjkF+WFyKB
+wMZv/sgujbTmxOn/3xDdgV5PxVuLCTYV9bwDDo47RgIydpJQgOiwCsmYx6mQ4vh4ZfEDLUpj/au
vwwgienJyQnB4darh2YAuKvkcBI3sKhQbPrQBn+wiyU+1pimKRMWiYiZok59AUK8r88yRGOtQ3/s
MzbaNu8/2CqzqMVy8cAzy13mft20x11yFuBoapeas3HkEJInl0p+9yu7LWpIqJmnxDEqymv8ErK2
sC2fEqeGVg0N9YE3isAsqVdQ+j+LGHYrNbdIgD9CABpP6AAqsnIuvc/tZ2VUYBM++CJIboOW7Jt2
qVIdYxfVnvz7KPbMFvJ5iawIkvtyDmQwpqhnt3cTISb81xZkyJz954o/Z9chUmRpwrPQLHjwpD/C
IR+6g6vNA1yFpaQHIwTcre2dCZO5uU55IiPLyzSTzwE0e4OkW7RI1+NgcbrQjJWwnzAXyYvMnehg
ltrd3onDoePOzV6mDxf3vjmMInPdaDnwEAy68Gqj0GFkPYJUsdRiyir9dc8uLvvmT8pJLkYcr9gR
57GFamdNgrGj05BDyJD6L9k6VQfFp1PR9EDOazlPrIHe4zEQXRd5g6NkMelvALYzx5wF85AoVIT4
OaQjuX3uy6GdbabqEQpmY0Df6aeABf6wCiXUwx90lw68GIJUuQWVp3g6ZVwzkLxLefjRC/vKzlEg
r5REt4QTXxM0OhgLhWS0tsI4sDh5FK6HqoEMJHyLI3dXLYNgbM3q3Cm7zaOw7+uHFYHs1rR37Dq+
3Zp4/3+xM4wFHNtmu94XdFMsW2G/WspnZSRIHbDTAw3N27cYoyQFLdcgKB1tu3OCpXepjPdt5jD0
8PQ4AfNIveZbs9YUk9hMwmJU6UyCeA7CkhDGSAWia8PuRRG+jkbW2/aGUBBWQe1SoItlecLXNKe2
N0lD3jmAeiAqO0S3CKvXqRWRYcIAM4PHMgTXFcoYitALpK4riLJSkNbx8AOjcicqHnXcAjFvWdTY
GWLdnhpDoaxquFxXF3Vvoiar16AoKHRBPtFdvekyqJigdPdnkriZJw3f+rF6KzSu+KtavDbECf6X
FkgstFCIhbvI+mphx+RGa3NPODW8Ta8smukFpkXJ6VQDWPmW2PZNc+1uyeoZ8/R6KBEIPIynAiNg
EGZ4RONZGbTqwiV8eDnWPHbTNudMEGsPIlCTzY1cLsT36biB5NVmUFKxLc0ADGk87fuX7zeeEHny
QzifGesJwt0Zjtu7hX0nMwzMTEjGY/wTKkBpV72vCjmLcKd/aX5Dq5XqJD9fpjBmgV6V/slMQysC
7qO865AWT6OpF41cP5eHyrrjoGPIFz1qcIk6ec2mIJtPj+c57sb7n1Uqh4rgqwbtxLtJopbgVA22
O82JJo1Z5eFBq3s0QblyymeEcTiLxyJp1AWkILNGnjYaDBz8YuOOEMR32gdqoKnzjgB5LcyfUOlv
DKNzy6QxUST1iMMJx5dTD7gWHhkRJtpYT60AVYSmG61BulXJSHi2W8KHQydx3Is9gN7DBJnoQ4yC
Ym256ds7ZMxmxKzhJarCzziOWBdtg2HaUo+znJ8bIA4LRLY+7Te2gl6sKowsZ6B4UFUKtVYo1beQ
PH4vyoazWgJNC6yBC3+5PpQDSoFf0htsCPhMSPFtCJAxwA/Gscfh2N2H+KfA4n8RWn/B7WWt62Rb
iDCe/TbI4IsHYORVXlMM1X0BBc6OUePkojs3Sp2ILIdsL9T1I8vP7xq+/JRXzAXMIp5v9rLdKr40
CRhDmh6Hsow8/UyUDYXGmYEsmpD173cWKUrCvDWf0Dr6l9rKgAvbBBtAIV+9Bw/H/XLNrdFT9nq5
Xb4i3sR0TIeBcKbMmyZUqrKdK56j504D5/7BJ6z30FmSLocOxIucqPoUX/+cajHmgYAIArt2dzL1
N0Dog8S4JsqUfeNb4OzEp1YDTsoiFgXhciMVufwt/l+/fRik86twwosIIdaUZwiti6XuiF2Cw+1m
SrhKIxaNfQtQFqM6qPpIQ4doEBwpL9HBAMTDYzGQ4p9JCvZxYfi3IfTE5zy4cWeKCQPX/W/mx7VX
GF8XcEz/JLji5sMw+xONnzYumlWftalvLTwN2tHGaj5VwKj3MvAM3mYU3v9mGvGkmHf0u+bQLWjx
tRxBI8Z+TH5S2E7neat2mT+T9JKw9cdU2FsKPEQgvT9U9bsgFo3KGf+FJ19UPofzRQjim2l1iesv
obmDawBRe++AS6Ve0SQZdoKXADIFcXWpdkSZP5kk36zmy0ESMeDAYst/WjEJE+K8TdGMq9D0iMYS
xHEfTcYdimLGC5Fo+1ASKDxggbBR3lhToIlt4vp5YptGsce1RyLeAJ3du2YdSqencY9Sje6nk+za
fJFxtDASQImxqkCtz30kpZnoZf2+egoNeL8oq8y/8WQyIHPjenrpH8wvKhcY7nPYW4xKRarwd783
AoZ4Aa5KcmLwdOz0tPrVDaJttvHm+KSj36hCAf25eB5r9wy415EyAm7HImON/VDurIDXJZPU0GNW
rsoILRWxH5HDMQdtheSjkch/ElQo46h9VEp4Bl+a2TW5te/KWZTdQV5AlByIfR8zMLl+hwYfi7S5
G/ioUSKYXF2JDhCCSgoJhAJiL5mAaawk2LYD30Q5k35SVPdKHMVRoEJXquV9BSicuJkLP5CpzDHw
YJ/Z8qEt23sIDSrIK7vf3KoKbaznTg0s+qcKSFcWhOc8yc6oHmOe1PTQiPQKwy/e8UwcN5p9PiHJ
VsikeLiaZUdnQ/BWSuWYVFMEQm38xhEtzPlJfegzSJ1HtAjALDt0arfjpkO/d00fQDoFak39v0S6
22+2Ljj+SqG7iRElveRY+v7EXGta4uGn6otKbzwADixx/OlRuqWue4kmBiP7NQhkwzij7WWChEX6
Yct6sA9eVfi0ulywK7YtiVzCoTEUCW0E0lAXIAJa+FBPIOTEyKViP7vCAM0njsjyGJ3pxuG7rjqL
o6wAUMvGvPsmidcM4nJOyZpZuBF2tYxyRW4x7efG5kRhe1mqrJbrZYKggvojTJkPyJ/iimVhzdXx
yrDw5qoLc+UMtL4+ndtYycgigsp5grtLf4EPlljfgPg2VBeq0SXwr4rhw43K/5lYGDMniLjAc87J
3WN9ILipDLwvyR0hNy9ZIZz8R50E0hTJEKkcjeWoEyFCxN7u38DWxQSFOmPiSdtbCbIiwb/Gh3kZ
bgTS+5abO7m/ogP0KJT43zkex34qOBcwce2ckT1g5z58wcyrTnUpslABCBAjrmEHP1jcRbF4ZVsg
BJZtH5x3xahG/E8AaiImsi5z5FmkYpqS1OxCtb4yVNjovoAiUBSWOXu3lL+mMlcnaQ0/WQF2O5yp
usdFAVzvOc/nEFB+Gz7zcDssiNNAgKvK/Zed7jUlLuGWS092hT98WC82F+qPoqxK37OS2JFdm8MO
HZpbrh0ltei88WmFfX2idZHp/OTWRsUw5viX0QaeqXAKo5bFhE+7f6+/7Dj6dY/t1RzvcmmtxZ7q
oqdVHuOEnNhlQEFYSpHqknbXPlXVOzjw0lGZSsbZQFhgGYTQ+5wbEi/tTiIP11izxlVu5MNNvA3o
VOGH9/XPnIrCwzyJI+SgbLFj0BGXBQezFwa78+bgAOzLw2MGTXAHmyaNU279e3vYBY81JfeOqvSs
EOFwEDkw9wx+ODl5OKnIBrPdm3tz8SG3bQxjutYSRPohT78A+MSzcKUwFeCRM3wuQAiwXYT4JTwO
X9zIJC07qQMXo4N62yHVZF4fHftzZ3lkcu/AkYULhxxUwp13NaO0w/72uDH2f/97OUIlDliXjPTL
6uinq46SCE9HR1TBvOMUaeqktb1q8nBmxPnrEho98Zfj/8UxZwTZdYXcy1kTuZju5zPefyniGCVu
7HjGLSUlVHTAEg4SM+ZYs/cSKjUq8smkXoDCrT5dawj2A3bGDHjGBwTxCj9s3zEma1Oswohn7ENa
5SF7Gry1yb0FK38ZHDq1FZfLs1KvslwNAvnHbEdnuNrSRzyZA4DsMp8CjRm8wkBvmtvN0Y1rqnb6
xHtf/53Wu/kdLoIga/EesO4PqP+U9OI8sbAhcvccyDluqozVEJNIb/ftBrexGhJfa4s1XM4fWUCJ
SFGjMx9sWAQC88q+MKpRyNKEKvaEMBpduesbyS+/VTRqRJ+KHzrmHwutd6FpvM1SUVLOk7+yikI2
l4XDGe+zqN6ZhEOKS2hx1ndPiTYtKiOBsgXFDa5CQA8WK9YfgC7O37r3+HGel/xhE9jnyaYZ2OY6
9mJ4Itm2JSEh81o58nzdt1lAAW8j2cU1rrkG4xmv3dfzfIKPL21Dn/noaVaItWNZ2BqjO2es+K0b
loFa1bRq1HxQPDUPj6ie2KpvuJCgs8j3FiRmNIKKNnvkJUG8ihXrKUWSYa+sYHVxYksQByU1XYNQ
1auQ+Dop9BejIzCXVLemRXWsKHjw1CfDU5JQYATixNr3Uw8QZwl/qVEXDYbQG64NGbA460XbhNsh
TXkgkmPqX0ilf3f4LT+/KPM3iImDwObt/soisJ0ts6cBVLjbIURrKXWQ4bRddSVHcpWwjl9FQi+X
3brDJMFSRouoQXC9KZBaek87O/x2c0VuuO3GzXhu+bRXCSDbweLW/SqYxVEUGinL+OYhYxWiYS8T
tiSmE/co+NvGjisHdKAw0fcqbtIiVbHfvi+3YNcXb0eaLdEfEtuIJQDdFc3mhByp96QzV5slgV8E
V+9g9N1LaISYTva6mTO3HPAQde2LiSATujworFS/mwKkEEeag3SQ+ZHMGc4/wGTupp9Yn2tcN+/h
d15EcnnuEXKl/R2JO/8mGGiPVh1KJWOSKmXxr8zhMFFsyWvHrypJ/4P/e7BOqJTvFl9FLVih308k
poFEWoBHLB1rir7ekVWduhXNJo7qnlLVvPjSXs8biz3vXp7QZR1r9YuBEIfdTw/Yo65pU+UkUORT
so/4GSwGJP0=
`protect end_protected

