

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e2VQd/JkHeEe4mr54dnWM16g2399v0mhU+1ZT8oWFJUJCdyMu4+q7oH8u3QZmAK8Rcnxp+2SrcpO
m9pYEpjU5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e4k3IaAaNAlNFkvmIoO4qJK1gZoF/VExyr/L2EnpV2zV6AVGzYp83eEX/q7O167vsBLgWYGwRFsP
yi4sfYl5lIuJf2EmeuOEauZwESJuKd6uc1klxaADn7CdEBB8W/rBSaqjDoVCuWxTpK1As0yCX9BZ
RkI2Kfe6mL0Xs6sQpTo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IbtPpkhRONJmgAFUIssZ5lSlLGn92JCOk3a/5TU0b+nZGM9b2fJWwwoGbY/OL/gG3eCzPWC2mZ4Q
yQHVXagA0da67WaW3vnZMDAL5frakXXSrA2s87T1FAjqJLmQF7Unh7546PBsqL3OQpKa5tE2Qt9p
EVAvDXDTdLcKhvmEciakrtXwSTthowcA9uRLxUPk8f0EUO4CTfkvluf6ycg5PO6pxfumZFj/0WGs
vgTtbHeVNSCwdx/DPIPQrx/2AfRxSZujtPeD86jE5AaqkaHPmVodviYONlhtWin/aHIYEIBELmjP
OfgBpo4y7pdG2K9gwF+I76hLDXYgXkS1E3SJtA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jYNHOo/XTSvo0oBfqkgIM6041mVNycidzkShFA7DjL3O3k+3PIOaz1gxN4XAJeVyBTFZGUu9UNpb
lLYIK0sXIcMhzqD/csYXqYD72yk+XSADEYXGdJxFpJfGamCnDtSyBZIo7PBWUINe2Do8h7OVRMiK
aS7bCOSSci8hvDiZE80=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZHkoK3izETxxNJyR8GdmtFOEPHd8+4rIb//gPmmS/L1BfMiycMWs4JZ0IF56rYeBFqrbQeNtD9Va
BKnGrhYVPTrxcjX5+asuKlu46CBX/iIHEmzrKpr/LAUFIgJgUQFePcXNFNPZEAJsYZmhuSrzc2sY
05sJlmShgR0KVQTbBUWl7mt1DY93aBIhdhmiaHpULcmSxpAU6go9uAbU3jUM00ZMhYA25YYv6AEb
gg84k1+xXW4rmxbK8BWXOVrPImvNZoYgt8qi2fdGpgMvgaoBCq3Rxxbaiti+CXpWZdQ5NbjWArUp
y47h8RokwLA8qG0K8OF44wzHSSkCcalfq4pG0w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26336)
`protect data_block
Azs6F9n07IaRo1ImMunVJxOeU/+RMtyXzjIAbSQMfes53RNKxEPnvakzC7Q4u7T6ZdrE8HyP3CIM
muC8kesALsoJvQ9qODWZrC5GJDK3YiimZKYYUg3TB8cF2rKy+0lpBQBlOPd44kiSzCHC7jS1qXnm
KDXCdCvz1tX1HIodYbSWWSEqeai3Bp5WyKxDHp4ibS6AT8uZiFob2eYnLkwk66sSTMdPgc7eTx0Z
LbnhD/+PG0IJ8Kf0CBWqRcgRv7xpudd1+te1sOEvusJB4Cdb9TXWsYmhTnXg8LxueSFTMCsaNrjw
C8iu4m1C3L8/jMImtD1mrozQKqLH+7zkdLdnm14VtyNsJeFDlUYLY+pg1RAgNTKBFIzIAf7L9qkQ
jluwN+hlDSz4iE9aF1LqUedPEDTcTf/Of5QwzXIKSqmNr7AAHJI4dkZ4Y0BVhYHI6TGAlZy3ayG/
Ux+SI9RmqDyeQHZ6DEa+lKYUQljGFsYWhtuS4FMG637svALRnS5pd5CBmSQ0UVqVoa5i+pCahMwo
JR47VodRbtMRuzxx6e/01xOHR/1zoPhhqI9Ed/1UUrRUwCcJOIUp3ll4NEib7ndbaSFPatp16Loa
A70t9bLTBd491mBY8SuxGvGYTSS53iaXexjCVjCn6+9m+jeYc32arhyBRFVBzFOHkwLIX3wpriUO
69V6+VRodK7mNE310VojEPfvnHadi2vwIxtHG1OiRSQbwJechMfn/jun298Ea5NKxj2YRmbShyZz
XORl8PhKfhzvE6aWNHdSPzFAXCNW5dEZv/39CxGIZV8VM46+3V+KhYRz1orSKHBXO9KKBDpnRVei
6Vd/r2+0IGmUu0bOhzdPTmwbfTi5kfCs03yQN2eahUl/bqqX8dy4uQFwCVeBSYu9RfsDTNW6CQbS
M04xsSvdlO43iN8SZh7Xx4o6lQuEN47ApcJ/S3bFvXbKz7FBe3OtmbrUdLIHYxEO6VSGVDq7TU8j
IZmdt36snj6zAy25cR2bscAdhQuuRpbgC8Z5QEEtcYz8Lmc1GzW0uHUCskHkZa4iy1OuPisJTdoU
mIA7imAQPA0aHaexTZZerJkKTbGhFs3kMw1nk9IZGeVCqlZJuxTowpeL2Dkb34wEkNJeSCztOaoc
KZMxp3wn/mRbzZFL6jWBhqyOmVKDkfWXbAYcCjO3S7C/Dnx5yn2dKA4Kj6PN+Oyob9AnrnoeWwjw
vJTXUYWE85T3D7mZfDqYtmzbjCDbGs+ISw7WhsrpeEc1+/KVRGjn64ysc0sn/RIkcUQ/rcQS8aoM
cqdJWeKKXbp2IJcVDWRImefDEaOUtmA63fRjHFBMMRzWjIFnU7eUjjwjsqiqW/bfAu3lRlJgf8pt
VEqFua8QolPUkacn6bNBXt4ug8Ra54Fk+w9FrdNxdevqNIRIjjdWAZ3vCR9Y0HWcU68V7qpxhwCU
xJdEssD9nZZY+XXEXUBXlZ5HEiHKEKX2kACK+98o33MZtpvlJuH3VQvMxlTqYLmHSjnX49knJuKp
JW8/NfRRA4HOPR2nD6qkP1Deg6hFui1WbA3B6kBMk8vlFbKsDWu8+DM7B2S0CRaJ80KhgBWdc+BS
QD2rE5ThTKpGbSzV2ikxcct/Fg+G28O6bUHO3KZfOih9zkIM04egdmQs+cFzE/PRsfptWKEj5k5t
KrZniwuMjyH9VB5JSm4y1JQVxzHVABGs3twk6CtbNMH6CGizSqWLIFR8c8fIUBVpnuSsanFHTcF6
S+UwPi2Uy/LH5W2WeaVaGipaAP2tWfreLH6Ac/48jNL1f56lXh2vtKgvNcsb3E4v/t5IqalrwKAZ
kI4GKQzgbKp0rHiaps13nTiz8jKyPBoH7DFvxcYCQN7td/ta2aWyvGTOoeg4Ui8GqjGmO27ZhOFz
M0NUpgIRykvqcrCjmDogNAC/t3Hj4gTUUyeBAggJ8HSvlJvOjXM4RDVUYM+ZgnSSc5aU2j7f79Dr
sfG6boxvMCzBZjL2f7GLJi6MF0jhwVjkowR5VPzR27VoABWoz7F/QV5CMy9hHefBoeHdwvPkJupx
FLLJClDV8EYLEOkh6ssCGPBzADaazKo8YaB/Vn0VzG+T+3SAzD6UoaaKX4sCd8gUfhRbQTXih3Hy
hFHH1gkVLlXy0CI39miPVfq38hd2sxeN7lG84ybAY/1Xp8fT/vV7huj45ZHV3gQUSAqhHTqS+53w
fGMEyZD1it4EJp5Dp5akIsUX3gChxn/kkdmNQbASWjAUHvordl2b/rHr6SU7YMiw8eSsrSWwppG0
Fw3izdWjeviChbVXaC2Ctw1snxhCa5L7E0wZ1uQEEwEYxQFsfGe8RR95EECF+TvZFPpmzq5dkQOp
RiYyH5mRo6/d7e79FsooJ4e3Dc0/EexTkyXqxagVjazQiBkFKnRjpbHsO5ZJ4oq66LV9NouNZ3LU
rPMbKHHJFgGjJe+/iL9DgjpbfrBGI4l7qFBdntRr4CrYqLP4z9McRcBktnQPCv4WCZtrE47KismR
V0Le6ZOSHt+X+z8lSsAWvFWr4iW5yQK6NIlo5TkTdz4o33wxFA7AC5UPQHggmjTECZIckMenmxRC
qNcUKsIzec/dbVGT8ujpd5H3haSAeOGb0iSb+JCMpYLXqRaq9694nxEaVhBKzypwmSQrIOi1z6iT
0nOL7CKQdg0stvdwDLvz4qB6rETjU2WN0XEtcHcAYqYYGrY3l+VvEbindTonAD11T0E4Vjf8jUkb
H5hJNdj1T+K94+FfvhaIfnzl5i2+yz/C94yVSprSnYpKT88AeKPcTGCc0zFiod2QerZFxNiDPN+a
T4ccp1F8OAJm1Mfynz2hn79s0+Bq8XAV++NrGg18pFaOXjoPfXGZLkn1knIqSRfPtFw1c1ZEJcfL
dppPD9POFpe9RPBPUqTc5Rof8ooZwNcWMbwnS+GcfX16X0CnOofluUYPQf/BdKmWu7PVFreHNlvf
dJy10MUu52+ysSfNj+rH46OSXEnHFqYYdi+/yWCH8SWp1/veQFEwcQ8cC1P/yXuZ/pvbGQnzKfbc
M6/IXTvrVPVTNLxQx0xzgoDvIA3TOw9Vy2teZMDOWYOIJMhqCe3LcNiTA6FPmblxXeSQBUUaWgVO
JmLe1GW4apjknA0amb7TeR/FdBrm2hIq1NUi6fslg1dZE7G6o8L/SmHNrbjMi7+oq1pkDQFluxMS
SNcPOUx7rB7R2ALQ90paGSPQxAtnmdKNjz/IlsEEgs3iQrb48yxoSLabHiClIfIdHDynzspL20rB
jEkqdOT/+7drzHdlAzrJGqIb6sCauU9yjWjGzfZbt1D10u9Iui+1i7igF5kUuNxLewEmr9t0PvwW
E0wtXZAd19NDmT6AU3ClEcuwU4ZoHFTyI8eVHjuO2ccvXIxKiqiZ1Ocl2bedvQGPw7WcaZnioctu
yfttL/aUNa+sJUu4Hm7jmMTLSTbqsq7FWkGKmoThI94Nqcx4Yp5uBVm/NVHql6OMMOE1kvJq96/u
1qMxxfCfF6WbK7sr1O4jBulMoLRbvJlPe/r8Wk8DIhccKrLcB7ir3Vw/ysLl75Y87Q1qae+uEusC
ac90nf7yLhP4Po5Px1TdJuG5LfpjP+emT5RiwWBnO7Ubkp3cAhvFIYzCnGGasFh+pdi85pIsgUGn
YF/SuLayR6cQ4Xb5TbTsxUjmqBwM2Brh6bKZDkXnDlrIeaeqEay2BUIml5x3FBPMc2+peAYCyDDE
wkFCvJ2OWmD+YkWuOi6TN/3um6iX+9/aw1J4o8ZyGJGI0AK32BfZIUPFILOTjDbcCZomfhaEl44G
B4GoJi/xXhvkqsQU2VXsC5dQBiGiM1T4Z4XpEE69rWLA4XjHTYMWMzBm2B/Y5ZwyOLV28isAiIAD
TPzMYh4n/n6jY974EsIL1gxQRdhWYl5oqricFIhRyaU92sbag73keluhcBNKe5LitzduzD8CgGUr
ODKHLXAITCQIwpPD1sfswKF0bgtxiZyABIjLBa9WeDcxw3PfC9Zlfz5CngBZRzin17PrWhprH3Uj
t0U6XWoC/DU7JXPCDaLtzv2Nlwir9V/5sjaRus3+M3Uj1InYMAgvQzfW7ASOQF+qBw1AHCEErFSR
/rui62XYMOXrarl6ZVvahjw5AMCxi3cPRHo8CeE1W+VglTGeWIM7/Lyox2bLcgSn652iGhiuFL1I
f/GzreyCXKFk2i0wS1PI9kOrDS9SWuj5K+puoMXk+vEtTKipvFciHuWcoqh+fgqrP+tqB5a2FOvf
kCvs/h/Pc+8mv7JZIxhUeU239nVbT/DdI2+DWiFA1dNjWHb+KtFAGUxylCqSn7AelGlKG1Qa872r
Y+n2d1WFRqdTjbizDyrc0SAxNISNKuJu/EeqNNfjMPnKOgmwRwyChulxZW4YEcFSw+r1zdInQwbV
RpgurLtZghX7z4WMGNWfGoBXKdoomhq6nfiuhQJBGcP/pNuKEgIcjAQx1/ZLV3+ym0iDMOxLCFQ7
PbpQ+UpF+vsw8qA9O2snx91vue9Zz2tReipwBI3sJbdxeaAyaw24yquZitYJLb/+EnajPmrfcjgn
33ukw4/VuIoVRjOSns/LG9nbyWiu2r+G3ENpYhjGGnR58m6GpSnUaS+hz/yS5+OwwJdFjow2L5yK
zG8m7rve9EctIbri4zbwo5QMfSOq1XVQIiEXSXsY7XTRQaAbkCBzN6e2WM2JygdQ9Di4cpaRzwgs
2J2KYKysQrHoG388Z3lnNChwwR52wJ1NmBDlgYvTBP0aRo0vVqd4Adl69ov/gAJ00DrMYH2E+wz0
nh9a5xkF6IA6iJRP8U8TK6e+Kw9iiEHXZIzMjElkWQ737NAYFZ/6B7NhgrpFllB0pNT45pnTGGGG
Ctm6tIsuEQsTZmMYv3WcFv1Zisfj4eO7OxJYu/3ImBnXXgHOLdijQShfdEuYKjn6+oQQf6xp7eaf
iNrdM+Gwhwf2Ym4pNCzbTxPxhWM1Q3nbfSMJvLjRyDM6gt42Qbo+/82moFSKXPjjBhQAD9aAjKZQ
qi01nb6ZuvRt2FWZvL4w4HdGloa6kpWPjtzy20H7057I+hkruW+M0kaXp3FxFtLl+PD5WLlu1vO+
LXGMPjlW2edZaqhqcgTO8bNQUZErux6Usr8474jwt+t6rM3V3aUOjuw9n1cN/tMQce0v/yxI9Al/
yfSU2V0v+lNRXaf7exE1bYPlqhPFiR3mBX4c9QxXXcVIJKwPRynBoifLCDg4KXyhdpvfP/BJGkhn
DvOs4Qwgm9fyRHmbn4D1pc7PghaoIRGDF3sokCN3WhtokakhnKQFLwQbFNw2XxAa3BVxUpCBPcGl
NOUvLJ3S0cth1RsESLCkRVu56C652v3W4K8BQXTaSTlUfK78qxj+DZ2YIGo9kEXohz6AXj4oGN51
TAraiRMDKy6VJ/tWg9E/8tVtwA1JVJl6s0xg+2sXWCzDbgq3zUftkkyekqNZ+ct1LiYdS50L/SR5
uOLvCHl/B7Du8aH65kyy45538waWDyZwArCnFZrbPOBLgOUdPlD2myY9pFZLnSlqTTXSoAWLlfH1
QifvQm6bAJ4fRFfc08LV0eMgXTVA3KAl22VpMDraYQTsNP3lDZgeMcMJ8+gWAB6SKA8VKKXidlbz
lCUuP61T4V+alvlBDYzr+M6LrIHIF6eY59rjkgJw6YZAo0z9BdBdW9B/gvRh9CfXRXYDVTprJteD
pXS7q+LM3j0Aw7HgAF3yaE5HIShXt98i/FG6ro/82Wq6TqK9AhCOZsl6Hb+m0Rjdj75UNJOmBqLu
A85GmsgST5cHLrGJ62m8CXzfIFlmTi7wnsX1AplKvEjdcCahHZgTsLI3uHP0GpRPREh4Alls32ls
topQoyWe+KHarp8my70tfmNRqRjl68TaXSvxs1aqwP9XOoku5dVbIIudHkZ0z7TmgBiAYVQsj4qm
1rli1roacMgc6//uedAW+s9pAxNe784Pfd4W9/o95/GhYYhrMTGKnmDw7H6k2HfiDfDnVg7HlQWc
fh5pAnO24ZxWdvtKIdCSYpSp7ozgqUr5cojAOj5Y1zTpTiiDtANvjOvs3sYqhN3D0jXRc9INKnjC
+LoN5b3THyLkVC71HPMw85zjAw7GNTo028ijIVJOqJF3CcEUz9kaWHpPGt1urJUjvEQt/YrT3Phj
/X3RMsSKqjCHmLbQxQ8KlFLtOmSd8TJa7EeQQKjtHZLAcWDAIo7ivx0BHve0SpElSFi0MNQbncs3
i9S7zLOubN+a9xb4oMPChOIxcO1hkytNmDmsBqpvILMIR/si8/G2p690ZceTUHrjUP51uvaRgn+d
9iXFHtHNeWVl93Tqb9/hPfZMZViiYLmNeImOPaWLsOq1RCBAXYiApzgOcWCqxLQJotwgmVBkv5oT
j1JqM6Z0pU9sn5oCfBNgxVQ9pyugnu+XdeF0ZAKj7IgZQoNI/+1iCwfytQlsklbPkpK9mJ2zh0JH
j2ypd4sKiZKAy9IFWzar/qDMvwY46Sl9nDXNcPK6VnMVgToV7xcMHfzizTZIHhP//yVAi0SzHETy
cZJFFiX4t6uhRA4bh9iAJA22jQy/Nm8emUgkSd4t/MvRfoTeQri6187HZRi9Aa9CmACKtMESmRAp
rmJwYg5M2IZZP4S1Uxt1H3d0wFhhMWdSlwR7RjouxffyQBUR1MVm/MHF06hs/wUpE1rMov4Olk3L
VN0ZSMed3OJHNKsvDbBD1phvP8fb2t/jXt9Y6OPHYo6MbvxWJK+xnMU9wgN4oEGqxbHowEs8Rlfd
5X3dIcUSjzD6Q7kwWnxBxz3OpWT4QN59Krwy4XOfIZNE/AI3CrCgPMKNscT4CeJDgXusJY6uh/8K
5sgT10aMEJ67gd8J6Nj7IDHF0yWiBEHC9r9dByOt2QV1/UH8Um39Y6hT4r4ARwidPugwBZ4Cd0j+
zLtUMmrjnPYZhoKXtcmrrEfRjrLftCP34bKRz71ZsmzU9zSr0AhkS2HkNnGN+LU1tSdz4T+4Hj6/
qpGBT/JWT+rbg/RjWPgrhaGFEOxMr8wMrCL8QghvaG0gSYfaJ3p2Ir99rF1uLS8I3JnA+lCjwDXk
S8OHdWcJ4XvhlOKOH3rNaataM6fnjP9TXzB1Ma52DoVZb5VJNHcEKRm5GpWp3Zsaml4AnHW138gu
jy9cTr7BLTL0n/2gj8P8OgKKXR5ALIzCxmt7cTq5MgNlOPC0wqbWPkOVTkaf0qxLbf4LZMfuXB+5
STG06GwMtO3DPbdDJIaxAeZzrFVDkBd+IKH80diIkwKCmUO2k/QhuVIAJsJ/aEBM6Jv9VsuN8xqV
AUM3ccIaY8RKYSKTkhZ/2URxrdXMBvn14K+qpsvq+GH/yPIfkoRNTuMMLjxoRfrBf3D6BUaptOC7
9eXp7uhYjWmjnrt3mk7MEtv0NJt2rFbi8owTdB8D2SavtQgOtvTFNIV4hFdICJKSm9Kizs0geY9X
Y/oa5T0SIIbHpokQ3AVnCsggYaxM0/QG414fFZC1YZIcA+dbFWRR+f9yZyidqIVE80FgsnHI9jXn
kGcNAfCFk9/npEZlJNxUZVXGgofgSltmiHpNR5iX858/H1eboyh0aSHHbrDgIc2I5dZdqjdcS9Ea
HrGbaBvOAA49sk6BHKVfheJWcVmJwFVKGh9gB72fqn+gXdMEwdYP9CBm8UmT9aTao3eaHd0NL23u
GVRNBnLBqUb2yvRaRg9n/PYkBKBGriIR1g7J5FS1EhFRcG7SzLNgSWc1BM5eScTrxRVYNtPsMnna
OVi5SqUqIJWvqxmd8ey3WnS8aAkDxLEmUd/5h+cCFQZ6k8qdiR0bDC/FbFawhcJ01xiz6zCwMV8e
ARYMV/AyrNNqRURCc/d88fPl58iS+GSs9V1d+A6kga9F/2A2jWXgmrftNurc0eQfIt1agJN8dkLu
twO/9RDf+G13Cs4MZbt4alkRaEdl1D7DcddM/Z02PaWu9JDLtB+bUujo6l+8hI5TYtE8x3SWse0K
CUIp+crhgFGfa+VAIdVDYfV4zpDgRGFH7vxiQ0SAWeAwyi9qnvCEogzoj5EtBPe3ol+wecFrh5rw
KUmbBe/dkyajxZGW4S1zBSF1s2pz+QL4Ia7Wp2TgOuYUV/SatdJNjTkJhsjjRB9QrREPVOH4Zdho
xHASpIz7ZLV07Fy42Ae03hOwkZEkAFVDOZwNitNLxigcl19WQrTERrLu2LsiZK/BTzow46wT1cS1
AagPFiI2P2zu8sjGDh68R8Rzcj2FvgDqDXnM6w8VoGs+HiSDHyN2uDLYsMkinYBLIVJWgSYOaupF
qwCvxRD+op9czbpxRuEox1fRmJSXIp8SUt5M86WjHOZsWWgNR75gSFbbuwQJ8P2ORc6H9Prxd1Mq
tCYE4kq3ir30Hcymjuq2vTvIVGIQQG/KO5+Tne+fB9rz1fDebG77CRweYj5vbJBJpPcaqQBr0GHI
qRzWKDMNNheOqG5haoDjS/t0ACsTq4g+3AKaZI3RytXCuVXIQRNMaC2L7azB1st3CranfmZA9/ig
2sB7OlGmKevQlJyY8c/brnUBg8Grkvfd0HIRWXmXdc0vk1jqBQ6pxCObXDW0PWBACzOWHYa8z2ws
EUSZXcwUOXUnS/FwVWE5xyvM61l6N3Hy4uROf75CN5hMyYxHVA8/O7b/KoZIrCeoR2B/c5aMUMKl
8OEcdy7q3KbFGHgcfEDd/YeBYa6GOpSo1FBqCMo6VuqUU+rd8eQ8p63k1TatxsAnny5PVyA9wjEx
I8qAL70EexPCd6pHvr6X+UrAXjFverx4avLWZrz0GmxeUjCtg+0SD+eiDmyYNi6btu/Inhif/qgK
+qT8vseDRD/5L5qraq8FWzdOgTfoa/3YfPmdMrz5OY/TfMXqKpFon6N4iqfNFe05PzaYXhPxlNCV
UboKif+3uCa+2dShEIc0oSev01F6FwvW7iVjXVT3D0WU59HqIkSm4x/2t6ABKGSCJzrA4xM6vS8B
9YWeW1GMU1hDfPCJ/d98gbU3p3A85uOHMIQIAy9STB9J9+soF471g2TsskR1kKhNXl1TJxVjcABt
WlFYv+CWm763sKvL/PJowUiJrFKdjR+LVugk4l36ihsWB6T1K7qwahfKNAh7C2lSfz2tZ3ur84fM
dzF6x60SV35gIvoav5KjLRCpJRCCBTfPMZDx1W4hXtdAsk3l7hZKE5QZ1T/fVm1vUI178vwLC6Z2
RQ4VusnG+QyNnVvCoWD+G3IAVraiZ7IVDv1a9zS4X9wb3ZBHBr+yKw0VbjDjjJLTsLhjNMNgGi/r
W3yJI2U5CA/Qtd88I5qU8yhMGGsrFXPBWJFeBPXF6toNqrhpnlTk4MYD7VI3j95WlEsGp7LOGoWr
bpIm/ISgTI23foSJL3wc56mP/RYem4NOdqEjbNXoq9s9s19QyaQT5xCMGdKrzPH7V0wZx1rDAqfy
sAKESxBrTDz4PLb7V4nakPxEgWdPIoZRTyGJl1f9defcfCY4gNDYXhT2u6TBA1F5+SY2/LaSws+G
/12wLD8p4S7+r1ebFmrzIxmg/ITVlA8QUrUk6VnkXXyX/RWmTrPxsxGMk8AoqBjzZWjcvv+a9w+8
hEk9fVw2sbp2DHadW7CYohH+LKVodmvVjfyUElOxzl6hZhWxSnU6Jw0qzaDyVQGQKCBHznCqBPos
IK+nIDcTbHBUnS5ax7ucLG+fv1m6q764WJ9UooNf6GnR34WvsvB01t/VVniUlUMbFadasP5WKmGQ
MippRQIYEI4ytND9ruEMqyV+0Wjv/FzCtiDBZIOT9pRRFVuJhUDOBViFEdhd3gW/lhC91qvfI4R+
IXbFk1b2BTD7pLsKsOBDff1ZaNuX45LZMw1Lcv8DTsQlqlmDalCyOkn8X2OuEwgdfrDcEtFlI7LC
/hulNZAd7QjTiK+5K3qCH52MkbekASXOw/fL3kYwPxAII5+WV9oedoibmhjCKpFb9lEMM+GaogXZ
sR37ZghxhAu7sCHSIgpy3SKwqnVbu6Us8Fn2W4vA7MFzNx85jxpyq8zvIDhiF3u7ez4AygcedTFq
fnceUOCAfdcfSMreYD6NtUyI5r6xMt9Jy0nEPIKecSh6GdOOPtQCAmaGOFPv7+sGLlMYv2i/rt9o
vaFNGUs8OA+HtFOTRdCPS+M+jHeLfARDyjoRPgXv6vnA4CUiUP/YxYETyUul4lu0RUd3sxtIobDG
FVXoXuXqMRbAclwadOKpxBFYE2ZdLZEboI3p6nr4dAN1Txa44bSiYkkCL/Q7PwCowbUkrsxPUmo1
RIXtKd++unyDPuynpyMQmrEjvyHyJgs/Z3n/t7XBxlzK2kZsdUtxoc3hp/3Dyf6199jJ+/V06bnj
Pbu5yuLFgXQuR9ZoSs9AIqn2fc07JwzZrVhQSMo0V6aGR1TraSVVF1WfQXzGzfitrB5aUhkrHgcx
liVVFAbI88IokNKdBMZBOxQLD1V6I/JYTQReTEqOwLdarzrmlgvW7peBep+1KDzrhCU7wv4gT8kf
2zZBtiROL27+pq5LPhxnPui3dQPzXQHsC0+oNq8fsbGYAlwqeA9uma0pSqe0q/qs63qq7PayHlgv
S66XR1D5LdLhD0K++ONHuBs7NUSE7AHMU429W4Ni5WXVJ2jgJjTQVFLIx9sEYZa/e4SC6FEr7GaM
DNjKoHEiZYrW6eewGS++G8oYEnwXsrke4720lkkB/G5k0SBYe8jbtWyN90eVTRyXu1llm5ArlwM+
FOLERuPE6L6fH5wVCS9wD9z0FrZgnodn5VNKwuGb5uHdWxVGFP2KWDtPR3wX+A7G/cLfwOGRfSkk
4x0et6nUewhZV0d6DXpkhig9CMD1f5TzVjeTCvYCNQ9+rQLL9aabYDlIkxN5hGmMV8CQmqJvND/x
4NiflFaol9bKfUI4O9nP4TP8KHvfmJYxQDX4+FJeOVBBpWvddURxV2vCvS6Hqlo1sCdmmMLe/YsP
MjhHa8eATuTgFMiPJtHxvYdtKA12bKQzq4i2zrFVTz4zl0VUicKJzdK1z6QhllSR6bszaKV9lWt9
uVwSotHCYB2c7FgER1RBA2J3FtOA/GWR7HkqB4So9OMQG7pJpu0IJRqdbSmKRjXJMKhrPEva0kDn
brVbJEc3dvCH2MIdiE+9taYJ1GyoHW/t2bCU/WKDCsE1yd4UtlYmYEw922MoAI6xnH3zBx3YbN9i
vfrDJzP9HdEh4MkEapXnwL7erRIGWcQTtpif9ZFPS4PMUs+6D/5uQascck4mLsRqjkhatk3krzN0
4EQNaOJxefUpzQjwGcRtkR91pnQ1v21dj0quhidWg1242/XxzRBJMWbuKXCK7qYuOubwWo0D63SH
gWRzCQ2paRjx6HwLfbUvtrL82T/ILADPDZiDtuJHpAfxOGo5SscLD8qj1nuOSj9g8MifqBgndtKA
B1XczbQ+HfxjkvPrPsvGm+dZRtRhcC4+kJQa3hH6juO5IWd3c03uxitdtr2P54cumvu4zHwsG40j
mUvpC1lbWA7HDc/12U0Cf9yasx6m7ekBeugRzz77p+B6zH0mgayeAyDTpPzz8k7Tt1V9UKIyQVA9
4PHN3ERP8cNHn/bAeSQlzTbCCUOTS//UVoq3KHkYBgLi4n3Vmyzrbvt1OOz9y8hFonutENYPkhgd
pKgQ6SAyC7mwZNalpbDpCVuFeBBXMyz6s9nBWGK0pNsAqUsSknjcGbn9quiKBpXSDYUpjxhe9LYv
wS8ZUZZz94WHkzCCYvxwLgeOq1EWDE7itA/rseyG6eGX59jS+yUXq8rFIZofMwCa2qeN31uRZuwN
XbidkAlA6HOXQm4vB1Z0rGWz53pPkq9TboyLyiiEUXL3QHmVU/C71dhXJQhN2em8DN2sEsruw52U
2jIqkyPPzoFYGmecSunfHhS+TAVjRNJYGNz5V5Cn4Rt3RjyMNOuD577nolYXjv5mExloQ7qEL80E
VMI6Hl+alHiHh8PhjtIxGBxyQRyr+X2u+Zpukkw8t23SOG72RW/Lnl+YPnzGE/F3cEujMaEtFkiM
DNeRL5Eprp1rT2+BYdRPMyfcXZ3rLWTz+3t3k2ETTpKOnxNJuxZpIPHIIv+WA2B2M+CUQQ81PWFB
yKdbVc6PpD8ftW65y7iO+IzOgLzozZ2otj9bXKQUKFuUcpsT1HhIurxTYbyx8TsgTlGS1B95oJrz
WozVIkjxOs+m9GZvqMNSKolAW6DPbJ7vXXKF3qdn1EKRUn1uI7QcoxMfYdUw3r90zDNqOfqdID3b
1yTY6lrA6j3IE8h/yMJXq/YVcqR2QwsQ2scRmHO9zbt9cWW8U+F9Qr4acX19i7CPr4GsvLjNIuy6
eCYiOnx+d6m2guQ/oFZL/MTW0oKifV5FhNFMwFKRnz371P8jIrw1RzuDpJhozS5miOcj2QwhU/rh
QOSqg3qKDJd5oxfd8V0KklY+8kx1z2QSa3NPwa1PrpIwf3fZGH8gobfzmjeoSZygAR2FxeQtBfyy
FE+VhbIAohWZ9l5Ep04ModOnRN1xWOMHbTloNbGry2KoEMNG1/zCp7Cu714havjFgakVdhuDNH4u
khQULk9YiBwBp+Q/BbvywF3iV4j1MFt+xPyylHX44vEeg6o0mAszxaPwFLzQ+lGc2+m4ZoqBq/Di
D6+O25tk1CWONTykUcki9Ry6MrhJJwZn+hjo2D7XwsgAdl/B65+SOfrRKCyeSRTiuDtf1LUtiQ7n
yZltnmGxZF+XFu1sdiDf57+h0542yLRdZXdQMZmZtxDQNRB/ZNGq1mRIn+lQZJk9Kgu1rSDl3P+u
8MU6voeuXOTNq594yZGwCCcMrkwYbPmnIEoWHo2Jv+8K1jQ6TqXVhNXnYjlnrhwFgTQbCeytxn10
JWFRMpCR12y9ZRLxbvvSKfNqd6AsDnfS5h/katQOBeNY85lDhsJ/FWaPVcyAsEgOqsZk6dnt1blt
UX4WtJMdsFIVwodB018oLa4LGLthLhwdsXkCW86Y4U2NZvYUekeqjAe3NgCbfOS+H5ZUxGqQ9/Wu
4t3iK8Sw/UpOJYcVHPFLaDDDdUBxYg0IgR01mnf6LC5ywlxlhQzFCqYM8SQ3/uxRSW2/Ee+/P0uc
Scf1HwNh9d/7ndasgkTUEN9U5JJZABiEdp9+w2uZdVlXdkax1GqvKj8uF3+46WGWc6uEMuD8G+iR
LRgqt0VbJK9i61uDmAwBlosAbEIiN5rjNrxrTZYsMTmbblWznSuI49sD5WlUDWpkSwFAJfqOoZgn
scpiXA7C2wITUY1Qk+gUl1fco9rfEclIkZx0fGFOIcouMtFCuVF7IM7eepTkm8ubdNESUf5/LNOV
xRWdmMwQqtdg96gkChNtfdKCO2HnTWnrZc4RvDyKeH3nmw+tVelDaFdTAiG8J5f5aWKhThy1Mubo
3H4P8k65nP9rYYSlc62vdLkn1dJfCq9Yz3YHYkTZdYUnflRBv0wfiql69/akdAAWofDkT5yBrNsf
lsnsPjLA5GswueLRI+psj6e53PEOF9i9rny+QWmmlbZQyqHvZ0cssF8zH9J/30HNk7lBQzG9MK6X
9vqOvtZTFJB1J9WhqZ4KsoLDB4JNrHtDV4AGb/Cv7+CEs5Jt1dtnI888VOzmXQm6Y/rHfZY8XsDX
6LC/w7IDi1pVQXs/r/C4pNAEEgTkhtWKIrnk7ETz9/zhmG3SeJkhElPjh2Zp9lZW4nSMe57E0u9t
5US2i5n28VLQrUR3OR24c9rOfOUPV60VilGbuGOTOsnp6vnDTY60mHm0jr0xL7jN1K80D3xxeoiE
loxh552TiwGCEaSa+fH67NzAEdysgKa7WmYeoB8bmXdQjVCQ0TzOK23+RmXhy3+5iOxYrQVd5DN+
gI+89AJroWriKTR6S4Gi71Qgjph39ts8vYlfftlIYnPb+wybxMDNLOBYX01aCEm6CXJ4ENTnkRRO
gzGdFzHunHBLavO+p+N4PjAUK7dSF+O6pgs3OOKdI9mvm/pMnTqwWhH9zLLHjn9nLm+OiDCAlcTC
JbnXf9vwgMbxkJkT8fRzyCKC/HYoMA+xHw9E1oXSqrEZYDyGEPt4WyFktBhfh36im+/R1NsAcZZu
TDhi+S2o+8bxGCPzHjfNPYF+b2Mgf2UFVuMpjCIRJ0TPeC1R8Swx9akEMkUJTpHd6X7U2P+ZDvfO
qmNX5FkwSmOG5joebNgx5pHMmCLA6hj5Oyc7znMPPSHJ4wuZpDg+POg08jxGTz1gBrQ/HG58eWlu
jENkObTN1Ba24geIWsHOCWP6v6bYOwgkhKbBcoo7dugY1VkszoW4vxPNRF0EX64zeZwyF6fYPPkJ
3jmt3qssiL+I6utrEq6VesXaLokqZdKNwCUyeO3GWE5Ou5nkPlvm/+NY63BxPS/zqLJ2VEkXIagO
Ng4C+mD8nHi10Et2nn6UMYV5t6lqYylod1oj0KpBbFaA0QaxRAYjLKswOqICodVFHfxIW9Zw1B/j
ECGXqabCBP9id4rsT+Xq/9aklgitqruCLyaItN3IJ8+rxPqcarqIg8SZQ/jexF8Cz+tYiAnP+uji
T5TSKeQmK48q4LaYlzDR0fWRgZUVIDLjSTJm1FECvV4jorvGFzNriiatqDSepsZNUwbBvHA9+/yS
Kl9W42XG4zLyPmyld41aMM5uBLzj2svbvM8iXAnpGlq2QrZUHpvFhje61YxF1yLdHPdUfqgWhVjS
dZAz1vIdaZAcsgjYDQS2XZLUdlSiYVARKCaIqqvwthPpSpWWJMicKLM8Tyfnu2cCYzuVsWhXOFqh
nUtR/czf4D9nVD/t7eBc7tvvETwfzGbwNnF3bkF0TOzIWkn9YAWqVUsqxHZMX6WQYlNtImfURL35
jJQl0/IhqXbynGDZGK2/M2UxCGuk7v/6np7qnNZlwvK6ikdps61sAdwJV+i0r44Tut7o75rQi7LQ
iHrASckGPDNNQY2VxA34quhPCO9r1i6bmNWp43cCZlUNzGAqburELHMFStR+HQQxLyeXGgKKJ4q9
h8ib0pvLMMEO0eqZMgRH+QJXwxaK5o2W0ioNs6bPDaE5LZGJzopJ01dbM5h/hUZSdTS4sM0rlsRu
/5s4cfshUjjtUbTSU9RLST7YzQ8ya7yeQi6mLOTBwmbFN34ESa3f9dkfh6wVejwpF2LMLBs2Z6RA
8PZEtaMGbE2BqYo+IOes9aE7k/jxWLgw029492jva16AVnxCsggCuVWyZ75qzvsF9TsmisB2+qdh
asHoGHU6+dOJvdnBq73gkGA4stHCVQSf/3P8jc0DiI4hD9FIEFZP4QwY+oFhVJBQ6oOx2x7AlsdS
RDOjZnRwa5BTipBaAt4SH11uIsnVGLXUN1TGa2y2Ac+UbknEj1N1IpRvCQMECp7VZcyAoHICqIoO
5jT/s5ScutUhRWnKrdxrA0vO1enaAFAbn7HoaachsTwWfnFvToZjDWj02qB3omLFy+PrkwkQRfNL
tHisJp8N0tnJmefRanrU5yiNw8wjSVK2wGgA0ns0M3/ZOelHsqgoxMzzQgtme9LXoO7es4HeyFZS
CaEDpHcFQRXlspcPa2zfTmxJBS5Cwp1R6VFqeFXznbsUxwsj63kkGDLlUNVCNQPLxys9Z9k55QI7
j7EBvQmuApF0dTP7D2TD7w1xlb0hgqu0J/EFwQ7iD2IQ4T+3ElHYwuHIFWUYxdAGgLq8OeUYZzGw
6yqq4aptC+M+e2QrGY8KeUDD+oZ5x/FjINx6s6Agc9dVPITJLwdm0VTdUHPoqZH6i3C0nEuhtFR4
g4fyr0/0j7kTb8RxolI5w1dIJ6jf/UCYBurzeIjhQeGAXofWZhBI1nPMQn9QDIFL1nLXdC0TQB93
8LV5yRlso6aNN6szA9nVndK7jqc8jBxIC+8Xfx1fS35s90oZLNA1Z5itHwo41lqd4ha7ZxS7WmHO
GwfFCV1Py2hGObt4yjRRbO/WR7rTmkAKdQu6Gz55SOaP4zC46FZFzEQVMobmmFwfyuMLAYyrejk1
eUc1HLubSZoUykMizvN0NFQ+P11E2Q9q71cuUiu335yK9CLLTxFNS5teY//50rhkhfiTUBhyZ3Vt
3AVBnoCqi8t+wThtIMmw0oWbUA+ue+TpD0iri6ZaIzvjYkGCYTt23ac6ssucKvbilqUIfG4lOiKk
du17qJ4ajNqZIeluxSHO8zpg88+XilYFAIYR4v+3BbPlJxaV6uHgPCSM2PRcT/GM5h6N3n92rfkX
mxOcnVZfOXXKiNDvItXEUvd58m/2sV8pSsThsms6c4ZT5P+gQc3tyqTX1RWtd/t320vpNLoNe3za
DAnd5Vg5UdKInKzVJsjaPqBYv5/MlomHLe5PtVYz3L8nved0znp8ehD1c7X2/s1Np71Xyg8D8wOF
khqmhAnCK5IL9C/04R6Satsr+UiQ5T8Tx8+clKwi7SEAMHSsDZAvEktZAg29jYQRpawzgfVenXjO
rAffqgmRAiXS7Ise4sb8OMOUfTQbG2m3UnSD4IoOK9eFREjEGqd7bgsYniJFrzEWnZNI/x/ebG5Z
LnS9ggmqqInGj1X/MgJt6MKItHfpFoamsHVlc/7ZkCuoWrpIAESmvL8U+hAGk/UnK3B1YY40d71J
4coHXgerIqQbMMSDpZG3dYHzXw8Tetxu3oQEJeYT7XQdTrF/pAKzvL+qi81cyOyfTFO/U/euiHPn
pW0AE2SzvpjcblHUHFEEMlVDwmywnWPqSz6sV40sb/6bp9ZuzB/fQsGD3WlwMggYlioUCW/9R/wy
Iy5CXcw6VW9CSBtj81MhNaJZ+z2k2njBHvB2rtntWPpEN2jUVBLHf2OJreYRliAN+QuSfTDoZPMh
sv01fsGDAVhQwXr1qIRim1rVL7AzbrxtI7hRnJ27xIVKQ6jT3wuim7jqVP3C1eSaiQPgIhBqQ/iF
999OykITj9eCDPTDvL+1p6iEnRvGVcVVDgm+2UGherSSMrKT47ZK4xEVAG4T8nhsyjSrpmMfh1N4
dI1IlrErPr8YXLiDzynmpURqVgnHe8GBtCtO/vwYY2m8S64Zwtrjo/ENsYy8ZAkSqDltf3mSD0sO
ERBa4Bf/PZBsd7Wg3m7Vh5n80Cr4SFVoEC82n0ZuDw2ktvW+msPhSwDcNLeiVitvtcp7OYyW/yMK
49X8ce0S/YagflenC3PENe0qUy6Qj77mMbZRKPuAvkxqG6XmGTOAOPtgf67Rn3PXOxuDpPe946MV
I9EqEWQJSnPoq+osx+I/zAGA16v8LdRe6SZFK7K0jMHeC32OfY2XKMjIURsNqkDchukOvwWLdIYZ
e798pk7A02/MV3etmjhSWcGKgwH7IQ5o/XgvBLFf5dbPdMclkbT2auwzrbvcJ/MyXHAvDcRHLH4i
EqHbjCKjKZ70FwdvXunEqwWSHuqT/Nsq2GdQwj5kxrzhJqAU+voQ9oplHJ8qasJblLNk3C2RP63V
uEsRuI1GLxbdOh/Awldu7CFgoC4xgLNL3aGlsMLfWLFOvb13tDdgzklz9z5iW/pti2n/P74GC/aA
kxoZP24c3nc4ZcjUGaGXVCrZNyoJuTVfcJ3nK366+FmDE+OPuP3PkJOsqAl+H/aaANqEcqc46Ufa
O4u5TbXXucfh34aha7EelMJAym32uA3qiIR5smBELEXiynp9rXOcosEFHQwq0LQv+GP4E1xSr17h
lv57XUi0uSg48cqrLqjm8a68yth6J6Q5z9a2KaAr/RXTlksg7zU7figvgJ8g7VPieBvidO2Mie3b
7/Q/ozdmf96EUC97noAYMBuzvXE49e0F35TEqjbiTAmkgn/tRCA4b5DxPK56GxwWfBnN/VjYi2Gp
x95qtqyI4BPmDljYIcuubnt/qIEGlPBOeIZVSUlhRgsdeBWgV+nFKiwpqTeIoeXTPNzkN6sSgOB7
MZtX+eSQw4oIQAXZxtSyO9cs0AXCN2eZVKGkmChnrSg8DLyiMldiJV+TjUjifN0M+ZhVIslzjdae
ddu8mQAoKZZkiLA2ZEy3QtNyZRlnGZPMJLpuTR33zwHRQgzrvcKRzegvIY0KQJhV/KB7jJSIefrw
7FZ3XzQyKI1TGjukcsntKtOL8GwvzPVXe9yDd3h3GM+C8NHhA93Kh8zpYvkKtiaia5Do9FmjHoly
BCnfunOwnHeyWbKFny0v60v07TbwnXj1K1BJuxceoEd173zfHUNkR3wUpDooxyp0h9cPbaQHfzpq
o8WYxnGP1ORAAhEcPVszm1R4qLiax+SeVDe7xXBIVBPv9dz2YvNsyQHkRYgIQZUDyUvAsyP83moF
IlsEOJvfWZ/tyb9yez81YJo5RCU3BLUZ39LtZAnA8CjpwAoXQuow71kgh1xnWQJIS/xbk9kTokSC
A8HhN2stou2lJyzgTleEd/LSmuwAILkVFWKyBGFvwY00T4YUqF4LLN6mahCdpM50Fwp1sKTxJId8
liuMP+jgfXwffXTpwYMpBF0U1u+HQ8SU0M322evnGVddDmehrZZEDJ4fkGEV/e8YsBanCju//VsH
N+tkXeVaOo6TkROpdUOFYf3hybLm06q+S5CS4ImKNydlW3LlI+k5o15Nvt01sajJ1tYZcGIQhs6L
gIs8Hf0R8UY25dDjsSDAK0lNePxCT1FJaORBJdWFWNY+lUxRKKdw4fM6c/uxtcyrX9S1AuKEgysJ
0M1/GSynM6tzkh9dIIty60GWIKxajq9I2idwFO0914NtQ2aQrE2FgocaFYcf5gFOxrDjlIs6JgwC
9lK2bH6ao11km6pyZKCfyoCmUVeJtjFaCe2p/eapxNNhL6zxEq5xgX5roraWVmpEkjDBvr+SYBiE
yZSmG29VIGEckJcbltsEd3qRCSjw7thbuOoFurjwyq8j6Z6zaexjH5csDynzwHeebcZ8/r2Tk4ik
Wj0DYzF3wR+/Gc8kBtOwupb6nAf2jyVwjr3nG5ptn1ZlRJuJaQdkq4dbL6usE7cpeYIM+dlyGNO3
Axs3ogMH3o6VL5f0wJRfFpcKyk4UzymByHnGOR6zUPoVkXIaYdl5Y3JN2SnkVwTmAKcMUOzl1HmD
0ZkRk7ncppYr1tdwcDE3Wco85gKLLGHMbgTyPJap0vCcwqawSQy70BYIeuj+CCrwuSHglVRpJ9bI
k32syK79e9S8xVlPlpweTwmO4MHw/3OFoS/Y2GPBJrbncEQ/kqw+quia+BxJ4f02EyUL52UbYV+U
q3TY5O5bzHk2dqHaCGPxajdO6HimXzORgDClMtXgWQtkyVn2zdS16hJ5QxdLywZfarWzDojcU72p
apZnCPlOLhi7Vo8KO/CowCDIythsbOwBKFX/Y333Yhorh59oLs7R+QfZWDj/XJ9I5zOr+nxqQzai
lI2MVOu/LcIqoc52NAhxxhFRdTBnl313TC+w51/+pxn7tdK8gWGbeXEPQUQLwNxB5PnYtf1lPauO
LNNP4nEaplpOB5+dHS0BoovKO2p/DzcgcTRnLJnIWgVcKfyNC4/ASFrJHq02lLYKTuLMOmg9Mstn
Rq1r9E8vBWjvBPPoF8JunSytTJzoHHlgNcb3FmEEaQDDtSekgdETT79EdGLihseqkYwtbB0SZnnJ
8ko4qS2L2Gi8DfSHuESpL7GpaIYBpyJdf2iMrGJJDspuTIZF/FZKWT7ti0glaPCVbWeGfyNtaFal
zWuRJfCgZv/DcKBxKRzeuErUM2LZxD0UUWbAoMFF+TyDtNZkRFqOGVdvw/QJcEEJWl/5iz4//dvP
U+aPpUHs8RNvohq44YgxOgwCab1/KO4yWGGkfKfG8/RWa+unAMmGVpEgcgN4uxc+X5C5yrcUVCE7
WZZDc/lK6+p2bGU5PqDRMPYRtCOUE5+J4NA7gVDTSCKK1BbjOz5SSKpbmIl/2+KssJtOrZanAw7W
Jo6cxfSjOVUdJ4EOjwj9Xa9AAewmS6D0rVhFXsx53MUN6OaNsP19PTlGm3BCln1r78lB+WTqCQ94
qh70ki6xdy6wiM4yiLphzUyFNJSz+xs5WxiX+wCYd83MK1xjsoXcpHr47pXxXKW4OBhYP8FaR9R4
lAljJpkX4xKva/A5yNR0RtQ3Oe2lbhuUpMIE/FJGkTWEO78TKiTxWNHV4/PLChr7b4erHKGjm6OS
L796dMNMhWIkf2d8Il6sgyUXNFzKZM/5b/LUZwBNEs1Uyjbh3uYiHMVDrg/n3O79YmtigkjOiBvs
BC4MydE95amWe5G+g57bAekXQrpgI4GDk32flk3Q+hh1jSsgrhmXveVGSNu1HrdUCfNtSSviL5Bx
5bwW+J3lmgCsbuH4n8x/f1EYNlCqYvPpYydGqrEyKyU4vDybq+hVP+XyT4FyTRehi10aA/245ipU
4z2TWmTZn3qoxh7fErsqSSybqzysl7vwglYNS3dGHRqWxOzzuMCmo6QvKXABA/M3jcZjeOHBt2oi
lI40mJiWdujtaAsP+L2/FP1331HWfS+P9jJZp2yUgsD4M9ZYQ3yEXusil4ZflKhBnMHmRYWxyVrh
pbfdlI9vg4LMt4hZOW3aLJnYBq6JoxWG0G1L2nryV7MOrxxVmtFTRi3MoEWeLkek5wD1sLGUVPKZ
jV4SwjMdoJZCAV0QXeo66u26YB5hnL30xBOZdsQBSOCmJ7GGvROxGREvH3c4yzHZNu1yEkQJArkh
2T+g8ZnmCCx3zBr2q9rc+qSQFZFZ42/i6e6rTfoF7Xs/k4vOnI2Jx88/XbzcsG4fFBLgChdhZZlB
klS7VEuJJacBHlI/KzYVBOgVj0qutanzFD18xHdv6id7TYfeK/hgHCm8DX9U0m8ZIkwBkfGBnG5A
8m+RMIfwxsRYcKD0rX204pU4YBUpivU4Bc8ouExnVerh9/oUYqQZqPYxc7FXANJeIkWmHzurmd/u
uBXv3aZZwZOzeOAJqsYeitlnn66fE+IbJPK4qO2Nn4APMYWhu6/Z+cKKn7yXYqrazwfP3w9NXS3/
nuOSi+bg9nnmd+5kbO2ya+duHdgJSrEIN/VUrc5AEHp3dLYgv1CCCiDLHO4PF/exH84acM6AlZDB
LV5VXZvncVM2KHZ6W2FHE4SDlWMtryPlpmrwEfH6VJ8dNojwQgMeRxxa3QnvN2wjpBPHUqyG9x+3
VvJZyMIQj2Ob9cs+rF/+flpEEIlq9C7OPTgwWm6pt40HZyObhZYlDZKjBArPdicA3XmfOLDza0lI
6kzOQWFaxFAj1q1YhkmCyGEX/eDk9Psx68YVI8J9AbgBwlJfLx5KOD3KVhtnfp0bbBPHPm4wUotN
aZAOXa+ttmkTSH18ejTF0U+OO1zbtPBvZIW1ACwnZHgKaiegg0swBQh3420vjvJL7SWIr09Xeiv/
g7LoWtrTOPmbbKwvnOpyB+XoIp636yxqtmTE/Cl5yLRf+wCrvTyJpndQMgL7wF4P17WpQPl5PASo
sBskGxrQppJgsPUGXZmKxknbgs5QugbViz9jrQnGr9H68+vpvbADwKtI/45Ir8yuGCgedPC2nune
z7X96lV2+cxZqmc3GrXnBtwuoNZsptSSkxmHTwbQrZuJ746b9W2bULZww1TgYaOHrt6C9yXQeWv0
FzVBQoSkH1EFDwlaNk29UrSqcrLwe1FMivFdkSX5W7Z6R5xYs1tMYEi+261CeUKnQJtEq+q09j05
MFW9zck05Hb48I4erMmko4nvP4xy6EOi6ZtbWLJg0Npo0Wu+xVbEALjf4iIHdHRi3hBzpF2jOEwi
0nc3mhwYLmHjv5BkzXWCFfAwfpbG0kXqccxnNQZ4LOFjsYXFwX7+OWot+XYYY8Y4NOrBhnX1qhjF
fp2+8frvrAeKIEAeBOuRZ7QIyE/x4l4Dw6ZmU52kiWAcRk1rWTtopsDunZeBIKh4eZE/F3D0uDko
+EkkdDSIyCwYTYcrZS/rr+zYGrP2SOmFlTRl23IHpjiC2FOngctDywC4YN1dpcHO//meHkVSE4vF
utdUJ2WcNUmn55usNGbTFdcqIKTTKyxQmAlsAt2ctXKQuZ+JP9D9OqMCezHZeJ1akdAjVo72VrUp
WpNYh64Gsa3EC2HhbH5xlyVJuzZ7WDUTIkQhNyeykxS4iGGVrA1KhpyTWcs1kU6R/Hcf/jIDQ6F/
HqVvHeLymtMaQvsLnTdLy0Wa/jUFOflHF9QWr6MRMl2UyMulYS2/THeruIe8KsjQWN6OUTDZFcfd
A/8QcoGK6TwPUvFK8/vxKShJcwtdpj5VXXDewmDZIo1g0flJXjrAzfwjM9/j02FH87E8had21B+D
FLw3wzPl9u9nfDlen//7cmmmqdlfEH2c/AmP3YtlJPoma3QTph1CBzsWY6X0dC4fF+J7K7xQWhW7
q7tFSHSES1zOC1G58vegiGSzSAR7P1QkBLEQEdy2U5e026hsuGgadPgQF5I99H0QKjwjXWNj69Mq
bQof8D6QBt6DZk9NJ+2s27RIJ8vabH6TGabknl1ii72GDAyUXIMiKL5b7XhYOStR9E1VPM2E8Mdw
AgnywU7omLP3wcwVYErc9DVzZTc2x/HHB7kChZhWOYq97sGxVz9XQ3dEH3miQ+lH2kJmh3o5Pubq
qd0ZDBg0anAoFJRJ+O8Ralpk/3+NrlkP39e1X8rD7P7u4GmqUQOx0vuKvKxK0VoCNXaeR8sWOq9S
oV/xz5cwDbSsInNShgpwSD3i2vqdPCNRT5DXWT3Yixk4iYbRsLeQzsOkgyklu/zlp4e3YLynZobs
6yJVuq2o9BDqauHavPk7aI6sVEFFBKQsBYjAE7xlmRmTE+4HAHcbUwhqNJAHuJeZqJngEbKmcu5v
gmRi9v7HfZahSofF2p6fLoRL8zs1CcVj6NKWzz4LZ4hsFsNVIm825EHTORQN6EjaV8r5Cxz1uHxS
HnQhHHQBMvM+P2ncyvn5VnYwzogRhkU3y28uAixYq3p6aoK7SF8ktXDWt6TDbvmLBQL046+04rtB
TUv3E8KVS2j7qFSN8GcezzqDk/D+lsTox1uU78MeM8S1tzac32EUPWPhOex91YS/VGi3II4jzCi5
BThmbhP5+XdGQ6HDsGgduugzewZe9yy1MstK9GDnkUq5BHVvGnfRnNMsqubehf21iUakmjxe6F6t
woxSDgWc0i1WXBljojYtVdqqGlGRfPF0bXmFVGJVukZDSj4kh2IsTp6VK3M6Wiv9TVmW2P9Xf2+Z
4TOtKiarZC8yps/0qmhMoVyEBGkRIfOzGniE63hu/QjZsFLT7k/7+7uW39KfaeZWizQ7Ebwx5AVs
Da5WY/2WNVDXvhe5MO3rpU7RhwB9AcJNdA1PXQPIdR7EwZr/1qeGpDlXznAOgdinhZH+twI1VLoy
vmneFMuRwnsCSkAf1vUkKb1RHjq8AvGZVhtXiDFAVE9YuxDnitIzU9fbs3e42Yg3GhwrPbdaC/QY
yTIbI05MasWZLQ1avV4p9e29KzokNhXJqJWrmxYHQV0+2I6dc013CmV2He3xW1fw7Q0epFX9jh95
tE/phIiBshPdT1cxlR+MqMOA+/1TgXO5cTjrnAsd+zEMjioh0wyQ3Q74QUORyOB6sWiGkNg1h0t7
EZL991T95jj53UkxET1mSb7HWl3hWRiCEmGaXqfo4Pm1vmqRd8AQgvpJlfVEBZuSbcx5nGFY+JY9
okxRPR8WmlchDkLPdgCpcV8AZS5dXH2smlKTeYZnBhLIo06cv/5fit7PS21WJFrJfepMTKrLqVXu
uai/kBjYQTybiRp4FHB6TtCZuZzff3reKSoKLVCm5pignxv9pc4bFryw01Zg09nVekfuWozkZF7v
UKkHr0t64S75uXjuL7C7NtnKF4jhx3sZuJPod8OxtE2P+bF5tEcKW4ng1c4Pe/1SxbrZ48K8W6oa
SSDOA8JjcxzoRilc9/dOckV6gUEKILMPDGE1zSu9NNyU95DbeDyxPu3z4ZYPx227kwYFmV8b9Q4a
Pjg3KRqsNd2fpiOXMy2QN1V84HgZUa3JT5//oJ89J/ODFFOnKMlkIWX4vgtD9+PUTxtndgdOmoVO
Rm0R5+gfF8Z/wts8tqmOXbBGpkz54xNzNin1UUaIEtgSpk1Ag96B49ZBfleH46vs0UgcYNYFy+Uu
CYHKl8h57WaEmQGXxq0qLvwsbwc15VP+FC2OeEf9/1IbB0zI16Q1CcNCknntT/pKTcImNrUty/FS
iG6/ZAivI9RWfDuYrGQbYfaSpz0lhy5u35dhFUDXha9LwDAfoInKuWm0QbsS8rtxHUNSjrUztg8a
V6IVmjxinLF2AgodLoKD6tsm/JNtPxyFgxBo/PQks5v9YCAkINExrkry2yGlNmd6mevLKb2lOFZy
dYloWieJnWBKbmVnlVZO/itL3nYfgKhRSoIYVbMu0/hXc0Dwn0g+YYm5QaK0ExW/+pmPi4xIi5jZ
LPwDDh/nZRo93J94XuIdVfQ4q0CgTEFlTkggjT0QkVJUwDEmhfCopMzifPTiHXXv8sXi71yJfJla
b7bRu7elQpD1j6UVu6YEFOCzaK2E3SSwy9sKYNAXqE8uiKY2YqgexJ0eOfRm8SDqzbccpuaIYV1X
cRcmtAfeHvcIpON8LxHQ+Pw/bbS/y3U66IVlkgM2T9X9MW00ln85k08DceQzN8H/LvsMNrcGb520
TJHLIqiwiOA4o0UOObkIdLkKmoOAww0az/yWo9ypawzcVWTsYIZHscxW5S8UdkmkAN514RmVXGZ5
GwbaUhlV99zixTPlGXyJHrgpdi5i/Iy6ebJJSoieRwmt9gbkKOr3CeP3CGCjn3HiILptZsoLbAn9
VNOMpFwpRm4gR4iPVjMT2jiCrhgdifWQe2inPzstAWtED6xvhYzZiJsvW4iC6u+ufCXbCls9fb+b
do+B5UdNSoNBG/pnkrbe0uXy47s6mizIRjEoYHFNgkvU70L5l2C9PKKpon5Kxt0LY9pBthN3Bi/O
QmK0dgQ/n9CcpfK8JtzSLt4pQB0CykdaFICulnYuDEAjZ2gvv949/TPOZHwkDGuPl5cyNrcMMBY+
/5vUKOLq5x83lL3AHZP8dqU5M3qcuqX0JJXvusPqQAA92Lbs7RBasE07wB/ReYYuEPuuGZAhAnuu
yUsyqJvXw8bMbYeGPOUsGoGIRWu9lrniIKEnPJN1wFH38n4Ui2iEVl65q+/ZDggOqd7r35KQ4DZN
tXPsKxeGBMZ/hhdIx0o/OAhn6M1Fk01efENPF9fIFg1rh9TCq5upRK8Tkb34BpheHpiZ+GrfxHkK
x7Cz5JvuN/ANAVXtG3T5w6NJEJn/+fz6Vyi7KNsSztFfXqhsqbJ/sThxMOuZfVb56NLeMsouFWit
ojBwYgFwVcUbjSFr7nTSoiTgtIPpbIh6ShrYAcfKOlSqGqq8ykhLLOKhAgh3uRGnKOgJX16DGU32
H0fMs4ZEKPBe1rdiu+kygqYD8vvyxO1rJKXfrAjqldd5gxYJVDmLc7FqgH8W9wlrmqfZxHv6yMmV
7T/XunofG1lH0UeJT8fq1BmCh0fdkoIaO4XWCajndZnGgM9TRaH+wDeOGtrb8Vg2X1oxT4LILONY
rLVqPX1CtosY3i4hh+HsCI1ReJrPWLrScNGBZxqqqh0UGsVcKWfxegFOTPmF21LvD+By7ItHEww/
iUqMh99FZKQJB9fNjJYQKEDeIfrU187F9TXhukfY02qYmZ+Mqqr+CMrWdOgnt/knMFNu92b5tlGw
wuGG0csMqz9qg387hBEQk3GGAenv4bZskmR3/YJAA3TebqZxJQkL/M4h/fgXA1zV8CcescUFWU1q
cP6zmzcCwXhEtFBgu8vpU8+JQtM5A6of18CNLO1HwKYa+/mBp9pzV/iBPgWUoYgkmEFdDHeE++Hi
zsS2w1DbwzYvZsixi0k9vnZSXEyTtFtK3T+yWCmpkSxTaSpQtOz08AS8WoZkg4n7hnctYFva60cl
3PmUN60AXak8hwEaHP8uuBiLzM6qNY0gbtf9w+7pvISF+MM3AvTTlTTdw9xhhItJcct+4EgQLTvz
Ot+nRRVLGNZRpF75q4+ZLOXRe3ER+FwW3BmPehyQ91VU/Az2CjfeKMzEZmAkM0hKh5K7oV8ne/5N
oK0elZmgkd6VISRThAz80f4kb7lgRVHPMHFu/W6M3lwsGkyK0JJ921xGRn5orCQ1kvRn4bgzCnl8
DRbNbl6CY+XibHyjD4SQoqxrbWYDsJqWVtsE8tb720xc99Awu/DuCWIFSJlSrAMki4o3SVh0I3LU
ChxgF+BswyLpC9sMY/35X3EcXeKZHzy5sbdvB+Fb20zj0cUvfU2ny9yUT/4JOeCNN01l6ilwxtbp
4TOhdo28EGSFOaQiZ6n1t+qYucDLEVnOTOqJc8e4R9cpQc282wX3SmdJfRSUQ4MhKEFxyR7OdG8U
yYz4NAZs0X89lLOO1me15RQq9Y83RvYP3hJyY6L02BI3sX0b/0LcswkmQWxoBXV2OBlFr+mYZqXc
jkTv2SSYRZcZ5Ms0u4wfzbI9+8C0QJoZINrWYzO+AIAusS9lCRNxZj+smXrsALmLNU3xzPFWg6Kb
WUPJ2IDwDeXZtJ8a8YQhH0VnocR6ACvs4fs5pycZ0KFkqeNJW8UOMmE1wfIAO/QNjpXdIYK8cJho
Ea/CTK20+kLiF/DtSuaDvapHoAVTvcRlMh6Fwi4/Qi1pG66qDzCSmXFvTSgiSpAgJWRdZZS4tXZx
UzEE5t6xUe+R2DQ+bavaukRZEHhE41YLpx5T/h4NdeweA3mI94bwtoT1yyM3Tsy2Cce/MbcPnDHD
gxAvDXGEiQwxqhEN25+kbil4CWSolm8xGbJ/Dr//2GCP8RTihEQ/Uz80J0RddC/sWcMzziJTNZ0T
+jhXJ7VkTSLsVEV7P2WPmBO6Y/2EPwJQACIATnyAbShOlqLJkYiefIIJnilijYSkV/1DqsyDaJ7a
BnzG4QZS14C6oed7SqWvIDdoguGDcveq+DJ24NRwUXVXQTJH5xIGn03KjQyhA6gAA4Y7w2I0J6D1
NmivG0+YCRBkYnbe6glJw1LvNqC109Pw4cJ/eEOlTsZXnUtiGuYIus/ziclTmcm4NqRfd8dHdaR4
rOnpDj1cDVLDlSqtZOenScMoKBjhgNd8CzMiUo8EaRHFhJN8DxvxVMLvJKCyE1cQGrm8DU9vst7g
CVrl+JuRgM3sse+Y++pH0KbHncOp+YF7YFvTd+ZzCvGLY3k/OVONpHjwsKoUOx9F3lIFDBVSZ2Bs
mmpvV4E3JvASn81vD7ZlzGFIZ5CfZOmp7peovRmbjt30anNNkVrdi3Yecm+vdr9XawuJmGjo0qEE
vpvnPheZYly857at27q127i3R/LtQ1YXwRV3+QPjDYEhridcRFvpls8eNbILyoCk+EnLyIlOX3ZV
+xXd4IQegA3S759Kv+xEhsNya1Co+/2Mim88awhy9WQN5XEahoNTNl7dbWiKD9wgb1X8X5k6L6qG
yncl5s4TxHkROWqJHjzPL61bxWTH8eVenL6uydK+ZvFGZTSKssZ6UQwSsprPGm2OVa5F38XOA4vX
SbY+fNEjSjKHHtnB96OCuvmVR2gr6K5jpYP4HL3wYZn5BF2DjLyi9fUEdV9/+svi+pR37it9m15/
pdBuQoDkoRVAYOI0zDZVF0PepfEQQbcau/XVQmDvBf6382N4TFz1oAvgcJ8q+zkH4fiRkT5Pco02
dPoKuIyEFaIuI8Ul8bh9o/G/gkah8ZBX+k5ahFLUMPSiBw+olJwrTNv0Z2BNRCOMTtUeKOeWPOyK
0PqYdtceDTABtLcaPVCiLPXKjvYG5KljtXMABnj938Et0dtdTMjeOiopCC12k4hFfHAxJIntSqsd
1uXoeC6owqSbaIgyrAAUswLlI2xverQTXU3g8nEMHezCOmJI/iWNv22OK3OZIiqs3EZXPwfvg3cz
AhpNCztBm7OX2Xm0LSOv2gMFQqvbovblGzB807tjBc2+zCNKzwbgLTqzMRuQJE5saQIZbt96+ZrF
r0ck1yqIaaEOR5Bw+9kEK8YtDYmhagGpy+9FMe6zER4n3rcw86jQgJjA/w33aC1Vlk0/ktLzIyww
HvaiZfNdtpRcZHtndobqywnfXd+mZj/mTh2ff3giTssibjRyTJ+1GYM3sEanN3ytn3A5qYYWyG36
6Jrh6bz9j933/Uao52Wwsx4Op2RcR1hggeigYwcYWsWKCh/8SrVcEcCZx57+/i1MRVfQecTUOjai
da0woMNM+qFz0nVHtLITdFyRU4UvEJvNp4WqhIBRZ0NZ4D/+ZK3QLrd6ggwkPzZrQP3ddxf8SmRT
D52R1/aS9Z65s2pwdmnZ/i6V5r0i6P55b0I3LDVwq6+flJBv5MnJsnNiCnXCIcKV0WY8+9wZ8O/K
HMAjZFA9yaugr9ic7BkIN22w/ggqch3JyLiLegOpGgrbIo24obyM8kOluRyEoQpbpla3awe/a8gh
FDeM5Iy0jqyzfh0nzWz8J1h2IG7G4EcjhxTPspoZHKz3gfABeNEvywukIlb2+FPcGQQE+SDysQq/
ioWi00dmpvVn/MHWZOxVqxne2IFDEYBlYjJYoBfPf4xmlZZWd78wb6/l3iRTzF4vGEpHA/CF9ZZL
nMmeR+u2LEIN+HmJ5D5ZAfvZCIO2WODjbnMQdN6U3Y3veFJ4F9U3qJY04PAVKBqkuhm4nKCe6s7b
hAczYj9f7SsKTQBe7a9XDv651ZCDfxp6S8CxvyOoLi9CHbyNKzpVKxoU5inx7JPe2OzOcoJK3AMJ
4xlRUPNpNnZZon6atIfMHKtkWGJCeizdTvmWh+nvkFxVjU9niFy4fIuw+GNzTWvJV9pltsK+8aXQ
1/lpgvQk7OAqc+jH8+yToVIIi8dBYgBgiYfO1ukk1P3wwNAjDPywamQOo7n9cmZlj5RCfUXn0JAc
mJ0l7Jmk+mwjh5H8iN5uZFDZn9yHl8y6LEldwGUYWPmTPmaKF8e4TUDiQ6os8P3/x+/uTnIsujgl
FOvfETDSQA+FO5aIb0x4G8UrmpZNxttDcPZnj7AgL37l7ZrrLFpc2vA88EK1HdhdIFUQHLbYO0yF
QubjIc232hj3N3Oj/3zyq9j2D+KjK4svqM7hi+2//X1rVtYcrNhLVy6f1IiovfetMLU0mJIQdyp7
ejY5w7ezAyxByz1QkoE45265n8FnIyFKAp23xDNrvD+5e+/jRdB2/WwE9xXt8HaESfN6f4GlbjHe
tn8vqsfZ7qinvwPA+vCyAf9ZLBCm/UXZWk3+Sjn6wAS76+WjucaLLt13qqA6nYt8BJqLqqznNVPq
8FZF3/d0TJ0DPFFlbNybtSce5ycMJV6+9ikiG5Iw1BfxjK+vxlLYSHAir3lWd5YDBYAJiwTm2HA+
Ox2RmzW8tl5YrwtMdaoCURzcmu2U3R6aDaduB/d5YmBOgRipGazlfsyEsSAMq7J4mw84zVtw3U3P
2nJj+JCE2YxcBcrpuR9nbkYmer/Nc8QT6mbAV5xe4KP6li4gBfz1UKpiIbKarb1TJcX+ICaX9hx5
ce8MoEExCVtufSbuzCH8hqbO1+3PK8xMm+i5Z/f4pUqPqI6iiB0q7vdwkue5XTm3imaHyuGxCFb8
SsLiW67uZDAFkdIOxo/PV/6eXw/eilKxLp32nUU52sP6LBOWHsOgNdjnKrW+VowLWH/KYT1iyJyg
Sg6Gc5CLp679W1nKWr/xVDlODAr2mTlEmLi0APfvl2Ud8YZ1Ng5DfJTBn40sJoLfOTCaPjgVejpV
OyVc/Ddo75Xqrof99hlYs147cTR+8X//tAB7wOamuvZt3zt0Nm+XE5FniZCK+7rdwm/NmPUBr2rm
/4skdX3dvIrWAq9z4fzQRVIQQKj+NnKFS84FkKMiPMjV9YdcpeymUHG94C5D5X5rn5RiJa4+DtXk
HB59k8nRn9mFOgeAFbchAtXybs1KBP/6r/7FwlEIoD6jd2016eNjJizzZG/sWHsaUd0JTxADt9dO
heUKL6eoGOjlmgxek2EqiA/FUZLTBh9GGw8mtkmDn3sUdQbEGzUNMqnZQJwxWfALxFdRAicuj4aO
I8PTd7Q/eipMhhrOCqT2V7suiJ9ereiwylWyzzKeo6aAsCVzCobT1+GtDDZi0ZLfJdEPQyLMfEUa
pIIrbTdPF4gWZUtezrT7Ofjy8uts6prSlckHaSsdWhZYuLslWkCXOG4MWBO9sBQBBG8nKAXrr0GI
Au4iG9qdT8J0++wMfWa82Z9f0rvRRtyr4p2WQs+Eb39RNZ3byl/fuDnzSt1KxdrExhZDyK+v0OxV
yWPim3o+Ei+hYmy5E7kvABzDETrltmMbEDPQ6gS9fDkBL/BXAiQtDbgubiNXwV0QGrP1P4lNCiZi
tDuXI+xqrUMSz3rcm5dlHOy0S/XsNsiCsAtVLF/E+J3ENuRkcDx318NDa3ZFyv1ZS258YdNWddAq
d8J8NAhO/x/yaM/2PO25vsD6LaoLXIHTMKKj53uXpChEsMAg//E/RjFjO36gyq9PdllhnyI/Azwj
HEMDSGMDXOgQChFz5aM45Co6k/OP3HiiH3zWfzNFeOZ+aNXO0hFyqtzHc2YujDl9F9o1OQiZbEXW
fokODp6EvtCP3iwxkDFpFzmzBlI73Ixjwr0I5h2nE54XwU5ihUgbu4Pz0AIZW5ZgDNbRVXss1+po
VtMqw8f7q0FnB2ZRGvy2JA7JSspiev0nWtUvlZGYie9UfdylVFwVYcj/yCdqEpjklJh3Jyt2nmvs
+tpqCd15Q3Ea6k/iyjROE5wNoizJ13WqFSt59mGrQUL4HYtO/cbNja3e9nAe1qME3XGSl8zD7vpy
5y88EhOVdqF89bkst9s/GxaBYcR10TDM/+y8UwBk+8fHFnc+K/gofd/1doatDAMvtUmwfDX/JQyY
1VzTeYPmn07q1NMBlFEt5ZZRewAtpZaehmFSpBbnyexkenujnfXpo0BPAG7bGFNt7auqYepEjYEQ
Vlzqy8hAbhn5Iy2TUGZUs0QgYz+byyt9KbX9kGCnY3kJYb0ZMieeGI69FaOWCcDtQqCf5okAy9xt
d5PCr2/NvUrI+r7e4QVKpCMgKRYKXr5urYmuGZqRWhiuGwG4TMa/vyHtnXpJHatQgseUIrnYG4HQ
+SUsuUFyPjVzhxyWWNXcLTJwXQc5OqwZZXooDtQNuWPb7Xw3wua/4xRDpzq9MUQRR7sZ+F1yA9Qk
aOPiWMpw2FQvETFdtDNLNgtMTHZWBbJ5JY/Wc+YYBJyMRdVe8sLJ6lYdHPe36gk+PTQoZMX+Kp0a
1j8vf9BSq1q75SYB5vJ99lNDj/8uOwRF076dy82hgipJK0x/R5aXdfUOzc2+u56r2oqYeLVnUEhW
Bs8iMNbmWLtbbTN11IX+d3OJGdxne5603HbaKlH12MKUX491aOtHjuk8ckhnS6BNHyW0Miqr/Mqi
3IAgmlOozT5ksTZY9UPzKipMDrej7HgofrX+gg38YHBEb384Af1RFjK0NZN870J/9dLJgFxLqpDv
YAP3M8TSR1/DGDEY1iwT5XKscBJwYi81W22ANGqs9dubtcRkjAvj4VAoBDQu+OAfNgDuyzmIXKjI
qxSUe3IMxcnuCd4pzwgvmaudSbqPjQT1vLtOhCu8HtMJBcMWGFxAv7PlK0Fh2Nvyo8FIgHNczmgn
pITFWJZTWL5uKyALfsYmOj4eKoD6wDgxnkgcXx57x4KFGTNES6UASjkr6IA3FJ4FS0k80KY8Zh+N
1CjFnuVX8C7eRKCqvNvb0BrevMuaUwQI0EYLilPEulmdZHlIJxLeZOHw2fQIbwu39ls3/Mk1TVL3
GZt+Li4Y8yOHeX++2HLlFO/4S14YmUSfQzeW3S4hingNO0FPchV++9KVasn8u8/q94M8BQqqQYYu
447PwU6szWogtuhrCVoQMJy2KIFuuH+b5BQTL3TjLKkIDzNIkSatsSD6EV4UvBEJCAu6jHQYv1MT
Exu80Bto0XmbrJW+QifkoHvVL4HKyxNc1IYUDBsMsIsckc5nQCGPaDqfAMJWfkuJOQeMl1TlAX5P
m8V5n1wSJHfIaKEVq9KFtKsoyAaG24kPhfzmT4enPHkjCuBK/F6Os6XqLHRTtV61CP5deFCXTtOL
CYtH+jh5x+ArVRaesgb+t9gvcFBokLMULItCIjvU2yBT5uWRJcwwDwlZlFDek92XlRkteX3Sdn7D
17N5gtiQ6ENUSedFCjyhyd35SCrW74rksY03sPjO3cVSQu5hPArd3EsYY/Mj4oMFVwmYd1yCGGl8
JNgDOPGLaRZ0rWv+cIkxuduqZgL8K1SR29maB791BKCrk6MfTHfafQrvAqUU/omWHDL/EBGsJ6ah
GqDV5RSiyzs0BMeCqn+9r/F9ZmT3FAyivFDFlun0Ej60I8b0/eCEiVO6FRV+EMq7xTgj47yWYL08
tv3nQooQnfAqqajbn27PB4RvFjLntJk80P3gIjPUUx5LNmeuTXHKlsYZ7TvY3HPzM210l7eQgb40
KmaCOJftZ8NHNoaxYjzV6W0/y8jwwNQDRHD7tuPkGthB6/p7CQJe7e5fgwfl78W5xZePl6o3x4w+
VyuY6Q6EAvLodg0lDNCHtxgzQ+qbOrz9FJUfQaQOI/Aq6D0yfqQmGqujI6RElKClIxzTWNc2q65N
OCMwwnAAIBOURarEYl08pcZi6jn+C5OmdQnXIPD2BatVAmX793WTu/Y5EwzYAV2luETmzhEBlAUm
+8H3pk90cHMkMn5XOqiyrwTHJYSMRg6kUo/3IDzFWAWaVTs9O1LCtJBwI8IdSm89nivNy5NjZZFA
jhA3FJJ/3WYOIE/oApCURx6AIrtm1gJjNRzQAJXW/vvzKHevM4OGxS3xPvOWKuFak9aPohmGgPCk
yCX+8OY+K+tVhj3HalV87nFL2H1n7VCVuqCYkxwRVCl6mdXCHHyNbpT0sGbicj4LpFiw/yJ4esX/
REUUe+SSZp8ge4mZ304Rh8MxAX0p46bF+1uPfv6Y7UBqWBOdYqetHmIFsB4pZaid4mIlBf+qwfzG
qnqxcdKuovYrRPb+plIiGVJ9l01Qvs8hN+PQ6eStvq2M9mllxVJG+9CrMmnas/kR3s6YLKBRVzuy
cn8hyqDKUO3859ejT0cixIgEYtiqCj1d53XVKCKtWis3kmPOAThWQUt887UcSZGfcfR+amcP7neU
VJ9Q1D6/BlWAtcqq4xSjMKdgN3y1NEXdAduk/HV7hUHWOwdI4Ot166Y8eXUJeNzxpjp3wnkoteQz
hcJxPZIwSp2o3O8ArBREyG61AaJinhHtvx+o0voXJsypdRCYJdywULx4zCSCHxyl/Xgyhgz4AFVn
of/iC0gOR7UJof5fbQKfXN/xmICp9H+WrgMZML5eXW8qXu2iCnAVpZz70JP5tSOOpNJVoq58QwWG
iLIY6IrmL+n9WQyVZS6DZLsjveLfB3B628rXDQamdMCBfb99bRQOTyCZx2aPbCeSdEzZDCchigUJ
RZNBX7PQ1itS0+9+8ryYOQxdpMewnELFE4ysbs8lBTivJn3pAoJMZDkmLP7iz/rtSMyPUrtpjEwp
f8KgjhzB53QWAKtTcotie4sB1VSlOXPtF0B0G8cg717r1K9rUS9h8qzl9bkDCZf6X4q6rYjgVenh
My76L1t/U1Um5qgCr1aBRi2WusrSXmt+y51L3Xv7m/uKF7YHwJb5cIujapVZGLOCaJtWiYZikSan
o1t086pUXuBcB7VHnousg49YC1FJ3u2m40TPZmDmY9TzkhIlzYuJrnQoKx6gBeqtPOrsC1pygCka
BRKqavuqSuAyaSUBBj6l7n2fsy/2KR4XIc4zTKsaqvTHP0oH54eaJVQY0JUsaIx5LeGX+Ne3q2Yg
02tLrvB66IMk9taYnBz5Luj/tRYjdIYMN5ImGC1DrYjY/0Vm7HnCjJaes3O5j3D7VMCrxF4Voa6N
0yLlU/NsPrmXPKie7F1BPQEMNbPBaNwN7tpAc+sMMRflQf/OtHV1b7S2fBKj8yw+1/BlU5Z2FDTk
O0VLh8TxXzOknWQhXEaL5oKxe/KZ4sD4j9K+Il2wDwIOXMWlA3/8lGbfb+w9Li++DP/sEfMMZjaq
JSjj+Kz4YENbtQi78ddma/U25rVpyyGz3EiOL0YorAkD5u6WwHODgMUIllUS+PDj4Pz4eOY6T8od
RDEvnA6zCnX8UZyX62yY01e/NNO36JeaNGqC5bkfLNaLhd9Bo8LBwdkAB5HVw8aR7Guecohvhtgz
N3fquYSJSzJlz5Pp2ZH3wSyDT4ytw1TEpM2Aa8amZWMqHsNkuNmzkvzPzvOta25VCxRLcEpmD19c
WtCZn3DnJkhrbUHK0CUYj6yytllh4tQtyv3+W2m6DTgZt/Ba00M7OiEGhyq575rfuK/O+kj6k7OF
S07xVgfDRev4J4epvK2Puw5V7CtcXt0x2Ft+vCArBUii5QfWBn12iMAjpwpOSVh2rVsy+zz8cDhu
kGryXJHTc0aRszI8czd1fm918i6V595Uokt+esoMMBnqxJoFvkN/h/pUmswY3gzLHzKQlSpDu/Ti
h+rMxonfySBmpPlkY9xs6YCDZFxEfz88wb5E3E8OolfVEUZIZW7iXaRX/tqZskDY8WLoSAb6wbhT
I9i+anJ49G15uUp5e7dSxGLj/7ahUVUGZvAm8CIxbkrJUgiltoIMrZNEnkQxZO2r1PnuO1iBKz9m
he6gszHgdgzHP3wt0TlLjWaqvaC/5eTOmWZ+1aRi2pQK7dNp+8Q8XGzvTx84zgRcPim9dNI+TUff
CN7nmKhwMyo+tVSI1LUN0wWwXT+8bZeRgVuDvAF7TXNLoNRKrPRZGSjCGxxJ9XkwDnjkdTYQGGwH
LFetygdqlFh9q6bOccTIxvLjoRhuZzRTvntPZ86d2rahBKwZiQuxjs74vYytwMb2TxC19KP2U21Q
2N6eqYqzKOYdZRbXEVS6/F9SiMWffrl+FiPb6T0LacqPAx4Y9iQHg+mYzSx1YBeSMLRcea7dh5Id
utyoFgsTBGKhx6fMTY8bXWHQptL3cIGyVILT+dCNsKveQhRF6inwWK/lFos41OUVvRX/5AzFTnLO
EVUIjBi8NNWQplTS/wygL38bon/5QLCKJBwQf0YesZMzuf46HZrDERsNrmwDVit1FqqehgMEIzdl
IXNSgVhvJABIMTYBpUvtcSEBQC6Cqsqvc0j8uU5l0zW5HYGCCRYcbd7O2JmiPaVmpsA548KAYnZB
u90=
`protect end_protected

