

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XoDvqNcsUAMVrCepxGZ+692mBkX+rCE8HMYzKPm5R78cJ+RMc0dkNWWZsdClXOY6y1T5UuLnfOdJ
4pIk+MIfbA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GQd6VykDj7htiYnOl+4WVHQM4hKgz1J8Md5aI6kr8/Lamm+PnYCv/9ATHhzH1x3ZwU/+Hk75nShM
Z/fTah2o7SNlXBmxO/TZV+Cu1NdyZPM9aMjSfxhjbc4DdKhbt2eR/JXlXgPN+qqN+l8aDRz6dW1r
rhTiAjUos5V3YtoS0kE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1H8fvXKZG1QF+UJtGmRK0CnD8bm/+01l6RcgU14qYFFE8GVuJpGQyW5h972p3ANLjy1WRtjYQ4xM
/dkbNa4PXjLXaYaHj221vfSd3lB0MAvfi3uUVJSvclNp9cIhjsynHt6eX7sY3mGpxNDMKipfks7Y
7QsvE6SpbzMkIaxn/W/Og06vrJaRobnXPbk5O8bulSLgRIfqtOFawh2LDbI1+cySFds9EMjhPXGY
R3cSwZrw9voRIz0AJIAvvOBrLoxc5eVp/j0gskNHjRbPo5Gkm/B0oz1Ia6kiZiwtS5XXf5fYsvSq
8ip/JtlfeTs2FRpXweWaPr5rFOg0LxkGg0mLCA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7F7hPxr1ObCyOsY3iC3Phcz4OOcedLcCp9ggSn92l+/8vc/8WokvA1XgYsChaRHJl3lXf2X6jfk
OU2I7E3QgZVgyd5+syjWVqouw27C41FFBeCuGD1GtzyBYnFEqdtK4Wi9fPab76EJM+QSrUTFTxOM
vNsxaERzJOCdVgQoGH4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DAf8RFZxkL4Com/8UijiDJflLxIdfhDldD1zcH1XeixMo5g8/n+Yg5p6ecx6wthzScLrbvkfxjSo
INrqjZhuOy8JD1hgSySspkuAnlB/pYzsB41QYrTQXDdhODLQLAYA4QNlYnc0Hld5QRA0QsNa7b9I
jitn7EoP2gA5KtAm5w8Y3SJ5GziR/wWC7+Oq7vo7hHrOsipiX4kUa9vhXNaEzGvrcPOJN0YgaqRR
HJt/OxiJdqU+tEWkUefOFMVnQWevf91iZ/Fb0oG88z41wfeJt8eTwCR6ZrUTPInU5uj9Frdns/GT
RmMrsalABVuwLraRXdip/IKnMD1dw9K3eH9MHA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94464)
`protect data_block
ACJuJVOegFbQHhCPzRNZ/JF2jtV5PpgAubfEMgzHbGPWERPEOZiPYY2YwD+fWGR3cSqfxcXo4hxc
O8OprzTjm2PH0U0718ASvNRNA6LPsgRcWXKTncxCDAyd+sth6oG/4eKErkNUFsb4EexzhUGiHSFf
ZRltWKfTQQQBrPKu3wYW7VVzRCtMrjQ0xlNJE3rXM2Ri1zH3olEb4asIQvX0FqJB+3UoMu2iG2zv
xRHgZA8BFjamG7YXmkKzBOKj54WpasalFfEQhKpArJxdIUcmRcMYjtVXLu+dzDDd7QEKMqGCnP1Q
8gJQzXEE1Mbo+lzDFS9STjtITp5d1Ur2WYkI4euU//FIlUpGmEGsrn3R29q39qZvAWmh/6C0gLIq
9G/P8peBuN0DGV7MS/uqwMWEWmUDItMeNhmEhJlpVG4CP+AJoz9XA7M7nyhqjH7BAw6yXSuvbq3O
2lQj+5cj9S5IU5aP1HQYcFDDrFxXrzQLAiKoDs7AZmC4iCw5ZhC+3Rr8lZlS+QjSuyqT/CCeX553
rV74SVTtZJ843C6n9qwHh1P5SGwzncPe6A3Orv564LcwNSjPJ4JoU/NwbX4JrxDmKx/Osvk61QwZ
mSy1pJxwT2+iEXyuMKhaCEMV8RuHZ1GgzdSnJEq57y+UKmP39oGoogFxNFLeoq+NiMrvrhFcLCnR
0ExlN4xggDR52E9pa6veADFRJQTY0EeVokwZtVm0HGaJuWzRxRTUSxZZSY1CBf32VnYeUVsYLgAM
OTyY+tZuwv2fERkPgzJVeEi1ZdjH8A5WRWoOqhRXEkF+GNt9I3RsDsKwvBI8jeDbOqS7Bcor1k1v
Ya0cRgE5oxd4XG3VeD/gH0+2M6Xl7GJlv3RHbo/aRvAL6Jp+d3T1LitI8F9NQ9WBQXVieh1eKIiz
N3Hc3VXHp+Q7P7HrrorJC7rJ18gYCaABcfe7G+vI7ymeeeEhniif+LlS23QUJ1DYSeIVh+oc3H4M
5t6dFQYZElkiq8J42S0nlGYheQTHAIkisWaU74WK7P2MckT7gWGyD/TGHskNCEqo4X1Zc9pIyrCl
1PJ0eWHBWbXVY8dbFDtBUQ2MY/9rYYaXIEug6Wgbicl1pf8B4nD54rjf7G/gE+QIjhYW9z3qfKz1
Lva4R9yrpK9ijMJqg6rEFK/jiwKc/XRC4pSLcmpr0noHOpjHWn4FPNkW0DYcnEzfF99WhzD93D78
vDJ0TV/BS6TtyvTzcQK/CnhlnJV3w8ZWy5RKQVoZkg6emOQsnaYRF/ixp58QY4iIj4zmojkzDM0/
rwtUXTW/ZJeCuQIbKzkFvbn+DUIdmsZwQqtw4WR2pWNNzGlZB2hkB6e9Yip2+Z7oJviAMVSmke4D
9NS7WV3hPLQ7om2DVshMU/bOkviH277xyIUbatER+xJRa8DpAt5MuD+0Y4mNbcE7sPby62CMiRmy
kACNR98tWL4oqgj4rjtE/0kV36yBz7rYXb3Xmmpj6X+TlYrmSLTM7r602lroPJ1i7iP5RgSt8IhF
TJqDQhSZsaHsLJGgfT13Q7dQ8ALfQJSozQpkKa5VRg/W7Ee8kCuIVOe1VSypcHqXS5p2Pq+SE/4m
HsRnNu/i6sIjySGlXQ9+bGalMv5b9xiXc9uVpjMbVc62qH/9Uxr9Oc2rFLhmTo7Rx+ETvN0OO0GT
JAwODdUJnQgIPWaCH5riTB5GVE6vibJFJ7+qH4xQFDtYy6szyng6aLs127nuLvp2qfKyre9Ia/r0
/J9Lm3Ctdqp+K9CrS48BgTiNtoZJ3no8dCehvnJWrWk0Zk9OHJb9XyGcp0O9CqgKvVXSdP2+LMgy
WFfaYxVtM4axmHJVg+9ExhNNo4cEtCtaKMj+w4F9Hq13N8/pswxNwmfBWtBUlndeKJyFFcCSdRBV
w50phSXYUHQ+iAYEj3wcFM/VsAu1RkqIkOGhlJWJ1elT9kdPnPudsCFnRap8OSaRAW2aCInIhe7g
qYUIiNGvh5QGcQykQ4EG+su6PGYGtAE/60vC69dJ/pXKxw/Pa1m3a+fuh4i+99UDBC14M6++N8ox
f9EjN9ZjvyqYuplub9YioGaMrWMOV9s0r6vA41PJz1nxfHgHGHbUque1g079g1qmpPzdM3eH1WoK
rqSCiYH2TuXPgm45Tcl8ag4KH4aQOUiA2vv3ibaA841p26irfwBh/hsAC7Pre06Y1H6R2Lf+49Jk
nEs0egtmz4/+bSxIhZGKtoP/PKbwTOYR6saP7bkfCfZs9CA4o4dgptSLWqkbfg5n6FwhRHkk7KQq
zfogHJpFfLUbItpUAXaUM7vFglwQFzBH8MtRxTs/BJCq9HrQwlt0kg9hYOU0BK6+JFOYurj3Gqq3
1E41g7ZocrVAEpAKYfgtZ/7u0ThdLZsWK64H6odK0UXuIiI7lMwP4TOfMrg0aNe58B88wX4lr1Vu
gccyI3vl4c7+wQuoncnMKQWQ0rBk5HNlGLcc+wXD+xp1YeisnZJaHnHrg7FL/JsZswxTvkOA9yaL
aWkvwYpUZeFvszHUoQClJ9JKap0w9c329yPSKtGNEPiKWhuZQZzobuBsOEbs6xfGBJXzfuNehnXF
jcuujWfndaGk9KI4C+CMANkgjjmpqfAc0o2AAelvt0bbku9fFdvaSwfEeFNjFvl68m19p9Dp2lYk
HCWJnrsKoMIDu4xgePudF3KTd19NjJe+a4mTwHGwmSjv/RszstHl+Rma9aILKlX8XX022jgc4RWJ
YqYVzeNcmZx8pxw3exD59oVstFJ/oa9v//m4Fdkw1G9/i1NQRkAbZX+/nzNAHPtCVvVF8QmHTG4v
qKRdWL6AH8+acG71LyUX4r1mZ2AK4y64mGHb93BY0hEHvyJzskp0A+z4KOHunt+89n7xaLpfeqH0
usPvULq+yFyHbMfqtjaTJkNWFOq0+kstFdG0r6faKY5rmwhcXuhM0rphhNh6YQAjNeH3fmhidolT
2KlMzCi0Zgcy5vhGgwAzs6/m7kOkVPVifrooyEorQnAaf5hx3lf1NE6+ePPmti5LiVn3UH6FgmBi
pZHyuwzm/Duc26zTtA8JPvf/7I8WupM/vARasS8ohY9A92tmevZSWKK7SO/nPNlPk+CWjMUi0wFM
jCBD7K0GRoLCFlq8f5FZCPpqOybXUyCca9t4M9HNYvq2ORcKNm0dhmht82PNfDch+zL9nlhHZUyp
XJahe7K4tLEFKbkCwX1zxCxkKnylxFIxLuy3nfr4ApFTZ3D2f9GsusTyPTERwc4+ge/qhJBauaeK
0oOYbfl53cbSPFM1FafYTbcBDknpPZ6j7ikzb5PDquY4RS3w9lMWHOHKSjGn5sjW3ojgiqzqVX6e
zC9XT5cG/eqQ1HoWoc9XRnE6qtk9pxXLwVU4RfvLKEJHHJaVNrgy0DMhR7MyZSu6gUPq4mHvSWgL
MSpycP2LgeCS0xTQiRihYVE5B9XLTVPs7RaDa8EHk+uqQg32doQJgIQBEu7BRA9ML8TPrxhO4UHi
1pS5jRKXPmNkVm/YQVD87HgPF9JWlylnlN40OzO9h9FmTpos4j/Wd/AsSKJhGsseQcd43rcFkNzx
1epvsqoNHW/zrgr1/e8ki3WNOXybo71y3CWsetjNpmouV1mZRHJ9zBcdL+M67EtCIstkyXz3CQ8x
JSm0Gft73EZ/jEIknpOuG0kJ4bhwHQXrouQiElFqQbbwOJvth7LnBbaKvfkvoTHjZXFmXZpyiFBc
oDZ+WvPWlvgqgvdXv/lSEyhurc4NY3MiuRpHReNLWKt4TrK4N3dYSOHdVeVZTsxR0k4EWTFPiEzf
J/kyGARXMMZna7d+z067MDm4vapgC9sTfiWz98ttnz8RQ7+8AzJqBTZ1wZvuEDm41hUmRieUjzH5
eNPRMe/IvzRT0TmXT6kTfZLH2LYzyCF23IlItdUWR2SZKT5mKQN/vbSBb7AdOLiP2AWsqj4G3L+/
3xnoF+U13im2YRwKRKXLuw9M1Y11HULRtb5lGZWYfcyKFmGeq/T0tzJrF4H7AX2htkoWOX5qM3Gd
RuEpGLB7QXeWi3f3I3DxWrpwWj7N9eJrAUIUKKZnHxr2XWwC3JEf/ELcsQzrFVIdPXAF+J8Qslf0
0cq2oSwwl02+ES2d2uvH6Ro2hE47UrdDzDfSk8M/flATAIymJ+cu3OUgG38SR8X9tXUGh8oblx4J
zWygCCvdyISb5J2J5oh5R72nvmAMbmhT4qXmCIfDZrydgWM5sRUApqWiJ+bxtsJMK8paP307UO+M
Dicbl1UZyoqMqNQyA4EY14IRzSBpV22QmqXu3I75usA/Zwe3h4IYw8jWmo7PWPvIUgwzVqG0NOIA
EWtWi8t6q8ydKaz78IP7k8CJ+u5lMHMkSqtbWCh+gkJIxdOrTGvoTxtKunQdziD3H+QQj4LRh+EH
fW9P5IsFiKScKjg0YtKuF4S2Zinwg7u7P35tOdFfRIPI1UHKM4mOe91hM/CrTu9mbCKXHrxfqtSZ
tueaRAx1MYrck112ZvvdOYQGZI0gNBYnzLJLwe/xwR9mxd0sBJe5SAWOgXrn7Cvc6nNrJIATgJNx
CI19mOC3tRhAWUzGXqXdYWm9oVtAjfMTC4CQAfyVn++tLhrJSheX5nkZJEtw9I7MveRtafkwgtL2
/0v6SMIgbDPaHs1leyBXFU0runfYvpEEKmS8EGIklQhazCUnchyvfTTQUuHs9yc3hxkd2tXWKfyU
pLXyTrW3Vv1HKrhdQ6pQPSjEMyAatbupBHbW+JbPtVi3geKvNQ6tarZG+xYjlDMT7gCeQYrof1bU
EbtvktaML1mT3c6Pex8vrzUtlnoq8Rxf+62tiPi39jqsEcA/1odvqq0ZHj0LFESYUIc2DdFLtm0m
P2EVhGUNSyBPNE4+AmzIklTPM8LUuWBN5lUY3ibzIgwQ1uGgQ68nJ8oCG++EKwYwFRAqIUhurETg
JORYZWGlFMmhNPZvfKzzMyojO7hLu/3VCaub1qZQQgW6unO+DNTM4Zg60qXRs8Uy1c5XddLS8jpb
u4u5FIkPiucAXM2WIk8KdDmprgnEHV4FGuR1PuZ6/pKohOlrxsN98ZtnnZDm2PaGLQ4HRYQJ+q5E
q7UGsRJznQwQFEPJd6/dIpCORvDV6HzSd9A5eJ2i05JK32pnR92+Om1hKc31Kly/UpC3lPcBlN+H
8qGJQU+/tBtUfzyZV1RhmdqKX8mjCQeAODd3LM48x1PmAFD5G158HwGHSQEE0w+B2OWDM3ZN0ne7
FfZz2UKiINn3gSiV1+sWigwQr9TbnQlBKoczoGijnN57J2EcO0qUiWQ289FXj4kP4BQIE5aVv+hq
U3PmAY3laVJyGT0HNqY9epSh7Ae2YKBPGQj+FmX8opLZOlq5FuAwJVPBcViCotXmtWswTmYHlp0c
2REjBCYM9QqvxbhP85ss+ijAK747HFtPjmyeEt16omqAWtpPuQw3FyWMYiVLyQHNECaC8Co814O2
m/Ed4RH6JKgl98lqSMKPFeGxGlrOzEkF4wizvwYXu45yE1f0dhlc65gfcXfqBUUz7l+sWL0Dxe+E
oaM3VcX03h4xDTYhUy7agHn/vgj01GOHmen5gMWIBi0VsbJ1oCTeSASpVql8V22aw+tPozqXHMwB
d/153lEUSxCQOzTaS2xBwae3/3RbQl7H2oxcC9UM7bXH5RIc+y686xnPQgNzZOTEmkhBkK7T1/fR
p6SYO54Wdn6asDyaARcaSDeVAKEgmeLpeMV9fuTxeyKSapNmrEM83siOJU/B/1/j/EopJe8URCyn
ZqrQyTqMyDzkzlTKIZqnvJFhH28g1ek53l1xeTfVcwlIBiMQO/6kzIvw6WBy2MIQxF8+c4iHWgL1
hr0ubQlFtx+y5/hRjP3laAgN6lTEM6j0XFQ6+uIUxxh8+Lf3OMFGB7wy1Ziyfxof9IrNyIrjvsRE
vdGNy7Bc2HL4v1xyFFwZv/RC13MYgfhiNmhSxMyxzIuuUuU9YTE36iAjyABhKCdppL7lbh3+5ry1
4egUIggc/elyg3umPHcifej2NDWehfanrLmx1nSKAK4LlqSnMSSEBuy9YFYBc3rolT+H1X9YpNQQ
v99kDIEdUU065NNKYuaS7M68X+cB6LZr1AanhjHbQCuvLAKgTPLJiad1pxB8fLxKJ9OSLFOY49Px
AVmZUgfYiNqp/XYvOt7efSZmxVW4zPc4l7dF/gwqaDOnk74GpmEv22+HYRQj152UIWQjaG9yKsZO
qdEl8X7knxQMIG7ZUWArQm0ebiciuTacXQzVZg3KZnq1y0TGSp8Ho2B+7293nz42WzA/XGRKU8NE
tpAuHR48cLvYWkd10lLzE0/erQBdecuMKiPrAk4Mmz4PNuGYf1B4NVJmU75bl+JYuyKpWKQF4n5K
SuKjHgGN8SnZ5NRNYW1RfbZrxJq6dzZtIs3GUg9FST0i+B76sgAxjfQnkijcRQh6cIArwionWxYT
wfpSAJbnq824Phy0KK5gs3JRuPxw9+GGCwpsFXumKpVV81fe10ZkNxvsYRutqBrlHW1qv+fu5TA0
s5zVnZ+clINDY9eJyEWFfvGLl0otjOzaG+oZ8aEK/1YPRH5HK+XQDP2USFeJctYv0XQdKuE77ago
JeFWCaPQbeG6NJg6JlBqzNrN69w9joBor0y5NiYz+kMPFHQODXBsVTvrCAK2z005Y9Iu9BhyBT0d
zCX5/vEN6G2EYxkxJGRUnpVOfQdirSHC0refh+E1Qp5Fl+RlY4gppN51M7VrT7aQgZYADe6m1bGJ
fayRBqSZ30o8o4o6dVSlAQ8+MAIJROThwleU51AylzPMdSzcrDjSUIsLq0iLAHUKdg0PHkEodU/W
2/x4cbHaWT+0reTZn4p955eh+jruvzUgvxok+0S8oD73FXfUPthOUgMh/ohp+4/kqgDBGQqyK0vO
DRXKzc++XnmZ+WzC6UrrUgC3Z0U+1mrrSNyn8n1CVPJHcKCqZ6O5athryY2wGLOavnkhkyzHXItn
SyE0DSVuc6GGPYO1xMwyL8inKjFTGGCKE9QKs73BY8le5BfAyTBx3i9jTDXIo2u+isd6i4PFZSRt
zXQJlLsUwvHWdpT14vcq/sR8j5IAR5fQm3uVGSud04oez4nUc6A9Yg9My6DlsNrhW6w9pK030FZZ
p6j856OiyjBWcoYoU34ertTfVJEMCPAwQr244Jbr9NRN2bKUkR7dxcoh6qMEP1gBrjJFmukP747r
6CxTs3vT2s9C016eaLy/VvtTkLgFLRyhnruhWl/QbjbcU69mY2bNeogVts5VOu5eP4LXBmbhF//y
oNYrciu4SoTvE1S/bxOB2aNI66uA5Sv7Mqka5DyldWNBttKRkf0Q5D2PoeV8H8xumu+Dzww5qmsz
b/1kbx8HdeYAlQfLFNRzk2NbYWTVJ4PFh9XoMVAKDIeWq1tM2NiQsHAf+wu5c+HuSUPqxUYJ6M7c
867b3TnUdVCU+4z10NF2HMZAmImR95iv83RnxC7E160dpIu4BuMiqBpMsURLxBeBQz/AK40V2x9z
VqzkOpeeFRWAbGIfNFuD6++fuR4c3Qrlagf+l2eZ6ZPGLcPHVwKatV4ezNarLi/8S4slV7t0E4mc
O4RRV77qsD85dppd8y+vZKmgIiEXGcERsQwjQg8AlH/sve67BF1JxLJrcm7jZmNy9kevC00K0/Bw
TmtP8XvHTZjg1ogI27OFkCrvsjXyeYlc+0hNTdj+9tpSHRVpVpYE2uYhVvuQti1Yzemd1U348309
VD1FkUM9nSt3l5U9U6lpn1WVORIymb1bNBauFnN0w/jTXP0vPWm/6kSYVqLkG9o2927hzSwyTS1n
8eNBceD6BIRID7vXoTy4eF1FmhlwCgHQdy9JeKCNP4Pc+sM5JHv1eWzaBMu1QTmSgwnyUJj3zoR0
8pX0ilhDpsr4wM4RHCpJm6K0ZCmQM5E+b5Ytrjp1uaPp9wQTiyqOQEtuFpRqN0HkyJWkXn4P4FU7
y4fmhL5xBVK6l2Q2ssDNn3mIUdAc3K8M9ltxziWyHWj5lee3NmgVZPicw7xx/79KSGYKIxAIkQf1
lMtQPE9V6sjSHL68OTUGTtCm2EYQQO6Gu/TeFsWhctM9toIn5QytwQcbrIy/HuSH+PUbQE6dvsoQ
BAWvqvfgoo7A1eApLHL2naLE3EoDJwbWa3IR6ZMpfdau4BItRGXYDc2QwJHKfO7EvMZ6yFgRP/z1
ykFVz8+qmxMq1XW6abaXo8lCark6QPI6No3hE5sWAOZDrckOjEP4MnWiTVzlOIB2idE5BdE5TDzR
RMRA2vIUyh/egGJfeV6hvQkYYl3DeDcgmt0bCIkZFpXlYgeZp0mMFUSzUOuVhsDNVM+tYCnrVgst
itJUgws7c02BmfmDiWil1h4+XZOE9QhiQj+deJWA6gvrQyWQhvBFnMpfdegeCnVXaOGu9qsO8LVw
zrDIpH4yb27EBw+zI6ya/TthIVdNHcadrvIpmjConifFodxT9X8A26TfgzMMH295gFxOtbyabvkQ
4naI+KPQZNmEhgUmtV6rOAj3hiNuyjM9xAWjaOPfSgaLa+X8wwK5Ojmfd12FA7vTe5d+/1wQpoOA
tjZLc480fncx5s2lkkqAlPmkWTvrPi0VGTA1vmQeX8p7HwBnSY/RFlGcpBEjDryg1UQa9+vilh9U
vF29JQQuQu2nYSdtmDMoqNsunnSVXHx1UFPylCOhBDVMzHD7LxCVTxtNlXEjEqp2P47ZBO+61OiT
DZmTHZZThI+FgtLoEj16tHrpK5DJe50VuaY1rx57IdJto68szT++uHhVto9/OLQBDnKxkew4MoiK
kxT01vHxlcdDvXAxNp8QZw4khzeXboK1lVUgXgJZgij9NBVTQiLlSJnbQwrPdPRNqimvp+GXP/Hh
dGNzUn4Nerpi2A05dsAfeQTltUQOpzKyzlZ9iIHsKvu3FSQ1A7y8P4dPw0uM34gHWKZC2+UGJqJn
FU/SAcvac3Rn/7Vqw7AELQNvExONvZyCC0TXz4VdIuCTIpK5hBolbvz3xZwL4xSCm/sDlscd8QZi
FlB8vG5R4ZPFwA9j5+tfpOKf6jOn1M1AMwDFygeCM8y87cTJOmIJAYrJzGwK6SzB4LNve/wXIiE1
ZVcVQT/NAt+WaI7rDkdUYsXbYO7h6D7w33Z9DFVyRn3m2Ep5peAcMGNNDFnhBP9GPWC+GSnlj/4I
WL2y21aN0BMtKxIlgfhP5GfMaMG3+hausjXpjg2pid3EZ6XI/AsaixXWlNtqZaehTnsn69GQTK6x
/YbdZY+iuTXwysHuESYXXmiqGuYX8TQ1a6oiwhc1Crh1Aglj+RjviuB1TJL5nvKV9SMzdMbI1kYN
csRUxHAm8+cRSAmdlLWqooZdYYEtclLyxmD1FPSOAFcA3iIC/yV1O4ldjkCIUulUewTJ93+NtIrC
fWZ5z5KwhjzeaTw59ITQUiRUm833OhjFYSOkBDCq1MfcoMP2vMSjEN7H+U+mWhOn4YmMRHPrUMqQ
7qQjDZGxApx91w79W8DKb4xB0c65nWQYe8eT/k7ZErYhQHz103a0rhSYDMlC+Ap9NYk5RHnBtlQ5
PzWv6D8THCSZqi1Utm7Ghdp0Gi06O/+C1vOjqB4HAF2z0ccCJHbwgG3FqiLlQW8HUHLr9E+s5+R4
SeuLQXDaGJyseFp4Ck7oBn0b2q1kLyABF956Q6AlAWDOXqkYMOG3/e2hnrBlmV0rujpLl78+KUxq
JUrwamRhe31R5Z9tdA96apGFXKoiuimgQ/kMbGI1IXTIa9VzqzV9BjFHb7gncOshVlwi51hQsJa9
YIqb+PLr9RUtkrPHS6XPN+MUzMLcEThaDUOWYuauMxpHdvSWWtEzCmtOdbxEIkI3NOXU5DMNPl5s
UjmFzXc3T7enso2u2/knXtwrP2V4J+sEsaq8NyJKnqEBnImXQOCkib2nm1ujO8LyoZDZfUcjJbaV
QQXKnOV0c+p5PdC05VOTCrPkOsEgi0hQQuCmW3ItA6Q74SkcpIKfBgIAsEIanB4ldoib8j4Hl2A+
dIJ/wY/vMIlZef/jwDjvIIciZh1rdvSYQ0HffCHReOpi084fBk2p26FpYnT4C8T09AAxLb5zUQv8
+SMEK0QrcfY9I8anElsmwr5mzK/AIz7Y5De8s7kkXavAd31aIZZa3qAt+xKst9wcT1jQWCrweKh1
0sTbdZk0sykMhl2MbuCADYVKrPzAt4Nr79JkApVh07K5Mvg7V5CXXMktZ66gBU0rYCl68a/+a3g/
KmKtXCFDyGUl1O5iyJWnK7syNHL3BCUW0BJKP4BZ6kYnnz26LUDUUcJiIBgOCTc4oVKTA4E9Vgd6
dj14cFXHNwYFkTYaEYiqRi+ki+/XWCK5lY6KgpNvZXxOeXpxyeiFAq4NKfQKzUHnS/qEd3Ul9/0l
m1XI4I4hzZlEpjCCcMlo4uy4Dtjb9712fGTj4z//TfUSxzDUDTQrqLCHdc5n0QHOIDccoxjh6riq
w7gDPUDisRm1u3AOmtsGKVj4U6X4LSrmgpLZ6mUlYEL1muJCjfcwP56PNqoESXoMsRGz3VxtLEOA
y/0WS2uldL0KUz1v31whQvbRg94LufOdpkdfnpHzr69i2IPH27IH3qlbmkq95Zo30WeJYu3+bwLx
CvZYIYizPtDaVNf5yLWOm/eiIBeY62cjDA9ltzObE0d16APG9DGv1HiYBV771ImjUfh0l36ffBsB
x4x3GqoVD0VNnQujTkZYBC1wOFIJI8un0b9cZx2OPW6XFEnydqGMkH3Ajyy7BfGnwBRJaDwSRuVH
oz8vbiGFSGKxnty5/ZanAZ01kgPsQ7Gy3EgpAUK5lPEpgVUFdwg4YdKJiYAM5KfsGUPkqaL10mVw
Z98NMQrT+w2yrrBvPiAiXCABEP2tuuQNkwFRGcEV38kbZOg7/jo/yABEH08/gbvSMb8FHoVMhXSy
o8wUiIFkJ+I8z1Z9vmEztwPxvcxcts4Hisn1YyrWJROc0SUDn0mAQf3YMe4n4EK4t4g+mfVl3Tnx
EzdfO/lz5H1DpGAx5pOvEJVuul0f+ODZj/g6ZqUEJ11sKJ80NNk6pdTKjPm3NA3RuUsbU4crVU+v
iOD0izDdCzDMg1fpoU0dwmG6mbnLm7dQ8RGPuJlwylu/Bk6ssArQm88wvxjKnC+md7c0ivw8JWhl
+J9eR9XdZKtpDBWuLihc547XFz3Ca2DCB3Az0ggwIKbtOqQ0DRmujNjcI70uOa7nkbZ1mT1M5kxx
57DdlUUiiJGEN9Od3nIQuIm7fvlmqsJN0Sz8Mf0k34TwDBF/mP/8zaisLMWo5orv7foFusGuhv7I
L/rVL7zREM2Uoqb/X1vba/+nkobKbBRjzIEhP0DKZ+e8KukLEcfEPTvyw8BOV7wx6c9uhFUPgVoh
Wg5iFruyDR5nHr8pOkp9J61wec+tbvq62yoRUTJSYJ8d0ekvrDcP7W1UvvKZDAz8LPzLR9/efOna
WGD806vffGKlNfv7N3eIAIMFJKigFXYnozKWFWXJIRT4e8b2oifxn+Numsu9sUmH8NhtELInomIu
Dhd80jo+s958+rJspf0rsuYiNhPis/8HTZ2F76ICWP5hJyCHganJlnOMAFCtk5rVXaIDjubbxWRF
9tIH3D3AKkTVnTARebGqhvvkdlu3Hot0f0qgVSqDBcIDp55s7weNTlzpleu7NWZMm46ci1e+c4li
apaIS+jIByzqLilGxazNPO2nrR7q5ZCvcSTu7xkF3yLrjkTa1h2bPa0CrUDXXy1ccHJUxAFqTqzi
prjcDBEHIBGuXJ+EfEc2smjYHeAz07eSQw5ddNp7tIfAUpFWbGosCZpedoPi9FIYsQ0kaqyO1sWs
Ps59rwE4GpCXUYD9cssEyfGHrr7A/bIkSHsKRibBPvHZoRaqTYKQuowZdaCuuxlxoZax8AMN1G1J
Df4cvqJ0bsF2MBQs7r5g1WqZAyCNIcuaMEbfFHJDFq31gtW7UMbKz1ZjxIUnC0PutN6QBfc3+sbM
PN3JMnZCKKuBvHzv1Z2fHrwiJ2eQN9u10GKQP6ktzqnnmcXk8B3RpCgoOnWgHpT4uwYr/XNM+/s1
JxENuV3q77HHRAU6EvYr0yBJD6uk8Kt41dQ0xmKUDIbqLAIMchrJA+WN1I6ToS/gb5S0bV6MBPqX
2shKH+xMvCpGLqmqaXUCwIGfYO+29strxBuA+TDj4QruDdSL7lMrKOxh8X7JTI19khDYHb1j/Pwl
K2p4ea6HyucFoxs7rHqEmAq/7O7Uta+etd5iACQ90Ens8Px81bfoUy6hQFLGxZLjWm+NtrpCy9Ov
9QgpqSkHRQHzgn+0xQv/JeE5ZVMkCfiaKsqUxWBpugKr6v3fiiFn94ouBXpPC52VMLUAN3LQjzXX
1i2/mRNEOxrUAcIZsY6xh+Vq/xX09FM1Uhi615+WuDUnnJmbdQWs4sbPoyrWJQ6N8idi7MD1r35w
NJ+IYA+RznAKxDAJMLKL3uL5gL4V74eW/+b6USeZ7f09XL39w0S/+Vo0OBux57+KNqYM3yYcaJnC
Wl1+2Y8raQvp8vZ867AsVdg3BxWgFGsbPJZq+2cApYuPgHltWjE4CNhCVYqMZrzSLn0Jvjo/FXog
Z0x5RPx55hGgjod9Q9o9MC0+sV37N+OA3rrJjFxu+CIzTbWPsvFd4YoL9nXhWGhQRI/05wqZf2dx
/3P0VCyLu2GUAwvjSvPY1DGbqmEBI/eEbR/6wK+cHdOLlD6trsiD4CPTTOEStEuRisJKb8ZEcJVh
hgdaYBCs1fHUo1YCkm/bcrrzuflGbJ+6se+Zwd/LZlNGXf/fNTRSGBm4mLXNA+tUGwDUbEBWa9hc
uvOE8Pmz0uqD3YcaSe96Yh9QvEK4iyjW/aJJlvk8e3hIJEc1hi2CZhgym1nuePYrbCv0/HQrx0Xq
+W9cHHo9ivSinZqAuOdAfbFRfB9mrH7Vj9aqkWuAWbkKTvYi7MUdaw0pO1uIpOmHFXxaeaNfeOCc
2D4eu/5Q9K9y1b1cNp6ZTvKBzCwUTCCxcA6+0Q68k/pgQFBcylh4kpBNb0GoqZmiZ2NeHgF04R4A
chXACDBD/KvsOWLLarlm9liUuH/V6yQnL3zd2xXKh52yN/2Ra6CWeXbB6eczb6q7aex2TUYpWEVq
0YuRA6+Lb6y4l1A2VMVGCJqMt7KhtsCQUHqFv+uYGMKt1ZwCoDUe0LpNSqmYFydq36jtmsKdJliE
DvQWYPlwZW7gQ1mEbMCR+XX4m5Ya7Q1CiunQTQzLkMlZ/9c4P1UipVvtKirEFpgY3HCw+AmMsJ1r
baPk7EsH8Saw0yf7IMXJ53o3p2PCOrJZlfmb+ajVIytdsAZcoMG0muWrth6niMTmoIRt5rn2gv8e
iU2MZOkmq+v+pvI1uI7YY91frlBmQ4AKdQkdOaRi4RBjeY/HsGFyB6AP2oCt+olV6qhC0TgjOmcr
/9uJR0bQOfpIHJ569QZh3vv3IqiDGrDHsFbnSsH7J+9aijZ1b1adj7IrsImcWHc8dcHhB6RXCz25
I3RmsmD2T8OfGwYzYb2VLLnk8H3DCvDNYCDoQ7FK6FB03xeYvjd1MQWI20UqsYIP42kUf992/DTp
ThTt9sv4RUhneAFjhkorhoOqaEeA4OB+PLTMvqRgF0Od1aqe/qbhX4PKeDpNI/8qcyC3MORV3KBK
C9D6ePkk0J9qQoIE5ur0RjamZKawZ6L+iKlHTYA+/ppJqCXpZdqgIolWRctDUyS23ZXfImB+Xvux
U41MfVdEciBX7Svme+WF/C68cEpwjGbHwSmX3ZLTtLnZrlfkUhJPZXhxgcVL7NugGfqW8/Jt5dQg
soptnp+eOmDseIRsZvv5RnopJirACszDiodsBZI4B3paeMaaWS3pE+LbkBB2xlwQSgsiVFOeDI8y
hHhAX3o9zWOVuBjx8Eymshz7eBlGu3wWDXlUxF6J1yXZ1jlfEmYNGyXutRvhjOBunXED4zxMdmCK
lc3wHsBvJcWZrvLVPhooHLFqC5EZEhULEYlIAEKmFFSt7YUa/5zViA5zHAp+0wdUgVfzcDFK2IC8
dRVqVUt9p0sb625MHUtZXeqXeBlHLSBv7FggwwKQxeSl6aK2OSQlYmu8NY47dWUy38iwt4gXA73M
F+cB22A2+4v26oY/ZjdoU08TlhQQooBMGvjneJMmfgK+hEaNdR5iH5NIdXmPnJ5pZltxTJcN4/ag
3NRnaLMEGLzEqqfCVc+/qd8IwSvORsf6EyRo2WJqjVH2zmvJXFJItweYLRjgQeALWXZ8z8CAtaeA
N/qZvmAtJaMW/u3TaAdremWtjTk3GRX6nAAhkXO1WMKpANeHjKEnd2pEvbl3/dqqsNc8+xw+gkfF
3KbeAVwN7j04hFf3gVypcKbSCeQ5f9JqkVmxmOG+4iFiKIxJAfA3CNVcQ2ZENaE773cfMMKvOUBL
kHyLwKQax1anShI//uABmDqxHZ8ii/MSV8De5q8vdnzOMID/2K9Q1PUzIGe4DY28/4/FMxmkRe9O
TiMkyDPyYPn9u+N0YewnMtl+bvlmwH6wGtFvb+0QJkJ/a/XlmjOcJHVOZl+vZHaqEoKH7gqSSFJ6
tiThyjoicfkXOFXQIEiHEzmAbHkxdvLs/DoOVRh7vmekwngM7h/ijkJp/emWIqWjqC7k+SoKD5hb
cnaWPSci95WaclIeVunUVDWrt3zWh0mBE9y+nT61k4bXZUwVn5IMQMGTx7Y7BTdVWaAKKX1YANWY
a5YTZsZoQjMgVLtNCE4o/SoZHH7SZiFGOayS6FWLd1K69PCyrq2GcBC3qsrc0JHI9eHjp3nkS+80
ECI9p8qRCHljT5RoAw2SX6BdnJ08zOGR2E6Kovki9XjPDTtaG9X7c5UHk9dPTyxlFyw6AYhRtH4n
yLvJ/H419j6M84q4BHrcIk1+tJQi477dxvHYjUe1AicDD1CnwybM/Xk1P8vQRdiagsZTVZ6N/tem
sXAIwIKkJnTK/lE2tXLDnnl0gzjCeEH/b/TMxUPyJSbHrG42ZiCv/VIWTotv8A7o5jKPfURIW714
ZTs1Zl5dA0E9VkELKr9wj2nHjau16UZKz6paZHnjStfR4BXWA8aVdtQUp2X1Pn7hIlmDA3BEUHga
OmD8q6INpYfQ/HxrJ/UISwkTljrkOTJ2SDBvNiYrIpajUpKyG8gMs+V5K8zX5TJUuPDzFy7We9Bd
slqSQQ0PVgCCDF1HlC1s7lQpFGNRB/AsM0JGbZiPAwqFPXtix/f8fKd/D1txkaHiqaxyVQLfeWLM
UWMzSa90/Ldru5Kx5qMYGuLmdTj0ffXl5NxMpb2WbzqRccNnnpm6bLtgo3dBizpICAgPxh8qqhUl
fNJReRgUbGM60jd09MHZxkSSMxkqCMzUr/ykZ/E4eFCraTV4GlEZ5s/R/MhZQZt/eT151R0gpixa
cMxCus6Dt/u9v1FZaoDh1tCzSt/zWr0eEuq5YEwO+DJ7ToIGRFJsFY8FwdESm7FTbdWRKYhHE934
vJRClt04GKaKMgmqDQCOE/IFFJcCDwndNRTyrF6M9tpZJ1UGu0Hcx9L8Dxy1RikFfRD6+cFSpx3H
tfTD6MJr+7Onfv7elnUOX7Eadw5fCrWUeHigNCR70WNtwaGd3PdmOCCM0EGkKPGF95nsZR/zxEcU
B9N1fcvdLN+ygMx5/wZ9IboU2ySdPl4BS0bZg2h5TZraicxBkbGl2Uer46V0p7sY6AILH/4sgOCw
ZXJ36P2QrZKX/X5qjn5KTUkQAX/gJov5g6n5D0SijzWirX2KAQXRvfL0LKw9Ob+RPDUA/wr8FY84
2snTTzJNTjohKi2JYcbG1tv1VCg9Ql/nYCtsf7MPrwSZpqeaw/tT6vw8dkvZgJoSaZzVz0IAhPC1
6g0V4P3FFcr9ylePyhEh51jwM/q2zjAgERdE2QaxIKhz0OQL5rsFoPgeA5XqgM5WXK8fXjyFVlSN
jUY6JTx6Jd35Fibd8i7JvCJvEVm+DJ+5l2nN82/i6e1uU3JQOtyFD/dpTt+8XKdKiwlwhVFwQELQ
w49R60rMP3DlYIwtThnISPv1adygVhXczapSoUnVDRax/AdnLtPDlvHFgLuc4puEKmtoGfg9JQmU
8DbGWiWIIhtLZoVbru/ABZ32h7O7dXm0FGk7QOsaSZT1aIZL8dIAO6X5zMXhUneHxi912QHre3Iq
rLeC2GC1ZfI56qvIXQPlZISk2yWPezBOcLPsTY6dn7bht7C7eB2ZA2m4IzGkhcsI2P4H7BSXr9rY
s856q4xJSlYUjtMP5HjP0FkoCixVS4pUaP7qiP2yA2j7tivyzAUXnbcyfZSHBNWKGH2hLb179X28
gjAlvp5R88cbInW1ThACIoYoCrDl+Gcag1uiQgKgwu/jRNq0Kgxx0UvvmuTIIXnSyo/Q1apuYj5T
8a+l4VaEEQF17rz5XXwhw5v0rJQrDt3g+B3RLzKjz5nOgdVaOTUtc1r9QSh4vzh9YfZkkZOukyKU
POofdp2oRe3ZF+AUMPC9AIg34CWNLZRZManjFFrjA3ZhUR5xkiryE3Mlpngpc5zYn6/SvT5zYBfe
+l6e6hh2zj70DISwAKFWc43+LYdqI9BRgDSiz2WyC0Mt46wRMbsb61q6x8Lecz/Vt5zMGfp7sHvB
ALKeIVvBqLc+tsCNTxPpWjb2yFWSBMMT7hC6hSSVDnfJhvfb1EWiNMViiHxfY3lmAFbxmaFgJJwZ
HWmMmX5Iibgmqo6IV3FQD5D9OjswUbeAJw8LlcpK+cNX1KH54r953LndWDtTJbNx/JxHCiUCtdUR
oxvRKeu+mIUjGBuXWlp0bGrxszjKmzeJFZPqDkwmWzIQqdF3qvksbNyxreMcmXWSgZ5Jaw5nGky7
o8KkD9NetVwG4TBsr40usEuVHR13QCkD/bY1ZguP1IUcGfAHQXwXXAMCsX2KDkSpaS5LIQjfSTb2
SxXGgIHJ/36nR60YTTWNjy3Ltv8gy8vMB+3L961rxXIsjCfR1+KX2JZ8KNZDcfZHO44OQKGOnf/B
O5/GiuT9qBFFOfI60OmxL3SG/uGzGHxXdzqghsv3ZCn++BHFUZHT9XCh94lj4l2qamS+Kd1MCkoL
A+si8aoclo+26sCs++NjwFwASOzPQtOEJG26JdGfBshGApZfmAHrlRuW/q017Q5UBmelfS31bGGw
bHvJwoJk8ew5mDtG3pirq/Clv93sd8BHS00Vcvgw824ksaw6MqEHMyysg+bJKYV45n+S8hJoHRxS
mUaIqmtLRpOKmN3SnmLl9hW10U4awgaFv8PB9xSyyjCqHUMiu6X9mUyGxmqppUrc/WITIx2MYNhk
X3ajy5dOvRNvv3C+kVm1aI0Y9Z3QVjxc40tJ54LTG0+Y00JmEZok0xu70DvjISXNisYmJvi+1KhK
gCkMXIqjl4FBHkETusmA2uEEoiAe3PM65rkCb/yu9dcdTgvV7ID77MP4wGPGNSN5EmmNT+ojqUg/
/gQW7LQsiiBb86EcbrDa/xBWXYqfIi9MvBHgZT9qbgZuazeF16IxEYQ3Y7sfSNMMr7rXmFVTeVoZ
Kfr1E7YpPIjYixCOS+aqOPIz3eOTh1J9egekgb40DkkbpwUe/iyItmJKFoS0n5gdXkBL6kncfHAM
FUPcZD5LFFSnWdBudBd/7qgj9mmSHj5VDoqhIEzGwMFH2Fpn3+I8txwMmJ6U5wTWBKWi9Lnsqyev
XAE1zbvtBtcjPvGbTmhDbfixxYUpm3nYAjqLTw/k9EL5h2QXlD4QwVVp9/vILKcSBrs/pjizFlZf
yox89jTj07ppKjDdT7ZQxb0ZvDIh1eED6XxkOlb8Lm372V6xScta13rhI/7pLw02mKhY1DIXDdfI
im7WEKlzihSTV29An+KpiGD2xqTVnqTJ3LZpST93HtKPlRwkOAJZAvEv8wyIjZKmjjd+UZ7QvL7A
EUMI8MhRKY9fwDUl8Oe/eTNIfiH49uHL3KJqYgfuOVC4sF/QjkEtq7n5c31tHP6hhNkvIl4+j5u/
0usWJJCgYWX8PYF4ESrgsEDdW2NhmWyaI6FDJHhK2gYpslpys7vSIRp0gpSgRDqFsM2gOXFYBosT
ehZdbD5f+3ItV7LmQsLL/JCSVgTYXkLPemb3YHX1cq5LOf5EimHDa1MgxOktDugjSn/uX2a5SIMZ
6hR3VGCIQTih+A2FgWaAsHGKFrmkx5OBzmUybnB7mGL0IhBLV+co6J1rG95FUeFMNhL0kuoyVA8U
llB07hHhBKNHxRI1Mnz2mSv6Ss+7TTRu8LdX6APlIHa8fkl8WT4WuxTWGNcSNGOC+owWfDbREZ+b
6ftsOJIR8SEqvIxhmVUOpFh+H6/uHgROTEDE/M2RjjHBChUB1JcmiavXCXSK5CLyyKEnmI7bMLhw
Crrpoe0x5+pb4LdHuH7zdCPEXVpsZjah/wnNV0ScIYpZThaN3kekQbzcOEx0kIx2pDqpNluDUVVI
aL/saZfB+34JhnHA7Joz7+MvORHS7RsD3WuMf1swfy+Xwt73kv1++iLjRjZ732EDq5d8Uu7Yy7yz
390WBZAeAMN5oD4Bo2rTKIVcjJP68jWZfdL7JghRX3qWmXCgAv2jri7cR9EbHG/kvIUBxlsUD8yJ
T/LnuFl7rQArmxCW/Z1n4oz7TrGHeHX0JnxicsF6X93BOttGvV4N34mhzfOm/uPBLb4CjD8Olo5C
Clw3LJwwWSxy+uQkLh4j5boarsNa3oA97sd1fEVZGG+nUxb0IjofVDfP4mfdCCquM00MT/MZEAq2
7ByJ9LMfY8wozNEOeAor5pSvm6AUxpnIpj3EfVMPcY66TKQXYOYEzEOF52xOSQTyOpOW0E4Q6Cf8
9+l/uMhv6uEV49lE9eSTyRl8eiRZ8BTEzWjTjrfX8NuhYIIFJmeD8c7qIRMvRdK/2PTqRFeGq+qw
bv8wn4GJZGHxcrRANk+lKh2OE3IdRDzvYBKWDV8edDEQtX+HHfuhGFkSx5I8lgL3o18byLdkmOxb
Z3RUX8778Olx7QjUcLY7BbO1uhVr1grPQERitylXm6BSQUxfkbXO42tuKCjIAWYPcoGZJqz3U/5j
vNsj9wkB2tWkItUBHHJJL/snxpFPmzIRH9b1QLNDMYToQFevTmOab6zIuMsoZRdz6Hpexg7wSjus
2LoBcmu9MP8RdelJ+03dtyQQTYuJZ0ezxOBoapTDtF2ke0L25EjhmT4uKDyoEvHqlqLRq/XBx7mq
+YT3EwNyb826+Ze0RkPvhk7qFz67gEqS5ExgR9PHKhGV/8EIUKQPevWA6okz8XyRnyxQP+y9w4Qx
91O/GkVV2Qo3QLQ3/GPZIJltmhp/Q3zO2gnQkyrpMNL+3T6Fukqk8RZYfXTjYRCX0QpGYzrW3nVU
CzYkXEZllYihsLiFt3DW7rgIEhIK6Mo4a4d0/OK9VeePVa0+1YInivTaPTS8QObvQ/HqqttBrx7W
BFkVQehP0SUGol5OrCJQwrWFW7qD0+dasoVLyETEqDMDRNeviygtkMUIK2N0s7wwPpE6UNuIVTeW
hOnf7WymJZtPAwXrcFrXR6Fw4i8fA3hAG9f+B5L0UltYjLodkofsLZ7fuZ+35qR5If+RXMxZYAAQ
e+hM+tXriPy2cy37sXaPfz6JbIFhXuilrsy+d2YMBXzjPoTQjda82VMotPuQuHE7lXnIXci9kjT5
I3ln8IMbr3DiJ5IPGvXwytHjlC5bZ2Vu9fJLAZX831XJeh8aHoSB6AD6HJkJMY9v/6D0t4eG+j5Y
86YXlUFRn9Vvqo5NYjK2ywHDP9tI91LeH7CSligHDVTJgQQ7h4LqQ8cU9UYMSIEsaAlyyeWwws/u
f5frFDl7AgSl8W2BsAL3UZXSloHFL2S/ThOnZ51zRC9Pb2llbRycOu3MXqUEkg19mgwHjwKiNnRx
qIvRtprORKZrlhn+mk1Szd5eBQuGZArHIZAWF5fJ8i0nOiwvwEdp0oU0TQfz3MIV6E4SKaM8g/y5
l4uIpMNGoCk7t4i4AqZxbQMXBZFDYsYye4UU+kC41Yb1rnVabLnhWSaGxXrPSzY3ErLQBaPfuUMY
Fxggk0Yp5689F362zUwl2wpToQHCY7ePuiKg3RCh/LTLIaftFKbcXwYxNbMDGRbassMyytkzU0Mb
mE2/I4bi359n1iHPyz2giQTu9DMxWKPVc/G1+GM3230MV+lhreuDrlAT9IeE/HBe2YxwSZJ+dfWD
MhtJbpcyv957ykPL+U6P+asraIJv1rbX7yAjzg2g5tyM/G07Ts/IXHs7Qql0GbEdkXS8ZIsgux0t
1FbhQnLXmAiBcsHX1LNgg4QVCE8C2LZaPD/5aiZITQGT3a/VvLU5uY9LbYyUrQyLx86etH9emV2J
6NRzPsO01QEsiRKKHbVoNicgpaum11KCquhdkLT7YgYQdl2FyBThAo8P0fqSIsv9cpmJy30GVg9I
1gYCtYTRt5Aphemj6Hrb0+fksc2UDlVbGSl3Fc75Q/+YKftFOlY2rdypLmJVMOvBbMvqJgyQEptt
vY1RtFKSi9y7HnkofLwfeAmv1wdmWuvKbimF+LnE63cpVPAILTD2pULGMeeVwWlcUV1vz/ExIn5v
QmuJQnSGGHp8oVcOeArOr+zKsypuNSxVWyTN/I+iIOWWZGMNrsDQN8zv6qwvt7sgD/0ruLPJC7OM
Squf6Qa620v3Wy2BokpHNRn/k/NvcOp4Lyp2BRzWGCktbvLohX0wV62nEMz1p/nyZhvC0imawSve
PES1elbES1GCI4Ngq09gEzpk1eszsh4m5GCVs5vbP/2PUwIc0V6NpIqUvnTuwEB0ElqHXAl1MR9W
Suqi++xO1OVg+GZtMjnJg5U92pCgLiIiQEszT4vE4RJZJAQ3Tic59aco/t+c77tn0I3dN18e+QBP
XUT+x1S3u37++gJ4y+06Oo55lgK2wgiC9v53QGB/jRUsCuCgsC/xZRvdUIIGkkYiNIVEdAQDiCJ3
33Vn6b/mETYQYsIe1ZnoFKRH5Lqd0AOecgKWe9MLMkpVWcZWkfRZGUMAlTmWXFeaFwt+5g+ZDx3D
rZaWsh7Tqk8/kvkj8x3Zr3r2Js0b/xLlUk7vuDb7kAf6lRhR4Rk3zr/IfQr8tFfSBOisG/m2pbPt
+KrK3Lknj3+4FH3JPoOu0fDrxOJErKua6xt0fGhNey7IbZ7pv6dwSP0OCHPI45wBUPQk8PBLfJO7
Px1duaq57hcD3VIVggkBS64E6a24baHPwyDl9Hdcj+peVTauvivhsuO2BPG75i+LiYBULA36gHvn
Yy23Jz979k10kTvSpZp8WmyJu3jcSjJVxwv3V7/6a8NEWIGaCda1zgBA5BFP9EoxUlWfF2D/+EIF
WTQwX3t2Xgxpn/ekihVgbuNiqcO/RiWcK9zIxlUILhtKKksmhC2CfD+OyBYwZwDPef8oH6Nbt8dF
cOBW5B6zEdbtzCBgLIIP+lf/zshO9fDjrrkH9M/nqp5dYdZMtTi1nFUAwLdKWyReAqYOlD2dQFzx
d4KWtQcnB+bYkqHVs30uCwEXhKoGNc9eeIymVsDtFnD2uwby087jNUCevYDAMAFc1gPgYsYWZERm
ZEFEksOHO6SIvNghGbvN5abF5ozbo84eazDHjPs4Prc+jtwErHR86GcU8FjujHz6fommDAW3e0YY
Dtkn7gvjfX7p3uE1Yfod06vQXkvf4rgplmwnLCAV5bhNQd5EVqjtRCm4yqlHb5+JX7WwYYVjDEJO
/GZRyNwksVcCTFjKYuzSemtoV2vhsMqr/P7QfusplwDwyQRIZlJBz/znw2JdPGhR8u5N9g/9MHW6
KTobdry26ZbvJ5gdcoSdci8/H6jtbIGHL1EyulxkPv3mbj67ZHogajE/Y4UK8nKHu3L/IaBmOoFo
hxgRa+0klWYxpgciNIMS01F28VYw86vg75HV3DFcGHpOO0tst99tj8TZxHFog+3aYnIJMSncQNAH
msk+4dqvXHLdggmfl8jrJpQtwThLEOHkr2ClIMy1UAys9p9688t4MmD9JQfxKbpQXYdr08XTlaVO
t6XfBjQ3hAvR4BGeweqCQpgRed+wasMji7BfAiPjJcRKVB79kZnwLPoeiy9T40C1ggnz2gw5/WgB
UmrTBZeKC/qluP39zMtVwIId4AJ/ttkiwUeRwUJ11Ct73SqpZ4KDt06NPSmmDpI+GRzs/5GaAuzo
YFjyP0oeP5W1Lm7GSCWK94J1xntIJCJJ8tIusCiBIIfz9kJ6WBBx+BzhuXycSi6lQk7MOpvJVe9H
mC/rqpJ5ECVcfuBmf6vUE1RijYrQibWvnK1kfPnu/O/krXfOL21AEB7oZ5sdvBWZ5s+nNgF/XuNl
uuTuDWs2qNoJQJUOSTJjXSAR6MZwZmIEGycAKdHwJ//HfCYy5bHEXORehz92dF3tbjF4EczRdAkP
Q2G5KAJjdIJWl8uBFKMvLUgGwTtm4slPNME6Q4LZ969M/lbbC3QBY1yqNnidIaRP29tFBuf0dKqv
pQgvBvOEn0v2DIf6Ymlj0bH8L7Bm3n1I3vOj/yFF+7hvH7dYDaEcYdUNwW5W3iZ86UQOjQlXwq5a
cPveV1rKZicrY+d2gvnkF3LUql6qOTPITfFx9ms+U4Fn5a1/wlQn+9ctqDM/EnoK4DhsDbI0ks0T
0OQookm9MvF6YetK4FK7nPPGj94H+CTBnD8A3AJLmnsHGnEjRtO95jmaEU+0FbpREdO9NIBEj3XD
NuK1Joq+G73pngV9uysTjbJcsX3n2afcwAx5S0o7xeIyt2LxX+dFhb405BEfPzob+jNVtroZfZih
ierI0zbM2vBJo65uPxeGXp0kSUytBPPolNVTOEDYJ+NzY0Q/HvVVyog22WrNBd7bdcAfMlGMMjIK
eCoK9ipXHDu/LSclhUhY8ozBz0SBS/gnIeVTKKnG3e0J+9ckhHDz0bpjPFCQdR9oXWTviqVZQ0T2
TBxQPPLwOBp1urRTARCSJaEHgpXJT230PVpdvQo7dekvTGreKvIMtfZA+QMN8Zs4C3RXiUapp0Rb
Sza0uHoNLJXVJ7sCtoLGrRbJVxtnLfg0EQ28BuL8cN0lF+Rw5pVBsO7+0kGK/M2XE5yG+WCtMsNi
qn9xy7KiN1d807Eo9srfqQu5bDp3lAulapCuZQ/Vw3uB/x3mS2Npu+7MRXMwrRQ1QG4/aiOYOMWI
eLSognSfiHrafiv9lOBXEKDJql67dzxWGe5JYFY9ReRsEdj7048wvuCAbMUQhi/qisXk3/ItErKd
38vxpI3dKlPpeh5ERCw/gOErqG+us50Lz5/RWn+0iXOhRPneZqtRUURwA+nltUvvLN1fG33/evpS
3kAO95OO+a59pfg6ZEQPxBFFJxLdPXjbibzQOHVKTp7ymf44CAYfovOxkYvYMog5tHylZ08lsDd0
qkcIkytKMbbJEJ987uwrUaJ+L8xuvl2Vfuadu0OTCYn0lIA8M3gaWVKgYnm8Ck7WGb/PS/rrz0MD
6w881lirApSE+fJU9SuIi2KHtGHkD3DpG8X2LDQENRNtiit65S8zELPzThS10iGF/deqvvRFm878
hpawplh0+a5taSDYcakots4XC2JbZEVdsmmDu9WNbMz0dsWkE/HZlHDxEFQ4aICBjkODpcw2a6iu
nUh0o4Q+uNL6WhLCqcbjYr+jrmkUtPSReyR19DtRgq4sSh792dnxk7Ka5WXVeY6rUTytwwjNjw6K
NeHmFZNIigZuIARIjQ7GGr66ADxe5Q73voI/5Hf6LHDRnNqJM4MCMCULfUgY+MtZHpkwRdtrbwR+
7uqlN9LINTFLKSoRxryU9qlFCzoaNn7wpoAB5TAhl20rCPePw9sF+i8MFl8e22wMfeypASbc7M/j
HcdEmM/5n8jZ6CWb8XrSik6VVozgrheQkysO7Xg1yaFjqD1qxdkoKWYqf6zLfE4MI19LvK8U2L4M
NFIgBInOnpzj+DYwZ/Wp+RijhiHIDw8kSrOuh1DUkPD2LZ5s+hHlRhf3bGSkvNTruprbCgMgsiwd
5tzTVyyIQkBUmengv0WeFm8/gAXFdN0xwlijFguoqUVxS0j/JlM/wpRxWL4QQ1CIgeIXvV7ku/Ri
BKUw0NNYhhz7AyK/+T+sMLby31zYhXsHBKHZFuom/85Tot5oR68+s52uUhB6/5CHtCGC3XMV/Wp6
WP0IoxQgwnCeQ2Ewjz4BwBm2AN3Gv3goeGlybQy5TEpTB55qEicZYTm0X9nPhtiR2gcz/uoY/M0W
SOHBhqGkrrk1vRKRu6HyuXw/pEfyxvS9As2nVRELqjKvy7mp0FJaGsHf6MvW4iprhWc9M7SEYWfr
/tsWYSdgoSvHlPXrdqTQDqdfFiSB6/L/16R647MpWFzflkYIcEgx4swkjkMmvofWQD0h641r7NmU
W0TIt++wrnMZSZDmebVsynNKwctp7SqYb45S7QEfwFk0bdB1I6W2RT1MHzVXF2ViwRo9Jwfqu0kS
caiKSaSk9e8J45WL+WYGWZdE6vDR80Z63e21SJx2Awk0d3lYuHz2R8EFuOkEXHkYuZrEwW9FaZcC
mLzS+dlB1xsEjPS2QDtv9hpb5ECFxPZ5swcmbheH7IYoPP/VZMetKKVHq8MIIwYaWMxCkRTxoW0g
6dcbu+XJuxnGfEQOqhWKeRIXDl1+HPSq+e/q9NEw3XzlfjgaLQyfeiC5fhKzWII9a4sy2Ndlypq7
d/NkAy254MHgKMw8fyzu1ebgOc/9HLp9OBdOSVRhfUAEUH/FwUxI+u/oXuulv/NMb/nlqDXvj/kL
HAzg+ujjwhN2GWXJgB+Nw0U0wT7JzNXAW5Hne0VC1f38dks8dyN3aomm9rIgWfkO67aYMbPO+ddG
iHs5YVjQ7tamrFVsdmqmvsoOQP+BeOzCuqXuLkYTKqqhv3xsuAPzoOC0R8DJmGPAoQBEQvZ6YxVP
qA6mNmAGZeTaGQkb6Obo1/C4GIPGUO6m3KnpXQz+hDZ57TmYBW9vvs2IpTowdsOVRsYqV134lwIX
K1V0y27LhziFj5vtBmnrqQTz3ulRTZxYAoNTdHeRVKtjra74zhJDYij7fxjqwjNHXMKr3SlffF0y
17Dc8wBbCOgufZ/AyOITwB3XKstmsDQsL24brzMy5OgC53hNozJ9acH83cTYwcXQrccVxk7VcUGl
UvkXpN0StnunCt0ErCfWtCCW4/2YpCZ7L2zpKpDlyYvHl/qqy83Te846wUtQHDi2/oUS6xavo71A
7XOwi12mhz/UuouT8L7VzAgDMG51rqsUrP3LBaNeWXQZ/DbKYTuTN6KhEuYbKtd/ksRqv4iSLozl
BmK/JC03JLK1SlZapO9iFUODfF4A2y1gYAKyTpEyD3f4dYRxCYPgf6RqR2lUflqsS5IkYpjjc2yf
VvSFBF7xFHvS9DV/t9Bj9qtXf2DdkX/Y+FZqBlEdJv4VeITdPWQX74XE+MUAmu/OTGu8IsIaui+G
00cfJoKNsZFnvkvCaEvi2zA8pjZY6xXOkQNs5DRxx2B4pJsMRCCW82+cK9Pjara960ex996Y806M
S3l2jZH+Sb4bUogl4zRW7tGvxSnDJDZr8d/y20mwy74r15FGbL1+ulEPtXektwprOMaPP+gYohF1
pLmHj423KHlSdsFhpI6xuCIYnVKvpQfhG85YfzTgK3814sRKWYgSg+qM4mTDuzFqDJFIBoP/ZJcH
krfBomVSxU6jsTAr35MzW5PcUJtMg6dNN874kaKuNR7/joLylvwaPYFNvCwrlj72KnIzSUy/cfBf
oSqwGxPjOezTA3S7x9YBkIxvAoYIHKP0gGHIuFKFqCfOA3nikts9A/q4apiziVfcVMhX1qn8BL0H
wrYBDPSsB+pfZIusYaWu6V964bgggVWnrukqo0JZCf2Vnx4wRPhaP3Bpecb4NonHu3O6lCZbJzh8
6O3IQJaLn9pWreDyrfav3qLuYAP7tbUWjLJis8mv5rYk49SQS3Cl62uwNT28iQu+TpUuJ4n0AGJ9
f51IQbixF3rRqsmD62IqhaX3CapWV2mOu+4ewJZyQZiDYzIamhAEBqBMiY6MVHJnPT7WTpn+06F5
/ZhXn2z8rOINCEuHZFiwNuKd+ZR71IMrCvmxaWvg+0glDzaT1spZeJx9n+SPStKS8qJJZypuTkgz
Ai1JZxh1B3WuGZgfYwOyLIHDtJ+2e3JF+lo2mVtSnmANQC3R14Yzp0kf6cN8HAgPJfomSoWQ9YuT
IZSZ4Sabh+t8aX1prkGCDnA3odyWdHbuTny02yLrjWhPnBqzCwI9IbqIyI1mu7XbVyWsPX5Up6Jd
r+sufJKVSwfBW1svLKbOEmj9y3Y2O5DeMET1l8moRnRqoNtQ5vnjpwqtBu9XrSgEC701MMAdK9pC
IR5ExFcXd2kI9R5Y9tXQjVFQSxY8ElTAuvEc2az8rkI0pymZaqENiajSv3xWfUFOJvN21SOde9lD
ek6+/gEi71Sg/hU7VF1XJ8gL9Jeloij3e7sUj7JjvXbkXGpBdXLlMPRH9gAjTrPBnhhhB06r5ZWd
XqjzrT5fnolwB2BrNBo/er1ZhZwXYqlcbGH8V3oNSC0hgiJPkCy72YAI3f2a4x5ncvG7HXd/EmFu
RmWjYCKFfqTKNX2mIEz3XzRaTC0Xd61bWhyRqTmVf2rIeJ6tR83dxY8FhLy4BQPkgNECiAjD9jhC
uNoM6biKMMhmK0pWwafvY5v97hSl0EkE1YRebp4e+frOr/FOA5D0a2dxy0T/eSP2e7n0oheCm/eZ
zdv2ThcV5RPAcoAa95hvpeHuVdQtEylN9hjeFz/j7jjCIY3QVTMvBPg6TAM7b5/mje8T4N1KzHPi
6E5Fl1qiLVFTH8d6a+BtxFgVYGBh9rNJtghJJp0pINq7+qAN7glXkJxVeQSzCLiJQr+CIF94WmHl
67UGyUuY6MQbcGpzoPbPgrC9XPhluR+t3djJ7WvvKShxGqoACPXG44sk7KnaUPXYCVRnx3U8SQIL
E0BREZJvzTZjShlSAdvgYpAeZs6HOWsI9uBVTSApW0OkAMsLrUHidi3xNCSIBwWCEVG2KA+P70rz
G+DaUlWQYKRNx9mc6Sqxzgg4k288o2EXbq5xdzKXnuxWIqMFlNMRBsnWVgMXO1MJPtp902Smt40e
1dYupiipB0NIUX0bzt71SFUywUd41wmNcZwOcvWcoFLcALgvIZ9wL4zb7QY/P8hdGfL3poXKfqbv
z2PfUhKBlY5bdtbRn6ioDkz1AnO7IS4iclOKDORf2NAQw22wYC8vN1pYy77I+HMAPX+j7Ff87kcy
BcvDyCIffUv3qfVpL2eB1N74Y+m6tyeXawjSKt/WDn++fBJH+QQsp1XtTtbrEAYRDtGbFdoOxJNT
MHzLpyfU3Z9XzH4+gfvTiMSxgyWolvRl05OjsPF/l39nzKYuFifyoQFQbWNs/TNLwWzLiCZQcDBB
N7aI8BfON4PJ4uafIjBCU1dIns1XKnSTX3sl0XT76rPf/qaMDhs6jROfurp07bFgKtcvrxoJPO18
CnYPmtCtSp0VBI4uxn8BQ1reLhODluqT1bupBlUoh0yKO9K6BGdzkVmu76G25wPfZWoQBflw4Gfc
yOH/hM+h0OUJFXNVO5eAxef1KBcWLMuzVSm88h1+kP6HiW53d1yFEdeON/DYDCcfcRazj0mcFw21
KpaQxz/lAxeQFmW3gFwZmRm8hvIFTBbPDI0PuAoWoivxSYhndJOraKJ0YssLcvgng9YaFxg5Ioaj
BBv85UHSFICd66WkUe8PaHlyh+3feJeQfdjzqTgQesPkg/CKVrWxao9XV/Mo39OcrTSrWARW/TqA
7mVcSynNehMexhAUA8JiWHQ/sDV8s/el1wChBM8zZcqqdnC5eGoVyWfEN+kS2qMfVXrE8euSf/RM
PWEfNitMFKDxNgB3N0F419r082E4X+qMWHUglb0q8KY0oeQUxEavbOU8JssW8B+WjKuWR8+2YZ/y
TeXASf4VeRwShUBtrU1q4v/PAohk9Y5jsjomvn0R5Q6dNKZxHNsoxetCPczW28amE3T9/8cTi+6U
w3Y7x1BaGYSxEKfJB2lPZWO8UHGWTmann6pPHQFTut6Y3UCIx87qWLRKfsiGNB1eKfVoUWeJOYoj
j292t3E2ajo0Kk7IEJYZQwwNcJNzuAxXWSdryvwvkhJJ9T17hmmNLMVUdkVYRfEdURrBr/Hh2L9S
Usjb2FyPvTPKPzL4wwNB0e4iqdbnbxWeGcuG1XOy0dH6PZ2PBfMg7Ojktj0BSwvtoydH/kjj3Lma
jrWMFp2iABBfspWujRzacLDME2R5h7ge74KfLX8suSUe4xVI1gF0NMKJvls2+DHRusfU2Ifw2ZD6
Ohcw1qtGeAhUKE8n7iHckpH/KBJFWM1GEEoC1ukkKHMad1jaKEqW8lBb18rBgx5jrHMfh6wVGupQ
JYmNvm27GEkMbLbEIYgttU7RsaMl+sHtRC73jArC53GeWYB+qVzAcyjwntlgRVPmYoblbpqHWSNb
h8Qh/isI67LSpsIHbPQIg550iueYfi+76VG2LcdzboM4CUaPOqoE9u/7e5YPuawF+3XKfvuqECS+
PRE5qDViH/1AdFrwhBSkcZXnj9U7lEtu7wzHXueileYh+1cfx6PEuJjDNIafR4aVLVwuBSWL5gKw
6fyzFO7fN8dgMsEp8weBFdBu4+ab2ib67Lqi0xeFUka3jnLzg4srmEN8jXdbzYRfvxe6aqEr++B0
bJjkDvrKohuvwvqbAPTQx8xMyazNbIUifFq4dG6tudI9ts3yNrOgemaTZYb04dG8mIt22PM2usOQ
8vEDA5gjJHWEOLCioUcvhnD0ekftB7uuUIXMH3Fi+TPHYy2zzSE0gtxJ4ufwtsRIJn7FKeRFoX56
VYiJR1k87qS24JPK5xwJ1UEFa6AUOSQisZwS1zww1sVWCDSqL+EOHduga/q1eCMMGyOjY78Azp5e
JegKHXb222YlUjIL0JDUluTNGGBwYZp1kk0sHbXTcAVknYVCaSgMnk9V9jRu4kr+rA0TIbG58Y1h
sp/H7/LTe6RRLizIUN/Eyvfo6ij/ARWBSHnxvMwV69F/ukhNQ10ZIPsJ+NH6Rb2M6YsIsS5Jw3MV
V9v2AdgaYNWqkwV/r6EU0ttIs5tPwo88+MyRXifzgKBOPGojzsCYrIQ4WKcKXJXCjG5HukGivPIs
RJnAtxPDGZHmJSn/0/0exz0kCusIzWLJmTc1Z0FZqRi0d+ir3igp6cksYwtLd6wOSzxb6dQxCyQk
cwDMeU/RdwoR+bQVtWjauP+80JfQvcoYbZzndUZC7yncYF78fn/evZXE7cEA6dOVXSZ+unu+RtC5
Lm5jB28H0xJtLYq/k17/ydxnpQqpfq0R2TCFbrLkbYuniKYj5S35KgakOmmung8V/QHhRbe6MOSy
37Wbs87TL+MHfsAwMp/abXTa/9OMGTD3oLEM9ImIN3ZDCRg8UXPdisOaDHaT5dMDByeWPqXY4JPE
Ov+Y7tLuZl5x2ax35GL8N/zi8onrAAdZjD7WNJUk7fnF5iuXB8fJAyzOWN2HJjA1T0TSlWiS/rLJ
qvMqM44DvvL+ejq0Hps+EqGAG1paUbagBGE3dKsm3P5wAcSNNn9cR1ZK2xd5P0IAOIokKWkiRBIS
OUmzmQG9XeEe/zuDeffUnngpKtr9PnS4/aH9DQtpha+gEfEjhPgEawyVJDRQroXpBwmLUNMURwAI
D6BQHcWIQZ89C5uUuQQ8HVGvya2C2z9rCttM0sI7Kj77kD/IHb4b6k9ZoNp/z9rj0iZRK2A9lcBR
1sSH/Lb0L15x4+Y42cHsgdTT5ky1ZK+thud9M9vh81Vy3NAJ70+XWl9K5Td8rru0xpuAz7cOumiV
OMvhmD7fKIaGmPOpjMZ3E2puOyXX/rwhftKaGmymnDQsV4Q9Emvype7nTKT7jMOO1WwKkVQpcfz6
XeCzjZCOtwQhCKuL8Nba5YE+KrZ1miRmqXIU6CVeE7AOHSj8h4zCJGKxAWQDwGcbsDJSZWiT0l+W
+1EmLVocAU4IvK7QlP3UDihNikC4+Q7VqiTKLZLrn1LG4dDbrf25Ys5ZiwzkCv0kUVaUCvgjudt1
lz1zg7mQetDML1JYHgzBiQur6c5DfCnDAIUWZcOKik3fYifcivDYH3+gpWag3fx7/8lqcrUGA4uU
nkQLJlL0VETFfYWal/atBpfgoIetAg/WsPUnJMYzcZJj3fYYc+z85EWb3uw+aONiRfV6WMGUmBx9
VVE3nGmtwWuqW10EOABBuiVg+0U/AakEsa1bAFtoyIzgtU5cSzIzYWl+2I6OvqCNdJqtFi7jO4jZ
6dqxmBrBggsx0ltDkjIw5nto2M4aLpgoFdu2rkuo8LW9uULuk5NJ0Nv0dqXnAgjpKqvnYBUXJ/5+
wkqhVVA4sFfJfmgPrW/BIOhaWO3sYVd2Z/+snPXsws21m548EaWRmTn10BjBWJyBvhW49eKtET+W
njIbGu7TUi94mL5dht1il3qTNEk7CRUCQvn2tD8jJHsnIt9CPfygAr5Y8pIHLhKC87JkLA2UKeDJ
664JXNK8vSvMbU/7jypbqHedzEmu7/dBiCJ9nGkRkApGqVg4MVpdGzEV21rFeq4XhNGQ6uN9mNHo
MVIszZtnHJDTXtAQenvuvff/n1Hnsqu7H412He6ot925MHsTuPmEpB8mlaklw9pfhiMGEQR6SN3O
Ot1Od37FQYJ36gF+zF11/gV0Q+twE94uOXCvn+7Qb0uAg/UbCgJDoNeOXCbs8DsAFzRki3JHmzQ6
3DA/bEWDtaF8yikPqWS8a/Fn+uj1aByS3KQJQe41wxEbal8pf/2uBBYvtaa85waDblPXgg16bfpN
aV2BzBRuErifKbQEb6qK9A4E7sc7Tut6I3ECxy5tYr7zM5vbfbl4+inKuFsyFiOF5g/B9+zqiWjc
PUcYsubvkCtzs0rS2DSZGogpbYeqRbdGtWlrpa/kVj4ISl5x1Tp2StZB83eUOttWdsW+InhCwl51
yG6ewyeqiaHZoWtzYpKywo41BXAUki7ETd+ZK73r5i2PCMgenJo19MMTz6nESo15ubBnoiuEENa6
9wNajI9o9x5hyUSQCkyYLji696PTFNmAzzKvERirs+BynolK+CfirapRJp1SH760pUH+jKXVMS1U
bDB59iop7roZd7rnIziZ07TfmdjscIm5fq1eu+SLtkN4zr/5Y+3IjvaILGc54y88gRvHXH/wcAGA
JKR0aO2wUgs5XJdYFym4BgDscX+mxfCqIBXqwhhHj+m27wt0D5iuTihnHMtY4/TnHoFGx2LLSeZb
5nceEnokl1AitPkFBbA9h376PK0pYtcdgMupJSJ8yJAlT+/POxSXN6Gy+S2FOlrAe4zItxZWV81d
4abOVYclOcLkl8HxT2RGcZ/RdXYSwB9/fIUImvOm29HwmH6TOgIbVLiM+htz+UNXIi7kA1UChg5y
qufzLNy8FGkfLghln8HtOqu7Owpc6hBCnRWICJ7oXdsnwBJYxFOXoyLDnmnHXCoUuKiC3sDy38jC
rDv1Qndzq2QYN6zRIts4r2GIZzyXxDw703Wut3ISdTObRH1lbIGoSnzA7MZn+PunZihM8omYhz5o
IlBG844YITBgK98t7fUx/2K5+grLUFvxgUbPrZg03jbZ0xoCldufDhC29bh+TkeuWoVZfFHDKrlB
CfNpmHRnulcyxh2af0OE1My6K8RBGHllKhWe5NLE3fIm/ISKFwp9ApB6lxdlmp1XqTmVUSVB6bys
5xyX4+c32EjCI3vs665HhH+yIYyiz7+QuiNh/DxOm5YDwsZEH2E4irpAyi2cUE9j1jn88cmU8SQS
rm0Wc8WZcZc3zVxDThGLZHcoNROSM7mYA+n3SheUXfFGE5hRi8iKefGKOP/8ka0iKs3erCHPgZhh
qiTUO3tZE4krIawNnVcn7EYZBTk5zl9ky3zOTMl/fITs8JqcNtZkQrUltf/6uZp0fx+AuE0z6/iq
umc52QclJelRUcXeEOFLoSJx5Iro/pPfWinViXEkC4KEAiebLTHdFf1D8HjEc18f4buNNvZ75icY
x1pATqZFC2n9r74Xt66Zh434cPOnfQ6GvNgKW9j24FVAwp3IQ49EmahshtvkquB20G6mHHsYHtvD
LafE2Sb8gGO3AZwEMXuLCZYesIj1K47/zs1vGL37V/RrsrGhOGKg1PNWH7sywLqiwqA+5SyZGC8j
ryRlSUOe6B8at/NJkDChXiFJKivE+eHwj+qoeUx9jJCbZ+OiNiUD97aaeu/NDRciWBYskndH28JM
QMkLyruOO5kWQC6zxlr3x5RjF8jrb/+fuSKBeIDnQEKpTCdffQW85GFtyG+1JO7a7OejW+AeoofT
hybTksNkETClL7+en6b52NGRJdFxUxwCox8Yi0lzkSNQ7I3i2uuj0PiNmLad1D117K88Vk4BMq1N
iJk2npMMGqPYcCfle8LBoNz7sasmt7esGwZqrROZgvpvz0TC+/0g2HfbagmMfVFbLej5Sw8bW4u1
YICdAztjF3MobuGXIWg+SHw17zQP4KqxZDDvVsvuF1cML/TdsqIzJ9bCEmHrtNTmuQCdmyobTGWD
wwVkZw5CeNq6n2At46ej3r77CNoClIOSul4eIXts4Rvngz7DzeYZxPy9wANaS/WJ9fzXv3B7uUvR
2qvOcn6QIt3Zt+73z8z4LgxlSqeR7kDvYVehGQnBB8jFaL0QSKB8NpOdwLswv+LqLao6S4PTHQmm
FklsSmRVz7dK5ziMlIlQAhlo5YfH9jbwASq3yTIbEXsWx/Y3xORDEUQb17wFSVFw3FR7fIK+ebwb
FFdx+VddVe8O2nnx0R4zyyqZvlcUxEysbvYfUnLFCyzRHmeFwPdoaSCNeGVP+t8c9mruBWoUmgPP
Ya6W6Vh1qq1AM5bEOjRCHvJcVepPhPmJ85br8uv7xc9gE9gbUP3Rkqp2jjYa9vflM0xfAh/QKjLW
LBA9RapVaOuFpOlWQZ9wHW6+f1gyG2Lxc0N8MSSmdpLWr8W4fUmTi9/DkGH5JS3zvH5Xro3BFCB6
O3a1wOYs6rkNizHfF4TaIk/jW/CJnbfQKCgrn5yQk2yq5MyA/accwRUPJn0D/u/DxAllM8B7/1Oy
rkTWc49+Zg3OUXLIsXIPxKaBuSai0ZcNkJetqr7ZJLcznhN1YXL13yHOTaRpHxb1FFWm5e2KyCZu
2i5/jS8mUMzuVS7UeaXkR/CNNXn4OW4ftJqe68TBHLSttPGm4ZrwHB6SdE1Lwj4HoCJxXYhjD+OB
ZEo5b/8Iz59dX7LGJhvyARciovzYzHCLtHrLx+/Gsjsl5sNPQxizTJ0VayCLF6hBDs32oWVlZ7S+
HkIuXb56Mf3RRoqLbjCeszn9znRwWgLLLAUbEra4ROK1qfCp9e3nazvgKKC3/I8u8TNQhwH57B9h
ZX6uH8bzSiy2krfwSLjUMMVISGiynHMsuMcawsG/B7daQ3BfiuRFwXhgogSOsgOu+woPi/sH3v2Y
rJKfLX8wN4+HaA8Cv8SkaAknJhykqYD4vopKMB4+LYqZ6sJS5GiluuFJf2z+AJYpHwN+4zV8JM3Q
HZ7IiUkdMLTG9+GSLBN34DMaxuP5+Jh1Jg3VTohiRzbO0cJjm+lqkSP+2pf5p74EV9nnx9SpFcR6
/+QBP9LSsfNgyBaSOuaPWHfmv0+BXD3RmTyxs6EZVCfSoc/j8BOEOmJaApVSedi8afwPycmc5U2z
Md8mSit1yNfFM8t/gA/WGU14In+HNnRw0EB8ZkfH4knOICQGnRzU+dxEJ3MF8XIdxvTy0ATwQqi0
nDN1sJdp/kztWvNSlvA1e4+91RaNl6F+3XSTyh/QUVb8z/LsbeaCmf/swipmuKZrvyA5ErGThDis
r2ywwXvEL+TqaeoysaDO6GtoktlSoOwuRI7pmm27JudxehgeKMIryfcQZc6Ds9S1i+KX7/LjEtSR
A9Ji/Ezkk2bvH1a9xKnBmd7TWG+rLVG/M8g4MQ7QvuBBYiLnshoG24DAYIDixQ2V5miZPzV2fXJp
9FeyG+dKvB+G9pyJw+n8HTWeqsAhORaAybt/aV2k5SPL9HO4mnr60mheiz4O9e2VnBQWYfqN8P1J
z/Bl4IO1SUBML2qW6pYAd/A3wjzvTtbjeWnaQEwbYugnz9a4j4Cbdd5W3bMPC7VUG5wWfZvP216z
7KIzJhAxQm57UbWYeyoiNtn2cHMMk+yBUoVx4MHrfeU23khX79Sx+DLfhMgK2cMebHoIFDhuV3To
em5pGxXupYBsWtpSLuM8FHaixcI2i//t7isH+Q75HakJ+JMUS8TrXEkUYbvAfIX8qfmjUMrt4XWJ
6MO/1cER8qJKhvB0q5H6/BwHQjjkvXT/uXSiJ6gd3A8knHpGglrCokO3Rj6woS06dV7ial4ZNr2m
3Ur9dPmJuLlPnRU9DkgDDA4YEtMQZbC/0klais2b2RvTI7gb0U7Mt13kU9O7Ly5xiGWYA56TfnSz
AXDHzFFDPhfBU6HLSONAeeq9Net1kvfT7WzE1J47edTkpwuNjKbPkkm/7mBvVAg2VfUSryqsQoqn
PJf0fR6O4blEGggpnkqMKcM74tuJTeMNgXmmrEyKnfiglVYz4Idp/XsQpKgyR3vlNHmucMI0P16l
+Q85xiilwlyDe7nJ5aNUObVaelHgYwKxE+ZkVmEA4OK3VjsMe/6BDgJoaqarAO4cIKSyjTVDbeY8
pFI/LfKi2APdo0NPyQByVIQimjG9nVy7S3zgO02O4+h7wuLDqkDR+u/cCjg5Q/IoSVgrNaKCxNtZ
xz1brLj5AZ5Un290Ue1IYFmk88EWbsmT6EacC1ompQi34rYxCfVn0nox6/HxUF2PPnePe/j9Tv8c
E1sOMnnhYFlpz/zDSVsbB/DHyWoSYzrZHcA7iLCGx8mGynMGGEmIFNOD85R0ZqVZ4k8oaf6bDh2P
eEBDwdmzltVMWMsL1YFUeNzE4qoVskM2/KpYlBtH9R+kDIYlz2HpXmPcZKIIDIkfKdpGe6qrSh6Z
jagsLxZD/qg9tD41++v360i8YWJ3EQp9UBXa+CuoAqBqFlhfvO6n/M203I2SCnZa2dehhUEHR64N
cs8oopXzuaYjwNyqwt1xA2A0KjiZ0noUYp+RPvtW4cFZNwcsksfp25UFjjEmGC6dvNceuMkdvvcj
IO5SPboAFqVEIb5YfETc2stom4RrxtcUne2qYjU8kfrmmsOI4GIIwYa//m/Xse6u0q/NhDghbjKn
EqkeftzOveB0f7cGetYsw8dNMURl9r+Dk4xT73eyLyDh8USKWm4j5JrUIeh976DU9iFUURBy9ohD
u4dA/GaXueMZFqQqdMXLhL8eDQxd1Ic3DewFCNZ2kX2ReWtLW/G1i2L+mk4OFzpRTEZ8w6ZaXKcU
/zjqbqBd4vpKa3P/wA8C9OWoxGF1oWDlL4Pb6xl8plQwlNfV9M4HewZWyqdX8aEF7SvYUsqbAUg4
ozQ6AxLiN9Ra+SYXV+nrhBJedm3SLWupKbwa6ECXpIKd+Q8IqNyUX81jPXEssROM0diJk7h5/Evp
jlAKVncF2F5MHKBvHt4X+sNQWfnDYeRqk/KwkJS+CdN/RhSLuZ5BbB4LBlo6z9H6246TwUNdHoqK
2dNUqDi+oWioRJTF8zmBFHonlScUrIJWLF+g89x+7vDFpTwmjo4uie3RPcj0jWAe0ZG83wjuF0un
1N7NSgcDGVOHWc6fa+ljHI6O3OO+rBNgHosCG4hrPAGiThhfFmr9M8ySLSdSsVLrVydAvSnbjhjQ
wFgL99xuh282ObD/4DO60UIe3A/oI9anF73Jxze27qyzwAK4jmy0RYdAMTlwpaMWly2CevG/sTpb
oDLk6cxf2ASCXWYj5BOHBIsfdDnQPLonkxQs2GrGpZZMbaXDwuUVWRtNMrX/WIawfcDRniWvC1fj
l2OumqREiJ5eGwQWHkHDc+XD0v2sFi3Tmirg0YtbXjInOLROzM6P7H16gSbACU3oZ0bqcbnpyaF6
HPJe490NtNNrV7qE9s3qAmod4Yb06MdmMdyZhp4Vya9DHDTCU3W8UeA+Iga55B5igNo1lS2ahU7t
e2N+SzNEIzJgOzYfY8fa87w3nEdb72nXFeiYNnDfNCeNqfNLCKr78WXasR2qJTUV238EEBWwbWGz
x6llEH/dyBCgKZeCLyf/3SXNzfC9ReFXtpegV6Vy7Hh/FkqJDkaGd7oT2znO6/ob+eT8QWX0Wd9D
sO6+ZbLts9+pwN6ZMF1zx2gxeONiariEWsKBpPgLTtb652vZdEpkSsZO6E6zcyZNTbKEqPIFek5F
F7xy97I+9KIsdTUInFtRY0mCrSFvgwEdJ5XVaPhgUFSkdVChNWS2VDj8SGcDO/6LusFAXRUA6DGV
UKJF3r9H92k9tFEM92fmVvAQ54TwpIT4iu9h/NoonlmEpEsgQUTomsHyTE4wm6INzEbc87Y8gLLD
IqZ+sjpaj6bi2s5tvtAo+9Rycnn0OKm3rpFeylQh/aEZD903DBFrZ7zmU85nMmYrEiPXl4eSwagT
GzIZDcx8EEvIz8VUKqpIwWJ2VwEOoCI7OQRcorSGvkBw7jsgbSKbxNiXO4D/i6jMI5ReUN5VIuC0
RJwy4RKOfvY4XW+2A0S5Teo26kgwePTrH3H8f0ZDobvn1+kVXu/JaKp+LG36Yh/zso2rLdQjSiNy
21GuKnsSTWwEGKeYAuLoa1BemgiUufRqO7uKkNlLIWZPnWDYPQc9Ej5omVJ5lopPwYiB1AH6ituc
0Y+Z9X9CtfWmp0IGKBNoms/RqKYKkHOFOuUri8vDLeSD6dAgRhnB5V/onj80U/eThr60CJR4bTaX
sg4fNwNKs93u+nRFTHte1bze9dwoXhFWQnnb2kba9VmU5ibdCNv4ZEcwKZco5/1L+aima402V5u2
EWW++CKBUASAYZAIBCGQqCPpqXL7YhAfFvBy3bRKEB/RjJsvn/6GRvCc0e9SQGzyfbJkZhcuDdsu
15pI1haVMdtCaxhsJkOW2PBX53rG/GcJrqNerxSm00lu35Sd/hylVnYNAC6ZLo2cA7mejNWBuZZ8
EcYHEnqBN4qxV9P6K9Japmo5l7fdFMAQs7fEvEJaLIcrVDM6ZkP7LTnSVWfmEUH2iTX4v9zQ6MT+
kl0OIF/wjDw2Lxt9XzMU4pv/uBrI4Bw24vr3ad2SlnIi6JBWfQpa08JxEFxoTX7E63OHGy1MTJMY
S6RXPpoYbO0AnkKxjma6nQzZHjB/V9USBniKH6HowywBAtuoVwnF9M5stBJzaV2hNVJ434ub2YyF
bVJdgoCoqap/ADKss/cb/NinKm0h0iqDm7tz0dHymn1M8Fir/uhyyOg0eLdrYk9ohOfM6oVHokTb
H6sh4TvbnI4Sfp2U6O1blZjcT7ciMexZip/tdxJ52XKXW4XE+uX/YdtrpFNBf6N2zF5Htd+nXvKT
/G48EAPWF27WKmMic/5tzqNcJIphBhwZzHMZN+Qa1s6o4I+bEQLgzjejfeEadJaoSE9aZh2mrIYW
y3wWt6Rex5oLfa3F05PcVCqajquLPxxrk16jI8hd0+jOVRIQqeU+BkUMe0DiUoC9XeQx8/2sOfhz
g/cxahaU3sJ64364FdXUUHgooDf6iP/FhFW5srT2xuka5ycj0engQJHYgpKW/dZz6KAaWXXE+A7q
fwN4ugUxkS/te8LH/UswIX+/QuXaYt6FlMNVGOWkSrQmu45IR1hkZAkhhZ6yDvSPuvVV8HPJ8vHW
CP+Z0fbs/7+kwGya8i9IUC/iwdT7d79N40Y4RXpMWtqATjXxcdwyPoM79n8hnGLBvkvZZZO648OB
BeQBfcFdsZsmC6qYHGyGJ6HN/KZnmo45HiOuMWiyZ2+M3uPJPMtHfi5+/aIiEPVOxV+ZusPvHtDJ
ooZMTv3gMpXDdIKk+8wojxsy9M8mW9ZcmJ3OH2t2rgxngyV0beVzd7SLA1PSrYW3ZXxJxWijlkiR
U5L+qO72VWfNXrNe1LADGxm4Df1mBNOKwJr02qit5cZNq3M27y2dDPq03wsgcg6Gwcc37dGUpZii
K1qXPY9kqFelFVDbnGJEiNwA/iRItDhlszvq9mIjON7CvC9DlXx/2XH8ZBob8ok4UA6XrLmOGSkt
6iTlAV0cPelsRosIIeKFWfMsisBto7pN9IqHBG/RSDgqVghXN2SLrXcAgaA6Pnuq7wnVkRL+RWLS
rWW0ek6Htdxcg+esir6GXuIehbgLkrsU4j3b8JwP+74BoY/6x1Do7UvckYEdAUae0dRGt4n5mYuB
vRTZ9ICWoewoEiu7ET3N2NZb38sP5VfDkzd2FOL49NI4BzZtMB8qAM+oaNj/xwzTwD3kBv2MBUDu
g6tqIdTGT3D6pD3sw4QBpmfjiPl+/D46CQFpbtdvMr2B0MmuhNsvyySRRYXgYhD9mPMfKKg/wRv5
PKXZoFecOBvJLWVIy8cu0PVRYsegNVVaeTuWI6K6gfqL3O+d8q9WESmMsuKo1lJWJzSwCfnkIMF5
JhjOOvBCagSpHQ40cjyk94Jkp6kA5TLRdg9QWPyg99ZAdH2fn1N0iA8OLDp/CH12qn4rbLBylc+L
SXUjPCJ/0Xq1FYqgbUHIEXCk9iEKcYde3CkK1pWsgdSHsYeOGqbvH7QTPEGtfJAjrq7xxv0tNDHt
bq9JQNHdo2jUhtXydRPDrSnQ6EuID7LwGXblkzfhJ+5zlzRU4xvoRcxV4JCZXuf+A5zuYg8V6quN
mXI73R6bbmuitKXDdmgfQDVAsVb/TQCUIc6WIPOZYG5ubJtlS+DtR9uRT3sNhOmCakUIFBoIVuxt
NyFcMu0XBkckM+1Bl+UucI0ZhmtuR5yGVON9kXFH33ygwXefLlG/olLbw3ggsWg+OR64UoY9c+S7
uFX567Gi8VQ27bxMcIzUgnK/GSznZeWFfIU3PcMsrgkW8NwSo+caqeeFj+Y/nGmagIvG+PU4iMPQ
TJTJan/pa+VNr64JmVFYfnIw4bWmFbWOFP7ylQqLsx9lL9Xuhm5mz6fnoHP6A8AX5A+Xl063xdS8
6cO59+oKaEJJemrrQ1c9f6z69hGtA9wgoHTzetmNAK2WQO4tVV4xqlh+48cet/o/IYRJc1LkIeCv
uzXclv3S4JD+0kJx8Q6LpVm1le15CbvsbxJ3KrjCxAs6u2ggkI5QTW9EpaSobX8aoWLazJb0IMZr
C7d8Wj55z0GhkSVbipK2FhINcJL1lx0DE02vD6pnma/8fXppAsgZAG4BNznsN9cdFMNJe8cVSmL3
OQx3Z+6bqvScy9N96X4uIDOB4OpGBEJbzkAUxWf7PM5qxHWaJgtPhAmfRxrTdg6UahnNtdkGns6F
EIxMbKJV8eG1FI9FrVYLQ1OkHVPZ+kI95d8LhPXONT0Un8rKf8eIZjB/6EaN1/GlOn4lTlGZOwjf
stVg10B1vBf/w5DnynPzKkjC8yY63KtlqG2rokwBEBhepOQ87/uN91r5O5v+KEXXUNcPLPgtFGH2
txbi0fd2mb/9anVYsECHNYoTNqSB6ow9B6A4xQCipfyrd6LL/ePNuk2/InUtSkz/Gza8+guNQGCV
TAnjQQNG2FRmIBCGXdThNNigx7PtPHIzKS/kE4nbKz/wJ0JuJ0HJamuqe/QEbWI4wagOxQD7YlX/
wNC7b570M22bjhuyUCD2kwqDWkwOe5Q/HaTyKO+P6Ldn8CKCewwHjAVrIqO5QPAVB4+lp9BbNPLK
/3pM4sCTNkA2+Asl+0xfkQDOFhOOKjYzNGvzoWYujeiq78SFsDfI7/+xvo7fUtHMi6C1cPVbAtVA
a725dyuYDt2sAfRvDq/Yo4ZpVxcNMOoyh+xBEdQKdZRTBQwGpK9P/9qqHvUED7SVBsZ6kfLW1WnB
JK4KV6IEOfBnMIwK/S9+ZbLQjkzm7iUSHkKzHIqtq9DJNA3h0PZNsN836VA6Mlha3IgK7VuIKWkT
S3clQkLgTo/ZubLfnStPCWgXj6QkC7wXTU6uM6ftLAU1iPaLn7oUrap4xKC+bYGxcaRJqRcEZSDg
kvqSPq5bIo9QdDBRZvRnL1RkaA2oCd6DeCY13sVqvlkTyH0z9IexU4UN33AvhJ364QqXImsQjnrN
G9Ih9mBif0K/HyyIwEbLN+EoFsnGRYAqUnChxTYC0Q4/bLegKyCs3h1tQm9CcxGq+RjppRBpkPe4
n3vVB1WmcdCsBYCMFHy1LbZKpYOxSLHUZXjPEAff8FXAFdtf8lO0zHcLB9yLd7lJZIrDV72ca26a
7W8HXRexoxYyr39+wJSxExzfiwVx8PXy0sJBv1hGHaAB2/rPJobynSghDGusk46gbTXFUN/OXo4d
+vpMA90GjVsk3u+D+Qg6cEyVk7ny9V3/X9IVMjBdZ2Q6UMWcn92WgPTBFWxQWZB2Epu73VmL54jb
TykcmsnsXhWysAYVoCjDROIggAa7K2fG7B3ntdQUJOWv843+CzIu6kqS/HiLYlFOjpX9vsHe2mgw
Y8v80/ceKquLwgDS+Mcw978bMEMsvkQW3V/SSq+ZHCND1YnkF4RUUbeEbnlrqzMEPd3yBr6BANEa
DpIRu3WG+GorkRfnvc2ltqcXZXlagBQ0E5ACe3Bj2aO0aweOkCDS4h4iv1Pw6vb9WBLL3sfU9JyN
jix3yNuTLtQ6kxhN+ZYYhC4cl9QN1wvljDsWSfUExU7rQfHZ4+A8zvKZ6WZkTXx2aDrehZ4qztJf
L04oQBr0LoKYX+e6B1jnYiAGJiXLtkAzgYbPsjT9aTsEENEQNzKvrLLQ+/GpK3PX7OViPkawls/K
z20hKtH1k1m3ZB8xoZ8nQ96niXmX7Tme8fADxTuYUSqUDr8QuKnb4bJkk8OEkYOQRqQISeNAlnR6
FVSZ2XI3G1MZOVF2h3m/+HTN+5bjeCD5PBi6qOL5VSSYWFyWblDwKLnLY0qXbCEN5u+1b1uRlIk6
IVZyUF6eWf9ljXy3P5U25Kt/oCVOMweGnZEoEY+3HGQAQPyPBSDUOybHOhobPtHhBqA1YvNkb5us
j9nvtt0IPfN3DBn/MP5YGyxHCutTsfrNK2DVC4oGDDZ4a8Wo4J0QbJ7or6NMf26URQuU771V0TAf
I385GXYFujK7mYVYafuP84geIOUgzHTaxVV441V45+PKG3eCViy6BVrq6Sxu5Mvyda7zmN+0K+n+
Yy0YNyLJTympu2AyNV7AH0x+UfoFekBwvASMCspWOK4yRIp3WJRrY9jMuwigb9tlwPW6ZdYhfBNq
KP62HZS9OzwhJgbEsYo+eNzgkcuwgk4bSmbq070GV4CWDe1Eo2lmDUJ0VOEgre966EElD64G5wjT
nESE0ImTEPKekh3aJyWmdOA7MeDVqliUAWfqUQclOktudTA5B/NyjLmuhVvNQf6046SrqVAEO5RZ
Foho801CEtetzyqBx1kdAdjHEuQM+UluegRiblzZkAHwlvmxUrvRYA0s30O0kk8yKH0t7q17sqjj
K3DtTQlIDOXk8ir1wEdOMMC7UDKWg7m6hyDX+EvB059rHohuUg0sE45yOk/sjoEs2X/SwnwQ1ysD
JhE6T1iGAJZblLz+5TSTaJB1TppugJ+uegqaL6Z+WMc18zOxHnmUTEGhOTu6jRfHYmh41fFqWUs+
eS6VCR6nTe8MjpkZF+1L9wjkIzyd+T1xhKwhkyY6qzBGLHU1pDZEOTJDh1P3n9YNDb8t5cTg1mly
w80SDkE99AFoM47HzuU3/hg5BjcwiFqoezrm4Nb9qoipL/Rs8nMBWlyiS71lhmSbsUfCsxp4VwI0
Jwyb/3uh11sqpPd4JEVWl/caxq7UfKGRSASAToiccajWsc3AYbnGzfd5dTZupcvwXZutT4xBu7kP
0/es4IYi45OxmX90/pzag6KMZof2FXc1gkWusenOjDiUluhOkI6ThMYwRFsE9JspoGZG/M2TQWbI
FtdTBLXRouV8eCFF+bqvxQzsfMwGb6hKY3TGcfyvx6fuSJEg1ru2bsOTXjKUc2vXfnKrYd+lS4qU
YO31pE7RYeA0cxsysuvW2ro+BdnKih2OT38ySXteU91mDZTHf96GT7l2HwwxfmGweBMCG7NgA+wL
oACMNLTUGcwNglwqGSnSjR6Lhxt+w+9+81Nk8lTT7SR3od33ogFollOjz3mqTOUKtUw+c0DqBMmA
x6Tmj4oL8X1sun+tAUiHpHNSP8PPT0sQ3N1c5QEfmFuVQcauLHiO1iT/BIRe/L2mly/JZGq1kDml
ShFa4IxI2GdCg6hUFQULcIPXLvpc2eiebnbCsEU+uinACkmyOY5/rikrDTKWyV+qetXDBLIMwOjr
/EJOJCr0WXp0usrBoTsfo9HWVRaxb27E9x/8PrzUV1gJXs13j/w9Klgt/vgbFsxWEt0g7GQ4UoBd
HpXR122y9DqZ0rvyxt34oyxx9Fss8cYaLB6uHdPst+ze3Z50mM95W23jstci3NWYnEuMQw/bbA6V
edAerrRZ1Pps6/wYZb62ShqYeJg6R07dc7VvHFvNdq3XQahlH9GWGIuu2ThbvnBIAu5q+b8wQ3TB
0U/Io0xXvXep87JsjMnOTS6fanBowq+Q2BlZg/ZEe/axx95+lJiHhxHgszq0qurg4mfJhPQ4ubw7
oXCBONMD8sodxSbS9+4+q9KB+dSy4eYZANtFX0kGoKe1ZzcZRof2RKtLnrSE9JsMPNkIoxTxtEzc
NUy4uhrf1SzrdcEzIUNvGhx6RdnsS2Mr+3Brstf10g1g3werz3a6BWCi5NrE+yQ3wYzKs5TLul/6
w/a3qV2z/+TJTIVEoZNnP1PPvbiypZX5A+nODoCaSwg0VvNfJWvviXjIxlOpsAmgSbFsqvxQutQO
hbUgBBfNPeakx3ZTSgrz6LVSzoeRQahcGnfZg2oySG3h3GPpHTLwksqV+YOi5q0EURQvleEXbnJI
sGgkvMZtqW0MFADC3jH6++2hH0c5kY5FZ4ZI+XfUsvJtUtyXHOOpu00qzk/Fbo5IadMhf6fa1RFf
kpVOFc308wcUkT3qVJPJMSYb4okMnc1lToudQ0+3tZnVGESI+0s6J6hKWNxFB47Z/3rDHBnYgxcB
NEOgQs5Rlha0eDaK9qX7Be2diLaxoSRK5yR+Fi4PTn6+Xhf5Ty+a6Hx4486RF6jPM21IB0Rvt12y
/DGV6E/3CmpaLzOYiW3wR3wDOPZO5DnCfYXsrxS0D6+NZx3xLoKnZD+16ZsRnOl3sQ6eAtfvXHVc
ZjcV18ewgQ8e9E6GosgMfZa8deh74AHRlouTw3tr1XllGJneaCz6ENAwnGz5MU4aydvs1lilPhW/
tNJTKa7Dvepf4JYpTlIodHeWgP7Ojy7lzO0TMec8LJf8c61A4Wnw3oad3pd1eK5ddaCUfCIP3JGY
6lprbhuVzO9cYePyG7y3c+ezjtmgWTCOORUcnbnqqj0y01woc/00TqkJUP5IXABZRHu75fa1xZzS
P6UMB1ULyFxDSl8Cl/Zzxu5BCiaAJucAAGOSDKMPpX+tk47DwqGt9mBzTSTsch12hsmIB1t/TNJG
7WWrVuXzLvT2a2Da/Ap6Fhp68eYH7E+j0pPHaRqivLZeMArEfM41cWyyeavd9sL6vh7cxYOlrQVA
5UlkJUN9gxL96n3iUEzjzIl2+0moqEplbvVBaDBECOJ9Tt4KAaqLDVJNZ3n5dovV3AJFnYePqUg9
9UgEQtiiN0Cojrmnt9ZuntirO8bDiw/faBUVTO8hIVaKSyU1K2UE2dKmuljY4rlNDvT6Pp25MqZB
vtdUdstsGa6m/lFxLk7l8Gqe4tQuM5xqAdriciq0pYbTnHnxwvF+I7OEN0TfMQGvGLps1wSWhm0Z
+F9M3s8JZEwMNsPs3u5W5e2Tuf2pYiazb2aCG7WCRyKfxbimUX3UTmN/LPANPld1H+tc80A62DLr
U30ESVDlRBikUAOFkc4jjeYcwtx3mpqFxdCyFadCyU3TgisSNmTWVA9xOAcFdvMDhCrzHCUB7G5b
HPf2Nwhl2BzA7M3/3eR9liplfXKuGM00O3BEcRsnygErEWUsmQeLeF0wqEsp+oEKAjWGUdGgAotx
FTcKapY36bOi6SArVRMYlil+AfeWMMrLPB0C4DfoNY20cu3NJYVlO+JpeySt3V0XoYbR/NKvaZdg
yc9kzGXg8fdVfN6lUFAs0ghVC5+olHimbKeedHNa8wZMmzIOG3fJ2aq1K0HPIWgS9iuDe6zaIUdK
RgN/zUmZCsYWVNb720/9IW9hV8KRwJevi8n1jZznV3v6Cf/xoKKWrKMCuEWcU+JzaUMiUHqu3C/9
6gZlW34FidEO2M2Qa7V6ZFaARsSWllyDlEOAooJjcuIq4NSozatcI4p4I1+tUg+0MostfyOzM0G9
+pfcbbHWwLMmXGyPbnup9jX+7fUBGKyHNa0OcvugneOtzJsfsJQBSai3ZyD8lab6gqjvM8atHcCD
D7mQDfFAmS6RaUcn60z2Bqz66PlXhDjNorXxF/OUIJm6uJrT+cohuXBEhDley9qVQn+iYq8qX7GO
CslOMJE6IZ7Eeqvt8JhRwRWRhFvYcRITiNYPgMol4b0g2m0EmsH4Ov3cG8X2FxLcTAiUUfSJ2m4n
fvnU2GKnI5kJ26EhEiNrj3mk5RGzO8x2PscLASpU8NPq/7LV61uMRxdg3sknpLFmCsENG/CRL6mf
3i9HRMxwfETvDAZ2LLqaYaKXd45x8oDoruhrdIRQE2e3ygIfxNSWc6rz0TM1oD/iUAfytC4zwdSG
Fn8/UQ8Mx6GuoSHx81CemFGWRxX2KgkCTjdAc7BIclOhd1AMZ5WRrC4k4RF/DvL1Rzz0Z9OL64hA
zni5XIW7fvlu8JV+vitsH/6J8bg36D/p0JE88VBwVi3uZxmiakUQg5Sk7ElYYbRgw50FqdvZ6a2/
+2jiOErPFB3RT/KZZxgPAHv4oUwhIJFmACE3H8PXKMyRmXq09IFf4a/Snf6sTzuG+fSQ/6lrGlS+
zx/GU6vwXDkYaBF96aVaNfFoHjfuS2+u6+1WzHsvrscgGQm+uwMNzza1MinVDEIfbNfrlxs9mckf
u+Ra7W/X7K0210vcrO9nN1I3ExODJ4ktdKbN1uXLqwcmGRfENh+Gnxuw9y4WpXTTO7nyvvLt5wU2
27Xoh1EZMrtRGtCqy0STftigmnldUjdNWv55rV5SOhn87JY6q+0xr9tIQpjmxuGpRJ/xzdhtCqQD
SNZpzhAI/zQ5CZYjyfBFz+TDNKMUuDM3Ej1SCbkJoNfiE+3lehoESrpvSOAQdHVK/8IsuNOrHaoM
hrCEynobnqk3aC7+4F4UsfBgX06gZgARQ4GMahfOGAPDDcDRvx6OnueJw4E+6ZwSEA7XHCSSFBJn
dbKKeMJ8ZTsT6yRI2EE+FvAIVHZg7wAz4CYahd+eyFNnz6xwQIxPHNx/BuhPqqJzdM20OcFv5PUD
rxguZHXK9W5rV8iNW/qVGH0tfAYzM9Bs94ANtX+GYaTTuQpb8XZ1/oEgrqVs+qE9Hx6f5e9bbKQw
QeYuhl8ykalyigK+ReMta+OPMRCSyu+snOWtwOw4ydBoRcSdJhWiMixNnbtdL3PcN4xcknA4bQYf
9Kk2usMkWjH8SMp02xQTEQEHYCMtZfDnizCK12me2HLQPjm9LeLX+XzmuQE4JOjLdUmMVWrB1QZi
WFSkd6FgrsnHaGnazhENCZruACFQu3O8iYew3fu4NEe3EkZrn8rVt4+N3iOAf8YCF4NQjYI+dmg6
rmWQd7HtSFlXuhoNu5Gj6mZLPyEYbtQyD+y+GdC4skEreaL91Vg/qbgNbPRY3iGyRDN6bh6I1UNJ
6iBWPiTEZzMfnZrbhRSMooLVAiseSYTo+Tvi0Enw1ir8pOGCv5600CLBdO5DMMCLQtVHV4VNAtQZ
ixgLuqj4STiZdtCwnV7QAiJ253IicvAJqrG6FyQEZjfxFxPpsMm9rdnl3EzolENhqDDNt5TS3Jm4
lRDpbjnXmsukY5uKL6ebtqu+RZt2JSFGL5PAGHvQKKgq6s2ax3KjRb43fWIQQbFH/0wV/uvmiutH
o7tMchJziBDdpKf0ppQqxHPSsPo30vQYPJPwJte4GuHnn2cF7X6ebA8WKxvULtg4UjxJ4dEEZfDX
TVNa0hQWANU3WQnFLe648X+PR4a+a6kaE05ova8+Y0bIe7nixPaymJ01iuv0OmwJ2eLIBREg+L4W
4mGKHx1f9gfjTf852e0093nTh/fv1pZwdHDDWUjHFZG/XrYNPSortKzbAHiIO4Jz2RglXCf4iCpJ
4DRJm4H1N37azJVXcZ38JI3Tquryvm78qQSwWbHG1aSMm9+cGjl0xeugUZhVnIsfs9qPlr3Fw6qK
7PQo+21WHy6WLobv0ax/o7Ogxb7M6639HVlgOe1kg9lOt+TXCiHqlucpdRu9ylDRaUFzTYj66Ge2
OrBttx6FvEcHFD62mDaYXjJNeO/GLdWW4puC9ueHvXmD0Ko+xHtmJQ5AIfkAMF3gmLf1inSoXRLq
n+P3vcOUu8Yo/DpRIV8q4LRIGF0ugg2TjRMhjVQAVDmX4KK3CdhzudT5oRkkph13HjchK0c/sjmY
9/iMCoArr0UW2k0doIlC2c/a/KYG22Z4BHGhUUwhPQ3mDbGSvQGiE0LML6rjxkHhaX6jcRwcql8j
HL+HDB5s9SO6lpoGNWJBcRCl98QLOgyNfH9Mjgo+Bb+ho2tERd1E/tzFUOIYjHNWhHXnp+tbsNj7
419xbPo3l6O3N3Bp12a/+6bKI8xrpjdKrfI85OjmVZGNtLIlJo83buJu/d7vlqK7tgTx1tu49ii6
bNriPEQezsD6GW8JbWFPPLbvxpfZ7wskZeVM1IzRCMPIivrWoNO9O38rqYXb4ujZ2Hvr4vLEgtz0
j+9lKPKv3bf9RWWvgSwjlyEEu5EIpTO/xk/g4EzT6/4+1bagzsCjGDfI6C8GRUTE9zWU2I5f5rH0
PdRdEfywFt6UMs+lHtDb0g2mQVnieQMj6TuqlnWB60KNacL/AtUiV73jMm9XR0VyX53ubBf61CTO
cw3FoLOLtw1Hk76DXY00NlgBzOCdS0Wt3i2zwwMjF2bIEpzHtjtxjxVJ/fnXuq2aRKrnRxOCUJCY
NlqF6ZSIU9R/KTQ6/6em9Tmu+qZK0sXUTbrac5ntv86RTgkQlXGcFk4VyWGzFPJrrMyWhn84shou
KBpIIfrdL1uT1HvRk/F40AevO2WvbtcxIFE1R0kbVV/uS/TQ0GpskAe2gMShzKIT+TaSGlmXhH16
yKvY9pL7aV/I8wHxbWnJ/LLcxFMT68VmVJ4ZmBHiuCC5JATVLf5BkfrzPPF4UrFwoRDMLp1mbNpu
FLE8bHY/YM5rCOoSYmyIXMVJf9WmlSgyGZZjdgCZpH5p9USeDsxEdYhoOOZl922Tajr+IF2m88Rf
dEkFOC42Sl4At8IK7Tp11/beXtdV8YlDAUh7P80nTCL3O+lqkioCh+yFp3QDb4OAo85WZauD7YnX
G1fhiWWdCFpf8nWaijBoySbuNiv+W9peunnX/G60hcJem/KZkyQXuJ6KDpmATi7BIKvkN1bOE4R8
AUzaZ7VhbcmZ05AlPKgqZspp6KhNfDsJOZnpnyqXAAAADPSgni4Q5CCD118cfGWm7I27zJ40pfeg
qOyUF/SMqAqu/tQmMvLB1Xp+Svf2EOhxg34I0N5lr+YhbkEoLORZ+zT+rCAYgCX2bv4O9qLeOZ73
Aj37+8Qhov3Nk/QXObRxwO/QaIuuTX8CAx85zga8JfhVDGTAriNSZWJ7exV9DFsAqc3i8q4X9MAX
odBMUI7dK8/Z6MYMhH1Gr7s5ynLRvvZMeKgSBFotIKlWcCYN6xPsm10miP2bG79aNr+QKwV8f7q5
eJoB+hNxT2BDzPBvMjTUmiH8dZiflfKVDaERpw39/hpIPFKZWSguRuSximlSRrpq2iO+E2RVVYIq
DIj94UC8c/wvtcQ8TGedvB0TQF1w8Ern+VgU+nLTWPKbZuAAmnz7HYF8GPSuIIt3tzQ+EtR1P0p3
JmJTlSFX+Jbo48x36sd+sWlQyDwHa5PVz+NTY7TXshwXc2iuVytIFjFRXaFTDIU6pPoOkvl0KdDm
2a21huLmU27eDn2mMMZzuN7fZIWWb6VtEkDGFXCurWOuK0wVQieEe1lCgrfIkBDjrxHaWmUwc2nD
ftFcXqcVnXSvpI5eM+8Jsyuyo99BKPtVXKtPM9oHJTn0TIXP+FKRNQUs3EpzP0dtwBb8TDOBAoCS
7IFAICYCXhuYGiFd3LCMg70FnuXu6LEFmZAtKDK1HQEkpWnleXoyKEoZxkO8AwoN34BRqqbX/WQv
qyC7q3H7VB0qUXvarlUFd477avfdOlGXdeyzJT/sTNVeln3DrexClviaLtx3r+xvmzvSgQ0OaaQr
ocilS/rPHtIMeibnBVUS6cHczAzEed929Si2gbr396SZlqdJmE/WyR/9IhgP7O23kL7e5oZU6jJp
6iunVidH/C0EjLlmN7sKzMHrYr59Z9WMG8SfSd0MXWHB4HMsfZfEhhX+JrQxRVsTaLAS81X6U/w0
/Ic81GwFSWi8R6G4OjMjYCQ+qC71Ci5KOTcsgiPmEExLn0sziMqU90Jz9Tq/xpqU84nRlcPdyyMv
asyhwSenUOVUn9ERccCGcg6Sqncrkj5+E8YtK79NHnXhI+Bf+w7Gu+X6YNs28idGQm3CJtE124C4
hSQRTify9zZdySK3lAh532byJn9QuPP2/2qFpKE/tlgEW58ulGa9KeQ8i2qqeDBZyg2hEPlW+EyK
1Yxy9ZpueF915ZIwFVYhrdKrBjMNv/BxKN2qXliztUe7Ln+1Y0v513EtYdPzv68781ZpfgxJsvPN
avEip4YVD20IlMRhGfL4IEC+N0J7nzzi1QRsreqMa98n71dmqxnUt5wTxtLoYtBFhjLXXMGadkMH
ir8zZzqtjiMF8Qdsz4kyMzqYBW2dcljwLF6ktIubDzqNYEMcBWA10jQna3RxfTFkdehJiGnNodMS
HkPgDg6JcyQbSxOHaLHhEmAH9/TqJh/vAi3B9OrRtdrtqU2tUzRimRg7pCqgbQdwcZrPoK4hRPGd
Xs/StElEbdwvg/Pwz8mhOWQW0cLzA7YPIic63cWtAWpc4q1QvTeO1kwrJisz0w80v3jfYh6V+3cH
j4oSc55muiK8OD7PVcXihGpHI12zMU/0ZUdhF7d9FrlfO1kBEW1yFZNd7a1LnJBtSg2f2A5uix5j
W4fKQ9NCt2gTgQHKJXice5sn27PnE1z66IoXCpH21nUrr0mpJ1taO0tewoHsNF4QObN4NEDNihG9
P0xtB1uhA/uR/OjVKZ3iPN4Tmp1UQTNdcxFBiFX0BuWvvJDbViTbdfSGB9wHJV2PdpCadNUL19GE
Eb8DEsqTk9A1yqhZj4VT+5hq1sapLjrc+2GI6gzJKNDsUoqV+h07us/OFWjmJ90YNbeC13HQ/FkH
aiNeo6UnW+JVU7bfyXSv9RcPqkv2PbgZeFSu/9xoHuCj6cH5H0zzwL8Z6KbRe+Rp9UO9zuS5gl9z
Zx0QgH2fgUUiOi05sFgalN648m1UDttzV14z9kJayhikVaYkLJjRmCo2RZCFBLLNKfgRDdvr5VmX
w1LSb00MnqJoSAzxoL+xXmKCd3M/WOFVd7/IIZo8pD4OxyBrFpPyq14wrcCjDpyPTIyhAK7fFDFi
c8vr5th5nfiBZENxdr3wOnGbaWd+oMaXyC100aj2tsljcyZOcZ8Ux1jk2dadbotc9v1asWftHmT7
DzUTbYQsF4LJD/sb6j8GUrvqvevbqvbSVqX6geHaVDJcS8TLeWz0xoASL+2q38JwueX46MlDnx0H
W3IjCbrnTMYoktWN+9mel0W9Ldm6IxejHsMIDgN4iFSbA+z9y9zmuHCPjstCr1bmEEYt6TCZDSdP
zz12NHVRtW5/pT2mPz0pYQBryZ9I6gG4ChqDp+2K7zpuyoyFWSP7X7/7ZHysKSd/XDr40OnZ3J+t
x0xBVQEVF2pwcdpu1+emWIEH7LB5wtbKy0YuRqz2XeXfJLTukCvpruVe4H/9V6WCoxhk5n5dWD0x
z6WsXDHGXpgop9q1iy6veBESHiUJqIuEKAWjbfbtNQ1FL3Z4fEJMMvIZmsaC/yYSr2HaGk1OizFO
dVoWP+qbTxvRJXrqLQ0LYKZ74j5w7Ph3CthMP/CZAHjGzUXnfZbZVxktwylwAE7ZFrjqccyTz9vd
CkDL4VWf5Shr9OAAdUYYWTE5eN6oFKqTluyM5L9/eAtzasFRdqWr0lRAqP6qb7FOqU+7ocC9LoAH
CeJNv6zvb++7/1wTRux3dvFM8Xmk/xMtzpDYfr5KaPmpkK7X+vGKzTMp6JOxZ3VIV602xD6ACjIY
99f14HMoY69EjHGI6Vm6XLs6PMzS6zuLYVLQkpS9oQ6lpkLlppkGerspCOHLQ/iNhpF81xXjwEsx
IHxDSv8iItkpaUXFi71urK/H7mybHidHEki0LKeHVCe2EzvlgRLi93qMA3L/hfI3e7d4I0FpQETf
tlAsD2KJFeaCu9kNdyR8Y72F8zSegWffbyBwY/JzsC29p36njG+1aMFGi0FHfwbTHkVzrl8Adwjr
Y/7ehBgX+INGv535X7dEQW6pjeP9yS88CLdzGshp6c2FA+X35a7Sn59HMgtg+QdPee5ZzuHeva9H
fvbZHZkyFwwYjO1Fl0GJD0VxU+tQWP03lpJS7JdiELoRfDgmOORUG5g2TAvCFVLWDq8eL/QS1ayi
MEwlpihK9o1bZVnONmrk3Uv7N34fqf4caVJ6C0cJy2+hMHV5ld6SL+5n0UVSSa/WFe/ejTAQcHsz
anEI8odGFKb8PUmIUhzIEsHalT2x+DhOw+uMMIJp87C6259oZ9+NpHzRcU+skKAFRWugk5KVa8ZH
kuuv5RVTXokrVosFjRVvGcob/9sLNgGLRPxpYNmJAGV8fuXN1Drrhub4khE2pwfD0XpN4E8shZjH
KWa9aKM/+gXECk6wQ7iAnjt9ZulsegcDk8F7sbM+fcU98GvfGMKw3jgZN537AU1xM2QvmOOuAxB4
P2affflMVDUvsnq2Il43Ks+RyzV1a6OOus0JyaGpQ1jTD7k/eJsNl849rS8K3OFeXZWxPeF8qjQP
Ydy3eTLwJjijB6U0aIPJpEGjphD5dq3bpTP6dUY2xQxOwXApqFx4QxXX+4Knvaqd3HRf5j2sNAqC
7xrhuDIAKvJyUq3+7U+VG7wMxzWYEpR4r0QZ5P0WXR0bNRvLlbAy/Cx4QRo4e+E9k7nQG6/u4/wW
w6eJ0s5E66XNFcvy49g0rQQHSUwZd3es9gLD+tJeKrsTufOZY5yJSdB7JG9qnxyHLd+EhH3tDJ69
oHzLLbA7++on1yMGc14r5ljp9ze2fiWp1dMzGmEJA3D43wd5vXSxaGea3RLKt/W2URN9GFAxoQLX
vRdwWssghnH+shyM0PCq2w3W3S37U7BNBX8Xp1/WHzOlIgvjTKmeG8AoMXOVDTVoatpsemSmH5aY
rsCIXWgUbzIgA8v1t0KiiXBfkAUCWKCeIBCKTl38UbPtHqSQ4DJ09qxbFRmAQgolt3MRqi/tlI+a
crDEOZzH069Dgo03t86jU8gihdM7Gts/OlC8NS9F5PX02qateTn6iZq/2lXW6XzYSyeBdwYChyly
YjEhPtEQas4+Lpa7/MqXB+r5aP55qy+lVg8Jz++RdDOExMSNIRjcX499lwb5NWL2mnYYdmC1CFZk
qEai87RqSOP1fhkZTn5D8+YgmUrdfYOLkw2xUiaBknlHzwERdzLBgp5pDMzHBkYUAmmz3vxK1S+e
D2k3ht5fTlk2PhsFHpeZnx/HB5pjuHw4/dgaXhTrVPTbNQH/tyZGhP1YKrpORIPpSQtctejYnphH
snDkOCPVykU6hMGRDahwOToZjSNO90jXZNEqGHKWP7laYJLLPyN9z7q0eu7u1KmkOB78dGHlP7Kw
N5YMVJZvQwNxyV0XDKa+pTyXpa167+UEGATA9ggC65o8lT5/fbBfurP/TbCk4qzQ7ovOVp2vI7Eq
AHnpjuz5zuBy4O8v/ZwUI34GKfCGbgGMqXezcgCg/l6WjhvWIbDLLqWCPxzqCSfwlFHw8PcTCSvH
leY0D727NivQI0FnbCgmgD7ZGt1os+nJT18rDL0ki4IruOs7uOjEulZk7I9NB2EG/YMmIpLbhAR6
+EXkAsnCd0vo3Df6wtee9z1veYpW9lLeU5WUv6/DY6MRgyGz0G4wyludzrZV2XK0sTx3d7BoD5od
Xj5JwplvbTxp5ocn8nO2ctoMA9hMXASu9RnHHfa5SDKpvvVzXs61E4ATanO2sDzQ/VUUnPFJ1MXm
LQM5bTDHBO8ovw0COuP6jC/ZDgjc3ZieIjv3vMjOYARvHxJI6SajAlOJWVH8077AZMwd2vS85stM
mrZcsfaXH1DQgVWvN+HBBOXbZfiSVw1+pTSjIwKoXhhZxEVXn3bfH6+2JUul8ktGnB/i75a0UNow
KNQMjoNBAhMvS46yKGjxg2O8QGYx+FVyYPCyqHfcrH3MN4BfOmahAcF6hl3mc+ai7s33XSKLZdW8
O9OyiDFQcTC1+QgvTfchmYx8Ie4Do7FpBB5l+KtzEBjW3fYmFPuOSO02+XmN8smul19epabdfhr8
TKnwQ/F/k01Snv0bhdLYZiJv62B+P0IM8un+ojDczYknIPN9gmjH/YS/xgAVRKDug+5IqTJUVjtP
4mP8gb5K4UnBZ92r4p+Sx+16TbT3oqr/STd2t0W67FXSgSVg74oKB5y2Oxzzu/+npxJ3NnVRjFEx
3+mxMqs6wZaKL7FtopWkbA4H1P/xOCPJ7ONn1bk47eSI8nJEzT68+6raum9uSFJxCgnv4AB7Vxs5
YgQpilEbMi9SMMXiR4AFXcJW3ymyPNDNSRM9NwL3KZ8U26XhwAwbBqvSopSWA0uUrtZhfht0Kgqa
aPWlnSVpTrZB3v3vAM2mgFtH6t1mPZqZuf0hQMWpw4y9Nrk7aax4tiL7cI8OgoP3B7+N/uNEPBcM
VdxpFwm3z5OLOY2ssmyU+Y7IiKi/s/uuRlXuzqER53Vq3UzKRtArFWw6mxBeOp++gEY5OIHUWo7A
NLmceVIbXo3J18qesartlA7uZLy/zyUTp/PRBaW3Q+wQZAoy+KrWkeVyTZfZQJCHxiqkQdprlsmc
i0RHp9LJKTNEy14/SXh2OvUlE8fNorALKsxNgoJ2QnxJdMvNFYvzv8vNt0g+BX7YqlTc6kkm+OCj
xQOLB9Fb+ViIwFMJcDP1/oyQtsfNb7QkbtZImydVTWzwNPIgDwmh4mIWqhkhIUccWl8LRPUOTPhe
oeSVraRN/CK8hImlFEqykDUmaKcqcR6agPdGK6JYg6FkixpYMCET/AYfX2JreMN9P4vC+3Afl6w2
H73CC8dzPOdSR288uarmEedUENwb2QY+pg2n0WTnJt9KL4+6+K3vhmsHfKzuOrdBtysfwd7JIT/E
dzVsx/X3Q6x3bbNsbC8QRXw9dbndQv62ApOPrKw9JxvRi9TlvhmDPvOOHpg2B71XgmKp+D+gCnPS
R20pZYzICBEfBQi7zgp6Q9q9cq/YKubQfemLUNGXvorSZagYz3c8GZ5QUaytMsoKcRPSlEp4pu69
y+v+G+nO8pk45sNz7KTccUUHYj/csCHH29BK149RnyB15sjVhzpg0CxIAYqYr/207t/y+6ZkKQZv
Kr+H1x5eBgm9GRHoeGE2Y/+zhZIFLwLgPPNUWHyShvuhsAdjGaYKzy/3jUq0sqA1+oumrdK8exJn
0LLC7CGLZ5m2dYekB0X8uwXgDHzINS5F2wHmGWdvRYM1WmJp6C+tOZ3UenxeSwJeXro8A5PjbYMn
qWmk0GDXFEDb4wii7GTrf6+R++VvcWEvT742G5zg6wpURp/uy/iaV9vdrpDix/hM8jjT0BMZkmuw
Gb96vtWcxxyOmgM6Jy+Rxofc/d9WfSnI/RLSOyuKo08VEmiZR7CtwantQg4mntguwDhlJm+4N15M
0BDsVXgH516D4F5xOjuSbydTA03hO4QMfIIeBfvOhVwf9OKqFr7rTrO4Wj/RxlKv4UCAm6Jxr3cx
fjbA7K7rzG0K/g+hbhkDsYRJGYNk+4STVnVvHrPoE/wiIN1MfN5FQQO9nn8TsEWJr6K8XVhDnIx3
GQjSJvB+SOzUkKn2YAGYVmwggYnN9hUONbAqu6YJXZD37/fkp1RnVSxV4gILmPwldLAYmjgD+ADD
2LO2mwjL0SzpksgJXNEals+0wQRVT3IF58jCxKz2ZFYat2/tzlmCVIINvYA7CFcEhAolEhUOXAYl
eKqOvgxOpYjJ7w9ya1RzSXMAtoblsPXAQJotL/AqAgyOwkNiCxpV644vWwzuiyQSpvbd/oLZnmMx
BQyIqJai1hLfS0fsOsfGp5RnT9qDAAydFhsdAIlZTh3lLt49grTtEswBaITQc51dy54vU8+WdHTK
0B7nbMRkV/ZJNKTDZeWjXY0HpH1jXiiJUzJ+VjsWIw+hDyZRNit7qDhD1PG9ciPL2FyF5jhEGTeb
7/g3kIYRqbht9OKQ0iJtbEa9JTfe6i6qsNjbFSWvMVF2523TSL+oV8uZDuyOucEaI6C5u7btgXcU
etgy9AdM8tLgWOiZE/3+EZV9NZpOsPNkFWta+VdjlXkEPiMC3Pa6IfyKXmbRB35axdxW9QOxFqKE
k0jdvNW1K8yFajDm9MIcoBqXftZ+fQkjTYaZkfztKQUJh4jFBgjpzRj+DXNTup7mWvzA7n7xyYMw
e1mGCyChj8Q29LuLEawZrASxp0lM76o2DXiA4jh7YxBQeUG4Lb0+fkq8cKv/COJv+xWAYthNnQns
5Pp97t7UGEKxQ+WxtzmTWF+s5+B9AaIxjNNG0GgNrNlqefYvjk9Ebf9RrLHoLmB7i/RmSaOF1HnG
hh8i6RXvANkzA/PAOij6/gIrD8cqjYl4BUi9XZ2nYuqLmwXTVGpMTDk8c2R/y8hhUBa8604d49GH
H6WXnipBGX3fedUIyHjxJTwx0bzLdMBSq5MGB8bo7eRE59aXOHxANNnLrbJsvo1Qkhq/A1R3+cNR
vRt2o3eecl+VVrUJVT9P0umX/yENTmAug/5DPqw5tOJycGiw9IX5k2D90fLZwVRmjDlBwzr8f8WR
P3qiUWPXhmZp5jYax2jGsXP0tZqHA9iW7hydvIdtidPMlVNBs9E+kP9LDTDYtfbaSPQ9mbc67ldj
hLMJYNleOFmrDZ4SS7pV6KZJjvy5SAUpovJsTg4Sb7hzrs7CX0FDAVbTOrl8v50f4ijnzEKD32jk
fpycER9Zd37LXSyCk/IDQS/ieeKNzpd899k3N/ZbM/YeUfEZDARYfzFb/MShMWnraFiYYNIjeSzR
1PrsUWU/7BUFavrrZmMAsQCv5dwWs+P2qtz9bNUw9bXezAYd9d8QELb5VJjOhABqf+fVu1F63N1d
jjfKm1cChT+8f+BdwdUdmfBLfy86zPecqD2mIz2QPay2A4m4jzW13FGDVRO3HDqXT7Ro2KwV4SYc
GeyWlZQYxKmT7ilPocOgrTzJTvD6lZTLhU1uzix13Zw8HZwN4iuZIObscFvzPW86eEtRpMjbRiHF
7ss62DPTVu/Yid7+SobAVYPzKerO4hCFgD03oPHKqZXUQE9h0re+PvEZ0ZuqCGX5ORGUOSCpGAQU
d+tXzfX/ekD6EKIUDiHBmkNZxN+jcHcsVJgwEKO9gIkYPz4sbIA3ALPGiMmHCfc3rsOpocAdzdI2
gL5upP7Z1hmy00RG/r8Ker6M0X69vtDryv/vuj8ftmh7aH6DO2gM6OC5JL9aU8PogP+nyspuK266
7+6QNHM8efiAHnH8b6STvnSVTorgmvE0yEA+vzBEECrzKqYscY1qSZmehLlv6MQShXW1kL4KtWfP
ZfmQBd1G8yfiExdJJHEcghxG573N9BZccxlA+kIlf+OdEgb0A/0RfMsm8wiV2+KA7qXTwaDyd5Sx
uMC+I8HmRSPakRqKZWfoLe80kEbVCeeY9YhwB7/uuXPNtC7G4b5BLQmOcPhkYzxFObBK67eltDsZ
VCk0aK2E4GEllWIev7dAjlvGRyDg3Ws5nQwEQUqn249huvhUNcUitblxhN7QEyKmYjJlINmv9SbG
qojlxBEVSAgqq9UpbWSaDbFdjdAiqPrpkNvQieoJc7muWDAImS3565FZNO33KPCAPfcERpi9mL28
tg+qpK1+YkZ3+oI+O/PGAVViunbkNJTN/I4YMRzW+CfLoeIs6olumHhnCqPFfTaGVAvedk+56YuS
qbuj3a4b9Bw8KVQdMZn7DsXpoMrG0GqAx0Ym0JZYUncX3LhyhCZLPhsNIwuHVeokuVbeKrKMWjc+
aFU3NuoSlsYdN9N6W23oIYqQPnXA+8pxUromM3NqPiTOwgK8QkOjRMqUHK2G9+AIl148DvJJMXOt
WTxa3DAUXRlq49/Cgp/W52ljcySEtD5IsooCT6uKy977aBNMLpN0YjEb2UYos0yAUg8fC3mdXynF
+8xLpC5vhBPCMUGcuxbG8GMLnW09BiLbPW5mg9P8SVERMV2sAgikKVSLZXWMEef5HMZcLPHjYosf
eGD7015DCgJu26HnYybT0VLOD9do+oV7OyYG+UtuFhZH01ZUGbXzqz3IQhfR9fxct1Sgg4V6f0tS
F6OApahmlxPb+J+ct8Pl8phgY7Ly4rOW4BAftxyVYEVlUUXgsxrjoLmQO1jbHP4uADgkYLzcF4X1
H51EBdYqU/MJVHjVi8Um9cIffSr5iBFNv6ZvVlp7/0to3oiTUA5Zn1gUcvTumVqrfpNUdUo82XcL
9Z0ULcLEbIIkyu7p8qiOvZ5M+ydFe88TnOHUTQTE1KbDqf0fxNzdhmyI68faM+/XfAUR5Wf/J9EN
HUk/50k/DIa5Eo6ssfQnQq5pLAN0Vv3p7s8ENQISsJH8HSikmuXOfUtGvhm58FbuIi877fyE6K8g
S0SXT2mW6OO7SBZg1K1K+cYPLsnnYyWBJWuSU//3pNZU+u2FEsLXwyXg8pqBgj/h3B+3E1MjN4ci
hNcGyc0LIqB6DpTTdc3BMXXcklrdOP39JkrqfEpg0BfgiORHqJbK9l5C7nuiBQlKGcWQHrfZzpzh
yHmu6JiuGkjwv6hkH9swVKhuJxRE6AQfd1AtitMOp2yg+VdoUOqBUHq7B4rhJyG+LFaOTro/mkMR
89j0CQ91C3W3cjcg5vWvmjphoOjYw0NV0hnJnwL5JgiE5k68WlsXw9oGXj6PY4vJeb1d6M5v4pDK
WcJC34mnxvupG3UW1cXADvOWS/pO5fWJsLb84vsMZ273OozYHhvdcyK18TiRiZHVFQyq+x331Fkt
TSmjvfhHkmTDHQXJx4GG3czaBsSifabowTR70r6Fc0sIIaN76FLiwmuRcVzGrB2NTNTrUL00Ioxt
ClKsV8hOioZn4v/J8MJ/Hz0zLZde5FDK6VhpcBqD0GeeBYlTr3XuQ7mBo/bQVI/2M2ix+zFl9bvV
h3DOVKdHmlxtKfsCAhbD1mC2+whHiwa2hlgTYgPYH2WBFhosrJ+02a9lnEyLLr88gYHCanfuez6U
t1NQlRkAVdli8ISiVQF4mffgY8H/TFA4PlQptRfYKgWGUof/lrh4VIwoRm0DcA/xJD8qjZZQnHGU
PvVD7vyYFLSBMbAVppkylnSwWURmTL8DSnBws5pNC7GmAZDSCASBnZyORWWLaHWkt6PLYk0bp+oR
RX4t0vATajJjN5adq+CTT/iJk2OZCSdIrYuzNvs2GvMe4yAqvColSvKU6YH7wFvqWAySxYsfHOMd
sXKYX3uC4cgNqxWNVKWtDbSROIoifLOejSEWwDq8gEUxkNtlPpU9g5o0YT0VdSaOBlIi9Jgc4n1I
FGHIgxMQPtI8JyP+nVjU4z4JewL1cKY712t8tJHmZX9fZ7P2nAEFSZp1WJmM8qPjClR0d0AWNRdW
rCtA/0BPS/adfyBPetkay6x/06VrczucQCuUooFby/EPqaNh+wipjcMVQ/OAQPiEAyOabMdPf3ts
ygb8OFYqD473AzqdFdU0wSokYevUt0attOugEI/cKk7uXBV24Cyqi3r3tI4huhH9OM8WTt2sVfM2
IXYGzOd7lwE4+4bzmzUTdVzbRU3Hcmoo4HMsYB3lh8JL+4Ywy+GctPP9v1mMWMiLd+6ngBmbvzrg
j/f60Orc/NVWnUvrsXMsz0k/a5jn6UR0ZPwGDM1hU5fAgj0/BuUo0IClMU3F63frNFzRw4/oC9Ff
BJw9iMJ1blKiJxeg5hWd5RVm5xfrHFAeSxca+ta7dJG+No7BWCMKJzXEW4VPdXnHO6znBjT4kNr4
+kB4vErh5louI9p5tZdBX5ZOkTqxd14nuCEKMh6aUDHvINKRMk9twzwFg1Iv+QURAsBLjMDF23PE
9b4EFIYwVWIxGHJ7GRvlpARFL9M/fbU7e6LdWjERLJozscnX3bGmdYFxi7o1n9CYwXZZBDjrR5Q1
c2AujRs2UIXsgmWfTQxvEwMWHC80CmuRg4lfp5MXOuF/5rLZPcbQrEniazwjSc++Yd2d26swdgRJ
52nQjoNtORAE6qXCSPdC3GtBQE0Tn4Qm4xdw7qIlK7+kNfgeNhnsx1BtahdIvUm4wtN7B1AKkIaD
27iKGZNxpmT+TE6qy86LbRn14wfPJSjZQkug+vpgK01KTQ/hY+4AQ9B9qJ7PjAdklEWsBjYHm98c
02l3xTHZ9q6LWYP3X4JLfmNq2+tayirigY8UEiu2qhvkn/XhU9sG7xlRaSzDj745ZF5jQ/F5gmw0
gwAXtw2V4DN5dAuzacS9hFzmC7v2uo8e0WTLWxpeDbHMERGCGF7IVU1xk0Vixy4LIjyOM1ZO4c8h
TQrdj8pN+5LTzn0hVgz0VtM+OwYqv4hCFv0SAYqw67GxLJzJdOBLGItidEZZUCqbnlz6hHTGK0Z3
acCc0HBzhyg8G767qmWcsC3AH7ma5LHOd2ZHhtzWC9qDZgjSw7yN6AJXY1uM9G8cshSae8CqMADa
SvdsSUonD7R2OWVyGQ4SKuhDOPwWlW6z9Qkfpw/sMNUJv2GNSIYj2vA1ul6N708Tzn+4GtTSmSC0
mfB8eyCnFZQ5I6QjdtmTfS7TKDTN56x880ScLUACaVaqOd8Epm8YGl0uj055AdTGK8GtOrNrbZsp
k5qGsR9LbdrnFv/RyxkFe9MxxCXilXUL4WVUCw9tPUNYnNUb8ecOb0opqauHZ1RGPUiPCQI+gxqV
OprAOwPvrq5TH4xXkCW/I3LGZDNZgrrqfICxvBqHEoSRlyCnEGfoFQaHrWyfX2JuZS49uHes18Ls
OnLJS/5rYmuksokCHJBPraxcF4Btu0RM7ePR8K8mkpdnc4GLiv8DNsVvBqCJM3x1Jql0BL+oB/u5
8z+Ey9gpR3k1LgGJFNHJk9g+1ySjorvwGe9hQ/us26n8JE9b6hw6c3MtkRdd/VYUpd/l8whc+FMp
dVepDgDaIL5ZxwzdjmgXIsywjeWc3XOhlbOn/pCQ2aneCe1ZjS0DAYr+L/5FWCDM+iARieJ+YRkj
pGniZLkK3OZu93XCYoNy6zd62rW1GyRH8sCC2Zyy+OfCaEmr1EG4hx3I2Q4Pgh+qMFIPWSg/5YYC
28/eHCFo0zD+OkuuTDOv6cMp0Ve4x8Jna/Tfm0zGA6Gk53fssH0+/+8P/M2dtXVBbdOfQU1OPYax
hZUm1vZKMEVbnshNRHLR3Ejpt3walneXoHGJReqQxTeqsXBFeUIXg4Zs7xzgI8xDGL1QTjBLb3eE
LLy7UNEhSbrBEoZbOvztv+fOdIyq48kVXFgiKvyP00UoIrS4MP/PADwuw52kYcm12OC2gNExkPPe
b/5xKIrek5quj0SVmRqnztpKY1Pz9uKQ/jzNFfK+bCwPxdvO4Sa0pMWtQO1qODK48gCayvAu0UyZ
kjzO1q0h8JDyghgq7OBWYxwttSTEREaQ19UzS5RmUdWiwxlX8SlustmtSBE8+2NX090cUisI+TKA
4elqvO4JI10pxay6qYGSNaVUY50hcyi1plGgZA+lp/F9XFSfw624Sk+8DzgEGBNYh6obo3VCa4sD
gDMuR3vAE8kcL0ayO7ZMUg7RRBVm0ZyfnbG2iYl7BJCzj/TTtkhJKO3m5w/hK+Xrf50gFqLJcoZ1
7w/tbRZwsPcXlgAq441fFD8uDOfgfMQ6gi5SFWRN5s5y5q7tZ0lDrcP+kBwzaGBSIDpGs0/pukBE
sqr85zqOKDKK9seZCq2mEDHY2PGD1msTGRGsywhmvE0I56S02WeozjGnKxBO7NXT/pnrj1VjyCzX
DIvZP2HrJjHppjgSnz7/1MJnLrocNDX25Rsb+W4liuoocfCDBqhJzx265mL7e+K3xMzsysSG4H+p
34xco0aQfekApIIXDGU0e7O31oK/DNd4/S27Y2sgbGLP4M5RC8jV5sGSWKQtPnq9jy0rlPh6xeso
b/HDlXsM7VTsJqKx9HDpee73xiz8NwGauGKYhH4vPweLlD+jjOS0p31iK+EpIk741jK/RaiCY/mX
imsXQc5kLJiZYrGxIvN7OJO+mRt8EwudlPF+mnsdM1G/QeAzVp7IGmSMLt/6iCNCpQrMhqEFQHoc
0agDotpivySvVc1+R5mEyJLpED2ZNDGb7PU6cmvjIu26EC/q069mjy6AUOCbuAkRrue5ELPgU5QA
1huCJeE48ZcspUDisSXj3rRccM76fINaU2ekhOeN5HU7zat4nPgIUhWx+V6UdXxp7omNsQsMUwwp
9izPUw+LyLQwIN+nlExQQqBq9kLg3g/Lzq6Gqp/3ZB2RDLBem/9j7pfHzgYOTb1Yq7wKwjgOpVs+
dzWHCDEOacKZtnCfZZXpFFcJEFc8ZdQJiKTtpqZYk1xlWOBvPd0vznCzYuRNzomTYPKedli/G/Tg
JIhLflZ70vZ1kwil8o0NtpMPijjgz12JGa3H1hZQN5ytEl398C98olgCjDkL365Nwpogp0Ym5iR5
0x0tYYO4FpSbfJd/4ES8m51DiD/dpTqHK171npAeCnNdHbLG3cD3co0sKqbTcXcqiV32dduZ+aJW
xSeugW9L0X4ShueAwfk7bE3M+NceRiQB7YRHeQm7gWLbroGv+47sJv+1JWVcFu3oDYd1jCgHU3Lw
vYOVUXCDbqJ3aoERXwhkwFuMe6eK+l3d+qDSaAoOyeDeLHSGQ/b7Y0sL5Cs/mby/vskNjQRAROhT
4o55NrlusnfpnJGXX8XLQ0dU+cMdzLe9KmiCSfCMrgey4u4TDUYprPZ9OObATBwBVZ1/gUCx4cH6
EVehmd4zeGyNloZu9THRnQvLgYeCwJjZtEsb0EQGRGjCL1M9Xp0a+6ws7e0d6HjNc0J81/9sClGm
QzGF8ZEvsxq9cNZyFaPKwdohoWvsGMEHWIuB8loU8jsZxssz6E7fEaquG++GS3K8JNxwnmOJIuOd
eV5BG+Aw4NEmqZveB4mDZf9V7Y/qjZOx0StaGqAMr4DyEjMAGt8McoBPiceXUVXl+x+dD4WoSg+l
wA6HpaBLO5i2gUGebCRq/JG1zq/uOJvbSvF2M1V9KgsVnyou3Sh71uSvVkYz+kkWwXkIMNQxJ+G+
edo/D0L/oHd83bIsq+hzXdgLlbHVmZxTbFoYKjxY5WvYJBiR7HUkedJyaRgfREjatQJHqJjMSfGe
SR/qRI60kIaXIC9eXcsWt5ebTrUmhbxsnX9OPlWr9r3SHovTv8IuLuLE21o2r+GzX+sQw3tFSdA1
+hKZU7rnacXslqFEANyD7Cv/S/rpdZ04507yogo/f/P/s7xg0atjGpSB3TBNYenpG3sCkCk66uq6
+4MkwO+NlvbxQWtTkIZvv3ZrlqVogtI6DmqSxj5ShkDA2bwbUhaUGvYMNv/jCwrrXDFXq+dSYXkd
ISs0F5Dtc7Y6BEidPuntNLCT1M9YWzrInEDqHbpdPWMl2khnp/HZsqhdM9TPA4mTTXmss3gJ9PkY
QMURcQkdcf7GeF/CKoF+ZxAfw4semXejgGMsgh0/f5A8Dad+7Ml9iTC7Ds7DMaNy2NvYZMbgHafn
mWIpY1/93hhCipWfU/4p0PRYajqpuhWpfOhHySeyYmkcvRCCfMGM51xvr7TqouS926bQRXXkowIe
y5WBgHcOvoUpsLvqj6Y2Lj2Vp2TAr14PbKXqr9Egob7y67AROOqbJhoBL4lGS+sGceyjJPja+uK0
yRt7EpjKaXEn5Mm4MLAhcbL4NWgZFkI218uuy59O8Lb4H58edrPRoOhtpEk7Cm+xhMSBVakv+B10
SUrrDcwvfP/eX0shSlYPe0GNXzGDm7ohfctU3Nm0mv9u539Bsygf4RoDCpyP8ge3WglIAt/3MjQ6
ts2wVps7uAzdphz4G5GvCtw877KWhP0G7lYqXDJyTzi/I0hBAXen+foWFpijcoFRxtFl9B5geq/Z
fqXJPKq9SEDJWEmtgpb4WxT+YKgI8TG1RgNQWy52BT0l1BqG+CpW/+cJwnsyi9ULMZbyfFNs7Y7l
KIpbG94P8JV3HDdmKK6q79PWA80t9idsYtmkcho1c2U1pWNiIahLOAwbuK3/dUlB/i2xrtLJ/wH4
91H53tYchPAVrNM4xIBJbt77DGk84a/t46NjH1z0ryCBKSrce8UZpkaSHfxtNWpqTyW2rbwU0ak5
nUV0tPFmeR/OrRpiwMAVy/s3JbpVnfm/7tzW/bHn8Zp4h/LIGHxbXA2cmWXuLDhZALoS79292Bww
9srOaZ2CwEmsMCqG9LbVidlvGH2W0B6+Nb22x2qK4jILa2EwQX7GBAdYSUKB+h5hDqj6f+g/0tFG
IBtpzFiuVoEs3QZhmGH+h0vgKH8SvRo0wErxaqG6l1XncEMa77QP9I+wMtFY/E4q5+AycZUd1WJc
KUap+yDJU+kaemlE8igQqKCmiIN7btZBR1AHTzh5Tbg5oRjISr0ZSM3QSj/7FO5ngaY7FSqz4Rc9
vcTqdUN7FHUJHCsSeNMnQxxVtxpX9W96uRSAD1Or2+xTgSZDAVXkmZmKpBApHanHgBbGJ78J5S+p
0wgPLSoydZ7HmZpluBut9eSwSz0CPJ05sXEBuBcIwdFPc0L0IxEZDzxEZq6AhMO/l5fg+lcL8Ujd
SZdR8fmkspL5mH4MCNzbLDERFzOihc2ndjuqQnsjyL8hWTWhoRzKqSC/nc6CbLCGzLSiekTKt68u
Pt1KRKx3+Ta9gmBdiEdnBPbNPkIIhSkfiL2DYzHOQ7sS803j0OUCJxz4bZIJxeIIjHuRNVaypule
mX3khe+X1ti6KQ9ETjtluKaAjb9v+PpYL8eta+pofAif8dWQQh4iy6vIZgFMQZBWGKN8mTdR4jjI
q9uPbPPrpbNAUllRb6lLCDmGfFG2eKzvw5A2ERygGBvoKNqy8z5fXLssZnZAAR5Q8NFYAkyCYmfV
+D+fWgX/zK9gkBzXk0PJKSIaDD0qpM5cbViqrgQribgSj5ZhQw0vJoEiK+RQrlPTZmliaKLKiGkw
PvvuMvdQDgpUNnw7IPAwa6auyxhF2ES044mloD/N6hO/aEnnpv4035kOdElsoDuWlR8MIzWL+z/d
RTMVkLBEhIZ2GO8ARJF2CRDn61Lb1YWg/5TPDyr6ofd04vbAI3ZYSryl3/mtIHJGWD1jcc3Hr84r
iAYRQYdWh0q3K4R8AWPpDlyPrnXlgkXqJPGlJz9ibXA64pD0FNZ1XzDlp2LDROqI9+AdfUJ3wSo0
2zBUMTpJlDTMsrY0A3jbdzapZirRr4Bfba5q4P6YctErLXPqc+7sVKcvZS0o/u/2vM/6lYH50Zvp
egCoMTSOdVvIj7LYRbYfxJj4HxLCwIPMb444M4YtSxOjKzsKp+jIwT07ewjALn8mxIMolyzYqXAK
L2Lfnsx5/SnfEPcI//kzOnjdVUBydt+Da6L5DaRf7kbkyfFhX2TaVoS54/rwcoU+43XRYsht4m+I
gqnXhctvxq8KnfVkdPRmQ4BIGu4hJ6WlpPdmGj4fDR2pVzt3sjiBq/5r0hWh8co+g9gYEN+ahhVR
UGTZBWbtFyqt4SNCYJ1lHvkrVhK9LhGAIQfcfUHTmAHKI84mdqQuC0yaqpdDI71jH0SFHpudfQbn
15dEW1cVXLe+MmNL/XcEH8iQSY0DTEa+OZCzYkXuo7WU5uZ6JsdECBhB1LAU2tyUnkic1uLclPXQ
n+iqwdIcC7FqzQHd1wuJWp+tAI61nW8rTiNbucgNeTquvMS5ir4yrPqvy9JOILI/dpWpLnVvVSzX
ADmK82ezwuUNj9s4aoX8DpRVfBlw5BtwyekaJUGkJmkEiIV+zVYOAey3ms+JWvs/9Qb7xuYGj5o9
x6/aIzjNaqb/jPmYVaJzp9MnNoJpbCn2JgahsHODA2bAhE1Dc/43t3oECBLYwtHTufZ1zijYGOSM
ZXEbmMarNBP4W2khSrBchlYEAB3XTn8IIydMkPzgID5n2HXWFiekC25rJ5dqyAa3P/Bt0XyfJKBs
Bem+h3EYyc5DmeVyjTyUDRBZ7ztZ1HHMC4HpAYAAcoTx/E6ggnaCpXKRCI7BAY/o0uQ8X8I6jrKu
UG0PzCSSqSfg5dO7ysYhKtA/TngczT42DP/03iCpPgGgnZS8BAxD/bjI4X8UnmEyaIwiY8WjdqlX
yFZTWltp8IiJXEhHyBwgLr+DVyz+gfUy/NuDzEXv1iIixdcKzv6/WzwPjvqlObnmZGDeMxuy5bEQ
Gs8qxH3AMb7xTWamr7LRbozUL0kCxE2GsPGzqrF/zGBThdF8o4O9OJoxIFCPmuQGeP8APy9EVJUf
tWR9b+P4cCAJ78IpmxhSJV3WSloafp3HwAjFsFheqtuy5D9oEgXEH5dGJ0S5wNomUfCqZC/4rOyq
JjtItG5iBOAzN4UGrHUR2dGV6PdgTlzoVXOgxsy9AyZhfSmp9kHYNgId8S0a22HnBhiuCOCG2Ik/
5ZiPIYwPS46IhXUp3aenMZt4muYBg0mrmOzFZTM+/LkJUFYWkpfPvyNDmUTX8HvC/qWQwcZqd3Th
VWyyDkJYnZKsSbfLQQ6W1Mmtk2kRJG7Hle/GWF/KQPQAQ8LJfOsmL5guUpVqzc0kp9ZuStd/SZ74
cJI0GLtWOdYXVe5oA7t9LgPDbs/oKbiYFls2YTgEyCfTTADH+343l6rVk5T55upqWL4QPBONvM3f
NUHzAkA8FouY39HX1aHNbAbG1NiE/JJu0hxtpvsUmp8V7wNkakhQy8C0Ij4ch8iqTIZrgm4PsTjW
ZXBqHcljXPFQDKHDNmqqhD62UvebdGozdgj/oNWY31HLuNe8cmLIg78kQstqh1AR4+Yr7XbCY+8k
dOMXdVbePwr+EW68yB804LVW5IRsF91DCFqzhu/d74zJ83poHd4dOD1adLo/HSsdADUvnpzrM/U0
CVK75pY0LVGdg+k4PW0s2oTLP09DhsgpGJ1uzSw6RN6Jy4QFMIk9XDqXZnVaY0JwImMT9begyiFC
uF8PgrR3D7KJt/NWpAwmVo776TCXFsviJVzRmT2GUyAJDrcfFK+WQcnSMmdVqWgB9lG8jvFAQfH/
UnltejyQqwDalaYab/rD0rN4rFlA/CeXQi5d/3KSP9UOoe3V40GisaGJs/5Iu8gT9LUwXTvgmNGh
7BGmoHmIGSynA8B8qV+5xgayYTGVC9D1MTijAuc9LnRnGiGC7ozeYQjbEuBxc3JfDo8tyzNTO7cS
r1+h0MEJUjvjEfdXS+ASrWLPpQOIqhNLrqSQqenQIrRx07Vzav+1o60leQ0lqSlkM8NDNTZQb4RR
35hq9mzOlV+9LO64BZFlrZBA25XR3q6hA2YOVc9k/5VB/wqAgPzmKRiuVhoC8H1wXUOTaQ1p5pOS
1hQdwSOH7qTho4qA8AqeoFlZzZbZ371RnpQc/6dWVHEFbsIGcFXf/HpIG3Xn5w6bOEKH9z5oPPog
mK2H1NGA/kvLW3WY+s+8PqR27MjCMZXFGorah7IPN4pPXS1gO0TYiuU6yRnJw47Mkh/LAXgl6Uuz
3UU2dJn88jPl4Uhax7/t4GB3lFkRSLP6LX9GEIUfPUtNDbqq3aFrW1IiydbrNenrdYyAg4s6R2X6
Ciql/X9rbTiGnGGjv0FPi4uAMTcDoR8Rwv6zOaRY/Iesi/O7rfoXSwlLDuaLq94s603bv4YSZj5O
8K1VvtrraM/eXUujCPMHk+SEAMiNuGQfF5gyF2izQJUCVPnVsJc8RPiwrrLd/0dUeKA5mBsErdW0
oogMQp1vSu6WuslfxOQNi5UluxZhzNn7JPTU8x9injc1Ugl1AnJtMHR3TED2AWKoHF95hHs8z27B
y//s/HFSFzr941fj6bu8TiItXg3x2pcAMM6ujI5vFAttxfGyKHn0U1bUEvJWx4FKKf5kKlkqm83x
0hEPM9di+85wsk2wTRxn0ACYNDtYjw083aHs8M2syRgsXGH0p5h9tfz2LXtdh+Ahw2aGMgeQh9hO
HSFrKofKHg0rpuFwzGI0EAXPeCf3mYxvu9lbIuc2sXI7R57RL+5zQ0P5APg1B2rkmQOYuuISnn7Z
D7FdzGbQtsRTCMKqEhdcCj1pjguuN3ULpF232MxDvksEMWZpGpF+f/DRWLLNadK5ITav8as64TTL
fGhA/+sOohmvI/v7V8ia/avjBa2jJKmdbfM7QJATnZBzzpdCG9VDwr5PQ9UNItGSn4cU9BbVsnpS
U5318lFgyI0N4pP3JLQWsupFdM4IiTgmbeh4V9VXHA4HHik425WZN1gERobog7qhkwXW+qtex1rz
uilIcRx7F0OM6/a8KeG/r8u9uYBmYzv/0a+HNWbkzDgT6ADCg/2thK3/IdLe5jcbWVn6W/Lci19p
q7azBmORWzV4F00Gv3AXBhd0qEB6zuDqMKn5erwqcH7jDk8E0FwwtbfESrTXUiPsptMmUqEsSv9h
y+BxyEujtCJoXNThA4cxDNRLES+dMlpdv7aUICDdaphhr0FlcRpvXSIEIw/IlxLnQoWN8h+XdIXo
3J3PlZ+1F8TEFzLszw1qmMqh2Hdmnd/AhJ7uhn8Mo2/qDsT3drqp6AsxaEL9DgeLiG/SFW0NQ6tZ
qU+qcU6kcJdsEraA+mTAkrOU2DcigbcniPlIyP2ZiPEgmWJCIlHpcJiLHepfB3ahXIOSAd4xB7EZ
KxJjQEWyVY5pvTngdANhKKTkSvFB1jfltTRk4xmGGCUVShZq0ENq9l1xIJfG3kqAc+jzKBhs+um1
4StrtDrfzt+Itz0ivNppDkijQyz9VrnkTkhrA4sInEKAc8RFu0MOhAq6s43MnwImxjxDLq2RW6ZE
uAAd0ZVw7mRy1C+8mskldYHxlnEJ49CPCsWBELYE1Zl0VpDLxza8mzape+juIgr1BAVKKDt/yQP3
e8dansHxbtnWcQQD7BIgSZ/sfyR9DysPVcktX95QFVKm/yrg2Ed0wsY9eGOhJhKj+EIBh2WA43wI
CweEFNDFK9/i+58B/GJQAQI1GiAiLsrkD7FvBpbeLqGuENtt0kubcBFbojPqm8Z0Pna1ROBajCJo
n83CH7TM9F9jxkixpUCoe0w3G0Q/P5ZXfeYdA7qCqcMfztnYfH0Nl+30kCs8+muBinNstN72YG7i
jQnOPzmN7to2hNS+7OQID8F+0ps7efWGGsWxmW6rLBP2Q6v5GhhUnaU8HkaBaDRtcmadepqipxou
Az1GfSBCR2Mgf4Bv1zhdkUqm/WVgExmjaemNg7yxdzbLP9QHQiy98jsSHsswHbfqYOqUK6LIhYgO
yNhDb8f7Y/XtEEdBFWG8bztB2LmO7IHAc927bbmYMKJWZwlwp6LCSegsZ8xOTuphmm6luhCpWVTr
PQJSbm0T+6Az7dFuueIbIwxZR/UDMQcHVV3rFShB3J9x0BTwl/9IHhi7WnGY2ByPLB5Q8by8AY0g
AxM0AZ2IL31T0dwk9z/1VS1ZShBk48pEq3BCGMP7xx8U8sKbKcfsf5LdGUVGY+AbollpETs5foT5
yD8qNP3n8Vt4GFh/rUJWeyY+jLWi/aYYfmMcYFQquF59SULnCnVErXSauHg5pmI7TXmwYpu7neYC
kO9VFBEAYMMlqm9z0auhVjn2hD/oJpPRBNb5haBxGGVIkBXl19CrKwEovpC++p6rKiGJkq/U021T
PJ6AOhaP9xqc2jTcwe2uHB0NPxX9KBBmBu+1dyqQmSLwVYlgFGwqtNtKCwGFv9EE6PetgB1Wyde8
eXrY3ZIYcYGBB8nb0mEMnJrNHZzsuAv8gL8Sk2Nn1TVOs8YBwes47KrPu2bfNQ+7LWMKPHDKrQoy
EQtZkwOl9S7bIOG8iGw44VPcA3anUtWSzvWoZOLn6z5NnDnBPqH0n4+9KFnlL4ab1I+nRPwrO178
OSBtl6ctK/kNLouDKt58e0DmA4tRnCxCYkDXG27ZS5f+eB8xSzgp7NxLqM4oTEt42SYidRwlOMrd
TMe+US8CBUwTVOfYLWbpLYthp1V1+R1hUIXr2HkUzntIcsW+SCfL0ikYTkEmJDNPSlCrEBO4uV1+
XWOOM/qlqsXPf071YIRFnIum4KuYy6oSULvNQmqfiO8AE0OqEA5KscJzttW73y81lDF71DXyBSrx
BPJ8F2OITYuJF5YqXoM3fCWskVFMV9eHqBVk+CQve/UtJ1QykPnOVOx0LLCdV9AmrAS6q2OTKQCm
Co0Bw32C5nliAwApeJe28kc3tA1G1mLXvAJ0DtR8qNx6AFXl+wgimQIhWCTioHTBTrH6e2rvpfP9
pLokz2uHuHo9EMQqQufM1/SVvyQbcSAHFFLf4Dip3dhmCr+Zc3LD8JE8IK7XyEB3iDwCjrsx/w/d
FKwKlf3GO5m6BpcIuyoEuTLhYz8MeZeU33++SkTO0scdoXliS2Kl9bQZbqTEIHTxvtWmzZq5YDkY
NYk/3xfrx2YNQxpskXigrKxKX9yeL7fMouDef6HCUbHMkv3tfrTIN3vxzV/FhSPXviBCYBQ9bt6m
q9ptpFXjWioj4HciOpvJs671WGAeif0pPj0VgjOrPJFpiWKhwj2AtxvIRc7atIVQv8lxIaVORQ5B
G+l8D/S109/sPX6giuVNYCN/ohqv1Ev2U5Qrw19GPEp/9baLadW745EGXWPelBRJKYoJMBuMiW8i
2cZ6HkFJHfyVqIhfeyevGBEYgtxj1sQUttQnjWbz0StxrjqhWYagu7TdLNqE5/53QeVVmNynvmah
mpjRlW44GHVCwPx3jNksKxhzq31wC2gV4VyBhWjJJMLs20Ok+FBtjl4023f/SwK+x+2eTaPjVpaF
7cKgqNSJy3QBfvpk4ViZ9cVfH7quo6eJCRuZoLeDVS1iOGDguhax2HAhr37sP2X7NkN8sMujBlb6
PeOQk9K9qzTQcO1vnEGjeApmEvMpT9Px/YtS6nxbJpCQgr0HNPIgigoousgzoz6vriFpFv226bDn
z8rFHf0u+gixD7c3m03WyBK7/4cFP9SDORPk1B2u79m7sbPcN6BtAPlohnZb1gmM+0PNQ+E+Kd0z
xd0sz+eSjWRV8ATYr2EPvPsbwMrCe0vKPvik/Vbl9Rd3yiMf2GD7VIeVXbhvecdi3V63e6Y5NZj1
uGEKdtA67oUntlSayJKOLNCiXLi5nUcSid/pjAW+2qlNnB1WFVoEtlyJdyxhscvUAnF1AINdkrvN
bDXsLXLg01w62KouTvNkNfoYuDHOrquKyivagh74eLquyiH5zF259fudcIWzMu5ugAYipsnJfnIZ
4ioF493XUUN4DE0ZpszCICFVaLEtRp49j9pZdy2+iongyJ7CYCEBUAQF83x/lEYZqqtYMSllH0qt
pPgUykMjhT1F10v12lWkE0mSJKNwfgWjftOXdJtj2weVMdJI1kkP/FzxBGsWuWZ1bFuq+rIuI0Hh
gin4kZwKqcfQCXKz4EcbyBzK+3MpatQIT0tZ4WThBM3Vw6kkFA+l3yjNLgUbY/slUVn6AVeETkYB
iYviY0EqrfVvqQcSYEuBMvaug1TxciSsXq4GGPeEBu8Mz81TCdJRaWjV3WLc5lCk1ZhKqTH3Uf0T
x6ASy/K7edLJBysMZpTb2TxlSJaUS59ShEFsBWwwyOhXtC1aZs5cdqp0ctRWXz5sSBupa0AvIUjr
gUKFOM0d1xCefUBqry61wQnNhlbTaFGUcOWRV/FqvfvR6xkRUbIOOz8l+swYD3yVgGeZgpcDuO1B
Inm/cnLAQQlAGbvtRURStW4o9RBV+ECTLaK606BaeymemrASRR/7yakZlHpzDwfXNX4olnf6lj2L
tz7jfhQC6CSLxlM+75Lz/AppV2kBfw3JLV/fCFvBvAN8im+EzmaNNQz/mr95ZRbUdI16DYgpFgQG
50c0iLuiIHMUL0i9cwle3QBZFZq7VNa7QKjcc0Ee5cvNHtd5N1jgzlPMNvIoZXs6uRp98JlO/0Q8
x/gOx+sPkHlxKIwUi+l7KSMo/BoX+944ntFIqkk6SIoIDLZVoxaqidX3TJxVdzhvky+F25Vi/ROe
rL8Re8NPNRAt8UyIUDg4zUME96QFgfj3x4bQB1OL2zGkaQzdQOUTy8EJvMFvc0l6fJccmbUCnjAp
mEz7PUAwrRvbuR+VQj8pxkCVDwTtMJrDvtDlxMuhCJWH2Sv2A1/j4hLhIElZCT1b/EG1Z5fpIBVI
YOqASpSoJkHkIzm3/WvM90jJz6Ywpr5P//oGfmlpk1R8IIDv8Os7nntewkC/b2qP4L7MNVvilg1p
VZDKdkN0Z+YktbhrFWIR4bihjJ6oM0Cn2sSgL7ypz5dgCEWGmqS//0bfw99h7cv9zi0esZ3jh3co
F5XtjwOSlgdG1Ny2c4DKnWG8cR5z6no93+k7j7DuiL5nQlcK+x/AWyLQvL9K7Ur+eOpFx3rBwlII
bxPAbSCuYG5JCwhbNLG8v8FjFlHniG0AGaAI+sjBvrvlyVCRYnIYogKfbl0BVDoB+pjCq1uBJvmE
xXb2303+p0PDU6yGlQPTYVNEd7T24GA/kqtlgm6t8yiIaDV70ZQJcUE3G2IGtcl45igyNmBkhU+r
IJGM/jzXTnnfnsj7WZsPFmRISZ5QHz1lnZ1kUVK5bk75JmV/gcxwu6N/VwPs6+b/V3fNtD9A6BbZ
mrA36pKSUA3iuL84/zwkutUvmyarP61xrF6kwZKi2F4FXpwDO7jDcg2xcR9hxXFYSbtuQwtx2p5g
sIsSyUq1bX22SsKIxl9wgNJY902UQLLU5zzLr+vVFET5u3gdYrOmDFlxVwQ3F/2ggQZgKUrPPGyn
hzMs2WvpUxyoqHDGBcR598+N2mPCYGDNfj7vwABK9Te9l3CtWuUIzbgkYkDCZ9n7uW7Sk0t0fIcb
nprZsE5MCZWyk1iGNC71RPobL67F+6q6e1A0ou4ew4xJdDp1I5W5uMGTKGcIBpF9BNbeMN5d8aLC
fM9FFAlES5XQU5aTZP0y/5BxhIWo1vOo5eMe/atcaD6rkBHA/ckie/JrvG4JoNX0eBnczX7ZRS0x
xnjUGX76TeqNDe0DhDVTjiD0ZElTbFd1xYapE3Vku8zwvjSBFbxVT5RedXMY7XE4/zNAmGIfK1ot
+iqpCyxLtRXTKwz+zgXAXUljxM5QfNl7yh1cNHgiWeNQxJPWqvvpFV2L7TAjFipmnsjpfM3TwI/h
gxQH2WqN4yxmbkH9P/qX8W1Bj7gv3kWKw59Qp6MXg0mWqPLrgqeta+l31wD2AOpe2VEfiT5Pib9R
jRlPm0j37wjdhDEX8Nj5i2olTPbRVEiUUC8BS5DNBNjTYLW3vzLkgmXFSPU6Ln6e0u6VfCQkXffB
suXK5jmGDmWQDeSVYOzVXuPA1v6dzDVu3eVBEAlF50NJyaOc0zaiaqw52jnnIGV8M5FDopgHp5i8
LfdLnv+3Zk5RQrdFanuaVGdOszR6ye3o6zXXAy3pVBqINjuDHZCBr5+R3zFnT5JcRABhDVPRzFx3
eh/Uhb6dO0W/PIqN2UIkPwpu9Snmnhw5ob62OvMXxbOZSM5aldqEaO6nWTc+/W4YgQwY+9u2p2FR
PoQm7kI1kCqoTGyKLtjfCtj6fEuozqHpRiDoeUaDOGl0/Qa9arDD/LlvoI/1v8t9KoSOSExHLy0q
01+ptUSHgE6/Zb+XBn3Q47PudjyApjrJda2dTcUq3akUjjTkZJ9TyGJZ7OjgW6ybKZwM+AIBnTKi
JUUMI8j/XxRE5kQzB+uMfYqQoiqAAj7YtDQ1G0dyAnPn6fJTlJydu9jkkntOTdfgbEpEN9cjdb3H
fjhpoLcQgNo8LIxJ3OWtHaV54GpmYjl4CH6HCJgMvdA8vrVchMjp0m8sxmF/wKVx4KAJKqVwJQXU
kT0mdeLMkCSbPmZu461edvisLJIBXua4B5Ks+neLQLzB9cCpGLM3sz1qlTJSoe+CXm63l1WntjMe
w/6XO7/+iflzSo8tML5Pkgr2l4zXWaKoQfEWbNO2uBtNqC1fNTiSnQwxrYbdGarCeusp5PKl6v0A
7Unz/9KRdQLrG7ULmVl+Q4fpf8hrybUiSHzO6RPjXzXmcVqW+proBD2pqmFfBqdQUjZSkAJsWAU6
2Mu6jTiSpptb5zVCBhdx1ISUTMnsh0lIwoEWyjEMSj5j2Xeo6SEBscJRpb8jR52C+iU/M2MJvYSU
pMmrVSzsvl3EcfsLFdv0LtxdoE+pYWj8SJJTs+ggpTIQT0ZQrBm4AN5Luy1Vfq3MGfukoEqP2jGy
VsiXyKCd2mrm86/w0Zxncas+yW+wL8wKoGR7o79tP20GPuFn61t+6b6IOxXJ59z9vX0+txoEzRng
v1hw1SUQyEDk27eFwAGPav5FK9nnRKH5dJ5BI/tTVg7Z7VMPStO2N0bweReknCGGhaeBY5vx2NXa
rdL55lnwUXdtwNlaSV9Ka3SS7dzbkLqEdn936OprfyUHSpEChrfC8TDYv98djnYjXTuZl/zJLh3i
+CE+wIRLBrXNUN4bycqpJ82rUu1UV4K2/0MU/xfZG2ce+zGrEmRANLUJ41lHeRjXn1F+qblAKz65
mfpAE2q62nq5TnqVO+76QRTNqhShyQu9WmkMX9ky36YmFQyzWdnqdnqrNlbBm2FrCYnxraS7v3sz
Wjx0QaiC7UOsJof/TP4ssIgvBvJt6odabD+qSOR3jrXjM9Z6cAsmRg+HW3Q6Em85vyf9H8autNN4
sB9wTyCwoZM9SgsbAfxQPO5Fw4OauCnpI7d4YupZQj4trRBw1cmx5vUvQMAfn0iM98hAnfiZRrn9
k7jBGSkgRPK74eXSu41EaSqtbsBlBsPA8RYvsTZo+/VUQDGoYOjguXBUBu+aMc7jNOudEXptHxDI
docJAIidv8rddjbC24z8JXHPG29LGHyFQQWmT3lEDtDjR5lIcVpGJ4xeujyYJoFegzMLqB5uvEmG
/xYwIyx23E7gODgMKkH+shpZj87lRBxndA8WIwMv9AV5bEVUjumGayQlslk8mmdAK7YzsXPRCIib
ZJooUihYD/tmCH1s19LvgP/ImceCRHxAqu9hZV/sk+qnPOTO279JY4u37mw/pXF5MFhxRb/Xz+Cj
DCL8w+zzEk79q2/nC7104f5VOFO0uJT6PMXWUmj8g0O6sYzC4Myz+6lbFZMf+1V09JPcFfUl4j+U
VKGKTIMSc0CB4A1ne6VX+FxWPQRZP4G9sxNKBWmDNUU5X6FMywUvSRldqNxVMd6YIzW9iBrqSNsD
WKr90Fh9hrXh2Dg4HDyUzcX/c38/UCAPvd6td33kiKiMpqX+Oh7p3ietc0gC3GMn18+b4duEiuJ/
QGj3Oi4XcVLLwAR0waWU3+WCoJSJ2t7mFg44msneP9K/zwh7YbVmQHccaJGqFSvpQu0h1EBVf9JK
fFxTWRCxx1yYFuAMnyKMPlDaIruOO8VZH9ST5MXqKPuWhReGBipjKkjk/JQMGW/OOVglg6fASNfF
bOygPHiiaU4KbP6qDRDLJe0Pol24p7xegX0bX72OR9FC/cZMRwD8t9bjaZCHoRfS2rZJ/tS7IDpT
kFDhnZrxbjuSGc/KvrXS4HxAwoLA+rtAwtVPIdGud8y4+NqGIt7sxswZdt0SLYBSViGXg52GAAMB
bb5LPDi/G/aR8MuJtemtkFI5KaIvG43y3AS+8H9T6MsMAi0JWQHHhHaSaqS3Vwh1nmw1cbyVGQgW
Cn4IA/dumIlR5Pvju8UF5w+zOwJdc5d6xX/ZL2vY4I3cwqZniwU0qhnYceXVJrf6pFJfKAP0HmRc
7WCgJC9+lmvrRTLOkv2VdW+W/0a4RH4+iB8CeqSKow67ANHaPEFw9InGGNYHlGdvzBHomDOOp+wi
2kc9jOpf6C0Q7hE8jotSAy1YsNRz5rEdhErFuDzLetIz+1aZV8zHJVnbE67RRjPFED/iR4b65pQA
QIPugSVSJZnDInw+9mmmblQ69OyUW/89vpSbGD6pjRvAyBG1iqwTjUFaXuYX4zuP3uH6V2UqcGya
q5OCPzbMCjWXW6bUdsL0Kv3ZC7rmXITopn3doa7HRpAzyVuirffXY6H0K30RFguroGw+cPj2rgN0
UcY769t6b/T2zwrI8XwEXvOD3rKieY804Sfa7NAGWFApEnO5lRFh3mcLbyzl4u4s4IdNELOk8zTy
zjGDa7jo5agkQSaPi3SHsOkWmlelau/1Z5iiyoUTiJV+XW8gWJjeeDFf+UFDI5WgNoZ6sGq8mD0k
gCs+DH2GG4wbHcCfdVXF60zFV1S6SCMrxe9ATObP9MmNf+YjKLSuN7bxy7mysfZGRRlxDtipgYSZ
HOxBv79GNg/eF90ATjanHo9JttEkSt/gmME991nq7BjP0ertdwW2jenBaHQ/IUZbDPurcLBy4u1E
3OW3HfuCZ8hkIgsNaVuHk0X/PmMc1pqjNU6zCNOx9znG/g+1d4trtVMPDH8zRKa4/9VH2xJPE9ea
/L6KgQjZPf0+zelhCRVqZ5JrFsLFTT0FvyUaX3XZhB3VgS+jilPTEPLaX+kw9I8AyIaVbhesu4AA
6pWqi5v0IVO/uGLTgT0rcCdU8K3lO1wCboCOqM8gS4V8SOm7hIAZzJQ30VvwYxj+ZqGrZwGwks9M
9m83o9CE9iDcLOpu/7GX0OJ92OWMBnmWFfQff3fsAc6tVKbCj10+UXGiLzePu775WG+5DLm7pnYv
hXusUudiY0kOPf3MCR7RR7UVxx76NvfD9DYqe+C7vhyH6Oz9AyoAe8cWeyIo0K98A/FM+po7yf9V
M1GSuddIjiNWhOj+zlfzRqwpd91eJQdAqIFXD2b8HNSbafGo2Zrq2C+BM1sM2vEW/hXoX/HTXoVq
yr4G8kZ1h/PHeWvKQSAikEOOO6yUJhSpnrjthuddiXNEuNAk5+i7waomStLSAIuesBVUDo94bdjH
oP3cbPlinM99ZBSTQuVcBiKcGBnT9nyEXoyViy/FTbcr2tivlT4bPeKLuv/xmoWM0NjDihvutXjg
2q2TcLt5i13mJsfxiZ7b5GnJdwojalwMY76ddZRTr5ICeTpLCgUOXIS0X6NbM95iK2fQzEN2B3et
OQGHPNlmHqa8ZQ+dion+nw4ZoCWF6hGhqb0eMENtV94bpp1lg7gJ/jwsH3w/mePU+bRBU8tcWNAM
f2KcMwpDQ5X/ZZ8WWBstbKQTQSJ1N3St+93T+tuelAvkS9KxjjRLJ0DOK6kwBPER3RUUc+FAagyW
yQFKcxU0pXk851o1EwoHBzdSlypesec2tgZFnaop3/aVYiwGY011u1utCVLihHQiqFZL1ihibpQ5
PACJxMgT0wtEs6iwXWwGsWKy+scgA8ESS9LlD2S2pNGKXzPTVQcZ2UaEJ2yPZo9A+PiV5tRX9DQg
8YxRFQLYpah3wrvAvhdKAZU7KdFDEZATX/pdnq77WB+sUn58flIQO9+r+G/l/ThDuhHdCg+lTX4l
RGHDEwHUtAqDRKARlEmhjaZvjmCgMlV8OH8iKd9J1S4hUt+p2svXInsuYgJmzbex+OeIO93G8BFb
RTq4hKW1vcAI/+0JWrXWtVKVXDArlugJ9vsRh8VTny0VyYYvSQmpWH/0G7C6FwEZLbJrbntmMY+5
WnprPrkVjuqc++yFlVTMedky5N3ofsv9PYJVX2T3QOlfYtm480XhtKTSUFvtc+ArEfFPJ0xU3Kwq
6ag552WKhnHu8HoppIaQckgMRf2b5edC8IwPo/UvL3MRt+tLWQvarW/SrF8QZei84VMNZS0gDjqG
slHwhRLemw5mjKrm1hpS7uq6dCXT9fIKwYyqVmDs0PfWay2znQS/CW74pEX8+reuGDwWJNy1cBsZ
KocxFKN0pfHofiP9qUtkUgOWHsJtrwdfS9qQLpPxaAvWbrP3YSqO4WGK4FdRBkY1oWQiNyztSfOc
9+eZ+BxWMG82/S12HR5WeUtCcopNwc8W8KLNnVhO3Av0T7engQXxrgUEDn1VRvu5UlDVoHkz++xG
A/VKAYTbsR1qUeR4C5hzC2x0MK67+mwbRQhAKL2ZRxf1ncDo+XZvaAKmrJ7QDpJ9g/GgA71ujFf5
5PId/EETpTkCHCp1zJfc4/a6FfnuvjCcjaAcqSgvNT1TmDTX2mbAH3DZpMF3nYlPHV6uTqRneIlk
9GDdu/EP8uNJmaluF0qo8uw/CSUPZDUKF7Jd1qsbSetTcUgr4Of87xFzXKBlFxhcLKxl2SwYsrH5
FvY0D+LQ8J60yEqhGj9N9eQuM84vaMYbv67BQEyfYRG/LxMoTraUwidCQHMfTXdh5DTgZk9/jaBx
QSeABkVEHN2xyykJ+pukeTv8jZAv0Ce7ow204Bfb1LyF1WuGL+kXLGNcrO4huLpxYk+1hYpBVDFf
m1IDSw7KFHOOnFTCBdDhx8Pl8Rco8iYi9I4nS0+eCc0M00xrqbhfv2/sSTaj0Mknzo0VwMnR6eGe
31iOhe6r7y6eLbsLsNr1v50aTCrzbsDMZqahaz/TboLnlulNLhE3nWbDzlshEiGwm6qZ5CJSpQ7q
/MOLRmAmEo4xyc/1w4arUUaJH9+RY1CkuxbWhn8zBKV21PlY6PXYy/KTUSLzyWNwyyleevhwDBoQ
5Z7gagq+Bw7aSOioxHp8OqeSmw7EAKskxGrn3z+jADID9Tuj1zx+EhRrPsLGIEfOpC0jfZ61aJEo
7JbtIFm7CcUG+LCuKdCH9X2Cl3jMHfSluJgbnpY8YdWoHLPGikGmMWxI4r8UvyzCb/PQe4N8lBAZ
bNbWFJCiVJZ0BrgUf1V74+XyN8yvg+slJffLNO/MogK5C2z0E8maOXHQWqmy01/VDN9ESkNjcoso
nr2+0BsBVjw9hKNjMi6pRvu4lYO4viDyZvRbyiFdNmDB99MCntwUjludT3omUEWzo0T0dpfvhdzb
W49KqzCUqOdCDPAFpzZeuPmCGq/ipTZlXnDKVDybKs7qUal8ytxBHO9qYLrQrhVSsHoyl68xzRAc
YWl+3wUsyIdnXCdQ7+MiSsIjMV/NA1KVtW2m6maJ+WKRKng6Yj0FHZ1JjaO7NGN2UY0T8lw8jAMB
iEotR7JERB0k72j2neoSa6gsCTT1cSjrxUeCx1dmhkzCVuKGjUiOgGh4TWwXxLm7HoeyV8fF3ZGS
jiqa31SmqlIdl0cKjg8CMKsr1NO52UG6Zox28+fXJ5z3LDf4wgOJDHkNmFbeirV9C6UG9dUz2WP8
iLzt/rMa4CZ4AgQ1o6Bf2tnta2CGkMiCykq8OIVsbWLkFkyZFM8067j22Vi7SFiIzhPtFNT+p6G1
kfJ6bwDuNi19kq+HZil04PaF6FJfItGYeAUip9Qy0AB4YdGlT7nY3F+MRvRwh6kjK3/OQdBgBwxS
S2tkzk/K25l5NuR42VoJl5ofspMIk5Ck5s12tnqQMrMRA3cinRzX5CcaBKcQE6mgipi97E7MqAdv
P9/vJw4KgjzvR60Zz01MN5RjSDigiXkLHoM/ADvqy0WcIbmKsa5Pei1S712aO1fZ4GEQfHBKLa92
+xkbzELQusRP/UsexgKI99woLf7LuoOQiiI9YVA3CXYzWqXBM4/gQpUq/9JIBS7SGpYg4tlHwgaX
YpfvYyQoeBmO6CMgnCjux0A7+jvWOkixyDOVAA8Od2dGJG4Fm1YqvKp3ZaLWn/dXSQg67v1rdByQ
iR+kjryzLX6QicRJGK5urBKX4cyE+R6HnE0mcJOdUjQ1J5Cel4HEDcfwSJNdJg8C8qJ1fGFf4lZX
55edDHTGbpwX9rxoLUEub7jA1fDEVZLAooyekp+qhN3JxmLNyq4DOUw//DZCYaPtocIv7RPbTg9U
+HljMrpY5+TGWECZoQOupmw9Oy3hAA54euXhmL0QB28brOkqTvHkHAB1oFw2AwQoPSnM4wNsnHOX
tv3ZlKVbrlRWpVPcgGErBGULdGL7oQNb7wA8lKFTo+h9umNrGUSYe2578pg9nPtbxBzROrEAhAj4
s4hW8A69B49UZbgAQviP1Q/BZ0agwbknVrgeXApe+F78hnjtq0ieRS92OaeEumSfU7612Me7ixoh
d7jLjv2YtAwpOV2Ux/aqby8/o3Jkql7MQCBy79FCLTNDtQuxisNvCvlLxunJ0uMrldhC4lVRhuoi
MAXmgDGfPtqwDb2E7g6mE6HJDGzpL8lC6BxKy/UI7Ot/cgmorkaKDPZOluHJQpqDSW2uH82rHnCO
N+6xFchtG016SFs7VbrbuTlj1f5TJxyyP/Ey/TQci4Y4AYl8qVfyazFCzOobqTePnvilmwqgGuTr
5ctrLxL1GnJJhRN4Vnlt4zIGKqx4qP8BhTv49MvqUP1j8vW3+/Ljq8ekX/5o/fojBlJeOL5Sa4ir
FyiHwssdacNT8Ba1YdxdSJg1LiFmF7ygt7uh2FOMWpYXVJu2nBRrXRB/q1I4mGdhcwctaJLOFNLu
LqeaxNyiD3EgTiqPsPIQCzQBQLnKQQgu37ossGZpTQmIZpxJbGUbg4HyxH41p42wwXBD3SPWM3x6
SZ6P4oUfQv5DwMDq6PhHT28IQy5saaC5UQXu5F/94KTHYOl61/LLseUAaB6NhfUcrhaijSVc0Q+n
uB5cpYd8BcQPsBd5QjW7JRxLPX1olgVKdByuzBMPYHUXq0k/2gjEhlKSx/tUN5sn/vn7rkPxO/tm
I2gm10jqEIxdAigSxKOyt/QQKILkng8d+PTkeQ5gKAhPu0SYotpnf9oPv/uAXm+UbCiTyzhy3U+M
Sx+2ioBsQmg0UKZ3KcStwYSYzvWMijlqEBtysUYO+dieoVqYtkGdxC33b28CqYACWyfDE2kWHDQy
rZImzA+VikowgwQsFar7Ou7unRzrIOBauYjpphBOrMSwVtTzRn+977tdMhHzsFbQIEXP5cYlyCRT
+NmiSaoB+gMu79tOFiY/GRPEdrIHdccMGwsEZ0k0LKH+nAUJoOj5tAvGEN1nbZg8ovJtfs5oMOlJ
y3PLTSZ/aMs+1CaNWl9G40gQ9I04bZX2CarhmP/sYuMpf1d18loX3xMa6XSC5KPPsJEAz8fhFFs2
kiWvlemjThnGs4z7ybv3G/6g7TmBwknvH3dFOA2MrxDbHsfJaBLhX/m8173bRh1wtqSPQGNUoWEs
K46r2xD4nXz7wX9BadVLkgz1Z/A9/FHZ2YBBabb5/Ia9EvDZYH8MgCemebbrEsFwHrtSD4rfiefT
54JU2/mdLsph6zc/a5ShXuTqPnVQswPvQGgewaT91qqsOw8dc6xXzfkt0N8hMGjHCzPL0DAQH/00
D7Xtw3OsdlwzGc80CRscOzO2juJZ+vz+pM7B3ULIhpTqGtxqHXWNmsMc9+BtiTlqrw21y4k5Ea7d
1APPB4ljOfPgW3LVfrlfjUgE9FmZROyNUySFsZQ1f/mHdghM/Bs31bijyFis9JWwe8pNgowCfPMa
lbGDmtzqKIsOqUGTPBg5wzXtOKo1hOVPy1AbRAc68YQZmGklwX4xoSMUaivDd737jJKwNFBK9bfT
iBlkDc/dOJ4gzKPtFV4FYNxmmaxYmmoPVYkxAs1EvxtAHt0t32Ax1yN0AyDYqPWYRWWH2QxtxOUY
eCTJt7PgrC29tIbcX2m6hzEoalQHVU0UXzv1MvFH1Wk2pxP4RiYLyOLozEOxX+G/XbxeeIuudv64
ncf2A7R282SeGJ/enVIz5wZbAYThY5Fv2tkxlE4aCA6Yvm/eB4Nsy0S55JwKsuiOC1MgnponJSS1
K60BYrflldhmDzqEU7ZClS5ktlxpOdVxtGC/9yhNsInyUlm4dZ53NGWFa8U2jSPiflm23TpONKKm
l6sejh4BZr1ib5GAW7SpDTuMEjNvVGnBX7t8GG++X8oZI8G7j616yPJloIFpbDFzy8hWmltSh8vN
Muk1dH7xKminpDQGYdRiio+2j20qsd/Sdi7JgtWA918fS0/OFeLOBVjEph9FIIGaGBEcJ3GVOUyd
BuMJBm9JP20hJG7SmyqoMe17/RkUr44kyxdQr0sIk8GCe05fHqcQkftj1APZV0JnuyMFla9lPwQg
vQsgQ2/pSxMy2ado5c2wTDJrCVnlFDIwmJgEEkUp3bMxuakic8ko0NDX7y49jBC+NYhk2gjPLVoi
Exz9qxxXKafY/Stv8J/t0PfrGu7URCLJUgPnZGfXV6ASEcrqL9x7bwJaKC3LndrJxPuT4+PzNYjN
qYWQKbKABFCRDZc66iXdbVdAminoj06JubSfuTbboR4SMj87wX2672E4xWcYEzAgJmJdttrlxF40
1QYhmzDVkJz+RDSx0gGjTqW91IPShn9krdlLjXKSYDsbDNtDPRIkzM4JzI69mZi5AY8++ZDYVTGp
hH8f+UD13h4+DD5IWyLrMUvzRY1+UBoOiuRiwPcoalPACQ24A23LJpDzjKdFWen33G0Gl6/OhxuK
aoT842d3UxnyVQ6tTz02vBTvIFmgDOIA+ROIP9arwEjcMNkYIMBy5OaSYgExmZenXmwKsE5+SPtP
uUq8oJzv93ozetghRtlFO4AWbawUWfKoKPWGsMePudf1TW84Ie4ec4Q5+TigV1liroGEq4vy/JTn
EdJQ0k5CG1exFpzM/KVTJhlVqT6elr/4964e6yjsmtOYS5OkwNCqLdY4n+3wUNLu5M2FsSQFiHAY
45xSou3gb+0sMijVNK0Kq8KrlqkkgdxTMKu0v/Wh9gMI1LIvoIINTMnn9WpvXUYGPAOlnPfTIDZO
eIdlqb4acZ2lkPfUoMdrK0yu2+WxU165pIzkjs+Ok8foWHrmMXIuvGHy2fJDIX3RvBrkSxOmdaAh
o1486oBUoLIfjjH3YyiOwA+q87A3W/2Q3aquihtDPjuTKG02nAgTY9kb5UQeXjnqO2OBYKqqPN4B
RZIKgeLF9dARNNrsMb156Lwtc5LqtGB60lRIQiA17wUH0kzIfMdgvzdsX5e1grAXlZYVLoEsZ4Uz
+YYOX8LUWC/b+yB34uHtQEoLP/bIiGcTseL7y4L8rx2/ryDYDJ+HxDWFZ65OX9aRHjvHEn7gxZjG
2fRg8IW3pvihtGBX3x0xk3JtPemMj2SiKNCOTx3Jq4o/Q64LARO8kHQJc1movxjAu/0zQFMdn5In
Ck0i7IgA2G7E6IzKeweA5h2PONXgzW1Q01Rev7YS/DZez98Dd09s11OfojaozvyMEDzv1jBfSe0e
im0Rot1JEfF7vOZ01t/rH6hTGLies76i4Ezj16r0KOeG+9KwsMPfAa9AlMY1Q6Yuv15SkSIi7vgH
88NXXsJGmzLByg7Qs1xWaMI6wG6/IAYbAjJR0BnuPGSwwi2jdhKUw4yoU+0tuCHtigeHyCSE5fJ5
zSsG5yDiLEjeB6dKV6uYB2vRIXjm8NCBA6mtvEhQDmGtnkqPFf0Td/YTEaGFbV2O3JB7M4CRdKH6
WC6L0lh0jm03pmmdSn09vZ0aI19Aw2zH+6Vbc6QDY5DlZbPCqbLXQCPXE5I41T2KQdWOz687u1HU
fnYr9ZiKL6E6hZKYcx+3xcz3G/JdnmnW+boRPX1ONLIDzb2z5NMLEqMMgAFfqnmCc+x7IX8Aa9Hl
oTxz2/plDwsuUIKboXC2zK+GECFoIc1YF1Y010I+Xvf8WszA7hzALQIWA8/J6JE0Y47JSOB9tsJ+
/p185f6Vd1k6/u4Qs26S0FWiGJNOb2oQiSo2737iys/F/U4dACg9pz0dM1dA7EScql1DZHq6HL+r
VMKyToK7MVnU1NPgz2WITCh0S3KhcQcMvrtYwUEXIsVkydZc/b2CKAc6IWiYu11211k6o7XRiyAI
khkV5vCBdG6k424Ji5KqP3DwxONAjvI6FO+bwUerMrc71R/utk4+V2WjbvztAZQLO4lF6EZdXwqq
JR9ygYqRGY0CAU4nlEF/EluELd93hFEkMq00OQv/byMrWhFMeCJzGBu2+VsVOT4eGcuXxpx01++F
lPx5xXRKKRTr6lbDp2DDmY4tirfrCRavzfInAgW4TmevsDkP0PwS1cv7w0bUp4TAYTke9SXQAcsz
25WyF49oSfTx/AVBnpkJLxplP4iAAhbXRhC6BeodaJhqbgu7zR5FkDTHZj5IIB1FS/U/ovdsBfD1
ulQiMFxWoVTFhL5f8ewR+xSLDesrUjJYxKQQuOLbFH7bjll6y6DY9XZU5VRVqTF6m/adjfkPVdmm
14e4V45PNR1OCDEDHkjRaus30jNaa4bPh+6eBsq9p4dhBo8Y0vPfGSaDJ8OBwcLa7othT7R+VNXo
0p9Ql2IYjctJkIZHa/UqZa183LZjxaIMXE/AQOWnj5EtoxumlMUk4JIodm3x4mPNFTl2SaJjONPu
O7RlWrWveM+xpNSHCFWnxRwjZlcnSmZPS5giDmp3Hcaef3gXibagDppvrFvTXWEo/ANV/5vs/675
aktFjtFvx6fx6rDsPf/8SZxH//8qcyUumbIMiKPWQnBbWyBaVIxwg1hy8147UDjbdNFy5KIgF5gW
ohs/PxjkU//mixsiJuWCYhUpNu2jrZRdoo90kTovveZ5B5qaAXqAil3n+O/nBkwPzdAeIS14wdGA
gr9aGm/4UJNCc6jmCh+nu8G9c+Wa72HB50euHuDkLI3eTGX/cXMGPHmD8/bIWT53CP/wrsow8sEP
KOPPy+3gzXfwl2VMlS34fYenRyGjA4nMkj1BCKNPFIRmZPgGa2dsgRoOthqjK202l8ygk4JFESa9
YgLOtrTM6xgD3UGUJoZp4lwyzo+K7RgzlNrpNl9HF2WvB4Wwo911iV2+/A0zRjGSFEkR/WQASmSD
7PTRFSUpMAdJzWEJDKXLbUDJ6Mza+2H70FKA4uYujY5mQq81G4xcjoV83CxtLOfAzB2tujFEC3BE
o5EjYmNxiEVE6x1I3Z0Jr0ESWVqr8aJxDw4cxrWjNP+y6qggvPzT+55G1RkavaXK0lkEKMhQkxYM
1qg2ZTTOI1mxqAzhoZO/+eqiKn+mziyNB+Fct8ORP/q3DA88OM382V4ibm2WC31fQm7qZRYNK5Nm
v2v88Xq2Aq/ZfliHxVtwOHBW19rYpSQbJdpMlj+lruETKc2odsAA0bgWDQeiEFBfvuxGyAag6iFl
9LlBo8JSB4CcK+1j/uVRh1qV2adNuNzeAoIHAo7s5q8rkzeGqYRupPd9m5hzhBZecYdMJ5f0vb8g
smmlztqOzwAF7vm+2CCQ8LY2ZLX+LmK9pQItkPkEzEOMR7OjljYu/uD9St/s5jQUocbiZMm6R4cR
mjRqfPwCcNnL7P+M7GGXrU8i2JUi0miJ/BFj655RUMB6aQae82gNz8Lv39NXZUkmhOO1+pJT/Ifw
ofKoLogfXfkolysO9ms3EwgJ2DzY8YJCnJlZG6RSisTp+0d+tyCmfNs7Ds9Hq7+nV3m7qhpAd+1r
9v8XB/rLaX1GvqyoCxPME0uGmCrWrfOQkVAPKw5M3rMzRJ+1SG9AztR9v9+qjsv3VtBatNJKbEXk
M0H8s6inNL0gTw5LHQkbuZhcXPk+FhgYfSvEEQmmNEvLV8Wwl7Yfh4yWcXZPyAQkZQQacPBNfF7D
RoBlbEGAwBcHeK8sKmuJ1Le85lHlmLdbEWwWxE8VjFaOT+PRlGYN98TmY0QTMNQsHew/pfGbVfVh
exnVtVqwQrNut4iZianNOh36dB+qXJBxl88hAJvnmBX6EocswPyLgyjzNT0J/YGJIa1dBiLDV5Ne
okSe8odBQjK57rB54OyJquTOWXwK6h2KXxRLEtKoJW2nnjO3cgl4DvXpNIELwdZDVA8UcGajq1Tu
B11YR64TXDBt2uFWXFD0yVz/T7dOXyLEpqOvsNFkx14AHCD0OG7MxDE6YxGUPbM2Wezvf22hhv40
CtLv11pr4HqiSfjY7PZOjGS5TDqzS75J+08fk3kjBz6l+2tria/bo+Evw13JJLjMT7eF1atjHEEd
HssqR8sWQdOk1U9UmZSoL5OG4QyGHw7Z7d9Zshfw1VXZ87OIdcIXRz2m3q6sggE2jc3Bbq3YMu1k
jlxNpCnyQHecSY6dINYFtqmHnTSGtuX0ABNVziFLLM/EfWn/fHp6sokTwm0K8nBH+9Uxnj5EVYEg
7Em+PGbw2mYOoOSAKrrHfVbzuxvhIs43qocqmWwiNbi/nM38fy0+YlYLtVkz5410iaFJb/bH0UYp
4du0dhznhL+XjUVUUGaa3JVqmqAYvio9iWNo64DIu/NppHhkuuSFDBQeiywUtOaa3Mo46qvFajYM
4iWI6b4a5dqayF8vngIo/0Q4ZdfvnCXeaUuMHYxP3vFApqxXPoeKodvsDV7gASzAX+MSi5rmP3tw
JPiafzvb1Pr8ugTnXlbwyaJ0hdVzL2sxYxEXEF1tD+O+wg81qfOp3FE0NzFzDqkXlNZt9+NRh0BC
kAXp+r7w6V/FwnuJJrxISC1CU8mbj1hYMhmSYpmiz7dpFJr5pN2waVMNb5KWNzF1CkNUsrRsdJns
kFm+HCjZQMbSAOvaYBtRFlTXw0xTjMigo788q0kQkVBb4NJzVaQdJqKThpmDGYIFXxfaFIQPk+eg
CsSuhu7XGnx4FgXTQ2gIY06RylRviC9vhcM6rih5DtI8qk4F5ZC74nii4SNJIRyPaz8jQIuhftno
CM0ArdTkjYKyy+Gx9fjjvp8Z6W39mDqPGIom9ScnjJ6aNbp1/P5bfHwlCFklgtY0FVHE186RQ34K
1miLCa3/NLTA9QpmKZsurxyE7qCm1Seb3I5TrZss0o4TLivALXrSUvdpCSftNnMyTEma9hSYaqMb
DISIE8I1jAoq9c3PXrjQNfqpeP0i+EX4njaTCfieMhSwaJl32B0v+BmDnyKSViJxokDK/roRzo2Y
VOfAikgZQNkz09CQmbG9xpPlr9StEeH7MHtyoSijgNJsD8Y0Lvl9/Z5RWHaf/7zk4XYMS4b054z7
5zNXWILIMDaa44sS5FtZ32N7h4n6Q94UKTnuGdt023iPUwD3OzS9aU0S23MfmzwTkmMPCALLGMBt
vYxPkCQQ8hgVfsv8ybJeNCfXY6mql08+rirUFpULmIF/75EfIn8iZv1KYneVH776kaCFnYs2Sqei
Xi8YNMZ21su/x7r9oXdPlClRd21o2uvrL3TeU1RSA3UPw9hJ9kgn3kH717k9qtX/gtcnMe+o3w5Y
bwCUefY4eyM4IBB8vxdnJDoNVVION//8xuvppP/zCFdjqtvobxtxaH9cShecpodHJQ9Xj5N9eWks
pnK71fTdsLs/GJbGVhO9j+vpEQ0y6sAXSxjbkJMMTHCXu8+V3eJBn0JEzDwuDjEE20XlridA7/nd
2mo9yrSx8oBkMJm96Fuo09Luq0R1aXkXNhcKaUhprePj/NKkNag5++lkxyheP7aQHbzMS9JVtL5a
Ddlhq5AW10q1VctZbPc7YNEILKCn1l7Oer62o3/9rRjQI9+ZgOuPrptj731P9VkcysLp6du1OeuJ
0G1wPtCh7nEin986u+Nka7T2PA4mWQlgQeQXyNREBCGx+ECCINEva58eEksGnwXcsf9xFPisXpaE
Luwn0ZF1lE7SGzvsVuDcAUGV/pFC7yKzxd/LDTQChc5lIdclhgGHzkIC5DtnakuxWRBqskDG4cdD
i60XA/dEHHCUc30ADtY5BbE+uoOw0XQOqJzF8ZEk2YlWvmAxs6YK7CW86hADlhN7gPDGzHdYhjW5
7UecnreH3Y58a8w5D2HWmU7y5OIxVZm/QlfUvjIqK9SbDRr0qG+2HXaZOuNoCZlNq1SH/eOweH2E
K8g8haqSckkkeiV4jNa1mcary+VIt7aU17WeqeMPJLFlNnx5vWbUf4p2vP/Gyn/Zp2BKFEF4Ux4I
NZd1CxXJdgqEXEn6XWm65Kjp4PyO7vUYNfo9Kdhb6K5Hngy/N6Rr9lk/RdT9wqtIs9CkBZjjrYuO
LfMWEH6/Lj1J59d9Snb7QbyPQso42pJW1CIYvOWYgLp5esE58YQoO1IdzPH1PeYqfjRcPZ3/finv
QJk5uQOAKiqiQ90032jvYZxB5lqvpNjG3liScHwcr5PPCvXrtEQyv60iucbrJP9XuMmG5UcBhQSX
ByivmzH+pSuIHC5mrbvCeN5WHorfnkyZyyfB4XSvXWsfdNSaSTgPgTCtDvtDPTIBd2vd+SP0lyRS
YfQusaD9qHC0ztXCBK0XuM41XB+nT0BYnwkJcKl013mG/UTIngU5udq5VN4/TfTg6RWqTMez9Ont
F3xgW1SwkWuDZFWFGYlISvBdsAuSpAqI4g6iuGGQBroRNZ6KiTaDzwXIf3igo0iPuxycnltVmoEL
rNNRgcmr5L79+B6RgXPt1iNt3ubzgW9YKG0uoB0K8trMuZA2M5ioafhP7MmbiqKGns2yHEWeLSTK
vb2hr/Wd0QQCJ6tgwiHRg/zXYs8YAoO8lHnZyTWmn7iMrO7fRz9ZK9LLPei/zJTKgKkygh/icE3H
IUVr2OBMNirg9FgXQSp1i4pPGXmMWol1ggAtvaWfRIQSDtKTadAi6XNylXUw2wldGDVdncRl7Y4W
H06hOHjZEN6H/zOvZdEADbaIvWuFRXdx/UMnCUoRB9qry2jYS3qMXmytLVRawW1g/TZq0wS+2mQt
GDayi9S2gHfj3km1ep1/yqLq5Jys+YuqQvgjZBpkl4VGceXCG3smyBDzgXC3hTLLlDd5ZPPZHnfy
G+1mRcKNyJl/r8msaMIZTnZe+wUBXujYUJz8WDAtsLco4f4+1yQs3LkgeQGIdcO3vZysqYtP3tHy
ECNIz8kLAclcs5ejF8RKpt2ky0l8vJzBNDt2K9tj7PBVNvMByUpEOo2vqT7f8juNGuNoXIT9icjr
J32tgYGfP/Kt40T0HVGruGK+PTw3Pb/LV1r9XHHLFskBL1Zt1arHQtCXQO56H5mg14YKHyD86jSs
ocaDSajJBM3+SYWsPvlmfAYlGwqO/lYFUkxAsyUtX1qtdjMcXk1vYO2ATwRsswHb6nAzVNJu7CXt
4tdjT8JesxHEYiQwnRp/r4f2Ohm4lqXWOp6NaNJQarHYOP97gCOefahDw3b4hy9IUd7gIOTLwZ+1
T3qR837N1BlT4MptqhjBmiuftPRRVXCpsIDH6BY7qKPcaHYbkIf/0IzpsFciyv08/eDSvoFThcdJ
tViwZUX0ysoit+0nE0p1mJEAO6F5y4rNrtoha/LzP0fXgisOa2ZYOTe36MVZpu0A/8arLzCYJQM0
BPkAcJRoy2Fp3UJdlEWpciIBxA0HRiMVA0uIZIUbXVHGrDRzgHVQAVgtfXlgb0IK0Ny4kGmZinHO
xV63FSEkLRzYlMpkL5eNNXrV4Henma+4EgjmoOubFYY4+DpTs+O29aKWWcgKYNx7/wgy4507nkR/
u6vNzFiMCnMR51DZv6M1oyAjIk+jfblBcJlvVVbIC4CvLpre/6wvZdOkkzx5viowsRojWvYcTvRI
a5AAEWSouC9DRzOpNXaXWuhFL3fWsVfGAEFYU9+x/ya4Bo+m1ihp+/5aUoS+tEQlHCxoWSFDk33X
fMComuobuLenzdKPQml11/uueKYd9AIMrzQPoEjmowkjwkjGY+MyfVfqUuCVxVwDOCp3fWzuF0Ce
ez0saRE+VZZFdzHibujV3n5ozutJ+khvpnMyLzd+TG+Z58Z0cLTNLLWFlaOj+JUBz5b+Iwhk9b/z
R+ZMBIIn4/190UbY+kYJrahmeZV6Id6rb9VLJG9nsocAkCxe0eDobt2lXTLwbsxwewVcaCEAMKy4
b3bx0pZX2PAjhCjI4eOValmuINc1uEao55qseAIVDdqIaluaG93buYpC/UGVVPbIBu68fxCEPDRJ
BvBkR/WEj2bvKm/NkP+LAzjnP5mcjfJLVwkmeMYuwqfscnsB9zFMHTBRSag+ZYNncV2ugYBJP44c
Fsp9WrB77vXkcqgp9Ri1vZurP2BM6F0QOzQU78PkKhWsyoaXkB269SJtsrws5fGSVgICioSCymd6
MszXlt/ZGKLlPeFvr8E1nOKTrEMiRs80n9fbxUYoDui+XtTOnp0UPZebfXeWb4cs9YvwzTX2uu5k
L59QK2oneH9LppvHukJ0QiIjnsUTYJhktV9blgz95+Pqgbta4hKr3C2Wv9pEYd39nzjJID5FQ396
2n0B17c9Wnj5Dw1Qw4SDFGUKUxLYaarwbVRX2SwyQoeyZyKTDMTZNSqrNVDcqYen0VPKjiH/3A3/
uAtDCqoZsJUHJAOt/vxy6QvEVS8CK9Rg1RK7bGFT/gXqyZ11vfFeSyNIBNxUMyk9uEi26/ueKISE
X21P+piiWsBEsk5ODYYbp8SnBsgP1754F9v2TqSNDm6rt2spMDy8Ed8x61OOkOvVM7gloYalhqeS
jyieEghCoGiIOEu22UK1SLNdn/bULU/YvYb3w5mb/maQ1sueBiCUawbH7PD3To+WFl6dh1p4JH4d
R6tSjNak4XPgnRwgdSVMlyRVfEKE7a6DMXnYI2F/PvzfyGXvru+HT8cwQIr/JbV/a6batDvmzlBe
s5crpn2cfks2gEsJO/U39VmvLWYNSMTRscSBeGUemaBE9R6cmhUvALAPj0w6g3d5F+xmQbvlJuE9
eMspYoFq6gCEbVwgUJYyKuI3W73a5G3bIwL5Gu3EKWhxGu4oRNSzAg37WTwoeEjWlafpQrnLodSz
dotQweE+zc0pjJMKRMg0hqJE2KVVrC6mHK40ltBJOrgnvs3ERq67f02glT1D2qPANdCMHC7xvUjV
31Mk3PGsvRVzxotDQrJPx/Zc9XVZVo6v1E6UDU7Z+ctkv6686IX1+AVA6vJ67QnliloXAH7hZOrt
I1j5XSUBcMmiFhmwexraxGhQeXsmq06RUTmQ3s5jogiaCVCwMlbYFS93kmwkU+z7kExA/w+Qxdg2
3wymR6KhJ4i9++77Q5wgMlJtRsrfyH9gYcXFrn/RxwLeZXaBENXfv6EXtZDdFzD78+nDLEAJLXD3
mgZpKu/OKlVH/2C7eKlYDO4IodA192Q58QnO5/DzrkSEiutRMhxhLDdN0qhPYggTDRZqgvWwKgVq
cFkj4UJtWXLkMEpPdBNiZ6OTHotOMGk1ww6SkVVL3Ie5t4Rzs3fb+rIuUYl6sBk2Tf77O4NjqVps
MNqwMagGl9xRwMlXD5qZ4szEAPYTdOtGxgA6ffzjhIfFVppbnp9ccr9vGzgq1BOzNrF8bq9P2X8O
RUjtH+xCHDq1764+WhTPiUTT+hYn/Akmv1wEENty6G2NQrzoNLTblUX1J6jMNxsLkI9pHHs+3S8B
+2X0ymTPwkxQ+wasp+JrngHeKKjTYf8FO2/wxCgk383VbsfOTUmC2VXsh7cEWkovvbdeEl9KRNXu
7eArIzUVnMtXROjjBtFmZqcs4CenxNeOoZc4/9qc/95WGj51hEH0auTjeq+3/g79IchEqE/gjYlW
H4NPjKDonGr1BrW84DSxGvyYRSBSuMzMc+YKrq2z1Aq4fv1NQX9qSsg57iBAIsd8TmnzaUHiLsCm
pwXGUpj8p1vMS9CfsIq7DqSVjV9RiXJrCt8Fu8Df0l+apoU2/cuPq/U7RApv5APnf2cbuyOzncBg
9S0uYHseNLxmr5ckTmkwfhItpGF/movafRFjAs6z9+MtZkmu9u9hbouurUnnogcfBc0E9pRKtXiZ
I6SOzyHILo5poisFkaQ7xi3F4EGMEI+SJuBT069jsn9O/XFQrNY5tLuGPYLedDC89DxVSp7QsjMb
upYYcFUasFYdt/4G4Tmr8Wvu+HxU5cu5aAqHfchnp9J7xoZmAnceAcZscsddZXDCCoVX8aM3daj9
YXiTOXyNEGtP84HDlg6ZlIbkECUZVls40rxjgAxQfkXxPwCyq9UZxfTJpRVS6VySAzPWUKvUh/Ot
xx0YsYTy3WM2NuIz+oNHkyEtg3lyVBnJw2TyWO/p7Oi6kxLbh2Lug+0wfQN8cr+kh3jT1pn1ltPo
Sp5D/1AjZhwNRHEPTjbquvfhLtpVrEHgIRyKOrjnZN9yh3vmOHbHqPxid9dDugchLjgTBolaxxBO
q1HBIe/9qBWCXM/VhfnxnbzTcO3VHqSKUvc7Tk1oJ5wOdXj9+Rz7qfuAunMuFUVd2oSZMyeqTgRC
+mZQOYkFMQpnysDGVMzUsTswNduCLBS4AcOr1L4gkB5moidRdozdf9ax7DWTBO+fKwH96gkZj955
VWzv+bqJyeN+34E5GitcxUGkLRSys4+fPb5kQqxxjhXXhcRmwnDH9Q55CVYzePr8b59pSWHyVGyA
grWDNyhgNMPDAWCbjR6lb2xtZTg8xMATWJgYQQ7Fibx+oosn43iFInQx6BEzPbpf6xYl9FOdxCbP
+z+1DLNaOZSkA8QSqURcMVP+j676/jtPu38jrGCRmZy+q4S0ydDOjAbjwA7G8w0v96LZ+/sVcb/O
t4RyDjdmDuVpMlM0nf0sio3Yvl3iM02nFJUTOBUx02d5kgqsbO5G3xG+R0DNSGejmoCEhDxkHQWf
HNUYfz0Knw4hBbIohNhXm9kbv22MlIx6rjY+g/a5n3FWp7Rur6uqL6+yVTWXjhQdEsAzrl+d6U8o
SVcJ5R2uhbF4kwR4Aff1Fu1FOzK8a2MEd5rqmmqbfKvsjYLIJWWEEe3NN8yDDAgIq5+6Ud1sZ1t6
frdHSrpTHtCJ4lzdhSPrbDE6EBoT8wL9zhs8tzIl0N7VI8LggidKCkvn5kE3v0fkwqyTsaLo/98h
HTv9zrl+zMlbCVlIJ7T2bmHUaMRD72VSxn6/vz6aRNv8QVzL1w7/lsk/zKM+UlCK51qQDuU0PnMh
rjsNX7RO0bTUWNKHLZyF9QgBU23yHNFrwCL+gBCGDb3iREXXYZiSiAW1/OvDnMS/UjVdX5W9xyNc
1FpJy6i6Alsxu8mjbV+cR6hYdTCT9OeLA/DxAIID0pfGdOx21Z/S1CgAwTHJHLEoDHMwEhqZVGxD
Saivz/h04/Cu9ll3jmRj25zJ/ABITu1jHXjevWCgYLDqnGuVmyj+E/Q6FJRA6iLSeFm78oKDGe3D
Jv007OUhaAd919idwsGX22dHZ5P9uPvAOh7Wk3mp/nUlg14K/T+GNS3zTimafnEENw4QqWoH93vc
TcfNySYzmC5iuRJNOx8UizIWUHhZ9rJAQTxOQg642HwoxWINCsGZbSN/fmdqCsmHYlL5rEVvwCtZ
PQPhDa/jaQtTlrvYM8J2fHsjykb9rRxMRytTp29H85v+Gpk2uHNv+CgsUS/7ZQfJGwl4x0Vj/pYp
Jqyt2T0HsdzZh4O4BHXUSBA366E9xJlvM2AXaJpWGLzpx2z009+W46Q+nUZKCqo5ZsHVEztSJ+wT
XURmQxpOIlatWFK+q0IDgMVgnt5i6bGHYHnmJc1Rr5iAwZ/vBDZH5v9CvL1p0X5gZwdv2WlzaUPE
gmtBCNTUrr+Or5wnoE93f3lK+uQLb0wL3zXg/C4wusdTbfo49w48qyycMlsL/qyqEZH86PhjjeOx
VGKwCvRe7NyNkKGLMO1kuupPu9UEMUfAK6lmSGTs5/32BXzPlLU6fR8akzK4o8YGiroH4g65JNXC
Yj5Z9CmkcxXLvEI7dQsmNuPoZ4r9ncWmYDYfSU/2f17Km1ilYyEuDN57i75ru2spQhGjeTO9R3z7
+eeZMBaJ9nyVQ2eO/r4wYahnrgK7OAKgUKmogWlbHpk+hSFVMmtwuOcJ8RHFsu6en+MVm4Ztk0U1
Wzc81PFy4DP/JWgxlOijwsCYA9DQvP55pQ0jZw19VE/t8QMXqZBfSl6t0qbrsCl+7/1DPJpKej8R
5hbTfyQgvnUKkXtLLyX6rkMuE3axF6P43QwLurSqxQKHLGBhufmetKOBYSQXa8ivG2zMx1WygiqN
gj6KjQciJuJ+cDo1qD35LstrEBuxnkjWGAhsupbOR/KrVntNspPR4RS75bLy6H/rYGhJusOvbMEW
YohVF6Exiajp1Kh3MFf8aSt1h9Uk771s2zjclsKoFKON4L4dU685xjeYk9RaiyQyoKue3on1l6nB
LiNbhimWCd0X5Qy1gGVZnfhQ8INma3qM0cvKEhe8xZPnYuXHCwy51uPh5w01W9ojPPyEYTSSHNC2
iBpERO3KF23vXQyzLUcWDdIIVDBijEpQMba7jMiEJz1SLFipEmFKcmcThZyBGRUM7BWAQnCAHMnl
AbiAyunJux3LlNx9BzKsXv7O7a4fDu3ypHTgFGkU/qx4o406kcZihXnHsj28w9oJXKZJa6GNSUm4
jEsLhiMgYDWc8CRpsx4zdIWBzJQ1NcK2nRnQJcuT8Uv2Dv8GkfKyfh40m/iuMLmYWei264rTiekW
yExjoWDbtxXn9a0cmvdIxuY9ShUxKQA8b6XHMKGBrMJ+naWYyAo5XTrCZkCt7RLfQn3Jr0+ImZeO
1hEVPBuGjTkyyIpT4h/waZeFtl9z/1p/XcsJcGRFWLIBN5L61zKsBVDa0pfpsB1QLLt8pW8sYt+z
jUyFGdcZxYw0cPJ2P+XNkc2UvGxjPuZeP9GKkIIz1Ns2MCIX/fZqujifUaSgftJnZ871Uu3RW49/
/eVrZJ4xXPdd5AVubFAYz7GGu39KWmiAKjSRf+Tt4FbWXwKN3X+gM86GQpwT6HibO83iO9Rnrr9+
tY/LaKWH+1UmldrJMXBOfkDQZ4ZHhdvZBReMRqp/MFu1JS/myQFiTMcupCo0uJMkC+Eh6X4Ac1zO
Vg5gunJNG8H0+pIhREoSbAYlptBKZ64xKhkP8sxhk3aTX1G2g5JIkwJLQsQpf2L3OWODREe9+fmo
Wpsy+cB7n0X0a5BaBShRxLRyhUW1OlhBAJMwzdPPfFeO4ay5pJdw0Bn9pmoRx73tjHwK2JnWXe4/
/d3gaGVKRv5RuW9uVwZMtuQ7BJDwtBmgBd/kCaRkKJphCzmFRnKdGfcKfCNkYx2Kf5ci1womv+v6
6RJ+EFsR74fwpCs668b8wpTLmZGDNf+4TWD9tzq92/2pNtpMpwVV/Hu9REhgH1TfwUso/7fyYr6w
eLcdLOEmi73y1g73XUvmXefr9U10zEtJrvsMpQbomCqUuLf2G1fxfbvSTDTgdieeisHN7DnOiCK3
m54NKb6yTiNxfDJd6k28PuFyU+RW1iJQ0X2TrUKZjRECqjKdvzM2xvf0fS5cI96VsNVrsLtQwn4o
mBAwfX9R+MFY7kIHqp8Bp5p0Oivw0Xd0TRMg0c1XLEbvtlOPood+2CBCTBQ3esX7p1FrP9BbGLt/
z9Y8fELlLk049YFXwfA9NOPSxMZ9of3jQTgX6l/Tx2j7vrb/uXn8N7qG4VkesbWofSyGZLlXuwgM
wk5KpG9ybEWJw3ib/CIlXNS9f/6MCAHED7cOTQeU0X/2pr81BLUKpfoqI4UChh1L9lcW+Ae5pzAq
sbCmvM0Gwbm91eHE9V83JsRgZqul9TEYjcX/xRAXpeMbv6bbeUkcG3XMs0ntvv8Pe/5RzE3zx6V6
zifq/2l3KT3wVTlGWh40A2fprNUeKpFJr5N4rd2R9mnT/Qxv3rd8OtaLAyXuq7Ft85tQoOkfWxm0
SPbA4SOrMFfEVSVlpNiEkM+qzKht5Hha/uwb6hDyVguuY/knFr0E8GrngJmrI7XMkcoLSDxiVuLs
mAULL/O+TZcTOs0TXsyCl2M+h3Ub6c3/UkWY62CKbpyrTtMv1+B7bNw4+t0ZElF1m+Mw/mAYdNbJ
DePSV/lGsb3AbV93rq3cOYp7/So6Rw5jEEp5Nn8sSBr6z4V3ScZhQB3UjJeE2cHxzMt4jPA2mPwz
J+IbFI21bp/fh03ks1PWU4xOARocXxk507/4FKHgyrYwtc+sTd0rCKzlBMQWOpPS3Ig2G/p2YFU7
DuLPvoAKaYYiC91vpQLFXMqikRU3/Hh5VkfWWkrBICD1+rrsnH6AKA8taKIr2NbIMLBOWRrGs6RD
7hm/4adIqdadTOBE4nvLkUJq8bnsPb63kD9un14m0FqS0gZcEA4SqHkzjKoa+L+X/7S/pWXxFW7a
dE1xoQacbR0VfdAQPVDfwDRMYVFRthcLzTiHLnfZtJcZcK1xYO23RK0uTrdocabmb4JOO3XE52vv
XRwgEBqIb2tKV0TbUBseUj5csfO1o5pQIH+2SyhF6GaXcpKgNOdrOZm/XIez/+l3nVBsOxNwS095
pH1q3C/mzEVYKkpi7yzn7NXi0CrtFn+g5zjO5CBJDRIxhqFyUt+OLLcr1f/CBGDvXi2jOodhRnoS
I4siXEm874uZOVNSy0jJovN0GRRnavQ727kLq7R4b3+AGuaJDTxCQhpp6N8wAI1ccLpITC07TEa5
mlibYfqcggVV/fNkeaAevExCEDn+Qi3h9KsHUK5k35teaoYSZUD3IEr843GXWePZ9rJ9Jo15/gHG
M0bF8OZn5YDIpjk1c/94RX4Ts2C1pv/jZlxku6LxtOJU8pxDu15MeS7uC6cjgM8Ukp6fOXPx+U1u
gXTVO+avXwChYT2i0OgAe+qflyvduJU3JGL73khAG8nQ1KLm/FvZ9aq18maZcji7AyUKytU24qBV
Gk70LOik3tqBu/x7n+KWYqm/k3jWDr6/PXuaUy35yM6TBkx2rYkdegS6o/noQ/lK2r3/BtCQ7Vv8
PdS3/5h6XDZ8bM00Y0RSpV0uzsRaULf7Xy923yNFOSDcGoEbhfnuV5HlK7J7+2ELrO4om20Ewjvn
dvf8Bx5gGcnagvw+nF7EVSc7l6TDSCZ/ngLHNbRT2OTiR932qY6sFyDsMJWljBGeeCdzEK+V58GM
DumEdu37x//FWqsJaJHrU1mKs0/PqRW6vnygkdX1H7roncT2UvaXejl4V78tcyg/qO5GQkUeDR8b
9NGk/Ph6mWIx7diwMonuIpR1K5GjzYhgkjXxIwX/6Vro06X/aZA+MS6K9tgfE1BQCeQRBeYEar9j
jInSzwij+WBm1uO2R5kDZWAATqxEwNzhnk75/N5Cve9ErrkjeTPeJAR9c/kdfVWXVyMHNJlhXUs5
at5jSVO669wx/P1+FFUmOX46uTkBnSSl6LvO4z2yRO/Htl/nPkbpUL5PCx2LdBrAvJVv/vFRoP+h
4uxHSV/sJRVw8Qx+LyP4KclfJB8pE5irHC/FKZd9uHdKiNd44/NoAiJMh9t1MB0oZkYp8T1hUldY
ljftcAzHx7g2jThDpy3rUxKFvLcoADs3TrjOs1+S1zqxwy9er5huxlcP/IagG+3T5HpMpFgfjn3d
l3dr38fyecYKFn7EyicjED/R6u1edBPBmOGdb1aVMp4XS4VKczXBtj+q2YcYBZ1mGHfL8ZCxuYCW
1o9SixCtGoQT32ryhCKZleWRcqVY3YXB97EWgG32+A7ATT/Q9U2q6TcSUJJussQf+pAHBWobzv4T
MUkJNmrfMLVN5zIMcJl/9Wml5xOA3CCK1/Hd3ZDNDVMCMwT60eSHjVzWjSesUVhFx4K9GutItRCB
KCy8PXXcjf18T+S+InAifbKeBnsppyYZRNE5guINaleODGAXr3phoDj5dN22fN84fCPqfHJKGWLe
TjAyN4PYY/LxzjThx+vKY1sAQquRdt4S1sZuDnYR3zXDgx6HvKFovqIOAP2BpuR6QeUJN+Jt5xBZ
//HwzadNNg4GSujbYQ4Z/kpH9rwRzs5VC1XQh1394jBFKrag94Ja/zWPm1SJ4BFgsaleOg0ZdbAJ
USjdG5nm7OCjxieiBTz7AUryjn4kd0e9klosWzEdYZwKE16Go68Zvol9YSWxKxtMaRuJonPA+jhE
x2sA3pQcokpywrrd/dsMDI91QlgPn08Sux7EfSh7AJ+GZRux2FnisOnPdaOhv3bSzhxoXpBbfzRb
6/e7kY39Mu6lMV44TmfvCw/j8FIF0MUtWYSJrBctLbsz0spjAO33eaSFC6ZvheyUGeEaf/3rO4g+
FTjBAC7A+EZWZ6bSFkye2hFltn+FDuTL6lJWR0/prT/yXdtQwswu9qB05DimtgZ97kLyXmZDdHlC
U3g4ACFJ6V5k8raAlHKHJiiM21DE8UmC/Idb4/yOzy58WD8yGcEanfQRb8LJBJ9+BJ7CDHmWpC3A
567SUdsU6zd8dbNLiAEKMAcvVjLJjsK9rUu5CiYP3Gk6A5vRyp5T4Sm2ZG21JchrnZZUgE4Bbau5
RnuU++b+XF9BfLy8IUlju1b09i9QkEm+XSIRxmbuNLiXBsuI1ceelp0mlz5vaDekJHT3TnapbG+u
w3WLGCkAJATbDcNwQDgmBoNFBnq491yu96D51+fIafLYJpgfdugs52/RdWrNYvYwB/qf/4T5kyyw
bJvV+bsColMw9a9qvM8RVl3nf8oyEpExyp7eML94GA9oKV/rpGWZ2ZmnGYsFuhBxhnECDIkyf0En
NiwHJPB36kuRrkBNb82IAyqnljYX18kpO+oOc+AzGMtltjbBPBegvlLQVey6MLlKexBvcf5hHufR
1010yLVch0FtpGipoEVh/abXO+B3NJEhJk0TvqmQLBltjS7K9yEK2loDzVHfREW+7pxSzM1/Wptb
p7vFXFRmXrfL18jJBP/dzbAvEzl8ugdku84Hh3xbzdlMYBR2KRvdbH6+P21dPpiQ6snyunOM8DWh
6C7YUt8uH5PDSWQwZHDxxQleURdOMzxJtN6lkv91XRV45ENFIu4Sr6Z7X5rnBHf6Q/p8kUL6HewJ
pAzHeG0eBh+8LD1MCfNod+7tUt9vAfiMbDKbZCpUIadi8cMN2NcBSqgZ1tfrV52JuPDMJXFarAFH
NYFdFGXFTgnJm8fTsFUswvNNT1I2E+93qbXJx2wn0ARYPnDyGmpU/YnmkQNoZk85VkSxl2j6q4SY
nce4I9P5n608X8z/6/gNt8EUVZWe+fvmsP7sMZcpqDw9NKjnrbKmeTvTkc+qzYuKj3IadiCHTEng
HS1LJE1dFilAi6tciSCMMPumD0B+7wzjSi/TKjFXE/IZB5BEzIBRZyoDJi8X60/upw9B3fDDH+MJ
uTgzm8LScx6MTaIC4GRQ0BKqA1Sy0ZHhJBbmSMYIoA9xotr870bqs+yVCP7HLK/n64NCX7jUKxYE
MXE6X8B2a49xTygtZ+4FDu1sVVsuKUFbIY38suG0qL3d67rKqaM66j28BZ8Z+pXJNpRYFEVIt4g8
I4nU1ZD/ombC70o2lYt0GeXvYeHNlypjVEoX8Y9GafPWES3pt9dN/TUf+rjrK4KA6vx1eZsThG49
MvtMKNyQ5EjoW3Xe+SL1ftkZQqcQztJVsWLmcq5Qp5TH4tbwicCD6UP1nhkcp/oai1ifylrqS+1I
KVvF+R4dqoNbPxGlVb4E1xjJjIIAiujDOhLO6RyGhJgWZwzHsIhzRJEQVh6xTJuGWsRpVPOJjQpl
gqUuGDIRBGL2apGv8mX+5iX7heD8R55AmFOoR0slo4xCz/JJcZbY8Hd9rvEkdYtr/kLSyqx4SJ5V
QdPgIHercDU6Yi1HIydx25Ruqf25T0tBV3MPiA08/qkyF6Lw3iPge6u4P1Uil3Bs4ZbnPEOTm2TL
oUZoANbTFRdN0bsiLsCqxXiDoDdArJiDCX+uOw+yh10+cbIZFpu85eBDlprk2jFboab3kNCXI3ce
pAtGnLu7t/EuTAVPKNhpETRYan6jlF3KfCWPsSX2LaeLtzurj7P7r5rt2ByEfUCEgwt9rA0d7YxR
oMOC+OeBnJHYBZgehDIgHtJzR/UvgZG0IP3vPxKJbap/0X520JZCXwPATUTGvjKWbCd62GArdJSJ
GyOS62VPKe2fnPYR1fFP16QH9yCp1zQ4CPmKqdkWDbDvCU9mCFddiZbE7gc7/e+3cerYlrOYW8yJ
B7ngf49loP9FQ+ZRSpnei4+QxM1SXTKgjPiHWB1c21OrnAr3TmDUky49smdUG3h90TWZT08QUPw1
tjX774GnrhZVPjg/S63HsPvb9WtH47MIolDQWKmGbb6PZHAmbBKJpGpuCZ2QInWsptuc/fQOaQVv
rxoLTeOf91rf564qYi8RBpHZdp5ZKvVr54IZ/40dawOFPAgKZ95XIoRe0swIWnjj4RaRTKux1NtW
K86uXJz9qjkEluHrSyFFtIk6pz3KX5PQ4o0YOhUA04Dj/lsR2eBITLSci25LToj9suR//WZBUUA8
JrY6yqmHGzDYockGYyC4V+UwhDRlh86JFrTtnArtLX+O8JTOrbeIEftOom3FcKr2B50DqGfBcwIn
o/yGXSKUKwp87QFnyuohlNuOtrbx7ValH/YCPiklFoH6VhyA68touK2mn2OXTJOgWBwsXNaJHhrW
ZILCbItiznYvESWpH4PyJSkobNotzBxoYebD9RKZHeNt7UQuRwRSIqvbZ5ExrAenFXHExduYDwZL
WmpbDVEI6kwg+SDAvMrkU/RxDyNA0F3rW7kDUFY6540J7vb4V7aW/0CDsJVxYBDBpH43jce0KBR4
5mZJurNNVMJd4gHCI9u+vR1rXzemfZFXfa4Xw0geg1MoixufkhrkA0mn/XDsU7I4HU9eSqcnK/IB
OEpPu2paavder8oORrVJX1Ke6MpaXxVoE32IbxKuhsc0CCNYZz3kTisMijeVFnBrYezVjsHj2h5/
mNv7LjH+XjkJgRDqi8wTnqXu2PSxqDvegJ+EsC+xZNK4raBgBS67uvD7MBgSXaoW/33cIDuR6QF2
2uBfngZoGs2VqG1QAOQjP/QfeJLmeGoMBvGZN0Vw28OyIqciowE6PWNOr4mnrbNWLzhMC/kVa2Fh
x0cNssLyiQmPXnkhxVMo85hF7PjJafo5CfgLZ3YsNno8aye/0cCGXqqM5GAt3XsCwPjMKT9rU3Wk
qaGTeibCAoa9vXn0osercGlNMfRwN3IrxLwJCPXiezTl4mHA2Pb/WCSti2L7UX4+aUr1XMkx0vug
U2ZslOxKt0AMBdJ3BDY4p4zqmufKdAna3bTyJc1hj84CMP3GjBKnPFd6qOyHIM9i1F/U7waiifCR
sr+XEnBIrNhq/xeBtohh8vmlt3BeJk0upUv0S+KUAYLJkoGot6e1tOyjSz2a4aA/bJw3QFhACIm0
A5QIZzZiobmc+5U/m+Egh9U7z56wel/vBNN9qQoJQs93CaiupRPCi4o62DkMbUJo2mDqE/0JnRXm
twtX3Njz9l/zUKs2PZ3wYF/X97Isb9CszmhOlpLsIf8W5e4vHVeVudAMgxfUglA4oNh4K3NaYySd
WGBLENHpyto1S2hFw6svY6udPU4nw+W1PJKm1BXCg1AgyFB9W33HQ8kvYu0wEbFryNcAoSFnBJBo
m8bpXpngK6BJoH4wvJxO1aHlSeLsVszPzvagd7PHnLfaFqu4XAIhnhY+k3eX8Jr6esOIPVYbFH8r
VaPVpBecP3PYNxZZmyH1mSAxcHzV82SXWoySebU0UUu+rZIxaDmRmoS4bwoMIzpvuv02JGgUL5Di
TMaNAdBss+ZzdqtJIIA9aoXyxGnQZxrgu2/EdbNyFWoyFhvkkkMC7yATzNF/AE02gFW8Y8kqz94y
vRfey3j4U9O4oSSkpwQe9hneQwe1Vdgkc8pLe33GdbsbJXsFBNNJbmF9fJHqaPeb1EjqgMGvFPiU
0UzV8Fqxfsml+vdcUip8ynxwlnAwJMq4lbvSMTOwDoAWrDEfQhjwaqegzyth8EzHGh4GNkXV9CpI
WhlHIBHxHsX2VsgULY2E+rP1koT7aouh3fJ5VP1lC5K1hXDSx7W5NchwUk7oMvLHzFXfzi4XDf63
EbFGOwxk/R/Sj5yd3McUkqWzW9319l0DGuSAfoqUHl74t8jFJd9yzi696lV9Or+hVof9opsJeKYE
X0SN2ndi6KFN0odH1f6WOCaEiPqnMRi4EfEDBls/pPfZ85XsEdk/B64+/KDRLPUvBHbqsUX8WsGf
IZjFtECB3ru96zRH2/GYXFmJE0/lvdZX6mgr3NoZOwfSSlDk77SeebbW4y0OU8+Qopj7l9s09m0S
0G61duY5y5k2w3baVlEgrgpYMJowqcaAJzO6k5/ofTL44AGqXt62t0WBziy624Zf5GIzeCjPbR9v
amFt5jd2dmfyt+kWZsLdFh1B+eqY2CLYoyT5dnkmZoy2BZCmx35n8YxgM9weNpIDsPOJIO+m8aHK
Fiy6RID5cgzB0aJZ9s0wHmgYf+urGn7j57rhTV/SREly2NmkUqPX+wTCE6qkjEtHLo4jROp/UIOz
1KTZuoq2gn8xzt97ZBk0tGlq8iSEb+zb/4B3s+hJo46w0+0HwYLOVFpqTnub5dr7B3ebl3Dniq8f
novXId91p37zBGbsEtjG/bgkMp5s14EkYnwMkCdwFbrMaezYmy2/uYBh0YJtNDRvhIWI8a0k1FAm
fE8tzGwqMaODgpd+gfFx0inawibvfwofNEZQyc4+RGkCS4LjKwD8Ecr7f3uZ6GXldA+QkqN/tgSD
mWb6DOR+MZZop/wPreoEyYKl5B3hu9K/lASBPI/AqBeQnB1sJY6czhs7frYdmZfqkTWy50yysB8P
dainH1nXABrg3C+3DitJWF+BkXqiz6J2SXiI84yDmQDk09eOxGsxa/lPXI8FpKGsLzx1MGooFy4f
KQ18DdkJoBfBDHyOru6GKwZnipYxrgYxfggVZNhmP/rgiNbku9L/uXv+L78WGG6I0JPNLS/4n7wa
jvIf6HqJWht2TVEGdh3NXoQwo3N0xGZAYIYkFtCfwIiNDoEnkmOnNLycydlXg+L0FQnXfKZxBOSD
ioHjogzurKtDYhAfjFgr1MX7EJEApT9rZyheJJ7eBlfoolmj0N5VDBKRK57jiQ2/A5DAL/D6Jc5S
cW/GVwzlzGiWTLkB+vc1WUrofvA9pQuIAiR5vWevd/DdokMSLr0v35mioKaR6ki0YA2pcSRDq1ae
Zy6JpdMOJSWj+sPKMY4lJCmUaZctKm0OphZSLwa8VMWwubMf7eCAE2OToHfFLJASVa3RfM8sYNQ2
ps9n+qjYdP8Sd/d2I9SNt03fOc0uHhM2eBIT2/tNTYpPP4y7SezVOco0AiCtu1NaVrdPLFj7KoGN
hPX6uXBe1o+mspNG/Kw7Fxgz0dWj0FxTh1lnM+zPe3vTPQrhLuL53jyu7TtQgo6NqifCb0wxbOWz
vCjYLH92shpNjEDQhhYhyhuw6iUnnPGFFOPwVQOCX+lmpYdJVZNh/WbPI7nwK2OPV3IG7+7ogx5f
qhYPSEcbwTnBTkpAmi/Q0zD8sBTJ7gVzT0O//fOeV+OuNJO59Bahajfn6NnOBx70BKU+zU1wUr6e
WgGTxRPhP4ZtRw8ooBYXKjZ/e2750YNSndBp4xRVGO4+vjrr4JHoaKiybCA6dZdj6LD4MhlzyPIW
y0qlqggErgmEFiPRLtNrE3zhQ8VxVl1RvWOmIHXLEx941U7tl95APfnsnbQHH+YrP4xrLqttFbbZ
LjhUDMrA62vMFxJhet0942DG3XHsf9rfazRdQH7KoM2fp1zcxn3Bl7AktjyMtkufv5PpNCxF7KQk
JvjTdQC8Si6+k12VhmlF4JXY3T8GjYd9qJDySz1ldlUo6oKEAT1HB0KOlG5vPg9vCbYDDn/3dwKj
/WWINq/Xf47tDcgdXlVCRObGif2bXE3I1pWwPzMCnKYqAwrS05hmeV5/GMIEIOyqKaLI9Evd2tSk
IZlOhhRzs68ybj3Rk3nL9Mq7GwBVW1f98jI4lf7i5eV2G1oxkaUFWc5GMYo9Jww/fJ3YEw5MXbRF
B6GKUfX8iQuNhcKgiPlJBJIJHrUYk7pcq8janWNtgiyklYF/i0tkXAgNsS5YlESIG0ZFE38L7IBW
z4TRBu6LNhhKsUM93YBxnuHZqkOcOq458V9QFg+TBzEGyBN/5OO06Ixw7P4PbbDCxiLE0ns7kIls
HlMMWyJH+Pm4Dc3LAHCYaKi85jT6rigHE7/oeIz1ueeDyYQbC3VgYNbbt6Bac3E9am/TZonLPA6J
JKW5xvAKaaWKbwWqMR6DMFzGPNHvQ10OotiBXTEoS3hupbIWbz04YzlVj4ADa4T2Ac5l/yDmdEO4
xORrooAlfCv4hAqdgE6DBd20xWPW4W/zSr+xsrsva2n/K+O1lncF5Js7WE4Ro1z06hp0ygdbBIYM
H8RMqYSIGrA+JgVdx4/CdC3SFWLUnCpKp+uDC9bNi+aEeUSwYFIvIgAfyl2f/712w/vVZ1YTYPlq
z1/eC++ABsTIJrFGjzsBX9OQSF7tDWJQ38AX1sqOqpptEWp6uB/i2FrghBKnQauei+q06fDpLKex
hayNq1wh/5TBdEuM5SqD9rX6BvOrZmBIx4YhbnaktwGC51A76xlwbL0mxiV5BMVaxyQKEJM1jr6k
ummRsLWnmyuck3bi1U6L/dhjGlej8QG8YTfVw732HnRhzqjdrHkN7mQ0RFq9XePq5Ya5XK3cwnTv
zbsvWgm0u2CpRHIEcFDPQ1Gfh2Ri6EW43mWPDZIWjRsqpbr9e2iLmbjH/3t/uJ1MRJCYTNePvkbR
hDwrgHz9/CKugHN2MTG4gIvvTKq267H/4YqMmTVMOl3AiSz+qwdTqg+Tka9dzSYZFUmdBC/ZEJ+d
G/r8OlZweND/fa0Rv5CQGBkaz80cd58FO0itCNdIsdbSpFrU5C9MoLxC4uBwLcrf/Im7fEPSoe2G
ato7x7HhEcjdb4srZOEjd4M9pso+2I3Msw7TIx1CyE2qwyPlEQciLNL0MpZ3TYZUSf17wOJN1rQC
2jPMlaBso5HzYnWiqVbqNTK3vrqk1DEje77l0N2HB+okditk0dTcM0Q0ralj3EL9P9O3FntgD11j
tw4mr2MQuFi9k/l0WwRcXhbq9IsjMq/MHhJWQPcdJqCderF6h2N9E4GNLrH7Vkw1ggx4CGzyNuvE
LdnA69+NTm4P/248v3l0PnzSizGM3uv5AGMRlSeExZoitp6xMPAhPsYwSDxS9cAR/qhUyt61PPHR
YQRQBbJfATawZQyXXzMPdVvyO5cVjS91gBFUZ36voAmqlnRyxWHMfWKwTAnPErpX/mAFDABHb6Bb
g10RvYB1Tw581Jx7saVq0Jxoc91i3z7ilygR9CiaDdP5FH73bXVBe9hYCiSb2lwYPxktRRc8yiWc
ncwZlJ69zr12d/4qqDRR3K5eIVyQPzZamAwJFst5zjwKuuaiOzjfMGwBPlPptpK238IMO0NxzaEg
/FRnDv/OEvfqq9V6jRXUBtujZ/+ue1NXu3rL67aXxl5e4DBKex8AecHxuCGJmoLYrk8Aty8Nf47S
q1G1goLZetKiTf+i8TumsnYuUKBQYWu5chuOpI0rilptHHwTlbysPqnzNvvi9Bim0cOyGSH7pZ26
8iHZMnRu9oeqzxi33efYSSzQEB4ZSY848oYlb6oHeq02eNkL9BNz9w0zosF9d+8IkIwUZQxK7aeS
rBTYVR+zzqF7FbsIggCkbhfakvTTjSNkotYsdrSJSqKtVut2kgVkqe4ViRf039EqaIeWoukoyj8K
ZOjj+uT4bltabPB+qWB70Qh9Bsda0Arhjr5O7TX07Ylch8PiLr0lmMmBTzrSDcv9Szeuxcq/i4Tu
1sf6bUvek2u6wYxOFz/STWICTutmlvfrfhD7RyruIVUSQGFC0hT3yoy2z0MkPH3/9AUQ+Eu4c2eD
rS2xMgBLGJloWPfGXKU9aZCVY7xCbNdOA/Q4nQVslC41tEDQ8jDYAZGUlQ1a0XnnMhZMfkaaUhkg
OrBDfljheMMgmabka4wVYTCuzvfsyM6We1A0RJwPWCRHG1q8qJu+FLatmQuuG0h476oVUNiGO0lS
xDv/V1n1u09RGzyi8fIZt3yI5alO+Ogrzi5ycWnvGYYO7OHLcYrIytLQ1a19IvhE4kKc/8w6Fxl+
+o1DRY72yNoW9yWKT7jejI77cho7OZ6um/epvwxbHyd0kjUR/Hk4nzod2He/NNLG3FSqQa5q7Uzg
a62G+ZoLEmZ5Rlpl4tigZxuG/Ngcf3LGg2atdIQ6g2HfLwWMXiRMx9ipE4aby+/Xd2z0u9gy+2AJ
dce6IG3HaecNymoEgCHuizfw6mHIQY28DFJl/SGlT8yr3jP7gcFMgrV61DIWIbbO+0nmj3cdd4so
upR8M+lgdZMIImhTfoP3ZJTtoMBf6Be2Cc5ytXHKOwL+tOjTftY3Tnv+DwFboXVK8Y2Y9xoG780X
+5HJV/z5k3dxsv71TJycnyhKyt0/QIA9OmdsCad6/ziud1Tu0hGIWeoElNd7JGq4RUmuVeSBv1to
noVIHMOcnsFbASO7fV6MxXT3nEr4YKnnOHfcdL2b/BsZ8QJ0KC/Y3QpO2ODs+nqCjmzXwjOXdGg1
dWQOIX5to1k/lPeW5gCEZUMHewaq+AmLbzsguzo6v/8EuV4oyfI8LH8vKZuIFPrgiUtk33WhuvX5
8Fizkne9Sb06o/7DHBuip2Y+c8DzI3kVSqTtntCLEIvC7w2cFtWQ8T6glFOWUzs+dNvPKTUGjI58
/6QDt3AMtgXMozNz5AQdRXjM5siXJnc7SCueijbSfryXnqZeG+FlTyEDcbQxX/66s6BNHVp5r8Wa
7P3S2eDM1llVT7a1n8uMuwc3SwBFTY4EYDbxO25Alr8YpMxMmVX59ZccsyYIXfV5n0sWtd1QEwdV
2fl1YqHfVjWTuUxmltANZB2E58oj9Lard7yc12D35UhklIaDe97AjoMw0zEvr46ZknM7cW81qam6
B4I3rrv1n1wxocHZJHAIMuxlfUeAAfnVzy7WcprYmeXfvjcBytSt2BFJoGmcjUaLBw1juzpkgOHD
Df2tJ4ahmTkXoNnPO1vZv0BJF4kmy6Y1sRRcbSPAkgZ4eQPKDzTykjbjJ9KTOZjfJNWwvfHmO9Xk
GYJqF9f2MZkBAlweUPEXnKXp4rjklYc49DtQ4KkWB5UdUpmTZsyeTeH44DkQCIRAi5sVTLV1M/tg
0yH9jqjixoo5fC1oV3I6yxBsREV9lg96pFLUjgVzbDLYyMgsJNIyDexurd4QtqFUUOQwR48CTGWA
XAw3I1llaQb5T5s3EzUjZHmCwh2v5/z4m5PT8IpXpj8XWmFmjFNk+/XmuLAS9OvWf6l9ox4IYFt1
77kzp8BklcdaT1R94cAJKXfPIyjmoEsP2sp+9MYrY6B9rrpKzXeO6o2hgRXO6pe60mo1u2gW0zYj
25g7TBXldtTe466bkngGrSIqzw/J1gRhn4wvZSrHd0P8Cagq+63J4K7/u2JNtP2U+Gp1aVZJ6YKt
FP5OGbJ74abhGuXb0GNSrZEYHn/XU5ijCyxAUC9NK81U1F9zb/RRTCy81I2VFDPExTJTPqNJAb9s
ysgbK8AERLRxnwEGs8Ma1ZYS0Xv5qtkicDloTe9vePwSzoO1BhBOWgnGqNqTimtq8w0Ts5UzJ7pX
6ArRcpQXk6SpnJ1YcroZiYJqBytGx98+r2dqSMBc5m8gipAkbCFsNmeon37sl35+j7ohd3YXtaUi
I47zcHpjvQtb/4TnY4vUP/2KZNSVAxHhiQcDpkig7d+6DRW5ETo60KQdGbX4bgBkFS/dt5Yz20Y9
JT5CyWQlt+dK4UsRMQ+0awfcVPs5gRGt8Bd3zfje0fQGQy62cjvClcWZCeR82s11HHHwR2zQeDpU
nYOzGDqXvuifHY5cwaZtpIXP0dkBEpuxtmX9ZRQbDLyALqrYsf3tJd7waF26YT+NVhP3m8RG+qOq
R5++CivQYDbErrtbvCXiIEx2u9cJPZ1XNnzvAjN/+V6EOD55unfsQrepFFZu4L0g/r9BHkmOmqNE
h0l+VfR0KGJYkYNYd24igIlwCXOrbiS6HYqmCVZkL2NTjZq7Nm9WE7sxhCD2fjrUES/4g/SGXi9M
xfW5jUReU+bkAlUdBnBldPn7Vixe6yecbjDLCc8rbAQ8s+WqqNQnX7u7M8ihvoZvCkLdcuVfv0xL
ibs99qscQ8sJfRrGXqs3ZOrIYGrx03VjGUh+TdAEtGx20vqarMRvVQAkvC0fu2muBdJ92w3+kXr2
fGPcHBxSPCO3b0bS3ll2i1LH2s85p7Mxw/qHJf1kps47+VVNLeUBFdje6hMI4dYSKQ71VcVU6ITy
OY+9lSVJjidJ0oMZLvVifbUl8P+jBR9U8AHl2g5OFEk1DVKR28+pzn9mB09GDM7Ekm3KwODG6/0o
of28oSmE4x+qOa9u8+jXLk7+S9xXA9qTTeevQB1pFlmiCaIyFi9RUZz7Rz5YI3CSyPC0Ff5JQfBZ
9wiaN7seXWDAlnrmg8cTNObTRQUyui2ucno05t8frWQiwNCVyBDWbRl7y+/I/yOJtkVshUFclIs6
AgtLt4KeXQRYIGTbBJf023wZr32/TCSiMJA3Jqizp9GCdnZUqzrntTp7Yt7+jTWV//f9in/fph1H
Hh6SssHU5OkB6ODr/fr/0ZPwvDEDtmS0YT/9adJnU+FFak1jnfuQiPrqYE23q+oVm8F9kSTOWFuz
MSNjTf5CJBE8V8T7Z3L12ml0K53QwdECCtO0GU48aVMbeov3IyoqL+A8wTq9qPHR/R4NRd7V9MA+
VjxRoSxKScTFycmt1wFQc9Pr5fUkJyEjmNPiYZ+LhUU9KXUrIx8dtLyvaGpvy4d8RKrgUnQi0T7I
Yi4ElMx2w0SAEr+O44IW/l5X1qsonKXfap8s2JOFZ4UK7Z6hP7cQ6d41shj+m62k5tzLHs1Wf0Vz
pPj8Qs1pWDlX3NuxBrYL1qe6n4jtfusKJRh0C2NHxcvxBNpJFzdoW9Mu0Js4bj8U84+VCKoIge8m
rGkxN/aQUqL4VVqtY2ePfkbVU6x+FiCuUTmCgELTZV3Jy1EjNZSqwPlx+8d7TOkGRrmzxs1uVADi
xz/F1zBGRn4CH0m2OnVdI4lBKzFU83Q/c7ud+U+o3usuZNnY1vFF7+ly158w7Xb5s+l1+8slf2/u
MxPy1i7UFHbGRjsO+yqj9Dh2UI852zDz8AqfqwdQGCjbcRYdxLtPG0C4B9hvBL9lp5wGRKxXVVet
6UNJByfJ+nFLovK9zpFz6Xw9xYoB0Yb8twPfPRbC2hV73B/eie5Ehs+gqnHmqwWTV5Vt24AzvCGE
UNNDuVanMZRIzvL4caPVq2M2O0nRg3S8El1EIyZDzWHB+W+hnjtyXECa/pzXwWYmu/rx/4ctIbsf
Rvq76JxpiJHxqQuh/1fWaEeh+KGDOQvX6dfD24919Lkm5e1fDK42ozq7E1V6FcQLH3btvr+1Vsf2
1zzH/LepmnqoGjgxop6G8xg7zE2RWLPEH2vb3dYSIhdvI2Zqi3HfVYkgSGxDrMjf5uGzP6c8hJTv
ed1R9gHBpVTnNOdzq5aFmvd6upaJgqZGz4+UoUNqbbYIhQPES9JOPlRKYI6t5Ajxu9xSkOYRl7ZN
M/nf3KQdIArPrc2rhWH8cMgSIvNLZ20XSdPo38lZLxkqtIkSRqfKfrPSjOg5SLIxMOkdcGbQAtvY
uW9/1JDD+ouIPGhGYQUVP+qlfUuYTjFsF5ZEn+tDp42hyxXR8hVuhatm/fw4SnJsNnL1GQHzwAU9
/qzymb+/NH3wkjiPCmzpwLC9W63HDcfdEkRpqAj4h+lG66hhwp0o80Chwr7QG+/4MFyFtIACnZ+C
7oXgprCqwi2tpn3mB1r5sOGoUMHnYNGzwT3tTEGoocz7URB6t2/knipFNUgln7SGpvcavRkWjon5
y7hSNHsOGL5nzRifDXL/PESCVfrFfTLYC/2Cit8kr5TkEDiWqBWoNEfAIOfWUlpbS2lVvlWEPztm
rVWuzoTyLNpIxoE15Dr0tvN3y2BZaKpdvqyUqTOrhNKECr1TMJIH5mtCaMjRVWDwRGJrX70AdC2f
iU8xUporteRMzTgGCJ4f9r5OA6YGo439H2tjP/004jZ1TvVwO7gAc4zs45S8uMZHwT07NrtEuK1H
RmA0u2Ip+LbhfTEbIbeQCWI+2bVQLhFRLs7SnRKnMSXU8nxY9LsbuSMqhaYSrfFxNLkiPRxjgNp+
dAI0/6OXXrm96GmxVYDU/NCbdKixmE14gr1YmlYhelQ5dVM9pVYb7JiW1ypSrJB9sWV+drpDwC9S
9VTtwFgbXZfh+CgMBGcdlJcCrEq9ExuNyAO9pWBJjNo+r7rLS9rFbMke/oYICFah+LtaJthi1j5y
WLhZl/huqQ/8IsMsl7vf6MvqjxY7JkrSFaq+CFKLm9cRjdNlBwpA3T+2fc2nQBWG3aKdgIWAx9iw
g9/f2QDAiB8vm6hDvz/0HCeN/mJeBU1KRHKZN/gc8gNam0dL+q6j6MEwIzvVd+vCV/TLjrkwWr9J
Ls7GWwraqH7/kg/20YnhAPXCEQUwNYiNqQNOzyCG4XqYD1kBb+hUAkQNJY4TEpODn4c1N0gQAbR1
nTtbFDD5V0Lj/UYF1F773SoTfsX37h9FXq074plwO1N8Ciuum0nLt+JTnI0/8RqajQmZOu/5eBJj
GzoDuIA+qkDY63h3K/71uIoppWjtlHWdIdMAbgmR9Rm+jcyWbBHylESoPd1h5EBcLaTBeZ4yhUZj
vhe7d92eMqcLr+tk/soYOmxKGswYJ5PnPMxGgG9nnlzP4YQ0OriE3j4QKwbf1ARCBy4zVPgL3WFX
2A7OAG9FwP+kcfyjYZB3vfZtFAjuJLTscJ3WU5SnddzdbJMbYHAallj3wJ21/6KDv4e+fUH3jI7c
QbtvI1uY8FEry9Iu+k3IvunQNUeDXZ72aWJmYdH5IIKoNn420WRVAiUWk+Vd7b6lC6dFTav6h+Xt
t2Xo6KowiL1ACLvF2SL0w0QaJKexKoLM0YwXCBlUGZdb9lZiysdiotDV+ZdGTHqMP+UxSJAopHbD
sRbe5vgPVxN8fwRmev/ZFjltAKTrtXzjW77T7JdhrRGUSexMfg44oeoe9oqOL5F/znhqmyxOQ52s
kJWk5aCBiNCDzSMY2q5V4eWn82WbmaH/7QzTeq22b7Mj9rd0g9Pcz9oenvbWYpmV2c9/1QPemgcw
RCK03AgD+nsZABqewAD1WOtEmTtx54SQgz/1tRMVdbCRDbSptU8lBMqMslHCNxPiAu/wMmTTBB8V
K2/dwzpMfQVgTevlIim0kIU7diAGKmBHB2s/Yp4esREXfvO2DAPcdcfQUHdUZYDExesQVWB9Ik6h
QQCxkcgXRCj7j5sMngeFrSrA2iE+116COypE/61q/kEhZxUmrhpsOuWvSOYegeAHD6l34ZFcRHhZ
Fva6JGheCiThVWF7RSjvbA3GJEZqNb125nB/JQovAiwlHxKwYbe9Qku73tZWZaPDfL+HkLCPbImL
wDKa9I6P7JW0vN6pOoFAyc2f8XsPMku6165VCMvymyQdJy/Rc+65FacekYojVp7uWdYVXVplSUyJ
+KcA1qxpUbSZkT6FtP1CX4y2vzODochJqNiTL0b2Wh5mVtcey405xTw8G+cRqhobQYUrQTAL9atx
NV/z2HVXwbLzvb1nsbVZT7cCIsf4AYzaOEwUvKW8DY+G+LuqBRKvpObNeT2rPUgsPVk7mRnTsumA
EZFZnfotCER60PhGGUJ+777Ba0ZRo8ycEnD75h5hO8GM/1lKPYOQXFMhzrdMcJ8ofsLH2xZIGv9O
kPDpusBcN7WTtfU9KGyQHxgsWHWLogsv/QajqysHW55yp/Ut4ZfG7v67ffrpbG5XAe+JhChKdmYP
3Xj/80v7jC99f26mjuIGDPE0xCXSWHxtSSIOi6oMe1uwLZoMxcrAgkgNcs7Zs8dyFyi9MBCgZCS3
BIsZLRVznRB7G54slnU8Fy0lF6ZEGAe0t4MMjYfzPfEZqmJ+LnFLR5CnK1Z7jBzlSx7igOdcHRAq
Ecl3bIPXcJ44vmx8wge0ZZxc8p2PzW5GNS2ejhXVngbtp7lH7aG/pm3S570DNVOz2k+eCDOppMin
dFK+wDwE68CkNjiJm678VcA6fhQlR5YbMcKzEMIsFc9BtbWyu4GnOJgZx5WF48EH1RqrdDYy6jro
ehdBl7Tiaw5C/bF20wpGyLA7K613Oj9ijdtiZiVUgWSSQoqr9rFjKVOb3v9Q1x9LoooMiqd3zpoj
FlRSd5/iH9el23Kw7wzQLb30jetflQZUZ5W5A1sNzPzkCwmHK8bpEiqenB9F8lGTKUfFMH9M+EeT
wnqctTi8aDNkYhYfqS6j95qRtA0TWHUg1BmA8ebs8iychORE+lETzfdhQy8wXxerEUfv+/9I8HU9
9dTB72X2Y7P9AHJzAzmpL93GAiqtsH4vAcgVLgffPOGZ60Yqa8fujyNLKj21ks0ufkQdBkfdoZ48
wbWCPEB36bMn0gspxC2mZIo7bcBtgQz8XE7n11ZAksDfOJRlZFytfqA29bQrZEyBox20DDYdcV0q
upKbhWPAClybMKh9eo0fhAmgS36RcOTh8GxctNOCuLafqi4/gHr11s1KiHE5KwrNhRQlnkcwuoDA
SCxB8pAS1HlJeeEJYODmPRXz5S5cAeQ0RZR0zIKk/RKTNE6qLB6l5A6guYuJT52QP9JJ7OE4SlBM
VjS9j8N2irtLxRasKfalZ7ws4bSX2+ZlfIR64HEIvh7hBUExJn0IxMt92sYzK/f6Gf1HYOo1P+V1
0OJIyTWDhhmTG7FEuASbMKuHquTPufLWR81I4wwF29HJ2grNDwBV1ZlzNILQkq1wcVwWZ0myMThm
c0IA6aQDCpAALExKrGsJCEUb1kfbp+bnSD7jLB86dUJ2LrjEvPObrMvMznMctYC3qaTa4zHOK4tb
70YFiwasZOmuXC4t6j5GLFb8t8gbPrJ1wFz+3VunmhcETiAam711gyOpscHV81HJEf5GIR/eT9S0
qCVSuixf6h7mVOxsdlexLuCoeelmUAWhEJBLq+HvthcXLBxBb3fIrmIV8FNVh+ib6zasX7T6cW3N
Xl8v+jcUDaz5pBd1gP5hejzIiQ/bOA701ETJcx+SHqZ5PavRv0FrOo6G+bydlGXS3o6/EVBZzd5l
wvAtMM9irs/xFdAxPepOLQZqHIQ3wl2NaLdAhwX030M/C7Op67MCbUDneWriFYWXDPehlZXzwI5K
sp5Sl42f0TVWDNmlh5mMHiuYMzTUBxypXQ+wO/udSQQaPVPb9cUlsygzWFftJv/b/eXP/f0+b+yc
uj0P+A61Y5XU/eQf4opirWIGgRv0638YewLKtPtFfULQwDNY3VEwaoCIK3BlUl4YqWHj4bFSvaAQ
tP4zkaE0CwU4V86cUbunSFXDo1qqKSsL1VQLYm1UdJUQ7+Z9x+/NbiNqMj6K0SxEHp/kMeE2+Cz8
uAMmFofxIlLGtpbbrVEGwcF2PdKpv6/CSE/TuOpq5dq6XtAmxIEyiodHH1PwVHcAc0mQaYyQu5Nf
ThJchRUS0lDl7uCpCSXNXz6vlJb74j/mU8oEUBKb6qzn2DQLVUhRw110YTSBvnt0K6C0/np7bcrY
asbO6aWFvwZuqU8qAvfqciYFvXjWu8cUcKzc3G+zNY8vDy2b0HfZAj6Z9h46oQptPgirY83CnmMh
7v8z9J7Iw+TTsELx2sv7Y4wz/9X1V0mvwITZ816w2EA91YgX6fVEvsA1KdFFDj+qpP8Mq8x+b5K8
ED+IxmZ5+7Cml2xXzGukDI4B0TB+cYMGtH4Qbc8EfYhPJgl9w7C6VByEY7RxgXCQcYoJYYsT4IyB
CLlAMYJCs6DQOuOIUldiMKin6wIhX7BgyvSAEXeJepFvoWscKWFjGaARLXA7fNvl2v5LRnWVjOSf
iDXk87FXWPczN1KiANO4/WgFa7sL+NduMZtlooc400V0R5EhlDsBF0tAYc94RC5f+vkBF+PkXlw1
Fv7VEk1zDA5H6tG5p/Z8OO/EoXMiLJHu5NHOALJrk52LgrraZxnHE1ilYwQp+vcXP1+Lj38WKE7I
fy5JwMOyYk77zfPUgwo1nYn9h4kjswyu2gMJN6vfcJGZ25K7yszIWmeQEkaHkFo5Qc//YBWlaTzm
8/1KQnrU+fOjWINUgXPmJqsHpgt+84nV6LjUejdP5Un9kZ+g94S2mEOqNGhIHDvURkBW0H94TQgu
zt6lYTfG82xR0rVF3cuSt3DlVou2JNcmSs0HkFT2AnbqgxUG4ot0bqUkftZqwOC8t4xU4/YW5T8I
/1klHrAROoa4vk9TXSGwnaprprig7dhi3FTtrIhsvVTsJ7byc7xpkDmzS7VVKReUYKDieBevRo7J
7HpUqN1wXvSQm4vwcF8XYWnoIsLZeYD52wszBPLUMuBauI+KAR7wpQAoRXXKMsDCpbI3yH4IsOn1
Mi76Hwe+01QDGyXuw+ewOALaoG0cX8kyeNbDnEjvqV14+ZyseBc922VlA+PbflsQQADpN25xZ2ll
yKRs3QYOKMTbYCdr582uT899ub4855qJGf9Y7aX21eww+OwDKJ81Wzp6JVcdRNZx1AH2NQYuelNJ
hwESH0Q6QSck6vDMa/Qx/eX7SPkdZ+UUfzUSis1vesAmtRfy+h2ALSoMJt9g1efnN2I2j7H+3Fr1
4vUWZ69BZ1xd+7apt6CJ5HHdGhIXN4RErdqRFFZGFy4YenNKHRalWqaZfoxyUpJe9I8LlQQrI6FT
Rel5vq3UnOdWNzMIfulthGE34ecfnpv1cG2oJPBozkX2jEDW4EOvpQf1DeqX/DM/GCEO7cduhIDd
qcbDkjcrPKth4I1NY05XHK8QdRzfohotSLt+8r4mXMcQtVqN46lno1jjA4nNL4zXy12daww5u02w
VJGWiGgxX/mGTPMpZrU3XERK4LcVcrWBQsijTesUHKiPyaz1XsaoOmIG9Grn3T4/uNFU/dyzJ2pA
Kdn/aMEfxeOmuvLndR8cGS/4sHsP9zn8Sn6bjUx8iKXZXNlwt/uOYoqsXGHFQl1icwK0po/p2kY3
jaU3Tf64gPs2mAVYFKakVfWed1jogJSBmXYd4KB8+ols+aTrOi4kYf39uEEnoN5EBPg05sCwC1Ea
ffJh21MHyhbgRrtazMUkTKf/x+ridXeWnkzA15niz9eXE4zlI6fV2LKP6lAZm04XxdX/ZlVvVjwi
D0KM4fTGFtuD6KWRIeGL57zJPKA1cSvx2U2MrcgOdcFXOmAl871+gJGSg4RyL9a1YI1eRTrvs+6i
MbfOQBC8v1J1MYYgNShdX9hdf/UaE0fQYD5qUgOGqI0EG/Av2YVkSrc0gCAwe/SHWY9lj8xvoxKp
bIdpycpQ8bhruccFcHpwfDD9oGNJR1Tyo4Zc8QA5nnhUIDlfp6Lb+P4rzs6d5oaV4el4DtOJJ5fM
cxBPAAK5bpoqc1bHnvjdBzG47kY4/x4Q3sqnjw05QhXM3MgtzZ/9RZF/yrz64KIU3yCYfhX+Neeq
snImCzfiznTs1uuDr6LEfX9q6wbUxk3u/ayK9APGLMKwGENTRAIXt3zvoBworn5TF/PEgsQ27fFt
5lf2IJcJFm+r3PKAFHHQTWF68cIq7LApiokZVjXSevsxqIrpV/Cf6vT0nNj8OPVOgXNKalce8ZSo
fXa23jMPi0+daojke663rGDGsP62Q4aCz1zFeWFwNsz+lnjGa1jNdZuUoYwqaqkdCCtxdCH6AV11
B/54XkUi2t/q89N093DWWT3deFxpA4LBwXFanOwYK2Xxd6TczAbSpzQzQHoMsgAeA+l98HOYar+D
fikBm8oqYwNaf1EIkT2xJeILSCP3efqzeK081hipIp7yi6KU1wZEAZsOmroyMesOPZ6Kl4rjCUqS
Dqwe8AjTankFaNxXp6CPKLCTAaGnsiaQRjqM/m9TfVB06gDCaSRtO1RGEqldeKMLQfga9L9h0pcQ
H3Vig1r5bTJbQ2IoCdT3Zx4sdZQQF2zUoR0m+m1AkiDYt0ZgSN9zLM5d1c5wfH/uVLXX69pCZ7dN
6yLHsUPlHxu8bZU85DQ86DB4352AAwO/HYviQFHwoLSf5JX1UiKr6zg4EHT9WoKZCs6VQt5ON1pb
cdFGMmHh9Ch45B3kzfZ+kwL0vEwgPzuq5Ej7Dr8jxjuVm7XV5YzkTycpP8Z9Yxg7EqIH1Ez5nhMO
K/bPdJbc7B4QbmuzHsMZYI9q4z2eJdQxKrRq3ZNCjmeoEcpbFkffN0W3nK4hz8oe1Zx8+moHj8mB
r8GNMSMVi+W4ldc3+JDuSS/LZO0I75Je1DDayK4RXIJ/Rhgbh/ay0+FYSO0+Z/QRScTCSYov33kx
GGzei2eir08faFFPSZPWJWpaun9upmFj2v1GS5QNWdBEH8/NMcs9PD1+hkGDlhGBKmTO6iovbJQi
GUCbASueCdg3VRegmUUBfjwWZn5FiOk6sPjBgP31hfxZwutazHI3JZKsiPq4grpaUruxnRObFNda
FtLauVWbnMQrF3HvxChNxNyM4syduZtYaSVNQJ2L1NSr98RTD+lcEj7OYzuH/AwhYo16vSNAZ44b
o1RDTEvt7wGTc0IC5cQOJHzZaUWrPfCdZb1cQuno18hl4bVxjAkRqhIG7SF4l3FqT0Dz3W1t4Xwl
fsg8tfHoMuANJc0hBe9h3fj5jUSHc26UDniUd9VTz+sxtgHEzbGzk1Y4uk+Lchprda887BLw7dNT
m9JiF9rjH2Fdkp9ZIxUelWsXZWKl5dsEPeMqMQAZ8c3Tz7tAtQ5GM5OtDUoLeluNH6DkPCaht9xG
udw2CH/BSVZe2jtU9myYp05PtcjQZq0M3rt4x7yoHYD6mCaxhg2gULjpjQyI4W86tsSXfxi+HdN4
HXalPoYr7xrscbj4l+vVaS7DA+p5rqWhpGs3mrWuAfhXUx/j3wj5DRtrsddcdAgnp6E9FPLqoPnj
u7IIh7TY+2N6rjZE2X6y07QNiLGNA2s7JC1Zwn+jbN+WtqZOj6Bxtt43xIRVSGArr/+HKRf552qX
ZCWc160mfXawaWX8pVFykserY6pN8fvmZV4aaPmuFPDKnCjLZ6EG7drQ/zs633aSsSl7oiBFroCN
5PBe0J+KlsL/H0u/3iH5yBv9HQjW7JB+kQ//6hUKZbr81iPPAa8AD58LA99/8+Jj1oRGRweVvM1y
xR/AuL3bzgTL2A+qjlE3qZ1B4HCruSsq3YMqTtJrPYFPXCJTMyp2NE2DVFjQjcjYVR1cqJuUBvGI
VtYCJbhfM4gtR4/RsNPQRMRAouX/VKJiBWKTJmX92BaM+iFg7OWNDXgMVTWDwy8WrHqgY+PbpEkx
1WTy1Vg5C2VGVx5pWbZRzoIW7mAq7ksZV8AkEOq6NGDO67n/TI1yPXCYz7DjgvLi2+hHOLeyGM1m
ClI1JAFhpbuEgq8KtPNf5t1I+y8RjCGE47KK+Q0i1X64dO0wxWzRrCAd1FE4XhjLLNnqIjOHrqiW
3121xs+dbbsS7dACW7jZzLVHKco9zLhPc5UpnXSyQCUwDcGb4FplJeaiuAXKvs7xHKqTKc+IxPwd
K1Z3nnb12ayVAXn/ssDnmFmbo4EBwqqN31rOlYlamZPHzZLtFI53gT1zERkko4aYubRVfazCbvV1
v4VCw/Xfihgmal+JQhyfW9DX18NaCYPz0CECMaFFj4Jp5bR+iKBK6n4Ud7/LvPTJZmEwBAq7SC4J
pXoGgCyzZ5sgWVEznMp/hkmitruugeR+gw3rXjnI2kbpoXfZnUPJziSQS1HkAWCO1J88d287sNHT
dJoYadsR+kHSNhm8KUJ144gLIVwwdSEBv+NrX8a5CWLjhra6jZ+04Qq1C8F4HDYEcB3I9lCHsScl
wr9kFtdEV1gRYhjADiGTyvhBPRr2XbOY98kMeem6b+ph00NzloHn4BnphSltnh1OA6cu/5TSXSr2
2CGqwT+IFclWhBpopIGZfCwJAt38td6roRmddaBO076x9EUpFZBxQ8dKwxFVE28LqghTwTy1osDy
OMEd9lSTpMNhTpx4mUJT7BDyDvfM0MKFiABIGRLr8b2xIupGSrU5K9gyWP+oZAHQ/RxBt+3h/jQO
9vpIu9cK/A9PZHabl2PIh5MZm9UBmNZ0UCwkd4jLjhC+pmLQLF1R1ndRBHbglrtbgzHxyr9HXIB+
RCOK/UCJa8zvA4RZA4xDeZB/nlvcNnFAp9AzKyVQNdUI4tN2+ycIkidyS8/wakpGX48oBOfJPfxg
09mKvf9G4exeRiJCrlF85lIpsHUh1m9tFww2Thaa2J9yEdgqwc87/Ve4QhkCC+ambpMeDOCP4GVA
UriSMZ0NeEqg9mkOfFOTM6gzxkLvu1WsP2d7RcEX9swpzBU4KNlRbsMjZsqwVtCdOw8p22qonIfu
RL58UZpobwxAF2eaFKxbYyIyCSOnIErQYtFLlLPEqXq0w8Cvboh0Slh+Mqhw/KosvsNPSuxgySrj
gFuNcKYky7rZZEMcenmKXWiIvrLwIY9EDQae4nZ+2TX8Lm9uG8jZ6A0JTCTrO9KOZR8o36hs2aZs
g/XTY7my8hESKyivs4pZnEU7uLAqANxIuKcmOIEJ/C4ttby8b8UuO57/mOao7pIwvnl7Rg6y4yYK
ZrIoLcKBsCxsk3sWl2xDBcWyP28uc8jB+eml7kfBeNsioj2i3Qhx6xJ4f3KltDuj4J4ELe9uiH7O
eKzZ9jZcIw+nTDH2bTlhEg/CZUeYCZDezQkUCGvPSX3Jg6XuPYyjpfi6OYKOq/oW+jWwrALVeAFj
hNvpBnxnI659DWqiSzXjvOc3lPXcWWSCNwQMKsfUO9yx8KBuKAp+z53WG5RBpzgsrYoGqzmXMsYb
e17Enooa13wdlpSKHUIFa+HoaYumr32ybnYyIla8iTU4lAvzMhgRFgXaFZ+Q6Smo85rv9GDGbAai
lFgP59mAREQXx6aX3zRqsz6hQBaCYNSTYo3/U+b6ukCw1b2ZPD+jR8PI+WqBNC16sDWCWzV2MmgJ
zvZJR8p70yubCOFI/KUJzPLbPz5Aud9wX/0BnGVhps0Wl4EuYj3/13uLKXHJTd7HCXjAMOY1YU+X
U20vOu9CRRPiCcKYLmUupgNlba9ObaOS0tiZRrCT2IyPQW8DawlRDCjED9dlXnRo7rKcpw7fK5Cm
s6i2TuOxvkyLwKpltKUj35HgLBt1FKTuayzcwc7woq98yAQtTFM8nWA4LHrbLqQWWfMGTlSPQ0eA
Y2E64aCYOWMdEUfcbE+qSOtgkKImJrWeCvz53rcSk9P6qvliFnxOXiP5v66b+DG5Hws4zPuFTbyE
rEPuRM9d1zpDfUTzRaFax3aLhaHGKorgZz1tFARPq/G5r5oPMyS/jw/ya/Jog+7G36YFWanx0WOc
c4ZkVEZYl6HzXUZrfwo2EB2xpcSuPvvNTF0z+zyLR00aaVXwepbitwsAhdQaSRgdE6VZw3dOBHVg
tMyyUZRr+7RkUZbIhIVYt8RW+e31/yuAg7VxmHihzLO/mtG7UKDrZpu0jezpD5occo5GdR0cG8sd
v01FoSS/iJOHX/mx+V920A0io6SHEUjrErTwd96Fh/R6+68Fu9/t90uD6M7416DF+YAa3UkIXYuB
looncTs+wVLvb8w+ILDZjTjKd6A7UyJH6ZJWlPtTt6b/yDhNftMFxtpK/TNpqmCq14sxKdW9LM7i
IvV1QLrp5OCnXnYl3iqtGHJv/t9LrL7hNjgsu3ZQeAL36C/qjDTsWa7YLm+cGbOHCrPuT+wVwmeP
CbnQASGoJZNFKSQU5ZdBMKc7vUgo8/SqpsKr3krkCMW5W9OOLw0bCMOWYs042lV6WpXW7u3slo0o
AdAe/hWF1iVRpZqdWGQrtolHtCSRDyjrNFvQVI4wAfhhD098FhVxT5EtWNquYeS1nMJTYzj5Rrhw
EUfL5s3cPh8cEpTOKzNfL5tKjZ/n3D5850F3LxnV1pX1YvjaOxYO+pZqzyeNyJKRc+yhDZN/K8de
cFj2DJIB2wmcKHdSOZWdo2ZVzrndnIrHvULFo7GwGww541CEZhfhr46T58dQ8SylhzGwrGizBb8+
LcCnIaLUXYh3reyn9sxPOmKCAk26L/+GMFsjojt1eaNF4WM8gRqv0fK74jgrLojq3Nh++dA83qn2
AHw2VK8yFsNNBi791wpOUYJIhtnGRf35bElQWn+NjB4XgC1NC/0DNDLEKamahHBbJO7hNC0l2dcC
Rp84E5N9EjvDURns5MhHPVCB6ZCtvTpmnyehckk1Gi2vAyHZciOLOAraus9IU1zRXvvTknG37ZMg
h5nuuF58PCFs7MuReO053jOavM0CCPKpUaIAA3zUvW/VuCQ89liOPojKbuYiJPJRPbB5hhveHMpC
66GkFA4nOafGooVSn2TCJS8E3JCZoH7GjisUV8NyE+5AngArsEk0VGKYsRV/W9FpyXj/kMkG11NA
Y4b2XziVD2+tNNZJv3IZv943KPmCFz2efSN1ZCv+TLUp3hxqd11JG6ba+8EPA623JVqktpSJV/RE
OzIEXXTXT18MFDhq1hGo+pxg+yTD30nUE/iiO7DsqijjZjwVdAhLZgDl/z4Vx4nT7wDp6AQF4Cq4
dfilQfEplDRo2PBdTCQpLLgNm/ySy3jKcmi8KnP78IGn3MuqD+9PPrquV0jIqKe5NOs0tQp/MHc9
1emLkGxOMmK5Zr693kHzA8VKMv5AV0CROrb0AjDWWGHnyeQT0r57aFeatik8VEXmxfzJ9lih4N5Z
bmhlCGVlNQ+SvoQrqqCcpHlizX3YznYU/GuvjZqnCNa419hjcssTtgOzyAElW8O/oJBoh0U5lG8X
m2IQ6CawAIukMxCd8ksdphqdTC7fZDcgNbNZYhcAfPDmlhGVrHp0EL/tdjRklfsWbZPNpEBV8IVb
joMcmLYOzX/z1M1kMC0VOPB3OOGur9Rbqp7FHGXl4htl9XBqNX4heQAt6iJenVGrwhTb3MkvCQaw
EwWGRorXElXfEtnko7Y7qQHM9k14qUAmm2mbFdboBXwphmsF6cNJE1+mAtUexkiu5ZCV0sQG/nws
+bhCFhIBbuCCKtZiOraUZhfFkhX4U0iCH2Rf1ERCLom3DjrHSBqcSdsYN3rLFgZgJfk+MDVJYO47
4dy32u3/OcOqHoU2ZhY6CVKqvU+0pfuJpppsiQFkkAJPkINXHM5+eAdmEdyu4qq7f/pveBYFuL2d
VVNJK4zf0heHUpeT9iKsnCHfrlnTzmJY3oQKQnweyR61INj+2bOohsCEQKaOFtF8V5qUvBk8/EVe
upYBVZz22/ma+4Eoxz777LeyQiHtwrjlCAemAuWqFSuB1VcFKONtU+r+9jYR8/sPszSXWOuLL0QH
FDnL2xGlVS63DlvZPjCfHmN5rlnXTETTNqgi/af/iSx4sngW/SCz4f74OcjSASrytCxy8G4G/9Wh
DYCkZdTO/5KCsCYE0+VqSEWak203TaBkkRnDLteppRE1FMgkB/gOIBes18v3yn47EwcklsyUVGz6
lO5l8LO3S16FDbh0I1ILpzsgLyIp9UGk9+Sw962Smesxhlb0auQvOB7EpOfnQYbpkvt9TMy3kwPw
QnjbA8Psjb0eWUxgqxnrgsO3tGg/LZftuZ+31A2tBv7l7fZF1HH5qQpzOhXPyEUcU0vijNSoepN7
DwDZgfMCs9/H6dSjeHJTps24+fYA0uAEO3+QRztNfgXLVTfd6S20tJ5a2KH8N8lIuyPpKvGRZvfu
lyST22bdKB9mnNHFuPYAN9iECfMSpjja6wfYSQID+9YmVEs/w7AzFQvu01DA9sydpFlpXeqGVUDt
CbIKuPplnWe1CknD9WAAnIBw4vCV5hy4OO7KDTTXQ1LAhxgmrfQnC+9nwMiJYYYmRFbK6c3VwSm6
eIM0ZG6vasyePDk27n/6Yfg+K7JR6DPQ4z9cVXUNdDcVnDcl2Z4ZqGDAs4NyfyEMbqURhdaFB6Nn
b2xIkVETV3zch3o4p40zZ2VKqSMBRgygZT4CLrkVTqihsKKG7xOvfq8zKWV7npx+uzUBtBWoykOg
YGvK3nqC7RlgS9mypTXVdHwebC/kdQ1D1/ZtCCDq81LqOjp0XbyfJsg21imX7TrOetDuayhXsRRn
lb+qFK9O0jITQGfosQZwJt/APFfOZzPOZVHX+d6rkuENcDcjaV/evmA1xC8GiVVz8DK6qx6LUtFn
D2pd9fK3/ncyRvy0bjbphgH5IQ8jtopUKipHFHJqFJwfk13SpThhtVxROG2K/w50X6FH804hSKYQ
32DWM4JtGRypqjvRZtrtCsGdkEosPrfKTSM9jJMdVg0mME4koWC95fKRWthmIq+oFQiu0Tneqkj6
EvgRuc4D+gKcnRJG5+JAB/2b0bAGEZNNkRcnpHLwSAQ66J8DjRMcEiIsKbUBWqNgA+Dv5qKafDPB
EldagxDwvGod9osbEZW53EFpaD1MuVAIyndXXyEHr4kqeMkZoR5oKGGE1Wy6T2GvhU8IP9lvWDnp
9UhQ5Hk7iUC3XYb/2wHvNMv+MdTzqEj9s4cpTlq3dGPdemA/KIuIBEW40qo8ESpczJJdD2TjbkLq
cbffzN0/yWGXeaSnnz+liLW/4e8qiIQH6M5xMobsZSacmugQ8mTFikelKsYYPqEUJqQUk3n+yc4B
vLKnI0GfDJ/CXagwf752X5Sv/HzZ1IrqRIc8dTrFH3HZHdBGi/QfSuedBx8RO8ADOlfzbc9y7Ge9
8ZEpVAX76ThHrxfNA4GfMNJdWuDzysGNslvGEKPqInrvPQIBdmeESORe+S/2T1dMyLfrY3lPh2ns
yo+w+zc8NrI0oY4ogXXqG6nYZFnwViTjMatwmglu6FtzfQImDT5zB0uA3mjFMb4HzGs7+NVPSlxK
GrIP8d64Iot/5ReAvulru1dOWKhywAooi6EkVKrkda/DuAHGLuMNaiISEpEJYc/+KXxFpdq2frUq
LuMCyeuAphsPLTWicIkArc58q1z3VfdWh8EGuQq6dSAWOyXyx9SsBJp6VR7mgFP5spVdYX3yUuuH
gj2GlhdF4jHvh8wkujvfnREHPOQqZea6cUhmZgDQoABP72kRKEEwGRi9gGG9G18uwU4DCrFeMEvY
BSYChPXf7zVBvZIKaFCcxhpkE3C2JO2fnJBL+5KhMPNFINQuwvRo9z+KxZZlt+Dv77lhKbMV1iNS
NZgs90pMp0s4GgOI1jo7kx7WKa5QNrz3P9Zu/3qEW1K4z4hlB/UZgQ9G5gWc2H9AoM59shvhg3QK
NpDRfDuyj+pn3h2UfVWVqNFlBeJLIW4oib+5MAFVOSbCN0PMTdmaLJMePe4nNaqzF23rA9/iumYj
7UzWx7HZBYfz5WbPMN3PIEdr3/Fklc1JgKAvlCmScFMjywLD9amq7Coidd2qnP+5DXR1MejaqlsS
JXZUXIbC0mYCBRiRo7lLSwvWHYSS3idBE3VZOk94YdSMl/dL6mPwkH7o0oyPTaZ5k7F+93MZYWxm
1BWaotL6/eNY69cCzbGQQeQ+lf7buBz7tguTxfAGIiUm+70bYlHQuLl311wzZYE+xrg3+zZxNprK
iEU2/+FxzICusBmO99f39HT6TYlygrWlBjKkgT5b5/Ir29/WvMaJbL9V0zlacHMdUflLHqFO2s8+
LhU2tiWfwET4idfIV2esS9BS0l37pGNrVgR97WT6rQWeGDqg1DTk5eikfRzJwRCBvvDPlzCmKiO8
KDUMVThKRlLmDH3pPxJC8b61/StjYyVsdhLwu180eL7z31UW+H4kRK1LmgZIXinjdY/wvAKIXv2/
AfFH6N3KfvTq+ux+HjUH6u/JrS+SlMkPw+BEk86RqXefnOd0tb4BQx1j/AHHcGSu1pvgmTo7ilfl
qhfRzPZ2CyRW1ikAiqpPzMBt7Hv/rZQjSzhYqOmIYj64n20BqYhJFBzGPVr2Et9pgXFw5PkhCCEu
4ZPb468cuQ27bF2bx9IJ+YDvnIDTSCZs3DyYPOQ5ABGZUEZ2d2wbLiR21yD+VuczI1jp3ZIakvzR
Pl7fhJDUrUnHYfxh5P4M1IDT+Zh67hmk9j6p9o36l5AC4iDNGYFpVD40sVce9FBG33q7t+seYV1S
ZZBz7epf1f6pgghDlP0G0rbD/4fXtiUMt444hE2RG6cadeSX3SkrgOPW8keGBD5L96MbwznAN2p4
xA3H1yf1U/r7FuDvVwUN/7Nv8enUTXCEA+UBxoQXlg9R4e8zyPOZ7vbKADX1AOSQsl/uMYWoSYjn
bU9m1LV3orv5I5OmEJhM0E/YMdAbnGGaA2mFzdnj9473G39kD8HGO/0hei1evNhw4Q+N5aD5hSg6
S3oqCeQxgvqYzU6H7r73iC2lqpGdp226fOMVyHqwkCxKLig1TgWWSHPXcRp9QWdtf4uwQj2xcluy
eznbf9P71yJj6ljtgYArIvjOJCjaUCfADI8LaViHdvPYixPLZV7XSUv2doNRh5eNFhXPOCxLRZ75
Xmv73L7BqN+hgzn5NuJpNk/9X+c3D5Dgupxl8QXKCXqYjK/F2mt6Ove01yDSvG8pfY93rZ3PqTLA
M6M00raSwjzdrc67E5+ifNQns7dHjYyQ+ILGSHACfTL1djLKay+mkgNXvuG5XUBPMU8SqHY8Pulv
lvNuv7k4SzjwwneCVEUPTA/LBFN7g+4nGzJoyhzWtEIg3fT+lS2kFB2Y1pDwV/w6zrkeY/bvTQL1
bwAhc2B+EZrmAIzl0kALPohz+p7Sm18CS2nVh+GT7Ju6VsXhi2DmWJEzTU/o9slvzNW5Vx3QAfUF
UDhswyrKCvVSvP+FxFAsqLX1Bml9TR4HnTURqYbAJQpsbbXVjtKzxnu9Gfripp6DX8gYUQzPg2hK
L9oxEvEZzeXvhm1iORp+N1X8thmPnIU2v0thS4ltUVAQCKvnX0W55uD3yPhyG5qby9sC8d7+ZnMM
X/wBTf3lwzSHFXwlKF+CPt/snpZB73EGIqg6fLOikIcKS3GjAvKNSoarSKdDst5yN30pcXmaB+Xt
mZiB0X85RhmHKheaF7Cg1PIaI7ohqpNOMjzStS6lyqH7z7OFMaA/z2ZCIj8oq7kxlRn9Gt5Q9Gb9
CC4b5pIT1xPp7dRWBXGe+iQl1mTjMGmQ9LxcaCLqtuuKlGMjG5so8IGz081aiM7GbSezxUW6sB4V
MdjuUUV/2nkPP6qFVOmZ9KwIsIjBEtf5sfTgw71MGVAfdvjku0jTMQaEwUq9V2J4CILe/bTx3TY4
idSPMcYXmF8PnKLbye/Z87bA7RREuLhOgtvAOAgYGqCN1v4PjNfTC/IBjgIKsHCqz1orGOPnv0s7
dA7sq1kzLmhNeo3XPgs9w+unrAF9PiMIL6QvPYQBjXvN6oei7JDL5oek5Q1T6Z3CzEUHAgU9+BW9
psA7i66IR8sE47XVr4X1y1qWiLbbjdbu44NfoMq0XXerUjR+gafCjMpCuPvIv7fT4riFNgItxAE+
1Lq+JEo11zyVZ0o7CwemyF8g7OEVrphjMXC7js+SP1CCaNt9ICqRFkzBsUOaTjJ5Myl7xQahXGg/
PW2j1SkxklTSv7a2ue3kyAhXqHowmKX8Mm2oC3G5XV8QdMuV7yCVA9EttKUB+vHi9A05xOyLZoNf
gd2kjm9vUsIKAxrhhUgOTuOIKgQljbqsVtYs0FelPyjn8brjOHq+I8YrJ1mZkB4giqAwyh6hiD5t
2S9NiqQdNkAmBQF19OuFdIKTtYCmR42ZY9Wt/k8fZOmTkIc/mWucJH/Erp/suxL5kH6RNf9jjWVe
spvWJLjpnF21ugDiGFibB3ztC74HwDZ9aGY9L8HwXLO/lY2EDp8Hyx25yBmc+FwlLBFdZywlBbk8
qEYVLti7ptd7Xf3mN6gruIY5RYFWzj532GaEOexcmEyaSAh59bZigB/L9/pbrtx0J2T8jSZP3elU
eQaQ7mxlU0BghGHGedfc/FDPfovgX5MydkZS8P7Is7BocBaZmvzFEmn86OwVlVklYuw+lgy+hdGs
A2rMUHAFJt/Nr6UIOMvRjZ9uaixAVNCKUexUTlgcycIc40vBcwzXPBMSQT8TdWkNDVxVI/gF+UjG
e66eHIyk70E+CilzuEBmKmA7cHisWUuCMF/PDTXVwU55kpBG0pQOgqZP213aU9G2C0pWmFY4jsoo
EHCu9rLMy46Q7pd+BLzwqqLyOriGNV5Avc/8ZBPj3j4n6sOokLWBcnHtXX49nrIqTah4GPCCl5Rm
pTKEYEdrawNIBlXMBs9ZmAHzdfHuLQH70JUh0QEqbuohSJBlGeob/q1xZKwqSFP98gf7OM0s/xRn
PbuVx96woeVPqHmrkqqqzYf6n5Ew2NKNMLomJazDJJqIhR5ftUUJw4zbgb3YaTpwHqo02bLIcwDY
kQLTIyPTUDB37NigfzIJ6OvbcgCiWtPie6kB4Au4MGceSidKWrBUvXUleT050i/H+SX2ulNdiSaj
l4gu8ljwl0lJAQE60Q+qjVzvbCoYlO8ZtkIrhBILTMM37ZPgT4OL7XQAvkMoEXTsrZJQ0JzmocrA
5tNlxfK6to/fbK5D2nSgpg7PqNLcBU13NJD9bI9jpX9jLCn9bzcT+EBbGPRw3EfJUxREFTaoqs2s
PJpCKcuwrohGMHNPqjGSRir+ys0Hvm1L92wJ/f6kuHO3UFuB6AYDObTeeYanBrnI4VpxRTlDNIlr
Vul2wm4xENqy2bDwZPoFehW6+FyizmL8g3Bgrs5mlA6CggFmnPilrSetf3pF6yVc8HIsjtJmp45/
ic/t1DGKi0XpAYo6UJlFyP+EYyUfj0SL72EMM0GXqDP9J+gHIG4BgbdObxTOV3BdjtxhEalPDaRE
Qj0Il5ARXztLelHW1mQdb7dVeJ0VNhyY9qzNIaPB1OoKuOgUFTotk/5EIO8gyOXOyj2bqZ0fUJjO
Q8EU6Ax5P79VK4OBdPe5t4wLTEDyZvQE0rTKbn2VnYuUuLly7LDv6u+70zdhqSwaso+S+bRi/0JM
0mmcp048teZfd6/HcucIKlgSVtNynT+Dl8RnedZ+4BUUIoxwqJmWHIjL/557MPDZExm493fUWbMY
DEk5XKSPyHtYpaf40aLUu7CNMAWsul0JMb7pXtMbP04twAcbutTKYmKWFi8w0jjeh8MRs6Svla+S
evXFGgrC42D6c5XCCNvHMyy/hJ1f+jWPX1xK0C7Jf/K8qqDx6oysNhWLzsREmLBowlRBpKAKFrWl
RDmfp3zpCV2d7FlfGEpkNR57Fci7hgzuO+3EHaWXGT19KPl3nm6AbnHbJ8LFdgsv4tLYb+Wv3abY
HGDucH83nFvnk1gfbnIvIvHrSCt4sKSKIuFacohSPjOSM5nrUN++cVEcZAox3tNOhMOFPwYbLDGv
3lWakLESpksQji/Nk1JHWJV77MzFOgSCSCmvc1WGEADjGRfjnPeoXsm9luEh8Hln6jrFaMlfd6cs
PuenavUKVk6qNu+qNlpselPbRHyv79Ky9GiG2mc2FUD0s7u83GCiJByUwBr6DV5UqSO9+5yn0LmV
9ZqiFzuwSxSE3omaZYV79SMd48+xwGEumdIG6voIpc6txtydBYlUVKUqVTUnXI30u8c4ZGkDDxWt
zTw+1lCmNoMEdtDejJYZZFALMcLWh61jsnQm4bhKUcAad7o0xB6XzlDZE3VDKnFcrBgAbrlB/8OV
khDsf8zka3Mi1WIfMFWSZVAvO+f4PiTtmJa4RQU9Jn6rX3ivzl04uz9HZNiBKpgRoxn51visyn8S
FTKweEfQT+yK9hWf/Eh8FLhKL6dKMM6UCme60Di7Ykvhxk7dvsQQ6EoBOCDCEyAb8NZm558kBW7P
2qXiHVmwNgGK3jYi9tHr
`protect end_protected

