

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SQUyeNX8cyskpzvvW2T3ssUGj6xZX5vHX5fJU9Ms0M+rWpNjMO6za6Zgr1K2FMwHi+buwP0Gw29j
IKEYpdzZOw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hoBaDPgZL0nmY18FE8yzpnxIEfx7SKisNM4FVo3Ao91EGtVywU0Wb7yA1enrW6Xd+oLWYcrMdoDX
JTxy8JdlM3o+jyjU7UKGIkB+vX642Q6fBAuo3SZKPKM/RE7lQknQIOi2Y5V60nbw/AM6mvYDKdTS
wiPRLcQIZpvU4dn9GkQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o9OFQKQt0GaB68TjFqZyGwbFj1TRgCs2FzlOtaWTgxoDRMFT9IEssmRwHo9pwJ5Tn3OigUlzbBbd
XTy7vthduMEKESguEgGeFDAlZPJdvm6/cpwtG3omF99Y9vBxA2K/3YI0+jDh2eyUvsHMcDbQ/C2p
zFKW1hcipARgm3A9Ys4mkgzXMVKYnvnQiSsmezjrXPsPy8jbFYPXFd6vFSGi/ZwrKMMLLNZt/Boe
k/Pl01HBEt/KNoY9VFx6N+e2ufES+vAz0H+DJSGPch6YdjmhkZUj2llujVX2dT6EzXeB2X9+1Sar
qYaNJFQdqXN7nDqoQMCiwqUZBJaHNrPJdzAMcw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gMFEdGC+ckR/NJmX/aszkYoB651qUCnYvXxq63Zrpc98jREIyboMJaogrhiyZ1kntx31alD51ug4
ZAed1vud+wZB4IN9oJ1STjbhb+Zj5u4I029j7Gy2lllPl+1O8Em+DnBFlaNak9VTW5oxld5AFJs/
EstFEKIMT8MSbegVIEQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I2MWBDnGcReW7SMjRXdvt63Rjoo/gu+NQcstRp+eRPxV1cdY3BaChhCXefqNXs4HwrSwjy6eXoRH
K9pkdKW/MmeSQuCCGBXm3SZnri7VuXOoNwZoR7yYcuzRHYCe4OVzWrXYc7CJVdShI1TzYNVzTc69
N+748OjVGLm080Ri6+7tnRVNASpwPZfo8iBz5hClukZRieQCUQgdHIAZx2RjUyVQaoW7cJ/urtOZ
zr2GA2iDsweYcuo/xtEmVehzY9Jjyk+XsH/W+/8SFJEIN/wAiWoW84/gDLItkUU21xaixyhQCl/Y
sHoICo/iHc8aTOV1SPHo9yWYmV0UZ8KJqveuUA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`protect data_block
mhGvRHZ8hz1uDeYOwGYU5qJ0V7dbXIjRP+cda8YydV4jqgPbfK1KbSjWOXb6JYTNT+BAKHH6gSw6
M62t3AU98aegCmUKStO7Nf0w4P92gpq1mrS3SYlgsZ5aT3jPDDZZiT5ZL2Wo2C0IsKiLHuBw41TZ
+uZVDEApiDzV6b5WYz84kENiEAfvQKK+eUeZBZ+Khq2nO9kDH0fzDcQUbWVmjakqD3MopadsYXxJ
GEDJFw9RLl4AzHu3kTEPObld2idmRm4oLS8GUBsYz0Mtiyqi23XKt7uuOrZZmtfXFhBXSLS/o/sM
PguxFGTDBpE15IQ7UkJoGnQMsDK3PxugPoZpvvQ+QiY+G56OsDnXT23v+g0nJ7dDkkanD8mHanI8
YELS4WFEGtroZ3VIjKSkMitNtKkymOL+hbfoHTP0P+C1EWrynhyZ/0HxnxgX0y1ycjepGDMaW+cQ
aB1f70O3oBfUPMxAJYx9vLxAsuWx5PEQhrmC8gHLRIgyTZsYka8vUdhQLlj2bCgmbT0gbA0FqkF4
m7Vyax+r00v4X8LRheZM5SqcqauORdfDGOzdlIFsGsqyAL5MfxrZYft/zAPxCeDZzxhQkcUZP/AT
EHMbF2xbFNF1Ayaei4+o7Mh1AsPsLBRRuoQwLuJ2SC2OgCVKXHHfUgb135GiNMHu509LO2bTjEnk
ro1HOvyTIa6YwfjFqF0uYfcODotigS+dpE0I59+6ZNctdq2I9hBvJfBo0yQ3YQTu7FI4VoRIjsy7
dd1x4moRBn7YoWZJ248OX5dM7vbsZggDRtklkozWIjCpcq8XAB410T0TqFmyCRk6JkPJg6brL0d2
75vzS5vN59Pg8dzEDSoKS1GpokWfEmYCpmAii39cSSgQ+wnW24JMnUfd16dMBKAoVeZ6qtYvHsug
WluJkxr5lKjSJoCUBoUd7TkUlJXelEsDS9L19Xuau9RCidmuRhVCUGAmRIinT9VBqxyL+pv95uKF
7H/TmcuD00ILTs2wYdZLSuTHh/X4d7rTIsZLlU23Vs3MqD+rxXLGEcVYf93ZUriwQaLMAKoujCFP
gcJXKRoVQSdDxYUV/nOJKQPmtFBAM9S7bIh9cXe6G7yYlBfZHCK2wPnb79pQN39WV3hsSt7bEf4I
BYob2yoekoOq4Y0sNCApA3YPvM8nH0hyFZcjkpf9HjnMIDh4FVOKM6GMsgHEBGo7hl/uaVD+gGXF
N4sSPGegjihwCbmp0h/gAjHu0JvAp/ee4ILUp7zmnlTpZwY+8nBRHM4xSnkiISpFkEVrRI9O11Vl
rz8mpV4vtgIg4fZVLbw4YMGs0MGbN/dI/2cfupjAdcjxWlR7HSHZ0O76M5qnJCJwvfaJv/TkComK
59GOxAEf1mqbI+K/FhamGJYGDMBmJ/ue7F/YrCGcYBPYO1RRAdG3OdTkjGhmQbsibazh5qSSTNg2
E+isvu0oczZD6OtLfmTM5PxIUhSIma+msvCFuPCZuK+U6R0jy75Xq4dVli80YbJzdiXdxPRaXh1y
0n/6Fy25dz8FK1lJhNLMdqhqVfeD08kNfoJn58usvOw9zNNRhqW9MlrpiPKZa2JEbbkgvgTcK7mK
wYq+qexBCAaXUJCldKmi3hGLKT50eYNSpFiGTMVQRnvXJaZgjDfduID9zB9As9bhLgt/L+uUcqPH
V7hQ3N190+NPLxp21Y+CKS+gx+V7iQktyJi6X36TsU3MdfVmO1TmEXDMnvAXcZoF5zHhKJ3bquKT
/tD9uBNQ1btPFJ6Z3F8AHK3Hv9rXECKSKSzYRzSkxIVDRAoji/gAzEwt+th757VGd40/K9P8On22
rlIrYORIgiYo7srsCKdKP9u5cW1163pWfJNQtQqSRglZpNM8BgoyT4e+iGJ5ZxcsaHNRVZjq6/o9
zxadfOKxDy05jrb09B4M69LGVUbciHD/jz9kgWhiSsWNsjAw6XYXP2Bz/LUV+GG+R+VedvXF3Cnx
9S3qH56fgG8jYQm7b9dBmKjVYWYw6X0wJIHDvvv7Runs/Wv6d42USczEew6rmeDhjCMtjqBN9tXU
W/tRu/Nu3m7sjSySoWnQVX9ypDqMql2S+nWBwZ50fVxUvp92K3mZyCRiujTesZHoDgA3NQHSEWNk
ZiZGnbAjVJrJwZtLqdlrJ4PUY4TioNYJygfZ1bFvswMO6b8LuF73sKou1YRKwA3X8LoIQRwWADrB
rtm+wRk0bSIK2jqvPTHb0DQw78QWaVXt6ZsT/raxVa2TcbdeeophmaY2mc/jV94SE/Hs/npGHAfE
d8uYWlNAArQzpA21nsaOGb84v+h39FBy585cc6M3KYtPEshtGJKcVx0Sx+V0tD9E8fP9e+GpgnFs
CkLiWJTnMJW6i63Y394ZzbteRwkMJiZUcLuKCbZ+KZgzQAhbvyaqa3nbTXwanmaORsWxs5jhXu9n
ELh4qcVyLMCtokJwGC97JxRGrFCaj3o0VlFxRJZANxnUCau/qNmq7+AwUrMee5Bd1V49oZnddljg
pVSN2nyPACTtOLH3skAuL6Wg7HmajEnzYGqpLi2B0pYUWEpxvlEiSIe7TvK5FQgH0iyEzQdTy90r
Niq2MC/f9U40hbhrdFGHZ/V2jnZ6zQYGQMTSXcGXWgc5WeD9YS6dJGKFmzWq2gPlFQe9CpYjg7dx
aeelLa5sJwOQ49UfnzizsGubic2ig57/9FSMsAYVgnRsbOB+yGczqz+tDbYvT3w2+CruzkN0O54G
cyKn8Qxnohz7ZbCkDtbIL43YJr6iEEJ6XVzOr5VJ2zaSdWUNo5HmAyAw25gG7msW1mZP+If2PWvQ
Eg85PUKsQvshZm3dDWX27xIyrSP/OjBHLm+8pwn5OlraqjyH3CytgXkzdPj1ZpXdvAhI9Zfx05S0
jcdyKOUI0JGffMEEu+fs/WA2Bg4sMf8ueRkLsF9hag9bstzsefLEmwwWg4LoGQEzVgi+UHopn1/a
AJOScZl9wsXQEkrAnwY1V0whcaCblQQ8wTf7F9VdEVXzrlNWrifapX2luPXcw9jtMCyxDxLf8hrG
ZrF7YaYzi4tFpfFzMgvV9jbkgiTpJMiag0k6wVcSKKzrHPQLZT1fsqYzjwaBNjia6OSe+gvCyUOo
okc5JHsi88QPfW4gFWXF7/p5mQmhQ+cOl6KInb7I47dXJV6hwumQebzp6ETHNVpEF/CeLp9l/7AX
h/dnspj986Na+gx7nElc1gqE80R3b4HSpSZLWWA5tho2RQejWtfOSO9H2VVWOeCU5kMkxxL9FaJC
XHr+lhOgmPq1DWqhZ0aT8C2OfeTGa+E0W3SVkBtjlINmVMrzNY/jGOpOFbEQl3E/ckoebIoPhB76
SE1VW+qanitjKJx4ORUSyPXsvOelPD93kqy9vvjweuJm2XupQ/ydG8cJj80nsf6kmsUlYG4MLXRL
ky5geF713dEhOl37mZfWA1veoyveINGNnceF4b5Sd1kvQ283iOyLAKpi/OR6mQ1kZ7gqZha4y1VG
l2+LsUng7vEB6HrcszSi8I85+zsTTGgxfTSTrZGUir+bUqHS//O4zfQVrlD6fVq6l2IReau6hTaw
z7fNoRvV5BH7/5t3xiO960HSTZUGh+HNfAhpCLGWGTX/9WGNlYRkaQyNbCUs+/xdSsjzC11a5VsI
Kb0UB4yx3CrxJgVJrdVyEye10aWHGEXR1f3KF3FW/zoxVnbNGCfXWbi3O5wdlVBRPSlIadeLZ8Ct
YloyDOsFvGQqKhhlFDjUftaYx926huCEESTz4GVQxBCtW2ed4TpS35hCl5Xyq0a46ZDRLF2yB/pl
hKTcEBpa4GYfZGainPkW5N/RvLF7rqxVOCadCuHQyy+z1gYDCL2TYAsWpD/jFlFB2VJiir4qyKLw
x0VF/cZlEvNLXwGmJfbfbiUljYpEF576V+aI7/75yq6Jrltw9nvRIo2EKBFmnLPjNpuUwY3StDfY
rY4jzAZNB3QqpzBjkFJ2JHErU8CtUDxnEniEWLfiNKtzSjyJlveGNhZOoaySW8qAq3UQqgFjE0A5
KGW3cL/QdLRSV+MFyo3ppkCeQi0jJdz3iuzTYv6m358uX6zYXFn4AEUHqu53PT8HR2E4+R6qjl2W
UF4mBJli+j5Zs1bmlVp3Dp0c/wG1TRm9F0h8+hjgU1WaDDgskYecu7kmaJnFbQP/v06rFux9cZAI
rnkajRHqhX+4ew77hFssk+cLrHITR0CTlOFAidWul2bPl2+VFSydqES98rpZ99JiZJEnXczLQ4UI
FMAJ2236cHkfxGDsRZlOuahioAYvDlrIOquT0g2MeTBXVdRblPfPx7EfQGDCm5uigZidu6xukkpt
2wwbpCz/jtE7ghac3GQmibEK2clxJuS85qTUCWrSKUCL8xv6gjMjEb4qyWmawCuhXSwX+RhTUHtk
/cXAqfwWNSylLNRQfhrVPJpsY8GuvHNvD9FgyyDfXCS41kn7c4DjutI7Ma64ytzzT0zA53fClgHj
jbMyLjPvDGdHLZ3tZ26XP9dwz0q/1V+6lyTbhbKPI6z2/7anrNK0FmlRlTWR5gvMaEz+HKFY3f+m
K1sm+kwXe6LnmkQJonelBrhHfYKSWkdIYZ87P69AuxCcx+en5z7j1UmjAV66BFWFyZSivvwAO5kp
XILlpMHFxZGAg5wlgHC0Gk7MLtoYJhu3/CUgU3HPBYeW0XSGlrvoQBnbxAdmAxA74YatvhEsaiNe
4/mIlgw8IhYKDDAiSxK9hkAhWWXTAbbtCBD449AeQ/AmQ7hP/rRb6aRlX9iUsZA1/8+HMGNwgG/U
qxIhtWFOvlXtwmH8fVwrDKTfgD7v0PhwZxALHYp2m5GPzra9SiGrx/K2XzqBs9P5MfzK0tN5wFaR
6cORwFRImiEtxirT3G1aL0Wy3Ar8qiIbWLPDSjfa407SGk+ZiW+XJpebjC2OI/btbnrIo8zyVO2r
sLXHKKOUL0jnomtmTKpBi/bBzYBTnVNAGTJogL0zDiyy6FgGLuvLTSXTNR0bWk6F2g6wgUBSg1Gp
wFcamaUjJwi10AmHL7Hqy8St8ydZr97yHo2jMGr34FlOPDuDkCJfJx42cM75oaaGHUbqvRCtdBsq
8+6WUC/LF36n42Qr3qpTzO4xYDVNZaCqBJOGrFiYBSiEpeJMe7OtCFCFfvWRgVjDEwVZQ++QDvHv
20arb++Gj5W1lU1gxsmSQjHTCuqXNfONkSzGcRBPOXHdaj/85vwKnIWCOwgspI/DZGPjGd5nh/eF
4o2j6V4W5Ij9tI3vSkDRIz1akS4SPklzXe4jCHzv/IWOIuHZbLb2CpVk2tJpyv50w2HupNNWL72/
yEUWYTZsA+Dan1gGV58YEftL1jtQFqSCmZnU411MywfSOufl2Y7JjyT8L6tJS3Mk4qQnYVLEKDpt
sZJzzcF8X73gHWmynmKIcM9qbmoDEIC85VmlVjvaXnX/CA+SXgTB/lKvWMT9d8djN2LzcdalpdP1
luHCsCw20T7iWQ86nSUF9Qz88cI2MmhIOax1Pyj/+1vlqmzb3jIOu7FA6zjemN97dpUgA7PwmC6h
PtF9KWmKw9kHlv4Fc+D49I4wmd/hiImxGQcpsf7bbW33iv1rBke6Wn4BKpRIS3gKQRWdAVDFTaaI
JEneH1h/BfRnWd5IQPnezdqMlrtNBmTro+11sCUBbc4NN7bFoJ+Rvfe/pA9TvSDttAfrScxn7Q9F
jFEa5OFSrDtu8czFEH6M7nMh2MEVwp+Zm5Sg/w2Nbe/6rHLWI8W6+z9IJNLJezuO5JWL+YpE7Hnm
/LrtJMFiHO0dpECSgkz0ZJQBE6ty0jlkgtFVVlbtguhdbrvkuw+mASbubsfpklKdJcD/O00CnOwx
KkVecKy+Rg8W5KCVKJcghYqP3r/QcCXIiNs1h9wrIVSIqsSWsW9Sf8V/wwMsQnkXg025Ef3lzhg9
Jwt8amjUKAOOf6q2/hPtaqbkdtmim1j35bB66ffwWNbFhSPhspnRjco/lxqOYJU6qH+Er35LR/OI
4eo7w+XGftYFxWqi3+PKkZYFAbdkf8mmr+BjmNyxi8IfaViW24eGEL60vrCmsdWZeYCx4wnqkYCW
v4bchqXkW+qkpTiqoiHwoPu3/UABWCZiObY1jobyb0BAHJewBQ3GyOEgYeXJVNNzKRxIKYecel73
OF+PiATtcQWchsLN9bKVw5pjTpST7O4Zptl35m6H+CAz1N4SWLgTH922WNzkI66k1z6AJ9tg6q21
Iq+YxynxbI1ANbUmmmZ9InZ5bO9vfq4EPI0wS7ESA8KaIbcOl2R8KCAWAncvCJJRWl5ZqoF/5au2
39KoyH4IaTvTbi3EmzQFfFcmKlIEJlSTpb5psGmY5HD1BPmmLwqEmsQQqkzs27NrnYS/F+z2fqL6
QJUD7QVpt8l6EBPTx9VVQfh4pAdr2xL7cfLz0VyP6b47HCiXp5u/R2TA319/wtv++I2cCAfMdNvX
+o5eDt4pO68alDzp2D6Y+DPX1+znziGHBzkKIoPHsdJTsYul3GRKQUo/dG2sIS5WQQQUlWuqhqCh
J8SqPTmmIZCMTXuPJI6ei5S5vmIC2U/1sZ+1q6Js+XwUrN9aMPNQOa3OxvsVNICj9i6X/nxGkAYD
h75kbRNsYESEJMXi4eFHThhDQSaZbVugEqJQCmUlwNhEoSKr26otWQyqkpB0mtXrUc+E8hBN9T5o
0pUATk9dBAxL/PTueZkLA+/IE34XjfLwO6kqETbryaHC7/YqbxblWPm4Hax4SiChFFz+R46V0q/i
xwObV561apIcVFHCcMrf26Nuhn+1dWZ41DqhLdqQzwqV6os3N7y4G9Z7KMtfQ3YKnDNcyGjn6HjR
ZM86nXkFBGJygkh8yvwe9SygMlvMhYTBpzY2uIFAXAwTtE/rA7n3Dljw+T0NBx38QFoaDfnNqXsE
XaduLN4wGJwHKF6g6yxkRKQIlcVJhtJSOsc9sN3pq1ah+qKIpqUFwSsCKHZYsVEfiAxTvVzyaMvl
xcZLm8NDjgGlUNm3/uWlJmpHSSSlkuw2tQCznaOnHgfsRE4eiGmfGbWin7v8CA28RU/zQX0/eOUm
1YXh0dQdj2ESwJX439bOPLfXAS+5C0fs4Qj+4JkwfeGlPykNjYx1bvWTT/Gfaut2O/B61Pq5dV0r
/DeFNVHmYAyT9Q7rltsfK7Eiqze/QPV1SRRbsMQn0ogxXgG6LvO9Qzy6LWAnR/b8BCGc4SPUMWBT
B8exoKC81yVSSTPNqqudE/eM1geOu0ivpB2nv+OosUoGCpEfNNn9SmUeQQ7g7pzE+6X9BBI5QbJZ
UELMG+UCT83W84hYYvl/xJ829M6nFZDl8JfUkUEVHFGHR1qBzZUM8SOt17WoHCvo2TEMuLj+uW0Q
7NiKx5C8xu0Pj40BOAd/nZ0QmO6lfoSUmrQPFe5LtxKypLp3SdPd9tAlVadjKgaQsuz1oxmnLPmb
jwjW3xAcIc+YB1Al4ndOimhf1MHpA94SVAYrxzBcjmq0XEovafl6odxh1yhxvM5ST3T+NOli4Jox
gkrtVVsckrS0UqLHAlf6jNGSn8RHc0Yjg50C2tzNC7b9szUScDDSkdg63SS83TX2l3MG6LXb3UDB
Kc6b+CHcUbnEMR93IKIIK+LyERAKeZwAZhYLysn2izdYWwbPTPldjpLoVRuvSHClzXUTdoB9bRxq
Kd6VyUbi4ipcDg3eom1hP3DDifDu0D9A+VSjOuSufjlAb97mVOeHLrJaqq9gE6a0Ud/JBXWFcNMy
/6M1qDAnH7KaVcUVFmryI4TAS1B4hhhSQjb88rkazuzpTEfpO9RKy4JEUnDGlhBCde5G7XRKOIVa
JJ/87fSmSY/IdS1puT7PaGXEgb9u7anSypNINSKreDOvCD//+XSKVEfSFWIZpVuxrSVYt5tRL8Ca
Z4hWUDL5VIZ4zDB5MpsoYcAODryE6BeR6HLr5lksAitlr0fdSvPReZeKFb6e5njNMAXL/xuZe5Sd
ajyiMKvmRmxMuBrmZWo4KIl9d87ImL7coOpaFJ92g7f2tZhLOZD4ia2mPTczJqtF/Npm+tFjI8Wo
Ljfmy2waCf6fQ5EE5wsjpVkZo5U41mGYLpcr8VOgYlNg27Gcvd0Jidw2A7czvK1sU0EUaCoDxEWT
JU2dpi7qbUPNyoQ7yy+6NC3AahqW25McFVpAsstNzlOj6Kg4cMWts32obji9NYBGqKsgwDW+TKTL
zOxNd4MYfs8eUKmUR/cqeUzxTjdx+UZUP9XioXfwu9LHLe7DNGrue5LG0AkJOVXGzDaA9oQG08uR
WwEjefuXVFgbdB1FDgsxEIwGRp+TFxNi5LJW3tzOz0ti/o/UzxhToqwFbePxDxDBGNV8Hh0ZUD9C
/2y6Xei9uuaGTYq/WukXusGWVH7nQ1vhs3+zCi4YvpCwvQ==
`protect end_protected

