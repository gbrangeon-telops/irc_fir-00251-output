

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
US2mB3ZU2xYMwSgf2KG3QONmAU5qxOR5gFmXyP3MzegSXblZ76jq0dw3DGi2XivflSREvQG+tGNr
93kJJN9RHg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cVCcDe3dO8A3aQlcacvtDrMlOeMM3iFulWP1GnL0AstVpxpdCCRRxU3UHiCxbevv+1Dnaf6o7WxT
G4MiJBrZR0NZpyZrN6elCTa1aex/x1et3mJ/kXtaSnXZDYRGWgFlsFwFLktb6kdkyrjtbx1rPCM3
CfbtCvTObEIGzIf/FJI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ybpmXaWiA2h4ouUhToF83n5FZ6mSwY7i2SbAGhh214jlEV4EAw60pDdsC9S1DXRUJs2H5ijqRHjq
O6r3TnjNUgOULu96coukm/eTQWKkKJe9Aqdi1COsXCRXpY/qPst8iFpcYgvP7x9BLqj2FuOVCOp1
vBc1X163t+3g+Wnu5wdB02cYtsPg85Aym4KDvpdGC2+lcbTElJIi+JurCHNEVSPxn/s/byKj9Aee
BWqSso/XFdRP+TM7huy2D0efcTINLjUE/2qeG1Z2VdFBpyOvUXxDlOhNEr+qAiw/pCiqNyrHCapM
TfSbH498t2P5uuhd9n2zpj2CUOFq13OvODvHsg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o4nr3qLm7Rem+yVuZpGX2Dwzye61TgXXpiZsrYTQhxAIOttLQ5qy48oMqssSkd1Afuq4E1AgeeLD
pr9heGHoD5AjWxk13hv9r2YUI3BND7NaVLyrx7mIkF/pxjMjFTBF3rI5FZuYgxY00aftrEFjG/AI
XeOeb4w/KZQIUde+tJY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dHlANyrutuNgAtytsZMPMatpxiEBkM3u/gDZ64fIbSRqU16FBJ0WguNKCot1/TeXAq8CSJHQCt8x
3wxDlxfMsEEJdw5OF5Pn172rV07Ce6wZ30zB83ou1uUKjnNgy6pYqTworLe5Tj4SYl9VY0bcZ0g/
rN0niMih/6g+8XwbbPNRS7in3icwjpeqxdXwsRyEX3dbCrKVz4LXcfmP+ybNfKunFSp+imrzoFLt
cLJF8o/HdEoH/59p1whEdIyNin1+Ra+5d2hGnILLEgUP28LNS8Xr0dqjxGFNrkIDmtSmsmF2E1fl
JbLYu0fIIENjFn9nAJCzGQU523347ABwMPcyhA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5328)
`protect data_block
Ji7CJgCMFWKuXoWoNNUrpOQhxiVNaNDAAvdIArBZJdm49UqgV4J13YnY4RGQlu+m30gLcNzOeqdq
mA+6scyeiGHfmrmUWOZU+eow2QmiizNAZWWe2mOZJ880wiDOG6pu7G8pC2LV58rSiw4V2qEs4B+2
fSc4F7VuVtum1GBi+zw7Yq4qNw4/tJ8w3OPjb2PioHQv5IXbmvWegaurSxGLixT52Ic9wbMoSLPB
i5p5AHEBiMUkgl3tnzUFrhVbWemQyEzu+1ZL0lqv2zaiDrLXptK5lXrPdx/cP5fVp4Xawm8xSIl3
3bfzbT7OJMJZaFqeiKdYXx+ohexXSUlFZH0H3fI9BkwXHTE9rGwrokNjDw2EHjapEAyFjgoHOiBd
nRlAXOUD1vQlsRFCUEs0zQoYpNYgB10780ovXGwcWL9M6000H9mBTFxS7HXTec7fizStfY/qCZ3Z
hfcpzKhlP2393LFWBxpqEyaWTMvA+F4ybdLl0h8M/DLZVUEha7ZpYOX9MTlgpu5SWwjp4bDBO13T
fhT0xCmCsLGWudxiWXP/Jj6z7GNMOHbv4NtUYfjyOdh3O1jNadVsfUjPasQaF+SFVzf4QWbKUzS3
cNJlgQRCVdSCB0x+FIJURuiGTtxIj3+yjUfUdYCxe1xHy5ro8m/PPJEKfOn+2iTGO9MTZI4xexf/
eoUm7Ngn85FKToEgKac+zhzssK2GH2JPUEfFrnkD/gOAPhPq9H3XqCzTZ15oOXpaKIHfjBA/kdJs
VBHbHgn2O5oZkNAKxiuhSaVNcf22piGbTmlRYp5LyL462IfzmJpi8pXAoeidoTUneVUAkx5/6RAm
xXFpu5Is52dW1zQtEwphw89AaeOclx001p/A6cq2kZ+yBaalQbfKd84cupneqIDiTA71O99ZWMxM
UFfSQ6d4/MQWA7XN9u7O17dC0ZZ98FemOv8D2fxS60Ty8uw77JK0A4p+VG3LbEqlMTISXWjEdlMO
tF/gAWZgtPQtPGEjhK3h5WhnHAyVZfI7Qex9yW6J3scGrr+/CtgH+nQaYudFO5JxagcT8WvGPe85
8IHVVwbi1cLTYcx/UctMS1O3pxWoBkSGVCNa16pEjDHypV+VGmf8IONEkuRQL+EbCcA1t2EXlIEg
ppycrIBtctSdBCTW/tbmIv1cDWLESyUezVRTJRO8WqkX/2ltsI/OwFWYmG1HHyaShYCdvgiePj+v
xJbKzrMQs7dBzDedfaa7rq7uHBuTcxRyaNeyzziTH6zMVPAhsWPT2qBE4VL180KuT9xAJc2Izt8C
XoUgVQEdCT4uDHhiejQ1gvODPy52+gJWU04HojlWF7brGl8VKqW4FBsAc2wwXQCkew+1XEjq8W0X
2ybINLuT/BduxrY/cxli2lDhO3hAaUriotJDGdlsxHi+ydPICXM0qUSsSeeZf4vGSY9xuKTjjnaM
84tel+DP7QjXpuM/9jR1ht458btbO5vEUMqSfVFjssD9Y++1y60ntvFgyW4UjuR74ecBWnSVH4yH
uYRnHm1llRWqWSRJ8s11poCqXfe5Bb7cfvrBj7FPWHCOzR+4TxaSOeCaP0gRgi0Jl1p0s3CK+IZC
Mq+wXy13PjMxvpyouBmo9ZyCjZwllcU5S8SKS9ib+XEsa5Kuq6srgz739nja9FFUaTwyDK0jRK8q
pW8k1lLioo9OFvdSWYavi2PjSNnXBuAYe1dpHgYyByTa5P18F8vhn5zIkQLE3WGk9VvizKKr0UlE
Yo5KYLI3HJ+KkvVBzaawDm9/FrNVLF0dOoeb/eOc6T/WsPgtPogIUbmKqxuV1AOprd8uYxuFyXHS
y+JJMNyNYCJdTdKlE01DyxCa6Po/4jy53cKsh7wXFHutZ0n6/XjErRe9bXs/gVgAx9sXV/8BECtc
6cGC9pEJaFza+HLCEKJggKlis2WZeWtbzvjjSIMTz562abzD0jHEpO47ff954O4ynIcye1narxdD
f/srtbK6HZ9NmaluKODIGYdSzkVtvx2xxCQLcS4U9x5b6mohK0ZRbg4OLihcc3lFWXj9kTcJ962H
uwm5e2apCbP1l2xJ3O8B4Bl85G3Y9gr0ZlmhRfgwql6K5/r5RpbrN3jp5cdEFyApkrnTquNibEQx
4+8pa2UAmjLEd4J/81gPFbef3gqyvnfAsBceb3q0EHSjh4K1dSOlt+TWUU/Rbj6EbUYy2a/Dyb0b
bOzKFwB+NyUBG2cpQLpCKWXZweJK8Q1yYFuE0kWBhsEinWmxrBo8A2lABpfDYxWCBoouYLcDqU3H
m6wT1AoFumagzj8DQJheTthRPnQGDtH+dnby1rWK643iaZCSL8HlH/MGoEwImxEfU4WCri0mivYI
envN2h2IO63kSyMJ9/c9Iw+iUEbQ73fe7b2TA/SfsLx3LBrBnKuoEv/R1j2OqDkcD0dNlTMuGVIw
8dpbZWKvyobwJyGJdSWPdNVD+C1pPsv8h77ed4NeHw0u2cXBuKkXZp3f6NrVKPJdA79i/xpbgXaf
DZUme4NspYmJj0BDx8wnc1J8upeZ6QKpC7NKv2UshEsWJ1ogTy96+FEEVPPet5QJu3I+AH+apegS
iq3vbJoUfUoqyeo/aGtPOzn78SynJ1fVkbZK9OdFolbWNindjqtWdp0sgDPlCky8utEmI0cRngKx
+KfFrZhLpBQDxN7Zz7GXKmZnxyhT9WGr7j2uzBoTYkqd/iQJQnDjEdk44cYLNRLpiJ404v8t4co2
TgvWCX7eGcDSBVoOdK9SWgXuxaDkXg7eCSsrVgQ3Y5ACARimA/TQ9MAiJN6rEZrPyQ4cHJ14sxAr
bwE2nrgjkogk0KBLCPDVOeuys52RI1Tl6aKfKl8CA9/GPqGdUBkP3nXW8SQnDUcOajL/8BfbM96g
LLgtNRHA0TZjaTJxUSh+ntRQEhg9iyLdW+Wrh0mCdNlDmqxy4t4IvGs48JkLsj3J65GTdfC3h9Tf
x1iauwUmLBGXAIk0k267BMMGVfsFeRRTqrdntU/tIQfm5PAfgYBnk9Q5DLGDcu9K91ALky7k2Cwn
eWmyFID1mERPvTcOBtp5A+GvaWh31TxzWlWyrjRCF0oI0B7BkiW6+AqjBrx4NF5VXH1gcrj3R42Q
2eUkgJ9LL+2A5Loi+VYCFkukfgjXyBMgXn1l9OknkCW9sQyuK/6CK9laBVrgiyAEFG3TVSL1gNiD
bj7NhBAHmBlOBtujDt5n+GJTq0QAn9O4jmxHWLk7XC/j3/odRLvRxErgaCezPw2BjDhYN131Q6ye
37Ac0yMxgYc5FPIBgSRiEcgHDsoU/0J6Hx0mL0jCZ6NTfW0XQiVw/MPENd3n4Rm6EEAAb08pgBpp
4QZua92HCP+Ri2vpK1FPHoG6BfvRhIXYij99WUtcqYCrqDCc3/b2KDPBYHCLVVU5jgE12BXOU+NH
23twZA4xu+Nb0z31/GJQpXT/oRqFFy2CenwaEYFHGdiqxtKa5OY+yzJ2vm1lJ/RRYm75vOAZto1E
jeMV4xaKzTwSdBLI3UvfReMQglPHw3Qj7Z5MFkuHoOCITn9OmAeXdLQIqDKt+D3EIv9OA5NRBWy0
5mR3nERnznOCeoQN63B2LWPFbC8C0z0bPq2JAUrzVX+Ar+SkcOs/JLOKL2MZjcBud7RZIDhwaIM0
wJAwTdZpklFsyXc63xkungUnUt/LDxqnAzx8wCpxIOVPeylqnPJjX43ckTqAImLQ6XOZUbzmhums
ueN9wHMFvZuYbkaHMBOcFu9ZA/KSQE/UVBkZ7Y77qxiKH3QFBsdAaknQ+Gjuw/2Ml0dQVT3oAVt+
XXX8U7U2HWR2TbjQrUAoCfzuSQtUTH+qNSiC9MFV09mhiIQjoNKcmG8N+fHxVHdwrgSs+fBL4J4i
qAA6RirDD/mWWx+Adc1RtA7EGq4zPVNMU0TqqJgTubyiD4MZaHn0AiAyF5rodv5nfboDhLXFtx0u
FVvC9uEjp2kSUXB3X3S5ycPaSEtLzDadkKDsSHulqqMCIbiB/ChLbssgZCo/0y4X1WMY19roB7RL
R25UKS/d91mJ8GFaVemskw1wBSSk03pIEGS/qugSHfYud4bjY7rXu8b589oHl4IdUtk1aiNDW7u/
rp9wY2zzV/VgpoFQeeUuv4a7yfpP/FJtOayzapnxfdaXb620ICCI5374SiS9P+tSvV28cSzmGYAs
Cj/RJMU7LYp5q5d4g9j18gITLHGZP5FI1vO3fGFhZvqY1fpB7kayiUPDwdjEdk6lH8MgnOenHuH1
5Ma488qD82pbSCm0d4SbsgqJFcLVrxaVW1sA3rSCd8gMSzsDH6fF4fpkV4GIuvUOwlBgklWagTUm
S2wEhXWk89Rc1vBnQvzW/8rF6OtwGDNEsEgTZTPHuuUVcXdkSFOIS0AkV00iN1cs0+QGCzD/7HjY
lQ3l1Gx4xPNoqrZxPu8FDWyrhBJ9CmMKQM7dUJtgYZEUVEQ5N/rSSzzwKmZWw5ZvmcgmzsBJ/NgF
7IrQoEKtaJHBLKTUVS+jbsIlfsKr+Ix0PF2Jn3pt7tULqGN+rRl+R6iaWH45CjqSvda0fL6FMql2
WOGMsQ85X7pLsog8L3hqaG4cnktu198KUwy+jxQburD0LdRXZZ3UmzBbxHvTijnVQdW52Ewsvmy7
qG7umcZDYp5kpHqtJXWCEuGGINmC729dueu8OZ42XjU4bDhwr8hSWDDQDnC+2P93hXoG8P31aLRi
YfSWkk7MmH4PVvXPzVTtC7ACco+o5RF3ZCEJ0oYRHWOl51tnxTo9Cue4AOw68KJ8PZ+OVOtSE3PJ
Gem13phrS3ciJfx2kBA0cqW3ULHBGhUSJQZRuJI7sQknV5Gvk7+5BiYrU4zsic2SPe1/MZvejb1c
Bm2Pnw0OydE1Q1tzt2Gku2IAZ8WYRETdHQSN/lpUGad2yYTIkPlYedMpfRFqmwPB63xybN3VLTOp
HQ2vdf5oCnQB5eg7jDjh1FL6mNEIpaXB7Yaalz+uQgC3WbhWBWRlI5KAXzebrX0E56mQxklGFXVu
gPzrxF6hPCc6/jVfUBKhA9cTUiZMTmsYTmCzZ3rs4WTeegw7WDdVKH8wQ1Xr2g/+N6wftUVPgll6
OXD5oaw/MGkn2u0xcEFrs+5q2uDqguLg3MyuP9cWrP2KHfb0JB5EdMwwn74IZZcX/unuzHJZEFUC
c+SvMzOZVb4vSOiCnPPGRCa9/5xoUgOxkTTCAsxJo2jeN2m/dAsJ76cw6RRL/A1GkHfdHYhrzLKL
cMnQ9NkHTjxN9xMTy+TzaKJqC8hz6NN9b7w6TRnn6/uqJshn/YYljf/ZcMM1/VAnzEeb9JVFUaEa
ykQrePpqeh9Se7I9Yxz2emUuGaIc5mY7PK2y/cSoFN9ly0fW2qa5K2uu5WX+/zHBj1DqwSTGG98q
RbvSvgf1yJX8R/lbn0l+yO/BymjlVyq2DGiHlSmNMLRtTYgRhdfj4IH+0LOv9otkjZ/HhJrrT8Ki
tRHM2zZxUL4tgGWsd7dYFsQfo7YqPqLD1clQc2e6ywOeO6vxQ99cafTmI8xUL2yU4+n1d+bLA5IY
SRJpxr5DuBbPS6YC2ycmmylkBPIXigklUvrkupaSs5VGEmf3twR7kwxI2SfJxhE4VUZiMXWIt1a7
cV0U5B32uufG1AyZysAY/3H7TbbTVXVJx+5Mwje1//OUhPKHetOxKw/JZbA7WX21dvhH3uCikNVx
ZjZF+w/omPvdcixeDhUE12PNMKJA5KlQznU6OQOZSdHfiAPJoZb3KXUgfK5VuccburbQnWCjVVcJ
z0BnKJ1s1/f3FPTMEsMLzJ0VetD001Ic3h9Wq4FulWUoWlHH2+Gx3rwxUjT6G92eq0MvDPmzd8rB
z9TEf4s8/qLe5PvVoAzDZesix2FXvib2wmMfWx7tQ0XBJgEYUw8ruerhp7L3D82eZnZgt0IBn6ry
Uy/yBP+kxBGtpVTYYtsXjzGLzbAuWQ40pWwea2dxrIO6cmMygpmBopF+bdlnV4AVvWgDyuKq87I9
R0kjy/EpKiDRO6p7O3Dgf3jR572z373dCcYN1tvb2EIGQbyhAgKR6ZTkYPSYL6gPIReqsNXAEiSo
jgTRuIRdXSSL67IIDODit2+pfwXfmU0zd78c0NPYu90qmmiBdCvzlq9xbCSjgL0a9tezw/T+OlU+
uRuXe9oRgPTAvDNGDWx76fyLD5j3TNr4zDcIAapZ/k2KDZ1UkzjAJQsW9IwKMI204DT8CNn0Yqfp
dcyKdQWBNmMmaot9yn1T8nrI7JZ6PQuT+gey65HQqRVf98edEmEaXhSvOAZ+mwdOitHgcAeV7/SL
ZHuHqiAL3MUIRh9YCV60LlyzTsng+FR5Qrvv80SyHD2yrgWE5pOT5YmXmMe6QpKSoeXJAZkNl7Mx
0r20/8/0fJiI1c68MxomUfEfQYcAniBCFYJ2ZicHQe9pEgY9kkAeYvGRXwuP0M3q4NwKmLKoKoVF
FgIoZML9bGtHzUckNL+xjLFYShk6FqqPH11pk/amrHr0eENRXPtMiErOM41gvQgOc/XJEJp6N8L7
0vC9TXu5XDSvaDml5eKxOpZ0RZl7BWn+9UpsEYGUsQa6LnnktRdotWRqFMDX3GxPqFasN+1mcqZz
Xirr+jdPZxXSIHhX6huCQA6JrLr2VzrU0HicQCMVEGPMqlEqsimY/Gro4XQBu3q8WQ/SDsODFlF4
0Wd7EOqYvyil+XaGs/NQHpLKSYZWVXuQiAYEg3nR+812g2/biGsYQQK0vgaXjqGdK1ENb4Sdp7wY
EH2yvaWwM11nik4Ssphh0ggDz21j3tHrHflTP/xxSF5AXdJwuzzcEhy0Mvus9IBmpq83bI2Ovu2N
kVzkvGzdWB3Htkt5DI9HZgL54kvFt4t1ORxu1x6Yn0+NnGi8SIIDC2Edupka16RfVEouJfly9Beo
ZULmmUvNT3ZLKA7g+jrEcnby9igyBR6ASLazrIMQGv8/BWnnHnT2kK0FCD2NXLhRObxiDCO5IbKw
zp1IneXXIBSY3PeQfUXaU4/FsIz5tjtf2FVlDd/2Y0ctcQR22sZuunx6Yn0oFu++nQQKlbyxYlmF
Y12RaByRp7+ol7Xl4DLDMZPxGEocbWXx7OAK
`protect end_protected

