

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gjKSpUobpdaEiN+EJKINegy9RfobWzPNNvSuynmxBaCaiXpZzE42DUdhJsa9nuNl5zrnRUR14CdT
xujtPqnMVQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VxmOSrOiNTkpjQCdEraeE2yE2mnMFQ7pRVDUX9VslB9rFCGD7dNvbneDVpuQoePUk+nSB0IAqnFe
/NakjC9Wt9azzGAltfbGlSpsCZYTQJMARswgnWL4Fmc2+3tN+okF6OFM1YLClj1yRXdxl+CDsxQ1
FBT8tPlhn++ZNTP2k9k=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aXqd6ynCn5cZfxJpxEun0CmjLX7cGy8EmIQDak6IkAJ5uWqWXRabnrZlR7iXAJjslJ8VJzSbOvYm
rNknXsQKfebDaT1iefkZ0I0Z762iOiWvIR0eap12f4JcJvz9RAzeBAaW4ZyAkczx3IYLwFNzh/0g
2pHrl6Pls+OFuVt68hp3jwzH7c003L035HPpddZ6HFBcZ3MJeQ/LoNxx+FWSqyEG8xTwd196QL6n
uNyNqC2ytbe6mU9D/s5w5KpomKyiSs16Q1gq8Rj3swuI/cDlyu2A84YTnDD1OVt7+ooOZIymcF7C
BaBzVPlYihS6ibZatAmcUNJ2pZYltRbTtDOOXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S9smd62+t/cc6T+Az0vn0kXxFJK9ox1swzdVaJK3ag284vMfjrlnVswyLQNkD6M2BaUNuZuzevou
xaHfzJcTFt8YvMUaEn6TameCIs5/mTCxVsde0MlJlF2crCf3fZHzWj5ooeKnlSFJXuUK/R6CGS8a
2vO0yBw4ZENNd3h5OqE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cOFUj+LOfMo1PTF/10pikQPB0v1eZ+hPEU+cjnPIX80Jf3IXfuV5X+QqrEh3UZH/0+YwNN5uc8yz
3GcUBcrBnY3TVkMqnhGUk3sy243Fxp5BXFf4yGZm4BbuFXxSAKu5Q+k+UOvWrFZfWdNI4lYLdSEu
b+Pg0ebBc04YBsQL8j7TFN2y60Hw4npf4Ha1Oh0Q36x952OAGQt/kpvEYJz+iBAv7Wj4b3IJAFhe
Hz1SVdnrXpsS0DFFqDApZsueRszhz8yuOSjC5Se+b7SzsP1onkP7OL41tcS1dxgV6XpqQDe6m87o
cIvrt9MVp/aWXYppakvqJEuPRZUIN54B2pTOpA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
JOXrZ/2fAkPxW12uBd3RMeUZviZvol4JXH2TD5bik/K53R5QpGHASaLsSKAcNqMLxLONASNZLC7E
RNXvvHzjVW8XX5ZW3iXgAfrjOuQl1dkd8jG9NJmVxyGStHgIk4ehdx+NIY/rX/FJAfJFxezqHUzJ
vrbySx9dHI1VVdToXxnrZBxZGxhObWXQLRfy81EykMONIXn4Rp5+FNVk8ZRBBV944svn3V/iWSWV
6Av7nbvg1kO/kfzKdYtn5L3yXqnCmlnsi9QCrVePln+ey5jk5HfsiJxdPuKNg+WnearU1fv9G8ct
122BdB6JUZpF2PF1m86Zc2HP7JzfdoO47QlwdxYqbr8e4c3VuGdqKw2YzlqM+ISnCJKxbWujPVWG
9dO+N87zM77QrClN9ZMABognV5zrxYlopwBkhsl7nwElAwPXv+aWr8y0m3gXOX/jyMO7r4kQ7fBp
r/7voSu8kBjsanxHY7iOyzVMXEOOeCizM/4zaurofkv/EeKjOSxU30dGRcizACt7EA1PAvN3bcGR
0NyUitCT8ZTY8Ej8mQLMME3cy7gRNKixPlNIOw9IeP2wPJ/fn/obn2vi9aWgqIWimwSqggojMuVD
eXbPUVFtNIYSLPlyKZlqixHa4Z8y/VGSxWqq8L6rpG1KTo5OxvV2adC9AC0tBM02jzRaR9q+puMP
Xsw1apY0iYkGzS+rj1wQ2KanrASmfbHoXITkPU6F2TJgeEtqme+KACfBjnxD21lueZkdMWfwhrhb
XKjmEx7Ul1rD05Ek8aVYQ0FEQkOmylx5lBm6N4Yye1UYiFpee0hWHg6xc0ACnKKm1Jgsqpjm2Lx4
qYjmUh2D6Gb5LG33RfX4sTewbnEYEMvocp8kOlxd8B4PXjumRVRJ0aJVt1k0fH1XzKPoD61cc1oW
rRD8/RTi2i4V1DF0F0Q1Qhnz3vIKQSaIul+H5ducSJ4aKeAbcJXkST8N14KfLZNFoVV3j8npg7G9
blMSiBqheMM9OGpPFX1aQL1Mnm6tz0AIQJJxcXUjzv5V8E287T2nn3xjv6m2A/bahRpADFUBC9Af
BikoY527BMFAekxEUHxL7zWH7B0j/AG/EvLDVLRmF3DGjfWs5eZXCh+Nc8QywOn/BNSBC0HKgT+0
3bznKmIlDVZ924TA17mfewJpyNuSwzbwnlCki3AI2ckgcCtllKcHAlqCkQmekUvmn/PRNnZIdHqQ
gukecsGv8YKzcbjgpuIzajrhWkVYtT1/T98qdygbjFvuBgNUKKcr2KFkyOQQr54nO5aoZmiuPLXU
OXWpFO3YmZrepMsWBE/nWhULhDJkDtj7u7dc9TtEWeDk9mrb/Xllj1wwWIkAJhLjULlDWVyEc6Ca
ariJTojawm4MlMF1VjvSwIDBlbi1B1cRjwwDtWSDRnqJU11+ScdekL7w76fYqnSZC2eVDsJI74d+
mF4owmgAqKs5Tf6gEr97zXkiQOs++wU23OdAHB89tzNinhQBQxymgzHrIPosINQwIZ44fgbhpN06
uyDmH/rawcxnLBSIJFKQ8anwK2LbKN8FlreyVawHjAFdBfqPj3i+KRGRxOfpUQdTrnWvreDvdvSS
Ha6zoJ+X8Q7dGj0v/z3gcSdV3haVUfgY9mg69576wTQaoiDsTJmV5kcKYhefRXXwc8liCgPh8i1G
wAQ6xip/ubZk955KCCCvfUrFw0WG5I2cPyjHwN8LEtDH1ldv3bwVNjPbRTPz/S/FWYWsti/Ex27r
8j823SMA/xt/+ciJeqtl/9gZpWbvG1vHZ0koz8U7gjxj/iXAwGF7RLFahUPwyhav8BSM5WKFGOb0
nbkfGh6SXb+rUgD6OFnTaIdkjw7H0NU1698gVyiHhyQQUoteO7Vbd2l/oa1/thk7OaY8byIeGooy
XD9KVQzWn0Ps7Es3fVsGOfJf00AnrPkEKgVlcfZyNJWUZ9+73gXWmmejRUZwJNz0vYmfiJcIehh8
yJbyh1o79tDkT0gvTw6UYbkgmqCqtBGpzlaJilZBgX/d8zirxdRe6mWrBcjNPBrp7xzqH63TIR6g
AdJk6TJ+kyKhP0Rgl1E0il7UUT+D7GZ9Np4DLCgB+OOUojH55RHXEmoVinIlHSNU4oZdAm7zR4dv
QFpKm2e5ly6uvkYBKnFfojF6MlTo3Yk2TkAhD5Ld2jWfDBhNuzemki1v1M2B2MUR4sYAd1g0G2xE
Kgr/9cawq+zhzQRzvdyJEYLeTUcWqMMdLiUkmpP8kXPxxVcffSxLc5ewpfm4m12rLLbqSzcUpxkN
3DSb8CJb1YVRWEXkIGqkk6cyNcNcRkKqh2b4nh6fviuQOBi2HqHXrQarwOdUGJORQMGl7BVd8oHY
emYbFQUtFn29OIwa210jkkmrG20LwX3cdmYVfvI5jLiPAJrpX00rwLwwjTjNZYoHBOYbCNi/MDD1
gh5Ts2MvCudFtFkjygP4IXu74evV5pjNIc+D3VIfHLo0RA/86oBlJvwtpzEdZXsJ6D99pyKoVme9
3jx5G0MrAn8VhIBvJJdpsjx/F+/YX6bSrFRtGpAawySdDgqVT4Bw0ghdn98jEYHhjIlizXBW+TLm
Ks1C4kwKpeObLYAAW5rA3yv5w+lZdt+6GdfnehVUGLy/ostHJLGh1nD63JtKJPBHKmhcnF7q9y90
JTni5LNdG+dnbSyCYj/U6ZZ2a26+8EDjE3sRO3nAuV5bUDPj5oPILYROHJh+lww5akP0JX5emN79
koW/ehBbkx/kJNIKdhGjbzQMVc/9hBlo9AGYSLblKXyTolJaqi/MPHyLZLyuqsBSS0PZ/F9k2+cd
n7Go1vkc+W8/pt3JNxuLg9sY07awf/BwCfCgmffiM5Um2cBlP9q3qE6Kb7l9HRD5b/+sXdhnCt61
6vJjcct3T5LqzV+DFVrsb3lpej6IHoSwwUYpenmWIycBA/hvUObfMEtgmC7Ff3topeQ8TLroMNVa
bNN8ylxSVsvEdHEbr2uMVuvfqbP0mH0j4LH1HJBfFOYqbTr4SEy/4QST6Zg9CY+dNiIeIepuXqZu
x2FNnkvdALCrop/TjyzESgN4BU4Zumdlsa/roemid3SsIvQFe8QNOlXYgtR1Mp+9SO9xO2vz2inp
0UmxbqIoqvNbLHtTcbgYpChZfJdIwh1ADYNGHEBWdSmmM5ZoRTGp2XuGsuKu/qbbsz8usAMs+WVF
LVlqRY0r6bwO5Rlk0r8RZ2O64/8CsoqKdk24Adm8zHYUUGxbr2UClOsnNhLUdnS/J0aboSmBq3Cw
XHRrm20oHUHgcSE3/Jkn+3YkKYAW8/D3UWgvKQ+r6ozeyDzBjipMcJ+KMe6qNolnEFzoaMIVw5v8
SxGbSv1lfVbb6F9zT1Y1Pk4tVAfJpQ45YA1cjbE/4/6SYgPf/T3Gx7b4yQ4iETy04PeWeXM7VZ7u
Kpi+NexJ5I1LhT8kkYvTfUA6f7de9RAiRFX5VpxF3peN2+wpnfn9BjL+a6ERPosWtjYMMhcgeimk
4WrnYI8uYyL5sI17/ErZBudr28dzdPg9JdApoBLnHX1eyBM7Na5ayval6qSs2LKTyiCZCCRW4uTy
Vsq2frlgiDFE0HPyXr7P9R9nGyPgk2s4dxe8ZYz9+WQDXei9XJWLssIQCfXIkLI91kvTVRfMmT+I
89cEAWVk/vQQP/EUblX5TXabq4Uer/dgr/L0cXFj3HnNFin5NkW17yqUMDBDKLMhRYo94NrP4voU
7lL21Q4Qnqm8DLtv8znInXwVcQV9uN3E4bQJTt2aKKbC5oostq6AKyKLIDaS6c74NcDF5f3PDXji
1+RXwC6Kj0UpRTzXyznQjxaT9GxB3djoBJIpYaoQa0KfH+Pj/6Gs37EKoLGtYxUkwi1khTit1pPw
f0Vm3xJM9Stxhrsyj+c0DwiTv3VLMg+1N+hFhMsBRZ+rAgXAANeg/pM/d899xqOziTxgZz9Ntsna
RFA6pvh/suj4DeLdwisgAqn4WdR1epVI38h17jfSgYR9VjgVk4ot0O7cbLDCg0TbOgMah79NqfTl
aWEGPfWmVnBauxCQN6o/5+5pKXINcdkyqWKoKxh72iUy0phlcoYxFwgiVal8gwVXnUjx5Jz4hiRj
WFxDrA7ik43kFa9L6As3uAwowl8aVYhEdOz+JBm7+OXb7If+8lqyWYygHi4mj78K9ykEShlb67Is
gP9V+aVhz4FZmeQ4DD6clNq3GfNJtAEGmQMuT020vf7l4Xb/WR0C+FdP37VamSFYqm6X77PuD3fY
iS6lm+8XgWJjebrxXn7VNOlyHdC5CfpftDxdyVWPaTN3BoyErvjl7Z6P6m7NUX7HUmoaWhtUcDsY
i9TC47UwtuolX+uku7IAVHgLzlGR1kLXW/kVleF71weT/Mgb9bu9ucro8UOlbsZbtzyukeLkOXB4
eL5bidK90wh2DVtksBuUUTiev5m1XSknDm60SRqI9SyEFt/ZQQThe162ekFEmazpo5IaOhTLFiEP
DicjnOcS+n+qjVKNY8hKGv2gM+tichc3mbdPwRmHkJV7Yus6Ms5A0CtOgrknquF8x5tB8poRkHG+
LUwh8DtI0qvhjqApKfA1S/bnWrhtRyGls9YSmCCxA3BSDXlwEDoc9vdW/p2fLXuEOXJbP91fnX3G
46ImrqHlHH+oE7gI7bPLrXCioC46PjMkZjp/HEJgLxySITcquc52Ol2DO4UMlI20K+Sg6R5nx0ua
kdHNV3hhSzEbT7KtdGK48Wcc6U9pns0Cl/D3/tPD7/svjawCE8MpM//q6FWO+9ML3CiOj3mjM8uf
++iCaDSCn4/9MXZQrunwlOIUXosCqYUK9DU6xrsNSV8d74wEZjWLFXqDDTiwDZy4/A+7klYUM7tv
4e6tsgfuv5JYNXUCtJs3nYaEq6uIfYCCZRgnci556PObpSUp3nZLGeiRJrLMSuDN4206t3nbTnID
3sL+Vt4YEPXzTzvRqMAp3E0QetHuNm6XvZAziE/AnCeyx9Mb1dA3c0FJ2JgH+djviAr7n5nlZjE1
7xhOXmUoiDSFaRK1/kahrDH2gQ/V+x124/Sb57TuYWwbz/T/qDNlGUylMjk0qQ6EdJZP4ny9xDtW
fgqQudTMkW/2/ff+qGdkr+PHGjU/BPyRaC0cDHococJxMG4Gd7WvfR9a07GNf92POfvJmM1dZzPe
08S+eJGdhBWSU6UmlFFXc8Rqr3bJ/amcEwuQ9Ntdoszg/zrGuMns9FZGGiP6jPUBKOok/GEo+uq7
/8gIFW+Zrl9d0lsyzWn4mQbKBko5s8YsBtBX45cw64PdyNZkHzk9w1iG/Ri4q0ohZp5lKTsF8sXh
GM+QtXLnMOQDmbidqM6QNdyD7pvPtDl/n/Jkoi92YZo8ogmIQk21r89eFdiAMTasff8EqXwGdptk
IS+a3QtaIsrUqtEafm3kUqMvvG0GkooBmcTyLaFgBJrC6llZ+vA9kEd0Ip1mMmMvXfMQ4ZLf7Zbm
JznD4D5eUkSSAhv1a+5d7yJUxkw83E6fylVTlb5H8ggiT7WlkGXRF4OjmyGJ+x7vm8szO19alsgT
Hdd91HghpA4zGq5QxHgPc/R9uoaZoQ6GvdMRhh0xmFSZmXKZeKQH7cmiYdqaBCYEu4Po87jruUH/
2lzlKr//pJDhRqm6skdv5fF89TMPkDk6j9W3Lj63Hh4MmaUM/jmtgbcfXXFQCEL1vtB7sHqhorSr
XgvExwR03BTDLaWylWgaKM6ZqKBsVM/coSqXfFfNMF6qQaeal7NVK2WYCKKgnAJ+O93ROSA5d2Vo
vJQj1SQzMkzZztpSs43TFtoN/mLGNMiPt0fvVBJF/o1hSgeKR0W2FSUJAG5KvWulepk9lUr39WSN
v+GevARScfYi5UYtFQ5MuVD39rEig8o0y/FDHMP8FQ7xtb/z4crNmI4u89rpufAdscatpal1dkRC
z41AFPLcx0xDXQRhDEbQFID/4xn7fcxOw17jDX5JjTBvOWeytqyBPRbNQlpKilNjfWKYheGJ99HD
GfGD0FXu3BGKXE+NvweC05vcSiypHS1fVhnI0hf/CgszjHx3OfU9vpKXjQukK6/P4c4ylYPm8sAN
S3Dyuxwtq1f62Jn7FCGHCbHlu7kNEdj0rQ6+7tra/68Ovyr1WXoXMHpu+FK+E0VfH/vPPcBJ43ul
WohmEdjohbKyPkFvW1HbR/o9XloWub8oIWpPa+ZSZWDzBCpu9q/R6EsZb8MJT/yZGqEF1yjrRt1l
RPlYVPeH9iIzTUnd+EBcTr61jEG1pCdrUR+rb4ejoePnno1RZhXMXVBRPb2qT8dTQAM5GcXEZEDo
dCzH9O6vCbVrUTtO92Y8yKfsg5utTU+Rd/ZuFCawbEgwURWv/gTzeej6w0hHKR8kStWMUBlDv/aN
lGFFI+/RGmHis8errauJQCGYDLZ+1E3b5tCnykNgwTd0BrphQtXRbu/4GdqGfFNcPLFL073jpBfg
UfQPo997cKFBYvZBfD33s8gq1FLX6dD62Em+Y1uQSIH/TertZ851sfMroCIMcCOfzj3MGVhPMOgS
EESwl+/gUBbZG4KfzJ2TSK27Axd/azfdwBWyNpmzGRKZ1J5m8XglhgtDUnCcJHeDguI8uM7mF8Pd
DVktVDi4zwfDLmrvEsWMQVxr0zv+zf3attK9pZPM9t82wW5T08ppsxNto0xwB8yFJrqaKPmnrplE
ZsKuNjZlyOO/sxkvrFrMYY35LoNA/9+Y0TpoeIW8XR3b3pTwpf1tucdsQ2TVd8P+rz0lHSa1ADSq
rqu/zMyJ3DQ2RLv/DWuGlnsM4XmH1q+cH91xAa7ipwHdclK4OjP2bNmKMc4s1vL2DH3jKHr03920
Ml9wsHOaUlru1SJgrxpFoXfJg0nkCvnXe2Sp6c/PqqEnb6R/xbdclDfb/vu9hWpwryZcqXGkjLaU
ycQmTyfAQ1THPH0boor1+UWYnvMJPizRCLjgouEEGsvC94fSOrHW0hRZWthF6xVNLgeh4IvFK2No
bZq9GW0p9DFBOvUi4KojqWDrluWcAZeHOhxqV+IXEI0t/uTunz+qVZwT1OS1BxN0F9iumQo9YGAh
AgO1g0MeH4j8Ppo2ckA+ogGwIghmdJjEfHNIu4f3nkIkjtXXLa13j5yE94ialW6KEhpad8/dpK6A
25vRmoGjbngQktX3uYe+kjjKzLlcl8eZ2+SmR7DY2AYYwZeBhIUCwPzZD8ZO0MJB3NYZVG7a43L8
vsIESioVnDUTyaf/s4Xr4Gv0ZtaUKjpr8yZ5KjyBG8CeXZDyITpKhrSezjzsse3IcdciaTGrIz9B
XvBB0K2ONp/DjkoK3+zCC/phCPGos2Z066GvjCaYRkBBKgVf3CAXBDJk8TtBuv5GHYyB8gxTnOWh
+wWgV1kyY/LtsV3STJph2+mII3gY+pTlrIUnj6RQ+ap8asb6V8cdMVDi7HeGbJM5AabH8fdlS1lf
HYz8b0ZEcuGlt+ex78C9X0+Eu6o+hVbfSgdhITm+EgLIrS48DsASDSZk6MFyjhI7lRKr8tZsUSDJ
itQWCGd8tpIU5EfPPIg/7v2cp2K1zLD5d/iR2Y3AW9bB39xns1YiMNNJ3753nM4uuUzoX13OTWm9
jrOYzMyVAV1YluTPJ+Gb8WU3r2GW5sPsclRia3WF58BHTAaFQNmdzAVFUDuaUSE7o337A1NMWvXw
9NWv7j2/pbex8QhOi1ba+yZjCkv4XqJNLejPZsv4xQ3Ri9q/i1hUB8+QzEWWLMoGHhlras6Ya2w2
TPF+ddu/D4Qq8FTxK7BvoetBIa8QY4mR81fxNqQO0ib48dyyq9yOFbMFUmlFXQtZMyYN/aeh+VeX
isUF8tcRD7WpCJkEcoY+wRXd5SpbZbyRK+aKR5tGqjb88nsFeAEDAMhxlBQDrLuHAUc152B1sl5o
4NrAGUXnCXBSOTDGDAJ4a2JkHPdXaxuCXoGCTYRYbr7O+b+dVKq+xu+e4Gs01zUZs+4DSM0k8SvI
xSDYjRQ1BVCBuGRduQFlfituQTltmnd1KxBSycdHwxCSoJE31PwaMy5LSY9h3dphrBg4ouat8D/M
e8DtW8jRXh400q5ll2JrkuiD6OoRF8SIWA/yOnKH93P+QhRkymiwdzxFsk3b70/qClOA/84asCAe
uGAEvTBFRxDbRuP6X4OVL98XMy9AbW4KCZzwaozdbDZcve2tbUccXgfjGnIm4geUnd4VVCWf3TzO
fBA7HmlCDSIKSp4XixHjJeAqS3fIsJpAt12r7wRdUSEO+rOIXjHTeQIQgkEzT1gcMjS7SWfC1PIx
dvUuvhJpBTrR3BvVCreiUMBSxRX5eRzMC+59c8T+CqDgpLP/YCpgbaPqyg==
`protect end_protected

