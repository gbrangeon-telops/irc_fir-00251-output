

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VqgplFNkI2rH3rP35CdiLJAesBBzx3ahYCWVov2QY8pnSpbbPHZzKXALTXuf8Lg9RV/60SesvL5+
Tx0kf3Xi2A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YpVJ/AkbT/7j7nP1FpW0u/1drBu1Ym0xSQcZVVNR2BH9CeGHgikyUixQxXpCsKnhOEb3pzk2wV6b
2udOCqgzaZfDIjjaxTt9/C6XIY+oMyWDycOTnGwR4Bf/A6rFEzTLA91kxNt5/tS1PVy+wjb7FCsa
mgkYj9eNUdtmSsLezko=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pSdvSF3+OBx+pmFIuKYX+lTRtc2CK1xqA/WmTxOA/9c1xuF8tv0giSEc/96tBGsFFqc25YHyYiXZ
gYsCabVJMk2jc2XaKW+XFrRUGrQYLd+QPrzsIggnGqpN1i2vEJ2/57QIQEt4pR4jX78IzCIP9B1I
Mief83M338G9aIgdzONBxsD1Z3XK2M1fqZBI+UT4b8E2guDKnWsCC9f6WqxH/+ijAu2o7kXfkz/w
wH4eaCjn38eBIq4U5maYpwbVxvzCRoB69hlCwEEVDievRmXHouMD407mzOTwKaIkf/tAbFyB6i0D
s5Boa+TiBtHShhLBGBRqGoq+2UpGEaVgj8o3hg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HVe+dxCY+VHrZ/rUbzyWsz5ix04KcDyyUrFaCcS4yZ4GTBKi9GYUFVfTsXMpSX8pxXieZIsbIrAR
8ATsmu7QwmViHDzOMuS6sHzr6e8dC4A3UKQC6xKKwbJdSWPz/il1AOb6t1CcrpGMLBXMZTBj00R6
KptQtwRx2C4sHo/bHEs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gr9tWfnRHlUz7X9jwun0huNacy2IvVfab84T3X/BBntsyGpCEQL6hR0/eLuvmgsVt+peH9UtRKIo
Mx38RlMVlftuoIDUnixeoGaAc4c+4+tb16q3/5V7og6YvplXdBH8LQEEDNM3+H5ouvTLLeMul2Yk
sNNMGtkGcvzxpzj7QTVn+eSHg5B5sba+LhJuLxq02/5r329tzFZy8dtsa4HltD5DQbMsj44UHU8g
J84rl4f5z2tzAq3mdpwIqfhK2vn+BHZu8UlcbrIJKEkQpY9EPDhgx0vX44IIfHNFCmG2MgNy3yn4
3WNmBdtLjzwOjBTyBBtqdvJWbuTYLVDhGJrWQQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4656)
`protect data_block
t8iq/Gp0bVqOJDpk97neB7WaLDsHnScncbEwHB9CLbWZ1d5ncY/92GRmt/u5BpX4qPOVbpVfgTYe
V70LqsdTVX8LyONrhdtpaK2hAZV35D6XG2dXLREsktF4PR3mMMfN64Ryj5jk4jWJChMJnawG355t
oibt4rowjn0hb2LTWPoGGLwZxtXfz5dqMH2F2JuMgTzkTyB3/+qA2JZeynvmZkbQUvU9zGOL6QsQ
/gBMpCy10QYlwNtX0mRn13Eeq2EHK+c6lIKDzez/th3o82sHf+Ue1GlJOQgsHP+X/VALFQEAliWP
V9da/nAIn1MZ7vo0c8b+1yIy7TgJhkXjNGUMLxsJb/WXAnQc6tpLAZzHIC6/Z9yz3UVOAe7xQXy9
l8NmCe6mL+BfX2lrO5/Ijo+WN4uNUo3IMvUpZy0Sn2zaRP9RabQ78iCiUiaXNxfC36L8TQp/o0GK
fR1hmovJYDyArSoLnR7iuoBWcl782GNHV/L2f9Jh8LOc4xxsPmf36gxgLdLn1P1Qjq/Q9xh4Wa1X
lKEqQi3TqQNdeUPYLv61x0oViUk3WlnCS4dp583o8ZsF6DtJMvxxq+s4u18U/pNSWdFiQeftnwIi
R90hquCeztuk2795CgMWpRim8DViEuTkGlCXDLO94H1YLq8UV6mPOpY/4EebAc3jBOPnVy4AAvNg
EQ7VOG+7GCJRur0uitJ4hnFQ3Ev6Wp4frVPQfsEI9R9CvD/l2/Lq7f9iWPwiUlMKZy59Ma9t9+1u
Nw8/CpGnU/aE+HAUFtWObAfmcGD5t2U4yOOSa8MoCBQt8Odtz0O1tgzugSNsPBgdqizYQw/yWXb4
Km2ek5t9tkXvr0cRFlT13/af7W6zavbBzFnombloHEGq9vXcIiEjfhKviMc6AYgu05T8E0JiM4eC
GE5VYWVmwnG54UvBgfgNCuTJ+6s6H9pLnV5pNdrgUVsuVtfCX93Y+MkjmbirOmihy5zrI8FtTmqi
mECzIyxBF26ziHq0aLOcomobhC+hRuuuOyYHyBi7ZcjdsEnEd6sx4UunCQ20eLGk8yvvNII0xFcg
nDfmSDeAttirNmUwd0xIP6MxOq83OcZAnIsln9h6r5YS6jondLdC8dN1sb9NNzgxeRUznLAU6l2u
ohrhBd5HUzM8E4Jj3eLvN8uFRVRyCO+izC1m94t4xZrS0dYgG2IxJFLxGK19UZ58vQ+5m6/ACOyB
c1HOcpcTb0U9VdrJYd/RbWY4iSuxdw2LhRPw3hIIrngBBbpnmllegiWW+ki+R/G18LiSH/ZLd/yD
WHooOAqZEAfV6JPlGZ0GNjLPYdYqh3U8bAVox9swwmf66ozQEX89Fblk/lBh7Fub9nkdM7mIe4TB
YY8CX73lmZJUA7ONHHGDa+JH8G6byzoaHKaoK8BSYnfaD1fXd93QEfjpmpdrRyfmVjyMC4fX9Z7N
ZdJ4Snrol/ec1kqOjK+OuoSD1Q41f5/P7M/qJRyxqJ8CQhZHAc4W1YBM5hf8CPiWT/ny5c+wEOdH
/dpYcWFSOdc7F1QrNXHzw0+5E9VAt+HjtYecR4ey/EHrfWCDm6PSeHzeEl2jddm6SMQKFXvwJq2w
R36oHvavpk6Xvb8Cjo4c41OUzlIPKL8O2H3+iWo0lJKRZ0Ivw6hN1M9SEMEneIbJcepsdNXGjwWR
1GzLozvpGH/ciZOlGHPMZlIRP+QiNSi1cDSleZlzU0rsrjhAUznLPNEgt/IvBs3RjuQq9ms/pFLw
HuiCTFIy8XHxXeEXTcGSnPQDjW2evM14NqcZo2MdZ0aIKo1oTNb6pDi6w9TctmSIxZXluDabN5qK
cms9NFLyJv0FoixlGYvLNm029g2DQ1bjeNrDsIn8P6kVFRlYeD22qsZI+C8FPc+pdGBg7eUImALH
2BiKnK4T6wlY9e1iH2zxzWlJ5KCn055m+jaGk2ePjzj6oStDpQV5YEyybkLdjOgtB5QjF5esz0QY
YswnzCmf9OezRizi+EN1Xd5yIkJNWecFTXbhW5sxdtIbS2AT8yR6NV2BRzQHv5cyD7N0aUv/mFsT
FP9WaMq/yof+Cd+q/fN7Rr7/MrlQzPXbdtD/4Mp4oYPiNkjKDF5/uidzJW5Z2bS2o1ktLYA4rdD3
tRSsu97xolLcCkzZe6+NFnNZ6oMPFpmjFoPB/05pr7aE3kiHgV7uJppAE/Zgc08N2NbH2IIsGrf1
C46Or6+jAWO+aiSG1t0kj1HEVChwdiOP2c8yGI9Yd7MNun00y5Qaf9G26uJMLdfj8F9ddy31Rm6j
9SOOWqcMNsHM0Oq+kpXSr9OmczYizRYA7/JvUGgQ7bnlVTbxSEcRgJs8dY7vBt8RK9pMmTp4JbEd
y/fyPzcMiS93hZ46OTRNMoKXN37eRhdmVsT+YNYU5VOPPjRzNWp7Ni76Aew/+ENtTpTz40BBRx8G
8CPtZ5UtSi0tobdulSA6Vs93hw0NQCFC9LKEH50DxEAKXntH4iK9a1chOHTPfOQSoqzr4w+emaUv
mKLSSypw/tXBUNxSrBIBKKAmO9JgpKx/8B67iel0BLxtE+A33fD738YPmlVEHtx8vf5wQfvlbndF
Jxb7Z8sJRFQA5Nad5E6yFt4QkjRaMVQSv6R14NelSLLitAjN7HZJAmNuCOwLemQ7tsaUZqZ3HpNM
4d2VV+Ky2iPxSC4Q0IWKtY/0utVgmuakp0cIg9zPvOGxA1oWjHTn7uYFap5L8jq8VU0MS//xj8Xz
+aYY48+S297hhwvbjoacF1+QqUAf0f81TWlMnMFUFfO4sKrc7Y4AM0S8FW5ykyEmINmTAlKcswRC
7ZuPXUwbs02dOctqHYJPIaDHLVjOdUITHw2YHZOmOGCjUFATF9vDQRSdt36F+07g9U/fEHIstBRH
qZ0nUh88DYiQVjbKOee+TzR9O0TmetHJq1cQYwgcibGi0AoRHzjhxK5rS0JKpJmev4va19fV/F6P
I/GKaOrkuOZUEe1iT0SuMMZeedWB1LVAb4YQ1fUERC6kQWuMPM91jA+j5uHjrb3Je3pSmIN25Lwt
8Kp35Io/2vc6XnQ2N0AkHwE+1NMddeuxhWbYkMvXH9N9MegN6+YPKkKSMZRCB1LTbtib0WVI+JCl
GN4FUOvcb8+HR5o31Rwf689uSoR772nSh8XR4ojhsx1nHs6NgayBX8PpYHH2bo+BhNRWmnl9fuEf
ibmpjtnKfyYa34VwA+Vf42zeLkOOe1K+wA3xw+U2zQR0Hqa6QJqFrVKx4MAh8TImgN4j283gkFRy
Cc94hmfbMtxFSKN0hjDBe7ThUSGs4AdRWyauhWELl0+nVJntTo80SeHpu7xilIe5B+05lIwE2BRM
au+FeCcp5szwOI7pRsA9Ep+EnIgU7hi1t29CeqoyQOGmDo/wloPGoa/qCTc+UNhiq7Hsktf8YSzj
YGXULn06cHE3+S5/VZ5u4/5xruklSYNf8/bqPIai5bYv6s7mn+EorZOBWhzgzf8vIhxVmRFN2zhK
u/mApgV7x9l14A1ZXd/Q91CYv+oiAz4qpdKQ7AeRIM1Ta3+mmGHBkTt+BCZ6Ue8WCijLUY9bmhUL
Z/8ayE7mu+iOncQ9XftOvzctkvImB3h3rU32TB5HCr+u43lqXM3Ozt1JNsxRHvzVp+ExjUA1eAo5
+V0jqqZGz5tDMF1Defw8YPaAo2QdllRjfMCbaNeYUrYMgAnOVRpYiym/EWV9N/cGyRP7wR+HhylQ
4tGfLHeud8L6dPvvQUyqq7EBPqeO07WbNvLiqxvE4lIva8nPhguWbBPe9qIrUCWuIaKhl6ZoODIX
s6cB4OHhOgulucGC9qTIFp2gB0lyzpbP6eAqBKvD/z4qAYf+puzq6bBzAwfT9KLxkYchJsmDBQSa
TNmow8K0p7RaF9uTfbWhna3+Nj+iS/7aQYPwmJt7z/HL5GjGiGYAj1Te9L5J6ORjFUoRBpQtDnX5
k9+Y7Aj47BZkglNq/wVS+3ytYZL1MikxZEaA2Lvuvfz6RtiBNR+8xphb9GYV/rNugJ2/Ih00GUFJ
o5krR6YyWCWKJd1zGh6u3TjwzMilYQS/a2u093F0EWHb5tzNt8QnqQ06iAyzqvvFsTGl8zkRbs8A
LagPhZDJD1rEAs4WqlICiY7evU9W0vxiPLLnf3LUBmigeOjgOGM1RtEY129e53hZL1FJvXVMthNI
ugq28vCl1sB1Rma8LuIX5OXI8q8fH9g7Qh4M1pOSHVz7bsgCW4u4XFe6SoGURdF8ZJkFSQwvorKb
gr1HvI1CQ7WdumuNCUJBUX4OAV4As4aKlfjcaZZ+TjqdaXM+JHKYZhDUFq0+psfVE5tfofde0GEW
jl04YFZGr7LnNDjOqEyelmQ7ZmQgR5hdJYr+jXMyojyw7uinq/jbAr7gkUa4ayNm7apxvssbPR5D
AzcQU6BpKtL8zNKTwykE19wwpPw4iVI8Cr5MgL7jYEA8CvZsRKxwcf5qNA8HPkME8x9lfI+IV37S
+4zIX1WFSvKsgreCp0TZwzrA548A/v3n4d6Z2SZduYVIPoDbAzRw48pw5dxUp0Kd9JYZPsK4Ybwh
vHL0MaBTdCPYyGtKfrjOZGYUaDzT1V8d4HGTM5M7vBYOiso2Kyy+lK84AkeWX9wFqEfQ7T1aYYCd
KRRoEVIyraRyIrrFbVXZXs4Km3JaLfFLi0lGNzXadqwwr3bkj+q3MRGkxzuxR7H3lsSEKHmSfnMg
jqNvcauRcCM1QAyMzxPV/16IwBTPUxp7X5+wizpaHV63DAwNiLlKXjCiwIfbXMMFo6+f+aoAltE2
XfoFmBKRIAhfRTi2BgPVkE7IhWkhXfxwrsZ16839+0DKAkCEbB3UspdySys4ThEKnQMfdyUIqIXP
YSQ79ptdN77jRBarIY+VkO/4NopqwzjjSAEr74zOpPGSfFI9yRsDHr9osArf8h9RugA0fbGTPMg9
ALx6DhKR5AIVu+Thh1ug/98oA163uV01ZNo0MYBv4pAV7tCHXPw9iq+jiCs9x6Yo6Il9We2tKVVR
NoN2dmhcA4zd/Ko0gH2ZimcmVXkYCnQ/kh3OhF7nPoCYzjahxgYSKeelg4Uo/AbXFVGVX9JxDwSO
SGNgoId9xLVvIvIF5pJITb396nfBLy66woZOrrUazIvhPi5PUTQeH2BodJY6CZG3TwsVS9J7d4C7
YV4M/L4pkvR+7oH2TCsn9KhhrS5DEqvEDzHvGS7OISrL7l+SgVmNht5MXBD0sduIUB4d8NaeMNcc
NCfkFjWOG5nvYcL/TmSIeiKelPc1Dq4wmyFP6aCRQrT1RIIfN6NlaH2lK24gN3O9wFwIzQ923Nn3
D05nqZuBMhAfd5WNz+XneIRsEu++cQnzBGFLIJtXkl92HpNc0oik2yKsf0T6c6xtOwUXh+mWcrO9
WU2NAxPVg8vCNP/NZ88O3xu5jPcq2THftVS+8Zn3bTHiP4v5AEZ6URQOTbHtWW5vtwWsUTlfHRwM
59bFc1bW1k2pDtSWazjnUwiMl6zwcP0wRPvMTIY2vaEs1HnGDj8eQCrekkKjbculYQnSOGCzKgZz
blXTTo0DRfaUICbLe9JkBlTqb2H7q8ofw0Ly+BAmDMstsbBAcgxEJhVfBC3eSXFBpaVjXIIJcJ/i
NvTe6j9Zwt+oU+0I0AUH0N6QusKv5F9t9rq2EPaNfS869Ly5ydq4zL0zDwi3SzfjfjXD91lJwLO0
QXzi5VahYAY0GQLF2KuxRj6JGYEacO0/oPMdVhNmFvUxEgtcZIv00sixyME8wCslRnE9g106Ohv2
/H17saaAqqfKTaB9DAgkGp+2YBNjbgTMXK9+yFq3ffgXKY+5VJC976mJcfkmBs5BJFpNQdSYgral
IyzmfFEd6g0ej6AqZMr42+Kr9A05oLHkhDkVtavzv1hFMV9Zr6NS5ye8mfrrqgPjll0Mu4lqoKyM
/xT9lLsQvUJXjYL+0IwFzdmfaB6BXKoPS+9YVKjP/l1if3RvamxaXWtq0921s4hMtCW6iS6eJg11
RWJsbr3VeyxRA3pQyqG3ueKaF29w10i7FFhqMk2QaAUwmw+sxVJx3RoM+TMcoK4Y43EI99TUaxWP
+EcUau6bunK7I0IaS7VcW3ovjI+JWT9xNu8OzWppkJk07GHUOoDGbSqWFmERISWO7cEW/MemxPPC
A/qkhI6TPlt8JczkdS/Xq9i7T26gjbDkuEBf9USJRWeic/0HJRkS
`protect end_protected

