

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H5lQJsJvaeLLGFRhK1oe708p9zTtXNXItx2KAtknEaAF2yq8IXwKFiVPbPTO8aJ4G1wQZMrKgMvb
6zlyKbmneg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RUvUfs9jruf9OSb6utxk79ymugfgdQ2mgDnw22tbcF4+w9YY12PtlphQ3EwSjE1BR+YNcfcg2ppx
nVp8oQrlHaYHLiZdJQiFcET810isTDBwI9+sjn4Ry8+ftUrGRDkzGQghSG1UFCnSyA55dNVCduAa
//ZGtYPCXRggO0BwEzM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GRoj0md2TTeeyD4XkfgAjr1JI8z1r2plHgATS4H88EONpa3oaJwG10L5TE6c5MDXVxHb/m1WeMVh
VBt3w5S8h9pf8c485G3a+NVnNsA2vHPB4cEC1yhvDIpNkeqj7HvAUARW4zUkp2MDiimsNN00ZMVQ
inLzBlDW8A6T3Y2b3GmoYzUXaMQElMyS/PaVNF6Se8+PIRjTB8Dv5G+A8K7PF3j0h0gW5LdMZrCx
isigyN5NiqJ/3ZZGLkd5XiuLlr0DetrgHdwfifFeF2dmLtMjIx4kUkMG45tToYmkQS3jwm191cux
eXIUgmzmvPZHik85i0iZegdiOZ1LzY1yO5OyEQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UnEKB1f1t5V+eYV1nijBv/smbMsJH58WebxNSKYwmtj2m6R5AlGEZE0haiR3VYCxPRjmiopDDdr6
uBQOF41DIKvZSm6YCypTeVt9WvkLpXTJIiHnLWz3IV+uvKXohhIry2Pg30NMC2EWPfi43aTNvtNH
ROJrUVVcDZeGvVPmgRI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U8EV7GGC48XxGZ3G4wShg05dze1bZdqSUw7dITFWVJl+2U1VEqYTGCRl5zpa3cGdqM2+nFugC+BK
YIux1TwcaF2Ng1I+Bp1k4H3BhUPfmkZlNiGri0KnFOiDYzBROYyyiUUX4IECNCLZnG/OtNfakQoI
AjU6WqtEEQ5JSpZpL5mpGWt7jGfdl9gqPeY88IdcWnasDywKSPqo47azQ0KIzwP9UejnEHChmHgr
3Gpvmrmywo7/+/EQRujU1oGF+ysfAmqchOGtHLtDFJ1h2OjLVkv+puXArlpXpB9wZah1XCGw2FON
8d2jAO5M9wEJ2bQpFyxmedBeZ1Qj0cJQKZW3Gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51344)
`protect data_block
+x8jxepAS+lGyoSdVfxUEyjPWjzBWjghoDnci568/VF8/xHRThUkQnPoCz0TBUNUoi15yVNzUiA6
JgxQp2A28AYYEzYUL3oJM0L+jgU/ZlMKsUlMHiSG2QghuBlwF2IDAJJPseeP7IflNF5KPhLlSQsG
kV8xRkZfq89UkdNwyfsjLS+KbN71/3TZ3PSUXrqN+4vlq+nuE0F8siiqUlhP/IOuNB6CIp+FEkWW
vqaCDSkR3GWhwicQpu1Ve2/LNSYa0TZ/yKwj4kW2LnRhiFHIfQwpFEWilQri30j5ttMxJJ6FFOdN
4Rdcx3YoYnMvsKBnwGh2LBzKVZVY0nbvJtaeEw2cJbOasGntGg1GlzVBj056Ezzj/y1W0v34kJ6X
biQCWgcLRhkDrzNJ54GepdoCj912tUNZXarmUW13J+JFZT9dEpGms2hwqVbbagzDNgxLCbeK/adh
6QQQLrWACXQmka4DEWjrX4IcffKib1QiStFVDOhOnNhttZpeN1VBeXHCIRpZbLEWGsUKQ6U6kmSW
SXuoJopKypLdlSVnCdCLEHK5EWc19UkPQxXFnYyZy8sjsvc7SzNAUb3JA0LjABAM7VmXbON7jyTP
gfkHvtD9u0+ZZBNi2WkeCTwv+XNWK3LwbszOJTkmvYk4oa/WrCbWo7kN6+orNz02n8NEcHrkGR1V
8BX4ByNql1AEiVvK4BCYo3NMPoCc6ZsW+Ylc1ySKAcGvzBpYrKaBici99nkdX45p6MNV0b4cc+Ht
JKNwl65NsIkyLzpn2+rZ4vOxVsVJU+clDewBahSLzez5zEYVQdMBLyWm+4q86c9hn2ZHUcHS0ul4
mc49f/XmQf+2xIW7/lyROoj/2OrnZXSUsIbARYLuHJgLlPxbzEWF2wDF9ohbdgTgN5pXwZ9vLNZi
4IDCFMNy+AiDarAM8a89XLbn1muemtZXcPHf3pN+vz4IqRuOJ9ulNXUVf65U2Bej76yBfDjCXLKT
cjN5IwPSyqSUPq4yLe5hYxH+4cLSM5fHzeiSlBI7GCYyW353eq5A7/r6y6zLFJ8YbwSfFaoMJD5T
ZYprigBuvedYScF3sG+aVR1IgO2OkI4IEeSyYTn2OOXn1qJNZ5e6abFY8LlfYtkAgCwxvGKyYEJo
6iEloKM5HUViAo9f07J2n9caIG7Op2V38FxH0Mf9vzoD/1WgumMGK83F5nSMF/VwWZD+eHYCqX41
uyLyjZmdxxpAtM3uzfSJWMRlnW7o8FhhNzHt8cFcREpMCk+qHHCHxJZmgIRuOe7pweo7/vK+bOha
CHNFSzyCDHHxOSrh1bovr1irz3f0Pv0BFcYK4P1dtw1MH9j5z0AV9XOVprjl/t7cxJiCtxrNPA5S
FRBPnBRRg70iJc98nU1MfjhUZMfmCTmu2b/bv5rouZFy3ujvguQF+zzHMtg2/VDOybSV73N6DD1L
447YPF4TEENEXmS/GCQDLuyh0GJ5nYfArbJe7lZMIiq3NwiC+NIb0pUEcp3xwFhDBUu+3561IupY
nNhfz01ikQif4X4FAOhNGeHv4chLpR9eAiqD6bLiNtkMiVlBMP0Da2exZzy7oIMnXkvQnwtaRlmb
KzFt7INEIP8irfqK4XXW3lJGnNfBpzfrIBHbOPm7ndSlj/Uvv+tCuqn2qU6EMA0o9Se+A3XqnKXP
fOZ/wjuFLARxO/4UgJAA4EDy9At+TgC1pCU0jTNiA2HzlIE6t09qMS4KXo4q16YsntBoDW7L+vPq
JnNXlnYMNgIS4yfwW2m4+70mVL/5ilXbwa4QbkSYfMlvlSyxZOeOAQG9H+UBEJ79anRRcP4+9Vyd
M5sGa1tr0rqGTBW7icP326RbiX4QRYQPDvg9/jEusWcrLdBRjnw4feS2QWcTLObXZnmTi//Zy2qU
tnqG/EbdMikX0UmLTrdurFSFQ5myzEA0nEY41UIZVTPae3cd9iCymYU3531M+UqR6cVZtPClrp+x
zCSnoXQd4XLTCop8yQQrZ9aOeb4E0FnAk9nYutdOYQAu2Et3nKwuDAd+kbHRWRW2yCieikmCycKP
UZbkhlqCCU09p6KrOdoHhpZneovQLpOwmN7sRIUaljUnTDF6hTD+h+0jWx7am0uZ94iNe04s/uJU
+hbJSt6aawS8wdu0BZT7WXcw86JvgXNTGZAf+90yLsNirHSDM4SMcacheMSvba9aY+yPfXhjoD9m
5RWCkRCZQ5y5aFHj1lSvwIui2q2aaHfhZ5KgDAAgYpXOumdGT/mu8EKWADKVv/pL7EM2LvCRC3xZ
JtjnAGvF6k7ESzfUEHiZrfI4G+zlvLlXuZHFoFvQ+LPEYEmpqL4qJyxjbxKywArKDpW+mF6K5z3x
CPLZ7Get+oSn9Z+F/Sd599VXfcdg4bBM97+kZqg1V/DHcC9exeyDQJ9tUIhR7br29m2gtkkk1USk
VdVUXBFgH1YTFeoNF92O7yMltX6PGsnEbj3IGTKttd1qf/AT5JfT2tmcBnuKFy6DTC9PuZk+W4xS
4zmHvKoPChcytzVp83V7N3UiEyQkXKNVElsaw01jooDmOXD+2h7LF8NCmZ584/oDtW7Qg2nRdS9l
DhDq+8toTm8pG0RO2u3KNyGOiahTztn5sd96P0mjETpzgbZ9DJl0wwE+g0CsgTRDxrnmRFvGjxY/
7UrUZ17TNjEj4hXPT3pOO0hv2L/uIBzRiCJubKRYbm/IqbYZdWujIvXK5Cg11TdRLPCSJ4VQNK9m
CDTw3NzHFnwGHLNnJzjXGyGotheOsg1DanEJtueSW+bHkVBHQU3gg5zHKYIiubCFjFt7ATnaDKM9
ia9WPE4gX44Rb/BXKBkyaW9CBKxARXAIVu2khqJz45hcHIwUN4WEfkeimeEmIBOvSdLKGF7Vws9U
fw/8ToK0q5KarjKcoJL/jTYMkoeguIgZH2eP4zxiffXg2BmLhl/D1h7MUrUC+plQ6QJNcqLj2avj
G/oBd02AC6W+4TTVANgefhFSdLI6qQkHN2Z0HrDgWU4aHMBpCvSZ6CtQK8UJm1ceGjtKdzxYNtXO
nGdEv5cDDNV83R7x45XF1kNqyGOSQv/Rqucbdx1vmH5bNWdKjy5B/6Q+n/i5/LwA8N5jH92Vdc0c
Efkjlf0wZ9FrtSa65xLRpi7Pck1BgV/lHArIVHPeQF73weHmwgItQHoPexPLPGfjqIz7NuUk7Jxe
m2Gw90KIjTeSbyiMsTHe2S6nLPMubVyk6hqG8raNjbYFmM62LibBln8dmM8j2nKdBnn4BXkm+4su
vwz2YhPBwIhPCymaf2dzqdCL/Uib6CRp+FsdXy/iJIIX4POx5fLI7VQeVC3uBPo8NbB/0t8mPyNO
WLt2aJ3B++mCwSaxGIcFfw2kr754Kp5t1S8k4gA6INQf422Tn3fugIgh1Zu4lkqliUX1rgJybpX5
l8TDG51f8Qr4GsfTp/FRcUasjO8a/ruqcpzOEigny0pFpOEtlue0L6NF0BBDpHSVuab4x509el3t
cTDbwEQsrvsXVczBXUW9a/s+mhGqqUw1zbUqlbMYgW4WA0wNxgWR8kh4OlnFiNo/AfEueMFlWDp/
Y24HPfEemNJzCh6+VBzoivnbKwcPEgPo8MFW60XSkZJyhzlm7MFms28cyDZ02wgBrwR1oBtunCde
vO7B2HKAm1LhBgkFtJ8Wp5/qUXhejnc0b0bncXZkLqD5/dL79hOfNEjTD/v6qxQsDpNnv+b8K6+G
IBsGOvz4drjiu8xBWGxkgk082w5nNFjgu7qZ1rTooma9x0FnRuRXdnqsblX4Ov+hGFT2//+wPJ4p
UXbA72j7LtnL4oId3cIgkozuM1e3Fb6w3PsQ15FgXHB88kjlBEolq/vTGtEzZkUxl5TVNCVxld9J
pzA3cKYYachDLChIIPgdFqQyICt286O64INH9oDa6dEkffjxsksPFArmC4QYFb+vpmGPMtVY4svo
FfdUcyAzcRjKareo7+5mSKiORKEmwnMUsMAak0SCF5fCvwpf7oPZjHw8lWjNrFcBd3FlGtNPdsw4
sHbm9QafR6OLca8/wLDNYI3Ko2caIEZAWyxU1eNUEyv6Y7nbuJwpfQ1TsLKwLs90P8GqJEZk+UIo
zF67qVW/it5avVQnGQgo4OZgsKzXahPMrVLyWPpcP6/itHmRNme7RDHuZhtfuMmUP7/wg/vu8D9R
UtNlgD3oAYROxjsJHehXy3Yg4L3DxyY5vpQWn25UhHaXAhFJozT4KlaEL2OtQlSHSXz7c8x7fVeN
9+PAMULwapzek9G3tGtmL6dpuTn5UsH7ledz3AdsXTXdmWbAbgkTJMvs8KyIGB/hg3Uq1SR8Ap2Q
oiOCPYaHa4MVLdkF7Y/haU/uPW0NIUbEL1kX0b2ZlFzwEHoOqPkSf3XdJY7XZdL22lfP0sEz435U
d2Hd7mpGdg6aRkkxY+HZkHqo0fcIQ0Lh2XrlMZM17RjZZmZs3xz0PdsEG/0T67yeMtmLGWhbVsIo
67SVAGJUWAcNwYOP0vD+Iht9ueHVOeXQKBkzA7yFaisoKDGDY5Ry8caQtQwr/LGfP0vTb6onC1j1
MLhaEc1JGOfo4q69uuEx7xiPbWUQlmmS2hQkJtmUe7Aa6ORZrYVea6oieGrsf2BuO8Fmw1qSZ4Fc
VvtFmg/4DELOzy8l/yoUAffnUbsuV+5JwPBL1+jW8Ubs7DZF/nHiicrLbNQHYR1w2a3IQOLjJzGd
m9BB1LEqHcqRuRvCO02ZJXSzt0ph+JUvf0BtDZaj5lsSE8dGs9QVdIjwiW2zMcc6Fy5XBfAti1Wf
B8gFPUFAUt9GmTV8HCHXiIrCAtRG50zaKj4h9wf1dxA1eMGJkr+DCeEvc/4Ax+Yk2JsPemb1PnFN
lv9SZAzL45M1AVhLuNGF8cs1Xli7ma+RQ0Z8wQjaPvqyhEZdxGTUqzBgUEJU3To2bglMQMY4WiEF
jJLSXyabeRcXUzVD/s8pDhhg29eoG0+6P8Mgb5yG+kLlyA/ufVEWxM+FHIVbhs40XHinH0r+r9fe
SHVxy2Pa/zA9UnOVC2opQEBTwooxer7/i0ZAAep7XcMVhWom7YYaCRXivOlzNkMivWjR7Cljy1MC
qkpLBuFC3GwBMRQRJ3XaQZnL+9cUT2WsahS21cIE7Rwx84oWwAV9JBYjx0vJvoUiXRwqXa/9uBFO
ter7+Uc9W49NIZKEUav3HKyCH5IkB6w/AdZkeBuSu4A7ueYS15gk6FmCmKe5g3tBTFtE8yvSQOD7
K8ErtU1+a4XihRW6fq9IAigl+NDSFKKV0+8bJrbx/nm+lqqb9vfjuK0fSUUPUZJpxuWiq7SDpP4C
Rtni/bPnh1TrvZ/WPM+94UrwtiqISM+Gv2DjNWj2+wKwMcH5y+fluLBHq0YZp/D0/pux9yBIgRri
BqFmxvGlX8PNO1e/ifAdR+FxJ8jUVVkzXAKVV999eiBylVj3JgtRzAJ3vcL6TbONJYYkN7NAYc3f
X1K9y3P94aHIKHivdZwXCuCeHPxZup8gkus+26Q3YnQubWNf0tR2dvjKO25AptTKs6kUY/1mcsoS
oYx7hS2zIulrwYNYCnkF2NI0v2AMfHuWHQE+d+WTonChClrmm+vyd7svPYoOrS535CObsZFqObCp
KYmVtosWR+JeyVx2ysJSalQyn7P5FhI8FsFhVqjpaWKE0pGiJp+ZxGk1JtyAQBfeJ/DAZqm2DG3R
ELuneVtsYWMlMtC8cqmYxfgOtfNtsbsdes6nvfJavbjN4GOd+wshj4Q9MP7Q9D1zaalrL7QYchoK
fPjYs7nKTK9tKCFOBFxrDiimOTfiaMCJjKehh3sknOLYTp7NjTeLZmC8LC5RyngKUrPhActn6l84
BrKTJCJHKE7veG+mrWBPMLxsHD91ZZFzbHL2fr/dbU/n4CDyYyxgKejIVb6cuGzqe7UQFCGRXdOo
bOBv5JMLUQ7HrQ31szjzBVfmYX2y14CZLbIwEMG3cbUc59sGut3bnVO6MI0d9m/nhhsS0+BUeVxD
6Y/Cni3Ol2nmGQMys1hAzO7mJeT8TfViKM4Yr0/Tc2h1lHvvOCErKCGu6Ftyl6TLRqi5Tq/kxxZK
6Zq57RELs8XzktnDDwS+WEsug87574fRguAQNoAixQ+7QWlOAp2D9S3fwer/H29aPS5Ji+ayJd58
IuoDChxJjDvUF4AbaMU+q0euCP97toYYy6QQ7YGMNdYOoIbIXIJkHzAGBDZlJLAaQjULwn+dbLIg
7+Tf0aE2r/UVOv0KvJHr0k5J1r6ldHG5/5rXJXNxuOr06dygz7XU/rJ1MPQ2ctDV4aVpSaKaoGvw
8izq/zyTJXcUPVIVoVZ+o/V/wSCSPmZSlTGJxgHPyl4m3Hsymq7NtI3dboFJVEdb7+zW+TkV4eHu
G/L/8pVBqzD9/SXm39ukjWqJQ5g/rFn6T+TWnSmYGuSLZAC/oZWhm7NxggDVt7uKASiLGP+H5WmE
8GIAMq1BNPJhTD2+VwpYNmEH3HsgpMz2yIw3MTWwW/EllD28vLbLcpU9LmlRTzQ6cGSy3NhNpzPd
cW1f9o+XzZt91sv+nDjPv9FwqKGihh5VrONQEoHWvVNPFTn50LErITNjg/dwEK3fF9cfq4/cEuq/
0f+OyKoXYhWIHFi22oyjuyqEmqtvvsLlB/khAoo60hPDsloMs7A1dyn1V1frceY9ROtM0wCJyBW9
GFEXk/Y4B0AzIkOphQZRVYZjqZNtllbWtbY1z+l/PcXjvsIH7SVVPAqdo26NemxJeIY8iVq4QpwT
jXtBOSb+XUL1AU3XuhY29wm1Ei/ApU4vqzgB1USfCSShIsAC1NW31ICBlTQHtTWFn2kT71GmZx1F
HFfXLmjtH345uovu0Omh0g+JvF69pMyDMi+Ckga29f5q7MPDtIPYGvQldE9fR2c/HvCB3DXfIj43
Xib7lKbglcDpIipt8ZyDgDfGHoIiI07GBthOjO5b23THXvFefQAlsfPh2i3TAsiRq4UNxyI8cbTe
OcdUXLzW5f31T9mr8aTFn8y10RaZUnCc6OsLfcwR2/DsBVmPiz1UKVNJq79LXALINRTxEo8sp5eG
xzEsJsmB8Oux4dO/OA9/XN6jNdxplE7aC4d0nJse+NvMiY/AwQ1IZ6xGG3Tj/29KEOwd92hc2TuC
AhnWeVfOfr3PBl8X4e17xRgFqR+B22DDUFGd8n8hlqMqsyj3rRo9Wvj584bChVeq7mgNViNRafbp
4Q13zvbMUjoWmeJ+o/chQ1tFZpsz/tYnmOqsl1FnM6Ywr33T5L7HBTGjgxOfhzAQv7OllM9JeKn+
Lzwh6/CMWZTagy/x8FR8mb+UKFgE9SeyEj8qGgp3FqjkpI0TGU/3YR6gyKhvdoWvO8lmEvE3MUZb
Ht/EXRuSgQjngUqakWHgg2bHOQjQpl76kLpva4bs6x9YyZ4Q3rjuhArHMsfT1TCJ0qJqIBDCXm9I
wg01cL6CJ07BsH2rFDj58CL9UOmMTchpKAQgG02sa0XGkKYjHAl8PsqJrEVsYPTY/dk2Qlk16NRv
UQtNqofLB2AFjpA57va2/EOpqCPJVF4aF9e0yQhMb+l2LnXnxxJeem9hi3QzTPaf4cC2W4l8eSrt
CFjXULSPArgnbcPdT9lSwiBHdVRXMRA6MIIKgMWX7kjUB/mRrmykHv4j4ybHe6skBlWm8ihPPxgG
sgkLVO1ZbBW/EEKe71yWgzDybo1Nonvx1WjEPKHpFQ2MsOExK9grILEPWdvVEvcpi5XIAJHZbk0o
ASwpec+yoA+5Yclofghskzzv4aUb8wB0sIsORh2du9NlwJH2W/PBgm9wv+XFDAon02iWZVRRcKXW
CdbintCON5L1MtPByH/vnA391U/be49DUPGwS+32MYDKes4I/OW4gQczrVgDlH4ugG6SrFOUzm/5
vedd6RxWLQUbYSrJiOXE6mMyAOlt5wIuOuYPZadL1EvIjRA9EWPUlnlIPYpAViqhgGsHha9satkN
ttGiu9M8eaLk7BUiYNueF+Z9KuRXDfsCBjjW6RT2BpJnUJXcB85sdwWRqNHYHzuzowvUuo7DabSg
SUbTaFRu1gMrEx8LeelSSIEQdbkxD3t6PU8YfY7XPnVlzcR8Djn3NqTD5NdzKtd7MgqBORmg4utZ
sgwkewIevCEtZeLt985EgCBr9TU136kzEXmOTcWgnUvwJK3IWCXsad4xR49ueoBfcLteC1q/GrRL
azlhQ4kcP8nObCvu9DAYJH964atVzDOHcv+g5DTb/Nd0UW92hYntua35OkdA4Ldx8IaI8iq0UbcA
/70CPVa74uRYx8VrIBn7fXP2FUNeaFs8BQNmvvHlZSZV2nles+3ayOMhUo9IuLnQFttjIqmkd+kQ
8iHWhY9p4bXK+0PsL/zgmI46h9SmV2YYvs1MFgG3zx3dg6x57nPlmRvrl5oBjXVcmDdkWCLMSNfl
LW2OtjoZcPbS2NRENkHdxxelLokGQ6NPeyzOpuzU6pV0YVb9Fo2zKVgEnYmwoCqIHzW44I2eH53k
ogLUcg3ALS0o7nsSR1KmtbtA+EMlCTNHoMdCUYe8h0BbLGArPcVdEabLNYi1igjy9gAUY3es+AgS
ZhRJNWXm9GEUhz+VSrGE2oMC0FPOWz4xWTeXsRTIFfIUEvHzVxNMvVqa9xBAbdmXd8+/ydNQCN+6
YOfg7KHg0k4WZqHc7VLC6Q0nXPVCrM32XxQdcc2/sivSGvnSSqmN0X3oiNGMC4LUjTtr73ASv1ol
nHEaT1wqjQF0Rm70q743KMRQn2cT/+I0kd6XDd7RTWBkoB0TfvYKa9DiVn6uk0cHS8oTiuP2p7zA
EhPGkeJDChxFiaTBLhejALZHApwlAxEJOoXNPraXAhYrlncGb3JrBYKPA2dnmJe0AmutmR6461s2
PF8hqBE1Vz7rAt75DLkczM8P1iFYeh+vlC//A+9Qw7CsgLb2kXa1+o3hL/jj2ZZhYfBtwk87vIAU
vZB1YPU4p9zTogX9Z3v3+edSkTTtOyZKBUt+RgeiZSpDl4rbln8M+6ftOcTh/yda7YI05oMuFKew
ondd+K6xIvYPnJf9bvJv9BEG7DiE9sn4ULoX0HXI0LkKb8eBW2yZYS05WVFsAaEnttq5Nz9N5yRk
eNAeWZeGpiipuVvR+Z/fWtE8CiC5cRiGzbY3YBmIfOlTv2Go6VajXIN4PvtFboNEHILUDjJG14Kd
4VnM6c7qT4Zt3rsSwjNfnvSgYXBIVswaws3EtXf6dypnvdX4Xpj79hSyfmim9Si7l4azYDHUaAo4
AtHAcDxb+tVM3b9imj34lE/nR9BI+YEUaUgyAlm5kXxdviX5QsxajcFBYg7CX6QSbKhdLpMCzD1p
sP1gtyskU1xLdKJsvZpjcI4KngAs/UVSNarEtDemcy6LljULrKLo31uveDeT76pERBhVqTODnVR6
LpQZl0LGi+yx7rfXnaB7eFii8Ew9dDBx0nhCk+5CdRBjM3vAWg8LZgPJ+GqQq0nGzi+9t1lwWWwo
lUDH1m1W5JAhByc0QvTrHkUNuNLsyPegEi4sdpW9G01m+n3Y7miXVmdZDp+gfxHsFi10+xgwOkjX
tA5PLse4QWqD/LoU9gma1H4dTCGQQ/hw4VO8VUil6e5qhmy1oRM9k4rPGRwLZaWYO2sfIZz+U10r
gRt2CutZN1VNkeSUS/OjErhHZroNb5SpzjAlLQDo0y5v5Br1FkT8ijupzS7s2OdDV+tp//KKA9Bq
Sakj4AoOvwql25Ug5zb89vCmAImw1b0L649dO2JlNSglEj7MP7OF7gwL3THP7LaAsVpcj7H/D1DZ
XSme+0Ij1eGOp/3m3BouyuPkKeC7uq3c8cCxky7IFCxsIuh59wE2dyzcamZ/K9OSWU69Wkr98dbi
wzYSavKDf8hZJ2JXUd+UuJ/CILWdFROjhUlEE2wu5cypFhsg7FLcbBe9IKF98B7GBBH6ecaUq3Nt
gTLMIcgwC3BIM0M7Dk/xhBWLTg80eR3unhDEKoexbib+2fkJ/c6pF0z3jtSeNJoNOXVosCyuDpZp
hBsZJxSFDKgXW7KET/zNwpty7Fsh08i3SZrP90lOmUmFj2mlMg/WPEMa/m1T5EY0a+Z0uneZxuIg
HnWKWeqcnW9tSyPcI4YJzcEl11KPl3n72RUlsRfXH6CQk79x7OB+tZBg0TnPnJvtgJaowT5utN9A
AshsrdfYw8WWpirhvK8uQdk3oiRtTQVHxTmR1+4cD4TihxXZRurEhd92/37v90TIzzp86dg0rr1j
QnOxKCNPoKuWV4WM0KPx8IK4o5xv9fqaTjpxYOaTQZvGu7nn5RFnB+R0zYoCogEEmYP22nnuXRuF
7SGLz+kXdLXgibqFI2S5vfKkW6hsM+Gf7vBjkhVcOhKPopeb3PgIsfJoVd4swGnXqYY1EPzkzFBg
RaP2XvJj0y0JG3I59zb5rbgHVLetJJQD1wIxbDsnMmyYGluwSwrQiO59+0512PrJpCVdVF6hctD2
LaLW3Xhox97orlReKalN7F2Y8Uom897fKjcuF5Ha6g4fItRKwAkjPHKfdbSwN462sxaA10nVKAJ2
kMhKRPmsC3q1g1eSOxQ80nodwO3Hi7002ePnr0L+QShs4Zer6wfk+vpHTdynzVSXyf02V/IQboot
usf5gnh/lMTsdZA9VmKve9qxbFcq9q5csQOoNOPscNKyuDeYvd9I1llZqfEnArF2JupewHolfbL3
gKvhwoVLfEgLagvLDXRkar3aT8rtinHJ3sJ87ksHhKzFDKW2wn+eF1na4xaerI9KiFRo8qU2T0Nd
+RP67xVyiX9Dd/ikSHscXzge40S/M5cYbUfV9bzQbrcaEBR/RSPR6CxozvZyLXGwhCWZwgtZk1tD
Hd/8k4FmfP0Y/8p5JgG2jtw/c6l8TzaHW/oSTKH7SBtDebpNWpQHUB3ykiACP9z2k/nWdSKVYDVD
TC37nygRAI5MFSrls910aaiGxSnOYSA/UpjFvaYm82wTIttSoCXpqsa3OVD47b5438tx/fyezej7
11m6/RiW3IA8JssBiaYbIrbCyfccgu9TUTaEwWPmsqErZIVar5c0UP5bDkaAkmz51+Flg1yd+H6F
eN6JCXbluw2U7C2G21ezb5xVKrRgwlhA6AHnrB7zrUjEPIFMx3ggpwBk18725Ff0NSRZePsG/Zqs
YLP/gUVSUO6JB7F7Y6xg5EO5g09nxZa2XNOLOLrkzNe6tdSthsXFP1bqPv1kpqiJcNQgNYta46CB
KoCn6KSacgisUte6btIMirQWQ/G/caHxztDQi1PYU1L9YDbPRSkd3YTAPH33wCBJ3Ch15L8cjzNf
sdXxlnRdSN6gyi3twJl3zhLdUnQiksNNC8NJktN+At2Kc1R//UzDc88dWV4XsYLeh1VfLltNS7lL
zfuH7D9JPtxNmoLY2ZrhkrZ1TNBbYTXxyHOp2gFDOKKmtGafwOoLXTteapekW/n6Z8uxo5VRxTb2
7JBMuvPbcwAymiMtiWiqZGWinQE9GhJciW6hKwc1L/GoNJHOE2T4Rs97N94AoDSpDGcedHCCFkxk
plrTVs4OdxAPXf7VVTnjFkSwo1Voi9C/WAPpNNcWOy3cKgYoJMLHusLNelV3ThcPNwXZNWDMJ05k
LqWKQRM65DN242p5NlXfP1CiwXLW7jA+WcA2baB7/cD2RsY8vwHGtWj1r6O9Z9NUcKpzkBD+uPlR
eb1pKiACYyAl6GCDLeaS1iHUEdtteiirO5dtSepOthvmkCxjmliZomNW3IAyIRR9NiGIZhj280Ow
3osrwyk7KI4pdqXDFPVPuYmqXmhz3201TXFdmuqeV0f+h9OviiGRDTE1gMPzLYvaXXgq9/Tq+euc
czig6zqLlens8niDwGF2c7r7kdlyYRth4w3n1KzqL8cZdQ6nzCCbFUSEyaIhsfrvX/2b5VKYAngK
Pa7Exc+zGowRRBjB8nB3Qj3n8LsFpV9JBSzSrOAIa9DTnB0XYOY8dfOjn2eAaHA57USE6XTSh2OS
6q386QUhBelA69+8d8COWH2ab02fqvH36MQtL/FTHWPhjITY98dFQwXDtr8RVK1UQj8GV3lOyVMP
r8ZpZ1FsZgov6qn4NAO6MuT28cadAzrDkpmtONoEidv1iWQLI4wUxZIJbNL6GsKkIPkXQ81frz0E
UI+TgHYysFomtY+jqRk40x3DpAtINxDH9cqqTP/xvKRv16dciwYCe5w2mOtj5S3ZkTL3H2dRkEYa
QxgUfyJbB96Zkx/iVJSBFPwFTg8fvfXM7WjikcIbag7cp3S5SoRv8UaTDSuy5ZGi/1I0alnY4rxu
38nEM8UJE7zRyEQhv++pEFQlRH6RdyocNF24aZQHVn3LqOibgrdQgcwpSmGNu7hsCJW2w5xVNStG
0zpPUSKkQhXpnUS/aqlS/irjn9ScJpsy4ahKxZXJfY7zvgg/HqZt7rqdbcMEyrRwjETlD0Ec+oAY
Taxxrkbwjfxs+AY/mF1c07BLpFxTxx/zuWnIR2ejVJqqKjGXOsoSDykKHnxxTnlo9T3998t91To9
Vi6OJNuzssoRTz3TVUJmzUhof0l19wuYb0KC24b3yQNo3SpwIh9x2xn6Yz3k9iage96rPIn65R8k
xrgmwqWRdBUv1ZpyGVgH05kAudh5rpvlE6Q/voEtbwZvPfhU+H5GnIAPycgqNL3DwoDG9dDWMYla
tXCdb3rOcUvQtELUFJoJB8YcGxf89oSK1SpvwIRChV4y8C2N4nTC6zWIE5uZ/VkbJKKsCFTE7LfC
4DH03/H53Jle5tEG0AZLQ/DXOfUrFCKB3T2jz6K54V/ecrjxnE/s7xwsv6ZzpSUtpz+CJJUtU5s5
0zat9yQ3TJE1uySj2324/3ocUWh0nninym0Ig3wG/uzc3Q4crql8Z6A8HLb93VaR34CZzqndJ4My
4sf1IRqGVee5ir/dJn1AVYNMupUWayuj/I47vgakM5i5lXRCLjmz+w4dgSm7G0PAOU04WnisVhv7
mbfG/cmgq0KxSGZC7MQt8NvMELArI0pLYyOvSeG9yMUsU5Vm1uiDimBg+U34bz19PWFvDskvdjNL
8oLA1cEd29jZfQOqo++AiuLdXOlMK6LSSkRQig1TszgYpcTZTqr334j3hbxOwgFLLlc3TpzXzWPy
JWHPoSRktL0ZcNLVCKNCBuCQNjalnqh3OeaKJ/XdPSIXRssq+M7Ouzdqunl5iWpK38J9FPWF5eGU
aDfsddE2spBQoKlWoE8U3xQftG0Y3cCHHDtjj/1utSlW9x6tgxiinbIFMprTtHbJsCg3HPMJfv8Z
gIk0rHQ1z4N/61nkyyLWmVvwow/qyZ4O6Ec12J96Vn7XcNhVhunOr5YJnBWvGat0dM4R7NcE1QqA
9wRHCNoKVC7kxvSkrTSkyK1KmJPKuEoLLP7BR+3TDddkm17BhwN3yyslk0bdJJxpwEPDKNeeiV5G
ksiDwG5EktSE5/W+MEXkvvJBuXrBS8DYD35KmKFz1nK3Y0pmtYyzoF7/U8baz5/5AYWzos0PwpiD
9ZQy/NugjERpE6Pd3kaH01TZcCVPXWo0UmMK1x1J0LNNREGUzsk3JklBQdYXVJ6uKH/myzCc01mS
frx9oCnuGCmK1eeaI9+ZoUSoO/N0U9tvlWwywaqr+xw6wIoabCFrYR2NwqViGrTIWDz1XT4pzgf/
T1+0knC+KtEWkhpuOjqDw9UJENLxnHs6ts0aL3mcPsnHpBUb90AcUAiH4E2h4h43XnjY44IcSSdK
KIqMVlFx1GPU1CDqPxSCDTiKSR4GQQBXpj+uMN5kbo7C+dlLtw+8UMD2d8lcQwJ/XBluDge0fEoS
4PCQWgqWV7mF57r4GYm6/Zl+DyT93XoE+gKKionCZn/VCh0By3hsNJpxQ070qZsPpG6YeJeL87Ap
KKsUzJ+fqzromdV1vVz5Dt4Qi2JciuQ09FCZR3fewsELZBHxhsLr58Q5BO380ug+QUi2gEagz9av
uoNVYZ3dW/F2+0P6GKddSWvysHW2k4eW/upCLMlyK2xoO3GaJh0ERF/KRFmv/9ATVNeLO/9WB6ZV
j8xaKfKCr5bE5DfFg9hGDWoSfvO6PnuFfUg3JZOwBilJQQ+ojvUQJbAR1WU4ujwtwTpfegr7Q0Lz
iVVCKB4r6bI8o2n6s0/+9WbE9IfSHcuiP7xMDeiGDCxybIEI0yLGugPYPjKQlN8CTWF3Ss+8KdSJ
FDWB24+Xj4aMZHXdsCVwtuXVhdnjB8GbtJDtVIRltmPOguufiOJr0d+T2bhvEQDTeL8DRE+yVvId
GpKfkJazeSgiQ5vsgRMzc8/kFEPMXfkfMiTqVUuuPPAlDykxNiYPYLAak+nDpPPsC50hGn7XZrv3
HVAqGYaEQ4KfVp3f3ECxiAjLieFwKqvz74cXhPLKSWod0ry859g78RyI9vKFzkZE2FKkQhCTEZ6b
xvoCfPSbBeK3RcW73jHkMps0R+Ij6xuUw9T0ejCvUyg/pdS1v5Lmx4FkT29cUId4QoET5DWGvSgY
d+vA2SWZyjn2OjLfeORE8/JVbYR2vLWB8pPR/qtAd1exmekHHvGeL/zFWRbLmB7ZNcnsr+59VA6d
GRF5NxX7rGK8If7BwqlLA4z3Bh3Y+YB3mhJvFUB5gNqRzo3aGnrCvpfZn8R4StxPfojIt5eN8o7S
7bhu/jc/Vfx+p3Yrt5O0b5Mk9bSDlvTuNCg8KC0M8LKX0qldGeMtpa99uj4EfwEsfqmmrBH6D2p5
S8soLQHNUvjNypzLAHbegtjs+F1MIIwEqxNSVdoYOAZ9adYBSE5G+XvmoYoguUpNwvNf8cdoc9CB
9o/+Nl5TXBRLxveRg8DoZhemPGw8LDHfuUcwR7gRzLZesZ5cRvqlfZ55IygqAHHrMZVZxTRHjNFT
87Qm0RkEV6U9JxaGxMYtJwzw1kcdk7eixPhZ7kUaFgHYdVBcAwbDDkXqIS3D994p/zE2ezc1fVLe
fM6GaHjBAUB2sziaI6A5bFFy7BKnvBQxRCxjP9bb5GqiSewcxT4Wk8/OYcAoqquDbuMCE2AnUUVW
XbmuweFFGPDQLtUqu7c9kSPmIwgjZyv5WWULOgLTFcELq42m9iv4Nc+VPM6Z2sfqEHNPM/tQ0gG2
hxrFZEpIQ52C0cWFDYS/b4d2h+1ETU16Di4kiHIEB9EawBq2DUXxYXWZ+o77058HQJrwNPLoQnXm
Xi1VvBkekpwjmXisYP7CqfhCUCmVMDI8Msaf+r1PIghVZbq7OtCrnYAezCkdr/0QRLsIExUSHEYk
0wD0Hzh2Au7tEb4W0I/bINsKTZLrbLYQ+GUyTY3pDFjR58rNhM2DUQ12wrVc46Tx7zNQuuQB/EDC
tmDp9+RPvsI5LaZSdFqTMjiQYtOXvzVakzOjeic6+u8bk3p+vpb3yMTvggBW0a++CCjGiDdzfsWp
VFwjd6VYF2W6DOOMlV+AbHb2ZdBbfzoVkj6zRDGF1nvOTQJi0xQtjV+jyirdqDyzkP7rDVimDdcZ
cPT0wYExbmL46QdHcyyAqNNEjBTXHSogXikzsmmlQAe30n25MFTErPVz5xopOn6Fhoyw8qkGoUMg
bKe0voC7jgMT1YGj7O+BTZnEYfvC8/Bqq0ZEogNPO5ispBTK3jUt72cYmbYdfSn0wE6r4JmC51Wt
XO0mx37Zn1ekJsfAjIJu5eG6J+ZsBtqMaiIs8zQ4KpmHr00SjgQCIFippWJkMkhwZW4+j2D9J72B
+9V7dM3xGQ5zO/QqH8yWXmV/lPYNQyApH15DLPxX3oBeNqWUEbDEW9fh2loheF1eSzMqpcoPfpFU
80NDlkjfYSgPz1vGpyOnZ1qAyvI+pJ5Ux/Whreu3ABoygCtL5Onn7oN/NbZwKxifGpcBo98q5H6P
bTJvT0olpOZvEeToq0xTMh6C4YM5TLQb4X51XoaH3MXLGwcSt34Kmb4Y3IpxcDin/vsGFbGg2jdQ
2M71rbx+kevoeok1BTSDSOu4PRVbs6ufqX+C0xaMMI1ooyuqh0oCvmfHFOPWimVwEQwmXwGuvNro
BrtEPuMMzr8kEqRxeutaPlXXxNUDCjCoknBBpYYwb8lKrIKRdvg0R2qcRCg+E/ErDvDiqdN2oAD+
e7pzvruy8zovJsqxbZOGlj4ekCmKgApmNhgaC349dB7FX5jaAN6yzqekpp6HO44T/EQ6ZKZ1vPAA
viWq2WvnjK7vma/57cOjdd7o8XeyCPp0+trkynEgfgCpXguCugVtHbCGSCh49fa0lkVMAAuUtUvl
y2CfMY90iFsrmOEMJYMSiG8tTDmAgoKwEGyr1SrN3jw/Mjm6siYtcfAR7VogcCLPtDX1yg0/w4d1
uySmH69TyRTGfHUx1mWj975/dQz8JXMDH7/NoDlN0uhb8iMgH9J1+Wbl+DTUReYLmGTImLnJO+GB
AT4RJ/yB6cKliEAL/CD9meHeQsMuvRhgSKqbYdfsRoSN42q7mazRnSeJIphmqDkeknxbPx7xZy+H
3CXjGhV7GSx8qdVfdxhEWriRWVO5O9tAkkXoqyn8m68htOD11AXYrk42UsicCudBThKgpFgDIVrE
K874WlEMUoBgWVVUDJjkhElsXBWz8JsofmkGXzIAKITQQZTsOeV9iWKPAquRuzXM0LYFB77k6Md3
GGuBC5lIq7p9EbtonayyP3zKRR5NIMLe/jf3buRceVAvt4AcnLTwE7Qo7g+9F+89M/XoQXdgbHYs
IuHEQ9xIj6NlEtHYUqm3Kn1hTMKkT4hTf6LJVB0TuocMD4T/15pC/iykHCjtUQuP45RnOijX2NCw
+CX+PoqBy+B2LHHUh8FBQyyXwuzeZSByG1ni15jY7YvJ95sQZhzaunwhh1EDweBlZv1YeqpHPpjs
y7NqgNh+hkWEMhxVZLJQOd0lp3Txg5ZcbUmmlH272vvpolDclii2tJ/zhdJjcm6tKMzPgCNIyv9t
8TQ4dlcl45uNUnLMyjaYh2laJvakwGVhxiT9MF2ff5qDY0CagBGoix9fJ3tXuJYr5uJDTxwshMxS
KPddaNkzzZZhNNT6luTrTarsLNKJvJzjMpaSOZ+LmQbgf/IucnSeYnSpIPDNz6NBjhKckFFiF4cK
Kkv+pITDDFvni4sC5gM7tHy22chOg6E9MO53lBQnO+1Q8CAOxhKSYQJpzmYaFRUdZQb8iSrhM1LC
WuHQTA28NAoyRVra6KkZ34LCj93tugmvoNhL/Z7kdGZTc1e9rRA1IF+w1qOOeE/sycEvIbuWibul
m/YdRDxkaMtqusjSnWWB0Ef1zyF3H5RVmQ7YQRf6B+cKt80msV5Wz21eplXNBfqBM0xGZbZ6Pd3h
/CGyOGkxMt6JtfuYt6dCa2fbqbVvfBRRy28in+m2CbIdjMWpmCgQ5NbhLyeigxsOoSCrOuWhhIw9
m+499P1VSY/CRcL1ETw7Hd2yW2kOXaTLz0Oo4ZWdmA1Pe9yhsSfO+T3DpimyayoeCCdRYAiZUT4z
y3G1SuS4sWUBIXDWK/Jjml8U6oIHOFhX0ukeSNo32lf7Wjw1jW8mIOrpJKNktpbIynQaoHpvlPRg
4wzv+yJTetT94o1wblChYmj1zALcVz/i+7+6V8ZJSyoMDbNsKugerFmWHjcXZ//+cHaPGhCRxeZM
MaUuY1VsE/oSpb3QfFi1cqqEOmfX0t3X+RkD53lupLcEJDrSmNMhN8HP00dONcWfLmdSDQBSuQL2
I4NaGtwrkhqhn9kubyncSBlvOfPsgNr4H0n4VG3Sbm4MpNOl7BveLx9f9LiisQ2yNBCpHLh+whTO
Yw37DR7FV21M3gbIKHNvhMbVXcuc/rWiN27NTcILJkDMvGRW4AlFQ/r4/UBeWrqD1DQTQUm4hBCe
tcWL8p0yOssPsDYrthDSUJUAmYDzqa77Pszda9UjJ1dYf3ghycNhgK+b37kwB9aHf/+Kqmfav+z5
pipznhs1fdExuB1z4OO5QCRFLdItt4QoOTjFZCaqweHLrwxrh07VMzYfBdQmwjkAkxmqmc5Vnssr
gIPbwSED8P1t4vRG9w5GZdht0aTHyh1yQDn/h5V2aZeL7PQ2y56Ii4tJERJzdbmosT/Vxe4IunZH
f/s27oRxRyg+PWp38bImwuhlh861lOQBq/yvxKePMrXry+Qy5Wyy6nGwcIsqEDnHgmyDtD6NatMJ
YgRZj0XEGXchwLBYTdsQwrtB2uje263ZkZtRdKNMSh3lV/wfJZnErD/QO/KU4u1ZkJr8P7GlLSLg
2wEziLWxP9JR2XGy4826fiqNtwwN9MsQvQ09VyEK4BEyNv78ZjII0ISIRFFTd3otjMFm5ezok3f8
r8zz4yQnyeAXEhB+6nkv1KaT79WjPe/Xb1rWzXXcw6DlXgJnXcIdU8GuxQ9IdohQ/YkfvgSo1yg8
1KFpUUKfoWLSL+Delu5Wx2BeEF25ysHfnPuV+AB1IqedcM9p+Zr1G7sjwLNbspkPb4WTHlFIWKAr
qWA0l15QUPJr+Nj+FsWk/BBAJ8/hqo79aTanSkLePnBPHYccnOC3NKlCiSeqPBZZiDRA4q8vIwFR
z9gTop4jI+23R++9m3VnXl6uL7DjrSSd662rS5TUeg9q/2gSZEQ8PdFzO2bi8S3/PJdVdfH32lsC
hb7vYQCP0d7OmiKkoBVd7oPVj9bkTzUnKbnbrucdN6sa8qMWMQ/xmYy0PqF7n6UbqGdk65v3Dzu5
RZuiZ3pYKfwEUgzRZXDlHcT6eH2JucXwglRnlAoW4HX6fStRDW4gbW1QitvQ9qr+LaewN2Pq+fF/
roas+HL+fE2MZ29Kk59PiHvgu65jNwgi7cU7tqHBoUzBhO+Dooe7lv3DQFA/+HxWAj/zq29MufN4
TdOBUqZov1HxbweCUbrNM5D6h1LR38czyvNI935aHucRmiicpxSPYce684yFwz5xVJGjnxFq6trc
Ij5MIuoXLZISilxHi4TFmajaJ7vjjVJGft9KPDszVz+5iAsVgOEsEmoEvQKAZl2aIHMgEqFuIwaE
4L1eJs3HhKEt77CKkP1/7F/2tN/WTbUDFBmhXYbOss+mfSkXxmZkVa4rKADhZd9Ux4cI/XE3oC72
Gx+E3LkHGBaSaotILYfjHgvZDaBtdxGshGsOyHWsYcoSHVtkgpJ3GouES8am0DZGTGTB7T++L7cT
mfIuZov9RrNmcnOB1LUYRjl8/MtbPONkZWiAcG3opYCXPKpcLxQWvwLYvqx1pSaPun0HDMcJI1sI
UxmLLylRDw06PuXOxM+fZ1JHACxV2hTW4DIRQtI3Y1qABOl+/AyxlK/V5a6z3iJzbJnGHWDKOKDQ
9222awA7IIiA8kqoESCug9jb3ewG4ZQSkpj1QIXICShWGsH+EODvBlq66jRBTX4CjHHmu3dQ8Dl/
NmWghz57SaLHPuC5ZLszFiEVPzvZtdzmVLki3FnMcCFWr4v9zT4dYAv2MGcD0pMJmr+EzXjSKvo2
PpazS4l/fAjRDdcsbcqq/3g5VtYU6yNgsORLqeshTtxfssthYHzzsGgOSTDRIW+tUxCoclLMjttT
u1p6VguuO+AAQgibYdWXr77eykqPPODXM1WfwtomLj9cGZ7fbwtgsxS8mYtEK61yH5F3k0ektzO0
xEbBu5Z8x5hO/DbMPsSYcZeHpi84s43Y+KkMl24fNDvSahYN0kFFBoH0Cwkx3tj9j4hW2TPusxyg
+KRuyJQmsmRQ90Bjz+iPLGnKm98DcxjZ+iWVgtV/RW709TgqQTmPwZKqFeAOwyUQs2fh2REmYxqc
NLaog8xpxLI/binWwt+CIOSx4EQvPTduyz1VNtnfAUaOAyBx5Gv7pD4zhucmQa/MIPFxYpYLkWul
ky4718s1P8q46a/uZ1dOIPQTzkPA8QWjde2udZ1y4H23wYKUrTvDqqGHE0tAWHBLXL5RtgCRe5jA
sPF9jdxbxetiW1CNX+GVvWyBcjXN1ZcHmqIyBC6pDZrdYJnZEIvDPuH/Y9bTDpLfmOhs0nwXo+Ex
TEIHpKJo46HP+LIA6gITjEZBHa4ewYK3nfrYUfAjBpFVXkRmZGSOq9BbtISE/PwWoOBJGb3kD84z
cYTblQU2uO48IpP7lXPEN0gX9KHYz0/LtThN3QVIq2aZJ8HBAcQhmfVj3hu+SBHjTTzUZV/mBbyE
puS5e1G9jSJ2/3oK2pm+JojwTHudN3B0bbR4lxilnuEC3DPBuqyfmGM2gYaumvLqSommCOUPXUkP
hGKiVS9qiSRi6O3x7PJtPmZG4EKGrTtQeduwAiJ4BvhGlTM2aLBeuCwKPCdJCyhnN4SGjiSn/UAI
b9m+4Lb4ZvnFD0gqNJwTRh3O3Ymm2DBPJPUxd3iZGG70GdU5xcwVuomtFzNL1CjoHHGmaO6bteed
4+5vQiziFhkEmzCNjvqNA5hhJSm4+TAKmjmTPDYUpH/aIpfxNvrt17EtqIB7FIsEZtkXJML/9UrD
+bJp+42km+O8mJ/iSuUD68cPm+5LaB7so17E4iC5g+mhLgt8dAasWOhEjEHRdqZ0AIIKHuvW3CQJ
zTuhwAzvdbRbg58JfP+XJCf6IRjCiWSGC8rDqUiny8838iHFm3XYf6yNWLGweM61a9gcl7Z0HfJw
Qx0IJ0vCisBzI8YYwnvmg93p4cFa+G+a1xpbnZRFzkQ+s+Js09DGihCIFDvUZ406X7/jK2QwwTts
9etFVSxNETmbdzzAzLQZfOi+cnfx2KjOAmtIHvqggn7KZDF7GiBs3kAaxeEDVP9otOBpdrEQJEOS
PDM+BKqadJIQzz9KsTVwPbtVW2mJ7jle9KRnzJUgCEgyiVYgmVfQ3UioOubD2FEppvwRtVoptapd
mcS5K1D5x/YdbKJhD730w8fuQk0fT5h2ePX6DhOSMpmwiUCj1DmeOCT1jVN9753lUOLmSZwLQqD2
fl2xPx4/VKpMFGyfeNKgOjzmKJyGIe66n91R/5fK3qWupMEtSZyxyCyJLMkauG0NvVMAScI83G+W
Iu6HApzKIfIo4OEnV960CmNWDOntg85fs8bAipxecnQ/z1FVURoZXf/sJX+yNBSX8DIPXUyTct31
hR5ZRW46zz2IB8avXsbzC/6o0NJdp0HTtTEc6p8MVDwH7R1q9gWRPpli6b75EMCUBzlZjK+hDNwd
tgZVLcClM1anYEglkkWS5pRVi13PvwBxTMD9ES0Qb7TOGbTfza2KCu1eJDvqDrz55e2QJTB9mL+Y
t8ZLgdIUtZHV7p56nVJM4j6XQilCRI5JTfWdUaiOpvR0n88wTV1akCz6EPBbCOANgygLwx13+b0D
foDo0V8qwvejmBKpititiTn+Aqxp5wNUmhpeVRyzMRdPG6PHTpP0edK23NWm8bgMW6B60izgCv1o
LLyvyG9igcX51bQIzRUmlyQHiiNNfQvYFYtoTL9iNBMTJAzgqej2m/+9dwceplMTCO380iiYP5A2
pmgW5KZ8dVVnf3GAvSKBBih4w7ClHlJA7QI6/f6UanpCP5wD+rsI+FB//6n7rMtA6Fk/C8Hz0hAB
+CtY9CYPptSRQKXnPLPUmM2Q4lXnEH3nqYEEjdVS+0mXnes9a82mr6JnlNtovo1ZUDtubpHyMnx8
6W1n0n2dIZebskPL1QTQiPr4hhesWDRBA/fg2wExjHbu2dluEiX+MCZk32NJuRABOaGZDnLJPXFB
ydL3Bd28d3XouqEcvm99Snsa8+oLUm5N4ksLI1yLDXRJZ2RFkIacb5ilXHm/mmklwYikI2LMvJZU
+aRo+8qfnJTFUuFnouvMolvU3iBAdMo7c49o6ZwRc3ysbspWyBW+dAA+xdkiOVVJv71EC91ZMdNY
zwBqx7WrWR9oOQdENfPEC/86PqlVRgrNj5yMwqFvS537WegQ0/5/TsxlpwyicCUVme+WJuO4Imml
W6WWT4TG4tos66j5ou29UK8k8Y1sV71H0bU1mfj0gMCrDtQS/NKehKN4t04BJl/A5Y5L4A4EYEmV
GsjN+Dr2SEg9rSvi1YElvbfFEIEPzuAQebRdmrdNWvVlLUgh6pc3rHAQHzh7qqr2ue9Q/rHnOkUk
/xPBtqA5o+KNt7yAa/CFiZKd/NRrhJ2q+rOP8aSCdNYm75B1X+C9eX447ZFT707GLnIOygIxzR5F
kRmcEpmKyiqSejRiA+wS7qWnH8NUoGsf6bcdfK+CJzRICOWT/TmQehta57lG5QoFpz9er4A7BUcK
OAsHNYfWmd1SQiMfhxOijSBgZF06s47FFvwYqXbbSICoO8pJmkSufXGmqEpoMMZBLmJyS12t7Vfb
E+5f8CWjULTdb0IcBIQqvqsj8ETLmeYLNeHhp5SxsEAgkEsx3KWwmF1HWfMQHAOL4gwt6euqt1rY
PRmNVQ3GYhofAmyP4+lpyooS8f1h2vYlmyAXdZYdIw+V10pwbOj1Gx/uM8IUPoEsyBEa78DRFOsK
B5pTHd+GFbofZdaSCu08Nfaf76P6uW/6NRrjt7RK09ZknTT9ModhgVTzbXWNIi0hA9eWUoWlOeVN
2VqJ50M938eUq/1bY9quDqlM6JqpWrRP0pw41824v10nuFHMoNZt74NjVyg0ee2+W7rEEd3wv4Os
9RqDZKFJgUHVp7jqYsuyqp9ncMfenrdshMQZ1g9uPgklgh5RVZaHZ1KoZ0a0SfW6ZrDU/goJam19
SthRRWBhbcyHrhdO/q1PfIEb4GtECWQkUgD8VG3U+R3Bn0MewvtXuDQ6c/sNcWZs7P6v6kk8T2a1
crM2Qo6tAP03etloKPoiq77Kwh1MVxSK3MmrEikXlcG6pJxBV/SL7OlgstCqlznnoV0vmveTWtG9
SdicY9D0elXzYQmSgbkuov/zDqsV23W34u8CatS9FPCuolRnRA5Dl/svX7hw2dIlb/MKjKlmS4EE
+BDgiXhHWqtR3cRTWqtA5yBEw2eOvgdHdhP3x2qQpjy6wt+qKIXOQ6SgXP6Ia3pq5rQRE9RiaTa9
QcPBJ2wGNlkAk1w0F06GfeoXm9eL//vlqnwKM+qGFKtPDtC0jCyRoQW5ugPSfnYsetYr4T6VY8HH
US8Ztcj30ru1mU4Y4zFn7sFu7Yx5nFPAdRaGquuD/qvjabWYJDvANpUNiUdy/qNMbG5v8+X087F7
uJBVBBSa0Ggqa13+n0xH3rDsgtdsux2e5tYAx1C4rm8XX5GP/QWKLEgRlEA8865QM6iNRBQPBD23
ax745E/RSdkDHpd/YFN4Hr/BxsmaglFy+CYqvNJz2haYwxJRMLXRqG+MxjDGzjqxW8d+q3AGsQpQ
WXDnhvTTMsImgRlN5sp/AKmIJbK25FtWWfdvTSOJwgVytW9JKo4eVMnpZaeClFKwV56iO4tlrffD
GTd+BAPw7TNTDtETvaUj4l/9/9Iq5nur4cekasnve4S0WZmAl4IDOevOHYT7CZzFqCO3Ai62auax
wQ1G6inlhK+r21Hjw0Dty/r113HS5CuBHvEQy7y41iCANATeW8iaig0OUaF3de2Z4aBGbRK1CEBm
nNFFt7hCOyT1ekzJS+qNodhyXRqKWGOFAVjAUhZWa6WIrogxRD0YIqXe7pdekUAidQcM+UaL0EFj
mk/Y0QVYJub91+E1y7FSRcI7yOgNw0l3wLdAEMRmKJndmUEUX79fqHZZHLpwR93XpbrBKwC9UyOA
YC+zXlWjAMZwL6CXvTFEjOUn7SkjS50Qm23yvdGK2gYOSJB3rm650pgHhbxpXTq6KrHyCgmce5hJ
vyBcU25LV/u9DidGgDGJ4NfKRyjH9pbuPzTeQhhB9YzuxAGLtJpc8RCbkC9mEAjNFkZgA/dAaC2a
3fm0Fk61k/b+FBFz79DdCYXtNJC+QPWR9RUaH3ofD0lrlaOMHUw1GRlDvd7PvslvNmCQny2T9lPI
IZqhDa6HLq1jO3qtVtn/8p44Gr5H+yQUfECNBsJzHUckTAxZbZr039rtHBgWzh5pgiD2J1KeYl6G
OK73Ht6Kx6WrJIrbnicXtIriAnylAW3vHpx5InnwdgWGsZaCqqpF4jOyy0QUA3l9NB/EfJc0Fa9R
nbg+5rmEcI/chojCU/3Yqi6CP1laa1hxDZ+HUK01npeLkeZtOQknqn7YhYmvWxb2V40Xao2p0H8D
GTmyAZRzrpcnAf4+5keDBr1BS0zyDrB0Ofle3+hBinf6QRUF4LCh0Sbvq9UsGQ7HV4BeiTpuXHoG
fxEa45+9MB7ujSJ64RxEbE8XkMAyI2VPHxeRMP0SWQY1BuUbD+X3cDYGoXoHgRncvC16SobaMFaI
S1G7/xCrnZZejmk4HW1B3J7CNkH+Ly+NH9OAJ4UxHIJzM9gnQHZZevMNGvQMd6zp0NSNAAiKitf+
2db9w/OwJe8TJBt/mu4sXr+7qxI34+OhS1KqDMTrawRtFDYvn9y6WIJm1YLzPHUCwIGe9T/HA0QW
d4FgH1RUUHPQ/7LnkV6AR6qtcuCljyzCPPX3K+5cHWrRfCcfrxmAnasExqruJ7VDVlvUdm0/VpkN
PjVaL4JjCovJ+QCbfUzfgfJVGD74QySh2ywDyEH+K/BsmZhqmS/MlgShcGt+u0P5j/OpThgQ7zSN
ztzGRzEXGZPwZu3SjuYmdEDFMgjcui3Oq/eNBk2ZkKIQYYTUN+bbwSb2NHhoT2fs2eRanP+Wpz0S
PKexRfrVcjPseEe38Koarcf6AbHVMd1xoI3GNKg+pSMT3GLWjuL5gdUI/ZNUWdQvPHjUz9LXIPED
mnkBtthZv+llynEX1uO9CZVdZZHOSrMLbvNvAi48vKV45aVUqEqAsEu9c2Y+7wFNfPq/isCjqe2V
iUqBDgvkhx9YHLtQWxmOWpWwvdTe378FfHZXzVKoj6yILIQpdZw00d4YXfeOJg/lcVVOdjGBhC7M
OE4/d6udZwh/QPm0BhIMurRXQjBXUmbvBFQPcwcuC6hKmWC29GhhocWNsGshpdwxxRaRMYy+0DCZ
n493PuYMGL+8sw6T+pRhPdlE1RTi/Hy4HtbFfgKIEoCWhWeMfMfCGpztCJXvtZRKshzhP0ohJSAC
rnmE65WyfeWCWWIufrFhHtCMVvUnxnd8XIZWiJQ/aE+NlbID8D/YY2eWRF1nwyY25POcAnFnUFYS
0LYSFe7clhsG9XA4J2veMbWNsb34ZOv4kNjJ54C6u7bbwDJJjqHPPds/fej5pJnGShCqfHvWLuNr
HwjT8wV16/jOvex/hYGIsiwNAg05LnMH2h/R0hKe2sCIxCYr7H/SjSvv/sqnkFCCADhsLNFGA3b5
UPVEhUFLuK7AQiDPF3EX1o3USPUCkdSgkBOCJDOINK+CqLHvBXCeQhPhte9tJfWWXE5iNl8Qt4rE
fsJ3pGHdXUvhgOr8LnX7CzpAqxz3YxmvJi36S0yQNRs2gWtAISTrI3Af5v+EUjF7UZHbnqAqoiD0
eEo8/LsYr0Cko84qQ+oVf8ITzNRzpT5pynRJUiznu4fvvn6b1qEwfLvPjm3VLB04IlA+rR99XNNp
XNeeaNbIIf/k36MKvYNWTUzWKfJ6x4+/bnRJseh1Iwf8R5FAuSE1rl1hJwW6U3rAvZtrk20+Mp6f
d6Fd6M6PCiglRQkGD3arblXyKCuPB8FRnTmIY5w4lqpJq9THa55zC8kpks4s2lBDSy2+olvjrs0h
42vI4ifAHWaiacrIfhRnI22RJUftppca50ceJ2og/IOQ4+WHY8d8Wi/zSuSzibJ0IDXikoYpFfwh
4PVvHKQkVFnsqAHOwSBLtRGewHg/uuBq0qEjozRu8cfYFNm13nzJf3fuzO965f3xe3kOjex8HNGE
GVY+ZvH1LvDaNDn9cKob/4tj61RQ4n/erwepM2MGuZ4GwhiLlqnLxs9dEk4MrKAUuAwGoRUxi+To
djianoXevOp5QDCPnEolJKMc+MWRoydCIZYsjUVBSNSSBLNWVxlqjrLvfmfk/gyPZIhHd8RqDMi9
TUZAax42J/psKD6rl0gutTNe/ucOTYf/W6oK228yKgQcJrMfzNbFiPDNT+Z1byxh7J573PCdunoY
bImIgXtDtKAW8C/sHfpKQcx6gMX0XWPK6YbN8f9NRT2Eid2B9SjwkKB0eezPhz0FYtIXVuMtd/E9
CYSpy+S8xcG1/OfxgeDWE9P7uqNviK5nJoILhuiXdf1cF/86w9LGKOk5YtCFCmji+as14Dh/9jbY
Cq2Gq/fKKHsnneu/J/+sFT1su243T+FoZM8dIkATBG/GL/gs7O7zqiW1Y9GpXCDhG9ZI9yswWwuS
YVmApA//OziiambMUoCPshqt7ZAjaZJxchj8MOonqeB/EpQd5zKGbK4mS6q6ik423STeCeO2Nkg/
N9+XhAEMR+KlZSpopyAhmpTTfYfs2q8b+xJ14SwF8jR1MyWn7v/Ibuv8MgJYXxQIVAHenVOfgRqz
dwfuH4aLMeU2cKQyrzPaEkUKySmT1WCfxshmaxF0lUzThSbjSUVKUqGc2VwRb1IlyV487ynqxiJM
cf0i+K0mtXkbLI1lk0oz+b+L7c2L2/P4Uqp8Ip9NYoiG6FROSwR8r0/ZMTAz6aKT7dDEsUYjKZIY
npJ+xHgLuTVdoJDHBxe3O0mDTmW1tze3yrNlZHrEZT/wCqWKdGfw8hDESSX61yvyixgksLQlmWLX
FzaVkbOrFmaCv3tCx/X089TrgntL/0cz0VQ4iyu3ewxAgFevjzggL9EpqEQviYuuh9uhb85lbPw5
Xg6rq2qOmvz1ncPCC10PyFTC7q3qMHGj5mgK2k1Xc+8AEwN3N6xg8fJXp9lAiOIgvSjM2lTVFw66
PdajXRffVtWGJmWZ+lpR+uejTMiOw7/6QtsFdL1ZVFO+QfdpCDb+678pXmfMc4xCq0cwsLCtOqQa
2PHqZ6o2rofs6sGM7c057uZf7Mm5l26rka3V6rPb9C5OiBt9x69G9TqX2MDQ4qISKAGftlf58Te8
GuACqbu7VjRmYERtTtfvs4Vg2+2PuEQD62pwxcZZtwlM64dCOMYuZiR+wJci8JZSbc4WoN0L6z/p
PojLVP6WLtou1XEzctDps+D3CDWZQusW1P83rmgASrqtvRqFF+QN6hoccnC9NNh8MEm5RfosA7W5
C4Rm8iyiujIVIK0uo6yJsezuSrbdnI97402sYBunpv/kDgqtydeHHOJ2UvDFowQzmoq4nttRf+1S
dqV52PbW7GlWUQb0ByZ+qeth6jcpXa1XmHDVnxdyfBjiFlc+IDCK0fvpam/5usSLOsyn0/YgkJwW
wiJNfcmrp11jq5omTlHZL1HcxPM6bf2ePxaJaRcuazPh0myKYbZ7XE+ZtJCmAcHUL6E+mX49hf5d
ZtmNSup1xjheFMjfchH7v4i3Pm+ONSBGhk9zHch4JiGceJtcYfhU7MChaezYDFtoIsVX/los/2LN
rfXNI5SD2RWkudDMBD8QXE/amtzz3ToF/TKoK8/VLyuCEp3q5Tvr/ZxdN6CJKze542qrg1y6yUZK
S7dzzYq5Yn2MTw1KSFzSzMYvv0/gHTa1V33n7zSkJDBTEPpc4H67CJdDpAQt/HtFt9KBNUU5C1j/
feQ0eINZT1UvJtu6X6nNfXw9CKmFfw38U0rVea8HkFqiNPO/9B+pmzKJmrBTVgtYoQsk2LGNeNoO
TyMwKIJtCprkkgrS3RQw4oqJbX3zW9E2jfnzzyxXGgXujppyBy5ZU8R5umdU1lTN+6qT7+JkXb+P
ifZ95sLHrPrC/He3vE+0lQ4WFQ1pZcFFz30yPSp7Aoyz7/yt4k01QuuzdrNXIaCBFEy0tSc5Dxvf
EWRv8FTs9mWAwZlB90BVCVzPAQgfn3YrunF+p4ZUTdRZUt9NjaS4sJhvg7IKrZ2HoA6/iDLvVQKx
jJUEdj7LK0D8k7pf5Aat0xC3QLDCm24esQPWAvDnkOf9/2/Ic7PGUbr9+VkfsfnvRZJno/PPAhOP
or1PNXPuqfrbRpIdw4pX8oD971z7KGKfYMrRPllOn0ziZSY7M+IEasJhscTDiyGIMhDRf54Bhzp5
93j9BYnHwbRiykT+8ar/TL2+IRQPH0P1LG7y5gQSn1ZOKAA9EqhLVYt25ZMDs6nlqf/UQybp0mf5
vFBE7G18XSgZ97q5f36k1KxPRPtb8zKwlQC5RqbSsGZUP+H7OxSAdIxgDSjslH0gBo+rTPVbCzhm
nbzxW+q5Gf5ckqzDvvYB1fLNnrNf6Le73pHey1hDWJp+MC4uGdrU9GT14xwCBIe/W57I/vCPkqxC
mfEfJDsD5OayDewbW5rodvJCserPR9ZMIiKH2YInHpfuFgtJ4oo0a6voPT+1HOQRUAlgTYWugF8W
oF7hUQX9UQds1ZB4h787jS6O8K3q9UzvAfAF8aBRhvAHw/5S9tx5Dru24U7lhvyV93bm+XZsMoMD
d21ofIQ5bDykyKkqGNbbTrZ09yUsoC69HcUVIqf1+UmKBPdNv1VCvpKN+cEdq1RDuSPy3nLK6Lq1
YApnZP+4TBEU45VUnSJ8GnrzJI/+/rJqaAg53wXioWaIk/lNU5WUqiGkn+6/tWY/ujhGkVKAwa48
xCKWmEmpLqtDHNbXN1x0UT+KktHewWgyXTRIWVfPK76upAo7WO6nrDNrtJtQ7VucghNF6OzO6R+W
myQ4+KT6PWKQydfl8vLOJEn92iMeTONd5GpUt1VJGUPOXO2q2N5RH0B6Kj9W/sQQcxNW09fBiFSe
fvltANwUNxvX2z6b6VIzFZMfIMjBo50R9f8J3UDZHrzqtqnMC6l59QPPPQ9ayu/tWsi2ez5fYnd/
BZc0uLLQU5F+OZLQ/asOWkbWDMmySdMM7LOw5W8/vnE61OgVL+/novxPHD9ZOj/9R7yJiwIzKO7Z
mpPbyJYIydqKja3Lt2aiW8vsS/MdjPhjQ1OhJCRA5+nKk7fZKB+FJhNb6sv26UwwDJIEVvt41uL1
m+KfaVfny89RZKNadbf0v5159KDVy4n21+U/fSROSGuFPppJJrzMNr8K794OYSBYWs1WjCL38O/a
FYQt2sryiYFsooLZ6LZkVbV06MQxGlNPKux9Azt6g8aK6+otqph7NkAuHbxef/rCNsryDYaASsi8
ZepFfDnK5nkDgj9U9v4NFUL7jBdybghA8ONYByBUPwhMPEVVfKWxtehpxbnkJFRoMTjCXOZk/QHN
GBC5TW2u0jBkv33Q3bjoE+10wgSE7pEbw6SADgf0G8bVF1E1rohw7rAhW/Ffu0EzaGMEvRWQ8IQV
jXKj9Td1Nqn2uV5C1shMrcbHwhUAv5clLOOYQWI1CiDxbxrGXLhyQD4LbBlicWq6mQjHRDyMDf2B
hT1jR/x5uXsWDb8E6zf9W5BVKT8KL6T9+7KCLQjwTRZFsgekVYQpbtCihndoFXXZWGOCIUk+3A7C
Neod1ltJpDCo802HwM5VMvdW73SoN70HCpi0tIO63N+9ZECwScDckqq2lqdgD94v4/hmJ+GJTNEj
TdcIjXyvPaU45lJLDzhR55p7lNego7E8k/WLwlFkzTCDpZUxgojGzO8I5BesCLhQ3JcxsoLUukFt
gKZ9Lf0F/3FM8CdBJqzHLmvOxFfQ9Q+H1hb/XxCxQAQKI8I2KlHxCppwrIQXCJ2VyhIDk2VgWVmG
2lyP0nYYqjGj90sAsndIcosdjfEHbn6Xr14eM+0LJy/muPWLq0CaWZ11LCN7xSDLrEgky8iMsOCS
DQVzFiuTsEnit3PAEsaVqrtEgz5ErXv5WJj6cJrbV3r7+yQOtOpuBpnnwaCm+1cR/hdrmlet3bf4
krc4vyjdUeQCwrK5aMb5oaXcPouQR47CemOtRnAmeyzjhoOkvgKh/wuNJ2REtbHvdG8uIVd0M14V
fHaa2/T+4BAqW4h33FxP8KRPe9UpF1WIhbHJ7kZZrza+gC4q75LawajUPoC7sirbq0jx55CkyB2K
DCJ29A9fA0GQ4/t9D05JOKmrBSySIDTjTSoj748af8Z3tiSyS9seVhKzPetTpEL+hLNZQ3VzcHpD
HJvZOUstfy3RDiGefKP5SoyuA2tgnxLvfHl7IHzz0FSSjcPtqf3p0Qg+qzK8Rt1abIja1e28k5A6
+CKFUG6sTGkNaE7A1YCKjX9kXuRFMO9HWGLyWRsw+jxKrraC66urrO0ihwfGaI8Nczs2rDneYcGR
4d3/CgjjNiiI8W1OCs3jTo1iLypY60VpF7+GKsUULzyWxYoLaZtvS0by0fO9HeFEMq5zZxGKHSSS
2PaiIwJJsKE9GdOTSW/C6MArucO6mpRV08qdUB0+4J00tP4J6yIjEhOgO9UgNb1EXQ24v+aISh6i
Cey8K5RBNa+3CO2kop/aeMi6lkLrTUlxDvKzmzQxeUTIpJ4AxTqKGGCIZpTr13Wp9B4YTf2wekxf
wlG0zwlysD6wNFoQeR4W8n/C58z3L1H7flmIAiC/UqrzynpTWayNolNGti8ar2XUP6gal31a17N/
FD2u+GBIQX5k9ChBxYpdp+FkIZkiYO35S1Aypd/eZOprFEhy9yF9FM8rpscxFTTJRC8Xh6pOWcKT
2iI244/C2ITBqCswGudVrLvUWIYJG48BoSKPuh3fQGLyuektvtgR495Yvejm0JWUy9tQQQMi/K9P
7aIk+XAj3p+ZIMXUmcZNZv/U+GTyNV31SZ31ub179WfddXdfu/vncKyiPaes5cbaEufPeBiuu4km
K3Ftvipnc6PrQeXBkoiZABMNAn2f0a7sp9K8QuNtRQ5Qyh+UG0RifbXfml+HsnJaZ+SMt3mpnPXa
rrovz4RLMTGtyj3jDqhqP+Rp5/vZJ5JkmpSJmbJx6DqKo6x4k2lbrYovbVp+iyVHtiKWCFP/YFOn
oYx7+/DchPTn6jcbizHmBagnOqqSoDCSHvW8gHi4LHytZrkLvS3PNBajyZl7kBIVMkVHwb8AiKko
XitL4lOJnCJw1iF4VCR4Jy3/K25PBw+J/zEZm4YzIafLm3YrwNXRdbY0jTxe02H1MPHdUS1B0U20
umNqES9l+Nx3PGHPnlez4pNhwGc7hFye0zJRxqtG/ECXKp3KWtNgAWYj7zbF9mlNUdwDj57PKBZG
wlO6ro/CXF9u09LcaiqG51MFQw0nND/aUh2SGFWCwgieyhN9/Ls8zejpRJ2HsvBXgkkaF/374SQf
s7YAUynSmyB3CtAEgT5FP95zWDG9hjuBPe3t+RhUw4EhhSvqCvg4gNT4Xeekd6lM8U7zgcAQRErV
Oxdr0jJD9Av4wH3GZVWY4Ao68Bon69zmgBYKt6MTIgzxfncO0n+8SqBVajfc+PL1RCm5OIdOnpfW
GVP40UP+TDnY/sIqn6LK5pyxpTwz2HZ5jMPLBX24BQLMBbizU/MCngJGK70ec0OxibGrC59pcC/b
dmXzqEq0dG7CtG58zDpYfP77EjQ1IVrtNKPLCaMr4IMVueFklPcMFW5HqnEXbhuV3ZwDvCY6kdYh
Luof+7YLnoQlRQOdfhqTzOcww52bd0RJ7m9MdBvLiYtmgKSVgUKXGqnuSnG9z8Pg68qCrXGs1QdH
aMw+kk51oNFkVhjtlAkfBzU8Kfa8Wypd+IitegbN1voaGvcegGjPgBYaP1N4lN1oskOa0+1wIiWz
NXG35csrgNUaxuoW4Xb1EJScSsspGBFVwx5Mhc0nerb5JyoLxxjOVx4sIBFwjHVIknHXX8AOr7G7
1Ld3k5i8yEFvnUQUL4b4TTTrC6KUiEmWJ35cDYECD9fwL4UIMysUfo9HEuXnn22Ym0/A1ckggt+Y
Pw8IPFK+3HCdk6uHMnJHld4Ncu6KAxFgcnnLqUEN7oQuUttthvKsHxhyX28y9zC8b2bJy5j5UVkM
P/CM6AoQKK6PljptnqL1fv7o59kOVCA9uGl5XMWH9AW32EnFlMWpLrsTnLIgEreOgwzbnXsaFrQy
j/6jysj7aakz/DT8OnPC0vDtEXds1jhl07G9+JjFqHhZ6a8FwMTw1l6HLDxIZafmIiaPsKXWvo1L
ATpPCmfXzcm0OTuBK+MDb5YLA8GZN19cTmqb0RPnPPRA/8pplbM7DbCH6j+EqJbKNg1XTPfp3vj6
a0b7Effcqq+GcW+LhVywjjDQyEGkurpi9zpiGhTrYnJhfEzxQ7HzkMDNzCzOkjlqJqC9ULAdBqbA
wU8QS+bxOvvDblADXqD/+myCHxoNo0O+NFq02T76+HeL155Ap2c4uTi0rWoK0u/b5skOxdXeNPnc
i5JgK6LwCo8YMpNe/gi532V7QPEJxjtiJosgFTkTc6NJrcHJhMj7HhH/2cjSp32RgnCZxGa63D33
j7t0tYtGHlH55ZxA0eq1mk40uvwmv+5QQ2ZqPptQvzlNaLVaJmI0adqtbai9di+TDkuAIQc7BlCe
mD+GrVHjrM7oDqVrx2voH/qkEEIruhpsg+XoC59ds7umSDPyOifvkzvYJuQtzVqryRkiHW8gvjRJ
GXHAtXhuDYW/BQ7aDaMki4ELV+eUlyTifAyX7H3bGVFHH1IBj94COayyJrchtECiYdDt0V7yOfPk
Li1dQqgX+Tmf5Md/5wIlZ3MZfPbdQM9/4lB/CS8A4uvoVyv9S7jW21lsLX/SAfCTjtq4UL8sQmif
Qhdbco9HGUg21Q06uRdl8b3Yt4tp2+T1Hodj9Gpvnm6Mo24iMFOMOCKCJHjK4IFufeODgyqvuLvw
E6LWBAahe0gvdt1M3HNWKmeS1lFvV7o3vcIV55rcgomsjbkiHt62I6ob+3etJZpw95nNI7kYMnEO
hQQz5Vqhc9d6xD17drXaroy3JqlqTGcRH+FJOcZ7zA3Jk5M4aVSe7v9nM8vKdy2fwt0YP+CxLRGU
Wivsv5cCYIj5T5nE0ZIoaV4o26dA1svnl2QpXgYPVbrn6TFtFAUVEWofog/5aoy4U8kfjeW16i+m
qXVPOtM85Ow6wm8p7p/Kx9yrJgxytYXNpi7BDTaQSe6qivNxNXCbEWxohntPp5kLuY98XMJBPxCE
BhgP3oPNaC2z/WgpaH/d9ErUlfyukdxfd/X+QBfNDeZ3uZ1T4VmsYz1zS/BT93088lDCWLIj3jAR
whtmhDl/wjwJDZyIQd8DCSjHBTLy8CnhcM9rDZFYZFyeIX4nnumH1RLuFQnz/spimtISYbT5827v
GLgJh376coqXi6l0BuBCQ5BbLAnNC9oCQqb1tp0P/LFJSvLbZJZVyIM1AA8gYnXzELPMWAgBmI2r
ImHhF1/+EhLMzDFBr1cADC2fcVi8nHdX/Gdyp74hyH9+JGsIUZYWop5oQ2mIEaAgesarfJvaq5lp
d1xwzyKqdG8317N21JLyzOiQNv+kzeO0F9aay6TFvn+MYBHn2qqFrGTf/pNYgwx1LLAzigY8cqG+
11TAVVdlgSO+K+LMYH0+BwfVb8lZu0FZOhDi3xmTgET1nFkI7RjVO2bVDelHIdHo+oRoX46yTYE3
2uQuEy3kdND5ppEj/dmKSyouQu+w8EgWlhviNoAH5wxEVcTb82wX34ZcEWhKZjI0ZSdjwZLTvOG3
ZM2naqdsGBbsmKzh5ja5ybOoluxcfDBvoSltYEFcSrnTh4vR8NLRhElm81BMjvv6YYkKn7yTX7zs
/4FrnbBEBJw8XEz8bCNP6y6JpOFtzbFVKs3E3f7XEFj/2ayix97gil0aaJgkdXzPFXgPtOknjlSl
K18tutyXo0sflNdnQol9KeLjW8xzQZEarM6E+BU71zmBxXHYErztWtOrmgz1xR16s+UqFS5sEm+e
SnBix9vXZC6U2gsFgLUTw+rsAYM4d/MgL4GwTxyZ026ItHRwkDH05UdoD7odVq6OzB1NKI/acy+K
Vla9j2k4YnKowUN95BFHT+yNA9jByFesv8heuHjnFQu5mGjocdxbukP/ZVjZcJ6LY10r0QT5hdR3
ynPVezgzcNcv2LE+Zjyg9VYCUv5wune6O4q+pNEYpS5aP/BGjQlIr+ee7wloe9HZjJVPBlUsnYEe
iA95wTs3hfw9epgRUrnSSzGAD//ostnkZKoskDuiIXvAm/eWqcIDVUT0AkTkYGZa/gib4ULr3CMO
fdqdS9jiuALiPglr+dgI5MT6TifddlnEeob9syQTZl2oSlics2U9oAmVH6vdchpoDnR08TVY5Wdf
42mRNaM9168b9ttqsq5Fl9P4g5PZFEOfKJ4UyyG3oSHsNZ8/Ir09ZmTUcOpmtsUd/fy8iTQDICkg
inBgKQ8hgcucAwZbsTAG5L305k5cBWmosuu2EZui+Haj3+Of1SqmqQW0wx29MXodb+8BCvsj8o6t
aCue5RhUVbI73dQ2hf0akVLdy7A+lqXa+vndFuYBBjrSDCTtD5ZPBAGZA45HQNxONcpGG9erEany
f4w7AxqkByoKjxGaH01dOQgTq/+OKrHTgOMQUIxiJbVK0bxfas8xT77IXz07U0Xha+MECuJcnmGo
/6pfXlTsRCFQ4ylcUB4bgehXNMvUU6aNnv9be0nGJTegFnKBigHEitl3MK1afbmbdx9pUteDIbdg
2zdVFcDTpu48agMjScmHGymShqJPoyU8KzCI+56AJCRDUf9L5JeYBBA2cS3eE0aMDWPmNtjG4/Ij
nnvdAfCleEUodrl/7k9g9qp8pBT5MzSFVgg1ClGwGGAKMqoD3eWHOcmVImHvgj/mdePYLdSelrCf
tWAUt4M+ELNKU5Bh1znxi09L9zs0odUDTnJ5p3/A0ht+QHOtuBNERHjWQVHkr9+Le4wV0Hc6kMOC
Y1mL7By3TctNF8zIsrCKo9EwA2T1yRVRs8VIzSIG4YQPoRJRGd09PxaRxrhyCuNbQApwqcFZ0Fdp
sb6Rmx90ZehQjxT/pBu/oiMWdkTsiEok33P8Cu4Wh41YWsbLG6XVDZ9JUgzv7ZHPAxAMq1BB+aSc
3rbNJ4ukY2rTTOQ9iRgpgLUG3uBvyGaoaz6ugrZO3nN59884Z/09cGEjwzJODOcOLEjfsUOgIXje
+kbJnFOLhid8ZC+x8qytLXGvziSpahcYg96tjT139ADC3zfLDmTuxu+FIJfVmAtsfMtbMnihc0ob
l3ghak8ke0f2lISILNQ0ekMGMZq4YmwiZhBHfA+uj6B3erR4pysQs4fakp8VOJ1UPSOJdNdzMGqu
r9E5OQLFWrSeuiEtan8fgsHbcPggPxRdTEgY5TYMWn+v9DjtsfjNN6QFi8DkzOqJX4OmitraY+UT
UHa6KNCo9sIKnDVIVvinTvweZOPOTE63TIDGKPuUTgRHt6CputxwdDZetIr5C3JGXVz+rH/2HLEf
er1qQMBgCWXrYFRbBF8cfJLai7XXJn+YU7NyXtzzxsZUuXQK5vrDBJsePoylg1FwqKg+8XWMJSrq
kBX+jZJUNXZEHbWPszeeQPK/802Z68eSOVrpipdU/Tw8mXpEy89Ep4aY5oibNvWhoDCb7yY5Eu74
4oFatnN1uKL5aMzws1reKikXYnG+D+w9HFWu6dX7s/PNGtoAyg/5PF9kL1PQSj0CI7qz2kpixSN/
M6qsFM+ZRrdUBh+ql/ZYhYKcjg1eimal3DLQmfp6pM4yOwJ3UrmA6fBgV5uxyvDOQX0liGVJr2tx
ROtMauGqwASmjeCcV+ElojsYHVgmczcFtAboqSYMmCfrKb1JWq64JCj/e3olhUrn8aU9hqOSJilX
1sYIhL11ktlYKsFC5ouNJ6P55ygZugyC0LxoIzdn52LtpV3/EoGjgalYe0e+erShsH8tS44V59bD
wlJjO6VMSlE9xx7DX+jXB4SwVs6zhHObmhEJyQdKFDWDsJaebxmmiRiV+99mawgJ9SRV94zhC/DE
7bH1JhtYu1izcZz9pUu5XJ58C1tQcI9WPJE/giwWMoGL4TXcu246bh0MvuoCK/Qq4rcgdE+94MX3
BxG+1ax2vftdK4OCowaQvGNqx5iepMlTDgQq/9X1AfLIgw/0pnP/GTSvmF0BpD4HTRpxShNyLQAS
ph6lhfd6hlSQiBHyiVdZF6GEPKhKmDJx9PZRaARUdhBS1LTCnZ6G+W0SS21BdxNru1o9MTGMNUnE
yBV4VwT0Jqb5UVACJ78Mw7im1VnOujXnGBXNaxaDOwxTK8qFJJW3qQKzII1P1zWAV92LDGNmBcPW
Ek/OdAEJX142OrhLDvjt9psmAx6d59QohMHQgPM44Owl6n82YX4cEiZCCc3KATSUZFgPietAH7jp
JXQE1L27kJXXokJLr+OHgNNKfgi6BegRQkxQFUzbBj3UYoEFmTuWNL+4UXuziruIxrH+JyJNK6bt
p8El8ajNZ5HgVD0Hi7EE91xazBqauo0hEmmdLXetlBD5k0ZZcjHPX8JawkKQhCiJmhpYEYMl11Jr
3C2wH9V+axKGi4kOlGm+co+ibUfkdyrC0ow8fONE5fVFHE+sXPnox2NVqbvKyx5LbLSMZipIkMZR
lDZ2UGo5qDVcIyG2myRbwZSFz7+XclCTV5VDM8uLz4t/7PaS7Kn3BgfkGn16Y7yDX2LMD9FvG7gG
8qiodQ3DjmZ1xyl8XsofeXXJaoC+KatmyifcFzK6cpt3+NKmqyb7odyOqt4LCe11mAzM8U2y7P/5
FR0KlkmZ2B4oYcWWDjJUtVmjLrD+pS3+P4snduWVWDNn+gkUWlcbyulsllZU6f74lIhIq3Sq26FE
nUOl+ZJGAWO/TBMK61cNIVyif9EsUsXXfHOz3DyI6sh/SK/HQ4UUN0pf8g9R/Bnq9DbLoeVWCqr9
EcAW44X4Uo9GGOW7vSICkwVqjh4r0K+/lVF3uJ3zccCpe48m9UXxahbjsngKu0d0744dh/QBUwUC
DqpzUndZXxMiHAUk/6Ct5gzgQ0rk4wVp2ty6qZ39BO4A/A8B2+2Cp4Wyscdx0N1J/TZ8WztrUy25
OHp06rhbZ//1ao3BzPWbIrZN+PHUOCWrRDzJxy9Rk1Wd1RZyUm2Ap56eoFRTLok3awnYtkUu/xWx
H0EiEt102hnsmHZI/bJKN9pReWsRolGI3Ue7e0R4v/ewC3uWIjCep5wyM3Dbj9IsZy0Z3F+466ON
ACeGCt84T031mpk0adsdD8IoqGSOqOmQ4c+N0y+MOIcRI29kcZXaIkKjbOXyZcD6JosL4d39EddC
jc3AfIbMDoSg84hOoBa8D5qOt4LIgMmAKLVHvqkBRU5JnkBNBRNsDxUK7Z/hZTq0+/vhq/0aDfF8
/er8zK5a4wA3G7RvVjJlbSXBQaVTqneGuv/0k/VTJogOpg5oXRDryDuGeMuTOv3RbVHdhBK3dPJc
ykUc+1zMJKmllfdz8b4R2WUuU8ox3C7oFwfm1x2VXjHuypJziOyEwKIFW37p1WQSdDuj0SoF6cjk
rQmSUub4OpCYgXsmnf8CSxNQCJIn4N/LRNJOPhlFyjmkaT3hnkT0iDfvXyIvG6Ivbn/KssObZ0o3
DOwegr960mKhzmYls7yphPfP1MCLYKL5q2kmwD89ZioRZC8HGBYxXqenh28SNrZcG3Hc1K/BUNvg
riCG8sQ7lINDcc9xnZEUJSQKrpMppBknaviyxcy5npioX2ilW4+8yV74G29Xkhj2GbUVFc0fxItT
xN1Mj7f1mt8PiTnW+8vq8DvOFLf4xHvj67T+c70eDlDFQIoXr5gyWTnhLveZVxIzCKVBsCfZEipn
MGPZH27KNkiorMin0UTl9e+Ph6CEuHC5KGuTtBPxPJQbDXa+4O7mEsoX6k48lhEupAwR5sPy5DGw
GeqSjcvgpiq0BH1JC6jmrs2lIZ6XMlEGnJmWU2Vcg8foKfMsBjBv1c0JqldmaHbtuD0srNYvipOs
Elj07XXbo8pa1DasqUDr+0S1h9ziS8o8xSRZ4SyVGYtL70CsSPKh1M/N/GjSnaGl1oaTbjBQahHa
D1m17076aS8L6kLMuRll5q57W44Ia0FxxeOv4KDLBboCrcHpNAsFkXOwc/Bhk5t5kS/pit9MBQ4F
SPeYJpFv7F3ozbetkbC/AuYWjJ95EGVxEe3CVm+V0MtOGkkhNvDnrhP2aPgqWd2RmUY7WWKhgh8u
fd/QTAD1xJVyqOzGZUP0PpAkMQnPXjNLv5GAOdQfB+Q07ewZzA28STxU1WJaZI439T8goMwPmG9W
83GxXcBCgmVXkqaJ/UtT1iqh6PmqtBgPPl1R9RVsPhAoHvWi8WKlXBjClxvfS4VFquNKkpJvmP1O
ZWDIUb9RxKQBBiJUXaR5NjxDFcIn4H3oUmWfFmisWD+2+OwPJ1hCu8dGWw8KRkR2TrBR3BDOIiZ+
wWnQxgj+AS4CwjZCecPjxxbFwINHvLzXfro+biSw1YDHr9OuryRrzuXzYhpnS0DB1W/R70SrZzJG
/0s/tkeWSLWyDB5GTsnDBgPeGOkF070DLGKCHwbV9V/kfU7zyz5bHxQgOd1xpMlSEeJxnafjjDq8
APyj1+AwAunVe7QuJh9rT2ZCO7d8LDgin779OOsqbXHZ1YyV5iFskBnxCqtTekFxMYj6dyv9Agyl
RHgM+Jp/WhMmWz+BIh4a58Ye83jvYWEKyjz9einPTmWVWjjsq5pVmgf4OzTBGHXPmfyi8LsvPEvL
NMEWGopVVM+khdY9MNFy6Bjp9GyobV5GF7LhiBo4k68QGEnj+/i6/nSQ4tdd2A/mhqUXE1j79MVZ
AHW3X8Rlj0PGjwrirAm59RCi90s7vpeKJa83utHFCbBUuBoSsMFzsb3/ZWxrtJsLVBHWktnLh5E0
yY8Cy1Y2Iv6SySAYnYProkRAj4LZLM3FZAGAO81d0SlfdgePXfjxXchZ7tKgceje7lD2E7HReJAN
8EUDp1YwjLdhcYqXKCy9xRqDpS54y5tL6GlUwgP0e141lL0+hLevkye2B549xu/aMLvBqB8ptAS5
wEvht5yD/mzCzV5nl2kHKk14PV+OcaZxQCEQE+aHEVZwaMmrxINxQp1TXlvAu/V2NG+wHBVUs6QK
TXcOZG8YbyWiOT18QEhIsbyrYjKcBSuadpXYuJmuXNt8wOAEBL5iAxRPNHo2m4ixcqYk9LnruYcm
NWLuIDhtIJlJJ+tdd3glx9e9YiFIHz5GSkWU4HcSw/kqs6C090R9tdyBxujT8z/zS35Ow4Knk5V0
f8dm+YluQTW1oGGlk3maMb1kSTYu3vuZ45VgN0pevGBOXkO6Xu47fSBEUMSspW8r6PsjehhZZtnl
RN6KREsT5wkaTMxYtfyMAqtq5s3zCuhxWFyCiorl2LlrS7pWuO/aSHMIHa7+Ge8wI/X6r9JfPVz0
b1Nz3GyjKiWzYNv0FQIvCr0pyciPgUXAdIcvRoFlS8wBLIGKdxE0blW56sk3870wz3t9Yq3sKEEM
x/OB8xjBpvY+yoODS+e+WUdjxTpV2GlMLijpU99L8OnwbLncownzKTe+tm0vpzq3ampjj8VKnWEg
UYwE5jan+MOXjkfH2VeNVO6ufqavcsCN7p/2GXkTOXFA9P1TPTPVv9CnBfa71EGtiWr9sS8eCBL2
L/c/6sP7utub83PVvkzBNMIQA8cyZb1woF6PeURhJKqwZShpqet5DVuxcfKgQN9nxQmk5ZWYcbeU
aZEiItDRuqpp7w+UQUzxxcugcqI104z7XcwTmhHPqmMEorcEqI2AfIY0ViylQHicWgBrSaK82mE0
B/7mTLEuAG/fkwNkPmTbkdrZEgz55dOBoDx58e0il5f8OLlfpyNAIhvB4eiVVsG+XMsjh+JLhW4x
vC0Ay19XgRsF+1ZX9vmlBudTld2J06hkaj9I5viQT4CI6ez4eW401PHpnn/jxZ9nf6urnbO6ZkMy
ZdCL5M9p/YFcRBUMkgAeTSb+OG4L3pyyBC6ONVGIdr8fd7xxPvi93Kmva4OVbZSWsI9eag8BR85Y
uM0b5SwKOBBrerw+tnriZZIvgUHQv/YaFmdXl0HW1UOZpN+f4jkiYc2TIBQYgefWr/psoCDE0+Lg
MVoan1c7iRb5BoYh7xF0X4zN27+jC6jd7fp6eSGaOcBlj0Br+EETEB+btp8snLgg/+2gth3a0B4/
5Cf85ALSOyLPq+AFF3UB3Psy3C+4NmZw/9YgAHKyRk8BX06Ob4Tnf5Nr65YEphSMaZNf5dF/CA7p
+LoT054B/aGeI+p6G4yS635xBsI8QZtIXvNN+0d2Qg8zkpNxXVk4vNZRBYA/gyGfrPCssQTP01Ug
P4otqsNwwfyQrR65sfr/lI3QllHGkTMgwNnV/xLoiYsqAq28dgnuPChHzlpJ/rNDhXFKuerSPtv8
YHnLMtaoUYjKGeS1EMlxzjy/oX2f3SuxzJ+i65nqAXr98NT9n3O34LnnWB5u1Cadb/7tfHVqnPMX
R5V96YiHxq1vRzozvoSwzIx7krdHi2u13atruie1i2K1UwSuI2NZCR8hfkpZLj3TvlmiXsz6a8er
WoatnChkNeikeXIzDMarMmjjoqtvN/A9ABtzu94eCiRU4mhg9lXIv/BJG5/+GulOj1qSc9VtmBE/
9k0Ea8xNyeClTgFDGCVfhec6tj3Jgo3eSCPcA3SCPowJdI/gwLaKqaqoAIF9RMSShuUJzy9Hcchn
rClSIe/O5jyfOLLn/N7jex7mzy1D/1GSKDr6C9M5gJs70El1Xr8KAcE3uP6mJVtxNP7b5PHLOTYc
QCu7OkYyRk5w4negHUyRnht0DfJ0d8xjEpaC3+z8RWNVG7b+soHiXb74hpFpEG6E/u6Ny7GwPXDa
BB0wYtRSrBRjVOoqlN/Ctzc4WWI22RbRNmXcvLfCA9B62HhWWDWce8+yLz3gWWkLpUM9nNkRmoWt
0JmoBPg6yeWxnK7p2eFPGi/gfoaC1clXp4ey2omfORgrxMAYuHXw8wc3HhFUdNMTz2V5wzNqrxyn
xomHEJsgm+BtxchiTveZhOyQUpp2YQz/ktswUQAZdUSBIS//5RcQ8/vFzaxTxBI6YKwKGtx62LsJ
qMbOIrs8ZqplNGxlk3aS0VkrpY90CddD8+Oi0EaYupuJVu5PWR5CsCAUfoRv1TiygR8kHsPZKR8g
sBdi85Ha0IfE2VWcivfvCWJC5OtvoHl6WrXjWtBiiabfDsifuwFH40fFzwDUQP/1N0XYWNYlo8gj
DEN0GrQjBLtrnkRNyY7pMqJ0YTSx7SYfIjf3vminucze6IIJ/dhtLkEU2jic/2GpCmOqAo3KB1WJ
vS5DKw4+nhh4eaIj/q1sdiRoSCcn+NtO/nHSlbFpXeWa9tM76KeeR6AfHsAjNOJr5YGtv4LonekH
RM2nk91YyOP6a7eO38+ZK6Jt2xsyECK9mZlOClW3+V1p5LEX4qzONFI5lwd9NTym2/jBUDaB4yIm
D1OjE70bGxCUHpZZFRDvI+24iaoDeN3c8LIxxaraqzpX7tbCviC+C2t0yFRXa1al50k7mmSTMDeN
xjUWtYah3QfNX6YQwCUfSzBXJt8AkIC3FCJEqy/YSQRuyfAufnajlo39bckTX7h3fBtiBx27pyLd
h09eL6j/ZXMlPOSN0t4gBZIm0ZeMAiONzms+tNhh8WRsqVz4FXcpKZNTWxC/6aEJzkDMpm7H4Rt4
mFB+NmISiHb3wNU4kO36LxLCA6tldGgGX7HJaz+HZyGEZn7bxoaQxBPu+y7mdDxhT06OL4p0L81G
0wxAxFi10nD50Pym3Bn3F8XgAe6lr0LbdlYBVQsWLYn12jhcIiXOXrxCOA/RSL53PBMojEvCZzyr
hMvHXxwxZjTr9PyQ5ips2kMHbN2wE97ijkauDSd6rFKPgecYSHqzwc2uLjXHTcAEfRUPUVAvBOhp
XbrQ7k4qPZb6jLB3uMupnuPwbzAm5nzhploZLk7GEUNLersNJGdUNQgOqSS4ewtr0PcvVR88yMZM
JBJV3v8ZvYE87ajyzMPrACiuM8i2gZEXi27esh8lhBGh/z1SzUn5WW4MesXU4EbnGTIPtdeqDUgT
JOpst5eBjtqE1Hz4Emr2ymMmjm6VC0Ol1fDw7ZCTa9xMGLmgqYPUE8zESOx0zJWBbfCogwJsv0J6
3dT17a1OriDn5bm/GMovyjaK0pv4VjyVsaiAdyT5GelQya9lpKVKIpZdvABIKC01SN1cbi4bqgDj
2aHOHJFqBmvlPWrfuqEY3x786Sx5MfhiK9tJLAVxM4+tSaGr992BEtQraBytwLtb4FzrL7Q8QrGu
6gmh8iGN9gpMuhdQyAjx7nl9xdqLfInKpAC+f0LBS8/H8+wEAnJfj4mjdCOCq9bs2nYFZgtShAeH
3Ul+J5IiYK4YBtG4oHoLw0aYYReekD8spmJ1dgsmnIiOy1K/+koT+qblSTHUpoP+rVCPwue4O4qx
MC771pxFv94GaR8o9VTQPfHw0PGb9R1xpO6mU0wRpwVKOj+M3UrwKyalLM3/Xi6e9S1oZn5963Yk
EkozxJSfYKQ/H4vG0bWjdoqixqFkYGDmwBeQ7vQgnuCTtESXcAAfHdXTJz4ICv7NWhnCTocVapRm
zEouxGpM0ZKBtQ651fum/GYu0HWZvtAbsn/D8prBDale7i6oz7tSWh+Bz65FnYzdWhV3nYmJnfg8
y204pjOQVNfQ09jcZWqy997+pUU0ZRhPtzBY6VshO77MU3ern8n5kswwxGsxtWluGNvoCS9WgUZE
TYPlbON308rhTt+VeSUaRiQlZdDT9mdcK323RKAx/f6Khh27LWyQYvoXuzdZEDNc/uEdOPgyK2Le
KPqYVP/1T2T4S4Mpds52su/k7Msp9/k2flv8im1QHb3JFZw0043zBuxNqNBFL4Bi4Wqqt4fYtDZK
sukyc655/IV3nB+axP51A6M/ZTT/OaYsTJGEeQV6I0VoHw7K/1UGcSrdknc2XqZrZDc256Ye5lJg
dguxpCqfkT01FAbFJSHianY1ZOmiQkg0ww5sUeQMiS2T97RpGHYsVTFgOXWkLwwDxQEUXO/cCsPR
8XDnEQ0m+E0IFczA0GY98lRC9aC2UOyczzy67TxelsGXIeCvLQhv2O4KBN5LeH7fb718+SajZ5XL
MvX2iNaE7/PdFjD4RZ9B++iYXPHzBotnoEL7R7db2znalc8LXe/HrS0Rrki6C2cnXQffpGG2uKfL
sFjKYhjnbLBSRYMxGRcem1MaMQjX2ptUPLeIB22f+X4/B59Ln3H+fE16hrbLpqnyRFXkzv0y4LTc
nTRNAqyjy+1sV8taa3bryYPVVnko/CZWUW+oqoozAbJnmBWd0gEUYDRe+p1ae3Oiht2IuJ3uFfCs
LCHU0PRIV3KsZ9tD9niSAfC/a2dHTJ19R1CmxNy99mRH9KuFoLyjCOfelPHlySCnw6JzR+AotfAj
WklFoPM7sMdA1Rwy3TN+OV/HerRc590sMN0JThyNagLU/RcJGHwJedAui0+ET9YPuiaNNcT2SvjV
xpnH15XDXLlDkHOTBaSrfoc/EJ5xrWHeVsAWWXWl6GhopixppLu0y43QJGtABbf020qLP2kEfNL7
IMB6r0xQNnBW9rNk0xkDuP9bQJI9GwfI4GEMXheGdNBZiD4JAg0Kz7NPalEpSY1g0QTmqg/cexPt
SsEn1fXFFgnO8J6eg4NTyJJvD9da5Mg8z0jFi8wSygTOb8QHYZGHQr3RfUC9EsBv3fPYG27gwtrt
R97wYuPJ+2Vu6IOzSVXUJG8UM1l9Bp7UTB1T8xRJ9YS+67Eo0TgVhIDKSTVcTdzzR6iKqpaGXcBq
GXpgTEBRQDxUIvu3owgf5p3Oh1tcAebYCcNHY45gyKtQaXi5I14h9OlnRFCmakrvFeLRQNPEWuUX
jDIaUUypvWBkREUBTd6RWBwME36xfyi9/L3cWKyyUGJz5OdrqlK74ooF1NnSe2KlwcsO/Cd07ezN
Hi2h0jYiVIkOmKI0PhDK+ohk5gDvarNboTR/qBsM68iDlZujV02Fu8ELF26RmT1d8j53xAHnH/hY
cyfNDb0jNRlzn9VGcYNlwex7eNUN4ZzXQaZhSr0CpmnfaY+Vpu0IT/MInzqtOvm80GsplHDRt75R
ji+a9saMlh7GYzYWHCV/Qv18ClquvKsGkFrpDzO0mPNMJ4ZHWs/IA2rPu/U1pBVFdqZ/M2wMdPFP
l36JWBQsEZf9/Job8rLee06JGx2u/58zi86b2/3GvaXvNCpgBmew5JmiW0SH+k0NFpmHWUmXenUS
7wRXTFjc+jzkxqQtuIvJWlXWgh7zvFyM+1zg7hkKUi1qmUjilXoc1v8xYgx8si1kGA2KD+n5lThL
F0mOjF0AypcGDNIUu6MtW86nB3j21GwVEka9UsWgursPK5Mykkjt/wK0k0nvO9vVXIs1Uetl6M0e
RThdBaq4+x8voMSMhUjqlf0EFpOInFZd9DWt9c7Mksld9M2VKKjHgLSug8wdm8JKwuppNLHqPwXo
wwnPKj96E8tC7gFZovHRkXHh0qtXrmUIyQ+hLGWVLorbFhdhwce4Sh/Xzq1/Vw+P//mESrUOhzZB
t+r9jTSbrfZk7IwycqQpE+CskmqII9jxNXqBFIOWnrNz+A4WkmABRz9lW6GIhDdDaOayUXNw5oT0
+y9hkt8JpjXb2PC2GmAldxjhzX9W63XAQkyN+tMSSK2tqJXFp1rKZl1BUrLtk5N4hRrQJy4rNAF5
qdKbnJPTO37kXZ1aBKZn9+pDfhTLTDncaMZJJZFvNiEVSE4RX8ltDeE+qjjlKJdJDK0CpYcUnc6i
FKvqqmRKoOha/hYjPuYQJJ7rI4eF+zOrFUBigaqjZb01XO0IWK8LkSup/NbHQoxqX2OcGFaG69Eb
kP/7xHDWnI2GGdA6PXm2WTC+daMjgcEcY2eqxWNZC/qWiXEFHvbn08yIyxkRwwa4mFy4AKNCgzBk
UosoSjaeerR+ATzA3Dn1CqTeoXF/nzOCJGaKRH33Nph+/Q7TeRt9kpyPtTeO8k9A8WYZYp13xbKZ
AmexE4US2xPODW6LsEi0p6XC5PNLVbm9BoMcdYvIXMb3iJHrAYyYlnmNJX2Ygjkcw/u+vXzhKWMa
0KKHnAwt9GwMG1jEV1ViROK3ze4cFc6BssvziwoFDWqhXHtNbiwQFzLHYXSuDJ6DiakQ9uoX8ReJ
TRgKT/eklpMzqrZrjjhN1nDFvhEEvVqjqdbFd670Yz0wkZTcrAb3YtXTk53ZItRcOxJq2UYuj14w
M+Gbb6CCMApGyt0+Z+fcmQBq77usJ50hl2tnmddKdq/jcAEjiYiBTw10mY04vQrz/2SEUXVBVRyv
VcrhK2pAna/zyXUNLVJ8pacPPyzA3gF/qRUpIAE3Kjwy/rCVY3Cc7U0RUTxa3U/3xaYg9w6erZTr
28Uqj3M1Rnf7qIsK6TmqAb5ZBAuMLP5SWZpw9MRD1Rbt4sDapiaoy8I6E6artFwAw1drIwCPk+Vg
dPnvtLX8EsIUgRpBXvhBTGUgP24hhQEmEUk68V4VIJ5mqnI2RG4EfYMELjlByu/nA5wkyPtRdWp/
Xq+mq74PEMdqaO0311TW13sjhgGfit/GHpgq8GpPzfj38dkaM94ZWFjLolMdeKNaFUToRDhGVQxx
MMYvUCldPzzcIpuNGFi0MFa3Vs5bKCOW5DKFhInMXUahHI932d7+hXKOCBMH6V56vmz+xvoxpX08
wPOZtV8UkoMyuDQriLgbzvq6rbz8XbkZPVGZFJ2mKgw1rig3RcjfHTqL9vuaJyQGwqAhDXrKGw2M
TMya7FT7Mi/jFsaR6eUJj/QOmm8w5lKDHKVGUZB4tmvnar88t9Rhdkqe8bvfas29ai0d3gYlXOiv
SSraj2bydyC38FLvpDzo7dG+KvpY2S6bGypLrbKxGICIfFAQcDV8D0p9j4t+Pav1XLOmexD4XxCQ
l/gHlAXMyvFmEfopuntSNBQlDFq/Gsh6fNDeUasRQXGmFOngLTLcBcUNlQU9iZL0I1uEo2kh3U16
69JIqGXZFhexIyVkuhfOW2yzDVAtaojO1a7fDkVfy2xORXNxHeYVwEmGt2h0mUe1kE+VDQMowesA
PtaDHPf/GlWT4TU+FgkOo/xi3MxXt/hMpc4DFOTx9fjEzwI+wlCuSrbiOHaQjcuHiTI1mSubqS3N
k/Dl4d1UYL75zkgUBUxFgDOsBH8zOLROWZIEj9NWYxQ3ijzlz6CxkEviao0z9Iwmf9x1vUV+7l9d
e1jsWlmYcraMV1OCP2xwIcKWJaoAGDPqFg8hDS0DVDH/9lLsZx+Yk4jKDUMB2GqVsmI4dVmsvAjf
V/jlCNHNwUTOJNBOiEgwaD6tQoifr9ch9Scz4yYg790ERFNMjr0qt4dAzmiH3I9YiMb2WYGJD0GT
J8QWca1/FhnfDOEQFAQFZLS0E3Ul+rvp6cxWh+QROgQOLOb9s1PJjdFkoYeKE3QBEIq4rpD9Mue9
IWAOA6l0sz29YHs54wTfCCZHSnkvICcOQ8Nc5pKF5VJrYaL3JsViRS3iucWSD2QUumPeCvklGHfL
dleq0SgLLJ8lGvm4ec9EdqIwP0vpu1OMzyuqRuCDxz0TBesYOwMtp9bSD7wRSxdVrUoqleHLKjxN
tYpS74/2IzsKihOQJlQiisl49Hq3glLFsaU3r/Sfo9s9Vy/gRfm53miERC7EfAqBabdsWHBTxppA
KiASGk6Dhz5645zqe2rSs/jrF1zj2U/xoq/EV/G51iiluS48EOjlGkL5mEhUUc0WFN1YtRIJNhyf
b9yxQjkFXBa6R8P/UL68F/w2dZGGFnmdb59gfHNoDEuOPq2TFUKNyZaSMEJadXF25Z1Co/iFybkN
3Vk2NuQJo/fZrdXA2Ab1fdJznYUsTOuxCn3Mxq/qIs2jxKAQVZmaEXtdNSIFaQYMaSP3IMWDKXTH
U5dc9Zy+ck71XxGhPt2RD8YO0b1FKfUcmgrOPjIzf3C565r9/ITgNJjMsDiyFuZnITAauEYn8lVr
DwHeBiXgmbsMazH52ed2RwumGCIXJ6F6ekGcRR4+lK++1MYwAfsPE7pl0MYZ3w6w1MYWq7WmtBJc
mzejoYy67PC4vzwyRGGIDL0k+RX5V/lDfzPDX/w6FcoP59lkgDNqGVIEWwRhVL5PiBMLZ6T5N3C6
jE/wFL7yLlIysmMFeH28BRCYcCvH6qwVGp2sUsTBqfyfNMaSFs4P+OYe+RmWCApSXs1xf0fehZxH
XMO3ON0J517t6/Meq5DOIJlRMDh480u5vf3b5RZmUcti9oszy92RkyS7/7jKz++HFlDXKM1a2SBn
w01RkIsiFr7KTDGntwMJ0/rXIIbJ4sc6iSAXMkJJjbB58xptUULlkID2mRRpaluZWUzlrNXR78IN
3xOv6QMVAOhklCPXhKUi+k8nPLXCa1d+xX5nCY3gSWCth0eTPkdsU4ZIsOD9dUK5wuvhAIyPRWCX
7rD1GCNY4cqfBQVA3hzKjIG1Qxs73jeZb9lSC0H1BIWOQrTlbPCIGeWFoRKAO3mBV9L210FgSGTf
i0w1yhRP93BIUPebrYNkm0KjgZJZ/z0K96MQTm28M9VX74WeRvHexSB7SHnSxexyEBq543mg7TqD
OvYznQac6c1+t9Ato9juJQSO4f96TnpTYlztltDIpxQ+55CGobqjxI/7q9kKAl2FS0TZPhcnGjeR
Bv7FbdK4cPqQTPvzxRQjo8oqTLNcYaNErHg8+9s444RCIMlNI0NLwSWkH5S0B5qRI5TeVwSikXRm
dZpnWZeRZpNYV2rv9Ep4C+Ghwy/fb9i+YvP9Pw3Q5F7cHsI7AyovolalwM7btWWNg6L/f/SLZu18
/vE4aahVF02telCQKNEkmxHIEd9xSswvZQ7xL3Cv/lFI7AmfziRiQz8WoaQgaebirRPTOZK7gGV3
/LgkTNyhjaVuYNaonTWffQS4I1AlJyuduiZLOHIGZM9iN1EDimCnvCJDqCYLD/hxpHLf+yQGYonY
/Cu0wQrcpM22c9IMaV8sAZ06gsXeqzxqALr4d5Lz/3DJfE8D5Uk46PqGMbwtiig/NW6DvGlsRUGP
x1+Uv1P7rT3vXawqw7mQanlT56IBFk4lLmNjUhXjqLbS8azbE+/ibpnR5clQ0kQAdCHUhCG0jEzr
AZphZTYXHcVrnoRqc3X5qZ8So2rkQro9YtBAT3hBsZYqh6iQI6aoeNwnBBNbwV9304R/otBcr9fo
EdynIdQtC50PfNN9pUjdp74peG/8dr14gf+e3mjOrygGqIY+Yf0lxJjr67doJGYwwxPpJrz2u0nx
9oo0K87esuW43z++ry7+xbLsINxxE92Aw7biaB3ViZlZV/emmzzuZzIp+YQSyE3L1AyRFGQnbhSF
QYTQ68nGV5qvoC8InlNXOdeJbhWIWPvTeZth2nYTIExSu+p8jJChlKHNsIiUFBAi2XxXdIzbmRM5
Lg7UEbXPSclYSBLb/VulHFlcB54zxyWm/IwZ39w5xtoE/Jme4KO60sDNSsm016pOfMH58m0mFO16
y++yRymx74DKs2s+/VJYFN9sBVqe3IFj56DOt58apPQfSpotphfJAfheMSruR4MknxeFkep56wEK
Fd5/rkUHjQhlOYxJBgEDA5yvlhcUdo8Y5BrLjM2iXKWahc1FA2ufVxaFyFXPLt8ntfJPOvvlOCD1
BwNWGPPjyMRhuYxxZf5p7Kn1XUbXjG0y2BwNJ4dwcLY3PJuf2kOfI1W95JUsk2K7j7jfImJa3rO2
WpYfvoTK2S9xi9l/mNhh/K8CCWkt2cdXeXJDPah3UwEqL76CtPs+7IoWupkP3hUsaPXgNJsigNp+
9GHHojEKY+JjK1ZtrTBgAMqqeSeMxJbknidEYr7TzKf0wmp6OAv/mdFYGfVdLyn1Ilh+iOkKJo5l
He6nMmrj30227kS57F+iVqdyRzgz0O0eE7r2DKrauytzwOFH+EOLcJo2oLtvz0m8aIKCOdfVE/2z
HE/Z5Bel5ZrYQrKgERjOQTfzU8gsT4/UX/cEXq3FJxlTvMuWN3+jUSHkugdSjs4aHprtt/iKlP8O
IT3HsYxedf6ch1QuQqnhxU7rolPl0t51GQnop46suz9MbUqGxDZPD5tlAzcAv+UbHaEMk5uuB1l/
xHWQSWxFeMPmuo/IWVQOAiQ60rPMu6M/QFduIYselIFqYCX4ZTa8eA16qhwQsJL6qMSInvySFVZx
iuVXy8NaJgQGKNKV1BBbkWp4WmeZRjxYQA1b1ZUyAYMymBju8Y44os83KHYC8WHDmYIIn6xtyIB9
K5gAvhvJER410pp8GYU3BTkCOHFqLZTLoNAeTPwOGbZHS1RbHLV0GHw691YHQR8iydMG1fY1L3p/
zdTrXFGHNQRYIPi0woDW0g4b/SvuDQoOluyt+rGX6tjqJpyznDpbrAC0nh/s8qCbOkG6J2rcOHP9
wjj89jbDFrTw+E9EadlkNARA076B4PJ1B1T/RYtWiHHo0WDoZkYflCzF4v1/S0Yh5l7i56eBX0hB
DBUKONBMMZyE3WXhBBcNXtbdFiKvCYB9+4h25mos4FXDOFGJF0g4BFQTZDORKfRmpCHEqJS0Ut35
hk8bq++DasNo61Vh1A41kBd11nq8v2wmYfo2NiuirRsW9sqDB+57NoWUN2p+75qZwb9BYmWmYrM8
xHoeoKvO+hoUK2PC4MfF1iLUrqd9Dy7WGI4KYBiOetdvzuC0QYH9oXZzPbHO0PfnoLKFM6AM9c/U
RA5q4JyMwSn+d/L15lrO52CxdpL9G1Jt/I3jMipBNgjmw+dIGQOQyuNa5n7tr5EZAqGSNeTaqpxP
C5aijQij51bSLWldH5upNJPgprDnvXb0OuWaIq0MnZSRHfhH7vYy5I1j6vsWAIowJ9uXxudkE5QC
kBu2LkMb6mDCw2d2GdUTKmdRBjHyNjiH7r4e5f5KyC846JCMnnkQhc2BFX8N7qVCGU/Of97psoC8
7SHAtii6aT5fLcJqLz89ZAlXHuczb6C9Xh4mtXWZ/4zhHCCQbJ5Vp9SNAR8m9O6H+6S7hgoUueNP
q0YI5w94MiscoZ1jkjbx/n3QaOQRwAnGXvMWzyetH/cmvM0rDVuj7EGUik6TtUNJJnVbkMa+FNRM
55Ycz461Z9JisvNlv1RkxSrK0FV+o8ajCOhRt9k1MA2Mopoxbcl3DnRO9qqEafYmqe0xsg8P6IyA
g3w19l1+WqrJ5jqwwAJnIwkVEj5e3zAc7074YueTSvcRNE63X/GamKk4mb0/u0CrVfSCZrYMd76U
OBmwIaeswYUckhgmQI5K0nE9AVFMw+XGO522xAPtsnfEuzVfdRw5eldV9IsIF/E2E9w9tsNKCSH2
LOLaMiITabrgBpMf7saA93LXmpJGxcnAM8bJ7hMkNZMVunLcnpDg00mGTrhyluTkbpqIYT176G7n
wTKDLw7hMmh9FezZPqBCNi/4C0qeZc99yUkwjqoj8Bk0CC7VXpoz4J6Lb+9CVOgYGuHO67VPuZnK
M3sELPP2zoFFDRgHSmlIjTDVQ7OhrGqAqbvg+mEJiNpRT/SOCqRAHQ3YDeJPmBGaGtg4jsrnneP5
Jl0LRofxLR8zolQ7fOcsxfStnwLqfOFxIG4qhH6FlQp6tiHnerGHCRdhEJQxOkyAqoyv3bBT9zRt
gb8dVxGCkcSkHc+sDj3ScJ1egnlCe3mHojLn41kzYAbJDfPwAlSAVc4f+gMMFpILcyHXbv0B5Y+3
4IHXP59MUnQvf6aqjxZTnGDtBSHUCet5cDVIl8W5W/zI+SS1ggvJCARxS44ZyevnCNPOpjldT+IZ
rSwleM8F20ii4OeoJw1r7Kz9zNTXrXVu4IChESuyMOu2R4cUugM1GSpHKXhifwcEHuArU9VEhc6z
IBquSDImS7iuF0+1wQAiX/wew0EX20bOdwb3+lIEJQCpNmvJMi2vPjicWGJvqoEMGenVpzbz4su+
Tkrv2yu6C62VkB+io5EYHU1MZfEbWJPfatwZ1CFBXch1uT+GRTsAnt2+PyBohD5NQ1SdLE+/sFHG
KDC0bsqGHnshHDHagfoJxwPDfZjPWh4ybvV2yxSuZp+bflIo+mi0MBPJGY6zbuGx9ibto2W6Ra6D
GvUZRKgOcRR4HSLvh4jPQpbzyg4FAy/zf3BWXi37KSYbyuIFXJd/dES/SiLh+U5aPJkYPX1jeC/Y
aJQ4pQ+Fl8O+3h6T47zekmU9kOJmgNafoLaZpTsVdx8PYKB/VhOBx+eYxEuC1DyhYzYLqLsWmZt9
Z0zeUORQj/A+D77I6x2M3lHSQdXy3RFlyP/ClO2kNzrUNeMgdoW23wdMIGnRuRbFf0xQrDesU8ph
so3wyWm50F8x/Q2QDpGlNOfoqsStnP21OEOtStusrDPhV92RlNc4BXsN9uUTkAeVl4SUexK9X4GM
NYSxvjHEDyoGKydjs92XYaP3HXR4OrAdbnKZw08GT3K+bz/47HBAC+ym/YdHusBYNujAhjS2mv5n
aLgYjwva+83qc/gqX+n/3rd3XsGDTuO2nyvbyjg6V0EVp83dPqo5zz9vkNUGDwYE8jvE4Qp2RAfq
mn8pZJ8dgZ6TUL4Kmd7EWHPGPUv3AWupp5t5s/6Ly/UFXgzaeaKVHNV7iXEpJg4MIBqxb/28PbhX
NZ1cdGtW6wXANIAcuSEC8382SJTxeXlqK8F/BKVcZL0OniF1yMDtlY9VwI4NdCrIStCzvufWFePP
BYHTKHLiJopRhLRnQsvY0FAz5umfiLoOnoG0GIvZpAbhQUpDo7QfnlgDYmflQmO1N0EwEW2SwKt2
vTxkGVVHkHp2pFZBDXPSWknlzhu/dKAtNNY4Z2PGQwWMILogcz8w9lFZS33mN07707hDf5DWB/KL
wxPyVOTNlFEFxmRVFxB43cJMXyGfIAUWJ7FaLhodtmU1WY3jq4Z5BNvydr1o8IgbO1+m/hzrVo3t
xnl4CzxszkSGmLDc41a9TlYmhy9svkD4TouQ3Zb/gFY6mFnIICd2PZL7ChB4Wlp835UL3OwlFBDZ
iIcbzg4IZYOzffL3hcqLuHsvQ+Hrlkb4P9if8lIrt082kELaNvbsEucJuSLeO8uhnCTmykFYvQ/q
jW1+qxLTKmyaIO/p5MiBQmP2k55P/H+2spWikOErfyFmd+8fc/CYDHr8vop2zh/UnHW1rEsS6D1C
6byajgolVBVsUuOHZspN7nuySSiLpkDwZsvEMYEnEcU1AKjtBhm/VpJk0HLV/Khp2sYwR1OOAL/A
DfJlyfH/ES0f3pzsYRWOQWQjJs3FIGyUvX5j0ZpIL5CfiW1+LDPJXSegPEc9IvpDDsBh9rUlFz94
3q3So2mIhFrn3BD466waW1yWPg9GV583Dn/7NXQ5h+Oq1mYYTZL3gqFIeFD5jxuM299F4qTdZzsi
IZrQAr5ce1PkyMktY0+ULt04+1BZkGaUXn592aiH0MMzH/dXOkwEtqnlp1zedWPOpJJZV4sfSEEt
7ZPoh/NMMcF/TPKTlHu0mTDHhrTbTMJzn2O1p/shSjB8xSP+xs2hfSQ9nfx//aXrJ6beF45uit5t
VYz+fcSZYJ8ZZhDm2mXVbEHlzdfjW8ad/cvNWOQ2F1P1auVOoRnYPJjzMaGzVh7AF8wNvmXaXaAG
D8+PoZpQLzAweLuj7LnyYYK+ol0KcyJAvzqYoUisayse4pkExLU5OJ/C6FlTrSknbJqhLNrGae86
tnQVO+nXZnHCeU6wl5k6XeifM/tgECVv1myUMJm2f2C9xwCNsvBIBOVo4ieRM4EzdFO4AuLJak5m
Yh0ukNKIgNKmnB0agXN2wgGwyfJfLqE51qDyokj6vtHA6HLIU7AuSUnIvwReQxMpPI+l7OHD929l
OsmxkZcG8Nzq3UMbeRObMdkKhD8JHEi6K3EFixfhnSVYJPR6/9r0Zxug4I9wtJMtTk31aApLp3ng
5w8ua+iDdie0D+n/p1afmWP/LOUyka+Xo74fw5m1n/V3Rk0HEU9bUCM++TKKxwxgYMVSmmOW5fIe
ZJzDvVczA32xm3MAMLVWklRq5HsiJLezPi2lAUNxttmu4Qn8v52kGZdtyoIOMAFbkLgPuqO8GpES
c+TkpyQus+qWhJ6y/+NAY4bR+wXSXHVS6SMxolf98XiAU3S7EE+T6OY0NKBRT7lfkdQNpbCc91kd
Z3fYk8h5s4yfR+Efr+QOh5hx5ERWIcmqnwPP9LXtx1ogDgpSF2vlp4wnd011F3m04K2jEuYUwJ8J
WNczmrnnJcEP40xGSGcfezKlgkAWjOy5z+k3hUldjEWFczI+zsqeMlsYfVbalaZtim9VxBiFvk6a
Hh8Ot3Bw316D4ZmALj1490AgrD0YRVRtVPMYnNCEzp30CZLOo/jHTHjiNKbIMtJCTopGOfrEONnh
Pj3lgyHOLb+JgYXTFxGN3OdkVid9ljJdndmQyDpqswp/JIg/vg9hgLw9ipWZV7A7ZQwcqIVt8ll+
U83nfrK0xiwtcHJU6Tmj61+43H9Of2Y25Azo+w5y1fhvI0TiVBFDWBnxlPEt0e/GR7v/G5jQj87l
K8vjJ6Ri1mnRbEsTidCAWhpw48CkLeAXvIjQZ6ekxV/QG8V+XDMak0iVfCAmybkG9bMuKZluPfSe
cnBW8lzgLfwirBW83IsA0sEZL9JUfz2eavXH9A0Oz6P3UTVkMt5A7hNNP9krG3MO0qerrUHGiEah
dsk6USDqSc15LP0Bdcced9sl4xNF7OZZ1Mhrwn+V6ZW+pJ8yqOCBMCeOnFX4jYPGlgbJ6s3ZbRBA
I/NwOKoEwhXdgHC57RqsQW9oTDLxbxTe1IQ+wn8EYtlYvMMgT3Dd2jEGqgN3jjYs9MA8R+ZC/+80
0ydiBGHFpmDSPfwM5ausP8SQm+g0jHwP8Zhty4nG+Sk8gQ2i9hw5kv4JOHoWn+Nl+bg5tqt76exR
UMjh7x2+XJ4Z0C1gUFDqRu8hJIR6i//5Zg9Qk/u0ONl0+YZ7fIe7WvPfjg+o5yVQchT6Zi9A+3zd
VB6SQlkYxBZDMc9K2WkliZDhb/Jk/sobAJTJYw3ZA8iVxWwbeC00xLX87SZHq+2wD56Oocu+ELE+
IBBpY+QTomlhQzhSkWHIzwhQj8AtwaI6vVm4bKRDTNsjcWeiCTv8VONZ/4/mwuzIbacQiOBLHRt4
VkCVZKuN0nWT6ku/n35ftjsOxLu1YHPIBZE4eXsKJV/HIpJfXf4vZwTN7VeY6YT7Z+0qHH6aQujI
n1ezzdYec9ttYiz/KvxPbPHrc8joRHZzUgJYnYCIhuCJ4cJnplMRZgQYPhX2P+tvJm3b0ZkRGoys
Ia6NhiyqxNu5zaX5j1vqc2/bIq+RrWn9bxZki8DJtRDb7hcm82pZzKd6mN90EgXcJwYspRC82k6C
NQiBOTmJyQmFWpQtuctmmpOaG1og2rBncgqvtYPUdT6XJZ+icdfWNBSggffymi2efBOCRyFEg8cc
Yahs6cDMz2cmzjPX1lZQfBy9KO731GgrYzBSSLqlw6PggtF0cg5AEHc+q93lMrSWPpUul9MHGQch
/OPOOhkeukq8bqAMY48gqiF39icsH4vQUs6TOM2aJQHhDsGFUG3KttpYbStgkPIP5QxiRCJcmLRM
S59wmqZezWOmvZGtPUpBsQcSsGS0fNBL7iC6fumuRyBtUgnrD2+dIqusx+idSH+lpAqNudkS0CMw
tm7UPAaUdxSex4ygHjkkx2Uewj16rsQ52ZcGJ5c31JNfMfJsqkE+TwcxCJtga8YA+by3YxNEjVQZ
ubGGvf0KDGVfYbt6KPVESNJrC7zEgDLOhj2Y2oNwZH0mu/vxSb5NLuoyiQgdGsEFxhefsN03abss
SKRDFA46FF0phRKBiwqAjezU5m30SEp9Mp2j53cGIvAT58kpX5vBISxDxgePita2/g4bLknFrMHT
75jFwy97S+2/TCliwXhKrvV164tdoneKAFyWBnKHHr9x3XBVLXrhjZKAYgBD44DArgE4PGx9jH3/
KEPJ9G6x8SwKDPcDU+WTVZmboQh74h8gtOWVp6dfQodwp5D8/9kDGA7x855HmK6+t+jXLQv5OCTz
4fSBDmvu42PxIazZxx+fJBS2l/4AdxLRNNZOJphMAQ81Nd+qDrCTR8gCky3sLGiSlda1keR/G6Th
umOBkiv9iSPuA0ew7+FieKhoFIX6FCuNnmdj5HiDzQeBax7J2u7/SSGoae8Utr9NVmI6j4feUThR
9ruMGrAgWPC+JoQdEQYjcN+/SyTfsRL79Hei15c58DW5295RNtbCqmjai5oVqzH1ewv24HJkoV7R
aK0rbpL+FGhFwBYQLW0nG7CZ/O3msma+ziwlIkjCMfP9ykPQWmsi0mB4BWUZ0x8y60A9tbhLTZH4
Xmvx2MHnC1LGwilYIrSUzd0TE/xSNXzKI6GmbGC3lIRGIT9U//wyhpF1SgvvwfQKgNKiewJzh3bV
6p8KwcRT2yWdHB9+F7H0kDf4/NuEGhi3yNZybESrRWqcv941UE42cQR1No4AOsfjMlvOxrzsfJBC
AveqAkCb9Ny94Uif3+FzT7WSqKnYhkJar0Jm1lRrzw5y5xQd3WmPbWUaJTtBa9eSjLfp4vVQ8Xyp
0tdQL47fPGIgUbxEmjXIZT44zGM5zN7EjGbChUE4IoXaX1JvXz45kKqXdYbOG3LrB0dJlvE559l2
DvCdr+4RrLoTa5pRsaivWIfKERjcYGBHiQt/0b4M/O6BLNscvQtMGcWiS9sGq79vEuUzC/vEHx7/
d9ZwHsgH1cLmm3NejuSxGZeGDJCqzeaA1jdZmFKe/L2e4X+BXgPAu5aBk6QEFbVnjr5s52g/h+6K
fdqvn5kQLl/N0065mK0A6UavBbwol/24R6WKN8O/udub7w5dyoPrxvUTb6ouaSYShs0y/qVkd4xu
xXZaHbsIgsaRf4Meb6RS25vxYcwpGfwgVU78miAipAjzIhKS+SMmO3/11TizXa8yc8j46h10B1vg
D//aDQ3nzrVj+SFmeRELF+1kAtak7zejViXJurde2e6PtjOH+53u7tQkJKvKrU0ryz3FIqBy9SlF
Inm3sxrzWPsyXz6g3R/6fZayOkEWPEKUP8VHxFyktECNyCsjq8YtpuVlT7Ppoc6XqW3FcExGNqQP
gX7RgGAp/NSoXzuNoHXJcAijVUo2THI0XQOfxggjmmill3MdplfSTEgv82Ek335xtoX3Ke2Bso9w
+9DAAC5b2jtALEP41qv1MlWgXydp+zkst6BrbY6DTupXb2P2/7sGZjCKPY2ojsPbHWUyKqN1wpxX
GUAHfe60cEPYMbGHhKWM90CGrkeErxSzBVHChvk8qLdose6xJYgVamnlJaXJHyyiEAqOz5KY7XXi
GV7QrxQcB4QYwBZLm/BZQNtkJWLdX4pxhVanVcLpIEEqD/cd54cqFWcYFiyCqWF2xj7T40jLEjkf
wSWc2T7H5LiKCTYb+34bcruQza6FVO2zyd9XNtGJz+CZJI9y3G44njVDUq3hqEht5lS7v7/lNjgE
IRbhmqpApsO8jAfi+KhRZGZZrHWgPQtiw1BgnHbDaui0RbcU97wUqMrB3HUwYdjSKwvnbxqJ0cTF
duWhnI0uCDShi/pCtUWHaZqJzw78ovdUeoBBpKWniab563Hsh/t2nD6NwMymdrRKOGmzO+U6rX5T
AmfmMMcYA1/+LGBEH26d1ecu//KBF0A+hva+PhO3zYdQ8prwxz0s32p/1CW68t1bVbIWk8bSYokm
vq24w4doJFmeLEU1Pc/8zoXl2sTqdyr1TrYpcSQjAFUI4xdh1rnR/aEAx+dF6LAgxQgeh5B2rsIR
NY0q6OI44oytwjcP/LkhSKrzfs8eStB2JfG/9N2g44iPsg1c9Tywjg7nDDin+eCy53BUQLSkIr9a
a+qKZVLs3zi6lpMCA2RO7SlISoo+rffApPn4KyKXndMD+QrlUKTY29QfmKmLQXyR42duvdCHzUxx
eysjPKMdfZIldCSzbx1hXhN8oKksgl15aIUxiLfni2jAIBldaQhFgJlqYucUXYYTxoRqyWDphPzC
QElvpPD9/3rTqJnJBQtGz13DT2RhmKXjRsMAwS89bm6SVX10E5+mlwnxnPQgxS2l0Ck5dAzsl1Pv
KNozYdY7oiX/P5vVURmC2EZoDAzF4LaaiPnlYdwnmGhjslN4KVsRSkozz6Woq3XM8OVkvlpoW4ZT
3rL0gP11j2HEZGZpwpwkQUlOqmrXUItJHCJeWsDXSB7FapIut7eaF6mEezsvl5DGvuFRHL/3Je93
WOw09piPiBoPb49zcdspUDAOHwrM8rKpuwoa4hlm4hEL7FFO9Lf4Uhr6C3Uz7wHCksHxzkQWMTKd
4vqeRofQLggR+MnHwyLFvPnJdfknp/f6oiZ1MCKUBHEkReUtyq+wEp4nOcJaxbSsP9yPCezqYQXs
D2gRA0lVkK/nMkfbMTsnDr6+p5I5fFvZdt7A9SoW/nSzNz5Bnx+ZTBv7j04Kn8rwUcO2Wlq7Ecwv
tcpp43ca6C7GgQ+DfWpkJo6Ku3gU2gEH29eRIwTOT0Xq+LJfIdJ9PKnStz6rfWdMDZHA0i4jZ6gu
NXVE6EV3sHYfB5xPHNqz4YyxzIZGwsNcN1o9tdKnuUrL1XPXAGgkfgbw0QrStr2C141sYx3tHKZZ
bUYbl145vDigyFhhRgvM9IL3VADeF3PioDFeLqrynEwoadnRB6D6+3Ekxq++RV6y2IHFi6vZpIOS
4foG7npBV/6bQ3Ed+vs9rKMC1kdikMGj8Vj0L1CGe83GtBinuQ7TWVUeuWgLUo9b1dLvD2N4yJOA
ZkwRI14QFg60L4bd4MnurNoPxD4yQx/RqWlUCY/mz48SYdxk8acSi0Ujb54zNq1+YW/ATPbT1DRn
yWtc6uqqi8gFDpwERUzmhZTl5M7N6H4dw6DF+VkG+O26gSrlYrxJ8Jbx15lzPUCMye5j2Uq0PfPZ
FW61fZY7WoYmRQFqe4E2QRaD3mYl4LQ0cdHJgE4+wubwURfwcwg6MYIvr0BTJEDnwE4cu09hCzuR
+EWB42JzQlPOP6WnwPiI/veQDxVC/OS+v3vgAcDAAROEVOP86tb659tl63jwL991ke2ickYJ9rva
VakVqV0oEpSHWT8DJLVaideHXBDmkSoV0JkKe+PeV1c4YyFPoC9qroaZZlSCMy+XHt16BtKSqnqt
30JWtYFKA7du6C1a7aRBmxcfKA66y+1i4/QVMTJIB6QqaXYtRGucByzUTctSbc/dP0ach9Pymnkp
AuIhTh6BKiu+TFRU0EZ84FwmwwSyw84s9XafM540s8L8O5X7+5pskjCK/Rn1PBm0pTuuttLOGK7C
Bpx34w/IunOMkAmUHXjG5JezhEuVe80QiENAXI68+96o72WOXNjoZ25AAqWLhZwOMi6KiOKQ3an9
xNDZRTvQzLt95V4M1scjoxfrnyGYfAPgG6wFI6+HtGM6n80AlaM41FW/8gLr5tGavMu/ZOxn7qtG
F+mzz2Qc1ZaW/OstU8bmOfV1besNU/qb6szxWxNkGZB0/Qa0lrv4U4hHFoZ+8yBhATPph/LdVpMO
RDE+jjdXiAUd7HQ4P2TnGyHB/vfxu27rFmmr7GlNM3tdivy2TQXV2n4tdmFx3GYRt7Rr//2KqwHw
gaAejMKnHuQI4QqG6VnZImsB1NfPcco1aoXNvA9PnDtJ+d7B83bs2qc5qdoOnRw+DfzGWeMryQVx
CAzdH7RAxKFR6HPKP6iG4zct4T9xWjcvJ5tGqvBHXAd/4gwne4cJcvBDTpJdq09fRs8SnwUfgRZV
myvTtUoB/KjF0Yd546RwXpT82fQQaP2aRcQyHzHvc3It2vCLQqGPufnUq2mLqaBI83G/xFz5IMzp
7kBf9EE8YguG3Rc4LHCbEjmuouDgBN3a5MhwkDDRf1lZLrS0Qq2HgS5HaPn45gN5qqyPhF12Hi6p
vmd5kn731JlT80hMmHRA9U2ElNK+bfXUs644pQsUubmoni+kTyw9xrNJmyteyB2X7/RjpuUiq+bD
EcRUXlAeN1GG0l4sWgGvZEe2QIiGj73DMbgK+qvcJu9KoOXA5i9CDLbqWvggKr5Cq38DT8ca8uSP
L1hgKbTDhmBeC3Z9Mt+FP2+XKJXAjyUksrx4NeQJTGfu6YrdkQI98/tCgpb/UAUpT4Qk+DdXXdZq
7179YGaRWHlm05eI8orXtBFSKMAt0ns152CVPLAUJvCwVVMpnS0QzwExj3oz1XOqr3a1PvKqobPn
gqapfyXZORS5tkeX5BNqpgPLcb3jnONDPeQrXACUTH+0Mc4qFJtV45IyWSnA2b6+CzV5GzblNxBW
0Jg5wmF3qQQDyNmC4+hIP65P/NXV01BmjFNcZ7O6NEFQ2k+NDqK3H3j2kFsUfjbj5PZGUsJPTSIJ
j73tpIdrZYQIu8QQGMEQFgc3+I15d6adfJJo2eC/TtkTemOJ0QaLdkrhWsHsV6F6JXn88Jm1YCFC
odnQj7jO0UxH/hw0zeUf6T8ZQXMtnl+3c+VtbvrSnLJV06uIzg/Ocb7jGIhWwnhyRofTa7E4HJT1
bD09vF13y1NqwbPFXHxNa6vJ3eYii/FjAUFXtBdJj6d3Duyih6n8Iva1ENhe4pL3B5HBryzBlttR
yQE+3eDU1lH388GmnZ09TtCcKhtUG/+DjoYn93jBnB9IIuBCwkadC14vMWYK87IWnCZRvi4b4wCu
xeUd3p/W22+Kc/YE3epnL3HCy8PkYJcPBX0FpE3xt9uqkPnMadmRn6TTX1p2toVumnvVmut63tWW
L1Jrkm6Tp5DapH0sW9Ms2eMKsWmXdfw90zvw4JMbqGcyfv2DiXLHYJTW5CSk2Ag1+z8ulvQdl5DS
YT9f9zXn4ZzxGPUr6e/716Y4lDOKAdF+B3+pEhp32yjOAEjEtxpkKvkBtJmxZ9nQrZ6acFj4caTt
nRrUvxMe4ytygvFj056jt5rNNCCw6kPBLHlGYZaJqMBHQFXK9gDlTEIhduKGF+vTtk0vgFh8+1gv
5KKNWA/upLYysWXHARbFFkg8dQlbDFS9/ypcqyDOcP5t4I5/xU+8XYMjvi/VaNngs9n+iD6RUxi/
ZDchDzqAyX/wCmIkNHQ1YZ2TnXLokcPRy6oq4KhAEGJ/Wvu5EryaT8gfc65pG1L0RyB5adwiHep6
3ftsFkWmqFw7bD3u38IamsiP5BL7z4UHtjdjiK+fOyrJmjYSGNH2TxEwnHVRWND7LSe12w7rIEll
vkx95SxCz/7gm7EqG9k1fC1EZRT5qAGtC148BEYZF3SQd26QBCkcJ+siUamdq2g5CTb2eocXhUwi
z8PCLCQJiMsCObqmOBSHTkpqryRGnYUjm5bDZoEjNN3mxTcgKJU5dPONq1gxNtyz0x39J30MslCW
4czoKa2WCKfDMO73amr91P7dYGBBeqRnGsFe9SQfyYTBMtETz3GSxqiTM1o4j8DoA0IQjdbyXjLg
e0n6tCmIQy7EVkG1QkxR8R6kbX/UJZCQSSvmnJVmQhqXan6GbtYJCxb8zpyTwrEyRhEwkvthEfI6
FEKVkc/qP9dGYg4dTQR5QQzEikD4eUWJxb7VJqJm6PdPChdxiqgdm92J3SZMpXOsRHwrt0hLyzl+
2OY9R/CEKsd3d9w3LcuVc3PR3eosqoahcAbvrRpyzzrYf6gQ73FpHH5Mp6mw20ksBz9bnJEcJLWo
bFz5hI0kxsm7gjz8xlWFon1QxT2IcCg29wubNeypvB9S0ConzBq/UxpxEygqDJ52Cmj8ve1/koEz
BI5oa+qYntV8Apltfw5oMptdyWrjUhETanB5i3ELh9xgP2aVDBX8No7FY5+TqFbFN5zJi55HbTsb
9eZQl1DElKFl5v6eJ1hjHrDQK9Es3zPAYiMJXz+pGAp8pIvjss/+uP3ZiVsND6E1aYHEWmGxmNYn
ey16+fk5ql2sZrzSCBlK0or3a+fgC+CSVUCSwIyZrwuI5sUSsbxTmeUchxdqnVumJZ9aeDGIXXOw
LgXVkt29BAknXcAJsQ2nX3ZV49n5UQbHKuXjRFsog6Op+8mvza8b3mWJVuDBilwDGBC26K1Mk0O6
iJUbWHOotNCAI4YdQy4mkHU13UnZn+HwfhtJ3YqdaJnTWyryhQMpMQkQOPWEjAa0NBPI6foXvoFP
2N/QRciW/K4C7yVLlKuX0j29EP3jZrlHeXIhkeYVGOdl0NaU8sJh0Dc5hTg8slNDRu0xu71UURoT
Mp89EpWVby7GZCg/TveB02lNcZfx3rPAF7BXXQrmhgBtulgqBQa+uNBqX8yHh70gKAFawGps4Ze2
T9S7bl1XAoMiK7kaLDP6oU+nTPKKX1+t9o31ywU9diDoiG3rjF1UPwFen4e36/uaZmv9un6g7pEk
4ooflBdnZ/jZANZGaZN8R7FQ+Aw1fY2xxJXQcT8tY2C2UUoU1spfXpgmdHf5YaA4UaeOE77zX1YN
3l/i4LxL2nbww7TO1Qvz9H9xufu9JIGPzuIYhh9EjHqIf14GA3jVnyqySp5RU+uwnyxOqemZ889Y
MqhtLgqoASX4OW8MgvzrKMdzBBiLUw7RqJpVFJ5GHV8Xn3Q/k6QQAc0sLXi44f9vVTeGolMcfsMI
0K54gwXAXQW/5tjswONYNyHNlk/7+f+8tWx7AuKrBQkAiedNEI0YAgaAmvv4UK0F0JakRHw4SBHe
RYZrdmGQA9wXaWxr2eKNYqR55c7ewTBon5FCes7PSys/UZ/j2oI9Ix/YHA9BKDUcoUXZsMF9iRPo
rCFlOMRo2g0ixVmNexE82psxbDdlM8fwrgaK/oTdJLuqj/FdYXGyk7iKpGfGXk+JASMKVM2wzO/g
zd41ubCUTJNU9ZNiLUq91r1OxrVXtdfFkrtf5m8wTzNfyO3gH4SOfcXYO5mCFNI5QujpWW8u5nzU
ZNDVzMi3oFOTgpI9bKlcy6Uhg80PTM3RLitQZEiMYW1+H6S1xJ+8O6PmTQJvLYASZ4JyFaLvdEs8
nNzCDCJTlaLDrjR4hP3gsDnBfY53mk3YN3QJ/GfOYeJdHvEOI5B3bYrCL1tOqgbTxoHE6jbXfzSl
v7ukg0Vp7R8mS+2v0NNOO6wmwRkg5wk0vxocCS2nmOFV19VyJbHUN6dv39kxCh0gQvNU2cryOhTw
SKsLj8TX/HWA0KAIohKcUdSNO6fixVZOKHXhE9Og4HJCwRSPS4mZtImF0nnqOdvM8hHYv/KeTWdf
Rg0jh2IoLy/najCIksn5oW8BsdVcjYXeDudfJCQ7fz1lwY4TmP67hG+KjpYAUBoz9YJXhBNTZlPE
bHJvD8SJ6S6VEA0aVokPs6Mmczi48HVo50i74yLUtG5/836lrbGf7lrz4580pS8tQFTOGxTyaUUB
XglWtRBualC/8whJM3HeGGnJGLwvc9mouERhz8fsIPcESH1xYZU0/OQYOqqMh4XUn/tlbgLNKjVy
bgknCpb/s3hgLCdQWOBQgzS+Kdr09ir+okrxpRwYX51c2BAZX72GE7twajuM/AdUT3xtWgqDtY3l
M0boDufHqQpCForczzhxKoYor7qYQJHVffb0Jq++dndr5Lg2w4c4Daajd/VDLq7hD/sNxl1DS2Ub
g8hOacxiF1SjJFcQfHsX/4gYpG5h2p/CDq+p/h9tRCzKt3Qk4FrWAyjeSIngERcbV60005VaDizj
ZQVJNchrufZRK2WCgJCjBflW4EFI2raNZDXBBC1zBQuxIi0yBeiNr1MgCZB4UD/p/mtSHcIHRq5E
63jVCPn+CMQXzie0w6d8mm0xrnKR+mqhneabGAK7vr/vb3qhuH1If7wbtBCwMDdH8fqw5E5nS0zO
i9I3YiNt4zx7wZvQ0PqX3s+9IMw5FdG57U64Vm13HYFQjxCbCHKa44Gaj+xpq2DwAFY4b/lxwVyS
ilimLZd75+/GqybwtA43RefpksnenId3ppVFOQ4hw7SLLNW0+HfeuDeQ93/2gcWHW8AxUwx/TfML
FZnzav6LhSPI/+0N17PFGiJ3C+iL5GKQGXm29MHxc8WB++5Liyjd8+NAwBur3Xjhdlqz8c0tvTYl
qUc+rqbwMg8DAMQTTCZL5K13LRKB/EgRlfSH2ht6I+xU4Lej68UoyOYrpdDny8V9JdK/oWbyjDcd
yZEWFQVA/YXZGJacElipPG9U1ok2MRJktlAJvQj4DkUEAeGupzmLz8UvfENQa+3jaNG7tgi2AuvO
jrtKA5Gt847KItJhHrPK8dTo9g/gaKJdIcIfkrqxcwL4O+pccQCnrRly7+PEplGzdqM08hOFqi8k
2CMOhDYA494EW0Lb3YTi1GPdDUpOieJpjYDVX123PJkwj7VzerjL8w0Ptb0m/FpTh1nDPyPX2YmA
xGsUfivy+UZbKpdur09lgvOBqWZ4Yzxj6MIY/r34RycjNBCqjd4sTeXMOKYlyFxdass3314QbwHV
jWdgkRdYWDDeWCn3Ynre/gDdgPzDnxzizrbFq6cqV/QDbYmfmYMPgNwIQrIA7ZdoFiae6jVfYjjC
FSbRLwaB9+V1XvfOEQiRrRc3wXrlWrvmiC3dxFqFUdnMWoxV2qx8U2iFJFu3Jqocw95+ULT9MbNh
EEgNmj+8UhugXGk4pE7f2SLrlpsoih5MJtE68a8f4rtw8z89EXsRVQh28Nk+3qsyVrb/OFuDIrEN
sHzQXhhNs6dcyhn++OZJKu+QfG+CPUUtSUDjlPAP9bOolfRELE88FUDqiQvdJncYT2jmM9d8gKVR
PfRtc2CcFhA/V/hlhO2yS+Ihf7ouCPUTItO5plFYEhBki+aArkY55XUZUzBsFORZzWp52Tuscb7t
klpBEni4D1ppl+vDFzfJhHTOF9aTeO0u2wM77pxkaUncpWcWU5wAWjn/b3O3IDHtxGSdT5SmWzAH
PHhXf2fzsf0xoDZZuS99/aGNtNFmQNPzePaTURT+DILOeloG8cihJYBPgcjrW5cZ8Csu8kROqcew
hV5+2vWmyhuOw1Hm3vxU7MhdW1g4P6NMiQmutY0rAO2y6ydX4kiUZE9yTtkQLxH2FTGtanLrk5kD
atyPx3uj3nHeHFN0ajcy4pTA+eJmdxtStbc1IKvm8iFH6z2mH4XCMt3B3Syee9E2x8a2rG7Gwzo3
qpfWiJK6FagQCxS7FOG7C8AbQqjy+j6LTFAZKY+a4YQviLrrbrJCbe5oG/dn8Zwy6jyj7+hH5xDA
EoqsG3BVy1N6xW8t4pRU92LhtfQbK36+MpTB0DupUtX/p6VsJx5ap8Ei6/Ur5WFOsFh96f0V2uB+
sakKTpW05WSw91PX4VHRLgo1JMNkBtx5lr9pA8GTW7hUOBkEhb6a8pcc9t1LQDvEycaW991sZfVa
xUArzApc2Gsf+MCR6bz23jU3ToEWeV1TXUlR/1LH4MW9Jx622oKwPzpX7glxj2MgYDldC/QkOfDr
JXGRYRoU5nArH0sRhSyighdXW5ibRVYBGokDGJSSk4HrAZ6OhLfM8UcXAfqktbFmo6dsNQtg9oHq
4E5oidB2Tle7dd14hr4wInGL2+pag2P452XT0wVQgDgertlT57yPHqC2nEQhtdxxNjNDY0RfpEAd
0rTSYYQt84JgwVysvwtDL54J4jA96gyPz5DGX0FrjdsjgWnXa4hijSKQFlaVoN5JYbjI9a2HRSLB
MLGyCLG1cTFGUSMGhkH0R+dW74u18Vyr9EVamsBRNOlQ2G/y2qygEgKIo9pWoWxDPXyPI7PVp49z
aqSp/jwK4ybpI2/upKVlBuhIJwzK/n4IAdFvjTJXxbSh2rDgg8GIONN9cYJrOAqp6EmChFkLuCk/
iH0zZbjy2uuwRKOG5yfMTTy38gbXvlldG0DUk9fLrXqP/WajPZbDwJRXl787K2bbd4xdPajB2yyx
jQA2fQG+h3aY5KNo36CbjRzhNQklDHYKVwZ3wjL41ugIX/FTaiwXkbvnnk+NiI5X+sO2y6Hcnzw4
FsPha/KTByJWety7hk2WTBUI9eeoua0dUH2hGVPmSY+kB/KFw3wTGv+xhv6En0kwbHP8P6Umk90D
bjmceo5PqC04jVvIqZYsEYi5mb7xyJYPP1d46SD34x1v7RY4c3oTqt3rGNe90kDG6sJV2ejnq/95
lPe3AQUDSV3pObvwTGkjCtXkjAaaOthYeO+aEZIg8y3wp+7M5Al8WwyiaBgQeAtdlNT0TBRFaeAT
eboCKHK7qY6m7ODVQaBSRxlMom3vHFE5qwxBIKIyU+U0YxLHsI3DwQ10EIH+rTYLXN5vmbymXXeK
hVELWw2tvFwOhHz3vtLtIZWn/xvEWloVtgksdxkrXKDzJLTPiR7eD4r8uCenkns5986iQ17zUn2m
h1qnZx+sZWFhAroESvesjCC03vXfwUB8+4u4d6+KIe3QypHFWoHXkxlzWLrl4woYkd9WI4iJxitI
gLgVY/sXTEfV3ck300hRAoYsbvl1JGe6nnAvCfe6QvYPMgosvBoQKmF/dwZklwoay0T5EdwsA4YM
5K8PVf7KtQsGcR5u+woCY0g35U05g+SrJM5itxnZjncEnwucPvZkoolMEQRHUtTMjIFz57gFs5cZ
L/Kh2m/Axv/xeGdXtkUkbuI0/9uquatV6ob4s7LIu74YZoZDyoN8kiWEv7rgiE7aeF0KLDlLBGyu
oQI64xzTXcb9R8H1Im98xnpl4y03Su1r7NQhGkE3hA3RCMqBG+8WEwQComZ7czD3YyEfLBfkONHD
hJ2mOgmGs50/uyHkeWoc1ZIpycSLh+rC+PIbfqbNnYGV3ZeafcvNL0qeQC3qhWREzV6F/o3PDnpT
wAnPchIAE6PtgDKsDcgPxdlGbkC+s6bo5clwBPTeAqJkgD3qtROqt1gyq7alpRo6EzaPRQ8Q+V8t
ylfQJPeYDROuXsriirsNKoH/GVfwtEwieFGfB6N+7l2FtNXlM3jb87uPb2QvBapRS+hbMJPTZA1l
L7gNoeSFcnj0I4sJghMPxEVwdns59/dJpol2j5AM6wHdj2uhQphFANsEjGVSZtV7BJWZQrmwwucP
JYUzXTULPYoj+dRONoo4ur5tePE4M3JBWstdThl9/Sg6ZyUkZz5h7WfZ8D1NNesh1m3UtsZ8grp0
82D5rQa2VOQ+o48l8uiZsy2tj1c3SkfHILLSMxGpe87FFU6yiCI6ft3ZWAInf/Nt6B5rhYfc7adv
wq0Q2bcQtK/BtTjMgc85J2Lhqay7d3hJ4XJuw5usKS+x3iUFIQHUWBfz9wMfl2INspasH6Px9+CU
LeaJfSk8RbHQl43OJAPD2iPXN7ne6sXuJ+ZbPOycWIOawEBOBBjesLUY0/ZBipNfK5eOzATZI0oR
SnL9Lbe8FpGo+XRImUShNDSt2dGmnK9JKy55PHLswL2qMbcj6bYJFKZOSLF4ZPX4m8IxAUs2w8VF
DJNQ31H3agqUHf+WWtGZRTAk/OA15cluLMeGLgO0d/VBNFo2pNhdh9NVW30JTL3fWfNJYpW0RFRj
xyRm4vWyNF/2UDJknSUBxWH/pi3SNp8QAOb+pR5732KgFs/w2kKimHYZAZb5sS88bNxpFQ2dqzA0
tLJJhpw6u5WF/9QEwkD5U7Ugf2bJpcj/65QEEf/9WfOhOp6g31l4BRMp721XXgNpnYTzGxnNoHv1
BpVZ004WTsoFlYyLystlj8rkWBQYFVOKOGdIehZ+/3Ipdd3vcEffyx6rjy/3W91HgSP8gfeplP6d
Di6NvET4cT/PcyglQltNUIkFXTeixOJcnQz9N6MMc69r21AHSmqelvWqMByIvgqPW62lPPfo5vIH
VIReYrFfAxwWFDRL1/T8KkPUdLWJkSLLj/lKDnS1q35PG8YSorqqqzRqSzCq68xH/8ML8HKbm+Qe
vD+6Fa4URPQWKu3JyQMTSH96kMLh5w+uIDLb/eeHvMwpSrgxzjyk1V4CA3Icot+Q2tkYr/7SI/aK
wG3WmvueMvqvt1FjSEfQYg7y7fOx7hv8UeRRH9hgkHqT9t1878njY2uEpfpcmqDA2Yo7L6y4ue+7
yXXdsjsh8b6as5sjtT1ipGtrMkzZAkRTnnO87JwNNpGjocJhYzxGKMM3lO0bd/J0g4PWtW40Qh40
xRcANoIJZXfYvvel1GtYykysWxxS8eNCMqbLOj7kG2jX2LEtqkhK5lmhpaLixb73tQdhwgU+Bm1s
5oIbZGLCN8iPl24HWfuhLFwJ8KLxKZcICB/8nKtK9MFgkP4/cw6+Wk/AixHmVG92r+hJr0BNCCVI
Y2i0uhTaHJHLZCePH85VBfqxcI1FAjCApILWfJKnLYCMuArRuNyAYgSva6Wg8i6+vYLRtoWxeAht
u5Bk/hbNMCGad9VwBgZ7Q6V2dUZUrsasNhK3YSSZECoHv4uLQ1xZLYJqpRBJCzeI+TkfJar8IUQl
8dUf87UHuYExikgauXzqCahG40P/3Jc1BJaF0tDnivlvCCcpyfjCM/eZrY68jzT+scaWO9YyRvAy
I4YVcrGmMJEdv/XxGzpK7gWjctW8ks6R3JOfNyR6PfiCYXDh4+OoYf3K9xkQxBeKSG8IE+JUAC7f
lIFGjk4JaJ1xw37hz5o27kDFkrrWfgX8paN5UKJRnkMuUbwGbsV5eO7/m5xs6Y2x52oYb3bgDAg2
iyR44on4O5gFsl5b0XdjidJINriBllcfiKaKKmH/SxUH7kev73CqZJ+eDlBi8k4OafUQhOX+R6uA
y5teEZ2xThf1cgehN6fWyjCSoERKBaSv+YROmaqxrvh7J8vYtOb+NB8y+Bgv8S0QptWA5lwkywp4
W/245NVInp0JqQFfc9tk3s6TLU8YK2ejmpTBrJKeOgFI1DpO7X+GgeQxZix8iqgfgRU4yDw+0tWS
6vOK5aeRSWur/OvjQxzXRYHI01zu1KLQbI5dnrp1EUu15U+0+3fWSw1N0nPapUMvn2gXp498AvFy
jPejC1SNwdxe9WvKaUEGrWGen/qaVcFjbd5fOUqwK6GMzy7i7IcaEoZswwzt7Gb1AwuNSNcCoy7F
ReEl2QJ9MxQP2XUwXMOd5GhFER9nfYUHeIRWnF/A+HbkbcMe3koYy0p7VhgaNbahcZRUE6OGIASf
vr6klvy4F0BN3+OHuhlcylh7lxDH6vJoHEZJm3CMzJYSJq5KmsIWC3NPeSszhWmijD7GpdytuLPM
tFdyYS3FY2uFymtKK/VBGJcY2gl7Q58byHkXSJ/3kL4H0R6Z/L8pF3+8C+A00Y3pq4IzxSBAwxCu
wgaglKMOm2bQiXbNAVCJUizrsWOdf9tgOQ/F12m0UOHqyThTMRxPjCZaH8wkZyQA5cqbJr82UGfa
Z1ohoFzkoHVt4IJDzx22mD6qOI2IagSSayMpKnGfHCqcnnSr5941JapH0hw2bTJkJuLDm25d6wDQ
Ij6DnMwrY+YOgLx5vMadxygkmtnBqFpyo9tO1U8u117d4n4Z3BUM/h5Cq1PzUM2Rby/cEXarf9Ho
W8AB1618G/zPitAU5cFwytQeNPT71XgTgH/7a14CujTCcxPNx4pRACYkcZUutuwt26jJVwzkFeWW
N3qQieRAWlgD2O5ejaXWO3lEaDpoy7CCN2tsMuD5BZLL0jY2rDImY3GJdErMSqc2XBEkr/wLuFQP
8nonmtpsK1Adaw57oMelH+NW48YL5THfuZW/M6Rzw1CPtoPOhegAPBtX7JdBqVzSkugTguf792sn
u+3k3yWnnUUaVHcbfcCd5CnFTe+0qZFDmPmIwaesUGp7IKpuK1E+5gP6g8c=
`protect end_protected

