

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VQBfeXA4hP5orKlsy+AFFAe2QBxKheQVMjP9iwMw/NM3O4tSdVMF5nSpUCi2zqd6Xl/0+S5YrDyH
MbW21sN7bw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NYnVtYYKs1fo/NxKyeagmW8datCnZRNIFQJ52Ut8vKAvoM6z9G59Louyi6BpOXJlK7hkOA0EyUcq
xnrhn5QTbG+/jjVXTRQq5boOLx13BVtwMvklEuJLJaUCJSI1mkPVMU1Tw6P0C7fzMTIVY1MXBSgF
huHBAAQ6j+Ca7SHEJMc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UdRiCUwOSibQJYHOoWlsqKR136XIPiU7//1vC9LO+s6bwL8gocVodj06NRrITDP0xKYK2ZTek7T4
6OlwV+xWr4k2Xf/sx0trTcVrHoE3bps3QkJHk441qMX8BKjF5fCXU+yOMX1xkQlvuWSD8+NvN82l
uzCDbBA0KjOv/IsJg1WHwqG44dahfC4qa2RHQtygQ4MsVR/PxcN8lnUdpguLi+YyGmh9q+fLgQBq
cNHly9YC9ZC1urY1hg8yqWcJm8AuonE47dIMtl55BTxzCygZ9uoRy68FfVsLU7NHg3O2kl94A2uq
uulT+/Y74MIANEyVFkVes/FR1hhgCPd7uNhwkQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tQM9oFLCOLGigsR+dGte9FyrpKbOg0a2HEe24uc9a4zzPMiWT4Zq+VUMyysv3hVDjsM6Rhdx2y1P
MMtJydYUSv3+V7JQyYwaG874Tc20f583mvfsydp9rtOQQwZoTUUdaw84/pibQ9geh55pxtJYjyzk
ltK5Hf2dDqQ0W2qoU2o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D9jeI9qTFJwFpVSxwOhVsb671/UONJ+BqwlU4oe+K/dJiOTSOoWnMaaYQ9Sgy96AbPfvmkY1YYgF
jNHbjBYJx/eNgXJH2lhqUlU4xX7po7K9tZYQraj2oMsohZUwz/eLwj91c7VL5ZRmCXaHh3hDU0yM
tta+u+KG7UfDjSpBDQDdNd7gt/bWHfns3Zj0BeTNOQ2o2kTzIQxImWuXKku154pI5L0sF72lK31n
Ls7v+PzriYFrSA6JTTtqAnDF5uCY0O6Lpa8FB2AoeQSutIiakkT+T39fToTawon3SeQIsthaDWDT
WAem4lxQFA8q64KvDBTwguerI8Z6/8BM0gLy/A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20752)
`protect data_block
XM0eT9qyMg03J48hUek7nGUORlBgaNiGmQQUfcSkUD7+RM2zBFCHv09oSEGRpVmldMzGZ/+3/GVo
tEPdNivIHyvjX/o5Nwbt95NPbOfeUO9j1DEF02L66ip+eSh5OitxHzPqWoyIJYabedjFZ9vWVot+
SLda0X7jdj8tsxz21Kz4+8Qw7Cp9Y+w2qzqiHVE/Usfs0vk/iXQI3STJL4O2tV6P/WzPavbsSpUF
8YW5/2gWyjmUZtNwdXvKIbW22oQIKmh8tKHZPuuR/rpaq5698pLSVFjxV4+W76iomybJYWObLsRy
zv36j7PzRLKmdjPV833LGW4elWXaOWt5c5OXeSAvadY0zuHO2huADlkJYCbFjRP5hK4t4Xk2PiXR
BsEihFw27OeSfzbxdZKl+Vb72AXKxoG9nRhcZobhbj0ncz2YjFcZTNHq3czaSMSJH3mh9DrmhXZX
nxDF13Kbd4IUUlBILUA1grFKis3bkXN96S3hHCYu7lQFm+3U7kLyhvFZzQCj3x3njgiysXC0RNbp
S3YSBToMqDLqFQNmkpcf39hTOaiXH7M/fFk2Dj4M6sGOPZN/Mx6/NP4YEQFRxVM35H2zVeZVTyPD
8zAnmsfSl4Ci2os9Z40pHh8RU4F0sWVoQ4/t8ArKZf8j/aMeEEwd6iKuGhZ7fo3RrdRRPXFtoqTw
QwQY0y2Ni4gyjqvQfV1zaNdPydmf+C/7n/JhOzN19QkypfiFAEe78cZ8Jl0sk4Lq5wjSPK1vBqLF
9D8ipfnD7XGXJ/WN4JTL7nefBF3UEeKjuwKtcGia7eZ4eT8SJLQsaqEq7cGCG6+E6POJ3PLhqVwh
h/DhZdLzHbf3Ep/JwT8qDt3zkiQKXctJuDpkIJXciRnbpOwNHebqy0I4GTXje6Ls1mcb5kdu5NTx
vgcyNpQaWMIEdul5NzSY6WbzLB1wkFGB3Vk87V3qiYBBnduESjzrl/fzDMm+6vf646e4PUvdJVrp
uKNhusY2smtV9kfKqRlgzlLxnKv9CE7ygkJCJOYmItLGZiDGZs7bLW9DY3i378R3x9oJHWBq/iI9
ry3kCHoXjBEzjHzn28tSrNqQ0E0an4/TdaRdwxjxLOffmJJ6PCt+wNCqgsWlWT5C0JzhIt61aoTV
XfFC+sKKpo8YIi4ts68vbYdb0JvqMDFqHdGGIsvcnY5QTowmzT5uF8P2yJ3MZU0XjJmhaPGvUZFj
ISOY70UCMMtAnckMfAi0CqZgKwlohYhO9VGMQ7FkEgqYteeGTCyk62Tsu+eBdroqXTEHHEF9FZ1N
jOuEVjSKZ1mkj8SPwUkA06mq0lqeUPuwAZSqTJ1lKqS3DcCsbNdh1JequrmrnsA5hNg61v35oocF
OGj9nH5fvJ6iEPiFj7YW0+XH2twOBZ/cShINC79XQPJgs+jCF4ejorJdHzEG3CDCIc3FmaHA8UEN
8uzqhiEyPEGvp6DvB1c3b91lwG1qDIu26Nx/5dMnwqaFe3iXvBbkinfHWhLe7APhDWLq4DcH4kpN
8v8IrORt2yg4I+oi2kCDHofKW+EMSc5Gju/nFVmXp0oLLWBxQ+E2iEyTCBI5ta4+jpmtUH1N8jz8
0Pj/PHUF/jNMwAIqbWgIsOOBoBb6Z9wxHpgJMuQ+/F4fZke4oxy7OUPgwLr+QCHs9Ggy9uuyaG/f
OJ2zi2dNPBggFJlJ3KJWklKMymzO9Vsq4/JLiJFWhCS3eHz60D6S9jnJBo0Nh+zw7vBOREmz7M9Q
4+e44nAi3Y8QK4odUeRnQLze8XdF+a3lOr+9rRGl6lzTKsvYW+vnfJSs5gQ7S8auBEuS8CN5IK4a
5+pPKzp5fM5kYEfQlP3xpqIKTFom2nD/6mytgJsK8ngJIY9k4LHHw8zRPTj+EJzIjGhP8DGSP4iU
aA5MB6PHbY1sGR788OI8MHfQklnQ2l/uIt3ZJ2EwSGjkR7k2OZgLfP9QL8YS3FIj8884NW7s22pL
l/Bi+hIJqXQLWvsrcbPAITX0ltVNrd9f5UJKpfU/v/Z7aO59k6BoSKiz+fnYYDPl7lkiQYoVF02T
vXFnuGCZXOYSuRj8uin52BpLBCD3HYoY0UqQHULAPIF29EiiGdBBmrDE+GYTPX/UCCKoVf5/KKUc
C08y5l6xQhcrWwDvcox+VW0OsrIMlciD28D6MFhy3yq+Shu6VFGhFaqb4yOZQ8FgqnSGHwFtNnno
Fd2S8rIMjzY9eabGQQ3H7JQOh/lWB9zqeK8+jbNPXSnYcyKayrfcFn/j8wQZmkv8qQu30VirgjHy
JVvl9CeRVK+CTvbBxlb91/CAYkOxkFas8veBvnCZOjkd4q2gcZZx8kvMb1ZlYXOv+i7/L/FsIG51
XMMNTJPslm+hTYtZvs+zoytEctZ5vfGPvQB6McYfiz1RzbxcHm9epdqsvdMnKmM1dw8AkSZkx8lH
v6jbsRMV+vi9o8QuMtR/u8RqCKguow/sSpjOOKYqsruVcDIWQNwZamL2L+zJxsfeYnHBlJ01jRhK
ig3A6eB2bv+3Gez9EIu5w8bZ+4XaKuzPPfpxCn/oI4iUNp3PMT5AAkgpZaoKHOBJHyt5qFIycjQU
NZbQ50E3ewE9XbxUfdtwxrU0ceqMvpgaBwTwvv5HNZLI8/KXZI1JjizH2OToYGQx4P6T6q6pfOm5
SQ1EZ1efoUtJigPCUM6WLB+OqtwOTFhcB6HFxxOTWBAuujVAvTq63npGZYaNOKr9Mzim7m3CblGu
Yios1tdJBM3+r7OkRNLbEGT5/8+HlOi5vxDIQvkTunDdG2BJSWdNIM6C5wH7b0VzuErIOHn6L7/w
zFCm+Lf7PANlU5RIxOB0UcT46IvNqfq/wWbxwzB2E0fROmxLo2upsSJ8aCQLczlbJ6y+xTpYUgLp
ID4Pg3LW8LTflWzvoDrQMjbvgfMIgWCIf8DwNFz4T0h4U37oDCN7yK/zA8mgI+NWvdXwM2MSu7+O
tLADJBK0WoqsQDjNOAi7+t100EGlLARAXxD5Cqkkh052Ch88XSfV9yuhjfOLGFIlxVIe6gLoN7Kf
JdMP4PcY79DZG3RgeUND7eWTDWDF6MUX9Px8nosgnszi/sV9Ho6jkitnS/ihMpSz0Ts62bgM2aay
QGApW720mQYLC1kOBs0IV3nHUHD9tG615FrAtQyqQJMQA/te0AYqLAHeFddzJMDup2PmRoR5dX7n
OVcWM0t8ecPFhShE7njuH9oDRAxG5ChKtXrGjX0TSezoL3SdYlz8S9KDZDoUeFlOKEKsbWpwUEGr
HO9FtVCZgtLe7F0x+aPtELy15ui1P50MRzS+a4pndQJRQ5pYtwYjbZ6fkgFOvzTSjjwnrR22k/VP
yu9z/g1+fF7N+j4ayNUc5fP/s3J/rCVbWr/lkBLIKjJav29JWrXmoOwp/978S8/VCV1pHKecJTNt
yFpvqhJvZWbVa+MWBB2OeMUR/EoM0/k+eJbqNRDMzbX69bou1Dltd2CVAfNKL3BkQnySaHT1X5vx
kZZIMYyJpuObG4raZqj5qAzoGt3KgTFl+PkeIpxYuzEU+idb81Aw75XO7DBFkVgPXxEcQuoJgChC
5n747zQdtZOf5uyA59+HQ6GnBmKzgKi0o5V6dHC1jpn215QCWDPMPw0dwOJ6DztPWgglCGwGySTu
DUgXKjgScjGMmrl9hbfzHXLmAHHq8r5ZX4bSmSbS1SDzDtkO0uEXm0p0QPv0RW+bT5OK3sQICLH0
N9yqtVjyv3/z77qhV2g0Od4HWVQsKsNaWwnnqn2OUCIESpc6EtRz/xGlocp0229+fs3tQRZ9ssfa
fbU4xEBxemcEEgatVSmIkluEsvdZC/7I+ONzSh2tgSz9gFXxVRLEgD2Rare/RnWQvOiOnZHiHokD
7jG8sqGalX5VFGffc/Lqs+IuzboxFDB38Jyz3u6Cii90Dj3douVd39Yg029j9pb9/D0PjN0Qwbd8
SWQ1d7zwTBBVamTjB8ztd05zjGvccFEu8KY1VGz2U+VWjqZr7JFFEDuFtUHErwOI5swjcJZTyzXl
SEJee7iXLpyasUOh6laaBhHOdcS6iKA3fpsDcMpyqayTxF6bp4wh0sVd+EUYh8rSLPAwF1GyN5EV
HDcVYAf66OtDbHldnL5YePVJ31DhyvpJrxrVY7yPTVTuQdT4gxmChx48UT8KMdoVA8GNx0XFAxTy
eKC6kDXOY1MqxKd6/m24LTw7lxFKlMxLUsaTMpIkcp4zWq1nG/c6U5MmET8jrpi2547tZJxzs7PC
TX//p6LzsovKU7WSJt9iB1uF7UgyuUctNoc+zLML5rbujX7tN24miLbrXU3krJFlVoYRHl9QSy1B
1ZVFnamI/JLF4PnRTbp8b3UgBpZ1u5cQg6eXv6a+c/JuIjpn+EcjIfp0sU/Zlrz8R2P4xNlFgmyl
U0ngkumSdhf+KIi/LutDOAc22bN2oQg3wo41U/6xsVISzV14XV3SIDlzWpRPxMhdgOr8mZxBe7ZU
vhHhQCCwQjwyDLMvUBF5a4ObgLgBrgZcXg+QIxBeDoKiSVjznaL7DRyh2Jqg0BJAF5hb+7lomUCO
u9P9qA7gPQ/7yh2L09ikBb2x2egt4ooCI2U0joVzMvT1mhNEcco5yTH1zPMQsfxxqUVXa5ATs2Yz
uhkWL5ory6Nh5som7BEAVE8r8GEvlXvFN1oGV9+vAG4y1ZJmk3E5Bn+P6VuQQjF9Gcx5dGhY0FYH
AtIOkSe7EDMqlyY5ui5tsn9mY4x16QA9KcB1QXD6wabcU6S3/AbOowkmhAvCFJsZoDMTMEaKWVYS
SnPJ98Xss1y4/4IXMGL9Tln0J0qqYkLO9pi0yg8ThOevS98EsV8L4AgYZmSJ1lkVNmwYdMAFf/DA
Gnh11WrlD3wLthJhVPpqhJriN+4EU4mUhq526EILs3018e1DX+nfWDYVWjzmd5Uum6qNuAAb33mA
ApZdTHS8XONM3Lzx1mXH3zxDNl5fKqBJnzxV3Ep/DKypij1T38d8ezjlYuCcf6ops9a2E5Wf6tRq
ixTqWZTAmK4SDonrxzDbhwDPBva3d8ML8i/ywhcYv8JmIooMT7GsZZdkoYX2CVsYQKqZL9THjUQ8
zsDhbtwH9PXEIy5nFm1zSOGrOfWw3tvD7soBN4OrM5ZmXhcrswm7OsurekZ5L1wp3ruAaX06TlGv
aWALc/Muzi/6shh/jDFwhHY8o5psbgI7qOnb4Vhh5i/8buzLKXDwKzD7C3amed1PaaQfzzc4Zmjz
cM59TCofjug8Og42N0SzYvCZj9x6kv083um7+n1oyAzZ4r8FvUaIW1gggKCUggLfxENDryStptGk
AATO491qvbVkHtvFL6NfE9FtaE4WHPlON+vMYIVpFyOXZipsVtHszlYZ+MPEDK7dgfXwCGTMrA6M
gTIgCFX+obnigeKpbnFK61LahHpYdtSNChvAUq6lgSiOgcOIBx3t44KG0y5SRKfd6ZeEt0sM1BYH
W7ACMiiDEGvDBCFiqFz9q/d7l26+vpwsav7gI8eA4hdz+C0WZnSXDYzI9wZegDTEcy4ZDnuOZuRo
kaODY3T3Ume7qQL2rjwMjfoIRwHayCc33oI/k+JuKzwQ53etpT3NGecGl9pZ5EWNUu/soSeqzIm/
SuRI/fO16AmqSxsS4pu0rW0omh4Qo91V4wV4olaXS3Yyk/GwjTHHFEL5y7ghcu19Xswv8jo9KrgD
wg0f44p/T2V75bzpTkcmYvQLTdQKNwmu5D1glN1F5/LeT+gM4Fu0vdmuMbXiDZwUilXboTT+dlp5
+KEGmB2ve+r+ohIMeYLy138fEeBSMxKHHRrP4TmEHK1jeLvEccqC3ZBx8xmO7xOsUFk5oYMz1g5y
k/LRoBY7RIPEXhm6SnlE6LRKiL4vyHmKeJfb6XJuWpg6fpeber/j08SS+TqeqbUhaltvALrge3qy
C/WOUOvYUvGpda48ixflTlcZlKAukCAanuWy+uCsfPbmP4vlHYyJ24IWJ4tTsyCBGduzyc1QjBVf
I0hxt0cRUEIwEFpYybJ4+573fKbR6ITW/VcgnzA+4ZtkCl6syRW+8hcTLXwTQ23JTXRgrBw/t/dU
h/aMb8GBlz52ETMy9HbM4TYTeZAF53qzjbkSpgnqC5R1GxX/uLZ5WDdO1Vo8qSW3tw7cbNyl3Ezy
HTkeC0AcF/E4c3DpIt9k0YIPRrooMMgKFLuLbKuT+5eLcjw2TkqBG/S2zRDr/TuB81Ag4os592d5
tvXiV1UdXBZSm6CjzJPGAuqr74ATZj9LTbpac9HWmZRVBHy5SrjYyMVJKut8sTyIgSJnNPnEkoAl
NeGrSrSTn22PYS3MoPHixRSXIeONOKEcLaKcjRYYH4MB7vgrVOy8QMJD9Dlg7XnozSy5SIKoMKk+
nzblMfiMXaGxkPu7Ul4L5trJ6lXdHSrTW2chqJsPe2YCbnEwZ7gnqW5bjIfb2QfLUxYXVBO1lTz3
GTUI2eSJuO5EarH7Hbu6tYhFC33qyS0l87v8OlWxRLIQilo3qVCr0vuTvbufDWNFJMVeWTR+kxPk
Bep2aJSjCWfb7GRNHdEHy5OeNvPYaqwmiiT8rfk45zWGBTAxQEIkNcWhdPXm8kjyG5wU+eKRGIkQ
UIv+0K5IJrZAb4QwTm+fqB9kPRHeCCWkpnePSlZhMbkjQtBOKGMoRk6rKmWAlcRhZdmYKumqFtZO
Z2D53JOIs0uH3PZfUXAR3yYDYRnIPYIocofaWlWmsaTUcDagvACNUJCPkF8Qu0HRfYT4mKoU2pqN
NQ4OUbdum4YQo2IQEi1DYBDvy5u/vjh9j6ktQGN1HRnyt7Lj0OYlCqKqB49vg7Qw7+i7xrwvlMc9
+clso0udn2uNMewiHY1QLggQcTSFxdvB659ko7jDCQkQt8WjexcgJDFPZTWOVtiCa8QpRUJkQY79
3+9FvZLbqgEhCP4USvMU9iiX2l0ll/nfdjSTeBNSOsl7TKGp224a7n7kBlSjopcBDluuAbERQ9Gh
9cg5LSHSZ36PIbgQkLGC+1/A3+Ky7s57C5f8FkP6WhBNMyDZRmG85fahbv1wwMBOpUedJRjHE2Fo
IhH6wHWWB15e+n4+f3/CDro+PXxNSQiF86SUNXu4lFZC8A2unAAbePmMBry1gm/sH0+VP9x4kxu1
+Jv62S473/iTd9sQx1KL318uExeNuvLgx3PR54WWI/27lPwdGJ1sCzHdqTP9HJTN1if50yinxTPl
y/fx/g58HA9b9GGBVQJ3ILn2mMaLORMYy80gWaYI1Ag4g+QAUy5vH2qWqDVgCEhotU//EYjiCaj1
KcU8ijdlwLNJlMBRqU/gGMZUEBEAsSYx+RVFvr2qvtNtvG1sqDcS04raNuJRs7+wZFwv3GNK/CvS
MBqVvBEJZZHIdzU6MEZ7QOgUMp2rnA9e2wJYyZXE9mGl6G9TOSqU+/hjXEbjm0kdBI1K5/HBaPOA
sw925i2pOS2EJJn4nqJI3xNpUxLdSkQy8Ao18nab1C+wDC9oU75IV0xg+A/rupxKaKBxTZ3uYXIf
HnCsNR9zdIML9ZQVDo+BhuFrHy8OWN+B9o0pFP6YOqa0aCApoC18894WylS61Wa1hiDeImHtNQwK
d8aClcjT9oDNqQHq43C9h3quaJ+fMyCrt+DhDttKmcg4b/A9MPiyyRXcqm7GjRCS0Kcqxo9yX1Be
/U7FktH9fmRFlGlxmxuIs+ywHYIbHVJTLVcjkAmLykhxXhEas6Z3NnLW+DPlLGgt6EZBTq59O6q/
rTUkgJk7+z9JG/4wh3LujvT88SCXUhFx/105teSIW025lOUiFubecIRW9lY3QczETzanpeeQPuBG
UaATy49kIuNFyM4MJUqnN5gx7InNkSyKzPLvceQgs/jR+B5Sb11TZsifTLgkNs9yZQ1LsS0vmJVB
z2IdA2Mn883pDyZXl8RUziaSe7Yg5J5ArZkj3+5LdaKNaKDcztqeb3mAVMf/zkPpjtOsnE9StAdm
hCQ1cUDgW3IAIEkR17kIuAeBs5Wzubah2zIv3Z3m5PddA7vBFdYSW9ySBJ5/yZpJ4C43nc9aADO/
JTd3o6Oxena+LM6hhGzTfoFUpf/wzFwtqJ7gLzB34dcFarYOeA9bzmQDR0tzlc3opApGsk5yFUAO
NPIsHA2D4MSDuIRtaXCH0F2XhIokQ8KrjSw2l03ucQV9lQkWHDArhCHUBgZqFhUhXCObOZxoFh2y
LhbgHUNmwEmzzb6wxtYZdw0cnib5rtbCw/7j0BSDt5yUtk79WEOQrKVDgv4BbyKTYJmikOXRWiOf
ilPPfyrR519HggK6Ey0MbEpVUAPMDB8umSqV60GpO7Jaa3MyQEyr5CKaqh2FPOU+sQ1P8rnczXZL
T2dOgdvw+scGSbEPLwRGHhLVeLJJ8of2mKrwiwIDBXmVkV/qQ2liXpJOKSOXwaE0O4ZJs7Qzx4JQ
EKxK/c7E0zkMVKyI0rkoGJN6SrlmTWuQwDacfRZlU2o1Wge7+ur69eFsf2FvY6EcDptLzTfQX8XR
tKWHPMbe/akLHpUFyz1oRay99AJvC0RETF9ZyMHP+GgP5xWnXGW3GR60EHaPShac5Cmxbo4jDecN
Hxijyt3qm36fCfucqukbLCym1wzAw8/SywNgLmjdeajVz3WbYbNBPO33vznUxcPB1sDBHagAm99/
DIFdJt5vLtHGIeYj8sJAsrAXAbxP+FIyHYvSn6KxY90/fspBlHDIkJxVPGqwKlTfCglQaqjkU170
c8p+0qd4BAduppuUhuUb30r6876/fBZ/ql1DAcdsn89hj11RLgBhpRkf//D5EXq+oDmEdPNkISfS
75UP4QV6JKmAc+cnwvrOieOtw3uElhe/7i6sjPC3QvSM0IhWpKEsrZnmfoiBe20FrVjDD4uToDFD
uGyGVXmzvwwgoBdvDwgWOAvj+oxjZZt7h0ieQBd3tsjowmUH6FlXaDyCqqdRlNsNQMsBt3SI7RnF
+hd+JYlfRsMA+1dstIjwXnW+1UFIPUfdSY59owl5Dn5Fsz64GHNi6Xe2hIxGLR7McoOVoha/tUns
mMeIx2S+wMzaktjsYZgGpr9InLFiASJtJPQ5Nx1c9pjed/Z5KHJjG8atDnRcvg36aGTe7IfmRExy
jDh6yfqeJ/QLlDlSw7595QdynkEfCDLIzDL0f91/e+DTURht1O360INOpJr46LXzyHH7Ir069vQM
xWdXG1BdssbzHjpCL/Maahv+NWNQYFY1OpoHGF9MKPkoyzNgy0f+fXJByP0D0oVeqYcFsb6CYAMW
+AKe4pFxBdFNnsnYp8MbXlL5AKbRMk6D078XF8Z2OwTe9UmcjCLZBjmkB9REnyMr3D7nKZp8FW2y
U55/3YiPBPqO4awVKkgmi2sa8AS4TrWFCgvPOeS14VLGon2Y+hGl6RrSRzBsZzP8kv1mZGdRPpiF
47UafRi0vj5GTQkXSmSVbnBWL3lHKW+jUK1qntF9cCfWiWccR1EgMS/djuIJdn4XaIIl7iwhm0Io
uiYZ6yt7gJ4JW7oNf/CTB2AXA16ToC53H3qGUwXcR3OaQAukGJUV+pU6Wha8rcyvXnrKrD5omnX6
FclhRg2f5lT/BtU9k8o/DUv/2FD0hfrNwPAGz0XCzS6qXc8NUfeH+HuecxE1IUfFUmmGVL4wUinD
dINWjdx1k3EbwLDvGz3dnXh8oTCZWG3iTrjwQn/nL5VpqV9Aa2CSt8jplX60A2rPFuOiq/Z/y+6g
CzNEeZVb947r1NE/5mTSAvgezt/Gyer8zG+OmJnm/El6FAUBYJbmLG/3DQVuXKP6V4K4ft9CMq2E
o3oy4bBafuW7rW6CGK2OTS9+6C4vY/8s+v4KobyE0M7+NfEeIPDPp9WqafFT6RzKDlLIeLxfs2wJ
nHyiYGruv6NvHVii/g6v0NiGkqDblfmkF7sg5TlSywq3FvdscINFOE6TQSWv8hzhPiztR7Z7H782
XKd9uVrKsKx/ZvCWFCjt9+M8FJghJUNI3y66gLTaTYFWuZxEzfO51qJZ8FQ2ujwrnQlQHy8jspo6
LluJjAsFKaIcqxr87TT10vJ14JsOnRxY04IGqxIUBiwNChP+YXkHcrczIfwGRbjxH4k9qVUydLcA
S2R4JTqK7EdBLNxJekXpJg8tML4J5v8BxLcswC+gKpP+r8eFD8W7yDKIFWji+n/b4k82a9KqjLWj
qSsC3uZT3CK+Cjw1Ha5O9W2tbhLTZTm/5FF8aNCeWXE9OnW8sg2CttKAr437f4JD6xXJrxJahUGH
4ttID1setsEWpxYBdAesjmT5YfdwsBqc+hSuBQ7pNULeUYAz90ipXF8aWmIRU9EtwvGLZTzIQKCV
spjxHM3OqGUq9y0LCsDY9dFYK0ADz1j3FUrSii8SESC9kM8zWEKtjcaW4HuKrwrrTmy9gd2jvtD5
v4gGsI6Glvzao9c7XJeMIVhrmYjKUZeY+hKpjA5+mDci2+f8m/ww2YwTlhCuDThI5/wN6aM1wUve
DFnteLc00p1M2BHuiBRlwXIfgwK2UeQpVbBROXTe8hQRuKrt4n0V9wFzgDvsLbPsO14ViYXcnMmX
+UR20I0sBun76r4mIFxCXMKLm3dhHGYyl3dX5ii3YV3PiE/6ttczFFfC6Giu0sB5WZHE9lfdDdGI
hOp4RXJy9j+qZKv+6aagd4KGcoAhYXYwr5y/EaNg5ZcPuKJ/ls9pu0FBBbrDUKx7puJhzKkaj9ss
jGBLOEhTpbJ06lcD2nvnNOVZgA5xc0KnyQl7prHkl+aCCgjaGUtDa/DhJp/CRVd5TUu76mG1YeAC
OGk8HwQ8OsXFibC3/7buYlSjy9tksl5ZzQPWjX3+9EW8kAaazLXyJiNqLzhNHlxuKw3AyUdjxcqV
KV7ZNFLA1N30GN83wediO+NyKxMZDXnW7NEr8piI+90vlT2sI8ougykZhqo22OSAOQK30oZjvl4S
XCi7OEvLSlpT1o/PZMPS/xHEPZ+OkVlDTxq6acm8kNWvMCH5Hr76FYfA23xZeAUkltSCdlHsYYFI
I+2BBsI4ewdAhXWlF9ckuj4ocSi3MbXV72ABo3We/SyQmL9GRajv2bluoSZ9n/J7nfIehZYauGDK
4Y0/pLsEjokJQxowzl/5LWMLtYZJDk+/kf+vQcuNPVvzN7cQFgIRbVjY53Rh3qz4MvipLDBAXmSo
MPyn8kc7jp6hBnvXSNChxFxk5PRGFC5zke+339QMfCricCVSURPaQ97W7vmPi5+pfv0aUEeEZTYC
bqp3YyKeSQSYCBCo5Xk8MIzNj5Ee8aKPY41Q4d1H5ckpDRD62mEFl0FONygXU6z11mzElsjbRacp
NDNxJB4lHLVgebh5WR/SqcmwKjWzSVnqDuVFYSXCtwg088KEY2aDZq0Hb3Xaz23jWJO+l4ol7YGm
N3DjV81OvQj1tg6kAo29kmSI21MlBNoA7cs3l/BbItIqKzbaucM4G1km09xUOFzoGfa+zqBJvqAH
5lH5g01znv9Sf1ZDt76RCU5hLqetZloe9MmSq0NzLaf0tK/3BvsFJ5Y0+b0lNtg2MKaYA+5EdVLV
GoitOpapv4FG4RxRkHobcoGBUFXThbn02pahAwjzP/2jsbddemk1yda0n4Uex5ATcER+9InLlF60
Jveawj+6zv1a29lKH2NBIZddhfFn8TSD6LDZdCTfvpDOnYAXmgC7xyy9nU13j7tMzgBl661edVfU
vLvOAsExEZZlH7rHIjIND2Vor9JNDY2thEBhIC11dDG/SxHcQ4uqU6P2kvTqC6alQ7ELZaLbf1LC
A+tB+unyCmkNqVdroAo+pc/jOvVXqaOwFNp7q1xlejBFLOLmqDNiS/gjhYMs8L83V7T869AXW4Ht
Ky2+zam7BNb/qffpMqWrjWHibOdyZAjku067wEDk9hoJYHjj2yfV72RahAf0TEndE/7WO5Dd3ltE
+YDNEdFeZGv05X+/LRnO2dQBA4dOOQ+bbqo3IgHitQbGW5Xq+fYyNvO06yTnbT6ZJk2qbr8eMPGO
63z9N1q64gce0l3CYhbTKqFjyivpq6AkLiCHoQvFlgP7hRhf+dVCk0TNWXEqNvqVagqjsJ86xe9o
Sxe3cr7zXA5jlK4ffoSalnjSp6BT1volFvq1WjN6n9m49zDsuaHEkyO8hDmNvkopmEDxDWP/AfAC
YYP5GTDSnDUdSzxBFEFEDsPYey4mRY0VKgLapIZgJMgGni8kDAwLwOFLv/Md+DHbTP2gmQBzIqh6
IOPMR6rZ2YPZG4To2M71kpwwm0nZZn2ovO0YNi5f3+SY/MIgtPy+c7SNL508XdZX48Xy6wMikrRP
ZMFZXuMNjcI/aiks03QxJEzUpj9fDcmLyac0E8iQRBuFSP+CXAosDEZGM61cPcy2G89f12vKNbck
Mde1SnZkJv5kXm8Eu/lvrv4sd56bcAvuADy7nql/10VfvY3zxw6MfTTXhVvIvIrvqSL6CVhySKRL
a97wxeYl+itknBwL28mYpNrvfl9h8EGls8eqyrBTj0LiNTt3PWF7vT5oo8AEhBFbYwr0xBct/32h
wA8VOkg8exE21XfqxFmym7Q/5G47qBw1tPhVjB3wlCaryOb7qHINbaNt9mY8naFDuQceUNZUQEtD
MXKF4NZQM2Uj0C5fHlzd6/AvBMCOrwfp3kWwdExxN8Ouw/Pr4dhyi0VLHySfHeidmcVWnTUWQTFK
o3UF3eaR0Owfx7kiF7KAUYJw4LqjDLetEQpmrrj5hLx1acvdbgNdBrpOQINkntjjpvqvDn2Fs3ZV
1fweIcLGisejn0LdvWWSMwhAp9Mk1QBqnBGovR+S6PNknhltFBWyx4A3R4w8IP1R+/7AKM8/Zvrx
BRJ2sHEp7eydd+3iBwoHg/awI8Ug/OjF7h7qkkZ7GQNjRQc6S/1ERgKmS6zugleUZQCvSbXdwUzP
ckjWSM5/6fUJzgZU+V70B7ZM4fZx31VdFQ1nIsmSaxvWR+m4SMeq9Ep69BkQ/xrp+QsLHHI6cDwk
JWlfpnjzgw+tGKdqudSTL0yog77oZBqMhzfmstsQ1xO0SoHoojQspuE0wQsMDTnbrlbGX63JsqJt
t8Cd0AeNHr+snXGw6okwZH4XNl8lcxzuh5vHyYM4dfTcd1kpoHw75ZNGlyvS4O/u0WVCRCYXVDTO
OScmswepIhGBVrQCCSxvw3N6AOmUVL2W3Uq+jXxS9MWiOUnURKLMi6gFI+7d1Q5uWXALnx25xndf
zq+hHeb+ZIgKnN6l1QP6J0p39fiDqIERn2oiu4eCQxf54VpJ8AxtfyTCtqEUTnhGQbMBu0DCg/O6
xczsRMaWP+S6pQzBYb89Cb+VB24jl3u8ZCpFY7Ud1wgylVDbFM62m1mAkepY24Vqq77xXzvHN1Fg
x7VQnfvL/eIlDqRi+cut6OGyVpDJkf7dXastiZ5PvtlgmxYi28R9deXJ0u7VpUtZTAfWJMd/AdY1
K5MCheOiRWR5qnmWfK8fQezcC4kP3zFD+hIqLQr+MPhTHI7tEO0WuSaop9LpyReWe+9gfzum+YYk
RWx3vyQjbJjr3zskxHYR3rtnPoZISkYFwoVX/cXtYLhLJ+C4twnTErjSDRLqcGOUqgd559WEbAaQ
jLz2GBnQp0lmaoHecj41HP8in5JlP13bsbH3z9aTS+86+6QanIbrGP8+OL4jum7p178ZluaxLRMl
TFz+0HEFs6FgaF5Wu83DLlIn2U/KLF+3N9E9SXRhJhjzqNzNVyn7tIUKJSYwkoHo7iugLvnPfoA9
46B45BCDuN8lkF2DrJRPxk6w5bJCdl/N55NR3wW+Xnl634VEQ/puZanWR2ldgtUWakv2LssTbI0Q
RzNf6wmXSZi6Eu6IFQ3xQi9mkhubruEVyg6C0gdrf+FyY6y6AJ0sSdO6hTxSA4ojL0ezlehbiV9q
k8MYWmvf8rD/p56utAwx2Hyhzr8C8KK6GlvurPsLs4iE96UUUHeHOSq1GNcO1iH2r46766vErVqt
6Mo2sHjm4Ci5v/clFKNtdcdXRiP8HP9RljAQ467bz79FOHmD7Aldn8Zxj++NQc1cGa7hLp8sZ4h6
H/rkLxaBDxqVOcN6SAcx9bw9tt9UJ3oK/8VVUUNvfg7HznP2VYeOr2Y+xC/c2PMGTVvoaEMwR/8Z
KnF1lJ7fav89qoWSb+82zLPGqQ/Ok8/UVb2eapfjvgTOcPzSSlKiuhq1j4x8Rp8USYgecw7PDztr
7mUDG+8bQKMJTAPusL22wIJVYYPktUpwepbB5H1N6xR1ET2Tjjm86ZRx7KDBX+9gKuU24JNPGxhK
8WZ6Pwb9KdIb6erPtu+7QDCrwKUNHPG3ZFrqCrTpw1W16qR22xDjqiXz/RbDRENFYRvrzDwhDMN2
ZX2+HSy7AQHZ8H6kWBK8YmGk0BC2w5rPsPKpKPbD7F0IwPBd/YkNAsk7UFOAWPsvWxQv6yrdDCIc
OoOmo4H7/53gTgzv49NXvEztXGA4PEgmA2LYFbr/DcOpKbrp5MQmnfVm6j9E80DzaUagdjsoHuft
LXlh8iKCtURERZsTExpKUyNtuWGx6M9jmf2/myuxRXuz7z7kJt3FunykbI7ai//RXlV2Y/QLFfvk
lk/CNeFJCtvx5Qf4FbWl9D+rivw3B3pwxi4RCj5rrrDG5LSC08S9WB0foq90Bp00k6eDhOty2imY
SpQBTtnsmPO0ZYKUTa/euogCpEj/KF9kohMR7wj83oQ6FN3yCU/rFnm2I3DiKOevJXAy6/N4AKzs
oUXW6AylOShvFuAclS+IKexBREoiWR2oP/h44rPm/zZouS8cePBEVn6PHBULDOxyT9frP9fNi6eH
sbiUsjQGEUSIBb3atiWh5m0NRRYBDBICrPsrxyWL+LKcENB8RJIe3rhnK92HVYTK7O4AyyTjumCw
sN6xcZG5Ya6cxl8NwedLGt+O2+CYFJ9/8QPbpD6eAfV4QimWsevlxq7W3kOURw/XbCc1aEFGfULJ
OvAMUi9SdnsSuR70i94J6VQpTwksBs2kkUFeFo0/BfviVDc5+rabyq9mqHqRyjuAri85mG9mXjQD
ddHN39To26NXGtpTi6sXSh9Vyfm3y2H325DLhXU4PAG/7UPPczGZGHL5n1Plt5fNyYP1tzfaEiDk
IcmdkePWeYHnnsRhOUglMx1yfqih5BVKAzg49ia8K/094Pg3kYFaLVAqKuKJqfa9TLWlxL+vhTN5
gfFXfCbMI8jfdE4OLia3LuF9X+o+JZ+pYYZ8O0PxKDllrzig1ezopCJ7twibsKRENznXyg0hrtsZ
KN5+m8T9Wvkfk1MbrIGf8J6hj4v2Al9jmkN+wdenJfmCc3zaI2cJSekHLAXyHq+kALrzmFtSTKf/
1W1+fOTQqM8JIZMx/ffMD5JJBUqz/J1HisXUfOfFI4lwDklUpJeC1sSSm2JeU1nCsRhG7vQx/kzs
TKWXh4rirE23GNe3R3zAgaMnph3fWDlfZE8ywcKofqoLkEZrjZytD0FvR5gudXS/hlyTr5g61wdk
RsCkmpsNqceJh9XjtLISTuyWgOrzaXNFMDhzs9U/rH96lVba7attKRdAU98lbUmH1OtY7SJPuHS3
pEqO7amu45qUW2OdreeWa2osOlU4Sx80A5PbZq1yrgEUupZHAxnPedHXu9WZ3FYit3wCXPrqmgZz
vpeXpFIJF5TxNFfk9t3O6K+M1IDHitwvgOAmBrXHxUqCCaQjqk2UczLZKvmkgp7g+P/q3eMwMu8k
F8z4xtMmWLEyIe7ywgMQvUu53cr3ZSCAaxGofRuJTsF4LHCV0pJlwrdLSDJEmudixGWR2W7oxnxv
yZ1S9ONlARZO48WM81WqiRsmHQpzjoUxEnULodInIuu4tvNJdWGLLJhbAO8CjUOSBkN//263JgNp
ATDnz5xIzH60tc6opvtam6rj10Q36Wjqjkd2QyurU+NP1w8P3lDb2iXVKZLd7SXvs7DVid5ITuKP
fdiO9pMXGGZUm0bywgn44NQwzAEyLN5GvudR6MvrjaZfG1NbaH47wEaDk4bpPDVKjG5em2U0lkma
ymkwTpDWcC69E1f2+5MAIkzAKO74NoCU+Ri6yPniBU8sU6tm5/9EljdHzljRVl/sXQwuR6IeocPq
yoTLvkMph6aUIRIOnKVg+nF0A+N2EalwR0Nybw+lrNB8OhenFxBav+2wISwn4+L79wFk5LWLYWtN
PtUBIPDzI1pF/mGcQFrpR0OCn1BmUUHwKqyy4/wDQKeCTma1JCVDYhpKtzOcrIG6N8EigBg9V/n5
ncBmx4F8/HjRZ7lulOSzJFjf+jrSB3Y3IfmkKx37LaaRcMhyTA1VtEVqJENcSYG+VLqJl7hW97Xx
MXQ8j0MQVQGimH5octrCp17wTNRHL3Hswuws4saz+HyaPhzALum9+Tbe7cuGeuYFMghiUaqeucee
EQkCyxCyyVcfgbAhqCukXnds0KO2HO0zp+e6MstGm0JUeYvvWRRoWUPCWwjkmCFBleRlPP0Ialhm
AVvpVuhF1j7uqEB0FdL8dFV+egrP+/Lgco6mMcgf9LnJYoKECo30vERG+jtSG3QiE3GNLvIYjLLD
4Wa/fA71M4Hh9UojQGOL7vRRdV0rUku892vm7UUI04q1zCNRXbFk2+BV1jyzKflPio6Uf7SBiT54
8BB6D0s1FndKRHvqlFF88D3r9SS4TBhFXKE92py6rOfl40OHBIjYRmuR0SO/hGE5mhclQrRM/6Sy
dp2T8Uib3ATK8vnQXm08hvL3gbwdNO+WRsl5kJVMd3b9jsrSIboWEHFvpxebARAVbzxZP/3tUUPa
gWqdinGqLQUHyDrvsw6x1eb6DM0YdLqOkH2CPnqpyxmMN6bUwQn09W+/YSY7TNqRO9XUH42s479H
7QtSf+T/mGd/024a363Zi7R3ZCG3QjFxe+x8uYhbR4zS0n9Qu6dP7pb0Rky1qHojbaaVuDGKkHER
ERplTXwoJg9ijdcHGOlE5waTAgkwNdpSH6ZSbM9ujYTnSpS3VlShCJsN36tdDWMefRTyh60dvo4i
3P1diD5iXYKP++h33aOoF0Dn4r9PGFw6YiaStBH4Rl9dR+gcirlB7guLWEG9RrMuBA0fC0YXHm+p
JyzBPZ6t9YLeZnD8kUYRmD4dBnkiRilA4wLc1c7QQFBHYvB7UqHojpTMCCwwYoRzffHHieKXBPjT
VUVnw0BjSAugCPSszPV5OvUWI5g1CCAzxTHX5G9u3cvLijq4dTp5moeEVpSx+0d3e/kK6Ib0ra+7
jZvxV9JuDTT8Dhbg3J24NzJILC/ZwLUqU7hdlfsZP+WtmiIB3zcXoJb/nimsO4dxAsN8wjQ31WKn
Wm9kbVGNTXIHj8D19BRal8fbi9O0uemHNV1TMTyFivRLLQPz4xMXWQ5vI8i6/VJEzeqFiGvqff0V
/RHZLAkfqgAFJIcW7ePe0lg18h9UVEe9sSMMeb17VBveLS9ZmYR1iYG7INcnNFVJtj+wRSVIyyPc
GrNv5r9nOUUyPAhr6Vx1H6ZQcSWQwZiP4jb71vG6FHWDBXw3nXEB+jWCRzNvDM/QX/S59TrGwoAP
z91yzuoesSzK+10ZEoKSTAngyeYRJNLcSUYHz15IKOT4YNIrEltzjF1F+PrBU7zZcMr4IUkXflER
FW2v/WHNPizmBZ86ouGzlma7ZUsiO00wRYac1GiNoc9A2IN7piGZyfIxiLCeeJBeXJlNuenavGme
h2di1+csRuss1MDoCHU2BdRJOyGDYStctRQHWDXlQxTCJyF6Ccy7aznQLMifDQR/RocOYOuEVYHP
2+RqN94MENeZzOD/DVw+bP2Ea5WlI0MPVYh2fGaiGjk/xUIAS4HMJZTQCCL+/R7M+CxXnBqX5kVj
e9q33ON0LsoLmCfuvqATTFUB3M9Z2522OIVvM499SXcT8+LU7b5Gu0iaAcWXC11o6ONRI60FEis0
dbRWbXXThDyVBADwfv/y7tXS17hkNvkI/XsjyBL6G/d8UohmR3OI4Tp3LBrOUz/iVa33IOGiqwzz
BoipFxjvTs0o78FBZc++VNNYV5Tffmv/JT1PCiS+SSjSxm0aFLdQSw5B8s8T4a4JQCj7JE8bur9h
FWW5vDc8omfMybNWpOXydFZJa7vJHvdg70dranw8OzjiP/gO9WvURHGtB17/WlUKSaRrz4OMphfn
p0UL2aRKU16fKOtyWS5hlh/chkCEY9apr7NjShFPxIjV2WmxhJG3f+l3MKsD4h17v3FyrCAp6qQX
Fj5778XKHManUYvuzqJwgBFwMKstOo/O4XQM0xcJjNHGOkSKtSDdeCxdfcfZYUFWm7BWhNkYhsCO
L9p33ep0LewfJwQknjRuPWs6UxTOKz3ySSF4QTismMlzaUw/WKrGAGEgEj8J5q60R1c99plnHR7A
tB4HrHdurQF5h9o1Vokp6iF6iJupQ1NpES3RkSBItR+ySaJGW6l+d0e4tk2AjQEvcSLcYb+2DlIL
WoIIJnymIHZmxkGE5DHrD4MLuHiAvX5+Dq7fluEILzDh9z46NGq/0Hbh0izsi0IsyqPk/++owlmu
KU6ZqjXvj6L9bmBuHPDS1R4ypd9J8rsldhY3aFvXdT1RHlXn9jkLGriY3qHNjw+K+YmxBsQpx0aw
SD7jLaBCcPXPPCQKPQXgNXDNFRxwcdvMymZy7lM2xVTstKkZuITWG9t9/vyFHd3tCu6EShuWol2U
a9TkEPQJLe3qFXAtMP9hO0xZiPyT6+o4afL4PBi7X6mbXvd2Xu2H50dJpm8U5k2ffIC5EhJj1B6r
jiSKgYfwXGd1TRy00WoZupQbQBcI2IT8czssrzmqw+gnfjk+7bb7/WhV0VEsGNRtAFfBwHaXxBST
zrZZoGIYOoQoZqIcJLKpjwtGwhM0erUtml3Jarz3QoWFCeAY82mQFkg73QHVbldf1hfqsNjNOY+7
QOkZO+F/zJt+rvQ6uda43Ri1VcHQaB4jyAQlVVXe8dSE1N5wyp4z6Fx53jiPRasb4tHSLBUdZT/q
B4oBDOB5Ziekv6xs6lVJ3JmQNP/9OWmz0XegB9QIlOk/1voj4TxB925GX1DLBlyAbxg10+xg45tr
mSWoEPwLJGB4iAuRhch0LbPq93ckawGR4AKcua+/xJdizNmzGkS8SYQgBSbQsR6JjJJA37TeQGnr
6spJaC5FLHeu6TQEs6dzXePIvW632as0g3oO07aguFG7I3f6xEpTbmEoQaJ9NDBsbymbt+vcBJ3D
wOVofeng0BYUGCnYzvwjfhSWKUlndPYFkC/x0GGK6MEMw6aYUaIbfZ2p+Da5ZTumEtVFkf/VZxiG
G2xxmh8aKqeRrytz02OxrQl2mUEu3P5fcDWWI8A3MVtaEJh3C7JS5HYTig4EDwiEZHJzSbxtC4oP
VgY9UBdrNDworAxC0GlFzaSZ5/7NJ6zuPQ4RW91KZT4T72sbX32fuKFvnCl/zp1wGKFtIStz0wq1
gylxrTWndafnMg2wX0PldzQ9xUW+ZIMl+ggSBmsBYt+EE4cSdPCQmQaQHqwjqEQMyTje1fHHDavv
sB5f1eeOhi1SJh0AD/TvQny2Bb9B/CfG1JqMDXb8/KSTSh44MPUJiY10U923ZKDu2kActxrBQXNB
5694UXvOkXkjxGWGVTL0xwAPeHb0vZhxXUhdS4/ZGxo5iBRw58ga6SURbvhF8QaMKy2T8SERokmr
S0ZeEgfv/eb7amkVI8qkclLQ7FhtOemYhNJKW+pS5Zu7DtARyOwKKRw1g9xyudcY3x2Hol/5kZSo
jHWhdohRvFYiRPcldeoVVZMvXi/0nGQelf20p8XwZPO5njAufZHym3y+5T3ZKmyNeBCPTsTihWYa
OEc8YXkriRj0/j5fw+Mo+cv1MxjEjVifOfnyXaqvA8eK+VnDc7Enn3GVjz5rlOgH8nzCJP/DjQJV
xSG6mP7ut9cXfKzZeYlM2xASLMLIkaSat2V/91x9ZuHCSm9XEDxRnVFt61kHunRs5VPgQGXS+LFp
DSECw0aPAdIUJFj+/HLdaXsBo/Urmb+mYsFbqozvVQ4hiq7GWmT7q9A6iyQIpK3DfDlG7u6LHXzz
XphizbhLup5dKyY7ByhO6WCh0ckAooD8FhQDQlYg1VkryuZkjqk6hlHDvanvh1K40KeIpohnkXqE
ZH0Y7GNuTrSkD4X0Dlbk0cRSuzSidJBCJya5fGq3uozkteUruRazAmUFLdsHKGC30b2nHWsh3cWA
cR7WbsGayRsirh+orkvJ8dH+EfiodcBLV5UuEViH3HfU457s/8mGvdY2ILNxzxfUCPxfz+FDum6R
6+gE2Tm7F288Z7Y/dqDYbnKRVmsfJAfpqzpp0KZN2kYg0chuwuOEg9RXMDp+lHCcHL+3tvd38lhe
7j7BiZdNxfklkyGpGiIuFn5BuREJarS8fM0Tlx9K+EH1X8T3CIpQNi+i8bewNtv+AB84HNDwzRgP
fLxkjkf1FRcKk4AZA8765U1uifxkp+QbvC4HOEPkwlwJ3SWsjw/rm5cEc17BS01kRCsRINn7ggK5
GhQH5vYiIn6PYu+mzHvR3hXdILBA60LgaO8B+j0IDw0bMXnUNz13AFQhdYgY1JC2zqZwuY1ph1FL
GHCuLbCYV2ydXQV/F3DcaNidY1x9Et4vBdsjO5NvzJVOxMBysVefI2L3rmzbcjPT2xGgXYt82Vht
AEyZqhJAq6+yBxqoH5853vZhgs5bPN3Xu73Bl9X112m6zE2NmQqrV5jS31q+8852s5TzXfCVChGA
NBGZm0C9d/TgT72VknxMu61flHzXhma32cAJ6s9YrtRWi5EFIKU2+w5p70GYwSz2ljlZnw7/rFDc
TfViRvtGyiojsi5IY5aB1mIcAgMRR+hn6kwzArUFz47E4Q/BBEHORnYM7kyLXEZ5Sl3g22EaoZ6M
sMcu4sxZA4xP4VZXeFlkhckNSUbt73y7dET0SIQf7EPwR/hoCnK5yVM3zizlivrFeQMjnEoNkE61
L4M65EbYrNQae5pL6pHy8GtB79MBTxcTGL/c0QzsejtTkDE/t8CVaaW0i0w8J4F/lWz0TyFEYUJk
tCgIdN4XywqvYKrgJkNB7Jt4VawsfQumKICmR6X51fwh1uC3nD5EUGz3rMBIqQrWLYj0+NJ2gM6D
HenwyfSp3oASE3kLPLFiIFF7opKAkveUhDok5fdq68zFRVHHZ2D8OvnUuFLV8aXkLzXsXvm42b5n
rgvNUdvZEx2aA5mRonxvVSOPoQMWliMOW37fKuMkNhp6N6aWEDrA6U99BAyyOHgrQ2ZFH/zB/DWf
m/c0DEztmaFeY/MqpJe180igBR8e2RAgT+9vgEEqE8UIbq+7IPjpJdaacmmLvpWNiLHqjCS6oASP
8SemLuWBcoWegaj+obf1IgtxNweiGQFmpyM0CbOIj+0tnBUIRmHHzVijIEH98vl42vdUMQaSTsxP
vGiMPLSyHknqdcF4MNX9yoC+dPqopVOJo/oT9WmQwgTHMHO8O08RQV8BcJVTedbEPrroFlWVP/ad
nDYqyvJAzFCkg/cOKLirJUarjgupWTrdvq5e183K//rV1LZYW3nInwOjfObHak9OUe2VYMJQoEcn
S3qKe+ZUXDRa5VF5+l56BFhPJdU4BHt8DxZweR4Q2xFT8pEBLkWMuvwd7/XYL/Sj0jHf32n6sIAK
pttItv2y3qkP3fAvb79msHUYG2lDFoD57TR2R/K07o9IO3/vB83IlRbyrtzh3qtzk3AQTddU1ub9
5CIGO6oZKkVBgPMqMt3ddd7KQMmD7xOjMb7DMYalWSCwqT0vwRdyPj6Zq/7qh4a1p/RwRvJPAOr+
JAlZP5f8KmjF18bgbC12rqnBuJXmBz7CDyxXib11rjMXDgDTu5+RRVbNRAYgGTCW3wmcX6Mna+8j
ocFCjq/ibNmdxEOxXd5pAW31jz3Q3/3HglonxoeVB3/pYmPtYPWIfddaNq6KfHjp1RSzpp4m5wSw
lf78e/ThzQdJWkH7vOMNT46UcSVlbaDzhD9I+xRKHoZk/TqMCpM1Po+jtzS2sNntRZyhnWivnOdH
0c5+NxNARltb+bbv5DWO2iXD7bRLWYlS8cwM49mx4NtkpabCRRZH3QKbHtiZKpycza4H7ptED0+L
AIsrAuVIjVVG5Fq0wXo0pqXf0/oZBpz7a6uGieX0HgE0S9Kzixics00qiQM+WusHV6f0hCbFITqH
kB2JYUQXgQ1DLIwalTqmdBZmEms4D+mMBwHzDWF8mEl7YllsU/4a6lvIdO7i3w4dX0PKNs9PRyz+
t/TOvSs97G9wC9X5BLnGQnGCxspkUgQ/sDYlrUhshjqSkYojunsljBzvXEqrIr5rskB9SrPZLrhq
02J20ZJWE5VWrqTdZhpEZGfeoKk4q6YLG00gz69vNrw8Jct6b/74mgBZXsx9oxb4lNVtxx9zwGDt
B5X0vxmudoDGQ/EzY3V0mMzmmK6oGu9F0LDlVTwkfqBJ9eWpoJ0s9/rWLNQURyNxPvZi621CV5mW
lZN7v8RG9HXCMwGNq5IBNcAb/CjT/qAIm1Rc7GlnjtB/61dLZYUfCrR5PWRd+51/DIbzhlV1fqad
5mtdz4rUjOJbxczaLL52P6PKz4YzOw3qAL5EWOJclt0IFREFDnU2q7hhLmojNegf9FI2dV5Kajb8
eSJ6c6AQWg9EXj3PjRpL5VruGDEOFSvY3CfJUp2Rh24ztWgYDUtx2CkCqdX6oTnYx9w4FHdjmLf4
XHyZ+pt2/ihlxzWkfUNDtEsXDjLQA0xlI+EE2X3ZJXK6lQ47CTU/QEHpw//n3GPlV3m38LBfikNf
o57Ec7GdeKDpm+Yu7yHeQFga4/ReqMdNXV7+m9x0eeLXVCkPSLYHr1qXOuLlkDRIwZ4ZaeSqeSjk
itPr+DJS8np5S6lp+gDrWnc3OGfp/HgTuEjEFCoDRyWPOZN6HyFvVyuaz9MTHYhmsAn3RZ8e4xet
LqJJC78vPrly041d6V3G3Hg3xKTeuKlMjTDFiC/yPrcGIKrMIF7s0dzupasyLYd3jeeflkfveaHT
tvb14yz4TKyishIrFsXhWmGRKD4+qrjERdWWFOmKpXL9Y8cvXwfXGfSUQyzPDelwV3UC/DnLBQ2x
LyvUe1Q9UV4ViHj5wmNTB8mkgDKyCkLEIwQAc6f/4zFyYuvIhOGVfnAxTVk0OROYn3d+NgJlgSn3
MTqwJTlgtwpvEfNlm423NS/st7zik1Vps/jDfVyaciUGMrHUG3jM6bA19NMcanJMfqam7Fxm4Tc9
O4wyGjkV+iL4m4vuvqW9KR1niLipls0ycEg8G9kUaVU2ygR2LMo7zMJxNmNHQCo4WnqBzBiw6jy4
3nS5ApwkZ4+qaxdc/UjthA/o5a6oYRCmUKxU60OmMrwOUEvR817IrEejLClnjMt56lOp5FvnC7hD
E7JEqKOOdnjgfI/Sse5KgcyWiNwUf/6+6OnoAEDQAsVKhwjSiir8OKdFTcX4KoxYgPoO5TtVlYDb
/d1Fn/57mrHlpbrjMBC6zEpeUnUxOjdpvn2Vz/19APGomtKhZrCtLrJyURN79ivW3M9NqZMqOJxk
+S7KB54exzb905mdK7o9+5jFvlVGe+uzxzsxh9XTHBtbEDY8nLCL6fnn1iW1rqWl2rLzR/79Ldzz
iqWzVWNA/wByq8sI3TSb759KAVA9WQeEFsoF9mtovBbAXfPgW5lmPzvAYSxozULUB+zdGqqq0ZhN
5wkZbIOFo/Il4ej8s2HCKyItBTMyT7mSrzZNrEiWuv0U9g9IfA+rqGA4pze+B6YhpV9S0P48fw/+
75NYqL45ycoOL/tXHY4qDEWxqFQY/dcd5GgdDebv/HygxyEFH0FNI4QNSHvKpV6NPhPQDxZ7C+ui
rawfPhAej2in+wD17ecV1xKgK2f7SlBQdhzVTs3vceW8Z9WdMEeC8vlcpF6UgOssNLdoMKlBkhAm
+k/cP9fXbknzPyCqKG4luA+LWKQDL0Avzcs+9/Ym16Z7QgbL5mAFsUHw47Sb9rZfR7uzTIvh2mxq
KHpp2sBB0n30Q1MsGgdkI3FUGqwET7ZDQIHnAHFIG5tnWJcOxtvOxebo7OeZt2u3NsUOcVg4LhNb
d+02lp5IwEECZwCl+Cq+S7RVRi5g3wz7laIVWqjNyAS//56wN7/qJOz6Bj+IsbJLfMdGWseGmcvL
l7tnrIhPxFVlJ/+orCiHdi6lOc1G/k2k14j03AzJ9rA0THJDoXBom2l9HBfOISYF19dFpDkEGyjW
7LWdhOAti6qXBciLapB8cZ+NpSgt44oskA91LvYJgY3+lpZlyTJ02nq92Q3rVv5k3MVpJWKxJwYs
RcJUHVF5fTC7TbvY++xV66YEjfnB++f0JQHKK5+LoaKQOkVESIv9LJ1w245HALfbp0bfSvN8Tb5B
5HJBiBXC6DRkriAZcblap+HYtxVTOLOAjd6kkUnje2CV8HLn/biUe8J54v4NU7wU/J/XJsg+/2fw
uoMozS8ArXbyaK/4iXoMQVdUL1DOq0zaQQj1VijCEc18qlbuLM9QzSzZprYTBZ3+YGLfRFskthS4
brK2dGnLK08oEG/u5dKI9y/bGfR/u95H4o4tWnhqLVNaMksa0fqvTWwIGFl1NVgsRi0YA5iiCUXc
SeLtUBnADOdm975aNNoro6eETPQL7k21YSUpFDpNssbjgfiX3nc6sb/9+JR+o05I3dDm3exo5RBR
mSyS6l2pNT1E76taJXCsnZpS9YlSWHdbYm0CMzLmurLydFWDY5d+oCyKvawzl7k9cr0XjRZP5DLx
GaWHQe4Li+G50EFT2TktVN07+5o09+igK4D0qn6M1FC3TjzfS8EQYRCqGujQjP/kb7lzrKIvuxC1
A9ZW0tgOHbWEJ6iT+3ag3w+UOghf0ifFQKj28MEo2kfd8DzPqkMofAL0x7ddzMCjNo3A2ZMdynwZ
OUEFpp+8No5aCJpxi88JjbcdU2IARNRbuXSuaQYUSMDdV2fB0jBlza4F0Di2egGNRhSL1YPJBnhl
VODo8pLQHGEn/0/wLZR9GXpnJkI5oII6mm+zSH5WqoZz0nxNzxuv2AoFpPCBXM1jIOJvFrjz8ABj
xw3C1IpzZdMw5QtwlVHxBJmIDqEepRcsSnqxpGaDzJheljYSTE7uZaL/c7kmTuHCVgqzCUMNJqfj
ghvMFxbx0j6bm00uKNuHUaTPVFAYx3gTGNPzE/dudDijTxrlaMu4vOEKdClVFElTcKctk8aklFxs
dYIYgvXitT2i8uIsNqYCskByJAEBpLxZoznUUZ6yhvzcBC4kkuVBWLxKYTf1xS6QGY9Q7dWsmFPp
6nIqSy2PtfMgnyFoUidQf1MR32xJQ/UoXoj6IBwU1p/7hHvWO0dDbtQhTjlJ43hX8Jj4NeMcUBIr
N7zXxa650tOdPZ+rD9msXtfhEdYoo0m0DbdJqQMgTGjG5Ng+NS3JWc6/IzbGn8i+xp7WVFU/jFpf
mBHFOJz9eerkZGI16xpLtSLpnhqwAq01ysYocLJ6jFTPRqqgSM8Yqt3BUfyjbTu7mK4crfL343sC
w2pz3+bC/WHSDkV8dIh1VQKzhCyHrHA94Nm8UWY1LWoZa6ES0tHijyWT8ip8WaUPjDKdf+tNzvtP
ULEH5CQB8TEcbmzv4f5QHzfH+wwJqUHZU7AuJsIHpeqGSbhzKaQTqyMKB4PkZSWCfVZl/2YowVYQ
3y5PizwNReaKGzD/7GBuqFSlgCOVYmB9UjWJX34Wr0gWbuU9mbz8VoL9BRn7vmFv2ENddJ0wLUGy
WDqaYsu0OCI2bSo0RYt2A0mD6gxQaaPE+QD62JXESFhcY3USCwO3ycjUB4QfspF7NXGypG0xpFRc
Txm3wM3qGrYr+k4BvOvi6yOxIpGwxJCDafGPKc4+RRQExXlH3TxnygwiZlhtTUOlURVx0XLnyBsa
rXh10so1M9uIqRLkp7WcvroLIBZVpGEHZvHILczUoqBfPkbawlJmdJYn4UOg53Byb4a7InfP4VWU
WW6iwVjloaYQTx0tnKddz3kqdGo44pG6buPAl11RX4EAQtWbZa9fVtG4SVK/C5HdFNXZuWbk8gxN
7CYJds9fPfue7+sVsbX2FH2UHcJWRLXmJ8SO6aGxVAYmAtsjUhkQPs33OylMK7xeI7osYZWE0ojY
Q0P1Sze3lWpEWH+akYfQ/WOuINYCwG+a6ElSfMuaBUoJpNKNzQ8lR73BPldYThxtqajpxz1TksBU
KNajbPa94SQ4SeX7kx/SrPfC+Ta9nx3MjWzpBtG+GFiBQS3TcMV7ify/owY5G1Ykpi6ekEquZkrB
UUfkqBG0q7/1MBKqRKh8o2Gw6ntCPoYQwzQ0aUgv1TOU7UXrVQ4E1IawWdwksNXL03luePlIgTF5
GoIAstKQ/aJM1+v6ABfegzDLxl/4EQbQPGoWdS90i9UHMV2b+2uJXX/1MUVWr+Rs69y44KJqy427
32lcx9YXKyb5Ff9jKqgiVzKhaf23Qj5gCBmca5rVY/zDKbsvPjJYLy4OYSYGViHJpvLDjgVwfXTI
KJK/OHPFhcmR0kcKtItmaNd8mXRZcjsTy/d+uG4AmfJZtLKjMFyvldphXhkUx62p8ZhR51r0H/yl
T6BsQl1wP/gyu8JukfPEZ3fXKunkw2fo45NFRH4rNl3BUxP5EQ3xlrcBYd2z5sFYm7gFTD74eydE
sebxoARfFdJku6CenjTr8BuXd4t19IIHeGBRtMiAq2nNqpdNRKFAsD0DABTCalEjlZiaiZRBkGxy
NQLpZS5VrIBZsPFLS0DRBJU+6AEpN7mjS5/lBPiCsGoGrqc8rc21WXLbdJ+lLNMGKULmpAGYxEiA
wNgmaF4Bji3Xo0XoX1Sm5YFYgFFVI/CWbnatd8r+fdPyad7u6FNC1vztDHRbJ13z8ru85oZ/AAPw
XDeHeR2dfXMAA+PBAgcrw31FtV2H4P9AFdYXt5lqKcDFNoweV104D5PAh95PpdXZUlXKOtw6ghSO
Z+rS3WFyEIbsNM06gqz9edtjmgpOe0u4uMPweXY9pp85qMMly0Y5RBiNibohgue1nA4ugfl1hvcy
RRuU9hNKHMO/e0rJono3zAVVEbfJPWxXLOcSFrq04POb/pHt2noWZk8uUF3O+VD8fCFnJE5JRpGS
WaeFnX/sne6X3StIw5RWZ/dhpfsq3rHGjAKjXAJoa9XjGrsOC8apW0tQJ343a8mjKwEqusebO5LK
Kgzca0QeMdxZOkLYa4YOK1IU3irshqrnButGW8pupYG7EQOGZNhPsCx/EMzIHoCc/lAz/a0e1Vt5
cDeZ347WWenw2WNKzRUV0vJdMnOvFLLgW7NBlrLl5mSO8UYEKTfcFvWdKQoQ6B0C4qBcpi66Lm8u
znpy6KVQihqPlwMQxDzQViMjNqB7n6ECw21sT7co/Z7t/k5fcoSBl92mO1ijvO3j4gp7MUB3snoJ
4UZNYzHpev1wv1J21H0X/8V+jLhrXCegEgJTY8i++/jWW6a3W+IaV3wdvA0mvm20jsO8tS51o/Ql
1ioE1skrVIBQPq70aoXsnuTGI3dQcRBSJcLVQtRmGGwjMzLoUbjwYZ5sXkr+CODAyrSP52B5ZbmH
XqIleJobXczSoDn3zaQmWWikF71ZJUkDd97eLtA0byFk7X+407QBsUwzX5CrO6yC7gr2NYSUXHTQ
p2gM8g==
`protect end_protected

