

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DYkUg37UnVRJ+X5v5iFDmCWObMw/mUCrJuxa/Cr9wGl4FgcJi6OQesLI1M+aH7+emQJssoNWrh+N
iL9trwbpEg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Vb74X6mc2H0e6MLiEAhBKZ84QSTgHhg3aAfwLeb5H8AGScZ7UqNDKDmI5IhuJ/LPpdHQCtOent5+
I1p5tELHTH0LzN6BILTKGZBdaGJ2AKKoofyljqaR51srCF/ZJLUOrn1XUZMkdlutYXGikghh+zK5
6+/HFEYyz6zhpfFGpAE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DUY8u9eRLqeXCDG4E2/8OtDIacK06AysbSio1XfMMKnofNQFNkb8eAjngrn4u/YZ6G16ZNMG7YoY
jk2Rx2Q3M5GrNkHLNcW1r1FM93KBIPYna3s3UsOdPXI8u/gdrTwtTwv/xpFT5pO5KUummozg1ol2
CfVK4phP0ptL6RF00qSF6IA3NotRdVSf39i8Abyti2fNqAeVQtQbe8y1/1WV9RrHHqEjarv5sqIY
6GslwJ8wdJjPL0QS11gBEh6rDpndqUhWIIFTUrFMd1tEU2WzUCNSxtbBPYlWfpU8e4/l9e5xSsF6
weW3wzZvwjgR473vdWcupdpbpXFjQjfOA39+/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p0GGQgjzPW+6PIUsMdZXTQnjW6BUopNyvt7ApHmGMwjrt0lKkYFdeq6NnHPNeKi9xrrloGAO2Tha
FhPoK1WSUQvFoRR4uKVUk0OywXYhciTgYL90XL5T7z6pvP+T2xdoDnAiUPoqzH/Ubhhi84EoGyo2
+zIDCCcTvvnznOBjfpk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m1/kaqW4ETEcDTOeEJMS5yQHRelnhe+7sXgpcKiP6lTf8NZHj87LtgfMx1Oh7TGMtL3OsgLwXKl5
B/MVSSTPV7z0P/OvFd/MWYJqIMAVI0yV4hJ8dwWC7KK/kawdL1h0Q4iS0dxjn9/392LJCmqkJJmj
TEThXH1uoH4tMKV7xRRg0/MNNOk8hPErcV0Sx7ZxMFsvJk/PuOEi0wzy6daa+A+gop4M475HPjAb
iPZ63o2focv37v9R+NETZc+LyDzZAZPFDxIiHCnZlRMpU+rYc4lLu+Wj7afASerzvuIcVvlJO0R8
MuDtSunchT2Nxfc8io8WUTVsWpkmP/zQb3BvSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18992)
`protect data_block
P6V53PQil1RAhvKekQyksISmZzluqzIBfr2EGYz3fn6/YjV24A5LlEUGX4OmN9styR1NDR11VlxO
gTjEIyBkSCa1YT65wcc17w9zfH3YcWeTfRYFRSk3JE372sxjJSX23Ar2Q5zYA3qHsV+u8iW499es
Cqip1NbBRRhWkjBOG+YIbo6BQnY/4IAqHXoWulkQf+RvhUQY9rl7EQOmnfYcsbhbCmbxFvemBbTr
LpJdG3K7iHfL3W1zEk4gWuhuyZ5OlP51V+CBTzm4ReRGCiPwQPXgAEhEEcDwQhW8pzwukQLmxnxF
Y5nZ7ilX8ngslYsxTPvTENAy81V5NQmecfPg3R6K1byZam4hgGsQ3WpTZyq8w0KKD+qR0DNLmuSS
DtyIatJtUL9iznWHqYhlDfK3mJSE21BGwrwHb4+FQvJNw0pSoCCCYbgnd8+w+dVkk1g8kZ58KodZ
q8RbUNib1wuvjNPnTkcXahfEFM5zd0XL7Lxz7fxAAmdz1DuoKPk7dxaD2RlFGkByv8AcYfzW9WZQ
Min0ABqWAlbjgVvRoI555ttsr8g49nTLiKxSY4lmWVIgQyXW27QX4SeBI6EXz2QIGr8bluDKC2Wo
xKG//VviKOmBgUQYnxKK5gbLppREe+INiIDpNYUv0NDsqBz42FoNqH50Pbvd4rlYttis8NW7A6GP
D9FXa45OOy2Fr1QYZw9RWheY3WtElfQvCKZk559lcnmM1swTj8EnDALy3Qx9DrpNhHVn5S8NMe71
rknWrGgGPl4dy7LCErcwvtZG/73cTATjaFdlgkyc+O0OrVDWBXhAK90/Cse8Lb/yr4lDTxaqNSEW
rVlc/7GEO0pZ7Hx3iNXq+O2LmGhw8c/1Yz/E2g4i3cRPX8kdD2DnaUg8C5K41qPUc9W86PWn1zYq
Ilk/y2QmCtG6VbP3dSwV6IglFr1dUwCjVp1RdJOe+RrIEt2hSN988EHn6ULvc2LqIl3Chmxw/+Y9
7Uw8Uc+utHe5Bxo/PNMXazpU3gHuWYYxaAxY2KgyOzsBrrdeuElSh58ilFX+mt51Dw02UEW/OGoS
P1xHt3ZQAuOPLABFSm7vC9hdqfNpcd93o27MW6cjVwyMFbInSS0f7x8iUxrzmdTpCv++HDMl8o4d
Ck2R39ykxs5+SwQWvQA3Q2aaFngkJ3wpCQWwJ/oo07Kw5Y9GbuxGoYKW0ClU5YsTFZUcQ8o/72Iq
ema6j45sFrNYdnefTo/3AlV9ii6JmzEfSjW1GoomcRq2nNe4GHPRAvS6o+4iVbVa3aufRkKwoa/q
oTpZrHbeGCre5QytlGbthTM+WesmYEZxCs4qAeEn/UXU7lr2cFKtQFgdQLo7RnMkgcelNuPt14OF
SGjFBHeLpnIdePlj98NV0R8sqGYMu7/zVIXv/cNJ0jhy+nt8BD5UDkd+9T2eOv9D4ekMvz4nbsNV
jARHit6gJsTeMNEQGc5dRlBzrSCr4bUEXKB+YrYLxgugrtjXuQzm0xgpbAZN/rTQCNwVWedhVSaM
ZrICTJF14eveAUtyPVX4gVCea+HJK8hDDgqnwa//MF226JO1y/+Ii3D/M744kZ+7NQvNWKUoWZqB
kLrYF4vLwa3vOaF5vVFSINDh1VdgTZC+GSbQzbTg/X6jfsaBci65MVCkWqqM7dXqUyAZKU+eCOdH
Xd6YNHbszCxYcVK1yDfFaYZ0rkDyLp4CWNxnH8BFSD2l3lzNfwxK6exsvHepTmJuGVeifw1QPII6
YONRsIl6sOEIGQuB2FCGltcOUzRTevXKusaswxJ+gjhc6e0BeGBrrcSKWNbe7xzZjJqHdOhZgrG7
5iw/PbBob/97Mht6WPmp6mEYwSC+mRP+Q4B/KCC48EvL/s3nTlUYZ/NxBSq0CJTUXeVWiWi6MxAa
sQq5n8bQlkZJN3gntNUmgCPnSbrnhpea+/Xx+VUu3gEIUIxd7mAl201lVx9DD7A5ZyDxI0WJun+c
D5K4PaBHuRl4JcZXVfK2PHFv2jTmmqnB+0KwR5wSbFOpkD6qrpW8I/evRGmIMAnzsrq3TF9/R8x8
X6TYzc6nAMJ44w96YnhpW/H9WJKddbULd12xrXo2TT0Rb51inXDHYUB28ns27w4DvB/xKYkWbIVM
OAkHXXENR6pSZEQg/POJuEEcky2VN1Q34okUhtIqZa9/h8/kOulYspx4OyQrLE6LKI0FJOcAqe+U
O8jiDD4c69u+u2KmmD5vghDzHiPuT1gVhY3RPtOIHEn43aGpU+qD4UDGN3YSwlolfTQ6zlsd8n7e
MzVSy0wYMCE1zJFj6jjTQfiLc+VFm5Jzhyz2iqP1Id62MoKI/Umvzi7LZTHuchF9lvHUu9VgiVlL
s3pF9wklP/n+gg4k1khzeRrRD3j1kHq0B8Dosv/iNwAasjbgjltAk14QClDivM49EYWnc7sk1IVT
+05+GASBydTvxx0F24TWgotuJNKGv1Ow01PV7kn6mRTU6czyxi1Xyy4p6GQqo5gWgHW1C429SSSA
B7d9SVWJJ/pSAne+BwTcA5L92jKCAqYzAA1YL792+jIMzXpUHCzsSZ0d8M2FUrwSXqoyvWou+eqH
GmXXsNnB02tTPdWCeOT6WhlIa2G+MipJv9MlJBk3gT53yojSsjucffKxl7jAOL92u34nQB/EfqFP
dVdmdH+snVnM+DdGKwBPdzeMdAGK+ZG0liUlJJybrSEu+F3xl+0WItGiYov1rRFOPhag2CiO5U0O
ycApRz40clsHbbJmiTEO4V07nDYu29NyZ3nL/u7mUBZ7LXRkHyZbYlwPOUbHS/bkeZTLN26Su6My
iyWzAZGMCVpOdzRGuPS+9W0IWcosU+5M5CfaWRNqyEuo3G0MCQ7JiXnKBd52Sm/FuWbZU5cYpLM6
nzsE3DinkrLsWTfzHH2QT0Y/Uz3VpVcQ8gLLDDtYHV4DseJljIBHRvYt+0d2B/Jt+2iGl6UoXjR+
SMsuVjSbBmn9qQn0PHCk19eeXqws2gU1uNHgRS4cYp37EH9c2anPrB8kfKfc0WqQfU+eUcWCNvtO
zqC4I1jXysnPqRGuxAhSL88a3TaMadtUM4Evj2RUTyXfPLk5vDwZOJ8pYXRPBWb+XspezXm5K6a0
KXv5h6DuGLBl5y9N+/OlnOx1aqy/ldhSi/8W/lMtPqmrK0uZFr1Lnvtdo4y74lA6FJ772Ba/z7i5
0ifwMM2blQJ4zuijJ9jlZH418eH19XJWGnSeIKF12xRIXBxCr7GYMyYleNkCnY8PY/fte3OlNFO3
4X7iXhC4TguJLO4mTi12j99BEjxDcQmSSsO7pK38k8Q6ASfgDtS32ieKKhpJxaBEyTFbvmqV2JM6
V7W2K+H8Cd8tfwZvlkoe0R8WyVUAqhWYYoLVLck5i0M7hgmOqHRyg2GgxgtQRNFMTpsuD9Wp5lUE
HtWLNjFqh1wd7//a+b+unW1QN4zQe7xcPZCfSyiBGIK1mr2y5ZFgtssmXqFg19fzuBnq/lot1TuF
rXYRZDxfl81RekcJklYrqO7tJEj2zWLBcOzlpap8JOt9tY23qcy8itCI9pg6uF9E0cPtUeUW7Vx5
DutU/75QPZ+A4Rv4SOrp7+Fc9SDqCwzz8Msg9YOcKNOljQLWzAKa6yU9N06LR/mQuZ7J4haEZ6Z9
zOkbVl1AbnVOdLC5Wp5QQqKCkoytCaCdWDZUYbPsMWKjV5DgOPWSDWxl39KZhfXnL7HO+c0awAST
KoTfGeVFvDZQugP+7oiB2S1GttokqG+3nZTr+VGkF0vFwAsQCHKMzkBHlawIkSHIKqvVGFgLetQq
LzDklWrwlKkbp/JIegIeVOrZzMoc14CIsEaxYtzA4l2qozZIL888vshg008/dK3dZCgRgtkimAzv
y19HeSC11W+/C+NU8M4v2Zz3jaPiYSEDGNFfezGO/r49j2IOTmnrvdQoJwXLEyVX90hqDenawoMw
A7Tx2i347UQ92cAWJ6UluLbQ43hxyuLAv9nfx1I4f3R2SmH1jmdddru2TvCsH8fSHJkodaHgOeDQ
jpePGNxTlgmRgBjYehoP5nxgKJ9fxXVPEp9sRwt1+r+9qn2l9LnF3JmJSwyAE46vwT1L88IMvNnH
xMl0iSQl9wWqdRVrFCtHDJIx/UqV+5/GLIYOhCEkjTD8iyP15nXFqOQeGwsx5CuZ0K18WPRTHPPo
EjAnW7eRwD+OGtije4RBt58dzgmQmcGWW2+d9+JUQGJwSiNIO//FliwVzyWTDNrPQW7/81n3ToxV
dJE24gXgmFYzjv0fEWx3OuVCsfNjpmgzYD2aJwxhlsTSpH+iNggoq4jxB1J5snPUmNtt3YsPhG07
X1uV1ePN1EYcqaEvv6WWBjHnZaFOXWkNKKyP5fLJXU3BHFE46vS7LfEUqQn2YAaZQiPYdRsZE2BW
XA03UFu73I3/gSa6TTq3cHg1I/uDbfEQLZpz8oGVj3U7RKzy57TIyoiKNrOA9K0E1UX3d1SyHcUK
vPWfMKRQTwGpzmVbcVLdunZKoUtpB/R4w2p/5fKZlSqbDWBiY6pwu/HL+hCzHktBm5NVhMZFANpp
FwgkooGSD58sdA7SJqTkpofR4FOzb+zwaVzRcfI6/MKOaH8XwykIm7Y3n0NifVdA65w9l1TF74Gr
OoK85yvmLWfBBMula8hS6qfPaerMVA69M/LnOkPRqQLhpyrqxjcCneESlrFvPo+Ci/uIz5tH5D7a
ufxyU9VzESTHDl1wtaCRJl/EwMDD7w9nzdF/E15xQoebT7EkagyUIDNdJMeY71UDppwuaT02HT7N
H42cy+dRr3sI+gOHEAC2nG0d5QC0d/kImvPPvkkuJYq9qLi1E1pF65FGRgxm4eOs3TX3ouuSD9m6
XgRVfwk/S/XEL5hTwyhi9/NMyRVnl+riZHupUIqrm8Orc9VWhyt3iTuFYKpfUYclhKc1SSMPDt15
JvgXVuCqFWifHJOabEWSEm+XhpOLv43WpiKblCA0T5RCne2ZXf0uGf2WotK+aPBfznxt8j40PqEW
Uu5mv/4qn7oegKMOmw+kvLcwyq4jkZHz6k777DQxOds+KSLFBb0oM+rUNwARDL5+iW8s+mgjrqyy
2r1mbowcdw71WL+pW39F7jzZfevyHhm7irNtlFvqMB4DNycZZU31taSsVnoUhQUX3e2lVO33jJSC
igVPo9bL9j/Zdp0qJtd4y+cEaRVwzVk5T6vBl1Kj3sZh6kntK9t01pSd1/D8HaOy3lFYrypDgDNn
W7hRJzHUoxdqaSUiH7vh+JgzruKZ5jXRLdPdtZLCYP2NPBLBuhaUBiTpAuUKRTlkK+hDpPgGQq7a
m0qDo3i5x4WRuFzRkyw6PARUejWSiDMYPxtKbglEkvH7EN0mV+sg/vlvRyqvEsYmgkpyrZ09fnux
1EqlxVGJltgjlzFdAIQXlARgijH7WF36EOsHG44hpk3KSn6YlH8rAhS++xgdes3KjT6V7AXHtknd
lnVBQZJTsbqTAUYcY0wLwf3HLHHgFLVFqjRAKTRKr7a4c3Et4z6u8sgcqWtd868jnpAQy1+IiH6z
ANHT7ywxqyk8+wOPAmdMLYL5FsVOfs8ns90Q0uvsWBEZbwE38KR0ju88t6Nn0vkaZFLTVWAuoM1r
K5M5w7kcOMzgPrS1hxviKiNZJ8YT0B/wwTchYbPu7Z4/89nihuUreqKrCsU8m6o4OV2RvvZCwRUs
oBsgtMldaWKJkoPulxkZC86zMh2vGrNJ5IuYvV85gtHMlNYPk1FX5mbPPt1XN/gj4RUM3XLlQqg/
x9JI+/laQMcTKz67XyuiHas9l/u2vBcHIAxWyio1ziD441CkB039rxtwzh0i5o6nnsiomIW/rePg
tcFNXE7y0C+Twl3fx9c+2zEfGJDDz6IbgZHDBztQ//+kOQydN1Q15gQpnFyDHYEhX1PkiN5ihbrh
FlerfBl6Lhv3NtqOIrT2U90OBazmh/l88dvAC+X7zTbeXtKCPjksl3+QoyQhkDjH1hH1Rtw4M4oV
RRgFX2aol0qmHOBcVfNb21Pu2LZ51DFQl47aHKQhVJRHxf8VY3pckyIDpsgwK9sCaFXusXsY0QuC
mbSp3fR8QDMNkY0nxNfEX43et++q8cTIPMEqwVdUeBdvFop17xBtY1Glx2arf5WdfzHA2Sg7UAMI
lJNW+xXTYwFg6HWuC+K6yyqGpeDo5eduakDuPfRylKV0108faBnztlwQejHHUHny/7AdCi4ZSkxe
gk9F0J9KBSj1qS5u521ubamzIdjb5mN5xJ0ASZoH5q2huUyet4lHAYCHL+54iDsvdDcXA7Bcy9BI
as7dmGZPWa5pJkS128I6YQjniZlMZ9+xKjezrtXkQ7otyitYA0IahBfiLHDWp7o6qp+FGMkkPw4o
nj4IOqxsS+/2Dr3YQStfEX2SrS62v6jeVrElx3nvLd7f8cUluF2C05tXw+LK79+OGXEXd/h4C+gn
w3QWBALDYExe9MY3FfMjN+iIB1j6AFiZC2CCGStbMioRJYoHL7/Vzyyi2TX9qe6Aedsz2gNELDW2
+hVlH1roTCoxubqkmCyFOKPQp8j+qW9yXWaekZW9uLPrObs6kZ+C0zW/GVODqpXCyaeDJpiHYIly
DOdBRQD0haKz/9WfulLzM3s1HzniX80jwNwEnHLs0c89llx42iETOjAczChBPu/hNHNb1W6GFZj8
d+Kbc/5VdpHS+8bgapvDWHmmgPUWlfT1A6uaV+QB4FIdaUylUW4nU8OnXFCY4oJZqn0Uq0FmYhp0
U0kseqt7T1HOxGr/tftAsB+/KHoSbhRB2qLhYh+SO0NCIfAUifYAq9RyLLWAHSHfW/pJ2UFu7CF3
NO4y7D+Ydm1Iuz2Un0y9aoXda8gQMOubdG0h5gNarTkLJo1zP0SMOk5EqeqYbJ9CNtqWcjfptgL7
GiNzWysJlswVrdaiECUgB7Nbz+LrHRjcXUmz/5rBy8bZpPKkp6DjAgLur/giOpWGTgCaHk9plRl8
70oWZwfxbf/59WT+BK3AjvLFt2hnLNOFV3h6bNNyFbk5Ds5wjvWfsPelgRlem0uLnQQQoA+z345N
Q4GhDFtMDKhESdL0hVuwjTzDe2poFwLSI1Vl7L6+00oJaDuH4izyxdRgHG3RdaD39ofFAm9ksu/e
cxHKdE3r1S4Jgq+WS/JkqX7NXWepjkShBh1OCuBDd+NEe3njmkVQnnHssxRfPcHDNNfe+bEOxh1u
onZp5h/a3sbiJO2zv+kzL4XFhAy6+7Fl9EvLSB39tmeqN90dQBgyGedCs0sFzscbSp9YLR6ZDuoi
Pet8Y+roLuGRa2JOqMzevsDTaJXiHeAxQwc3YNzXj/iWDgSiTKLsiCr3EsEcs9MdBWOEhZWaj0IS
kXk33cQ0/psfgjcbeaQ0TOhW0BCjPKky4DFcuBzsDbWTt2vaBwML4cGcg/2cH33KhybyqPAf32eA
ux2JiWQOYrsKxT8goNIn3GXlNFtVlWECvf4HB5WVwF58xhiAWb05kUFoID6LOXP1jz7TB6u4+neQ
CK4tBakr+pl9H/YnmtQIlGo/13GPeFeZCWEuXIevOO+vjwXEJWrRwIwvJitfZJuw2c0uMpiRGKhk
5wEI2mL/J1XFvERYlDUpiV/hVN58UssFwpqq+yNmxjznv548+zPfaJ/aXIxkAyBudsxslsqyFk02
i9kER+H8wJZLxuNwjJmWNUyeZ9ckRnI/Yt8Eyj+iuVFR9CZ8HEVrbF4vCyoh4VxNp0sWUAgdG7UU
slzFZTTZGM3ATh/4XjPIeh3C7lhiyfO9Mk9e5WFiinP7c13TiVdxkj+bU3pNPnPKlNemZvTPVhDY
YUmg3TIwM/AP3B1N29HPyH2Ad/f60pI1Ap+7yWYJ9gF5vt9tol3ZwIh8sshqLYZD3GirbbsaQRmM
K5RGjf7AmrtcEOGKAsCVDMf3U/IE4C2iA0nqgHLnFjJi0ZVMCwa1dHE7m47FS8TCLPaH/DJyE1HF
aduiEFt+VYaWCTuea9NtyB3glFe62MSCTG2RjsszMmcB+FrXSNLk03iKLjR6zvp5XVGlvV5RXp5Z
gtodIkwkoNyFJGb6MbIe/dD2xepgYfGgH0asFkxAIL7qAaWPh7CebEuVjKnj1N/RUlFZOX/Ae5Dt
Pk5vMhMI6bUj9MpL5EuH79VSYWCmfaKLcR/PH1xpzoTLYW58rocKeWRZ1UFrbd7LR5lemjxnDccS
K6LrTOcn3bR9lKqPxG5hhhH4/eyIAUEQh2GE+gb8UZVVlMlUyuHq6ve0587xiQXwf4QIKvqdYuhc
TxbZ9KaewNp5dyAywk7y+M1AK+1ojWUDoCecqYH5vx7619Mor8aHzakzFC73ltqxQCGS2GFuDdOl
u9m83GPAqkKm6WgMjK3qHb8WQUH6+XyBEA1qLVfiqYJHKlGucnYF1lQbD+nygPh5SpX7B+f1hmJS
3sNe6mJD4ht+RNQ2J5K39KhfT6kmFiC87PPJS0e6lP4k4ZjV3OI3d1zRbsW+jqd0kRskeGGhsgbk
En5hCSLrYLlrD1KWPy20f+9Fhhb5zeiTAMuazZlVKUEgiH2ShLtx69DrS1Cw+/RqswX+5OGOVyKS
HMfBt37FmLLnBBa3E1r0hLQrkPcW6KBdhNzOHGZ4OVq/ZgTv60JvkvO3Z9AOBLmpbMbCrPIaoRq2
Mromv8bUlzActD9Xbum2Eo+HkdKybZM8T+2kihOBWBOQ3TgoYuON2FwYpBGsRKJqPLcE7nL3ILK0
33lWRyFkzSIbX/wXmFJISbe5OUQX12sZKA7q4bCliZjEYOUq0KJVYFCUbGcQoQM/PgP+eOSmC2Eg
Dju6Wf0YSmyUJirqPFiUY81beLE/IjB5XHRpmCayQINDRX3Jmh9vWF4FIkaAiSz8NOhnDzd9iOBe
hzV5sbKksKSkrfqSwbVZimq+l2aUx+wIGDVN98o1R3Xd4iTnZ00wU+64Lkji1I5Z1W5rW57VpCIW
Fozq2qrgzUXSgcTs3mCK+ixI06IrtiF+MAiCiN27l6omIYdVlm9tTJUAW/P++LaxC3sKURHExjH/
Qr1fiIUvnCUyOoLM1Pch7sdWHsxJg6VKEEZoX5l+XDiXliPMAymHl2hn4aGdXe0DuwIPxN6erOfZ
XJmxFn3TRG4M/nRwobhw/jJq5zyxbvmNO03eNIFO8XK+vBE0OtgrSMqAVoWCLNIAAR6W3Txoa+LJ
lTNnJJtPVyAu2iokHxtX+baIGsMns/JKjQrxJyya0RIeYGUQOqby0+iMrGcSCe/vnrSR0dZLAIDl
n3SSUUF5WNVKbUfO7PrgKls3as5jtGRmw/TLBMC8JMVrAqLyis07BdgtLgHGUyeFk2asPJj7RYtj
jKIvkDZjxBC6HXqsMevO0YhE2yUuAE0UUplQBaJa90hlUaPAUduVio7fo50NjiCxBUN7qPs/drIh
KA+9zsLCSQOz2Wgie8/AUP749ChQJ8H8zNKRKr5liLzHMSs5I03zjISq7AwbYrxajfNEg7d6DwpC
qBKMaYE1T+zGAfH7gMXw/lFrkWc6ctpuPXjK6RysTlr8tHILPLv9k7a158+7mBDI++kXMMe2X3wV
YPYhAfktuI51nlcUpW7FRvd3GwOZWCfrEPhLPTgVNkRKJjiW/5Ncehtr1WyxlwzUXpEqIc0o5DDO
MS1BcEvzrsVlqBoZmKFH4qShprWD0+18RmJMDfGqYmzVg5a5362uGla6RCYoIMIBwKaHRk/96UhM
GVnbueMQK9dpNTJFn0snq7A38HzgUVSQWWQEdEfuuAFUX+Uw2Fr5+xLqYtom16S/RaQb8h5SSbWi
VKyd29Z2khF/d0VpGjAF+YR7CTr0/9tdNmcKG5xAM21nAVb9bgYkN+rjF2qXtnJwWS9LP5wumWkE
dCqXyFeqx20sXtFGMjHCiJUL2hUQRLbXnl0wNaf92XJFOwhNCu1hkTkGVFu54dWTRIEvV++xRABm
P463CCvBc2s/rmps9lMGmBuNaE9s54RAMi61UwYl5FtfByMdm+BoRse9xQDg34EKiW9+yTJ2/1NO
l4e3ymAWbmULQAght5WoIcqIJ3o2iqFjs50CZFm+9/hMyPftj9fGctvhyF0+CF8tUUH9QIqWfYVZ
beoWmmcztOriY3qzNWniLGB9gqZAUE7GP8FuRvM1YzfFhdAK3XROqjlxf9U4vYTJ/tF2k9wGibed
KraP44SJWmFFYDkQDjJHzfhhd/SscQULlj9wu4KVSB2M9NhEJferxQw76ieMTQUF8m7DqbH6QEYQ
309tsXxPUfPmNMRfRbt48adea/KV3GYI/6DO9mHOSYip1NdlpX3y8v03i7b6Sa7LpR1gu4ybviOt
SftDjhuZqXnSM7DoHThC6+57F2QvUetO/xfyKbQNmHizQoQZlJL397dPRjfjlKxDTRMo/EQEHQ52
krWDWUNiaSLzRpU6OHYl40kJ4kWewR0krHqmJ2MXVd0i4idqDxgpDKwNrX4Hexe6ReXvRD2hNzEJ
5P6XeJLI5T9xOfbpG7DIwC+Gc/D1pvcyi+4sGN5C6KmXaBskEPIUyIAahXxVMY25BfeeFWRIE45V
rs/4dvUJLP1slUmqF/foqKXp8zPItn6x9aSmFe98268CilvVLZNiTFoCGVcDPhqyDj8jPKhmT9gB
HceItl5j3ao6HeycYbuan6FBwc+K1rTZhEW/p/6spaRl0AuHtzexW1HYj/q8N2zIEoW6rx6tNCiO
H5ZNfND3ZHNciSJpWkCbwHaTU9bh37KZEscEXH09Va8IMCGWvD75UxOjcxbi97THC83QZ0qoE+wI
f43769RlLNn9K7gGdxd1hBXq67ke8HT4hdM5Nl3PoqSa9u+yg53l9FTqV1rELhsOKYHfA+LYpK1F
MFb5Z7JNN1kTUgEMF5UeA3oj4HbupS4FZYnfyGH0S05aXcvrh4fUt190aqVY/3ZRlvGE9ktZ09+d
MiMrvobL6fVPNsTN4EI2HYepMfKRsbpYfhcEnyXKNeY7jVYgr/WYxeB9Xq6d8kJVdYrkcdB/kG58
y6H6xio56znqfIc3PTmUk2vG59DU/ZGcccP4bI6a/X+NliBsBml7nHUMvuoLIJliuZoeCxwikDrw
r3pD+qAl6r8FlhI/XciPuJ2yGchKl3DI/2tOkFSKwEwRHCPVtJMFXhIfArxwyuYihZK9wbZo79QZ
Nx7GX4mYqG6ap1Wq9N9XDWOzpN4GfPXznJ8jtmp5zp4q+X2weg4jieHrNbGc+F9R0EH+oaoXSXdm
jiPulVD96yVgUlx/o0265f/WWJ3RmxdQxGv2m4aBt81pX587yhk6asP3dYD5Xuj/2J5ORIAeHDDa
fhtuCmAfwS29Y2XW2Fbt+tOFojgXHKdBUAXnxbIH36wlkGceuoFrkskXi757b3xeg2Z5igKUDlq9
Wnnt/A/Sq1q9hBrd6+dDs7s2HeSUuIlx2LZjkzxL7/6zv5p3Bty8n8be9EaPi1/y5pABdoWzHqBw
OB+LEcsFaviK97XXzoLygaaKXTzyj1PiDDlAA0MFb65Go9bL4c7TiBLZYuJVuFYPPF5JyCaob9Gw
GzvaPuxY2VTJTshwyudpLq83FgAiawF7lYt1AxyqbI49xBiJu3l3XXM9DGkNdS01U1gk98C0VpWC
vtjqyrlaC7AEMuO8yR8xgo1nwiMpqcXLp0jkh/mZngJeBJUn99acLFdDmTYB9nyngPl5+mEY0F43
q2fc3G+ECJtWpnPdneQRBj0Y4G3sKKdpW9OlpH985L+t1+sbWNtKbxq0Pf+VPS22n46AxDB8gmyB
iPC/ZYBm3EDuuZySAMom0FsTqEQ7BhkizC0DIwjkUYX5/HIF8rCSgpqefesmuhUUmwFMbfbIvebe
/LlJ74stehpuATv1uDdbJUyKfu8kNqCBRoQFuMM11AELX0YYtZ0WjODkkaMfIC9m8KY/t+abbzm/
X1c2Vy8oCwRJ9os4rF93gSyi8Y1Le4aXBbpWc8L9BsBlSCjZ01Jqlq+DqQ06zFlLhwiJcRA6Vzfd
spaPyAr1bLjaKUkpJjybVnh22SU4av6GdQbcrckGuVd70Q2xheNzQ0yEVs2bIhP14Qal2K+6gHQr
8p47upPHipFWEOlsI00jspSEDgXLM0pmx6yONFxtbXZZ415wfVlTNpMp2mIu8QGmZ3mlHHnT49lQ
kFdBEGsZGGhgC6pBEfEIXTNEvLhkSZdqeRTc4PDgq3yZ40zDdgFJaJ9sjsMVDonvkUFCOMR+KIrB
pTZ/shIAKMq2QcsvradtkruDBEhqXwl2UVx5JvHfxubb/BtpqcWXmoGuLlLXze5eX5XTME7sSHgU
YjgN/z+Nz2wdldyVKZ1g+aeWNHVn6bK9coaiKk8CkVxQ0oC2RlLn8oHVz0e66nO0Y17X92I0U3hx
+7jEUrJCOmkLu6gMLk6K+C5SwAh4hTu/wrFgM+ZIP5/v7csbgeUZqKhm8+MTIwkwfcYZuEC5TGFh
UssG5ExGwpe4LX9t0vkwgbtLufBR86nsd7o8qRajxaTIyWA+2X1LHN0nunGpdjOo5wkupfHV58iS
mC4/2DMskhyfN+LnUBsGQSignWzorf5d0VphSB1u0jpT5AKFYirpGLBbGYut41+feXcuwMXTEzVo
va8EYfRGFS5oNDtS5ydvsMK874uUp6s2CfMracES4aTQZzPwot+YFyBfiQNHc9gYQzotZerCPHFa
Ush6sYYWWb0iB987H408s1Y29hHQsBemUbFkAgAYrr6kUq8WK32EYRe3G8L4LzeGIXAynQQOlTW6
CYswRz2DnLrTKBv0Lt8M1olkQVHvLoCZvBvXJCeP2k6C7Z52IWQK1CrWWlS4Emddgp1pgM+R+LdB
LY4HsSVsdIjWeu6Z2BcT1p2q31Z7ffotkBiLpKG/6/YujOp9jvWhMSKhzlcgt8VJxd6U873Ir5QM
SpRPIbF8rdZElGmvhymQohejx6UKruuvBZj0lgq32FQj97c65l2hmLU1gyIiL6RI+kr7rRdTrDG9
8ZfUPSDf7HJtD9Mn1qoSxqx8nRRhhFI8iJt684gZm4EwDmj803IzbjaUq/rF6R2kkDxC2iqYsiGD
EqQ/tZM28EQxxPiSvdRVYhh3hDHkUO7DKLVyUxFPIhOoth0amSA+RJ56e4JlQxds0PPKzlXsiJnY
X1c67KZCKEmBfWKveaPRzqsli7wFeajICNLRE1tvD3EMt+8suiSpTF5CIbOioNEg+6yTw/o8QSj1
AWLziWyOHIM7S/rtDf4f5IxvuilOI4nN9u5DoFg9SgymFn3rlnx9bGjzyVOlyqRYJWSFEgMeF2Hf
eU52kAmlNqxW69j6uFBX17lcuInKatpZuVjFlANsbhtLcDuGJH/dQQs10lteJm4vDhx5UUDEsmBU
88AlkzyjcwQL+eKmTe6pZqC2XlAhJaKQ7+pxs0bs3QOQxJ9R0l+9g86mLElQOH9vFaN6X6zyyV6Y
4Y7kwArfrUJ7d6+J33QbSKHkaHGw2xC25LIlx/u3tZp0T1I7vsTyGpfOY31sRgnlzYnToFYC0ya3
YKbygvEoylfPKV2PESq8uuu6P5HmXTbdTRk2rxNR/Enri4ozIpmmJUR13weOOCHOYD20QczQvWoX
4rGSj8N1SRt+/GPMTu8ZZx4BFy0gGtDf6+lM/8iW9rBcw/6NmlFo1+oUPpIREV/E4kSpwLXgkqhm
Awt/FfxaLAXI/HeMw0UnSNQ8qrdT3QxJxRZLRZGQjjHItIB0DwuANx5wbRHjKfm7mOVifRi5jULm
rujx8fQodpfQeqquD8vMjNA3DwI5MpBkEFCcd8WhhL8k/3AZmKnQWjIHT94bKIkZijZwuAooSO3K
/asvriHXN8KBAapKxz2k3cZCaGPU5oDuHQFsvE+rNzU9dlwlcVovz81FM3dRZWW9gihUDK+aw/89
z2f+xPkpsBjhziZTUMVIMg9/2cfttACMqvThC49gWTRjOxpChpFbBTmSj6FkMA4LqolFy7gGFkCt
CZlQevIpIMQdpC7YGY1HuId050L3Ajd9MgvQr+S92ofgrAw1Q3qc+ZYE8wzs0UmPfMCVI5hET0CG
T7NxZqBjEXEgQ72/+4hgY0RAaD3zeMhPjIqLcmpjRfyyTA+RvQN5UVwIWRJXWlbK033KoumpAIVi
QawAki7FVT8pvnFxV4zNvYwDu4d+vCgTL1pgfMWiyMSmr4kssAJhdIOFLws+r/Up7MhrJs4J0Byo
4MIfcnYEzQL33KC5cLsJf9cBiZOLp0RQjAMfNdF099es8hwRkjwnVwmUG3QbbZTK+VrwasyFAtiT
toaA6HFSDSCkGxmCAJKQyTMCfVHQl/2lgNngleAMo+XnxywZLCqysHbs/6PilMWRgh7OxP8MWz0X
2TjBi129M8n3EPKlzRJYxcmJIJ18TYheObl/zjspMNzjHywEZSUAVitu/MA9nVUzJojOO1QqdGxx
XcDzs4iVge6A1gQDxyFir76dMBzj9XG9qdFxScd/yDwBthmgsLXceVUJVT0lUlZYG8yTCIRc4OYy
H5gtkgXKwgy6Ynr+unuXumsxexWs78Wes218RbmWDeT5WBWxHj/mlZ+KNvwUWZ4GylXCZljs4yAA
rvvaGIp4YK/PyWa4CyP30CzSisUJkuw8foJc7QTRzZq4LLeL0F3pIa9q+W3hLo0pxGMPkNemeVtZ
sJmxUWqm+mytb1shYMqoj3TEW+I46njad3hvvcHhhtzUZhlY1SJfTNAaJyi/kBxgwc5ebI2vpCi8
CDjy+LLadjLNWkGez38xBF6vHgTxZzKlc4Cxd181tPptM6Nu+ZZrQRVAREw/2Jw0VA/MFk3D+5xX
TYnp/edDWEEA9ggNV3HlvxJYYSJr79sJV2Mwy7nRulHDv4ujQKZlBeqWHFdSE5/1TAd0PHVoAZsA
ANy7wB526OCY8xgnwHmDN412yG4TfmikPlbxDl4ChIncrmbEoCWLRRbhsMesbJLNdRrjqpsTotGt
kZ5WsfaHRZiOUKKjfdsRni3JZaIMcwzoAapQTeFlDa+fEb8zpH3uzGS+Utts5RTJlaMnQXcV5Ekr
CIJL6rhc0xytVi6vHVe35d8qt7eW7mfuj8QMFQpo3m0GlgK04sakVGhHiZTRBFTaZWvImRq6w6LN
xungNDAXaRyw7dngDg0vYBKQiwTKqCr1ll/Y/kLE/+CizsgR4pbEvHcxdIEhhwtCR0kn6ig1VabV
WBHUlw1KjgcvvBkjSifMC8l4szePtLfng8HV4yYeKaQDcohijpgq9BjDxBK1JA8r2E8zKTPgJ/3p
YVDriL9JdskpKWJBbzNw5iNtIXa263M2XuP6/za4G8hVGN6PyjeEjQciALULqltG3L9wH36Kmgsj
JssMNRPQ2pFz1Y6GyNl5+Y5uJnqdEzQFb6CRhSVK48lYgIdF9grMSQEXKi1t7NrkR4xOgnLysJru
NzFUk4yABZCZkYlyyXqThWNkBpFg0+5hUEcI3AZNACPwVFNVHIfw6utjI0KPQVGM5gWFZGctL5aI
mhss9zUbWWZeyy1HgQUsy5foupaND2U/Hxhf3UJBCRzYwDw8V2a/LjglvH+f5axtqdSX132ClQWo
XEK8Fn1W/DfbQsH5vVCrMBC+8ioR05jJcsZcOStBJEPEZB6qzMNi0Rs5M9xKTt8caydL09VsP/pX
/IbJpP8H8HgcsWqerXjwbjywjMfEhvU2ZdkRZtDqdgpJ74nLVXaqbFNZgh54eq8anzCCC2SSFOZd
7iJe6eLKV7MvVCs2cHWbbwLarChYa2ZIkTQuFfp9AzGBt68lO0y4Gic+hkgKQQqU3MYgjaYIKePo
DrprHPTjwkkbo5GOXxNAcVMHb/PlnCoaw+cu8wvIbFYWhwP3Um9y/zyYQlhCkm2WTToPAHKmEEm5
pbPpxuJCpfhEK5vweKsR9UOepKqONtB7iiPhnVL6v8J9/vNktWC2M2kOy3Lis5VueNvTeUwea5+N
XFPItMvEd3zyAd/vC85P5nDsYH0C43VBd0QqzbIdsS+49Xenrs3abf4tzz2euXldMnJSasSGg+EZ
hCQUu8C1xgCbj8oriBpDUehFQENbiXFE1KHuEmTaHSQ4OmWA6a90dDfIn724BFi6LyvT2gQcOYtH
2rooJ0MAbPwh9jlz9/g6RFA3XwdmfhH7jhgsjAtU2MzdyLqkw7Q3xMxQ54YrBDU4IKV0yB2HX1hM
q0LIUdof6rcoSoiCjwVBqHYjdsyvwXsFfdVtiwSWrgPzRlK/UXeOWH574xJE1oCrKJtwuhYXfz0g
zXSwL4F6COAvvoMjeIz3zWnKgO7GH3R7WljRwwTVvipmLaIRaJ7KNq+pGZje5nQF6ll7gf8k8KW0
sU4Aj4YIZbwx1Z5kmE9rwKNBPTiYjlWylRPvCcrvIOGh4yscWBx7JROkGZO2hNrnvCed8Et6IYst
8vwmEDtnYa4nj9NnoQ9GoYU3WbCK7Eid9MS7dXL6O8hK3rsw4j1/bGjcYR/hEc4EJEkKXhGO3+Cd
E1pB1Ucj6kPgqRHXy2o4Qk7tlX1G7rSpRDJXP6Fce2kqDn6fHCmgMl1NdHmgkbzg+OyiNPzkfi59
1RSW50RQnYI1qkWQ1RJnJRsmP7jl98OoAOVYf++PcZ+D1W57my+9JtYglBtvMI8i7x4Ers/hw/37
4A8bho3gPQEk+EhkhmP2p7tw3M7XpFXIFUxGg6vPBMVIIfBlVvSQ6FQ+dkgZ/uAfWBgnF1q8GaOi
eBFgwfRd9YOXinvp3jaIi6cPlUVVaQPTt0i9uHuIdVVzfRMq85p3v//Sb/obH1VnvNdCQCoPcM7w
wcS5n/8lJgLiuOJ0SBLTfJG0AqB2q3tpg09DZiDcjRYBQVzMpoCBpSGhUYc7AS63VIh6RfQqKXPC
4zYo8ADRipdAQoO1qLOPoI0+jguk9A50+5taSE5kAuF0gVHYruVFNCEVAJ/ut3RAwcG0tPh2aMO9
K/uWN/TQHth4g83ibma8THEpQqQ6UYep4czSu5thwP8LLPFJD3qtLuhS1WHihMCQXhG+/1tyWYWT
mTidsrJwwSZPBiio8Gin1ghsQ7a3lCa9kEAHbyoDu2vhDukDSkohGJ6iw7YR5I5TmV0bxpOE58GG
122d74isWrST8DcIlg1QJvecpHkMwvRopCPwbu8Q3pzA5bA25Oe2vq+odH//OK92NFjl+IqrTwQD
hib/BLx716EETFGP0Z38bi4xTQt9GstawCTGxvbMrgO6o5XFvS41B80KwB3ms74iCfXXfuthkq9l
uQz1K30RXDcvWh7rGhd2jTkP0qKsWqFx6SZzXY0TnokjGRZB89zHRforlaBmMdoyMxgxVkjUDOPj
4LaJHtyP29vosBV7qDCJeZwFCGA23BHBFYkUOvoqyOpJLly6/GHAgtM7lWWB1/y24IfXTBZGnQIk
SPpWLkSCgUvy9/j8MWkn4Tjz/qDRvmwQVCatMwZb6re8in2isGbbtazJ5q2b+nTuOmrS64cNCUUP
WPU8s0VRU4qkPQm0exYQkY2mezXNpYTOJlWVuFrTRXtdapSEkbZgLMRz/8bBxI2KB848xs9XThWV
Tc1ltrAnVn3EYfiCAF/+7bdKmvav3J2Ggl2CAuCvOKNnn82QBOr7RJCqRmDdHNfrKoSRer26IWJm
kO8EY6P6rXI6YfWZFePPb8yZdqNMp3WBOukGvyY0mn8OTDIQV0YlLPpz6dyj9z/YS5VKAB/GSATH
TUqT/daxa1Xz/k57VECWWSbHXB/GzNN8RZZywQfxpSZRrUhH3Cvu15ACqAnO0H9TkKpNKQ3h4Jvm
sKZ4W5xpiwPVKBL4L6Bc/qhi8uqNtTouQ1jiBtzHCJlso/hDcRY5/Z27AbNz6nOIT6wNybXPYuLM
Q9A2veWL6ApD5yp7xiVLoJXOg00uKSqG03iUAeYf3jqp9bbi7UVdIJPJrK6QJ0fQHLVjvYi3JVpE
WJiSluXB8ivkkB2ylLb2KJnhwCTeyLVKuEc2JBpLlR8tv/L+yZIqybcXSTf4sydS2KL25rLIlRUR
93NW+q+es5QOVKaz6sTUEZblX5U8etWfOWYVn/fF51EypKgeE7OrmWKJkW7rJlIS+lspsat/LUqf
iuHxFTi+dlxH3vk3YzQkAMjKe1wQ4/l9XdFQs/6lfjT7I8g1RE3bBoGHeBp0YpHvm/IkAoSbfI+X
NSK2RhD1qUq8jCrC+nIicGIlqs5aXFJ+2JyANpgA6PkuTD5n2YL9f83w80NTCLLhg9Af3DNLBfAy
3HxWbT6qv3unUpJpg3bHgbXsZdkdR9RstLv6avHgTQG+wLG1oXbvTslwDyCdZ+50ZHPFnucj82rk
C4LR3GgpcVY9RQKrdD5XlO+Xg5MCDXJ3Gvjv9gKuKErERZ5//LFbAdoiKudygTci2uVmAthQIqQ/
IjcN4dh5iwlRFbI2aEVbQ8rae3bNJ5//xL2ydRcJ+PaEhdhLJqNQodkVsTZ9c9AVjr6gl7VYQRA3
sqKh5RcDVC9vvfNIg7CU3fJvCFOccJavTrokw9VqyZsrwsTm7Hwx0SC/nk2AMDtmDOjxfAcS4NHA
2nn5vjmWTXiWnOWLt291dPybcCdwfl9tpxLsyLJ+ShVsL5BHrcBEJ/23XHXzV5yqf552+1D8rcst
zZKVmRR6aelZV4o+qLG1xJqoIRHveC33MCNzuqweF7QXzT0/I5fvBgd4BFuyTrOnA25rY4s79aLB
6IVglZa6+hmIu0CC7SD+4YChvZ2nlLXWZ4WP+hwNL/vhCrxv4YcPYxAXx48DGCCzD0o6sTagwCae
TT5GDm1LPB3YCWFL7vuIPNuFWobZDegXJLQN2I4CmpZKGxj9vWIfolH5Ih7HjHTR1yCNlR1z36GT
8RCyHZSre/pPKHmnxJlCXsFswzVMhRgZl7uCakIxip0sIC+HrG2ZJKuVS3IlWJ88DBuogWX13x2o
sppWm3CfoVbf4zYJ7gUBU4qD29HXGbmMyqdxOSPUrWusCheu6L6v0B8up+bp+s8mwB/oVQZLrIFS
UgqEGZL6l2sKOZcOpqfd56QXO8uJve6Ihc14cU3KTEhjukCZm5rOCbve3lyIaIL44egNTj0dDbCQ
GzEQebeknaqgB6XGc0K54c9tDV7rEH3x7E7ljOnwFkjJjwGzwwPFKV7Q5GltBSD9arWM9SGufVtc
Cv6L/p6/eitsOrum077tBO56NqkRoarZe7Ggo4IUEWXZaRcTex220Hgo9ZPo+UVve0880nxocwcb
qkgECB709NrFbTg3aXqJwk/9TtToUtEhPIPw0YN1hF921wNCc78Brfid0ojqrV5BJg1OvF/ebDKJ
U0xBxUvjRZ3jx4+HHhA8mRUp2zqfW+UzMk30/vd3DTg+VspEyzCVutWAzNzpmEUAi/Ii6gbE8mGw
fqbzAcCg1q8xTPR3cM8wlooHtiS0eF++CHwyMUwreCW/GI2yBA/7EXtEGqDQHW+EVzirViBXm5Ak
xzxVWqnruGvXlM0NofWnaU/rgrcheTpudSCa76VkOimYZR+P+SlFXn6zSoUWAfZw4Ck7u32Md+YG
YZoz8i9W767pJF0DjjHKXCVAp0TU4AmMcjcBtBdhbUo8o0CJuFB/iQYFKrl2NLWTcrWnQYdl7KQu
+QC2CY0sbgGd7zR0nJKVZrvEIutGU7qP79ciIw1NuXkHQxjYrZkTxqpLSt4ENz3pxUjIuD4H1VVY
zPqYnY5sl3D5NOAjWucICcMHhVd88rsudIukj/CoMylNEZfYjY+E3sZahty8WKcQ+9L6qEHe3Gt6
LCwuW+3WoAMud/Pr2saN0Wi/dvRgNwCDsNGKXuj+EF1H6R+8vPUyw+A33bpS+PI9x31gezAs7EYM
UXSnBCDcfWDbmO0ZRgsBC7Wdi2cx0bFy4fFFjCWfeDOqfwgZUjMVBE10eBTOZ7HokUxlwAKDV1FA
DakPb0QBuZeoMqr+C5QyC43vH1T32FSDkq89MswLyzkDfT/v37h4K9+0xA7K+4JtJpJDuMMGpDXr
GJ/OFa6IoJ5BJuYiFS1YpQEtPB+0HfH78GLCICSWh89bpID8pxgNhSBLEZD3KYOsFJNSfuOQg8be
n0JhF1dA+94yU+059MLkmbxHUaI+g38sjzN9wgMc+/vlMUwcD6z02MywNWZiE6TlAUwlB5+reFpC
oNuCl7Z1ovPu7N7S80LjsOIuvXF2oZ9zGc9rakjRAwUqFx6LsU43p/4ivorYxYkAQIijzOKCfDyD
2F8S9yJ0E0a+kAhlhxrtIjUgCkW8jwhIofvCM+46sWjjkfeEW8GF8vSAK8oFYhdMBcroM3HRtj8q
6ZbmTwq7PE0FCE1gFzSmz97WNBf3576fNbmgvkesoL688uLN6AkxUeHDFDn6Crn4Dg3w1nTDeJRC
wGOZfkp9v/fX43pJ0kjpPlwGs1I8yPK+8mch80jnzUz7a3TjcjcAraz1G8fJ5qiFXLTrtDfrQVeH
OnMZa+B5IPHIGoH4UlAdvFzO/JAu+ewkcRVZRDfqqjSRf8nXZZ6WxCHgrTaEeIds4T0AYyunxejO
5b1pOZb/aR1zGQhXuK5JIQZFO8XFrc1TyOw/94rjQEjjgmJOSX4a50Zeyv9upVqyJhJiDfeT36yi
MIwhptJj5MqELwL1QixnOu6Moqn0sgm5yrkStHOBjQrkhWWlvePwUU+bWj6k0ryNhSG/r/LBLq+n
G+ccrvu/musuV19uEZc3XYuxQ7YcK2Qf3qBtTaXlzk22xzEkKsIb2WePGwHn6J4pM1xobWMFPsnz
L0HS7jpXyBl8u9ltkTXDnLiLD16yOuVe/3/pdX5W1IgNyNhX5WcpBTLS9I3FWe8RHbupkTb/kcwG
onRJy7rKer50W2skquIZgrx4IjD9rLMenfDOTmlapgV2tlXSJ2vt00Mfae/ol3TWHbGQNMl6Jpzx
4Yf5O2oPfRUrHDYwU26m9ND6WcHYHtpW0OOaWOUMwQrwAyK/DoRqSYESlf4Sy8MIVOdPejR8/IfK
YDm1L9EuNAUkacFw4pvRGZo3Wsbscqq2t+bVoXFQG7YdVI/oWPvgLxeht4HrpDp6Dw4Bpg7gouIr
3LqEOKfPb/TYSlhtfP5jkLIi90po74wpbabUch0pwUEnvclNf4SUTvBYUutEm0tIkkCVSm9QL/42
13DPSFxP07O8gB8f9Oal4llHzzvwjYugEbqMzqSXkun62Qyl8H67oe5naom4JXu9RdS3DJ1Jay09
qltDEmh+kVIX/MkTNtdXraOU/NdpBhUdoW/dj4irhQqI9wa8Yl6QHbQ5ubuWrlz96sTWVxTh42wM
S2odv0Am4ldzndArAcwp/+7Mp7IZssj2l/f8+wVBLq2DX/ytCHSAYuVJSmGufEVDoYjW0rBtR/Dd
dgGfQe0tnh4guQuUmiNVdxerS87efYDiTfP9Q20l+a0OQy0tqLhTbtOL8mft/eiaBXDVz+i5DT1k
COVMFLFISYJPLRj0rhKYyFujDZ5m/qsEIl31PdjQ+MHXvp2ynXKWSG5D0uJmAEhxDsM99e4qZzCM
fa3vv8LLSrUV1+zki/6Vl4JE+20z4MD8V6F+/XBkOb2HxMI5vcxhmboWHx4To24A7F/qGU28l0QN
PxJn5Jr4ezn+5bS5cKMko7HxLpeAeAKLo2JVYfvMk153N/YtdWlaBGDe856YeVVUYCL52iABGAVC
kL2p6+Vgu2s3eL+qQJRcRspmZqe8NhN1Ay06d0veyr9ea1Qx0/OZYHCHKMioyBLj/a8Bze/xVEYM
sXzHCqoC9Qs/x57NZ0CQABjr+jNsnVk/BSgwDhhDaiXlfM7Qn63POgwfgpAmoGUrVFVZvNI9nJqZ
NAa3OsCeYZH83J6AAWbh0KLBMW+6fOWWtvS6ae6oUh5uGforLyQ++jzfT+lM5/fVQHX2jdAWlMAq
dIlfYk560hoA66L7iTkFSIylwcuY7RQP3m+nD+n7v63zZLOvPvTP41n6fZEDDDyVI7DtSUWV+G7A
anYZV1Kwz7sJ8KWF8nM0iobSSkXD0pgc+eIvHYOuac6RFGtwy6mDb6v7HcrMYlh0/Qf+BXELIXgi
xaONuk4LeXpkroDMHmv1RiR2YRhB3wmq5lOqqg8zmUjMtt24EA1GPlOn/P/oIZqGp2dgcFAWRlYR
zzsCM/biQeIW69mrVcNY1oO+85StGaelOGVxSsw+vgmtGww/j2YduDLb+NQUrYRTAIIMpEhwVrjo
VLFyEqpqEpelrX2oiEhEH+ktgXU7UVMORjGlYtTlALzwGFh+iR1Rtuyz/UzOQJbuwKKBzAYfuR4A
GqEsQM262cLopI3gE7zNX1QQyJIXeGziDjiaLAhSW2SmF/1yCXoQb/5BUdrbwAByCmwlr8hKY7qL
8uHf5u9tHA9JTgSUUhtMWqOq+Co5H8z3X7KAPmWKCuuTRwHthTXfTAT72MZBlE49GERJk2ozUi3E
+rwp46N2eWU03bPB6JeWplTRaQpFYMBLdoyeuYp6XCK4QHph5BTlxNUjAd/QpTLb/8hxetwEwaMy
BQfuuxZmV9xfvoUUbkiYAgcNLFgbaEDyDoPzdfmbl94YS2GtkA2Px91NSPfdUZYnZ52EOCz4PGmJ
MiiB1HGQtxa6aUSm6yleTam1WSN72hehFPKczwUBFEa89dIFBchcKN71HA0mH9427TpFDdHV/6Eo
/++ma4bY1Pg03U8BLbFP1DCVG4nWCoaYZJupxapG0w8YL42JQ1U4emHVNpSDdde+Ypsdm7UKNcVO
/8ASg7b9nelCQ5m6Y6AaX7FlDsUwdFgCdhQ1F5Tn7cDM21NphXpKAYS5lVu++CLM9DpQIW7BtKQd
oyxlrZPN7LN3n4KLN+Pi/Jxt2W7xiUKAw1pUwuH2YmDF1bf2gFHuXuS3K7plkNM3A3fMNf9StbfC
K+1afnbMJTyISZjYyZPM/9e6bHLPh4+0GETrIkc5uVhKN0Yx4AwiQ/WaYTSQ9GtU/veQ3HT8rpmw
VE8J5M/JQ+1yH+O9N0Mq0Iu7TdbU51OggTITRbTz9vLkNbAgZB8r10H4VxaTXoc71p7NMfnk0uKW
dkzRcxwekBYSabRNSO2xJg9ibWHDFmuAQZK7WfSLbV+ytxjq27Ffmgob0zlYKgDBzHW4TUvtu9ef
IyMN41J0xP2tzFw3KkfUtiC6vDDnw15vIFNu3k+F3X8KxkTkxuK7AG/tRivkyk13rVM2DzVwmfRn
Y/tCI58otxnJ6DkVSp9dT7Ee4aHg2zK5pCXN8olzN3cLN7w19LKvQ7buwRepRY+6jS/svP2pC7/L
AxCqroqiO+Gh7PTmArD0OoaZY/Kq6MicqvM0eDQSI1RGOaE7Je6/lzU8TXIevoSeUM3+lbQTgrgV
QPAuMNH3QB5VEmSljVZsTNuf0r3Lj1diwm2RE0lIw9QYiNyUQDkT7Dn21CQ9L9LLgo+ToqEbAeV/
qo8NzPy8Cxj3JJe1mb0lKOTVrn7lm2vqL0kkE51kUFXXpbL5Ol4je6HPvM8Gk7DDAT0HWd9QfZiG
ymFPDZoUDWe/X31LlwXEhtDQaznUS82TxV9jeV32H1NJ5E+PGkIuZFiC/wrW1cRWQ8jdm3pEE1fW
JiGSOPJYfIxAYgCleqdZmsY5ojTWgNUpnHdmJUUNVTy3QT/SPMJtU6iqVqEK7hevShgY/FbbiNDd
TaTfXD3SqQftXSZ12cMI2tNOutpRwPDsTvLSkO3fd6OFVA3r5e5Q3e2jQmXIrdeXrd+Bss4H4y8W
3/BeLOnbYd+SyfTBUsXIEaOGvnxBDZNPf7wm9EcJ3vVe3h6qbW2PEcKHDWKDvDKKcDvoii5Antmr
3koMKySOlSgpmLb2V5+KOIk39o95/5udAmngO4+Ps4OHkLeXa4FmpVhad2sbkxPMF7BDIBPM/QsS
Xsamo9KNBzD7cGdzR07XzxLLnS8cVxazngO/aKTGKAUgBVpROIvv47zdtPO3MqY/Ei15e15ZYNzv
VCf+Jl0UqtjryF/TxifjMAfx+fCQECNb4tdwYqRuceAiT15a5iaMVqCld3vbdzrN+b7ez07TT6Ax
MZqeE6+eCki1eeBIBOdysbdTj/aCV9hhm3J8qVnRkiPoKcF/9Fbw2kbYC6OGX09YPSoTgZBwsiMC
ajlX2dR5SSH1Ti+CinOl4lFx0HMzDPKx8eziUP6AFuvbbM5Wp9tmkO7atg74xfKRSzyu5vDWTz4x
YpDWmK0hOnCQQQU5/BUTy3tl2ZEnjexRWI7YHSdC5jyK96i4RasIvFtl7wxqZMKE97bNXDiIASEi
8+QBkj0fR4B2KOa6V1UIDpkwAlq4c4Dbog+2PL6SgfSTEG2V0YNhUeuSpKtJKdwGruptx/wcxnnh
BgSwLPk1KAlRvTO2sUvtauc6GkdZA78p0prPijWMs7uX/TIbnoJldGZ2sqh48qxsdSy+vZx6v22Y
TN2Iimmhgw7TNtzqu+1eJjdXu6JV7Wv5Equ3mEC/5VUgSFxZHsVzPPXZVmL9jnGHHSF0hC8idtRu
q+GwkInTFtUXe4kRdWp91p/GyU/6DOB80Qe3XQ69rlm+Z6XeLVmSatTtbTSxHgj2lg8HIojSmzHQ
AFQ6ghWdy7dhwcV5nzICHNf7NV7UhNWbA10YKXqQMso83jfK6qxOoNYN95QMmQao+OSMwGNmNRAV
00OoAoS6BMhqct2W8FtjuxEv6RYHN7fsW+Le6V23BdgrC4zj6lE0L2dS/xK8AbgmWIE6/4HDySWW
l/nsv1nEY45gqiW2hyvruo2nS7z6u08mkRxugEcw2oP/HhGurnRE3+yHFtKO6zVE5ZAUkOWP53nA
xSfIRoA8ZRNRHkZ+QDVu9xOAhQDLUmLNdRsUflNmZNqrVgCSA3Z9cg3ikft2ygRNzo4i2/5WVnZC
qDS0eYRfqZkqX0CnCzFnJ16KQJjfpY6nwNu3MwM/HrfAmusma9E/jUr7KMB3rgWAlnsCVJxq+PXo
0MBPWykCsZ+1EHRoUSKBrQHcvj2D5YHvSCAJqDhPu1pwyOWWzo1LiTKAUexX6opsuPDvOQ4jiozp
z4rJ8fA0JZkRLXpplPAYwFHP4e25k5tDN5yqLi8HGkFFaTRzyBbZUZGZVIvuMcJnWNi1AWg2lxXF
Mla4lpAOhplbi6v4wCZMPfFHsV2K2cZBKef7DculGowJhSlA5zSf7mQiBkMstqqgKkQh3vVYFGq7
F+RW2Pg79fC05K1MlzIvNFyYISApql4ri7mgYyrJywy425Euu9ZjqB1aQm0E9enNIRula4XaObwT
jsBEYqtpjguYBb3sNlPT05q3Zy2U9KHEo7apICUyBj34dgszqMGO6kxpWuNtYB04//KX9KGrYtdn
dhApNQrzjzWS9WQ=
`protect end_protected

