

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IkKQ7UnyfG/i0Gz2KESfn5rIa2XG6JjMuNzaLweotYfssoXFPRW5MF9/SJXIBGc5jwrrtn7ZIvXw
ZMKFyJ3FzA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7z8fuAKplZhDCneI9mNA3lof0N+J7iQN1H5R3Mj6yF0lZ6gCWQLLnnmsEoxkSX05NXSzlh4gcEg
7rRfO6LtEEhf+XGNB65vpBYpfhGyoq59NAHhGVo4SvBM+mv7uMxOGdpTeOCZ4JbHV0AkjL28mjov
93MegfTkvdkm8J0Lvdk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xuMQUwo0GDzI3cOEq+tu/2nUcDmn/7fhQTHPWWNseJwSS2v3l/iZo4evCcnhY45ESTueA+ZpjAko
WVoSIubelzbNSlntY2uMGs5oczMZtiztniKkMtgrjy3EW9dfGbHhtmNrOHGIHH4IdMr3kAy4Vh74
ZigAJ9A6+7kI6MsJi8v3mT1ARZHCR6MWsQMcVGsi2drnsGRWoYryCO5xQR7B/cwBGzMymTal23NM
pQKOm5sZ3P6n60ZuBiOsJmbRp0+LVYxKNhFdxlNXd0mwyAZQT/UOuOuVbjlNnKY3+syFmjH1X2jU
BRKqD7PfkYIVMVQ6XvOwQSNLyki/t/1FG9LntQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2lTj0FQ90PRwxkOhP58Pis/0pnBIhVIOGqxXo4lWUDsJI5sRS1Q5L+Q6i9o+BNlX2LRPYus/9Dnq
5ATglZxA4PDv34H6B5xWMxj6PrHSWzf271mNIoMFrjsSBdzp3H4BqkwksoU2N0BujU4mvFktBj6s
VuYwP8rZjGtZ8cTr2i8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WKc7lQN7TOvrS4DJ7NNUxP98rrzfIQuz4DIZ8eAY+GKFx6NuoyinV7kCt4N2qBg8IRnkz00LUdTl
h4FZuBrLJJyfOOGbqIiZNIhgdqVi7fXcxV2ef2SWPHLvr6kIV0N1TmRIBZht7FPZCej+/BNW8QYG
B1Rd/mmsAB7hXx6GfVQ5u7NRsVDyxlcEghLjiM7GAdTaOWl/F6pDM3aRwjjOmid8Gt7xmiYfPT0B
Gzk510O+OqDJRqmdMvwBmv3K/y+M1RxYsLOpwIle5lGrJoXR6zj5dZS3g0EOtylaiuYJczAHSe89
8ncn00hUVfz/5JZCkfgcxZH1LxGTI+Ly2xY+5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8544)
`protect data_block
9hT+1J/QfpbAtUvHvp09UZyXeuP7c3GJPDP6O5igAOPLQFWG6bzjkvkKAvS382FP/8mbBnqeaOCd
xM1eTTAiuGk1wSx6jpmULq+E+C0kM3Mq6hpHEjmLW8hpb14E4MbXeKztRCKx2WJJzV8eXHZo5QrG
MA5DDdh4N0nw/e6HZO1ajW3BBU6Mr43raOP9vDEKHD7bKV1dRXRQyEO2PqLIUkc1kZypZBX/plrN
hHB+AKySCk8QLYtHwiN1W+irfAgqHvaqwARSgYvVrg+RRONiwxZcHE9n55RZ2WA6ybPbinmPXDhQ
aXmCBT7NZooplNOIHPjAu6asTgA40vHjCaYwsjY7KSKW5ieHxd4Qc+mt6kC+BcACwgDatCTq1RyC
Cd+jTTBRp4CYzUDqNMQuhxHpSz1WahW8lhea/zH68+DUAF3Ad89A2XuwnxoQjSdasEqgF22TJSKb
Re3lAZ61b1OX1FhCoRNNUApICHAOxUl6h1e+YNA7ksOfTSXm3/jeezCpxI4q5HQGGjPZcMaSqHwZ
cC3xaSUZtWmSKSFwUMJczp5zKhESVZlsGxSMdFX03I1KshR09JWRhxCDXjUt/Ip/ze+cslU8Uilt
BRWxG8wTUPaAwnnNpgaU/8k9dBcgXktYtpcNbqE6bTRuXWuSXWMxZFnn+NZDc2Vy7mH9cwR2ObFe
c0jsHp6Ymw++5/YDQixyfvLtqV8x6dwFkxCA6RnE9c32kgk4m9mxbnO8brm2lNz1E/cq38Z+0Y3L
Gpmui17Ni76RPHa+vLV8Nh0FYqxdm0AO9jYzOCE3lpwP++0AX/9E/LFtaxLN4C3G+AW8tGhLRnqY
WJICe4ECdl3TB/0Tim5fNoA9QkcwD3q6B/iGc4YXTOk5ehB3sKjn2jQL7xSNWU6U7aKt9wc4P7+6
inc3TjRz3UyYwNbNm21Vk8GzhiePEd76tDoUyIeyl+5b/7tZ0NQPabQb102/UDS2jQCLU+3CVbXV
Cjz3d1qXM39QugZPTNfU7EGozW6ARnRdosVgv5og1WzqZqUtucBS0uqFbMya5va0b9lic0lhvlJE
CdvHKaSW3jPkIai3N/9XB1w57lmeStBKDuhL/oH5TzeLTSXo78tWVLeHW0nLgjtapDVjRfd2ENtQ
isEudDRCQ4MOCajI8VXRmiMTsUca6JroFLBAkXaL7c9lwUqQd5KgZNcUOASwVFQyliLlxilQJ0sf
wCtnnaxCM1Z5QIlYAARuSrZZLpQnGKd/Z/m7QzxB+S96d/rv10p+mdSN3pmbYPHehYyNjcjnKObz
0Yl3jImIAsbpnYxIyvQX8x87AAC78hJJvRyXpT6CpAzmaM6eiRAu77UWJp+NsvkhAgdy7mp/L0MS
SL23fHn7LNde8ytmsiGIbjNcz1Mxob2cC1MnEsxXTuDfPJc27foHlGDDepDGYtSJYzTnMxX5v4DI
FjOVq79x9qy1QuvI6EZfRdUgEKRLUc5psc0gdJogNCPdzJPx+eijXd1rqSdAEvOUBT85dBdKSDt9
de1e4LXHbvCNjor1SO2lPUsdcks7X4N0Dn5ZGem3XVNSs2FscwcMldEIKYOVIQ7nulciqlP4oqs9
g2P9yQnp0Yw5w5CzWMj2KUu196u9zJjHBDcX/QclKBqVLlagus+E2YQ7rQ0gSEZoBgZBkyd+mX+/
72tMqoK/QCXhEy0f7K8QZXFQ6BVj8B487VA+dqCtNOqkPJ98lVO1X6CeJhT34cR+OIlIKT6Bbeyu
T7cdXorzWf8uo1rw1OZd6uwX0bTvKO745fDUnSDw2Cb4CD143B6r3r7+4OcjV44ev9q4ukHTCthq
v2n5KWalGKyfvAfdD4E6xS8Nl+lPGO+wVcFM/ybtsJgfa+8zh5/WTumBY0/JjidMGTE7RU8PuMy8
51VGluvaoTMouscKMIxpVdAJAr8ClLbLv2NYt+0unyECsoFRUaHSW7GnKT0NWAk2rBsF4HEF1nBc
6BfcvBJrz3cvXoFWBV2mmvFpLczWmO+wawMeSJJ0UNcRMbNJbUXyPxdhN0vtHBs/G+QZWzWcWvHn
SLsmsW73fCLzDw8DMTR4muEIWf9wK2Mfl0fSHU0e85rWxVZf156nCbmXoe4/ZnITvURxyucXKtnn
/1ltPjWtrZhXYnV61LPPasb0P4ZgNATWI6l8rS3asAZ/utzva4iBvPB8jxK081J7ezoKjQM8ipgx
BR58EwFcc22ysYhSJxeP/DGHMc9qNmtSNrMAZ6Ew3RBiVRsN/BZ3JX/0O4bOWdFNgwFFDB+VoO/w
u4aFZMQtf2j/1xL/1VykxO9fOegAWc9mbWH6maxcB5GAHZhOSf1/IyAij9hHm78dHMRkV/A4y+XT
QAUDmEG3wAumDCMQfe4axIqSJ/yZZTdVTG/upmHZnzkqGucYEoiyIf3bysBuMqAoDO+exhtUbqMf
r0ggkMNPjSUP3PoEFh7E+HjprhICBYYpehIdEMtgw93jpSBMZwykzp4MQX/Bus/eWRcZ5n8J8frw
24kalh27BwDJQVnbvUWgmhqTDKVbKkUS8Nsn5w8Xprw2WSWEcIBoz8Rzm3n+K3Vuz8ICZaQOiry6
MrALagn1XeThPZjv6XJGQ2xmZ1HR+1EaiUgllw/V32kZCcMuFBnajiYueCAhseuV0f2LQ3gUGYLy
xNLrUu+91g+cGOyrEjDDb2BybgVtUtY7eEfFBZUFkWrzrwEiFhTMpvgOIIWykvDeBPmQrEcuBifD
wThkwo8IhPdhBcpjq6JrpRGAdZKqpwE68nwhrcqnHK9eUWaWi4MbkkSQtoX18a1APaKhpKyewjFV
AwK7rTtz5pbXF7dmvsNZMJZIe3IeUAyTPyk+Y3r87JJY9xpfa3nOw4CHyeDiIo/bGe7AljXgPUrh
tY8pfhdfp3sXZToucz2a6w7lWjqYBIzbKixEnOVot+bf92bgYoyDvxEpC1isSKPAX7IxLjYkFEJd
riL5pXUgKEEzm8VyueMOuaI/vCCJ4q4l8dmnQnk3qrIpoFcWE2ZhDwiiIzZmtjjmpWuyMYjIseKv
WToHQ93RB+1GEMYnUa0EAYYbn12F1rNVExzgMlMhe8aIQDKAho2RvBLvV97bd6ZPZhoz6iQsEeuE
gJ0F1EmRzYmRsfQBwvT4C5nDWesCSci74ZJPg8yCo1NPV2YwdW6ZZHQe2XS2+K0unf5CMHZX1KLQ
hwPESPsJQBnmWVUM5zFzTawW1QY+4V0Kjk70+tjS1Qu56ps/BTZSJ64LGMRY0VVhsDX51VG0tLNK
gv316JJ3m2WqYGRu44TcsVpqEiPy/UUHLixPABkHobxP7s97GzOpUkxMNrW9YCSpJr9XboazvnX1
6x9A4ZgrDr8vYRTY6F7VA2LB74pb82f8PKDPraAwq04K99gHZ/B1ee2LlFQDw1ftF5oZ5P+Btx3G
oYpCocZ/rG3WQ3yZNu1t9Lon+w18g67tISlBRjAt18UOwjaT7jYzY1TQKfqPXjY8052FsB/4FaiT
thmqbbBf4lMgyidH0X00yEAE6wrQ/dw3iIFpxQXYkydIHl52vHchtCYX21IOCOK9VfLqcwqjFIYF
dgKtnoUzeBkRPVTZPIIX/Ip21Rw8mCz0MofWrPR81a8WGeBjhXoDAoXb/UYDdcV7VOQoa8WnnpRj
1l4DzjXYnTZY7Yr3dVNQEm3PCzLTrxbAbwxIfL61RR1giZlPI7Kz2ZLcVj45LxfusrUg0LV8b0aw
oTEm7vYcrZAbWnkNIGj35TO9eRapkt5gkHyKFCIjcphRoGHB5ZsXoXMYsfSHNpTPanFsmQMcDZHh
c/xbfryXUUrxVlg6ypONpdgkO5VeNDHxtQrJ30MlPnq/snS36KJRTvgLW7d6aPooRkSyPmHvFBJN
1TBh2aE8GojENBVGqd+o33G5jmYmqeh4dNw15rAS/ZqcKkJroIEW0MalY8qTw3JFxONyTfiKs1rU
YuNFXNsTixH8szy/Ht9YS3vWu8o4UpQURNLOK7iBM+5mC5lMnUpITsW6+NXQKhNKi4zDbTWmnZRg
7ni3mnHfqCWMm2iYWSgT9MWy1dpBBs2xqnGJUyZWeEWRv4tVerKkarE/ZLMs9/IiEhJBvgwgpTrX
Cq3jg7C0b3y5IyXn0Q4DLrEbbcT+Ut4tO3dahuf/nICtVmdj1X1GRCb4k/WCj/Hw2UpGuqvFAXl0
dTNP/MioBQSxHi58D/p9gl7KMaQ0Lv8bIFMc+DmDqidI2JsWCBCeZh5Auw7ONa26tRixRN+Kru5l
QLq9oO3EtLV84C7Ym1BZBz1NMe4MSaFGwK9LyGzUAZq5nt8ql9R1Vf+ThlpYPNZP0wsGbHTzgmfU
2n66/IIPLW8+T+bSZvL6ZIh6NxlrasWTEqkN5YBKJ57uwoHEvIL8R2qfh0Z0jGKxVhr1ATMMC0qK
plHHA0Lvz1NU+OpojAvjnhUMgnBtyuwRDZZmm422UFF4ZL6oM2p4y4JcTjkpVqvYQFsqwxy5dbb/
vb+vJhLm1RIv2S8KlaS9jmo2KZZuNwT4zxrupMixSqaGJG1ZP3Pkc7x6AfFq4VJrcmaFU0BliRej
CiU3g/w438uiajGkVcnrMXsuIWXmGiOh9+aDb6hrNz7nbyjrI2rhAdNoubddgCPpeXFLx89apeY4
+SGaYlahAv52xftbzqFaT4IRngKfd4luddo5Wzw4dh52EqhMvNZltl/ykPtmF8wP0TCQrmV0VdIX
RAqvk2enMZNdiOoloSM++IhcgGY0qCOJeNS86C9OUQ7kJF+/iMPHww9oV5KeOHboOzimCdxe/olf
ivgHiPAxqM0qwwEOeEBPwfA5apb65F7/kcpx84R2XMtd3WtL3G8BdSZrgt4fgJHL3vVnsFxS9IpL
pR/Ca6hjE4dOljvdq6A/nZZX9XfB5Wa57WeW3neiKYdawjkVBujtgIm4b4IGi7E+OtNUDrsnBIap
tApV9BE5ciB8ZSDN+0OlaSjIIwa7AO5W7RPazOg7KqX3I3rHePoFwuU3AdGb/pBXJu4gpJEA47wW
xtfsZTgL1UbzohRB2HgEv96qpRX04TnObdgr9InMHEvb7CHwsjJLfhRUB9y+F94iAKKYD2aRT3gb
RgkYLL1VBUUCQVkl7oxzoQWIO11S3mlZhgU/Bw3FxAtyMiJwKr4QQlSQEpiOSlqVyqrqsCsROlYO
fKv49YO2WWp7mkjce8lCt3hFKFi6Ja6BrTCPvmUHlzErdru/UfWYtQ4qziwS0IPcOrE36+lkvk/2
P/D+lipieoc0+nL4mo7nXg3IlfX+slTyguOP3D0vVNiYoXErSB93Q59/NbfYuaNIeZyfMS01P6Qf
R2EL/WR2uTUyQpgZds7wv2GuBHBNX2rCOsp20+Y9RRbO5amypKrP04T6eBxmXRivkKAY4Gknhs4z
ws12froUR0xViEwom4Zl/68cC+BIWvBuWaF9+9NVLyWNTaYtoCrqud7yCIFfaWTn8Ueb9H+tw1MX
rcziTxU916WQy5s1Ai4N49kcJSzlR2uQGGn2q5tRAkOIVlg/3O8/3lCPR6FTi543e5aMRCRWp4Z9
0nkVv5ba7qhmgY1cU2rdw9e2WqOPGUlK09Hv/jYgFBq0sYlwPRqAbfh/mOOZibMfourADPi90sT2
pohYZSbtE3Ps77yQbad8AW296phPHmA7ckn72SkqK+5VLH31qU90OSLMSEDshMIVi/lCmdRKRGsB
J/JGrUxtE74ELiG5qcsgJ+RvBmZWfj5+DucboxnEBhH/ZQgKQWi6Nh70LHh4HlNKFiO8O09gsoHL
P6h/nskMUjEIojPFdcJHPrJ+cD2nLf5kjrWzCUVSewmWZzx7EyITMlhjin6SMMD5g5Uh59RYlXcF
vIm7Rv/a85sBBXA2St/3YrfpUV0QwxGNucy17z7bhrJoD3OD+g1IH+/rZLj/0f5j8E3bArTeDwKg
OY2peZrKl9nKfbH9tXRWo9PC+u+pcoX9cA3UdA8V0pOiLzkyV5dcv9riCJKo/L5wpUROUaY7xT7t
bSbVUNMEhbf8HBx7/aYOfUP1AACqNhybjDA/avKaEvTmFw3F3Glq0RUsRyK/Mr4TPRWiJHP6HVFF
Dyw248A3J0Fe9+Rdgq4D1rnE80A0yL8K9eDNcY7MlxambLtG7dnJp7/n02QLKhqJZpyjvtMgMZ8f
lpk2nFJHhtGxUMsJJkHGtRI7JO0gQCes4sOiKnDlJ1SYvRxGYGtToeG4QL8hSaf4P+EX1JGXpRsd
CJqZ1bRrqFN3Ro4Qx0FgtV0WxvruIH2j7mvat7nIEfEJTAwSdUO3UfACnX/3klzBnVXwNb7kM/ix
1bNe+nhoMC03WSM8lbn3H16/D9dual0akE85A9MQ1BqihvWfN3UMlh+i+rvWDfcTHcr+vpGUtMk0
R/7haN3+XH6Ro7fOQ1MGbWVT16vW8lEZDgtuR84+J3dRJ2SNPIa7MvrlYiWBLgqg122mArMHn/ab
RdVK7mEdnNnFD5eomBf2uMLO5P5FYHFFl52Z2pZz6rAEPw5Ng1YJW8AK1kMwgrzl3vGw9B3efp/6
IGOnSTdPYCgSvvQ3ITbg1DD5ReBHkC8VAXv1XOM48o7yk2N+jYAt3vuCnNNBQK+pDBhpGQ5pbooa
b7dLKysifFXdHrpyErj3jna6jF16i2zv2AZEnbQoSDuNHMtR63w2cvtuaI/3LIRsQUjfyxYuE/wD
Yai54gpRgMrXaLXp1SZqFVASi6OVg0jOG9WKjIH+WMVLAgLoRviw1iCjWSAsEdK4R/4IJRS3katJ
XbObw6loLVNx8eq85FtegfvxokwgISBvyvWjax9yqHfNj3z/f5o+WbEv5bhhK7OkbExhDVvCdtTr
yVPFKaIWk5ED3qp283k8nAxr7Rca79aAbbffUKo6UwL85UTtqy9Lbf5vDAc4nzgjie2ZUmdmPFiZ
+3EIulYW05b+NP/BUAiVfJYDbhZ/Xt6FzQgLkqxXKTuTDfkhGTm/YDxHefKS4CrIWP7cuDx04Soc
trDeP/B9JmuvLRhfROyHqNHpMGSSVZLGLEo3Kge2ZpEzJXG9Yu40LKXFIgWNSvCl586H9DXQd/Ce
Liw3E49lr4fzVH32woAY5oFqnA024evuJ8853DaVEkEau7pIWGQVMlQ5uf3FboYDlHEAFIIaYtve
/3c+A+e49BZRLyw4mZN+nHECiQRDpVXyOJpKK3/xOT8Gc8C95/lvvaBIAGLjwaRfhQeVlSDSjlcX
s/UiFJQbhGscCbAywcznScOTk9Ell1VVbw76imF7ptXfp7jmXa9Ovuc9hwygs0OqRqsXqBIgU++4
RBXJfQaxHBEQxa8rqohWQjpEskd4MaBEI925NEa7QXXbi3wkFYLX0YLvlaM2gr3gF0NtnyapXF2W
G/7bmETrInEaLwDsKHVqVOxbuDy2CEoxED30zGI5rXz1E40qoVtNRMxGwpB16Z2cZcfHjw7YNhfW
llb4rLbyGxrr4Mnq5LsktgX0XggtUdfMNlyVv3IOVUPoFFRM4EPh8FP1wnAkxYhADgoqRZcue6Pt
2FpqsRNf3j2njYnlwTDja2r/RP6v/65KNh4wtyD1fBNE83SFgj5cfRrcMqd/qEB6kOJwmNUp/3y4
En2xdZiv/XfU+gIuZYO2wW1Oo0MndBbC/wnnDL1EXKI2z+BRmzCrAu69ivuaMA1M0dq5SpoqEhy0
CLBTdsA23taGR8QCQFgppaWgIQxezS/2nawXc0SbNir1oQ5GF6B/liDVJDljlcE/t+9hh+JjkM1Y
BhLrU37aUHUM5SlaNH1MGUIBMOk10uVfajYxYAgM4nP5RGuP41uArnxzw4j9klT2jf8Ofc2g/YLw
MGy+RQyAMEy4EAr3xgziqrixe+zoYWWmEHIEzi79E9JVKxfEOO3OK8tZL5acpyCxSSL8gt4pAz4r
bg4cBEoVrHJaJr9hmu/AJQxpS+gcTpiOGP/xDoul7vUWi2d9wuyC921gMt3hJB24Zo2pAmTvQdyq
AOUV+z7eq4DZMYmFYu7huMhZd88/AVRKiphg70qlP/mN4SWPFWkTlxW1q7pM1VouTgeajFoiZ4P1
0Po7EIap41PFZfQ1E7HXIh3JKIEwlix/bKB6MUTHYq0vzluXkh2Myg28pw9Y2rDe5CnQaF4iOaN9
cWXFAMaUI+1CXdLEcpHRhFgu/fQbNZ25nYOZZgQzCSUkCgwtOgsCv88hfpAf2mOY0RxHmlJO+uCz
vmMS1+Qn8efAvNrnv4gcJ13907op2DdfmCRjfKEp8zZlJ77KzuLUlAHd3J90Qf45DWgr1aJwLyw7
IjC2TNNfrvKmMjHSTmO8DI++wcqt3WK64m9P52/AoWrfCKWe2y+7VDl1tkRzYvtKW8hsPQPlZxNI
F23FcnX/35LbTk40pr5HVXUWbhR4KHwsv3oJ0tq9EBLZiRt3nFjLbCzmuqXeAaG2PER1Z4YbPZdf
1NgJEfD3f/nlIPM+bmjEd3izEIkXm+APZDec0uXhTr2S4Uy2hLXD3URLgOoMd1ymd3NmnbJbnz9R
AyEDAf5iVB00UwZjKSx5kHyCsDbTGUTnF+E+OShitkxMWUvH5+5z1qlgWdpfobr97bDW5ZraoIht
CVlC4n+h8M95qvlAYEJY6TolJmdUmOXDeQ7GQZ8NU35KkYUWXPHkwz8rPipS/ADgaFXMkpKpxxBo
3ZX65KguN5+9oluSyUXQF0NFPfe1eC3GEfrhD6tiZgp8I058wP2iILsBcSWp+hWhe7gGUhXHGhpa
TH630AT0nAaN1QSQO42qNn5Uwjf/1oRPP0jNz/9Ufp/F8+tioIpw10eakyYQPqYUP/sSBF7kUBE+
KbN8kycgnb0L8IW3BFY7q9xYR+GVbnb9YNxQ+Sk9C09ZORfhr1J42K8ueTp94z0NO1nVS4ECnFMQ
W4eRE5cVrxz9mB9TQ4U4rNhd/7hMy/3QtWQdqNW2U5kLbzGWnB7KNckogj1veVyB665gh7B+DpHX
cg4Sh7xe7sO2HCZK+ebWCPkRcezlCFoeymhNQw/cq5Sbwxe4s8B5gYgUIdb6WpEu9d0/AVSfgqus
RH9A61q4Bfos+UAg/s6lfFbaxFTcNR5ei7MExE3fhU97QnDC1ZmdT9kKLhoV42aNmyxQ47TsUtBU
N8uZ0qrbbuy5Ei2I3oCFF1UtJkb08wqduiDizDTeqTVCPF6ENy36PovnZhYEdU0OBoFnR23xucU/
QDeOPnYip6z3AJbac+CzgiiYlCUVcu+wkyJvOBg+ZysNJ/vZg1xjafWIaz/pUhv9MNyOV2ad7kqj
nkvXqgBITNTX6Uhy0Ly62eUu5SFm57iVvEYRBPhw7XBWSTSmnC0scaPFKI9JTe2YcG7ObK+mSWUN
a5oEMMK+d5Cn86phGcZ3MctDgfBRzfOQPlVjjHvEjmdPr/iIjuhmbzeuUsRfdUa9WmA2lRuTJTbj
azP0PajmglK7S76Gf7WLUwogcAgX9baElz6L5b9gWrIYI29iCvS2++FllPQ4zQ5pQjHxNBbMnNIq
QBt/SQD42GEceSQ6bycuQy9wIBRRmS+0ida/tAzxZQD1VJv2S+hyUw94QQlX9mK9jdyqonz94jGR
Sku+OIAlJnSonRzrgTjK9yJfjjkPAs51JglBF8qRRvz45BbekaRwA0ajP9rOfDqQW3U3jx7y5+k9
cabWboSOOiw6Y4P4KNtIUlxg0dKXKLFm+60BSgv/rxyxOgSaxaY0YV3yqgSq8Z/g5eb+VwJJV23z
MFzsTrwSVaIU+MCQFn8Ss6hMTWA0Pe8isU0Mr+YWPZQIYYD2cgzGS4kvlxui6O1Pi18uIQJ1kpKS
NaDdaXx+QqR7aoFd4gvQG+X3ZSGoDSm/cqXTSKfsW7Ncu4LaT9FIKZGqmwF9Q3lj1sr+NoeCZCIh
YbK49aZYoVCgncqGjuCBL12vM76jHdP1eFL3g7cDt5T0sLKJt/QQBnDpJseUiGAfkasENTDBHbH8
5JCm/apg8nH4xFSLiIiynwa6rTj4VXFtEEdcz+xrM+gmu0L/Ho+JjrSQNMO5hdqIdDtnmDTonex/
Lo/Ueya3HqM/L8g4Cfx7QUpPALsxK3GsEhskJu7lYi0B6Dwbw0P1fsLD4o9VacQ7OipNi5tqycR/
NdYDVtSZr632HWkqLbKmaSUUFiHiiqNmaW8bTotyYiN3Ur3HXuWUrWALfb4TUqIQrYmA7GTLDl7s
muTH6uklnAUIyGZdiVhQCguR5EvwGzHGx4BbMH0CjTSiKT39K7TXQh2QfGRNpbNNzblTBpN25s7F
9uw84/YMv54tR7FTH3T5NZBrInfWv0T2pn2MU2ry5/Py3wUy+OzKZ8KQ2VaD+/FnoFqAZAmVVfaH
U1wE7+7G++QiTk1xZ+2IC7YepwGr/DAnDJVI7fhf+r8WFQ8rCWv+8lo1a9uoMtqhKg6GN94L2r2H
9WWF3jRThfzxHqxxHhj1yqOxIv/zah+U3S6vknVLx2v0HS7WXC7B6y9H/3Dn9kehCyM/6Eh401vU
qstPsaXCYQg3vyvt5TRILqs4hFL7Mekk3O1mAcb385Z7jR+lr2ZeZeysH6QTl/DuT9idPkmZlZl3
cxjVIFqQ6sF2McQiGMKhRnLD3EM5PRV2qeiBNNRJoiuxUpnaID5sfaH/I/PnuBQiUSbqGq8Ik507
M7RQKgSeuZsV0F7kCK5pC3XAVhveeHb6b02sYhFe+0fV1B+KQL0kmqsa2O9v8XFV6kqnkrj1aAE7
0cVbEQAqqsiQbKL1hnZpM0LAq3xpA/HumHxV2T5MlD/CJI5dz2Qm8tEWOvDVq6KI0Rs8J6rjSyEV
sZwY3EihzPAiAYze8JyrzCbsvlVRS4qvEtDuMGgaMXXgx+2FdTL107ZSqAA9VLVvlOSdC1lKYgIl
MlXxXmfH4J5gfLgCpTChYfcBUHYJ+6UEn6Dd6nPzouh5pEF0yHMc1gtobrv9rpA0cIJXK1u++MVo
knTGRTwD5dkJ1obrBlul+IVGls2slCS3nv/MhIDm1JQ3qX3Of1Z2QU0khz6Mtx7U9gW3o1gkJYQ9
9BC6EOHFEIK6Bv0S6EG64ZugBAc4TW+vQfBBDMRPBZ+Sr0n8XDurI80kMGo1Pr7G6uGZvyQTMAni
c+9ewd6Y8R4AhxUnGS17czPzoHu/zcoYn9ul27Y48DYETG26UwhuQHIg7VVfDNjNjlz78yv38Q0N
fw/mIKKlBk5rXGOjwvgdtsYtAs1vVcUYG9HgjmFM+grSdZ2EmuwUydw0rMH3+agdPm2qMZe2CHAR
u3aHuNOfPl6mZyyycKX++f/DM2h3saP1BG772MoY92TvIxiUBzW+tV0TO594l+dWD3lzDqR+1ejP
bY/1UGKfOnMsH2Ics7cAPJNB3tVOnHbhXsC7gSZBYoZ8bDf3hTC9GWHFOKp+lMT1hE3M
`protect end_protected

