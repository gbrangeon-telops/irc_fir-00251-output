

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WH/1Hfau3yp/7ANrlzYJ6lp+xOi/gEnoXSHu7RquVCgxmSwM+u6NJ87pS5P1rM1REfM6bC/4VD/K
djLzpKr9YQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K9OQ7UQRJNNsqlJeKiLZja2cTpdn/7D08GuVLJ2Q7YwPyOa9sKS+3g/15LJ/yRa/zU+A98tod3ce
QlWEn4ue+HTvQflEH+MpavwOpNzd9uaRdRTecGrueadi0jZCWhKDECPBSOBftTcItmWjS+iuOrYA
UzNSV6gBgTESSUMmlbA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rfuGizF/z8gCeFD2+mr9MbjRWuTPDiFayAy9W9SH59KTv32ja3WRqyFVDNKefGFWmFgyXwscsdSc
S/STQk2WVtfaxUn47IIZV3HVYpgEROzZ8tdQyrDPMbi2HwmCfaz6YD5xdrfG9Tlx4ToidJJ8M9l4
XJdd32TWh7NYEzLxqVy6SlnR9JfF+0+Nf5C57mxaFcf8i5qJ+wGXhxEFyHFj5aPx81iijRBXdTZB
X7F/NtLKVCgLQvWL22LQZOJhyZVP7Cypy5OtaouwesfLnz7akydXxvJf1kqXrAdSNY4YWjxfZQKZ
dY2m3KiIO6F542kNq0ktevUOXRqWTgZJhPauRA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IUtntTnFOD14laEXhqBklNwiMVlWXctApP9259AAx8PFHjFAnJ8PvitVWk2w4ALBNs1tWO3QG+lc
7ANJMKcNRDw3DKgO31xMYxIed+W9fGmJO2Vhw+W2lfZUNPYCZDcGN5zCsW0hJkR6oPg9+0a7K7Sg
VTgdoWPi0vZlEf9gd0Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NobNPEAvOyayp1TtUWqLiTt1wnKf7VjSBi0esOl6kg2wXxaycO7UdL9j1KzK6yLaXpPqGWArWcdZ
OHZWjNgANQMvd87WyNjFR+DZMXSGqH3lTJ+rUOlsySu0gV6nE+CIBmIaadzXmtjlUXyV/oEoRCZr
rq22ZdRXEi/z57ExJp2QenIf48qX0mmYi5gFLdknqEc/38ewzEWm4uHsakTPzO6DKZ89VmneHDI0
7Rw0KBtgnhcNeggKkHBNrVAExbuEzB7b9xOHs8SicGFL9UTrJpF8NFV5zuKj6z6MHtvPDvJ2GC1W
BJO4/x680qEH+0G3sdhClIkA5Ln0j075tcfv5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73072)
`protect data_block
CTcRYliocX1Dgtc+x8/6N86XtjwyA0Lqv2bLko3LxMntwcc3QDecFmSEyRwYBni35VV0u79LYAkf
IIBGzYzSsN1MfVcXbYWpJPGWni7C47TyLfK8VoRGw9NmgNnUYNe96jOCuf1qyCmh94rwQFxD8JXH
gJ+VrTwmM489MJxDsiBU/7uewpm5DG2hJ8tV4j0tX6Bix8CNnG0gB6sbZs53zq0aMaYV0qiVITYY
eBqCPjePtpvj0hCT25kNvP3IOfKLtZ0J+1VdZzgZ/ps8KuyIZLsPUP834G2XAHvAeMpV7DUw0voL
hz2yEJM0NAUaKnaCFEIo7fqm9jUrqvNbX9C1Y2ew3PEPOMcpWm6vxrE4jR7zo0/Ed+9ugEryqXW5
7SmbWgC+8sO4l4qbj/iAI+nL9YmHuNJc53AqorW/+ZCTwlTfqrd/eE34t8XVuc4wYx7/B6rShj/c
KumatA2vpKCIYMHVMrI1Cnae4AEjHRyWw7YwXHk8jQPH6DMAoEZPXWCR1B855/nxh77klC37kHBy
kL+sOW7dM8tRM3eSkeCftmu8MRcQixGTwn6xme6UClzquws64FWCQ0P9wKKxo7ctJ04HmvK2srMK
FY/3hUz1G4q3FhPZZnnRFP8p1IzL5cLrRlfo0vDt+mvm08A6NfE5gu4NkpMHmZ48qcd9CKTSvKL+
/3geFSWksAG+F28xdr3A4Y/9dbgkbrQ6vrRpv+RlWkLv0aQpbDy4FvgPiabi0x9JlQByCCThHI8M
FAsnCXv3kMy4jjyPCEQ8nBoqrillkG7ug/tY9yKEHXtB0JYiNklnApxJufI4FKy3AXj17JuHRnpS
nsfUI0gRDUXarM02a7WD82Fw5OvebE23rKHYYeHUURCQOQee2lEgljL60Vju/7kHM/P1e8Sio0ri
3LVwtzn599YJrFpa2fESgceCFc586mssulKr1jDbWEg2tmqCe38aaOzSCjcLrd2+2XFuWiEgf5Rs
/+8CV+KdIJg4eUxpQou4TI8lwOSIz/z9QHyJks5tVnI/oaV9A8QREYn3AC8q0L1XheFaZOlRQKio
663ySW2k8H1Z3G0VkuIcbgzNsuP7DYVBP022WENrzbD2ViC49Vc6jCFupxsIp4sa0t7dbGIeA/TW
Neno+KSAebgQ3rDYRIQxQt+1p9Zpmiau+NxhFTo93bXoVJ4b7nTicj5+gx6RKDEL9yWbFBhyB0Hf
PwIhLlNDnuC7JqdBsvAbkumz15e8A8YpF7XkoSSsu4Y4Fcx7k3rOwXch4grBg4g+OGm6zDuj/9Yo
4Qlkf+2y90vyz2VAg4weoPNfiYRM6X83/7zEvlqMzyc/Gs5aX9xRX7fWewTGj3MqStHnufrubmxf
EfGUuR8Uyp7fvCR0AII217FQYzISoftyKnIKX6jxySsGOjnyNSMnP8rJWQc6JC2tg4sRm2zdQ7aJ
cde39SgyWdsyN17jUT7Jh6Kprq9Uiy4IiV76eSk11yGMybvOu2MS4/qv/bym+2krRhxSS5Cf1Gv6
HASnPSPdzusTnqyEhhC93v/hPWnff/yeb17d8T1HuhXKfFjVKLa0XlsjoO/ymaBtpP/Yfs6DqNBr
OWz2jZ3WS5GEsUI2Ozvli2Ltp+Qr4G5LnK9KR9/iOUfk5vyWqMLYPbnvbn7xBz783dLnrSSBPQj8
nQs+SRTftiaJVKa6TMVBORu0xNmB9s3AjKkPhycK/aN9PhPY7Gjxp5eA3LcJi8vbs4o6cv8XKk7d
TldRsmxRMAtI9aiN9p0kwy+xB6TWW2HXHzEy/eAywV8QzDDKTNPZhPoFEyQWzyORvUiZu1rDWoiX
Caa+hb/xqTbuGBIpJQi5COQAn1d1TFxgGopQHO04yn4kLpzsvGQaMtOX9ENRNFNVEhueoJIygz35
C/6rE7/HchOYBVBf0kl4zirLp3i4Ph6pb7Zh2FzG92nyrUi2GcKXbKoy3vcyDDn5gB3khNu0ZD95
J6GPUTcVLbFP9AxGMUkR9mfuqRa2lNLgeMDcqEbBrME9BzuGjQTISPnFj5ZVGUBP38Fd9duptq3c
UZK7qcQH4Phvb55WQazKfLgcWNQKa0LKFAeHE8WahRT6AP1otFRMuPMC/wjrgIPD5ZLWSqPuSaDn
b5KhDAr+WfjQB+Cgi8KyxwYsoVGIjajnMJE9mWnjpn/1XWe7TNV5CGUCbtsKodON60umbxnMeA/h
yd8w378Zrfeaz8sFMPGCkM1ayk1G4yDQrONZE6ktqMf7LSFY0pBCenA5zZc2X9UlaTkr9gRjMb3i
A1fBuA4YNNzKgsK2CCIZTD+0YsWq3UQklrUMM/SfS6AjYgfOfh3lnVusXUsLwsQaMqlihLIpAZGz
8gIcQQpiXhJdNf6rhCb+/UwE6SM/acon4Ug2rJcjtzi9lVhAoa28YtL4KyFjiD3KLMbxzcRiuOLA
WmLuVLSXOv9WvZMMOsowYrSmu76sL74HRiwZsKGBJLnRwkMHySkSP+GVP+h/tBcFdV+1R7WlBgaR
DYS2O9TgeTFTfVqe5k6MkEVF4EfL0ktacuNXKpwIVKsu9qTfa44Dl8qErBmQ86opfMCG/4gbgPIE
bm3986xaGXtApbZVsGJcm1nB9TsMCr1QtN+ryPFUBWLl/z5MDJ5TVPl28fjRYv64Qk/D2QvE3xNT
04eb/1RteyOIN8aVT6+CBXFaEWcIu2cTOWIoy6kP9ySxbv2HfgEiL33eL1wMdjAyXDcxwi2floN7
8bzJcygOGUFHIIsO42KoHJf1CLJntkZsQpyxb5GM3OW34t5E6Y+QLewpZ5EPr1LJHbrMeWy4YpuV
5AtA9JO2aEg3PvUVnaSvkeN9UqHY2xZAyiKZWWBTaCBrQhCgCQW0PPtWqadp/tnOspYtuVCf+rtf
prbkpnuJ3xC8fffs13QHBuQi0q52MJaJIXG6ITF9XNVXRSFWmgMTSBZ6JPI0BNsK3ULBfrsieBMt
e1G1yowJ6eJLzzvKUq9E6QoUfEAY90aK8o3DL6ctz4AhTTVpMQcW2knrGLRACCY7z2ydDaLoi8TC
kh7ojp61Jp+UrDZXGxPZCvJ+ntTFBicCvyxwpLhQMvkNnLoNpgL2RDwI8TvQ+OVVrI2VUp4ZkSDY
IrUC2A/U8J8QznzMzP01ISy4llcxRVb98nr3ytUa+Ztzoo+a14pSRxXnvq4fkovRyfckHlJvXkGB
rb9QAgVa7h6Nhl0/2yRSCbontXUaGyTkNEHzORiaW+t0gpzey3wTve/vMW2R68Rzbq1uYcBC0ODk
is3s7E1n37ItLEeNgzmm1V1f8QcpD2daZ3Bu28HtWdIbfrimBVfP1Ki14m5fw3mEXntu1BYHdBOZ
5da8/GRw+TEjknFh48qCISMQNnIcmanQhl7jw74o0rUKOExsUn00RwV+zDTN1MeRs5pvYr+lye3c
FDy/35ur/OuLpQQP0lhQt/5wyK312sXbYoB2Wz/nTos9t+zfgjeu5KrXHjmJWtnOu662V+Xch4Hg
oVbqBX5soelPMVT1K8QkBec/RD/HRZAzeBp60USwF1nkTp74+QcZ4e7WvkCV41FMi9DNoHTZTQGy
TUWKk4zbtEnB0/FTK7donpCsjFABGlRscBBqVxTpGI/nZ2W+vcCXZedeqmESR9POpooePzjtmdPI
sRunHoKYClmoLFPcYPRRfkOCCURe/d+vbxUNwEESBp86m8HMlcj7SdCFCMwBWwTJ7uMmX7dLBarZ
jyLGWq/dL1XFF68u7j6gPnCLjkIx5Nr/PItXJA0t/1VCwrR4j0cDLgog29N1E1ZHne0SxFFJs23D
LenXWFlrIC4LRh2CC//8PPjop7fOZpOFHE+D1hsae9iBIAk3Wr7ngW/xMvPinAgl+kFIwt3kjlUN
NKx0OXVCEOXNguL6O9gtYzWoNkaMF2+petRlObYQDqky6Alh398ANGMnS75dEX1++0Zr4z0BcO1X
1A0dtvWFikUmdJisPOLsxFn2mBVaFkjh9ynS10MCzLYqDGFFLWhmsxb2IXQICUrc9hszkQbPbMlf
5fbdeadDw+9HCjDgABAmg+F21z1XVFKcav5obw9xWvWktuw41rip20QkfOOIqTD5bK+XAq0LzYCM
0BT012eSzgmz4ReZRUHXRIXG9BFwGZwXbKmClnPDz9Nu86XE/nsclX2CWaddg/k3X5ivnB0XA2kE
rvu+f6MkTerGVF2jtQh5+ma3F7VsM/5TqHROVpkhKXkykaXiBBoqdoPip++VRw2jelhjsCWEk9ni
0AJUmfQdhjKyPFrnuCYqmf0KLWaEsaBAQLGs9fQsL19soJQPZ1huPo22+9oqf6vHfWyHThytMEeb
sOs5w0+SG+tFTaSl1npTOEq5kxh3mFyyxFwBLu93nv1Em/p2rEkpvqmNB5D8iOPkvce7Fg5gNPZT
0NshfKaiWKGSRdhQtyPVT5tkrO8aZykxEMIZR6QISGD5o3UR8YhK3bnU2xpXzZf/p/9T6o0DJCFX
FDWta8rCWMyZmFZdiLXYY6KBCGZsUc92KIXEJceqaj3E7bpta6uNX8xGB/onsZNUIk0qfciYl9QW
q6ra8BDu8G8To7wqjRci4Ylc6NLgOw2Ct48R97dl882aeuOSP/YO/FcR9+G+y1fo/APq6dmO3pBr
v4QmyW8v0HiKot9XnahVzwt7OZ0bIENYBaKayQ5vf3owhPLASQ+mf/ONG0a1cJR/Tcpey6MsfHZL
yUIyuw1pZBB4NxWEGitX4/Bo5s1qoMcH3Y4PRnvDSLkQgKOORtmpAiqNkEqIT3ckMBVbrLftaSOV
d7O1HidT/u6qgwyLRwT0b5NT3jZ9PuFd96iuc6dOhGsi0wDnmao2uXX6WZBRXL5kTHRiTQTna6KM
fOyhc//v+ZW8ZDVKbdsSJaLraMIOeXa2CTtBkSOstplkf0E7HdqgNRYul2RDfFExULTLizf3i4uq
APF9eiUr6xd0t2+HmwKd5HmhWUXpTLOVcbLzdKb9q7ZdsTDhN5syyTyX5Q44KFb4lfZ1sZURM6cP
pq1UY9ZcfZFMjW6tADtQR4kKD15jxWG4qJ8gyj7YRiruXfNK3j+ekD49qs+tTrh1KRpNAzY8X4PG
W5aEkWdiNMtER8kcxtEShHAmyVpE9jTfJXl0Z0+XH6jvwXQYyJbjp5EnBD0puTg7UKdI55ncCpnP
dAEo2JC/0Sev2YXoBiunq9J9mSDuMQezDa3zhdd4yHKjYvlkgxbhNzMSWzn2fl0Qe/ECpHJmn5OI
XS+Nkhsf1+H0SEANaFuZQOpOPNiRtHji/wZ2a7PE7xPtn9Y7fW6RObKmkU5UAb/3zIXclgcz3VW9
ZOdrTZfkfZSeL02RdVng6/MUcNIg5Yq0IySau+xD/+zhcacpfGRV+iVqbsTzJTi0cEilB2xEXFnM
8F/eE39QTNCh+HjMwuPqsVswdbZG2jMPbFNDpcHkMpGyU237b+1HE0PTEFOyNlQoutzJbH0x6DbI
KpnqKVvp+oWEkjobJcpUirXbMkT1ZtIcE9UJZwfnXfcM5xun5y9vmZVchr0p3T+vnhy7hjWm3MYo
IrBRM9IKoQePx2lHgIAKF38lOC4O35ZHemn3tkZcF4FFe8bIT8pEivuTd8tLW43tFCm4QaQA6TLa
2T8D/l1ZyT2B5+LCMFEYy2+s4Jh8aQkBgQMcvXyasK8wH8TdqiaW7aEh4gvSrJk7LOYqK6MDjSvO
TCpoJX8Xj7c2ZjCArfEsZD85iiOHL4GURP9oHkEC2K25LrU7IVMGeSEGwHYLq2ExL+YvLR6+2bQT
xy62e2bGlgztgSX/D1JPOEcsMEOB7QWIKX08MdsGH6WfSCza/eGReiOddFGoxsCGvmh9SYxx2gZ+
SE1fc2o5FJPv9wMrrTTepIUCc20HPLLHrZDUQdy4A2XTKzMdzEMQ6jjKeBJ5PSci51r+U+98RUFx
Omzzfh8lq1gKJGUUss9zNyr0bKfEZvyEHnvg7ZVR29et9yQ70BEJ4D6aEVf4htu5jOmdeMu9ajbC
oTawtDLyIGYddhmE/3hSok8HXN09siX4EYVfIm3zrNbL1hjcDK5yiu8faf5i/eSHu92g3EzNeeWo
8wGuNyrQzBjX2VZDbO9NpG/ckhgrlCVL9MAfplEihKP5tS0Ma6j2X+HgGNBUtyZfs6+HoYVuUtG+
+GGwXQqMsTkTmwa9sv/ovYOClhCoOp5gvClVS1P8U9cCchAn7/aNDbu1V8voMonx4skp7RH3a00M
Gbv5jk7QR0yW/n9qBvWf+FpiS+F7K6qp/ek4olU5isb4gl96avzwVPcmjKW76cIeIx9E+G95xhA0
TYOPhohP46GhXvySJaRdlFZrx8kJbaiC0kNPh2M8MQjxDpbwcMjOcdJ/FeYOF3v3hsnx0ukPTA70
CrwPTUYLTsLoJ2eub3tFqxteKBlSSQWFU1utVzGuNWFsHFs5zcqqchLGWCg7gC/v1GjI7FWXE+fN
PURPFovw+8NFaMz4drEK8km8Bv8bRcnMaNUh+oBf4ra/IJzL7YnxrXh/ebyP9cI+/rANBu+7ea2K
jnHk0ujvYmFqlgC/2Y2sizFaZ5T5q3lx/Vq0UhpEfUHqCOtNZDzhSirQ2S2U02BPzLLdJeup42GX
qCysaADjknbD5KTmF9Mv6dwzrLcuY8OvtpE8NJfnynXUaI2ItuxJemRKH/tvYL5CF5LR/2gnyr7c
zO3uIevR/Ro/F9o1rUI1XVZT3SkKn7hDHlkxHLnkEzW/TL1CphlX0UbnC1iXj+tWCO92RtiwMdQc
ZDQyaF8ggvXmeXPYbLgULK61rcYsxW5FoM6qNzOUAmfphAzU5qqRWyJ8873PB0o29prvSQ0DF+EO
q5VL3zjQ5FAvFy2B6WjzIkC7ikHTVzabmisJ74SEsZjbmGHNBnF0fjO+DoK+s5Z5X4c+uWWqihE0
AzYcrTBbyaQXuC1sMYbHWunMVCpqYdQg9zXNW0g2Qq1lqeQlmaBrvfWefnpL+LtpSyADdXXUVnZh
cCXMXwKb2EMtcrUO+QmdJIpbrqpMpBjK8p4N7Fv35InsHUSY+cfdna+DjF8JvUDH2+Pb8gJefv8/
Is67XE9hrmYPg+MES5N2eg4SQSPYkyyWE2ERyX3SO0wTEMrk/ZgxUogIYbttneTAMVPXXb6q/MdD
SoK7YdhazrFO6VDPhA2tAGTWi4umIF4Nk1Rzn8D8+YZ0EessLVPeSjAK2ql24ZKM6fTDNzq+VY8/
itdyOt5/zibMGUD59K0YXE5j/jg2YR18lHdRkf3U4k/MW6IXd/mjAEkO1xlHb5uaKRav/+m41e2r
V0nj8hQNgpgFiJv6esqO1J9OTVXTTOzLkcLfcg0hBOkZOd1Gr0t+qRiZsllk2p5v4iRSuqntCIHa
VfJO2KtXEjWZbYuRBUfoB0IsWRhZvGhUIXa5rdBYHyBBJ6TdQAZKyjunSpgQs08z7znC2vzOOx/c
//W+ikvhLR6ysx+Em9dT/sOA+LKIQ3EL28rlzj9LRqFB8YhDYafyPcI0lkCDZfErm+6AuyQCX9rs
Hg9NyXhuIaBzGQ/WbqgWXO1r207Tg7qUZ8deIhW3dmhmq5JKPiNFHxzRcZUowIu/6le380Sh0xfo
ESBm8P28crdk+DPp4kyt2lqdqK91lX7svWwzsQbyEWj26JhC6TXHlSDm/ZMhlpGYFIMJe1k66HMd
4ReZIjDcDVF/7kk/UslsriMcE54LyBwcrqr6tLONV6yLCrymyrKfKuNbbIE+jX7Xn/WwRRpWDdfb
/EZbbxnetPWNwqKxLfHpmq9W9cwsB6Zww5xvjJvgZHpLNoPaMEDIDlBIbxt3q74Myj2+FtBBU+N5
1g8G1aQxqJMlVyXQ5x9C7TEsB8AguJAZH6RBwIdTgKRECCG87N+n/+9kiC33kgE/c5KtMJiCHDqs
OBYUTmeQAN1Tyc53qVHHwFdqRYlNgwpSDgg0y4rj01kGfWppl5EvH29wKHZkO5QWQmSIWwdvVr9g
v0kguFyoTkIBQBenaYFzSB5Izu2sBjHnpmfUSqdBEcvIAP9jn+rE+BimWNVRPYfGKKT4UvqRbftw
LO1o4NKbhAXGYXbApmiSw6FKOdy/5uWPg0DLsVpNjeX58DlvbKw0rq6uKebiX+dl3jOc9ZrmqBZu
Lhd0ukMOXpr5mbSoBefbnVYyadTl+dUXNkbYQHKUpzVNdc5DmEMMW0QSD5jRL8PSMhpXHSV15TYX
CAKvJrSAfVWDaqtexRE11Wy71TpWYNgKQ8KU+HmL1UYn1nF1JWkkmOGDCPqxNwuS6nfnYr5MnWot
lh7nnrbwOTh5Xma1e8xCBRMv4UfMfRS19KZPe5nbJSDWS/cAFwTqz04MigZjdAek2dW0i7ez8GUN
X/8Jm+0fhIGpU6bVJEIaS/8DPXrWIOXVwa06tMRhPbIV0/clPkvH+7Mmb5cqdVyrkEW0LBFr89QH
lhkO8JpRwoDFtQdgAzOfE7s9+yVK7wTQAq3C2udTJhYz3Lbfxryhxmw3hoG31b1v3H5EqXFbswxu
1a3tyvwF3X9t4KZ21dE4r0srzjsNEk0enqL2/CRbBGoxZEhwZj/D6tPQWVmNP9MEo8mw/2dKunPK
iz5veG6HF6ClqyuaVRE5ntpN/RfiZfEU3lFohliU6k4V+yF37aPShXmOyccjEdSKvujtcBhc4G13
7X8NAf/um5yfklKgHurAPb2pXBqwdOl5vHmhLys5s4t1JvR8m4c0tDbgH1Y+EHmr/5FaVA679+NL
HOHPP/a26oUC/roxTr4YlCvGHI9sVM4hvO9w5mgFoaimoWVqnJ6pwf3e7oZvOVbp+XyVvDoxy5m+
hHxCuHtm5UmyIQRxadEVz84LDH4VjrXXg/uzr3bbp+V+lgKpBVWzKYyGK7Frckg3lUepa2jvYfMO
3nUkLA+o9YTafBQp3AVnJSOn5IBD4Ut7CHfrtrEAK15epiZr00bNG2gPHpacpQAwg6FzQ3MyoX0U
ttgo2hzdLW3rlEdQE11R8ui1kPSF481iwDgoq2pMtMKfbsRlVMEgdqYvZN+TQlTcTZd0lYam/3ay
OBjLgvVOHirW6pyfDH4swep61tj/ksNob3mpR9uBdWP20583/der0YslVKIbQIO+VTPcPyr2XYZk
RJJ9xmvWs9dKmmFQK0TF0q4J6UDClxANHioXIX7cNxgbpXOb8SEEPK/AptFtfhR73WKiLayktqN0
PuWDddbwchQW5aaJamyEQAzAp4Xc4khXQebFN0iFnWlhywIidiQZdz5OsILKzAk0BijzUdkZ8jzc
qkJCwQ5d7m/IZmMBAeIu5z/rFmKq87wOfljZWIyRUy5S2TcVNkkJX7sk6qvzjXj3W1DrN1HozqoT
ig70Hf8Wa8UTjSP+cGiegf0QJUDfDSk2Rxj9T06IldkOGeUt1Utawm4TFvAC2PLI2jrZfvrwTrzl
5/WZG9UztNlBQTE6PqJeqeEMRgTtE4iHsLwuDjF4uqzz+mfGtwuzgKOMIPgkPZ78g0XoBH/7h1y+
oghGrOroSEqK5VfjpGn6TSF5ktJkvG2TyU6xHAFh/HVH/OiyJ8GaRjAndYsq/VZAReiHPRhQEo12
KYqT+3EOWxTxMvad5NWGk/z+iZv0tau5CJaRCWeg9PtylixWtyl2f++jOUEN95QBK75Fcm9VdF2z
/Y2PGK+Tb4asLI74lzGB5hzq0cU2Mlb+ZOOSMjc6MCc1zuRuveOuj7f4ICPri6S1L3S5B3Rk2cg2
oo7C+bx3mJ8kbFskAVKCGJnypLzqUPOOggfoGTmhMBWWBiUd/e4tJRoQ8CxGKvn4Cd/hFZKsld+G
yUeOV2F+yjwck4vhqO81qcxJr403pEDM2kek7jmQamKoc6S7XIHAz8Ds6pgKLhGx5Aqlit+PZijl
i9v7hLhM/8QAiqzKoWTgf+AwZq2TS+IIXLvMl+nqBPA9KNDFuvTaYmdspX5gGuCJGc3WM030GuXv
Qt/0GWwQh5obC8E9V9+B60F8xjjS9tDeKuceBJBklwDOjF3GaezbU+SfRwvRh/M2V+zrGRP2dysV
gcGKPxnkjyc8LVJ2QT1aMy4Egev+9gNEhs56XfFEymH1FOP7qFE2NQIe0kON5y2d5t1TDoKxRaXg
yrwUdFk5+pVowNqO5uZA6lvKww77jLWQcgD1QI8Ucf0zxRQStEoBmidqYxaFskMbgnP0QsD4YzU6
Yj/hShRTmKL5kUZqYygUTktuZ0js6NXhedjZN7ZhENLMC8CTwzFW1UMCe4RLfJtMlG0wkLLbEtW4
RZR4quNOOYF8+vFU2KnXBZTijlicR4paCSZeAnWJawxgfgjhp41BwxoJmrEjXWXQt8sAb0q7mY6J
DkDemBBLFyyP7f+yAca+XoPFl5caLvn15NYWaldxIEZVUs4AsiqA538xmVetCc9Nri9wWbFPMd3c
lt3LLksrPFqj2kiBnp9TY8WaBqZyGtsIgXryJJWJqQSYYzMJDgUR44BGHldiiaRXN2ocHaGUN4mL
lh0UrSTRYsUu5z/XaK+44mpDt8DctOViCw49qu1zsrHnZftEgMoPAbp46yLUQPv6x1LqyU2DmAmp
diqAClZckmlkmxicbIFJrjAwbiZ80VPSY2eZgHKsxGKKHGXvk//X8HT4OedReyPtKrMFngxDrgxA
LHUwtCkyBJWkjJ+Ygm/pTBMTQKX6JUGYh+P3wRput+3i0yuDtDv2M0aOHqoAac8ujewwz57iuMtx
n1fuBG63SntH5rjSmKqbLuc9EyHaOjL3jWm/3OUfS2KEgItdJ4E5Iq//wf84dVZQDq6SyFfUr3HT
2YwHpeOZF7E0iEnP3vjlTrhaLSULHuOXwKitGisQDG5PJTnMe93DXHN20SieUMWBUf9UDuOzJ4tZ
HvDEggpmI+IzsOMkjO29EcFAAnV9H9GDFztkFRF8h641Uym/DzMb+2wmMX0nt8/sNqatPjjk5VxY
m5U23XIBUs0lt144PrmJaNXUOU6d8qx+fI7gE74iQ83gPnlQ2sgxft3jRPipUKFZP3dr1YxA0tSX
HWiUu3eVOOc3LEdd+Ao3NnogCjAMAzVL7o+83aU23HelY1fwdYBBPFNUcVxZDS+tEIrrXBDIzY1l
6Gyp1BjSuxA2xsMWlL+ZKxPSlUaq+z3NlXrWoVfA8VF5GUcBp4M0rUUHK3FuTHEuzTNhE2yNBLab
1H7kHQHqG0CjmaYp9TveNS8B6StN52Zg5g8hchQx/kOS6xwAzNVKKrGrwzR9xo2PHMbBXnbF4p1X
DDY8Fy0LvxZpeEQAVu3e/UuOx9giW2HkGf9hYJIoVPtt1GiftZ95Q70C/dB/susr0RDf39B2qyKX
onINUCjqbDq8aHu5W2f4CkuAqmfZRQWmBvGcZUkECVumu8PsIDwpyeBd1kLy8gU7wDHFhU4pn5Nk
o0F0xtiht0NaT/PWYyFRg+P0Nj7lDpxqcL++PpaQk6w1t9bSX9MQLhVUX1NWGqcRP9Ohd6DAtjsT
U3VDQDXjqxPcHLDPVSfIaYl9SU3+WY4WHNhQo5zKL6VLwofl5V6jNCnglWVRL73K1huqJRareE9p
60w+t7Bp0NrVa3+sQypkgcL9gxtcLNXDSXCFo8tRA7rPmJpvFoHU7e+2MaXhMyFku0u5SsQH7biC
w4367NmzRfU140YJ5BCabdhiHE9cNiQEBuxeq8SaeUluOqvu8IALAeAfeIuuN2USc3n+xGglsAhP
TiErRO+x5o6tHXeBvBz219KtQ7HdwnRq0HyEDpSK8wf4SK2v/XargBludPpDTbg4u0FB0rLpQVBo
DiEsc5ZHnGLExHixE0umM7l7FUx/1XOHmePW6vzn3fhRvRFu0CcHHFsKdpVtrEXNydIGRPsKSR9Q
uzh+eZRkS9sPkmAeVOlOCfCgUeU19JTCR7r1NNMtarrtDkwzk2gUIq6Rks8iZFP8a9fyJUWVJuFN
u0RoNX6uTM//qIoC4b/JjVz+rxzx/33RcUHD/roySf8vHoqbVYPnr9R+ICLXkMuo7a+98ezir7IC
aiZeBdBSXh5woGGAIZ8cfSyCKdFI57mzl+r8cwP284DfVmzvL0x0qxtR6KLFlThGPV388LrbhOhW
ZyfNipg8tZEpRUgWQog2vD/d+rvHhLhkH+dtysLcTMgtwKEd08yu6JbXPdLHZLpvN1ZDMD7Jr8VA
5lFOoz/NYdnM5gIaRcNa/H9kPwRjzfoN/JJPc2/ickmYUKCF5LDxmcHjenPmapnTtoLGbUl0VSZl
kJsZ9pP7zN+5sdYe8LCZ96I6Bb5mK1LHHpaIyhfKgMmF84RLWzb5xkVI/NQWZmDYCT08WxhpbzF/
wEIBBcQyF1/NfmvIj+ZRMgGZDMRkTC6Z0kHROOPF7QZ2GzhjDPs92Hg03cXzYTiIw8RXm4fRQUjm
fPrKk377UgI+PoJAZLzIiGCLLVynuA8qBkAV4Ec9Ywy8JCd/Zy/Yjr14aLWtprasyi/HHJ4eIKcy
PN3meupTB+BvHR0kLKjkWP0j0MVkmd4qiBghXrO9urBxNdINeJ3VWdixhyyS3PxZT4DgjI06DQk2
OTKj/QofH25XtRrJNUoDDSM6C43EgVd2NO7j8N/1uNnN4i2PQrpe8ILA7OTbDjSkMu7qFDP5BPye
iwd452MpoXwm3TGbQECemDNW6ndG6z6fVH6AJ/Fo7h+xrpzvi5P4VA9GUr3cbws9gHPkYImEu0HP
grrWckIZC68iFnbQuT2WMG5zBPn4efd/LG12KXckNJRrKEmwy7gbaqU2Wgy/ZJEUgDm0xE5kXs4j
wgBd1yyAHjid2cnm8t+Uv/Ac1zGiLp10Mp47XUd4dCTy4mBIEyi1ps6fvO6nNi6VYzjY4zgmDZkt
1cJoAB49rzbKi1g8hp62sCk+EyCCV1fFcbRCM4X8NNPz0yLj/sN4YkoYm6BgiOli61T8GGDGgCQ7
/3LUj4v4b1iJHBFk5p6PhLaxJmbGQHjP+TC4QcsuebIYS2FkwDRKo+KsvD0WxZowJ8UB7SMzn+0q
39x8rF2B5IzF0BHsdKxBr+5H+DGrWgTht9rBYgBEg0Sl99guUd7vwot2q3IZW6QpylQ23N+/KfYx
79hxoLAXOhPvHQo+YVkdQszASMPzLaD8IahbJWsMDMGLLXZ8iVijfPCGnEUAiinG8lGZl7rNukm2
hc6FyUEyJK44wzXzN1FkdsyFpM9M1ecxHqwxSAbK72cRwwMLLKLX4xr4qVV0+28kir+GdAcqbFms
zwKNFf8O5f2+7EOb8x4ZlBNkSnWDxSmCNBB6fvdjC5vXX3QHFd1Hqlryw5kFvVWGbppP6dIEL+es
pezAhgy3srBj68eZeyrWS7l+UNRkod3+QjDxh8DWNc05BKQ4i/88fkYaXhMmCT4h9lUA392R82SL
Ie0pH/zmYxr8icj4U/pDs02JamEAZILnTk8TJc3iUzN3vRpVosWBmC+rrRkmK6xmV1LLaGg6GtuR
UVhWaThLYnza8RsNB9pEMzReON1bh/1jY9IF2bXrv7416wjAhS+PNKOGESg4C7Ul0nA8HVnUOACO
3wGv26JikSZnWzSl4nhMRDo3LeOZ7/GLEHCOtmR1HGPw6fV947D/9+8POiU/I6KOM8YcTOl/z4OC
SLzMA8p5kOxgBDPJolUoh+79tLxvo17k03sbr6t3F4orT4xfa2dD6XT//fZR6m4mZh24AL6lmwnw
71A6mK6ZDCOYyHljtMj/mbgHlkrfXSy3FqNptxwdSYdHkZL9lNXElV9KLPGFPwlP+3dEOM3GNBKy
DbtYBAQTOniyEAiwVpLzvEdEMNg+l1Gu+QdQ5vYspKng6J/iQHD7aQlaBSjVXHyu7138rhNt67WL
JWZwS8oNpvRRO52PhtK4BqO8SxOp3RtX7FcvSUwcp7wWJSaV6STzxt9M5uRYKFX2fjBhDkRgxJYB
RpGVcxvY+MnzEh91naPPdHo0KqTgW74q9pW1nlqWgV8Ejj+6ZDzfz4Lpayd8CiOagQzzdIxXQndK
mWn0oQDFkALvBlg/snqrXf0BF+meRay2aqYT1h009s5Dc2jEbOxjOPXTtgIdSLV4w0gTlGy7HFb8
0ZeAsGsDNEA+4O7VJUIHvc3kYZAwBonucapcsm6OtdKy2j4RaqvrH7Pv50hReCRXo5JCtQdLD51X
wySgKJyq5aJ2duVW+X+84FV1vE0UT4UitX1TYxglhfapOMWNYDAm0u2+FDd/sqip3u4WJL0WI2GI
1G3fqoyXj3NMKgFerj5dTbV8N02aGhKKAHa1fTes0B99dvA+BDPrXC6ft7ChBVVVNiOEXEljHSGl
Y6XmxqCuodYnW1bSLzcw6cLpKQGkEkFXKZjpXxNfNrE0iG/tYhAYERldDqxVjs51i/uwK1FQyayX
AEH2BuRlwXESoaTah9PDgK37YPt4McJQHYv49kNQkjvs92ph8r7zCZRx4J9gC3R4FRJD17pD2Pj5
7ecSmAx7bXNclEkEClh2Z5kXjpDgMmpLmXhcPVDtezoHVAijivYtHZmhvZDOJH1zXNfUTiHGW83o
EH2o2gapgjs9AIPef9xlQMrEzBDOsDEzagRpBGN62mS+Qm9pxeRvwtbegddApuIasJtPweDap8go
SEoSbpnXLOsURFGygbxEfngGoRFyj25BYhLsI5s5A10X7U5cUosGqPRXZtx1Fp4wfsZmgK1EXmYq
pwAjEu42Pvqr+ue5E6wUySPY4123uMIcSFeYJOB+uSCPzJ4gIZ2AcUU9PqU/oTv4G/Vm/QuNP/bY
k0plYzFIT1g5BJXRi5hT0vrgCUsj/IaCzF8xh/ioyAq2FKtiMDFpsSPtMojya1jngU6mf+X8wfg5
wIBi3DsRzTAd8oKk5mkMRJ0tW+rbZePtOUXXxv7upnI0wcOMDSc/87WtNDbN+WMZ4bzy/Bo5DIrk
23f9in22SH9JgkwFo8JeqHFOAQtrotuR1tenxOwikGl92vZjUdjpQoAFZfQ3s76q37bvQRiIQutf
HBXe6voxoWeaLZOVHwYBZx5e5SJP43XkRme/xrNt901qbcp6lynKK4ptdRuj5HR7cgPw7VLid8vm
pbl/4v1zZPEl2Y2RiSt9gDeWs0AcmDeW3nNxtulWpxvMMKmECiWRfKjVhzgx/wWr5cN9u8udqwd1
GGDSH2iTEY5P9XbIBBWtkwsrdSu+j3kU3mmrjnbGjjrA4VPiO0f0WCz4eaYiNtt1ocFmKOgRhdCO
BLQwiWsIkFAoxZzbdopwe1aB/7Dqj8jvYNGgio26NXiITCCWaZ5te/9YTMxvh04tl9TzDodsAd/o
fp5Oh3fIw3PMKmAjjApK2fi3ALYttTkwtFbSnVKHeBfoLgE+kxlW/FGzTzkIy+BIPpK3OMp8uefH
2+p601ThO5HTGGUQI6ouKm/HZo5/RfheOFIY0aCg5Rt3jTK0Ex0BfOAGbgRv2kfgBC4pmm5XFZ1t
NK3Vw9zjH4Zm37VVe7cwjjvOS9XK31aIiIjQD5lk7enkXHkXumF+PspyH4ERAWAkC0uKmfbYqpWk
Nm2OBr7MTgLIILdY8RK6c7w2GyxlgIQZDO6HJ4d/rXE6VzHHoCYvDqhbK7ohRYfh+7v+jOFYfoaZ
ORns1fjx28HWZmLNiT6qn4hvte2qk//TjZfqb8xtD5Xqnc4iSnGXVWahSqkjsqtqVreX3BLqyrar
DNwcCtu33ZCXAOnNWu+UHFVj7Xx3yXs7TETBxJQuvOenj/56dVTtkfvFZO2jTJmH4AaEblAXUeP8
HtjSzLA8+EvTdwnC+ZoGSNs8A8Pc6palN1nlvEE/XOfH/I1WujskVUtpETuNI3zMVh+QT3ql/k+O
dm8CMa9Q/LGdhqwQfvZNrVtV/itTEWHmljdlGfcGUi+1EddqRkoeEJKQu8ceRFvRoDcqeIxCG9K/
d7fmW1R7c75sbRBYu64EafMe8A2MhkWWmoX8RN54O25s90m0ES5HNAQJfilE/3c1HbtNJAc7icvh
i92et42vPXRXSb949kHmcx69TbaSJ4dIlmqhmj8LPTIbrdUJKfgyTuu0shYJMlePqNRkCyOYnDAT
Is0ZBFRczFmidmWZpUtUOaBPcmqTKUXQB/vB924vxMQgV5/l5/lKA71xf20YbOv0rFz+HGQiiw81
qxcOaN2H6vQaGoOSMqk7/DrfMuelQd1Ls/BJz2nGgDQlhkArnUBDTqrzMOizaE4xw6NMeRXlR1F3
LgTQEDAmbd+ZHOaLDuKRgE/OKsXjpxv/cdyGiL4SV4nUHaFmCB0KX0364Q3rYBlbMC0Kqx31bJE3
AcqhBAmL/Kt3jMWMPaqj5J484YLW2TXCpQ8eoLxkeQWQmJS7immNTxMU1qUeZQ/4lXv0aMbHHcy5
CIydZ8xT+cPLhiZPRd0abyls0WRKoxiBbU0Outgc8CBRJqSbeJVrr0MtW+RZRre5mWc6EcbJ4wV2
tx7P8xUpsTtO3ZhsMw++KrESwwKDhNGahIU/x+MHwBkwsuomvcf0UxMyKD8xKQWEaFlgDQTII/gU
+snB7cfRH8zoKpeurDCh6ZwGg+FjfdccTnsF3G30g3pu8vSGnbcvrpMGRP27CGRJyVKDjkX+gFYY
yvatusNRGCxvYIMO0ROYRTXHnSdEI3jczL4oBFUWgU1eYLxkOCKZXhX45dAcJk1dpgQZKM1BruPl
Sh5bKkc2tJjXkIzVT3ReZYvi3YjzwHVCLT4icuxKbEBZtzSd2ci5j+facSkvHBRKmLw6gT1rqu14
KVP5KcF3hGY+8blQIPGyQLaL0UmBeihFUIAdkmwCYZL6814FxKZtsCERm8AkyGtxclhX+5PHbEA0
5exVFN3TUoB9BRQyNy0nueyN+cPaNdEHVJpe+uchE3gSR/S7ZEJjsfERW2tT+Et/r591rm4leyyb
VBb+eAEc1p8HEJiSf2/fxeHF5WTTKppUFSp6TIADTZueggLIGpdCm85+yJknOvWdoqdW1g+bxiRy
6yBcVPzFL6HbEE0AzQRrc+nf/TD03+wx2VT3JmLjYmIN6nPhmrvQ89mriaZ9HmrBavt1z0NUUOvb
+7SUctuPc3JD9xyRVkq1uD4f45e4uq0N+we+zaa+e2w/apbPpTTRGqPJYqUMER2wNWVuuE2zZnAG
jbxHD6bSmny/dEoImDMFiJRPMDkUii+j9nclPTMUEPkLUIoA0A6JFDeq+eg/oHK3WC2ZWOJDOg18
LtsMXoHqZ/qTcL20NUyAGvOyQZo3rlQxfvWDCheb4rJwOh4Q5YqPp2ztXRh+AD7sC3HURzuUBAOe
KVHQK22JdewxQL+Pet08zpMXgKYToJNXWifirHE9G1aIlcwT4KN/7PJq6iuUCu9iHh48vT8bl8CH
G8tBwQZNt3TluPSq9kUrQkUfEofKBY2dLVjX+6f3scALPytTsXnz456g5MukP2dm3JMVq2Z6pT3M
x6rd2zHpOXKS4eL8/XL/Y2R7MFvhlbMRyHCSegQf3c4EzFGfCBrBUz3+DRNqIH7S/Nj4Tcc6iPey
u7zsHdEs8LzhJtlmu0JDXW7OhDXy2+q/txPf9Gfqf9NPSKNJO0VDHlS9c0NJafg18/XDPM8DkRLJ
uIqsQjLOUyaenS0AkQd0ywyWbFqswv75ii7KWjkTGfczoeDfS8i5oR8tvUXphRDtRkK77X+F03p3
F+4R1vpyYRBwe5GVSChiQQ55xUfDfrX613YtUE/EMNM3cySkYpKA7umKekYTcRf0UtBQBIap0X+H
nCpZHcxhrvSp3HutRyLve9e3jOuiWcV2cFAGANoIjJWR2Z/s4j0XL2Bw+At2JTwMY8AsO8QbNvtM
kT4FWcSGvqS6wTxaPKBnWN3gsaztcv0nO5pMlWItLl+7bDvfBfX+h6CxpajDNV07w8yoz6bsDAg+
qbKsLeuhD5IXASGIppCs7+yIalbnDdMqTznwpp+XDBL2/lko30VsqrXhLQMA1EKEYzVgkCqR+ffS
usrL08t+xgoneC/aFiKdTArRjYgZqSrunECOA4mVqVZHyWPGR8hAApG3ehTafFiT/DH8wyDFT3kQ
KFWCOza5IXWkmkk3wLhKVYg0fjUgi9ar9rUFY8q+gmJjB2uJmZHhbZOW9fw3uqNK+m5nAArA2QGw
WXbSE9NBo5kcEnuSyFl3cpm+WkL9jqGXykfasxx9XVIcOko90ZrlH90s21m81vfF+SYq+W4qlKXm
3JxZxofJCrcZiNr6COI2rkI/C1QXsr8sz4fbjKiRvsC1X/ns6JF76pk8O0JqkAL/JkPtgR6wC36R
UnCaPYXNoMjkMNy6VeAKVdAQuZMp6qHaMKSk0pMufOsDEDSSI8937JB8bKt0i583OUy5wAa7JoIB
D3wkavSj2x/eMRHJ5joim6E+F6Va8j6A3P7BeQur1NEZx8WoumJc4CVYUypQHW8KEoqmbpj5GXz0
J440OU3swTnZWEhNANR63/Q9m6IFq+FxSAX9qjPoeWYnU6xG+gqKoxinpl0gPnnSEANGlHggE5WT
zHHQeYckdDUEaMCp3m0ksgt8u53+BIftHWZHjPkGUTUCgSjzo81IRZyBQVSgx7aRZNdp+bfev5wj
5wn7eZipMQyxuTW2d3c4NipsXmzOdE74CnIpJtQJaCRV38QAA2rzTpEEPynIUUxjbiV6MWU73jxI
e2vWSJvyraw0iTbDs21/cT3M/STPSaMj0GXKkx3YsgUtwN25CpCBtbH4pLYPyIGA2lGQ2znPiZI9
sLXSAVFMclmHuyNw1fZ+daGUNv17uApmNI4waDdAjFgJggkj/Mih7tPS3cyKJmDZQUHRfwDO6wxd
Wb+6LUZuS3uSj8vJdSWpqXymJsa9gxUJFeI9aas6CtwUHBFi0RcHI3xEUrBs39dPeVfmfDGFrhsi
YcJmxaWO6td64MU6qg42AJQsGv9Ds0NLtK6u6JrRRmbSqRyP2O3lRFfjbSJNo0boYnXFxz/VCq9B
e+pebQ3MD54m4BO5EuO+tTqczAWKMC9E8i6q71fItjw0+B0/HbpJJsaAp2AGbp9uFgOtAk6x3qNr
YlY8C77bTvW4JZGC9+NhFw6smJ03ZJRuky1Ob2uGG8B2LePD1FVg2hibS/Xqere3JKnYI8+xChNT
K9Spn5mDWdJ3T2OlHWcXwkCJ/MXe5+jBmSAGcXI8fVlO4X5JiDmjJczJiZCfS7BvQGRiFWQwWeu/
3Ip7sAR19lzLL5U44YkonWqVzuAZUUjBMtKEFBtda9hRk13OpzE0DD8tjf4NFLL+zzpomv+Nl0LY
xxHtGzYWt4QFIrWGOWPk8z4INc9PxZCwJtH/MpaF3QKUlqxDmvjvf35QLCswkB+40CDorEAnidkS
o2LvWM56yTrf3RPf3Tk+wIxP01AxYqayZ1Av9Npopt6IqcU5lrwRUehMoDxdzdEO1H9FQzYz0zuJ
ROcp3uHC7oUrTrHpe19EMLx2NnDQ+w/ydg3k6pEPcO4VhZlaPf1jWV+Nzdna6/TizcZbPoqQ8B7T
jbwlRoux5nLxkTKDxPtyglhOQvgCvVM70iRh0nduDOLRN2IsJBjWaZitftbpOqVFMXil6iiOzba3
/SIxjd/zVkhKGtudH84nGnFtdP4AOx6a/ubWAxUB5ibmO3/u5EIZfYlWQtsH9a7S1TkHHhlNoLNu
A/ddDaNYYCXEmp/px+juHhMbglsoKWAqKdTvCfPeHaQkv6BrfIJrSsFH2/HFsqi3qb2OazDtFj0H
2zsD1Vy/LZym05lHEvSfUDZNFr6P2Qz9+8+zrEb9aHzACnNCDkw4ssnJRAUFei4hoTfh1cE5V0Ck
SzIk6nW3/xtygteKgt1yh/zqOQhDV9rSsH5KdlgU/RKzTEb1U0TT6iTqmB8ECNMM4KxEQeqch3h0
m37rMCJC72YwX5uCI0v6cLFXKHaXF+KMsA/qF82oFkOYXY1JtDIo49DN3qtE2qsn5b4SzWqEgmB4
qVZ5FqRedp5OrOMzXmOV6WfeNvMhuVgpRibeuux/NT00OrOrgV0yC0qKeSvrviMG6iKqdi/P1sKM
N9TlvUBWChBthPGABGNVRTU+GpFywu0wmupsPJtnJOO86za5tLbgN0ikIkm8lGD+qDZ5UsmCi69s
+XDC2Zn7Z5/xE/NDuKFMkCdLCz4cC99lJCrAJXfPj9YN9Kw/PZSSLSyqlv7IlnkHWIxemZD5JsGS
X+kqThxIq8fRSq+Wwv0sYybKcrjZjhIerNt/pT3W5rRzgQi2x0G0QG0BGfX/16vDRnLyufpzvlFs
Mw7D161tYz3T60j6VvY1KhQG+nD7gHqEb3Wclg2Kcuoszf6BCA/XIef7h2NofEbofUI6tJ0+Dsh1
BTON+tBobal5cAWAPy5BIsZli1E/CYsONbfnpMvVKDuQnzkBCkKibzNvagPNur6IVI+kt8ij+sJs
Dm4CuX3jTA5XIFLajeiJxEcsW+jiXWyzLuUiWcRERtpQubuQ0DezMfo0uODr5/xjqyxGzMItjkvA
a71/++PCW8Ajq4HNLIbC27d6os0CQz6aC6B72P99UdrLVKWCFKskFfvmF52z5D9vS+cjylRPFlN/
QpIcz73GyX+5osA/s0LGO4kaqc1BY6XPDPQSPLPgVzJaMwm756c4McFMbIM3i4txhSJ/O//geVvd
xNFQKJr1LLTbD3kPQ0bO5hs9+IW9JBaDEpUjxIsn9lT4HcfsXuT9QstAq/lnghM69CnuFLCJZ1CJ
d7xQa8yE2YnlkECtbI6exkZcv/lPGNjvNXq4WWVvfVy9fFg0JVcOPKixxJhYpDBYtmKLr/oijvae
EY6iYjRdtq+Gfco99vjOuqkACPoWltdAhCIYTcuXEwmG0Z+x2lId84kfZJfuKCWU2HuTAGUrEw6t
hGTvzJYPGaFKjeGUAUj09I4Q99UHMe6eo7XFTorIyjFWM322LzWx7IEu8X2wK6AsTUDoTa4dbduZ
qLl7CmV1aHhGgv097kPeQCqvME+lpbumQQ6iHoXQpnC0cTno+ZZ3QcZL5AuyYridlPtbc7BqmcUG
wYMd7lJtnOIbtIF07dTAfPAIf52ZaC1vATDoAZE/9GcYQq+xSBn4dx7be2VD6srwGccJSw9613bF
qA+03Sp+k9+aH/YwECsRugp3x3R8iEkHrRdymkW1FDf9rt8ABUxeRkIaN2+kup3Dh17SSK/N3Hl2
hn2/VHROIaFy/dNGJrUMBpv3Wy7BS+yW+rOGqNNo+qOY5szn45lIYWndzrlXHyjasrMfMpWpQZX/
4B7Zy4/PdHTrQPRNzKjSL2DApStpFLwbAy1y+iraktNqZFzM9UdM41cauoqnhyCaR121XGeTkIwT
/5APA9JaUMdUke2SYsqzxclqi7dkDiokJppTp7QGYDYUhUpIYR8GWQ/oc7TAq33J6NFA3O3n5yAX
OR0P1oskbUMgxc9VqhY5xFmL1hWSl5LEhrPa+60PkQuRXkpD9cjyKd3Bq9P2wQF+BUtJ3XH3Xumn
tXHa6AW5gcW7I9Gafk9F7IvHSuhQAKDEWyIp29Zf9WZsbwXuzJ0qi/YXx9EfoaAgLfCxVSAHahlV
y1pxxWcZF2uyfkWER8a3KNDO4LuewkMoIAejnqkSuyJr1dVVy7L/fFkZ9NWMaEW0jwNSEWNVVEjz
0tGkRojmCKGpLEmgUdcil+u9xfOEJwk9i9Nd9T7hODQa8CPE0NP04aely+4gpUMgIYiVSwGLzk3Y
Yab/DkGadzNdI87SL7ILfmKDV/W54oX8xIV5IXp+38eDzfU+BbHC2jYZ9Mtyosaj/oOnRiC5k/Aq
c/lpayQlUh+jEt0YuvmUxCd1xFoXCnmR7YnT/nTcmsIxCABPMFRtpkfmLgP7QTR540QcgWTgktji
4KE8U0A0KLt3zFBpRo8CU/jaNgQ8Xvzp2mcvZ/XoC5O1naqAIq1dVQecOoc2u/dEX8Acw9inlQnV
Gw4FrwL8ASPee8ZEmH4dKuUtkvGN4tPofafcbvSOFc4kw85QWUNJB0xLlWoyV/p+u9c7739CvQYS
fsdWI/V4it1KtU7NaxUL8FkAMY44q9FsQVqF9qVBlF88AP7MBPks+ilGjsJRJie+eP/VPQZV8ChV
Jyg1PgqU7Nn8WI/vNn6bBB6E2Ta9z8BLpXH/grTAl6mrOhFy0GSi8Il+YycKqwE1NO7A0LItXWvp
Q6SijCz8WEwgm4Az3pRZzMX7/cHDpA1cDmsdQ6Ve7GuykfPhPugouiyPfh2fh8EItBZ6fBpTm2fX
UWtQjzuqc15fhTp9u+FG2s/chaAuZ57aj0RkCvk3OFQsqP3Zhft0cO/G2GhK0RQEGK3Ux1ZJLS8D
nOeQXUMrbaYVjS4HlfBiKMBcywo0ymS0wGWWOpTpVd6OK1tpro5gMEJCzEQwg3ERtHPdiTvMRMIi
egtRKXEL3jal6mzisaAF2A1vnvPpzzQd6n8Kj9uFWZkDoFk5T4y5jVVQ0048o1GmQuBYorczyHjl
NLIu+QEIu4nfCBE+Ng15PPnmmjOLYTrNyjpzhtK2yZ2QwZWcgLc+DMU9tnpdYKtgvmEv7rRrBxOH
llv5MT7XTDu4Tbzz3DYDML2zd1Mbke7J55xZHFxXUA4/An1UB5nz9b5pMEigiURaGo7Cq74txoh4
3i4pt5FRop1h5Cpm+/1VGgEAI4vg/34moEHhbKRyZgSvsIPNpFBjWdduQ2NXq/IQnK4YsAG8DhOR
KYu6PiA1uiAnf20gBelufyMJpfELXpMZQbugZLaSjXKNjhsBxdQEQGDergCv+mlX3g6reabEt6yp
54hGS/IW0txlNDoF8/IuFmzIQWrBcrsahPIMaXEaN2J1p7+5kN5Tc6DZ38DPbTIUFjY45+xdp+Tb
Hu5wE3TWHpQG3W7mZ+Lexbccbk8wMhZy2DnPFhBZLUTXmooiSgwWEbOlTEnEOILnbuOGpJociD9C
IMiY6ax5XOkg6xGDX+Ji2SOvQRyVtvF0xqYZLekyC4nfSvS1DA9DzmnikM//Tzw7GOQe0No/jvdD
36hv3kzoPMRqSoikmU85vJbYOtO3nnYEuVahDzZ6C8iVcjCCxsv6tAAcxurqtzdWOGr9jBI6gzQg
B4rfVowNodhpo5oRFzcp1vlVSWe5PrC57ZHO6O6QaRvvjV13ICdrs3iFpzVi4AASLtuMP9C1C76K
QfK1Mhl7piYzaMArhpgqEz9ckx6UL0Cd6q33gpDxWV3YcY/EzJt5BkFPjm9dWtv3JlC7dgspjvTb
UPCpBG71rUp4Lq8D+qFprU3ge3a5Yp/Va4LMuW9QpFZnH2AqvYkBvqHfiay8kXERDz2TikmVV5+z
3YZd4nfc+6fvuWARViOFqQF+nast54LqtLAdEpjTh5OWtMryLJFQWCz+N33LyEH3mPtwYC2Y+ov1
dvlaorOQagMH2n1AMxR4ZRgVWiqmCpGYZr5X08ocX/sDuKAYxOvfuFLKl0U2BWNVXCn1NTWvsIma
44AjDkDoGLQTnITP5qsxevhOQc9pI7g3hDP7K4IRxPko39c7SIeY/2uAdsMRgdy8oSF3V8uZ34Fq
u7gxSJTRSy7KvGa5k77X/SaUoPkJUWBGLpqHftPf7VmZx23QML2Spa9E90mIBSQ2VYsp2EF10YZ0
kdnaUWJP2XxpOldTNyABhq4quoFmKYtbWMAbD/hBv24vxGigG6XGQkx0+YavmtRZ+GykBzv51uAb
q63cWlNBBC4zBURpCwjxY1CzGXuy1LMWRmfjTOfIx+LF2tFGes0vooXPRr3VEZWienwF7J3yg5Wc
5sQv77xTa5SSqCM4eg+uWT8AuuTDgqxj8GmsWQoRvrOXPR1A8cxGQj3fcdDPV8njWv7FJ9cH1DMb
8sPJp5saSNFTQbYFRS7OYhgu92U+Pmq679rpD6ncD7BfEXnUQrVsOmuKxNtOaUBdyQTVQ51/djRw
ZkDry15PWr/sajj/c8xIvIEe5JOKAAGbxs3VPkVSG2wQtPJq8lNDLcKiYpxmRCdDAYylYoHkXnT2
CL4jC46v/VyCX2lbgedgt8AFjzcVQcfi2N78oBsRuyo1Xqhup6rFd1Ta2MrKGn7CM5FrOnw/LWxZ
2xpkBRQLot4UIXlEJsjo3v6TWZO9AQ/dr07YNP7ay6bab23ur9UFi8e+HmQQcCwjRKOBxQSXjJNe
imgeN/r/8gpcNkqyoQSr2kM3Juy/rkP3tHo+9LPBobDANdKHgcJW/yUQ/o5RNwylUDOy7yUZQdHK
q8RVHiUhF5zQ6BgGU6lGBX0jeHMGT8AEKsZLWGuAbxLfO6PnDVBWd6HnymSlCCgEQhgWrs+nb9Hy
Y/DYvp7cZ74zEAF7SoP498OIamiA9DfYVQbo/rrNkbljIYf4+Hdnu9e5boT8lmmPa6F1vgYAoIzl
e/qTg/5Nn0AzJreAtUSPI8rMidz2CVWkrpiaXCcL8EfoHS12BPiO0vUOrdu5YaeT33pDg3Ru3bOz
+lFbhG35n4RU/xWPCI7SK3lJPkVMmwIgvgQ6OP01XZYoN5JRRvTh5FrqjqLgjLBijotUgMPj42ER
YLIlWsRVNKmoBwQufaJocolKESaQwDiLKD8JpDi4Fp7zBpwTubed3u99YvWxDtgYycpN/Te/xTSm
LYeJJB1Q1Wu+cXbF3SJCE5xR7/gflbLUWWTzRHtiKde5FwIbbLaJJBvC6vQFUpLFgN4wShHd5CUO
LeRuDuV7EIGT50TZ4hyaKWka5q++7bN72yyhgT9cBC+RmjwxDBnvYz603JqDdELWXIdVbtsN3TGc
VG0Ds5QyU+xpVZwlYfcDE0a58CMaykCR9iPBUP5Dmox9CVE80QZ06FpG/nXeQI1Tj1WRdWAyXlXH
bBFgOqKAm+iK7OIjSG0J6me1V/XdepcZl/Y3ow+n9iCcvNhLh/BQSjygJsZpKC6ZWTA17SomgKIU
+QdODwJRIlaE2qcWhd1LDriSDB6LKIj+vkRCDQJzbiEgSMSiL8ONXfpLLmH1aYNyfPm1fbZTQVh2
rHPslOMuIcWu0jQWitKGmY+SdsyYRRrDShb5gv2yAYQSXb7aj7U2Be26eaIIyM/RioJPT52UmoKl
G+hxO7rSgG5kmBpOWmEuSPUVC//sKVZbNFso28aS226IINm87SLlwo6/KCtxWyxea1AtY6UbKG2L
Nbe/dYYduot0V4O/R5kYsjRHnn6w1ZJe8Dp4hxKGbQ7kRFQbOEnv/CSa+NVX/lhLq8WN9yANX961
q9olnH2jhV5YGt0KkarPbRN0lFLo/Lh9G9PMkR6klt+PBhrKtJYx0cPrseNrWrcHtt7HN5kxkXtl
nk8EsecimdIxYeXQlvsCmbEHivud7YEibxkEb9TRB3LXmGOLTbJNvM/jgyod50wdvd8+gAyXZzMU
PjYMYanMZklzRsT7/vlwMEx/cbeUY9nsBHRvTm6zzHAYA7x1YZAAc6VUjHntZoLAiFJm3WUpkCwu
OytGem5GZraMo2giXcjXTGJAxHN+nOh4+6wiJnAwmw7Nm+vaQ2krsbIvQoVkU9XnGmctVM6lcjHB
z5dt8fSlNQVEMqacBWFSp7ChSHdS1+LyK/GZUzGFmNhd/H8N996wU7diLtTpmtHpNtSVcho1WbYA
GlPQaYIf3pUEARxQsa8f5wbdXTc3k/qoREViIaSPbw4TPDlfkpafQxG6s5WvA0tZiuiIo3oH6kzJ
Jhvwmi5IDPuOpA+SzcJq3abQkUYENUZQNE99hJ6Bm6z8Wrx3GVRTF3d1aLGXnsobxT6AWmfHX2Xl
AArXwILrrbdLS8Hvo58hjfG46DlFaKQW6OnVyg+e2Y0MQFJyUo6Z4dQsFLsL5pVG0qPeL0276M93
nIUGBwlMRI4iSE7yFd6mRzmUIx61DmVRrW7HBmM4OZXZa6AcqqY8Inv+QH+z10diYtdjxpk8kKY3
TmJRzq8kjPIWPGpOB0miHbduGPDS6ewrX2128f16GE9m5lvm9rpB1RkIy4JBN2E236LCVB3sRxOi
++D7xJuwxjFormqblWb1wTICnK58mCqvot8zjr/XOfFpsoP/O2Hf67AffQ6JAcXc1/EidBd2cUeA
PTtdSLBh4o4IQQhrT36gDLVWrGzLdEYR0IwVDIGyCo3KpccP011Kf6Ia8EIgODxm8yzCupAGwRfN
moRQ0ehaG4ZMmEsGHZTIhI7bbi5JWDMoIAGxoem8OETNeoSNIf1WSW+tK++MtjrxRb7FrsDziAd+
f4i26krS69esJsAkqq4eTHFJvfdf4+DrikK0W8aCONjyrRiyohgeg3beMwnOBlznxyStXkhT5J0e
x2+bcRBP/yCAGclhyCL+72JxKZ2ngKWuWIFKtanEFoZ5ttCUfeBefC6nDmrhOCfv3Q4XN5rMPlvp
VDUzmqgPabvcw3yW3U/lojZFsUSbzUUW1Nriiql1X6ePzw2hUbTnwy4tsQBeCUGY0q+eiNr4O2Ce
IH30VGtLB3F7a63FLxRt6LVwimCeLZHGUyLp9N81Zi7ozHOAtT0ScBppaOed4TkqR3bJx7+vswNm
6IbwDHZ+oh6rgltjX0Pd6PjD5Hg3Ps9KJME4HLVEbAOH53aaQTDDBBTDOMgGK4+5JtG6OXv1FkWB
t+jzjQX7iIFLAPstkQk0e2JmAg33yYI7fchJbB0FHcOvmxdOX4L1EaXriIRiRQ9D8y48zqoKpjS0
hkdnbIqPNUtXh4JlsvtZ5Oz7M0pTayLB83YTbVcRfw7XNd+4gZeFXCQoNIxPGs14jtFRs9btQUmp
xHOfQpkvLC7spKIUzS9Na9jt+lQ+bbaKhPQ8VAoBJIGw09evrf6jGpx1ZtRPqPsOXYjJp5DJ6NQV
ftwME3Us87VKO4xFbu117ZTkVCh4Rc49DP9QX+VR0NFf301Nt3JxAcUJqjMYaCiXYW7S2sUKTney
62AheXBjf7qqNMV1B5q6EnHrBMlUgBfYEEv240WpdWslnUjw+OSkD5Jbic0B/lJc2P3oLGpiAZrK
1lr+YTzW+cJnZAGTFBRURqLdDfWOErycHbsRKXGziBLcnZXj+2wX29h7y1Iqc6tVNI85/VT7pS7E
Jvxhnu/MNusrar39sIz4Ly8vEqaBYR05fK5Hk74dlMnhkTYSWzq+G1Bbz3D5FwA6qE5x/IVigDO8
0bDrSKAqJhM6PRflMI/UyQ14mwC3kK2j6LHqr9ztZk4RPlGnKP7uuHAcj3a7IcgelusLGUwBkHB6
UJ+cvStvvKU5+siK1UW+eGXmRbndbs3ftNPQq+fUvBgK5nFuZaqYP/OXxZmK/A4Ne/mi9qyI5N0I
gtA+b2OP2VWRvSsK4yW43AqrzohJaIwH1ycNNcULO2q2qB/o2EwLys9j1DLC4Gugvp9nQPhIBbca
17mfAsT9z5IgpFuvM2GA5waDpNLopG4nIxD6I7LdtF2AozpL1Ua1QQF8nm/CEEnKadjPCRWWZtug
+wfN+aDBu+UTtG+XvMKtnhd22/fFTlOyekli8XEJkLohhXmtAqhKbjS21FeHSp4ON05gcY1GFpb2
ccwuJtEBKEnQNnkpPhwpijMrYNI8QXC+bQM04Re3CSNReKs/GjetbRjInSkPbbDqb4BL8D7fnouP
KdQwQkYrLEYd7XbXl7rpQFmkZz374PpQIjvPFw22pPvDLfMNAdjfZwwhroz4QmYF0osqzRl9EWN6
YucsZwu57Roxy+Im1RfTOY5QNVPFWop+VzoAuotPWCNfDq8f9C7ehDjF3DpDj9B5W93Enq1GYx3V
jEBuzEtCwLrP1Uj0O0kZHEUSqaCJh4ZpjxagSHVYYB7x4+sJWrCu40BIsZUMxi5SEFv1Ih9kVbe+
R/DFy4OdPa2eenTMvfvmA0XmZG3GVEvZw34AAhsuvdlFIoeDISVDj4z+WyGlz85rPxWFTNvH2X4q
Q0HJzXlqBuFjIJJfFc9nVkA3s04yvAQJyiQlEF5A22S1D04SeM+3mzQzfBey96eIeNOvDzGSOndv
3YYot0Qd1FqEHNVEGtUDQBxsab6MEFC9C1/Hkf2EVsuw/DfuBtEeyMTc6KXwOE1dURFR6VI1EVVT
+HNGBd6VG0Mk841tnHzwk/rPLXhIcikOV+Cq1UA5jldBMu1Ir34K4X8iaojb7XgCHBPYkJKQPP/Z
R2//ORkIKDnR7bXyLF2xvNDaPWuaj2cc1k7XzsJLRrFjBtMnYh/G3hy476IxVcm42pigVyZopFXd
VSBqNuhRMESBzL257LucfzAaRRgZ0+vFCr2jdzex+Q5HjrnWVTjQ8FmFoJeN78YHWH9xz8U7ySqI
W4mXRlc508Tb1g9DljICGU5SVdpLyGcNAtdhGcCbYQVSdYag6SYWSXc1bchsT01GPg3cE8SiF4jt
ScuTfzp/fcDF1TAJbdWnCDo1zFPCJAjrwg9NpcGgBE6Vw1QerHI+aHzkeO2jMswmkDwyfEavjj+m
8VyMNmb+J02J/QB+FVoKyiexOYryKk3og/SoBwPlCO4WFn40/E+JCD51FOXysH8S9ZJD8g/LJ0jk
2zv9ZwT0iw6nRFjHGSvoNVwVR9R+No4eolzNsJxQpFN6JIbqtELZN8ojaQQ43SA0jFF10jWUnXTk
U2TQrJVK95ia3u3lDGWkNIhSwA8g5/KTzR5ThLpW73FUuurhVt3ExhQyw7UZbjty/ggDmGGbnYWh
qo7MX9ACjKSEv2m3ISFNhntA5Y5FgT/i4FsHFygSoSRRsyUNHR0msMrsw0cMKZacXoTGClUiCKhZ
S9/C4yxoWmS7KNf2EIyf26CZkco/kHL6v/uY9N3TBtZ59R5x0pjk5PvcZ5GzSYt9/XZOFYRAwE3h
P46blArXNNaTJ2sFbPkK+crOWm3whPuYVYDN0YerVoHSSt5tVjsGo4zU4QOEa+LgTnrGmi6MVN50
cHtRtsLmuNJAmy1bPs/srmoTOFS7HjLTtcMHvUYbtnNfCeM54Ln2CPaV2F75BP7tV+qvRnac9vDT
7UYd+MFqc9dQQDtno9ao0lI+mqjo5SKDXhWbNcPB1WXUnulTa4eIyExcPPWoJGcvcdua6Q09GWLB
8c3sI+5yd8g0HdyQHXju6aftP9jJ4XQHaALvXBa0JYOQSSSOXyfRsP8qVXTK8290m68FNOJ9gXHC
/OhsmWp6eW0JCJTAh1iGuDiZw64eLfX94TwTcUblKvpQvXcqqV1jeBLdMQqeN/TozZifET7iMduD
pEPF5ihpGXY8T/129Z/g9K85Bn9hjEHL2RmXUMLLoFabTnGyOftmwhegQ5KmnsFJIHFMfkPRpTVx
6uM6Zxi6N31tLbOMfcxE4uIscr2Ig2L1wr18XzA7tknQc9bdTMsLmWqPephpNNcGPDlRbDa/htqD
PbSJ+rgRwjLIiRCj+6/kHW+uPSsKvDtKZZAwzI0yQDQCbMfSoIB0JSSPUVzU2BX1zfrpaX7mXsyQ
Nx2ytO9gX4Hg/qdSgMJDRqTBxCGJwq5zpiAKSsMvYJfLbGg217EygygwOTnE0LRLsed+Cr8AboWa
fw1fRSz8XyhWAC0OX1gdxKt1D/uEXV73u/AyJp2d0nHtyaggZl5iqpY3HiOxYDwy38WpP3BgMJwb
NVWCjNE+HBI2y/Q7H9XtA0udoZl/0sK/YEhBOzyFT11Hk/XyIhC4jqp51/YPblTw1+xkkrXuTX/m
3yOQvnMO7wDExa2+J7QmqEei9jsLxpnXYVsEdxspC4axYJCHVeU8757xUEQSFU1FNXRRE5G7uPUn
z7k8Fbv5xcBvFBY7a6cCiXCyJii3DAj136bqs9ow6T2IyzQ3Q0hbY9BXWwBe3bApkjDvhKWWDkpI
/mNPeRBjadePychoHyRlL3AJDQFfdSQt6ZUhZtkyPeaeuv9iKXjnJJqvNVCPzGhrbyoaRodqgEQo
mnvYyaZUALNdjgpWyGYwR0VUYpWtbqTgo+zafzc2SdPsPfYng3Ntjxziu5viXQmmOmjUgvANL0cK
AYCeQOnu0zgmRSi6gH7qbcfEhbp2gmUZw+XLFLWpqNx7Py/6d81UoMYsGsCMN36lK1hDW6KsNfaY
MVXJtGZsSnOEnHBn9rbjUWsxIniSyJAVpYUE2QPeOVU/0mrZMRPDZg0X+B1ga9x6aO65CfdkMUyC
j5fAdQaAdCZwDYr1XfWvy1hNhLdnpn0dqnxgyR4nwcDcBsMK68Rg9JnhYFtZm1yhPTp/SR5nP2Lh
xHv6ZnJw/zCzNipycLgnoRHnguP4SsIp0bQnVXh72LOHJ1q9y3RAkSUFWsdRNmYdsxEEMYwmUs44
pF9sEFWEmDsk0BP5dZcSPJrin/dEHJ0G8xLHcjrRbPEWFDmfqA0JHms8/FmfwpJ/uuvPwDxMjV93
URznlJ5/MTG2HTiWRXqcrp4yL3N4XhFZxJVTQY0Qcz1ElT10HkXXPHU9UFHnnnkSbgJ6rfKK8VWE
geZ/eRLPmpbFKdjBhnuOqiNrjw/z5aUXNjzDZcqbBmIRyOYlfksZlFtnWYXxGzGl5oFUVm7CIDX8
xr7PJgKH8+5aLMlSiRX3EPPk+wbayf2oyVcGQNCfzSd0+KtkkV9NXry4DXJDv93DXYgoDtoqxM+G
accPUuW7YX7eGjIVp2QAX5Ijl2BNvCmRpWD2ma4k8Qc5Aj9p/veOtTrx3NZr+LWhuWIPlyFjYh58
KnpPCSTKBQylYZnnrOoO77SjRf0Nnh9FWKwjDJWtBOhAIUmbqNljP/n6prOdqLZe2Rh2bv9HPIUs
n9am5m7pJeQVsVQPLYU/tmaWrTzDBOi+Cs02y6nFvZESG78we2ubOHLRP3Fz+PAxWZKkb17WbUP1
RxUNCxWp1XObTFYNYgk7BVFC1FDLWzgS2rutUEKhbexny2otaCnKDMmdgy5AuEdYWh/y4mnVFOtJ
1dLQdnC2NrceUD4VBhzaDKXi1gpZ7V2agJ+/+Gu8U4BfcviDmBpmNj2VksvWUibfrpDUWif3K57P
RYCLB82ZQTJouOjD/Psk+oTnXmS5sPcRdU1QdM3c7NfpYKRyz8ltgjA1LyS1uN9epR+X95PNdibg
3y9hDf2kJb4+3Rbwtx7bQluvXWBhPzQrrIAzXraBJt+9OQbWDkSLO1AP1L6xf9CeZSEiwOHLKEch
vSEOmopqqpJzd3NAfi46i50N+gAiZe++Y9U3FNsHtB/HGg3u1ZxwhfFvU9C1Z6qx6eSRBziagos3
ENoCs8GHbCHZpV9VSTzVZyi5tVIqFtuH+JyCH44BbxBN+SXdNQ8V+8CYeREK6731MMwTOGM8EnG/
L6xERHhVdU5iq+0+LL4we4mPJMCktJvA/OB0AEwkGpFRmCDlzKOq1KACutqIwxgq5bs0rHdhRVay
tHGHO5H+8A7Da+ImMq+YjBfmXW13NWLShsFq16ivD0jdcXsyQ0uiVDuWyC1oFRjcPD0k6AxZ6bLa
vT8paXy/ak3SRURvvOafm5MC/Byn+Xha38Zkor/6QfCvog2aIDkAbtzm15V9qZ9cLSU9E9u0wJYe
2B9yYtaFROmd3APICidIGGINASTbi/QvnTWAKps0V7yg7upDBfg1EfJoKsW0SU6ECOP4FAAqzv+f
PEVmJFXkhPdvNHUclkVdU8I3Xkjx5tR3Z4rjkzR7zxLZxyzXWwK5dBel7W3YArjFqg03jKBJkQpB
ud4ID9g/B5TLbFMLVecOo2Ar9g8eqWU+pg5Q8ghbm1RALo/O9VTInno+OnUhDyi6BLrN1mUwCPo3
Ty0YeyAfYok/D6a1jiH+aaFvg3eMzxXbXMT2RGk1Ql6scLQTq0DQKFjbEmHlFbevsvIPx/0vwnq9
HILRyddkW/VcefNiN2fcrJQWyvwT5L1xBYw7bPB4PVPkQGL9/hIxUctictteXA/vfukzM2qDbr1i
MFUwBMS9p1VqpWoC9Walhu9tRAyIeDRpF5MccAVlGNmumtNqt753cOrFv0XwXpzX4iph8eKOyvb/
ywbJdXJnYMnxBOiG3t3PoX4+qNdPm2XGiUsRI7EDPKs7wioUjnghl55qc9yLH2AkgmD3I9cuePCc
z/acQSm+0s38sdwFgrcm0KId1W1TKTZJoDu/UglGMY8WGJmwJTWHc4IgYTc/Uw4hthLIcNoAc5MU
dFTPgg7qsNbAAveozhTNhnaLu3dyao2SSuovsJhl/BUpjsO7fx8t5xtpUQlRiAog8semf5VaXUvB
DiorV1oF6Tx46+TGBmvElyWLEW0jQi/rsO9CtzhDNJoHrpXmUnpsK3dlndxWBOUkijpoaaTpMHVn
S/dndEyc+AoKxyM5CT0VTwacYBzl0KpDo94E+LlVawRaq6DLgb5H8yNw+5RK9beXzVLlQRPfXq8I
6WD1bawdIESYyzvvYFxjcD12kYPAYnRp8RljbNIndgPFXVnVj8vWY0JIlvYifgj02/fu0xGmwIAd
1iCaiBcuQRIahsl352tvnR2TkIbMW3FvF3TTlnbwbPAMWD+CIDZo4mgSXSkkBpuUKCq4ZsUgIOO4
cojQDqrprndgsYwaxp5mViIewUTP7OyuJU78EhsFFh35Latrc7Ummne8Ia5MBG6uveSfgWUY9mJX
yw4i6XP8z3GOtpBQu4+GwLgyn7jM+AIMjUklPi+WNlrGbUHVaDZRtd1M0s0tV4yekxn8KA1Znr1b
VDGnD4B97a8n5eeFYS6qvsz9hkYrKNX7rb3POZYNZbjvhKIQXxp/9M4AgXcuLK6IHXd8i2gv4Ls6
MnKXQ5g+5ec8vtg7YtTOWDgyF4H6IdNLM7+e42JRBmt/R4eFQAanbGErgwFudW6rFl6vTB43YXYp
b+KLICRDZz+7Bma0Qbe5DOOUFZQ/BDUBT3c8yn/UqTxb8SlCfzmFmZvIPeBxdejtPWLjO1mtXV/V
8i3/XcgZkzNdRB9LTVdJJPGsZQEyJrSW2PGV/FPF5p7Ss/PkhUuwgz2JidBhpUHzwRoOouffDvnM
Tw9nwhCpv3jAbyKhLHY6lnHnAt7GX0PPaFGOCyjBPXy3L181HzCfl1H+gzKjDG6iNAA97cypdHLF
3D0JsaXyQSjTRqwBEDS+gay9sCWl6v9HYsT3cu2JB0WI2XQRVsr9KFK9NCJ55Y8zrzvCfXVIyuXe
FUXfWl32wikE4710oXEA1LJaV1IrNsyGj+Spx/hJpViMkOGWF4n1yeC+AC0sFBU6XvWEVWR6Du8O
cf9czdORdJD+YvMbETPj2i9MY5fZryd/KyiNaQhOJkJ5ZQT4zgJscJqNYzJnz0CYOLixUVZQIAtn
296tcsdKW3wAuEMF3KMBNMzbLhhvzU1WKZ/joMnb+mtnuC3MpbtI9XZwN8e/hjwpLt87WyYrpJZN
bSWRmy5RP7TUtb48mKHzwOj0F+/mWA3IPo0lHnDb1uw6Ecau38RaWixiPzNuy/f9/xnXxdFIaSRh
qWx3lQi0zZSsJEl/6Yl5R3JPOHAZTUrVjUPn1xIdt4KxpJNbM25Z6gpBbiSXsVY2qGoaqHf+Dlcx
SwxagAfGXg4sikhJuGJ9Bo+DLSO3DXeBBnBRIV1jHzJCFJytYjAkxp2k4RPqTJyzysRdvg4EXtgm
o1/6g+MP+P63Hg+KeQlzdLuQm7lv4rwf3hcnwXe2a4EWF3VhS7U/vOuqfXFWmkZsl86onLALuP4E
bCigAnjMeS1TVcjztQLz5pTr3nq7MGyMY5AQJgx1w2QauZjvBcQN+qiuoKDkacv6Uq/quuuNuu8F
uBEVPo4HyAFP5E+jQy2T2QSfnscAASBWG0MnlVU3IDAHn0950b5GprcwMfJQ+CSoQGs7VzVyVxya
FQNQ6TElefjzgivHT/zx3pPhq2GHNu6raDBsbdzjySIOJRIrfbozwGU6QWqz/q027akoOsNGImUk
bsVKSRkAOi2VWfNja6UFhPHVFkpHqJb3oA/K/92ddvgxlG0ek9o5sCboU8/HWatbhUf27wv8cKM/
lhVD7ouLgNiEUABX3B61xbpkPDQ91isxIFQvD7brjwoZUK4G72qvclfKzVc3Q8em3wOZVjzFfiL3
Gt8wvRRNjlKd0lJtJ+WnY62KeFh/osVAKPNfa58HEy3aAaVE3mJyNtEuAsZWV3XUqKNv8Oj79HoA
sRumfnytOqSsDyEqMZ5OLf1rn3Ry6YrkC8kWhiPULFI/J5ExeEYfvEf8rEE5heL+V8Mig0RB4NgG
Vun329iMMhxOf/VZKfn3qTBptNzglnmzcTYpo9gf432SXEmCb2TYgwLFqluA93a29Rj6rlrNikDY
5072YXhlD8SwstJK0VXotViE1YWxyWLzQYu6lmoSUpbZqxCvjHV4jS4IeaqXDVoi/g+Ac61JgAWe
MEPsk9FNzRtRxWjnmE9PPeIUv5GOzg67c5gLVE3rUTDWuPjEqdYkS/0rm6C3VI51I9faO7KltYF+
ccRKE+eDxeCk79WjKro6a71/x8oJrVlvAWr8WHtcmGt90wHHfsNYdeybeOIvoupop3/KvTufX6Zx
Crp55rAuw+C7wjWqkMGL4oFW8ICycwrbGlurRwuitw8n0NZmnp0MMGc8HrthWAH5niZqid90Xs5U
/41T0/nriI2LjJDJmcDbObjXy11kE2rE+uQjhEFmvjvLFCEde95ukQvpLpw543VGXYKRCETWB+6H
/cnsf/1qS3ZHtxQiVUrHfkdNkxb3bCnA/gTVfXjsTPJZOkpJftVxjsz0Ix2SMecG287seXjwjbtb
zRjQ++OZ9H5GlXIegj6NZPwJDniZCIz9K6zJj7z1r5MKpYgG+Qmu8DuScFsUKcNTX3p0msNX/3xz
xWcR8eV20aYKpSbVIOHLuCqqJPML3RGp0Uq30rEePW1/DS/8bAhfhmmCDwFaH6okuKH+FUVU00UR
hM0Y3wS/7jPB6eGgGxUiKkPTtNMsHUB4/cIfzImc7ZJYWCIrS6wG+1LVqzdbw2t2iHnPu2nvjI4v
Jv3Brb/kP+BcDN2wkVhfklVb9dD5/gTpe7dzfEHefuowaShVuJ8FjGdbIZfXeMeQ7hydKYbnQqLp
cCYm7Phqx9WidRJfloRtFNQL7CEy+3RZ/Eeo0uVx9F9fwqJWyHqGGoZnR7uPVHX9ips+tIZDfGTz
9gGzt7gUZR/AfSb7bLjrSOxbXQ3VkKJEFjzPp43rr9i9kfA05x7qzUT8aXVauuVEjpEORciHIJiY
wp8h6GRrqZIfll3Y2UVyWi+au3aAcx1wRofO8MH6+ZhlNKRXfTdriDxS0nGHiVscVVzpBaDOQfGG
QC2cKNjhdN5OWeWRBG6LZPMVCnNnDH8/ksFicao/LN0tabdxC+37+T0F7kLANb5jk6Hh8qNuKpDv
2BUVIfwIEN1UNxw/VOgZ3ToUNZ/Hf5Lie8RIvo8ziblpzY2tIVIxuwffA8WkPGe0MCHZ/msFV9Y3
d4YNEXVWuawaUU+HRpWpI0AYDWQGNq7WiGoCFQvDDfqjFzbKGvgAx2t648UYCwOpzJpTbj2dp8+b
lB5coQTlYGJjeZ54n++tWGPFAyU4z4uku5IQYB2m847E1mT7p2BFkdZuNemX0YUnWFpsCuOc+Hja
SUo+kDCkuFcaLiWVEPrfqUGD9o+kcj6gVcJtGG6f6EA3Hr0e7nbl5zevMSuta6B8EUEXlRBqWgaR
r99r+wF2bBDqmfFwp4DNf4yVRiaoc1Tez0Afl9JMBdceyl9u2oO5VBbHOJ3nYsVSKftUxItDxYJg
kMYvHQc8h7NYRIzBug3fobH4I7wFySQ7mElncsO05p4js5yTfnB1Eqwzvd6IQgdLyZ2hoAsmttSS
iXpgXpL60Pa+J8U075cKZ2E5njqUuDAYLKEWNBwjc+Fyp4708ZGqtQVClJx41kfIxCmHRgyzF9/C
Qw1YBYfHijbb4T1QhYjXi8yoTpQZJr34l9igzHOEFeam6zH84Dzm9HA8FkNfQGnRXLm73CKQuUVC
Msb0OrKbq/kx7VGDDGRsKHhm9/o2lpkNZe4OmiQbmkirtnUnRhwFu/l+E1hc7Sze0/iuJy2s5WSv
noNXdIyRCG1gUjfzdNRsw9NVbC8AqLdemD5U7nUZ1dC+fAusv6sqoWDTltdOUr75S7nmu2bieNnJ
/zz0MpdwBsVtmkv5L1jPkP2hOAFTe3P+pY6rSEMZvm+EkL6YWm0zawgX6Uqr3hOai6iQZDVi2oOe
UJhgNOq4xTgqM/ndfEwbK8GJJ2aT0ezNyxCJEpGOZH2ct10a4dN79a7zpgoAIfi0+L+xQgkAne6P
NT34caKDNhUrw5K+k00ySCaV5xuQB98x4UnqQFSk6CsIhRCJA6RH9U3P761FnUsdikYSW/RqlWNC
u0itU1YhV06skeUqfYCKYRr/Ll/cEGdgkG7HD6EEGIe+J5TKJB+3Sc2VkrxPzvd6pyWfNwnzxw2t
G5q79NPmoaoQKob/C3GsP6qrj0yW6WAIFsKIGfwq6pbyHk9uDEhuFPOOIDNLKyIrbNjbaoGmDNl2
vu06CaaXBBVqY4i67mIQkDCgmFH2rnKV9K8mKeAY4jaYVNDhs5koLP2XZeh4QKPMQMUz8yq31AiL
sLldOwUptdOGA+w5yJb8IZLElRcLTpltPrFCQlaN9Di1g5C2ZNIONWVHbWtjQzAXZJLazigp/gqz
DbXygI3TSGQ2zApHkn2KgEeMhAT1c2hbeIWfZ9sUs0ub5QVum9lCH3wVq91wdFeQT09ckxZzorPH
wRzN3+cWxiCPFfupl+m6jFl2N42Uta3ouDrYzHppr5WIk1uaw2W+mG0XSIXb42LFXG/lO/vnegEh
k0vDpQHFz7N6uQVYns0VObsQICqdbAN3mnLG7EHs8Vfe2Mr7Nzv2lUJK+a5lnDOaalIQBRKXvSZn
2O33bMEORsw2Bw5Wp3FDAxNUC6wBqPGgsmrnvQmkrKfUU82lIkViYAPJFu8U5BSEXqGY6YN/ZP1C
ZcKsiEyHre16rQdHZzXBaR1xOL7C2cRcx6/E1hROId+Q2K5nr5KHudoeqHzdRevLkMt7Iigv5dfs
l81i1Ht4opgClZLSeG/p5r5WNeuHSAHnnGcM8YG1buyJt1qky5G9C/P0qvLBW0j8FJ/MM0tnCVkD
HUfmZEr9voiKqJOl6x3v66AKIpzDj8TYmNi4uc+5nkc0AiG0udsyXUj1q0c9uUrqKG0lsIMsMG7A
2uAQQZ6g8uPDQXx+1OFAq+Ewpm25uUnP9fHWMOXX6JcM0wmNcdd2srfSt5qclnc6VvdUxght4ONd
66WtpBHIZhGT3lS8PKJuzmNeDpeXJc9ZTALc8ZhleksbzZ0onJmM2ch3sfNu1pIq1xqB8ktC/2VT
sBFADS9xu5bTC1wFnaxTnj4HongubVBuLMF/K8oMDiVqCTdkvXuX6KwxZLkritczGtO+gDTk7Xk8
y5sZhY9sP+FiXL1SzNrcYCpGUo6wa3NrO9SVDQPln2iEUYJv95rzjh1UrqI5j5qoFzmoTEW/F5LE
3dl9fmXdsdMmkJxetx6146rAvKu0nFk4ETXDH53o8J6EhwwFWfyPL5+jZpgM9atPxATkiRGvOHNj
RfB3rbG+pj7WLc87dNXxqsaUMxb/zsYYZbuk8zcHXWCbRxjh/lsOsJImwFs3uYD+HreHnHpfZF8P
gWMqkgFQERtJNMjVl65NwIgHH/WSPO23eVU44PwLyFbsKjDwrUKgWmLDi+i+n74Aiilz3c+NGs6O
WyW36tk1yxBOGoZEWGPuktVtlWwyNHQTza86d6q0vMUCF8jyva5USHC7yjc1H3TVM5eWw0/XhWLa
4tT81jna5yGcNZh+km4U/+g6GJ4dE3zmVW+w+by6BGmtIg5HfPIOcs2A1fh7YWqRGbIg16zazgLx
U6e4B3wVAg9CRS+pTZJg4gM2Qo4J5HF83VIaRXFV3eIEfUx/Tsjv5/kY/WeDJi1fnUGeavym8YBR
ey0cavYRx2RWsjmBGfBtPUczKtX9LvBN1Yn9xaL0DEmhlTHjPwLIToZ3iVO6fIvhrLU3LBW18Wtl
dy/0VbZqNSn3snJqR06Si3EavcIr8vOyXQUzqKXTcwLXUH4ghmPs+rXCVABUJkdagQlNyu71WR0W
gOH411vQZNebv5/vXilwk646nXVkuobdNOEdfb7OIW2f4agG7tWPWbEXzbmXEUMWKtL+MZkdX/Vo
BiU/56D5EifvGVL/L9RBTZYMR0sKaxV1CY8TRXafEZAguWzCPgVrX+msLakllHu20t8zoBaGw2FG
BmQmcH+ybLaT65u04/AI2cNyWmhvrm56GicuDDl0stQNLeEhkzNmZZ4HYFaEefYRcbxAFIxHPYtV
gaNMoWnSNlBYqsRIRYGnoZB2VmAd6gao0P2kilH5BBa3MHO3LHCBRWOpDajEuA2+93aNiTBKvWLq
PyVI1JVFq4dOQuTPS3pDAu0sJfl2pX8UVQ3tcJRvYREAruSdzOplvjLmgenpZYDmONlg8Ff02mGr
jyK+4jpfij5vj+DiHllCdoFn1mGZo9YGSBrMlanEk6viBc76aOVTMGfC1CH8kxp51e6HHWeGq6Rw
nEiMwHjbZOb02htV4BoU1N22f26FXj360LAodvivL8pOMFDgLWfBXGuynvCIqBiM1y04eqFZfsgH
qlQfXwyxqnTUkPKja8Qfl4c5nnEhISvTCzkXq8CWKWMn8Le5aSTHjJh1slNzSRZvHPLzdWF0T7Xc
ZEGHpvnmM7kvP2T4bAHtIAWN8aFR9pg0JUcQexV1DgM95P9S+ict6OVc4XT8SiYNZfBpcLSkWd+h
nZYiuOiq65jqBFUZHCl391UFeu6dBB1loJHxlPlqyT1cGbUdaCrh2c0nchu1h9tmnCGansNQAfRq
XO6NhCfkiP4JaQSThhbKeexce/Vjs+K73Zfgv42LaiM58742c/OApFk6EF6HzGwqgO84C7Fepcnl
H4Z2DYVDQStuh6nDKfw7l1C07enYVq6tE3lMQ8d/ZaOWjh6v7uUmHit76D+vyb0PUb+Yl7IN/+4h
muECxk5A4ZszUAmuOon7OfN6qIIQRQwoaKFJuXcVIuu3K60nN4My9IC9OfZKfo/w1uKqdEUrBrUS
aPhdR/5PWByrolAX1Hzc1MgLew8ANoQ5VoKUqgXyJb9aHTukBGv28YelmQrlwn0ACp4d9J9Y5zaf
HDtK5lEDk9+RHKELTdcSBO4vxTWCuXWTXmgcGZv/yugz4L6StjMdA5n7641vaDl/vqE8HX5aEfb6
hctqlsu1I8svySDgyGx//b1iwDkF8IhlqbLBNT6QeUqUPsUvAgK1wV2BWoAJEwv631PQu1IS79F2
+j1QskiWUu/yCxbR0mvYD23zFNz+TA7m1uGSol4ckxKbqsFrHkY7gqvp9q4ByQ9nmfv5TOAiiAmM
oGlulPZ4AWY5SBJMaYh2Wb5yq+k8tRx6Ux8X7iALzU9GA7xrg3qqcoeVxSI3TwobgEiPRlNuDUJn
rkd7KdqtthZA3QiQ+XpPKlS9h3N6kwuTNPOP2VuMomAtas9ovGifG+D/09mqSqG20RCcX5jbbCqj
OnHEW3cJLL4mkqIuq6c6OgncZaxVXtG+dbpS7WdluVqutJviMqeP3Kx/7jjSRh2QVTeMOSf0Q07G
1ZvQvwZYXZcxHT+TnxeaGABndMFtibuNRwU0GnmjzaPH77m4V/RuckDJ6ekR2fg30g6x/QmxUttW
g45je2zLIRonG3smSnwDpeuRj327XuotzmJhQMaeK6SacBdYd905CMNZfJxXFr/UIjj0v77MeDMp
82TtIfkPkfb5bo/6PwMOJ6zm54CwWN3qkf0ZC0OGFNdrYgzpbm7IkabxBmHMM4/ttrMIDe/Mtb2b
St/TB7iRZjgvkUTFJjlE4aEqWmURr1VN3Rt4b26vCjr68c6UCdVfRqH4KPaovr2dexIFk+RqmY6+
3J+6SrEh1BM+L7wOAC295t1hXbx9Hhq6ngytcC23YIOOltlo8cBBrFp6lTXxlKg7qeANkDQr93fB
sn8Dhdx2kINgN3qfyieABNEbdp0KgSfAt/+iP7u0S0FPNFW7asE07FC0/rFK71uh1frAqbwmM/f3
1YhtRn6F2X5Gi1zufidSx0ZnRVUggUvznLQCCD+6tkyKzzTJIDQU9cZSzWMbZ018PBHj/mp0rZjp
CvMJawsV6rm6sjxdjH9vgO0kNtGCd3jih7hm6UP0xZwcHin91Yg/oVVexHzjtZcWieqqQF+LuAiC
/j5iVfjVinoxRPQiQmaIGJ3sOJk8ajxH5dr3oNAEQNUsrQw5G6x/OhIj5hkwnPdipFzRsVQKHu32
qIR3Xj4My6yV81GTvsRviV5nUGjyvHvBW2LaU06jRWHasSonEyQBzpP9zobZKmbDfPgeIPEm0WyP
XEgIiDMYzG+ReHfF3fBaGqIBO2UGb7f21xWOxFWZmqojJNgj+gfZDzm8+1UQC4wM7iqnI3f5lkGU
v/8Yjd5A7Bo3s/bsfOknr/JtlKNBCYMfUclLdUCiNk12JNvpjDBP0X9R6/FkSkMyA3TVSUbhy4pe
VNIybAlAQ9dD1yYZWybNJysduAjPLLuQ8zu5vuk9TldffcdhKXkcAyMX+E7diHinCKWTjNK4tHuE
Npq+McYjkeyIehuyW9sWWiW4qvD/Muo1bO4rFZM113KDz5FA25/x0d4lasLqGf/IkB60oWqkPrjD
80OhW+1WNkmsRcVnSFm8gtne4f+DRoT6EKackvjKx5gVnvrMqiZxFDjP4Ne8a6XJ2LtL/33nRviS
GxPSPMrPaUXb/qED31bOPZK8qhmuHdM7m1kwhNDdrWgiYYcktpyhMTCn47kLAx4Bd4WY6rARyT+4
PbPtC5l+/0w5+DOwcPNBjM6yJmAlNaj5Tk2ZRkRIg4bG5OvX992gvaCubthNIaBHXNBvzU8Lyc2U
8GLhKRYaZuPEm5zqtCQ3wyLx8XwQeU/N4aQZck8HzrBqHLbZc3RuLokbWoq/te+WB7EFKDzC90iL
upyibkndc4fr6xCShW4mhngiueS9pIeGchF0K0hDkkpI50Ls9PGgkly9VVg9NEkbm4Sa4WQ0qJQE
WOxPzLahT3I3aWEjlW3TMtbb+uL7eLS2fDKSTTiogwaj/wqah0aBq1bso3d9c4B0yEUQ1Yix8qMK
gLB7Rq+oF2gZ5zTUbYk2mJ7BqBEqGz9vIRl69Eek36KJBPh3CSYeVmwzxSA/xP1T/jBubBu4eykK
Lt/PkbV/kq7XnOFtGeD0Uhs2wH8evDJbNDroSPkJAbHI78mye9XJawNw9GSZVBDLwxmjNlPGXQkb
gW25E5S+grzwsK6pQB9sMJWVMCsQtvoVYuIlYjeUWMl2GRusZ/JYPK4zS6cI8qeDvKFi13d7HDuU
WBioWC9G34i60oEMrO0GpvBIYEqqltGM59bkJLaK/BGsaN81ju6z6m8RhDGlCXbMSWs4cgj4Mn2X
vrgJshw3JlvmTGj1g1TljX0Rkd4hFAyh7TqsczEjb3YbxVVh3yuh9vD7RJcnQPK+3VFmWoCrM89i
ZxM384oFNm0HjufiMAsXZ2P7Sc14lnTP4kfcQGUM7Xqy7j9XvP6JJL0QVp5kjflqdACHelSTkKeQ
6BifYvDcpih3+RaF43JtCrn16Y3DAxffknsmrMfgSesbwzQ/dfUw7SwUhCC/CwvHtfISMP0PTKSw
8IdKfxQJALQP8hYSzwWXxRcdpwXJsM+mb0g+P0OEJnDNQTShI6Gpl0+hagkfQWBhLzaw0E7+4HJq
oLSx5tt8pPCR9tnV+vJr9hA0Q+RAMpedur3ts13w8aq9YUSoMjZfkxwCl5HwIDjfz6o+3aDL4xwD
Hq5oBV3k+B+8eJIHZwCQUKlaAzowHdyAeU0N6N/EOkhKkm8XCceb9MuQEB9kV8ygXIjwWYMV8j+h
5Zfi0jglvxqYYkGwrey7npvgnumrUU8WZzJ9H5ABdA/NPlyocBsxGnSdIx6gCYkK1lISZYDSAr7N
x6XAO/b6q6xT/+1hJN8qeb+q6Wvj1DOOECAmueui4LneV/VhWSejXIrKfyBrc28NFK6Nl31WeX3V
HCL6PbrKGlnZ/bcfo/eJunt1ZifJzgncr2yAdYI7fsAL9NscFcKA6VjWES+Wh1Y2wlXyusB9oZQI
HssWXzBh3fBZAcw05Lc/8fC2YlGb0V325JKeI4o3hmXVPkxDUJwrSuQm+xQEGv2Vcci3B1vmXTdu
kZX/8QNWXxOTwZ3NYYkqk3bP2ZvnBM3tJleUa0V4FUMC7L4i4hYTc7TRJ9rex3jv2F5BeXL8D0nM
fAdF3m5ZXVGf5cmC39hbH7Qtt0wAn5ibJYmMPBA9dcpFTYrrUa2Vnw+gTeCZWzcd06IJ1GF6sw7d
ykM5yT4vlWQuZjVqYooOtTfdi5DMh346w9Abk6+qmBkM33aPBqR1UabZ06IlO2Lzxgu6beBBrU3h
FCnEG9T3kN6gcN7IvsE1kAFae3JsBh4soVev9XzuRGLrqGnpTkY3FOmFBjNURmdFwRhsY/5SgudI
YqrGLVduaCDGUAHPbwsJ0cLzKCcBv+Gu2rX5EHIp/8lKXn02RiQyrrfQv0BtWE4lk+fTIeRjWskM
2f0FLyUOCEl8Ux5pgY55BYF9lZfQb8LVcIwvbsRbEV+jGOpwpdW1CLHolksY0ptrJubKXAt8a6ul
Lx0qJ/SYtAZMgzR8BEMPD5Rd9JerJhxpKFjmskaNRJnKqTyKXOrRhWOImhfncRfDxGqIohZFncFH
j+ZMwXpzGlTNwP/EgewMuc4FRL7zKelhotIB7WMfLa2N6A7WalF1lNhmyxU8VlH9PmQTfhYy/B7t
0hNxwV7m+Cp0XM4BCCN2lzdhNNBaJIWd5iDDyEO/0FBF/tr7LDgc4TxygQQ+C8DKaEf6oT3GMKYI
dCdzNmfwIw9qbK7LyGVY556qJ9kMsAUpNf9tKMuLq6P8QsIvSTVxKWFNPYkD3jDokfLRarLn1KxS
DyWO6La676bEGgZ0Lb4/nEsU5j3msUcZWLGzcj91pqlMURdib+nUABpy3jrHZZOrDzZW2gZHUTFM
lmM9K0e4tV0UgVSxCH6fhy87gi+jGEPuSjEGwhhACtOqOYf9FE+xo3qxpa+yH7UpB/CYVn3L+EDS
NeMxoIMklkPwlzeDZ4JxLZTGsGphDovAR+DJ18KXO6xIlDUOnjM57sytP8aN0e78zkdHx2dLS3Fa
GWzVdW/xJXpR675FhDSghfFxbymDMPlRgIVxD6HpQF3Rf1XhxarKmuQDbZoHzkMkRkAMjSzlv7pc
kf/HbJ6xTDA9yn69YCnia3UXiHbpuMrIRcMhAjsqQ6PuYKKsq6Ny/Scb719NCGRhWZYCiVUWBiZ2
UX9RJcPYXkVuudgZ/3YaxxuBiZQGYgd27bBwAR5FaTzt7jaI8zASiVxAyb8Q2BMu7jnED3+S50YP
ebzmB5y+7AKDguxyG+Lb1T31JkSXVGfWYA74vm5DCt+bWPSY74DXk1Sh4LWjpuf4LupDhwmcY5Oy
b+xgYLQxlhZ3zKvNdw5BzKJrEi/NUqQcu1IHbV195uSfc51IYrBWil3MiZZsnOa/MEBfR29A6jux
VKthmAeU5xAIkZUieLPnaK8yTjYj34zRTKMBNEye0EE3RGn49vt7BOn6IAXRs754r1PLRSx5TutV
X6fqupPJIOr4oC1qwhCn+A8XXsVbEAqL1vb8TifhV/yD2hliYrRAGxbdQRzogK2E+pBA8nffOfee
z5N1f5AobpHYGbhpJC235ptxief1sje0S0y0d+spR3oA4/Pv+BqgO4dQBnhbVZjls49IdRBIBmWd
gyI68oDRJKPmNafIP7Esve8Y4LBtwNava5FE3E8YZr9wk88AeAiHOWGJlST7b2jbCPOdogDwHlz1
EvinrNbibJRxVl+NR1quAheTbqHlItZdjVDZEERPwvWbtSXy9C4Hh0+dj77vbSyNkeKzMUtkD3iJ
U6cG/3MH77LRr/q0bZ/un5BpUXQk+tcej8jqH06879LLdBxm0b7ZmJvcFvVDAh0idYsTiKKd1guA
+H6n7RExc/H5mWDxig67nNDtEW7fchvfn8rxAu0lPgZWXLzxtFa5HmkFsMfoLE+6pg3ceUwMyPyd
SLpBqT5iYaV8XJrHOr4wqGOZXXl4zZvbgMqre8xmeledRd1Jbj7cotNL88lfuNAqwb6qdpRLqDi6
ya1ensELOJuIWQClOuW9aYUP3hIPFzYhVVzlOzCQYIGygtnZNtjZB8GtsU0zkFdBu5A1tMzRqZuU
fXoPxE4ZR/CshisZUbi3op79FyFgaWk+G86CnafLxrRBecUv3iDqJdfZ82QcR53KQoFu7ajSGcCJ
3qdxZA0vYaHxpHWKjqFtUCTpbZ3p87j/uYsX9gW+GlKmpIhzs1ilp5c5En1VhZgf0irRkxr44/we
vSbb4ITHMY8AoWp1SEWudCFGj4d8QFG7I/wd5UR/IzxcxXaiq6PTdA4BIZZPc1AAjxX9qkCLqYC1
r/G2L03N01/+feUaXySOQC5nHT4FalZbrO84r3HeFvVmYs9inMpA0cEIkKt6DRw7O9N22VdsYT2v
v/cZJpwx7TzCJOTC/XPCo8StZOcVh6zOqnV3F0t6RLJVNRNRGpkeATkkJvbXzg58UEKQTxkEQCPd
x4K9oYlBJYe+RJ0pREeyPlOXoyIDG2pltfTzeYLtDttcJRdxcxwRkze3qk2PPcXcngPZU/eeRd6U
gBpA1IZbxTmm0rvZ8enT3N3jreyge6IEYja+F29XS10GqHU3AwKOTLjY/9BUdTPal/th+oInixs+
xmHRtIthoDd+zeGzg1eKnHnG7x6r5ElEy01m+RwGKErp/sGOOwXE/YhbyAFp+Xnb2Gf8ONcpZBFL
+SXWOXSv+QqhOdpogtYrELF889BHSy0T8AavjrsA8sGN8/7ZQqxOKYRQ4qLjIkyEscXRFq5hIwK3
soa5/BRFH2+ZX0abRPK1jJgnJSZkn6aJuUmX5r9QzHBMpiG2FeOmanz6GiF+AyonVF6aW8TrRKaU
LGwTQXnX8pYBDhGEcnq+c1QbTBkChwcoyme5YgM7cXENX3cHQuZTEajqLv5cdvHH9748WzoXrcFj
mvheQ12++qum1AJGAV4u+7LAvATy16MI+QiL/mMdQhCmoXD4LoRdnR3XerM2GzCukk9rFzPixYLt
LEZ0HQNWa7K4tsj24ODYp8+S4M3SgFf2qVOLCjL9W1BLF0z2XgAgS1mKi0GD45gjnC7ARNqpnfv/
qhdkYNNH0t17NSVNe6ymEC4kjuP24sojvU0ixQhggDkHRgiDoFSMkS+Y3SZX6xt6NytwdyxIysfQ
cItQ4S67Yq2qCbaPM+lN4z4cVM2KIBCia+t+9il9yUhybv459+UNwugOmBRslR6iPDsrOnc0xxzP
UcoHFz+2Lmjts1MTtU+vGuOPqv0KLHDAxWk0DBs9U8cBlnC45wxzVWaGTAHzaLLzby67TVKnSD2L
r/EzcQM6tqErxAZ30wq8OV2m0irUNOjhP01BFZg+yjq4QLyroma3gGKrVK9XvKqxcCyVMQMdN3BG
YL6cJeg+axozxUXtFVQPi0gRlnxzZaHDeoUIK08uIDquzy1oB6TuSy7tnWpgAcHBSV2WWjRTsqH/
Jp1rRV9n3YQA1yJJBWT+Cg2jsVCGkZXH3EraVUp7D3ISuaZQSQPikzaa5azUVVVEHWSARnVKOG3Y
eTsX/LXOOxsLn4uvBZO06klkCrTut7cJ7eu5D0mBtYo3wR5gFd21V1EG6OAC7VH+Ius1WU7xIcjG
szPVDHbsVKuNgaT/wM+J5P60OGhmH1OuJ7cgUHPP2jGb0VionObFkFgYObPjOu/yqAoInX9rlOs7
XlrlD/rqmsBJX3TB/AqVZY8lvqG/TV62O/s0chJ91MYWqBCfx4X3Qxy0DIccPvl5Do/oQwEJLUUN
Cj/Gp5LsUQ0B7ChXhCB5Cx6e7zXbYL0mpZA0smzjg+KdW8mo8ucJcdNgs1RjrWOlY/+JFm3XaPN2
lQdxdRSG6W0YphUsUW58GvOMbjGXgeWPoOEOcWvgYu3YwMjIUlB61M8YRdceusPwEEr2aqxoX/JZ
ZtcuS31sEW8rX73gyq6H9d0FZ3Thk6+9GAyvqCh4mHVQUPZDfy2/6dww0xVBDsbnEjhZQF71Bs2b
6860KMVpt+XUYUgkEmEl+fYWQCmVhNtAGqIWAywHBMxN/dPHbYSlCxud69d2jSKaUqDqoiAp/41m
YehYyx0gfvT8oKxan3RiKP4UU4Lm88LDKUORJv8pKp+7IUV56x+OzUW2MpC66Qsg2lG12qPdAxxz
hYMR8fZ/aitr/f6Euicg/7xU9b58d6Z4drbYr8coRT6zqqGzJyFYmfmWTTmAci0ACwJ9yKSElmd0
6E0voNnbrUO4ljLsIUZVGu/nJxkVhcSsteJAsrWT85ePE+MTGouvcTK7IA3ybWUx+PfWqaBhZsc6
DJxqPKODY5IN8gMht7Ftq/+EPadqEzxN5gSm0FgJsU6qiD4RSc++WZ4QLjFLxSH0u8nzamhjqYn7
dYVb7OR9bbI5/ltdiSFAvRBF+NTdmQERl1O9MRfmd28TjtX02cYUTFBcjS/QRBEmWQVTx0R1pjtz
VBogUSeRDTGmMXzESNci7yYx1oRpk8gActiRnBETOMnkrRfoNZ+YQCCBP+qhZEJxZfgIt8LyH3u5
H2OJuSJUBMbXd8wEHC6Q57L4pt6iQD+ya2qMPn8z3A2jzy6a+QcVLelLk6GsccCyRwnZRhuiDCLk
D6pU7Mwu/EWl4u2YsF6JkXqJaTlAMLkZ9yO2+5lZwl8hjJ3X92pRRXK8dgKTqSwwOc0/1aqDZ8Q6
ndIcuO/JKo3FjI6FyFUVZ5C26mrjYQJtyBjge9Tpr5qd9VaW8C3KpEDZ4cM0Uo+aB38PaX3kD2NL
maZFeTV2A88MGllXWtm2yH7kOAJ6VMZTZHDfKNAhn8Js2pi2WBeMFDA5DSfQFK3MInL4RrxSC76b
8/1dp+E1y26S9UWeFvPmZieL6v02IBW1YxVdj5y7W1bB1HQpMKAJ8EJziBIh3p2ynsKaI+z5G/rt
R+VQ/SkmC5COXmFhIM7WA+lVWbvod/Kotn3GTUi5wvIunjSUPX3AQ3NPx7PeFHEHRSJIHXYgHZxK
P7OG3CeMNuSHM0siMDOh3J8W7QNTWnLoBCJMukVJTc9o4X3BUPyXFJI81KO2kBEEFof9WcikxCNl
a672cEEGTl3mGn7FYSaklsG6vwPaeLdNWlc8vkN5gShgaAiiaynU4h/J/qMBscst+svL2ozVHQvo
QGgH1wO93PvMFR1CjNZSCwrj7rAwSQHbrhJhoIIr4NE21wQv40Xttsu6V2KEhfSREe25QA/icbdy
ozODK7q1c9ka2KhcR90+dOUfek27n2htQJhcxYLfEeM83T+DqmzXTFbn9+OHP4CvMUf87CTndtts
xQlHTYfPAGxG2N5/BQxzakuu6aHdS1z8c1UKkwAbBVBFgRdoljqAfy5PJDGNJKedhmUDUeCZ3c/e
697ig8qMj1wHK7+sFwbh5tEsVCa+LWslbFfuChcqgk8LvSxN3uBfbS4JP9qRCVCKT+iT13Zv854D
1LOcUyQGBKk/fDwu4z6loDA8JlTMV5YePSE/aWTUufIQVAD/RwZPTOVuFN1hL6E5GtbBvxVEewOB
zgdnxLYFdyldeb9Vzleoc09eg5WwNWANs0svvab/Ha8Z186+BUfbbp4eFjjVBoJgcQicH8ChHv/8
QY13chZ+dpqENh10gshCoEse0k9YXydhoGC0rLq2CVcqdlYoBRkV7y0GVF6rMDGLpi4qpEmzuuoH
YJqBoz3+ek6oyJE6EUCi+plb7+iVv3zrtyIEP3e+xi6Ybakkuzvx8h8EKo69JebrTU3bpHrfV/td
yn4hJ1nMJBEmNnOb1m7anCi5impZysxb3ZXppE+GsdhfeWMlI3aTFcLXqX46tUoDzNiSDQoUVV6T
hFHjD/Q2XUEy6PoX+veN/PxkrhvillU2bnPjOiexSPu45ftuogQe0xpugz/JjiA6LarLxt+F3lC9
uMSAzvgIt7wjl3LLM2GLACaeDmZteDyI0atCRUfgFE3oB23YbdQFNuYqo0agzVyUF1Sk3GIk8PN3
0S1hOQzWB1FDS+fVLDzC0iO9N6jUiTlBsMgcIbCA2AV0lFXmWuIkjf5vH2yd19ZRFjU6Gn9w7NMN
ckkULE1nIoSF/qqr/RcCv1pgWH8uw7MWoHhY+Tr2hIOxp+idBtJY4lHnT/+Mg1JJYiy+hNfYxQp3
9kXtAN3cTz0jP5unA/x+gTGYV2Oi8voU5RAQTKZSvMfIZw2EJRTuzSe8V2+oc/J9Vytxw4+rJC77
k5uijAUHf1QOc6STpaATAt0ZxnQEMaDwoSD3JnSLsrPaCXem16nyk72PO3F2BGY9tkv0LkTq4F4l
NpetPfDiSXBGgPW6Pq7+8LOCM5Di3V7cu+dlp5eigN4jr+7kVMETTKBE+vjRoVCsfmXTj5rr3i1b
YdZ5xw/9Om3SM+ln5jVM6swYdUP1AYlmHiN126Gyj3qdDxcPpAVtWMyjB1UPhbo+WJIl1YBSwpZ3
KBao1AS3v9PYiMPfKH6AWE9ESSjTKOwR7Ak9mlgMxcOj0TXKztd097SqbA4lxJSQFwqlk+9S6wRi
rXm7iQNisbMTTUYCEBAB1JVmRI1fkQZrPk1obF/0jw4lWOKqG5XS8hs31l/R33+MmY1wgjNuQ2qe
xq3vPpfJCnbEt2ySaty/3+KjRNRW7lsv+/+w9VTCrIb8oA4x9AsP4Tujg8fr+bbmatWufqOrU6aX
9jjHqR2km8MsvgXSMONVqtchqWrY5ezbCm8ISyRq/2Quom+bCIuqP1x//AZT6lUACZJnkQO8Rkmh
ZBK6KAjU2URJTZZbPnGV1CgF5LX4bRr78XA5ry9gkcSI3DvsRaWsc63XcLpqkmUFbexn+Y0WYHrx
EQnNRKYvBF7zwXm+TryVOyORYbDHcEuaMB0jrMYtAuZPtqQx2qrexAYPzDzQFm7x0uCXYsFsllrA
2L3d3T0TT1ukMTcaT7lod0K0idUFzlcYcPk3zABE6edb7a8YGEz0XQ+qK9GD8Y3crRddsEDOfcck
bfJGWK8KsvsoEZjpile2aIvB4GLT99Bdh05o+laH4zEXKaeeNz6K8tdwgxFtTWZ1fpJnTEr35vKy
W6BNCZi550E/OO2DT4ONoQE1KfxBWxyIVT4vMORZ18bu/sRABRla1mLte/T04xEC2KrclE75hblm
Xi8bZsV/a5PDXpubj/QtGKNrAjtzeJd6HXj76Lp0mudCrsfpa1+MYY6+QeuxQugyvLpdLOWqIz6N
pDYlMu73SRj0ljk6qdRi8x1Wy83lHN2Kc+NvvmwmJF6ZxNodBrNSakilCUIYoAy/4M/EHodYNgrQ
bTHBGSGLlX6H7pTCP+BvlrKAbfS5szX8gmz/wjw5Di3X3jOmjsMQgvoCamDOSKYrISoA6IPf+oav
DhD8HZk2Z5FXynpnZWw8u7/IOiqYbUG6BbGdGjmWDVk76y0DZ+iebiaIvLcfddFn2JnXyVroVX4/
1eQJXbWFhJmtC3wPl8TzMSRi69k0hnrjGc4pIrfN3lwZCI9uBU/yuA7euXCGWQUmIEOTeOECE/HP
Tw7YmYH/c3L9bkGxFB3ZS75IjpHfuBMjss9+JmEzCvAxrz/5Jrxxr7rCn31j/3ehym0ufLAx6btn
ax0eCIBz4d9OJWTpSyA9fkVKViKYo0JZhw4Nq/MXy7q1szf1rj1Jc4KCpYx/Qgo+tHMNZtD/SRK8
2KlsZJI8Ro2yIyfvts7gbavTMLtTF5kCHIbLiVa0M3fzxnYs9W7PnC5c5UjLj6jyLINVq5cnyKMn
65mMpFlHRJbY0nLXE8kNzWxFvW16t1OtHyKUT7YQaywkXh1syWqxG0uPRR73rylEHKUQTIqV4UMs
3q7t9DoBuGe2faY8m2cu631lCSBvrzAptjbgty2QUUhIoxWflZ3YXXXj3iCk53y007Rbims5WSGX
lF2P89OoUwSyfOpTGmV7DKZzzqWL7+III0ziBeAmvtor62rfQblL+XuVm1fSaBRXatE7JEA3N6Se
NV4a2t+VsmsOUvO9/EbBy8yuy0OBdaVH2FiYYcnV34SnvbMTO2G7NR4YcbiiB5DrPIxWGyd7KBPw
AvEwzeXZPrCHNA3VGShPUq5Q84+8lxhQ6YBLd4kxv6fIfNmKQ29+ouEi6dE+svC7gm+ejPSlU0tX
fg/tWmlw6adWnPlkTtQRQOAG+CDGTccfCH1ELtnfqjMmRqMzUI3/8evvpjqaKu0I9qt6CUKy0a25
ALCdhRtVSUzHHa/e50xmgxFwzSwQRKU56FiSwfoKvOXdgB5l2Jg5XqZ4fXe1JeajsE3pDOl1RRlR
F24jEQl2aNgXSjNJ1Xq/xQWzysWo4W58VBB5uqNM2i0VzTqFICZW2sfY5AuI+//jz3UqkXWs5Q5h
3JZ6qtlQYGfzRfAcf7dmxW3+lfPMksVioQgKVArWaVOutR/kONf5NQDNnyDYdruHBdxj3tHCmLFG
Fxx1elVwxYrnQMVxPZYVOAz6FdXyGBCkMdf6rL6qWw3GPj6aoFaQ5yFXvGWsdgaxOtDRzSlw/yKj
p8sJjb6p6aY/0FUePW0R0bCapX4A7r8vY51N33BR2hrMbfZ9dXDU5yF9HED3odXcoLS2kwIv7aa6
4uRtH9qMpi8EFemAERksUbKQ9/G0/nUlPNW6QcJzVDoDOCawE9r5JsjZfXIPGNz1znRhj/0+25Rm
YqV7Q6+QVldSsEoFo6LA+/HidcVZutIqbYz8MChNBPdBsGMtYIQR335H07Ry2/9U36aHmmtYiXGH
l9QWGxiTKx451JvIyITRiKt/s2a3SiedEMQjPNQgWd380Dz+pAd6LWYzuDxcq9BvnMydAgix/+O2
qMcoNSNfgdh2NBmz78jG40VYpjENel8DpJgNCNNSfozGEJBLW4QLfxCblcEVQFGiUWQ744rku3dI
wrD1kbpus3sJkJS/rSupReMOlUR738aMqSQ8jf1toRl1KJM7kFuE8aDJBdpipyo6tnm23CRTIxGz
IUEhSdgjAXOmdsfafSfzYWVi6bk91JBj/cS4On//vvHM/fvbKW7EGc4w3A4SJyPBXMdFtiRgevSC
VOR4VPISdHEkEwIaMS66cO1+fW/sWxsfl3GkTosYNx4B2xI3TZiqZmVLSsQ+h1hP6vYv/IHwi77O
CVJrJUkFGroWwzMxrduRErsv5ckM8jWeTLu9xevAGJXUApkT45kgziYeHcAHFA/CQ9KRWoiXF+S3
rXBPBQFav6EvvMfJs1nsoZHoQSYZqos0d5wB+Xb/DW02G6o4P1yDzNv7ExqplUeqv0H+5xWQhZCg
uUOW63Hm2RmoaTbKPt/uL+G7VfLakC6jmA5rscVFV4LsWpquKpebHFdsQIsIhWWQRz2tK3sPfXoi
n1De+H8HeaSLr2IcxyaqH7VMLC2jkTNBQCbKywo07PI7JBhvGjXITTDOsLSkWduKEa3Z7q3KoaMP
NrpStkix1hmq9UncdS0BhZdaqol06rMcxhxaO6aX97U2P/chhA8ZOIWReh5nhE8WuoxUj5B8LyTA
y5ovR09zK8F9B5Ydw7dxt5yzpuKZNY0la+dC4QufCDx2AIcymPsxTkBmzv3NoBuu3e4EJyXwhzXz
57WAaeLzT6Tfe/Gc1yShbvq12Dyo1wi/geZ+Vj78r8TvE1bL+YDSkCrEmiuo4zhEdVgMgiOKvTKf
xfsQdrcBCXLYx/Vkh2q4JYw058Y6MaG2MWMF2aOcQspjhaZQrNzD4migHs3PaC9ECg8t00Wmsc9g
Y1KSscffZyVzPYLOCyH26NbW/XJNGY5qVnkhjOR8c/SOLZUAAIGJh2HWQeUBvveLxaO6K0gaxN34
1M/gOHreLmrnO2WYaI0VHnn/fwmTCjK3O7K9HeJnTbrevTKZ7lntE65rzrShJa3/p2/8NL54CUvg
nfvXkr030uAuzSS9/P8j0WlC0fVX/rInmJMo9Ysf3Q/WGC8gAiz4vDDY+uqZ6aCs6XQ3Z0mAuPxh
qwGIaaDbg3abw5aYaMXDvslDqVSQm7ePtXBZrIChx4GRn1+6PJJngwv+itFBfDSHt01hzVTjWFkI
3G/ybh+d8vluvvxuqA3qeBhqYrSi0qNMhw1t89RzE1Ek3INK4mYjFF3e4dv6TK2/jDMjhzcVLCjU
L6LynGAT5cYa1wi7axDq5Ylf/cVpzx/hsO9y2nl6yve60UKlOE7g9NvBPp+29yIBCIXKziLoFluN
i5PSdVDjBc9SLe9FOvwo1CRfUFxLl2WVvY2JWQJlFNnJ9qG5cPZ62ke78zIbnPbA0HZSzHT7ZRLv
HUInqulwYLnn7c9/zEuP1/gJSV2ofAbKb4fZybceF9RU10SrZaO2S5nR8LJaEr/UqeVnDO6VQpsT
6H5GPKMkT72j/NnEDKfaQuDdGGiahDq6M8P6zclsjwDO7gfqMQ5WD/ld/iB0X6QgH4tky1mddo+b
vXElCM2mGS8pchd8e65KC2HZkvr7L6tnFapo/hpG5LBdoGGvL9LHQmCqZoSen/s7YzCIqLmhb54y
klzre3rkmC7eyBznT/SBJtJ+rEme8SMk3pooFJCdkjqBTKz66akRi496tXEB7K3FoUAuuRvTixEo
Q3viu4aacAjxgR5NPKeDOuctxEiTRvV8Wn3AJzaH9xCTZe5mD6Jj9cEXhpgqWP1fLRLEd83z+FnM
Bsx+wC6D6OasDgpc0hqZOrZ6E0ipVg+F/Vs4aLdWFphDW9BmjaETlJXvnM0m1YMpbNe5DJXgFar9
VWHNtHAo+Iy8cx9Hxl+KKmyhzeO30Tjh2cYrhijnUCf0MuQctCbXyUGwV7391zAqQ8BwaVEqYfxE
OooTvw86Ff+tq0P/uDg4AvRhxe8mBkIE7sqduMOZ9vWhsRa4Hys/VzidX7tk7IbFHPf/D7FqgXQ2
hgs55eUJPZLllTFShjZTwZN5eTwGiUC0lcNSm+OsTRUnvEAk9ZVqLiHr6bkrbLKTLSZS/yxhP1s5
FCZsv9S4+22CLbXG0zMtYP5cqSMVowR/RGtii94sjpXF+0jN0/ucuDnnJ3ZNhZ4puYGXSt9CF8qn
wN0XS2MNoa4Fa9nGZvjGvWvf14i3ehUCQoLkbvQKsoQC1PbHQCQKzDqYFvHc2n5Khfzzz1M9y9FX
vzu0s2vDmiasLttQdNbwepPi9WcuEVsKRB4a0mtDrsXU9AGSO6PDwXCjZaZva0tl/ssWF5dIAO55
55nw8XxK7Zh5zvM4wKDl+B9iLYL6+3JvmlEp8rzRZzbPmq+0AyTPahlNkUNcpLbIW3JfVageMojJ
AVkqoTtBmYqTgBHmTHxf9lzl8trNIRPEiZBUGF4+taJqlPofWTdlptSHDEsPO4z1WDYdIIXmjl7E
b38ZURFxkTvAup4C/iLNrSM8Rj1qfE/EgF8QdVH5O0w/i1ZKdFWnziSUq2MOcqZLdREBNsiTh4yW
GtuAVyd4n7Rz1eQQFwXBuKAgYjmYz32LjZWYPi2uXmW7dqYENk54rN49ZRZTGhvZjkYgJdJLJhSD
+Zt2lz7SQ61sEPNha1l7WAMEdJHE2hgR2pqYH3XoLVA2pHC6/ay8U11wqN0yd9xfaPFq29x5t8No
MVwj+fFbmAL1iy/KU1QOW0UjSNQf6fIf+3dZRgNdk4MB2jijY5g9CaWGIPMtRJ4msNKr6S6dEzeG
GxMyp+qTcbKRzS1m3Ccn/PheIt0BzSF0pCLXvlXN5aXkBwtiEBWt9i8k4cTkilIo6sYY+mzKG726
a+x0Z5+okzwy4cJ2FL1jN3Z7EC6Y/A/LryEAEgzo79oCgyYcyzJC3W4X0CZIP6ULBoQ3ecRr75kK
J0vTuXaL30g4/2CVD+S111KPuZ47J29WCAYwYM7Emmq6ewwFWL83eQV8Ebcr8F+N6r8xVLQoBkSg
QHUqlPeQTe9DViVknHhsOkEYgw1GPvshco93BptaM+U7zYlGh30+Ar6fDnHbOBMH8jxeVRRWMuCi
srvIbwlKVWv8aNVLchQNQchjCct57hd1Zcf2qqef6iPYgCT2EBD5fR28bLIfGOx/bQkqkNF/dhOz
fv9cXs5b6bp1GbX9ET+g4i0MbDJe721HpIJroRyhygiF2dlbegPTnBmk+Iaxj89hVj932DUz9rQk
87BwhG1wi3UaEoZy8bKP37tW86K/yXIX3fX7xVKs4XkXzAoL3JBfv4pYDC0aegyIfyKBXCb0Cb4+
3c1uM4CStI5QhnFLPza5XU/KUaHMcJdkm63BqrIzKb0KNUNRbgwwFZGEUZUwrptjcItHNs8op0Rb
JW0A5OanGFp0bfaAiDyi8p7C7RZ31xXueeSbYX448prLq/IiWKZRy+KvEXgpknGAN+kj8lXLbUsC
cIOz3XC8FNVqcPnGUtpickd3Z7PTBQZe6ghOSVH5MRoMKiN6gRxYRyE8oKxDP8TB0YUEYetcanHB
crSp7RvE/kKqjYISFQN9FYdiaPC366Ij0nqr9Hj9feBzIEXM5CPwjQkjag166oidhzWnELMMkmD/
valzfaA1np89bMosG6aZGMfiRPRWqx3wnSurTO7sUAf8PkYl3r0LvPomOYjT4l7tQKguDnZcBtOg
iSkY7BRy8k2ONp6PmGTB3M0mWvIrKoWG4RJIaV+M65QnqY9qJJu+XeJf5LXM9JLxsSjgCzef1vw3
f23LxJTyHGv4PGq+n+Qls349BKVhW8argN+AqkouoX6aJjj8Ad6wPCuGkTlqmSPXxbUG9ahYGE9U
X8pv1wiRteelJ32XpXVqDahub3CwoEBcY11xw8/DG9+VPSERMtkY0p1Lsr9jH/59YbNLuaYRJ/s0
mqrpZDiSpc3k7dSk820MfMHQX3hHFZsGOaKb96/kwzzpRtKdjJ7QreLVFRkJFf/xCp2yWuzeOEBH
VNbJpeToa/5joBDw/C6WjBDXgP1iO3eOSDgSPaUt00rrC3yvKn9eJwe4PU8K5QCVZmE9VDvIOE+w
s8E8FzV8brS5C06DtXnAYSvMtr8LBCwCRS2WDdNMYij3xQrVodXFxmaJAwxSsIOnZCqpI9jDOvJI
z602rOMIcA4me1AdK4hXmaA9w15R5/IhV5RYEFyNjepu9M5N3LZyqPkF2/0WPgy+F2S5EfCevNIg
BzC1TAhOHS8vchpv0k8iaafCFmKbUe0pQwX6JPr/pfs7sdbfWne044Ki9cdJhMlHbXn3FyKlZarw
ruS3yrusrz/G8ZaY+rvSBU5CJBNkDi2ZLctMaKDxl3wQX6HTwP7ycS1KG5mkEv7y2Clnj+Vf6b8s
kmVpIO0z1elFz3udp5d+Gaw7IlD1tdS6NCXnghOl45EbcxW2Shhd6i+Hs7vs4ptyMzZPlL84rYCR
z84o9RrjQF379g9ZI8z4w+DjmBZJR8NgnbmW01aPsMd1sIZitjndlQJnxvquHJ5Vr9nkjOf+uhNy
pncVh36nkflCsk+mW9p7q/N6oTJz3UrUbB8KLzKFAWIPbOWNOwC/+31IC7qVyiPLAZvfAi7elMhs
cQx0fKSUhcTXCkgj2iK6Dzl0ebr1pYSnUjIxYKYV2heOaHfybDopi+gf7Khy/QFhD1eV4+yAiPzZ
uotUvBir8okvUFibZfSgnDkty9/zIW/czJvwfSjLQwq02EsJNQVhijmiIZ6FxxFnwgERp4wqQQdj
F5GTYQNzlJgQp65FIcG61MDmYfiYWlSswAslz23y+inw70xATCaSGlGmNLsuQWW8PvEflt6VvRnM
r5pU/Nx1bfrvUxFgXo9WTPjjVnViyPugeUJFn8Qcn/kOPXFyyEEgIAa7IzwdHstutoZ9LYvOzRAW
wDH/YLvGITXaGq1YjqUGH+urnOcIJynb1GwFIBTnujAVSNBa3FaMQbrPBBw4mU29Vbi9Dpf01jI8
BuAGLiIP4Tr+Rs8cnbUuEX7upU8GPq+wTl/YoOupmN5/w+QKnurmN5nqOTsiFXMwNadjz0HoJflP
SaCsfMT6alliAiCPqkqTb2/fuSwilOhheQkXLb7K7H9q4EPbmdyTjMSKpmZqXxe5L9uf3lfeBROP
NFxmKiPvlqcgA087uAUF8958yMp//AheRE4VDqIMnvTquJbSTAvlXKyzZT67LEMfd7zhksyACbaL
Qru2wIFcPDOV0iiwh9glpr6mlITrDLDCnPuTwqnmrRXB6ACn6u9oN/LvgUVT1FONyJBVCOMOVzBl
roRNTJ51UrrEYl5F6cNzLAYKxV8bMdoLNo/OVyd3XuABzZk+f547oYYIDtSLgKf217ITKoTeBYGg
ftRN4EHRsPCtncIZw865VZ0ge6QsSdXprvkQVj205EvBjLdcDuvA+WDr3cmJAQcQAxcHkPJu95UK
vbHg1EXSQvg+dK33w9DxXHewiEbs0SRyXTQMEGEs4gV8UfO5huefVls15+EDVc0cJ0LDJv0Dllfp
D5fbVG7eI7hkFDetKcplT60Muy6uuaANA/Mi0fRFSBex1ZeJA6rAQxzXFILjhMIbMCvRxKBgsV+C
lG7bHB58W8jhe5mTiqclu9EPXjIVed0mCyHqKhCGfp40+D0ORcXXCrpNnLhJ2UlZC2WWdluEBhQV
HrAdTq0B4n0reOkI0MFmFcyT3ysqDQ1BX34IsZ4paTtlOOiK9DWDyEY8spWrj7h8lrOeTqlU/Atg
HgEwnAuOdOTMi2S49Nh6uGOF243gO5YLFwxgf9WZZTentCKXJDN9WFEy7c7HdAW/CyOgt5CXlhl4
0uwjSfAR7JeGfFtDBj9uvuBRuxdGGJVymDTocb430OAQOkOMY+VzIRgnVkT1MEs/dudccCsvSXiJ
RmakSu9OJxG+Hsb4HamQ2lBYesA9hmDlOgfw4pPab2gzMZSYlzfR8F+4OyfYKEouIRbw8srF9JE8
7Q1+AumOntoHvUOp1p6fnOy0tM7+IC2yrcg3euI/V4nH8NNJAZrEt3sQUiglTulIXx0EQstE2pLa
0PXgXSySGgRN9pz1LC3HdEzYbDwRgKQTI1QMpPY9g/n/rMu5j62GX6I6YFQPMhxuw+ma0DEjuJd0
5u3ITGWpSP/SLx4NJ17MU2jWibztWQoRrZYpePMZxNGUP9eC3bv4a1NSElpov3mIYS2B9xStMZ0u
ioO8QSAZZMg1V9ZxmP2ZOOuTQ4RRWQ5xLA1Pt/g5DMyKPeMP8LQwJ/imxitczfMyyPjIHQ3cshBS
C1LylkyOzQoc7VmmB8/tgzFcPMdAmIX/PhSWQhnNxsn0h+WT/Jpg/9agA9qVkeXteh6fKqNy21Wp
wjB0hPEnupHl9Pn6n5EEf0xgxg7dCEKC8qhuarsM5XTcq6ju3KzGtVAeXvu6qq0X9rscreWfo1an
ZiER9NQZme3ZigDDBGPSc/DzrpFfemhz2068FUXOt5FdnFPxeQEq3cS1gHpLjqWG+0IfEeas7Tnx
yDcMMRY8G98/9hI+TTDyXOJJ4xxZkHByoPYtRAUQ1lI+1II5vBmhEH02gpNgwg4GkHIcSJQNpy4O
IW+Arbfw4+TxrFpm4WfB3ISK4QlSlrAfNTOfDhnDwK0ZKhoEGMBtgfgraI8Agok4eR6SZQf7JS6x
C9npb2sp3tCUrgn3KRhKDTjzkjsSxZCdqsFxbeXgqvQ8Mg9j9T7MBgaz3Bh5pPmCq0/SEKt6gbvS
dzTE41xPzb82xpmnQEiB/RwhFlOkoYLh3kMJzFIMgLQGu6FDR7u8MJunwqMgzvSThBiAFjKrC8vc
3lvKoakcWl+nrTnMN1k1gm97o2I9OyOHny5zQwUsnHrU9cIEiHFhA1+THLo2apO+gP/A/iRBkFpe
YTpudxfCwkgnGXTYSbLZ9e239ch9o5y3sDgWWAhV+H9e87TuzWoUNci02yIbFDRGyIADMn1qxyLh
b1qfzqCy5ynUg+RFnSR8H0vhXdhY3OSo0dXaDs0PDwh1qG1ijTWgzDwDJkJo7YEj04xrV2F//Zsn
l8ES9YGI7XvBFFOVZOjoYyLegyahLduApEjzkOybL5+WyfgekPlD/EAPnBMPy3yJLmAn6NeSLTgy
j4xI1fINiv20DLl6b1Izuv7x/5R/34S92l54E0xxUqdAggPhf3h66SDPC/lKUtOkATIn9QX4ty+m
PrZxVeSOFTKYyc6mnSVoJS66cajN7mCQiSr7yZG367ngIxoYBs9iKGBGRD7f5iio2JnB5BWHdPaS
ss2pjmxIKnIsvQnbMjrnzW+F9kVBN5pb+fXiWwdeOHT33bjYSLQkVIn12gH+xtlEy5fcvklhbrvz
cMAfCyb8I7Yq9Atxjns3jUVzViPq6V1MgzESCujMEcAg819kHilOqj9nvFTBTNoVIpP+36hDvoSH
fmLDZWUGspEuuI5abuIulZwKJULV0QferuTV1IiTGuzIzf8lUU7LXXbCGZCGmgDuV159C32aRihW
j4pCnjicbpeNussR5SFoRGc+oNnE57i8gDfMSWmFK9kWJ+lHjGCwYqWJizmcClUyttE0g1mMQje3
05qpsA73gvB1UYgsbZBs7539I01BrG1jg3qdCJY7djwLt43Oa3y5vjPN7CKUCc6+jJsd0pCyC+Dk
3iBFpMuL2bXKftaQ4ryXeCkr3bu1J0Y6FFSJ9yattjUZWnDd/sy3ncx1bcXw0dmcEOIdmBVDtc9h
VyNtZ5F+nqyskv8bzDJJ922hncmwoQ8+g4vHDxOoLkTP2hu9fkCqmf157DNuZ3vJlfAD3wA3PLnI
tjBGrcVs9dJe0CzSdhGf6Z17E0+iEGTNsakZLeMgPT614SErWDArdhM/Vvn4jQBNcruUDfsfZJs2
pVDMcm1LByVwdcvuGlkCydP8JBfREdyp9btDml/hEF9TPGgeDsansWY0S6pJrvjZYXXxcLN+KIGu
5Xc0hRpeu5YPYyvjIZqtuPQCeCvWHbAJwXbU1tAZ5ZaEhbBa+5CouzGBZOTgt0I6bonGFFzh2lJb
/denya5h2JWyzPf/ZjxnOgq7KiTz+v+AtRKqEGBloUXumfGAoLDwMEwbHG9hXiI5xwhq3iD1Oz78
VHzJXde6TIgvtFCKoPqXBF8/iTGnO89Qmgw4114VdTjilzeLEkmbUZc4ZTajG7N136/NvtxFl0h6
GJUt+r1AQZk6RDl1OqG+AcXK9hfGaSeFtI50ILIMBkfexqzErUWXD+nwYEJ1VD2JvD51Wla98ums
Iggws9PFyyg2uUMpuKk61c7y2Udj7mEnLcDMxqI1VYvXEQoET9sukHOSi1p8LLYvgXBHNCUKVCWG
ws+wH1QWWuarOR5orktCiYVgQnOme6h1WnJHC8t5F0z4/XUqqPoJN75NttVo5waHXLEk/+nkg64F
1he6CFZY68q8I1SghVs0ccXXhRFbIN4TrUrC/ViXk270S7wtpu7ou4ezYE5vkWuTQOfRwOcop5an
+AgSU83GN+g53qRPiveih24iUrKWo5U4Zp+Z2vg3ZOquWRrJl2NqkoDtJvcK4r95+qfsMcnxGcDa
MqaEadaarp05DZ9tx6J23dqKw+5AmtIgIlEQE5kbUKF5/gbHfQjT6pd7O8O8I3hap/wdl/WIp0fd
Ppo9XGWAtCTrSwO3PVgnpZpnqLIG1b8e56riXrzg/OZLFY22Wn/f0h+oKFzxyF+a/A7Oc8D9Zxxr
+nfSKGPRCP/URqO8ifpWGfW6uHh/Hahr3cFnxIvLMO7R1JwGQ+mr2hF8V4X7ONJD5rwMhyFx1Mk5
mQbX8EWGC/HA9HjlMQdrUtKPGNtzpiIE+tC3bv7RfnKiPgs05Np0asf+7LbU46BhcclOTYz9zH+y
lKeILAcCI8C+pgbVPpVLzLyk9W1zv9HfKzi9ioNn1uKPajgE5McOq0UoO4EPjeqxNpdctbPH0o9B
FA3OJ3IHDp6hN3Ywjpx9XERVAwR09m3gso9we0ZAtINWDCnN6iTYIQaH7EDiUjaZ/Ia//NEsvq4O
Bq9hN2KiDWppDt4jOL6s3KduEvzy9a51J/YKuHHscAS6+nWcyuGCpZEGy+/oQob2Ne4jHeq04zwA
GTtWc/TMnB/xasvj5KSoZc8RzQTCfufxM5o6xbYeaCUnNh3b/PlFrk4kDRHRQ4dbGOTQtYvsqrGE
rPhRUcuGZN/CSLb8CSQssnxjFRMT0FsRtc96b+SJ0UcVkOHLd11OOxVb9sAj5qG0PPlfhKejlGsH
Y3x2qJW/PsQ1pifupMd4M3JMbLP05oCO/bAYO74TTJiOaEGlYGlTpejt/4oprr4GIxD8svtBsAON
BoWUyn/PFmTYRIOVbv+KLC9zK74qsc3Uvy6QR13H//5IRlrmDc1/9hy4yEgoYFjvFkBP2VhK28RS
lqelPDmBIX1yl5LcQvtNYjYGLTFI3FXfmUvdE/oW7gHkzbBJ9z73KH4V6zp64+5qNtjI2bf7vf6B
GJSghBmzCv/XbJ+zHc4o6fJbUWVeowHZStt3Ey8HBkAByfqVmJs+5XrKFL+5/enBoC04hYekdWHZ
oF4b+YsKH+kzvL0DC2dzEzyWCXJ8F4JH2B4vCobeWej6J4peBJLiSYC5dLejRd/JMU8KUH84NTGe
zuovdUKJf+gPhWuT89qx6dCiBQqZVoKTUY5n6oJYYNjSnBm90Mrx6/VAJ3JqkyLhSFRKsiZDMf8u
NpQHNMAOe7kr8RNz1WUoeHu6awny5YbLV5SixEl4iyvCR7F6iSW/Wqr1Ojr6klLkyvdoS7MOcr3b
BKeVtMowLuA+ugsHebB+DBNdJbyZVVLOiEKMA0UrA9CaHD9483ISZL1shEamewCnQLDol/NcPaMo
aQ1Qxh1na8X0oYwUf8Z/iXzUFG2tWuz6UfVUYWF8U1ULpVteOfUu0sd+hIUBOj0AM8iaW2KseKth
cuHvyZ5e2EN0lxvlqHK9Wdk7mv7QLKsCh42phlHcVP1s0+7l0/3e1eix163ngieGfrWehD66QLvG
rxNMq3+GAK9cVSQ30fu8eY5+nyiXF+xGxYxLqh+ihTEKZAHus9jdhOJhaZuNFVQvrxhaCIWNsQTH
98vi+AUVJQ1/W0B7gXAL2pv0sKifRGAo49EY0rqHGmKLJcLw4s70yFsjnKA1rH5t9DAoMMFNYbHA
Gcw3UZ1LoVFKcGHE9oHb2MTQUBkYIfpoUV5kPfMUVPwU1w4dSmpbbhbeb5baiS4a6Y+uF1n/CsKZ
oSBSzxyOFZXAhGmv+0QzpS4wz3c3y7CX+tetBscUYcueiNLwhg3vNtG0QfXXNQVjGcRQNnWPJv4r
IidofvecmICEGbOLhJJknVnzmRFTULMX/NMttjKSL5l6gGRtd1JmV5B/VgxeB4rjWOatapTSbuOt
6UvFSYpzP+20WUt6yPHs4FjrcUX4giSdPuA17qG00rNayfxl2xMLK33rEOk6pi8//By6ndacN2kb
YvLkf605Wi2zOVFY6/TbU20PWma5zPy2YtODKnj0rNtCazJeejo04oNQ9A04cBYGXh6AlJ47cPg9
R5l4TkToxLuN0UE3q/RpbZX8eeglF9K7vSHaSqHWP+pMHxOyu4d99dDDcQdE7MbfZdnBlJzjRGXJ
nIU2wDc5pbDL3b4/q21/11cvi5mpv+0BvD6dvohUoTj1htzeTXbWmQj/22V9WBowiu2xsidwsPJO
I5Q4tR6ux5eBibQ4xzn5os1G1QScYkTObP8FYf/KGGTeJwRNAb2V25TbbRMzkAGY7hk4p+9/GCBN
QcT8rV4WagxeMhN2nDYei0InkJ1a4l1n2SN8tvtL0/MVIjM3fIa+vs8RfhcTPDoyATrtFmWePipG
OcBUF0w9BGg+1vGj/c4MZRK2UxLwpYcJvXSRX2UYquhJvw4Lh1xxYfiliMHPWee7/pcEb0TK5LS+
yhd1QCv4aSJPEYEsN9Wvk5NnVXVNm8Ersrt7Cty5EZMdVo3iGeb+CIjJzLLjB1zEwWzakDyfVa0Z
NMAoQEam+EbBsmpG73zKHUs2nXwf5xKrngGbNwpgWcmpPIoujSw87TsTPUE4O0J1EghCm6SZQA+M
sA9wPSwKieUBh4UUdbZZJQRHEZJP5m0j4IhDOJSbw7wmklfzHVAjcDYTkXn0Wh2Ykajqzae+N6gy
hxDCYNomIpWfCw3IM/Jbr5NTQabI3f2B5H0vT0ie35jAaHAdjay9B5W3LXDj0Ot8Sl/CDHVuvOZQ
7ZuwNCFc8yQby0VM3lN35W7h0B/IYxUitYEsKTnkdCHfHU4VZt1k/bKCKnSzlbd51qD9EAhMB2gp
+yktMpLWQHFRFVM6P+rXbmMsZ2FDFzgdFb2wsdau2llfrNv5Ys/Rng10gX0fvH9gA1JeOGPX0rre
570i5sfvCow2cqRNrGSQySWblurho2VRR/VksFNBuwbx8Tm4jnsrpuyGRi/2ZiNLAD1eRi8tW3/k
osF4Y8zPPvALztdZiau39wd2B7pAr5IFPz+ZN9lzwIpvSmJziZSQHSr0/Qdzus9OE5Hh+Nh46CSx
q2tahNkfxqjtdLe52MOd3AtfpaTPCoajH1Gn5QlJuh6obCDa2UZzAg1eYsgbHLuNrgbUe7g1QqtA
qkwhx2Nh1X2PTBLOMrHjZiTyPwqD9Mm+alH2BoXicecIUlMCXXGaWrJqxe6KHYJTBrP7iXM6B2Eq
xDZefYq7eIkHbGlNxhJQILSLaGGo41SlVDQmehBL0qNEYCxfNb0Lzevi3KbhM5Ts7WZGb5BIOZAU
jrcgU+NlY1JCPIC9LE0sxTzB1tzFTgdDjidzw9Z23mhRz1YPxeUsvVROJVQeQKOjoGJuUri8A0W/
bSm0lHLCPIYS8jFSmc5B5AZaC5ZoQjSGB7D2uJzy4ZQMkL/dqXaTeMX8IIqSWAX/JYnxFtQPwpLs
UDy3n93k4qQJE5YjpD94vrZXluT00PZ3I3IqkWhoMfT57dIejBszkPU5KM/laBFZT8bN/aKJguBU
4IrjvKZJPRh4O1UoRnW09B/cb8QFgY2f9k5WIJ8Rv2mibCXdyWq1Gq65Gd8yhvDnNWffZd2dnvRq
2jpqdY1Uv+/mJUyZej4GJRLWO8wMErd7O+K7hM/2W3YOeezfYZZG6diWjAobCDiZympWWHPfTm86
nHYIQE2xJxYroZ5VB8avDYlkKLTjX4b0zyD6MWsZGnxpn0DhF0QYcEiVxuQ+Gu/ZxDRXDGOQXHbj
vdNs3wgQlxSs8kaVZw3IVasDbaKzYoqsgiV6Gg7bMNWZJU3RBZuuhQrwv/IJ7BwvC4T92F4SMIWS
DjnVGUHfyinZL4ltLTqpNYQI/Kgnfy119wVXaNfJLG6Sm5OAF5LZXDcurK+QucnF+8DljCtKZeft
+I/qi24jFbIUO+wSUHj0Ci4Bh3Ew3RwROaLHL7bBhIgi8YU3yc+MDuzGwjULtJxRsONC5S+XQg5U
tXy0fvhjB2aoyMv5MRPg/HD3c0TYSnO1HGZGZK5PfmwKW+VyCs16A8EaVrfpfeaIsdae2DnZ3v66
FfWERqKupNFgkz+8o16LputBSElmdznzS3X3zbaepsFKr09Uef4sd2871865FLyNCkvYAxRNeK4d
sO03dByXjJGCNsXcgUydgwOo3wBeI6FJ53+cAsVREvITYWLzdazmaxM5VSsh1Te2L7WHKlScvizK
crNDBbiEjKhoqxSP3VN2meeWnpkjzqDZj2iBxSuBek7SobJf/JF4dh5eRR2chLG/qJkNuN9ov4uk
NZecBMx148cZ3znT5bDKZkfoUzbc+jLXlSMy5boE3vOiBJCW5TqFkBgm6xR2lNG0mrpddwYuXA4o
zLQCwXqj4Vv4Lljg8G8KjQRLoxl+PO5q7jIj6SQVWJi4bAFSnCWkrgPQFsY5N2y4gRN/R1y2rkZZ
BUZjRlNfg4wst8eGFHI+pLm+rgu5RfhpuN/+0Rb5LonjfDPCUXf3hxa6+rxhM39uyo5F+sS/B9Nk
27UvQx9qPBHAjOy5KgGQqI01Bq+wPlg7akNsgd0xoEL06pZtaiBrRZ/UxMLKsAQ0hteTek84yfLM
2h4SQVKYy94h9ye5FwU2nuHD5jgEPtvATvDbjHNCxGZ4UvQlvXREMl7YKi1nRk+c/0LsaMTnf40F
61USn9bI+29dyicUSIB5AdkbeUINO8G4vTRYutMuz72SSV51gmExy7mmQGdnrw0+qpNuvXG4BpOD
oQWfNqzhzvQzZvVLlfaRlVitXROy4fF01pSJTZrVGl2xn2yasKXCKhFCJHCi0TCpbtcPmqYx7ZFR
UfwGlsFkJBiIZaOEXyphMXF8bv6dRTA1nmdWgYks4fvSrKoaUAmNA6bcMkEh9kD3tT++W0JUixNC
PtVCk2XbNHYxbhsZpi6CRlKOQy8BwOQuPd55suvcRa90uDSKyIJtyJ4ON/txVpR6f4MqK8pBE6Ki
9HJLJ3eQLb9nAzgR0L2plILsFKxWEJev6v6kQEWEtA/BWNhhU5e37eAs/Sa4Hc+/Zo6lb9zfjTah
aG18Es+IHtFMjwlTVNa/C+90ZNk0bgWCjbW7gfyQzuq7ScPgfdATu54Ze1W6nV8+oEFyj6tdKhte
vGRpJIOctlF551Di6mstshF0HlztmXBA5XeQKtCew0Q2Tnfx9WRZd/ugXcRor+cdAFi/m056/B1S
Xssi+04OG5Ib4vdq54F+51W2yJInUkjz9/v2wpE1SP6R5dc9OryXHEFSZYLg2NA2pL7VmOL7nSQE
5J7p3TgeJkWBcEwmauFyuJwbGvfekqGhuLiM/zgfNwAhqhW5FxhpXy06JaW3veKN74t8p+2Y5FsP
RJZKoZOFcalm1tXTtWp6RPYM517u2+pvUzuz0iHWZ55Wx2XZpm20ibkv4Xg6/aEiJpKlyCcAzfCg
otj4xx3hTvsdRfJ9LbcaEyJBJahgQCw8KqrUSRTHl8lYyocYswmnf8VimgWfgZQJN9iaToLlbOpx
zMwKX04Bu0VluO8i/VFOsoQA23Y6pWkFORrMXZS9qM6p5vLgiI1+ycreI6/3DgLV/JmQtRWTh2Ft
uAFzqRR8e4+ItTh35KQahFIQB7JTRQ4mzL8/8ZpFPP0A9vDKUevd1Ief63wu2I7W2yj8FGRYh3dp
1WxVCFz9wYjTzUdGxcoTFTOzEpOwUOrj+BEFOp6egCDML85qj+vDQhXARgYa1sULnq8HIo3mAQZ6
UgzaXrw+S+RRdKv1RfF5oWMMXjOqw3FyIzSbrqqri+wGjL9xlE6wqF9EDn/o6Q3M+U9aELq1RM8I
7ojrjmszZjfRBO7L+NU5yFpSzEtVWitLSgR4NyPTV4pC0TPXi+57GQpSFdvb6D40nDjr+eE/pX86
o7AhzDRypG7tHQSo5Td+mUjU67lOKpDT4kZvrm0EHBcachgWD9TESROKpXJL2VaCQcYWGVRk7GQU
IMF6jaNCo9cIJ5f92nr7tJM3eVknOOQRbqhOgP6YbQoVz2aCUbeyQCVNtY9NibosyZRqbgb0x54L
QHStmz2Tor/Wej5bceNnhqqtn5z4H+B9xfqzrwZC3Tg4Y0cQJwx7wRSB9pKa/FXdRMWfs0miT1Kn
LJ3R79lINHXsOTJHGANCq/K82Z7Zij7+wwarXZ+7rVxHpd6tZijMIkW8uCJvQUBUoaCZnpPt+VlL
1jGqeXzIm/3/kppauFQufJUS/vmFUJz38OSekMHxa+drdIrwOjUsEE6pw0twzkkPFeR7Z5k72xOr
PR4GLOmRO1ofxaK7/jWzRqdCKrBnMIfEhbk38W+hwIuO83PyCHl81qspigc/VQANqBt2y+NzK2lw
EIJO0wzqzbuOVm1GVRnJoT3bnv7eSAtTh8mR+yN80+l66Qk6DhUkgvCNG313Vil0vUhLwXtGIVJA
fTNaqygZbBFLBxJRUKBgGe43/aWNt5iEkjcZtZkSjTFKttXP/DI8k/lmmOM0q+ZgHCZ14EedZ0pc
OBmXlkBrTjPx/KkkZYAVi/iQYi+/AgkiTHBhasT+0N2DhXOPBZIPJi4izk+aBjEGAwjs49VDb+pg
tgH67pMP/v+p5w1XeTlV+MjXaJqzPDx7SDjHQgPCP39YYviurh0ia2uJR56c+jJLW9DWSan314TJ
fVg13jjJA1jTu58f/7ahM8IJ8OdiF3V18glHmAylQDYLbhDW3oYurSw2ufNtNm4Em5rmA9Wd63yf
uIpAwXDwvj9JQoIY8ZDj8HrRT3kh9eCVxSdEF5i/GwuzIuXuuoTMlwnQAqhYDCrTJWcvO5VU/8hb
1uJCcKkWI5AdbAs95jtwRrnN7BVAIqGJdTvqG3QNm3CXHC+tUPzrKaktgpWKOHMwfQKyYsgMlnFH
IAviRwpw7WugthTCDS3gZs1YtYhFuyfGk3EUcIWyDJN2hoCmVlT/NBVVfEqteAXHlEuzMTF/9nb0
Bxy6N7Oc81QS5bMxSELWiXbydlEInL6YQxCH+Eu3Rv0aJV5HG9aaCFNWDMr9HVp9ps8dn0N9EjS4
Uvc1ftWp2h1kH/Dh5eVhWXw50E+eTDf6OvDf+xUFqlzHMQw/8GxMzp0xOJrkJvm2MaMVWnej9eVl
wLt5oC4z7y2fV/iAkSgtuxICvUFfbFply7jHkJJSYD6gPk1TQKdLYuNDgZB37a2mx+D/kCqxqS4a
u3zVBFoYSszq+A2zArdL87QgC+fOnyd79072VkC/RlMVHQYcfwMyvtsaE5fNm5tYPlXMsVZ2cyx0
hmcdiPYPkwN3ITQWv8qXPvC1P0jifWh02Vjg+8X51J9u/ufk1Y/2fkcsqZuBeeLtZposRhSUlq/Q
0+Atcrq4B9EpDSsrNRC5u89WDRVhDkdZeagfQor8tzeaCPMg2y1K5T76YJoqqERJIwDxWmX+uDnh
1HSraBWm/Aob73spInAmXJcMnPp67G+ishU4CvmIh5s2XgL1MyaoroxBz1OMbJjSZz6vw8pGeUQu
2eTaI4edy8cOajH41Pn+UesdB7whiapkpbkqRPozBBB9hWdXlc35qw5DNfqUiLAz6FNXQU+1vbz5
EUCIXkZTdpkIXngjU/zGLHYrJ9mUiFA8xv5ZTx6/3twyWmLw2brrzzuoDXgLNaHC+2Tx4v5HapXi
rp2jhcvbs+w5hmHtgS1o8weIpZOIPglBlc9Mc2X3T8uNSaz1lNhS5VjOzvxJXnryFJ+paZoX1TLv
zfmC9KCz8Pwwm6wLztq7c0j5DcwmC7I+4qfOSIjeo2u5rq63rrW52M0E3nGKMFrcCYfMFtVQxWX+
SXT/4JXBTeW4jrLR0Yu61IcVsJk6uc4WMmKl1/SpEY+JBi2cBYPlHkb8JQb5+O2JBvTMsE2SbtDb
fBfXvbXNNYoXe1wCFHrSpYXNGpc5jimR0uGh2wEq8TRanGCUEV1gZXbg7/prRFnBuXU4PG7E6R+m
Zc5WNU6NGQeekMvtMlmOYI+PQZ+yx/GYGpa+0rvTKx2tOTxSvgRP3qxNWyDjtKyAAkpSWK8vWl+J
FC0n/cygAiDmtmXiGzYO1CIINgYj7nMem+bB+RvLZw/9OrOHuyqUl5d4owY8nOiveErkov+i2fG1
yoICVZifVe/0hesDtT5D5KLGp4dA0WUHtHFEnAUZ7wlhgMoRbCANO+xTUp1oNS1xEQPM/J8LXXEc
Y9yJc53YIVA1jLqJSGErS2OuHvjSvrNF0sTPQeiwSFvsr8xX7n/lkAUveUJRrzvUFajKP80QbQtZ
MWlb3L4j3T/ck613Wk5AcvX7wyhCCkOEn173wRL67uI98i5auVLRiTguuALpiomJheAHAmuojmm2
+jxjnvQZa7WRCVHrNat/wssuqnwvuY4kr3pL/VUQX/lQPO9sfr9To2eSyDfTN5FeAEqY7CZQdRgP
WUUz7v91GeeHq+nAt2/ypE4xsjPo/mhOKKkFqNFCa8NuvCVJN6vaHN4K/WULGdbakDHaNY369SyS
eO+2xz6GXEr6m9FoxI7/VNqEvJAv3a6TTTsZBEjNw3oeIrkKZ5jRQpvLu0t9xgo1SKKPuFegQ4lM
MhgkLMs4TL/WoKvXdN4TC1OBeZZYoK+5dmw9maHnDTDqN89xIiBP9mCPLdawNq1nAfuJq/cM9bHq
FCaOfhhZG/SiuL73afiy5PUUyEU0BGRxNJpaFuk3aNElquQU4v+tZMnFsGy571bde053OhFF6w5T
w+kOLMr+4JP9iXK7HS0Vg9A+FXwuNog+xTDTyy+0nhT3AUOXA9lm3MwZILNl4T9W6iOWlXMUOeN+
I2tW9YrNlo/OEGgGzY58Im6YSu16zP/Rz8HZQQfvBUgG9gZkMLrBxPpaibtBduZH4dkyJSy44QGE
rA6JazwMYtd6FPaQOHKQEh9CpmmG90JsrCfxTzNA3kQmFZyXpTCcSHxrrKhOomERTqlCvIkkn6HG
xzQDOl7NPoGQGvRznAHz7sPZowyqXk+l4CYJ2Nz1m+0QVtB9vQ5RGFZO87451KcxjSbDNJzw0zA8
ip+pb2reWUGH9lpSu638+bcAk1ofUy3XiG81DSAU1qVSkt23CmfohxzvmqZTE6w3vh6hujDKKJh2
GyDYY+/8in6XCOe9WUxlPw19D4rnBViPg90if0ktKsD9qGUHYJFjVd5/oBKdopiKjqylOKGkstGl
BsgJFsreg5lhMtT2yxXCAPa5XXvQ875F+sXkdZGLzPYm61VAoHCtmXKH2WJ3MBZ7hEIcU+I2kzLQ
byyRo4+g8THY/RWMni98wc7MLvy3Q60tLXoL5jSyseFhKnuTPju/eHQJS+3tMgHAsaAJtYroH37F
ZVJQIgPThUA89orp4u3ms+iwrkeeVr6RTKE5tlJMtDaR2/AHMsENdA8Hy1HvJiX5HyEtdDgahMUU
AqxIpEsChUyx6Z7f1P4YxIGDD5OBy1TbiKwsHBQBTuIfEj4XEc4kCnI346oDd6X5UWgP6ypDCECT
4cSuI+iVD1qz+akTJf4QkjNW7EG2Outc+ti1Iu4RIcUMB4yre3Ch3AsFBBOV9G1ClJ5Zyn2EPm/6
seo15iIMxBPnSQZG7fCP9eMp0l0jFNd6fzHKl6NxTXo4rSazOCHpIapgE3C9+ZVp75bbIorss7Zs
u1CiTZ6Hw0kLl0xKWFcVNmY4JTxSubJJmxwTRvgxL4mOQg+3pohI0Qo5rTSmFocgpOudiqE53Q5t
BfABDsdQOqL2VsfNDD5pg0fv1qwCQEAaiJk2eB2WgCDP2FnbRbmZ/xJ8txt61n+hmzT6nZNlm1oU
4hqIBakloi8U8wWQFsA1RIdUES5sQ/vffoquBEJeMaHTpxq7kgNqeZ2tBziMzHD8jQOvW9Ej+XUq
CqdwVVPlcKvHUpdj+/bNyPnbZjqqaaB8ZPj6L+qzkYF0cbzdXhNmKEAMMRqWgyC5581OPZ9yauEE
+vmqWTDpjSKVGmrER2ykdK73iVp5q80R7MtdV5Kl6jnHfCu5OU3WTG3732mQJs/T4dQqZH0tiz5t
SlR/YKCltO7JbZSgO2U7d6g5gn9NPlg5Jx4Bk94Ao9LOexR1bTX6ePnTm3iuokbOW6cxFTw24JOs
xrrfcfve+GSOpKZaD2yirz77+ES4uiQ70pEHnQu7eEN5/7hPBdvZhM9+k1Dmmbq3yfJRnBKN9AK5
8QoF/wsRM9xt5RFwE9Moeq02TWROcNFu98zMM9zAcXaAf+gOjUpHroq96FAB4joTEUr5Svua0hHI
UFgXv+p8JIN70ergtAV16Orskg0Ug5hp1CAk6a3hfNmiwS6Cjwe6SEnLbZ+mz7u3lMJ9uTKsVscc
gNuEkWK7pub1XTGMDb/0RaSg6pHCdUVITbaU0fcXci8meAUEu8cBnIMrTJGvBkNsGie/j34sax4f
4994wkCplHG1QbFg+uPzXfR52QgjKKaFY5zxbVUe9xHcInTa5acURAYfxX0XVHCRfHqPjSnY/ifG
LPz/j75mwlEK0xqxFJH2W8UEu93vpvZDQBEVm6h2z67v+Q8GQoI939tnHO4Z8X3r9VIhHQdLmByb
4XRTyszh/+7Mhvflj1cZ1zFpLCymdW/s1SCvIUHZmI541U46EQQyGN05CsN7gmRWEbQ2V/03C9rz
KfShHVqaSefRqQlJTZmgmeBCH90LhrpeChciVR93zI6qEnM7jd37wTA7lyuxSrSnYyuRgug/+lLR
oOU1dxx5VwO2buTQkWery7U/+6MLc9Qfj+/HAr+VI94Kv+m2v1cqrLk8w8fL58QYGuKKfOuYIr3t
h2NZJhZ1u6gtT0FVVHxucIMHDRsVs7PHYVGakpJ6GoV1QVvOk4G8osH9MNgMqUFTN08u6jH3tT/J
hsRlvh+0InNR0fkvvXZhreQCjswuRIuHdZIUZyU2AoGYIIbCF72K0caT8GuGxm3YFAePQErU2zRY
EqMg3c/3K2Ykfky+YsUktBPmvuxWf6lrcSvuk+Rg6J4xg1VpW6Asytkk8icfmqAHjc8uNt7c2X1u
lLP1YGeSLUHS9iTP7VEhUBzebXMT4q1twcMSeDsQcNchcJbl0Lk+aLvOjjEbMN1lEV82JXvqf+H/
l3EArWdQzW9Q4bpYUV2OxL5V0AG442nOAHccUyeMwPPfYbWI9MJxI9uc2O2/nnr/7SC2cjnMSQ7r
EagJdJ9MnMLQrgTl4LNt+VFQSXOGDNuKSdCvZsQo+BetlRm2zKs8QiN2tJKEYWugnZy94ent63aM
TXIRqKQQ3NB+4s32qCRhsgDiA42YJHffjxBeu2Mo5ydiBBZ9fJGOfwzHDlkE170ltpXbMGXrvUdp
IeAbsJNEI3dQfa4x3K8AK7XuywLJVTze8Hd7G7jibMyyd6sEHeoMjgSb7StlTsnVLfbdKJTcDnN5
Bu7p1MSiVZ4nVLDpo4bQ75fdIhTFuOv9dW73qRSIL6BbCmtgA9KZOh92XGnjB2fqIIEdD7ageOiv
vdehR4bCfTOPo/Qp1FABbTl2M7Q6vvUYtU2Ro6nTcrcLXOuDxLVVahl6MVtoKK0a+XVyBug0XqiP
9cZ79TqlLVgtyjZt3tTczaAlenPfaA+2pobFccmd/gtpU4533Z9QnK9d7aI79yVXR1yUo+ZRvFfG
/sT1pOg+2QshAN95v3UedTmK3+jsYgbGOI7M61Z7qk6Y3DhwnEXvciU9J4LZh9peZ/FvkyCaI+52
wqhfTbI0501KgIJZ1wSzW5QjpqQ8yF9NPq5GTAIPg7vUFp/6dZgh5JgczhTn50rtIaucWraAoqS/
3VGHI1IDUn1uoGyvwa839u+YcSd1EdLfe9jrzDDzY5qS8phIyd0+euQlHmIDrAnxYWedU5KoehO6
d8CKcWyxhN9O4RFaQFhrjwhN+WqyIQeP7v+uGm4u8YWHrcevUKFhpfkd3VqVsqAXoOWlBSmn68gG
l39CKh2JCpiI0cTXB+AfsXQHeJdRtnLmwbXfSrqnhfyFfmp9T0D9q/2dXFalkMPJGaL1i+t3FkT3
XN0CpuTLmlqUWWwiwOkOozIXKPDioerEx3XtqQHHQTTSodkat1/OlubHVbdiu/2gnKB6S/oW1dKR
a940iwbh8e9Ccj6xl/uP9Oktg0ydPYWH3ZfGHwLGKS7vZMyOc/vxVbyozsw9hqBn8xgdzzBa4hKp
HNaIy3t9K7gBmBBVIbHSsWlMWDTGNJxqga1HZyRguZULcheq1nZpA4FHwECpviW1smYlQirQyFNj
f3eIv5CFlABgBglfpMCoda/pg76hvYiO/R7yvrNkK8Cy5rOyfxCVwt/tqcO/hGUjHXKjOh8B4fX9
+X8A+8MnFzJPQ16spywGIRk6f2CCH/68gGh8tqmEivoGJyK7OBfwhqXSd5oDCvHpAC5k0l/ej/zy
P+ApienGpbVXuhOVhbVGf8/bQFmli/WHvmWvQgk0DwhZ0GROf4JMALlp/XSPT7dQ0BLrJi5o+AJE
Ed7fvNr0WXptg1seYjmhG4SM5ONK9Zk9VhKuSQcDSRDNHyTLS4j9RzQzzLLjQD9Db9nlZiKxprLI
NH1WFEd0r0lAyBxutvce8yvnjylD+6tQt7WpIHwYb2EpHo3xHNngP3iT6aOz05iXAb5Vm0wF66Wh
30csTBBgUogHXxh/bz40u+9GTP6WKDSu7o+38h/KiArRoxjEDXxbsPTDeuBqYwcQ36k908A/n5+h
ynaR4E0ncGJ9FEGct9j64fynbjXhpJhxaO8dU5x662wBUqKDYjqFLe4VHk0sbQBcabVNbZIqDqPA
HBYhpVJMiEXjgmBiDLVEcuJ03Ok16YiPWkyCFoPAH3+s/HW7dIpyJ5BPNE1+eY4QJyRe/AfE90oX
+R2AOX3yPGieTdlolYQzGIldav9+Eso7ocSTIuT2LfKjveH7eW6f+RHRRcFt/INxu0HXMO/DxAG/
IYXTW73YEWS+1DvcIJRCCXQdPH62YrDPOZVHwpN9mxQdTpDOTj65PuhCEXcDE9fWM+DUbJHjKs85
HLYGxz5NRYAol1ST3PvDNfgPtSIvi3lqZlteqPpmeeMG0zwoO7/LGuoSLD90yCh81tLrxNOZ25kl
91lJ1t2z7eVoDpnkLTqWx0roFJcvcogTXud5lBwxT7+/jfFt/iLIDW35f7zyMEzOasxjqTsf0PZt
kQO3zmriy0vI6Rm7mqfA1LK+78UoB61D0vNRxIGh5YO8LHZGQUXYQ7c8QXwUrL21Jj/rCrv3bJhU
xHPqdQvC+zfMLgJ+SnPz/wUi2/TjJWMmibdr2537PJdopGajG36wXajsP4ZE56pkG48WmBKWUrha
CdxUcA/zSUqpFmhw0PgwIaP4I6lQ6rX/nlvzPuDVCOl5NHg5I+Q3b7gUPgeLY2DHEwVAsYaiC4Pt
5t9FS1o8mDiKBERdKhay0Bi/jJCkIvjfbzftCSJu/JwTPOxziyywcL3luOw3bMEkwwS9X+6iiKQ+
3Zus1FDHF44J+pD7hX3kAQ5KpfaE+moLj37Bw0QmW7z4TJ8UjaZ5z2ZoyK5e2WML4OlgN52Nam+s
BgnpR3nK8WR7EV8nRn0WO/3GUuEioEt6LCCkzcOrbmLYySs3JrfDtX9WVg1mJGj5OTkV+TWnKGhQ
YHiiKpCOwLrMriF6XbbhV74kNCJEcGTAe7xoC1kBNUtaaezaEifTml4/3EDcrp/JiMPzelr1ge9g
eiS963uI4kNDfH6/51mzJDYOORfnXChnEVV6QmyXIBlgshpQBFfXXTumOajn1LQG5GC5ZvZ7uqNg
LyfZ9e1DCovlXa+z0stp9Dv4FuUqWgmxSRSztltcihQKvBj58CtXBiTJhMxG3WgQD1jedmvMSUPt
dA+LjoduYt2928WAUEb0Wx465O37HxMuY10i823+ppPBYP97Sc0E0YmFNicFQ5frt1ufB4MJImfm
J34fnWgB+6nQNYYfbrcHXCnEb8CjrKkFZpYGLLMxf2ku+AQ4auLacVkowzAVStAu/JvFJekq69yy
3oOEFPbR8ct34Pgm49KZpM684hGl+kKUyO+AYgcHuugSkS7EhbywxnBvGn9O60/s6sIgl/TJk34D
4dpA7m3kWuulU5LlVbb5q7scRV+UW4qU9tm73H1FwRWgW92Ou/LWezQTeJ0XhVBgRZBph9Bc30xT
KbPgfZlTH4kno54P3Sd9tgiJ9DajpiUMQwiwRp5R+mXHhqek13dld7yLG2yfTyvxx4UmcZabg+bM
3g6/ef/c/Nw+BphsIoP72tt0iYHITVPNNhK1929G/eGfNsdb0L1HTDZQ333HLSv2CoVelwJKynF6
N1gy/YwgIAJloNfqTu88BDBdtXFWb5SgtCDrTyFOzw8X3IvBHKJlQD59DDJsrdqx429QvpySbRcI
iXK2jyvoHnRNPgvQ92dvXEBm1R1vS3iwcfZqPBjRNDbjn0agD13RJVrkhzNR9jtROuYGDUU4y9L8
h6NnbxHZlWH/L4RpdnEwowOHzJjXttjOT6cb+wQEOclekxZN5m4QE2vHagmjINWnbpiQhBctrPxG
EfshiH7hF/t8OqyvUBGX1MURbj+klRGrwtJOpOBU7ktVBVwWPtIx9ID5w1UbMkevV+tLGDciUaRg
qP/ZHixsvs6NTT4cYI0VW6zxNBMthEYCOjaXfwhcm0MrLv8CSFaldI3FbTRmWhfJqW3Qs+DVKfol
tSuAsjoJ2wbJs5SwbelKYRU+HR2CBHz6wjll8IeyDwjz3bLVNE/cv++MX0Nzrj6JMgkWQGyc80dh
4sf28JmBqlnEalMyIqWnEtqoFOuCnu7oRWlHpr8IOWJSywxIqDxYoY8U1lqSzO9Zi9hEdGy6y7u5
PY2+rB5hCFdoKKSxmlzGSBU9xqpcUgyb+FFliFjprf3oFF+3dcs81EtkYmG01cnD+ne1G9/yoyNk
XULVd5R04CmsAKXOdA9TEw47EoCGtGXFwvsCgm8sT20mS8TXJs/Igce18wgbzUREcpjr8FnyhF/u
FR6lbVp9Yqps/2vMdmD6TE47ff6MeUYWGsA1haV5DNkhs8jdMwUpLdGSm5AyTFteMbFcZyFp4WR0
PUzpn2kX8GV5g8m86GvtuBz2145ueoUH6jO99/cvjvqmvokIuC9A1Bn6pT3u3dSG2bz8oC/vH7r6
pkkYaHOEoHXi4m+63+g1o0Oq7BBnuuft2fhF8Qv1m3OruFTfaWiTg4Z5Wx0h33At1N76nCTuLKOZ
rBz5Wn4JnCo4uxZNpF5auNfUvN81FIPkVe61E5u3PPFvBAy8T9M3i6jtuaqlXG/SZMtAe/I8aRLJ
Swh3i9eBL/W7JXNdndafHxin6ZS4hO0SwyRkmUVcQfYtSEz8VNsYZqfww5ybN5Yr1CeqCDAqAM1L
drdVGkqL75zk6Lb7QcAyf98Eg7Wj24Sr7UGLQEO5u0fR9zrKrRHE02f1I1FFZcnDq63Y68YlzgSp
KrIBcEfBaU9KjNWofk23X8VLcc7L52jdLRF21a0C1sFFBZY6MQwSVR7HXnmugW99AA7SjqVRqltz
y2R4k4UcreaDiRMziw9AJN92qefYW3t8pISyZs58BQNMs3ZRWPkHCeMvzWIaBCc0W3HUMWLUN+qD
KV58Ur2uyffqzjj+SFQ68P/BUBlEiFOWArZkKOdUtzXqypJPj3JgzcT+BTZ36TPAIAESinsUfJN5
R5guMsSpd4w54Ql0r0Rapxw1l2SR8ah2bmNE0B4bzxlo6/WsJCTT1yUpdO2aMXNzca8vUJ3x3EPO
p0kutKFw8I4bYJL4IAFy8sJOqgwQ2djcZM6YjyH200V7DUdwRUl9JBUcakHhX4LxkDIrdbLz98PB
xseP9PJGrFN7aDQixKO1JLgl7EJEN66R5JgySf4mSdboNrTjQx8nNykoE6s+BtxVRDQ5B347ZTq0
yGDRwiaUhBHjXE+44P1G0yCR3rkxi33DoesISLuwKHB7i2s65aBKkFYt9bxpzkDcdCqpkovCyCOe
Ymfe2SHZUcx4+e6oyloQSNS5qJbnNKrTVaYXP1dLOZoQYvv4Oy1AZzli2Fey6Q6Yclh2LUp2zYTU
spMbZjjfTYMqPh2fvGZfBamVr+OAEjVkX+WxX3Qs3DNBzbBwhMAELtzRvXI2C28TQvJM2mqzxNdr
tSePWl7pD0UuF7b0jxHl+bNv/+pFmpJRMqfK99rjkudciGwDxFvH9OSvUchs9KZbSX98H5aJn5gU
043FBxFK8me1V0LsvN87hLSQhdaURDrgwCDr0nHPHZlJOq6l32KEdw+JD5GO6TpkuCWeWOCAPirI
/6grp2WFpvCAWB4M11KiRDZt2xbL+U4YrJr+amLlKSSXwqE9lFxs4icA+c2TfD4AiVKuEJlyW+kT
xu2UwNHxGlGReX2HjQMjvxZk6THN5l5tZJv6KSngPcnk4lD9sm7ZCyVzBhexK9aOfMNNksa3tsru
FDbEQhM4H2lsJlVx3fat9IeUZuzQwhzOr7tYV7MAu/QVz3lQVNklmorIiXOCx06AYCWzQfdjhRCy
AIwSFxsqtT4crv8Vf++twj3G0hyyG/y02mh+Z4HOmCV21NxLybyH64D6o2zk5ExbMBH2YY0Rn+ij
YPicfVsydUTiGr7LxcvnhMQAvrxU6fNlNk5qdbZXjlSMO8Qomm7fhTcq63ZTPWDvkIoDrAfa3mao
W0ncDfij5FvuxBYUpzzL2twg/D+h0HHV8yA52wEVc3n02DIDWYPHhPdF+f4FWgRhoGAuopzV4kKI
UFoxdGBxOcEU4NCsFpJHqj3nphkS5lM7q9c/u0AFar89yEWG41QrtVT6Dl005fibRRwbi6tspjfx
yFeY2SB4Q0XbDfKk1ZZOv5xbbIEUXZLnJzX28Kw7nKf41VSr+dIlOuEvFr9drwZDdNAuQ0hjTAzo
NxupERHnZv2RBrdVUlROpPAjANDUs6524KWDcaj56M18Tfay7x0fJh83ubYBEsvm5kMr3TQYco3k
UKsHKePvtBoWoKpiN2J4ryrI6+uJmGwoGtKeRX2Y59iR9YfDgZ1wQiBC+jt5OGOhUmxQNjNo+Vb+
JwbT/+uBYRZs0r87YS6ClT39NutBt5nLuYpKmEKBf6nswTiMUzDCTU5dGVatvKUKDutcAIuhPUVI
BjUUr7ZM1a9RTVaoANDtYLfmiVUKajbXjKd54TARbQdcesjdcte5mBohINTYKS9nAAtvH0ZQnEVR
4YXN3H2qd8yPEutm3MViFzvDFVxJI+JgZihjEoFteX4fIhvSSw3MSZ9Qa8hRtWftgeTu2xO0gRNg
xZlMJaGtsAvUYHmVhd4wWWKlFF7gGTCR+M/2L9rS6w+x/VsPWtFwSmMiaYqJcu0eaQZoRUijM3jZ
VGSlnO7b3qZM3bTgG4We34NZe3d/JBN5GMUpvLh31gjdzzJyef18BNHerc+/d7R+iInmRkVuYVM1
oxWb9rn2t5Bmfx7EGiumUaqxyUw4hykHxW4bjY2VASj3mpgkNgkJ9ZVFzfT33NbHdFLRYxa3YJSS
STG94XHu09gV+eyBE90YjWp6v7xwozHX3pz6WEM/cPttNf6c5QfAuOgFQ98ziJsdyCFuVxOdpMDv
Id0R5rTWTjK6OV2dgA5o/MJGjNCASud5DTi4Nvrqu9FGU4s9zvU8YQFEjW30La+8YuYnXzR37Bp6
a+8LkfZfs8qR29li0sQ5RxLZW+2ovJHHXoRvdITzIjh8chgPA5qII8m9fj0SNgVdAR/czJNj+Dg5
YdSQDbh68M+F5181MzuqWmDtNbro9uW9G3LQcihIujTLvnF2uLdZar7qp0rZkgzEvaP5CP5Mw76L
8dgD2ZuyxVSC9M3FRyDtdHbSKB9fuYqN+OY1MMTLZthe4T1gOJjiQJs2dysRohv0v/JgnTFVWjU/
RpqzYATWL6JGmF1IINHOfdoeZj8Afnb+UPtBcs5b4deEzhtCbJxEQmDR7yDUdH8Syw6hcAnftXYg
EA46Hy1Pxmpb3PFTBUlVZ1cxv3im43GBjuy5ZX0+92Hq/3NtjxLYfsJJvQGbnslhx6cdY2HEKdJR
O1VjQWHE4At1Uw9fjukAth9Nccsl+5M/6Mg1xCVcgigVuxwNxJEB592lMes/Z9SByWz04MGbvJkx
62vbUDKt15nxc9qJBYIDoRxT44RKk2bpL1wlLCuGnJLHgaS+4Un5Oy/uEH7QBVcoaxoujHMHkCzB
yXwJ6paHY1gnVlQCwlMR4Mtz8righPw3L1bfnoWbej5y2nDRJIfDoPxh2hYnBCh9DIxqUAt1zBV8
r+mZ3XC6xgo86+YuMWrvSK0l1jb5qwP0Yan76dcb8vTOcp3zgVrjTd7eJvsI50/oGxa75kv8Ed+F
HVFXixVIyR22Y3vQWHz56GP7trk9IXNTm3Jq6P1hu0AWvQjctxlz7MBuY8iFmJKx9u5mTRfcVsry
9GGJPiISt+SgMwFY13fDgu904VN2EK2Zx9by89V31l3W+T6GJssrW7QALfz452DQcao/ffmVFOBX
AkK9M91oEj2TecsVdDM6rsc2FdmNmwGqcW9D5K76Lf9kwKYN+b2SC+/sA2S+SaOty79wi82eanxn
iuWpuQX4XiXlxNG543HBrCMxnezg38DEn4Rud5bE6E9Y/tQOkeQa9GZ2XAvfBbsk+R1HB/4QKZQN
TFqnMFWpqgZITbtkkPy/TvRCvDZ1qoIykUO8b5jjCM1ftJZJW2AoD4dW8I0HPi2yL7L7jyVKhXrg
JVl9LuhJmTp8rv/Nu6bEk2+ULF9ArXhENy+3A78UjgB5tLQQmMkvZK6zjnhr52ggoSBsqCVaAmyF
MHGcB4XOGsQLijsSVqYVzrqO/OqdRGi3FvDqAlozUjeQXNHt5Yw3jrU8AYP6jhWypuZcOOPqHw/6
aTUmhmjHZ7RzKZt0AJCieISwZ6LeWY4NtGh2HUHQDoU3f+DKl2WitzCWN2b5rY2+BsOEwI+yqXoe
EIg+QWVi4EA86aZgjswRqMC/ZG++veMgYY4x4cCjOzYkmVDDa1b2jyD/BPmaHDA+A6f0Sju8t/Pd
UwZSJFl7omBBiwGlyneAOb4jLJKetlYNAwIkgRplso1eVteDQtCskYl86V28yu28ti140fLz0YU1
c6nR+EaX/iih/aQTVFa3cLOeYeavFRZInJ1kgepk/rBVodo8xEWBQvPS+vHYK4+6LC2sPT53ZLt+
CsXkUnCfkKQTfqvJBrW7Ct9Pr3LFBYO2OS9EGXxE0U/HqapbjC5FdXhZQDdrhk5heJ4ct2dkk+JD
EwLjz6exJIa2jFRT5mveCMS7aMmFgMKXfhRvpwPsgVaZMzR5nUIzGdYzrMh8OZPN2LCLk0Luwlfm
1NiXCtYajrgHptqC2kcf8Mhb0yroVDXRzLhZ732mGI3B3ImqJ/eWTYydvOfDzDJGkq0nheHEqgzV
qmOjiMSWxdQnSEBVn7QgoHcbdyRy+JnSys+vEHdKtkWRQ8tqwX3z3FkVo+MMrVk84JvJLi5t60Pt
soeQcKlddYy8CAO+1oppBsBmlbgQAePtXPpVGf7n4K3rgRMnykvnLk+hF1lTeEaLYz0E9TqmMT5S
pdBBwoo8EvDYNMHSDfa32lalgdJZt1pkToWUEuF3THHmgupAI/CHR8yvCTA0jIVs3GBRqqXFAlq5
kt/fwFkcbb0EzuXF8CBAen0fZW8amP/A+cGN2DU4P5Tppc+ZzzUD4uLEjqeLWGfBy2V+4v25I8CS
uouEH3dE8gGZQm0BIQ7IeDbdkbban24HIVE24NQRvSc3Z6j6gG6FBVyqa5qaztppuym1j4R3edl5
vjs2YbdjavA5zBWm2zbfivpmcDXAhWbODzbqpIerpk344iukhuZ/trW3uZ1RsF4rWKA3Ba5MhAD4
oMhmPc5MlD2oh/iQzDcTlkVYAFufc/Z1KsWpSogeoBLdCbzuyNFwe48Yrvhkv23dwPRzpJxoVe1+
90HKUzAZjS/MoLI7D0fJcOGZyyKBDeugRbfjpbvhetKfgaPNKanXXhex//sM4/LNyBBFeq3McpAZ
UQnSN4qL92/6rF1EQn9i4xbPrvXrnMU3+W6/7J9VQ2umXDRXaHLZBIb/Uu7zZAEUEGvdNa6XErBd
ZJ/VzNKUV0aM7E2jhd9LimHXBi2hY/TSbF8DMtL9GPC69wID/MHG+uWKzrqAGsv4yV0GnEN1tatC
uDYG2OBSyKQkDnB+lPmOgitdFfSsyJJl2ebXt2RTZKRflhv3rc/0aCpgsjUAgMGjGqVU1naBj5KF
dXgA3ht2/uMpIdoW/vygu0EGapFnYtv1MKqOYrbJq/oZXHSzZEoymWj/DT+JNyXQa1ZuhJor1GYP
5J9GfqgZ14B5V0YIDcbK+CRT4cMraXcT9rQsXAB66eL0D5cdTku7xzJT1JT/5o4vGwEICsCfJr1I
Fr2kRRGTWIWjTlZyytS+c5dVerpWT2uWcdZoaXtsB6PqNSGpc8AgE5S3xRqeUph4hxzi01obF2kg
T8Xe/1bwphPQZqkbsXylqf6bnF/lv+PVkmWqgO5HeSIn6GgIgi34OHfS1ll3xkuEIurbYL5+9GfP
v0JtvM3qQtyHkGrhPZBz5OJf/oo6JsE1dUf0WYWig3dS3ZeEqCE8WfyLdaJbUDVs4WBFEHrZalQL
SZ9oeh0VJKnhw3O90FVLLqckyVHZeAK/rey4/iuPptzg3hrnfpNxIpXwsaGicdntLdD4oLKfdDu1
rwO6GvWvwD8Nr3DUu5sea+DSGSf9WeA4jnYbIcUl+R4VUA8WEtDR+NtNDQXXvbBgaXeHv5WCJNDl
VXKvMv1tqXhkhncasnLCDdAuhhk0CHJBRRFn3hb9kf60bg0l2fwJKQtbWXGb1BH1cuwHMAXNJALY
dojH4YRIQNYMkpMhNpkMEs1oLPa0BT/0RTbPozWxPGgMThMnTSypQLh0hXZniIOGyGIDJMKM1BKd
d1MBMTwR3EYTQP081pVMrFXAUNA9yacOQi2Y/q1xm7ESEoJqnBLHthWAvfwwIBAYSdm6MtupKgpY
3UWJFvJF6/LMm9o6n6tntVibgtd5m6YdVz4L/LmojheygOV9MhV116qpVf3CgRzQK5QvYm3UmmQq
coZq4fndlhWDl4MX3P9JdJK8+Vx2M+Xinl5PYeA4Ku6deaZsvGgZVsARX8PCuaZYukV45Wf8pb83
RRAyzGtI8MU+c59cPcYSJp7pgL7AN/g7vq2J4hAadUfqfZxeBKloVMlTQop2E9nELW53F96EBfVi
yO+7xoOl7dYo7u73bp/rQw4YxZJSni9ueptFUXkSHq4nqd9miyyATJ5FMwLClf0wH5N7mWaYJIRW
KpvTUtQT4ZUkyyf/3rr1eVr7OLIwsP4g995HGlCqwqMfbXXplWYrVGdwnDRU8gO7Mam7Rf5dcHkb
cET9QwQe4Dg+S2jDS5dhiGuz+pc1naSQIFFRwCvUE5Rx/eZ5F2jDfocWpWbMIDL9hED3H4jXlUha
BuYA3c6VAEISt3UNX/GLITuLFkllqqwSl7Qlsay3EUMZLxwf3YR0JBDDxTM1ZoZ4j+s0UhMHzsF7
4a2URQL3YFdmwp376hYwhb7hWWuCyFFV6QgEeDF292dPtKiqNYmUT1i9yxvozrWhrZs//4TxAMAg
fyrDYQz2aCd1LEHocpnXXGwbgNoU8RalPPPw9vEMUc35ugD8G7bvidZrKnPCxPgRi26ZQPkNgIod
AhTaCqlQyvsE8xNMu8t5F3Gdx/lBf4EEJUC5nwoBq+tC+2SvNvQV6T9vLnAeoqZPXBQ8rdaaSK7U
ir6np1AlzxXlTBHIokMAl3sKpushGCslYaZ/fH6RP7lWxdykr45q1upfoG+ktRT+W3JbI/6efMpp
p2WvMD5NQlQ9S5LOfFYyD2tJ5OQNRppipVXrYbheXuZHGZBSc3hWkKqBOSkVi1WhOENL3RGH5zrB
FJNPvZcIAHJ5VybXt/tJN3Y1RmTqxN8BELeMcuVt0K6PDDhdA7Aqk41FWVereCpVx1vVZf1sOdgy
br5LeGdxqZnRG6pM+YnQRhC5cahQwybgjE2hBCbjKPCPJA2tURZ8TnB7M4ODza69hDSsPSugpsMy
Sau0n94kWlk4/EebiuvttiwQUB7P1yGrSgMRizV9f07o7pYRGukCHI6htx+ZG7y0El/gwaN8sqa9
linzGrMuLjna7hjlzMoWChR3+v8lj3Zt2K3quc8/xantpaD4WDhztj+ZYtBG+8dRiGXsyKrG/ugc
Pgtsyw1UIG/G7YK0RuZYTb3n2AJmKwQlkjHFfDBlr81rMmylN9kRd5snRBlA5gyBs5AzZ1ajOxXm
bWGWaZSdhoZp6/ESAol5nFSsrxXXlka3csz1sdmMj1W1BtW6y7ikBpakZhLZt8TYJkTxcwVbXFTT
LU5cBDtJUxOp8Hk1cewlty2CyR2cgxZl4z7V9gb+osEKPIM69nzTQBWzvWuE5hvVE6ZTXugN5S+7
wia46x1IIFDqrp0gR8ywc+ygIJ1ygfSmqQOGMPShnl9lWlFBIlAIWfnz8ZAQnspsY+dJC4JP9S/w
OCt5+LwcMYjkhX7Qz3jEk/dTpIZaowFgxNcRnfa7p5h4YMTg6bpiT0sxeMigYmOnSNkfbYCipxRC
39PP8Iho330VO4KhZL8QHd8gwD+JWa+IrJ7wZwQAh7HEqmV/QW63ZmSdeUhyz1GP7fdTcM6eE3LI
pYMGzLQ75gBWjwrRKGiDZYJ3u9DhOlXIRFarm2OZU1mXC/Gzvjcg4JOSGBfuAnN/MYc9c7ufvBir
O8KgnF4rKf+srHeyxNMgU9UeZ5DOUYwwFCVQEVBEj3IXFsq1AVx0pkNO0clxKlfUV93T+lVDl9/P
BLkRUdTuqWxplGgHVigwx7Xsa4MhaMSVBr8/IZI6U6tj9SSmAC4MRRrW4qzcDtFnx6WcOU7CG99/
i+dnw5jk0rRy7vazIk00vIZ+4BEG01PTf3sUZm4zeoBdhqUr7I+pEdyLDCAwo60ldyv5DmdDiAjc
fzzDKJBjfQzoN4gGRdbRJhhaCWW2NJ6eGi4Q0FAejVZGIyBTfL5JW+nSyHwY0XgdoDLqzkfiooMz
S/Ol4+zT05gCeL9S6AFsVVRz0FDs97ay5m1rkuUy7ibxeZX02TUt2iw19MbICAdGiwV4dfzMXLi7
AOXLEuk56UFLpppLBu8RDEZoRxURtWVhVprne96yV1ndVlHxtAT7pYhx+IS8xBFV3ci4F51cv8Tt
B0qJATPZ2ZWEDF2JDjXB8XTTvlSJ/7ow2TTPF2uw4qH4B1pr5nbxIh+aHFM9Mxj5KH1i3FUmIKYm
3mk5xZlQSlvaPKYMEQu6JxIDE9ouxzDcynfEPOAk7F10HNOsnKYArV+ESExJQ4UMPStn/f2UDioG
7l/BNu/0VjJOVdmhv2Dwv66iP23wfWPETNcQg9g7HmBbvoIlo9aLa5u7Zam/QMzlF+LnTtfuvV2y
CsfUqWjHB1Jg+ghBZiyBpyzYaYv3RYh3411fjFg1G9QBRhwGUlRQrBE9XVQOsvv1y785VmW+oLyI
ReoS9NtG+H73HNI+zaVRYzq7mUnfLaOCADSJs/fgAOXppvtn1eDtvjUIErlYT3aGAM6L/RPLlIlv
h/eZi5Qndt4w6wTCpvmf/BwkoyIelr9IMsM46RIwaIWqRNVp/k6SdiYbbczPTHEvwj3HlBHasHaD
8VLnVpWYqZ+0odg4JTDIz4O8YOUuLQ54WkdNdGDGOPbnoSWVQAQncwSxVrGovKJVce0UZGnV94ws
qyePFiCJba33uzPgNC38QL+YLWuDHBdh+GFoBqEUaeTftx74H04AxMrR1DWLUlPt72Pp3IrRj1DO
aDNRjfNopBsQfrpbHjOxegKn6fVNcvqagEJ8Pw5cmIF+GQZaNuDQSpaylr3QDOcXpnIgBDxPNxnN
eKodTaQgbkQDLpO68h5wjoTklJjv5Bv1uVei/kddQXSLjLIUCJRJWNEDdEMPKIKsjgH8ttJr3/gc
FkGSgkkZCwEHQomwjdqFWKs5qw/D9LYlqWdeNBuq9Uf9a4SGt71FAO/x/woKUZIUdJBA7IaVJ4Jk
iznrJCRVQaKPqHOudm5bagh7H2RLpmRIhsNi9oJLT/5TMwfmBASkePI13ji0fGtd9ov6uY/aMND2
SkcKbkTcOQkxD6MUIRa+HtUptuQpfhYOq+nZmqq3WpNQrkUIeP93djvMDZdOT+GRLk4bCPgh0Cga
McbNKzPjPpBsqeOzHsco63EJ2WzEipnZlDaBonzuUYH0gUNbTQD/Brxs7piL44xGl9XAMTU6ypCX
+dIs4Uz5Hw1w58kbhA0cu7yyIYPMb2TJTTojccG8Vih3zpwoz81ZR9FVxAf6DP3MBTFcV9IBxvfS
5TQh4RpafCDA87SjyO4RpF+cABqtk8eVJkdL36/jB0pRz3SYxjXbTjcd5WnRErEDAp8JOQKLfODB
TSHYVt/D8F78ft5AFHefCyh6rfwFC/oFuX9+dc9IYt+JrtJHdGudcPNywCLcltk5n0Au7kil7pFA
ExZCX8Gmia8MvmCm7Jor66nyJBhGJsHXOGeXTsiJNBPn+UAacRmHDwBwKViPT77Ch3apSR/IOCqY
TtwcLc+tM7NFpynXqVOIMBNxB6K8mWALedjHddr/SZcN6SgeMNl+T23Rw1eh/efsYMtb4GDBeyjg
z//y6eWOMqNEjb/y+mU01TqUju9fidWGMXozE/ofTQH9E/tUIVLuZyNC2JQXr0NA783QdsTF2VVn
owcMU31NwV7fH4lprErcjE1ypbHdDaN0OM3+MMbMgkVJCXPwRkRrPAuOEJxTi+/Op51I3waxnJg+
b6Bg8ls2F0JB1fsxlwDcOLaQjSTr0QfBVZrUAdWTGI1Nx9BkWQPgVb44B97mVJV0SotzICUGiMoZ
anln9jDxcX9oTWFQlACRvwWbDZfQXsisVrKWWFk4A1lYM74/irr9CupPxTj7bWN9W7EUejP9qzyH
QgwZR5PuJr6oYXv+TPG2FRLMm+tYQiHZnKn1UcsOnvHHQ9FDGt3L6F+YR5JKRO2Y9wsJq/njQark
gV4UQ1YAIcxE2KzSiypOix3bsgoq+r0otieDfUQ/WH73snEzlwCc5z3cfKckgpuAqfeFiJzB4l+3
ORXsegOCcUQea/di7WUaCYkYhDOi6r8UnSQ1sm6GonQSu1ARDb4dbxzYHFvPtn7Zf4U3/SrozGB5
kJxR0zZ3L/GXeqoPMW/dTHTSDwdpCSgCZWu3NfAepJMYgdlJO34CCOeImiioaLl6Imhub6PuUbSU
egXC7zdaLbAiA3c+qbIkMXRFQY2Xzbc8JJV8l25Cnfy7K3JNglQYxzwwYmxUkWG+w8vXWMJW+CyR
sDdCz7BNYU6sG1Y4zbE8V0FhSa09Plf6HU7xCON711g236QkRScRzfYqGT2riOmjU5Kt17YxqP7n
9G/i7ujQzvRvAAPMnRuwPIdJ8JYloSK16c5ToVib8GIczy/Yeeh77r+HFtThePu8Y17DozfD4E/+
jm+d0gJVh74mA4hut1U1ICmgsS6fwpHJGdKzxlBawBRoD9uNXu5f11hLbpS9nHpw+TyyJuAnn0pE
xygAfYHU5zNRYFlKCP4Af1fR6Oyz02CfNy/hSnyLuBif58rje7cuDjge2TzuWDZf1jKJw1cw9L7t
InxVcluUmiBRLqaZokiEwGRo2/vmIagjMKxaT1A7SlWUpDpECTd29u3Mm8jb61fw1GJmW1Dak5hg
EpJs8XbDeJUA1WLqsJ4TiGboigth13gRIJ1CgOfI63kwbjcmfwhwgXC39egFkPdxM2p/pq851V4I
003u31pm0pTnAGspSnlU8u3vpz3SYadZR+3Pu3LxGcervChTJHFPcdE1J8orViHOp9lsxkXbV8nQ
dekYXSZRagYQDcnDZf+yWwv6x7UDfPhSJnZx9sIey5dc8Jvh17U4998MEFtfSWTXSco8Lk8zAZNq
kHpXLy+WQ8aHAg5mu+QvM2uyg3wXt+/lzkQpZ7pz1VdBregtTdmYOC0sABvj6C3All6XddvvR7Hw
k29cu9iJAiIWPf4Bfv17QQEtO1Grd5B2q4OU964D9E4li2QA0vV7VyZgSRWpqXdEQ51V142CFbfr
jczQI2ppQPcbg812sumNmc7QbOaUTRo+Gs8FptEwCxCLnQfHEGuB6kKzHUafLh4Fn6oJg3sT7FIf
B+iSH20fqpujYqbgHJY05osMsGq5pxPxIn3wNifbvWC46PFqUQM3t7PLmlA+Y8HP614d8Bpn5OTA
if1FXXJ1V4K5d8blLBcVVu+8Hl+KZ6nZBiJz58aELXSiJqIFXD0SEwVHjMD81hRL8jU1REIXT48M
F+gmrEXIEjL5zvsYh2Qr4mUjtZfel5WVTP9pkn8bqck9PdRvGK41ayX8YLcldguWqOsrgW4ZRn2I
uE8y34SxZq7bjSEix5cljIG8jZJG5LrAJwYLIY630fYuvPkN8HekkvdF9evIgmYN/QEHZvo6+S4O
6ST5F8eBTJRk12JsFLMxcfPgjAhmUDlCp05kmGMrU+/sagCrudrsURWX0sYG5+wK8f6Vv8JEq5Gj
HpiS3kVPrOaGGL4HlktEoJMlAFeCYQpIgWGC+JwJghe6g67m0cihhFV1FtVPpOgdi98dKZEYZLnP
0igFgxSA5b8LrH6ppj4HQeDl2386gRlkc4oaaVw8X1dUp0RtW0uDvkpp8wHEc5wn4v5G0ei4Bohr
BYU7+bUjRK4rPqudC6v6e8XD42HY5jXsH0acjhx+JPP8i9dTR/VHwf7GMCJEcpqWphCb4qDGrK64
fmHGonfxcqwwjP68kvkIJV6y2Md5tRXSHjHAM/kxlS0tXbdfCe6O8p+yhHeImnvq/h61PS7yuIwB
6krso3u8gVwJzneSbcF8VR5D/OPbT4PwjXsgxX1SmncT77FCGgpjJtgx/P8AJUDqn9DFdrqub36B
Els05ugPJzjW99zD4YkV9ZIRZATbdbMpI9dN0X10MvSUVENgCWjn+GpEN1XvXXAP922P/4rZxAlk
xQLowtVIL3xMSkkLC9W/n1PXqu4EfbiUxAk5dur4LZWD/ZfJUBbhE0vU4kO10CKeZFyVaept9Mi+
Q7XHhNE5HRMfrzMmse0f8tTHUl/ggh76Wiw7oqadm7NR/rOy046NDyx2AeIyuxEavR5KIjfCFbC/
CpIavFHKiIp5SVLWrsyENfnQx8XeBRTvx1RYauHgeyuzetM4N1wE4l7VVYGlKy7D1ArGMZ+FyHc+
RJvCcGvyQs80RX7M6X++7GHroahGYqY+xMIxP0JRKzldLUx27GzLIWguX+igwpStU+Gn9AQ8Q/zq
TgFcsIpFRUnWBeO/8feqn5BaU42pcUfUs/T94sIRl5NkWfOx8gDFqw9UT61y1tGyDABoL0isHDhh
LcOOGUxkNRGzQECE8WF4suJpZrPt0gijrbMlPL9EXKkLTKL3+KdXv9igqgF0aAlT2bpBC0OCe78L
XIZHt0j/9e27pfK71UaLRJL7PfCEIVycUoXORyFTOdX0o3MgqL7khomKIEjmMXseNyrl4LvxsvPZ
OLln6WtE2v5ArwCmmHpaR24ePEnryTO+3Ci7mHHH/xHTMXT6GyJsyZDMPwjgyf3yWPSjF2/sDDG0
u3TDpcCJ5c5QK0oqvCwq8h4ajpe0brfq1UCH5dHoci2vv2ZAPH/G89Rs55R7L3fvwiGgDFHpDzOQ
vjItuPShVlPUigy61gXe37sWlHnpAFAYrmTRmMLGT309eIziiVN5FYnw+PFzyQny4vQ1DWHL1/YF
BCvyiXVO0lO54Dwr7f7hLcRVIHWUvyQyMElt5c5mwcuoeSu3bO64n+h06V9uYyPzoG5avjuwHDaC
+TbPIT4obuTJrYDzQ8qCHXb0rE9qiadcm6p+r/aisERQ379Z/QlhGzMmkujO0dT/RXAMwRJ3QuAq
s3mFz3sm8QNnDORa+r2ZSvK0Y9wjGUw/OAF2yIRuJmhioHa8mVGdFIhhH0kzn69KeuuQVQHTb5OK
o7tw8/O7GPDA10TDNVkuYQbtm0FIxkOx3CqjgF5r9x19oreXZ7O51BeHCr14ELZhrvFK8hu9MxOC
TGCtvLBhlWqNjM3k4WOx9UtNzV4xBxkwQmFQQs73jNrYYZmmyHKN5xgaUgoesE2SfOKuW160VdqL
ctu/BViU1TOEs09KN/ngL52Ejbj3HjJwDsgI3OQE9+hCUEKd/WqBEfQ26LIEePs/HdnsSZTPfOLa
5ijKWvgohAn1Ah8NYLNlzn7QBAGRL/ZdWUcJYDdht9Ka4kJwNdFTNzzHn6JC8PSPBCEhHIjDJ90N
OMp0AU0VwzotXf201oiwkufu4OPW1BNJ10oJqi+tEUQZAmxjhmqIpaoz0rXK0ipGOqWXfHre7F2/
QD3IuvZb5JGzVGSWpvVEmIjHFesJWjMmjxlPUwdEk7QENeByf3v5u/05h/ZvD3wr6vz5bsR/cb1y
UG1CRnYy4vHi2tBb+FCLkuLPgIYDFnsi7ssuTdAN3WOtb+o62SottrhggOcq6+pZtNZ7IxHI0F+R
tCmmmbvHVw6wOautrnW3/qgy3EGO/ka5+LxrRs9tfejiZZ/pB16ySbwET0cTZXAbwv1ywDyRrGsb
1MIN3N/u2E8k67WXoE+9oadifZRGA5r5zOTkLPfkQA10ZjgT53U/mJA74vnIUoTuWrLfjbuDOg4A
Dl0pkArvVGtM75HjPxGShrlKV5LDeLQ9nrcFIiEh0TPmY+xGRL4Gl2/TS02IDZPXvu/NlNwzi9x+
O/1WmNqGA9x9pNELB7ket4+cT1QsSYiSIlVSwK4JM5uoHQJ3P1NO5tfL/qCWTKwrpJD9IfaLhZ7Y
9yPEMu6CueBg3IYHHwf7EbRDkktmVJzUwo3uGpBlAPpGEcotN+Tz6jb79NwwC7AwlRwu0IwogXNu
UNADvX8IYywop/Csd3DKAgiHVORHLMj0F2LQICPRnli4fON6zDDRx2jFUeSY1QRliD93adQBYGrk
v/f9JPrejrw/iFQ+8MbAd593wdKwEOKWDeBJ6syceaXU2FeqSmTnJ2map7vvTW7Y2gxk5vGraDto
SIWLpx0nvyBfMl4xOF7Rn48Z35XtEUYR87Zr+7xLoHxbAJYgCH1q5XyY8sRQ28R4tlhL2fYudT1e
sTphSGeMaH2XDthiwWNjXODzrs9A2fZOUO8Yk9M2RJLMf+UtxFrGNV7ANcEO51P6PPSsNw9JaPo+
hzRyiUC+G6ycMaCg6yTK7w3ZUVLXWDbD+RvDz6tUTfx2MZO411sgL6MxCW2XfQ9769o+Fositktd
HXuYBN8WtVEfVVgjuHtRbx7DrYx90tbZZ1nDjoLXums+yq7B0A0do2xWWboHalXDmIERXhO4TEHJ
V5LzGhtOnpHhpsAzKd33NzS1KVSlM9pJhEE4DziAs9hFqZCX8JexABNBKd6XWIC5IjivRjz83yXw
xuVME4A6FvVRs87ePTHCX0kcXPi0jDrCc3Nt6CEekdW5SVubiDGhJRSSK4md9ADORRsB+gGPfFZT
aFx/BmDWWwSQTQs11C6UGDUQJkSFlwF7NokgUtdNT+C5j4w4hLG0ygsVVMZEreVdffzGfSUC8g4i
WOJRwbc+6GC50OvkvmQbK5WtdTAS7ge954LyZK1WPXhpTpJm/Juj6SbfsbpkRKcgKqhThZiUqeZ8
rtgs8n19JOUiwdjpw1ktMl/ECMQlhIjFtxT6Q918J4jqh2k6Xio728EyJpI2tbJH5B1sLAeD3HWQ
wSzcE0+7Ju8nYQfNKOeC5B3GN3bwvg3JsXj7lxVu7S9PL1vwF4jWUtj9A6mDqkIlgXMVAKulbvp7
PgG8LBL2Ms93m/vjlcTV9exgDLvSO2Ed1hZ25JEQIHAf5tq5Q3f9alZulbmwDPvzB0Mz9jsJgDy1
sPNNbxDft3GSN3KX6cqzFx59qS+Im9JzOJoFBpl6x1MDSgw4adld8WXVMbRIR8L2a98Y5GLH1gWb
iE15lvUCqCf/9sB2uF3RiU0y3jTpejEVVRfNHUYeTeywU6HTqpc74hNGu6pPQ2L+ox4dDW/76qgL
T7nHIYmHafkboyoVHWZ9o0bWDwwA6Y8UV2/48F1GZqypaR0fK+iXQCX+vd5IrKrd9BVlZcUROt3s
G+KX3p9bBe3s/Zf8i9qsaMnZPcsLAdnMWrDfROEZMOYapwQa6qapVx1w7TseGezAlSZpT7ebnT7v
/MpRg+igvkGepjrVMkk9xNREjJ9gHFpmJhTdUt3vfKJ6uLgf21WHOJEJQL4Kpvq325qSyEnARVmx
2zqSOy94+7WJ7U4GP6243ahxI0hus9d/wF94JzQmC+dDkAuj5Hm/GA+MZwQ2hGTzIPX6EVu0FfSS
3kkYW0pCTuQwGMBUBduf7cyQZqSbZDIQwRnj69ANWl+8gZlMTYgkSOdhNCC1jOp3RFO6C7QccTrj
F29sNqqe2MaBdq4YfYfpDc+ZGKO9ANK9AE89TB+OWWHHBqXEz7qf4RGjO+nbvOUM2Y/1pVLK7T8P
cwZY+FE3qTAlMNA07U61Z8U/CKI45/0FUhytrjJQkrIZeU8IxhSv8HsDJedegPyzmCa+xyeKi0ny
W7VRn++iDoxZuQ263qt1olLOqnFSxRvSluCOqILFhTg+yWAZxCnaUZNUTegy/Bw1H/cd694bGzqX
tNz+kyMZZTIIkUxUhLYgxDJtgOFwwsIoTTd6qVKl07rtj+xIKkcplYPHwhxKhXqToStdK6yoW5Ou
nn8Ca0hK4Gq4uM7FEBq1IGkhyuKcsp47FfiY5rrQbxddCvlxDTDwY7LqG68o0cuBSjspcd5zak3w
UJk0rD3XVI2jUfWUPLJTelvEbz6XbGZEb4hL1TP3S9pupN8adRH+uTJ/dkrVkNr671TB/KuWfmng
YHxWct77AaGzf+8Tm3UzKoVV8vYpdWr3Ct2neGN3M+yLaetP7myhRuFEpy+8/Hi5ZDCnXNuXrtpr
S7vIPrkpPfrgF4ROE7yFoc6VRSnCHoe7p73J6ux2mSM9y0LBhoQQeD1Wa2OMA6W2Z7y89gLga4Ft
g04TFv/jN3CCPlpUiqeWHeKnY03ZIFZI8YehNQHK0RW7Z3ZSXgSJouiDCvpIfKnBFix3OQ5bS+a/
WtGEhge+ZgzrwEUtrgcqwhSPZuRv2GAmSh6Jcxh/7rNxL3xI6krpF9lRmKhPDzuExhz0kt6+rn/c
hnn8VQ/L61XT9YBUxb43SCvtbPgOR2RDU/Ah0JVob8+VhzaoYzoaN/ljyF4nxTdrGF364Msc6MVJ
BE/OvEHCPShdxKD/q8mLObdjz+8lUJiTwdtJgnnhAGyxndhacSzxRIpQdXuzMbdfUYYBdCQ24oEW
L62WQ0LHJEe8rEBILao+qn3/rgSBNzIxYHjlk+IJoclk1eg5/NMk+4ElD+rZtoazuME5sItHaMPw
OUqGM94Yoq+yu829SbCaQyNsQJFne+7b8FrmK/ucWLERwzkGifTO3REDNwjk4dtdjo04H6WqjEX/
/0AtGfXpldiMtqyYDDbtKLdQIWCGdKL7QzR3eqAuEFuihrZbAT8QSv8umBsI3eHXOb6Sv0hn0bC3
WIzKF97kwfAgyqJqgKvwETdKjXh9UW7ioNqjS9X+b7X8ryGy4HacYAeZKacKkfMetyk2TKe0kkI9
VbTH0EyqeBj663RKGhN1O9wy1j1cGH490WAaGfgx2LEcCWtSUbSoflpHdPNR6k06u8QG05uoDQTu
w/rp2c9OVR9Qx7uayzx2FUB7LEraAq2lGh//qxRrBe4xlOCvmLzX6EDRxTDlakzm5dtUNNqZyQ+6
9KfLyvsQq/tQuTJrC48vPwVrQ9DldAPXRvWOfkulMn9tnUy6uyGGVf+t6ZZnpQMoWWb7h5CqXas/
Mzuk7DnPERTQ88TRblmelk7cV6lAElcOu772BjLC79QIdUbeqNmP7dSY2owdjQCf7WOQFuZuDf/L
6NSNTFN+u1f9Iu1n0ZRTitNE6WL2FdqPa2CYAWM69R2MmkPzf6Crz57tbwpDF5x9ISVNW0j9T06b
7fDXcjc/yeCf6DuUVhdYuo8Ws71kbJH7jnntD1NSnt76yZjHX9nRqVa2BBfm0upc36bxWwFZ2gur
wWTR8xxTB7pkn0M+6cKPFkYjk5IBa7Sfz7CHZZUoIWCAY8wvpCQyd30HKD1DiPxLhqailGkn55UL
mIpSqR3YOWL770Vb/IzHqqyB6LOmILlgbCLuEWBajMugnqmwmjVw8Z10EIWGY1PTmKz3ba+zVlfv
Jw2mJl3fkZcX4hl05inTD6KTfJNuJ+A1khXmOL6JQPsJhC30/v7s3MWMvz40Qk2707U8lf12/hhv
7cKhG8nE02M4D5c+i8YWcy+GYeIbSfJfSlq3L9jnv4+JOFqkKLsKgMKjhxFTKSCIpYMRueJE0xcy
IVMwCxyNgA2sD8pF9LjSZc6ShgvrgNFRHNr9T6c2OY6M4pNi6xDCNqdXtYYibf6MMqsOSgTbiDqB
l4rvq3BK/afqYPM/qF0weUA3idjy+I++KXSV8q1ti5YN/bm4x+rM3Pz9Xomic7TkhVKMP3mEb97q
SzUqItmfQfsWMC2+vchvaeQ2fSFHflJYjg6GPVQIom6kElzNvughng0sWtbGojPFNAwpfK5KXamJ
Wus4P+Tcy80gOmZBkE3iqD/PZutGsNyvn4w6/O5eft8bAHp5UvWcahOau7UwXUcN2njxq3tPS0CX
1HP7RVzmO+JPgUM+qO2b7Bh1LdL027PtGKytGAxYD+fkYEvPCRm9MT9RplR3HhDRWvt/PLqnpTP1
NTYWQZUsfGL8WkDHTWPimTCZnwjggrAYwjUTpze0Zm0M3dKAgL6lXq7CEO8HqmbiR/ZBdjQxHmE/
dlgtgytuhhQM9dJfSzWsq0vPTnP5hI1fJAGz3Qo5EhC7Yn+V7m7nHpE/OI8jbycrvMTMI+pL2MVR
zswh0e/Q5aHUVXRO/V33WMyEp0WXwB33vY0IosTWS63noqbYDAug6GbWYZMV6iO7JKW7PfgqhdM3
nLyNoNrYUEf23GZ8ByFGFm7HCr/gJbb5ZFHcbx17/xE5u6Oy+cgLmDAzhaOc83AAHwWjXvQPlk4O
XFZ1oH9le0yP/nOgcLTzUePwtuRtlEpGt751vLWegdhQltGgGwMfZt6fM5BUZQUGZPChjFuFwqkc
zZq0ACYAr/dEVFYfFwl+1r0nQbia1nXajOZouKyOBc+bmT2RsqhCC9PuGrLC+3MWxNzbFP5PPISd
UCKhVhhYY2wG/AiRzncZlq5XcVhAKNYC8WBK14Evxt+ToSJn/Tq7PONTff/iOAwOszcfQpowD5EC
FKiyihUJySAEYB8TYpmBbbi3EZTVRGoGZUIt6mSpbi+DQ5kseqwJPbJFIJVyqIKjiaoHqluy14A7
xoA0XnkRo/okJoCF/liBt8CrdzUsarrZ3xxTVCyHN3jct2kMW/JJzZmjZAC6JBcdyUA9iMzr+UsV
X+5WXlE6X/dvFyvDj6UtcH0YlMvMKdxwS7EeKWvYf22I0HJUMd5FKfH8uvf0yS+1cDgZFPg0Xa0f
p+quEmAIFyhpqNgxPVmf+4KLBjJGixHWNirXdGK6X0zFOdnQqI1mJH4zG6aUW1Ck75QzePO602si
8/mNmzTWO5TXQv+bgQknfmM6K9fKOfAn3T6NsntFpcUv7otaACbEHRZEfquAYfDvaAQkq2eswogq
iFniQiG6WOiWA5ydM/6pmXg78/sh0VtP/4hXrWBh0o5v6H2Hz9ZhJCSg/ZBPUaJYUW1x87MJbFFv
L4YWW/yQCqp2FLKQeYKbUf01cynscLh6VHZD0CXfn9dunbHHolGDQcDAEZw9NF7nteK3Vt32Q1Ec
424OC143UkUW+k7Xe00adK2rLA4evRcXlPHSF6d+jIRWQjHhLzoHEa9kmajgEYkdAADb+aZAGJKG
4KPn2J9iOdCS1NAzu67QGgLMfWe4hQo8y7DdFTGrMrxfczqXKCipWEM45a6i7tnZ5/ce0v1paHhz
rs6NeGKd4HwJkYf8P8/aIpz5+IoGv5E++rpDlknHTGPJaFuU68qHw2ZVfESh2CxF0PDYcq85sAK0
XAkbMIXeWAXQxIE1tAnpokbQb2tjf0+jIJQ9UiyNUh1dVD2YNWSjCCUbtaAIIpSnOrslMviQzUeJ
vF6FPVjKXFqDIdLOCMcSTjpCrCifSvkeRZ62wseGqH3qKtpzcrKLifCQJFdJIvfPefrfCSjO2FSx
LKd4ME1Zu8RBC7vVdzlOBdFbRRf/z2knnOgJzOvALX59bffyKKwQnZn5GjrVFutaHOSybTq3Qlvo
ND5z4e14An+AxViKNRIT66AXdnr6I65vdZFQ4oDJe3au6+ecYl9eR7VZ/NMB1lQpLjB4hu3tYILS
OOQCKCTvk0xqYUIjPLecgpRWURvB37bi7lPsFv6yM71yWsYDilJkcWWr0F7a1wtj44sQKc6m51cs
cNv4famcu6XqqfvQWVz7rDKXDZZZ0tokaXbi9HQNncVYsP8Ja4Wx36lRm39Pdi2s47Urz0Uz4oa1
GRtILJbwN/jFgDx8N45kLC6/mBpBdzneDipPuUCoLGrWXLVuRs2mxFg5FF7xX4rtqCCXCwWd/Q6K
6juVzCoFjvJTWFxi54LUwbyvuzFVktAP6kehngpi6d9E/jnDCENAqpJm9oZ/+v2Z5MvHokM+Am7h
f/exXRdfyGbDiX0tlttRiQpP56W6N+tUBFXWTJ5Ch9cHCY2CAS2FIxzlWxeBvg4u3cw1RdZna6Qb
6IFI02NVnULZYYZ1LRJkU0LghT4q87yUWJN8g5HnYXZsj4kh032SjsuTKgg+/eZoZuCEF7OhnBQx
abuQpWlM436vfC1wth6Anb3khv8JDapGgF3ZRDL62eqhUJ9iWUXmmAVLZg3eT1KmBt392ngWZyBM
1qngzS+vm5oy0DgjTRR/GE17U8JPu2gnJxsL9vmfbun8jlnTCrrbBUV9Go2JC3c0P1pj2C1/fzVh
G0wV6VVzZG7542EFvV0i6s4LPZYkAdOs4I80mNUQSiH29GncmEDJnV2RBxnxYwQUIyj09u6CsNcn
zJ2cdSo+UaREI4fhCuhU82lS0DFGmWjgAfSW5Ica6/tdg3L60FtxdFzT2RL8YYxjRgGt7hdjgSga
MQCoMO44K4I55GOSWTz8Q9hjfOERsz4wg86o0aOxChpLkisdJM2qRR03//8vpSx2VhpUEaBvkBlu
NOtrgq8TLWtY+3dz6cS5aze9aQEMMoXRW6UIpjd3HKP6NYWkHiqGRHg87TOSybeaPfJiJxQNH9Ju
Ja/HeTNhg6lCKqOBqb7XJscWvAXFlGf98qc819Ot2wSbMMyLBCCpYmPTtzJ7jocGTd1EIsQXBIuo
fcIlsLP/4zMK5xqF/d36R6h8WPdB0bYfIE590xVwPbOTpgDo+AsmqaZ6aosnro0tBtphHYBvD/Cq
0G8Km2AibzzKfweVtOiotGxeZeyU265Q4M8KhR0LaTy5fBfv+5pbETEayNiAOIeHj+cbR1jHzpLj
sqOLuSXTv27btnpr+aKfhPD1U7yw2zHO9HSFefxOEnFXRHeVC9bNHA6fEshP7fEy4UGI0Gzc+VD0
MiqxwZeo058Pdlufjtd3BP4YCEqVI7RF2iALlc1lA0v72/A1AqnvWbpAYKiqZ5H0ublTVUUgqcVP
V4dlgNMTvS4+7jkb9hswMHNx8aPqRL2KOHMV4y2BHy3fYrX9BFg8NdtVIQoG3KtyFsDSOmDEi6Eg
thEQA+CyaxXhQKYPvTrMPgnfmF7OC6xsO4Hp/Tt0gwKHB+zo2hNAe6oyjhcofFinNT10mpPjiJcJ
OJDEW3wSx5ikKK99TYb54LMACjr9qFH6Y7kWBj1ObwyUYfwrZ6DxUo4UHo4kdlotkABlhCx2wT1o
DOVPHZ0x51itdXXC5/DS5m0r1VS3sm/BYEBL+8LlZD8hMHxcAgF9dmyo+B3P+EQ/rCnT4DF7CbWj
vE+J3hz57wBUozqMN9Mdtt+sYDx+hxKFwLcy5ErLUOyd4rw8ws/ZktntiiaMTBu/lxPwH6dr5F+o
nKUM7tM/Vrlc42yjmVx2dK+xDFJoQMLE42qRR/N4ZWLy41eVsBHwISvhHmSuG7Yp1dxbHuJRnsij
qB4W0bTxWkbb9Z3m9OGcihG/dmYAUE0huyXjxcDic6NF8i1QX8IhkecoG1BWHRbD9IOHnb/pUyzr
Fm9G1ntIpldsk0PvEa+LQBVsckVExrRXLe4q7hyRxV9SABs1SLYrBSsqyA5tqIWseCHMtNMJ8UzF
WfIiEFlQYS82nKsWnXn+lOIsSgvsWp2P3FMZJUs4leWvUoIRPpZVKmdLUCkCVnY9NhPRm+Y4+SeO
GaN1b8IOfgcvP3qVY1hiPGWkL+CHvqmRGE8vMYgrLa4SYoGNPts/lLDsJ/G8RfwLQRgOXuUJ4AgI
+kEoIrHgrHVuGweZAfjZo8eEcHAQPT+cmG8ZeWhBNcOsHfwZJj1dNhP2ssVTHiw5/iC5DYE+vIOC
/NgytMHliqynXFzVB4u+g3t1sIrVLhfm6dALSZPbHVMoCUrpJOv8LyqTLNAv0gn0T6JPyEt2KCH9
FpS9YdB+VREqLfFffQsZ40T7GCtok9ds0NPaMkcl76fz9b2xRQ0JGPmOCPFydo+VfklEbxC1770X
fVnBCST+Y1jOsnhjhj/Eai85hW1bzQuivoVgWSkw9jdpmYt/0PQTFBbZeUTl6q9AZ8hX85nl16gF
rAhUMtct0s+thVBYSvmG1j34JEzubRK0UO2hnOw64pdn4VaJmtdgSqQUbGgU4jM/UqdE+wIzbxcN
Uni9YXfSLWSVizXCmYNATPpSZdJKCPdcC/jpoFXsbQv7D92EEou2fozn2coyzggCegIWR40XffO4
z5pfgk2+AAZNCqDUQ+tDM+l4WxRAzYg8fGuhEmC018+JjM/klvlI0GsYjvygBc2uv3fDE3rJE2Vr
zvqD4QJVaIPgDGkiuBPH9/J/jUDIeBKjwDt2KDKgjyvi8JnUzvdD4BFSKpwokuUVkRc8ovKvgULa
nKBMm39cLtiZDTzAmib/EWVQZYTmYrZD2ngcwPetbC2Twga/egFDoILkRsaFf3lTxgtl/mp6jOsF
YLgJk6nFDBTceM5z9krmiti+aMjo4a8DAEzJFih78KmtPLZ2EhMN58a/7c3b5oa8D85kmGQkH61f
XDOQFauUsyIYgKtAnOYGdvSWir+Eh8X4b0y8Myp5yCAR1oO/D6gEy5dL0jcNSXBS9PRgdhDWxM8L
ZkL/kvc0wigIemJkos+RNS8aO6qQTvVWzxC+gc7mfIQUD1f4Xg0fZhDEScS9sORm6VyZK4XpdS6h
Z6g8sRBAiwR6C41UQnHu1KQNEaPLrpRLlz9e1tqprwh3doGep7Pk+C1+SgjEndWJsAJUHppF5scc
PlNaoQ6etmsA5GvHNWN3/yDoLci1SpNNsSl9N3ROJqp9BjkD0aMIqTwJyb6smaSReqRrKrpXQ41n
E1cFN5VrLr0/fpHTimXy2+k0CNWnUjCYqqLkRnQRfvc/BX444A/05SoxHQIdOKvpubdgsSErMDz/
eRT6FgcxH539OJYVi/x7vpzq2w4uDf0HSrvMa+vAKPhl3M62ndpkfaKG3eyq5RbKcZCBRbr9QM7k
scfgrH1kOgqjcJO/0plhxRodbwGnkP++JqIGbkWVN1Ezh0yucftyYzTlraBvdul4LhCUZ8DPTB9v
KraVxkNTJ0ArHusuCzldrOBlLcYrLyOKsNbFIipXTNKx7Mn6j96znPqTY4RmacMXFJA3xCA4f0lm
53h/8wszxNHP9nbtgLbsaFT6j9HMUmaLgnly/Za3dFER1KiHMkjm805GDCjSjkUbWlmDp0FUyQEC
XxulfwQpV3REF9d3fonbATM4q3mqoQFW5ZM12pG8BV+aSO7ntUN18dJbgpcbPO2OHlCdD0A+pcPf
O+nAn2EIm+4+WVfmWjiJJd94+EdGV5HXsr/V12Dds+J8+bCM58kPpXCPDMoThfgQDx7ekPpgtrHi
NoaWt8FsNQp1kLXZbe6VhNiFoF31mMMwqI7Cvdp0yWuMW1ruMNzXFYdcWV3FKjNpjwqBTQIHjbjE
nh/MtIqEN0Jbo2sfhCNrr6an5T+hly8h5mtD9yw5GW8qfsARVAF3LL1H6vjLXLDXsV+2LQpxfxfT
dYQOHoyBMEQgOgWu1PLkDf6C/Pna+Sml1aQZVxeCC+MHFEFApfND2PnmJ/WXw+2E7L+A4nNsLg==
`protect end_protected

