

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iaGK4Vux1Zzm9gBS3KKNmBXNdPq+lSqE3Nnx40zW9JpQDS5U0+JlSB5O0czPvIZs1e6N9M3JonU6
/VRFISTQHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hnTIGD4PF052NtQspkoD0qYNWsnDfk/EZli95x6g3PoDiWDo2i9hfthnklZPOTwcwwB/on/PGVLy
LOGgor+yT4ZX8UGtoSmScYDFDjshoGWHhtXrHczoGSF01e42zFHCzF3p+Kqif4EYEFLVI0b3qWfo
JoBwVA5mSGa7z6eKZ08=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jM4x3jcOa6ByCa1VWDPoU4L7JC2eupLAavYhTE4GTMYrnvE7xP73g8zjlwq1G8Zy1ODZ+0DDopVA
JY2gdvefh3SJisXvlbuH55643svFB8C9ZXe+EMovXErk8XGGsVfWZZ9248m2dlrUXREntbWGdORb
Fvho+MXYXuv0DV2DKImT+u2TQDacpvX5e8ltSYsMmjYxEdkZrVMF9C544bgDvuCE9PfD8XjA3SZW
m5oOMSMtDQabvtrFCxaEG4NyuxA648giN43WXdidnKPUkuB/HxDMEcw9NxHOVNuLeVs7mrwTNW8a
Y8nkGhyssdB7pA+UlWrXAfs2U9Wpi6SjK7D2dg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l1zDcM4+iGcttYyoR8HHgtSyP4Fiyy45WEsaODDzemrDXcJaURYpyLa2UgO2HmqSNgBK4XdlSO3S
QC2s2wdlVLq0nr6twxtavd0Mc90p3l2akMlkawzSfWC3lR7JsZexWZNEb6frZfXhesr8/8i8wphW
9oH5nUnhDJDdlXi2xk0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pHbCg0c3yWoABGhh+X5xmKdWu54K0QNaj8yiI7dbYcl0s74Nnt3O7DJj12bDcjZRfdRoiT43bXo4
30QPK3Jr7E41USUv0QfI981OyCHaIYD9DzkFx/42CQBEOSHNBrRTW/rge+4hugPE8z0ogrEZGdei
kB3oPw27BqROJcBQEhzDTOz6PP5L7SaiUGBsXkKo2TeQ1sLfd6VNm52eUhSewTFcPcdSylZU9gjA
/KlsPUnl2PskRWTiOzVvvy7q14ROz/8yTOqbBslSCNrDfBQA/bwCsE4HN784FAGU2BIu6GH0W9gV
ySlMw5kMiPDazI4NmLxMcJvTd4Vi8xnRt0T8Dg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5728)
`protect data_block
upmQ7ofiIpIjuhb3vrb1YnXSrcQjXQ0HrrlwTHf5T5Or/M/EOBT9fhcipqO+vhuPxndQZNGW0xsh
xFa+S1B0K1Wme5Jage9d5ri+RrtUH7MZ8bGeDdJk4a5Xeyi5pvfZFPOnZ4uAyMlIcnI7dlrzcC0U
uni7dnMOMQ9lun3C8NV1Zr/NniIYrLliaYvdOLKMp54OXR1DtLbxTJOQe/wTT21s5vwsnBYheY7I
rDS0SUJpxpcuJ8LNsCoULUIFgScMSbz+qJx25EJso6U1/Id7zD37hoo54iBzPHaTjNPDsSpo53xQ
AWzd27l8gVY68SrPb/3A3BRPb6lNxWH7iADSKPdnGqrPqtVqgC5F9PmNrqpfmhUu+RDb8RnLGjzz
ONREyLXPslj4GlR6uKM0jK6ZtuaVYK6hQTY77LGQcVREAR2fQX2RLNzW8aPF6msMnsjqCkN3d5vp
OCU2fc9/rxxq4u2fYrs/I+MjUY4AiBNAW44cDFpjyQioq+z24aWGrAyjbsrtZoTVEhZVpwwfh1lz
u0kKzuLQSH+u8cLskmPDkU2LfP09aXVTMi1J94cgXAi2/kA3ofCA+8KLf8K7Jqlk8ieBvHZ/65ZQ
6V8dnxpH3GYUXBZsxEQsZj7CutEuWBC41nGzUrAdh+gBiCg1QA7ED9UfKMGa2yTapB22p3Su2rtE
I5aA/dSJ25DLZ3yR2nAdzk7SIIDZkACjNTFgbpG2RIVDuwzYPdTe0RcP/d2q+2bCtUH5P70ivxQY
IIQd8ijXoE0s3ROqfsroXdZDOWPmCx/OmgrD6PnPJvKw1ruKxlUNnpyJ3J6vC7o+Ujng6pnphz7U
6hJrSlcEFo6dJYypcdkDImVxLXI8F0yNsL6/kpg+nuEtcM7aF5DzhkJZfz1tgShpBqvf8LGPzGLt
2pHAJwdZCwAK/CkTp7Ggm6Yw/WffH+hzL/qxqrcqf5Aaf2h7NnQ+bGjJKeirARIyoEl4T7r6VnDg
BVXGyIfJBenvM09hyB+zxjJZBIq4EVxtOGQw7AKzgFx33YFU5r1izoURA/rWUKimzMAaU0u1SonD
f3SmrShscxzzVG8rT/S4hvVGLVbe5O0xntoln6i/sE5z5wNyyE/K/TmLf6+FfhLflD9NZyH+yail
4D+D65eA4efHMZANh44QGUuCVv7mVm9dd7qm2uNvwcUHkc+BGUcZFE70VpfZBlmZevZBWuzRjqdZ
ADb1aOsulWgC/fxEY2chse9HX7EgfO6G6NzSHleWP3WaSMTveu272BD/+U1L28eLfjQnAW9Jyg+A
iADWtJAD2M/IeFxMn16PpQUy+kocHxH2Eilb8wk9+rfiYdVYS6URK6iVGsrQM+NxxcxmNjM4ybJ7
+mcVoSq9wEsgJKeT6VW4aGYQbzVSjkoF5MLQdB10rVCcmWBOvAmRK+e5smYf8oPMDSuXCzD5hUF3
SaBnl8mKOBYWva1V60mrLbqNkXtRs74MaAPJjHAsCvUdvWmyJsm6OirzraiBIOijyOQuF7EZWEOw
LFzyGWPPdI6GdEgynlN+dWhRyEi8EL+pN16zwrYFnfYBz3+gWgPF1jv4bLQSLGp4/5hVE+e7bN2V
nWusQQLzSRDxMmsUWCh5xiFFhlHu3k8qrQn6s9rcaFQMjbsOJHLkRyMBgJp9hF59I88//F2pTKLF
wsnnt4dAEOGVpWD/HOg4tORgV4AeD0KlBpJqZ4aDVcr7TynWqj3RvbIbIzxH1M16zxZzr69SrYag
J315tJbzxldzTdDLpzzBcipuJD815pkjDnAbYJrztLLog3bQxbgp6WoVjiUOX/6d7RciiDkdfK74
L7gsc6Cg2Nv6XdvWpte5DSGAuyY4Q7V2t3vQlcpSiWRUtoXDJAADtr4E/jjdGsq2V7j99gFUmSXv
LnHUtHhZ+NThXu1vwnj4+Cau8EMXOb6L05AyFBik64/gx5W0sKLvJNkj6VeT2muHOxXeSXvgbDRe
uXElgT+3g2/S6la6VSj4GuelonaoNkzvXPbSdkbnR281QZDfrXDsZ4deyYbiT0yePQXFEiGVowOK
c8tlD5AMSv4hoHvAPNcuWrkKvqRy3do7bWXNukvLETSwpM8gaZ/SDmwn8Lc6e+CT8TnJ3d2Kkh5Y
DA/4fgZY4647RSYv0Go58KRrCthBphvApw7KPCvrM8TkeSbOEuN7jUCb48B+QR/tt1YErHIbd6lz
f0RoG1WXXOwcZwSX7+Ct86L0dx9DJSGIh/e08c5d0xwg9tkiECuYU+NkaZccT36Tm8A21TqGN3+t
9tNWKumjEK+5PPfwApIY5GrPhqwLGqVopO6mlwbiIHOAmZy31Yz1Ury9wOoLLV8gBS5oqP8G48K7
DhgWOUHVavlM4zpRr/jT2Ei4alxq5EMBc5sILLKxMxO314CdyF2kc8z26dD2HZgcHgKTPDEXI6GG
/VXSzZrEZuKnmoh5/FONkameQ2fFbUhx4zQKO34H+tiseRlhA6cgYEJZ5Ta6Nt0WJbFccOPGUosR
x3M3InHtVNcw52qRfUKzWjft98SFOHyvznXPottzizi/r/CVWt42nQrB8O29D6H9D1neDUGF7zAC
p5vIsjkLpqvaXiBhd4ylYKnG3JTnFNTUMCTx+N5JXygGUXKn80r8miQxBfE1J3P5X+q8BzIwqSba
fBXYdQPUwnKi8/adWQ/T6WSB3SZnMfP0AJnf7/mZTPMTsaebU/iBYvmFLzeyQ9wWMHgBxA5eLvX1
kMpTM0piEQw+wWukoKsJSna3y4G9D2B5Gz8+OTTTMvh+LBrkIvXpqf9nxDbcVyyI9ziT2UIPdTh3
TGgXzPga/6/GKwmKhSzZx3Z9PKD4dxROtsJGeIFrv7HqpQL0XVi+ItmY4n298+XuJzJ8/1glDIbn
g4K/G3FmHNd6oL4FmiMcHB+IdsneZ51lFScBa04o8P3MxQa0YSVR7ElmhkWT2uiWlUo67almAKM4
64y+t1aAc4IfKX+eLu9UgIPaCFqxHnH2KTW1U18ucECLd9c4/X2jAtG2vCHAxrsqAvpYXcd3TYwR
AeoArnTf1YcTSFQPI3CgcaKYUAuI26Nw8kg2e8UeXUyK3E1QSUJVp7o1eKyfOFbGkgAbtCvts98n
HH2sgDutaJkhW7SXHQzsrx0sHSy4UjoMpkiH9y620geUGIwKK0JhXnw48ZYISe4y5UBtCcIe6bia
5muNbUTfX+X9WrDL/Z2qhKrBb4R5dAMcwqwiNxn/M02YALFnropwCKrOXGpDA0VDEl2ib5zhAMOD
a0Gn8oFSZuzgQ8iUNKssKOgjgk9/qVXnhHwJvLTuGG2l2Hpn+lfGJkIrMK4hkge5EEqlctrshaIy
Unw/YjwTeTNGhOf0jeKptsIgFW/eEkfYnd1qzotZCjzyf7xRqWXry2l6muAAAoLPkQIJUNoCXNcX
3PN+oJrUidiXwXUud2nBxnrCZSAulk9co/EnigUh+nyt+iV0tHphXIJmohszKKrKQh11Qna3O0H1
B4Z0owDnzaAtemMOlKN6Vqt/8bQnSlPxzDK7p9QHbnvCAs1/qDQ2wbtuT47zhW5eaTk5IrtSpNuh
MSfhs/ZaBGeYkDY8Nyf3vyAFK+4pKpJecdtiaVQTHdDcq4TmAeq9Kt/Bm/acchaEOOj4r4+NVfUw
JVoI1Gv92y5VrW2LKfI++k2jdImNzsCyEFsFZmzK72i5bUvjM0z1yR/dUiLhqCwIWOpb7WGG/96j
y2JQW9zqE9aOH9Kmt2qxDg8wGkqHTRFP9npa3jMjILe2f856ppxI24d2XS0FBF+BaBC9OgqLCOYe
dw3gR6thVLoo7s4AoPmzUNCz+8uK+6oPSSjLSoKDkGPC8D9CcN/e2h7/Ny9Nh1FpVDGwPQt1RFBB
UH0e5tmolRsRPZo2quTZuKFpk2aYO6FyF3dRUsWSeSLv7/HYNTxDNlXkwN+CDO9atGX7eWfcjEyw
ZImjF4d/XR+IfGaGRuWlJ1WWAmG5O/zmv/rXk5WRIBzJqqKcF6/Op7jgFQycWTOeDp8i7GKaC0GV
67Ebj0vwEHNQeOmilYF3/vXhtVcVqebE1ALNptZ5WtjEcm16RuKC5hivTFqNqk4+3iighi/d3n1Q
VM5OYZx57CUtGzz8Z78on6BKwnMCVt6O3SyRrsGL873sfhnGVIX/nhThobEXrPcpcmZjfxSGy1Vo
nzu+4BtYETDYuzueDpzgs3BE0PAqfozPruJmHXyHaNCRN5QC22C+oIOc+aUzDbUsv5fqQ5KEhs5+
IagdMUpDXsmVPWRxKjer0DPZhLVbmpL/jhuUExtv7/+QiCDKyIMGk29B02aCZWq6GDBE37lwgVVp
4dchsZPQzhXtp7IMr+NdRmEJHXALqEtT58+4ZtcSLICnicSpXvyRCoPm6GGsGPWr6eizn01XtLyW
D52S51WIxN7Rz9g3z252Csd6sI9TNQvPbgJ6+rUoN2oH9A6xtjfK1LFt2I+eYb5mddG/hCo9Lb14
fATRvma/V6YrKafSgqDesUoSR302fXSiVznh2RNGhRnd8CXFT5xx+nnXJWuRVKghSlC1vvBLgkwJ
sUtiGoz+NlnLz60peay9Yxavz4QeSEgCxvvpdb3co5WMyZuSGEb/CLY+2O2MEcfebvtom68+jlax
kCF4sJiv1EYKGbfmatA6xP8cKLdWs43nOkhnldsZMvOXy5JH/WgdFyewQNbZIhMXqnbtVVvy73DX
T3+3Rky0jGK2bSMUXD9jgz0LI5Ty0VSRpYIBot5cThvnOZeoFK67k8fSPFUK+O01PGYM55QDxwiF
BAHxcnWpew52zrnB7qCpO9vMaXgso41705EOqQ0UR3odpeoLXVzlVn1rrrPL2FZ7DzkkrIPFTbmZ
nt/CQz1Hp+/01oN7Rgjgd7RagneXWq+VcQT0OYEq1qBOgCvphwtFAPxKgUFwVbMDCu+oYe5PD2Vp
mGTXgzqEwPZZ5QOqtrnJtkHZBnpcqUVlNin8Ilzxn1HK6QKPtvyrolqpyTnUuB1gTxjADma79rYr
cuFzbvBPO27OTN+UDc6Y0bgsNfjRuKwUA6PcNzW0MNI4K8T4/sEVMtjcWPIeQrlCZVfvZ3Ww3rAw
5QwLlToN37vlzL9dtMePvhZiWqYiHbYUnQ46UuNWYGml3I96wV0Dv0EJXLtNRa5balazXBHcfz7h
8BgNHVfLqy809DdfHMRyD03VUlLg3Q5UNZU6J5SekSjKRiD4sXK0Y804JRRQPbji3UU49UrQ2d8N
e2yzguf5Yzv4xtf6S2tV1ajA5HRpxISLE4Dp9qCUpih6LaK010LbrD9pt58UVff68xYZANxTlIfn
Om2qBY1tb1EnrfdqUB8NR7cyKMdQyTNDRjaPtU3TpWZb9NovvyuOzNBLQ83Kjnr2vL8xhNhWma96
yykO3iCm2whqlMJanx4RbLEKCBTFPCTgWJW88fLGVRdTsI1/86r7MGtwwyXzGx403QVF28nUBxaK
bwRWPtKsA8M359n28rrFZqJBVWbx+jfAkpoKa7luEjGuoeJPtSIrnFRtnhWcFklR9m/qyjdkyvhd
dIjo+rtJw11j2uUNpL2lRiXAowQ8LJorwWEsY8ie4R2Q4yXqYjgAYu0GjlWv8Ls+QR/5QvBebYMU
vx76aUPEr5jTHD3ftV97uC7ARERjxu4rBYKELAULXOkvOWYjWofpswyUtPkjXy9adoGWndlKUAoi
/Od+P91dB3oK4Hg71dvMP1JB5C3bjfCWlS2DxUEq0eNXCIRmFtBJt4FyWIkBCoCviIZjYuzrf1vw
GVr5y0t4cjNqXCUyjJ54mT0Rq6yHjlGjVEKIOc3pe52MfkWqKkMOmniad5nde3M2N5iJ1CE2hws1
0RbiUprJJFgafRcScaXJZWlHXnByx4zAciaNGSumGsvM72iKxi7PuTai3uSvrD6uzYv1XMnH1Q2Z
W3poyWPdlYlM2RzCH3v9e6R7JK2CfN0mn2qp2eoearHQf4ha9C7Qtbv6lhL+jYKiSXK+oSgFmZYa
4zBLqD+fxZTcS3gaFTt321CIvD5qYgLDVP3nQTDiIwgk+Yti+lmf5UEfbqrZZ4jvI7wtQ7ojT4Er
NVYjl+gCJZwKkRfmei7GUpsAed7CmxJFs7Z/wlCcxZK4fz0KxmatKqlvdu+KiTRmJFFFMNyUAgj1
PfmB9Tbsz3lHVE6SCNi3uuEXXsQVcktPlDD784wWwG54dMsqWGt4arwV928Z+RoPWCk3Zo0ad9uT
ac6txCFLYU7h6lK6mxget4L0SdC+oLNkMM1gshL4qDjT/Rtt3MHrmedy36+tOro8wlyHKEhf9CFp
KuiOxfWelaDw1im1fTT6G2LIoDZhz8EYlLSuqrbRuFRVeSf5APU0NvJd+iUJlc+zo11BKHGd27xR
nk2FLC5cdL4ya+pVDTXmp3SUfW72iB6Xjoz67m1wymmJlBymE48MeoXubE8RiyO3m/4SsH5ePew7
2bpokAUkkTgoCPx2wxCQ2JqY65UTVdUfHmLjUrIGe3UZ9mPaZKr6WMAXsNOg8kn80p2GrHQ8gmg8
gnvg82oYX/rD9uKs85el2TtbvRMK8LnF5141rYnyroBsLxlKplRohBtpnp0lnPuTB7lMbPr/PhEv
+dGxe+fMbepb5Ra9N2GVrypiZdctISmZjAUWLaq5FLyGs5x1yetQ90aiJQB3NHOX1ufHnJCONhrV
A3jVah5VJQ+4VF1FA2VU321LeRVQSWBjXUpdPusc04SymnazzocWLuKEPb7cFcKNABTMZBYAhbZg
YnFs8O62z+nZR9pRAvAq3O6l9Qz3CFXVS0aRIHP2vJuJRwq6QwBOYgXw32NHVCxI18nDdrERxy06
fcWhZLlCGcSiBtagnMAmsQaETUbWtNf4ZbdaCkjf9FfWk+Zpl5rCniZHHcvTV1ztso/Z7EcrbXET
Zh2mxDu4wCAC0cp5ZeZaxGIEgK9tC1jOEDNidozFRGltjuwZm+Pzfn3aP1s6PLV4TlSwWOKQrkWv
wv1QnbFJHIIf2IqiOpE1P7PTvY6qWCTmpOYSglfqGxnAMk7TErQhIsEHix+1kntdcU2e6Y6IxKLB
tJUacSvoFTPKJCopitHv3nX1lCaHbDBofCQnzPSySwgmsNLkVK9o0tYNkk+jOMOOJlDI+E7vyMun
Wx6G6jD8m9f2QOZ1826dQILJnRvDio49wBW+wHi2cYZacvsJJiWJMvSg254KRW4d24HhwQHfAZFO
E+44O772q4UaSlxUK8Y2za3BpKAhFMTiwTwb36ydyiK4D1MVYRCrg09qGClLAtOSZSULMKRLnaB5
TmbwO0cpwjqEWdZabXbxhybVEseqMPGZd1Vw/bWDQWlprteMsZ7xXN55TgrGoFo9kOUmfczzdtqB
mTz5nj65nXQTifFfIjNWPQGoXoC2uJBcnlApqV7FYDeEk2uWedoqiWhwdMlcpS9KRmQPQybEq58C
220rtZfv7/yAK1Fg1mxi34arE3H9044DAotGFt7tZs66EDHpXiDov6iefgSC4pJ4rCyvBW4KRRx5
NYIpHUynd9Fjn3/qQ1n/1XT3R4XWNOJ0uUbgQvNuGxiNfUBCBp3IOSUlA3+DunC81rPgis5TboKb
XHHUzY+NpAGDED2sERA31nUmOoZ6gZAZ8LU+AA==
`protect end_protected

