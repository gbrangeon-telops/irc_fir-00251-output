

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EHhlU67zSXzve/de+KpY85nXXvMNuZL7tYgf9fn2xs2MMX6KZ+NkxxVYV7RC95SlNzgUt4DfQ4/9
3ul1mLnDjQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UlAZFSxNoqgvPPKliBxVt5c0coSpd2sh9B8mE9L64FOLOsIE10QbDZBGLO1c2gEWIwuQ23M7QvQA
5NLCK/AU93Cer6u3Y5Kw85Zu7Q3cTJ6gtsPScNo+F/wtG37D/TBvZy9QIxLBvCRLOZx77GL+Y61M
X3HQ3kaL5tpBN9LRA7Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BhywTGDm5IJZmP+63CSoL/TDCpGJVG3VkCIbV3f5gGTJ6iLDPwvtFhhY8681GBR+EoOyUSMbP3AZ
DMFHBgscpLa8vafzBYp5kDkIAp6zpVke5p8WT0T374mfT86d/rJV4lUvVArJtTXZ7Qb2BRu+oMwW
4NXsxCdhgqbldJw6uUCqk28aEPgcbivrgwKY8foWfBnTw+EKHyn/oWDvwghTokcxfEnmhIMsR0T3
yD/98FKNKviERlHfn1BhQ/aqkW51Vp/q5U9qrKs/+lZwoRMsy8lRZRggDQnNmQrFO+0t1Oq/DlpL
Pzgpskdyam5KjVkaaUDiD9LunE1mnunv1fkvkQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M0G+I4o5qs/wY3cBNkJHuC5SdvD7yJrXn6vr03zDaDrjCzuSM2xSWnhAroxnc+rs8YiB5XG+kxRS
nfrpZghhDmt8SYAMsT5eb/ToWHwFcmxPkOwf0TCRf7UHox/rcVr0f6gppZYuBp8i/HMdTy7/9hVi
Jazk/jJ0qiENaXH3lhU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
II8O6ksX/NQP2v4t19inJMyzBruYXofFp7EnZduWuRh3lmwU4/uZj2tsoMzEFI9GURJGr6OGMrIR
LHPoTtEBaHFBnPNcL2m+mOF2hh90g7CmgF4J8nr08oNvCPZORB5fd/Cj4ujbrC4saBHdapCX/nOt
W3mratI2AGAl+T3t7Q0k1PLokEpC1hOrn+eLqLqV9hKaNBlW7DfM0Swj9M60AbHp0kL8sQjj6PfO
zKNcq6Xvq1JnJLzZ115Py+hhtw8g3az1/vAI3s/sf20/ggZ0t1s4m7+wPif6Tf6IZJCySXPmKW47
LjAxEb+MGgXZe5eFDZ4nbVPt5Q03mtQWzOAzTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6240)
`protect data_block
NPfvvz/xMN05rCdckeJthNvyFDlP7VQMCn9PVEKIQdaQ3zahxpZdV+Ham1dqS1THFkgT7cCBVmU0
k8CzS1uGHANiML7uqpUj7rCxhDWcqGiCnSLJJBuY3yTtXmUKCPxSRUUG5aGDsSIjl1SO0t53TI5s
+yjzpQfoa4t24eOKzYBEIGcw8WUK5erulFa1H2WpaCBNawsfi8wVYXlK99yE8vqhBXo8es0qjPuV
G/Itm1ED+I18ByPUATBau1oTfQU+fThfo2j55svoKSfpejOa/t/B8hjfY1CA1B7bsqqBaY5naCI+
zRcqkgzHUIo/TPLbxjTxujZnvEn1h+A36K7uAJEtrOKg9NEVSRhg4J6Rk/MJKm9d69Y99PbhJBrh
9TfK1bAB1PDKutE5KIItjjuAK+YnTt02ou9zh9voqHj9M8AY1GoSlR6OMOVKe99ENqPwTDlADftZ
jjh2YNS7tA+pcTw5pEG1zWN2CP0EFImsV7QDQDW1y7FgXpK86NeHM6fyMrNSR5yT2NaLwIsslfMK
FnsaBJqiRHRpcEY00yoGPzrE3Kg9lU1Otl3HjoWa+3uJAE4TSjD4MVyRuH52rtlIUSiRuocuO1Pf
wPo02neKD6Qj3waPU9IwHCgK/xREbZJ+xVzELSXoYXVsiBp7nSiGnigtlK0GyIA24Uc8nAXaG6mf
MDHpZHgbouFtK4BckN2LWyS5gjYFlvE+m8l+IrRY5XS+8ENjuNii2TU6ndtxQbi9cDK/iTxQSeRG
hspdLyfHpUs6ABjATR8zu8fAqAX0Ml3ynLbdizlv5fqva+qfwvKD9wr+N9ZB9HfY+xPPWZmrotLS
mIkkh1GEnOvnKXK8Ib4pBuR74pUBldH/F/gOHWBxv96RP2iJb86FUVfhinIc0IGZNZR+G6CfIvc9
fi5DwctiKmKjPSYHJLcmNPxvtzm+wYsUsJiJUSU05/iqjyo3mNX6zVVC7IGAmhHcbhxqARa9UXmp
73VhU9ISWOtQc5C9bPoo+3UJdsiX6/phMw5FTFYb/aBsTn9pHNRkUyhjp9G7dwAw0FxavyevhJbn
Ra2MluuTDKQ40iTHvu8j4aPEjL4EQ1mHR+eGziCS8nEmZCMBpypygqY7/CiV0k85E8D5vFFrepMS
RZ3WDkD662KY3XToEZUAhdfM+SuHzMrWwDbcleSkF0BkMLdrUxaEj5Z31x+4L2r/s8LQNleD5Is2
jLcOvzZJNXEEydOm8MibOKlS3x2p50I5+zlDyp2HWCD9Du43IVfFAFqGqgPqKWgQY3yrCmMC39xf
LRa4fI9X0LDulhqDy8qINgqW86/Uc2b2lDiwygR/wlgTaxg5FKIJrlhN1/fk7Q4sjOdzC61LNRwz
a+cEPVOAdNqMeXg7Oc0kzzMMXzgml3TGtfkyC17/PNsylsIETeqDl6NBSZaVvkboG0YEXLaOcZlN
hn/a0ISwEvZZL50VZ8+2ySaI4UMgv2Mo3gcz+T9XZy3D9wgQTkwxdfDv40zHK5j8fKYNi1b1EeJK
E/j3LhJUkw5mIwTk69ogD06OGeiH6R3CbWcJpel3sS5jRqwlqrpcjwpTfdblIwtnqbBEXveLKeXJ
hIwMkl4ESGUIA6V0QihTj0titJGP0LknG7tat5uXX4mqS5FQl+2MY/ToyNaszhkW6CafgADJ/vu/
E+UCty7s1s8rMh6/KRq8xjzGxdj7AnSpG2aBCrGY4wLpAXupPs4r+ny4qp4yDkYZNGNVxBgamzz0
IHMp/bAOILcmxVi5m86OzPMw12cI7mfRzgspi4UWujZkfEjyGyg8FB58J4mLEsWcOq0qrDVO0NZm
GNyxeJyEJfr4Qlm0AMpM6j4Pv7UbllZ9PnmacfgBi37N1hltPfs8NNhtyeDu+M4xcukzoogV7FNa
KykG8YsRbxTf9ZK+aTEEi9bTU59o3CeMuoCDwCnfPwNVYmNhXQiLayA9Xiuk7O5X7T2znp/lCo/y
5uOvg2IKsT29ucsYGRGHyfE7A4IlpERhI33xf1OIxxuvLxEGLASIqehiZTWbrtGybXeo2pTZAUCC
iUVs96DIlrPD4+nGrj+E/xj9xXiCn+xxo7u/nIZSOKmAdxqPdAxBCkCTDWonL8fUy+b+DdMf7VSd
Se9o66QEjg2PHsyy+3XHwo57AID6xdNI4JFXiulzVWw4Dc8EmXA8aFq6WLrk18A/PJXienZx2D+L
8hnFBg1zdEIxmiLJWpBRySF/aXQEc6Dq+DDZF3p/c/+wSvVwON7Bj5b5fXJYbWOUQWNPSHQwNWel
spEId3TESu3f0MIt5d2abbVUvjrTTE1BCR13uAJTwQeFkfDaLtgd6LpxWys1Y7YqE8dW58Cgtq38
X394a3A1UlkWUxTSj2kWBunuAMinKmQEx++iotTgAHQ3Pn7I+IQG0Sxlss4BHt7NHA24N3td2sG7
qjDBTBb3F5M0TAYnRuJwC+X/TdGyMs5D5hbHZYlf2eHjyAEhYkbpx0KQCidK3X3dKuj6vt9Tokig
XxL0NLoGOs0qtdyzW+l9PcSbt3qSWG6ChU2lw9B8PEvwSzex52NBwtW4hEoDUi0yYUtlKYS2me4Z
F0l32cMdUbEVBzkUfxrwCKQC8Ua4TJg+0o2Rgq7RgkHLYOQ7DfeOnGVMbcF03e0npdcMeeKSNL+w
PKMGzDQskBB8Czp9L/Zy3BnK6KWTZRrYCWzD+Gc8wOVj6iBQ6WBJxASHh48kkiWnAjDYoGBd51WM
QnTswyUjYurrH/UaFpp8yJKeAcyZMRhTYlIZe0xjGIjfqoGFZDuxsARfFljxFIDC/BsuSOdqd6Ou
6+nfJH30yH7RS3CEZ9HrT3ccBNYL6fGe72+wOzEmUbdBL6rU5mQKyN2up2cVS1eu0e8LXRrLug0C
t8zhh97CEz7TpsaHuwXe3XiFy37WIeriTmVsbDm17DOiGU/ZucaAboT3kgl6gfNQTjqAARdu6QPh
qt8r/33p9F4T4vL8kzyC89EKpU71lqx1EBeSWkIXxExQtAiv1AG+clo9PEmDSuwAPU6GAKwVm1Gv
iMAcjM9IBdsh9F3WaHNIfHd7PEbbXtDyElGGw9oE45Wc1pYrWEDBzXPXqYoSblHHw/JYsdG+m4g+
FBhIZq+iywptuJ3GQQ3mnGXXpaY/zoHimd9mAy/66REw7hJhI2GdwxtL+16JI6xPKW7MpsX8wJjf
9Kqrc1L0psqsQJur7yz3DtRIviPoRTXeA2YmOhuST8Nk4xOd7hzlcnPhnsKy4IDsOX4KUREpo0os
s9UG3gLO9SMWnQacilSg0s6wOgMYIqGQJncX1TFEBDWZ+2RiAVWMLM7dKl9mQbGs+9BBRVVWKBmw
Gvy6raaVXrrW8+ENNXDK+3A1j+Qu8ByDAt5OzZTVycSUFLXErQPcAR+4WFHj123PnT/uP98OwYeM
dtUGy+afmhjEqzxIcTo3uoXM4/MeyJnxKzoBwlC09dHQPKU/ZRepIMXMG6IVfR6B+mfHEMfxlHsj
bTFf/oaF20OndNYwQuSEKA9H33c1Rtsw41C7lLKsiLxPD3tbfWlDDT/WvDvqkqpJag3EyKlQdCLr
CNy0f1R9ewLtO6TQ61oT1bY95hUKtYaqZ92y3pI0/2tg0THuunYN4TFmcEpy7GRc96Bc9DRDkaFt
qpSpUJZXUJOZJHzHuQhXl38x0bnXRIJkyb31MO6fya8zomiYI4egDYQnragAoSMmHkxJL6w5eouR
9vlGtVHPEhP8q9CxNc/29frIMGoiiZVQvqNwzsiNEhhnDT00wcnNjYM3Y+DaPYBkw0yo7uOatyfg
TnJ6EeiiPHkTNX9MNfVL7nVi2E2loxTR0mFtQzmHTNxKe/X8ibqBHk8Oe4H+nXit1KfYaKpHoL39
1Tmzn0JZRX//QeTuhcBsbvFrmtx6ls7XjFf8LCjbIpf7DeEYTd2iGM/dyJEWb/HxB8NpOzhO2ROW
0sliFSkVh9LWt5QZ71Qw/6NBntYMdBf4CgdOax0VJqnUJxKqPY10y8bzZDQbdLI9T2T2/gB6wYyI
rt1JLFQFwjVlGMqLs5hY2b3nG23IZzBDV6EyrlYY+EiZEMh4v5C9PyrsDvqdfHSdfLxUbfFDsMqt
Oy2OSF/W0HJgRX+eM6s+MnU2k4VR9761zGOV1jH69z3rTB6+3LDaC3k7TZ/mRucGgNoyx4SCUZvD
tac3heGgjfArKf//loybYPLR8ZMVjJSHUsjl8pOz6jfPB+N3YUd9aJmdAft5mhD7lpDypyj1Bjc8
qON8p//kZ9Wwd8vvlvW6MQTJHrm6QbRLvwQtzR1jM09BLMz8lsA+Smjew5Zcab3jGJrL37tYNvxC
id7XrGq9d00kUkwDccxgkU+CEBS/lVTW5atwHxTNPugn8nR0c0Uk54ImTSdBwiDz1UUVjYI/Ep4s
18ib0UI5kN4jZvfmi6yYZQSP/SXy3/6X7zHHxMR5l3jGIYkjQVSD1UGob+a8nX1MfzvC5JxJwUzC
Gn0ze6z2mE7fQuLBqAp1Jy9TMczbLGE+0ZggR+i3bI/VfEBvF1xf5cE/AveYef5ZjAraMCOBchAm
PAPWhhiATUSKPv1bv29fHF4NB5ZlawZ4KpJzVnCLbMy01DSmWeDvrhHbk5opCsaJBMXqI03qBuko
hU0BKX6Bo0Yk5vP3ENyc0CzxhDdO8sc8nSky1IddywYECYZuIL5pEL3Wuf4S1N+JVlBgBeaA17oI
mQpDYcx0twvo+5Yb+ZwuNLG9WRDd+Mns74f33t7SiowkhL/8HZ2QWcwg08NeTz+F3cLMjPUl8POK
LDhetF4M39HLNR8qAMAu7JUBSTH7HWBtdAuEX2e3BsIjiXfBy3bpof1y34lMU1WSIrQCbdB4s0TG
CrvNzRegWzlMKrA4Z5t9tjTAj73/gCE6c19Jny5hBL1LO1iPcUSKn1d7YIPEndfzpnZbaiyybEEl
Mnva4nFXVqzT8pQaGvJb4dsPcAq3JFJsp6wtZEIxeysYcZCeSN43seHycKx/C+LGr3sYdddxkp4N
b5N5FpD53KlTfKuakM7nWQAbvY4Hza7FAYf+ytd+sLgacsQBdr43azWwNdQZOAPD902EEEiqIup7
VxNnigMbbIpS5h6h3v5dta4qRqeA0WcCXRzDzRHQ+rHv2/bW5wC0uDW/RZXoyZlTM/rIXe4zYBrK
fx13ko0cGiCf7siYBAgma3L8M4DBn7bSf0jTkL7S9CtT6Im3yZ8OZlWoH7vhvWix1y8XuYv9+c5P
cOb1X95TF2KcYIJb8Ubds5KkOiKfa4aXA2dJJzBsPC/8GGJu/NxYwSMlwpPf0/XNT/IdqBx1WMxt
skaWWUxKPtetjMBUhPFCLvfz0+DE53lpoIcedtwP7RiiVo5UAzdM+FmyQColSdNWh3T47csJJ6AR
Id/nI1SLAf4W7RNzYiJrEcXyRFe1Fh6e5h7i7rwkrS7FP/CW8/6/eqPVsjnTKYQkMUc8fv7qodCz
PTCZmfhD70RpiFu6R6PJjTJ8g4TIPuyQJ8t2peFCv9FY/JNCZbu3bKgNlEHA94c7J7219LLkIyrb
fmROToggPExjLaCnA1YwdZbUzKvC/rn/1pzL//8fE1987e2EhXFLkhO+fohR0fTACB9plBEAW+h6
J3gplzkS2iF0nryyTPYD51odizGmqnhn2oMl8vpOgO1eN+eYj+xokrofo5ie5pumKLwoWEIUS6n/
taTP4jC3duQwJcatX6XSjgAQheZhS+VoS+JZqjYEbAHQRn3ISk2XIe7sZxomtFZRjIyroRh5EmdQ
Nae3pI2filNFnJ5P5mDc6xEIev1qPqubXzou6QTLRhyG+MmQuQMRoEOf6wgWzabQaMqFa1+vMZUa
mOKc+fxDWGaZPybyf/c6QTAqrHH9MVE3ThUbZmpBiZnYQefbkISKqmPjWGigsuWqpM6O3jcWkWHh
w0RcuixQxI4rrwl5Bu0KYrGrU1C0bxlQJ5lX30UrC7cZL8xICEmaEXV5ZBXTKknZwQcQ32274aQ1
KQ/2IsDByGgZLdq5fuhEAmxghshPj6a0B5fYtFmN6WeCn01rmwP/p7oppcGKbQAaIcKthOE6r2rf
EIrua2LghhMZclluLvWNM//qOQROG+Ix9Cn1F2kbONgX/YLP8uwXv5cMpTkjr0ZcDejmuheTEFjW
s+/KtsheqJpGI9M1pi4PAqxMSoPfND8brw6PBfIQZVhIF2adHGRkkP6/x6QbYn6EX3+GMp7V0IwD
htxi2evVFdIhlLJZuIrgb6P3JUcve04pOvW+euK/vCGj9Wj3ebMcD/LvkWU7M0AB1GzEHSf40SQm
3fjQR4CaYDtXLsBMJz7mqX+gF0M+MV5xCsrJm0JoexuOL9fmAbXRz35kHxayr3gfPd3iYRRUTDbB
PnwymHKC32FgCKplLpEiBQ7vYRDoqKoF/mfV1DuiydrdN7syOgnsIQC9Ha66FkGGgfyV4YfLPjY1
5akFs8fr1B2q2Mc9QNYHKJOYGRtkH28zuKaA7yljBtA+5DeYorH+ToGxwRPszhwGp7geYszilKJC
WqHHuHnbi3fBHOKUJDkEBSCDuwj+9lRaSKMKIot2NEqoBG7Wkwx7MtEM6N1/DkR8rLOquhCi3qQL
xGIElLxH0kaymllLA5JNl+e0vT5mr0L3moxJeF9EFaqGP19nh8veSdH0MuMRHcMUj3KgrtaWp2LY
Ifa4ViZmi36OX9QGc5UOuPIqQ/pHVo2l7x8jBP4s2tjdWM0kyUtBrJEGwwD6nti8bpxIbsLt/xSd
RvEXJbhQxUTJmY1fF4IP2Wdza9GkjJsFXEKEjgPhN4YfIlcREd4NeVlGuMAfX9qzxtSiUu0kTLfy
XbPZProDaikooPfXWjuMiUqYO5qB2qacxeJ5n5U3dt+r7VI5zoXwBZXhVOccsiy2Hsedn1pYi7iz
Tq6yGW8vAJjSjPZfve7TlhOMLESNXfckcf6Bh2k8c9981DBckA16rN0kWAzsgA9A0BmMBuJ0WtfR
8Is976jSrw/pzmPSKHJqPKxXsRKdvljU63Bihlzewon6npMJ8YjfDgkwDJDeqh2OzlxDb/NvkhKp
xuFizoTFhqGULp5OBPG4vAnPLjESM/wihwwwXRhqcbcFjVzQSth5PUDzrP/vsYceH6UYiBLm89Gk
WKyb8VzYf32HPKU5PPCrRQUscGcbOnH1iY183Cv27pjYOBfREeRDh9LxvkKlMW31UhsTG4f38U83
C8WBVQkf1Mx88nn72DbGsEGO8yfTpk4B/hCeOYylfYAW8MLdSsdK4CAqi8Ng5ptLepGHW2VPTqDD
AWCe9jq2VjBKihEJLQQyNHEkQRevzgzfPVuQ/TKDjs4T/N1QZWLOc6X7wG/k9MgAbi40BhtXaV3E
5hOu0fkJDkEWo/qkKZmtuHr4mxgd+Vqx0xsDBqI6YKOAFrvL9joxeYBPZElocyF9qlvo7AwQ6hA2
w4OIQT9QtlBMHuS7EtXg5miqdsPDnqH7Zngjq9tFCZDEVCVt585kzuU9OD5m+5/AL8RnETNt0MoR
M3V3SPQwV5uPzi4N9wpeLbviscVgIvURljjL/rC3bDkv3QbvijazUkGllXmqhpV38gYGomOhggCJ
fn+wQTsvMAxNP0K3ixWJE8/VaKri1wXPDGnM9XrI60OYhk/rGVUIeDARzZI1ZOqmf9pJb2c532P6
+Qf/iG5KrbTYj1xaJbtV2qGcQSLsq6roZKEHudPWmIcIT0gtUk4eYykzk5jNSciwkk1YwTqvX8sX
bpdgB4yymnnF64wJJVWnwsOJXo+fYAFQMlE1p4JcK4H7MDXpmOp/EhTSZCJeliOX3mgqQHsc4MRY
W0ev/VrMzf+ExjH857kdHfm1D5DG0VckIXfmazj2+DjDNtt2VqZOMHCt6FbIzqBit7BunlZyjw5p
tYoi0Lpkc30McFylCBJ27MI/wk08aom8fiE2uredkY1At5lpInjm7tQxAZkmQRfAJ0bGfOUugN1A
AwS0p2sDGp77fwV+fzsdHqw0gbV4/1oi6KzOx7bfJl8U3mo4piwH9H7PZjmXd9zficquV9JhywuP
tGrVekFojuYpuKKwVMzMgccRVtY6ntbCndFudPBrsOrqAMBvLe9/sgo/SmvNZd5hetzdwRXHz9by
FpkfKhajGTahJbcCLCxIB6zjvd6Z+3NFNHY+gbwmz1p+6yzRekPEc9TdxhNPzJNvpicA4ixb/k8S
Xwzx7mcYkaFFbRtwf6jKn830Ckoapqg+grt9Y816vdHBBlwpAtDXZr0mNckfJOH4JUCIyKgS2Y20
+pGNE7rXNjCimsSdW9EySEnBvDtAJOm5Kj4E
`protect end_protected

