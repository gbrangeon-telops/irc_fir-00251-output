

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rMj+x3ocDbJ+0HvlMPtFLLYN4V3iOWmu0i3VYcvwPU8r9dUqilqv5BoOperD1z/j12cu4ait0bNC
TvgieQY6qg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LiFkBwHJvbvIRsrs7TuS9x+hbpgzWqPRKAN+86jD7W/DWOy2HiTI+Pr3kejl0F7PQ/wd2Tf3u0hB
l5PFI7Uciy5uXiQA7fDmYLdPcNoMNQWm9hohp6Q8wB4H3kSwMFgjlrwYcv97jBF9K/DD+f6kjMEJ
pjxxREwM6oJfyPhyhBI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mlNr/JQ7BAznEw9Lq2hOb9T0FUxDG5TxOJH6VJoPGS12EjdrVMK5Jwy/CrH7dSOtWY2eUHhpsxFO
HZJnPHkoY6pnOp56kFqNAyiHJP+z5BexlWOYCHMzTTDXl5ecpknkEs/jFqX2DjV6R1MuxPdeXOjM
JpDfpA+rd8xFCgAvhOcvKEKjw2lJmNukB/NqmGdLZU9Yd/iDC6mJcVuTrR2gzFDMoFjQUitH7TCG
r1krtYbVQjkm691WyHmxufh/qSc3KdzrpZqycBevqxjmEqCq0nMXCiMyQRHMFNk9XLymhnx09LIk
8Ck9EeU7sTUKIMhZ7oB9NRbr0Jmue7w3V7zoXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jcrZIuGwyVPSe4eEqA3CjxEN8wKBf64m71qLvmqrllZ8mLFeyFjj3f796U4fol5LeUOSCUITklpk
5B0LZiT34IugfACCFG6eSa/KnYkpqdaiyFEJag2zBthAbQTJIoKzv4hrVDSwoJffRhWS6ZAZmMOH
9HJ1Z4KODhrBj2PMMOQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
He/hsXsp9htM4v1ezeHFxTi8NbCInK4GRCTZh00v46syUmSwf+mXhIjhLm4sHKCSUqmWt1TLUp0m
CWcpoGxiawBF6wEpl5GgUNyVTq+T/CrlV9Oykyiw8ESh1/7hqCFXSES7D6yS14KOyEm1cr2UmC+u
X/NTzDDvOd9e5R6zaiks/z3Qdqxiq6f6jnMuQiSiMBsAMCHxpq5kEezVTATURKXvDebBjGkSTomU
Wve9JRKQPSiMHuUURnaiqzi8t62PeJzIwk64jI0DQYpuyHeGDNIZt8qQokGYPimAYp9IilmsSuGG
FM6CnM5XioVenoNWDUkk1F8M0K5I/5eHgYEnkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30400)
`protect data_block
WJ+jOOUadL3kfZgSoSj0ZAguYc7aTTzV0sKkUcQiB9+4FZGwTUmt48RrBE6RCQrkPvlW/hBLu9Ve
tiBMnRj2OWYpln3SCgZfWEVNzXow25ZGdfft32iJa+oW0NeiOpySiPMWFMsM2REIJ8U/j/hznv5H
pTnGlMvBpZ6ftchGwrTJo5cEa5DDt3MjanrFqC5iQK0Nbr1pxK5Q2Zkgbs3bS5A8Wxrhn0igoPU3
2o+c1iT4JpKlsI7n0AR9ooDu10EFRwN8LmJ5bcmWRVeH6/+NCQN2ZTxr//qmu5vprCHRNEXDZhq9
+wrty/R9mFInDSMUTKCBJrdmeVwNVvSaw/lO8aZuscatoZ+6x8NPSnbLx3tp+NBjOqJe3wGLLt9x
kec+fvC/PyDis6gn2NZHLkKiZyNRSgX3oixPuhiUUlbsFf3d0w7FWZvYLNYlKIvXHAiNUnem8lw1
8LHDeCeLTAX+oqs1Q/Q1YomnCNfR+7sTCwZ5B3JBqI6B/sqEqPScAUDjDvnFD8P3XLSmKp/ZWXux
Gcr4uBnKeb8tfoFVZCjViGQQQifn2cWKY4BLATdPheqqZtUe5OpeezbQOcoHOSZixjha06fpgfIx
Vqu6hjo4Rq93uf9HWXgdaoMk0T/RQQtwxIEviT88/Zjo08K2R5eFLVa5OLMPavXC6tckqsZf94In
tYd5SE1QhikP+f21ZYtpQ8W/Jvw1PtsLGv0zwTJMPH/GRQMFQFWVtEYSQzysBnXCUqFnjmsFPdq6
XXQEuT9OjLJtkHRZs586/XWluwRZQ0pq23Bfh/MQby0xXU4xaYhvO2424rLd1n/MaCDlePbD9Nc+
GTgIGCLmkNdLf2Ir6EATAoo9f3D1kFibfOndw71FSDCqC7ApOUoA+lIE/TC5rNLxxrQ75PpHd620
J6G2Iva3zn5XoS2vQfotPuRpNGASZGzgZvR+oFdyzC8OsvQHqz6N8nNmLII1qPqTxyGprn2FYED9
NMGhMojHZDDSc9hJSmxNeoZ/oyyxUhOtmlwqNqQ4zB6/BD76Ks1co9SmRzlzqip7W40JvmAqOKWY
kILRBKzeg6GYjjhK1ID7WoW646ChCDGqmjdx41oYljf7ZuPSNZXVbBSkzH5PQghm2gvT47I2Lve9
QVI3m0/WNwmwNnSC6HCfSQFfHVZKAlTQ+vjmA5PH6F8ITvHkIYfBlPIHu1qiG/Lvnzp8RyP7aQqD
Rn8Vr3xOomY72a3uTnm++sRO5z+D2GpU7jOGAIlD3+lLORCnagk5bxT7Gy/KAsw+7BGhq3EG2BeT
DTo+Dsl8UEmQeVg3QA49AWpVuSaJb6ADW0DtR4R2t4ET/UvBitUNqQK1GQktTxbDJFiBjDeEpzcf
G2nIK2dBknXFl+EQPRnWxxUugXwQxQxOD8LYKbhBzew5YoNVfmW/fMdW8vR8WYITIkk78XKbvxN/
NltVLC7kV9jyT8RrSP4leZfZayHSxjg1V8H2Brz6+VD2pS98agO3KWkPH7ZzsTN8rBgMsoAM1lDy
rQe9za8t6j2ezFKqGCzgb1k6FdBU/qqVKpgfrvzyPjYnw9nMTsP+QsBAGrHVeaMYVsmP6k/i1U3c
t5xifgkbWWF4+RWpJcs6yJh2a7KPe2lgivkImVh50PiVYxSDYlVQeharHYjF/H9q3e+fUQvC+yBo
ByhS8rmDoT1bR7rCTBGGN7OusziMV01rNaLj8eitRYkqNgeVRvJ8lsXUd0S73lDslNgI3vFPu62B
D2iTwZeQ/5FBvEAxTCv1RWokSZYoIYl1sbWwAgyi1aUPuGLcLIr5ox4qUMxin2/4UkaGRjgWRJXt
3IlLsHFSBYWV+q417e4xgKx+eLaQQKlrY9EFBNdGAR7tcHej7HSuXVgizK9vLlGzgBH0b1jMZu+N
ZOGgKJCYEW0qRAy+IMOZ+W9pd6xbgrduPO9htdjXz/xggW+EqXxDiiR6wcucYRqauhfnvmSZRjMh
ASFsng27REtUkpzxf5GL6jiPt9ZCpCVVTygZGNHn468ksuGpPQ7vaJ+ohViazbFzWDAhkgwgJSgI
AzZyu/uuugPSsGoJA/QcoVB7t4Bo4iDFqxduLhq/bqfFcrFd2Ncn0VS+WlRj0YLk4g+8z1pqEos6
SfLG6rombLdJqaUNzJ+an2VKJ3QSpOXaX8z+yPNYilwGDO4IsHd+Z8W61FefyDZ+Um1zXTnZDE+v
yWW9Ygcy1lMLBvYZgJY4C5VoL1944b48Tc7EmGCi3lIcy4UsuyQ2YSe5WBb1CIeATxDziV++csYt
/mvT1aS6QN1jX2Pf5x7yeinm7RGPQXRHleifpsgGZy9DqXUdVzRPauZUNNFiuNeSZsTpxNLeRpal
QfBLfidqmVItjZr2PvkXIXWqtHPUF16F+nvOQzNWJwsQJWFqnk4gasdckqxEbFxkMxmUpxnAWosC
hATaT5O0s6oAROVUgdjcG0GU7ijecmVXqdDexuuO0yq2MvT+8NwXyGAaids7cm4kuwOqsjePEQQ0
TNoK8q9yP2sEj67BRPyJSqM4Eq5da6qOmvLUBzx18kYofnk6jWdkfsZIhwnRenBGmNqNvw2xdeDE
kyipNBfMbdJLAQBzHrAFGqGAQV0pQyQI/t5QHqL2KTe/q3Zv+fYIqj4JfFgxUh4tVlNII2i5YsjG
V0lJpe07SWkjvjZqH0AYnX2IAcgt/mPeuY74DqyV8bii8JuJhXIZnbzZasG2nUGKcEoN+b0NWIK3
7Kn8yjrz4j0xCeP6+XNveIXG8M4FDgXn28EyMtASN7KZib0YwbZ6pQMpz8zScZglB0FEz93sfpDs
FO/Ks6nNtCoeNdjDMbJNqyId5yuIb8/B1RFbtun/apB6ptXqS8GcxOMmPPEwj+pfwR3xY8B1i72a
Sx4S0XM4hr50abC4aTsq4hDkZPqRDoqRK/WZC25X9+OYmJ8fwElxTlPVsQPr43mjrrXHPV/LwUjC
zeG6g54IUC7uRCh6VqUMStVhR500O+5qDPxf+qmqhsD1/0Elfg9eoKmTunCX950PluFBNNTLesfP
yjbricRvHLU9zv+XlcB53wl4qCYZ/cuEXPCae1dV3whq3O/iwEmaztHex8DgXArE2WqtrREWdOCK
ohYJj+BJgQHZyAbNZ2aFQN6xGVCoC4+iWe2LiUAt88MvWxw+JDuEu9ZUH2cwt4ltHI6WCKPA7w4o
3AzV4halX35dPQYZZ+6e5vtpVjC6nU7HmVw8A5a871XTs8v6VAyzx6uT5xHSkK1V9jIDd8R5G2BY
X/WCkFqPC0irbHmQ6N+sNaEyPxAdzJPd1Pg55bsEJTJ1xJjCN5tSnwKI7Xo0nC1g+BiGeu7HAoxb
texbFjmsDbB+uwO0fVDCu5Vx2Gb3pVQrHDbLMQEUDTd9Y2JEPp3GYKfez+595pxKxpjrA4qprZ5O
oK9++QOYeNZYnWjmfV8f1m8zs8I5DL55vy+VPEIwrwc4i0pUKCIRNDT+o0IYu5DhdQQc/QoAiO13
AbtM1y2B1CnOWHn/SqLL7hkUsLKLa4wuxPMvCH0ccdsPe/HZCaUxb9LyeYCENUz1tPOY9fWC41jM
BSYeZMVX7moYnOFziSUwvK8Ck8cpFjD3itoozTV5TtLsns4m9L/EUVA/GnTVK6Uht+4nuU3o7Vis
s7Q4ECeBmLYpjAk7mlTXNBanugaIJtiiwnUQm/RCT1K8JQoiiyF3CgHURHVC4aWZOpJdGah8R9pg
gPlSwJrAod9znfBFaxo9DeBdZW+qGO/hDRs11KDM1Ow/Jhp7/QWnF0/0s5v/d9Ac/oABjX3uLk8e
lEakHvadoEMHN2YCaFdpDaKqYqRR05aoThxm91qH92FeyyKRTy8JrZMSElnFgTd594ko5uudj1DV
iS/DuD0SvfKXRpvKjcMiFkuWQONTrRJtN2wg9FL9m7oyCPAS4pzIzDvsNdaiQKVny15pSIFO2ltH
gkVSelPZuOKChX5aOPHTbVQHRwHiOAxyn5ZKTEIRx9//ILmLvI8BEXjewHbYhUsAtNCintxHTYwz
RIiVklVS8gON/1yCwAGih5a0rukSHC9AmqTvCyPKqwYgS0QpvjkE+BZgeSQLxOMQHbg9n+uIu6Xl
44LkN+Hqw/cXvdUJCWzzQSh0k93Aw+vV5xHHTzrFpsETrzFphsIWd+EDsNixz0yQbi/q6ICYBHXm
y5SUgGldpn59hsQSmKOsceRqxO42e7t1AElTDthAk21toyzirIc6tEP/VU0/+UqHYE/AUH7+Fjhn
j1Wp1NjAtTTifrJYRzSLH8nV2Pp9Cm9uen0/Ru75Bbo2c4ibTCMtBSB9PNn8/xnV6+jE2PDXAEsv
GC23LdGOpT/Ev4aBuUm3DVf6MebOi4ZWjZOxU+YUZtFLYc4FWWVtnX83v77BoczTvZjiuV1JibOF
YP5OOMxhjITSubuVDBQSP4dqKXRk4+nYap4nbrPHTGeFI3JdRCGfol806Hm3DyiPRjnxv1E/rgCH
J+bD12YMilmcwAYY+r6fULAh5E8G/uwmy/wbsxMHPr2D4KxE88FwVi24Qh4sgGTvz97Swa3jSFmX
or6tvoQkRwTKtxz6b83x5YH6vpjo/yMXgySZjKykDkxwCaZHrscfjVjx32yFA0h3npFDREecdMLG
l9P9WS3kXsrRRngiuWYWswwnRYq+nO4LDsXK/LqB/pwcrea5ew/X402+4QTfIJcjkztPrH2fwmLa
pYO5PbbJSkDEax4g9mnV0ZPBh/7st1k3CB4GaRdVNpkGoQH3k0flJM71HD3Qw6niTpZndkn+5ckV
VXWcB3HZ1JwXNGIk23i95sn8/y1RN8enXLBQ6cp4Ijh1XwZ/bMkkgIMobejsE8/HP3PkOW9eP7xU
4xd/QL0TkcKH3wcbxz2vzdQq6XR8hX6Zogg6OA0fxzdO0xHDkcfm915hrtRgtwDWGT3WddRuONU4
RnCj3Du1yxSMjpvNTVhDGBm66yJu/dkNMijenbsNsjsfapKk/1AtJa97fdv4TuJVHB4XvhtQPV1b
j0YW46vWrng49rk5zMmCbMSnB0CyiyPQay5nFmDtySjn1s9IAbNFzNGM0Q5rJ1INc3aPTZfabhGn
BQuhvukgDHT2OTq5+RANXFMi12ViPTxrY0BpNmg3+yI11SCVQId9+wYkU0gi1ZO9s3CdnEzS4fLW
uJOFCUhrzqkvveysGczJkBbe6IbsBxwD0tscBKpJy6oNKoMoZ8ImLyi2H7b+D6xLcK9lf9tFl7XS
Xv92/96I72HZALYloCm94sXernWHUssOY4atK3ividMP4H3rnkqebHBdgt2z3hQycV1+rPb0/nYC
Si1UoIYXb68vVnh56IlJeoiqc7n+hSjJASU+Ocga3Q9FPJH2hD047IJ2mf+6Tl/g/sV1EtxtFgjb
1YxShJYrsNf3cTkbIQ17EAsRa96HOpZjB3DtZ6vPaToLCHxeWyDLxFBvEHRKyp+yef8pbLhoEWej
IHzIkFbj09vN/dFTOFKhLH0nXqmmLZ0l4ERw0AsGtlPJ5yZkBSx3IKQLjrXSXAne6dRxNUMTpEiw
kAyQtsq/SEJXdNJ6C7+uSZhIaBLp2fkYZxk/sbdsmCLPRFIGKR/gr/EKIbbxvGcUuoQwR+gorBar
hjMi/aAfwGfSASJF1qcybVV+oY+1xY42QzqavUNxAEsA0+/vFABMjHTD3qv1JwLPEBYfEgYQcrft
K4C0KGKgG3MGDnAyRpD/DcY7ntJ5cn5lBr6IzIdNiauiuw2TMIiSWyl+yeS3XuzwgdWgQYlT3WZ8
/vmTdrRjtheSwiBD4n9633pWuPfSPF4BXv1qM6W62qM3Uk66U92G26DGIWzcVl35M4I1o1CEmio3
j6lcYAO+xxj8j8A2CfLmU/vMCgPP5evVqLYYtMWKaKE5ukk2a+Qx1mkISWFoCpaqeoJdOSBcmdbF
fSoi8QGAXpSVyDWkp1KkmVvgDpZHCCNc6lHzxBrXHZVp/mFsNn6ugzV40Ba7QM+k5xX5otIG2ihF
IChFsoBzghCSEeC4h8V6SGgqh+2smTFehkKfRouj1Yb+qwwBjw1dtpWXPo9rQvoz7Bysq1a/KoTH
e3w9swVu9vNKA5oaewnyQXL7FKJ5DZ6GiQduuoVMw5wrqWwg3iSrX/iRvptxLGugnoQ2fCq0ANUX
2mHUfZeEK+eAfDn9UAeqvLEjFPcetmRWEEoq+K57IdaYJe+x/f1Q7IdfSUuYN6pyw4v3V+nRYDg3
sOZWZzfjqzMVbl9+znEecLt88GzJnWuuhZuZQ2CbYlfp3DMaA28qxP6NdSd/SeFwlzyAnmbjuV/C
tZYew0/Q5gu1mEzIwniR42iWx3gyi1fknnQ1FL6pgaxx1TjtQgzg5upOTHm6k+TRMjf6NA2GlF89
a2Fme0EcyZ8KZ1on04LDbsWoz5J73GT2ZfzIos/sNf9qZtNo+q1bikwvKrEpatLAM4/hDe2dGfOh
mQg5gPIHLPT7D/H7AGLTPaoMTs9qeHr7mU2zrjDW15IEV5911zNWpovX1ImlvH7Rz+WEEZC71Imk
S6L5/lQF8YQyFCuta8APW+oFvdMno+lI68Bmes2EXSy2RuI5OwCsnftyIMmO9TxYcvcUJk+c0no4
DmszlT1buBZWpmvwyAI9PXFT/c0Jc1gxPXHxmnS06pPKcwA7VognF7EY6FsqW+1WqGRbzyk6LzOa
UkVH2fIeBWez750l7Y2hkHUThV80KUNBQPeIRM2KOHddOYHYuIBYI9iA8xXsOwou9S9+PXW276MO
8KweJlvY5fOIPH+7mdlSq84Whog6tzSeAMJ/I9zbf35lVi5vcXmPsQM5W1K0ulRtXHJbvylghTAk
mBL8dJaUoJih5tiBy9OcYZqv4yI09S/N0TzHePEcBpoLNtMeFFRMt5/pUCrlrzinQ4GxpGf8ptW+
iBt1/B4ACRT2dg2Y35qLJGZoPjvzoiAqJimJu1nz6g7iRCVTF8QE4iuofQ9YEMwTRn+grn2hJQ91
/1HnW9YOO72QeiX5RDL+NFOQEUo8AOwkaANwBPQkuNyRiSbSI+b+Qyt/h////3OBHgAE9xH5cRHR
BDhT29IkHVLwe6k5POAX5aP7Fr3tjfWvMjWV+In932SQ/L9DLpq+GoACMCw4+vWpYi2CRPGmPFZq
ZtVEHn2JwiHYunY8wHrA6/zpVJCou2nWXZr7MiLlpD7/eFFDrirObLCfJsZPzxy/+YowgWmmrDsY
22lajexkD0fOLn6mhyEX7cfkdHMIKxaJ+ySM/yefMwxo//fNcCwCSqs5qTR/aTERKpeXywksuosW
L574sWA64cVYU+1WemHjQ59vhhy8wlOg4IyD2/Rpl+AiO1AhbAXcph+zgFOJTl6zzDMqr76Xsodx
Sr5DOZzse2fl/bXiBfP435aNmA6p+yXWOWxZ0gnVcNwoBq0d0gNAkF7WiHbRbdPJkMDi0cKu2tfi
UyeyAIsRNquF2n0ZauiZtM8N9AOYo6zohF6fFcSOdHWYt4M912rLgKgnvu7kti9U5M3L7CyVrF4/
NNo133GU7v0M3eE8TXjTqQb97CVHUXg0sFAX204CpaniJPRNLNG9XiSgN62mReVnv8EHPYvaGhWx
EmNZYmrMdu9DIMCfKsS0An/pgA507hn7ciPXyRYO0teUEc4IXtfNh4ej/vyjtHupKR6TGNmuxaX2
IMGZWVOg64bInt5MGljyXn+H0sxNkCcrnN2QqqzluBHIALhVGuefudNCT3puhli30H+KDi8Oggsx
VSKi6XzKjl8lUkI82FjDpmQaNcUhpMBJ8Y23rQh8vr96bYtAnYAOgtqh0+NXd9S8ZN9Dbbty5zbE
oOE9A90Kzw3HesBURa8uhwaUjRnNPKfJ+9inLfsj7TGpMcdY5V7UTk6/DLbvBP/NCi9UQUsceiRE
4T4GaKMj2tVwOeu9vEEeev7dQv60G3UjSHwcumBxlrEAfU7r3xRJQGedfeZitbh8c6zG4D1uLZn+
qG/FgpcJFGgtWgiRtEefWhtaappmUnnC6JMPOM+JvRk1v/VXULLiEuH/+uWHLuar5/36pb4N8rgg
5PR2mn8aKO8micMs3PIx9i/eknPud68jeCnNdnPqE6HNfwQA8zVbUReQPQyqMCbUXCpWgKjYPKbs
peQjy/EiIiQPd4LUGFo7cVDLk+KZjMDnbYaZSJ9AD3vgmErJbeEaJ3sxMb+B4lTnGi67dRnNvJqU
RfbQUkcfVtdFQBAnUf3RsTOwI/RUZ8t/aeI2Z1cM7KNnNZq5xhsTJqZYrHDTM84J6AovLb1pelMK
0HALF+bpHhkMnxoPbBFY3SeRaMQtHs10IJtbV3Rm/MkkzlQjA+Qf+S3Jqas4KquuRTC1Xufe6jcu
OcKygox5JcUi9Dq0j0Tp11YXYw/OCS5pu9YWk75DIjeHcSBVkkFW0DJzGUkCRpfS45yo5w6VnG0A
aYQeG1lQn3UsJMXMtIJj4ZyzZQzvCtOhXZFt7WmSE9j81PV0f4reO5cAVZF40D8Gi0JAbm0RlurK
zhePDYMMSiD5GqfvTr65/C9iWjrtBBkKysAhHxF4IPCtjoTV/tXldZA+ZhaxTNdezDd8E2mmEbe8
KH0ZBi9kucIPpl3Zi8SdX633zh6hXfjM+8YTF3Kh+n99eJlWk1Ikxg5G+58ClbkK5N078TAlRIhr
Pzf7+FY+cK8nFdOuTtEc0yuW8xHAanyFBzpaO3Bbiaf+gYa4W/UmY31lkmwq3GEJ+wqRy7i0/aZc
BHSsuw+O2lnMOt8XgjIgR9gLki4cAjOc1ijA6X3+5/iuiU96KxzsRSg0TyHx9V/YUxWuxtwyqUR6
Hp9G/e7IxKeG9amvTcdi+0LPm9KMuaArtwMhA7Q1eCzFdnAghiqr3gWCGEYGYPh+NVmH32hRt+W5
/FYHkcC7HPDaeKWLPWPb9HIs6CKHYSGauZA18PCMUuXcwQQPnrx9fNZUl5l9ivbRgACrG06HGes/
aayeQjRpzZbdoafOkMcTay8oc76BmV/tOyAbdTF04qVje/1+ip5LyeWlyinzoENCVMYutERq/rvP
tBn/PxJcsEW4j5TLcDhdL1iJnTHHMfltaJAQRuMJowFsTlXUsfXuq2W6ErwTnV3/n1b3SmEaQAm8
ye8R4Xk09Epkw4jQZqaOCUpA9EueOhX+Y4l4N/DkQQ4GtlD6B3cRr1/OkWCF/GJYTUnD0CAsqFmM
DWDc0POsHCke4o+AqpIZrxYUCTab7cvsP7adkepFqYtr9YfmMbFrDOORZ4ta+2PzdAvGkoTQ/Hoz
nM6girEMsaw4Lcq5wtc6tyDYOm4c8JNIAzYkXxXMe8zq/aXiriNU9WLRARSGHthLaEooS9j+b3zF
n/22VSq4Z06tWoLO1SbWd2M6naUR+GY0li3bTK5VBLMtB+RbT2g+v0Rje6DQ0lb6W7LGc7S/Xvy0
kKcWBdjoX9XB6pPKMT0K6GHOA7Mx0HxI79FnsSarKc+/1l8f7lfbjKJHeWseiXc40xk86wwH5ur8
F5k+Hxie3yyWyiQvTxuZ4ypO9EYebcd89ftPaIqMuTzu1J8GXS67GFLLrkG6hoPO1pBBKHTQN8CC
wrgoEaLqHqH17rPGpjb3ff9N0HEneSkp+luMWEWEt8r4nxPDjphU4dhWVMdO7aHHY8NyM8Bbt1K1
Y1LYBAwh2QPrbjB1EOrtlGXov6OBXzZ5fbmQhJ5gXNA7OTjrd5N/5cY30zICAQv8HKmgV9eByKE3
8ZFiMjHGA41Y1aMtKbRHEbo06wpx/dEDmBoF4w3HzhyMHXE/gURAGcTjxvkuV6AWWlFS2ShRCohp
/u6vYHAjlMbf6foq4498nsqG3TZ9dMocYvwW+WxV27Pg9wus47onvIIxpBAgYaviKTb3G/TG/O/b
GrbQ5WUGh72rpo/iV9pZ9n7LiIDtPAR797dnkAe0tZx2szv4KiPkXDbgPfzDnMPMBTOExSFIbXX+
WqWiUMSmV0U2VJP3ooiduITyuySx7+Xa3I0kzs0T+NGv7E14tbNvoAPaNPm1rxpQVNN3VwrrIpaa
v89kutTDkU7QCR5JIw7RXh8kwxnHrbDdmWYjbK//EbZemViyzWhBmhzR1utk6ScTdeiZF3Un5CaN
OiCz+T2UUz7XyR1jEvCprxlpjoL+ZfqxAguY64wBOKrcl9kZY9Pin9dRtgvkvx0P2G7XbpCL7tgC
pVX5jvzIslJveNnjEpoYhgF4KQjEWOrZ+Kiw0UJAPgbfClSkzcxesSg5rApIFChJy1fCn39JLig5
Tqvd716+3Q1q9gRnAeF2PN8+tVGKz2TB7yICfTC+OwOzlKj8lheDl3G9g4XFHq8WGDJ1joCGbHWg
ZjpW6xfbf/E1hLQ8Oj64XuUf1lVr5COu1RgrGhqw0L8I6u8Mq8mA3eK2Pyd3xV41HUACdgbmJ7XJ
cWnATTd7wohbKK58YaWjIVdC9MK6zGUUtsKQPTwQBxYJpC9fPdLJmewzo+mKV6eXv7jagAGDn9Ei
FMeYB/7iumI3xreFKCSycAbjddqBURxa8+R5zfKggG9kRTFet8sCaB99oAdFDoe8GEjxZ0cwuvX7
VwVjKLTvVzQe5OUERoE/As0KWCvpcZHHt1VCCBFF1Uc+VFSRBuprN5CW7OV6qLiWw5TVdZejyeUM
9v+Cf7gYkQ1Wv9+xOLLrB8G6OvnFVubAOvXP46J3VE5Op6EDDCYfidaatclb1/+KtdHliaBlZzUy
08ZgVCKaPLtZgBRoxi+q92uT8bWaotUaXDmdOvjbEmtGYfBWYE3m406GK/Ycj7FOA+KXLEb27Znw
OGbfcNTEohN7ClUvggjRrA/hCDCFzPgPTTFbCvaan67AbrDz/RCL43fth0uvJwrBjFPf/MqWw0bh
hWCLsDa5AttkpD3HeNHJr8cscYpg5C8sHBT43vPD3H08Li6CUkFRGPOCP9b4e42EB24tF4bJYh9T
PDFBlVo8+j6C72ijwqSthx0Pjn9qijQmAB1hvJ5j8rsmZTAZ4q+alsiig/mhrBIalKc6xtL8KDcv
jQ1w9JnYtYhC5P49hQHawdEvGrXXwH9a0pEwI25AdVYrl9ikOmKtNqFQqCpwbdp6KMgI0jo/WmPJ
zkqbdAoyCjA7AAMxVVkbjstzMqIIShxTc6+sbJJQtir5vvFlJj/Qo7l9xazAE5/Z9MdIzsNYiIEt
D2Y2X9LZYXQ8iQR0cBNHWWENll4PgsvKnWw+f3f0WvDEM3DIBb4cGTYE4GgQkgvYayYZMOeZXCGu
3qDEccz4sV3qHXPWB8hxWIdWbQVHE+Jf3stqYktKtCRlYww7U6ITIzt6seHTQik5xaiWa00v0KQz
S0howAWdCrGtsq68Itrp3nrKM6YHH7zppOmBXpmWPw5NFs0KyYJbu0Q0TrGMMbtwvTo5zpnZNw2V
YMG6x3p4csJ6nREWqqS8806QOwonf8LFFEt3b2bl/8lOWoXKF/419aiS8OM2fvG21yBuCF/dCoiC
bMjw2mqCn8CrYF2Ibz9dqP/kr8OxrY37sRL409c4Y00mTB6H6mEi+T2GnUOwr4QmcxWIiJ2JM/b6
NEIBmPXFfmhUu0X3ISlzNJnrMZoz2nC8hgh5CTYHmfjYLA8r6kfeYmHazjmFnAUMwcENUlYLwilZ
LCXi3Qyf60CDK5l/ED63sbnDl3UfNGPVRb+IQKpiWHIidXn9wEFbVawXooQloi1qOVnvKImHE+xf
xmrl1+Y+GiaxQPJcmS4TtMZh0oPlBjfHWzNry/mK92uxMAFY51QcWuhPC0VSF5nu3S287J99QWra
6E/cnbqrvciV4jyC5963/GT6A4n4OE3ulxyLEhX/9em806DqjrUBbI29MPhbubdQRI8E9qc0B0mD
ESKIG2NENkOA3QYf0oYC9pEvi/y+ye8Uxyot87nWakVXcR7Katixbo2alZzO1W6IZVCXbQgpieA6
np/OUN5sSQUavPmnZe0y/s6RongzVK/2Y3eeyKGtVD1MrCKkYJCTDcAXxOlQZO5GLNuv4ZqBCiOu
C6iOKh3gMd/ahLGf+hCV6D0kHMJ1QAUzJTeVL3eUr/mpXxpqmf0tb/nXH2PgjhIPDsFgFP2FF3aY
LNHR3vN2MDtiO1ScKCcwlmVFq1hVfhb3/Q2c1I4j5WktqjRm1pQ80Aaxfcqzl/ElfWCEDApkCB87
s8HAjWQl2gAX3wiwbv8hXl+aux7GzJE2NOu7RlPRfDO3DgWL9Uly0YIUQzk0Dj1cJeUvD+E7wYhv
Lq/3VldM2vA+BmXz0iWhv7nNtUtR27XtiZvVh+i1rs4UXfp45dXCOGdtYcn447OfVYmr7yafYXLA
cf+FOLL4Ru5jMkI6I75ritEgI9C2DxFJFpdiU+mB+oXP/RwxyIw0DC0YFViQIa0T45jaNuj8GUgV
NiZuKjlZm5UOhbJua2rlsGUj6lupDyURgv5scCitwOhLi/Ao93LLLOoR/Yyn/hsugFZrZ8UUvHYK
nYyC0BYGcILx3WTNgZ3YbM+Xg9EW/277d+h9qgzPZAjM12bf1YpRXZ4HqR+sMk2CWBRapV8R4iKe
RMb4U8za5LFurpgQpUI8m8f+JzDPOrfYEa47gcShFQ7WGaFW8t6LCPxmebFHuK7BtVgn+uyRq33I
ubifjoQyLyKX44p3OPbqpeJWXV0lSRNe0FL3ralaf+DAlWC4aAeYGrm5bMpUZ18BJag4JCtjNDUV
xITX/H9yR9TEAzJvhJfThzvqFBAe3XPAeXUDUw9YjV8gtlQRXdFa1Bhw41vAMo7Rs/O62GgRdEau
7zjCNnYN8ndRuLAQoXf04Y8wMHdCkiyXmk9Kljsu1Iwta571ouREqaRUvQwP5JybkDjpwl1IHsWj
afMc2HKytCyKDgjRgQH1eR2xwAaAj9IC8uJ7+McKwNO4SCu41OMkL+8o8GWovQi24BKvA78ZXU+/
KQAku2ZJiqrqmzoBnD27/g3JMy0S8JQ1pxiUUjI7oeXshOkU0UuwtdvdDXj5UAqkF5PASVE8ijEa
AQdi2oStwQ6R8nfBIL7vCDrijNhK6mHxLF4gvzsvoATMAHRNSbveY0peVXwfrkPYh607Vk6nuMj3
nUCt/iRHi4nyKVMNUHFyq2M++NHTTxZLMwMJVGOBd//vl8I/3u/9/lguLTM9zNtR0oo+tFX3tD0c
FxladD4xx20cOif1hSjoRik4l/HyNkao7jSWlI1Jb92i8BgY9uxDEDN6rV709eC21mfVQYM3q4nn
bGv8be0PRD2BwC/lXh0TZrG0rwCEMV/iCY4dvFwVSL1NcsH9U9OKIwfdPo+jJ9BGQ1WpbxZPfRwB
i80BvdwtGipqZg9GG5Y830gVgfQBTMo2/bTJ6Zntz+8K1+v2teaBUFWIsl8TYyRFEfJPC99IZyBw
mKjz69KSEcgdwad+xW3Qx23gzFQ9MqGFANi8cJeR9uJoBZtE818AJBz9QAOxQFTMzKZ6hlmw39ey
pzEf15PRkzF6yg59yXW2CLvh6MZytDWFGa7PltRfmhpKx1sNWRTl7F2t1n7lLg8iaSH8RWAWDml5
BmC6p63A11sBSPXUiRFL1W+z4NGX/mRTB+GWICKU01JNEXqbg3VX+5ghvjHQ7MuOkqbLPBQdKP2e
6wb/ACM0aF5gyb8JcRfMVvAxUpYm2sMRudZT/41tKH1R6lf3viJosEuiOj8dAs8+adVomK7MSyKU
NtOr38A2sJc9C7f/0xT8rheY1Gv+IuYaJGLvqgfbnQPbaCqifqs1GNeCXDeDGdGtT/q0rRz0D47i
uTzckZfQY/unacgDFPZwW2WRoWnpbtYJlGuuq+hCZtFmV/Cl2ZC0cDTYpAxIhMRST3zf+GnM0ANi
SNBCmgGmPu5pz06PmL7K3TjtZcNXNFzGqy+3in0ScWU8R4Hpk1Pdq/O7/6chdmWxgXOxfkVRcQTa
tVK5Wp/ixAxdQaNyFZFDF95VlKcLcAx1JR6lfRdsyXpJUbJPEItZDun8MFTVaxhmmoA9yC5R0pLz
YPW4uEnrZnMYbfHIhqUAbvMnLgPuG8uqYRNu0q+y6QRtAlUXAe80DT3uCjyV3960M/jomaTJ8++c
P1mIF88agpp/AlVjPQhRT4Lho/ope5pm6sEmtk83Lw5ioOuNlznA/XSRk+QkExcbnR44vziD12cE
YrtNI5DuzKZRHA7DWw0pDf1Z2GT6xXNogRRFP08HdDH/4AsDwkwQzAitbiraz6SMEj2gsBxjBP/U
RtxNnXqPd4Y2KSqJm2gh6nxhL/C9YZQwaRDGzsmdmlXDLSUX9mS8T0miWiLEWwbTrKYm5nNq0rEV
y80VlqZNMyjRdwqTVrcDxJE+MT32uK9Yk71MMe1/W9y1QdEEfuaI8yKpnn3IR1/tqP17c+yC2f59
UyFlHnadqZLg7FQ7bpZcYwi3S6kLluLLuTrcB1kB6m7UhG08UujG6J8XQO+xlQq2thzCqIqaQx46
HWfKnOI9U7JzvtnCpX1DracXtbNcy5IXGaWAgs54tBzRoUT2hiHr01OqVuw8uLJh6NNK5Gdyp8PJ
jnjRbJCP7w5WUc67XQVqkypBszuZpMNz3s2+eXxLWG0b3Ifjer7azA9H0rioFMXClC9vNFWfLtE+
E93ruQTnqT8fmL8wpg6Vj9qr8A6mVNzXrG5KARvl7ouD4w+L4+fOeQa2s2J08tm1YmqyfRxdIl/j
Fzonfu51G8eyZTHI5UmyNDVJtjf4G8joUzCQd1/+zQKAjaDmGDKvoW+sZp8moU1IzefDs+TFGLxS
/kULYpu4kZhQe0kv3W86KGIM0EWLw7eIisb2fA8fn0wcwT8PPQW+dABeBd+HDHi8NWGjFd++U0qc
fmimJeoUYGb4bg1VSKIXqSo7WU6cJrFIcA8+PqbIOOZOzG3apPcAFaagOUY4i/xiD5S58inHPl+F
vB21JQE04tNZ6snJm/ouI4o/vVIxqAwcLQ9W+QPTOY6MKTF6T3CVQQ8xkFldJ3REFZRpmkqrbmb+
ruU3gI3Dba8+OxrRKRe8W39JWKPPkyu5W6uNZlIhZEQjVEj9AcN8ci/g9Dro2SBmbTPkeqRIZUPN
dQenQB68iQKvu4bvvVVXFJdik+rRx94QPYNdI5TX1t/yN6R6y+ktcIatzoe9+RPxEYr0LtAyVT7M
ekbcsWjkeoX/gXUwyPgv4CNqIzsm0v/cFJswub1DEwB2EXSEYL9VgIaotBPnb620ijqznL9GMOFp
kRcoztUKdEz0Ny8flQJ/wNyvSMzKma1dmb8PWvwUuXQBrJiCjf+U4BeueUAYPHaMQC87JnXSu8zO
pkUXpyxJLk3I/KSr4EiBSXax2eEUSecTErcgoVJJ+6lt892YnuluGvFxHNj03Mjx42pNZnTm7Tdi
mS1BFymapsINoltHQKxZCveiM1cnFJVQuLmcKND9DqaVioDkP6Sb94LmKYZ+mCtYPRP+wzYpY4cp
237kFNN0D63ZGW488ykoO1lLXrELQSm3PabQMwm2xKL9YvSz5NEz8w1BED/FferdZx2kLEXr9SXd
KdFGgFL6igED/XVur5ont57GVNUNqANo0+6aji0TgcpeWpalfpugURj/r3gpB/X5PHaMrKY6IvvJ
/aYVTm6xs/HenH8UAHIK/eKd3EYw6xOVrWz2fQ0tkGnBz2FZpG6zb9NCCKCKbXPb4MNMpNEakD/t
sGGOBWOsG9vLXEtOIwhnDTz9zI5aInX/zjxxH8HUb1EIyq8oPQykpJqURJWQKDaYLy8OeDPprdBF
bWgb0s4/asAEXYDSdRkbGqaRzKrNULF28SR6NJ+FtMSUbmDb4sJ08H9CZQ1mzAFo46H7Cd4efCm4
RXAKvW8DiThUBANtAsoOILpRgshTvvHN+VjN/eDiR8QpDkXjBnl/mRqAmqE9Uh551jdl5Ul8FWDq
tZmQfe6BWTc9on3/xpqkDSxZhEl36K6LTksqj7hkChJtrnMsns/B+QbvPEZTXS6jQOelOUlelcMK
I1BWvsHndPcO45LrFyz26qvVrxsMBMTpI0hYluyGsKV+rvvNZLguI7QDudNYI0Vxn9uLasWcd6ki
A6TVg5zGk2Fm0zuZKM4hWKO4YIQwRLG7z2qfrd/omYZZZYcxbyr58h6fVoJuflmrdksPtEMHnbH2
c7U+qm4ODYUE/A8cOIEICmth5+mtCAv4CLxieuEGNh+cYvMTP+J3Kiz9SImxV/DVYSs/rYLUIbzS
rfE0aVzK97Ic3WnBqzxlx4dtYgUMzQMr5CVVf2YP+F9jwWC3nYoORKC5a3VyT1qDjOnLrd9Rcjof
xdbdXNF/vJC5wDVLa6xg696mrf8O0GT8FF5rjf8QF4GDEclBTGZzV3RnxMVrmFYcORoAaJh7iTA3
ClUQvvNhQkREI9wzXjpcuUe0BTVETzzijQ1Vc8I3Y2F1spA88LBa0Hwn6ADX4pjYdqoHCBse5zv6
mtW4NiQkgjuyLzFH2CQvuGpyBM72ImUcb42kXh2YzbITxNipzrD/2CogqxVdfuRoQrSv4z5A5uSU
vyKHDnlLUItVrIfZIqXMYTgie7j058mvVTcbsLXsgMEgB4EC87p6ysNrrMBw12AjBvNmlz1W6+h0
Qei8wvmAiyoHT0yBo2eHrpLKzhxeh4aAYV+rCUfnUA3kOf3vwGk4iaBz48a6t9CFGH9jcbchr5za
bU4G7AblcmG90X2d+3jGGt86NjD4VNQi5rJVfwchC8e07wSIe5zMRTYsz7+DxhISpCAqfv1RsBbZ
K08TXQD4lW0u5z9x9IW3m8Ksbw5J4PLJ9WlQNUItXqBhdINzoZzuMuM9a4A/ou6PQIzOM5+YCtIP
s+vvkA/9FAkCiqsBzpOtbwuq5KwLvUh8vXjhRVnwFuPVBUmRyu9v2EmqNaupiMeKoyxiALDJ92XL
jbN2BgNR5D8gUvrPv8JiY3s6tgFOHNN5kjKxRQqLulENvAJxvszLYL7Vk0Nmq3y2UBHzqTeHQ7hH
obkRL6aHAOG4LZ9Ghz/TVJQ0q9T/MccaUnXQTLleoaTEoVphftgchMpUGNG05x1DlpOC6lTqwg5K
4z1P1gl4CUJpSkB2n418rz55JBh6GxJpUhYNKncH9oQDrJkIvnSb76QXzntUc/qqQ2DMCTYk1w6X
ML8A627DnnXTEDTFJd68MuGzD1jJBTUABx0X8ZPS30+MuwPKHu9czgYY+jm6GJ7G/YKhN+OXvY6N
GrnI6da8KG4eD0WD8jBcrxfwZj+p3BR0XxAUE5BMB8uFrT5SdGZesf4pzuOPjWnUhxz5mNgIrE+3
8+VaTwTM772EFeaYZMRcLy7/nKTGAIjW3CpaOSPAx3tUdLvB6nrmycH+yKMantRIbnhM5FGz/k6g
5oFODGXLAvc5BYw50/j8u4WNeU0y0Jyuqd6bz1q8VihrK5+pG0LG4jG4qXO6h3yFEkJoB5HdCDwm
bYk0C2V8eLubXyP07NQxNLXcscujt7/l9f4bJ0Lp+vVYtL+Qt9oLZ9wLO+DPKvgGa16cb13DKN2C
BzEQpXzzzZ91lwgVXBvoVD4hFqcq4A/I0q0HZEJ02FQd79gZFL14jB/7Y0Dvbetk/DnlB8ipEsfI
9CgigEOOZ3Aq1wBT2+I7zda5oIlaRM4jcabuu3T2+4Eepzcggmiee5YUZhO7sfUQ48oMG4V9/yys
4PTHv0f35RIIQ/KzPyFDw3r2lkqO4paPoxZB3SSfeKvYgOxPG7lgxXm2CHw+aPlAYZIExVl7HDeq
gVR0qzjClFH6u2/uN7/oPC0oDlsF1/MBi1aYbqE7NhPMo1q4oa1EZLRikeQ6oaS18EkcERZ96Yey
LukTS7cP7UrCdzorE2li1L3M0ZfOD94mBetp7QameTT41/EEs6E+uJB7fxcsSeKjOVF7ZXvMK38Z
IajjJiXI5doZKkzGKKYappjXvhbHq/6IPpjW25oB8fWiBcSGTQucDyAdM6hGxVIQgkdRwq22Zqwd
jiZMeTCHQ9h9MAQnTFjUisR+0OLuQUouKiV9hFNL2OBhC3VmL/TqHcXltZkE5LomgjWpfLQvz9h4
gKUscAY6UpfBJ/rhQD7HQO0uTpmN3TCy8rqU4jy9UFiuPZpC/skzzd4Qxt46ZeXyDM3R3hR8cXtk
v6aKRbUcc/cARortH/I86vPrMzeeXgBy0Ff+5IP5fGGkeQcKG8XwDqXwPf5y0fHBAvLDZI2VWsRD
Ot8JNQV4GCr1oaJoijkt75dlh2+faUfeR5XQ5xGmcHOgOB0gbHzDbz7fDBGIN445NWOuX+CF1IR/
DInfmUvSBdJNBHyHrbsRo6UFwOxxZU6aI/4rqzrrNGs3gQyMgeciSBZk3Z1J0rWOPKpf05myWeFK
YT7FflMgG1ER83122bHbQVBB5yPF4TCS74C/c8e6/pmgNFgh1rJRI7+ZHxeYEIGa6/HUMaCNM1pj
gKxmZ/Ig02i7b/pvrCREspkqTRO4w4Nko7g2B1afPsmoqJUQOWMjctnCMuAE6dYDXjJhRmwwNA2P
Hu5qljfLtn85XLsYhJxXcE0v1smoOmj3LB9n2BODiFqaX838rCjgqcs8SHI5ZcAy0dVRKgoMUU+s
wrUlocAf53KXxgPvmiylEFFVV3lkVazyqvQmjbjRXf0R0kEUI68+0e1Sk/c/XTQjneuq/3cl9J6P
asRY4+a+eLC1KE03SZwDVQNkPyLN4lJ4fREoSGqD52r1B8Y09DsDjLory3/plHCODA+/dxVWG1Ov
5PmZW0j11baP0HTlNhCWonzueM0JKhgwQNMHgEjO3dJTj/SRg8Tp6c3QURqn96N5lraOgEyJjH1m
hppUeVAntonmFS3LIlhLlqLh+B2XQe+Eek05ixk3CD2XEi3NHr1oa7U6uCg3J3pyfloVO/WHShB1
oPstoik5etkO3EU+bwzo+C99mIi2xstuZCBzS2Ugj5JKCtyYZDD+KsUimUr3t2Im/lGUMfQAX3l1
4tNV+ouBgbtJu7AqHDmucDQSeZ8XPaqhUczol8mtWE6N2nCoSe68VxNZwOoXqB6QWeoTWsoVSEos
1uR3kj7vCwY8Bt73bNe9T6pRgzy2fIgFThFQsiQzGo5naA0Ho8Ao7PfGxgrFyOnsePSNWfluU7aB
nobzvW9J4qQoSS8jIL0oLNd/jG+YKW7enIhllA/tXtR024REDB6ep+U2t4i6mBNb4DHFam8gTCGp
cnxR4R4qopUvU3c776vzTgWDadsWZntZtdl9yW3CMXovLCrvCo1WWN9f0+ownEbYF7MqcpY2gfLs
9oIuTVxhspL+Hx8HYLOl+lweinNQcOmjRYmuYIK8kalfU3lXCEkwAiSGORbKDp/1WpS+/LAWPjXw
BUvdDStAHm3V97E9RvWBxFnU1FldThbinFlM6F62930kczoXxBNuBqGORJ9spdnym8pIQkOLOzGr
MWDxZ9vSinq446oewMDN+QMDknVgbUMmZlHT6AGODsZhJKcOprWcYhOj2bswRYWkWwyS0lHc6zqq
CgpsdD7/CElObfjOHr6lR7ZNl5qjku9sudEFRSac3mHMYIZwmAwhEKemrwbDzZaZu0ggnvUcVsOC
z8kZsyXvhjcf5cS2BD9/sGrH5k5EAmXEpBRQ3d2PCbhF+hEp8U+j/b/yjHFef10sHbSOQDYsCday
w3cLUHNNYdCjXRB3/SHkL262G1oYFofGnzEcuxIuosIyWFYYmvR5Q8geD5z+8vU8ebVId2SpcPhk
IjVaOjrrw5W7VC5u32XeNQSmUi7fWYTPlLIXmpYQB1yB83l8ntC2NYMMV+Xw+TAQQGpO6/Sdn4Xo
9maXTKJu2zeE9XlzlxwFkF9MuNAlQXlNno3w1e+N5PgkXKTMmUl8+9ZrNBXL72a7fqTGYkPTTdKS
wkh+ykBZCU49J2s+g9qjxr4BOri6KhF3Ff5DAbtG8g2TZQtJbfZe7pxAQ9M+HuOmOdnaJGZdCA9d
r1DFBwLVGv78bfhpxVv725zHBHeRbA3vuHmVWSNWG5A0JrdhvEc9N3VrMFZW0TIUDYDmvM6a6aCW
HHVVWcUzyvqNDRRHE7ClMG6WTyJRhEsb7cnVs6PW9BNmTJIfmgglT4Wf/dDG/wpL6c0AIYRg5ddO
DU562wHQWCONj4/YSD7jld9iEOFSHtb6WedxdHFNS6tuISaPL+3Qq4e6PaT0UTHPnEJvteilmFny
DQ+Ie/6JaveeS1Pr4LMPkqcC0pEfB1EqqzVnhViVFoE/PH9N0p/TT1L28mEfqchvE5BUCj0rvr6A
eji9jSUWB702gAtEZOG1qs401naXPWwnmSgtqG3ZtrrOHYcigWoDNEbmmZCWeRrvjMQPDCVElBUq
vkmh66WHbV/87hfHWrZmrAD4xXYVXGWpruH5qsk3cb66X+iCYsn9zXeqf1UnYNaeYVQmvYROwIqf
CRbGSTy8K3pqZ9/GQWQLa/QnKlijLdgu3BzaMw6V38OdlwCNfpm59Kl75cHmNJG33/WLxiiWIzia
GWUH0fhW8GdXHIsBREwvYfOM/zGoVrkYkLRJ6w+SxXwgPGhZjo1Z2+pT/UnAOC0X/r8VMpFmUvPi
unW0fn7a6y9H60hId7Shr1/NHvra3fF/t9jRzdjfhJK+lB2Nzj+iX5Zar/+7MArkw7Q26XQTbSlG
iBUsumionBnQ55/TM9X8iPlF3ryWjuG6Ef7IkK7ltQifskoG52jwz8rAvU8snJzJ3snUC3L/MHx9
6rePpaDOrfOQ1+ivQWdbEYYyHHisEcT2ae14ipC1qLNa5IO72S8ajuPABLlmsLMr8c6hRuFhC98K
tBwuVtg/Bx+y6lgZnp0posbesOhZoYgpC8yKhBPp5m+m+MofqM9LqeiMHJYva8kSk7YnIboDPpJ+
chDcLBnlrFcMwAoGg9HTiATvVujKicyPgSbeK9JLLu+inKqX98Xiwe1Ws0zgIHiZKkVCqfPxXQzo
6khxum5gYItgm+6f/WHmx2cbSFCHrUTPpJdaP3G6jiZdyKZGAC7xDND5fopWfHPjZltMtxx6pzss
t8q9f7PTSYMRf0IuFKX0tL/YdPV0Y1UspotCK80SnlXiHAuhMhA2S46+6fHhscCgJK6RTn2i9jma
0VU4obIfb1+sZuU5I8gjRwv2jFUSO3qoJ87Vh7uR3zQGmb+4ZloijNUvHlCHzQfvtPvbX9P4EbJE
N8Y53e3mL7Mc5uts2GZkXVS9FALdb8OKwF9hC7jaO4+gC4BvxFCjxpsaFtgpZYxp3QPVSmpWOkhZ
+1nUrbOuX0CnLPKRlLfCePArezY8zg7YFl3xXIzFDBG+gOGAXN4udrrll0XoOOUwCJB4AW044spg
LarcU5RZTEeLBPSgih7iOTf0WXO4G8nmUOnT7CHijBaUViLmvsqAF2uNLOLnr42CEhZnB4pEyuCy
h7OhwrzM2P138nVHUR3KWFHUGO6qKpV939aoWk0aULGrUIj7lT4hLACk5o+EpybifQb3yh18VYXI
1G/Yl1NB+Mpu8elwE1RkraGz0Lk/SAWlKtOB2iEM9eceOa1kA4zwQbxPWpGG9PdUyFxXULDdDG2S
LSUa/cmz/PjFPV7AWH0HU3qZzMY96MKCCuWw3J09DDBuwf0IiuUX2kzmBAy7xdxblDfHpHdXdaR/
Fbe3ODYLJJvyOI69SiCkGpdCWL34DsZCtIKs6q16kHjj/UzK1r57UK2ElRok/YU5KnhNhgAv7jvC
2m85FoJGo8+0iV1uyKq12xHiKJSlCxmD2BpUTqMJRgP62S/AzHWmhd2hNsdAavUSqYc+30rp4f3F
D7ypVuGKDJhqEDh1ZA02sr+DczU1RyppPtc8qGWdyIheJRKRU5EH5cvXyLCF3b1wXO7jxEsxTzis
6yglt0V0NHtXMXyId/lp7EpOx8sIcKK7e6VGkgAJ+xvbMIQCde9FrhFoO8JQ5lzMIr9Q6NnehOGC
GaOdYcZoW32i+29QftID2UEgp1SQKAVi9YtX4eiZx/Z+O6mTrXx44EaNQS7BKbCISFdkog00N80h
shSNPzyTZsitDRQB8cx2GeWaasd1Un/4HNIjsAixx54a8zXEQ1Jzlbme7tRPEmXc2yaNAHUBSUxt
Y31BPnJEgNMUU5HU6zX/peYyGmtuxxrxj4gzQLXtolK/WPe6Xklf67d67+pq/Sm04XbfVauHBOlc
0DpPdjEBLBQaZ4I0pHA4PBDUVtahS3xE0FbvG7osaS8PbmI5KvQC6mYynMh2XadwLQ0LLDh+mlnI
czE/0Y8IKW/Rdtn+2f+pNSpiz+8AMR49IiYAL1+Rjmp7Gt0bBFv6mHwI03IaL/WvR441SjwBo8y3
/uiTu4ZKJnz3zD02ENbS2lSy+JVteThUzqcDZxDISB6FkTsoAxIdUAtKIVCsfoKhCuh49O2TyhiM
Lj/nsftLZWFhhnUFvqIoy8g4+Nx9m+qZ3MynlhdZClkFsLv/Uj8tpcLDh6wtj4ycJwCyqfZE/d8f
ou3tzom+iuzsIxQ6NEKF+F871EorS6suIpkgjuuEOPrvOp0B439G/kTBUChpPDMhuPuw+RsWB+z1
7//ZHPVsOBSTgfT2p7esWL1e0y8dXRfn6fngrMGUuShyE/TrGvFmLrAbYCnWvLRRZ06Oi+vzcs9Y
RIgP5SBH4RasDWdUwF/52qEUSqqjx8rgfEzS3Y1f0qQTM8qeBsIBhPw2esM7D4HkrBQgMwZF/5iT
fXSFHYv3/cE+AG/y8Y4k0pBQBVsMUEq6UGmp45NNW0cy5LzJvOzuKxG9XKZ8k01t0Gq9LPsFYl4v
ggaejLmozXOmawfalltTDoTd0jzuF0fUenJkski5bUgxjH2Dv9p3o1FvJ8LEruYbu9fmWxCIlaWB
ZEmVInsOser2sqO75PzVbORVYa4khUmUAmWIVItur2WxtxtjRiARyAyEMszyXVRW1m85dDrpyMje
enSCsndnAhF48ucHJgTuUJw5UgnYdmzwHp/E9hT5Yq/pqKHZqVr+7n3ViAZazznUg43KgdtDmx29
wfmUFBtXRZB0ffLYMeW29H5vWxVNiF/1YOrIE8VFtrJMeuUxuJ8UkUzdpP2FnOjmtAqBQIHFCU7W
qSad6JiOXLEoZ71TYhxO3xuQlv7EtaaDZyW3a5l7UtAF9quTtffh/Mvc5XBBR00NCcF9vyPKahnV
O/lUcBGl8SuQZaOY0LCSUtr44NZcwg8DL0hwMRBZfgcDKA04eHFchtOACA0idTFYLgMt6kvq94iu
sKqEZdHhXelUma69wmki9hihLJ+CbHpf5NqHZrEJlQ8pEg5yl0ssLEjb0bbY4f/tsT4mvB3ouBvn
+z0cIgt9LWiEscKDAkONakHVC457+moB4RxNA7c+6j6rPc/IlkwI0hCsCOw2rM555IAYddvrvuhe
muWMDsBLkMar88Jy7XCGS2ZUkUVj3gVL4lVLz3SOeDXbW12gyV+hAiSOFKgsZ8QsmCYbNMHa2jHr
683QjzGXyfeeJ9wUnWpvFDxuF9X4Yd7kt+d1SYxjmtV++wg/qkhK9clihMP222htnR01KXMYl5Ie
MR3pLBYcxC+EuuPChMbEo6o5ODoCBOKZjMULnnxpxdIlbu3jQZGk3EQzVR+IM0TotTPBPIR7cSPR
mKBz/PZH8yLOKeBnKpZf6A4Fev1K0c1j11gu+aTjuoNMjPLf/gIS4l7qIxyEq+laEx0+V2TQnw21
AkXqe+5bTc1TWRhMl4W7M9MlXJLW/bcdo1mEr1GRHdw0IB3wZlJdvyIvx/4v7sTOeWWtOog6hueV
8IGqFn7Cug+zvtQju1sBMMtF1IMZDI1q3vD1x73rrThUPEXNBaR87atplfRfvwHSHZ/0SyazX1l4
NiErYs1Z1RkIbLf7ddgxcqQ6BoqMH8EpK4LvWuqh4V8/79JGio44dcwSEKZoHzr6osuBcQbdDQt3
CJbBaWoOAS7qWVHyhjI/JhVNLMdBAc3VtbLPpzntdnVZr8oIEe6IamaOlNn+lNnJA7uZOGS39s8f
1naLfwfkAZSEri3yxkDUB3aqKO2ipB2NV3YEn0DFnfF9lML0Fg52WLkAr/oledRAfSm16ILCwHF7
9bUlm+lV6qVk3wKwbWA7zJ7P6dTArqzmSa0e+WIdmC0+Pjx8aE7RY2BWwMsjulSpsCPUH2VI/q34
upJ972c0jq1jeQZ1uPCk5inlC6LAu/m5qGL9JJSHNCRHbKqC2X55KdkG2ujrePOWwiFn8ody1jhJ
1lSAUHP0TOseXO1QheAcSJcIfz1prrno+WJnHrgUzeGRsHerpa2Ro2X8nwhzEaSPFrNEb0eh2jKg
Uve3cwQITbwenV88+epNfKLTSMaQfRjc5qekWAZyGrc5r27Z79ITUXmiJV6W1aTp4SRchsAPRyoS
tDjsTIVsKtzs+l2bgdd0yB8jdoCyC4bokvzgK4SrH+g9rIWO2J6EuCbRK3zoWevbGo+iB9l1vk26
lp1zoyYeNKW4wu8P1EI5p4DIAsYPwNBlasTWfRm6tAJwzqrqR8kWYe07ipgpVtxN+RF75sU9g0IO
OiPK/nLLMhzcoAWDh+ZNwZicSO25aIMVFp0mBBtvJwNazthUig4X56CwSOPLmZ6t591+plMi4E+f
qSCAcohImWzX5DF08S9BYCApeskV5SFWThP7Lk3mUW9UX4+Mb+QlZbxDGdcuFJeYxnhL1F13i5Np
59UzQu/gySH0gom+KJqP0TRE3bz20eBBWLvAWw4ssxEuQl9726YsDzcH8PzcPqIN6Qq+zhau1XIL
8S5N92Uy18r66xHedLXCTPwybO9etOE5zzld25Ck6OTPjxd0KmvUywY0cVmLkeOY1NjBjCRmKSQz
nVUkAPYY32KmhjGuBW9w5ZMZm+AmCIowIX41yAtoOZnEnUdSUKDlWUhbm/h1W2jpMcWNqYCpYjF7
/Iudqqh7q0J99ZcURbGTI4qoqwSnN4vJPY1pq/IUtz3gIZiPWCLny+Beo5DiUTqYNzd3BJTOv+oH
CQXqy9Kuv2Adx/Q7ygueo1bQ5D4EdozsDzH+ZDcBKDaIQQt38t36WnKrFccBFESUHNDAZ9CYA8H2
G8M+sOC+GsNVXpYLvPHMbByWDtha5H+00i1WVFOU5Ebe9v+UcpNerXkxWVsgth7++n0r1FwiaXWv
MA1fZ51Y5eet720I1Bsuvxnjy37i+RlwScZcuOzew80wyPLwKBu+fpFdLvnEkHCjJj7jwoiz4oMO
y6NthPLaWZpz5WHGjSGEPFay0yqw3w1QX3+JqoVtYkMuokJihGMm7WWNk6IZYEBWrlDqw2t6kjQN
aBt/ZkoCVPLgyTwUnnoLAmWBdtpopTlQhx4vGkuOI4+j1OHnwCBm5Fos4NoehEhP6AVH9d+RgsOv
eUErOJaLo1dEIkATUxfTTPB9C7F1I8gag2SZMW3cCwlA3pIf3tRPbuo22YlvdpRzP8w+7soK9k9h
3oupkCiIeA4/4N1FidsBJoHBDdPVYWC6GiVEVwLADE8KYPm9lN2v77N3LypoJ3Su4j072PD/3OrN
zOm7o98f+H5NYLIN9d56tHENjptJKq3evovjl9gJDuM+XZWfBeQN2UuR+6nJH8VGuTSoWy5LmOH+
gy5UtLtoBV3EP+tTlKGty4lQv5SpMQjEeL2AmAQl5MqX4Lvi5yeTNS2gB1Ygx8LMAr6O9pIPhOVZ
7qM9wwijBr22g2lWJcsKn3OFku8yQZlTVqAVede5d1DyUSpzyLK3PBO1mBLE5r3B53s6VTcNZW3l
EniwmiZ8U5+eyKX/ONcKIZ1gz9ksdLkqeePa6fWk9WCKqouFbh+zYVgQ59BkbUS/Up0XLAX01yZ4
xp+QkrXgclKkIsnQUN7djtqQBqHW9Im33zeDvMOYB2Z5PL3AXu+iN7QI7nm4tkBxbxrC5dJkw/CV
/ZFvs4tCUbILtQRxMhgZb/OtEG5x7CS7OunzvaE5bO0iCgbRMRumG+JLDwcVMQDTfJG4M675zPkt
RSsygKsL+bDQi+nOqXdFkTYK0/Bkf42djy8uSSuyFG4+QYPRr6PTG5Yu/z6ffRaawUddQM0KOJvW
DE3PinaNW1RHDRKn+A7XW9HqoJkMXinbbtvT/tjs6o8tIJG+N5lTmbFTh+qpCU1iSEE7zJhoXn6y
B1aixEYB2s9AbW3gXfPsOL1G2/3VWAIJT06BwkBn3KxMgtj8kvBedpqLDez3Gxhlz0RBRZ/Lpmc9
nkQu3rm1m6NpIUENV9dlsuL4YFVtDwBv8U8wea47KezVV83kdpHxGm5Ju0x4pULAaV2FHfGN05w5
TwPpkW281yEv9J0YQ5xYR0ISu8wo7ySMIIXMg1pE+ABcbhdVb6YFnInn434nGwJz37EVTCQkMxQY
Fbc8RcRiSNUNcQDkZ2PKpSjlZPsPiz6FgyiH+TEuglPxRPrLslvkzmcc1EPASn1AznVgxUbnCL89
XQBjJIx1dgaMRFGsJ6T43/3DDCNZcvX13emK9+Z1Z6s28d60UenF6I8nK/Gi3DBm85gR0Hciyt9u
uXrObtqSciMmFj6/YNRpLGqWzeVCDQKz2WTmfSg3Bq/K5cOkXwTEmSTbq5ZlIbolJg7DSPmFAXRZ
/qSSMAF7f4Bt90MFWMRJ/OI6cEwLmiglBx8oISlkT/wCqYKVw5zEFW7s4cCb6FHkAlRVdCBT9coy
drOMUFf0elzAmjUF6JmH6gnYhpe3Tv2C4Fpuxbv4L31TzC7afsVzjQRjzePKgcVnqJW0U8yHwtVw
Ja7xDu/8JCds4GXNB78qkbLth0PyOCa1uqwWMCRwFHd6YRtGvq+MMq2kI37XJNtWNgdRbwvrsmfp
zJ3FF4cNtWylKDr5YxlVhyv8M+Ru9S2dz9kREqCozn+F8Mp19ctWXLtZEuQG4UdVl2HSuYEiq22H
wdD8QDETkK6lRQwWkmrRXxrb1xTnKFVqSoPA0y2ccv+NI3lKKv/QE6shnq6+NA8dkr6aTN1sZqjT
8hfzJ/D+c8H/eqJrTvM5rYmNB6l/E2jrX5sEA5qhErpnJVu3JsZ6dEU9uc/jSiIrECi8VfkWVdfs
xicij8iNY8P3dn0euSzXIiBi8kVBVKOy7l5NRvRpRdttQZQqYC9srKRsDmAFjbqHcSPBamMB0TCD
oTS/XWYqYKrNvq5G0tf1NcCDvofR/W/L7ghpyNnGpT/g5wi5T1AEaOy+QzJID3rVGhM2F4tCtC6/
GjIaojWt3u7j19wknsxfzHZKAQWVsnozE/hbMZ2UDYI70KiR4AmncynuhJ2vwXjUpsXjHYvMKtYA
vjcxBoWYKrL0QAkpbGzjcJeEEWEKtzhvDXuKsHgmsGv9OEjilmK3UWPxm6Rey+uqROyNmxNTqouw
gUKwZZWLJIhP4ebrOCtit7rLNQiLWzALc7kY896b4TH8JCuEmtpRFEewR6nepCbatFdXlNuRdbuX
bD7vkLRu30DrwiyBAkhyAdPi6sdCrVve8YDbXfh6u0/33YYVRsqVF3fY8bNqJR1BdljuA62HQepL
ln8WNmiJtgl5lo26/Dqa4yLttTFbj5+8+UoLygGiA01ZWpYOL9xprqmfOBsBExIP3WxbAejm8dUv
0lSXM4hznnigKkJiXYbARtrzF54RhVWzFe68osNqfu8xjh8yhkOrQ2RHwCQMVoPuNN8OrQGRispV
Cn2TruAvM3BbVoE9gPLSs5asdD0a7ZY+p3ccSd/NN4aW4nFKqaa/bPsLSsqkoGKuMTnUUtPepQZU
a6M6VFATWa7O+cfEL/x4/pNPZNW5Nlvfpx+tACdKsZFEHpsC5AnTpfYuJhHIg1kNl2T9OpC2K5R4
Qcd+RVv+fJpSoaMIVjaTeexUhSy1b8b6PFIW1xQThjLjohcTu/mnt6nYhqe/ppfGXN50NLji7xs+
sK2mOZAN0LezPa7emkHS5gmmjktsTiJ74w+vf+ZO993DQ2hiWVIHdV68T9lN4/nEgpgFftXuYFzT
rtA/scrX3p8MSviU7RxfJ5YuMiPIDZ+F9lIGmhxG7Iz3ipIAp5h6PcgNkkFwNdsSfM/C3leGKypc
w6lBXeb/6vmWJNMUHidii8ve1gm/kDshKpwjYejQP/Ux+ZZR+UmB/1d52GIgYvWNvs/dSDgGilxE
O5NOlKcuBpZPmSdNsPPgmTplbs8k/1W2oJu6AKV0z3JQ6J/g4oj/VPQ6PzIUyoHLtg2usn3CMUAM
8/Ev5XQuP3PLE5o38BmSjj40OskJoCjdidTKC6SMupnDI8gXVgDn796lbftHnS6U8Tkg2YZyKh4X
4qOcdEhsKGogv0BICWzO7xWAH2j9T8eNlivO+Ko9e1pka3AUQ9vbkSWtT3FjqyVeB6EiUatW5V5j
llwIOpCEp1Iop3DhNsTlnR6r+esG+HWEJN8c9jS1yR+27DfaFT7XQNiLnksv7kG0E56AOHGIE2+V
fAXnQ9zSpnDqjsiPAC/YCJ6BE39+TbAemHvj9dJT+HhUHVLgwQwaZeGxbIbdj18KatK60C2Pyiwd
aHYi7uitUrKWMU4kE89vUJLSj1uElHkVE5QBdWb1ugAnHhl2bxN79PYqC6ABgB755HXPpg4g0FKE
T8L6h3x26RyJy8xO8YjnUIGsFuHwuq3pXNFq1ZdEiAPMdc8JWLUn+SRy8k7x6aA1hpjSjMH7mNCh
GuclWJ3lgkKg9HWR4zNBl72aZOfEYEASrHABZEMfTQbLvCsz1TdDrZc/x/+jfgt3cp2iYz+tutKa
CTogn5/7Bg4QsQbXybtSs5BubD0q0lkgn2ISbKZl0BdazOQfQllLRmzbXLFj9xvwhY7O8z70o5jK
3ayJzGqHYsOuUisiu54e3EYER+86jy//ow48D+rHKt5cp2CJ9PNdWcQUyFlSHOIiUbK1jAjfLhf4
o5QQ24SwDuUFAVVp+5WwS4G05JVq7xNyonWsesGs2r0EC+dhjaU5SI1kqs/06BcSOjntbs64FjJa
aLzhv4P+lh2VRN+UwYN99QL+ittfyibbmffY9y/nTnlgtU2M0whxfw1RM6oZLG54igiAbV7D9ddp
e59Fqi8ByGEObERSrpv7RWLuPAQ75nY4Ujp+iVYkRKJkmFdBSfthpxbUW+T9nc6TV8z5RnmtwKRb
QIKI25AfKiWNEXFr+5JS8bEwoli9PmwuQMD6vAbukAfwERQjeWxTNy9hEupVhH/QVgRp+6R82dfI
HNonTuAvPvJ/Fr8TSYOzLNL7Pcehmo7EnL+9JhFnJwKdHSgCHBnzHSV/Xtmp/iudllHvP5nwiwiG
akhjJRHNkRrQhc5Q+k553R4PY3BE77+lO2Qbkj8iF5q1LGwNpJpn/PffeI7oACEPmxsC7yk/9SMH
24pe4Y59vgkIy9hN1mF3C0XOSKgmHpeIQIIcQsxoRmpOu6duFU3WNPENCOOyR0eQWINMLf5ybzkq
aWNihTEVAKijsT4B2e8iwySxwyHUf36IGoq4m5sOtS5diFomM+jHQuTwvVKcDMkwdC4gVyJsxCBm
vPp1chDnm6LZTuJ+TRzuPubxPZF0nBK/cfa7lyRKU6ZKkaSvOlIjtDG30Tzew3JPxo8zsfvu6ME/
yVLGyoNpw7ZFq81CTDCacHMNlys3zHGr/u/svY6fqs6GyLw31Dk2N/laOV0xdpJpPapN5c/vef1H
xzPSIqdI1BtX3Wikp+NHzW82JdAbFKWKEuyDEAvM9HWksc3mFU/XUIskq72ifu61nYydAl/SzQJ6
O2GGbD6SHbPyuFUtBAJNmF6LGke7rKLlv69L0uS+jeFZKnHub6gITHABO+cmIkch6C8/oNNCkzpV
ZlMTQHHICDZtGL2cPyZFNqfd1YApoMbKn/3bkI4BUqdHdT1BeYkFIK/bl9bEAVenrG86HNh3Hkd2
Gepprevyj4rzYrzqGpq3VzTJx0A5qEAYl4zfEjknwyhhQY7CAOf3g54UXwzzgFxg3/r16UEq3TiZ
28XzrOP/DzsalDbwPxUJsnLcD+Fm90M2NjhtUIaFP/NAGj00R00dNNFWFid9yEgsJ6cjXR01iLe/
4ANoexoQ04yaTYL7PKT0dAZn0no+OS+rnGA/R832vlxAQvKo21JgDO8hWzLJDNgQS9PDQHmcm8M5
VLocNbbYrAoyx4Fy4D9wmxpIYqxwlFAogzWFFoq/SBuSn9Em0HsfupykQKsKs0kZOekeO3q3ltU9
TxwUkKtp7P6ZyU86ukvFxuqbmf06PBgf28h931iP9t0YHTPMNvN0R6S5IXpeU/rPgrIaup8XNAcn
FMASXlyCOGGDn/ZxQ/0ALsRH94Su1DIPuRi3bni95qZv/FMPdpJ8hjWwdslGNKfKo+K4MHkSEcHG
tgFoA9WNw9e1xFxO1XCM6yeg0pSmTJ4HgIBuALBxPrWr5Gk7P3rVGgqCVehUAEeMUhUHOpU2f8Wv
sNJ/SRIauPSynRXoo93mj5Ez0bv5pu39GGhNjcyOqQH8UGet+FRDwP17pGO/6e05jVBTXtJcDWi6
8vVqz10YQBMui7fUauCmRH2EYl0uYZsPKWjUceGRXkvJxt0OCSOBaNzfBxlhjCfCV8KW40AFC5sS
THZl4Q2xg7sGZ/tKoDKPIYXd+J7HcCdXZLLe7RVv5DqYaiqI05X4sPb9c/kaGMb5sgaIicUFt1/K
GRX2mOyXyBUio0At0diS/RZRGEYsEowln0kW2MeDWPH8yRQyPfzwSPENCBMZF4zPE4f5rpfN5Lqq
S/ffXuaaL08V+aCcE39qcQEKthsmnNdC8njcw3fLYW48pEOaHcgTG9mPdYcR1p7iParDZxzUJyvI
x9ikyubjzIl3NIgtGMAuDpRxaVU7Ot5uHLZNhrf+YABZosPKKtHhWSfiRHrcPx47jTUXcrcUHf5X
XRBbXzoP5k4lRhIRozqyLC96HxtELH60zm+IQZfbytwLwNcRTqwrtFmx8y7AGMuc02H2uEUqORF3
QphvxsJUPGH+QWk07dByY1ieyFa85cjT66aU6xBtMMjaB3tXG8/+D7byhHXgsnB1dvQUtIfdohLL
hQmt/ZNu2OvLPXYcfqBcaQeaBITIVdI+k1TlYK4WhszN6pio2aG3w3H3RHYHcRsm0r1jHVv2HmmZ
PEZAoHmSY6t0TvkQ76RBdvpPJXRfNSZOHzBtWH8RvPLQc4N1ZZ/1/g8hdnFTPyRz4Vh3H/AjgnZT
whnTpVQSXTI72xZIwxSkLGRZgEp2Q7bFC9ryW9HhJorrk6gBJxSkgoUqqYvWiWYQ7L3yh2bKVprt
546L9mZIkQ2gfj53PleFWwdP+dLJwghu2krSFUDiEGOe/scE39/tvRAgD36yB51YILt5A4ec9o9T
c7UXcRsySwbNShwVIarfmRiBns7TstXw8ieC+ueUg7f74nEprIcEkwPiXQgkAggRV04WQx+NU5TU
eoXecihPlJOXoS7S20U5QdwaCLK2ZUYkiSk/RL85tvhW01BB4C6e1Yo6KoP6OfeUr8dqa4aZ6686
Z+m/0xoqgiSKDR9l4NWqrFMopT7Y8tQ3ZlqbyzZbntvjQkqL8rhPTl0i4fxQtAMLD4+mcNGHJHjl
GrO8nuKRl2gtegIGYqzPcswMU0T5aDWiBhRG/MHqb4njkAEeiqbdPU1dJ+i1lrjNfA99ylbcJm7q
HY4Y3+E5rnegWGc8uO+1Qrc8loj28fBTZAnkthDVlY1VOL7wczGN5j3rPbS65boAupkpQGMfbNeU
2V8u8BUlg50pPXuYmlZJAfLh120MeAHtgAx3h2c+QwSmrBm0A8Djy5YQOWVzHGbh3FnsyLw+L3V3
8BjKl7HlKeL5DieBDgUJm6KKR3T/IB9fUFshNEgJjFFKcoXy0qKJMQe/DAhDa3054nHraYimMwfd
lsl6iBt2my/0Jsmhl8gytRNvACL8MWL7Vio3levnfaYA9yRudWDV1biiIQaFDXKr4KA0qnoeKrTR
mRdxOqOqYHD/vsTgA5wlxCSJwrfElLaeIjIISHKaE+kKFxAG1+Lm1yJAAoQeeqn4jC2G22fncSIA
BAdc2wOA+a+zp1+/MZZI0zJPetTwQddvaReQF4anoxUz71hyIoGeDyDF36IceL68xMpYKPM0vM4+
TaeeLatayR2VmhQH/mQiWj7rHF5LFvT3hYnMG3p+YrjS03ju0E9oo5/JT287MRg/dE/6Ng3zjHaM
VG0OQOToS78MEPwhSJ7iamv+zC9E4y2wHicTWPLhy19NIFcXO/8PeKOEwmgDT8RxHXVQfsMT8sty
YzaPSW+PCw7pVTDZeqtk74GTgfN34LDnxR3+gkCLRwdOy3xBp9PM/7QAXgCAFjssKZVUwJJ1WimP
9Aev3zue0eYnEVxkoperIbAZ+jRjv3feMRS/V2av3LR32tyIa0DolBTsAQH7/M5SCPazT8WONTZ2
A8lS3roCjrvEEN7Th19JHSvwnziH3TAHdgKqDVAtulyKseSnv6KUNC+/RELk9Lp5aW6HI/C+j7RY
83YUmoHJqOhivOXg9VMXPW/Xnhtty4Mvp3gGyJjN29KfYBjCjWfkmVWyx4kkwgSZaMaihzJQbE5k
vcRwUytMqEeBs+G1vj6hQMLauxUUS2ZOzktadZjBBRRzXFDJ4uztHG/UsVC4YprmJGNjJhgHcfDJ
gbtSwXCjI5RcCYU/LQLfib0EqZ+SFPfV7isy9dDtRuR8r1bzDyBdA0YCFfAE25kMVg/kN7JxJkdA
bdJOqw+muhMXYqPt2DA0uV5SS0R54t7V10yynEmL8USLhTKuAKlnwaYirLSeTwHSYUERlpgwZWpU
8yUI42y+owi/2vvMmIMRTo2SVdLLL6tSBJklCZcvH18oWSLrq2dSTzxsHYcD4iMXjnK4L8/Q36Xr
LR+PMBP2KjiCM8gPE4ExyY31QU8qxaBTZWwhTCvcdVRjmwZ3z6Ocpc8zH/zqUfZTeDxY7O/zssU0
4ZdG7D3ZA75ZMr1fTcZvmT7uAOKw2qHmgQDnQgicUEQmwJWH4xvfKm5Nb2gb+ys4jF3Y25UMdk1u
lUBOM3OPmyVLmtGW1kyw3l22w6ci6AoC9Hg8kky9cOFIQ+GT+L0dge0GzI6qVmW0suLfi4k0O5Ph
M0rfr8BcitHfbNrhYWrePDlllxF5Dhcv008Sv13GcGjIxF1WWSFB1F/97gjDVqv4xLKcZ7kXJpte
fIRAn3myOyqdg8Jh6xDBwi52b9Kt0ouRVsguz3khV5u7Gx1wf1QYb6f6dsE9eIoXVLWCN/yXhS2b
xm4bPU0PKA1y+cJdoMHsKJWG0hSg3qgw/BHzz4vfI7MRpGNHrFbAnmOkhALfOoFdrmMKJxq7q26H
blX5bPD+yzw8F9/h6zyojYvCwkhSRVEAuuERviVYSVSeMsRp49dW9l/3a0nhUSNqvt5QJHEhqpKb
Cp0nCuJaLUZXgRvL2IfhFttc+8QnQ/PG1m0smhtVVGtYHEKfs/gsjlyNMTuP4XuxbyoNciycYTjA
MSfukw7xKbkydIhtkt83ujCcr32gztgZvuvbWVYZrYpc6jE307ZaWF0A8fK4DaJFET48SAlvjqRf
9m8PWzMf4uIYJJ+vdhACaE7mDEOS2idimBLl5tZpPayawytAgLkI+NqbxJUpHOLKvPnewQ5yCU95
ipaSNvczv2Z70MtwhjZzlgL6AWUCenmUN51nJH083sSourHLKFdRNDKpI96nocvNYEira1V1xmYE
+/jkUg6zUohNAbwfjnZu2+3N2ceObKZFdnB3Vl1idWR2jVKA/G2WP0TzSRA7UouaW6i0b9waAySg
85eJdwrepXJrowD8ugbJ70KBoZgDi4PSUmoBDMDIykd8cfiqla2ld5GT8KXUBfxatG73HWuSIqrM
v14OcFc7gpYB1mwP814a+j8mN6Ai5vKi8W7+j8cfkGog/RBzzh5CCLfB1CafFSBEyhDp/pSN/nAW
DtPCZ4h+reFsFlRD/BjMR/gYY7YmXftgOtsyRhcA4hXFUkZzQXJ8D9cXsI9vlM7J5WdXeKDZS703
or3iOLjPs+B2LgQwv1YjGeE2w9POBgKk2dPwPBnX+ymONwuWBKwjAILH4JhYCf2Iwe9m+vVEpaVs
TNu9ffPj1QOIT3QE6iIK4oQy0W3EWDN+vrihhWGhAuuzwC9YVpiIAGRz0KNR70VOZA5sTFpisHUo
OY2Au0CKxx6TKUIE+ktNm/4U/WYog/JJq5wbnra+7DxeQChR43hobNyzkdpazz3Fd/2wpTXjKQfQ
k1mcs/PykOdckRpAkHiv0DzFlJTQqNJ6Of1Dv59y01ig4u56cyvlmrxz3I7u5ecEJSIOkWaMW05Y
sQzlJtXdbTIKJlsqsmgsVHevNI9Ovk/15GVFLHzgb5sxGpTnUgfAZsVM7qOupZS3sgfLkT2C4f0Y
gB3TETg6mIsOV2nXFLe6h6JURjhjbxggruJSmzEcCHisSeaSjBaan4lcZ8O6rkka0FiqcK9mRpL5
gAxoTfx5v79PUt2D4lDuiMAtm3gy8+ZTQqmhrTKwVqpWronxvl0esorRpMHrpmlU8Uw/XFKdDprG
lDDOHfG83/keATO0joMA9uB/9lBiUCy9iXAS+JXJBu0gVdlrLW3rUr5qYUbo6dmX44AUz35KQyJF
HGVfvrbIx7a6VnPKhdIXbaxS7ZBzJ23IZoPDdbg8zx2rvZyOHU6cGSaa/LKJMFdkiwAwjnioCe6Y
M3KnH54vOwxnJ63RBro4uHdsHuTtExaLiS2RPABLSPJw7Tmn553BdjYzsY818lLgi9AgkxGCWX0E
kZKcO4X9vJO89UqiIL3ARl8tGa5dN7Zn1SVlQKl6iGCLsrBv88AZEiqRwl7ZHZWqVJZ0b/uFe8I8
nIu+NSXNDK5qe3jZlHkXKZF9eF/1+nf3rq3Pj8xQr777dPcjt9EN8s7oNEkac+fdRVqPpvNYJrbw
8Lge8G5WJv7tHDYoVzg25fdDoSg8U/0QkR3rwVVfw2KMcJ5ZVRbwgF9rHMAmsgoISkOZzovLmK6J
ziLO/iJ94y9D2UOXuSVwm4RVnWvI51pOc+M67Vk8Uw2ddniqsxFpzG9WtgAbmohEIB8zWvaa9A49
AhanbUU9L1GoM/qd0lXwl95L4d29OfzuiAz5fDOecVlDf/kGBeIEhf66gg7sfpzffg04LPrFzDHH
2tkAAlscpp7qa06XDjeON7+kuBYb9Wml4rYigtgfzZzFU7kjtZck+gvfaouxKseMtxZMgtRBVhaj
whPerWyykGiwD5cY9evgR8es9UtRSxR9uuFEbJj5HRyXXvXhqU7FSxjH81KHEpzQwZoso0bibRKY
HY/lewyCmFI7hjUFsfuFEI3iywuXxlVU3P8cE52Fmsx7fl9cyMS0rCZus+pyoafTMqmFb8q+KwX0
qmblGPuJGWU6O+1UFJAnwqtQmBtCQ6ElKdsDDD+IrxV5FT0LsXfsEfE8qqrGE9E9xtKoE8jnQEbi
SdHEuuSft97EXs1vHVhEgw5KYkoQ9Ccbu0Wi2ovw1Y0GQjYpEN/465Wq7pzU4Pr1Xc367wo5++u2
N9oy1uUzYTYci1YFdQgNWoxrEcot644YTzem8X/A5uvC6n9GedrcoxMu0DftxqDu06Hj1oj1/A27
bBBq1ySjuySVLAiz4VyA4tVTPzCz4hglADxL7HnMoOmeuysDUAyWbD/Nb41Hb1QScDimX8FKR6gK
xQk1d/I3hjakLTYzmjDL/Hnkkt4QSEqodn8hzm7OIXTbsJ1ZzB2CjrYf5J9jThE5NLofvhlFfJhs
AVMdNkQ8hRTBhc/X8GVe3zYGhO3iDoFLUn4BlLwnmT2JHdmQxHIAWtHoAspHBQjw1YgF0Rx9/Cw+
UEdTzcHfhQfRAyfygMS9+a+hg+BnS7H/WzghbWnEWlF0839xQc8ULbjwHHCcyiUP77R46ejVSFD2
zTWerIwWlZSAA/dZkOpvlzYLG2DMsbLlsviEZ8MlPTOItqZqsxO/8YbJ1jDeV0ikWlfUnSDkSTek
p0RqU1tJ7QQudCtXzxwaFCH8q89593EFcU1LEeZQVNdwWjPZqi3bcOhAjliCyQDRcPynG8Gzq+ZL
B7lnccywmiKJ66w+esVjzjFd5Q5VF+VG9lnLgofyC+VMQvQLu21NlNTtMKZl7GSa3U4638aLYtDD
Za6CmAqW1fjngzW+Kf38r2J6TJ1p2hjJoOpARDyXXPAYkekXPCbjTcZjiKfwXSx+rHVkNzJK2IyM
tpi4EPractvOHFUVEcv2uhae922yZIDct5vRSVlGyomL8+CeK5NnbXfwFe9WZpDaZ7OWQ7LTJsms
wDDCJPQzZlKQrt5ISFm8cl8Dm+JEVuloQ0X9nGzp03YB5KuectWfset+AQq8mqbzrtLEgglWxcb+
1eksjP2VtSaf6ZlKcn2IwuVWP34TxvtJUGO0ADznn0zIPvjXrwCGZ66MCM4vKLe7BZMEkCjcpUtd
MxIw5IE33KVROlA9bWmOQuY08EGjyE2KktjfwvsR2jvEoa0Gv4V6T6dWVqtO24OiGF5tAyeF9fK0
jcTEbVp5LBnXMzznSRcbj/FAF9ksJPLMLiXEwncgMH8KIT1EjdtGAaBAXzI/U6oa1C0BKvlZ/pgX
VFmdPC3BFe5G+dDC11PzyWF+mQuXkBNExoMM2AqBL1gyRfeZXFyQj3cGV4OLXvG3x/ga+ZMVn9bj
1P4N9Lv3cNdeiz4MC8T04N+9At972C5yTSdUjJ4oEPGu4DcbRwEnXNsRKOze5mQ8dTYOWQhD0v9F
6fhLE0yUyt5UiApBUTmj9rAaGTuyT5kon996+9XG+z7uUH+NDcKy7a1jpA8CUMwm0UZqK4zugC0I
RCmJXQASJV1c+3Vz6RJH5AV6pPyUSSPp6kj9BeUrLNZ+3+D+7q48M2BGLduX1flavdlOI3BWgECR
v0c4PJnnwuchAC8CXJErGGv4ROe4sNT/TiopfKqQRKHi0RZp/DRh7l9pq2ce/HJJDUPAHyOZso38
VQvxdLSrKGhdfDOX+gACBzzwz3X012rMEhqSDLOKS4D7HCZmpRv+fElWMhh4bSCtPQiouaKWDMu9
iIgUg4mZjR+CLfFWoxlPX8wyg9zW0e3v5ub104BT/S/1VtvVm63qmo6szROeQjDUc3PWybGTBNdp
KLhCpdhcwO9I9jMVIF28TlvY/9aSQjeRA9LlUPFbHBSnY4pAzXigslYAmcray12WK6cWQArQ0114
RAw5PaM6IkPNCFtrrqAb+39UMnhSS9UHVhk5qFrxEmPVyqZXnCvixBYyoTj7sfUtjYzp1AIhNQB8
ziOfTUjxypyjQZCfPDgL/tEhW/wpHiKZeAFKngACChTZNExIRPQCfAq5dfNMYJMzaP0qujjrFn8w
nQouJyxD6IbzniqNGphg+kbsy/k1zcH/coG1aF86tYscJ7X1kYvqs2unO2NqmTr5K1txYxn2JvsQ
4l4jEsHAxKJEWk7EdQwR3+yoR4RTLxMPB6MDAJZ5mVX8SrtoVks2h6iXwp4yKmCddLjG1zjnZq9S
gfkOvwUdzFRFcu3bvqNU4vVeAatmvUeCZFcMPYGPzZpuBJ2z9K4XcWgOV5yCZ2QdDz/OpDQqR9rQ
Uj1TWxd/ajhIftWWQYqKln043HZJC6T3ArI+dVQKHSPj+UdbOBfnFwhuFjU/I5HjdcFNCfhBTR/d
TVk3iAzy5uVVH6c4U5zQcQSnErgnJN2E0niD/RKkAAKK0RxSuF5L4m/N8IPcJKqWPUFPR2PK1QEz
A0WlECLCRppp7vLsYO9d5GwPyGrvHkAkS06Se8Ozia7NFIKQEHF0sUxYYRRO17Nb75B7M2mlmpSw
2oUa1zTzltXmTnYjzOKOQH57rguQZDV4nvqXB/oJBIDSlDEDveAby4sLTsu0gAeuGvRJDDA4pN9S
w045BhnyF1bMRI2JGiBQu1Mqqbb0Q4yw6B5jmpv1+SrEQkLNGOgnhxcTufuRLlBRNManZhOT/EFv
SzU1ZjiLFrd4y6svFUSjkR6mX/SOnpQkVq/NB6An2OBIjpd++wObXkd6T32U0p6H+IQDq7sFb/c5
b6xgTM4FLaGdd9mQSxryk96MSALgspKvulF5uyB2GtvfZtRUAEMIGuQMuvbUR8NkIpxMKhfrRl6Y
nHf8Q0GD+1ItJUbUlOC7PNK5f4oyqQAnng2+czrb/viw0xXwFHcG3xOG71HelNCGqtwXcVGUOASE
Uo5MAn+MiMEEshO5X3gDp5Xa8tU8wPDLISKwaDvL7RNWWNtNx3Y5q11EdbHsXtBqZVvUnDuIyF0o
KqS3+YZ8jrbSLmmOurGddFGjXoWa4RGD4rlkK5/6QVByCvotfaJ3uqm43lOaIY+Q11Angh46qCQP
B6lqnIqSLx+t92xoxVKf/xGXTpC9paxMzhhJ+p2cfPbX6MqZD3DjMH1ehRLst3e9bAbZVoqFzAT7
OFpt5hoLIkNIXTWUNtGBWHlY0sbY+nByU2kIA0yOsFhPJIlxWbArsGwo8hlgu6DwEf44Oq9BdF7a
EZdugRllovhzHsxHtdpQC1gcNR7DWp+Zthm3IxlEkUU/e2AzbLG5DNeD105i/Hw2CI+Q4TXHgAPr
dAPRQwQ97S3FDMSncYra+gjEXz68iVIJ6uu6rNLAfIt702+TNxPIYLWUovB1UxlWBFOwWu4oWfnL
INaeGi43sagK9zWISJ9ocPtqhwVdj5bnbNlXEOKTly1fjxEdBWGSketgmxKHxoOBeS0aog+lTjKW
0hEQ+XpmCX1RbyfmvjFtwFZXRtGsNHlLChPFR3TfiDjJxG/Wo5DCijvP7eh/pMMc+/NSRSlmwa4O
qYJS2ygBcfKkqp5H+8BntKsUvbUlSWtu9j/g1GuvuuqO4ElHDaCCm7MgVPMUyA3zVYTSH9O+Fr26
3JxgzxE6/oKOv52KnJS/eJ2VVk3aytOkzFzAsndGeyojMnbXA/KVEItiUrtLZB59O3o9fE7t1UUC
z41pl+CwDyUls30anCAxpwfvGN1XuQHUv59OHNwiYMf0Rhlw4r66J5NDYZGqwFALwNUtR5TcQZwX
fsrUSM0AxB7gI1BVtShKNnz3/y47VMyu4WdU7Dp/au2xBLL9iZh/WiV25Pb1zMFErSY8xztJHDf7
6z2Mcw19nWLXhi1dRqNAdyUcuoj9e/7D8S6bZxv2e9rss/tNDpJvQIeenKJVTeqSZpzPfQyISsxG
4vTqE32nmEvlkV+wnnrDLknRdx+r9DxESQ0Tx0kQLaR2vLMf86BUYriUut4sg5SDKSAnQ9ixN8ar
FOuIUxdQLyWMlSAeLMBkaCrU8A4psAiXYlZVAj/QKCtcadXqSWKeapv4Rxes9J2yJ0gApYqFwfDF
bUQzijG8agtdA4Bgdkl5f8sNWroDIS9wKpGDO2scVvzjNsJQ3vKGsag8Rn2F3ZCfJE6+xHfuK5Ia
vglBorgtUqghfaLzs/kO5qC3GtqhhB78WB2+l13eIhP51fgiOIhLI8kKK5lwSRyRYz6GmWXROZt4
O//vQ8J+EjMxNJKSL+pjux67jQXHgVtKOUYk4ygNDTFKFiP7jh2/KkMNknagm/5BwcklGMyWQ1eD
q/GaVE14ACDrhNNRPneUBJ8MGiqsrHRIL+K82hkiUuX+HFGV0mgrv/9+ZbxuPaWxhueKfX2YlpiT
8Q7Ezzuk9xpapG3SsZ+tioXIsKgZQnvnyWPJcpVtAwn/sGi7JdrIQpdWWk/IWhVDWicfwlsHbtNb
uZ1SYrFPH+7v/hlyQUJQnZmPrNbubiVjK9ofzPB40dBHQ+RS1js8GdGpzDLDiiQsjISjEi+sAXdm
EmKR6W6iq9Vt1V7EgZ0MF38sF1W3jdNg/XfwM58tUc/lVpGDRoNGpN53nxZo88Q5a3mI7r+RSCwi
dmanRFtP4Z02xPkOQNSnGvNX1rqP+wHZY2Ch1QI+txoeciiQgwco6o7ZfKmacRqC86TOcOmtiXUa
gC/4bDLxtealeCOUplYhU32FR0CnlKbcyOzCxLqPSFum2hqIPylIH395rgNfFrAYFwPWtD3g+YnO
Wwq9TVIS1UoJntVojc61P1/tXHfjMiK37C6FjJdw7+3B8vHTYTIst1CsZbtN/o4ucpYux9xD17FW
tdntNARXXeCvElZsFyZOVPjFdlhRP7hqotCfNbViIn1eXP5/LSAPcPClMhFBMue9wGUoV4Qk4KAb
PLxUhmdS8cMDIiGPrlT4UcKCmlmwQvmRs14cOEDCxfcMc2jEL3Ko1/UsstLVQOmphdYbohpSmGso
2qpnMGQ0GE3MHbz4bRxXEF/lGPzQ4SnwYYgRkTKlC81izda2tP4dHT/jXPGYaGeSh1L6wsNrdreP
9kz7f4a5dMqh126ynVXELkp6d5UaljTzSNFcJaO04kkMfExJaAIRqiwVisPgTRMP2bWwJXXYY5w+
PcjKFJWroTEjZgH7cRE9X+1AT5QDC1wOWlyqrmeHoT6s/jR6Im+2kvWGyAEKGe4nu1tA4fZkdgX9
spVlK5Tw+TaiXCJs/4YurZyZMHGQ6oOPmaQNJw1uh4SuWhv6+KUjpoSgHPCd8WHcp0oemmDc9PAX
1ujtMXHOLa0DzOuhYbl8nKoCTWC7jp2unNfqv5vdfVoeXtcuLg6UU9QU89bW20rZ/n0hzoy7iSVJ
fqYu9zMyvbdXZifaMOvoaGh5qg==
`protect end_protected

