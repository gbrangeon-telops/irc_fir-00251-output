

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WrSZEf64fUAl1kVl9HWWVm9JOgHMmzn0fv0uusEaRSoZ0YHKAX+sj6D4gL2WXWrV9+rdMofvPwNs
9A6zs8psHA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R/iTmfCVAo0uuZTRynJ9b5Z2gujQ7+Xxv1u+96JME6mwR6F6/MPV4ayotodCx+xcD+9l4Ktib8Ml
C05jFwQ5vFi+09RjQvyvxQAR5CtE87QE5Bg2A3Gt5QmE+m7ZfJiQZgi5YQHL3kAHS0jfaofTkZIU
6VFVSW/fcrod0Swq7VE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RAfB7dvLyt2uCWNWspMeHiLYPG4TlOk+8Dptz+NhWH6nMzYrNkf7IWIjXk3hEVf7lwT/X64pynoh
QoCCtl9AW1iC77VMTIu5MgFRizuZMUfXZ0crSPULV2aGonx9nQ5JKx8TiRv5BTWxeAsuh1lT/5p6
2v08ZCt1Nwa8GPmEeFnTZsTB1B0jFzZQMa3GGdV0nEcSjDo4bLIkw9sMEBW2OdUuvE5yIHF6Z7++
/wzulmNKOqQpmeHrq3r1VKkMUHNzsDpLkGo5HMiTmEUJr/s3uq2EhCIq1agWSVbcEjS5uDaYcwdG
D4cRvgOxtT5sxpWA4fivRX7vvCyun+C2e4pYew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MsyF52v9pEo5RpJJtfhlgAJQ/9a172C6pJMP5S/aXQMuRuv2+JV5wCeynUZSXHj38Ger421EXuQd
EmO2OIKWiz2pShaEh/NwF+InGDF0QzD16vAgn24LAOYAOX1lcCquf4w2rs7e+0dn2PO/GYRn4rxl
E65F1qdRiZlUeVoRHdk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
klspBE6zapxwDIEksFW+V3vEj3afpsQxyK1CWGpsw53FDriMhZB4hONIr9yRSN9nitmQ+6cnlGM3
S4Cxnkb334zdXXX5YoppEYaAdCcB5nDsYhSpn4PyPhd2ANmiSIXxEjiEJ9MDJlVIobzrtkNgFEWA
QkqC/Eky3QLBOqPuDJIgkf5UFynGEkI3eWzGSyuNAHTTYXfoLlYBh8nelaKS5vgYh7jpllyo5l6k
hn08k3sWZKuN1S8dwb88eFGM6hwg1UoX7pTnUY5yGPZZS0JEiN6WVWRmh72r5l3yyFZOFNcvByJJ
z349Odlh9AHKI6joGGP9sLtbKDrZfmu9y/SSsA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22384)
`protect data_block
cepYRadAPzkI/8n7Nysww3jPhpA91K1FTHRtBwYjy1qqh+aFj14G+FBYLZb9VesUnx7DtfHsupXo
SwmzoLahGbn7ftffWs+iqtauAN1mGoyuqbbeJ9lCtk6waqVc+q0eS+rLieCEZzXEk2v0Lu3KTEBK
KOZmlfEhZRWrggAG5q/WrgUyBof2BIdthkvLFYB7wXlEZeDgd0ObLwQU5/zQsj3z/ya1VtGFG4LI
ZWpHzwkC6CfX/CzTt8S9t+5U23hKOvEzaPGpVe0Cobzb5ducPeCXbxe+3hOn7D8R/mcGPHzfk6p+
X+AI/He72CwegkPvJtXOMl3cmYra5kwfT7i6fIuwkNT3Ra1ULHRz6eopgq2V2JRKEqNvXwsXH588
rHGIJ9zw+NHFyLjdPUfQ8xaMxZAql6/Nw91xKtzt8Rzd7JheKVhJj24/FG8MSMWMJOxq5OAv9P9E
P6EpWIYN8MlNRr5YZQyDeFcSk7/G5y8k+wqjSWxhQmc2Dw+VG3ogSkLGAQSsWs6s8E3fa0QaXt4Z
PCr/biCxqfLY1spwzCkbmA9nsyyju1IMNxUpCNFFCo923XnJ+YYxKkViSN3OvF1gGvMiZqp/9wLX
zXdbzh9tEhLfWcD0Hf5C23XOR3uH0GoOpzzsqoqKP1LdOZ1Qx4Qm4Aqs6qJbhX1fOrHaZ5clePgI
uJZqMKhVoNo5z0Thbki5ZSi+MHpBYagjgxAlhmBBdKai2HV743ht72GgrJptGaNScBZDdlvR0pDR
E/T9ueZEhWWOdbx+5xhcGha90kkA5QowUjpECQuPypi9QN3u1N5GQQ6n9zZAhh2vTaTWlQM80/yu
yTPpISW1gAkENlD+7BHaT3LvfZN7iG/8mvTexQkPNypMdIzjHEu6rEAFecx0ZRydBLi8bXjQRmZl
K8om+KxGzmwdb0FxTMNGHoLgRF4EvhciyzBLgaZF3V1bKILGDk4y3RsH1sylgaLf4goluzrD+BbQ
24xmx6DMsLXxvK7FS/YCwy1BwU4I+p0uHPhWEAvFcDWmb/jnNhqvLFRZCjT51MbIHzJWVzxbJ0Zl
lF/nOrW6KlVoWo6tUUYpJcPaBNbo4Gb7ourLTrrsnsBiVUBn4LoDnlA70Ew7ywXuZoeCOwGKX5xe
6EayTPn7xkcwrV3KC3Mo01FQ+3exFoDlC+I5WUxJDTnvlbC35/DqKZc/RPr0+tGiNxxtQMCWi9D+
Esnhb0FczJCT07y+VsnD+OeaZlO5M1aahxk7VZvGkQ6OEv8dzftntQiX2bYolvtYMSVoEylja83A
jo5oHoXlTlovCrXmY9jq4ZVY4QiWlCIyMwVbqorUhhbliJySVnTKdVVzGwsOXHIEaEYkG7WN/MaS
dzVfD5DrydDqpXAOdwXO0Y1XhcJL32/FoSYMxJ8zbQCINpUriF7T6mZ7S5rqLCJwji6BoEtgGhSk
hVSujNFIc9SJVMl29O2Uxn5YRHpme9h29FLQI81RNhUddUGxKtdDGJs5Pa++k2d147LQHpeR5zOH
Tq+BQZaeW8VxzP7kRu6NaeXyyO4fs63fV/+unjb+gkyrguLZO3E0zko6EmundmgipXji5+qrgFI+
Hp90D/BdXmwDJelaBX638/722ckofE6euUM1JxG2xnLJr1jUKzgx8mMbaOkf4tbaxRVyA82qs3Zv
JX923vB7QyfT7VQX/yICiWoVWZQI0xDgJkNkKZwGT8091gSUrn8Qew8QheMkbKuJD7ImGMYcWceO
17RdCnI7iIe48JkBn06NKqf8OfmCaYrsqAUkw0UH97ECGWMo3mqfgutsyHFrUL/fJmf+X65S+8VV
t8pt5Gju/MiKTuKVR7iEaoI2r+Hbm7opn+pmNZ1mbOMH5/ML0BHzTw7tz+1C0aeqIOA+7DIIPBVx
LevaUkWmJsaagP6eBsdzdDYGFLM/Z3Rh9xO1lgG+XDRgxaNjGdrfMCj/OjumZ7NV3PdgrbYk813q
Wt/rsbnsGeWRdRsY5Izbq5TSdBAuVmZAE/IaaIpEzBCKmigF19iHsI6LQ3ZLUh7w99gDkxTcWmyD
MtEoQe9DiEVLghDmcFPIob4JKdWYZKSvKmA+bK2EQSZF9e8HFEHeDDA+DuMSAaxR0vDz3s1DTCks
3WkSX8CT0lZr14F1j744XWReop1qfs8hhnw0crQwPMqwozv2fUlhloLlTYaSLEQciE+8Sivb2wvW
HLtr4AtpwPOK7ZyCNyFyff4QLFJLKQVwsJPVJNBYEqx2M+WMO8J4DoyK6XG0n4vS5U9G5eVidciL
uwi/hluDzea2B5EdavkFzFL72ZvbYLxwEpN8JKMMCFejdIGpkDw/crxQq2ICA3UsblGMAtxeSzjz
RMjpwWzFD0et2p8LhMRAS1C6cuqpAe/0uYNXWjlL/bvN59ojGfUB637EDMuZ4idpQHdsrC5bQRup
F0IzjcsF0/DKPEaF+w674xLPtAJhYabpqfYp4aPWm8RE479xxtGOY3fzBf49ya+WjhIDT57UJpPN
skc3/KwdEvzI+/dUsZ5CePktsod04PIFws4y64vA2Xocg2fvAiHSswTGvxa6J6Vw5BoDXf//ot+P
D2A5+JG4fNcpwDn97FCVL7uuK0EXalVsrekq0oJ/XyHsmDjvj2bHnzGMTsFNSJhtrqEg35RpUhvS
sp1GMTxVm3e1Z1mokeZBOi3OOLQvOcAomhQiXJsfZmY42Pk6qp3YGZ2uT22BaWJST1eK9jtdsYdw
j/bOb54h01CqYeHRCi1AidVgXb2vP2e7obZGAZSeJAnbhRNHmYoazie7eiAFqdrhZuHM5uQ0MpAv
sOKfY326hjVpvOF2DSKR46h2Cv6IylOWCX09qqErjhsDl4qZqfAFD2XTCyGaV+k3pFpOG779tN8x
R4vTVKsL/bfN2/DX7grP1XmSBoQFlwopaFcwdwga4Q4GsktqFV+rNNwmqWGIU10C5/dKQKE55FU/
6wCxs+hBJT3CIwWy0XCfj3F3Fi5gHwIWvgJH8JE3ibKxbaXoBbYZMIIxgMvgHp4jJWgo1F/46zeH
rlMDYCwFK6r+XusHKJcA45fAj33Du1nxAUUCyVsRNBWLc7U2rUwe97cQjRT1n4RLYojp84vAQfov
0VnB1I4Oy4RHKIBprM3XAR5OVz4KewYO+JzVPB9uxmg4nYAn5/e0hdTHMTPvVzo1EvgTAwmq8qCa
st5VHRGa0TVUErHgyrji7dQEF/30pt9fuP03204amtPzfLcdeCmPO/DoDirXxMH9bNjMLot/jfJu
6jNOaKTrzQTTVvgcYtIx4LoWAPYyt6YmpZWfqVrcqfGPIMFpwJ4Isqilx7ae+V2xELslo5a/QNYC
tkhjALSZlFyp9MEnMFJ7bHtj8HJo7iUaBz9sf6oc8aVs/8kmB6AQEEEVYz6GbQWgpDtKziF80Kgx
yBdTP9zoFq4yM7UqfptYr1lXyIFgLfNudf6q887/xV0pFPhhEBq8Toa9dO2naXGNmABHHzaAM1iL
TErSCDlYtqBz/cfujU5Wovy3frQDhO0bc1z3UQoRjUMmDll42lyn09gH0ayXzePyWIFKO03rmbxM
BX1UbWY7dkVv3JuqPtAY1o05485ivV34R1cI6ZBkqjelxhfcz1fbIY+6w3IUjmHiG6HzsSxl1xYx
NKgjO28gnfsmOVCKK0Rg5neWuYUmmiD9jmIJM5A4EfUzohpSs1HHbqNEY3GMqHVweJITllfqZtfU
YBR+E4LbkuXzkMFTTuGxQ7Jv879vvwy3vkC7fU5E/4kLiL3tTn1only0Ju5x/PvOo+vgYWJaDgOC
1FSBTsXkcX06rmP40ffeAMFJmem9QNhZelrbxQfnu84iLkC8r5t67EFYAZuo+gRL5gQUXoFT2kXl
MDB92Zj6qYLe7kJxccAymxM/6KhQR378PG+KCBBsm4f4072Kv8GZWCwnPCyePfW9jlf8GnOqG/cy
+TkUH78pzH7lbDdtUhpsZbKH7U6uXWZa7NGd6wqpg/rV7BiYfF8XbceoKYrFhqRcL2v51PCMGSS2
9ZmjU3w8q9r/ZjPVaMXktSVWLKkRtBXuXdI/VSYJsz8SPZQKIVBUKm/F7OVccor4+5q6hhb6XVKH
ysoQSCP44uAgVe7cayw0murswMMfhLZwVXmINz6/x3Gyho+1BC0T8wNaGmR7oav+6t6SfgqVa0Ml
DmkmWE6nocuz3TRwYTX5/SmcTRAG6XtwdxRUula/xRklB+SakDASGCCWNVO+IXsF7w5xZvquXCSm
3f7Y7HYs2yCc4V0g/+3tXpv3pRmIxXLXDktQrz+hzh+bIYrzhhOKu6S8xdlASyLx/rLhPvkEc97b
cypVJI130lkTeiiKETxqe75p8sm8kd98vxxBHHsWUQvfvVqfMSagZtPODgpdDLjqn09Z9FIqjwsA
hLDcFJICEzMmettXvByLmBPdoStK+tSjDFDqykOp5D/yBsnj2lBmWT1axivLyX1qGz3isw+8L8oA
5x7Z+n5vJhhwa2u/CO0wuvrLxitlrm7V/FNAz8S6XWQHNPzrZHQCUtG0LrKWS4S6jX9Zo+wsVecu
mida73MnP7R3ezOZ14fpJ3uij22rXp3zHvlah1sYkzMgkpasncWAfdPdE+bO5XZqukTsh6bTFRZY
HDZtpD1YfMwe/2SgF4roCYntU4+M3iOwLTthii7x16XqmGmOX39vil2b16XKwK28pQdOC/4UXxSs
E4itCSraBHlyXcJXekXNtmvK17Mhj3hAbFfGNEpFjIm0lH6iKXerRh7NE2jH0qg30EnJzAuLkIoJ
b8PSV7HzGRsnxCGwrKhttTqXhquPv8HmVzReJbqUkmSR0plC0lHPd3jJh6XsKM3SXMRYhbHsZh7/
HwhJD9pjO7uRn5OqP7YcVbsDBeSzc3w4Z6p4FSVJBv0XB6+aB67ukA0ldwq6VcgV/tWqNFuBNdxE
b1qviSiU8Ru46QPmjfwdVZuenJd81tTGXB8gM3gwc3vX2snertfITML2ZL3LzdR/9iiwdqz6sjVx
R7XxxvieyHYsnOOKvOOIWCKLWZZmvJmJ9QmA3bN0j4uZCznO4FO7AbdaPrU++/KVVcaYYTn1yvZX
dc5kWiKp0xfWe+WIWwcdasevWAMbJ4CosmVd+XT+3rUMCK9LFrDKLLPv1iuMPbu83qp1O1p4YN3n
VhUKJGk77MkWdSan2ubXXSZYg1kImvh5AztqCr5MqqulwgBYSJ6pGrRBWft6v0D7z6oHDs9yk1uX
3wkjnUQIa/ygF6kkuEtFnVN52x8o8m3SY95va8LdPxTc5PfVgu4nKGvsN5RBWvDaIe2VBswh+9wU
Rxu6kUkOBPlDKPDLwMPSwwriV+pQOkSOVAb56US8XBecEwkEKUug1WVJncK2/Z91iNT4pXfTQXID
cJSk4ocmSQ9Sh6vn2ipxd5Po2rwlXGOKUp9jTDt9S0W3unHfRpoWji78SqIlFbYVDDDjXbzsQeA1
QZJ33InidcfhEFUkP1PhEGkqO7QYt7QoROr/bryLUwcPm1aBbbSeFPeV/tKes7UdDgAAJjfjXsCE
as5o8u76UlPkc7I55u1yp/yYacrlrcOGRbdsjX1K6UiKnqMnSAbAANCpAx6ek20y4PC4RWax3o41
dLUXjQXUe045Et+oZf4lHt+vruNwp9olvr3xW710JPV9o8dWyz6C+ZUiuWUeI9qK/Qpt4XVXEXIK
kEdB0zlPG5HNwO7azM73QqRychisNNXuebpEcegpPWiogg1KJc4hfyzOYATbutzGtZ6J8nvdvU+Q
0JXKBcFzbmCGB/e6eclJ1l2vnVpecmBFQpChJkEonaZcBCVbcIoOS9Hu+ak+EjEch+/7f231TXjL
mqY3QxdFghLKU6ZXXzCPAQdvOsaDHzoAvFXWdWizElOmJH6STFlEQUwBQStfCL9tLtxAxKGzfpcl
OaDCqbm3nTik1MUkx1xlKUePnUham+LzfGtxfmjmLmOtCIYr4N7ldLIC88z3CN9DYJvIJRM8HGAN
vpZAP5zQnxwcgXaKuzUCT+/ae8MCbZmkoKUuWY9TVmxNRR6t1Ic5QJYeUz3BjI5v2k+NdeYVEF52
F3db0eq8NvLMMeUvfg+6t7DX+3RnaO9eCbq4UQn8O2WT27apS7pa5FXpCWnwf2NEiCIhAdbLHbfO
wA9kA4WV8gc7jE/J0nhiUnwQjmFzCcZejq32aItR0hCJnaY91JPph7ynppXKjlmOaUIudAubix/G
cAZtCESLBgqm9G83w4mf67nuBWRa1w794QKJpUp+s7zvS8Q2YT37TqYt1ymsqtokazpKX/5Zw59m
gqM6tncyYJuGAukLvJ9kE9856aluzAJxfegtN4OPEijaC5hE+QhaodrNihtYGhbeGU40WuyfeD1X
8dVySzcATIEXWUFPVvicRXB3hkBuWVl433dYrQG3XFLYvTLTmUCcew6bQWHib0S0CrfqnqEyG3RZ
teUhQRAWeLdo+NHhv12Tibj1+POG9H0Ixno3na6u+x0BFYb/kN+f+dwKvCUh6C3YWFS44+OFL7pr
MFuAdd4v1nO8TpiuMzx/OTFEyEJyPXAIk4a9oUEXqTuP9u6RprOPPtC/UKK3i47KqHsd6TxvNBY5
QyTd2c6FgX3X/qyuh9yuRhDjnnn8SuUJg2/g4ALOKI7OGnVXQ3zPgWLMnJYrTZNAl9NfOJwDhQk0
/LmXzjTYCjmviaCB+15ufYvjP+sdIvisdx/uVDf3dAJzWX+z9wN0qv0PcG9gUyOZai3ZfX25Tlnq
DH0MinaBAzHvXJ6X0F9eWuWy6gJWPAC8LGTnkbKp9tE/KJx31KT7bswUA0+rrUwD+yrbCxsfH0Dc
jh91q3tJ6DU80qOK17HhKR6E7jIkPBy7XmDCS6CZXyT4+6zf5l1W5zXo0sg+hJ1Tn6TmLuOaFoLm
j624nW4rVVwRWcsVBwJXHZfROwdcTWbOuC+E6UKJc4ORyYo0bp87ByxKvmX1eqDtPPiVKNPKBZxJ
mnP3uzZaNVGw7btapuojZxzOQ7/pUURjRqumiVPUvddaIloWV7AvvcrdLegJ89pH0K7NP8LkPRIO
6D4BaZuUM5qLpH+MdF7uYPx6PbbP+gYzmq2NAgJX+YHqpmndwY1g0PpFCuGRcKIiqlaMPIuLUvCZ
MyA6K7vIievgUhuSEKnZGy7X4AQCUXqF86ad2JIGYWmKVW4kDI34tk2F39QVQ3BTsgV0e3/OTZv5
WneZnMmNy9Sj08E0prdKmf2YjNU+C8AdOIOwEnTetgZ2MUjBod4zL6tmRXJoCmmgIqnsIa9uno7R
/gX2HVaYtWVKpP2nZNtlUlCp50r7dkigajOqrDsUp8fN6xCHdwVrpEYlPMzG5jzF/EK6vlHkRWu2
UDjLiIxYl3OSDMFa8RePOXjP8eAv7xLAP3+7ynmOiffLyYyCxr4z+NUZqktoXWBwAS29LhWkyjBS
Fjri2xRMs9Fwvgm4SPr5Cux1fbNET1P5x2pFodJb3Xogdbs8xAcvtMr8hk4U+P7Rd56HDVjHQkLr
oKkBuXfGxoFOqJ8TJYZziw0/HL1/QqRTCjHN8WpZClWju3tuUbp1XjtLVMcBtXYNyqoba3K3lhhi
MibpQnxsyE5zn2JEa/VVtNlPGzdkNInYQCa+q3skJvweNZtxaA3CDy0KV1y87Bq4qLiuJztpKHAf
lHpiBpU7WyWAsaTUjH/DJ5iySWnfAj79ddsIYToi/MDlDmOQeJ102k/2jTAls1XtdbV6zaJVixhO
veGbt+NjizWvDlWir86Bm4t5mX/UC+T6qqfDaWGU/MgP3B68iVvzRxw5669v+a91jX7pDosIa+Cf
xlGM3KeQpBFEfpDdr3yJtNduHPgSiwtiIiN0M+tLL6EWBegG2UeeK9GwobTDFPbCPntHnqzc/MW4
ruKAf4dgIJccypSer6Q67IgIkpTDFxO0f6mHjBq18E3ZRKy7IEPESdMeRjQxGzVIU7KdNLA9obLW
0bof06WjNqoP2pUaKRx+zcCRj2o8UEYaZH4Y1hLCZgC92gEJvhMKMVHoIEQ6I3kn4mQEKTcI2avg
kzxG0XE8EeRD1iPH/Tfy/GW1AwQAztswWwbbEuCnFQo9IW10t2vakj8nwrXpv1UhMMsUDCwmC2Hb
h0RN/FVHVjt4Ornx7fbM2cEZJk3c68Z0Kwda1xk5f6kZpnfS7Gwe/2xq9U3qj/TgvmxpS9eo9SAw
2GsDEsN8a2rzv/U1fT3rUbmC5d3UNPHrBMy9t5SmXG9H+5bRqv8eZCWvx2LgDUivbLQftWfBCpq5
jyjtcUNSAISFMPh+YEGu4PcMz6ireI3k8M5ZOokXAYZcre/doptHX7GCVWGdX7wrWTf0wROjPvou
mNU200dJzmQERi09eu02Ke5ci/N3wuM08ScyX5VhftpJU0fl1bT0bIwQ+/j3EYOVUgG3RZhvPF2f
Y6BV907m/sO/Xx/oZRJzWXI14S2p2s6UxOEriT8VnLpIu6v7WaQCBoVGdn0C/mQrvZYHMhoZatbF
zf9pxdU2xx/dpv2B7VH08kHghZtryl5WRBuKLmvr5Z2c8HPc6Zp40UyBXPNUEH2VPCd6bk9Vlzbc
gZQGInXIBXfPxwtaDXypB9SBBcS1Twe1qOtgsA1t4c0KsjxDzhV2m6X/Qt8/9yLg35bgXbK7chF5
uDEL+NtWNqDvahkWrIs7qef4iGYocBhCOlx3KN6PpB0VGB0siFvTcqW27vzaz6hBpMYNPCWFc3xt
xph8BI/oWxgzh+1flCTKhLDJhedpfcfzJ8cC2ezxcLPqNZ1+v+rQuz9x2x/2iv1JZP79NkrT5yi4
brCmMEUIqrhxGnyTOFqXkBMDHedQw3b0FjLzfvDrZUnyG2s+mnrgFiQCkX/k5yJ79NQa+bMO9Ra2
DzweXpVAwNZvn3sxNodCH/qFi5p8e5WJwO2ymzXGmsWkYCmAH1Xm71l/nhecXAqBVIOPJE6XuF8E
OsvhHFBC7z8Q70SRNMfvI2EsBpEZJaqi+YIzmOWnCdtz0XbmkoWaoTTO6in6TqwvmmsNUS7T9y7B
y0agnDZR8UB6xcZdPVGoyeFwAOjtcnkIC3trdJ46mqbYRbXOLi7SMUXLIJJUzYq17dFktNYXePfw
G88WKkI0gWWpqbz/Oy7qLJti+edHZg14mHmVCUq1dEBiD6ZJ+byBTTslixE0HSqKXWY3eKkzarlB
RFr1bBH6nN0IFtI4HIF//Ah3Q9TyC1GNg4SBNU63WKVMwZq78Sd2iEDCxDz9wGqnif5H26FKtE5N
I9nqWxvrMTMdRX0NtXoO+ps3HH5cFp7IZFh3uqujkgnooChgosQrQm9xJNlMG5cMb7D0uIbIIL8G
KIHtcu6V3YAg1ZVbFMY9zynGJn/4Bq6eGFwRGu5QWdkeoONalDUgwhlFmG3Lp2gep/hghV/z+4ge
2Cvvn1F0iXPifeip/uGzWYSE6Poc034XRMx+W5O1Amzu2Yf5HKd32AbX/2iDiB6N4xuxMe5vpS8H
D5NieZSyedIS/H1IwovhHtJf8513YfoaDCLiiXl0PI37vyhMgZYXZGZINWez04l0vFLFYhWI5LLX
RYvLR+QxELeVjutE1fzFvKp56YLJQgvE9z9VqDeRsG+eVX8Y5MvSN+EyVK+eqYnQHHOHT+qMadpF
L7Cp5WrSYR5f4sgoY9fCBBvjIbbeVhhBoxtcDBkExAy2x2SNfE/xtXkdqBLrJmJL2zY5D++xPyDY
Fy1ZX+iyVTlOW2bqfuwcD3PYwSA+GX4xYzknMUmpMuMaj2COj8cgPccfyMLI4rEQAyFhuxW21u3B
+FJvlHHac4tKklbKNxXbTfKB7ZsyWRzHuUfnn1YSSmUPpfQQ1UTuALrIduK5Ch0T3FwBH9NmX0pn
etlHcdy9UtrVWY9X7Peo/lb5/fNE0ejJDZKF042A5t3X7Itnr6QsRf2wnFvA5gpqJtqm2wJcsyc3
XHLkf6O3BaaTO0+ApHU9xv2P0//uywyOltA0AZOfmStkvwyL+xDm+/jfp49iBCyKrdzX4fYM7xAR
Yp0L28hHQus7jClP9kBV4OM90ASaAqgovKvOF1/KSNtyh9E6bxRUox5Tp+WQTVYJJEubzGBwBwRP
psTAENLtJBJMrtUyIoxiBFrvVLysHk4CsFAiu5XU7aDv5DGZag25t8TZG11J6bfUzpBDKJawmy7U
b6mDaPrm99N6vbEbeFvMrTKxKopiYBR/IQzSXUTTdWOQj9+jgGBGOb36tOd2SSv8rvS/EekEVzwQ
n0TIywT/Q9z/OhdWkHwCNp3LzwmsMwLYtqPFqaRWBbKkeXzcTL8Jk5MLMYQVmf8ubaa8wGnX1aFA
VO0UT3pPYlEyjt/zOJfQ0SMBeRmNFsWD0+jBDbgdAX167JmAgQmOhBoUraxXTMfnyIcVfmeH0tIP
SJ8QyVqGQg1eR2q+3XLEf+8klq0X4g1N0prG775daQ5cHXG00Scw3Ci5rbr/5apovDTtpbi2szvR
Vkj48vtRP0i8X+CtqJBsp0dYcgc05G4qk3drvvUc9lNzI3U437j2uBeJorsGZoWaf/CGlXvbxD4J
LKSYU5wnD6gqQkTu0iFBFNWYffphqe1WHJFusBteALrYi2ZDedxvZRrHyHpW55lV32xjXhbxbdLL
Qev3jHcVs2xmbIiuPrFWyjKEyf5KJOcBYOc4g6VXLOAkNx/chdljGv2qQaOf9fNsSFOFxsJXJ9j5
xE84QsNZDYC8ct0eHJUTzkEE2YHI2+SD9Gfoyew3n+TxiW2inr4JxThNggID6+hbiY6wcSsswlVt
T4Zea7KY3YxZM03eZqGfdTOxdwJeZ2qfWPySpXb0rhgDxXYZxkk6LyBl/8TBBCajerwoHL+Orhcl
zuxGaGGqagTAuNobtOgF54f4NVlub0KvlYFXqKubET5ScgqvFGSpYFjBA7egJd2pnbV/3TiwVBV/
cv8E5IfxqEf9CsI6lLCsbtmapU/mE4MLCnXfK7OVEMJw55yWxsmyGChnMbuvl9tQKj3jcAzPpK/d
bywJCpJ53qwrnIepvmHs2wGYxft/u1jYKMsxEQXjrFHMcubEiAF8lxCnheVgF7LSao0Ur9P0uTMh
TnXKwy2e0Ja72HLbPlPraNNdmzat1oEWQ6Nny9o6BZclJU+FJLB2KAAI0M0m5q5m3E8PTNSfCTpZ
lKmjYBILrAXxZEJ5Q9mGXhAEvqfflLDp2PgTmB+xw7oSneDp6m4XvsAG2FzH0+kaYZ4RvxSxUj2W
v5kkkXtL7ucb+042q6vsxEJ1mVL5pGq5XQeflyhswspYQtXW0q2sF+pUM0qI2WYc/LXv0AR5upKi
ivr8JcNVpzHlHVErCydEkp6gYptZleBgknjYncLHznzcAXt1J3wcOiXXQJHnpxG3pbs2zsf39iAn
L14SHUGJMLJEMb4o27w+W608XdWk0KmkdMQw8bRM6DjX/PfU68EfmHZ/sNiQp+1EG2iRQIJZXpqY
LqJOrWYxdJqim63y4gdV3ltEL16CObqT78Bt0jA6b4kB61O0a4WW7jXYAynFp/EforQBXpsIzHGc
8CWlnu0I06HadvkaNXwPa2hybc2V5ZemM8CnKojgQDZTezzIeWMKJPmPFmupa8CJHbtT3fK/HBSo
/SLcLqdwkrr8xX/XU6yzTQVrXragpnZ0D14DFaecy4DugEdPKAKVyLAnAwNu1QNay/088bJFVIIf
C2DXDDcD5AzH//q1V/ByRjRk4xA5mz5xDGFMhu4Sd0E48VZ71JTvW/f0HzALqqevKhRxgTeJ/ZrL
TAGvOrysvPlYy7aP8g5WK7M5hSNV3617pkIJokVRk+5p7Nd0shObfQxNxlIL0XWe8dGmDlQmXi+O
4xlOViydpFmGio/hiawZicT/Z8DAPyVdA+0Ng99clNXKiHD9JGS9LWqaoZvHAUQfB19UL2kbcvM4
Pkb+iO3JpYwcfYfWfs39fQfneNmZ8V9KN/4IuHwkMjqR4Soz9Teo1j2zzeGfpB+u9YrvO7QwD1VR
CuzDEd/gamtByykJGhyeJM7KAmgr9klMHvu1K0pogDI+2ECC6XkWHinjbUnojpLPvmiD9AE3gA4E
SjTd/YOSVqq568bIQUS3wAWIv9m2yxOCaM/jQiZ3WeT0exNxowVKMhDo1gxqQ1fz5oO2oft14fwT
EJf5I7qqv2DfLQczPu2EZdmYZI+yvFgBAHc0kIMrG2z3qA4SrsIxfMh/t7qdpk1uT6vHlGaD6/Ug
/TZqOhQdoc2KP5VMmxFh3LDPx0FheycqKx2dZE9VKXdeyFolJAvekwoFnpq9bcZqWTJ+GpEI+LvB
vKKZsOdINoEKWvc1flqOJs2VJSWkMZG/9bgdbM1MT54iGSc3eIbAm+YGTDu1IkHvlO4BUi1kGP+d
/hmrNkEbS/POrtEanHLpdFghO7CX/1+iE8W2GkjA/ne6XUca1ZsDew6EKWIin7ZxRdCBJoxT5o6k
M+6YZjskKbPYn1dHnE15FaQllJI/tDOH/EBXZkWMLjDjEIrJpDjx5W0SOhKxFZ/xsIgNwxySNACI
1AnlX7TQwr2H+VLuumDYo+ZfpZBtZPkdsigdgbOO/lyAYD8p5b3CTszD16z/EALyhzIq44j/k+n7
CAHOJv/kvXsnYdiKWmYwTMHEG26T8ZcJrT5xtWnwYoZMqrxYex3HI3J9UEgWBmUpIlGVfblEskRC
JYGSZ/n1/3RA+6XAcKxRuSpjumNrlAqmtjHRWMfApGfv2l2ZVdSUqi9cJmdf/VyquCtXIbRBt80x
lgFYVfxsIllFwxV7dULGN05aIZZFB8oeNffux/2X6/gvZ6jIZktsCbXzSLnOBOgdccOoCd74jbX0
Sfk1UN+Zvd4a5jVspNmdSZ+WulRKUbb7VCA5INtQ0w9CVBeSHyrY+YzrkLQ+9Q17WrLsiX9w1mDI
3L2t+JIFfZqYsbJZsf9XlheuMxV2f9QKzQ33ijTxrYiPtn1wWFBw5vS0K64jsTiP6usO9BvoZ07E
yk8YBFsAkkv676tUiZ5oxqXQLr7aECtgR/gVuJa03m2s6Tufkt8ZYVrmS5PgICD/aMNsTbR54aQj
d6O5UaQ7gUtHaM069suZovCudU4fynvhSU+uCH3Td9ItiqkP4m9p5GusC3cY21Ea6gWsLKijpSXr
bdIf0UsXJJW2TffF+cCGp5siCHsLBvFYswwb0bHAX4r8+e78P0kupmCvJV3YgL4uFlocvy3uoCPb
RIJ7KBWWDqaT8hvtwW1nZ/7rr5/hRCz5uwAXU5p1pP4XVvEJc+aY5J1u2Ys1Gd+hlPCdHPC1B0eN
gH8Z5J62HPFh3MwHXlUoSw2roP3cGPDxzIiDmwoYCniXwCT64dZbACzTkU3/SOP6Pgxqq0JuXnnJ
mgJSXziSytLsaArLNN2OGl8aViICT21tOVtY4jvNQZflQWB+Itf21Gc3Pj/ZH1wcCaTOeGvwdNY7
/u/8Rr4Ew+52CRBZaenl2+ZwhJINWvGc7elQ5wpqSpN+CDG9ujJDK5eL9mIdOw3JdgjJLTmCf31j
tOogLoKOGCmsuXovcfXP5F0kxVdMSRAnloG2AtEwUKpHZB8Xm7wLwCamgP5GMoo2FnVrP24JOlwd
fg6/FmGRnWEcRTdVpr/uzVpu/hdD5iXgDatcSKitx5V0IQT3RVQzxntOnIwz8tm7F8qafEBIiHJi
Ewj/TQr65YCDJsayNyVh+XT7vyzjkNjNCrB6V0S5TXpBo7kUyUSG++9v1hIXCDIMrRh7tS4cradv
v4T/6btgB0Z1LdH6R4t1Us6N0Otr68DV1exAotIDnohfZldrZsKw7zXbFI738MGFbX4yDejMtheN
D0FDGqfwgnJUTC7ehmeFAVPxdjoN8EWVInHgpQEQ9x8zGAs/ExF3kpt4J2Uk+TSI5txHq2TpJYyx
m69dOkSEu97tBBGMTbR6di/bExJLYiT72dSqh52T2ltlreZCJq5O60vVPrS0/RD1pPbdm7xRVAIx
GJv1Dvb8jMYfdwHn5RrvL7oIIFQd02cmz1ODWoTkmdUKQxo3acavTjm5sggnn7OSbLCM++/fCACq
UpQTtOHgExml9GoGHpVBQ1zk/5wQlyoCbSLWM9ZhPwZKBHTfawYcMo1RSZUjArpODoyuPF6x5zDe
jIubUvcsfe+1p/gwb03lhD3+xv+F75WDvumFsihWPVUCXFqel1AxFSYQeB9LqGN0bNuLkvvQlD71
K+dj+4KkT8ohLJwAbme9BR+9yhg8MDWzj4xiTXwUjOgQtQ3IyFvLL5UPu7Rp+UatLyNmFIbev4li
88jvHvWSl4ezFCkmdeDlzKx8G+76ZOFV8a6CQKQ7QT6EYAC+UGif2uymVNYZ7KALambRRjxxA1RR
RnCNRXeHUB7o1sdIRLqBLHFrGhO9s/MyCvUAVcczqbEG2yLwAHpH5b+OLVTfdzBbsUrZpA+UXdFK
/POxiBXkfT2fxZpg1TZdF7v4DmCrprccxhVmSZUXrysf/JvP8qr65+h2KIkR0TNCnU/umRsn47FP
LIUR3FOvl7VyfnkZBVtsS1Q6DmBHr1u/6KmnSazzgFtJuv0WxIH5C5UvYL53F8C0zv81el3XVsM+
I09aThrU2eigKlJZkYIJhTjRN4teRyJYDDhoH1cFZr93RYfBWKmT36aeiGTlsZ7krtZGVhvthNzA
9yljhlfi5Sr3m6u2wkvxeIl/VdeHC0AAshvO3N6xV0QrSNvKKbnzoCElMVe1uiVytjm1LF/pNfk4
RllJoF+g+GzjmQppCuluZe0Z8zqQL/VCT53dOClFFmmCqI1rc8VIxGpM7XUPGLNT/Qy1Wv3UC9pQ
XwmBSwPh4/RBgH0iRAYhHv4rUHOtkiUsGLafgXMGz+rBP8QHYaJCzgjiZnTQ63QlYKexwpEwiEMJ
+s7KOhN+k62U0FlDtYIWt7QIScDSiAqhFGQz/ziEtPaiIhBc5E2pcvF1RjPC2fqfG1nl2bjnp5r1
bLXUHlJ2TO65O0Ux5WYxp4sZgAXrKXsX+EzuvO48dc32jC9EzebSWTjgZIkJjfXeXaIT5dH9i3sW
9Aw+4Gy13wzjsEVcjkc5YmcRB3pR0+5TQDTZUcscJIzyGRk+3S0IfrgBA1u3bLCP8GVrkWNo6sj5
3gKzO+EfP87BsixrJk4ekLUu9ro8WAwYwTuOhzscjTYhPcnmZKyHJEm13IB321xsfg4/l6Whow4j
2DfflF3fCcjoQjF390dDzsnqMUG9i78XlyqADzrTQVyrxhnmm5aPp2kct2FSGoOgPFpJtkl2m/ue
3/rBPVxlqeDNHGpegW7nvLoahaaum91hXSYxlM5vf+WRzB+hEWUoX7itb64giL0chEF7JNrb/BHO
B6rhlrQgpMFNjw/xPXCZW3Xh0FTirvVVP7+Eu2NlhFA2BBH41I/xsgvSIPbm0yKFzmS3h5dOLE3c
takTrINS52dSSA9EMgVtiXOI025FUyG9/1WYgD5txPmLp1zrHOGiH8eQctjov3Pg4dSpxfB7+9Iu
p7Pc1/SE/XrS47H6YAX0s3QsBPPgctxYbbG4gZaYp4LM1rnOIgAT6VdEMpW97GpkFMmUAuRSWR6g
U/3wBG6uAbeSuZ5gc68giud+aGqmyuEJGEHrXNrMo47JJQ1XXqjcvbpeAagqkVe2ItAx3aFjjk9l
yDj3pg3kqX1iFMjJcY4AbHe28wPXY6gWgwi6jyeK2suZYz7HOw79204HUHSRC9bsCDsI9+n5+uBM
rB+xom4KkiNQJ3MtxboQTTqrxJt+TF0GxmzH9/FzRZZddFvR1fthZVGlFy1+6V3UxXpGIPJstiai
bs3aZBrpgnRAPRlbyWCC0M/ExW0zje1P7cqvKMTeJd9+HhrJBcAjLMhU8Ey5bbqV+Tw4IdRWWztY
hihswZ8pneaHYXqZcM2rpOvT9uJNXlsYFbczSn7u1QsZTQhbaHRXc1F3DdJ7QaO+fbOHR7dpoOfr
RcyE2zAVEaMcBB0+TQZMLgwG2MXMYo0TxSX6YgK0u6X+BZD2CZMXGYdh2/VMRXQaARV4wLZIac6V
eq94Um9tBGJp31IRI1axjQLXdQ+Bppe447FEOzuPTvhsH1Nz4o2NEi43Hbv/yKyPP2RrDRAWVTAs
+9Iemv6qLjFFUj+QWeOxDTNsGXRbvBlr3JlkctWcRND464eIunzMWULr/GSR88N0LG9LoOLYd5wv
IukBhxJ/N50ORxWEf3McF+cUrfwOwt7/dIGyl3TGDC7oOZW48SvSBE/3dZd5ua/UOO/g4uGaGrek
t28xQrMCRU/ls89TSYaLVLc4xAwyylta3c31dUcF8aGqVUPKxsNe9IkB5k2Val4VgXkLlqPZdkZD
9fP+08/p6ie9vfksdgwUMX4n6RFKsUMkz7I0SZwtf31VHML2fto/B7IA1oKQYEZ+xjNZFG1wMCrc
CeLZlnS8lpXZ33ftXTy6WgMKlt4QS2Az74hKLi+jH6maSIhBCENZW5ZNMFcBri0r/xcHEGrQfBu4
c3amruyKI+Q8ifk4zrOCtbwxRAcvkJ588FIzn25+uivCkEHoS76+8SOCr3Rp8IGCzfTpZWWkKRF1
Xas/FnEddi17Mz8jM3mPGiaEzargV33tUenwsIXB/P4DVbct1t/rg4y5p7Y8v4PMlIXHYe4gpiGd
oeuP2E+Z3zZjrFh1S+1niQrlra1u0YpETBjgU2RegxHzUcT94T/DVkMds2gwbNcU/Rly56hgu84k
Hwq562ReNbxpFkJL3yfUEGiabvFobVCMSSibm+stjlACYJEj8q53GAJju9DRqtv1KeMWyIz3R7z7
sARBxBAToga19HjjAKF5OodExqLHfwkOllooPr1GBzdpqNm+RLuyUzBDp1zR8IshGv/9lAa32V+E
F0rLqktab4l+Rl8O8iPw4b/l1bM1LgCRSGOj3RA2ax9vHIfHERX6KxDQLc7aLpO9VAgeAngYUqo0
Yubm4Pxecy1WIpUqYjNB+pnj4CJROsIzZeJz6PRNrq91z8LduxhPGPytIzoqhU3SR6PHNEm64TSy
FPgKlD84SonLTrI+Ayisw9Duom0F0Qtnjyw6qX+E/MN3TZFX7tiMo4/q6MkpsvR4rKX1L72i5V8a
bHAHMaSsMfrgCh+dCBSgT0qhK3vBQa2OylPxYLdvcO3WfT1zFClosSi2eVeq5BDbAY5VcSoDG26m
i71qxSvZu0NSVu2aP1BChfdzNT7Ev8hJJvS5QxDDLEklCBClvHUexNYmcjEXf9xIetq7oX9YG9/4
i/c0Nc/XvnlU4GOXs3BTFMSweiUDZyElPR9RNaJ6kFFt3aDyMd6HUk3DaQ/X9dDzn2BRPtGHjLlf
yUSqcNWgSsBtUmDfvw1Sc4r7JraDcAuy3o38EL7MZRcVcMlp9T0if/EsgRz8T1kStlxN5rEmukXJ
1G+BADkCvvMhTbeL7OnDKln8cZc90Wpi6Qy2FRfymqWxJtC1UTC2j+YZPmyibAbtdMNIuMa53XXr
hUtlAXrO71aG4RV5VAlghm234PrdhmVg16kMfYoiW0qh5G2UdiWg2sTWQamj2670Mt1j39/byGXF
jAzP6SKGNVSsU7TJ+JIOZ1wT4bM+IC0Rg1p/9PAALpO5C/WpBaHB5roYuJC9LgaD7+d+PYgweT0q
uTH0Gh8cUZC/EU9IIHX72RhlTZrndJDEDsFzw4owwQJfPVhsoOUYLGmXHflydLnc0S1lhASfyRGj
VkURJp8Dm+Raz5J8WZ6v8ck65AI5eJIP0AcZkJ+pyis4ZsYe89QSWGwCg81vWLU/IuO9YmGW4Wek
+3bUeoIzz4QvhcIl8UDT6HjHVS3VNi+e6n61FV01pJvtHujBbaOl4VHCSiFtGpX/mik1OikotpDj
FYpsV9T9s285TseoGY7yu4x6WUQvNWHa6csHl37CBD1Q0YcwaVVZv5mRVIYF12SfriEGeBjIQ5X/
IqykoZQp/aCSaehGcVWulSqjDAklaKWLlXQWeRKE9Z7o5uZG0cB4/fwJ7Zo0Fu2DbWN3HX1fu/3X
ngaeyigBCnxggON+JGxkHrWvFp+Rkn+5FryNm9cI0QSXMmMoRzHk6KpWeG3tRFxR6/zhmpxnfOHb
/XkBa9PtyDk6nJrxzKXnRlSUh95cbuKZABgwlJetHWD1rdaE1kUS+XzT6ovrzjR22CqAhR6om/Hb
Tcd9UllHl0oQo9WNeZT0daySc0v0AaCqhI3o54u0r9/B75AOemu6MICvZV8iRUf85309cJ3SdM5w
b36o3wcdvdMr2O3D0BI1zloeq9ShZUuymISZS2wEiCvS+6pHMsbk5Z+KTnkusFKtThQoKSk7Z0kB
D2bfHAH+LtgYuW9N6OBHDhF6TuoCZs1C/ICpOPCi9ryeWmcTYUbIEn69w+2tg6ntvxvF8wRkkI0k
8fMA/zew/BEvSfly5OP481hyPzxNQCbm9EM3AB4qd/Im7h0ykSbB/L9aYER9IkPp4HOd+mXaPhTE
E/vz9s1l/WW3Sxp/j+9t3/xR6z3lw7etRNtOX1pAdSxSUAWdkBQzbEUcLXCs8kt0qAj9aMTrEKLf
+X+dw7YVfnMVhw2VfwoWhZZdyTckI9MY8m0Zm9xUdSB4hJa1ckDiSR+5rODxCMAlEzqIcTJc2y1p
tGvR5AEAuM9yZF/XiuUIwDbxN1RFzzK4XK05Z88u/PvpxIXppt3HG19duHk7A9Ygc47Ta49JCLUU
jsm2k+Zyf1uhTG899lkKPXXd+j6MI9709FRh01dEQXkqeE5yYxQE92Lfq9IG0s5IovcYtCdkvHZT
+OIH+ifgcfYml+pgUL9G2wi/Te3NmrDkir257QmfPUmJwQGPVfVjIAv2vX/6qQBOcrq+d7ORI2PO
87TauQCfYl4+hbdeHtgK2QzpKOMiBvFb/jn/MC8JklZ03qqlI//EIcUVkmHpikRGwoiYp3Un6LeU
lwxcGYMokkul7o+gv8enQJaDSR8lCUODkfgbm1lKFe0mtZbyLClsGiB6+HM6lMo+RlF1C/wemPbz
GIQKDUGE43K8j7WlY5n4Pap7aSGIihHxS/M+QugGy0xCMihSdWooFvzw/nalL5XcG+mnk+Jc0BDm
jN0LDvn4fDbQXjHCc2PfDC92EpaJ/jPWAFy03CVPh0RITfZhMWX6fnTYT4vfCaG31fTxEysO9LMh
SZKIOnaF0qQFciDE6kiC7TrI0N02AxP+DWllY0TzcodKGCfG0TgQUC3Tp132MKjkDaLrlbKFluJB
d/fc1WmBhNv8dWpqyve+46PcbJ3sGkOWhrwH/cATbpJ/wYRis0/rPAyz71Wxbn93LG98c8ET1zAh
KoooHTL7XsmKPg/jVihWWuzZ8hJ/+EqQnJ+k9xfhQJtDp5b2L5KEXA9hCySxx2JJE7tGKWtAo46u
c7AX6wlbqUN9ZMv0APTp7vxTE7ragonoJhZ+gdwJtYDgef5UqkXM9CX+Dw/M2kBv0hzyIOC1FPE7
nOPlG0+TGyvnoj6mHeznXmezCERvChJCTHjGVsqBZluSIiwH8TSOdaFb+WixIHmEo3Mrwpo7DMXf
v57uhd9TRfi5VE48t6WeBREjbH3dZBoyRDK0/PGnUr3Q2bpmX9KgBuOI3iA4MsrgPKKIV13qa46u
HQ5xrN0PoJyj8RqX4IH8vzkGhPjI1F5vIyzO7AXPgrRHBeJ3oa6EOLenzem4ATf9A1NcmxIPPYw2
JNnxXsUlYXYgXvY5bi7jZzTN9UXDUygYzCn1cAX5fHIhNfcG9lqTH3cS/HNJHFQRuTbrKqpJYkFY
7g8vDe9kQKV0TGdIJN+81Qx4F5Tsc57ZE9Mt7qjsOJGa4fhehZBGk0WhPzFD72EXrquQQgSSn5rx
/MWZmrgc8OS3QjZ3VAPhO6odt7hPYiJEKqbA6Mie4RuOgxI28Bxr3bIhwAUIwumF3kC20HCHSjwy
mzSXL2r9XgfuBac+FdTR5JUq+qad9dzvY1eV0hl+OgmZ+bfLtsW1wg7m4SVptne4OlLtmNRH22L1
OLdvLmu8xsO84DRyJjIN2VDM3uXW/8ImZg1eMhd1Lenp0r2xtjnLNDr4e7Ma7ybuXiYlIky7BGJf
QC9lcNalEl7zrXPRHWZ17UTZGHH1SZrcBHFg71ry0YfbnsBow4cWR/GKkBKW1hF6hOhXEBSr0PMt
Pql3kYZFbRNO2wbEp2d2lOJ9aXRj0QfzUB5tv02eEzl49VzTfPO7qxAviLuWINpq/okzbaEYPkrE
oPZoeWDB3XotaAlxqM/10KLswP7zENQnGClob7qpxEoNO1Rv5EPHt9Tfx93Tg8gJmKu/2hdshiJE
JLWhu2Y4rF2B+QLhlMFlIRZ/OyVnZ9QuR061w16lbF/nAR4GCqhXT0hbgIA81Ej1TtV47YFyEu24
634+6GgSDFTqtVDQLJlr13B7ElQdQDbOSJZlNtGU3FvOa9MPe/zq3o08TFbwdRfw4uahBixDM8km
Ymo+pRUQI3nLMF5KzRachCkCCFodY8RKdj31OX3N5mceVScabrB/YWk51bvCEMcM+eKYBYsh8Ewh
w4OQK6JVP15JcXVhlY2hggxLPhb+3qc43cX4/FHeypbKfMvXUX0SHhsncQ2Heaxcw14VmHmvdTXZ
w89fyG52+vkZfzR32CAEvRjrp2tHj7gXPITiM22i1vEtpwDlqoz3F7F1UVX/D6Vpjzgj4HOpUTIq
U6ZHjN3Bcy+p6IE3uk0RkltgEZyXFdsBXUJscNI4DHIYCKXue08QIX55KDC004EJg2fcACIPM6ot
g4BqoPAY1xwC+EE5WPL3hkXSohARbYod5b07vhEJ7XGcYyFCStx2eho4m6RyrOTM9h5mYf/jGmcB
vsqYFHdXYOi2S8qLUNib/1hgSQmmFkcplQy8ZCxqu465aJM+ZcmZ/02POcO/wjchTCo5IYZ4CsQS
RJn1ZXwXB3oxxvD3ChXkRvIB4Y/hxuPk23ZWuK4BZ2p0RRDMwbZ4T0CLu+YhfSVvvERu5aQ+zIpd
KRtffu0DEN5EV6G7Ql0TdS172EtdwBDwhjyWwfgmoEWay7+qngGLnMjUjPHDQjrRQmWpqFboyXLl
QCm71oc+6uc1wfMwy9GACbcxpYlxHX/e9nY4Vox8xm85+CjfVAYE1trJaWtH0a9lTpfVsYAtquFe
AJJQUP4StynBFNYxift0QT04jtNr5VxPGeeNXKqfCv68uHm4dvH7nadx6cEAMCRD1QkZPp2UREVm
742YU1kBTNTTil1R3zQpFquy9G1T4XnwBM7fu+0GgIJWloAM/ONViALo1wxtpbCA5C3U6lYAwvBb
PqUX8gEdzoQoHiQevzvwVVpz/p+6iyv6CRlADTru4EATAbkKHRmWFPdIy/+fhVRpuL4Gh3Da7CRU
bJjgQM6vX7YuhClySuc18qTiMRjEUvAotMX2ZaJVf7vGeDoNNIsZeiNUXvApibOLI/4BtPEOwsvb
3cyTj3soZf0iGfAkUaMtahGboNQhgfCSv7e+OD6Yb2qbF/2AbyD6RALbGsZhSL6w5xoFjQ2RKLez
sqbCefPdxVyjoytxQ6/zT4jZsTLNgGsrKCPYhqzuZafsUxX+smQqDYVADLXUrLxYOkHcHl699W74
MKduWLIXwHB93lK+RxibCsv8+vwLHrEN/34PgTxe0pgIO9B1Jjb3/2xJKrK6rsJYbW6/pCvm0Dw/
p/2PlaD3gE+A3hac+ubo0zeWmQq7uuQxk347POMQDXsJn5hqlL7kITV3QntDiOaHchXojhIqdA7M
sh/Hs+lajwnubc3Nz+zDYutBMh8BrvY3DzuAXo5WOoOUtHTE+yr6YEVyYpwjhyXI9ZfC9GqFNwG2
toj3nnCl5SxSWEsGjvEK4wHn3h8B1QcGR+zBcCKJT4zg3mD+jHUehj9pQ0pcCJVRBAbVFDHG+O4C
VpmPnxTuMzm0syGyxMPMv/SWuYO4+kUJ6CuT2Fv6wAFcLf9DG+5J1+mfqgeY10dRdLT9En3OOG+3
btkWlNQHKTnDIQBV+HYv/xq0vKi/m32XiLFFoY2x5Y0q6lPdJDur/0vYKCHm3rt5roAiO7j9KJ1I
TvU7VdxPF6p0dWYMx7/rRBXvPiArb4tVSGREm3EF1u5TZuWBMSw0+p1DHldMzYiBLHbESqN6Aglf
5JhNNu1Pt7YT1yiesgEqWjJ+lWCzD+tNH3ZFqqja4WersW3/4Amk7K1rBf8e1N6hQM8HQlEXDd0E
8tmfWc1pb6cOu08ieohlSWetNJ50V/RKnCcW8d/X1TCnBXsKmjjJP/lYxnhrH6yitti52E9xhLnx
vitSHAya9UxiUd1hCjHwLXOSGmREGEK+G7V5idwNaM7LUiag+IUo/3n2Q7fIrGtvHNvU1z1HtAMY
vpE60UBAP29JSSChYomAbzLpd5WyEgiw2XCzftOWCc2qRA9pjf268ZwKMQnihDE/smxXkXFQtWjE
mQb4MT60wv1cuiw5tkfsyVZpN7hgYA5L5leCdui3RXnF1cxOUU5lHzftk/lxiuVYgJG75tm8eybT
6SX+FkQDE0LG8QSXN8dvsnHEWX4HW2kcC5wqWj63fMmk1bgVUHxWbIgC3DoHRPPcznRfC2emFt4/
oIw6FQBf7K2lkLWNgP82jL0QH2lxn03PqkwgOrDtUnx47K8fqR9WjRAc8u5BFFsxY4d2npsyJt18
Mg4pp4bbmwYQIg9fu0X82sNiSPwCnrQhoXtlXix9YRVaKk3MnzK69BTXUoQMY9JJomkqVDCvmlNd
n72F5xPxQ2dXYCZBmjDqKmku3NOQB+qQzwYVZV51tJSa7rf8K3/0QrGG27ten8dy0N1KGZuL6gNG
PjaXEcKUoY/fjtPGZW4qg9Ec8YvryBcHpfoSHoYCxkb/o7ohY5dGthEUMl5nb7Rws2NAmuo8xSlx
wzANIJOLQ1wKAN3xMAf1iEe9v1NB0zJWmR+b4i23v3IvN/Cns8DwqjDl6frU8uamx7+nGqFXOp4J
v4e0hpWBVEOo9vLm9wwUAXDxD1wUhsC9hhfM83rV+O9KvOyp0S2sBIju7dcnRpSom6Su1ZkW/UOQ
R1ra9YQSTbUTIWN6qFq1wwykWQqeaZey++4aJ4+bcDaRT2uPrlQiEZrAbiMepbqzhEZ4KZv/mwN4
jtoBd9dnqV7HnMiG7G6G1Vp+cwVZEROWPnyvyCOq0Vv/46bPIC2QdwY7JdA/3a6MiRce56USh8rI
okdStjC1iki+aYlA3vzirGZsgj/U1N3kynZzbFSEj/g9k4tk3Wbyv9CBmxvxhFMAFSHjajUDXl8V
DMp26H1+UiQLdQJOo6YRGc1BTl7ZJ6Sz2XmR4OrRKlOWhSlrNUaJNmkKhpzar+uzcWzpSQp6VZYi
8enAh6Fp2yXV/G6h8cDNYePsjUH6ErTUeduXkwqlztmDJ7jCyIXrV0TjUPne8QWPh2nzC844Bd2h
BXDuzLryY4kfof37Dz/V+OAuTOJ1sxn3zHrXLCjUQhzofTTQWKfKeWNBTR0BGUjPdV+fkZIv1dyU
iGdJpE7toyrXeEN2zIKjyhFaQ92vRGqoFBYYMMYYK2D1sWpTPfbkasqGiPfn+nxc1wYFyvkduZx2
ngLBWNB/hId7XXmwpiYy+kv28WFfTXA3Ts9W0RApMjYD0R0MsMVnekSVbkP2XgZZXJDoX8y1Wj20
GkrpnzWas0B0cxSNVCP+lQjHv1bxt2D/G21Gr9RmapkmHb8CTr3olC8B8/ClgCJMV65EOhQCJz8q
JHj1rRki5IEKYTnN4MzBFxbD8GqIBMm87EbflK54+5Dzw434MfH/KHtjkiXBTAPOYu5xI/6wcKo2
eXsmI7CaiEf7MxwPmbtYffyU5nhl2t/kjHH8uDdZQgf97jl4w+qiD9hqZe/KP3fldvz6KeuuHq8M
hMhzQ3g1N1/gpF8w8WALbJWOTQh1sgimVWt4BhN8IzTbiwQJs0mQuA0BV54utnDjlQp3mE4FUtLq
aEUBGU9WAEbsBQ3g99CEvdQkt2+DGBSAMW9DAI9nGO+wUR106Yio3QqSauvKsUp5p5zhG+Tv5Rzb
g9CCqoqMNue4r4XSwvgAIYrExoX8wkwqff5nND70mQ67WdsbmE0NlKA7rZCxkEoRpZ25K+GL9b8U
FqF49GWhbDCITixql+MflloCWy89FAVAJgPaWr3ZhBI0Fa+5st76YS+iz3yt3obJVDuLQAPvEA77
xbyzNno4UjQL1YYHPP4sFxEyZ5yn0luYdfStscX2lgWt13Mpfa+ycnNTltv9GWXfuHnVHy+8/JI5
L26cDib8fV9Q5E5HET9O/QvHliteipdMAlTCYzQIArt/kMiYt1VbV17Bwyy+AlvRjEEdAetO+iQo
uQsfFFbMk4OHE/kyj1l0/5y9cMYY0U0S2AomNEURtHvpbDL1wigvsCmNnqLOZjRfs0FzCsOUe7Aq
TMTWzCGjSds8/68c4g2faHIqGiNvkFoMCVvtmZpwyAwLuOxAlY4kBBQ9j//+Magak5XMDxNjJHoo
OwpMdFnuwTkdCx34xr2IQMzAJXt3VHfnjvMFy7y7CyHL7sXyNQCh+OnKN0eX3LWfb7TP2rHf+aAV
dNIyvQLhFPaHoCLk2COmS//T7/H24vzGGJSbeGzXQ1+B9fD7m3mKkFcewZaui1ppa09o9RFixyfc
Mi4lq/NWcPhHsHRK3ZS41hMTmbtHSQwUfC0LsarPId7R/aVnvHHY6ICM0lO33S0gN0ugGh1uKv28
yXWC+iYa5ZmCs4oh+ZWw8lgqedStG217Z5OhPoDEXUw2Ph+6XhsbkkSC0D0QpDktiZxFicKADqWV
RtH9qX7EcogO6Lu4waeuXcjNQ1OKUQtBI7n3NTiOQwC3jfLNMoqONFZTuq8ekQehcYKVI5PMt2KV
Zvmas2FBNYQRAWniIG3H8Eqi0jdij6xr4HgBoi6oFBOCECg9siw/ucUzWa2GRth8Vx29fG6BAuSA
Sxt8KB31QHDKdSyZg64hfYKPi4CBbUGD5OJhTicp7ntqejqo0GgGFrbx//itiHUA+znUlVS6fszn
HnsiN32Uo3EiV3IjU/qHXKB71aOoHAnFKITFFWUeym7TF1HUk1//91ubguafX+z9j4fQdITqC/9j
DSaOaD7mDeDDRmC7R2GWsS2kVPMzcikO+/UqQO5+oB6L4utqS+krasFeTghD97IM4yBzvjhzRwRG
p4gTuuowlx9zh2kSTfadtKNBzo1HIYwN5SdMFBXicmNq4+e4oKtmb8pIx9LfAovv6YGcA6ZU7G0Z
s2Aag1dXxytppWqiPGt84blEAatQhhSj9YkRl/o9UZPBUkpKmEG944Bd4bzUQtB5zFnbsumYNsa+
Zk/DjDHNdM7MrCWPIi22GuXCmnIPtYQUzFm8WVBRoPF9cwgqnKNO05xO4fFqbtDJDNcctuZov284
33XjA1K7OIbL70rHU7Cqiy1cHYbqlxndSRXKWxwmHLYzuCZ1MEvrM7IqpT7voh/6CJJ2cVjarX01
2GQabmiqdpb6j6dMDSi1WE16nWWLspfzoNGQaW56q0GSXROaya4zdLj2j4uGT+uDBwgyy9p7fUCe
ebpQVywqTPmBiQ8KvaW9b0XWkSjZa/aEDcjZc5DUyyLt3SFGxNwr4PwPSsh4oBx6QY7BN4RQHY7L
w3T3sT2M/w6N2Q3iijXWrSSHc2GiftE5P4JRa93fedi9wiZVfxmwpgxH75jm2KDmx6E/gQRzeQEI
TahLS1IUdci3YlYWmUa/4/ZPKm/+tTjhyDcNKQjcvP3cV6D5il+DhluE/16OlUqV55u2tikT9sHO
2v8f8Fws2yIIB6hZNgc3t8gwUGk1lrm36X0jCO77gUhiE8EFLDqkxYjZfiy0TgvQvzcBZCD3X8py
9v1F8UmTWYZxMNkPFsvqY3KkN1dJe2sIehZbD4Dd/BEW7imNAqrmPdvXqL/q+7/NLKoEm23kqkDH
pVf/xyeZNIBHc1F9LWe0WQYyHJA/OjnkLPFvZ6aj1J3O94xy+hRZ0jl5/5winmNYBMLbtJK5zyht
ZLu9maiDcQq84nbxXvmF9CByKWgxIqYjkdhCyBD2HvnalSe94THpSe0xP/9wmIe1o4cPPQK1Uwaa
OcUXj506UgzvhuopXikkk1pJo62vWUvOuqMLpvzs/FEbROQIYtsWCmgiHzn9V1KI4ryT9HiGGep5
t/UN+FJLhzZrFigVDB2zw0vmrV39u0yfSvasl948GibI+5nyJ9qaKVkGYRQlwOBAfQF0oBrkB9Cc
QiKVcwp4a9Jqaz/N6YfHIKiz0L/wFwndvUYSHyHWdYR76A0VNQ0nGO35dlMAKOBQvfwC1QtAtWji
RmFh7goaVDakjxnOpUAgo/ZC4YzpTk9fln9GGWneKJe54rAixFD9TCeP2GGzmU08y+eAZarb/xK8
mJNIpHOm3ydu+QfVK/nXZeksH52zp1vkW/c3QNrJEIYzwKiLtcb5ijKQ2lV1Sq5tH4TRX0gnOd0w
Ylm551JfjFLZFD4ayaDoXcjayjv5vlKSAjFS6djsK9Z3UXbC2GeWi5jiLuNk0SQYhdTXElR+E60/
luKKXrF6gNJ9rG1GVbNtsdQ/MRtgn3UDjcu1ffefqDKiHRbhQwB8TzrtLwvDQVu+4xu6Ne7/PjQY
dLfUaUF/o/CVE6zDX73oPF8NP/r0uSh9zNnNc69vF3wDzIrPa5qWtLfQ8K2qgV7MKaSIQO5Lj1e6
CmoXqC6IppA76d+mAn6Z8EUwthNw1tnbqd1nv2rvNhnnoR31X/HSz6haDfiDZkasKDCdZ6FVSrwa
+1QiXyvDOVFuMabeuP34Z8mYfLaMrxsLHSEesoaJA2j4Nc6g5Um51o2jz0bprYkZMwrY5GPRU1FS
PceD0JcR7keK6bCG0wGSYgmft1UwwiPXQp1Usq+PqmF8+RQ2yyfcusu8z+B9kZxTiy+sbrg02DJM
V/7fC4hevyl0klDKxU3CAqYOyz2PbYXAazO6vDsLnO5NhG/7p3XYBprGflUqdjaJmLOj4G58y7SN
0YCSOuolfC/8XzVCmkjxuPpFN5JL11peqFR9hPwH4495xA4e4u+jo6lUjHiAfjA3hOPPJ/nIKd2l
brfSu8b0Q4mSSm+Wd0wvgeonujLxXmwhmn0ie7DKpBvegkxtuPAZIE1zgzPf0luQ20jru/Nx4Xah
CMmBeanfoEOzigUm+5m5FqP0Xsmsw+WIj/wagxU1ER/c4vTsgkes2r2ZkYKe7iTP6JN4l8xIVsOE
29Os2mJRDQO84JFXhaEMLCsti8z58pi7OtBJcTAO+TN7+Ho3RArQshLGTNVrX0DvATWNssuyKTSH
Py5dkm+JHzLADDebHiJSBoatgoiSgv0p3ba6z6WbEIT8Zre0jSsQrqaY7iNvAhqpmhTcvodfFcBj
FIWu2nosNIJFyc7ePtAFTrBz5rMzgyu39sf+bRUX3rzrZeJZwpvCBMTNwtbHOzaXdflZhB0c2lpn
5AMhW5OTBeKiRHUnGdaMJe945xZudL5rq1pQZp9ZT0r/5QFzm5Bn9tkvvXnllYf2I5C22o794LEs
VghpFIxHE5LZeeEwrudVBafIGeUEUvDuv47obqu7BVAQekcwVrqLOUGknvp2t/LbRggOoeS9Wdos
HNeIQMyfkKmS/wvJoMBNnZ0XPMgfUV8Z0xTSOvFiQWxNZX68m0Q2HgIz+Lgv95Zl3Q7JjhtSjZaM
aEzw+z1vaumFpguehd41ZCE5h9ramLtPGj/hyLSF5DrlNeaS2o2Oe8A2qeZRw14A7o8Bwghc8Kew
Z0Nxv6saoIm8BoOrHJDDI3UMM7KyU8GBf+XpeI/UtPjiyCZHxZLhH5cWSod6A+3CnSxrSplcNGYz
QKQDS0GDutCaFwT7Q7EyZyCItLEnDtRKnbukhvndOL5Qv07SWOXGODlQx/PxT57vXP4wS1tO3si/
ZYKDaZVrGB2uCkJiSDYThds/VfcmpRqzUp2ODABHDZEjF9sCk2/D2N7agyDpkqCr3hOx1Mfex21b
/lXJH0l7oTB2wJQlhFMVG2YAKLsNXdF3XuJ6OD5deHKouknfgbNQOpsPpOaKBqLDw5qLWm3Ao1Uh
2VvywGl1Cojo+oC4rooSPefMUaHpGMVKCBG0NbP3YgnMI8GGjyOZSqH8vkAtRuiHlxSLb7awmhg/
3LTr35673UyBtLqw1KSmMQ6fGKsiInv4z01Xz+cRmq9Pq6wGR860B+5mgs7vNGKOZLaCVhcxq/42
D1Mk+MvKh9lmH+QW7vlF46mvViIag4Vhse35iktP4mp5+X+zxjOyFEpQSjgrpybgM0hAllpWzaia
/Z36AV8eJqEfxCAwFJQ4lZmH5+JRKnvno66ffG634obnUsHShzodGjo+8zfbBv8PtgpnU4j/66TL
2aPDEaTZMoirwrANnIim6fjSM9I5azNRi2x/HavM5b203eb7eQgfWuqEO+H6mOWUqIMLbS615am3
aKxIfmboZ46lTGmRGDhJNL6s4qsx3jatChkdy5zcr4RtD0DnobiZfEng8vnK9egtHyiBWTJSXGOF
SqE+9hWDOmxp2oVZGR+L++qUSYIj6WyIgmMYIHe7AisY8cwAPuVRF7kqLgEjgSd75sIRH8vJJ/1b
qLYge/u3EYJxliCeimTZuo/qwbz5DT8P2sk/SdPRRqvTeWLWDDX7yE8/wJv+1FP5uRK39f7qPiPo
fciYoMJH0kKW3Gr+8yM6bkrJuKDe3PPROEAfB5kRvZHfS5WVlZNotC9gPfN+eCRQT1pt+VgaoQwF
c3z4XygmpNWB1PkuGz+wQQHwgItVFAm9nzPh5+6E6FzNCETClrMotTjOM5Q+Z/RBZAy+QVOSEvsj
yo4qtIIYkRm0F6w5whKxD4h/l+l5pp1creMT3AKubR1lJ7UC9bT/TwDIsiZCfLJIAgEJ5AfzA+4i
PNEP3jQDutbu1J60yY+NR64b8Mgxf/x3nxy8+c8wDXQCQDS1LisQYeWRT7Tfwd2tHKYqY37f1EFn
bUGeDMcdV8zcoaI2mk+evH0YAMo5g4s3h5bevNniYIXw2Ylg3Xh9oXXmGHqftqsWFeAtniybVaKE
5UxcvsUzvTZyV69ZJQNQumlndbw+rKiXwQkEkShVkq20vcv7SiGPtgPdExI2g6ECMcLTeHu7/fxx
AYw/fmMIIfzLO9oAe+PwN6f6WXKUAH4WIfIXSQYBHNlNAbDXGSwD16H6bBUryBPQnuS5FevoNr7V
nWXn3ID5be9+AYSdyMrGzx6fcDU57xUJ57YYtl+JSJQRXsek6rWrGUV/0GHqDlxIgyZv8tcHN6T7
lcU7rv6u81iwN+LsOn/PIhg2Llw7j90gxTHQkZJnyXD0Aeawf+VKUe5sWVdl37Kl1p/zIL9KzypH
Q0I6YcplbERS0GyPsG+QvsxcjG0CsUadj5TzQk2jBX3Qyzf5FT6QmhR9Gl5YVQtFBjWRfa2u4UNF
HG8T6mH56FIsIU+pXznVin3sUOZu3mpckrkvjTv1Bbl1vIcK2HSbUveDPMyLmExRhM/7v5fNajMZ
3zbNt1gK/5SHwV9JOZRcBD6sYo+pxA7KMuWwhs8ZOekJ0vbiD6sBOQzVzB6wXhykA6qFyQDTGpTM
5NdyRbnqSVkeUx/FDY6m9S+27yxzMijm1TmpxSjTrnMHUj0TIXG+/5fjx2mGSL06JYvHkqB+HFzz
RG2xxRahXwR7R0JxSVqB85KbyYEPPf/Pgh+2N5ZejvwVCyb50kVZi3KrMfTEn4A+jgz05mTujyya
VF3pnf6nWPoaZ65+9zspmyOFJjvfiI6etoyZttA8tHVAYKEIWFQiTvTczrgPLPKR4R5V0sUUcjcz
0j/xuQyhPZ8KZX/eUAsPWOSrkFJey4KkBLlFoTHDw0NfLzNJ8UGSYA==
`protect end_protected

