

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YeJs3h9nPnCnr3aRxIBZUXmhDS7WeTgKjgxxU15evXAwgLO5UoYuCJb2fGld8H5MyDQGWc8UFp3Q
QS1bcwQeLw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QMDnsLueMbfhPqb347LcBnHgrgkl6fbZ0QORe+igLd+Fn4pMYglXhNwzAsr45PWnZnHEuCtMe3Am
9p5sJ/ms8icpsPjNhMihj0/+LhkVUeJEYGJR6AGOi4DauCIoKWFsirWy53ZScEPa2MEe+a32HUq7
sCpglfzmrbsWEab4EEg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F3FpAl1oCeVkGEm2PKCJ71S6Z3CGasBF9SuzLFWQnXwmvUuKd7HyekhOce1QfyX+pLQcgfmP3XmZ
qpZIDWOrbZbtPCk3pZcRYdM0rjk3gWPTq89GN09GyodyzYH5nERal74RXFzqDSlXYzgzDvsSzAku
WQ8fc8R6wi9d8ZzaPtv7Mn3RMOg32FvlzTpy40zwgHFS17RZjspNh23gqb62COtY3bIw5wgzOnnc
pwYSu+4rxmNM105eSJdh2TJiSEN9+pTEYMITQ2PUZ0OLL5Qstj3GHFD8/78u9ynXfzh4PnzFHX+c
DtImYoh20HOPJeCFpBeWPHfekXHEPhbC52n0dQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lq9ua7Pc8cPhzNKkRvioUx2DGTzaswIzLnIP4rJJ3cLZM5wsk5kiUTKl9rdBpb7G3yE/zCnmkGDT
ZEvIhQ4CGdpOb9ZjoYg0BIc1GhYnGIexWpvkFarqP15NwctZCibdBpj579M1D8fvQ9Xw1j6ILLQ5
gUYJd4OzxaJCHTNx0vw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qzr81pSyvLThhRepJmzjPLJdFa8x8hA7KFKfUSPL+CaCFf8sC6XyXYts+1DRzPvdthUp8ISKrFAv
jy1EBIdnZB3D8J/YmjzA1s/E0S3V/3tyfjjyCDrQgRkpjqKN1zwlXCzBMyGSBWpl8ENwa6XmbY6s
fYy2IxFIrKpit7mWPaxU1OjywKhHRwk63dw93KzE2hJmtDZhJmXSPJNkgusdN/mkZzbIYUj8bMZ1
mRTDgqzRIp9L2zyHSB7GfUn9cIiKtJb71ztIZtRMoFGfKpLMWPUiRhyoCIz55vgxKfE+F3ghCh2A
ig+nnH/YWVIR6bKztafV39mEL7utiMvwk79iag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8592)
`protect data_block
NtXbBfknTc18wtXp0zAxc7ebs8GAOS6Yf3MFCOdYBcsylK/yw1Ub+oOtPBoHmCgEnTo3ihDz1Zr1
3Gp8wORLcPpTuj0VUT7aJVOFOzyXj/SV0YLfdkxYSQOjk4Mu+eDJ0X8/x8keAuPTkBOjo/b+VSVH
RoT5/vONF0kd8C+eDwzYYLDfr9+qB4mMdRZ4jUMqBSx9PRqSyQK5zURMcl4enHVSVNtPwWPnghcL
ohziNpDTxH0a07OKGts3LgyrNpptJaRUpVeo5xtITW29eyjRPbYCQr4411RBXfp8CuDl1jI0Age5
lqvOjdYkUdfAG5vXXfriycXlc+WfY1z4PqAKlLSPrB6RJCq8H9iznl+OQ32YNzrAl9A/XX+SW/1E
heOjiLecCDQlxl+IkCY53Gew801fg+arInZu+bXu3u56egAagQzduRXUDsJUfEHOnHMut4T0Msl4
FZmY4kNm0Wsj5NqK0BYvCthzyDiG0MQ17pGTKWtEWmGxXMgEzJGoMq3JhvGlGB/VTtsnjr/46QEm
BxzrPYo+6pIlwHcoIki+nKq74IlT+3Qzquo2Ani1fTkbhB11iVQj6QmFqhaoz83e6wxS5t6ofRCa
arvoUhXOjO/Exl9tV8Vv8rYnRTkyS7xS+N8CXytWOLTzivEhSAB23iGav+9CAdUHOC4u1w9eRXIQ
6qgASMhOO8Trnnjg9pI5rhn7x/x7WVt4haqg+hlaE28WVOM40Xyc1Wtum+lZBg5btORx08Z3a5GB
OFJ/MOsEzvDcty2Vj3hT6bSS/t2ZVuOQJLhMUgePxLcuU/AdB2Y0VE3r8wKNf/pgUZEzGhjUaYsk
9igCnczJapwD0HHSS1IsllSjT7MfN13ZjRVRu3M5AqqDbn+gUN2ZOlLjwQIVvP2PBnRPiYoWMNLa
X6RcdIF0VzQ0OAX6QU9tlKyHrKN+6XmHDoG8gY1ufAoRf3Rv6bv8TciqLxxIdijUThnGO9rhD03J
BRkGgbOgkru11swFZBSK8rKkOVKx2mzEp5nD/5cH5U5Cf89n80PEOlfX8U1jBjLw4Owzuvqlp407
YxA6ORPUMA6yupZi582yDNxr0UgyDQ4v3f77IQMkS6+3qZBiD7x5UU2jKDp9Ih7squWxPfW36cSM
LTVXo9ec2xdLe86fxOZcheTci5VgPbYo1b+O/1kfBX4OtQcMEf2TbdvMHjw8nHHPhTlgg3iMOqlK
m6X5QlgmHwZ2lBToV0PGZJ4yHa2OxSVrdsVurJDDK14cRx6NNc2rTAMyWVHzLrrwqOGsXQuE9h50
RmhqJ2pO0ZmhGKw31zgStM84mbhaRlSqrJTzXRbywPKQgFsltzNo9PXspZEmtKwy+FNzZ6r2xGFr
H8NEgVXfFO28Efjfa8XN3i/sDQX9rUE9RduDhJurX2veN8jPAG7skYa+P6n0h7TP0sSQO1vV+Abp
jc92Vr3YDgb/GrHhfxx2TDUDUhyWHUmf2+SbdjXlm8/kVhqG8pnzwNZCUXsR9+FpMREcTE3jwWu4
gpHIeKPOjEhlEi1c3NlNkY70SUdlkEMLaBejnnQDgMZ2MdXAqPUGYOk34nNEcAo3n0UMZRiE/7DP
bXE3fg1tjXajtyE7xsRQHW+G0Zl1azToOGIA06BaNj8DYmpMeKeY62wo09/ur5f+HvPTuYXGXRaI
L2j4AM2dTF8sA4uQ++gpPL7i2GSUr6Jf8nCK4cHH67P0qDj8mxXKf/Ev2RP4mTgYKN7rRHSUVkE6
5CqirliIzlcVK1aIVx5ofpBZ0DrtwArLvP04l+cwP02ylYO5EYZkjBrxlrMoLd1vRWU1i66IvrAc
15brOQkZXevflKVxI7g6zl0qeUR7Iu87qEws20Do2pauFNl8GGBQt8OoUNdC8Oq2AYxC1vC5QWv6
JE57hKrI0BonTHKZIzO6YMpF7oUjLXXFENH3hM01nFKTv1ws7BH59KfCJ4ijTke40kc2QSKg6e3l
ws5sWmxWvqVj0AJ2CJ90FZgcmhqBYU51vVaHzyCG5vdUgs1kego3FQhI8vOi18dLsX0bOfQzAgyC
sI/+AZq8VRshgXzaMa+oIUyNI8zZ2LVHUSx/tVxoIyu0ySDkL1ULEHhKw0Qqe2tNIkTjzz9KaTCJ
I3/EUmjzm2NljY/GMV4tWjy68ITK4pCxuR/mUilhqAnWjzNhzsCdKB+jxGf4JVX2d64i+0qHcQEY
v9G1z63SUoXUUbSFCxI+4k0n5IDpna5BleniZfSkjfPfmqv9cO88hExPt36o4vks+XlYO+nhZyvs
BA4K8HjOM3nqJLIxgM3MRDBYbf8ISg6uvJz2eSlnMV1RikrkpLK83eafpgrYGXEGd6t2L1xkwna5
tTt9K23Fa1q9HgGhtm3t5yIhcx867jG2ybflSMnW0umdune0IyrkACy/lekKK+FB0geZ/xlTsUYl
9XEQ1Ue7S9G1p/lVVOO2JWwixAOv4MVMR4qPaYPBC1XgL12HB5FLKjMJICAQgbVeJ12d3iEfodTb
tNryDG9xn0uI1AJJTBVvZaGnNHTrThxH5zdFOhdHeQf9QKH5dNBUIIkrbZSdd+IpREZZeoaFQKy3
W36BgS/LI9Hkwz/fK72fc8Q81GtCL0RNLEtICeeXroJOZpJAUHRLhF6uRl41UXJ7F6r+C/xq/SFx
4wLJH/wM7z3ZVmn0aNyczbTYQ+samIYDMuMkQGpNh7o7WTw0SU8TtSSGI8ecr5o9hupwkRXMK66x
hoUgeGo+KZtr6Unr5Z5Qflf8bQbtHLtpgexuHPIFcSbkQl8p1cvorrrkLutt2a2HfLCVHqx+4tuW
gCv4y0Q8JQXcs3Nvf6nF1A/R+Tccyt7ctP7i1EIKDu+D+n/ONXG68VlmAzTJzLqbHTDVfUdS2QhJ
+SL0ZBmNvX9m7Kc8R2PbfSBCkIGZR5EjQ+snKqJOe6J0MucBavv4vCi/bjudMv65eV7ktU0M7snr
YH6AAMK1QmKNO/kP9kWL5mHBmS/EstDLz3TVt5FnfcRkncbn3cTvm3wmEqRsKixZ3kliwzPtIvHk
88i/nBes5QB+5b9Ia/2koXZfBU1z4v9FTQdfdLRwT4Uexb7z7Y6xPhHQ+6dd2g4O7ID8bkk3KeWg
Q7DrUTiepLR51Y//ewbsBWQo2ehiRSs3g9Ns45U5UAe+jZeufc9Mr121i5cvQckyr7fPpYYX6RIA
c06B35XiuSkLwDQXvzN+sWA/GK7FOcW5O1bHI4PUWpYHDIjT4pbgKmd+JBaSaUnQzvuxdTNnCHiP
kLARJ4D6WaUChwV2q5/6FSG+l3dUwn9cGQD3DjtCgWDbIGAL62vy9ifbX/HcumLJ0h+GwO8/CXMc
UYLfaULXHkHMnAPASFLiLvIaVDnAFUZlDteHGAardbxA7uyX/akDZ68UQSsIwsiiZ3HIbA4FKjGi
p1y11YWJB8d6jRLrTLwhc74MMZBQrW7bfi0XHyNHylQP3UlK2f7EYk6ozB+a7L0P+NlhaGOrz05q
1HKzqTRLwIGWGSDiDRFW5nWByhha6r6Dv9d0cGT9rwyrXPyOPMHH80Y/hDh07aHU/qQS4l1KA+ps
Ic1943i2+X30TZ2eh8AvWywvU3AwLzMqNm1gYrgdSXGPnoA43JxNZ7Z/qicxl8cUaX/eoMMJ4GIh
PdorsT6OoRr5bxeihceOitNH1rMh3Y1JM3kn80rzymPH/NDtSexAWi0NqbpWstQeC9zjJ6itOEWh
n/ct6E+HJq0Jx80qy/+sbVW+30YNYEy19ugl4qqraRbAj9APjRaIBFtfdS507MxgIDkF1xpSljpB
M/sEEsATp3cSDafLB59FKd49/ByBYGhFvAch5R25Da+wVna2590nxwQnZtzdU2RX0+Qg3ApOiE9M
1hKe8PaSo9yPN/lr2wX2ksL+6vwaw1fHEYFTmDbPTBF2WBgwDz6e+g49YlqhfY6rj08kNgskabsd
wowU/1in4+8UNNq/y91q4fvIsi21QOCBPsk8SxUfMeT4GFlx06aDdzHArHIy1bar9kWBYRm/lHEW
jrUf5mZDhAnOkouFNsIXNn6Na2mGwsPJSt47NpLQeXqh3VB4EoPSH21iEH0anKJQ7BEbS6dTjwOc
8eIbxVKmTmFlDp3S5hyfnVHxWRUNsOl3yOzRhhobqoxKYkOBwr59KnS7m0HfFV13LZVBCRUm6h7d
g236J+UV5WStka/358VoyHnvl1JMXx7ynUaQsTvSArBgA0rP5Uo5Wbwp/yjstrUtpx4jL4ujzbyo
f4nIeV/P3hn315kbJiKyPhNRYE//+bGRxYncALSVWzePXgYhzCyCgo1GgTGBP8oS8GbjZn9exUBk
TTKE0nX7yX5VIB9WOJmKKYyOYE5kRDEocNGW2fLf4nKb9bOW/ydS7i4lug+AAuJaREhTacyqwEaM
l0at7YwZqxWal2tC4wpJvTd1FBkQNxhFWc9xf5K4JKCO3tv79JSuCg67HxSiQ0G5m9OxItKwOiUb
2YJiHpdaccz55doCJiVBq6VroDSCSqwRMW6gwuF83bDLTRSqeS7NW+2DA3rFTV0JxrsR6IXTWNnY
1+Kd5ia1HUoWqeEefFvX8ZMbymniCSN5JMZ30LqZo/OgMCWCyhrPWv35JkpcNJVe5pX1+pi7AeT4
9vL0bhYVnWhR1CQFvIQ4MdBDzo6gPZzSxXmGtSyRoq+FoWKz748cx49mXrXVKV3XbsPXfAgHXOq7
6rD70rE77B0GltJQQxN4yZq2VMdlJOXnSkWfLcN1KTkwHE2dSF/oYzpyhBuOlv8B//QCEYZwmr4b
LOgsnFQH4F1ul8mcJJz7uM81CM/JQP/AQoQBZlhIbVhKpVnGVxMXrJAhIjgRFS7Yq4MQeb/dlEd0
UKn81o4wp3eZbK4v64Ldj15JluRljKZ/Vqara3P5gNdKnox9d/QLllsLD75dxyAHsFo8sw8U3Wgx
kmAikk1OXbcQTCN4kuR08Y2dn2ZAiclunFvWpz6OcgCeQxMT2ld9SJc7/F/yqK7KgpTKw6bcrEgc
AlfA/0bzeKBoCCiCZFbgWKDS0i369+PvFt2hSKYuk27ceGypFUPAGaYknOPI0S+94kFTyZNZbDDn
UzWtQo0un4eZ/gxwcux/LfdAoHzPhVgTOXsy/xpWu3wKBcAzOXGGMZDdt8MOqyR8ogEZpZ9gcOp3
cR0A6gxHJTfwetFDak/bBygoeYOisPeO496QpXo83MpbjTdli/H+B8WjmMQi0kdVycw4SFAx+i5v
O0QNrtK7iUSBcjf8gB44TfL6/IEH4tK2mIz84IChcxTdrmvPRjqqPeyo7qy+LsHBgrwQNB/+Cv7W
7M9oyKbV/72PY82/xBpPCwNpt8p3UOefkgv2XBAEtd2Khnjy9p2aYVNZFgXsv4ss1xAElYriWhfz
O81rE1YUYxpsUhTwuRAzP73PdwoffYb06s9papE970PZ+YemyJkL5ffWIWUbqXnHIRb+mUIQjXLg
g4+xZC0zKCbfiZFB+VCeQ1dnc3KJzmYDI6ZE1PZFHgF+QOwo3Z4xVPdpzslUTmxybs34j+ejvo2w
o01ZpxrdEB+rV5pVUUfUV1glaA8VVGAIDMQKTZr61F06TWa2XwXP/40sOOTwGeusAckPNctPXb4R
jlHuTiGvGCBTIYhYHZEus4SZ3EDXHQs17wFQvsM+A6xPZoeTieCW/b2izMoMdWp4Dk+hDiGzXN6s
TGhHtM7kMZ/T9cUtJKxMMCh/TqsoJcZPdRGSCjKj3kocXPyGm3BKSkKJp+DQkTXVSiIqa+bAMa1K
naJxQ4PiHyncKR0NifiRcmkGM0Y8AOZm5P/nkbhVA6lxMKvN+d4LbRMXXK6c3RbsWo9EG5cK+o3X
mfpRW44L9r9L6+bBfqtKPDFzeiBArhkp+C+yC51n1mRdy/eNcdqJTd+K8U07DvD56GxgThE2qCza
/T9YT4b/Ps5xklW/IisrxkR95koorEJCBTIYRdT9+MZKNJ77/TABFkFsn3gKH/Icov/MxPKQV+yh
QkhRdzQ/EKm2daj2FZtwJ0q26VS9yZuPRVwUwYk4BL2I5zOfLw8mBOBTin3BCFwVL9LjA+1hbBos
hduxEG94dJWzoQjgzMSZvjEOv0I9vL5TVNQlVOIt1l6Fjil0wu6BTrUkG5mpI7AMxEMXZYc/Rbyp
yuPpWeAWbDeC5f7j2sJCffYPzmqjPs3oQXkiQ7De/+jBa3Hdi4ReItUkZu826ejDM4OUo+0Pe6o7
bLq9EsW+Ltlr7uoJ6exrFCxlaHjgCthrB2cqPQI6FBGhBIsqu2QJuhzewt+lRtzRQy1ktDa/nJy4
AVVRhOZkWmlsbl2DMrQBrNuy9z2DQYkC7yGPr5lw0RXswNNZeTCJXC6H3MdA+gW20B8xpODzinFh
cgeQj8M5B/JFhmMClAxgYf3vElUiI3pUBVhxrxsGWFIHsbCSACXOR5Lgsb+qwrli65WgYmLGDlii
wPasPO1OuDx1YLAxmd7B/ywOUz/AZ0WtXx3iseh0GDC32iCtPvt4IjArt1AdPpWOhh7DcRzyghd6
SGg5beJgPAab9G/6KFKFfQwIOlXNnJMK1KryOl1Hj39I/8s3cxHMNqH3bHb0iqWK3rA7GFvhRD1z
mIckwPqPVT/eumofPi9Xz4ANh2ALnSl11gnm9OeA8NEg9y8OyXKfhEZffStx7mTcHUDRNTJ8uUgw
ehYn1GWyP0dfr66BeDO9ISHZ8JJ8jbSil8HnqO//Fx5Ebg5zZiJM2os8wabENRYjlR9U8sHisW8a
UK0Dp8fwE/ctAD0BJkP8vonI8cqluEQiJ8IfoM2XUctUaPjTFzIAktMrkbG8ZEHxd38mAgAoUkMb
Cj+bHbJHSGUeqpT54GK9XOx5GvpMHXvodh20GJcAnpcRmzx1eHE7dEb7FwOZN8BIVwfVrKU4I5kO
ixEiBAXWVhJKI9OFqIeHcAzhQXSyAIHvUGEPwzIAFmqSOkPZu2BgPEtC3p2ikLhd/oEvEw3PpA0P
47lN+sHFsdQleNa6YGYMdOkrqv7cMCPIao7g4d8uUM4ED210WN8Xno0vN2DWJDlB9pSuhX398RvU
T78n152BEx3Bxj0rYll7vLmihIUGV11cc3WTV15VlQC6Cnt5BpEFFXCAmf60uvPt8ED9e8toUxZ/
DE6pbXZ+2poBneW03eqqsUxuxUScJuggHm1t9TtL4ACmoYhS6O5cak6Ln4bEhkzqwuT89UijQbGV
/5HA7mxfLeTc4a4k/PjrRnCzyGRmb1BDOOpddiupL5QwiWNCATMn9l2+1VWsCuUSLxevQ28OQpc9
GpO9k4LXXSd7XUd3U/XYA3qFwHytvPusLkwagyAf5CH9q3iOX5f+etLjBlrhVx/GVxJWf7RjMtl4
GEBexCs884GjPi8CNsQyf9XCYMNp7CZDblZ3mc/Ix4dH6BSTBJnczuc++aAHoUMqm+C+gbWefURs
fkdgKfgOsVWq8K9PKPKPg4sD0DhVjxqXpBIVHnUYhBYBIXixWyOE8xePfuGvCkLlaawhoMXgI/ha
I65PlTHT51Fmr0Psn91bceabPO4UrRTgJi3l4m11H6WauasCn4ezV6THgaun70GbupT2hJXsU1dH
Yab45kLaMMiid212mUMD7KU+3hO7uPhCPU9ugsPKYUWh2CnmL3wxR6I7U48DVG5dkrvlOMYS+3fL
A2izdDgZOSq63M+i2tCsSQ3/OyIErs5N5c7X8MSmPYmVtTad4J+YeB3zgwDInJPaFJ3ktQS3SPWi
eY/HDpzuKGErY84KTzaItwDvOqEq2Oy0Y1NhRWjpBmWDtmcM/BdPMbUSE23M37uotb7k3KXS8dpz
W9aL7xx2ze98EU8xIdoaZRJwzW4lfVp2AmShptApUkmirfHa0BvaGdfW9e0drEXGtHxoud+hykMe
IFLBcTMzlKMqm7/ee6+Ct2jvyzlJGf3YCfQCQpHmcsfoLgT8KVgyXRy/O3scAjjcPKQQh0JpyGTR
WbfrT6uHLiRpMdHnZPPQfEgDHDxjpaF2T89fNB0YCQsjJnbe1hKh/QaZBTR0u2uxIOZ0pdHZkYLZ
JIOfPWEEKZZUnRpMGUxXI8hMZRmtdG8yNaMEYAc5HU8tQiT+3xtxwFVuK9yhBRdyc8WbfM0w9ovT
cdJP3afzCrGs5HKv4fIVS/me7WUAEXo3m85YPtXHtRjxDeJ+XMxeDl9xD6Nz28win3Ag+XKsUz7v
JND9w2TDMibZHdmicqG9tpktGfVGZEbgw6Kz7rFKTQAsdQoKhJoWDjnBLEmOiRAjvabx3OLefQ7S
VZiwqy1SKC3zfR28Mpb5QyFIJyqJhTI00kn9idYzzOWSLcUDyDVQ5sW8QUVdIJjBsHYhINutdbcn
vWUMIvvGFmZQ9w1CM/ai+lPz7YJAeYfp4WN/XhljMyMhn7KQwJmnct00gn3tbOnlGlR6CXIlhHn4
37/qGCv8AEN1HhFj191AElT3Ulgi/nRWCN0rqaJqvSRQs0BfEY05eMMul3eUADYwgxenOlLH2KDi
Pt9fOaxqE3ogotdqR8yC4MVlInbg8ujsXgKtwAafPVMNhBTA4WTPHj8M5vMI9szANwIszuM3+n3w
owDptcmtqNvwEXHh83G8hJwDiTIIszTqAMZuFGyhN7vVXRS66oLUwqvKC1FCvDWlYxgh1KVuczl2
W1nAVl1m8AJEAlmazJsPKHpVkbENvLKJY7+/8hv/DSo3L46HYeprzLzlR95ZWi5JldfpdXse7aGd
+jWBzVjEAHXI+3KLvYbBY5d7HB3160/3wjux63JdG6eM5OsrSJzELffLv+fEBhjPzk+cwNWwrGbY
/N2icmMOysUJo1M9HjYswKPYm87Sdt14vTtSLwe3p3mMwxwFNpnmjG4K1qPBofl0NaSZGq9ZdwQH
z0xyycuG40Wyx7rTp1WhD8iTbH8wfn69nT5xjtCLIgJzJChcpAGG0Ug1EPyRvQobmhTWYZUuTtak
oBEHKjdNFCkiOha0/K4aoWeXu3kjNdsxPqsLjLKD5bZenndnZL4/osrxNls8Atn/zUNbhDjavfbT
RGMLH1hHaEJsy7c6jbq5WHikBKdJ+1KYLA2MCwy94C3ziBxt40YNfbke4K/MbQbjJ4RzGcY5/Fjj
arcO03yG91VYidHysjFqrjhpRr4CxH1v6nb1s+SCckLPapNT9GUEvMVFwUJtjEo+fE1o+buwZDDv
d/CATJmgYNI7Tp+OOXs/n7dp9+4meO1N+OrDEdVbd4mpShYZPXhpjYtgL8hVKyPH5zi5gieKu075
iILKKvcuGhzed4tzmpqh/JuSE8Ma3DVh9BV7eLaTzhPNal7roB2OsyZrvjgtIVyutRjjLhuwP3AK
4uIfLRiUvn+67kgPTLQtAu+5M+A8k87JfOsTRP1ZB+S7IUAJXhl1uOuMRNHgvdDCRYphGNSgX7ZE
Ofb35PqttsLfHu4CnvGhdFoHaRTqJ2jJ6mSequkH5g9ss7n0vSykbXWnyetpXP9P/6edndo9OoDB
R3lngxDLt0wcWEmhtOwlrVUNNcVBSjNYYXi9e9RHiLF8lrtpZbk40UyCQybRj/IqPRe/080yEszz
jD0x2W3Q3mK+7B+FBbhRbz0UHfhykSJGgaweJ1vxdiMXZCRf18h5/Na4YQV27zgyJWKhOiPuNhcS
6kYmBsmynHgILe7DFXaIP5ENhX+pptcWXVHHSvnPELNRTdUyUe7g35BDX5hft9PIDXAthJLBcoax
naZEMR6acl6NwdQSX4QB0hQKtlkVzMeWFDChx8/5+m0c6uk0dNNM5lEI3l0Qc99ZpXdzTRX25AM0
78voWtqro1Ykxqo0qtn0FButvfV4AOrAaqiXdtj88htpIxzPCo/E3PpZktknYAApIqYKcsCSUjTr
qcaA9QzzkOicVWigi+laCGi2gDRCTtfW/W4egHn2azRiOfe11xVbHe/ZQJGfpVqd4eZVQIbErBeF
RJdN2Sr71h3wr6bx97kRCol7joZXkhGdZUjCYP1d5FPOYjk6LP2AZhOw/9Epk/wwUVUVmelO2cyo
dDDHX5dPEqFoFWoN8/vbkLogBAFI4vcsIvQOP2cneQSod0U4p2hgGv4vLjl8boKeap8KEz0DqB7w
u8lpHQaTzOON3/Qpb31ISQ6NnEGa4mV1u5fW/kHcrD7M9JPup9dRLzjT39RqWxbWGN/TUM49Tag+
oGu3iVBAtALsj+mfAHCTt9eWZOQCPHkQg/aJMExeLcb2ChhhxpXyjSCnoB5KG41ArQYVFEDcZ76x
bw7N9hjb9LySuYPNGvbzW1OtuxmEL207xl7EEFvNfYJ97EVJcIG0OFwA5DJWtW5QpkZIF6Y7TnfS
HFIYEePQ8swZP519aftJ30l+xJqk9D7J8+bHflW4YgsMA/yoDsphJIkZxBQmmxBtdiR0z8XHu7b8
fkkmVHidR/H3lpEEQxieX/F3eDtmPHp4nq5Htsz0T9pwoWeoGn5St8Pu//O6ZtheHJ8k9lxcTDio
xPXC1BR8V3xbi3NlUz2hNZQuFll0HWiWVq2urRXyaNKACjA+XmgZD1HUT+z6G9nRckJNmbQOkr3o
nPS3E7xvXT9Y7hGf6x9J2zTRcnd7AtxHkjjd/3HLBI2oeapCjAr9Duq55tzhWB+ih+C/YATyw1Ry
lmk8Xo7K1434uu0S2N70loifTKBskFh2ck3HKk/8BizWqZ8F32jxFUOTnKCdpeU8crGVouoOe5Gy
0izUD33oNT5Q6aZ/4r01rInKGjWNnGn54pt4K2F74IDyxdbqOJ/AnJNY7ZWZqyQy3q7uZwYBHRnZ
X0Khr7g9x3Cdl5rFEJ3Qg+KjN5J973jPecOxQD96a7dbb8ysujD1tgoisBWH3pjbC3V15aRgS3F/
GuHcxgXIEucKpdwzNYygM3qw98yQ6u6F3RounXUFCBSlpH7fR7P7SEKWioP6/106SeU9iBDKzOSL
foPKFKxoRMU9ql0eDbWU4vzmK+8BmidBNW/ThmaoGgQNuQbxO93FZKocdLSO6k2/iNqcy418NYxt
jypgP53AfShhu2tCbn2eQ32ZM1qTyNHdVCNlAnM2npPsrY9iyEjGY7iBZ7B29drPO55VE72RtJq0
4Tksf2v9nak5WaBU02QHGTrOEBXGQt7l8MLTsgMNyenyjkKPfqJsRP8gHrIboJhFiwNxZ1hj+7BF
gjA8/SrrJbouN9gMO3LYFmECX3igXY+jWjdBYofYRGKTaSYfaXuCgS8uoHSYETAffEDMrFgEKEOQ
yslYyWGbvLtKXGOyOKP8jeo0b0wLFMnpANEiCiZ7v6OODdYA0bQgeOKCExSF5vONr7C76l2bivE2
YYXrtKHa3vFVRCS42S2CuTNxyf/JZi4kz8aP4R9xxwHvZhBsihLAMfI9n0meo1zaYPCTZ9PEM/cG
MJ+6U0/3syJGYhg5l9s1hlFCUZ5zUZz7RvudyRD2GY9QZPyGA6DnR1FZ
`protect end_protected

