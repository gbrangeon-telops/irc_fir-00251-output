

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
b5iEwcuh/jbBlgyw+948d3lvWBbFsOTNVYtA4pJb/+7lAHor6DKhd4akfRWg+MPGWaTgwtrV3Hjr
bBdLdBNTBw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VtyA/tLK0cCJJRwkcmojHVnJYFSH/hY10K0O1xHrVFcESK6dXqpZL9jghTqU0K8Rgfgyj2mbpSmS
d3OjaMJOT/0rjwEIwUBTQhpYCQbUdyb5e+tsu6Jle32rY2EO1nN6daySTSkOW0tup2zZBsIOCr3t
+ejm/NK+miEBBu1xCLg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sf+0xczGTqZZx6dcqp2GTylMp6ojNl/Es91rC3p2Qk7Z8FK5U8FSMHtByvmeihj5pitp5aOxAIcO
cjVP1mZpqkA9QTc6UkTBmHGnHSpwqkUrzOtsT2ws44zFj3ryr3hssigeWwtnVK13YgLrM+5chsUj
26gA0jBZIt1YnLsbFPdAg3CFuuIkHWQ39NEQDeG2BTbW5KtUVyDTnpctdLn+1GQ9lYJeC7lVtfwI
4B4xEL5dhZYik7uaLaobO+7jlipeHv29o8EQsg6BnOj1c1kxrXtTLsKozU5mRUSyPYYAw5cgAAvI
P9ELz58Fq2bFhjjPjC0ULrxEE7cl3R3lE+lEcg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qzj1t+dWRPGHMv8nVaAMZRu2BQPWmF3UL/i0LvBgsHGjHy3fNoKTLAs04wnbPCVtn8n3ytCSqZ9j
YDEGkJeQd/ctkBALil+9bfKGzVPGZiyWs36ilhf0nuaehXbM+Zt3Nfkh/wd1LKqVrJhOB/A/iGYL
jRkozXf4ccRU53dhQZE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eo3jj49OyneaHUaTvAS2/lR4/3L9GHwLzRAoxweYog0SBxlqFd2rrO0OlKoc3GfXgogda87o4tmz
l/UHxih0uJyK1snlhQ6A1EHKpMBpfD++gCN+S5IJFV1QgpWejKXt+0a0zp/A429l2cS7KMD2pUZc
B0C4VRE2SAMGJhfx1GIRczPJREH6ZIkDU1qmMs04rSp0PaGn6eV7+euaxeQcoqowg8QlRFnxfvHh
5JrqhxNCP2z579eEXYXH3AWOzWM/EnKEFUTbEaxMGP4W7RzgRCZvuM41apmXDWTVjEj3gQq6xKn9
0OWO8TXN0ID1dcJmFJe2x6yA91duGkuqWQQaEA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43760)
`protect data_block
1HmfGW+8QULY67vQR0EZg5hXVlO4R/SUAKItUECm95Kl3+KTwnY1hOGJ9aSuuxyL0Ohxuc2kyATI
xhPz2leagpQxN2SHAK+ZXU7k8z2ibz8ffhgsDBFOtixekoZ5sw3cgTez5vXhE3qFq4bRowE7jAXz
xJJA5Iv6mkJCmQ5BXu2DW1aYfHb1lCUpVS1PdHjeJsLKefFikHI1foitJwwz15h3ze6+bGxPfhp+
rmI1+rpGUJF+7fcl3JlPN+rsWHp/x+R0srJtCYKAVdNkNBkbG7nJEoZ5XwRv83PtW0ATUlOCLuSa
kK69gCAZGoENL+8PjSDwhSkMzfgdAq95vKlfRKphQF6SyjSX024aPpBuPFOYEn0ikfPXfUklsmQX
GDRmEi3Ya+a5cMS0myfiNd5nFf06L0l/3KunsmsNSJIBIJhYcStHQev+uL4SqOE+oLQoNAPzlvIK
ibxFP/QXJsyFa32tFsx1csdV9QwfNQgCy0LxnSDAXxGNXyUx7fmQsKtb+A6kqipjGf0j3jziR24x
zM7vAQDZ6x5n3gr7w3oBRrcJdeEvZQtJGl2OugixsjXEHy6X3SatDJB2Rpn5QhjRJcWg96XzwewW
d8hi6WxjaGRDyY0GjIwXnrrUv1ThK4YEVwGB90gE2TLB9xPu5lOc6RrExg/5GZL8QrjLjlQLxbpz
dS6cI9NPeQ20OYRZCGq8CNPeabz0VxqBw634pk8RJxjd6uzps9pebSmiq4YEVl4zAacC61hZXBc+
9svqucxDrCxVeDg0URChmEo+apOjvsccy+S6pvyLgjqVkR4mfXoyxaExkd4okQAeTSuc7OLBJMcW
Qlouuq5kZdABPmBxCIZVEQRVBKNOKpIA7RPZiEHOSU8+67aC+3vQa4oovBPoaWunLI/IMelutPBh
k7JGng1uQ9BDrh+5ys73E7IJHy8Fh80/9occGoYJ+24ERv61YqAd9pPB4DsdIbD8zLgJ+dm3iPhM
U4HFOoc5paRADko/DUmjrEs2agZZgGG4BnHo3LjwJrOCN6m7KjtsiZav54k4Cpu0DDTRx9D3roSE
i0lDqQSuuGlMPNdFqgdnjx8BcCxZaovBKjhXLp0xlt8WetERAEyLTyAuqK6d5La2EWGI3ILjke07
ZciUY1T8FZe5iSzuL8SL5RjTvG/PlCdX0y8rcgJ1ae2VzWZtCc7GbMKppztaCZlX+Zdk6K5SndQq
yauYX/PJCH5K+7Gbohl/3YZkOw0QVoSyRNoaB4V5Ax6R4QJlFnJfwEOHEZBEPluB9d2aDa8ztGgN
u+kQeLwqKuTWdZHu8sT5ymq/pC+fKd0e98oImcPzJVh33DuZYzSD18KbIasXKFxkWVhejgBfHkyM
VBEuK/C2Oo2wyuZG4hNwpzOhkLvDoG1BjMbWG4hdY4Q6uDlFoMlE0HxfIXWnwljVUfF4Wf7KzCyL
ZGZCOq2tLsx42e0Z+bZiqV5H/b9EEXrZCEPCA/3P+DzPH6otPdz0TTh/NFwDMdbQhevDiFW4BPv6
Dmj/9SlDEBHc9vq9s7hNkK4zwlfnutM8Vc8L4/hLrQZAJFY8AGXIPUsEdI8IOT63E1E+z0I6HSZW
gQ9uL8IURZnYYrTpzoB60dL2VxJtEOGiR5NkYDXZRfmT+N8ebmUdwroxxRNNRukQ37TcyAYGJTEl
dlXbt8puSBAoekcmdQhpeec2f+LLYSOVhQqOGaZm8HhEQyhdSzOKFYFi+dmSWz9meG9WXOLhVO6l
XJgCb3ytGW7B+npmGS39ucD7rgFQhQjbcb66h0htsBiOMvTZ3K+u/H8poRf1cfe50bSr4A/bqp1e
QpWuwmUTMLoXOnkPQmff10Egqmkk6z/B+pNyN/BYQaAcYHv+kdEqwaPV4XsQITTtv3+zVO8SSuXJ
NSKaAtjlbh3LMOFI3uueA2Xk5bcCXVbUMnkRN785zxaf7cV9ArHzpnft0ph4HbbxJk4WiEWb2Cic
qBcQknTOyR2RS5UikRXF0P+gz1bBvDPajsUniTm/PzuVIHPWljEPvGWj3PotLhukBm3NR5QQAzhZ
Ebx8OTZLmKdHgNZHGl/xW38mAnZXMgoF/UDGqhxo+EjK0EejenvaDWl4B/r27DtewqYSbixlDiDk
4OMkoPSQ6v9rtFbNbvY0u1o7kxYoqNS+pSqHnDYgtcgJeRUqRlpO+ZPNvq48hoQShQUoczbbdfwn
r3PLAgfyyf5yz9iqM6XSgN/FIkh7lVyjvDFgcxo4tJQX+vBw5U9k4gtACktvhNAQU8LZu6sXDNOK
iI/Qc2Y/VRX196ZaDg9q7ZXTWYpXJnzSSITl07/8zXfs1o7Q3EZ0t0IhSNxRVINTjkL2sIgIgYAT
ahoXxVVtL+VVHpEBbNhL9yHcmTBRbk1PMZCHSGiIyL4/KgufYfimXrhR6GC5KmHjH9xRoU8RskOV
in0XeP0EQg5pPmMULFmYOSgYU8Hzcte2AVFRx1pWHk9ST+mjW6jClglh5jOVNy0wEyidrZsliyHF
jP8qVc7Dc4+rxbWUCvHxtdFQDgAv44yEC67NLhJAeaLKAGkXQXRtkuc+h17bysRmiq17OFmWROll
zXKy6rMCvGkYgmD2CB9yeOmltMNdXjqpyojvLJhBNNXNJB2Gn5SarfApmtxKApyU6jx5t5471rOe
AzExNi8G5w8k0zawqnppxuS34jEXrcV9YnZASh9Nb5GCAM6YgC6BvsWEWRb1FdiPaoPzwgFzVSGO
czYt/1bcnrC+aKU/ieaWba4sKMYZEIkD9+VrjfoaOFqeo3ZDOz2drAMM4AA0z522mFd20COUlrDz
A5J+alSko3j41MFi20AwadzjTOQ9wItCWxwMUarNJGS0anrsf9rrFvw2Nl1y/DC8eYUN1+yncva8
WGILCYM5cjaLCwuuUKmUzlq3JSws9YwfMwXpcwdUzee/RhXDkLxvQaC8qbgGsC2xJ0LGxLNQ9f5j
jQlpXaQ9squRnY4QpkRHc/IHcd7X3j+FbBddWfbqZNCM4GClNdqcsTLKfpHWI+x6SlNGSzFPAtU/
rf0/cYLS1ENa1Po4ayTUN479069AAIe0SpHUyryF7KyCiOn1jEBTX03wRrGV0sN8Um84hORaUKIv
t/nPr7NPD7Mn+B7N5H/Lh/tcUliDGz9eA9eGnT3XWzx/hQUdFgmJzQbgAWntbhDk5FG/bJWo0oIk
vRpPRkdoftJwjNgBgTX7bDqdgWYCSXG+L3Pv3wLz2bB5TA8pRFAnvV+YeHIouC0eoBR8ft7TUKdX
rOxf/gXWRhA7iYQrW15ETvoHVTsLdnVDd0QqVGD2JSe4r73UH5rZJmhECq+hQfeQGi9wQ/ik0+p0
1j+sdimMl9AUN/K1CF4UFgQiO2zs2aMg4FQxw79Flx/ybZlyqS1BukiMDavf53/laT1grqdD3FSy
wPP0vGIuCEhSak7cM9cCj7AJdcTLzrFJWsG0UCHjONMiREDeYpz0/ZaJflfOLYrKai4KSe9oTGuF
/UOeNFiEeLhfHD02QNyalQGDm99FpF4cQx52m3sh82A+gacGbBd59en8m7Ct/vH4LUetAq1dcb/y
0f+9UsYzW2d8xlZgXMeo6MSIzVfiV/FASpU1ZkAs3om8YdB7xZmVGgCIBRXeF0kkVqOmTBVkccOS
Xv8TC4Ml2tlxR6yJc8JAZS3ZTqJT8nCNrahXGzvmQtwYKigG3YRN/qHMm4tGwqII0j/1elq7jg7L
cTnq1z4EOA+r6pToQ++jDuTa8untMXxwGCSCcTGeELSupz9N3u6abuWiuLxB1qdOhAfVZWTJvfzx
0eoXRlhd17OMKxXaILfX/dE2xHmbj4ho2jWoAsx7mJrJdycOrBTAXsq7pKxzeGYnaDrjHXtAPPeh
LiT/c8Kn3yvn7Tb1c9kjYf8Z1aRsfx5KivHvIhf3phSAZlRgMu3WLCSyrfVxMyGmBLPU0PhKM2di
VbS8LpylOuPbrqyOnkClExjVzcDUYCy5GuOzeazZIsZ14Y1JOBr4yz0oamwQsa+0fr5FKZ8f3U2V
XLvPvavfeq4ThdPUNEmmHb9yvB3OdbkQlqswJCHDL52TzkO5Aw4wAtsQW7UR86aSFTxzgLkR5eUB
/fXGLtYdzYPe4hHlq2ee02owhOTV2P5r35dm0oceSGTT1tHaCg4e/YSvhq1XHTbVCdaOIA/Wc0iQ
dl+IikAS/aRmnt2AdpIz7Tktt16XES9BnkiaXWHM/WgZTEXLmEgWM6B28ldbaw/uTrhczOPt4Xba
fQhMc+MYFG6Q9xayhaoAE0K6DkBzyZd5GqNLRHPvn89d7Jg8mEcqykgVgc0DCFOAC6+KD7BIA/XZ
qTOyHA0Y5kGMNPvQ7tTvJDEa6FKRL4Uts2fA6kKdBFacMeAnHtRCfKLs8dK44VEThq5o3KNue8Hd
lpwoNrdFyPtMhIW1r7eo++8K7I7UaOOE4/Z00Zqb0mCQZDFnH6srXPyFn2n6uAXDJ6BNR5XpGiVu
A2/8DliJTNaXpFbQeM0PpCsBu8Nh123pu7esKfn8RpizOfjnvvzTpYIBe4MQjli4awb8YCiJOk1e
liHYN17yFz58Vf7YzPGrMfKdKXVUNbPdhhHLcCuomTY0spmYOKtCidgyKWIuVoPx7D1cG40f5a1G
HrQYFlG6xEeH7LfpNHPdPbQO+LMRmFv0Q2vU3L6zP/MzxndzgjakOyoyiHA6+wTZl7syR7FYrFvb
6tsVFXcCGxtPfGzxxXqQRUFIlJ5mvP8spMbYQGtMNR86ab8xkXzGPUx0eOKjshlY/tf8hlE0Jt06
pMDrX3X9TDbr23z7jxlB5YXc8Xd1K2sJTc5xUiifJ9nsrcMFvJIxyd4J7C7S9RkqYn9TxUUumR+Q
Fsd29NIvi4dygV4T5+3Ov2M/+uDm8OoQgs7EeJQAwJ+6KrtTZdfj0Mn/UOzTnDg0vZVK30gy9cGC
VQvIzoEoBMQDn/1wXoJ5x29jwe7tHSHOFp5OqqMxDjr4UPUvIykTRtZs3huc1BYtZro2Wa2MW/ys
WlcT6p+kRPjhsOy47VwupsrAiwoINACBnU4NqYbEAS3K0JJr9ncq+eIxgjoCv/7vrTDs72ubeU6b
T86sa43x/sw6lXc/mNF8UoT88L0fWNThK0BdYpxrj2x202nAAkloidfBQBBhRTBpV+C6xnaUdM9j
qtXaaY3SsWnQkRbnDiJwSkfQ/eaxvaEBLJdOpi2C4dPkEuFCcR7F2LjK5WXHHPr7rVb0J6Y/s3lZ
kCuy8Tmpl/3zOkjQb+YwzzarEL1khQsn4Hl4DNSuEX9jizPQmBLsXQv3hOnHqtwqSeAZe+qrzoSq
/0LR7HiCX12KoQXTBn29+VMclMKX0ZymmRdQC5s4gDHZaQQsyCeh2+gZ+NsPs7iW8NGzbXePMjHa
bpoCLS7tiOIDzKsyi1KTtjf80jSVdhAMwcfi+QehA7LWHKZgI5vze+KsY8XPq/2f9NgUA+S6YwXw
/ZeaWfDuCizYg58xVEGNPzbrL7Oif4p8kmp+QSAvjyGAccKiBbfs3Qn+hchWPWDGHSzXeophwNty
RqZFmPIuKODWfK6FLPT93kXDgmdxuCkRLPgQ9jP8QsDZYeDlHN1dIVbrfC6UeOIff4JniiOFKfE8
hYGoFf3gL9Pd53c/pbawUZIibFrVDbgHKrny/ARZ5p85d4WwzweFHYbK7WUcYtOf4HyeOhDn59Ob
kcfJkBT+xEEhyoI3BN6D1gfjdsG1r7g5+pR84OFLXY0xZRyCix8nV2hqUj2foChOKfguqR21ehQE
Ljfr0EFSvqKan4DUoCvPM8y9KsQJbadlr3/ezTrAd2r4Gad6apiXlvE3cBr+bLynQExGBDPj6q3i
izKJKoY/71jninguNqfs/cHs9/htl0AD4wMxIWf061TqEG8zux9rAaMp2zUkRuTOaBV0VZ/t8/x5
IoO9xnWA9YgompHBPHrMVy8+H/08LLB7A/KiSuU+UNbYqgbkUY0+maX6uQXsKpE0xS/+r4aFjP4H
E2c5i9Leuc5O3Uhv6TNokT5ohaFIJOfBXT48YOBAcr04cMl2Sygoamd405T5bS01DKh35tVuRaqE
fSBXkrJGaJ3n8xuhUWEDk8HPiPwWiE3pfuFh0CWscontpbq9QAyagMlwdE3PupQ3xWkSPHte/pUP
vILD56Jzima/P3gBd5AgySSQqBN/RzHFUgenY0DnA2Ofuc1a508zh6szr1JAJcS/04mcWHpJzJfN
Yv+pqGTxFUG/n7g7Gbb3z3yWBluNgfV7cKqxzLnxplKoTE+3DMeZ/4zlg9HpZhHx861QxIzc/rs1
HzJ+J9qAcnaGm5WGw/ZZaDypTdwsEeAPJiZAbv5ovxkMgUIyOZQLI63RjZCacc6rJ+patKLmkgiJ
nDKsZSr5u5hRTy1sjNV8Lqek8KuC0dC5mGd29gOpI+m0a7bwL7mWhK2YTNXiDpLWBgOGcKY3LcTv
23iQtqw9j2rRLMCYQLqdpmmf95B80qPyPW53WmhoXr9kKW9Xf1Fo/XpOc5QZObiOYAsYHr9Qofhb
cyJFGeA9logKNxq233+n2t18GHhfHTFU/xLah8YVH5rOpFMFcKtLG+Z072ythiWT2KQxc3Zz4/vu
30/5JiDfaHD82p8mem9xCWKdPejA1hx3NUYIKZySUK4Ag+8Pqj+8ON3wTWrFfn0/PyxVbiE1+8rV
gvWoloXiv+gAB8mVPmqn5TX3l/IAOd5UMzrTE1vdXeaJ2020yPXYnThAVGGLji2UskzutOC5lbLI
3zH6xv8KlhVKjs6JM9r335qLfOoOyjzverpc3rWoa54K0EcczDFqbwx5aXrFIsTJCNakz/A5pMgf
4xwSa0gS0N7/Zm/sNZFYlU8jB+/ZJX2MqpnUPmzV/xnCt6a8tCsG7qUtIAmr99xavGP5KmVDGd1/
Fsg1fnQ0e0C9NE8UPsiP8nmo7v3YgWg14GuhuU7H4pR2sUziMksk8moLLUKxpHblZHSR/Ffvcls9
uYKkkoW+O+cZSDg9vEbcvDgp0JD3RiHeNJbu/ozn+vozDlRUMoPjW7Vf0Qr2Rf+d4bmeTzjP4h+Z
VMlBAR/YcuGOKtitkGLHV3c0kh7DkoAX/e2ct24HGUVKh41X0JA7rrxUAnLqhv75Gfb23Xqcsy4Y
Rg9EtmuOIL4kaVUc3QQYeBpMGswvhEfJrmmwRp07VfHcmXEcsT4lBWsmHRt/VR8WLF89d+t419TW
9nub8uW35yY2Csn5G4EzVMFOLw6T7rKCmi+bRmNFRwsjCHO3AAHwnOR1zWueZwxFSNgrwfkvT2oL
d8xhjRwJnm5AHEcVitMJDaMnqALmn7c0mnglugajO58K5EDVjX9SPpiMswLlL+ovQ0/gsBNs2LYU
D2WyY7DJPSuh65mO39QKWSKC3AxVzJiVEWhBCLatl2R7hXgOMr8yr0ioFo4Y2CHRJAPn5aJis8X+
MXmngxp0LwUi0doJoYJEiaEG3nJf5zhhqANvquUikOLGwu/Zl8bfLn7JLtYD00tYRq/n/9ITv3HO
yocUev14Wc+E4lSzwkK3RmkZp7VoTEldZTmq204eNeLNCib4emh3M/QpqY/sJ3viXGGBjAvwkPlW
D4ghGfPOGR/I/lysDpdFuMGPCHqpUaIyg/8uQF0fYPDywPgb34BNNxeIj12h2dNabiKnyevTGFsk
/GKxixF4cwhVDBXFaugabObaxQEWtgOlVLYBxxm9Dvmmz/HKISmYzNRKuN2b5L6I4G2Ve97p+ZWu
4UGIVcQD8kJpQHtkIO2Cr6KcA0Ae5jiVp9BGpFPfzojUWAxCDVTIyBI+2BYXKCCPSioj2ZfXlAa9
5YtlhBPHdxVR6yj0nCLCi+IWhGZRqwz3+IhP7XIgYWL8YlzBn5zroFXjEmE1gd4VFi+Tkhs/v25W
ts4YqY8U74+lpd25FQv+G2+xyKeBwPDKS/yAR7oPw4sslzPd5pwoLASqEjQnqncQjCRSu7ClqA3+
+naOyvl/1RTTO7AgPmsIl/BpBk00tMuqCdMl/mOqMhq0mvExBp0rI4203x5I0inR+pAxXeV6e58z
2Gq9nR3z6kToJGw0rzo0EzeerKTj1TL+vncdUTMIfnyOJMeHhZL5VzFirIe1NcunE+uE1ybCOxfU
dbUiEkYiEvKToT8EnXRNv4LZs+A3tvustGP1HlbnKMHpBhCwv+DMNWX5Zgbw8h+CM0ykIQ57tcnP
7gP+UGc5aPheTEkUfAXDp/g3D+nc1MEbKcCMPvSkSjwoIAKyWx9wsxfCJShCJ2N6eEIrROJVQ++z
To+39q2/lz8rvzHLTceiMx3tUW8EIebEVSLXz9c4XTQXBTU0Yrx0N47Oz2FnsuE3BVUCqvMSYxCR
eZUdmei7NGNFeQBxXYNAsCwVLd3szS0hbPCJSPyUQskloRN/ClOcsVrvKDlieiizAfy9USwMX6mj
ec7z2kvOIFygeaK3cOJUIW06e25FlwrBsW2n+ymjC4zSIPBOByqj1G0rAcTbu/p1WUBu803go53A
34f4v/PCBGwa5CAPVCCTyBnJyTgHyx2arD8N+T6do7EBAsm/XqXKscG3S4r3CMCYiZlpePk1/s3Q
LFa6a4mygKL3e+49GwPezLfTGlaNbOdRxO06ZVSQsLml9HDbfKKqIhf4P7q2s1RIS/aIvwUu7Z37
xkUFx7OTYrlW2ixVA1kaBrZIhxRYhJYHJQJuRsuVPll3xFY7D7wWGtvja81OJi8hsrgeSSLvMDkM
50sHo/dpQMESL0cGNQAD4GLyo+WI7As73hjQ+VaX5vxU4LUgtmrTVwvW43AwebCkL6Fb5G/gWmS1
XE2a+muNdkPf7Cx7Er6QltZDk10my9cQf4GLPhIFZiX8q04Aay6b294BdqrhyGylt1QBF0GsDcm5
to1O/Biwhqoc+171DvUw3d0sAssxHQrNlgxt4R2ZmPx7cd8ZyMBnJewK61MWs2unuJdiUGR17RIn
+SrL+o37n1a5zXZVjKKl8PpZDQmlB+omicXRgDcAEZfOvU/iUWUPCTbruvraJDrRmEvhXtTKUUBL
r5DcN7lC6qkxfGqrRRyWcCJfVME9kGsgQKLKFd/nHziGb3k8e3CoVq1onT2isOvqYJ2ZpWajhj44
rYh71Jh4Y0SAvRmEJQqnUIDu1+CT6L1nwe7qlyIkazgrkyjD3ontUyJTQK+dzWMVrmbJsZVOccmv
Drp+lo5AnmDjvLu+0/h0+MhXkgYF2p855ythTR5SxKBeJW7sQWnFG9yPay3oXujplddgJfrzxEdA
HXig9niPnvGiRAxMUaFNJDJCVV18JiIw904Q9wF6W2nEBi1o2QL6cdybdw1mqfmRSW8Sb6VkhVgn
CFSYzOTopMhqr0AZbZAl0RyOVxSAWjlXsJQd3x0mzWUCWdBs7RuBxM1+kyrhTTp7FhC5Y8k9vacs
u7T66hnwxFIwZ64Oqq3nGxtBb+owJjiKdWAonOQ1AMVrhEzRGUdVt5MDgzX52G+XqtOQh6Szuc9v
mfxfqe7DmIrWgKpWHVi+q3tpx6+tTPUtEPBwm3m+E+i73m6SY/at7JG/aIpw88rXatbmfdJ326lj
dvumvzIzkH84DfvTS3ISfEWW4Z9kO5bJ9ojOhXE86hD+slY6enQO4qqGYRPC6GSJua4jYODLRErn
YSsmTzeEFTKw9XCrT/4mFkwmXq1lag7z3NfF+MrQyYTKCiKmB2y/FDvCXyBN6NUqkZM4lyz+Ugki
TQTg6Q0fC5YWrc0uHPCq0C65HTQcIFkVXFapN838kovaR8KP7/gYlAxFAUphGOcewFvjJ+q8eop2
B6YmbZLEy91s3dv5w4q8ejkQP+bIGwg48v/KLdjwZpQY8llo8PG8/neWELNdBxC+gPeO9cVDrLSN
h7hdntHpsvrfIN3owG4kRpy67C++Fsx7nLRbWhPXES/LafiaBXpbduJzT0/rHGoa1tugg4L8KMvp
4dmBHCDCdOAv2W8T05HaKULOm2WZMZ50F6v7XeCtSUZLtnknW2KiQALfGqci3jfkTS+nHW8YtxXF
W8H4Colp8cu/TyTbiuqecV05Nho5EFDg5ha2zuBWjiKB8KYx/p2gp4e7LYdraN4LAldQcGOE+dfn
hphuler3bRhAM61ubeUcSUB/3fTLy6Oz9RuvooBp5oDeU1dlc21Ks/WotV7wJjGIbkxdRd9susum
5YZBiVogotWr+DJ0pUNCdavjdTYBAv6xAy2k+olsMktwFa4KNZbqVSwIn3XHvSlj9j4wwBzXkYrV
cBfRYJdLIxIuhQeDWVwVve5nUFPPxwHS48sqzmJQpABcs0RkDXFbzC0JzPdl2ISS4/1Ugqq0/dV6
hAvz7TKNEwcDGeacnjELLsyWnmiXq0RsaobDzrrMdFouhmLV59bECFkHHV4d03i5EPTjLbZJR1Km
0xuu7sK1J7LzTonrDixORLBz+XgrscsOrIcmTh/Vmb58Hzp2h/h5RtylOowkfIljidG2zkaBpeBw
+v5mQ3rw/r/L92PvLCeRINs27abgjoLJrAyMCjOOZANCufXwou6sBglI0IywtXGeCGWhuLZuXFYO
EVpOUc49xgGsAMO913f4pG6KU0YdT74GdQFu3SQNu6gHYJAffIdpp8w/vkmUY4KzpuHH43iSC1e8
wxXe3KeAumRFsVQ8CfY4j7lp1G5nyoKlK2PeyPgKuSG9JHSOlYfsTXHBMLIoNalaxEy/soRGHcjl
9fcrqwwuZ8tT/5fUhSIJAGuqVTx9k8wVuCRti+jSy91eQ5a5kjvhs2T4oh6S+rqFnT7MhOp+ps1Q
oQhEXDe6Ygwbr5sXNo9mHRbNUyYTZ9v5FjemBm9OelJAH3or9JKUKZnbrtmzr9iCYxIAYnLRIZY1
U+vlo1s5WdEE7xmRhk6ClXJ3G/e0kTTgUVF4CogJ89CsILCOYaX2fEnT0WYkvcF8w3cBReThDQzu
ZGAia1JwknYkmfT+Ff9q+nzKASBs9j+RRmEWyot+dYWkMgR0gRHCWlDVXx7KM1WEEwQMJEBSjIaG
XNj64/FCQheeOZRXBoG9qoEDWRoTsjktrtrTf9H9YGb+v6BH1iLqlRepncENxo6xq7fyKcoFCUpS
OaUKf/5+6zjo6IOEZMBimVL62aHGZHDjHdDnVWS+hYQLyh27ejqIqo3glnenpMIm4lXfoFyqGVNJ
PCHB7gCE/XFCWNTLzq3xLAZosbf9dPMBSaEgVkKH4S4FYzm6UxZj5bue0pxgbiQEuSdI/3gwgBhZ
iXwLfhkYds5Ftw79CmySOo4CcKzv5l4Hb90YifHQupdMF1ds25UtqIJ/58LrCf9cm2gd6NU7TScP
O0fx+eyqpH7RDgxBhkjn75+NLW/5ulX2bLyx8iU+/RniGDuNhTkni3gGfAzOGPxJ3/vcGbA/fHnz
GynnvdqmlI926AfZQKaK4xTTb0ME5T6UsZ9jnngns4a1lbh0qBgaz0/X13yASGBL5JWV0I68V30R
0po+R9shoFppAhR8ZMddkoAXUKaI3fIXNTRtYNwqLTdYn0susDRpTXrCe23d2U0/NMGkxho+sa7O
nK/X7bKqUu6iKYfDQKfeSL4EKz4Q2gdUY7duuGgZDHkCnhCv2c55HHA8hlYzG1IzHinxwPRhUW54
XptaZodKH9EB7n8WxakqUx7nwQ88seH8oX4KGflhBKGu1ojxJsj2IRpFcAHwe6a6OHdGKPCEQjrz
wOfTT8XHIFNrRRQj216F+B9g0sYPbGDzWQADv/GInUNmvHumlyLxaA+voi5S+2J2FX/xwBR4dZaF
glUgSmsqf2lKk57VC10ae0vlWDNN+oU6g6tR6uqzkSJG5OBgCg2jbD3mLIqYaXd3oD8BnLTJDHBf
bASmDi140f6ocBbxJ6sjAb9xlM79vSyPxxY7ziU7aEJ8CV8u+O3IOYTLDsQQiLhajos01EY4Isgg
Pdj7U60Vv9qWGXQByHTuQ1TOnAwhBus/hB4vULmqT8HrDQrJPPexCJjTE5uPjvExLBraVylyxCRl
mmtmVkKtMNqOQstHBI/JDwgKZ6X5wzq/Mbn149Yl/kDLpMtt9HM3VHtLbYfGRTKn6muEf1/BHYVW
KuP1HEd7tvVUbOe1G3wjnMSKv8ArTBXxJKSMUmkaKIxzfnz5CiUShAJIepHE/qX8sAJNL+lFoXXM
RObQHhYdtcAeUSScEqaUHfOeI57YR8N7mSGtViSCwPX772gOd3AKHKL2VFAEtCmXp8Pu4xjG8zzY
zDHK/2/XkIAChchao5D0loH0aepv8Heve+FA9B3msJbboGyGdZA3k7PA1/It5lqIiI07PnFf6BRR
nE6FirUkfYWCmUR4O5FiZ47GDfHs176d8IVPku/P5yC4b0xHMxHcLHTg1D1iRf/44leWXRKjaixa
CrL0pCPyue3f38MD7cO0ItOdJjYdznOKgD7UQYqDl7OMDjptVHeEiWPZcRvs7xtdv43iMvjMy+VO
tuzOWi+HwF+3h5jI8jFwbkKZaslDjnDwCIBI3lDuxluQJzv7M0UnYyoo2oS86jFf2GrAf3ly5KBb
olB0kijLjaCKgdZAs4vZbdokLiAJZ2UR6ESGCiICxT1oG/WfiaEUAMqTPDUEqheSJyjAlJNUIoRZ
H70WTYoaAu8QSVt5kAM9IdQRCR907E4spGWAPNSi2WCpr1YYO8lSR09t4v5ULIuqYS/StB/ieoVZ
2ObZqGAt6ECGBQqEIzk51UIvKri3eHnYDxEnuA1X/dzaoWveYbWZzaZlqqiDmj/1fEILd/SR0aiL
+F1GVAPCV13gbNiEQOIiftJV5wAyeuCMMNH8sIq+3nWQmPv6oejKO+YEOAz/kTACfaclLslEGJnE
b3W8PCv8RW6LClRJR0Xk2r0QGY/scmFPFiYrVrvoNKLN89DBWhDkgqJesnFILamf4onqeuOByEbw
nFCATaJyms2V218tVcHJDd9KmfuIsHbwX+TKsFM2g4lbl7B5+CHcM93r6RO2qWGOtHCXIcVtsyWB
w0KdAJghTN7BLb8k68ELITT9anXI+dBFw+jhX0QIbvYeC9BuQ0wbPtmvk6J+MPfZmKD4lhVHAG2q
CPnqlJRQJbG1aO4AqDdZhwlegvY92vxoH6Q+PANIwSoslBIvN1UoijZJ5wKnJ7yPxVUvm7QGSBua
DU97X3rrG5ybho3gQMeGbk50X3VOLHS0B1vUJThkw5N5SYbzFJo51kUjosnEv+IlK27QJczu5k58
vuwAurlFZbGdFMIMeizjdcuPHr2Yje0vhqy05opDFaXOPwAuRAi6Bu5F8wdeMEmzMWgsCT+6JVNm
8wTfItMlbixzP71jsU8GteVKe9BHsxhpQk/Vew+pq/RLma7Oc+sxnv2lkiWEe5QJLAwgW+Qw1/qL
LM1axi+5/p/Tdy1P/Q7Hi/hdAe6mUhctbwgFm1U7kohH2iVo836r6lC0HJgtZ769yhMKBf/A1Zhk
zl7YkSaldieIkAjCZ2hNnuh517xejoddO+L42yxB40ZL01zuMCG7qq5oBHX9i2d046SMoWuU6u+t
0qtyPAjPavJ28JhCUkEtZlBxkLVwiN6dFKCHQcswLdxQdwiM4lZvtaZwzhqfcwo3AG/f7xwsPq3R
VZoazEG1YyiphY7DXT+6bgkMa24m2NHnRaiwfvtF4U+fabjKsEBrq2wGtebfH+9mE1ObGHEAxWiX
nZeUzeVvcktqC2GEJ/8emohKUirgsAu74kUnUVbsPGyjEIrBL4bMe6w3JgRJTieGjxr1tiwNZVde
dCd8pptGX0xKXf44C7SqLnwOzt3dx9p0ihUQUJGkJdcJI8vYam4ZiqQZU6TvjsvRhElqalA0k5Nr
jGwLuDL+Ac7nJRyXAE7kJ7JgPbAIZjTjeKWqztlEoTeXIVgA188GaligDSor3VTijPCfG7FNJ0yC
ynJF4uGNAnHFzCE2KSx4KnDHTgrx29KOBqzUBnlyx6lMWwt+4KywvsN8MIeDtg0TP7gLSU05uV8y
t/cTX36SXY5xgmvu9HS1NONM/Z5kc/Ag53Xzuqm40BmBTSzAZk/m4jyug04CpxgpOO4YvvwwcVBz
X5NvoVO5QgpLUk83O6LFzQhMYP285nHvu7aPZ+PWfKAv+GouhIrJz7RFwSuXkPrR2zpJTVfEmL8J
JTcOcOusv9mwItLZW/DLn/yPx5GuyjAObedjBnv6wEAuqc1BplNqaHIziUT+4ukjuxA3cvPJmieY
M4ZFnoK1+EUmdBqix+/0b6WoL+GPLTn7onENSgYYsnWWejqFbcMyY+65vdPvrfKcY/EadmRoHsm6
8hDGWF47akOXIQYCp/IZcae4JadFIIIx9uMce2NFSXAS9l3vczQ31e/mZl5rOp9Bj0qQfGip3dcC
KJr1nKMFcl7eyWiVL11s43vHz0X+d4onSpn84U/jHZaMHicqBPeuUq2/4kekWklKfXpYbtcC+eTE
8eVm2vccqrrlvAr6E0fWWbC1kVh9yqk6l1wl+UktKOvOKC79ljJTnFFQqkA68we0yqMkCYuq+NWr
CTYC9M0+LyXnxvo9LqqEP+eOk01IUNy9wzI1OBiIYIz6Rz0Wh5RSUc0PKOnVQ5SktmYjv+sYTihf
0qSO2fr2hhK+GhPgU4cMyUZvpojLwzEQPez08Yj4Y89Y6yuXfsHZX9FaNk9XDdUc7xCqqiGq3p58
CkJPOLo39REaLUaKzL9i9VdLF/UcNGW07AaHPPKSigmWwPF+1VmyzQQVmlvnvxNRgd3D2ivxd8LY
AWu0cyzUTalGU8jT10ABtZ5PbUFDKip7MwaRmW6r+tEpIqNnwUlCfz8d5HatMWmtfOOAh+zpGMPj
FnLIY9OmVMTYw34/VnycU78ARhvTQ37GBdeuw4BjtJDovDJVolfigI9Jakngwzg44NhPmTGF6+pm
IYHZCUHo2TmytPekKaH2Pj5xvfLvdC/7fJHwcIdSc00bE2QPASq6VmcbL8753q1hWS/N+QPqIRC9
5w1+SjBSv/t0+cM9ahjmsQxy2/j30PmPqzp3TDnyAPzdEVkFB4u08Wm3NGLB3zcBs8eGA3Rt/SFB
MrqmprJx2AviQhw7NrLvjsaVOsgTde7GvNU3cxuyfP3OuYiJXoerSv9TkHnYZ/MUfkixJMYjrGry
K8ZDRBcG0C1tjAkv5A/cqdmVqsQydEMVaFW2ruk99SLaEN+WHxS6RvN/C/IQZO25dV8NEG4i06wg
m8CWTQbqMSU3AtXf2l3Og62t1jSxteVbd0SxsDtivbyq4OMN9iuppMgnw+noD1J7+RkpA9BF895i
Q1lDetm/HG//9wed58LAX7Klzawv9toKYjGyAukx3Np3RQWm+t+YUvgLeZ3m3j9w7Uf1erPGLIt/
P6o94SQR9DYBuyLJsgyTk4PAGnmNr/rwApZ1L6B+qAxj9LmRqJSDDf08iSuqGxq1Zoc0d8e5C6H8
O7IYtqMO80D/bsL5Qtz3LiN4v5kCinXaL9fPLxVctIpUw+XEHFckLu0TssA2QH7ZBo/mODiRUpG/
gkJYclKvDsc7Of1pbUDBVbZ7k+SyWomVSUot7DuSTbtT84nQ8dd/WoQvKlT47iN3kYwMrNn9a+En
u7nVg+blfBF2Ck85ZZfIKDYJeZc77d/4zpsK/jKCrOvpYOkgMVlL/LFTz11fgPJ+rNwzvim38/4Y
lfP6ViRSOg5oN7r93l7QtUcT4tGFHRTwdmDgUiAm6j9T1XSeVQkKXPWmawXOa+uAIwZTkqHfuoSV
weUGVFywSsQpaojj8Lyy8SyPPu5z/kKJjKNVLK2QdNbufR1imMIQcmIuPBe+PU1oe8jm28HHuf1u
bUu/KUsEFx3a9Cz0Zby6WWHptDYyeBtnsKndRSDDa9BYvR2UIIEjYT0RaNZGU+8VUgFel5IbUoYH
r5EhkEAKWDEnMvc0YeK9VD14sr7QOGDa4E0dtBtnjY1TqqdavuCfH3lMoYZNDpOQ1ks9jwu17DM0
DbXkszU4E9P8phaUlCnMfUR5LbQcOl+2aDbfovpYZIl3JLGYhb6nHJH6vX5JNlQ7Pkx90pCzenW3
zLzW8yhyyK7BXoU1zp0vmRDzQccGUCWYN/qFjumR/2ZHjBozMChYIotAKLDKvCkPjaM4cA87HTaq
KgZCZ9TkwQAP8zxiQw7X99tnCpq7uRftYeucxaI3zLFuWrtSZCwDo4apO3h5U0e4uzRcDGV2IuFJ
CQaO8LboZ+mRgkug2dbqEzaQ4hUIVt18HMnvqog6GpAWO+rEeaoxeqLgAaOZGSjjHYZ7svybxieG
VUbOGxx8s5RAHCLdlPJO+R1lFPuUshOLKdENzkcmDodT2Fm+D3uIWBHyUEtRmke2NJ1CKWlvaAoa
WPAaCuUKW/dhwggPwHDti+9UAiCiAG4cjQ4j09175Sd8xroDbyP12zzQoDlJ1Bkg+8fRQSOLVJ99
AQijsoThfpXqPdkob2ktaLdYvGUQkjpiQN0FpIF1HJiXTArF4rYh/eKfJ+ok6UJXZ8y2RNWMkUyV
pq2zHLCgm7abyKwPXawEfHEA7ARNQAZ75dNS+dZgMBNPkpZk7XS6aZgwhzX/3aDQkZtQFey6hyhp
W0tUt4RRC13E3kqoixfF37JQ+zG5z3pntqRacHnBRrHmNO0TJzuaWPeTCPjahpQvCjuZ11SDwoQ4
D09k11PhVr3zfbHtP9oT3dEfPuHu/OALWe/DFHUWz2z28XxYQCes8GQfgD5gOAbNmnoDEjcpUnhs
KbL5+E7OOWGiMG1GAzRrLAMFbANkxBaarJLRnB4PDG4uKx0ltk+VzTMhI0IY8CHpy8MQDQjEbPqY
j6fPpPrajqjNGaOzG1tQ8tk+6/oJOJ7/t7WueiVDP0heqsjBkiQV9ptBuEWHrRKifIcQ9wwkOmR/
+iLuI+SvlGPqD1vMmYZhty+2YArpnSnRiPNWRW6+WO3P4CjyxlnAtvkwYGUB/ttbQ4PLNrBbGVYG
RbhKH4cdVUJlMm04n74Z271Q4DJU+m62pZ0Ecgn0Ws/Z7Q24KPNILlUy3NBHiKS7okbTW0RyCvIK
ADtnUz7QqNBnBkFKtZgsmqNu03zEiY0Xoj0xIm3pJAKMuOo1EyEho0mqmad39WFf5D0ScB/sk5bc
M1YdQsl7dI0LiXCs7tvn/RuG5H546/QcXIl6t5FJMfw/bLPTuu5387pNxBejpfp6sLK8OLMFmjUc
6T9BADi8iZBPmjZNm0hB3KLrxXfGlCo2cMsEE2qs+UYdqCZLECxKt8y012ufOZ43lykbkZqh6NMh
k8aAj8A/SJiYxWr9hCCp133hy0eKlzVZeTFZrOflOjCWQLOy+yk1Jp9qAnyPw+TVQd+AlNApCyND
GK6ifRSgq26/lK8Q3TyBr+GqOwYH1nFhaZEmmPXZLxdCF7w/s+dVjI4Rjr5Y0Ff8q8GUt/5Wm+vZ
xQ2LjjIyoDciVMwGpBQiSflskovr64Hr+F/qdxWL0eNBpE6LAWHDzQYH/ktSCAUsfY8QdIerp+mZ
0bZvM2Xs/WamEARd8+siq6q7WpuCvqdWD6bYAdIdPHEPVPA4fgugs1JIhrVXhm1pSv8eEZpI9Pus
kQnT2FWigPjAwjE1jHHxWIkmp/Z5dYSSzLrgJVcX+XKoVfwMjodhNQvprGtpX9cIMfrtYYs4mZKo
dC2I8OUXHy2dfNGaratq8RYScVX34tR8BNjcW8P25WFXrgFohIqH5aqD74CUGX1xpYJnfK9ZBPez
wAQ7W6kk2/iJt55egP94x7wUHSBhRp/C5yTMwAMD2OaIn5gNatCGAQL6iZ0FFsaGJl9mOfFX3Szs
vhNXDXIt+oBWzLHnmLLJ79Fwu5WQ0rMAJRc9w443tWUOP9d6JbH01iiObs2+yP975HzS7Gd5ggqf
tlsA24AzO2Du0WNnOvnKMZN/gxKH9Mi6v3leYlfNy2mf2aJgqZti3xbrmJ6+fU4QCy3KRoXK7Zao
9+grJtOW60FaMw0W2wlOdxLLzFSxqlOh7KzPIrjpd3xTxwJ7g7MxEOGvlvaiUzz1gEFJacHZUlF3
tcRv/KqM6DNumYre+851+NxFPUHylg+bk8wLlPeexaoRcVdXFcnAPOfbarTInGNVmR55838pLihi
njtN7fRVrZFG3jfXIIdYalFfim4qquixKeFLf07fTzZxjhT0alp3xnFrxboMQZxMPc9YI5hDE9ZR
S7vJ8DOzVNZ6Y3olvxpCmYicD/nEPEYq9Zs0UYic7JDu6WdTYE+eoo9F60BeJaXLJJ09Ckt+sa8H
1klnVRAZNmwWhmi5Ts99jAQiP7saByieXTQiyoxzadngX0eDvieQlkVk4zXJvG22H5+L5uI1OG3O
93BIWAAkyblEWhigPGfJ+wFwtbGNo8K6sXPfnnEX2n059eSinWgT5kH06gXM/P34NNHE7cdLTjGI
Ix10if0QZeKCneBMRnlQsI3BZ/k25aNEpdgPIdqspKK/f0q9yZsw4+I3nCONKX8DC8fvnzHadnY8
RceZ+Etx/G0osCZKeforUiQ7cNL5xxdH8p1LtnYasQkRq4Ulxf3npEXhJ8Ow7UBF3TNXhNy9cb+H
YJGEf15vIdGCMFATZ20xNj8GNY50wL8ElIIa+b8OOZX+XryJe4GChwqES30EWsduasm2DL4eBdB8
BwdHQlmMJyCjr77Xf9mLUq476+hHIX3noXQoOj4rUwJzlm/+kRANBR8bchDA5iqupSJgH0eODSPh
8R1tEtZr8r2FLo1ZJhVHR3MGS0iPilUwi4Y7FkPW6OHpIqqGma+zJiJOI4Wkv3/KQgUjjVhGCsV9
bQUwvl2+0oQqfPzisreCX948fk1QcuyRypEHw9o3/yu0Ci9vVXXu8+2Hz5pFOqT9KOFEpTlxfY5S
x710qzDmwhUAmKBpypGhHq1OnGmVY861B+rYl6cKu5A7qK3vblCjqp76NyAG4WuvArXn4PyZkeSZ
fIOBxugsm8+mHlkA4wrOleGo84bM9234GOnrT/Cnt4ZXfEvekRqwVwKuvV/nFP+/iu424GMw2M2o
SfLgokioIL1TgNXliQoPDDajc8zmuGlcqpNr+2J0r+70f63XjZtGntXFZkJ298JSRF+qXuz7JAie
aIsfFMXNK9Oh18mEJ1cblE1/rlpnrccxM8/DAxUs1ga9CbaJx5WcZxri29jvhZb3JE9qtKrnnQDM
u1c2f8XQCIivy1P6AM5TebD+zTj/TaY2/7UMw7QyCJ9j/bVWRYVlp6bI6DkYiPNg9nze7gfCsyIc
R+m28dV3iKKsq3G86JuYO9sYBMZu+Z51PKOXocfu+BpIx5Bja03QcKplYmYT3dfn2s0AN5jRRcrn
SQ3FjTrwjemZnyy3CovclsiZPam2uN97/9AnRnfNvGaxJ2cgTK7smqN5I94k0YXYXcAmMDWIp5Hf
jHRucKCrcsWQnmay9ZtA7D2xPPSp29S+k+IMmbHC9frrgIIFSBv8iXaQntRn+ur7bXr+fMSuO1Pf
cUJaU8MK1Jt7Rh/kMoqV1TrMbcth84F2UwO8viynDgWPHdZCGOQbkRbfSwgeRdiDkWcF4YzgT7MW
cgCN8dAPp9KVHqF+h6Xoe/I1LZY3cM1rVacDn69xCQxjX7Fwxdw2s0f6KRhoyvAusxuf5aYey6pB
bBCSAjqe8z5oxyrwGgWAA1IJ52FInbvYOZf/7MQvu6fbBc6Ukx+NfRoqJqMgPhQ12bHYu8DoRnb8
i8PmatYvp6wD8JyUXIJHrpAUUPuBze3JL4Yk8PVOYuNKA+vgcn82eMVriWFbn5xNH8MrOQP6HHkS
ZzutVY9yfu/UYO3eTqFtBZPTOyd6EsKsuguab2h39PtcfZqccU+2tL/eFw2mGOX/UvRZ19SlHXaR
wCZ9UzurZx8Z9j6xSLNp6HbqdY5QBfG3r9KwhVV274EcIkx3vj+TYZQxHy+zubfI1l/zpdYQtDeO
Zu/clCmdGXs0o95K2cXU+Az72TdCweY8yjv024Xv6a7fn+0eJjRHIvOskSBUkXLACcdyWvYpfyw1
f/HEnLT77Vx7qWv5oxQiSpjDL8Dlvwf56bh2b8Epz/XVSe620EeWfPBo4Gy+3MtrMGKhENc+Cufl
fEpBrnZmcropp/BKFCdrDDp0Wxuo6O/Z935I78nJ+ZPhJRCywQ0NpjDNilYzyC5G4ry8edTph63G
JG/Io6xWLyorTioaAEIoRs5HiJ/4f8MaSAbCl5a8F2lOlrBfqj8k2/wTlUqWjmSGeNFJeWowKP83
HWywpTKNDt1oSzo1oadzsf9mI4hc9b5aAhHinhLPchpMeKvr/FNyoL24cwWzyVrWhqVShzZl/FEI
4VylpIl89vWvULi/17rMK4c58QW7WCtMd/stNVdTqJKYXMhoHqlahbm69DQSTtrxtYTDFRkT08/y
MRUQRo/OJUHNAb9nJgMGjNi+x843VvNTervoKX35orwqXqhbb+/1mMqmPcIiB4DC91VUDfbH52qH
r7ynoIyhKq8Q1AbdT9PFJwys0nSvMtZ469WJ1Uu8CQjh46SkbflzI2XTCDQzzbWOenWSGajUB3g7
1pUDIN0b1jIX4QeI/Gc4HexISwYa45E8Bov1icONDwWFOpiRI1l7FrMS3fL/pgezqWOc429zxm2A
ndJTl/61+EK5eHWX4VD6CWQrsBNVoItEjY1inSWuq5hUaS68euTV524zDfe8DtJaDHAMZiHds1Zw
KcsiDovs9uUPxf3vS3wEm7PvPQr0WBZ3tCh2OjPB9yf6u5DhW46150el3Nm3wAhk/Q8wr5UmrnZU
7RkCja8xKiyuXgraN77m4ZKW2M0jXQ2sMaybUEkbBR0qZaP90ONTdnhcs1YiAkT67Yu/BDDydawn
kGdSxw0pROSvVmdP30eXsy+k3WsVVyh7vIccSVflFe9Z0Sm0i76lT6E/ftnqT7HTBmiHTYYcIhCH
Hn6GvfI4w0vXxjhZJAVEclmag4ZqrHBgxMaUSNp+2/7mMsOnzrGZmmWd4xMdvXZ88YyQKfG+eIxM
ZA7eVUv68ENImOqEDDOrvh4k1SDLJgYKQfph2t5881EgFrAR1S2DpkM9rLMPL0d5fXklssqCAZTn
SFRrwc/rGh4voUAkmq/dc+2NRlKcxniW71bl4QBHWf+yr4BPPjoJIZBOOqXAEOzAXeuJDhppqVt7
LwKwU7Ne96fmehaI69WVWnOtXkuv/Y3H8t13XgPrsctyKh7HLKbM7GJsoWjHdGDhBZyiLrKkxUQ4
+z3t9VsX5isaMmbro2OITZl9KeZU9F0kTNm7yfygvBTfB4jCOVVEYiLjA2gKuHcK9A9g8K+fTGw3
AfLfbClnDnjIepVGyKho2a3H3vDu4WExZDkRh9yM6lxJdWPkTpPbzKGEt6cll5i/elADMcfbDYc5
f+ba9q+v3bhJrC7Qj/gajfJzU+NR7IgVo9ORdYq3X63W5KhrdyIPVhS244Xz6uRfJ6vLCjLI5S6u
Yqon776Z3V+8HdBUi85uwhdrPyd/tdzLd2nPhWkZDXpLa8JjUw/9FRuQx8puMf3esVHXjGT+WKdB
FuPb9pTTC0++yCKybz09cgqbgn6Ldb6Rz2cADdQ37KiQMH2p4CBb7hu/QQw8eiDVayXlLQzlMkUa
JC2j32eBe0KNrvKBmyl/SlcA418Wzxp0lR8gT4fxSIbfNpgAvG5aXv+FU8BhqHjtWu0RA4zsGfFv
uNqfa32hSFruQyOoWuHhPaQI3zxbKf1Pfzf8VoupW76qE1b0mZz4OvyN8tbAFtDg2XL5hwcQ+JUM
u1pfzEWBqfhwkkfRE6NRVMATW/3CnjxCZ0UirXSNDl112Re7+yTQF5gpMFbfCPtBOYtJmJ8GQZoO
KcLEO3PX9XNN/GVr5BgYLqaV7NYSQbYEVIkYDkRUniBpnKVNmkkbV5vZbHba6FGX8G7rDGo3eM6T
yMkf5NFRzFphOk/+vj75gkRPi4syX2NoMWWYwVjPu68oPbYlajvB7FPoZJ7NPWYqH9OvpaJor3HN
5o6BGgJRFVoazHpa0vk8xNTX24GDMrEkvp9eddTLQGO7rLEAmP2k5b+1WgZsbOwV+d3ii3M3NAk1
O5LO8/rPdoNBWketAIYKeZcFaKQPEJDOIAsU9H5MomvdTi9H7580NSwVvico39DRSquAvj2NnxiO
9AR84Z5gMOFROmIJ87LX7R1qWQ+HPpV0zbkG3mqjllpK18WXAzW4RRbPZ9SpZ88aHTnFWj4m2DER
PucX4P9k0e4niqvjPISlWT5csgg70xQqkyljv6/RseNciE3nAAGjaLR1NceORUYPRmJNRgZ8iy7G
w7a/2MjjmKI8M8gDPEDj8ID/MVlnFDLhGVilOqusNbuANfbygG6nwbpjQheX3EC0HUmWae6sDSo9
05t8kPmamNbZl4AKeqyB2JM8gK/JV11HZ6ItGEuaOZkmcT8YsZYmTA/il02TMewqsmoMMYBh2uuE
BbGbPftqMvocV+EbnYL0U6J3eqrJ2/GrY1UjqZV4IBFqMYAiXqt9cIbDsr8VnWjxIB0UsOBN+zd4
+DvzpA1KMQfF1Qfd8PmGjNsd5t3gmx1St4fbGa6rHFgtbhFuy8HMnfnFOQwEGyOJkmI0l2BaR2aH
vvHHFQWN76GFKenESSytGark+3VaNh61aA5ephFKcIGR6SevGRHw7xuT6U2DmGRV0CJCQHiwcFFh
z5aN4IKbf12qCiSclRG4+qbRdyDlvGZioZKWXElRzZsNnRJSjNwn+4TUSDeBkstbLzxoLScm+7g+
CYkyKsXTnanRRnI4L1B2Hgvew3/ryZ9hzIwlQV6MAflHn5vdyqA7zdS/ato7QZUF5xT6898zlwAt
ypPc+fosfv8Hgk1pQ7XrzOX0gxZUeayprGi2HISVCtfDHIUSIDfs+km5cGslzG+5c3uKuhHeTVxG
/i5ajECwtgY7/715/VI5VvhLrKfRTNF036fLoh8svWgkYyhijX5h8vNxJwapEucCfOn+u6iiD7lH
AJo1FelSspAkfVA09ZW7riivzWtyowL2EyKKCs9fqpfEssgs6xoZSMTc/GnHK3RfALdZIPVLFI0x
GfkWKERy7t9hx3r/pjQPrTcAt1Pc2WJkJy9ZNEzcn6s8YO3h1x+U4e0TWZXK4fwWrVPBXQ/dfINV
gBU+VHzN2+wkcWy+zEietPI9geicXkU/Dbi4+OFK8u0I/BWcgq5A9n5yspPBKgiRCVp5jc7TrHu4
kHmmUIWdBoJGrmYFmfP0nFlVOxGEJ33gIeewtXV6eXOKLnjDQvBCGJxIWELFyhuJoM31AGa1ZPnr
st2UiByOzWX1YZzAV/qBgJ9SRDuV0uXStLV5QA1CaJ9R3KNva1gm2D4erRcxQz9cIYhe5Oormm+V
A/ksQ4cdOxkoaL3SKj+ICjKlmZE5I0gLyP1qxJQisjbjL8T1l5PlYoE49ZMBeS0gHCNu8pqDzXr1
DsKThwkueDFmmYd+bSXUDV0OQrvo5Wo8AK2BbVWz//cfdyyD49NEmIk/ModBBXmyo7hWepaAMuop
/kgo2IHec+BVesB8UELo/jRcI0UTeLhivNuGvEBR/Fm2KvMYJxFQs0KKRHAT3zgPcRtEmdnqu5Pg
ibZ7duZvgxPcBLclxdm+38zcsYn/PVEN0Mb1lk8nvB52Zxih354OYm0R7SzBtV7R16AMJ5PW2RUK
/8r/XbvGIIdD5npc8LarOHijQ0ZjZ5NfJVp72MhxVgfb3DtXvswyeYx5KqkWjYdq0mhmOWjcCU3N
KMqaqQjmOceDmPYNLXynd3UoQG0s33zYYFIR5qwQx3H8iYel5aWCV2bGB5szMvKeoYPwQBNVigKH
j1NWeK6/Ym/011ECcd3SawkW0HOt9/XmuGZXRjcVZIN8Xbjl5UQ+VSQ9a/fHjJ3wo+97JLacXIxb
5yVZR54p90I6kSEkC3kPui+QcIm+rqEaG74RvdoFDeCED276yRHj/78SylHLE0n53YNuQ+KlkTz/
EelS4ss8IXGNa44WAes1LJ2ua4dbbJJJ976Hg6vXjjQKJdufMNktdajfpVHVZt2BeR060c+siH7z
jqr5koE5a3V+ci/9czNlN+D9pVt9kFd+bPadnIuM9C+Iv5ei3NpRpXAuulOK5z21CJuM34nkYVAK
Jv1cAMR+Y3E0Ol6qn/ab+GTUOBjuakMM5+eEuNa164iYe7vRaYneHEGW+M759R3oqHsAGPAUHN+O
MDSTf4DxOGGXJH9IxGvE2zPH/hrR6tCx05OUrI0j/NN3eQdoI/oxHb9jV2q8hZDlqxUiuVk47Wv9
xZ/VdV4d4O1jx9JANygpcpoCEDlYCsuPvQRZAf4xYalzx9Yofb8YZvSj9ljTGLUo/2Zd+jSW178h
jd8uQmFjY7tqp6XhQCgzlkCPW4Sl/0HBZ16jM3HNcJWedj+6x2uSH1BODQx/WSg+SSzVOeIsMF9T
X2qZBje8wLBvshMNfWBZAd15EJ/Y2zL5N/mjoYWzhY0KgjhH3xqkgY5onqVoGFzFwWfa64Nd5Uye
pKkNL58e5HJFKnY79AnTfJmiM3U5dxojIIEuKlUTPvx0uEuhDxeWhDLmaLr6h0uRWLz7R6YO3QV9
h0jnzZ+ZLzIMSjzGGJsG6sViAefgphw/TiWvOu8VLSDSOs6SbhLKYtFkVz8nbQf6fokA88TSf0oa
R+MhzjUJ6yyZOylZgK8OsKwJEpMqcJF/wLO5j3kn12dQiMpDEvebZsQraeUhePPr44vRDlVWV1P/
b4ZRGRFB2YltlvTIOWCJ3WW8eLOP2DBhIjHYWr0ANRMubYNfi4lHxhIlfqeqZKncGprUYrBLzrn+
uzcSlT+nrIhnebxKN3gYY4IyU92dBO9yCI7kKajKQ5Rk+DaUSG4vRljqdxo52g50/mQev8poqASa
4cghBNj+lBi6XOjN5q+Vd+dVDchdoesB8gMwtfZnAlExA29o9YdpKkfd84O7laStbhe0XiUtbyPq
e0OePiz0E72xG+ntTCiAPtE6EoJhwnnl9eo16Fk3huoOn7mwB716mWlrDUBOCau/POTmnO1VRiE6
j8Yt08Q5g9efVacH83eDU5Fdlfn9dPIENcmBr1hX8UQgRMcn8Ck+4BlaaNFwJLg5Wa4/E2HdtqEu
0aQgpurod1fStCFaE1emH8sd3q8w9Zg8yURzoXkcobCWGD5/O6EpXQy5lQrqkMstLUUmNL/N1oFM
0YvwzJicxmvTWH8Z0HD7J2KbZlY2YSMAq8/4pCfbO9jPqDZAVnnLsHD/P7HISP1WW0QxcXbYTuqa
GH2ZE6An2+H+pKh+I0lGRGpreLkRPdV4CCLjQIND4G1+0thyGDSpVwabFjRlX3NPNUvOplTRIEjr
gFhv18fgaY/sMEW26uzWm/bPCVvZzH8SrhrosnAueXsIhnirxF4NduzXuv0PERLwOCTh8wXpDFlV
IWCWdB/ypxC8JGv8pff22jwqqdc+xP+kVwsHIVMfwwmeL3oNktR8ILwMcWhTtSHVcB11CDWnDPox
K0IZUh7HUAS56NlOj9377sVErKxpLi2l9ofax1pfhHWThxmIIneAPs43Sc9Bgs7dFcCh6DY4KJ/l
cbfDoEze+debBI3VyX3XkLXcrAa6CAjt2DKX+HVwDGGmiJJvU4n0+IE7AT0wLRvylANiBPXruNML
d/DzwNq0KERsR0JosePxE4b7yjqhvRgjwSKyD0V2XsRFua6yZ71O+fH0yMjz9U2biqJIFFrQLdSE
CB9uH4h2+woApJtEBWDkP5Xh1RObA4V1u9TLjutPG/aPtfsrcFM2Zjkw0MdfrdFTIE29qI7n2jlb
KK45NoP5O01p258LNAxjq5SLSWHGZuXr5CibRtQOK4dkQ71pMwLaBY4C2+eMelNwGQtPt392HBPL
AwZrC4SxJeFSYb96vPPMHritEZ7PqEIu+Yxtl/7SGvsVvL/t0MA/F60AOOKo7Dtakz6MDGi+mBL0
u73mduUUysKxBoqEXTLNIx2xQ/0XEdEveAlIFNvZ/wQB3yMEpxp3KPx1M01M8kiYPKIn4mvDPsEz
w2XO1XpObbHAqTwv1IQFFufjFWOs18dn0QtyPXfSS/4leYtwLBvzLds+gB2Y2V8o3dKHhRHajS8g
dZkMORVhMRAEeZ/JQZ2PxygU7tSwN1IYde+2z26AWyAJnicyY8FTUqPw7gAihiyejMiZC8+m0hfq
GvQuMFTx8jSK0yLAa8kn0qDxR7kLrMJ5EVIkpQBtiIS38CJJTtTdJ3Xjhpkluh1V9Btv2wglvZXa
vOpkS6NAezgqZJweWqbu+UY3V/NwQNSPMfCZICyWR8Qx54GL8uSMYg6dmy6Da1KYv3n9lS1LX62n
oaLUPKE/BxJlci4E1Qo+Pv4P212v3m7Xq1OGhkoxrnJQ9c98Y9wgcvEeHp0lS17DYrtVg9cKra9J
Aw1YchgFv7EoYw8jC+z8nX+e/Nr6UqapTyqsE3Xkjz+WYbv3DQqrdVvYm1AKcaKm0KPODxwUDVyk
IzncMKxGwrkkWAM43Ww2lvwXwW8qfMfLOXUCIF3EtFr8rCHObc0ruGXhj0ZoyQ6gkgUCUJU4k59O
5cqB++BNk8E91MO6NrA30Ym4rwIRQ4FQVcu2p71Rfqu23VFxQI2muXf2v6o5f+SnPb3RMIJMG1eR
RHZoh5RJSp/2mwwP1YIquJr0VpHSIP491NdEQg2ejWQub4Kss8XnQD371F1NvHJItdMvwZ9irS7N
Z/14g/vNf3zEUhNgEmL3ffC3RqG/y1QO+aDOyCBC/iODNUPobyB1qm3PfBbFbXK4+avnqNUJnPGm
osqRdDeZuEYmuxvgktOxm7rZdpz+eouDH3ETAWVBBvwnF4Sbue1fb+4IAtithZNTyPLjjhiY2I6/
CUbW0MWMaI5NQegZj9cd5Ru7c12IUDBn0Ax3Z8biMHxum65L0IcyT4wBXicVZtTiijW1LTVRmMqS
u3wjz10CK5Z01FqwpwwYgYcA9m42twqAcdAhiIGLGGlTkwSdxFV3yIGsSh7bN58ITVhRtn9PC/lM
i3CFs3WZWRwVfulpKz7midn8ehQmGPDfy34BKSrrkxwBndAchI+osaydcnE3XmEZXEEEdDQmNIRp
Wk47FVtju2b5SOhEUBkmcGd5bpwrnugfvctr6k5Fl3AR8FEa7iryOv+J0FTws3LwgjKuHUKDEjTp
mSYxKuixsCPIlOJdnmGw1pYJBWtsZSUGiiX6ZG/v7rc/6O0MOFAT69c4VeS5XhwgmcTz9BBuUFwg
7uhy/Rdn4yJe6yU5/OgEXBlHtPrckkN2pgJTlCWcT5tZtjBmCNEZaMepWgjp0toYUYK6B9ytsgSJ
Yfb3PHeZSE79Y8qs7Ah2Gy5wqRnHX4W9vdvJzS5xusk5Y7FElqMIoI7v4poBMn7QuVBkWbjHm0+E
kZOuSjqOpVZalQ24h17PQ69wnk8haY6bEvXqij5IrlqmMD9HGa5An+Sx3rXABPvouQJgH0HOY56F
FkG1sYkOmZ8TYsovgPBu9bzCY6BvHiK5olokvCusVLgiTgYxhkFrkuQ37ZQgMixwSQIGX6o/SUXq
cA8n7QrQWM/zOL0cQDzPMj78cYadnRL+P9xYEZwiN3c1UDOtpVvUZcTMEcvzeBI1HL13BUW9HK6x
IDOGfzlC0IcQMITqZaECyiVwPNUrg5Oall3pxbotdr7jpWLYiW4f8IgHw1vesZvH/mUyC1/vfGcm
tBqeummx2mIhyTT5Gvum17TAykyv/3EQ4qUtBbRmC1yEaCtffUZ6fmoIJZZdBmctFrJjyWaC5tWH
Y5Gpwwpc1mAam4Q/KgCg9RG/4mrhyEUzNlLkpPd6XAKK25Z7+cZAwSQKaCOZH5aadg81O+87kIUz
+u41R3e2PBJtDlkKiuwWpFgbinJ1XkFpJA4M7DCyR+7SBx+n4gFbdAbIcLsggUWoXNsa3C70hYu0
ZpBcn7uGkHWsxjLBCQgjC0ekmWn2g/WHCOIX1NdWeWnhZS/o3rl2ulz0auMzixnsz4g6Ap9O5Xqb
o+2Zu4VDL5jj4BikKBFsXP0+m/gsu9vN6SjU4ihHPe3rSYxU3RoodsJLZ56cGoBxzPwY6YZncbhv
Xj/a/FYPm8Bbe/06DQ41aXDtOk1liQUt5NUmBjMTiEeocGSJXOeD+izf2I4AwMGQE6QhUKzXGSyK
VmwGX/E7JnVh3UnVpo9D40Isq/dQv4GnA6LLWK5B+GZBDUMK8WJ2Wq8BkVDa4OwGj7m2NZJpj9jZ
DU35aZdWA1Svpy+Z30W2zJiMC5uZP8GNNn3MBokqBVJY9C9ncNJ3CiXmBcUL+xL9/+Pab9vBtONj
AbgicOiA3vxE7AQvv+HGPudbZfNvKF55yqueo4vDyAmcD8HHKIWOL4wlp79lLAoPyPTaLzPLGT1o
AsPjU7P1MBEprpHZX5ukA0xaOMGW2bNnddhvljxcQX++SUFxw5Bkv24GV4CXy0PZBu9XqjV9+c0G
r3DcWSmxzDjNvZF0N6ZrsNu4iNg8UdgYgAd6p8XoCTlxvrs5z2nDTbJ8/cBPm/+BlAayFJOkCZ6A
rQgGuyEJw38dIKgdpVHFokm23Pdmr1O3y5lZEPAbDh8SdK2875w+HD6r//H88SD0RdupjVsPjlBS
MSB+myXQ+OgCgcnec6Y7POJ9rCg6Bm9v27HmssVSUA9fSXlN5juaf7dcqKExR06v0B2vHzBGRd4m
XsAUMvwT9IyfhB6E6lDPKiP5U8eppJ0Di+lanVdEjoocgCS3Gi4ZSBUHk69OFBlTUSEUuG7sSrsC
ndRny2I9zP+6vzVKfsr+/0n0qWSL196N9vPaQJCQKT/W2jAP95pTSFfJdNvq9ABTRRDwVJey7AZq
AlVhXWp+KqTPaY6+vYQVE6fRM3xC2dGSHGMoUqx1GaTrFrQz04Tc6OJkORMkTgEadM47m7aScBy3
EjEGnissgSewAZS8HSd4LLBD4QACaRbzB06Y/KtlkgNZcyQ8mksHPyRjuO+Lz1CfZ1K1kZSrFtpQ
YzTGCijnmmFmr3ZXHCoP9qCgab2lS0try7KCr35xnKErx0Lqvk+aB4zuQjc3oJWZwyJz6qUKPCIV
weorh/y2bNZTWEBlJbtJtMDbSy/gejRHiLngc9KcMzB2HnnCrndYybWEuNkwsfgxFPZV4m9pjT8Y
z4k7/IqttHAlY8WUsJza6VyH80tfLkMmhdvroV5yDx+3VXUJYt7B2zTlxYfz4yX8VABzjyaGqJoh
OXAhWC2sU4d7b2Mb5H5Na6Aa/IicgAWoyMZncT1JgOdpshHvQ/ALiOo8FmM8jltYa9hV3IpLvL8D
KLZ9qx8ZWw4LksMk7yl9PL/vTuX6FAgf9E8HhEQ8rNXNexfRlM4J7CqBgMHNR3TkLUSKInepp6eV
KN6vlcFmXx41uOGo88MX/sPSfdBr/Kjg8iPA8069ZVMJZIFP/szU+fwji5BEWaH74sky40Q+bWbw
UmtAWNg6Qe+7WkelzWgxLCL8x2tzXajVtZTocPjfmKiuZFDm7CHl7TJonDJ2NDY/CqILKK1Y9dBu
Vij8JsQc4lONFvoIdS34dlUyHRR855J7tzwPQBH3vrjDOQ1adSCwyYTj/O2ZnjBENLFj75sCo2/P
MqXf1lGEuqXNw7h+NHB2veTwD0R7SBAUxc5Ck63VSnkyP5IS0VewUnB2B6hD7HraDA8qPHY+j07k
/lLn9NJlYg2ghiQbisQ1jYS0yn0UUvU7gk0rE1jY7VtPgqY9JgO70jnqI7roE0K+p8YH9TY++97q
kbvn6fhT/mbalLDN7wcvX52E/uJvniYAsaUea/WfR6Oh8R/9GpP/Okg9nPafmTPAHMQNLuuYL9pa
hHF2omHz7AQ73S+jzvUDegRoQLL+KlO09+TUy06PzrevgQBZgZZ/+ltx5CFk31NqwLtIVKbggwGp
RqBVvrFMTw0n2X+grSrr89RNheN20KDMydyz1QxGiV8Bxx1Mu+or7aOoql0i27tjX/PxZ2BLJWN4
rOnU4qFQyp7DW4Bu2UtmZXwgvsg/x2VH+4eoTAbwI4GwJBDfA5zWQ6oFz2TD8UB/+rhhl0Xa1k4C
klqt1mdOIEmEw+8vHMr2F26jIHfdyYCzFZyJsr3Qf30EDE8cVBgn2Dws6aW/1DEJTpneCzUnwDcF
pnKI1yrlbiDpNpjnT/Ty+AUsrJjDrwFzvsHGA+KkqzBNx397xEsdkasbRtMhx7JZQXSvNcc2bb5B
CHQu798G4b25A0Ngwd+Yar6rtYRHbgkBBbiQb/zxzp0cbIOfqvzuKAo/sLprlONF3C+x4SkP1Apr
fbt67IU3e5kEZpBbCkc4NizQFAfLaNyi5H8MD12R7Wuqk5o7o73dZfoVnnDVPNzRvwYNs7AIsRnp
ffWGFxpWm0hSWvkjQq6kLaBySamFkaH6Lm2R9w1Sl3JjBFIHLDwwHcsjO12UG1lMc6OQDh0NWFkS
3u4GugHKrqS7AdaYEx9eAGybxC9PACUUCX6o4DWTRA5Ze85OL/bGH6z6l2PR/5kxphq9zY5l31Zi
9kAKm0YBo6Ydo3dfze8Wq9lHvt2vlt627s4ECzdaAsqKobJpuwiqtAJShIcH1GW7XCYTMm7clvow
Yc9+uExdbUe8pY8KmdxITaUaTGx3CYjx7PaXYHYQkqnTv7uCJx0DfQVP1hHhvw0dsWyYzlRuIvEu
ZB1h+fIA5NZbpGEkrir24kcfkaeYdsl91QYh4MjnGPjUiSX+tCEC5F+qMUAoowR0MD0dfrOIpw7G
Ken9xDciGHqrskctOcwOJDCr2GVDglW5rs5IWlaGePGYj9xGD3Uycs4pdgs+S0Se0lX2MXM+iEow
6CXdr2Fxb0Mua6tQZBme5D6PWQ9JsLVbFSvAQzIpeiSyhURaPfdeiBiar2WIeOpN0QO/7fcIUGRs
QTmABC0NYhZGxHS7q50NhH3x/8YTMmoBVICVS1YEB3k0vQT/NwkLoD45JnJ1z6gKLkYJzd0z7ZSJ
50A796ipZy/MBhgCNpoV8YJ/HA9gtsU0Jrs6VE3s0ZUkXt0eTcmCByUFdBlt+oiPZNbegrjurint
Do7gwCXLqYQCtHQEswbpUFv6mdqThC7VzIY4BS4mlBQeCl8prt2YS529Jw47NkQgTg9WT+PIFmpp
MW5lNm6XpOIww2VUw75UwRL5W6iq+bkqQw55QXh9PtKskmC3pyTidMurXjBKD16ig144o56CTvX3
uQuv/zTZa91eWjWac2rD+YuvdUKJGZmdSpNNUsPD3Ugr0mD0ji0tP8LRr3hmkcFaqvjbBjZwoRkM
/ZTq1t6oaNiGcCFJVvg7H1OXwV1ioNnR7ej6Xx0QMdEnhQTUtaBrTOOx0rk6aVLEtzvVww6ZDdv0
z+0b8Ui+/FRQ6aqK8P13AgGmPb2tql4LvjGPzQg6iR7oBQpamYAd0wfypnBhgct6neCb8Mxxl10z
f3QmhsvK56vvbl9yVxQrOjWl9PVok9yu0nSHIFO4TwfdFGSpknUO0hX6MP06zbUFr7hBy8Q4dJlJ
LJ1qf/EA8BBOMlQQbCNH4Pb6W1FklKZ2jxBla/VlniQv9PhR9z5KozqVdsQS8LDcq0aqCcbhkq6R
JvFj7Pu/nac3c2jXryhTmsYr6gGDI6SfIhA10U2ireNpj43q0V9hsjnNNdItTwEkvrZuoo6/ai4O
xwCGrnlnXMxb+gB6AYjmXv597zgQeEc3ZXIAaT2qulo4p0gj7D4VtsNy5L3SEm7wWXYmjdEgj3II
SZfWdq6XLUt9AcuipFPLOsagjDK3oGVYqz7ea1m0hx7x0Q6T3OotKQS4O4TsJ8fbFq4QowNayJKk
vXglrEOtQmD0vG2/ys8Ka3wGNfbbjRxbZeCbOEnBYO+GCGpdL/q4902hOQ18wtV9hIiu9JjQHArk
EX+c43RpMUHVtFmS4w1fXbg7KovdLP0rgppPtI3EIlMmyZDeUfSaR8gpMSLG9DNdsi3jnxJVJ1j8
rN39ZOhUI3wKug/CYsEa9yKzi2TteoAnPOUG0QeuBnz4mDa772AYWAL2NIhwp0POioBG9YOI7o2u
jOkVHdtjmKwOaqVWJBVu+AyQ2kS50tQKXNCOmZJiO1S7bqs/OBzh0iA29DIQKnMAYrmHZ51G18GR
sYRS/2Jgsx2BABdoJ+IdE2MmBp4ZgnoFaJRQJIuHURzgkpXapUCoz6vhozbSbuWWAUSzHXK0S8Zt
YGGlBqLTP91jQ+5+pUfLB6lEqT1SOsSuhVndtq0qF7cURu2blU8YeABN7EaBETnC+WT1lbJY2uZB
SG8fhOm27pIjxi3I4bPLLEL7iJiEm9WzrVmCx/JVrEwapjo+76PDg8TbtWpDiQ1cfsS4vDYqKv9T
1F5ZiHu5nSwILV5paQ19cjLx0zcGwdPC9SJfsbH85MXgqKcb2yMDfZFNzN1UQ4rXWI1N7b77LmHi
v/KQ7FO7aDckTeJtiXXK8q+kVLBt8o6XZUja5CMRfsAsRtXf2kwZjQljetMR5L+cGaGAXATiba0Q
EuuUbGPVjYUDdBLh+oVJDcILP3lw7nUUtN4s7Ryu/kmRZNtzxo9156OdKCA8Q1XssVr/y/qej8Vl
GfVrDpsWNLPQrit8WTq/qM/7+Z9/9/m8BkUuNiPITLScwdZieBuZ0he29PJaqlraw0zxO8SqqsMV
OFxQ/TWQVgjXwMp/tl7YDE2dRA7oFBEpbHRVUkSlyz0VM8xvhXI2a9KZS26Ds02FCWX/STjnawIj
aD1KNoZFUkBSsVZxs4mXJa0xY781Kev9RTsh0HwBuz7ZVu3P5LyXztYE32BBmZqJoRFcSXzRWNT/
fc0VaZpuIHOeJokwIymAGeeJl5wIA7MoXf9XhDptLRCixEPXCvThm0yOw75QZB2aQ5ImEb2dvktA
q51UQnfYiGGIYauZ6akpTt8ITNwfwmiR+vkTxdcLiNo2D9RKHfRUofZgxKmLvsIeVNaz6yYV2ojm
ziCLFyTmxdDftL/3avqd9EiAUkypyg9GYyd7sYbUUyxjS1NWjZsiaW3j0qn95uDhgKPzkpzw1wkO
7CKq3kkUxrJvEDYlXzmBX2oUUFrYRDQM9iRKtA/eug0VCsFftz1m8Y4/ylL/iB6gzK68v30jGphh
JN5ne5Zh0S7tVi8p2vjeX9DYfbRwAJAsp4foAJqSRIExkvRPonwKNaCtvi8XusoUb7pagNqCp6c0
67oCq7AtilBE1Un4GS0zHwI/3zWE60G5Y6AX53Fmesusrw6RH6COqdI22k4BeuYhKMM5ZfidVF8Y
dx1Pot8aLR852xy61j50cg3dC23iduutA/qazKI/oXiGUu84J0QMSgoze/CVnflDfyeh6KvkNLDU
V/Qd2ELtNFsDb61C8PCE90+c68txSHRKdp6+5c16Y87lsXg92BdkRzeRxWqnD+wu2XIzI+05eTZC
jVyvU9mrBQeR6nm4rWgoj1VCpw/fBHyclQG1OZ1GpNpD3NT65mPY3GkW0TM2MzF9NaHSGLcFAULG
8WBkDIG8RNDzYGj92tEVq/swbY3KV/u9S89xBCk1EV4kNHMlqC63cBu7PyG8X7UDWAeRi5yin/Dj
UsMzRpTHLTnbN+8JPIQrQrYz9EUxkPy/T1GRzhLpKBifp5VkeDjx+8MVdudijjMyX0eCnRyixxJF
3t2RhwYLqzUwqDITrBCZLmJRHFslmF/KUYBkbU5cVV8VIoRgYzTx0iJqCwhsUVX3G5Y/kI6wFS1E
e9hrDoEout5CcDKlYnHPTOJKIbI4iTCtM2GV4mM/jEit8AqezyA4s1h6eFVydUz/VWa+JnLeuDyS
sJJXWFbYgywNSKUqcAgowadhS/3Oo3w9E7x9hUOpHsZTqfhaa86bKx+0yiTKO+u/hd72eTGBHa1k
ym4FOaM0iXH6meMxWGl9ZDYPRiymCwFXk5F0Yhuvl7fo28KILhI6E4MQqjyK877mCU/U/Ss9k6W5
sObXedzuJQ8HsIi/20zuT7TxW4lWMzzq8RKWn58CEqzifU5J523EchhQRJAW8IBi3QaZdr9EB2Bf
6CbFxwc8l3Z7mHw4SGJ1mWDDDFjSjPbWMHek7FZwokT/FTqXBSqcfcYvV9c7zDG0kXXfdePuUSg2
KflYtNFMw8bD9MOrDGWHXmS7CldILWB9DVJD/xryBcxnw2ZD2l33ws8MuPu/4XJnU1WsYihTEfEX
S67yPl4ebAtf/hwRsBDL5LoUy+h993kl8479+1FQwE35WpVYLjQKRIjVi+iihLqAYsxWtgQ0Wuav
3UlBQmaBxNK825FYQgxMCcyWrjCpnnKcFqzseO3gqNSWn58ZQCU0wclHnZ57CJsL3FWC3Go953Fj
e2EZNgz8GzKE2jgK7FEAzmE57toUuPT9vYYevcb77bJnkSl7TgSfepsIbFbWuh1CdXNEt4T74VE9
nvU/RBM6VBVOZeIUZ43K9dwBl5PrAx4fg4DPhRq2enylSL999Mo15l9Wo9+ZYrtJJQ1logVhfh0M
6Dbum6KCk9K4jcAU+TcmZR2bAKF9W6xjeWKiEmmP7u4bhD3kQYbLy3IAmLy/WMPGTorupcqr2FYP
0cEs2ME94l5v7K7itSajN4DWxJ/6aDdqLgZhk640H+zNRgo55IL7HQZv99qg+yQgA658iTa70psU
OYmsC92X5vt64u9eqaqDE4Mhsp+UBLY0mdbgLSqrkWQjzWExQXTvXW89TmTiXM6M1TuZHUnPxRGw
kvf01uBUlj5hDWPThNMhoA4RdQuuVVJTjFIhJUzfbQ0ueXCHjqx0/0Kn8hF9IEJ/kgmXu/ouO0xX
y/etYuSkV1JDXEVuBxSsPvw7/M1gmjJSnV8ufqCpWyZU+sH6BWXIq0y8ZNgkTk69XxlPFzENtlc5
vQysaCIf/ak1e2cd500VDj8JXcmdhEsoABHydbcVvtgZrPxZZTF0qBoSHFuqbxY3k208omCocSc5
ONLyZCor/YuxuiXvHzGse02nIHKCoSHmYrSfLbhsVi/LDLq3wbsE/26LHS2UdPP/FqLJlICrpKNe
eJMZzloH5ZNuX9/gGJNQI8jLclaZ9Epi4zHEXhE9YWzERAIhk0wIQJdpdnylHPM5r5Ikerm2OgCZ
2HGJpXXlWEyCDvD/qO0r8gGqDoR004c3Te1meipnDYOYwWm82TV7NKGRoTaikZgDU/uqD8YeOy48
KV0o9rlNYd1GFPhfAs+8pS/ooGJgvhx0myqsxwgOTvgnK+USC4SIFwwmm088JdSe26Jzs8El6AOf
s2wTY0rHjYCeNduTjVS7LXu79V0odjPqUvnzgB7CaK05SqI+UC2uL9G/ImdmgqBjSHYlkqzDykrm
yal7kiAHOweH8bJsI/+AjGPPUPl/RZdGo5Tul62rDeO820Jjw3JjNW4kBolWGXc4MUFXfQInXD2D
up5bhWSNHX8hVkmPkmZRr+xM98kQduS6yt5kwGNhp7Cm/6mAA7ajKcZR5UMiU6kfswrTJnmy3xOV
d5hC5K0JMiaP4zCskySIp4ksv5nrc3o+I+7unUkhjF6hXfC0VnA/oYgu7Ig1r7EHUF7OPWKuy/QX
dNNcGUA8fQ+c4c7K+IgKx5ICCbREx3AAl/Y4TTl4VdFbxtK1+XlIsTn8Sy0KCmgDFQNUIoQN6pSR
QQWESFj33rk6V3gObRhrK+BtL0KAvxyN1JEdMviDLEjPe05sKjUzSoBb5XJikan4MycgF8cjKtwA
ClKrkB9E+PwqBahp2y3lxClXzZ2lkiT5bBL/CYw+W2rchP0sdbkh2DSKnI50PHNJ0q9AghnZPWAl
UR1el+qhY3bD40UsKhhgkY8E+KBadInm+j++a15YWenX5uZTVsJT232kebKKTBq2zDbroeZiHtWC
jVNbCLxAvmAL6jwl6XIlws/H6SBTT5I3l7xrGrs+/SBmCXym2I9N/oPeHDzSkTpR3sKyB7ODX1zp
ClS9Pu2ygW3IuyI0UrTSK/eAzYC2o1JpU3gnEJlZyIDxPsJvywlaUd5wkmdSLU2kv6ac7f6kmImp
92mibqAREm76BUWjXBL9og5EHpy7OVYiNr0fuFQBfcx4ca7tfnp9nUezor3iprmMirxitZ9pQwVG
U6jCG3Zg1iY5llIahIyZI91OKWdy2PnrVUHL6IDrc46KKro8jwjXdjafWai5vs0vc9K3WIeI2gj/
UerojBZIaxsOjFAggwrIfMjfTB46AnR2YKJXRaP0OvpqsKPlrsHdjpeS1+HKIF7tG79ohhKGsH/m
lkc84vvsoq+3PZh5lvas8MAyc5Mx5IhF1Lr5zv3MOjYehGzkIuKalhEhZ25rdl1a615WUyqGS/Ev
UqpPp62stnbf3Y/A17qBcv7kMRA+C9MkTvPu6EMICJ0SGtmolqkRlmD+493apNAam7edNF1xMKf2
3YsCz2FVkyuNFRPLpburcb7isW/OMBB4cugjIpqMPTVkeFW/UM9eXoJglDwKwM4GiRoviArb73C9
d25QJ3pnQKG5xYbwWyvzjxtkWcXCE1v8eAxujX4XR9FLyBc2zcGIVNG55CJcYJYyr7kWRlf06MaY
xUFDbj8To79dW0NPDKiUf/y2GMp0hDHzgiyjf2wlHu71Hqo/njrueABlkzKM0oFmepRdtsxcDdVn
5x+XHEMeYZxhACGzB+051+R1oq9Vue5Kbvbsq9Mu26hfQa6f9p6tZDp4o02/ko4KV4vNEzoMG71s
w2lDMBKoRf4ClFK1675nO1XmB1iCB+l2eX8m83GzaClXL95WQ+J6p7ZY7uNXdGb0XDeYITYlhjvZ
HB/oj2lg9OGpnyNqgQXB1nItG125Q+n5naF2f3sjgtByxzTeHV43wgZQLMvZjZpDKyU8S/Ara+bf
39YqsJcAq60ArgQdSLX+WqQK5RcVl5aWwWg9SULxkYoNqMJ9F3ipF/Hw2OrnFYIv/CCbMxl2Lebz
lejcpdVzsXjJ7tyI5KyAHbr61O6uJ5lO/JeTLXcsA7itG8hW8PXgjzl75K25e+UEqILar6wPsoQ2
O1oIXO13fOpRTY3GoknHI0UvdgXinMn58C45Dk2XciGY1O13J+raKkSbEe967P0lbqamxsOoWpBz
pVh3dsrFG7hAVCy58KBgTuTOikiNhxD1YJ6ysYm9lQSM/9Zdow6PZXyLMKCz6aLqfSjZdM8SB8wu
h090AxPdO9yAePbqjWzmCVbuyKRxzcZLUxKI/+1HK8rzYSetMGChjg3rUtlckV+aZ/Z5NzAzPQFE
Ae9/CtC2oBoa/i/5pfhlW3z+AFY6+6vCBVSbvQq89a3eBxwZeE3XqD/Q0/+WARNI+kub3B9k7nLS
W4O9RHFLbam4zVZedHcXjKT1mKXKuKjgb4AbVuH+u8cISVF3BItriIgWw+X1DOQkQj/++bS5hyGE
AyY1Rf2Lz7EBEhmSo9akYh5kPLumGeIt75hk6tyIlkb2hqN7OZZK8uGqRGbKKtVa5HufukqMiUEY
ISEq6GU0ziBJZYUKYqKpqOP7eNt2Eyfd0MKO8yy3EmRzToiQZXMF9VnLxm2nj07Y6G7DMV3lQyyD
Qr/42HU3+5JIbhkKwIOLUzsOd9JEFEpVpNminp+xfc4C0gjbl9r9F8Q8T8HsBaPUWsj7H5SzXROA
3E/vYaXJUajGN/tRHzq6jow93nTYCiO/SonNVdZ5mF4reLL/yHLLmlS+H/aAT9c6wQwDA3cbg98b
6kly74OllWElkNXGmJOK1CAzbE2CnrPgk93yg9YZNr0xWbPLuqv/Nsi/qunGF2JM0C3CTyakwxIl
p3f+YMWiXQBW9ztuVtHE4Jmvw1q9wH95QSJwj4BxQx+nTmL5CqUn7Pyg9Ky5t5rqLZ7ohdgFoGd5
YndwgZkTMGqmcQmTGPLC71ZYV8n9tp7r64mnF4J+qtQNH/186fTkzw7H3lX3ZmrmlmcM9vRvEg2V
Idlx1KsSUNTgq7I71iexunYqOa+E/6fSL2+PgcxkSMAH2m0vfA0U7YH/4+F1Ida4BNT/pMB8C5Aw
wx6fCamVUBhnL1KDYvfMW+SyRieCf0qjh8l7fr86o6eQRWyjF0il5aeNbRRxEjwXffKUpAGIzuY8
m0mFl2LrL54aa5qWscNFa/FVqBCZPSaxVqeXmF4ZOdNLYkB1TJ68PezhIHaF1mQh1lLi4Qh9eB9l
rIyHfl4vKaDnySUC9EbEA6/ZX7t1co9W9rIQOcYvjqKfv9ScwzDNeSgJdDlDU5bsdVMTnDR/NI1s
Cr0GDNaq+SK4JnnHMxywLOqokUwqE1wXU6+UL5ihlswSL7qKGAFWsrPcGV/MVCavofUrlVsx48Ol
gwpNnwNj9o/7Bu35pEwsg6KpEpvLkmPz8EpFvzps0GDk0VfPnqhttievOkXFC3Ef+sW/KGNdcWmL
xE8dcjLoGmxmfJQT6L05igUjhHagD/DpZQXBKkKXVqxn/dt83dg9js+5zJUvuhZIoFrMTLPKqIr8
FOFurE4wvD6NaMxSEOJUIhmk74U75py8aLheEarc1Vpuwj1kzYr9n1vQu9v/6jS1XMnSSMqQ78pi
iaGSufYGAVP7vA3K8DFvacqTgEH12azY1TUoGFiVY14YS0uAstul6+PCOq3bc3W5nYPyMZobAZPX
LMJfMqwWNHX4QTq1T9xSSqRMw5uRxzJlPNLYCX1fJnTsXfF4KKPc9zDJttzW8l9O003WFMUOwRH1
+jNV9Qsqjj9f+6ZreAiQue5BEqYJGpvyPhEoxUdCNhzRacFEj+dKcFiwYLro/W8Gc3WWxobXpwRZ
705yzIcQMBGwJ7zxlQmhu+7VKPyn7ebjwEr3nJ1kNX2Vwrik1gZ6LFtgNTJTwAJIKN2smMiFaiDy
enb4RM7xluNep4LJrKp0su8wGpZQPTWlC3ntXFpV/SZ9qZmLXRPLLwaFlQAuAIGdcaHe5tkATKK1
S98INK67qXRn/W/8HRDlE4Df0CL6fSs+MveCF1naBGBIIdIGoOINrC+tWc4HGak5SIkhKoawixhy
r7tOxjIjp9MnPmlaFlr6l1pA9BwUDyY4+vJybQk0MEPY42d9cfdCQL9UQhzfc7Md/zPlcvYn//WA
zOy/sLcpp5iYpD90VWV5kZjlJgXaEYfzUu7omiKzcxGHGigjN3a0B3bmDsrjZqbq+GksiqyTgz1d
QkneGheAE+zE5jjraV3bL62aeg4yu/2Idj48zpWjU3CE0Pi8auOX3/wHmBjSiKxQdh09X2R5pHR2
Cn3PLjfHJdlyy7iqpFrRRGB5OD/T/vKhRaXJ8WTFAVhjNfIae2r0tqp4JIfp09+mw3t9v5YN+jxB
jtQEe6LAbYU3grvO6DJ2FTrLo+0m7ws9x7ld5WRNuNX25dEeg6n01UKIYgI2DvjKe5PAIBj5L2D5
O13DFG1ZETIuIbOvLEMKt5fxaSYX183gxvrz5+TiqUIoELmP3dmLjCtKE+wL/glIr+7joGMEf8Kt
t9eDKenkOeX0IN59obEQADeQVye+pOGzVObhYniLcKLiQPQrD/uZ4ZOlrjRm7I5S/bTeocDQGyqZ
mAhOcLpSxfmxKVtNLpAW6RjkxW1YM9QUfSjrbeyUf77M0otlPdhwD1vCTilIhYOKsYCCsDQp9X0H
Oo4CY7ifsxw9ARFRziEU9eLVVaaI7LqXKsEk8bH6QYp/l8YPzFQc8tGZMSAEG1X2btphECpqTE9j
QYTZSIg6MomHj5X/X/FGbQthoDAxUTqYqKX81lnD4vLBC9g+wgO987TVE8QV08fsG5xEg1Rydfh9
aLZOwdRfcVNScCQ0YTog59//OXMPO+nWHIZ/aXIdViCvFORfc68s9EiwHr1NmO8sRWcNGx7pHUav
fM1m/R5j55a88q7kag3QppNnjOYeKfldm5VCF3BhtlbMyqOv5siRXEeNPN+GpJJRJ1mtm5FgszyN
rWhceg+HU9IxGxZsEQC+reJQSN7OoeAUNUBj0PZIKetwKmxfLZwnWGdnUmmkXOVNwA32I1G9p9cD
hb3LCfoRgAtZ15Y9a1NzF7BH3qihwlNrUt2FaXq3caUfgoN0PTnZtzYC56Dhpz7F9rK5Dct0kbk7
IVvZgnB+M4QohTtW0LPMXfClExmrRaW1neXH1MX3SvQMNts9Xcx2M/q3yinKEey46pQuSU+0tPKM
nOZjdoWrNO7YpbLTwqkKQVaax8+RWxpRaN9NBHvlpOpYcBRihBaaui4gtTCplMxlcKFYBZxaQK9D
j5wiNT7FQLAoZes7nUowIun/Mr4oPVMQAczt+5Wbo0dqA65oydyoorj7St70PYM1RoTNCwmDZ3OD
s/DLg27ThRIG8wfNo6QHFfcSZGyA9ZDMf8FxsjbdjZNeQHmp9OQKe8zuQgmkfUZ1vMbqLKhhjrDp
eRGKXUuVZaZZ1v7sJ3hGy6Z1Dy/67D3wMpDZOaQRxPcNqpKS/4zIiUSkvyaKcoG1ZjMtItPFUU9l
LJF/RkfeYMQs0zUps26yhNyLvUOXdMr3RE7/Zu/aVE8B9aYagAPX40DWmZyBEjKGzQtcYyMoVm11
CmInQo+45GRcEhHkRgt0zODYovucYSujDfnQH9x8TLZccD+BiAYVpW+NzKLWfeFKPjizdN8kCn0o
XAjTHbsJDbjmqNS93a1wf9mRFHFA1RPfNVLh85ZUMNvmxbuDCVCdTcDpioZCuOLweMROKSwKtjJ4
pVqck545MTecYNgI2IKaCJLKSDsu4xH2LmSKTk1JY1QdL4BaDpr7ALT0PrtkbowE9UGURF9VL7+Z
WXlPzQX2X3T5GgB9ez2WHy22HePeexabXztM8ih1Tr3jQATf7BdpcLT+MwEXXVXoh0A+n3VYmvoi
SXD2iaifyxdUD9Y5x9cDdpCJr7IzYAY+2Tx/NY6Yu/cuiw9wgtOxJAcUhjEj0BTufsaWBzN9ZJbG
F1jVY5CB1dcmLhmKxIuVa3+vqWB8DXyyiA+/DjfJjOvD33/+wdGa7i/On8doua12XFi3aXMpZyt/
IPD/c3Ssr8kh0WsmQsH5PxgeJ/01KnxpOQVTi9Kjf4vdKEd9NOTflARwQgvkr6fG3U8iOv/F2nzL
g+L7+3whfDFnlneavseTIG47j3FYGJJWr1qHksr9z7Phx2H9IStNv2ontQrBYBl5Bjj9Xf58Nf1g
dA4ciJc8S4gvy0ZSY2bW+QJVkDg52kzJWgrm2XRtLzgYWpkCncChC3OI16SYFYJC25J2rms2+GsR
2Q+sfK6yDpRUiV+frp1k4kjuq0R3RVo7f4ODpPvLsn8tENgN3Kszpg0XEE0tNoJNebDe2rdQUbn0
Azz9IbuHucs3eSzz9bvA8nEG4QwCU8N+FuTYDoPpd/5I6Srja27JiJjgaYX5LMvHfc3u349vPYys
RZARbZpMYjVqZC0uwf4vbZ4FdOcXO+LIoHzOpkRuQip9pDy2H+PEcIXWLTTh9cFsioG/B7iI2yK0
33kGEWNpEpDOVKhP8YedtaD0Pu20QPgvmOwcI8HCDGYK0VfONfs3yIK+ptnWepboQe1FQDJtZZSO
dkHcZs3w7Ybe2dG3Uh/Ll2JkkUzlcB75la/dy1VIN/At8qMOPk9/guCyOxehQopRgxdBCo0ezeRK
DJkqmUTOVH0sUT8A1npMeihTE15GgvxaxII7+IL7BC2K+dNVrAloJLZL6r9GCOlz33y9QieYP8nQ
/wJoWJYfMe4hsJXzST8BPVksN5G/SqhqbcepU/5VfrguVDBuH9Qekp7QRKj1XEMIRod+3eztta/b
B1XC/fAtQjw7nSaCIX618PwjQ7eKYXL0Yl/MFpwRnVcxCtMCOC73PCUgaYKqUYlH9GgmONNLbMKY
6tVxEocFnwUApWqReWdJ6rRFP1R4HQsEvHxc3NxwYmeFe3ePZMbit0rg/wAeti6l/qOxJo4a+0dQ
QCnX92yKLqWL2SuhpUCidPvX6snJc0CoknckPpiW8qvSBC3njrYOhlQKSzSQTtWMy22cPXfGlYCD
a5Qy9ylxEfOhkkpSdSZVZEfYjohL4P+cvYI5pK8r595d7szAUAJD52I8ArzxbhMDkL9XQzfGneWw
xmv/WQOYZ3o9UK1osAeHTrH7bNm9mh4GxFzYrsA6L4ru1BVPwm4nC7Y2bgAw1ibf7yslxiqXnqNR
WqQJQnABs6SAi2/WsPQV6osmP1x3db1DG3X+DaN9ipQ/rfCSbMvc486X8AsWHu/IoNPYJJe9IrWs
EgDcDXkaD97bZslit4Aa5eUk7UY1PAqXDi57bAG+yCXw4EeQ46DlP5aijJp200Mn81e2d/fGJdzW
P3/4Ni59C7yTms9scTwQ1RjY5JEstfcXFZby7i1KUiqfJVJGQ729SVVWpqxsggqWqaTQ/ss03Fxi
P0wWd2Z/yGgiaSw+h6UbF8tHFVm38BpcEKA2OpvbUIXzGOgZQyn4fbwTIFDcs1b1m+KfkX7DTxgr
BrcG3KjM7FCPAzEtG2XtMfQj1ASw+GaZgRlz/yK+fGL50t14xr4bXwpLnxpgl9HxCvfbBTiDFY/k
bcAr8NButh/+rmR9z8WyIhuxLAxg+xrB3GbIbpcMgy2wWKlYN0DjzOU3I+G5jtnEm6TdFsontbP6
SfOfFngcuQlNej9Skl0IaTDTssRzTI/SxNc9ljnVLQOkdHN5qdXUCCNRi7r+MUi/1kWzXWPtpzWo
8p5sHFMymZKI6Esp56B6o2KU+zqKhkKWuV0i0UBoTx9hsIE5zcWs2pP1zhXQr8cPEtCrbFJVnLk7
RMi8L1+IM6k4Q3XAcogtjtaKO65LmwHPVnEDdv0Dw3JNkEDj57cr3F4pvR95+RkJC+gi4neGOqVk
UYVANkmj+TC+qRSvB9A7SRnRLmmILwFzsRnQqF81VEtRPPSGSOySwzOoY7zEWmz50+i96QKq7Vsx
G2tISI0wg4qlcYvaTtHqrsdmRlrjpVfghzWAj9IvdL0gifcVG+JYn3yMEbqJeI+o3t/7/Gflu1bY
XVNcjoebDPERWgMwyigewCD8sJwnJ7o7B61aWNJjl+amqyK2nG+I5imareuB+xNwSO1oh3RIHoPN
s719ZHaCHgMw+yTk9LdkYzHqVJ+werYCfuLOWDw1aeTj01PAl5jRHT9AIIw9oWCEKhSEyf1MpXpH
JmN7Wj7J016StMu/W3CSc4LHzqVllWigSgC4MNzTTcKoOOnNfYMSWxGQnFanWCJC8XJ1YfyLjnCJ
BReGVAduviGaMYD9JXeuS24ru29bKYlKe/o23z3wMgzWEzpziUHm0I1IjbDpXNB9sCUcELxTn/8K
NjdrmR/kcq4i9okmfhC4fYLtE4EkpJx7d55+qImCs+cmtyW75djV3ryUVnFlO+3SINdtugqhb0IN
i2hM9h4JdhskDMB++60XBWTBeXptpb6pbGReMWw5AdCnGEc5mmq9h/x5qOzSLCc30rE1t0n3U0jR
SgeeeFapWm3+9b8M6vtmEuJDhpc2hB/WiDuGfd51SuBEdLmqWXdPJZD4dk2mQqti5rkSw/a2b0r5
3I1FhNeql1i7asOy3KMJvn8ul5zvJP1GsKnkbaFuYzsJGXwYlqGrejga9BJU4lMaij+lAoeSQtQS
zhuB6R+QWXSVXq82bXeYVSz5bdBsbS05YUb7ur7VBlcOijMKuuytbEcWNdDsm2FWZsG3vuwi/keg
WGZ6PLOZtT2E2J6xrOb1mtRrgpBMoicigjW5gTUllJbk5Vkf92robE3yNtjLOzZLgcUNxhmXzUs2
czlDYpCBVbELZ8/blHaqDxVgsHdZBqAwxXoEYJxoSeCBQm71uS6GDk7FoJ7oFtGF1PdbiBdKVWQA
s76w5w8vL9VEy+r6tkY5JQxkxfkfr440JGDBoUO2411Lo4M9JcQYEIcP9yq4HPlaWVUJdOX9yt9/
MaLYOmv0LyeKyZwI1R+Vw616FSiMZr/62wZYixgBFSNuv7BUBTcH5BMJ21Ng/yugpqwKU/NCtlsO
H4j8oHDRDL33vufaqlbsZg+8Z/FNH7x1jXSo7D9Ha02LutUznMV7yMK01ZYp2QTYo1q5c5Lkz4/b
KbaVDoRpLyWf0xgOrD+D8jxtEk5KJ211lbVoHlyjWN3p1yyiSTAa/HTS/WE7a7SfN9F3LDUt8aEP
qEuclYbxt6gJdEfuARAwZDRNHJ93v1vtw/eMiZzGoMjjGfaN+fah0wRLy/BW780LVpbVJxOzRwJ/
Vhdz1zDqjKzKzB6HmyxOa0p4RrWiPKo7jHekB5glS3q7h3c16kd+4ayKR0gsIlcTjfx+9K98sVlw
j8iv74mWTDbGwAI1gOKAypIzmTGhip3fEIeLfG5Tqy6+C6ULII3mtF0/j5x909+26RWb5iMrBNfv
xxaY7isQj0Vh9rOUkS3wnL6azW5uDlTCxSkWY9jw0SKtaTBzxOyECY6pY8Voir2bn1tMfFN6CxPd
a4n0fYTwki4Z58b8VRnYt7dPTj8yIZ+lvUwSJilEDnI0U98XrbDPxg6cyfXXYxDzgCw9ZeIJ+AvE
s0WD1cY8vJawBL/gNqWJI1C+diKIHnr59Oo7TB5pELcvWRQXTeNdqC7gRjfDK29YznQ3A5yBoZQ4
/D4r5ipKPAiYGoYTrHk/oaLHawigJF0W83/PNhV0BIRlIdR/iOQMuxnU3dRYFOWAx0AfIX+vnEB5
s3t2IfiRU1MTF1xtL1nvifYh8hfcv/uWrdsiD5do2K2HxnpChY/wrCJnBp2oc6kbu+UDWvVttCBj
ijqht5NljcegLFK5zL4DRGINtpwzRonlrdrAdJ9evlPZ2T79FpKU60ibCjAbNNyrrHLa8lNUHlea
YJlG2t/QLbqFHRufkHZWcqi1E2fO2TXyP2axrqSSP9T/oN4cwQvGz+PV+nHo0/Pw03svkIwtMNNT
NzqnAMw6iJ0zK5jSElmweVPnFzbIqRYvAfnQnAupOQgeLOmAAFkYL+14LYUTmtkSJM9JzWHyULOW
KiUj9IC3KlKgrcKOVN1QCg/Iv3vkCzLmgEZpWvRjp2L9BJ8jsTf7rIpz1UJGo0eKBiTLCxcMIUhr
3p37RnhdaUf/GUNlaoKLEDjfKLzvvveFdAzyYIrwcxbaqftF25ZsjFqclkRWuNIkDST/SKSggrxw
YFuV/BXAro60ooMTfs6sVBqbADpa6VtnvIcNTfJ0q6dG+XRk0QjLYUVjeguNyDQrdU9CMM1G1Ul5
SkzD7vb0t1zsPekB1navXqaAdNf6VW+YPHza8dne1UAZfzSD+lIKs91psP4Qb+rlzejCQj/ejfC3
o/AvdTrp4KAb/xo8yvmCjwkPJVvgMhInh68kMV66YF5ewqg15TQB9+RddylaVExp2oGfqN2Ldd51
T2GhBx9+0Vi1SjnulgIqjaNeY4c6O7pRmRFtZN69tQi13JvEcvQ4HQeySvU6oUC4X2zf7XTqoedL
FDKlizg7tt20kAiMAFFlz0LRXIljmO3KtqbowyuxoMNwiSGjduhihHKLP5TTk/iaE5WxX7e9rkli
rNVWt1ddl73sxhVmBEzjE5zkQ9CBmtZyChQsRBKw6ud4uFeAAkmcG55PQxbqA+pvXHD7hqFXE5yC
Q1s0jb0vW73+lp3/nxV555zulS/LWCw4OukLEO4lvWZpdJk6LIFV4QJCKVg2oY0HaMvMk6n3aOB3
OeV9WrhWZ8hREm9vTupjdOz2N99eg68i2F4plaGzYPryXKQreWseVRG6dHEf0ANjmKXWM3g5fnhM
PfE9wXy2wZeEdqyuXsVsf2CDVaxpYYQxJyDJaOp/o9qVhx+vPiiaHvYCCGEPVSJksXj9bSD8U3cB
22jBuPndWlhyqp2uWZgHaPKlDLend6e6C7pGFVLXyBmHue4RbilI4xApvp+JYfOzgOGdOialuQas
3ccoewXgBEg7TyyHv8TM82MbyXXDnoGZgRKKpRIV9x8QSGPqUvrPAd/4phcdLJ2Q3Wf2jj/N+08l
fwTGBgqXJd17wqVMJKipXN7CahPxPuxacPrB8WM8hQ25a0U4uv954tw7cIP1AfgyOwSr48yNNfRb
x6FU0NMaeADP3Jt31z8NHhmaKpKaPksOXZLv6x7q8j9UwB/txqG+kptIfTERdIru1Tw/DfuR2uor
lugeCZPo/kcP4GiSqHD6XwrlcJzQPhGwInJPV3ngC7H8GmNKa4s3tugHBWepaV+XU7PmRbisjjEx
R5EbWCOen5txH0xUzo8OGUN2eRawI/9UoCM+OrZkEUx2uiUqkC+yjo1eW7HrmCiImLAaKlyixXUK
5DbsWHGnUb9QTJ3V26OOxbLla4BTbgthvVHV4LzbvKuSTJpfAAd9ejeFeTy5dOQbSJgNhCgKC4q4
+WeikGB3wYOazyTUoIjpkItDYSZd1fYavQNB0K/mBp4kG/LPBD1rwAzNG8ZC0c7q+J6HYLu+PoRZ
NmptjGHkyfduj3rS12NQZ/CuJECRqwr740H33K1kKu9uAnhNJzIUCI1I025aDuU+gibfbOiswi4Q
xFIIGos4Joc3V2bbwAiZ4ehGBZAT8SgvX3oJnu7AWTpcyFSX5kqkTGMSLJO3pVQhGtpzYiFoRgwJ
PXBnBJL9JCyTKiMFcojJZQBiufE+D+Rpw6aNDm1J7tWihaR1e9mx07v6pipL69MRHwIm9YdWMS2k
FqAvUcQQLZ4HuAdhb70BWrHOTqTTnRd1xTi7jKlPZlxnA6xKi2nhZinWiV9mY/AqRF4ojWNvOD3E
8HGA3TwnzxbhcEmjYVO2PfjczYpZd8yO8tL4hdgln4+JOLEItWTDhtjRITDA/uJa4xAGYhoSXrW4
rC/PDZ7X11AS/HMqHcSN+zAfuPqZQmhDns43emPEomjJM4dMzxqs2DIEOQMMuxX0/3RMrZeJQhbL
heUpq7AAiQFpqSbo3ZNk4sCl/4QZB7Ob2hBNjCwRpPSsVQpddBqueArtkIM3Z7jsiix9oehWnPvW
yVDfY67Mwh6WmhonoNYsxRnEsEsrqr4ebgPPWYLdgrEsbxMpIGtrCxVw4JeOoF0wrItdxeiy820N
GvWsYLA+abbERv7UgbNCqIy1XvhfMzK2w2PxnlJd0msy7H0EtCrAtwQgOA9ySGNj1qytkGSggL2B
9UA2kSS3wpjplcw/9y8TULuVxIbounyWHn6d1b1WP+VKAsXRPAH0UCxA3mNYnob4u4nj/3fe5MOO
8xE61sYPse0WHiI/yTlcfyetkyDBg7VRIScXwWPxGAY6Lp/LuCzNAyl8J/DM4hvmrCCM18xPnWwV
t877PAp81qc8iU+2I+rI36pnuG+umvmIC2axzeoCuUUk+mTDfaihy5SmHp71GxvenzFV7vLPXJQz
YgILTFy02bd+WL1aGHodFpcdpo6OAzV0SNFhPrTh0pfzcPp5cj4+Q8HilREvaPtyNSz9KpuhVnh7
CbJXUjA6KV6ewLuVcXhxkwEnJPwPDbE9ExscjxLLdAJg1dD5QNM5imBDw2Ws4K8UgJeWyEqRlvXF
Xki4wLxpC199C7lOhnSZgcPyKAG8M9u1VC9/NApS1UwgPjjbvQwkKwmMpCCunZPxWKKKNW5gpD0e
YVNl/h2KbzVeJpnh/u6tbwrTQXDn5hMPVz98ytHociz6fD/Sqm1VzPIM89ewrIYAehZxsLnAbOUu
xpghcWNG+MPb3X1fnwhKaUKr06YNVlicbnG8MA4eVsJ5jq1J2/ikKDrjlGv3eWOPE3jglmb1vgNv
B0TcrB5iR2XW7tB8fbBFajkbA1wykBRl5BAobgBJRxemI3dCZeoxAevYSpcPGzThTMtSE/Fo+zQo
Ctk7Daf5jyGIbu3qvSW8TxEm3ed1fFQevixp4XktaMsWi92nwl2tOJM4bgwh6juOyhVRjo2ySPDY
RJICDa6grOYzK6p+y2+Jyo3DlIOg537HyGARk/bwF4u/2brRCj2+7UuWQjaRWAA5FidF6m6G1o7i
H1S+0U2xtyHRFSStmpvzO++sM6MEBfeY02H7xc+soqRQttDZ4BJf2FORQNwGGKYMZMsnkxNRWqDs
3F23gnCKrwO6rJa+8Q37aeMDtozd8pwrduSGA2e1YV+5DlYFSBZVH81uituDb9Nq1+Po4FSet/Wg
duInl/tDJw1zllIa44asvogEs8qqXOGGDAMBYECleNworey+M7ZXh6LFOzC2O76pyzAe8uVJGE0r
/TkMnp0OUfvzGHkIAC3ZqxA9mkMbvWyF5DYcCt368Shr2crgDGsFmAgWw0unleZhxEIYP28JCmLz
VFZyAV/QYiVC7b+PN9aPT82UBsymxx8Z6M3kgPT1/JH0SNN/Ky/R2F5Cf9Br6R5MIFFwrD4iH3uo
UI487+qQXuhBFIiJNI+ejVOXnl7NiWtFU+CIYCnDA9kwnTFREEaMh9lw3TBE27HI0TVNrayFCa++
/yvAhEe3C0lCkCGYAhPohe6u2A2uzh1s99ADDF98aBxvOAjIo2elqhTC6VNziwCKMEHsWDYFcuIS
OvQZnRmyDOiTorNA0LyGQiuUPPY6peHEf0tKAFlwHip6831XYoCwkqILDaH85as1PyxcGLxHj49k
4n6r1gCMFlFuHSZrrvXl371IiUsZIpqygRB2vnj+wjOozFZrjqXhPgJZMteP9Pxh9yIJYA9u9LzP
CJ6eHC8JQCCveQKBy1pl1XEcyXhsrFh/wQBMaC0JgMmcyBQ0H0T2j5qF/Q0edlvdB5YGsVloVkzc
ymPhsOlfGDA74l6FanbaStyXuoD1xKu0dtUS0NoYMPDt0GoWMoNjyuy0XFKojzv0exnN+HADjF4C
vuzExOaUzQDQKpqV5OUHTjkeR2je7K5Vc99oXiq6KA6aZisoDyJubi1dQKMl9N18L+Q47aDD4aeX
GcXKH7xLoGbYkQSvyOOK6M8Mh2SfllttLkMxPNPWjilt2V/Pa1wO/MxKlWOePbn3w6SnaXRcg/Xz
UDNsAzytJE2tIE35ZxIFsr6d6rIBcta7MjDVyVzBvWPbFXwLMCMg4ONaMs5iNviecpypy5R3oUSj
VKIX1lYgo2H7vo7zlXEhpChWBs3MG8DLCXPdCStaeWhC33YQ8CGiWsZZUpOP6xzmILMWudCp69sX
WJoKPanbGbojuHUCjp2Ejim/bFLgpCMdxx92mjqIl18DthdAx0sKsh57nR2SzkuPVxE9+Lk79u5z
Rzg2+F9cIIrR3DBXGcdZbvPYerTj6vDV9JgonVXjBSC8HP9CGPDHIbqHmmcxnA90bwyvMOgfZc7V
/vpaeFmXLz9zFCWEfSzJFgzSz/qknRx/Tm9RGUWMAHi+3YYhTSazM8mHBQmEkFN5wGLv1FreyezM
y8k9UNkIgtcUh3jjpM2xLVe9WyaXCHdtZNbcHZoPWpeO126rqx/EzVcV+mI/RC6yEc/h7JGCMo4y
QSbhKfP9b0BVKicc/ai5QQqzG3NiOTSub/3EDZj12hrHfUtT3EX860tz3EtdYgAVEZgARObJIOFU
rqd2kAlZRHJJo0cUqRKcZW2des1KT00wscS0itZsjytJUYGUh40lWT7SkCKsQYZH9hcHVFf5lFtH
Q6aGdf0S8ipnvOwYbq5Mnv11t+5p/eWDGZ7VhPs4WYfcztsePCTyhUkeuXgWH3O7JyWcZKe2m2j3
ZnyzRfWfK1Wh0WzSAEzMowI8qMrGmyfRQ/k7j1qXMA8ubIBh+u/zk3Wi+RFrwyt7XSaNyLeq6Rg/
ucEdRdb0Pfg3YSHXIfaxNFOrYi/V4ksLq89PdVzdJ9n4e69FiHsc2x5G0jIv+NwCLM63ud3M+0qW
xg2C2bxanznjpp4pTOMIuRbXadAyU+vVR9SgWWWAuBHhVDVURd5oAAVCUxF4FrLj1fpMKfoA3H1p
hxWf9/8IWNVoUXF5xCE/S82CK7+nQlbMqKeIaURHZbbnfEElR2G4Uc13YGnw72xcoY5R0VBHok+u
Ki2j2i+iH5oqwiFblEjRxMynQvPR6hqZTR8xQIEVkRTBuTNd+PTGYPMvpECmpFS2fPlbh9GWfpks
CLcaoGNDaeJCmjsHFYd9US4/9sRT9pVqzAGtDZ10NY31Zk+lFbADI29lUULso8hk81XTO7o3W70B
pIuwWhN9x2eQ54lKLDtnYOnNun+W060SI9R8He/n6NKVksI5SRNxgpzx0TNd3ngqErIAo7MrXBpM
h5WUzZWn6am+bmZJizaRbI9KmgFr5dOaxUsyoICiTJo1JW2NxkYUqPo6H6p1u9ZeaUa9Czfn9JGd
Hw11Bz0bXAc8UPWeV83vRZnSTp9E/BdV8duWZTy2Zh1kQSxk2S+NfkjlyIt64OuV9X4doDkWMvn1
M4/9LX5omaR6aWZq8Xbfj+0TQG5/8Dm6S5O6XCrqhwuwM4mUQGSQnPp4a0WOUSQF7a64abwsNRss
Ls2a34JDIIddkAziH9FNI5g8pI8FPtR8mqCYHN2vCnmQq1klLp1+Pmnn4LRzXLSEruEZncIxMkCg
Jgha0egUWwqA9G+mZdE81LjKfqde32Lf2A8dJDbSLj/iGe+vzK9qnbZ5hT7GZ1Nt5Lvohji3kwc7
h54DCBIwbMoiGHc/SegXYjZ2yKh7WGvNxz5jf2c2vSV6kEDGe2YlZ2N/fU5BVklwlWvd/TONPfBy
kPtRupRE6iEvdJwtefd6y0j/aSIaW9p0am3i57zJ5e61lkqPXy/M60U7lMpAFbooKNT90Svv6avQ
Ygg6KcOzpgPH/4ypUujueIyH54DX6OMPoB7KJaS74tbUpiOUALuvxpTbYJPCxE2wTH+AGeZLUPMI
yMyiLpAd5r/4kXxT1KoqeJdIlnlZXSzvv37zKy2Bp3ozwbWyhjQYJBkC376QPfUoS4RQaHJ25/RO
yRXfM91KCIbao5ByOaVarhJKuCIHtvu/4nGcjFcSOA7VYOhMrP5uP8vt4vYjq5Epiu8Q1ImPkJkq
UC4uViLgwNlxFSGUxjqd4erl9srOC9XCMI24nIL76FAnmGiPzqpApY3PXFHzb+9M4RgoOTAInh/k
+H3nJ2eBsQA+8lUNNln+LxjBefXH5nBD/iZ1LNzcaRaxCgfKzC+lUnuHy/5b6o/d6GYDbz5QHzX5
qKAzucsq21w6/Z8+AO8QraIYmeeQl1uv3qHPjKEfEgMyINaubVZJer+reDwdLzJDKhZ9XohilU02
vO7RShTMU88Sej7RMZqVf4cAB0XsQau+3I14O86sXySRzhHPcVC9x6+O7VqLvI7SiaW/Q/KRNiMb
HK9s/FwObeaITW0hvQSLYCd4V8IUiCWHgBmBZZoaluuaSdU7JgVNKcvkgcUE3nYDYy2iuejDb/Ti
s9q3n2a0DRLWA1kcnq5JrlkDjxopS8ZbwEA7bj/QlbsRL7pQaloJEYuxo4qAcSfmzJznpVN6droK
5g4NAUmwVxEbt/5C+rt+HBPhSEjqnalEyIDsFpBfXZOPOcJT3aPBsDOxwwgp+VrZUUxcGcLkchyb
lm7BUD/InsLtbW/SxzPKNrxSs6Z9PoxcZXJhxQlDxtfnu8NkMVSWiN7AufNYxswGXC+Syq2orId/
U9e2k9+p2jli43p124nCEuxEPbMXyf9FlVKotjc93oFt2q+au/wezvO39O/MhptOboVg5a8jxMul
kCYq1Go89F4catIbYSLscAPSygSceiP6w17GnyE6lREBTxO8HboVi1kj5dEv2x567zYIgDre+Hdc
2cNtz4EijmYor01DaQ2vkmuxBaxwdrpLcZ/PGa/mO2sWQyeIo/gVITeTikBf9wRv78OBoV6OxQvD
NC1JHAy67NcyTE86AhhH1hLTf1xU3QicrYIdSJ8Q9OE0WYm3Y9E9eAq4/0DttKhigfUL62A9hmCp
tDP3L0A0PoTqI4mtnzz95BuR5Vx5kNNldENlUSED4AxkZ0IvaAeOAhU/4ZQD25cztcPrBt6S0HCo
pzHWkzCOCQZA/7im5KaKx1h/BMzzA+zlqn+bZ/vwa3OlnBVmHtpG+lAvkLW05BotpsEoDon3UvfH
31alxkFly/hKpITPXyao51JbMuXB9t0QnFaJGptUtjz7ATJYU5i6VGBXBG1ult0LOlTdvk//gzoB
MOC5v1GLKd4XWu9Eav0OIMWpdJXgznbrcWDwfsYv65off6sPf9VFhj6yhQeY5l8b5X5Wgaw1RpML
aPGD27RRaXLqz4tYFbOSjk6cAMOkuj0jgI04sBHoXJ9+0GksojrTrZQeGBavW9WU7aD655W5aSm/
TCkTpB+tEAvtYDKtrBcu6MyyVEFg7cE1Rasd549mk4PImTRjY16lDcWm/Vtx1vtBc1h+U7N1jRp0
RqdethCC0KNhkcnBIG+fgyKQ8GAhzG3/YuDqtDiEAvPedy+zinZeuD550GxPuTMBJZnHLY1XpnwO
1Ux+ooujFM6ZRcqOVwoevRWfcLKZJAyGK/804JOFiFwKRkwez8/2rq8tDffVOoN6VRtseOSEHKyS
R9fBw4dWV8Wlw9BPpha/mSDrtWZXfjgFwwoQVAFeAcjdJ1GbipgwAThUfJyYTgfKUfwfv+BesIKr
i4dPeE255PzP5Pyrc7wKfSaXoSvPygP+tPHCOPV4Ck2vamOY1F8nM/xddC/t5Ej9nwif/ggQee+d
7HT5q3HLFWthyP2Gn2q754c/Dc5y/XP3UHYx6oh1xW4bnwqmA94iMOy7CWQ0wpfsrvgwuD+pGY3a
KPFuUlJeieF+8D6tUaHE/1/nnlTg1rZZhCPjYwHNEz1MMDRgql7lmiN47GLxY+vnnmvrmZ+kEEi+
oD09rS0fTp39o0bwAKC6B0uYUHhSTGFZdydVbNybTnenIOKOJ0/y3S9GoxDJfICLplVWc5UpdHdh
9VIShBS+fIZgo1YVLA8xb5EcVAPw63L3eJ4i4M4vcpNcFdD//P8Nmg1XexfYyHPD3Lg3U3Mf69Ut
Y+mevTnj9QSARClNQn4/XesUUL+Wg5HjmGTJQXlhr6fhfiI8wXgu71yJpJiMcamXrd4A/nc4FR6Z
SnJaMkA6OyQpI7gqMK1ZW0AeVYVOFgi8OKihzVpsJzVQ1fapAr936v0tk9MqzftslIwDmhb5Cd5C
chRXihKJN93JF+IcXEPal239ZtLSQ+ZNjoiewLkKiqN7iZr5p3hF+250Qz6F/bHusrAkZrge5Imt
38fYzD7KGqbqQ+4x8afKNgOUd0uznNABIvOuTmp4QEVr69qJi36jbfL1XhoM9BRXKM0akFogt/c2
E2kdhHN2/03eIJgsqepyCzepd8A0aXoVvllmGV9szIQoThEP8h70elKvjY0ITqupros6JQvbHR4R
B8OnsFR5cMDbMTSVLJfp1QFqKN/yr+X7MAYKxMIzGQ4k0ACgOSxPpM/bR/XWNxDL7lVkUXP9SJSk
2i+5cZNzlbFeMQgSDB7JanVpxMuCnpnwhF86EwjSYoMHTWmSub5CrRySaEG2QJp7rjRiF+ZiUKOh
QFOHmd07fZu6AcECGxzCSB5JDuiDxsR1ol5EOUcspsRr2x0z81Mtu15hPuh4G0lorZE8DcqmpRRt
CqXxnx9M6g4rQRToLQ1dJHGeztYBflbSzIXe//94sEsmnjB+LguquCiy0Ad2AxniLVCmJBcSVcrg
RBNMxwfFLI1Bc3p/dX8mYotI7TP/bup4+JoVu2tSjxy+M6tS3RqTYiBfBMZQQnC9SzB7j0FwXloK
9X9eeTLPpVUn0O8qIe3zP9GjSi+qFcFeus2XdeN4ijUoOl8n94nzIAB14amEXRm/CNQixdp4Fx/Y
u7B5Fhxp7wEug1jtovmSYBkQPjJQio0rdjZt5C+lXETOGuoWyzCVAzsHd3iyLrna5kIDPisiXhBd
06GNUtPG3noAGSgcFf3SfGwSR0xGYuE62Fd+LxerUfW5JWmFUxsszvsruzTI583DzgnigtJp9kDi
Vbnu3Tnmyy8dGN2G8OHKdt2r42zsfB1ZfsQgDh/gGTn1rBDnOW1TKSkDwLffp32EGW/3VpUJgcF0
W9DJo7dkVC/b3jTcXb/xZWQ02GNEyBMh/6uACdICkIwnj8QpC/nOn7HEGW6Y+TBkzy8U+cH3JHC0
3Vypgh++DUUy97GyRLnQDeFEOcFl2dA6u3BaSSqV8mbWKe683OhIM3UcDq4r2J+xw/P4z/2hYigD
ZcSBfZ2NReDEgZKsRmqjrZWph7BpP859YzWpzlFb45nHeYNgXNMOfWYF7xcmEpTmlC72E8KiMf/L
sSm6p0kSp6W7jXnnXXGEzhbo5Z/RAUrbs+b5URG2UI8c+9iA+YfK6caRQV9UZXOdG5qOgkDMigGS
dxzke6ltUGDR2keJYTSY14EmCu6urx1RjRu72waPxhjuYqqWkwvw5QHPlQ49XNsM9AaTCjiBh6rH
BdfYVljkZR1E2w3ThBY7KwtiWwofFzD01NwDnQjhs41y3pPl+B8Ci9z5LsYCq9l2YGmxMW9JYt3k
u+EhORlYyYFaCUAG8WR+A9EgtatGwMKYM5AoBw/pzOzeoI9gBIPkQz7KNvo8Pm4n5+/LpT7bjt9A
pzPWE9iobSY3ACxh0QP2Zp/VwKzQAGZZuf0LE2ByyZXFMOLsqpqiPXbGO+dc6W+IiubyIPMpwbjm
eYASX6LlUcMPFP2A5CzAsU3Fsha8IXurKZC0f+QbN+khfxgO+q3q6qYQ1eH0g1nnMLPupamfQ7gS
aQA9NcPnNFdOZPRVvMhYJl9TMIsCVAMDbYFJjGsXqNPsf5EJ8MG0xDAe7ncuGsmwap3rd6eAHZi9
xuLPkwaRbRyt4CUpxFRmvWXv54Gu2DoRdu2Ax09VTPpOSbukKWAT3gbRvZWXt53iK8VvA6sUcnfY
IL6WK2JXhwNKWsAxCP9Ft9pwVFqLYQ1xvNlKfn15o4lNZSAEW9pUsTSqajAWScWhqu37vAwd3Uzh
ofPtArF0drhUG4d5icCEWFAeUL7lL3TBMXvL/bO7fVTGp8zUR+2eo5sTHbOnRgvvpHo9smyLRjJK
EA1fPfzaKVstThhv+hbQNKb5SYfAiS3sl+zuPVIf1coOoLs6MwKuE/IENRFLRHJyneqW12Tt6RaP
jk9FX+GuX2gjr1TNOPFf4b3KoyhAnYz/YDTlD+Ru9Ihr1sefqNOs5CCVH3VW8ZebTN/TCYVdQ2ge
L0ssRrJbzOUhHtV63c6JFwcrPrup1CLgGIcNQ2oVZVo9YoDqohhZoo4MZ/K58YMhfe9hHPoQPr9E
SM6M+mFQhE4fRgvhh7ufVPmggPoGxtF3TZZWxyrrvjytjD6m6GNHQSnrTynUbytHmTkLx2bq/Yoq
3xjRk0mKY3j8VeB4n64z/kcyhjz7HdIl4f5navPlcnnOoMWRL3DGHODjLxBErVnoasiKv8dkO01V
hfDSpolQnBY9GdGCTpsdhna7DewQqXWRRa1R6FLQciQPKrri9E2TRVaL6g4f0YYCOirHGz23rmo1
MrBa4oyr7GsFgG5XZomPMbinsZel7mT0EI3semCJsTa7JMGk6SbkWZU+pHIx0n6p/mc6maouTFVr
gNOPMSBe225+pNvxy/0yJXdoowrCxtF1AwLiw0rS9PG9WliU6RaybIEv65KV+DgIFsbztxTnLf1h
tR5NaSeYy3p2EEvW4cu9wDiJm+1X2ta1cYlJkwRV9p7mqyHQdHnOrMJUtKqus0/q+kSH2nyzD64w
bLboYRfMcZ3m3JesZU+HlnJug5TRNrBQa8YZ5TjugKC9AEMQFPJkV40Pu0Wc80z/IBzrEwzzU0mI
yWGaqztdcnVslDSiSdzNyMZ9w91jqhXWq1hdz1NYgyuEpnQ15zJLzMnSVfI+Oz17Y63nkj4o3VPT
/NryFqF1hjFi723qRMc2z+uc7fAosy7vC7l3NGXO7Bwymw32+nlkBrLC9ZLwwH9Me5xbzMYvEzP/
/BKorMGmCa6s+Su5o8aOEflm0VGsZGeVM45oWyAX9sHcs1dNVzQ+999ZCHkjhnmzt41u5UNB173C
/+lhUm3wzJSb8yEMosUPF5FvN7ScU6QPZm0XqDxnHQa6qBtbl/h9IE5+O6KN7WNoT43O43T2iCHC
mk6q0vPGEq/ejYLJ1HL5UvvRO379vqMn2NoPjKEA81MuoUwGD5pN/u06H8Y0DsLvusEepJuPdmmL
tyor0Ofz6IUoC1Lrww20WSHhS9KEHC5jCkHmqXQ33quKpjlKaOZuNSI9EX8I70l+XZseCSHifAGm
+WNu7LARp98dRF6kv3ZATPDg6pf2130dcSrkI8uCTed+7Ir6+9wsLCGpUuGYK0Neppak6Vx+eDSI
xevFKCmznSYuQRfwoTw2U8aYD7JOY0QRAs0d1zTk/VSP7uCkpIUPTqhkXwhBQtALV3KKlAvsfzVY
aZ5mku4EpUHpDJDSRxPkhTFq5ZaJqD1cLfvfgo0T1sclICPmWdF7+UcqQhG/ozoVCkMGZOkO78sJ
78M141xKl8q3aZrPtXSuFQBlLpheLI9tYy8r29vACBPcyqF5iUrRxMtTgBTRXV0JMlTeOygO5f/m
j0pYUhitr/oPHwb3z0eqBDYkI4e/VmwERnUbeibWum+s564oaqejFK/wLpyItbDMzvZFP2EihLTz
LIJLzPdne6Nb3e/qTsByi3+Eigf5kvDg9Yup28dq7EMUHg+Wy2zn2RjPuZvR4e6haXbtj998UPse
MPpXukQjgLUjpH69jNndDG54qApZQkV2Xe11gPYcS/WsNWq6jxXa9M5HM730srIU7NHCBvf9C38U
X/2+nMAdkgvU4OKRFWbx7dbkDbe9w0bielZ4KoIiJhFD8tqbGGh+UnwDPIElAaBQrvCsHMxY2hhI
D2vV8E+jCzYXPlJcaAD3jNWvjDxWxVF+xfJNfzuqAvAaGSjaS+vZHWyj6NOEo4S2qK+OIIzrLafe
sq+gprqTWYax+s4eppTlWGYjbhmLXtCTiz2fNj9CCAfJzVM8gx5GAQfu4qYj+1l18fqC4MFD50IH
RHKowUqowMH6al7Ndc4WOhphGwYAMqzrcGO7jDiI8vbgzwVdrhLjXaTqbS0a08IIljkimpOm9d8o
PrAbC3LCUWHFKZ9wFIc3JU9rTPeXv1ohm6lREx7X7zGSD2ef0zyAbV3DxQ700bEmJmPo5ZJ4YMQO
e/3PlBI5lmrBKUsCLf8YDyL9fPngEzgmMTLKasRgtQtEXUP/YJzb8uw51omuquSXeinm7lJxbOvW
bGvrOnTR8syGLd5/bDFJIGMIM8DpM9254SzwJn5VCYedLaO7gZAxOPSft0acqNySQI6knSYtmFrM
EczO/tcISXonRGeSI0hrFSB9Lj02r/MT60G0XmiBqH6wuETDZFB7jHhHbkTtrQ25TjHFYhCi7X2D
GOSuJEgfqN1j3EEVaiCvGjSWJccRdPkZa0I0VRRybpyRWfvvv63ztOW1Fu5nsKWg77sAzx1ZQYob
tnZR93z3Vt4npzsLu2XvGGlMBtoK46wwmTkMHOWLqgB55mUCE12xbWC4NF4eBP0vBtJY6salPxOS
WYreAKev8kdDRId/YZbPt1tLC4YZ9M5pTt+iWI5kcqYCrFRF8Xqwuvvhl3PATRt6V9L9RUA9kXE1
8buwqNqsS0lrPpMa7A6TVlBK+JHt9Ey2ykwwFjGXg460WUFx4l8KHgjAnImyvwvXyhAPntXjribY
JBrZvdsfg6I9fS3bo0vK0wPu1JYMGbV0fyv6391HWOTGO1rJZaY8sDDXyn1uE/yApoWBMsXtJaJA
/7y4NGG8KRmrGFyB/6/lXO1/OXWtK5BgL49kIGtlrZDzSVGlgYHm0oi5E67HVHi9IsKxThJJSFhm
i8dZW24QnuBrKMi746tj/oisEUGDWGJKNTV/Q9Q2PH3T2RPoqKtv/X9KkvIIlwbHuVesaXE7VHxy
VExEl9W2cbarFjx5GRFvdTEu8i5mRv6QM9NA2h7NG6prLwig7CqiXWMaq9eDwLHEGzGp8kmDR0B8
JPkjgrIMIS0O8XOg3YscBlJUBvDajz6rN4IYidWYIgY5Gu5Jt6ss/Y/CzqO1tvi7FSwQI82mRGcf
AifaPirZDAUh4b1Z3fT6J6fNJiOqtA05UoU11I6eY62vl6s6L37nk2oEt3e62yjLZtwiolb+hgW4
Tblmqy4fo/ah9td6mDhJQzHkYQvwzsUbjnh6Tu4f0kEZ8s7xCc5ucmeRWfRWrdqHEU6G19bcHpWm
1aACMreRPvQCELPpBpRJUsOw+/0qOUP1qq5HUa9ttCPMd6FpXjYZAf9hbcQGfGlWXrfa7e2KcjhT
Q0IR0d6cdUT3GSv/7KaxTxyuTebTybfU1BcEeGIUmaE1FF3bSXj6nr3+8BzojXXkb+THJMIz4PbN
DvTD+Y2NDQEAaU2XOI2M/ZPwbOgn8nwffjF9RWh4iAfGoGGVCyAgaT/2Ct1R5XKuYLT6fbAR9XVq
uFN2jFRtPkEQ3x/DKy7HgJJgwmqPQxflckV+N//AavJc2UNr+hsJQQqWC40GvAJOi9HPjJuAXoi4
GCAhiyFdnvcS2T0tcev5/Q1ehlCRcsGcV4itM3ifuC50em9H3X2oeXM=
`protect end_protected

