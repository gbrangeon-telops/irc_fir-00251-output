

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
To/0Y2C4coh8VFh6WzI2wbA/wXer17nunFaUIFXEvO3kBprRAlXyefibFdeqGdMCN/jPnm1lnQge
X/HG5CdHuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nnkNk6e3rHUR8DaNj0C7aWkCs5LBgvWhHhtsF0DtIcgM1egO9JMHLS9VXFoTsIgw40ekMylMZAif
7Mz04TLeS83J8LIkLQIVFCxUoXkTdVbP2vwAOIuzbV0fNimpIIdRDB4Qyrb5oJF0cClV9EVhM+PP
xrslkcRoMPftZWbNXzc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fa9acIf/jWyoTf/ZQQ2RdBUZgeC1x0Ej+f6KiTiJLxfGAO1lB8jxkDwdqife8FqrZb9GuA0CC+35
3eXgFQAQNKjhv24q1nYDvGkg1xQe+JaS1IiyitufBE9Oqujx03ehRV4B4wJ5uK9qxFjJm3WBZQeA
cWZiPDwrU8E27DqZYUHGXiufRSfFhYToep6g7NhnZGCmAfAD7Cg9pLa/AvxaXAS9nnGeBo/RPlyk
G/XXEB6YF86+MUOkeRMAxi86Vcag14njI42hNh7J8Lfa4beMq2Avi5tz5eGJq8y6uRjal6wz33O+
m0Nk9SOLFKAmJ/ib8Fpq77uCjrQp1T7Cl70Ebg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h4sQ6/cKFAjr6toNt8WCtcnxvbT2RbQqvunqru/ZMP069wFljAWXbbabme1u0tsoVT7hQ/OZYU4t
+qXe0sbPKDx8M0x1MxaKDasoQ543qKQAHxR7Bn28bTi4sQCu/+YxH72mTMVFjRAGH6M6e+MhTnGO
FYX19oeiewDQZSakDrY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C8DUdaX7Hd0diH5RVXOZCPD1GItaWr9F/mVcGAwJsPm7j/BsnnF1JwcYxytFDkPy0E+fcaWYKz9u
7/hZwJ449yH3vkp0VWbVjDe3BqRjhnTwAc32kEGR+a+f8HB/6hGM+mJkcuw5DhoveoZqvYIICYqz
iQAjheEs1g2k4DBWxSdaCPNW8fXVd3J/pZQSuvaNRnCtPGOVMt3rO5k/WAzjiaWwDL0KdanM3fU6
uD93ZtkLZCLilGdf0EAax4p+pGVd1C8GYV4+XW66vJmZoT9LNfQ7rG/mL7dKp2aZ5DJPqw3W/O9c
HVwQSloSjbmiN1Fhr9Mdj7iCZycwuy9BYtMK3g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24720)
`protect data_block
R2WwFQS7kiyt0F41c4NRpQvYgNel5H5ko2A6kFsbxjuLzRW+K0YD/wNJf3mXEgdGHCLeU2lKVOXo
HFNmbNQdTtjekQP763e9hzBlIOecOkoUSlq1l6W/g6vfWeg8hgZs4XNBt1NW0Q552aYlcTj4ZnKh
jOFRsvNeYJw5CTlf9b7UipZjvh3Kqvh2rpg/Np8jIQPzCrWAgZG4GZHXEfErgamVxGmk7QCpX8+g
eb/XddOKVGm1fxhZZ5qdTJaG61z6jAe+mwCaSCcE/SbWnLBJeI2wAHX6jRQ2yoZBh2OJYnuQjeTm
Dj+XdE7hZk8EKpAymu02JO8GpLlg5/o7EFt3EJ17ttgR5UMvwcFAKooYUVmhZeEQNzxK6vQW0Z9y
sLvhwc8UyemV6WEUROLnEGntQz3awV8zTI2XeC7lnpN/z7EFPsLr/W5TR4l2y/vMEuyNaAEjt6XM
XtEeMwf0tSgEpUubNr8GQ/vL2f8+4WsXE1HynSkgoB3MuuOc5Hk3n8166SWjYKngbv6YTqjCKOeC
nzzzMhtzPfJzcJQz6Y+MG2VTBvOBaD02e3RIUCGEYqEbDBsKosNwz/Lm/aA9eg/8UgO7dKREluOx
jrvibSiT2V3Kx+Mcq2DHd4WEn8xIMH40Mhns4jGAcYUQ8WL7KQf1NpOSHHjYNPq/4Mdgvbsr8pEa
HxUMTN71nBhSBdWAhb8rgdBMND9ktfJEs7sYcQxdNcYQAs6t5HJLiAPXT7mKA4TpBSKjIHRORHpi
4L+F8wESDRJ29UM4Uun4iFGMWyvCwBzU7gPNdwPuH6ugNNeNPfLrmcs2JRRqM+YkVQUOuXqC+vxc
S34ehUWhe7u+k7bTKKxnTQJsdjykALjgSD9Nyl6BV1XdOz7tPIeXejMNRfIr3GvBTNIXRSte6fIz
Ub+ZgpoSzmZSdqlQrEUuhIOzV+gn/0peRN2qmoPTQ7TY8Aurv0P6Ljxd0kw7LEe6eTqwSg5rRYSh
99Xe2jeaJax+C4LkeyNIDQh2UUKZU6oLzpfL3+t5xCbNEdcqBXfHksoT9LSm4wuCYHfUp6TXwGCZ
q/prpLHU4LgcLisdo5gj3Vn7fL3gBr2XoVER+PWSda1yJ0CzsHtkWWDCoGXxib4ibSm02uMtkzde
HmjaUXKppscbeYG1ml5ysnFg7oKtDTR7VPe/q1XbQOAsOLAL5OoOjXGp/fKA97RhAJ22aB1XWa6q
WUaQi0sTcjFIoy4BQ38g7uZbJy9zHWQx/y0knFFTIQZsludg+9OYyGj9FZVO7g0D32Ei9s+L7pjR
lLjY4swlAo9b2cttXT89e4PJUr6EacxkWHe71nv6SuhAinuXEHVB7mEFWGyIhKv3G/RIC+aVNv6+
3QNLCMvktjCIlyE+wQWuNqt6HWso6ZDCKG6tC0tUI565XXehk6fpbXP+FeDvvU05l/nzVdQQ+IUT
AJrVJxGOtO7fU74hCCU7VyO17HyMZPFUF0AFlUvoAduBXdvg6h6VYnbFE5kfex/XiyHPUf38ulaS
CO/jFdnrsZ1Imoa04h9QLIkqVprH9YqGg3KV65WftFMrlDnchFkfILqZxdgX7kGSSQgkSq5Mb1Sh
PYY6sB8CZSTxSlvLbqQInF3VHzwR4AbrlAeGp10k8DI4m1vSxORbIqbb2Ol3+n1xTbWbT51yEnwR
6XSqqTkDMNDtLOw0ibozOQmUk3GBApLAP3Ar5Tw7taodIP5pLzHTItXVfAcCpcgD3VrgnV7DMJZx
N9TifAWm5quelZWxBGxSH/UJ3CN7apBtXRis0j8hFsmYWv2W4tZ+gZZw2dk4K6apDZw19mj9A8Ec
HNMysRTHayrkkgswrjUqD+3CYpmnBmJki1JDiVaWxPkyw9BoAMIV9Q0XZhiKShocM6VlKZluTT9E
niK+qbggDaAGlTGIqjk9RXBDVIwndKNq9gGAdy4Cxf+9PY4ULex3ksI3vnaC8Rqzq8sTjaJBygD5
H9/acOcrdEeHeqFmJpvYjCwjsILwqWsC01PUonM70rtaBQUt8wq/lW0Qcvi/bLVA3ZTOMMNJBSnt
g1GXzEBBKNc0tu+SEDYo8vkamQCGDK9iZ0hNoItuDNAomDp8CadfsARjmkDCF5sE7Z5WbiEEqymO
6whalDJOlmQxsfOochC06qJn9HwBKe2LEdriIvJHpEe3b4zO13hLbM3wTJSY6TdJvD2dWeQw/6q8
yfmj14FUxqiwnnkPULSMNpsvaIdh8yKlpzADT/gCGGoYe88vLTujSiI9lB+LAi6jO0xC7ZYAXUoT
oMHDcqcxCGo/Cnr8Hvsl0X+jni8uG2YemdTe40J2ylX2HYMRtfA7DOxKwHi8rHztUDQs7x4nEvBJ
SC2/yl3M+yyCbyIldCyltpbjXv4ytoNAm0GPcSSQXYYO3LWN1UraF/kF6f0OtwRLn+tr9nzazpVD
IL+d8Oz+hiMNqcNlQSFZ7gIziQg3PwdA94jtsFdC8hzDGNQp7cjDfb8v2KhO+NoSvrJBqNRjrEvG
93F1PPFRO/Wt+1ih+ji+mdKFCPH9vlMt4qxE9SI5VfBG/40tphyGR8u1k5iYJIUHgbw83hkv+FJJ
NGm7hcprhHj8dg6MyJSkrvSCiyRxAcSv1A5q/vXtuTgc8UTxVVzLnefICIhO0KhfYuUU1aVvA1N2
qGBTHOOJ6A403pNl5M2O8Evs9fvh6jvpF5CTLnqiKnRu6KLpFi4TeluAh9gTw84kwtvGEqTfnccp
QUOwE3g4tKBvHPlFMBKK1WRi3wrHZINSaFdu/M2Q0ipzX2vSMESqQb1XqI8IYw7xsFqf/GaCNkmH
w8bo95lQTIwsYvSnN9tEmdaaienWlsiFrnXYkA6QQuPTpcVNAf+URQKh+AioJqgdh0knR4AY4GLM
1hHQY2uXR9yPnDJ8G1UKvnrcFEYAAOoEcOZ0cEe1rX4R8+35iUmsIfJxMUgK1qHlYY4qfBm9kViL
gaf5rBrltUKaVdc4lsI7fsTlfeWr7iBUmHJEvX97EQScT5dLZlK65jlTsUe593JgS0YhOcoKd9+W
FFiDEyq2TbEG5ILXCcOPRBB6DfurVBqiD7wHz95n0ZcxsfXvrw9GySYflDjXwIp8ao29rl55KC0/
uaEDq7Ez1rNaNN+cdb3WLk2sA5PP+7OBTRBVAS1N9zA729BceljR0whPjWcXzd8QzSz5HrP43hfu
KA3Q91fwF60sBn8qlLXwGSO9DFCKeld2rOBtwqxlKPP80Dy+6WJnrlITz+gk3fhdl2Qz3G8Im/4y
p5ruFj8y4dtpb/h74MUz6COjjPvPiEx9mmomimedEweMLLT5XzQw3XrXJ1249ox9kKx+LMBUMrDa
5U2EByjoGJ45TNFrKzwv9S2op6gSYYqSO5I1wN8yI9yRq2q3D+rtT0dBtjqzGWdExN7Ui06Ahtvv
waJzWKoERi0NyydlIL4omIWi/GUlzIPTAwAx3Ii+nsRr3prY6mlGsFVP4hsJLkk4r1NO6pFeCi//
6Zxq76AoUhdypT8pGSnWaBxMA9Aa51Pgbk0qSceEH39l0t1VtmJhjVv9lvsTt73vOfj91vHPvcAY
pCroZiTfSIx0MtzRZcRKUtrFz5QrmWNCR7/QbGRJMDhV3vxHPjrZ94Z/Ug4gplCNgMsTqcQ7EoFR
O2hadBde6XR63R1vUDX8Xu2cPnfrepF/zytzLh6DvhMpPjcSoKBpK6wt5q58CNWUPexOOznkWpaJ
vxD/VFZWjpkt+b9hyrf7CH/zBrSjtJJGVoTez7/DfxPWbCoSHFTDYZBuguPhEzSTu0eGNue7Tj34
iTbc43qFGOXWT9/ZElSpxK4yaygnL3qXDcKMW0HrlPD0CCl4401G01w2e/IqySZgI9BjrYOTRIfj
7Zxe41gNvf3lBUyX0Sqt3bvjRV1PM6AxQsKNGKKa4ib6T1naXJgLB07Fl8G27aXf0JFQJGDSoVSC
L6R6vvmmBcdfwyNjcOTQIvdNrv7bQU8l/0PuVYOfs7DhcH8g1RL9aKAWE/Ns7X3MVTQnPuyUNSx0
LQ8KxtROk0iYgJLKURvx/d9cwgjTF3eHQrdd0ju8b6Dzw3hQpiViQcXFXpBqK62aizbCHdfDuMGC
4w9th4XvTIqgYFOAKnpgyTzFiOf8xtkX9RoCyhetr6ovh0Kso9B6VvdBIIHbrCgxQ17CcvJWazCu
BgFZJ4qJtainV6Yt5bYOK0N9aNtx4190MgWLce3W9Qe6ApLAw9DBP3Ttmc3sbEU+QidFfIK8Nzf4
OsDjoZZJUGg5Uv1Y+ivX4Q1TI1Ncop10GfNHGz22gEjfXYQKmoSi3Bh6sFs2016Ug5bU0HFvH66k
Subk0ud4ioqHO3sK/f9NJRrEouqqN53lfuQaxEA1j2nHtP6YpDdx9manna65sKdmYg8KPD7LJCh7
rgpZGvvSRx864Tg9KnAu1q0Msnr7waE/EnNxp9Wab0VTQbDdj1jYYS1rSUKc5jJ2U/dmv0ZOFZ2c
QnMbXeXOq8/y0DXdcDuVO5puzoiFKpY23m4L2YWiOqzHQY6+iqOhu6JuNMywH7uNWsDdkIuqLvXm
KbTMSUyavpTPe0WrfNIkDQC87Udk+ShplqwGnvyILPRE00eryDWhSBpFF0f8dncoHTujYoRIJp5E
Nnk3yVh4MB57eIZpB7LLedc/IZRPw4ghntI7SNPV6pJ0/nwplUw54BAW7CpTIlHmtMK9/JIBHVBx
pIJ9noHHKLhfnIYctbtN9pMyUe0+oqPPTmOmDVJ4FDmHsH3JCHz8o38m2wQEbsSkDwwioYnd6kTg
7E9Gab8F1mTZ4LLvRdsFnRL5xBLCONNI97JbuhCKo9CNoHQ/3+tjtmgny+mcZ8092NFudoIrGA1M
qKZUm4L9FG/Ahg2PDnF4niuWjwMADC2m9QCTxsyGy3g5XmVT1rE1Q4B946mN6Rmk2oim7eIsijYr
2axhl+l0ordy2Ue0zEly2HmIV4cRFgmxJp6vDUjAtd+r78aSpL6E1Joyvex1aUcpOaE/GFUPymK5
ZKiSDW8JtWEHt4qQ8/8QaohiJFOfGG6brrQgBP0jkR+HjNvo2ntY/7C/2Gq25DT5CXrxPMMVxByT
D32ZNRDJmW65ouvTYILXANilh1x42MHV5CXRPYiVxl6jJ/uTokzSQRRyVUOOFg/2tmDn1ok4TZ38
NpkvzFgUJhp8UZRu7qlatOi0cCPmwnnBGXV9xG7O8uqghtt/NmewQ3ALFJ4DFyZnOuYgahrx/a3F
KTL80/RmqOtI2AkIVRh6iw7j1rX7qPZeCXeciL8ZjjXuz0NAZaHO7naG9GW3KMjNg5EE4OIHNXDP
gHvLsvmhcmhgDH5pKBmSIQlbK9/fC/sRHJi9ZV5rDw+p/IgiDYhvW+2bCn9R8YrEARMr3vLd9rMj
clAYE2jdCSwpt3XGvF0QBcqxRWRHfh12z9Htdc2bvAj9Ke0/3mkK/iESZkrpCAXUe6Tsm7hmjv2b
uN6foEY++pBN7zZUxcuiplmuBYkj+A5UFEMUvGcdMYgLJ2DfOdjFbAZuI2WD8YRKqRXAdnWzrEl9
d9amJQy+Ix55Yuwj9Gke644/z7slLMcEmeuGLn7evUXKvRUM2Ny55ZM6Fe/LK4WDZ7uQqfQYtTCs
oVm9/01f0XTXDqv6ysHe2pyYgsREbqcDNXWII4Z0oKGQ97R+kQcxaRa8J4JdQw8Al3wxcUQpeulP
606OCoShU/kYVNLU0jkoNvTmgkwf/vJCRf2GQ6h7CMkHiACK8HHN3XVxIdXv7zmaxMLp2UZpJWmn
ohYcP5AKTu9CZE8tAgLct1BnqPu14sSstY6aXpWC76uPMW5cSUQNo1Ayk5zsdjq4c/3e6M8xHdRy
nU/ZeOgetpiQGYqj9qfCiHYtaxUpk1VcsCNT2MqlIggIihuSAjoWmNq5H/m+NnUtnCsAqHPmnuY2
8l+sf4EUUPl6cQynfz5J+pDfRYpjZ/17DaaGNoVoA3mGnqPbKdwWwDhv6PbAdNLypMpd1GSJQ7ik
aYcmD4R0mijcjSPHb9HCNShgeSRE2BxUaW3PevIR5Jm31LzQsvRutngDsVSSKZIS4GtH32/vyd6L
EMJj2S/mQIdPjwzED8Bf4WCbv2ZB0Yk6zJirqGG+G/eC2/5XaVZIifT0uKwdTgM/EwDG6gdbd2mD
jP8Q+z+L9jlZ76WFV/p3jMsqSd7TOc3TEATQ2uKPOIvGDhojA1fpLxZhyx+MNuifTrGL+oOAiS58
OOnULxbLXKm60WyjabQgJLpnvL3/8zNInjRp8Ul2qBS4/ht2ln6vUZTTmNpgMv1xrv1PaxzqAAe5
/9uXRlY7SL6p4YL2lub04fRXPW/7rObCAMxJZQ2WypPo37zIKn2auS/g/rkiw3NR3oY+ZCHFoXr8
6m2trMgmmnM81GTmfw5clFbZEJEm+bqUe8TtKTq8yYa8kZSHsmzZAP+cuZaNgVe8xDHlQMdt/iCk
43WN41Hvrz2B+6+5Dqay9PWKU3mUCami9y5wgujmtoMYqQ5u3q88jV22N26G25Ii29I4n3JcX7jO
z/uupf2oxgDpBhc8aCbaf4amgprmOtnWVuQiyA91egtG9XJHOzTlPBi25ktgm7KIz63Tva/Wigfu
V8QQHBTNATtCyAks3WCV3GjP5sYExWaG7A1TqRUsoRpcw+l3Idii83YXclLeGcFYj7mjXEBBfwmj
C+nxu5jlzaVkQJ399zwjxnmOrK8o9CTsCMeQWiNezuuNNEMt5XZTMNEpwqoTpcQkwXWbEmy8x/jq
3HdXCLZ+Q9NAQTzA2jtJcKik5lDSefpAQn9ZFKjnWKSJe7FXHbPyywHaRU5S+LcSUD38G6noKiQF
m8MSbU5e2fdhrY0dWfY6PZ8K6Hck+uUmxAquJcyIbeGb+on/cYzkpfFhl6eIM13apcVJHCQIAHNo
y79RZNNI6BT3dLRXzvAF9F41JTqnSK8EOeBGyBHdHsMN0pk0PWCAJmCX8UjkiyFLsGpvyQ65jzIe
wim4QLrgIQbvJwyzHTknyOZPwEyAdtSVFfqQPLb/UF862bGZpSPKHCdKztCCtWCCz/0reVFPwhNU
ZbPfGB7pJAl6oERVtHjYRKjgvY1SJAlyzZK1s3wa1/8miCGJs9adG1o6HSn8B2FkV6glZSSHHeYH
0iEegCoYx+jlts0BFyHsM+FZVcTIvCG74UcEOOf0zjGzq0n6rtCAin1OLPpKIhEas+/+6lsHivvS
Rt4sfAzNkCAQjOEsjg/gqffsc782O5tYhpKtyBX2MD8eLgeH8DNEf3OrkX9A77ODmfxUj+8uI+EU
Y66UQYkodHvOaNsviOkLvKMxsrPQqAZA+KfDiw3t+ebdDaL6hcMGB2/hxRKNttHAAIqUUcCmkSh9
aoi0ny/qNMulimh2eKSc+52q6sWKShWZJ6j6QQc3cMQiNP0H9dPVK/c5Em1J/Bv/5/7H3s9U8k1k
ubz5/rrCoaGRuMKlBIl04e/U7XQj+Ub1NxWGf4Z25wdNyBJAPdMvGqq5+nStn6ZyuPT0D3WYP416
rsfDKG7f+URDJ00Q+XJ8hYaRiu1sCmpyPBiKSpXzULhOYO4klq3PAUmSnLIV9pNBw9cD0I5igx8L
1ROyGUtxinX54F3bR8M7HniZ7YDB4G0LykG+nhHIM+wF4wpTo/5DhcXKl0j1opZdWVbugQSpl0Db
X2Y+tWPrauVifClSDnlwfKBQf+4K0IlUTSJc2iTU02NfZgIKG2v5+JFNNDdtjUfNQiJ4h2lGlcFW
dIc/5wwcldgEWthnYATH9hQ8n4HNt98mnCsoSVm9ZgcJvCROsc4xT+Cbyj5NpZLgeG+OjZaMrHET
UntjjA7mCYMQVSdLyJkKMXnWnGav6d126KCaCIAzDsBCJDYla+z1CUWcn5AWq/8/fxYOc6CgW0oo
nd3xuobBytsnGs2XyqKeHxL8LKX++37AR4dMpSLOCFxhaQSDXdXaIoWf265zTkCb5Jx7XCwW4OTm
ImUO+dc7ulHhtqvmSzfr5EaQ4Qf8lRJE54f4O/22c+RjzncIXz14zZtwyTsc3wpaszKiijEEVUSS
Rh4TtB57nVb//CtuwtP42Z1uIWm2D1gBy6azOLLIL/X6i1Hg8UsNS08vDYpQMmF5/d2HnMun0cYT
FctruDqd4jG9Qo1EXTOsOLxGClEbXF9XM9nOe1moreWBQkjzvbakxkIErN/rSh0SqQ5ZCJwaDGA3
qDyFOVPtt2XRMKJQ2okSnPpq3brlO942U8tANBNPICr4uazZm2EekMS+gJ+2YkrPIpYKuVZSH1Nu
ZlEAftIjyFPN9Cd1RkDMzas1VtfLLkXt6XguPuCWyB4vSYiWzG8inrKiMCI8i0ej0BAfmHc7ko+J
wlGqZyW86cq56L6pXj0E4FGDa6cTbT16qb57Z4NQ7v2V7eTdbtAdoRwrrLPwLwd3sJKAAXtXqaNp
rNMLFTI8tjFZcYODPdUruT42b0pCVznvvE+LjBQQwMmshtedZCoG8Lks1z5jL/OAIOhFxuqFhsdG
/Fc561YNhrmQyjdA0EgBQnKW+RIweaAg5AxtMsSJTUPFFHuHBeV8/E31sEA/Kugd+nXgHC6ZWxQF
rGTVFotVRngpmnw+1vaD9Nt37keX8It9g3YoWHEKLAGy0XL9mPCZtEzRsMj92gpUx3yp0sstUgzt
eh1jK/6bmTBj1xGx6/+e4OkRyF+xwT1L1DGFFrcAnut6xGVceC5dscTLLyeAuAan7FIgpl63x1o/
Ac06GVZEbVxGCNpct2FDG4tfRyvX/0n5nxBI28iARfqT20KLMX7LV5NfQAK867a+ZWgUs6Yd9exg
bkyooa5neqIzr4CB6Z6tPZiRss7sf/z1HpSOgytu987XqW1UfXALvqqLOCZFXZkQbLl5v9F1TsK2
EMxGkdaWNVlxepz/q2r5IMIimmZ2ne1zSpV2H8e+S4HhFFnMKdzjpHvluF6j/9cHlizbVBHijKHJ
WxjINsujjuU2YxfIBL/V5BF29G99qyQ3wvqRydZSMJ4zZfetw0zcvPmUvIfoQeVVTxjxO9x7ObpC
aGbfyUf8ZAA3xsFt4GXI6NjvAs1I/RXrKjN2xK4Udq4OzO6u+NQU655bEvPgJJz51iJvaGkpipiS
uOTLKF1GmnVPqcZ92aqRyXyg2g7+yeA2CeMxb+ns3gkpToYXMFM6Ovub7QjiKQ/88cLYwxQZpH+L
jx+Uyz2yIWvmftYXummtzFzwNtDGyx98sETHCntxNlGC7crTnj9j3Y0A0+Q2MSqLULdMXtjmTkRi
vDR7dvOcJJCjx1aP36YsE+E3cOl7b3+xKETLJ/xhu9i8+UXeXEMHWVqFLBYtBRznRzVol1LxKQR3
iVTm9AmnYLazsgpAyEfIyAaZxXopJvzHb8+ojesHwVvMgl7MyiZ5TyRdRfede2pBaqYnKpqxgJCm
oZpQvoDloGi098bTRL+Y++usmaimJTipHhCRQOIb25v0oMQETCx2VH9+wM6y3w5lV8CbaJNDJ1bV
h1uUyRafXqGD8H3DUf5zSVu4Yb+9wPegDM2wiAz1jNeHcOTN36Q/wP23xtk17XeUmYQsc21AqSSy
fE7FzIknxszsYspVcB/ZNbifg1KKm6DOOGob0DIL8mZriV6DccCKoOJq/KbftQSRLirPxAr72KfE
t9YdsCp7gK+e6ZGWIlR/RpinQlunepEZbfnFkMgi382JvEXqW0ZKYRZc8QUFitUNFjWsYBeQ9QZb
BcWkux2osrYTknbpT5Du65xJLNaqMLyzjYonGkaOtv6LOClIiIulTmOnOGHMSvOyHIerHYe3sT0o
HVycFS3E+FLQCxZi0j6W/vjLhOjd901vNGoRlUrEwu5qCj+ARNr1eDJMKt7BPRwpVsN1C+9RWFZM
Erp/9HY6K4XAKvYk1RGtPF3py/1/j+vhmycBVLS/DLMS0bvTmCEcsnEYjNd0Ojc7V0yYsYLZMNCO
cGXwrEOm5WT5ORIUBHVMf1oNzz5CFVU3aZplMqS7pqYi6pY+Uw5KJ7YHj0lWi6kDpCbm4STxwlb4
y1rCuPEtFh2ewIaeAtHE6BIrDy5YvDmsp584rMrnAA5XhjDUCcaz6m5jeEHYivcW5QGKz9/CjCdC
MMZnvvcMOB05juCSTppsH8BvforBElVteY0IgW3S8YX4iN7T0AI5VBo+ZURpm7/9mr5F65WZBKrb
ZB0w5eKs3ZlZ3lXBvVAs+JLItayaIK+6xpmjmtnQFzbDAPEKwSE1bb74zcrw+tf7//vD32HVihA5
Uu5UNazb7HKhQIyPIPAwASOq2zfEOyYoBX9C8TSKJTaQtg3IbR3WxPvkIIHTbbzss3kQL672fDBV
Ohj6qZTMUl+7A9VT7/U20yax47UCMYX2gqVoY8CRkONwNHLSJqzPZ4QfiTjOsNJrjiLTLumiictU
1Y/dwhfzMFUWDjBtXjR0DzXwkJPstOkykLoL14IdgL+bTP9flB58NLfKGvLKOhqxEImKWd7NZsOQ
fKNXuHfZ1eOzewynYrkUVp1sQstwmYOIOKJo8v5f6c7PQt3r3H8O/RFa54TwN1qDxOURijg2YWrJ
9pd+B3YjrF+gLCWNXwdtyrletgUA8oJ6Ye+ddyVSQb7ZHNXHKhSyENodcboDbDwy0L+YWPr1ScMJ
UIqMCLzVRvAoC/X3vQh7uzsYgd5BSAqev95R4zwOTtEBRx6dCSuXgUcahDabdF4AT66nghfHFJ9L
QpJwFntC2hvJXHQzHYuPJD76GI7fWnBxxufbaz7/qF0ywWFpVvtHl7F9/17qgu7gI61w5DFq5Tbw
G8iyDfsgHYpCziyqG9Vh+07tp4EIx3K5Qhu+cpx2Cou3crwck36UuPOmgxr9fLMZXxBVml+LI1ow
WyAKaRgRMNzR9fITTL55qzkYKAJPljSh6Mctz0C7u+2BLeuF3pUOyK2+i23m24Cb8WTcy5WC+n8Y
VOeeWAaGLhZRQKWfjUKSbqhGLotWC/WKPFt8a9n2VOTUcgJeHkL+dsqAfXj4cfn3n/m/2uadGcEa
ksrEWwMQwTFu3STbq/z63LTt2EIv9iVlKyIXbKbjv6O6YfRfD/nVyhcb1TphCDRxsVusbIde8NHh
kHd+YVEwysYd1StIk+Bllz5OWajYfJBQQnChHl3Zkb9NAnJ6F/piBcqfwpSAauJJsXWX/WxS/RQc
QDjUf9H+18MUv+0Cgj0rtCMhXsXzohY7NMtJazIAtjTtvFmALTE4LXskTdJ3RCLIOayfOmmjhEys
AGNIRXD8UHvpubhDJXEhoLpbBZf2toyK/x+/AoJo5Zp+4T6Lt377fghQZnZQ3CUz8cRXG6r/RdBv
HRt3AiFbcqH8CxyNNJoRB/3GSPf0E8gL+gVun/2B4UC0CSMq+Q/WRDWssahpHxTRs/pomvPODJ11
xIDJxmD1krrQXwhgD/qTHkVZLX1FxI8KAvGiTuC59u4JwD0smMY5WjlKC9DAcFYlVAEsI2eQ85hj
l47PfRLA3a+gsOR+TXRjrdEmq2cxR1l3XttUfKGeQ/Ro6qLHKATm/OrSLG0vWyV0OeQUkbmGFT6u
bUbTfvchDDm70kSiL/CfDiJqdZCzqcZodOnQRzfckimpkiQIAGbM7u8o+oiP6RAG5hQG0LL+6qhO
/9I8rud5u8nNfrTQODIyB8o5OXpBQl85tsJCxPQLnkfDgwXNuM2ExERVrQxCj47gIUJuHIEj1nG3
ugsYqpegvHPDpc+LXXBWpAMvcRTto63buwtCn+ulE9bCMTxSEqTnIAKlkiETwS9AbE9zlWfAnV7j
qi9O7dGZKctc/LuNsu55C8yDLFbYKQJmmw1/XoKKQFH9M3wH8cruseX0t7Sp3rdyHvd34xWK/0+u
7gDa3ITBiGmeGl/VXHn8n1KP3X41SjAX4FKsyLTVuTXoJIhN+Z57sR8dhNul7ngJo/yHsy9Pt3mE
ZWdiaQOqr3yKt/+JOV5j6uayzApCvmgQfMIIxGxPuCc6R+bnHpvxqjiGi4O5QcURmdGMUhnmC1R3
7I7vvoRofY1MnMtkVVeIz32ZFMHrLl3bXqneGKSmpBtW+JBgm9OEz8vVmLcelJirVmbZWLdDgDo4
GahRa3uzTGqQ0v/SG2YnWfqTkvTzyZZbD8CUwDJWP1qwbKj6g0WoS4dE+9kMrI5OpH29Tg0XyjI9
eX/81CBdmQy8sf75fMgVpNt3HF6mfyVUpFxcqmm02H5fIO7jd7BBs/pdl0CkbEf3eN7ECERtYySP
X2b7ppJ2TCxJ2+Dls5HzVT09YRPS5h+F0cyfsJFbqBGQ5TxV7joLwwAjQWbc6FCXP4wi94gwhRJ+
UbMKcYcZrc+JoiZLTaVbX+JH1Y6gpKkP1FeAgImbcaCCOaczJud6WRZla8NcBBbm+igOL/hBVVGR
/rdTHs81Sarj8V/snAYrekk7myUjPGn851e5uc5RghHsYmYzMDF7gzQwZwexYPP25lsccB2w7IqO
f3WNXrSz22/vC8rcxiE+01rzF1yc1B6Wl+ezhfQFOEHa9aNZfYzw1f5otQ+DntPYiNgzfXR4XPZb
i32i1I9pF7r+UlWvfGYZitXvbH8crqTHiAeGHEiASCvhfBRFHzvf5aKXArXgYg8WxLPdpZq+FdQG
Axy8YBVRCYKR+HaG7zXcFvMo7LPjt6vecuJPwwg+4Jj0zYIunGvdMc1STl3LeskqGbphL9nJQa3J
wX4aR68IzpXYyadt+lMFh+61pLNhvxkvQjetq2eZ12U7y5UPeWf31yuz5jz5AaFCZRFJV8QzO6co
vAdpUBZQH+1KGAwIajkRAsi/ewLNGrjm+RyDPTymqnrhu8mHGLcleoyuUAbjkLno4dxpb87I9w4N
MTWy+2AKAqduEdp/d5K+6Vfq1GukD35FKaLwV2DaWQVgBTxqTYpVziJaRBxMItDACNa4c6XzZ2fv
Peso+7yAHdqFj3YZUWjK/1TpfbYKYMmAV/hJqr4WCESIK3jGlOAgV3tq6LvZ26oreik6EHgdot5g
ccKQv1c0L7Pp7K5B4jqZjTlEiH5VKAENHgzN0YneNiRqIQMneJ0+hA5yWU64oahHKaSDe4fcu0vN
hvIf7YByj2Ci6YJytmcepR0gC2IoU5fT4yQ/1xQsKOz3t+8wPI+W2bycPvTky24+bfrJwD2mIdl+
bXGxxQ+bVfu5+7hVxn6ww/RNbDYKz9z4oCUbpEiF4BaXUUaFk611Sfq8txMNgqh5Sf2MXCawVsUj
14uXwV6EP/k2BVo7C97mxDo5eOFGmy6B3A/vR4VGPUmb69c0uY5smjKbZNoWZiK9POOS7uftqQfb
Z/Y9S5Jg6CqMHyDdoHxnyvHCwF1tjnDLCBZI1yeRuBHFDy0xQRrwErPrpOz1umBoQFsWmV0ipn1U
V6N0ClikXUA1vC8U+gWVporRoLzBWozNp4Qpa8ffSDByA3zSxtS/rFbPNOhLAW6rFHWOoL/rf93i
DZ8bbT+TEJAm6uRaWAgaiaXwuRHqd/4m1OixiQpXDi/eaN8YbEPBosOWg6hoE+CxYn6C9aO609H4
+eNmaiY/Tmpnt4/YD8Zp6hQdKUyrwWtjAfDArl+UfGvGGIpVhqj51sXHnOMuJVD/sEhj6w9u7RqY
Lfw3slsgaWlA/n3lDXc2WLRNQeRVi85ImSQ+lowuZfuGKtjRqsG+MYzD7RuajTLjmZbb/ksMF8zA
UKwvc7Mei5S8V8bU5U29Y34RMo85djsfroJeeZgL1as4U21NGk+qHfdIP0Ds5oYqPT4mID7WX3rR
vg2vGwdxZw974ZkgIu154LmPXLDo1OHM95ptFF8JyuXfbR4U3TgJ5xPjEYQPVwEkQl/XUh/qodKS
0TrMufLxqhjAbZ1LBXeEI/3F1mnq3XMoCV5i0YUh08MAKF8jDHLla8kq05VZ3ce2p4Hl+IBermiE
KLWX82h8qqJ8V/GqM8kdr8WqQV7Yd3pyAEM8SIPYy++gkR0QbttZdm+XMIj7pdeAE032wiblSVus
NKww/aeNjDGvTMl4fOStkvAJhKpB5XZt/kmp83d2ppwPDNS1AMHX7V/xM1n7Lflclq9XeTtYuhGv
BEYnz3t4Sbf1FftFsOqyFrYNqONp2yCfTQK6MaQPmQvQa+4hjQiauqewVu6G/1rr+WFProBn88Ph
iaJbNAaXLAfk5JV9yFkl4Kz9yOtzifEop8p5UryagT3uiESAAvc05vssMpSAEIbw7G/m/vX4ycLj
Wa4rtAjyTHI8LwFxbQAESQRgYGJGTAMLjER0JPT3/NUKejPoufCOhbY0lebiAbcttSnooCTHjxdw
BiUUIFhUQzVXKHIMJK3a3sYeteMu4VyZGuOOQjBfu23zeVO6hMWwdQIJ03AOYg3tf0nUCQir+njp
LhFGM3HIVZv99Hzc7GXekiE2gnUAyZP1ZlQCxZ5EbiC0EBVZe2bFNvJF5lXxn9t/gSy80NQSkyjt
V3eSQHRkVwtPOdPw0OccE0t9jn6THCm7G4c7PzCAvo4ABSJWO5F3CUZjpF1FdEcYUYWhlHn93cAV
MrqovBmFo4vQbQHaLAbPFlWi6dKcvS9828GFfaS7vOnAvE0+cpXLEcQfPtDxrL4PTzi8MDlFFP94
20QH01CrJ2aClUv7UDME53nlLMzoM5nPIvIVCc+SM0o45tTysDLQ8u+Zc/JEsrgRE/JIAkE+9/u6
nw8ZM7NaX+Pd5By/KH4RwCnezbWcc/gBAUs6/fbrKn4PdxImwFo5J6ME8ykNnRP2obb4Bof4LKjG
nWfUsRBkeTqiltSJDCfko+71DPx0Uhoj6ORyUGHqY9e9cTzVAXojw075O34k0pNF/vyK0nvexs2f
0E13aAflb5dTM8AJeyeWz2QnULtbDUuaLlyU+MSAfS78KD8prOlZa6Uf85txIF1oh1k094Kmpc0z
8Kf9lEggttysa9FX+GjZfyciX0skz+B0ouPuLGYlIpt7ElETTa9NmffJKuROGAlNuMi0pYgDs5AK
5wWS74uY3YbFNHzx8Ev+8ercHKE4CIj26xVx+nzn4qJh9hsd0WBV2XN2NFzwkD1qsd8B6zwk2+CZ
xuzU22R4Gvedcj36UTsDplg9zc6cHTH2YVZTlKEZAoUKpJ6+fs2Y8UO8p8vV+ihYZo/+CXuJadGv
H2Ex6QRaAPtPPB5Hja2YH+1Zo0DiETkRiIaeibuKe30YwW1j7FA/ukiTw7HpPvWdMDCD5D62wY1b
Wg7q6i2XQk+g9cfavX+f3uokuGO4pKgDvZ4lwEzBY74yvayuQSMwX8F/zvFlkKWPPqnpODv1Rl4Z
GMznR4GeAc6AHX69GbN8YKoe2BTT21S8mpP2ojZ7/QcRzPt1JCz0/1sIQbu0ttXqjDRJbhyjIfqB
3Ur305Ws8c5PiHXKNXbVbqryh0WSD4HfCBw8QbsbXbO7G+5/WoZaFbfzfFfKuNF+m9WSaZ6Q4VDW
jK82Iu1BAFl0orIV/hEGOnwK8BLfeXdYITpFPrwe8C3ro59zE321eJnYpOsn7cJnfjxPo+LglSyO
XJgutSirRSS7lSwDQHCUNurpfYM/YmILLqZ8lQO04iepUaRboE8pZVAydHvlq9RHTPP18ki8urcr
uDtR2/+mbBjBRc7bfCUsx0qybbZqbN2s2hK10+eXuLnMyNwFo1VmqVStnvbdz3JuWAtODH3ttXak
qjSoRfF09mUfcwZvmmlHYI9CKM/yGAV4flqFS4ZtCQYXGj4lKuIVbDtG7KIiNPiwFb01fOs+UC49
hbLjBblvj0S3qGs6hty6AG4fhi4kn+LzYQIMT+oNz7nJ0/gcy3DOPc8zrDyhxxmjlIEG1G5sx1po
DSDhRpFEHIM4cV0WswcTSHXdrHrwEFxQ+zdYx4OiDJ5QHgffvG6YAQ5RB3KlfqvpHCmxfmDIQO0P
mYXgeM21JsO7d3FxFSsIrc8isOiwoDh8MU3kK8PGjJlK+YaN1eCuCD077OKCCtVEOv24OtgZ0z8J
XZc2U5A8ATOIZ6rbvA2QWicyLwoLn8HYbr9d1eqvP0D5RrkuvbtHIA9wmYUwOYDd/fzda47zLPNM
I+GGYUklvr4slTr8hvQ+DljRuunXounxbL2qKMXdxgxa5RbjKP3UsznyHMnX5xeTYLfSU+ViSTPM
g8tQTl8xpfaIle/bRmfz9A7Wg2kpLoRehPcRJseQZw5odH7KqrZSuOdkhW/Ww6YLCqtp5eTN4ZaE
nmJzAwE3rfDmubOYdDMwqO5hI+TTXkzz3ZGl24xFo69Uhx69W05lgcZqSy/9otO0i/vAwj1SJsvI
C/LRnQiSt+JYgIwdT1p0+u/tNeZhdSR767XW3gCCFwnF+RczxEgiQi/B0RhQBy2SzMawUojG9cPR
0S17w16hs7fzHWk+mCQwwKWo8BslMbZgjxA0a8oXQAC96ESM6boYyxVOOC4sRkckZnCnRNVt7Qc/
YHo0dPGZXCJXU0JrMGu2hX63vie3ZiScnr2WwjtMaeQe2ilZP0FFV5PxwO/7SyP+gWbEaeiGI1nR
9rX6MWpln7yqnt1Zukw0LmMfuMMWc6quiUAvUEx6ym9U04DbfagDdF/b4JY5Pz4kzw9UZBlr8rnD
9XepNf1Kyfsts6mXo5dUINh46A+WubbH83cWe1CjgCr4qlV0qrWGvq28CjcD6FqPrYCz+pPU3GxG
ST1tm8vojunbKmCeib3o5Jah7/xVSB9wYSndcIHC8ddz8e6nbvHFiKRc/aznwyOODfV9Tis9TV/K
ZY6ptj4b+joxTw4fy9DCVAa8j551ikWTAmG8X1803DqWSvXojTUG2ympx0zDQ7LPGlxVoNrJkYIP
KC0fnq37iKhQStyJb3Qgt0mjb6iPnuT3W/5K6RkL9zkKUnJ1KKPZTomtwwphqwWtBHmENYx2/uqd
chCJ9YPBLmmrjrq5reNbXQewRhLJwd2rKs0b306o7qLMJtRec2+v/J43pC4LiFA1lTYBnnDj7tih
imihxaMKHOX9+RubEu9dAxpvePBN9mGqRK+LBZUGqiDSmE80U2xVR4IL+QnjrfcX3FY7kUKWexJK
9l1HFXCigRK1iWn9DWhnZvAY5ezcdcbZjDxJ0ip3XnhqPEroieeH45I2WMgVi8D+aWK4fpF8AUxV
v2bh1p7R3BWbcEOZ/pGbwg4hVkdhJGK5TNbbRYvt1Dap1iubJkNRTj8iMrqVksDKGpi6emVxP/f9
04zpVyd+bhUEN4dVFHiWdUo21tlCgV0RwgV8rl5FTsS7Sxhiao0D5KJYKoK4HaT3W3YYyVHthHqk
E78HRqg3LPGJ5DMyzSyqcI0SCC2JG6Da2y9vQQ+81Poxq+WaztY75Mvm5KMTiANo0g1KYJLRe1Zr
7Pu3ryYiwF/S67/fIuGy3bVLU/DDTOatcgtP5D4Tf1pa7ZjJX6lYfF0EBrwGfMxolTiRucfRh+TU
jHpcucf12zOddSs0AAHO8G6rUEpOa4c3wsuD5+aWtJiLghf4/9T5red25sKi2BcAMc0+vzf/OrB0
vMu7+fCp1kYeTeaL+8QgXNAzAzJ/zQKdRcKtWGZCMmhn8Dc5aErfXfSlJLA6na+5Be4Z0Ybhpboc
9n0e+347+jNp6QsYGK/EVtxctZOyK7A8j6sHzPypCnSTrIF3i7dAor2U8fajv8voAteoNYWpChCs
AY6IB9p/OccnA3SbwxQoyr3hd0SE8Sa7M4Fnb1iB/6ZiVPjPfeR7MC8ZfgKcpWyx7qPi7AYzjdHj
w8MjjG7+EiJYBy8BcPoiar8Qgqli2ufUppJc5haQM1Agge+Xv2veLH7d4vfY8HORepqjW660sw23
JbdEbmJkXagelEFZ1SXsXkw571a14wwEVs1d4smdQAsY4JVeBH5Y9g4VzJZGcXmILLZSos8k7A/o
wXpOdhq4a+A3RLCCX596GnT5Dsiepyl7vuTLxUnMedt88HNfysIayszsRZxYijp5IsPXOjRwcPaV
lpTyqWms15Vd9MkynFeMgxQrhKLcQoiFCluf4LtJcVcdL40gK2th3UgcelW78J+P5VazB3LJy5IQ
BBcYwkzCYVZMgJjAUFP2dszzGei+JV88P/KkQjCLPrQScwm2cmBS7nWuyMmbZbHvVtq/W2ETx8K7
uBruwGIH0QOZMBAPuyOVm6VqnOaGS71cOC6/SWVQodLZb9P3ML4IBAPtbDiKHxmLKo6IzjPP+FoD
7m6oZ3yV5pZZhlkDNEN1o/QMV6Ek8nR9rmAffoFoiVwsaglThvi+CjEpwOW9RzbnnU/XrA8IPDfW
ChI47jMmWSGHFnmnv2sWxFsiX/WUST/uY0oFx0HYASB8CdNofED+NQvwKTogyfXKOyXod5LVeK0Z
VIn+vzd/c6SW/nEQGmGgXfapidZj+vAmkt4ZK7UuT1Pna6+1tOzHBJDh/DXr4XIUKUYX1y7OiKB8
tIWsiyHT/GvOfnQyv02UtsVBdjwcv3ya3Hj7rno9zcjsP4sQ3D60DGmnqnlnhL+cq3zQy4Vgco6W
6awpmUyfrU75wGVbxoPqLYbdRfxpBJQ9mP8XtmV1TVDlunnLrf7m8CCSa9SXT+mmvBKXWUYtvGW6
JyvVsv4kmWOf3/5VhgXqW4T8gmK/NX3x+1CGSM/C4lhiNtkLiOOySDLnHfugdK8b7ELHLHpQYLtp
Y/8XNTgwRQTFAEzEL6+wSUyVrG2sf6Ew1CwpepEwHAVKvYFcx5h3Tl/xM68PL9vlx7lgK83L3Sbh
qkOJrlwhFfkgVAGuCkty+begcUXlLca+/OHnBwRUivp1KpsJxOC7N4McUuculdsfNd1VF6mlGiV7
4zcZwagrEHc23I6Z+22s8LZWvjXOzTNy0L96JiwfsnytC4OIc3KTCfpzzcNBIXKBLTFpbJXuQmQR
mR9U/tr5GamoQvyVI+337tnunRAGBp9Hx8FXxWpxnJwxEvpk/l3K18HQM0nTPc5I1pXtNbC/eWhs
zmTN+OssuLUTKRjmf2TZPH+dAbqePln6NgximWslu++YTSNKCYhiicnbCYEj9KvkxPxlLoyzIzHC
v596KVcaXNCzewaIfzwu98tSJ3Zhw6S0SE6+cDHTIEMCKV4TlS77hW5I6GfhfdHsSN2kf0oNe9l9
ZGiU3Odm0lzxKai0TdTVMVrC3Iyi+2ti3a5qCX/0A4wzX7862Z2hNUCcXazn6fKbiiqnXW5uUjCK
TKxxtqQWL9CRj0luiJ5n1Mecxs5VhpajAiNeurbfVjFuOZIOHLx+mRnjX3J25hbhW1rUdAJKqYt3
5ytsg+i1ovTxnuRa6XpDQ9k3ZkYp4z03UAjYlgMt1oyUOPe2O1SQZRJVDMOKqTllPAHlSGYDGAVY
yHCUame0UcgNneMJEuyxZQhDxyHc+vSyIuromATDkF+IRpP1VBnDjZL01ayh4xqFTRLnGwJ+rwVg
OXFah5FsH0nWVoAmgn0oTuIyrXlUI1UJOJPsupUEBZHyJTkfBmke/o0L/qh189gzaUQnga9bxCKm
Waht37L0zCAK+KAUwSFE2LdyKyQnblZRdA2tkeiCy69xReJuVPndmpPcDwPjZVPbcSO5MS0LKcsi
HWDHtW7dcaluKRy6U4+ZwuPjHngveaRzi67UlM5M/2JRVtYa2ZTqH9zvrhe4VsAFnEHy+DQdry3E
Jg0n4wHpRAaFVW9CoMQBRxwkB3FRHekuKFoDor0N1ym2kN8dU3zNnmkRXm39thgJA5Y+6vRy0TsG
L3MLT3o1dxYV9X7MlX/+83L5kpg832J1+59Bd68mREI4vXh3To+2JryVegwCoE0noBIKbGegvT5p
QogRpNgp6OM3EuxnNdTUnDaphEVdEswaIDqr3v+mZqnYxxq/dUNN57QKZY+zdCXBSNoz1rZBaJto
UZ6B6z9/Z8QpUhrGzM7dg15fLkiBqq3w2aofOsg4KGrLxd2+/FCKw3UGeaXtWN6LIDZJCyX2+9Ib
fUOxWhLttPxNXqx0c4Ua0Ikh4+3JVechtEUhL1XAtsVSMnJAhgmF1TyPvcwmkNZFrcxIZkR58Day
sZvFnQJmKFxsWxdFTmzr+ecER0+vXoLDXGubS3CY7kxlvSusngV74k0CWs6VmklVDoPO2g80TUzj
MsoeRNntUH4eEZTypn77LUUFukdUjP+C+vd2axAJHCFzo8QvqyuIOFKzO1rkV5HSjBRu60tepB1q
YdRM3X6qzF2i/hoUh9Ed8fljwaKJ63IImT7rm8XGs/FlvSufQQo+f4H2BHaxXPq+ZjvOh+4UB5iS
m6xJJtOk7LXn5hWX5crobjyRrYi7pivXdfV2/1ozxvK/4IAoShBjJE0IsgGdb4Lb1IMOfmDO6iY3
1VKQeOrdho/ZJ7cybbNR4+LUrP6+4NHWVqfO//W8m0/VclQwmIo8mhcniLzRow0R1Uj+6DX05IvK
DJiGWdWjYIpBFsCUmTTITn703DC0FwI8mXo+LlTOeRC70SgbjtZBQPYaG4lQ8SicFuOO7caTLiVW
TB0aHqaeNus4HDtAivWhYPoHqkpz+DidqHB+PZKeAz6d7qSDNSEYlZRfv6Bd5j6HJDitopS/t197
qt2OjQxUHos0HEA0SJJ3IPjXJzZuPCYV0xDcgLdWXRG9LRbuxnpqdg6L0GKeHicVY4LAagxU9tBK
Aa6plC/qxPRYwJQPdxizE0xFYQfcOo17jAS2HuwhiAutKqRXhS2I9TCa/egJ7BN0dyLGQ6+hLjCy
eKX59lMAaaZD57obEcj++G1hAxW0pNZWC5fjbJhl2vj/71TkyxuExmpCDp/0hV8GISNwbaAcYiDG
gwLnpXSCUKJPkqsZENe2cCt8jaXvlOlbZwkGzcySIWsC+7x7wKXOsFLQNytiZ6AgT7qXurbjqNO+
Kl07soru0MhrU15kPx8PQfYwMc0XuxNC4R13Dqt8KSC4wkMlDK1syXMKR9ucAUkyU5lciHeFTYY1
+2iwAhbfomjF84gyooeiSYqIsaQSAw9nJhSK9aADOe4tl8b9r9KgxXd3lfyaea4WupwumYz6l1ko
v8HzP3OyfwWw9JgmxUvkoAaIe0RWmyn9VQvo8Yi27EGaW6NuZfc2NhfU1lq2Cav9XJGbZ/kE9WXN
vKng42tZOAb1RHDuMxQQA5Sz8UEbDmz2uSuzQStDekYvMl6KEKgALEXFjhjcz+suxf5ephelAY++
VfHRtOlHs9CTcF1IPQTrJwz2SW0R2H70K603XoI7Q7cbQSk1EXFqDcHaSQINLAWB2rLrFYfIahU/
6c0j946hsRVk0Rb9Gipy6tKNgyN6t6uSjeJp2JB4wy1dDE+Yw0FUqmoyftP69c8Ao8waTLEfJ4s6
TdzVDDiaA9PaBflZHYZ+cYPwr1zVkCzmuwUigpQ0zwzaPz3yg6xQ3+pku4BqjzMhPjtovrXCrIuw
d7rU/nyQKxfvJMbrA55HHql8iylNAJZLdqVjQszC7cWO31sSkAlJGOIVbwEgjeyrJpmXQU/yWH+1
DKLOHjQRgNpHEbMcT2L87uJVaHMQjs0AuhOwTY1M2dt6aaaamObVf1nPpkNdPHy/b80/Q5mzgZfn
HSrVVc31Q3zui4agkqS2A07ckm6yuHBuf/qn6gOhzoH0K2UOS7/vUZGGKoILRDOPEPo8R+XVzCeN
xjzTLEqYHYfOVKqVMbDV3VAhcmb/K9MtBP4UWhwtYWuWu1Ul9CxegAUR0C+rBzJnbGE8L9JX5P/w
/H9TzdNq9mvQ6cjeLk+2P+1oDVmUZlijYCYcsd7NSJP11djXGFLecow6V2mCKUnXnxuoq8jHI1mC
ZKvqGYrgkGeKKbGjqfOkbg8+bFlu7TT7X5mXRb+/BK+wdhFpRAmuJrQiFcfj2pvivYYYfE10WRYf
+GDF8ckFNgDu4mq4tPQ20K3GidcwbB9ctDhhGhFQD239hKZBhg6k+OacB836rtj45iLmP1BtQ0mf
eZM10YTir7vGRqO0XmynZecX2AZKAOUhNqHSHBJyyphtZBgNr6LM4ZFa53glt1gWluRBO7YcvxTD
Rb8C9YK1xKzilNHJWVKPw3BDyUKjc02Zgo6HclyIt6v6tVli+y3cwmHHszthvnP0ieJKj3SVgxM5
RMerH51K/96c6Axzw9SLUMEk3iKLJkjuQ5JCmT7PYN6XnWRRIfoVOmguorSXdU5jepYf/q0bAJr7
qGoLuXWEyizB8PDZWHjgRBEoW6aFtQssI5Fl4DqqzUPmUO3VUiPBZy9ohDxDm70UGRnTXrZIR5bS
e19rN9/wzvLAO65xMour5GG7IuSicHz5PIvNRmf7jNb9LyOZg+xDUdGPEm17e3uow8OhYn1OoZxn
wio2990FywYQ2SIsO/Z+soFucBjqayjUHtyLcMyDAtTMe/rKDkH//uapM+d2qQmDshd5roS2D83H
OY0qm8zBlYFPTmAwsBM7klT5e17bn3AOCTfqkf/BpKXHUkHSnmitWe/hoWVlQoYsLOmOTG04Kgz6
hyprYd3qO9pZVElszKJ1fUI2DxPiE+czt7xiPfVwVgyGyPlp7F2vvgVVMgq0ZM+597+C0Si4hRoY
T+KNFbOaRsuVqh+1tYDxz5kDsnjD6ketRHkuGpIQrpGm0lq80vkNeJzSCX+1GKBPNcMZNzWOXhOV
2FhUSrEQof/WfQ+JPYjUDlgHtdIAScXfwmKMoZD6v1gvpySGECoI7nxezlFOn8CWg8TzTleRiwHb
rkA/ISTn4ZlOJCqtq7LdenJOABNfrkY1b+EuVo3aQh5UQbKnZwwTkduQXmSZuUakqzFFmbU/uQqT
1INJovLo+DYRQZiNtn6n0wWmbziV7HXFq5oLi+vJxXEQt2WfsnI0N70k52gfbuyFMjm++cHPTu0T
M8rsr4bah4Wu8k9kWjPfOQ4+bs0POvMUF/8iOPtY2IN9G+YyVOU+xEUn5B7skiSLSb9Hl2pssnib
lAHHSRVtH2rK+/57ReKa2LaFYsBNGsmEEybIvFCyjuyQZ4ts03ijiK/elObs6z42a7UpPwiK1R42
jyf1Yi6JE86E6PzQrcdtrtS75q7vG51guJtWspAj0J1vLkirJ5ERjJp+lE+V3SSaWBle6ErWUgFi
Ep57DeinJuP1s5ZkGEnPNqYVsJr9bw0gpb7VVC36L3USd0c3LS4vpxoksY4fhIUWPUIgJsULBHQB
732XTrpCUXkTV5ChTWUMDh8ZVXjp26gsmADdORT3hTSvy6cAutnx1/aopuyxX/P+5lRZ5w/bO+6I
xdGIBriTF7dKqEYbyuV0TOX0H8tWiWGPJyX/n3Lmv0GtWiIlVAi59c/sy1T73wjZ5s1mcqLDdxqo
z9k4e43/1YbTMyGktZYFlzWWqdwZ5jmW/h2CwAx+ohG9PK5bWNVSVNBpNM1n7b9iu33wdON25u8Q
I9WV04G/4vB1nCGTirLW6KphtAibf2VmnI4TtLFaQXagpcmhFlBuakUt26JqVG38IjWjil6if4Mc
IwUT062Eh50XK3CvFbKhmifFvQLZ9MfDH5tyIB6hWRBc2f9IpaG+lExsjUC88prbH5g3NtTKongp
uUIrkpn/t7C6PbOmpaS1TSAUlMLMeuBAvrzfAofD7p4CfeI9V+BDRk7SOo0NAjQVZHRVMi0JlyQP
0nluakPGa3dXOY4MauNuchGQfaxJMqf5gnnFx7+zAnK6uf496APm229BEtUu1y6DfMyKs8MpFN4A
a+H+up8pRakHf2KLhx6Yb+qCccQMGC/keSBw4ao0jYV8F6L2Gyr1hH0g9336ISmusM1W8+iBgcN7
qjKXUDu2bR+K43pexQgC+844m6aScJTqn4EaKOuMt2Q34wB1Qba3gBP7uou5eOUXtQqPQch2WzGv
Z7BEHmsnuokjnLuxkCxTnaQLsxa5u6K1P/eJPRFUqWjt3Cc0ouos4p1qYN8vcQEUs4tYEgh4HRcx
dnmFZH6RdcTJOkWegULYpwDOauaQdptHq/gApgvVkfi1/xLyqQ4kq0LRin62oku9l2VPrrOrhjvQ
/85FCsTrXxZB/xVJnTjdMTntukAOzqd5vZ/w5mastrRoddlBd/gkje6z7aOwsst5hYtPWBS1KHtT
W6HmJvWEPMhJkoZYIk68XMVSTujuWGzvSh8RiI6NJjJgbooiM9T0kjyB9LxO1EJreOIqszM13IMJ
Zcw+sC8xnga10P+QWtYWiTrREHMs3cs0G1izbhjC2A4ilDhsPlhFOx941evIidJCAF91qal43GdQ
aNvSlAejcGb0zcoOh8XDpbLDkpy9SrhRKqzonnpi+XtLOEAn11nAr8E40EJ0xXIWueZwXJP1x7UP
2sRGlqCUR/4pG2Hvot7c3s8rmy/QtzU6Y81XBN/kRLkWyyZ0gsBy6lbRET0awtc4Tezw1JnfXeRw
xkPiwKiqfU7ceJsXKhGtFh8cwfAlvAGvuHX8mws8AVvcuQBwz1PjF2iztsJkmQujnn4i3kgw3vEv
yI+RknbXb37jT7hFckPB4pMCPcQ/G6RT3vY/AVAy75XqM1MxUCrEDUHzdqv/5vPejkXFqakm2IqP
Wy8H+bGo67j9dsHt6hRbn/Vyganq69JFZC6AgrPC1M4E/Pjdy40GoQ2WppRHeBLUmeVlv1YYnwuk
dzwrexUs8tmTHoqHUtjqUHtmqszpmLsB5zV6C69m3vC9p7EUunvG/49cZKj8zzgxSktSBVk6uOZI
WNQnBOApzmEfktP3N2Ckny0STrS+8nQoUfAQlyx2rWYlJq4Y8onE5bYDBF8AycnavEORYX9P3EvO
OcG8ho72IFFBB+UVZdSRJuaQ1dsP3VrRabgP01WPojBlAIfaxGuQNm6KKvw48CFfwibDwgdYt/WW
i7tv8f0uhFbTQBsa4a5O0MM5PPYR+gKE7pX7FMWx4ZyuKr/BwIyfRr60p1lwkb6z2kn6aHHRzSYS
Rmiaio3H30TrAj1RRFL66SVe+OgL2hnk/AfKyN3dEcFT8dAt1qnCGtv4lJ/+ZmEzZRGVccwl5W8S
A8wC6thQ/uN8YyyxZdsOy1cdbkYYvMnQrz0px1zshGCXORh4+3+O0ZUCgGmH8Eqx6rWrGjFCRUw0
hPmZGIoAwkYA0vYWGJBYMZa3f9Zvf8Z1qv6OBlVp5LPTTbngFV8Vn3s9HkEoHpg05BhcvjykIYIG
keMeXg5drveCncBkm39itlz/5UiZo2/GBLyFLE4h0iHLlRUoDbmL37XvOwKmwJxCOG/CVsfR6cQ8
rFjMVH/J9/yrVCFYgEI4TkOyoVik+d/SxyL3HinHm+RYii1xfhTaEPe0f2mdH1PAUDqgKIxvgVKM
F/HNa0roybyAwnV/vgIUUgSf8mTGIWj/tkj9MWjIyIetOpAjXxRJ1ir0hISrl0s417RsWHKWr9PT
UgwI7QMrZU8sOQeLSDZsmZU6hsQ8mvxfDdXTy+MQwKNVEqjaa/RaZCeFdGYmBRB7vae7JyOBWD0x
R1muVmtmDJWwTGUHmhho+/eqvgS2Y+wfj/fdGRM8omsC3nwuZ7UlrOcGj6cxTzuQtSOxDyUnNvZE
maDljrWbE5U0ZnaWiJZ9ks0+8ao6IQuSsmkr4ebRBeFOpd8O+BYRter4E33KrTgzXCpOoIxqty95
gzitnxR6RNwTrWg6THxouPsMcRfVljnTQ01trMzgWjMdZXlZFRLdow1jOKrawnVTCXYBOfVixHeI
0vKOLpqyY4Crb0UJGHlJjxv5VSawRx+biXmtd3hqHQ7sQJgmvFsDFHu4B8wGxPx+hd8+29fc3p0M
3V4oWJLCjDlQ/mHhCm0/ZPLtkvn+H7OnG4dmz86uE+fNQjVGJBqW0IaDGV/QQrfbNz+0OmeWHBAg
2ovaruo2Pheg+lXKdPGyMoyTsCqM+xmEgdDRPLAv4kgzqrfQ9g/H9aJ9sla/v+vqk1yWW6FTBW6g
l+MSGfpP9bDtGM3dVSVtH1qTjDlH2ET/xI/J5NxmHRRXClCXfEMGdeEPoxEq1nF44kjLURCafc6P
fovZB85sfeX2QOGz87J107YBU9wuqFf84FnCNudEReH06Ppc9wDK0oJwXaKNFdSRX97aBrhVND0w
KKyMI6nEsmt6dZE9lpl73v5d48L6yMvaAzVqKcgeSpX9opI9QtELXR55hb9Nbuz+lOr4tvuwXbFr
bxHVIs6w2C0GuDViv0jjOwH8T2H/FKibg0dT8Pz1eqw/rMQB+N41pEgZ/4tCdSUUTh+41EbfxI3r
WjryaOiTG5k228OO52h0DVFvmwnPQImYG2DgQz7TkAZs+Pfp5Ba7ML5Y4n0tVF1oQUN5uQnc5a8e
sstJ45cxp2W+m1t01oEfdmHCY9T8EFGTOfvuriVinr49zbfF5w6lmGoqP2qMM56RvMP3XWmUzkER
aVEzelzMYYLVB8SlWm1NV2cf+wV8af7caNX+Rao54Zekb0W64krRW4at8TlVloiQsGgg/PC2ygi8
JGoFMo8g/l+Mt/H+nXFJZIxqYrddrycvpbsg57Yn+W1Hxma1xx/Apk7n6PfNLq8rvsk65zJeKSk2
ZNmOG3u4CV0BXc+AeEQeyJlVvYjpKi+Kn3TyTBYCNJE1QmunE0p985m84NhQDvFIV0t9jiXw3Z1/
OwTR2zb8UOtXHqeaTmVVh570Qt6HsOD/UGuCM0ALfyuBUHPx1beCXfd0cGEVSw4bnF4+xy5LY3aD
wOk+rQoDxiJNp7sJrZOtAyMi6nDIT93jBChKSI1jsMUWZf47nEVfOlk3anyIIAxe9Si3GmoDMkcp
efes87aSIdqBI8Hp9ETJmfDNWZpWpYcwJrwuZhHd/MDdrfwLM1lEu1YwkauKkXubQd6Y1ovO2BV8
qt69V48CNnCFkGLSHW23wqqcBNVS+9dYke2d7b3+cF2onHw4T+5OUknbI7Es33KyWNVcl/swpm0v
1V8VW1JTQKzqatfcc51FoX/t654FKqL1+14yS1lzwnl8YRayBribICtb3EOHLhFNjr35RVbo9PSJ
MD/InKdozFtJkrtCmfzb42IL3TJS5b8n37cz2QaBNopiGPM9GZqA7S/f953GaTwHoB7wttiuZqOn
4EOy6tqL5xK0kog0q/L4h6+OPad+scdG8Q8Lcm/TH8fS4nPV85tlFsoE0DX3AGQ5zVbSlvrPqFHO
Zv39YrbU5+RcmZ5BiCU8MSXs1NHcPtYnWd/KbzyrpFzzSbfR+9VJZcwy3wEd3WHjDpWFYAeVqVg6
FRP/HP6TeHtUFoB2bAsZ2rWL5/iPqJCVzk/WUYxQm5bZXVWriUu6oWdGle7hR81QQkXMCWHHj+Um
ZyT0sx4Wgthd7NFGG+Sk4xhpTaSNak4hylmU3kfBGZELo1zeYnBJPFC+hOeqeXnICLZHseddgSLy
N9oTN72W3eYflqv8v6SypV0E0+UQ1SesNthCarF9cHJ/hkp0Uh+ZSrSP+bAvSKvmsH74ieMnCoJl
u6LD5fqPi1vyFdafqDo+YGYDPflUBmtu2beiXNrrEa5SCbtZJz62O23LDp0ZSFLS4Na57KVXnmQo
497bUuf3EK5dhE88SS7KemYJcVGO14uF4PxzQq5m/8os8ctZLoH4tQ5679ZABjqcJGTEyWnPs3uO
7WKKW4lutVGFBcmPOMrgsOIAI9gjsSYGcoZ3w18MglfIcqwJVmJGltXmEZyFbo8EJfMPONgq1+mZ
zo2XDGTSd0d09SdWV7szVoiMKVhc9UkYIOFsaSsUNeVv6ShsLuxCxjE82G08dSqVBwCMW81JQoHT
C60T29+En63pRQ/aRtw3RM6goXD+H6dhuM8DHqfO9mGcyhTisU85RrjebUIslZheok6iBeYuj5/n
CcONGdPFRyeD6H22bdLFSDwx/4P4mvbOOSdfi5p+UL+CMrZrQ4w9tu1P7gu5ifdWi3ZiljiLLKwT
Pg/dQNzU3W03FlOUxW7UMY/3wDd7RRo/TTbvnJEBL6BKaMAeQolkSi6klGVfWo80YDUN8CYiGM3p
BGY4v3WtQkFV84pKXcRU9CYSTV5rEBcGHt5Gi9fNS6p/Vx7cmXu0jfE3qsJK4n6oDEq6HN4kS1yZ
R58PldFbhcrAdaK5A605UZ7cEeUGkAtDorCdUIOIJBUCMyXKgXRvYAmnIMKKBAhbPAry70HQ1ZBy
ULpfBNeNT9U1fBHnLUQf+xdTbBDPEbjf2651KVf2wQelkgswlxGXKoQra8BqcPrIR7Z1XhdrMvEW
MavTJ+Qm2hukGN6y5xgf5ukInk38pd3iBt5uq3jXWZA5ysv3T0Q5eEiTzj6zcKPUw0LTC1wxQGHo
LQf/qZ8fsmGF+SkvjUsC/XYIqu1B3VCOk4JsH1wdkZivHEo+EfPBFfDmNZKCcO7XXPQ6AmDoW0fe
1eTW+Qm5g6yVZfnwjfF1ph8sFiJNPyJzJxaYt2xdkgaz+jTxxmK6N6gKLYALDcK07bjr+pCRJb5P
brzTER+BXafTKcw6a2B+Jj7coYEcNSlGSjahev/vV70h0p0QWp/yAYBcpBvkMCdhsPslmc68eUCA
libBsTrWyBCnKmrELGowa7CoKkiNfUT4vcyQ58QMgJxm9rBj9pIrxagD7X7r//t29mokizG4MS6P
zwhRLS/CwUnUNYZ0sLlVaC0wUwN2DtOOXfDLCEg6WQIu2VGI9UFNQNeovSuqpiog44EafiwHoqx2
p7oQZFHvHk5oRqgxIh9kdWXYCURlP3Y35j+DQvZRWD5kqbAesIDdhkDA3Kt2HnGBukcT/7wsIjV2
6WgAmB8ufyMP1dMQN8OEO+qqfOISiSvyPgVWAY6S4iEzDD2wiZjjEEfuPfY9N7mBLwvYp0LG2NB+
KjVYjqgMQdChtKTiGptsIos6cIKSVYqsCvtpbPumDZxYbU4RFP9Jp28tegff325IlL0BjI5JmiBl
6m0bZVBINa+HFyjR84ApaMPQJp3rtVoYQJZy60iZ+44DP5Zs4vTDDHjX0rXJW0x0n5NxRyC3qmV6
02dd5Ljzt7DBH6jmaA476ayq09ZdpNGNIDmAst9C6W/uAXtwDjxNsPosfWYcro+AAwgZZHzCzUuw
UgeFJYj319Hl6/X+Vbu2fmc6A3bNE36u+ORZ8TP/o/cwZSzfYCTAlUoLKPKpRjTJFSMwaUYhDBuS
WBA3eLsllfT+GjP6A1UlLIe85AoN+nNhNetilFxqmVkv3uxz8GeNj1wC9lHI33IN8AaW7AKg686n
Oon+jn+e37N3vmpyQtgXxsBwAQzPHUmxV/Q5RLRHQJw7qakjdECPPJDs9skGLFjYNY3FU/e9T4pg
On+3pzM18TrAbpHGf1oEUZYHcFnO+P9TLIecyhxxjnUBIH5+U0XM3tgTdPiXfHHeMQR7hzDM8PDl
1Nb0Qb+pseDgJ0LiSIGTbkYpyhf0hZfss709r6atPxPbHRRwUNVN6ckt8YhK6whx6uMcdhB6VY/U
v0EIj0DpMO2/wW3mTYRgiv3R23jQ8DolTBuaoY1AwJoUR/3OE6KOWm1X/s0Mcho+EjpGU3rF27Ab
VYRUqxBi9QYQ9HhxxozSTh+sUza6RsJ43Zou1VOyiV1S/iBhTssiCF7Mtmj0D0/PUqn9DhR0rEBa
IMn13xSwZNJdTPEzN9qyqY6rqCr755JNhYZBjU/vH2D+a6w1U5/IQpN7GuswkcG40OSFgGqPB/UO
vIkGE30JkE0B9oQ0fw3VLGaib90EhKUwhyxJbdaMNZksyEsRC5OS6O8OhrXKaZQzjDgHyTfPMZRZ
7znwKjPPQcRKyXEdN61wT5amwe0wmUFwqGTdIshDTqiTt5cBNXCczs8BiuQrTkvL9Kv+GR4DDFNT
D9rHUSvRtsP6S5bGjV9arlEeZHynZwZyjRJxjFfHPdhPj0N3oRpQTMQpOfOQq21MODI2ZezjkoOg
qsfgDGxrRX5RWe4AoMUgVohA8/btSyEls7IyaYaf4ikCQh/NZk2OqaygZS9zDBfr+3lYL8KV7KHn
QkP57m0cM8PU2vN3zzGwcer6FYFwqVv1tjsVpv7zgMm3WgitfV+bsHdiGZ6PLsKZeOnpwjXp2KBa
q54RenZIG1XyB3q0wobbRoAeNVFFv3jde4hO3TpqYVqXJyblE0+opFl9eOCwDklKvhQXi3/EXh6v
uVeu93D26KYvJS4qodcdlLknTpgasAlRNpW8Yxq3SvEq5RPGeikQ878/GEfDaNsbM4nNkdAX8cSo
IGwaempmjAMSpivHFMAdemxZOmZZhwVCYm8YmT0S5M0piUBb9Ka4MNew7oIiKOhj2k0uE2Lyrkq2
KBrcuJ0Q8WlLhfIW2+yI9uqB27xtLYKVz2OnuK7SqaBfa84PteV77xN6L0AlLTSU8jWtKOJe0/MX
M2YnWf5c3rEAk5MdJ6v1CLon2B5oOOf/MbwZ09qhl+x01lU/Otyan/4RRThj6QsLysGYq8BDEDGg
kxQyJ3uEmntaixTFTVo8ItQuVMc4mB903FcS6Vgrwa17WrO4oReTB0WU+VTg8eTe8q8qOEooFj7L
qgYeqKgj4SM6hSPdNSWhauVytS/p974P5rKlMErhNDbMLceAo9YeNg6KhAQJKfnCvJreQBsgPN0Z
jQWcRDlPW7VVNEG7e9oAg3THpVILQ5407phOPSpQFjmroFwD9e/xTj+klrjMPc7Ewh1d6pjdnfKW
ncAq7HgSFRIpw0O7V2AKwrokkPeZX124616sQmNTFdAFEKYJSxwnXUyVUg3omMkjU2MQ8gQARo9B
lK3ZiVDLeuTySoONimgyC1shYWc4gaGUW0LOWB1m4M99VxVzLJJOATqbCW8iYF+15FlZ0O0XekLN
LaH1RpudlZ1Fb2c9+H0hLmd0788jpuDOCf7xNfYyqrHHTKAsvXI/v4IZ34IOKFwiuy2RP3jPMBcE
kt9pGJEnxzIcvgAFLEDzs6iLvR3RXJ7jTOES3bHcZBaPgReTJoodMlIZ3g0+NMzIfJBLO2X9ztQq
k87FmpHFBQykT3IMHIJzVG4lHer8sO4pa81FgzZHc9Y4gnVLFNr0MIwpL7AkzHVz4I8DhK3Dagie
4aAkpZXobaZ0yC8fJoTArS1eftRfCnzPt5PX76HgjBcm3Q29XoOrRVucYOOBudHRbds8Fg18lkHh
jU+hIP1H+04B8qWP9ohyNFYv20TMuRdE/G4XyfJYzkU8aM7/7KhiHORFmuVhSuX1KQNXcS1FpYr/
Y2lD4KYQb50BiEdx5zjeVG/9jXfMrYuCySg+RER7WUiQmWw4yOI4B/9QzftDtv77lz2KCB5EcQDh
pjWEs2wHosFYK+5K/c0icH2tDd6UtdRIHNqWZDz0XAbIwS84IgFt158ypU+UDUwWeXm095ghkUJ6
l1rzys48V4Zthd2Gv90g8Dm8asIOquhAjVbVLR3E+QA6spZGs93wxe6PAP1Ieix/YWursgxZaOCh
VHoNrFFGCSfjSyEqEWGm3w6avDTUsGxerlq8FPoSDZhD+r7AqNdKtYX/9u96lDMoUXCSXnqkPMwj
ScEdEN8tT1ERu9V3qudETUqW/snCAYa30rhMqX1RfS/yxouZ680vwyAGAPH17i8TiDzjj/YPa3r8
rbXIHTzwKy/Yjn0b2L1b6v/tCV7c1aULMLEk7uR8o1HwZJorPjh3G2nzesJMd8Tbd41f7N4TWtzX
ccSK90tMXTxwlrTIHINuFJB4BBtTJR7HBxezzntGDQz1bsIRWeaOxVDrOhZKuRJoWkxE96mxRshz
TkcKdd/K0lPLlQXso1obPwNneN38KWJipdErtAsSkotaPjbQZsYG0LOyD/p7EMo5rO/kveV+qHuU
bI8BiiiYBmdWQN2nWLjD5QFxuI8lupDpbaGabXfPA/o1MirZeV1Yp8bW/erB7c4Oh6izc83HvAf/
2oxV35eZtnRVyiRJQuQZ8sQtWrY9RFHMLvaxYQovpapGaUfUxFTc0h+ThIT2B8/NApcm4/bLGVWA
//xu2DYhWKjkx4RBlUGV7mUzAHW69NwRFgJrgXBCCHarKLTJtO/qHzGF8K9MKEs5Xf5nCrYix6n0
RpjBlTQh7j31tXzg4iwBXK4k1EPPBUAKA2wXxD4GI3YN8aaTEB9Md0TYxb3B+nV8vMJLFMPg+54B
q8yByX9FyNLewiqABC/vTB1sVP/Or0m0tGSg9vzKT7hguyGalqu3MNr+QJ7aCdLwsmJyUSB4iNSv
BZxWyoZYTwtMCQbNGMR52rcKxj2x8okXRA6PNMkF4IWfho/t25zoXYzGG7XpZWNKtDBy+aE2DHsd
FZpM6VWTjVYSMQ0S6fqNh5G42EwOflFyxGM1WZQAaqFrduuvJHVCLX+oI9VYtKQEJPl7gj24JH43
K3IL6M8oPoPdRLYYsqByt+M5+LdOvwt47XdW8LoDhgzcua4tNnjmqtgKqsOWFwFf5/w9c2VDvBAw
HyIwJqNcaEZOs4Vd1vbh5H0Hgi81OBvjjyTJPGVCQ3f2jvZaaWTec8vuJ6UO4ghHgNko4dit2gb5
t9KS7Rb4/FeagmcpGEBQZzCzqiidFh+5liRQ9m/eOGG4rRcZIzU0o+DTbQ9Pj4ORUHJp0R9uuE5L
lzVTC+X5xEyk0Lj5xKjHb4YNp9loXg/lcPHB6qGvdp4ETwfzL0YAB36gj/5x03KampRKx7Frcsa/
ZEH7fvT9G3g0tHrwF2hcYyZjglKfWfFGHJkfJPx294JwbN0sWxetjMZCjxN8atZSAlNrctQI44F6
7jzgqetGPjMbQYW/AjU+5mnLrgIPRyi6AZcaB9LYYAhRSLMQ+NvAQZ9R9wZo2xTQKwCy42Tk5s99
Y9fyK+Jx1cMAU6mjQySkWa7RH99pglhovIL8h7uKCiVV3A6dblFAFRqVv0d7TMg+jey0VovpkJk6
BQkuR+8+F88udhj9PcheQMz7isfI1pSA7I3lVy6YFDVQfB/IcH3lcy/WIYFaLwB/3VEFJ0fVqMHN
Mtmam92fIPMydDLsJA5GfQJPbL4+GV+ajoOESGgJtLGFbGrF8HNYYIKOObEG1dlxCLjotUf/rB7y
l36VpwpC0WBh8OFt6JKb/qekrF4MGzqGwxkBuLfJRERxp82WHG5u
`protect end_protected

