

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n6SxQ4cZpYT/ILbURpz0n7m3/CtPg7Srwf+5G6B92ASMc93ahDGfXsRmbxfQ4itjqNp4bImRWGHp
TxDOCQa4ZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T+03ThTlMB5LbidY7dBVWlYp0mNjkvlbypoxh4ls7n36ZTLkklcCR9ZkGKPsYI13rJYYLwxb8HQ9
lAxKeG9QmQNzwwKufgYFwBDRimvj8pMxUUa5UvV+Um8vyzZZSQmIWtsYrZE6EEbBovwAJw8AOtaR
U6gMXGczY3zuLvGCvAw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xyeO5Evu10M+3X2Afou0ntsX5ZB/pwkUmxi6MkSVEZEp/q8vhRIBXtucD3zi9CwKskciGYDIN3V0
Echz03lkOALKA28V6TwxpTDjOCcWnPUs+SbNU9hrNos5LOcUeyT/Umkuwxvon+y1+GmmTNBs/HsN
LDp012R0drMTXSZtr1fQtCR1xHLj1REwEGmrPANPbJm5g9t7g3uQ7e+eNRUcylifmDkL5SHkZMiP
o5a6WQY9gEml+rOEV7XkaZKFEUQnZO3nxTVqbYgCz7Fr3B2jvSfBBfXQPG0AKW9Iz7aUGng8TS33
LFSc4gt02mCKBH1NOkwuxP/U3rpVs0fnK6xENA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UaJ6dwyNV7zPNxnKVFOwTBNM7GBgDixNLEFTEeGL4zxIus/wUjUkJRcBksOgUQrjesNLi9rSamfz
a+6oBrRU3NMz/a6LqvgLX0FtqLiIT69wj/tO+121sBluFxMRAbLYxwtNx0oswICZG6ot3kY7wUo8
MIP1BRyvBE7h7gUe8AY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iLkN9pn78C1qipOzfdJflxHJTY8JBXpf4rPYSCaQgqf5yt0IOulURCvwg0EGtXIXYL5OVuC8GGss
Cxal0AVlk6DQJUg5tnhgoani3XqnRusVYV7ivY3j4fNdUj8iyFUm29wArxnau/1wGXLQIbXlD+l5
Ze35HAoJRWjnvYyl2fMDrjYG0QtBEQHUh7moVIQ+kI8DwofjU8zFsu1KHGJsBje+80Fr1j2xEByY
nscMu+13hzF1cQaS+Ce+aroaWDuHJWx1kJ8/T+29qUQ8IgrJDtRVEWayMxcA9x6qrZ8JHoIeOcCa
xCl16mCCnpbqxuPBt6lvzV/n1cAzp3w9LmCffw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 87504)
`protect data_block
L+upHbhqbqII2yIqkyvw9bXLj/Z7ZWx1CyHrN26MmAyFa78ufhHA8Sa7X8J2KpQ21WPSwdUQQXIj
UduMdz2bg5RkNeAzNOTTEqnp3+OWcJof09mhxFJq7+mJYsjjl8a2RSRVCbNb7GY2ojYVW9iy6stU
d/zCBuhjaaZ1igA+EP+e2Cl1KxH0A3uuaCjA3r/lJlP14lmGfjF/6F/gshO+r3X/SJW4IqY7c/FN
of9n6CHfdfk3O2pSkAumLfGeGDnDrqwWuBUdFWN/wa4ImaUB735KEhZOttudUkLiPY1cXLgUO2Hd
KtDBvqTwG+gFbMVSBkw8UDduwZu+keRPsPBQedpP6rI5mpvut4uwexTrnnHQi5LYJaWzalljsneH
SRsuXJfPMvvDs5QLVzciUMgjFru1+9X6Tv0nyy9pRXDMdW/u5Qv5OGTGBl9unkbYlQm4YSq9/Zap
81tbOT2N9VZ3XDqVECFp2QNdfvIMhZdR8OGZ3eTKYrjQyJze7S9KrVlE7EFBXLipWcXDWvw+i6tX
r5W318yy85yzambEyfMLXGYD3UHCs59nRN2C6WEyRwnda0wd/TGauVuFjZVaj6940f0QWltlyIb8
Qdt/S/N2fSZDjHKDB0Sib0gkOyQPFHc/hzm5w5gCeoS/azpppPU4ZvlTB560ndPkNf/xhQ0378tX
yNZr9XqYWX2bkfmlzxVHl/ttUAXMfneRGI5pkxpU2e4wkZukSvVaB89do9Un4+aW3PdQ8H2G2cbT
4DKxzCzQUVze6sG7XaJQo8Oigg+Dny7tkx3tlJmli/Gwb+1Cn1qeDLEswBIO9Ceer3j2FH5wcY2o
pysA47GLjyR/RpMdhl3UZsITbpN5H/131+nkOH33oayW4LaHOpqTNVFi3lHrv0C7xF/ze1wrZjsU
OMaNJJQorJBDSRLEK1nGDTPZVnAbX+P3UqbNHEFBqY0qlhYje7yDv5vWekGPaqZ/g1MXkX80ly+C
WoiXeX9VRDRXCrrmzhUaPOoAg3wWo4ZTxsXgok+SZ2/g9On/H/sR14JsN3sY5INQyNFp4jfkZFfn
696A3ajnQCrJeFIbjfF9MESxWfIoAS2cvYFVGYEw2eOKQ/m4Eu8ycuLi70OL080ZoLT1CyjmyBn+
BYxbw54ms96ARdymmJUrKeLU06SmwqPEL+zLffFq02UB2oLtRf6cEist6+CRLJzH+lyoZpbO7n10
LlK7O1k2CzjfBT7MnLr/RNpD2L+1zSwznUu6DsNu1Caj9KlS1392qXTnWyTSozLwjk7qB0rqW+BR
6x4tCIWDuFYuynBMAHCQ5nC4osdZb7R0JBCxBSNdjJnEsMmti8ls0R1vYla8zRfrp9dDkMXeWixH
yz/8XLnnj5g6skTZ3/yT2UVTkjTX/I75znc1yxySP14ka88doWtt18X1yhCl+6Gfii17VtMqfzfM
46vho1j45ZmUQanPBVSHnxTbycwEZeAwR0PBZwFX1O2WiUgKgIk34CtGEl1KtDIcHDFDKwkLmk8F
ooHXLMzk7TpScZ0Jgc0kfWDBUV14lzrv7RtP+90Jd779jdvpmPOePgT8J8st7+LJm0dZeGOC3zkd
R29TyeRCzAVTPDG63V5OiCxi4moYWOWkSHMACq1Jnc14jm58wS4BqLjIhdxDlQ2QnAMoEZCLMGll
4RaRy2S0RTYZUU/vMPyZJcH9qjGHBZ6t5lzR4K5ab0B7DL3+ujkXKpDblWuq2rgHsy2mhC/g+kTn
Bae8BQrBWRGS7pXlJZgxPO3PzKkBePrTKEyOwg2GmRIxVimvDz9q10LJelArF9r08E2H61tACJRO
XooEYUqiWGl31ZVjcdX+t1efzKFH4Qcrx0WFJ9a2hLLLflpLmqb3v/c+7ynSzYNdvQ+frTYGdBzy
bhoj2b0gO9wDVggVzG1Wu3J8r/CttllT/bYyLInxJ4FvO7x/TFzelL0oi7B1mjzwTiE9g1d258Xv
bZjeR5mMGhunm4LFwYscnDkXqvx0hqIo22FbULmuig1CiO/jil9mkShnaPDjS0KhJxb79ZPadO/X
7ELUx3fdTgAAuvVSvsgyHneGZ99vL8CrY+9X9IvRzvidG0toeEWaBNuYC5AOUHFoeBjdS1JgI7Y3
w6r6jGgtHenlMU2xf4fAp8eiUNQlr6GnLSyxcKlXqe+1Zs2HlXBky1VNWY2/PmB5BF8TNpMiQjZP
fummFrCVq323wgiLj5t5Xn0RkgNmMhBUpHPt6mI3MXcuTfDFZ8q9ZCHtfhXkrNmeF0DYlNjaSYSL
WgbW1MkyfZ9wsJmkcpcvZwLRP1xSelT4dsvMS8f0LUoLwT0I1Jjy4eBfIVkoMRBrzhVWHYbowric
fmgy8JDvOkEY/uGyJH5pxpdM+Yy9bBQqBy3VVF7l2Y/CniGQHsHYo6QjUdcG8gtzIRoF8sOAg+JK
tBMq/Ho2BagRINJvG1cpzo/+M7RUeNZtZx9c9b17qxHfmhq0brmwykG78RGxEzIwH0Tu3c1AoEES
nS8X8WgGDcTLCUUZwjv7yFk5NACjqGiaKsk7YXSEaQxHuzyks+TyNEBwORHQWVAqpVtA8F+KmEl2
mnOidx8ZsEafjGgg1U6eGtN1VYMrSOl28zwoj8aYqrdwLcXizfEwO2nb5p267ZRQzDjRu2wUWzbG
x4Qm0pxxjnKS9uv59Dj/cN3H+S/PEYX8tf/eJFJG4R0gywxIySz+w+x09UWdpJzyCRg1n4AIK6uX
wuqnp101/KS/06kqSY5kbmV7q4gOSZSq8uEdjTq5pBPet2N/cOBXi9RItzaf3czEq5WhunenyBP4
Nic+V1wj7KZ/n1FC3KG0X6/p5jv4Njm/LxoGA789coXSZ0O8PJKCHS/mzLaNfH0fXuWto/fCShYJ
BDIzmzZivCaULJsIfAA3+fFSJ7IvLX8novZn1R9mB3iu4htKwC7YY3+jnDPC4HGBvhr0R6EDoHHv
Tor6r439o8/I7aXR3+Mgms/+buOXzqY0qaCMQFm/8NZkeDz6EeflR3VIEmjhVk592GLi8u6h/7ba
lBJnZ7Tfv/om2CrHTrZUPttVfRpEk06yG+OjBxJ8d13xVepxhKn2rgNXuaBGgSctWsw0GDbBcZQ5
d7ZU+vOrJog61xQENy3JAPNq/B0V0YzwRcsdFOQy95cyiBw7fkc6YjNGbRcgWwH/O1ahkxVQwo5z
kiB1eKumh7N5r1khyg7Sq20wj4tp46u7pcIRxt/oYT3gIfZAJQeunZTUmR00JuCbM5VsHrvojurR
kqDHthnJQWlwJNO51PMNbRdbNhvTpCJcSqFXc61ZdBgUrGK/OdEn7raQxqoEbS5eyV8GA0q4WuVs
GqMgorpCjSGza4vFRsvtLBD5A+4c4Hxd8oOr3+Ili996dtohzK0aKIZ/qLmOcLfsImVHonpgcAM/
Bmd4DB/79SNEttFGShZi6ZSeq27F933bq8e3ej/1ADVj700IaGoZUvro55T/3fCCRp3vLW4HMmxb
eGKeMYMfCsXv3TlxnXBZet5PGKZMXAob6FM1HCRMtSm0G0zbotr1gG+SDg+HWFvIGsnYsjW9bO87
SFCK5M5gQs7F02MgHVV2UYa+LJ+OoHfA9hSmA8XhOUEvt0DtvkRTAFwDCTl/QEdKxKo3g7xIonBO
/AHBtkt9UuRLLo6DIMgXmaXLLEqK6uK+AcF/i8uS2aHhQZtTn5sqo96MBP56PsCv85bbz12KrLt+
f+prvQquCCWhNfluoHtA4INUijQMi7YOOto9SVaBXr6QfanFb2oWs8glfVSip+k9XU1+3xgdkQ/2
4CXaw3T6W53fJgDofhRkZTiZqJISJAQFBkIyg2jXC7CNpTxtRhjQp6ZnO2O+VzEGiTmpqYH0V7AC
f/7+XK0+1tCRMB0MGWo76wOXm0DN/VSwvHc+y8aJtcuUNyBfYsPFqOhJHJ+Hhwqa1MXuG9OoXHnK
0zT3+o46g7pWPOhX5vVW/mMi9T6eLOhSx3YOeph/zX4+nPQFeqFfERHeAyVz4oUW/CYUZrb4S9YN
G51R5ctlJtLrms9BivZgl+uqZnXuxfN3VaW/O+LiOBEXbb6BH//Vz6peJlyCJUwAggtWjcjB7uiv
fuGEoVlLu5MSzWpraYWXdmXmNu9Y1lcYuLhPhgPS/YtpyMYy+f0u5tzKwrIQK7/WUqrU0mM2aGPR
SXG4ggzcqERL9XTsseVsVtNGJuQgNAkUi6hP9onvGyWXB8WZ6T1mkacPrAIatgp0za2wO/WT4QOw
8tXqHCrsFA2isgHHlDBxGQ3fvebxTthobUX8tvQPn49sXRvvZX/zIBGzEocqsiygsrkaAKcccNU0
ykc4KOU1hoso7vvMyeWzDUG3r4cQfCgL81wumcfEaY3L24Hn54M8y+DduRZtkC9OhUsA/fDmuNG8
Y0RWxVPKRwlJp6kEQqarH0JvJ9VpjEDBNX0KhEaiyJ3l9oV63bjZrq/fp4DZTJWzkt0NRmGRW116
jLE5nbOCb1sDIUL2YMQgJ9RNUziwQMGUjZZ5zNJeUZYeN/Ptb9SkA1W99oRoSMpINE/X2QZkbi1q
COBwCkBfaXHhcI/ArNKcQLFYOzQ7lx6vsKaJLUPIIdqQrIesRJkVq8SIjrA/SihFZgB/GZAGRolX
erWhBtpVD+RNavHoS0X4B3mzMf7eyFYpkvdcJM3CI+llfnwfLB0J5rDFZr11Vk63CMYMLUMcXdJQ
En1H9n80jWWgotAMyblqjnfmLiN/kbMEYmujm0IJvNecaBHhU+qE5sUorb36/xE3diCkNfr2UdmO
jIHLbwmFk5hOMfS9COG/SiiZSPOivFsdlyaGWjN6V1RLvArtcCZ2CpI6v45xZoiKC94aQ7cFB0s7
HpUNtgyIrJqrAuYYs7F4iIQt4EQZB9cFxscNSgYPxGLqR03GfSyA5JNVBLiMaxAT+RirQo3PDWUf
nsSHIu4lwi7UKalX9vyR7emczD5mIvwI1bXIia4VcrxF7pD0quyg5j2R1jfgwAoJ9JHVIG04rUaX
laNWr3o3m/Dq3LAb43Q3puoLcH1NtKz97W+xKT82Hwo3FXvwx+LB6LmlIa6/pK4bRnpI4B/rGyqL
Oj5R+9o5DGGnL7oluNKCQAWpZXq00fnvDNZDLl3lCXdA5SAOM5YxoNP5TZxvlggXGU7aFXtr4AUk
qKb3MFpP89dFQsMtasN+6Jc5RM5EB7q5W/r0w7z6phQvPRp6X51BiU9zcMsLFvtc92hN1O9Z9wTP
CJDHllQ3tI01diRzXM1juPvuarA3Fqusgiv6s7427scXXwDfsWmtMURmJRRot+CBV6QdTNLyMyz8
A6AttnL4Ef++27JW+4wYTb9ES2FUjpHd515+WY733cUXYCKkF5KMivpqn4MPL7lJR4Q/qm1Znxwn
jBzxjsvyVIALc5QSil0Hy0i48XvjSSgJ+A+EoWpVu4nZER5wX6PT/Nu/ico5Py56OdXDvezPGJ3J
LLN4N9DLUJQTFpWhP8ycp1zyDMDXF8kQ2UYgK0ix5tGfwTWsTLY1O7yEubBZ52HHr+w+r9jE4DdJ
2GnCVVPj80eKORTx3cnn4hgkCmnj931EoF69HOTnOKPDSr30BoSVJxJVEeFN7fJ+0ebKXzxdobAD
cZ6aMvhsK5zHSwvHT24Pdp9upcVZGJ3ug/FCjGnFM/Sjdv6arC1crR4utyryqYVwYUS/gxaA5jHR
xX4GSIwIE/RdJpnRAPX9u26Bpcd+SrMspdq5OcQSae1bYINbZZt6Ng1jUPrNPBB17/3mn6bwaX+T
owNeuG3cbPCEZYNstYhLtDwCLknz87gqLwLkKcTZRjSFzmFUJ9KyW+uszrEmiF9FdqUIGH3DJJOJ
sYARDF7dTmEGQhTe6F0uQAhZ6tn6R3RwgCiirbQkc1Vi6zKuhOJEpiQ8c5K88eJyNUt1qCptyRPV
NyNmJyKpJ0kzYysUXR96JjpBv1X0fe1tpQvF9aWHqE6ntDkrr5sTEqNzZ4rO9cfpfnjaMh5/6Uxg
1FymBPhR4xLskJ3TIpvrr52/vWCl16PIRVk/k8HBb5KCLvkd/s5t9fLrIa6L8K4YX+M3EChgbyuy
WlNeYmEgAdwWOy3IEmY81SB7FreJOlIs5A+kQBvPYRM0ecGds0Fe9MFnW8ripujeUn9T9EN42WNA
3jI/nyn0S+yZ7jfbEm+OXVHIi84PPHY3VvRCVwD0sxZCpROpqCTtEKQmugTORLV3v2DVo9/vl/+3
vXJz7ssn7IoDoP98vDbsApjRJ1hoA38DtDFUrFFUiRvWdeGYTChFwC7d3Uq/Fn3ksEaiMH5imjjN
AxumbA01HGsaVK8FbLoxvhNVU5yiOzMxlyrHnWa/rSmJUiNH+FIdvorSdxVKW/bCVu1iDnagVTOH
nM1331v/kt0uw4zYPPRlkRSmnoYg41MK2ONjSg4Gp4PqWFNnUQ61wpDqGbZDn7mhaRaKeyf+tfKM
+6cijQl6vzGDF560uiEi72gwzRnzdMdZCIEJx052+9a2D3BTapBkbubkGSjHKFdwSCqAAr4W5LvT
Kk50xYKl+PMUFzHJa6yQOt4BN9q/eQy4o3ynYNVUdTU5YjpG2djzPF2nFzcvfLS5q5rkBLbuzutB
FqW5KFI2OYCj1QWYN/UTfz/zADKEpfh0ZERgeOs7CtLIGZ9pJ+PyKnKEcxEb36TDwEAkVflXM/rW
NiaRYxEUrTKp/dQVnsAfJ4/IJp0o63oqgi1q9NdWBozUdMyZRKA/B1FLqJoXFl34CuOZfp2nR8tT
R1j0ouiVN0flhtxgysd/tEPjIkgKzArTBWy8zYEK1UBf6IsYfM6hujV8c1MJ5Fl/KW3w6+O1+xTT
9kZgiTRIBouXwa6JMy8Nwm1UtRyafSz9+ITybhPZXscgBzLZQgbqS22Qbbi++pBC52KHiSpi2ws3
TljtodMZVWSARR1MqLE83BkK4J18azAyESK64qWauSTqvYrpY+Q1zRJXRles4PRsVjKTHQofk/ZB
oPup7/wM2WAk0UgEnvPGRqtfLxmEe2powVzfkmuTyc1hOVH9Ml7h72zXxCI5k8luAotJciZbEyap
x/YHN2Y7vewXOwJTpSCY7+D3vQhydMJPYIjEuuB8cSdq6Oh+6CS+MPpYZUL/NH62qw7+A1WfeQcQ
bLxHYWqj19mCwZG2L4MQ7GIA0Q6vBO8WDclFemg9busmsuBF8yL2RFdvw7/aeS8QU94fxQQmxFM1
Y0njdWyILmRDpZtFWvH1Yz2DvGs6+uobJu6DcVCzlPbRvLBE5bPYTLeTEcGlz9ZpPUHT7JEt3rZo
gHCoSW58GfUz968IGwi9F0I4uHVDTKnMJ4sgVtjnRiuhOzGrmqyIPKYsQqlFScH+Lr4CVmN8wfXR
pmERFJEoShDH1rqIguv9VbkW8hVjo9B7HhpRyuV+LZ6WSQjVB25OZSH6jJ0LQLVuBWUEoO7qmAMv
Tmt7RFVzFcy30nFnscfn4pPhwvpmDmnH/FwhY62Kx9eKYjJL3dPuyn48TVRU/9iQZ0NqwaMBZH2+
CvgOT29tkS/Fhna5AyixuQypprZ6TlQ1Sc10BAtwGlY8YReSjORMeHp182zfrR7asFD0U1yz4HgA
9Fy7ZT7Tv0xAWurgYaTuXJpNlKbCJ+mKPsoW9tP5wuYrq2jA6bHZS9DvPf+XacXp0R+jQTLO/7Ua
XuOB49AIkB7h5fwSKU4N+g5iIJJVXysN4ates1NqbMkY2if0OObSbnAVXsxcgGt65zcGABgKm/K6
nSLtQWRwQOCMT+oUE7kPjuAyNxRSddv08Lyi869CvDl9gTVIJqQzoNI2w57kj1JRWkZ3CrItb3oO
90fCgK6McMXbAhcVLTLNJuy+MHfGO9+VtLlnDrHbqr4LA3c7vsLe5doeBQJfWSAH0iUcYG+lzvuc
YKucvJ/UIvdb9OKoUgMc65IVW2Y2p83JnS00M+3rukuhHboNmd5j6P1dfKOSEhaODM1FVpVySulg
i4Ef06otfzHek3n9Uw9vLqsH+LyHU8X1iSyRCmPlKsZvxrMzlXQ4gRrk1FTtlGRGAX1c3xu4pVHn
YNQLnyB/eAG/fW8fJU7XlMtC8s9iLLkYmJQVp+srvRp4CGDaoptLi1aW1iPh/gIScq5qVs3Sd1iu
1elgoZlIOOnU8eaJ9oFx+sSwhvkRTFfCYCi2YfEx0nYvt4l6GffNhp0f3SFf2DfRWg7T0D0eGUva
IJJ5uu8uN38bdIP4Jpso2djXbT+ArV5HmGOXCy3V+M1htecvHShz8DYOaHt9AZFp7z2o/aKIjUQu
OVhxpLKUSeja3QUkiH23CehaUMThKRFh+qcx4tWjxpItESycON271kvQVE0x4EsFequq0k9P2szB
SxyhdZrF3EEgG8OhtlNQvSl4DFP8G5NBkbAFCVQSp+S8fSGbKHO0ypKwM5oHE0EwlyuWF7WGzySf
Kj96kkHIY9Cix6mSv31ZqRS0xNW3bI6XQ+WCtD8QcB7grlcpmXo8ExDV3L5pBnikMFSMgEo5oKMj
9aURXxXHfZ+/mXnirHotJ8ZIIbhVUcelERK4PUZ6KcD+Xet3e6O8Jdl++RZOib4z1UT4C8s68qte
34gjYsqDKZkGiwRVqa2k5FYaGAkptRs7BukCVmaP4rsIa/+8rW1QStwCRvI05KYkvhp4h2+vzQCM
lUBnkvKzHIJYBsel//Lg5D2oWYE87gDz9F4BGVZBfybXw+pQXXIIDzbPgIG0kRKHEj18stD/X+VZ
1SbP5hsdHQQUJpp1GLHVlkVRWD0Xl+65ukiIlypsHg0W6rKkU4x7dkwmnV016MttCDEvbsLjkHWc
B0PU7frv2zWJEhsiFwwqr/9MwsVgywSPkSJLlk1jmQHEOpQ1rj/w7OZY0HyrepWFM7h37uG0X8oW
bilSURdKHx+jPVK0nXH5ahRxzZlRaZiC3izxOEwEmv+4PVaasLvoAERg/Vv2MZ209HVS4JhgA1+9
VPfIoA1KplPwjC3DhH3Y3rji/X6wW1NUqdnk0zhuBEKJM/BfThjNUiR+Z37nUENxj+azRlK9wAks
v2UvgLB+U0lw0HAVhUlefe686PNkhRr3cWnO8GCsor18hmjOaIyL3SxgA8JOPuW1fk85Q8j0w2XI
rtJzKiViWTpyRSMM088gkCcubH1EJNwqhvSNP6f340lJuaW5KmsDmqbBi3izJdS+pg242p+IWs6Y
umC0Ll8lpzWaT9sKUUZALQI0cuHlElhBBph9kHFLijyteZzUaY+N0auab0MlG/+pgZLxWiwbYAUV
RgA/5eyXMOdgwVyM5xNzO/zah/2Jh7FYfOyxIj3Lx0f/CwWiLIgP+eNFiQqMYWHgzDaKBf6nsIPO
ArpB5gUaUMtsJ3UnW+pYU+VE4B4aLjD7C+HwdIITu5399dLH+dYWFBjDA31yl+M+uGaoeGlVbiqQ
0prvB8TERjxpQra4O2/TOOeNJM8jiqb1qhBsb/OyRhvx81Dl+1uJR/ZX3BiOODbOudn82GpyXWGL
ORzqf+sxIAGKW4XkdrWLmAwahfRptB9s+NozooXer7vmlAFU1pbeyvWSUrWpDAW0XslQoJS1676m
eKRYxn4NRbqHOqEGEhDNdDb9duSXIi30JvDJB2wedPm8d0Xo4Tb2774JEXJxTnEFJWJ5NYexhu7u
ddnsPQ3BatzY7m5e7B5qaG3512B5STLmF/1BBh5QG189YIR2WJS0Ub/UXDLNHM6G9WN6nN5X7u3x
Vwbx91+lQf6d55E2Ly7636waJn78nOUVfSB7rnya5LYMUy35HkbV6ot1JOSbbNLAFIUzzX9DisxF
yZQnY0aWe5Jjc9GiwbVVusDuS3ANktZxsVq/ntnJkJPURTARk+TbI+lr0OgKHsqIFfAB8dIYWwsr
zCRZ3XTMpV9H8jXi9mswX1pf8KbFJUrRZrC1t3TZQ5kEMXJ0YXsf4ZAf1D8r9ABd8Lly59AnMQix
VNlDyCB8VzTmpFZHW89ApiuTDcOedu6tsSookjbFSua14w+SwF5uD/NbIA38qtSn6omDM3oIg1Q2
Jgdk+0rJrXv7kX27snOGxjHShtOd+QYHJ0Qo1jA/bUpWkkZjT+65ARMJNmAiZpC0q3yS1LOwd6Zp
okFpFWgx9KAb/0xyg3NldcfHVkYRvQJoDJJXORMbSVZatU5J5TYoH42WR40fEdyAZOzbgRJ1deEg
zQaT1jAmOlGuyIkoI3H+DKzOPA9ytb2xBpDvDX5ptGY2U6KGVI/9tnNW41J20Znh1NxZz6266ukR
TpK2PQvM1HynsPDLKklRu5aSmQLq1P9K//0Xeob0Y+XPJqDet8TWFVTGTUt21YrfvQdz2rQssrOr
9XDA3Cv23yETB1oTaTI+fKVnjJ4oC1kT8Y+po0+9AQmYoHMSYTyQ3quPt+TWTTTnCd1Z8WKECgb5
8UWkuQn+vQNcem7vtTqElPTqJ59MxgbXikoh7Ea2NEICmWWmrwmCvNOvMg15VSBRvfaUHffUqmAm
Xl6uVof/hLkpxhbJS/SMUAK5DKFl/wQFMteI5HUmnRgAeoSXmuObZBPNku3GeQiErNHSUQCC8uZD
93l62p0d+W9J6cwfC4FYI+sbpD3rrSwW/8OJEFm+i5LbvqLczoPLLNf9eQ3C2JmCtbIbPjUdZL1J
kwz0qTLNLSB/Cs3s3c9SYsY5MJdL7gCida7PAD4xIQF8JxRj5Vejns/O3/iiIw636zYihd0wPjFX
G2XoCTDAKA8Q3++J+YQj6VFpHp+XTQeksX9A18KB45NuEi3AIRZ1P+n06q6KqJIoEzwl7szsDfwu
/CR7wKkmmpfFs1W76xXMehSeXBeitNbqYOeIZSylMCkGA1qy/EU8NzmobVwZ8KZwjyGu46lW69V5
ieMhGx5Ivc2oqY+v7hvktWM2/aMYEAuK3P9lDLB0p3K2VqUuR4WdeOGoF7VyGfXL6kFnRwOCkpwa
eTBCFRM1ZlKQ7AbhhhjrT73EJETVmblbsrje+JctD28C2SPuujxcLaBqDU5aa2hoCZ9n6S33Vasc
JEB04i1svjNikGpCMVrtzyogx/H/C2RDis+oTKiHEHo4jOonMVhSwPmp3hiddmFmv/Mq++DuFM1b
UsZOWkKQRGJH/+Vq6MKVQdcIb3jKwe91QmbWFye4UuAjzg6gcENO9ZYS+ePYv8eg7uvMvMbByIXC
iDvfk+qO2rVTSJuxd7U5UulzIW27PQ05MdvpcBmCWyl47AJyl5aJMd4PkpNEPYXepgsfU2mrZB4T
F9jZ4xZ7j1nzQJFeoXclukTKLAiu76Bi2cFW+sZmXciJX+TjAfxf8LjwMGn485UFTfitBW796t8p
NMh22lL8X9bXZvrg79BZv251KXoZqR6alDsnuWQSKG0XMM6+UuDgIrUu5gfQcAU2Hq/W+jhRMx9T
PSnf7TQZ+d2Bay4TOXDv99U2uPGG+pIKr/gawuUnA2WiWFi5fQl+AgVs0uSLBU/cL6KJGvoW37Ia
4E+cycMRylC/kTpHLozbsbovkUuHfg9TVcWFxvqSBhmByXPoxBj+w2WQhvd/xY+rcZQkWOkKTg10
0H+VB2EZgUmxUpfn3JSFr3cf/lZt1RiMWesYcn1ycTP6fJ6I1lYWWAlW6GwTopMa35NJAURdVEUd
b+euOHIYqquxEOO2JQ+4JGY64OB/f/9XuPjoGz5MVJrASZCRegLx36hB+oPNoFvRtxexejx5sKI5
W5l3BlclwYbtoQCZ38kDj6j9w8un5CWJrykh4I8+4CsFgWO88aqmhszvYwViT2YLRhpbemIVBQc2
zOZ9TlDtx53IGzhB1WIVL83YQI5p7cA1NwlSOkKUL5FKBpvJ0eEiARjSz4DtyhI0eHtjgUvKG6Zv
9ORzu3f52zbLhxD+TjzmpBDmUmMtmxDUhygtUMTJsI6WavaSg70rzmaNG28ahtj1bb38l2UIpAe4
N8ky3WCZE0gessa8Doc3SxtDbixL88mW3F00Q0h1DL/8JkPyaD6ER93K49oDiDNXLXk7OENj2JQ1
7/p7fdN7GlZrRMt4UTGl0QqXqFd1gnSDgojjGx0t6O1EER02fTLlQJry0i2R6aTG+e/extIz6BFa
U8t/Ycj9QlKZnuU9LBpfcI35b+d5NwUJAqdcka4BNdDFlpK23TbOMW6jRWH8rxMV1oyecZMYTpIc
G56tC8adIf2hcfMtxNBMN4AIOQIFijHByLsFt/1s3OQ2wVsn5KZ5W20wx8ijP8F1eWEOt6bjrQpT
7v/X7kP32QniUFaP91g2+LUMgdSelDzyIRTjXqBenk6jbtDb7dQJZm1GZTUFo7jfqbAi/ppvuZ9H
q5aDn2XkMIAb0EqmETk0izBkAlsLKqhAjFQvlwJypyUdFXTUR/Fd5sYRjXL18/KlcnwVa5/fO2sr
ANUPSAsmDiIlGCfEpvf1di6RDfBJUH5vELpT8WylHmPc6lQBR/O7D1dfNw8CE77SZ5FWr89i351Y
kctuVILEGc6cHdOLPtiqSNiApg9VcisV2kXwj2+k+TgOxB48RIP+M+K7/yhEV+LiHDTdqplQvX29
QGlyss4KrKnC2I8VZUpk1tkxw1gDb24xs58jfWHY+QSy+xTWwCA6NFBbdSekH2sXQ7qtdTm8mbHp
s7GBL+Sg0C6kAUyByCHWFyCifZ6+qkXlX1jQTWeTlmNcZqb8wh5kL9G4wnlSq5ISZmHIcMG0roVY
te9T9qKmw3Dmj/LTQvCWia0giEnviu/LqGAFcU+Gp2L3tbsBhq5pgLuUW5O0CwvPvi453Ft5YCMC
bPJFNlYvcCkOozmt5pam2Z+NtayqehKrfu7x/ASGbe73m6ecxzarX7kjkJ309EBVf/p1I4MrRpss
qT5E2N1coyjh/PNFv73X4YBLlA96ycgnv5eCzqdCvfJljGXa9OtWIrfC+rodSYaPMFoToKeooVUq
irDkyLo+i2DjPNz83b4vclxv9OgjlCuIfiity/cwLjYd4VCm9m0a3XEUk8ymovpGYyDBzDFlAIJt
NCpuPcKGs26/6U4HbmYDX2p5dOGJ+BhioT2BjIhzpOYVSZ/y9IM7craRDP8w/+qD2gxDtC2dLaxJ
cyI2F+iF94QqgS8toJCTSeK4YC41zYspWB5WITuVxni2882vV/vpZDf4j/HSdySCXQLSg6yK9IvI
CdQXNflloUNDQxHM50MY6+TGarN0Ls3vxL62c2zMRcCCvnmBkm3qdfFQFmanDvNL8+aXMiTqUpHb
UMdamkjgtI85YR1zOMooV6aC+/sJr2z1GT+LGPH+wgqP7Bps3Yme1CksWGJOOl3yLFlK7AvrXrz8
yMPc5p6+SqUp5pqG6AFxh5IJBt1FbqI0sY3Ju+mG7yliMDqRaqaqo3wotcr8yuffydQoHXQxwjny
Owqy3LtQqcv1DvcjRLpxnC2ENCzDhQJxa11bsca4NzcBtEnPuKIVaPNFPErRpguvm9zKwNzSZ3TA
nYtNz1PpkjQclzCung+nIgEUqVVJShj8g49tjErXw3hV6KUFOPxAUydNjMwOjeGME2egy5Wkgtmg
rverpzitQaJr6m7uObrmIDg7AFomyjcHyawXDucv7j6jjZE0R0hjMw9LUG260Tz/djMqpiWvVH4b
gCEjJyqSoE9FY9T1+7XkYW756JyBSGjR88SuGrbRFkqgw0j0vfftih6lJGC/Y0R2Chq5Ucpiz5j1
H7Huz/sM5zgbxE0SPkhWk12nGrHECdCnSiieaOORR/NJvWqDtCxX87/UCekyMvvJaqnineK4aNXO
XCEgdHcVPuqfwqJXKTTY+6K6j/b9sDWsLzWWMJQvOrGrJeQSs4uO8jPqUQH353WI1zQ1xahyEZv0
yYguxsOyuWW7mRdKtFrJd/LyHFURzeMQKbKDe5XFKUwhLuIMLU4oVDp6+Ni5tgV+C8Ad15NIUAvG
dOVKz4eyNjLFjiEYSh/EE8PoYTH1djl8/HlxNXg5xWgBq/GkZvei9766zK/A7DEFJdoan9+XXiHF
wWlL57f6I+quoTQUgaj5JOfoZl8gecuF6Lj7w4oknJIaSZHYGJSs9/uGi2liKk2V69DzgI4h4NC6
FY24nc/enQSy6q3rHvHe6fOov2nYjXFPN8//Mb0Snbf/2FpMT2aYy/NicKrL1T8pV+Sd7zNAPjpf
orl822+0+clwdVNFEexpx9Az5rPpmi2tyfNJiZfDJ+0qlgaEOjPgoz+rhz7obRivddxVEKy+Ra6L
yLsECtYMcyGtdOuLNj0H9rKTvCjiiuRgopaS42BURL1+smjHJGuwQJAFdIfJ8p3WcaDzHB9DGQEp
tdhWnohFLi/jLOemRk5UQKf95VLOMhaav7XePkuIfCNeG17bm2TQX8TSY6vR8uBDN7jIh13kBy6k
YjEolngOY+oOCmBUXmPHMaCmW8+RWTLX4ktqZhxNGt9SNxFs7ezYcXTvfY4nUoKjRLq7r6JVssT3
5hyK5UdIoHkpCA4T5S9ETY/oJlpkBCfjpr+jKojj/MdOutUkiOEsvlB4znzEYYLgPX+VkBu2ojdu
cbPl7ezLKrgEenKcyN6m0jQjKOB5qi8d01Te44emsKYozGimNX8j+H0foRTLGR0Gpn75f3Qi8RXn
0WnobJ5uRCwtFXJjClAyVcTRij/ejnUzApwok5DV881r4223ou8U4uOwEuC+u1o0Z4waa9HQzHQy
NoCSgzsSanAQcp+QISV333YNuogXJmy7wJhBsZSrb9BT3QKfSQeT82HKcC1gVjyoGAje6oHnZTn9
ZaOE2qa0NzBcmYpzaU+UxFB46Kc3l/xD7vLjYsYCxPn21WPJ+IQ0Eon2aMEWhcPPOZ1ZL2P9WbBi
4hGanNo1pjnj1hR/JVYBAJ4gimtrtMx+aBbo8bBez7Y21tdNSD+rIlSYHKBmuv4Y+s5X3Vr74yqW
2vxX5snnciU/xBKkHhjtCS6ejj2Y31IXRXF+mkP8a4/bFbz1lNlLA1bo62Qud2dZ9wBeM2xL9Mqo
jWcEBNKNc+vPX+ufILCqBCvBwwWazRF66TcSvGXaZu8mPPKdBJvxoxmEmMLxOFlXlQaiWACqHkWO
XesFvGZ1hjkq1wj/uTWOmd4m8pp81obdpmA/82UzxFNiGppvGmYHv+kwPeN36gUy62ntDL2d9Vhs
X4fK6VN9LPIekEDfn5+fBhyMM4EP0/dHxodX9gHjXlmXPaC4m6DXY+u2h7Evto92RWruCrxlzE95
4T7LLxu2Y+pvXfBpzJoq/+NihnCduTRhtO54J9J1KEkvIP0f+GfulzXMw896qSAzF+E0RfhUUgAX
fVW9NOokFfNdWMhb1H+BRk823j0kckev0j62dDfbn1B4BBvtVLQ2JMn8t/vUODXpQ/z+SNpHPgXn
rN7oAQFZWIlzUJHKfYLDyg6sGM79AKU+qLQO9yjdlDeL+VAirylWtx1nApio/wWX+4R6uqFyi17n
J0Zf6et2f6AsAZqiRUYD4QZYPrQ6BbAfe1p6EBxI3y3pa3+sz+v2EorFTPWw4Np4u1vuxaTGvpDv
V61Ft2Dx1srqNXOJuZnFz8+JFKg3xndOCidY9SNR6ImDx8xKkMaG7REShTzXQewZmZZyEV/qCmQb
5eX0L0nci5y9d4cl2vkw2SuPpRmul/iRHuWkIKNDzRCLU31MwwWCQTFoO00TQCawALmLMA0fIsfP
Y17dthswJopvmAS6EwUDC9tMFxxl07jOwXFoLubFLmtX3HkBNmv8gQtXv1e+4JJP+5y5r4FUhS1I
FyYsRigLuJ9SzSYAhPBHskhmYRkZoXuASovwH6425mZA4KwMK8DC6B8TcMX0k6L5zTRUqQgo5CcC
bOwlha+1FS6XAODxUZCumDAdxMB6ibtQUyZLUp/ayI3qPyojDT2ITyKfa4c/gdoze/5NQQSHS/LW
0G4CBtFbwQ8i82rztZwdl1u2dN0WZ/SZKpBDK0hqBa0xu0lCEbjGiqBrBkMBHKDDDCrsQr8TDPfx
cyDWxDH6DaD3HvFvkEOMxpTM7Di2UyiHlPvTN+FzQcjMqBlosmYisCn+qO9qo+IhCThhBPs9YFlQ
32T/dgV0A1ou98vSycU11HgjIOKPQAKwn53YPSQCsjd86b36bvwoVA9qWv4iDKVkinh8VvcLD1Qo
RPE1PAlML2oaRvmm/3JKJvgbSyb5c8UkrBjXWbvGfK5IGopkyO9Td8ML4uJOoEvY0JX26pEv/Hk1
YoJ/7Dt4nwc/dCaiaeu0j2Wk1Bpz7k08owt0dsJiqmigNjijUzYjAS/P0CUJkBZOO48E1tPmM46q
IkTwgHWvZQy6DppRb9w1ZCEX1hHqr/Kd87DdP1luuSQbifz/juKYzGMDag9rAE0kWUXfILk35Cbd
3Z0dewSiiIqI8ogw6SN6/fbl0Y2gP7QxzbHa3tlAIffIwTmfCYJCMKgtkTRV/a/rGF1HD7FX9y9g
wVe6BQOmXtTuw/pkYU7QKH0+6vKJwkY0ltAVSmfEX1qF3U/pmZYiZTxC2M+JOErsAuBGD4MkKEe4
oqpgRBt49d/6jVchPhzMHpcZrY3mlO3L147+wyEKpZOUAOP8xjQH8QwtjIrAq8v2BEV/DntStzlK
yEOdnoh8qfoNW7F5NZPFg0/qvQrLTSB1RrOwCxalPpHeM9dgR1uewCK4pbg67C8v/Ec068rQ3gLl
0e0CSPF9UiB5szkEoiDEY1s8ZHFfWeY6KLgYNtLUQ/OF9niuATZOh7TSBSOAxPmd3PZEP8+rVLPp
pZ0RgZ1Bs71IMClxtg8DwViR4hcp/S6TouJ7VVG4o/JPOEmOddDJW2KE8Qz1TZmpnPaSm2no+1tQ
UIXKTnV0AR5pYsJZeoEUA6yHJ5c0dWyCWt+ar885/QimZlxI/NNCgfHLtFwVXzjsTvdv+QP9eiTY
0NC4MkUcFcCqKAa6ZkBsapJ+DKCz5Qfu4y8TFRoAZb3sTB54MM8BMC9WV0FxnZQCNDA0zyGvwz77
WiFBMHezClix+QkZ/yCZDU/R/QZHWoLfmJvBYx2rNw1Tq7+Ao7DYEL7WdUTTbj+0UdaW8RuX7rjG
Gfb4B4x+cddHO/ay2/HaD0CgOxv17cJdxZTNplqE5a6SqpxFZ+F+zAKK89d4Xr2rgjyrYb3fdrqu
cyC6PJsVwbHc9yxKKT/Y9Gl0oW4znnYLnmKkrJVDc069fqRo6TgvIqxoSGHOKgajApnyhrsM1yQX
/aAZiPSUi8WR6tcuz2VafZA0/TKp0UTHrod3r0AJMowdZyBtOAm4NcH0xC5Sp2drbFUKzOsmvg48
CG+jiiTXXK72r6bZg3yEhXsDSyfapMqHzlRFBQvUQpS4vTZpfOdCFERLEkviqqlnWmg95S+vq/zm
7ZJSpVKHxqDxO9JkTId+QthBRuns/AZims5IGQm1wgCCgzlBmDUcPweE9rgDUfjo7RWLjnT/5A3D
k+tFgQDAhma57BEzzkfYfP6UdyKaakfAOyagcwpPtcI/QsPse7abH+VLYEbHTqQeYVMg4NQWYYtk
voY61wpjwcx4nd9oV7W1XXl7OSHDQOIdj7yP1hLLRWr3y/xw0xIa5fbAQ8tlBvGpihjQMvgicQuv
HJ+o1KswaStBL1g2R1pAnw6HvatZGJ+0WLT547YRr5e48vtmRsiYbA5wR6o1mTNnmO1l25dcyWpE
b11Yf6lKDTyvchNE3h5Y6zpyLp65RsHy2FjER6JKBaIVa1Kn8BSmdhP5fttn4v4E+QoCm6zPKAZr
NLol6gE+YlbcGK0stq+eoiaHvvdLofXRb5x+nNDXfP+150nRc+QI90Xj/itQDhmCvN5axk54x4k6
Ap9Nbid4eeyodRllEffQ0THQZpCz5p5LOpM5OFXhGGnQ8eVFwObCuiA/5LLQrDUjKXAuhCNshnxQ
mWJa5h0QiAi72giZ9gYiC76J9Fs1gOoMZ8BzF5bja3id+2EFyg1gK/KGBB5BbugT9pLVPXMthW+u
EqKl481thjkPgasjY8bExmTDOiYfhXg7G8e9qIDJwDlweXYnpnN64ssIP7amTyH+Pjms7ryAVZ3m
R8LhzSPZi0NlVG9FWklV6vDexHcL+dv3Lr9qVbA9a8QERQNlUsrps5o9G2RdVRDg0fnL1PBU6eNG
rVG+KZ+2m0/nfHO1LHPOvm3FJI1n7jgBUD7/z5YYDLy5mNSUizTGPWLNyAgz6kE7xvsuE/11mVnX
PulvfS0aFAjxUTcXjTqwCZwPWy+9/8zcbdh5OuXjQ1P9+3bsxmUJOK7hllSlSrfmjB6NK+JvYCuS
naD0D0h/h+oCE3IAr0Wjal5u/GcFaCXjoZWHE9W3rJvsWs1/7LbRxC2RRRMW3S9eV860L3uxtHW4
TUyT9Llr32PXAopHCAhhPulS/wMMgP5AIec0QPsodBrkCy2dkD9ugUrp5GPQDQHGVOYcquqoCqF3
1Ei+vDo0hOcUfLvBpCvPtHawRr/lyJQ3JZEUiQFi6u62quG7b6SY7ZfCQZu7EL8CL4Xz5oD2QvBX
VRN+hs5SikdXVty2/qjvlAZy6zQr2XCknsfenbKtSZPzORX6+1gstIheygSV6GGSRHYkLjAsgREg
WPQxL5eO1MLMPPSvrCN5puQBU87Aw3pxqXVD8aPBPIxp88B3tKKw0GMd4uabFWT2l70K8N/izTPx
3Husm3zPk7IQr9Gor0yKUPUCf5xkFVCI6Tq6JhzU5p2kI+Xq18BXOir+IOkxJQzDocuCgIdhUMF5
kioT5rkGg2w88ZBzqEWC9kLVb8eM14CkCbAWem7lqgIvbSTxnfdgZJcl0v7f7dxz/6u6TVrTzjLD
HgrijEqyhs4Lpp5x5hzBRhOho5cz8ZqObayXmgkpzturRXKT28Jm4QWXR57MN2/O/LT52Lbt/E/x
G0j+N1yRwZuHBkZB5LdHGEe0g3adHOnW2G0aSZ7rA4+fzDSZEngoUT/dcBWupTJcG9f4J8f79xKi
TLmHJ+k/iWkAi6U7Ti20+z3DkK63MuklrCAyTdFfquVWzC4YY02o6ifd+yrAkgbtFjvC0lNEg/z7
1vPfkSxHpNx6uVgnVpesDZBzVoTK9P261CXvYyrmIpdmKwpaG0/ULG1uGX5JQ+ZD09woSA06s5jE
q4lh1GKR5JEvjMJc0tPE43FvZOsndM1x8aR5T0Lats1G/nn9ejGp3FUbCvkMx5Crc0Szyw0tidnB
d1JPjvDfTX7t1O6D58weManhTaOPI21mO8apY1yXKNEbYKebzf/6N05nRx2PloixlycG5KFU5aAe
C1/CnJr9YKSUxNXlA/KaDnAOR2tAA3w6Oweg1KrQkaiahAnNQx2E9FIOLf7rVT4nit4amOrPoZtR
CIOkqzHQ3AAZOaLbe4YqRfnpzTiMENHzVyLMIloL6Qvi/ksuYC1K6fZ4OyS2wNaxKZ0FBWUrSB0k
1V6CZ7CS17eSXoNtKVlze/jUF0WhYEFVHbWgJGFJcN7EA7CTaZ0xiR0Mw1fFUbhoret326tDqDqo
5njjghzyavWrARnpJgpEUyRZSxE6vR3jNpp59QbTMPkf6GfRbA1tExLBVI2CPJa4qEtpegvCanXG
GI9Ma47SxrfwJyl6y38cwCZNo9DGurt/zh37JKgz+p3z0MRa/jCkMybsdm5L6Q6TH5zZlc/VIL1V
kbPcnMgjjClpR8OCOsj2gyUItGKQ+TXv9mlMgbXjt7gaACLIZS4rFdcPk1tVINW1JlMm1EO+iV45
anoz0YF+Gvm4ole8T7+cDbMZDW0hVndq5T69wsbzWt6Hgm+LCD+/u5TbzasEfeaWQLZ8G1GjTRbl
taAdLnUonmsEvm3xLcLuIWnj7XPW3wAKHcMB4Qo83lgZM+UDxoaJp8bPqnLyleonc7FKfbiteUOw
Np9LwmC58PvRwRSXwfaURYmA30eZetSAixc+t39i/z26vsX65V6sra7pM4oY5oCiKV+9bvEZMQih
xVPkUbTQ9TcvV5oicUg4o5jbzp1VCFb5YmdnCuutwqsL8rFWU3/WwLpBKtOqMu1qcpY89hklY3Fc
3ohqWnYhQqOCbl7kTChu+D2r5AF3gafKHThhzoSs5hDFygOibK0/gInVKyguXpaXDEEMRvZu2WST
aB3+tO9TMTdMrv6VCOGcxN6y768qk0ArIzGp4TUYgtebB2mTrICf2lnC6KN3ROMdKb0lYyKjURHu
hn1I2q3Lri71wMTF0vyCOrQBqF0gvhZDzvX7iGNGpYA+ZLsrNRuhAsBWqNzbmPAN8YLPottzp2Xl
R8B0N99IkeUBJq+LUdhZQhath8xa74Ft0FBtwLRwDS6DgkGFSzwBCXeLf895xtu3vEFvoVJHnEQz
Bh0c6fLy6r3jkZjoa0xNZC09UzceWbjRyTjgReBEDglJ+NpIlF0+awwquiLiXXlQXO9Z5pE4edSL
PJsE4xamVO66uSE3caHmPWSNSdaDzk2iO6GzqxwufH+k209wfo7ccXxInJti82fNLT8Ytj2Diy2m
CZy5rqAiGK4JFfEObERxolqx1X6MRA7zsc2+Nleup93p4lSmsrPGqohslhD18d3qqJrLcI6R6Vw5
0iBifgFCWVoVpTklt7USRC0bW5ouzM5xWcLe3FRWXM31Oqcjo/oiPWnMdKxQorE8q+TefZrY1VJd
Le128vY5Zhi6xR2iw2Ms4S8oOifzlu2KMejLkwIYVbf+OMa7KdkfEZpA8BofKJB/yE/w/IyBfKeA
ZVAOx//XgsbjoDDKb6XMahJVOj4wSAbs0BZ52hvejqekbfssI4b7juA8iKGimUiMlTxSGXZfih/k
rjHz0CTV1i4pfbIUp7p4FOrFcCXLX3EP0l+AuM98eZfXb/Nl+9XsgELfOhoHo2Suxn1Sr8msUpIr
NXq82+trL6hOyaDtcUDCGg2vX6JtkIJvGg9TtLtqYSfbOZXdWFcDZxMhhB/T6NhcVFoSbyLa8AEj
lF7olkTj1ywT/Tt7naucIy8xUAEkc5m5TCsft810jSEmPTsbNx+p6PbQtVPdH1iIU9vkp5q6rZ+z
8XIii2YRWo1GsWRvmBUDepxHM2u02BV9LoHYD87oaTy07ZYeed0KsqnV/UNHLrXTePmrA4AnYqD6
RZ0aDb9gzTQLlKnefiCf9nr9gZYCM6njU647QpUa0V1CFEEftDVJhmRvYpIrxnEl/8ERWsbACCgF
0oHAHKVt0/CWwR0n3P4TSIdyO7sOpA+ZVImSw3wsi4/aolpRu9zP6V0/XkGOmU7/KghFmkmRM9Gg
7PPNozFW50GJNKgzyLdWbpNBskiYeX2dL2TZoblqeqnb+rQtbodMXWZWhow+D4yVOUCKUFdbINyz
pcEfWBxnYZBRxAV52CAaT5m7JcUCw69EdTkpJrqyRJbeRXJtsQ9LSOoIZk2147Zu2dqKV1txuaxS
+GG9+o1NSklsO8EX2cb4Zf7vbXMRL/zS850PdvMTd3KTy3eeUyBGte4CoVY0+/JpE7QIxr1Qpy+O
OXPPCtfU5OZ68vIpmcYq9WFb1uFGSQuywMFXy+aU2LkdFVewO9DLPfYO6hADEAeq7qLfuYHxIcic
Ljf9CogjzAJ6LYDRATjy0GuJpozg/N+D6s5Y1PG2ArfbNdlWUnjj/3xYbb1VrLaspJgWhHlLeVmU
tmUwLj3Hrd5z8C8jWwHbQuv6riSKN8E/+ev1ZiknFIrSEkI8S6j5Sucn6kojkxk0FadK3Jpbrsko
5hMsaITY7K3FXOeWXZeeNdJuld3Vkk7q2yyizBopwlvpwCgFSgY9+X/Yx0cKlQftWCK0kQz/+bJS
nhdJpIFCm0JUsX5aDkDHFpJnLEbEfo+tSmKUrKIUrPyKeXddI9IkVsuW8iCaWq3zxCqlSnhBvnPu
3sENBL4zQU4iqM1BEy61n8xGlXo6sMWSLOTeIGUPRPcnNxcWAaCiboJSUs4IyiQ+PhXG8ynJ0ENL
7I+o4PCDXSs64zS7nBZppiVwOmrIWpBXzTuiEnLrwqMQGRJ27mkrMUEjvXZTM8MUikvCJKFMKKn2
RKQ2/0SKiVhAptmJq5O/zbAr/l4ZE98KrwPRkh+Qz28dxJfCAv8HAQwFv8WbKkhBZaNjSLmA63cV
sm0qdMhhfVimcjkmZcM7FEsDZxQWX8FStt5vFDA8R/8wF71IzO9Wty0617KziN2pVa/JtXyi4/gl
6NtxmVRxEetubkywAvwt2/YuD0q9dHrswRRQi30U45gly+HQ67/pUs6lSumU/jS0qirj6t1isd/W
PYUKs9NJNqC7JRRv3564MG1T42oCT762/+/MdOJHc0d2xwmDPFvyHDMZlGfq10FqNSJC5CVYl6YO
XKN2DEU2G03VSqbTY7oLdHexoWtSIhffU8t9RrqoKHbP1675hYIq5+vQXOdLyASJc2NO5Z38FLrt
yVCuo10LtX6UCcmeWLvRsjrhaUZuChulSlkbscW/6BPdkVThoclxO7WLZKMYe6CapN02S+qVjQqr
qnj+/P0p32cy1z6LUDPTLXcgFxDPPhS5uatTSG2vNSIoPDFA7fUKC4qzjBmC/jIiws2Oh+rUuGIs
lML3BkvQRMfgPM/ejsIC/dZRSawoknyBrtiloVzk81mfoAFL4WZQ/kdCv68TCG1e+3o70LpTYIIq
01LweHusl1EipRezDnVkQSwzYIWtNokAHlGuSeGF8gB09LjIzNMdGs3OsSLv9vSidGc0xyyONnor
ZqDhTILTNlQck/k9TEUI6lfUgrzQlcKqFU4fFfKvWW+j8PrFOjnVk/HuyCHyXf+a57iRTM+Y0wFX
wbrangkqlAMG1VCBM/6G9CSKWqghMFkGVQ4l3WGVC0L/4zJImwbya1U4hnu7x5Pb+pHQUAiDmvhO
QS46vO3Dcu5c6ETwzKOorTZfI4umSnoBUmzfmAkHN0hX9XSCfpx3ATPtwPm/2bKEopxQ33agi5vR
Wd2sKYLl9cwgXWKtMqqezMBApgLR7v00Jam63DyucUVRcpfQKamS6FYzV0mMr/U+Kr+2bxgsLZRM
gW7kZx/qZoSmfPO9Zhjr6AbfgGgKhERqMOTm9dP95NQo3sGHTDvgS+urEdTPpYY4jEIg/bKTYOg+
qOFLZiyzirZCcqwaXnXR+3sQX3i7Q88DHGi9R9sqMXntW53TWwxI7Ldfh0zw/yo+w+MEXRRNUPJ8
GbGLF+e8ap50S7zgUwsMlaD3Oa8iMGnCmnyMUm/edZ+s+MIzdc0xT7cM0SAv0/ifC5vJs5Adj6qF
g/fLkdQ6P76pmV4MwP90Ggb34KnDvqnTeTygI+o+JTaV96VnC19zxuq9CRcFa0+jQA9FUQXyf7nV
Jswg5GYhGbVvnUqngwBSIl1LXYN7+AzQN6m2YOmhxRWDeAfblRKjGFL0zo/gTrI7JhjYnO3HImqi
5/GHXAfl90YTJvJkQwbtvnntX8YT/22ox68PJes/+OqH8QHK+FLozxez1/x/WdvsLth0oZZ6iHUj
Dlzf6vxukez2cJrZy6XYvOblJHX3JN3MrejgAwk3laEjftLnkMreBhgs1/+rRuv30IiLSTPD2BKb
7+gmXfhwbKupp+z9HQlL9dx2lszEdVc3Jm0v47dG86geyGHwfjiYA0UrxIWJpXxEcwQvHr+DD7FB
BITBUnCoRac00zPValylnU7GC4ZcMG7HrBXfgRnfT4XUPcAIDdfhIWkLhYzF0YPBLIliK5cOauVn
NLGiLX4sxmH2mStBht5X/cNXJFiljji6I+Rn3EZBdebwtm16sXoq4Dj//Ne7//hPBvzwpGg/8lUK
iB/3PSXZPS/fc5l9znrYwGqjJ6zFKOHRBJR1WggmkwER55wU5FSmIwkc60NnZ7Ax3P5Pn9Bri+3T
j59CNxlCcsIatqwy/6aK3qsHHau/rRxHbj73Vm7BAJr82VtkffISAqOa//Y9B/Gl9zJtENIGUAoG
KxSfauEvvgzWLh+9S1IjJ9xX3UqvKL2U66A81AXsjp/8wgl35SVejn4UyVNsw2yGFOWTzy1e+Iv4
GIEHaOVhEbZgKyT2jZLLXKGrw3yIZMPWaeH1nOHP+Zgk0WgwHgmXUbN41IhHj8OUBjvs2QBp8A8w
oOZHNgHl4fD9FLcPZpmWkqpWLzXPgSeRhoZUPR3zcNds8tYtx5Ek7Nx/K3kI7L7E5fSeyheDuZUK
VoiUKfDir6MxjReG86IK218y6y1K2ps0YaIymysMIyiIK2YqOXriJhqAOexZTpJKZR3xxlNu4CYe
/oh+vWKOQ6gYfhcIVJJIER7NciPNouUh4KoM+BDGsglnyHT9wbyMzqSDJLjXr73lFLz/2+qg73dZ
rYIiEcZoY7Y38VT39Dn7EHbqnnaGqYt0cdq1TKUlSVgA2FoyTUyhTHPqeLJgaJnT4GvkSs6Qgn+M
936Zw+fHh+gp1twWydWOF3+TeHK14MwUY8PM3q4dp3/b+vWAYIG2XPEkKXFx+E8JQNRuh0tglv9E
kps0LHUlaGm/TGZcEjiuQKhbRq+SdYb8vf03OFfaTvc2ofoe5PI9bVgY2DuEQvSfWSgkTaA9t9ly
okh++Z7UzV4GmnFf047+A8dQxyCCAfEmX3zHLHxadQHXkJYBVaUCzNsqPT+QYuDjES8ioA+j2+W/
Lpuxopskt2yGIJOZdehlMLJT6VmIv+x1UcW0NhnIeFjefRw1uxpY0lljQI+79Ysgg4t2WMYKTJdb
CtkWkO7YBN1sTVM0kEr9+b8Oc1bwBAzizuE1jsA2dm0h+kaYM61tySJTaiWRIqVD9Eo3CbV0rgQ9
Df35yGqPzQ3grd7RESl0JeO5lFJjTgwJK5hrrVSbvCwHrjeVyrQ2IXHgXgYFgnRhi8jWDExycd2r
f7+Nd0G72zrOb8O9NJrQICyWGpF2UMtL9tV5+906ZW+aLvJsGbBK7tpHHJ78Cl1qq7MKgBubBktJ
2FAAqTUWrHgyNpyAQCozeyipUPfrzD1KbBuJMpZ+UfF3aap0KNuPhmGuEo1+rgPun71ezkM4Vw3/
8N4jPJdknbr0jSu79QgmkhECqv7biKeiq32e8e9dVNod6FU57dbqODURvelJsNmhMtKrB1f/Eg/z
k2/zRdMD5fRfHU7FziyDmPyoc3xZaMupLAJ4cO3ORZA8gBGWQjsfZwIDRMqY2XM+1d75ZVMcslgM
4DM4vbPbtdyTpCORHJVkKkUfCmNrTR3dnUtCGcnMlDEJ02FsPlVCqUCgUsI3dZDJ5FmqdvjXjiRU
i3DBX5O3VrveF+RHeX0PYQ/tJQwZD+ZMuFHlND5VllOET8bqMtgXf20ADbQU9qKo56JtwCLHNd2/
LkjYHqe7JTjWkniToD9KJ3ZZmosp/T2BYi8gTxUoy0L9Roa63zlpYu7mhpW7dxBnNNwT9f7ux4NV
lGmt2n+7cslwzBba+9Gl84I/ketW9Unff9JtySiKSgzSInUwUXHZ0GvyOueCLMgTPHkVmDJxZ9wT
qS1rxz0N81BTDkZa9/+NHOVCBIQdRpw4bSpMPFmMIvdSYoFltYhfQTLQZ6fRss6sqI6M4BcfN7wt
+ja8DMU85R9YgdN5AwNjuQHnCUReymmhb2UOdGeSnQd6ZQCO2Ti/lknt3KIy36QTgjyD3w2OjZR9
4HNiDcrikfkUdhQKd15gCyLmbfv2PTDOafNxImfc/mffEuGPZweaKh90eM3GRvxSnIoj6UZ+rBYi
gz1JyWK9ErSbbIS+GTBfmalpNWeQESwzHd5NWxhAqOywsw45N/dAhcWmgd2Of6eaIU1nhxoyCDbD
G3t49vz0kR12QqE3ikPqOLjT3M3MbLmitL0v4vh+6LPwOQUX7ELJgEhd++Aox435zXrHnT+kTso+
gi9vXTY8aksnmDaU96UdbpMK4t7vp5dE3mwB8kNfgWxAKW1/kcuF16dcpSxGN8jkcmFfmrQx0Lxe
393gedKU/NLT5tmC3n4BizjZPUHPBE+/z104mUoxRgvDCK5wpvoMfhnj6Ww9hoAg8pwIi4QGhnNV
R914AowR3vdInK3/1S3uoZFA3gxgPLj2LkAfs0gSVFtIc9sqnnW8f6seqDRotAjhG3j1r9xErZlk
WEhOjADY4lnaYPOnbMPC35SYetz/fppDfdUsQHqRapx+NtOPGC2YzcxhwP2CGkrBoo/6iXPuwLSz
/YexeKVVB9UBHC5BV9Z7XaqAkJXPMIRHdI0hMk+gukQq8G/t5jDZ57cbKY8Uv7h0C2COYcytqQ26
UnIW7K/mhDMOysn6n7pCu+MHOJK9DQwSRGJl/X4jdDhJO3rU6kJMvGeu6q8cyLizRVLJ36nKb1KB
n9U5aUVl1iuPecEN82SJheYdOiokUw+SG5w4qD2KYVtcWCmtXrAiO5Gm5mrGbMyDmJhHvzU2znNy
qrEKeGrGEy6lgktj711IQSxCWg2yA3U2GZUazjLMl2TYIsgvvK8vGTEYiMfPOq8xW1KzAt0hoxT4
QVQ5aiNQSVaHJxnR6JKY1CpryvfqLht7J/fEVlMzhApAa3fYjmS3+24GFabkXm3ZE0jjLtzwAOwg
o8hBTbdo0K0h5utGQCR+qYor0nU5fzhok2C8cuUn8Ss5l1zBcaqsAJdIFV0W75zSP+OkRic/vZ2x
398PndPsVVz+3HQh6vCjxxp5Of+zCOfumftLOZhH9QVJtLHG/BDWM4jdeQYaS5z7Y7lVLqxS3Nz7
Y7oHTxMuQkltxf+LJ8z/yb1w8N7GOVCwsesaVMiw5uEGwnyJls/9Azh3sph3Ymx11kvFOhye319c
q2l13v8p4EHI3LjGssMVfd2VhviO0IGAzWXZK8J9g70zX/tRapPietu+cJpj4XqH8ps2gd6Ao5yr
BXRUZDTdhlEfPc4qtQmsLOeCcfLmOGW4TEPfOyRavla7TJsEXEfRzVlsLfm3w76bizTBIpWSNQx6
rRGSWJvNZDpOyn9RdTPMM2anjz4PzIGhoGIdWTmx88wCX6H6eQwxG67DVB0mExVMVejCzrClD8CV
x+XcwBiFEN7nMUom3vZ6y9fosGPSpanZ2iL5Zve7Sfx9DB9vH2nryeBTjfqKD8nFuNxk47ke9/b/
/TNvNRkvNNpiTxLlWLBn/W+lQ4Gld9dLNb4P/Kj9o1eiXJ2cZns1N45g8qpbCSIrvWczkg5fLIsp
P/ZAx43zYS84A0hMwW7L5FyNxrqIZuR/UMUO9Rf4Aw6bxfVb84N6QLNB5VMCTY4tUFZE23rkSHht
XaxWu3BYVpAfzZ0pAafUJFwQxrbFMUpKYcifx5xWUDm0Jmu3dLR9ESm3iAmTvRbiIKtRLPGp5+nd
3dUvfsoOe79JJT61lJ9MGoxIvwTG+6+SBQarJ1VP2zCzztNjH34zPP62I3Vd/q36hJ0bjxqP5LGv
mUKucA5mNFpy2iIZ376iQzJNzwvoVH5CK4TACJhC0oTMkFimhhx2IqIGtkv6oXY2ubQY/mvyz/EY
8xEKVhZyOiu72xboFmk6UcXP6KQGYWXDOUQJRakyrxyPGDw6yP/HpVCFOq8GFU/Wb0lROANARnXO
50JwUH0S5HV+uB+BKI2I2WzB5qfs6bIgVA02UvZMdfnNPcukHtiL3Q93SwIJIeol6OmT7N9gi8nW
KmRoXOWyV6SHPykwcXSEzNJQWBGTStlXzuFA/3YBPjXGpWJ4bHZO+8ZIfp93Osws5TPXwpfROzGn
IztbJKnwCle6d1GF8NkV0QyFqqwygg5//aqyn51+VKJx5L8kE1/cud2Dt+aOeOuwyunlZluRF9aJ
mOHJbyOLRtRjFQ8BCCNfLjyH7fuNYJ9Z3jtsN7Gf254/LAP1jY4//G4BXTlCUza3EAFsogEPuBDz
rybzCALvoEJz8PkvK7haz2FJFmYlDtaHMBjLWqbPi3hDq3usNJbo30ba6CbbM7OIYQK9BnL+0ofL
6CBxA/cd1xS9qu5pNS7/yERY1y2yGob812ddCSYhnZppQxOYoGIRBP2rk8zkwfjSurJjVTPkKAo9
YgqWxN7Q/h7vFBzUTBJlkTWR4jgKrBaBirSstCYR1I4rfeYranhV8TvMKAHzFUGqdE90ULfjvJK1
SWhEPnC9WmabV060ei1A60co28vF+hqUsX4DC0zzGV6djK27jLeIs3OohSgd5Np1aL996ph1IzTF
uGFHEt3xCNTUPpPCa3dlIlGy6ln0xWkKcEOdubMeOT/PgwbNm+yHOXbxz7W1um8LSnwYbxsrTndy
+HkVV3alUxsprf+BYP7LiUa6i7R/Agcd8zEpv9EPrHsPJ+oAFEqRlFTP7Nk5d6s8w/C6QBc9W5zf
o3k3zoNnKTMG4OkIdQUzzibgqX3v8WTAdt9TsZuZvDaAy8XZ0Bv4s0I9MNbSdLbGfzWYxn2/gcOz
XW0w9ExP5NBE7U9mFgiyfMjK6DdmtYnORHZPcYhx/vHFZVdhz6YQ/NffyQs1OBssP3x5V9UnCPxB
cbM1bc+EgoEOh7OwMBBS23B1fqtYQGeeekW4e0i9Zi9w3l6O1yhl8M0L3ZfkDfuBjhAb8IHrpUet
0bOosmyGz/TUjMDQ/Z7BxeCIv/R4i3b1NvhtIYgSo2mnaPOqpuVYGKeDaKxPK3ozUrc1OnkSzUnV
1bnfK6SqcglogxYHy86PPl08F27Ql8wQSuQcSyAfLiUguMzWS3R/zf49rn1PiRDvkFnlj4RsQuWQ
/3LZzedWY5d/PnrMsdza908XdvNkI7oM+r5MY3jj5YF8B3NALwKICyiyJ936ospiEAFsnFS3SJV6
lzxaOWqTm4whntVPDHsRXKPe/SLmBHogciBN1xIrFu/ilY2fDSkDmWv26iUHT7PVQdgBHeKDblQ1
hkvCSa7nyPIr3mRjTYLtMTyck7s6QFjFgF3fvuV1p4fKs97Uv8EvhWYcI95Hzmh1SVrpx9cOLfpH
CQs3fwGDvlm4p69NRKhcOlBQGtmwqmcRCBZTrEgl8kto+hAByS3XrHBp4rk7CQV3AEVpzdIl0EJa
WOisQiSUPYQwr4vxzWMlNAML7A9bv1D2u4gM6PfXvud0I2Ye8qsmZ2aHyc65qOAyH8cWxU6NkQFg
9qbE3dzJlVAioXj/61t5cQ7roAUIC2h64xQFi2h2btZkwtU8JyLnKHg5VJWJd8Dt1Vw7y2wBnbBs
TgcGNZVGNCbVADC7A5vub+fKWD4jueHUm9Mll2swKGsVgPBq9G8SI+tma1U6Wy6DQncen6crln3v
6AeECZAENYrXyRS4iMaGAtQ4aHuxzNZo9FxTppGY1dhJNwInS8DHOFuqREZwMaFvYExvTZuLlhib
bK4je69v/1vUctEryi+sxMOWCvowmx4YxVW+2M8cgHCVUdyNhzmVxW8VzYu/DXoun8B7MP9frb3f
I40PCdDrurzBqLsk2BB29tkVdaciQygF6SA/3oxOgzA8ZSu7m+0zrAr3oHP95obYzxR/of0YnDxa
TMTUQ0/jdN6zNvu+czWnDMd0OANB8uUQNNVFD8HqLCTvIVhaML/INdba2WI1wGwD5Z1LemjOqecC
agnj5PPlKMO4MI4NMDZEZUyL6Ir6/XGXIVW3Rj9gNvsx+dNldraUYdjxXGVpfJtsfeumzX+nfI5s
wDPCYi5Kp/gE6zFFjq3e+LYAxiud7yPqG5IHiot8Io47B4fKId8hgDV+HjIUPemWdL3T0U6OjrxM
TIIjMF+fEQ4SPyItfYDDLl7/rv73X05XaK3VmohwlKXqR9gUTKPvHccMzj8KLOj7HukfKGjFPbuu
MMfIE1yqAGVEK9H1gjx/5zs3qOGW9/6H7yO7VPYk06JbLYgPpRQF0J3gLKkJamhLebS9+tPnAM5q
em+zBocMqMGUXMTuS4ZjhzwFahcdmVfumilgJE8Nj86+1cL+6lIXxyaNHJGVWuPdWnZPYRyl5yri
YDewPvd0Bl8GhJQU0M/xVnhfLNv1ytkFB+0P6EP+f27M1BAzlZEmt1YLChd0E262hpHT+w+B8+7n
wUNFXV8fR21exrzAzq9P+WeqAc30EYLsOrow616eibJCr5Hcrr2uAD/rytaCX/DKK/hcNf0I5iIF
Yv+jlpddTpqgthyRCtWqH3LwZYT/NnzUaDBeEadH5SrkVuQoTDBrHFTCqT2eqb6tGgFpUziLpQBb
k+lZ+sfo7t6+MsTj1HCsOyYhbbWlTZFNdvNENeHNQV2FuzgjkrjbvYDdrXs6vyJRf5ivnPzulhIW
MfrxtEi97RglckSOrkO/ut9K2wvstktW0bUutUD76m7eTfvq0fIiQ3774gxo692l7hTIEalRR3El
+XxWoCN5z4iRR9hnWeZWAOD3sb5FVqJ2ds4fY9gT6MTEWrUXI5Uix0wvwBoWW0m5OGwKr4vhn9Sr
T65Lkq5DnNs0EiXhyIh+ennT8GNz5wFWpZF4DOM5f67GK7Ev8ruZdrOo+DKmL8yuhI5bi0oh1Rs0
FaIwjeVJFQv0wMS54nerrQYRSC7mnj6PWGwAh4p/sC7RijRzgAnvhA4SPON/uM/oOOlGR8qLYP+o
qFRD1GXlG7xZyvRZLYvKxIavO/KUWdEDiUvD2hpw+CFVnoX/aiTLRIdkXeg+Z/Ts/K9ALM3CcaDM
VASaEJuhepCB7DOWEtq7grN1mTW49CNf/x1XWSCi1qy8DnNNWQPdCPkOyFc004WQXpSscF8SfIfX
/C7pt6fqKI7d/hf3A8pWBAdypNWY4xjSkUuJ54T0W4xYsqVEB1ZEA9sbHLtumTrTAtAKdX47AKMC
9JU0YuYRCi3q3csz8zjTJ8Xz5o4YHgaUo+fl+V3N/+Nd8eVymgk6bJsXF/5IKmrUVB78MrG+/jtE
SNHAjhR3KKl083THkQ2HgnMMR9YSE+/7r4EiR7a0R1oBthgAlVnd88yftd5qPFtl3hG7BIGX5Tkv
FvWWezFr74/8/kFUVbV03XPktzTNfi8kkOLUPawj/ppp4Zoz1nVhn0IojbnwSRgtnMybGaXQi6Eo
GlLgCpVkCmm9yzZdtYUG+zrTfF4mQ1MwA0l9A00DJtjXEUtGvnL+qqdsH08poRQ0Z6mGiTCLGcVJ
hT0A3cBnGJ78JkuD9ko1rWVOPdq9ks3Rjnz9HJ3/4fVy1DyVxsiAbIRjNAaqKFHYthTAA31L31OB
y7A2ceqDFL+F+2Ct8kXpyrSSbDV2fJBQg/d/tCASYLxP+U5T0jkyGO+88rP5H94LqnDm/cw7zZJX
2dIPMUTTS748Ab1lvg6CfmzL6SyZgBzYItt21KAepIg51413ArtMZJmyFjwU8UJdNbWYNw4NeIJH
7bNQH0xBy8uX7J8Ev83XxSwJsA7VwQq64NcKBumtxRStdmOjlMJ8Ml7bIuQP0QNI7yAGo9RizSf+
By2/ywhxqpHJjAuu9nOz30qNHlDpAPJMGH0QsK62lYDvJEcdceeS7s3f6/JaVADmaLei3R696mVP
td6AOB9Fhq2Hx+v46g2aXUHOFEakrwrDVuHND+fcGfl8VdY6o2VBmSRBwNplSF07GLqiqe3cNnhJ
WrNMLyN973WaLcTLaOIm0wyEEEaL2Jau/NnSejIPHIva9G7EqwFMyHS7ihV9lXTW9Pf/OPI3qBVV
CWTSDRNTbJcEOXC0qc5a9RAXkwX+XRUs4OhzKwoH8Eh8vf/lV8GogVXGcwRywFwMnN9nFs9KyjCM
s/bkF2l4SnQo5AVLc+TSxmuyMo4eJhOACLh4ZL1i2xXTKb2Fdc0k+yqtksyIyOI/et49RdHTd2dB
LUjowqPb0xnQtmE25Aqt/hRjuIeyojnLZxfsNKEBcD1zeNU88CWPvV9hMtnyjzBOHnZG/fzoCUIR
GFHgrA0zEPOlPgpmm3qKV6FTm0E4Z7N5lygzk0eGIcfUSgLEiTTQl5p5/1ConJy1CRjGpM2UNF5y
ILq514jmylwaP5BINqVdcsNEqQ2/t9Y3LWXIMZQCU1MX7BGdPNobMwCBMVWIjyw6TWgSXQzl8iCp
PMiWq5XoJ4TBxn1xT2scoCYKFVdYAHCYUR8iiNbR/1esQK43QXvRfkDTtRTe5Dx5Tis4J6tGXUlu
w6q1/1ArczrBCQ8afubGWtsfJXV6rIEaG2ysXer8f4NQZywt0Y53L8hjkE6jjrjKIn2Ev5Oq3DpU
bOrvr5jPS4zNfKY63dAbggAXKKBkHvBcuoRB6Ui/ayWGXDRQvgftZ9uajSdQrEOVfZmRvjSrq1MJ
G99+1zU6hR6RbS/ILWzyqfQwcTpPGjZa5nsnKwLA/MuwYKLTe13J0qvdRFgtch6AlW33HKwnurmu
s2ZLaSX/+LXfGYmdRf0vvurFJ7w6vc/amTK6jud1Ko6YM/BiwgBRW+VPf0PvfAv8faIrbGAhj6Ol
MtE/JPWRd0w2IR3sMNKadrg+kMlXyz1ica9NK2G6lNhVFWTj2PcjNx8qGEi2PpnySYGHyJeV/9XJ
1t5nOevyWOZ3H1zSrIpK0Qyh9TDn9tSRxhaYXP/B0A2Gz4ZeSHhqfObW4FWqc5+2RgL941tIcXO0
50u3eBcsXqUvEbvvxeYxCQYRPoXqxv1+OCkAoIvF7SRGuMZBZxsfAcU+c38Ur5Gsn+fgKuG4cb+A
13BO2NyX8Hsh9kFmrxiyuujAlCfbM+JqITmDlWGHJ8ybnF04OJFIR+Y+GpCzDElt8ng8aa6NBrlm
lGFhaO7W4IKy1N17TkCampOqTAyl6zJMQkkpYnSXABMgBRhi58WeABQM5ihMZjG8xUhmLXUe/COj
i+fOd4jljgLWhvy0drEQpHTNtS6ZPEeOrXcWtNdyWBeAj5ckf2Q2egMZ/Ci5cGBIY1OErZUwav+O
fx0/E/JeA8Jjdlhwqx/1F6UmIem+LpTzibaCwvgnTCniS72MF+eZIg6UPHRDyU7ckeKcY5Iq6a3g
lYNgHa1kxL89o1z6tfDhJvU3vPve7hJOUZAqF3VC4LFlhTKlIL/ry83ZOxEwJqkAE2PTSJfM32RE
fxtP+srzFEPs5G7xFCTxgjzhPEjbsloI5+VZUm231xKZUn0G46um93i893ctLJXBw68i+UZgSIE0
HLyYE8BaGOUFr0JxVeUzOOvA7tHE/Qj4i6EHFwasPivGa13ZLFWa9m/kYt+k8JRwzRU/t3GJNq1z
J85IDWHOOiDyA6aRuTuPK9ccs3AWv5mDeTW/lEHLCK6Yu0FbGRRo8G6ke+b3YhN9gAQe5UoVmvZd
a9ueiNqBlMO/BPuOn2EK/Gn4LpLq0Rmn/eqWpSnhJMuJbjOb7b2zvTbqyliBxP20khHTnYKGS6O8
z4zrmYEgyGs91FDGt9HGPNdezfiv160jhCbROW4ImnM380D3yrJUN7Zp8uuZJZaR5f7QWIDNVeK6
QQABqVKix/IvES6p7E1dzXZ8NPDx1flzHACZ+6DwdfdAC1S80obNLu02GV9YwBo4vJLnkjggRWwU
q3vwpm1DojCw+IdgCuPyx1JSePCmPwIQUO0968y47w0HOOALfzx338TAH09UeOhZY4kIeYNRAWCW
pnGuPCqqpXKGHLKMzPeK/4mp2jJA4E/I+h6LiKbKnfwlpIYyc/repS1Wwf64yu3e76dZzMPPH2lY
8mar+4IQ0PeXCPGSOTokrrzHa3XW3b5bPYuC/JvRbxO/ZIwsB0Xsx9aUBiG45ZMV0afMUfiTX/vw
tyMVLprFJ3sTRejvrSPvTzakWYv/Z2nZ2GHWx9klyRDDc6FesXRMjco12KysELcjmP/PV3gzJWLN
lF43j3grYt9CR2eVOoiQ2zRHGYMU2yi5jIqBzkRuESxvTWvjOAzH3LGmg9AwhyMAxZzejw4vpsf6
234xJ/1Sr2361EAHgg5yu2viioNPIqyLRzKWjKetUsOSm/ZnjNBguAId2BLred3CHDz79mHDDMg6
KACOdp4FXrvTFNy70EQiczhO4SK5FNyn8m0cG28i+7ISEQv1OvVggWH3pkOEMsk3UgFLKr+Mog08
UsHnn+WXphdP8NtASMciquVYUIOlw4242YVR2bxUFB70ROQEaee5jEmu16NjZ3TtQXQTZsCTX+3I
T+A9vCVF1sXTWxrAVFVqWmQ7BnsD1+D0JOmCDGNngAWTZ0dqnLlNZwZ5jq9HclJLdnxDCjVajiGB
PQxOg5ALNAgZDcIkoIjJPmCBtF17kkHB0OHC3ACf1YHesgIeRGvA3pHvYONqGJ8B3pa3wAZ2QVyz
eQ+TE0vxhP+3LiKtgO5ZuOd9l+vg+XM7VkVYVETQcV2Nb4B0VP+ioMNAR4llVOSjB0+zRxvEZH8n
uEiPdphqSJfApyca2WFwCMBizqKzkMqbramfBGkdPJ6who4ey84T0GIMEqze4zmBPSiS0xCpbKQ4
1ybqlKdMQtI4i7uCJJ9Ps5GzGW0cQo5hr2UD75d+Eh7kI119qazUROY92VEwGY5KAPLmj4MpY1/H
Q18XwV4uZMWyj/E7P6YJsVfPuKokqX4OfvfdASA7YWimJVhFwfxG785cEgXVRotiXfK52ZLwX7Zd
TukxitnicU3MzxGAwVdwLKPpm/XEzvBj3UII6ndLpJeJqOYxbhGHB5KPPAPIPSLx6peGJY2UnRUw
pe89Qcb/6xKrHXL0FXrfznEZtxaFa4V8c25S2hA7UFQTUCkRVhZB7YWUEG/8FcMq7uHISHRcxGf/
DWdE2mUL2EQEwsQWuBMTSuM1yv6qjAnubi/Kkgo7NRVpbZiv5PeG938pWf76DJu1h8COiX4S4iSe
VNJxQ3qv0yEX/BXcQaZKZ8e3tOkkvscZgCCRUqtXNkfGCfpcEGqyN94as6No2I2WAo/UXQddoYHg
NR7e2Wv5uqrBt7lzW0blS5a0cfsZ0n/3N7TnN0/YfiqCpApAi4CSsdFpUATAgg9oBdMuNBWwA0vx
ALPMUj5ESCwDsUsz9Ov2JnCUIUMbi6EcXGYJZQ8VyqO69aJMqnmPADTVnh1T06X0C4C6DY+S9plm
07qvDeXwFx9Uokd9rV5hUB1MyEJ9aK3shQFOHiSaip17iFBeEfey9WDJBESVW2aXzdgRfMjbRfXP
glsytm77Fafm7bR2Eu6FZVE0TtIKFChDaUZCSiu0vPAFjJec1HwhTu0TD2SITlNmGlMWOTCaRN0f
GvCyBB836K++zQNzltlyh7l60TUPRVTLsgJYMsTcQeoJGoUh+IeH/m88tQp4QUJJsiQ/yk/m0mQh
4RnOsA2fhjkRxDfw0EhHLYbxkXQqfd/YKbOSYE62xt6kiEWsD6jdZMz56ncZNSh+dtk8bbWy4lai
1YjX667sua+3dZHZ0KR32Fm8Y+dY2n7wInwlU5yAoBmvHej1HfdYe9/NEvozogM/XpK90zdGzNHa
0ntLxIU3yc79iuFqUbPqeFnOdCpFbquUQLUc1hKm8+j1pYetQF46+QQnmqLjFHHRsypzks9qy/XJ
cSFzPPn4o/UobdyEpylPg0FXuxckoWZ5ATdtNWX3FYd1pwSvUVRDFKap7Zh7g1p8CuVdO5D5LAXx
bjw53LmaL7sTaOTewLcOTlKm3FWZ/lOV38BXLCC9IN07Ps0vP5jYjDRr60nvoXe9QR3HV5gPkLUs
KsVvLcqeyLgBHzsexQXIfXgeeyavpg5RjdASEI3rAE4u2bh9xtO+ODJKOao/xcHq9fGmHsevbw2B
V7zHz6ivUbqLogoNaBvB8CqXLcl9cDIqezlFx+a8gxzgJJOuEKJYS35rPAMwQxIKqBcw8l9Kd2zb
ULrXhxudHOzQiQEg4tTJqoSs3x3u2wypHsixma6ey66yqHsbfZ2bfNu/QFJaUTv9lngfk44lI6Y+
+m0STNs2BX619YevgmrJEuxdO3xeF1L8eZ4hXjMU4dRS4I9iVB4yCgxER/kbOqCi9ATQSB4GqyHU
ysMDi8u4BeRMLOSMqwRxM0bR1ucstcIvGAMz2S1LB0nqveR8IdcEuMJIv97ebMcD1kIGxxG7Z4bd
tGiScF3tyHL9Hg5bxkWwdNpWmLAgqJ0hzJPFPd0wZOeRxM6W+rMKLog7555TbosgHFJcVg+eWYr2
1cGALuchUgTbtH1ew9FDnXMQ+qP76z96lgexpwgTL1SNsg/C8BSt/xd1SVlqFhclViCY0SazYhQQ
E2qulcSDpR2OtRElLEwodwia6tjCbpCm5A3lNQ5Ig6wLlJ1VvGTsNoHkMVwCgNioAdJaQGLhj4Z8
C6Y7VQUhVnlv5Nu9PGbMbzGu50QWt6IpoNRscSsbMY8QsfVDJkIyxWs5VSJXcIKFkEnHIzEvPDYb
6+cDo9EIqU9lLncoeQpCMFnZ5DArWJv9mlQ9bSEbPP9h8i8z+K8WPjB9vyIjhGpxWckGKcbnGmXN
5nc+DZsXigcsUYhMswo1ac2kv7BW+VJ00lxrFJdpUj5xsGHnwBGHM8vFNnbJ8Fttf/5YD2nJW2Wc
DxW5+ZWJRcKaGpRa1Gf5Cb64XdMTyHSyqHWbIS4NAXhJj1dTpXBHLHh/GYPf/3552D2BQ/E5Fy3/
To4P65M9h5rGXk2Qa3PVaLsGnur/P5giWZZ7IWs/3FHAjojizqu57Ic+sF99Z3h9wUEo72VjOAmG
xAhJo0S307trMODaE0NivpNQTZ4h5kAx5RbTJkE6jDGVI7ICfGQ/uf4xRGdI8yZEffX0roBVmOXb
DJiC+p1jxYL/prIIhUvNEPnJBl3/3IPJOW8C982KPdTaCJ5Pi9e39eauW+JToZHvDKhofnZwvDtp
l8IVVg8ya5FMCZAMVku0WP9uFgkdD2A2bnb18Lj0cMpyFECTrl8/s5uPznvM73iwMEiO+12nKHe5
3k98llSyl6RIarL6KBVHvnS9KmgZJJs0ClSGgxe2lmKNR+WR5O/Bc4gx3nyH1Gb75XLPt/rsx3tu
9OKUM8lLWhax+EoDiUoiOa9Fmcq/4eW9QkvDSFky59dKFnwyhsO87JlHD8pWU5jTiZr1DRDI9wak
Xqm7G+P/3mcGjBTeYYbEDEgKihrogGZv5n00ALDBnx3sWNL/u7fBh8n7yaQ2jncMn16PIRrdQt/1
iXglNTVQOk7pdCHKyf/21nwMNG8+FZoYsNZogejqFY8A3hN27pB4glTog1LIUAcaRa2h0LBQwW5P
4IA/e5+qYqXrncF/srF50QVdmjQ9it1KoB0fqBf4HXanjMT2OV7UghH7eEwATIsyRDcDomcTIEZl
1eOyAV8yPBls1+ikvVA9nGdG3vrtlnuGGmzL3e0XSuU46G4QOGAktWKejv0DZGdHBEXsYw2v91y6
aGugI/28/8CX7oK0La5+HJj5PA1wt4PxWsmAwReGEcVomRh/08dzwNf+PVPKWPSKvln7tOwMvpy2
/JTSMKh5Pc9KKgrcEDXRQ+gkR/RCZcO7+qe3Pb/dCfVe2RfJaS0Zs5BsESzDio4bYf0/CtsIi/5Z
baiDexnCZBdLFKzgE4Mj7wQlmkwhJvzbizFOrLohQLgzdNJ5M4uFOR0LGXpS1lTfyl6RypCa3FIi
a5stW9hNT9YkqfiaZwhb2LKzRr9w0HavgFPGjYq4FJf01dfqaFhvRgxwSdabDREfdJmaFoCwfXPZ
idmBuBTeWzcsoswSxWnQu2owKuYOgNXZoeAWdUN55CTJ+KCnJqQYVYdxhL34eF21tKybq5vqvdV1
raYvjXSZgjbZyHKK9IVJqUy/rhcZnC9LqBpB/qbLKCyctWaMWDUufN1IeijTFNTuFmtJhvtjcpBJ
Jxl7A4OOc5X7GQMAVGaJyUdoHEYuuDLvOkaZFM44myN6SaFjdCY7z27aT/oMvhO1JNDAXEvWBk/u
p3hNeHOyX8cydOMF21zBcYZgijfBkpePAoVk4f6lBFs7GYIlrF/lkjT0hcAB504oN9IznmIkLDLJ
7wRD3eEzMK2uWu/J+e5VCYSe6HIpKPuBo4Ux/xJAYqbjz9kya+VWzMlwWo71SRNN0h4cOm0SIKXa
yJy//pX8wIuMtv1Y7GysE03mQX0Ub9E5z/qfy3A3Xz690HGotvir1uZP0ARsDYk3pBP9meb1KD0h
Goc/gGyqh3i3pZaEMZDDM/yO+RrFPUmF0tVvc5bsft9Mt2fyUAlugjI/SeJoa5MPLqx+dTrgCU9q
Tdq1nCao70GNQeEbc0vBMPv1w8Kj/KOEZvuRvQqfIZ5YoWfxWFDDoDjEp57XKyJ2nAcIkErTyIDg
oIirBkv5DO5pFHb35GLuiok3xcSpHGvoW+P4n/2kXQcUiIoVzsv9JonLN8ZdsXdI0YF3y2Llxe0O
Z5RSFQkoslWBReFAuxXfuSKIEoxXNCib7WJ1fIGNzUbeBDodcSFgOiojeSoAZmkzTfJCvDCxP4nG
cZnWEU9SOrQYHvRyGDNwG6pTa+zXoBiQ4TS+9DusJSH8nKKUZ/gr5lP69wEGiwVULeMC/nTo5xyJ
v59Nc3YmJak67lfsLOsWW4A7pdmgmexiLi15hCpzUpnn075/gG6KreCRs4ApeOMPvZ+VO0lK+xFs
ufWYZFJRxJg7gST7tjy/z/KmGyNguvateNJtcaO6RjBz0PaxgdUPr4ApKGKKkw0Mr9MjMXWwJXIJ
bx2b8SNMHNCxcU18CJimTbJPEYcAkxdVykoaaS/pl+jjMz7kANm6F+xnH/vSMeCHyXaP1DJuNRKo
+PqG3n5wWKMrxYQsRqijQfukfYyVcc+llcYePYAtj8Hs+JbuVpYDtRHMKfQPQEYTqgmhoYw7KaDa
xU8LK4eCNzhTw2UkqW9S/6i4SmFMSbpDoVRjq6W26/mX5i5NFFzDWuAIksLHeCaqAfMnwlTUsWCz
gIKGMzEyohx3wY2TjpXwUZc8701r4WOOaP2fTPTFIEkvuopU+KcjgTjK7srroxUFZPY4AbSLDrzu
SnSGKkOeQyoS1LuD9OLf1IVhJV8PYV6W6GWS2LzGwa4sOq6S/T+cILrcmvEFDEgQljv31tS9i8LR
kqybUguMZksQCZ5LpIk+jPT0LerSwhdDmdY3+FQ5CIzsCUOHv7Ona0UTAOzY3Hj1oEfmSdmcos5Q
AlZwzrJ42/vhlbbikmpoWpqsxBEdBDEjfGLK/gbCyZZwaGAl3DXDJsEMQ6VwtuubglafpZItIsrQ
p8Rdk7XZhS9m3ALK2IV0pKjjBrCxyCxMuVrbQvvrC3WFs0FJdEwkPuuVkCNKpjHqsuyHLlXLwan5
L1wVOf5aEs+P43GlHPenHEjyOmOsYz1FllKWpuTEoVB6zaely102OsTpDeEZjiSpENPt4SiQ2IjH
G3ku6byf0h98bzQTjoTkFmWZ1OKq74BegRQZRqCypr7I8gMPvUv3B82Hr5Y+mDR3BLxqA38G4mCZ
CvVD8BpPrpBDZb8qv38eb0CF8U2a1EJtRQfyCgQiQIOAzCf/HT6Jv0wxLVcnG+gjHMpEuCexd+dS
8U1zCs17vO3QU5t0ZUCo5I/TErxPVfhPbTS84K0j+/0sP43vgl++v4mgWV5AwhX+2QOnoADIG+R1
wfN6zPgWElLTCCRXFxwcGFtTtL1rsTFE3cVnEzQ8sbdiprFc2qNuDk3G6p81lVTYfPG6yYTiB7oG
i4HUSw6CTP2MbhasCCqjMVxlVDyClXFIUMNALVwYgVoPnv4xNC42d1GqUCKF6LCB6SP0hEwY8W+j
/xQLts98LnAR5e+Q0mVzKgV//72dvkeV76Urj1tykaPEniIsKa+sarklYKrjsLYM17E5HtuKKZqa
hjMVD4jcUmwKqNjwYWwyZHdmv2jobZo1HJuDaztCY3xCtJXhvJiCM8nfgQ5nidEYNa5TyLvoy0vv
KtAlZJqUcPsyezppjky4Fk2jVcNgwiRBB55j/0stnd6MsGZdAdAbCiZ2fcI6XCcAtSHIWCMzEdyQ
MOgNrWTFRJHSv1UW2rsozeZ2lDxdTsYfrycw5rbY2JObXWJWdT05xj09bybXjuWSSSuKXAzD/+D+
2xinoZ8rI99aAZ49tU7dGjzX0OFYRfd+Nz0fqBGAkojwPVgYu+vRF3OD7H/NWDEzrQzPjcCg2Fg6
0i0Ho/2Vc0DujfwIgf03q05D9cz4d2UHi8dKN4Hlw3oUAL9nE3M1h9FLCcG3dDSD6trjUbxwyy93
LYfmfIYSsh51382jS8ZRBLklC2Fi4tveKa8KBN3ZcsCu/i3HjGEQDLLZQvf/iGP3fNAh4VwVc19j
4LGFUwCZqtVE4sfsEQLdRQY5OHnrM800q72+AfUzg4h561nein/O29D52q2Vlo/5H+Bf7moTSV4H
VgeFsWA8PxByTwj1omQxz7S/CnZvfd+oCf48WsMNnqmaE53ymyGIPRfVjDWr7Po0lddW5GUSl6wR
KPJslWm5x77zKzluzqduUN3Nfu0HWtkxGq5JqUSNg5w60+fWxDibwne/m/f5kP4QLsiuO5S7GX2h
iqDKTmYh0g3fqo5vBXqBXBLYI6jDqUXyW61B4p33EzctPwl2r1pteVpLlpUr4gkB32fjwmnGGKrL
z6YpUIhtQ6yNjZGjvBTpypLdRgLt7ZQv2vCl76hjmF3YL/Yos/iyLsfjHY6g4gappTGIBkJVt/9F
lHHrd952k+ANTSm0eGuqLRJAzL+56UUygnMjLZHl2t8dElyS2K951TwrxZ7nSG3YjfZZVQBy9ggX
swJQQaymJPPrQ1zmpsFxq0ho+f0Sg31J6q1CHpG70C2rhbhoIk0OD4TGI9wCveJLqYv0GAA+MyuG
OMoIeb7/4PCdGnxg7GqqFGZlrYhwo8kLJTO6oUVaLplcJOwy2v8WBsnwYg4cac+DkXFwNIWZ4fKq
oAidm/MkKU109wKiQn2szbKcNO+Sok0mXykHrXWquocEbjsKR/VvMfVY7WEhLG4harBdnn0OC5B7
fjFh6ro2q7if2obfOND7xKi1A2JNlyZJ9s8wHhSs2Y+rvESBflPtSg6rH060E1AAfMWQhc4ZJQz2
ONebIg44igHFE+bEhv/QZ8beJ06T/ydvWg1i00rlGwer4hf1kPz4K1QJpMADiRXfADzO320UWDuI
nIvcse1lh9Kv07UrM3+ql+hBIl5jcoGguhnHl0NIQlOoVC11W0qLro+qOThsHnS+0gurEKJ6shvz
pjIaMBk4IITxnTMjwuN9GXLUAmJNEcHIq3Uke9VGDPO9XRARvMfj6duotIs5aj6KDSkGzlQMYhuM
A9hce4uwiCHq+bXFjbpV/HYtwqrWBnujzBYdklU9LaX9kB4vQcSdVS5o2zs4aEL8aMby7Tdzajle
f6p7Kd4WzQoMfI7zDjAEeI8dzz+Z77B8C3lS2w/gawTsFH4Mfs6bMx4u3+pFtr4dWhDE6HYdJHjK
XgrqN0q1mwzRfJUfqdzc5jvLaqOxfoeE14G/bsUGe1yPWs3MIcTaNmPyNY3Fa1PJmGe1fypEbXVF
S+LLKtXMHtYQN8XDiqwHg18CtIXHsP+silN7PCE9sPYZfOrv52djIO84IFmL28FdOcJaNn3lVZ+C
TSEpklGkz++KEKnLtxX9Xfrd7PyIiU5bP38sVLn5qbmDCQwSWqA9h9FiA/tAnAIfKPRuHI5bbeac
NOERDDGEpV9IgubmfbiIF2C3YF4TVURNDZoYSM/xmefcGtKmuWC0tWYM4b+STvEO3Bd1WKgnwmdz
/4ZVHsVil8AJ4Yc9AqnpxR7UR77MlYXbzc5xkEvsyhVVr/zWCMAhz2LR9LMWrOTn20vHI+P0elyv
nWa17B+/GQ7jlyQbQLUIn8HmiIGN4dKgVw9DRpXVVAfDF6jjwNks6si8boPc2ptudk8pKbdmHSYr
OOjqhumHxvvICJApxD9VBh+O/9rCkqtfNwiwGmLPj2WZUe8wEFy3NewZC8txypulGtjKOVHzfZo0
R/YCRVChHqTbCHYn9elvdHsJr8qESdWiOEb/zirLoRR6IcO7mh6zUcb4/rpRAWq8hG1yJjnZYe4L
CfAXiHGPzkCvCVvOkq803gdk4pnwmquhHQ59O7VLSp8ELpRi6RIf8U36KMFQYO4UBfRNBmyhfTA5
070iUoPpOiLjplgJ6sFzv38qONNO2nDbWT/yJLkhvFEaPl9B425xTS6R/eY+DM5IWGiQFKPW+aiB
iLeOZpioNN+DE388CyQU+hFIczYkb7mkVaMNW45PPKS/616oq1y5XjIIRW54DeYkRzEBvOOowxaX
v9XSXN0H+H3cpkXC8m0xBXf60inXwCzeLzboYrDZfwwH+uTK2qVAwZx/RnVuse0xIRHP6toGCBDd
i8mNTYZ+lWACRIfRaLmC3DFYXUQr4dPM66R2IP5IF8Xy6Lbn4iYvK8znhHKqa+5y7gmUmiJx9JPZ
Untx38C5KC0iGRWFHAUBuM+3fPxu1BzVFWjppYhGOIeO3UjfhjkfPhetRHIYvK8uWKeSLAbZf4qv
aiVd28CtycRNkESDiLdcgrUfvfdOFGOCO/EXQCNQy9LVe6VTOHr35vSyCwTUOswFYyV6bNCzREU5
nqdRO24350wdrIrTKOvDuep6cNqHXDc6J1lwjZAxCsPQq8AGqgG8AhHZlfDi0w6Wb+Dd4gGcWsiT
ZtYnkNo3Trnr+GYo/wtcBhB2x5m4L37vAbMsbOb7SNdxQv6cnjCk+yZT49Hbv1hpEHeAiyfdHMIs
UlwhTPOnN5Vn6vghpUWayx6CxnQV7WnJejSdimEb4t1JkOziwwt1hudMo0utTx37dYmXoUI7tCsJ
Waqa9nj0nmoDM1dYLhDOiMTlNAasTldC03PvoQSxaCpenORHp/nLmZbLJdwvaQJKWk2MqrTtooj2
CVtk+aAvQsVYZLmbqKUX0Jo19btHUKnHtxbtoZMF+gLXMDYZBZd8riqfSsIRVfaGTvQwxIQ6Obw1
J0IMTc+e9g/+EbIfS75yqET+qCxrVYuSS1W7T4/I9h2xJQ0kFo039StEm/+aodjRmO0mGLTVwSSc
hjTu1tIdBXacL5mM/wPpRee8zw2kZYFmx3g8uxM4eeMS3SsIfV87Qb4ImcgGwFlcejyRVeBxdf4V
cdDJtO8Fblj+QXVB6avLWwEp5IjibFBx4sVyYMOuXk/unsNi26qAt1plxZ1SQM4KVSqs+/0derZv
yPAA8dTJBMIQFQxd6faSqLdPW3BlbnD20e9dXVnpvTqXuZMS4TVjVdshumpVJUwvGd1hMthYP/Mz
d0EvgtZDbn8K4EqXzFndQTHFEUxwp4mcuvBwfmG5x4Zm1L8kuAdYxe760SW5ap9GplXn9dqqBtA9
WHU2PYeC0dN39wvo+yaduPiciODVUe4mOcQ+ZkRDcC549/TpPblekNirVtgruVoJhuwpO4C4bbU8
prPTpnHkWI1/o5bYeqFyHgI+8biAjGmOHbyYVp0C9GorL1T8/H7rOtBXAUSHmBpl61KWERczJHBa
zPfmtAvZKDZzwix4+vW3RhQfFyWK1ykbPYMnTDXXsAszCkbHPbf7XtfuziJPaKetKso+l+rMa9vf
htMx8fHO06V57UkvgZdsKoMZKIKKdMv8IMY4zM8LBP/cb4oXyV6g/8QM7vZAcKTxafq5vFsKC1Ej
61LHoLgg/BROSnAxlufeH1K4bIR60ZWRjZNE2CN+x+zeTSOFy8SrSra0BAKQdYTYMQ7Fr0QD70rT
AGDJwgvwCHoPLTSw+8zGyqbbTdIgM7mhThcpA8EgPDCVQNM9QgJ3mWpyoEgm+5EMd++9K+28vqoQ
t30DGD6+z1dWMiuawFI2XaFaWkMZd4/ljSM2eNTPB6Y25qH2WY782ybcXK+9ly6/W73kx95oUKaG
Yky3/9Sw6Rk7ihcMeJI6Flh4pKPwDMaG0EVee3OyiLuBEDEFyqzNu2Jgld+MaZNCuwexhTy/0PfZ
bZkGTNumJUGN/7QV5HBKRe/PmHHE/2LXSxyx4R5cFQUPqCvKzYavGvkIbz9fC70Jt7pcmHeZmiXd
0Fgu3WWfBA4WTbs7zxmRTb4AuvwB/UzkZ0QHnti6YGrCtf/Qitdvv8/rv/mE6fxj7WkgdflkXTRG
JVbV4DRgYt6ckfErm9TyBbBzoc4s1TrNDwNY4nvGUqbXr3xF2B+2WRET95c9HoZWVWXV8lXJWePr
gyKSDfSXNQMU9XEfqiXARhWQzCYoLf+MkAKNZbt0e6GbvPAJuZaNtnQ7tC9+ehuYOcCTZUT79KV6
VAJ0gTAYH2HMPliZ0T+7358Lg4IQAmS+R1ujyIpg7Y9hhjYEU7ZBi66lO3kzbzL7b9q40jEdS6io
yGhEUFAa+Znez94A83XMk8FqF+XVEIeytqC9ViXNWa2OWYbN6SvTHTZT3kRUVvFU2lThDmN8o+ff
3ksv4E/Rr9xomjdCNHdV5OY75oCPNsJ8PjkNFgTAKJLk3b0kjZwBTuYcZqpw4cGZo9Jwbyj0l3FP
0T+GNwSEPB+OHMVt5ki8L3WXJdqDa2ZDar6yKwTVBzZ6C0/V+sWkLz+/biuFOEJ6YDrQOmXHve1E
6YmbLUQ/3fmNlnz7Vzyeu529Ez3TsL50f4znMEcK6kYkGZvFnJQQxoD1t1clnKBkNJki/aPvzd9Q
qSKGKOfC57AWtlSKn/lDAMw7kuGY5tWpa3d+Z/U2knJvSDsXYKTQSQMLYc1Ox25E6k7qxfGeXlQt
u2Q0+exED3gxmWAfPTrG7sa9kJmUt46AVpKr12Uj4bngAoZBiMD9jPLN0J1q3QFiiFerPyf0c/L3
ehCSWPEN3jzEnCu1NV4KgjXpmNDOuHUvXiGsmuAVlcbCi7DV+0uBGvekHyZW/ltYuFtVw82RG5Tt
J9Yja/roicOcP+bTBiqvQ7+C9STBLiA+iA78MpNf/8YYwmNH3cT618ymQgJjZ6qxTtDwUeBBF9JD
jr6J0kLiouSdKSDsN5zAeD7UcDt1NOLRbZ6WMtMO2/t9VGie3ngxvHKYLGRlQyNMcLxMgrJApNVa
KEMsDQ4Ct2KABNiDRvKGXqf77JLF3qgMabJiiGOBcPGbBF6pKyjKtOnVvMXSG8KvMSHQz92NKeoC
xuL57+GAm+uElkuB+JN5P4eE3POctIZktm5DlU52lTVFkOZpAI4hWopQrmIfiDwHiwxFVth8xRm7
7egC9yYa7RHGf+55rrk1t99H/lFVHSrxaG4X/qP6pdri9EsTcEA2gXet4qnNeYqirZ7rhatBeler
wBWyD+03J7wCnsts3lJx4H5NlD6tYUL38u80k1ETA9RzaHtDdMp61o22hNuBBIVblLq2MEUucnVt
80ONCRaRcz/ygedrHoVgWK1gKjqabFqiv5Y5W4/mCR0fsJ3jZSnIxpAhAd26RcjNUSXUlzTXv8VE
f6l3C87M9PXWKg9PYCfPF01HLhIEC+LLehnSFfXtfySlUJ2f7QOS4tPI3ap1r5IbYvGNSpFR1a92
O0X3+kOtRmx4luKZvUVFp9cQKg8kF66h5aBfNoroyEYR+GFGh6M9kvq9h34AYREfQztjQKZ5qB0c
d3xgjwYn7WiHlZl42ljOFsZV9ekYM70Z1KdA5YEDHLmZZP5YFUQiVyHSmXzKPX7/ZWssx11Ty1Us
sLSj8zNw+5vBiVPTkKbVLh6aVvhCf+ne4muI/FMX7FWU5bo4ilsCMrlpZitQlAgKRJUOKv34g0Uu
Lr1Du0z6PsTwKsagB2+Bl+IajIgjg0ZQ4IMOIcOQR/xs8DN/gpzsNugtqYhEFKcYuFhYC20Tpmy8
INUSwAGyuLHRYfd8DFmzypWca/895RddkdG/cuJ+Emw2WpdRMCg+7MtcaVHH1t6SVGv/2QahIk4I
huk6KyyghfKnizel6ZyEJzV8EMQPji7Laj2IrR+0nOZdBL8MPAW1DYUncW1lVsnYGfwZO2dQ9NKc
6wEXuWtuyIi/+zx3ZNV5gSl8nUI2f2UP7lCfnQ5RPdThrGYT1XGA8c1Lw6lLRS/oTxeXvz/ZukWO
/gJTNijQsrb6oSrUu/KB3mULxn3VCIDTneG5aPFEFTMUC0NutIvKMdyJF10OJ1S28R43t5vcrkq0
GcAzS5vt4qobVF3vt27JJwSgI3mUNnU408cze2npqQoIZpUdWGA2xvwA06CqlyI8IS05LtTOKGZZ
CiqXVg0BytRc7aogO4twr7CLTc3k5IPYOrfZwQogVLR0tUUh2+fYueITAPfwHey8PDkQBz4XVdYs
ahYn9N6KlLWlRorXHZ0bqgfvXdvWbUc1a/f8GX7qPN/3bs4zOSYvXYiHzci/PH1jVdzGdeHDX1l1
Hoz6y9GDkk9te2b2FOFh7poAkX/bzHT1kGhI0vGvWmQ8ffN5IYNPyfzcmY5p96ah2yIgaG7sJW9T
dJ87NHkPH35TSkHwfkP0sANoifNcDoPlOPP8ieuIJjrBJK66HmMnrDgqYhpY4RJDVAYIXi79z+HG
mn3lePx2K3iupMWOMV2xJXC5ASWk2hsODcXdGiONw0eCwDy0l9feTyEXfIVFNcvqYqFptUiNl68m
1xzpclJlzZAuntZSYacs0BMYj6R5XKof3zprSgnwDjc8+nBev+N9NmxGIeMfDzfsWs9CkLbC8vRy
ctGi44J+p85DsBGYRJNmELNKCgyBs5uOkZLbszQVAGZzvADhe01mPRMfiduwmkpupYvY5n31hh/j
lkHXWm0li8aXxPqP4csrmqgN+UWtxDSV/66nrZbhVNkcHMtaxoyFYCEmjGTCsopP37Wn9VlNJ7HN
Z13JJZ14ioWBJtitPumlSZ5uTJQk18uXvEmm3B+t8AfAeZnFj/kBtIN5rLgxtIaim6kQs3/8IB3B
um8HKNiI9uqXBo75BeVJDGfJ9a4jOUeh7P4c+XnnSXVNu0kkWzITEFzMxEX7bPVtG5n6jyJWFAjN
XbAITlJt3AaCj2+wGwLNFWJwK5gfCg3L7EXT+Lc736jSDmkxtcpg9g3AScVaDgsv6jqmi5Ev1njw
8g1kNguXc1KxWtEQh4VPde23rjal6rIS2EEctt7kxopfjI/tTCupD182rPISHwAxm3rjoE7cJaKp
m/NoYJUhHq09t+cXMgF9w1N4yMPpyb0BTS7s3NsKLUT6PaAUOyPYINhSuedER2Q9p76qGaTR86g6
a2x9Xb5AKcCUBxT4zzCp+PYxsxLeK4RXN4d9hq7Avv1PGfXp1WYXOTLFjQbtX5XQaR8aMOXg7D+Q
X4zWtCl1zaJN56N9+piqeaQo+w2UVg4JYjnhxU+LAZBM8U2mag3+N5YdTW+2E3kr1JSz8LYJdol8
vnBXsmtUBxhZyZhag8AJlhY3CcuNlMqXKWCO03SHbM93SqEXKEvLnf3UMFzUkOoU0bCPazQrCWTI
YdT0r6hYtBPeZ8VdJX880FVfAYNKzszy6rdXpBL2L64E+fbLYxxD9FfSImWsTbvmaRTJuHRqyDbI
j1mn8gVlwGC3+Sz15I0Kgst71zAFYPCSfpDKWm48Sx/DEydCd7t8VJBYTxNjOpyMz1DzdriPUN7f
+jQSPmzkNvRHt2kuqJaIV/2vwdZOgdOxD0VbntPidhFlfWWIdb1r3wZd7xGD5u/I9VkrP4pQsZ21
CAA+lTf1pjKcb2a/WaVRARqPywkd7NFtiE4SkWxMTbdn5ZCHvRFSXtBYVAQ637bAQPuHPG59oeKO
1FPpNgbcf5vzSLjDT8tpO4+WMz4vgBC953gkV1oEi3WfOErWfWkcT0agzkCLicw2f5si9Rozha75
ihtu6CnTSbWzEazrjqvtDIBC40SPbmHQbClYXhsbCshfbYLyDj5GeVzE1h8bB1Jiv6MatEhqxGz2
Rgr9Bkb5ZiL6AKQjiZcI3C5RmsbVuDdty6a3A7R1K9K46Mbpi3trkH2yowMkzFdmru9kNOh9wXUJ
P8ETgTSacTMRRT35lM2waVs3yCSkDq2uIT8V96/W5oEy7c+dNztvkSZB2KYlMDgVT/PzAH0/Qpwq
K0hWDl5MhYcqo8atLmUqK1w1wzB8b67PeGZ9+3MAVNrMrwjbtV511gaiSt1QW/65U4PF4LpXDAaD
5UUU9leRioUgU4UrFyEU+KkZNIU2j3Ri0xyqo6wBeiDOnpb+KgeiM29VTr45C3rz3F5nyNyPBjvj
cAJJp2KRPSGzdzRNrV/Otms7FRm20BgeckDgdaXSSAK9z716Ib4g+CsUrpYo8T6nLeDaumQJ0m+o
JE3zXE7udycaWrcbqd0Y6/LjvlKQm8QNENgyEOL4YUVBVV0THrfOLwDcGf2YsRcC9f/PemLZbP0y
3VK1eX0HzruQjtR5KkIulyQXpOF/wrLGXL74ACbXR92soMLqrJ/6LJ6uXYc7bBz4opUKPCHBeuVD
g2NO5pDTLwttvBIEN0JZc3lt9XktcD6mScBcQI2RgImkGgBrnHy3O0itPClDfRY/Gefst75Iq71I
107DBA/2fSE2c9PBxUkzs3pLeQdkh03W7drZaKzW4xg5guDwiQ9C1hw2H2IwEyA0DbNiZYos/v5p
6EoSzfTNb4YrXFWtBiuXfsZBLtGyDLCcMiNQDfzdn9Hm3w10fzN2LrVm1ChQMWSXJex0R7yRUglu
XKb44lvRc08bzB62XxWMrh+H9owZBibZtfuw+TC3S7pVQEYIo/MOnugVz4jIWyOqtJoQ5aoplDV6
mW2tbIJnsWrYYbQ12v1rLTrhpa8NWHsTYH9/d5LiPTk0MupwnYor+DGn0dxIl3Y/DJbrRpnEspKf
kPUMRXXjWzSThOL3bVA6dZ5yig4VariwNokhAYHAp/TxXRzrMOB08zqkwI1kL+pCpkYsYrXJtotX
oGMzV81AtRx1RGJHbxfQQFM2vag+/p4m0Z8PsNh9WfBeJt57jal5uQXMvTc23+O4swlXSwCbh3/B
XepldHD6sbYQvXXqTXEFQsRUp+I0cH8+1VQaZyCj23Aghhok9she9zjKRQwVfcFCq3Y9jTfG6kLz
gPxu0KX9K5u3HQG06Qm18YZj8oDViNCB1oXScHQTIQwvwhUa0Z64PSjPV4nKc0ux3d54c7mbwMt/
oP7cW+Ad1TQpMIdBpJXfPyXpBZO6nOM50ZtDtjL7+k9yw6GK8R29H02qud1ReOS6mglIXjpDmYGu
afS4Nkx9uBoMMERLOdQzzzLhyokqMWQbwHjd32Z4yWMV1R2mFCq/rVw0lhQ7mFSHeLJ8fNxiyt9T
7cVTiUcT3n7SZbQdfXXo9ByCLMlOWaL81V/nXt0fsfMordQqUUCjP86K2TDpSxliGPEdgL2eae2c
n1sikD03Ah7c7EUfua/wwr3wYMK4zHHG53XTpzYAotgq7D7hdj4pKcjyLAHidadOWmfg3ytcXb5U
d4YdU3fDA19LrpopPsqcjwKCf0bt1vi99m4+5pa8WrvCLzAFFiecn3SdcbF6uTZdNpJ5ZAh6EojP
Kbx0wwR5Ybu7GJD2foJlnJDPI8IgJQXVJ1gdrR5jtDEBNhQUnmlQLLdTTpijdix/wlkF+M023QPJ
4rE+QLZuJsuat3TMVO6ADWezMpKZ5HSlS4sJSan/rxYu5YWjjPj9zQsTSC5F+U//MqUmXULrXBBt
G6h4Lz+Lz2QEscNPaPd0j7z7u14qygMatNi072zUbxvuchFco0ld0CElnTrPvr7c8PDiLlCrEuvc
KR5NEObbnhh6eYOwr6A21Ro94KkXC/LpBIBuSA8X4RUTqWDNGRClh92kEX436IfGs3N3rhZeNBC7
qys/rBgetX18CN2d7bDr+IgyIqkIqkV4ZJf4VqYCLAYxVsajed4IiA+otL01EdahxYLVQS2anySv
9AlQx9nAOnDl328NA9ItHuQ8fEO5+CHePLNnWmEN77IaexvZuXRD9/7bLOD/wzuKkOWHRPe7ng7J
e0MbKpfjtRx6ZG4tlglgpEVrhgW4cWi0ff2MNYRcANPS2HxbSLBfqKc0ErjgPIH6C5Hvhc2XsiSz
CVBOlQDc2QQpQamTKM8gQP9oUC1zLClDwZQv8mlJGV5is/HpO7fy8msKbGNapBMDufnT86Zlrzjx
0f5qeA1YfJOAEz8a2PJBlR0kDzhhExFxENdlANfTi49dTr322WJop14Br+YNs7gYxrHPbYOI1saU
4kEkVmQjmIqCF+P5wK1SRR0nK4gGvjDeQagYinNZ7Q7RjLAQQN/bNGiXql6mLzecs4KxVI94M8C5
ifpZ6N8GcH92ttqy6blkOJRf2zS0v65lR/oYgCalhQ1+iZfqDzfkWpm6R1rHx++kdWQeeUyRGWbA
IZ4yfq8VIoiFS25MqD9lGsqAf4mDLvbLATQBFN+BanOkk6hH2cJWzYQvra2R7X1yzANYhqGNCisp
fbrzxf7RqP+1956dZvmU07/Fei8xVYnQ28fN6TOwOqxsBxM2qhEpqI+BNlHv0y6K7fmZx3S+4C/V
4uNbZhSqAFstvuPRKoRFueOW4neZ14Kqc6L25v6mUZ4Y+AkwTun6kyz5JBFv3PcRx5m5+83MbPRu
HSpJVbuohXwatQ0D2PMwsr8ye0kRN1pQnaoz0BMqxcCYuLryke7jmH4l0WshHPNSvOZKrKBDWM4p
DD4ad4PL5uzok2rpYwbfZ66vcKrzBqTTFKO4joEZ4e8SPiYNqgOl+XToGW/HKEhX4CgED3aLADON
SYGdzF5YPxbHtbiw8eQQvSjL30x4TUivKgt5GRBiFmsIvEakbw3S67k4lUy+Z6iy0jMbFioMny3F
eALarXecLOn1MElPqnxcYCDqokUdb+p7ApVH8V1MZqJCPnsYZI/i1MFlaL7lzZMWbSX71yOHDiL2
pabz4CuTANx2cjvZhX04QX1odKvim5FKQsMKYS+G7r2tCWepQXwWYMqcJn4sHsN7D+Jpn2/UgjGz
qU4cwxh63vWFDdlZIe+gUvPeRxmbl9A54tcSWT4L1sqbIo6yyb9Geu/P0BFgECEEwo9fcEMkzGY7
jCkFTHqx05F6MNWk91ssd5UI+WRAzF6MBg+mRBn07m2DMsYuKj6HLUsCjWICcdkt4GhuxfwxJN0c
MvJvaA1tW0cTkPWRq84HFnnQCJ9ZwW+lhcAj2ESpe8r+hhwBJRa93F2rYputGjWNsCrp+1shKB6u
x/yshzzf53mwfqXaChrlGFj9cwcyVDwbNs/7CXuDks4ORx0RVAGJtJ4QN3s0Yt14VMNBIUJ/6Olp
mGpHRE8dnpkZ0axWsj5sNDGcEMxj1d1QVdQ3VfAI/yDhBR4lJTRjWYxhw3dWicPg7wcWZCqNK+IH
1Ag/LNBoPtzANoCejyz01gOv4MjXyaq09yt//UYMOEYIjQb76GBqUgqI2c4364tPWl8KINu8i0AF
IY3vPud4Hw1AQFfafvBymTJaVXtT+EzmokxIUqXIMi3keEgXbU4XTWjUktCD5pXYhLa0/nSl6gg8
7UFEZ5QTWtVUOetE+PaH459ctI5t/huUeerULaTUSnHGfyfRPDFgJ2e0SChRWIYrGIpJJ9TLY8D3
DdH0zpoiADbZjes+2ByrSz9kuOGSokcaCTXZTGs3QXffVmVMITbhfVtUZiQ8Lx4Vr2JS0sBWLZUr
ALBNZS99ekVpYkE4tobqG97M8ptp/nibdnEAiu7v1mWA3Tcpx2GDhGM0yuM+mGyooRHL8hlXlv8i
1eu5QB+s5lkXBiRUUbmn5a/85eopEmiHw/shP5cVmwiCXGZtcctJKIs42Pnvo83JSaZYDJe3YOZn
rCL7lIYtPKHSnyL4D47PtGwPtmEJIQzkn9MZlmg++vIgrjsyY6X2iyup7HQ6KoKOKJgaSAfHhYzi
JM4MrSZALeCnOt91LFMBzDy45uLFOw72SELkOXY0Yvc/dz/dgiVyqXG/ILDRHb7bFExLzcrn6hBh
kl+MhxsGgNxPdxoTU8zdKhS3c/+dTsOxw4mZHY8tIcTCu5K9Sab1/euAiJrrsyPf+dVKxNHrmg4i
3CIsfnbxcPihxOsrO1Pe89ggwYjsqLgfxvGLoYbYCRlK4dYYHbAib476aHY8ip+tq0pAnPUai7Sp
S1XFT2UPK60OZk1SEYrXxg85YlLJUo/bmVdXmmhPxrl2pDUfXo24rZIa/xiJtnhTbrxdXUX5K4i+
j09jx9kdTwTjukg8SlWc1/gOBBXWOXqavDz7sKjm7Toi0LbQV5rWHAEviBMMFC7JyH/js6evVoPS
VPQJBu5UPurkMWpgIwTdH9An4gY5BT/eOY8+f1ZMWS9tXywdUtFdfrT+RHmx0xCyrn0wfdCkGgxO
nAspG9O/qhIiDdOHB69UD119NKdAQuVBd9DUFyvHXw1mJ7Xo9qBtQvqzHvdDb8Sh//h4an0yv5j8
LjK7LV9We48hxAPPFS9mg14hvVIyXR9OKj9Ll9isSwRn0ZtvHPw5WZ6grTMpuKOM+GtA36LlPZlJ
qJjtsNz2WHZ4GdRPUTxAnbD6on6AfmRzMPnk0xGAq57xdehF+pjxRF4kRNuBZ2BQNmdv3zZKUQL4
iuchoFG5/KZftZJqc22aH5Lv0Gb6WPjFHEwczMJ2iiZXInHPpuH+0wM78WdXCuIJJGRzDCjjtkfq
v4D68HNm8WqoHelRab1akNfVsM+51SDRDf2MGzXMvtalmm6E04ss08Gr5swAFIi/ptdY4T4lT4Oc
PHiAZDdSNqCmoaavUED/mTrfxTUkornAEhgJg/tJk8w9MjB9+HIUkv6Og8IZehr2qIG222K7NxUq
iB7gg7yQA8wLefDx8+OuXv5b1MTG9ocNYE7PWuyviMkgJQ05Q4ch/e62QYKx65VpuuJWDQ/MpX5k
6M7aMzUMS/uFSZ81PJIdBvm7W8PhJ4GgUU3jttAyWjd0q4M0Txbw7gU0mTMr+xhR1pkcICauyimj
ukFzT3GqtYtfIJJnDqdSRSHxoIaJ2VvC4Bh+TgKHvrzVpVbeGtMW/sE9Ao4DpOIU0uMIKR4uuTqO
37tTyl+UsSbZGVP6LLgHutPUkYjMuePslmO8MJWKkRCmFqM87E/HHcHIRHtLpy3sJr0yDwjK0s4f
KOygTz7VW7Igf/pOuV57tHRA3bP1Yz1H2PZVtarfUJ9GyXQYsaO3rIO2Py6aPTQpK7vcT8SwIAJy
/HhQ4TYx1kj1847glt3hJ8ZjMLcblejtVct8I9QrITh225HGkZ0m4LKEeBhecZPJWvcdgMPonFH1
5iTodxtXEPPtr5rQucJSwcySW2Y5pbQdKbJtnY7vYxdjRJbYd1KyRbYIL/kQ+POqfJtmRMecFS/g
njsjkx/BCcFA1Tgs8DsYn9S0llH+7tdZiRWX4QzONUBP2RxFbqrkLUblzS7FPC0/Ww5SsQVzPlgd
/t3eH7oHhXLJQHvW5aLIpSR4Ck5fXl5yMKobzoqX7deRqsQeJZECNIzEZhkPjxVyN33w2Y3oqKR0
HY6+TOooRDBLSgIMWMOs1YAmOKmOc3jwCr2jsEl/4/1r6zClYjq98PbC9SuxM3rGjzvhphqCrkn+
hDrth7kSJgQ1Lhc8PSHvqb89WpJwVSh7LyQmQSPFxjDzgVQPyZ42xavekDrLu9vTCZENdwR+GtPK
UM6DQdK+a7qKYx+szKB1Uqx1wBMlXXrE5djBVvmc7K6naZVxYhQlhFM90bjzlBNR0nfmYaeFUHKF
d87Oh9VJS/cFlkQXJYJhA7o2ssYv13C9AJ8lVF2ZHxkGObd7Fu2VA5TZ7+VGmVw5E2hQIFWmcHrk
6uOsCstM2y27hpAD3pCsd6LgySLLll0Vmp12uUwzObr227pLbJQse4nmD5BWvMAekEpBTpaSuoF+
dLrWPftYddFLY4D82RgEhfgoHudgMf41Vki/JvR4Wq7ZhZjbsnZkOviKkS6RUteoWaWpEVvhxLzk
5joZ6UJCKkEKC/Oyn1SESxtIP859l8JfKfVy0ZLBOk5nSnBtV6YBmMzwa6wHTjaUo2TkPS+ClsI1
1qbu/J25W9bSFsPYawTo6g+4ChK8YfV9XDrZzOn8tP5VXTNSWWVYBr6lyfEH3a7eHzGhwt8vkJts
okiFFAz6VAqfKYkpN+ii2ZTGUgQHDMYwK4KEOwbnk3U6NcDykiNRj0/RvyKG86WetsWWfXCKtoWf
lr/yJbvt8xEWaa5NbKoOk4hioHOJuJT/UTdzH4y6ukzzCpJbNBouoeFmqZCav8ge0YU9w0c8USsb
xFkcHi/2651SUvArlapTBRtWZ65lUM7LPS+qi8aKJ+T//dVJDaJh0RzsDPpo36mNDBhtLtz9HjVA
1XREWF1xMvkIhRqbVGDZRCTrrKTqCm/OAkbe9RGh4hx5MIr41y4GthFtAorz9E+8Q+/VBYsp0ou3
8ZQ/BBAv246eIXysSONsAOCEaXkf3eXpmQR5LM3xJ1Uu0BOhEqAOkE/HwDDfdIAO4LkALcdSuEHZ
aXZkBnj+UDLYWzY++rmI6EXY7vZ+d1q6mK0K0d4dsYNy/6FR1ArYtUkwFbwEQpiynh0iXyDDmIyd
6LPzoCdcz1QIprnC1EkZ4XA3l8idJdn3/GMUrpA3ZQmfwV46aTV4VC5uTpx78AbGYjG06DJuGJwx
5PDW40mfnBLWZEt0vpi8WT0kvIAQVYSc2V/+X46uRP+5GlS4EJ0BRd1ISxSCtN84F4RPc/pa1V7z
cEdlEfrFywQ9xIALmH7cdZPUUHL9NVe248c1gqL+kOPlDDqpZoYvyBom4T4mfOjHj9RFsDn/tbEC
nT/HnbTRWm2AiJMBd1ygnl79u6BWzKVBdYYmpPu7WtklnQ/SU3DFLNzfuXBSeSPlOtRX/SMJ9x3G
JpIqin+fB1tNyRrwOd3bdnvwyBTwS2+1uIwh3CJP0kT6q/bi08QqBHPs6/t6i3XnlGh+XrvO/Q8X
uAeOWGTnRqjK3HIk89JqyEUQpnvQvITrytvEcVgHylTyzbpCLsdWlBOAQdgOEJoevI0Q03qZWTIq
S6iNToZK5zmwwzqI2NhGTRtYKdjhjz8CO+YJkNnmfcY7hUdtQWODf92Ug1KrQdDId03c8f2LqgYA
9erwPxHgQwI/JkzM7WMFOUXIzPtX2yAvRUGAPVKbzQ2SkxEFcWdOQvYdzTnCod6FJEp2aS4vgUd0
6iAdNMxmF4x5hyqH7t0hYVsNUNKyGf6kMGbIInEVFI+2YV087UyEiwXrVs+H1/EbXysN2miw+EYG
aSwNJ3/h8Vlm/UcDj+txGaqm1oGA76q0gRBXGu7VFAPlvnOEU+xxaY2q8pkYV0jcgSoYLOPJd68J
BUQqknoSETRlc0HCZSTNQiYZNnSnalhrsFOGvtE0+wm2jDldaGG19UvXDCwHMZdnkUq949nYLHE8
Me1dOcBmkGHtvX+o0Fbuf3KPX1c2fbylBOUnWCbjhCKuLk/yiiuon/SJeprsvbgHOl1Q/zVvCKGn
++mDc9taFBQ+txILAscxC746gIy/pbrjmltc7XcAvi93qPbl8H2jtb/TAsnrSItHnGprv74BJ1Jt
1U7KsHphVHoyPu2oFKfZ+ufRCVCXQ1BHYbau4Rr/o0muFVa3P+RsHHNefhtoXFBbAUhhjgx+vMec
kT6Y514qzN3W7lw5QrKPXcOC700jNPOvmhwZaO+VgRcqMKKBq84rq2UUcvxEDYnS3/4bdyqd8gZ1
nODiTf3Az+RQ0o+W6Ba2gBbenmwaJQWD3g9iSER+0xZufMjs/3H3D0bwkrjyflhQwYXHtpmaPRO/
KJNKOyq24BleyJrHGn0EAWGYH2iZOeeAE6HP6OHmHp4PBeYW0XQoPROqk7OfrKXNTBPiBTa11MHy
bDgHF3S8UhZP+v5cu4karWOYDqt/C1P9tb+LyS1sqBrXfiN5F2CkrTWqZP7lhQrtqKC1jT2PfDc7
z0Lon3Q58CtJNG4OWuatE8l3HOY7eBxMF76TSrtXZwYvIhvrbK9IuN2ZCbvtd+Q00vedFQXm7T5c
Ng88dBGW1kT9ygKSnlYqJ4Uv7lwFkr1QbrCPbCIer31oyVeZcE58KanzKIMHrXrjl7StKNzlCXc3
H8SbtiNAhK8hQmPraHTR0SR+j62gRE/yvsIJvltuTQnLTqZ4OAiCJYtvsnXZ3Zg+nxJmbvxDYKSO
AbwxOjM8vZ26eLkWctF5ZH3mMu1uqQqAD2sQ49ESOMVqY6psdSJyly+lpOTuppR/ZVrROUnqZxap
S1CNHSMODMsTdAu95axu2yuNbo8TnZ0/v66VJRRjwnNWp8K3+cY0fMsNaGc+zmA0C7P0HfUxVLvB
K04GmdzEVv/2i8mXtnEUVXaOblhoGVM6Qm0HgWL8gwLrtnTwJUBvJeTJLSPQ6Gw3JXXGMMhsrQAK
40M6FX5bOq5rkNnwAAJRL2rKFeN+ex8lhR5c9pt/3QJPLOqFyOP0SLOehVjef23szL1X4j70AWyr
sGH9ak0kIi1BScDDLngrNCFa3QIiSdSr9zWsT41fT0ox+iQ+R2054nbtpFs0sggGUJci6kIegt82
BvRyvx5A9saAaTG6lv4Mn2rinaVOnJnWtp7be4zhH8THXqgmnMkb0ttqqWQFL9BN3biZe63EMrwa
54Wtxdq/nAMF+gisTwxf6Cr35GKxAJwj4cKufqyp5munou4Q2htLbesANmoruJGQetwBRkf8IV4c
eqAy2XIMzy06r15R89ksE7oxYBOoTVBCkrYhM6lImGiKwYF5N5e8v4ZIssOqHpTcVtSLioqQP0It
zD4XEL8ePQoJVI79pbfjMyf20cfHPhVrBvXh6s8ggwmH+zUT9/mYZVkD6o9VBWnS0TgeXrlL+ENr
uVA/8fsXlvAD3KgbD4tz6ezr4inwamr1rxGordxZG6En/teSfS7qR7IxkKgU/PSJwDhcF/KC/5Q/
r9diZm1WyG482hVUu81Ki4CxR+WB5lZsbejtKR0yqeoafJvnaCjOhsxh6e+yq3liYAXN5sHA3Tcu
eKT/zcSQMRn7yBl9jErZ1yEP5M9rpKs8WIVA/buFpScVN5unQbKZysULjf4wl8H8nVsRgz9WhlhQ
N1qhYWWl1Evhg6V/GFsrI60fFs9StW8u9XVUFnSAVT6SRNIvx7cvNxEtn8/KYRPNEjBwghPH70Ko
IdPeAF72e9ipg58d42tiZIZyy9KeMIV2vzKQi/tdkDQUz+AucxtMUk7SJX/X211tbS7Dd4fyRC1C
fUz4NbTR2TH1zDNID0u//sMYS5zy31lpP9M6btxusVziZAYHXLw/E2UQMpdvYQSEuZQGGA3dAOo+
ixqBMk0xajYdUpzroLyyITkoXKwYOAOwIEJliQ/mqxeKqLxp6/3xCWNeD2B1lWJNHEhu6DQVB/Fl
OXFiED8bhxuPmoRyRUmEo16+E53gRdwqUKoRUe2oCuP81v7PK/H24ChuQbHFlUwKfgYksqZur/gR
Y3ojw8F+znw1sI6coRJ/zkDNUdOglvxXmbFsj87nLaGqc7x7klejnOce8j3+6jCL5M+sagjKbwg/
B4+sh+FtYJ042fc5n9XbQZPGvlzZk/x3KcA22phY5MmUPoaFE5398Vk2V16270DGn9tm1ERZ1Koj
PDetu0CUzdeFVgOr27sdJ6f9MkvMBhbsI7/LVavmQwrfh4uaiR0Ox/Izavz1yOi7o5Msg6Kzwcdq
tIoAUv7dLLwPCSqM594h7EZD4Gzs9gEK6BPdaLgrC8mByC0x536Y9n0m7eMx5/iiCrGMgveOXnt7
xF0cFgdA/VVaiVdQ3bEIfUWdMcKYHSfJeK96YYwyv3EQwcckLpNrpSJiqXPU9VSajNHEQkMLKvMU
KBkXoFq3ZnWSuKG6NFqNQdV0vzWB/7WBTYgbvmJTv2iG4J0Flx+3TNV3u6t1Z0aVQGqI7GJUSZpU
oIMXZOfpnUoYu3R8oPLigJ1EnpqLTcZY4feDjc1WWIMEjJ7vwlYb6i9R+ctuTxO7bSS/U/oxtKog
GQsClyD2uAk+FcYu2RkO0q9thQpOA40qbMG2o9x+dxuNUZRd56DIqhFCcP380/q4LeVX26aspEF3
EL0BDLRK8kvcDyOclXc1oENBeALcmvQwFaqusXn14SKZD+1rJ58CT8wYiwq70GgpfGe7C8cPmC6R
rTFuFn2be+EevLdBK45eVSh8NzrXH7rb2XXv0gPxRkPhxCC0jsmxT7yFLW5vgtYNnMu0YczX48RZ
2VYx+R8pJkAapnl0NHZ7ys+sGNNvKw0s3WTOXGaYhrH7nZlcTAkVMujqsVGUXLQOArIdPfd/B/8S
Vur4BkavpJctgDtAlptJhf1HVWBIFa0VQtHkXp9mA6uMN4VJIgRZdaJkiHqPIIdZ5ii6AzCXmOVx
7EXXNKbtI2uzVjUaVRsyDNtaLMO/j1wpUaoMVPh+q0HZuRClkdWYZAEPIvbiBAYELUwmGBs6NwK7
vZi0Vvi37/JHRaHiUoiq+RFTW0OAbb0bvXDCqV2nNoCK6ZNIlUIRA77zNqmlTA67iOaOzWe/OcDd
WfJ6JJugAZDVDdeXK7a7MKuXHWsJ53k1CsEYj0HE1COp1z/+DdalHpCvmkA/Tug0auJQIza7E2fP
TOaMMYrV1JM2MmOYj51Wef/sCemsX42MGG5EpxBRa31Ko3Qy3omrO3nakN+i+mr3HhQVcpO8y517
oaijUrvVojwrG3ZpEwi6dQ0leXdSTQ1vvy7MyjnbTYD0ZGNhZ5rvLMpZVUSjrxjHJAveaLOleXe6
U0KBmaf9fg85Uc91tje03wOAHbhpBi0eK2PGnde4S5oPUREoNbyeJAgiVGg0ORiL/h+iEOsFdSmc
HYGrbBX+MCyJlWiWqwa2QAgT286FhUbyoLhT3bXToaj1p604qcYoagLfN8NVjhcbwepd7JHmQRu9
ioH9YpxqP7VQizWDyG5OQY+GYHcYdqUjN67X5c+AQk4iylGlNu76OpTBzyH73w3+grfmnmRlVe+s
njTChlWPx2r5iHqnTv3CX7NmvPiFs5aEnvTES+B4ubw+muOhAcUrf4yyde106pU6uv8xyrghmk6H
lorIrHeq3PtHtl3lvxUfm+2dVwdK8Ib1zkbe9FWrLAvadKCDBx71gDND4h6ISXSzTaqsdHKzv1kU
9WD+B1X3eZo4kyr7DUFsuZcGPKuPDGZVEeqe48JUF/LWSQucCVL7uGIsfyuI3ro7dREQPLr3TtSM
2V+8UypH8ROjkk7NeDhLTkwOJepHZXK5cCQNePBxUy/G4xvoHjkNf1p6hAKkmLjApwy3AHhL2M9O
R+E0vCCMeDm55n35HadkHA9dvtTQTLRmRqhw6wlXF+lxyNvzEhz3Wcb5tpD9rKmRuLansNNAA1hd
UL75S+dyIq+qXIsHTy5nMHMs4Cw01UZca565Q/RqEH35eNQOySwwIIw6/EK94z4cEUoYMKOmZVLR
7P44BtXK1vDV+a1A5cYlDWaJJehPZRp4X0LyDsIs3OcB0l8O9DT2qSrkHw65WMkgKQdT9V7tLQEp
EzFP5KgcAkJLYQFXl/V4VVDJG67hOhLJb14nuCuEwEjQMS6Z3O5aBsGMYs3HREnr1oAj8adqClUW
FFdSdZRj++EEWb2eU0Bwgda5Js6TW3JvFnAaNCZ5EiEzV4tG6oexmitzsltvGO2QKUgHpv0xgboD
TF9KjXQRLxA/38qh/cTbAmxyHPSlXHCFY7srDG3VHgI7i1gCWcc2rqjD2YaRCCFrLPu08rTUMC7z
3pfAiZy9n3D/zCJG5a5HqrBbrUnGhniBvaZaRDbFw0joaXpr98vdTmVZtNS3ygFPOc0LD3Xf7SRl
Z5n8wsOwoPRS71v/BH/+9H3KZ17xPYvw3+Ilti8FUhVNLA2RpNWco9eo26+/UGGrxnxWHkG0mfiO
XZZM+khZEWUsC+vNbL9DgXtv34qid+ATwH7S7eYMd15NsoSqmk6qNugrFTlseSMzNPZBMGoVI5tT
JLyj2UWwgtHmou13sxwSRzhUIG7P35tUTHDDpsSApuN5fpG4D/tf/XSQGckRPKwMEr/Xo1HqaOjp
4phARTDnPH+0PNVJVXEynfzKvQUGpluSotOuIfZLAdDZvh7tn9MA1nKG27tVbEzY3pa0Ef0eaE7R
GI4Kno5Hvr7S+s2XfyOe9b6AR5n8HGlyetCtTKuq4klmtSH2mxyoiou4J7bT/3KqwZjiQyQ/FSBa
NdKYSG15g9+nVXOrc6fzHJLtaKpMexo9Oijmln5yJU2xyYjmSSN2q4891HE2W9ljSHGwKuru9AiW
/EOmzGLUnD9k8QXSDY5AxFzhKU4y1DMmXvHbWtcyS6XddpI/T9l0fuJwI6ixPoCpvYVubCrI69uc
1JcLZEzXuNHhODMio+IjoBeVa35yc79CO2411tivSTrfZLVGrrJb6r4vzpxU3COkDxnlDmEyUbh8
28RgPw1VqvdzDpwezsYt3AKzw/GH5BpRhUGLiT9ntGlURfoiswCQ3IjpWOV6zXpa/Rz2OmuLDaec
XkkYwo9sMJOnuEuRz7ttXH//Rt8/5QSew4KgR8hWGGsB04VFu99wItjCRRnf0x3hTaYzijIB7UMi
YbzvkAYlgJAdkw8NMgYpoMlFca3ggJdEfstlRoa46OWdf5pI/Ca0KV2fjxVHrlPwmNXt95/AKDsN
Je7VqBN5XRfPV9B9NdbvdYtyE3IqqoiMW3daSFJIsWJTIW/WVbxFcKXGeAK5q55yW3ahCXnDSMsF
/dCowOhIzsZoCBH71W/gsG80XtPD94zPuVXrVI66qe/pOmo7/quf+lu11Vj+rx/rsrVrGCAMkLE0
Mg0D5ggOj//P/91wD83Se5N9fZUrfg9XDxxMPdDt7wuY/9SM2Xw5zkPHz2K3LnBggpoVXDv7rmzJ
I/g78ZHaXQBE/aP9g2ZgVMFTTHfMNR+7P1Skc6nbXLc/KIi+m0PCPNMkfJHj7Y6X6mY9rBBqyYIi
9U8FKYYHCoViXKx9QeYNsDXA2IdtlWzn5EzQqG1ElDu0LGMnog9S1ZVJkxTAe9FUivbGYHOzSKaI
MOe3aUmaRl/bEMo2Lc6UcpO3Es9bfam0y6tceT/WHeozpvykAk/x2AaBXpDqXcTwrg22n6Yb/Yhp
A9TRNZJ5UukcKIXpzYXs5cTueiX/eX9aJFOfADmoQTr64x1BC+7rOkJaBg8Huj7Gmg8fecqfiRT5
TRH7EkEHiubdeLNBGramjPifHku318t92cv+3JsO+hWds7JaoQzhrtDblONj5aJ8Sthl3OgYXXYv
q+hzHuFCoUSq+KQQRQnJZ+be1c8fiqxe2JwusWhHIfLHNj0EjbFP+/u5dYFzdUcoCDXKlj9lXiSN
fZTBrZHm6aauDS9PU0LF2Dc2Nl3Jv/rBQnnMxPtpEnZClvN498TGHFfWQJuihP2BR3XH9f17QS4/
ZTUFR5YBjQIGLrBodZolzGvX+F+GXpEcOD1QqFiUkX6l5aiq/fniYyE9YV+ZzPUfn0h3vFwIrcz8
+cPDxQVfGB78dsIbaO9NfeeHiPHp/lPr+FzK9SjGkh3f5gRIzICLJMcI9nSGIY+82SCaQTWsisCL
yNha3kR7rKpVAtii7nsMsvDuUceH5g97hN7p5RLURKDiQa0ifBnRiFHNA7h0StY91PrEdPQMn6gd
V0HANiPDWkpW+h2au3rqWjtucURWDO8azrCwTOkQfudRFhueFeSYX0nAJxwiZnfo5Yx18RvpRz3U
T+6U1jk3JTTuIIWfvHbiOO/H3U4LIkNYeSOKHkLpO2puXTdXC81hzJwsuCGO2TFQZx+9ZK4Jok/T
bK11dmXRXuYf4dTySdmQcLUilWQbB8+8BBk2ZEeIwvOW3SMV8ow9wcsVvd9k9/zf4KPcnwjnYppg
WN8B8SErbhaVyerFGSYgMaA0CCGhJ0tnqtpwmfvUDSkiHJRLXgHhgFO8mTpqQvnefowLZuPwxH6e
bgUgVZL+jRXc2omuEsccZWI2AWhA5L4Nz9h02NYeQxjomq/hcaUHwYtXRzmBFdT1coWDeMYBLylQ
iCfjzwe/wgcPipCA8/3fs/4CnmkHzT1s6zhTHk7npmKPTKwLPbfj1S6hQf+dBdsBSkwxxTLwMpLb
FP2k62xIK/EnSks/9Sfbg4eOYwugTwL91g9IZ29L06Z2oTM3cE3U5nakPFRzDB0oBpccp+KHK8rn
2b/wPvsS0U03ntBmjAySjubRWJMhVguyVJs20zIGxaYIWn0J0ohqDJ8QbNpgh2NA/1gLIwFHbbjy
W6Foo03uURAacRL+2wfrgjFfqmOgyyoytGmm7bC2Hua4Dn7vxZe4h3wucAPVM0i6MFW/WljtQLRU
ZwchjHEjDtDLjg4cu4nSQce61I5RexJbMxIgcS4R1s/j5uXm3aJ1IiqztNZDf66TVz4XsJU8nvFp
RNxvrTHB39LairrisKxyfSkglrcefxgWhRGzcQlB0vzMvhCAHsrY8ICEOGVOyp/hIEYoPw5l9SXP
BLaoJwEpz0//+W2zEg2jDzn2drmZscI6zYOhTr22EccR9pZ8NYUIkN3JdQpo72IfqhmCjknaRe8t
u74MY5m/Ln5PbHsBRVqrBxhjJPjJ+XSSVPXyTI5KZ1aixVy/wlBK9W50NgfGnnkRBL8wm0cJv6y6
s7NxGlaUGIbmeO6swRfezaVGAXVfpj5G0GU484uwIk+T9+QeZbmE7h8ZGq1mPYHjGrDdjPzHj4vu
IeBYTO0oPzG+UUkEl8qX0Qq9wAUVQeNydBH5b/0RWzeNpvxw1HnjnZz1S6IeYvOw9b0rwpeCLpbM
K0QFS8JGGpRsLK7Eaz7ZJ6dAXpNOotzemiToBbqqh6pRy316D6RJtH9eOgg2Yv3SQgJwaLqpCxma
8iTftEUCtl1hI28HxFSanCiEuuU5zp6V3EJLGV8WHjDlUiL4HRShLQEbdPRxzF3ONPmxScRzBJFa
GHydx6IWUcz5QXUAB5Y5gxMG70dKegNZw1TYX/mDJY9e79eSs8Po4KjecfiKx7PRbOBk2MbddAfx
RAoxqwsNj84FWV9e6PViT4rTmnV0sp++TMQwcyZhcwSJ2F3i1OIOyJtwN1QFyfLf3evxl/lo1DUM
QOOyHmXc6519mal0bYn/9VyyLYy16nDSi0xZ4M+TAkAdVIAh23ii9bLNIgXzz0BTEHA+8+EI3KTf
Zc1FsZjE6k9HsrtxqwdNGFuATtlyvzjNekubL2YCXsY2UmMuqrJTe2eSwN1d7LiNv5LHdZ9IXKgE
99n4/ilpLV32GJgZ4m/k2dGnPOWuSyE8E4WFqVKHr2t7NFhGhXoBA7/kGILXTKyK1vpODPRnkZGi
NoLzCXLagPQgGrq4aCeWnV5gvJ2lhsr+IXgY872eRKur4PPUDbOt0PiTM/OiCv44IbAhVPuX8gtA
EmG2o16RWs2vSyBfovjAcgEbNiSRnRqz08/RqE6H9csr9Fs3UmZvB8DdrvdN8xAmXP6MqSPaClZn
GJeT5g0UWSiXF+T9MAxXQxLuIYUWQdaBPfk6EbkgkEyveg4Z17glYGTfr1Urs/9RmKjAmKpu3f+D
vTNo9BYKC1C/qsjylIsXmd1llHmAsC7pvZ367S68scFTvZeOLfLkWsg3hxlwA0BF277rMbdFY9xJ
RJdW0tHdoq2PhdBBTbEm+KY16JIkTgqAOan9WVIo/80mqJVPFsVWTGMUFwwMctbrdCNAR9GF739R
ush34FJ2c3U3lomMSzVoKhIo0mwZ/Ec82Q2bAm1cvud8kJRH4qz/vo3CUTxrKaiQPflxT+iuNVma
aFf3omdlDZ4fqE+teF9IhqfFdwCAm95U9Sf0H4qtmRTytyI7MzlYrwz6c/d1lrJHjB+HHmP5FP/+
iPZfmnoyZn4+YE0od/N2S4v0BJv+E/wNNYvlmiNPXcXyNlnerf5LYRIwmYuWyhSxB+I1JyMda1pm
0vKXbbDnUnI2qxdHrot4jUQjX7qWhS1CkCunZC+5QHqcuHRauxxHUrJ8YfcRY5CZLEsNlmjqMEjE
1trIV7l0lT/r/UcHORAxPeqHpNSdxkjkk692qcPnLqlBi0MQkJfYeEqODtQiNZIF60fPJAEwwedo
SqeZDdO/KgvL7GaWQKcOYb/126D1f66KSXX9EuJB7R+RwIDG6rhfesVHpEtTdI8bLqHdG77edpv+
DATZIQdG4Feg89RKP5MFk/GeGjKF3t6+inQ35Bt37CbRkHX68WACdOt2+zEN95pufHY8luAPdl2c
pd7Ui72a5itFrAsxQT7uoX3SAs2H1Xsd8YJ8xR384gs2V/ngXimW2Bbi7n8VwlPPAmCnSGwfajAh
Fvzt5LMrp84PfJxwokuJ/5pMgoEYqT86CCFSTDzjUjBVe8TZOY7Ym2wU5VI20JA9H4NBGgmKVxfs
931SflwqgkGlIn0t0RNydXWA783RUwEGYcUDPH4SwbyYmb9/YVQuTmgh+dVtsSD74L6Lihhtsh5B
zZTN+DhVx/3usN+gekk8WwT2atz1apwxnZWBECf6XnWzdHD90LxDbauqK3FiubiWN+xrCBsF5gPS
49X5KXXzYg5ppI99AhvaGDxQHBeZ0/tHXUGt8J8Aj6f2z0dF2f3/UMYLKr9iPvABXGJFOc4Z0SiG
t/ptEz2bIQMA31V6AFEdnG0434MaGEXnvf71PpZnDoJ0BZLjM9Wky4osyMW7eKXtXLN23JmvLzAZ
aNEKHW8pXRrOZ5T0nocwyq4sdw/iRSwcIETWZ+lAe0xPRjBlsNkB/bpS27JZs3U/ltqeukM2V8Uk
3dMWtdM6w4Tk4WknJLyCbcRu4WHIZybWRoJF4HyIffVIzmwpr5MlCp5n5bkn4uzdAqJYX+pZ2iyR
EZwkCIrU/chF+HLhij910S2c9xFiGzDrwFBbtr8M4qTwSpOlcEcdtxhskaILk2YKqctWGFCtvB9/
5p+j2ykn4jiGJbiNoYHXtmt7TY/UaCfflZH0y/8doHU6LtG1akwBNl/lKBNZuhXg0ZBKeOMnW4Eo
0N7A96e0dAyD2lwA6coOJv+bZBXDz875uG+sB8yPtlDxNlVPYjmnY9GTfqgZSz6ECIq7lwm9DFD7
FpYPRHNG1HbhPR/DXifHYGJyrCLAWiRUlEOp+T2mTyEk6FpVgXt6Bc/yOonxftszA9qlvrt2ntEw
rTfFMtC3spf5zIT4j29YyYclQPinEFVlk04sQcnujp83fTg+9zb95QHid4PiQMZo5NdFnw8Yi8bz
1qGG0IEESX4CYAlTwaLMf3mUbd6oq4Yb8N8xEH/onOIhAPGsnSj9BqAje0dEbf+xvjqTmIM3Uv9m
IKlStFGhImZkBElxYI23Gg64qp8pYRSl8CKHnAGtegJ88xSw/67t6QqwWZGhNrsW2ZPUN8UQwQ6Q
zdugAUF+hEFM04xOIlilyUdFUIf9DZ5Kr3i6iTIgCSxa0u+2yIP91NLvZAP9TVjd4ea+wZMCAR94
1rOUg7+znTTFA9It+SMXSTmYBDJPYjk5GBUoKS8gBNdNZ3ahfkT2kuuKHFzJFHd8sld3dg6TDS9S
o5u+GRinyCYp6y/ARYaErGwuPNBA2NHKwwTZ0tFgjckELhuAevYsBSVsPAqKQVCuR1ZPAeCbBaN+
XDZ7qDjgGUWYrCt3H+zwWYXm8o6sCg8DMvlGxerVu1w7tnUg71Uzt0DIvi79XoLLDp+jI/22Tbku
xN2MZWzrE4Ec/OM8YFXseNpA/Eju3E5Lp7FflFSgcZUV9ozqqKxJaeevnaw68tSXNuYXh0uZrAWO
/+T9HBlOCuBW49bUbkONVm1ZNGYxwdqKrE6sFNYqTukFY8gm5wQ6iFSMXvRBGbWCLvUoP395vhDF
hHdAnoT0IHhQctc37fvrRDxtvX2zYWbpjbrbqAJOSi1DmIS5SPTr9y4QcptHyOA0jrxu9mD+zVK2
kDXX8W9aksWrrJEJ6J7aOq4np7DFxkLhU16G7O6Du4rSQsdqp4uHcwzLuslihEeMSRLXbMtRGMQz
i/MMv4mm15gjmSm6LEen/h48QOrJIEDtNVVViW8jrhRQEGx3XJYu8pm6EXlVzEbVIjgz7qHGeXhZ
jwb6yeMysQzsl0S2I3Jb+v/Zte/RlQqlr7JqQMRoaHDymOYuazcYde73A+8cB1Hkd2fuU2JTc9nU
m/RR4xsXEFjatoLzxnoy16Gu1i0UnCYw+8PYYeC8s8TZyTcJGJ1W631zU4/zhP1RmaFtQKyz/dMv
2BSzZDqpY65f2/SkVUb+dhiLkKzF9nroD4LePZQypYnSCuP2DuSNBIvNC9kVznDwXF8EwAAN1iSv
ZhdXGv+T2x/O6f8MGwG8FiE7Tsq0m7eMY5cd9RZdgzElDTqudpRFTXS8N71eLAPz0H73tHU0V1Ka
o7XRPtnMOI77I9Nax+rNtXNaFdDKkfQog5iunXByEL4vhWdgnJQQuFt/wLgAkFrlXcAfOlqnmEO6
GwSM+fjoJyhzqX9+fPBLQ920XxIG3ss8691IMcAOSFnw/LkTaF+qEkArRzfDna6qcJeb9xfgus/l
OccWVCWcrUX8Rpi1JCUC6Fdo0OideQsAg1Yq+bsMp+2FZ5FEdhk5GYSZo5bA1oXRgo+FX4LYjZ1x
TV04oNL+UlHxMrYEW1WF500BnMWgo9g1Fb/hlrV7JDm7at92yE51iCCtQ0GnBVhnZPbrE5p3SuYz
MY7MXYDZ3DJDuH81aUh9htKp/Oe/7ZZP/ownxm+xyWO7wVnyZ1Ntpd9N7YcS4wdzTRYDzVvjZnqZ
zh4RW811Ktm6A2jLAmSxSjYtpOsdX9WVNV3+P5Bqun+aR8ao0YaMYUY7tqQ9Tj/pSlauE4jQrVxM
SCCagFLuwatiK8Ukuzxutkg2sHuD+LdykibfoEzGKP4GSF5eztu2D0nYTNDkebgEFNzmKDEJC14p
fNnUcs0Gz5Dkoyw7tYnqFTBQ4IN/PBgiW3UfwNCaZG4xwlnGK3DPT9Mea2jNZNwCWY+poyoOLgqj
+3pWfim1ihcrG95e1UOWc4UKfUrPscq1kUifuDTRKejyVpnMhYoxddw6ohiRJfHibeaivfek3ZlS
VMwvHhT1xlw6na9ThNGVZ1W3EI60X5XV3N7vzwWHrhXY42F82YQJAax5eDcNHlOVeQqEKamaRPD8
8dK2LTlpIEhf1+Z1Tb5UFQLOEa4TqwKbIVkPVc+p+SmA5fGQeEVOplD3fnfIMsWcXegpxwecaoML
FLQtloZHxfPl6ogzunZa8SG+frkH/owIS6MSsQp7dtIhIVO3KOJuKr/om1Sy6UvhYSUU2LEyF7zP
LHOLowsPe5pSJyzUIrvmJspwphsp++YtlR1ghlk+U9ZIgquoEK/2B6GS12cjwerQEL0M46gkPsY5
85Dw5IykHt76EcCcnem8vWxJgGbvzxtsAc4UurGSo5lABYSprAC35ZnfDYsExmrasONgzJaDdwKH
gnLmIVU2OdWTBPlU3ALfX7uXQ6k6IvieGokICHM/aDJsSYCepytywGsfkOvpXtCSnHJ2a894ebnt
TPV9akR8cgke3LQKk9JiUrhAMK3VUPonHMa17C6S5CHvyG9E3fShC8hlufjbgNIuPWUmO9vg7AyV
+TZdT4EerK3NVjj8fDcrT1nPauEEp8bMeoV1769wBT5ku1JjJras5IFwEujo3DJKeydcw4Oq7d1o
5ZbuRYHmqcwjzb2KpN0uKvomFUUuj684fj6XgXv9MbvX5XDVgEi3ng0+sDRfKGDTeyZ2aL6PT/ne
t4q3ShYhf7SqrW2XhjaZMxWwD11DEysF/Wj/HhZFCshUVWdiCnDcmDKhbb7DnmjSx3D0MLLgEp1B
Ogtz+284DChVcqcm2OLUSKPZtbvXA/DPNvkun6yyTj0WpXb2dy/HTjxiQFieNSl01720rF+5vuGd
g7V0fmgKk0CuYYz9CO1RbTDn33sbav5q6mftW9Xx0n5oAV8AeDwixPpik/+rEAnSEgsaDp7wKrsI
mhC23ciEkZUF8BNCQYLRKrUDZRKne3RvhWLzgNAKVruImys/9SIJCjbJ9XQrSAnwKe605AX3oovZ
IWe2cZHp820IOkFdUQLWBkq8gb3STcvWaXv3r7uUI7KWSJ0F+loYZKkgOQBFvPVnSAdEKJ/efsy5
EJXiYJzRFeoLqowievofTIpZlOL8nHxwWyB2o832rYElLNqi+PKo9/FwweMBGGJDXeZ7ILX7O8GL
2dEJbBcHwr0A+ThRYqYRYpP/9GD0K+kCkH9DP7LHUswU6f8YsSZC9MXlXvMG0j1Jw7Y9dT1P/Bov
ZqW0wx8qcJGTCSeeBb7rrXbE1k0zF7SEtK4K3MbDBY1alMLQaGKKsf9ZBKotn3Gs6IOAbA08+9qZ
fzP+ERPhWqqgVT4bJAxqLsDFzuIP1Q2XFPTVtpuDXM9rKVozew/Qjk06tKJcH0HXgh4Lw3bNK+VJ
2JQEXKMDQrS8PdHutuZKeruQrwEL/rsY1Uo+TJ2/l6HLxVcZlItTP0t8FkvsCyBA+qjpGyhbLEdJ
zJJZlRLako9Ju9cNcxd/4Q0l3+GtMePMZNG1y8BhnWqkzHBYjcOZefYnkghZnONVbQ7IN/Fzekdn
Zs1p/JZHyBWep7uiGzk58emtqTeIfv3/aetW7GwFXgeig7AGbv+YC0wy2pputn3Q15nzIk399hgU
6HnA5xh4ikJposGmYXjHMCVAO6TN4yV2Yw2No9/cW0OlHtny7yLHv5uwqUo4T0wpHzaN6r2Igxyw
jdG/ctAye7b6UTBc2RYqEgmhhg5URRb6/FH4ay4faOd3PsQB65MeGQw66eRCh5tphald3m6xXd3F
0IjcfxjPo/yBrluWBz2QV73TcaeCucnVGJjQlbgThf+N80eNJhNZ4amm+0vuNNngLth+DbezorPT
fscR+FmJMETJ17asjQfHiSOAk0mj+BDza9nIOayWCYWLwE0tMirgZSBlFfQsB5LtTePUByasMSuY
B9dXxD6C5JY5QAqHr0zgFOMehVrToFS7jqpFHC53Wh9xMvo0jr20nPqdRY9zWjJhP4PF+IxYsBnx
uhiLrW+01PNshRqy9sGMjk04Bkkgh5PNnLvQ8r8JszthVuk1VqYvRrESKTYoMhV8Enfb2JEv3cDm
Lw30ANfZfVGHDRBmBp83VgdGnDFgSAJiEaeq+NmAZljMdmJyYudK0LHnJa4lmYrhG3DqSwID/GDE
9KhYq2TgomR/1pV+JixwlMDmg7ODXpJzQcsG5+2D6ooBSU6nkR5geUdWWurqirFCdgyESKZw5Z3z
lXbsxT3pEZBQgyaIt6npvu5QMLXe1xXe64IDmXThlQ8Qe9+YzItksMBfWu+Yy0AO2aTuRRJX1Oli
4beAuK4FjY6U/xllEXKS/Jh2SYXKzSyy0gE6aEp7TbMdKkxPoASiiFbtJqoNji+6HVWOzolzJB78
K6IC+M4GFoFOhTH5VjjqbkmpBqMJ6ra3ymzLX4rmoPSofIeuTdMPivBrUjBlkwRzM5rrmnf6Tdhj
bAnThSkjUpCCqV/c9l6xusHt7q38My2HEHSF1H7W6VxNfgpBp/AxHCsrc8dr2Xg953eS6jz9fet3
+hjCW+l0kznl02W0iR4nib1AYqA7bsWE4bfYfzlk3KS41lvdjY/s0+3W6UaES+s+baRgqdlbHgoO
wxM9qWfR7M+pPONLj/4y5vwD/ChlHIaIYwC00XTQ9JkwsJVHbMwrcgMFL/On31Gq0HtKECy7eUPy
+mkF7EcDNVlY+U0nyMSqHZVy8lon8HM6he72RciBG8yq/ltNKkqgOeLmWfyxCvyTNE5rRs0HoNJI
nr9vJIan7nhKDTrzWUNeXL95Rne/rzc1f7V5mtgEFERTfbYYwzKbkileZE1WEb9xVreu6kfhway+
JV+3oZNZsbeVp8sv1K2juFRXhfFTE6t2AJ3GQEQMQd7v7JNOu77iXfZ/YGQO18GxB9s1PBaLXubA
7CR6rkB4Gczgqa3bjvPhWHmD8BHWdi3dQ04OYdtmjkVfVyJl7k7/onAJGYCGICUS1YGrA+SQFMBD
JfRYFK9N173TwGIzVYiF43S0XMWX68LgersVC7QQhCJNLF0YUPHnObeOG6wx099/qidk7onbVByG
NNPKWby8p7cJOhiKzjlCARMc+DGNtoxOifCJ9WpK27HRtmLr84QO9Sml5DWZksSyN4VUP+9jV0N/
zJnlLNDsF3K7DfakN7XyOZPSib3P7RzDUQ3YEZmwo8FNkETtnKngNCHEG1lol0LdnPjIaWRpPnuk
pbxuGjVzlZ3K/s2UpREb89oJFzZdtT9YDxrHU/ib8+qHh5wcpIMFULXV9LZWNNkibSkmKjqXR7L0
cUnjD/8OJ5CmFAPSsaa0/NnE857Eoe1ZJLkqX0K8Q+WhUrP6O6VQL170EAklia2npz0uj54fv+pO
lEXQEABlCpY0lQMptqq945qMpvyDN8lmRLCPvPfu+xC9pqR00R1n+/Fo5nqgiX7af7IQg380Gk+w
BwrvA178Vg7leqA2qsusbXoGvxsnE3kCp31m4L4ycJvhSw8st4mJkOGGng8gdhDvJW3KXOHln3DS
rqeo1vH2QOBRqJlvxnD16WzEKFwOQzzQ88ztil3drN2rbTiqQ1W4sKzqlxr/4gf1TEV2QaDmgSf/
oSul8KLotFVynmL2JVJcTK0XRfEXRGNREYV5fNpxeciU+rDqMt5aBJSbDD54WvCwAkaD4O4aWqIX
bI95HnMuHWHIIsOUvs1vHrxPLxsRXomkXK2T3bWwhmCo+j6es0S2fSOspZ1e/N3rNeqvF30mroKJ
+yrzbuwU3R1rlGlIioz5qoINyjiGv2sUP9BF8BYmtEth0i9gJxH1L9vvvj3q/YUHdPfQsEURoseB
jQHGobEjgXZEaSZlvGHLNurMNjL4jw9mMLUUEyGO69rimCAsbubzqHs87/9w2fqIscCxIx/JUfkV
F6gCWSCxDr74B5UX5QM/OBg5ii1iYLWIdomCo0Y6bPO3Qgn51D57HHnOO4qAUy8dYAq+9AqyrGFw
AAMQixKJtdb3YDbu56tqAIXqWsg1e6t8nPK1wvgKbVvsmiHehI2t4L1rEREBr6SFAXlsCeaMJMQC
Mbk056AWQ7ZOvKkoGwq55MMM1MKwYy1stFxl/hty91klR1MqfcXmW/5nrzPob6e6gPlcuS/X0h5i
1Dv7ntkByo7lhAFneR/XH5sMnmbHWqkmtv/en2QvD1Pqy9JqSkwXrXxLbR6acm+lQDKqY1eNnh9N
bHX9qBG7q0EngOHhuI2a5y/7dYPOaP0+PbwzOTe2aFLVE51btxmZLGZaDn2yZJ+1D9hEkn5opEfh
LwC8zJ+edYx2/Xz7w/hHfQldzrMQlGlUqd9avFrV3eMzJNJvcohndLh+cWXzMHv0+jS2bSwvuaDT
F0hSMJL2n+KW7YnBnW9XQmB7oYh7XLUc3/FyMO+y0G+Gt9WdC1so1OXVv4subWGo729hXAGcYujH
0e2BCBi4H3UJ7BweL0jJvnL8vbbrNOHcvWbgD3R+j+pxI/i4/n9OfI6OuDhhQvYzo4mC99ewsJSh
zyJjsqwEuSx1kXkf30vzFb7jDmNwNU/IRtANYlKKqbnscw9WOKecEUujk3ZRlcLWXmpLSUvhp4MJ
TKMYXJq+LkmpE4p6ZmF+4I+SupMrpD//ZrvDNMXPPM8C+YdFoA8OOaFjYRfLbrU725khLDh3orVf
ruFj9gPc6TRn5cqFalV+m3H5zyfLcYG8X8JQNqX7OXla2+ZoZkjOPpkrBd9sBM6vl4zf+2wpPfgK
MPtmNtlGik/lpcJm6f0zL8Ij4SDZKFpF0vOvIzAOuH+sVPigC0Rm5A6KUycEuChWuQtyKHJ3wz5O
w9Ljm31E2mTRDcGgFyE9kAJIHCWUns4sEKNE45azCLbOQszKY0EeXJDaTZMrZZ8cPkqRwuOFCEV+
ysEaMUzh7kCBWmOFxJ+7cbK9sOCblJ7xvsdlq7KHUiSdOWZPOL4S+Gss7s3FVSWGpQRA78uYXt0f
ROcz7I9ZouRIQq8upCM837HiVWD8p35KpkLD1eaCOWtMAfuty3No6lgQCYMmhE5T/KDlXaENzQ98
uO/DjMU8eNFOpiIiqBZBYC3cbVfaunOcdjwD2A7p0Sv5Mzip4g1xZMuHG6aSYngiRxSZwUCV3CPu
jl7+VIT/Cy3ES00LByFku1PZ6TOyiCK8CWeLAmhxkQCx6dfK56no4FWcUi3nrI63ja5++fqlZv4J
pYYATtOZp+MV7uC5n6K9TRqmwUqZRmkIXQc1pZTHmmo3CC6uEbQ4IqCvIt15YSe0LbcF6W0sIXBa
QajjUlMBr5e4n6YOZz9+uOyQ6MhIADT3UHsqlPZavJKoEyzOXNvvPa21qwRBrxombaVp7QJDhgNk
voDTGNkSdba/mIOqBVgsSGqrqo320rkv8ZZZxYjx/udin21NnA9HNChD+CgxuzaAMfFbRsug0Mp6
UAToEfnqKss4VID3u8Oin22/4ArXqCSKl/xxwOvDlwb7RH1hNH86z1n/t4rNenx6qEnOKcijKYb0
l+aCTpsOrB/aq4iIGhcc0m63NuDpSYLKrCmnINgk7K2NwkuBrf+IZg7s8Kwf2rN2Abr0V4mYyYWX
AvnjjTEHemdbTOB3z3b/cbegp4zx9ncMJI3Ir0eSDS2/6k43XC995OAtHJpwsjIgD345aEg+vq+L
1F3ALWAEU6X5MW19sYBQcRYKiuXa5PWl5SK4cLKcbeqW20/iCjtoupvgCI7EqqZ4QsE5Fr9cl/Wi
0vAK4+DodGM8cgPVvAAR17jR4HFl/Hbp/W5NVMDSORsrQvb9+bRJU4QxmIbo3HCYk1f027L9ovgn
x8uzOjbAJfWgzqjq/RD1DcbCa8QIyxPG4s5aS85+IiAO0rl7oTQmva1IuOoXo5N7HKkldiX2LuYL
QwldAFuyE5ZDkc/NJL8X2fdA+cNcjdhDQNx7xnHXKwvAO0AoMLp+1PJztsKDp5RMHBJe8WA/HIiw
lh1gUxmXFhkOj8O3WNRRn2hq+17+IYOBdxGJr08SaPdePTbH7iBKgrr/sQK5/VHPaOob8LUUdPDL
re9hmSy0IS9JU9pwsO/mLrgqsv/LzBTlF0Br+01ZtWip87fDWNV/hg//sBm+4K71hjBbUMwEPNDU
sHjDE/J7C51i8ZFss3vR7Ll3r/PbY7Jevlf7ErIO0ZL+ipvDMKU7O7lldtdDM/E924UBgSkvL1st
r3wJldYSeBjHzY+OhsOyy+D1CUnj2Gift3eNiUDoMru1CQ8NnFVuzqztdv6PTRdgMlnD/6rQoUMv
1PhPz0NfuGB9j+RD2IROaKaeFWpcvdZSrwbgHdNRCyZLT8mcRGgqiXAaDIKOMuKC8HCP/xEsTZ0y
+OPY3yVP6Z1y9M/rtl6ibmIxiySSxIEs9tgK7Z6uHzGO/A7RWqZW9jg5BJqpCVWr0hQs2wTmwHgV
W8+/rR/S/N07AE6fmyyEAmyoZ4mUw+IOqNJynK8qO3UyQvMfLXoaEutFojM5+Pueza73tajjABFi
BdReYKTJNF9JQvr1M+wgV49GaX5bbhjWQwOlPEJlth/PIC3AcXEPaKG4CUOc6uB04i0L1jc9pztF
GUTMzq/G5QBT5pgM07Py9FbYBNOg6i207/xsgOC6JLKsZTMC/jWeNIefJW48BJxNMB/TPcJUA1O9
QesoEX03d0Qxg2dK5IE3RsIfCsDWF95+qjMXiDgdHi1SrjdqRnqJxTpe4nQP4uYuy7s+MksuKBws
4F5LDbeQEklIMegVcha8duQaetPG1YEwpXQGfTiAN8Ha5LdfOH0X3YYRWjNhf+v9NXdJpTuWdZ2c
BrAtuOIyK8wJLjz8/Vx6kKmlDKqGmWSMCC9jFvbHY3Yb1ICU7uYgDaaTJBV2rmOio2/rBRpvgezr
iHim9sphzQRbBTHZFQiFBN339CvdrcNLI2RCEf2sS6S3J+zny2p1LAa1ALNX5gxU1ke0rKogqDaU
InGkhFtWakRAu2eWvvUEivaw3pY1sCylNv7lzP4gvNfroNvdtuOqql9UuAuoYOrMtrq6zt1c/kkM
Zkmai4FYuwbnpE72sckGXzXTZKZrvuI52i2bPelIkHWp2pU5VkF2dgV5fNQGuYjtJLSicJ1hxjZp
Ld88Sfz7q4KHws9CtxlxgixH6jSAcPiKJ94KHu2DMSLeX9BN0M2HaeKP3aVdziAPE+8SBkkHgL3t
j86cu7abwtG8TF5MTIQFm0oPKDUw4WsipXcwB/dUccXJhZvKQ9c2RxI6ygrBVNvpcsfv/fS/CYEt
DT/lYn93VDgwbtf03rwSw0Zt6ZQDJdSZgxpNh7pkPEOafnTOJ0fjkYjo8t8bugYIwVz6aLrTvESv
g7PKCWDz5lKRAlh6ps5APmnrSgQLyUGnsRY8hvQGBEc4Ps+5vU2vOUSKAngUb9qiDQE2aIuGCmf9
L1lOe4nqbBifzmRCfDagaiUHeh+rF9EyUxxkB2qtDRY9jX0mfDCb+cuX7xmXcXsagMW5foDz4dJi
S9HJzIJnOeFrXOyW84OILI0zS7AQOyf5LLN7fEmSNFFnw20TrNkDP8XL41drUBobNPs7cNQeqYip
F050NmLvQu3X2Tz/p1OsTTU5wiksaaUYNstAXol47oFM/z/tTOo/j5wUJ9vPFyZWK5RcQGxHrm4d
DAcDFRe3BchVVddtpiMvYmiQ162zl1wGaWGbCIqBK7nx1FwBQ9hBYFO7MkBW2MJK11uCzNA3PFAT
HMCBnuu817wAzD+HBHair3fRdYS9rkqrTyCAQjoT6Sh24Kw7iKByIetOtrJ15VCQoIUFoM4iFwcb
84leOcGADYdcqhjOpZAquMHpCefYrZ6DlX41o+7dLtb50/112gLw7u0v7ZcPfvAiFJEzKhRaHzch
FkgdoZzcWRzOiGMuu9iFcnpOrNkkQzQtMkJrW+GdQo7SLt8kyvKD/gBoq0swmo7kPbYeInykyVXE
k/wTb76jhssob/iLoxJP2g7+TFaMlTk98rgFmfcqeOC+PDIpaWilqZBwcwX3uGtdTdRCW1tll7Me
JqtwY5JD4oKMqlw2N2IzT1ziiP89EeQQT6MLWvQSyFutOuMjpAQDlVDk3EMLp3ZC7AmYO9d6AYOM
+h4ENULogXO/DmPnoGIRE9mYX/xY68S9EywqSxGco8ZlcaNB0J+7M1E6U70X2WHwAMMKdK4caMoi
tDaUxleGucMF8GUFHoV99Pik3aPl0BAsoselMDlqAWSBxIv7O7aCskgiO+YKabhr9AwBNiLbP8CB
PfNbJF5WrIhurltcnnAlYxpK0XOxSxMVHtYlSMCfo7VnK6JMastwl6e7A+Gf5681Kq19dWREEtEE
M7GBmeodRke89z4bxP2xGXvw1FlQCeAv/tY+oYAX9IVEyatvdHtTD2w8NF6H0RBZG/JcYsAaL0qj
KG23yotl0383aIGstge2TmaC9qjFHz4xgW8WgTxxWqymmje+Mlw2TxBuhxKYM0xss1z1o8mHeZl+
QBY1r3KFZJHhER/rLvxkfYAGq1R4utHubt/vwnd+2r1gH23rC+9/EBcK6U2ZLwbdDeY7BEpBszDE
a4aU5OiB+hR9uvRCA7G3PVSSyXs3jTHwigGLtHGsEdRhiZwJOUbB+ZOUg/jP8qsD7T/fkbmHqg8/
tnxJbtGV75jmEJY35MFnik3FiwsJyL3dNIgttCGnRQn8r9uYaMhzlZQMa3WoBnQWCqqfn5qY+1+D
0IkagNb0gk5tzz2uPKE+2pnhKU9FkIPjEB1TimPey45GiCzEhYJOXXg4ieTinycE0lfOK4F0SLnp
7v7j9NIweB6sk2kZG383OkCiHF7JrHMvgQadK5EPuMtgpZVl04jOSIKfN/CWC0fVOoTzYWDNMiqn
439uVr+Zi7zDbBqEJMODYjZ4iHhhky0O6TVlfDalEdwmVEcvkbvYEy97y2ZAO6F6vStrJlbJfNnP
1WfGHaGa1dhWFn4OuSR/LRGnROhmCtlfcTU0/2cth5XGI08rCRRZ3QIcNBZLgnMDwfxDhTpHbM/7
XwMtCS+y5NcW43Weec6H7VHZ0o1ZZ9kJEP35krraEpI4yzOs61imh+HGDK+TJ5gN5oD9cBiJwUMj
c2JAEReYiwGJvKia00QRIGdpABqvR0mKU2vmN9unwTdAAvpmkK+W1EC82nKojq6VH5JFs/m6n/kx
7MklLyx8e6T9V6fZ7YpyOU8+YtPu/Pv+j0ImaewvUIj8bGXEv2htPqz9APeKDeKxrmM/SGCRvuv9
2qwCTNLQDlhKQJ+IfpK+aL6e6ivwcooXitbV6SZWVFwsLZIU3RBUgm3O3VN0K/bPKnkpdbzLgz3D
kVmqmlRfWDktGE8aPmaVfvwTDAKQJlQxM3Qgej7Z+YXhqEqz3dmkFSxDel8JDRlyoVaJsaDmt6th
gPuGFSddpxxGN5y0oxzfUNEOd9LXDZLHnHPR3LxxA9xvIbWRTskdmR1d41X3S1znLNMVb4LCHkVc
9V4Rd/8XU4bEAkxYSMtZvNIKVjWRKe8CkbKmvhIk02AwLhcrWzEaMWRXq89cEt6r7dIiroukFBrh
WTX1lmQVoXn25Z4M1gyUyl6UcpBeQvaOhSLVDYTaBvSW00uHBz3WVu5C1RK08/Ny0OapDmUDlSAJ
Oht5HB8yOMUd8Fe13GK1PYkxC3DTDfMPQ7oLgdzkjhgaHKl4JZR2O4mNf7rta2GWagCuRaWxDwY5
W+DLaC8Q0WpAoZdG6nUuPlpclxFxi9bEIBGYcQsZisXGYIiVwtkGE2YO6b5DCOHDfMys2dMeoDwK
zDDZrksjvK87o9xqwXr8T60uLU9322xAQKdH4xeXD2WQeKm3jo+UQ2tgmUWUyMkR9v/wPJFBprVT
AzWM9SW64nNuzEkhttyy+iReinm5l5sWZpKaXBL4ZH8jARKbkcUll3wYfzDnTEBtDELVA6ICEvE7
jfhRLUbzQP5tCCTdX8CESiMKWcUHVNY+/Q5qCYow5KPynUFyP8FUBbUirJM8oB69RINrkjprIU/I
MxyTo4oAYZuY1R5E81M+aAZA5Wcbw8BZIONRHAFRHAEuZLFIORoFX6MtBzAbl/jqPainm1k8nQAI
YcWghQMMM/GZo9e1rt+iCmpcYOpJltH3+ukpRLDm8DO281r+ffHAvb64LTxaqlbcgoHrsHwcWo7a
McPCRaEuI/dpeGSy78B0j+Nbn++xUdv+x9dJTQxbmwbSgWG6tO8IxW8vVNPN+0HDr3tzA7yAvL86
dDQGDnHurS8QRBpDbfvi1tFiIiwixLi2TTGEBtjEaaKtRtI99z9/V2Gqoc6imRUi5WNZLj1NkrKo
WvDIG2Rg23MJYtfaIZN1FfimbrlNdvOPzXyJArdaxdu1UeZ5ZqfZe86AbVa3kjPKQISMpFEPn8ix
wFXh9dtq45luh6CIkTVmND9XXVJxMTfVmFBtXaW14qYwEWu0TFBKSmN1PRG7LS98Xb/3p2V3Y1On
v3p5J4wsWs4HvIAsDPdtu7gZ16SJk+PishJEJBvuyjtOMDu04pTGZ6nx3Yo+MhLvTe09CN0mERzp
Laheg7vjQkQWpK+nNDFgC1CGPMVF6UDBf32hQWNp+Tvge7lC7FmuVq3wxu8XlWv1/wQ0zZEi2smm
lHYtvS90cal6WnsWpvR3vvF2ICjeY6aSXRHrwWe6N+xslo3aMWwn56ZcZ5DjCurpM6V59VRH/oJC
UXJwMO/cSFWgwd570qFo4Ft2akoQCgsFAzyjZMTKhNQ2bOOyXG8THYuySedzPxpE+MQ5FudKF2BK
/JLUNMyDRD0Y0e/6RNCgeddTR0Ak2ruD55tbt5W1ARerd/R45bpMt19M4DifwUBpCsxST4XjGt4t
F8IrsA9kIMQ7MVOlcppRLOWoaLLceaFRTPvZSo7xTiUOeONXh6x67UA2o4i5sWR92YuPIl5AJtYq
kWLRU4T8EhBCa5BGbILIie5qbZKoFgANzXxjMzeWGpDw/SypBH+GwyXYrGMW2sFw3bePiulXzLNT
1VMNPJyLWwKuzeQHRjs/EWK52x87Nbg1epnXwaJvT7whfAqLhzQip1MmbJ7UZUahFWunCpQfTYKf
a9FUJTD10ylxxU2LPgKm9rNucpzKO4Brw6oj3kh/I/F+tXBNr8tgnLHMnp0ADLH4ySZyUPiBgsad
gC8vsd/y/vOAKHqFu3ad1I+INSrEFNhTH7Q2BBxT7fc8kUcYaIZHHSGZd7BcfXxbrm+14dIC9k6N
LUk4PA2QmYW8qxUZDwMbONinFWMUltMmf868mtnKK3IqQJEwhx6la656Z+wVcTjSn5gysegjuHWr
9wUevgT9wAZBMOw45Tw4o6bqFXsx4bUKtgQmUA/bg/J1HHtAPDIdQQv8cvdFDuApv2SOYm4qmRlY
8NX90q6/5rOjR7WX7fwrKR+gOckUI5MX52JuzBrdfSBVpIaOxYesV7hrqOsie3NgwiEwWw4LN3IK
Gc5qVxydlUly8yReuPmZXLGjXHkOhxxbvdrhwjT/QaiasDOSnoj+3bPAl1woAv4iKlF7UiFw9Ng7
540Z9EL4eEZuYBTaiHn7BhEcrRBW9mtMKwwd2xzwuFyfgixDqc+yCxBJ6K8BlKlnMWKQ97CDnLVh
MBgmVQfRB9qA0rgG9UP9itnGm/aCjkoAOGrX7PSVubD42qMH4ia3ccKOYiQkxp08bqjpdkr9v2Ns
1KdLLCJqB2+6G9FuanWOTSwPN1xWe7HTlSLqoG1MBTZCg3vrq6Txhzb3j/Ff1TRyUnsCdzhvh6Xu
wZW5f0j0/pkXJMvhU6baMtRo/IaG5iU0XL+H2rBt+BNIDX99prWRXDibS9vUdfOMB7IC7Fa+hUTf
i6jgDzKJXi7Piv4SWfsFwEQrtNyJy9s0R6Q1bTYC07+0pSd1KARbCBlFpEYBSCefvAZxE4EBt2o4
qozHz1pz1b+VJcwM4256pNg6qqITt6O3eLl306nFv0uhASdLIx3JusgliQLe6mYyVq43GcKHbZLc
zv7G/yEaeTKsYrCVe9YbU6xiqOxqzVWvhbUkpOUhAiVYAfFxdt93iUTGApIvfpRGMEYP6wUMvKBw
OtPaPzJjtPFPIyIl09Jttg+LqOE45DN8BpMapwM1bnP2qu2TqNL1WU8IrsmL+jZkzGV66IdJfk9x
E8d66VZofn8wksqvHFazhHr2AYpkCkgPPA9NvwvrUc0/Jtc7Uj7EoidnA7nvqE+/iB5yCVaAmEQK
1BNwabDZ61vTOsctFg78u2VdbECCNQuHhmrPObbyjYfybi8LBPjKU2Ie7CoA2MrU1zdOrLynpXtu
w2nZyDZtzy0f61FGBO2/qjIn6hDT4hIH/sbH5vdhMRSYqQxlFHNQVF1y9+5/YCq8MorWoNEDF3vD
wen9mzwDj2GCNXH1pnV7kIIZxI3lGatuFfXQYO+PiqXBo0OMlYPD1pCaCi9NJ/i41UUL3CPv7zrQ
CJVEq6NYtqomxEpsOaLkd7I+nDsyt0xzS2e94ZSgjigxl5YY117pkwRPeL6bPz5sHfOFk93bIgkT
Ya48JqQ73xN8KtTSQy49tYdpX28bgc9fWemcSoqynm9vLhyt3vin0n/E3wz8FNFUKFrBy1ppT4JV
kXD2TEl3D4jmjHUb38rQWe69YrEed2gHrW9/UeZHPrtxriwv3v7B813NDaIfzPVOFuaOM+ywOrSI
pqwxBMOEkBzDJKmQFDquAK+zuBiRV06FbRhCcpPTeshkAkGAnUjzf3iXa3zuRgQSNrYIeHfxRHKZ
TcW5iCiqB8U6MoYZBTqqfD45WoH9ZLZxU+ACP1tV1O+I4jof6HjME/Q1M8vEPtzVyep9GQp14yat
GZlHrLOw6ZcfQQDpIGG6AnuZPI35vSmcUDw24G/Ei57mc6my+nOInT5gj+r4cUEuIK99lx7Pn92N
9y4ojja0KI2DdnB8B4ngF+u5lqCdcoxzbHyowAqLzYFq0Ww6p8QZvu4r5W0rtqpulL3W45soqguk
I5mLGjwpPr6EhuG8xhHy2SezP2bwE4UoR37mx49Q+GBNYAFzDI7M9DT8cIRvO/U6Kpx6lb7vbN4Y
S2i9v1UQjDhHjQkQVU7eO4S5FUQymhO3qq245Jyi23UYIEXkzQz23ssd5Vqn+zrCKSWv5aefdYp/
ynwWX8hUZb7o7crOxeH4yZoXq9ytxlw8MzL0uPiBkcMkW1V4ZMCef/2iBqgeymM0Q7e5SgqH1ucr
It4Nxu8tdjmmeuKYXIhQeMjz0s4Jp7QQ9VAh6IklM+FNiY77K1qCBD2NvyzoFDMQWlTRPf/f+gPX
mk602JrV9xqVeA+6iwFR1ko3ommZKk2GTqRLxlJZoPniZD1FRs2jDkmDUqLPnAgnMnSVnNS3CG13
5x0gMo7y4waLnPeovLl1ckMH3kMgON+o8HEwJyRKQ5436TRsS6RIMXZg3zg6RP5Qo8T88V6STF5w
Se08FiakEnePVA6h9VM3ajMo+Qc6rVpfGTLIKrJdgQhagh66OL5XHQvmS1ke4NjVwvKKyaBiDAfg
8PAVmaHuyS6GXfXl+lFTk7V2JLKdL7XtGNpom0KkiQdMLlId/eFmeiypGp0tyTA2QYCsP9IRjVfU
zafaK26T+Hjws7qH3rSwOvpQW0WH11jY8nOoeHYMrm08JXboR8WSHsTWPWtwwkbPWd9vaCm/cpXN
d1tkuDgfcAXsfiQpVH70n0gUoSBastOyn4s0I8uuu7IHhI78/LY+QtpsfHDoaEyvrShdPu7FShmC
M/aO43ev+N0gVWImgTU7EsuO+clQXxcSP/JIssNeVmyToUlFesS52K9zLHircS57jMj1l3gmtLTp
1arNx7ZZIV7eFDB1eQLzm6VEJFRQQlL23jqn7A3ewrGAo/adjKOq4nLFb18A2p2BdhKC0yvkBI+Q
+JcAuaZ6hrCA+HGhQg+cImiDafkWw/gMS5ss2Vv0HXI4hIQGk2fisHdSS9cty9qcVKKtkP/8MBjL
QSu3wtzVzeOfKZ3EHk8+WGVp3G8q7FT8Ig63cQa58QszpHR8cVapVEMhl3EQaAreEnEgDZX9BXzF
m91VMjNXHSNHH/Gtndl/6LaD0G0xY1aBPmBwGKEltz3g6QaO2MVyDyvOCEXUMVDApx5io+cyS3oq
FFmjHZvIu9sTLWaTFiPnZYfJtxs6ZjPQTrgaMR5OGoi+9dZW1qHM2oX7+D84PH3B1hQWkFkAJiOJ
A2zwGl4oRHvU8mCEDPIfo86jkyvN+wCLH8dDCmcwrIanDXQ3K3qVTjmeveIr9i2EP0XwZxQaL/az
kzYqvgYsRMxuxJZ45unOgF9MtEbT+oYOMQJn6xHsyZBkdoNpEBQWra6am4bZMF7uOHXBJS+lDvcQ
1km0FoMtmkqKex5b+u0MO9FAWS/6o6cqt+aP7vBSNEmv1ptvKUrJAuQtrTJJcdorOkq3g5nZDB4J
4+1P5MqqhNIRYWV+A2/kb84jvJfLZPGPVzwRWv7xRvU+dBjOnO8SqrcJMcuB5v4QG/x3WlM6x99M
pF1KttNMI7jFNkHuhyqJEqwC/29Vn217knfS+YHOhU54FENAt2Ticf9Asjki3thwV2ZxyH2YqV8B
KohG6OEWop+B2Czki7tHYyy/sPmimkmHGtVOIoXSh11QzM7GF6Jug9tWiYPig9UmSI86t1t3RamB
j4eGIaS84x4oaKAs4T7v9zFzC3qt4IBYhVfPtqMl+ssH0y40SrkTiJIBKfnzRKEPpH3nGVty+YJK
/4BXRw8qk9hI3GQO0toO7BlgWaKdL0sYgAr7U4F0hGMjVz9+a69WIR14Qb5Hf35T2j2mdZpOt92M
VKXkPvtB7mWWz4K1mpTTrhvUzPHYhJ6JVpjoXlrvNkzDBoRm0gVJDQrMr8mqznrX3ubR7Jiq9hjd
YvxP5lhuw2V8NRwVIdfNbSldpghNw33TsN6gvDhn4lz8Wt/isCP69l+rWdyUJrTA38Q+KbVs7jQW
dP0UTEhp6iJ2H3QP5AegxfRtwjnRJsuTuICbShUj37vhhSMkgaUEMcjUzG4Clg36tqfz2mD9qjFq
JFP2+jOYISQsGS1MBvH+iL387dhgvPhtp1bKOnkBDfJuHHEXPEk89Bciji1Ikxnpkf+/dCC/fEmR
DsXWKqp4gOKGAno3R5ea+vRcUww7WyjurDl7oE7DAEcn/xY7bi5FnEVuzacj9fdeM3JDLdE6PQWg
6p0EhUpdazkqEnQriH8AaYr/rK7k5DMa4wPQXmI3t/hBC9oSYCJeXMpN1W07iIkDOqip2u3omKTR
teC5MJq/ZNlYrUbhghxPDhvOgVcdvk/Vs+AHjStJ0EQaf3Psc9f2x87FGJgUtm5GS4VKx3e+V+L7
gagX8sCuMtFAz0DTuFj7Jlr0Sp/p5+Vm1wFn8MUqn/fZpWAVH8H0c4DxykNW8yswJArAC4oO5QX8
1HQtUXV8lmkFEvfU3lcrUnrbCfwCTFLAZkVTKpr7RNFozTbqXrWFNdFd2jhL8VZV0VzU1MvUizJM
t7mW3clVvDhZROVQZbHmIJySDuWMuYNC2oObRCyZ+YB6Xg+ThXv22Y/UYEAWDoJHB3p45akwfkdO
+2t/4mV0HkCxoNHjeClW9ZBHfGHG2y4AvZT/mZLEmA8ruBEoX00DjG0hmSp2e5Hjie4ZtEtwmEOv
ji1Q2icfd3f8AiOARenn4NyyYrlLSKXC03BeXw4kAVV9YkzNrd91GiuED3R91TKuhCc/VIng2LT/
QSspcjhk+CCtK3/Y68+jjilJS3k1//zZeCgmjcr+jiYEgafGOkWi8vXeFwgxDDzNGZX28cpHRUdG
dv8RYP9P6XibBgCSMbwVhjIFmyS6wCJlBLnHXqf7vAeBLSBdYJ05N8P3ZyGZQsOh2Bk/q1waq0ue
ZikLjg6IRX/qCPYCIJf7vluf4d9fzCUVa7h64EaJ6JPEk+L/TEFSvaV45RqXF/jxrg59mNTzJA64
UxzJJNTRN/FP3BelusW37ThuvFL3J/yunT9GCAlxz4OXn+UOvP6HzLigHJdp+injX9MSRR8oKzlG
QyPA+6o7nT3MJHSL0WxuL+L59Sz5PPdDvrc6HbSRpow4dZk2aWJcPsQ4+3CKkwt1O3blSo8V+HJV
qwwiSD9rk0/vIVT3T08a/rgqLy0GFwsHd0+Hil3djECnYVLyTJWigi6FlH6dR81sdwANq4j++9e5
sD2ogVOwi9WOuSPXTRugVTwDr+1NiLAsz5+SgApTWBPYxsCQIzTKOG1h8jbnLq7qfe4tdjcPItxs
omp9qeHOdsm5Cs6CelPLUCt56WgXZQsw4+dltM3jN3jVtCfOBLl8WRygK8wlC/qtFTkpoqP1McYr
NeEiUe/mOyCdItLxKQ0uC7ehrXXTnbeJn4zyEyY3HaRJ6VDplaAVvNwmvhNDFFyGELX7H6dXKDOh
NAUKwEd5GOw8LTiq/MZGUEt1jIkzGRBjjI+J1NfEoDi6tkMLb5wnaE8+ua6jBlRxECiXwdniCsis
vcUBv+li8g2jkqz8iNBP00uZ4ECgRlG0ln1qGavGAtYU4UwmrviQpw1DdVAeG5qkOvY85WgvgBq4
0BA3S3nsEDnLgnsBo7b5uxAqQhNMI+c+IMSU7hoPzFiuuGY4dUlchKKjrVruJjlb88MJyV2Eh2Yj
J1+AxeIo7s/2iIRoELV30n0/PX7q5DM5XmCgm8FkVnQWbXK3axu96LVKJgVsC7Z8FPiHZ8QBgcq6
XFmh9oozGRBWZlawTH0c6fBXRPgpJPIwui3jZMKHKrslZeMT0O42u5YYhCOfixVZEvW+y53UBId6
TM4CH6FdE75Lm1NIOBgI82pLgAny7nXmBEcoFSKaJ2+cWP15cz7w37GGzHLU3IrDnnkEguSM3qKN
LdwEIZbzS3E0whkIQlj+WXWwSDl09a+fbyRpxTE0ilwP/PzfBNWR2wndP8T4csXDnN+DWWmJOKAu
DgJ2zsakHbz6e9MvhSDPLrPPr2QX41SVIKXv75c03HHwPoqSsMirNQTW5Cbbojduze0rJ8qQeQXr
OfD3TngL12aQe1/rdf9NYe+8EwqHrgMBkh7cRKwwmt4sQGZgZq2ffjsy0ngAX9A7K3BioPvPVr0F
nLZdAmgtpoa/wguHeYzgyM4x4IchXgSOIYfyB9nTQsDiW1oQK65sbMV+MhKwVvYYyI7zJ+xObCVA
9gyEpQBYKYY9QPagbLBd6ulLU/pApXiexg0A6Fdlj/k2EY67Z3penVL4AN37tFk0hgW8MGatrIUJ
R5k1DHBhhyOkPmC1PAgmmcfIInOIfDd637KZrNaOcijz5WKEjDv6oFPF5IE0uagD2K0pRJx3SiyP
dD8pq9ytwZRKfr4PISfcOPWjUoMg+k+aWSSN8OFJNuko1Ns+Ox9HuDCC/WITuSBQDdkOI8ZvQiv2
IRpMjEzmjBFVCSPo4KQ+Ximdd0k7aTslWcFwBMabcm6F2Ig5vLjsxxtdOxsiaCIKnHsI9jOc3Syr
chh/ZjGBMXffP/U5czxRXK0i+rAJ2ciZ3WYcKQ+gHO0S3OQcRrbssTO3h5afkTzb2eWkrrgwn12M
hUaQ8tivRyC4w4QIhjZxTpVRaHHEnMKQiJozkXQD+6AYdyuQw9frcdvPtVLLihdwh3xrJrAm6wxr
z/8YbMh2p10X2L+Osr2bebs7Qzj7Qx9twhhamDTghKLqqYb9RdY6dcCesMbIeq+GTiH9ywrgyXCO
C90liYBy9TtrNqHAT3s/c22vlQCJGppyTNNU0Wv2AF97dQgYa1FjtdHOXtu5CnhAa7vxmHDIdUsV
8vZdfBlXp0qADiKhpMN/gvuelUMB0FE8UtCJ+aA6e6UaU+d8y5SPTMBemd9rBGAga+JEsJmw301d
KZ1ZUGaVHVlUEOhR/anxTaiUVhHcS/2kHQNm9ipM9htaAZBdY4Oh2dNY2BZ7Nbsoayijai/6BjWl
zjWmjhy3m0RCreNjAnuU8Hm1eNGaP8MwQAubgDQKLmry3fXBPwXGup1a1Q2wJjrA7y42+lthd0hD
q4wA/dZpZjKhwgxItKLqK1K0z8RC4al+IaIoVgSAinus0KkCEZ1pu7ZLcPfRJE9v2pNoWWcbipd3
Wmnpd6QhZBvAUBVvZ3b3/wODVi0cErn4YZgkOZ64b7Zx6JgvaiwDPHfdxznkXf89tsWVLfp2TtxR
8oTqISkACaCb+lV6UP6LER+h7NdIg4wokpgBxTfvWVx57suWacm1X3hEPyB+J9aEzr9vhRjuYN4b
4IlIZjmZZy/jJg7ImOVdY+HpO1CqgJVVbroOFl22HrdzBhNmpFbp/t5uayxg8Jp+tRTaPHsXNQ2F
ljM7k+UKbaJK2UmGg9C1kM1lYdxSisCMl4MWhaqK8jn/ir6tKsaTEkrbJSpKqcVIPP9vY/IzZVnP
4+61ryw9j+F1aEY+f/M2Z3zDcFp5jIR7fC5ZnYG+0raK6DZNUSqIGY2nQM+BecKYPfkZ87Hr79P7
lRuVn6I/Fe+87zVHAY4DMMcUQvVGD1G7mTs4OyAWFSi02Qew9z1zlAERekJhx07FgOJKvHZzJSZ0
2mElnqJp7SHZwCHwANM2Z5VY9KjlSLN0WxJ5vlhor7Jx0fvNnwmjdIXV/A99Joz1Oo7CjDneCpLe
+AkP+NqJFN5E/Ki+1P30/nrSZ3O7f3qQWZ8QnaiyggczorZyNK986JzUkN0hLFt1ScpdAP525kso
IZEDsj15tftbz5J0utpJnwOJkvnG84cCYZBZCCetABBOlgPKSxbHj4vm0JVTPhYiUTn7Wp6Ojzu2
92Ysrlm0oDr+Tz21eGJidd14RqgXEmIFQdlbJNYGbihWhIAUXEZCJ5+U3j8vTLeVhBlxYHEmuUa6
2AAD77hHJ9ws47wxh9IoBKQTDYNl1qwKBEfr1OosJ8ivmWTkz0BQG4sXAU4t13OnLGPosTukGJQy
xXDCZvCOhaCScer8qKd5HPk5jBcpyfGvd8eTJ6dWXiAG5HAYbRCvLOkoOC7bKGdSuC/GEAb9YGwc
Dr9Jong25OmfmeU0m2Q+M3a/WPOf87rW8ackDTTjdI3fLfIe3jnd9nZlh9duS9qcX8wTpzip9FbN
rUDodGc2CQyuSWCMbrRBhk88UMRjA0m9wG21yjMgg3pHxXA4aitLiGBUhM04wZCOQ+pgy3gKE1I2
PKQ1dvp2Ij+iMwnQKkALTop0RQBDMZQK2AnTSmRBjy4YgaIJ9x2ZN3L+EM5dxetuiqjL2xM8gUqW
P74srdJMWuyCUmqzG1xxVGxCdxW8IgGDcgaL0pc+KYFkmv4PfSr4ySvGoIPr2QeqaKNxtKXHA3Td
6ztbyLMDKrBRhsyYK7ttRi8IAYplHUWCcMbChiUTgyLkAlqC/1hKtWicrXqynWY3PE0gJQWNu0XE
5/leSSGHkn5Sr+4jSk4MwUx0DOMdLnUQ/HrIwGcbdNJz3TzqUztY/aP0rCCabb19Vhp9GyfEg6Fe
kLBYBN5JKGcC7VBR3FnyQoz5mYLEEo+WXBKPfAr0vCSsN0tAqgYrKHcFlOoVJEUgIjlXExzzc0Gz
0fnmuUoa44e+dS6UxfQ7Ab1zUPmbho7t+cqXPWKNOHsn3A4xubGG0yW2MNSfvJeuvn3bK/kOEW1R
/Opn6eCZQPQhli0po+V0hl5NsNqnzMP3VXP/hcKXAFgoFcgCW8kHVkZ8KMy2eoMKVZ88jNFdoI7u
B3JwzdceEeK16ozer3KY9fR4uOkbUV7ikMsLfH1BFyW+V8paH2X8pM/GgpNrwiBz4pVrxH+DlpGM
ntIqTv/2J6EmN8O4NQw8clvt6zVMjh4vvmoQSZIS39HRaPEWfgPh6nEGNHIWrRYUed9UJq73HW9y
jL/BVFAmqOznen9v0MNmZoWi5AKfo+VI067WA6PUcAT8HCbemLZTRZMRNFnnEn0Lu38nusYBt3bK
YlsWKZFXCNmpryMJvBTyihny8o3Newa5SHHdQw5/C9RInuQIlNLD1/coHYVzO/ZSGkHCYB/2dk1h
6KZZfkoDWzfs8Mn3/RJ/XzJDFtNbR4EJRs5rqfPgAdm3bDyYfx7f6lyta6MY+YfbhEapmPU+1gFC
Lcx6xz8n2CGuWqSCiWbqYq4Q50bjYG0lw3YFcOVlXBzFS20E8A8p7twJ1m1pfFtmWHFh3uoJsOB9
2So5E0rJYxxwerWiwNufPpoNYJDU6NqCvB64alECdfqzJWW+RV7DfROmIdtLVhxV4pzATpthM4hk
4U6t7IVPmzsXF6wT4XY93pe+f+FDLkj3mvgCrsnwLGVQj5A9rFympchaZg8OvNHH9XXSrw47MeZ9
ufr8eT/SvIkmmFwjVkQE+wLOzWdkhHnCtmVatu3kB546E9S+TDyMVKyLmdd8NHfKcmimZuMeY6CE
3PDVpeIUD1c82kbkSKcyjuvQFQ7ukTshIdt4Ag+cEo/dM6QF+lxeFQIwJI9WKuhePdRxIeIW73s8
kIvKRWq0+dI59CjZjyulVWOzqZWfaCOix6B8QCHjY/y0mdKGxeCrNHeS+JsBONKXuYW02beKdoup
5tXbPFl1Dt4NVqZEu3zL7rlsP05ktXf3yS8XQ/ocu05949yPCTw+r8OU8mhkeWBoA95c11I/KSOL
C5kqSmODQFJSwCcC/ZTdWqXlkAkjDhi5f6JXb1jsPgnTMpcld7CaDH6tcDnAyDFDb2kipk1/TfZo
YH+UskLos0bnbfS2SaLZ6myZFozVl3E0TLBS+Wo18vg+ViIzU5KEcEQx0lp0F5hTBlmAd/5jxJAA
pnzWzEtDcGS4Fm5eSeMi24deGstN+girY42jH/aQ/4YZGVXdRnxTDMZwKGP9vfQvFyoWK35+9/fh
jRuoWLQbVsRlJBqy/iDJQDdQwHRkKcQZaxb7jMbA2lNUmVXK6ixL04/ZULedtRM10g50X+y/CUeC
S30HD0sBZKhq3qPY4XhpGf4QPKGfZjMvwz2Z+y/Qent9pfpx3Y9JfKqP55Edok1hDwNeEjNCC5mG
xZkuHUMhdvRY7bcYvjgbRC79ylWDt9Fi4KzU//iTZhnXOoEYG5ttNJmaPHCAcuoS51CfIEyPa/bb
652si5yDqqOvL3qD8FLU+afT0LUksZaAjPNXHg5HRu1mlSH379pn9HYo43NCLorqIfg4wFpP6Wbh
h9JQI0N/CwJ0Zl3GoDYDFvlIMbrEGZnq4AaAVcUuSj/2P5I5DjMpF8Y/S9GokHlsOeX8i6IefWDi
VHcmBOdCX07DCKqz0ziJ9dcbVLJQCZV1x84dysH0sOW/ikVY562mWyZArMVQvJdmEq78PXGhAn1M
8HNI/gmla3/J3SncOKmoSIIlt/3TBS7LWlWXFwI2o64pt6Ak7IpiPq/0+qja0VFc3HEvFpudfadk
IghYZb63zHaVWP3wI6kozFClaRee2fbQ2LyFTLC4cJ1rt3lLA0/DbwXyMkCxC9+7IpM7iitnBtKR
pPu5FbmCONynqbRudFR1XW82OlMXcB9yU7Vjj9Cei9Q3JFR3vzPNphMbQepiS2ToRa63ZbmFO427
vehL/mlak8lS8nPt6YwqvJdKdPA8yzxGtGdxtDfeh82z8fmEAPw3EVsUbgBjvyFb57g28D4eVWyY
7y3QI9EvQmPgfR9RLn90yJF+1cte8HgJBfs3hYzcXA50YSh3boNq8vnDm5Z8XpYmg5cbLFVq+u9n
Ovp9AVHN+bVk+fIaVQM24HaYY3ITJePMiC7WAGxHg+wb6RiMlEslDg75WBDDDSwTmvAtnUZ+xp/W
Qnog0Xqgzgu0s8JpAIbP/+anVDISoRGHZkJhlbTVV4jtZqfdg7SmkkqPLB/ftxk1MASFzrDP/6uY
+zuaNiIaHTupr7FqPNbV9WsOV1usWZpe4PMqUPliXiCAZ36VDpc1YY9pwU6PSFHaL5t72pfiLJ/D
HKNnnCCWqrjv/DGFWoVZiPuW+nbLqJnTIwryrNEpsw96HGqucqQPXJBevR8kApAU5EKfjEAMMVsP
h8MKpkURboSR8uKAdyuy11qRoWtMTmmHTICMDyKE+71OCfQ2LV4F8Mo0/hEjsP1rr+sdo8ug29G6
6lqdrT7cA5H4OulUV20GRukbkQ9E2wAOAcDq4ylzZUO76eKY5drPGokfzFdIGqmIwzbU7TP3998L
cUl2uSULo3f4wM6XAUci7zPQh+ARYlG1u9LuNiyehM0dOU/Ci82WWjwcsqiyGxIYuzeU40bKrX63
Y6DWqvTxAnsWRtvDUX2YWZR6Z1eB8EcW15jj2NAZLwOjc140m1751Hl4ek3hVpEPaLZ2Z0LhN4iK
S7jc1GB+SfaU/otTAenUqrUYjbMO/FmGvfeXKAsgBRSGqmmWTlNfU4tSGiWlz7wG5abT+OOkBaIC
9ksYOygqTR2A6/cTIkEgT4VX8Ug1r2o5O/8owol776SN9lVmjwqlm+ztLTjoMo/prOwwscV46IiX
dsQkrKSo5jDXmib/2l5gYrVlzetLvb8ABwuW/IF2y4LXB8iYeX3syd9dqG0wm2UR7pNefP7TQq+q
qnxFLkEHgPMawY32Iln08xO12PWYY0T2azGmp0ehrQgGa+MhrC2Ju0y3btn4ozH9jnFFixsIuI4K
6MWwlbOLSsVoygmUjWjafT3gQsRt82ZlV0a4EtiAcYDhRCtba01JhzFsz2rKmx4XYfNGe2FxmbXn
NC6zp8h5rWf/OdUekAcmpdSRm8DmNBPJopuLPUSij9fc6PloZyVoY6ak4GQ8w3X1l7z1ZpBYuSlN
guZnyv4LwjJQaYgstt9WYyBum1CXaExmB89w5UOok+88cQTA7dx+Ny7btikHkfRcpZoD6iOZZUUT
15rkZpikMAb2HfHBMenEtQYABToMhEKnhTX4gcpg6IbQcFHtHaJe6WUvJ2nS5kT5uisIkmFnO8fG
jOt5vQQWXRtPVa4IqfKR7FFfjTwIyyc9tXZY8iI1M+GfuzodVG0dW5LUmoDLLI2A07d3Jl/hzDfQ
gnwFT71C4a8JMBHKglP8CHXjpbyMu02N/eWCNfZks3lx3Tz1hxRgTXwGafYk4Xhgnj/H66T3aKCx
po75/scE+EPjbKzk3mQhj2aiZdo0a6mX1NpLiWJRU22pxtPkDWYDJf5RffV8oLMRrMimftwFsik8
u9ljGZA2B6VwTACKTxc48EuYfzVewnl+QpUWhxDxAi9P9zCdwBnBtk7AB6DwjBEBb8e5MzzVSc0C
pB7FRIHH9Ln3/c2DQlAkyrrbleDS2qAj8dKBdWFLQA0cGUU/JAsrglZECXWeWZVrLuJ/0iwjPmQg
+MgVLX+9arZlYLJ3FEwmgpFhnmsYpc1LYCMo4n11T7KkVvAOjacLxk9UJBOBZpvWCoHOaimP08Ky
W4wzYz2WzmquwlSpS2DnOcjiDY5a2IOH/9YAgprnN0N8j3U3PtV+/Hr7gCmQKOx/tDIuXmkmVaHA
bqA/rofNR+obppi2SuNs8gh43FaGUz6SktJuJwiq0iMJpv25B1uqsUmlN2j2efjpPZzAbkk1Aks9
Y26Vj6tQ27oyaeVOtA5dIwy7yUftGovWd/h7n6c3P8spaU0W2IpO5t0EXy8dd4aSCPGMy79h7ES2
neQAwkouD0/j9bbcM3NgdFkf36DHxlMgFb3SYm7ZLhAahzUjIfoyXqHS4el0iPKhz8trwGLKVMvT
zvofJ02Jt1kLtusF2k2OT3dOpITdqk8jiJq47I26vEgc9RH7ZicKtVh5YIdZePGrzraWIUY4PhBa
hrfr8FxOD8WbcBOGuL2G3wLUNs7Fjim6y23xFHibGRFkuKeoikNaNfaGeRv6E1KAEp6Df4AdwSbB
pfBQrJ/P+JnW9eMn8wO+PKkOfS5L7bdZGJQZK4advddyWPwkXFsrB9GmmXha9Z4OjnmxJx4A45lT
zNYLNuKREg0GX9VvtUpTaNF96DAAnZWPEO6SAJ0ZGAtYqcZbY47qGh0eOh/NKqrXhOQdcUTvWrrq
kgsPANXkG3PAdMnyhpxpxbZnCdn9VUF5R4NL/Vqs28k+CiRlUZyruQAxPIFMUt6ap54bg+YwrLIR
LuE/TVkUtzwUN77F48+kg5NEjef71dHKfr/0B1Q09iJhb5RQt3+9G5kvpU7YS4OCm6hm2QwbOjjn
3BIdw8rCkk/kFtKsm9EehAE7k/jk29EorFCMfoTDahXHKkFuiHNUH/B1ejcjOS5UHFkzWak24NV/
qkQHyef8BtabwV2oSE8BGNDOWVRffpruoGaRZJj50dXvVZEatBloYY6MI+jHTNNatLCD4T0uKGtC
KpBJ6lRxcQY/FdjD6W/Dy+sbfnKRCsc8PV4a0QYyJ6Hqm4PpGV/hkakTK6EgkfHeopW2hhfV+RSD
YcD/oU6yKP0dg12kmVopCh1X/LFoPblscfBs7qndX8ZWqjT5BVSiZ1QdjBqEMFhp3Hlp+isOTVuc
viOsT4lT7yt1fPZ+kvzQPfmm40dvcTngSmiHa/8dRnuXIX/kaBnORTRAB5jod9U4eOD+6mFXw/OI
OQzmoP0jgLs5npm1F4KoLHFb5Td6rZqPLCJq6aHcwu76YXWnSrvXF9Ig10x+5cZGILFTWopqL8Ax
znIJyeiXbIoQBvKxbvKqSoWU13nHQmwMKXJ23WiGmB83q3LinP5KkmdZZuT5aryLLVxnfhH4fZCE
2zvb4OpCr7vQWl7rh7kwmJS/VZjq/hlDLm0b6NlhGDGI/WB4APxg9lzdkyLZeiRWcEuTWpGha2cQ
0X7TCD3GG+SwRJfOIadDcN6l2Fq+wiE04SLTC4U6MWIL0HW8yDzxKoWLZmKVc6weSxvymVT5MKX0
tzOQcdiyu/ZrbfHlqHxcDznO6jCBAfJbbBggKWAxZ0hw16jepqgTEqeieFZgZPzdsbZlesPEc9IZ
5E20FO5h36NdEpKqQxlE2ekq1SfCQRfjn+Tb26hygSFX/IwcI8roET1rAh4jYITpnTwZdd+AeShT
4wFZ//HHDOYQT6NJ7KIK8GXNdCYIQko4bcaA8dz4wMQTCcQP2VxaqeCdh2Nii+/jLb/5a7JWTkRO
2V6CalZL/peFyGKV352JMNccdQx++gk+xhJCXQW0CA8XLIVKi1saMRwGf8jTT56JWAOd2O7D6Wq0
l1jILVtvI9bPdlwPx1zH/TvC2J6+elD8IT16k/QKsOIT0b6q+kCB+fx6e0xlJX1fnI/mhYpK8Lzr
yABLfNL/5MSHlyrw1bI3EiKtmdCFUBu9KIv6gsQfScb+wxiGZ1xqyu60cWor0E/gto61sWZ16Ozi
EawsgDr4BnJMhApKTAcvmlztZimzkW0Q49TcpagyT4H9FlhlGs31MQq5JicKeatFQII6CgSrlNVz
0/TOjaeR4x+rEJeN4McZqiDFIjyuYbrazfBoseLV1tIbi1wVg/rHp4glg52GsiYC0vGgGMUu7MKi
83jECEwkbPC4SBEJl23RS7G5ru7hUM2acDOUoiOyjhF/LkzGyjbdmR9gonXU4dEf2e5c/XMVHS1f
bQI7bb0MnZf0jECrFvdqhsh3tZEiowmrSF5Sj42o1iucT0AkPwpazKruieNpWdFZSvlHXET6EVwG
RgdgyfHsYpi5TszfBd4WIPc1TB0xlmrmDKyzEcdxAyUxl3r0fCyrWIPFuqemB+bGvBX6QU/hIbUY
gWJQQtAa3eUaKAKv7+No3rEeush21UsNaTnLrT2d/ql1ecsM70d2fgRuIGoDrJyUfU3fl4y5yPcA
NZGTd66i36AjjO5MIg350bP/skL1K+x3opQjPnXzkVkrFEH/sxqNgY1mP8DTaS8k2V0Fa9hC+FD2
bgbZ/sJLYayqiwJYCBHpU/DfEH68aFCgHW/FbyzDLSkgDMavvP0A5bco0dP8lWGGgqFAebitUOcZ
9yLoS3SbkEw6j+whGc1nf5xaryMrTpKoWGVC8Lg59tI/PwOCbarZOKCBnboPqLEjwdfV4QYHsTc2
S0sydU4fHjRCL9I7gJMob1RD6iPRDf94g5nSiPjAwQ5gTZUD4r7vdEO8R8Kduy607c2HzbsHxBOq
Wd2UobWO/1sNAtQUJFAjeKvxfrCwmzWvCcIr+dOkYoMjytTznvvWnSEt95PrvyCLwP9HEzrNsZ63
Li9kModvq6IE7Gtf2vmtOLRVnuYUYiHK+DMOnO90QSuwkw7zuxMnr6cTOdWVaPgNuDguHwSzH8Nq
1/E1POEHr1wn+K5fqFtiJUS0CBr7i4muWnJJ4hf5ntKR/z5TzKONMUe16HH5CXpajtjiPMvmQ9dM
9cFXvXdQz414MWC3vkHIfj/tB/6tnWqZx5SK8IwjIaNH9kEFoLH3GTeMo9/+g9HgS2IsSUBenGBD
fEKh5FsHHWlb7i9NFTXgxBTJZydmyW5OZOr1vRFOoh7ljUBHNAjHbD3StVB439xZRRhwdbwkzjyd
/pLFAOP12HNVaAtP0j0WJ0XeJ4TI1S6KxIjpsNdIsWQtJsbIXNqnXiXhB0HFYlmonMH26TwEnXq/
DQHdnBHBQnKOsxE893fsg9K8Mwvq79NTvjPuLy+pln0MgoANv1HkN2E96IYxG+E5GyevDmG31psL
vYQ+rTVy1pzzHjrSK3MgZ152q0le5rPI1+EzRC+kJBeZyXIBB1MyOmzhgo+17wDZT3rlX9xf5VlZ
vwy8+sRGgu+VcAMbWgl2vnWpOCIT22F5Efi+O2LNdalzqVan3C4BOl8zK4DeTX6wCK6fE/tNR0kS
L32Prsr593Rir0vtUZqgHuJDndWAG7kYojLAmjrFn4W8FWrEQB3fjopJgu75CYSeS609vu4h0axH
lol+WoNdwIzMSYVxToA55X6D28KtMdVdV2/jcFyrkfeLVp8BViCda/TCOm4c2gah9Rpj+iKddbzy
bjNG7KYJ5DdMEOoKSpvOubIRKkyvzSCBGmLqpGt6ru1pYkHv28gkL0DInKDP2lMR9eeqpQ9bKeZH
lTbOCvp59JEL0QgDdgx3NO067l59j6zBE3aCYFgBavWlruYpXbK13iQ5wcXEK26fUHMPJHM7IYcl
+F0Qt8OlOfKkc2LGiN3sgATBDDaAFOB2zliz11MsfjE4jRmUn1lmY89sHJVk08Wj/olRHe3InVww
6SetV2/fvzmIXRMCQjZamvwbyJMGNYuR2Cczo5nlShXocl9MoGHTvVCi9VtoGI/AzuYIMnp6kr6k
GcsUXK67RaWBGB6I3vuml4nplJgFVq6GhBeA4zmAHN9Nyiu4tqpOqiyyBDIIB/B5LttLZUzaiPa+
4ofcbo/1vkzpVYQYHTlbUjbhDyIlG8HgnzigcbCd85FQC0gpK8C9i60EDb827juT49ZvFYlKXLPx
A2wR3D6oRTGPI6EC6WksteJKJ742z7SDW+Lx+cPtvJVgzIpx1U+v04A3Nie4Sr1YT58QCPQzwXEe
DvM5TsoWtuMSH3hgYs+cqfistosmpcdNvzh+dGBK7pQS6gyF+/nkIpGb24m0v+O+WbjHbXXgeuw1
F6oWJeY+vCW5PXxTuqtvLyTPcmLRAF1UYIod4aJvYc3kK0SR1Zrnhp95aaIyES4x01jOLMR2Gymo
ELyOh19NcbmhDgTYcabwINbv7lSxrVX2C3PSf9ibSmeWGhnEaBeQ8PN4IwqZ37IKkJmnXXw9BqWZ
YUBlPKHNAlxgfnQJlk8cOg7g61el84BeBCQA9Y1+bDKw/AxUfmrolbYZIN4++458O86/CY1A2LY+
I7urtm5MmEhdOkHhcaeUA25xOYEb3FmZgfzDFPqB6YS6yMYIPzG6Hb39MsUGFZadd2Pz7FzBMTT7
sw2GPWTAGj1AwdSLOKtb+fu7ulp3j4SRJjJ7leiBvMsjD0av0FOvZBenb3fPSwjHi0sO4t7Z7qo6
B0fjR/xdeRg/yzSagdbDRBUTY/5o3NKTL85aGNEFBq7czocoXYZ51WKr0l6dBsnFKCb4JhpSUtgk
9/j2OhEjViaQpFbXmyIqqTrNfvfXHJpSwSozBrIGpLt9E+IaLXLwIG/9FUbjmQGlmWpJzIABYLif
Zstb27Bym0gme4Rg5zj9Paj4NUGLAf09pVs6oxsrNCg0YEj1bJ1cDPHFpEHZid4UIZO3WfrQ0fUa
/xiQBjBQRSCPodY03t76aXBY2YBDoid+IlgG4r69NY4XUh09b6bIfpBlMfDo2o1IPcNKtayuO9Xh
2E5e2o7x9EzmBg1clHjD6Yx7uDhzjhr6RyS5o9vsB4wYzj8+mdekkTsFSUA4eRSZpLnQ7gePgMy+
j3qcOCk1LmGAUMb8Ev0Psqxzlj3wzyXm5hSVTeoU5bePq34Na4MUnLQ0Q9zFvjuep6dhhTCbRoeV
uOLvQzuObIsOZt0pvWVnfN433kQlS3HDEf/AZVRfTYU9QUlPMAoc0cbsHSJy1zWWvMUxRghQohBD
nlk1tDqvJd99TMTYhr9zJyJdzoYFv4eEasYR+4WiX63/3qT2qjOr9EzyF0YO/yEUg6oAonkgeoKo
S9A71B1+JC0qZ6CakhVe4eqru2dVBW7wsNzUSA8vp/tqLymOpQi/vY48My3zPVzgg32nDKhtmTCw
hd0xofMo2ZcSoY0ux+ETm5AUaXOqO1ZDkhSdoNdsuHNs+M2npeGqQ968UHXWpjxxSI6Um5cQ7gvc
OFuJ8WHeDSzBLWV3RlPT6OiCYK1rZpi1wSLLBTYHRB7K1rFhDx2UaNrUJun6zZqaZ8aZiVPgeLCO
SXG6h3K4Q6FZWRiUXn5qjo4t2IDyEqcDk7cERJDorzwXfjQecp1GBb2ax++1JugD6JIWJ1yVb0Cq
pYS/LG7enpE2loAHW2/3me5ZJl5zNH18l1cOrtimRDt9rGV3FRDrIRD6jQRv/fH4R2QypEvxSmhW
02DaLFlzxJEKHhSz10sIgi1KPSg+Hv6BsKzBFr0X3hf8dc0jXVhtBcKt7/FuY4DU+WkbOCT2BGda
ktt028s7ePJ5GtlIKs+pHmRzHRLcAvpPEyYppoEdabhLp34YxNQPHdBMXG3hVov/LWnRAi8bhg9b
Z5kyQJ3QYqkmwIbniTIv7/N0g1WviaCQ2rGwKeGfEphuUH4pQpwlk9AIcL9Lj9tCcoR1PgtdbchD
tlt+4Kd35hp383XkvDz9usKYo5mDg0wLEV3GSyNC6cVo96CUzuifpjAxe8xapqLwL+zjrq6HmZXA
/BAC8pQipnq8XW06PbefgGkyg0NoVJVDZ1nsfm5DQ6hWBy2vzLUkX0qxmX73gdQyM1gphlTzqti6
VbKL2dHa5lR8AwiAC5kxF9g1xu/yao1ESlCqdQJnzayHZ9bzRFZV8FvurzDllEFopEMq4J3EFmGS
7UhHrLB4Ub552VHq80ZRmT1PCytvdfPDqNXw0iBXnK0do7+iI46Z2KhMXSVniWyd+lDjFRCGqrjU
lFHqqOJrZ/e22JtEU7uYSgWTM2g4N0yL/pLzFdWDvMRinD5AkaM3cjVIvlFnnCMTHtKCWwFZBwgJ
aVQwBcaCSITXA5qIUbS5xcGS1FhEoPzcbDxf8DalJmP9VpzPFs5YPDfnH8hlDIqixQMnOGVHRyqD
r/dqXMr4Oe300uPo57F7xKsAuS5KmpQW0E+Dz4QqjJPe+g6cYzhsFA+7BaXnBSCmYY99ad48wPK0
Z91QqGep2Vhj78gKYA+wg2f2dxy6XVp0YFJZiQyX349tAtpew3Svv7QSANW2xMDgqDbdVj9G43W8
OlIJMy8quf6kWhm1lsv4nuPs/BaxScY+fCrTO8d0rZOJpd3E+HQjHwEi+E83HN4ayRyQU+w/knd6
JHN5UnEyCo8cU5RzA5auyfV2qqf6vtVgIvTLxcClViYCiRhSRYMjWybZJiVMpNwAaE55QnY33Zz5
N0nc66S+eYV6axeG5B+kD5S50Foo8pqceQNxvBow0U+snhAFlnf3sJxVDYSgjTwJO6gIPEN1+s/q
abtFi/HaWizGNo4TPPX+/8vauF9K3CW4sSMiWphP+SLZMTlfeYZ1InxGZCsjr8eKzA+nzfYV35y4
u3UUnIOJbAhq/meP29uw0BWFr1B2CtqyPOZ1fFipsvkm+1TErhzyReSsuMebGYP8bPwN7A//yNAA
Vo6p3dc/4J1Ah8R4Ka3mAUEoID2NlZEin1+tvMe7INxWjpzAX1+TYSCkxDP9mAjFQFfjQG9SnfzK
M7WYJJZPPkMEFam+VqzIKo4CKZrMmWxGYvg7qrIyzMM1SJv25b/CcWzmwR2wuGvYtVmbpoC6+lTO
z9Cwy3SU5yBY4P6pGwrf1Cee2Mgk8wIbxmoDjZGV3jxZd/+/DYA2H4dH83VZTkL8j2cCajYST2Ow
bAYCFkRGiU0CTcErKEup9YMqMc0WYLCk7RA7YIE2EVx1icmsOyc/rM+bkJK+3nbZ8xLLc28pPI+I
HhJNrzxWoQyTZRIYKpIE6nt+gFaWAUVipFGPvpC7W6XtzwAAmOZPUXGhfWP1wHl7t1ieSq/ZnwPe
enAz7yTwYYT6nKdWSaDciukovopxLWNKr+EE/YZzoqlALrtFHmwfXZ8nYcXHaw+UdMqN6Imsd0CX
xI1RxtaBcb+1rqO1nHaoXz1qXqJJxSXkjQnsh2fztq3d5WaVe+wn68Tp/3gXg4bX+jB4wNee6dvG
+lIJbJpaGp5MexARP+dKlsapE7LAwpC1kJJusTu/2bGr9sC09qCA8EbQk0ygDhRPndwWwpdmm4bm
n9YFwMDj6Lgqx7fsdOlduT2CyTbnc6C/KqupZ41VBbG7rkHtNSZvFofFq8eccaSVytAH5HproDfJ
xf/HfkuBSccmyXqdwguhSTjHtv8OyRbNN4J2QiXZkgQr0ohCKRCri+3D/D3u2QioLb/gxwXYsiEk
Fzugv77BV6MEnHSKjKVEm0IVPAwHJ3zxGNwmH4p31B5blL+0EhRkvwvzILQ+oCBwO75xGzXmHVqS
xsZDxhsetjvaYoPtvTrbo/nj5ktPqSoRIqk54lfTjIs71CKEPZqyqQ6A/ur6M0OOnJiNQbz//fHR
0GubWasluK+/nJyXODMnEWrHFRnoKlCs/KZEP6/bxFntJWqcZm2EdQk21KVCsv9VB+Nj0n/fxUvf
oPa6DunGHh6VDBnU1Gx8zp/SwTnrnrFFURlQwob3BLEVofrSRGsz6kMUu3b/8exFq7Rhjob6GhnK
r3517mpxDvyvpz6kQQGRTZ4VyqbCETzE5Sv2MjpYfeuDef/OfjhkIQX5DaleblhV4f7N0e+/URbt
T7Ii+ukSKu9Aa7pP7xdOySC1dPHuI3NRHg9tIGVjEq6hZJ6Bie44T5+XPdqWbU2EDQul/5MUWvMA
W5M+mO8iLPUbM8Uc1ONXRv7Qml28H/BgQPSBJRw0hIVq+Ts/LR87ZyeGFk41zLCVu62wRegYIa60
yC7Ddbd9veHjE+Jy/JnYIS7p3XfvtMGtBSnUqrIOlq19zfeEkSJDc27tphOk7uimcVc99bAq4Lb0
dpE5T3D/C88AW6506PINSCaeVOoIJO2v2aYfw5I12YOGBdXB1eXWIkcNUp0nRj6tAGzlp5EkAr5F
QAOX7ca2lcrhhx2l/U1Ht3b7dzAozRqL02quoFy5fzgtYAok8WLRMBZsNBB8LzI4pZev3JCrKfmS
szsROg+6jib6VdvMkpsX93I2xvXzYVvlLZ2oLnUnMgfA203P7rrWMx+k/6Q7AHATGq9oIH/nZpx8
qMoUWKRjvFL/u2lgHVuVjXiCZzDTqJcWz1luaEj6PSA7Bb76px6I7nHPw4fSdXxBrn4fEKoUQ944
Ut3cu20J2FzfIlhh3g4po003U42KxtTiu0E3KZa5TicN2ZE7up3c0vACUHTDegjDpCYVr+qs7dp+
vHuxRvfhBLGkZzWOws0ZQ9/lyX+R9h63Tvd9zWDSKIrJI5vdxYWgngJbJbXGQPuiSuocqF5P2Itu
HXRR2bQ1BiVKgcoko0QmqLt7GsKsMld2oSuX5rwQxEjwN3XmXz2Yiwd/SLriHVW2SJITUhh/oXag
pIANod+vQW9GCzeJJ+sqwcOpbTrXtFQiHf8BOMkmte/X0gRxRzj/Uru26lXl8qoMigUSAtm7aRcQ
cddmwQb2KhuVgWbm9T/daDuZoaIWEpWWQOdogc3p41My4AeIKRbdAzxBFdQJK6+qKESerwCfko6d
etYox/F6/RcK5Sw1zWFYcbtpe2SwmDPXhwrHZGr1q6Ef/MPTNclo6KytqiYb3BUQ7QgeypfkNjk+
EdbNLo/mUaYelaKoAbc0kAdfgplz+uL17BxXtICSx24LCONUsTt+uZXYFDu5XCMabkyqGwiNvVFb
v+Qp7WXUQ8VrSEYIGaug2UX9PSeAkn7/G7Njgt92KI9cLAhrIasAXsrQbg69S7obaCdEhw2Bny4P
a9bYTx7etR9692HSiYCP1FoLVf+ahqMdMWdeL8oR6Fkq8NMOjyBzDQ66dMyQ2hb5NMbHhe0pt41L
D6ZaxdWABXnPAxnLFuhGn33lgujG7tUmXbhsqzJGRwqVfELLrlIH5bsXZsOETbNzBNwRz9SmbXuy
pfzjk6IejQuNXU0LjBIYQPsuwkrVS2Z5eHGYBQ92LwwYcNkmpeg+mMa10M3VzlKorzhosiTbRKIX
vCtQnCCpkevedyTJ5RiZ/aSLi0JzNYX6JDm84rKnFli60sapl7E7Ub+xW+VCOB+73M5a8Pu8xBD4
naahcutb0IL/zVg0L/RrdrJxOTbR6MuakiBzOG5tg9HHetcQY7Jixx4/OhDWpIkGMnTuZZ1GVDSC
z70y6+DdOoyewIpzidxmqFURrGnLxVVssPNQBh++lpPZmHwqIk5+Fxn68ZK4wHXFmMIfX96mYgqf
/MwNgENHvVNd36g2f/cVTCgf0+jt6VPSJNP515/dCOF+WoZeQAq/cvpFANdnPmNNmJgWkAj2qCWc
chMu4f6h+k4ZZt88TCKCdZyuEEYc/POobpkcKt1281K9XjbaGmS6hlRVkCsvI1CvU64QK6I48vT5
7t2T978QXj73tedvsuBGJlEyNkgUNOuxVBCyia/dQ1ET94gPjiOq+ZClklA7tPeqLZ0UrTDg4mS0
43cx8nXpQ7kas1egyMsCEilq0p9M5uGTIub/J6r3TYW5YXAuK4GN8EJxiXzrvu4NcSuNt0ROcRnU
tKvjT9aMJg33SLjv9imGYXuD3zxx6qQrUdBsefr9Bkp5dC6aw7Q6ojYqVCvH0em+/E/u3MgTJcXj
Is1lXlCpC28AKE809gbSHQId6rczAR/3KBCLKvsKOUlHrL15j7+Zuzt5h67B3UETbnQz344Wt+mz
mYxE24GLm1NkY+ZiJtc145upd39XvIBDQg4gZx8+NLBrQtW2F921EutzHo1o5F3mlH1iD2ecnxME
981Kr+SkAoN9j0NHsMOOUlh0kxDFweiCwZyU8M/tjacLNueBse9IAEfnfvDGKdHu/WGjRtnxjsRu
DMn3CzsawaqgaLIe67fMfDUhObBA4d0Vw+URbr6Cnb81fhjl8FNqeyR3+XZ1FdIEXMzh0GALbJCb
Ye4oVAyLEQ10VS5V0mkzNEIpol7k48noPDLalGSOypd/CqgXPxDLEzA3k80VxVWRQhrtf2JXfk6v
BJDXMMWcUpl2ph4NOdUC/W/oN0n9BzVhqTt8UnTmHivWGpiUQsVa3DtLW+Lqy5l756kQ3rJsYb3c
IbvZCrNgHKP+ZQxeAtn3xNRnawQXxJE/oqVA6sngNcooQVt0szV/UTIHPZAImItFzvtmsWM8Y7mf
DMdIBoOen/0lCIAmcg9Wrrh0rv1X2IkwSGdGyYXxkGUjDz8nU+QIqvuBa1NoHL8lpAcrLWCIInb4
xOFexdN1xQu1Juh3dT7qvILuC6wH5FCF0nCiedh+PkMo6EkQFJ2AGakpyafvEQ3pmpRdaQZxi2/7
mqaYPmDnGhV3TKPCUHCrUMTuxv/d+1lIqUrQNe8Yv6aFG1gWzU83Ce095fvawuiScCsbSpsFNXWc
chFhX7D7zoRrrgDAUz1k+Ha94kICpj9dcYz6LvkvB/PU9z8sEof2yWDB7bZrGdYReETvjIliKfZq
kF3lfcPWO3NwcGHS8OL/hAdjhbztXuAUZz5ma+gaY0q6VwTjpbqaKuW5J+l77ixDDnlxvYRAo6JG
6CNjr1bl1dsOYfvJw5bTQSZ+lCWmwe6KMB3GpRzLg+aVXHtIznxJxrmyrbu0lFb7MOlF1XsOb3AL
As6Y+2OMe/7SXEagXHo8CJju3olh7ymDWHThpREi+Kt9M3zlpYhPdRTlmLtgzo+Bx/sEwpPTCQaw
z2Oc+LQAygnkDVOyunnfwaWdFF+GWFeD3aBOc8N2ZZrqLPc4LoOrnVEe0Qf35sm8po67eso/cG8O
78oM80l5BchJ4hds8ZGNV29qT8MjxG7pVqIfwQlCu5LzE9JFAaTGf6itgkgmyoqclJQAbrBZmSle
EbK7CzYiLiDICL3bui4j5N/Qe7jn7mvYrrGNlDboDP53e+TeiimgoHNh2RGV+ZuQkJsUNykb7c9k
jEe5y1CIRCu3mVHr5rFVYS6pEfx9hvcX30KV6qrFLyhtAtpPEzHwv4zUcohne5XV5iC2Tgzhw5y4
yhAHmVBt+ZeRzeolnQjl++4IVpmZvakKeAAQ5iY4C6iPUiBAdTSizGGTZ7akHaUtjJKxrCzOiY7A
jLeSIJdBjJ5sXg9rXDU2sDrEzyixYvA1st506T8UozrfgDqOP4mKQCscBduyfb+fmS+XihayjjxD
D3dHAqSRfGKIbcS/OpaHUMaXXcJUqHLI/04px5FjtfnlLJcZTnNWqia7AoSikeySduEbJX/XUYq0
Y5N6th6W9GRgia1aCXQ4M6Ct7Pn2KLteq83ThQHCEWsuKgc9JjNK4OFXen0j1+kSCVwA0jrcMBQK
rFOduttFZLiW1bVchFqOWoos60im9SzrXKpYm7BUjOf2C6DFvw2Y7JKpAKy29mw5hBJBWMycNSTh
xgzvAkG0GHTtNkte/bp5ZDsGeZchAyHMQD9N5+9KsShD+0L1+/WCRykU9BzMAME8K+5iAFydkJpZ
0NfOrFBlmG+A2Ccs4smW2sOzEybrIjzyRCmv0kBPNGDGTmgcFJKxqwH234TBuS2u430Zof2T9ok3
S/mVBgUIa51UlRVkVYvV2NOQ3G62RUYteVx95iNO2zrj+jbwoWdPOyUFrRBXVhNiYfk5puL2MgEo
y9ldSVywDFp+bg1rHlK7W0y6UaBS1sAFAH9ucn/XjqfbuoNmt4f9w6ZozfJDLDBeS4qK1cZ3UAB0
suheNUQRuaZ/VoMMECrdvhc0Hducdi9jlObHpwtRajDl51YSa3Pp8bkxxsHv2kQdY0iySZKVrr5w
QMG03QSDHFECY8WyzBPlAPl1JY1tANHD+eP9WM7vkJ2y4NVknoHji9P6NSlmQwnFbS/r2T3vltjL
kuDpDeBrvGB7sWs4ZoHJpf5CwSKHU8PrlPk09zaO+fae1q32O7csuirS1INeT6Fl9Pqo9s3rK8La
FSo2CTGNB87cKl4yhWe5oHRaEHVnfzwMbvAlIJ26VCSDEOIWx6I6pHZvJmSuGF9EWo/Jy3pNQuk3
Z8OspB5MZsyskcbmQLjgOiw4TB7C3jNoaJWPR3m0Vqh/mP3Bey/vNejFjhFJwySTdDZgMojVjrKb
xwPdEM2N3r7GYAbR3EFiy7qR+6oywv/kOIYZ9LhDxmphJ3fgQrptTiQu9po+hkoFqeyxqqaL5euS
oI1diI+MmDUzrvjdxTMakB+9PBlX1R3Jp1KdJ/ZNHq0sHQRVs6nlunYeqR8vkuIUhgISvXMpS9Gc
qf+M8TBig52gZcakPC3af0NgvaJ7C+vKTm9YunocZwZMuWcYBGF10aop/NR5cFDtX7Eic+4FxWsj
UYu+TpnbPsw0Uo+9WXCgkK9BrIXjQ1nJIYdC0ydYpXsCEann6RRhiK5hxKMGs31WjRTQAVNUI8rY
YjKqhZPbOAJClqbruVA/HSskzeSAraFK4CNzIbY0+JoqAA7kB6g0fevz8AvRAJMSq+GMyUVr/9CE
tByw6Ul7yqIitcien5l2I9yIRX17mN49AFfAgt8JkwFEYVUbnPX1989bZFwUclY2msLrX+IU7mYa
j7O6oUQicwpwxnHrO6eeafMwPngjfpLJVSSLfx/RKSuQcua6Kj5EnttRFw2li0btAsMe/fZ26ttJ
bFqn+MX7QJuGinK27+U4RLWPo1rabamwSOH2EHtOqALmCYQc78x39B4MQOvD6c44++YzbPO6qLr3
ZplhM30gP/fSeVhM+GTr2UEMC66wfebOMXS1rrmd0hPC4xl4XnUjhb4zZeg9j2DP7qBI7Xdch/iP
O3ajyccjekFC/P5km0UWKMWVUwQcdySk+JO9hhwCzGnZFeKk0eJ1IwCe2Z6ofFdUXXHByr5gpP5m
NFb4NtxfygJYm8MXmwKlEE58B6Q8SCVW6aNqRc8WxribOvdjVlJvUpZCJTNWOI1QqzId6LVB7Lpa
/ieA5nNDeTPLMQApyuZmJVM1KPq7rnMNTYOqa3TTHKdNfETrdJd+++tFH03KQgltbqVuv/baobC5
XwHbfqwEPYr+iZEDCrWoWPMnAveXM1+7CalTjlTnd7qpNQg/Phk7Yx0fqrLI0TiPWXcpFt3mV1Hv
VBG+4Z9hKU0jj5yQFScct6AltnHDqMUFqEH46Bh/vmRNhexXhNcUchgVHFsnnjhpy7hDC0HI6T0a
VLPbZPch6d00jnWb/PeSR+PgyXvP53+sZOxNQsgcSmstEKIkUqCPKzzAImwAzxMFmEPAgOQ5IIGA
o5AaKyz2HWzwP1yqJSojWWnBLaseDujVstPlzQShjTvqszl8LNvh7r5I8jM96oQwNz2SlrnCxLH8
KP5TlrNLp+tveunQSLM/ngUx/FqyXqgpkgeiIYVkpA63kMhS5VVWdoHThryQsphQN5meauuexYya
Kyyct4hfS1fQ9xEzmU09jNFLA9xLZCzBFIm70tUZl0Ji4GT/hHXT4jgsRg6Mmjeok5nOV2U85wcF
EQYezfHvANXsq39ca7bjp/dvyKSfHbBAp1Fm/V+SpTSFAZWSBeG7FMbX9+nSiki+PkhQSPl+X25i
DDNQsFu4DsKsv2ZWapd+NRoBK8gOfKJGhT5dIldAcawFM9JxuSqhflyu5F41xis9WxITSpPf0nh0
+gEmYbaKaz3BF0sGct/kBK5pl//UtuUgIXpYQeO/TJpTZCzvEI6il3tsM2y+WD5eylxcYO48CpWO
y8DQmcVUqsziHuiEyp6ldFR5Hrsxf6HO7yaWkWOzZDdJc32glMwBwAIyoliA/ij3Rayh3NEbXjCI
6tEjRcckPj3kOvh5ml74w3/IoMfJh1y/0KV6h+wNr7rhneG/3tfc1x5cjOCmvrlcJTb8W/KbS+Py
jQgFHq7kGy1Nv9sADh0e6BUaM+pDOiPkCxxnYFt2x6CcHBN17TiWqQNq8OXhcFnbjQJHcsiO5gMu
51nSRXoPVQS5IrlMoFTD+RRYpC2KYfNtaCSg3wh0aIHf6vd84bGIF4K++KzAs8jDN/njeOi9VDN+
oSs62r9lDIio04FuqWvyKu84MM2ZGY1icWFXn92Vhd9twbOMLGsxlLjzRDpct/Ka798qmVwMg3bB
uHu4LsRbT+lYEj/HTwkZNxETsWee8NggNsdDFtq3ByXaKCPNZ0JyY6w3edWQkRol0oDYg9SaYXRW
5/e8RH5HJ3S8UOQ5tJZH/SnrQPd38NaAoB1ZwmzHAUWtTJLZ6Dp4hI2b50IVY2KOCvwF/3xfl+bD
Z19jqGu+HlQbcwVKzPKbJGpj2GktwM10styDlNFwEMBBKXa/CNG9V8RYMBTjeXpVbU8Sl+AwCJdQ
Awofb/ekmDlpUx8waaG7j5ojYbLzEHQAAhC790g9YTz8t2W7o6h8M1RcI9ICKZy13kvJQu0GXxTe
NXLyzVYmFkNVXA2v1VJtHAvrRjUn8jjzPf42GrNreRWg9EV32z2IV9f4/qK6xqdipyazVOINgNBU
DP920AWbTj0xFrwEhcQHQorW6Wloj3zcrQ4U8b4V8dMTeNAcWXPkIHHjQcpeWm47eSMG+QUGmlsB
0hxXJTmFDliIg7lUQ0WvfPbeksPU4gbZ/aSNmCZuzXhtWEnRNhVDoRnhsWGfoIqUdMDN+7QhNR4a
S46wetm3v4f+jo8mSEqjGRzYYzaLDgFhxo6qW/CO3U8A6Z1qMbP9+UNvtn7Bem4rXKqgMAuRUkKc
ANGj/P9AdKpUKO64vY4VE2yWMjCiQSsAKpB3Bs+nAUF0oanWX8wnh5zPpFHWu5vYEKyf0tgn76lT
AZnKh7CHoJmEKoJm8UF0Y8yy6eXMXqhDQKBX6eyR4o0Gb0OtUoGVVVWTwYY3IAoFnHk+ckPXxrUJ
5lNexe1a0A+WqFdf5EXNQSv7tQM4PNfYtfpSQ9M3rC2oo+64GLe6mXUdYamETWPV1DAPIhL8mvGq
hOLX0ywMmriPfxLrUgSiOZJ8x01fzxdOSeK7RZv7LcVcUrH2w+3kpwoOtovNh5LK5FoTn3k+TNpa
EmppDW8F7QeGPWuOK5j1GvW2e51EiIeLhxeA7IZnVLjenrmgMohXzSW5obNMGzRP6vf5DD6P/kIs
Vl66mgHVbrfV1ksSlXJ2E4vJxzxF9iAqfq9Y5NRn/o56f2Gv2oflzfEQbJv7COBTbxNdc1ug6sb0
3UGFNUg+0gNBmY8bExZn/IcgdJ6SANdBKk0Lc7D9Qd9kaFD5GxXs6SlqP1l43Klwhr73Q3UfgXaI
SPOFA4pNInKjKxTvSuThsEnEhykdEYux/kmW75qGJQrjS8Q3ISiCoAJL3rB6xMjgSkg5hRUvDJla
d9uCWacPP/R5lR3S8bW6eIdWtmdoktMiph2QrU/5Mv+beNNXE+RZukB4JnfUtTFYGxOXPp2a6sy7
BTK78CLpQpaoZW9l2DuI1t2ZxFN597SR+JuMAjXcvChRunAc2hcY1lL6YccRLwVbbxGxLfZBsO3O
VKiL8f/oDjyYCqlsvwOSvuMgpbdmMBUV9Wvk7+Er8OigSfdbfz0ExPy6hbB3GUmKtjznScExgSVv
kg6HIj9kwJNgnAWptEh8fjm659pWyklzABumswvmoosmWE1HYkHVPjirySFYNA9dJW/Hi/NHDF5o
JsD2snXHLP/yZoZagYhnkfvGrsdU3tHG3wNMDYDu3YSyp7CN56eC4YPFF4hTr7Mrah5Za39KqQk9
As+RtLtcyI2PWOgSXCFLE79pDuFc+2n+E7i+3bt3a9rkij1LinsVtfd/rCILPuX9QBwBrPaay5JA
RosVV00AyXQ/WQG1bKIjuB3qngOJVj6X8KuiwOi3oWUHW/B3/mp2T+PdfXrGeZr/915mm1KGouCr
W6B74PZc/9BPIzfdBt7U9x5KshneUPv7yeaipMB8TfY0DRQB/vtfKAblsh3JeCSzXsa+XtqLxlFK
hcTlp4sdpBT7yfBsshRAwXQVanukmL8etjUsScW233tReAZ7FAkm9lAKLBmP4tZGheObMqs42QHK
p/if797j1sL6d17t2Lz3Myg6ZwkSCvis8gMEJAVLbJ2UCrcIBY3GBEfgeWwA6x/2cCDM2TogfUPr
ImfAdFwlIHRp1Lv7/2LMJo+WaltLM31uug89bMJehy8rv7t7M1IPMLlfy/W/SikwMoSg+EZK+El2
aw8o9pMjEG7poNfnpkeXP1O1+VmS/eQMoC5S+Pv1Wd2EOigoGP9RsbKHgItVx9fvlEkqGNaulkBA
mlX5+dj3FnciBcCKzIDO45HH2EVRh3YJ3XcyOAFj0gI+pbeGosasbW/OEUiMRKXH7myUXgZlycM3
+aWgeJD0mu4JddFmATjRwWA4wvlIYM7hBz2APz3y9foQC2sKTdAMb4jWzOptH4o+ENvhviEbyeOg
PbG3PzwQqgRi0SKDNigYGLAau/xiO4z4eVii5wIwgdf5QxdkYXYWEjaW2vDXDx72Jt54Jllxzkro
sypu7V7qVhiTvWyDJJLhwBmWu2JERFi7nyXuhZrZLHnDpF6XX6SsX4X/Gi30lftHVamwHPG8f497
pO93FCYHWWJErrDBSd/7OOfzV3YtPckX7Xwm2e7m+H0KuYUrwDM/2G/lZRXOsayQrjvNBt6auUq2
LnJ4clQluL1B6xKEQ4t6rWmwpw1N6trYMCyhWdupQYppQU9JG7m3QAMP4sYDxHaAUQssKbTASB2P
aC+cUSTmRjiYze8U70gdDJdKovojyyHhO+kjIiqksVPVsz+EzbPMKLaAqBJYL1s2n0UAGSnCgG37
MnspKyuSD4AEmXPGOdXesbhGLms1nCOIa6R2Ml8W6NwwfHYmuWz31rLAXiaDL02cHwUQxQrXHivq
eqNtR9jjEIv6C2w6W7udXGKGigdsQtCRKLx4jzHGbyUdMsV4tb6Z26brDvrc7iPQhbGUHMzTXSOL
EUevq+TwdVtFl385spUoUkAccnSaATtHWul7JUfUqF2xPiWLo8KfT132k6bZah4ynt9KQthDohI+
W+rPrH/aGAihUGWlrm4FfG93eoRiMp3qWfLedkZ5Npzj8AQUW/S82jHpNS0vcq/Jz1jT3G55OSIv
uU9eew4OkkNHUyn830oyJoO3Fi3qvmyeX/rqSoCKH7YbAXp9gRXbYBl1lGG4gJaT0JYQRcxS1bXj
rYbH8Ri6eYXPxlygKZjPMuNLzwwVJQRCM6wtgskqagzAE+3Fks86i2Dt4WDVHPhZy5qDufXxcc2t
qQ/vAcpHioIyckxi34RyTN4I5TtcJbz1mLoOEKQoPdn67bBi5AWqq9876JFnWX3Psxn/zBvKepD9
evQaiHOFWz6RygmS8GF5RPhjgSoPUoCKLwIhwU03Sw+t2WqCJeDaYCkxRONhGUvPsToJVBiyvH4O
NtNn1GET84+WnyONR8jFdkanMQ0zHYnHw1WEe2CKSB48jNaV6gMoV/PrpB3FB3JATSgVzzY3845I
pZ0NYQzZPL3fcvthR4tvt7NYI5hj6eK/be1Jx8bukZbY2LxXakwdOBZz8vChZcIU+cOb9v069C3e
aAi8FAow2WRi9MXojOXTW2ZugezCpLx7aHymMGJNusumG0DN9m3rxG0Be940B9/ScYFMbtfuSNxZ
4HjETtmfgpZxhjgTKfm9ThKRypA7CQCR801MhQoinTjAWpULeKxdUkhw5XhUWWJk3O2mG3xHa+aU
jnbvd2dnniligf4S5CDcqNQn8aeu8KwVxxHztSKk5NHcNBpmeUQXILi2adfmz0Tc0KU4oJFhodMO
oLIW3THWGghRe0+BJMRBs44X+W2YYg4XEcrQ32P3alHsLMaJ5Hx0a+JPMvLhT+vAMQ0V3Half9rc
g6GMD0f1icLTeF7CJl9uk7D+eDRrdlV1+mWa2FzVIz4x2UxPVZ3DC/WPGAFMP/bKwaszW4o9KA9P
fy4e4WaVPgQydTrTxB1mWbtwbRmXF1/u2GYHj7nhuktYIU2d1Hafq5/eztBqpGuRKtz4UXbE1htW
+1nlDVpmfxeeylEeTUfLdDYvPwAYwcAfIu2N63QcaJjK4rI3RMhlVRgZCXqUUssUzJZj92ideieW
jHrrmvjYP/ytphj6KGYpzeso6aFFxWnUf3+gpOG7SuVEdyc/frWJdWHc87xMWwzhZdULBX++jdaH
11MqMgeGjj3SHL4H7LAUFiUTygT3t06UDzOqGy34J+my7SYuHvbqMHYs0rjbtf6iyQacP5h+oOPW
Sw9Y5HgeUiQDLuhuKGD4JdBZxqVDndBOxJhoqpu8y9pKNIjdESmXbA7CsfnMhkmeBeXEQfaknnnv
+BMOzklRGAsCevuHyZJR7jqB7+LWWGXhRlTMb4hRytdnkSiQ2ORtW98C8kTNF8CKVIx9oTbTKrw9
CKeGlAnZ8UMmfllkBLi3auqycnD4OAGcUCdw9gv3a/BCMzGvAbqAxYnLk5r/+1SKYBrQZYCjgTDv
msRSIZD1DH9PH5mYiz8QLzyLmu18sNl1U1pwwKQvB/bI7lYBHSybcJshqaytZ8Mc4Hfer3K/T3iz
lL+gJf/HmJaiHC6W8DaKf6G20GokMLCwKvaN/AurvXDZYtBaShZ1Luw9DvaVXm6EmOF/3dHmYrCk
QyG6sLfVVpRotAP7xbVHmkmCP6yOZYsmXla+Xu1RhUEuiSZSHcc/VNscrhiWSHFDb0fdeP8MoUkF
9OaAzoHssE1jS0eP8war20Qlb+oe/86zaj9qmevHjB/WcbyxDDEEQgIG72v+gimLTP2rTdzYR/Rw
YqApc3Bms79xnJZhsG3HiYI6bpQlBLev32BM3CAq7xlHeNG08y4zl5fXZeEPWfLxbInxpUxMTSi6
F3/2S4+ZL5aSXiBDUAL/sa9vRdlOm8Lgaqk5+GIgayxto2Aau4irnYjKRcOR/sz4wtGfGErwJoKe
8IPwHoSdtdPhFkooufbxBRcODegd1RkEO3u2Oi3ZvJ/iSsYTHRgzfZN6rOapGjdL56Kngq46ai7w
y9KlES743KD0spr9ega7DVP9IiQHALFwWZUNjPHAlmG7dimvV46s7DaAlF+kzYz4lhqT0XyH/oJ2
umB64rl8x+ErivXbQwbH/UH+/IExKUxb6GDYNhpF1tCzOLx8CQhr7aox9eJUTBMruezfbNMigUew
dyusuHbQyR9GURE8xre2VX4OAFwbXqiEWgvAgV4KUAbSwFeEY2VKIA4jcNxCzRAag8WQFhkD0UJr
3uFLsOXcTAZ+HV6yDP46GieIxVkEos4ndDITjgfsVw1Jh2IyLjmIwTVAJvmzKP0FJfge2WSBVWFL
yfWInz8Ymwdfhbg0p+Qthh3u+7bP/rTvgfI4UvWzX3ytkX3XfNlcS0eTAFcWLadZMcUqsEpkXlWL
VgBbKVxEkBJe5j0urTGxIDCHFcfWlyfv40b62RYdiQVvpBeiixGVZF6RHZqLTIvl90lK3/WQtTVw
MLIJ56oOxHAFoRcUiuMab7EIgc6fQ6n2TrDV+SEWEtPFAMVBPyWCCDGQGhpzEML7kwZ1SlIqeYc1
r75LB3w6b/OrF8XNagGkd1rLt3RF8g/89GmEfbqNDyW5KB1RHRoDoma8nuIZn66LYeLnlxMo4+tW
2Igu7A+VUotYyk3Fx4VLMXzrVsIKnUn5UBuJj80S12fnS01o351gEUmW+6nI2u8h5LXoMEt6D1Rl
tGg1Ib3/GqviBMj4IjWoX8LKeoYSR9WkNfFIIpSo9lRzDioiDuo9Ao7k+cH3DgHh4fycWQadLm32
XnszRBhjBc6rZhNqujX93I3nEcg2nQG+X5UsOlWMzqpkFUAdVjCpKu4Chkw3XqFcA8uonBpfPJx4
sjCga9o5uecCVY1p2IDHiF3VCIs8ECQ+KRkx5EBlpfPLcyRa79Z/GAMgjZvjrinkLcup4aEalSiN
RfdgWVZVMp71kfDM+aX+PJPRb/G30mJTnZIBjDJ0FiohkfrGVoG9xM1u86mVYqiGIF8T5dmRqtJS
J9zAj/yPEgFnP64qIcfNnnxvKftqSroziMVpZaFEIOcLSFgIH6o4usUzF6qMGI9+ozeXHE1OJY4r
1Jz8rQeOTArepjlaM4Cfzl7Pi6mrMsRR0I6j6LfyTTUylw+wyjp+DZnEHxocJZEWddqtX4aB69OG
zn33b3dRFlB3tgm32WiDXozslaYmHxE5B5HF9ghiZ3wrhs5e67fTAdb80kMme+UpW1ye4MuU3tqa
ZgTvXelnY8PlvwD1TnBYBeCculvr93GENeOgB8QpOguFHKhHbrGzO0tmPRUmTHfvzdiXCpZryr3n
pqZOxhdBSysPCR5/XHKdPm+0IUx4JtWSAFNxQX+Ug17/8ZI5wSYY1FWSNsfgUI6eu8Ko2ooE0EuL
wRaLtKBymStvwcBa4wjVxIhJle8c3LijUZn4GS9r3iovLpKSAvG1p7xWjbNHakSJR3Tj5TjIUW6E
HPs/DUfPkCcrWDtno0tRsqPJOSb2+1bUFM9lrlKL9cK03nMyiqk/xyaz37UDpnUZExcyls4nwOKA
JsUNG9P9LwTc//DQJN6vR9uhuNnJLyTh9ZGkQQRrF1A09Mu9KMeAlH3AafbsGOGI/5sEihI/6KdL
rJxHLwtR7SkJs8oKBltgsCBsbViEqBsV8WtOlDso6+eHPKYCL4D0NkD7hQbl7KHrE0OG0G66CUFl
htllouwNHxt4hMF++hhiS246fAh530F3nI8VdG5yKzGx4pL9sdeaGz9aHjrl5b+p9mQuqcfI8lxJ
36S4wlY12xJfpTgxDmimOe6qSsPLEksP0d/Q020CSd8Tqru5lxmB8iLtj37yaEWL+AzLs/2c1tHx
yoTOwz6/Sh9dXv1SoqCsOLgSQz0KWyxz97dxlfpjoM6Yg1dLKZCXg2OKf4PT8NTmnS5VNRdKL183
iZeefA1hvB/pPLRNVnetXzDT9UOKdj/X7o50ZfrYW+AhjtxPjUBgsSdPU7PBsFzUFwzilVpJMjcm
nZwFfN/AlHlPQk86495bthbOxgW5WoGxuskxLmdPNhUTbvcwPyg9hn4Ply5zEgw3mpWCTtIfOKK9
mHvPa9dqOlx7p5lmW+ACXwCP6RFpxPVnjm6231woD/hwHCPmDuAam9KClFBlp0nX/QyIclZ+XapE
Tj8hYT6EMYDIxgM7o8kSNGMh3edrgpu4nA5cnfMnFUHuJT9iKIGdmXkTXnqOsl5zbEMZ89hhmGTb
uYO9dskCUUQC5MuBqPf/fCa6zQCcF607lvnToDLHr7CR8azenlNtsN3lgF63coc6u/oILIk9az2l
JN+VQwFPH55Y6qn+aG0imWstjs5jWodb/KzvkOa4aRRYUHun1QX+mqX9XzmVKeuDNV872hRbdt1V
/vjAVuvERh/5lkjWhhcniwEncP4xK9MqTqjstoIvjlx9Y8p/GdrZaPBinGDswKBlIvMsRwAlKm+F
tJlnFTnNAVj5NOrKic8fbyYHx/AobCis4CqRRuWaqATJuRKQ6q7fvxlDd9ffUVpXNfTUKyWoZjdH
eT6hCFmwCXh3vN6WPCISIxDwp5R6PzCwIe55BAHJSyVmEKOcPsf4I967u0rAehmkmIeN+lrgXHcj
0TrH3YoTlxqoCymBL7b6igPWcVvit071b9TfKcb3VADJqkTVWw0fPeFZL7lpaT5AgqNZslyzHpmW
cKx+yx00b+VgGlGI/iH7lJr9nxGRmxXoPgrArBcdm5ylufAQSD4G1grHwHHAsZfr65k6kLYdYb37
fE8Z/afyiFUmrgF6MmpjrzQl0XRvJZdpGns0CBz8DHjBIKTgVP79n2cslmo/R8IuQl6L7SQAATrl
j0oaUF+W09tluYrompUsYODfgdHJIED84CmA4dDMpcIG+EkXnALLSn190QCdDAtkx/NGwvgmjg6F
mjpXPnDZ+xup92gt7G9OAdSF1tYEPzid2HgPCBPPK4nyaGrhZkj710QHammA4mB//uHL/AZIMSeA
p8fCv/sqlCGJLFwc8zv8sSnivYCBSYmQukpyiEmKdiLnhsNkurwAQtZxbElK6PWdixhvN57Kowuo
5BJO6/fZPk9JWi0MvwekNWfZDdAipzA2yZb+i4DmnlaKhRujQge1mx8EzrMFe7AxDcaa84yRS3Gr
Crn0BQwdqiLhVPG9+WURO5aqEFp/2tZmfWES5U16tSNPAn8GqO7kHFPt+zapRRn50SRGd2YVPd9w
oUGaq8+X7Fg4Lk0nt7Chuvs49RFgZgWiI/8rnykJg67U8i0kciFhPfNg06jTL1I+C/YbRogpXSzo
hXq5oFZUkXPHmvU3HYL3UC0/pQ7if1p/VbeD9lzyHV0QwBHBXupRvPSZGO5vbUUBvFliKyzm1Fkw
94gJiX0qhhQD5Ket0hkLimh5d25HlGGHXwtcFKiWOB9kXUptNiHNmqG7hApxEdbRFOi98jNxmBr8
lwOLC92ln8u5DUWWd8yG4TwFmiKi25kZvKWcTkre+x7enMEminMCJGJSRtrlDsP4EFwsBly6eAbC
KfOfSWKIoDC3WRwsXtaIuC4AzgSQQAXGic3f9u4IVIeiprNRmumLCxWM06/WOKTRJLqxyWomIfAH
rWCjIHFK6p8eFmQmbZM28tXwy9XeNwnnuonjv1wF4L/+eFlxYk4PRoBmZsLUqsa2fHk7aQ/b62Bh
eVuoy/AlFYoJv4gXjyOR3IckpAsqEO/Pwhpy+UGGjAvmUiCwxILBo5tdZ2rqFClMUz/Im3tjS8NF
UGPu8QOc+jhi9uLwYV8YzWYNQxkjLa4fwzEzNrJz4/0FSP/9HvUBGUAuaEEHSmaNHzWrnPLGnuYG
juORfxiiscjwbD7fsy6DX2kqzPz9wNeYUok5zjEb+DSvrwL2yKsthXk9noSuWuyFUQx9uZ+x4S7T
4kquVB3pzThMu0ms/GJAxp8heOAjnKMfHZU1FYOgq0GOhi/vqAYZTC7xA7hbifuZmB4VlWhmatEt
278DxYFlxEkQOg67c05haoki1b+I1xOUcbkRDDaZUvZ4cFkWwiR9sBUzL869KeNL3CiFLsUIlvNu
oWYcvesaHC+2ADGWaP0xvg7AjOszKXIxOWxVyTH7jqyCOZJZ3zJxB1zZ+t7aZRcLn2LAnGTcaVZi
uFqUn8WHwQPzdSpHj4Cov+XMWKqcL/GFkyyoyFMbdN8hgqtPM7w4mbQTMCJ7zgQrCu36YvqzpLLR
8A/RUF7ACQJZwWpRnN9mACUlZEgaJs6GAVlC+R0ZkOVQUeXDBoWul0cYn0VOW3Me6+TojooWh6u7
W8uvx6fopL20P03OR79UIvNOKo49ZK8+URPJGMmNp1NugoLESOf51f20WAdwBR2ghmUrU+chiQfD
3gS6PFScFFvyguqxOLJGJBahfrjj26Rn7oTa4uJOMVf9u8Rs0JBYD1U57UaW+Qv+SXyDkN4dcbh7
2Uj65dEqDZYlDLFPPlvqiJGL8NwRxEdZjxhZ+3bCJuQHUCCC9rfFwi1hRteppbTBP3Q15wa5jhu7
YfRm+6EArt8jDVMJvXFDWJjpXa+hP5yUulfTVS9cJZntQiaZxT12at/oBVqOtVGirL8a5r8gFFQv
Q8IUT62kmKOhrK3x8cFMh4wZYHGrorrN8pnhrXnvHzyuThgbWF8pZ5I4akuuY2KDJuR7XiG84mHQ
05bDxfbEhgVHppsOmSeSlPdtSnm4JvG1bBVdyhHSFeeF8uj97d1IppjET0IZ/Eh/WBuqHlSNrVoR
io0rGqns3tmifsKd771p3b7ewL8PFcil332qgJJDQ7+6+wHkfxbG6u5oTBA4x6aIJWaIfbgbMfc/
Taqo9FNVs+Snhx8XxcLqk8WZL0Ocf32hr2ku9o8Z4rCYioptd0+MD9qokuaY8OFa1cFsy/YEAhmk
XZaoZFbDlf2A8lZPcV5Rn9cBvGx6vIrrvI5a6rQZDCPqol7Hk4pswOBhtgIkcsZk4pafbgtnezDt
PCO6p8mmHtEtiT7ePMOyjPaPSV5nb+ZNXHHYbDzUIOSkSJNvdLeAqz7OHyyZ5f6jU7xNiIJzA5cP
7cqjaCmdpF4LG/ndH35d0rxZ+Xc6BICydiHXAcxSRAfG9BQFJgrRp7t3hP+67sk27NiDOiNUnxPE
+7+zLYzhJCFWsbxb56xT1htGInSVbIG94hSwGhy+STT4EXaudwuvLXXc40jL/7IGQ/dR3aUSHPZ3
qBR1qEuRb0SYbodo0Wsy4QWrp5/r2uqy+QWG5D/wFJ/L1GTtP5izEcZhVR9JkK9yWoRcFc4WAVsM
VJxE410raoMuZ3a2dqRInT6Xbl1n/oqTccmTc8qOwsn6AzkyaYSas+ZHM1GsxIp42vwPcQEUdsoU
0TUs3GHoNxNgjQyrgB5A9/cyNkKk3gvXeSpbHxONUoUSLxO6yT+d5TEoei6+6j0y9+v7XnBWhsoU
/fajYhFmHiU/kUqT8rdNC8Ny+O6wvQqr0cX7IrPMcvIk3u8Y76P9ja2TnwcFTkzs9Ajv/MLqtvE8
zwzX0V1qmeOSrm01R8imAAKiLMpuX5uw3aCqSFBmFFN/Oiblq+Y0mv6uMK0Lh1oOKnPKpNHt9A0E
pMqjl1WJPE2GaH8zk8Nv0zN0LTKks0ZQG7nGCLEpBMQ71TSs4mT3g7EJhwqEp7bKoJYTto+PUite
pe6V0ClgUdHrpaOhq1bLbr88bnDCxMuJPkL2SSkXtyFlMHKHr9y7O1dDiqz+x3SpagTCDADAdef3
s6+huDBjAyHFZ+v/m58kI8wSGVashhft/22nNY0AvlW3oMusNZvnGEDUKL7w1doc+O+091QKqvNR
l+S3j3H6AxmFUr5JCa2EMd55HuP9/NynZt1P7zfSG3cAANnmYcQbd5y14Yfq6Jgr9e+Y0wT5SHxf
dCnwzD3p9ySCai0PLLIMFUdJczXTpR/6Lq6oKU928Ol/YXl10efXbPV+eEdAf37eThSunmuDucuL
II77eOKrB8BKZ8L+JaRg+anz075kYtb2B+M7JVeroSpradGgTrJsZ3J6ULOt/7nO+jbdHb7TxkYa
e5Thb0Pq6kdaa8yp1l20E2QDHQxh3gwVuvJ2D8sSZNazY2BY9QxSa+ByJQDzrTW7tb8jBZrfEy4d
+Yrhn2Yk1sFaVLsatYmGjVf/FC2bb1pkkPU2JREyykjSUgZq/uqsGh+XBVyo0IUgLuiNIss+lssr
NGS2PukN80QybUUYCkjH1BK7wwouVrw60BNBZX6AFKIiQenLuVF4wcEQ/jBLth+1GlW3imnxw/j7
6WdMc+aVIsSI86/UqrbUJZTHZYrxCgyT6XqUvBKCVCZXQIk+loPYrHtD/wC2aiewTimwqS+bJtc/
HaPKDJmWS9OPWQEq5dJibJ/nvLhtNy7P1hJviA/knL2tcE/cZEGxdDmzNIN3lCoJXSDZPVa4A/m8
7aGPvtY+W4CCJ55dfaGi8nVlsUIJsd1LUR/so+BatvaaDiliCsWHoMHDfC3w3Oz1bJ1tux6YQ0Vi
qSQtIMksdCjrvOpCEjuwjw/L9oRyzTK519A296F/Gis8rphWiuLHhqV8acR2Z+po1PO6GQoIiWYU
gG3zrrGA4I8lJFicQ5sTXIUTL5t9BNnW+FABQXs/drUBoJArJ5sLJoldqT2G8jZSNYeAYqMiLpyC
2630MP8tirqmSPuZK5J+yeZnrI6Couo3lQ7ki+vvNu9hxYhe5YjE1C4mYn/M5gE+iITrDRU2odfa
AEfkmiIItNx9HAt1ikZbmP38HhPIjmCrG07kGKUY63hr1lFFBQG5xGqzcAiAPxtuqDjjSHuJq7l6
nXAaWXtvM+2JneM7NWjuEXZgI6zHIuO9+FtTctvwMbwy/hw4cqTRsYuoUKyhxBj3By6KpfgcqckK
1EkekhoLL7ATUFMfJg19TiSNLPzSCgYcQ708Us35wYX/KFim2a6NoVG84P/cFie+H6EgnEEGgjxF
tO0ig8BWu53Efp8V3SXI1cdb1pmL3GFDWLQuCG1PQ/2EuNzBrf8D9dB3VXRNfKYqlFVcMMPqurjf
9III0+YL5hm9JrPn3nFk9BXuHUFH4N114joJKv5s96RZMJqCEKFxDBQ729WRY1wZV7OAcv89Sf7v
A3IUwJ+iTvP69nBk6d0W7bLd9yoolfx5gMtch55Onuj7SNlNVjsXLnxsRmfbuKvBulD0uZEn7JhS
sUnf9H3qnFRFMnbA8czWCiVmaeciw3kK5F2KK7L6UouqNBAeu5WczhSywTPBGvac6m88pEIMNfzE
QN7z7PBxSLJ5Sk29VGp+7TepvApF0eo9dCerNVsMG5OXTMp040TQE3MY+1X90flPnxLWoDhFmTaK
hHYtU/T3zl319xhHSj/r/TIJBLFw6sxkj19uslxVEXsEgRJzJuKvACu2RKH9wIwEAbyEibODTuzT
/3fDAxvFNm0NGfP6qkqn28nht05l3/AmDieDD/o+j4QapgUuCb5w039VGY3kpID/rVRTAiDBDq26
rTANrsUUOm2f2BtPftaBy08tvtLYmFS0hZAmjA85xfA9jzbX7aQkLfw/aJO/2O5/DRdGxMcUQ0z3
ba09Yba0rGnsGrbbEpFYkjbO578MxnTTB71Kt19BZGjnMvAk6A9NHcVG3cpcpqmCCr4BuNt0RwmH
Vy03PsO+aIrVNTBLU0aarDpThvUKc7YyoVbCsOYxEfaHayV3CBLpw80B0DNoObCvCbtnf3Gld16O
BXjaLxiUNBX1A2DC0ElL1sbJB4XaguIM7VjS3QjI89H0linQyd4YaYQXIab0Jxbn7jRZZH1UXcaT
rQTEFSzdcu9V
`protect end_protected

