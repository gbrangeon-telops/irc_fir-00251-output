

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SPpb0sHtYr+7D0Z/NdHkBGKHFj6bPnAk4zCT9Qd9jSi/NZdzqHWXjKwgFh3NrYG/AQMVJcT4R9KU
T1kWm6bsuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PM0w38wqoKZTqxD5ZMv+He7u+x4mAKOhS9vNWqYsLtlMu2ni98hkp4Js0D7iFCQdcFCu3Jaj2Vqe
E0m1H+UGB6We+zPa+TnTKUC9+mxtEW7xpi8i+GVKfIfe89n3euEibIBIS0WLtZypuPRjuzr2TWw/
TpBFYS1oUTQ1qwWguI8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OIEbVz6QJBHT228fhImFLc7Q94gbSg/QOSgeKpAp1zRCxot1azeNL0EHN3pwZU9Qs6kuTNEAn7+w
agqdilWN9rl3uQlRBfW5KbIj2khza90rK/4UYrbcPGQyMxF8l/LBS9RaSzH8pqlJgQ4YfgwGNaq6
EHHkNL7CBEprP8VBO3A9geAIYBWstNirz3P/01jzH8PT87csZHkt/KV+1ancvBdl8zy3Pi5RrOtK
WdR5qLkbXJ6m4DjaubrW8HdK/fqusuCVkVGxmajuQw899iRpx5AiTEwKYKOor3msJGxdK7STL4ZT
S1m+Ec1GdsxDwYBgiKT0A3c1/unIYBS6y17V2A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y9qoE+tEhAFEsAZgxeFxNUflksEoY80RYly6rjz4X/QwncMYkOdY5w8AxmW4IYZfWprQfyfkxMrN
8JuXogLHC84iIPhEFIhJ/+RivFHW4gCUIf9NTOGEkQza7hd31B0/7LZttbZHcfTR5stmYGMhB9xi
VCriwe4C9iR9zFvOJxk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eCcOM7HngIZB2JCDRQ//SPPOptJbtDQ6WJM03A6xR3t8OhM7+MFavTdB4aR11UrppwUsYiZCHTBc
4AdaSSNbTEcILhRaZMNZ85hgqiNgFb3YTJu8ZIWifM+Ad5U1zkzbH1xsVssRl/Sl+cf+TCDh9Psd
UOpjIzWfsyGgyfaSSbczC/DMklBqFcyspqzOP0YGdgI4It3e5xnwDvYeewRqIZggj0RyjkJH8PxJ
o1XlyTZFQZIIFN0x8sDbcPdsUekU3pOCvI9JK89jigNzKmLJRotLEgZQt0B8gMiz/gm5u0+k01OA
f/7Xo9TSexSaZ5evmswsNTBQhg4v8j39bgkh9Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7744)
`protect data_block
E6+SSr3h845VCNcI2I7WT3LDbD9pP1FzpP1hnHtbji4TS3ovcIcR1a3XBiqBDzsIL2O51AvbWzKk
fZkSNo0clmAHz6NYw0I4s4WnguZ5nyceiKUSZRqQ0G+cCKhXmtJt/31Dy4ajulEFx5Nvg4NHpQu0
BtKr0YmAYAYYPfhNPKydSMZUaagZ76knZHEmGIop18N9H1zAy+iDAEnMswIUJlP5x/5FY/11iyBg
/xKCd+LDJjdqUACbOwvqom99YMfybTWNsZ+6050gZSJY4/7g+tFNzbOVim8akDDkQWuxPPWEVXK3
xkHd+ckb6zzwhnAfOljuoIx+u2oVKojE+dtFRbY7SAnyj4BAg9g3ettkm7WSVluSGS9iVev4bfp9
O02xyhceW7HNJgUDSH10ukC+ZcqtR599DIC97ygrnfuLUkTSFTqiNWy5HwA6tK/qWwNbNNevV7kT
Zctse4IUpeUxPtpuC4PkzN9sW+y8unJkb6dw3LBcPgR1zdNr8PKWltkJ/YR7ElRA3WmdIEJBJ7yH
2cuiafDTBbHqQreJuJ+AkxqB66Dbtdo6ClYjKsPF5Jwb8AOvorai8VwmrQ8SkoqX2qfm5beQL85A
1yVNXAQf6NDCtB0l/NAozGIuIlNCLX47uHmlJzen+W8t3g/3rjEHfJp5YA4aVP9DhknDbMSkor/F
tbLnf+x75eMmxuvw7CATgR84/KU5xuKJOKhH/SpbqmgVY5VENVxH37CjSIQRNari4QTv8qW7pUNw
bhfdGWGX7Lfz0ABWIhTW4WhWuHnjM6kg8q4hixLsKT/9VZO00sKgL6dOi+IM09exN9bHNF8vdpcV
PcxTIjvy01GEpb08zt6rd/1s9AI5aU1kT3/FJlUqhumKKfM8fqZNFt2ccwAeoi6dfF1NOcfhMvvw
kbKOBxuk1xeXynLuuG5Sij6+dFEGIMuTLnUsIVMagDID0SOpUakOS34WFKeiLxZq2tih0FQ+4QdZ
N/jL8fjrP7vgg22l3RHkF7A27enQoTLwBuiCHUjtePVoClCdV6vKSGPdCztZJmeFo9UP9VncsI7P
lOpee++n255hsZfNmq2tyZPkosu8GpBn31vWov4XlN/f85i2TcYBeyxca+cexKuU1JBbm4nm6kpf
CRZGfrA4cGhBfGr22OE07GNwC+ph0mALnYBy5JATQ7zpefHK/r5wLOse5q0G0IPg0Lg/BdjGileB
BH5t8zXe/saKBtw+CabVg2/r1lH6pWSRMxkpVEftnYhIAm6m8zomqw4O2/ym2E161d59Nsb2A/ZF
m8eHY+hTYQM1ntn2td/N5CafKYFfoetGsj9CyepX8Fx6i6w1bxlFUzw87/CK9GD09W+ZfgwDxbcQ
HpapjIEGCLaNjR/aeJw0TKfPJ1b+OZeDxjkb6YuM6/UeV9V4J2v6bluMeQlzdU/ukk7yD4fwV1a7
By0Nz6doW0/WrZIEbRy+ac26ZOkbAOQ5e1j5DQZMoOja1TpW6ho2deSAXXtX/B/rDorSAzEsTAi2
Ss81zusurOFR13UKPQLGef3k4skH6aArETeRum0fbPPHJxqDIeVoGYLHaiqiiwCQVfNoWsALXUhP
/ykmtpbRxFVEda1XeA1iTey7LW1j1xhBAc/ZX+EYDkkUek2jpMJ2qIJ5TdNDBMitgcy9vDblTz6Q
hjnSmVzENolcdgj8jtSrAkO/LOpwd86P0N0QxGyMmRjxmu9p1N9wSNKdo8Q3Ual4w3jq9jC7gVw/
BpEqybeLx+zbLqz50aQEQCNo6WgitMTxBgIYESCsprxorHVlNc9IVj8UNAtNhSAb6XT3A82avSx8
HUjjEREAlBNHC+9Df7Uz0C1dPOHF+SNf4UlOAxHTdCAA5XpEI6yoWJreZP81rEuqSXs6/LGOmzsj
yY4zndgVxO+CN382QRg8Y6cUbSh6NuEfAm5uh1fqKDZ2q4N1pDIGqPsaT86sCGiqBm/c3aRebk5K
FXSmjtyPYFzhGlDAOzbxQxd4gXZhRoLGL+7S3kuG1nq9gOtheoXvy6okoewuQXbjIQgdnMdJtS0P
kPgcYoNj7kQWghQcxw2NA+nuDIPPUxeQJ7xV1FkRfX8kqOwDuj+CQLkrg6/FQJPYXz/niQ8Ek54s
6mTrixhfPiP89PaSQ44CRxCclDgeZsfZGfhLM6MptXDKIcRZSwWSO2nOoQ45JbuqLUlmfyHa5AJv
nmsQLdiyvk+kJexEw2bAuP7K7JRyi7A9TTwBDipTxDi2e6HTywqnX6GfTwxHuX0cTrPTZFPK/+SS
3tp86p/AT+4eAqRdHxkRf3FIQoHv/wUdsitJxMHFkaJLgF30iKEHL6LdPcMz0tAITAxBeb1i2iXN
oHk8WpADdEwIT9+tr7iiKIhLQrsJ6lxFVnVaMQcLKLgSt4lx5bDV8dq7Gy2LXSrRc5R6oVhVKGss
qAd9l3XeRJFNzK9u/njv0lbhpyNLplKX/bY95wRtjN0OnvZXJkHYLK7pm38kM397NTkpbUM20/PS
wvNS7YJjs91JqX56jzZuiLXuQ7mMyR+A4XEkjdhwSm6YNNq7ueKvQfovV+ehoTJe/HBjPuD+1G5H
oRbqWVhhCLOuoWQojHIDvZ0jYDnlGNQpcubfGIVm6snXWYMkJjark+lBi7sKQ1S76a2LG0bAuDcc
O3B7RUzV74DhpvdO6HA/RIHC8/K0AV6HaFElytqftGlQxb0d/uSpA0fSmFqlYIgOLr1wLRwYrweM
shxkUTSC08ds7jVQfQtXSJPqXfEaEuNNBukJdqOxxUnDjzGbtnjuxaxSm9fG8jlCu08AwNsn8+2y
unIQx008/PauYdUESLVk814yBk5iwwpCawrsKEBj3WKz8+55b4MNe67M1pnFkxm7rfWiBfnqZmBp
9pFRybKL1IhY+M8gOeyUObRIJZJ0qGEpnQ7rE5NtfZNrM7ZtdiaNBQbuHZafTH5hfvRtOC7B77Ws
EaEE++hMDus/bumuFgTGuyPoilNXtgSsHOCbFUAIgF14c0FBI/NPAHHtA/+35XR9U0UuvVAInfPB
cARdp5m9jW+Iu6rwPbeJLQ1fScgLzDz6BQE2CvCxvr5SIXVO3/LMeox0vDxiVHg4imj3e1rZE2li
RiZrLyzQ7fvqWzIdrqDjAQUSbsX8bBv/yRBhHAX5EjStRlQTov5z3W3kEn2mbPvP7Wwd4qe3GXyj
7hEUYuYNnqgzuwpxeWm9cTvepoXTiZz7m9eu9cNjtKQGc3PT6miNGeFv59O0BzlmL7x9qqgVVg1m
zEJk1Rz1GFr+o6xEv4Kxx1ezr9BLxEkcLs8R/EGD63RRxZeFrRmhhhxyM1JA01+N7ZHEjV4K2T0L
+ypAhOZlE75XRGm36pGipT/ga7m0NWOSOhouy1grhG+zQE999xOE1VpAU7CAvpy1DZpyxhf2DeZZ
1Bhe5DLN42mlss0/EsO519ZSqsBOLOGbG9Qo7vPjlZdSl+nZ0P4bp1xYH4xMxlHkvKAEvkU5h31y
4MH8y/rAGAK8iY/DK72vZLF6dtEi8oyZcujgKZDhsf1/FEBnO+5xYt2tKVUPUJWkKdFJ3vol+Wkd
xV2mfuybE8Kp340RzgcX12EU7opxn5DsWdKAD3qDa3ZT9NrHCYaQtlRg8FPx9esf9pOjvmZisTUV
KPS0mgONq6LBeoDPhfmnwQQqCAVLiFfoymd0pw3o6qvdM1u0F1lQ79K5+KpA2rtMfgPOz0akGJnC
8MbitBbfRxKJEhFDZQEHkexQke8M1oDoKaN5K0ovYiTfZgOVkNpI0ZVK043PwZdSEWKla+1BfHlA
Hd7Z1boaALmfEhzYtY+PsJdcLpb3oLzlzBW3+C4LaZA0WWE6x4PiDssMREMkrDQQem1luXf9368y
ipFBOgd8DUmo3pPMDmdeLsG31HTdZiTXioKK20Ll4ePESlD64DCNHUkhOzTGrEz/3e6wxIxoVaSp
vYXlbFsmJAp6IgHIRl+ld1lrroljFOl9ut/SInqbiJ2lLro1UhnfdX8pzrRqnVAemY28Or02FNV5
e5SwNL4u+i93g1O8+1t2lN9quTdqbWcwKf7v0Kewi27iP3DxTkgNMv13hSbYrt9a4kiGz6+tIrIq
9VYh0GQykGrcz/SaKCIPaCF1I3tk/cz3NSWPBAzn97D/xhC2X04JO7ZVZr55QrCNMXvpS6MJIw/V
VU/MBSwHBbtXZejp2O1LPvSD6EJOboGMd6C6nqz+5/g1yhHZLUoI7jNeHvKv7OZF2HIVaR6haD5b
mz6yv07Gnn6SBSeWb7VEe1SLv3vVaxi1OLhw3KFtRRaf5XjOfup5BzmrMj/RKc+LPQ8E4t6DgrTl
D0BNkAfqbEjVGQR4dKcrmE0j20NvzNVq56lsLDxdyvE+MBEd1XnMb1/p+dSzuq7a5puaL/v+LD+a
0sxKfA8AuzyPDxgdhmhHT7pXlebyWycX0PQlLz4LKGwy9Xv7kk1LYmdyGiHwl/S0JeylLQPuMJ6L
xVGMCsLJsVyh5N95L2CMPmGSoXedTe40uhjbGtdg2fz5A0/2W+LoM2N5Wt8pbYqiyuJ8yl3dqjUT
tflO317tmT6pdYB5nBem4xZj+9hIzCNShnyfprx+sZiiB6yUDWCv2yLyzSIRdCaDTAnPyUWh7g5h
TonpRoSiUy4ZMKn4Wi/occW7M+eWIRVrH/K1luvy0OYxj+f9kJCoxDF5sNZiG8eIorqUoXwNyy7T
ecv1LiElO3gxbtWCDSyp5P7wZU65fNQqnLuAUPdg+WAWEj8C/KGcCirMlP+pJ96ESpPjUclJDyVd
/QwAZLCeJeRQze/CmebOx/yz6KdNJRFAIGt0HBzmBfK1d+IbSCxrxPQxQ1BSWmaHS36ze5YWnJbu
W72jKpOh4X4EG4xdlCv8086QWisaQMvgfxOo12LXTfTtecAMwgippgIisn7ucTQBq3c17AqpowpO
ybgSiipDiGcY4I6ay8mv5VSdPO+Ak7HOl0WLWSL0vLqg0c/lfEBHyamYO6Ye+m1jce2UNX3I2ubS
wRsoaC8zWjt5EzbKHHshDSfBZXrcL8cneGbnIQ0xgYgnjVOmsgjhgK/6F0xMDGglRfAJpZ5FoqKH
pwWTdWcFqBRQTZnC1CbnzT5hSxk6WgBKvxOPaLSVRzNeD72kOrilGGQqrk+2lOIFy0Di8pC8e62i
22IrPA43EHAJ8986w0kexj/XPBCqfXMofdZSWVa9gfBsuR9J72rifGkQL2TK1lmfLUrM7n0DjMwx
kld8A5y77cY5H1kw85TNHqrUPIKGI1T1wDfWLX08owbQfYnANEQhWSrFlYkL8m3rQDuWE1t5tbjf
tzwYiSewEpNDLk22KAq7X3HWzozulxIsoAEUYvaUg6dEzZtoZ5OmUoE0xbnaGRgU2EvhDa284Osa
g/t+EJhDvaux+0oXCzPEK3jVpsdRAc5YEYziLmo1jztY1D5BTfhXDgBDazZlnAF6sxL07CVCWb4c
XCU60YLywE7nXmuzkQu6djM7FxTqL851QGvmeg92j+WEMIggGSPK85Ms4WvBU2suPUyw6eYdYZMr
mzGtjt4ZhELTXMF1HpC/rSZeqsvSeis7BpBZLwnU+lLisYH+COTJy14snbRdlEYlgSVAQ15G/V4x
j4ooXHygNULaiFizlSM+aP0ptbHezAh5SxtVM/XQG3aNUtIjA1gBEP3Klr0Zpf3pb9+0FkwdeJ3O
KTPj3mtA8M6GtF/I9X9nmyRLG1u8IRPJ5qOuu2/IYQ1aNLMUISwpIDn3MUJ0eDOl6qLKQhinR+QL
IHOSgRi/LtWX/93J3rcbFcYRFIMxHX5yS2yxOHhf0RXgRId24q+ypsVmslMQ35Jvruu0Uv/NlSD0
zNTbHwXyFk27Nmy/y0fiZQ/GTdlDDzmI0FZig+2iY9vfvl6jChm5y8q3Tp9Zjf5UAtrvv0XrZn1x
oy9hnS7NfGRbu0Hnw85RSJn8fv8LIAvp5PqB0IbMVuptpeH+oxtX3NeYIM/5pvJu9Kef205xqVqY
SqroSVLvmyTCkLL1peyGGKi7q2Fyla629FvYrYGtpY4hFH6fIFo3LqsHA8gMzDKoicRMvTf+5Kay
2OT2P0dlTMUR9YXYoBq/q8AJYbQ33l4CgTc/WPTsBmhfhvpo9v3t23sJDqy5gxEJJeDdbcsULore
W0ErJxEJyfqe5+GKm8RzBnQSZ+AMjvom9Xt7IJKN11QEGIBaiWQ7Rrk6NmPlI/z5KJ+tAEllDwg3
IHdA5F2fF6Z5y+p6h0LIdqw7TZfBQHqHHqfIhrEUG/TdTza/ccl4M0Q7HVN8BAufhe12fcbWHUFi
watMga4cYw5SdDeMPQJyDP1dk/r+zj5RIOevtednrYMz0Pbr0ajiIOixGKjOm0GurXFzZTTFGOWu
DT9SnkHgbShiKJ1p/YcoidJIR3719M1IuCikmXR0upMjtviynELQcCIDsFeZtF/By/Jb+eoQTX6I
8XqHpaRsRHjF318x2T31iYYa9jQfc8qwiJ6KFe0OVs/AJFJdYBNvO7zNH64RRhsehs7nmZj0ak77
j8rBsKeFPnWk3r2wtFZH1hxjFo5JbdBCps/t+PKhsnBrnUCfBfx9asvWNEkDJdAvTQfBl41DdekJ
ju1+BKl5jlSFRZO8nODbffCRTc5EUU1uwKBlGUHczqE3aokIGTGpJY/NsEE7TwNfAZN1Ob0PQQOA
+O8H4zrRLvkxTBQRnZ5GTuDQ0GWoNGvPswPVRzebdVcBe5fIjJj+w4ck3Mdelpla44YO7Sv6UOKN
n7In/kSuRWsT0TpiJeSR/oecknYkUFueryE5jy4MKLyR8MHS4r6beNUE0W6CnWKMIXGI/gMrm1Hm
Ury8QVsHtTx4QN1+LE2vSUNp9ptSseGFNOZc2EWECCHJYalj07zPz+byrnepnWe675+adQh8Ghhf
1/REFwep1NE3SUV/9goCR586ZoXb8q/r4EovsRC8f5NdZKCbUoqUA3tZrikyigx8w+VC4rvNfmn0
SdKc2vBvCv3jt2xyI7qQDMgb+txvkQqfnADeTjUV7OCaY7ZEFoOTM+VkXLgEQAMnEK5ikP72bDyi
9RuALCffN1PBZgZ1zb5OD1ta6KXUAEKPXASsGg0NLwcLoaZZB2OclARzFrgoYbMGwAx6t2jomIM7
dOtzBCjLU6mQlnK5ucdekKeX0JslXP5GphmPe/cJNM3Cc9b3lNU5qgCmQ8DD1hA0o35cHp7eX23M
TN18gOXet7DI7w62XvdtwwZN/h2/ue7GHXU5knOBm4TpoBS5/3hooN789ODsXNONHNu9YO8ThdS5
+lpvDqR1q4B9L/Q//FQD7rF3hXb+S7aI6Fx1KUeQjfkcmv+NWs0ieLkD5BEQAzO9NpAUwbjIKaEL
kbreyIFVuO+8/lNwSgkfQ3YA798ehqhj6uMez0aaovAlZ4chpVTgw7jdxBQZr/BjtY749PqES4xX
AV7IvsXzzBPNuf5WylFo8Q3PpCgZzO1pxFJEWTUkpEpIRdgwMIDesfv2kSgbgiaqE8L9/hMCQFWx
zgnc1g9qQ5PAomOOWnfX2NIX/589+4Pj0L34HbG6jlAnqnO+U0GJB5wsCkRP/yMgUiSuJiGSxwpD
dG8DugPFPrBlJkmO9UVLnNYMlnCyHL2QsrX63QB2+O1mhzBFUcXNooDYNoUarOmWt6/LRsYk9mdb
bD2OvieVMPUKlWyBxftyNuowzisDj9qTKtvBAJrq6fuEUoZaLYXMZ047pd5SAUc9eGOrBFuVfFN2
AbmcVrLZuoJKXGxEmODRhMrHIbaglRwtdCb2ZJTaeJey3UwrrhoNyEHy4/nqLhYOAR+pg8nSlTd2
hIsgdz9zQqaF+r11W9siCqiS8e339aSkwDiNQv+bylI4dhx7JaKbX2qwB+o8BBjzddAe+zlF5Rq5
8LdiQx+SU9bkZBiryKMzP0Bp7eTEmEFFekI+/oBHgw6poIAQNu5NhmVjeESBSilosEqO8KLEhp65
YWCy9/GgpABAuosbiG2gH0cN75dsvqwHEQ8WB2ncQ+t/xAOVRVPHJPYbO1/hSrovu8ynoEyerIRj
FN90g8Wl6ty1LUzpWzNF8FSjkb9n2SSONny0mHP2qKUEJ2vTN3PvOvMCgyE8KVcSjpz542qrSi34
2Dfh3CL4Mw32TyKF9cH/kBw06tf2hfBm9G+gsTIOflk2ufTwIEeDI4oWKfimArty2/VL8PWJ+JTQ
6DBK+5qZI5ggoIZxfzBYdfuVAHUqPy7dtxeGqisv/9AsN2YmCSCxyejQRKSNOxx5oZo7iC8fpqfj
IcC+TtjstMahvlEb+w+l+JGv2ZZeJOSkqqjm6DqGAzGkViCzOn8e9lwR8sAhZ7QQfs288DNHE/VQ
ZOx9qVt4A1T9F1A1qKa2g93EXFYfacuEMPIu9sSwo6/4baNdYu96Sse9mH2o22eAiZ1SLzY60tuu
tSRFILVvUawN/nD9PaiB2N2624uZs3dOVdaAS+jJyLKdXozrGWQtzMmg2i/rABTW/lj2ARuVV7Ob
AoT0/3TLhVX613uQx1T+9VBYrrmhBcWFb+5RnEciIGyFEW4xp1yfhv6HmJRK6o2ssXzAHZHP40l4
fAApVExt9Z3qF5GkXn/00arNDCMQqqN4iFlMZD/UBX5nrwB/A5Kr8csfGmOqCerAksGAwq3crDxN
2dhDlMTTOkEsldgJ5MnAetbRyTYeOdE4BVcdXxi9Cm2c4ri82CXQApFsZyKJU/NbAcrpH7LdqQaz
IWTjoDgwNNcFSGBT2m7BcierpIpbDy8X+doI4MNiYeFMzgrQVQSrrlU/Vf8wzoA1Q9OgXAg7+gi1
zej5bBa6uOeiEyWw0IN7Rvhww6v6R+/keLRhiNLR4O2NOMAKZbuustQ97Rv7lC+cPNEAQwCxSjGP
ps3zxAWxnx8ncbudQsYd4ebqnZ4ZbnCMAFGspPNXQ16heeLHjTLlN83s3HdPwUhfZsCpqe9l2pR2
SHoJyirhFNyBrQfMX7i0GXTKLIF1v8MhiH7ADXEOzUZCVz4Y4q2lZn8QCth33Xfi1fMZh2ju8Fy8
hrBgllx3uEDgisOBzCSviSQkHcjniSM6+YckJjH2y1w0LKbGSOl4Z8lhUzvp2dlHz3b7l/xSJi88
jbekD/9d+/QlmNrrxkK6A14o6WcbbbUQWiDEYgkD1RAcu6YxCQ39xlMElrhk3aiLPIfd/lGMglod
ng8Ljso8c/IaSLhU+zIweqgfinDSIwsF0/H0erxnE+1Sw/n5w+UUJLaNofqpop+/hXyAhxQ3Ir4v
LePQUH0C8dc5u9KYwgpuVGmjDk96r4iorjPoVK4bUslt5v7z/l0+gSUSjPWX9rZK0DQBSxnWtsVT
5nngGfFX4syTH8CkDNq0+kSAb0Um/JvNh4tuUMP5kKcAkCKN6HxT88fgUXmhrk1b9/NcATJo2ftT
C2ubqSrBILHNXgL7BEEmwwDUXToU7MLszTfJhkY/2OPsH40DaZaV/l3NQQIAlWrb9LbhrZjHwCq4
h5jpNXMqTh4swK5MSAv95lPRvifLcwYQ/ePLtD66rhIrxqjT7eslj08x8NsuF5M/+Rx5ADAUs+An
ckBWhOJ/eU/LXU1Li8r5XTKEEjdUGpnr9TcS+Pf1nKSLCC4GqzOrNIunqY0m8Aza38SdZmXDba/B
0Xwv8lRo2t8TW05FR8DRzUZFzrEUEuBrak7B8YeCti8afWBEN4hl70OCyg1FiErfSIab4k10obAb
Y7xeNyGwwQs3gMCwxh21chMNS7CzRfac3mG8LJsZD/q49SqMfoF24dKEm/9QUYrn+rIHJ760h65N
pj16yqk89riYx0VKUTDmDTUDomFk5WyPLSav+Vp//VRFmv9vs+2Kf8S5b/jEMohh1VCJYdOxXZDJ
AiP39PqR9jDvX7Ew0cyhH9dYqQqSaVqz4R6xI86+c+3u+elzHDps+4lTNaSPgX8xQIlR1Vpdinw7
uhrq2/O/Qv0+e8z1Kust9z8A8dX9G4DppI3LocwLPFTnQ9I/b7iHNUjHoYdL7MU95AFRN3grzrsE
wHrHwxlSSm7vTv1k5rAr+COwROKqLm/a84ll5tYachpXpDFwK/CDjgSPOPYLfLD/fHmnwL42NPcc
VwTnaL+DTlnRCs6IfvIbpLZ8hky0xqvSm4CszzzIrurEf6iCVrxjRefLznssrMBsiG9yJi/1IEk0
P2RDRTM5Ls1nF3/bihltNYu5Lk6MsVyINTZA2kXje3gyAeISTTs5VNhPOUG5Bm12fZjfibEyghJ0
U5yE+IrxYw5OYnwy735uuUdkI723gY/YOLky2z7NTQJpsZIoslSldnIIkKg/H60EtA==
`protect end_protected

