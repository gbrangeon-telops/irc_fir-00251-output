

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
E82wkdGPZb/+6GZoDi5HpckkoDtuL8TGRb/JCIEDYKunG0ehlHY7rWSAl7AxBVkDytYXn4VY0NY3
tD816aZ/Tg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aN+8nTYiRF19Ga2xgugxmmkjykOIKDSAJe8CuGlE1RsIGMA/TeZJn/LIOmkC0L4RXBBy5zkZr6mC
39gWvg+KhH324/pLiKCLqvJkIObctxdk1QghQFlwGyR5AgwumO5V8XR0wkFrGx5lcmF5I1Ic7QCL
4FCmeVtU3m0TggWFC7E=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aDXP5DZMSmAZ37R6bG0c2an3UXXBQ9f2UcCbZO9jybJiEbg3jaEsz9OP8BILMEuM2Gg6zqGospJo
IL0GjwnUkhmqiXNrUyuU2ZA9j5Qfpqi0cT39WDwUPJ8gireHKMW3Lk2XSOOhzAT2gL6kjlBz97a9
e5WZk5XJ4JpzHsyykVOoT9yBzVvTvBYrbMxRFsaT4GZ3NCp2/bL7FcAdHRGbG5cNEc+P//C3rwO8
4GNkm0wKVMVQq/2HclGOKJAykNBN7fGuG7zIF27nKqnI3IBVFzw28uEsxwVFMpLMQ1Amv9lQcw/X
S+F0+1sbjSvaH4de4WOv3cOUzYKQ/wzN6fSahQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c+SPO+b2cpVqItr9nAdAKH8LRjqZZjyv88QHjXDKD8kCd5SL0IXE6XqQ/EIjme3B6XJax0d6vBvr
92G/L1QzXOo8P82zgbpcUFM1hqtYFVROwwLTcIHV5QmMcqgWTv/CxjwYFY9l1w/ADUzzHakm7vO5
G+sQHpPE4aud4403sjY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T8GeY0or01NdwqMo6UKJMUTsmtP7APuN0oCIY7KzFu+PsK+FyNTk9rSPzJS4j6dAZuNV0qTymCiX
Xbb3asOZtqkbmx9Ts0TBudlU37PFSlhj9aboLv0+uBJsltC8lWgypATvI3dldUNiHT8HwKeBDDaM
ge1f8g9YSSRm9Jao06pgbL/b6i2WQcOEh+n+/rJDy+mhlYh4b7sJni6U+KkkIH+Nz+FTmo2KpEia
kiQmZaPY0KLlWtwgAmS9D9WXDnBy7lDRle2NygR7a23rjPwxBp5MqpWylPuquQQaCFWvB6BJrqSH
TxLzvd+PYmz3XQMRs1MJrzzaNEb2P8EXhMkKPA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12384)
`protect data_block
ZVyHCwlZVvjF2qiXC0gwNzPhwQQTA5KDSzBwcJNy0Q1dmaMulFYdkKqvJ5m/hs0ixAtWF8etGIGQ
333xsU0XwvSPC0Kzy80f11atL/ez9WhR7CZxZtYImxeixp/qBR0o44jeWaWjyqb9kzaSa0wD3J0c
29tPj+wIwmv+eUyOLe5y4jMvnE4T/ftlM72aJp4cKANUeI2i/FZ01vFyVLkBoNP6j52jdx8Rzwws
ETSJ39i685DTV2U9YanU4EqRI9HqdSb7EYSkJSToREppsXRmDeo27uwgtlbOYS7mZrX01oslhT6X
8rWB/sJ7OkBjI50zVb63iRWpESZ0ovNKm8AZWkgKEa+UaWMcK5rkrGo1lx85sHQB/4Y4G0PeO+Fp
SqW0DrnLITsK4CpOKvi3WO6KQv8MGWdbAfQm70c3FNSddGkstCtkQLLVRi2qa6VkvS6Tyr10v92i
XXsc3mnWwgzkGQKa6qoK01byT3fwdz1V12jOfsQvXFnZKYrh7EBjCCl2he4HCabATIubTAKPxjO6
Wn7KYF9VfTzV9IEcTtOFZtiodrVaY4mEsMTguIVq1Uhx4jphBgJRtliQbS9sozh18ZVWB5sK23Jr
+XFV2pHYfwAPi6iOXCpM5OdbcNTwCciq6kESq3NtYdqpW9TX6Na1aDag8PCRRfCfcRf+6mRH+NFz
b+9FBLTwx11AHe+oMAa0SPnrfqPmczdr9yM2lJe+wyk+VIJN7iRpubOwkFt2c90IBpbLSDnn41K9
Jqhqilr379/NtvcNOrPVrITsWwGOKlOe+CYTpfbwnTIDc+NPQjL6b/bbLrKqLugFw+yJa+yAIIO9
+AeJXLPKKBSUqkh0Uph8dfid6xE9d3vyLNghqbnQSN+qfe4zgiaYIacdiy0en4DfzUH3VwLxxq0E
7Slm5dNwNqe6VoDpqoIBZKPLcMmBx3eUTwCJILaflYI+IynuprO/dwe6dIBR21g5sz8hOX4lpPF+
qJ61oUkKeAUQO5Ujs3pYl7naKl+AEAYz10zJoMkfNyppJ+9gUZp/QogqPcHrSnCuV4dFy8P+I/Vv
rFU5qlBWLrCVzOYquGFRzIB73Xj/IplmtRgnleagcIcOdNKRJzOY4a2zdC+2NrQbCnkVMxfmw6rh
wOkb3jR7OaB+j7IJy49WgtWV9ErtdMldjZoIxnaVizTp0Vt30nwop9L4UlRH2GVdfyxrrO1SBf33
wYf2imDvCTiXYS1RgnzyV9njXTR/YCbtKA68Bhq74wwpZTsX78rgb29q6VH9OmG+6QBx1IVTZL3n
eOsClj0V8lE3LpLMlsa/EtHKeIyhVrcScl3gUjnCNEuFa8k5tPoaOwiv4PDURxxL81+nd+pIbPGZ
fUDn0iDGRLD5OYXgoCETOSkqJmcXfrEenyOX8SP61YITzb4ZM5SZzrzWcDsHGO1hu18XeO3TuW+V
9nxKtdZmdkrcLABJyxF7GzDeJ0uG2VNFIeGf7AstlrpFsb+ZisZKv73QTLCkVrmzrtCiS1HXo9In
tamKpqBbE/47JOtdsMZuJPsCmovC3L6sFlDSe0tRvzrgFyz6XpAnN1rLQ/ufTrpctllPNh96P63d
ZSrA+sNE4R/ofGOSmIWGVQOBpZojLTebrM075TNGQdZAwcjTaraLLjqdanIb27un9sV+FZbeqdd0
UgasjJbDwn9yTvnS8bStj5kXB5Mzu06HTCXwepwKlwHazKHwAKfa5FZfKrJTnyVcnY9DOy72xhDq
ARugl1Z+Z6kepEd/fRyCOukkutOQjiGsJQiJZ2V5z84rI6LRaCbXmOO8J+/jETH2uiyVR2SdK6fo
h/75Dc4lVuKqzXpHHksEZr+WW7OPkwOFRcfHjA0CeBN+HlYvTCRESgvek3f1CXgTSktepIf6ICq+
lgpajWrwHQhWalzSEAUJZ7LKD/mhJUj6qHf/U7NJ2KQ8JckZegZRnSyGPuKzLJVM94wBmXg5M4si
7232YJNOHy8UGeMH7dg4vY+K+WAVUtxgWIVd2bbbyRO2bboTxWME2BMAKa4eaIQQmOiSpema6F80
RMLNVLRNBirRwA/FjLdaQ7f8LVjjQstBkAbaTJUxk4uPRb2/wFFpuK+Dy3kgcr/fDzXfiTr8ie0R
3mi+Xiay6tBaERW9YTY9I2hhYuUjCVaSRCuPahR9t6a0k7MvFykIaBU3O8vgBQ5qCd/BvGTUJWLR
nW0tLHOFECxYr/bJS9jel+fPH11K2fN8dDIzliDzLy6MgBFcdmcmhs2YR5Tdf8DDRqpUpZfokDgk
nCt/HJd8KdIfpxkaDx9f/ViYGcg1HbTlRCtfD2asvC87fj3TktcpCYWII+GOkzMvpWM6mWDQ0y5/
PdvhFwITKU3DXkFW5wgB/1a9dD5JyxgwgZgdXngQkRx42anEGXCnqamJmD4OWC6kNF0MQXHDSax9
neSVfQjuAzD1iCctSYgSs59S5UeJjSugHMDqTR4Xec1N5OqOhdsdVSnmhsDTILGMnF4VjmNRcyA2
pZESLi+zyYHe6dcWG/h7OPbai1311r9Ax6mZcLdfqE9L3Hs0gB1SkuGitw5NmEZG1JZUCgAgPhT0
XsdTU87B1/OKH3wlydYlRgdOBkZBk4lnaA2Y9GriP9YUxhjif2zgKbnAn9W7WV/WXBD4qvdbb/aU
omdqdQHciNWX+qvr5j4WsRb0YMgv/9+B0xreosj5VUJCj/8All4us9zD5SPlwDfFcQ7hELGn+6wb
d/co3gJvZEFfd3G4xeqzqvsFxOazvJ7tap3DCWGI9VBnx78BqTBvYR/dogcqFlA7Vugg3dheH41R
I+AiIVMuxf6ajubhTEgTDZ5GxANVaw4h0qa3RmYPzNWLTJeAZ9QZNVUX/MkHcFzBKCrczstkuuT6
7XK/aSq5ChvFHKbjODma4ozqkoCCkr9BhLFuhxfYbLfGsqK8oMLXhy4HJ7MupeFregpAWV2RCHdt
bbLsaF8QJyLvL+LNJYBIT1HDZc+FBggstovEscyR9H6L/tNlo5FYWPCDXpzVhrCojzZ7FCcOPbJq
tcw+HivC7fbuCZpmL2BbUjSyUYV4kY+vWGjVUSRQKApRU2LXDx3J65/P/02ZOPQwZRY+9rxsM9xt
rClgs1jbR+XTTYqD9ykweouNL527CRxFxEv83tswtfK8lhCQfQQwqt/0TpbNiMopPLNFA/jzVI40
D6Kl4Guz5EsRFWHi4Wn7TxPGofMW9WNOssHQrQZNxJtBuVcddyASYf0lEIf3zDFbr9hsPxsOLbbc
Zso8voRm1eD94vJkBk/4rRgAzJw8MXA6TOPuJKbINNB8dRx1IcXwUmQbkadVBGBsIPi5B3oc3/7a
M9kMLCWByiCmFUFEy4zbtpgGGHSW0BNt3/RuYOnVOZYODclgWT9N0VidMsaSoH6clM8opXFlXEHR
sq4Yic8FaTsTGe3rO+giDDX7UbaSVPbk+Ha5+HpMn5ENz4teQKB+23Q2UHZzykO9qP78SSqkc5uI
p4jdt/kRcicuqFScTiyzxNaTHzRLxk1TdvMREb8AXYAMZRtm30BbRHYnvLzNMYnuP3iPEf60nfoG
071d1fSDkKddPrHPq47lAp3MK7LrRm1PSAh/VB/wNSdXZt7GMs8HlxWqJZmk46S6M7DtyXBrSmk1
YM5irC2fGVwv+q46ZqPhd5nufm+ptDQmMkYnk5Sx4Vfl0PYb99v8IrZvMKFCCTAZ1vk9cCgSlzIZ
PCWa5GRmkvYh2ZhVTk7OzwD3yHjIm67baUnPTyw9wSzvmJh/BDxEq8bdeojpF54VlDM2ki/zqvms
ToqDBVrtMWf+niIx82due+/wxActd9/nEb8MJ8bHCM3zhBjg6qTK2pWaKm7A5AxzbhREpGAcai8M
dQ7CI1SQlsAY+RVMOpnJkalrj/NNXzIn57kctPLVrytmCyLgNJXmSH/JmMSJlng5LLjH1vWRGlhL
Y1W77KT4OveFaswqcrkHDDaHZ0ovZIEvk8OtDetfYjDRU2Pdxl4MMoGLWzCkxaJgExm4ep79lDjR
sj8M2FPMNARy7Uqcgk567JQkOR584eRVj6sLmN8fc/lEwFe/i1BE6IPQBPZzMRbQbGZF26+zmQ2x
fWh0mdqPcfKaO8mDAScP0epPWLN6FSufdCZEuCqaDd2MIgKXDl3ZGT47/AsAnvJmg1yfIA+FMUDV
UXhbvKhemeiVA7J17fHtrvKCFmGoFh7qf2Eq9CncmUyP8HrCLHqSCsVGIbGhVcZpmVmsjIJBszFR
1YacdI78fN705tYzUfiEQSEJFzf0TbUAiX5zoOvUxJn65D0oLUF919htCPHDpHu48MVV0xPP1awC
KiXjM5igWwiZaryRVW+68U8wUHgXL1HhZRh/sZUIBCFFbxnjIFqATFLCIPqsP4+LvztFnUtwPVMY
oWOMHoUaajRv71hBmR+cTrk1WbPDkfz/XEq3AyqREg3TrgK/C/kfchl0+32mVCv4Ca4SMyS/8gKW
tlXxx7lpydzzlsv15RDcXFbwiuMkdqbZ2OEdyXVkyjFlCekLkv7XyHkVA8eASIPqpZtI0mmfVaSA
wexFexmWfqaIrp7cntfMEzRA+Ch6iHvrbGWvNcluQipWmeyXXkDA0drugomo7vb6ehBaaoLUHL/6
EEXoHgxQOzBAdIRwhn5osqALiPzCvqB8TfqDYKuhXQKl1FDUlls4KSA09euNZW8RWSIHY9BriwzZ
19osAAk5SNz65WqLKW7XfuIpFoArjoxAPR6Y75xv56bnTq1L/uSzuJUHzSs0v2JvuHNyMR2L4fdf
o1ebHrooJttnsd6a/7dDWec/EVsfQSaPMmRScimxLsUhrE7mfs/mzJMYiIPHCd8fCD1U3aO6e9gE
B3u2uqGF5NADBptOMims7zdc1LNMc7ADVb02+Wuskt9E+XI3epnExrY264pdZ2JUkgPcPsax+dUV
eLLYOrmXwr/64+5wIRpFkFecWexCseU5kqNbgjJHB7TBhCQbl+WvLzUL6ZtItfkMLffBUx0Evl3z
KO0UkOikQI8YcbEgu7SM8OpojNxlIl5ukWbbOHxtttJeQOVpXG08EhQix0vcYIzTrRwv2nLjeNp6
Ar7ZnIFOu5+2NbJMjr5RcrwX7Dzt5PhE4MNbx0MGVnMwzMDB/ElFBRgYdxybjhezx7XLgitsoa9u
RV1MboBjPw8j0V/R/4VwSqb3x+VBh8WcHMYySjmIsiRKcIV5fDuZM7QKiOgm9P5sa/T7+ZSTsWjq
zL42cVidKut3y+n6/R1BdDQKR0Qjwl3hnJVbyvLrWKnsqo9Nf4nWv50L9j1BP345CTkbOKE1l79T
p7UkzEtBtbZKNImQFVug7dI7gMt5KXZV5GMiB+x5gvHZP2dhhj4w+27oGi6yG7MOgBTiv9rbOzXK
Yovs4y1w1YuCEapnhjscHaVKChcY7US0osPPGfDck3NN7M8CL1CAj+TdUcQwQUOebaJp/ZRCsIc4
HjlP2XfArqX2WvQYYAArqaLhvuQXQdhPrgP+nudbAMYv8tAUtEOkedcmMiBuLszMdiO5qlh8y5jX
n1/6c5uESka3vKFHdXUlMyP11Gz1Ft3jYf9mmxmgojlPdtMAUSaazCO2bPz98P481zdEmdOTyLVV
/H6SCOZq/1ob55o79RE/nG4KrKcmKDyD9myzatdQSOfUMEAV95M2PbteP9i62W+InICkyKIjgAtL
KWKN+phzbxsawfWiM/vS09tR3+wguCfvCVjVO/YXVho7PsC4TlofvJVv0L5V2r4r3A7gqql/5nnM
aulRDgrmSlLb3veUB07dakDSDbHo54iHoNXtyHPNCDeFuv18ZzYg0xHWvrn5gsZTuipUho5QLgHp
+9uywhMmqJ1VZCb8uajkBbmNshtw6WxT9Nm6uY7lytHVsyqtJ4+ZQyIvztYebn28A3zhStJXH0u+
YjVICgbVZB7ArQL8/TI4EK05PI8a/URzsKs/OADaCVn100fBbGQx15Nosa0GVMGBlYrLqz1beTp1
p0xbafJ44EiXxPJousO/HB8UHd52pWHOvaD1VqrHbResFWThkBV5Ky8rlN0Q1oBZmGIlU3pqjxFt
7sVotUMXkEDOBzLYi9oRLc1Vsq3jB0suRi7RO1VlNuqe4iVlRg+spQDw4h0lthB1WcwUhE+tiRKH
r3Oj0vsmRS+22rVRj0daQDqeH6oreop7Qx2yfWfXAH0lkzFj+bA2RhLSMW3bSOMcAMYgq9iZzp19
z9zqthCoEP1HEsH+fTffGIIfsOlVwV28jX0AtP2idrKaWipfbMD60ttiGUabUR7/wuZGlnMnzP5w
8OYwwZWUZGBnKSVoYeMIpQ0JZkYPX8Yyzpt2wu9LWg4RbKx8xu277IAQiYG3mlAB3hz+bFubkT90
JE1sF204mglTBix1YNYPg7gXukdDMDwMe8UmFID+jnd8ODZUWAsjUJ/5Ot2XkY6rZwSx5X+EVD7F
q75pBls1QT04extEEZ+I8sU0u9BcKGuyNuo0vZksWprUpqCIxLdsjAgi3Z14Xj1jvjhRYoDBAzHG
f54o8AHVqjLvm6LH0sxYBO/rHKzaM8aRdz5cHspUMp7wuf0+fpPm1Q7Mi6Svq5kwx/kA5apW4sfG
9UF2LmnKlKnLYZiuo1ArNqinBoSPdNv9U/SZ/1uEliUl0OyFGm+NqMFcHrmTNS5Gy828aimYYmd7
Pm9BuLxqNLaWfAV95b9OCCpHgoEaonOJ7/gx5kcBYnXFgqXskaWSrvVHEgI4sdqfSK+mJy0VhnDE
X6lbYdcuxUs4XkxZQWYD3IvKn0XvpgORpjkLRya3cy7kUht028lgbdgWBUUjwAE5Zpig22za5itk
2Qx7vlEDDCWfbSaH39+555zXE8q8gTnzgnlwHb4aQl/5rXO7sJ+eya20GjGRb4QUy1k7fsclq8U1
PfuyxM/aSbFq5zdPapB4/+4O2S4jrOF+ryRy5QGQCr3Ze5aAOkalC0519lfRtUd9VEiwXM8SISfq
qDQBuPl6/u3udnGByENY47Fql7XSUG2oWRM+whBtiUn0Kj3PdwMBqIc1NeOGVO7g8XPeF7E5t2I+
jmIKuYDCw3TXBMgTx91ZwZNxhCmDK3Y/IIFIvgUOGTPE8UFZ0QzfNSu8oO0QD+2dyUcZvJUzKVI+
NwV/UKH3YNbQXbTBZgeTrNWSciZuPmXerguk6HnEvnuNnWyeXWRTlwcIlw94mDcpl1lm5hw//IJT
EetXe/9m/kBJcKmMB6qAsjUhk/s8bvKKwRf77MMLjBRDE1E+F5PZVRMBXi02qYGC0adistevn/go
ZAvlEZ01HJ5DZLWBhXq6tGQ1QjKn8KPCZxdNoEPxDUZyQaaovLKEi8/MY7nf9tn3IiFa4GduBq2D
x6+MorZVRSF6AAHlfDlfPgQLHpcJU/9866Vn1G5JKWNU3eaOFXan5uSQEobkiCNhKaNTKocpirJY
29MwDW+Mx94hCVsH0O4Jv/OW+X89Z+Qxbv8NcVCET9klzxkiXXMWyxx5qN4kzs3QVKv4GKZQ/qSA
P3ojb44wOy08Pzxs0xe/ioP5TjRhjyC4T/uR9/MJ5g4/51SJdw7w+XVUvzN/J9VKZtAehvo2or1a
5ECCy7UZYFa9mLgQ6GolI+rLSy0Az5FNyhkMnN/XQC3DtXaUZw052apYvRs4K6r95KO33QL72HdG
oLWbYMJvuhrcoo4lYPLaYnkwodYhMT/XKeFxQcMuCNELLvxQaKqTeyzH/VoRfS2Sjui+wUanndnq
FiqVU+tINAZWCJBdzPtcj5NCy1Qt6hlbGtMg6UaKKGZTmE1RYaVXBNVkxMZYQSbFo6cMu+M1hCM9
N23ZoXFLjRnzVk9z2nP4uGSfXjsT9744pmUSlesPHOhTr9zI2z6MQcV/crgmBgUywKsKQ6vZpj00
TIMnTOM9F4WxxZ62mdXX5NxGP9F39GCYwyabhsu0mCApLQC/4Sb1bRHiI1prYnkzuQixG/sAOEQT
iH3rq4/E6EYXjZdmHhzqisGDG1VkVtdx+9p0I6qa7uyOd+kE+WBEK+YxHoE9q/8h84VPr92crfkv
YIVo61NhDpT1W6EgWQM4tCeSJ+3O15vbjYaeyQkiprh6drq6jWKiK/hI54qptVAGneu0ny387C2b
gNHcUbi6KO4VsRegGWdIhBwUkBx4UbB83DZiF9Y74adZuNdV8nBLyQX04vS72+3aROR4uZBmq9aA
HmsnMpdj+xEjW/VDxa/fkTsMGX1oDDR/zdaXl9unBjtUVDzy5lYBYwZ1VDpBUBCs3b8N5lzNycVc
Dp2Ax0FdFJ+mp46l6f8AYQ5slelwAHLJ956Un0LWTSJAQE4/00r0I7dwo1YOOearii5zL/x73JS3
F/lZdgUOBO7hjUBfsMtjdpVJYvb0+gQ0xlSUvyfwzgrSYN9J8ThygtQOkS8k4dE9wcUoP6BZnFik
ALArtYz915ksOuTgsbp95p6gOsqPrxA2UhyCDY0F2NZseg364E35fFsrxt2I1X/rfX1zNroprsWA
Cd2llkmF/ExBYxQSe6/m4Ink8dqL3TKZ7ktQIUXBhECtMX8XQxsaryRBjt+GtG8kpzj+2QHQLn3K
4mRqk3pjUpQrZkH6F5Ws84x2CwJlW++OeocS2OhuoTJvVd6rtRbBDd7MMfyLy2P5BOSsRCqpCZK5
Bt65/cr3fSHWJ3TgVxM1ZdSEC7ijIZTB/j421tG7iO0BZ0Pmm5ZvFM7Niz8uK8mSw41eGKlsSPnH
j5ZlHMWaZC/q5DX5cbgYeOFqumZLV6uqVMYtlQ8yL5F6cbUoqhYBrFYIe4LZInXgVrRdQFxozn/m
KTwqsfGeG3xGaMbhW+7qjMSR0ddIloeuuzoVHwqETMyTpXcOsV4WRFr9rcA0zUTiNuzJ0hGlvi9H
57lJ4j97oqkNKOlcXQTcHyBeue1tjg6uZ7x+ENQfk5meWmmMFUE7lAxaI6CQneUdeNeyygVybRpt
bj6wO4Ypx6DyHtlSBoLzG1EUTNxteILlNgFAowi9R42hMdCILVxNcr2H4eGOUuDxr/hTmQeBhplR
OMnweNn8x8IfUotvpKKRUcRPxG8Tv1ADm22QYUOmrHAuI3JIf3Kcv741JcWHyXMeTDDk9kBD1a/i
Ilbzys0nJcN+Bp8sq6HyVu0FRTn8iGu5Sgw5QFxqCM5lr+nA3AzPUYmhOnmxAIvjuOvReJidLSub
p8nSR2VK9PhKrt4SHiK3kSc8Oc2Uyx8HyDfKnQIWgv190onRvoL8kr+ZQrvb2ZFZS9jClo2c+/7a
tMireDPFg60GSq6ZqUb41cPvHY7jgu7gFAK/Ua/W8fkz7FNeRPPLJA4r/ptEARV5mYcEL54bBKrb
9NTf+2evs0v79IVlMr+jZPFtl4DZXXXXV5LsB2UqELp4R3VCI8UF3qFj4eqaH3p44n0znZlvRyn3
QGpCOTGXfd5IqtwwUY32LIuPC4q/QemOx09FPLbzOYJil0GwMVQjQeHgirVa/j7Z7lNS9FOS460+
G3WTPWoObAu6436rcRwOed/9qSClr12wivsOs2uk1RTerz4M0rC7bngVgjDAj4uNgbHHFuV+jdv8
2Be9UJy5VwmArCyrHk4/Qlh6FUdRkzZisF4DAoeZUUlg9ClZkeMfUfpbnJ12emtU1VXQSXD9hUHq
+VnfJa35sa/uuTQ9/n9q0nCfTU3zDNOvUoLxhRsycr9BOB5AxEEgBoB9shXBtN7aSgHlr+Ue5mEN
AjKTLAMtSfC9+KwA0R8Th84k/g78O2ywYXAxsZlFaS2XKwoF+pCB3Ky6Pcve6tputZ/PRb6NHNE+
XI/0FpEuoQtGQaDlIKg3B5feXfII77lvlZRJ3JnKVHJqocQ20JbC2tpKAe906V8fCNF2oJqgDB5l
npyTFxNU4OzWpbJvQmyX+UgJ61EoRDg+V0K6BZq7XHuXkCcB4zKViztqNDLbHkvwM+C6yksxCDAj
JMK7gx1ckPjHwkKVDG6k8uj2DfLXh5N48KFqCyv65ckM7H2qOQY43LWMayvqMmCuPY8GKd4vy58W
jHwOXw7ZDhj7jCEsMGPhMyhV2YRbG5s0jOnLQN4nkYES0mHkVf6bhEq2PQFiQGdIDD5c13/OdTgD
1Tvln2fVsPPggFrIXxaiXSNJxVdjeIyjwJ4zFNJITo+AMskYv0fgz/OvtPK1aJwrFtm84f51psxr
JHJSkLFEaujyG694fTisQyFsTXlRmwPzwj2up2SKvbLiTQR2c2RubK3dDYLmkDT7X9QFMWfK13PI
fIBr2fwfjymaW0qDUQj6J9qVK5zfQADpYhsJFAhgpVvFzWHcgFGkXeNUlNdlkYQlV7w0Wi6WnOH0
QLyRsY3B5dA00Gn3SQA5OpJHcHUkNx3mw7Rampm2U3WPND/zBRAEbRabYxXybnAYHI9lgvJ2ZoBx
SQ34dGxtm7sfrvgJsNTpTmd0WzPYgrplHd6ZbJqFGXnQkk3Q9mJGcAf9Jngac3sDhLVNevubainU
x4YZNcbaSzvu78GHIpzffMLgO0LBGauYSYHZ5pdnQKQMQ/05QamCgAadqIC5l4pufWEylcmsUZ0i
dqtjvcufJLssl751ZRz0Bbo0qOul3ajlKlwiUMCXs0Ew46VZ1+LE8Nsp6Qwfn9oAuXM10ZW6R+ue
PQtM/RBfCWJUqfM6rBDG4T0d2u+ZUESU/Cizw8qBb2bX0w+o6MQ66Ch0JE8O8I3YVdFwy5KLUZNn
Vnstm7/sem3oashdKnsE6/+kO3LO/BwIkcStT+LLkDpOrBQmRAJ7oVuuJ1629G8Tt8A5INiGTWJ4
fQV/hy6DgkJbeB+9GMaWXjxMHYfRVFPyj01ZXMYfKlv7dZmsWXYsVUh5mdrd98j2IzXmUazfH+Oj
xppYuayifrmlC8v4Xlb3lJtO/zcK0uX3qd8YSt4BSU374HaMQu5NEq1quKslKPVkgwxtvr6jDtGC
3VI4Bts8blmiHTKfHj+nr3rosww2I5OSascMWPi2P1XVqFy4kSLx5tsXT2E2JVjswPFJN2inbO44
YwxDyLnwOLXa32+Z+/0AuJeZzIj96JzNy1tg10wTzdqwEK84lHUJjzrYr5m4lnYNbsvsn9dFFa8N
kk9SdWLzqRE9W5VJgdB6Ti5ioS1S1a3lv/vm437V2ZOd/yLbrhtZ+vhG4CFqXMBk3J2ogonn6/V5
TdLKZmUX55wPGY/TtaU3BiEyJ1K9ctubLhhADyutwNtJRXZaWRvXdaDr9xsugC/BYO2hUPOE724L
CS/K85Aj16zSFuZVBqUxSqhd4Ge2bLrEPscsf7Mhs2EEizeheHigV5s5HWMh1Mbpio+fwsyZwntA
Hn8fUP4zcKZC1o86CphNYa186mDAnhvC+UFIQg3kEdj/SOcQqITLb3iduRo2ohdH1drQwVwr+dfs
ZamZCud+G+0WaCZtQT4tLE+8IkT9dOe7USMHvEFym/9yE+t5pOErQSnmRhmPTvqCJolDZD3KqbXy
vKifNJUdkUeWCF5+DcMSumuyJzNl8ApBre3Q47B1UszuowZfPG/8/cOu80INunSAZ7Tddj2wGQCC
VNjtBjjEKPBHzyVfPnIk381cXgp8iQYlYn/60bL2ezADYnHbZ6vI1xaXHbSwEHm9ajRvqfh5MtwB
HsPZd4ijZOIks/ZZ73oWVeQRzXPi2ooMHUsFn78tUtcnpj9WcHcOR3kFPWFGuyMeyYWzHg38NeyA
GznHcoV0LCDT5mOHfNo9oO9QJiR5SOTIHpG9KUqUzpyK89Iu5UAu09aXBH7Of8TcoJTip+FHfIed
R0AyMJsy2ATKFeGquTBSM2MzmIuqKgq/IuZSCCfM0igzGRknjF255OB++E0em+3OcPbkNvVphOUa
8+b4I0EM1ZC+KYYiPF0eJwz/nDuC2WGQMt4Sf8c3om8nxWktOjb3rMfPhD7QVrDoHTHMUTICd8XL
54oGqBaT2WBM+pQW0XalwrP6p+lCl2Mm58iIuMZ/Qu7BjCIeQG+x6DZnnvDNvpsS0oDGlguyVEhj
SfDOsf91TYUwy4nBB7x/D0HnHkZf0ZGIcbmdRqOKXU8uoqVxIxgfPcfzJY8Dq0gyStoLMrb52Ze8
kMrOVKfwnbfTFR+aJMW3DZM78VsgigpDqIYfDbb52Nv5ONfaNFwBL/o25UTwa+0NCznAmO0gz1t6
3SKJ6ZbW7wZ5EFz+Sjmi8KgdmUDBDNY4MnUl82wd2Drnv4sVLQXb6wWjru2rh90NgucYdH+tJS6E
hI0BdbAyaVubL4Ry3cun7wqApIsu8B+3cTx73ccEhIgRkas5EjIwa0TtxkuMmf6ii3ajmVBaR4tu
PioEtiqFhX3qwQte8UpfesKwVz5yW2SJHPho1lz3FsRVJy9Fvj+JqnB2e31MxOOwtGbDZQkkL6+V
AapSa4W4ivxie0Cc9SnVZKVJYKjwkJdlDq6l3nCTiqYMKkkdAlZBrQL1FGvNNPSYKmYO+FdjsCHE
qLNKFIFSKTydbxILkiZMlJWrBYoSDl1ebZze62UhPA8GaThYCkSTgYISTJtZcSGs5DdkQgXYvzyA
V1dXP9YdIkLZ8A1b/h0ONT7YFGYqPJogNc69/evczm76TpfR0rKQHYB676kV7bQLv36Zf1u6IRDQ
ciSUZdWErL5Nw+o8ZPOXx1clO4be2tJXd0nb35M/wNCpws03dvUs7BGHaX2ozcVgflGf5aVcfnGv
TZ+aprBRdSF5Oq2BSdj+bw7mXZdOJ1/WVa75Bw2SHVjepaJHbulOHG4x9c4EsaUUAcYz1nTG+kOU
mWWvi905ADiPquO2yJZNEe6HNiJdVnz5yfjPhRcwC/0siymdbxeROO1I00psqr132xsI+i771kJa
STuy1y3z2KmrjuBfPfyTa/KdlD1hYmwqeszSBp6qF700dwfUIcGwbkS9U2D6DJ7wFT8dWYDsFa1I
Tt7fiWIDhAi/pRkVt+/Mb7u3Ntmno6VR2THzVujxHgr+WyLgD4MhxuCdZKGP0w01LTYLo2/YpEQY
GVEC9zLj3JQxOflZ26leZWIePbNz7VqTko1RzWvG+C7+670eVaW/y6115c/x9c+It9ETuVt9MkDx
8KGurcozFvGl1bwMzLManO31hFbWQRBkNuL/gc+MA/63U1LOuDiCOOPjZadAodcqO9/MNSh+tOmO
j1clwvXcd4RlvwDPZtlfyeMnw8XN6AKzzdcSMVE3CYuN3domnXNM1ZQyd1BiVP7HVlmUVGCcHnKu
R90rd/5KeXsZaha1RgQhT+R71OZOtPTL3/gj0W1fYXOR0nrqgNawwI5XLzA0jYjOW/rC4ftpg/sH
Xx/Jr2NpYIpKdfAgDI+iLg6WEHQjjMlB/xi458IBm6bKgrbEO/d0wrCArueGZ44ZOtbOLAtiUKem
jMEuwkagKNX0i/ep2MKY7djvZX1hWqBunrhX8iPOevKupw5JxLVCgr4v/KEZlIgAL+mAEbzUdy5v
T0BwlRd8Z+JB2Nuouya59y6NfwYW1ohU3zF7s1uzovbGxWILu6zcBeY7rLboY5MvxQJnSQ29LcqC
zuScJEHj9/LSZQDXTAZ8/p+er8Bjb1N6Tmd5c2dGYDmdr83LIqqyaUMTeCGYAlohtsV+jPOW6xjb
Agwi5yZFGSjRF/u86AXA9Vu6kPUqBAcyC5CrA1ikTMNqlJza38AwOQXVBzpKh875Rdz92TWqus0u
UoBVrnFG57pOmVVty8vCGK6zsQT7eKX/+gcQoVrVbDE8w4O/RNdxFTaRB0uovRATN3elAHwCKZET
MoO+uLrS8JJ4WiJxBGA27gbqtvgFoSqAOsGi8AiAz38Kjvu3AyparQORarZiHl2JpIXLuVJc6dYu
nybeKlSjLnXzhSaUb8ZZYdiyQe50imofyoOqfPC2fuL5oAA2azRpgzOoHEMUnAGEr6VQvx2UN+EH
FnAInn0cxJIozsK9D4EjbqD4gLfC8Ot5ZvxywL3M+J9rnZmRFe2KSXHtlIJShLedUNBP8hmfkgE6
NpRgqgCQVabF4oIr0c5UgfGMM0lwh5zM17XRXbSVs7p/6eB6pw4D6DDRK3oXnqQda+f7DluExP06
7aHfbBHhFyXDeW9Fx92jeeRgQ+ev7UPKVllj4lrDe/jK0mHoCOdwNqcEn7iZrTaNuT/qKYOIyasw
qs9Yp6+sPLfx35jj+uywGsgm9cMFwHV+htSr4T8c2tnBzwjTGgysI1W9pAP/BTIXfqR43h2Gi53E
qikIRCOEznxrDCRVVSYbjtXhbsBMjLVj9ak++9zu3+zWiUSLk5vDl1yS5V4n/lKA/4EM/YfUX02G
gMjnu5KZ+9CD2IA0VZdjc2ahDY4aOFY6B8WwSCP0Mp5oV+qqXl2aCGPHykQcxrG+WJn0MMORtAZY
hw2gcLv5mGbyfOzE4/Hm166OgtsREFTpKrr1CtSv6DiKgrfpVvchWefaHKmT7PtzWJ8XvqrQxPNr
mw1pL9Bm2GpbGyL1eKCrSvFxjB0KIu75j5BHQeibNkg0FUK6KY3MkqgSWq6Eu1h++6fRMh+1KVae
/pbR5WxUn3wC7QlVCE8bp5tc7NAbqSM+H8bipG54/86BrJxTt0AUpADyhKFuWPOX0AApsJEuXAvJ
gqvZLuMo3O0oZKa+e7xl5nIzow6M/a/1UPp3YOgI8sv3x/zNGO+RwWOJUYWKjwoudQFycnUK1LIY
Lg46bBaHx7vT7ommWujeiYbQyy6ABgrjtuhLwKtOleQKOrScLcyfBxIyqhjP5tXTYp0Nb0IGxrno
FuNzSme+/XF3qDr2wZXWro8BUGgOM1dY9+U6OnSSy5aWCC/K0Tc/uLdEAt0JTHaSMz3JOppk4yff
2KUjgdrWr6Y7M9RyM3jwQ9913atOCEY8TgHcdypwORvq+MKMo/8x7EkbW5WVwGpfhWSgco1BimjO
qcKzgrX3HusSTaFRZ+tKeu/6JDv21d4e5uZtisirFovfVuXwPg/kMP5aDZM7Z78RROQ7yXMpecvl
L3aMQfHb/Ip86yhjx/e0ES15tf2sVgDORsSZk7CbXEXd3kwJ2vHw2OgdgEGwsF8FyTjxHNSME1bx
iKsq3CSC11WYfma7esr1n+XJJ+J5ms6MSHGmJchaK6KKG6nuosqFRRn1lO0kKgRgEodtxpNixX/D
Uqf11nPyGjjqAJPSpnvh/UHw1lG0YR+7OHzYBwQhJEOqiBrFnuFXtDtnLPwbbe0cOg61pl9RGcy7
5QX5qOsKe4owIkQTAhos5unuxs1BFR2AsyY4SSYIVIT4aq2CtYE4feskLSTDFAuzru+J5r7bXEB+
QggqqqizqZouOoMVC6K3kd4XVCNtTbmMRRjmgbHdoEqj+vE/STf6/4UAdiDfM2Ou8A/JXEY3FpHP
c3Rc0PUAFz/4/TRe9OK+okF3orQ+y9E8qvqEror57yaQGa1CYEhndNM6j08TRrHw4ebbb4NFQwls
wviB2QgI3GHtWtHcTxDuYjlcM+bOu4e2nkwVik2tYMEFEdc/E6U22GEyRE4cfClQ6Bg8mVDoSGrr
7kaxdp7x3145oAyiDXwMQVfvzhXpQ0pDWfE/yhw2LHi2uAR4zHCaVwGcOTmCKawtS+Sq0x3YlhQ3
cfgsQNz0XnfllZycGuCXbeKa+aHJ00B8tDCxiA0/0szj4owFZ1ZQL92FeA+h0TGu0WNrHhXj/IBy
DsXtKTdo3ntcWYBDQx0JWy39680XALZ1CmimSav46pIbVG6BlMj0fhKoF67rZNz3XINLl3BM7OwQ
iTFDTic5wYl5XPQGp4KdEk4cfhyqAJjjwKl6IObBFM7mbfjMlBGRDDtRKfu2twDeiNuir7gDVUMp
S0OqyWfgpSDWCjk74dIT0WzNiUKOHWCj1lCs1lTEGQiSlm7xITYGz/bauD5qzgywNcBJ+fXxqZbr
qhyU3EQTPHrHlgsJX50g2FBRJXMaXlQFuBDQzmzTSJyqzhVr/7UivN/miAAZoGJ/M5BYqyQb2BVD
9pbC6SIX9zfrLwUkP6JpbTnZrP7+z4emDSjPa7hZIF/bPQ4l6JXfXvW5HJV4nN6YKJKSKnqDFY8T
/TDvTVuy2BeJhL7GHeKvCRv9YONx9N95n+HzhDiSQbDhJTIXoMmYHQpdFWJ+//Ze9nXg58ykmRqG
vRufw6Sw02JBkKXkrPs1d4ArAgdFPJSS1lekoVBs/LypWG2hVienkx5bokSNOtfuHBzv0sA3wF64
trU5p8rQKgmMDkAQwG5BDpwnHP8fnKFOxFgyZukd6TcPFQmkDthAuWo9/81uEWq+wE5Pp1AE6ihY
CM2XaL+qGUB8p0VBOj5JXhGMYc5V2Y4lm9x8+2wi2JFqVS3x5z+rkNw+NDlh9WtA4IqHpUwmdiqT
1dhiMBCyg3mphP5WHzAM/JQnpQoymVQoq2HaB1eIhcXtFExJHlP/wQBCVpVAdZS+gCxqcHMRv6fw
uyne/oXCYLjLo4031W65TqMFAzG962G3wnkbm5E3tonTmzmDUQlBiuoLCCh5KrVa0rWCyDglfq+u
S0AOQNkUwjUGD6RQxIUd
`protect end_protected

