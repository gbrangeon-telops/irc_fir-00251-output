

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7Rd+JJS6BPhm3C8uEMSjtB2IOpOZImN8ABL10O7dB2/wknTrPPVnggIUugEe0Un6rsHScVa0yw8
WbsjeU4skQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bancDuzOXzE/C1Vj5QpW3wyih2C6ymZ1vv70urQ985WeT2kXc7KQyN00fbod+1ycgrcEzdZs+OxF
/cQLUqqV1PAWyHyEqXlxABFUHjs/nxBl/f/B9V0jlBhAzKCCHBVtW+DFv8KpHE75Z2lg+r4JTjg7
zQiXYHxUisemJqUJdhA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rZMEEzwWFXOuo5snJgtfZx9Urf7eZRBCxLhuSc3DgaT16zNB/FC6Qo2PLk9pQbhTwkt+6VFrAqaq
rIuJ+6NqrQaj6tzRnuILLQxRIcZaZnlaNGPM0QELT1/pgSpbDRVs/w+jfcFf6hDgLWdb7+lF2lZt
EzdkUS2z3RzGxMw0dEl0kPzX4BrObwXWpUb1u4DD6JMZb6O50zBS5jLIs04xzSPqxA3PuLRWpuc8
zAMmWK1PCPqsF6JmUA+ToDlUTA4DP+Qb/r/OItKXADHbpGUiJXq85NgUc8TOMYazRmcSDk09joNa
rvnt13K7ONnKnXu7DU1cLEZpB6zC/Q33/JmxrA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fSUvPGwGSOzh5U1OjbBgxWaXchd+ErSm3+d+gvsNPzEzvrhBDlsbz7cjXesFumQgP32hemPRlsUr
lFspe8TkimNAMoMtRIt9Rpr9MJxdvSAJ2AckK92TaQKYGICYWnAAwRZdM4hFhKQynq8onwVPOItS
8G6qhIBnq17qx8rO48o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MVMseSXR8Gidb6hUpBeQo+a3Ho0qfbo2cQ4XmaaPwOf5p+bpngyRNVgFStTGlS9V1Gq9sxZR8m59
KVYbqvyTG1F7VywlVWjcCzm53JiHqc7770pyh1TFlHFmlBkxaKOZI17/BbAJVPtrgC1AFUgqJIKl
KWFzGNfBnaqYhwSBpkZVKTp2N/RCKh6/dORV7jPLmH1kXSt5iI647oKA/xzmV2IPvCjRau9wfIMP
3BcMw9SliL4YOeA2gPuyEVJdJ+sinBGqyYpGCshGE4syCgACrJDHcCC8bST8+Ee2RwROkSw85PvD
RmNqdRJR8yBkuN8MggDeHwsPe2oFAGN33DaQEA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`protect data_block
WXCKhBsPj9Y6XcBDfqwZToZ3iGDIK1uE5lV6OSYJaWWNbF1ZazneXJ7QRIbKX341d8I9Tt1aHgr0
HScr8pFC9M1nCCAJYm8EZmyUr1ENHhOo4jrH5lo0xKdOOrbrG9J/fMJ6vulAJrsPlig4CcsQFaDo
xCh6GIf+NGewhlcHao6xNlCKKCnYwdWYz4DqChw8ARv5DBh+3XGPOh7E6JMREI1cLFSRQKuLp9uY
Qroe+TzpWK0xg72YU7JbYPjWZCdDVITAgmKu32cJBZsVnY4aOydz06zu9oMgvnMcaMsV4P0lyz3j
0gHn3vIt+HicXoZPN915Gionb2a1ayZ5FeteOyckdQUlN5YTE7Pv9jI/cSqvKtw1JK8preGJwuEY
AQDTFTdwjaznR3jLWm4sDiltYiACrPOK0j+C1vHcdIdsroIYJXxkPOVpUFEsSSiAgeA7EVXpuEDh
3HiM5NXYgxCLaHP3nbujDcz4YrmOi4HM3Ro3E7TnxHqvpdZZ1cIT8NkyqbSse582VdMfoRuEQvle
Zdi15DuPUnxgwW2F5kprTUUznj8yRBcxOl7OkPdGZHun6r0QuzVftaSzNokphZ15cnshB/ACKqOk
SdFBo34VD93rssBWdFfPZz8tcp95xg4AlGfiu0b3y9f+QCXKmkaTKOX0ns+yYcoqMXEUgOzE93QT
K2VkAhCU9GngD6g/41Itf4jAAqBk0M43h2WG3ULC+5KZbBpqXZlZ0miJuq2C3iQsbjfNEjpmS7E/
55Il+q3zZ0uecWq5+8VOCpgj5zy+PSX5znmuLkhGGhxSLPKlpEDbZB3/TrzT8bEdIuKlxPFwQqmA
Kl0VjUhSUwn7NG+mT+4/BUa0fl4JXRhP8SRVeHsUSk4QyvadOWWmMqWvJV/c+JRs1qeL9UVrapiM
59KT5stbSjFXtu/JoFsYZy9KFFeDKAfW9+EAjOTT5IZJlv+EYmPJa2Qq/ZRwnehxKnEYnbFtdshE
8p8/c9pxygqYAEcbu/6zVBbGjBgHpwc8KSQJg5VUqffAPK9Q9Osr8oyzZuC1DWkNfR0M+Zs2Ufwc
cnflZ9VxdvYU1lUlxlnnDjaKQ4H9IYFEsc9SKGA7LEORnnJwXusddaEH1WziEc6sMN1UtCJ8Fus1
94CQkm6grEo5MIBazrhQw4q9kdHY7Or+e+FYV0B7r6azZ/g5cB6wTlL2QDcwaq3sw7NsEsLlMLSz
uInNysryV4HW1ovQlxinq8+OxbfT5nrwW1aILPB0r02mG0JqDcPIeL1TBKBEg81z/HGKzMQFwuXT
+vSmT6uVf0LGYx2LWb4mNb+2n7uSH14o8qk4N3yKwB7xtLWEU9Vowc9b7/btJtuZao2HYCGcteX6
SUWPRwuJKBRwVuVQwDu819bHkV3Psu3Manp7ken8Jc4PAz0rNBiSdp1ZK57CYpitoXvZtOprITDV
JYS7mxwjC9i6aE3dKm7tYMfkVIhBT7bpn52+25dtw3nvdpvcvTYf9x4Z5FNHtbEqGww1xH+0w9z+
MQcPJVcngR3qNgm06FIyM++hqy9UQclKmHwQWwoFXIfUK3b6HjGIjCEHpnOk1k/q/e0To3DDl8Hr
8a6dSdEhl4uieNGgCgwlLqSEy8/YvfaS5lFRAbQ2k979nozj44BXGh8LCFWuya4bOxTpEYGdx5Fv
cuEXXWp8o9bGWNvJJLXr81FMPUsHdkgPCjCbSXUeAJgzig7Ff8iB0pCgRRPsLPNdoCKfK+G8YrbK
hc2Q/pC26I0tC4YPf8DxlrS3pcAaOysNBYbI02WsnvAg7ICxPAygg0R/7qtR0WsmNrab9cCLLdZj
TZQv8b6Q9VsJWqDqxC3Cma/g4mWd3jdXtES5TgNEqZzwXF0N/BYIfiWgaEZ4ygkEl2T114hLHDXz
wmq7MCVF1QyDT97lmz5wIIgmuB/0Z4O7e4znqWkaraGa+Ce1Keg4wBw9tyCfczgejRPCkgWxmGnP
zADT57NI2Nh1H8v5brCsuF3v1NcyLVcL27xBn5Em6atv5Q/p7vQN98KwEQiCcpGEnvUl6IdKUjjY
/01/EY/Ikv7sVxKpx3XE0zYmxUSiHGCgnPUo9CZeuxelzOJHXBQE1A7OT5MAV07Mp6jTKB76lhZZ
W34dssljziL6mrUwKlV48Wvs9R6qdpcKo0WsMM0uRUBRbnEDugTVqnhYW0gHCM/JUR22kdGdeIhJ
WqF8qGIyH1DFuQXJ1pc+iUgX16yDSZlRtzBWZ17wBEl8PgNJM+XTlX7KoEtoL6KrIpdYw7TK5Lki
ZWECfa8kiHCRfKTkGjsQ5nO1xkKiK0JNrkZ8cM4yM3vaVOIKcd4aSKvWrUPZPPXJZM+pITnfD/pB
CvNE4NfUihWB/vfK9l4qPmgjbElLoCGPyKr6U9y8F/qBz0sK8jhO58Q7vD1vjQpPSlvG01ic1Wg8
Xa0iGZ+C8Rj+wRpY1IXT9RcRwUI9hQ8IHNTtxmW5+tjmesui8qKGCVLHJrn2Iz/K1SGa0U84b9yK
/Mvja6aK+YnOUNjz8Un4OP/EQfYdvjqtT7NwfaMIoromNqeYirpIs4SQ8W3W84CpLsJUSH9o1jhw
is1/iF6G8ev/Sk9JKdsvHIECTclJk5yvCWZw61yJAxkyGzkhVpCcovWsx/TUwr/bSVmxbibgKCAI
9pLpzFd03a8NSjjhjp7+bw4ZV8zj0BizOohBTO+ubYO8OzMtxtEoakfN73l30/t/C5Kcylsn1Sjs
Q3xuLKzZn3npM1oXNGM5XgPyyVnQk0r+6MLgi0SPDkXddE5GS1l8qCJIWOckNl8qyemkPBg1ulxa
pGuh5WtdojxEnV/7Au2pMrQcKX+c+0OLSbAX6KmMs37zZ7OUbjWOIIvPE82IlCvO+lgOMNZtiM+d
qFxfd27leB9t0U4MA39AoIatBzwACpbPoyU8KpeWD+smPDBNROx8/42lA3gL+csDQL5DQjgIhJ8S
nYUJyO69ohDcxxQGuHa1K2XeiQUQzhzHAISe8VljMfBKZujAHE9RATYKXlFwiibYrJ5wgjuH4se4
gGcLDewh56hZsaJyTiZOILs3tbwf6GaJrjOJAXi9VKWixqVanFOyB13tymGy0icW2IWnej6fWmpM
Ofo+gXFGaRVpcs645qqy8TQQv4WX2GVzAD1xi6RNFPigFy8jRreb8P9QcbVBJZIxBvZARNSUhI1X
+HlArQ2rPrHrG1OmXWtWZJFncUVpxI1Qq1Dp0x46UJSYlkQ+QNUTrvq+GCZGUaqr0YyTNY1rUlaN
aCHD4ztlCAv4H8OyEBuwMU8pHWsiafZva0oH9+VCEYAjwHcywC5IgoI74wp4BP4fz2V4zmhh+qdJ
f8hZRmAKu422NPAJ6XSPn9IyNhi7Soe67R7Vy+jrgh/BfZO8rvtEyO+u/Y9EaClb50rC+W2gfWc6
7GOw5XQeXjd4w/rSneIEHsV2E1ibccrOJquv9iID8I81URqnHHL/NpGVqUYSzdeIuSKtnYfvSZ3M
6VUpMnerEMVhHDTNK0qyI6c9aW6LPfcR99QNJ33ZeM8UKxnVF7O8m3XOSVkHvBcqGpdFuR7IBwLj
N1FUZfRM2NjWBNigDyx2j3DnC2p8iKNJ/bZ70h1ur0QobmEuHK1DZcPi7UIpe0uop3Xb7Ml+hu1x
6RXMDlb/UH61WbrdbxyN5UZtBeX9B4uomAseM2gY7r+QYdR8VLBRiw0MhV/NOkCFg8JYIGa5TX2+
51qu4R015e1HOh/RKRHfCa7k6CoouSQFIAwpsj0210A9kVnjYSjorcbxxn7dkvyoMWw/szA/M07X
J/MI2efe7P833R1jvUXz2fJhPqu/nf1Bc+1VAZUaZm69muPeFIKHzcvQeR294zKpLCPVaxklhon/
RevsxKgGEoTOm7ZFrwkXBBrWfKqEgi8wT5YgTrTXwiSuTWRgF2t4aayEP5mdAI/Vsr+lasPS2Lve
msYnDCefIpeM8gyXjNhD1zpM2r6ajeh5GWPqaQdVHm03WeEO096EL32KCIeKu9uu4xktkj/sa6K2
gvKnxuLozYCmbLLrCzH+uBpJCzVlzmoITTddyw6PP67HYZ6T9cHVpr0lhlZsCp6Kn5k5AdGMW0xe
sZl2E9Xz9T4WNkZEspucyPO49WaEis0GLUiagg9hQAdwI/J5cP4g3Zty+Fmkzx+HM/GwJSas8gkE
iT9dowZAYImfm79NYHqwg5jJU83TG4DM6WaBW68QyPtSyzjo2YKrT/o/TP48Kguw0kloNTFf//Ue
JGl6iNTF5zf4CLySyOO7+dLagaoXUbfVUjdvxuZOoxwaa74io5pt29R6F8rMMtSOsXY2A4g9IyBS
XJOJJNkHkbHR6Em+s0vu1Avt7wnrNr+0a5r/hTIkp6qup8u1FZLUPLGnGxnITthBUT5C9lF+IQBX
/r3QL9mB8llJgbu5OU70Awm+DefPU23AYMApOC2MGn5WGmGTyOYRr1aP+/V1XRtQTNMY9bYVtxmd
9FKUhBM9qQRFwa2PTfrAgRbklDKN4LSdmM+a4tU+F9REi0nhcm5XojXpQndbfidjO4XiAc5gIuyb
Xjw/5s+WlWYVKMzqOQ/vqbexnDBwpZ4STqCqEdbV9c2egmMMK++BOIUp75RQc0N4p5Boj6+D5QPW
Fy5ggl4cBBznxfwXryWPJV43/shOHhvigToRB9LOHpn892TP4LTPc33R75iZQLYV42TlW0FR1wVx
3JgJvl/9LxGNnkftH0P7E6JzFZrXLb067rPjMZX8mTqPUlH67peqi3b2IXtm+BpiXttuN9j2zrjR
uO7te8QCia4JDzxhvRi7TLqt2I2qIfKDbke9QMYGZwQ/EgOj/Tk3g5SP/YsyUKt5gT8Yn+irojE0
9OEqb6mVCbVRMfuow0MNNvprRxIVx14y6UMw8BWLO2aK/HEA110vxSBOIDwyw3dTWq6hF4PJVCKx
AwWwFWChmBQUxAgfqKjkvwYpehgFp+NvZm4SmzjebS14dJhO6iHMq2AwN2SArT91AsRs8+Dn5nFk
RyJsQa2tZMjeMvcFJqYD3TjM1Kb5Fk0+s5eEWNWQHk9t0nbG+wLAS4KAdlfU1I3Dtps1+fmYapPE
uSKj34IEDPZENJs/acuynN3FbiEqgapBPo+0ZGBXckOtO/2njSQmZs4n2/Qgj5231Osa2U9yvR+J
hoAApmn2FYKvEQreZvwWtdpMFOvjn4Be0TSbF2Csyor8AhoLV8uIx0WfuJawE5rtvgohxtNPoWXB
2npe4V0FSvp2olFEDe7lC+DAD8ajgtv27Szqhiw56nQ7HYTpiEVh7kMw4AnFc8iQy2haf09uYqwb
tEni/KYb4ujUEt9FhQqsJlYV6luOVwzL1k3gyEG1MDBdY8q1B+4Pdhmaey/Hjdd5Kdc14KBmrXDl
47++e5x0lfwgxEv3MdYNi3Pb7YvadK8mKgJaXhSQD2uV8K8Cxv4WQaAZ4WYwq5YFJQqno2fwZRrG
dweqiTFvMbcnTC4t3vYO1yr4xZutOSbkMvJ96jH79taLjfQX/VcGXkHO9OCgHaxhO383RHIqaGah
6IkElqsMu/FhNjxTskQrQco/dv6/dqb/d31456+Mq926Rl5B1fxGRgFdk30JjeCj12l6fRlyG/GL
M9Voz8XqIXwnUQckvueuqsles1cf83uM73eWwtStUc7EGJt1Ksf123w++BBGCCtLWUgH5d7b3KFy
zsbf18T7HVa4/YysqYKHi+T2XSNCoF0ahSo+fJ19GoBrKbBOnUS9lbzyDJqsBeU8AnzGU8+pOCcc
vnbOzLYM+bF5jYKk7jXwk0io5aHkuggIMRXPMv9l0K8i6II918aE/RitbmAQw/xh0pCE/SxOC60U
JbZsLVveqnryYTDcVBEShQehlCjMD5iESUt0S8XaAhAjRLKPEeIXfGfCZzQJZl9g1ya7pH2C0Kbx
iSY2gmLSx4TeyJ8QTUeR57BtvdIUJdkZWVIowGHQJYsqnGd7gX/Oh8+VciHpEqGu5qvIx2pd8GAr
swtDfaIziMQkXFqDaeF1kgbyiB5AP5h6kolJuk5/DyCVgeONPDOiQF+gCgcbjWw8CaEtXljqSDpg
mq4YZ/ccF5Lns3ZepF4ETBJfrCro9+vogvb78VTTwyvpJ7ExiXcB8NOzZ+/L5J34li94zjb7wml8
DMg/ujOAbnLJoQCMZPySC7wpV+/Cr1L3Vggp5iLAsViI++7E755UYVUeOuEvmQD7ecvP6ADWtaV3
NRZW/gvV7iNy6IIlGDP2sgmMhjphw33EJrXYk0bUnqQ3njMeLlDvxe3hDXoPUfS/kKRrnJv+ge5L
ksiKvTiUV+TTHI0ErtlSBnX+pDNa5TLrwhRIZ3TOBWDTpws90ONlSAhSrXVzmQ0St2Ym54pqjzlF
8yiVWngAca86ndckfhrw1cDJ7ZaKTE8CubBcGtSYSDn/UPS9PPjyD7aSREFOEiGuFmc13is9BOG6
4wnSdnuB5lRPha7XRla7KJjmNLv+E9RibNysAe2fHDDVh+KdYMH18ujdkAAh7xXQvKBjDqMqdkam
+/4342Bzlw6sZSEoTQZcuT9eykYnGqTnzvTFz8eThHIazwFjxmXN29oicLeWwpmknom/RMhjbZsL
sq0MJ91aj5q0e5smyiqm/eATqVco1pqoI3GtPFFJYmZpPayrYF8mgI4GJ81tMPi6whkdAWZapZ12
KryF/E9HPEgFZpHbo/G59XmcUvIgg4uFe5C50gszvHovI9CFpd2tMzOdBEMcYMoKDDqIao+S8PQ9
S4A0wBPuacaYHkJ3R9DiCOQrDUTyn4pdZ1enHJ3+IiLvXbECon9lfWHG2AcxLm+ymF/X7Jdv8eO2
FraKQpoWWIKO4bj/cKOw3iay4GscgMfJZ7RejWFHahp20I8Rwd0iyG2rFPN1m31UGwoqGqAQc7kR
IytxGBP+FfzGiFifq41p2ghe2o3DV+gNHyrPyjaqCVq8zn9lzV0jLOZGzMBJGOORs7KXtqdG4eki
YVXGKc3oXPBjy4wWE7kH0qY/E6U/Tv32Ur9DyK0/LmI2ssZpo6OImn3dkfPlSvNHPc3dSVBMovLF
qgT7iFTunwDS0NtRdh+WRMCBJCqNQHm60mQZrTNC75csQo0ocXW79giKkdowlTA15vLhMjG0XJuY
D4xnZu7el1GAXjH2+lR3zl98/JGH6f+YkGyK1RZapjMoPjq8bjGNMjKKtsX7hJ7yabVTIfZ9qnbQ
Sa6eU+B/FEmOg1+GIwTA2w/0FUBL39HVaiELKaZwgFIJwFiI0RKl5Z1M1mSXoxpnjG6+y9F9wAaJ
tCS9ZnBDGBb0eWAM1WDjHtOVa+RPFviuFvE4y7ng2cXAZoPi1i89fpxEc3p1UC2arb4ljDuHjabt
95jHk19zcKQXLXMZDdV3lHEQjFXYREdB/LMGMpzBnQpYGxAXz9v9QYv9+dfpY4DWgV8jRVNX2N7X
G0HJekJM7FxIHtqi5wX5DrqWWMrD20mmkO003Hj7N4gqRcJlMwDn1KbijSrQIeMVTqqSYEfr9fug
NhJcjSrT6UAVbsZloQrZQ9Z70jL/AgH+chhhu8Zja/4d43HmcbC48uBIEqc8gRtQcZoX4+j05uwh
f+bJO5H4/35eWdR+5gk4glVfpHb6pzUcO017lt6KxBYgMFxHDHx5dnaVcLGX4y2mf1LxOXrEa3zh
zSbHsgdVXWdYsZV4VP/Cau1q2lLPLPBKgCpspKYo/Pi4sI4Qjp6MOYgLobNi4c1BPuaagG507q5M
nUH+zSe0t9kz7vJeK+GrZj8hULalAHYrTkQvBt2t6MGkbi+NPHEMl0y4TUSxI1PZPu0yJgpx1QM0
QispwiG/NObunaT9t/mkrmH+1MP9tdTpijLZoQ3Vca0nmJNamAAcvWUAFGOApvsJ+dXbqAaeAaFL
cR20TE/b9KoLGKJawjtrTRFQoSO2p1NiC0pae4B6k/kygTX2waU0xaS2/4g4RNNwWyBLLKyzd1W5
Gv2NFQfTrvUAb0iVYzyPGCyfoaMhr0uJdwCgFGHkcJFjYHboKssX1ZNwc2DoOojoo7bqGrzqFcpc
GSDh0DZ0tZiuV2/q/MkZGo7l4Aw8FEB4LQQFsU7wAV8dfqd7DyEE/nOMwcNVhVFtROBGtbs9t0F7
IjaXKN+fM8ZEkp8ff4ZTIOfKYuX5GuMTz2QvZJ6cH98V3A98Zbvxf5+FW035M8JERTzwz+23lvUs
kqVqm2/maUskofEmn/7k1dI7cCuqBKVIUTGsFvpRYeHNIQCX+mjCkPlOnw/8qORQzAxE2QxvBZb7
t9LAyigXdkQCOENbjV+Iv5OZS8TDjx22P39ypNZSPZxONtCc9w8Sb45rbr/hI+T9mhDVOTyPoayX
zBGrqcM/BsPT39fMqYxxcGQwgvgBUFCOXO15ZHDQhNyHPTIpN+AT9vZNupjZm9fZQraXlZa3xq7r
6omwQlbRnqSLcch/Zy4XRQLUlvhrrTJgvDJxdT7KajXWaR0bJA7n7/jvpT1FE77S/c/0s9g5sYEg
VwMs9fWytqlC7vvcTd6FCobcH0sAOECZ3UcXfD7v6uKYjBKIk0iQtNVVKOkXeuBapUKxFVRNyGfa
jukiBmwFrbch3FALmt9ik+jdGLY9Ks5z4EQyMfX8MDAd0253vJnXnqYibp3GyVC+73jRxPhgFxSJ
gbWt/hzenJYTRxRHQhS67SvSEcYTde/NpvKEjC3GwxgzSwBNg24/zFYKCkouJeoByunLm2Qh/OoG
nUT/5kGbndi5Oj1ihJmEIWMnrfjr3Vn8j9Cta5ThKR5y1EzOMbR+vWjkhP7igx0kvLTsC2+ME1wp
9QxO9ajjyTgUzplm2YcyICEfvdnNcCEbkEeQDU2bLG7pBi9FfA1egoMTE9JlUb0EnZ7IFVk8QBkE
xN2TaCnRQzRQsfYE8bV4L9RajnPrMFsxxqdue2ZO1I2nI9DpvELxEqaWYQTmDNiW5NnX/0Rxd7rt
NoVDeBVu8A0mD1ZrBOLCD8aiVuESbcDCEdhRyWswR+4WhymG5E37TWu0Rs81vRlsvWZUGPa9rg/L
k3+KbaYJUOH7UcfaHXmyXUzbAA9pVQf1nUZGB5XT6vPrIn2EoYxZrFL6qRLcslPuCjOSlYI022SC
S4PEzLzjoppOTTBRZfioLJ2wALeyGVXPcUmju+MEwENcI0Zrx58m81zSUaEDuSNM8oPBSVgeWBI0
bq81Erx5LIhAhfHiT0Rn7KavpbY6TPAr8D2j4xG5oa95EUr9Qi9ka4t6NczqBny5+3AxpNXaDWTW
CMxZYg8TQ8a2TDBFb/9BvZVmzWSHRFLHI3VMaLGaerxyQggSi8xesNwVRWhCO6jlVwIpKqezVW4r
SJl0y9eX8Q6qoj7zj9hrg2/JJYpYBYyOQ9iV07K1zZXYFp1M6rwFO0KI7to1H6a20hb/EJpPywfP
w8DRE6c9bXLI9ePJqy29fhahmR6gOIUS+Z9fxrCfXH0lQ0pn3cIf6pNvPpH9wSvPM1xyGYRgD2VD
z2cnU7b7EAdNwyFFS0TqjaX/l+kGEF+knXNncjgUAQtFj0qXGOWiCzcoV6TjMwCu3+dWrEpxvSGg
D/M7OXqKgRFKEXwjGioMzF4Hgj7+o6fsWFBAyqy11M5G5THDclxqR9HGDaDJSJoiZK6kb/wg7bMg
Q8MH5wU56yv+M9nnwt9WJbIDQze7bxHdkSCha5HfEeHeNS5VTRi93EBoGYqZZFzeAqQ+xMpGSnXx
gery2oQ9VpdVXoHZNpmFDfhtAuzBbVjGhDpfYvDduXhgK4nNNF1Ks48z6OmpsHuoPfO17/mVsu+U
ifbZ5BrY/8ng0axmXoY5P6uhPmFscYH/aiKvsKV9nfg20B4sKz5f9byqE1PeEolRdYjphc5djint
Q6ZWC/m4nXXFGP8uH8gdDtnZj/ZqDsMCZtgw5vbwYPN4z7wlGAc7NZL5caQ4Tsv94H1FrTDCSByF
Yi5h/BdhijdeP4mAQBTCpmJWdsAruAs9AZ7GuCaL5KlJPYNdEWdRLI0T5WSAyAJIbdr6FE3y3KW0
WoHpuMcpw1fpyPuYS1BriXgGi2OaTIuzka4V4sajgPCXexnnNFV/Q1hqCvSDYRWBqRQy3iUJS76d
lNCwLsFt/Rh7LYcf0bt/oKZ4NpMfYpJSvx1CMco36UuejNMw8SnSlUMfDxBu9r1GQIfizEd/+DyV
vP9eDWI8gyaM8rgp6AMdJ74N6eJiUrwOVu5HZKS80pMLwDK2bUBIrTQOlzE7hh+8aHfAfgwckk9t
G3CXDOIhFvUj7BfLy9eoFOWg7UA6ZArKDTV7NB6TiUlk48zxjcC9Dn5fZNturrbK8dKadV8bp2lf
zdqkINNwW8m9EGSbP9qaLfiz8qfBHPbCp6nOYUn+LUGPV9wto06bf8f6Du3cpLrk08fRdt7Sa4At
iPvufxUDPL2/BGg9HJAbS4AucBsNcDeBZGVpN0x6iCcC0gkjOPT0IaAXzvCzrgDV/hcIqWYOBL2p
o/vG5Ksg7+Jjji97dt/J/dg6QkUNBcdaHMiegVVlJWSFLBAv1gPNB9XLTV1l86k3fXu+yPC4DWNp
DJeAfRVGR/9WbyALWSdcpuNuN/ukqjnieeJfKqTiE9pYJlir1lXEmyxBOxPt/zngotrdWseJ9DGB
NDLlYNVhHmKTQ6+pkXZZNlZSRHETPt/2E+wqvKa3cho+Efjo+i70Mfjosr5GQni6d9GVLqKes58d
meLueS+l9v4i8JPmUFi2+Tnkc4i8WvUJiXyIsLXPne40n7dx4dEesVPrMSDIyelrEhVi/B7zls61
EHVMXU+ngID6gUDdZjSJDiIC7GMDMQO4BfqGbQpDcky/AhCYPd+BkF3iGma3h4tv3bCh0j2QeCxa
8jc+RQcupxWpAreZLruT8U8a4T+WJqk8R5b4mXr+xIov6jxBehaiZiJLfICyDF7gKcbci+BUkQSl
kO85+9fnA4CTHTRdxAxKef9xoTFdNtpjc/uqDuLstHQNqtcpjuAZD333C/e8W7oMuCMySXTO1D2k
mkoBC4H/sjajbzep9POn3jwVHWTzPsxq3YPECbWCzGSgyqze9BzHts2HhI1GpEoQc6LMDNVSkj5B
gzZaBUH56fQDyjwX2MMw2jgYRjtmUCNW7ir/xXOB2aPL0Bunm35fbDYSm9fSZGtIQFyqbVvNNqsC
cP1bq65BjImcWhaZEoAVU/X277xglEEgaEPnUnrHtGpmJhe8Qt/wiyyhIDwFWbsJgYvN0t6zaoMW
Y1clfl0jKML3XSLHtP4bDi+i6eqLnjkZBlNINxfFoB/ZHXdUKfWz+CcKNaJuwr/ovcHXzm2FgdrC
hbpXF7MUZxHC/oXcfQ+3EPsuL/CuQD4sdQUFJT8cMPVAim+BelgCADtavC/OOFyH7KbES5l9PhU4
xqHcWG+tStU2uC0C6LDlmIo5NYcBJl5bXJ27MSXDQjZy2OsClR5+yF4tWtv7uccKQ5/03rdjVrP9
9FomTNbeRZtvBXztmy7Zhpe3B1c3rKFY1aD/9rpoXDzahIrmauEuRqU0ZyNZb9S73yfAci8+taAB
c4ZQ1PZrD6k+l3pYT5ib0AAfcdNss0o6IDTaTvSsybjE/T0UTUI6aVNX1+D9A1t2vDIBCbnl4790
18fUWRxfbrKJVmFMJU5f95zB4Gy6G1tV5cQMY07ZFLgHN6JFdl6tgtvziXWyYYhzJeUA8PfGJ3Y7
0eezIBnGEu4XhrucJX8m133hP5uufLq2Guy4YhATXR2NmuKd9wp/kzBTiRkkvpjG+I4HPY4e/5Ja
cCpVwmGNgVHavkSFWxSArNObtI8TP0MvuLnqGPCy9VOO0IYoE55up3s0eRMjCq9e5oZliCjcJNUb
n8XGrDv6sgidbJasho4vZe+u2DvS7YinCmb5cxtwoiBHvuksmtxmHGHphMqMYG8Lzfajb6vJ0rj8
k5K1g8AhsOctzUFOAWSt4QH2qb36vATOY27psyLxiroBMZDOZDGlTcWo18OgRHSg/t3+UeXwKPa5
X3OLx89LGKE1hJaggrqDwxrvIluJ9LE0ogWhe3lNOq4CAJr5Hl4f6n4s8mN58+3MIR19/II5vU5t
+OOseU/GW/romtc57/gUXCIh0DIFMsb5CEhDgY8EmrxCGG21pvgNyVyXlj6wyJf0pBBLNgXL35EZ
EY/nHgt/F1ZYZFwPtofRZvSRHPC8wGrgPWP3G1Epd/L0uGpB0wAbujQUyJEtGQcz2rR/k62L2tvR
H4KAEhWENrM3gErtsgf04b6L2XzX89xUsYuhhgUfRwr/+arHqxbEO8cZLLzQMf65/jpnfTYGpgnF
RCzJ0MlNpqq+AOLUlIRC2LXw5baMKuk7pWiu1xbOEihYSd9H/u42TP20RDUNn9emUGWlyMH0CPKJ
Q9jfhMZLLF0KBlZ8QFVwa18jt5FpDB6ZtJqrYfeTRAJksa/KNyC95Vw6NhsAp2/ksa0ln3Ff4YCb
0xi5lr2RAC/402zfirTWTdpElH9m8w/R1kONC4f5aKeifhoJRbyxh/VFS5gH+JqkWaOV/2rRm3Xq
bn6UT1OL5Vw+5M2b84Np3PRlDhEFQ+143YmqeeNuD9hsTjAhpdPKQkxHLxJbz4JStKnpfoz01wrV
ufx1iQrQB9TCns8V7O3PheqbkWNMKz6ufbtw8fkPgzaRAg8lgmgVH7hyMrTDQUmCQCzEdVoudMqn
aqYaajCL23Brf3Pm8g+GakHQVhQq1BxUTuFfV4D8PveCYweVyO/bdbZpnSwLQO0Jp6NCf8/Z5vsh
kw+SQ2QrtTzbC4B1AnGSnhrFycp1UtpEoltPphyTgBy/84VU6+rU+Fsr+H7vjkVO71KUaYZrglxL
JlndsTadC3RcDmVy3EU3nGY5e1r/+GItCMipBEyk5H5s1cAt/MKaFRYj2qoQvDsbeQEsONMvPDoO
9Vu1kkYiLmhDHlyNHc5o4mgU8UyeZSEUHvuUQ7L+rlgaXs/Ic9/Bv4WPDedqMhfKgQvPAQGyWXV5
Nq3V5FvvC862FnToT9Pgfd6KBemihVQvFfVW5Fs5q8nWQRG/fwRyxeg7bTTUDV84QC3zqgWD+nKM
sFAYMtiV1xdfnnbDdlCYpVgpayyQnrX/VX67VbH2cn4Rfw/1DkOjbDqkG5qB6Hrjm75Qgx8StdTN
++zl41ziHm5nKRLfo1yKOxLicYEDi3dv8GgkDhPXTjlgclLyJNdiffNqXtFvP/0wlPe92RLJHi29
i2GUpIvRsUTiV5XzkUJGMsauTBgJ/oWeHqSiH0ZAAsGjY34g1sZfRYu+RUZjzx2WFDlW51kcDRya
6+MKl11IWQREgO6/g0QbLnEopEzsKyettEY7ZBa/LD7SMP1hcKUM5acpAQkgSGPjk039sdmK5xWq
u/GN/FQWAz2ZVmogFv8TuK5Ux5mk5LxJQPXCZ/YYpoF6lmwOggyA65V7RseXZH+SCNfYdVq1wjtR
uayfOCQUgJV8Q1pGwhU7f8TmRZ4QZSCJvyoPEExjIBFWv4uuQVi+xycPkgOFx8Irxvh+chz0ssDY
8VfA4Iqv4C+G0Z8lG4mmNxfiD/cOUpyMKDbm8HBqXb6dRIaIbWsHJG17re9y6RNmjKCagVhl76+S
ANyyNLVbu9Qw3ywwoWpjvBSupMeaRdq/27mwBhMdySl55AzYgojUUmsTMSszw63q46pGUJ3vzQhs
xIiWTKwGDDuGxYaoaHijtz/ZdYmrbAipQgqS67I1o5RFczj2nQ17T7z5M9cfWZUuEE4EJAd2Diuq
mI+4oIt/AxQKPGrLTWdGRQU/MdctdruODl7WLkyKq+eFU01C7kWOgi/9tqfDoak/XCCFDkTXxUJ8
HIUGK0BwEizzt65wDmpEWFx5YSEXuwwpHvnUXbirmdaNtkS3cwZYwKcmJj7/vT+0quT/VZTky7Js
D/VTR8e7lC3FSBBfM6nEX/tFLbb5H3zE89654cPgoG1jPnSFC/J3SyS4i+8QM/dXuYkTwDm2eC4c
5HNKSYsThqwIMyZfvgVbWI1gWCWuTn939sjCQLObIZ13p3KuXrqk8pvvLKQekJjKsi1wyMbj1CVr
9ighpqB8Ek4LrGHA69SR9+tvNWl9Ym9luJomBBJm4WA3LoS2z872sva9PBkXFE5C8Eqi0Ncdx2j5
SXoXaINVV0FmTR9YlXCooH4CXO5BDD8Yytn3+FEJLfNCEQfupi6Vz99SJ5dqcWiAvo3NNXw6s9BE
Lovb2N8+GYnMQ8OKMHcjeLw8BEE7qCEo/Ffl5qQ3S8uyN5fwkB2gPFn2kMH+eFmwyHszl0shzpNO
02RC0cj5jLsCirldyH4UDTYE1jMUcyaDihOkSPNsnNdzy6zZJ3zD3BkkJ0vdXsH1577wE+wr8SKN
l0fQ3ZJ2x2ZwQIMO1tEukyo8q+rQf94lC2bBX1pafjPeXFrhVBAHgQ41PwSH31QIDEJsx3/ohxUb
GT9EY/7wBqouPTrUydjsGpsYHFmrtZcmLtmwO6GkgjtVZvmyBjKiDQ9Gjcf+t9/IdtSc7QcDPpUv
l0CfqfktrUW2D22cpEE9PHVffp7fx8pLL6ltUThxe5UdKGdPuGYwpVuO/Yrp9WVMXUn/lLaILE0C
Pyu9zg3YU7YO8FXwrAxYSxLbUv4L7rEP0qGpPjwTmHYHChlohdICy8NA8LjxjZVu2pnOItB2XJgo
DOGzF2u27I9Wv5R7HOTsrTF0oZTqQ+nzmGfq1wxmS+WT9Yo9vjDh+X19ZTUKxPPrDdpZADOW/86S
CRENRVqCPG0vTS8+62vrXyRpRXdmjDRtWOY4TDG2ZXLZWIGV1mN0rS90rmMmpJkdp1wBVmjY8C/k
IICq6MKM06vcTwhWDxS4O3hJKhcqshUo6scj3v7eCKNZSEMstYy8yyO5Bcbvxnl9Euw+xI0J6Jk0
phRuaZsRRWmlSoN1QnQnVlci4k8HK+FFhuFeqqNFi9zS6zhZCUZDS2xwKb+Ux+K6X171eooaWXSx
vF5mECIbNOssuQdKMH+iObbnRMn3gmADx8oMYjpAyWooEhrj9lRMiTT5ZJrGGfko3wYXdNNV2nXU
fBThWNwiaDh42Kp3mDQD84gMCsNWooWLGWCf6cE9sPXcZCWpJW4WozOc7nQCFnplF/GnhuaGhlUD
tBmeKATAAs0wuSxWlU2jVOX+E1CoivEbDX6J6HSTGhjEF7Lhup32EF5QGFVYFBunxhKdwCjjC0d4
tyvFJRW0vqmG49ShvPQy2ls8t697BVA5rrei26g+gHMmGdcaJZoafYuR7ZY5EQbOVPYtuOuJ8V9h
3zw7neOU2zFUaWOVADcMyUqStBi3GDNQaEkQdGS2A001cb+XIFPbuYOdZ8BwmBP5wgctGlKk/gdz
7DMLoRkhZVXCmiqyUwHnaULcbNrnLe8c640srhah4L/TaqrIROLOdSntBK0ImwKsQbPKUBQv55W4
PoSWIYwes5XzrkRi1wQ1oY8bkKHs4IfNmOb0S2v1Y3kcmapxwKNSAWRd1RnEpfGjLR91o/drsRWa
34g0WResBLJfBfQdtVff9jzr3c7kuP6e73D1BkTn4dds3JH7SKh8bBFP015MN3k3hQDwVnN7Dxwa
OVvsXGHdCFT9I30N/Wzf40UAQf12iQj1Scno1rPHsINwZo1PqE/WgHEd9o0pEnNBCazQnrzLcYoA
TzUCXxEsp03Y/EM478grshGT7AYa+SW+auhCz9HmwHOE2116fO8rVUOQWXKfH2g+gsITZZRucI6G
45+IFBXzH4MglwK5k8RyEvGcocd6NaSAdp5kzXoQp/sCSogry8gFko1ZL4Rxzse0Zv86GWC2g4lE
w9Y6NDvpWuvE0XpzxErZD1Tq1TZR/DAyLa+i1D+8lv5yRBFlNQTl7uj13PgHih91nXFEycaim01M
Uqszzylc9M49l5FTwzIEsZVUySJ33+acfBFVzhcZp2WE9ObQwQdFFMJa3UJf9XdOjJG4CLnyFKHj
xv0Hnq8LUYPcOOwm0fOY5XOsyNdYKsIQirLIZj2E3NJZd9QO8khOPAZjeLBeCEW/XF8jgBrY+5AC
1xsNCWWSkI/bwaQzNDEl0hsc8tbO1rgF5jYuxzMIZZKMP+GHrc1XYPi/D/fJHfqYA+k29oBIvyHZ
Mf+fUreJSrPvkZ4qtMXtKP7O8G3ytntClFB9mjANRxiDrPg4EPn3/O9iVOm8/wiEfFqH0i/pv5Xa
eJ8N0suIVRHXykenve2Wjt12hTIQK1b36R3i8S6gY35jjq6x4cvWK48/fI2TYSlS+rH2u5Q5KXTi
OUC6TROpQu4XnUwFD4oNpYnR9c/wJp/L2a2mwUs1C4C2R4NXLVQ8/Jl/dwRaa8F+BSaTnX6vxVmH
EUMWWv8gUGrWf3+Z7D7QiI5tX+14rwOHO29rOMUmyfDNLXUMO7fcX2IY8aKctaNSK1+6GUIiH9VO
ROt1g/QAbIobUxA5FsHD5ysZbJ9vYcAGeIsWOOahm78xU6RRcv/toQ6rs07XIKXXi2pSHH7cLoOX
w/IjqY7jhWm7iLkIebW3w6kiyndtTovsNMF00nEYh6MvTm1Vce9G1cXf7zRaY/rZSrFTyBCK5+L6
E/vGOKFAarefDFepM+jChsWaR6cAyI7/5D7DGam4XaVzUzm+ZwacniTEetDi4Jk2gd2/aJg+4ugH
ndhMqQzkZbnqANpm2C0I3i2L/UpvCLEgCc05JabtKZzPQ7HzPZSvUfZ+DZGTXEcB5+Lc5B6UBuRN
Bk9rugOa+N+ne26e/TjLlwiORXeMlxPgdggmI5TTU8NG0X10XsbXqQijuhuZBrizEAcCw5JKDj+L
txx/ZrBnqZofAyWS1qSqV9KkqJf1IZdbcPC1gMLobMS1XvDkuv5srUDizbc9+IiH8Vj/FxYsbFfd
F8BSkWJ1pXaPq+fdNMWh582+8vGr0VFn8u9nFtSONz0douPB+Ot140cI+c9lCjM76fRgWCIk9ic2
67IZjdxXPcyfih+KyVXDL2qNn9Tdv0XaCG4ax0SPJn+NdX/AqZKGfoJcoXCpN5XUccF/ArRlQ0Mw
CUHMlADlPvfT4zhM6eqBPFFTi+lzZikGT6bEUpSW/S854XjKGUsDMfui5aNKdECfr1zzhiBMIHb1
rqBkD6OuhcbB1lxqIrYnt9FpT1PxqtheGD55sq3RB0rs6ivJA5mWkGgqOKzQucBnhNCBDcfLRPoN
4CYEroRiQ/Qd5uGSYjIcBLlxLclbhOdV5pnsw+znfrsY8hPzy11vBd8y5n2vUAZfTYicBdTnkQBi
qzrg6GidAl99V9feH4y8+FxD9pgyvMEKbkHbuLn9TDMKlNiKMPfgkv0lX6sGdx69Nmkdzve7OOQ0
5v/fmufcqORDGF9H++SxiiJ+Ro/wgAFwg4DpTm7+We8nxM5qcxjs6WUoH/BvSutzC18/G33KPOUG
Ra4tRaueGw8oyPqSyUfh9RtkgkR//EulhOVBuVO3oDoBijsVZnv0cDLbfLxGWQcpSyCafpE/K5XF
dpQbwXh8V4TvUX6tir3K1v1FUGBWOXYhsWAU1nmPCWwlhlBE7krP9wGApUKpSxmNGoMcHLXBc2ey
/Na6AwXue5E0CSEC3Lx0nScEQInYV5aQ7gYsVoqCXFNr6gEntfenaWOkVDJ6iWinS0kVP8vOKV8m
sCp8UySiO+/nIyRt3gWXVsB2znyOYZ42Zft5jBKZQUyKI79kNPvtrsBXHIG67FSEfsqUKl1SQih1
QN57CVk8BiosdMkixyHsgIlSj8tOmTi972tcXoGQ3TyRBIHKN+WuhU2aGhzX70wbWJIGOMb/i7Uo
yHJc/38h4zuSS21paJHTUdsCvpc+u2yZL6ibF2SaduU2XbkPICwTOMeFjAwJxRquhYr+eEf5D/Zq
bP6KWoXRBG57ayu3MnL1ezjHiVpOcVaV9FNMjcCBN4BkQWn+CvqW3+DJ1SFKOzmGe2Y2/nTP790U
6CNhDp3FDQXw1hA5c6CD3n9ImhedcdivNpC68EQORZg/F2aQ0S96EkFKybv+XfWNWv2xloVBkvVB
lbbqmRuwavc4UNuWtWkmdTKOvhCpu04aFuo9ZiZ4a/v8KmuJWNVhc5nwX1Jn88UJFMwmj5n0WyJE
OVX8Xs1vCyCERvaF5RHSANs8ANELAkoSaU3TamN0YPN8i0PkmWJXoLpVfaCI4v3UP9KbQVs6v0JU
JPAzuUimSCUZIaTfuGczSAOaYIg+OuJKDDZYxmUQgQqesNxwcPgzYV9GVeZ7isPa45bvfxVe2EyW
A+Efpb3vFiHlCN4Erngc+SR9OdPhIDhH1/nzta4ExyW29JBH8Fy0P9ytDzyquQpPX3yCFnjnvCRp
XxNFP0ckwfaxkiEjUjiCm6yCRHYX9wuo5f0099NTAMM5z6Iy+Xi4SxXb31DKmQw4E1LDSWr605Hm
UpVldQgGVCLKrUgx+u+CYQ4hRH8F0Af23NYjmV18CDu4eMwly8j4EV2tT1og17nwt7bOC6dawngM
7TDh+QJGBxhtcCOnox8dH5K8IspSZIsJ2nqdJpDoP5DCvokuQsSHDzuwkK4XQESnsTruFuFLXbUY
yM60/IkjD5k+ycg6HvZgEGBBWiQ84Bq9xvwFuQ7dR9+5p+ti6lWd5kHhZUq/Ic24Ocxb8bosFaXP
B+1ZJN4VcugbRIxV0GWQGfrKvMGaBZrRFvywWr2qfiB9m07+Wuu5Venj5votXAqFl/GlelkIF0q0
EJSsKW25Qd3zpYQybS4UEXxW/pys6y8SMntQ86zJVVuhYFDdYOEu1upGbAhkREFdE8wDz+8Vq+pn
GmwXcLAtdvG/l0Ve8Zml2VdjVQAfZuXPQVUmNDsdht+Ne5gY1ZIUGsbipYapskh5yV0TetMh8ApW
7bNySYyct7nK+72DQzV8ZsYMoXyEpVQP4/qqQP1aLKanNE1oKrZDjrqxj9TswXOO4eYIus8i+2g2
PNO3rRZ9N/1iuZgUdHPMno/TXDJ7AaGZNXzg4IAdi8iCfsEdbUGrlZZhXrg86OWwqcC0AGhugfrl
Qbx6FbBoP8vAM9KxO2Mf0UKzxPAjBko7i0hPmh4jQ35/KJr5lLs1AbDq4pfrDAIAcZVgLx/2GP9E
Tf29xEUILTYNfHhadCZjeTqy07NUU0gJUyjWs09JMaY8074aQJdvA3U3fU2iVJU5fgI1w4kzpfe5
Nwjk+qAWfTIfMdTNLub0ozmbQ183l/soNhbB1maE1gfjHw7lsaDJwy5HYnMOml/qMxcxxckqGnnt
JL/7y0MTR0pfUVV0QvR6XJOzQk8Q3DOpliKwjEFIFXynhy0tSIqQoBA+Pm2Vj/EORf0CF+5KHqX8
ytpcHLGk5aoAelhh084tKdYipbkWYvcNmJmsHbiqUDGE7z4A5EJxYTv9kjE5s+jlRkTYndW0g3Vq
zZcigE2JAMoUfO9UTCLpxdUcRv4fsnmCamDF0x4ShtFeR4Ph+KYQSeayrrCY/3M3Yf2i1K77mzkI
6qhPR4Ownogq+SaSsZMRHNbJS4Q8lyJ+9nNynDATmZlF5t9sC71QaMGjTN0gBqF8imv2c12Hzc3G
XcpGtrK3vZyUUnLkpFvEMJPl4yfR50XdP9C9DnRTH7y6OLEyDR8hWtuhJJI15p8PCPxiEJubmoXd
CwQzyXpkrGSFSsgk5J3D2oakNRmsXgLYi5RaeNjJHZSB88VtvTq+MYYDGc8H0BFoMHPGuNv3lyXf
9VtcRmXJQbx0bex8G0CReISq/lr9weFZ3ha4UmqWm9ctGPU/PVgIfwcdoKPUq1QXR4GIkFSOWKLC
WbeC5N07vYuJI27jfYbNNATof7yiQJFJ0kgNehLZK5rIcCq1n6fdDhXNc8T1Yj8Cip4HeGbjt7dj
zH7lUbJwCGLe9d0PvWv5my+yfyeXF6/UUZJ7oSRhEoihaNoKJ+bxdzxSGiovqAkbmlSOidLnwoE0
meSzJ5Nc8rnDL6AfZkcCNlFXSJiOlRgdyPWpCjmXW1cBS8Plgh5QM+kNE03EZ3omKrrYnoDaubki
JeH81Ce9sVVWGjIBmCmwM+Cp1EBCZteF9EiQsHkv0kEsFEn5cLIUb5Hk7HHTBxLarhebP1ADyw6/
c9Qiy2PGzJCZi5GGoR+rwBN4QJEN9JDoSq/w8LMwrSwV8SL78ygMuNjhXpyQQzJEoDCPOB/NQdNv
+ULsGTBNH13K7Ti5EkTX/0+/XthiabXQcrw3LXP5CAzhQWmjJWNZYW0wRcNUoqdYe2sr0Gi/n2Z2
0bnAYNGn2fZ0w8Sk82sflhMrFiffiWCzs8ADhliHTrhvkoemGdJeCOKe4BgNrKrbktSxhuNSuVZT
qj5dRppuYRwLH+kKaobkS0aqEMEqIlQkn3AQBCkABJTrbBBmrVnEBmgSa3sFxgRkzvFP3fnEZ9SE
oj4Ma7rRQwwMWUNvgBrveFJGq0T77CZLeT7Ky2bJ3ZKACoeQNk7OzW8mE+egHwOitHBtEG9eME0j
8XuRp9wiLczbUwqO6AjlHxwgeepnk+DFQlGUNq0zV0914bSZC0R1UuCOaUdos9uDxCuzBgVeNX6Z
Z2T8VBAWS3E3Q4WxnMH8imYg1HVpk81GbAtkMxQrT6D09XRnCCADPQ9RiSQXlrGvJn00D5D5E60i
Wv/SrzWr75IaXraRVNmtWqncTPXeVJwgdBHvpNwI6d/CEtI1hdxbGXLB/47l0hF4YY9ug1Wdu/5y
53MnyH3QlcZ9vd2ljh7xnw+DX/ptQm2lGAVsedeW5vvjosJy7keuvl9lWJz4eUz038i+L7fhj2O0
HI47O/NDOPdI9EH+QCrhJ8vJUdXDQo1nUJ18fKP8+mekhtZ3HxG7IKMEWdyfZhn+zEoDZIRmWqTZ
umEF6HqdG49OA9dkn/xEo41tBJCpvTa1PRjXSkrA4O3qUm0EujVPHFC1jM8rnLlAYlNSmEfCTWNx
ajZ+EkAxz2Z4e98ujwQz8N1ylnzPT3xEDTacDbE2p/zCseEHY5E2DLwRzc6vBNPl3aaY/fshadON
asQcLf8mZO+FlivkR+VtS4U4cRgy/LQOFGmOVMjHC4evOKyWf5zXDzaafGIa3/1xXOMSORaWUq/U
BExZUlQ8sQVOh0Mcq9Rvzl71Il2eflgANlcn1FXwkoKtUocVd56HeQJDsLk7kjTR9xQRlKaWckMR
x5kFHjYmrp8NnMY+8F8/N0Tj62wMxVO2KYKk8pgGwbK1ps8ozWSUQs+eUD6nt1gOF8PSXtjFksqo
W+u+2vMmUbDpNP7zkt++eHMLooG2rbsBKZ7RrOvIYw7QNqehetA1B/LHErfDufWInJrdoXQOJLzK
L9HswEGPLxaxDv2Ilza4jpuACE64TUBiiQ/JmYmIKBzJ3UXzOGgjhUHtYyHhjfZ2YFr3MfiV3vmj
xUZUPhwY6D1uRjJlviTZDv1tKfm0ojN5j/7mS7Tq/jOaURvzaAh/+S+PtK29DtZEZ8WGSweHoxu0
1tVxtKvD0M/XD60mZWIQGyKWcpq6SmKDyE50kRVBma92bYkz3q4bfVKOUH8BWIdL4ZmGgPky9tmp
kp39TOszHyqEPvnPIo/B+5GUQN0MJoWmzFWutNs2dWTCGEkUgz/39J1Q5ZMJsPiq5kzpkrq8Q4oN
EzEi82zb5E5tQGwYGG6kQWWalo9jHgIFEmVRG0El/VTxh9d/Oht36pZ8z7HfhwSPr14bJGDkVc3j
oA2++1/aiD9hdvQZMyoyTRG3lIeLTEnoC0AHJCIem94TCI6AcvAJ9lMT2nExf/CLy7LiwWl23m6M
VRI4ksrcqd/qsk6K9tlMBktJQRwC8FMEKJE2aZ0c+8rIcor99Bps6f/pjYKHe/Fb2248F78GYYF9
TrD2nvOyW5f66PN5+Dvuyd5p/jfmOSOZ4oWPEhFKJ7TN1leSY9pjhPSiPrGN4Aq9P0rzJxI61WtO
FBVqLcfuJdQDVhEos+UlL1xIDyR+QWvejlXlKGZxGWtSmmvgkoJFh3ujKeZyzocZw7LevTQptG4H
hiMHANcXVxffgIUJdlGtmmWX0Uu5y/123LbdFhstrmzy0I26paJyZWUYikNYKGPs8WnwQoBXUeO/
GXSbcuLFpzK3odzKwfK+R7zhU1JM1Uc0c3uQTDUGQzljc0T+eu7CMXxQzeXd00MB84W67Hg/+7b2
R9AioJlWAnK+wK8GjfDb5acqOy53qzkUuRxi4QSnHBfqnrup1oav6LhWJjA5/qEDQQz2tE4nR1IL
u5FGQrBXSCjAol5ua7ww/v8fRZV5FXM7k4aqkDc2VoM0WPF19sG/7i4nsIVkQyZx/Qt69CbuKeiR
IyAJQoLRg8iGEJVM5zDlTsmhT1D4wN6A4jpKJRdBLsbMV8+tLjiahneMGXUGp2i6pwkz3Ud6MJp9
YxOAxGuMR4alMbyVbEwGSY5dHlQvs4P9x3Yoj2tHUbxl2ge9+aG3xEMIHxc1BuTc4KR0/xx/eavb
/aCMfdiInFMrraU1Lz60kMkMgByZ8EBNqxK1T3o6mZZghAZdiIHTqJL+i3XxnohtwBT5ASXXe0uC
oTDQrkSlRqHpgz5+iQjewYyQ/j6v6nSdHdyD7SzcmsgcBN3kH9BTkFNahu6sCxUfyrBIugOcEkSj
83ONc3fqme/B95qFfqR6tUPeq5qbFdKqrRLBt4lZy3bch3HmxA2kUHEiiKAD5VXPXvCYO9zMYY0m
GGLO+DOS/AbB6aSBkuwImrV9z8qbpYWs4ldF7xfuCY6xfySSsOM/g8vhmBcc/WzEOpqTg05h9pll
wBkO4jlj2+6ELU7L2O5FWxyTQgzUocO4+k9hxuFwek3sKq866Y4gnHks7vyKxom3+Bt22iYYimpH
4zikATeoW245LB5RAL1hKJoQY0kVj1FjLKuZwMHsiu0OQhOrzdE1RyOq/3vIKiOOOJi2NZAf+jpe
MIOMDuvvRP+v/o0NyBxa5gck+9IMH0BEN6KpPKIk00sV+gnGP4TNgs87D1ZTdJKN6X+0ymMpb9jq
6ns8SH8aqxAXJ9cFLGLzHcfQsdQCG39XYkLR0pca30u6dNZKCcdOAu1GfTdVCXP+MHR5zxPEPd2I
YIBxkgxoSdz8Hg1yHyJLmNem3iJETBUQERQjvXCNv9dUvkk/KXjPdqzhhZjP7bHMkOH7IMiNuvwi
hUSRzEcPfz8Oxwz7VnK63XlEa+TZSyXvki+0EhELmrO/O05aFr6nuEdO96qO1juqdxnwhu8OyFBC
heNbY3kKT628PeupOSDVm7RZxs6bkIUBOnxZjRqRARlUrebakQmA7GSug6mbl++pieJ3gP4/W4tZ
jY37YU9+A9cGtOjA7dyEI/v/LJyV75oZJyydbJr3rEf+UNXyqbBTVqSSmzurs5DfM35bdF1CkWkR
ua6ne4S06UXFTF/41OoJosNy0phuXCV93v5dW8wVGh6rryPBuz7oPjkqZAyiPV3tcmjAQ5jMkjfx
iqRngj7mD8IrbtsGkbxKE/dujeG9A3p9y4LHpzWlA/xdAaWZcJAi7VYXECY9vqWhoyRpfZ8b28Ig
CAE/OT2SgaAhVQSyYh21yOH1Dd5TeH2pfvar8mWzFR7mzKoYMDtp4tV8VKFRnFWrQYnkJW6XW1Vh
knSNbRpV/mqTegb4PtjQUt0S8vOpCQz2MfPO20phRSKP7NI7Kb5GUg8aZ64+CvPbHva3aRKHLAu5
cPJFSExm7VemaTNDwNRhB8d4DUMQaakzHEerBO2Gh+ZF2/dFrGZsH9fZcPbFOapDK3xXTFqDbcpI
sugbQPKIb81L0MiETTqGg+vQ/hcGksOYNIzEjDJ6OUFjTDILC/jEkhoGZPN69ujdzQcPfWg/k+qB
5yXMrzcUuHk5HwPb+Xx7h7kRqz+zlC6ty4l2br5QHtif3eZSSmwVmQI0FAhtIV30DvLZd5hnVxAG
bNdcLvnzVYkUUpnYG+vm37ooFkVwrKT/O0Hqtp6FDhoaQ/iV3jb++Soqd/HNFmQeV92XySzXibaq
7MTSzeIY3Uu0ibgVfn0Mo61pU2113sk4bEfUNwEftd2+x/cdjIMDZCJnAVEUcppglDvPqnXDRom2
TfYr/39uCxzDufkB18+tXZVAhz3RRw5gTvMYBHG+9lXoYStcQwmi+icQcRL8KmmEpyMzx6Xp3ujP
rgQ2HQp0ZQ/4CfSfupkFqjN8X1eqHLy22NDTLJfwA+U+KyVyPtE/Q77jV2hUtX2dVR3XldTcaD3L
UPLk6mbZvrS8EymPQi8nAlPbvO/XePrIKpRh/ikubtM4tIlJYicrg3Iuu3h4AoEp6Noa+8Ybw8xO
4iGz3EFZklw6q3a441HMJ45JJ9qBhQp3dw0Wr574CRt5sVAimR2H2EblrTqs6EHqOO/ojdMx0sgi
VadttdI16e2bO9lA/M//0FTSffkSIMTWMvuxOymdEdibqN2b52OyToElVtmXosB17rUqnuNLfiO0
Rsw2WS6/ZJ4qH8d8WfXdvAT/saDlcnsiEFrSkRAG23KrJVkF8KhJzRA3fTbIgJnBLVmbbPlwtVdi
q1j72H2sXRLmH1aX3Zdy83kALzPtQUKBQuAp7DP38as94T2d2lXbW8BhX3IgUZqPk7uNbDHGVqY+
Uvih3vuDekwPvNo9kAiG6lnitmrMUK+0fkwtnuI4w3r3nE+VSqk03zL+m7eMudN0fJJGZu17f76S
7iyugEYVsJeEkXrGkcyBCD/xw3h2CY4IUChlDfsOAx8Ck+aaunmEh3B1p6L6Oi1XbnK55Glumxb4
8fVrPBKt61f4h2Fw1TxV8GX+CASdOY7y5VBHhveb85umNvTKTiwL0u0TFyvsWPb5c5KFw2F7nC/a
aGHXIWCWCRiqbNoREIy1FKrCX79GRLjaR/Phw1FWU89gwumYbyDguBUOVxHdEXXqBYkvFclwMOcJ
Pxy2Y0l4BkolFXYw+5sO5GsBQ4tGltruPRYAJwGvX9w2bIOsK15hOywq+Ob9VTXnNTaLJWBG1Umv
wOjvRFApg9DAJBI0frkl7vY+klKbinutKj7/zwJjylQMmFe+WGHs7EqzkPql3MkOXq5CHPOzTito
VW8HZPUvj/bsAD34FvCBdB3wtUlzel/6eSSulfuwId1IDznohsqJcn+Y27dZufFoySRDOU9+r0nc
JvCVENOLlKIX/yX6NMpGghM9FxdpHBVH8XBmkiEwsVeXfnEwZ2gtu3T2Q2luGtHrm7K3pMf4Ye/i
DmyhfTEVTqIHikMoYgDOrm/zTnOxGhNl5YMF89/Z9VzFPPhH1Cp6m+6uf3XQ3kFQBY4ce5kqfx19
bOOTLyZAfDzmp5WayTfysGVVC6TP8Rxr7iU2fXi+TT4rB1Na2D80255RhpfkHY9JnhN+p2Czx0Ww
yJjHAv0gYi9I2bHPAI8B42FG7XgXWVcg8u2SjNAI2DBncK0hc2lsonpTLEwStK/+4qJFIKehZJ9T
FPY7vxMLCG5ql02IpEoKcL/itSwYB5Vpq5u2q+fQUyMFN3NXWKCm4jTulTLQBIa230/dT7uQx1Te
C6XqrJe6tgTSvv0LCH3KcBJ5cjBtLQh+h6ROJNwejNXE5UXwAybpGSB29+AVRu0XOOHjacb4qFSh
k1oR9oqJ0sdwocPo0kTCpmZRPDTNi9CM5EZV838SctRHQDiLbS0voAy1t+1iU+echdfp33Ye8njE
H8gKuGjUCLZy1bWlZ8aBFYFY7+t+rKOUU9XELkFm1uTbX5Ch8YgViSwHi5IrD3m/2zNl3iIV0A53
xjj1Kyigq2BnC9DC4hpQMObGk/VDZHMr0jfTqjGf7ItQ/fVgB8gGy9DanQi8Vv5iXOhGk9X7aZyy
RwvS6SS6kJ5KKrdGDffgs8SJ8MxAlfNesO0zLzIUOYQpOGEOte66npqvT6XI52FHd0pgHshc6B3c
W2F7e/mjmhI/nihC7n17l8TGFemgWfHQVeH17yKpVkiK4Yy83t8kY7tUxO/13+Z2AjfK9UBIARzc
bzOHeCYRvzicBVI3IpkZieqGCvauRRZdQu5LfnlzJCdc8i0+KGW0sfOeZGZZCmeThC6YMPoLTsST
kMisEtFvOFKFRxTfuOPxrAFP37i/6OZ5Ac1cBkST4YeH3BlhZfVKG3biAvNEeiw0DT0FH+RZjd61
eAGQ8JOt70YXP1a7dzTgesLQPYAsg4BXOl8o7xOVBB9XHC06wIp4E9p2WJpz5oJntUmrFc+YgEVw
YFWVCUTffJQjSRSZrMlk5LumXrAHtAHqSxLOj1uz9yLWoYNPGaPwLR1TOBacSJZd4CUYSdAknvgw
C8g41/m8ItJYD4f+LY/AGyxhRfJlnD0BRttbE31KH/f8ihedDG3/cv3xoRJ2fhjGbeF7SLzBUiEn
8vjqrxrsgbRoINSs8PHrnN4z637V5eBQgCspeMdMkhGFEYctPbOZj51EkB+hjicp/Woht5lkwdwU
QHt+ukpTnqso6l4BNtN4XPh5bg6ucr9/NUAzCwOaMGN5TOj1HlGGW81bF0lJ5IE8LUsN+X8G8Xsy
SYAe8LtNrVCxKwQA5Aoa/2fh5wNdkvPOQiEzzNA0oL6o2zxrBtd6pjASQAWwmMZHw6V7aAkE3+Kd
kEeLY60TqkoZdyqhFbq30zTlEMYWwone/SqWRYgDC70uHYH+kKVKBJKwZisrcN3HPgQ7vRGXw5NQ
ATH2Bmywu8Qa8l3urNNmnOOb2W/oiBZ1d+IlGYa1epCqJJicYCaEmorSZS4/5ftp9O1RPK/rNo8C
I44DRmQuSTErxFlxk9W6Cz2IBQxCBE2NidOqNuk0rJ8mF1axFY46crQJOnW42TbwrojJ6jkYftLL
6GPFxoVYMQl4fNfSBhJ8rnKyGjBEjbH+Dh1/LqVBTzY4EVd4KHiWyetCA9sgbBseh35bc34vsEzo
vgd7db8/6BQ0R/Ap4xcVWEzOxo6vrvA/2Ea6iaItmVwWawyxi3gBUT6XZ1LT4HXXDQOA0iVpgXya
Kem9TXBUvppPo7dC4XQ6cqA9pF4cwjMxZ862x15sPoeqVMQgYw35rOLUYQbtb+qcH/l84HvigzfV
KJ+06mnqfzW5gjSdi5wYCdZGVGZCNveePpM93bdQ9txtrX7uCOA3iIbrLmPIgxtN+347tH7aDz3w
GMYCyd2qkAMbShca6xxU512ThNOZ9cXAHwLYBhsTYR6FznemHBX2PZRWC/f2RfJRxODMY1fl0tFD
4RbO+2y3fjbbX1p+gJqxIYs51n2xemZWjfFY5AEufOjXuMVxh+qfzoed54LNfiOK8izfHxbVNIRM
dsBhrVKUKPoANg4VI8wq/erABmATQMo3Jdqq4vEprTf67RTl0pmtjNob6tY3j+A3ILdlF/t7BnNt
0TJ/XyH5YDwxYtV5wVpeYcHw6fWBRgngcTBYwf/UMX5W8y2oPGAhO5TcvkOiD372GRHIyu77b0Kz
kYshdS0jiKXAsOLy8y6QoFEB7WRcH+tIxd2ubb0zkEqXUN92kF5NnxcYSg2qWMvJzg/0KaNNPBxQ
BRxVHOOACcb8TcpJSHJiX0V9TkVQsKQRMzbArfcA/e96LoB2vtacUkRIgDr7sp3zWqPIWvEW60wA
k7JI1IqxoToFLGRqL1tz1NDWMK7Jx4FY0ovoe5N0w3BTu4J5QBsI4YnpiJG77KrBHFbRNtxYnJg+
rE0bg7Nui9frlYoOca0Jjk+HpK0gYysHJyE06QWew3QTcHQ8lsswi3YBEX8Sjc2Uh2Ru+ABEfJ7T
wIHursrNMW7KmXQkuyqdVKiycMDsYsqpOJdY4JCiUByseQUXm1VfV1IjBprugEM5mYDsDdVnnvdM
CCZ7VkkmSQbmiD5NEb27nEF9ODQNFKhAz1HfXnqwzlVlikRHSHbzwrUH8/ua479sGPoU/6OP84B1
fxYOQCNw2NAMSNVGBq8tveSjdB/nkKnyIcreTKenFA3AdFay6nBd5ahj3RyCaRxs9q2MYzZ41Mc7
A65iQPrh2UcFZDgD7M3yJOhy9GGTY6X/pl6PoUwYX/qLJnXVqywqpIMD8U1e0jOyg5TNM4AnAc0V
+nZPzoTFPcocO8AlAuDRQag3WZes6ca0Ij0YaqVe/bExzymHVZeK/66KIi6EHV7jyqLbmFkn1MLe
ZCR9F9yVTdJi8mta9Fzg/eCPD04HF0Fo7lQafr81uF3urFAvIyuz5F/pE/MTsSwzX9h92d036ZPH
n4XRAwad/+RkSDjkBtiZsoRubrvCKKmzaRS/5b/3B8BP8v7DaqW9bJE/yCApKxSuDUdswhwgy7bx
BBFEyW/FvjDWj5K7SNaZeK7LZWhf2MaDUO9234hd9XPMBIevcv3O0fEVeDF6eDVYD3fgspTHSL32
9TlnPk0ZxT68ZLksR0K0jD9X2f3knj8HOsQ6kVn/HRqP8up3wAAgeZwwg/54a0zLQFPOJAqljR2+
ap8cb5yMr/0+V+GzpfxlaktjXCS8Jpr1z1nb+tw1PTQ7CBYt6ddrnQL8QNEOMd/Kbx5rcezlSWn5
5f9hnQlkd5Yk2TmaLbbKjoUyPbirhNSqoJSnmllH2nOxCAsT0nfsPe9yQr8TC6ShQ2ASzjkPbr5P
U3cMOGA3Xo+iq0ffvg2eo9pFiBwEJtk5XXADeCZfAGJUFUh4yHLywHITOT1knAcDxITnIH2L5hMC
W1DN0lqpMj1pWLmnDnw6IE/lrhke17rla8HkIo4hR8bHdQzARMB+PkZ9qSv/BVmuBvQA6Al4dNB3
S73pbffxOScLO1szj4h8KvyLJYIvQojMb85nw4QCka7XU89LKuKgH4S/X1YCVQmQ6Sc1GpKk0Emo
rLQ2lhvOgprcltvIX1gyjYaYheIP5Lz9pFENzG06FQ1B9/65y7SDAEW7nWJZluoyLtvjJUzj76Kh
4kr4hkYXy5T/VriC4wyaYWTqqMMr8mV7L5N7bv0nuHn5gYd4JrvrHanv0z6srkKPDi/NGPyZY8nF
ZdCw6AlIJLfkUdaRUty8QHcyhkJrmqqX6QGGc/1Dd3rzgW5CtKypiWAdEAmi7Kuh3anz6+mMM17q
qWkSWnDXG7pBpz9FA2xdNlQpkeeh4ZRobB5O1xbqJhLopCIOa2QCaqLaP1SfQSm+JkbrsZ1JTEGE
obPDuRVJOFL4cW6QSaH4TJFaeSn8lm36Ht3DlclXiSYyoHjvpKUMJPzGYeJuQoiWEH4kW2oiIs4S
21kGfnC3KHaJWsoKP6IFQibfGPh62BTB6CqtPWFOK07jFOOmM1r9pCtE5ip4iHnBEGhCOJxZuTrT
VmYA7HNvAeSVi58UefjZByr+0xMEK+svbX08yuJBgHpsHsUBqB1PCnb0p1hjnBaTi6cyMkDqBM3a
tgnKK4KVpXCdncZ4LpfHYK6ofahDUFcpYFjXcmfqsVU2rg+HQID3IpplXjVHqt31FXcar5bAm2NF
sNgG6E6gkrJzONtew7k/cj+LU/kmu1cFOQqKrHu7+UOX/NYZOV5adnUo/KU6lN10xaEw5m+EvdWz
s8BrV4ImhqzLbTcnmkKWZLQnxdhAduEFM6916BQk/4Sk4dk78lsC66YlOmLhCu+6vvsc8yXlizu4
Y4Iy531mUfp1iMmg/ttNeEcM+fVe4CcrA6LSh5iEF80jRPe9wSQh769egyMrNYKDrM4+/UP8ZMXi
dztzZi1+Loq5SVNjjQi7KdyWTmQ7rCmjQS0TGbJerALeXF3SCiPM3BfrMcqT3H0wB5H5XAzkFBc+
+JNZtXrxsrSsIu8+YwoFQPho97+NvNOqlgAEROzIDMUEh5sUZzCRUxhVklkfY5EIIGyfcQ1iw4ha
PPInEP0fVP3u2ifmfnc/LAWvSPN24l3flHUPqMqV8nWa0TBNF5SGn1TaJJHW9jvTjLdw3ybufgQy
EMfSE08LGs5jFhhAPN8J/dr2hCMJy2lF+/DNmE9pgAwcWoWXtFikshOc43J0FoXqU6prXvSwPGX8
43usw6H3bnBw8bna9H2rbrNE0PxCFfudpDXt4edAv7ZpdSmfH7xZ7+ocnyeoS7muqVpE+xJdJIb4
HqPlKai827VlZeJbmZdzqHREXDx9zcrwS623nfZJmBT896/zov0+uqP9F9hlNAKY4Aoz0nekTOYd
2qN9Sf41bB6nMlETrYgnc0J6z6NOFiOIKRSYk/7t2oll7v+1VCAv4/qUBINyIM+c07eYMSOZF70N
nQlUrP1QUUy1qoMx66hyDxoTVbGu8ADJ63BS7eMkRoxV1f2rKUxV1bPsSWVZYkQCUpDFJVPRF+wP
gR0R0d8E2wNURnbtKCELVHhNZzxHCWMLxvu8EKwnnZFV48hYoMveJ1TzAS4+FCH3dlCGbUA/Wg1T
wOJ8Gr3qGRewgELvueHhfVR7phto2T+H+i1wuQCqaMcYYPmy5S30sHArBlGfSr/v0Qg0v/BYTrLj
hGgjMTrNamrxgX+366AdWCFA1w/A5a8p0Iapv/bdaRkbLNSoygZ/MmvLhlVDNanpM3BsWRDHFToW
rmlF7SknpozXML0xVt5FkvIgnnDb1UahAIminB/1506QhnacDk85zg+6/8wp2tZWkQbmGVWe5ooS
F5Hd8XOD83Nlvc4efNtrcGx0fKiQytguQ1pm5VLDENU6lHmax7cfvPOhegzJhTTadi/m+zJX+u1/
bXZp4w37L1afX5+ROpYtbWmpr3eRi1r+ZVrhbvGacG0V9h5mP0u4j+fvObHivPfevKX2btL/89YK
ZE0I24HWZX3jJw0Zsy4hKrAEEq/kpiQ8Y48HarsW018/kVyzxC2wSzZ1QjXX5VyQd4+sLgdFqfx0
9MqMwMZXeG6sb+zgY9RO5f7m07ip7qapg5YNf4futTGQpcmlE9/kcSK5L0t8tWRGqNPUVPM5LNEs
dOfYsyVPl0BxD0VmdjOHUgqjWmqew1ekuzwqfx+2uN8DK/NNoCqXNthneYeyhA3Bt4svoAX53Btm
Xeajai00AJzIv5fZyCsX39m0fkXYlS9X3KAk1KGYOQlxkjUvexX/Qj2BB1EgC/0l2p3rgV1t0EtA
VZJj6RcFFq7dRAwtmjZ8DiW8MEIYzAr0yKRJ4JsIsEr+ZlRrCsl4Lbg4QzUbpr+aENjSacW/Q8QO
ncSGyUA9/yreA3+86h6UOte5Guq1ZU67ev0TEOxblTWyUFayllz2gpRWVZUkgPeVQltROZdqpXsb
b1/3Trs7VaM4aAeB/KjM9KNRbO5vxQGDePPyKpbboFILYLWKVK8WAYgK8peZ5/ZcCXijTw3TjgpM
iv0JaoIuZLWwcOiQp3LcPoDuNfqQuiIEAEZ4v4nN0CeyogfemWYmHd45vrUTPABsXwIr9wbe6wdz
qJGBxz6Mw0Ncs3pToBTZGp6B2uiGfPsIkHLvNHcBMFO53kffsHPsa0coNYxUXPidzDV21F5VvoMj
PxMYRjKYea6XVOYp46gikZZToq+DtYnCvtnp2ymHZr4id/7IjxJytp+ww6UomODE8qNpVhshWVPq
b0vAUlALo2/JgGyfu4ZCwIurx0j0zb8XDq/1uzaMUf7+JA1KN8vTqwa3TdrLYDMBm7vMrwIysDgd
3xpQU8Kx2T9A9FPtegTridb9gc4QpjhRHbaAZlMeCIWdpuQMYBN/1oTIwogx3A4Mpw5WHv6sSYR5
+3AGDDaZOekqbpVJCtftjrIec4yJ+baMw9tDKIs0y6KLCLpJmoikh6STSGyye5mSSuWG/nbJc6yh
GxtFEdBYrYfiSI496lwFGeVprucDzYON5XQeWAfrXdS5s+eEl57gigr5ZzqcfNOdcc/0PAFfkxOo
ts+JAeo1tBtMdd/FIz5cJ4lduY8RkiygEnUEU3zqG6tBLaRYUfPRyxKb0sgAmSpFO1G2SSyLPZ0R
fsA7LFx/cCVXpPVB6YPCKAmahh1ImVnIa/afc1AJ3u8hlSrIjT/PfZ/6QGV2gtCEB6QYfJ2Gntam
G9Zb3H2NOg9gihQFegL6+/bgpZHILOTmzJjTloO7kgfJp/jJ8uiR4Ob4Kj2kM1BF5KmPybY940A3
iqaDb0fFtif9b2s61q4SX/T2etWwMboMqFMdf7TlFCptgzEfC2sev+tID9PLea4ZiihBLqnnTRob
3D3pqjkCx2ZnbScykFuNAroL0+QUhsWWVyy0jskYcARibJyXDa/Z4DpTaM5eOGyu8m/AtUY3xkym
bDzFV6+9gfReRACpxFR8DQbCmRJvFE6kFGBtA2zZbAlNMsuhaW/AQ0GPVlNzEdMu9eScO90CYxFg
9RlIi6rofcO7553rcsSMpU+PWfExsGXgbORraaMAOIgYspjXlUIbceKb+eU9dd9lJHSl6T00RPVZ
8+UCJobQExVFVIQ1DEUa8D0ibG2oorJX2MWiBCbKIlIQuL1vCGX/imUrF0B3gZkS15CukkKdJ694
1DluuAu6bkWKUcSYu+sPmhlkUEAJs7LuStKVarL4nfXcsA1k6IdMcJ87q6Nxvw8/7P7KiP9KRRhg
CuCmBlnl8vujM/isvMKeQZXTbaRlBMuiyqqncZ7pa2HYo3K4iFUrw61BUs/Sc+7Dq+27Pk7jlm/1
REuQWGZIaqavKoJ+EUGHYJ00En/PE1FKPwgFWBLe7ypa5zxih83szhvyZ5fv2KFSXYqRuimY9MDp
ol4SNWERC8hom0YINRgceacBxni1Sp4yA7LeFqNPxInASC+pNcyprnx/A2hFGm5Zuyknuqx4dPUa
vx1oke5zimZ+SzY1rj0jN4pWIb7LUHpoO099mZauTRLKtDjSPWDGl/0Ipi/V2rGsoyUKToMdZo5y
AgeBl/rl+nXooupZm+bhL0QPPACK1LhfWI4F6Pln39rOugpqltzFegvTcF1OQadkjVaynxxpt7gx
IfzXVp2PajZhDaTgfeblkre1Vcovdk5s1FS9iPWcJvn4FWjcvF6mu2lqm1C+sbzWguuMR/ogc6n5
GPKRvJ7CPoibCA16u0GdV2xewm35Ba6mu6CEKJLKP2LcDFNWybpjbGoFC6+5hj2wNrhH+Is8Wtcq
lnF+fZAShakI67JNFVFhRAA5rCoYJgV86k0YRmE4ijD4jL0n9GkOurRxJ1saractfRI7vOwmm77c
4yun2o7b+TbOan3cijc56QlerFDr+CaDR5eEyuT19sEwmKM+cTK7NjfoWqWFsX9DJ6B20kRQ3X7p
xKpUK+JUx9k9bPIYSkShSD+d70IYggYMe1K9H6Ebxg8lnXr59Ti7JaL6+EDANZlcaxSNXFLmypdZ
MGhD2X2vsPNW57sceK9C2278YDyNg3vAGhDaa9RuXnK+m5i/KeiubkB6q9KpEavhUaM1Surad79k
N++4rPGEeZcl6gJEe8qyeGdZP22q6a/LZMm+ng60lhSFZsuwpiIhX7yBPuzsZjcrolb6ND0ezllV
9TVFuvuGkrgo1LYN9IpatrtbqtB7IZzDBKx4czsXbsX2T3K9bjvzH65QbQjgoEqZe9rEgg/qiI8O
7/mxWknLuJ+mU57BbqDNNBdv9DH4NNPLEydt8rW9m9csMWvoEPOwGeDjF2/oarm3coKFmXujjgla
ht+0l3Agnrfx8aY0XU7RkEdwc9XkWbA4979/rFaMqgt/kTLPmsY96lJsl4iypZ5jVIPtHZBJ6606
lTJghQaIGndQ3jsuC2A7feJJ1EptRJ51OIJgWi1jtenZzPXqB0klPtcFxNQtUhEPLqj6iQtXslk1
6AHVyT1UOHgo0bhkXK3YaoV8Jv6UO1W6IgOeTNEFZj0kHYRRoGHnHKdN15vjz1Cu7WBgKBQ/dAY8
egjN43/5Yy/wKcaRf6O/1nnU1KVnxDXaqDY5yibAmmi3rWQQyBNaUi8fxOYx6ybCl02bftYeCzYu
NH+RgEO0RKfz1uUQ7uJf7Dr4aEHclO4oVOhIb0zNvdz17ARg6hqpg/irnSFuIuw0zP2lHGF8/j1g
N6BBD7ZNF69n7mipN8grGt8TKFpfWhQaP5SA5tZVTnQOx0VOMHMFEu4nuugLzBEMpbyqsyrr/BQ2
BCkEgfFT+j0u62B5a15zfObRT+3ITBtRT01SgpazvmOaHFqwExkOsa7KbfWfzqTPRxCxP3PbLFty
711wdv7s65uAhQ5YETKez5hP/32ht+iml1PoJZFmQQ+GPmnGjlSur4Ey9NKahhThPawUYbHCTKU6
EgyYigMZJAif06DQWfSr0qb2dhi01AreiuxW2cQOr02s2JZot0t8AN0tiKhZsg102HmKXNHsawIf
Y94TfB9Gn6OGhPsiu3BD+uMoGxP6Jc5GA1LH7hhB5VtoiIEL2na+SxRHSptEsPavqC4x6nrUbhY7
+N3Aa36xniUwwEGT2/WO/ZTS9+DgivG+nm9pHlxpIOcEsP7CPvvdKR2ggfcBfc8d5gl42a6zEKGT
PGI2k/BT4xJHFi8hxSL6Llo3YUVvbmNrzyT3Sd6Hc2ZzPFiuUP6wfg0W4hmESVCboMVx0EDdzE5L
8f74M+K/9Mjr2jXJ9JdtXvKWXQagCsUFWR5v/Vsb/F4AEQGmkpx6RBQ/p07Q7HTkD8l7sldsIHnU
Ic1P40K+ZOvFoZNMWDLIAlYDmB0Xe60gfZJSqZNQerPR4UhY7LvE3U7GuFRllYtDEKDk+x+E9BXu
u7W79WasYJ/s2PVqqtkxQ61skDtJ93vN0N1oJcxu7DL0FIGRnXpWQ1m4wcsYK1dXavmkuIPBdGqS
a4ni+65mh4lAN+6w1MvJzjdlGj/WJgrz4m6KDMIprXTigUvv80f/BpjOVfvLW/xVXSIUGNdCSpWY
f3fdiRG+deauYQe3dPEymfU8hiNVT8lyVaCDd1eY9UkSYXX7Rew8UtxItrM1Ahd1Fxsil31MMg/D
R6lvXkW5wmhGdCFccFM3CcFD38jtoNONIT5VGMXCwOyefEAvUsrd0ou1HogsQfmP+gJcgIgcYXRM
qkWTiwNSc/s/zBDIW5qxhPwdj43U+wo7ewjm/MZw3fzpmmoOLnUI+Cn7Qz4VL7xnzjkKSZ5XtmcB
+y2A82+vJT9PW7/j0M7NA4CsM8jqhW9RukzVAYij+64+IoJZT3cSugsLPGxERIGTDDPXWJCHbwSO
cLf4KLFgEjZKjjKrFIBkid1sxRm6jwRBm7ONDP4aHDEcuV51oTIIJ9o690zUosf9U833KxiJZoTs
UKl9/8/olMcAT8GCciGFL5b2ujMzv3EpdJ0/+CmL+ILK7jMZmMmGoY/LE1an9F7uKujRHPAGBMEu
qadgPZe4culw372asSYUfd/XRDS6aotr0cUqsHMcJmxhEujoRyFopNZO59U3xPAPi/xv8iUIFFwp
LuqUuAwU2FAM8XHfTeoz9aKJkt82gscBNUV3XQ7qkFmP1/owbDQ77lv2nLP49TmRHISCVZZWaF3C
S5mV0TqiWmpFPhTTxQK8uGvWGSUo93jQRX78rZWTLLfpOqd++4F62WUzNct3YU+kGgwG+/lDScIl
1qaBeVgW3DN1iKFG3IEU5PIUJMMIKqb2Y0XMkZ3eA68Gd5mA7K4buAnBohLCHUifrOlksBviBpRF
Qq8RG+82ryPZ5zh0vHngM+8XZ5vqdcEFqHGbefH5HJbLJHcM2jovki/lTLGqrALO4WYlG9w6i5Ac
KhDCDNAp8Wjm3Gmwi1O+aRO5ShjKjcaOdCwamk3il2DlwrQN4Bg2p1dzahyLACpYfEigLcCJBwuI
5e3iOWSXzY9Rq4YRt8d0EgpqWicOhq1LClmaGkIWIikELXNydFnt2kWHTqFk6+bpqliQWcoFgDfa
TtU4Ed2NyYTKcv8NMiTaSnCvtvNmm2zNUXok2zrnlwetunuRWpS6t6l7+vphu8IJsnaQOxo2U1UX
VPJQT0YPZhfoThXe4M/3tNRw6v3rTzbN4bnRQP8EJkaOXp6it9tt9hAxpDvSjN0AuPhYf7Vb06Vi
xDW9hfgeE6jMGBP0oreuvkGuxkas+Pyf5IMcRPZYKB/h+xq/uiLVkfkaghdC4FRyQqVMK4CXRndN
ALt5u31sg2G6HkUmAN8vRs5yvXQIzDASynCRtjvq4/N5i4umOCNvz9WdNflJ4lalvSNS2YYBY5lX
jl5632IdlYBsoxYLDh0ZTM+i/fufiDROhbUHdZTkpsXet5GAiRz6ap4DjIg5RBOdSSoVQpq/Vu/E
PUtEu325LX2UHz16o8z+MrkpwVnLufIBG4vbT6h/grFmzlgJ/3SufRELsQidPXbd3HNWxhrURDHz
Stm/60UXKESiFtwGnbMUJN0Cm08C8sAbzcblyS2ul0A6aTomUvG0UlUtmkA5efYFziB78Pl3ncjW
Hd4u+O950FduB0SE4w5TFWhAQYDoZumvCgAgCi6d86II7+rFcAjf83OSqOyCl/EvPslYUeiXCjSo
5lS8y2TVTjIN35sM8PAMdqU7JKjNZOMmE6HNsmJagrWLJAvFqQ+N0dCl0b2xLTtA3ZBy6dkkqesr
opyKXZE+b3pX1oUSripMzJ4ZGC4YRvnOPrpqApR2XStqWGifRWFtk/FxaCB77k0K6PaXjzShckxO
6Bo8LRHxCkxC6hAZxzelulMo27+g70TCy9jD/5G5eX19mrjYpwU7L6OxSJG5t4O6iLrTS+XO2GQ5
Ww50Iag3pdc1qDQdjetg95SQ/u3YlyVWhc/UnapxPHA7YUe+6nObNc5thDNj3hsTqT0WwUrpyH4/
u+BlISAbMgBBPqDgQF8VrmpmN8+tVkOMENQYtzlfnpD9gpzOn43lWhzoX3CwrV9m+YTCNOpoUfE5
s/ojUI9Ub+jAVKznjbxKF+HJob76i0qGtIdmZtSAwtOEHWuAn1iT/lUIef6UJ3o6QFSz5C4VkoXd
Z/b4pSWqcjnrplsZkIAJ0gSaQyWChrnGncrNHQgCyT0QcAGyJtjlZtOvPh62sSKRGkVp3bZXmSf4
badqPLQ0iPuLtn6cefE1SnwVzxU8ci7JEK7BFd4qeNQxiFtXvYGJ+50kRsmpQDXVihxNJqyfHx38
wCTBsq9rZQL7XZhgdPm+xJC1CI0EpeY9bxnHVz3/VXZbLpalj/WLOVO1TclYcGbAMkhdhDxeNRHM
/UcdaWRV8ucNEfwCQVeSq/OXk6doWUToH/95hNYlIbJbx4m4dRw5QTj5c5iu70Mj2tXlWF37LN8M
sqp64pEdwSARE6CelxetmADwEYrCFcvuLiNwX1u98uwxDYj/9CtuG/N4USg9iNWLksPmByaXs0zY
94il1S+FsDbw5v+cMwPfDy0832tdguXlBEcLOfPec1+zoGrV7G30YUFR6go4TkQAUlnTf+O+p331
bU7YedMQLQhPBpf41cFkrWBKguv7bz2ubUiYncVdV4qjhLyGKrySnSH8lYH91R4U4c+A8K2pXo3r
1FNVwcICldWb6/4syVjwlmYd4k/7O7IalYo/dqqVGZN87UvDj11ywWjjuKkQUcrWYaZxVI7n+VPd
QQZYfZz9UH9y4cLB4AP3Be0uSgBFTZxOK546q6tZ7Cv78NEJL5hirwsRVbtl+5Dey4nOtd0ssWwc
TTOVY9uuTxBCjnhUZr43G5JIgRtwTgKHW2ZVtlpwGTUH4YIrFLzP7MaSlfMftz95Na7c276gXd4A
o458+fxKBBUe0fk36w48Z4Dl0HCTuc6ElOXCljIBYBWAKtq/oAn6B0lyBtcizqrDho5iSEAUgYkt
qYqPj94MRcxtEA4syuDPI+6sHSdQnZv14tNZs9Fbcwa15MUT1iydroFh5z80WvU5Dbt2wENdUgch
okpsU6e0hfGLhMWKUac0mZwp548a8NrfRyRC+fm8X5BtavUTCXqlSVUmAVjNL8c6zGWrnwJEGTNo
3OYylcb06ON4Ho5oBgdF0H88aK4xexB8uxOc8joXaiE9A2P0rBUCIdIaNJkzyDp9Y7NfSEKEtEgm
8q15bKiT4Oe+gFcs5+T+Uwwywu04GvaiEiJVL7o/TmuAk4oRCI+Q8vYjAjYh4+BGdhLzodB8ETYM
tmbKlVnX1948x7WCU8OfHIPQTqJQIDsjXmKMrp7ntpEStGZ0ziDZM1Hud/p8ZEqNPc0CDnJdgqf4
KvwEETEeKWkyXzJEcxCjs9wPJhlUKNDRSPGvDPywD3kThS8r0hbwc5UEoWiCPYEb8I9mF6QZkrBI
q54+09LwA6j269tMYwySRnXCDyqVEWlkwxL/MyOBCsr5vG85HcBQCqFbypluVuNOdZKkv7VbJo8J
F0HSsIKRKqXOLBOLONLmplJkSycejyVazNyy3PuJdWmepSv8Ea2gdZXnW1Xo0nuaVXlUHXNkSH8f
36zYejToTDCXIi+7GNNV3udiiVmDBoKGqcL/nyb7Mu0rYhX0ol2offYvURIfvzB9pTOfGhpcU8il
0Irf7yWHt46Ul330329n01+t/tU7ozGzFhtyG8Te0bNE+45cleEmsZsR8hMgU7KK1nQ3/QmSJMMw
LleLdbj+j3TxclFQxUKiH9GuJUNav7EEPujOy1B6Y6aIP3H5mn76cJcnUixeqGJKnix0t8oZtLcE
sN8hRp7lVV+UXl8qHjqN9fqsmT7VMWNcqebM7NCh5ZccGnpGAEbAEGUkw+lb+sd0FA2ZnqX8ZWsC
TqjbVuAOP7nTusgyF1L62PuBhF6bhu6pPv+ZDYCH7PNPkAJB9Rtc8UQu5+h0E47XCtXuRi8u3xoD
bMI0lJ2PzqO/J42xxSHhM5WpfN2t77tKoclp2PbcJO4I+aX5I2dDQjYBYvYJ+QrUooqaSeKoKl9+
E8O/FUTVV4JNpLcSH/h25kVAtPow3LCBPx2frN3uTYCkKF5It576ylNrJ/z2wlTd7c72ZpEjT99p
gCnswtbNZgGd8yNSbrVldlSoh0MZ7bb2w8Xd8hS4/pFSJtvB9Ra4QfeIorhB5+jeeGUpKYa1MbsJ
ZlxasUTtJomFvnzZOIHJIWzoYgB1Xyj43/k5MNLFGzBaXyy9Bmm3hiPCyO4gRKHZia3ocj2yV7xG
wgic6V5j9RO82BH8NEJirqDpEKun6APJ/wTEVndJ9W7LWyYxZwtmVwArJKQjDOwAGXGxrOQMXnmm
5QDdPLYATY8mCqjnfvxO3tx9U4roY8IT/+2UrI23jbLNEXy5mMHlo5BciD2vTewE8/nKJrPA2vv5
Lf8L+cbaSPwJZt/hFE85c6FfqYGb79HpUfW0zt1nh2Ja9yZ1YXu9PAZFB3DpJ1v9Ty/aX4PI+LXm
ouUw0oTnYpQeqQ+c3ZeejAcYGiHa5WVMaIaQDghXv2PdYHWNAYtint4ZWLVvJYA2dk9B5uRlyRgB
bskp7Vh4ocAGD3LS5LojXPx7VjsShxJu4n9nz493XLkIm5CjCOwbLDke12sqqLr/dvldk/vbLBRx
6yBSDxgF3C0vactjxQUw4r6C51F9+EXr7bPbqOAyS+fe/+OJXG8c+cNpZwAwtN4Ds9+7P8fldwKK
l2VWursO+NAonXr19VCxPUJOE0vfdNQBJjmSbBDtA0zqEbUBlJRWxG2tRaJtLkvKQaT+P3PXfrJ9
5pltYqM7Nj1MJgNghPbk6qIjYMMjWITtjWstYy+X8hVCEJ8R1snt2rbmyIBKoq83wrZltP/lNbHf
i6VtozltWlLtatECA9uLemZ21amfChrvTuK7mCeiqm774LI9fsZ8pNZCnhpaYJBgTPRxT2HD3af8
bw9CSI7/WtufDQHFuTvxBhZQ4VkO5zPPAbyjWv8/Ae1sPKcoCsnhgkzpnilq85jNr7JONDUPDs0O
AFsHeQRng11SD4msBi9GNV5PxG7Oi9fpv9mbvwU1F5NHFHj/QUYNrrQe11rhHRTAB7N2klYYInup
JHWSN5lUePYNZc9py6PHvLF6FOH1k3n8qYHr3O6fVfzQoEHefkGFg3D6olYRw9p8zTt/9a5lb1/Y
ohWXSDYUetTyHYiAuSWvXlz6DkVHuBMJ9FiKmWgQRyUeB3rnbj050/nLQOW8yEuZQq4lPvH7+/Yd
fhoiMSDkZld7F0DhpL0aPCIr2G9Jiap6SADYppxq/d2gcGTjefyczdAI1v4YDKV38cZfRyvvcvd/
MblET0ePS78ycyRwzwCEC7NWIqs1fMb8O1a+XBNnQRNL6GkKvVd8Dg2mEfJtV8xawDd8fTA4At5g
elY9I7NDjACGCcVGnoD/8YN01qQn1tDrVKyjrg64tStGmGgkXy386jl8cM75MxUkP7tqWN022eYT
aabMltIdktAYmkUmovb6NwuifRxPRbusEdFUyrh1bVAWWfTHbGYoeD1fW/dVElcFsKWwos7Bcv7z
hfVKXpxtZlw0KK8Dj/cEKQgpO2lqJM/rdjyDoKwwnrxfVWOda9UgGdI/53Ew11I5GI89y9yhRTG8
XAO48QLLqiQ6r+NGYLX3a4haKnGs9ddiNjmiOO7o9iJqGUwfKzV54/n6pmjEWTe6pp8fwy3mFlmy
PoF8qjqnANmKH4vkacNrDeSpprxrldYvGxSE8S7BbyjS90HC65pgN99vjkyqzhlK4T9m1zig+lJV
stQGfBSU+t+UeLS1N9GHHMkM0LSvpHsRvp9ksClSxibAIaExet37HDD7E22Ln0bkHrZntWYyfkII
Rg5bSrIjs3HQ3861itRPhA6C/6vA+dtrtejbZMW9546wP8Z56oKV50o8Q1CGZGhe1zQ5C2ngdnCu
tjUlpxzYiANI0kgyMwHgCoIe4grWHX2HwAYczw/EEbCf6dkNwDu/G1oDLPhSTEd6E7/O4QL0927Z
5QYlYr6AfABNJHlh2QGy+wz40lfUIQk2z3cIv7brALoDMilInzCz9rNqnQEA/n+AikFOXDjCuerA
h+HIxeHILOSCuyJh3LgCcUYo0kaVj0aGGvVHJY3Tha7Pltb5XX1pcLklVChfhdzwnvrsfGvUorQy
DQetBYyjMrZ1b63NXa9FcsRqeaHg34xEGLN4vz9tJzWbWKsqjy04UF+J4FauC1oRAyhcx/GPoVss
54QiJg3P3HxqeCECuHKSndZPq0FjQKvmXSb06CFx9NwndhwIQ+OJ31BMxRU/+WJ7m0B9laK4n3NF
Xn5Shyncm/uzvZDHibrXTbkTvejuDeenWFxR0dB6dvyp3UbiqKfO31ePdHRbVpXNTnqdhSYlw/Yr
uFquii5ecL+17NYWjP2Nhu8nEbJfnmcvhbdyczbsY9M2hg9iR93o7h4J2N+xQICtDoNIM4nT5v2E
bg468mNwVqUE+z22SnA+poCZtda3QUXrxo121LYXoKXHrnaESHtwLoO0eFDHnp0E038rymnn5TJw
X0/2j7Uq2d3RaeYgOJ+VVOMkYXwAmOCS5F4vO26Tw14gCS/lCTVNHcICd025miOAP0RnykedzTFC
GjaAaYtlN5Gj8Vz0MD+Gpw76sd+g1rDY38D0pyhaWYq6YNEwBe6/Kwyr9I7kJIFaE7hIwsO8E9nD
uMG9TGpoTEK/1iKUshaWnbN22CQHK3NRmQ2GnetQ3AQZlk2TN3ZQqsrShWplE6yoCBjLZrAMoB3W
ED7BPDZqBcD6iUozqPbGbn9hu4yHNhj5p61JHEIDudq8m/BGjkracMtJH6d9eFFWnIredJaA1YJn
/tlj9Mk6HXojAie9vWZje3mzC/IUJu3kv9DG4oxLFVWmctEqH/i5/VNwQMpygTV1knWJvkNqyXZm
n2nKRUYyqlrQR6wuirkPHXRWuosa7tibK2i8Hwf/lDkbUOwhP2sFhTvcHgSDwi/pzlsyBZJxwQhA
C+Apilsd97mnKY7i6EF/Bjh8//79cITuTKHG+bNiAsK2465FIlayisjCGg3u29A+0Hkl8AOj/gok
HJJrc/Kvt39byUb2A65HAUOTbbRxkTnrqU629CT4EslxHUZXUJGe+AHriiCoxTG0xBUKE8GQPNpl
D7WysLxbY+oUICELqMe0O2suecHpazORcvjW4+RKwa7t4JUnK8TmMzrEfr/xRBw0UY7fdxEdjnpg
p432c3PqeV/cXgesZ29wOhIP4E8w1TbXM32kswXSjuGtD/6s68llDkcZpxM2BgubRbzjyVKsSeXi
du5stI9uDT7UU3M0zWDQLL1JJl0uO7HRTo5WmKvSEwoKWY4cPqhuxea7nz1WXC6Qi5zKG+5QXrTw
PeAdFcQ67V/ovzP1iakcQLikXSjPck45L8lJ43BdFMSWH1cIPlad5lNs2g9KEDM2ZT/IjuBbGjpx
x6DA1fyeeoV/cEhOKob9g3jaVlIVzZm5kXVqOaIuVMaWSbJRHrvUCUPRo+ntH357wNoSQDuNkxli
eGhhWR9xBiaAGdI4A/8+Fr2j5DtqrLV87wzm5EPJXhxBOMG5aeMezAxHe7uLdnNt3z+X+A7Q2Z0Z
A8W3wtoi1yyS4QnJsV4ImAzha7VhkYVeVmPC1IlaGlTlzBp1JATW9MO5Mo0jH0oqkFOv0olTHoPt
gWiLO2Nz47PIhHQK0ZSW6ah95pjWIC6dZSqVMA82gjaUztFfjoWLYzeTotn5MbNIzo5/BDalhi5b
ojMUVk7xBx83yfEwhgi7ZHDP+djrF7Gih4B84I1yNbvjW4smC5o0uHJQR7A7RkFA2/KzPP694dZR
JRXlpY84n7V1ndZX9HhPcfFTC7yKv6TV8J8RFqSfQdY0EnQO5tJhvF9ynIcLeYyCRqzpVq9Sh0zz
eF0XPIiukOQlncC3nE9MA+BeRHGqWnVVAcdXplfgKHOtFdw5XclsUGc3Xau1o2hMxM8hFnl6MeMj
pUM5ydOtHrcZWJjx+KrmD4jXCThhsi5x0SyhFX03lkxt7OnDXHXqRor+EKe2G94fSJ5OveizGtFh
iEGoB2QWzAfaEVGZrzVfscXGZZ0L2XP6OgxCM+E3xX5OW0bZGfhvInpvvKaWIEtvGudMtwYI+j02
irRKIwXk1z4kfEw7LNb+oF8h9qbzshO0LExsJOZYUSGK0YYCkbb7K/viWt1B0a1mee8s0ZE0y9TP
iUODZTJ7k6nPcuW5FiS4zGm6zhFGNg6m7XEISgI8T2ygfty+z0I+gjqp/Fmi2Vxgh5TuaGByWKbI
mvVHwQd1Bns2ZDfNo/3vp0bK7rZ5Z/YeW2lIV7JyIppBk7JiGAsZIHuRzX4i32DkzCvzRsr/rtSG
+2y9K9J18iLtPL477ksMKRIs+bLH0EvCbSJhf0c0btWRAZwUyTLmsZhIvpijLqEtNYijxka84pPI
RwwzQl1PUKf8fnjWRL199EJWFt7hs3TTokox5i+KItrJ3vFcRrRiMvSol0klpMDrXcAlDfDZCOvk
6++zsy7zVCxJr6RJCo/pn7W+2eiSyfBMIofltCMmt7sFz0eFsLTrQ6KjkEBxaTJmXF49DHfZ5FoI
k3skJFYA/1/1DYWrNIU4KNpqVwp7PmsLWETvs298zXOLDeT52GyCzROsnR4p2B6BtGWwWnqG9Avc
uLaiwotLX99PJuxO8I7p+IoqNZZfhSG85RV9IRHlGGpI32b80vvimHCq8ajlq1HnvKT6KtQXwh5l
nmnTuuZHUYix2rB7a2DgmxU5/pK0nfRsbuSwHecjL5QU2wWQD3dfh66W9QMLnT0Ead4yu5koBHFk
RZtO/hXon2ZnTF9sLwv+5zbtsbAMzM8t9ffpyAbnd33fEFWQbIQTfh+8zx6jwD00EOHVc3NVO73H
3Jmlige9NyXdKJMcBVlkJYCfL8SVrL6XXoWkW5lHuz/ekZ2oErvxbGcn2JVUwqNmwOuFOkaBjfRK
6qIdeq1yTyqBpf1DOEkK89J5ZBd5CsDdt6XQ/8Nol7y4JdIime1FxYnmtq/XSGrE6PZVwOSrqMQh
90RNGd9fhG7QVETw+uABbKc/f0d8wTGP9k2y6fupP6cqGvlLQC2Wo54XqJ/ir2ZsZu/dALpfGIbP
gICd2ZHJ2YW8+fDgQ6VcJ3PRJiDWhxtbZTyEZo+mzYn+BnfkNePD8evYAAPX7FxIzmAYSTdcEXYd
Zo9QUNU9ANdMHYn4ClSSNMrOvLyHI6YcEpgEE8c+LRbgbMCbBvikOxF9tcoizpNN4Y2SKw/dp7iz
MAYT/bhDYhYGHniJMkWr/MQL8ecqti0zYekwWxIjIaQVqLBNssrkJYKEsKh29rz1fC4/K59t8q84
yjwaIwk4sVthb8pa9jBAP0sntZ2eLwkF7fa+Plli/V9fL+eJMBXlnc85bkjOeIsn4AZKtTUEyuZw
JiyUbzVvOIu8iSujcn1/++OTNYOyqFmoQjosQd/AC9pIulb/eR7nqqCVvBAQOFCFaBZX+ZlxSm7i
QFLy4LGFgiI/AH/RTLK0qGlw5QthEZFibLPhuVMGPGF4d1VJqyLdJmPp1g3/bMu/7egAUgNxI3P8
iVqOP4DlxiHESQw3fuj9m6FF8BwuYhT6jHvWuPaOVAwIeHrxg3iNXf9mNhhusOhsScRmTcGa+LrK
S14x78zTe5Bp1dBXFr2Ac2Krx06PeWzn3ji/FNz5xelWFCC4aRPgZ2wtIjKwKpvU/VhApF3ioL9Z
iSk2LbcKNrLEfutOeQ73HbBW6o70RVa+NfKUCk7rn6UT0xyUD8YbX/y3BgTR22m59Nl69xqij7U3
4AxJeSc/4SS2iEqF7ZW5+0Sp/m/g7HpUfQ0nIp6aoZwP7ZUnFGdLhAZR9kbCbAPEQ4QUp5T4fw7O
SYW3DzHEvvlim/lTTaMQ6sjree94/dvPj/n4EZZR6ytvSmNqPUbn1JF+Sq8DGztCx00O0Tb6hj8k
q8JNszz/Iniqk5A6h5iZweADip1cl3kcmjLdCb8NmD4oPeibd+nCukmaj08ChX2byqdg6YkyGoFX
+GvZSgO+gmI91no0aM11Qpr8CzuoOE1s1RaHKQU8rYm0y+e3PgMJ/9SZzFL0AKwev4O4zXjyiMBp
P5LGugqfYwdQpD2/7OVhCiJHGwV2W/BHzp+fTNUaotBIDoiOkr+/fR/6fgRcrLfLDR8l23/Bdz0r
Eys4XkoIaOcdwl5EhYWj/eY5eu3cyvbxcHvh9yIcHp8mwd91SEkpp/ij0mbEagn5Mx1dv8ON9/9U
a2mhpllMfFcgeDJuXbuJbllbHq4onLrodpmEPI9lTGVcc2kK4+JLfks594vbVaF4kFOQAGKOEplA
9hFGrCb+GhfYN6KOnoQProwbaTkyYl7vGSL8rqXqTSoEfTLJVfC65Ta/xd1CSAmIGFQST0Cox8um
BP74RKeHKTgT9bi8zMfqrNnhKFRJUD9AwRTZch3Zgwzqisjtpd+HIydqv81hTrt6ovkA00K+eTBu
0ngIRamfNsL6kd3v/Eh1RtslzjjlaRrBHMjCmuWqy121av00kamsDOQrWdO2zOAdFLWL2SCeJFGS
K7zIKLPmxfJGL8jefBsSdJPP46F0I0urAZipQRkkbPTsI4iCwSjipmJN9OM9kZFtUhfwl6JjMZSQ
9BxvoGt69XBxYN0LrDXqUv9wl3SYJAXq3w85h9tpfsHkYJLRY0qJLTbPee/kZslMEkUenQequA2S
CkwZli8uvQK5NIpXimAjv/TVAnNfyRzOVqVc4m3hld4lCePHGLscCS3G0ViUdx4IuCg94zuxhenF
8xDMsK4j/dPDLkd9Pf7q4VeTI6YZqEGTp8g/HiK7yEQR7pyReUMEYAaE6BzJtitwCvUlSn+H90hd
bCXW6KHGA03OA24OmWwzKj0U5o95prDg166VGgvY8zNrSQhL2UDzabuZtZEIJHD0rGKt/epRAGJ9
t/Hm1PKecufFsGUaVI0oJsmolRLuDVGamK9NaaPjKdaFt/PWmhazRBqbQLWIJ9hF+4NQ0YOyPzkv
vXGxRygdPIF/7sL20LSdvsDw3/A4GSFfm5IoKjY4RYHPVNrQF98lfut9LK2RcdYDPuj/Oy9uwRSv
cXfLeW3/KzTHE6QyXjzC6KBQloF88FZXAOGbAZFrW9zUl3v4SnJTbTnIEwaOSoi+NRjf3klqQz+u
L4DPzuxperkl4BjQ9ZhCUy7qZHCimKcbCo1iBIgEyE65TTs6+hRpmCoJItgXKGAwdRrje/eTlud4
ELwODdLAVtO0JWxFPa1tt+WdTvgKZil53B+yl5lU071IFHGr3zZo+UnulE3Nc8e4sAsUbu6wIZaT
Bkq+L3ZicG1EX/maTal6o4W6ZvQgUGJZWi0d2ych/mpDZyIjocrWafRE+yQ+6U2H2Hg1+sac++rF
sD/6mLKz01va56ctGWqTv2tfvgvwqrH5GTI230141NVPe2k4HmyS0cxXQ+9zWm/CbKjpD8ELfgo4
Nw//42O8sVrv7lmGbNKHRq4XCWkleDGaVHbmqUZZhGpBJDItk002B3MlIJnZbzrfU8X86LQebTRi
uD6zesgxBkNH7X/m1xzJX18+CQFdeo0kANstrU3kG/Wkw+4gyU7gJ4jqHlryEyb2GcWdMGVIFUYz
t3ljP2TbyU9hqYrGPRQr4KJ7K7B0lSBp6JFzQDebgW8ji6FgogGpD9/uoZy7xdcp7rZ3s2vTYK5M
7nqrNLTewz5T3dHeWdGgdBdtlJ9k3MCb4u50Rqhq6DrJ6fA98rBAzBi6Vx83K7WfKZmCiP8KAEDF
J/Vfu0jhg8ASmJbaP06XrSkoZJKUH15TX3OVTv4f2nE4FkziT6VHBmkX5So2MOOuJV4TCGVhwciu
4moDU5s5gw1jdaYnM/+28dVsLEdp8l3WcHh6eMca+U7hwfs4yyn9jyCbL0O+FzeU2OZQJZDod4P2
I+44mkmr9uVZCORCN+PkYgBv11wMMpbzwatQBSxqHBQ28QGhnyf7+IKQ+ZQsjdPjN6csbiFaGNIk
58ZDlNTx54G4dGpczAJmYWDnrrhbjH46OZBG0QBmMoLzfq30iJryq+MrJ55YxFxLuk4TJ9optGmj
l2sWbqCFWcO4dJq8TT8wIOLotjM/F781Y6q5uMpBk2xnuRkFwvHpvT/GsT9GI+T/2xwD/PpFfIEn
kSjLsd3vWpIAkid0Ay2gaQooWoXvTlcxhuzjHHKpp+jsqfe/h/KKlKRkrm+eWN0QHUvsFuf3DFOD
1JAKjz/Rb3zOpIrBr3WkD8hScbWblOYS2ttBKeOLQrk4LfcYscv3BapucQABjv+jDAVoMJmtd4qQ
tXhip4rjlKTu/dmMAZTfy5Srfvw32ZL9EfuTPoJSIDeux/RCHEplzrU61BoVGCWPmPp+LEKpMSj5
7AIRo1BnwHCBertgl54KCdrogcVKCmuftEwCNOG/BIcP8kvmxbMiL14EeTwIpNClq+7gSx6NmPcR
kaQa+uaBX+0kSPCHDzssa53jUjYKWT+Xdh3WHPtOA7DABRPpjai0CoZfPTXc4ZvBgP9Hur+F+PvB
O/D6ACsNi9Nz91YXXF8STu93K8jzAvgl5iqWpDDQjpfE4dCj9oQ3YupblnsajA3vrRhqTowCHmwP
d/4WGqQjAmKcO+G5PoeAupxg9CR+UnPKP1cbjQzX+MTYlwBCdZWT9r2K7PXjIy8v/6ObVOAHQrAO
FOPBtX74IzkGwARB5QlALHdzxA6LpinCzpJQrSzp9yAVBZKfV2jIsfCSMopeSXQmwJRikSc6ijtk
zMWFwEhWXtj8Ef+GR7jdJYGcKt8LJldVDoEEnahUAwGAlQM76lnpfk8jxGkCYn7Ucq7wXTThnvdV
eAZPpXpHMstJ+3+1A5mKI/lzkjNQedh5j2bokcG3h5/HFWCNJBuwANSktFTGa4loFqWmyFkX/Yz/
Xy+cAANwh2ynWOViJQ+brLI4Bamu1IbVL9Rb4wglZRkdqYhXedUdciqE4RoxWQDYF3HjrM3zF6HU
8wVsO9KKKLskO2Qvh2TVUdc4+yhW/6iMGD3RKgJtXA70aKC+9vWhL2iHjam7ieqWOh+37To8rrt0
h5+Nmb5uRjgUh+dRlmW8jtowjVHjJcZxLPMnnvJEvU5NKwqz43/i/ntrkrbqQMUI0NF67wBdPL7r
ZtlEhTOL9PoeBHxIYyZTc4phUeDstjVQFFidNdUJbGoWJN7nLQ946nGwjb5bIChx3vYAu1VhfYFv
VuRd/C8M2nz3eXfD/AwRmcjHeaWH1tGvAfxJS/8GmjTgImkv34d8aUrwOJI8whpcwb5pjm6oeo0W
P6oMy0SfwJy9hdDlzWKuXcjgVd5PYXdZ4JHNz40kqrcRz31+n33z0O7pYsU2WmCFBHntKEYf5ogF
ud8RgX+b7Wr/j7JsqAiSRVxuX7+0wF14676ocTwzBfR3ZY8SbtfWyARtw9+FMykS4mWvs19taBCw
6RfXUq6MvlQeB5dABK7SjAkMTu/TwM5qXDNjParEyZjgywR/NRB3Tx2R7d3MJigklTmROzKY/HDG
MtR4WfIwEk3mMHQyNXtyhzgoSqUE/Xp6VJLLHOVW3a+I4ADvIfUHAHCzfZFLHhp555bBGv+WiTGz
T03GEehLyC7mVuH4b5EXaCLTCum2PuCfW2NX2B0OKCXMRfECXrkuIvwOwBDotvVRFVfZDMS+KXTV
BUgSktZ7uSm7u9bpcWkcDW8PzYpn0z2RZvuK8Pp6NKCFRLptd5PuiQrpXZRpICDbfQ5MSFAT78+y
AKTAw4tgsab2zEMS+3FCHmGWjjMj/3Jver72RnOszSjvsBsItmY33gjUvjVtvKA45QOD8RizFdOw
p2HoRkRF/9FZn6HVBrYfIfJyazte49+O1jP1TnMdzHAAJ6vOveqV2tTnjX2lyZUnrlw51STuV2W8
W1+9GiHLphlFG4onELfGEah4SiC4RExO6sVVQuz5VyKGvUaR5cAFjCJaAC9B3kpOTVBGKGaZUSua
7L+4AHwZiC8oltY6cb7YyzlaZzDNOTBH+Q/CoHReNltbOAW7sRVQUt7mnDrD1TK26pibmu5waD3S
uW35jojFJMYazQrJsWyWSVR0Z48bX1JiA/WuATyuFs/cvZPlGkUfp/9JGMAjb8DhdkvbX89SDZzF
fzSNnZxn6CRhc1fbih3mP6OXioQHMFaB0I9s5T5vsdxsn0tjk71tgy+VQMFmXpkmi4KCNlY3759S
fqDzyjnuLm7EejtvYSY8heT58y5rt9gRDNeRSDHoEpwl54711d0V4sjmFBQe5tnQFebyez89XQHQ
Ts0QMeuh5KyJo6ApIVsRNxFXVeh4zU9FwWLHErZZUkRy7i4iUcPvn0jOPKuhysYWltdx7y7gCVqW
3DnZeWNDc5KHeGO74t9AqrUFLURemNnYnG2+BDX3OOHZHHfERGVnZqATTM+oHy8T/0gZ5HUQlTjE
eqpHZYlV3I2SvtWN9UqPm2OTMPenRF9pOKfj0sMc7kSk9eG8FERwg6Ow5NFSWr9QAzA2QXQP3315
lEhHqKl2SgdqR0SNsJput8xE98Fv/obIQeasLouCjepa1LLKtOejjwa8Ec3bQqAPrq2EEjW2qNGO
1nrAXx+uQ34bMsACzFzEWNyWUm3pfahdjr9A7m8WQZYGHMzQb1nTrQsiUzKugL+WL95VUTr8nFU4
RkPzPagDVGBG196isywTlNE+shUwHp9V+bpqZKVMLMAQ1c2FAtsrbjAC/rTi+fIDlqfQ3eTFArLG
XYxrERqHPF4CSFkaFYFbK4i+EzAgN66DDF4QkqQNsJLLZrvJwROgiMK3oObBdl4x8r0/D9ZJEPy0
3g2DfABD2cQ5typiGLlQ5nvOceyHrkKmaRmVVdgWWkDMEFkphwXBkLIrQrL+HrsUSv6G42TFNaK/
0hNsQf/nPHUohiHdb++uCQes00+n6JhTB1nuEfmDxsmEAO1xZbZQnS+8X897rWIgqEy1Xcyx3sB8
WQXXbLIPzhwhl7Z8fvAh9KwTP+wli7ZTPwMhTud9/2f9LcxDGNoZ3pEmrLcoWVVY8nOkC1oTpmKU
NbCTXvXqNlSVKRNVbzmQUfP/ZlkImxIrp0G3LaAQwPul/1OnNDptYpCxkKBFSHjC9f65RLU2xHRX
PiUYfE3x1eQ1fMlnAojfqgOxLw6LtVew0EkMaWTX1BzJTNDjlJ5/XnWaY7VQOBZNjh7RfciKgb57
JiB9J1IbgnrxW4rUfasdYnP9Pe1wxHTstEIjPRF9TZaz3NRkHAnT7J11CBfKEfj1C4YvXdn67Te5
qvNM5tJdRRYNOCWRSZov2qSEhoRku1wcL5dTO+yiLdP+NEZyxnZnOmSagiHAUAW37+0whSIUavTC
LPvgEg9JA9i333VxyeFAMATe2yoj4iLtKFpQEgP/gK15s260zZ5tD4IlCKywscri2zXdem4Rqrmz
2d1NYxHHSuyKMUqQaoQRWBeHWn3Yoa44xvJyjLUWMg6W8Xo3OLyLi13EPco0Qu/2tJysDuhEKsGc
oDiuIdog8O3U9UeNcryu4H6ujjeloEjAC2PyQKxAdoJGO7RnN3QoW9QY4LFOnbI6lRXxziJvB4YZ
8ZgGlnv4/5i5tAwBaatG3gHrxdZ+N16D614PqCjQfu93X2QTsPIqozKVtqDKZpRJOfrHJjSJrNnm
58DymceS56Nt5eKEeDAX1Xs/bg8hII4pbQCdduO8wLIXg9aQN/J5acAl+YbPkoVclKf9uy7drwvu
nSWaLmqlt6r45F7Z+z9kzhbsFBTGWXBTU4U+rLI10G0HuPGDhQdVM9bCgeBFyLzuXIivIRHpbL94
xwHfp1G7NA4HPf9d4qKJrSMuejFu5VGyi5cJ2PnejwMyXyhBd+eotcLqlMhIeK5Eca7jG7RAPPel
iWA9wcgq6NsoDQW3lWQppAsYVCOKr0ZZMM+j8KVP8/JESSztCjIzBkAwyuc9vEeCiC5LyI8GINdw
m8PPUIPFRIBrG672a6qUWUcV9/BUys/UjZ0xQ2rXvgimlN7Vew+4j9Id7HUV32XSqWew8rFhtYXl
Vg0MUn+Bw/Ih/bjEOhG1ipl080NS5MvJWP/Xn2xylREi+a1iG+t3MDEhNXtyPRlZta7GXUp1olvi
2ovELrTjoZVO0J3pcqVOduAb6obhA6l9ClY3di456fDcZHUyA96PLPx25uzM1Au6XntbAwxCH7SI
X2JQaLlL54JX3KUc2ro6ml4BL9YgVp3EvsPtDUnYbbm++6tT7ahGXu6DDN9ZFc62wIKaH46AFBvv
6ADMg6kEeIJYUwpCL9+3ZuOMwNhJlEe63siYjqTroZw4IloE9vAR4r37+8XWkgfGHy+79EJ6BLdK
EVmNXfaq/0/v1ZTTEvDBX+xfLs0s8prOt52R4phqiuyyTWaBV7thytTp49oLfTHqptFPLEJZE014
z0mS6t9Ol0FhpGcqmbJ1SvHidu+LIUzAIFqHyrE6my5NjqEAPgKbEpLaBJvbseHaMb7IKZICPjtU
xWoasM1a06lwN8a0jVHEclkaGCVMbuB6Khq+CvgILv6q6JMd+IlNVTKZ+0IJBa4kjBdXKnxa8h5/
rLEmWegWvmLPyoiOd8dOPbW4qgD5BuvaOrHyxWmKrMFPsjegjNlp3K1RhrQVf0QWAVtRCE2pnQgI
Q/BgYLrCO8Ryf712rqw+yjcnDL1I0Ckj8ytLcBhPnCxWlQDsvaRxQvPrSr16vs7Yv0WtdkMzTOdR
QQdvBJwG9o+F8Jn/rh5VL3PnY612JwR4I+CYSikU+5Xwrc3ibmE2T67+Tp9JgxvxnMLCEZDGHoAi
F/dJNcyVBAvYSk/Nsk073VK/N4tthOe9Tb310wkG8qiEQEFuP7KWviv4zYQOdB/XR0dD6gwu0yuf
pDAQlv5Huxnb+I/K4JzuvXashHCBEAcQ16D74r6P4uIs7tOfeaEM6Do/TNCQcIeZy7+anJM7TAbU
dpHsuFoPyIfrpd+7mRiixc/WeBESr0pgXeGx8PmO49Htk30W40a3jvuHBSNwCiIuTuSHzaBYaMX9
gILJzwL2av5TvLsYUc2gjlUInPlOC7w4LG21Brwk5g5eeSmp7o1hP3/x9Wrb68qGu4vrq5jid4W3
9qjvDSP+kAU9YZ0kYPRfR0Qxvt4GtACg2qDTQGXXVmwqzrAB+yvaD4YYBP/edIuXkM6Vindo7No0
0nD/iIoPD7vlssaKfy4xG/ji2AwxdtPJPCofMXsuuoqXaZcoo6yjDsW0nIWrN7Fy2BFaj3uzFBeJ
etRnRmpECIsnRjoOkh0Md8ch9BRh17JhUAUXp5mQNEAJtQsMMmff2BvqSi/HoYauDo2xoLVuIhBF
XxIdB2wuY6L1EOZGhLAupx+dW8p+mWN6XnGwj7NfuZsbfyy/pNt+OAJuquBdu6F/ydPACEGekALN
RmKlw7B7cqsNrlXKftTKKlQ3WNnIn3vRIfzp0X3U58io0U7Prm8kQU8Lq+LnmspJnG6OnuTWnjIr
xiDpV+Fq+SJsQdiifJoLd+cOWQQhlSYMhL8YtRoIoZ7ywcAimFx2NVdOnyYhov77EVTnR9py1imS
0pJSoRBa06RPDpxadvXWlXPxD5UiEUBmrYSeK8I5NJmZH7cTg35q6iXSawRltuBGYdh5lp+33r4E
j2CN4ywPKjCrEyy8sqoGW+qlYF1I75ewJ1k/drSxNMm4lXa6eihw2+aR6HKbsuIpThnhTiQabkq+
V0B9LnIovOluQLhIrQUkCbijLp8I1xDMWNJO2wLMjKCYVuZ/aqtZ1cRyn4Ecpz19BJKHltbGY5lB
2igVI4vK5DdwxUDfR8xv9Anmbfzj8sGz6WG3qGKhy2g5R+McYdUxeuRBvIbHquG+eEnd8jp3fKHO
ylSz9SbCp7hYiSOKm9nLjFp66oTLZ/EdXKXlS+DhCYYBBD7Y8LTsUVbJXvYc3+EqjrF3AXrmGQFm
Ng8/vqXclNAgGu3IGwouJ3K2+6/W/IztGZcpr9GMe6erjkCBNDEYDAfEB6iq88JNkEx+NbrHggT7
9ENaStyAr+V+5dkRdAPHBKOauMudN0sPr+I/2oIbS7edXP+E2883PEq4jIz/+BQVRa0ZtzeUWwSM
mp8Ue3pbxZGd9aWWGtKhDT5UbxNW0OTrLlejGe0wN2rSWB842hIcemo2AzCoTnjBtw17j1ZddvnX
Ukez7suNbYhcHL22Z07+GaI5Yn9paA9+HTh7+GrLWw5Fg5cVBxMHSqM3B7QwYASp0BuxMt0gBh8+
C4anjN48dIHurwUC0lXOPgRTZCLDvWLk7Dy+5tMHOrQN0lC72LemsUbt26fNC8ZaN2/VASOPq5Y4
6SMPyHetWf5BXN1dJQXEntX7NvdK+nCJF2935mRZ4Qu4rqXPxxgQMNpIzv8mVOX9bcGT2Om2nSuO
g6QHBEWsaL5cwevL9m9ScDUsQ+JbCe8LG4H5uGADn5+Z5zk8KBbOM85cMEK91nXF8h5Fx2gnzvM/
r/O2srLWacqQsHYZ/MppY5JMUZ2tkpAtZw3KvdO/s1wIWezBpMshLkzj0b0xalMJ3IkPT19rgXEJ
fSprKs9pqFsp30Ix/8KKKif7TqFzA2zNJK7GwOPfb1cgvl/uUDmJAatrq9Ldlux3CQ3Qhfihb0rn
OkwUsyWnqSZoSWkxXIOdOhYCAfEGsBgyAP8E1YkBgw3NcsyajQWAomD/DhnmwsG4qjfpnbZuAAyS
qe2tdQzg/O7A+qV5zScgMwCc6+lNbk9+hrMPxgMvn8QUo2OV4la//6hFhi0bKtKSj+tonEyZXLWV
8YYQdopbo9afkS8p5gXIvdZFijxIoSqi3gpV2lgA7w6LDRplDHbefEnKshARa2NL51t9tZv5k5Tg
IlXc5m8TY3gZXDZ7HdeJTuTTMhSjy7QuLnzbkebfdh0avixbdMzUZ3ZHsWpkvSjv58wtELedj7j9
iVkgRJlHBG1X3s5aZe9cNOuvjpr2i01G+IFo9kL4M4xDL9FmYRb+ZnL3+v5YhNT8gYcLduLbtIRo
fluCi9O4AshmmvC406MZ7vlvTz/01Inr986gt8CebBQypkrk90nmAyDiO9v9tftR33zGIMnVHnsz
jCiWxrdbSn5cTnafhJ1b1h2Th6Brnl3FEH+lXB0FebJqK9vZt8eojwu0uxkEKcsl7U3jMdgMWEsd
/ZqD9HH+9ndun75ArZtPIgBWJK7S71kvTetg/eBEWFbALjdjyoUjlswE6XxaVsB4nryV6DdsEd8q
Z9cDloOVfawAELg+Wjfu/plKyyYcE8wPhRHT9EShdx+eCmuDA8Fkxjc3pXUHuBndqMh8hb9t8epk
8QhoD1oYCoeSsa+vg7rp/sZdRhFCHPIMhoJJ/qvr638bGTNId5liM4ZKQNu9fCfZHBLfQAjI8caO
SZnkAoZPiQivzkIQi0dqmqGIAJ1mj483wcdWQQMdUOqDZCEDKFIP+unrpKpcztP28cD6E2GD0JhZ
p8F5AbLSgHPLJn18blDsDDc6l45HZe/JETabZxQQD5SYieOkCy8Z20jxTmZ1Zh0xjopL4SrNgzG9
e6/YYpitKHl361fnk9o3xoQxuLiqmmHZyvhhRpsL64SdEGwP+ge8kJj+wF7PM2+DmCyU6QA0u+Uh
XkyvGo2p9ruu8p8oFHmjY+yQOsm439h5HKLFacxu6o86l4prtT+I215e97jls7fjNVbqSn01upSy
Umw75Qs5UMcgN008GMvAepWynrEVsPUdHxX3RBn5xfjwki4d1KqPin+bItWP5Vqm5wgEM1Z74E01
jkLXnzFBwt69MGQNx1w5EnKgCiC+xW/IM9rbAJz97SMrPjA4GXY//ulkg2vaBpBwJfECwcphcVpx
0cMFg1ynuMon3puqKwEhQ5Z1EYnVsY++0qeQQRcN7M+Jz8ad5VweV85bg3/N3WtpRY/Tk1m67fu0
pQNQHOz3LK+uPieXkGXd46qvGMSA282BlknaXWJlC1Hl1RXkG8DZHrshU19REO79HvDg4iDTdsWJ
zpUlf2bjD3x43Hvm8M+Ad5PenfRPkYc8ywecBLZLfy9G318VsUKK/SldwGAvt0JwVqsPxjRnuKvW
G3Yd1pp8tG+St9IVTJbOx8Jl/dhGhGqnTjzp7IKWlVeiX0B9014VXX1dWPZlgwu3Ar66YkdoMCa7
6/m2+cgOSP72ymbTqHHi0oHdSjaYvFBxDv+ivWuH7V4lKDKYHEcfLe9xTlWKqFZRTdfx5nLGWjhW
OAhthOwxAOsqMlEo0xu9BJg0E/vpLmfeGJRhYYK+Jc96YAZCdmrpzxMpSAmoqLZkZRbHLqIJGp/E
85buUp4xLsjUi5IvdrFifiej3+lyZF0e/Emft7trPE5+4g3/zk/16Akjf1T5kxtuoZSn2Ah3bnsU
gfbVawwg8xx6JPUS+NORBOmei+ZBV7PO96MGW1ij5ND/g/KfYnwS9sWHGxiyRTTiMSi3sNr8NTk5
h7lBprKUv8tIQ+tiQL1bi86/reUyiMK6zB70gJLb1AXaHoH0aDFjyYqg4W2imeS+XDBw6zPvtysR
7Be548c8NbtgUjWRM5vVlYSCe9bSk6BSkPBowqAm+G043i8N3gCOmmhwBU94dnwcZTMDuNOYotSY
wo7IoZmXG6PzlulhcgOOJbHyt/x7NRj/GTkSFvO1Ff8f5bWdN5tv+Z6bQi/ntP8/JY0TFngNjRi6
NBJ5BIK+RqW/o4dyjDEhghOJetM/f6om+GM91avMj1YgLQ6/goAzbiXydoOtIak8h3mcFO7GNOSJ
1wxgnkdzeeiO8EdObsWzwOO7rGtUCu3Dh4cQEDVPyPRAnOgV2QDaNl02v4MKyPXDytcvLSr7roDa
UDpMbnY6SBjuMLfp3YjQWAHPjqb7nvi1ND/fkzabwZ05VcBIhx60wePOEFeSzRKugtfhKzEsmGCX
8sy5SdxdGEmI7N4abYzfPnyBAS6tYKDwNvcZKnUusH8OWfkS2GjbonT9Enr6l7YAP5eFxDi9ttDM
j+g9U+bUQwkp13dAwvgZPu9SPLgTOVKn+DgETAGTcFMcEH1OF3wdghUsMhGk2aWgE8IN7M4HLx7r
nONefwdlGTp8xZx4Vg/QLHRV2EwWssrYMgG2o3b88dfNVAS/ZiupHeKziTf94vRuWi78YOCWmB+/
LK2WWKtgzxEG4bEe7QsMNXZgy5ykRDUox7oekUIh/gR9zcA4na8hv/vveIe4vHk5GPYIKY3+Hbko
HXpbQ282hUgKLNdCJ64q3aNAPimvw8z1CtoY7cTiVCFkFrP6OnetNADjWJKp0ZfKQkLx/0pQ/dSu
L8ZN+I3kzZbzljJ+tnWF/NOqZCPmzosCxhGiEPZKtAt+RoNPAsOSoAfsppUWmgrwKoXtpYq56SLL
1D8sTTsL8dY2YrNhj8MDwADHXIis+pR1qiDvSqXhPnRoPZjErsxudWAhPYAqMQ7F8teRcb4btJo+
888enGR/gBd7gAKxdH8gftq1xthEovy7t6ihbyVprhvCUhKXX3X/JHnBquceFOqVe5oO8+3GYT6t
Cs6PLRGIVVKR04Jwk3qJQn0HqedpQrteqd/jDOM78sIdILpwUruxISIZ2ck8OzhbZ2F0FOzcGqkv
Jnx5tl/mq8NntbvjZeV6Q8klx0O1LLnzdEbN8FcU3ajNCzDIG9vwt+hyheXINoRl0FunSa71x6nR
AzVRvnhB4LkxaNOOHVUqUdrv+XA6iTTDDs3l4gWdUOygjcpY++OXdSjwBjCVBhOsAkA8T1+wWdji
YT5sZIw8EmRBcUqUUCEKCe+X5ioy1ptrTl7gp7rnPHw5pQu6LccF1SJOZ8ax276uXUAs2SpRZIgs
hDacn4Jz0cfPj50+xM9saWDG/bN/P7zxK3fNbu7ZuM0nn7CmXNA0eVgzUPry7wQXQ512lDaLAv7i
QysLoV3AYu7bJ2wq02yr9BgCEtv9uCZFIjC/6oL+3PAYCknlFQfoFo56mFUqYEIPSZPAuXdhrMxD
VBDT2cOnnlc6yfPlBnRQSReSa8zOwOzD8KOz9WgDWXPWqI2tW/jw7EK2iTV8Y5DleDhBN/FEM0ph
GqLNhsKX2Ae51ML1RmAt0Y832ANLxPkQ/vAwtuRz3YtfmF5X8SBPlmyfgj40BMSR24QqdOhPEIgB
hFZJEhA3ADArIw/erImA1xnfjhBNw0h44dit47/SWyIg7w+4R7Xl0uUBqVNlj31eRFn+GFjPzO5i
htYsGoWw9gFOJIU5iBku1iqQe0I4aOMeP0Z0jWJx2h9Quj+m6o4tIN9Pg420zdng9b+lrnktqEJV
++5IJhgDguvVUjXf8UTP2oZDw19zQdXPo0iMLMmMEOQITVPhb4XKm/6TOZVNPlIUiq7oRVdRw9iR
UyJIMJs8sIIDy57oREEN8bZgq/0PVwjwPa56dNTsltMalbEK34yfSui00LJYvwuME1xmBVGEenhG
CG8bZ0TB+IjGYOg79e8osgJ47BUotgQr/9cTQFZ5xlDYhD8tiuJ9d1maiSxUofkzCOd9E4EpY3BT
lGK4r7PcyD4gE91hy6NY/8HTRbUyDk+o23f/Fgsab/RAcAhVbh5bOV/gPFafBoKE02SAkqX1VGeV
C37q9HSRtHBhEGKybwWuMLMbub8OEDhlhBU4H1Ec9fvfdiKLUZicr80Hn09fsQe5XeOqzB+iLOny
x6vXtpYGA8FaEZACivi+TiAXKWMgJiF9rbI2i1djYiLHNL3pBeNi7ih9EaVfJFH4x16V3sPlKEqm
7MmGTOTaTTh48gNR4FUXP7TMUTGzdwgwn4TIGEZo+v0ThyvQGqCMqperaL/GT8sZsYzPrC0CFChZ
nheD+ysz5OFiQN4swn5QSJ9xIMn3xRt96A4LVltjme+cLxpnT2g2Jx3r2BPTrXIQy5PdU2kSiF3Q
z6ICv6+Rzdb8LYyykvWQla/OsSz1KAD/Kl7ERQbG5ZJcRl+uNtvQvHDUs0FKNZ+ECrin27tvTfTx
jR3QanjAI/9MoA6KRW0n+vK1YwGa0+DjJh01SL3rF1QhG9QUZkXV3XuVHFcvaJTHSii5EylToU9S
mfnBgerL8cxV9O6A1okSttzpF98DC/g5BN7zAUqHSNsABZmBBly5jgr74J4U4jukipU/z1ps1CHJ
yM4pq7bMG2ZcC7+8Cz2SUfjAMyMdZXBZWd2Et4/VUOPZmU6ldcjX/y57s1fCcqKhb+6jjWCEegxY
v/X2i8I6bAM82HXBevSR7XBat/4orSgvR5p0S7aWIJ08Zgzim93NUvY/M26qiPUt9nLJugntRhiP
syAzGtXzIn/RaLrHwKbA/m9HOMLacoTuPaUZnZjR9iABOpCVn1cfrJ4eH9ctxeRDhYY7jkot3Lku
9TQYB0bKRjLIQmhDR9kAKsp5s3pvwZKARfWcT0I0khwW9wCbNapoLL5w1T5Sdob5yGPkvrGu4kbP
4wehlOEQpIFkUbzL31BWcqfj2dwFu3yPQjUC3ylUD+ot572A2Gw7BN8Sf3dLL+bPkNNJ8VNA7/nl
yFsi01SvjmyZWlMSmgxnsi+WVmVvIFkiin7yO0Nkr7lgv32LCUGoIkcT4f5VlMtP6N22ph+mbSiZ
drasOPnMtueyNgNl7utDjB4b4OC2dkKdidRvDznEBYW1ElXQ7nLaabScqkLH1hfzHaT4antY+U5C
yqziDVgOzG1Mkw3ZBHEtWehj/38PG7o7om9XU+3B29A70oJL1TduqedMXSdEmnlBEyf/bG/mak4b
hM39a6Pha/ZRCa6pcVx03e5eHKoc8UCiMZsT9B7yGJYhvBJuLGHB3JTTkG0PUGBSF/++s60xnBBq
uYKO/KVwlwLSwUVSYn4PrOvvtes1XrzRFb4abN8RfZhgD2BFQnRYMApHOq0Yt8ei5SYpuWHcDCjD
UzBOmegr9+j/Whv7666AVOowhax1vp/9y7om+RUQ/I3obsyYBCpy2jvVhmzQwrzl2VYM54ybbwDd
OqYFj7cCW5U3BA4EcgzUbw8gmyCoEU6srfptFN9C0NrYsu0eaJF89DEO8zzcgwC8ykTriBWHJs+T
aruxxESIU2y2rX8MdL7TV6MjaDDEZ4N/CPIO5P8emme0UMM2QaEF18xLrIHr4c7UWnN2ZKa1xDh9
7DW4QYpJllJTGIgKZliaGKQ/4nFtsE2PSIU9ZzsUtL4ukmta1XhvhhSYpvWiH+JETDFYKny4M8eY
NGvgn8T2NmJ/4XV4iIKxN54fRvACFT2CzBIaqeUMNAND2oHeUdgvJGfcMwt7MQ6FPrjnyBckFdn6
/SA7QGAgV9mPvLVznMKANiyBX6I7ktqdlxvHijHkNYkwA4/qgPUTvueQmosUJTv6kGCnFcO3OE99
X/6BhoblFdUMPvvS9tidcPUNsEWB36p/kS1KtyQbxtqY3yDI8NLmJRd3XwY5in2lwDbvNct4tZxd
/IBa/UevWku7cPcmxkOachgFtcHyQTo5MUZrVXIwarxKnjHUknveArGannFcL/VEg4GwHo2VaKs3
pJy70PdyjOdHZl1VVRr1RhCF+kFSJSDfxtu0C5R1jKt51zBI71GGiY18rzKQFFrpHAMf9A0BRqBC
uzQszyf+VKxQIiHvxvPexC91ldNif7+aqbwdhDkedoR+ss4ct8JTQ8Smiytcph4F3RbOTSzQJb1Y
w6kgEkT3Ue8DMiEuwMG3uoLDU7oSCxfHa+oCOukvkk5mf4PR65Nl1Ch0iC9gLrFHUEtu1fsglASF
a4ZDGN5SsgdDPmMnCHNz/rGW+4C7z2yxLg5W6g5LVGwIcqjshdAGb/2yCNom7dpWOuEaN6LwGlT5
f5tfBs3RWOvKGw9EiULxJwl+gONePXGRVubga00hdtKKtZS9E/juWLM/f37lGnDt9slX3T0py29l
Pfqd9uj7dRWdH2AZqDP9W8wfgfKpnH39zIe2wf2yXJkaCWSEnWX5elegdKARxZSOpKgJp8goaq7m
MSoylrzF/ovc3QOtEtH+8P/+T3D3w38iI9o7I5YL7nnIpesXoadlLSDV4MP2y1yY+T0Ro4bw31kV
2qi2YmGfdNbY/qIVT69WnEAwPMjZ8PaICaPoujxAKKYO/9uK85FHraQPat+znzt5bCY8lr9DRsdi
g46oNU6hZRRvIG+U7JYrT4L143QlaWNNidVzC54CsXCdso8k1Y1T4dprzvNBDlBkYg1GsL7eB4q6
V7jdCemWwTMrZTJEBOwfqQ9xxVfuTewK9e5w7mwxNUO8cdlaPPt01WeG2S9B1wufBmT60LINmEoQ
mZlZcUdo7ppYw5ec8TnZ3CCOo43BavSIjI2kDya68oc55RnTDElwzNat3AdKB6BOm/JZMptWjI3d
8KdaX6Izjr6nP6ui7raMpHgl9FFw8M2WURPm00w2b5AuQXVfTqIZ7I+DivKYRh48HBrTi9kvpz5L
L+YlHqwG3mb7y5nkghh6oPKxSTLe8snVP0PmmqBgtYnKiEtSW5vBIpTc6mtU9rk0k4F3aRWiJ25C
vMcLao/2XMVagCcE57B/4gxPlrILGPVfIN+rwIDNeHJoCi4ymHV30z4JCQH4kdYa3Q1Owuv5Qk/B
a0K17DlIdiQtwNA8abg7C/kV64EI8lB+/G0qkPevdpUjYMZHbvQuM8go3GATzJTpY3itb1MvqJ6n
JUUBBj+R1CsSwjnZAhtm4/3ZBNE3K8IxwjGlc48uD3YAlz6zxpYrXzVjCS5Nr7M1QQSDpGXf59Xm
Rbw78nH0VTSwtdU4Lur5a5R1TmGCQCbmTL3UBdn34CUd0hnc7X/+vNsO7VJYroSx3FcT+zcEZkiX
AaJ8AzkGleZUKsW3Fkv+mF0CpzxX9ai7D5fa/NM/+T5BEBX+sfoPL3FvC0q/azQeTjY5RrznS6Bb
XSNiwYCRE1auL5LIAbVt8EHUvR4jtb0UP/H5Er8tu8wAZAkJ4eWdZYIVjQ1+1HMLvW53K77IaMnI
uZCQ3H5JTNEEuKTQT3kOIn/Pe+dzbTvl91/+ALsIC1AOeBmQtTvSMwvaX+zwk0th1CRZ+A08H/hC
kzlK2bcwtYETahQVeur3LzYhD6+LhX5E4iybKztGkALey9n7kjtPeenQBoZeIce9QMCGUsxmR5lq
Q4L2Xsbq/quIDBEDuPqQMpu/Ugg0opAa1xM2RnKxwiGvNIUd/AIPUaUy0r/jnDWQE0F2WMYFuqXg
K3Vvd2AoRxsFs9YIL4AxJ97BgSkrErGRciKGQE4dQRs7ZkxvA/MfOHBhq7++1PHBdjryjTW5ZHLb
Dl0iPafRT6lV4OWcMqbD+dB1pTKgd1BGlh9iVqC1PwtSz/ZvEZeZZalW3uOSnoxytIUQm0M/bxwC
DPZ/zqdcTlGvE6vZoe2Py+gpwm36kPOBP7vs2UpMVcibHL3JAl1eSWGN9QgsB0NXCK4u7PDnDbDh
8qNz0dNefyVPXzyZmasyTz3QHUhJHOYjJX4qlpU9jGgO7/LmZuuPb4450fSLHlB9Fk3s/2boVKzu
13kiuoiJgxU9lds8hXs/kODPnbSRvpe7N9sYpOzP5tjtm6NP209m5rvCg3+IU2a1+1tadNbMW3cY
i2N+V3/h3AOw2kGJkBDonc66ObY+nXzww+U0u1Zjhdbw5una1KSHdzdnhkZtmkA7cPL8yaHW1fx9
LTbBzwreuUMbAI7bhjhhtEWffaKIZ2ZgFEPIZeIweHpNKUMSLX1ER7BsknfORpT0RS+UQWT6ZXpN
FAfEnujCLis2Ns8qbOXhO+79hP8QVakqXEtvVr0tDiMMwdxqbXBSmKUaqPNXDatB/oZolaQfv2y6
lWfVyE42ZJRfeiW7caAupDl27enTz12KellF7ADWwFv11ze4Ke1LjWwpN3/PN5IpOI32SOafKOvo
lun/FVpvwa4NjxHHVsxzbdgl528iIsmFQSR7w/0zAmIGqOLOZwUc1bo/RRzza1dESUd4Fl8geljj
4ppLgUVzfl8cXxh88DlejX0kZMDQwLaWbrf2v3c9wuAZ3aUbKQH2fTkeMrxYcqLp5lb8jcmZxsRz
7aXWjcFHfOX0F1ewj9lHamdnck+iG85JxxIjEt4AqNuW9t837/Gd4yrzgCcWUxTfIGj86DaLyKGO
VEhWyE17iiSZyrf/b2A6CNxrqxoHSX1GgZA0T4RbujRPSuZpWjqbeRPAirPB/n2gJqBMSY1jHxsq
fVC86ug8t9HVdUFwnyvhG2wwfCnLuFlR5gY3UyCSim8AG4xM3XhEHmcjvTZO8nRhFYNgshmnu63Q
kvu+Q6BL8YgZlvG9SjUQxVNdmJEqUKz5XQneO+09MccuOBHAlfyNh1FDvJiMHO5T/EZPW4dWX8KZ
jcUwUN+/tMXIS5tEaE2A9kylyRmMCiMYcHzaBzvP8v8M4lpxnDiOH1egTqOS2+mH7oL9GHF3AdQQ
oedQsPJd9HoUMTtJYXZg8GaV3II+PICVkn2oaPET7xPGjhGUWSJq2vvdEOqllMFikJuNn9w6oXZj
vhaxkstWUrWCNlIUEw2dJRxQdlne72GK2N/VwtiRNGzEkddlTD3nD9KCemcEJyejQQ2STRWZAuko
8eaRJzI0KznNTBDtDHACabWDMvcWTRZCSXquj8wJNnB8EZIQL9NcuOen1dhxI5tYyKfuJn62/lNs
5cwaIK11ROM5DWDVH2tkOSYdifusaZt3i/+lBsXVlalLuauvEEhBe1bG5s8PwgEvyEMDwSn2jZR9
LIz+2FWnBX/WxY2tZtE06MVdXtisv/HUM1bhxWyUQhNBpcmUww9mnQUYDiY38tWThLWS1BEvIf9b
UQDNCt25Qu3HDewEm31W0FPVfRFfZ2WHlT1u6h+c1uv3eyWoIrg7X5Cy1ELHJQWEz2UmsGohTbgP
gaQOW1xUmim8x8jMV1zZWC350DPLSZ4hUFs4wgflIhwYuNOn3oDjrEoqli7JrihIdTKefWRXUrB1
W9ND8KSl7pl6HYxOnGLY7MCda3LwQTmNfnMaBJujrNtzdGJ2wlIm5+Eu1HmbcQ1U7+odI2w/c9qG
+PMGrR0QZOi2fqjvy7kUjNsCFTw06U2CoZVNwKt8fSCuxS2FlVdkI7p+xOYIcuI4TYOyyZHfHeqp
r2SB4dVlhfTFGHbkM316arCRVyJohNqu4ijTzcCtMHHm2XRzczep6oZYsIrMuLu8soQmKSTNi+FR
Z7FnYg7c0ZUDvJMHlL3eQCWZ25OaTyztCj3CAcPxJsJqc1Ny0BcwOCJLep/xlQdPBn1hkwCgijnx
9hWqE0rc63TBzXsbL/lIZsJqItMrX7ObzpvzJEvOQgZT+pMbYMclQWEMHwNYY+lZBGFCF9TAPx6g
YXQcNcKiPCXTLbRTGEtuStCG0KqvyCzD6ydnBDFl9qgdoBv/3whFMgdKTTXOpu1L5eNmTcsKYwcC
1/vkh4D1bBPCvzIRbIs+diihcpBnAPR1ZQdckGYAsKE5nhjizBDUqlCj2umVH2WFgoQpDyD8Ei/c
u9rmZxQU89BbtzGPNLG1iEmh0sCIgMJ6Y89DmYvfLskKv7ELLNkX/FslPSve2khblmZN0dRWcbNY
asEnz0eHQ+3Q5s9n5a+nkna0orgu7gxES74a7MJaxAMMJvP0pTZjNBI3btnFORCZEjJ/Nb1cUoVu
5sqH32JfIwU7nItK3z+3G4E7tuIh8k/0kvUkxdxNVUSD/KtJkMFo41oi2w4p/U4PZ5GnjdoLea1c
HjeII6SF3nQtnCUpy8RXXOi2dtgfnZPDeKrnA531+KtmXL25vP5nkO4MfMrHZFDXVL2BoIy2FYJf
0npQB2OQ8ME+YI29962mREXw3O+QuuLsL0E5HSAwS+5PO7FOjWxcR7qPGdVC4d4eLCOP/ZFRGUnf
An4ILBJQ6aiDSGgeW8O3WysKJ52YuFNQBOGOgSmae7iqQxaiFCPuPJBs2p/gR1xNP3em5hrSP879
inIa+72Hw/7IsCb9BE9qDiIm5tMxsvnfyrqH3lHR+zP5opifeJnTe09stIV2DHorxPGZkCqat1S9
jcmiMcfng2IrUTdc4fSvjNFj5ZL9Ix1fEi0u12zgG+aBvZmMJRrpHFL+oW22yramZM/aiYboyFvO
Bh32H0ZhlH4pP1wap+YM7g83sK3NwRu73+xqpq0gDIi6wizdptcQK9620QcVxbhc6kxCr2PoBE2g
R0xoMGmmOJ85gfgnKVS0xHcA8z08OEDMME2StxUlsRx82xPlJfnczC2m2HxqE4dFh5snMJYXv7No
w0OEts3J7d6+ODCO37oMeAxTHjlsS/ajUjcjh6rvkWpPPVKqGPTxiL0AvxZJ6Q0tMKx6fVL7qpmn
D1Ah5fYBUUZtVhfcbOg3YPworYhWgG+8P1VYhsqZzGBmSIh0+x1/dSCbqSjeb7rwk5EWp22iJHF9
umu+Ei93CmYbFc3PBQO95/14qW1P0jC8b4XeCgDh6wKrb0Sxp7wNTxvaym2aVUpEcbnANXMLhjLN
NQm2xwdE/drf0PlidvcBcPOph+Qs4ulk2/5XoXlL+G8dXsAYo3/2eL7JWl2KZVgqXgRs2ULUd3z0
68BNNb59bxaNX0QgGWJlAUgjXOBwSYxs8kYWjzHwQktg0fUZ5hALJ9TX7uEQjg1yxeIvCLlP2dw6
sdT9VPLSHDhALQb5BI4e/qAa0veVptOC59rvbM+6VN+HR65OcVeGl6zJjKOBjVCOsN3tlvRaebK5
zFHU8p/N/mqEwqI2stQeJpSmB3mPNExcgjh4z2G7oZZVKfGFwJ5aJLjeip6sRy2EZ7Ocn/2uH8pi
zw4M/F4Bnx+zNIDNuV9pJ0M6NilkfWfWcCDGfvkinrL4947T0Zx0hA0bYGEGx4B6opsU6xSy7v6P
6VvgNnRuh5apfhd1POvMowplXHv78TBfry1yFt6VHh7cJG2LSibVwYDtOJqldSlfv/eP/abEQ1b+
EedsPEvMhvD0CWlFAGts/e4iPflTv/Rz5tlR4n39EtXwEGxPLYumwJn+UQXbRyOO7fF1sIAe6wA8
aZF6x05bCKE01VuJNj6Qk489VDahEFZYI8wYl8qr/69ZeWdP1X0EZzvOTg5ru40Ds4aaRpTE6A5S
Mf2sE0Tbtsn2MxX3S20bb430ocUfZ+wH7sZ89pM6z3t4ATpGr1kqaLqunEWpvYx78aLaNxh20Yxt
GwrWZ7xj0BJrKKpqDesjR0P8BPlXIqkQpdV/WmcSpmVOfdceuXp6yOo0/exjIkht/SxPKAZIhtuj
B3qsmr5ALFTO0FEba5LnZgUjyCF+PePOKbDfkKXwO3//2cv/0qPnlTxPpGiTQyC2b7ja4Ug3PnoG
0fpvEAe4k9lUUz3qH4QRWEE12K0YnT798yQ3lxDHofMYZ9LXTKKHrEhd4PLfQa4k94RJE0ScvKbr
j+8qqDg4XVSBF4o4Zrrcylmp2qSmDKCqL9d6sdiNBZtNzEFW9WVF2iplG8jelYgvVCOKbkAtGRIU
Htr4dYkjqqyoZNbus+QxI7B45GIO2QhfUKfn2qrNZXDlBlpBVkbXHUuoljuK1pt8hkp4eN35NvuX
fp91Auju5sNLpZpfBia1QRorUYtVhNC6s/hGFkC9Zz7UvCf6eOMS6FhhUo5COejxPjkBXkwI0Zp3
3NmukkmDctoBVl5xCNoyhQ82ym/QjTU0Amt1zcAIz5XrWP/TqqSZFCoPfOvyWk79G2229Z8AXdoO
OBHPM+sAt1/DyZfJHunq2ylERCBBKCrK5YbP7bXqyPc4pJ1svODmEriVSBRE6IyQJxrRc0J/BYso
N/kPpva70lcqdAXrc0aWqAyOnrNSVp+sSPcttKBEtHLp1/zMgRmy6LZBSzxO6Dkqftzg3PfVV1lX
PbKrV1rQ7mQZRxdNT2YXEsnkPXYAEFHWN85uLNmXyv/wRxbQS/x5CntruYmDaLU8SQcT3sL4mNb8
Y3HqqYcI7ItagCB4gMKIpsNwpvZnMOBPYx7gnFs83TYM4G7EIQ7DxKMURezNLNKS1LzyUjUlhlns
JIfUenGt6+c6YKw/B2G9nzhpVrm7Y2lC4hiD/BPm9RByd4DE95rUnDJYIJkQXp9TF1kDcPjGBJoA
euBYIlWsl9adrBxE/DoEclftHMLHm+3TCmtCnJWlmk9jlKgHjCm35NZP1mEZbhsewHWhNo8pr7Y+
VX2Qw7+41t1meDNMjAKfcTsbcU0uI88Bfz/GHZRI5ZiSTjlH+w8YOnKwRMpgUQ/xrbVirLaxlEy5
Q1ekEPeIp1kl8Xt+IuQZ1HZwy7QBet1Ojfs3b+lPALw4HTeTkMTwVd1/Lt0o/llCjThU3SSbGlsw
pyy0aIKhI3f1pP3HJg7HabZFsHcIpdYSpPkuyozMT7usNIn7jeC7LyZ6+RhWnoVRpzGWVMBf42HF
s1+kw6cHBeKDWgClyzDXB5pVBVBjHE1PDNdEPkRUqsi0xh6xeteaEf21SuhxUTt4Uq83jsplvdov
n5cj9rnjQ53pbXSD78/G8lOEqyf8Tid0fBVbBNIJEnQ7vfzUBeBf0dUIEo3diiBjAHSaI9uwBFsV
+ZxZJuJ02qLuOJqadDeqIk2sDBbr7xIkEc3Es1lXhxnYp5h/Esmz1b4HP4B98fQB7tgp2sxrB2PK
CTqGP+AiKujr0CZUmruLiNEA4h0HhAfY+Ie0pT3DWt87e9viFHVeysXXFtlqEYliNMWYitJ9nonb
1BMDthTUXPHHlzdd3sNJLqL+WlbuOPU3ESxviokgrmhmMLOCS7wG8EWrYKrAjmIbMDPqPywztCLq
PizkgCeG1isFVW8uXzjzbuKOSFpSoyj8hV3rjsyFRKnQN17uIQC4h3ZGrpuAgVQVd2RX3IUUVhrO
1pST7VRfelRnM4LjweTsOjsL6u1wph2L/im18QpL5KjQvJarOxhq+A9NfT13TF1clS99042gg6YX
xAI8WCOuyCDsWzpHU0WTOM76ats5hYz7vd/+NtDeihjfT+5acCCUVC9+7og4PGVvF50F6O8YICza
S2NQbx/B5A6aYhxkFQytJgmO9vJKWfHn0amosV2Axob2V7MkHyyS2dVjL8sNyd0tgt9UXtmWcSOA
dJM9KLEz44dMtd6dI6CeMPJ6kwwqupSDS+KevE/0+X6Xnt2Uz4XxAccCfZGnsl0PMTAMfZRZO33F
DcUb3teBqGWcu8P3rCboL/XltIAkkfyOtf48zQQaiE75Ewi4vV6jTN5HoUJOdQMdbnT6GIQ8sLge
HZoZkAmLZ0TTcdNxPuQKuuwrjhD9Dzr6q0Fj+grhO4CssxgTlj13//CRARuHTo49/zeEUc7VgBBf
VUagEbXQjs4sUZ0HpIjfN05xUNATGPXKiuvka2/KOIga6b0ynbN2LUyra1ljdoNsj5GCZgKwf+GI
q4kvVlyEWNxBpGrBpWaoTuc0lCmygap7o4m20TOzr5gnkexoz9ruCySPSSJmVnVIZW/8MUTSsBTJ
RScEQC//Ak1MaVA8HaTHRgQ7hcTg7/FRB2HDuuaD3FKxigZAsRMrK8porcOYS1mDP100fexNMvKg
5mmfS+/kuyBIt9p6kvgzoKrn6Z7s5RtK9wHCFbGZMFFRs/MDFnX07h3MyGTZgcQ/e2kiHEJ+i9xc
Y9kqvS2pYlAvcr6LnhG/Y5n4k8hLJlr/bohMe6Pudx3mhf3P/X3+zprf80BZ2CNx1crfypLGTdme
FLyVxbYIqtSBjVRmfyZTjpxFTpGK7BwnqY6w/TM8vT2qClc0T9ERV0VMqjUJEBj+Tq3ooxrTT/dg
rvkMpKhyplZMoCREldCOuXTbJjXOaYC6QPo9CodK+WZTUf2a0c+9dbKuk/jJdjbMo/llR33tZ22L
jhRbgMW820x2CwoKXOwAr4g0fg2+cCgwd0zVgUow2LAQPijqdz9Tu9gWKfyhTgqDLI+U9AlZrMVy
FYin/E8V8ky0gmTBMdj4lBONUZq70T9luz0XenvEkegCBr70LlwFVuZpvjX9CNnn2jm86STwiMIj
z3M2AQpufk9vHuGwQ9ohYhGXhXLbyjM4njub+rzNsxMfCe6fddoxxRcHrIsBttVRShjRWDwteD6l
9GOnf2KxL8dAS+oJTCMsi6Ps63ssnnDM9OlSqp1zbTGRxyxAPmPherfWx80VOQQ6KuIBjYYB5p7E
IPYUTkPVlnDh0EgbMaiJkAfdTvJzp6WbBofMRI4Axtv000xCHdm0Lc67kEp71HDWfZKBwk6LO9r0
qS5Ld2tW0DZkrItbUG1KLLTWWTsvnFrnHzbdgJJQrimt86uw7argl5Y9QBwnjheSA7dp6wzl17i9
Wuk41zVRfQsfxDeI056oA+QL+Dfm4YN5s8Cd3xe2KJT0TrQcHVZvxI002ewGXBoZzAsh8RWPxax2
F+MiatQoJwelwOiYxuxmlp2iJ6vVwGV+VJLo6DME11h48d9lEgshOzcYl/E5fFErKZSMmRHTeRpr
LTs3D/OmPSbs5B82d5GHBBcPUiPX88hPx74KlpuoDDbP7GAwvIjtl7lO1I9W/h5FgQUM03Ts+2YE
sVegOb62ItEtj4cDoIaGGaRQF4tTROmcPCQy6GQtB7cTG/8/1M23r4uhJ7W2fjA9QxGVYyw8wny2
HB2ADZcHpb/5kRyAFgE2mtSS4QzK/Mdt6FwhnwbRbdjcNRiQ2Sh+RuucIdPs/DGb9cdqFsb5CkIz
BJCIE4wPzqFlaD5niCkmVs+MmMRIWgXm7p1G/owwkcwePSUPZe+WP6sVGzewjIskx+I44GQAktdz
75kHfx4S2/Zx4ChxN1y8DIgVOvr3E7tfASwgD6BCBX3vBpRoF17UBvc25UVx6Kfab6l7FVv8FmJo
wiWE94lOTsG1ZyqGe76AsCUyb7c8XpqL/quVQ8JtAw3b9Bd0gWA/CRzdpzu3H6GqjztbKiEBGpL7
ciaVIS822FNre9k8cQAtZxXKZbV/VRXLMwIPBUazOxYiu6NKd0+OoJwvqOqdbjo7cgzaXFkUl57W
v9fciUa2+EvvsciKQllhOxJqYwf2VBzswxcMN0xzW5eMuoB/tc2iAKORXzz1DYAzN2x7zWihj960
YPKdcCM2hIrzwNw3HG6GFHBCN8eGNd0qufTgagV8driDwGU+l8HJe4aeKShhu6+OvHgXvVKR6JJR
OQfkdrQ3A14EET/q/yip7WbjWJC5Lxo77N3UlEzyOdVhOisdZeiZd8hJZzEjerCpFwcqDMp1dwAM
XKrKqB8hlRvr4/P15YvwmIuRYzkKzXhQjyRCW8Cq8OnW5DinEmZ2LnNc6dbxAowpff4nuBqe6CyM
W4ynpjs98YsjmAICYFVn/Zn6VJ7/2MMgtqdWzR8VSrj0PEcM8+R/mRsgYW7dmF8n3AEEbe4919ZM
IFBqOT2n/z/IoRi+VlplYEFPqeZwsv3F3/s/znPlqk7XKlnMMg7GqEIsSVfD6LtKOQ/FdiNNgsS0
lRYBOgq0y+KlgcfMfRN9vnOK+rUWPrdx7pxMU4tnJ18UQiWGoJQezy/V2cL4fNTvVMi034/mMZS1
EDk/zOh7GFed2ssvzOMGnfMfBUlDSN9zcmSbsRmc1vGMFfG8/qo44QFWBUUV/oKKSehbGSntiF7v
jQqmUZwQjLzEUT4+mgPzk8EndX3R4e0QgGE0yGchMGiQMfoPtiDD1z+E4SVLfq2NkrghyI1sxnFi
/sbh9FvrVPJPqygotB84cfKcS9tmf9qQL0GKM9hV4Z0E0De1eIfUyq/27C33yxsoj6unDbE/thWT
kqn7Q6nrU0g//gsHLFIfqoih83dCEYlxMaPqYvv/ktLKwyFqTVdzDHeiCsRVdww5TX52U8GNJnBp
bkV/1yaIAm9xz0vyEYXBKCI5ubpPBKTyEj/T51zHJxMlm+HA3SHdHUZPH+1Aj5sz5zi+drX/pfUd
sk2RpR9Ov1EydqfzkqT6q6GsTawuFQOb8czhJ7y62BPeNgHIphinfPqUOPUFulZcwzLWigRCv20O
oeZgLA2bm1HW/z3fV+KQS2HGhHVd7xOmXeHBZ0ILWN7zW+OoiRUu893T4fpuXxJvFRTf3clBpp9Z
+to+uvz5yalojgS67XlmYVsI1IuVOb7kGjYdH/ufnTPf0JaJ7R1KJxV2jwJPPAMYrAuu+QR32Q5x
E0wrW51fT8RJ0zkgdNKPWujHrjCuwxZpHoVqk6QrJvatTpA0TBBplIgqK46ULdgBWX+kEP0gZY5n
au5WdG0Xp/Ofqvu4+KOj/kQp0FofIcOH7j7tuQIc43shKvZgHl4UXDgp4ZqHjnVmyrVg3rZWJL/h
V1NCKtTqkLH5LOYK/ltAhzjhroBGJHPjdcQr8HpLse2ijw78zexSQaOp3wtVLLbyD/Ncr0Xinco/
Niz0ut0D2AqJQ1VJpRtJH0toKrnGaMdVeHMTdbOKrc/sQUuVkMu8T73m7jp91bn3WCxl6NFXR9ZF
waYD4KydwrDSPku1j76MqbX8zqsz7+JiVHVfe4z4WjwmnO8TJ0U0jI3Tuwq/w/HQNYWSqF3ys8c7
O7KBbobpIi2EdUOS7YFIREqZSOmhdlgytoRf43VDWcHdKPDppqLxLKLvdmCTiDhJ5yEohgRk6D2Z
Cq+v01nk2uSztmkGv7EIOexf1RO5r6SS3cSDFzX8XDxYeZeoVj9VJVIDY5Fvcj7HbBmQxPN6PUhe
XHFcEnhH+crEuEoxksi98lXwbhcXMvd3WtNnP4TzjcsmdqPoa7aw4FGNuYrArNa1uAUpiNp6uMeg
cQ+AKyCldzK2qoIT9V/a8DxJR93LFb8N/UHxKq7UYzkKuXzNo4TeQiv1EiprevPQzdRgQR9jjpDz
/2ss1iLIK8CuaWseTUtVkW1zYE/BseMH8b4f3V1Szx9rklYtKoarMcW4ZbLzVVkV2xRfxPshx59J
frvfgKCds/Z62yce30+mROMfbNxvlv4j68lBMCMQPyWaScQYqDYTjFi2WClelV1b+Knir99/z/Tx
SAhbpLdUkqiXFhRAEquntFEEcnlhtQYgQfwsL1EpwdgK0cRA9aGrNm0tOCVjBhpPNrehpdferbH7
+nOuwR0UDAmjc5xwpVxivnEsW9z/JxKv0I7vZvqBaydjZO0QeRqnaoYF7g1a7NTDo1FvIAZdPYQ+
/mzB5g+vx/RcK4jx6GxxkmkbVFv/jPmGnAkR2L61bVYhd3/HAnnqI29eZ6Je4+LIzBpli6M4UDph
00p+s42ozg4MBK5D6o0f7mw0VwPK4Yx0gNLiM7oj7bQ2DPI9JovaohJTYBr85BaUmG2ULSkGpNpD
y380Zb6tRkwxDN5HN/W9q6gMXD1ohSNzssDiT490RNxsEr62O5yh/9G1BtaJD0FV1huhagmD3LN8
4+rLclf9hnqzWRkwcsYkg0RMco2qYUBdu9TGQ/Yk3noBJX8YCzC1OJ6sS9oocdTusdHLvsertw56
ImOfOEM7CdSnCAl3cL458gZTCdT/I1lNAJo4kL4LobeAUx35oRO78rOQEn3sIJQlJajFMqgXggWw
LT0nh75dTw7cgmJ92ZFjCxgNudnTFiUJIYxwZZyZOvE+cOGxZyNVW4b53nc53imGUC33FlTVGex6
iZOPXwf3snzjm6XU2lJ95T5GjmafSbEqWufpe4nSm5F+bJ7kfcXNmbL5m5Nb+LXdOWTlVtLf9Jbd
sGTvm9xhGYo7Yo5v2/4WUKcoctRHLbInFIcbnb9zZdeInMOOcQyY9mlAMtAL2KFtE1gFwU/HywNU
TsKQSCeMBBQszNgukCfRLrddbZQ5Z5ec9+I4GeXlqrOhxwKq8rAVDAPTmInQgQ8hs1JzYWyER2Wp
sri1txgEU5EiT08rGxYVT9Gg+ofwT2OR7n1WfOHqQPY3fuSgWQ7nwLYQjw+ktMucCU/ApUPHE+o0
GSLeVmo9V+zDMKyHjED3I6IMOcXtMymT0bG97Hl5PWrWQPZPP4Fj+W6HfBbOWJrZbxWPjF2CM24/
kDkPGvB94jqUtrQdBr+v6mUjOaxY4Mmlq+ROJ8Do3ulrRzoZIYJou4p4687iCG4NzOSVH/86fLaW
c7iE2c1MH8eYbar2zcHEXMbV3CZxb1ZxAG1e41nny3UfEDxeLa8TRL8+xYKD2hKUgpK4WLoK2m6C
TsAw8r53Eav17/HnW0Q1mj8wpEzXxxHlQfM+YY5AS+3oPil0JfuFDfbIiLg/6sYdIyUTVyIyySZr
e4cOjt10DQp4extuKCsdR/TPScQarS4RaEekcn9V5yfB7euT9WpnRLeO7ENH+965wJCy8rdACiFq
Cwj6GaMJgwq4/aMXupBUafWMGNs6EzCy9vhvEQnsSieRofgsQ/HdU8iKhWPeMHTCmF+mJo04OSPE
aKFLwIn4fK2acobZL10K3Xx4/AhzZe1QscmKEk8t9u7H1Y9ROstxDMI4j0M9f0jD8kSKcA/cdYVF
3R/UWk/ev8ImmyUnMKrvkCtZYbkVf9ISm+Qu/b0+aeRaXTSwhnaKk4Vu4eaSCRBZTeJefuDgKWXp
PPPy3oX271YBQeyleMHZzmFLwgx+zv8NUHPlpVmdAVNJoJHC+G0TsYto10nrNbhzjcCd5J71sVZi
wHF53YH30dkEfaOGjHg8k3KXvDaQ5Y3zd880nIImKllDljpX3CjWtNs5D6fGrNljz7o526K9rtlz
cuD4YDnq8mVNMZ4eiDJ+mYxj9nO70vCuekJwOk5bmkYkZQapByArGJjcrD3loiaqi2D9gAF51OXs
V2LIlWtm4pMe8bwKbqg28S07/ov4JuaythLkcmxZJYVJx6Jib5hvmsHxlej0j4d0/DfEtIKepKqD
3Ub86UWpQiZ+SE7+VawXQG7zSMgs4eW3irqbbCjSsntcLrwuX4+JrpHvArlfAmgY9pBiTPv+fLWQ
MWjvSiUt5ZbKZUYsWl0OAjqJJCfEyA4Xigb79TzMMa5lwccYvyO0GyT4/B+pkM9qO5w9H2l7OT3u
MYM5Ezf40zoJ4bEuDofMgbxT7gle/nvhg4k+yxh/WAJzr7cj3wOf2+ZuMjJoXZ6p5lY24YDt1pyh
rbaOtvLELPe7wAX893nc9DwITRK+Md5OrT1b4ssIs6URezuQsjrl2fZvQvvUNiwOrZuy7+2vu9lu
WD+C6WajkeBWoqq/gLT25SuBJ6uiBg+sBEDw5zAcFOvPauzxFk+2o/tofJ3ydMGPCQguFNQwJJ1w
0vKW5AG96IksirOrBf7SrLfSG+KqPVIemO6RluUpCbY0uwZEU/j8Wv+iBSUN3jGqyOyKiAw2V3Iv
AcFfgJIIoaHeA00EOHx7Ss4OXLsSJiy4/S1fbouA9lVj+2hmR7Uc/xc23pFM1+sh7P4UqqDlBj2B
PTylSL+F+dSBvfqlNJUkwcqdiQZFuKR85JBPWDQ38W8rCawsl/qRf/XrNxgnrq94NhaTmdSF48ky
gGsUBLI2OLKnJE6u7PY73t3sXupuajbzqoYDZyBrq7EDUOrH8QkHN35ILO/VlMDrSEtSlEd6j4UG
Qze2falY6RiJ8X52ewubPQKx6JFP2/xwCh66Der5vxuIGS0jB2hsbhImInz0DUZ0anxz8X2YgcCH
gzZEhofQdTVH35RQASePWhjyNkeGjwh7ArwGCYyPEJ7gGqhPaIgnEAvPP1EA6gLF2dccw3O3mgnv
rx+DZgCN09EQYgztTmgvgreaF6HsOMNi7A+srYD2vgjzNlvlxLmIAqKvEAAtJWMZM3vRKKuslMMK
q/7SVSRq2GAZFet+X4pK8SBOqTu7As1eGz+6xQR++ISGna7kkpOxKdc+hJ6IUdm9DuOOwMsrJUGa
8bJYzRvWOao4gqAH5/gVZAiJuKT3KAdvgkklySUGeJn6a42Z4NalbqvZYBJLNb8L6F7EK/iK4tIO
BeW+oYFsQPXZ6IeYM5/PbpVOolz/BfsYYhUin0H94xpJ8qWR1i/kke4UZkNVmvABhlRzja7xUHUA
xRS9qDy8sZ7xHZJd5yrcUCQbDTgePlqyTHcWQcTR1U4nCiYpESMUBS0Kf2H70l6yu4CI4hg9OHCY
gRLWtlLS5+DpjqZenOcj5ELKRt9ZTPGM19OxCU1bQNZtZvnEITgBJ8oRUR8DuxvYrZluxFbR0q9l
BactgQRuU3DnjOZEQMkrg9K10JttjQue7psoMRw+8MzO++MELt6mH+cguZ4O+ifQ2gaefdlby1hX
DhGzrpPeqRvV0c24iaI7YHmKQzVMsHxPwb0ZYUWTYU08RVwnTP2FSHwiODVULr4xuVWcBJFVhIdS
NGmm3mrpWaM+qa+l567BpBYjTmz14/wyp1AmXy+bDFBv/KGFOt3J0f5fuzJSxtV1d6UKSabbldzz
RZ+2UTAyO98BPcrftSypcHsY9KblpAnW8aDmiEir+teOsv2etOjHeuXy6w1C2h+6lPDtssZER9P0
mHxYlDillMj5H1oTt5xuhnF6o0ihnK1/LKEAD6/5xv5Hr1YNR/6ptj19vlpGTbiParyP2vInXytc
Xz/j8YR0pa6rSh6nKl/N3Pg97A2Spyo0TDimWKGBa1K6mEbf2w1qVpPiIIZYsyFctf73MaYAptJF
B1YuRzT82C1852ZXBXv8ylbLtAIQI5P6okj1AVnbx818wlmA4TAg7zXtev4ojbLhl+qvAv/fZqH+
eFi8MrEJkxiSoi7YwMyfss5toxo10n71Zrwa1MYg4ZTLvyRI8ZZyFRYkVLGehvHfDXAO97dz/0M0
6iJFfAtUz4w0KLiws2oyPkZ2NJ0TWmS0WQ+qUo3wS3FUsD9k/0FcmKboEnNcWfQNGutc7xog9T8/
F0vqO7k5VMh8qootapNbOVzciAirNxH79IwL4xnQkRitNR2eLb4dHInqBdaYWBt3NTQwb6Oe/If7
Xnz2wclb9awkKTO6+RLq9M8MiRe1AgKLvlSYEDOLPnHl2zA6pw9akyqjNiNgPR/dsax3WByIZU0l
Rh/c+IMSlLENdmk1WF6PN/TKAEkFovGtUhhd8p3Eb3dyhQwhbKfu3iNvJFKM8iyj1K+jFhdbWxZo
7n/DFW57RES5Lky7AvcdHcbWzIFQrWEqpp77BpBJ669twutCiAgSPrJs7xNR0VtGERzGSJXl0jL3
DbxroO2rsQKJSUL7qHWrtcU0jIPe5kT3rmOSLlnJURyw14jqu9ZtQyRsCmVE3cLWJ+RoCobbB4V3
RctW3KZUXUj2adrECBRJ2xd1K7tLT7Lim6PQ4sy8PMYdzCRaMA2GXHkav2eiV9Eaghy5DhJ1V2gC
ZBQcCGtRZF1xgE4qMfSEhCjilmgEaD8vINJvYz3zCZnwVRXVPhWhkcxTVNmWYd8FljjM3Um2R+K5
87ruYhTh1Q9fzGQcir7x+5riQ8SA54DJMpRh7dOc/hmOskRxEiwNmzy82J1Q/xNRNch71o8+ghLf
UcE5v0NFkLci0DKg7oHcFw43L0Awjjbylw2WZQdEmFsvCefzEkm/1sEf3wdG6DF9bzr64M3ABR6o
YkErtN23FAKn7Kqc0VhLCDBuHc44ul/5qvnvA7fTBOc55NpmeY5Is6m7/JJW6bjH+IjoCeqWH1Lm
ZKT4pofucYT3W6a2Lf7cTd7QROSoZbSPVD8n6m4Rw2H2WnFlIRgQbIT8Wb60
`protect end_protected

