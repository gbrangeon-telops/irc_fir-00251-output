

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eRz+leRSRPpou0Iyb6bnhB8hg9kPbBirrzFUAdKqw/be3+N8ZrhDizYaLfXqnwxlgZsSWJCzRfM7
HvMw/rTLhw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rl74r1iJC/bnSjzA+Rx4NZe56NnmjoVRFzUux12uAkwgT++rVuZ0cWQxVSY31Gff9TGn02lNxavo
U1xWF81U2u/Zi0XY7ZHmbpbdUEdpSv9huiEIrpuLuTgWjBSUwsGYqRxHLx1vq4vioRXFlAhPk9JA
iYodwxjKI7YbbZElfVA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lO1ylq105LQ/xiJNZcB3fPTy1RngsQ3yQ/KJ6FM1qs+SoXmUQjQaEb6hJLPAypYN8r4VdJAzSC/U
5nFe27DWNjEKmiIleROkH20okne+9N7+PhPIZQnib521U3SV/ecBImKKPYRpHhAeqE7OE/DzQFWx
10ISqR1I6WBii4R8gkz5k4dkFHhiTU6fgkIHLUXXclJrpQ6fHHlk7MPcpQDjK7bXjIiQ81qfpVmp
P5Kh8wiY7VppUj33GlIcYsNio8GAIV3e0kBKLoX73uDqdvJ/2zBzKOZoDd0As7C4AHF8YSixL0MC
djalIDRCSOBX8Rd9h057rIe8ZIXNMu/BHoKk/g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aJoUzTg4Ju9hNY+ZPcuNUmGg+rCD8aivgSTst8VRB5/g9QHuzghA24ad2z08gxWDFeIOT/HFgT6H
g4nDsyLlbHK2gxUijkJ6ORkRfGOxb8UwHTzLEIRJ5zmkHtJXYM250JOsiukrgEDT40HqdtSgre6O
kXXliGFm9MU0LwRby+I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ca/+TaSll/KHF7mIE37XMZRKDQpSdluwuJA9x/CRPHNmOrubSxRKoPtbXlxVM6ehE2hXp6yB6qBf
Fup9ZI873BFwgulDsuQHuOSUPGo4bBHwDnNbSi/4G2je8uxqj4KeP/bv0RKunNMT/FTascQdDh6n
SVSARZi75+ElUvhBfAjPHB+yugMvSxDk7TRPn1RomvNtW1CJTL51/PQt26FoAtnxmwYDcU5wo8WT
ATzZmP4jq9ClSvjXHkf/VnlLenBFunDj22Ef6vdvxByXWMZrDdZyqqIvDvktra69BBPdtD2LNyW1
FCI6v17qDRdmShLAB1bJHs4PPkDtQbDOwcgx6g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5040)
`protect data_block
bBlPcmPUMjm4Hx0pmOlG136Wn0WGqQsnzXVMIllZmLcX/JKsTmKpQFUlJ53SlBDWcAjMzQvzT/Dx
2FGmAfRklGKj1EQh95m9qHuDjxWyvuX9efGg7w7TxCt4d3iRVOiomBIZn3hurxZN1WDD9lGN3dCp
GemRjYJo3gnvOv96BfqeNStPSs1epnW2eIidd/Ud71FA8+B1Hi8CnqOlcN3QBz4HxSZcVw2zeR5e
9cC646tzpJPeTD9KHt8U40SylAInejS297RVAufdN9cIsMds8ituVlwwV2wbuX9hqnRRG2vBkKAl
hibCy1L8VcJJ85YRqL+PIAPAEL55nbbaSbo1ul5y+7Okhwd4RIr51bqOGXBorgiPZ2LsfxiNKKgP
LBbo4WQpZe085AVB87kfrFIGL2jCZvLrJu/c3C8pPtJkh6KJzMUzib0v97xczlS5QpjxZ4A0Yz0/
aXg9xhCBjVc1XtfMvE7F5D7xWcEo7wTpm97lZ3HzIGzL9DGVD4PpOiwBX4moNQQErfMSVPAVUKP4
4tJLdrzk/62dVmgHZGUUXbXSWmkJf1I2e57XmkHFxrGBqbWrCNa3hs9LzK4bEeH137+VSmiSGzYV
/b1muLezKkIV9wINOAVRDz85FDVJmv0X0DFViUcC69C1uB5xZF1fNVT8xBsj110BtA+TwE1Fxzak
61DJ+woYVOS5YggC5RStVjEuiGlMmfOY5P6OBI9UAklUT9pqh3ecC8DixpkfL/QjUiaqpHBPueRv
TSzBKCjWC4lLOvvia3GBlSRAiZ+Ns1/KjeWUMQbRRRoiRd+o814kpXGLW3plJV8rSIQ10Wok7XLP
YdPCiPrgMMRUdQQwt83OsG5bZe7b/FzxHLJkSyq6wsVQBNLUjRVLGeJkLISenDTofV6VfM1DGJq3
p8FcOM9YbeGMpRvIGMbyJyckRzHfnd98zgp1JVxjV+EDdlslmcLs0UdzwpAZ4OyxPlNP4KbTYBEU
coPyEoc20oqXakUgxpWvJuRrrg/Or5mLIZjBCtDmil026DLwe7EunTM4wwK6SGVr61O+CZUeir23
cZEibSz82gejWSEl07V1xTFQ5yxPqpOxI5qePrGx2f4xWsTdz+JCwmLrusqHZInPQPTrjm3Tg0Xb
yGkiPPi7WpPfoFBXqHFzbS5dB77vVJL8U85gYJMQbv8fQjSO841yHrF/3wO0ZtBeaXlEl7hZwDZl
BP8N9hk1O3Vtt8tEFTB7ENOQy+5kGzXOWYs/oh1TGP20uFwXItGg7GIPtFJzmv7QIJLmOrey+vul
x3bThGfEmuiTeroXHYOc1z2CfqVEmVkAJqqrm/vKFsJFxhGzdUPtK1o/qHzIkG1l9lckzyRWdrKC
jlW0AicpIqPCLcxbgp1UoZQgEHvRmsSDqsu7hcn/5WIHz8Yk/OOQ8QZRUFL/4GKOVnN2V/yyZiWs
oeNJwPszDTWJNJnBeH5s0Y9fv5mfX5lsxBUnYZ2oDyBQqkHCw2Pop/FMaRIOqUrpH5HUMw9FE/F1
Bany0lrvXHzMCUfo5f6chl+05WO43ojyhVTKeW/GULx8F5/Di7neeyvQcTU5cZ+zSb9sr7JREp9s
29QyTjOEx3XpdgM3k8dCl1J+jE3d3TBajq36SukEiQAlb2eudh+LTEuRbJbcJYfO01OvzwPVSe1R
yV2cQC7micPCmU0WQ6bpkbEpKa5N53GtHxMZaJa2lG5LWBOIG5dIy/e7lka4EeoO6PVxwfBsP7Ar
xs1VG5cr974JFFdylnzK0OpKpx12tJ+ep07yJqJ0QwJ+pGdQdtdYamj2LYMIn0rlIhJ+Cs96SFkU
e+b1l2dmtC8JVc0q/XqcyD3jjl3jCtl9UwsGs4iD/O+x0LpdBx5WPrpqkneazP3Jprw2seVGvt4t
WWjOBsg9yLCYmD2jJt/ejEtbvB3vGsxa0rM07vZEQHc0dcaVIRhoQuE8l1eisls6m/fNcxdCIDV1
4y5bKPAz8rrjoZt1SdNCiDHwSY7ttzC+VYK7MHslDlVA8LoY3G5RceBK63LRlXA717LlQL/4UsPK
G36QBl4/KWtNtZKFwiSRal5flgWF1paekv0zTHZVU0FwKOpFX3mrWZFIVwg8rwKITnh3Tzsg9xlx
sKb3sNU6QlfjYAp6lmqx76t0JZeyN4AwRifCmMdChTOZTSVeaaW9sP4Kphmx9MY8PrNLvXrlEg9S
uY4c9FgpY6lrcrdIWy9hnYX7L1XwHnZnIZt5hq2dK2p/ZdjpEQalCTcM9R70oHvfC8gYn8wWPoXL
FBLYnHPX9myI248ewpRDbWueif8V9SQM+ClaBi3VniGi3srKczP6fjD8/Ycr+ge97aVmH2FQsIDy
rQJp7/h7acu4FJh4d5MQqbux8touUYxIDxkCc0TA3N5QGRY6fgFw7h5xkS4JnbqvFEOJQhxMUYia
Q0NuPCFXoKrj0gHbsAGoDXju4fw0VXlzBXvaV9o9URo2Gnxa5tiJSRhy/0hFm9GhnnqYSirD6pal
um7KxThYGuWtzybvdtlA4HdYTKBCy6rqc5Th6tso0DMjFThUb8Nu/z7s722B/wWkr0lTj2bdPHM6
N83F0RDTMiwazpkkYcTKvtEqhOGrlbQaX4ehxG96qV0Kr1zRbxxLrJosci3elzquByikOwcsUCR1
MBiUdMBDRrVjAIwnCH8PvYOuw+AP+KgkO6IvQwKYEDKxcL9mRxz89qki4GxfY9Fx2E5ZOs9KSQm2
a/kWG08nOMFuROT53QzsvHiJuIPLbGEpDOoWI8uEpaOlPCy3z/zUFfOKEtVCkDVIXAwt2z2OqNXw
UAN/951DglE8A3tG7RGiLaN5XBisHEL6vodCVXmGzZiW4eYJKQ0AwnjdDRCRuqIDmZsc/RLN+JmU
oCavMX4P5erQnJ1IkA3qMQWzxUc5Z/ZbpGrnQtRsTdp6eRQ5L1ssTl/90vaiwG47YKj6m5P6/gb2
oIeNZFOHjp3UM2w0DOuijCkxK37WzuMUtCnI3EmQyiT+rg3YqBM5202i/j3OdWHY2UsZy227mHgl
BseQwEgxI7JGZEA+SBgEmKZkryc7W7hlMVJNDEE+pjdU4Z2g/cFV49IGlLkVpO+gkcj3d/VxgFuX
jBOgHUyHv4kt/tS8O8kbUfHu5vwGYgSfwFAa2ve7T8KNL5hkLr0rhzN4iQuJS0NkeAUH+WGjchmP
GBTKywf1j7nCFG0ZdJrFVt3ptYamAxEs01czs5tIXKIUrYlNUU3dU03As4v4DA1XqTGrCIa8Kgxv
MmUDdg94M5u0RpAXFL00chmnZPUsxLmWMMufDKbXupU+vn7dGV0Qegx9gCWlzrd535B2BN2+A5rH
AsaH7eLJCLHsVcLkZQVFQ8p56lfLNjA+ydszJulHLdKiyCUHgLAMedNHRQ6S6OqE211c/o+4Ng4q
UA/9FjnjH90oFeUyUcKH9Q8XHUrRc0FU+xppEusc5uiXfYb3mXE7gY4B60iMe80iuqRsgzzUeURo
SWBOcO/BbKrPd5TsIJc7BWEybWYdwBbPdxVEcAlzRH7zz4z8zhy7Ab5SvMrFZtwRQOPr+lMl9wKk
gkFjLUaB53pPQspShTcIjMA1bXE3FrDcmlbuMU2z8uTrAYOOEDek9uy6cI9zrTtYUr5keFndGMJo
J4IB1STFIhHoy5Fpyzof9IqviTqtbMeOiE6k4s06sPmjQPEYvF7c1DHhf9SNWu86Uf6AfQ8QZSU1
K2mdvDOyodqn+xin9p/bCoZAP0s7ZD3yln6uosT0tOI5PWdLt5YzcGGzk/Yt0Fxq75jINk0mMerf
gS7jN4tzE3cJc7AhAQB0BRNyZlYlGlCY6UaiD4IRV+GhRXdx9UukD94dptkOk3UxyrjxUye3RHj4
SKfFQGnBZdtj8/YBnivagDiiJKIqVzQj6loikLn7XVvae0aZGzspwimHTlQ8RGubbBeAvDSEBFRt
YeHb4jY958xp90onPJI+PKCH14hqNwXUPDOmQIIxIzyqsBt9DyuLZ+i0LGnHNfqexLKpnSCbqIH4
cbxbKDJ6Voaz6bAHMRxyyQbMdjZqaii2LKeyySDAJcfPPI6MMyZCc0/lTVIoes7bpAED7TJWNoC6
U6Qx+RABQXAAldWugVvWBAbwUTImvjXwhUQbnrE/GJlFaG8G2Vmnl231HM8BqkyRWvUsD+zBr4tV
rUj+RXlIoYofAdFspVkgCpGdgrOzjKg1Cy6uyiKqf8A78CG93YkARZgi98WQm/3x2bzHfgczfJN0
ZK+kv+2Wjo+drMQ3P2CgA7qadmoYdnyE1dd7g98a9/yjolRtvVWYzILZlZ2l97dt6KeWXtgiQiEB
TtH46QQiVD4s3/onCv6C6We7Iyw5MSvbolt1v6VjiwsONkzBwZvFUj0NuqV9V6jcI9tsRmWReqRV
Pcen/HVjHTPnHD6C64xHOFw6PcqrfTtY9JS2UHLzvzurt/hCTk4JsEDByY3Fkm1QLs0kbblXVEmU
xN9M6Y3iT7rtAW/0VR2t5tCAAVynM0Ydlfs2JwwV48s1uPCTq9X+cVPmauBEimlEHFOcHnH5TPIR
2KslTbJX2xAWdwK1ei0eq23NCOUUJ1LDtO2eCbnfGdxhQrd5U1tY9fXbRRwMAbiE1Qd8FKUpIivb
b1L5ey1q6cJBGwLi7fTQ/8NElQm0/+Jrbul5C08IqK2dn0fEr+mvkPUNBREbWes33NxMjr/XbiZg
lacHv7ELW5LoZdyYUMBZCyFdijinnVCUReg+dV+ntgyRm0kYm9FJoNq5lA24618ROzHenBXz85Hs
Xv2r7VHxw97M4CViE14VlJ+UPeHTnuzeemWJZgEjg4pa1fXrFeTuqXhxDDL3K4knT/sY4bUsWQr4
qPYR83c54cLnl/g2uBxKv9+ksSFEleuMwrvWvtM7hDQ+Yh9u2asovPhCj3PcipMxxEvT65Wuvb5W
xij1drHodZwbOLMX4CHIlWPySIvIbOqYFxs2Qsuxq4LVfgx6AM4kW0HJVDa3S50nwy/P1AOn5prU
b7daVWOs52in7Gj9wOTsWCB9GH5NulZb8oxFNMm3DAJiJin+YSW79bzsniu4bsFUTDITRS7GKNld
TZMOfT1D1B/ir4d3PNqUxhewOoKakG8PiypwMR7BElp+vNmmbpH+nCj/qSZ5TpF4uxjNtWS2IYEe
mv3UHZ6A+afpGPz6zAWaq58ua3Mqy5u11EblguuQ7ULP13eBp2c4W6PfpAG9+30HIA2DHWcXtoUM
SON8waSdb368pybxf20bomSaYYz7+63EWLPRD6zk/jeOx2n9QAJenkqK6DZLTsMJ6TT5vn19r0kj
t79r4CSUn0/vsOkQYmTy08mV5Fhmrr2OliFiAJfgQs3lZjLbjqU2Bx9UI01XPBj/L3ItmV1/x1XP
6XdRPtly/VPbSEBiEKy+EP8QXdCHXwgaNOwnRH40/tu58CvnrX8yk59X7zzT9lONaGMeQNhbciVE
iwCvyeGTMbFFzhevp9YqfPpDAk/UdjdteQJxkBk/IvVXw6tSEaqzqnicivL9cD90EHTk7+wmAH4W
AgYPvawcJYWIISaTS7iT4O8ldsV5tQWAKqaN8sLRMV4DbAOCmylnCBBdXV3lxJwgwBmAg3BxV7qE
LXGd4Ccld/F4R2Oe3ngx7teyZQH1TtEojJos6p339j5y9KGN2uKeOrUHSbyQ7gM3er8vY5p8anoW
YIDr6t23BmlGTOcrxz4lYHwfFXB7n+FD5kQ+7+iNOZI1VaqzirE7Z8NBYZMapG1syFZdy8TAwdkv
8zYi8wTVb5dTc3h+H0OC4wuSn4/zJl8IfjdYYSfLc4HyD5BcpXYEkiTSeYItHbyiA8OvLl5fZcNk
fREhyYVuOfXnVrZbjsfFf7bPM2PWlxS2/EZ5O4x0PJam0O3RwQykbijSTto78PQ9hTJbcfGSuXpZ
cZmqnXa2cOcD7UuQruoQcor05jMr+nW8K0bK9n3LlbV4MpTF1fp2nW2pT8mUaPlH0/0LXO8Qfxwx
ldJitWFUBlkOGBZ/yeBd46ucOjTUibugtOa4SYdsmLlPbkzuaA7xFyFOf6RdUaNUQfV9jV+mRUEx
PQM8dLBU8fxabaiYSdCMc4ljA/LewFziWL4Zg3tOPvcfXRsdM067sCm7zTFL2LrJuL7rBGKkkR9T
oNusEj9rod5EDohp5WggQ7c5NYsGRb1/M/1RLDCz6Wv78aMQ22W96okjRn0QEKZO3HTpz5FGSliz
Q5YN4YiXnx6sGHbrNqzvg26jqwnuPHtPeQgagzCwd2bvd3fqxCBuvL4IpSkmwGFIWZKIBEEefg5i
AnofV35FCcY76zj9v40PEw1g4ryFf5axTQbYZBZoGdfN5TxoFNxnpZM8E0CPh1XJ652Ma29Gi0MH
+7MbfoMttqxINQN8VadcXsesDm4lH1bj5EJJa36L6ir9RpLj7OT7dPBUq9amLCHVL2jitf34Q7TO
1SJWdUPlAZj2CviovIlu8ru8kctOHJH+u+caUTFk4T8vIVHdN2hXwJuAimPoCfk1BECsesQf+Z6l
jfAjJ1LKi5oeFzrxPJj8CDP3x+uHSdhmiFdB1bxrijocUL10IaKVG1DZv/WqCjDE3WUQ9f+SSIl1
kR1svj+Llnlb30K3fjKYbKADxl65PvSvrv2YFicBW9g3JCQLpFvGRsDj/9Q5Aqi83UDdDni/FRKL
efvwAKWh1G65288LdbNxd7XaI/x8wEEl
`protect end_protected

