

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WrSZEf64fUAl1kVl9HWWVm9JOgHMmzn0fv0uusEaRSoZ0YHKAX+sj6D4gL2WXWrV9+rdMofvPwNs
9A6zs8psHA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R/iTmfCVAo0uuZTRynJ9b5Z2gujQ7+Xxv1u+96JME6mwR6F6/MPV4ayotodCx+xcD+9l4Ktib8Ml
C05jFwQ5vFi+09RjQvyvxQAR5CtE87QE5Bg2A3Gt5QmE+m7ZfJiQZgi5YQHL3kAHS0jfaofTkZIU
6VFVSW/fcrod0Swq7VE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RAfB7dvLyt2uCWNWspMeHiLYPG4TlOk+8Dptz+NhWH6nMzYrNkf7IWIjXk3hEVf7lwT/X64pynoh
QoCCtl9AW1iC77VMTIu5MgFRizuZMUfXZ0crSPULV2aGonx9nQ5JKx8TiRv5BTWxeAsuh1lT/5p6
2v08ZCt1Nwa8GPmEeFnTZsTB1B0jFzZQMa3GGdV0nEcSjDo4bLIkw9sMEBW2OdUuvE5yIHF6Z7++
/wzulmNKOqQpmeHrq3r1VKkMUHNzsDpLkGo5HMiTmEUJr/s3uq2EhCIq1agWSVbcEjS5uDaYcwdG
D4cRvgOxtT5sxpWA4fivRX7vvCyun+C2e4pYew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MsyF52v9pEo5RpJJtfhlgAJQ/9a172C6pJMP5S/aXQMuRuv2+JV5wCeynUZSXHj38Ger421EXuQd
EmO2OIKWiz2pShaEh/NwF+InGDF0QzD16vAgn24LAOYAOX1lcCquf4w2rs7e+0dn2PO/GYRn4rxl
E65F1qdRiZlUeVoRHdk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
klspBE6zapxwDIEksFW+V3vEj3afpsQxyK1CWGpsw53FDriMhZB4hONIr9yRSN9nitmQ+6cnlGM3
S4Cxnkb334zdXXX5YoppEYaAdCcB5nDsYhSpn4PyPhd2ANmiSIXxEjiEJ9MDJlVIobzrtkNgFEWA
QkqC/Eky3QLBOqPuDJIgkf5UFynGEkI3eWzGSyuNAHTTYXfoLlYBh8nelaKS5vgYh7jpllyo5l6k
hn08k3sWZKuN1S8dwb88eFGM6hwg1UoX7pTnUY5yGPZZS0JEiN6WVWRmh72r5l3yyFZOFNcvByJJ
z349Odlh9AHKI6joGGP9sLtbKDrZfmu9y/SSsA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22384)
`protect data_block
IYmS3hg5eiSXEu57sVm8F4YmSVJeYf9bKxSS40P2rPQ+QwyoaDM51uFTwmpAQDpwsMpLtAJ1hZz0
MZBKxIhttmlW4nEnRXV3paWlYsrTLKXzxcqNki39kRPFQ3o9CqnnR7nF5oL4J/qEsKhApxxo82n6
Bw2Ck8fPVYwEoqyFUBv/qZSIqkIPhuJQBHiqPx0hRYThTqZmQfe92s3TsEn6jte2EdSfcSDkVccX
/fPsw6ZA5o1xrTu0ynpTcwZgtO9oZrV4wqt9IcyTOTsnY2CsvmYBufbNke3b1tABNuZlJPvrPTPq
LIUnJsUTXy+IRw6IBXCuu89RqOZovvMM0mpBZJ47P6LRdjeFHqZDPWP1rGnLTX9nCyrN1MZ1R/4G
Gzq8J9dPnjXwICcQUze8pxRfXeypzV4o/mcSQ9b85Ak9tl/cpUZiAVIBetSaQvAK8yAquoRyHXA2
NOkZoVuiJ72M07bUiNw6hHzy7QzsnQJdrvn135Lic8NmFSiA3YM37iGr4E/MDO5VXy5vfvBqHC29
kUkIghLDkP226OrlTF9K/c1FQStJh+emEPwB37+4OljXRrvn3g+1/J19NQ6qBXhMfXx/jY6NkU+l
PUgGOLAknErrmh+RQ6XjhnzjFwyW+Vc7yg5M10cugkeGnmM4U5qE7hi6GWh0dAaYiV6et+JTApsi
ZvnzlfQAJLPKmcbhmgnh3OFHENOfzW3wBATtWfx+LoYXeSX4BFzJiPZgs1aUCfYH2MDA/NhMOKbY
OJyPXIiMTxgajpyZbBmPbykQJUFuLOvY8J2IaZVeFpGUXkAQJX3PCQ6ZUzFGUSwaRTHHjdJQLTHq
WxZtzEnT+8+C9IUMx/snN/Vg9tpcUW4s08iiLKW7ZL1MfjfuygOjFpi16Xpp7rOfeH0uEQVal5YB
/OI3SCaBB73qFksl4zU/uqwUQ6QLtCz78aWpV7XwmahaI9H1K/IMAq63kNjDieOK7/1gxiUjjD07
ZUgMFJH45gE/FKRX+RU6JVoDzGIKd+sZy1MJeUpKzKde6RzHG/pIaHctxdVv9SXFWPILJ6RJpVuA
WL7jB9lgJ6EGoHrfxMYYnUMetixz9MaeG8VdwLOtUXgAWc82MtC4ScHy6Azm4jjhJhafuPf7Pvth
3mjuVk5k1EMD7RClcIR1kwIx+KrGl8ZARQoDuOpCtpGgSiI1Tz3M3bzw75UUNBVDIhl6xFpGL5JD
ShJflUnSFlYZ3pi6YLng9su8EcTKSDhuM012UWJasqG+jT8T9gdxNwimwMyJvl9x6ZnxZJzKtsjO
CmeGwUDACWpLGhWmeXQYpVcoGUMsBoG6/YHSChuA4DjQMv5REC2/NnxI0RPTiZOZ49Z0TtiGp82b
AFuq/SOAN1O35+lij74kZpnyS536i/zH1NDznymKtHY+YBDusian7VdeYeGcsRD9zFMic/YYRI6r
k0qe27DzU4kfcDtnCbmykgr3f38laoxPpAUMSXr+5j4JV1LQfj9d+lzVoKh42vx5omMWYFve3eep
VHRYctcXnx9Vyd4pu8LkPW/nWbWdEVXpUPa66VNX7y3dEGTxy+DgnRBJOCWuTCR+w2JZ+gpvOM5x
KlyRtHBAdvRCzqcYYPPf6CtNBgr9L6RuafqHi7PFHWdEsIB6kV+NGkvUYhAivT2eNsRIp2WEbCsF
WkU+KxSmxB+C80vvgcw7IWW4mnhqmyaqLXCkNwtnqvjMmxgGQeXJcVR764R8kSzfQMOuZYg9EUJg
T9NnCpEUeER8Ah+3fK0goOVWn3XGnzUUrwfm1Y9dfGbcWmvdAjVZIMwfK2nkkl93DAsKFb+ka7dk
KqoXNRjMZrsO3vtunTNGEe2MQzMkFTvd3BcAmus9Z7mw1P0zohr8eitEe1TtzyoGIbeMQLHSvoiR
34oz0FlrkhRFamLGd/p9DYtPP68ov8jKyW32MQK7/IAVRgCw4Jkkr46m0TWR+ynOyiYH22xesC6x
hWSiCTf5+PfR8pIPT7ejH8zrfGuexKxgpUAxJ89anDJXcU8iYjt3g8gNljqrVac5OgBZylg7a1tj
N05x3Uld1+E2lg6nBv2w8MNB4rYLy3oKK1SOx4XruZSg1u8jk8kleCdYY0JoeFJYsqoJ0PapJRRz
gGvCP8itb/T2oURvbNZjqkXpqgvikiCtN27AJXfjRwNTARew8az1TgpOrqxNjdOsHs7OfSSEi5Xw
0G5fg4n3Em7xvBXZyWKGCXDaAKk5/qNs+xSL2FOKZLQgYwc4yORNt2j5Bgw/mP29dfHChPOQImHG
BmTjAPUJsc0/5ZjE9GFFdcCfGXwhXdWuz17c09hQKXFRDojhTX8KlLqCnrYVH1MnnI3Ik+XamvM+
OYNe/fAMRBBPToQYsXe9hNTIlmyKHWzTiu49jNTnG7Z0WCBhCMCwUGssNG16GPxJv6Hvhynpq9NJ
BlMwVFCMt8Zsp88OvKWulHMp5+n4LEqlSA7X9fmP4igq4AKFo54oEYj3tVX6Fy9XGn4pNd9pLFI+
vUwhUkCWrqTo1sH8T89EYXtGOYdP19R7huQE1zqqrMq68SbJPsj0aFTDyiV5ZRjBO2C9CZnjT/nu
eRYiatQeD3Orqh9C8i6H0DWqSqjNtFwV/HPrKKXOe7rJA3wBGqvV+kRxXYe3aje+/6Pl96ClViCr
fldj7O2QkORcTxY7btGGlbeHx4ukDH3ceR4SHooNszN9dLVykfKJmNbynh4tmq0M8ILd8OHxWOXt
CdmOJgry5rMBWJwQJLZ33M+/q1TLCxusldQ0RmqiiMW9FJQP6wyG/Uip+CdS0bd2oKWRa4VOcrPA
oS3P72yAziQBeeLnG4zpSt3WI8UNN+iUBIn5XNTKKvYfmDJP5piVGoG0Cqj5XSn80wKwvw4QGEOT
XGxm41Dv2Sl3lWmQhHenPclJKxDU4OfFuHyKQil+HvnoSVskk8QilLq2IdEMWvpOnySBU6jCzfpc
cZFx4OKulfQLQHl9iEU0JhndziHE6X2Z86KYt8clJEL7Xb8gZlxBfbfBA4iOrKvm9QZqGd0HwcRf
dYWNqqdbtNQe1HibSyef4McF+hu5weraBUhah9Jm7ceqL3Ij+T4uVJLYK0M0drAFwF4tfmbXXs12
YEQYuS1jlzd4RjL4q/8SYUqFVB6TpEbfRopjd8oGjcV5eQbqMpK9IBlC9PDOfTEyaOk98PDX7gyx
P5TDP+Rce6gAg6sRV1RutOegnvU9cIIv+l1DyWM3/XL/iSGnFtnQEAScEbC3w3GQJPPLYOxhE1RB
nOoicangku9l/vfk4xY6SGmtKJ3fR3Gi5OzbBX26DniXcXb8d/lpBwA+lEdaK4uYSjKFHm7Ba6If
esHuFITGjqDfNEfADx0UEzt70jP8U8RnJTdhQVo6zdbc1AhacL6mtMI6oz6cPZGVW1NONYilJFki
Kbircfg9grFJ9XpufDCnZ/grcRIPhg2nCdBnkXJ0Vq4Lcg0etxb/1p0A0gbiXIHJzKd+1FxLg7VN
BoLNs16B7Ts0o4I0yA3U7mI4dWM48pc4tYfPE51u5rk5EATCSiJwlyKPhDZPYCMYw/XIuUliGX7Z
S7HUn6/gIN6af4ryWQPSBPEIdxNyWgs58iiEvSoVJ0hvRBBNFiP3YlkEGn7lLwXBDBwzWUuM6j8c
Lq1VgfrilZp2VOdv4yOXU4FfOFy+y4nhLPgOIPT38bl0OCUQqZVN5lUluKu/eltEOFoeiI7lomKr
vEKHnFgPalhEAcOPUOvrxOXWm9GvsI0NwXsYDxTJQKdm8QRbMiNE2hxnlUCVazpnJvqOuqBKgoJU
coRV1InzeGnWaZg8e5X/gsxUJwydBG5KrJQ7YcpgowzYn4LnWIDVv5CJ3wPJbwZmd3GUyGvtPLcv
7P5x6BFRQDdEMYYdNWQZ5sqp1iFOTKYMRPKeXOTI/oQ8AnHZD73ZAQc2N/+RJmOR2qNCf1Silf20
rpzW8JQDM4h57nRnAYMTppFaNMbKN8KL4RlPIsWFL9Jn5L+TcT+aO2GkIEDP4825lEjcDJnDg8f+
+m6jfRl0oSzzmufwiHKfS3jJwz7AxlS/zQZpsA4RZn5ki7shGe2Xv6ofiNhxLQJ2WjUweR195ncP
kTqH2P/sEYGaIngxGISA4WbCB2ElfsFCXfwSx1cboxpu4l/HlIsgC7ZhNzCZSMfgltBMxrh5ceDE
d8+KMEUYcLWCcs9BZ+Ijpp9XjuGi0N63nwkj3mgJxTAcWL8OWI5/71ff7D/p1a/YWe4bfW9+qje+
fID1E7bMUCCMCH9BGKWLU0XUc/t9NKljs9C7F2lJgpHPPIGMddFmKCaEw1PxUy3r6w8INkhj2Jwi
kbtCOc92gqdzQCM9Ss8ReBJNfiW8baZhmiz9qh8+eZGd5HTYvfJedgFqpZBM0FOw1tyOewQLSTKG
cMGEQlnLcITskFtDNFZmbzf/rXOMeh8TkXTrjYBLHLv9b0gZhiMBC1+IzODGyrI8V7/PCf05qn4N
zfRnhBSEi0DXpU4ghZSJRnbDdozmBFzqZQ67r9cJnfFhRjEqSr6pvRGZ4FbTggK0TivivR8qO4G0
dxmNr7RuZnupw2SBBgpiCzyJfGiQhyaqvqCIT/Eg/IrDBm9L782aD6iAXYNu9COHJ39fVusIJsHr
9gIpdHE3yJxfmc9ayziMWAxefHl6GsBvXsCGS+b/gdJm03YzXIPWJD192XeVRf9q7zqSyv/Ve6uk
4q6WLc0KbzpCFyj7JSZJ2kh0nO+DMb71o/7lNSDnnkA21LF67B/dx083qBGkzxu3KWx0fmuxHaSQ
c5+uLAcmAr8Y2+/pmZcZd3G/6UVldcTi+p/1I+rMM3/TxK4h1PcIQ8J2BQsN9BJi7vTVq7nU+9d8
O90zHfSVTIkL8+AV2gfHQ7JzSzLJ85sAfCPy6pWNVz+clwBpe01vmT8xlpzOSW2QuSS7Z1ZlbBNc
0RtjjVM3TqKs3YpSxN2lNFc0nWjfZ9l1ncom9hvKp+7RZxmtmTc8/e+h1QG74fEYWO9B24BIIVfc
rP/ibLPiyfQ8NwsGlS+XZkys7uDa0gNxIVKpWoxcblcoQC6JzthJBbH/zQ6m0e3tkeg30BxNrtFf
Oc53yn2KaSuoVDbRZFIhAW1ws7Z4icaRZ0pWX4+WUfpYmZsFObckDlTUi2JrhgU58/uJ5hmXwpQ8
ouGb+8v2a0HquSp97EgOoXy50qG9QTAfg8w7I3ghJf8r3rtdCRpeDuGR5g8Id1bQcNcXPf4DlSnN
75b8aMI+kVZrdwactorNmOmc8AtPfH+O9ZoSAxFxloUUXkUGSBduhT3ZI8kg86HWJjo7w4/gzYo0
D1JeU1q7FmXIewx2+xS40JDSFouqG9AaTkQAfJAeUoFejFC5bf+Ry9ZGaFSvfYE4KvP6bbRZDPfr
tSYp9gTm+gnCH6XD+ZJ1WKgtNF6rmUZ0rvdPUjQb6//uhS8SOE2O9pVimhKq507bBmgcoVroJ5Np
zBtLPpfkKbBfHc8UoqDSKwa/jvP4YecT7+mZi7W2ytHNuBIMNBdDJN5LVGeZUAra5/608lj/4RJB
7DHzYZhY44VY+OhHa5BWYTR+YICtNRu8ExAwZIyzeZ7AJrRZ4kNTF4ScMi2zbTZkFNyYj/ci5MJg
8PxYdhcI2EBI3cTFd09+969SRyCKvdgkI2ZxoMytqnw57Y3PbcoMiEEaPL93lF5sIWoYNPrApmvd
BQTwelym4PveiEI+xCnq09jJ2QPAs9YA+je+ULP1SsLyEJQdqjsNifoYB9RXBwQ+o+/Q69xKBaGu
zjyc9e0Pux3TD/aHvK7B8YqT6SBStl1PftVRIIRmRDUX3E8CtMo7XQgHV+l3P49h+6P4D1Ou/SAm
BFv5u8qvvUlix1O54iIu4GbEviiFidhyyZ+pmOk3ch8YIJ6pnZ0X5FdnAnGQ94iPAQBUlm+J+H73
1g437OicZq7hwPTPpQBGjjWltnzTdfZsYrIN9lK/qtbfst4ncpASAV79cfjbZRqT1tzYdUEUBkX3
p/1tCngu38hnT1SPfiROtujoOytMhozpXTIdHCbylmmrm1s8n8bswqqHIMvhOxmV4+YkO6zZXvfM
T8NmPNLNaw4W7jx2r886TQOZspEEt22qtKfe9h8kVMx54LKDxwUg1wOOtahXJCHcWdxKOfmF5alX
zOrjLjkkNOeBX9Duc98gEEX4qFgMvJubW8JVon49Wyq2lKMpg5p9KNiTqqWVBkwy0O+eyzchwN6C
jEKoPtpOqBrEwgQt/a7SJKfTqB5ca6jnym7hLXwMAG6VggnDZzB9QlSZ7zpJeD+a9ldNOfjgFxpo
xeetSxCK1Xf6PxXfLBN6UZBelO5dzndAim2P6oT2FVpSgL9Ieo9Uo/Pfyy/yP8wh97monUqoPqiX
DC/7DqCmp6OyXUhoeizxUBfTCETQyqTtu9rwW87Lk9jlrixpIM0Jdiinuwv+amppKQDZtbCmXVbM
meR/S5VpqtB0iCx/hdQei2FwseZPmpGIp4nRs+/nY0ZhLijw0oMp8bySdmjaz69nTyTEAEl7CxIH
amH4xUPz2fc7sDQQyJAiEafmq9p3xrigZC5ZrqpuuvaTudeMSySyp4CTyvWFG1bVSok62kw3S0hx
JaYhPFTPO6k2GK0qrvfUac5QaelnxDg8s0tEv2yrPNo/XxYi304btLLxSu5qsE5HUWyM6N7epPK4
RYUiJ9fcB4Y6P2VYuNkLL2TA+bl4Wo+Y+tPVpWpSoEqBRSXfEGE2XIGkNSi0N/QoY3W4zL+TNLGm
3IZaQpKIuH9nMgeT79PTrAmVEJj54q2Wdy9mlI5hrER3xSJu0G67ph6AIyTB77x5b8PN6MfaCipB
Kpf4Ktzl17oIxIvkXAGpeuG98UKCEdJ0dWt6TK5+zF9wIX3iVSW6GRKdyw8BhlDeX5VB6RczeQ2j
TnnAleV4Db1CMHUl0EGLbAPsxgi2uq1bbzdVdnuI6XjnsVYt6LatU5xCelE2G3ROzehQQ7TpVrl/
dW4+LdOHKJ3ZChiGMyN1XH/d+L7v/3hq8smCPiTgDq06jF1xb1geORQsoP83/qqVS5Ombj0ACjL9
dRJjwbMhuWBqYU4ChIO7IZhmlPPbEeUmLiUKqpiTNNhowiHfmlom4AjH3M7KWpAdt+WZhz7BR++h
vWlAOGr8ldZ2u4QS/hbepGbYBqL/iwMxROR9RyIkJX68++cShkOejZRvyXwhE67/4wPhiqSUY9bX
4Wd9nhjOOxHebcS5ofN8Ki8vWYEq/guyI2nCEYZNtlwTDtfTLlHnIN8w6zdPMUOva03VwJi5gdMZ
VX5le71Lv+gmNvs548y28/MZ8RpeEgywCO6za0M+HLSuWUhSIyI+1ehqCRJlhiyNs9iIIHOcFsxn
9P2o7kjj9qeg4RH6OYxA4iwAXjQbEQ0QkTLT01mzJ6LY411b6vxR1p52h/EVS+NpSB7L6tvT1G+c
PXLuICb/+sEpRUvwOOo0Slll22dzc1hsxkUaTa6jn+0Rik8A4to0FSsgqT0FUfmC7u5JFsPa5d9v
wSD97rS1nzfOferMx1dHV6gm4eVNKGNvezgQgoU4ZngDAvwJCdpEePoaoqaJhuWRLtJmbizR9YMp
kkwZ82Kls9fYutRgA2Oh9mpVIkFfTFwWCFfUc7qENnB2fDnrs/faz55UAMMd+Aix0qIxemZ4P1R4
v76Qa+7hRx4krJZSCj/A2+coNWpvlNYCN73sG2WOpXnCChLK0GAGrbpEOsdkquyEMYAs0FipRqs7
v6StndZZgxJESurD8kf6hFETgWIEK5JUT/hAhOGszMDCIUPFJ7o0f7kME5qiMz2fwzmeH7yx10No
ZSE5T1UCT+6Uzsvj8i6tT9EBysi9VaJJEU2VvDU2heVbOl97eI84ZOIB+HHUXMWcsTF3LVa00n+A
OzZhJABCJdUDREd6hJUJPQZNkUtfB0WzE6JNHaALoUGWeqiS889YHNQ4FwVKJoKioXsFyQku1UkJ
Hc1Ued+3uxXe6PwlPVKnBN8Nnhw/G2vgTmh9yUOdOTc5wc6jB7DoESCXey3rlAX5CZ6XlprgwuPw
fJRsZRBGcQfKkTAPfe2R873mjDYUB/kF/nup0U3YaiKi9EfqLEHma/8HdW74O8XNP72h7saVuow0
cJJskFwY83vLhny19hmEniAXPtCQyqpzYpCSyvoH3v3fZLtU0jrZE9k055WraXmf/727AgEkpa1s
PogIKm1YP90iiV+xr0RR1ywXY/EN/+K0Om0f+wL58mibyfNXcDXVRO5Xye5DenEYRjtz7umq3LhG
F152No6JjcptACO96Ix6of5mEOi6IiUOXvGwSHNCbeIAf8S0VhddftDYPMBTH9jI/Vq3T8OKMyxh
CCK4PRusdM90wHCTibwBnuSf72FHZI3G5ROOYQ5N+27e2MejP0mc1U29QMy8N8dHspPpj+oHlM1W
pPMScTssMr2rowKOurCjvgElxYNG8EwRavcEczaseV90fv/MmiT5h/3mTo0LFEb4c98mNXPGgidT
2cD8fKEihsyUavkgLNNozIzncwLF6ZlwstpAChMmT8zycYmLn2UBLjspioWny9TfBDxxJTZI3LuE
oCcXxeCfzyLh3Qp2t6iMSmRqvLo/7sf6DIbNuI1mJHNPdUPrgJdtNwoSdaL7BtUTEToCu8Me0GdO
oSNrTx+3b5JNEB6WqiDfrS04Ah8Yg9zi8mELrRJscZFHvg2GhT532bCyzLuG0dFfwhrEL+kxklgL
40c4YrxB5prGAcCRXZklfnG7tnNeuXGHZEZpPgU43HakMkUC7dtl8KWBDv4TwR9fSJDEKvPRrnWZ
RxnO9ZspdET0kU/PM4kW1y5C3hEUmo/jztnU8eGFeJ3Ow22X4uN0040BZ3utLWXBXYw+NRZymWOT
xQkX3DLwIby7/IC0bkeG2CoUgyQc1F9tw9NT3BlRKAZUXzmwjqCquHBZDPT5YFVLh5clZLUtrwJZ
0pjw8w1YzoWyDh8HeLSt8d9GAmpvCSV/8SQQpB9T1fccq9xzYDvPkyF/54CJnPs3uASZ4trE0KOY
huggAix/npuSYEtLAYxk8p7sUrKa+9uULYb1GpWGeTxLiKoMuiUwM6VnKTmqdusGA2GDheFllMsl
o8YasMCv9ABe4lH1DcZFt3G2alo1ixJDqa5KChd4n9dEh5MvKui2cyjQ3JwkC3S4MdQzBlrG7NDp
0nBvYPTUcrm7Zki+Cx6i+hdcWa+Awk+7LUw4TCaE2VXUGuDdlK+MDEZZhvEXeGHVmPKTN9qlhr9r
xfypO7FZ6fGzBa7wzz9xtm/wgV2JpkBgZyizxpwZ+/kCBRea5FjlvBXVSv48KBhajPqSuCmVNzNg
NqpFeQt2a0K+GjR6uxfo67qtVNamuUcjv5RbY7XrjeGZ6aNoeLPKYvHO6CXpajX2XxMYw8d3LNcg
vf2YQewcVRuKwi+piwjDvYMmYRNimUjIiUtqPa3jAjzzXFQyGasN7TH3ko1lgHZuqlrDaqFOZc4y
6eIRTB+W630itVXv0AcNaIczGdfP6rQalTiqHYBve/YdcqjMH5QbqNjjvSih6d1+UwFl2t4MOU3G
vDvME7wQAWb6C1oyinkNYasxrfw7ewmnbq/qK7demym6jGaobTnkQ4hexkWbZMpAja3yGmLjNA4E
//SKRC/5ZezrPpd0Av+fgDj1QGewWEnYLVhDSYbK94otCYJLwEKL0GUkQ783cPxqPpQ0/RyWYCc8
dZw8Pv2lahF03QybVPYmw+iPvsNgryLQPpYiBzXqrFfXxsYiAKLN09WUoeKdc7K0dPpO5fIlJmJd
14qw71ECjPSHkXs4Wqx2kSGZqKr1plrjKVPoHQ9fAHjKDMTdBy/cM5waWvnqhGjRPK7a9EXQWtE2
/f4g+4dXUtgn9B9v65bMEzvDZFtzWHGlHCZk/ZK1poiu7JG0PSaOUVQ+Hr6rxFMPq0NRvn6le9yx
LKMQ9yu3pbVZH6SBa+/cI5ei9jBhfm6XO8cEvG7Ht3EPcAUJWrEIqn7k4JYJMZj7HnYQsWLwHsBK
DRfNf9nei2IRLmTXUUW2uiKObCMaDceCKPsz4NwK0WtpEnjUi2dpOb7A9tO2fD+E7w1t+LoVufh1
5WYsnAWjCOos3hiQDquIxVja3zAUkOLBjAqWdsQw0NxAFi/F2zL9+me9bg8Rf29PnmKn3gY1wIUc
PqxFMoXL4uehtxmQZ6+FVjq0KeDbrpVH9PEoyemQxejaI/LprwnUBaDnmomQiL968narN1Jt34HZ
+WSraGidE5lI/zVAl1hHPZ/DO8DeFfSNXFi264pE8ZD6Cxvvqds4yig7B6M17A4aW0K7vahiUxQ2
Jh2Prh3v19pjbx2zUBYJq1AmwWF1spBT9dAcB3JFm3m8otECR6UjgcKdoi+oeZ1KFzXXno+xqMEk
m0GhXT7k4dc+ExpGuvNTQXsK67NdlnODSQ6VgSX7ka9ZuGOBuuOmoJtDHSOaGN64XNHhIXZbZRBl
SDZuxH9acxO2bAvoaw0d3O8SfoqtyEkczSOtO7l1Md1EHq5tMyEsuX+k//N2XPRdE+QW+XiBSNz1
U3vV+CcvRj8h/xwTCnUVQGO0Bu1eyWa8KLf/jxBjBvzzqS7P8Yzj41eKSHDT7np+unI2R2tk7wHx
anhrOBvPitbC+IGq59f311eaxoLh0Nc9u26R5ggi4O5QyPdS7iI34my7EZ7lAG4FY8d4HKmVR3+V
dvh70YscFd0vWk9QWtv1BlLQ5V9Y58AsGPIBgTYXh1ffDQ/fHO4ZgmSe2uMDVGxoMCpykEugH5Fw
BjHBUTvEDopWejzXsTFRENy2yfcE9TWmvxUcJOV4Sak3WZMCqgD/n1Kh9HelrBiJS/kNM+ZZ9fg1
5ioZnhRp1U6e40te7iFtCvQMj6Du+1IpMOJ9RCBJbkP7KsLjiIj1XNdN/JeN9ThHcUz99xSOXVnz
/OSS5bhtiDyULKLVKDYzDh1xJfhF4ykVShugedfXzx7/k6bO11n4u6xyL9lTczM+h6Ilx8ThG1KD
CdVV62wkbgLIDTMIRL3sA747LejhYWm6amHTtSjgkgKqEVfXmtuf/Si8y2QfpWI+yZ/wNduKmEbZ
mihqu6c6XUIkDFrCto7++NrTJzGQnaYkH4qw7otpQzHzErfHU5mGb0PI1/hXXh8iZjWwWmyB7vj+
UIa4V4Nu7BErn88ldf5XaPaZVuZDU3Hrju/uIfVj2Kq9Lvhn2LWY6+tJPttJAwyMCAbfbm5V/N9q
MD9JxwLOQiTmt8waU6Ja56uRgipTQksts+PaXbUpH9xPfCeBhlUaUnz4iThrjWLu4m6k+HUXFABo
bhwpejTPVnuSKARE5pMRInL5EsI/J1SB1aXfB9x3rCHMV4NSUxZtKIpypCyaOQQmUfiopt390kwQ
tdUZp3XjOd5rCz1qvObImBsnoelKHTQHAzUcXTYwzH+U0286XgLGabUOuXdmYKAblZGrU14nnKtK
hEbLs9eot+/6dWHVCdHGm08gdPnowTtzVg7/F8qKUW+exsm3UVVncNCc9H7ChbVzchAcqUB6vQpZ
zDzEv8gVSvkpkomXsBhELq1wLb6DhSs3WefP+h7zPr7NHW+apNvUWYFgfbCRidePKLDM1SCme5Vf
TgpmOTFmjPHJSRmdBuWWJJBsiLAZXTxKqtJV1Yf2oqEQwCkbLa/6FohPhq26Rvj0pM9kHQTf2Spi
ziDqMB8mTli2Z7O+tYjCbeXqyXlLjL4/g46Kv7dqycqNHf+v4rIMjyR8pngDMHS78t/xwbSXXUv4
dmXPZmO4KvAfr9OqNHjR6p9soSfhYxh3TyknDXTWCHP/xUhNcH60nlzg4eVCHQ1YNAlMLhHBOTAa
XKF3IWWQ6KwO1/cbv2G/HSKhhGmIgHBDqG6jRYLtg3V0X+V+m63bw2nE3Vlnp7bCpYHITUTVIh6V
qI67OXC1x+kMsb/S9vkY8fbEGY0vVm+U7yIoZiYtbJjzVigkJiiCRZb73aut1xtmANycTFsgkgfa
Q8kDB7dSO9QRd36Q0aVwNO9HA8sQ9OnsWSJ59Hvdezx09fKp/WPwtP5pafaZrcAttDQ3Qga4wbK8
4P1/y9T2ifJfRH9Q8cwBrC3HkSAYZGd4/oGuWpwwMbXl2YXT9ww5Erm0iB27xZ6XeI6vMnjwBU/n
5SmG5VC3T5u3ZeYxxmuJLAaG/WCsKg9J/uanVconf+D+RLHcJhYvsGefE5RlQeus1Mz59jqUNkll
gDYOWTK1tRPhfymC/8+xdZ91Lzkw70DeODT2Dz+1Ew9nbtWC0UrGcJCNKwKrZmcaFw/gU5TwA3Rp
fq3GlH+GRlTtz0afpkpqgAdZAIe+GQaskXIWioc1fSjGcvmatUSRdLJFjVezHaTZO2vsc6cJU/Lv
LnMTFsOBhdLv/XZg8jw5K86a3x0jZwc5OXH88QHXuFqfYLDuTyA8mmo07wLYBfx9IPMTU4uAk3IO
zKMM9F1nQH5e5FDLx1luQuiUn6ntnQFqY3wXq/zOomelZqB6gpzOKwg3pHfSpq/WhcP/KvLnxU7J
MkBiNQhz9UbLSIomdGSAITfquh44ou8xqf40GAToFo20+cQAtDvHIY2/0znR12fmRYZ63iAdz63V
8zQQiFiobpwQ/l0zOIE8j7DPelP9z2wmLdBg/tEc7dN1CrVon/dRgFfD8JGIE0A5Gl8CXFj+mvSN
8XPY0n3zyw6iB/AZsant3AsssgFZy2DUdpFZK8JrxFvu2evq2cjNou2cfRMEdurh0VIQ3IqSzBAQ
PrsGOjzOXaU+FcdwqIHXltTMH+9Nu/NpaJdC0OMqaNLU+xlqj8n+tv69p1MAEYyiwhbMFD8ls+Y7
OUnVIixx/8iJ3WvGgewYZtFblTKDAu6rhjHP9b8raljGDJTBoV+lu7jSXMyuUYNkfOV6kr1nLEDa
zz5KPkn9YymK7w3vjPxVTvjNp3XP++dvpDKZp3n85rKoh1c9czPYN/PHua/o/44KENI1PG1H2bn+
R6nS8ZSBXv2oLm3EPeFFvbMN6kD37NJ1hJchv07NjqTWjLwfD41AMSfxfkJVitAbstaNQuiG8osF
GZ+lhYVVrR95CD7Q1CsnMYWtlC+cmrGQhMWXA5/uvofTPyJd8I5HOYinc6dm/PT6mZ4C9Kl2B3Q3
HQw9Os0p/NEcMFhcJN70lJWe0KvWJTaiF8oxeiiEc0Nl0oJR4tCy/oDxrpjh/Hm2IAFHsXaq/JvO
TIQ8DE0sWGYL1ir9/NBQN8SgCMdq62tSKP6j0DshQAI0yB20rFv9YJWT3I8iJZ/7ethZEJZw4Q6m
CfVyRGdLiAF5v9qodlKK+XTBUNZw46EUEB1tt6PTbF0Q/UTNY2vN8pVjX+0HyKC6cdj1C9xPypGg
1NNRa8BLiQ52ia04RmXn4JXeZjZ5juje5HN7aoOpI8TPAE1muMnMS0XABxp7Xp0mU95ATdCwJHxK
5G2uABimhsq2mQ2qNeYCFzGn0m4mjVkwjyQ30xaCGf8S7e3nU4gKbglW2Q54AeAeBRZoMuMGbpOp
hVxvHWsnPW3T59XOJJXxNVOrR6wJqi4LRYBthW2UKDgdTXatb2FKqkCF9lT+5lU7UY5hFdY8Jf7e
ahfGRiHCDqzy3M1k+IdEqfbX4Wmov0U3ExCbY4Mp4YfMwh6tal6lkQL21MKlcrulINEZZh1n2bGs
biELtJIU/3Cv1bApaOKnTWhJpaAv0d+rH/ZLkedX2RyioyJkCZr31L43E1SHcegCqa7lmFp1pBL7
qqdSPGd82mhdD8Kq6XbQDRAnKRxrwFL6Qhiswjg5OJZE2OFvNm5TYK9WDC3qPSu0hABKG4498IR9
ChysPzuoVvetfQs5vTi7S2a4/E/++dp01HZxxHAEND67CKXuPQr+X2G/a4+W7oC64geBuuB1/j6o
JBZdyZ/vfJ/GMJvidPc2RPm/HlOl18uZmlYPfZRG0EJ+x01hytVkKB0yvkiukU3gLbB7jR9Jdr3i
bDi5zrutFi0H4M7DWvKw44jCwlAIc7BnWlIZ89OmYYainlnlg9rMh/JQP9G3NyagBQHfJqbd+dlc
Unx/LTUrK4YKD++bU86Rln1h4Cty5oDlk8/BxdxwCOQ/+L3x3j4/5AgAPi2w98LzlojBMQuP8qzl
ywkGPu6PK4q012qV4eJKrC2EaktQaeAWKUKNnAd2ylKkRjEGvk0tsbyxCqLSCwN1w8S6MwdDHFfa
ytaQQCbBoNRj9L44qv98zuqPR7y8Quk7kVOVOqvGvywWxdUcVVYOAMaDAyFRUvnpqtN2KHyo8ZLN
MzzsU1Chmr5kLVkmly5I2NXR7Zj/6VsOId+ki6WJZBsHrr003Httvkg16OX21xi76fzEZyjhv/Rg
bD9vExU/FDt6Mu38UJPB6evAWwtH6EEW75zFrwPGHHmilm6QbC7Vi5sq5htZlQVcZ/TLv81Pct2l
kwloMvCBJqaofmwr2FJorQFeNHc8YF2pG74g4r43AOGnL46mYw1hcHzjC2UCyDz0SJddowSLaxV6
Eg2cNtl98GoqTXxw7M3RezYvoSimY9xod7sCIvscsqXchBgaQIHHDzo3eF8VW23r1fN1DpvVTVXj
F2QuK61A1Ox6qpiAtVXybA1ZbOwy+qQ0lcnBxhluxxbSbEXK5Ef8PrggdJn2YWtXzFo4qCAnj1wl
hIDLq8Fc5CgcgMaGmDpc7XLX8YuSc3yW5W6cgTfB+xlFS8F3K+ZCqCQI99cXobh9URfsA0KjbFNt
vefslfDSt5MHG9I/+vl6Um9ClNEQzb9VCrtPpI7XNBVnmQUBPsK4T9hwoEALnZACsPotxhmCxsRz
it+O8RWQQgFdChlUI4aLYrpXgmD7ffCcvhum+uHeF56O51uzLnJS9gnxpLZqJxm0GI16TGzIw7aR
laPFmVO0xyN6YoL/9AVmcv2BISzXDkvexG8zLgMFZbzW3sMwNsIBww62MFMarxQXXMEy4PiZqj9F
GR+iG3UWh/UcNcohu3n56oj8nkNVbOJxNkkCTR0euQsjzb5AQNo7qbnY56Z1lV5bGOkQ3qLfOLoW
Jqi39AlIOMx8i8zqkHvb+uefdhvwv7FI8HK4qmOquTPwvRCwRoPihvCdmWCq3pOQh9d11OAhdtBr
5VCKBymrtz/zlzZEVSTCtPSwQRiKXjHV2ZTce5UTIx86zazUoi6Lii5W9DI2m9ZLdNfcz8yufwxA
CObG7HWs8OcEbnRQORs1qi9x7Tl8nZoL1NWwN3ojw80vU62rf+d3PJ1qpPuErD10ZmFeWwUoDjCO
uMR3sb/mmr2wX/1pA34XhSfmg1Inpgilzw0UETxNFGzIyZNOKcrL2msLCZBUibVc5Yn26B6C1cDo
jKpbVpTFq7dnV3ak+rtq34GgR2aOQOxSxm6UV3+r5m77MN+VEi/Psuy2DB73YntEWtCgP0RYdWsD
M3zzaYK6nXo7AMUGqVL+6qn7Cr49EPXExCIbb31697/E+BNkKAv1qoMLRUgjpGJjH53tGnnnobsh
hN9//rPXfh8A7R8SGYxojszrYpStDRuy5AnjdEcRbVjZKADPk0sf/NsacfTKpXAx26qwCH9hqOAv
eeCUqpNOgXyOICMCSg4z4wJyQ+9j9S9oPUCl8EMwpUbNWw0/5RlhjydtlKAzVi/9qj0Iipuuyf/t
ibxbiBmmN7ufwSaU4DazEi1FOUFga4AClYGy9vqYRDyIzZWLLtswSm4wPAk6I6mFvjr9ZI2Qfz6Z
mUijz8cCFYb/bodaFlYqxEfwcRjpwcJmOoGYZivA4BAdECzDgz/Gazg/rwgUPr0JMfNMF8r84pD/
uEk/aGLfjjG6yRfvtbZ9sy9cxLnIEybJWMz4KBDWVQ8ZZzKhooh/BLBzktBjDX61N7dfEtx8Fj0k
2Q9AfPXrRjeVZPJuj2Xi+XTkAwehSaCVuRvDhv7gf8iGFx4yWzpT0yewPwzFT4SovEOUHTCJXLsb
sYgzi3WKcNYS7Zi+FIFejKx2mRbMq7xOsJboJ6V3UDLVvp7b38kWnAZP761Mx3W8kZL8dfyoHRli
VzfNlDAkN8H1qXYkJ0JBKajB526fI/J+P+e1IrN5FPsJvGrA6OXxqFJQXFsgl4sPKV2xlhrLkVBv
keKK10m2e+cKO+EOUbSgmTvgRliQ33zX40ZR0y3WltDPVcOlXjPAzHw1TsXmItr31XzdEQmQPO2v
RMUeROpYQw/wcOsqjj9gVwTc8Iu6Rac/9yZyRW9PQMqonmBGUTtiClPR3yhS+OhbnmCoj6cztMzL
VOb26p+t+56ZcF6OIUKiPzNYaYJBztQmEJPJUwQogVeVfhif42UefjsHewoEIoIzD02iwQS09gW8
CX9Ms1vL7i2pop8mZbA2Dv27z4AWcNU4+r6rwQPM+jv3m970YwgCXyThM9uCK2RE9nYnLiFcnllu
RSmtBWW4muVLPGMu1H3M0rrWPWEXRqUE8Zfo5nySaJPz3HxPO3UMuPL7Dven76V+cwtJDzioyW9b
T7W7BMl1BtF9V08O1jXPOUouiqXL80Uw/A7RmsjLJndjT7o04fEPbJwZwPFpKWpqwioEmheZb0tc
yWgACypxPG+oG5YTIjvXCaGvXEw1bn++hUc7wzizeqBqhLwnMITzOd6q5jFOGq8GzkL9e+Z/JM09
rjXilVHSo6iUqg8BcJLcYruSNGzwwrymmSoIl4iQuNDCfo10aRzMYCFiJvdmoFqHOC4IPcfkejAC
+l699Kh83GxBdWAC6wuuFcHStdk3s7OIWxK7PWZEX8o3SGpJq9LaK/ghqY9wMmarOEuyC0XY3rQ9
2f/qYPqQFn+rCJ2+Ya+EGTlQJooyJ4LOoBSk9zh17S3j8bF/bsjUPjij+/bAcwdYv2kkrHWVOuFH
dto1zRbGLi3lcLEY2GDXB29C3b0sh9A7qbj0L8xZpM6yRrEHidihkUFLixt61BskslHVvJHOzzx2
vJ0cC0xTRvbspMZui18GP3Y6QCM9P7+bCfim54MgyJ2oyEBvJuPxo/9AJ5VF8iT0slEQyFWm2NeL
Dt/qn17v/9NMgSC6BRf2HBfAWeAOVdmUPHTQj+p2cud4zcV7VbMdCK9MX9UsL6+4cl/zzPkoAb4q
fI1Vm1byDxBTPPbkj7yMjnHDEjHYvZfu4QdOcdZEbwI/m2sHCJQOBMzgdF5JcZrlP6bdS1QehR6T
VofW7yuY/PYi6pGQfPdZyEatDXRPh8CK85LuJ7Yhbc7FGHcvJfl00REXHSSM0kBV5LXpu5yvVnrn
baTWPObpK2IL+Rkp5uNLWyc34cFtQFttMTHWN9L0/N1pP4q0lf1U2FI0PqDAbhJJSg+oT6X/qkaE
2zOLly2fKKr7GzBMq48CfPnuqifrfDvpsxKlNYXBlgptjmSDnP9UCOXFKs/7wMqV7Ite1+Pr+bmJ
6RxoeaAaVh3ZObqQsFTi5WC84oVoGQprVUy90lcKyV5yRm2dVyX+RvGVRHIp8rDRsFZuSp0X1v2C
wCKfgyxzo9taj+rhhuoDEpKicccKkrYLiDscTgKaeoX65rbeufMycmknTeeg8knMbxkxhM3NH3pk
yfPtKl1DfJa+yAcKdNJqWh06DCNHUwAfC3JxempGYsqSCFpKKw4E/MsETnRTOpDq/kHp00TIhkaL
kh067mgjv4E9nMZ32we6WCCJTzWGxX0XxVCVB0OwoRRZBmezhmFaXDx5gco5dwUZxD6lU2RkqHmx
SEkts6oN8ZJcAvMqGuDA6hx7+4smxmILONBPOW20XOjzpPEoJhXvpQ40x7O52mISKsGAYBGsqvMW
IoAUReKLhM4iBxpAmv+TzcmDcN++wsI8Orwlf1g+TyOGTgD+yUTW93BD5srE8ED/4EUjKrUvQGUu
02zHpSi/Gy8tCDOvM4DllgHDdx90/4EBsDzjZmp+sfLVkaKGOZxHhSZvnNprL23FRPzj4RhLptvg
PbIH4S+Eubr9qcXgbKosgDZJaeujFPMyLG51vcbI0nFFAhLuGAJZRcT2pQ0x8zSaRit6wQ6cq783
pMenL40NMw1z5wgGDtmbOQKv7mMcYXI1d+akl6Tr3lcMtgZIX8YspcJrJIEH1ezpSvN2PWA5GWws
LT05iIJ6JnsDRQy+ungbdwLQ2VcCn9SCqoz8EJo5t50veWLSwlnbzjEnXgeN5HxfZnkvR9CCdrXn
86nErnlvxfXg3knBSVlPPkVtA9Qh0qqNFapmFtvQAeVMFJIgVGAmrKU2F/zaPj5w7NO2sGkZbRQm
pOe8QbmySipCX0a+QK8WvNFpJk5XEAvKGRo/TQXCb1miPr6qARaFF4MzRKPl8FGG8D/tqTV6x4HQ
2OFzMxZ/M8VnkIPX2XsizEdFBdXWSoz6QezBgpVNTmBO5nTwIkblHG4h5bZNenyaakMGCp/TWEDq
l/9Nnx7yFoAyEdaR9sJHpaYH0+wo7BXaIMlJz7VOUXAI+MDORx73wb7YyQexNRPW7AZIxoKJEahQ
3vM2BH6vaciZTCAIVq1mXKgUYOCZc4tysk0Bx9zMKGVVCNhLlW5x1mU2gyIUyCpHgKoDMK0ogrJb
rhK4C9CpO23hiYbeoYksyR+w5wYVF24SpT6tEeB+avFCOabU1WhVmMtaVTZzYMeTFAZHrqZbiiNk
wAbFgaNcGiU0i9PJDmeKzoIOqfUgMrtcQIeSU8yhLPbd6WS9fsQqrVmMXtYtkJAFcAMf/L7pkpqj
phv2bluoLNJBe6eJbyS7hfrlaGJkU83pqr1apUSqciQKUPvBpMa5vtPZKhvfVrz5qSw7aij5nYiS
LwTBBFO2j1P6J1Nbg3ay6TZBzTibow50XBFZHjuyORESbH7rJPx6ic1XZ0numdkK64II78Ivxt/4
FYx3Szrwr9syZ11uHsgvmwR8+21AbT+gUSDfiymkOUIt+LXHV0ADEbMD4nlWue9RD4EILccuoa67
Lh9jIOe1b2qwuK+yN5YsJA4+YcvudO4ekLjsjPPoEEUdyw4CWYZGEXo3FdrWGKuzCFW4qFvyb6O7
AeHElL/aBRIDQgm2yxDIe5TCqx7UynFrzhvuaD/gZ3Rw9Gd5GAidH+6cR2c088dxPvHl7s9n0OzC
ZXrdNhGSnuyTZ/vmVAwOD37M7bcTnYt0I1L/XftaldVdd5INK1lAAqPIH9x2eYBTn9lSRueEMQwp
4WpGkLm5iU9dS/aH6AnhQ+SrP2NQJXz+dzNFB/p9qvkTOxW+1qu8uxlLBbN4yIUHx1/TqzOhAJVK
eTiu6XknLzbnoAUoxhHfJZzpNPxR79+4d07c9wW87f/A5cMenYuYuuioryXygyiG/WGo0dL4eG19
gdpn4TIm+5tm6lnVJIcbGLMzgx0C6gSik1+L5bablm2C99d/ZsM7xvIqxKhvmtCFnMY5a02r5FP/
DvjCGuvdCKlpRvKxx3WDYYkMdxFNHDM8YuPcD2GhDSNaTjzbMTkskZWapFF0XALQej+/isKkr2vj
15GOzEc4KICViJJHpnnNj1XBGrmkkTfBROh+spUJ+iQoZdm1yas+ha+znnONZ9lkCszNSsleiyvh
ZQLiIm6nnV9JjpeI885p/5KdY6QyKSI0Oz9Vi608WXqkOgy3or2LggQJfbc/t9KLkktBQwzJgoEA
TypN4wplmEivGKNG/r/ZF2MmeCxkjo5Vn1E81zlhcVgm5fdcajCMm8905uV0ethwglpXPclKNoeo
tHfS6INpW9EHFBJPHQBEgY8VyWeVYP1DQbJkdSP8Nl75eU4Cf6y7tfUUwIc9kS8dsQIEV7J1esKL
vUgpDCOtEZgRTajnwXQlFumJIow+tAQbopekXGfY96koLMkTcDBnUctZ1lfpzfhZqE1pbLy8LN+F
NYrmI1+Xj6FG+kO9S5i+EBFmGhX/UO8ORC8cpkzrl5UblnYnHNpYkjASryA0+Rf6l2oOVRo71uZG
7d19gXGt2ZdW6r33DOQS9HvOlnDQgnLJvGDO4nbxUZts+gRfztC3WeMkZWr+H6pe4618pqj5chCe
/AKwpv6kd9Z6gP6hjt7oXPRODo223qrWrSmvDKZZF0LNUNzb+W1QJR7kJrL4eKcX3DtIH5syCDJe
88/B2A8FNZz5blUQqdW/C4iBoYTOtsCK2zapyX7/R6Fr8G0/s6wK2+AGyREMqLrl1B2RR7lMxAho
+wmj/GMYnUTnd0F1o/PuqAoCeJXi0gmgfWWTYf5Y9sz5DFXvxoaqKYzE+0CphgAvKnE9j6Ppba8x
CMiQ2nl+/+ILv8Qg/zNbULCaa8/FDwkEnM4Z1sdYY+gITeowSZMFwOXEZk+QPXeb96zIqWOGDtoS
Ayls39fwAThTwx8hK5urkquEajRDTBbv7Ps9yQhwjES4UtCdcRU3EgsjTUL4GMEoVtx2GBUUpcy8
2WVFeBBvTKvXLoRzZkIodtDYmi4Y0E5L7BBBmD+XYUbUH94UkVG/ucqwwEpXQtWZSRCKEpaR51Qo
jJjIS7MEV1/apL4Z8B/+3Y8cDvQf7+oTYbcbXbWtOwj7OUEtiUOf6cqpydORgrIiQ2tdJa3pyPEZ
cKn9VbvCkZvVO0Op9r1rGRnInOX5vslPN/Idw4gkFORcYlhNQDMMtJanJUFtuz/VC88auh1yTlLn
mWqdH6wqXp7z1x192CxgABiT1yZSdu5Pv7x+x7FEvOR8PFR9CKNqA/khQ/Rp689XgkN6JLz3ZXdJ
8VBOI+z3A8Vy2BZB13Tdzk7EKvsqc5TKCcr5w1/7xKAB/6II8yBDM16vdwJ0qr1/R+klPq6O8x/Q
2NhzEBhl0BVU0K/rglTE3Dwd/c2aMebvTUnKJ2+pJhEsWms//LzDwVeEZoBAnek9TiamdUSOhnXG
tnzUVrFq/TJsSeLFB1/RWlaj+t+rA15CfQ8yIzxVG8iF+T/z74yqLcqyGeBVjB7UzcJW6FChWzfe
GKlnRhsnXojIRdn5Ac5V6KUGbEHbeWy0LFVd7OP1LZTkJfuqQHuT9crUQnxrVnLtzg6RrGQpsjAJ
JEl9VRvuJimLC+VghaAANEDO+70gXoeoRD2hc4wpFfCEMGyrFMdW/JbLyT4+xNQ2UDPXw6uSR44f
bMJN3vG6RCtr4o0eppL4EcfEZk4wa/s4mGHG68cZ5xQ1gmVMp9CQxFbQrte6rwRmePAS6GsiAKDq
4cdUxZrEzu6TGRozr6gNhAWpJs2E0Z0/ob/wCkKp88KZQEJEWyWi13SbXMll3meMK5VfIg8m8NqW
2TUkMA0hvfIODYX1culVT3N3U5QrrkeAXX5DHCcDSS+z2EHWgVJG5Rv1L+r6Mb1BwmkUkDA5lDHO
ZrDL3st/eHbOZroKr3A+vPb4//Uvdkbt/dHQb14Ag70eXv4bR3WkwJa/JsLEqsgb20o03HIl2QfL
KNBg2nXBmPBDuKizrwYsWodZ6RvdSwAGaAwL2yCvbWOvmHPE8HEEE5C1Byy1A0KrIPVxYYoX5G02
tYzVH27ff4qrno6fwy4GEs6PuYysgqREOQp9+q8YI3Oa2VHMhuLe8UwqSm+EiguEibosSp5CyO1c
o5/TW6oYzlY9rifmSxDvp2yaKAak2gTIrH+R/a3sNhnDmoNFTgr7eQsu+xrW2ah9eO8t7gbA/oeo
me7u/aTX9MJkC7B+3Q5Os8qIFEnEtbj9vmRUS+jw07twYw8hXS6v684I64VxzXwPzJjSYjlX4tU7
uAg4Bv5q6ZgAlxAszyBFtevOBwYnWsqV6QIxH81GvziVT0sD0wtlyMNJ617Z3Pm93soCqtM/Sy6c
8ZsCSAZvLxhGUGz7U3zG6QasfV3J3nRM48W6bS1LvoF7cMMoJOP46CK5cDLH36WeIHY7MirjqDGB
o035Rcdb3WqWVs8beiE6ukCmJj36L9t9eZg0VTNw170YcyVPXi7RMPw/MO0/L3wOqeiupjxlxIFW
cf3zV/Pwvzp/4whFlj/TMzzyubm0zilZ96RPxQPrSEaYvDTHBx9aQbBJ+OLUITFRWEHAqIFROTrB
HH3Tp3zuWut1629buIuZWZ/KDX9amalCOJwXZdY0OQ0218uwpQFHnVUTY8ffI7cwKFFkg56tBumR
OMjbAO0vGPdd+6DQ59OR4KptPx/Alr82pq3NbAmKNinkOmTFoRYraYMIhW6435V8DEb6naSCxdMt
ZTbpi8ikh7LDaYKqj30232yh7bn4wUA6RGO4b+IFXRbNrBQ5bwB7KpTwTUyxszHX3KMcjMcEGB/f
RdGNVdY4rwLfrMrNabMM9Ax7Gde956AeWcOxYkjEFBblhRnA0sDaAGNR4f9hgGHGsaVJZwfK2T1K
hG1YZqstLQJ9OYPfoXc9QT2GLMJq+Eb+iJPVlQGPqzo9X5CvsuuXaTPkdK3mi6W6v7fqKz1Elxmv
21UwCtQSHaN6D7AmM30UeXRymclffL/4x43A9N0bbB/xsVExAecTnYyFOH0B630jYysGc/R9mAsZ
eVkH9feQJyYAdir9RW30XNfSw2M67Cr82l2p+ToVY/Z8uUdDVZ4H0lH/MsMRBltTsrP0sAwpcYYg
1YNZN1EY0YN+FpJBYa5ohP5gDYeKlMF6KNzBpbxLB1+fDGw8H8lqh93VDcjh4KN7Pbe1jfhVM7++
6pN69vC2RSFHw87opQh250MNGokNrXaoI1lM4o09huf2vAD5n5z5c7F/QE6u3BekWNCDDIKi9r72
SztfNOFAp3HHdEEBOFMDL05O3BmKt9iQ/NvfMr1KACoNgP/hUBtM0i7rtQZ4JCXjdfZeNu2lgCgK
zNISFfQoN4ZEJ7cijsV9rT/PivgZSsDMmnF7WE0akhtfMseTg1d8D58rpkqT31GIdhpxQ3KCEKs4
Zp70IUQCD1Up/cw4dY7PjdO0FqzZoYZEfFBbrgUPL0bvc9uCBBLcRARlAs0VTgtgL0aCZrOO/wad
8eissPxy/TQaX9lFR5pY99I+TcY2xSXgF5EcrnPMrZ7NRMePTLVbLWxDC3xPRNPd7/GJfMNt9qav
D/GftIqUfcDQLFWWnoRM8lwnE2I5r6aLCzAUbqdQN87LnNDAPKhYE60cAXizYWMgJGtcTWBmmIhQ
luib9znhLe3S7jVV0szHvFuKMs/cHE83Yj0o9EzzCVWMoKzo89+g02U5Nmjx74ymske0msRDRUaj
L8mTEFstVXKb9kt7oVv1Ca8QSpOSX6qzl/aQrdRYKV0zgviqhFA4lyG9+Mu7geWF4SxtS1bqk2e+
0d99tXMJSVIa8AY6ubhA7ZtkYrjiuwt2t3dW+ODfp/aQqfGuff6w3OffxB7eF4yyRXHKaInPNbiS
fzcqhJQ/tkoS1cu7oclvJKr4gbs3TrAtnW26hNN+cVit3dkbys5j8J4IgPjWGaD2+bZtGSnmV29o
Wh139GSFDa82PB6RMhAwATvKYvD4jlB3cVy+N2fq2PnQ6m6efgy3vFK0yfJ3OoIrEuzz6k77IzG5
CCJjID/NUujL22Qq89VkC4Q6n7SV9HvzniPaftcKuaPUZzJwKYvxM5Xva6bo14DcY6kU63dBOdwD
vh0yVUxtD+7CQTBXlyHN/0cST/mcBAe32FJ7wAzsSRispQGuumRJ9JbWgzUAZlTfKzqC7nWR2Q41
VnhKSOu7vEsS4yoGNi6H8PAWS41mMRko+xKntSR9qQYtTrsgZtejFYuhawy2EjwaIoWjb00LFQF2
kg21znY1IOsqrlvPpGDbWn9DLiaNAWpC2KIc0nlSA/YqzqpS89quMf8tXXJKymmfLfdON4pXbqWT
o56n/xZ5LqQpp3pYUuuKSvYWrXoNirqpvhJcJBUMvMbYMLoq1p1OSYgEV+wy8QALbEC27X3BwSFz
sv//jjDWb1m467P0JYOHv4aV+XVuJ+iVUo0+5LHxoRlES8UN2gvLqp5xGhMRoxEg9O82R6Z5DywD
Hxig72DzvXoZ3Dv4NHE5VysA6sF1Ell4VFJxx6vTkhM0lTh8XovMh+o+lawVta/JHWqhRYRQ1DVy
zfh8qmi0GB0bNJxROkQqujzdpthDWn+CtcdWbkiE3vN31w/o19hgj0hKM/i1LTfyG0OGMNqQKk73
MUy4MVdGlf3STfj8q7c0nGwK+a/BGrP06bKfoCNFyuX5G6aWdzDDHaB3nv80IzI73kuVbD5vaSKf
nNdc2A8ovVXtGg+3/7Ek5y6GTy1ov+zhUVjvDMcSSHSyTqp+0QyMMjp109P5keLR0Vf8Ts/KCybv
PgtWMoGnq1APWUIBjs0AHJmJlEs33fsLnerNk/PaSefIEbZtyAwlXNHib3YS+BwdWSpp5fwy0qZS
ik2jGuICHzTgpNtj8AIUj4GvjHNYwNLHoHAHMHi+c3VjMEo0xa6ogp/BS/4lQ643lvdm3xEaHe0o
ZUTlUKRNCHMBEiDCGNM2Zct3X7XtFo6j45et9OngV9kKsUlhP/FSjTRMib7Vw7akODpWQj3FUlez
Q//tl/JVB1bmxOTiaTHLJmPg8ntmI4zR5iZupaxCTaO10yIlvzZQ2DTpFS53BLSh/ygiyZPL3bz4
Y9m/AV8noiZxql5twkFk+PwijuSM6wW06IW8SxQ3kAjcMtRlsMuWuiW83fqfw0m0HcanZ/QBGXgl
JpXzFYTVLAsRnSyZUm9SfI70m/UXsZRzXzAy+B5PyeRQWrTT5tIru/79PLK0DdWWUv8FSXMSMr/P
dnzXSW/Li02v+mmi8NBRufYzmkGRo5sKhtDMD5wN6yMExkT0HrMW4sE6Dv1jxiy4fmzy9Or0MG8d
LfYRna86q0+FfCjt4nqJ5KkwXHDU8G1IFCA/eVGie+X2nwMnTKK07CNdOGAIBwsFinpVqarnj6fw
O3uf/PxFpT0HxI/m3cgiOwdFb4idYDIzOgx1L4+/cmXfDrkW6q+eJ/AeKoK0uBoPKQWE1YxWu4kg
8i/Dvw1I4iqSXvDfgytzr873veQK09p0UvFJ0hhNyKDjKg2fdW13IW+79lyT+RsrHgiIhOrR+3KW
+QiYFuqx99qFpxi4IuvyjwORbgWPCoNIfV4iNRxpGnhzzoC1ZKl9AJIzjvloRiC2p4tT1BnnvYlr
7/d9YSQK8jsJ12oO4iYJpH1iutXBqfJ6FJVhLrOjLp5SA29ugyexHcbPJGkDAbwEnc31WIOk5jXT
TbGP9WMHHF/aEQYREb52znDTQ0WskUA4VX/P3wv7EvVOr7CmeYE+MzzqIW0rjK9bUOlBao/UthRV
0CXX4zKJxOqSfi7c5+wWSWYor6DOC6bBsm9sWNr2wCz8L4zVHWHvFr3Y8g0Dyh2vxVIsMlpjgPPq
pwyXcwjgIXJGqdPQB+y+Bje5qQ27im7Vzaa3EfPVHWUh01dUnnTxjPIDFOnMKt8Anm9KdIfYUZiD
0CtG+Tsk2yILeheSpe+zvsrkywkNomBhXjFGI3BFz8j7uA/NVYeqX3BbOVmG18ngF0UwqM/gh6Nn
o5DA5Ofts6nuNzkSqypV0I1H8leJnG0itAcaKSOoYrCqQc/QJ2Q8SWyHlsurNJY+/t/fOA1Z6XhT
/p3gfYFesDkPIG0Y3pwHHJVSqN6zzuGNnXUkfxAwoCwi+ZG5ta8ywalxTmYCf4PyXbB5UAgla6tx
tsLs0AWZgK+MgEndJeAkSeXNXGhVrIWl6FP2IpWMKX7pquZYZfUD5udi4Mli9OaecZJLpQfcgTVp
T8TWSVj1f6HPNns32ZEbLuG7bSGH/7bQS+DjPLEKJ3C/DSKgv5OsSxywtsJda86HUspgvlLSTOxi
eg4jLkLB8dBIgsDrkkHXUDXGQakTVVmy144A+bOgSRG0p3PzfaQI2RgpgZp2dy48pnLNkSYEsJ2V
44NHPFjFzKKxCTLL2BiG+5S8jClLViCxjin0ca3TSXi+/DgapqHEa4QMQGcEzp3/UWIvQzdGmRFk
yieWdsUOfHd1/tDJyoUNVBspgbOTcuPWWOjo3NElld6FuecfapQTkWUAi8c99OKmmqqU8ezNw20w
KMbF9NHISrJII9u6h6guIIbvTc1AVRTSP/3sHItPbLwozAwQYea5BVnzqEii9PzwH/FD3gUih0ij
+4G1aUukQnMo7GT6crPKlH1/F2tvHKOtglqkftlf1kgsOT/PEHQZOI83Z7TJhR2zvMCNrvWxfFKx
+i4eINbvxbitItz+5a5vNaErO8L+PT4JGQ+eu0qb7dTDm5LHapEE/eX1iNaRrZrn5z7sI93TNrQJ
0oaPWnNmQVsmO5Tkph9A04jWdKXP76Z1cK0SECsYBvdnXtSxBQP2F0lMhRw+TK8NXHZ9T3hZgXlW
QZSHzeZC2/FaK+yHn5SbCWcXZsZ/mKcACEoVecE/VTxn6+ca5lPWmpAwX0vUs+wGfNbOQbE+Vot/
bpgfPIevSrMnwptSYbERr1VX1ZhtOsWCQsNaD+e7XPC9P+oYF4sbDPEySpah1Y+7RXcJfdB6NE6j
wtqy9M0ioD4dxDHowR7wjH4Xv7UAu3Wzb91Ed7T69IMr7y3AF2yjFHzJTnDv8LmxT8isR3E1YB2f
r+DcF6maaC3hinn4Xf7cRrqB/nmp+OrXrKqTxySBVn8XmPcGQyaLIyEGvP3ob5e4yOkfv8f5hDeN
OhE6efW4f7SuJwhHdG2GG10/BNc0XNG2MiWmITXhGR8DkfcAOG/w8mQeJ8F/bvfAeOfUCmMjb+Nv
wgADU7xWd/HwROwYh3r5JvGcxM2hEieCI51mQeKnW8AB+JPQI6YrTCQ5WDiKqkcxEJN0Xj/74Sv1
1UqzY7/xltAETbFH1XiqVL2lCcJ5YSuTxAQnilMI2hZ92yQLhwHV/3SAQwHLQJQzthE6u04KYI9q
L0nuRHmEqLlBRJJ5EZ7Sgwbva0DcCZJxCSOFQ5cAlmq+As1+tSzryijgEgEs2r25xx/fNCU2rbws
wzjbBwm7uUvr5Jv/9IT0ctm5u8DMRRZvbDRwx/QPs7r8t6VBKt6KpvhwEVRcDHWLo9iDr9bA+kXT
zusc4d+1e7YGX+xKOq7GzPhr42QA0JatDFC3HneAUZkMqf0HCfVJp7Rp716eosk0tb5W2a5eIQJo
abV5KunBQCXYu0qRnesGx5jOHBHeRTJRgYfc5yTNPPHCTqhcTUwAo+/1kr7/2kECJvmhgGybom3t
VXqY4yNCdNtykRlsCOC+vO8nzB1HApDBSpSkYALu2mBv3lzTASi2qd636lBeEjEe88XebzmMz0yk
fLunXf96WLgC+ZHSgUgTOyTLjwcUO/JGRP80OT39yA0qdsHbvHum0mg9OL1ljJ4ZQsyqQcq8Xkvg
tqm4zfymxSqPSHFxt86EV418mJBoa42mUaIAP0hcMK2MF4ccVECFSUGz/jhvC7H33iXiWsjbJSr6
WL17MX8jn4RV/jRE1NMnc2OcsX1+AATP+qpaGFr+wDvJvwCR8oF8aRnfyuOPevNIE77/b1SLaIKn
pv4nTCI9bm/HmK0lz6HfHVmchpuPDRaKQc+kWnO5WrEnAQptXa6IexCRub1SvBymfndjUr5R7evp
IE/VkxsGJC0/JmrcK5Q4gMeoAW97kiJgJnJDsw6Ms2fpQT+h6kh0yDftpML4rTj4v7xD+GKo5T7W
/azp6plFm7QF1ziMUGBYjjEE40dOEI0/jK1Px0NZ7cVwjmmfmTeoVZJG0I1tZZVKcY8LfdBhk/QJ
+brOEfp4h+FJfIZqRLvMBsfJZvcf2PJqOcJ2YFnlBgGTOXUnr4AqzmnLG56A2LThUeJuJ/XqiBsl
HNM2/hHzEgKSci1L8obdDyRGsPlDS+xAFS84YCNluqpx6rrc1cOtwD2GteZoMXYb6trfpSMDjxRh
pPKm9qUvZD3MwtCUw45pjAE+L2BSeE/f6Vb/qaMdPeBa6K/6XYQc7tfX062t57AtfAOkckAAsq6d
PZGTK8V4t1jmwnwpJVSBHT2Lh6GSUI/yS0fpmAQKCpqZfDLMUWcMrCOI09i9R6mBnm9FWqxTkrex
lUM3uVgLi593kfScUNKmavaBUaPvWen2VkEf/gvHdzKguuwj547q80VNzgJKN3iGFohx5NYBUSh0
llj51BA4r34knmn15fdQA+0//2w6fbTmCRlzSNLFf11oE29AFuzdWsi0mwDEHKYrBE7qf+Qc+MFH
391Q8z89TAI9WwvCC5uULm8FOH/D5VkuACrfOF4z2XrxLH3aBHFf5X8oSVzQ/WHh9EHJETxOCawX
fHAo4YivhzETQXQhd4McmCAM0+IcKDWRYcVGke4n2pcdqAy8bDQqZiNLDSauFkIZ8G8FDKxE48Cs
b29Dn9YzSr7znsKdrywlIrjNSBW8zfSnf+zlil7/jOE7kSNIOk1tmIMMB6f5Aw5zN3aT63lv+U47
7S+1FdU2c+70OCQKyTopZ+oZuWQoffvnblDDsmz8gAgwGLvS09PWAToz+uPukItqALryHg2a8cS4
XPHS1eANsa5hEbbFTeAetjkeDFX41HWhilePUU8jU77ZBVU69kcxUpY3pJDV4etPxolGkVH3PhNd
sKzSCRSUU11vCu0bBsAqUiAqt6mbTEc0sq76QDP54h6DZphdTAgPGfEq5Lk3251xLzOrDBO5pTRH
vKTo/Dc+axaLC5YdUbwuJeHcprb2V7teeTlmCRndeZ9Gqp77uDPYGpo6YcdIUosS9oamGNZ7FsYK
REly7GuDqiU/cjCY1bjcSnypp5o+bANylDjywNKawBdqdR3sFwmnWID4fQHS3KLtEimXrSk3/ZPu
usfEoOzZMPIJ6MabUnPuWM44s/bI3hGCUkxBLxQAKdDNH+nnR/2BoZgUuCfM2sfsulGE0BrsRjR9
ebSbPjCnfaRz4BfvdZqJCTOvZlG+mKV5tsm8pJkI0xkATdcNhoJqgQGJogLx/KQkVoqRJHCM3ul5
UYRypu084qUxFwNAGB5JZKsxv0Z6fxsxLGvEFh3fV1qxNGj0aLdjG3e8CMGUxZQnihGBG+CpuENX
hDTiLOiGR+VO+jPPimaJkUqUH/3jzPkV19dnsC/5D93EfHTeuW+ef49yAQbiy1CB9YXXhEZK1v9e
ndv1m8JdhiEHK4uadcNNzS5Owekoa41Fw1px8gzDqfb1DaOK32xk3CMRM9HtEV+Zl9E8IOXk7qq8
BTB1PZl1bdvsTX/3lo//syC53wmhmQFNoS0X5uU+Q4SEUyz2V4g8iue9j/4D6iKVWU2Krea9RSyD
eNpWrTLJeBz6vCk77WMmtEUWI+Cr/TkoUzVRXbiuFn3nJpV9G5jiEeFdu5Q2/y/bZnRP2/DFJXQ4
g1bRnyPkqYumgEKm5MGvEZgC88Hcjvo8ZsTxmIZtzfkM+Pb4MuswCP7c+q8c2w5fmxx5FtsgVPTb
t/QQFpTLQ6dxN5ER10VRzNB3C3eva3ljMNOYPYo3yWlqJ86cKsEc/98dLKlKbxBrxBSbrzB0emmE
Jdq5VawUVgX3mKYvgQRQy3o+Bgy5sTrXefzpyN2qpS/LpGUb1rHIzLq0wtL3fEgD81OL6Ksy+lp4
21+jPVeuQOujV6szT4rh/a+sT3UQqNQzp7zll4/J2wSGRuRi3g/JS7RUx5eyGdXEXql6JFtbDJCA
hKEwRWjc/EIwNIP6wEBIQW/RolMwrEiIXEyP3acYfsfCWcbefD4e9nFIxwBnCFtQuAmJ8sCoqFKP
Hnzwj2bN+wGxRfDsomGHDGf9oDZVNE4yRAFHeFDeAvQQpbS9jEKW4sGcPw2prCCIKqueBM4CBY8W
UUHAyNeU8K3VYU8nF0oj85DbjbvH/CrnyJy+Fh/e14hdvUQ+MqPGSbfKD8mlZqhUBl4RBwFaxg35
Jtrz5m9fmd2vu7PSjRu/wo/Oq9zsJJAtx682r675bYOZQ1+7kHlmAq62cUHJOltb3m8t2oNu63jm
Wfrmhj7/Y+zEzZntAqZq/dHkm8LclMnQ53WBKcwn9nfolk3gNa988A==
`protect end_protected

