

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WOJX5Fv2S0CzprysR8KMEndET58Nnshq5G41sUF8nyr23cEOOYS3xFWHzDNrh0BglAkKcA2/EcsL
0Mi0zP+UFQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gc0ueCwDN9OX/N8ZykP2NxXOhHr0aqi823TAFhXP2T3sZajOBosaRN5Om/T8R3LfwK7+baNKGGz+
UJk1ogy8JwdYWmJV85/JpyrrDFtvClJsQxdfCiEg0IVlJhvJlhs6FCZi5Rj8qwlvbn+/sc8hT0BX
IEC/9Hv+yH9f2HZIeiw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gOAtaUsYvJmoKivS2pd7kBeODY1Q4VX+agLZ2/SaxV/BkQgGuuCLHYg9eGdXBmjxTqXO35IrXGnw
8lzEMm8YS53SBgfLbyNKtLJ5Qej5jTli3Hhz2BXRqoQonahfpMOh6WT/32Mi5HxamPl3+Ad8Dyj3
AbqGosJ8LBJRb65Babsp/E0dGGngj0nJjmmY8NHpqNTG489434uBxC5ykK4ltOheXkVJtXSHoR2s
c+RXEPDO94CZYlHnY9b3pUqLafSVqXTeYuw//0PIJQNmrXYuvkdozgm129vQnlKXVGzYsK5DUlRz
Q+VO09C3aal1Ga70326sWIG6XdhCFEnAfQoucQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3INKfUgfMTydNk3PjPUP24H0r2p1C85cOfDxce4LgEKtine/HDrFDahWRWORtm3mNUVaknW/GXSC
5KErdi7NyQ5+CFdf2MMmaC9h7nGYKW8O4nbf09hLlm3blRBSd2i3h46PihYy7iaS3Q+Z7JKvWuiD
J79EKDKw4Kqn3mmg3iQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YHV/PdEXZA1kC+N7hsk5uDSJPgfJRc2Sgeu6l1dsNtZhWFmXeBe9vCszID1P11I6wOICxCc/uQgT
A2JL79m9I3kuY9Ji47hSGH6+xG4kfTKsYaTVdl+16SjuG/YaIhBwQfN13p/8IGQ6FysnYNYR5siA
+0Lm6CwAYBXVRwsuIA3R9dSPKgq+Sbk3MQCuaqKXbxHiA5oAAI2R3Gz78f9hrvy4Cj5P6dJ+TbkJ
j9bOdpZE4W6tXHasCVI4EqJlfqQQ48uWK076fFPDGpd19w+K6NBgkvxxlXDC1t90ZvbdFgDD30L/
SOFjS0BafCCf2aKaRk8VIdeBs9pr4wj9gMwZYw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12496)
`protect data_block
A4to+QxsJrtUjHWbL/V6yR2+ol8cmczSTJpcdV2LvMCib9XopWzydU/PNTdcmyRtS49QOIfWSzri
58Hg/jXHFQBCc/5eHDn2M0w5VCHvh9diArVhllHffsNR2RWrBqMZ28rA46I6wUP8raW9pGlATB40
Dm/X/GnGj86Q4BSTqzaWmVwSe2d+xE4A5CqwlZL4I7VmN5UX76WB069wKf1lpqJ5bw0slo68ZY9s
r3kDG4VXMPSUouT+fQyKn9dpmUCCjfdSgCwKPby9Lnb/K1BcSgj8H0u7Czy8pgpE86w8BLRB0UKl
uq/UrOselH58oLdWihF8I3V3m6UDvXNYotCivgNhp+BAqYLQEu3NUEePJV80ls3iGYjKx66a1aDa
p2peEUl65JpgapUFEAfQCZe3MQXjAo8PDoofrvfEHR4DULf3sKub6jwT3tlS7Uf3FADfzo3hUs34
SbnQfzXFf5//U9hLKDCTvPhoCbN4+vxmWT+SsfOPTBxe/YP4/kZSfkWsz+yGyVCPL8OLKNrqBR4C
3dvAA+/eqaPRwUYTLyWkrLeuRJAUbqaFtu7agq/h8nP5Dbt5IC2aRLyfHHNrCsv42rjE13NOz/4s
xqfSkLCh6uvZ2wxR9Z2P+ldfvLqs4p42kGazHIwSmeyomZluXStXY7HCmrxx55+MWOWJ9kkJEriP
ROKeXOTVVAmT4AslSxDrmg/J3j5YIEgh4ex9i2IB8l2te9klyAz3F7li6W2PvUleNgMUV/gJTIjY
xdEmuvbypzo6sLf/r9VsamG4s3Obcv4pJeMNpaAXGfOZJiG52x/zenZtGNqqaqRfVkYizb+h8fk6
L3TLdens7K6OXdTeufqZmyETk7xg9yurB63Eq9/FWQlwJ/f9RLZsYhWCvDSEr6oR0Ed3Gao6aySz
nNFmx5Atfqv5s19hld2E4i3IMLbua6tIa6yzJTY7wDyuvY/pnivJCtdXB8uXRLmss2u6VbTbggxV
WXXzq5ZePszqEQVF80W2/oGt8B54t5R99htfzLwQzSqogiI729mPDwfq4OWwe56VSdLzYqAWMOoJ
nT4nX1ZHmua6YYScYn720AKEOjmCMnnz44/7nFZaLAyxj3u6sAPwg4caelzX9LznmtOAEYHKGE8q
hMxyaWvSXCPMMzw4QJGqZmBM8zk2SY2Tfm9ZhTEGLVI+ipy17CRUaUVaO6slC3PbGWclkv65MzFL
XiPc/+O65QR9+eQtRkd5pE1AvnwF+7TwaKRin3vZ0BME50cPqoPA306xg5CGzxOfrGZDJO6FWTCm
4Xh0mVzSdi+D5X5SPSQAFuhjotUCCJGOxphlgSDG+W51W+gdCpEpeLWwOJZxs5gdVkqYaE2rPCkH
c9uOL1LmswYQ2IWxd8XOkn7NfkRZEQ0HeLbbXCAeFbLVSqHjPUc1u7lDNm4CXCiHkIH+/FuU1wex
rawxqmWMCrMhXe+5CQDnIKKVejK6Yx1ulGFf2eIrs8hWbaT2ZYPAcKJfwyFYx03/EPn6uMgrOcRz
YL9wx3ML7lZIvPU7y9Cj/IJ4F5biGkDBPaP/6kPowgtYtTBV5vBFOK8YMb8FkP0zslCXbvCu53l9
fC0JXBT5N5Qg44dj/jHjcKhKmoEoGaADZv5ZD7jH+uLewwztw/MK7O+RVhFNf0SVWN8s3+jnbqPJ
1z6P7tnzExgxQtMN82kkZSHQZrU5sTBS734xeqnropP9dHq0l+bujdKi4kRl/02WF8IM/BX4E0wv
/khW3pQIsWtym8ym7jy+DFeeUFFP84IOLZkMzamDb7lRaEFabCL5uLo++PEk0rgPJGDwbvFYQc9w
iWadsrWn9LGFvqDTPdJsNwbiVYOjAiSX0mHvP8DCsvubn2yPBGQN10AjZsjDhfeLfhkQyMBnXA0P
3sihyMb62QGbAvgYbsKhop40bskHqZJg1IUwoOdZVJD1Tn2r1WGMnTODHW/Ipmo6XckxboBFSigu
5McptFNzwzAK1RVjptd4f8R3rGiu3d0Kvi37NEMx4tHmb85pC2S9mF8HAVT69JPzCXKrexF11iTo
DU3v43qaGQYAZ7HoGXTZAHWU/s2AtMs5lHqyx9iwHpPJ4rhWAo1OXveeV3rGtlJiKhg+tw8sfKv+
+r9If9lQrsmT63NxtA/8GxglHsmOnnKj6jiLW2371GrMgqaORno9xQmwPIdwkBEWAUL/MQXOIpSn
OgsAZnkcWE56r9IaTD7f1xCXyzOqv0+0V4Vme1hpugC59aQAsftKbwTzCBn6dhQ8Qd2+oWSfhS7H
PAqA7sH5YSxPHNG4tlxk7sJ38kHbpqJDIk/Ovi3F08Amcm2mDuTvRP5vw4HCDeIsVAdMv3VJ9UJE
qdp5j0y7xpkEZefLX/jzlCOiFWZ37bg+y1r350JbTJXleFFRgnrkqmCQR5zQXmL32Kun2tk+MxdO
ljk7ns3Yi0o/9Ertb0UrN2NinsXfTiDmQNMzJOmr1ta9eSWLMhrbX24fGtSuZu6FaikYIT+yoDDV
f6Q0iP2EvDybrttRkSLDISbaAYM33nS1n6AdN7NyTjc4uTPgseKB/suONsrLAp8LM/775vOiWIp8
o4tyCYU7bNFcX3lQzlNFDobARkH8qWq3YQVBmS+MvAejYXQcDIEZDEPbObd/aD1hEo1xjBetTTXT
EdX6mYdC8rX35Xj3P2EI+zdg+++Baj5lMTKAnv20VJeGRmBQ89srQ9+0i+dmgEdIz0ofuIjG7Yce
wY3IY5iyWl0acTU7rSX4NBhyiR3qZYyqgD28M4mRBQbvaF7seQd5rHKOwcdfX+nImAbSVF3Wdj4m
imKtu+KisapzTO3gRQYDr3qzLn/14rYmGAX7L4NoXHm/9pLqq3jZGVIJORElf02ZLXA3RNFnH9EN
rJ52PiawLCFMcpl48nB8eXsi/7t4kqzm4Cl3AR+acKKNxWll0PNAlv6vCbN7ea6ozkeYXV65tEEa
3qS2b7lfvRvjXMcQlJHXKGUAR25giSAmx3mu5YDzI4+dov4eU6+ol88o1tOukzU85jAD6iMv7KB0
LzoU590iFRcc+fcr/h2e9/SD50Dt1iJiBedA4cBcY80oWUvJeE9hcmExar+yvP+6Hw/f3DQE6WXv
3bbrvmjb3ciQdeTuAi0qTu8ZMdT5KgHW3Y/boeluYv0A/5mtZP5l6wJse++gN3mXk0RODeDKyjm6
1rSN37VIshDAN/5VMqgsS2uKtXR6n3VFp0vDZDzue7iAaEoiwPDosS1Mt4CyBA3SbxZlC2QSW+ew
VrN/gzKQx2tZ0fkLgT/2x3MhtDNC3z07iOowLHUw8yOuEVXAIlNFevEUaRDuv02Kc5VIldusIXv0
vrv3X8E0b+3qc8IQ/y6RwEEiPbKdGT4LLL1djEcoWTETzXTZdWkwb9CSvtSNYIuE0tpLI92d2PnD
OJleThDIpUDa2bkqI9ooYy9snJ7RDSM7JrNojG0CSbZpwcnP+EEunSB6dDiCct4d6woMm3AF30nR
IcqRJ017GZ+xazadwJTPEsYnis/qO+GnNv6oW52Jew/sNn16/IoL+gv+l/0dnkbZdAd0NsYU4nvY
FGD3DM8YCFo/PTK2QnhqzH71vz25MDer/SVx/QQljlxD0Y+yE8KItjPR0SBc4Ipp4TxxMLB/DSAz
ZmDj4lxDLBin47CN2gVMT1A+dVlpvF3PXvoXsns/PgWQB4hLEPOOeIIVwlPnwdgi+7j7Xdm48DKz
0GBXE/cQcR9+OPmzDFdOPIvlOfmOYlLgbJfhMU6y33QQCfQtEf43R7Vvs8v9M3nenOD9akjowmxv
mygl31slEQ2paIPGfxWUubkCOBLODcGxbXz42CH/zilm7YDPVgHFB8DjipQ8BkIplPM0Qucb0yjc
vtPXMc4juetLryQNM5EfymILXQf28v+fOsL0HDFON8VIXQ1LfaU8lLGShn2wyJ6fczZ053ERephu
5EEw7FYKG8yxlo2B0CZ3XeM1s7mBLHxaBc3vRKlzJfxSSJShxrF/l2+zxpUK8wzQ1A/d6O5eafmK
h6VWTLa9DRIbdxogRoxwZWG+lgoUFmJojtEMr541lQOJbPF4A3tW9EdKJ5WcbWRN1fhxQcOz1S/Q
tEIA56pUpEf/r1dfyrL1qUoEzf8K2wffdnxPUtQuF+BJRCNW6uUwCCZd+Y7lBLhipK3ERU4mtBqb
IxuwJApzeadmYw74FOUrPC36CLQYIWeVn3tBdSgw9bhJWLJYmLUFBM+X10PkV0UGfSVawkxJqInw
tXkTCLhRRqVGo/0HFQrW/wLw5fHcOBJIDUF+tU6DV9UmFEUZyYFDH5tLnlebY8pkfyNiwOMYsEMB
R13vlf8ZPAQTtIaHlrl2049/ZDVw9c1rB/Mlo4RGCIVuCj+gTdI8e8QnTnkq23KFObzni9Ov3lvB
JGihReWTSqdMTPCdomQR49wMMyWsk0wSTW6968z/U0jkaCfHKpLicbnxkct7OvpF1lagvkvRDxa+
osQLBduap+H8x20uvu+Y93DeKyUl+Q+lkm06KYDMXtsBB457pzMnHFkC2Haop57afWyvMixIYmL4
lIgXVH25B1S1vmrNMps8XiDv08Kdv1w9Ptc63m8+G7d/hyO+YMjUV8fpKBp/Eo9bnjSw68nalVUJ
MRz73E4QQCY3sQP/+mr4lUsTmhCCmFGxRC2lNne6A7V29sfM+E5TLDd6rBSeoaFPzL/ISO00wwn5
wby/vKR4KFkdHd+UeQLrMVYf8CZFM/jvxg7rYbP7iFqr7bHYuSIwBN/xPAbqUzqPV4G5wv69WmKB
PV/xEiZxDX92z5dak57F4t8aeZ2YeGOrp+lbEfbpc441kRCczb31NmE6DV9D1kpVB3fbxsRXeaF5
1FrxXCy4/uyoFDdV6WgVKiACSUod9ZOdxFVkb3Gl0TvqhgqvOEth4AKfvoDX3CQHguu6T+tbrs70
h407KUxZxQktl5zOUinB7a219HGfL0Wu5+LEt2FdVoZzj1K7MsiIyuM6/ro6QAomHFnW44BSNDji
qwvtXm8JvpJUZb4nETaTM26WE1FT9ju71ZQzeMvWUfLs/A7PvBeJY6B1zncQVD4bIpPds7nnWR1m
ZYjxSuTNqMIUXLBc+8DDh+8EWQgeMVufMLaoljzn1On6K6Tk2JLf8S7bp9firRB2BJX4daJPiou/
InD2Kt77ib0F4MS0b15JMV7I5aT2hCGu9Y+PAJj1HrLQ1kJUXVfyp5ogSYXGLBlwH2uVkAxZiXji
P8VpU7PJg/bd+wZAHL5TFtDJ9JD+WgQuaTQJV88zGb/Mvgp/n2ZXCNb2VOkSnkf5Q+UoYfemmn9c
WMnCbcCeDUB8Ci3v8SDHdtHa3gJzvRRiZGPc4icPjtbrCZPlkNKE5CHHNxAq/W7J7NFMH9x5GQFu
I8cXrf05AMj6KzN3x5+hR+8ZBJ87E5DkeRbmjvc3QPbnEtAmfrfi2Ic7xVzoQ5Xk0DfXn9ff6G1B
66qD9dghfX8BYoqAkOUcA0Zkk9gpiwirtLXNLFUhqsjno+6WWfBuHbAV5w2gKTDTuH75NwMjB/tm
ye+G4qAZ3ep9qQvTExo/2Ha7wrOHy56OqRifurTBcpWpbZowQOz/a9ZLKFKjRn3A7I1k/addVCAg
H5Uiq60CU+uk5ypPCVpXfxacpdHfeWiaEfUvinMyr+t2LJlTPxyj84YJK0gp0dgUE86Xb6xkbimI
JzqYC7xcd7+lsXgft7v4K1KVTKW500Tq0Fh0IwjWb1kIK8HysVSlATflY4C+1EtWPYAttLPPcZBD
nQc444ahgkK7H3cYcsJa7LRD6Li9tLGl/Gu2DUPdM0ype/D+omjr8w8JZM6evU9Sp6++WvOaPndi
4peaaB6wIU4b0jmHX3xqW0TFWE1qGF05/ecgBET7liVmgPxLsQrgOQ2WCmCz/pm/Y8QntsNzd4Wt
8GYcLAvzLqp6HHUcYwPpKTq52tmRkv8XZW4SSIQ2Flt5c2fnIfKkRoWjQzqbNHPK+FwWr5lJodZZ
JYWohNWFgntQ0E/CTZkeemUzXOdyz37hYqCqCKRl0haJ4004l2UechpJTOaNRrxKHWBDNb5N7HwP
+zk15ME5Jr4yzhsbRMgVSlY1oFyQO6+g7A3+ad/Hyhp73xs/tFgLH2Ku8VqFalx3pikxl+E0JwIv
81G9ZhkoGxFYiYvBkQry0rNaE3dK/jGy3CqUglZTMj/qI8r+8Tx8VnZ+Nfuyw5bObrkesX6D4JJA
kvavdLuiWG22E9jiElPqCH3M9Pvbs5iPPgooklC78EOOK5x88/uNrKqM9uFGVidImoV1pRjhnQCm
8BB8v2FhYAVm8FN8xjtR1UgszTlus5CqpikkYBrHd6RTICeTIoZ2dHpR5zApfcu3RAIoucFGQpnz
AWeU6BzPFR9Zpg0T1a/puQfJvx7g67URLw9FWst6TT+BJMMxydQFQ7J4mW4bbh5NutIdOZnu6sEV
aSfxWd3pCFWPwG8n3TAgYydTe72KsPgw96RUbiH1TH/Ybna+BiPbns3F+6DQ3RjxtAjMObITyhV3
0zaH9lH638/8yMLae9TWIGlYcm4lTCakSKqs+v0GIlAVPZoVMSjbqXxi5o1IK0cAA23enw3hEbGO
0Uk1RTj+uZwQYB8DQcTh5KfLYId8T0gDEWLN1xp9h7K1v8d3BoNCMUIDTDJBq3MsMpDHDMs4QJl3
pRAfT4ciLaTxcbTunltogX3sLDoWHDXuydXm9xV9KBEhpCctoHqJZ2ZYx/VO3IDGWm4MWGfwifNq
hwmp8TO59KqpbFNGw8x13WCHwnPQdx0LQM7K2BU2I2VYpNpnLTpIzXjLMZeKccjSFZcZuDGcnU0D
8zy6ctjMAmmS9gnbL2Exv86cJsVhVy8Ik2YSPUyVqWmQOzRmp61fO4VXJgvzpDpgS77WY986c33W
b0P9poL1ZzcHQsih3ad2o1ka6XKnIRvH+oTVzxvXInpxVu6GgT8ad1XKQ0TlFSNtEAwG4AVGe4Zk
RzuKERIr/HLzGw0t0F+15mSIChYVQVWkUTfmM4NPVKE+148glFC//EL0pqzqKZtGL3fK6D3sPk1u
eP871G7cxthVHd6bYzF/KBHw5PTBxfkKuGFpx52C2XdEI9gyHDLnNisRasDKsgjQsoHq9fmoGbS3
btJVHe+BP1TPDQL697P9k/VLsKwuSTUmd2zLuivSq35V0bcsnhUUYLHUzKJ+ahs2FqDFNaEW1QoD
ddgZZ/ZVLETpOaNcQDBDHRgEz9W1Ex+loMniplyltH9oL/IHeLAQMCYUME3X2pK2Q+5ZmJz5EoJ6
hfBJbaFpfEsnKBPdY8Z7kqg3LIfO7WPUQm6d4iLxHR6h7/b2I5jk99BB+yhc0hTLD3ZFbk4H+lZg
+80w3HEI8OGWlJ0iZ7j1ighdpY3VmKqkVu4ijmXzFfDG0xwa3ZlFomc782Cxx6soDEMaaVqiyW4u
6KjMWJmNfcKD7Xi12P3tftUVPAp9k5xUHLVUIq7vif0YhLEZn8NFpq/HtrfHUz356WhqFNiS+bfs
UJap8+CmV6YP6pD8dCz8CYrANZCgZMgXhTGotHC+p8yvL5oZGLhu1LToZMSn7V7T+z0r4KePGVj4
AMmFnPAS/+8OWNalmIyDyIefyzzvU5KqGP6Q3gJPKnD1kYNRWladd5MkMYYnldyXgTvWV0PC/uzv
j50yJHQxQYYi7EPo03Oj1p9VZcfZT7Ie7vV0aXQ3PGqHxc9HwsyDBaBWqZ9UzcreInG6ThEBdJ9n
ssBm+RiGeoeO4K8T8ueNxJKeaQSDCQF9MyAC85wXedk3gt478aoP5TEZG+B7twiK7r0avbdBpDvV
JqutKmssnV9ToIY146wddwdJFrimxMPo+esAKToDre3b8VGXRUJoFIGm7bL+XUyJjweFK+ivh4wy
bvk46GrsqII0G4VCzfptOu0/1gfZIP3P4kZ7/Fh8mT8rYsR9Lkie6ScSa7oI18KSCMidVOUohRu8
TfnjfoZl8r12alP6ksMjVxMHkGa03UidfACPR4L+KW1NJp/Oeau+jZF6PkfapDI4LpiL0t0lHojp
ilQllXp+lNGzft0uzYuyQU+UnGVwQz0srdzwNbvpi+rDGGuTeV8+Za1AzPm/M6VGfhMK01S/QHkY
dG+nRnUtiD8Pisp7qqnwkq1A4DH8Qol7n9ALFcEDisaXmjYWhRUwYO0zT8RLhQ4G2vtRuoEhFQym
wt+gd/XmlrISgcWMan6PgFp6Ryxqpq/+x7NOXtvenlSWc5kjQkUuth8lM9sbJlXQAz1FqtVuhbTC
DYJDKcjLixRkT2CxZMm5VM6b6sjadzMgm97YZwrUedLIhrZcBKE7NGwVFytVzbeH2QGKUWW4E3Bb
gemfgEwOtS3oJMXKrGeGAymDg3Ynk8Fk+lYUMvDtY3IikKNsyGDfxrxKY04s6HcxnEb8oCqPXva8
9DoP8Dnh5FSLAA6A+UqXBxGLT6QGllV46WOdGXS9Qw4z10U95q0bP6K0FvsDNw1nkQL4Dru5HSXw
mbYHF0a4D02NdoJ0fUUf4GLeYZORRP8/iJEsshxCZa+I0Qqp3lLmIv0qZ1X6nriSprxd99KuL64h
3+Z8cXV0GwGZiaukml3y/R5Usn8LRG67KRxP+BL6FmCZ9EPjX44SzQ1cC5+3yXr9vJeS5Lln2PBT
yme4Umb+0RAti3z+lzpIzWpUIc6eVcJzY3QGAv+911WPgTu8PaFT7vRMUN/M2zgVVfcX5uERNSLd
pEO0l60YYm9cX2K6KmAQnTeGt7foXB27Z/0Vmm7YEtGGjG2bIvAqykFy63Uxje6wileXOUFo3nb5
kDQBXhdhOh5zrHLN4/JRuFKsEzBWOH7YlyWT+edOWXRmDbordtXEpW4FVoJvMKOvCejTYLnTn7p5
2A+1TXm5DiKJsYrVsfHSi6C1twEQPd5DT7mQfqD4FrwfKhWlk7vz1HSNyomqUzhMrhOPGNIbDUbC
MMaKqTTz62shl3EV7Mv3L/2jObtJEJLoqHEkgSqa1ecpM4O1mACpdoJ1UqiRuY4bs061qxsoy2ub
PP4uc9HAxE7/BP7CgDRwiOvcBlAwidkjOU1hQiI7SYBwlx8ZzXxJC/LTQt3ygyzpml/QHJ5YXGc5
G6ScV7EGVNdJ7PrVV+G19E4l8bB1g9GeH4nMmbFkLCl+lQbtnlapAwtcoWAiIaeMWDIK45ukZqTJ
zHAQH3L4Lwyb3tcBwFszM3OErPJvKqDwoiM8Maxh72JH2mXPyMpCZ4+C3nRnf001V5yj/OzpzpAh
uua+pJ49UIOVC4vqZy2K2YRmyi77R4HmdL9MphZOvudCxzN7N9/DHqH7kqW9E3R51WuVucLju2GM
CziO4cgyEGO2QGVa9kuvmck7PLWQLQL9QLNPXK0aoTuVFnmj69Jf6dc0nQgNZ3j6MNAdyR2WQiPM
SqOCoELOCr9mNi06aeffusPpEjyn3zsM2U8R4dbXVe6M4aCcnohB3c+I0sTQv/hXkf+3H+4ArreX
/xOJC3/9e1QGtSMyaemRZZ2IhTM4zqU31ZQ8RG0+ZjyGlMuJi6YW/OcIN8IiSHE5PmMeVuL8KHco
EDdzFKuLyEo2kDwPOSygrOh4NPZAk95xuulJBvOHO1RpLNiDdakmEhJElXBCLoVfrFFhyLCVs9YJ
jLgsVN53Ln3jyo0rW7IWeemagZorrV9Fto0EMoN/kK76r8jq9A63Xb9RcHbboltDL6lVrAEWqw3m
SWIJxL41p56+dPATAsBPNSAgQJfVw281LRZwar65IXY2d7TbThWWnIcpF+gWRWn5oLhnl5nAidh2
I+tOxhxRb1YDyiyUxYMB6w1Z2Ru8a2uAgfpEU2Wcg67gYNT9JHwXei8gSAYq7A4F9MueFxdS073U
OnZb8i3Ud32qGEcKKJxjcVLT5Y+XHhoKzz7BSwvVrrsQGbIRDZ9Cf6cerryKvE4TrxwVmSDPCN3L
u0pXvoPcrGVn+SqoMWdq2D6aAqdkcwkHz3IZNqPTjNccbMccSKursRAsxazQVBNKralwBkMKi9D7
pO/RBAj1tWEsfJ3qtjEPVaXVdd/R5JURfvWhpfAMZdVuEz/JnAK3SW31diHuOOBhP04HY+GZwtrk
91/i+7FjwxHFdZSZBL/7GC9WwN/eo/JZ9q3BaGbEm+Z9CGtcOBujCGocJRWYhnp9LbrbPDB3llqX
OhN1yCHmRIUunJ+HkVP0UZoJFJxkYc8CKIrGrowJBhaPeyde2yEPYB9Dns5FJRbd0tvVilpChfG7
OWk0u1SXA0XYzsg7hn3a95TXk5yamV0cr/ybnDxkrlAuPHRxq5XjqiX5R+MVS7k+5uGXhRP7iZtr
FTE4PJOUzeHRRfSVWJ9mwlZDJmOXhxPlELipMA1fJmsncM+/YZOQCtqtHa5z6qDfFVdu6AHs+J2q
U1L7OKBYMzar8eWfDIp785rU6UAPEYMhy5oSSpRV5g3cjB1ATcvt/XlHGS30bSePX+XAqPheC4BT
iT/fC6dqg1BPX8IH98FLdue+zgB2PbrWlbLcVkuvYv4NekCc2cnpfIiN7+9cdL20oKYyJAwbT2F4
21anzj2Hd0T6oQGW8FQdHAXV9ezpntTYVLl2KmPx6/yZrZpRXI8wx5K82hWaXhBC/1GcgHJyh0aM
MkqTcWTyHhY1dG5FH5ku1cqFVnXRmwXpogXjnU68MsP1rR2fF6qXYeZxSgbRtjsf+YlvNJnRJgOS
iAal34IyOxRAIWyaCrVDAGSz3OV9vbcLKoFtMWXOAtNGcRdZL1Zkl8JTUUBouOyh0GDKjq0FSR9y
FYUvJYZXuM7V6iBKETQ0B6mqjck9no7RzSw4BoLmp5Ml3ggrntQ3o3k9SCmGvYJcgrKg39INEKBm
+wv3Ux4oLUAA6UrUr7yoUV5cL9b6IxMZws3puITT9ZtLrmSGqbDFoJkjSu+emf1uCtJyTk7cNrV4
GUN0vHQcT8NPBcGaNvxtRgLSSdO8NND3XZV45tmWnDsInhAoJ2M2egdm8tiuQD6D6bHcg0ptTntT
9xYxCpiKucmAmGxEiTtinDkTqRFzz+JOcLJoEw/sn/mxCcnuIK4IpJ6lMxw77tRIGZqPSfLDTi6o
aYOGpHf7SJlzxPb3hkoQ3YxBpIWcDtvsZkRBT9dZqQI63soNFBaAVenwBDke7S+IBSJzbOzTJoGY
+s/+HplC3Y9jLvzCeWLk7lmkwmXtjFez7Sn5n6/00PVdCBmy22Qj1Y5qF+fZ5L8TSWPbenbTlVli
OqiymJPoMH4ReMmyMC+mJNzs6C+5nRuG6FIQIkem75J/bWQeXf+wd4B1xJBscCeq9T6FUS6u38Ss
oRmF43wn9dw/EGAAn2LZjCBaS8k/U/dCqlcK+6jd62cGovvK6HpdLp+LszBQXokJkdATh9cVxPSn
5WsEuZWgPaQvZnFxtZuLb0WHPs2U0ncXi1GIVYEaGDKegIATQpE3kElnEDlsXhPGq/6RTSN5yAzg
53Kqr33iapu2/77Cam4CBAx0La2pFGZ0ig8X+KoxaGetwgZvtPG75dixhV2IkeZb0ICwJkTd6FhO
Vf7TK1BJjisZv5ZBrs7WOcRnCKV649laNKzqK+3zEzn+4VyyAyp4lt1x7Xk7y9GuRn7Kr+FN1Pq2
i72stBFg8vwTyTLDj1eDXVgoAoBXOtJa2QeYtVlnylmG3xwmSdvwk7ly0JySJ3RAK55wBSGIhCrD
x69SJNR+DNaeUQo1GPTXqZLbN/tExNuaM6Bmu1WE2y5FC8cMHRRB61629Si0YnxQIkZYonJ8Qt7e
Dg5cJ2p2U+BT0nz0xJhDw5prAa2BuQxUqFxqjmXbbqIhXM5H9uvmcDnCG1UnzpSNujzgL4lzx4VU
+P99/LySn867XyyaOUKdR1aP8oD2T4Iylw8o+LHvz98eIat5aEYmxb1EtkjkzeRT2HKy+OWiwWfB
ZxbGpn9H/EgSiFmkiQOUEbEKoldbdpIHAGggA6p/FzNpiWXJyr7eLG4XYdwfbST7KXfe/srMLCsU
PgG8W8PzZJikWoKh8cOaTKpDMCfzQbWeDDPIvPFHalsuPw4Za40AxwNZ7OTrKDM23DtzfHL4yGk3
vLwhvBSEOjrQlKIaUubJN8qkJQ3Em6MGY4VleqxRymqwbta3tmyyLUPkXVrxESK8APfhS26SXsoy
TWPDQ/M78ytICimfAUhuawlMtDPNWfR+/ru5pmHhkZmBS4h1I6fw/wyIEuSAj0SQkMJwtFv8xZOR
LBUKeRhM3uzDtn9v1wtG2g6sw9IQq9Do78ZKzAY76deAdVXnwEt5bwEiHu2dDv9f73vBmrxFRixx
C8AZpt4LDqFpSabqnwwRB0SR9wmc7MgddpYVmHEKMhajAcic8rA7fQNVzMqtnD0K1j2g8mB7dkME
vIilRqEra9Na7nxHdW0zFc7+DcFOXFxAh9kpEWFKYlSkkuZ5klauKj/QasE2/V6wA0sGsCwu0+nO
AAoNWrlxOBFUZnWEgEAFvlVcfPaO7moi5CyW6YVG3hIDg2KGVWB2jESqiN9CTjnP0bAJtwHMHoDr
o5HGeB+8mLxC7rLOksVDDZ5xebQ74uFEmEcU3Nkq2LRtXjyugqLKS2GxHcKxTbgOfgbZ0OXxS1b9
C/cKGutqpf83jeh6Gcu8itEzgTKy1Qzy+fuqNsvvr4V2MPW9qRh2tUgchuvK1fhfsQqF73MjR7PX
09HmEomdOJNWx20NEozYJ6I6EZcusBdzVF7ywUxbBlYShjPIPimDFKvS+rM6i+NFPt1pQS/mGqL8
xgyNT3B5Wbyw7+t4cgmFrmct977RPEaUcapvm0YoXmXUE8Yes2mdKYNVQyB+li607jLXYGMUotQQ
LmXY/xjy2xLg1Q85n/ma8KrUD9hE+J4xKpj+EC7AXZgj3vdWc5criJ4dAE4uNL0+bE7p5oAr+JEb
wEvtF+3Y5BMokuRzwEvCklU0cpXmeuCAVn9g+Q3G6ACJK7YAJn7tMUxZ6IqldF5Rqz/PM3SrNtDq
+JwP4fK/tKYbn7IGRlR25VvCE7eUclngfyPpbTNq5wQmZRpNRC9x6t3rr5A4uvHbCO9Qti85q087
oeSsyOnBFuIduXY4lFUTuV9qmiqwSihu11rKOV6aC9burP+HzKZEdQhIqzLRH8Baqs4tmVd7lEFN
cVrbhAE0vzBoXy6R23jLycHX4xYU4wNmVXSHNJVfZXWHaJYKxPKM+eoIQHGAKwjqz7UebEk0cAKY
I3b1/dAMLSrqHrNwFLCQsJalMK7rLfZ2UYLnCOJA9e8815jgZwOfRZVi23I6xs2B8KR4mNJnbRDK
fCSDaK5vUPJD9cSBTkeyQyB7JOUv0dnM2zdUx3/B00nvY1GMKzNWUWLisSq1rOFJceCTIw0umG8C
ly7Wr2HwbOfGoki/zA4Cz+nUYSlhUya2lmWhi1gYbJbNWdHXa9bg41zBL2xw1qis4ys5BWwAlkl4
YR7dLHIs4XC91+OPyZcpy7KKg1kEAKyTS7a/RTBwcIxP1hqT3hIfoPOWSs8v39u7AoAJb6sY0z0v
bqE+CeLFZDBRohtdDf8P6TN6urDP9Hjd+uOgaDL58PY50MWPy3UDeTbnmf4OnYhN83bfnG2Rkykf
t/vrPt3VWBzFcDXfYdLKinn6qj63HpZ80wDBPwlxTIWqLlqTPl+fX8/xkQTWahVRD9ebGeWWzYM3
88gGC8xkEfYHnJH4UooE0OnbM4wMPeSmqFjkUOcmB0Cg8uFXpDNboeXYHdFIfIDOSbNQPnXtFD7P
VvA0w4bAowbb1ludeqHC2Skr/sEUJ3Z0D7PTUolYsKp69IT9mAs4VwwsFYxAvA2f7Uknq1mSKRLR
TLd8biIgLj9ewvXzogSTOLtjbheY6/Q52xUoi9oB6Vf9Ud+estN1fgKIGXo/b25j1PHtTehSWp9+
uP/5f61nLX8k7lCYraKsVkWXm/JKGwRxSmEYqHSWV3KyWKgBLu71OsOqa8NFpIcr2K5T3hzsC72p
N7Jwh32wLTEYP2RA4uYWy7Z34LXn48vhZ8Xtx/+cwI/XrJhz2q8y6m211cl3l37XvP1TqIDDQCgY
U96Rt6ixH8KFXrOP+2phJSy+n+I4IgbrOY5Gd6YDvo3UuA14HzP7gmQcY6jH4gfUSkb0oKLUlhtM
6xFyfOjl0aXwF8YvpskjdBLIyUCjtToGxoURbMV0GYCVt5e0ru5Nk6Tj8kamtBd6qkza/h1Zm5aE
AX57HbNZV0XnmS6j0Zi5gs0aPw1vOeOWVZRQaev3gxBusms70e6fjhciKxwLmT3kF5nBtzj+/EY7
/gfGz0Vbl3KluDpZl8rI/yMV1XxJZBN1rnzd+zLOpxDUsXhJJ035g5LmHaonv8oxeb7vGT0vKr/1
oeAupGWmoBFcRc3+bR+zCUX6AqVxOYqrlDTV0shq+dGkll/BDNkA9oOvDBoFlUq4ZHg2rW2Y9iyi
Krm5j1fj3kUZJ7LDEDI1PDFg1LQ7miWq00x0dDW5sd1Y/ZnZTbFW5bpuq0O3XadiO//dtbPmtbmn
1nbP3aTee1ERU23jY1WEdHzgFKS0B/iWbQublSKt+xraww6UNNOf5zzkNqrDw0pSzCqoHiVOfckh
YKvOhlbbto4UqHAu9ct1qFO5StzHqQ+ry1NPFf1AhwRSpGAqvvXjZ/zwsTTkI9GVj/cvr2xDuxH6
953IGd/L1Sm/jjcesZqEj3+eoDvkyvQFiDQUgw3AIbYcuMyVrodER32qw67aS9JB2kaxKhjS/sHW
00wKG6Z+6patLPFhZTn6M764CemaG7kXiE+Q1tT1Cr8GN0jMQZjEMGOPWWQ0130TYrFkPE2zfrwI
mWkbjngQsw4w5pW5YmySvcxtq+DoaeyqbSTfwWYU0fr6+8eyqgK7sLv94ItqetwlrPpBS7eUF50a
mCSLsNHQSnTHG0okOL+Z/Rnc8g/8K190N3vDQuNkiJPj4le3iYImn1znDTDWEyDWB7Zf+BB6kVS7
0ICRlI81ntSO75CqBLacFI3wewGfh0jFfOFKIJSC2g3O6moUtVn+nIB4PqH6HipqOeDnAh6oRCOd
3FkmswcqrIRdJ6hfuP9y6Kognkca8cU2v9x87nla9Xg2PrLfyuDnuxfgZrwr0sGzBI/sslTIDOTo
KeKH6ogRGG5ktE9M+lwQ9uU5kyk9xNywxAgX40UlR4JJd6lNsMQ4jk41E30emwzQ2S+uEs6ATO0w
SaYcNpZ4LLrXR1Bkyp7zxnl7tQgC7ZaY5n1KGKysT5V+M4HJ2gDBWn2UPih/zroujDoxAsTG/CR1
nZSGsud+4/m5joIRMQYpg8chNcAMLh2RTF3qMeVt5TG7UMMUYozI6Mz1uKjygwGMvORj7BsJlUcm
OIRKPN9vau8wCnhBOXs47jVBiaj42D/bLqHKjU/3lYKt3M6b19GCtcFPkX0sDoZ2gGELPKWi/YW5
B6OPEXt+TFmCCB6lNmi1kvVQGKe9ce4tnMqGaR62hhBBEq7vGK4XUAgxpQhoPV/9RD7uy8CK2HJs
IaS3EKGkXrW7UQOYNy0nMBSha8Rn3zhtYt+upuD4p2uP5Nu960nerxGE/VHMqzcYKFTT2GfUu+NQ
YVF4eThpVfqwVoWZ5hMn/sJEZOx60isv0rRz65GszfTJDQW80yn2kjb1Dr9DQDVjjm3KFlNhwkiG
auIdaK+MFaza9320iay/YWjw/GfHA2Ibswbq5vx04wLd38AZhkJIheiU1AOBPkcXoSPqjYgowC2y
pR3rqOWZiN0DMrsXeg6LVS+0wusiQxybO/BKwUWTMpfOdph5/zqFmRDNmaiZ4TVSze1NgXCwS0ci
Tj0F4JcXDGSJaI1Oxv/XV4O41qsuySNcfBQuOu2C5qj/Q1F9u7HThDIM2CQWAmJ0TwCXVb78sWuL
RsHAafcykU5Gm9hGJif+Y83XoPBuuLJhRIeDTTdAcYnzC3w5iN76oVQaywub/CXDW6XKC6wn6UJ3
VkHJgDI1wUE8Ih+FVnKRwtlO4P/hHlY8Z5TuwFYrd53NfsrI3lQUBm+evgn/Sf/Dmovaz4M+Eqes
hHCEtgiKuRQ7iSEcidOeOawm1wiEkbVsMA9v4WQbyQ7pDk+ga16lgMbPIPzWjzpengD8rqV+Nekm
tS4qIW4WXHf95Hq66z9SdEU+3mLrpA8qdEAbNHG59hzgk1e05rqIDcNrdq12HlePvxaJHXftNqOq
O0vVy1ak/dX6G9Zp85sGYRlaEg0qd0bYyV5n1FLK6fGcOTDfj1c4txYEPgqM/5XUp06nzW4xP52z
CYrMEBvAB3/8I3x7LZnGKHvHQq7zDq4tQEm4j6AFIeKRd3/FCHZ3BhR/OmePJFUAss1cPg9xwRFm
uBeJ2UIQO0oyhzwO9fQeORU+uFuGg5sEy1th5GANdS3xra/hZ/FLL4tMdBXUlj7hrcZBabtuQYko
vmzXlx+JPWuwButmcmNZAF86jXkpDQPdzjaKf8ZiUhcBilKUTMLjY3ra+LsMaLOh3t+OROpZNigK
6O6+X73gpGfU8RdrDuPkExhpPCo6/tUIYNfs5xZCioLKU6vvAViPjEpKjl4VCyHHzAWlcJjVc5kE
/sGJ9LGLoD9/HNvtgWyDGsO8bzsNIfQJKYHgwemjTSAhQz+ttk/jzYZ8wMBoVuDsBtv/Dn5s/9qM
xvTevbTywvlnHuPLSw==
`protect end_protected

