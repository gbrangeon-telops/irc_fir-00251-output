

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IkKQ7UnyfG/i0Gz2KESfn5rIa2XG6JjMuNzaLweotYfssoXFPRW5MF9/SJXIBGc5jwrrtn7ZIvXw
ZMKFyJ3FzA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7z8fuAKplZhDCneI9mNA3lof0N+J7iQN1H5R3Mj6yF0lZ6gCWQLLnnmsEoxkSX05NXSzlh4gcEg
7rRfO6LtEEhf+XGNB65vpBYpfhGyoq59NAHhGVo4SvBM+mv7uMxOGdpTeOCZ4JbHV0AkjL28mjov
93MegfTkvdkm8J0Lvdk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xuMQUwo0GDzI3cOEq+tu/2nUcDmn/7fhQTHPWWNseJwSS2v3l/iZo4evCcnhY45ESTueA+ZpjAko
WVoSIubelzbNSlntY2uMGs5oczMZtiztniKkMtgrjy3EW9dfGbHhtmNrOHGIHH4IdMr3kAy4Vh74
ZigAJ9A6+7kI6MsJi8v3mT1ARZHCR6MWsQMcVGsi2drnsGRWoYryCO5xQR7B/cwBGzMymTal23NM
pQKOm5sZ3P6n60ZuBiOsJmbRp0+LVYxKNhFdxlNXd0mwyAZQT/UOuOuVbjlNnKY3+syFmjH1X2jU
BRKqD7PfkYIVMVQ6XvOwQSNLyki/t/1FG9LntQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2lTj0FQ90PRwxkOhP58Pis/0pnBIhVIOGqxXo4lWUDsJI5sRS1Q5L+Q6i9o+BNlX2LRPYus/9Dnq
5ATglZxA4PDv34H6B5xWMxj6PrHSWzf271mNIoMFrjsSBdzp3H4BqkwksoU2N0BujU4mvFktBj6s
VuYwP8rZjGtZ8cTr2i8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WKc7lQN7TOvrS4DJ7NNUxP98rrzfIQuz4DIZ8eAY+GKFx6NuoyinV7kCt4N2qBg8IRnkz00LUdTl
h4FZuBrLJJyfOOGbqIiZNIhgdqVi7fXcxV2ef2SWPHLvr6kIV0N1TmRIBZht7FPZCej+/BNW8QYG
B1Rd/mmsAB7hXx6GfVQ5u7NRsVDyxlcEghLjiM7GAdTaOWl/F6pDM3aRwjjOmid8Gt7xmiYfPT0B
Gzk510O+OqDJRqmdMvwBmv3K/y+M1RxYsLOpwIle5lGrJoXR6zj5dZS3g0EOtylaiuYJczAHSe89
8ncn00hUVfz/5JZCkfgcxZH1LxGTI+Ly2xY+5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8544)
`protect data_block
KVHpMjETfckFhwRwQVddKAx58f/Cuya1g9ARSDcU52RZrfu2uKW7YR+mTyar/nPYRNTkLIKw8MLI
6nIYUv3+BvXiS1ErcwThHJlfN91xDGgXhyY9dZmawzbw3ZWukJVHkTjm++q9FDxfbhXCPDBQ9rA/
spFAQ+905AuOLxDeE3A8Omh3rR3qtIpDZ9FFbJgiSssnzXl65zdSYGyPTN7xbImK5rRDgt1awkB3
9p2kWBbN8DV0D1SkVBxRZE94nxf1cQupFtS+8yFq/zTO9FvDFJcY7C+T4C+baro34cN52XD1vTeE
/WOfZpKFQ95GgFBZV/zgNMXTTJ7uvfICBvUl7Ltu+SzgDJTT6FLwDLuz3jK1FKYuk+dOSp/rNtp1
i3UD1uoTtCsnMfit6OdVqQ39xCxyaP/4yQuaQ7g0d4B2YmTBhbsR38gBnS8qkm/Sz8GRL8eXOoCw
C/Au7+SeAvGSYRkgbBI9yp2Zw/GqL1q7fUX6/AkgYR0w8otNGz1QKMULr3QOWBN/L4l3qNTCPGK1
pcQ0A0Jx+S3qZGV0jnW1C7WP+VagXUC8kbbYZS2hASWpLYjDHbFx4UitBbH+Sh4XfljBAU3R12Yl
XtsYbuhqJU7gLCDM5gyM4vOsf3M/P5KBHRla/lhNJgoXHuRiicXE46jT5GyLphBx+2J5moIRquLA
2wKDL/+EMoQHDtg6orOjF7wAhFZZ/YCaCz3wFOykRXSNNUqO3Feq2wpHzMbJ3SFVTkMTrpFDM3VC
2wiV56Wv+SqIRSgloU/iUDCqGBOAseazlrIySZjF8KkTVBAXTIfGCEqSZHSBBs7ttt/tuh7T/ijM
uAqOCZ7mdV+yGPEIUDJAYmZw13wN9O3/BmUAsjgwUS0uoqmKy1i+gCxZhnWXzlTzvEkkf/Kmgqzx
fbu+3tchMnhIYjujQBXByTQD2YxRbXXWSlW5IH1PZJCnJcoCr9SFH/pCcddXhj0nSl+fIwB+TQx5
9bXsL1LoGb0BvgEEnb2ehxpe/c47vuH1UO6x9KwTsuptNLdnjxCULVvCM+8Y7QUtAFRUh06VNJf2
I6Orbc8Fy9Eq2kyntyoi9dBNJDifHM+jHvRgD6ry3EPkS/vrP4rmTqpexNltZt9jGR7nzL7s754q
401DZh63tDftVmUbj8+oApxZ4YtLkqSjT1owmXw/PJFSVM6DRRUuVihi3eb4+/QeHkZGDNEKdH+A
7yo/wiCFzX2k2y/m6Vfy41D4KVfJna4qP/p3YEMlvfphAP9Tssv9xcsQKk26YQx6dGeYz2YUq4ej
6KnrvpAaW1IHzq8U3RREDn6xbTH8bkDCqTlAgrQQy33MVBVmqD4XmNx74cgIHFUKdzfHNgWCD1LJ
JsHR7U9iOgctTt+XylRVPYDj2dr7IzZYfmbSrbUOAOm7r4rgY+95pdCEDVi+ljXqC3gFg02i+i+X
W6uPuApjqtc/RzX6aqdGrlNxKhH9rkmy18IqqzqpRHWQPfOTU4p1+mUrnGQ/zDjzNyQ4+hRbqLYo
3h1l80Tmc692D75i2AL/vHl+b4VNzLRHldtbbTh5bA/2G7PW212l2q5Suuo3aJlh+/yzSk/+vFad
RTosh3T2RNoxDSim2rDEWEZimCufKkuBpS7HajHT/QGH9gNsRBGTMW4n6D3zwKEl1n4GPbKvQgPZ
754kJ2RwcVyiRYUoYECDA+ZZ8YyAhooZGaQs0LeaNdiKJsKymuDSTdjk8oOzbt4MHEmDy9VW0VNQ
7ggppN7pH+/Ix0AATHXR5nXcOkAZ/9S3aB+CQo6B7F/TwXqa4VsHSj7PpWwDx5Q4R0HXNzXWOQXn
07qqMI7hSgTNCt76rFKF4nQ+bh1vTRoSB14kqM8UuVZt7ZY5tuy39F1A2J/zkr+xxB6v36DLsh+X
szFRbZRBiPxLvu4aR7QaWdqjR7Yy5ab7Go5DZrMI7zY2uqeQIPSSRozjDQGhxQmIR01xKhYYBbwU
b5f9DG55YpIBv7Q0IllWUI93euMnEPtspATXBDjEpZ2OCWHjbrJvQgshTaZjSvdCs+jmmWOG7Bgp
P5lWsY1Vvv54tO+oYoLqyJYzxQrbEujF8JeS1gvPvmC74JkM1xLkCRSr9CKhQsOzywbp1JRPWxkP
Qniboke3I+OiW+uEhQRiOa22k7CF4xOeGB9V3G+A5w/NPaZdEW9k4noF2BsV6bmrwy7ibYFdY/gB
kTPAaymVrqaw/z6P3iuL94hoBOqtsSTy9gH30OICNxbhiCJLb3uz+mDPEYw/abiWI3BK9/eEjC/7
Nux9vMK34pqBx1nHKn00sVWfxlFl6kuaMf66EhaxRZU5qVBf6geCFvAET8NQCp+NLmHBaPM+jn/J
XLYSRsdQQ+skaAfhdCQwcjjBCoH784jYJzzcM1O4+WjwJcmVeygm+ZzpV/BAHOHcBxGSBSLeZjNi
bAX/SpOV7heCEnYUSNzID8v2vlgtI6xgEkqUA7XMEo7QvJq0ybNzOE1BzQ8/kZKDERTEgAJ1wmeD
aUXSJWssPI9s3kRQd+itChCMdN4M489mP0bJjn7+VcmS1xFX2xdha6vB833YDJPIV2gaKBSs0/k2
JQRp4SAesns2j/wWSue1J1/WqJkgW9T9bGJh15H/NW7XHVi/X5YHYR7VvAUNJ4JfN1ac7BSUVfTX
PzAa8MDeYtzBa2/np3y/xRVm3BwkbASIzz7gI3Ve2iSquqczsBzk7HnbTfluIoToIhMx5SdA507z
zgSK7DbYAvnBM19uhcxU2wAuVAYLjXwdWTXnOr5OO25BXOP91CenWMvEWFtLG/cVeeqyWRv+BZav
K4a6U4fd3gxLdNY3DL4v773WuzMmuSRdzoZxB5iJhvJnPL9KZc6MlLUQkigWEn6PeQV2vxkAYbZt
bUZAvZzbt3sU/3bBsOMYPd3QJ8StQt8ONGvWSKUionwrJOmL/F5cE6/lzSYuNxnhMIfuHn8sAQoh
Kvn2wwDKm60339LA3QvoPBPydgNND3qk9WpQxbYR9hDraaWHeDwhiva/sWJ8kDanSgTZBvibZHSa
qbiump9n0RvX0NaF026odG5ygzx0JjCZZqgMA3gkVfP3vLlFXnpiXY/xF6+R0PxNnK1XNrgJHB7F
9lQISaU36JxF326GGy5riptwlTNvmYebj2BFLr54OlpRlQueHUwPaH8PxzfL1ZLUvywjRPY/aIXg
A3eB4mCMwRhXzdbExxSjaeSNwnPInKOq88/kX4ffknDAWAUPnFi5guPKsSKhFr3cvaS5CFoRR2Ws
yagwjjEzFdo7VNL3wpI+ATTqPt6q/IbM3VmprfWywQjEXHn3CAtl0+Tfky5z525wXBbKps2U68EA
4dMvmJYMeYRmgOJlwFwfx+MoW1QZ04pBuYax8KzdKZYOBSfyfwZY4OyBXaQFUxVGrwRj0aMkWI/0
8dMMgGI3CGAHYr2Avg95xOChTiAS/uVZ9HDox5e1K5cvr0B5Hrtc+V00vAbkkdEt+aYjKv0716kD
LRUy7GLsEQupCSUUH2RQVU68SbBiZBsa9LrT2xWnI4nohKMSQHJHs0Ak2PdXABqRW4yYzx/cRJdI
SHk3kkb2zJnIFG/jmyypLI9QyIqMEE5/AQhQHG8irIAEZyy9jQ43IjgcJm54wcn4ygJR+DXebgjE
O9l5im0Xa+h7r5rCER0gm+FTH4jiRcPGgzroGHVxYxlMBsfyTFw/y3zFRHO338D81azCPWpFnBgg
stlwra4yZIf9H4HZ4qKDeBmg/1x9YN+fC7WDpLbWPzaO8v6oPqR1/ji23x7voir8HvvoyClqer8Y
1RpUsYtVBzFbKQ5u6UD/OdFpdKTickff5kYOPV43D9i4De0fgXZwpK2GZHr/qv8c4URPPwMSFWQU
6aRaUciLNfnqSh9LlO/mIJRjlJNnNG+CI4SaMncmItlzCa2BdvlIf9/drBoNKhNI21TtY7XAtFZs
cgDHEjyARJLZUlZHt6t5t0UR+EFmD4W9gEjzRbKHbWpsCBsWKdGzRYUp/Jwg8BCdsdtyZrzf4xEG
vw+UvoqBgBK202LcZORimOgPy3dvubPqAaON4NpgU72AigZwiN00eEU1ScSi7OIlQ8gnZDKpR6TX
SKaPaJAVccs7LC7dblZ2Bun5iCTxqJTqzHQCxc2u6PHC20oc5+U3A7iQO3xO5F5LZ4eVMipfr+T3
1dSOeNK83frDGxafdWZfDrMsvUxw3FemUmvOge+deNk2Fy8o/6RWBU9GrYK02AMj3hBNFrDthMQr
B01/cW7O5j1Iu+QG4IbyhjxGGOLPDPMex7ux8jn+8x/9QUd5abEDQfmzaxDsuqd7axP61pRkxJIu
0Stk57UNuH/TCEP1I4xWrwPuYTpqnoh7UWuAHczMn51Ro58Z863FIZhwxitUXK14UV+jxh5gbh2l
dpi4V2rN07B4YCeMi4W5JqPFYPIFr4qq84ISEhgOExsrYukdge1i77GfdN1UhJ0T0lLSVAZwqAib
ft6PQbxJCQtek0HMgmdYVe92/ITeznh6M31nDpDM4qUVPb0C1MbAGiEI86vk/8bOuj6GrK/4ZPnT
DjK9T93vcxCEf8rjucL0qhhVxC0BKd8sFKYmCgN76B0FHLt3KD3u/QAik1575q8ZABd1s3TMotdX
E3ChBlWVqcoO9hOne6PQ23zEw5MOYVbbjLHCy4xSswtmE4X4e7Shn3PqDxjAw+rnimva9NTSFTi1
dm/AFWvxDJLwGKy1gaAgXhpNQA1P8s+z8zzb8ZP2ckQf55sAuJBMx3HZQqaaplZw/xTZCKv0lRj5
6lGvbX3T9aREa6QuEw0lYIRm+afmQmGNFCVnyWUnAD7uQbeCeiN8cUCb9dq6xUdeyrjB49Vqz4Zq
0XlEnHCi1cYyDRdx2RQADcAWU1NaTaYvzgX6sKMk6NquwqcnPHKSTES13NtpOZWb30drjd4+DAkJ
coclnDV90L9MNoa/oWuR/H7SAaJVSRWCIE7conro1i0WhUsY5nUUgdAeAsMYttyWRaevQORK6Idl
SZfxb2OXqmbULRU7ZwenbFoWC8mwshVH2A2Q0t/DSFkwNDt/6p25zyXf3FWtVST15Q6Zh+BINo9e
fZTM+EZjLBMk6eTJVgIFfVSt/unGht9lNcUpr6J2rrvCcP1OnWCOlt7eSNbmA6EOQeida/QL86o0
O9Q9HrMMM88/hpcmKSj+aW4d/s1bqQ5XeKgCLWhs1nyYe7ONAPHcAzt8WCCLQanBaNuc7EJs/H9o
Zp9Jg4nrCpuxgLIAxsYbPysKBM9CciaO7mSZSqan8LwWJMCFCT3CmTnWG+eHIw+5d5Wgf9AfPFeM
OkYE7S146NRD1libioEgHO3XWZZ/iml941w3fwTCfYJ1Ie53dVH4NacndaYMtYg2k5f33yd9/Ozr
tJcCpDPhtFUtmPlHENsZd7EbPwltZ8J6ELUcAYnQGHhPa2IIq2LVC+o2iOSXBuCnaYYsPKaBI87h
OnMu/H6Gpm5lTud3F3mMQMqa2uQhWzob1aruU7ikw1WRdCo6bmcrxIsY87WK9wjqo2OiDQT/n57e
rvcB6SgYAvxuR9ip3kukD4kxXbmfmAFLjB/AoIjx4rwy/mdQVsVwLtXlb2CQpoko2xwZex+GS20Y
WK8QVNHMf4vLUXuLLZnNO2BOku7PSaw3lod6k8fpDpQ4D1uz7y5x7nexnzg2KSo2zFzhYclGlqEw
8xDXl0A1E9Y5n2jy315UOhbud7Jpf3uxKwobggqMb/a8ZVMyII6mg738pqIMgIC47KyaXo2tYDp5
WEdY2VR6cru8EYMx9cilsURQYs0RZ074Qj2anUFR+5rjVUZU6w2SSWx290j9Q4OOFv/d2Md0RVkX
4Kla2YnKWnFyPKHG5BSSyN2cfcEXyGoLOSy5tp1eZo2iO2gK7iSG0T+oDvG4RAnzyKWo/6NeO5e0
ayWr4ZI2SdaxrW+kinV7AqBhugohG85KE+ljPTA6NM65nMu6BaoD+NbotEgJJY1eqfU/CocMComm
VhfBqw+uiclEwPy3C4K7yeKSwvKtC2W/XL/0KMThXpiB6GRMeGvw9DePXCf+TLSKdXy3I6RM+yK8
1FluEU5JmPP0MzN49/Q4gKpcXL53n8gZSxycj6kF0p3Govp3vQJclABv863V7AFT37lLype6v7ta
zGmhcsjxg0pkVXv0ldzdy+a3SrBQ9d1WMXZSRmL3oxF9fO2BMrm0nvUAH4dr1KQQuhgQqUSISqQ7
+breR02hqO0qDAVwSAedAy2HXhuhAptxVFv0kQ5lLWg8+Vpc7qnp95hlbhDkiAcepuuav9o2mBXB
WpLeAruV1LCr7VS8HNeYGJ3SDPrzqhdDwqUnkvO+vKLKVabkLqyVpeFZUbR98inwYfINofg8KBgE
zSOyLr2VqAK7oCzlNp8Euh57sfac8bRaDcJKrG5VLlzHvlWelKD01muHpy3etWAXK2xLpIbpo9D1
heD1NrVJR71E4A73j0efZnxhViQU6HcgXcjvImE3gafkWlbxHx/eZHjjs1Epe/M0l8fxkCdJT0d0
IrhCIdQo7NSSjwWiVmoXH8MS8c0yYTdF0mUInFXZBoBtefHwsvJfdVfGFzYjaap7r9D57n6nw+Ti
Q+k3rt34Hn0iXH03b8FuF/f60JQKyFBdTuL7Ov3r0UVP6tfeyz4PDT4djPz85h2lsHu2m+nz7t6j
90hpEmbQ6ae4xDLry9iwFohOgQts+q8Ke3J3Fq6GLQ8v4V7naSLGMSod5rl4XcRrF6RcrLieS2sA
srKNvcgvbAjC7OGcYD09Su1ab9mhg3kdiJ7V+9C+AIkRr7YHQV90n87ACxSX9wUNPwU9nQyduIQn
5b0tJdjCyMvfS8hGAEm41zOTRRCkDsv77aCDNchFVlntiPvBhCu6cWjrMZYYihUM3Gac0ScnazsZ
TVx6LsPfrFO7t7oZkv8mMsSVolWUVwutjCuPOLY1ote+WyongaVfPlRmm9dR8nwTQ3sMfJSWM0yI
MAZ10E5ucUwy48dtfw5JUSSYBY6HK0uIYD1zjmLYj8VepxEYQAWuDsqSXkb8I07eJeY3ihyCLIz8
FakoGsNcIvMKOJUx/QR/e1pYmHPxhvJPXcZqSZ+3qaSqxXf3uo6eZQDNamDyvu3PbYSnUyJrqZYX
d/A9arl2DW+kA7e3vyO4sTTUDh8OI8pe/gXC28sS7oGt66LsFV9RPfAG+bdE50jQjO1JBRaH89nU
2VdPKdHvNkyqj8ma7lh9pOkYF/MQcwa8dIoGqkqB9QtEIKHAThVT7NrdmyuRIZFBHO8oAxYohewK
A14DUwDf5BncXv9rIx+t/3ajJs7kw30bs6GYrT7AzW9IFiRct6nFk2FHrnFvEdpsMCMOpN3fVTJJ
7/BqwVZ29bwEmPWgAs+mnYyQHVSkHSGwdaE10SZz8iBTPKnaXobc1xanH7uZRXOoU3ec/vxBeRxo
SiY9qVJZJrZquOGbwcfap5Xf6afTFTG3KEqqzLjZQnntfup+4w9hoSWFmMx2NEWoKVt/PuyidqtK
5UQI+jGLdEv1UOEeuJ6ZzzFGe2mIVqDbLyZGMNFa8/cHoQYijkS6bqoNeWHubEVLzpqZD8EmeyEO
iA9axY/UX9C9M+Cf7vTVig4j8fMUKjjZKPfa0rWEDt/9VEpc00ToJglV9YnSjTEp1066kOOvPUlT
z1GJOKcOJDiz6zi1zkI26mp4Ghr5OU5FAe/GwEgDZwTQ5FFTv/GhAgzXrq6akK5XhyKoSCRQVUJA
+7iW/10as0QAOdIgBn63+ccr5hOBP+8llDzZgtT2qzRBEJHM8IjS48JGp2ObYPst/9diJJS0mGdf
6Wok841abnVlwHSlKriG5Ps5cBO6gtG0zCZvUeqgmC9dy7w+zKQJw/ruVY52ZD9/S5W6t7qnbLku
rW3sGTw7bhJ7g7Ywxg025SATParfsumd6Tn4r5Yvh2NHETEWufP2pEvkQYEDDZlDuyjVejr7vu5G
ELjDRRq14U5TxcCVKEMLXCnPJClQcmmSlp4/vpGjJiKt90ujn9W9cFFlqFlHP2tgVDNls5R00vfD
xygZ5z1xxxuJz71N3HvMEGNMu2Ljs3ti0SfE8jBks8nA5Tqyw9E+i/pGMBY/sXGSgPsvF8L3fYbF
hlP2i0ehH9xEGZt5rhKO6nT2+c9zPI4TbcFjw2fTpb/N01K/12Osl2+xRKRx+oGLnMFpG1KDgyXP
DvIgp493lCC1yl444f9dTZQojcZkOGrsl+BFzc2BU1NjkrNgX1EdEKkyNfEoaHwaT1HW8SVkFdkk
k7YpKECzCjXnrKvHWMj8XwfsOPNZ2F1xjNuzR+m3oLlXmBR4HLk55kcGL+gKR45eCJfRb7iX54Qh
Jka676iUej10FxE5vNiJYojfTkd0w4lSY7/bpHHTK4+mYY2VyY2BOAI3p7DKw/Pt24rKhN/+upx9
ntG/+YVeL74SpRNz416nY6TuKDhmt+hl+mgevqvPGoPr6FEx6bfE4xwqDbWBAAbdmnHrxVwNadBq
HMO1BuE4vAlODIpWQqPPLBZsHv3cEYbXq+p1vPioHVhWSLIQA982Nxw153MA+xunj+GIijUXS3pm
BaQxoc8moHE+uPSgaDNv3qQYeSHukkpGbO2XPPXTj+u2E8DtKhLjpimBmRo4HQ/PXxd2XfbREIc8
PizMxV1R+JXG6T/+EcCNo8wShDCY1x0G21tz1YZJh88KUvWS09ynnBwb0gf/4IRxao61Gv5G0wNs
e34sypERleYzUPu6JyhJbdYniN4TCzH+FES+HvYhi4g/hSVUOpnEPtWN7cVnYpGbqWh90VuoGk4X
H1KncwKd4LLwXrS8h9Pd0s6rifWvEOeRbxavDyeykPhqqGXIiSatGgnM3D8e8SB1of+yIEa5NvTu
2cAN5yP3az5aCZsUCrJF3cp2FMsPLfrua2OXaE9Q9O6cVqaXS6uKuZWFjkkvyq9GHM16WKgiZjZk
yQIfuvoZfDiRd0ILm6S+9U6exIVGYaYocnGQKJqUsHU+3VG4pEpsoEZTkj02grOhAWq6UxaipDVF
3OOW3Y7OcYes9KnM4DPSTVdcykWkne3YXkkjhi+hCplp89wzsyFZmHbjI0pO3Yj0Nl0EvPVp2kn1
kKbI452xXJNERuZ6UD4MUoqtj7C97kESf9AB5RsmQ/MMO/rgszMG2NnZ1MHg5XqR6b83/RZ1X5Wo
hL6FFIhY8uSzkPU8vQnqsMycwiPifJErXQbWSUTGOGkYnHNmMPBUQtgQERltoPyfJqtXrUitJgug
jObI6FKU5qOSXIh9+Uf6Q8s2MI1bO6txwGVFXAe8oqnrgsCxgl6t9iTQ1yyThXPE9QQNauG/5NaI
osxrx+3asOXP5Emorpihsvzf8NPGGj7JG9Pi3EGG6LItzgJsws+Rc6CwrRXv34EnD3YyUQB1t+Xe
JS4akDS4r7bPxtXQYyhunUdY06zii1JEsjxqfU+dryCN8Y5fB8mCyYhCTlQhZlCbNYrH9dY/qmqv
x4ldBAOJWTJrEg0lx1jvBRa5QTHrendfFGFnQWz4aFZi0+MNPx+zHql+/L6CJH4xDU4o2pTlwYhl
WZmCGuFm/XEix5TYB2tGixR3nzJy9z7L7+2MZKKoqzxWWriZQLBX6CpMQsRPSvLE2eeguMeXVQ50
zwRkIShuDWmyWS1uc1JuC4ci53QxAgDskiDSTECAoabxf4MVIS4s5wx6/o0ByJjkwklNU3Upvwfm
WFs1Xw5n2ArNeCN7itKwHExRWbHqqYv3JDuOvvCICLPaAoK0Ro91oNQb8UJDbs0MAaddqpVG4nbE
ryVyCAILfg75qieWNfSPf/NfvX42Fwn063ua/rjP7Iyl6wiZbVqPGeLJybbAwT3rG1/FXeitphdt
JpCj1mXc5hvEs2K2/13FgQMpabLq9VqOf/vy91dSLRBBJnRXHXGWG+SQGCwN8YZeTeGKuzbiI0ZZ
+pvqObpJWGpQDBlOHzNWXws3dFuU5x31YP/Mji7F/YSx7/+keQEHXY2aJwHb7zbuP7BHT1vk6512
SiZ5Is++xMij91sY8LhNXrUKb4bBWWHa/vNEck6cDoJEROUp1h/ErEdsQLHk9CtTqnvDiWJZY2EP
w63N56RBcP1i6G8tA0ZHMRRsP7hMVaVzakAQCh4rcLEs+e6Lq25wuJ/1VStkaWy+Gu+/UEIFncsu
jPv9v0wZCVE64sPCCGSq7qYm5I9QqksVtBu04V4vzMNq/gLkiMhnzvebbBvUKNRsjNLS5vdd+AdM
R1qeE5Ph2qxSwEnENLZgohg4KxcFrqY84BiFeNx3g0GBmLasmuThAbZcEUmrm3yDtMC8vkq0Y4VT
0Z8K8Nmu68z/hxUXdeSxyBowJ8KP6kIw0RoP5R5vW4xIQLeTzATMVVXmO4vqj6ZKz5SV6t2T1a9C
VNwqBjIBs906Y1RI7WSCka0Hzdozcc5XTePWz+TnsaLlJfk4h6AtLy9nWOExQbMk/eDrBRrifAue
BZs15zYcIXJS8UwlOohjxlOLzHJA1rijqB6l08vm7qQ8i/QfTkOv5zmTISRRfDwDa8YXALzIqfuC
s+l5EWhlrmY5Uo9mdCRKmEGYw8RLR7foBIEPSv75qZZ3FKyyI6HIU8HAbZC6LbjEnlGfF1jsV1z0
trr7QTRUZSMHqlJKjHKPSNf4Ji8P5XqoGO+XeLMMjtY+5QjCHXddSuT208+boLY/pjg61TUFTmUK
3Nkn3uD3eEoDmklDQjHWQKcYPsv0FKmJPGIe2sHxDXT+sZjC7+m6mtqxuzmfDjVgNk6OZ88cIXoY
bwLUCPfsUqqC1sbyYWD9x6YemmYyr2Dndc6TzCS0aw4XNG9bseA2dhxSBIWpb5w9BrOVF8PGTXjH
HMX4b0cVOW9SCQBHg8wr4bjbDalqi4hoh3e+2HYpsk8s73Bft+mkBuNyHsfgylO7zquR0hlM3p0V
Xj1qNxZIEkcfWz9UiFBS3Ce2kqftpPEF6lVWbNLsNkuX/YJuehSrVuJGJu2f9Dm+g/SflYcHwsbd
VZH+nGCYjlMrhCuJe2SyvaQEu75G6XjJr2uA1Xd2dFaaPZKuugIZnAsNT3vdoJ8IsBLfupMuwRTy
ugCbHEVSCiSm7OLw6QrQdtwXHY9gAc8SBH87YwQP3onxMJGPuvXihFJEI6RVpfYN1vM8DMFUKDpO
gQlfjx0hApCNBCBZbzcU1kMNXA4ZL/S5sn9beFllBe+2YlEsQzwt4iK6LqGXqAFie2f47N7BvnGb
rk1iT4rqULaaIBQlFQMoSeVTqwZF3iRE6myFZhzZWkiuWMberSJet25XAM4tLd374mACWojvVxWf
KSR5PFWmLqozblDH7q9yZiMDLTXJaVesQ9s0l/Sz5QIz97glyVkC1H+Y4p2N1COdzBPt
`protect end_protected

