

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jtXjITQ50a0ecf2Im0hc5gDMz+eLQYg/zzqRdEOtUonTsMauUR2I/zDZca/cFZRkz2Bn/e1TcNfn
wKr/p3+6Ew==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ANnTEQ5JJem4BDOpiZXGW1BGnlByArgufttfMLkwemXR407wjOM5c7+DduQ2B6Rws3h4VtvHo6rO
wrBVcL7VsvPq1+tV939t3BGzv7HmeOgz+bF6BolXyM301AxlRkWo/0oJhXt9sAWYr7zYDeoXtQZb
l76HOHad93vrCilEPkc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XmwNj23lI8XFGQYG7vF9oV5Kxca20ebqjV8UOZJpCCCr+xVAS7ag+llpfkHEOHuw9tSDfsd4Eagb
WTNoLsXhoBdOAYPEcNzU+W9qGu9/wjx0qrsJ9f6NyxsR8o/IzcMAojV3xWACKEn/35hhcf9UXdPw
jFtFMZBq82H3pspBY7rQB54QzJyh7kwXdtgWfJuR8vKgpz2Bgw+sWz2/D2DHqFf2M9nR9Jj5wsYi
jA2guHzbYFRqb3Hyb8w16e2ODRs1Chv6CQa8J/8jZZjpfNE9JYFfYFbj02jB3GIgpxkUh95YsKVS
nyG+AAIy66AvGO8wjxEaZssb0O8bFU7NUeHAaw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jhiEXYtW8X8urAKsC5DlhfR1BlhyMUwpr7b+LLkcXXJrwnqMhkaTCeeV/MLdD2fZlxbKcfLK7F9V
JGPVeMHqW/OgkDKoPYInFHgV4dQ8+vVlaEgOkFd21VNxhDMogpMeEu/OUw7EcrJ+uVFRL9Y4CZQe
7QVrICfnVX7/1Uf6PJs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fOUx+hBZ6Yu+THnpJi++K5FNQDW/3h2F0eesEGevzvwYAUzmUKIlynhcf5gdgPU7azk/daFeo+yk
Krq/01NBV0vQpvK8q0FHFH+ghuL05juk1koa24QZKqKLJESEoqe8+SMhcjfeA/1/cXTmsbZU0sOR
598davhiRIPeODK4SAJwb2vC+fldvr29ZQPfn7IqVQ1mWsnCoHzWBSYPyy4Xw+6asrFDW88G8kf8
wyRSd13FqmDW+hKwsLgtlOhvBagW21tHVBbEEW2kPEAMrlmNhaLMf5utkD/lTPuEPBItEC5xgDps
hn/cW4ZYOpIgB7hTnFioHxnAEnyoEZ+mfU5gPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23952)
`protect data_block
Hi2BpWTZWmzgd82U9hDdvLaPpk1Fvsl8ET00tqsSVMPcqtKTc6962xqCzHKfjjqF8j5D5eTmoxrd
pgBeyC46q8/1lC6l2beUU06dz5SU+0NXT/N7mXO2AZ/5/Q05KJtNiLSSdv8TM7GSI0DD84GuH4cR
yimPFDThkOO4cqnJMsA4z+7uaHZ+2aQRfzrvzhWJlL+pjhRu2GunrV+Ak0LT9paHrLLWq+VOmvE0
PZe8IF2lfLUj+M2cbO4wiEjNioGQWTb88gFcj9Lsk57NzhgsT8tr4fWkgXv8a9kFd82j7IB7jB9h
wN14uSmfODAy4WnoWhYAYIYj1gUlwa4i4JSW+cUqfPvbdu1R+Tmlu967c1f9czIGz2op0Noahdox
Qzffc3KTS7ptjZSQC1OQfb8SDhpgbfee0mFoN5pCIWgKcV/lpYLCArbXrON+dEZECJxJC9OmpnXa
NPexGIkEv4mQHsBvhIGyQ7s/n6kR26IaXOKNQX4dhAaarYOABK8FIuglvPszud2tKAcjM3FGwBDq
Zkz3mtwex7RW+dTULeBtyf5DGEIXKMjqTqrA3FKgpgWhEJKnprTxL0Nhxr+5TIj2iD/0CmNc8Mbr
u4AEDmSV+yn8xqtztpclPtaNx9fUtnd7NCwgiwf9yX308RNyCzZaZ2OP82Ujq80n9VST+1COuARZ
zXZ8je5n7qT/5GLcGLey9wF1Tb271g79cp2h0bgmD7nvyWHQqVglwKebkNfSmq4X1AvMAV/GMHBE
f6qA3e7DWEqpuVGo7DN/8OEYyGLjqJFvFVf5OQLdnr/85sVCqz2krCrb++dJsELc0Lzz2BSKFtjN
KOiC46All05q41gGqT/ceinpxPXzRfZIaxdx8CJDJfVqAhKnaZMFzjdEm6IZ5vd2j/yaQLFdqZ1T
i2aw+YLONoYXG0IO80VYd8J67QUP78Eu6vyLeNpXNB8qgMgS79VEK/H8nuh1uqrGnUFnOiR/gQSk
FBX7y4m/4fxS3IZoNuAlv8xvRHHlgEm/BwU6qLH6212yq5bWbnqvzb/5sPbEisavO7vAPrilAq85
9lvcwB50lqF/6Oq5AN2Bfi58Ui52dzAna7EP5JyS05rveP46Al05QsdgWYD6DL4pubp89fB9Sm0Z
JQJ54Evf509cZEMYpFIed7QNrJf6jqmwl6Jsd5YZMvS9EQNcSotswrM3hI31ts38PQcI5aTOEec6
k8HR/Lt9TYfWUI3k43rI3E+KIqWio7cxmhxAIT1CxvkT15oYMF/74v2Nij+/ayLiRSfL+C/i1aMq
KUD7cVLJ5Ru4ZKAfIDxiZX88TyjOCu/s0TRyBeir9cQaKgn0fB9KQe82qTINvVSJPCU+KWT3syvJ
81vjJxI2fET5vk9OnrG24R3n0t1ojJkNCyuQtPD7rJKUko+2ePVVmzjqsMQCl/5Txl8eYl3h5xZU
WCTom75haN03As9dx12URd98+82fSoUZ5rQ1ubYD/Ra0cuXTlpvyCfxxHXq0sFs26A3VGR4wRxBL
2/7/9hG5j/WMp472ASKrhp0G/nMfGHfeVHFap/PFrgUQqCB0MOfC5Q8eH4kfV4FAoEYg5ojbX243
vWA52g/Gl+e9h1DE7TesWJ+o+J81WOADVP4j08Wn+taSwjHJ6dV9J49mBpb6I3OXkCn2jZI/TOLP
sTNKIMOCY52G6GrtX7w4eJZvQ4p2ySDgntFawsVkOkul8BzYO2t0sn5kIpuYHHegAYS8RtcbX5pz
6IzJ5vnTWtS4IXOy2IE7cqR/SPjeb4xEHuZWXoUicTVwxEqt7HEel/8afiJ3ffNXLa07CzpNySPi
J30G/TunaJxfJ22W2/BleDJ1WY2yfhywRYStn9P2Wqxn+FaR/5ha85kw7v9TNyES/b20hWXR274r
gAhSiKgDHwqulZlqOGlrvDxOK2WIpRuvn9qt/qmHb9SXeXC8VnZi57dzh5IWabll0JFOsWt7ZPPa
wmomsLlqxrE/qmKxijwuYJIj03OLPqsP0u7rUMAtFMqDA3KajzF9WUXrJAV1EF+HBSFwvhhC0B7u
51oU8m+IWITiTHfY1ZJYiKxLGsMklWz2otE4MzszHhxJxo7HUu6tUfAwJA2up/OF9HPkGC42RsoG
9OTUgsm3jbykG0v11BK9xNmTZqEIjjHmrjy2isK2ST3ML6btj8U/Aeu3Ov8621yGNz1/awePbiZE
mekqEHT9ZBvo6Bu4Bzc67L5v9CNi9VKxQgjVWfCorBrWOW5JvApOk60lhaDilqvsGNoGPdCNVAll
QihTBQbT9gokuGin0w6MUt6IpWa5jYAf9HNRCjLv563LXZ+ZF/MqnL4cqomaqGgYhZEinX4Rro6H
rbJY7eZ77D+xAYTH2t2O2/aK5cPfN1THVQba/fy4ydKbLvxJbdzgg5VFLQXAobG7uKudWzt1e++D
x+85sHGCRs9JG3m9AJyxikDqeZsUsnqmBPxUdAu3NfOew2mOpKycSMJdzs18A8raJkZ9cx2/bxHt
gbc2YCTRC2tblUh3E6zqeqnLHuX1U4Gc8ZXY4h0ZVRlbgTd6RcbfJ9f8HOSFOZI6CXoWs25rg9LR
vA86QwqnXk8Xd4Hbvc+6pS+YDYb3DI2vYz/mBkUljdmYASKySTvZ6yS07UpoEhXqn1imZ+OQTVw5
36E6iJcp10WlVvEdYzEbaMBu703nvNl1AZXWKLPNsmZHHmL2fZR7ZjxpHhy9JDDQ7htRY66+k96i
UQhpYhhWsT4QEzlzKr+/ByPIX3kp3jKSJC7LUeIEMZnRwkI1LgdOfIyfLVeJJmWL06mCiJBHD2yX
EEOU5Gg6NduzpBHNQukCsc6+QIeXWRkphKPqt9GDyPBs9g0e3HxWrtg2whueX7szjJ4zZNJ680uX
69aUgAc1K9Cs5mTWT5gR0C7jC/Z1VJGkbwocVPEAO/GyP0+YYwBWrS2zYMpYIagjDDjjeZtVsp9x
Ap9mOVgwO5tt7FUxz0FxLNciQGmw8Ebbv77ezsxZ+/C0AoxKyqCtRbguTEuup+UmEatKGcFj6OQJ
Xx93mnkEC00NGWhtJVlZQkFI0olEaTyI2RcrrvSnfchU6ph3GDDH1CuV3/LOYBMrlfyLt7s5oOQB
kId6LCvPNWQzj41ZS6RFX0FF+WgXdoQJQewsjtnoqimTGhf8UOOcL9mDJBrPL229gP118rO29XhM
zmkoheF38wPieNK7hkg54CE0m+1kbyGcJbtMolORWDvk3Abtv895h/pKo4fezdUjVidOYrT0Xnci
8JZ+K7OIIjjUVCjjS/Zch+sSb6CbexxfRj59Cqyeel79S8DvCa7DKTTGtbWyAl2AOvZ5M2Cy2N+e
Sz+SWMSF7hQIl7Q1omkYBJaEqnJbsqKDYHf/JdApvPPot5C2F81mC5Mvlor/GTL3uUrTch6dL4yv
Rk1PMUky99DJGlJvsYri63jvEez9q4i6MwF4G8TZi6DItf5k3e4H65ES0J+o27VSYQyCkoN7dgxV
C8wKyQ9Anr5kwzrga9PbzZhrN/JYFbNwFfry82kjVEiKddC7dE068qXgpDczVch/bcCI/LnhkjTM
8zsjTPEcqKAesZyn5ga8wsVMTGaCNoB3Npm1n9urm+X1f/d0C1WXlIkf+4PcWXn2jmMZUb3TnEV6
UfnVviIx6ABfICeLb2H13k6wTZg2Y0ZTieqICvnqIn4eK/U9czpZxbgj9RDU37MyCh58QN7qSktx
FSYTp+TPEw4iAMnzGZki2xcrxX+yY56ObE2oAn1F3Quc3wJuckmAQzpAz1i75xCERLp9spNdoyV2
rzQfcU5AEg+bmANB1ZoPlN3hfKCAnGTD4/Kq6rCIwhcBZEmQdsdPrzDaISlXpo/icRLKJuBAiGrR
GI1nwajbjSOqjMg7EwiHEKbZHTr+C0Cbg9tFD9Bfnhiq4yMDGqeHlxI2iseWyGZbUASYr11LgZ6/
e8yUbUUjYsUpVflgx8fu+OnjeHyEGcWuP3Bl7lxTFv7g1Pxt+hkNTB6wuOx+H2/mqnfefsITeJzZ
esTQKpfjplU+SrUg+DCAcNvKrYw3MtgAQnfjOn/Jp/gUEf+bwMrroFJVY79n1YFmj+Eha+cfN5UM
qUni2OAFewAMPl3j+Qr2K1LNnXkb1dsiwhGBiyLexEMKRvHfRGQsLA06l2asq8eh8xBoPD4jqkFy
0t6jWBFHx+HdktjA2OdQ5AbTYFxrplJs/6/LID4LTx8HRnUISIGGku1ipg8fl+YqcOfXLth728hF
bBpfJ3208MDpdNE+zTwmfDNFi5i2ZiLYuqTH4CVTMRV8ipqoABdpuid/WTqmfghd7yOrYLCpkQOm
/qUjKjv33mdMT962Pl7QNh+2H+uGOuqMu5/LsrA3Z8nsqfeWdg1G79vM+ZmvGYDgQ/gzv1KHvha/
GrKChHt1h6L+BSQmjqLxIYUfH8EgZCu2F2EGyiDbhjPF9WggdRtm7UI8p8StfHhNU3dKceqz2Bzb
pKOYg88Vre8mwWKcicyIszGZ27tEdp1eXDiwosjv2jigZWn324bVz4twiMfU21Ma78eX2OT3tiWB
4RJEe85EUbOpVJPsvQ8JJR/SOELSnegukW/JlrmObp6SRL+hC+NZGSE0mcB1QLR/5u4Arp1wQmlw
rOugF7igSezdVJUQeylEi+wyUfjjpT5KZhiDBf1ZLLGuxG3PgOvKI602Y3Ydy8ukLeiEnYdc6MMP
DZF95hbRkW5dSy/9p2A+f5BhmfLTdxC9ZwIsiqB/totjzHPJUsqbQ3R7y5+Id2hIatGIEyQmvnzH
iGqetK0KKS+a8KC5caj0X55QR/NPNcLOZcpVkMCgHQYUzrKhgSjjTRNJKuXOMHEXUa0VtMzhe1C4
aiGlOxG4Tmf/bUM1SgHEDWunWSC7SMR3oMNKEEkrA+dWT43BsCK8l4Ap85GnG21rzGUZuMITN2Pb
C2Cj46fDPmW2YFap/x0faTtXZzzbeDNhvujKMG07JMQeDNO72jE1y8ONMJLNN4U2iIdQbrG05q5V
WgSepyeZLQbs/8pxZPIMGEjwej09CkfJ3fJ+e0BM71jV9AKw4FjZuA0v3vzEeQlvvFFe79iCSZgx
mfXIw7uihbU9Vp1CKpZ+hzZtRClMM2KOAxZzzdn2kb8DYhOSgt9PbEVxmom+fRXkEQ5YOl6YKp/o
2VWU2h6dVsQdmFjnA86FCH0NQ22JUKddYCqYvlEvLThppuMYX5lk8+cRYpgcvrXQyNn/1wNRGmG9
8/YFF1LfxMAItj+TgnNNhQikZ9a7nGForSmYwxjduuWYkR1Io3OPzZZMkLlkbA4dGP3krVHXJiJR
yhbj9ntdK0UHTsE8fVvMr7jybiMwIezNeb9AQyKc3QB8mn2SKap3SduA8NrOQ9sGzdadSsER3tAv
Afg1gBQPdJuBe0BCfFIjcfRx76JfQ6UtXsmC484xOG6WpJ/Pc6lkziwIwibC4etuDlc1coFaqanX
+++zf9r8LfcYNmi+YnNSkevURwUm1qPM3rt7ut09prv8kEKjDa32y6i6Oj6OOPd0C9Y/X9gYdMf9
O9opn+WB+JPTcJXPj2RbaeO6IT4+AplsFv9ooyGN5H4Xd0qkes+fTW69szw//Oytv/FX19OkZvMK
+/z45TKr93IhUKKVA4yGUzoU6FR0/0SPoikx1UxijMwiuNstSEgCOC2eMWUthVsEFWKU/XBSL6Z2
64qxPzIP7y5r0/i5aQeKZPll6y0dNOpxIRiWt0cKKBHdhe4Nsnsx9WVmikiPobWmcunCTw9pULaD
8WIonB3m7BjZgX8Hx9+fIyfM1H5aSMkvHaISfCpwnUI6xc/moe5bkoKI5D08qcef10X5Dgca01sm
DV7oShdp17e7WY6hRVtTRzN4x7BmSK1tlHS/Q0r8Utyl5WrpKNn9e3Y1FaWFxN9q0XLVAuFhSYod
rAuwtmh77kmky7TlVqDe6lolM8FlhIzSNJC5+597AdjhgZtAXBCehAggOmd75293N3YwS3GAjMc2
pk9tqg/caUZsUFlUey9QpNy03BkKfZERH0hsKtEX9apYP37eD7GQSBY5eOrK3H/TzApgxOI1a5zh
gcbmB6iOksP3+fF6ylEUqhCvSCWzLt6fSZIJRatBL5Jbjp9m18Lh9fxMaqkPY1dCyhE2hV1KARfm
rRw8QkokJL+7cEAocJxBxaohJzGgJVZSg7TFHU2cfmTMcrSBFrQqqMlIYjAn34Zxi3cN9JuiY9WA
KxYBbbiiZQXvxDHMyyBqnxWL0zKwKk1lA78ywEhQzmN7FPVZdmKSWMCgi32nJx0USrkQW3IRmRKg
NI5+F64JmtMR5GwBRDV5KwZLONGIX3eT+AULfMKzrag1TEivx/LLk2baBz0Sk7dkmDQWIch1AayD
l8mFLcKdkjsJV9iToIpTTX1xkipUJ6Z06xX6gmq0+7+N2rjpvqqPTZocPaVqKqdViQZky9gDecQv
3eYkeyN2oiHUbVtnW3EVUuyw1l5/EMRi72eMWu5k0XNYZn/eyAGGg1De5sQSwPLRcM6tP3yhtTE3
7vN8RE5lO/V3tk3yVU8O2IYw1v1quIFEi2kxafovPA83ObxXgEM8Q7mfwM9+z7BUVVAITe2I3LdR
Hb+RHUffO5pwUSUrYR3DjNQTKgS+9+dmf/OQoNgXB/Jg/NqXf6oT0kwrJ0Z1BbDZEjOcEJ8lHfAj
8i2G1i6MamF0BhLM6GEP2D9LJaDPcp6yaz+XfL7GAt3w9PDH+4rSaH2rlaxX31hBQixPI+1mQ1cx
DlzPJSE2pO/86+cS/c+7HXgsNsfXxdZkUDNspruBZm2ZOmTzK4coXe+hQmH5G0s6EJahVGy2K2kk
0cmRafCwl6tkkBeWEnfAGYHztFEPunM/dyf6RzRD059Dq4SjUrIWmIRfVxzGYzRJnnR8Dq4feIYW
lJnS8oMLGVWvCX+EhWn8tNhLC03nbUe3R+vJwjAlqmtO8qCyg/fvK2Sd2YGlskVR9lNexj7jVckr
cVc2Hce11vihSAM6lBeziXdOMqKDQxYxmk+wM6IxD93L2fB788gxZqS/y+IzNYs6qbjap8SM/y70
P6jK9YsYpYetN9g7xU/thvipjzc1jvqSGwZAFuUzjO+xZYBC4TIoDLw7XD74dKWRQ4zSC+vxMF3H
vDE0078lQOTb+F2A3wSHtgIVTVCjswM+JjpEhGIR9IJ+wO1XWFW/Pu5+qOJ//1gAM2jYiGsMDdXL
/UVGftgxde/cuAulWFOTzaI/b880mAPbLqN0xtBQ9cmyABBv8+tvjBhoJayk+xy1Yivv30o/uNv4
7h6HZaFIzyxB8sdGN6P7Y937dxCY1DrsQgbDi/nnv30wLMlOCNwSj/aF0iy3qFOWHyP1wh/a60tj
kLPEHiTuEjynXzfcuN/hd8QLmqgx5WUeNn1BXJNzhzy9/29wEZY12421CfW4zWbpv53tPkxFYdXE
V3wwWaMy9KHgNevKp1XoqyOrFaZ/TwmX4v0khCPchqMS4irGqTb4/Dc2CvXSZJSGz/Br4uZ3/Bwp
3aCHQVmtEPoIFFHkVUt1yp4Vk1uQz+OsLjHcPN2RzFSpMxhkpezN+ly38n49aE7oAiNTW2RRyITK
BwXk9vGBie8PeZBET5H0tXkQWoN5EUf3QaNQYjy0gH216/VFjVCHSg/M2Qe0b0Qc/Vj1qSHRluQA
vQuk/Abv72mHMMYIO3OX+zO8S4pk6ZyDcc9QKFF/uCIr49uEWuls4B/m3lVytX/bAsoze4D2rYIe
A6fIAylfzfeyJ2wIkHU72totWLl/iPwH6A0d0nPV7KmRIsCriraL0Hgq4mu5d6lOJidNnrHH8jL7
ppHnyIjFYNC0N7y2FBaU+TegX3dfBOIParIvXdBHEKbIR27CAraFZb3sfcWbPvlhgp4jwwBFQyRC
mEQWWOWjaEXXTJkaffPNy1QWS5fgoA0jCIGv4s7MtesgQqGyjqwOrGpak8QIJYo6ix6vc1tAwq11
sWKjdA0CYMjuGCv6TClzNmiNRIiEk5FAe3xNa6XtWb9faU08dFl86X1086ZOHWNSFZ+XSd3ndt0+
q2VnfbpC8pghW5PrWVA0m66CpRmDQCYSsynZatnqRFjGfTPc93NJ0btW2ZU1QYrGeSPxYKqp2mlH
2Q5DUdpUs4mVOkdBEk3imbZ76pYUDAyNnlQWtOMQwMcDluyumlWY7yWNF052TkWh+rwZH9WMuzuF
l5NsTfiGmkQnVUjeSc3h2Xghdh8mAsPak7mlN4XmyXkfZgtKTYsLmjcL9c/5ZD+gBGncj/fo/oaj
27SzTcT69hSRmIUQA6pjvLBq1EsbbVuVhryMo6p1LYKjO+MAly8ctb3ro1oTiPyX/hpTRVzV6otN
5Nt64Z74DERPNRkAqki2cSJiPUHhgPExjx4DC8uS8aLKZ2RXnAomk57qEepo5HlcriuN+vXHAs6S
FwVCfwTlTrSQF74exMfC+Il0V4tq8WofgPxUU9lMn541LoqXs/8a1/WsLPABLzwJIiH0aQvIo5im
8/H0kbELy5xkFb3v1myrA14sGHItFkqlgs7/G7fpH3xFFzMb3ZPN6iS56K6Au5sXGJ8E5r3PRk8m
aI2uNdI4y7C3fCtZddH+bF0HP2WyhGLPnpXbIKrq66KMMkC81ElqQb1ZOZgJY/LFARV+TCI4n0eA
DMpIyjDwUB4OViqF0kaLNub4a1wTRlvZ4ceSy4959SK3NzbuZmiv4ShnRO83tT9JdBHjNb93lcqn
PSS6qLPDJQEZ14HQ02/D1tcl0YQvuMxu1JtdLIYsOmB257lM1ozYUB09WNiI9L5cCIh2RPNrJH4u
f1XMls58hKBWf9A1uIaMq1p/Nz7saSb+L8gvnJ2QGyeurmc9PwjwHkqg9TNkkN2kaslu+S2NIYgY
uFVjwHEadRjJlDE6jotKuU7y50utZ3yBhQKPf/3Oo2M1Tw2CSy2FlWNNr6O+Z0NSCU85vfyt9ojR
e3GJCcQEE8dFzazdLYmipdTDA3AgvSjTVp9vhgKaRpkQZYioVlKE2/aAhtmE2bdkx3VTv7woMjlc
vAzKA1Wv4xqnwyHTdyLRMkm0fXXS/NUsPlcZ15GxET/M0YUB+wBu1R17/zxZCkDSwMcIrJYZ/w8P
9pahcAz7ClECCFQp3zY2scu08yp5blBK63DeLQOTNBaZUr00m5y1byYOW4cy1ZcYoc8kqz6Mcw1w
gsVZp+4SeIdX/z1flD+plBk4KdPi/vcBsCrJeQNqap8F6CH1VAmtH0ByqIdrJdF0pzcemPpxkFK9
hmWd+Hy4k4IoNHKHsYShGThDmpO5SwmVEjASRNHFPgw6C+JBqazFStVVDPdjbIAyZn7px4K8MK2c
sg4xBpHSBLnqOjipChEf6AG5bxQnkM55crUG+V3BUWz/sQ5BVdf3aoxIB+WABhQq6egbWIxv4b5s
+YW3Qrx+mJGyr5C4kJhzupOIrWu1uzNcvo7Hji1pJ9p74ukf0kUBa0KnGdHS8fTKjmIvZpjWVd7K
EjKeyDXhBSCjl2RlTqo0oLSPcINm+dqyW8zEd9BpL3XkPnBC4OwB1txQ398id89Vo0C05G8/6izY
+CcSraBaB1DhDJjjpuNEXLdoTrQj0IGgsg1BH7Zt6B1k8AyRGycVXRYScUhdKQegmAT+py7B4H2t
aOUHKcXWFj1XaMPYBBnGETnm65MNz5PFSmPZnho5/kxKlt1YgzFycJjwUehkIVZVDogsg+LK32cu
c45DOU2+2Y7MSlg78ztsmcjcIYzZne95IL75fEPKDkwun10bmqZZ53bRWgQNzar4hlYlq5bBinB9
HotSs//cwR1eqL5MLHjt8CpCnt58s1OC+DBwKDBTiyyefu01OXh1IjlvKN5PYjqBrX8w5zQh9NcJ
6BM2UOslwrrliXllm6rA6SKqAMBtjppbgwOsbdannLKG+I7dLRguYDprid6DT4ATfSFh3bzIS8sO
4GMkJoiZmdQP6ZqnlW0GIunsbIKSYNxB77NFObIHrzEKonX/B0He1EpoDo7RU+Gzzyj0W18Cw65n
fpdoU1IJ5kIFIyHcfWb4z4TdDOabKl/73B9D3MMaecpb0Ip6JpZJNTlNYf9qTP7bxJrOvmUfiFxF
E5IHzs/OoTY8xvx/wtVy3iZ0VgtKxnslzbt3tgQ863T06oj0NyxHdQXgx39pHAGYG2Hsw3h/nQaS
+MpSNHmRpLzHkT5AG9eyrXVj8LAwf3lmV+QGNg9QKVzwCz2ztj5LstHWuyDyLVCB3obmch+pVg32
efcX51qffUUMl0w/1yQcM3rN+P+cC9mReIYdrUK/QRK9YJ5yd0jSBpPKBCFg3JCQAQvMAzhzUeUq
YckNsqNohX4dLEm+GI0kZZBi9md9amomXI9GZ+xs+hUi67vyhS+lH84i2SkPlw3CJqyK2dtfrMxl
KSW9eszAyWWkR4ajzoq2jHeYEpbt681UPbe5/D5fHrylVY9lEtVp2WEkf+T/77v6D6Tuhz7IETmU
O4tIy2hwHbxMY92V03s4AI8+PdyR8Ky6hV5J1n1jtCaFOZfoqZOYm/8eyoV3c6oJqbQVbnptTsFN
2ijYs44bUXqpn785Ipr8x8u9QjaRfcnoL4OCFkdxOX6FsqG2zqRglSqyAg0Oa8LgGvwYDN5RymVV
81zzsk+S2u4p4bwr1qX9AkMPFNrQpP5xe7cdw0klbkIl59QJLYJ0qK6kv34Orbzm6iHyXnQFI2Ue
2Ml1KEtzbeYCVSk75skyB0vysojSL6dpPTfSrlGtlkImG4MMzcEQphiEYLqtDFaMOYYbbx8GUjUj
h/sfvTzoU9NvOVDl+RmM21gQJF7cJlpuxk/0jup9VJC/avY81nPT/i7HU3YxPVbHtwweQqbpHTjZ
hgkv728t3HVpWbbZAS4bGDssc99AaDkKVTKtV85DwpFSDF70staPzohYroTkWNUNVkYkRSd5Nled
xBl6nbSi8TylGD3IfXgZlqE56rbsdQ3XEPu4hTDe+vooQVlha1f9jypG1XZKcUbFTtw7aTGhdqkj
A7+SRZ8OdeIIz6mi3C7a/9/qgqLfwl6Z4M4fMHdb1e9HXWF0DHDxnmXSJAJbs10LD8DS7JPI5W7s
e/8HPi+e0GchOLo74Res8gkoIa9glYnY/kzCOmjGPK++cbkxKVkuSNx/N8u72SOYqXUAILHusDol
Ooaep63H3jjQOaiSEwhkT7BrcG0Qu4lcat8OBlyJ6uDjhtsI4pxh9eH/yoq63PyX02Va/NBHgtw8
GoVHKQIQ8om4W0Ig8X1oqvZmdwf0nmqtur60GgVVgZThZh4N4zdFto5hhswRPRdb5qdlXAafRHey
Xu55iAmYKtZSwBY2hXUervROceOJ1DPKw2TpLVhtkKzxxARmIt6xLR9bxszRkW+yp1fF4P8jjd9c
u0mul80zGjfnAB6V/sBqxenpJmNX8zs5sqNpouKpMUxfqHTU1zxCY/j0GnYOImHMpZhctTj+PSIz
4derk5tmpVolJSxJlAg2lmxPsMikCYPyO23GTvOzpe4OQPF2dkZvoVTHQAjpZ9yb1IiFwbxr/alX
rIuHIVyoiHhegq3YqSLfBhCUWrocjSpf+JXHbFe90KUaXMNIzV6wacLYl7WHQ08OlDtUblwHtyDh
PTM5wnITyBTF+FrKfxyv3o2AWki/Bk7jLinuzbD8aXFpvsZU9sZdaC3+i2HfOFBO3W4LWqV3KAFZ
PocfhMDSN6zi8SJzzoXvrNJlLcT9UVt367c38IxIct4VibCsOVAZKQf4UpKWxPbkrNKsBlRQuCyS
PuFv0goZNCoLq2T9SzWw0qp4WWeYqW1Urm9nqvGLWHSIK4LoLIsnK7SFIXE1imjv3hEgNqeT/rh9
GIgZ+NZjIF8/tlmTmOiRItzThEEXlrXO1vpGWP6V6YZbRfKwZrCTav6qc6Y2K9jlpSZ/2LCt78M+
nVbqX2fFq6U8fgQt/vAq+Fs/lD2FHWh+vNzJXVkCddMNQl5ADtdXzrIXXWbihFQzIxTyakx0XUaK
kN5kVap0gtpB14gho7Jlrge7xxx/yqE44lVoXkPjr08A8q8Hvr1z66aFJRibB3AKEmA3S3wPnQyW
Zpwq0lT5tYFzGpzdlJ8x3zriX0ozGtvCt4UUuu+pgtdQvkkjLku4lD/Z2qqin9YciVIz4FGjIxml
hXC/6DF9Ovf5VgFpClkpViD26bCek5fbOUZ0xS52x0SgdMOyFSC4mLm4F5l2Q1ju/SkVbamjSb98
NAvtDFYXAogOurPbKAkn7/l3wAsSK5g2ZbPnLf81Ffaake5VCZgmuSG868i6GjgmkxYNu9mfWrti
Q6yGK+oGknxrrC/WbLEJrBCrGAdurBqPkJYpIAaaJkWpyaa5ObPnVIYl87ELVg6HGlu42l2a48p2
SwsqdLV1gywFi3aA6RRRn+lZdLdcNRBR3ibQazmSMbQqXvlKOFJ01Gw37V/ESYs1aYw/YxaM340a
Lt9VBUTeoRQsqlOhqZ36WeTjpcGTy1PsshkUQ8IxpFHzP7StZwzhPqsgULIsTww9w8L+bEYNqdq2
CA4DrPXz0tNthaw6qezhU6e3dfjOgl9fXaQGj3nHnf4vogpBm/AFZpz6H1C+JV1Xe3F7n0bnOwLF
YZNFhan8TdsKflelGyTJacKMuhI7z4k8acJGLp5+fpIRo6oAfioKn8HyuqGzUuLSo8VzohZZ3i/a
vNU4pIjOmS7Y6Lb1Am/gv1U5AllUpYm5Nbg3Q1c9wW7YhwZ/XPTPF4w6JeV5h9Pbe8RS2AdmYuKb
kqSpkCGKw3RZlf/v/kCGzGtnYmqvm7tM7oYuMyJ+jv9HQFzFP2e6yd9itK6pLNlj9oVhAdt1km/J
Ljwl5WgfI0IPcBNbLZuiiHFpVQ3/wpYd6bmKv1YooOM5/NXCWUpuuCRCppB6HAKwhlrjkfJWBY5B
N07hmGfa0Q13VhwmB6Jfj+FNdtGyq7wKfM1gAzOJzmSx1vnALHRhOwyveuEhjJ9INy7OZ/57j6F9
cXIYHYJPu1JQk2JjOBStx58bvchNbwxIWic5v0solDbtjOOU66stJujzr5WxbpvTQVseQVb8QN+W
zVy95r+i75IvH61ZrmVjZqyQg9p1yH+9tEf2pFqI46e1WygvpLj5iNYh7PREpGa2etkxfHrFP0/k
7f4B8JTeU7LzNkw1vvnhSNy00z96dQQSj7JZp54CreX+9qqbigufOz41FpHQeF4MOm9+UFfRuBZR
sgJWn6jfKLlhZiNSz8lS9uuAHkjBb2Wo+/aVEITnXJl8k/Ox8P/usZiZx2kC8mr4WAVrOFHtvvHd
XSPuaZgkN/WLlUpl5UWI62bOorKPBReH8eDI2sLabSijxeQtmi77WV5mnktv2evlJiE6XuMb3r1P
/vV5mi8iAsW+tZobdkkMK6q6hA/H6ymjjW8G4NtzVwxFbpVKJqZSZt5bHC/CG5z9CacTGT0bc3qO
PcExwgm9kgdo7BDnwKNCXT9ZyGRpWy7Rxv9Y0XFVZh/jGCFGIfFt6WBBv15swekkJ435u1j75E5w
0/6bvv0afRvqAP9kH522LZ38ojPsibHhWFzFvjzV4rh9HvN7EMbO0BOpc1oMwSSWMZMDEa12gRhY
OcxL8nXITJ1wPpRK+2+RU/en3CHRCMKhKgALIzbOH/uvCsNk9OcG6TswS6esC2THLAlN+plf+A6Y
xefXk3dvJ3G3UQuZ0UVuyz+98wih6WobLF1ujZ2s6Ss2qMAVJs4jDAy2gK8MItS8/gmpEvLEMtyW
6T1kISDk5c2ymzLzAQTAS6Mdj4DjnlRfTE5HogVlU3fhaBrcxqUkAjxCDK7zApqpnT9DFFxyJdC0
Hfv1yOdWIzzia9ciwUMwx1yJ3V6yvd9EAOklEX3cmmEZIzSAERBo9FpqZAMZGN0NSxlqBSt057ur
o0mt08wJ5ipBB6YnSFi+iknZeX0JyC1rxh1WV2oemlGAKRbIk1E8fZZbWNge4wYt+JZQNFWZ288X
OFaMRXzkUt4Ug5dwzUzmWFbGALA8ZB1pGRNAcCvJqs498z07PGCnvxuH2SOVsWXbPZ2IcyiF92jF
ycwZ8HY9PgIj83wMId5aOHWr4aJob1p6q2IpV8fkjIu7dDDA+ybIaRfUDZ/wyPxQa+XnGb/LWpCC
qkLZSSGFdrjLwtlnW5cfbD3SMqIOqR0olPlD9WIxYdD2/DkqmI0zcYbS9F+aKWTC1G7iP9PxuFsy
QmDNXqQIrG0+01DEdVlGFSakf6QXaa/rShQL0dowF+mbwqybYjGI4BKD+mfn88elriCd//jU4M6k
kg0L5WncdVqap0auc89MhNToqgQtOar2pdmX0vP5R2sdHVpPYJjS6BP6iuLIB6UBDiyb9FmxT0hv
XnrzjSghWJhkCr9UHTkYyL7ysL2ZfYF6WU0pUrwSfmcT5Kne5jPOmm4E/puJjs2KBTeXByzn5MiB
WAOiao/vvpZcU1V9flzTCNR9UgKJeRoYU/jfVatMdCnmlnfXtjTsnRiqJuS8TviOxKVJI0cbhKup
8EeNCZZzPsilExTaGdBuERYHdBy8kcziS81TQZZ2KJXA/bw4rNIzDdUikMBShtloo/O1e647uXZ4
H6EoYNoMVm8sW+BaheYreSd4PD4YrjmtzKVxq+tl4GaE1rX7fBwsus7kQMDQIUiGotlfC/7D3fx+
WaBY7ZYeuzp9mQHyWVkyw38S9vn2k/04LkMcAEEkzzprELENV8kfXLwyIyvErMYtRypSYzZLrK4U
w1L0sGr3nS8b5XvGUXD39SWxgP6wwrPCvJLEi7Km5MaFw472nKEWOutL5lGyArl+zbrYqfWYsY57
nzSNDq0ZZxH4+BQMYC2G6IGWVP8Uzo6MD1ZxsKNZvH02oqODCxn+sj76HSqgU8HV7eO7LtaywSRA
/bQK+pPNCT7Gh1jm53n4Eq5wUHd2Yqa+EIt9N1LpmZ5J3V4Id6X8yNi6pAPv7/DrlnVtsBG19GAw
NJGRXekCHlLXjtM8Qi97rOJIhlQvdpA5ABzrCqdY4i+07PJZGao7atBO47TeZcpjjyB6GcIBSGXP
EtqbRr9DK6Uy11NEUsfbePFiMuO+FRYiII13nJWkTFFFW3KuLQutcfMS7W5F5/Vkzb8jzPF47nuA
C8pd+WfIcB8cPO4IW/Bwj48JNJsXyytkJ/sb5l82PhC88v2kHcd8FrMNj8pFhsYKQXAGo6CgZdXg
T3tKUXJbL/Xj4j0gdD9fPMcF0nJRT3BrlylergNHr+uS8S/A5dM3a8hxXsnvR/AN7xi08uvUsfDC
SBjh0ngnL69Hk3n3SzaV4C8GpQdcfdMF78aw31T0VwCPhnWLjNJDhMJ5YzaX5cXexIJIv3cdyc7/
eMEBjTAe1P/zrcbgoY0ywVoKaA7HPTSV9ZUz1oPN8I6DPRPcii1OfiFlSSHXLgZlK+OR5xYhsxq/
Kn6c6QuC3Ym0p+GR98ZHYOuKy8q2DbvQurkDcwNAHdTehqNBXikHUsG2era1O8lfxf2nriXynX/2
SSDBXg983cpi+DVAGmQdvnJuxLj5MWGF29Yl6LrMQ7BXut3Ha8gmXilG3tBbVNkyUuxZHyd6lkcN
zGpdEYONqSEuxgRKXu5v3fJcA9MY1abva85geBgJgYfKyg+eBtzx4zaaTMZgyNC8azCo4rx4V1ru
nZWTcIfxuZ8rldDDD/Cdoqxi4XomZ9eTTJLyFjKiCpt8SznmbCsbSiwwwJw20y5GioosidJBafNh
7iyGz+6Srv18kS9vLol8Fe24tsGuYEPy22ml3LMjMhG+FBVGROwXXyDcNhdQ4UJ0chrpAKWe9Skz
KssQS+MzSI007gdhKisEaSgHCK5Vcpd/j+lSig+9G3eto1+ydAsn4ArmS5DS+JlrP3H98Ob9Yld1
j6z0vhSgCYQzRmrvsi1YKOtB102xtv+wdXGxMAZ/CEohImaIte0GwDI+fk0CLLWSABP7OIVzQEPU
8LD22LXrnjbnY/lrauwXDcuk1ZQC9WzGRnLJpHPNHGlf/sx/6lAtljpZVR73j+4o/oGuOoG6Vqxm
Pe7tRAgJtNa51rVM8RP+hkknXBH7MUjK78AucOWBheR3uKvEqrr2UMQ8bS7iUu+DVInQP0mYnxdH
t7lEYfrQ9rHMtmOWfeCzoMz2FLivaVd7INi1rIwrbWOA4g3JStayOlflxnTR4gy93pDJkiT61ITa
3BboK27DKsZEhgnAK5pNMquQX4OonI/7PwzkrcFx33RcAirUHQ/bQxP0buZgtTNrY2x3mcTkxRww
MAMLFKIgfNbTo8uq8mJDVNohg5cOAnLQ8Ww9Cipiqmy0PXpCFDFSmYO1X008vxcCF6/yTEB3gRHm
uToSVnP0T1eNvmuVSFPn8WsqKMikwlTyiOcpks4TzXHZJXOIL9LYk/uj9xJfZXyRAB33n3ro3tZ4
Y2raYKBh7lkqLTSsgvTTzN0W4KZTUEivlTVI4eGN51BB7fQYAPUfPEtRU5XKphQuEIyWN7FFChQh
jnW+ufEbaAEagzmtYcI71M+infAz9bK8OIPoLnKb2NppO805eN1NHrwDhIVHl0uIXooxG3Td+pyc
P0PY7jNcOd/jYyycGmFuozoweHMc2huSVGSrXxAgX9tGOZmTbIk2q7NSP5SUidtEKhs2dpH/gvZd
MGvJSQ7Yz0OzGO4N1wEmuF98O7XfmtW/69imavzdRwu/n9Yjsn+GmLPg+d5rWQ3eMBnrIAcft4IN
nob8yJbktZt7PGs47zMfvgvbUKCZprdbrHW6A2WmiQYH3osrHl0C1Z47zeX+rwwQRpyckKfAb+HD
lBBnqfcWV+JXG66cDUM7XLz6SCS7HnigCXKnbPSlxdT4qB2umFjdFgVxsT+c9Eg5vd/EI6lYhbAG
9ZB4eh9VQ8WqkaiRzPhlh+aYVQDAAezNNWos+3LwUX8GHLu8uMSRE+0KWHzBfg44bTf5Ikx9Yu6k
X3f9YyUM/A0QEQ8GaL76w1kOZXuFLiLGNgfYrrDYBs96iAl3/vitpqym3Ze7pGfWYqt5vMmNGuMj
8qRlzvK/fcLbXvFiP9c81UGClGedqEW+sB+6YDzA/CNz3HD+FlbzVINaiiPSg+vMXgiSIO4s7VR6
TWZbIpY77yHuxxfFYIdrxQWV1DA/oXmUXDsofU2fyxzZl8UO/RUV1mz5WMCoSr5/t0k9/xSPrkdX
2DyC2q6Am5f4J6P51vHFyq3aENjTbAek46dDqJmj1qPOuoOviKA5JQGmDDlBYs5AZJbgggxW/9U5
3DTLOzEp5cip/28zmYe9rzm7OgTWsaSy6xXAxYe29OewU0jEANa/YPENlKH+Paglm7Ucgy5xDsEL
7O/0XOGfOOwlmxWulewHdg55O7qy6zviZXCYsN3lc90ePON7quhpZDIxG+l1rguRTeZIzZp4CgYh
zxdVunctsXcq07jQj3asjAJHY3fnr+j5f7w5qaBCEXMgR7VB6Wd2nUd6N0hJUd2M7B3s2seyZhNN
KnN1WGgnxNYHJukGsQQAQUbG4odRryt+uaYzKLt9KR02G2bTgpzOZMR3IrXDfiRrb+tIzRBI2qqq
uiz5zdZ/oqo2Pb1lBeLgdGmZ/vMSv+VMEZcQpcDdvhG8pHpVPxMSaaDjKd+Vm9C6qFivIJCsa8WR
I4gfKy+/ArxVeMKWJKjdibqenYN2JO5gON6gSg4QnAwNC+FPGLBrox8kakX7XGgBu+Ggkdf0+Yxa
3/faK2gEyQJxJKl/6ckXebhihAC36T+RFa4rrfbbcCdmBHxmzPNclioKXXlW/flDItE7v+rfKG7y
vQTSy1L+zq3Bh190oi3F7K2qgqHkZm+RLeo0vy9aOvagBEFqW4hujnj2/VgR4eC+lsmoNx1eHVQx
D3W/KKooGHFyd40I3mO8TmDeEvu+BPQxEo5g6AQ733fIL+lUR49Q5KZX0E6ySgLGbo5WV5ZOdlty
nOigUcHNcHwSnFjRRr7DjESyRkcQcaNJzvJY5gyovv1JrZw5izOywc6bm3XxuXEUrE6hZYHjtABG
FHgJWDSqye8tn4ZXTEDnFuprRzk0RS7GNOXViPQKS4wkPkB8pq6dHrK1EeLp2dBkdoVzZeryE+zt
bcooEoyWqJcgaTI58kyeKzqIu5K1aL287no4OVB2zsW554R8dpSZGIt9nI1GTOVV/2a6bMzB/+k4
9wOSCOxijCMeRT9jwqFCfMl42/undqLRac90WmqtYwr46iEswShNHuLvST8LPnSyluH/jaQcV9St
zri4sWcRqXladOyicQvxysFyi8TIaTBDexPVmzojkOiromomFE5CRMi/VlFHo9uLc4pIotNlTH1p
wg1VRuUOwhmueU0TgVv5+9DNiR6rrQs3YfIcTh+3628MamQHnr10fgYotJWBR7h1snH96XIFySZM
DCfq25cNJoE/cCJohHIx3aCyu0VkhL64EU05Ht+u86xm+rOMaZYCKAnPusClX+qnI6kUFGFeNlcc
dH45KURYPbhfS+RTPGmSkLvXVTZqbpv01Tyxz7c4DJ/bSDoDTURAVsp6oniXyDpNxP59zME7zmeI
hfu4eRE98StpbPTMtoV4cdrZ3XgHy/tU6fLFhuQxYRAX0htUwkWLW8W8DBOi2e4fE5oUBF8VLAOo
pDR7BS2KfnUxwjvR+GgjUbOK8cb91TbC5qzRe8NftbFBU0x2XaBewwBf5tR9tMbTIi5hdAiBVj6f
UUrzAD3Lbq2RDuZrKq9SCKduDqErmLIgqh7lm3fKj5m8lN6hAktlPY5di2BbPgCrEQk6Nmt1FsDE
btcZOU6vRjQpHz3tIOjTDUpl//BkzRD/IRQ9szp25VtwYYQfXMUJoBzmD9x1lK16uO1/z8gVQ0sh
27xVKMPlz+ZK6O1bzMyxuwI0CDMCmSznvOG29lHfqvej9ne+15j2OYytLqMZDQYkNcdxK9Mycr8M
aPlM7IZJJ0gzZXNpKSMJfOI7hAaQsb5PCtN1LIi/NeVTKKRnK3iWiGN8KoZZ9SWKPQNhvtABVDcI
Lt4FzzpKy76bzOgCEzEqpRTBTR5H5uGg40CDKuVTNX3GmqZ3VBZ5R9oYMhg4mEuCYrTJrXNe+1mP
quM3qTXXk2Ka6gktJHWRWh13+mcgc0UbIrCDhvY/V4iI+2nF8YrvUI5kA4G69RydyvMJ0OvTVeVe
GhlsGEa4cFmCDhvJhYUDLquin/St+mVwUrqpPW2bJuhol1U9/lbl8PNzm/4iSDPAt+MMlqNNt9hp
FVaf6d89QhRbOS+cYkrDr1Dor2QgBD463vkt3VSZyaVi7O7Ti7jJOOxPe+HaSfsCJG7QeXDmHfT4
kb2eatMgmpQu3x7h+GytyH9RJQs9kKTx8owc0xYvPQ0ap+rPSqBPvriO+GhgUeJzAizPozAUqn2L
+eTCNHravZRYTlKOMaNYYuUxd6+QFICYCHeYRebv9JkrgsyflkrelQi0Y+832OR377YZ+1Zp2hkp
dpIaYYhOn1baW/jaVeEBjDFe+KsPFa6W8pSvNSj6OlLeiSSB1ksVAcL7d6+ilxYzjdUcHDD9Hd4R
fwitSxGnRxwrYx+Sa05ExENr5PNY4zKC3kaQ1T8oD1tbH79cswo0WRZz2SrMSlTly6UsdYtp6gQW
omBwML/dFrjihUkhrfiumw9epwlcl4J6edgk0uFO95ee5WNOMXN1bgSnPvj7BfduA3rFY+eRtmKN
G4Zo9ZoiHAaVEKzzHe06zzEk2UnKKBZdv1fjcn7+Raax2QaUDNhjtYcz8e3zLcSB9gqQIzlCQsXv
Dg5UwFfvhSsasHz1kSoaGCOEC72YCnfGEUzZoxfA/dXjO0YdNrPOT0NBwLXT1wQig6zO1X7FT4eC
ti4ZFzOmU5auMktEebVd1LWURdnRfRIZxfGWbhvRVxmQkAv8hQuq7dtVB6JKy6tYx1nomtJJtFHE
cSVVG3rsW47NCRBVlkq2EUO9BC5J8w+CitVabmJO9iQ0zhijoMLHae8bip4vI7Ap4//DgfroUjq7
p1EuiCgvK6iYtKU4R7ADJ8oAZYlqTcBiHmFK1H7LV94d1EY8gRV60JIKS3wxcQRoF3GuYTv4lq1c
kmbVtkliGuFF4oUl7eWs/UChjSwZqGQzdnI8cmQE+p533tC3PPsvn1tR03s/J1cq5gRrID5Ee3QB
uINuA0/oI1zNxj9x2fOkfe86jjt6ShgSmnhDFcJgQSSjVF1gzDxS6u+WqGa+I2mPh7e8+8OD3IQA
xVz1SJenVtseptfVC6Eu7Zd9svvDEPfDdlkFI5+a4RIncYXbJ6L9DcHFHHp0HrA7deNLaxoqfgji
DCAMyQe3D6/n05dJUm57U/qLxPhus4Sv8XWPYGC7fPVLs5WiDWngzi95jHw96VI1xqymDZQV0bUZ
dZigLhTwZoZ1RD0DuL4APMFsh5e8yhLNYSUKFMiw1gLKjMMb77bVsztTwIvzMz67SxmrtB9lYMSF
V04Ik+B2ufcBHzxOGINefBW2xI5+z4E/J4ym+1C9cqpVI2F2LP/Cz7xRQ9liLAbvpgXB0WrwpUpK
vUUWkgEg3aTm73HU0SjsLuF3wMoVswTl9F22TEHFhs/fcqv22sOK5LjXxoYpiP6612O9A01s8Am1
8wDgt9EZMfpPAmomw6eCur6milkSJMCospfAHHKdOoLkAIpqZxXgg+SaMnNgLVyMmvtCKXoYBBmp
kfUZMDThCW5RP7B0VgIo6eZQV6BWAgAJaYYYolcw7wL5itxj+ToDakp7UDjIPRFPba0RQIL6ofD/
EUXj8/0fNY4fvARNtkRZ07ZMQFEiMEf+JQSQC5lTYUlZLE/c9LLiuTpWtD1cNK0SJZFwdRvEMBYk
XyWKO65JXFS7u7gkic/dEeW/s2GG3rG5PNuiJe1zuZfwhUQOdwRddVy1K4b6tdqzItUJZfDI6jO6
X9LEaqN6yp9KRv/6+45tQRDgC27Fzao6UHN7MkzotLxEIBZQuMrZAcuK73RlY7egfpKOY/HINN9y
tlfyYXaoS4IdRw/pQXWAZ1euZ263z2QE4Ci5AYmjQjYxXONRaipQEYmTmm09I/iDGjz6cThYq3N9
XBJEDG0Lnh/BVHMu1EuiAJR43sN7o2S1K1zhATB+IwZHlKL5tr/euRUVD/l//Dj2AuihN2dcSC/P
EZcMUEJuIzDJ+cZtto5ff3wUHqaqeUKNqHRdJppVOGSokb4HYWF7GoGERPAkascH/F43HuDFIKtl
8prkEf6fZ/OEXNx7T4rZlsENo/BCa+HWzEeM/hfE+qRq2lTVTH4tu3UtWsP1fOmu198nzt/4TkXx
3lNR9ghMMHhoVR8T4PHM6gb5W6eVc6/f0xpRBU9XAEOm8YYQ04ElAjm91FysDFf/kgCzVHgw4RMn
HbrhjDbYtRg5aDhDWSzFGCv2WTQ5Z3kCaidCHbBXKdL1XrIUP3/gwvLpqJNSFvy14r0XK6zthiHu
6JFoYQjHXvl+lFqn4yrOJ682I3jQX3jWmGr3caWU4+lgQEGkS/Uo3+W9ialcvP0yF2E/k8rEQ7PQ
TKGo424Lltxy8yhRx1Gw7OqA+tHGIvLLfs69VfHKkpcq5gHyGnj5k85/Jz/9UaRejHMFXBltKway
JueuvLg80+VLZsGmV5zXMUndrlziSoZnMUuhYHkMO2aK4ZRsOdbiNxMEQFxkJCJJWDFiVGmbNR/t
17u26aSnAHqQ481+cOvfTFlhgoRAjyJRk0f/TVxUZCDPikCyK0xg6o0e27USNMdZqhaKQFzGSL83
M5J3JLjWRO03u/Wh5oojc1VOvbKryMXt64FGGGHRDAAOOqkA56M3wSmArkOgFHhOE5rx23jWqwsm
PwLjN+vAgkjHRM3cSjh7Z/HcCO4vpkxUliJ0H9cslBTCdUnqKzX4USRSzzFvxzk6/W34u1eqgdzn
fbcNZIYwwQLoLuUpUB9W20UJVufDQXekktK5tX48yx1PiN5OnsC0JoNqmvq30qC2PjVRiU900Iw8
/CW26WTsBiMI4Duf8ETA6xVkJCZBEh0j0581743vukLGy/Q6vdH8MPHl7BKzCShuObxUWFUCo9r0
3KtGVdTksPtDlZqgVNpFo/BpwfXFbTAo3s2BCOvEaeTWabd0DWPaFM1zzbB0WPkArRNPO7oF7DCJ
RW6gvo9OgteB1WQBntIl1dAMdB3vSlXKZqbfTuoCTjNIswuOHip4SY/SPFwshm6n8VUF3FvEljf+
ar65WOeZnhQYcIZMP3+SrhkZdd87ovrer9RxLnvcMJ9fN8UpO0x6FtG+9HG3MfyO9p+TECVQ5W2H
LhaYXvt40NOdCrOiRcgCVoWy1gMYdV9ZS82c0YX18KRQ3B/XmZPAK5hj28WPKIucx/vQ1iYYVjQL
sbZvk/4xtajSgnwalNz1qRQ6Aw1wwSmD9yFYHuEhyhvjCO71MWf1vQ0BM94etle58MWs7/GlJN6M
h5RQlh3LNU/IvguV0xiVaja3YQ5KkYn+vujvqge7GxeLjovL7xze2bIDqD1logy7Mc7A/DvX5+nw
7llJ0rIRRC29NYmL8vm4AUB6CLDkId+Q1jcjvpTMciX+21+rxz+aI1vWUC+Wae2q07pJOhTz+5Qj
26am08qULYFbi7dIEKHcyq5Ol/Avda1/7aC5bwbFoxd/9rSV0bOmbHFnF42nt+nWWPSIZ3HwaDgi
qdlh9k1Lz03pSPqBUzBlKgJ7qgfXlHmJ1J0OUyoxRTHXeouL8ojUNWet6mNPMlB/FLBYCFfGe73W
dwoNl5L8vXGFtsSE9O5UoCZjM0rxQ6ZiD+XakB1tGgcDUSg265ScrdSzhO2EcceLix9cxrqfKL+c
DPW8qJ5tSE9lA6/9xfUXPZyIXcl9d1n0S8zuUjLwuvnJ31/cHF8ers1T3RTwyBaVAzd3IaHHWB7x
7DYiQvSuRxdaMhfkUsUlPZ6P2kvIixaKf+mathA9gzH1sLvPKk7+OBApnaQVzACn4emhjQsJD6un
au2zZ6+PamkhGcuYrFv/POVFTG+BtsonNHv9YK7796TghoF1+k8LNkE3pX4UvCBBmsy6TLwpRYVW
aBSVDZ0C2bkiSnItSi1S3x8qIfQWqpT1efbJnTctKtEO4dD9+/LxTz1YbErLjjNj6AX74iX+S8pf
XN3an3YPXpJ8ddSwuAoglEdGHWv8SEXyOB4Umd2B0ffpCRPCWgiU23vn7sXBkFckxH3ENJEml1rt
aHgYxEjBU/PMlyLFMk/kJE4E/iZZD4NSNhzrEh4re7tuoDQdI0p7QE0NA/pW1HMxIEYqAfAiIvVb
Cw9Y3eL3Dni/IKusZOn6CZxcNLVHqy4KragYsA+/9rUY2FTv9/xOlk3kh1ZrbA7PNp0iF5qI0uQk
vsJfAhBl1npHn6UQkH+Z37U3qBVLHY9aJzPBMjkhpj+3p8D9Pg96ih1u1UWaG3hE80tyxp73HzM2
cHHekBRwSw8J6vWWKtyjVfoQ+1Hw08tMk9Gude/cp3SlNsx/7bsCInhQQNJx4H1hvF7aTQRr1PR9
jyL5XE1XngyOnb67OD+Sai5P7rozH/3+F92H0Ec+wF9VDaoPJbIMztKxFUqbBCKusv0zzgUL+LZh
iCq7LianM5sQsxfTg0i/fbDFXuSaCKCoE1aqCs6dOzo9QrWku/wRFX6uDlPr57Ixg3IYaxsGxqNz
MwEw5GW0wM2KGfSpAKc6YVNgL15vIcO+TIJQhYOoC2ysKTB8YZspExyJ37keq/IZFN+v0pttS4t2
qzMn6CMO0tI2H1hKLPUYmnnGwDENyIyrtm8a3M5dPXD4RzepyQzonvZvwqIOL7nbo0Q02DeQbIKk
kAiCdUmenQTIDOXBPU0jUSVCTDyDTvLoSDFHMpgQHVfBRu0OiCt6IuukFJnFUWE28ahXTrVA1hPr
7VIw8BlqdsTtspYDnV6t5/yomRSrp3uf1c/2dS3bcKhIXjk3p39vjmtpU+lwyiyaMyjrlBh1/rdQ
lyqwhaP5fB5gjvz+jiM2af9MoiG4OJIS+sQjKWLWESS5TqPV0PdXKYeUKsz/VmzjgXcmQOwodTSS
PUPg8bHoby+MqZsQj1Q46lK4Dja9NvHxzk97wljFBzXM1GbGA7HSpSktLZR3z6BUYbcFu7XtnQ3+
KBbjPqlCuLblH37eOBzUsf1BmOTiensVZRuIkytZG4en3TUXz4tFADGZe4O7M32SU66ElhSJhdvJ
0DBtgCN3OWY6O0kPGDZw8aKcnVtISPo7fnbjUI20yw7jd7wihpFa2ihrxbNHfqlrYzYrG5QvBNIS
0P0tGrV+H+au5a9yJv3F4cwkEP+BuFaFsuiIFR0X+HTC+wwsL8VCcW86X4hFW7P/CjWa4Ec/hp1y
UjhEU6VnMxfCqaEzX55OD+ksQ/vDS1XEX/tutZ1U1aDRN+didqLjKSqKJc+dJhn5ECoAtVk2oRE2
QltuvEgmCIhw3KX5jZERCdeKH9PcUxOzZ0GYYtdnvXQk6jL2fmH7/WZwqzy/9Kr5HOP5pnk/KyvG
MvIZ2uh+LLkWug1Ta9BP3bkys6PTkWPTZEjM2gqKWvemy4s6ipQlzhFFPwWcQ2012CEQOSfAioJl
S6/MKWli0qJBfeyiT7frSkpoZPIxYRQmoYXViqPPKxkI1XNrlPm+MxlHn05hIZH+vp0fbi1YH4Jw
gvWol4RDenElhEYJBXoXXKzzEkl6QHWMdEp7nG+tijXkVewiJKCc76jIZle2dMJb9d4J65yyw1iq
+roSlBRHGETZ4NBLII1Zx3co/OYDARU298IrC0sO/AI6UJ7snj0dYx0wCrdhjRokMiocnXsG1UTb
pKo1WTsuU6bK3FNIXzkXMHvoeIvU5ch5kVZWlXlmdcUzP0g+5P6zahBYBUZ1ooGg1KjbvINiVSut
6i2qV81GkILzmNKe5guJYSZMPLD7wlPjO4DDax7XK2o38xSC3khfCK3WyyMD+F5UvJ0vEHBYXM2V
j8lQlA0yHjZ6cM0mBps5/vxr84aQwAHKUQeFmtBRWohaSkDXxcRbY51C3e98DHxqlJ46CzcWnssg
3043+ThYBqLXy6+9hGngi4JsKZ9LERHN2HWpYBpMVKUzw0cCcuJzENBK0KeFeGsfOLQswWOkkK2i
8q55yqjHOOKSzfyBdf+/b92+eDfySogKWWhZfA1Tor68pAb8Kpg+iAbxevB3q4NAEFZXO2gclMMP
0zWrG1yoV3ioK40TJBNsysTQSOZ9OyLexsbbrv4PiYZOTiRTQP6LPl1GZSgL60bJy+Bhj3JVL8lN
4/AFmr/fz38XTUYGcJi0gg88Jl1t7EEMb9w85kVr4olwvALFB93KNhETLdYth1Xo3tqTn5En2EwR
hHDZOIh24dy77bYkn3VkF1sSjvmND/jROtUxi3RmlAusNTuTbX5iioVEd5GudWwljvHMdSmzeuKe
9rhB74oTDqITrh+aLy6rGZMthtZ6ssHly/nKBNvRgmHlp6QJLcH6HjZ5B0UbPa1ANCoe3hSDv3uX
21tDqmIA3FoqGZ8Tq5hhyH1SGffNkKD6ig+plfUkOA/1fkXbCeK2e39ncbO/oHSs2yssCGC04wuj
YbFav2hY+j2+Rd0atBvXCFVVV06u5OTvPAuAb+aokrHYa359ehDvXmKGSvmSCPxfMWQv+m7ebuCM
36gQx4rJ6O9+l/h4NTI+9c8BTCkqazNyfk8DvaZJqxalGay3mUyJpOqghXoou+G+kM+pp2UdD7aP
k2xpPIq/O1j6Tn/DSpVLQaHDT1E4uK+wPbTJk0fXfGfGgWapO/IaqL/uIK21SIiL6GZSzRFUlLfj
lWkmRepnlaqNeEcmKbPw64ZmFpF7iCKqVQ/wt9ddAgh2meLouihX9j2NTzgJqq5kDC8mCF+yTRAY
equ69xalS1LrCc5oUFJirWzzGTqmUPOYsfM4kTk0eujCS/Es0m2SqYkQtugnOb791QJcSXh+OtVK
I1NmwAyLIJ1tRg4g61WqoelL3lnryhwwpynx5yAagXA5+7NFNd7ol7b9pfWuOMloBlT30KUxwiod
PsSNEiAx6AT6OAmRhryw+wPboFzU7iCN3g8IKTYdkyQKBy/0i+jyc0SaPhw9ueJfjUNTZHNsK9B3
otkpXp5Hgsd3qqJa3jRP6FSWRs5RHlqeh15KhTTSiCsLKkr+b+c8AmYzuHU1AULOCsHaEEPvoGfo
V7mdd2XGgVktUGGuqC5OWSy3ea3hUGyC3lZBW1oB7w+Hiu+HoFOiqj3avEGfnulK/+5mn+OVY/Ds
tNigfMsQNf8naNaFz4gOqLenJvp2xLmR1+PiDav+7y8RrxlJfrHt+Qv6gTPJ7khxxR7wq1wcuqCF
QGtO01Inz47kwa5NooTxrde0yAy7YEo2bna5MdObIzRdt6u3KRnCWo4FXWRGtPCbuo1GhDPexnYm
mcZcdOYbi8xvmZiLAdtpAJw5RbFuZOMAIw/o5kFyQWgT4jtPP8aiaDmwoBEpbfUE3lp6enFE20zC
XwESZ5oawyqeWYfBVibQdxcd/bvTXUv/JIDG51CzEtnmDDisbrWucbuwjuYoCUsi66A4qPsWL/SE
QTwhC1nRwooewqRzazI6fIOpQ+kOzKKis+VUQhL6e2oTBUI8LSwEReDOy6Y4cEe4CUkhJUN5Ll3g
pq+vXJWmOUnDKKi+hRGT/6bBZIhFaOytLQjgy1wnRnRNrJcs62ReThuiqGSjnk4BPO5UO3qEQgDB
xVQNUBnDAEG4JTTmdLIMB1dnqptrUSj9gWsHBfOEn029DI09wxQ7C/a1yN5lZJJcOi/5Oe8pVvWw
/zg8+poIfDWnwcEoPru+9a3ZOiB7f/MbPFjp2tf7r34hyKhtAEz7ZiWGWkCV8k//JRGffOAmJO6T
mw90Ip0VwN5i9Xm7EZCxg8f5b9WulABWxihcv1HYrC2ENtm403HZ7nJnmRjrTqrFZZJ0E4pcFxoj
4kzjyuxfE8F7zK86qfwie9seVakP1mVspdCKMwJhPUU5muuIvewMqR9rc/mQD9733mGS1e+8oWh9
O+F7ESFMm3cSRIv0KdBTkgfBC+BaSRqbHuOWHX5uy0RgitxZmFiIa1PqjjoqcBa8zPVz73c18t33
E//YnaW9fT6fqy4mIDm0TJ+aJB8g2uIdyAl8+Sre9jW73dzQ/o5X+YP4PCPhs2q4twk0C5br0OWq
5kXUN0vM4I2hASdPXZyhAol4B3H+gx4IaIni9t/ilX48tj4Po2tzXGY7jL2ZMLolgcfUDDq43UU9
TnjfzrPyS0twK5ghAWAbCqZ3iO/xUK65NyNOVDrXRUxHf1zk6KCGho6EF9xwlpBbPhVGMkyRMzJp
iX9X07qao/XexrmbciGQ527C+5ZgJsEecpi5huRHpLaRMY8r64I/KNHGbXBXjR6ANf3POMejWvJX
lInG7dFQwc1gu2DWjIpsqrIJ76jE++a9392V18v8nNBRa6g9hoRPRzAtfLWtWf1WFod3mGT/poz4
aZmKjBlhxutxUNOiMgCNcjG+00otndhmd+mkmq/0TJKvdOaHP48jmeudlgaApb5Ev2X/wXVtOYY3
HPJm0l9KjeDs00SK1MnnsZHAxyZp13rDVIGMp275sIap/fULx+5eS8xoXNLHPEgOjgXG2bvmLvEr
jGw+A1Pqf5cBmOjNsmHT3rStYPguoRyzxU3luWWO8sVxs7rjnyFQJqalicQ7GlvC4hm9UKiA/4m6
fKm1yxxpkqk8eDiFN9yTXIskFzzzEF91KLat1AVkGSM+kPnyXt9gCIE3KvXMcnPhAt8aiNBy8faA
9KdK9dvHcaq/Ozv2zHPtwa6rxjNCTYLbbzuA1jcX0KmyN3Tfkn7cL8avTvZgVUoxP8Cbzi5YK0rm
p9RI2qC+OAFVFB2dtRSJIHv0CsUcmeNoHwLKEABogwEWfjIajgfA709HqB3P9ErDfQ6ACX8/IQdx
UD9Hb4VoZ66jaBLZcP+JW0xTbdRuWU0qcvDkh4PhxfuD5lKiApxjHiaBbYWmevsX6/WVJGV7p5hT
nPlVxaGZS1TPu27U7Pq9xwxn5zBsMUsYtM6A6d0e03A2uNmx5OBiQf/slRzPX7NkDw7Q/pvEVEoX
GLjTvEF29E594l5bLz7vyYv1K8rNEJ9RB0id4mWMLIFG0noPuZySJV7K9Bun+GUllU4ebEIB+k7N
zYLqBTJm7P9upiZJ5IG/6SDnZfOlmE4ejBoFag+EVsreZX5JLm+Kfz8bj/ZEB6UXljry1tJ0d9XK
bK4/ZGIXYKcBDVxmNyWFfHG0+ZA1QnYJ2Lzw2NfL+nr8t3As8i4OQiQB0J1bfXMXFrMtkleCljcA
5xhxSKBjhvB7DCeMOUfzaJhqBkJ9fKuNxH6YaweV8OTDcNZgSx89kEBy/2d/fjoJTnQW5MFc83+M
lJph6XvdVlE3n3TaNQJD9+z94cv+ttexCJ9zf76CD2FpbADIO/uZuRkew9Hj6mOQCFeF03wPk3OM
iVfdhiYjONB3CGflzKNs7FT6dd2Hfc7ulz/98rjLn2Oj1bf4Y4nWtUUV1qX3h0fjKqx2q4SSRQlc
bPrtGjNln8+olMcP/mMjK5x7HItk169DDw8KdTJ9Erp0N0gvDx1iZPU4oFLBRz6JlZ8Ceorifucy
okTdqvl9omxMQhHcX8emBFrfkHDVykaLPmvmFhFnWsiRUQxvmDqzK2wV9xEQTNLvufetC0tee0U3
IFsFMlDzy7qwttV6x4/jpo2ndDvmODs8Yy70RjFFGrC94Ytmd0PbujZem1WpPhIOpgcc9/4KwwTT
QRrc0Vv3M6+7C7lrVG9OoJ8G+lI7NFhRFIQCQwPR6FfxDSdjBJ7Pz7Xeek09karsub+5dLlPlkNl
SCQ3NMqioAWjIdXnncWlnIHAVmQlYwNg7EE94Wn+SU7n0pwkqySV9r8fjMKH2SdcLT/g3xBhJsXF
CYkEZo6PLiou5s5a4MzOfbs3f/u9puUVpU8/gIWSDj7PZ32MrLkTpL8UG3lfi5KP+r3r+y7k0vyb
YKQpwmqFZfOFVLaa8MSUYuB2J7hf0KMLWF/WCiELj1fgPj93iseMk7reXwHZxHGY6NDKVh2VGAQh
K7asXmXMOAxE/EHZnmfMk01A/89T1BO64fS9eUg3Kv6WBIBfkm27qTIkCej1R0Gm2IZp/ZUHoWPr
+MHbwd0ImA8+81LLyzKPXK820XBw0wypDmfICwzawru/9TogGGmpZQmJx8wlHL4vaFWYeLeGKryZ
lmI0wa9QVvPydq2aug1S9oYQgAcGBQyrYh81GzIxmhgQS4vF7wYRh07h/yAyLFeYox7J9vEuomoA
O/mSHDgJ8E/EsqcNE0+Ef6s59ACHxab/HKfnZmnOxh4MBMUYk10dtoEghlCAN5VTcm/hn3ic0Dp/
2hLYzZqpeOfxRGLjPRCs3rZxXI+q2wqVdMdWsYGaU9tOBvZA1+00p2MeGZfr9XZoaZFyYYvF9oil
emMynQxO4Qse7Da2zB3tME12CrdzedZ76KQGhWvLF1Km71Dd8/sFYg1wW6J3U0v7xDbUOS3qZ5J/
LEb1YAVTmtg4zjTqgHK7ot+JoGcC+uONWYGyOE15lH5iNN0zoN6AKteeyagJvptD1uWTdc9NursZ
iTuKVgNF3UXPLeIhf6hxDBwymArpUNMBp3UqSRvwby1zG8ZKnWOhZIDKRelk+Zpu1kdvvzFxf77t
eSA/0hh1i/hQ45vbGH0nQUxNG9AfWikuhUU1mWCHaC+aYQ6IjRJihQH1h12+u6FBTtQIrFNOmo9r
wEbFWvbTwBMz6bvochJeVlg0Bm2/rZX9EknYnmt/trBCwylyOvazI2yJHhxkONFXMkGtQnWWlIYg
5eaQlPjVF1yxJPSN7LPKYDfmzhUrWy//m1mG+jZEKX/4DuNi7wGWADzinmrUHRZcNRKHN2DN6qPn
t471QqaY+1S2exEZziX0qXlDFcKAud6bY8xW/ydhoLb0UfHGs4ljZJQK1R0Nw8qfO5DgTkheLrsg
DqQYWQCSwST8dfYbxKVRS2elOXvTLCEqER+my/3HxkENd2Oe62A5FfX/q5r6U9NYdNPdRJcebYuH
nALjQ5e5Irh6Q+FjhDnDUsB9ak98VDVqWTgCzu+6nO/Hu79WJhE2bwiI4Bx1tro9SfbBfSunE1+u
22EB2e/ccOBgoWUUNQ8R7jm8sjBF8TsE4htsGQTmSgwcfU2i4eXID16DEHWtMHRcFCAdP/4jy4Dg
MHjMB42DWbgsuUdBny5oTRMlbV+DSGru4tmpN87pxyf2KhaH9MvUAakMvWweJQf4pLJeLEBh28X1
+7mVg0YntZGaqlJFUFzIgF0mBJMojfxFktFznOZbJqNzzsKfszEbi5XDzKyHTTreEzmqlXESSkuv
stbpqnId7xa9CLMGxKmn5IqCXVGibg8/B0WWUcdXls1SuErs8Pyzi2trhnmlje0jezcSAmL3M117
M0GunOl/yhIr9+2Hgsg7uw9rQk82lveYQWRPM5qF0COw/Lt95icTnffwfA24CG9GNTxqOeMksqkZ
LviNCk5e+HKCVcdHQAowTAvp+3JVWWam/aA6q6StAr++UEQf6nURoJfvtCiZpnMp0JA7sY7wdfAl
MdsK2SGudo9fTnulS6AJetMMHas01ZbVLv3eneOYFSsJDWlXdsd6LU8SXUDgtS8kQ4v7+HjnjeQV
BrMvGpAlQKOrSQOSu55rOM/+zJBPpt/vV4/evpiUvR5aQ1W2KsIVc+NIaNjRLlaB7FhiceiabQVP
Ca0nEoi9EmdM60VPulBmZML8BJLSvaCmsCcUGp/UWcO18qy83XilHlrs4/paGXsSkvI61Zev3bTr
hoNTk8OETTZo7qaaJmkH0ISqqsjkxum8lQqt8UgdbNQuP3VMUk1HNMVyln6VOnjJ4qn/Jk2zv6/K
a5KAas5VMWfi+d9PYuJUrXM2HOQBVEfTOJ7dh7EWdX6Elf02ztznxZK71SmzIOX5JSwLFrCtrEZL
zTSglrGuJsX7jIqT7iYLjZm0M5fbXwirv5B1fIjM7zrUSRLBfcDkstP3O/j+YMtLxaz/wGR1QyIn
ecM3k9d940xWELzqi9b7/YYnabbkR02m03PwC33TwAQdlTtarSeApjQGG2XPY63JO57gfltkoO/Q
mvonWR7hZFA98n5Cw/OHZnObZ0DlshXseCj3ONn9X9O961HWeYHvQAi+L1KVUQYIWAZFhO0t+d7G
LPnuFspxzFlOrLKg5+mTfWgS/rWar+UzI8SxAmjjsDlR2bVvr9hALaElCn1TZpcXVi98FjCnzk2L
wsJHHVnjzrstc2rc48whfEG00VNPi3mkH44RXQd6fKjBOi4Abm+GWcf37GG1t17douQc61Wd4XNS
2QW3hVhHSftI/9ZUh3WTM4mTHPEf1wd7/2lH9xQr6hGrZ+DFmbGma0rUgsF0x0tz6SJ+IXsSUPix
naU8VNkDu11iFHTujhmHBpmw33ouuJ19fITJclkNB70QUlL0EB3GdD4ZJ+cfXFah+qWdPDCVv/30
TKWv5qMfCCR825Qmu5Imx2aT8ijsCJbZWAt8uovXIzc0hp0LwnQTjrFjcE/fvGLxgL1rQXreTq9t
tN1JMFNFWX4F1o5LY40uH3OB5uK0zg+eS2giWdUKocUBwZ3uY/ZitGOsKP5BVskA/aVbrC2lvkvJ
esdqhdVnqJJwCO+iwqpen98/FwXPBsYKLBpfepV/Wn4tXlZgqqPqR9JoUwM3hIPsvPNJ6wu38SaD
GUxiy4oCazaZ1cL99jUQMfPnS+YiQQCuuE+lr0ogD117comoXlJom21zWaNPShSpwBH2lBpsn9LJ
0VdzYa8xFyNGJRsLUTbIG8ogeUNpOzSIfGjuZmPmcQBfKVSh2z8naB0d8uzXJlXKear48GbW3Wro
LQ7BN6iPoWw/wIIvwzDbYPkwD2nvIP8KXzQrvaI+WDRVxLfOcB6UwsSL/gO+GtKHLEfEnneyy0n1
C+rVPImKziQCyIR4
`protect end_protected

