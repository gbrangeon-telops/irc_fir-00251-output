

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gjKSpUobpdaEiN+EJKINegy9RfobWzPNNvSuynmxBaCaiXpZzE42DUdhJsa9nuNl5zrnRUR14CdT
xujtPqnMVQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VxmOSrOiNTkpjQCdEraeE2yE2mnMFQ7pRVDUX9VslB9rFCGD7dNvbneDVpuQoePUk+nSB0IAqnFe
/NakjC9Wt9azzGAltfbGlSpsCZYTQJMARswgnWL4Fmc2+3tN+okF6OFM1YLClj1yRXdxl+CDsxQ1
FBT8tPlhn++ZNTP2k9k=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aXqd6ynCn5cZfxJpxEun0CmjLX7cGy8EmIQDak6IkAJ5uWqWXRabnrZlR7iXAJjslJ8VJzSbOvYm
rNknXsQKfebDaT1iefkZ0I0Z762iOiWvIR0eap12f4JcJvz9RAzeBAaW4ZyAkczx3IYLwFNzh/0g
2pHrl6Pls+OFuVt68hp3jwzH7c003L035HPpddZ6HFBcZ3MJeQ/LoNxx+FWSqyEG8xTwd196QL6n
uNyNqC2ytbe6mU9D/s5w5KpomKyiSs16Q1gq8Rj3swuI/cDlyu2A84YTnDD1OVt7+ooOZIymcF7C
BaBzVPlYihS6ibZatAmcUNJ2pZYltRbTtDOOXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S9smd62+t/cc6T+Az0vn0kXxFJK9ox1swzdVaJK3ag284vMfjrlnVswyLQNkD6M2BaUNuZuzevou
xaHfzJcTFt8YvMUaEn6TameCIs5/mTCxVsde0MlJlF2crCf3fZHzWj5ooeKnlSFJXuUK/R6CGS8a
2vO0yBw4ZENNd3h5OqE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cOFUj+LOfMo1PTF/10pikQPB0v1eZ+hPEU+cjnPIX80Jf3IXfuV5X+QqrEh3UZH/0+YwNN5uc8yz
3GcUBcrBnY3TVkMqnhGUk3sy243Fxp5BXFf4yGZm4BbuFXxSAKu5Q+k+UOvWrFZfWdNI4lYLdSEu
b+Pg0ebBc04YBsQL8j7TFN2y60Hw4npf4Ha1Oh0Q36x952OAGQt/kpvEYJz+iBAv7Wj4b3IJAFhe
Hz1SVdnrXpsS0DFFqDApZsueRszhz8yuOSjC5Se+b7SzsP1onkP7OL41tcS1dxgV6XpqQDe6m87o
cIvrt9MVp/aWXYppakvqJEuPRZUIN54B2pTOpA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
mOrMfMVDGTw8wf03+bj4jnI34FL0ITwKszRZa1xMDGsv/+zSxsUSjS2MSmAXwJeDi4mFMoEXI2yT
FH9pRiYUS6PRu7R2GIk95K1vNOqAj2tn3ytPmnTMGaI62kC143RnfDmyF4J5MPWB/4p3RgAu6o/Y
HniM6aGDvvv/0+42P7/Di/98rOcrrjz0lcb0r0nLOmkTsGZ27j7eBALpPMHFCfDuYPc8Taqqdmd2
aPMGX83k6t/HKt/9x636rOFM0CinAyA82qFZuhf05ayCvlAD1bzqLeu42dWajZcToCvU45Zogudn
m0TGzpfEc387woSNGVNjGehqUzMedeGeIwwb98Ls2v+TRKgo0+6S1o2JfeYArJivEoAslWGmeM7g
pkC0H//sO5ZLGIxFfBSJzIJa627XsuaetsBrJmWC44H4eSmBOSxi8SCdSwVJee5jo/OKeohcHLP4
vMSYWi6IKYLulFxEDbV7xuP18EeUteWRutFXdaIEsens10muQDYGHO8y/mI6qXhGcstdUoe8lYuf
0vQi1tRvrL9N+d5NMw2Kp5lX/CbAUM2VjC5RNmK2UXEUE3/LX22BUCvlcVxsR8tsOfqC862NAjSo
yWtAWeH0f/eTD34bHFm61az9YQJNbv7Gs8c2fsdAvQSqn2ICi+5tq/H42aQu2CTc7S/hYTvGeHoH
PTRb0TIxTwsgHpkjq8XQgEKVkVWa51H6dOYBWcfdipHbKV44pW5O6s8GeolsQL1nPGOtB59XyAzB
CYhwOpnXgYO0dU1+tYaDueydFbgO4sJsGIPvxfY96NEb6MICxeGeU/CyPly2MR6KgpP01WFonFhp
+aAaQWuk7j+etFMtlV6os9M39IcifWG3EO9XQ2cLflq7zTXOeThCDQUW4kialPtTpabHBZsshMJX
5n3/mXTRdKru4ait+uDl6Yw4FtZPPdZJNPwazs0qSkMvRlPPjj1D3lYqtuJeY4O0rjP9W5gfuEPX
UvbZZ/1H+cxc2X5rJfcso85O7qItUgcn9Jqq2jzh1sDMFP+xyt2wqTueOQNmTV9T75E6NUr9dZ+h
i+oBBIZliKnMgMiLJAnIk3jZn1JRhkVCCfBfhZVltBwYg0Hr3yUSYx1L8N8LujVqI3tdRIYtIy7N
dOQsgnEZcB3h3sgU64QEOADc8z8dCwwr2UlEPCWqomo4Hera1oE/dv6+H07vKMUL2bFnUPbwKjW0
qiY3ZWzN8k2QkTPmRo8LAYI3Vp5+Eldy6/XsPkVSU8o9yGAm1kzOi5k3F/LywPeDvIPrXIIOQP2n
+xRz8NS1MIKK+qTwNYDG7veHJkBe1ViNKswJif9gn/DbhH8hDs2wXtkcyQoTNzN0KRbm+8jVQWWk
63wnmLWRGeqaOeprsHAdpsUvEQCIXHLCAw6de/CAbQk8xuI6hqUOvQHVO9/BIjMbaEr3CPl1HTKd
FixHV/lDuybfDkXrVzkcuLSLu2cE0t76ui5qtJmo0MHjv4h8XpqXk7FDx9LSPyFoV1zGkkvtMPoA
+GIjoKfbJXW7mRF7QCVvzzG33BZTe5TDUnPRwFTuHizkTEYhdFOAjYkRST/6sjE4/byujzg0yaZA
/wepr2oN+NzalYw45f+lckrqqUFrnNjHWsRtDXfzGQofCOND6/xYoY74TkluQ8DDiVByBicASOlv
+zYEIQyKmSdh3hKlcIbHjNcg2JKcXA/upraItYn4pFEGNATpVRfq3iswKba1A2VlnSdcr4siXngF
u3cyF/D5Dx3QpUm3sakan2QwV5iarKEmJirvIoBB/dsKdeH2yJmo6q6jc8E3AuoMZSHRcXGEtHJY
uJEEabVADAYcK4p20/UJZWLyEJtUXEWUB7m1cl7fNix7K0OUYkiBdd8yU6PCeL86FeCG9bDTbYtP
6b8D8FGx94aA7YZ7z32tC7bNgOecwfhcnMZKCbqA2qtu8AOsFW+lPK/13RDJDNSEfxidHfPfih9d
dirP4BnT9BYQnQVjhAv0Kx/HQoTjCmgppq+sbVVxcjbEbi59PMWv/FuRHuQ20UBMDAZaA8eXolYY
A+6agDfUI9RqFuF5+Vbewe1mdN6gz40U/H9ISwpJKC6CSB3GvI3GLFvWfWQNe0DgU85rDLXpOKhg
pMr70lSD/wZyxee7xPsMfCUWpZvIMmBRBX1DhKtfDt5btVJkC3HxjlPQcUoRdddy7QpFzxSz32ML
JkKhfs6ojWBWOX8heMiAJogWI8ZdN8BgWIN/z98kCismqv6Zm1GLwlJwDyAcDeHCaVaBaSLaoXYd
dAtEiAaeUBzxMN2Fn4uL54+JwAcFSSEgGK95Re3N/SGiPEtzhV0qdAreMmIxJst8+mSI2u7R0roN
pgVIS8qcSl0ZBOn2AgCki32WCk+HGH4AXrhrF5HcuCu3lT/2QalAnjvsyNDW9v2EfaVrF3olH72O
LFZLSqyzxLUKNaKXIcfnETp6SgKaBqZl09+vqX4xsZGCVyoM0q4OYaFlE/GSJ8FbZ1iQqievHMCZ
7bs9iY8cqtFK5ZVVJKXYqrGaRyRKHFeJlkM1oRvMpYp7aTK9izGEQ1gV1TAgJ7E5U9UiWKECdRtU
KqC03eUTHtE1Up+A8x2oda8M9kjeDBkfnTbmOpLH3LHavEheZYhxWdKUt2BMLi10XCDTsM19Sjj6
1t26N+L4HxaOAT3uhLvRV/OrRffT8aOugF6iPtTLnaYv3m6pA8l/f9wfj+0ljjPq9lWdAhxGKSQH
0UsamkTWSjnqnIeqICbrmynTrzNr5Tsn+ohohAkeOASNMWwsa/GY0RNfm3uUTShyX37wo812edzZ
Ngj2jnwaXQEWpkPI5oP0xpQRSjML2HA6PEJqkUmIe+6s6kbs5gtvOg10NL/ZUpvkITdZ+Y6j3sVA
ZQP03zEouelVLK9lOKXf+RaHDusU4pjdobnALqmpnn22hGNXArewGThuooZZry/hU56sHE0cL1ZE
GCZZPTJuAFYYTfG8j68RfAtsl4rbeP7LfY+TvNnf4BoicIJU5WAFxUTfex+gS7AcUhViufKMXeGG
j7eAv1eXoVa0M89XpvHMle7wspueoSNs46mYPRCRs7X36bplsoAh+8FRkkckVls8dGQEH4vCeFAd
OFUmwq0gdGRcJLQ9wJmKJPF7X4l4mkwfBQzx+T2XdiiePHvZDV8TRi3L24QYJQS0AOeRQImWsJF4
RVLAdSAV3EFAHBxR0KUiQNO9m+w3YSq+xKkMlqZEAu7qLVncMPYoVFb2huyTlNYsEzL2LOnbN4OX
wvNm5hVyIl4hYbUg9w3Avlu8mvWWIxPZBIu+j0A6lpUYVleQzJhWoABUGwU8bROy5h7UNY/eOiRP
T/SLGDMShYbIXukUsjnvioRfSQ10LolbvIXb0anu0re5Epq2UoasnH8D90NqhYNBXiYU8heonFLK
UkiQuj5O6PANSanbsxwlU8vDNxFMO59nWp/Q4pH6FHju9q9sokCAAWWgr2rGGVuk6b/luvx6nSPG
B2YBTb0EyOkICKx/rI2jSmNvLOVlZuXFqJFbTwn/WLlZg4G/cCPELYUed5tIPdYHSXeuutzePtnB
BL1v5Uq0DpnAy0tsjzqVG7fB5O9DuBJlILHNuqMRix6xE4tWAPlXe7A4jYUgQlRnN9p73Xppbjqh
2xwVnZ7xg9HdtBgteQI6FECq7fj2i9Zk0BW4jWE9wB26dKUZ1Yrng+cucMZfQpGgZElZuwAswcTO
dIpApskvrBtsSO2P57kXp6bORvyJS8H+ZtdwQeDA0FwiIHIED+g+TYf8DW9Qb6M8bEgBc7u/eBP1
GXQZTBh9poJOG/XxHnHvwiBEqMJal0e+yvVuokRB8DdlfeKP2F+XoannAfV4Zv11IJsMisvqo4hw
8UYkaZgRhovWDArn/OcUnHm3JWI/252jEBh8DoXlbV95AfCPuLOBjswmAY8fmg+fBYVLwwDkUJvo
F58TPhPT83+HjHgwgi6d6YkksSGUYImVRWGhM2A661R82XqSk8x4UGasGHf+n4EhCZB8qJJQ7ke4
jiy5xLef4V1L7fR5XVWXyHY8LxS+Yd6scSeaw+bpUYyp/Q8ArIdc8B6wx/OLq1EViNhfPEa6SdDF
iP79L8fghHDmbeiOa5HfyX8APAhDQN4RkSN3RjrzJvJDwCxuV9JhWdSrTHRI326B9Kym7A08qaFq
WOGJoJLePzDpzOy4Pxg/L7EOyrMWYJF40VpPFbPBmAr/4/TQBs4g2Sp4lrxI1FGMUZ6A8iG08eqe
dFblN1heMbGIHSmK1xBAjaHIjNXCKPRFM/JCsqO1iRpq5u7SzwsCOF2P6uUpJ0UjL4Xh39m02U+1
xH0X8mZjr1HOeSymcg0OMVdGCVvgVM0t2yT0pfmQMLb1OHljPW2VBW7T6X58epkzkA8qu1v4zH0D
lxNIR5swTlhqRioyyBj1l4Wk6M1iYGhU60o/xtdNu0MGwaBoAOrhBJ0S/5njghJpngL+6p1zr6hw
VUKF9mUGGuwCFNNZOIepjXCCk2wFLzUpTMJt8bl6qoMknS9y5RbtFuvIKyxIzft9kbTtvPLy2sv7
E9y9q7TnGR7e3RqzZK+3hT3W33B/NL/Vv8aGE3cF+h0jJavmgu5iZyVV7UzbjzAMa0HMgha6QYPQ
fq3LbmDulZR2SF++7DyiPMDRA6GagZYBw9zpzufEmcurvPdZK1fC6qa20AsUM9o0O2QU2zjsrOkZ
XGEO2jQTvpDnrUejYUF9Mly5ly1R+JiYohxvMi2gROngpciVxIx64xQiYFeQQaRBJuF/3No/Y0FH
N3gUOKDcTgzKH2oMTH2jK1uOrUnFBG6V4/8pGMALprEud7lGzFZBIPM4+pwDLTpxA48wcHYBweE+
Y0W5RtAbZze4U79lOfs3ZtUS4ROdwNhIWffE1LF373Wd6FlUUChR7YSJ/TR/PppFHCmurE/c5Cc1
HEIJMS32QWH+i3O0O1AzN34Bh+JMPmsE2XAS3HE0UXJ8iWT5zAHICDLu/4INuTb5FHPP7fv/VwCb
hIA8becsXLNhtq0WbwsibClNaxvoANOVZo4e9W20JbK6jVT3ekqZcrZGI/74pNZc/2cUz7QebbWV
bMoXVuhlXxV0jC0vVRTkDTX686BqVFIWBIaX7KB8oA+jBnx3Y3XGNYRHrePs7/deYKmWlEtnDh79
HHbSa+9iF1YTrWKW1IFPdvgvG4gw+8/5/YtOcugneDYafW2mW3umIVBz33vAA+L7zUeVq14e91gp
zL6x6Dl1AZPmSGfwz5rWCqcKdrIRSu+BYfjVbWdlOL7F2mvuIoohESySsgjzv2rx805jsmkNg0/z
mRowTk6dZdbQvY2uR44AV/BOtm7fcH0ivSpDVisX5pNP9UJgwIryO+/pPR3TLTo4dlKOKB1KI+1B
u8jThdaSTs/5N+fkRTxXw4k1cemXheGHhYdRitz8K4zwGX6l3XALJPdV61OD7I9anrwBrz8ddU7B
imXIhA3tstQVG2VMbRPVeUjxgSonFHxWRzTBGF1Ex03NqRFBtd5vQEygCzKR5ZEb5U1OhbzbuuOZ
guYxJJyZF3ZTJQGwcF5u7Hg+Gj6yoB0g+hvVUPE3gCxCaKWRDk2FUNLkVpyPaXHw+VpmOSMvCU6Q
0ftBcakww7SfjFV+cURB+TdWC69tMJ2GMLG6sye9NBXToCKvkv96vqOpWy8ET8qF6PRQg5bZEq9o
diA9gQBa81GOkn7tQ5B7RDydUwm7TvvG76PZpXeC1DHtImX2ymFbl9REPA06X8eN2bJ4Hq0Dq2w0
iOOOSeBWOHWlCyTC4xBdsFzieG/NJwCRXNwrwf4FKCp1ms4whblAkWGl9Fa66IyoPduFCA+gXo8P
tWilS8hcifRwqoAEqE5w3O3R3i1nQ1hf331PlrTsm7OXl1eMjuoGzOprBqDgTxsK1HbNr/AdbWRs
2uIt1KCLaW/lZ8xuHq63TvasUOSYaUNaLsuaa+gylGLUYgpg9Ip72mnfjkUpnyKns8rEiKd+uo+5
ZQOMyc+6B5OUrXc68jpJmzY1ogZ+zYujkpNqUD/cHnnPuqqhahrWeltkswNpsIZrZf+5UJT+1kA0
O69P9ZiONKnaWCqJQbm9qvqTtrcb+dAZP8dyk2MJ5aOnzi1Hc69RS3zfeeaNnn7vZAPhtcW9jPYB
mRmKCKeS/o1AVPEc812gGZ2Ay6Z2ph2Rr3w0mDLBVA11LlryOvSQEHR1ajVXGZDduI60uMIZbAG+
nvIYOYZEaBhJfCmwBaVTbrUdzNkUrgz8TsmQatACDDCZ1nXi7wCA1namDOcJ2kthoM4IHlwS96Is
HHVAzRvWFWg/r4ygeKhlNOmO4VBVQMclgRK3c4z/3Nd8CPqvrmFmDkV523nbDggpBqlXNcn2KqFx
chGC3MVji1MCSWNlSzl0jQBJ2qHAgsH1ccV22mdT+tbejU6E+AUd/IOTkyCWpyxVSCu+w4JMLHAH
cNnLWaz2qYLyd13JEK5vbCXKuxQL2iYnTJy+YrNL09wAZ0mV2Rg6m4CLAmbROPR0+RhZKQ4V7Syx
W4j1tXgDPnfEBgrsIpo5uzSJ4HPpwu8uEtBII5rt4rEtYSJtcq1EMsV/9QA2HFt6vVyY2Uhn6ILa
LY59Bn4bR33pk/Tn89hb8T9mAnZQbDDEq5Sx7je8cBdH3hWYg9okD4BoWzJroXj/YyKQqXx1UpjI
GeUjROxFLQUmGNP9jq9NCB49beTHfDKDftYDB5PyAFKGVjmRb/MRYxtuYMtLI27XnomAQpvS/VMf
Tl3+TD3ZJ10hehnScRik9P4rV/0lnChEGyxtCzcQE0B4gBAwBiVsbgSDPp1813LGSqimHa4+0Ks1
s+J+1vYgEWCqffWmDgo4Ul31o7gI3TAdWKHOfD1VnaQHDELqjQo9qq56Ag8KIoCAgdOT9V7WuW4P
NN5RuICyrmNRTUcluIScBQyi/IgeLuy/WdFifT3RyNz857odPXMuo/drWia0Tvsz0JXMYxxxNzZk
yiuzPNGp0m9+z4KXdGwcJDRloqzMmRnwEhcJUHOLHDjiVjsmnYyq+LLwR8CZEkeYInLmI52op1eT
fbGsO7c/SO+nFHabVADks0n7yVhJU/5wC0JHJxwxCgtux7LaQnlXagYaR51qfJhzSsOZQ+MfyFVr
DVnqP4+QvVgARalq/TMAJSpanHYoAkF9sCtBLp1+1/I/kZoIvghdvZbdgxdytGHrOh2Nl1NvaNJQ
DrWiNl+4sGaDpRcjZI7nXwREB5WpZCNeadtYegDEEk01eKp8tZd1mWnr7ckfgTpysCK8dwfULJJz
Kax79NrAFKrBIcDdi1FOTdaP48IZQNor7RS8tkSLw/QRINXQj3Kc5oOnNVBjiL1OxVBtjlBZNu31
m1ODM561qhWDBSK27717eu8dhlFaTiQPZeFMtaMz+W75bShTpc9xD+N4THUTDkMSGCFhsDvtvX02
yxalc/ZdvlfIjH3uDNWhajNM4ARzOvRk3SlrkZxlZE3P+zSc2x7znc8ydN311FF8PPBNPvuGwxfM
4leZ+oqsZAMAMOh2rSgqUNw6MjHiAtEEoE0qjNwI+4ZkHplIbrjxp/+8DGBXmNulbY9ai1c3JKaC
LuvRZ6u+o29RRNgZPtzbyd3cqAXVxH8Mb7eUH1xsWk9JkCJDbKjmDvPKCT1PP7KXQicVi0j5wjWD
+w0H4pl+A+2dgFMMCAN7caf6nXNAf2QZS2HXmFB0AAPI85ygERyMT9gOaEmnWq8bk0ZgflbX3bTu
f95I45nekesjRHYxBJnzYIjo36GtbqPwa9dvvx5+FcLlz+O1vAOJLiLUWGNIE62hZdmSneZTSTPL
3bm8RhmIAIZ1lly/zs93u1vM397trtaA2H7NEOb7KFc1FzAqIxqGDdppx3t9DsYVi2afEvQW3JXT
sL1SDA2fPSdlYFxZMtdjriTAHmnT9XhnS5KK3tP8rOJ58b8LOLoxZW0xn1ZbcQLA/RrzfHDqPdVB
m7LQv3SHLcvZ6lpvUSc6gShDnWuar44i1e02QCktzIBm1H/A6ugbvoXpxoLN346j6qM6f+V03OOK
jU2NHTICrA0I0gahiR14T4ZUwGy6XzdGHGmUPiR9VXktWCOL4+aVxdkI7PuUkF1Rs4UEqeWKWvqV
2yhaez63azgxNRUtQpfe5KcpK+5lx63zWUX0lvRKn7b1+aZyjwVyea5l/J1TdszgTyrI3ezHPkQp
z1PG0yRgQMW4v7aJWcyuTWy9WhHvTJtJxTCA83OLY7B+a0GwrIMUbzvhAnFfwx2b6AEWnPKTzKRP
0ENSI6lycZphThAlsJdmmAqfN2VATlMK9iOUUdzfcoQnlVwQemJ3RqHLgw==
`protect end_protected

