

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AAcalZ8o/jQY7YVFFozBN2W4CJ7dtDMmc4qCXcw+X1HsQOWsjlnqJ0ExLq/9HwwPaBdBtHuX8sNt
9MbzT1NoZw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eb9fumGdx5oOSTot8dVQVSjhrvPnjy5/uUjD/aIEqv1QEwLJo5EU+m6JllUu7ONkl4q2pMcv3yUD
DaaWMJ5SKNM9IQtYV21pAAxck+unqu58lsMHcSYeRXYcYP0huhB41kbacBO7fQsq8URHfGRa6NSF
6GxQzFgW9OWA+QBW/NU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EWQNTRM+yXYG4PYEP5SycD9fkQkTTfcM6sgjpG7m3z8pRk88pPYs5UwluFbB09hVSCMPYEKLENX1
JIPX6A6AjJm02cmQD/SZk/c9uIP6nVMvhv4HT2PqiJbMwRsRLnp0RV8WJNl5IwtzQhAltPQm5tcZ
c9/ABn7qb82RSMRxfzibhF2Uc1QWD8PnV1j6nVmyG5zwtPXyKG+iY84QCANIn7Soa/s6m+bpOho3
0pAI7CU0STIdsIAbeZ3h93cun/ow5TnTga8aw0A3DbHVrLc+5xM9M4rs1eiVbJSSdL5Fc7sYK0UO
cAQhBC40rZd53OFEkTfLRVfwRFeSU8VoPsBCag==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EUZqFPEsLcyFBckZdNISKg5E9SpkAkJYhYdYkwRh/xgSz3PN8kMAAO+ttVMn672EPHPSTTeJWt1p
AvumrJCguaLVBM7NIXSVbD3Ckha5a0glBfzxCIJFFOPOOxZ1B+rxQ2W+YUfoLzcw9DE42G8bHsgh
CvpFN0Szn2edsSc6Ou8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OK0W/E9mRq/arn5PVxkw4+3w3BGYpl3KNYb/ZgKXRQbbZBHdfBtfu0H1VHCuj27qhD0QdkPpdnd6
gHcvGTEag6clv0PLJ5PHHHzcIl4hIp/MStOr0nGLUPNhqZtLAZRqiy0IB5ktSoIvGu4wUrWu3P7t
D9RQYPlFcbj3tpqdazX+5GhWSHnpe6FaCtaWmer4ZDmYZIG1oGk2h3p7ggKQ3amLtCrg9RLkGQQj
yEO/bz1jhZ65yzQA9tlLPbVh4inksrXMkvmJzspRm61mhZF1ey8gENJN2v1TzCuN2XD/gXtMbo1u
8igS7KocN9wbd7hsHdkLAK4mTBcgTG5pa81agg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 998320)
`protect data_block
Ab+8rZHho1PKd18d4ZkwTQjSb7iy/3ydJgbE4AV3oBu7PA4RovadEjvgZd5Remdfa8XQRGAiwQ2E
x0L2pATTi4KRQq5SY8ckMzq5rCj4od4it6WkvqAoK0rIGryBBlW1cOjtWHBUJSzXiKa/Z6K3nstt
gndh9fGZ27lPEGm/O10Y3pCgoctxmi3qw4TabVwfXBb+BuAHdSyQcBTEwPJfk2lKnTPU9sugnR88
KBkyXheyyhNNhVc3TzuI2WHnbextz8a+91blu8JFCSw2BmqoEjbLJt/swSeVsPT9TrIOWqHk1UzW
rfIQvMUQ6zir3QNpKhsA6nUen9OrtLXXuK4olzr/SJkGfyQsErvhdn8Ge01fa+0F9NzJ/JfmZj0r
Xvf1xg0MU206+q/pYxh+aCKWh9lO+G4lBA0Tx6msw7duE1L2VreSJ296h7zib1QfGtu4PCcO5v4P
rP9lT2ICAl1ViQuXnMiPvN+qn7u3RP1HiRyLX/TBFBSntwfYSYYygS2G4AZBaUBpWaCS6Vb4yFEw
svd2cnrMBjW80U47dhZ+z1AFqgTnTk2Zc/CIhzLhQBffof3F2GfuB6uJDbQAeZUSBebKer3znMfO
+o+HCyO+cyEG56y63hECOLjRhdPShdyxeT6izwuu3ewtyXMteMZqeOrME8WWJ90OsEghnfDKmkFV
DenUcy2hT+D7Oxxd/wDtQHDI02pcJwyXN+Rz1VII8gAYYmjl4Nb7/iYry7DlMZQGdpYDMyPUfX9J
8ZeNgSsrvg5t7xdco+EgSn0ufYTJR17Qr4qbm+q/KO5O5a7jug7Nh/YGxfywkJGpGCqgRIyU6mpy
qErfXBqUWgDrMmqbLkOepHV/W59o5am9QSu6g3Smvot2gm5HbY/rRyiTVNlddarixTPbJspfvN+G
IYwvIw7Q8+EcNEocxGaCBuv5e8Y2mJxKxkQ4oVzURUstghfsEuR1lxfWqg8ShytIjM9mzKlwXPQI
a4FKgVCYJkhR97tuWmsIa2U+1aHCfF/j9BiBN+UejLcNPYAbalVVf3kAIKrxL2M+1XnP337mlQbi
KIv3Aok5LIF20dosHX2VoTKXE5XFqNKyc5P4ntlN1sshKMxc4ddzFjiz3AQ8dX96uJGVGvHF5Egy
2WZQ/XYjdgC+BKW3t715x6R/4M0CIw8SRZbfa6YZmrmteD+kiz5D/27o4Zi056UQJUtNP0hq3qNy
sJC5XvCB/eqVZQbJOS4OOW+j2jBO60LjO4hrIcZbqAvWJrLqSql3QQxLLjdol8qXwbldp5IU4sZ0
KJlvzG7oCHspNU2FzJjOzCndNvjIGJLBFxYZy7KvzG1PQk+D4oYnJLvlTao+cIpLAQ4dzjePsSRO
zT2jvQ6AQgR8+CgxhzLeIgeRKOU3/Hz7zLbyY9WSQ6AsryAGkPMTm36yEX0Kz1xQNVMZdsq9jHN9
+Bw+nW1mgSOq6z6OB4jqYlvUNchhX/3EEFWyabzqwGM4+OkzyDy4fb+wpzKx8cse5gedMrrfYluj
PkOPg0BsL8K1pMGiTs9rqfKA9uuDorlzzIf6Or11MdPDNpFeEyKORis65niHRA2wOdbuIU+U/f5a
P0UsBflEkbgax2zOGtBivx+KIKxiHZnKGQwGImVLqrnaWP+ntbyrBxXtuMO4V1slmO4myO+VeLSs
53kGHhbze6bGP+7TYFTwXAAzcEOBdjrhbsILABdqIaFiEY45pMXNg/l2r910MwKox9WN9WejjmEG
UayKxPw/aBZZrqFoXhbW74IdIUppVvcviIEZZTn2TuTH5nDW7hcMiHZR3XO53Aoh6g9iqpRP/InM
23yf7fOAQGAlugfbUF3X953HtQbUMgARy77WKNK6RN5ZVLdb7xpS2x6DndBvLZtnZz43IwIP5BzJ
byTA8GQaPaGUCEc1LA2S5FG3JgS9r1Xz8sGB/Uc0/oK3W60GubxcpNOJ6zolSrSJrGpq5HhXcjnX
DcBdjg/1fxwlRciFZc+HVnEinVpPEb93wONF5T+tMcNXUkHpiKLrluow0xORdPUlaN7hUk7SRq95
ItMyc+jDVEpdlUKJ7MON9XYy/R9oQeu/cLi+FLv47SyXitz6OyDcCtFxBF1baLmzS84IzZLbDTv3
/KMDD0hpr6Yfdk/rtsb/g9mK1ekVfsEhBKR9sG39yhdEzXdnJlPFRV4bm3UzG86a6Psu+3f+pEAY
h7uUgphzb74xAnJAS6aOqMqtF12ZQFTAxEuEkV/FtYDPJG97CvFKyY6N9MfZTBJepIhxHMmiNj5F
EUVZ3foPmOTDoRU84pu7huDR3f9MCH+cILNAwx0isXYFLV3Pdr3erXCypaaAfzbeU9GdNQFkLum9
QRJWgfBUQGWX4zsir2/dLOXF+6kLK/wZIrFfEeofy9T2+WSV+0inG2aCqDnmCUiC73qhUTOZM+dZ
OFb8ZJrolBeFp2pSYKztBkpQrgxZ5XD9tBNJmwIAGGYfQbNkKsubfhqPxhNv+meGG3INtQTeg6xz
DnZ1wGN+5jZqe5ombs0ciF6dDBvYVtq/3hMWc12bqOdKI4MPYsz9POXNz1Fjb9cpo5qt+agf2MIR
6yjIKRz/Ko+6LvtPV94b8IbUwWMLDL2Dba0SstQIOD7UggyB9FxGolEdJy91isJdTuMAGQZZb/p7
hIookAM0ePOmf3Or7ENYt77DMiy5VDqvRVVXygq+ycPUGe28wpYbyWQgsobOtA4omLGI/s9EcINk
nyoFlnz2ghXTmcmNyVyzg+uRWMu16l3Ya3PlNUSRwPUBqkcUpalNrFlRuM4X0745kVSZ6/OlK85P
92JoVfrOMvchTzi2MgHZwHlBz8MYpUTLuu1Xcf7h7fiByqt4KC0z94W3d8XmaCeGblCZ9BmSC/R5
vifO/xYGPZcOWePIAsfNKpBYt0c+uxOUEiMsO/TTvld3WfkyMqWHE53PE6unO3W2R6Z7RND+Nvwb
U4h/HaDhMslW51QF7MYC1ZQe0XCkguhTuIa5E3EIGdz22hPiFuwBOFzC/pNWWOVdyuDEx4te+mR0
L3id/zspHADOkgxUHmh3RCCIoasm4wW6wdNFpOF6PGD0nVZDuR6gO0YzXjvsW4aOWE+kAiqDXLQC
dr424fHQSj8a0ogRhqeafnREgsgKpRZDfKJu+bIcZZ22Z1OLmzTVpOte5PPOfMQNInGQPA1Zvf1u
HkdWHYBK7/F59o0WO6P+XpdIGnbhara5/86jFB0aiz5zDQbfDKL0u4oO6zNjI9LTnpmC3DE8vC3r
9motfWks0ZdjWQ/9lVfOJHy79j/YmvFFMp1moE8FFCTnhVHeVL57g7PJXnlqFxOPRMft7Mf+Qq1h
yzI+pLq1kJztBkeY6ZnOmFKQjyfX0G+cZlrc8w4CkudGRvUJAvTQmYa6l/RyUamcldwDb1hXztjl
QtpsT9uM4o2OKEnx2c1k7LjOvzaToGqpU4xCf4IydMnYwAAUUCG22dy0xVTgesi6R+u2E552WP7K
3OuERUkF3U2/NMPkV7Y9rBWuL0txvDOjS2/Bhdfyti82jQe0nmOv49LM826C8EXqp7lDPx746pUD
xxAushoGYHCKo6HD+lGl+DsKqCRJkQxIDcEUGNYAoAVOPk/fv6Le+g7Uu8hLzULIIoDywP5wJBbt
NfKF2uosqLGacGOI5jFwGERKFy8lf7v8jnd2MyrJfBnjKS/wWEiqDLuq98qNoXXapVJxVPNlizr2
gFVyKhdt1eouSO8BmKdkpcWOEVnBCprtgWLCl01B0+MOv1pbXn7mQy66LisLCO+FkzlUrTg1AxS1
f11Rcczc2kRcwaq+BsrP+qU8PEXWaZYPDXdtHjcBA9r333R3i/WHZjhNFKwMbmvc2leNAbjxI02M
HIKrMVNQXwn83gLZXGvfB1RjJUzWea3Sd1GpqdUOnj09z+wHg6Mt4ETQTSoRDtfiI/sr+QqD2SCt
X0pwEWzVTOB13wL+xsH5tS+EFHzTbL2w6ipR9JvgmFqYalsqoYXZZ7dnxmle16irH+RGngBgkqlv
LyH7kuMB+BLRkaXghNaXiAUV7Z8a7VcUkvQIyYnxqPrpbJonZzTzYM9rQoBFr228kJHfm9ZKuqCC
lkigUAVJjz5c3VoA7/wEd0hY1Mz2Kw0wBdpT/fEKP8s+tGSJQdelt90rtQ7p02/GGhS4iy4Eqe1q
oODL2xQKUUUD4umqWFwLl0S1v+6tzFugl0Be9FrqQqe5qFk4k6GBeLPFtqNXjIu0UV5HbKlfkpRV
vMCy17DaqtAftN2W9kQrjaeMZt7YnKUYoVuskQt8tb2MG9i4WfWAUvTyIzYAiBN1xVjGzmRFXlHR
3gjCjDaWGe/KLwrtq/jhdjX+qJgDLRDKpnmaa4GOXbW+vbXFAV3Iik9P0W5KV5ZHKoB6VAsPhniZ
Sfq4CFwDK2p76hlDNOdpfb8wKjYh8sHsYXQ1Xs7uX6FUe5YkIpN/1PBdas5lW3IXuosKD1/wAtzA
zAeNj5Ke56gv7wZQXTbmZM2JELzuA+H2oq6qPdP59iZzyTA9iV65XwDIlh7Y6h2crolgnHGSxzoV
pD5QTM3KCroxWNxVEjZnQgJM4ic0uwuHHQd8UEByQGklR0QjMa7YStOVK/KbTUB/4IERc0BgKPIE
QFB16OzcYc4lBqyMt81MpBGoh1hBpd30ZHAqpEIZXA3AF1MGVobl20+uSd9LwlcUDNUkoQc91aLw
mAPMdN05XPJ+o2IjmVRV7j6558BJfohafpgB6UPWEQ0TQcbsyMiJBjrLey2UDVFBeqcXwy1THpz1
59IXxMwCt2NfbK6ffaNxcveojc3XwmxtcljdT5ygzxKWw4nikR1XGMEg42Bo1FMHyVx3BXDLwkje
Akw8yER0j5FNcAXYJ0rRec2bh1HL2+m02B4WkW21M9nWVxHqzVYBhu+FPuFjHuP5b3TcobUt9vZT
aIkE/lhowZ2p9rJNVHqiOnwbqT67vg3DSuYCRU7HkoXjhXlEzfHTktFwQg4NURDLITOh5B/Ow8WH
xA76Np5RzGybodPcH0Sf9DiMVrJ3c4kxp8dUD2Ptpn0zPns3AxB4y3YknbH468NASFL9zx6PeF0z
OsafUmqgVsYcp8aBqHMGaNuDlkDx6+zJrR8YbK6f08akoPVbUQeyV279yvQqCYXLNfqTXu23uvR4
pKZlsW9sXABHhkJArFwjdDYA4d2s5mGt3zr3lkFxWGtWpbzg1o3YCi1C41hGOxdvLALQNDlLwqj5
fF1vQaBeeEqbjG66VYgYzaXwDy0wLydIibDZaEdGKaVcm00pOYHCIVWJQ053+ajNPFp+Rw6CmeCu
6kUvc/PdkUlckmD23nbFIwHmWZmDGn+qQLk98SS2v8OebGtZvLvt++m0dZxB42lZpF9xjn9ZioZU
LenytN6uLRgnpjbDmUY+eYVvICMJstzI0CP7O63LvoyhCxGGR9ymCFiEl0plqV4mqaXchxxWOfoc
pjlLEkbDUkhoFffJvREnjyJ9pRtbB2jmQgeaadKgtvwtdKiqyyi3sDtB0SB1UcWyb6kUN779641T
b+jCsyVcm6W9s1PkXz9srFcKL2lFIteJ6LZbEzmpYucILRDeTlVzjIcpCw8IdVrJOBZHIYlxv4al
yeS1isB0EWxDJ5Z8S8CRFNpapUpaThCfHN+Ux6tfT4VXamlyQrut2c9qkQvNIIgJ0XsodqpFNgP2
YGCS4W1q2CvvImDp+lZO7lTdzRIc4to8RO3758FX+fLW6qxRzPCtrhiV/iQzUcXJ9js/cZazR6L7
POTD5g1m5oa5QXaGrVxYvokq1e+i2Id/FLD7gX8IAx7eB8RhAFQgBCZD/r6s1ozivBmhftNr2Tsw
7PHxuby4+n8r7g/fXdrBV4tjBiPDVh/4bpTPWJmE0ZqL2+ZaC2cYtdNAS/acXkEu7REVaE3XsItA
kitWCGCbqoT1e1jNjoXKZ0T0hfVT6cimqNw0JwTk6+8gWXhaynsJ9x/e9O+RN5a9xtrJah66/Ikz
z6b16AiGlc2LZGKY4JsGnlGH94/rYTkHl5p0Ck/WYd+zQ2D5zUi6peerCvOVt/oMlERrASxqt9oT
fo0k0gFyz4jEPSIyBUH/Fy7HNWqOtF4581xWyf+t8/rSsK79ozgcSrwnEqYGL6en80uj4O7P7tqh
idmeLWLYOHPPN42OaYmyqQ+D1Bq9H5MBpqFHWjMnnGvsgUBG1qKPZ0jHd6joGJZkm61RWUu/koF0
O++vKcxC247Sm/UkDFd++3a5mercnh4SmtL1qme1a9dUwCZK8yvUuqa5g3nhVzLCRZQ6CWPRib2J
vowWhKpTeAyXMOAZcjI4Zj/jkKi9YjE8jrBnFsL0W+sF64eXqz+OmEshY/QE8N2WvQ2rQnBhQm4y
ceb6P7Hx2LNYJpFF9pzSEJKzbGYB6n9JYvV5I4gmj3uImLEqnNACFtbxVGDyV6pKVe7sXJ86k05+
tc0K3NbOnYTjd1zS9T2EdOFvcaafwwTbwCwLziQjV7Mnt+Xss7Is+JVreo6LVunESCDa3ZRhgpnZ
CQSiffZ8QrAf9MjMjp2xOwccg6KceIKJ8jY8j2XUMVNE+7v2SGyZ2KQAnSZFfmOmf/sPGs+SQ1sT
ImWI8FDLFyOf2mCv/rezlQhzI3KR5+JQBNx41t2IP04I0ns3M/iNpCANyq134M70aYgDdMfIw4sO
LfK4a/4QO54tdKjcxA03qP/JM1r+y4mvY0J9ISTvRYvVIMcS3LpkDKie2A0kuyBWRwuQQ8Tivqwk
iarKyYgyCQihtoAmn8AEDmCS6xgh7xhmRw0TgBlGWL71v0qa7b1pE1Ra0p+rvQTLs4Lk8oC8sKzt
TNLPqC9u8ITyS2jh4mgNvtHA5XUTzsHcyiqhrHWPtogeuh1BjbK5a7q0HS2NVoTtDzqeOyPifspD
Mt7p4Xi/3pI403Y3NWfmmiH8BIP/rB73h61hghARMqOH5P9HoDHiM6gHqdkPlrtgMb8XLCrZrA8l
kK9o7vysT2bPlbvILjuJCrrZOsGW/4lDaPc8vlsUTLAQEgqORt6rNAgQ9/7+AUKgCldGToAWuBEV
93hj6XKGRoEnfWOpd+v7MUzBrXoKpn+Kciln8IhGTHTq523Y4rpdUAIvb22BBk6N04lul8yt9c1c
iIclEzc+LZ2sZLxQSTvHbelrp57yL8TFfmmVJMujGF6tTXApd6dfHy76/qELm5Pw389w1ag9v0xj
xBdzJHDOmWIkQptCD8C0YMJy0vTBoiBTDYkV7eEOctpZDk+tfBaX9q6v8dUXDBCUYUk5GDEAB19D
f7JWbsqb2nlO1ktyXncGfc/wfg+3yALZzN3BAe1w25sFsobNIvNAxynakXDKB8O9++ZjHf92/cdR
itQeh8UFL8rtagM4VAi9sVoct6kw8V0ig6pb2I6E3XKuc1DyF/QQbL6QzM6cj/jMGA/IIcsroB/+
OHn6RatCA2AXP8q1TaydDuGL7mKuIKuemvy9TDWB5YCNlT0Q1/bIXhX5cOqFl/HNfnzcXJxd3f3V
ZpDvwP2VpcVBqL+Wu+d8LS5vw5/FQyMoOYrtAxiDdtbl80i4VwgWk3M8/y2ah+E1mRYq63gpLEGB
/cvCrCgFVfChcP85mFWOFSRoYnr0/Cn4E6+JfpzeTPNkgIlBGOtcZLaWmcxJreckrDXPEdP+pox4
bQmvlmGQcFpKIgJReafuwvoOsRke+hIP27BG0q9nGDRHluOTNigQROhgXOan6LXhseHtQiE+4ZmV
EAWMjW5j/J+mfDnOLMZfZfXnNwTkNxJkVmx4VoZPjoZHCGhOTEV7kMzIus4UNLtLJKgmz3qVoIiQ
bLh4bTpbWQ+1RkW6WCkQoyfZ5m58q40jkeeeSuRtzXdCppLgnVStOyEBGVZ9DQGtzkSWygX3AK6c
lwYOkvaSWVSwSad9QHvpq0Xd0MQJnQyUVmEvSAg2U8Z6xUy1o09FUQiJFIW79wbCGMDOyl4DNN1u
zB5q0I9p/TRSOJeaHnl/VmXPrmkzi4zepWoQ041hk6QgG4wwsnAvN3yMQQ87kv0CgDRCYnNKIlYy
nAdCrQFG/dx95fW+qp4bt2Dc36QZmWd4cjmjOhe4BEeWZQD8pf9g+Bf+It75dkwQqFZuTmBY3ap+
W1WxXQ6L/lUSjZRWssRqKPVG0d/UoXusebnOBVpvhpjgMFOG0vig1Fv8SROA3DRfOKhDheCMx03J
fYV4D3lw54NTVo4hlaLdPV2qoofNJa8KBZgP59ibPbxyMcsUVNGMbjecPj90CbS0xq/bkPh4BC8M
/kuuE1rv9kHB3jwPARAw+IbqqNYlqhbJmq4ZV8R8vPMXWyDKzRNCVYZl9lTxJq2x3iHwxwEgkVKf
Loz5V2Hrls23liV1cMLPsX+4peT+IhCjptX1kY7m+MJuQrqZVG6JP/xumbppezEc8oZIS2fGkxgt
rbLjjpSb9IY6M33sVdBez7kyrR42hvOonRD6c8vdTDkFEeAm5h+U6LNWLlPi4h7/dVVAUxieqcpS
GtFIYuJNidbNUDUHHLT9F8RpqYmOYgqDTbQBjOtwc2BITx3tL7hih2op/3U2y8LgoQAGrhNc+0bG
NgxFBFomydIiTPBSRWw1FeOVBnchP/NYjnFBLo76u/omCLLw34IVHge3S/sjCr+d77RT0t43JFfW
Jhd7fQdvteV7IrtDshe5X4QNNRbpww74rNHKap+P2b/e70KgiPaKjsLQyH2pWHCPm+oOatcKyXx4
OBwMSuDmIoLdfn7NYLJoiqlrjvvw4zmBlEk3nI3Hk8Ud/QywJ7XOoSt3DC5cpn5XHMtY88winm3e
he0qJOfVU5VYYShJ44TuSdQwwnDqT9SJndKwoXHuPnBvqiUKlsJSZ9yeDC/3WlHUIZWbe6Xf2I8k
4Dm4NmNHIf2UiCCBvhbKkRy4zoEhKjYd+UAr0kfDkVYQUNXDVJflzsVkrBTvzg78FqVCwEhycWCc
6eRZPqzKOFWQ3EyP1s4c6FleF3a41a5NsZO/CkDUD2+Nw3huOiUEvac6kuShjN1Yw5jaiPka9dj0
zLSndFlCAmkSR1yV7GfpoqNyMJky6vK5toFV23Jooee+3FTAjFgKWY8N5mQmDuzI/Skb+nxyLTBG
Es2eP0lhtOUQeNhDfM9WSWYtcEswxCzzqGZGsr+qmZ0Zif4e9ugZ25f6/PTz7JKlhvwXvMMN6HDe
xmMxxIIDRgRHqca6k6N7xczDkokdikTptwpdg6Lx0eVc7Us16Q/Dx14zII7g5cqANwKnRijM95tP
V/CEyBQsLyziDjma/atStLju+TnF7RjOOCa7J2ijbZv481Ty96qTfedl5nQNYhcbUeYkuwIgnCdr
0WV5OoJ3oPk4RrW+sB52FnBsce7Q4q0qjLxvJeECczONwzNP09uutbtqR5/V1UWX+yKbFT/YSWHp
A1hhWNQXvPsSL9AICqJ6FmFNh7EoSGe1yepT+fNu81igiG+vqehFAC0KlQ9haJ+nv38rIDPEw/mb
DdN7WQUY54teWVFYCBn1Iv5A0z21TAkCSNlXdAZfIppwb3i41XxOPbWflBu4KBbSbmZ3WOyvbXZP
3Tlb1sMBBdaZs6JCK5S7HqBPBIc5dhL+/toPoJHcL5QTO+CWAtPlA8+f4mpa4XzjhEQ1cwwarECE
YmU8OXbZ04R8o0ZKRXk0jNpCa87L+tnXr0pIe90Krk7+27dPHVVN1M+JbddChdf3PGP5gLrsWTqg
00zh9UON098Bpye/JQsOBy+RJaYWW0Zkak8jpGhneC1yrgCg83QaZKr9Nrx6Tg2o0bLotr/pGkYy
vLFatOX46U+HJzgFw4CHf2eXQem4JW1wonb0LCQu/xgPGxeiyvLYPpja8U79cnTMroNflHxt+fpD
BBDuu94j7JaE43G7ryYmGGfvB4f35uotNaoc+1yEtx9GAWjdtbDFMgeQjtQQ4rPKU0NwwRFZnDba
eO86Lhe7kfY/BvCe3ot8ZHXF0AWy/3Babh+ETMhnMxw/qtr3p2wm5u331gGosMT3/BwtqEnSoyjO
xOmOjgNRmyzVRJ8cRSF/Ko5RMF5OnDmCUW5FTWtNGJ2LSw3Ff8BW1kKiyZf5qWyzdGqwBoA8Yc7O
c1OHpKU/0AvNJjj3CzIKMUVf1Kga/+C6WtRvRANJMKatakZrA9SBoETxwKequhK88JXTZLVyGRe+
Cih/SWV6RMIL7km1nO011IlXUWsLS5eWn8rj4AJKZa7rNbShkkvdDEvPhZ+YgQSH9Nmg9aIAnLIV
lhDayEkxoGQrVrrHdEnT9YO6l18wArN2mFia6l5C16BI2oWaa3i/uDiNmVtuc4beC17/d3KhuGCX
5ihHlphetLl+hl26QLp1Z8TkG1Ou4e5AxlyMVZ20beK6mPXKHTxjUAbvs41MCv8dVs+1oZDlg5ZF
HgXctnaURyt/CzaTOeSOFKr0ijXfL/JR3ROluZvFCR14R9Gy5jc8iEJsb5kGv6WXXJ1+L+1X/DYe
7kX6N9c8QGZBhC1D//eoW6bioZ9RGmmb73mfHbMjNVXzxr6L+/1HB41LL2NpfdMmSfPpCrd9eFZu
cAH5bfZhKec4kgu7bswMCi8kYqHBRRdJwK+bQy3YRnQ5Oyl7z4IfCMgjbLv9RFCNupBcobBMSWKm
73aiDK3twwynItfQ69F5TiH/Yrw/reRKYsrkYUUHyuJ60n7yg7EgeqVuKnq2nGJ5Y+FuFvBNoxA7
F6XX7y8V2WUUCAw4AfXiyJ6ENHR8D/Zw+p3LeDeq8ptZeW3AAtkhk6pXQp7S+F7r5YS9X0EcKe5t
ZxdhFIud1DE3BeH2JQbwoHI3o/0VWvETczPWxv0jrWK4Z8Mri4cs2tAwsCq2lrZ5DcJ7xTGF7Ky6
0edHzRICnPMuWw6SVfDj0uR9Obp6YoN99X6mn4JskhS1WsZ29yrtXs82n1epoXXLdwUqJdT4idVy
y7f19TMg3V1Yv7zvL8FAS+wBDt8FBVwpPXPk5/CwPEr0KSXpOqwxOmGXukJarAegXSIC2eOb10Ne
zCGXpRhZYK5CYVXNbGxv2CpxxbfD9j8WqcZDeT5Ju78zRQ2rtG2k/iz3GpfNO0yF0GubaENdw/xq
/bMz4AIbLhvKdxpdBphXsfXI4+7x7IbSsVeF9FE7AMueJRW3EO6HnDaooRMSOiE1d/1S9N4X3T5j
37AwmIGJ8T7TUrELOCCLqIeERL9kQcqEQsk1Gxnxyukm7OpDn4PMszFIBLAW7OK59zvJ/I/wBmnZ
/6NxrinpjZcuZ5ViN2+ckmhGNBnsl4NLKB8xidrdrLhDXO8IsKpDYjb2YZaQ9HpmBVHmpMYt0AWl
9Ok/91LfAC4VbpHANdtv7uowXOtKIJvI/j8zzzkaU++HCdmkKbGQvIK9cF3r/c7fj8Vc/iJbnTu1
PIiTnnkpp5KoYzN2pWwEn7AtnAmktHGSu4pWDrnmjAYE5C9DM8cEb7MGGd5CYgA3RwirNk5Hj/qI
PAvbJM14mDL3qrikv4iUTc0cU2Xxhtm1gkx6EeojhJcdwul26rFqbX7aVTmmo4sDoZwErHx7EJM4
uxMwgEyv5XRh3dfe2Kq8PjHI0Ogxi0/+cAbx9t7ccWgNu9G8B/6iITPLbd/DfBuSeu2FZzj8eQHa
How5Us14uc/KfLbDhn52Z3gBJBcbCMHWDk7ljjb5PYvr/vAbsBub/8+8gvv5un3y1xzpPixfwPKp
V0CHCVnOVBR2uhduMjpRoMkuy6a7vRSiro0P17Buq8vds3bpgrigcqzbvbK3sHQYiXC8ylKRUuYd
mrSu5xG9h2eiO5PFn9Y3RNb4sS+tmFJ1aVMIzg/9p46acH9zJgAtf+ekz11qtyM4ZGZSlpomIFnr
PsyBkr1egtJCVCgrejMvxjYd7TMbS7Do6fTC9UoLYPUIAQwut/rJXeO0lzrT1/QKtZjKJripHVYu
HsNAUuq1/Li7wC7JwlOkdyygRPN7rk1Joq49NcFP2FvC/SLzPddSEcunuVO6W/vUYy6XSWSVG0s4
tFqqK+9BtZwQkVEkf1fSbLgh4RTovjKkeRiBWjoEjZUr2+igDOm7wpVhz1S552OSvNFo8BXUWzqE
EQZ0CVJ/xWKjAWHorYRCj0p3oYjmHWhBL5aFSFmNbL4nsrkzPdl60H8kwfhh0qgqAN1I5+NGzu9l
76eK8r8yme+9elCHwMIzO0v2v1SkvrH79XmXlOABEP2u01cc9wGMpo/A/LXzA57Zp4cNHnlpYNtF
pkgOWhTijVACWx6JjHOW12uGLNfOaBcapvJgWyphuO4aCQImCGJo5kcUx3DoE/rPeYM2AYvgwCkx
CPfY+v76DXKBCLiC6CJty5Cp4UkkNf6v+ymWN0gm8S8kAS/4wBXmSs41TAsPX2trFwXhzi1n8IY2
B0faFCzCu24oVcoA7H3lC/VLFPJgTpp8uRgZ0TG4MRG10bYrlLMleMwutmf2gb+JpSc0GqjXOi63
h40hmSm/gy1kSdeY5b/LMCXT90NVdsgYAsP0qvxGlDj0F5nDhyL2AFGMLAGvh3qW8JWpa51oxvxb
4muN0+HRdADyy32wZqv+rSf8NqIto7oHgmnmZjk2m5kXYFnreTTgY8tCfDB3IVAcXrRUFFRCJ2Fn
x36zNVTZPb5DWLSTBtTcY+YQ6Givugzw5E2X5OAuo0ceNzXyMIxTznh0XfCAA2jtMZpvAxVxeq1Q
hgDsZNiU+ilasqcLZZQE4wiOJFXYVgmBCJZz0VjxZy1U1mkFwEgrXUwFPeC4445pMa7+8zQCF2FK
HfbnLefsa4YRHbMf8rzPqiRzotPYGAPv75BO67U2c6Bu4d7tpvUd9HEXtBvhrufgLQrj5ns0i/wi
L0tRTgCv2OWyKedzFrK/434jx8kVb3677xPGMIrG6MZKQ7KXWYcQaEtL6SaWD/agJnnqXSWYIyrC
3YkBEDHwfEx+wskrHIRhyt6q9yqFMMlyfUdCHZDRSDJ0if4lGHpR5QRBNGPGbl3wWR4KOLCjEuO6
q1ayHC/Q3ON1cIL11N1AWki2G5L4omyI6YY6f/T+9hOnTsb5pxElOKIHkUjOUTKMWjQs41q8PP9i
47dZ/oIcUecm2dzaX0AMFh2x2HDsjvXrjuZ1Q2/LJZEb2WyA5f1Sb4jIf2aP5TfYedYQAsKGcgp0
U9N5AD6O9DzYwxVqx5Wh6g39+HMBu6A8/3BOPK8Tu/dAtbOn+/k96wASA8gRu3Mql2TZazlF2Nw4
NoUD7EP4hLhSm9hWq7kM2bSXrrFYggCU+1u9U7WTWkDRITRYNLMQH9E1DznX7u8y0mWAcEq15Y3e
p0Xv1BlaXCZ2uFgrr/SMlLYKnJ0jpyQc77mYRi6CUkOvGawcqysglcv90Q52rwnEz7x66WXJSlFF
+ldoB0/697I/AydlbFG307r/D4BtP9gC1mcCUMqgh3V5TQaZlk15wVk9dZihkMzwqD+OVzlblvnw
09cvS5doUl7LBNOSs9I/u+KZRWq/ekIETECUg17b0L2H2b6yIIRRNFJ903+mDsP4Mhucs1Pypvto
Q8QzTAOy/SS+zg0NEx+MapDxbI/xG/4QCetSaF17Oe1NJeM36jtY5YYfP4WD00382KcFDbvjI0T/
9w7wpCYluZ10oFYkcQYAfQXMMwscPaQcZ1EjujlRgU/dK9qagEU/ryG8iJeWtTOWEY6MrUknRK/Q
oDm/fp936xMs8pxFPajtD/RffWEFb/Vz1aYkhKXUWa6BKHohdkNkn62m/QndzbE6cMGn7+OGnkWJ
j46Na+l6UJnJvzU0ujeH/hsprKsCfk/jn0NyIZxMn5whpxu0C+GZfuqGnUBOKoT5+9k6Tojgqznx
DnymMo4g7pdtdp6SFv/sztLCcYlgUdDFkaGzxy3/yi+r8CP921dYpNZcTENP19S6BSZasSMS1z0C
xqlA59NJPn34qwyJCjyT/CQwN3jKFBbkdC1osuUnzvBXBAsGO1KCWaw9egp9kkb4ibzgL8ckIwaX
CgWkfEU3nuVz0ZlCh3ROutEtt3+L2ysxHFzmWs05fmuYxdvMwUxTafyVEORSzIPQa5kX6irkMMhM
7UgB6bySJds0Kr6EeCORuALJhBWkuF4MxPHOYjnHj6aLsKcpmMaKH2G0wPV35uZyXJ/LLzwbCQco
qV/Zxy6i+wcrkk0PaKTcx6xoCxgKI2Taven0wPdJaZ3tMXuh3a6zVJls1qWumXH93cAfUtzvu9gb
ufNTcc7AbSqTIcHkMT8dfzvT1fczFJ1d05IHLO2ayNRBNFakFHJIELVYMJQ4uO5Y6ykB5yw+YQdz
rVDcvTsRX4yieDSQIpLNgYtpwm8SbgffvgZl1DOJyrUtT3XNnSflnVNwYrQ8CxQ6ux51CwkpbOxd
mNs4twg/LhvoBEwl6++hLQqQipz3LeaFi8WpfHSGQgithw6mcXcwh/DHNZSCmLA8/RPxkYP8lAKx
YvqrFw4r/n29GLIX79352+NfbliLeon+kSI4WMagxWzYaM3JJkheZqVLDGKfDFzXCAecI4F3MfBy
MPCL2y7FNnborHicZf0xsHJNHD+bgFF1yACU2f0QYR+WUW79IPsvF4Wh4ObVVfone3Bs9UkFujg2
CYhfheOYXLtfG5ZCeWXFPMm6DcQUTZVqRIilaLMdOFxOpa2H+YB5ldCGQj6dma19eDdBcKaegnGc
VGBlSCjEth2zt0EXHBMxMFbBzBP63s/iCYo8DV11cuhaMaonALvyqmk9C1qK9RALrh+QfDH1U9hl
Orbi95UE2OYngsFpoqFSZVWEKaY1gFBrxClhRX25y14hxoLHuQ7XXH85RZxe5CMoTSV3/FoFSgIt
57j5YEP431klQWVad6QDvgepgTbiX0wol+kef+QPjS9IWNoqqeVuFQI6a1TipC9dSHbn9/aDG0aq
85RMxoSH+8hrSDfyCBdYEMgQ1hBR+klHfPD0ilayF6Q/TfZLvONqoTcCJmRxk0NUcf/hhBe6/9xZ
bkXE7Rhwn3X0wJDs9/xzdZWux9LCf5cQu05N0QP7uto+dnOk/7AoqsKdPEgA3mJRyDn3fSbku52S
O4ToC8RIvkXnUhl0LmS+fOXrgE5zLOUDdUM6KZ9FEbZ9Oqv9FR35TZOjh83gipesJAJd7gxEhEs5
Lc0rGQLW5KifjJzU8jVEB+S15k8fYxDTioJH2t8hJlNtzrr3rHHhNsfhqM83RCmckMYvaK6o6c+F
TpVgqn3iieslHLP0VbM+kwBlvCsf7niwx2q9Cr4UeqMf9jEJfJg0boEva9swSbvd4rwsw0/cujTW
sbaRx/XVXiXBIY7DLHgIuUjbc/okq+iqoQmc+cinaNfrVX4ghjpYTya/mEBciytN4KCCpubf7opv
aU9/pm1yV5K5xTsOYqiLQgXAkGO3PzlDv8SezipcgyUYqeCCWmOzxRUEEQA2EhlPc2voUQqqW5Tn
YoUfC3AmY5F6Fq0N81vsMKYZKro9HJgFQb91vhm2lqdPcPm+Re1oGuPQXlVEbQueq3EW4DSVBR8d
motUflHmQl6vg43kAp+gRFHadwbZZVXfZLvUXlCTnnr9nqdyHQqED7Xh5WTzFs5oU9IGyKNBCiH+
hVuIM7dGW9owuFDH6rJqCfrdEt07Ws9OA0db9317S5TdZr97Gl4s+QniaFKbUhDhI6voGOdB54An
vEGOAWtnNxWoQ3O6GkbZZaEe7oYVzl9ENz5K2d7MnQzT7Pq7JrNFKLjs3TPdFeezFk3jPxtIOoLp
gnU0OSZRr4wGbSmqspbt27NLlQEgYVyDJNK+fNv5wNtq7cTkmpqSeIqECA4VhMMQH1X69viiq39r
hy1qgSo5CDIwdvOo8giMjpknckZn/MkCVkxp1oGblgnu6INwBpBNnfxi6HkiQ8UD08p5FupiknT0
O17YSq575BODHlOIrQfnegCqSOjo+ecwpAuHWhLQE0kT49ZPnz8ybUJDLF2yb6jdzmch0QV6aAVy
KKuoL/a/ykKTXx2Is0Xs4+iB7ZCNYonGE77xCHYTwIo2AVKojTwQgBwgT37XfWZ9ooSqd0LRKvrH
mCw0EoDNLF0MErbQPJ7sU3ovOqh9HIJdziEbBNzQAsE7inWOZNftNQR+iWSIl7PL12mC10jbIQqo
k78+DXLHvGbjZo7FUaJYE4bBeK9jXgl6sgawIYXI0cj7yhwr8jvXn8Zju+HyuR2+iqj/pvtM51Bm
KIRwm5I9T908ona+wnhs0r+sNQuGNv7T0ex61yKml/tKXTnw5wh55+owCqi1JzETUbNzfPyAGHGy
E1XdrttcJgXmUWmASWP6Le/vtLQGHKVFYn2A2p68fO+l1bB3mgwK/IG0XPJ4Ea8OlX+S9SIIM7dC
VEoy79HmKJw9YDhGlhDenw5Htc/RgR+NFFXHlLi0ws40RhYlCXZn0H2VYdikjelTPP9QH57MV4M6
A6Xzo1yErbQPyIam+Qt4kKrCJDrOlHmwMMMuKP+p1Qi4NJKvwQyqR1J6RHCVvN0wKEH6PlfGZfni
Pt8UXXZN/LbM7WVrsYdRT8alxPR1M5fgKAx4XKzWcVZSokWDvwYK9GeKSdpsH+4jjtCex6lZ1iHv
3ET+4B3WA9g+hHcT5DceQJjFQ2EDnCCfoRwy2RFESTflnXMM8z4pD/z2kvzYPVN07ovzSh92f3xF
3DLaKOo+VO5EcoOCb7teNh9WxZGG+MkKtZNewIdSwwYtI/gDvPyHz3XxXeg/+mZA1D6hYYJzkRcq
9/tuf6nm0IFikkyiIwsXF98qFFgX4PWcxegTUaGPRDcQfGz9n4F0aO9K2GiKWZXORUyPJrZINGRm
6aMhZ8vbUYD4mW1YLXJNHNycVIhyOA80Exv8jonVGICwUbtSSCP0/q68H7yoTF2hwLe0OhJTJ4qm
YxN0mFNF1BjuhDQKc9LaWe1sEiz1oK6xyL303CJNRGYrkNnz7eEiTwziaKbqS1J1dVN1esxCiC2M
vJ4drOIgusP3fmjlz96WM6FvUPB7J8VzvNii20krofcqDWyp1j0XApBS9tkSwH3xO1bOjSAK7lp5
V/oASbVecGXNAk9eXxAwV3dfEKJcyL/dv0lXAtE07yK/YMzCCrvle1HgrS4e6tjCyDZAD5HWPz+w
BpPrL7UlCYsgJFWGJGyJ4LhaXfbtlUx4sEGuf+s1HmeLRtXb5+sDaHpPxDNEx28gJf21mNdONtT4
LidKQ0J6mDQLPQUjArU65xSaszHLa5idT6EYuzce1ZR66p7lJF0jn6UX7Ibme2Bdnxob5jNjqsPT
jYJGQiPLzaty8Q6lDnS5V6BK5JZvq9Ff3YCT8/G17Wf3/Uc8o0KDFXn04b3KDDtJhwdlScEDciq1
jq+IA0JhFWRep56qVajcqTyE0BzNg06gz5dTa7D6oT6Os890KS4GRN9kuVV4U/jnLIk4Absb0OWZ
rQMNnnbmbOW7YusTcaRn8JhTG2otg30Yi8dwsUXa8/wDZyx3buD3OXQE6yQNTu0oQWcL+IsqufOI
ObsPvchB5M2V0J2RBxr6+BDKi9RatZc5oi3WzVG8PIFS6/iIf954emqDqugC+0Flva0mssKtRyic
ayGkiHZj+zQzmxVkDoYXRah9w30pXfsM9kb/SjmTPhWigbZ5nXu4D2yWEK0JzsXHr2NKspriOnq0
bUWHbOzJ5ZkJBsgmLBU9NhqvIZ66kj3n1yPCV+6CoGs8Kre0469Yq3c4CM0fRzcFyMsGqvmmsexy
7LQA2f9ycFkEMrrIeTlhpElsEZOurBqJqJ5ctRtaAZVDYWPUV1rBlhLhD+lu2uVn+mOwiMdIg2Rx
Ng8/WyXp5aEoTFELk4rf66cPpofvqKycJNaDR1E8VfH6SrpPdm+sj7myiev4+nvTYxoeB8umtPsT
RIrGpz+2NHqORtkW8r6+GaoUpb0EOx7oxp2biCFGj+hJsDSUdiPyOnJvYxycsCBHGhZSRJq8D+9D
KJ8oIzTyHyRKYdX+nl/nMikoaMHDsMevI+SUdX4l5uLaybtzRYggma2Ts+oRijenQdGVyuSCMqwX
RpHXH1loDj2UekJcoK3PKPr2PeI8L6Tg/1dvo2sYXQPdHcSrGphSmk+y2xCvWTpNGKe0ombnKsSZ
nkFt4XCyA6zxv0bJ8WHuRvvGiuOjM08PZcN/A9NxzKN43pf1JKdhn9JR8c1cNxrm3xI2iySIxfVf
3OHRvT6dpAZsd+tYyFyfJjrFjWbNqEtZmwAAvGkNo2+7OaawBKGohbirODC2Nv2dJMaB81R0NgY1
6dFag9z3+ZuKs2vPHHfKScAyVWyqJ3UYocstfEvmJZW2GDyJJPwTaj4gw+5Jftm1m4KRoqEihaMB
hrGdrRXxF4ljQJ4EnjbkJiieeda+KofQXBjhLOM3dXOlY9niWog2f7Gp3ggAUWNSQhg2Udg5UqP8
9204aONGbyMfiysg6BgvSD6zHxMvwvtgEdJ5hNTWiHjwQjD7QSx6BpsYKOVaNMYNJBXduJMSS/sv
cYyW5hFW5JvOoNRH2mXjsW1IPnLmBjYscVe7deLEp0HTYm1+l0/XzHVSVJECEp3OaLy1IiK0Rdor
2rHq1NpyKLi210+BozSQhzOO1f4A5YxcgW5vTwPgPXJwE1iZqGQxNsCqwVf+spmArkBx4D9Ljrfu
zXcKy/+UT2dalpSNlBmkQBJNlIGQqyeQNUrmO570bwpJ8IT/Uv9WlEnRHEPbOeEn1Lm4XaU28IeG
/obuNAZdDAV8ZLFAps7dqHmZy3g6m5MMMquKIV6jvJeevQ3aHdbCgd+tT8e6AFGb2/EsR6NPOUAY
0+dc0tK63uBjnkxv6hUDs7Xrljd/io2HWUbgy2U95KSle0jFKx4wrqe7/xZ/EceoiPtkamQziouP
wdwgRXMNINYAJ200nJGw/olp6ZWBJZa2E5rjnS1VRyPzaswCRgZ/yKgr6+dnoZh/BdVfAM10+YOm
9oBUka2bKUCPYOa8gZZU4ImW/w8auQsQND6JedaS5t50EtxhyQj/AHH8+OArDLY6gNIlEb2jsuUk
1/08LPyaOzxS4V7GgffPhFFqWZ8t0yxn/0ahHdKqecj+OFyG31eqVWd9ViaRMQjarQt6T0NwZ8sy
j5P3NFc7T1RQFnUNVpaGqeFiAOo8Gbxk/+pgeVLdQdhX2sp5WRJrnTYx6jEQ3IUWtJ+boRn1RnZx
JMo591J/xmOPKfU0OHVochQ3pIh8KmGbju+M6v38QDXKauyVY0YgVnoWB5StpDuULceI2mZznqGV
8dL/eTnwVJniYF8lBI0BWFyjkeH/CuU/Pg5lFHRI+RDAcGPir0bRHrKTnB0XqLKvfs9OSgrNtBGj
8sQ9WWZJr3WHzWE92MBhqfBSZAxdifGwbWCUGmWnz3ibVw/uhqgrmSeJKSY7JAFb46sPqZ0B60Qo
ir1YB5Iai4f/s6eRW3gDzIS3Y1ThyxTToiX0hZ2qLkn4Y0OUzLmwDDr4OIfhX4leGts01n08OZA5
CMCOLdBj209eg903vGFW9KSTlRuY+EZ2EiSVAsAHWH4HjVXD+baWb0fyWnFf3eUleUN+RqrQcdvt
NqwuK6vhhpMtT/2rn2Hp9ICxJ46S6Z/N8ZDlfhQjKh3Z48nI7bRAF/RqHvO+yf9VPVPfOUflgpV6
A+7X3U2QvyktZv5q5j+B+4GdV80azr1+nsbJ/8Ao3MELjM0UU64dIaBkiqdSSxPptyfMT+Zr6D/J
3pcOZgvVxKF3dkvCeC9QMadwgD0XBGrRJL2fC7OoC1LH5UP51qUGIVogv7PqF1xXDCs5dGRMbMcV
F0iOvE+7nxhx6u181JKjA9zpps/FZlyRdWT0KjLW1TY+ECFaqzVzzoujxU0wNQPONUVHa05E1P8L
aINLPsmuG+fGO9JNJ9/I7TJiS8tluSQlTB3CYnbLMurLfVd4KNBDPc+Z9v4C9CeKboK/xMGNaONM
vrAMKmhELXs+14Wy5YmP6wQZVzu8XJFkejs9eCF05G/w8pcpUSrh9tCw7lDbdMGqsP74E110Irpu
gRZmHkAVfOVHgSjLcXTzx7cHtuunGkfAkSWS3VgbPWM+H16X78GT2BIqXgEYOO0J1+LLF/cWi+q/
CXScZdKAPyN1g2Frwpk5arBOR2CDtzUlLxy8jAV1RewIjS3w1omUQMYuZVryTz2XSAzt0s9VuaY2
zb9A3SIXjtwzBheVxCsjKT0dieXb2pjhAZVkNepLKaeLxu6IkDd5My8qeO4d/s3u83I1Jp1op1FW
XwiYN65RRl9e0lkS1ULbzk+sWQVwuj/ij+OD4UUgB4p8L+zQ2ZOOmBMYbTmXl0DwdLNOcp+7Wi1s
X0OZC0vXZ1llrL3So/OybcVlxpjS7q24BtJyZQCNt6JdFJRcZ19o9+SsBPYNMAv6/M5YOP1RDzM/
AW9jynHbNrrv8rpE+F0fUHG0yQbGbP4CyTyUNnLsmTIpP3NTf4vRTYOYA2HF6VAi4aec9sOsqMtl
jTLSKCJsHueVfjHdIcWy4u0rnJ1WR6T5e262MoNXSVv5Apxi9H+l+r1EoiFOjnAdaGwJeASoOmG6
WDApNao9jqYzAreM1E1GDiq1s9Qiv9COpk7EK5qub1qcW0sJRuQDcat61vFI6P13lQG16yj/hJ0g
v6aGcAhC4gMZfxHh7IELxkjR1+vFsADHD390Y6UYeyIAqWJ9Y5eonta4qhKMc8qXYMgSEFmNCCk4
AdwdurhV5LsADMgFiLte+bOLjmTGka6UnMwpcUvW1tmnbhkptyL79/qLD3TJwVze+sjhNEZXisnD
HjG6aibC1Y+U6rtRYqfQJM2FAnTCa0LcU3hlPy6DKcisfk+c3poosBph420CzHMJ991BX1qChXJ9
4qIiS4Jk/03YOubKfcBuTsJEKkwatSE4rYSmO+ln7uj9u9gdxVmK8+WoouXFSgW0nDCzFwTP4v0j
uWLOFZvUgInkyCWIbU+VlCeqILll1JCnK6IT6w+AYbNk5x12xesMhLVPbUsNalOSaajX/YJuXHcl
QswNVmVyVziPymsjbUEm5nEmZj6XsPGmxcNXO4ViY+DHlihNuLgKKkktyA8GsLnj5X8HbihQN7CQ
WuEjHtw8HVOkyizEhn/mbg37W9uCAXob2KCFbmvmiDvy2vq6nWt/1M0oce2a4s0Il8RKp5QV3KPB
gUp9Vfwr+wb+Tka7X7OS9XEP/MfF4ph1O9HXXOm5bQpBazcxsOQd9+akKv8HV/BSqz7jc7fxB3Ea
ligJmdJuqZAx/4i2KejePYtbYW9CwEz8Au4HXr4u1gE57YaBl47plnw1g8QCtinQOYgaeTjVEZJS
FvP3PRMrTXBALcE0/+a98qxTBmgt86earWT0Yeva6y/RVmjNjUo3odRfFed2GoBao8D3RN1UFavL
v7axeb7AGcy9NE0fXO7ep0A7k1LnnBlEm99op87KJ4E6u74hDEqI+82BmNU/6S3l4DSQrFVpw/0+
Um2KKq2Er6V5IhCc9rpvUIk8XNUEHt71AzY8aIE+K+NnOEpfS9WCINWeu2rocKNbMRZG/IY39vxn
VsSuxw4gXeSwJQ/8Lc3VpbMzbh8tuQ/xGNQqRyJxuLD1fO8oYKOwrKE2Mbp2sKusvNz60YyAIMdj
2xhv3pKAZPqExNsmClb00aPaRMhJsgnz/N5Rhlwicvw/Q1PgWbsD/jGbfvRt/qQGxWP2hgrH5kAl
4N1N4PDNOXybaqCbE3PGOCcz49UooRwh8ZNN140zt7SKbSYfz0bl60AW1+Wlaopyt+4vtoy9Qnzs
WfHvdm+oGPJoBY7WrJTO0eHNf+xejIITIY9yznswsy1sR9NK+byA/3KuoaxQX3NBCmKXdYtGFOyX
dY/9jWh5RDGgF84QTCKM1NwvVC5sNApHs/b7+Hpabzfy57vF9QmHhxf34GCpnLLTgfxIfPDj5Yzh
BpnSokgP2/CR0OtkiZ2ioU4BEfv/qz4NgK36sl5zZfqAMGZrQsUloMOlwPictw3msR848ugju03d
dFW5E4NqEJrYdIJLQ97/SLqkJJjxAJ3MsFBtn3oZUnDPifwQTPp2Nqw8VRWZLPP5qshSPh8obssP
oWmmUrq3KZt8RUZa2vKOw7c7hxXuYjQ89MjdFQ1Qcoq+m4MPuowBYS9J5cfvWttZbkJ/jE6pAl6J
blecYwEfvEe3deuqZIraHVBXTEW9LA9r8uKKLXeU2yrtOTi15uOdr/7O0W8hmQAUmlrwloxbnF4o
SZpTPm1bbCIhvM95Cmz7U396U9Q6zkEr7Fn+vhkDUHhbZp0Gpw1W9JlDzYgNaPpbi7fszxlS2Jvi
BoiGDwLEb9clLqVjWb1SPL9eDtg2KOSGfhkZeAQF7wP36TFr1fHPUqvzz6Ew1kFI4IIClVzlykdx
XgpcsyfDpEhMsu2+hzj6cHj/rJ9y9TDwPu6OR4aynGb/LQ5OIk0oM4upuxZ6xcN2qa3aBhL1iyQZ
2XDmGUuKiITlB1UPwfL2ZoBFkyoumBRzlk6FEmABgMAdh8UURioUndRcEIOPZdoKRf2UR2FKISt/
KmUEeaiyaiI1nBGZObENTo2lDF++lej4dBr7uaC3kDjVtDk5Gnh/ZwqLzhj+t3qT0TswUbfk/NOC
xCnSmRukCjyOByk/8PKo7LIQOqLKU+KCPnoHOxwUfB5d3JyI1JZ54hS+nUUp0z6HYXDM25bTJZ0K
8+TPhWYwICoArKhkaaZDtlQORdfdNhJ3UNK0Cddaf2XxFnAHYwPnInfDysgG0lMbg3sjqEPk+Mvt
ZQ4iZQ9xIqtBycS4O5i5voacKns0lrnu94R3DmL/2FPphIAoU6kfRHLFVo+8HhVVmMwy+KsDY4A+
Bxh5KPpuR9qG3IjDcuW7/hWQj0WyyPmjkNH+YHduoS7qyLjHAW2g9+4yyH5KSu3Xc8Mx+SIVJBW7
OKyOrhUSFns2iXWGyr4Yurp+UccGEpg4e+Eobk/n7FOmtzYUq7RBIQAz3/QlgEH8XQs6cJVqHEmx
XjOkrZ9bXUtzXarNyrMXQSH8jzmVjlPLK82j2EvV8MN3K+xc1JSHy61VdHNp9wazC5NO8CFW1iVC
DUshBidgeGj/nWjuBDrVFumQTzSf8p0Q0ognK4Tr/AmvuhxPj8hezlcyiuuLQUgMMTqMmhE63xDK
szi6aZkXuLhmbW6Uf0PArfvanZXjut8Btv0S2i3cFZkYvJGAuLPpnN6x24x1AENQGZT6h3CGWX5/
6rq9Tvs7Zfo1WuM9mqWvIzozmxT3V7INEX28WUklNBEqXpD9ZyKAw3n1y/je1X0VGIjStoZ+cOiU
p8XcShMdt69hP3KgGs+FtwVsMA+5UG3z3gB1qqPabnki/vfG3ogYeq3hrVtQ/+nJEUeYeihVnef9
E72yuvX1FMKtRRpfueGMxDnpxDdX9vMrQRrgJF1WPJoyV/uTERjgU63JqS6SzXGjF9/uQzO9bylg
ux0Yo07FStZUl4zO4/ewbxkpw46hRotIgdPC54RYqsp5h5GDGx8F1dZOt+57E80d/SJ/zFsfNe6U
AQgHhGDkUE8uoylu5UthvMBFiMC0MC/eMuh639S5VIBbxnQdNTCyABW3Rb9b+HmPEImVlTOoZy7T
9NWLNT22HJxM5ZsVk+Ff0Nbt3MjEeQa0YZx2b2F1XVDNxSq22j1RMTFJF2MIWDGXn37DSLbH1MGW
ohcWIw0GL9GqB4glk9ZwViIwGybOZC6ztR8WbxqzXJJ1FgyVH36kw9RUw9Idz9rViBXP3OloI7oG
yLXYuwxYQ4nhkPhHhhXh0E2qqUIKbiEl0tpxCcOLVNI3+mvqmpnXhzBz6lgVm/hT5H9RjNPMK9aY
g2IqqfaWABeFDZfM8S5t7rY3ES/VzKL6Z7lVbpVeaJcHEZjokE+V119iq/0fbJQJQZd573Xadmrz
by4YG6hffftcA0LXl199F9EJimGlAgLh7PZc6JDUYotfcFTraOvLKCHzDOjk1Ls10OdMAgO5oHA8
x6gHpRBswXUAsCOGK9U+ROHxE88sWvxBuDbDXlrGLk6gLiRlNk3GKx504VcUhBaamBDRyFNVTl+x
Ryp5UV5tzn7rqC7eFjeveuHnsNCTD4xvPohVOOfrG8Bulgbsc+t0a3H5xGJq2q+EMi0U0ktDtvB2
AZE5kvexGFUh09zF8L60IkMWRNTiGUrQKSLdFJNRWdHVFZvlUTZiihuCJ/CnIOuEjCe3BTW0sRKq
WUAybiryHotPNtzpLvyeC7XL6pFqdZsGsNL7QCbO1CXEW4kUnPAHjaNQGTgZM7a0lAgHfuWkhetp
miS99YlgVmPM/WXAgDiT77/3HuLBP0T/aAVUsigqIGd7bEcs+g4CUBIThrdn0nIdH+JhgV+9qZ+N
r5BB2Ts5Vunb1RfB1ZO/dGi5kuuXx7GVr/br04cqzonQ9yvxfDMmWrERnMx8GOLdLHuW2c0QzS9T
RxLWEs5MFJE9oEkEovoB7pbCbCzCuRetqrjtO8WctpEi6cOdJcpqDm9ZZBfa+tkDyCcDZty1O6N3
kVp7u3crVtpJd09fCeHm7nJSLZfLY73PZctJpnllrmPEPT9zzYsjB5c+HD0tRSMJDl+EiE4kwrP0
NCVNyf5ONw2z1KNqfNNOBaKnnqO8Arqse5FNdU9ntAiTZdAPyeyXqhe+ExHQwHNkScpVL9+wFNS7
NBfPHCgZ68ArEATSMeVVn0O7MEy6l49vJ+H692qLq/9cRJvLNRlAhe544Jdt80PP0PUUpd+YPbPY
GnBF07k7AvonV5LY3BUiPCaifoPv60p5DmOtGdsibO5OBKSF70VEq84+30eKvKbTfOEA7SG5tmhR
+HWnK1kZbtUjFH+koWa8Xu4PQyBVifklvzXTdxexmmIF8Wcpvq2xe6XglQZpnVF//Ub0gv06iIvQ
WxviVbgvtnqZqIHjcYmDKbbAQlDLIBlQ0A5iUTxfonWy81pDSTNFb+K6uuDKL9td/tsBik3xTsfw
+kMwuelwOAfHu1G2MMBrIR5gOostTqVtDuSYYAd99UAU3JYnXXXm4soDgR6DVtEGDnMzSKUXUS5n
zWeuF19Pg4oDXn12yFtAO8zxCHTR0MW4CLaHIQBx+lgiXzg4UFEV3YPs1gQzGmdVzQR6jwW5BZYC
Ho5FUjItScHpZj47tDiiV2aKSPu+Y++CJ0LnXYBf2iILrq9bEvdvtvhmJ2nwTn1/COzFhhg38YHg
XZDkKFS3R1j4a3kuxC07KkPeZPk6aRS1KlfADpBZjO9bqB6ng3qhsDJQILVc5G4CuncxOgj/FSLV
cjn7Ct7oEqkRG2DA7luaE9FfuUQe04A+0rURAQ7fvY8SDnBxvXMn6Vg6iW+edia+ArHLYfmM8Sav
rii1sKlpzukf39+KGgZc2fgd190LdAFF8+6ZHcZ7GnmlhfLpfjbPLta5y5wkDxSdDzzeVvWtG/iZ
Fy0Lj+itLkfib/t702ASOjPYjROlBc8Mn3rLXP5NPyAPjjlB1UPnVefP2q4bxfF/RrjQr4vjRFBs
zK/Jf/brQgk5ltBN/gneTaVmObUYbGWa91pRsbOYyShhBY3cxTkt63bTsLxzIGl50wTe2+OiarVI
Dh9iG4V2V06O+1R9NdXitX62eqAQnu1XR3g3M3XNtKPqogqyiN6bj0jWzH/FNp9ZSmMASuRZ7klt
Nf/wEaXzL8EoeRf3BA454WpIuI2P8IqdtulkM/g7BZ1fYIojafL03MV7ExDogyBaSgvTLyBjrBhj
2XZse7iFeN30rdtl4RxNicTfECVRzAum36SIvxSVSjbqvz1mgtFSjxiOnpj6kHvkmshU0e+Hh58n
eF2bCDTvkViSiZwD6FSVLdodMCB6rQoJYXEV40hkyujVSnGrfdIWm5FKiW7KU7ycQ6uxkaL129Fk
Vi/YEttWJCs9RBSURx1+2/B0Wg8MP6tiPepYKQQgypr3yt+SCIu9d77cqYNA5huwLup3x71ONjAz
XHDTOURyTI23p1Et15nDG2AZ234ENTOQEnStEv5GBgepxDQA1t1fOmvv96031m99qwYeyCN0T4jR
OivXiVW47SlyYQJpgMMjynIaz6cjZfTMKHQMjQKVllj9eN6pYgOcgcxuuSbSDmYjHx7f/JSIM2FK
PIc7SabX8AMnBD9wWgT6aPGQYtyZY5MHTVY8vWiQKZb+/PZZEyKKoaeQ3htLGENyfjMOwz+ipUNG
dCbZ0NgufiZJnu3GeKwQxtcmIsobaOQ53vwlQB7o0iPp5Zqh6EbuQ+lwE2288jaYqZgKPkVE0JYC
+6ocE3MiDukTQ62dK+/ZHolx2ROYZeKkJqimD0e8fRb6tCIYU59PHaFTfHdc+bREIg99UGg3VYc4
sjEfqro4bMDYZxIrNrXzj2CrnxF8fyv2F6aY6iDnrrLo41e+EocRZdK7qfnWNP92gYbEeAINGloh
F8ZAI2UjCZl2NRfzOw5m8V1COZZw4ZU1ZfuZ2KIyASS8xQogY9pmeHREwJ70ky1GbPlMj1OySian
SHenLrulkPvrN1a85NASDnexHsLEhzudS5qxzZcSOnJoLJN1yBgS9ip6c+Xc58V3Q1L7jFljdp+s
NB6qB4zGjD6Y4OwhVucXuVJ9em3kxXpfakFhiTS5L16+aZcINJ+/M5lb/LJ2fMWNsD69tN62KcYO
NOI4hE2XMKXrdLTa81uHO5OSvyoNceAX3q7siFzdpU1f8GQSI46W/Fv5t8DCbNGDu3ZQicJD965P
TdGrO2qGsZ6IT3hoJ2sOzlDkANFgVN6Eya3T8Qiut+P9RaHqcB7oet2OwH6aeFkdxB49DfDVfcFy
xdGmhQMS3BXcgQqdyR6QJnxoSTKWVI6DEOYo85MrrF1e4vySKuEbP+GhY93aeGtiWvHFXMiy/pRC
N5uYkB66EIwoaG72xMXrG73KkpWdFMSvBg5oYbX+5ibjTr1vWxRheQcXkSCHzljyhHEqbPN8pl28
3VKC1R8jRPNyKR4JGupuibTHbd/1KtaqKDf8dsqXifXXXoEyNI4WC6GPx460aiKWDlx/42VHgmpy
m/7QWffgcgLA/pShVOLPgUKLOn5g2SMe/cXE3LeHosQT5WRrMswDM+R/yj9e5LpAAn16f93GhQH9
QhoBdNjUzWms0MbLr01qgU4HIRagJrqxnZBJEfAwlsgbPdB3UMME6/sUYgrv+pRdzOEzoMvKAQfs
Y1IA8yusXuzzVXBXagJqDTHOvbc38drKJqgLsBsQ/5LgbKzfbZU44d2c88PXJODkW54/TXDMfjF8
qEBmfFOQTfdjzp4yT3m2nW2yyIqu+cMHKYenjwebewU0zLTes8S5YzErtRcnl4WchsHZlUcuSkDD
FGU+JHjFbQ7V3DiLAVtmHQvAm6q6cnpc8OpdIyCgoUnW+dUgOAN0U4vBydpC09iE0Q0yuvyutkHW
AaSI8LJmF10Ii3Qb2GiJoZauquAfXCqsIO6TcjEkAmv6ur9aBwrQIAAMQm7krCt4tfmkACCDriph
S0QJ0+ozq1rafLleqPl2Nx7zce98v3lSND/qPrIPqRcVGWnvUc9dIXGT93CeLdIFbdrKoC/JknFo
+ohqHf/gRaHDZjBGLdW0bWxIOItz8CshPAyMMnpjKrPbe+lAvIMNOzSLs8dCfGCvZCWQKbUt0Zw7
DCXNIahxSjVVlLWjk6GRdV2foUXSdacSOc6dTpxsDTxXC2X2Cg3DjuMbxGXtaRsFMYLGIKKC1N80
WWXm92sU1t4coLYFAU0CZdvPWIV6clGpBJ1f5Cnnss6Hj9V39X6ZlnkwMERtvcOWspvGKqLfMRXy
Xm5wGT2A/Wvi7k+Fqacm2D5Fot0zG/ngvzHefKnfwfTgkoH/WPrqaoeqpalm58sdyqGW0r/tlDfL
4bnArwaeRCNb1PAQShUO+aC4he1loeX97qT9r0vrdCKg9sam7sOz4vw6XRqcwGlegvz2AgcKbd7k
LfsVt61Gy1cK9I0NV+AQ2JMZ2UlCZ0PZUJ+icueemBCKIRBJJjTY8WAJrBZUvyILurgHAnB/pj/C
r5m2lFnjpd5+XbTTiOqo3IIHGp5SSrshBzCiS0TSfJ6/Vw+KgZNq05Lf9Pg5sl0cr10JITdv+iO5
zEo0vqiyQvm5i3etDHUiClLacRrTwN5LtpxvhHFdxp7mtuCjZBZkbeYZ5Hkzwxs+DhhpgwulnIxM
xY9UtMd1t/sLMQTPXQ75fKBdnfkTycgVhoz9Ehc9W3bIHZ/uTVbUjG0G4mjHjcLvIpVPjDPxuB65
3koBHdWNnFEfB5GMWO8DYmY1XDRyqm2L+kTPWmCGL1UaoGcyvf4ezJ1+Uvge5SNv+a6qn/8YTNh5
v9mZmZhOjI4LlOzSgG8+LZawDXf30TEMT8lLd7LbtqegIJezH4AZw01PuWGgCmKBs058N+4p2hS6
dHeooPuGgXYmxWyi64xpY5JaCpP14rha7GuRq+fHu/9qnXJsA1z4IiTD63+2oISUXjXMAx5wY04N
0Rr1LGNz4eoif7av2p8xhpb+a8CiNIH1RuMm9I+YiJF7H12XUHFRqjC7Ga+GqYt3AkIFvWINH1lm
FArGBtIEze2CZ1H3m8S5G6YstYtbQ3JLQ8fuF0RjoiG0i5mTH2gBOO9FvIUD3mmsXY+l+2q9EztU
NceG+hoOEcz4n7xT3JRu9LCuGAPoRD1HqgxVyJC+mcDl8brTHvGa3DYW576ND9kpkLqy4ZxBWIzI
bOzlc8SICj6ARawegGsIW3McVYxJifRgRQ+eMGVmZIpRNdz9kZwubi1dHfPCUjBnPrj4LXrnGbtw
FvU8ceIJpmJiiGg88ma5FmYnRoID5xu5EBMgFfwW7mRbanc2WGXjW1zUG1lCMkLR7F+hs19h9rwo
5emE4rEI3NhlqyHUphToTjfCtMtlizAUUzTzLyId/S8qaEkKIKrizBd0GGPkuWh3/tK49mUnuE2U
7zZltG+wvqLyFmxy0yfcqEFRgQVuKviIaM3IkzvclepRE/57semp9Sr4jellAyhiBBT42DVKwL8l
TVTqykiim29fhTLyIF2JRWggdqD8RsdMARri3zYz/+eWZ9GjRBthTvEek/ezY70TxZ5cRvw4VYQW
aecIS4uv4Wxw8yvvkB4PWNiwwjrPFSBUR61iMtNJNwL7GpWN3D8YDb9QZvp5bN9FNlE53LqlIJFm
IqR+Rrl1S18R14snYEPHWHQMCm7oLwZnG4QqYbqYdZFdvp86ef0+6zKECM/1lbpZKy6khZH33rmr
2elveInpvBCTwBMdhsLjC/FjPxqGX38+++lU5iBOfxJ3//wesELAXHrC0zZ9txLnCtnnhFkWlMvt
VmowygwH6oSZf3Zb/1lkhRQyb35FEXOlFHFB9Fx9Y881PKo/WVPhFQt6E+axb4gGXWABXt6QMSH+
FFh+gapxBUkTLPD2Y6q7PELqKVAK6/PwcF7aDEmPhlE1qsW962icfdrMDkwFEstOw+0DOoKB3Sl3
pYB5E7BgCqZt8+dx5n6ESX3bWsdmWfN27/WevX/J/AkY8P+6MRk4q+qTSoK1HP0j0oid/QHLivMx
7BsHJiNqU/TYEnB89qzpzsHT4pqg4j/Hg2tH+H8ZtaxjstH7wHvV54bCFoKgJ6xzf0YqhFfiht5j
q5/1beBX/kgYQVj7cyFpGFNyjUaNUrA1itF8GmDV/32791oVPHJqZRta6GSHGJSLbVFnZR6GOi44
Py9dIia1/zWNtdyKxdN+2SmhKvpaJpWUSiZt0u0HTVeYftSkGne78GIrMghw23pzrWjJEqMzihtD
GMJSIXdEznUQW/JEu2uJyau9KfRA6FOCVt7XVlrf9Pg13MnnAc4v0Dlp8iXYjFCA6Ah1Yi+IRJwq
MbUQibA07t9IxxZlH98bZGkcHi2QL7NGUNEZoKv8BWOgmyX4Sv6qqwkj+EKTvJInkbJnGfGIZE3Q
gm8/kWKFeHLAbjT6Ojc3rxo/TlHHB7JYjVCV2uEj9ZS2YwbgDVkHvkeDPlOf/Ajh9hdAkkSC7zsN
viWncdzvDsWBkPf2baysNLgh1QN4drCjflA9CjJm9iPSMUxqNX56D0vDrL8hAK03G/26B/9z22Lq
sIrF6Ri7nEJq4nnMxSya3xcI8waXHlqLV32SVYWvdsYnCeE5K+yq1CbcJH7VubyBjqI8gbQEmR2J
vp9sRdsNBjNrjWASKM+KnvdLfcgUqA6qgx9jV8voIfxckNGmvqLDmRrOcC5a35/hKaKIWJ0BvbWB
HJbffoZVUQGdl7pIdM4b5vkZINezaF3kmi7RCwjtoSTZUuLdA3UBmJn8Lur00J7bkOp24AkiWp5m
FBMG07yp2E4VNcIupEa0If0uoab2A4AnbzZXpR5Ma03V/RrYK/2HIL6V463v8sD5L5vKFsMC7xp0
/u+QxS3VV/LXdTD+Olk7xdRa91K9l+WZrNg0dQZmJWRAIwq6GbHt2PJI650YvGbgTxCCrrKIzVO2
5qfdQYoG7zvZH4Q9PrJrLy9CvwxRu6pxH4k568t6ammVFfthqRokfKVRvlLweSirtbdT1FA3vId+
yGYCU+BJvXUBXMJ7IyJik5E/zM286VAIenoORPuk6XECqyThjit3VxV9kUl1ebn5ODFeGoQBZErd
r9Bwm2v/jKQBEfMi3ycH/MuVsv71Ef3VGaZ00cWXIiFPkkpfjwlNcF0jSNBXs7VYszqoTLHO6XMt
2RAy198N5UDd/B99vUhZBBGVEyY93VAZl2gnEn/jowIvJOHhHuhs7W0qKWBAKx0VfTcEAuv9e/xx
bwS3OuGNosv0nRlyl760800Y0/PAa32wDJyx/Lqp9OHPrh8IpzXKyv39CfyBpa+iGdY4IcJAd8Un
H/xfRp49a5LLcF2pQA8szB012KyroBW0ETCy1imU53Rnd3eh17CcsUQI6agXYU4upq5boySGZljM
MzKpIprL22skUY2MpFUTY/N6BXLYMh+iQX16fWn55Gyk71ByTuuVqbNXUn9MaxZTuXNIhPwzCyrh
Yf+yOH9CtQM97pceQ8J7xqNkttlbdlSD+UFVeA1IPyUTkPI0CM7F6UkfvH+nlMkpDgPg1Te/AVoW
foxv60dAEkyIQdfYGZA+EBQEpKPHX6pvY8dAgklqHosm6NlAERJzTV4sYrQmsMbyr7FMK+hiCfa8
1aNKRqHMdUz6WHXVAa8ViC8cDx45s64qGEhf2ZhBEJu+PPNaXNLxFTHC+I3HQpybN2ryhvMFOscx
zYqhmQ6Qgmsq2R2vFzZupECs0yOilAoiJpZoj1VZyfcnBNaicg1xVrMg68SYsugRvD4rbYlUXea2
2QeQmrQPqQaA10d6zJrzMoUAT4AAevyhqAWbQPugVl6MT6hXO+vpnXvizim/rHH1Bb6LtSUqaYIe
77ut95sL0S+YVE8Skqpy2B/nfuBDkAi2q06TOouJMdfMSqxX4M5AKoips+r/wPVF3lXKg7O8MVeJ
81Gh0Nq55YDPsgzjQvpRY1/xq9Cj+D2VLxzf/sq0uB7s7nKsiijw7pFwrucP2TigGu9THlNc3EX9
K8cDU09q9ea7hUIbTc+QxbnDaPdviPMXpi2AbCZYVljsByBxYShczfPbv5e0/8nLWkoqgT0g2yhj
aXqjaUZIN5SO49uwPZy/8dPpMBb4c6gTIrvz25ekxfkdRLB7ajgWQg2EIXM3I38Uzo/3BwdTVEab
U8gebGATRy7OLYlW0dPYgyQ2tO9Y42m6szyQQ3tLE7liVNeoi/ILSKysh0RluNmYJoCefeK4lSA5
JaPyXxtZOB5ASAcn3AZp7UJwFRx5VF7nV7A/Fc4zPKG1faPMN/8xenIviEoIXgkpREMHaKz31Fj6
ccFMi6ZnHmLgFQ9iGQQ1H0KLDr0KePdY4l/A2lEOvqtBbTK4Xed7QaRXda5Oyv/GU1PsIkzhAlQG
+QczZg+OifHpEuExUZfDEE6WA4kptX/+xLUm3FfNmUA5vAfQtAeORhLJ4rg3+hJ18dQ5mFQd6T6R
vDx+dXnUu2fZHYWRLTKIQAbz3xCkL7bRCcYA5KDfRQXGUd+RholHjg+GgaN7YLpnhytangAO9A82
DLz9DituP/xbv397HCigMpV1aJwQZVM/gfq7sSUiMfVr73t/8LxmZ2uFNqdjb8QOI8fTBEB9Uc9A
IepDDcOqq1ISeegOS2MX5ljvtRBDOjlSwMP7UZMNwNEmC0rNim3FcHH5bZ2lviqLwR4e8qETeyTd
Oreu9rkF5dfRqT4vP6ciWFaiDEywOoT49L/eRVD5IAAhkaDSWbdW0x0zMPP0wJBJUiWHKJgL4n/0
ey+XTNHf5+58MtqKG4XS7tiPZdEU/IQRMfw0mL98YwM4TCyTAgNrSk+Ftr0Chvaz0YUIHrWqy3CU
TeFcwS7KJAKl5+0WZvReggZWP9yXeiK5TztP1GUV1MVykxMW0oZmgodJPE8aqnlavQ7pz8gknibs
BL8QBhb7/1BFORTQnVWX6epwT9ufx7MqOPbQHCf+wwgeDw8MaEDGx6PNO5gOM5gR2FeTZaZJErWb
0Oga51oT+7djNsTgjldGGTsUPlpqEIxWt551OBvF3fIhqmiwYIT6PXtRHZwJXT6YorPbFQAOnSun
KaKTmmr1Sd7PspAVzxiDy99IdbSEzeBNbvbiLgkK0y3jbg4BXlsVnNcY1Rlq10Zl+2MFU4jDBHOb
2G+O5PlVKahVJKawvbBiNq7EHPrhtieZ2PSQxD2tEd8TWPHOKiVcOl+ZZBoljllv0nOEnnEeHW9U
oLDIR2L4TxJcYyjKEbn6H8Aa1y0L/inMi3a96TFiHovPxOe0czb9O+eCR6T/SFM1TNZWOo1CE7BT
67HCGU0CN21or0mNVqGhxJMHzhHTVXcPDmOztaL9W3gW3esi5BW+m4qSsB5BASusH1mUxuvtMv8W
MLGXZnXBbj3PpV2z1Y/uMutNuHYbZB7uTIOFYJBqX9Xg49mo3Xr3yvfUERfZfwXdD6fGlaiOE6w6
sd468PnF1ApQ+mrwaDORYGah52rTdga37s+UUT3oI94UC8gukm86n1F7lv63MGrTErJkpLZmu9oC
+fyt8nv5N6jMSAdz6iq+L+YIFA/lbiHGYkR8MKpLyZ30XLcOlSWGfJ0SnCGqoJOMM6pZnScceYA3
Ae0zvrN8sIIigHGhgr8RkNrYDPvKU8AyjBeyLn7ZNhOVrvUmZufpRTyGl1vf276+7WMAX67QRdzr
dsIDf9nliWPwsZmPLBbw/arRiXONzu3SuUpg0HlNcHcDtX803m1gybj/r/pUb74blo/woUC9Z9x7
jBFIXr2EUnzH49hyqpW+0+/UEUEXakdkz2bad+D+VkWsi5rhz6b2RkE8oRenwXCmhe9QUreyJlNk
caH+z0t+oUF/LbRRx9FtB0vEGd5KsvbKW6tUKjNfTqb5z1H6Vj82sELpKCMYFqN5+uEtafEKm8/3
5TYLXlov2n6zK/NfXWelzNirTYhmsWEch6Uohj4POIWj39P6nLtRecZoiltUxYEeraArMXMU9Ve3
XPID5ZDhU5xD2vsFE/wgvmp0Oc5f7ZLUnwt4vBcY09HyqwekGTB8ACFwf1gUE+l4ZfEH7Cc9xvHH
6DGKI/99EeGjMJRmMw8NurMiCyZK6spC95dDNgq1SqRmImQ//sfANSedek/l5q1plD0o2tsck11U
j6xOeHfSpHGIhYZeDUDd837vuAQco76fMmHK9q60J7WJKLRFo5i3y8Cq8klSxS0Kl0BVniufinFw
2Yqs4NVKuLxNmC2i3UoxqQptei7GlKGncxF+THQMqFRQKegkHEHI2tHxidM3JsShpeti782GehaZ
xA2wPO0RF5xLLHELX9VIC50vo2SLi5CjWTIF3249aguakPgtebwSq4PlnP4yf1EnlHE3DAcunrmX
iUCm0OkKXUBkG/zblqRSsT9oUOH3fWDXTpWajcWadDlhRSO01D1/FKtULBuUy9IOP0Qg7DrVWTSV
XoIv/v5VHSaT89noMS7JAe8ogHq8f5pIjs4N47MExfs1J/QCo2RPfke5pNS24TGQzq0hWAic8MkK
xd34xXHIIfDfUD/d7GVA/8KK0W1H9vo4pKRImTlmDhtSUEzriq51V7EYqRjgr1GLKwNXt49xzbj4
AaFivaYuq5BwIZ3ZdzGXEXDyUIIph4ru4QOc5s1tY2xoU9wKQZZN/fOb6Oa0Uudy2sQjapl0b5ez
7tTNAE7b26cUB+gyn3uP0eeRS4WzJ2b9+5LEW60oHnT5WvdFQpt45hzF3g/D6dDSVmMFKQE1MCb9
VZMtX7z1t1/c/eGEO9CAr2VSoW57RucfohfVSNnezJ8mIGPW7TkW7YtmFiLIPhuFt8aw4NVXoC3e
Xy7qfZIVG2livKnh3hJNntHBAZxw72CFTqb09lmRsL4MzN11FG/HEsCaCIUxoRCQUBmZNvcgXqZ/
K5WQJagMnHTyFNgHBh/tRcZj2MIeFdCiZeWdgn5TBiLB2l6CA8Ts+wXRbWAwT0kVrDQMhOXKoGHh
X6iD6KXm3mTuK2B5xs7045sloQKlLF46x6EfljQ3IlNoIl0KnMDsPpWDQ0yHw20turIDIYsNs1ui
njhvWcCJrB9BKBIX/MGZiO8AywUYvJQwrZOpIK2tU6prIsSpfFlwX0V8ZdX08Q8tWOxDsHWB987g
8A1sPZcxn5QKFqhqyzW+n1JP4JFamLNxO1hOS2pNdCkLuTFRx8ChdBakC6OO0XU8Z431XpOK9b5Q
oq1+4WatQ3NzmBBsQEyYkjeFsLSsCGLgP4pKVKhSdGuOyJnn1ynLr1R5orc57W2Xo+gJ6BXajHjr
c30uVxJsIBtyhDO4Q0UaVXQiCSUACSokyZQy+L39JITsyY75f7WOLW6tJ9j2ucbjeeZUBE8yZnZ7
HfbRmugfR8XaBWcjcH9PvHL6qbnKzaYFae2FZfaKwZfd+YnxbkG2BoQjl3JAk3GHbDCh1UWUlq2T
K6iw/dxYE7HuqgrSLmW4yhJCSKE7K1nUpgrNc3//udLvqNo9yQQfJUWVjpTELSGostTKYXA5ISog
UG44rO5spLQi4Lp/ZBqgcwtb1Jd/BwD1xGBEIDUcfRLlrYTeSGXRTSCZe5ZJTRtHdBPv9yKrDZ2k
dxDfkIsSw44oIFS+bgmNILqdBIt4nohkn5f7Kw7dHtjk3m+Cq6b4z4Hp8WPQ3z3Qb1+/ICfIK3az
0pbwdmfwtn/Paotv8heJaLnK6E93nu0F0MNFePw35jCPAv8n5ayH2Avnt313FZ4/5MCeUSAvKJG+
7crrtMG/bDrcgxcjE0bw7MThvt4tqLUyt4s9x4NYYD7OPjEXg5G74bsmN1I0LlZ4MbHx9Mwg7P58
PDDMk9fuwwn2MQcaPsN1c/Ysy5lrfuOx3/+RPoZSVvVkp4HRbTnGyGiDY0ceVOtddg4BmOToG+kf
KaIQS2ykFlf20fIXiQMuRH20x9AoFCnoqGaBVq+x0ELb3mbiBIVWurEH7zRSgdB/gunGT3bscNlc
KCYFrBzMIxBhPOPFTCdD/mHQ+8F6XqGWajvSBpsPoHeVf0Ybr/MdbONwlctw0zw/26dfy/ZwKIZf
fAO+i0fBRNiI6JnAqZ+WCATYp2AHTENTsBUP7sT9wnPx3f7Av/LxFKqy5vbPHw2jT14H8OEgPFsg
lE5XeH1U6X36flNxCIhzlN0xBUIW7Q05V22/ww/d6GQSaUJcfHbi+XNN0WvHKq7hO0JDLxwUab4W
1DAdN++UFX9MfbX1R81YCTmIuXrzt17Gc1EHYstbw93QrcDCClkU+/yGust9JhW4XmmdmwNQm1Ww
Pk4Zb47SlPs3Zv7PUFYKEIwbgoq68Y8oDj8apotI20BgmCAZ6rYRMdxkEtf2BDKl/1XTedGBxAaE
domlMb908V7k9acYn4p74DtECb//tu+Wda56gBS8Eu9FMmrHBC9dGd673sZbC/7roS2/P6aLJOXI
s5WgNPVUtfpX6kAt/kADv1yZ3wreKhGTodmsgITGOtxoY6Rn9k1A9Qu3PKCp/G8hUPeykIjeBnmg
PCCN/KKIqtkJo+zut57/hCBXaMcMPzyNI886xbK6ZWhra6kz3gA20qwv+R3qd20gIFQPzg+/euoL
WSFAhs8nI+BtdyYqT9T72tccw7dHB0CCpooPPp9yjMy4+KW/EI2r9vvelnJp7GGPc689EbF+fDAu
a2RSya7+81WT2E6W8XZaY9wHvT4unCWhR7GY1Stqca3JyfPdyejDdoXPjC6B5vCcsG7Eb4af7zGU
g7TEB6c70DhLUKtUQGXsPxtN5nLl6bYh3NRzwEXKBX86+XpA37+rCEuarmh8xtvfR6W04ssNCKio
GVcce+H/wjRsVENmCnLecUloAEkbcUZXXxCwpBdr7q+c2/xwtuI1HSA+H69ibFkdBX1dWbVMA/nn
jRnMNbUNbf66j329y6c0cCuB0ni3P4J2BnLLqrfymM7x7Fhus6m8/NedzIV96zXIXnQP6RpZEsTs
20jhGkJGh6IDtRMpY2riKH5PfMUFvI0doblOl/R8Kz4x0rH6QPxU8ef8NQIub+2YeQKHl70aPeia
MPYY2XUkuF+eum+OOXCM3jnabOzcGTYPbol5xJs4FpF5NQ0owJQT5GnFLSWygL9UdOyfJFZjY3k9
r6jhzmkknjmvXO5i9z3xIN9usx4Sgbw4bFRlv/Va8pUG532fvks97UpN6F1aa7Q5T9nFTdWPTyJj
+MTJ+Lj8/N3cw7g1xt0PSd/N9ufg76IM0xOkzgCR7jv40b66pVMjbbdUymojkqbaVkz5SIV+UhgA
UnruE7WSp7IARos/J002e1EB66Jwj/O2FPeiMsZceHHZBZ2jqdxBH8kuWx4P7UBopmJlnXD0WXuL
e07DVfQsThmpc3/OoYImZs1L06tiygEir+MnAn3QaCYD84YES3P4by9ChydOmMOgPLJyJNdkuv8Q
H+R+I+2KAsBmgg4RzHzSbOFldK96OYLURaDCjkNawxpGn/dx2aAP4grqhbQEr5R5N9xHNa0BTAhN
WYZ8RcyHOLa/HJlR+RQH6ZzOTW70n5Azi+KgVPOyY8qCqfI22DpjIkbPPxZhVQZg8NZNXQe/Hdtj
Ehlg2LZPWAU5gXpTttASluao1CLYIcxD9WpiUI2wSJKLFi3ZJnrs7lcia3VahN6eMk+jRNBNLcA0
DpVMAeCnCXDVn9/dXD41oQSrLi2oWigkGOhFvfjgtnPQLZlVE2d82DGtaI61VK2U+vYjzinJC74P
F7VBw9JkMxKGWuSIQpQp0bDtSzyi7pjzgvQPUIkZJY7EMNcKOpCk5SoHYO9pkjTtTNL/2FVgFocp
M5yUYwa3ML1/GjEt6mlwLI4tZVVxRZpfIk7SKVn+zt9nJ+hAvFajDGumLjZrI9JCve5apEi2w6QF
/eCmTZPpMfUjHNSQvPRJhRcykujfYJL7H0JIMfxBCr/Y0hK7NYXEq/6i6l+4IDFV+DhzELv9abkb
eqxiSVNSH+5dy5pkbgYcZLAYihq2qETlfHD+C1YRMnkt6wR+CQfV2t/aniAEJGyzzlj0H5l/iYg0
sSQdpbsKG0SH8S8E+ThbzmHh5CZjdOW70gusEd/RYQvYqI61DpW0aRG2FLSlL/DZTISzdbIl+xNb
T7PCLTP9FljUHeyRSsTJB7rsCk1GlMOQbUD/925elg6+NMgVJLwaa+COyd7RYjLKMJgtvv2aE6Pl
UKCEF+UmV9ztUrw/yUw7yZyOBqk5WRSsuhAArzGR2wV0//KBvShkPWDiEheeaMB/STnWKxPZFwgd
Nr8DbYS0UyWEKY9AcvIobWCIrMT5vy3UEGge8JcZZ9KveS2g4mBscVilLgOs63DC4r+ZClg6BF3i
K8ghEDKnLQ+O/qhEt1gfeLCwRk8XaT4lbvlxQ1EEOfjCzISfjFmVPSUwXHcWP2FNMuLaLn+io+yh
AmXmG10gOHoAE2uxTei3iO+SjbozPmvlaxAqgUKESfmhn5q/4pCG0/dzf3ezKvYVOiHoAQpGqWJi
qz/E2ZpzFdFJV0NRVqfBEuFskLKcUwdFSlZavb/D3c1QIvnt8ZuOAy/sEQGyf2wW6fEfosGNVCQu
CaE32VuwPHzuDUVqywsTxUaaPOXHUzFDLVZ5CHmllgxa+diwBOz/LrV5FKIhmXW4H7P9uTi6YTUq
8Cpc9RGZPFc20vLYFR7sOfh5iCf4vhbk5y08S4SDYwYhxUaQCCuEtRHqI5xOhx3hOSnM8m2OZMsY
pztjjoDYFfJTg0m6DgD4OwdveryMeM69fmDP1vq+iVd5LfpzNE6mfGvgki20OKRkT1hFREbUKrMz
C5c1voElgxKnD7HN9FE9HiA1KjX4IZ4TUqLxuyls8gAvWU+u7+m33VvnpZY06oJP7kVsjkkeTgR0
1yd+PVsSrx40pUyANRV1Wbr39hJduChy5DsMZLizBGuZBiqZaZi4almWZk5MXOiHP+G1orUw8eQ6
QGiP9PBijz7sIcOUa/J/GFo3VmURO07HJ27XJKi9unEC8BvSwkSID3BPGbKefq4EhK6jF0jZ0yZu
6wGh//snRXc7DqqTvjerXjyTaPDgxCNJSOMLhw/k00Yi0j4QokQmoVFerVkczGAVyLzPr0Rozaud
lN36CVrtUyByrzgV6GZ0p3CjvdmPCgFHVxv/YCNnGw+cNMAJ2DStgKaXVQiuARtSNQifwkBuWsRs
VyEyiDE15gQRAyKeKILj6kSQn301fPFuQvN2Zpgphfnq23CqdzRbigLqsg8lNSqkMVGIZsmX29u3
NVGTWKJ1cRi5WUi7qw6CS4Gy7XgBJZAlXHwq3YDsIblg/8/7s6lJFltcSxYFGx1OfmRnMbfbDx1J
uCkoK4xkXg45glIFA1pbpq2Ti7x5obh+2UBCGfR2fYasZVb+ZASAsp6h3CyoWY7r0d3bVPtaGFDV
x21t37r7zpB3tdIJjwsovBppsY2Dx2Mm/u7H3ZNlxcpaNZcSf1Lwnm9vygpPlrfLC5S41LZ5OJG/
YyjdgsnNGwRyUBPZ9mFmAeOQO82+vcgDTxlzNk5amhVgGVoj5S1jpVQbxWFWPXw7gTaFoeyS48cI
J7XrOgYcOrGbRzSg5zvXs0rlrQc53q51geZL41FW8O2jpybVNzUnvSml+Dvs4mawD/EmMaMRl6Hh
HT2+1gV+Vu53fAGUbMhg3/t6hqn5KXzboy7p0NzYjbGXh5+0wYpFOUzfTiq6lhGEL0X3BQ2trSUl
KI8eeQ9Aha8MEilR3wNHawRto5tbE593qsZ5X6MzjB5I5RDJcgqxeS8gJ8DjRw11QW0Exp//8oCi
HiENetZ6izLHABVD8EMXg/KQ6a+Nxh3RMxp8o8OKmG3aek9cGV6t38C2RNZHYLMRgDEpX0XMGV3O
XOfop3FLUraPxkOTNdh3HJpktccvsjpSJNDt48FQVq0rnzEhwSs6EvriY/NGioNe1XvDDWY/RuvQ
71Mae/FpJNBiHLtUzIpwPPxyMdl99ttOXVxMPxesSkw6AvGE6nnhYBR2FP0nm5wU6Ewl/9l4nU/B
TTWMPMH5SWE+oDTEEJBnBRPRE6aTm2FLZMe3nhOc+qNyCwMdS8fvmZGQSH3jFFh3vyef7akWUpUv
4jESkOFpA4B15yenRMjvvA4sRWjxeIbD8HDIsPhtOhzPPZ/EuBug7gou53xrA4DiwaWJ4DxHF8Vi
QeAoS/SiSz9iGcNdy83z7PbLzbfB+8mANt9NV21LctZghXV/4lgUThas6qCEgqiTZtY/Xo5NH2iz
DYNZhfwxrJFQ7I9OoTkOxW9np+s5TW95ZIj1ODoDX1bE1PCrX0BVZ+y1Qj+1I528yXUdbERfgA43
kC5Q6V28q9fi/gtB+di6AQDXq54cnz2JamLusye0O+0RmSgtYrmI/DpqX1uxVDMBYPpKnXA9RcZT
FKCnDRuH8r/0eTXPJR5uu/jEfm6xQsNj4A9PEAJStw+0r8CpZlmHYd+q+jt2C+6mxD1IAsXmAPcu
Q/gJKl3pCnTZn0p4kxBV/K/6XCIAbje219aYu4p76dAURQyD/IG3w+XTP+A+otFRl2Ze6T4WS6ei
TvTmr/6E8HNUrmyXeAEYe50LNX3BM3z9dFZ9kvx7SJvQPVkik4HqPBCQrTjPAvocgFBKDSM0SbjW
FliUT80fDEkTfzs9dtUl5Lmw9apsDlcRlNt/uMXhzxScWZfr8hOdU3GcwIR1DmC2x7duGlvEzKgO
Zk26CQ2FUOI8iaL0NMMgfdRw7Ync/sT+svZZGJONDwzo23O73GQ3BW6mGRM2jI1ZDlsbjPTrDIMy
aAu4YmVsoRTlJ8EaS/Sr611ZsY8sdvYWp6wuScsrGbnALe6cUDEqVNACFdenl6yEnj/umS/MgrgX
4nHwFtNNYiIa2dCSTe++tVkNZLEoM8yxhy2l8d+1xSNNh/ZQWMXGW95jZ2dZhkgXvVGQ0wWi8PIj
GbKfKFuKmVTvEoAnlwJ6mtoznDM+4l+bOypM1r10mlPFhIxO0SeaC0fiQOozhaI3YAf2JpCRzYTg
zevmNIaqcdrz1LBzOaoQJphlZvkmu45Q4QQ5DiIL0Q8VDhRA7Ms51GiJtjV+2fDbgbjtK2tnmuFX
Qgxz8I9sLiC/Xx+lH/ZSNC0JAzCZpxtq8wdm+j4oKM1scjBnepWAViNhouEuF4LsM4SSaAG9KMD4
NrNJyj08NQemvDB7YQVvRZFwLGiWaRwk5pcf+UcDq2wRmwShNTGl6AdHTvgtIuTxMUA/EFBL9bvq
QkKosxelH+t5tI5EtVwfl3FYaDQlkssYD+TOeZuidrdu9ExQWJSXuvF/XD7gZGzELhzxogq2U3pZ
L4t9sa82G4nlvSEeuDNsivHmvkX27DU0T8ZL88uN7KId6KJBEB/to+xb6M9u51Kes/glTfH/NNJf
8Mx69TQuSUYhLhaLV1XMXBuLWD74+3Gmt67U3nGNbS6kXXLM6tBtmVdTyKwCO6G5ODZF7A1Kei/b
WbahELhBqsUfwaY1RNk4xIeXEXTV44EPKLiz6m8SKhaEknEI56fENqn42Q+3Gfs0/XMUvAlkPask
D1kbMlObJTMfhAcuTBfXR5MbIe9MoojWzavk/RKdJzJZ+ARpOAMJcKXDJ2331BLuPhhFOiecsdyO
8td/64FS/H3zQxE6P9EwCXSRiLSZxOLdHdx9o/eT1IO3rFwBLjA5h+UW1suCe0DAgWVIK69j2/sS
XPosxTYQdFUFWZ/evuQzF5nTEo+DAj5AYnzwpzpTOWHpgjsAqg51vRHwOxHX27LszEdNBa+HJjgD
Fwqj+F8hRbLhDVkpnvgmjkft7s4ZBZIIQpHdD3RzjGbCJ+d07LqLcN5xMPSYiNWi40NIfHRVy/MY
K3u4Gih7UuEJ+KRq9VnduLUBZoTQltJRfg10dHo4URKQcjvtZFQKo+EdtgA8DXdNGiRP8pzh0Q5e
9x31Ceek/IVQaldE62LeObG0yJtmINAlQwWwE3T/dLcOE6Q+FbtTjdpX1QQp9LHoAGnr7S6HcY0d
wxBGGhB/QZO3/zTInU7Yf0wYX6kHx7sc49Hk+QcVE446slxt0A4DSdureFEcLpYgH1vigQuR1B58
nE0mqsktXyz8eesq8yfAWkTvQHO7daUc4CJrO4Y9V2Ip+GLBQc7lNzoi9LXP3sfHgSJ/2c3u1E29
p0sll16KfSJWkOMJ3rn1vn6yLyDP7lmnwXKkwLanleF7J9glzBVmoCPDJifwLrLvISwokKsi6KCQ
d6enPhph661MWYLZkZdKkeOm60Jsj9xy4dEctEoY6ltwwX6/Ej3see4ImPTXxAHLFrBpQ7ykxlgC
RK91wztDfQrUq05Jbn2g1Bz7PGsY56yEzdJwT6KFPK43HFl7pY0CVsD7o/weMNqPEwvEwPePMr7B
9eTUb6Pon2exxnFasch0IJatGjI3F2eg3VCEGp6+UD2ZK559Dz8GD6K16eT7RhVNftR+AUzfBQpj
nJAwXjE+Bw31c6pKaQThqWF4eenoiWeKShc2aELZhLIEeStWwSbGnpXo6FC2WlfAqudN4xGut7kB
oPfCmToTqbKbWfIj2sOw6LTw5v8UcXJ6kTJe+SNnQ3FI9/segxu9WiETJkHm20u7md2gGrL6ZyNO
vUfbtZmq/DJ07mulE6iJ3/145O/T3x+B2maobrwUUqYJuR2uIKiBPdCOBmmCLu9na5Q+u+FgLw1T
/C/yghK3dP3JQSrN67/SUsYi+akelaILHefk0oRpYeBemrNoXYTrkdwRhKc1aWSULX7ZgYnQpQ1r
xDvQ22Q+IMBWvQrr7fTmTaxamfR+d+FPxWzgfD/lRjEQa2mW6k4WhcvqFubKTpF+zcY+8V5nIXw8
YN+Gn5VrZhy6vY14X9bwX3r9fnyLsSjioclvp/mFpbw5i57GxhWO8PnYUarNvHNBuCEjbaDqfPsA
I+oSeXAhKJqJRZyJS+03uDBHt5+uxltJI/m+7kf1Fi/yT+/8aupq+M4AXmdnPFBTqHzn/cTp9tMk
a+1KnmAjb2PmGdDFI+ijKzjKp7dGxOOEfdvZqW0Ab/i3WRzgFl5kkO3NvD6UNRyqLQ8ooAz0l97S
OD4dZOVAhaTHD2++tUsSkZaL382EZIQBDpZFG6rtznJUsa4tH5grUPI4/NnUlm2qw66WebF006Am
ebyyoiYmtuBsyZ3l6wEW7hspCY2mwN10qS75sDhrn7U085FJeGVLCZiozwhYeOVdEJixYhCnXFh9
GE4e/huYJcOWl5MQF6bNtHi8WkgufMj2kr8yMwUyfkjjTrovFvTd909FCw7l/fauEhWyA/9EAs+1
D/BFKEWIh3TolSVUIiqyHes5EIFZcDY2R588TJl6OwMo5xPjWEM4wdCB7wmoSSgTHTUISPp/G0wA
wdUE2wmFXK37WPQfrt6Mnu9JL/Ddr2cOFy8FCFiAk+3zc+Zsv3b5HbwpHwVUuoV+A4D5Z1Q0SaT1
Sy86L7ATO1xUfyGQObkd4PZYRnCWgGiUZAtcCcsQKRkU8LWNK21ue7p8Q6Otd76WiylVrm6yL2EZ
ZPjJNd+RAfPbXY6MhqKaG04agpJ2R7zsls0BDDDH6aCt2w5mSfdwbvVeGX/2P1pxvX6laII1eDiV
izrnZvd+DdL5K11wogXgCZDCtKyHl7MIa0cMx3xk2fvDr9l4q74C76eP634+sLvTt5LSAnafr+jJ
/yegupeAH04CnCLFIZF2sU3GLd+TXEaVmZlV3Nn+zFvdeUsNwwmlXLDYta6H7N79CbZ24MBJ7iWu
jDSYwEHCLL03cDMQfdjhtvR1iZCThlKdU8lwx/G6kLspoWxzNRAbGbugPrHWxM8v1FWpG8u6S04T
zMcnLaesej8ukOz7Bpie8sxjrkwVBbwqclVvOnv9Tjl/iCb15V6R8O+S88wyJfCGz5gkBdXyWLNS
zEL6rShtxC8xLkUAEqh4EAP8aN7nz0RfWOpqXZvTWEwVjkRC4nBLHPyS5e53y5ER92oI9QqXLTd4
RR2xARLYCfuAXig37xQvLhY7c5+HFAg27pqC4pPwXrqxoxY8oFqe1pj5RhW0foretseiUICWrmSD
w+cZ+Mllq10pweTS9l6n2FtqZ3i7I29S8sLUt82sDoWLAjA8jo+bQ1JLf/u0ED0xGlecFzVqxU0M
oQP+5zUJd3B9nLT2mk7KrB2Gj7Ztfkouu8tFQuepCwf0DO00B+2xOtNrZ3DUazGcQ65KHI1Xarea
BGKscd1vbbD24QJRrcMRBYe/S2om/JQerEphCe9xZG72sTN/1+dw/u/Nqlsh6VntZYwOyWdwlf21
yZvaUfnsuXxcCtu4HCgGNksgd848hQ5/H73UTyrj48pBDs7oW+M2zCXdUtiVmw/NiORRVs/5baMx
lfYFdeLplV2PMscx0mGw2qv7L/AbaNY6dvl8VZrsPAHv+HEkpqsmUZesEzBwirXURgP1Z+d04Ow0
YzKxJp5RiOhPBo8Yv4dBaxDx8/oPHMVOR+8/pOAP3JD+foDuKLN7V7DGmhAOHbYnCb8x//+lqxr2
JhklPrROjIfwFNSzRP/+DcQSNMBCzCsNYqyPr4BT2gKrkxUz1nu8CtEiNuCuiA3JWXK40qHE1tD4
JaXPs7fRQtNRS5nYDKQrF38dVZB16QdIa1o7Jcqcdy6Sfu1GFX0Xym2T8c+9RGKmgKTgiEXV38Ds
J4xTCvvuqY6uXt3MQcr+J1zAVBMUkiOP3v1B/0QwgzQ7IL5uO619HkvowRWV6Y6mCCy0898OYKAJ
Oo4FWqzaAya3YFrLhkjLf6td03u/StRymrrdEgHQJauucF+X0Y5ZgnoGHOdjHEfGMU8lsL/x4oC2
GQPfEPifYJ+H5X+eEkszpIlYebcMQtm3GO9tkJ4SJM0EZRJJiDe/GY4pArdfVNhRvbe+b0N3+sst
WBWs18l2DOpWmDyEsc6XcOg0SkCSOgqkKzNvS7bezY0Yh63dfi9YGRANDA5l9RdwOcpLLerzaeLo
aFhIssZgMDdwX2QjB6yP27+59JAz5JJTfH0AUArnruvNPdk1a67/iH1c0meMACGmHjFtt94ilqU9
buzOb8p+Z0kLMLRy47oy5dLmxfnMepWCl7eWzGklWQ+ruarE516o+cpBYiL2Yme5KcHN7OAthggn
XA5vjof70sQkSFtVesj+NPizeE+hpPJ3s7QcfbFuRG4fIya81/vMdac0Yl9uNpffScu3kz+2xm4U
23yZux/kkZpHtUUCZLhmcG2jRLWnvafqvT8slxI68bWlC83jl8+ALLtrRqcsWXpsLP3BaTiB9+PT
cu/4zQ2qg1EQsuMlkkKk9FpqGBcjs6kSk46Gch6TyqCQGQHVdv4JzqpiS+w5CLrooGZS6nadfEPH
K/JQZPvD2NBwk40HPSTH08AL7Q6tMTTXj02tY8CEZPh1ZITa17GFIp6JXtfKCcaev7WyIMOkSNBR
ocoxm0le5UqnpfeSBS1jvaks1QZ0mYXY6fbwi2A1PvVZ4LyUUkzxxRf2vj15/+rd8WCCO9eDwOPT
32Zsu7Eb9jMDyaF6cfxEbCOk9i9kQK/d6gNC7E+JovXc4qsJhCn12Ln5ZnQSm5FLCd9iJosR5RZ5
WTJ3IUHR8Ft6F4BcrU8aIaQ7GRppUdZ6ozBaiNvpj9G3BlKGjlc9rf8Y2XhFDrAgDggSJeU9gCBA
CgdzDiL/7DrjH/XbLo1YnDAH+UhifoRext+laCfVOWWP3c9b+Qkx9lROyFrcm9KQLNGH7ODEGCRZ
Zh84SGhotT7zC2398FoyrDG7sP9vSrkgjE41Dmbq7k+3SsIcYt6vugGQFRFjVSoErMl71tPkttaS
ZVhl5ZA9E7C9Aae72L2WWYr5tQlRWZifNHpW4X+fH5CqkBWCYr4PyGO/MSeSJqjAvmTgIjrgAeD8
CkItgZ2Ymp/TN/oXgpbdXRDpRKDl5iT4hbHoiDDvFn2j5H/P6VPmYBghKUvp6xwTHaV4rtJRb+Zi
p4rnyVPzp0lsdg830LipUfiEkLaR+dB5IYo37oUluXHAXBy6mx1IO+JFwKd+D4+ZUS0m8jvGxsOJ
KyhIlX3KansXDvGUtTKIeEt3PrEyp3845B7A7WaXGJDXDgiXsBKdui2r/OZnivPI8rWigKV9tl91
Oco5k6ohPzM55dd1qh97S4TZaeJaLiVQ2NBEZM1dPWlaTdAFkRpGfvSVeBNIRQo8etZd48jZBSzo
T4bSAR9cFuhUeikS9Gg98pnK3zQBKi08JnIoOLuMBKWPyhTj8AhsxcXAdYSEft1OZs3Pn2aeUwha
BXD5Rov8PKKWGPbwHMVaFBkk1+w0uozp4v5jBO4WVRIsAhM9J/2U6ozdyhPiaQwPziC7BbcCBMqi
Nfph8QINrWM1MyYtwB2HqqpJ15GPVZGQ+G4n31NDv58gaCPxmJy2xLguXe/SWEmyTxriOdjSnHoC
e38SLOHwMWy516lzrnhdl+42yk3AaBrhjmKTFQemAGnsuPOlIg2lJ2VRdR/zOU5l0nKsSbNTIGLe
rx0ePeV2ORgKm9e7b7B6Jk6SPwiX3FQCPHBY6qN9Q2xWyXrZGCGWqWaACTprPCHPgd8JX3MCpGel
C/5UpuXrAmYnSKWHI3OC+GlWDCi01IkDFmPIpoYfsTy7/7N+nEZ4g+CkEMeIjG6QKBIdGnVs7jB4
LbtWWAcZ/iadG2dzZ8s4ONPMec9GN114+2fTSPQXT56GCF4xhBjxZE1XRZAlLwNRwNOI1YHwC0A5
bggCL7s9VycoMvDMZ+2NL/tV+gUyouS0rdBN+u3glhgcmfDaMD078CQayG9wOapB1jC0H9v+MmRj
bSMpdslsEuLg9zbhvt5VwRM5E8UnGMFUTIWYU6pyImqqsGeN16nuZVjMU+nW39qn0IQnbQbiR4lZ
G8NXaYKC1chBek/nnj/r4+Xk1AhTbTIDO4t7fCo/NGU/PP8eD4ktDwMCMHwY1xMWLVRVNyp8qNUY
aUMyDyWGI7VYQ+fddoF7JDOQBdNQ56cT468cUTm7onmFtCY0/+eS62JeuniwYzoa+Ycq3kT0KTcS
4bcRLAm390rJ4jLou3TDTiSr9wXZrDlnIcI2zGtCP/L0ITGQr0u56nFUmDIBQ466arOZi6Cmo11H
7odt9GYUNKJU2kVyDgzFnqmeYuqK1+1mPRZ10lTJ1KrGPBJuobQCt0HjFsnCpWJYs4JC8CliCMfR
s4xtmXKO99EpEkt/N1HijlWI5y1xxh4G1JnkigWT1Jv7CCZ77mabf40cYMnWL/b+AMz9P7cLNSs2
on0oPionTn7B4MzDUmitvE/8IahOgzVURc8QOAiUvGum1QymIiKW4AGsu7un41+UbGYSCyjJuvuJ
e2eSgViUq7PGVgBsmj4rreObX0iHuDfUMCZO5gkczRxY8JHavVHkImGNjO5Wvfx3zE0/Of4QhV07
VRC125DmypB6GDwAlNRKhAOewDD7N3pxO3sgbYQq1WOt+gghQg1gFM0U6wtPLPbPQFyLiUamPAn0
IVNxjFiuLOLnALnAn3cL7yVkEPckwQ2gCOSNyqjt//COU08VImrrSo2kmZtXlsbSr2/gROAV15tF
Lu/ZeAztIxLSHgEdrtKtS1GYUk0kr5Z0NTzlpu5LUtryRvLLsXiAMBlYD0b00cylAl6dC2IwjwcQ
abAieCP1pPS2VmH1b+u/Wa2LgE4TJc7S617wVfYVwUJtE2Uqm3AxLD1Rstn5s3EZVqOFomgTEgSr
b5yXjcVa0qMsYf7/u9aMyqDG1NomrkzJN32StZ1uFGJ+Wv6QJooyqEAF7dhiR2FVTXDZwyrzQQCg
iMnQkbysVZ4ZpxfuFs+ayKXD4gtS1nu1RjSztn3ttFoal9xzlZNsJAu8pWjh+pj4NWOLMo29d3X9
Hr8KIimG99cxp61jZimXD9NPXRVOK5l8yhX8zViEM76WybSoGYDQL7aLw8Hzg8K6hsgKYDbLEoer
aMe828c3MZZ4yfgZGT+kcIKy/WFtl7asws02PXp4Z9kjjAzP6W+JMCkgEBCa3JFg0bkje6LR3x7Q
t9HKg7unkunm2t6tUitD7SGes2zcjOCzYy6hz4YImzJpyCDXTQ87IdFpXxJYHrU8Og/OgIw23Npu
Il40MyDGUfpvjmDqSeR9OBtCwjYajO3idNCs/0NW9WappIoewQ6QoFtHLcBAPkR99qfFO2LRGbPw
sBj9VsldxuqgUcYDdmh95vy/VRliki24SlrkJxUrECZgPOu67MyejlBisfFEiMY9nTBaS67wh8M6
dIr4qdoMp/0IimCRp2vKV/wCyNXr/jUCePz7bJl7ZB4WANFVmjrMMarcaBgf/zesckTqpEnRlCy7
Tji7FOQ0akH5HKrp0JcTu+BP5PyLU+6pD7WgM6XFuhw9AlNqj0cWPIcaXhWRosx5NRfxSX+AaQUa
m8ffvblWOr0KKbBJ7RjdEbaMmWHvO7hrUwKo20NCdwKSTjHlrnBieM2jfr9A/pRIcQIXrKtKat0b
QH6vUJZF9p71mEPmrDGRouF3kkpmaKWI00aSwwagPZrhWajckN+5w+D+/zuxHVUqNV/eOqHY4edA
TxJuym0gNXnS4AEfTc+kiwV4GzVQxz09qtj+8dhd+Umv2Zp/RcmIfR3qZT/lMOpuatETCOpiHzlM
22HHgOj+rnKntiDe+GZ8jXHAziVmB+3dwETFZQ4ORIwJFrGhJS29yqkQst2Ok9UQOMXhQiEFXT4o
T4Gqx1Rk5ovbe7xsWp0/XJINp2AXY+AUPseYRuSRpTIZXSh72GumXv772nFTwxOg1ZqMyev6pT47
NMAvh+3VU/K1zcPJosN38YMO90jFWhbkM2P36ORozzDAyfGpuUCyIfDPFFDVnowuo401T3CtoDsh
tFkEePBzgbGZd+NDsp6shIoLg674NXazM/FgRh3JpbxM3NZAGu47sdbW8Wz2j0dQtb++mQ5NG+hW
L2B4h7IMk8/IlkgeabeE8P6/ep1T7HZlCGI1y76Kdi/IkDm7+JPa7EHG+1Vfh+EJEP2ZHdyqfXJU
gTkSAUzOv8y/MJhtD3V0k0XaFTy/wGxewM6k4wXmvc3Y4MARpvsu7/MQ5a0J0SUxdDsKcR/J56+I
tqzjQ5nll9l5eYyDVTzQO6UpvblOxtAw1PcVbcGpsqxpWGq7NvLF9062iBXMLL54kXjwJixEP+lp
gTKr5QDxMl+t+U49kctmAogeSSxOSNLic9OwTc1UceZUm+4ZkO4IUmKctCVM2nt0Sr8JsHwdZ5T6
GoQHiXXlmKb47DR9e2s+fu5Ofj5s8Gf7Zmawn1xJyp74bfseP7IprRANPmTKCYuIac89UE1alKpX
0/aAVDXQbP0R5c4+BHB9hgoVaQBEIu0R88Mfj7hKeT7PbqKFKedG1e3MmUtAu+tJtyZnp3JbtLP6
HGdKYo0kX8f1mzAPyMQ/8f7jbN/34OvxcmT7lc79DyXt4L41SLFxI/DP3jmZjMBL8DrTZfNB2+bk
ZX1wlX1/YtXGaMuv1M963qQksPZT41oi/Cb2tVm6NtLjaxToemSs9KWiotSszy5RE6rVXOFZXLYP
a2sQfF2KGBCPxetOYTpDZ9v/TLPlaBXtMXsS/+GlBPyHqnQkc52pC3OvFzgg2kZ3/l+VDca5VNmi
4sVNdJE9jtuBDAYy6zCrQJqAGtWjPLDi/mfOxoTw3a2EMUecPBhjVPGqdlApnAkEUJMRADXgVpwF
2YvWLjeO+E3w6YY1ZwLoipPe64We5BEsN1io8vsch6Sr7CMEqm7jxE/kBz/vEYw7Z55L2kNuim4Q
vZMaUIxQ6LcQUjyghV4y0X2hTCQZu0nguLMaRBLvBipG2PA/kuiHZlMo1qEzxHg69DzXVUIAR9gx
WT8HF2SGkCwjJiL3fQgUaE56wIYSL76y6FZhyP5XltNd2g/9Ln4zEjvFxXMOHA4vMFjm8W+CpYUm
cUArZ/xb2ovjx3uvt+E8qJr3XbsT4uuPgULfm7olz9BNastMU0EmMx1pjKFlgokQDiRDzYXtkOht
mXEHFXTiDoY1DAmX6xNDD5MusoxiqbaJD/CNeInSK0sodymkV7pUdai3nDajlTyvunY7RD5aACXV
N5TzeJAw+SnlKOm9887JBbV0k8SJNoxht0B6iZoe84w0UnbrAXb3KwoOsq+ozcoDjlNiQOMNecpD
0Fx5U6hTTMZaI+CMHaAdQY/OK0+imiMDGJn5d0bhGoCvtEgPI3R0eS8W2a9E0seJvzFyC+XvUK8o
4Wm7OjY6aQIlYT8oolso8p4VyOlSyYnHnHgvoSsCxT/UauSATCXJmum7qX/6keKmKv+PfA2I7nmT
BPnd5K/gciu/zmK8N1zkCbXsKsv7v/h3V4m1/4dG0b4ICb0yHfcIGArpM1KT/gzeIKWL574/PIZF
t4qkuzZ57b4iNrt3aYOom3nWjZxcoxKuPiOVAOgM3qkvVMxmdBdacZzfDyiZsz/F1e44+xs2awh3
auUVuB8YZK/V476BQ8xUcwEyfomr/p0nb4iiHmgnJoJ6LcCXrm5YWqkzurvhCQ5grP1Zft/5cjMS
CJICKzoXBmu39DU3wGF1pKLUc1iL0qxyKxOjpbdCW/kSHlcSqTbcEIxO6veRovnPyL+IOYxfeQL5
v6ZsPEM4gFxUGrbejiLBl2vc5YQVYJEoFZhqD96/PHo5WRasEd60mNlRuuRfFC4Fi9ZmQ95NjbZb
QVtDG9baBQi8MFqwFbIPP24wf/Y+sZAADs2prcdbFukBBhDPLKfDrQ50+jrY0l9F4lhStbPHEHkb
hIuFkippiavE0jc+ZXVjWiBaaBzVJwcJzBQEbAPi+cDt6BUrUrSQdSNzwIpxmGOnOjPFBy5PsSD4
Zd3EReOBd/QE7bHgElSRFB4azQFSWZ1kthDw1UK+ZxxmqZMLoTlLrkpVLq7BtVbr8Jl16/1vMtkz
eZF0wNc5ufWdXMma6pAg4KI4n0ZNPkYiR3bbGIYrSL0aZtCagSblodkyFiwFOkEKyYYkAGTBW/UX
IKVnT9fTN62TWayd0ENw/4PQqaSMAmd6uaVjAvPRaUX1Bqa8uoGWb1qwexAiyv+z+kz9TL1GPqVx
XLLiN2DqX2EW/grjhDoHjeQFE5XDXWYEh+E/COS7BrOWHhFSV1oP4n9gwJ2EM3k0lbT2BEB9I05i
jTAZHDpH8JJvzkG+4TP7LII6kIsUSI5fcdhtzQlnVJWCvS/C9yaKYVxNfsuXfez3XyyYA+l7bUZC
lPymj8UjdxXQvLJbu3SLRqKtMSdFzVFhKDek4PIuis3U8uRki31mKFxDg3TePtYEDVTtWIjomnxy
syBLphdCEfI/wieKMkst62EGch1K0g3MgLJ3j1ka33vMOIe+rKj4L5hSRgmPa67S+rkG8ClJpYDe
stXiEa6txoyfj9uilEjTIR6KDRD6hjrcZt+EqSvNFNqcFI11TobQfR3EbdaJZtTHVZCSw13Ytzjd
w+SByi9wKNIsOVsIDbOchGdOQuk9xrGK8WNuTspG1mj63dKgD3tIENvhIGj/ny1WTQjXYH1IETfr
+BBIiUyQyRre0lsOH/G8DSu/Fxt2qZOfrBzsf+mtZwM6GkW6xlkbHI8O/vKEgp6Ff4WdkThzQxKO
V6jUt2Bpm1cBPJsDwFqAfPLQFBctXCuy5knTvLoPUJOPh4IgEAJD+dmfIEu3td6FJF1UM4uGKXLG
atSPBd8kj8mawEnnkX/dbzNlobaUePi4C7UDhAitvdewhbfPvONSyKk6amZELJbp75iRIt40OGA6
CWCaRV7/3SFf6fTAeDjW7kFETSCWGnkZEuELTkqSwl2pVbqJr74ARd1b91bZejfuiyQsV/vP8fM7
g4sWKmVDti911Zm4Lu3vCl1YN2on+GwsmAtX/tZLWPMJBohyEbJEePxeHkJVEHsImmolbCrSFlAV
AM6U128BO97ZhtpgZQ8MzIytfZK/hzlR0fyF4JiULUeIjhaT+ey3+gsM0n3oYeJmuM3SCe6HRZBr
ElWXCfH7cwE3RMhpK/HEgUa7xLYnXsZaVfKoVxN4fEfs1K+68vrjqaoN/reKwu6TnZr+Bt6sdXf+
7T2QT2nhXZ9vWMjKioeklY9aLjZNXB71eSwh9K01P66UY+ri4Pas7OKN5jog6VQaZ7+I5z5IQEv1
R/zObmF3PWlerfBuS2thqPGSwfWJwluJF5yrVZBf4Hx80a2NRa4ER8htuCiFgCA4sPSOHifegnuo
iH3C4ZWxzyymu+OcjE0qlSK1db87NNKeETVLiSDy0ZjVdYxw6xJpEAzl7wVVzpN14rQFU8np/XUF
tXC5Bkcwb0H55JsRHzlT4xqL6mIOvr16yofamTuCUz32rYvNvrFMdpaDZSMLdtiz1ciHbLAK2hLB
KugfQb4EMjfNe4P4t9vYiVbvna1JhRCe8f6h8pIWw3d/Cw9Hes7XxmG9rJCxElWwvG0W3aMRhj7K
dL+CQJV9U54XQlJWmGqfLg0y5xNMrqn6mds1YhMH44WeiB9/Jh211hq4CU0PbiRZD+sXNuKtbABt
mUeRawlSw+iReDPKglx+QTvg20D5gNpK9iaNXBglCs146/OvV0syPx1XPyc2pTbmj/E910GnrusX
47ZxrS5EYj9UwdpSW1fHBwMoo/gcpNxPOEl9Hj9U7wXUFP7gxqNMdzMKtmpggr7TcFhQlHZieh42
X7U228LGHLYUrjCM+HHW7WqIcuP6bwgMDNiKZTD5y7XkJP2CP/qPj42cJZ+bRBda3LB6G0/rUB8g
FnwTqGcBkbNt/MGj1ePHneoDQYfryrJq4XQF4r0USdpi2O5Tdzo0WzYgoJ4fCnmT95rVogFS+NMZ
Mm6wBx9gIRPrL6QKJLjLyVLccc/akP3J+SIFjOgr/hM5US44YM65TGZ4fqLE168MFQ11q4l2eiIi
h7vkl2f7YAgWlEhH2aKlc1vYmJMu4zUwnyIKqqU9r6skVJKVZ3/Ozwn1vgNWU5z5LRBk/1YREfGw
o4pdqX0Nn9Yv7SHqWPQyPHSyQGi0dIKvpDHFTs00Gx0oPNQ6e6Zacm/pbIgbiQVASMt65L22dsrr
+Wins3kdNj43LBwuvwNEziltd2qn9uqhChxz1XaG60JldM6+LYbyRFQMgHuFbN1MbWlqr/YFXdhE
SC7XPcAVUZD5pCxFjIwCau8Z0NDeG8uEWHb+Xb4J6qnj7MHtKxkhqQA4Gqi9EBg0z/bQn4bmZZ3b
xLGjdtPUBV0WZd5FjDv/EyAVJWE8jQK17y0D2qJqWcjk5u3nmYqx55UNKdO3MMffCv/SCCAmV7lo
+KSmW6glObX8O8gLiIXHsq+TcwS8pAAawmcVlCRMybCPslz7IWntg14WaILjmov3w8kJUyX/4Ria
3H5UHLWiqpjcVGJ7cISuoJey1lKaZ/2BEhUcw6Aos/9cMbQAs2gxeId+t9RSqkU4W0zvVSzGVEn7
SsWKEL8CJbLLtWd7p5X3CJH/SwDIJWm8Pmr4vKqKd5x8lz31CKwPz1ejAVVH0sQFicJCJecoL20R
oBOdTiiRK+GKt+bAKQrsdfzX2EfEmtjX6OyRiF9Wd708+Eq2bEK+sk4aDNLGKHfAY9lXPsbLTWtS
x752j+0zpC/bTG9fnzbo1D8HeOMpj1WhQTVKYPwNHW3fAnqHbLEBxodcMWOlB3eiJXjrB/XWNuWP
XPVG9QVdk22p36gSBqoqlb4/sBrspVk2r6mU/O4CVGf0Mhl96S3szQdWaNdaqVqRkGvou5AAIdFL
r26oPJ0dkmbY7pJBfXGbiWJQPaqCj6eM0lhwgWXwmzw8NtPdW7mn3oycWoP5kwcIalgcR0BJRCCA
EANo91o7bU0RcyA9PFX8inC3IKYqmyO6RWM8Yz5qqquUisUVNXslBEM58pU7P6nAGDMosZwgFmZs
57lEUK7vJUWJj7Q2XiySgcPDhitOCdiJyfDWwn98MsKe++hqrMjWmTWsl9tbvcizZrKXbbIClfxD
0Nk2N8VjRXbeYi+FK1Bw/IdnD5ojCqi3ojCnNLUUR6HHWB6UMmsZtYsSqtlmfRAHB1V3nmbpJweU
9cvvsHvc5vmZHWSaZiLkRj0TnGs3BV+2WeWhCshmQd33dSJr+0ySIDNsDvJlpDxq6JJ6jijErAT8
B71gdj2ohX65Dcej98pJrfz7QegAEyi0fIxjqQWryJElOb2CxE/KlCxIQc3uukLTHDlXsga0i8m/
o2hsEvERaOruc9jBY4dRILvSANmX23SayXqMwIn4lXXdcZOTCNBpSN8G9nglRvYfDVRCGlOKReyh
F5VBHd8K0J3uoikx2KJNr2iLwJA0OLze4RdmTKe9Vb0qjJ4fLrvEdiuda39qW3dAkXmudUEqjmeH
dOfqCGYv33TXceGfk1UFQk92t9iMaCiTEnG27zze9VQtM+oVjhkaHhixhyeZB+TvRUFWlPegktve
Rz93ACNBH52rdPjyjjZXt3eJYIdU75G/vtm3MgM+ixGxJkmWCQIdnubUqzzE1v0uqeyIBO5HSjdH
YOJRV8XWcvmD6VOSGPmNiAlBUWMphlxT7WeJoHgp/QvQut9ZayESHnrQKcfyfktL0TQT68JhQ3NR
Hc9gGnrP9sZManLb/Hw0+CrjMFIoIeeyL55NQK7GNZrd3BWx9Q1gAd1AGVE/ahaIOmq1FTgBFyEr
QHHk9kv51BaHjMjHFEbThHtJEDCAk+OImMFJ83CiRcE3ZX78aqXI+Qv5mIvWHcuaapE+uYHnZRKy
r3wd6VsqlO13hhT7xJ9kO3xcbTCvy5h3OBYbiWnOVogGLMuNSuU2catcgMJRIkrvqghByiFurXsM
2Lz5gPFLeWhFR1CPUz9XmmAcRKCgAtYLHHYkdNJLWpAXfOXxTkya4WPnzgy4Vbnf22utXdsnRbbp
myX6BntlEOx+gpykz/gV0UfkDKLqt3Pt4GrKFUGu9GvE44gTcwNMXrqqE434JjK3+C2Lo4JzHcc+
UBVu5su3ialahV0gHCvJEgNEY2ZGwgmiV55+moS4nkcv+IA4v+ibi7V5out8pZW8cbMnD0TRmy6s
LHNqqaI/VhlnmwWeDiDagK6DAw1zO2RGsfEaR7b/QtPV2hVtekNNr827aWO2Q6Ukw0zeDE6v4EGH
liuuAdJSpd+rOtOoJaeHQwdP1ojJtk1x+xOYQte2ZwekTogLuVVUQdGc8PRo3IglAJfnWNQWPxAJ
npYyu6JHRY8B3gKDYDk33K7yHBjrOEZHpoWkvyLiA7ZRhx4XGK0erzl8BM/f9rK0/UJXklamvFjV
A5RM0SfwHVvmYE9VHQp5xX0VMaxwI01neHqLRBMC/sTotYd1GtDCKGpoA+/fZ9IJQ5nsJYi+2UBb
Mc3YbP2Aw9jYowsUSZx+djuIifQcmUIbL/CtvT2hX/FdTpZL9UNeIv3FcU+AeuZ3QyAEissS5oHD
FXyU2obad0WTV5lAymWtHQPYn6VCpLAYg+gXcQXomAyYmGEc4Cg+eckxrinbj4CMdwos280ncnXp
8bEh5aF+tJZTtpAjBYxd1SdMUdkI1fi5zddklUqVb363oZlyAwLpM7Jc9Zs+2jCk925PS/sDhwJU
Va2jJkshSTAih9wpLIh9VhHF0pq59ruuL6sl+OZWOFMXsYaMqQ696f3R4CIH3l9PxybCHHeoL3jb
Zb1LTEQWrbAvNHE904ogu4AANu5SGXSP6VUQURhzDoIH0DOP4HzUWuPXcnBJY8av0NPml0NrBsiJ
SCfUtti/irxp76NlMTbDK8TFHavtCAd4cjxcyG7glqesKZzdpHmnmsQVr1DuTUaGMv5h1atpmbDt
qODxUIqisInyc1yxq9U99D3PvgEIxcfpkCZJmCCnApw+vD4vsSMnErZZYRa+rTWW5zfELUVIPsmW
1SBrdfZjUN3ZXkqLfPZym0gGp5uDGofdiDWHoObqL+GEqpUUFXRqLKHFFg5TB3JH0LU440k2OKHW
SlUg2vituCyf2jsfWR4ACQC5isW1mSyv9erSOEEchZWbHFBS1154kWbyO9rwlKj7zoIU0fNqZs9n
/k3kgTtvk/MOSc6r1CYopqK7y84Xeyd85nnqCU3lMZrvijqukl6Cq7wo1B6RzbxWqCn8lMyngBvr
TNIH0WYJBnOUVY1HN83UWxD0VN/g0G7wk9e2povxPdF1a64gI7CMqw0bnlWczTY4qbWm2gARTbOm
t3W54YwKlVCnbVmK53YHIfklmFafRLJQ9B5b9khu8gqWV3unNhCjBxY8swMHV4zBq6fIJVNVOxoy
CRHW/siIJIwt2loMmtNIn4TNRZqGtroiPLHNL4KuNgOaFjzEJcpDANe14mTQgk4E9t8JY8XE7UzN
hfdwdNBhh0p0f348BIO4jCT4//7NdNhXosvv9nxKtKWbiqa7kwFc+u7oSiNY9OmxeQMbcoG0VwP6
DNIc/OjWQRh61eXeAvKLLtidzxD0V67KLXL8VfNc6IQMa8w9D9+yZBavZ/4UvNAL9k0HQJdJ+JVf
9btsuiUBzRSvoGoxjQtNVhc0JJ7xAVkv2jEQBN5y+ArGvaKx/yEHPTiRy8j5UczWfrskC9iufVTf
RM+Jk4GGIhAATvMyTiPzZ4Yf8n4Zp4cMJVxwIAnaAfmEk56vUk+Mw3BDtrSgfEVUmhrm1zCh2rqD
lR+YNK3cwd+zzbdLqR+Qe4PdI0QtpXyRlUYGWAjFnBDmDd8TUDooZfGT7/yL9EtU9JJjeecSd7Tz
oNsr82J4+jaNrWBZ2n8SCZsMTeHHCgFSEz1SdZYcWrDtck9GwFSeabrM909yT/z22U7gg9VclZIs
lPdYEAjhtMVNnJg3eisQH5fUqbcEPGAFUCDh76IMD3QB0LwFlHDguPm3Id/w10HMxALW3Dw+x5Rp
tRv9U8TRPhrjMBdQ+MreOwsnS3N5mH57UDFXps4r6RfgItZ28aiakO0euRgqdfxmGPPNICfyOJD9
XMfOeDB9CDRY0TAvJ7ZA+G0JpdxjmnNRc4hEtEhoDup8j3qGWjKBLbyEM8hPXgSVqNLRPpUr4aot
EL+17Ej2n3Ey10stDhKV7YjJnqjywjgaE7LPtqFdS7B9QeQCzKwrRma+k/fU4A6Sto5HrmeMKMPk
w2b+aIniBY1TZDHRQ1P+Bbav7takksCU1OrpaZuBeCWkFCUnHhdgPMTMz+0pne40Q61mU0sXEYYP
esRYsSMUgzgPoiZkYhGex7sYygjTXoEVOmhjKqTqT3PMJlQekhRQw91MFb6QeRPrJ1VUiS/D57/O
l3h48VyBFF/W7Pj75DdrEKmlPCQ6nMphbJLPoEdiCLjQ+jaY3+5qV6eotmgUeAN+Fe9P1TANrZAf
NgEABD+cr8b/cygGpHimqzsm0oRWTP0duqfORwTYoDHIp0AHGtDANkgUoTCp2I7yaVcHqRs20oeO
R4O1C9xF2b48tWXZ1clZRRyngHFq1ZVou6/jmcxO2mtTrwrWqpdt3IGE+NQHr3VdnC5j3zq+glrM
ckYVb+wGZRdtZFo3kfxV23iIKwCS0IO7R07EbHTP0j0Kk6n9/I46ryv7U8kteHHaKUV3lNyojexV
aeDgfYZR0HmIw4EGJ5vhBmEtoPk8JJ40631QvvEMLgx7i33DMQ1GIzq0sD6419arSHTg1mBPGn82
uAbWihkVZCueKty30tVhxPXlKcpc9D87q1e4iihmurY2u/ViZQcbHOmZP5vtG0hcna01rG+r769Y
/35GI84rCsvSoO2J0AOsrjwMTa07eqVXCAIVntg9kSYo/uKE+EYq+lqet68HvtYzyJjr8jpryVkS
fwscDNhUHxk8whAthhyn/m+qNfhs22ZDQYAECPPLmazin3QY7S91RJUSAalewsDrTFA02PxH4fv+
sOkpDbdoZL9vBI//DIu6NdILBmlhVIA35yNfbtyk4RV54MndKLl+g+NLglKVjPsZ36NmQV/llVr1
iW9VHRZqakh/Repq6Y/K8BduZcN1hf6HS8+9warUPMCaVLJkC7pxNQXgvRwoRuQkgE7bK82I6SZJ
/7UBXtziOEXXcXio2lCDuZAYyaDx1/mokPcQR2DxAyyh6w3v4LwGSnhRgraRn4DBEBooltQcT0Pn
c+C8mHAec8tF/+lJlKMx+0fZCPQs/BFNn+uDfX7xbdfhOgSjauCaG+aePsxA5Xoaf5Qyf+1tn4x9
yg8oNnaXqgW/do6QqP8h4IW/uqQX6CGkVM4pD1heH8oJgP58Ro3aXhu0o7Y/KsByJnz3Zyvly6R8
H9/SWv665bi5fknJGEt2frV3PwEmhVC8Pt5+bUI4td85ddN7shxb65Wie9g8/Hgpe9IXS/gTD8d0
OE1/yCfGlMrov+wIOZtm1Fk/u/+/ajr9GkgK8GQnh1hV4WTSPQRTviT74KUQ8Prpfxj49gb07tZv
dfd9T9i7qhf5TiRkqccfZ4pBdm7UQvU1KU+i+/q2LSMcccmBzwI7YerLY7wpLy7XIcQwAyjVVZOU
jv5E6Dg41r7ybuVrMqhlV8MaixSGJzbKnIsFvclT9j5fCN0lo2ilkJWMNWfF2p7UvC2tv4+/z0CE
PLHQ1gwvvezYyrC2JhtfZc0Tl8bKr1OLnJfKgyk2fpzfpUeVoEyVhysU5hkPakQNOp8jQN3/feLq
hegiMc76i2nAyHwJX8+EWf/JZWvFBOWixkRg7mvsfEfUzRMgUaXROGKg05PkfmIy9Hk9Za8O9qPp
UqHiqhiPgTuPnNaAbrwi0F+JxVP+YbdTRmHZMropzH32bmGCSt8G49ohh68XgJlqS6UzKxx1nH1N
DEAy66gj4/IQRBahn0QaQaFer7WURhOv/W347ngAw5NVatGjJO1GqbRAlfPcIpLqQ61eGRT6fPO8
/WfAM4+nhTH9WMfLFh1/5CYTOTNWx45AsOIbxDOiZ5eL3AGCSi5Wnctrx0+U5wwtiCU2SkaKu27f
dfWnoHeVnYdg9J9fFK7zEYOXE6jmHd08AwX6iU0afE/kQQSu8Yqn5yAJgXOufITWT68SjXE+I59p
IZZHn25iA8Qbl6PfxzvNAHX7IwibR7vbZzUSGTN+R/8c9EmJRHwGnC/cGcev23yTIT2f7sSQbnUZ
zmQhyt6F3AcHIMlT3JJa9SLqNRy6FVsKSQD/3dR3QjrgsHPdpoLDjhaDNLLzvovp+xlEWXchAn/r
aF+4KQQ1uYpC23iQgZRRVh5pkL8bvfAgrpU5Jl0BI69ebaQjKV6Uk6rJFtqYYQJFYMR4xmUCB83d
n2bGMGnzdGMNhatM/hy22BN2pLGEVrEkGWCJuzK+29ZvTm8YPhREyp02Wp/GxgzjbIlKW2k8J4uD
mW6l3smq6c2uCqkyoC4b5cjRLHNKAJfh7vvWDD4LZ2j13ty66wwGOzmdeGR4+J6N7FXJ3dOTDnHv
36b9Yqw8w4HbJPgxgmOr6pQAy5yZ+Q7+kDe66uyrbofCVNcjASVSdnEJXS+Kq9efzU6I4GaMNpn2
wP7cQuewYt1XMEBZ+uQgXSI1YaFaIAK8tQh9e3MOPN0Nh/Kjh3NqYPDKj19ucvGjs+yWlO6Fl5t9
XSv6KwkyLxoHCoWqdIxrZPDdckjsqIPV3wKMLbdN6f9vwd2qB4OrnwoZlEGfsmbOfP5EIzdEHcwH
hf3Np+RdgDNRQovj52l74+BrqiR4FEooAMaEHzTlMktPvr1fM0V6Gt7FHh5015xL/hwCpYYPWEHv
bBeeanaCU5CtvZxmXgZzx0rZvYU9AqT/Ew5fxraTCYYHgl6DLELaO3a0Vj7udgxygvQsa0baNEF9
y1ufOMlVQz6YOv4uoAOzL2sKhTza7pzVRN7nMTDTlgn+sJ37KVDvsLnd3aLROKmG3/8vlqzZt2Wh
r7W20VI/WhdAkpT9l1vQgo6Zi8R/jr0BWOTfnSGJ9gui6FaYJAORG+6cCDb/+0CZ2FHFSrXHgM+9
OQR9SSZ2Xeg0/zmkzBvyi07qvYYK3YQZebntwL31FIkkGVQzRHytMp1uBxFikbfX4j/zW3wDR8kH
Ys1a5CCPC/DAc36cXNYyj/KBjg/ryu/fbqChJayDt9w9vzIOIIrSs3pEQZACiCZRrzGRWbr+LPkH
nvalVJwOj29L6FMTllN9GOlIsT+PCbVZ/8h/hOkpz1T1DfYXXUGBKJ8X+yfq4HybuiwLHXbeCJTC
v3MZF+FWXfVk2B2lL0IfJ+1Dpm4UN/rdu/LiFiwJw/39Ze7MuCbHS525X86oY8HZkHKRuV/3M/lG
T6cKSrV0ad5LpiBfMcISkV+Ux4k1GoazbtTkBtNQBLhUfQV0y/k5eZ1RJ3QijH2W9K3YOyZgZv1v
44/lrUkDa9ihH8C6sKPsP5XEH0fp+NqdFZJI+sQ8OXqsi28hEDfMRE1IEbKHmUhvDdIrvYFvmd8J
FXRlp6SEn6mIAUmv3luyXOJATigBed4hrGhRY9Nuzw56MEMK32E6I8DdVqophiuBdYEuN/EEDiAG
pXf/nni3uR7z4a67Ymxa7uMepQ7EPoVa9n5hXDWKVmM5u+q7rqGg9gzv4ViTRnKQSstP5LbO6Rmv
Nb4OjW3dohG7wQ3Dq+Ovsng8vW6AEGRddrxuejiMClupoRV4bIOEv8aRtyI5b4manvOaotoCVuBe
F1kZppmL0j2Z3rt0YOJHBdZZhpWAOFAPZX2dtq+yr/FvgZELlEp06x5Psuw6Iov3w9Ke3TdxsPXo
pxu0AjK69If4tkSZrgi9OhN2QSiJ8oGf2Le8p+Rj4Jlg0WYiE9PhQvxBrMfDFSSO6ERNcAAl/lu3
4yiK59dn051bYj264wEL71BQepfsu2EaOBGxLjPWbBFCWXPUTjlcrANsddnzlsVe0g10LId2mGmZ
iO26+pX8HXf8g9KKqNaWn9DraHbljLYCc8tR53eUR4nqiAeuBCSfUhFwvbLK9lmGO6JWaz4XEF82
hRir2rM3JbC/7Ua/f8OBXqsIcOjQsgVaF6Yi/MNbJEvngdRymiY/BiLg67zmIE528mPQW/FmuGuO
kym5eoorBrAYiFsUiBOBL3LcXcYHtEeZhQO3+5prdU1T11hJq7PnJQ/6xb8HpOll6vMStH3eKvXt
oPWbx5K3/3UeBqlew2+lk7UGFbaP85f0MwOYR9p0hMtN1ZSMTGSMKBZFopdcNhSpcHDK2hmb2MMR
cHeuTyOaj93jytIwRb85Ysy790drjw0jcIxzLG+7DY9iVPjiAuv0qKdHivBOB4JNLJSTilStxJCZ
z+CxTHzXftiOnmrP2hNBuw7fuUM0WxcYvc94PiMeBh7sy5L0hyrvn9SMQn1f3nYskyDGJOgg4x6M
kaKl4+FhdXFnDkW4/z4/jk51AaUYZQRQqgMeM+jLVvytchMXrMq+CnOt3Aj3xTLvKs4Woq268h0c
Qi22u6SWtfIJhQw3qzge/iCrkHTezU7TYYxVIJq7A84SpnUG7Hg9Mbd8Acu71kVYtVLuxvrxHAc7
3twxuSx6cMx4vXWuRCc4vHnY4MfbuurWaG1WtIzLpDdmB7TekB1dRV0sGf7fVbOI5U2Rt+1tPaal
szNhs9DO83LbFI9lzNBNKHJdbDw6dXYT+0iIUp6zBbSJXgFUMQUwf2yUJIpMuXUVosyxQShtcEuV
MGyCV+QqEixu2D98F699tQpQKuvE0zYVToJ6i1U5VzMIyLpkDzFDdrjQjo2FrYpa930RTAbTlrNE
63KpFndkaTGM9bABKZs+k901An78KM6pFEtDUkzDDzRfycFOLUuzk0ubd/1Fod8J86u3BouxXlaA
l3B2n+u/jO5hezAAfyJ7uTYIvJjXSenMo0g5WvM4dnY0dkRTkBzaL6K1uOVrrSmXaboLQO6Ezt19
BBfyBz2hB2v0hGhVXbaTC+UJJN2HKpNjkJeNU+PykZobNOM+vxgMMl7vHcHr1uxYwGNrCjz1DS/b
rhA4+lQLk82cPQW2RoPOXIsllObljPBfHwMjTHrALxXOrIm7qhYialpEDs2befcq/0MIlfmTafrP
S8PgYZ39v0mxPSQg3Rs5tkjyVQeFegOVHENWCVolt46O8TDv5+NRL+l+0hwxOpVeXCusmOM+6ZAB
BXbxKCQIMIRxQMeCvQCpNiDq7fnv++RFOhdyg9AsXDjlQlEv+FDxexKcVaTWYuYIbDLpM3kFry5v
A2BjF5ufTb0XYvcv/janL/fuE/WlAaTFW0/CvGlHdMJlACcfYEWJq8/MK8mPJ/c2yPTsAdbKC/3B
hH7iPyJtMrSIGx/vBmh4FWhaQdeK4a0E3j4ZKH8Fg9PQR1SOS43N0h0DtzF60l2r2B5X/Ox+ANH/
dSYBAM7GgaB4AQ41FB8VjFGPcJAnjDQiYGvaaeNa8thAXyTHTxOUTA2o+pLwphG1kWx55J2WB+mp
CkqNaplNKIzHVoOIsQ2qPPhu7w5UfxYbpy4umRykF0BBpHebf6i5cq5rWIic7XS0WsU9nY2nPL0M
/hAdaBn3e6tS5dnNGO6lOUyePlNAiGF6mdtQwCloQo3mkpqaRfEhpPAU28p1vLcAW+1y1BX5k/MH
sPkPDFaV+HcbAI9Mlgqv4hFXZLPtDQQ9yqD7LAKLot57YlCm6OdbDIoBeNTOfNonDTi9Xj7AE9Wh
tmpfHOnYaHUR1cOWInCEXZKDahCqe622GK47gvMJKHQUTLAx879Lb+8fog+Hgjk9QFoa7lzAWRBR
Eir4eZjY9pXAgtGUEVS3sfagNg1CX+z7ku+wVf6R3FwRQX3edARFof7+0fszmJmZE9YntfT1AcS9
Q1XsmnzRARXCZ+q2QC5WUewMyCtvNMZ/kYupybxOy6mdjfkEIISkHnUyk7U+FUy4GydX6jr3KrKG
rELZorATDgPxY3rscxDsBYQk5HzUTeVkJahPcyaIMxqDSfs0GChjoOaDcCQytwt0blXKn7sg2nni
mn+0s64fTZ4I9t6aeAXcWt25nXGhHMVEgC6HQKDETCDoKobtdySGmUa5xDjRskC2kxaPGItjrFwA
AFDlUxTDtqECSI2te00iZsomS2/1Eb3RAQ+IWtchzlwFz1EGGolHV78fmwR0yT2eSnzdum5RoSST
nOC6r0RXia1c6qAneqjObusUk/cTlgysnfW2jhS+sK2bFnfSpeTZanw5AWY8brEtTXehVVUPrDsW
QBhGwqq4gzGCEXYuHXb157fqMnZUFVR/hDBWjwAf6hT+qhg/M2LlkmDZJul5cIwnsimdtKUQg7i+
gg0vSJdmrvkuhr0pF7CBGpNobnDs37dDpCG6F657+c03vnmIt7qE9LscrEOluf8d0d1rMbDZARZA
/py8hDHvchDLbs4OuipSTem5+QDKZOJqgTLrdPHQS5C9pZ0UEN3FCmeX6IwtZAekddAvzx8Z9k9U
M2QhES7KCEbkHwjLjpdmf2+0RLwTVzYDRhvHbBX1ATrjQASNwpLyHwlXlt4SBNytMXkmLd64EMBN
yq7+JqU7zVfoan1dq46f0RSwlAuVBW9n3AzkgjLdBrjORr7n36LA4rWPUl+VjSs3RVkJJFywaTvS
df8AjhoM94L1ikHNrk9831eYQCvOSEOlOvPNJtFMJRA1OmghypIwUA3ruTP0XtK/aMYu5Rt0EJpR
SMW33mgGB5SoysG27N6g/db/OEDDwc0AbCxcg6STXG+31PdfLsFHSii6X5jZTcu8vR08eectPYMN
1V0yqOcyOkMl+Tv1LzR4z2gQQtmGcrFpsB6cqo5w5kbo8WJ/wso5Opoqw/tLrVYC1XqsWFgPoC0K
RUQBy08vniMO8mJ0dZI8AoJEcjdpjuoRfkD7EE3kQLEz41XThxp/WvQ+D3o69teNqXoPbtUJ1WmN
zdQCt+0+R3pqOuJtDK8unJLTjw0SnWJkIvBH6vVBp8SKvA4oqEZHTm7RKGn0GDZAooDoRGgLUMRW
jndfakqnTPhvYuMUsw9kKojtJYFh0Hi1EUiOBoVaTnnxoI8njfucW6fQusFxs1UJ+dwTGG3h54ja
iHMHo0CCRa5Drr5AcfTmT97dpaE5EJT6+O74zQ667o8K5SuGCsexcFX0AwUy+hq0JLc4psmHm7ei
CcOlaMzPN/dQmNpybwlJx2YirtcxEwDlNQEcdQKJ4yTErWUbhC5xGbtQKlE8O4FAQOwYIG/TYF7j
TQJO5mnC3nTHlkLmPyEN36Bv2MtwD6LD9RGGzRnFBNW4sff/jt6fmwT6aDs9AXZAkVvftrATI7bs
7hHCZa3TqNUPpLi1QJX3sooJihQWdkDMvQ9ZyNrkclmYFgbl7MJ+JIXct8NktJRJL5Z5kl7JOP2t
ON0mAbKn3r6CFMSZ5tXZRc8xxRb6K6vrtxLG3YV/wgXmTjhWoEHtGwRaQJ2B+PNFcV639rr7yjmq
qa9Uun01cADzK6Y1bDVxogWu48wrStsb0eAWLCT3/0+VW3BRTjRvYHJ9fYNd+Q5c54IP1Ll545gZ
OUswA3uFLZZaNSsaGC5UVUVpaeWsCwPVqo5pDp2T5Y1Uu9l/CivDRygPvAsmtbvq7iONUYSbbn+o
/DjcFAuL8oZUKWvsO4R0fjtmfZicNlT/wHyVW0BhupxZGo1iR0yiFoudsQE0+QKZX9VbhR2e/Xl+
RzkF0Txa2jsAUD7bl+Jd7z6xs2LFJ3Kml+pNPlxNNfc0e1nRxDjusJW0EauvQUlRccKO2qY+WJ4H
+koxlz2QIYAIPaIeOXAdNJ9rHnadoRJmXmSJrc44JRjaAiXzFpppaQLPgpoBA6GCMNSZwPwmkoMB
xXWCpqXLYJ0oNdVJlbo7Jv3vnIcLSdRMRYRVfr86kx6IPn+TX7fQGkA8qhfv63iP1W9CeAZ6d0gx
QNWVbDps4SCC77CoVBUbMZn2ROc6bNnEETWolp5fMJx4qLWjVSlmSy9fvSSE4AeYhlvKADTrIFNm
MddTS0qgdwJhdL1AJQbMWjcrPcDq/GrKvub0ibylMnnpC3KEKb3sdyHCfncFCOBLw4wvahqhnjPl
fBxTHZZ3lNdcrEqa0L/pVYLiOnCEVEBKEVfL3KfD8chUx/gEjmL5CgazW/A1H4o6ljs1i4jkeKKn
97kwPOTxqgU1DNLAouhGIucUf5fb5j5OuZQ43FmEkhlCsggJ0xH0THGR7+z2CYVto/94cLMfgTMX
ZyVRS4HRViOjQWJ4mnP8I6xhYINdu0RzH1SDyppr3aSA4iuMhXodiYw2tl5LuIeW3Rv8FoRx572s
SD5OkjJ16C4+iQUgjcemGQNWMcBTcg51lnHHMRre32uUAQqjGniCQbclZnz7lOcDGLblpxSk2MdO
FqFInyX/eHzpY0rWUvb6pF1m89q4+bQRon1O7N3QAnUE3SZwhd+eNk3SEpbtlSWk70JdlphE4TPF
Ig+pwWuJfKeuCwJHzUf7Sxvq4M63vAJluLYuIpkVNMevtl11Po030S7z5EvhwaVpvsE9wkPhkJa9
Bdw8jmGm05b4sQD4+WEs4MoEKd0rnT1wsvo6ZvwHFK9FIJgovdwVoMi61d7r8MPLxdLWuymAZyjX
MOk2YDaSZma9cqhEtqIEb5UL4sDiIqifhsgu9KBf/zkPsdq82li2UiFG3FM7R8cIStlRa8Nh7l/U
hEmdkbMTcjVyftzRbA0uRvr8RuHiapksFgnei8PEEzmuMZNsXEhIJKYjcKVbKkHFzfRa8jpWZymh
4/BycmR8yqhhHrFaku/yAL/haJsqy7CWunN7NNWawnaV0LZ2BOXgKAVdPLN112hq5XlP8GrDHH+4
f1mqajrHpGVjwvZ+AhPVFRKCCBHuCVvn5cWRQCfX7n7B6r+EyRNvsktYG68LL7lG0LkxwHw7SqFZ
eCnkqgrf6SX04qeOyuf3EL8UbAzKZWODedbDz5WSun+tm3oFeTP3TeBzAKKM3DqQaJWVA9OKRy8/
gcJNTcfzJV4xCj8ieEnxvJCL3ATSZQl7BUNZuIjGkvu8RRqyC4Z2wtS42bI9oUDqiImKo4uwpsmV
lp32FLX2//3GTgNoW8c+CW7nqL2EvAIqZttXYzXFCoqpi7KGM2kLoOQwd6QEz1N8P0F8jAFhLA7O
5MzBbXzjAg9RV6yG6ICE8nsKgQBRaVgvO3Q5svKybteQeyP9p85TUdqJ48q5YL+L3aiGGkSk+ccy
HToHYL3Rpu/uUaTnSJOLRjFjvO53Md8YUekxwW1penkiIrK4zU5im9MW/l4rjqG7Vc+Ic89HjHkk
76er3Be+lS7sm/rOYBrLTjI9py61MFFi4EeRxrAJMPvY/zOe88bnyR0FQpUmfjTCme8dwgqmnFqu
RU9VEAjb7Nl5dR5F4QA5P732wxB1j6zvz4lhFB6Ob4t945Ooc0MXmRM9osp6Jn+tPqsZte9Gg5AC
K1wAfJ54zajvIwMjEcMxc6PPiJVndxY3psqrSIGgn/t2JD6XWYYcLBBfDVEww8kCe0Fd21aBNqG+
HMnu5DK5DORidnYwITYDrAaIkiyVnSDXRfVd+mosqIY9xZJLOisvXAiR6w+itLYGlJVsyXEZ15Y6
Ad7mfsr/qWOKIH2dHsA+s4PXkFoxONMAd67xbtR8fcn7VtYA0xCilh16pPqJNretEtxS8gDCBxMA
NTo2Ke7MVRIZpqWNgqWFtNQv7B2Rn3Np2Qzp2v+Ly7pacHsqcgw9L5VFhVWGMzIAyyDqlVBoV1yc
ZDjHTAP30I/2fHT4/DXceg5HVBmXuhZEJc6kAVggS8PsiZjbszd/CgIdIPCDTpzduEuPRVz8gWfD
Ow22SJ4YfsqorL9QfkL22hyjuBrnMpTkE10Y1wwjg34K17GCta0lyu/UxyxtAZChFOiM/owUp3FZ
w6oGou/jjz5U8Qr1sagveRcYjF3JIC/ktL+3A0HyDbxE3UdIzuZJd+lt54BpfKwcJZsQBCiC62q8
r4Qj35W65/mXx5hmScBR0WBweIu5vxBGHZ5nog4MmF+gvtpEnVwhUC4esbuVRz6mtxStW5UWwbOG
xXt8MXyhr38g15tS8OUQuLwdX+OoyCtYbkELAEfywqk0mdBWZ8/gXtoRhIbe0kT/aI/R/AbmhOKA
RN3DFmp8JKNL3YXiz0JCarhel9ChuArjUvgd9mtCxjfNC1Bqm1EyCdtNclly950TQ0ixaJ3Gz/Yf
8dCgUNphRLvWBELF1rX4AZSsWm1YvxGphO1mwbUKxW/SIztKorNx8f0BFAP6pqJf+lrI5BTEmFB8
pr5a5hDIHhmLkYcXBhD+kNNMAOOsZ7ganRlOLs5jG9VEPbgeALhxlILR+oFKhXijfjkqGnj3CkrO
rZfYwrXMiDbn2+hiBEN7HUl32skCUoWIWy+XYVgpL78WI57NW7ciQzkozVJxBoZ2/9TWLb9HykNq
4Yt1SjncSbrmwwbnVkcSW2Ao6vlLHr20xWEUBvKn47U/AnOJC6a/d19bzZgZJETZZnvVzS+dGl2Q
WeWYHE4H5WQry8i89OuOfr7UvxFVzwTYtYIcfp5hSPqzApA+XNbwgQ4A0FN92lOp+ipRSGQhjqhI
b0fKQz9HhKFtkiAgxWmGdbXB4Ra/n/x1VgBekq7NA4Hez/eeWN7pYj6gmixlm2CnzkMsXyNVe+VA
XBjImkaNzTjc9b1tDVxldw07VAAjr7RoE1lX6pgNHnRvI7NqebHEDDhs0FUUjrsvSWr0TudvkTom
b3pwBI/HrEsiLdz8fmvYwgXmDbhQwDZ8AIHpx840KnogKu37FqCbAKOTgWJ6ROk/V/UP9CHwDe6H
8bpmnKivL9Vpktd3JSjNMWJqkmOoX3w6LV4uosu94eH/XlHH0M5bnsC2iciG1RtjzgddpCptQ0je
yjGByyzEczvXKd3sxlb2lbedXne0sPFJySC06U+oBtbwSk/KPZRHW6TJF2/86l2x2W9twsxjR19D
E/4IjfBWMa/qSaKMm0rPMZ+CiMoj0uuL49mCZAg5ILxI/d57T73QA4dnWt5lN62mZIZS2iqj1n+w
T95MOJQtixMQIP0WKaho+pMLfhJQvL3tRubXtGsKIvMsOl8CxhMPZlkGTO+sF7W9DN5BLjiPSiGj
QEHxQUw9JmRd1GZ+voN6RGh6MpucIOTw91JtmwP/cQ+S37gSiH3XRcWFSq9eJvapA7ZxC0StnsD3
+ROZo6HKczbUKPGfbg6va9KjC06+ZtXeX5QEHdq2rf0Vl3X42cPk5LVxjDvEa8NbtUxJPdpPD/O0
ISgElC1/WQR0wuRLj824gW8h6NWtzFHlrlzjTOqE5tZXXI9tSicdFdcJqZJ7rIEjmB5HNH3uC1tL
/TkQJyLtBo7NKQR80xykQVro/bhTxaRu29GMwtRIf4zxwSEsXKo0d9rFHO6hNakg153GMPpzpT9Y
20Mfw3zXH9y2o4N/aduY71e5SDJC9bAaVOUicPf6OkcOxHbRWOkPl4Kg4TGgsPkQhOmapPGONmsQ
gq1N/46yXiwr006iGLT9mfautSCqJpANqhqyje0S0AzvUovtH4D8QUOgdj1AhvQDAACd86O2Fomy
sycgr5wq588FFWCnZAQ7L7qD/rddJO3cpTJB5FkWQf2xSpv1CDRQZtqw4qRHQXFK1mD/qFQCMpCd
EdHLf8fe84idBOyZ36MabqT1eNWoim8w50F4TMZ6he1UT4I4y0p7ajRPw5uzi3lXdBsnngqx7Zoa
lD5tLkIytsprZKVLkWZHSF9VuMufsfEVVq/AlWpwKJrp9lbx17vkKJo153izzblrc9xz0gQCy8PZ
nFLREHTRmpWqwu8KumjjQHcbV4QnDpwhFglzZ6710zwSw+Yu52bpNFd2ynYRKgzy1wNtZh0/an2W
H33NkKBsErIHYpyBs7qJMayi3ayj3ELxNRnZI+io5cl9zAc73Sw50vFarKNdIBKWGpaLTLvmFaOv
nAgTN9kjgasBggS6Ifk7IfNi2vWlyJ7twpFL/XE7vQBzGefyBE6QrCgVJxYbVl64K5jCth7OObjv
WEgW/Qyi0iCBvRuF8s1m74m/yMDo6EME8d/QLpPeu9pLAcVrF28obuxMyES1FyAf09J/3E60t16U
t7idHXgjKb7GG0sjFMpHjiaDzY8FRqpn+TATAuihuRaaoMsB1frt1K8Pc1oDLnKjHO3uvAiANQaB
E46NpGzLe/rkLWAKrLImBHf/GHpxb5Y3b7+eN8KXdUjF2RVpuZiw++AuHem+CmXWOkR6CLoAgFO8
6FcHl0R2OrrnZ6UeSawV9/FuId1RBFXKpFXaptBuJdGNQjDbItNIdHE+GqK/K+k+DqLYpGtQHVFN
FdWc543Rt1Ww4dRYKOk8JBccBphJ7WrRcPj3zkIQRpGg6OyTh7Gb2c6AiInDusC8xf6n/tqnNS15
3iTzrKLcnIf3FfKIC7F4kiOhzc/FUqfIpzpjms6Jf0GtEn3lVD9TnbW/dL9RD3EIvqO9OUbGaftH
JxfdnivKe8QQNXVmZPkM7AeCWxL/pPsm12DOzELeUqX1gy0cGHLlr2d/WSleSn3KcxCtfEbJc/Br
deo+Ee1K+kQ/D95J2fq0cKCQZVbg2goSg72QryeRc6G00H7QdoKahfSmZGyplj2wcNTzKY5W7ZRZ
k0gjM5Y5d4fw5Xm4MYVl6T/RXD8jlgrGJhrDTULcn4eOKf9W4MuF/EKuqGoMk3TVkTN9neQmhsJt
1szELEHOyetuum0ETlYx24R50LvLT2NtKdfOEE/ApHxRAi+ar9B/xCpUsH+SKJQ2iRPPCiAueLO9
wQbZ/lue1rgJLfi56FOV/kMpsmrLlgP+/HKOuqxrnJg6GIALr7E8BdUKcw1N1ZUsF8uPZcqpIq7v
RWUAIUBZHrEGYx+5dF8pSpTHkgZgGK/EgDv2+Ond1yAG4X//zVOKhkW4+DE+LR7Ge0xaOonAAGky
sWW/roPMfBgEToT6BMYWKwJNFrnAFcjifbRhzRzNhFbdL1gpstCDQOMUFBFbeWPz/SYBptkLsV+Z
77C22gjZRUHFBhs0pdjXK9a14SxlpH0kGoZpAk6WByyPJmzNJRoQwE96OcgeRfopGL7bRE/wr3CP
ku3eru7k1ToxRQSTwxGVc8sWBqAEKdjqRvhol/vco4jck6DLHWLaV4as+r9gzSNYYxa+38qwPbRN
j379PW3pXyWea6aAD36JF1r/iW+mdW0IS1OIBkMlaovWoYZuil+34diZMSEMf1aHwZfbYwpDV6IE
SMTqSduLYkKbQ7ny/DKvCzBc019uAJbCNNFNyAYwiC47Ze5S4TXePzELm8TOB0Bfa+887HlLGt8z
/77QGfL7YjH+3HsUGkG+20tdKoJjos2K/xe0ZByLZ9gR7D7I83+wiD72wfLLIyl9ODrshI5BC5YV
6Gfvafb6M5mVgoHzeqj/QYGW42vVYXvmMQGln9XPRWj+6Bi0XAojLb0QVYc+sG0O2YB1+pIyRtaK
PlY7Y8CPUGXcaLUOTHapaP69xI5JJgh3WSsx0rZQRLUBFd2uQhEPM6lPBjvVkQ/2PK3jfeO2Ad/R
O9h5M62pMy6dt+B6W/xMPldwNJAOOkGHV2BjQ7DlYkHXbn+t9jN/2yNkKlB11ceUszTgRLTGa+Nj
hhsc+HONeTYvAIAcIYIdpE/CH6cSZgvXBbipQPUVXkvwc8Ji5RiVmmEksgMmL7pNOOUjONiy552j
d4+Ez9HkpM4kpf+ruZqdJvfXxOEMX1MAq4j687c7cjKuJMOBjqKCrn1jGKE5agAMi6RY+o0Tpl2N
xCj7AU2A44eyAcd7l3OLSJBw/ES6+lxDB2s649O2XZ5eJq2m4wC6udTwSeqgDesw6JL8CyBK0CeS
6qTx1rCAChNFttl5uNp7L5Ra8UMOUEDMrplEDHvXBrzJ7vVXUqqhT4945yFEEqJF8ENnZJohlK8V
NtpEVuYzDZw+dBiySKG0+noGCuG98mK5irMS65RmejQRytiuoTpsR11ZiVVSC/Z/AEJvRVi8WDDe
06ZF/fdc6m0tyqYgkP7aHJhwk0r9HNiYKw70amf9NztU8W7ipCGHaaRpcPhLw7c1iN/TaB6SKATC
kJu9TicYtXPRHAVsiTHfVq8MhG3cl2MdZUIUhlmHNFwhnm2FNTOWF6s4vFPjf5Zvqrk3D4w4uQ2w
8CnJQwZY62eT2oSOtw4midkF2/FRgIX7QeLtl7jbattn+Hs94ykcN+wQ/hWIdYJi3FypIpaj/Kt7
faZN3yoOuYzHViGAeGYJ4f13LRPWYo6JYydf0lvxJVMyhExXtEQNy3hk8yXab6xGzNjzv/iDeTW9
gUznkHvcwsZlqDN8nzDbBUYM30tmyhaayefioI3Zd0JU+/uEdBReQSMNTyA2cAqPSyX1r6SArals
RnZLu6+Ta47rom2CNdvQMzbUVb2lQixEVQlVXJkukPWqfL52Dm4Q3Ni4wXQ3jGGS4FsW3zbQybz/
RMB6mpFFQInuqST1OK7d/KbPxz+0B8SnOnDjTfUPH+JrKkP6Ef78eqlyeA7meu5x+PspzGpcJuDg
xzJoOyxqoTQxLufn8rQKr7fB9dhhLCVgqKaaxQGnx4/eL9tgT3ZnN3bnke/U08nB2o2be89bppwl
xx6N87dURb8zs9ZfbmW6FlS779hRv/0y3taUrDFny18c99RCWCD5mN26Zs9f0ygELkoLFnZ9FC0B
Q3bDpCtQhUizL1Xs4BpoCMOMJiG7XBPqKcPJ2927Ujo8oirQSv8+YI80/Bl5//R8EnHDpnyJF7gQ
SYjt40Pbo82wm2UWYpU8BoMBhtftJDERW6WqQ/vJ2Fhp3yiqcIo4Xdj7h69PbIFoweiyS56/hbg9
DUGrdrTvvTPRZMpizPYnM6UHsckQdgzbaiv6BWazGIa0f32yly3tmW/dhoweS6V3V7Dp4k6OWyz2
75z4SeE8KSJBnzoAv/poYiQtezYdegntpN/dEwKhdJ2hj5wAsp2lVUz/gjM8xEVSLH1mxCXZvA0t
KxLERND2PHCRftwyhjtuHLJbtxz29NhWjEnrd0kh29lRR6RJYSDGKspmEcMAH6tfhGWksTtuNjDH
0Jgy9WsbsGSxizbaGlDE9b6cAJju0jIfBCExnu/WiT9hzqxw6aLCBtjmweuBs6WhNv2f0TqFijwi
wH+xbiIVPd/UT9xP+KHERBeBFowW22Nm3iGkTiUqX/6zvXdw/q5XGIjj3fvvg3qmPDH/yeEI3PTj
XsDS9pESjtrVXaqwNKF1QifuLf4J/Lw38tEOij0FDTSmiOxgJZufGozzejjE39gEvVMQX87SW8hk
qyCWuEWTKr2DygE/rEfetteYab28aP62pRElVwvtgljws023z8xcx/gwAPVttYnrVwm8+B21w0Tm
0J5bZwmJfVMMz0wPh32TP6xlnnfnVs16TsdEThvTf0hPnlUmq10wawTjlkzIGZL4WHMDWYHeObXU
BeKBaSBzaN3kAwhikADRLnE1VoPTfsatAEOzefJWdxDoKZ1Ds1zmUTzVxFFajqX/OGdbGbpKGbnD
QUT6mxS9STgiV/GZv/OmuNDjZ21DHkAFt2aIGpqLxeT8HUlEHA8vnrv6MQao/eZ8FN4+z+0WNv2p
aW6Hr9RuQW7dJUD5Zh/XodRx/K3IzaRgqUQsMLreKaE4eKhmKH+bxmtnmIMzLeLsz8JYIfT2Eeg6
elz9LVDP425kuRE9OsR521b1szY3HWKNLFSmmwB69sA8UWDjq7kJRJNzGFTSXJKhudN1+ZHBBq4F
XNytrPsugsoxoAAlYxFFMc7ZM6CWPGIvkccsVJUUVyK7qU0Hkg33FGQNNMOvIULtd244E0tkKwD+
wz+s0G2Ng/d10CD8JAQNXMLd0oKmrxkU2PaaArdIclYf9jQoD7OcHk+QpxB3Rv+OlSCxNrL/hCiz
eSz5HIqnWVeKOA+q2m2JYaHIfobXUHMaVTR3czMQqhx5Q4RVD2j/VnMkwdVihCfoewSDE3Zd9Mtv
Rw3VOyLF7vu0VBhG7PPrDzk/qqkPPKcH8MvEhSsbsWyztZZVPZ238tO6WbhcIIQGNWOIZ3/03CXS
RERQK54jPsa7ZydYEMyoR8b6Ol6opMNXtnwauAd6cocSr/VSlWfi2blZ+e58BBBR9aNiW11SSznb
8OD7zer4/t9q+GU3L0k1yKws2JBijBB/YGGwf7jqmtFd62mMtOfOyVB+RzSnvbfkhhNu/afZaRya
Cmc0VmpjWGIhTmieBaPU/Rqab3up9c0S15Ra/cqZwG/SGobfN/tqUY0uwsYBXZbE6+dntd/6kIDl
XpTEPBVHvLwsgLHwbp2FE28fR2027fdUO2Vk3lzlvR3DRYgKtBoGNnv29HRDhzLCRiXEpCrwV8q8
GVPzpaP7naYJAhk6BU1B4pEofv86v7OjGY0CZt3ih/D+g2nVCyg9oRhLM2FuuNSnM2Cbhk0SHPTw
H+nlBju0Y04/mZp6oN6Lpihx5r8u5SNj5YRxIhOn2km+pdWlvkZNDKfRCXXJww7QuGBkoZCnRGIL
PvWtfsGqhpmfO5B7IKYScowieAXky9KokhCT95fVa8kkHS/mRWqnJsRKRSmNMEd/ntTjJpubf6aP
ar57szVLVg0n/eEFc1H1gvICvb5nVwyEdWNgVwDzuOjtJAYyTjB0bux30R/jnCKrHQ+jx1iogp3M
PvPURr1iMDeznYB4NoIPwlemmvRPZH1ISLCyPLyYWbUerX8bTNGMHNKhY4qOnUe2c7wNrQG7qxA3
ZsKDClrb2JkR96EaPtJjPfjw0YJa3keQKQHY008H34n3Q/c+mXN7SxfdPwyXgw6F17rE043YdE6T
MJnAsIIkTUNHryOoy5+BWyqEZLd3v+cMJl7lW9/qxdULpQ7i4niJPS/M83sbiFxbQPmromd7fT+n
k9wyGKImAjT1sz/rjmX891fu53Qi+PId4ybyTU5Tof0/GLagUuIPxVXXP8Cg482XRx9Qul2NM0Xk
sXT7nDetHGHFUpM8t9BHDi0E9NS4JCZnIezsiw51lLjmwD84R64NTiQw+BQ6yQE+pk5wZc3tiM1m
MVLPwXmEKTDsblpA+w+zP9iYiMLF/mggyYK9mDv0xqShKvufedtpbyFg3+Uv4R1rpMFhfXGEFtaE
C5Pq3IYuEM4ILBL+6TRModnjxVv8JGhcC1aO262staIPAxOJhDmqYVRwMs7o+p7a+xVGWZVhGBTZ
wjkJ2u56NJRw3vK4SJzcZY6uiBolWRL5lSWJOyzxb6mypc/LqnnAXJh3nr8IcS8DGn9jSP+fb/yM
Vks9K4sqT14PbcWN2iKr4wimxPJZLphy54anPZ3Im12iPyvsx/xbr3LxzsvKBceM/LNUbXNC8caS
ouaHcp7sEk2TspLHWonou7S37/Bb7Zm39Y4F3ba3wbGYiBIipPOOTLVC9f+C063UzUkWxcHx/+my
sI7onfN+NsrP3cigXJNT5RjTWaSkozw4OY43iPmArlPlpMQGPPRWM+i9g7VN/Kldw2J2aSv7DxrI
3nebgxIKDth5p2yTtUyPNhuIal+jRc2w8FBvpcbINifTTLroMLRelzX9WhncO6JhlDOAGoYitp8O
Zs/xvF7MnTJhF6+xFXSZk2iPey3Zk6bWzYuyU2m6Q4LnIG/u3ovj9TgKPKJL6iNZkKac/aSv03Ws
U++UqDEfAikQ+Sm2hUNMMLYsVOqRdrq2esDKImbFlyk2TXhlKcSMxCGVZPiAk9l7VF6aRfpmCZfq
LeC9j2xfj1XwXdkKF5LLJKHFE5SORZDUTlBy5NuAJcL1FhDS3SiubLrkjVg3V3IWX1wZIKSXWxyX
aZw1Xc0msF4d8G0h5CgDd37aFWtiid1R1lLYnfWH7DHzapJVpHNT1b0C7p1IVRqH8nzOpNCwh45M
zsew9H5+JcBpgFKP6rMNKrcCn9V1DYq9spmfYIh6/9kiVxsJiv/3gWZZteQyEXEPHcEDvLYpDhJc
Fvf3pSq94VnwCpCJPTmRm9liHT9l++suY/zN7GXa/P2N1ICNIzPRV4eUeJvUiWYNIuod0XZpse8c
quPlPOmiEO7rMj5p3ZBAyH/23ueaAfp66XJwozAF4FV3MWJFa6KpZs/1zKy0LoUUl92san2+EnA1
Hx3azQGjinkjFjjQoteCtJFDeXuYpUJ9EZrBPIrMdguPCkOwlf9xxOQLO74TdQG6/cqsBJXXchQu
T10YHkEvMw3+TOGRjpMx4Tne/fxs4wvfyXxbogYZ5/BubaqRvYUtfbuZUPlIs+BwGCaRdwcUvdMD
55srXPqYBRNVKxORMLvb7dmCWbWMjmHgNhfvUQUxtTCkW7MhPViNoXruu7dXZXw7gim8m3slRW2X
mUM4Cs3torlgDoBzcTGW/0Zj7zKGCF51LAiJ0aS1tu6dCeNin2O7x613e9JlhE4Qky7IVIZUp/02
yHL2qHVBjQjWrG+2fHvSQasDswyLb5lYD/n1DEKEEoidJFvGguob4/8D9Q8l2ejDMLmPvFMcQp41
Bh5ia5VqlFBKbpNM49ZBdH/xmiZyBsTHDIHXqu+w7cKPmDVPZYcFdFSmUf+w3tcDCZtpdSBmUoPy
AigIv5OeJozhORZsIT7Wc60mQzJ0oSX99NBC9mogZHsipUcbU7t6D97lQ5DVTtBBVMGvqvXTdUgF
in+hqj5tXYcwCJAVeqSXWWkrVsYSGvpVJyk7ZskGQ5xp7E2PYvaVXGyUE6SIUw5n/O3y6Yxrog+e
nF3Jd4Xyjvy2+LT3ssbc+cU4Ju1uJ6dIjud3mk+NSk4Mik9UYK8YQ1tMpJC+TK/FZIsZVyyY6ZZQ
Z9fwb65jLKgGxmSro2gIH0x50NSFJ23o3EMWtI/+PEKLd2iLyCoe6hP9zYDGaVVprBlSt9EVD+Kp
z8PjKbEApBa1b7jC2ndZIXWEX+ML057h3d1m47yOjqkdBeSJAF2E+gO7xJ/jHRN9et7zM8O5MnIO
6oBEU0SFlApo/aAbJzMbR0W+CaT03gt+ZiV5lnZ1Ue0e4WbeCwN42p2N9F5EDVaIve58nj93ep+C
Y0WqVIAB0O3nKi1vElbG/BJsynZ3zN0LN7t2Kyx3Yv/ix58laAyuemUQwHpiaLE3Vmx4oy6KWevA
xgvu35wuDyB25AjYSgDMx7ZGSDQnf3Tah2g2ct0Hqh6VFGqYXKRLymR5QreiPiiosLA4l1/ZBpYG
9VlMqFSo/vhU3Uq1/hFBFyJYHxsfM4S8C4sZx+UIDSeKO39Qoh9OovhB+o6hVBUv5utTYpNeRAII
YVD8lS2XyAkp548++piVIDTCFyJrYvCw+OtSCA7nOk1UThm/FbAAb5rs2oWQe86f7QYOs9HUc4B1
iN+7Rgx97SBP+go5WOhotBF+uwJZ5qMfrXqkkmSEZJE5819rFoB1h7tXbvBfwO7GOQ+7mEurvh0z
/c6OI1kHCJ5NVCzHmv8D6tIhwc6G/v9ApEJIfN9Q047E1qhzRclKTVQFA0sq0u62LLNzGax2K5M0
+kjPAgi6yP9Yxla2byV+fbptt98lDmUTZzE6yvmZ3AnaPJYsd9jSqkN9G6H/SXLUi/XhKRcVHQlP
mYuznLwR75dqA5Y2NIUetbWoo+uL6Sg0ZMI2c4u32y1VJH+/ZwgbpHtG2mKCa7JrWQu4fpNpRf9p
ML5nlIsbE/0ub25Sp2R0xlESCUqKHuPqu8sByWC4mydIAc2OucUXhvYCs3MAqOibkTUwlBaFNc6r
07tX1yptGiL/Kw/iYOVcFNhko85RH5EZVl5k7XtpPRxrFGn/HEV8PpVBYhVHD8Ou4tB2g2M+p7T5
7IkDKs7DtAjEf24nl2rf3U8pg7ulsxIjy6S9BfxL1cJSUgoijfA81HNsyZF8H1T0faSagIv1UPSA
87gkvBOcj6rGvcA6GyLHA3aF1LT8tlNGD7C6PQgFLW56l1s+Cdl8bJ+JgMsEIEwcH8BiLhGMr38u
Q5jcEfBKDviqYVLjVCDuj2J0bzy3MR3iJgdTD4RK6wW49gz9lAnOMzcQ/v+sTjYhHxGYhTUmojbd
GPcN95z9wSo3YtM+ml5KWKykDFNnaAa3eAf6JovEKeG3jhWRYZPfMRHQodQ1uYJVdWznbr7xXRb0
jCQVSIgTQ2H72i3NM46y+1zo55yOmxfJmR6gL53qW6Dt//jE+wWlrX9JtJjILMM1+7WxSilBym8L
MHgadB3fDU3ZyH7RorVVHIcOTqop0oKVcAZ//tjxuQ17K+xf5T5zHYCBsVY9Rt6v2SEMvTLXvmRM
9kund6jwcJJHWptRc/sja4yDGnguuDy6V3iSh+vG+TwU3PWyC0xvtVJPmUUuhavEMZdldYghB0SM
H97rKvdolC5faszcND2Ly01/bpRdky2aWxL8F70x1iCr3UPZ07anIFM6dExibuoPzEVLumrGZ4aD
Uji2ju4CQBtOU0OiAx0vfbTQumCaNr8Z4dsrr1HPJOsps5sIKkiSt26HVIE76PWUTWP2LWwiThT2
RO5RBu6T1LhX8WpcI6eQbxFh7ZObfDF9hMvocxVhIXi5V3pMHb4dMnZbVoznEV5+frYFVJCWdqfU
wD5JSLuvhkIBCXJ4xGWH6Alm2JTy/TDywQrzWqmhlGMREtBkTM4dT0zRwR0T1aiqxfabxZPoRiaE
8atuq7ex7jMnWfyq14zz2KkI4hHJH0Uronax5tkSnsRVYMrYTmrt8uS1MpIldrPT7toJa8rxlu5t
snlyUT/GhBkOZ7FOTaC6kEzKVw/8N2NpN1qD5XGvdiG+/z7iG5P9zEA5mwMi7FnyEpmyxdG82bCE
vRb4i14zfWC1JJcXMSCyKYLwz5ElfwwWUSFT7XnSI3JM6juqRi4sAUI+dgDBYdE7PO3lOnQmkEzm
o8GJxXNLBcQ92LX0ApaxAk2g5Q+/L3fxeYof1zI/jSrwiKkchTiVHSTt+mkYW51BqPl8JwFcUup6
bF1ATEQ6uHI9p3+s1267ikCc6PkXgDuLt3Pwj9JvOOhW95Dzg/eG3KFiqKBo7mTlxorBHlSgyU5M
TQlq/BPVM/uebAhut+AJsLIOU/DoBnqXFdYdFoUanq0VClu6K1RQs7r0Set2q3AQMbPVUgc/q4Gl
+BdWeQ4aPf98M1/Sd8x8i4HFH0Dkad0kb6fLqVXe38sHdUI5Zg9N8DRcnNu1RYKcDmKu0r5TFX9N
UKTwzbWWNmRMyuAQ0u6dmTSAGHpVar7YR+EsJVLQ4lfdIFObo8Hyd8qAonF6CA6I+fYuiJ65Zxcm
JP41VN3C7rouJ4dRN2uDnNwy525BpfjdNzgAcSYM4fmhHlDph1H2L9V5EBbgMCtyPhrvjRRqe/H3
FwKN/sn/UYEAFmwJ+V0jGAj3mYAT57ErBzRD+sTt5WrSCoHwpbW3a0XO/LCv2QhHY66fc3lqfSHq
GTxys42Wrgsb1dZWrBIXjeIoGM+OkgAjlSqwJlRFf4mEPhpjbFjp5q7915kKiWoRMXfNrHCWoc6O
poDipd2fxopV0eupcPXCBi9X8MhyHd+jsOCHDUQ7Y36Bo6RrWsomUP1qdkeNk1cbV/XBAJjgnrQl
UnLnIOT2U9qlT50RgQcKOCC/6RWytgIdKVF6/EL0VxbDkt3eraQUFcvi1zWJ9RK8YoY2EnCulXno
0q81mJCIpwzCwA5nIp6x8sezxl+2X1bRLVG8AyoLHmaM6Vt4o9BvuPeudJTKOQ76cB35N3dL1FUm
u4ZTJMX+YIDlnUuN6ISqBVOJLIs1zGnbzreVhJx7x0q6sHMaxFor/+297aX6NqusfhbRGtau0nEy
dU99kXplAe2lhrJ+gR65VLtRe8fFm97rndCghcnXxUh73l7p+ktT+5qmglo+wKvUxIjH+7lgRdV2
vBp8BgwIhhzfnm8yTWemiPmw2KqUyoEb2uZFZDZpiTXs01RB+1bqnI23+AeJSfwqMeRahRF9TSoh
xmVXFFULCYdO/zUPWjpHHDfhCE/eZnINtwn9CDOER5+4ao57wAJ1gEvt3/VN2gjrXV/AuT8E9Auf
3n+BdLvO8sYSzYGPcU+C6q/RfJfl/xrTrlS+SnYFhmfUWx12MDcinruJkSCMFGZwWY7uyb3mNv58
c9T1m2B+hSRA7f3Ngk7yjPGC+G3FDSOaQuj8/Que4B7Ddg1sXQm/kH/RC+zgk3e9QPUJGN26ni0P
zzr0X1xEkZGUbswO4yRtNaxERCnAbssTmK9eMar+iS9NzLw9qk1fDOkoK+gJPz6anxmvrrAkma1W
iS8NZHqdcwV7C8KxnC4if037Oz9RtUvXzQmBrpzCu7VWRZSqD+mY4/uQFD4dqD8+PYEHTyzyu89p
Exl+ns40lPW/Wm9DelQm97x+yZrMkAHR3NuDNjtCk9UxgEKDnsLo1UIH/5AZJ0YuUds2C6KlcLWq
NIsaLMR2u6F3CDuTvRjKzASqdlUvj6bVlmtkX7B+j/HilfBHiQAcvrTd+16hmy4Pa+UUxZOeooTU
OhzqKGVX4kLuuxUci4UGMWQuPoZrLWLIvaAGq6xs8cLlk1VK9e4MyZ7RqLCpJlzE5kt4GAxdIHRa
vXAnIDP5I3Wnu+WEmXuKjI3w6qFp5YW/A8Y7me8KP9XDQPbC/NQz+gWR6EXY+B/qPKOLXCDV9Ol/
xzIYQ7yfFWlIc6ytI3pHxbz39Bxai1faIWyQzIqFAOwfBKoTFIsiQf4gjwtlt8AwRs+0w0xbsM7O
Sf/7XFPQAsNqyV16apIucLlsxYryF9v8A6tBLcqnCCEOBFsXLQE+NUX4TQYlC9+z6SHhpiNrrG+a
jQCLpsP7W2o1rkuEbyutExFA6A4IqxorXgzSZ9c0CTDhf1utDQcsxfPwj3ENFaBmIjJ4T7ECZuuR
d4TrjraizdKG86lfYCTKb99yNMUcuzoZiyXL0TgDpuAIcIulMI0Ajft/AqcpB5cGmI0Xis47EPgl
MpNg7dauHqrl0jE2kzYRkXSw39dMlF+JsqGidrgT3OeYBhcciixoQGcqPy/xJ3WEo9Q+4Y2Rs3ne
De0JE41muVuz06Qd/Zq4X58LFHwmPTZc0cGKQghbDFOdT1yiWNzAXYzlMWaoEHn5oyS/eDmcHpIJ
qElR/j5QeHaknmWTKnMrKJkmP6rvNQEaeAfCVXItDR9hjO3bbnMODd3yzIOabMHxfFcIg/PF7rKw
2tihtpJIZZlWJsKpw5pjQQn24GJx30o/W8zajw17cnPJOtShs18PKN2avvS4+m4J1uRjEs5SUwEX
NDoVBXh3mXKSRz0wVFxhCANG9lWps9BLtG6mXcqhycChw8YrORqbdouXYO7C+RW2E4OlatJBSoT6
ByndA/6A5BcNuE+kabQxuhNd/kD0jwUzL/NOxROnHD9opzYg9APWy/EjNlMP7DmCH6wFNPusDjdd
b0bXXPPeV5F7AJpVmW9slTmnDdfPH14h5wFRobSsBrCAkI5gK41QWSXoQ5g4/aWOVunxqiWgeEiw
snXwYjvThtPvlLBJspZJ/W/KWysVfEBoCy6/zA9BTdYggv+gwfHqdmPWO+9kHc6Tl1/WEdbHyWdq
wGPZZ1Xh0qPcp0ZyX5zArcSKeQAKyiW1wVE8ztez6+CHjoFpTk1GzPcHlb6O3l9CZpyVXWltEnoq
wpHGnrS2reIaK1fj5WbiPp6qFOMf43cNXiEVeLSJSeeMxylE7Go4ZmB/5EEzzYbblH75njPBBtvz
zi8+lubje692Rz9NronlHaiOry49jRBcuaE7csKnjkxY2HX4xFNlFcjfi/AkIPbtOQ69jaulwzbg
dmOjlYNXy2Nq7VNh1m9V8DNRntFmiPD0sZvJtrFJnCr8DDFWhP8Eo8JZjSX+sz++LOyWLOMrDq7B
S8defDoXXT5+JwTc1BWekUteV/KsDg3IkN56fz9sumVgecDdlCFOhLa/0elmN+wVASOX2LqO+dk5
ghQQ1iHzpfHe2Uc389Te3jxq41SmmOoWfM6n0hsGaiNs2wa8BTow1kRo6jhV4vyFIO3opwVJFXy6
5rhinxysH7p9prCERI46qWKhDtDX5VvLnJ3fZVCoexXr9yZKSMsPOqrOob7LU071FNg/JNCN7xnV
wZuxW3zienGQeLHqlt7LwS/XtsLkTNi01xh9ZK8+lvOaX5wXLExSCVlgyNEcmEF4RZVFo8JhDSZa
SM5LRhvJG4HtNY/ShMoYggEDygPwIEbD6sdtoUrBYkvNSaxNG1EW4H3ryXaoHw2j55Ks2SMhbMDU
jx1EOjnPK3Y4F4PNS8bm8aJteBUgrhG9bgEmqeigh49V8H+nmr7jmIGDLVdDFpFWXs3tJ9v1IULu
N46/xbrpxAZf6bPdgzK/x1GsQlw2SEOf7ksGOok57KxHWbYwfTHhzk94YyIFfNpio7OusiU1/Ui+
iSbGOjmo530btSgvkr5WaxUDLaJFrobjdIaKN0mZS8D/IT7puO29ctu6yEgNqfYJkwPoa5we0G/D
j/i9xarzyuonyZi6UEkcUH5NcZVWAbljLsGqv/Umankveklc7uh79hMvwyzvpZt4F17t1TZri4BL
uHq+nKOjGQULCPBRQAl8xcwMW6f1mNFjFL58yrlxfwyQU9Rsd1FA6wfUvxXhqc8fS7X7rfk/QmYV
M3yZQcj2E9A0Kx1OuJyWM9zil8QWT8FVRk/Lg8+i0GHAAAL5iAEzs2C9dkR1/4n2DgbBLFYckJgU
ZIT+TKMrfUI/2ntuqLynDHB79j/i1sMzucu1v4hKiqhhyngRT1Ih08flOxv49waU/JgbY1uE882z
sJDQCMRp84+KUmShweT61aIhakEHweuk+U+g7a8GQ9aWwx9I0vCBsqHfRFC9Rgp5EgUAdNc8snQn
q3fTW4MUvdjSVBObV681PAQB+poyxokfzeI4Zx2U5J9AkVeX5ZITGJmJrIJOC46ECGzkLH9Le5ke
JEfnEiyFIofoETapR2YG9N7c5ysO7cIze4Ugh/iy7yEzGyXLiZxX3a8yZaY+fKql6rkgysxr9jsv
ptGAl+UKOneXbDZX0MM7/NiaRBE1lTBqstL4M/MRvPsMq5LJnjutnPT0GawrXNifEjDTkWcsKZ5S
4Iwkwk7gXywkFnIhMN5MUJZ998VX41bRS/Vd7+KVTxEiUSDEBDkkE1Yuv7wYmRuLrtwubtGTz+6p
UzC/Msp9rGWusAisPjgUat/gFxAkIa9dtoEOysg4Un2unqCfRnVkzS3lewdYyuW3/P5d84OziGqk
AifaPNpGR/TSLeicKJ8s0EGjagduJdTHtJM75EvJxl7BI9Gs7Gd1MybjRyd3Opfu7v6L+ogEjd6x
U2mihJZ0Onfv+Mhxg3/2GxMRRmmeWn+d6sBVzH3JF13lymPUIsbuwC4pFTjvDWYJinUOhV3p5rZL
+MD4+kUsyq+V/Ws6/sO/1+pQej+yTxnxCIizn05lxEor31Vn8P3Qgg79DgUMj5eAgF6VHpQiHD8J
yyqHw0gFiJX2AzGnx6o4mMCBl5TH+C0pHZo5mI6nHbsffrl/gVFBA7WblGyiYijeGQn/XYkKzmfV
VIyP8a7F5m5fMNvDsSvK5tzjUbmb6rrVlBGj5uFUxh9XMHoqBgz2XUKjSnYSoX9K9S9zG/IbIHjd
s0qXOBXYjt21rM4WMlb+tNz+lQVFHZViQXhSgjkYBRi1f32GU9v5ZH78WCsBOEpTjnl9GJ62EKp6
M/kj6WeTKmqAwtgoLH1dmIm2qor3gzSsQ+ur5btXWQSXY0ObzxUuA8OS455UoKuBE4yG22t/C4P3
KbTN3l6pjKLYEAk1HtIt58LfgOWI3m+7QHzbMyQsjE0vKD8/9IC9yjyokHUH4ddiDEu56EzfjcE+
hsEzJ5+Ir6I/VOStBZB4K2Kb4NomVbxS7xbUFbR2ntn38zt7t3K7rQYh/MgLf9gFh/BooBwYIkkz
ZCDCtYX5Z+2ONoEMd4AQwCTRz3H4KaadMvbyKdVvMPzt3p0x34ZnD/34mjnzGhURTPHPhGquhLbi
z3Smbl+bDtauL2cmYx7ga9dWL0g+GmSWJ9FQmjWmnzHiRfJAQRGUQgfedl09Kj0jfXZF8tL0KoAS
noKMDlejXizQs1byGHbm79zSQ7BdqoX1z/syB7f6RUUthiyUZmIvdoCK8UW4wQf/lQK0bO6GRFnc
tWQFiaEfCM+mWWIW3y1LlhyRIJnt4PUAKcDhOBpNS1ohBwXmSzDroQEB7VPWXkmjHF5/WBoN6Qhk
kYug9UZM7sUxeYLAQHHg0tauV4o3JdvUrvrL3gM8zeXVHnklCea3IzuHlu/yQ5+Ux5fN5bLCh0kI
yaKrWxt+cektTaii8Vf6vLJFjtuNECCj6KlBMzriTB+AaBI62pzfU9dD9VoA/xIaCUBINqx/4fYX
CrD7stqrFJDbMdsR3LSF55EPWsEAnoZOPsnazUjf9mGZnIfIKoWecoQmSL9hRCj6NV5x3kSPsUbb
Fyp7+qZjzDQu8q1J5v4KAQRMuPSerkfb3FlHH4OtMfo5j0zp/F6RPV9GW1f8kyWM65kqCvkLrmCw
XqW+h65zOJ9KdrV56hjTq0kYs5LqnRFIr9IW0XNxcagxgB9btFjAPgiIU9lXxyuAE6FwW2ZuTmSb
6LakHa4Y0JtIIiwMmvOz5zgudmVBJRjoKFMptJDcjfDID33VZ6RKyZ+Su1L6vESHf4vwjQ/5AE1V
HvZYY53KUAUdpbPAUyjTArMTUASOKYB3jh+NCG2qagTEsv1LgS3iEzTCfPo/uanJ2FXaBcPyQFq2
LT0eXP3jCp2HT2jJK+JsG0qWNBKbOuQeOGlqHid6PveYD+GiH8ZE72KdDfppsoV3NRlBYYM8/5zj
tHuM8XglmAXy1C1Y9GhkFFZ7hcLlN6/BCtVPDoRqIw0cUqlwpVeHJGIrEvXbJwGExoocunJ0iiE0
X/jdm7P+O+Twu15hlMUY3rF2AWq7rTHTi++Lc6AtGtBeOacBVuOZK4HleYLjVyZD8zeKTalG+qFh
54jplTDwjXXKuluMJj+Sgi60hdFco7Pmysxaeb0xnJkxC+ySp19pSiUdWtOqcuhvJweIt+UKCrPg
EoT2+FtElFASnFD5TM5rePII5RXsKWwbjWoB1DwabIxBz59ShG8E+4iys5W51QSL2YsSK/LKFlSQ
7nlMSbwTOinM18KUP1SVGSYK8GWbfS8SeiEHDg/8+nZWoufJsNu/0RiYgCoIdQelcTDebpiFM6Yr
Pc7XRPZxpHhoB9eCtkaYliwHJRk7x78CJvVTL/3DiyZIrsqaZ8iaYjToLWPDGOKgI+U014Cq+mml
kFk+OMywvq4FRHVeIyYlZSdWP8nZ4IQgElKw3aFxJHIyCWW4Nvs45oQ8MgyptWC/Xb5twMKpQa+S
MqIN/OeMvfjnh9F7kp8JfkkAvmM1nm2gbxJYBwVijqOComjZb8dwSdt9J1ZDhJL57PYzzsiBtwm9
G0LoBYXv5Scj2k4IdRArbpTMgPuENBF/htdy82NxO1YIb/cjsdIrNBn/VF5EO4T9VSHqwB7Jnrzj
04xISkIGMIZTINdeLQYJHew9WINanAZ74+J0LaToqYuFCCREi5FTZNQDiOAnIvZ6WGBNes7sm0vQ
a8Jl+c07gKkCiz/y9GnGF2W4pZ9yxFm78QcKrgyfZ/Bl29Q/1TjFxKPOgE32c+Y8clxOSHSHCMOW
TV8RfIYduZjMydPJmZIXk+tLYh89re3zrySG3Ajg+YvjbkDzxDup4nLcoMSd6YJ/nqqXmxjydLqC
e52FAqjLKa1cUF/Tfj8ugXtfuoAf18652rnf5X1ieDyeYCDgb75+G6KU5Jp2gh6puczJYUgWafhL
7cJQes6aPockmhiLsp5NQZxQH9wTQlnUyrXKSZsTIY9wug7aHlFgGgLmqLcajL6Jzvu7HoCvpMB0
JPV61AMXdin/20X1fDNn8zIaJbJ56MSEupYwSbbM1KzPmTBx+QautqWObodT1VMP042X9HIGrM0U
ngZe4kKpYV1RJGrqJ60W4QZfE6OXY0bdvkZF5dTfM+Cqxtztos2APy/6+o6fNyWJeDFptPtJEmS9
0wm1t7uR5bi1fst6gHAYblBeAsQZZ6iY7dR6SCrRMZIMHsfw7Sftg748/5IxDdR0fB9EcOm1mvXt
8VMLerGfMmGT5sUptp4omCq44NspJxGA+lYE3JUqNDXAhTvJwUQQDModc2Fo/UvEf7g6fhoQjHfT
j/vQLr9NnJNJ91BZnGbqUcLuyVBt3RNvVekORONsGtbV/ZFzLXkbRbgczYWvaSTCCNMYWcLNClWm
/Z4a9Pv3Cl1C1jdTRLB745Un4t/uwNUzGvx+TjXMa/6tHNfmol7kJVVGasM9wFmvj7+O4/J3y8af
cQ/eJ3UH4iHOTpANxuZZ5jjmJh9gCu+kcWRZjzfaddAHgtC023AeqqtzFS1zhWprHW9D0wLAQaTo
4McbePxtGi+ujKg5cCCFzbrCcNrLQNYe3O5iFk36mhYtERje4U3YIJGoLWSfEx5VkZG6YVg9zP8I
sdhY/rbYh7W+VquxufroWgfsxofc6qsAYB47dyMZNqTihfT1NBMaj8oxTvewD5dLPJjcsUIqsSq2
nfe1agdHTsi+TF8c7HXTV15DTut/QVANXheatz+sW1ngOWXCHBett96AllPxLGvg3204trEV+dZm
BOFbPCvPm9ACCvBzdP6Ho9tLAr9eFrAKdhcnQfCJFotuCvk57FA4UzRhNofqH2OKTNB0irAR25fW
gKE3IVd6zg98FRKRLzFssMDDO8Sdmm2wr+7GgrSOvnghYxHvoFBmnbfmViMlyN9Crxm/UoSXeYfU
s4cAzef7f82iKsMOCTJqCSfeIhPR5xIO8i9RyfAmxGYRdbAeIuNFJo0tFAv8b1MaOo4J9GN5jq+n
gUnF2+muLw+gBapp6ykbneKqqMvkovtFiW8F6T8nv6wRYG7oRjkg+goPKD84WKRFqiCUjsB6N4IK
cWccpPXrYCh0oF6Z8wM0AdeEom0Eewq0h1md07vY2K0heSjJFyeFiO85jGh5P+z0XHjWTuGMXmsY
QQnR3RZ30j433iDj3to2LEkIoBTTeEDDL2WEaWgRsS8bt9feZtBnvRKv+0+ju1feM452l7YT+M/Q
rwgvzPziHHWWa8bA+/YQ/GDevjMlv5AQ2buUWYh7E4BEmAYDGYVllvKVhfT9H4aJaGj9AjCox22V
3GjjeXS4sgby8E4Dol2y/LVme4L/L4qNY8FzgkG0KIwJmib4xlJKA+OVnzrghLoC4AIsykeZg0sJ
wt54KdV4MH3ofSMQmYY/xtDXJJ9pZ3xlB7PGi0uTC2hK+KzCKYqPbEq3EZyyuPBMVYpphiOrLqbM
J1dY87vVBh/OVysKOGhUxLjhjViZU0fybEFAz88XQLdkJQS1ZFSs2pxZ94p2dxoQy7LTSahBDzuk
BZmP3Z+5LTqjC8l8aaHfXpqsfqM6SRqDjCMvbztDh93BzhHiJNscl0FgPTBeKtzdMSFIjE7KHXFT
tDuwOMtXiyyvKp+fpsJeKp/Jf4TitRnE9y3kj1wNXUT+0J2UCCi9fWsgwFmSsRBNvO3y/H8nX3Gd
iyt49lAtFnT9a/NIj/PGjElyTOh9dTEBArHlEwe3h5I+Hzx6myOrknr1jeGb2NlMa0lhpp2VynRW
WnAOpWEiLeseDTTaIFpwRjXuoQW4LL7EzRqKzx1bpEWf5XQrbS0xOdmId8B1HTMEEkXDuUMdD4eC
yvsDQpWIZ2Fprrt+7urAT81+ye7vPY9djMo45YDG2EdZKy12Xy9VxIeotMURgCnGanzs7zY5wQsq
LJFQ7sdnGzuleYUOLrCeYVCxWS46R8h9ffdNsWk6g2ra4IoHxx/KyXCZfURjaKSDeWrOLIila+ig
vkjUbCt4d9Gip+u4i2M5vBKBcjbvxCbQ67YzrCziVHtU2mSyLZODHlxKk4reGZGoC+LU8ZaWvF5f
UHXpKvRh/C1bA0ywU2B25YZU8Fy2uix0kCSv0SEi+hjamDR8tmEVdd6qshaT7kgyyYdokZjlqdfA
125Qme1pwl0DcvRprd9Jmm8QWuno3ggxdqimiy+TasqQA0BKfxRDLUEsxmjdZMnwGT8FE/VCylrK
Ruz0tGKFyrpbCrqZgllTlKxQFceTrZcMeZcXUJcU3mUs48b95CIZtivtUByl6NZdhS64ZSgp6YNA
TMxZzFwsyLaTNVNk+EW4R525twgy6oBrhhVCAGOCuzjEoxVWsHG3hhb6e1Uq1WEiD+Jt9njMF3aC
l97YZevzIR9cfO1demVoQDWx6g3WSIr09fkotHW2SrrxyAw4TgTK0pJkGciEgSQzQPvYCVcm5nNL
mHczwSkV9raTF/1RI5mSaM7/q1p6tZkOFMPAkb5gBg73I0Z5b0rksVrHT1rDjxgk0bUJrDTi4bxR
+RTra8BVBNhCwjCUUhkuJLC6b72Rll6CSGG+BPbtJv223puh+NxbSEgk/5q4GdqZYnL+CAUSHEnl
FGArQDc771JEWrniXIeuusJqWWpVzDENqW1nRkytZLVSbFwvZkLvmMG4zdWu3rOlZOZAvZx1VUI4
GCWD3RLxHg0jmz/41Bc1kh+UZ27w8NM+pbcCn2UGs007/Qf6Pvo1FiITwEeP0yuMughGKRxSTf64
IT6lXOUmWpkcLWrfS4PmZuEgJjbdP44RwXvCJB3ixgpkAnlHWIII5k/CACvVIW9WvpXaDEY8FOcs
68W4K9O2UlBO+HRilErBGl0GtOAYFJ6vVHzXltzf/dDel9meCdMg4SQD6hwcclqWC3sR9lZoz5H3
PZFqHPAOiSDKKtJdj0fW1hwfpaIfDKMFyXcqMTBvU0ZsK0O/sEZWcoKHTE3yOB4VH2jh5Mg6lvbi
lB9R4SqRQnu8nSQHZenElNUMRyK/bkcGONRGisYKBUdj3rBZpcwyf8lhqZL945ZaFHbVzIzLnyQ+
go4rrxuZBerkfPqPc9VxZ6TDXX05KKAKfsXo9gm+aK/Zvm/QbFteum6U/wp0LoTERp4QTMT2xY1b
LKh++E4/p8pHq1aj0yD6OHuJLQBbeslGt8ZVZKyify+vOrziqu9BGusgTsQKM7+YxErN7NDbqBqi
AZeLO7/eXWsnfEfpChapXwJqG3bWTD+Ik+FOzoMhg09qxuaSxQh4hAwOFbKDY+fIBATjPD6ErfVh
N/qO0NVZQF66K+GbHPJgKH6OFSEISYAUUy+MZLgpp+PsOAVY0UBWpltV8k0M833MbOGDlu1GVpqw
Gr/TCn1qP7Uf76ErnOHKBjhBhP+qYtQ/WquWQylKl66zFTLQ3P0VKu6ZC/aaFGSeVrPqMzaP82Ri
iLheeXdWWMAiVNS47TA9IFl3uV3Kse4T4G8Sok93DaplSMLtB4sDxJXjJnpBWl8TUNKXdPljJ1B/
Yfw1p8sbUAVvvrlrbmsuhiDYNTOVi3/6FTEOPvD9I4j4pef/8wPO8u4qUnj/LuJBZyKSJ+X4itAW
cP3cZf6Eyy84n1T0P+gtQ/nl/IcbZSgSBOtWvyRCXcRuXpL5MTyf4HWoQPmDKUyCx/EVE/93YWTZ
1zE4vnNs3/7xuQbDqmwM/SrgHtFP3zlbNO3+a43i8/vQ0UsDrECtvrhW0BmcsBTLfFP+xlYLHR/X
Fg1V4Qcj2wTktha92G2tdLv9Og6NoJb0PITCyyshT5i034eXb9W9zVNDThrcREE07YY+R7CkHTHO
44BBb2lBqjg9Th0A/Lgdoh/eCj7U3U9TO2cKYPqyTZPlq72z3s2zBNaRjqrEaXy+bpgSzggO/M1U
jbiS70Iiv5YAqSrbqkAA/hkNPV33s172hFNbv1skRcgPxWBwko8X83DDHfxrP3mmFSdoh4/dNQas
vj1PIwS3R7VPxPIT94VriQivmfO9LH22YLrKFgcZEUxNouRMl2GvpXiA7J2x1mRadNscD+oWUwRv
RkipLq4qLL1SfnlLWX2r2mKUq9gii5AFYk9CriZmo38acU/tf3LyF7VlctXlsL1R8tdLwvrnoz2V
WkKRqZd+tj1LbMx3AKNpLgeZ/5xpIhcJ8Q2fP+MYNzevaCFjhD+Twlu20x0Jom893z/l0vtIn5QX
whfPjNyeQiagUKK72b7tNXj22xNRuZa4JW2ukAVOfGypnLdRsT+17xSWDSOwPFL0qqC3L5swEVu/
f1glhh0Ch13bnRunmJJ0saLNFPfpMnWa1OI8Hy07JNsJnfGve+t6bwUJPKz8cQh8GurBMSCDek5D
3Et4Ny0kZF2FMjTAFbYQ2bLTuh4tAkpekklBqceH8RIbeh/gXDyRNkfDjZwENKVti1+woCMYN8Z1
bIXZVIBikopD0swDvsB/nU5G4tlTNGtpEf1dc6Hc54v2IkvhBw8QC8Qg4Q18RymJl4whhK3y1uDW
LAzoDkAy/ZBmNuHUPkNKNjRGLTfrIRNzDdc+NqRcE2Yq9wWZV5hfh2hO0kj1b44IxX55A/sqqikQ
RVqwMkFqzl/tONSM+yU2sxV7FdIPTdbXMycAQuWyP6FkJ7Iz8mungi0y+m3DWOfbrwMjqJYcOKgW
UKrTSOs1ulhBo0Xaa0qbMAp2omd1a+HBPv95OqC5RZjOdMQzX1pyKy29pHj+QsPWpmIHmIY/lURL
zfBhRaYJOUfeH5kto5UoX5U7c8UrVmtju/7G7LaG5siCi0Z0b4aKn9MTQ3u9I9m+WLW1+5Gfdojg
rMC5zlrwnPLN84z0Fel3nuuAI623U8DS1THcGiV4VJDEjSlNcBmRJ1nwRznf1nrIjh0R7Etv/LsC
13b87HZTQ1fX3pu1YwwikVp8jp7+KVAUCoZ8AhrCKEd3ot1nddwRIdCHmNeGOk+w/Hrgbr+BrpB0
Ra9BcZs1WkZCzjyZSA1eHnUoLNuVFR4RSP/+zFTNvu/yYP8n3OKFHNljcCM3c0cX2Tnft35y0W1L
kfP8i3z/CbP2lO/lvyBlnscKp2Nro1EINKo8WTSNupwLm0X+GX5SdxgZ7QmzYgbpWOOHUR8gqoj2
RxDrICeUSLYwj0gffMOvtGexG4IF/GvCfHLT57k3Udbf9D8hOWMg6SDQD46BlK72HMWsUGnssXey
/jYlEvrT29uo2YsP3h2v3spmsnDlN5g+w+33sl1YUCG2MONXqndyAeuJHJqMVPtc4KgAa8ABUF78
wEovLElqC35nnlRfVxrtI6jf5Dt6Crtr2n9qWavtU23iwedK9v/KTnIEuil0R4fsW/WHv59tIm7v
WEvpJB/cx5rxrCulB2b3DyKtE6KEE4pWJpyun/6SAtASLNew6BGFqnkBpPRacex0XHIXwncERWpl
Y2wzFi1oo+WX+haWV4NE7gUK96WvIMSxWl4GkrOWGul8Lr55S7glb9tEFKiWs8mNqhpFLH4QSxJ3
FFYhuNqUiaUSVYw3QWut7VD7D/PD1IWFquB0ngo40HYWjqzTJi/5DYoriL5fz/K8hnnEh+vMUkbU
zefgbLOAtlSxpLluKMAQiptKQMPXcO4+SHvprgP8zgaxYmrlceDYFdh3mbl19sLPKjQ3t/JNiJCw
iqe8/uiObvpoToIQ126umWnoZR75sUpokHb9qR9Bnd/Xk+Q3c5DNUtPE75R5YMd7B0kTeXHpbAL1
NWlws3kEg2r+46jnqAo1JvSlA98X94M1r9nzRPUJwPbDPI9kFrxLRV/pb2TnyGUQqbIsZz+RsFpG
XSXVh5nnJL4nokFegx+mrkQEG9BoA1WRMU+LaCU581TsUkr9x1Qd4VHDJsznvyIRvbWLSkIJpeuO
/D1b7AZCqh7JAq/OneSIQqGxQwnrvqXLqBn6hQj/BesdjCQPvozadV194W9p+ghCrOSyEVaZ4P6d
HaYpG2Yk2sqL0LrSFMBItnea8Ia6LQZAHs7OHSE0hTTfE6263ZibO+IguP+JUzPnpeEDfO0/2t3d
fb2dnYzf5TYnV4rfQPS4j9VrpkIakTQyvDuchgL4HjuuKAkhXGwNe6+4u9rZmtuMTysiztbETVVI
XI7ZG5iuiB3D8Uz+00NjxxEgf0IfoZX2GurNK1ex00Z/F3VR/myVeg355URXMrvNe+nIaU7PDob1
XaYhjN9sktAtkttYWOm7z14vJnxdnsgB274k5lkHR5eSnKrEz/TikgOMgVf/9TObohtZ0jPUmEXJ
bGKIrigkOMhzfTKaeLnjtblzSB2OnumI3+aamjoOmBzyoVqBSCEegRZ1evkczefJC12TTJRm+xI+
aN774LkrYWrfLBb4QuuVsVirRZ0A2wHCmLsok3VhptF8WJKbLd7EFX+YmTog0JK9Wecew/pUXpqy
70/FWNr8T9A7+R2u9DjDDm6SbSGvLyB8NKUbfZAYWuPNeXr7xp6T+lZiIFyZtudRjOToKkeSdg5T
ufS2FsbcaElcSNNhq6i+cnq+rqv98T1WlC5jEabE37Vtwz7odb6wakyJXuP3mZd+jbUdrZf9/m++
ZtEBZ2/eJbZaFvLKJEdfjJAqmAj1n45UMAcKyMUnQKr3D8PW8iODuH0CSKaXq48EbcQzop+/Q2G7
xvDTXmeUSXLACm6IuEHItveYPktbvlD6GRIdemE+doeUBo66kl79sJeyXRPeS3OrO+9F/dWMJm7o
V6qzasDcvkPFdF+/gnSUCG7FZWQ2ec9oWHR7lRC1haXPbYdPO/lUvPGL0BxqEi4XJk2YUoi3Yb4+
FwEiKhMcp+Qvt+FHCripWUpXjRZRH5+ukLjUwzU9mOQFJANzpx5ov2jECILPjViIin4GHu9C7al1
WF7YDQU5fzSolfps2ttdIbriG2GF2hhELY4haxZ1r/m+2mRyIO544pWdMNvqIVvTSSr9nSIjpg1o
lVqRYsXC/GukxKfPyeSa8cdlSbpLwkV4P+1zLOif3HASzxZOTSItUDon/5jNFlRyhOoqSMfih7XT
lXuGZl4OesCqgAmH8DbMXBiVLZIhkhdNbfDZB45Mo6Ab86w2MggpN1FOd2C4EojMGcKeyADW2FyC
rkD8mvzcMVOLWBTZfI9uJSv+t6JMNSwC4GLMTgSdIsSr63SdLxJDuhBcX4ud5n+MNlFKv3lMisfG
0UyWR0xz970+Ih0Xap+zLbvrBrVk3TI6Jyj2qZHdtdE4dHZmAwuFQjKK30J7/G5am+nllob4bJAD
HJirU/lABV5v8D0KIqI/+9/2PETCVG0X3Le93HhmE6HAMVjl/Ib6h0RLxxBYzJbirpVK2w08dFSv
nw5sjtfmUM+QmdHZyLTmAy4MKYGJ41elmSu2SE57SLWLdf2BSWHPknhQwxdMHaK3EBjqIQvyTgPh
YHt3oKvfpoyq90ZKJKXGhI5Zvb6nB4WwxFQypemyfQNtHTesFl9D1MXR312CvR2QU8dNY/cYIOjx
YGW7+OTuoylUy7JoKbl5OtZoLNU0Kq3YOeh8J+pLnF6ksEyU8uprwQaHVbLY1B7W9W6sDilgisXr
6Btw2JX6v65KZEmahHr+YPcsrbR6o20T+11D5fmLp09qJyXvsWMz8BoEtm/B2UVXdvDoHklQJ0Z7
Vs00cG+MQcXn9uZPJeTnG7v10Zr3lurDlpUTbmRrnzBsph1u4mymO3hwOgjDQDI9QpFfdz88Coif
KpEIJL6LP9FUF0o3p2/BWxlsZ7UWhBGtikorCXV3gBjr63+cWlFLPQa/V2AKtbhZPIkWaJ5eo3YT
PawYl08HXFY2O0bweR16PfnvRsiLE24kPDcle6CLPf2oEKPExxr6c0VZ2IMVQYKGIF856wl3Qi55
MDY8iCRvQUpWr8+sSEtmSXcuFFYvOswNY9IqsMUIdvGmZ2/G5WhUSy89qPWGMyFLnYzx1xnRGOuD
hSIwMIpLXHayxVPajHNM9OmKgXCJta07m60lVSdcdGshlMd7r57hYl4jh5sh7gowMjesrDemLSV9
mZkI1Gc5fumlRd3+oz7Ro31KwT3ZkvjQgb/MDjsYMmVelA5ZvHMr+CupuI5b1tdruu22AGGGcuKq
/TKtYcEX2vit2wwQ97hU5wOXw8uZCH4lHs3UVUPjbWXU1rqN7dfI575MAgk35K9A5TYgSy5ONr8Z
RCCKJXDWriAFI3G9HVz9S/y3vRjn7mQmTbhtGUID26OGeGLY4j0eolIG9Hv1Wv3eMiK0nB8B9oxw
kSJ3SPUxThhofSBiCEikNq/tBklSAHp2TD0k4norXWpiTWFIkaFMdtV3B3YuQMHInAWiXXkLQnjP
+bYyrRLjfasgrnaSx8bwM9v7HR29u4OA164cN3wIUQlnfU0Dz8porrwuidyaEp0ITGuQDY+ckMG5
3xv4lRwJ8syKi4ZizVE0j9/3nKHrzMFE29C7GOPvIWhAN0LeJPRrvgyswtVUR1M5P4Q4Kt26AG7V
degZxy3v/gbBAc4hCW1xiWf3huv9dDgBhUfAQeSw6/XZwVb8FTe2ugwpWjmzumvRIoTOJxcNTqZS
+lxCW25xEeY1WoEyyEn7+fbf1QHSt4VjJadJvt9IV+Ft4iEHUPG6WdqYAAIOIpZrVZW9RQJZDb6G
SSS8SOtTM23DvgWTIL8oqq7evVWeuIbw6rGG7YoSq6YEURTL0JYnmN9OGP5+oIiYyVLD8qiw+Vnc
rWcGoBNyMX5kdOsdtETwYj1yTrcjrLEomwK1fY49fup15xppjKlmC5qQhffBZ9q/ZSmo07EenI+/
7iyJoigTc5dbAR90VZG69KSShwDZ6ILuOTFCCaZFlb627vIKMvqf0lkxaQ6FctrevJW3RCvCFwtN
l8nBRRDWkQp2RfQidiOvus/h7amTo9Qi+Iq/I3YuRUC9WJPNKq0esOkoCiCMWcVfrF2HkCzlFG/T
M155aMSv90cXaxPeavb6RDWqZCvj/WqDIOaNP+9UDM9HW7QUeWfklUHXdV1Rx2X7k8Vkoxn44zGO
54qreTReKxoOuZUPy02PeX/Qgz4VtBr3GQHFIad+ZsLuYJpTOa+oaULFjc4vrEwKFz/rO2lz1meD
6TDScNULmv+Yw3egXMCovOoAYaA0jx6pb+6bkF9fxmVprwX5rDFVslaa1gJyP9SSsdevEXb1eef6
rskjXzvk197CqeUzimDXGZtFUlRxYbKZGWIcuTRIYG/LW4EQTbFsRhxGdunCuefjGYihLenvs6o3
wUU/zxSDOZ6qTasLxUHzHlX45CI8eGWP/8XH5ZTpYe52RHcuRIrkJt/rSEwWMsdgYsCSnetiFSaT
gs6sZqUcYOnlXaygoCWwSNk/BdJ9i8zMmiap0ngKu1lSFfmGU99Lz3e9jdNZ8LxqyOm7tJoQfr+C
BsTDs3ROWmIXiWE/ZODDMJwBYO1jIiSOT5U4TJszo8ROnFZi5NbPAYhFnxR9ubyNo6Tu5W7ePpiy
zOEEHiNXd2Q5+GtwYeB15iLf/caTvbiA1Jot58VHNMdo+4K7FtzOP+qZJ3fZTdaqr3oW9PGTq8Dd
6FfL/5olMR31bmEazabRsv3jZmFhq5U1Dx4nFhHgeqCGhDcnenMfLfuy51ct4yicMQDSvzj5AWeF
7DtZjJErDPnQ/+Gh6P00SweRP61DDcLwlV3EHLCqmNcFEx+iJRrJbwsYqZCdfVjDQ+1GneLDPtG1
O79woNavdb04pVtK7TOEA1ddEMj20vo5w/taQP3PHVwI0G0ABmJCwK07Qprg0UJPr5SbTx3pvYQv
v7Nl/o3r5CxtsLeDG54tpjo7Hk7HSm8ay0lMZmMYegpXGWjf3VsLF58F7TQsyDrNkyBEm4lLODyE
REUrI413NPGtTKNbZ67AFF2QjXKcKiOz4B0Wb0upLYjw2Gjdv5wxtELOx+T2EfEFx+dD6DVgJU1w
zQ5Qh7MH6nPPVmm1fEv1lgbbJxsxJPCzkL6Ja0OLUM7fU34G+eK4ZdBHB7+QN7fTkxo7MvhsZwzK
zaIlkhtSO70M+MJJOi1R6gT5Xk0iBS9ONzJNBiKP4YURg7gpuoLSVXesRcaR934JALQRBpOW+QGL
YNzO/lRcDYIcGAeN4APBNQYbkyGtgNb3BS344cVba481xi3hC9OjCKUsuXtU8sW17ynHLYPpDGAD
eyP3rYNNqKErlcTHS0MROiMVTf5vYdzPwklDPz8GXA1bly7Wn8MkxBbO38ZXrhG22tyAqXDi+Uao
Q++hwDMDcvBOAfwoDiPv701gWpq21EcmvKxUs2JLUj39tDrKRQL4Ce9NBWKeCzCxhYPrkr5F/JM2
FBiXQfHFoznSOT2JfJzaVm0o3hwUohj8UL4d31uAFxfYB3XQ2/50QdSZzq1PblTJPvJI+pzRhuo6
tFBsja8kRSLKkoi1SG4RZSSLp83Tck9hzMaSSg2YsBUxOvkS3Y+47Gx1wzjzSG6uJrWdXxkuHnoc
L9qKyk2OD7eEs3YL7M+cfwxINaXtStHBP25F0HU5eoAa64iGQcR/X27NC5EONt/6D5c1T+t1VX3i
canFi538x5ssWRJXbQEmbs9RnipKknjBIA2lZa0Rx2Nt8/4DNfdi+t+tvr88gqs6YWYrh2AjJXjT
Pb65Pc/4hWDhZ6dK1NHvBGBoxF/xVXMJ7QyDJo45+txq5edCH2UNCqlvBTq7QVrQk1/b4e5LDiMy
Szd5c7o83viIhbQnfdKZUsO7yuaEkj2mcRikYA+CeB/dX2WkBSWYaiW/+tiAwtCNf0QRP3k0ngNe
fZ+AqfkedXHIwhVwGinci3YPqiWz4SyFoaNKoAlrV5utp0Uo2NO3rJ7zStz7XL2gWhN6vrxEV3n+
lQh3w0o74DXrfkDfp7sYLqGXlvR6y2LTHXYaHT8clMrrCAluIKNJh9UP+67oGbEEq9s3bXqeVh7y
9vhYQ6V48zMItDsNUYesKOGS+ToCjaARqBXfzi28ZbwKAzhGBm1l9F8z1VM1KPuD9rBt12lELnNe
LV80hI7fe6itdRKXQGvgkX5ah3knCSetC4PDcOqzWJvsmS30Rc1/OXrwkixaCxTiqr+Pk0cvAJ86
TTSIjc061GLFrE2sj1om80EeB2G+mKEn019gib5TcEYlwGveUYGVnMHRzZRttjK7aD/OVgrXLu9I
kdRDxaPg4LMPQmvGCK2O+kcItGl6r7eumcWs8+0Ys57Y3sVLaA6UHnjwncbfOUWvHmvnndZRA84X
eQSD11daMu8noXcV4Eh619eY7jfsQl6wQla4bY6majSNwRYbQOXzvIGtgugRtfbETRmYFWvtfBs4
1oYMvxScH6wLYCtlM17DO1C7GJDVF63TfvJjREZKSN2v+JSCwA8/Ap7L7f6nyUxC6sS5k4OJ8EFE
cVsSusTkR39iUj2gjAmnmOgBmtPvpKCkHb0Oaw+fbHUUvmM1r5HX52VxHpi87oQo7ccWiuRNkKkW
UbVwvK0MYxG2fcjb0RuQCV+IMfAcAwHErSm0tQzsd/4mNn++3TXWp7DsFbKS/KgHSwcnfNNYyHHs
GdXe0UaiTA1ij5/cLKI18BjIfwV3JET7M9PpkI8HA+f5pTmfwT2iJ7FFJl9OpPXYyyUQjlEBfu/Z
eNRIyYruFWsmBAGwCzNIW+B3caSRREDEoIqvL3C+DXsCIzey27YUmcd+aixD2Dyb20NJ1ZZiEIuf
dFNEU9sao9HikjY+fpkpkuJChKPWaDGujQ/GTj7mJ0LEf7f9l0p8Ayex9ZmyA8YgkVmQ3GGKbgJs
xE8jPpcx8/COpjVL9m3fMs8fk/+Tn+P8I7xBIsBuoiye/wz7gFQrVfjR7gjl2x0kWO93J3dqojgv
gZBgxVQL0dfW279DfkygZ7XV4s7nzrqLMvlMEcTkS/l3rT/I5Ks/MJHytXWBQjvLG8Nwuv8lMTPZ
WfFwBzroSIsWFNZLMNpzaGEPUigJ0eoztc53uVyeuUKhjbXho6yuqrD5kqzfml6McIURzAZB8jaA
eSnkenyJ7yHFm9ZjYFebFIl+wWMYGTthhGVtqzo14FLHqB0HNACp5v3QNaQQz0sXfYc6HfMw0/AU
U6kHSGMY62ercuThFYDu3IkhiwScjQh8Fymzzcq+GNrKNVItgC0cGMJwamsFtUTl8iUTt4X67ann
0gdwWtyTLS36SRvnccleBvCdn85xtKlMcRTztsn0EgN3EqGkz2rbB72UvgSteH2lmGQPWx0quBb3
DYbO+9R4YwstXoSI1D8n07F47LyhMkgKqiLpJEE2VKKVBuzDhN42TkELQCYq1G+KEzH8ZKwmmlQ+
pTFxBlu4J5UUpahvrwXbpAuX21lD1tmnbjV8upKIMoQMuI59assqyR2rnsuO4soy35Gpq4VmLSdQ
oRfLi29mvzFz9bpeNfMRWAw0VzQiDZAWrlrUoSoXuNMuDySwLyog2BcZmFNZH23TYckQKN82zJHg
moLlHuNAz5gEhYZAuTANmAV0Ipiq5FWfmOP5VPI+kjNSkyIbKprulsmt7n/6OU0X63HJVtTXCZ+G
SoHOKJkZ+6yYdOHuvXSNdetVWfvJDu4R9oE7r70IaKI8RzWZ6oKlW8nIRJ+5Bp+6f+/oqdVcJc+j
ioIYVtSHKcaAeFain5sX5S/+8DJ4nNwkY2/X34JB99VzeoamTUzGv8mjgfmAV5ouGQNkNCqIjTLd
GdvducFEQcFUMuJC6N9pc0/MNaCINRkIxlzqBDGPzrKTxHBobtnldE/+DXWTICcTcGxD8XlFu2dY
ntHvaCrAVmpx+YJxMZ8h+x/iSffZxy/xRm00aMgJHL9PnzKax77jUz443i4jgkXEne20bfxS1iru
ev6pKkUl7AAmM5glnZbzQHhT2rnBPSU9G+xgRnmiMpcGGaMgpYS8pM3zbU3M5gnov9WlBdmdHgnK
mBJq8Ci+0eJK/Mv+g8j/Trow2DZU3Tq3VzW9mun3vFWqbwEDnTlsI5HieDuxMOmNAYvLlg7Rk4o7
3sJRnafpuJuIqfw62GyRIO2Fe6YgKUTTD+etNmAv/aE2qz8SCZ4apsCOp7mgU//wFJb1m8cPXzDW
ZdXpeNKAJq2/i7vtLjNC9NS4rjN3p+LwvG45UhqsbLuj9wHuwGiwu5jP31mTbLjp/ygdlmAnOfN9
a2id6IiRFVyX7FJNaNXYNmkd49QdYn4VSauwKb4uM1pY8/po4lzohtKS2v/OvBjwDxiTFY3/bgbw
aEqSoSIF/N0Mg6DgTEhLe7n6b3CF6+wfV8hWGIwoSGmgFD/wCg6laipSrsI3fWu8JERrRmBex62U
CJzIFqjxwgW9FSgTIFAlVBhqBeWxiZJlFjwyim+gnLa+LA7mqqYJ+UWOvCGcgh5RnXopxcMS1wmR
r+jy2KU7b8qIy4ojiB/EvIxraNTPwvqW6dZedvP0bzwEI4oDV/kVZdDTD6u7Wxu/v1F5MV1AnC0c
l9tb5F48/YjLeh51s+eI9GSu4iHvLBrZ2SZTJAybxsPxKH3CLyWh2PoU1WqUDwU5I6CmarkXsqjO
mHCFDUEL+0FMe1MQiYlYXksUPPaiV2+4B/IAqszKxFx4sWinU1cS/tX5vDWXntCkDvFwmaabwWjQ
viHX5mAOpFmD108uKKFsZ9xjY/guRMkpEH8oCymyNMkOo7sw8cWYWkahzxK3pr8LYLGDZhM23KxN
c8qW/7Qb/x/MbjZpb+IAhPB9h9ksZMbC8TVHaaJa56lNdQ85BwkZD31BzAFr5DEgmtpSNqqkEcpl
iY9cinEdswQqJk+GuietDHwudxkVlGKRVgifS/o1N+A+vZoGHt7FKKQXInGOW1lwZkxAgu5NQGDe
V448/8mIxpdZbNTqJIY6pUAGohYAYgCpB/+kMkdfilD7iJBv+ZYhv6rNggWTX16G8LxWEPhvv4r1
FUNP/1G+jN5sJ72hGfFiEeQi0nccxyowlHCYFFZ45WQAhR4TThsVKp0ZPyTQmoa4C7tNw4K/k719
3Mna1af+JemauLJ29sgJaTarYtQKqAdazYxS9Z0xuFuEqjdoEn8W0vb6+fDdaXRJX5yLcGeh9ufV
EJkd2AefT8hdAOyEizNnTwZXfbSaf1Y1KlWeNYThsbXsJX4HWKhTtJ9eT99wdWBVEy3RACrfWfLt
5cYJbXzXRrj4jQm1RN/Wc0X+xAPngtN+tRQxLg4HxnRDZQmENpBqxmjV35a+2LEm//iwv8gCuEmz
HwLrcIKBTJWzrUpgsF8nELgEALgEB+GAR2qWLWJoRuEpFOAJjUyfNdvK3D6XR6auVPm5M05p9Uiv
+fcxXHTp3k0krdCwmINdyny6/oF6Ol7c9wq8pY9aDSQyhxGqMWQ2qlFADKVC3Z4ubvpJrmIUJGuc
ZWn61puK7zqCSVsE7hs4dAxg1lWyaMSX+aOp3w6KLqHHEm3M1V7MnfGHuSZRGj5OyoG6LdJBVoab
gb6ab9ugj7MuXilw7JvouK3GrK95Kpq4rLO2JAvRv4lnvkbxtXbpAr/xJtfZOiE0EoXezXdCk5bb
ejfmG2LU5yOrkDYFRf+nGo7UN/juR1Kh2aIihXV/mWmG6fnReqrDl8DWM3yl76i/A6pRpyOESUPL
Sk7mOVvujS2WGQ44o6+fFiOqSNwr/0RoUnKBOiSY17Rvz+Vf+4G1ranX4mLMRwgm81YukkHAbhMQ
3FKeouoAbydScfblZO36CSiFDPfmL5BJSOhVkWxJMc85GpNMceQJ6pTlb9MZybx5Poh0JcbQuMso
W1WvJHIAsKRgN7YgRJrgagZSU4kwJuFTrCxD07oGjPPKwoWVpEJcbEQIK88+sdfF+m9hji8sku5H
R+tLv1f7dhjBKsWa9/dWLqPZyrH6us+JyTAgAkPc4Nzd/l4Xc55CUtmNyYKUnYSj14Jcaus1cD0d
BH4adAqDbaoC4OM4J3cxw5P1trQU9ep2zAxZOGrDaiJgqZm0rWCOVmHEGpwzQ+sRMZS/jOoGOIrE
ZIhINE1j/uwC/cwaDKTtn3A234VfeEBXeX1t0x7+P2AHusrRQGTvgSWgjEnssOC9iOyyNhrVCQuk
K6vtY6dtxo8Of585W72DPr+H3o1Tvgb19XWfX59GS0xEhbxz1uIg6JKGx5sibvIhTzbgrhgiR4JD
V2D8bMcd/tfOfF66ahKBTEw7vbRNE3qK7l2ieg7juJLvhId7N5KprvBO6H90qJM/+rQOJFw5TNWc
P+riMiYRONr5ntRRE3ScqBLGyYa9Q6s7U7owpAm0t0EBw42vXYl3XvVq4LuooYRWWC3mUlrlV+K3
obO9kq9igPsdrkfOyfTnV9OLdFrpcdtFJrmTREOiqoiMeW03XXR/TzZOghO4lcwrDrxVy+b7ZuyU
fa/gc5iY2XXSK7iK4ZWyli4y2cHWwZYnuRw8fzpJsvLCpZFIZ6NcswuxWFfc2KlyGN6q240/Vlwi
TrEQ3bILyezRJfoTxVk3sxzS0a0JJwEL97ETABhgGM9vSgLO2OAIWhsR61RR+uO814zPi0BePcrl
e8A55E4wXunst7xabG/yQBIuqUjJSK3XbSWGZsUVtrsuBYI+ryZyDuSgs28O4XlGKFsJkEJ1Foxc
28q56ZJet+s166Pw8HO4Rpxb4fKbfJg8YjEW5jst3Hj2yzoa//HF7wx3Ea1FSq7C41nUBuEc1Hg4
NYw3MgZmKyGWi4zXRv9ULn2cEoqnBcxh/93NOI/8+hS3+WuJRZWc2Yq/Hdo5Gc5EmqZtEBn27QpF
fH6DZXNH1+E4VZdn28GqyjrKuG5zN8k918DP6bx2/PMIHWo1dettACTKdTxbKbR0GqrRAznKvOZ7
WVlk5WNvNLWLjx5N7bacm3az+Wg1nG2dHPT30SOjH6NBICJ52QzrKSl5704vHdBYHERuG1lAI1Z6
B6/TWEOtCuDBDaA8Zrp15UbxrPMsvaa399+mojmeegMTWsUZ+0epKNFFynLPaL/BUIKix3q7sQew
3E5WsgnFXemw4VXnjCWb6gTa552jLSpIx5oqQLth+busM9E8KupK1YI/lqq4vpMDzplYV/UJAxFN
AovPBHi1ZemQ7AFtD9xqmOAwAEdczBfIUvQmjFQQAhwlCawodcdbhp/BJ/s0c9onGJL0pmGwVZCU
zLh7jjqC7c1x51ne3IavK1PoXskwyxTDEot5vULIqgLx08O7FLluTrkWqssVm7FUQu71Z2M7zQpl
62je+Qc03tJBUfhRa8Ya5fW6jbDRTJUtur2AE+WZb4tSpqe5q2KFpFkqv4/tlrVckIlE1RnTj8D1
MA45/eArJbwodBWGspCrZMrUl/Jwp1mpbNYpgdzrTA5uol/HaHsCsgUqON7nBaPjRmN1G/t+8ODX
W6FZwSSX1EXFtCIdCBNRlb3GwobE4FFDskXbJlz14LENdLzGaQwLGeNozfL9IREMK6xfX1Cad2V/
XtNu7C5Wkiw56CTQhKYXeuBWp86tb7wfC599dTl6Am/Lv1x1zwTDwyXUjlEa33Dxvs5Lhrfa49ky
mY/ThSNOH8l5nzExpLlEXu7ZoUOAYCY37MkAlF8bXtyzmCsyt4yCiyV1hHJE2Or6g+/I35WtZlxd
QpsCuf7Q1O2iRgst6KkR2OjvpeHYNLyB8oKtfqnaRt+pep7wZtuJpvpbQUa0Fl+3ZKEV2VgBAInL
yl9YVwrDQPwud4CCuPtLtiC1QcuJ69xhqviqAUtPEhceppC+4XDgH7M3vOKO5F6KAxGtug2JNctx
LSVBuIBkG9Cj3br0dTXRD5cpsDhadtWxuJaAXEOXkp/nCuzndvrxurHxIcU5hblUvWTsD27v0JiM
FYT5B1N5CaTcliCJHgtLJ9XHB5fd8GUN+IVxm5WN+h380KL4GmaWQ1kPKE4yMLiJfocfjMutcMO0
UPZ+E1qLvAaI7ySDm59MiTQCLP5OpISk6NfOW2aNxteJu7BJ6VyzpDGAPSEY8GuMbIkGxXdKJRdD
jEzXcDkkTylmk3d0JiAQSW4lrsLtJN8Bp/QtzuC/jGQoHzNYQ5qy2OTu8w8nandPUssjvSmgORra
vwkE/HtdXFtrGALu0VaSSXdYPlITSp4Ey/rPOffaTJLtJsipEeit+vBj932o6w4LbM7ky4xLg+Vj
yEHyb7ICmUU3lZdkwY3yZP48kSj8/5t0ZOPv55N7QjDyf9VZYMGFxwq4jb8ZJ1vwJefkRg9C+z78
Bq/q8WTP9+0csRVd2/hh2ImrvOj1Xl+BvrVJ5nhhIjilt78Cx64mRjTQSsC9C6sA2Wckx14XcEvX
vQ4Ht4kHPZpNQDlvPzkdaaj+e6riH9gZ7uGm7Rmadoo3+JO1gCpjd+3vWNYonN/YXoM/zCrFyH0z
OI6um89AzWlAIzldczWlZfc9BTh4AInQqc6lvCzMusxeV6Susa13T4LXfnE5VBfiGR7Y1ckrC0me
Di+PMbCuTfHwmz36Vm5oHky1X7Xob/JpiG9le1hKNWX+knCmmuCN9wNjQN1PGennLRNFfw2X9Zbp
GKGTrUDS7tFVtHgHECMGHwxUL25KLrGK/HEy7v7hOpTfATpfsrhkigxwsTfwUxtbD/CfeSGWq2/i
vRdly8CFne4Wb1ARmKLOg0eJm92M7t2DSl0BlzfqejtzT63J1sETi4OqkKztkq9rbGNH4Po6ORS3
e48GcIyIDrKvgx/JLjlcTL3ENnNF0CV5eu2FH90FOS3D+Hy6Dyq1q4e9530G4xP8WVY72RtpBkeE
vaRP52caD2wyCPPh2nqKM3I+5l6RVde6dCIWmfQKA1SA/j+lWbSd5vim5EtTY+u3kxPZBJUeHHwj
0HZ+H2FUCOtGLZv+pudgrX6ggpuCgft+w+O51BjYm3EXSGdihZrpMGvg4yOfs39DDkqrJmgb0Om5
8oxfxhcuwGk4pQ/oPSh1Pptwy6AOAToFntWng5mUauVnEeTv4lCNddRB/YJHRvh8SipkyMW5jATZ
Bte5UsInbIdC4LKP7DvJMnsIyXgSYte7CocP9IrpYA46xTKnQOCGwag62+tiPZ5/WuC/iWLR1GDG
Ztyp03jiFU/e6HI7XOn/56urnuOgdo41fei7e/TvIQBw/lC8WLcZL4K5KarNELhTLj4ByMhyL+FX
zsjKKL9v5f7s/tEdzL4LWTFh/5nBo04fG4+v1u/52mGXAuFduEw0u0kxuCV6WEqk7YHGKr1afPDD
ReBD5sJKD6NbIPL+qrGCG7YZtrRXOKZfKu1KQSM0K2WbIlxMapw6pxcXIPYko/lyZq5VsdY+dK//
Kty8pgzHGexm4miGn294fbA4FE9xDy0x+Tr9kzThjakTFQ3W9lkVm7BzjcKfbJAhGYkmpbjvOzSE
EpBemrSN0I5vy9hr5FC7H4sWY963mWsitQs1m4qfbc78hfENp+M8u5Kct3AsIbhJNZM6X2ZJrgHa
WnB5Rp20F+fJGuKuYpMjpkNplpX7wfQeXcMicqX1E+kQrrQ8QWTgjHzBEWiEjbL0rco9p0+FueXa
6lzwHkv9OYlO37eGq7nYjgzyYeHTbx+c+jH5Wln5Oe3S7kJOKcK/9S/m1QyIFu1DhB/ZZ1ZjatXG
NgNThPMsBFvXul/txLqI1D/G/TpGJmBUYMjoNSpAN3mBEVQMlr/oH3pjz8tiQg668XoumX0IhHD2
vIkpKucZKy94d/RPYZfuE9W2tWSJgluVgN7OgpeKzCaWQsfPr9vaCyPbr2FtaVVrwfKCK7yu9WvJ
5emQ24VEViBAwBwq9wm29t6I8HdFDKcmj5Ci6Q2PWCiDsHVRNoQfp7Bx9QrqDAZ188ybbT0oa/Uv
vqQSYQrZAVgespzrtTO803UBUNIGrqBnx37vuWoirHVGZ+A9uBGcgJKkzc8XPtvEMT6FqfLE5/YD
SWUyabSL5GdxqLPu42XHTjawr/ZytWHUzjmfoA3b2foun9sTDNsawuQQslpK9BE5jQCpkzsGHauW
AtY+MeJLUN+/7BGeGKDGXt+P8yoF0Nea/hIcMRTGb9fnOER4E7USHJkMwuqABhtHVkol/W4Xxxa/
5se7rStVH1gNCQ1lfymER+i1s+CE45wFz1ojIci8tiDGbMpCOzOfxRtSDW18Cx0lKC23CAc1M9SN
VE099+m1+AJoQFy+y2NxuR7ZOiCCFTtS+urfAvasPLTqsuXzjsiZ3DY1Hb2cGeUkMd9MVLtLNnH7
v7uRE6Elrw6zqK2vrb/wQj9KzUG0AsVQhnYx36cdxoAbJvDFblhWCZawzqLSA9V7jERLgIqhNmwd
qTMc5B8TZNZPnteCx3ZVeBBisq5mmpJULp2TZiK3U4A5iVUcjrMcAJVgUZ9OojE+0fLg3cr0UyaA
vhOlwG0McAzsbSwyaDw+0s/3MRb14uD/DnqvYZE8AtEhYlm8e216Lv4qleYuHJ489Wtdo5j1bfa+
dqz3lciGepwGUPzsDWfYmhSA3Jd2CbjX+RBxe2rRn0LxyXKl03H/y0Uf2M/VVqUWQLuY3mF4lHv5
xzVIou6EGNRxR8me3NvDQpl5IFuUOfHMrP2OjbA8egFbjzSHKmSbxPTuDQQS75IkBTAZcB46QEld
eefn8ECIVzski4dliWnc0FBVOYPjxBPiZPPHwBXE9xDlumdxNo3A9v/fHGwqmOJb91tY09WaU+CX
0yPvbfsziX8SrBK7B2/X/dfCT0z15Zx4YMpQpLgyc5nWMFIVoRKHzEd0wUBBt/pEFduHojVt2i29
ao3xF4E2+r6bMiVqL/630VLRQ4ObBEA/ZYZq4WQlQn3AQqaeDLoLjX7kTvKrboT4m0cZAJ8n2jDa
EXtu2WHYPqFC9AIDuUFYocqypDtKBa/lLNWDWd3SxQxau7Ob0FKJacFEr7VcPNmYe3ikzkYIjtzn
ANavmMHfAheqodbnhr519rd7fAPz9nh32EDP8Y01jJp9VXD1rEBxG2b4stsd++pg/9QbkMfBRvCi
JBJm9r339Ab3v4s6aD3vNCKs0uKhLakXmV/xdWxDSJWgreOhGDlaYLhk0lTtWrC/+vh1dkXoRof4
e0PmH0LnVpRnXsDI7TUcPrQV4LPzM5TIDZfIPH7mOzK3yHwjjeCdwXms9IBXVCOYVPZ923bmh36Z
NJTEQ+Q1FxocBTgGznQ04Ma9v22qoKToro6FSwSkxnOlo+esivSxw7tbZ+cpuTWpYyBk75vYVG3T
1PclsBTLjWruh5Z5m8vA91tvTeJ3bWaGwMQmqXVoPf+53zN7V4JYniWpL3OxiUwzaIbtpqU8G8wn
MpKaF6oMZ7AgoulFSpdHwU7/bT/UtB91i9GiBIRsT3VcwsSXm1JoTT3D9RlD8QG5bakHZbP90uHl
d79o5OLKkVPh7VGb8BfVeLoJWlHi/RxvXsZZWtF6tvpNsTZVfi6Kiy0uccp9q1AUabIb9ta2m8EW
TLZojutF12Zd269P0lya8JHgKySBnR7FF/2LLuFKMrN/IH7I7GpK4YnGBguAAtQpxNxChB88LfMd
BFGdSjMn58+9BLXxo19Gv9hSAwKu3qHGP4Fr2KEyY7TjwShcu9XL0e7zEiAy+518iuQLKgdkRFbP
IpfyCO/YvW6btzXSGBdQkY7ke9YXD4zfp9XXtnwWfXc7nIhW7dQAoDWCSaE0eZWZgfsjZzkLQ/hY
gUhDsCziGtrVTvivv2xQ/taJh++dP4VEJeYCga4J0HjU5PfBxYmYtMYRjDaBR0AVKHxBA45qLMjV
lOKfVvNcZdj+rXTxED+4gpBaSjChyD9RXvzHogN722NfyN7dIyhl4n4Z+6uSHGkxvSaST1ZKDggT
K2NkHK6MNgx21Q01DIZC9xB8nnIz4URP35iSplVWO4GCjLyqpX0UtRoiXWbRg245L9CHDSnNwq7D
9tPASC8EPJ7fC79dW2F+NAwfpWlD6UcljVqxQQpKjXmU38zEtSAXBDw/1U2IjoILG/bSbVMYjZeN
D7F6AP5ABbmxdHM/2ql7h890eMrHpNjp+tYRkFtLkAqurdK4cDyXoNRfhvr57qe+BEaVMoPhxts/
Mz86j5HkbJYGNDXlaoZiVxTT5LmpNzN0hSdBZewLwZYXQoghRgVZaA3lqSU9Y9S382NrKqhm+uf6
wohTlvHVVXlmxYyh3qy1jzIaZZhdwWsXmvD+dbdfBX1OXKeazegZkRRyPPwSBAoYjoumNT4irpQk
e7YUxxfhAndXHacr8GFPdJiKTRH9wKFEXex98mVaiqrLjZ5dO25Rc9C9dg6sK2kN/8ThXSIPo8+U
dt8Breof9024qT/EUbzoASmL6R1w4rLo15fd5BHRJg10iQiV3KTz23sx5Szz+8bR/qD2UlN3cFxr
FQNVjtD0DW7uaGquVGLtjs201hYvB51NRUlfyjKqQZAeTGlRMn6/yCcjL2VwvHgUevhgIFAkcdZI
/XW+mmzoWz5MZmqMYPzxKsqL0NIwWTSDlFd9GabUaMs89cjdfgNeupUVTXsXCc7octFumZ4WIZYe
3hOuxB4UQcJ8tmPjn+LNXP1KGejbPaYEOE9CM5ah7Gbp1HqJzVlllqdToa4TGVkji3J1N+9GE71P
TUy+3k7ro2/BjvuGvrjmD/cNk9aC52Th7qZLkQkBl0aVVwT1zyeStu1kaXCcAqYSKabFyriRFpha
NK8tG7oWIsLyvQG1qZnEEYpv/IKp+FFODGhbZAX8+QQDhxkEd6a1GDA4UFH+DdNKstVRLp4tOuuz
05vdlFfBUYrsOgCdwZ5BwpFvEzWQKMb3aa1Xvu/QxRfxXB98kkmvmeFa8Y18tdz+3wBlF5YyDYy6
9q383DbLUBxiE9x4AXEWwlJrtlUgM8DquXvq08JsMpK+F77/xSQdwnjTOJj8g20NvOs3BftDsSXM
/phm4jBp2KyAFDvXGWkODz2vquTvv2cayDv5jkPXLra21RLX/HHkMM6Yxa9WOXQYz8FsSjyIsSuO
vUWH84iI417sSaw6vdxSuvZyvg8YiS8aOZTG436qRsjt6ZhFBBEIhTD+G1r3YNbpMdpUmJfJ5Cf+
5v3g6Vrqbh533UynvW6vBIaRnkZfMu7kgZOH7U6hdss90aHKwAbiX7Qd3r8Du/wi92D05B+qiX6U
UXWnpEStAW7RsLwWG2ah1uD42kd9WkvKX7TIvsxSjbI9HdbLvzX/kYu1B71JP8saOZFf0qhKoWOb
lY27leEkWLcdl7BQOjJIDoFK+xusn/SQzgxBgIWj0menuMVHUajNcY1Q8G+AK4KqB1XK1xUsssvR
hzc5DpI716g+GoBdYqqPdTegZ8aPrOCRNnukB7/OHZ42Q+R+PlI7/VcalBZjztQLO7t60OUdvBKP
CMI70YoWwEzOm3bRqWkPAkcHTW355RpsH8ao9BCg0Ks1d3D6bVxiZg+fcjPzp7wSzBp2bZWbnnGG
EDJh1G8GMffP0j8MZmQnqjgdMKpAZzQr8HOZ6XWaUnm1wJyX9fQ8Is2rbKDpsQq8MuCkPrRzsfr7
4Rd7kHvFcEroQ4PFZOYmPHLfnDriXh6R15k44DZZ+RCNbaB/5PgAwv1DaYmV+8BvQN1OMzld3RfI
AknTiDfj7T/1DgjkenDrKzLQPDjn2tIcT2x708O5YnjW6XPAPWgGXSgCitbts/Ek5atreHyilG/X
akZUSkH8I3l+Znp963QOT8dulEkR6SavsjJwVQpf8qLGhqnpTxI4X0jjBICnmukBtsLCxBtE3pjI
LWCXE2kmE6OQP/67ym0713Tothu5q1rwnusThfo/UkpYPX0BdEQZA8Wbw08irNEVPC1tpt17bTTI
AGit7nZo/qsdQYLvGxdVLY4hDdVX9Xge1mGROaN+nVcQjafTdOSqlgZgxPzAT8kK4Ex83Ubutj/B
vClYfpusxYQLKRQ3+wzTBa2NUwMxDTG/prqFZb1x6EEGPMx4gpE0IwFA1xF0tKdFpMdwK22o+Z0u
inUoNFr3B7uOVFrx0QKhP3EUZ9Hbk8vVdGvcou6hWYtX2MMXAhrRlqK8Rmjh6pyXg2kbvGbRZUZV
HWfznr8FaTbD2wijy34fHd9RQtP+S96OGkin/T7Lwrjw5xAgQ20yA4wuWTNWlqGjg8xnx5D+eCjb
7Sb9Yy7gyDWwRM6lDxSLCfIWw6Tx/EW//alaqSS9j8SDu3TZw/cny/j+HttFc8sfrQyM60+O93uB
308sPemVkxnKkFMET4mmrLJsUOaSD5ipf4j07zuKBSo1T8nxZbXINRlNOW+//McayFxjFMCniCFt
1KlAkXNtz7rAndGiMTbz6ZOguz6F8dINdOeizggI3DJuxFBNoYxKFSuvel2zoBjjbUvW4kggDuJN
I+mylg7JdyVY1zBGPyWm38k20ORCL3uFV8zrTH7b0TAdMcOrRFLSAOW9TqnWO2Ehxa3YRFtzVcQj
vErxCcj53pzStLp0EqhQQ2BSxhkOThtrLEk0ovbJoHUduliCxHg7W8QPky8baW/WXKvyYNwvmy5A
9DMwCJtygJtCbpDZzuTNKIbMTHsZgOl57kKZiOByrVzERJunziz4G/eyZHgLOuAD18LBjINH/Yq/
xTsmh7RjgfCU7Zt0dKwoHRbkZwbOcVxXH71QDRokP0x0NE7R5asCPmB8flLmNVn6XMBIXG9ZjwtV
jG4UtTN5Sq8CUYW2e+AxllTUrfBAvLIgDbL+oos/wULVsqTjZrK0UaPSVIrvoFHJE2BFB9IyeLWe
UWno2J6ZOCt7w7WsB6AqeEjlQ1HxzWEa4e+PmH+gQmlJlYgCgxkJ7BRyAWOAqnynQBdcQQhpMzzu
5XY4+ZJWMWKPgjNqXGJN+FPJwVJx7pVGX+uz7FyJ5rBC9+aCGcgUxRfDlwuLbFPWgxfLhATTkhdV
YZZGspL+n+5ZzpASbqQ+kWsORxHXMehQeeZ7ti9BE+qwdsRT+h/UXQBB6uATpfjsUKGVu/TMzsWe
zDZn40oCdrT9F55D8hPgJBuNNnzICrF4jlStxIiMa3F8S+DiP40T1aerAIChjUORmHhFkX4ET5Nm
pWmpcVe9PMAw1oBjmtMHc35erREme0Av0iGMt85MrrBFTSdWRQCSb468cadJ+u54YeuASjDgnlez
ACl9tDEKdOYfudmyVbEohBVHwd0yMjNF+JhppCjrB254Qg3R8XR4RgoLLNZYnZ4JWmW1tTquynj/
quW+pXpapVStAffW7ESZ/8Z+1TV6/STSden0/AZK+otwOO8DG0QNuEEG7Af5wbh7u1CR154jw8al
Vh7YHBCH6jVIMQj9LeAkywKWWAcIihGVfpMwmvu9f0bqMNuQNkYkGWx6m9YGDcUymMUNY2/jsN0i
3hdRoQ1qemO78ZsYbvZXUCwJeImc3bGek+TDhZyZDF6JUB/tyl6cYVvyMTFimCFaD6jjk7Qs0zD2
zBonYbcPF7JPKmxzYMZJg7Gami/wK7+3tRgMdgKQmzpzcMy2cU3pOrawKHIXMcgPYUNL3Og++Ijf
MkRY6XethfIGuk7lBO9e2QC79gUY+gpSHiwuoJ777tWh7v6ZnupJHW+pGWbhSbr9yaaxiqfpXWaM
qvgiZhhTQGmouqxuyGN3MVzvbl7KkVZajtYY6fmSNjdrlv590e7bDlYyU/jq69a00ahUuNj8dnqQ
dOfxgdoIO02ztxs3maqEw0PjW1ozEu1tnkjJSMoMMqroHP2aA8GhORbBvB8dsfX01FB7ZTTT4KxV
OGBMK4CEfwheImSdMGrRzgLMdQBvG6smLoYXJYMRWzwVipTpF/08lfZKl/GAzO5DTRuB8j+/uEOg
KBtWF2ZZWlgFFRawa9Vf4Ovzx9A5FOtCNIubc5RLVjRn4FWbrlt1t8mcFc8NUeSlHf/FiWstMIet
lW/P+VFQb6v5xd/dt8cFkKauR3sYjKuu88Jt7gEaVzmS4hXwZcnF/qVwwFegDLsQD8PoND/l34ay
400Jpg6JcgxZFWJ4WuZOT3ygMD4WyXmhIaVevfMx+negRmOlje2E2FmF3HF1K1fI1GfsHmy4tzFm
9p3buBNZ/6YU9x0bPpBmob62LKdmtiaZdqA0SZzoFu2rKBYkorEocteGkV/1qUqyAu2zyLi7x2Nm
WYhDxwVU2icM4ooqXOahF/i0HE4gpF6O3y2hIAxgIlljwAKYp7Qt00Xc3nMjGUSG+CZCdZn+L4/o
gv7fJ2mtdqe3k4YP51RbX5zsJnIHIvY4+q7JocAPmJhC8/SxvfsS4WilSBa2/bEM5WqsuIh79SF5
vCr9UA+WeHs3GyGAtEW+mFiVqZc2cfT4TpisyrpZvugAD0gibqW11hSURwwFFhp+6hTfBNSUaVWs
6wbuAwkxdjP/iE9FJMfXOEwa6SXdvx4Gb7PBsCVhj6iYUOoryamm9Qp4m3gowmPB5QVaCU29M6vX
/jRhCQCFCmz0Sc+KhKCKIp8gf17Te9AxC3a8DDO2alnIzJPVVwcaKQLhnIm72CT2+1Wim0vLXLtM
NClglIhgau1XSd0j97eRqsk7+Wbi8tX3C8RmtNP4yS4dGhwqRDvubwfdVXV0vtLc2SBl3IPXo7zQ
8aZ9dFLEOznJr2bHKSyhbM6s+F4i1pDNUS6ilazE5QFxks9cCBhwSMgAHLLAQ3yg+cYx8hqfA7m1
pJTB4s/7rHGF2z8N9ujuIOo/yXuAao38z8OQYHzaUBmJpl2j4P5Lb4WUpgXZ6U0cj2iiFWxHdnf8
wT73JqGjpx/0zQNeSwTWPPMzn9LzA87mImdcBSM/2UZFzY0qOIekqWCn2cFyrQXl0GDKrdE9B5gx
ESvZo3BnKwjcI3Iz56XKfQ88AQZYY2yGRusXVdw8XdeFjuEHKzm0ML5vHFHLuGYsR79S2fQSv/VH
DQw7FccPenzOF4eKjJRrnOuc6/uB8mD/RJ7ZoSEmRz9nroflxTpv8HcWzC0AZS+IEC6qBFEFrvJe
Slnz4v9eY9V7kGIfYVwhEknfPpC7PO7CzTLAvjsFpLlE5mnuYAIzca94r8T5o/Dx8RjWvgJq5GGG
CGM/ne8uohL4QrNtY/9dpmck84kgDFrJxE0ZZzZTNc8z1PkwXOFw0QSxhj7soj9iY96c3d++zdp3
uSCoj7z5NWZjehtA9Sq0fESZRIx5fqAoXRSE5DHDFLRn/6Okw0VwCfyUbzT8jvCImQVcL9l27fyB
YMD4A5nxA6n3C5aXKH7UkExP8OVqgoWULQZ/uRacRKkmpV9UalRyHI+HtbTjmwpU3knAPxFlwJnK
6I0iusxFP5pXegX7VpnxeeQsZhkQRZ5HSmdrhF061vzQfaUKYaKEly0G5WOokkQB6SdwEgiWgBV7
WV3d/xjPEzO57qKbjrKWHOmTAD80E99kVv2NN8GkpDvsCjVMuikB1FpjaYan86gdGkANtuwTQCOY
yfK6A4rl6XEqdTRbkG5PQU1sO2nNAg9PmqUKkgwKAOXAl/HzOuqo+YHdcTG/uNTmpHpxfQUk1CYs
Iopkx94Hdia8DxXVyUgX+UMpQzA0XsNkXebkVw6IKGb0aidPZRWOgKFy5d7PzdMF3ASzP2E5nyjN
rkgOvxAQ9pJt0SNqdMRGs7it69/rwi5n9z5imHqQQTTpnvgOIZfy1FfmC6PkoPeZrgM+zN/hzhrW
VrXJQ4Q9smfFF1vc+ERxEGKrFkm2Mcx+a0JdNaQulV3WN2XxBwfzbkUa3kzix2bL9PFHXDhUh7cd
i0rdtmlnSi7ky0kgNoPQFWQLEQQoruVK/P6NkONb2p1xQ+RsdDoh5teUtwWBCIddMJVTX9nSA49T
3lHmDoyPBLhKCR4OTnHO1oOwfT6D4R6hM4bKEHf82G+xmrUUP7wMazZN+i1RzBIKDr6L/5F3N5At
qUgsE4P0p7ig9RADCaSRLNk2j/RnPlyWfmrMXyP/zkNKaN+mCsxAZTKZWXBOo7wCG63tkbQNFHmD
Gmwh6tZZj3+JD8IXHKct8Uz7z8HZWFITNfetkc8SQq/mvRHPhWlLajI4FMmYIm6eax4pqrMjvxsV
zUNGRwWp20euMclNLFeBT+dM+yt0oO3J0AxR/t+VgumAiVQVzJeSRsl6gBd8OKrjEJQBvLqhlvfM
nOOhIIK+ONeu7WGw9iUA3fmqhsT2lM7+WxOPwGdA9JTUUQ1PztTsFWoX+5YUeoPqMdI15imCzf+G
/PYQk36IR/7e9LyAc7x6jo1xdpXbAJFSueYChwH1OzE8FF/P1k/vwfYELltlkJlJFSVRL9L/7sM1
VU0+7qa1Aigt1BJfi5WZy+giz2ADcBhynPR6+ADerJHqPe3E9usyC/Bi29GiC6+ZeMyRxnYvSA71
F+uTkj7hgf1ajnDAImLztx6OHsLEqIzXFvEW3qimQbXn3IGsPzTyIXD4VZ2MOqNviF+pAT8xcYdc
78iBV5ArEQlHfW44TWIHnjJy17Y5evw1RiEttGj88famr4Q3zjYkvJw0U47LH7UxJwKvJbfTyusc
50D3k6EpK20ixCYDV5+YIsd/vq69+y/4AmvyvYeS3zFdbskzNPJEJUXk2pFY2rhxY5xfXkAqTbJh
I7aAv2dZAmU4weMFqFpGzZY1886bXrVij2NYc1HOW8y/f9dZXDKfiuH2Jh6wPgbqc/8R9fRPK+bT
ZQMmtiS+j2MMmYTpPof8XpbeS0xhFIpz1aHPDSAwmQPOBs+JiQ/9T5qzoEuQf5LGAjr20pfGq5iC
uXqLM2/FqVWAc1qfYy7CAOgb1PhckcyBNYxoGxccqdY0GnL9D9O5AePDroRE+ZNtbQ60mf5mi//j
7hijyEvexhRHE7A121qgt8HnewNM8dGY+vONLv3VkdoWeoZR+pl5eBqEByvi8jlhC0rRTB99Ysi8
Oes1BTQXvdxm0RZXYdqtA/dN9jeZ0M8edcmAifiHZjrqem0EbtKVw/y7x+ZBDMi7lbRhB20TxjV2
SNX677IZrjExy0CpmOt6ae7VnxY0iVlOL61J7I92Zuo4xJlFjlNJHSoGyguI62JqD6y0SjhtbJ4V
t95Edy7SUPHqFWVUMDGPUFNvKUa/kHFETJd6Kp/xJH8M9FfrAkSUjq205SfB6W86cw8mUh28qE9L
ZOuPv/I0x6HiChQ8U+2cfIkwHNfVbR4m22abDKVIK7y6ZitKJxYuldTn5U91uJer/4l1Rnm/3nD8
X0v9UnYnNah15eNAhw7A3a0cjcRPIBNx7B4gauh89Mimu6/tiDs6HAludl0VSOZw+HMTcoQwwZrW
SVv9wAiAx2PLj/CAvVTUAsoVTe3G+kyTrud6dOc6fHZs6Es2Ee5nvEfDgnLoLWzkSji1QMrc5AcX
By7eko+8XfrAHBL/cyNWekr/pay+dx9KUUQa0XEosqQPqjfPDMs3DKg8RSJ/aLL41bDhCwU+tHkM
teUvnZTxvkyZOiDVV0KZH4jIKI35nBjseZC8wF3n7xOe22o6WD8gE2TmAqoXvdGzKEbvhApZjSxO
+vvKsCj/t1klpp5wTIwOpeSFSyMXMwL4Lp14+bttRT9JqgnK277KM4d6FGbt6BpbY5wv+5aZhzL5
eLSWBJWtDyRaDMbkzqLMf2w5Rua11OxSdiXmHUzTwzuMiHX98vNygBni9+eN8ygUL9FKUmlQdH02
AkA+ffsKvDBG5uRDY+7WHj5WoJAfr1VOALN8Qls1/a07J2mXIc0vnMfZfM+h9liiMvkKRWTHaous
9a+jzKzEfMs/JuaLnv4AIEAiJFzK9suSGgl4wOCMEdFmkAJA61OmI51QQgMDPD+p7qVB2yPVwZaj
lcgct5F6RimayrTJoU6gtPCzU3+VkRxnXmkcK7gjIrkCfxoagQBR3RPDrzyANN7exo8g6ltPMyvh
w9jSGm5qUJnID0XzHXtbUlg/7hNesqTBuftrhWtmBov05M93MW4CtYqFeMybE5hpmzO+Ql+eHuwT
kBurl0cDe3ghjOHWyOuoihGXnrVQiECD3LuLZpZWrf5EVr26ynI8YedIipnMlszcvr/AZM/V+uUt
bf31AshgvdeacrI6EXq8Wj8cyW1U+NI33hHthPdgfjipN77/ui7xnLJ9umIuUTbkETVGPL8vQBPz
TYMTDV/40OgQYpVtK5renD55hOtUryEggeHCooWS+sYftuNHGDD+QdXxG53/fafsUqotPnBGew8r
Qfb09tlqWUXxt2osarLb824VHDxzpnD3UUJUKqjLw3A98ftes++mHXMgVN6GkXVBoWBqNbh/ucXO
Qx+vR40uybeUf3i2pQCQwwaX7ra0U6C9R14ohKx1XmBUteQW7iFORjIRpMfQOriudMCL9Rzv7IeV
UucLstRS8aoOixSULku2bg51hzZnhUuF5ov5r23T3O2X+N2SAQLu0z0eE3a340KmAqX9LKmqB1OH
mI0hxS3o7/aPdXW4lzY5D+DfMyR/CRB1bHjj8ht/Ee9JJO74AmDHH2bHQpJqzRw8WvQwRQgIt4bN
tVDbte/oCISBl1/x8Gg8S2IaFEQmDUoPe7AVjmi2mc2V6vf9dY31RGgukXMZ0SI59xYq9RozYGO1
QcR4Y8EnkvpY8TI/k4r0qz6umWkNc+ZWRgUAY2EHfOaFYLUpT+3l0uUBA5bwM7t8AMOZfjc8HULe
60j/FER/+uTubcuSFB+GPepRT2D0e5Y23pcnejXklM+vT6vzrL+dSqDou22NOiuVj0yBHi4YuHx/
JRV+MEgcMeugzD1E19Q+IxfkFih7PXdZka9u+Z0uGEHWFYZsxtfK2KCY0JF3xyZoJvvqZ3HvkhmV
6nNld0qDfj8D/MqsfgDC4RRFB1bET0N5lgVuvcVf1Q2AQVuDUhU1KNWGfm47XFYxtDYdj08Z1NbV
t34fvtWlUa+s7w/35WlvWgQTRBARvN1oRqvDuocgincDt6z/rYgYSkjrzbVTag+R+sfA+lMp5pui
c7oGFlwCHBXUob6NT8l/69fV4xxLMEAdR/Wl11Z/hKl4HvIDRnM7iq+pJ8Ct91olPVZSQDEO2aHg
o8HtDfRewpInaK6cLYCT901ET3NyWoOUj6PfrUQ3Jhn58aH6gUhegdHFXWmOPwn7bRSGT0weZHK8
+3P1JdxEVi5mJE2Sgk+F6GlhF7+d8w6W1PMLaOZqyruYaOIWlygEjbzs8d9XGNcrqOH/Zejstj3u
NzQ58esuJLQtyHe8puVaROxOQd73ydbmORpXD6MisOY/Blk5iHZxz9TNy+0fQFszIwI8e4vWZBvN
JkKcVZfQAuk26t7NtMjL8Hk+YLzQjEc9TMm5y4it/R8///Mr+zYEgbrGOSfIg9k57Tj9lcpTFSbc
rJJC6Z7ZK93ZN6hoth6IAHuyGzu55unAPXgIJgUhLC/8BWIX7rjJDLaOijmEOizv6yPzNTqcEsv9
Rix7HPRYncB1eaUTq/pcTeuNfhfxWOH1a0mOkxt3t9kwmVF1zwk+56HtjyPd7m/9UvHZqIwuo+X6
aUNoVZ1xpU8F3C7PTsb6qph46PFMGhYGIsYVgKf1gdRGzeWNa5RMLa6+pcZN+H6wQkXY939zkbNs
OVT8xu0MJwxVM4uYHD0c/fviI6979amV+UY4p0rOgqbFr59bN6pkRj+cHwdTkPc4aB/1WkoYSHCe
b9+pOLHXe0lJxfPN1VHSxzobX4rKa2fn1DGtDJKFGzLVLQexS12zEaS2jkhJLDvrQmCzh3+1vyWt
4C757q9HziPfH5K52/2gxfMRJgLcN5A+GNSudhng+aOiCyaLFPVIrHhxVZSMXk//HUWKphRT5zSr
PPe015H4J4yPLDqrwFlWd8J+77MW76vcAC1AdkImSsLebgB8GtgR/FHgAM9qBYwBeNRjTmfinFKv
pk5RiduBK3sFzcEoJ10YKDtyLnHfFgOSDvIvoAd4AxmYri6vnpilQnld1vSt7jIgKOweT+dP8nh/
gDkGK6f7dkArs8fvwj9pt9lJzVq4n67iywbMQDN3GfLpWQGTweLRNBbc3E9FpJTCiQCSBnTiBViK
bVhlLNBHdpz2qYjUCX7cNT3P/pcK7Y+6A+edzILqCFWp95timCRcfjVO13t6GOOldalrolBUxANJ
+SxLM1Fw+sR8iSOCGzqlA1eyfo5fo/ogNXQdSJJdZsvArkthpudTbTXIacpaIYqtSzTvs28w4oOq
JR+E0ud1bkmjLhbpWhVR+mjRewkWojcGo5q2h0x8+OVLmhci/iL4oMdQBGVREsdOHxVT5Ue/crrv
4ZyBRTrxhI8Opljg07GEmpW9X9Lx3Op6kLt1N0Sv6rZCZVMADwejnDd9vaBy+1oHau3s7enQx15I
reKp4Jqw4xqzgnrOR87PADsjjxMPxxIoQt2tR6ot7jw1GVmF/jC0oBerg+d4ifWBDZ+VfAZ7zafg
livYeukdMKT0Qs0fSHUVeXCq4zBaVHPohFgtqdofpuIFEDNkYwcWxZfS9o4mAVT4t7Lmyff+k20i
PWS8GWORTYEqgW3liQCKT13HeuHXUcL8XsBRnJOhCoW6RS1i9A2YO+R84uiGD7zS3IRps6hKSSxJ
EcWLKDzVi6SIWmat6yo0Dk1FDAm0YtcLXIxp1ikufozZTQ3ns/9oyxiHZewjVrFQA3I30+80spYh
95D2FbdL/tjYdWcqGlVPCoKFQfn43aneG67wtAwCVE4cYCNTSrVExiLgu3AlmZ5k/9ANOOgamIbQ
Q43JOyP712LSlT91jhbMMpmwdrqBstaPGY5CZGz7Fbj5xA85lA71tjCclvPC0HoDZ2Y4iuQoMFaf
THFeujIoqnXL8E7dyqvuyKBsSWZ+JoD0P2ZhKasjOu2sLWVhmgON4vKzx1b+0s4d4OKPK/V1/D28
ONnX52K0WF5/E15/HJ2yoJNTZ/jYW6GICPEkzpV7Qt0V+W0WdBfcKnjcpK/fNEN2N7+hVjNCYn4g
JLQz3FsVBExdtKusA7tY9Zbdhu/Pxo1eKolqbeDFUBtnG5fX6OH9GCFtkPXf6Fi4VFLb/it/n09n
2APJSrhDsm5x169XhXAWjl6hxMdFp5jhLKxdVD9Br4WPyNkPNyvCaPb+YuDKXK+mAPJholOifxSg
o/D27sRSHEtNIDXuZfzYk1Ug3qYsCtztkEIzPmNuhcuao1IYyaHrNTUo2Upami9Qsj2F0nwbjqZd
s9YF8Wpyjf2+6moBTeJb3++l/LH6pknpHwZ3I45OAKcPXKLCGOTnUTYBtTzX2keFe9IHv1EXvJgM
4LGWHQ0Wzy3d1pRi329oboDwZrvEBZlFeXeIbprG8REem4jiSD1TicvbU2oGkzbE/heSV6Pp3iJG
11I2WidDFn/kEAxu1CpaFHZJ3dLMytl4EZfIVXqIKUzB5TzYdNDTsJR1hjl5uMH4mJByhngsmKJQ
9Jq9tRkeDnqIVcmJLDiNSgODOXEHm3X0ilJhbvd2XFa5Q14g1JsIvOGsbvN3S9MGwq8sPjwU/yS3
S9oTTPsAi+ARN9YAJGuIbOwBIBtVk5I8ZV75ntiiXNopz+0fPg5w7HkNgwY72xQ2yZWuTSs/9F44
JmvUHzmZW7xrTPwlGlLVA2MGlgOpkAPpJLPD24vgyFswAx5YhkfxsTfunTWofVLO8n8VKr74ZeQd
YwI2AQWFkxiD94FQiFtvp+e/e6ekRR6YKGVUq/dtOTmlpdnXo0tEF1cFWqM6Elh6MPAneb0VjGuj
meKharDMxzI07cjlsPRQlIK0RMlYIaK+t5xj33qQm8rgvZvEWS4cpdisaDg/g3NQVslLqdg/r2N2
dgSaxR0VWRbnXkdALgZvUjp6iE3knlzm9kXIO2jZNIBT0Hj8CgUO7sPpMFPBjjsgrDn+myKqbjW+
v7WFApKC8m1ZmD2zRHs8y5QPm6qru6XEXJzPRM5Nq7+Djwr0+jxgPyqrcT8yOjPt4d27hulmOHCi
UuxsQEWtWPS8VkJKeEXInGn4UCt1tILnLB76o0iQ4jh2b4HpQuJgTK8he1ux+7nhqFlNsVFsvpPm
B81jDjfdv4W95njv7NqOL3jgOoYAkVtDcXDYzclllsVqU63QXJazzAmmKmxx8n15KEdWLV6himR5
HoY7qZoiNk72h7NDO9D/Q163QIl7+VVHVmQuQU5aXwZSq+VoPjb0fV34yiW6/U2QBc8DpOyt8v9V
PsIO7NOSpddCVrFSIBXyPMhwW/Klo6/KnwZsgnosJZWvOGAM1bu7qSSM+eYSkNB4SuncSD8K7BJa
TDHImf15je+rbQlvw6+iRRoQTjSDvwBnMU2mXhoXhEPQCXOtDTXKYiqjjOf05yMWave+BeVqlGHv
Ijut4Wu5JjtnNCZHT1hnyEUIvq79rKQUm459dAwqs+ZAlL/dp9V11vGIk804jukLO5ElbPJqrc2x
0Z2vx8XPfqBlkjjjPmUEB3rUra/d7DUuUH28nh9oNeUO+RG3gDUVY+behk9dN4XJ4dQ9c5Q52y8B
kI16pBHoiEn2hbdm3xlwoAkt3Z60GxXUgzXKOiCf0MYZx9pmu3KlM9HleDGd2yi9Oo735ATUAUEW
+o25ypk9GlzUvteKJw4MmM8V6aJcVIH424k9Y9x7nuwAahTN9WEBU/egLBlAlGuH1GV+qa6uPtuA
vMweoH9qGJMXU/KJrOengnuCBCU3qUOKc6rTfMIVFV97X1U9WTZixyLgDxvKfMbs7SPXIRa9lBmI
Wbb5KW5v5UpKOt3pWNf2oXwiRUeCa8BpemTsZ6w5VK8o0ak9Msjiw68vZFmjf9GdDRsyb7Ju9M8i
Nsyho1W9P1oQ7pecc4LSinuiVnNMMcVGLyfaXiqBNRCsyOh9MqhzcOKFtSHNI/+v50OV5wrAKUfH
cRVh3F+DWo2pFC3EYo2tSbRbKJ3603KkC8x2Vns+Knp42bp/Jdvs897FXtFwgMYdV7QYILpZFcm9
n3eVynUujr/1HZL2adCtOZgYVA20It0yQm6v4RxR+a0oGfTW0ZmxIc/9J2s23ISPa3FzYCATdLRm
0Xf2MV403uXEYASZ+1nn5fzfo4wDeMsX2Q5eNshXXB/RVCihgpCtVyA79Jplk81EqA/CSATEf9Yv
jPKf3dZ/i8cCUdAq9uOjcftSmKAPe8Qoj07VxnWfTDEempdSxA+fg0rf9QFqhCzF+h+1/U8KhWmA
t8JbS8i7g9LVJTUYrdKWeNvwkUJCHGBzqqoRhaQ2hSbvESHqi4ZAyzBS0G52WZfFb4ozhTVGZDVU
PhsWpkzpeIoGf8IjCiXhAZ6FWEJHzF9TOlsLOTKFS4M5QzaHXHQu19AaWDOqBvgaAZPXvqLGkD4K
MLSlcbuEYEOtMH/+1k4LVAeSnECaqynUTb5+UVBBfHe9S1O6xRqdtv82KOCE3Os9UxS8O/ptioyp
Bd/RzXuOidAaqsp2vcc2Tc9B7F0FelK+foCOxpRqwyOBwQhZ5Y4iOxMC6NMfRiOY1xO9Eely1q6Z
VhPQisij98sZK2QwjHfSv9ckobd/NJnBs9nKlLSwOGSnnqNPVMqrZi5ks95nZ0JHnYQUA2tjm7Dm
4Mkb4+OOCgHaopp1a+ojA91PAbvCcyDpQIuCFe8OXstynDaDE7OmAvJzY2Z42M0cAkSvhoc4CqM2
m9lXrA53UjwRb00HJdGeKIInTlLRUYDPZCkK225w450cQ2WxIlfR7+6QeOIYVH48CK5ONu50FCz/
zeZsolLVDDl/Jr8qye/Sjg+eCd886ctcd9ZtnHRgLvpHrlnT3yoZheqO1B+au6X9KWGpiw8doHI9
+JC7ZC+7o3KJecy9dW/OZtqdJst47f/tbf2UK6u7oG/MhLRe9hy/bIvEyTKrM9jhLE3NgZ7RDGr9
Phu06TQK+8fpyKTji4GSsHKL6i5nhjZZViKtrEjhSmofmHewGyezAZ2xIQ8Rqf92CRWcbKp3QXCK
xJMAcPrQfaaICEIGNUur15EeOeO3kX2eJPhKwgcPxNSfIehTrri/QVC6hP+3VR93+Cu5Tfp9CURI
S47qrHYzmYKUgwb2givMZpSt9OzKn6OW3DpLFh4stiEhh/RFRxb4VAZDf4E+UZSwFrLrOH4o+the
Io7Ya1+uRofD5YOj5CBokcGmcznJSjwbOYK4Ijai2FvL6ayLqg9oMDYQXtd6J0bdTl43/kHpMGrT
J9rJfBfYwCcr7ZAARJGn0BNpssh+xP3u8JFmZaZ/prjcm9WZMgDA5USdyPA+67zzQylW06W/SLLB
IQyVlVYw5X0lnzDVyvQV/uVQl2o0J4Fq0vO1zVbaidptFqpMImYVEkM46DYvisEv9FTWZfIw8mVZ
UkuExjLHDXxmxAGe3xbmNLd8HQVyuKEkRqGONWKzNC/59g5ThWO86M27T9917eTXe+ANuGM1EtH2
vZjIx3GX9PZV7emqSvB0BVG9JBIuubC8UItj6smQ2Rk8ubGtuUukUZbkKGlNAgjsqWxOXGzeRTEY
ojVaSwPnyjHf4AxtWfKaCvtt/toLJXxjIdZHmBltSYKmlPa879t5nthRcr4w0ygHwwrPfux6xZdL
s10qEcvVnMX7Lx+ajaBJtM0htw+8ytrYZ/JzyB3Lh21T/bvNCged7RJm6qLsnzeYzck2kiM+p4i+
5LIPCcDgjhOapcuHWbXFS4Lj7rskVYdHiXT2FpXTyyGgg4efcaOfRB66klAEzKbkNrCQHGniJZwY
1wAesYrIy9OykL5LY5YbWNS2bU9BcF2Mp2QHBu0NCOjeUwrhkd590ozTC6PA5KPWrtLviFBayUAQ
dJ/1CAONAMv6TtyzNJuWngLVGhXvGhydwyWV9BTm/BUMg++KDWiay5FFCIU6e/fblhcTd5qO9QrI
cZ/eWdgYZjYPN1POL+hKewfTqpdbJxWZHtdxiZkfFJrJ2EA0xwhGbT4uByC6ChUrnuRNLMRZo33X
kQJ3KpqJT73uT78PUbsvj2Yj4pxht37DQ/I5Liah+7hXp3KVgc9EgogZQIlQC5qqJWLGs01gzU6d
E6rc/40g9sVTRYOc/+e+Fs1PGxJXSk00IjHKzawMK1Tlp6kKPwlyFx+BNa+ouUxdg+dIl3Jauqhn
GuaMZ8KHTKiniDz4P8UIA1QMYk7fiRkhqv1y+Qyzjv86x5n+qbdFlWPpq1D6g03LmGEMta4j890S
we4qQi3qMObEiQTaRISslzPFEjxc/s8S3VM9HnHyXBLRQZV5JrAucXUYL5a94dzw8w1QePCCyAAt
ZpBdm79GE/3Xz0ocQ1ew+jykFG6dCxaKwvfzcG71mKgrH4RAb6qXE64KzGK/bEApjwdQBxHdb+kH
bmZk+prwqvaTpVckLI7wEWz3mdi9fKbGIWxTor+lz5N2/FRMlQ0sZ/w9RHrmG648Tmwfd7HCoLcz
ybNQlb+7iwOIx4VeLL43q+dFklSEw+EIy2nc5zlrIzAxeLnLm21Jz7P3WRPbpbPCqSUh1p3FvgB1
0d2/0JuocoUqxiiXkkXiztmW5LFggSzFecCTwPO5AZiUiNA1/vj7f5InbTsq9ZwqGJfk7nbb+wFk
C3+2UYrN/QDKjA3ZgFK6QHqC6AMLWPFh9EIBpn6wsKXQItbDieelKOARQK7t1pVS/A5hkudycbJ+
0WeuxMtxzts4YzDZea5p9WF4DQYxgOhtYWpqm3TL+sjcpImyw98vpsHc5I9JSzxafR91WO3/ef3z
/NYhbfq3E1I7pUf10QbumnuxKJLOFvg+X76rqc/e14BUYjzYIxt8m8FabjXB3LzTQJAt3IjKY4fH
33/5bEFWJlizNSrBOqZWB3g+crPEktuis0LokI/g0TB2/kZ+d7VffDh/Aad/x4jm5JtDDm38Oq1/
9UhspO2T3ZrOv7txFVMmgM4mqEEOi2q6Qd/cKVYreQYb9LHSVxh0yxc6W+TnSE5/ESyU7ug69hCX
z49L1UpHFRThwb7oO1k7MjcY13Z0i+uNc3wwuQ4/UlwjCExUJHGb3x/ipTzOEWkjv56sT5BqH1cz
v1h4rgif/4RK7M1+faY92OBtGQCpVn9RDUSKNI+IJDLSwX5iLjR8H4+JEIXOM8DanGYJZTWL+3Ol
i7DEecYi+/jooHQKSgfqjJArbQLLvW3k74lNiSvZHV9Nfz+5Dmc0rw2mFAB0b+3vOvZ1y5SdfZ4Z
cnYBmGYKWRqwQd3C/jnBPw0IZ8cvTem81Ia18t1jkw7OMkEVY/r5X8e5O3tR/rAmB+hl9dUYaYZl
a3Y0BEJ4tJvunMe9GM/F/j9c2PiO6aVIA7SFzByqDKUuiw/y4PKzYbr00ww7eXryScLLqbBRX2AB
TT4nJABfmeGtJAv/XMIytXtiQRsMahZl3puDvOfk5q8E7TUwgZeLwBrm+GciBwBmAX5UobqD8qae
zarGzpy9Z24TuN/R7v1G9s4oJBNKaGh37HBQQXaR8o9FGUEZ+QgQIdkPaGIlQxN/srwWqu7hyJqD
jVtNQLOWBCi99qiEHFPVWXwvqRJluvM8DHL/f9NVskJjr5dEDNUFM81kiQB3Dsmhqib/F/PyJWOW
B3TWJaDcfUC7UfABAwfxwkjhvCj1xMFGL2aU+VFBNRGhNz8XBJRmqR8rRu+cl3144jBwS/NCU6mS
08UG3w8oG0sOJVkW2fnVULh6BRgHPcQmmiRdXOORbQjpg4nN89SdfAZE7/7YoFrzh9V/Q6PoBrVx
09xLs7A3QHxqPba1FDVJqys/nA9k4mb1sVvNbvNIBgraB4Q7j6mpxM6K7wMfIRARmMUkz3q2Uy3p
CQKYXR0wyKEgUwgx9FQbokAlPhkQMt3LVJo1B/8GAdz7bqgjfyu22dasoHvmOwHCgMKzdTLvOagP
HHe5U/AdSe05nVsYqsWm3NqZ51PhgnSy86lehAEh0G5gOlfpnhExEVh8cyxkHVyNsprduC2AymEf
P8GR5oHiN4D8ggPvpcilrJxBpNcF6+mauj8RjYKOAqk3QXJPIS+hTP8VfKosH+kWkegbH8RJBoff
VgAi8XA3SfdZIeNfHjrxn4UWmCGIDPjuo0WQakYOW1u5v4mja+tpqXJbBL9obzRrQ2KiZUSxxCqs
fE8eIrpZEh3lj/QniD7lCuR/PYFlWKCW5NxWw24nN8lTnPO8ZxHTVNtkOBQlY//OzWUdCqpHHoKk
jts2iWadgbjg5PSdAFwOt1y7yg14QtgMkAcjVUsCTc/WqQ6Y6gc9qKwaLNjY/OVuTQ5npYTKoHCQ
IYVdtEuZqMnp1+j3gLBFcqLaJc7Ax5Kz0ozhfpxCuhkunnmnn6ERRs/W8RSE1lx9OtWP/FJfyOCf
YiD2NOKP6e8KHhKPSjjAH8+UKTyB9VUgaoPmx6G/vE0JWuZBUtCnzTk16dbtq8spNCyQ2Jy0OkQh
mkl1krZDSCvR8dgq5k2oQmFvr7cYfj+9YhlNlP0k/hCgReo86vtMpbbPgVDExzi7Q8Y16sTdw6Rp
Jj4WDzq9iJmIAkAFFahcEaCRXCD3uCENQcdNnbOvfIHL77EW0nnXxwM5EdorsNMYbPszBvzrfwNI
lwcAigtEJrOktI3+KAGIoYgHq7rpI48so44Dd6kHsYWb+4gZTYq/WvvO9BT2TFbEroH0TLqdvr9S
0DG4RMarskNKEW6OMnOakxWWIkaVLuNDOqSv5XWjMcTnA73CVbv6xvIYuXeSqjcr264eb21GIYSt
JoLUe6b4+UCq2Fe9FLkRiDDPWNKT8UCGQbe0nJddONaId2mPRhrykagBU5K0OZdz7oVGH961M4gR
GP7QsO25539vu9jRQc+ZeaVgn6qO99tv46APHjN9StZ9zftARl+EQPoKAM5NWN701Wp2UwjZQ9Sq
zVSDHpF0SKQfcJebeXMhZusuYcdi4jh2Grfiw8ls/97kvPvDsfFmx8vfWRRrChukXdVHOTGjvzGQ
S1TrVUFpMaWteQqbFj+sRM6bdvEK+++7SyVAwBS8OoDV988oUfs7SUp9JJxtvVDevRzYUj6Z2+K4
ehPOoUkMXZQICmQiic15RMFb3oV7HD77ME6D250uosdP56ntdoRh2CeD99DS7XRkHC0gV9JZZwYM
OLJOXbqd5wd21yn4+YYyIw5AEKQH8cc9eBO1SK0jA29KIyoGu/pCjGaI7eknuRMPikBFlmOT89Q0
jGTgUedpJBQDCiEfzduIz+RvHbVYXPRg//kwg8hFAKiTEDJdMnoGi/0nZ5xEo2in/uqMDu9/TOHz
Bn6WaUxETJRyRMI8MONcPrC3H5PY9QRASW7rGVTRzj0DAdbpzQhsAp/AaRGlDmvh9BeIcfqiK5py
J2X0IDX9LNfDJ5cvEoKpUdXBMAMsn7qIEisCMqmJ+kvoWY6tWROZmPgn52LHClowTuK9zi4OmFnX
XwNG2V4queCFxlT5MgLGjvtUmdC5RkEWBtmcmdiijdDNa7dWVvBQvhbkW9F8YNwHARVJ41D2bauY
GgqCxyyh4h1mcTqB/mfv8Pa0kdDZuPCE0aVxs0rhS6uBx4wWx9iXulUeiWJD3cq7YpbEmH9GS8fN
5wfo5syd9i0e8G2ZPl9AQfQ1YKSB5f/Q3l3FpORt7t28KpoAIznwsCmRsoKc/aLGw6ExIB0okR7n
SG6ccNkOg4ESpSqlBzSLTm85OSBps+LRvs9uqyzT1arvQ4XzWFNfz6gkmOVIRWOvsX5G+O4roPlu
tZEKLCACMP1MsakY9dN0/HC+PNYinqzPCMTBTOUCeGFxwhfBtqd7ivjILz73uoMP4UeQ0jqA75dL
bKEDnC1RcLIzG2gLb+n8TruufUL5Hzc+wyDV+FlcBBSp8EYZ4eoVr+UOxMY73bAXZfSwbyHclpcW
JQFsybiGMsdstpezQKP5TbAojBW7kd4M4ZipXsoRBB3I14xypjf4se2agustnRAYoUE5Zd9+HZV8
hUVrURrFxItTXk4eIeOPFjoz0AF92TzYL7h6MDwamnaU23mmq+47QmdLr5U9LxeYvh/y/+yXa06v
1xy5DEzSm0drr/WDQl3Cz03OMySwc7por3nFjnXM3ziXHj3MPf3OTj3cak3PzCHC7OYBMqEEHdX8
URMhuzEEYz54lWfKRAfyeY7ULIjawq7deeR3q8Gzbq16djxPwygvbkzaJ9aWWtXHNcxw0GvzspZs
GNXZTKMt6whYIzeDT19+RYuRu2JR2/qVQMjzNRrrKjimpKO8BFQSgozwP1XzLwym5avEK5m0iaR0
H35vQ/ZGtnAtsY58l1IE93AYqTaPTLcmqUL7mvCWmE+cFEXlPqazNAWV81BygloTg2uEZ9dRWmPD
UPRUCnYQOgilPph1ucIxv/Lh5DsnSGK4MqMsezES3WMBNXHRVvHRC9lNW1YM5CwkasQzpEbV9Szp
LyQ1s92d7h74Nqd6Rk4M0FS2uw8gX/yIOGfjQK2I4/87qrnpPaZOvj9XXfbFUflL2izWZb3R7lW9
rUm7mLQyoOeRNSLDqczRM69yKo9MSvUEhgG55JaBMWCMoVq8Dv9zuX+xksd99kiQeJV6N04f7AB8
uxn4qQz7+9TucEjyq50Rd7y/JlLi3j+klJ3EnfxJi1aBrqXBIjs6FclpqhPNdx3EO2fC/avi79Sk
OODVh+/vWRROPvP1X5NtnOrkgaq/E4jC9ZF+TFrS6Dzc3+VNils+f3sEqfMiSwktrpRRNuo4bECu
aFVEcmFGO8Fv40HpI0DIot4tSzEpUXw2o5HyAEcFXKSOp+Tym22f59JrUk5FNDJYfZ71GGr0nlBb
jsod0XewS0j6yoHn66iiiTctecG0V1Ebnl2oQP87cba7ANLANJp2l8djEjVmGkVqgif+We6wjAcf
uSL1a9odYeDWBsP73+vk5CYqiTK9yFXASeKb//CO4RGnZURg888ol/+qQicH8i5JJ8G4+QInNJa1
aa1a7CzeDcpUXkWdkaWXK4D3OuYRW4bQzSFuOu6sGxMU7smzNGUkBo2FHo/vmyFx2xADas6MaFa7
npcVUmCHTuq1YSQBeyWrpdw7swzrQPTOV8CajdtT5LKzGcKKzWT+QFxeE2npl2BYTlRFAmznFQaq
q7PNDUUFY89NzGlyHSyuYOlFMkBqXOsDKm5wB3o8vnHYevqjQz2I8WimZYLdFSzEgw3I4zFFDPAD
7qn6IsZ8cpeSWzKrbPXi6+ROStGMmul8fwiqaZcYaINkXo3F5+12CYyACJQ6zZNWYXf1pYP6ZJUP
s5gQdwLS7x10hYPxVJltO89AlU/3vJ+6RG+QszyHRZvuPEOupaKzntU7KCoTPYcXTIUAHNX2Sy+c
yZd+jy5kn+6Luew/z4jrfTSwwefTlrqavk9rVSyrNx4w6xJnWPjTA7IK9wEvStJys7bVZ26e08R8
YppObMRZclVJ+5Jax/R1uQD6gNhmLTR/GSuVL5bq0rLIiOO8ElvcT8ue37L7FXNpewQjP+YTEVsj
Yaj/jm3U0+kPWnYSHV0saNaQMJu0AzPMZFDnnOzMNE/C3s7pDXOBe7QwgtsZb6HAt0Tf8+kznT3I
5j7NY4JgOquIi5acqe1crXUgwh3bigvFFXEmImnHsnFJzBWgPuzksyiWwktivoIwk+HRz+5IJP/6
JJumWyqNl6zwjs28N8e10fvuwnkgTRT+wkb5PG6pYjcqQPGL2Pu/jk9ZuiU1AI/AjAptxXO+/S6b
eVLQvm3f3CQvjAkXJ7IR9siCCEKMV6AsNHbzlsnjQmvzLKqArDqgO0U9fO3BN55cFjD3EcdDm4tT
mIsyMyaLpmBp+/AYM1+eRez3xLPpyXJkA50cjCm1p+CfxCuu0chy6PuMvStgzBJVLsTikBIeNLWC
WDTN/SxbacRCL6MCanEfA+eIdgK+X2A1dLf8Tgk42pOzzl0q9wxsJTxVI+uwARySjeE3Fs1pm4ug
KsKt1XY7nhBLlNB13jCXLLhQOR9EF5LrNUoxTi1C44iDG9N5aJSdcN8F/q3ykftQ4pBH9pvJPXwt
BG8j3+caOtrqsc4d9davVKCFRXtzq3Rj83ESVUsGkUAKjDWEOnDciZDdsV3lIMlkEXz8W7FnMP09
fg+mRXGHFGvYNs1Jzo6zGmvDvFvnQgF4YgXoKl0Oqm/PNBgiw3fqZxEN+Z+EVFEj2XMRXYaAnmVi
+7QvsQ79wDvsafHUHMQOUo+4ymWwlz9QTMJlA13XR7Z6pfbgJFPmZH2UhbmNuolDJcSHiV4BcwSL
Yhc29o+RoBwzmansbz4l7ygFdN9uoGFnCAt2PmGWlb5jA8Ljs9rECiyarkE9Wqv6Wub42VKqbsLY
O2BqWpDcREBRE4JqbbahFC+FgpHLfEv/99xJaEnxbIfGSUHdGLwH1WsNs1E5X2UYogsaC6/31QbV
ra2qzG8wqSfe27tnoNh2K0MD+aYsO7itwf6FZmVv4e3mb05pYSpGF8WPN/UL2fDsNb3YrEdusUeY
w68hUR7K2Bif8P/NDvUPLhZ+5kBx5uOnI76BkzV66s50LTkAyEFFenaezR6XYVO2+RU+3DefNx3j
dZIyPgwwNDZjQiiCUjFP5fOs67amBpA4Asgtw8TRqg05LCewgbqmcD0HM2u1wvWiX4HuwD0saQhQ
ZDtLNwHtg863VqkhQ1nlRgpsz80VdRWoRuVd+7uuQDUD+swy7q2oFVqJa2CGqVfsPyDqDVHEP1qu
mPsPT9epzUX51pSD+yYYjVRjXx+0dL6M8Q5HUzSYow15JSKbWWNguD86CIHwBxQnpX4HNZWubRFa
+Rvrrse8Kz1z27K9btkwEpxbPZeVwWIN/hN7DWekgAtb9+/tSrk8DyR21Mke49+7qrxwhAeaiLXK
3AZtz59+5rm6gG5kk560KNSOOtoPo5hs2KrU/NryN6UUrC56L73TAckN5nl/GFvzvcLsHWbuqg4V
vctuSi7EcOAX/APLG69oIjLlbtj75POVWDODgkbaPtCKysPGMcW2SrKd0UPR0PGBLevEOuMmx8c+
sZr7BHOUfLKI3wDUI2MMkcHgpfTRQmk0QaawJ7J/iqimWaZ/eEN0sfx1731wAaQu1nf1ZmiR171P
dDE1QxORYDypoSwwuw/51QuFW2xMze2do9ngA5Ys554ef8ZAhoJg/M2yDDXn/Zo41mRSZKqMlkK/
JryVV2MoUTTX7AOb0aXMoUrZfloftL0Le5zebYJcMCuRuDOxcoiBu1uIDi1hraW/cfKfXaV/L/F/
rDbtREBsN3rsbZAmjTw6SEH1hOGvsyB8yvq9BFb9O3UtQVjarCKv33hMDQm3U+n0Floj2mIDFQiy
bAc93x5/4dfgN51tKUk6L3wVYRuYteXKEJRj0zjzLk3UDKMRvUSsEmRxR0g4xfgBh0Slh09Ix+l6
FDGFIG+tAOHjAP4oOdvN2QEcjyxRVJh0u2FpBItCqbJQvRGReAZ4/Wordjqo029as/euDk3oh+/6
2ylkJuujQeCixHica8bjwCHh9BdPzcFgZhnKxq2XPm+yKDeNCZDr4FEqJJ/+kA9s/iVTowArju5P
J/uBzukawTWve+ScmQ0LfDVWjuDdLTpE4bwB1eULK62Kd9w+ARgntgiZNmDOuzvZA8oHAYbbabFr
Quz7JWWX/WxrOsQo0IVj1XS5AdvrjNfn0974HW0/pUexIWoeqqSgjRflA5vgsBQ2hWPbCi1tsFH2
/tYHBE1srTsrc9tIgh8+ccdX45Nq5ffSuifwoprvpXHJSj4nQD8F5VCd1siVZQTL4pDK74oyyGVq
EE2Fg/LLb6CNUJ1P9Oz8phvI44ajXBcN9JwJ0Ft/Ik7JzLsTm/TpstsVVXZg4EHVbH+oHI18KCMH
3hvxQE6KDNYHUG/IjdqmYjyULom2xkAETC2vtirbysnlKFIs7xIQbyKZe3Hl1D0385ANRWWtz3rk
5CMVbQ9wg2EcGVQHUO+zYMfCilMS40hBBv08eryWtMVifO+O+5CbaSVZmbykml8uKDBFMzIBCWvV
8AdILLiGRpzkAZ1UsgkkfY981Xh8v3uTpiIaQUlqMZ6DggnJbZPl8vWHFzdJW8cNr1hKSASHy87P
WkJN7zQclg7S0FkHP7O//k84qE6U6o/SZ022wNGewOy4YQ5g6tqWSXUZFkxsYdfEgIm4UD18YQPI
qAS/9sEOlP71quzqxq4NAQSFVjQ6yFP3xASAaVLsNNrpUDZCSAo55X99fFTKw+8Fk/8J+OAjBOxM
a25lUZ80RC96yYd8GSeGTnpRqAh6znyMCBX8QKZGWeNat5Lp9ybtGHrZmtm3MlGg7G5avk6rwERZ
8RxChUCvEwKyy0zZNkKwJpJ2AfAVjqF6gDA78Cx5pMi1RJJA+M0avA3wzuIRpaWlbBK8we7LedGc
4vgHZWkqY1Ump1LiamkYJTPu0aOBsVmmso6yt150CE+FsmTA+jm20pIrwC8QGRq6nrhYzJEz6EQW
TxB2+gqnjiS080WlxcFboc6e4eJIw/0gp9UIULGPNsiaqhsNbDB8fWYgzHy8HP7bjvomEuSFRfzS
4RCKZz6L5Ms99MJpvb2iqa5Tv6Re4fx57yvXIWSOyLkGSi+2KtQqRw0Mqy/iW13lZIuzfK/8ErnW
TXCnqQFjT/ioWs8AQmvYmX4GnSIpVFccA/4DJYpO2XgJatfX7ZDNqclmnKFyBP0Gvytl2nHW1uES
v0Q2PAxFj35VPNi9s+BnTCdcF0lQbVnvzcVXbzgyYsErQFinRTVrkbh1UUE6ULubALYCQc2sQP5v
kpqcQFfBv8tFJ9HjRz72aYyyKsQUDuHq+wp8RdUvsUWNR1H3/5uiAL9sJWkeDr5btxuUfGZMcusv
WxsnxKxDYvxdkXCoMNYxGuRQbpNBNJiH/pI9j5W8B/bE1z14cXlOAiGZJ0N4slAfiPTtHYRRDNyf
mIVUWhEneW0SqAiaw69SrTSOLVTJulKsusxE6KhVOGzwg2Pwi3gtLl0MIErrN4MY9pLkwF4QaMH1
KHS9LYOjESrb4hqZUQhVMqj5rLmn0lGUmuk2CIkiSJvluYex/ySmWN6/xhPFfliAesHzpo99PdNF
SZ9oJlpLoQnnYcpB0p6Uzd4/OASFlFL/Asqi9H/xnB3kpY2nVofpO6zUYSO9Qb7FSPojEn61+hk3
ytKpeyN+PoDRgyGqdEb1dSm5OZApxLfuRW34KInlaKBUCIVDYeVLup33+pKNSOno/gW9q7dTWpEa
YOCVmo3eBlGouFDUQ8iEjEgGRYV741rOyX06lCGyA0FS5odQJkvs5bBDoxyjFtHD/ckgfofy2b3i
lGxVc6XPZdQNCnduAyAlknO9nHYDV2KzptvAAOaUvK04qQoKuWKwylN7eHpXwyPVUK2/0xm631hf
2qXHtscN7vYpN7mdek9ZBLuJ4LwC72wIEtbdOX2F5iwDjqUeVRFGjPX3OlLqlx/T0ULmV0XSHpMd
YKf74US2pQo4VDSxKogqLCYDvk7zch//gQm6pQUj+yC8lKYcVCHgNRSatz60A+tdpx/iNs+aoJC5
uoujLtKxF4ZWs4T3R73gVMkgVU4ah1PA6lMmN3ecl+PGDnOybM39BndaXmxkevIVtyp5CUOqHnO9
WsOoV3kD/pxqXXpQZu6eGhTLUIvIEZmSB7BrP0+SF/xH0B9O6VN4HkwwHiyPFeHYnhdPtn7c8mhT
95JVXDJlYhr/dH49hQ52KUmnsDsmq5pvBXrIy55WR++MHdT2QuI1Itq4MWXjZGRMWHMee5d8RyL1
zEl2rV/7nvaMRGGir9YOVvxqp5Ib0JbXrgeUSNGzk3SyW7+8GMTcKjZqrDPodC5nbMk0AePTfHi/
7An9LmqCPG7rQ2yHBjirQv5GJ903kJ/tNwQFOW6D2xJFmTChTHSooYKGEam8zmlb1DzhC8j1B4Mm
V/F85US5Q3TyclplUW+EKg8dUfdGrWS8DpHFR8ZF6/fYbj/BbvI/Co8GdKShdnR1Cw3bjjzhxWUz
9io4RJP3kT3VbcgKHUoTPKS1bMYT5corLjc/HKCaKnrTzT0Uz5wyTGdcw2b0VbKG8Ov0kP3LxCh0
KnMR5mxaLbH5hPzljCHTpg9jYzhf6yZvmu5xfSvhQr7DU/AdT80TVbJUk5bW7N3ARbl+EpRHZgwQ
P6HpAfEXD60ZEayOX5dS+3GZrms/hoMgExskdnDRxCcXCEUMsQw2cKiPohCQw4FrXxfO19f10Alr
O+v9NW7K0zQubcdEIBFzjj9Uwl0H91GqkzFqYWdf0mA8+ay4QT8qvh1LtR1OtxmMvOR3Wz+5Xcbd
Ut7K7tHKO49QlDRnCYd2YR86g3bDc1efIV08HcmLqt01ABV51QAuMvBZez5cYy4XrKMYBZQg3/RJ
0ZP9aUw2a4svZ38Ne2MC+4PZlpCv5WKT5vELksqseu9kxztxz5o+2ZcPb7kqkoXD84s0UI8fYGLr
WEsGM6dV7V2jguqA3/Yl1Sbmmj5aMjybsfGsJIyg+vxszi45qM9Y+xVUg/72cOmIDjb4CMV4JMF2
SX01xp+PwEdd9m026m4CdvgqaXI3QNzpQXvd+HHFO+zF+vqVq+skeP2y3oqugvLzBy0ykXwOW6zw
BfjjMef9SQw68zTKDJE+CqlbMRyMH1zEX3PP1rPaL3dKygEy6N6vuvQdpy1Re4AacdMIbO300ptY
3cCpEwfXv4pV5TzwQUVGuhzcRr8tG4PXtIukzPti0bhLk0V6B//mafrsHuKko9v+dIgEmeZPTIAQ
k26KQvaiNTwrNnaJPn9UtTSVkAdHJBtkB6ilodhGeLOZq+Y/V/kd1i9VmOrz5kNrsgvv7QEW1N2X
yXDm5HBGYdeAK9VI7e/NfLfS4r5YwFwENYASYpwNve4UsBod0nx1PNpp6H7NKGGK4N1HGlhS3pHK
RqyRpE8Sj5GoCWTMeDcJVtVIQnRp0JgVEIZ92TJKhR4kmshl4uSkAdX1JYp1gsq4nqnAyQpiasfM
47z1JvGPTKXidk4jHA9MjqoKU88X8vVv8PHStHkyx4pqUPebG2OtnbtuH8ifTPcmLGY82w4Bsfng
cWgV1NwyMq5EMYeARpGBxPFSOMxv6UcemPG6GFNYp+qjEE+yZmrO24TnE5bx81yOBU56x9JSKKJZ
1NO/ef1kf2z8ZccYHEcEO7sO60Cp1LY7QLwI0WmvFWn+jqCQ+jT6YrGzNcEZj6kIrGV9oJ/79NU/
9NBN1OhJ1ZutLSBjwf6DeE4wSkuYbujZBqtdAs16TLxQqtCjytYvajAXWEPXn6iCO4leVlH5w948
10KINFbK+Pl3NhhKZSphJl5N6ZsrQ1oAW8scK9BnUEwIgF3I7JUroCWBwEWlfxWl0C+vgO1pHNSG
CmXAffEfs2T/xRAJPGeA5qPljN0ZBPXzPl9t9slnOt3sxNgJlseXlJ6kjAJL6W0ydG23J0C6lUTt
0HwV4Y78qE9IpUQ0N0ZjOKleJl0BwqHXTAtL0RdNTklAgCA5lSeERh4+lryh3O99I6wM2kgkx0sC
nv/y2cCzW611XEJJK+DUwZDK/caRp2PGcMCEiHivc7cmP4i3KIt0zBbO9+5JGqTh4vzOLB9xtt91
UfpbdqV/nVVOymgCVg4rfQBb0t7URuWekJW+CWQbpXDS38PVBiqeq/t1CSgFvY6HVmzlASHZnjFR
OiBpWlS+SIkO/np4uFm6U8R4wddnk8vAC2r0C6Cb4Lk0LJRXnv8jfPFdHaZb+PSaxeqRWZCxkVNj
iWvo+55+aktH8Bm2/GxKvmoh7Wgq33DI7BfY6njJTa2P2MHGd9pG7itivKW9iqu9Uc2V1a01JMZd
qEkiNV9o8XsVfNQJNXGBQJOS7erWyOeJxXEP2xdkA7sY9M2RCFZDUD1msJZqfoTxqr8MGx+GmtQr
pGacEUDfO3VUnESYHMb30pr5/Jt6sRAq8eQ/4j3NSQHKyUw/krA251M1Kwau7yM2MSUP24+Jnuoh
BZXtH2BeQBCnuC7J064EkTyV11FM3PKxlWSY4KgXufxt3apj2TAq13mKVBTw7GJNLFjclB/nMaXL
58CWPsbtBn2TAI6F3vNOcerDKH4Hdu+dq5l/Yv8BV/Gwg91NDD4DO2pFf9PGUwP8uqsh/kXalYBj
bUwmJbJs+B+7hcsZvySP3fQRNNyIJ0UDvUlR0/iZ795+ErNB2hwDh/dwQ34NwLpwjOoWalrm0g/l
0fc2ZVaz0m5bMeEqlVSeqYd8Ck6PyrJC8ntwuP2xM0N1rU7tM04x2H/29BoQhNutc4oj1G9FX7c8
0FqYvYMOx+5ZkCN9OjNmZDZRtKqlSYAeehZ4M0XDUp3aIKvVjieWgSWwa7wjlbMc/BAhSMILgfIo
tWzZsJo0twE7lHeqVaOa2qq8Wri5owfxF28S8O/B1hAsv87RNHYnM2j/sUBOcxXH7DXjO8A03yZo
HwCPyOCMyM278vLLCgBvAEkufYas0F0ZXFQpbHyzzaE0oJIl57RxmmaP7qoErrD3vpUqEWfWVFf5
Y/Nm+Tvu8G3PYIrvj2U4s2XsTVPivP59VtgllDpXEq1bL78a6cZeaK8nyrFoOe2NO84jUCwEmOEg
F7eVPUzXRZAiQjPDwt8W1Ss/ejyBgdalj58Ko2C4Kz+N2S7ZsJ0Gz3ho3inDeNjedbT/L19fq/kU
lRVZOwo2T5nMYqSCj0ripDUo6ggq/YIXL5SJ/pPe5k7EyHFHDSPIXQjkj0ALbGyDsd2BrdtZACtO
tev92w599HkJFh2cIgKlan9rFnSJZCV/R9++EPJUTn0rnlO/+JhUcTxZPizv0CkpC0HCAH1S+Pdp
5XmXTO829ABZ5CUrtS+oG/Efs6Lfk7lPId5LyI0nWVlM10olLIrLcnX/n5xgteU9wUYfBvEiT0gB
6b5sibn6vTvK0doFdzACDXkjIGRSCl326oRxawyXnOuLeFRlBr17KQrmTIwYPk7D8i9VSwewEBRL
TVjk5dClkRqoZF/aOLZNGHuXF7m/G/eUH81bM2tJqWEp2Wzb2VUToA9GGuzWeNCI+3zAXgUdyT1C
zuzZUlHS4vHfpWFo26dSl2ZU7tvF55eUGe/VojGT1goktsdWKQoCojT6+UTwLV2uaFkQ2kStQkwS
elLEV9PqWNAlpDBcW3eRy76BrUtcu6Q7lPDgE5FU1/XLGDJExafKPtJdmT2aIAsJrip7cprMGs5q
JXvrAboZFI+lTzBoFZoFQrAmmmzrHSeYRcPpcNR/xbOXV2CzgScZzJfk/70eRYyDY5aLnp7ukGpQ
kFZMvNIDcEfpwUsj8aebV2ygG35OzoTlvMjAr4vn1AnbV2CS14D6vhw2v3T2ksJaTMPQ2xvXwf5y
yU+tLqWS+CrXnKqObGMLcxhhGxPtuf/hFGULZIvJhxAi7TuXhF9ypoXOaE1a8ta6eUUpR13W+kO9
5WHE5KpSiC2jQdnT+YcA2WPwM/0wmVvjlZ+4vwdyEm0kd8RBRTsDDtljwrwbWYYuRcOrUdQHecKi
5FWGgMAwh6DkVCXbQQE80qAlLU6uXbia84aDqz2Y9ZkukdOUKrl/CppdEkKeAUGOQPcQ1gp6LvrU
iOTqeKQgQn48eTKQWhyyHX+htqp/HQcQXnjbMaQUjy86kU+U3s1fKFUld2FlO50RGxYlTOZde2Tw
ng52g0LuV655357VjGSlVBszkyGny/OA/Qu4zzDYvKqT623gY46xmQF3AqXLlLQXUDNkDzttuEG2
yZ8ew4PRuDjrE5gNq/0y1xmG7Kjx45JDwrJ8nS6+HtC0Hx8qhH6cGWcVwY3sQ4cBV2P/jUU/PGTM
z9BNHXFsFnsXKMDOMLpB/sy9wKcBdHqhXglaUTRx96aLhGpNCBJ6yovSWIxl0JY3bMvNdkRulu6M
k8rLnvNu7HFSwZw2GLfsXxbOm3mKEh4PtKpNQLhzbZeHp9xp2SZaSnvJsYfp6JvGL19uFmcwcxb8
JnXYFglvqqhcRx7CvpWzzGos8sREBUtbT112iepQvkkDFVCIoM+apSnhwbpDvtHwVqxFozeykrc2
o7+mgB0YVgi0zZwjkejxro+6Bo6PVaAocybtgxCW5kM+vXUII8aq1FlckilamP7ay577T39ekI+f
9Fo3oNLxzXjIRliD+zRXWeX4xH2bYglebo92IguEvhGBnVA94qOjPC+1nGfEQ7/Gi2X08FVri+IJ
Sj956qeAYBnKuDt7GrDogbQgd/PfZtQwA26kbuQR6JeQ/T3ZAVjAydK/nzU59FfxkkfRbsrHqJs1
WuUJwdkSHGkoVMR9LlduX+EQK9z5AhM3gnzQcRyb6+p3Vj1gA58V9Edt5JlR/7xpoCda6XX8HJxs
H1XBYmm8BIcfCenSMpPoKSMX3Culg7ulYej7+s6RLCnk83ck2buimRGXe+1aoyTnw6djbhNC6AWI
3mKaFMp7cKoD4t0VEJZ3xwr4+0FGOKWjyPbn69yB1nRUNCBSMYXUdN1bwET7shX0xjlreF0Vnk33
BK6rTp+26tGwSssm0azs0EYOkkWMuC8mym7G2qjSqaDTswzGUOnhOjNUQ7FlXrxW3tR6fmLaQ3k3
LQ/92+VkAp+5lSnaOfn/rYhsAK8iZpnQzMZ3EAP3fUCOsuMcxk/ysut1jq4YbOnksat9xDUtWuBX
7lWt9tVpljpF546DG4oCGyroyRRk7FUgJMwKVPm1uh0cx41pJrESiXQugfVL/ZlarbyVmAEiNHKI
83qdTZwXZLdW8us5SsPsdw7QtMPb+Hhv8eFyUYk6QKWpSgk1F3zAAVyRhAYzM+pBh6GjXhzk6jdI
EoD3s3IfMGnNXKgRC5n2HWJZS+fFJ6EN2Mo6juadQ5L2qeWSm2NsqeI9NBzmQgzSO+75/sB+aD5h
NZ5pdKl28VIP3ZFTJiFhG09dQibileX0oCzCDJZhY1QgolF2V9fzneEPbxZG3nTpYlCaoPaoJ/1O
ebmjf6vk86H7u9BC9fIJOYVjt2K1pDUHqeFxIyilS3FN2R/cinwMxn4HuHOn9+wJ0FKTdkRZhFOs
Nelzk1ZXenX2KbULlzqsfkHFdktw6qW/y17blSML1v1xXweuBjSzVQW2kN4391u1TkycthgtQznB
utYp9f/BsjLeTzF+fcnqTeF2w3AjpNYpo0mX4NVSnNJSPwqy4aOz1cdrfbmHxAP0BrdKgnmnUcXf
g1FxkhFY8gczRJ9DeUCp/h7/5//zlkCok3pYoaYCM77q7jY+rQ2S+z0MPc4JlOXSS7iJdvAJKSiH
GZMOYY7ol7Y0iRuRWKjVFapH1MOieOnlnWJ6o+awcJBQu3OXI8oOAEI8vOt+GMCuDdWmVu/kgPaU
z7dtrb7v1lPib6Y1VIJH6kna/0HsOT1bGkIHI1YrZHDJDZUOcMq1JHy/FLGmk8OttHR3Og2nVTS1
UBxR7PxQcWdOWuWQb/YpWLrXHqTOnWO9nGwJLefzW7HGEZ9m4zn4J3GfMOXxo9bLXc/leuvSCd2G
MSGl7lMo45kLye45PJIGGJieN4W8pWvs7U+PTQ7+k8N4sgzK2Rnf7ja6+PVf7rqvsA9vF2fI7Og6
hnV2H7o0X7nizFhV9zt3D9Veg2IoK88SB0ZsJAUfLdOpvUG/zMJ9wnbngdvr2TfE3lWEiQal505X
pec2TWxZCZZsJUREx1zIbMMfaR/cyzI4GmCH6fObvgQEbBlOPA1J5YcgRKbJO0MJCRz6Fmb+cPT7
lzJ71mPe9fIV4UCrMvI0dFw8l027L54vRzA1Ub+g+lcIkLLj2XYma2X2hgcLOUyegCrzcN//t19f
OAD9w1pBlsT0NPN0rzzraNj5w2ObFCbBWuDYK0CjRCKwPXbVP1ylfPpQn/HkUcDaDK5vlRnwJKrI
cQ9zJ1Ra+ae+Lkfg3MmEaYEk+SHeUtbuI9y9u+F2g9/Ydn5hM/39o9buqL0JGcF00JX+lxTHoE0d
Tw8I4Xohr5FZVVmVrbnBrDqc7synx/uTv1n04v2XxXY26eo7dptQ+gaQPJpsHkPZIc4bSWlHicEs
8YaWmgEZ7qnlmVjEqxeYEdhGeZZUh3M0aavKrNnLkxBR2ylC7VqTLZ2jUxBAGa3fnj9lUqpFjxPA
iqnA2gJtvOl95P+FxQ88FfQC1DN1l00mfW1tEFem1eLji2z3/vbYlp9SM9ao2ePS38vI3ILTwgs9
UDEIPB8WplDnuyhj5w/NIoqwwVuPRvXm8UnH8Uf9+5b0ZEys1SfmudrEU1Kg8h37mCysl2EYVJtt
Jd6+3GPgkpIhzw22puVRgLLpK5euL5xnntT9CVDEjW8E/y72C4AuYHPCSegx1vp8up/DftaPlMqL
sRhY64Yuxq77pCQv6CE1jPVyEAQHerGG7asMiACH+8xe0M7tNOAAvRWf+58uOzKX19qmaYlYRlsi
bCFyhSqa7SHohVNkiwJsVQ441Ih+xAi3GeunIKjqcXpS1eISS8MkhZx3x39ReQI74ZxZP/uiAg83
VHnHb6/7W7eG5WzaSbV/D05hUDH5uptI1Y1MpwrB5yRcxwAFTboM6n7itwYVIcMFxVFgm2q0OhPe
o5WuY0lY3xPOwJRPniIID4BBrXFvEXwBY93U7ooYF+G5x6lZY5WWgZZ1ysxWM8ylzBbRoynvs3ia
atKXgAwpDmiLk765kLcQvUDgwexW76MJ2GY8MInwGpKOTrpOsjvMh4cXBS+Xb4GH7BeXAf93xlxS
dkWjL0PeCuYP4vCx5ZUfxxjp6s4/VRXbb3IpB3BFyeKdg5PkpNDR5Ib/vI1SF79kfzo9MR62nkyN
dt5ZcD3I4S/BjkILVW2AAuQmt7CVskath6pXfGfonwRWlvXg7pidysTgseoZDwYKQ4UQkunhG6o3
KnAe8C+d79zFv+10nm6OZR+oRpsreMfFNbEgnwBbeIMK6ziwHwWvzTxLfm03djg5SJggAKkzpC40
RdaeKUPcTDhwWMlB/D4j6JPizB+oafoCdA3PjTxKYfN4mzMlzIHGe3gg7W5nmJ2Kg48I4lYfGjqG
pxV1ykjs/SR6cNGpvG5J46NyQYmMqkaiF25plyEWJYUXz/N4L04yWZKBEQRku6+Vu+TUpjTna+4A
WZCVZH37NiwQ05arsfmtb7ZE2SMCmvqxbYy3HP3/zVsS44zXuKUjIION6DsSAlaJlPCI1eb5bOhV
9wZWXGlUxm9pjfDYmRw6zZt+zu9xBD00n1ceLgQgRb7InQpgv2ik2Mcbuo+BuF6JSzFP6Ht/7UmZ
xUBKOvunvOsYnN/Xv4qNQkaYN2Lri2eZJIWBJdRaAWzz0+AcmhQ7tW3c8WHGQVJ9tSUwpB+sMjpd
7y4if1jBeN2ABn4HEa5rAb7SfNutqYAibZeXxwK5a/NAJShRqBybqxAu/zk5EIBwaZVMDCnXL4sI
6nc2h7+1HQ3vIKDhfw1JQiW3uEFeWwk8Q0uMrX0SnvThw/bT5FLWp+lM+Wv/xrEWnhtR2K8F45ad
SReIpZ+vUZFnHIZ7MQUzCTL4vT6ZUcammHDVyg3dCdJpNRz7XViCt3tLG5mMC7kIXzkp9Rnun5kZ
bAmaJXItMMh4GbXlfyknlsWlbZhj1VQxxNO1IDL6EZfPmIMdjYfyph7XRggvDFChAW2mk8gkRGZP
LHun6BJSnG1d6+XB3nBfcenUdYWPl9CPt9rMHAaQGede5XCpcUwRhrUHoD1I6U6Zo5iUSzLh/nJu
Yf+69QcpmdU5iKhA4x/CJt2KYXmE2aR8uowN1ISS4rGujrUpXsjLCe0/sUYkSiOLJJQ8A9gmJapc
iitY9k0A7x4tSzdKef59cHSNoEbEtQSVBQnZXCSmzF5FWXaUtWlHkKCbSDtaksCLpTlyH2SNfxQx
7KvmOAO/Ya4QCk8/vNqTxLUxsXncEiGu25LnWvuQLXuGCdaUAjQaq3kugSMRDGNyW57xxGy1rMrD
TvaQx3+o5iFG5Hff5c7L+rGoKuObBjxjX/DuMIgCSC3Q26aUKFMMLBB8AcZ07MHQoZoIPrgqdzIf
BBs2YRBNVzLgJEmp1rTRswd8uD4hk+T0XoyQFFfCNI+96bcsWe2mqQEFnQKpq4hSksFULk/z9Ije
wUSthwj9oWDsKIeLsA1y/Pm1l/jGzzqUWNOa98RFb3IIaawysJ2eMC5NDHKNAvZ6pEsLu4qIus08
9az73Q6A/uSqYEJX4NE8lPkxV7VQQHSTYXZkdNlGOSXqDBRuWCTBruuZlKFr7fBHTUQ+QDWJ6L4l
c1B7CgRrXsMKDfdkxb+feexC2cUQ0DlQgY0ZMcU94rXXNLQaJ2dOaHByNno6qI9/xvvfVMA1ZdWf
7URMTJoQzIrAAHzk4Pi2RtYSVqxPEl/g4Wq/JfvUddBeNziqkW0hlAsPkPrJdKRzZdrGFdvnV58L
8hf/HWY9XUhPPIxtlgnZpePcT11eVkNzcg9ybRK5Oz5iNsFxRbJ+X5iGgVQZ/c//CsFx+PGvZKun
MVsrN4m106DKr4NqGKjkHzviLylZ9kaTDw1DXjosSGdfVC3zYqfw8og6Awx/L6PhmZsvrnwtfNDW
9RCg4RYacfWnWWPGMlFzPPpla+Rhns5V8VL0EJA1VrI7jQKp5FQ+Lc+gIxz/KAJ1tqB3NKjQE0/o
xkB67M1nsNkZWk2PmYZg5zCc3shnPL1Pf27DgG/wy04gO3Ii6HfroLATjVgbHy94zA8yl/xTud1c
s4wcLmGwsE4jXAmx7fPQCto8BT0IzBbfRWAkxqVjIeCtHz6mkj/859SgXnpcCegZ7JJGA0E+dQwL
PWybkHvPjwoOqNhB/BO4FUm6OvNdQuDjI1ZMVA5RA0QDEzbX7e/1ntztnh4zFIelbYiX12TUwM4J
NZ0Ymx8ZZ6/Ugqw4LRgMEtfzMdYFnHKye+zIMC0Eibvb/k3jqd4hFZEa0XNOecu55jDYhwd008Nj
Xly5AcfyjMCGDpysWtoxia7/DK0iwSueqOZpm0sKa7m3/tPKRSpkzkz0IOfAsW2b2AVvsG5c0Pgz
bn8N732SIqVrpw4I8VrgQ4JiER/l1S6oQDM420iLwVKFBqmICRrlE9jdogEXYPzX4cq7TMpgvslU
/zHew/IRGuCAJVsEZtNo/GPwBa85D0sSnOX0VZDFNHgpdF0HV3afVqnXt0ySTokhBmn+IOOZs0SE
pWC72heZFwyshaNN/u+nmedab4xfizM2IaCN4s7emOXBaTosZxgZhb44dZiz+7Y+0urPsFqv7qz7
pR2AWjkC5JvJWnvr9t7JTu1HgKlW82WBCF58LB7yZvMvEGcrG09uQMnDTczi34VIEMuqD+8Ehi+0
rkPOIBt4SX/Y41vBx8sWCtoRHfG6SzAraT7B95WNWtGFUG1VAm6Tdq9ee7Zf+o07j7F4QHy2YiY/
L+tYXgPA9FuHiiOPSsOSfc5Wv00fMmOxG0mSCwUK0mtvK53kki5/hIVJYHD/TWZAaixy0Q47vgxo
QoTvW8oEu3V/busyzs/dGy60ypljDcxiisGBv7aUBPKP622BcN4h14UHT0XbDKsrdXgpn6W7oHu/
0xbLZMfNm2436tQBPvVgv1FkQhmMWDyR+8Pn9kTguf5DyeVC1TaoCroxJ7f9kyEIJf3ye2hwoQPn
muVGyi0qz4ZADJkLsM6jgIUA2Nwt2/GGMlpfjhzL+eag6oQbXBgS9NZmd9k8XB2CLbzvr6aIXvWu
Hcyy8cUiIE1oknqxR7pMPcGGmGimQnaSFyllHnsNodqoONFfEKXFs6CJYzRgrQ4XHO9t7pGLwJPm
1k9qKww2PWq+FB6vgCl+WmavIdS3kUis/dTJv7Lrx3w5eqK7QE9jNe2zrITGJKvTkG2Sn8BfYY9t
xxK0/wyKvjU1HpWtq5pVYqwQIt4E/djLAp8SGcjYy3EXzD3jNz9EnOK8dgfeflSRcoXiAAehS2X5
Z15g5pNyLWCSE7fUb3yl2pE6BKHpD0PSzzw5pbhg8sqz7P2Bm3LvH6riqOU4xf5qmaBWzMQ3kqT7
SVcFnN4Zg0vy/+MmY3sIDJNC7feJYha6qDtg9cONGu1t64joim7i4GBMlsEPutpVWgyub+uV/7RE
MIos8yAI/9AKgFK5WXK3LRxWkrdktMyqyKhOLgG+si883larSjvweQg9g0SK63FDsJjY21qN15hE
hCCtOR//thajpCQCtamgL6Tff565L7c2iZZKueHxRILENmGlGGyIL61lpKkcR0T0DVC81FGoYwbN
8cwqNgjKinA9XFUDeZJzqQ89Ts0QQelnnV+DaVlE1dl3DgSUT2TVh9bzRiV5KZA6faY0NMMaMBBF
3QFyfDuZt3Df79S5BFviUoKdjcFxbIVUN2PonGaHWxh//mn/0rk/gIL98zpdpweMhYAV1ZYyp36L
NWO1r1jLWxHA3BC1fMe2z4Ir9is45YQpAp1Q81BmgC/MpdSgJ/7YhsC7WgYqwce2+Jo56JnYkC75
FHpgkzAJNS7PTKfkybopnR47qbW/14iEugjF0NW85UoyCh61jZV7DoftzUKs6Y8I2dkXQK+PsZ93
1XRFmI5c0vcoNf00ipevG5TIjY8rAEMUX3IlBwvyEXSukGVaeis/Mz3Wlv211MCKV7LSFHyn+8eP
pHMPZ0yvNNavzZ7Wdq4xVRypZZc7C0cRffeaGRhV+g5K3TjwKJxuvm/kbEKpez7eUUB7KS31tmtW
2KDzUKoNQt8cS8pEGxw7gnIa9pCLBkOI/YSYOfZQBhkMKzchI38/lVxEHM+zaKdlX/Ki2qTlos6e
34f6IaIQnXwJpDgIqOFZUPZWN5Z3L21vHwIAW/6AR1Jx5cD9A+Iy3FMXTn3bJVbxHBYTYneBNoKp
yqJ5RNrJdR8Ne0rmuhbSGhrQXCm/Os/At4Ks0eRTC8iLZdkCJpW5AK6LaKtuq8/p6vDPogE4JNce
yPYjsJH2locTDxErC9gweBhzLR/LeP6zXivty1sH9gSLFOn62sQof9rNcVIRi9ldaEOoByj8QR02
+Vt1t4RI+mJ6D89VMMFw6hm5qJb4I3LWt/Q8EL1IqNHJJAVefMZO4NllwrCO66Nx+i2mEVVi03t3
225OX4RHtSsFox0jcOxLouGoQwB8Wsye57xXT2OCQV8Yf9HcPZ1Wcz1dHNzWx/C1sjPdlFAI8sy/
rQbBQDj1WiA+jyW6Pr0wcBe+9K8tK+dO494Nzl1RhPiMuMu/FufgS5Fc8sRrmire87QV6I6REV/f
CsuqeGudAv3vc6xrLIJY9BfYwvqAgIrca3k/D4IJQ8N3/le9LmNnvQ22fMB9amnwn32I6DCXrlxp
R6G6B6efNjUfiYFoguhe5A/sMmDHCSsEkMrlhOYWBCinQBLlLUGR8mAVjTASyi3SyAWjD+1ucFP+
4PNrlYuD1viLLJNQsPra0U5h0M79DOemw1YVoaIGh0EIX0ByUNGUzztdli2f0fkAeHGaaxXTwqXB
c3i3FI3BqaEqqWfOLuxcTK/Zr7iyKppfVJiMElld3Lrj7DOzq5uHlvYPunHcMonJYKi50pLHyGd9
/0kaWjDVG9GodGiKKqX60+rbzPDs06AXzAwJnKOJnYIbrsYF2VlKTKbbR6tiNlBa75og37hoKBKe
Fp8fQaVdQ7oIE/pQUQezUgpDN8EnJOhXAEuiHTQq//sfOqknBQqIot6z6IcXEokANvVutTG0nzve
u/7iKg4PQ+pWWeajmAMtqPAuk7A37fsjuR8I5bDYjyJHWP7uf5j98c/qr9l07o2yT2vu05I3yZyb
dorrRPBV9S97RzvpXXUvUsJ870HVjN3So/JDSFOUjpSlh+u1oyRm1Iz+WYdOziXeohpnwDu6NH4O
OUbMTDiSSZHWr+cxsAzzg2LaBYLgRoqSRTa8axsM7YkzWxv6y1ct6zF7J6gjpqYhAoYOaDBuVcT4
pyu6koZ1jiYrf3TtAoi6xmSAkKU8fgW38+yAJJE1J4i+VX0D2R4tv3bOYKuhXXn6O1vJyB/9kSk5
dEMjKBZJCEvYTpEp1lv6QroqfuR5b2Vi9y79TZocGNHMleJBKZqLLEgMMU2AKdif2k4VxIYH2bsX
GCVyPvyfR9BD2ev842OF30T/t2hHxMFnsuZO/FMovDy31TdWUbyVnZUluL5Vmb69yicVw7NnJLxa
NoF2QGOrniG0yY3D3s/AsdvWunygO/TvhiAD32s8SOTeCDo2Rq3ONVee6qjluQTEi3hOxDOROqng
3Tormuc0CNaFyR2peuIE8CjvcxB4FWmjCwk5St7RdONcUI8Lxo88TKtd2AMl9wme/+ANo+LCLzou
MrhENcsKHGB8CbFfvgS30/TKc6UP0ovqcRvLxB/rotzEl2uA6xenbfRGN/hvQnGbNbZ51rvd+rui
KOS73tbLu7z7AL+1GDB0ETmetMsfyzPVNgq168RxfSIo1xnbfYcqw1ZwyA7HQ2dB1wbO3UHvvU7C
j0kpV+KSS+PP1T+Xa9ATOn0Tus7e/J2E91gI7MCbpXAehpo+ymliKoXO2h2PnlbrpMGeYAKRRnmh
yKrUkV96I10tonllfLjrUGQfKYbtUtAlvY2weDm/zYi5nxpfSnTYYiCNSzYa+QUVXFARxd5iTHYF
72xa0od4DiUgOmjyYa/Bk6CaNRADtiyAckNGbIh2nI4mOv0WErW6PrfXnOK01fUMNQ3ZBNX8hLte
LeHofeb+hSHJMSObzyVGlmqclH5vioUrOFkU4fj3WBB8AcnaDYrkTsUcdJCQngLTjVr2U1jp5HxO
okktWLVi2GKCBlJYYFXnSfqiWKefvkvIIqnsOPgBKnB52wNoD9kzQ09p7C3APTY9E6wSn+tzwcRu
2gWjAaWB/vHWrM4e8eWV5NG0uRgJcS6yur4lq7oIxgUbvGrpUavDekcqOzlvPBmDHri7dSQDSUrr
YumuI0581G3sKRSFiz5IvklzkKp8hwEqeOXu9ZQuWbTSGREX/4xeUMn2ha846sMvZvYfmPIrpJ10
4V4KiKAK++J9qmPSG1aMBKSPO0oxV8lCtYhW/1SqjuHN1/c7UjRgMOi78sgPQ1J4Dw3TJOH5WEts
N9PCEZsAUINpYkiDSosw5KZ/5kSDgXZzs+/8EHda7Q5aom+r0Srd4PSiNBPAy+yOHm782Eu/PIz+
LjpLqeBOJzjJ+ZW7F3QTq0kS/HyU6sqnuSYiqcTyUhfAwqZh1oNHAlokwggIjB1G6eXLI/hXE0CN
VDfUSjIluqGqLNkn5jGdin07vZKTWBjCaMEdkFRP+pOQrg6YvcJnJeufyrQZOsoom9gZk8IjbJfU
y9knGGhzrl+Zmiliy6P4pmXNoRmnSh5fAqBxrwMUatOgWd4yFqQqNGPV+N+7lD9SJRIUQ8aZXwDo
ipX/ni5upoj2SDXiSFngaIA5TB4BDlO9IsRGPaNe/x1vmRp/DEhnz3UeDLhaR1wvKwNlgXW5H+cv
55yfT93l7sVaKTcne8Ok4j0rMnU5OIA6LbaGaWzryzUy/qfpqe5FoIIlcsn9Z7431bsdfPpY6py4
6QbCpF1UB/i65sTCcK7IxuucIb5YKC7rNQ3QoBBOiz5C6v2+1K9Gc5eI0Mi46YnxOgOy6t5dFH+I
4CmwvpZhhcm6XLlj8AsgD/4dMJYWqwX8OAcCgzL1DR585oZWvUai+LLA9dt6t7DcFaxjhqAnxEy9
PnABXsyzH2oQ4Ct9zAWiJWXyoLUuzmLSeFfJdov9jy8Pnp/nQLOo/niqy67Md06ufm1VwbH3nFpj
VN6GX0sO9XacduFeT8Soe6xwKjOAmd3Lgjqn2YBUWlDyOGZgOeuuiiKv/pCbRJgUtHyNYhA+Cacw
D5yf5U2NuHW10CxgdxR1gjkbEcOVb0IIoG0LOuHHIbffCE5Vu6TVmkv9Y7V3OhhQga5daOz2Pb8E
M4UwMH1/95trSGigxzYK1Qx004GP6qkFVE8mtYkM/t3m3JFDgoB1RAb4nHyzQ7Rg13812OkRG/zI
q8eUZf1TE1ALpXfhEc70RZOcmAQM651/3CEkAoQPAP3IVxzAWd0/FbAIM04X3Lx5W1hpkuVXUkQ5
ncA+/DYAQqyZ/CPFP8eUaZ5EGvhdcGRhDrAlnFhY1P6jyxjQfRhxMUJROZ5TpmgaSAVbol2xhkrV
mxGw/kdw4FWcn54jPA03UFEjIFy838yKy9DK6UyxJUNA2nt0bL1/GQ5YZ9yjTYNwqgdJNc5Dedv9
8/E0Zyf5QCYkTlKmdDsewtcqwwX5lPbeWFCbHGSWrfNS9ROO8zsoQHwbkvViTsgeq3nSLZm5SL1f
IsYLTTPPQP3ISB1OV4NrxTHTcRWXsqLqxmEQJT082z+ZVwDUktOUN64omWmDqmhK03OTSRoL1EcQ
U/BoJcgJJdJaGV02het2sKxSM83Xb3pPPo/3GKka3z6lgovq1+GVVrsGiVdo7ZxMGXDeS2qsJcXP
xI/adlIr1TTAjx74OCSq2VhtvyWb55e3O7zwhgmVskpSTawGC79K4ibFOFjj9NmHaK71n+GiPAsY
lPKgir/2QFW4zqFmd9tdfh3XkzMK07LdpNq+JFgurp/n+U9cnAPFvMonmWDVJ+MeHISiAnFsA6lX
fVOOcl2Ej7/ft4kN9/x23W4mOkaxNcV4sTqMv5zepGNr2EvNQsjYN5S9YLUNkdtfE/9wSlRFnZaV
TZ9v8TOR3W5fBnw5DWueLc/MZlmjyYiOtNro5Qz+KVtmQTDmkHFE4CqVG2DUk9oZDTis1mTWvz5x
/s8z5NNZEf/mXlVRx3GulX9nQkuEHExAlfvlI9ZJ+n7MyB4ptPicr89VKY11zsxikGUN3mQRP9C1
H+/b/NTk3F5lciNfQ28+j405h9k+39g3z73DDAkOUGYJhpp6e5gRCsd/n2KxF6wAUcsmKEr0MYLb
cueIZk25/bqZzB7nN6M+D5nj84ao/MUPHvI91QcIeif5wppdWzSAUKWKLhp6gTeGQvGikV3YgjFy
NYceMCPL5TMGK0HE4NtfdsgMnLdxo6Qi8DKhLbybrawrmt+gaBmqEVsHCTxJClL8JSgbAlOXVio4
VmQTbw2+izZF2eULvAMjl6zqEpuVwx+9Nn0C4KYthyFs3PJt/8VJYtVBHpSHLM+rhLRi+fuI3DYq
hkyHsBg+hbL9p3uH1PMDVv4xWbic+iLXUROD5HJqsU8HdhRjCMYDEtc9g3hARc/3LM1kIbYJU6K8
AVC0TbpjGaBl04ACravSQbpdcHIz5j7SUZRwZnaVj7djLFmaB5kAVdnBaeFtAPI//G14tc7EOcXz
GE3yKcTvi6zu/Ee36ri4A71IV2h4Hcbe/S/Mw0sqbh7y5fmlgv3Yogn07PqSEraxeUj3DcltcZPK
6Lj8TXR4qy9ClChQTywU0Rw0CJzkqMfZzhgteJYnRQaOLKleIK2ocBGq0N9to+PQeIpwrgS++m5C
EgkINzHCVNsruydg+YmykjA3KlPLZiquLQKGejUorX5bbYpH/bnNyEahEnfuGL4KoCeBNwvp5gK4
TZcyAwggHyUUr05mn6oVhtPfX4tOgfyHWEtiYJVzJ7hzyG5ebpe8c5aeAj2qGhWYbXMe0qg2hBqI
ZC+D7EW+es6w049R/w+zEjzJ+YpQu7OKH0cOwMTZx9hS+UpLOI7Yyfhb/EBJvwvf0cz5RFS8dQ9s
WR49RqFfxtzYPOTFfqLGpoSQlnidLhWrv7F/gOnb4UFL1bKzXhvAKgg8QnC4zxZJPOTLjWz5J33m
AR+zoH99WDpk7pd3v5JcB9pOEPyftOT4LDJWORyy3KFkGCIkLZVEeuA7ijIflOaUKGrMkiVcGZ/Z
Cju9eUfAYFS86DqXOySH8/F7vAlqJCuuSOIFo1Tn+pfFsID78uJwzJJbnsTrLnRS+PFcABnslcn9
5t7odUYSEY88kB+T92zLYqD/k9/anvP8nb8ExoPF7KPIJqLnVNTA1C4FH2SKsdLDWt0X6Bk+ritR
mqcAIyA/lLaePM+Cq9xokggMf3cx4KTANmqvh92ny+adG/Q12uxeUsESdzetx/P6rL4Sollt9QN4
4WqkjTZ+5JQsJXLlJtFnzneAaqrkycAiuPktTc04xGETP0yXfvoaJmUBBrsF5DUuocVmlDjFlpGz
U4hTLwndvB8QKOkn0RBAnUQ25X7/YI2az0BhxK0AWroAPdpWTdd0X5ie1DowtvGvCyFy/w1PrttS
Fz7UDoyrS9teOj1jffGea3KkuNlJmTHeuKsS3bbdQkVeoLungfCqx2sS/yvcXzvAmAYR8P+2cCtb
PHoARSQrY1zt7NrneNviQsWt+AQyIRG92pI+EiD6oj48dF+h2L06XoFOHf4oxA9lDWpRNomRhoVw
+yTMT1k6niP1SiJu60Vm6sB7+WFac8bQna5sENUv/xsCRwITKQum6Jl8tdXvX6H29P0Xc4NZvLmI
4t08LyaszpjW7Xem0YIbRpRNrCRUkgx515QdYvHxJwC+gIEMFzY8ycORKZ9e6IxPf/Lsg87oIgvR
Ksxd/INITSw5jzEKiPzlizhuMMBF/AXn1GDhsaJUIvlU78wHDi+L0tqfl657/lY2udBFwXNvv5oR
P4me/wPNT+DlNad9VHiAs4eqylKv74/nTzCjLVZJho/A3drTXc9bWxg3/cl9xBLrNDWvuZWGM32u
kpYIchqEEev92lLP1ymottcQPuTpuYEC71e38bIKEbujKZc18IPy5SxPvwZJt6HjPr8N7LjtYYp3
ifU1/e039heV/2YTWYXRl6nvtOEbB6dhXPoR5Uc7K0xXBOGq/dPlzw6yOWSQAnovmDXQfESZ+e6R
PzKbMitL/hADloDMDHRbaEdEAWB3NtujXGV5YdGHf3hPfV5jHvp7Q5h6qgY6DdPqvaEl7o4u5cTM
U0bBGMXcQsFodtIxE0aQbTf1dzLhDDPPr1xxAepM/Xud4M+87ZcHGPxt4FjGvwj7nEfoVwB8hYQd
DUxP8SOCkBKvbcT4ERmY6CbUWeCOALYjyV5XA9LopXT4/ZQO+CPCdcnqibzlUEhWN1Zy1IkOMs1B
HRxnrwbWvOAlLm+b7RiVxmuUAF5ulZ5pSSweb4OrjF/fSaMQNLDX+kQRHw5iVUhvq5mLw+oqEinT
VY72+YduBB9RT7GUhrIg0WeNsX6Rf/m0mo1Wrc5Xk1wajByA3p6fFfg5IA6yXA/QJoJcyK6MNwYa
ZAFOF9wJfrX4QNeG1HtuO9HxfPibPx5zAqaDWwuqTQqBYGKiD6zFo5FR6mq/SWK+qFWWvMEDbfEs
vWvurkSd6UCcr3HDSEW+VpSbV8EV86gvmRH3KYM8NofzJF5zsFcZWcAQffraqZklLOwWqg2+Ayvh
1TJNNXJjdA3ImeAGLDLhGmTRKGyaDLYWTpvuEdWA5DEn+r/wIptgqByXvhdpFB9fXjOGBRWaO1oA
bKeiyCBDvRV48VdPWFR6FMgXSJ/g+iVuGUsgmnyEDFyLnuJvnmUHaSsvnvghDSRFTe7z3jwV8D1p
R9GHpwrGY7E4p0YbmEYOldJy0AblFGhF2gkANUdmD4hgPGaDWwVKE7LM0OXgmwGSkMrPUkv51ojl
B3uHNDo+RRWVhpCTbjxbtEMixUAmNZkjBeARgWGcNg7jlKJAglxH9OPZ/61/TBDuejBSpZm5fWtK
dTdcZX8HpihEglqUH1LeSq7M/vGht8UbN8M0VSIdXjqyD8mTPvEZHfL2chpdyiSh5WQmRd0PmInJ
IqjPXPcZdFkIzd/ApbKeodxRQZXuMaUiCgrdLJqiVBGRnk1jl9dI13i6RTtlDwiKyLKWrUgjOTlM
d9Wlbtgb/jlKi00ehHBE897Pvp+Z5ZPQKzKoiic0AkGR0NMdkW3fKlM3zhQF+RKCxlKjfRSpMMyt
HoE0ZHOQMBI7wLRR34afdfIg2oRgBUxYK8uqqZtN++9rf+gShqJn091NTNO8iwiGQUWdxtrgvmgR
Pu3e/MLGEbFbsciXucod2nJEIE4qPVE37sxRWkT3YLE2Yfdn78P/mhN2PtSRTM438kJkpjNdhslx
/TKm89NvhtnMG6wKhI+R/0l7T8vVIHLVWi/ctyLyCgrwyaLFArogHQ3W/uJImsqAzcyBLsbaFyRJ
MULKm/Y9vPS+MmM8ipTtrHNIDcAwf/Pp33bKCYkbwruLCz2GjXSDL566nqmKF3ZVyQUZveEEbweJ
zgYixtjIm+2AprR4gnd9XGksKR9LLlHeEWnLpLtk68xUtou/Vmob8aaXzvJTQTA6TmA8sPoH9s6t
T+VrFc/lAIYAWejWUVcs9jZ7tz7M2xsmu9ZSeO7ePTWCXBcJgzVXBBX80CiZ0qo2Cm/8g1mXBmMT
fXLvfxeZaex4VxFYA/WEbvxi3Fy89ugP7hoa18jvsIociWyI4hON69MQhIekhWuxYdXJgIRUNGOl
JW+HMoz1A16hmEvu3cDeMwYCI8eoyi+SrY6+MYtWn13LgAVl+hRUYkwtBM+3fre2th9HyE5iXMHE
seN89yEW+YMw0NBn68qn7V+mX8xR1jjhTU4lT6nTq531ykY56ZPYnyQWJchX1LiJPMihx+oEf5xv
r/c6V5tB9v6AzwGso/gFgQLtrd4apzr6fRWmDt29+2mh5WqSzGm/RjKYPeIq40ZsCio30RRVHi4a
6iqMoBg/QAjXsnxhsn5QkL5pZuWUnzA98sziPTA+pVgIzFd8VKduxJWunSJKLQPgc1g71602xqWP
6cwjPLt1rQ4gO1/ZpRqNupVM7UWATZc/jz/aprym3BwDfX/nXNU04obnK4RmtPMffivV1QJHp0Pz
2eB972aUx6jmuSeZzIq6jGqpEFRAIwgO4aQo1DQrPj85nd4hoQBHPt+stJNkav1crSIpihN9MN4c
CAuvjx1vyQNCDy806Ih4Fp7m3GTaiyfObbaRjnjXxLPSZGsnQssdqz2KUOESgkwf2NryIbwzNp0L
ufI9ObNtGD9s3A7R4KkhmYu8hNNyQgvvNKmnfQuBQN9NXkJ7Lt6rCaonJJG5RMlVcmEhYl761JtV
mN/cXRFv+Nr91yci3kCpl7XFQicKpvRnV0nY5u/17iWJvIL901lICLzxp6JVfe6dKZjqbT8NCGE/
gv8j8348bU7cyIkrHKeVT9cbVxtz99FnDErDTlwtz0pIdlomY2gNjR3vl3WE52pUReNGTXku6Gy6
d3bhkRB1lS51EXp269H8JqqWliuuvvn+Gv4LOGSYFuLmtkU3cuuCAUnKJre/csQwJb8TgJidB/Ap
Zi2GNz5qw8+ikLpyxmEIjQFGbt9fNbJiQa5XcqNe4IEmYrBndeU3+SSabSvytq4B6VduZXcHMOP+
p7x/OGsTIk3dVkWz8zIy5eN6r8voEZSlMJWCutfwXM85AQI4Mzv2lgCT1Y7m5TNEePWN325s4E6Q
PDvpcLOR1N+8wcVFMmuGYhLTRCZQtq0cxLnlmpiqR98w+FGERC6wSHJo2fc4o/UnhbyYRM95Kv72
HgtRgReaeW/Lu7OJQ0DZev118CmLtSJzLob+35h9lfmb5q5GP1Ie+X3w/J9HCusbd7lc0vNZjV7U
bSTNWAJSaIN6qOhl841mPA5p7yfdPVjPdjfAgHuEHgtZM8sWqipsJx+ucbHYAD8wa4QshVH26UUr
yJ6V8EXGkoYlwBn+HEVhpuDPYm+Vvjo1GKs2GXB4pwadwAOwWQ3+UwqIixk+HRe+ALCNX52R+aId
1mE1DO7QA+EzlEk/pImepx0mtQd2T7XnGErzWcLO3CSlhEt08NVSMXU38NEI9zx3JQvCirzH9qxR
ACtwUVjjTwLK/9lPPWg345CqFr2WgTzK9DypHVWSZYIAimPzLs6Zf2GMvK4SDuC+mP8IBDfKUyXR
E9OwQFfzbDC8oZ4ewExVrvGrRqq30EPZqPsjV4CSmdimJCmlN8gcUPbpJvbyydivghpYN1Kvtb1d
/GESfS6FUSdCC4rawHH6X+Zj/2iFHbSsDyla3O4WpBI1QFVcI13psyAfWZc6kCBV+IUy6m2tQJrE
J3NWOLjeD1CRzkuhVWTH7fnvXAx7Y6iEKa+ffokoQECm5+/gSKp0Fu/WzO3VG+9x5skL9vCaLJLS
JfCqCDF18jtxrAbzopAI8eb+gbVhN20Vn8AF1qJaK1WRFjIY8wstf28uy4wfdPVBHZ25uDIMQdA1
MvBxhwZXNgrg/EVYDWj86ewsK8WffVT2WIZ3+ORpFLWle5fZqWVltxLiUo5wJnZ9KVNwq/o29I8A
iLOIQZZqIsjl+qsQDDkAeYP1xYftXK4QMF9zjtItLqWgULTC1H+qT8+MNwbDxd0r0pnDZbssTmye
GlGD1abOHeVwaHWDgUrW98xhgo4jLJyzObm+cpSAJcay/Tl0twkqLILwb3Nn5imcKR0wfTlJtrNs
shJLCKkiL3o9PYUYPgMp4pasjL69HI8aMkGqIK977jOjhUgAEpYqT9ZECiB7NX7iu2hlMjrbmX/m
XYmpHsqwQ5hzDmFr3T0XT5NuwE6fR8LyvPm7279I/2zNeU0wDJ+OXDIkxPqOrIE5kUvMzIjCNDkn
0MQjcPB1fxLX5cJCY98lSsJOg2fYelW45gf+Vox1q1IOdXH2j9b9BEoacLM6BJurwvdbOyLFJ4ub
CZmHD+EAddRkhUFT5jjWHf74SMIdg2V+1GhkuD4qF38e3RLCd+/Loo4XOWNtwwL99LLGUpuqKgS/
dUr/7qHAtU17h7KZgfhkppFGqnEpiq1cGcMB1yVuoKIk4VREQ3uQzbIHKZlzYj0XZQqaP4gMVmaX
bG5rszRWU88hfNH61XFj/UjEY9glm/+/SvNVY2YZh1zLThX8ewavyhfNTqKXAbNPoOeQTNyYpvao
Ue6yE+tBppc2FMzUwXqyMW7kJ8oXvaX3rJEDIui2HQTwThcBIC82QnAJ1gZmdDZ/D39RO1cOitsB
lbl+vVVSkCcDbjCgEshVMems4SKE4fBtU9Sc3IyyCjuHGNL26lH7MhNIv+P1yu8xjG4Trm0MdGhW
6wHQnthDBTIGjd/IBibZtR+qu5+tKjfQn0agZTPX73RuLAWMyeokY3R5WTbAVijvE6WuXUrDXOf8
6vjsGa1lkpDy9TaWVlxXyg2ItfUOqORbRlu6Cr688+/72tQpt16fmD+mG3S8rzRtSxodlnneE2m3
C8Xz4T4l6jUD1rnynzswxlDq+I9uQegjqGH9dWatAVFXznhcVO4/M5QU914XypuG46btE5+zzTHK
6RunpkkgVDtYAWaT4LOp4ZMKyZMTrVUq+wxfa5OB/WfWNVBQfCyodBxxFMi+YC5YtVRXR8zJXf2j
xJsx0ejUq8sevVZQUT/3bcjyeub16m3C17fc1xS0kzEFdR9dFbGbWWQzuzHLjZR0OOwsGU1gr2Rr
+bzVzLlEZPw9msH/Ioi1G140roDnVgInTaKSE5rTW34KYv5PSlYAEfnegJb5PDTBy/Ekq2WNKLZ4
SNc8iXtGRSQL65bDWRdDPf1LDbaPat0EftEHPsUtwd/XlCfr3UJmTCMBwUY0ap23t8mHkD3DasOg
l8jsov/MIBSt2tySFW08gGCThVv4pmXd3J6Mi7XRhS6vbH8iwCbdXVQG505YrqKyKP9KKvpk7/R0
YWvoc8wrzk9g7zhGS6kNp7veGdTkdWLZ3IEsgOjg3Z4ORkgaZTnHt3OQhOOUYGSu3RG+G1ortIWB
HEcgJ6ZyG39Oc12rKh6L4YzG/aHpzVPeMeCTN2o24TMHIofTzpwXRJkd98i6sKMScZyG6GTe75LW
B0CGd2/HuRQumDssLIWmYCooTCqTUQAH18spl5A1DPCs4kIyyAhyKU2/4EeD1pDSbWz+mUnNoKfV
iXA3xyCht1cEf8yxseJtyevpgflpKn7ckqEiVseDbQwonC6qswx6rF/iQsddAOQNvuZ3Fnyoezkg
JbNAJjGY1vTPFMmcImmo1+bD0+xPJSk8sv7DjloyjZyHDlcx58U0TgJ79fyIn3S5WQZxcwQ0MVrT
08hsqXiVRgi+dduY8WeqnFiz4+N9Ya4WcIfEkWXYjl+vXEwNPFAxMQRZgNUxM7Z3WdYCwW2h1h7c
Zdw6nGrSfbJvGKPGPEny0NoaiiUkFpX0J0wmJeSrjPgBTyD71IVOWv4vrv1otvyrFO3jR1BxqD/k
ZcwY5zMzfZ0IR1pati98ufz/LtTNQHSueXe89H5uR3kH9WVTSk01bmoA03i4aQst1XG/mOnZl1fn
QKRi28MN8WAFORtjI8lCH+BaaOAhmn5irPGKaRMiGv7alwh0X7j7KmB3+g35AdCM4xEysfQOSU9U
lhDSvjmDT4i1OqBkbGLAb9IHByoNxGDkera5C7RCoDuBBSVH6RiU1ycJY4JKgI1z3lejEwBf2lPQ
TuJeVj384lS/tDdARTRRGvJi7wzXf81Fg2uGtMwy4iA+FYC8FA+ocHtFnimqNfmyxemRddK2Oz1w
5R4pgIdsq5g5uXxGa+6/DPycAEnfdJI/f/pdDWAhT1DZlOjNp/avWWonjBNh7KyVjvvPCvi+ywxV
i/r/+aR+xEn9wj9quImP2MDDmQ5YZVKGVjQqv8xwFozw8dlUoJE7F3R0E07gNBZAIlOSSBvzzS0m
zEyyIxOqhACUOZZLJC48FZoCaqWhS+8uoLkLANqPaNC/feaOE/PRE5P+mtwpvKOi4YqLA6PY4LSz
ikmISQJqkiMJN0Kg+7cKPFZUqnL7/EWOvD3tLpVWmkGXgVGlWzOK3i3A3BZLQ+G0ouw9scDP8XU/
qTva66BKOlw4Pid9VhAIdlsip7HMBmooKZeA7nKMleS4WBgLfhJ9gMUdOXpENBbWMIp4rUtAlCQz
1QAfNcB2ytd1ju8mBfvhZiF3TzRQNId2YJ1ouQeB7/3msngTQ5TOMJ9PiK3MRwcj1jlbDxwtkE5v
dTZRBHgWR2iiDlcNJsfjx828A56l1BNPq8/KywEQCYNGXlQApVPRof9IQcQVXwDRtNon7uq7dpxe
2XTTQHCEPkLxeq7ixZALFcmMqIcj7gQg/Ezdl2cKKmm9lcVEi+QN5agfXqbE6SAC8WiUtxtbJR8o
RXtT0k/9HF2y+h07iWUvi1Wise1ZScnUZdFxj4tuymXhSbJy6CCCFOhmQicn7JIcGl0u9X2jN3ST
qERCKCUywsEeB3IM+C/IwvoD/J0bh65iiUAZy8EPFYxAh4KlMA4MosmNTo1qZ+BFBxZY2JLGmR0o
TM9o2Ls5XrQeisfBke9KDb9Gk829seSNRZQvWmZbIelY2+Q5GkH7wwj61mQ4vr/i1dLjm2/gyhQm
h+gYoTZr/LeZyCL+SlMwmF4TsfRxKZnBx7/RtTnJiGT7Elllzi01N1QoPnluB8UMPpigQa4D4uGX
PqOMDGJ5ATvS1g9ULWCzofm8qOcrBlGXHCHCvkUhEZfZADpUtPD9PALCSyMYLmzLH8wyvg8lW/9Z
mGZYUwvabzJe6m75iec5bzWxdc+rqqq5dhvC/KsXtxASPl2xX4uy8lbAqUMd6u6peRXT6oCjh3UE
f6Kqd3mPgQ8jjQHHulQ7lBobNnZ4kqwmPxnmzTCGFZxpBmlJ6fGEgaANkVU+4D0a+AZJVTqqV0O6
bhIv3hV9wny2xWwGdwoDkM+p6oFcAdGzIzEzfArbc/vIUZ8UM4YKaVKhaJWJknFGxsFVWsv+iR/7
KBwWsac17f/X/IrTc2i7fzuFlxJtLjZHkmPa2yi0dMtTnycvi38OOQu0m8rhCKJR1EAd/yOgpwoI
2u3OEbnyhTFqafCqgw9SHkHiU9gkLhGRRNa6+2NZTKDmjIXlny/XNfCXR6tNyttnLQNf39EKapQR
Fq26EVqJuANqZ5rjDg/T+4llbaR4hn76qkEWi7IaPJW4KAFoan6s0y634fCY/aavfJJ4t2gUmDmB
Df6JOVbW0kxRdFhvkkG/KUDTeJLBD4Rs6Y+zW9cDlPDU4pHBeDZzOnPPvRIU6GDRYaI8vQGwjAEF
iMvFyr+vQ97Ps7Te2Txay2kE9gTb8SKOf0KAyfTkt8NhNPUGG31H1OhhiY9hRAx48LpLtbcnxlsK
/xrf7ZJ5q4oGPyxKmOPqzv4YeklMU+8d4RDJbuaAm2F7xU1mgUkJPP+Yz17ZxSXd9leZj7IBZxeg
IIYjeq2AGzgvrBcVoM0Dlq9hnQTb1xfImwTVDUNcbTM3cbRNTX+10NcYT1Yv6Cxt2WKZUGtjd4aM
2ZTUOu53ZBt1Prb+y/q0YB5yRfId11HI9l8eSF0nYu90P452ivxhMlR9xJrvR7rUU4K5si1s8YSc
5Fo95YFTeLtXbEuNh6sJACDo50u77hBz4XHcUT5N7AaFPYKUeReAJU2RP5/tSd/N6JXQuNcwQgLk
7nt3uEvEPnmKCvgt8yZcJJsR+VIaqRwUeT+PRPoY/4JO2smj2k4+LN0U+zefGHvxkY00nGwy5ast
FMQ9AfpyTsTm4jkts3gP5UoYazp2l+v8TQqnZMPbAQZekxSyMEQUYdRFI0jfkVEv6WuXmoI3S977
5VODoAb3k5KoeCL+vhrLkfJhRUnii6KpT+zYeVvnVfErilVXg3z3iHjMijUqB8lpOu7wsXDHKw92
Jorr3tMAg1dEPe6KlUrtrazyvZykjTiYlVzZodgnZmon6whkDOjMgtyFqamfLRcBPXL24FXt8399
DVMzPKi65UjQQDsW3hAt3PwGaId4U6XRS/IWKZ0zhDDHmAyvcMbsWOAOL7b/rK+y7enKtic0jvhF
uRIQ8bQvoRzSP8f4kt+ATddbilyBRtRxvk6q6hqIuER/riXSpEGut82bQWzGMY4UErRfQ0N7uvbX
3duc+GeK5eitfGlhm+ITl1/pEHEt72SDF8eGID5ypyFDWSInp8ZOznb2fYn2DMjyXcTqmZ7HXcfj
flT2hQ5poSsjLemuQ3hsyN86WeqkyxBABtIpHZx6XgeHKEY5gsJf7/pML7Z2UCt8qCXQKiobAGuY
/LBWkFHovHKrapz5a0fUZQhhse2LRF2Bi/dUj7uYuKZSzHxAuU8h64FIPaZ+fwRSsMQSnuA0mtQK
eThysYdwZ4U0MCzVQj0dH71jowsy5zk+KW43/REyFx7V0R78LdZyipWwbeD3Zsprq2x2DDp8Q5j3
2rgaP0SFvFdy+pUtWn3H8H2QCqvA0rdK7huK5Vr7xK8BF9z9dzjFAk5ghCYXax0jDuzZCmZb9BW6
xIFKx9BAm4C4KuikdOC2NW8xtCJG+HVAgWrfpkKNPm5mZ5TLmZ4/d9DPEBKdDCVvKPEENsX7+IyX
805IyULhPOKQKlitu/qRBln/A95r8ptH2MwvNJzGzX3cgZuXPfN0b48Q7sm7zFdViLJ83B5ok/3F
i8Manwo5M2SUKrqK27MDkVzLENwikohEMjAdaA2nObY2eYbf/fVo4R1QIfxyd0E5Vk3FGA/WzAAI
oXKKqQpteI6DfpBGhpUYeEO7IAk3K2/BZXdx6xUcH/rS7JzQJAiQafNs9BH0apysTpiL7C5blZs9
zxjaOpT4J/t8ZcbZ109k6YZNgSomaKUy+BZdvaTsFxHzpSkCHcscWrynxGRcEzo1N/1ANd+yKia7
JJjIpNc20fQzmsvDL0+OBCv2f07/P/yyW4WYkTMldSCHQUQ4xESVdRGyaeAXkoxcbs0dV9es0WKI
T1W21ckh4s1jcvHWlCI1i1W0ZVwka0oxy7mrV7LxQmH9uIbhxRYv0VurOUJQB/E3fZlz6D5ZEVXR
LZEzocn9E8N/q30/sah7jNRya/cXa40lQocKie7giPE+P22uk2aAT5Lanx8+02gyBwSlDppynEG8
moFSv8b9Ym9tJeIh7abHP6Ptc4+n37bAPVM1h0PyRO2REGlIXDow0kOLmQqHIlrMaLA5ZkAL5RW9
sVboBkx363O6FvA3v/rfzcdJRDHtaYEvw19VPDKOczez/M/9Ec+Ot826qEyl7YC+ffCOD8StYUgd
qE2evtZHwJ/eKTiNbQPVov0saW4qw+XNvvN7gvrwzgCk0ZmxGSpLibmtKQO/bz+h8AjlGOwx6JHl
ItZYm7WPSqxOw58plU4N/McKeYsNjbZQTr4jSKNPNeGq3yPnNPR+t8PVY15ImvFsDoSWA3I3zL1s
ovJEytXKuNWivDmTog1vDp1mHjXXS6+zEQ54q/W7FuDQ07O3vn38uyHrBdldFoNX+y1GWKzfJZvP
ecX4uUmgcd6qsT01ncf5yToTD6TSMYYHodvAgvvdhIgCOQbYZMxxju7NapBHs5yZkrnuokfr5I6K
0NbkSZeJ1zVUT/20Z7SSQ0ZUs8eHAHiD/u4wcMUzsxbwOcip12ljrqNjFohec277gGDB7/Qs2mKe
J2OLQXcDQ18QXFD1GXOaYyRLeVkb5VGPTn1UK9O+2hN7doAF9g6Wr7+5ihFVR/zQ90K0+S1lL/vj
ssiAJPfbfKW/T8L2vhV7PjcOqtY+AKwpaRnR7SWF1vpI2gZNK4WYWhTDMbW8alz43l45OQdbjKTD
t9GOxLpmisVYWh3G9ub7P9y6dcQBU214rEGOlSn/WPYnJM4Ox6ttqfiSzOnfXhW5JMuw4vzueuZz
kTYucOrz34/Q4J2Rvtmk1zFF2C7M8EvFOIhKmZG+7/X8XDXJr5vH0AnBoHbWaSkMcLwVX9KOhuK7
YnIxA0Y7neKbNnk4Zy8jj2AZnWv3N8BY9m0unrRglbdsPn/2LdwObsCDwfziP6FCSkNDlTZWObKt
8XeeSgKmS8fGX8AiACC1MR25LGnkf2RXAYfPvQdbI/TVVp6K2YwLlrdQZQ7G8Ih9XKEbKTjRzcJT
LqhBCrV4oo0TBzom8wx7vYq5N8YvOcAv6Bky+jWNUeF7NZ6hgma5wtu/aEeaMvtLjli0hCy6piXV
iwLF2/icd1fAFZu2htFqwKcSPrGUOZD5rkgu3hCDetizwy4YcXlj0YbQVOxTsVYzSfJVjmY9BYtG
KFkgXIz+fzuSVP4JRnv8/NPja3uu7OVWcy1oKp3Q3AR6PFiIhhqsEgLMl5e6ipOYKCa12zm5/uCs
S/R7Z7OQu/yGQnMqGyn3DxOyQo1vMUzL6+AR23iBU8n2UsCLGtOEyEzIVHZXwa0pshk9Hti399cx
Pc37TSb67pk02ygriuMdObYyvNrc5YfFnwlG6GulvRnSamKW5HvsYBxUzy7zxmKncbwV30aP+pN5
jSH/jOxcO75D44FlgVzdPKZ5HaKsF0ixXiwURLNKkM/zQQO/MeqiDqpVVybJYV/CMPdVwW5qsMYr
4f+C4SxIJXMCqkYmVq/yqlm7SWZG+6XWX9bOSYxUwu2FWyvdotnHoQuXmU8iAbX6KXUBPbyQ0pxC
lSOvCntGwueELspjWzmsz+wWKmK+W1qt145stKYXbCjJ80MLyLXLRgz1QVM1nZQ07m28RxUS12UR
5LmN5ybm7JJLZmdqX4KuL9QdTOJwixFvyhz1+a55ExGHDoM+u7gOCYXYTWNEn3YZJaIzTyamqtPl
FgMvMvZts4SYv8u36etLYyGkSAX8ajMvnfJQPzJXeFpnRwpzjx4ieDu2D1hm+ZzF/zU8N5YoKUFV
1snf76BBfR3OtSCrY+LdRxmmA4DeLWpKkVo1t3hus8K8n7WIoXFWv60CwL/sjhAOWLjyDfjTVBkO
Kxyl/LgtARfyu6kR3EwLaf6vUqc1IRuIz8sYDZjQcGhWqaaxzZlwkYUyUu9B6vMhr/BrqnSPgknx
pCbngxxA1/n+Y98lmP5OTsPUK/oF4b3kfha+P/6Dlx2HHo2UbA22GuYSFeKtXnYsEUgkV2vtgN2S
jOohTHW1/6cPJpaRL4s3oUHHOK9Vs3FSZWITH9qS7UUXnbYdPUYPA3UDX5RazZHvCahflmiYkv4h
ZzxaOubWb0fB4jZyD+1+J7HtVMDhRKcPFFu6uD/5hxo4BF/d6bWlRRV9Nn00vrWqQg1y6ucJl9E5
3JyjRdGbxAmooHGvDlHb2NhImYq3zjTn6SU2HJkRKw+RN4ZQ8MaDBr2cyatpym3bGEJAeIH/ky0D
Oyj8E7cUSvvYvaS9xILjw1UqV+J/+AbeXmJ2+onZWBTne6LFZ+h72ERTy11AYrU/KF9+Ff6xLZcc
MhWjXsW5m8DfAxNK1GO94BhNklSZabkck7jsDCjiulzwDKZEL46aFL/f1iBHUfZQN/yTGd3I4+f5
Cj+QcbFX0Wq5AxnrOOb+DBoBAJR2rrEzXPX9JkgmGD19/9RD2kAqtna+kpZKYEq7xwC9F0cN5nx1
u8AlWrXOmTHh9ZluBSCIloZsNKjU2M3AYfc8tXIN9c0Xo2ctMv0iVJ7C0JSQEcXEE1H1xSULScLn
O5oHQfjDtOw6DtGguEQ0aGf8b8bfxNWXQNvOeZgaXOJIjaQW1OdXxLkoPuaEEr+aUEKtghmbtl7L
htwUIhuhGhm3RZhRca94LqgyN5dFAOR4V6hNdEowYI3u7AlNNdFX9x6LAKVd887j9f0U+1mw2z9D
mVNYLJqKU3ylaxGPUBTfKvVhe8+TkKfgOv7MlD9du2Jh044c7E4Ib+fCDmAP5LNQMOe1YCf48NKM
x07umiLlXZ7saSmjkLoffxFVPtpBxIlmdDx+KaEWWwG9A96f6elQz7cEcKfvKT1iZSAolCiHKB6q
xUvo+90NVlAbfqpYvMthxxJezhZ+T4DCwQSQS+/kZTr//eIIMA9q/35abPPOta2gbKmo56xe+8AW
h3cUOvrkZBmbM10q/I6nypQAjgkYFpX8s75pyiuuyKsFnzc3hbUllse0TB3G1Qk4kwbLA1IPzmkT
a8JsyGvldJZwPQwxhoWO2Yt2IeLImZKA5Ulvhs2HEQLsBGfcDrfqyL50dxmTuXYZX4kdnhLNuQLb
pFAozLvw0D5nT4pTQv911dEbl57ApX++UFRwirHmYc8yZeDi2/Ficag/h1smFpLsZd4NIYMwvg6l
qlQImrjWfUhSJ7Tb3iCE58/7tNW5TMpKzdnTO3SP1avBCqwjCmcGw/kF3+p5qx2Dx46oly++OKqV
BMKa+i8WQCX7JWQYh6caQrFLsfPZhrSXXyDGHZ/ShAd0oB09UhEu+jmtEi5810XL63U2Gf7boA6K
ayaXZqQEoxcIwluf3HRIkiqJkNnGhGa3VJs7wfzMAxd2YzEatSvSYmK7cBUDtZLKHNDARgZFr3FI
a5kiGIFl00s6mdkKyZdOKzZ9A8vMgO19MhN7mShSeujQH0vLohGBbfsrAbyZ7/iQQNkl+BJ2VWKE
lZ5T83IgUsbgsKk/obvNA34/yniHpHJVRqD0AxIT7wsGpKpOD3WX2Jhel2KIpcZtVOMyA4g6NW/n
JNO/Kbe955/NBFI1sOBrig/KNte25bVO5sY2Uscn2XcTAJKebIbPhakpiWHe8xSnuBeUnRxDJhET
ev08MNBCdRij3/4yUqF5PVW226wu4dEVbXIgL6u4rqoEeTOLaDxCIjWEZAh8VcOLWfyfoVJnHnPU
AkwpZvAqW/nn6YH4QySYcjTZq94SXZz0UyYyom7Dm1l0F4DsJ7b4rBueDFHayQ5yYcba6WSJnK2E
Yh2E/VW4t3lDh0SWLTAgTVF1hJbQLMOvpkSV9TusrOJ24MUGiqN18ZR8jm0QvbyljDWNQksHHzkN
LlRPkP79qtWd7pPQdiyilUKAMJHZuV0F4Z0tGTuF8Ab9/LY0dKy6FXIxwY7/9UPIkrFxmGr8lL39
xEAdo8ohxPKNWRWnv8lh8iiQfQ4QehHYnGrWdbINDjRsFgdndzQyga88dSoAP+w/f+N8u7kq/m3y
cUp5uWH5x4Oj+5xQyI2zJT0oAe5hSJny54B+PZ9HiVbNlpbsR3NQkTa2kU2cWqlvHYSLNvxyiWL2
68eKygtOI6Z0gE3o3ZT7c75ttTZB9WGOW9Q8EXTgF/zabKh2n61CKkPmYIK92kJnKP41OrQ/dypD
nBKU3Qp3HXAC59OQDSoe5bQN3Mbw4CJYDFMdvKCQpjZdj4yPTXCKOaGlrk4x3lFOSL96YuXFPiFH
icU8rd7CZTj+GVOY4BaHrOAjai0SVWyZccqyJpS/CJwqcanYV1eunTrMI0FOCYCe1qRW65ChYjdv
mKmmE4ljaMU6IpLP6nSITDV19lKOAwe3+1i5zI7Rsjawo2PUNaGGapqw54sjHfKHzSIh5cBYiVKp
v2MkvMOBLyTzepLVxyUn8alggVY31PLxF3y+r8MhrVgpTBg7fgvF1AJ6NI5glS9jUumUwsF4uS3f
S8/0Y6RwV2g/GdZOmeQ6wbzPoeE/NEuxIxhKca4U8xUzGiO0gIZbOEyzGeb5pVqEJLoJs1w6dHwI
lNI6uUVM59NrukRcCIKgtqrmiA2uStBUx8wPuL/p5zEMQntUSMTTRvjCzv2WLn8HhJeHk4rkUAUS
+hwInEELaI3MSKidfM2pGrDDKYlX+zcT9ReNF+HQMAtxOEwraNqTta5gAJ1yBh53+9FxoMrLJRTw
MAw5UJA6UPKyoaqBp54AJw4ME6fLCGdArc+yXwjPoxId+9PdnXJ8hrvHHqcewRlrxz+wjivsqNb9
WZIIPEq9vI6tJJdWj7XEz/4sya2/Z8dC+eFYgcXi2OJpZ8out1mDDhshuO5CIIgUAI55Ye2D6rKl
OjrY7MFmsJ90FkHoVvGwzEF/yWy+K6w52s7fXcPi3k3wwMScExr2dfZBdmiq1sIEmLqtroFv3Pp+
nEtb9iVb9c29Qao1aGQVA0gm7nU6EKm2IurMSO7BOgqfHKvzBI4gMlMmnRknrExaJrXW4Nko2lE2
SZ4xLSPQuyA936VIw0fY89I5CDy298mlbxNjwh9XiWh1yw51p9RW23MBSNDLXdAncQGYbgiWWcDI
iUo1icAZczfuVYQSE4EZ27g8Lh9FaDGZjEVGcuj682iCuwxjGJJwiu5FaqABRtSGB4A/jwgEPQ3M
DSDGoBZ7v8zmtcKwLmbUDMCg+gLVhhRLiG8h7ApSOgNzky7LVvPO2x2xoIP39ws2h6rkWNu9gsQE
KXk2sMW7fgRnGmiZTGXDw3moHiziirzOErAN02ZaO89erjr2CGxmgailnpf0dWH8vs4hl0RYvC2H
NW8sv9wJHa+FpcO6+liirKtFOjt0A4tzxcsZNjHt6H9Ws+LzjhCurzK7eTesTjtV7fF+9QYaZnrB
Nh1dXuMyjCQmiKIL9r732dkG3uIGTteLXYAtTSYoV1R+bb1knDUxKcs4colck493KpfHddst4iDU
xPukzwqw/5KjQ2hGVfztGkQmJXNE5ZQ7PNCvpRp97SIHuStwNlNxWzfS+YL0vBGdBId8H0zoISlQ
0UUPuBMbkwU9+vtpMBRsW4MVQGn5BlcbubsbkeXqJ+baTfQrCzYbc4HXY8LUlpIbH0IQJ8x+XiIt
D03RwTdq94b2URqfYp7NAyaDDBGo+rSkRbNASnF4yXsI0mi6z0BJd52B/WDREvDSpwgnx8Qdk7O/
b6b9UiAWqZ0uGSN0FbPK7T+cL1BhEiM5TTMVMeVj1MOnf/LEVs7wdVNNb2sSf59C2C2tsVC5UEeK
ShHuoinql6jxn3oJDb8l15t0Daa2Z9g0dRt+1CBQj6WoLg3CfyP03hH1VzgSv63JzahLsQHeEcmS
F1AjClrRUr4JrwSV0d1fA800JLH/zAEj/JFp2WIoqokD12xwBdIYIM9dRECLe9DTo/pMd/3yW+nh
S+IKzPv/qFxfrCf5NiiyOFMw470xaqi9l20mwyxrOFnfwsgVKoaEhzzZ+i7xY/tt/g+yg/uEd9wt
oJw0S7D9KPjv+X6ibpXD6quc6LDiRuWgZ/j83+OHSxlp96BacIr2sh+Eiytw9Ve5TNKCgzND3sXZ
ctXEArDBKwV0aY2dmOj+d8mau0IFeRuZ79T00UixtOsmcilEbJfbAhYpe6GnL40Fa8LAX3CC7rj9
SCDWa6g8c9EFxHQMV6a6kSzgww1FXEkqZToyOY8YQF7IukJ4/xMWjXxvkThG+CtzkXdsOW1cNmGr
XG9gMWR7f9WL94hthVNuwvu+bf2nh8LcbXzye4BhcArF0hszQ0ajEe017Y7L32ZH6Vk2f2VIUrs1
AV4z7pWzf/WIwa9W14Y9NVIohTcZzlPDGbxO/3u3EWYvoNVCuBPCdVtGB6iMIy0eSDVxdqQJFuSz
AIdZt0EKHx3HAn0gQqxqjCqnhbtLLOa4VWbmvaGUGYXlpjsKwmSEC+I3bJMl419P5ZkdpzpX8RcY
jvxT3o8447SE4E9OVSlYQVj+4J2AynJ26jprb7uCvtvM27HjRVUOzC3TeYTSGOFxsU+166/yibd6
JMn9JlBfJw5Ia7K9M2Tiy2dy0WXdeOKpfUFI7X1xFHbIdX3vJZrkICsE99O3dtb4K4bJqt7Scp40
XU0RKhOAEI90tdKkjGcctWBE5Jj46891nHJUjmNeFiAX4Ms/NMemuCOt5YdpKQ3fu7KCrw0AQ2h7
eocQFGqpvLhqsB29jEnZ6fEATFLCnoVynD88tIuqFg3YlfrSz+qSteYfpBRSuVe2h2ndLk4dlQLy
QhQCY39/ev9L9yG2X2BhpjolSULjrYQESyry7HkgaE53pgq7aABG/0BQ5B0kjTo7t3OocCXmc3m2
4dYqRNnybmPjoqpa2nb5oeD1g4Cb9Zy2XX7EzrKm6hkmAVnP+fSGc3iMEksBh4MzeHl+30yfKaVM
L36Wpt3tjLEtJs3lWH1yPyTZZiKa6ADtjeWYHvPyyXmUi/zqtHY9UBUO+MZtQMCo0aPzZzkvuJnr
cW+I46zkKY1rma9ulo4jmMs32GEldrMy/soc9teCzBaWtdtDb7o7r7UkHrCoS4GYd/M4Ysk8y87h
9qCICP7oQTxtkinZRHzVdKQh+UPlJzjnmKhv48lCTuK3+F8nTehuO4L1uWz5thr/K7lnjnjnHcSg
P44fS/t2QW+wHfyldN26iOQ6ekBBitz1dOh8LsAtDZsiRWs0uyZDri5XcIhdGaEQYGIXJNqicEJr
wYBa6FLdoLL8y6shUGvaJb/x0CqIDSE5gmWO9yzcrSaN15JxCK+EMCDub59wC1LVJ7B2RAlF3oMc
o+tZMBKpTMxEF54dutSmth5ZfRnkjdIB/eFI7IdFj80KY1f1EShEITkSCYOKgcdpiFMNxAadsNhn
JFK0+xgCxywRS2lbbZTCejj4ExrIKl4B8IR6tB3x90uMmxvU02MikMF8JeDg4yYGr2ZK0Mldplt+
6i+o9+YHx1nKmZkPeHVrliiUz0h+SYtjon+FoBkqRB6EtkPrmUo/aPxLYspEbAQwrgJLVHfQTiIo
EJ0f0oXkxyLV8vMjwbo69JcPY5MNydYU6KBNx5YXKHksHrKK7D92TElIWqROo8mxHdRBD/mc238B
PmNnOIaF068HijYRDIR3eggJaXejuZJ0jE7T4QnJRgoC7J55zUby70J7Fp52Sdqp1IN77hFsbNB7
yMzx4RgyThtIYxKr7wvh4op8YVjt4u9qNia3L3rvr9D44J2uJboWDHrJF0afo8vF1OL83Tv0+ro9
Rmh6v4JG0vlbweTmsY3MknxPhpHpvik7KcJTZohAC7F4QmEcJD155QtVZK7q7veeDAEO3WSZ4Gf5
4keCNpey+yutDjJCPWMYkGq4K+eKk0pAOvIviSfnYjz3+hucWHM0LkZsrPqy9v+F+w2x1hPjVkXw
u5+IUMbx+j1S5G1H/XeBHGuF78waED9y2JWniwHhM7MIMccGxW+bRIlHBhm4w/7PV+repeQZ7T3m
rs67i3al7F6wDU+u+qO0qpxB76oaRTI6yAuJ+/YQOVzRhCq3p6wgt4oprBroZ4act19HirOoMnC6
N3ee3n3Q8HIKW/JZDONxOmXKIAhAieWRknjNM36WxjekabrnfKkLkbmoEYmPkY3jWuITDfuuOJWm
T3OygD0yV2Nv7t2r3wOO/jP7nwBS/lKXco4PYrozu2w91oGf0mnkbnOHF9iZVS6elOlimUSNDeRk
bh8bHvv0TacmuHbnvLM3Xu/NEL3W73J4CoYfXinQ3VGGBDWjBSYvRxs/flP415FyEjHW1FVzBRa0
644yfK6N/lhl/37JJhGQogxfc8PhhKFc239vD7jaIXPEqiQhkbgI2YjWgDChEIhVg5j86261fwYu
J+uMzc8U5h1lnqTvyszgoXxFy9hP5SUNhNHJP2zujF7YkOAGPL0Lb3cw6ca9tpc+jiGnEOFzFxFW
BXeigoGlfrlcf7fJ9l9A4Lv1aSJvWaCuoHb+fCL/4scQDxLjEEHLdhFBinp0Zp6eB8/TvnezlZcF
KaJS24Jd0wMfHsiH2AkxIqPLtzfOw2ojmwtpLdXnGDRJZUVweAtPqC1/fJ8qmeNmUJGCTiPeqEor
JzK1VzvZCWaUSbe5ndiiyIsxF6wuOSN9e7N4DZ88jIdchmQoVBD98Fq++GBg1siB3YJeONS6NgMX
YCtqS9He9mX/fsgezl06o+3kqzgoUEiwKag+Xg2yK16ZGhnBKZsott6WEtYS5Uba+hE6Pr4zkhs2
uBlqO6gwoQ0/BvjWYVliqbTG5fpO0WGe0bVqcUm1uCSsRE2HSiqZZ8opO6/SqAMsKsz27GWGTywt
WIk9W/guOVPw37BBS0/jxyxsyYuqiieypcmWxmqRq/kCvImR0CR4wrWyykcVo+ZCyztCMJmdWOb0
BhXjbbGpQFKWV3HJWigKVxVYFJzAdiK8m0HwkDQBYilkv5Im3CLePPVHmIbd9L59Z2m5Nonsetit
p6o6WuzSQ9DzNBN1O9l4FTaTWc6FUpJj8r5Cz+EfKhSaCmpRKRRAOrlFfF7rxUPNhuPvVP02ZKgC
70HNl49jlJAMidtI206AqiDlAIOX0Vsnet03BFVzziAttOM1m7wgLed7naFb/z9kqBJSZZXSwiIR
t0RFA2xtdgujOPTrMKhFfLfHnBLxm9ArmzwSN/X+4elevZ8SDIPnYGNBEyF7tCWuoFzidXEM+KEQ
/RJTK6B8dbvG9cGeNVKNs4pu62ULPJLVB0HIMVZWhbkXsWt4JnYYiUyMsVVdzTZhyTloMTFHJxUf
BtP4msDCmoIp0mTjMK9sZbz21pe6EIfXF0yggu/PdJnlTzTTL02wpoeHnVFZ7ZkYhw+UxydOV14i
Jedk2aX1Vd9xNmAR5bxPXQbGix+Eevq6izJMO8Xpk/8q+A/Zft6m7ojs0ct5BbpXIVo2/B8RraLf
NVHsKIl7x6yhwroDq7PIEEDGs7gDloHs1Ya7/ItTT11Ixj0GajQh/RNxhw7NW/MHXybnx5nEBsak
G/XYJlkXqsfoxcol8hDIF4OpNPpK6mcBHspafTB6cVFF7zzIPkgpr/uRHvXKUzKmnpg7ThRsLaQ0
f4NtGX9z7nn/ElDYCxM0aOTRhLlwC3A/yp54GxlELuapaPbv5FTdTUjESZ64sZM53+mEQvPtSezf
Nt8zViTEApKHqBor9zoNjemQxrrfGBInDr9K/+u8kNmRvw38wLtKDSg4jccqanOAkNoE7fYL7mTw
YeF7q5XGm+HG3Ntav4ljERVgrj7eXprMGvqwr9fTM4Xip6+uk6KQi7k98wVLGGQVFlPu0bSRoVQG
ww7ePukLDDQ2t1RGjT3nS3v9kGfy4KgYhKwWdy5x1c6Ofz2Kuc3FkZ48Lx7VUFIKDbZ7CD4LPV/4
Ra00UpdBid0lcuLllnmGNaahezscukzdHGmERsNetHRlwIgVBweZjsB5jRvBTYCYLFkpFimbtgqQ
6JJvls6TE8J25VXi8I7skvJ72BAWxC2N7Rv5tbezZSrv+o9rYn2Y0kqBYE8cdbbJK2uWnNn5TBGJ
gnM19mqURpQ0KmhLJegpRiELo3laJk+H+T+FM1lITPCjUELlMzT8f9iDmRnPLEyL/+0HBOjOziV/
azH67EgRbvXH+PYyp9OlaBGLPkiAnqKZx9Hyg/BlYdwuIIHYrn8v9SrQPq1W5m92+xSId8qFBKm3
FVam62pFbU9p634MmVOokh3/Cvt62GD1cUDTv3nnO31YK9Z28rLjxwd4uaPmfc/Ev93J6lycPZV1
Vc/14gbAMlxMFqOi+iyh9oTOIqsJbel3p3aJNZltJ1FlERd+oEw8P+CKpYJ5GaA7xTd2exaEd0au
HBY45MLLLPeLQi9zODC2WNx33kbk+IzaxaTpP4AqfGl1B2XQSv+UhhrJf5XqX/n2Jmx7JJMasm2E
dILRzQPtcd3uZFzsVIqADMA8iGdevfs3RlDd6NeEOt9bcICVsg18Qa8/1HFAXycPv2VXN0U361Cv
bGhRGYGrEVAyVBnGsj8SRIZiGog13bQ7JMRMf7M8GzF5sXzx9NgumUooYITH75GAxjgCrJVaQear
wrsxmpPbCzfwoTDKPnVp3kw9BVCm+5wOkyq2xSuOyaMW5R/+cyWRw1ZtVK1LBoC40gNK8uGjQB6Z
LDvp+8UfVtI3dA5XfcHEZsI9ieX61/oC5MP8TnZbxNGqRp4o6N7FpOPRgZRwFHb+zZOCvDJ2cxrh
JiH5pdQYgRm+3AcdfIsJXs/0Jb2gOh7yB0F6Rpbd2upkqAU1fvPiH8h4mjOOqryDPD7u2RYmsAjG
m8uQnXolMhfREx4KLvXeM3lHZ44FX8R1CYQdqmyHHj6bIU/qO9nuDuu59PkL4r5XTPk4OzCCOKzb
dMpyMGi6+LTH15/mpwidxEt3IP6WfqtQ3Fxf4JfVPljQlJsmafqJ8bzkVykxZ7IMDEyIy9puJ5j4
+s/XsxBkUnnIWz3vDS8xitfiXKKR/F/GdSJTFcrTGlqi5sgltK7dVnHJ3uOazp33x+/rIrZkY5tO
RkoaQMruZcD1UFnngBSVHaqAn2KRj6j2HGuCFq5hLHwgXYSuQ2RklnQmyNA0bfWP/aeOUlzp14QD
DESrLBs+2WPki+ZI8P3xmGzY29Sd2triBSGUz/coPFgjRivdXCbJCZnd4C9RhDNNes3sqM4PCIXK
V8beaI0PZyhQkQRzXakugzBQbGZJG0nLGjfmr4W1ZsDiT0Z79bqXKcsxXmaF1YHnqabMJXtR7fLF
/nsWKMzF53UL4aM0BaZGAN5GcI1147eJx+bhAxNZtTQBV/+YEL4d7b7bRqEQZ43O6cV5peu4+bdx
i+2dvnc/KLgPRDM78/hr7kjoEdTC9zeWxaOgIdh8NA1m9H0hUQY+EFyLGlcstBluPzZBnjAkVCjV
v29b0SKPjojdtcekSpSHBu6Eo/+RjODI5K2/14ctN7Q+pPUYQIr+CuaOkDp9mar5jGZQB6Jo63Re
EM0/xO5t1wmqLpSYEcgPUGkJgMezcymbNr7UBbyuohli2AfLHVf0OF3o2Ce7hbosUXD4IL3z52IU
9fo/esGu29huacst3CRudMMrfKcsZolSH9n1ACEvrHs8VI7tidQZhDvbR5Q2Hj++mOm2ib3StcTX
ncj4WQ9zkcPEZaaTGGosw0FfjFkyMx+4YZDXa+uj73FqgrFpLPTGdZMZd+M5K4oGucpaclVtcRp5
vVmrt2wiWMLz3nw6GwPye4CdBeKCuhiVN00FoWSaOINRI3TJDRPFZ2auklHMvA6myd7bWA1c/z+u
Xh1AAB4/0htjXZOSio0sbEtlUQDrWl8gUoozjcvZl3lkgjQWXIqX0i9nWGF/gxL3C+8QV1ob/SBl
0NeQ9nTzKONPglvc53R2DX6Jwljl+6bC+oH17onXq9ohQQ0maGAwnwZbL8YRvGxhlhajLWoiCFsr
B+I3Y2ralglA5LkD5uIPzAIisMjCj8aybis1rI9WNKJXDsaIu+6FqeRxfN0RTMQTTkjRJCHjYalb
FrGdeTMcG2Xu2iOo4RspIha4Lm27G40i5vzvROvUwopTDYRHPjYtDjbQUb6hkkiPWqgV/mP4Kj3U
QoZUNahEbZhDZZkOY6EgOOHPcv3B9Wm9GiQo0NTJ+viZqrYfeDm8HFflAWigAXNkxjeI7Ude3aI8
FP/gAHNYl7nX1S4oFAC1Ztc9futYFcndkZUn0qDBKVgHXm+nXNFrNRCzeQJuP19tbDpAHIO022KJ
m5bxuZwuOlAwRPn+w277izBNNfw0d42vQiDc53uGoRFKH3otPSpZShYOxIPtMhSgfpT0nhfm/+aR
lGgaiGOyupKDfF9d2MYmVdC+2rcgrsru9zPaInST+9+KMa3wNDTlAxQMovyl6JQ8AHq4NWuc3TLA
4RhJh/npmWbHUrXhyU3re2/GlBzwZf2m51UH7mxzUjZheh001iU8EnBZY/uco++j0CrC1vEL6O0N
Kuz88ch1znPftOa1k9fIIO8B9iToFb4aFcMjUnTeywt2zW+K/XJMBu4FYwL+8NyoELWF/WcE5K31
4jXOqT+zsXNpnA6eP7N/4uGMNrSWwqgFQmzJnorCM/aWbSXfn9SWd+DTD1GWj+H/B/ieC8cwUcJT
ZGvcqhmyp1bt3y2SGWLwis6Auatv3vkHIM/betTyrIH6o3TzjtlfDcoVaXzSuQvHrRlrnvpb62yv
45AFLC+y4Kcl4YKJM0BYtIyKpB/fkFOAKJEeMssgjMMi5CQ6zeH13pL0CLjJH0Mqf7JNdAWhS8Du
RzyONWlkFG5W5U8VIS4Ckgbl+0qEmglxQyI/0HtFYToDwMF5FYB+UZxzYpyEVhYFydaK1Wt0F0af
VUq0IzoElJHkJ41mtYV3qnFLpeRb8tnvVQtdaavfcY7c+SYZQHNrDkToUoxvGonDyUx9AVAkDcZz
CjAhEou/wb6Xbm3Unj6AWJ9HYeZBKZvNPOJFYaMmt07mCZDcHr4Fdp/8iG/Zp0zEiC6/vtTzgsDZ
CrWf6RCTrYQPF+4eso8I+OPHGU/CwLj836y9QZHl+bnpl6PCb9REyHiMTXci0yEC0bqY9+uLUFU/
R+XABl5OKB1YTy4bEp2VGex+/MfbigShIPcVRqjADnvg4/SQWXTCeAcDb6EB2H2tIDDBRLU5e3eA
ypa2Ool+u+Ob+Kr5pt9XfZdgFjiIQvaAEgcrjaOzPrtdVnKrVNgUCgCrlPBPhGYbzNxqi7aMB+QZ
1BfzFd+bV922SIptL+Mih6MYAGwXcMBMdsucjJJaF954rIqj6kj3HfJA8TwxvFo3dG7OmLd4dqMk
X1a9F/0IXnm4PGQhTVO7Q45lu+tDqn0f87CfFUQDBmrmsWo94R6k+PErrHDpEZzF6RCot42cXWx3
z/2BIwkZLAgkwprIGZpOJYpQAnmpDq1jlWPDsjHUUY7EF06IEqIb3xQX4mx8BlBViVhr0ApCIxP5
K3Q8w/DgAMxifvh8eWReizRnhf6or6E9aiEieuiuayovB4PhQrJrzYaj6Cx8AZR64KypP3bFak1x
Zw1fs9dIIQNOwKhlLpJYQqFJm8p7XMiKoPWdFRf/09i5On7Z3mf1PTgjIDY/bw6a2e2kbM9d7j4u
05WqsgxUF3+QFxlTDaGDh5gAcP3T1EnnGNtaY5yvQxae7Qs7bVwPjiSyRgIwsEjKFjM0aByW9JZv
peAtm2EooJHblwbsBHX/nU/gkQBpmwxbWKo4jq1PHGCw0u0jGcQM/+bOC/9Z/fE/PjU68WqKHzd8
vNc4iSyvU+eNE02RQPpvtfBjOwa8jPmEGWaEdoeA7JlAAzYM+/lTzH2GCrNxZZW35SHmGNjyrfos
V0l1/8/32mFMIzgjHIq7ev5dX7mORT8BJnaxfeQmu/Sq8QDg11X4n1/sXXzEgn8BOrpC7zCT/kLg
BTH4DaO88wYSKXJs+aCeSir4EjNC1tRk4D/lX+2/WRHD1AbyMQg9wtUMTj5CKY9MaQHBhUgpyLiO
JIGltq4kBLIr+NV96VqzMPvhElbzZ/RwkYsromfur9Qchp6/zOcGja3JzXIQxWflqkysTBG1nO/i
wkja0lucvKPQClkNY7Jl3tlS1j7o/Kh4kD3GcwdD0ImNsGyxhW6XDbFWnK2r7qsUAE446rZwZ6Ea
68mZ8+lR2vHNsb2QgqKADRXfYLE0GOb1G+j4FY+tO//KaSyDIv27MJKku5OIHU8OnjGfCCyzEmsj
gRc009taTdkBmzIXtDDrXbFPdrcwwOb1rCvdTlTm3Ch8m7HMKk1OSeHfoZ8tUHZJ7AshnSjoaM4S
BNSraNKCwr3XjgOxcL3qGGb1gz7r9LFoivCjP7KFP9TQCjwHbVLH+czSorM0hgodF14Vpa1fxIsb
PQqTnkpdyTFrtxZV2LC5DR7+QVnTRklqz3QlhAzBNO8mo67GrW6OpzZkxzloPdyLcGanqVJ/1ua3
2Y1oLaa1qvMuHuwL1cpcb9/9699h9IXyy8Ic/geIArY4g3eXhmZBYAXkK9tvsA2ZAF7rCCld0LAn
iE/fB+sSbyb5r7pMwcf67Ga9AApjvH+rrvyij6QBUAb3srHalUbCS6gfVz9hdeT+0r1LaS5pMQ5A
mTiJcwQyr3do/fsrnmllCPjnBcBK7BY17pqZJhfFXST9g+UshyCdgpHtoMDWZK3LHgj6dVPi0js9
DY0W4KVuts8SCuVHB1O4qhYceerGUmrixGykAeUXs33h+QQYb48wFvCZbff6qK7unB7MpETZsohk
2gkAJ8upAwtma9xwMZiH2woKEilQPzm//qx9kBt1eT0JIjmRN8KdlbYc9s7eJAtj7klGlDjEcvJD
gG4YGTG5UdyT9lCHYkRE8fqaKdq/A2EspHYY9GTFeLTEC9E5YjC0Y/CKmi9EcFXuDYlNIsJJMa5T
nQscvRQDPkwiUPg1jLCp0UFq/brUjWYZp5WpU4lxAlrmZsO3MxBLJyVpgx7+n27GPqJUHgJsE+PD
c9dXzg7KWPt2JyFtP1uxgJU9oO9IzZFmR3jzZmrbEpK4zZBSv1x4VXlQ/GGoIWxiUQgYx7uVgO8J
1JWLQzabZhZQaO7uMIEhl3cpZwrbCsMERXrQmjaCZtBKcaVA+AVfw1xvAHPOQxac7UoWTKWnCQGJ
T7a8bl+Ni4Xutk9iUXLCfdWlLg6x7g0YTtkWGJXJwroKzd5kY8wz/13r9+w3KhaCYXDMMEgVOFfI
3M7ceRRn6I3Pormjyhn3xtL7QD3WXZUAnN0bqlzZC4qLgD6IhgKdWsXo7EU0LiPcefv1C4w4d4HB
tSBUHxFCTDUwEwIEXVrPg5HpspMKVSATofBUFncGiUZPWUgKEcp/3OXj40Twj0WZvo2VhH8a8zH1
C/0RfQ3ZnZGuk8W/Wu5351PF4vHaiilvzUjlKxPA0psx/+dlcJhiJzmL4nCZzM/EbcQTyxMIhf/O
ubZgNAxSn3jR7iXdRKB6AJrm8MFGBbC7dZlEktbAoyWttETzC6fd7VBkX5HjBI69KcCm80Xt+CxV
MblfVIjpAui95GuyBUEvyn0A7MJujMmB5K7rk9kTjg6KTku3i3h65twBrsrjhpUWNu7T0cu4oohY
lojRALEyzqpmKVJ01o9Ao3Yk2m7DSnA1U2YPhvqMleoNT5MQfhh7fwHjuGgDkR+8q2ziNjXJberC
UwVLjoeo70Bmxobq81qoiceac/G0u7BYxVwJtHCu4PEJEo8CikU+HuVRG7yV1cY+/vnPIydTrx9R
g1GOy0D1fP8waaRb/0USD8on0Sf0Y9SXgTeCz4KQz5ztqsn2rduauibkNf2BzyLOyU+atL9bqoan
y9hmP71e420DwAJBYOULRcvhdiVCo5HkVDGtbEB6v9MbAfhUTrM6jRWygDdGEhEoZsqaQ55t36W0
1VAjB31fPdo4ZgDb2spJo8XrcOUjkD2aaZFULpz4pR1CfsRuOm9qwNVpNI3s7EQxeDGy9LlPYq4P
+KJaQD6iAZQyeWkXzLKHi03xWFthrjKhdyVQPKikgZYXccWFJOY2ZzcYuPTCcsP6CLN+foB14yYE
zUR1k28QsaFAoLO0g8ef9Sc1zIyYf1Hc1G11KCVMmc5zLJ6ZNs61ip4FolTqokJVoL7HiZmDCcrb
J6fBJ8CtpiOJRpvVy5Qku5ujrOSHwM5Yuv4I/4j5Dj1bnVQnqrJMqaMNWQJNYOnMlWXb6PB8Rol5
Y65G7rkw3QOp8dX8g3sOLFq3FVPvNRjvARevf4KdwFPndpNxx8gxky/LNvzEZqiWXui05t12fsn2
Ihw/MKg6HNIscNofT5PuNZc77mILmiiYqChktgnScPjjgfcWKQ5htZOqABrDqJdYaDt5oCi+Cn1z
xZZ8xsb4oBwpnoXhAGTwkIvZGmqH9dboxWinwrxruW8VhRJoh+aq23vkRAYFimcNAOdvqNndgMT5
LVStU6nrkZGsVTUNU9yKQv2RYKBLSx1g3QcHgnSFu6534kWBUJGX873LSV7r7fiBXDZoPi7hA8Uo
wygFawlFtvU9wsTuZsbCaNfOc5d+HgRBFrQagCb6f8LJULgSA0p56EMdxK+fh+yWSE9RCvKXlWE5
XbE0/UN+r4zGJu+aLbNMW2psDHBmXpHRgmEPw3SE4AST2l+3aa/BGgPQKD4LnhXBwfHpeE0/JuQX
UwTaLP/1NWEC12IvEp+rvQ0hGUBZosxdbgaCrzaJEGnw0DMlMRnGTOEclHNQqtaqjFTZfWPgbVna
zhAU05gkzvGYGhBtyrQmMOLKLGmuIAyPNwnK6JPbqh9YUI9g4aE3qFc6+hL2ykNiqoJ/i2HeYG7w
tor/2cmzRN2+Jf7/qVr5gotris1fM0nTLOUTR49cFsiWzVfWGZK3Ef9mGkF15IHdvndyr6z7XqFY
1dUqY6Qvsil7OWCnM3Fj7fsrebM89rpTcfDhbDJxP5kc+HsVIQZQ+VdSYcSrOPoMZLWF8zPDPOBn
9GZbVkh7PkN2nQnGYs/S8Vbp45DkD64aZwNnnkMd2BPpJ4DtdOv2vx3OO6+EfkjmHNhpYRwZ9sZV
ZnTIAUNaYhGnZqrjvquWWZMeT7k0OU4phC8Km5w892KatglyCZo44wJlDaBflHRrvQvbJ9vXEuD/
9gzlEHaDtKdKyIdgS9+2mgW/XlQ0D4mvftmbVObNWjtQjkC9eaS2U+ovyJoLsRzwpvFCe9a5M9mc
5IwA+KEs/UFI3VvS+jyq5DeLfFnXILLH8oROZIAX/JrUONPRfzVVc7uIUw+dEj2PzhHH6oeYmGr7
gz7cMDFnMhZup/XobsaS38fE9QfYM85XsTy9EcguLYIGkoYhKO8yOdrj/ckTlZjUtT13nEWSyBcs
Dqk4G2V+URFr22neXyKhfCk2tsUKXMLROlLWcX0p0IPSe8rmnmEIQedmUYhCJ3qogTI0FxyLY9mI
ytr1v+unnIXFtgQmTQvTaYHj7uRF9jmh69TGUWsz3sR35tGbQ2XZ/JUFYYpVBPgGYEM9+czVk4v5
oSt3Ca2GCW9Knxaw3WQPdl/l8EUH+rztELwgpuOJHsmOD8qwpc5RCjKjLdt+G1HdLco45zxmNcSQ
D8OJrumZxiJjG8CLPlocYYtKGkxvQR1+tMGHUnCndYTQ0TtMVcNFoLSqc6MSFfU9TAcGMJQ1itrL
o1VL1Usod3Ir+JDysFqQmOGIcjfoQq3dmRDegvqJh0MLlLeKSMfW+5TQfvM175BuMr63986/vIYs
J+QfEfgY8JxSifys9YY2lwOTMrNcTa/ft3OoE6sFm27az/pHMBXA5tX7iFwH1+ULKfJVAKeAX6fc
4ZjwC3u2qbZpb+S8iHPs+u1rcW0cxxGtoVJTNTas+qTTfr1YYnvqu3ZQjtIpQisaULnIGyYkCPb1
A3SxhO9ODJNGpSPLNHySM+kpulIJPWCqlOpjXILMDLUC+xojhWhVKaKOdyKGg6EyWOQCMk3NF9qC
5nmXF4o33uJF+XxAkhjaHnflC34SO74qWlB3zbzMCWSX83Uz004UpkayQF/tnOcE9t399vRgIdVm
C0CmreTTZafGjrS4VblzaJKqG4JA2E2Bs6GNFjEpt63OxxW0nbaUWIxh6qalbPEnDZ6MOXW7AQKa
EvVUVjl1vbSFzD5MmRUnQovxQtEG9DpdWcplyoQwGX1d+B/ViI37u27c97tQ2VXoHek1xW/yS434
AgHY9Mwg5DxGt1xH81Eg6AhiNRQI7nB7rMulCuL4MuURzRSKlyIj7NNj5uJRywlOyNDb6OXPu194
RWklfEWT6zgRufTgeQM0MOt7/1SaXOXa8G0bzCy8+FyVR15n6Bna2BdDl4WalFdaxRYDZTG3LPgK
vj3OEhpNco5jrLfIFntF29ESOB8kwpvIwA6qdwiUbquhfMIrgV/4Lz22f3LioUHr4Ox/E2MI9gyV
Hv58DlGugooeAMtxZk/14tUn8xEVX54QQvdG2NAx7PojaiGGRhfXzUd7C61Ti3bSSgpStpNBinr9
xfVwOAZqvORkf2J2shjAGORNkXNTYm5akIC95SVDqJjf8/4hwj7pw+EywpIT1+qUe2lzgSVgkuvS
tshG1MrI7xbtU80ZvfxvJFj50AxbDzu7tuBHXcmce+6T117GkQHTxY+wkhv3z654f0vbpmrqXTVZ
n9qXO9gxONlbNU8v9WoLSyuvLYmDBw3kAyqVZI84Djd1IMVHFF+WtMfwObXKjbtQzyY9YDfNcLwq
ZnkffxcplKoSOGcHCghQitTcpNaspvulV6pSN4X9rC+jX/z6oagXrTnbBdFfs+XG62dI75qLXpjh
wNR/ToH4teCteuNgjE9+zqbhXNx60+HajzYHblOEYkQ31V8F04KWrmQqzrLOWz0tyfXqbD78SU+i
TIEjyOCrS2+YQVZwYPd++aQdjKr4tdphyODhsv/V780IrX+SV4upBVVoQrZIkW1kTTlXsGnCfPYZ
vvw8BhU1fFewaavfejJfANRKQrlIOMy8KeONM4x6wxxDnUGbD1F+nQ7JLs1WLtkDyqDNlKl+iiIE
kcB/SsLn5ZiKh0Fqk/S1gd/F5JoWvBc0j35IKAI5j8c4SLdhMFqN//YwCpA/fLctS30bdDy0L91B
XdsHtj4MvhOF6ca5qn1l2XUfevxYh8DV44V6zY+Atu3vBC6EevCHe9I1qryt9lGycG42EhMy5Txv
UO6gIML3wNp6J1TVKdfLCTtKC0LGoojo/SQH/4bFrFJPKAq8GzMaKp3qsAFP8NDhb3f+CzL9sGiu
dRH0l0oXJZb5rINynzLStrWg327vxUiks/JzAf2LQ7pJTAKF8fGyVFiUUXR2L+RUkXirqgkPaZ6P
CLI9OI6JSH5Dar6NkyM5c1zUTjI52VbVCAbLoAoa6JhPadbbmF/3Gcf2zBQHl96NpAg2y8RifclF
AkX/n/zt5L187REUaxvjUPvLTn5OGkyQJF+PMuF+r3KZTmuIJG+4Vk2Am5z8879TltQ/JOrOPX5W
wx5S+c9rODwyBeA4ZGqSmsKqBWnvx8RMrdcOXkH/D1QtV9me6K8+LaaLfVoh119cXFmKLS+uTX/d
CCs9FVo5sD2X9onk46AQ94EdaSBaECk/p+PLdt9RZfg0g3H6H/Nl+uLzD/iBM5ujY34g5wwoFVZX
ho+GbnXLAUEf2Co9z8inC7b4AOSIawBxojLnBn37Rf1OaQyvKiBkT6R2y8buibatyv0EneVFUmBx
Ga6ImOhE13eRtYGioLT8J7A6gPn/HxLxuMYpN/6TIGTIDlW5ocemuAcd1b263O/sZn1BAx2xE/w3
QVm2qILdrK8LFbQqestfhfRqVhd6grrcJfTDFmiqzFhUBmFf+DOpMoQbR/2/tNjljb/hUHScoFO6
Nb44+ZXFTRMDDlggWBRXGD5PLC7zqu3V56bHKx8Nz277JA+gAruEAYRGO1vLiiwULoKYtURH7c1t
KVwdJJisVzxKKBl8tIdDXGYgkrsB3PneFXIcqDE2nBD/fdOR3/IM6yTe79LJprTOOg+5VtwALwAm
cbhrkNt1hrjtoJORQ+tg94XX5hb+9/QV7bFeUQa1wk5vKI/WMovf4eAK4K/ZmA+6Brj/yup4pvHt
tDGsakQplBFAz/t0r6WCIjNd0U31LYtieUAbQnNUhzTQIVsMVU5FaWwaLGbBx4xRaLt7lfBhLdzi
If3guMC0tc5FiZJ0JQaxaBkIkR3669jIV2lJPgrhINoAYsV7vwdqP4RD+N38o3jPkHqzMjPIU8cW
/KUml0uW2RJ6MAzAftm1yf4QKfJXREfcnO6fPZcs6u/rcJwygBE2UfdtEcdor4XY9e9LeZmoZBUO
S7LM9W9dCrvr0lXOJDIF/nFQ8s5jOFn3FRNXd6kHcjphGLPdjjN+3wgDpekzi5d5XfUjY4yGTYSZ
MokuiHccDWST8JzsIf0NdO3ctfGscpR6+vM+nqLKFHbYsDdKRgrG8LPOFPPzvrhhmr8/fZEi1Jq2
rrg/cChSwOFv7DMVIRw3IvTPC3AFytor+O+odh96tXeyBJkrFxgoAttyPI1n3hbpLKNKDUjBouTv
XChB0Y5nf/Jqhy+fD2SQkBZHFqyhed7Vf/XvLZzinK1XajV6pxIESBiHcTUK1r259RfNkP90hqle
7fGjY5a490yDUQ58FseiXD/AMN5KbSaDb26KzL3zybVny33Ec1oHe4Hzi6yULUMI1+SZ4NQJm4Z5
R7EEajWxUn67rhkX/m9gvIVqhu9anLrggbSEx/yLAjIaLVlrn2RK3a9SyGqTHrhtRe+/lhBWNr/k
v7Rx7FKg5aTHjwd+e5Q7Y0dD8fm3kJm5dTaVDwt69QBLxBq8ou0G8w+rVRwqeW0m+VX0jC5xEMy2
ieN2M7nB0vpDney62WXhjGY9kMr6MGchTVe/SlaUqWT2gyi4Yf6txwcCqfjik5t9EWkKnYMWf4q+
vHS25PrF86f865j5ur/6C/ex8aeY30CNJc3HOXBrk8AJw4ANk5H2x+IXQbq0y+L6tLt7Jyp+CRsj
6XQypbOjUof2rHLNGj18OqNx1cuCCgx9xGZtfcs9vnfmH39OXJQ2sf/f5+J1jt9bIHoHeuQBTJ/D
SKKX0fqbNHNFWG+AlNfK6I9Bhw5TO6Gdb+bngY0ytSGkzXRB8FRGYXGp2xVRF5+qqd89omkBmFTq
tfVVmADp+zch6WjRcNP/H5WUHnZsDXMRGvX8Nx4p7m+OWDatbKA6w02y56Rl+9zB3AZCAmyCUnBV
uDKv26TGo/Yl2D84HTAtXnlY/8yZC8ypaDkenXT9Lj3bWedUmUzKFBH+cOm5/n7VQNZOVTjjuM52
qehethDpHJVyaLJb5PcCO9V0e+hqr5o+vSdIKRgJcs06KvyBuSQiwiZ3kPsPIwlQVfS6+edXKgNi
lExG8AIsZgpA4FB50kpNYsjUNmnsHQW8YISj7zX6GFLLlJuNMujn5c5SziFtc3QnE98tTUZQANJS
NtjpEdhmUnTR29Rb9mS3yOr2Lf6DVIUiNOrQwaQIsiT58O6gw9IKbPFHhvufZOToFm4NAjuS3bov
QoLbbkz9q80DIvEiLEUuu62kERFP5diewUuk7roJQWMiLWuGx5xdFwMclnsPnlRbq+pkJw0eZUiB
MXuj5Z8oNjiGCs2Disyx407g35Kwv8tJ3QEWvZREelDbCqILlPmmPigaou7mHv6iCXcoWSlBKoXs
FQvf2+TW4syoj0JsHYJ/WddCFCJeZOb+UyAy05tqJt3ITlUlm9jN8QxaJOUUCjfwHzvQkqMOji9H
G6KkBtJFbXlaCHBmYmkXzD3wd4816fbm4p6NeS0mkvMWVd74mMIuFYRhUi+prbxrX5OOujlOkbXB
O+18zgP58N2Zx4qCgQQCupj389Qzt5bMDYxJvjZwYrc4o+30YuYQDp9yZuCGpNEQk2L9QryFo5W/
YFuhXQi+0bU9MP9FwwNkP0FW896pa5pPf/QmS3+UWhtLz5/M3qeJ0caWRTQGEoQgF+hj6OFKsjmH
zGA/jfer0MH2+eo96AX+8Z5ETrKMa2aKq1mbFy4eLlzIFNpi4DP4F0fKMIb6I3ombXQ/Pi9rhcwM
twrUMwUh3jLoEJ6ex2f/ISfTfdI6uN1fIaNpoIJBCGiu1UA4vM6dKlxbQgxxA1A7xjwrqstP6TiH
4yNwMUjPmKREjZte+W4Ss4Ims2PaZB3hxxLFgvF7wGULl269O7Gvrr6CZKkQW1EqVrEFZMDXLHYz
awX4L78X3r4LZa7Q13gUu4uz0Lryms8osf2pefiDbsk120dLGk0MldFzb1MFAoma2bU2jUkch9Tj
sLA22qwAxr96okhOxxFm8eUyWBUilMJXDdnK19LnOElEHBI0Rvu8ZJFKvdix8rVwmPCcKBQnw6ro
mgIHo9SWJqbBwYnJgf9uADKOJP1hMs95aIS57un9/thpsAXVamDCGtSz6xihOK2/reZEWyIrmTCl
h00X8SCZ1BAlqnZTMRb4b4vxOpd0021mkEL4ovcZe8gxDtBQL5/IMHnIPN+KZzpnuRkoAC8/bIiy
hQsU+kb+7NIiQ1B0rrPNQt8wN8MsA8X0RegIcsm71MCXPwWbIlP78rhE9zUCHp2G9Q6s0bDuuvRI
Wbhjb6htK2dQZahATXGcWcNcQ4nrNTPMukcNYB41gmZYApSacCNf8bGYAMEOHtS7fzW4a8liTrux
u8eOeERJ1dT/M8ojt1PG9eJmkKfrk7SgPbNiU1C9bSZShQHCHuWe6CNhdu/CSqDuakTME87GCpX3
BlTFQE2kxZOYyuaKDRHMopqQFmI5JsFIMdd+7Ft/3gz8RK79z9/1GIYAKgcmnSwzWfKBvDCmqaQi
yQuLSRFEFQtHJjhfisJv1J1Z6x20dYByYDMpCJS6CXwwTo1bqopckAlysGg7lbmNODfTGgE3jyGR
BGrWGAJmu8HFgJpsa7Iw+nHU0UtKD8+y+CyfJr9425X66QhnQABXsQ23J7hSf2jYcVGqJzQ/yAsI
nKhibR4z+XarzXq970nyF4QBLSRJ+jxnrkG3UgmyYPqv2Ew1viNTC2PWfUXLn6ENRIPrXdeFU8Uh
lAczYQmgfs6NSIvEqQCMh48WRX6TPx5boSbY269zv7aYwZnBp3ItM1xCPLKEAvUSma0+hUZRNPt1
ruSjM4nUcrlI7yPSOCehaWoTadZ48ylrzPm34Dy576Bnjv98zCWp0cNr7DEFXk8AcCM6YkDJ0Emz
6z0bmYCgpT7Y5nKPnHl1Y5DpFjsEU9gHoBfXSGS1/n3PTds9SLEDGbAcIBIXU8ylvA6vT1GoXJcr
nKKJmzK/AaAIJyI4//qWRINPE8MSVqdr6TtN+zsei1NpSTE2XrasuFHhGCmqK4Nymvttuv1HKEfh
pkSfCZkjjQOzo2GOofS4Ky/8JXYl95ArLdZNKnI5MzNFeYMRWXpuwCSWmUQKI2szZvV4HPSHHQ+q
iPhBHbptl5kl4nFjh6BsMsCI2+0brrVuXTVQZdfYhaqUAqt2Nsqe0mG+y2dDL6m4yGn9BVJEkXrY
bzIP21OIZtuUzlHdAeQf8uvynG5BxcOIUlJ6UmK7/7XMqtzJL22CmUENS9FU8Coj4ynM71s3hB+W
gBasKl9llcUoRCU8qQLNceHYGI9nBzQGc+yMOfXcyOl5FyomnF18I9QAmFi4B+JkPCXlw6hSw6Df
w9ilkZh5TSAKQ6VtQzOltfniwDt3Wa6gZiMaBPaRtWHjHnMw4wDvvhf7bYczJKe1bEIUgTP4sjK4
5gVxWhZQjmcUJbCH9ajbzY55RSrS4ZGaTs3E0EQeOY/7j7QTszKpZRH37vySpiBcboblEeNxrydz
kUzfisJl259jprehqBJ4luYlzdGag944NvxlE07Tv2tOsfR9LZVlP4X559UlhxSp5vXeWb/NMGV5
R104MYGGipxGNIBRHhtehBmphC3uqXNlcKE/oQkxkijKO7M19IxsBHUcWDBQ0w+aepgiZX0vrFq5
yDZpu8wHtKvqXcjv+ePPqAuG9WyvIw7LVG6XJ/Tkm2CV/NemxZWK2k28jOGL1ToRvycEj4EDkCSb
fEj3jmW0wN5vH+n09AEaXW0dPMrPyM1HZ2BvJ5eYBnsxPjBL91vgiRd0DOOmOtTlTJ330d70vVW7
V+Dab9n5zvR6kR0sV8LofRF7VdyP/MDdUw/Y2ym/kGsfk+cX2Vc4hCHVNlyLSGLsJB+ggwGH8EwD
xFtI89mdqFPYsAdjZQ6VqfqjbWbkuVElP/qhA7Mel8WG17OA12DH7uaIk7SxBrLJQu6HMtGnfqYi
VEO9/SUtvL59MRjylCtoY2Edg+9/rSZoyJqST7at+bJYDtZFO4KcaQBzuZi11ESXnf3oAeMo0PN+
dlOgN5Jm5064MV7IONaRYye2HRadR75EAtkVg+uNfHV/5C5XMJ84pLfs9pc9j7JBL29zhWO//u4a
Nh2sOMbjqZnEP2tVG97ms0WoYsE5pu+9iHOtzw9pCxHxUYs/dJckO7mmqXt55GuHimpSFFmm+Ofg
EByAoW3BD7nekpxEVTftAWAoJMOHZfnwrYpRUVwQkAPJcD050+DERpwiGI93LiMFOviBd/G3HtTV
K8abhHvDOO1qXp2p8f5oZv1cc7UPEPTyEQXQZ8VRffS2XJqmj6yFXVtLAgOwbLrwSHnrTx+C2G1T
KU8UueyT3WMtMDyDftH8hjcDlv7NbFkQ9jnYkeAnioRImIMs76k+TZmgqLJrcDsbp2En2Ul3V0w8
xMKWjkgWy98EbZPlOndadrnnbFhWqkqf17RqKXfodt0LME18+5B28xwupaolF44FKSOserkcMCW0
zka8D6fUfd0DC6qhYTmJM5oUua6fNmFXCgpw8Hn6smMGA6e1uQpWfot2OTJii636SBFxayR5qQfq
pMYz/0HcNxrQxD9JWzDWYdLMzjwBKygeSLnJqdBTAR4+WSmh5YOYEuK+QK/oZhUzuKW2FBFFDRSw
APPU9tRlq2MrgQiv6pdhVu/DdTMF7o5nF5rUTMZ+K1CJcZapCmkLpJjMJg0G4xz7EPpRn0VHnQHl
b9dnpLDq0g+oztTfUKX5FL0e57UQvaK9SrgjBfEg7g1hhShljf/L3DJ93f1sMN8ybg/nrBJViUQh
f8AhF9lGnXFn2G144knIqtkt0iVuSFzBtp+A81cUQNiLFm1ACeunj7Li82usYbm2Z3KaP4JFC3Mz
6RgaX7A0ufzPI0Ddlsc3/54g9tHOwtogVveWpNtYoVyepPAaS0knVCuHrUbSk1AtyyaYrhbOVLwO
QoaBngGTJAQWJq6uWaj9baAGJpFyXPwKT4hISTvjzLxuQQmahR0ZFWK3r2b7/QiZA7ny3cNBAwpi
i7PMlttoifiItVefuxvr8Ath1F5LIXszZkiRcOO3h66WyIYXRbyhLZnw5iOAoGLwu51G045bkrvV
WbzSbgdXTPzBwzhpHRRmLV45aBcehlgv/BszKnb4Arv6tj2RvZkAOjzHxRjWRDphFgWDxs7vhOu4
qvBIYumBMayEloephv5fqOLjr33G/ZVUrEg3IFMnQmNiquOQoGYrjs5LmHyNXDojDtyAQ0OK+AwP
yUPfMMiVmMRlJjtNOnCx7Lxri0YhhNm9de4ZhDCDnQtMkBKG4upVLJrTdn5VNEWKRR0snECVvm7r
ySMbNt89SHkLFJu2XaNiZU65iYI0p01tXgVEkNSwi1H/uYFghQkowQkBxOwhM3mUcJ5c8XemN6s3
YyEpEQBb88kHufVYSDCdUYhV3euNbLxlcU+QkbNwZMbZAH3VmtqIQs/ES4pPCQ4ACJS4bCrDMsPv
+p1+ufNLWAkF/kX+5bnYonno/13+omLYhmgMs4DdhLq3m00AChgfN99jYQzNVX17gq6XdMLjnA8/
DK1LoBufARTmT0DgjuNi+oQXrkR2f8io6YXUvJBeCaD4Kl5BjmG+OEN+gSwn+7lkvOxHKgWYNaM+
KLzAynD5pu9rYCk7NL1nbGiHd4QNB7H3AglzVA8BVlygiUIUgTtqaA3W+QabItnIgsuvxXXME8eu
PAm4AY3jgWQreC5wZlZ2/hzLuAqyQZJJUe+K2PxaC6IoIcX4bX6ehP7qgup6NYuT6W/n2QcT9Nvf
UEKJ8Tgpc4Affd3oePWEAM45tUBcHuIyCHha+UZInJ8AMA7/icX4YGdVmsYHqNsH7wPubcyO1eKT
jMucnGbRJTGaiZDZOp3DCBt+MY++kNvPOb6IQxHfDxAMUkbVYGwrgKQ8RkG3InwHYZo5wFoPJvfw
xgtI4GI6JpTreKiYUzhBCVkHOr/hQR1qtQ+q3RZ9AFPC4jgUqj48Wd7+1N8cYfApUMNP7/9ZOdEk
2DwoX49PTwJS2VkXppY+Ct4ki9HuSARyYr6+b9eQQ0URBHoV2QaYkgTHWfuOqFMo7Q1/U/LrhAtX
RF5oj1bdkULC/xbzTSf5iywoZPzAJ5YZzOQ5tVoGHgIYu6gHtpCSU+Tu5n8qROoyTuUkaTMmcXDl
6EZIRBDk56HWDsCzJkM+ELmG6aSWFGTStx4viS5jcj6VKTgYlAyJQk7UojyuPSczCG2oucknbA4A
xkYBcB5eUxUcfZmyB4H7kuy2UOR01nJc5/b5gGk/86zkJlN9KU2G4LgJJcsziLJn6T1rotY2x5Jm
SYRcem5ujFhq0zGEZ/z4Z12Y6PfM4/tQjUCSxxqUczyo7gpWXw0MBh+pZF8vdg4uYntZtn7/qvXE
+fpSYj1lXmUS0cnvXLWnWTlH+yAS2pfDcxnpGhjMmm8NCVRX6NFIJEXQL53OMdM1zc45SA/emwuk
Q0rGepTD6Odzl1zeUFTL95ph0dDREYeh6IY77qXx2GsfuUHGVjz2F6lCd6ePNmMyftnwV13YDyUx
rIV944xQse21VFrS8eMBLyONn31hEs4NALKqiyer7MXL1t16S2bHqnaJf6tYJWnPPWR7iMIibn34
uGexi8HEYYYip5LXh4uujK09Ha5IRh017R+DhCzo0Pz0/YumbYlRa+5k+CyuEMdPnuUlPl+ily0e
Qk4CWrRB3n+DMjU2Ujdd3v9+wIf+2rzIF1xB7iYzJIe85kL2JSpDGeol/NglUNCkii1G44xGNKVV
Kl9aOXAIcNUyMdUIYkWlx8WmoU0UBtYFDtz/oKbC5v2HIVFPOz68rT/aKEEamBMKGS6rVZ4sfwMy
GUYXGVxzaFBo8nc+N7ZrEyi2bG1JB1bseUV+VZTutre4QouDSl9F+lWwA3Z3rur/J+C5d3sbC+UI
BhO0kmlNXcT9S3Z6clEq8TkdhXRC8XHBnZlC2YxmE2lF6NGTME2MIAKhUD+HexT65b9CojjloolY
lyMo1kmJXMSJ+5GVEMednVfaZ7Uuee7VbFktX+NAwOAQewD4WQC5hjn3waTsIFbMuARtbmI1Ilb/
ITG/+0Ov/GtmekmXel3qulKsP+UvhEChVXZl7cLu7GaUQtysI3RE6ojc4fryFbQD5+jcdBq5GoMG
de2Y1IqCODTIhVN6k28ByhGCCKRHPnV0iNGbEeXTZf79W9D0xaW13jOvhMB01HSpJG08ldo4iCh9
MsruIqIMi7Qq/tD8EXiUnaMQn2NYMN8v4mdxNUv5JBpSfGzt51vLPg5f4Mg6Rl7nMuXB5zuXqwFi
c3uxapVs+EnSO7s9DIc3gn0bAjMy1uYxnieejnGyI+AtaXXINW2Sw9jt7lr9BuRgZNYxw/M3ysky
4aUetm3Kgi0oardHz8zy2czqVSSG3gz7WSoNj35/sxdUaYhtizPdbziduQWOiGy9FXSSYTEPM9XN
S5FZb7WHGAiT7YCDgSa35YGcDlGsgg8to1NMvGn/5WmamhZmMcfJ8bquoUoRAkXDNUPQHYi4wT8u
cwn+1L0b2pik4KKljDkQncJVPGHT9ICqZ6zWCx0Jg9nAQq91CEsuLWkKhLD+yUz+L+79TlqgIInA
67AGV0jekth+CPAT9rJ4VWuSg0iK8tm9O7mQni1Pi5nf2xxViCT2rsrcD10+xnwbzsdtn13Snnwc
AWAVDDGesp1E2OU/fH83yDKWdg9k1FrTw2vfSh8IE7cBtwNhu2BT7qCntKn2ehjXHkmiBKNlDZfz
Pl46FQi3m2dRRfexiDuP8UEDatqiATF1uXCStPzX864S0+DvwOQe5fTaHRlTSeQfrJEu5/ikTqub
o/te6cm7oDLqCJ+QpIjodknAGdN1Alvtb+pdaX3fK+ES+SChc/gQN9MydtHPca+5JL6Hnu3YRl70
Wj5sOW2y21xDpHTYNyRMZmkcGdlVVpz8r4GGVQdi9YiPS1gmasaPcBfWUE0hB/A5G2Z5vmxsXKz1
BY1s4mHZyRns8BfFn30kLmSu0yPAnX3z5wm+t1owWYNd/xK7zV0kdrzx1qb2hRnYobx7e1Lq++sL
xiHskLhlKVtlNwUDFcIbMlHxhrVbdr6ZyJ+wZWgsTuslZjAvA9xzndUnukDuXrd9B2fh+VI3wkqF
d1bogigPDxC3DcIla9lI3iINI1gvUcHguh+oCcIyNPzzeMksYom3muRuUA85nPAZ5Un2AAg+05Ns
sNugiaTMeWmp5Q6d7qcP6joEzgnZU677pJaMnXfi+ipbaKV7csoKOYmxYY4OuSYoJFW4ud391XOA
D1XVEDz/v++3zLas4bV0+hutOjq2ofBO44W3JcaHt7tIrCMLVmsvU1cwAA2TpLsFoDCvX+y5Pm3t
a/Q2cyqgmz/vcTKKIjzLXeNWO8ns0Mq4OcE2C3+gQy5v8szMMKEdIihnWv2bSbG4pd02udm7yyUi
VlUjKga2tq92OLbbUWVyss5kZtPB6qjLqy+lPqUyYSB+/0z/cu153Iwnf+yX9x6LhN95xDMLf8MN
0VNtRuLb3vhxuXuPzpUR+8hGm1DLE2KNZhLQ1RlHBQ8ptH/lihhbhLgiSQBX/D2Djp3dWkfMEfEz
5cl6EhTCWgr54f+g5ZOLvGlZqRv1z09KYq2wBsbqoHsleupaYFANrKNpnAfP2/n0D24JEJsMZhnM
1SYigqKrDA2Q6DK3shRIBKz18g6phPatyXNY+OUHKpBPrtaIokuJlc2bWq5xlaqLLw6g/8LscPQd
6kACI2Shaj2GobnR42yRf0fHnIHy83rFb5jg5WvDOYAvVCFLk/sFzL3h4zWccWa8sEkTbLAaE592
kOueKsv7IYMYU84i1Vdi4DuebX9tCyK0CUqUHNS4T/H7rKqOISo3QI/prKC8Pp5U4QRqDT0dvU0N
TXezpAdIwzohJryeg7wWATR8ked4kjihYUUHVA1LAw1V3PgWfVbUME7Tu/ABi5jOqRa64iB6VB5u
ztPrQksOq81QYeFqkqkytmiI3N4yomFXOaFm/BMQUMx5yI9gxEmSeVfqgrzUSyH0icvns+ilELzH
J7Ck49zJEhgO37FUdiafhuQMRoH1CkONRzGXLPcvSVraGmaU2x3wuxz4etM0EH9D7ebdlAz4zede
91SoAQuX5c2b+AlAUhSDAgmqdpCL44YeY7YRuMQaa/+f01g+dOsGJjA1HGXiYmei/rgwxxweoK70
6xdGe8uhx67BaIMmWAXPFZZUCSIXSONflHRYTWetoXNdSJ3HU3dEPqX5kai3a1F+U3C0Oj9G3Jar
LtABtOSLvx7q5IDWeGYXPfmDwvviuIvHwYYlDYhiiOnkGN7FgygWjNbQnXjpUoO/ij6VtV/HdYYZ
cdiWby+Foetjq7MpU6BU83eMhyEcMHjHc3x4Z4+/6nKlVUieUIlcnY69xLTzXbgPcDyEOvlNexVl
7TkiqQ+HZeBABbH6Nxoi9HAUcj61ZnyVdm8Pq3OQPyc3pi35495+cHx4+Y59sAIPh99EHn6rX101
Pk96Z5wa1L44IwyrGVREi1RmnGD2Dd6Z5OHKAmaq185EAJjpKvEMQy3vkQDm4h05HX+x5vH5BDBB
Pkh2GW09tNnPYSDKtr5k7QAoPeGsSZEbG+9DENqsT2B2978VYOTaV4dlQiyHzqaPou1ed1XuFYiU
eCVlJNTx2NIrITojy/+9o+EI/eo+i7qze+lEFPy9hgh614PjbAP8fUtYYqsK6lAF7NsgEsH8zeqX
An5R4t3eRqyB5sdNjXxbjhX1ncu/gSEjCHYuF0zziW6wjRoWU6u22fX3GlQla6MTQj910GAphoNU
x2bBGIQq1KxA0uiJeBcKPrBWuqwepP0euCg9PAV8luSSN7Na5VLSEs24B7DRt0dtxYXv2l49MihX
MyNi95eRdV5MjFQMfxWM+YA+TlqJeu2CobpBaEYfPhRoestxpv+/HTXhQb6mZjqZ/C4kqtY3e8ul
UbdOFm2GjSag+IYchENWMC6YyiOI3OlIkEZ5z7KWqlPIRu21EYR+1ZaaTWV77LuDdHvjNEJACVrc
2bJLWjti35sME6rRVsWza8yxG7fn2rDIg8+ioCYnMh/Me204439LWC+qKokddQU0ZL3rE3ITEXfW
xi6/BWP7eKckTR/6hAYqITtuHGjypKXED+YNMjzO8/SqsAneExYbg8X0G8CK6DgseU2pVizHiz67
SuIsZ/giGhXSg4mNyeAzvCYMzmh3+CZbReJlw5RFKY7GTum0zco66o1ICQzvrySsC1dj1No8j9LD
2zqh4J0MH1hl+9SrQvpVkl2kigKVBmMui1Y0lR5KO4Pi/fTFrLzRb5KqIyaifHtsA3nmfu2YV/EX
7XtB4epZINupl1EcpcrLfYEND9KykhhIlavOTwCzltXBa+TvLZKuOq/kLdSRoY8rdJh0vf/2pzet
wR7zDHvqPZGU5Yo1eJxToWNnQlhTyJKpVeXf6mASPaMkisatdKYYWn5ZMrosyD20POqWC8hiT2tI
iPuCMu/C+sCcVauOJeuQ2XJYcv6jhENVOHX+dn4ppajRl4ZH8/RG9giKgq4CGDrNefaTsg6S81pC
Qj0zSYea+Xbesv+4WpwFcVtRTwZzEvhiuqxrmUo1SjGUzBvyWDm+lhgABEKT2REyecLwUGXpgS7j
JNvryJ5YxzwecrfXBc+n3wP3wwcRCpHmIxYGjlMxEGVxrtNTyomIiFp70WkqpvkggzDVpxC9Wl0E
sJ9pCZTH8gDeqC6XOJ83RqXH1HQ+7NG3vtzaLMCiHbSyFzQcJX5D6YIcRW55RXbvhr0darCHyRCi
1wG15Es1m5gtzYStRKSZqzuPd5O7dMzmE+3oDKK+9fg+z1pu1p9fLR53v9RpBjd/w2ove97YZoAN
fDEuL4J+ia/w5abfLOv9d+b0hTmtq0wvUHDzDQCAFiwLNuyqY4ym21HkzgviCaqbThrmxUWR3l4R
iB6OG3fM+dEyw35SjKRqTZO1SD7MTYY9+uGKUAzxALP9HP9ZTsE/RRkgiT/AzJXBR8MNZpqBdvWK
aHlt8ruBNtBVVoLXuRS8RnWyIMrb1vIEwFuSKELr9gZ3EqlhdEIFOqYpj61O2HNfQthJ1lmb6rku
eNMR2zsn8fwTkk5WqUuYbwLVfTerTPTnFnDZ745jlS8omwO+KrVotxSLwoNs6thBrydJ7L5h8AWh
N2vGHTVULmShLUgJEl0aMH7Adc9Fq5eX5jZUyXoRA5+rePl0VYUJ5FSJolG1BA2x8U225MT7Vz2d
IQVKt2y0DYoYcdaS9d3kwc0ecxv50R+/M7dtAwGzJWx8z6rR/w9mJ9wGfd60npa5vElsqCwGngHx
Ono5UVRU4Cs1kkhpan+3mSrTFkC/GlcYu8EoMMPNI1zKjOGBF2QlIAQ8qWg8ns35V2+gtFBmGtlu
Cncw04ACpxj8NJWdAypIugpaQYxeq8GRJGOxnqYfrxifuw/a/rhlS1OZsK1V3ReqMig55oZMFJBM
4I0At8h1AW++sARkK0DVoiWDwvzPrFnww80jM+SPebulyYRp/GSNbTSLnTCP37HWOyD1P6f1tcwb
q/UR5pebP5dJ1wucxqUy1O1RrjcK3RhjzCsC7/WRYLJbPbMSH3AIGawgFcyJ4wrM9dt/++O6E4zM
PWarWypxpxW1Idt5U2Seto6T0+oyCa7YMgbP9ar+zNvRra+aZJOg7ZF80wzRSVp6tirC8u4AKWHL
fzf9WJffmh2LfMQk3ZpJTI+YkWt3ZunawQgXiYvzi3sb6ExylazS2fl9uhWD6QRb/JgyFyOmkHg4
Hhn5FLs+qp0OqRr0wPmF9pN8xfQiTuRx1L5L9VnbB00YDBCNrwYd7j09p8qGQhcak6hhOprRM2g3
4Na/cPypxsO7gOZ/cDP4nAgWmN+ImpXUf2tZOfFGpiQ7asB9ajCOVYoiz6V6IFYw2RQ2dTj5HLSM
BiBdLdC76TytqLOFO+ALMg/IT5zoogjJyHruSQ45VYXRhVky5mcJQk07Udap3j5qVWnS8JG8Bt0k
pqxvWWdaTr7Pk6Rjvg0h0K3/unpaYnU//5kw53sm0vW0KIpQ9i2gykvFFqT8fO0tLpMwimP+Dver
APf5xbLztifuHW3jasvKThKKMj1mvbMU/OEJ1rtwhRf0zjy/qeFh3yeb5e6Gig1y2I8QiQ/egAlV
fJ8SEljch2P8zvdqcty3U4dc7CVDJS0AQ0xaFhF13v0RIbM0+ykgH8vvm025eJlsjSgKTiyCyEc2
WSiICOyHUGYTA/2PocpSZ93n4so8AJK1IIHQOTBT9BXLc0RwTi/48JKCzC+fdcYrbhhc2hROS11u
jpieWL7vloXF75S05PnCq+CqbxVbqOALk/rLCQ1TPI9f1p5VNbAXhqf0Q7V0nCeKKnHDoTX1IRky
I7z8F/JOvDYWZfX2sey09tsH9F5WctNmB3FD9Y/oclM5BoOOfyrKTRX+IgV5Jc+vd6AG86gYHYEm
gzKIIsMtjb3vcVNsRs3WPmfxREkiGTLd3N8VmqGYzswY9dxtf5X+AvraeIxvzS+TelZKOXP2d6Ea
bKT+LVqKn6Q2XHyEhHP+Q+exzpnHDhwbXNLuTHw195K2bBNhAQO/n/xAcr20BZxWbdsvh/3tUMwL
0I5sATzxFXELI97oAB3ACdMKU3H8zxkpe5aIFOY0+iQk3lLGdjECVGJAc00FD5uxPRfNJfEHGUz8
N2j6xZX+n5ipcJD4O8sWDK0UFng51mVke18gg5uTEv6pKJmvmpWtkkeddm3LLpHOAFCTxH3tkEmt
k3yHG7Y3crCuVS9JXzlKL1VPzWOcDIcMLhx5kiYWXjrI/9jDpHCG47ili4mvSnF7m1kLmO63F0yg
nHkfOlBLBeA1xsj24inFE9IKz90boMHo61lWt1kiz2TL+R7n28IhJWX5mcF1IzLYwLl17O1CCjXn
pnyApaTYEcbOtgL+cCPebZdbhgbK+tlrjx1SkGKAlgoyvEEPCDYwSCZjLpqtUhKOzFdYLtYrmMPH
TpuZ0XaBXpO4w27wtndndORTtleIAeIBrpW8FdyfaFJaniL8nGGWulB1qNufG9Mr0L/7c1Wbo3s5
T0i9OrNVgoe2VgNdvPksMnoOdntMqQN06FhL5sN29ivwtVICF4TKClz1aYrCStONUL/D1W+RT8HK
h4HE7+S9dQ+BcGMNtkDQAp6CWwLkXHSUV/ogNWb+m1dxSprG92Kcdq3azJHFojgMUSH0jt6DtCuY
VrMZoZH8bZHH/ZlzYws3ULsvyN7avDH3FzIwGT7zb5ZrRvg0jSCHCDxXaQyxSoyiTBG6NhLgtkbt
HE6ScregB4AdPlQ3+eAypJLZ2w8N6NM1IUNdBId9meHZZDHE2QEnRHk+f6jDMOlYEQlSKwNiVKBk
xhcscmcpK2jmHCtsKcWcDGKVV4nMECo6UZYgqrUk5HXgFWYBgU/qrubBlk2sUFRGP/yaA15JE7lo
8KZwd9RWB1mgoIKIm/RuXuo/iR+mZ927uzcF6f3aLAjUfMOOf4X003Vgm8bwdZHKURZulp/R5+zT
wmn8M4DhESP+xpMRFBZPH8ObdgOj5P2HQwNfDubOvh4+hPaZ6qiAt8j4KW3Dfnx3RXvns2OX1Jz1
iFO6+T6ajF0mtZSuhA/doyyXwaZKvHsQ3d7ioKT9Mw4/rt9vpE8lysy5Y30ogzj3o3sd4qUyx/3r
JbTEJXdNQJ1bw2NqvInIq1gMuekXjdWG7zOsr7Z87zz51d8+y/a5aY2vBW/8OGlEMGsz9pfjsvWt
Or91cio8P8h+Fl98eS0ABd6xuJ4BZgCWMdbhSmB8bbaUAY3RmX0TdivhTcE2AvIJ+SVo297thhr7
8MG/fkHkBlYctQEm5aRGK9OBwpag3WgLWyBDBGo2JfUB7o9qu0ZvyKyuWJZUYCv2LfeRJ5uNUIqj
27Cg7/BiIGRP+1Pk19Rz4P7UnbZOG6vHw6Un/Y/4hwJxn07v28TzZ8S1Z7g7Ofz8o0S8J07IEw5H
tknpz/TR2Ah8cPwadotnEUW5+ApVyTZQOHzeOwiQUC7SCZIF06vOEUlFFyoF7DgtG0j/kDdjRle9
6r2ms26NYrHDBZ4DMLDxsu0v9IsjfH1SZoNdejtLxuZdHea26gz8UtOm9a0MA/DB6MDBfljwHMSp
eGBSpiL/Hf9yWLk3IX9oyFCyA6iq8j9cjzO3RxASfv+NZFgYlwa7JlXu0Ks5PuKhDsvlyTwFR1Xg
osXpHNyuyfvOrXyhU+kussFP39z8tu1GiAXYnVdHt76txSM1EzxwZuKeIlyrNMT1Z1za0j5ICTWM
J7hS5MnfweCBo5P6Iq9/7GKPDuPHRNMi88YwN9WJ2+BVQ/8wpLCm/MZoZWsrWUFsY37dH8emgFdq
cMNPs1JmaQqs8zDFzyGewuulUliSQEqa2Fv93mtjr0LhZHx1HBPsoZMyDmVezyWsuqOfKJEBKRPy
43bRlkfI+1oauUuhMzeD776CzOorIfjcmnoxI05BqdEbFSOrJkabCObZe48ix95mUkPmUSmp/ySK
v3hURrXTbrYcnRNhtQVHJDBNhPKw08DyaFqW1AZfpaKLck+3Jut2YUMlVlLGQut/kwRxqSf4rdsd
pU9IZwNhNom6wQhCq4hl06B2tRIMoEnT71FNGlu3ES6h81CO0+wKJrVyeS0t5UZy46K0gGsznuVO
pOK4rbBuEZ4/11EMhfzmnieJPfGGAGJueEBqU5ul3IPUYG7WxwYhBbEOAv8G/f5T7UXUylwQK0yO
hdyLRP5L230Vw6QGY1KzMmBToPuykm4xnT5yNI6e+Tf0g70ltl2JHuvSHbsZRBaexDMr39gyVl/1
auSAgO5x/cwLiPC3efsMOAsHNxjcTMU4fEyq9QvgUGqcaKHrxOTUsR/G5JNPfGrqMMmBaB4Aa7ej
uiE9rQUBZv0EK8a7n+DOJhrwwUHa7WkcetUtOwRhhZfaOICFi07XpNUj6F8rzUjtn++6NSFm7iFG
2EWL0Wn3v2UcVRQFBq3CrYsEgRHT4LN1GiS2iJB858yaPFy3n0pq04Zw0kZxi43tYI7aBzsaLP05
EV8h7pnUleDMZ1GiplaSma4QxFND2h3nUv6UOs0oa6/L6tOwUtIMudPcXBGYjCCVkTqZatWzUdVB
Bs5N1l/Ni/JjBrYayTd+2h7uD8g4GUJ1cotasKV959afzwlVdPeJ5WNveT7nsFHvGuhC2fYpURgW
BQqOzyn9gdgCEQvKlL7eBrbJpAz1z2owHBjmsFhqf59W7NVTSqsiHQOeilvV6lCGW5hmmZnYWhX3
NLtNU3sEqv2tw3z07DVFuUpHAeuANK8kPf44NI0PUjSnqggtkhfFSsp9vu8PiGY9Awzxd3mRca6c
iRCWY0AJL28s1firrKKf1X4FA1u18qntUkvhzLrwVPYOwvci+LbdllfhXsP2gW5YUrRiHWhKHZBD
3WF/ve4rpmocULr6SPs7699wrGdh7kUnljjCQM/X+JmP4xncLdP/ys5mx7dit5TCsAan/Ai6FHO8
DY71v9lQBAVd7/dE65glKvlM+TBepXbILD1z8ZzbqxbVCxJPp5IkzC5m1BFEf6chvx7laQ2eejPS
Uoaqmjc/2t5MfKZkzjSUrF+kSC5QEZuaue9uQeBQFXnED/qkWPbJNfGU+9GqZ6S03t4DGe4R2M7F
sfBn/Z0kywAOhBGG3iKPy6e+nJyetwR9UU/K432jXdmNiDCVKbfSGAe1mQgJNqnRdOi+iR8fGopZ
Fzf7wkPgLuzgbPA5d8nAS8+AzvqJ8/g1ZOnqeyv6Iz6BQEirwu27foDMJDmMmAvl7gyElm4ujier
C9hLrb3GqPRasRszdGbP5qIpW+U33hj9WAIO+5BMB5y1BVQgW0yZGhBjxqYwml87nltxwACYw8Yg
l/wEqMS1qhG3GcloZ8LGbp7EwICbwos5Q4G+bdbtKbn6BXkiHxcqGoLeG/hEb88hrPzvjBmCnx9R
SD+KJj1ef56k9gBfarYxqPWd3FuRVwQENQIO/BWH5Wx0rZiMEbsvLF3YJiAddnMH2KJG9pcmTGQY
SO9OPWrERYm1MXkNjYHZgEGoA3Crgnemqa9A6dQ8/tlDk1CT32zyfSYvfT1CD+HompAPoKo9msJK
4Un5CUzz1hHSw0rp8D7/hhF0R/1D71rPMewUY+0O5Kn0jmsdzoRja+gcTOccd1ACDLCcy1ZNkW2d
9eOj+rZyDxF391/0k7g02q9bCEQjB4xyt+gZK/cr6G2UkCgIySSrQefNRbGKpXC3yenJ+eKagLCb
1MRyFnIm+6VOWLRgUxUVAitMjk0uuzfv/rajwshB4iGjEtTEPhhQi9JlnbBY1STRIrjxB49NAbwL
ierdQp+6nQl+DrwcvbAbXdwgYys9rCJKu+Q+1pHSzHRDcu3PDhgNxpp45QZQ2f5zZgkf5iUtcxtE
XG6C8kQpkOC2QaXcxnCX+ZCzgU3Pq0XV0k1NcF8SXQN6i7kWhXGH0Md7ddkR2aANzEImbRhxRHCE
HPDKtwtIsHaRAq7tO/hhHSSiq1qFedIOueWeZM0sJOeXBWM9ucZEpJkYMngNPXh4tgYwMGy9k2iG
tW00HKAv+5EXlr36MqE8gHvhYJ0Fi2TCURVfSkSKAWYCxHxR9aBPSKAjfxqcLj2iv2nZfmWGzJJO
76HITGsMnFmj7C31JwhSK7xTDnKtEMfNULC7hnHN54wcipXQBNFI25zjR14PAEBKKcAdTJ+Pi9TE
VtE7u4Kw2AWWpgoXDN6j57CBdg8ZeKFM2xj3m0rGN55hcqzHtanCNhwgRH2VkrJtqRiE6BJKvyMT
g0pON7CCV0e92ZgSQgMK7u8EFN/zumEiXpiMFkj9qpIz52rKNcHC6mqNUpgJ2ISiwwlOruoGE+CF
XcdPQhuxLvKhf0FAxvVPeInb0j+6WMfiSgqDrkbttr9JcAueDMtXs5fL/XTY8IouIxzss9zZP/ef
SvCwBKSkCjSHKISLKtJ0Q/9ZYUeUTvT0E+QnBA9g8qPHgpYTNPUGQaxvCkEOR0bg30hW8n10Z9VX
UoAN+yUC3nHBKOjhHBEBkX8gztcKdRcGmdLp+jswLVSuGN3MjlFtaQW0rNeyEhWnH5+1zqPj/PJ3
o7gQmHtt/lKjpQPr/h+iW9k2xSazG8RxLF8q+VVvKSZGGXnCuYXUbgroTTkYJtivJEQxdEaX2SWj
Y+cFIAfIsmzoYRUk1fMrvBX/vaEBrsFx/HELzsRTKxqYIByuRwniJroM8c7YpJSapbx0toFIKTVT
1Ja1iVZ6U394zqIb5Yd31lcV4AZyH6PZ5iMkKr3aXhIKslWkDPZSJLPdA/FXX58S5G5dZcVHE3zp
XCdyBPCLH4MjJZGpVgMNRwslNkoL/k0CVg6yxlzkadegpPQMUHHY8PsUy4CXvi9Wgib78COxzDDs
AdSBbwTHcaJ/mCng91+igib/AJqDd/k3aXJT9nXUy39JRFpNHYuA8YOjY876/MgsSqn6VrswrItB
ItsyuXX7NWjyVrenlRGKSU0eitJQN0arElbpKB/TSPf4mICnm4uPpDroSIbZLsOSV4VZElLkrirR
k8LtIn3wJ2bAo7qmxuE50tp06bJup+pS5/Z+36tCiV7Mx+YczHrdFUvsx38HjDxEq7euxpvvlXhO
d+QtvFl7boe+LlSvhS2dc7dtdhJp6AVhuXnGGK40heXyBH50toBwqRiCV3D48oF2bNgabV9qtfUs
QCwKRGfWQWfFi3rhrXJ67/JQgEks++f4eB2y2INVzgEe9uD1wGlAEYYUbyd/eC9TBSC4iuuwmrK4
NZk9fxra64F2eoxAKjxrMjyy0BUApjG2O4cQaXNWhGVeEClbVdk10oaWDn+pX0Fl0UW/Mdt4SswN
yQQW1YeIZJJTtE8JOQ/Hin33L0oStxZyVZkwh/zV1OmqsBYaeEQbUJUEWTa7C6MtzNac4Vta5Hvf
oIlb8BccuY8TEx/FTqHFu4I3v5slgQgDopj2aX3g3n+8tKWzUcO0OCSYvZ4Qh2+q3YZlqJWvKr3H
I5aWFiKHrpBA5H7Xen4ml5RF7I9PO6NimpC42OR2hPi0EVizXH+4ihhBjuvQO2fhIrcymbqbyLwg
+gw1Zfa5Rwq0oupLo6KDBwE1rzoqrie08rbjs3dYcAAA8RpCn4Lw5LmAWh41UxZX5jlIroIXjZn7
A9+xhadnhkEVPrLwfuLRreVbaJ415EH64eAeBPTEzLy0gsJzBUtvMBLpBuZINktoF+HHAoUFCHqd
ANBGAMc/uplIhnSzo6rV4tYxopRqVrZINWj/jNC3yODnTbjELm6tZECsSSWAjwLSh1uhY+qKZagw
QrXpT0c448dk2QlgyBrkrLLMemElnIEShru9UKl0AkrVh24eiNU2e//BDw46yd/leT81dFlSf2cp
IY8r+5+JzTtx3qnOi5tA0AQVe5l2VcIe4rcutgiaFbJaF1VqN74SgzjTVoG8MxI6oP6L60J4+CjF
KG+j7VR8kL50nKr387TWixXy3diqDCK+6set2TcAYVXZ/Nc05vlBUlduOcXRromQsfTRJM5t6bzg
TB1JqAdWTZGSbHXaEZr1i1Q9+WuR7OJ482JJPsNZObkkYNtEXaIEJuDf/nAS44ZLTELCRT5nAq4v
28xjW01MVKY3WbkF1/WziImbQAtp5m+sfQj6ccTpyVPe2tHUXsq0NrjgUKvbT1THtmBKjanqV39l
H5FpvXBFnQ0Ry4F3srMqjD9GYY95shMaVXFeQ/gb6lwYovxO/+sz92xE0VJJ3aLFN2y8Gfm3ATgG
lILBnBz9nKjK6H+Z1Tvmnw5a0aYzdO9PSjN5FdVwD1hk4HNBgOwHTkrJaEE9y4d92DN+h+TnOllw
MhZhPdA6eza6zwjVNsVjF+z5Ho+Ois+8XUa9jUzJXv/ewC1SlnZeF/uD7aZZJqPUSqCl6JNF4BpR
ahA9z/ZQd5kDJVzfS4Icbf1dXF6/ws2x+YKU1XHKIWP+C2CzpFgUzejHqdbLT+9yTxtlaVRqk2Cn
ZuX71fw0mK5k12DVHKloQf0YHRVui2tpG7M2doNkojV0R1luoBelw7tRf5LZLpLC8O0rVD1JRPv3
Ixa8hhRBox6F7rVI6ER0MqrabU+nQIqQ6kCu8MNdBw4nrtNaT1TiJq30xoCPw9EWE78P3enRlhYE
Eq2sYyIetj9lKfXXDdjYJlaHabd2oUO7XAn/EKOhHR6wAALZ/bw93v1Uiq5afEO4IyzGtgjrOsdL
sZxwoq0uXICItmEs97aoYeJqMXy+eik3qRKLhEMo5bvO3V7ODxXRgH9FBjMDo7DHkymU4q1PcqNE
lZ2dFxNhgmkr5LzTUvx7tbZ7BCneC2sKFoMjtJiF8wfNUKiZcNRQv+8Rf+KqZzJTqcPwBth6ObCC
CcIvYG3T5LiCQ6tYwXjZiG835z/kE+A9nwlS6RAIRf1pBoXfeuQMNCAjZCRLv23LNsHfqANY1KJA
XHoShFTAFiVxVaijYpytmi9pkp6ARJFRSU34d3TC1MwZ194VKl9am87LmWUhD05AYAMzip6IgdFZ
agso/74gmchfCZTpreFK49qWH47xTGyNE9AfQDD/JRs+VV6BLfMF3m6o6Fn36mIiO75n+aMYc5Fm
/wHTJppO2625Gqghk8DT7R0Pk/DDVGWjjN7UG514Owx++mWtAXJEFFyuLFurCyDtE/jMvnERMixH
xWA9GZIag2/ac0CSLX4wqn46iJ3ubRyFZJfLi30HiwERWqxzRIySJ7q7Qgei0V+epkGXsnYRyk0J
f+7DVzWWD4pyJePqwWIFHvJa8onVapUknB+LageVIRAT9Q7XQjk0iZNrugQ0A9fdpRoDHgb55g25
oWPs5sqSpOebRC5P5ho3iNYsslCYO/Augl+YqaoX2Dkd/swf+fcGCi0lMb1fu38M5+4rY8GMLc3H
LkrujvfnyKzM1tv1XapZ5XSPYftAToVzipbQcVRfVo0WR4N72E7BWiYiCr01OY5WyHJXQCTVV1Tn
uwJeLe4nHrzHOyw+FCAVSZvTPFjyvTzQYE2LeQUEHKChyWWHw//q1IwI3WWWYkwmJWADKuD4Hlgc
Vc5MDEIqqrMX0HXNg575jGv+qBgDMvzU5pYBrpRgm//k215HHevwoQXLod9h6LI2FalwLx4/k4h8
cmjUiF/rf02563xiKaZ0t5EDXrk2VzZpLJNpRi2i3ltk79UWgIkPtdu+TCsszHN0lvVg3ZgWvSdL
iXGi89jX/H55l7KyEcQT9SXk3SFzWvu5T9RLdmUSPI3xUq2mFAnS7b1E7TG4X5+WV+QOnudviyl1
GYiV/Fyah3EuPU9LODpq76164tHWuXH2KaVe3Uci9AkjsaDpcCu1R5OdkHYRrw+GddSB15bkRoNg
M6YcH3tJNni9MPWyg1J2LlelwbtXZIdpFqfJPaWEUcSmzVpe7QKzqIyEDR9I7C+JqpdXgNZtGbQo
GuEYdmG545qfQXmH90zSX5G2rPVb+qqEydlYttJwYQyJTrsumOLXTTvplDbK6hSR3UHgh7I/ly+m
gXT2lefH2TeI/2P1CyXQIGMfiALQS61uUlhZ2Gsb6w7GvPAGNRDTBkORU5cPjlmwKDuHlds9KBV/
rKdBLRfdQI4VZx3Tz+TKlcS8htAcku4ehT6dTr28OhAaWQ8Ol86ebo6N8VWwzGSJR/Q6mRTmN9+y
8pr0HdjPiljwtaW8JUYERtEHrqGgnfSjVQ5N/meHwr2eeL2hc6yjNsUFIB0yI7ZYywrSP5wKvoGz
raUmqafykIeKt14V12mv0OIJJmgo47hDjgAIrC3ivCAcalyasEACTqVIEnNbyD1GQ4auQrBSZsC2
fIQOQPMCmPlwwUtzXekMt0/Rfd1IPOZevcqx6dQmvU/6K5uzj7X6BBPEX4IxPUZ9N2LsIU+n3GBS
2cHi/DZfp9qZnGmCfj2ghJdzcq9ejiG2irv7ec2h7/a11BbSx/hJh8eWP8MeV5mXaOqGaA+l7/sE
jaA/W8kYdhgZvNvUVmX4M85zWEDCoVqBfKpsTyfK3QnLIoLN3vHpnMBqgX6qNnWgV5VdHX+figY4
DtoOwqY7ob2bWYH+qRCJD42l0UuULy6kJQKQ6X531ikilya1lMcPFtZAKEVouV4P8e3z5fvc+xhH
Ts69BLWPp/9sVk5NCCCF4n1BZ+qKKvsWQWBKpJTeSZa+J/PTeTdZ7sJOaZ7wjfcEuRW5q6YypVCm
dHxJHlCF+mQ9hU4ZpEBiBJOr2ainNN3eZIjGiY9G5lNdQBeqiT+O9T1wV8xhSsvxs8+H4DSYz6ym
J2XpGpCgpwuhjorUUVzKLAsvkmhW27jc2gwImxdWl2lilADYBtPNpHNLQF0gzioABApk5kgyJ5gS
09W3eZ3IuRDnq88ZS878u43wkG4arihc5NN/vgWaCDmi/FHfck5q52raxr/xGfDOcsiRH/yYEUDE
0TFUD1waFBzCyDD372H6KQugsHA8Aw7LVB6S6EY6elgJ7xmD9hKs/DXAhOpZJTD28X6WiIOu4Igm
FgicAwjyxtLr2Gzyh6XSfrw+bPSm7nlfDyiF7MSbQXjbXf2SbyHZDVZvGwt6rWQ8FVPFMRUBJLei
KRmccaLvj6ICvvzXemTpAS/vrHQKWr32BN8EMmvSHoDPkMbWfUD9qWNE45JX00MDD/Yo/7Vdonn6
gg8X2hkaIPE3j2z1cJo1UgyUzeeeqgajRAqyctkgwD5B0O5eEhznfC2KbOUcvkB5pAcCvCH8ZnlO
9UnjJ8k/XE8aFUijRqHAVtBJZ4/598Huja04/A5klEoCHWHGjkf58GY/WQlQapmsSlNRlZ3qMJfG
7XL5eqayIszig+prqIZoQIK0/FQCmRaqWEJ/UkIjlEP8e8Dk+iHyqOoN0DsERCdRWsf9yYcBpVKZ
M8n+5RcKjkK7PIOe2u6y6QYgCVe97U4VMTRLFuIUOijjnee2zmsCAuQNUVreQlN/TBMfIVF/0gBE
fTv/1ifxNUekTsc90hevzMXI6bCgqKUvTVhFymRKAPszf0+hUOBze90etKoekD/jWdFtjC+bGKuQ
3FCMmJCr4AmfHBno/gqJZGJHmLQ/9tDZdtAVFBElG5UkP6tFEmjdfIFUHY/pV4WU2xj53KaB/ScY
z9YoaBjwC5hN2twMAc5G6WviRaVEvFf39B4jHI6zuS3IIA3v993AyvvBUhXefswNCyd8+D74R15z
1d3h7ePLDCpStd7S/fl4QnVWfIQslVIBlz3WYPbFw5WBEt2m1U7/BmlPyP9yfp278Bn5eTUkbdYi
WpcSorD7gXgbAhezhspTmaJZoUIFRP8LfBfKkouNyaMUsGuBrrfJHnEl4hLqSnZO0Hl/M4VsT7Qm
IChRfUHIRAKtUALuGVaH1AtFv12FKUP2gaEXRKibYcs+oFOagyHDOavlbwL6e3U8TVVWWq0ZTsn+
rorUOu9HZaaG4jRsq28J7YVB1g/I2ao2EqLBjNyN8ke5LCPRie9hGKFKWPgw+y1mNGgCVXgxr2Pg
3e7Ywg+Gvd2huJcX7B7p4a/oolMTDZiU11c0pi0P2LAzNjFQR4XRPDFEabFXr2t6EW8HNTDRDo/4
ne0tBUQKIQTJ8laKCpA6jGdAfdS9rxwQrCps0fsV9Yqa0VdaufgMMstPAWD1EMOKAFLqiyQGr17O
DgA93ZiT2167NM54TGJOpcw8cDrcoTwFvTV+0c4OtiVE1Z+YcbsEwD/Zv4LRE+kKYz8SUClfWLWC
ljZ+3nqzMZRGKnDyzuocT0EnLHsJ0Qq8LbxqmMo9fraUEKlG1kPyMLxMGK4FVGTjpLw+g0ysVSce
qsXDmYlSpR/CO11eIqbuKtmKEnh/w4hk+wVBP4K8rLf4iIdiQHzDDuLAXg8q0ZDb1ZhshsSamY8P
AzGtPBvP5p8Qujp7xDVtMVmXvrhW3/RYz54MeOwRrS0kQmApg+BXSZSDyifpR8DZr8ZW5vXQDTfK
FsIa++Wo2aqQ/aS+l96vQ52j5+aXKRSH8vtRMRWoaC9hDoaeupfQnmgynDnkGXx5boCu7Fn2+KLv
zbMm2c8uy7cBvQ3wSsfIR32uaYuLytyZL7I46Zi9J3y+BLxgaW2hwL4w1F1INHBupEJLkDv36uO0
G7yn1EKItC5W5d2I2ioSSjrIJ4aJmdUlZepVx3217bBVdduuIMOeAJ9KPyBj24bAHqbRi/lRbn0k
5oxvdfVIQ2OjK3hPgU0a1/hZCvN5auTp/ONDE7Pk+Os0THJ3hNlS5TRWO8Jn5/RlJOox1kg5smdK
wogja4jpvSSPCWf2qfGpYi5z7K4yoqUrKnGZYvVwjQ2WqYvtojSB+tlw/RCUdztSGiBvC/W9+JhK
ZNRfrnkwj+MJQs5eUxDID4vOHL9/dypyAg7V6NQ+eN43JnYhas9YHC4uWoLhcviJXWlaGQmn6fA8
qLqN2qbaTdbs3lbAnJ4Kcq89dag95rx+nSCiHirAJKOksV6ToWisfZ440xdnnFmpn+vUuuFK8nJH
Osu43c/m6fj378uebcnYLzdFi9qQhdwkuHoZIbC9zBrI80Fcei4fUgh1DJIwJ/AOKxYfG/mIYmDf
8ADDQ4nB9s/7eL7h61/pkEnWzgGYf83pzafAneYL+JbqmHYFfnuSsKLpy57P0iad6ixYa8oXSm9f
x0ZOuegrjMv+t9tqM/daq+hjXj70wSVUf4dNcgPq+o93oxXVx6vhADPcpQ7m3nLfmKkdNu/cnAWW
qSzind/+M2Ho5ylA6/ESq/i4Ykv+0yxde5OUuiu1jKC6LyRkco1iSWfLKxwNaTuAHYal0cPuJhq+
znZSVZXuo+MXEofwOtwnCKEm168HEUsCwWwjQ/XjpHIOhj4hmqceZ52wJODV6MKuRWi0OFe5e2bF
i2t1iAO7UtRUcDoCFcb1MzWHayuSEvTX4PJp1L/AjXwgaQI+1rVJ8KcqLvyDs9iAOMEFUIcT6SeV
4bAGSp0OInXpdqm3+TtYifwY6hqTR3ugXYdG+HH/hk1Lv5qFO92CQ3qOBgmmJJ6c7O6oypVbdm7W
6KjlBheK0WoXhrJTI2LTlRQx/1JHvSIspsy5Al7udRnD3o/0qVUvi3yRD6zwYnQRtU77R4Md14v/
3VmQ+z5rCQHqTdc58APPI51qa+Dz7AlVAtstWGqO6HdHYUCUxsX8dYoyLmhBMQj4dSku9MUT0hgk
Vk59XQZhD4TnmTtKnaOKujUI//0p9V4UFjZ9N2d8dYLkA4Y7TafViC/RxWdHjgdOaqlBgl3TVsaz
oeV3dYzh6QCk27xHYP8i94JeWRWD30Hr4vsUzwSLDkyDV3rdSQ7+I4LTc/4dm9J1eJUJU+Dje/8c
a8hCjvUZgfczAI8q4ktRN8G6cfqT30aAgTIZLXU7B8ij+xyqY8xsi3+rvAWsDAtoy59OnRHtDrU+
rGd/SJ4NGprBZuiJBFm4RSgtFPc/Abk5C9TVk5AB+6dyIcQSDcZLWPCoB7ifqLdh8nhKk92gk887
vvCauWbNGteDcmW8gqFFLlUqUpnYrocIbhXptQhlh0xMDepSQMYuBgqOg+qJgRpCkfi4sP+ZcT2E
rIFyeRYLQoBczkqQt2KbscLEOeEyBfZAkMt65lepEodlr4MCbNLX8C9XIW1ruRftebYTSQZsHKhe
M8VPsRXuWYhYEDZ2c/LrQ/cjlI2j9hTKfxmEsRm71NXuwqiCmAyFt3Ut8iLCwgPMawDd8w8mdLkQ
JULvsFie26supT1pncsucXFtGnZdWmE1N1+/WvNgCeCfOLTTLj4CcYZJ5re2BW5aYKg0S82oYXIK
DEyc/BzzYmNMkxq6iZUA23yRGVz2sc2p+CzDHOdai8KNlLuLznvnHTOVvTH9kTHpQhu2FStWZM4r
B8shjin4Ii92Y+1FUbgZIAv+Pid5cguyQtss4tHwCPY0POhy8+vHAZBVoOYHGPIAuyD2vg3dsFiA
IpUGc9FUGUcGdOcnKG68pS5nBmMB9+C5thPZ7NaYOpIkrGMnJAQZ5M3hpgatiQBU1sqONfqqIdbB
wjCZmEEVk+LfaArxEtsbgzFHfvl+ohfWzwFylcIadlbveV36KRlOyJ1S0dFgLDtDgpXOvV0fk9Cq
28qQT0A/V9L2hsMMHChriXvGDmr7LMJacEJgTAC0JU+KQKpPpzyBmTPjn845NDvaTt71b6R3AS44
ZgohcsiKbNMF6afdnlCZxyoVekJ3W7dxiCdO7wRqClsFB9l9u4eCRLkqGZ0bCSSDgOmSYCfTOi2k
NrkQvrmriw8S26ILqFPgCZVNUqsmlkUVGgakN7wAGh/6OF53uZqw120h4y7Z5taP7cgnnb85HB4d
HNc/A1ic45/capiUMvF+vBhDRRngCAyv3im0bSEDiSHY697TFzF214bOSwReX4pXgb7A9MffqQuT
KstZFXiJVo5s9btpPSsRveh8/jiiXa2CCaXdIzgyzVfqJHD2rrxfSq5SMB46xv/vsjpkJnggac/d
IFi7RtksJN1IESB8fV6xVduulszxhJl7HozhONaVBbPKzP3FnDSp2QCRFFXYxAOdti0jCwMgTn2m
MKC5Z19f493dGH5c9PPhF44Tx+lzz5mP8GOpIHxpmraShx49JE6zx3VV2oYqoBfY2rxSMPgULNJG
tMf7yH7onBJnNnWPCS86klZq1s/lhf9v9xQ93LQKq2eC7O9DPENdR+HAAhvlmvBY6VqzrN3dHw3f
TjVPG4lwQ8ynKUFO9CV44qF+zBgbJIwOzPuieJXdbWVY+uxZoGoLV8AHvaHTFcynCqJZ4sBakfHY
i5hUwx8kwBPd4vyqiKHQrjQb7HsDJ67sbX1G4KjyCMI7AmCLA3O6E5X2M+ywLHU1JLbTpyEGJrHd
HbJAWbnpU9WzdM0J8cjt+PwdcMo+XjSDRF0PwRdkZaSnYizI/dEBPx87R1WBbPibnnjmYdXJnZRH
dIDPKl+uWWyCvRCHH0kWgsAcIsHicGNRBmSKt1/FxK1qHj4eYXj1GTtqNJNYFCm3navRdSSz0SDa
H9To1n2ItOXOEIUiLfLFvKnnE1crzKcetZgPJX9e77kYtAWf+FMzqujpGksnj2U8tpO8Kl/ND304
O9z43aKYGPqnQNk4AoygVPMTpxbcUiQ8ul4mYbcocIUPpyY4DxsrxiEcyFBenPwTX6BTGonKLc+o
NjVKFR14v2+yfSpi+JW6UDF7ja/snS1qN2irIElXFdezHO3I2XtRLUPg2qhJEZaTJymJmaUodneE
PZP1SZohJz89Iyo/GNJCYJSmS9n+RogqbSBWFLWBFZyea2e8Tn9k2IUg77MVDWzhJjylumW6Wa8Q
Itxa+m2Er2B4m5dzjNWfeXpZZOTHIMsWUX7I8KOEzNk1Qm820iBSGtZoxEtNLz7re9NXCoi/pV19
W3whc6CNZycEjeHtws1/9y1X3fbg1a9/K7hs3jCwoIdJ0K8C9gYaHw3klO7zug1yDq37MkvdeLRc
q1N5gIAUlb3JFPLiCBrHkHc+/2c24OBOWEFc+7RyKoZvuol8yOHBo4PNEEZyVmBZSvVGAXpR+ATW
orT7fswpT9UmD37jaIlEuuwDErJ08mmq7dwEfIF72xZNkjUmhjwLXfm6ayn2ee9rhy3CbrPmQIOR
DRSHO3xeILnfsW/dj0FU5TENhy7PLduDCWXfg+9En8/BsYFIL4ruf9BXsodfjatJKDjGYFRaLd+B
gM004Cnr6kFidO2jDX/uVaN03aKF7Yd12hBJhs1SMOpqswUGJju9e/hONxpsQTRHZPPwJS1Ccrv4
qmELeHaJhTTlQIGgQuobep2Dueba7iP42zoAbNeu5k4f4qyRY0xWvKo6MWVo+ooGsNsQfiKYIXLi
hVw6sXYA/N3TIJgtTuNKY27Q+bHASKsHHk+wx5fN6gkLubNvAO3JmBsTuWnbSinHX1zhDNwrEBw9
EF/YCOCFUI7rw1fy2H9+HOwW3A3yjVhV5MRbNF2tkyM7Gez/+cMBRcNHi+LHBCjVjtYNQtMW88N2
T6JWnvPWB+JvDxKHr2cgJo0R1inxcWfY/bvnL48rtWDbJyC2QFgCviZUQXxQ2A3D74wpkSxJRXeF
A2T47azTj0jtPxUB8MC6J9AcVL2iDXjdIVomDokpikUx3KL57XYgZmvIq8ztZMFvU+pFtFJYNNrF
1zl2RCJvHu8jMQ3mCRmY4h2KZom58FoM8+JpeMBCmdBTSta8Z3FisE04H8OhwRNl5fxi54jQjKJC
r7GLLqqjodSX6fytUTg2X0YjZkvIpFh8buR0Lmei7r1jPOwGAGfdYuHf436wytf8GU1r53f5rr57
xkXvm0kE2q7yw4QISdIc7/D38P0gNxYUTt8oSAuFjBxY5kz4uWz74VI8ZhzT97lKgOd63u8eukqh
G3euGhMAjzxihw6oNRDvKk+1wyg9TcYZ9iXIY6sOPS4wUsxCqLImoisjWroh7ygjYNoRneZgAEN9
nah7bPcepRPeVwQXzHq/cBCqeRxKZLajLBMAwVh7MEkrWwutfvRDgBH+3PVQ7ohYXGqCIYfHlNn2
BXf5SZt99DQqQgup1IdFoHjLMC4dZNACTK0gAvPqYIttXZa0WZ4R2BqibhrVNb0aFhXbK+o2zymW
AsBQ0lbFCuwAO4Od6MqvArBMip2Q98YhEcZdtygrOeQ8fEMp48yI7Fy8UKgx3NGof1xh6NuFTiKg
V5WTCBiO0bo46GPMoUt6peNvbUy7gGq9eDm3wM1FVUMVfcobNigqaekA7NN513EecKKuXDI5WNIV
gxBw+obvjJQMh86bplGqetO8nGPRmrI/NP7twPNzEKcvD9PN49JrW6796VttI3ml2fUTyeFmr5C1
lDqGMkZ9KYc0CPm+7Lyb32OTD3CrbMsEW3ejoLRNw4bo+eWC+pACFrMQJorVnbf1Qfuac3RLiGiv
q0phwVRJLt68POJkbG4iPh0VKYjk5VNgbqy3YwbizKmQURAaqkMksBMP2fAMD8aQwE+jO3d+zQkJ
cl0CL6sPY59hSRrf2HSvSfInvqXKfudFbdfNoTBxIo1SWb5iBwL/t/Rf0rUHAzc/9qUQN3XAGEwi
CU+0XV6rte4yapShK9p35/z3ENlJOeruRdGJ0i1hmGaIXz1NBUqnhBskxyZxNqyzL7/tBdVFbXYh
0oYQ3d1WKnSwedpQvJMVRcrqJvMyRxZiONczHSW0BhzkpRRac2m+t8VTtJ39xxv8zgdVZJ0dfIQn
fK3yaZlHeApEseYtgn5YUyxeeMaBDDESlDgjXCjehB/No537ikFtyasC8oB5PyMCUjESrp5c4DU9
u5EE2ehkqNn9dtFvTXsSAhXP1rP4V7/OsIZJou291nBthv2z+qvhpeOL6ZEBOcM/au32DNdG2oj3
jPz/T9hfI6uLFADYxPT974aWyf4xUrmvQmexdmXLiO48wfmiNtq/z1B2h0FopxWBuaLfaeX+mFRp
57erlfu6Kf50shePTN+oQSGV96OUfTqf1YQxmDMeB4qDEw8f/DynGXTNbK43Ly78jI5ynxYpMZ4R
hg4frN6Im4/DkOKTYwDqnvb3rD5f/ixHvENtCJFqMUkVcjCBpyMPmt3NWK58sA4jdt+DCVCpdMmN
YjkzAkAKgFhupR0TFbc4LwDaNONOGX5n2CkYn0wVFInhNjrYL1Swkl8M1Bp+ns0EtLlzVuEfHMnr
gu7airbPu31O2ckO0DwTv62QKL/MO5zIOUZPqknyNkZsMU0EY4HvfCRRtAFGGMQD9+PrwLjAVMP/
nz1A60zmlA+CDHQ9N52uGBdtQF2tPD2ZjprWLWXPvdGrMf8FqDYodlw1tE5eKO8a6NHtDx4po6M1
A88V585WNcn+qhPn7iU2+pRKqTfBBDvSbYew4m6lUmPPfLqFfR+yl/WsU0qTCc9f1m9qPPyCPbBA
6pP4B++V+PsN/rXfJfNpuxi4vf21OT9dCoEl4VUpjUpRJTUBBwtZ0s93IWS2la7Fv9hllPAHRdX/
ZbYgThKTNU9QcGmwcc1IzAnN0bWfDuMag7cTYcvmSjPVEz/jd8fG6IjCxVKFyRNvJhja9onn9YCb
gujZS1iS5ay2PdYSmdwEhV4NICUk2l1pBqi4tnpNSDNFNCE8sQQVuy2V75oENIhKB32ccxXCr/yM
ZbI4YO4rA7snw9Ce85OBKxuzBMimcy+hwtzKPz6fVTKH/AIc/HQe06lWx0hnkWT8RLoaH/Culhn+
1lzgjXKrxeVIOIc6BgkIC4dlQPXsqPbeHXBJRCFDFpgglyLbzPCU2aEJGN6cwGRKjZD9XRykuDmF
Yycb6sEXTKChkvT+3MPNbxw9mUo/KL44ybegu/kKUwX6GA1I/dvnydVB96NtYut6SEfXGz10F/vU
LL7hK6LKjLStTi0XgWsymYYM372fjQn8K2xY1C9gow3Ugh4Xy8sTc2cvmXXHQVlKgX4gJQ/kf5iL
dTzNPktkcVkk809zEDDTk2OHk/4XCXUSpjgTZhE0lNTDKu6tZWLREwAmI9wBDWkHb1u/jwQIct1j
9OkCahuY72luvsGulOm+HbAovVonE67zDT+hz+35xTtL1EeVUdrfiHKKJeEv+k+am0+zijwR3oCt
vTdswSvB+sjwD1Mw93qQt6unqCvZlC+W/Vsl0/K4HfhmOw++C3agVJPw4SFgjuZj35wWVmj1qvI3
utcKsBaMx1xWzSsaY/PAtkMfQR4B6qJ318SuLQS8wUI8bPvOXvqTRUhvtIiZgTbt8lbBOyfArUNL
PfrLZXOHQMPlfpcNgUR/rRhB5eyb35GcSWsI9TlCVnlN5txLE5i6W5dOvbto99ObepFn7rOIvcWc
NTlVNbvk6oZ/GGHpWBDx+7tgkXEudjBWnnAXgAxCrN3UDmRbhBrt25d1SM0tNM6YvUi5v55lugZ6
o2FMjB8HMTQyH9ohULAy2nPLxT7zKPicVUCXFW0sEWawyVPnntcHOkA3gzS3J63QgtrGE0lcZaNj
AZJUaeEggrOjkMR71erhXslf9NplnFTxnXFWlQimz5R42vhFqEyXkUF4w5ZvtfVuhyyF2BE4qZwi
/0Q2I59eBeVfateuprz/9pP2/a/DAi7DN6LW5e1gsvXUAG1JGesH2YjzFohzlkADiQNpnyoP1kDE
Sr83o2x1Qr8wcmYeCcHQNVPyB6hvgjVG2c7+smw0AI5rRRuWaRiixnWZMmLPAfJHxPE183FdW7Q/
+irNVuagdUGBumvbscOg2KKk7af7Didi5++9aD9HGwe9NvWYF/w4NI/op2pRtiU0c+2xPt8zvPT2
ArNxZmNguvhvhc/Egw8sCZ65fZvMSUMynlbdhgajcTj/v5BXkEMwpzzhIrMnjIVZMGOBvJ5MLkEK
8JLnqKtiljYgPopOjCWRmFv1N4fte9kJsXT5uH06CCpKg72O9Y8qRDhIVn6XxQ52QGuIGqG9qT3P
nU2GJx5EFhIHq8pRFSWKC1MzgIzgV9HH0r7fGZlBF6ACNON5x+O+m8A9R73bDGwbgDDS6Zl8J+/d
tZf2OAWqGz+qywioqOHRr5EHaHvVMPTKx22ZTpZiBjQ/NMKouP99dSprPnOsQDxlh5nM3z6ohDsK
gwHhjKRkUO4vH4pfyRYaDHj9fWvYkikW9tLl6BByb5boOz97PIA1c2Y99d32N8MeJZoXHfR+4vZS
l9Ctl0EWCp65+/RPsTZr8PRXgjqDDilXGsDhjcKliHHnevQKRphXwKshent6JKfjjFRlCAlkBilE
Y/m5W3PhxIPNmIXI9iN9Djf5JCF1e0CB4FVSQqx3w6FHQclgZS5srxdzs1ttqlG+gKgnG3unRUWp
54Symd/PXT4BdvhuGS909KlcSGiEcwVTA40nsfGACJNxnY0xAThDmulj8hw2TFppO8VMhvblvLn7
ZRe3r5+uXFmFb1kIS98ic7prr0ij0PPOZAbzh/4qemVY6VF+YVG0vTzOqY/5rV4ZLKxiXi0wyRph
OUmjmGWxfdzmxLEtsYeb1HdQ2LcClGNIKIK4h+bARGlzzw1hUVgt64b9hKbt+i0S/ikEVrpWkFgQ
q8c8Iti3Tn/w3GRBWv31aDW5svnVADu+ayY0yvA3nAY3u30IDoNDKZMrBdAKMW4o0TguWZOGMkqH
K/BoupFOfQuQtFiP35wGWTDXGmOWvUph5MTvMbCazh4ardYNMhtoEDuGFNqnjfL9dmlUBUf7hfpS
tQ+jWUz8axBtlx7m4ltT0obzTd1qGA98IksCcj4wOe+ZupUjfL+Qm9qIjGdp4WQw7CrNzWDIrZJf
EsputpGFT5BQ6oDKYtY/sBMXlnoRJmR0Z58fcs7OU6BzXrWw3KeK1CCkSxuM1gGp3y1JNpz16TOl
sunVV8wpztcwfmFhKPfaiELhl0SZTWBJOF58erg3Q/HyOBaSFgcJOXPYQd7B3O6uZosZPGAWhzID
tpBaigfhjZh5q3FoHK7pn+ibfiNurGVglEdNrGO4wfqjnED2t6RQogE//Dc4z1HISaWQlhRxjZsy
KJTOOxvxWr7RlaUev5YdJ1i3FoE3AB2ATYq0NX1vAGopG8mHUdOnn9iOqn3SXfS3gxQcJVyYkvZu
VFeY/WffKB03DwpqSFkX6aTV+Qej0rfOIW17Ppzde8obFPpI5PayND2QR+iSNdOG4yKoXfuW9sM6
4I260QVVfJlN3B4B+YqqxCz/9nYsz6IbNpvzv2fqDaGChkqL+nVCNBmU4x074rQQNDvpRisZy+Ju
2VxsyLxUYa4T9/pVnGso8Wz67Fei1gYZwjIvf+FoZQrus6feSAlyUccgWiUWESgWnliFx0JniwKg
+ipcUwze2XrJzcpaU9zlNKXFf+3wNqQefqeoXyfHhK5R4Zp63xXBSc3D07l5Io7vbthBiM2j+0bO
fDfjnZQvY7JB75upnLo6yZdd1R9Z8k6e9hOVwsBYMmBwSOsuaw4op+nLBOhvo6ORh7szCLfziFy1
ydmCKaQtk1bDPD1wf5yjq8DD6OQ3aJAbaISSnqz4J/Nzwq2Z4AX4Vp/4swVxwuCtN6dH+blvdLO9
2dFDYwbc026hmkZ906EN4oRgWpgTHbbjQyy2E5AZ+lCwAGvfu+6qt76r6UhZpwVCae7j5YAC+3Az
RLc64a2r88burjyA1MAvk/ZWxUaL9wutnp+aH1j9+ON9pxpfaiPDA1dB/Q5DOGxtSu8NjQ/UejXn
24pAT3kNGl/4Zg2dGBznF0fXeMKIMVEuCOzGAyR3edbhQIsqnTfFm1KTFKS1qBRvhK172jOfmh/y
QD7vYnrngg2RXi63Uf98aoH+Nq538Ch9AFs/M9zxoB7lKfwhM2F7lNrRxsE9V2nmHbF+dsZmuEEg
Xq9V3zwqCOivTrm9HVAp/2qP3Gdg/+p9SYdMC6mZ52CUXiGA4EzFrGcWOvVqa6ZDZ40znMNjeMAV
Uas4YsorKS46k3PRbDeTw98biXMnwijqHI5ukMqoXGE7QnCwidj5nRIq0jdTaPGWwAXiWMhd9DDN
N8On+K1MTJ40uyohb1OGU0qtWNdNkH+4Rr45e5cBhsLK/fiIM/5EyjIZtiF4Cfic7SOh/pHTIZbc
hIIXK/QslNDWwUhScNbglz2leStT990ATPYbSi3Rh1lz+K3C9RzZJxY0a2jSo1gt1A6UAzzXaeRa
Q91mMo+BQkHJDidew764kBitDZG9LsyYTaO1GI8FMDxisnhbU+2JTpyKA/tt8fRTgMcNJ9NMPUgd
mkh01CmCaoRkgob/obp7FngZ2t3Me85V4GCBBV6r/5SRvFj6+gkquaq44+9sZYcp/JyP/IMltS6J
UUUvqWlRBd7wnLDd0Pk4SQSyxhs9858j/4I6cAaLkn4S/UW2lM3IkS/WSEdvPqDczH0K8+AOiyPo
QWPDQ/S9rXTJ1PiShNApjBDPiFseIrXlN/n7U6j+HdUYAEW6vxR/G66Bb5t9ImQKJQskMPZNopDb
jxk6HELYxSb8tx9KrTrpA0oB9MtNtGlgvK6Wo3fTQdOTJ1J9CX7Kj0utGlN1kgnk5zYNxSeMo4UP
Az+EnBMk3etHeqJFlNJa8vvmAi810Qyv2f2JtjaXm6uMvsQNiklEUzqm/mzHOl+NcNlC2D8tofiC
N8e11kI+iP0GGo0DUt32KL2YH6cIjHRGN4ymi9pbaAjX2ZQqiwyGa122r60pVx0Sl0eZVf7YpQgg
b5bQxuODVqZNVhmIAPvWiuPYo/HdDCr80/Oy1Hf0OHidJ2dlXBvxPrUomdA2iS1HA+k2ByWlJwRQ
8LNMMjyzg3Qsdio6pa5jcs/15x0eNaK4qubN9UhiczPdlpaGC+SrbI1D4Rozi3vVcLxOb93ErMUX
vCFN7CJBAOvqowongS/udCeWyKoP15Wvve2VL7gMwqqqbKH5FrH4AKEMDkFKBlrgkzj6xW+Zn1VL
I3w2vKXqFX29agQeTfKJVJead+6Ib/jY7DWQkbSL99SbzK7dK0ec2RuoirMJLhmN3u/fmtaCWKMF
QYC7BMAopITPMyJGuyp3tCN//MIOX5ikkzcSsypbt5HStO0TbOdFeNwb3vIMdc+PwANzORGEnpeW
HoCXhVykGG7FMN1FlfeRfO7imqW1iY4tz0PJLIpxffdO1r91fq8S/qnwSmwuzUb+vPy6cNExbqJ7
Wdlp+CN1mOF6bCa4AdyW0aBdgAfBcL+lyaiQ2Z7JkvTgVPuSdxHqAStlhP/LUliq4ynPX+nCv2+t
JjACvvnbk8ZbBsJCsFf3rExNrZzrsx4kJ5eB0SO0QOYClo15DOPppnGtouT2FFEPkxMcw5bKZVK1
Sl6M6yVHve2AVVXFUh+xr0U0UQMs2fiLn1WcdXWof/JPD4P4+/REtwO49zoC9/570LO4jSE1qHK/
2hYIRL+Fvn2wtpPWFMlF1M0p4UzxQj4XrUtk4AfNpZnLY0jxrPzB2/2mQeVnrGZj0wwj6IpOXxd+
2iVuQvRLtbBDgjPBe2QwotR6MYOSZCqieuvgqlMUwWZd3x4FikkIeLvk9kC/43S60+Rz0DNKVOUy
+ldX49tKzsVe1Tcq1CN9Bp0y//L7ilh8IbDmxJACFC8OEFAMLf9grwEWbq9nwAuCBURvKu31OpI1
cY4snWQk4tkMq0fvUCGyy4UPPnidZ9TtOqzFPfWdV3g4EqE9HIcL+85A9uvmy/4u4W/jzaksZf52
tkb+/RzdiikaIG7zCRuEkyri0i5cUwdqPdVMvEnKkizE19R1NLRHa2f5h9ePJAcqJLKKrjfUP/BO
/Gt7cz4r1d47N0Hexx7XPk8m08Af+jJU9BzyYA8R4KzXE6zdHqVGO52Qo8Oww1ApvIhepeV2uUjo
xHy8Dvc50LNp5ZEg0SMeJmu30jISrithDDhW03RoXcpgXGTfy2BGoy5byTFvstL1T+qldKHXW5+C
SR50pBab1cACudPPFLaalBcTB8UdqTfxV3iaWsS9BsAZDcelRzM3SH8doaLH+6g+jFWgvb5tnOuz
5UlQeQ1/vxmbezh6ItsHSDD1Vd/T6G+ljcwiqDYZ7nBIx6g+fKw58blY8bhfVhZcADHdvsQKi1K+
hLRoOfkX0JOv8E/fzB8wpTFbbOZyJE+WcWPFvplrgHtMR//3Wy4wfROw7pZ6bH/TFDgar03JbTqc
MW6GRauSY67YGoVLk7Oz8jVcRmwjKC7cIQtkSHsdrT9C6d05IP5rLdxcuxX6EN8neTApINLwTXRI
YHhie1Yz+QHOSanaLONrOiY8n4KEtUs5zKBtrkmm+1/SVfpruDHwIchnVKFSjUFhmBfqpycVsDOs
73NkxucujrUIgNPoG1lt8gVqwyoTbqqU+q1mdHlQyXxKV+mDFxDb/FvH7rUvODCJMBlz1vyxW5nt
ZIh5YEVeduo2YEqUK+aMLmLV0srCb9gwIStp2bfwb1uI0y9XI8FSg7TzQZabczNfFnBaGGsDXNTr
8poHPuoV2hutxJXaqnv39kvnyFEHkHg6dcq/qJaSbHyoMVZuPCrbIF/x4uEUc92jvPV4oMwuDZx5
ouC4CekOzXoDcgmhrZ7KoPlVJoI9QnAR+E+mtmr0VFPmfVMZLEpd2W9TYUSALmBp20y2G8/3j6GY
qKJWnsEYNqBK42CsGO2+T7Tivi0FHsiyXG1qMfUk4CjcbM+OUMLQh+V3BBN9Nw9bV71SlHpFJKQo
kq9x3zBmvX4pMBrZdiAH0Mco9oWt2YqrQjbj6OemEWbXdjIaDz6Y44pauoRZjBMl2ADRZFgdb8Nn
z72dnDCDHdZ7hK4qPUfje9oV7e/fW9kvXse2go7oxOkY4YzN8fFBWgzGOEp5Q7QGRi2buTngl7Ef
euR78B9gAuYf7cf9kZ1qqEOnxtPX6rYOirJvOwKHozSxMtRIn1kTJ2thn4qt4Iv7YzOimaH5hPkr
RFfghNWHVmNRl25OFpyzIHbkWNU79QnCsCsxmPPqwy7RkRHFRoW05vuQm2cL3Db/IOfUQGQrDHIA
TlPTczJEU0c/jRvh2HIlWhODlETLVjJLC6rF74AjaCznZ+3cfIR0Vpf9frVeaVn6iXvAeM5R1VAU
Vw8VfVRWfmud1iwJwaVaJTFJBw32MkiGhek6dsmSJEymJYBBZir+0n2T04LGddmXE4FJbIKWFlRK
Tmd5FGEDoJB1dCjthU7OjYZaTfY5J9hZY46iMBt7tcIhcw7rTWVfdKTS20BPfKupl43PoIkxmCRo
aWuVJshKD7dLOkD5VEKgen7T7Dn40D6no6kKE2cLxT0ZwMx38ktnp2CKYmMDRrQCzgs88FaVZvpK
7P1/9FCznJJ1viNYP1+t4i/tnhQM+RHdfIbsf4MFk9bow4m85xN1RZZMpsvEUoQH+pdcXRGWMf36
jNPF/UIxDWVUSntYO7hS0tq1ln1h98OrwNqoRqqD0MdJegl7Ts9McE650kRuDXwY621gn2EiAosk
abPCssqYtZXimQn/0QReS4QMxF5OypurKXqOTWAOLSLOGg9lN8JAjCJK5NjmPDcxjhnm+uJPO/GM
mIfSHxeDongml7Q2ZzNuziBa7432dQyp1a0k71vxXdJh3WDZSxx7Kp5gRiNfwJ2b51S5y4iT8w0h
KX+fHfTEvaggl2ScLWCDCQh//pwMa+Axw+6x5McHsNzk3YoUvKmYne2WWOoXbbRvoCnNdbtNQdhf
/Dd+YQjuxIPEgLFdHIX2vPr3/t90RGJfRoQ2jNcM6Jw6LadUqI5+PSPpi/3ANJMbLBEKxv/ALjrC
Yl1JeLTkX/x5FmPiNPKltl8tWXRKYptv0wvoUIWLO9uM2RQMQX5smYEJwWada18jMux1NdLPb0o5
RINTMBGFpyPmlzwg/oiRViJ5Q5y18uDN3uSYxGHDVzWIMZhe0/ULis3jVu9KzSehaPxz0ACL0qAI
3dR9IT0SRiyqQP75oF7bkyf2/CUlmazqUDvtRyODN014eSkD94w1ujk/r6wHPAF12PE9SRa9r2Dq
5Xj5S+aaqIg/XxvaMM+DOVxCwFbDPuhYnpwcd7J1SyOsoiodS9ag3YZtGu9X/ZQ9VgXp/A4bC+tq
3WnJshMVrkgEJN+v54wpZKojLebhnwZUa8pI7GC1H7RYdVLqXCIxxkpkRwg2lGiYdaBGEXOZBiJb
DmQlbNY6uFjpmfDUhh1GmRtrqfPCwD6kmCNa6Zz5ttHz5rJvPTjMacydn5h8Bx3viU/d6vSie3aG
FKwbbK5mqDJGL2w9yimFny6x9+IsRagXUfFua+4DnXiHaeF5vTrPFzCNsWnQd0IB/YUG1AgTv+Y1
oQGMA31WSTSkncNvibdp8cbNHQh4s2Sg9UfP5rtvS639MzeiivfDuV/hyBk1FhclENQV46YzTq/G
phxnbK4QWvLOt14UF8tCr+z/9FX8pPPzlzUe9TK1P0ahhEyTw6++2U4/lWsAF+85jEal81ZWXxTJ
CidKHucAvdrR63zzu32jC9LViEgkC5ptzANpAc8jagL8CnZN8diDHiytzsw6d4JGOLe92yjIZw8J
gPqjMXDNiq/sw+WvDIAh0YQtF3hPPtGowiYoWcyP58BK/ZANLiiS8v8zW2I2m2gOl3HisDme8gaT
b3o1Rys5zio9EZg3euZgNlzGIlUH0HyF4Bh9RTvNc3p5C3dleCkirx5/Z6B0Ry+IgWXWVPfm+bDL
RETmsT7OTQLcy01S/K1MtCw4CsIkNWrjYbX9xLWhrXe2vsXKAAi53cu+4WbG4cVij3rM59MxQDEN
XrGJT6fyKFWZdF7ZG1+Uxt88nvz67lmNTln/mcoE0ySg1Oss1muF8xBkBlUF8qdPdHzpHXd/mAOa
WivSrdYIapIbOefEVrQIjuVAW5mSBw6KY2XF/O0TnC6ZL/Zz7gw8F6/H2uVDbnwonYDnGQ2k2gGV
xyGH/hyj0HDwg6a4J3ge7WWJPLg266Fev0dUgQTrRBgwHSfmsh0tk58EIL0iCXpAcO9Ode4VLeTj
xmZTLg/vh31zdnGczolUWkXlXsJA+xi9nmCU2qszlTI4kWuy/OGv0iXmqupI02pcjjDYR/tw1/vw
bMPlbWkw1RgOXvNTDjCUiBYUJPNTGIJG1LAYV41YUnE2+CMzMlPib2B/MqRKJ3lMraSWqc1lRrjI
Agrze7f1Psjs0gQY81r8tgKHYsKpzD9svE7K1OWdegx+UqxI8pGUsGf6jmml+rLstYQVcP2+RPxt
/lgyXhufqLG5YXkVvzXXWdVO2CqN7sJQfjejEfjd62n5nL4AOxqHkaAfw55fUd9r7IhCyRfx5AZ6
PlJmHGbA877l4v+RLBCi2BaXQneRSR533OE9XdnDWw7NfMMU/3fYmSnMklbxka+fw4GEIQ/NCvOx
VmR3+ur4dZ+81Hw6miSDLgvUMf16IC0TXUpwlafA7mdSHMvxJD0yEV10req+12xFPKExhhZ6NQVI
WZnWayTQ0SMWF1WZDiqXfxDR2QLwM2Q/cZldNliR2+yrP9AWMQc+T0jwWmsFe4CgrCF0MQ9LaYIQ
5cXazNojdc871HSZRPLfgXfWLOPkr3FSYQfJJv9nWz0FuhxGn7HcIGoDAI37CijeSkvJgQtLNppr
G6zqnjw5WvBHKuAbL71tZY5ORriHqiXKnwJukioA2W4msQllVzFkoe1cqaeuBXg5vSZcjopS3/wR
J3vqMfTz9dAnJlqOpu5fU+lZM8p1S5Jn9NMY82G7j6WLxBh0f9qXPjiO7qnSEVaklaU9Gpr09V6c
Z1O8fZ7R5jV+cwmJFMXV/Kh35VxD9m8NXpZnPnekisA173xAKHFm+MPlXLxcftCN+mCKV23IQzDi
oSDhMlWLh91MJbp1iWtnKE4g11H1Y8DqoDIy7Lp9o5Wu4U8JL8E9MOPwuwKBGXDSvGo/8R+6thYC
cIUB7j9QbIK77UYyH6dATDUBhykTyLDkt4f4QrrY+elB/RPKms2EDTNaJvzUiRWET/kSNRL3XQc0
YhpQWxDMWx3TWGyMQkUcgv9UFGAplJedzIPRRQGlFU+pDcHBsm6B05eBQVNUzQUBJwofSbKIHy5l
7D9ThqvJtGjpdJ/xj2SaUcEoD2IzHlEkffmijA3aGmo1HsUclZNPxXpgFoeLCQaUdgxXJ3Ak4zqO
weRzdBCJ3wqhBq1+4JpmweaVPYbQ+p5Y1Zo+VeSIbxAIUxluGhSHnMMzX6ee0roVWOFxaTUfMwxQ
3MgK2eOLIu1PaDGBsm18iulGHK/Yus3QajHLMSbGydxKbhFRNTx1P6hoiQ9GwvH+Zpv7osXguoM7
qmQtqggAMNmiTIlTo0m+FqVRB5hq7GTXgB6csAm4XtBTkZzZFxK8I0eepBKiDvyfdggPODKhDQ/a
aTbKvlkBMv1+e7o42wJF5OQ+T+UNx4dhsKL9OKU4l3bz/SwlU5lzzyuE+aU0A8Gts2dowINHIzXx
6VnhSG1uFMgcGuW3vV6M7vjMw2aIke0oDb4BM0s5fPNFYIyJXigDwoKe7M9P0Ihk86bF5zP2hZWI
Ap0CE4vIOKgUP/JbUCkozBcZIJ+VzjRXdlEQl7vjLuEtQMZCNKdsSbV9hvDwiVmCzBi/nGlgfdeO
mmu6ey7zp6lmh6d7b+82pweMrOZatwPgOxfB+0ex7qHIYkMy9BR8k+2i5xdolZC9MtLtESPnjb4W
DOMSykpyTHAaLZ6xrt/EBKBWSANuV/0ZaWxm1cdhPY457LM1LNwv50Pbc3iaIj01yf4y/WK1vyZV
IyIZCjYgPrgnk26aVAMnq1aB7QY9pWQt01tixdz8G8kbTvaw5iGXBVwdz9gY32rcl5A7lgVb1aGd
ivUTr83LGzX8zGS/qk9+Bw67NllBV6CJw7ju6kR+Cb1bPlv64lg8yIFh5yjhNGBLObqVpJoOTfjP
DLQ4Jig4hrNxjt/wxhkmyH7q4DC8w419E4I/MRKOlkYUvAwCSZsTbLmjdW7HnyBXPOeKPUcgBcgG
Tj19TfWj+1CzSGFMReUFD3HQGCb/PWjMxjPI420Q12P1gXUG1zLMSEuqWXdjoRJJ9+3U2ZBy2VSA
yc3fY0m5J3YFW/9cawljYGZc6sn8+5MHf8TLBZQvNP93Hf+CWQ+PWmSY5IYhE0ww7Q8e0jza1suQ
O56iaUj5kEK7u0hh5ZaL5GxAZ3hh6EwGzXKDQnk6UXZ3sfRP+r+4Kq6osCPEXnXdMZ/ysBbSzzjr
IjeDGxB8+Sk0yfN3Y7ACnFs4giofdKahZrj7eAyvVZnUsbnGuENikk9FuYwl3Wd3a7Hsm8uo8bat
sih8ax9DHulXZ+aqtzLSoMfrfGlZDPBr+Ojc03ThlgeBt4WgENYU49AWbKARhat+YGpkX2raBR0G
xsZ1+6xCEjNi6xqQYmdaRlHx26aQcwsLfkbLtTV93vWyv5qvObG2nihv14/OwMzNYDLzoHl/HXdJ
XMOefld9yMRu/jalmtBWSRVbaWiyvuU5MQ57tKSgKXy5g011YDaweJS1P6zbLfSvNUHt9plQObGZ
kc2/bvcof5/8xWs5BRFxJVm4oTxQMiRcmDnAuxvwIvNcB34ux9PHOk+mQGDpmNeWGxULv6hqF9l5
lMG26iL2dVdUKFDmFVnRs+mimfS/+uGTQ9bzv2F7gGj+XCGgGjQv4qhmfUbaqMV7IB9TH0cN5ddo
IvqIeG1cUidaakXCMrptlvFHFhM/SON3S7b79P/mJqywr9SXOED7BfEwbyo6etn8sJJauENYWwga
7+KdYQMLdTEJITHMQ/KUh9DPr0/liPPlEMR8Uqj3SRhMMk4V6uP6WUNDoaiQyzLuhwjCgQDBYwTV
zJGGzFgxCcMcTJHPsTItPUn80l15c/+f/toJsiKKIt/PFDQrZG540ZrivfWbF+o0PAEtBZ/EXiVH
P9bF8xWVyrg9VlB32EsdCdXkSeA5uHEDSPsW8qox7R1tAqQ9GdLh+eX71jiislWFN+9IvYn70Wkc
YzaCO4NcQPxM/MxYs7/4hayWXLEuUqK9IDB4Bz40DmYyH8DK5dDCYE0p3vSXoEj6t1KR1vGk19jN
z2/vV2bt28jrPaBfbuj1u5HkysJvFY5YRXV6TtMbvXW2OWkjxl70czwAi58XFjAF8DYUt8nhAFzd
bGe37xh+K5SFcUrmFVjbpNfvuZeRmCl6YbqwPW8y1MoG1wkNItdeCkv4A71kpPTV3lxYkXveFAjl
Yuw29sIF++1hQj7g6g5epKQhQO9eb2Pd0v8bxYNftQjg1Ndlm8LLO+vOmyDKMnuNs7dNeV14Bb0X
TxPLtLl0nHI/41lfH4EVg2LtxJOdC46RWSY1JbHMFMd+vSfQ82SifvPPfLw/oN36bvo7M/Zs1ybF
6of/fgQWrYUVIZKfQ7FyL4xkY8CThtTf4NxcDC8jilMQbSYCfkZYx5FaFejgUMoQ3HmKGW8vAdwX
v6Y3CBG10/Ir4dONlo/hdnD0OD6YCdHu+yz0UzhUCHjcI2ucOtsLo+ixwPe4kAyTYSg4OcCsjoZi
vTaAxDDGblmER3Nd6IszWv0o+YUNhoEtDsq4MKAxacm6xgpL9OSazVv9hjbkRBKbpnedp3HtLAEA
SHFVZYjcHT3STy73UFHDXxZ46FXq+MG8TufK/oO7KOKfj4eian8LL/UsQdsrUhoNiv0AnBKifKex
SIZ/nSmVBceMAmDH/jCm711GDydIG3O4kagXXTV695igxHl49gpt4inejWiBYP7+S49FWW5acy8u
549F1f8yT4AosOUSuY81QcUbWyRNPT/jBOr+olMx9s4Clk5SSli9sFcAKfQm/t37y2t6zJbOx1nU
4ZhoPydryTn+9Fv+BC8tqZyexVwToD6FVOaiaUUL2nlr1M8IPbwd8/YUrCBl23ECUEoyDxC7vFQ1
zArQIYFyeikZlD1/oXfx9wttrVz4/p8jCVWBupoCmxB2eVk9tOuHYeljRN5CXtegAB/9CuVlZWdV
rHIAvu2LCdHbCPf8NcuC8wY87WEVNcuMR8/TxA5hFu+XxdfK9+tWfNkEbTPlavmw1USbpDefH2RJ
638LXMb1fHZ1/nfgHIImlO9a1rANLzqrcgWqgVcmmNOHI+8CWjOB6+xjfLScjVglg6Xw5ViKHnL0
AbrzKPb9wO0+AzC12vWnyQQ23ot5bsiDTsS2v28v3XgSL/kGVIWR9npUBiQ/9b5NHYxUZWCcAOS9
YJgiKJAqdJX9vyyhnuWHosHxMi7wH4xnHfNf9rfyYCrT9aCfiDznokEDwqHcbcExGuQLF2s1glf6
yrfSGZdZRdEEeJFCmE4apK+M3MGzhG2qzUSBVqJI2iIvVIBnGWGUN/tHwgkSdrjU+7qWTZskAqad
KtUQ9JfJWmDM2VhdBAfpBrTf+TgjWV5IIpCnmeGE03j3RayRVUfkH9Dsw1XBT1i87yD9/IWEmxkH
uzPh66oJE0BkqsOZfGC92d9q3bf4QFGXsqvJog3beOoFNWniEbzEu/h1SzPqk/UGfvsehC4AwrOk
+en3V5EfPKJ08PZrpTKc7ZMOJfBhpJJft0tBws104ygiI4ElW3sSjGTNGGc9r9FHQ4Nbyi+ePvAq
MQJNFoqrB3BOAwtYb57iSjHR4mLC1FTERh7KA0iOwrgbJAwyLcxZ2i+xVinqS+9K4qUoMXJwv7ft
VY9jMh4FvJUOaxwWKK5eBzeOFaPrFMhtbcIhbJcaz8eRb179MOhFZusA90ITeWusq4gm6Mq/kfe9
dohiBNn7YQN6fekt4xUQN3XjeCnMhDUdCKexEg5e6/5NbJslA/0A6sWHXjydrcCgJHB5316+Xy1V
AzX8dEtLYiD1YhlWOi8ON+U0IXh05VEAK/f6qYAAX9d9Qq5jjstHWSThh7HLI6QL2HBZ24m2J1lh
2OYl/VwhfTyVaVyta1Y52DRLcCnmXnxNGDGrnd8rvDnz7H7HBCMu0EvaxTlAVmhkn0YbCFc7jQv+
bNm180X9MK8vTZnSQfEZd6foTpCUSJDJowSi1WlM+wlYhIuvlZb/KnHcChJeGk3JrskyIOULPQpU
PsKxHhXhTIDRi92iCmlrUSDPEquWG0BZo2GcjDWKO7raHxFyRZmF3jXkziZeVPLpgy/drDV2OdEp
Q/v57Ex8zlTTXXuOHEgCQSeHpz5FptHDLzHwJOyzNgBAIleQj7JslPTzJb6pjuK424SqK6rJfc2x
h1Q+0jx4zKvwq7kBs5geMJmHSBxiZSe7QsYP8oG8pDoQqQwTVWBJ+Ua9FmPJM9tG+PYnOKV3HUhq
JV27XUBFrA7gACrolNzfPavjZJfa9hAsNmR7GqQbOnkqlcKzvYfr+Ax0WMtJoxdDeHrK2SOANsWD
9NUl5BtXKjRxHmbOz+8uIN0zXYvt9KypiI5neDg9DB2NFHqDSguerdg2IH8/BZxcER4Zrc9JPv0S
uTt9Kry5p0puHOh9IvvNI+v+nDyhxOazE031d82Jsd1ieAxzT8IXi+2Vke+w3sPJGWWshZ6Mpp7v
+oLGFJEnkuTLqOxTBAat65Fvnmd4N7DCfvYBdOGFVBvmeA7odgeKc0XsRl1d/qIZ1HQYZuU+mfpY
RXxHzhrAz85goN4dF4kIjnszwECELlY9jdwqdYbySzWe32ffxCWgg+Lx6wQYhyVqj8CFQOhjUGPr
xaKQ5WIEdHMTOkaVeaDBgTSxEWtLp7c2KS5Dp6obpEfBES5maHmyBTq3g44waogF30iXdaUQGlfM
tX6w68nZXcqtsn+7uIMKm9vMvKU6QXsEhGRyHWB0wK2vbIm11jW+xuEZ8d51JXFlmaG4CaQ6BC8A
lZ0frLfxeObpGODtdW1l1qkNWVRxbDiOwMjos9ZzQsl1gfH1a5grZw/66Kx9vHNEUdTLU8zWOFJo
pTwbU7w8x92lFrWf06fat5XiHZE4mLEth8UCwGzTk5+ZOpxTXVteDi06yi1IOaJdMda3Q19OcPwP
4c3uunB6M8N1nkAah89m5W1Na4o2y7NXGESmcaZK8SPMYWMoQwhZ/crpPZfuACPzdMpFZiJWT02D
GLAQlK94BScPFLZBeoi64B+rkIQUNBTJICzjnHw6NpU/lzjV2xVn1rGEJVjHA8rm8s23k9tRKn1/
jn00CXKMvpBbY8I8pX428QG7FLKZPTSsF6pDi3i7aKrNyNfCJWxYTUHjkpwyIG5IyLRR3TD3l+4y
OZEZvDDVxBbqUFNkC6hqcu2F0sYcjw2Pq9YcgAGzS86sDCZZJrggnB93Lp8+wQhHfq1I/84Py1Wj
9Ya4mWCE/QCc4tvnUyvmZLl7ye/cBu0av6ozuz1gWHW25rMFvfdfr1CrszFO2J7SO6+M5FAJoyIc
R8U5iWLkZmZs+4X5Z0zr1FWUqheYQ4p1ze58FTaJHff2vqJOgBHqM/gi743GGBOyGtxo37x6/MMX
Pfx89/qn/PPO9qL+neH2C8BtiT5JzPNM1xF5JkdDZbhaKu4y20MA1UyLDOoZaNF0lANu2/yFXO/p
iCNYdQrpiKP+k4pwSfDIgYAZLJ3sdw8M1mh5Tn9uCz/LHVTApwDHBr1/Pnx6dU+/II2AYbeoYsxO
ta8ylvAGoLf44RCyGpmGaTHhyBK6JXHJE0f5PH8SU4H8DbfQNKI40qwjhXeIyRISWD4Bd9UXz5cg
6J9jsiwkZJqbrurBXBLlX5sy0i9oIS+sRGNtGl8xcLBb5QYgHsB6xwCFeOGKlB1gfLI2JsPy7/9g
KdxJEdR/wH0oVrWjA+FY0tEKXeKJ4Mp3mK8+l+SdxX3F2sRYMCzBcswA0mLWZiKoTvnFASGri7Ge
fBs3rITLH4itSEvCK7III3t6tZxQwKoS66p6JX3fuTSx1oyOiIwIQjVvFUcJ9nuLYdHfecsn50B4
9//MXZ1SzzcfAkmP/GMeI1S8nCWm/u4xx35AOR04bKGcppt3Pi4LB6iJnka1iZ05HKweZpqNowMf
LeE5DmkAiaMdmHpnrPGRSbz5SZ9CJowiFAjWw9/DsY+FYNEz7IgfWxLk0t3r02zgMBknkJWhoyMV
XnC/HqnJ5n1/3M8+QwMWzsQIUmv2ZMYo+YC0oLA3KJB3hUX/KsE54KdmyMeP/BLbDq270x2pmHnk
6TQgnFSQea3TVbJPXcdhsTB5W1lOR3uB0Ar9jUs7a/KWu4NizP99y9PbEDY3vHywxEr4YUqUUxzW
o7bMjNeQSB/uWRz3Qb7j6Ce6E5HsXuWj6GJzi45A4wWXC2auD6HhUVI5rQupohzwlVuMsXxs4etK
1EnLYh2XsTMuipidkY9+0wjDfQ0UjUvY8iI7FszwlbKrOlA+O1PucVV7d8h3t/KO2vvaByAvZois
VOwU6qnFtRbesBAGKX5IDvdqaCk1ogVaviz7V6hYsn0meliXAP8hhTZAc7PJ7wDY/qSHn31rZ+Xg
UK574ypnPRc/F/WojZDU+EgFcj6DEhCEgwySt++RKWsZU0yRNMHT5s4YdbPG0pwOtHLtlsnBlnx6
n+KE5l+4o9ol+dL0ZvRjeFirc7ssCJ2ZGOO7oguluKRCZiIPJmxqsaHNLgeQyvSsNZjkSqCAt361
flIM1E1CS+kXJldDbNPAaE260ZSsM2s/NsoKR8WKSNAapo9iNz3LdNEo2xVPiibYFK4D7xMutJ2p
QTtIlgilzc1bn3zQ8m7fh+tJCK9iVN7/5DN7PSKXA5EP3GGZ29X4OT/n56T00JvnGIqzHxSs0fWw
kWgpmFMUucbkxXNA0H0EGBvTVziyHJ7qxWNRyIzhiu1DiD+JesoCiJI/uy3MJDtu7gTPRgI0524w
RsM/dpB7D1zKKQp+hJlx2zjtbXhnM9QlR6kF0Ph+dP6YSqmv5Xbcj7zXjtGrd9gEhk9AOqk2m4hB
G4Jha0n6va1t/mXCUVkmHkvawn7WcnnKKB6PJxug7UwjnNG6aas4TRtzZo9/3/JIGP0EdXGqfk85
/ROAljbsyprWHwoiuOZmRDChxQ303ugsMQS2Q4yYMyqTjoeytFqERzPCTy5Kup+SYM6SmXjyJx7T
g6umTbSusrZI3t9ogpe0smNuYh8OI3l0SB/zQPDsbm3TJ9LcYT9mAhYXpemiFFhuueTAn6kWP5UT
dcwOpCyeqS+DZn9L/9ttEj8nPbyT0xBNmftXm1lzJfMphpb2IXS9JM0w+R1lgSON1kUk6NN4ROLA
wb25fNXp6gHYjuySGfXmIz/LDyKyN36itBmu8kjEhYAsuDjkD00IO2YJByLty9lvLjL0AQybVeX7
Pmx0gwHe8Z7Gf83cnwB0HX9H1/c/NU62mRG9J6SeYYznPeQVoVT0KlWFW1UZU+dT+5C+19mD6D8x
UTAyyM6swfEgActW6ANLtJIOFOMQHJPjDw00tXrfXIYzyW/yFw7Il5w8dmGNmIHy/WhmGF7ttdr4
Hw3WHotaZtzfvcOfPtE3+ghoVMG98llbySp+ijIJBHoHjN2P2Bl5VvmYU79x+RsOz32TOOvuRsyN
onQY5A3hOi3wzJawHVdUiPoX06+mkom7aDI4iCwEgw9dTpl1I1dKebZShuli3hyovhtQRaUjLDoS
EUKvYezQvyh40qR+UCvAQ/DCX0vNOHIcuiiRhWNLoDrOpMZvGdaVlaLSa3FvpKCeuKjed3e+EJG1
afgeTrUjDMpW0uCURgFJNy/GxmOfnJ78MjEkH8ruys+SdD+jaYSIULZySwzqh9dHDvv+AKQywB1S
q4trO8EFTXsJJDO31uarrGVkMLqZs9ieetFmWgjTkmAtz+zfCDC3z2tU7wWHhdPwVfrfDi0Dxn6D
O99gLQOiLySnno8QYWd9m4sR2IhNHdZlbCZ4/r9fxp9/3uU7SBQEQasYS5xzuDTN6OlSSPX9w+o0
FPPABq0MH98fcARirqUi+/W8Hi4joJ9DwZE2xRsDpioYLkdSQX1D20APpYq46bC6rcSui7ZFgMXs
RYw8c27W1IqZ5mY9EUKlPc20T8ql9trXLFi0PhyZqM1qmLimAJWKk59YKd6SlX3AM4pPN/F4mrR/
XzSwgn3XCFPNxJ+mYp4lGZFq4pfktkCIfbKZS5+oTAR8S61ThfoWQbrdM7K76AcNir4xFyE1dCh2
6l1EfeSSIZjR/1qTopZ4tockxvAbHy+0ELb3PLfO5fK+GqEgg2J3+SvItOGTTB/c0XCZ1diwZ4px
HMH+lVj+MnKtOPF6cYXAkKnw5ce8VtGo6LAbxxB0eqTKWrr+bG/TsR6/0940Ahzv/EHgrkNNbWVC
C7XvjODHX1qZFXxTSQ+99jIRNllLb0FsLN0kYEb5S4Nb9xL+fe7KsNUVXGG+OEMiDdveCKnIC8oZ
C5Ho0ZEnRWxX4+0e/VPqhj3SF9GDkccrG5PE+GtgIfZQw45kQbMh6xnj5Q/OPWn6igLFiYQwf7sd
EV5x1uckJmKQIh2GZlhTh7EZY6zP0h7AG0ZrcroVbVVIenmMei6X/OpgGPB3GvWteQBLSkMt2VGc
PYEL1tCnla5NaBrFeoBN+xJpnojNXOHhknzGSAWeUP2aepPcuQKk+/J1gVvD8K8D1jLiDWM7v61Z
5s4pkmxj9rKMi8J2O2h9zQvNR/vGSgtAteicCrZZ5WoZvG5mckQPaHH6SzTIcM0e48YEbXyci9rN
//zRme8/1i137ARAOLtCv+kjM5f8YEoIxjRRkDPkkInj0GHjpG0+Hd0g+jVBJsLy7oHBZSEc3ovg
wb0MHPEyAJx86qhy8RJXNi2k73lb4SEOq98sLkyCHaioEn69sXuFcgKx2UqoaKR2iaRhP0+VBSv3
PebeRxhC0PXVjtdaFxL8QE3KLEuEti6wqpWuzFyE8q3iI1OoAqMTJrxeAOoSBxMqeQf69oDMF68O
/bZ+InHmTRBijYwY71tU8+lJQAHT6bjZlk0dnGfgEKETb4uqn3suxF/2SBXOoe0DdwDatXI+JO1n
vzC3/v594TbqvHN+ilJvhMjsiaoM4ozQilikRq5TUh2aQ4loKUYYT9RxPxf2bzMqfOkXz0FrD1rD
VZuD9k/NuKqeUpbW9L41NUWceU4sh/yhij26c6lssaMq/RMHHwxqTxUeHFRKzP+ylQWY0S3Yl4wo
4bAmoC+bLORba40EU24FgoaGiHlPY7NZnbFhvo3DKnX0vwIf4zJ39XLwudKzyeymYdIdOrRQZWiX
5TFKqBGB4QCttiownm8ivJwFjqXU4b5FXo07A7M542vnqICWZDfuqstRpQDR5MA+lLww+yHE1uen
SwAA9FNhi+o1wV0iCXMUOt7Mr0ivI1UOQq89+JIC0TuApSNdTKjOfrWI/MONBrVSuo6QUUb22ekv
0ZNenvOX5G6KJYPWIHyYP+mwDVkdloQqyzzXwxr+A+BJgCwEwAGTiTtpJPLnhgPut+cqiMooLUkX
OeHYKuIOUZ7aopCGvsMXa6z41NxQvBUheOj2fyqtDt5+wNw62fA8Olcq70Zn4UysFkoCWM/EBHI1
ZKLKaCR0dCTE1X/S0cRtc3ocO3p91TxBnabdeaIh47M/BhtT0EqZQbsrucwsHY+li2UoVQmvMYve
Tu0ZvFhfraD+nxAavZgQXVomyrbmdQ92imrm6YFbgiEQiksfrWpzu1ppsGZyG6Pq0vbc1u0D32LX
Y5QcvMkXrQKtIhfKrV0DPTqdST67E+pTWRYcuqEjk49zSk9MDGS79Td+DPb74g+ae4x6KJeabJC9
Q4EjNzbKa/Y7Pajpr6cVWk6GbWRb5VQfzsFYuAarDPYL+LmHB57EokUlQUPrTwbPd8JKmTMAojTR
YxP28mLCrxhX5zIv2F4SP9jxkf1EJYWeBd1oXA5ETy84UgIOV21uG7xkSerZipcr0buBzrO8+c2k
R/sWkkubuXAchfdUEOXRE4EI752clkJMNNriDefizIS6IbJIp0fxsWhrlNxs25G5g/yMo771/+Jd
FSfZjPjOeTRNj2x0VsSsBD12NCQcA+bJ4YGsqmBos1aA5bprgDy9MwQpEL+R7LtTEuRf5tcg+oK6
Ji01GML7XFUHms3rfxMIsp+5g1uqBnj5ZhtH5Ucp3x7+EYwjkXaDSQc2AEJ8UoZRf15mbGi0+jju
bDKUHmaVhDAN8x2xy8ESPJYR0IRDiCPQJrsRlCH+51lRyLNLXITfIJEgKJ1TORMeBLJalV5N0ad4
7KhV6B698l6Sb5hJwcBrLUD75Uua4V3R4gDsGEX0UxcQG1zG+EbPauVPMq6/d1qVQgmR7o58cAqC
bGwIVuyG6AiwxG931bV1M7jOPIdX9q00z2Y33dUEgP0aAazAHu5QTVqGTVQAJMcUaG6nKgCrPwRd
ZEGgOtjhq3uJDxke0hFs9SUWI6b/jC3mZHcyLxtJPL7fWAsT3c+ksKpHlrHJUo8UPic3IaAc46YB
3WSbKh5E/dTljScxin/a5ArkSLYyo2m6Es8fx4dE02Ny01Xu9pzBF23PYMev+JM9nWtR4T9PYlcE
QVuL9nUWO+l6gmCdOcOFSMfAoaX4cuYjtnv7vsSVq6tbeaB07F+4gzYnojpLCSovc0AGC8w/9LtS
r0nPjXnpTjsSIaQBtKwUoNZRo6m54XNGq2DXHvT2YCeHjQ+hq/qEufm0S7nxpyQigDm4RH5qHnkE
4p2SMicXjVrwe8dvA4FanUbD+nmc+0VRqW7l/lHVQjNo5M+8obUppdyC/SjCDLFTPNODO1PXxHOE
KeE/jHwFQRaD2MGaQ/QYUwvb3r+KS/Pp0A8e0DH0aYjYlf9t7G8ibThM4GKZZL+mbRMg+k+RF9kv
UukJjs1wpw7UxVVyT+UNZyf3re7vHZp/4NRyv3Om9HdErnKcQuaoeRd19smn8i96u0eUFF+XEuif
j5ETWNaNXMaJDgagtZDSIiW617Bn06vzypR12NW7QRYvkEYDAzmHNrjKF0ehuLfXpowlhDPMb1cq
HAKS9bCaTOlOmt7z0luk6vqMyts0wLm9VYcEd4sxccNQGTddISF42sQpVmCQCgAhwVCbvLrwOAQ7
/0rxYZo0u/Kox6nY4mf4MJTmthqiTl9ucqH0GNxPCUb1klQohM9Mn3wc/P6YNAQDBUQIOP8hzSXd
VtGEu5Hvds/qiT6pcneWwrmI/6Qth47NS3oxioo+uqonAuuH1ALMyyOkfXnQ1VqJc/vhrvtdFi/K
a/sF7Musp6HaUOO1CpoJV83JcpbfSRIflugRP2HYJdmwT3QOeuWftlawqGbA67MsxWLpGo21oOt6
VtuHZYzIW0gT+BZXbBUxnCd2Gqhntu/HnEtdLXhgNWHoAVoqYR1CHie8J3JQHj0nC6DSOD+mu37A
Eaezpzgg5Z6RBj8ZAHsgxYzhVgRDo9xyT3Gj0y8PYKdGSd9qlu6xf/xD0oocn7I3NCO7s7UJpCDL
NWgAlCANVw3ykAp4/GxZF+aWIOkAJQloRzwDReOwgFudjn586HsWrFHkEupI3iDW2sRyTm1oO78v
BorDPze6aoMEN8UKRndx7EAqOJVjIddvZZ71zl7mYecsrjhYByKwBfpkICWvp0Qmrh3XL1TBFiVe
/vN6ozzgHTST7kwnH/uPMhhX+9Oc22X4WeKjJ3oJeeGXrgKyLuA3BRbot0bpUIkrU7LWpPE4/5WD
TfR+7iihDI33FWS0+HVatzEtFlXSRSX/yOTwwMv2HwoK8BoYb8PJokC3S6UP6wFOAGu+r+aPtdmb
gwuzWx7p1AzTTq0mT6T2T2r1zi+qzmcsdFvrEc9aP0a8+uGkgv/SaxBAK3pHDyRNhluhcjPxraB/
8ikgSoMOb9IqduPVlHu49klrVZ+yKYYllshH89S0uJ8EHEKYub6/vOCwigECvRnFkuokraup74r6
vQHZxzP8BxWdpYVLTAIDP9gNby5xOLlC3365HgFbjBtKdppT5QcSus0clq0FRC+nG85Bo/7ZH78P
5TYlBUQhMO6jcrCkUT7C4te9C98cLGhqSH3qiExyPJ85//8CAXeRZorFJUHN0IwDbnXMo90aoM03
ifPsyliWjTEJb7w1N5BrsUNbKazQ+RNmd9DOUBqytEaMY8UCZL1ryAhwsG08DT/zD0kVd+S4VZDU
N70PPaahRZGvqC+FAjjGLg2JlM2HNGEWlWf5SCSWd/Mm7PqJJT6i9IxhCxaC+SZHivj3WYHQAxtG
pNf3X0UZC/zkJKUwaG4ehc7Zq4ukgLJb0iBjaiDliQpWSb/u/jueE0k9yeT/E0DS1ECiHjv3omCU
yMBThHYPgcw4WpcE41ycBLKSKUfyJ4RLJHEdkN1sJAY8lcNGtOl+NnKkGAgFEa5RO6b/ac9IjYfx
wlFbGdQGONalyb7A2oBXNG5D/yV074z5KDpxV8JGLidrAh1sJD6oeY909WN5jwJhurShbF8R/Jvn
lx5Lw4j+UX8K7wT0fsVLGNyrR+ut+KLN1xs3kUwMUW8hpQ9YjGHlMk0WNrLfWGJihh8HWrEdgusG
TcjcbbrxSiq463oBsZkDSkwQNo8NIkXf/j41rQc9HBp9gy42DPCvAMqQrCrsSeH2G/FzXqhzudHG
4nGDZodLswSOT9NAxamJqwngpvncMbBFZ/YUo3ypMm/vX615aFSzEiaKa+NoQDdEJ+ZPlX1k6mM7
Cvfo3OCwrAWIhBGx0ufQNlhw+LX40FmgZhpe7WpjcrK9CU3B6boxaZcFYZ3qVafHH0L2nHlrfmdb
g4gWvn/voAO12jMcqAVD9N155WwvCLNp0U0LDYgCWco3Uo5xp+mKBAW/aLYWdMNmyAdzrmAvA9my
0RrLpFvaj+TzHh5Zt9moYAMtZ+AyS9qVFH13vE20P5W6u7n8HUqnYN4+jP7feMIWbUTVJQGVr2lM
fxZkHnyHq7uWJ/t3zWAao4Pr5UGOm3A+W8fOy7zXg7a0feG2DUINgDCtPcHfG0bECUa2y0ar59jV
wg/4+bo7uycFnehZjSjTJwm+kGF+HZaXK8MbgqSvFn/X08mgsdnrrXyC8815xeoQNF9jnLMTqjDb
SA+XBSgkqomHHkUlMPDhugePIJkM7PStAkVmG3XXG5vF5lZSwp+Be4mNTHIfw0xmPSBzjRfchSiS
8TDOLOI+sRlKQokxLV1tM8LyW5HJLBKd0P3wJHxURSKZNRS8Oft9H47NjI+VXKThTyy8RCTaLaUD
l0UMo2Pgn/7UBCtHihelUPX7CWKvOTP7Q7btEUK0aZdIV96N4mtZGjeTgq/hc+3f7rZU/RDvPWD/
Ba5Nth3ieO5kcTx2PRfYx3jA/0adwghcHu6Z+Z6Gs2YbaKYI3Y0WTAI4yHZu5Pz7mVFr2qpkS9/H
SiLQfnF3cW32mFqIYUDo0HXmPbISwpeUYjT11v35RJGRjk/dQjuq7e9KeswPexVhmGwFtBO1sGyh
xOkiQe5Vdd/g2sdgVFQPRYzWlPHiG6ksb7Bmsj0wMNjJquXGbxy50qN9dIiwb8lNpdm8cTB0IsOF
+m3Yxn0jKZryeFZwEmQ8gQj/AGSuNR43hm5XMl9J/R/br98qoT3NjgUJ2Uk1qb4rLO9FtovsEdhs
m0Em2QKqxsPqA7BE8Ah5Nhtb3vukAheiOeD2udk2a+1iGwqkmERixKY6fdys61J4UI8r+ocMrJCo
ZhIIYybk+kUIfYPHot/zeWYXOitf4MRRqIbtBvCLNXLDPGE+LYiIbYj6DV66aqNpkec9DU8n4KHA
epVGD3dFM7W8OZNjWYVXZNsH6dRN/oIp7P2E5TVXBSiYfzjFPD6/jMlVcUiHfpP8zs+237OpDqE6
wjAVS4faQqoydZL7SB6zHKUA7eqMYfvyfSh+eb9/mpCth3oLZvT2KiGjY1028d1U9WGt6CXtflul
kf+qNqs917qh4vWw+kk3yuvpoctkKtSoCAXQ4cW8/T5Y4fsPU43Q3rzNBKaIkFSTYkVfLudiE4QT
xqE0i7zeXntKAgDusjSYU+E0gdr58Y1I+Sw3Gbj5tMIpnQn9GQi8tIfa1JuLH1UVbDuON+mU8oXj
p1YyUybj4NcZp24TLVUXWmfeKSbSFLpHmSj6K+FQZPcb299RX/PeHO4NTQln+AaGSsG/hAhcXZ7O
aI5I98HkeqREIl/i7HzwjYPDN0g7r7jTqjZ5LRtQKZppQzwm+0Qwd4NLvBwUrZMtCGdEf+xyok+E
e+GzhbXDh7veaVvFTpA7wsTNCB7OIxibpKhemH3Khix60bawpFcrs4cBMXdQ95gznxG1K4yKPMQN
92tCi7DxXvxO9Vmq5NJCwyg0zOWiCCd94RhhWmiM+XeTfFkL1cXngj1bcUIBHGNqGmN/Bp878iRN
FSkNmLceDrmAyY/ZkphL9Rwj1Hjvsfy8fw8y3y1KHG5iRM/42jXC3zOhDF4ogCpasH+cW3Hu+GSI
1UoEwW8X/m+tk20yfGZ/ZJUw2aBDTbby09sF233qFv/cHj984av2O439osd+IRiYqAgugNVFkILF
yZpHSt+RsdIUhL3o5myaKE1Qs0nmLU1hZoqA2Jl99JfsvOrsLoeNMqW1w3DzxEXTLbAhOg4AN1oc
VyuVyxk4xbZPfXzJPYfJjixKpcBc5MjTIHRXXOu4AXH0IW0KjhXWtnlFOWn5fhWTuhs9JiHhbWsP
UXsIp28/GtCueEnlGgn/bEvoQL2Y9S5/vfm921/9cKgLYSaO0KHOYrj7jlizD+8B1Pzx+fBUBI6K
N93ucknAIS+yCZmR9Zy6EHpXGZdoq2aULWJ2KPIOXV4paQmFBJMaG3n/gfTzw+PkfjvnGx1Qq5+1
VbK/uS6bWnnfWAOTR4evItAJEc2ZGpMRq8icWKhOGsiEAvgHhd9nxsJL9KMP8nIliMViXH3yDCM0
KMeRGNy8aQZnAppHokBNpvS9wTYS1b854BzGp/szYjqBeeJXsz2BHIAK7e68Ki99fThp+6oTCzoA
1rSmoX3ixrHAvAe7+0nPRVD4RIFxmtXhhf5v0CcmErBnIyQsYgznIXMZarepLqHqRTYcBGa7YMWY
vlT1gJymuMaphccHmccHBKewww4j1jWyKg5Jxtc5VHJKuTca59l3ZtGYV0lilki1gaXes93tg47k
irim5KRW98c/mzWxclT81BY4df1GD/FqTsEB3Gv08JVh/guXNeyaeXDPok8/6HqFbeDPEzh2YfEv
4Y6yZtHSL+0lzgpyoRh5SZptSJI7mVWZxs0jVZD8bqtP5whNzl4PkfJDAHWdpqCelu8MPMKiz90e
3N9P8dDI8MDrrnS2NwsCyZ5dx9dAXG2HKf58/TOoB2N1yLh8LqEqFJOnCfqadr5reqCOd64To7qn
d+Q366zDpfRoGrnu5nK1ZAZiMRVa5WO75M9FQFd9lb/s8vD9y0BoD0NsCEstlUEqSeX9AK6bpTLW
yHeixGAU4mFzt6szfXJQWSsHp2sO6XIsT00hak3fAjTdgIFkEGQOv7Dsuwb9hrbhciLnqu+lsJC4
rJXYxDTsyzYEsbvv8uMqOFsafs3tzhEuLUbu1l2AebNJwI4u0oDQkP1hIkYyTx99H21xcwnt+FiA
F/LGQZeBD/sBRBO07RDdBaAqquqmt6PcdTC/yN2kP+PjT9C+e+ro+S/LGPRFAli9FTHH6k8Noiyg
efN19oOBIv2CcsO26Edwgsk3CuOuoIlFGD521KbZTo7DMMVrpuRDY0aP9BJSVWrkEm1ylhcSKFJ3
enYI67Pg5UiMZytEh4700d3HajtQSp8gXyR/BbaNAqmN/GJZ57SxfZMHLoxYM/rN9Oxf15for/yU
BUXr+/5zHClQ8GRU3FWb18HpPz8J8mg/AvzFj5ssCLxs0PGx3YQ4kk/88wRKE8oZ1g7mHr443AMv
n5enp/dN5WZPRy6zIQBDIVzhnbKE943Ye4LJ3sbP+Ar5Aei9S7q8GtEWQDXAIgkl/F+zZ9B0Qed8
Sum7XpX+2ebqiXBAerAIn863EGtPPPWL8d+pI8xzIdoEFllxSLFdHMziTbHQfsNoiGnvEtzOF57i
pCG7pPL8w3OjF5DYxfNhdQbhfVK1nPXlf7gKebOqTk5BWmz6Abanyx7AtoLXHiW1CCztFQxetzQI
aRY3/aFiQXtNgyGyPsGnYZx6y7ri+C59yxNnky0jxRBR4N5FlcQOF4iqxuSONZ2Cy5YqTC4Eqp0+
KnWBSSnqlzsTs7/roNUpSUOGLJI/mh3V+8ynAwvNGbhMQWPzyC9GF54I0qbKZEAuYI+y1DbDHxIz
eqCcrdSx8xDs8GJYtHAjDO/cAUl7JIPHLwvDLahANUTxgcfado49tIhZJTb4XfOiye4kidLBIXsu
EipA949pY4wEePRherjWdLiW6VBS+2YJUb7YseC74R/wloPw7k4aTCMKG0eMoRCfvx9qlOEfnR5E
b/MGy1jjwKqIU4ZNcxhRatwvGSKeaeZhlNeccBICbzPpKfoAttsDAkbW/uTygZhhYqYD3HfLeFgh
iZnZVV4MtYNdMyccaQ3SLVu+EwQU8r+jmWotTc9Z2ZWgjcqqWk6y8nrqiF1owNZd6M+o6yqDEF2D
57io2r/fsk2GJT5N2sp1YDZle3sEqi7I6jXLnsNMIQp9XLgqHzqGjhT47Q37eC4f/kWZw5d3gFiE
hpJ0pN11260FkPUsan3tICHIAeOjTY5PmdxdwDPOg1c4tJYYf/ACz30gJzGKOJtKNwOjbzL2p8aC
TntkW8GXGZLS7T1RPOf/C4iFac2gTWJoYnFNZ0iXH32DytXFjMtaIrGZM1cDGx2OLLQzuqdN9/57
BzKiyWgjRmLYoKm4I3fIWq2jdZXV00DpBGI6gEwI4aixXp/Xt6XwUfyJdnDWYH2QhPBkoW3Xs++n
chend56220tDLb7lC5/p+t9sPzWV1LXv7tLsH6VSaibc5qkDwrNFQvwAAYIcu5/GIVg21WeHlXQ+
a8vCu/733aiFFf0XcCxS2RGzdfVKv7j776baTJxx0Vo7Jp1RX0Q8QYfAH6zaGxN1DY32X8V3NuEA
ysLRAAnxt5Mo/rqp4R/G9BevbHFqeFlxK6Gw5iIpsgzi4mI+LpHIXBp58p+oCMtvyXj3kUItjy7w
IHWl+rcH1T7m2EGmqfl0Ui4DWGHJDomCAJRDWpXEEcexzyxx+bp/JdLKna5XsWr8SWDXSIBJz6Qy
mQpMgxMXOAy5jq7qF3FUAFDLgPW9oQKnLgsCxSF8rkfigrVYbk2+8maMQ3btOFqOWcyinY+GbbNT
cbip+nkoOwwNxeZ8M8UO1MNkWVT1a+IXdwn5ZqwHyTK4SURbQyo/1yUuFVdYydSAR4kPnpk1ZO+e
pBwxjYI6+uzo7ESl66OA2DfPihgr1vifDSXIatSQPh3Ek0fdtNvSo/cMBaK5mLm5hztqJsy+YIHl
FCB3wbpYQDM42ZCQRSl65EWby9unXPcloQouIBMQGX9E+RCN0sKMwTHuJw5mzIfciGtkvJfQ3Tvy
PjJs0JrOwI9fuF7d8SDeBaOuMUWjas+KS0jOMLZylNaOizvvHzmXZEBmfUzerVIqCW/9URtmnTw/
rjrelf2MtIhwuusWhZHWkGFr8pJx3qg8W0tmvNaC9agtD0oYX9IP56HL/5nW7Sp4evaCvPZaTYVU
p41fMGaotfpChYjIB5wx7OxsH/ZoxjLPObkCIdGXslxrIPqfWs+ipKWUB8RqBxST7vFElWk9u8lA
EPnAdwe6JImhS2vEY1tS+BsZa+dOtc7o7fMycoS+WtKWwnsT67i8JTVENIV1AuvbdmEtmnS49CDl
KLc7r78qzAJRxr/ncYeUeOKqiwSNrK1o15qJEagsl1r91Agh1HX66P9Rlw+6i4gChj9Bx1qpgPsL
llpRTZ7p+jRine97kzfg73WJaAnJI9f7GnaieVWO11MajPIlD8F1HGLkOfzyDblaSVzLW9mKO67S
IfeY8jYhPIcSp4wDQx8tdCDgz81kj5w1ydxWrUf1dXju2gnqspfqfJcqUwao2t/ZZ9i6HJ8V0FVM
t9I0sqdVZ1xVaEluBI95wyZfN8zzLBY5Nfgq6CNgUx23WvbzTeL7UBO5lr5f09x20z03ALivZLUV
n0TdTq/7emSHW/C1UPxP6UtvzltU5Kdn2uSXo3TYb9uDAMtkciqLsJ8DE+hmnU9+4M8SSSkEcOg6
i/xEQq2+XDt22+y5qHKOU8izrblbDPbdbED3fVHIUBTH1jicyGVX5iYNAfYm7NbPp0A3eOdTu/HG
Gw8oteGVv0igDkyb3nshbwwTp5OYI84YOEfSq07n36VucUWdN/EBSzYH91DdFtkw9yejSkQtsXcY
7Znr1zw4z85GkdBBy5fK7HXEJlqqjsYMxt5u3kkCLUETsu3DRCvNpzC7v2ibvPkb5bUjxWmXhaQ/
yoclbQo9gPOXCJFBrSlNrJy2EOvKVK8tn8wxZJX6mb8wdtKn5u6urkYLh1TB79Z93UpQpMUTVisP
Js1f7Oay39V8cjXWYn46D4P4/OEcvSFljFsRRwjggLhNt9faVO6Oct2Zq6uZTD80eENqqtYnHAY5
NnyO4CFF54dri7VnTxrRA3SapA+JKCDEbdCAoaCBxjPwqPSZ2aElk/0efIaOYCIhLeebkcgSvM8M
y7mOck2IS0/h7TWYrF1ijOgimY96qqmY5Za+2mH+6MQ+jsDT1w5zxXBQ23dpFBSZqk2scm6Tnj9L
QWqRaaylazymLf8Hx5traWt6ZnMEA8z1V2D0luhOVKT+Hm67ZiMGcsSpxLQN85uEXcEDLFPVDS9n
0CaT+VROM0WWGuwvBSeMGve8A7YqV/xXVBOBTVxQ1Mul/qM7pShW7i23xhH27AuwZAnYV5MBDwvX
+0x9qaqceaoDdlGS+1QcuP9mMC/VTIVVtXJf4ye1AnuDaglv35tIWC6b5J00eEYdJmUxThlHsKii
eSidowj2rB1eer62VhF2j70wCfZMUENH0hdii+WrY7Q4W6B0KTlCU+/mc9IcYql3rvZT8J1demFq
Jr1ayO5IesGfOkwOlQeu4FUBl5VJPVLHgdAkZz7Nm3MX1bMhvuBzOFWrOIwn4fZfZz+OUNisyj2D
j/ST3NA89Z9IkcrKzJLMaEnOmnX2Dt9oaRzyUz/S09h0mHrwhsgJ8+9hJPl+C2DG1zfPFdPge0mp
PyfyjlSuI+mBseLR7fwGGs+0sJsj7OgqXzEu63l86nupmBAKJz3twmIoTb9G7ffpKqsyfYIlUyLt
JDIeP0Dm4fvEcsnau8xM1Hry5hdqLQoLi27PisxopAClsLO5pwiiJnYx1h/Hcm6gJ3YfCqeK0tBS
PzqbPkcN6OtULzRSzAVqbG4gs04KXNpVrqcJVfqaKDKIHaPP2a8ynBZsecXieM6dFK2EonJeTkne
l65lmDoQ7F0ey0KlYzdSc6W4RI5Fh6IMPsUUdARRQEIVb2DBBhR0izLy2FZ3PzvepZDDluG8G3wT
AjpOS5FAnR8ff3uJrlSMstvp975by6uKlMLxSW0dcYQOFzH5ohj160xMt1bm57h/XkhLnOVlnQ9L
ht1UUdKJnfBYlpluQuRN3wLDKsDe/CxySflq8cuuU55aKO4iyZIChpxYNs1FSPb8DkXKGgFkLww9
8PoR2FRkkA8mlKkji+n5HScaWmlS9gwZDaj+xusJ2s+2IKHWuA3R5DEWOvksyO8Bvf1UJssLUEWt
N6fVfD4+VzWJYMZdM93XPasQ/MmGFvOhvAN7MyqiWBTNo+UNOzU0g9rWn9la92vCXEYTWh9QDPdf
dO3eA9xpy3/MXNa9jeuo0IGJYV8dIu+YoICjtUYEmaxOUi9djYzcVtyx6QO7DRLLUGKZ/P4c9Yuo
u1xRnxEvsyTR91EhkMR8/DYywADEJ0+vF+9TSbIrVKL1sfGVl0VbsAdYgPlno8uM6PCmaPZyoSXW
81hnEUqb4PXY07LH1Gr09FukLiY4r/aE5tClUSQD5MJFM3eq53ebND6RXg9Rv/L4LKOS6Gwj6tpo
pDfPCbVYCX8K1KXx0rRgiJzkc9bh9La8qaTtbdV0u8bZWFNZtMnmd/7a4iIe6GcIr7GyKKX72BuN
MzUjKsu6VeZG1pM/uOiOtl/XtVsLNxhp8gZQwknP7cSMxXNldfG4asJHIxFD56EA1vXDuJeyR6zq
B/kVOVLzwRVm1N8wMHKbdxmttBPElpMzCtjhlMcu0dD9MYwX7A3v5th8IcVeJafnZYFdZ5LU5wZ6
nRAY4QY3n3Ghhg0MK2Wz9PoiymEyDxxYgyqLcWH38yTx/Rr0jNteS4+l6JBK/rkHKPo6KepkxK8A
85ZSlj7U+wrhXKMXRqVdPLOXcWH/1QOGJ9hu3wgI5vGI2/xyEEsK37QBnHEZJ5Bo7htNRf0vR+Z0
SsdcOlcKYwF3N6U8YUehCEQ/2nq8DKyRLsMPaI2d79m1/VHWvBglD7UDmhIS8R/8pYp1C/JoTybm
WLfmbo7hnpJHjguuWUIPfDhf1vFLzNH1hLr1CAZOIMARxVpKz+ZoKbfbLn5omGg2CaSyRH6gGBbc
fn1pP5tGqnjSs+h77Kux0kjPPgCxhVgY5J8WEM1z32/MKFF8gIdpZMSTnUCI/nqui74qReh9WU53
vxmQmYbWsocPs45O5Es0KmHh+1bIo1M308vkvgt5Dd2if0ZUXatX65VklOkstPlp9nkjvFXQ3AIW
Xrwfk6+EtE5mDIScQLkKfhyJZ+IRev93WOnDTBXOs3gUrUvOsec16eae/LXZBYPWbsvsCLlqhAmz
fe5mMJS5PBN2311VmnqR6Or2FDWFUkwACTCnii64Yz32Shs45tqZTesfKsQyXUGon0YgsDZA7PMG
g2OQzqyLXvEqS5SbRqhMm8wdT7f7mxbxMBGcKIbpM/nmLa3W0fSc31h1fz62pG5sGVYBhCt4xdE2
m2Wfu0QzP+z5+Iyj2Va4mPvtluTvfI6f59B/9vYXlqB6kHTYo1bbvSF12qK1ELaUnak8aOiJeQ1r
uP/Bajq/WU/kdCXSHBvM/iwVcEp6Uv+1AkkDTcizm97KWStV8LQoaR4KENKUKfIA6auAIscMsIPo
1HDly/pl2j15zUBjAMZF+JMIXvbLsx/AE4r9MU9pLWu3mQQ/7khW8Sx+AhFYuBRVfiApusYiQzpj
zy1SyHpYMJVhSse16+Y1Spax0knhSa95cVjIADqLQ7s8hfYQ81UhUEkCdIPLkI2FMmbDHalKEfyj
opX6EzlmnU7W/ycEo3TOZ+xLCQKkC1pdcebqzK9psJclnfsjUHwMfOYFOSWchVRXrcg5mG2yCXzx
wG21V+9Dtz8y6bJ7VqS7obLpk0VnKNEhUgJKl0MXbkuzAvsFl9VXpBhU8fwrrvuQOeRq+QU55jPU
WH+7awUITv232DkJ1vy7KrS6NyhK4A3yCzyOKPF0T1ZOpSKBzjAp3Rpu2aFeoR7TN6YU5kVOYWPO
EzcGv7O3/zlOI/wPHpwN8IUJ1YpfikuJStd6TYB6yT350SzhUOPts1T4D0OVhX9XLduwEsduHuPd
8K8MEjK3u27O1E79buQefHZXV6hD+VkrCnqJ7vVoy0l3z3a1RZwIdRFQIYHaFVW/kZzzgRq+JN9S
9Ug2YrKKoiA4/nHh+mpc/hBp9bCU0yyENmbyc/VvhyIixmJK2H/SruLG9UnW+JfhHnWOyo4vrZjj
eocc/HrRt4X2QeI8v/YkgYGQungLWy4cQev2fpKL9k3WVBv+ePu49bzAfQMVt3pcNsiwSwphsq1G
dFCggdzoQbzRLpaMT19fycYY6iM1YLLZFoF6WWtEtjlQMa2RmIsBGTYRdtYwcZpPcVHWuIB3jcMy
9yqOWBvNj/wP36tWK8pb508JN32AF/DX1yIzDPtnPzKduH9ZQnfvkyXgkjT7FJhkGgH6SB1OQ1FW
J8kjaxpilZAfQoiVXEfje15HhXiMbE1L6RVOhF0vqKL0YrSJ27XVP8POCscr8FKZ542Aga0rRBIN
16YSb0owb2ebMaCa1YWxrtt20SkBLiEXfs5xuTHNr1v+pf2bgvcI0i7Bk9JWZXHVKEu+s44cfhxW
M9y4KQfU6gleFQi6tdGDNAbEn0JN3Z216t0qdPl0QLtHPIqO4DcVVL6uNbHm24GyIhHo9jWZf1sd
uh/4XdqIsXkleC01TOKvnwPcdz3cIpOimURIQctLmYlFSSZRbR9sMrSo3ILXFpmCjXACXSZMLVfq
B3wONudk+PfqKQ8vwl4azRlKrijHHCWROafUqWo05N1xQ2dtxp6WUy1j5Z2vv5lAEi8pI+2nBlQ7
2KkfI2E1L7aTfxgQJmRhICJK+SCFZvp7BelAwfx6M6NOZPizYDro3NFJYA1YkYSP18dfncGQUmzI
j6sJzJD9FbFLmsveAWjIlaUahMXI0UUVLXoelrdnYf6PecxH1uiC0MehlXOb26Wd/Svc/YhGOR1W
AuPwt81jgLdituha1VY+Xk4Gh2DS0Do59BqesqGAzENQTTuR30nFiItfIrRubkG/xQ5+tWrA+qJ8
nimXd/YhPVi4JlalINE1WoEPTReuWKYT7lPu9f/xpnCSnI3NGsjEwp8sZN+2Og3Hzq6QG7l9s/Iq
HrhKK/9H8RNRnYKAK5pHLd0NTXh0qTwFzH/qfKWeXHHLF2fYrdXq/qxmDUM15qYjWxrbH6ZFAZbo
Dgtlkn3LAio/kOoxVkXy0jz1l9ziosmmiVezpckq8fDQzK6Cyle9RnPmfiWRcvJBqyW+3+oXmW3j
4vHrkENZUej9mnYjk9shU3ea/k5836w1tVrU/l+8SNGrfzrwN8an47Q+kUo3vOn8+/Yc6EuBO1OD
xYpWfDDSwK5/U9hTM5P4a4SgIKzYewWhM+EPAgFFZrKoHzHKl//im1SeQVX0dzbYIZIGOtlQccm8
OjluflI1k+fe6+dM8/dZJ3n4T6c3bR7IkIZIL84/H2Y7yLIUPX4NmLr4RxhIJ7OCmGUpWELz5EyG
jzjx4cYAr/nkPu2hLvhZm2B/3Dqkmba3nGE1cY9oxwRCQCnW4qNlxRyqa2uua+8E9MsrtntHbZTh
f+FSICF74Wi68MkNQTSmnMz+5jRvQoUiRz/ATEM+FM1bCAEYISSjNcRiPwMQGSHU/XzTLXNT9d7y
VrrUfvSwgFHc8quT3VRMNHmsUTJ4Lb/8/ZmOWO8rrCs0m/FcT5pmYOXl2/8V9GeLNZPJrHQPMG97
19CYdMWagnA8e53ocQ/iaAJ8hBf50SWWP8sfU+hglpdKJlx6FlvyK/V2hE9tXxWaYENoUXI2Grhs
UgTayQn1q+sCrtoqtG9J1J8JGsXjj8t+aCMGhe02pv2Xccmwb9m6rpvYnYW2fibXgdm+tP1BA7de
y7fOTM4MOTNaJcXVjI9PBybLcMoJcq6zZhcGZGBYSiJwyoMNzop13ohb2At6YyNa3hU9ZAx6Ihyv
utD0PvC2L9yyRDUnI6f3z4wVu8PR9vuADbtAUVn3+uc5YYdCKlSEW28/2Vf7eStADB3w0y4pxWgl
h/w2oB01nuc2UZe6ICRqSL9J6RKYs/Zjid0BZlbi9Qy7zgzLqMg/mtQMx939aRwH41z0CBt6LK0X
yh+1Rb6Ag96H3LFfjVBfrEAf4sSZMXTw+IigPPcbTiwU5BEkzWYN+udm4AGM7fCDXguYa+6fCUlv
2fBobMKZ1/4Y0qg+Uh3wSbHBDQt69cu0TUAyC4ebSX68CO1/bLMH76s1CoLtfzVecJHbAoFRLAHO
i/diofEeJ8f1PgYSwY6nFpHuUbwglmk7Q4G2qdweRBYITuEFykFbNF94spAROYlyIYj0rvOtmp7I
ipxIh5VsGYAdfuOse/1aR3D39Ds1YUPXq6/0SpSGIUMf6p0HEkQI+3k5dgcUapwvtyWNh7V/ugHr
MN2gT/6Y5YU+sJEcJ/veGiOPxgI+DV7y2Eo1aNaWXGYXMegAkduIaIdni70NcslcnSyIb0zhdhQX
CjXt2Ro9wp+9qjq5w7MpGcGzxsfRwozp6mjuyD+lwGtFbpZ4vnOt0Hq4brEo3P2EVoN7YNYurZrL
7e5BL+CIhD+PuiWc+2IpcIqXXGbRLoNN2AsAZno5P5KUDIyt4sYauqkZ7NctQX298CAmRmBmeBjH
8YnicDVZYDJfArJEbWF6tkQLxMbsHmZ8vbcRfxPgJueV2+JS6EW7xu9g3AKYaNOYB6B54X2+GgaM
xG5DgJ5WLNrVmBjA/3XrpPm4TeAlBKGVbT3C0pVzMcJHT7Ej2cJea185fFyrvnNpp72GVUXV0/oG
S1yx/njM58290bxXByFAc5KUQjeT2C5yblRiHtbo7ygQ/pdQgYJpYLj2MDfIvN1px6vNkJOJGVtO
ZscW2PQoeZhP+FxPib9AcECFCVctdQzrsc/W5aqXfANVQc1n88ESCdcwRIId9cRyJqrdPyeOLl//
BWZ+SBiZKp75xQAgTUzc07T1NAigM8yv9GhxN9rjJodARoIcbEjkN8IXY83QFgGZbQV3Cv3v5dVY
l+dTN2a6hKRzVLXXc4wfXTuQABFJ+eTEwG0tuINSCIKKpBIQmMwIxKwE5tIfYQmqQQDOJ5IWbklx
zRxf9XioygLxR9cMbmfmCAUWqA2BT8/66T2JHsx1wcw0HyhPadPbZ6kWpq5hQMUeVeFiLbsQ7YVi
bzJCs3expgn9xVZNHVJ/wCUXn7kDJiHuzUCjmMzrteg78xf612asPCsVHd24zMKEK+OhhHePr2Yi
Mnv9QhCmb4b0GWEUrmzfQ9a0IN30Ivnf8F4Wpiw4ctkhtL31Dm9IfBQMWawy1Qw/+aYNykJ7Tojq
O2TiA/GjpLMnqW1mB8KyhSTCjsnqRUNPqVHjFdkgymPtpokR+qSzPdv4A3GxAoGYgZ3bCkvi2mft
WTqq7QexLBnYzbqC2W3Ry3rNYULxPvOCz84g/ZzCEfyi23OUHCt5Pbo38+UOmaeG6kqsJCgSIOE3
jyMuUGVb6eQWsgpcxupPL5uysbAL1OIdu3Mc8psG6Wel4iTP+fVKinVwbYRunRBXpyGAbutJSfTe
yUWR/Y+9UxfevnQrs49SN/b/tNSgWF11YUhntWZNujPWqo8nQvmg/2ErMgizIZDmdPIvs06QPJ7A
sK1bx6K6i1zP935uaWCh6yaQn2DGyjH4Es6imOx5vPU6z/tNHcCHiBR6Alv+LiJo9n9zo4KYeBFv
PjoEEqZ5hSeIL2GVcBATBbWh4czDk8G6tqlG//p9sUNJ0XJ7GGUiKAsyCrFsGqZqidehSRhBQ/tt
mT7+LhrXUgg9+jloXy4pcyAW6s81d4XEWf5ijg639q9mwjfCbObfNwZBWpEGsRRjQ7ZpLpbNlU2s
Hq7yCIZamvjY28Qlp+kct3AdRBKgUSeMIQ6H/WEPLxAmeu3vkWhOeP/ou29rMz5jJsrOo2Tk2Ccz
MOfi/ZJkUxCWEtyFFdXTHZOTYjj83ARlxagJoFrkXWIANbz97zqbjJGpvpNtG/xklrH/jMsYN5d2
oGsOMX8toQNPOD11q6JStsAcVXI9O3HDAd7jqhr2GvJM9thAdRp4BKKuD2EESOmqcIRyFXkNYrCU
uznTVTW8QcUgP7luaUixpSjnatb+N3bUcwaL2vKPQWodFsKNBpGJiwB/JXD2j+LjpWc/zE7vIUOq
rI1Q3jAskW9kqscJsT7XzTRgq0v/oLVMbwmcJ+qQGE44RmqvjiH0/vjk2gH/GB3Niyz8dSn7KZYe
o+O5EKZTE1Yv2RO2o7Hx0HAi/xkS6fQDV9euECXGwtf/G99LG1s9ovxjPQBkTQUBoiByWxjUoAHq
tCYD+KHzzBhJYl5hHW+cgaBA4LRPQVznsDQWQ4T1CiKdtLf+C/Q6C7dcKSKouk74tFvwNGy4f0A1
gJ2csWFKZRwfZEROroTSt8boMf5JvvptH42ZABZAYiK0motVbkVdjdOPvQxUWdug65qk+GhI3r/t
ReQaFZeERWBNaHZK+oHE7T67U9mqxrvtr6EwRRuzLPOEJdOo7hWSRYYcWwgGzL+Eabk/Bu+k5T1R
kRQzT8c6iP42Bbpyk1Zb60+RUiZ9ybpoX/E/s6yjTFNjikNGfDJrxRFUUKcC/vdECkKAOx9rn08G
yhdt1SnWHkEkJ/VfdOh91MEC10IAdT0SPiZR2D0GUMl/ggCsh3t8Zzs6aAN8XG0+isT0PsZFKNKm
1AbU+j13lKuOSWf+ud5fG3Y8ed45x7UYCKVF4nq8AzJZ8Ox6w5jPwS/JvTe7FlpXSBWQrDO2G4zQ
Z3WzR7t7Gt5e8qbznT099nK9aJRzRQZft9lvz7rIEzM3FLlkW1H7hcOzGk2QRktpHftj5XXk2yCq
QIZ+kHEnyf283jaTWLXx3pUvDrciFX6/O6dpVQO/s3SwUgwsx8HfGe09qPbZHlwJIrGMvJO29oWi
nof19/GxtTpW+Vo2YkKG+qDFSAlZvVgN7eLO2rTo7jjhYAOsnFfn8+r6v6GzGOEAoF5A6vXeN1y3
Y2TPo1zO3c02/8DwL+ABJlfHyjK1jF5yX/VlHB56M0MqOCV+8N0ps1WcXtr6ftgTPE1ikRHe/ebu
/Gv5CDElqlcQcFetxFyYfQRRX7IeXPqdLGY9SLf96KkhoRsIX5ISkn8OVXTChNWFyOzQJoL+6MlY
O9wLDLDGO+slEna2LMInf0Q6IVP2/F8aU85SUaenxFwMyoWwrqklaKdov+6L4UE2vozKuDqDci+g
cXOCew0nH4LwklbOpIYWXw4r35Z+xJxlY+39xFJQxYhllzhhyW3/HrWG4+IEjFeYLlqtnxReupPD
PrStkXSqn0dTlQIhaQmh8JKYre/0UNltpwSPjl3F6BlYQt0Pk/NsIbsw3F4o9SpL8Xn+HVzyIvt4
+KHtgoJvP10AWkoLJu1Nw25VNcRqd3CrwlDjWGBte7cRkBJzO53a6lMJopd16BPljarDS3hhLaQe
e2wt2BHeyuXELpTqApY2lToe7WQfthMiqUSwl6gPLp/hl1DQW0b4fkJwjncEzf1R+M5loEkPyWUj
sbQi0EmrVAhPMeqaBI9jSLSa/zXNhcb/jTzF03VeTgtyoK4wSycCrsG+6jACvXiVn2SxRGmILfRe
f09c1IXPAAedMt0J+HDkAcT1AS/OYhJjhvap9C4unHrs9K3GEytYeMjVh3me9Wbxnuzx636LeTj6
L5vHW7hl4ijiJhnx9hO66lKhXb/Vs9Yy48Dz5EUK6itkAY7KsNxLMLpofz32g7KCnlxVpFzPWz2/
OOzwWCdEYPx/FV6J2D9SjOdHVkWVnY0t7XNMYIBAQvGYprlGHNRsuGfjrO/TRCp7nJZuq1pUZkrO
5icTByf2xFcS30HZE3NmUGpk7bQlyPlw7+G2XVUg60O8mD7mXFVn2JyEFe0xrCMqPEImi2Dnpsc1
uc3FaD1K8dABCs3ppXEklf4j0zAr3+aBBtRdYMO1GCoUtboW1XqT22k+GLrD8TDPR/dr6g3kLSKJ
zhNNPcFT9KttlLQ5K9MZeL2HJfLVob9zNJUlhG32looHgbQAzIK6fvzkXshKetDuhK6AE7s56pu4
NNtaDhhIqCZiuAsWmJLdlk7Z3YdayrmkAmLf3h21ag+1y6sdagTOQ33rOHEVlYV2xsXaDVbSGK5H
CX1m0srn/vZKt/VLDB86fJyDCaAuPbkcCT1xDgIye2jS8rMSMNWviQD+XXUOPi2QRyja7x3m2udD
mAuyD2OH87+k1dWXplRwQCSqFpsv1ONxKBKyEUfXOqGuuDBwAxQP0BUF+2CA/Pb61ebIBqiaat5l
t3LtzQToBI0rjsOM8GbrjVw3xh21hDzPMC3y83Gc+sKqEEAzSzgzw5C1VRpvE9GklV+BWV+uF8Ax
DdwENBu0xEjS0Y4kV/optNyT6ybGqrib3j3Y8/NRTAWvDB+rEoQ55f/Lah4/Iw+awekHSVNAPgw2
JeNXDzijE76DzLepIGjHvoVy49gCvqVKXB1nuMUfp58Zvn77ETTdqxFOJ3HWBvAe1DbPI6CVVTSQ
SDTor+R+xUdg+oqTyZTztzHv5QvTzuZxHI/MkB2yx5Lo/UZZsrM41FZbIJwGiOMGYstVxEvWxSjw
eIRdlSytSWqI7kSXP0zTQ+zYqBA6ZB+jkIhbeVf+X0fH70UX2IIwAN0sa+lC6TiwyzUihpxaegs3
5yYX9YgAirxrfc/GiboIs4rMdtQ9N5zQTLso89hIeir4UlC07PcWGlIyHHsvDfmYssWHsQqRV2Lr
yALoCytd8ik6q9r7kd3xosRv+UTw8AnaKgWpVEJ5dXDiVsA21zSt9ud0DGC/ifVKxi0FIZr9jYGG
EAFnwPBEBcjdzwe/AHksn5gpWxUb9beNq4Q/UrZO8bSI78nCrPHXmaarIzOfvIz0hHTzXTx0Hjg0
8rTuNLvWQw4yl3+uqHgKpDrSi7VLOYJfK0EDk97rxFClWk2zwzGiLRyBxoTejUOj/DNCoE29pzuZ
YfKv6Ci0irhbiyuVXRAbO1UE0bB4WMx3bnL0+b7sI7Py31yfonC1vhQ3xKqT4pvBZTSurUgh/AcL
D07UK+CqjCwAfCaiG+QB4MrUSy49HaDv5SV3mXyTTKcm8VH9LckTPPonFNyYZBeyd4CQtOW7J2zM
LP/t78ItJ8GVEsuNxSIg/f8Lfk6P5VidlfBl6qN/xIlwZbknFT5DKpU5nWa+bOLoQQi1JQKbq5jo
t0ItmPJGvRWECchx1H2AvYpaQg8JmH0tKd8BYHd5s8yTzucBikvX+e5/5ENc1+bXhgaK5XKVv4ow
P3NnJBmS9RjBcO0e/vD3mmbGZysxupSWu6Dj++CP+7oCmtiwsvp+y6aq9CvL44cHMoE8CY82FCZg
gcnA5uLuM1bD6fHCTrHV7jY5DT2O23J/5rWqP98Jsr+aUrsbtl8/8/gocZBSA/Jdey95naZMp9Gn
CRvbf+MJ2c/XzYWmIKnq2Y/HfaHOlUFnTsDNIvNPVm2DG3qLEqe5X1k1UNj9I/u1rL3RuYC8bYuZ
cHJoh8VmXVDMwGr/+Q5UIFwtxEOZ/cnFAwdtg6dlz6ZR7AeNvqcCSOh9n9uofUGuBM707SW5tnIK
80G/ZSrd9R9q1X5DNaN1mfboavJ30O2RjJyKgwwJ6FW+HQHJtiylznv0AVhqYd7kvyg2e9we3hAY
+lCzos+ri6thCa2BJ4ahNkW2v3b02ZiG2Q4UAaFnWoqtq3hoZczz/aCzmSNR4vU4i4js+rh+p1tX
+wf/qX/fPQztkDaLU6iDp5pE3H+pYK9g2PCLhRpydkyONb2bjvkdbd4K8l8TTKTWQwb6Rd7jBbmC
rT37KecZyat6654pmcjdADF+toEUYQISpRMhwnuCvlXXssPYJbIk5Db9tDLK/AqxVPjtTN9ViXcA
Kj4E7xF00wp24OXdBZIRVSYg8nTvmKt2GzP5o9KlT7FZnH84N7PNoQ5wO50b4Puxm9ITaNXD382S
73gzmN1dEGN8X894IdGEtUsP3hzWNGdays5AV+qXvhWq4Wtk+L9gTj0qLKAOVLjx1I5+ocMsWJJe
WbA5+TH40QeJiIcJM8nmz4gXcH8tyNcI+Qih47O3gkIUDZ0NR2NIlXRVL8Y4IwnnpdrBWCgTeYWw
gTl0ZBwNmVcFhjlhWrXKsscqE0752GgqObVBKl/nPtACU16UjwrbPqPZ7Nw+DqhgeiNkCPYgoHoc
xssFOHKvkRkCdagb4d9LMXbP2qj9fjqMJA9dPyyXIG/N0NXU2jLAA5Kbrhxa2JfYHL97DteHn9t/
5IIwuF3P7YQ6n6YnEktsZdrPsxKdKqhTRcDgEXqFB3Mq4BRDiyEnm6T6JU2rRcFoZW5zUWDE1UUE
UvELbPt2PLONGj9AAUT659k7biydEWcPEJ+1ahnllsnPRD2j6GPBU4Aq0mHwyK26y2AY3J75vAbU
QlBv5YveZFYNzAP4n4BnNg5Nsh80c6cedUt9AkS08AfP+JN8N7fjR+O0vGQnL65TMFj4bNI1U+rr
fO84RAFeLmfUKAHBge+d6b+gVnES0jb/teG3QLBdRx23GIDf3sKgDQlK2E7RgzEAX/V8Y95z+w7i
c/fGvyjaP3aq0Nedo7tKYchud60naSN/RccLxZCt+iZrZzYrhgs/6w3gq0jYqkv7GWVhfHviW3rN
diseKdM0aLXZcxyWDRQyC1LjpAQ5iF3WGEarB+YZYhrK2Wm9i9jTYSct1yX4eTfcuAHq7N0PE3rN
u+r5bLoWidPm4z6ZgM/0JXa6kuORqyBJqwaJVqh40VwaHbtBdAs1uLtMa40RPOzaGji6dS49RQau
yoQLxnb5nKul7jWZsvI7O8a0Gyl2VD17NV/1rmNlBErMoNBIJcIyh91/srayXN1NXGLNoVqM7t+I
AB48bWPDayX9iZ7befhBKN5hCyyAT0BBJgGR2C7lXcOxiLQxMdaLQotHgwBnMK7G+7Tcu6aFh3gF
z5TLSUPVyTL45o0g3/3IuRcRIDQW0w9fRY4/L3yCJXEnBvZ/D60n5wksLvtTOqY/bRo5AAPFNy+V
4O8D76HVRkaFD0CMBwVjAe8iZqErl+SDUTNOV4AyTsiWrs1T1WgRQWlO9rErdHHnBCo7N927SB5K
YK/0Dvm1zTPIseC7J/xCm0M18uHr3Rqu4TmWjoFssIZDLvoLD7+e+2Ir2UqxihUguJR+AwknviYb
AujRBtdAVm7rW5nfWAJw6jTkLstBWtzPdmCDIbCemHA8iyUr09Vw/hdKxAkel6AK57McE4ZcE/qz
9jfCHhtl2G3x2P2YCjtpY4jY6aOg/oYC370FbCgqWmUtUZ2pcDgA386H/emG5E/McxMB4e0xAIqv
uXpAHm14ikg89h9+kBXVeFQU0mzsOjzddlnmgJsQChcithYn2kHSn7O4xTM8zcbdpED6v9t3vkxF
4x8dBQpc8JLYYYO3irCHdYOJIq4OLdsz7ud4s44D53gSpag4lq1+FT9ywNIlGDZxXnRp7djKSPHj
cJ2BjBTUemAotyqk3dHYS72aVm1gchH3pz0/2R/3khL8zD1mv216eIHjPbYqxA8KP2DD7by3scKN
x/ng0SPqMBq+H/RcCFm08a99E7yKoV5VPsnQ67zaX85Ft1+nBs+0A7eRMeMPFGW8giekB9mEEeJA
Xn4vz1P0h9dd3Lbi3UrWZXS4bU/kSeVv8uQYqSdY1laLh2ht5m7EGc4FBis9tMzyjFnx0c2LjzkF
IpXqqZIHhjkCC74rLXfmJzQqVwlsRR6fgaxiGHAakMCCX1tokVYeGlSQB8kmQlZWGH3bMjSqLuK5
dqJiu4Uy6EsjdsbHiyh+Je4CpakRrKDAIYBvqGMpAARdwYeTsZNjU1uzX0difh8Hva6rTHL7LX8a
7Dol4uED8M/Wk/PXMbAONJTuzjxOiIGYbt4ivWqi6UpDuz2PvR1cfDA863ByY8zJxI1r4FgBK0Yh
sYQI33Vj+H351cONU47v1z10Zz9ETXl3kc0fH1sRbzOMGzBm8VI5867sVFRdRcpgqOxuWrVke36u
c7w0u9A+NXNOjfzlb3Cw5Z4S/B1OXVArqwxLzpC8wG6fiLRmpGeGb/v7/+evDJWTIJ1dqTBlaaGJ
9sXiLfH4S5St7sdKQKcX4gTLLbbkgJMTDAv46Ivv/6HmzmbbBOOizJbo/ttz569pqiUK72puUoDD
vlsPne1w4kIdaZANn/f3v5pkgFZyKdGlTtqTGfLjbY1bmBr0Qhaf10XJJoaaMia0JsEvsvTgy/dB
bFGHCuC9cuHyYEF+gsK/v7X40v/JGA4kCNOdyDVBYBkVbmkYHPHpeCzWFpPbP4fzjWsSmm/sxcw2
nEqg+QtUy+wxxGfHFgzrlYn7SsN8mbU0pC1ofE2Mx7klGZxTilBGFxV7cpMuR22jb8xNOhwphom8
1m4o2/jq8tWbWD/8Z2DDX/XgLStdlBcpBEVZO/rbIBgmC6KC4fue1/WUyQUB1VRiGgWMmkiAPyi3
BRwnMPWlrHJIkVkUcLGOnXSJq2nPwgALRWaZuGuOW3t84VIs094sHR8uNuL5xWZvnUEZpSxScr4X
8FUtsbAb7XCiPJbDCEsqtH795P2K3cPUhR7YkueP4BsDY0OG7h1u7bGCm6DZ4+DFzJ8zbkWaEEAw
jTC/6vbXOTbxYz+fNMtrAFvEFh8jPpkE1AyAKjw8Irt/Oe/K8pgqSj/NM/Z/ysP4oKIi73qDWOPE
AltYBwDek4SfTn8Dl0ptaJCgheREg2tmyFq5xVyK0KhjIehY6G6tAT702ScWQg7BXUXjIqUEGDtN
hfkLQcvKJWsrT9l4d5ctcGpd/ZGibPsskexWt+Iga+m89jOH8n2Ye4X3nmMnTZi8MLcdyru9E4e2
0fhMYq+X1amGy43UhAh9rbDD9cRquHw6rVsZ/2nRGwU+Kcl0BF3734FoLHqdOLV4cQJpTSKrKiMX
YfaQBuvhMFa+swn9Vo/ktVZNTaw4gvungNOA6/cLWZWzemLE/G58TWAy7yFykwmJTkMvnkuki+eG
7emNZoBg+Y80XGM0m7i0ZDkqIFs4mL3TgcIwaJKCyC29ollgShggeiFWEt0DVu29gpWAmKUmzmx7
PMxPxJS8PEgE5oFbfyzUmU4Nhp1FkkN8gTGR4jNG11DSPJ7epWA9bih9qIp3o5d1glNuRFOx4Cc9
JzTF8i45as96hbkf8zajg170P5wcW/rj5ULaX/YJRjexpLT9LhH0ptWNv7iVxPeZ3hisKT3ve+Ip
G28M193q4QX85hfRBEF/shhPiiX7V7t9HONsIDuFGT0MzQM1MGOn8hkW8JXMINmz33PD0smYvU/n
QOe/pzP7d8TqfQDfda2aALX4zpzuyOvmiY+6gqr6NXq/uXUqwunkseVyA4aiIRM7sYcAKN6N6hu8
cwhwboDp9443rrr6oEa0fHxAaXnEciKeIwbShEE8zowW4if1QVhWr3fawL8YNz8qWzF6Hmg8TNZJ
UScXqsL+Rra+gQwGBP/SgdE6l/KbmU/oLSjXX8DZfh1EC7xaID1vo+wLotlNLDxAAgUjrlLz4xrG
Dj2jn6ipSK7UF3jEP1OmGglIc2wlXk04fE8HdEqA1C+KF4z/nmYvHlHYXjmhZcBojvio77uGTvzH
CYuiZ6CyGGIka1khGqltWyYGlUKDHOoZI61pvfGdUlasFIfg5Fx8C7uOCOFU2QShHNnCmcpF8QBj
rVMAAAqBjveyk8q/0Ya2z5KQBv8XJCx54JMrfVydimuyXXDxwM10UN9NLFM6heZmzsXJlWqZfbEO
4oOX3EoA1V44aVbz9NUfUpOVzROmTMem7thXBFR/3Mc6kyDx0USjgkHzW+n7CxHTLZhClQEfrzrG
QrdKm7ZCScC0MbHYKArqEwvUSZUuuyWogFSfdGkGpeP/Fant/mXqqrr74TPGaIFHlfMrAA+YVbjK
Wtv4cCQATJuNuq14YF/Ythk9xgMqAi2QDh0+wcjDAgHE3djUxQ95ep/9z9jJR6PJmZFUY3E0u/5A
/5+vMPFZAOcCl17+LvG6gAb70Qrq0Py/tDU8+PrxC+KblxwgXnG5iZXwvmrRfWgiPnjHDjkR2jyY
muHlgvcq+as5rAxdANa55s/+as+UvbPraRSf0GjQRXg+qu8oho6+fM32l4rPAtvzJv85tUelEEfD
IiH1V6rQFV503908Oihfl2T0HfYsuGfJaNoTf0KituB67VJiQIbsbdbb4BwN26Lic24UCFwRsByr
3FMtWEbR6XE6IDJdcmrxs8ZhLypfWbVCUCnhZafqhBO6kzl4SeYiojYyLpzu1Vnvo4GTUxKI/3ss
/XfWSjnltTTw3pLVX4pN6M9wPJFj5RDxSxstrAYzM3buBEaxxdpxrEA96y5PXDtS9PV4r7bMcO+4
PE12q9gfYa2qAPCwi3K/UvpUmcJ2mmFj8cKdKCk8aHamfFxzmGMaMRTjvWi5UD7eG7ynTDnQ8fiG
8dAvbJpfyjijdcJ5SxD78ZHTv6sKzB7p+53GxaHwDf26BsmnSZscBhvPae6l/OUNKdk+5pOPjKE8
Y42HQnyfCI9moIyIEUiLu05ypGwpPFfXvb0VyD+cTP1Cf3XPxyT8hGUZvVmAmZAFzPj+jzg9wT+N
bbIeVaBXdfhJHk1jUHEVoeCBKQGwMAqNaq3g9R3/lrBRor3ZDU6HhcUBfoe4JGrqxjh1WmI3jxVv
F+49S2i7Blv6IFvMevrrEs2dHXTZ3v4ViofnGCcCcWrania4wmQlsbCiZbO7Kw51bPt1NYFzXAWB
pmtazwt094+5+MZEJtDONYBZsJR8mB8PL4rkuCdCcFM/EJSxGY7elwqBARd9WceHQ3SQzVWUhNUq
8OAIMlf5pdrCvyVTwIf+DRBh2cNEmrHDJt79KXb/kZN9u158Sab6eQdUDaeqjHAtaNmfrxCPJsUC
XhAzh9F9I8bU1rLh8g+canbw7CuNEOlp+Ks2bsRbI8bSL7zaiyeJZzg/9S87VzWQYF9/Ro8f2t5v
U/qVii5O4caWZI6I2yTawNsCpUlLN4MzB65mZW402YvtKd2q9BdghnVqEmw9xkocly6o97oCgzQY
aqrnbOk1Rwclbl2SDeHMWgmfP+G7mOVptKzefMJdgkwyFW+ro4nNo46ZeUGmTpt8Y0XnAzpZXvmD
aRH8gLviNMzbe5Iw+UFTpCu98KV/QwdnmHRt3SFs6zWZhO4mR6FCDJDuPsr1Um4T+DTQSaLQUPoK
jOiwrtW68u5+5j4sWnCsRtv4d6EruVFjComaMXmb8WOqsr+Z1QajYmOfPT9f7fHkVWBSHd82/RS/
cPAqhFZi0NR1Ejf8agLmlKd6uSsjI54Zd7sSvFcNO0IDXX26aTX9cR/Vn3Hn1LPNaybb9ivHWlnY
bJ5jE/xmhjYiKuXOqWcLZlegSEMYMA846fWjJctMnwgqeG1OkxQpHc7JyGQ3m3ua4AbIF3P3/rR9
HgRD3DmsrX+0v2r4q9CIcfM1SbegGe3fn7A8Meb76Idhcw0KVhkNa6FwSQW75agWIb7AiVJfJTNU
w62zu9NpttaDQgs0lKhyMkHHsPILHO/Y+T41rSOUh9vumcUF5FHuGQc7/YWyBB23tuqFT9ZF4kc0
2ZfMxjAGERr2JSokdyAyspBl/oG/7YOLuHQzhQ1pSaEogCalHJPgvZ1v8GtmaJBQSoJGA9h3A8d6
LLgTn5bz2UlFwJssQHBf/r7t9wtfBwYOoFG+oZ+4urIcEO274TIvMqY4DMykkZ8buqscTvatRfzu
B+BxYQK7VLSEVTDfIbCvr4cG5E5t4WyO30K2vK+zsknXFto4oaf63SoqcFiuuYOefMjN54fP47xy
Z5Dy0mqqTmh15rGJpJqJKbKQ6HImGkUX+E4J7a2i/ZV1yuckwvMe3wm/+TGecvoVANjvGgiRjmZy
mlha45ks0kAYsG1Cgm7Rnq5iazCrpuRH9Ep1UALTq0P3IWKB1po/Qe22+5rxkjrctYES4aAAELAo
Q29m0RsDIzC1fw2cp3VT0mwZ3FimU9wWBxHRURvlNDAOI8l7Qr0lp6wZQLvckuPJyKwlGxkiXL4N
kqi2ejBMcNGgfuroasuaTcFTE6E6xM6iRyhlOADOcsIKeHrIBhiWcZkIafHLQLhyZxWTuw4OloDq
XbXWnyeasexhMR63YTmiwcfOXCrzMYTY4qAMggHZgh+d+qiH0FhQY5ABXEiCtY5ld4L30sHJ5nIl
/n5U2EaT+EWK70Hzmpf/FizPTT5zMmAogyC4Cy2S4vhY/U/fvE/2jm80nTrvCd4l9D+lTDh+sRjz
wEEHvs+FNPd6+z/XIyqy6QZDC9Pnmo2uMY4MOeSvddsJWTh0vHVJ2ecSI8tQzTEO48zdyYhq6xgc
0c5UBfO84KdOGalUY1J0Oy0n/i/JGxjN3wtrXsoag3m+P98JxmcM/JrJOgqnHQ7DAnCBPGQuRbbc
4w6b84Gdp5NwjVICddv68HXh3fjKhr6m+DGRwHEscbuOzhbFOBbF0t6o1kH1etZZAPoF8xSd/biB
hvs/y5o2zOCqp/Wl5ir4yhh7pbvtJ4e1mJrR0ohtuidZKl2JnHcw8NANDLZ5rtNzt2JTV9e0zXcM
Oh8VblRB5YuJUgAUndIV5AqVwp9evlr56L8K+urZwfT+vHVqsb+zDA5iq2X3ZEa4rESRNAJAmRQ2
L+B/drTk9rGCxqsTdhuDoO40ek9vhl+V3LvdXegdFkj2O4FVSX8NoEP4X7jZRSmn0GODA6kK/4Mq
9Y+UUpS58fh6NESlLIlUuFO+jzvb00Hvg3zhHVQZ3/q3dhdpI3IavwQ9BfX2JSv1v4gVNpYxxqD4
bAFObaGmMo61MB0LIbAr749tTZqoNOeNTmfp4PvLwTKLQLoRKEeoiLxuEf8hp5TQ/3/gWtN0IiOx
xvfurNn0lTa9RoyUKJwAbmePS5q8TzgvVlRO3IEQcLb0ddEIfSQ8mnLDyu3krJP2rrP1NWoLSDcn
h2ICZ0TsbInAki9lmcLanDNBlR/Hi8v2mr4pBISmjrmBfUAgFD6Hc3/dVVzxt2qHdeMwP1LFL4Zv
/iQidxd4NLnXpA5eUJDckEPMB0HaAHPOHF+epdflFKGDBeeAfjr0Dqt0utNuHxC4NqnJlG62ev2M
97zE8ro96FR08NmktLyKs52Y/PLfZrYkak+lgK+x+ifBdZtloWuF288uwLDBf+6AwomoOIjl4Y/8
E/5VoBVegvswqwdKj8z3K5EiZR/8FoxezmxiE6SwI2N/rO1apZWs9Nq2iTfeD/NG5jw1xZCE0J6/
U9UZCjZRaykjGuVCkWFjekHyRtTGNA7Kv9PgPxrhiEKlT3Fm4bF3/Py/da89acZjzshaaj5E1ocR
MfWSQKdGjfRatt9p/Ik/F2Ngfg7TQEfMv+b6ogNj4LA+AyqR+omALEszfFecnDejzO84viw4R/ah
wfZVyp+KnWqjfzm+tvuRQ+92mklS/qg6PeDBmZp693AErn/sap8ekDCBSoAUifZWlDS/Bi3k49ai
QRMm3TVCupyJDAgHufYfG4g6exgykypB9vn5xgxf/yvGhv1aZgRu9Thv0/sB2PQA3e1ZaN8bsJMs
fTTmnI8Bh1JlNq4+dQ80CWmxomGwwyguHFof343iTw2T2TXa+TYUdhC+YD5+F2045/MS4t+aFBKz
kieWYCZ/UmJRllvZ4N0ZvmDV1HJFV+pYKFJC0jyCsX5RNHIgWleen0HJO8wgCWF4NrcahDYCTJm2
mEOBd6YshbL6wqK9fYgbm/jdnfkMj/7n4kq5SYEoQkfWGkSVvX1OGOu/ih+pmpNKrBYAsmZsZmBB
beaLZ1GbsVPKSBm+Xkgpux8WSmpj4xi/huh7/qcOlUUj+Nda4vjr5rX1Ewin1f1W+10CW+MoeONM
p4FRZUT1fQNrO3AR5YI10Xt4jgVzBuXphD/wJl3No13kXLtJjjusQkuF/Zh94eeRfMUuxU7SWNBq
dIdlZODXPPYDfOfrhk+GFQ6w8hVcq9s91nzrIZvMXizbYlUM4iEJvIJceS0rFNlWx5ZjyGL7WSCp
br8NxbCoFrncbUB7wjdmKiEMO42dtCIWEgeJLG7p2Bin+vFzwPDtzcmedU7nmNVF2CiNhM9rv7lY
48VON85cWhRXZ1zKwZYL7uy627vjDEndJysowXDgrzp8W+GLyjWZiy4p6h7IN3jl8L+MYBougyQT
itaKvgiSPSO0DRdw7h67UELWsLxhequi6Ie2k5F3LSLXRQ9nmdjlJk+bOoEQ/SEMKI+ERGvjvtqO
KUAeKicdzGCuzJtE7v9k7JO7yI0+ZarP1uWsHvomRWDBpXPLSrK001KNMC/wCmFqKmcW3MWuvS6S
Mb1VHyaHZUYmnrKWNhfsXdgsmpZZE+U5jsaIsJFrFhViJwg0tjNJVvj66r1bK2o5L8dj3a3B8sBd
gb4ynOkESFIK13NmCVj0wcl0i8T2j4Ndf57YSa+lXo1eUrITTsNZkj8EWBdlAfMYX1zfhsXPAQ2n
2ywsCpp1IpB4nuf1v2NXNt2RieqarBxy3j8dRwef8dhT/tF5/ZaH4GN3z8jjceItG5wKUh/UpXiA
yGBfsf8eNcZ1yzcv/hfuMT6/niDSnaVoDwceCWoZOF7YAI2gru4REmY5HkRAOOLkVOgTa/YqZOMQ
lvZ7vX9Y6oKBU/nFuD23DxgXJ3hS95le0wN+3ReifVQCFDTeeCHAl1z+khOX/7ft/Uz/V8t6x2AN
AOCwN5kvNMZVxT0sFO/QP0bwC7uScGrVKK7pWaN8VG/VbJcEV9XnhGyVf+RtZREJvszJnkiUkWlO
uAUf7P7FABXK+ikDyXUUHqYFT3uo9xNaRDhkHq9u0ds9Qmm9DwsM1GYUTO627M8h36v7wysHyYkZ
9/zOXM7Mznd5Oo0bPj2LTB7Wsf6dHgbEW65KVtct415/BCYh42KwCbDttldrHNM9/zu06qLogY0/
ieSImIYtyiD5Iq7SVjCACG2WrKha5Yf8x5PWYto6IKnAdYUkBLx/jgouxK1K9tJBg4khlUZdasjW
F/84jNLITapi9hHNbJwKYt6Bv4ZmRSs6lQJm2Xd2B8lPZbI+CjtEvYuDxOSgyIAGCnmT7yDx1o+b
pPfZObkIcPiVFyjsOmakCs6gn4Itu4yKJ3Yekww4gDt+cJXHnmmQ6gXtmpZM14r68EUXkvSvfgm3
SDBkJas1jamPS+a+MZToJR84Z497DXpx/OliRoxiBiVM+koDv8s9dNb9lR2UcZhI3tWr0EyrKxGR
gyAv/Q3D3yi03+hovFsQboIxZ906jrBmYdzwGe6ODOujaquFLXaTqb4PAgBiemFHzr/BJ7sYyC3x
F+ttrPYXD8nlfpZzPvPGybOEVfrLlb12xiMSFavsAvJZiruWhPzFbSQ0zKFmBd8xTi00X66bW/ik
wv+L76rFomfCKLJLiP85iqHBD7ha2VBtpPi6X8rwVi+NMeWVLv+aMt+FAlNrE45CZrr/RpAjiFN1
Qh4WgfAahkiAnsz2wOSpGyKs4Tep+LqNyEl/CO+HqZGGR1WMelAXINSiFJ++eDUQQ1QS6rBY4PVH
AC7vqAEQssO27Xyj/yYYGnphc7WPilYAhqkpCtKjIE4dvrGelVxUpGHaPn2raeO7/HsJlhG+Hnvl
XxUqnvfh8xxMRqIy81K9/oSdIoFQ0sRhiKmJX1PPfkdoCCCtf+IpNvpxXZ9o/K46Gu+m+aNS1Nxu
6ahiLUhjD5K5ys4iC4UuyAWQYcTZBH1+M4m0fwoqZkd/qgPmLKtDd/+O5C2B/2gQxPT/NTUTlb1A
QSg8dQxGkY0kcORto9dPkPWfej9s0unuvWA90r9twoVin6cHZeIPg+QrDootek8J1n7u+v08On2C
EvL4D5iME8FTFmZSCkDhHbC0i0lGfJyn4P7CEGzBU7/3m+1k4DTBJ9E+J7QX1bxZfkoixSctAYJ1
n7PiToFACYYOnM3J9Q5mNLY0aZVNp1/GLmVNxDFVsUGEWpR+dCyiM2akyB+5aJ1wRC2UioQaQ79W
aVrV0GJmuq1f5atr4XDzPe43Msx4Su2Mj4oOmmKWFffQsJoQkfe4Lr3TcF95MRpRgi7FX6C0xus5
qdNizYc91FJbHlqUFcWW/Jz6ZNDbS6VH+3MZIZ5z7nemlYC3P1pvVCbXkdJMsXfjx8b1luc79UHR
OuYE9qoBCvZAf3jxWOShe5sj6ZQg3jwhrAyawItg5WFlfECQMLTkitkkLTuxS/HUZYi3O1Rssbfx
DwqBLS4ruDICrRw9xdvf+BP2pEI2cB9Mm3tpMzOngIQkqqyu4mlf/lYViIKKxIvC6r0qlYAnfYk4
kbBDB4Z9yAESRQjTSM2ZxT8hecbR6thiOSaAwdUTuuORFQgmPtyPNs/sCPVXYrxsmYme5hXj6x0W
T8ODpC4DqTULFEj3gIhCGiLEzWifY63QRtLr/1PWcUblz015qyE0SLudcPQHB5J95vw8oKGRTdur
ic7acuYYmvhvZiWsW1ydBI9AMc+gJcSBEqWq6S7i1KKsyxoerYI+HyVbRNZ3+kqDI4FpCVnCVI2A
WPUt2r5UnTYczsUJ2+9s2cMt4QHYXU+9bC4b6WYam3md0sVfYuzwk4OGjT9G56Rfm25wFeVjKTJS
arjmo9bpPAbP+OgEItRF+gHgfLhspijzCe+4pNke+lddB2htf5HtHop5d4Ez/ZfVvI0leKGwV6PC
48RAkstwFCrxhK5YvxcxUc3r7lAx51dVXwi5ACZaGTsMxfLrwbFN6obGF4iusOJc4Lx97FJlNg+j
sVtQnlGAdI44zuUu5heZVPuJ59wV8PkmNAyh/+AijnUoghYTQ6kEdefAbgOc6HlLOEKv/Rbr08RG
Pz4cMQUdXDTCJwayUPTapwsdX1xQytBFNvcxm/H1IgAbQ02vOzS5Se+AtHp+JhkSapU2GleBWdMg
XTOsdrhLt6UL+BNguaylYZrUAbt8mQvyfmrXGIgtTDoEC7hNhbu9boU4v2iEslCY4jiLBxrGaS3n
ey3tjujZz4n36l4A8xxcX6147fqBUQu258rwkjZMBYCQ62e7DbocCy6o+8GhpH7ygDfqngi+YSTb
SzIac/WKmCN+GSbBgjANxI/hG9bvumXYYc11kRNns7mzdtIVJoJ7MyOT1T2LYl0yN2TqrqcAbe2W
NUgCoXQX9jOW8gMp5Uz/AJ+fR7+9Nm57VOfQVbCKw54PDbqRy05kyBX0yBOuI+4/6ji7+bpDggOh
HJOmUSeHB4rrBWcBpF1R9FWvYtn1sFugRW1q6sGnCuIcKQkZ8xJzrfFyhLycHGu9Oj0brh0OdU4/
kRymiDZjijwsH3IPu3busL3lG3pAlHosHOptKXHn5LZJXUo+t/OejtG1U/8XpOrNgLsjA3HUyRrW
MT7MMOKKI4/b4ShxhdRPJHoMXz+QXhaq+Vasx3VIEd4MD5XGU+p+Jx8Ip475f2kgIhApWMnYu5DD
pSXX4Kys1UkeE4e+sId4aZwI/9gxFNnR+g0/CQCqpnv+wZW/euB9lBLOjj3anon0BG4DKUCQKWYC
xT4pwZLbYD56Kgjp9WALY+uaAyXKAuc+5TuZpumVRcsDBC0x4Q5s+pWqdYu/qt9XT4WgoUFrOOQ+
OBm8IS89WHxPAh6bQZHYR4xDyhDZjoSd0WdyMpW5s0SJwnBTbvQmMSdUZ3hWJj0Y5fp0oxRyNmRr
wBrCyrTD9e87rsZeg7/yUs9T/ju8hc+E1SNqpbtJOWv3dc2D7Fja1aC0ZtY1hCcGxiPAZ9whkfYB
o8nFDpBGYmMWMDQnVadTtBs0zntGK41yKngy8S+P63lzoQ4Eo98XQ9XNXrCYYNgd2JquMnhvbHex
g/sY9xSDqYxwa1PhpHRx/8LLw1w/0qFzQXQW3QF+lt0L2U8CqR/I7Gxl6c2a8NaOHaTdaOE/nhWR
x76uNi3yLDEZrC5cqIQvl5OE+80/bY38c0mlL+1xRr63JiMD4qjbD22u7iCh7d0CfU3ZbkIJ3HgE
pmE4iiHnwzhJlbiJIeNH+y04tro+0DthyGSIQqnuN/+OtZuhyECMc0meBMfMqsA4fsivPlghoulx
TTRCAS91v4oSFkXhDTPpw+e0x4GXlQZkJmeBfxws/9Iya1DbsERUu4M/Qr7WhZSjI0dTc+xy6vWx
pMvLSOCkf1aYkFDZ4Tz2dy2+UZgiAkzjMjvD3eOFYfpHBBQJtPvjPzfS93ZWQRrWNfncsVj1BWP5
jVxnsaaU4pN7YaYNEDHvPnThDYA/yCSOOGcIn1XDUL0SjeB8P7kdrrPwh6W1YeYi0vs3iFMsBzmw
BfXoHITcYVuFDp1XrGO3bjyDcY+PHM1WxDeSP6lU3U6CsakecCvjG2LADKDrs9ySUXwuxQpyk8DT
UqPHLH7FL4xqCu5PxHxXLpN5+LDb+TQry6DHEv4wojO1APoPFCgcdHbb/Jt2vhuJUs7M20zZ2YZO
zocPKr5OUd13jfdVniovzJ9FnT7aXB/P7d/9ynGs3Fcbg3A10qU3mGY4AF5kUSjMFUh2scNTi2J3
7lghY5ms0tajA/CCPl4X0hqbJDQsqt8zn1kYpjhG3TYaHw63SqMs5W4YKIAJ49Y6N6OEJZnv4Z19
+1zffbbEf9XRvmNnmXWXFGPAylm0ZHnWv3oIG476E8LwPSfT82demZCf9M+rJieNr3ZcIKFZ9yik
cJt1qhjVziS0itiSNe5u6lSf8rLcYXEigmI5PoP3ZaT4GHlWoamIx4eOfg/OnLELETLTWdXMG/xw
Iwx5kO/fJw2ibjdGCZ0+wq0b3CJ9cK55sStvuL2GLPm4tVRiksMNURB+D3CuL/8oR/DX8HAYisZs
+Rm1ftlsEBwpJis3O+TlQ/OQvMmIRVUKgMXbgJPkbWGVuIn84oAult67Y/GEzb8betfFmq7rJ/bd
4XvXARzQZ5Fb69JOQ/iowJtmyNiPKhB8lfP1AVtO+XVPs5/jTsWNG7XTxzZUwQ56ouCL+YF/2f2y
VYMW+fOZtC0NzSuvMav8iMmV2Vz9TKie6KcBXIcERrinlBksEKuwhHW+IDNF2IKWSEI2h4P5kv8I
9MDu9wcQ2ErfBpnPh8iOGVTsDJpG0HRxXDMfVgdnqZzs5dTuEZVXxvZln5b+qmcI9CzrJvfID9HX
WpRnoBni+brwagLleDc8gPHeSxvrNMVclFJpWi1HLz9jFDin4i3T6C9I6hkqEH4819ftSu21QHB6
mJldjkNkPPOZr1rgnvcQOPLsanvtWaFvinhlFyduyDhNkOKKq7za9luctcaH4slhyZ6Qsbh19B4e
S4/ZNpOsocH9xU7J4LTSnILeTS1JXJQBzzfHXEwhoPiJVDu19h1JYy1XN8eaN3R/QVsyyFL4A9e3
szEIop8NEXq1TeM+HpBv53lmdyO09yEvMvzNYIk0yZQKVr5tvBsVe1RntyRDy5r9mgqo5uX8dNzl
pV8Wh8wSpEGnIzYbkiGp+z0qaSUtFqvwwXtTcSvWtDLHYFYSOX/k3AFdZkcHLcO0F9LebdXkcc4s
s1Aq4dUXlQy4Z7YY7yvHG5pTsHLHLwGrjFmcmtfv2N26yeJH0iz//3H8drMvXLOu06xchzEI71GH
34A3rUXfodiFFuC4N4C/4rXNRa+Evr0ASXwuQ93bi7RuF0yItE28Ceg4p/VMYq1ntonB0rqvnE2Q
9iqXEMrCZbCyg5qI9R/4wcsMgigEk6rIbHe5jikuOtm5be1KWtMvQyJplj9dM4smajQ8CzM12fMD
oCvPjbPeX7RF3RPyDB19WMpJihtDIg42VNM+dRynD7ICtqxDRvtlrSC9VatXMf9DlbgDAF/JHHed
kP9I7SjBPh7T312jCrt+bS9sGtYTDOrRum+CoYoFxwfLMXpOsxsupZr6d4GZSMZxSk1JM6zOI6PX
/e+JUf/rWMpo+Ew7rDl1QQqH2/dTLSGdhdaSxstWiSVPekkLoUys5I56aOBmghEDLlRl/hFIue0p
4BiwAUvLf/RRsCHDvtkPn219Q84cmrwTuozFXrT39tFeJabXLPx0xauKjO0fWTCsOauR4jI++m6K
Go+sqZno+3oSFzw4ozlpTwl3KGZtXZ5SA0QXPpL/Rcsw8eox+OQFZ6mgHN6crc3nys8ZqcpwoWWn
7PSeUbTzH1bRKqquzWgsl/8qQ6VbuXb23DWAkXojIj5IJIFr8RLiASnWpZiXQ39Fu2fYHAcy6fUa
64mQMeC9wPpewECFgVXG/D8NWMvlRlDacU6t7yqlcrh4sa6d2M61bbnRsPPJDNrieGzxfOrOKUZY
S1EBXfCi/s1s4hb/4zMl8QFKUJq3ca7Y+42EK1baiwXAlKFxjS9e9kHZnjjJQAt6prPEJl+0EhRW
UXr8yMOetk34S74kr0+V5bFp+tMBbobeupKNzyW+/F32Pz9sXpmm7fdQaRxw4aS3Bl7Luww9zqUR
n6GhxuPjGu/VXVeS4VLXvcrybMunZkpDZtK8YLx9rL81BIQ738beYkQZEFW5tui2uf2f64EvJLm4
TJ5k4KYxsCc81EdpxeTmq1IB1eAnKn6CzwK8DjPk2nVOQUB15tgrdxqkm0nItN3HuyMAvUxZhrAJ
vv0oMbZLXmuymMf/fRkbL3rLDIh1IPExdIlUP0k8GRSrEaEzlQJq3vJOPBCFz+rYbsXx8OzgNM/E
TYDpXDProEmz1OINAkjwHMsZZ1Uz8WQ4RzZnj9OWfqIewBfR37UbT4v0DHQkBuKlpylwuWe6U8T+
895oDmmLoGB/SzIwPjNb2XRX8CcnH3If2oUIB51+gPjRRGdvHS1UtyWAqu9fxPJhzIT5GUpXOzgX
8pWWeO44rUT8QAvEvsxuiSHocuxJjNSf2KMX+K+bplIT/SGTRV9fs1InqgxMGhq+2nHqpe+TqNT2
Xyqc3S57dxb1a70hDtj5223XxWsu7fK7eR0PuIyr0N9Eaj+nK2Po8DD9QRxEQPbunGbzInqV8xds
yTUqLFYX9EgTOGfLLmCBunaYtV0sxLw3UgPm56/bgMPQpYRS6TtOo5daV1RD6GQZCWLdp7BTLNid
rZY8KzLpFalUt7jcL64/wbdzqB+EX0TNP3vniMsCiZr1dMkVNFIEqatmTRKOU/Zcdi5C113yDjhY
RX2DJ8PfCilxs2esfIoLyopVtS3xZuArTTUJ8E3YHyCkdQlDPVuXXzHpaBnnouckIACn0BonLDig
MrrZ1x0COos85+AvTTUhODHHdJJFXfVZTSXBpbaR+fHJ+cl9abDF5fb0PKZwnbjiWwtSe5UK+1Cu
AK72uBJO1TxEFrDoWxvY0KbOJdE9vR4V5jBmmgRCQ/fqQc0W6Q8Rucu6KYjpGueI2HugP5ejnmNF
2+ir5pOBcGSt6ViKaPRzOfo+LxtrQwCgrCEJDh1JIfiBrTpDtwMJD8LP3FNPKmgsYYSqEWuKD4zb
KC2Ni6znOFhfb2+eVWiY/Jfx+YMJOvNAa6bncteXwa+kqY/AdgkBbfPZZQa0jiN96EVY0h7TcWSW
12WWA4ho0tl2YcWLwwxAIVhPShaJ1+Obmo6bHU+grBQ8xUhnVT5HWXgy8uiPDTxrOhxioQRhfQVD
W14v3zVhVkTUPMBLrF4mWlw6MVtSHX8tbYEscHa2oTQQVqZgvFA4MnxD7dQk3dmeorqeSS2S/iHy
UJY9dn+5pSl5YZmjf+Z2tswSNYyNYHnYZzx/59RSTHZl7yOMT6ttIGC+viw/wbWwrR6mOFuPKhfS
S135+rsTwjdL3yTQNd1IML/8Ewiy1RYiKxr+m/loh3id/NqSmqvFJg2N2A6BGi3qVZuI5QFFSfL+
9tvsBPT4PZJ05znQr3rVCUvsrSrr1Jc0X7U/f80VmmwZ7DcU5ihBMO9xKgdalAEd6P5qYPGXVsRg
i55hwvKjngmaKzY1lKBQTxsjgaQGng2REv4Vv6awMsFABWKcPMUTApgaUSS0BYdqJijSHrN/DhSZ
jsVvlHhjO1/sMO4X4vly8K58NCkrlgJyFY1vHmwFHjr+q/Z+AnmPWItndzVdPB1Vz68cHdKOSdiv
AtP0YGCJu/OmR1sIcD8ymeF9CMGWnvyBDQ12walKDG2Z0pg90bGRBwDKl0RyKt3xEkB90eddz4Ou
YhU0zkHPEStlmt3XU+rSaACgCG67QxoNN/IoJSiyyX8FhPBPiMrB6ausiWFuSlVG21lciW2/2k5l
eadvycxPy7f0kvE5EKZo4O0XQINb02J63Wrdm29Wsbr7PpYmTVAIuSBMFNK1Kae+GMANMS11GRUh
dynbSPDw7FCLRuDBZjGASNBiaChdBqI511RiEqiyNizu8MTv0lqyU0iQVDJhQWUCqNZB18crVyl/
3ZHYsdqV6JriF09mBoGbRD5DGXbc8fWGo+rLS4ZRfuxIDpTc2aAr4DIV6DYou8hjwFk3c5saqR4u
xHtr+B2QRAXgbbiJcLHiRjFQqTI8pa1jA/sN5I+WPeXkSXHENEEN3gNj2FyNY97RnUkEOazqp3UY
eOtMPfrFDUoT444HMiw78dJIJm526xdkrDhF2bdkuxz1oNJQDtNqfoHiZrqY97Dlu4iX+miJfV0H
zi74uC+WAbqZY0NG6CSB7ggo2teqm2rHO8VbGaBACgVh5kJcZsbYt5ycs9keFOyvlY8xjgVDj0+m
TFq3WChRhycuqW28HUbKapQeGY8ihwfpiz3ytJqGvcAn/iwIXoe7RqfNetefvDY4HoTaXvoet/8/
y8O32Vfeh0PEJjxxmtBkoQitSHczUckhDqIc/TnIqijaA1ZPrIdhHGlGLJL+4dbm2E6AmjiWs2Ev
o4lqtqs9P0eRF3NMifQjyp/nbwRnvvo5L3Xh/SY0q9tEoayuv8nPDPf4mRfpqU2DzkNQLFPSVhEM
SwTtp9m2gkH1eDOQiH/BPIZNUoDw0yrek1oINY6zOXD58Q0YX7lTE9htvAtx5loHOqzpkQkGFVMB
tXzsx8/gMbf7dMjrlcJI4FBeOvCxS7dOXdMeAbG1vqvjAU4C7GiEozqkL+44z/rwueP90YCphgbS
RCXEF/hJNmUTjn8BilTlbR8Bjsi5nGpWUp/9JF1T0P2W8KxEngGWkhcM0tyQ/8GZBub84dEKxRR4
78w/qpSyM6/S3uj6JebhvHrkk5bhgyc/Im6JNOmGodwV6jScWkzdKA3hshlkOy9osTX+SyhExPIv
PAqc+UU678to5iBAu8qiJ9YOYwzaj+UATZ8J19AGa+vcL3u/zM0K4Aaw3ZMq8BT1hnCg5Nn0RTZn
gnNHXXKPBkLSKNiA+PB1Mmod/fAcIRJRPW/4Z24PEj3WqJaY8WEqoQiXzcw2qrJ/xe180qRLRI42
uDCfrquJIrYp3gyTRPEOJwijymdvZvSGiwCoMCruzdriiIYqYcFF9fCkgW6ZerYU3ZZts1iDLS72
Cz3T/1JrHrlqUkKhnBEQi54YxpNA2UmSFqwUz+F7680cfYL6zG37+mPO9J1GZnTCAxcmXRIY78+7
NvxjjoaZe7pmw+dij5cRSwOT8l+Wq/p4Kh+3AP03Dna+ts5b/czpbyIjChYTaYs1nD28jv56sNCs
NBz6wO0uaLI491YanDiPkqwO4Vxz50ZMVoxBiYRkB1cUAnxRCZQx6Cs23uDwF9g8T9WSiOH3gcq6
XucBE+jQAQgjB368yrMZdlmJpb1epz1bSl21+xZpJpe43WqccO+9CAMbjxrhwCq56FrG6bWc8e8B
qeX8tdXHgHlRXuXdA5VgR5JDQWGI53k40dzhIuj2ZDVLIbkvxWc5hxHrGC1k1r6wXI/9MkygwtlY
fMq3iR601i20475iXYKXfUYowYfYOzaTMxQRgnsd+aqzVQpLCy8pgZM/T0EAS6nMxvzRrPp9zpcG
oCVE+qXvQMQ7s+R6hu8LGPsocC2OlbJ1gcTLPCyiDaZwaWH7A6FTygLRYQA8NdfR/ZkMuvWYaIEj
NDHx8jiDFbCQ6OqOI8bXWqwAMOk2bd5Q6zbTaSasQpKTLcLqde9VpKbGN1HUvlUDyLcCnUakmq0M
qT05GGmaMHxbQ+Qj2g6tQiAkrwQ41YJOQFHUEEQsj5Amor25gHdP2iRk3E2hnbu42/gUlJywhNru
Kui0/D2c0OZRyplEtdHhNk3paGtePwOpDrpACNp4StD1zBQmAJzSsTrmDkraru++v2D0Byr4eZfA
zbRo/HB6tUjxzwbmPCy4ib8AufGGDyVW8XT3Dk+MRHnG59jD+rLqMXFGl0CfHFjc/xC8hfcI4kNB
ttdl/8zH7+N7Ue7CY5lzxWT0NvXCh4ScwCAQNj2YpVaFGYQnIM269o4YdcsBSBKvgclU9GgJkO/i
O7g9YJ5cGerbu1VvITUxIm+Engtih/MaRsupwnUT9trsqraLCqmH60H3bU5bec1wJsBh9JFjvoai
ZQpmW5jCz1vQ2+XO1AC14e17KR1oVVJbbO/JIzEZVPtK9rUilI26hpET4/c9hmR/xAoQ+7P41QeL
L/T1QwcWLwXI+AMzbVRo5pljJkjhT2ML9jvy/nPGz2S0WBnV4eYxtYTrfotJBdOy0bhDC8kyM5hi
UtiInIqevFZpa355ssLoFb7r5uUMuZNeoKXpMJAvtO2uiAtOo5kxsU1vCiZmW69TJVai46rNjl3Y
Vh41TtrMkJ9lfV45PxTxWg3vTZkLox4N7/Jo40064cUARH7uQ8ibZNyJ7nhwppJeir1qrd09tKEM
U2lLmhpIjBSYSamYh+I1w/M9qKvo/vgXFLd7IQ9qOd/y74SSFlZaw9zrmphM1WpglPt92T1YP/OL
V3bM+viNDuFYLiyIZYPdPcUqH2LUxlRKjarVAde6YwFz7i+0q65mSqFMZ6apjV9tfIg61Kr1Sqg7
m7by14i8nM+PEij2Q0jZHrkZhv2iwkp2jbbewlu2eqXqmUQlF7GZy8FXWSEOuiuBr0SBR1Qx9Hr9
KHfLH+TECbKlgghh5pHaiLSpzJ16XM4GnMiKyhAzIRuyYwWal4p/aLlYpTnaumZf6WEDPJhhd9to
l4S4MOkWhrgpUx5ZMHwVHzGphKa911subqqPPWZsCzxTBrzh1nnpY/GnzImnJPu2v6MIcmJiLN1v
TDh3z346Z3DFMXpLjomtP/6CvCphDuXdhbsuePUhnMFqr7W1Xfn79hLSWJaQD1ZAw7Ie3WKdE8HV
3kFnHeInryCdXpflLF7oSgdDeSUdIU5hJMBy3+XxJxXydx3emtfqJ772NTaaeldP8b8YYn/GJV11
RCrsi6y16a6GO+F7daXgyWWRrClxOfHv77AS+QJuAqqlN92TEZRhu7sGJFnu4AVK1aMQJhW4tZby
4amHJK2IRb2fmDiEYgcaKqBd3Jg8qPMYKiMbX4GQ246D03RErWDhgonJWTs9xt3V68mNZkvsWKAn
hp/Y10M7Tlv8cPHSBrIoO6HwlRiIkpg6uM6gzKa5UMq1j7ymll+v6P3HWN5fEXRfx/5Fgd90+u5N
rJTF/GmGFZ0J7Pa+QwzyGtVq7HXXLZZn8+JiNSRS30T+Y+uh4j13/4ZFb9ThgtWA6FSjSmF6riz5
8he+PchjDRROJsA1xBIDEn8wOZdk7e3WCSr+nn9CE1GQFNHXKDsz2iaZC8+8Yz/ac4amljv8SyQv
vWHvP0xC3IUhpxVPHMmmXYbUKvRXeFn1wSQNpKwTWOHCxj/MIFcFW2VjU9lTDkBNIXfvPW23xkdE
NMrdzMVewQo+T/39npib5F7CGq2P75gplWRg2y3/k67/eC2qz5MhtMzQdjOvgQx9sXcXc+lsB2X3
kbXgZOrMZRNNMmh7dov9omu7lnYGrOewsGB+dpLNjWAupPE56FrkBIZqzzG13tsnwWRVSoLpU/nq
ubLSOSxRhRfe/smn5EIzxJZBs8T3mscF12P+Ibk5PIBsq1z6I+FZ5yrVo+VZSfUj+fOC2N7i00qE
5tf+sSDZ9GYtUDdxQZ5KBLD/Mn+gKGAZtNcuAg0kSgp+og2G8pNe9/fooDZAHqQSNolWEUJeO/JI
YJEXv7UJ9MwVjTDI5ec29+6Cb/3MR4Ygox5X0J84YyMYt0SCyy4G0i5sKV79dxLcb0NnpfdcTkF6
uLy7MiTBAlFy1lh8i/Sy8D6olearQVkxQJKX3kyBpAanYHf3QiYOI5PzioWZ9cte7SeA5FmJSh3C
+uJiUvNdkI86Qnr/XET+6rmQOCJyr21IrPHg5DehiwNAWOKxjw+IGGYWvwv6LIJSvcbFsKNjFF4s
hN/3GzJMg2xg7yUm6O+D87BD138DKs07yPt1gFKJUK3iHs+jLAmai4ldnJPul5uEqPIed63VBcx9
h9i18suY/tBBqKBnPN4AKjrzu7Z6smUU4xlHNuECRVKQineNsE79u/ofrF3x77OjRwH8wThHpe2S
/lx7umNIs6WD2xoHFZ0ZNm/wiqQpsJGoUaPacJhMXdYHSJpt1b0p1pH45iCESeQRWppS8IcsO54A
MpZAGZZwzBaS3rf5Ex8VJBreLzMJGqL1VhCTeQh60tbOxj52gwzCKgrga8k6N8L1xr2Z1hN3Czwd
rBx0ZZ183Yj+AIR3shpFqL0tE58fOg1wmw7QVIMLAJbqerOwTMlgVgNkKBbnYgYntgcLsNSpcMux
HuSvMaA8qZArWJ9b+T/QkaphadRSaxIQF9n3O6EmOrxGxQD9Jb1WEJCReomubnMFZ5S8pbVNblux
opUBHHZgMsNsJdO51DqpT9S/6zGsbqvrPArd4VW/DzhF/RSoW3g1FA7eyW9HlgNjugurkZ56Hi+F
4bfHPBkRCJb3lDaWnXw+gIJDu5WdtlJVK26U6GsATE+IXRTGitIO8MD/3q3Wm53GlTLL93dsiUO0
ZoAFVrT7RRs0TDHOML5+i4t65tSjRE/nMyicEKVjdBaAgvOrnqIO/KrSnzYsNfN1vb6ou6SVgpDy
AUQTOgeGxThBdyO26s4dpXsrUsprAhqERCIFS9z570XS3Ccu9Gi6JdKHnuO0B+zka2p3wY77QH16
pizy0ysIF59ibsvPEcKmJKhJcsnbx3DJUNKtpbyqC48IiEYbOOZ7SuvuVuzEhI42C+2GA6YzsMlZ
l+iOMmsz4ZtkvC7aVr2UoG7swwwIbYoLmmLfOLZ0z5Al72JzdnQ2ihCOkk3lIc4Ah7lpRroZTVab
OmNbAiaqhUKZQEZVi1oWasRNcMEPX6M4LdIb59fn0ZH26RqTI3vTDuNngr7XpeeoccbVpbuNnTBG
LQgm3ml/j9VIGDjpKHvMayP624Hgs5LNLQHdbe9Up2YkPmrkTTdrhiCHjZOvv+qygh1EdavEwnhI
k0QhFIvfJHgQMU3Zqt8eeF2gdeu+EVWTuA6sblnj74O+eWB6RS5TvuXquMJr6ggCE58N8a5ZS+Lx
5tyjecLkVpigVuYD1fqvdzdtstHI/xNwQgVPRcH9VSs1T0H7pB5HQ3q6//BhEGCwIIwffyXoyhCR
cSNdBQyAg3BkSqGxv/40nFeyhVTkAPT8knoPJN/J4vA81j/r6Du0XBTSHm7TuELHlVC5ULUDnoaz
n37x7c32WzFdbnlLzXfVCctgZlyza+PwU03ewGDxqGGjulKJj1UcCs85XX/0sC0Q38hkOsG8YXRH
ZmntnbiDBh8CZOZJCWm70kAX/siwTQFQT7S3lYxJ4n14OikysLw02lqq0zLkgK5HnvnZHVzXfWZV
R0QkupkrKmDSN3kR4aP2H5Bnz1tW4Foo3KyeFSAO4MT1XAp3ICFaMdU/wjGl38bThTkD4SNp+LLB
n3+KRjwGnP5yTFjkxzyF0zWHJgv6htBSfz/dpC4JQ7lNiGv+D2dsLH2s0o/9EohDu8mNzEPx5Xqg
2T3CUkRROVr4lIj8IChxCdgWLDCK9p9bFrh7NuYMxlxd4KWu3ztfpZICV+L790wFvC8OdNwas6n4
fqTuzHqq9vrhFy23DqAfEuj28lVAOOukhWkKhDSdUqPi4V05SoqOLCtkFayGbJ9e7nKZsjuU14YE
poldUXLtTH6Qrk5G5WYJJ+ybmXg2BDn40s0NEG4zEyFYokvkMnH91vNx4aMd594k24SH8rXQ8MaB
0MOypNdYEIDrzs56erppva3Ko8YF/13Gng/DuuL9q7oE8rCzWESnjHLnQaog6t0yRdWlmnpqeste
GgjH8uJohLTdmdt4UQMrw4Qn8KBoB98Z8cElYJo33RKw38IjfF5EcGjK2iIr/mxjPdf+gBXlz0gw
F6r/LK4sipxCpVGx3rYTuZyK0Ge/GQKiB4Tn/YArDODrDXBogoztLg3lrXjfD3toIZ5Y1xpix2UJ
+0U9j2ROpmAQDd7kiHpW3TZai6uTjdFDdw1IemJUGoO2VnGjDpaG0XQlGjfmqzgpcf9BGYtAGbmd
lQ67cuE+2WP9tNLMuI4hMsUiFRpYmAkiGhmEu6gtmQ8GhV3jT+KfuYjr20QiCBCWq4qWeWB+GI0g
mI7bsFHMVNN9Ptoexs0vL8HyQfTF2dg6GdKtSxv7qtZcOeuYJsabClTsiztnQTRNpw3v+oRlIuk4
DXy1WYeXr+gxeQazEDCBmcgW3ZPwQ54/irolNM9eP8W2d8h9JVaiSo2jHvYxMJ4naCuBrO6RtnGX
jNodtiRsQu1u+msDsFS9AlqK0ghwgxkhGh6i/fXP7A1te9jJKgh+6qqNy5J1uGSMmQzesUMC1SMl
ZiYnU1XEXkEVhu3oEXN3vPLJf64vUfOp078mIe2UjuBC1n1v+3Y9bul0sZB9Ry2ccX7jpZPHB9nX
90TCf7mOP98lAvit27dhYw+nTxaVFolLqyvKVlgwM2Qw9tIH4dEg+sJv2EHXJNIniwXukSN3rubL
mJPoHW7E2yj844ELOL74UJ19bJoT/Jeg0PoFG0/NAKA5pjBB9MV18CH+cQzwbfz/UitRZRaFJFAL
0gEySsj0kK3HdJ2qAm+gnVP8YCnQ/ldI6bEgMb2ZrDDHTZ2JYzaXhOLS74iyJyzTGyRj2MouKu8d
Uo9x0sxsOEOfBkmqsAfpsPLlPyT0gXRXi+XL5gZMy325gRlVu/aRSFuA1SsB3ZIs3KcZtwHLaS+e
glgpvLyTwIRsCeV5/YlI3HjO8LchsoEX+caA18DeT/vl1fOs831r0nymTvaQidEJ16Q/OQCjs9Ve
OUxHTde19xE4/MyR5oUOqEdFpC0PaKrkG+0ln/zdCIWuYIaEWBWztOvIOvCe47wA5iZydGDjt3n5
JmFXkWJVoMxi2FiVwk15U9xswNwFtxSh/QoGIdj/1sE9UglGTXaOxVqw1dajwhDEBBgKXZcRbNGD
LUCU58FadpKcUtj1GpFiW+H3QvA1zwD1HbCWa3VU+8Rb01Wd+okRo/DA16FLTZZ99fSsZoEPodTN
cDENuyUjHL6Do6yeBh780O62JJJQ0zQqlSRhcIhf7C/Nj3iGZfwSpmINghm4k3QlEYfXrmc9ZPr4
iWTpZ9AlEYfAci3OzRh/bSb1nQy0Y7LQrxsA/PvJnzKKQmuOJmFEHcoKTJN33HFQAopb3PFnkK8X
TJtTuHweZgSz4H39LnvTYlRpsl6hg4+wJH2vlLGCYNsNQh8PupgGJSpaiWEFK9EoTjfPRgiMIAva
6WNqUwsY7CJKEDIVDp9Onl5VTw9t2uByrmoVDnWnqdFf6baXyan0uJvtX/jZQyMmw6D3HY2zI0Wl
e68W2tihwkRp0WQ+zrUznUaxwyTNiG1JqHE9+TVDpNV9f80bsmWd7y7OE7s4QEREcZN/10kroqDS
hhqv2X2jkgbfrTR4cuhkeut6FIb+SbVC8SnOGJKM8wYv2yKBonwX+VVYbrC2AGcJUErtw/6oHWYC
Exv2wiGEvBOCgm7CVvaC/HOXPS51gEJErZ6cNEvrrzP//+Rf5YAhCo2VVIN2fMmUuFNUhNx/ss4T
jviXGVa2mkArQ3tHW5/LdemAPBsJBl08ijVymLe/QLKyAJKHhm6YahJ9qcg3tyDjQVtxb0H7Uivc
Sqngyf2JsT3i0GjPY+c+UHkgnSgvJMTznQUZ58nBW4Tl/jo6jRYfLkoZFfroQnki8L/Mbo86bgvz
WjJzDLVtWTPe/4RSIZAQKHSY2WP8EAEp5YtY3oHgK/Kgqv4XFaHqflYSe28ZAfC9PYw5iJvqXjMg
KN57vSAJ4h19RyxcJB1LzYpIglD/ixcpkaHYrej4hvvf+venBPVyM/+p6Ekq7XgHCmm8Rjs7ciFX
eeH9lz9/pIZYxmnFd0xlFxTAGnmr/WtP0QxB2Z7lneTiQ8e4YwG9rK4U+7cExcub0jSiaRtvwZLV
HU+/hwQYRKXTukFhikj6v02N6d8EtQ9farpD3pakxjYpXJtE+vNPQs4P2n9gtmK6FEJdQZqEqKgA
9mYm77R6/g5P2JxgCfjemLB/NExW90OVcq0lJhd27r6cGvaC1zL6Zjg6+/cU2yP073YLHsHua4T0
MpN0IOjpqYU24ou6MEietw/mEoIyBClb1KOkphq2yQsbuqbhWwN5TD+n7XlTpk1lLqmRSS2WTln1
ysOSLkwbcNdvPIGv2FP0ka09E9mshcvUmou3jHT+YipHCK50ON2QrdwW67+jDK0dj8ZUjpmK2qu4
1+U4CI8Od56wqdj/VkBnb+Mow9HLopRpyjPPReU/fYHzN0CiRaFdOatCwu/FLxgG1HQ1XsB6eVuc
kULSOCkFViCBmVl62s7KoUC+K5kYJcwOKPG2HzLKroRHiBu3cTPQ2/ZW9IFBquRHt/UFwAf8Ihgu
TIVxgSrI9vaF1tsTTm+urDdsI1g3VGlsDvICFYVmORaDAFBLWZbQIuiGso+q66SK5jFB3fMJqvLd
z87nMkNO6cqQ14TIbLThv3oyc/9xd5trq1EsDbD9YDS6l8LL7esRD6aXW8Iu0yEZMV/npK6iI4QC
6v1OUSI21v7z7mIlB57WDamk0LmbEhFLeSDCgusc/W8K6fZWfi4CGOnLnRyh6kn9AZHUm7KTFajB
KUbrdsV7J4z//yNL06yIbiBXfnbPRo8OBdiwmLq0YUfU9nJGMufGeOp8d2faXHTf5AEchWhylHCr
b2up9T/hmbRBL2+E6EUIu+5gYouy2eU+Zy0QrpX1or2tkMC9oNG/90rkIdgzI0TeF10aFQbYDN25
FJl63bVJkPsi8EdoACl4N1D+nCVKK3JIp2eTpdpMkaIE2+Tvje3DsYjiSDi8OrYXQnegPXVvvS8V
6a37kpMIkvFVfpYSjveNMRA2VD8AYjyOQzWQTRAwDPIDZz9pH9MDb8YuxS6T5z0+nLKp6DMeLYAJ
Iew6LwauIXTR6oidXDOVO0dMvjwTeIbQqOsdgf1eK4R69AmD54mFxwfTc3pCPBMja/bOmqC+og2l
s1o4Lgcewz7a+X+0VOA3kiiBK8yzUYFmpY7mMpAsrbla2N3kKqb504pd1kMks5nVODfwUvQ7MQm8
IRJJU932rmQoPzr1Py7OvNK++6UCGgtKajN4Mk4f1BlX267qTzp8VGqy9WcpP70GJm9hMKEw7eBH
F1+8A0Cm9bpEc4NreWHhiEv/Kcuq1MPtSygtKjtmkeYae+IO5MqBLodB228+trdN3b5aBb/lRreF
ALqM0xeiyWeprTFvfbCcfvtQ+N4GMvoD6HdrEt2+sCg2uFEsXpP0o8ENrzde25GRQvwGH8I3U9rS
xbU+KW+xtOFTQqhBQrY0KDd2vA45xPKo38Tt7GOQcpM5ih41ccy4EbWt0wmA0/uStW+JSTTyqU4U
P8xyjRo6DP6TbtfS+id2WKYs/WvKfY602DJBj+dtrHwAgPXBdWSoHAAjVgbEMlLKlzmfOTrW4QjS
9Rke3p3rF4TDhsLB+nJtHwLmVw/gG9GbZDP0KtI8ijP7ACoNWp1gyg8c8pa6td5I/YyH5fSNqYDw
FaFN53Zy6vjeGsHkFU6/TbSA04yf+U7l871C9JFCyITn8y9xiRxtQZwwVc/+NHIAotAQ57WjXF6l
OweFekq+wyAXoRgOvbBFjtmoHA/OY8j956RjgbNJArx7hSS8uF3t1xIyQXHHqfL2oq8FArMwcy0S
DZteX0H5V24OTonKVUQv+xiMBHmWr4ce0wcjQEFuRLN6FsCWDaYv2FHSIKedRQPFXMZMbZ3CfBOr
dgw9rEy+bw16ZgPuAJ5HYnXOledLzIOPwSofgNS54sDI4bH0ohgYn0oPSpXXLnkLyJj8Q7VpYIxD
MexWtYfo73VKcnEIgHFA2AIQtwUqFkrz4kJS3ecjSt+VvedwgAFmxDfbGlQ4bqTm5ZONdbpfq+XI
hGW91h900Dh8cKgFNmFVEXi6nSAy7IYcim4SKNTLGpRHkoxOqjsA4SV/zh8r+/yp1So89TG64yyG
5CdCuiNhFZIy5QLKzuly3bXsXps3pfB126U3nDzYwYmt7UkC7m4LmG/KB2H/b1vkDBwDzD8Nz4/h
9IHMbYuVOCQFRc0k8mQALcYjeN/7+m2ne6XQBqw3YHiPHeWl03wtNASqtMcId7dPiqQb7OdlDVCh
mCxdkNCDWGDrv+slwsq2ERK+eSvczEpOXzkny5k1L+SJv/1c5xAzg2h4PGvhDF0Ft5E1wUYQ/U6+
MbHaDSdXJFCkiSGVmTYW+yKqXWkJ9heRm8m3/4XF550VxhqiWwtcGimGbph2cWJit0iPAYHzFBrk
TAN2UPN0uB6o73C/Lv1qTE/LBf3hRPhfm9y8rPORJJem3XqdxRlrNPs8dNxq+/Sadtxh603W24Ff
GsAkz717Z1CXGDU8Rk+wGXy79+0WqBa6CxU+lcd4HpURwmDAgB/2SfGbqin4d8VRAwXcbIssFP8a
zcSua6xLfw48DAVaQbkTZn057+kmkzOAI97KXkrDyQPqkheOwtHKkTUw/rczAcTz7ZuiTrM1eZSL
TCKWPmBcpKZPBYZDyPuKzGEbu4Fh4+ShR5ZwqWW8GXqzShsm/UqTpVMx3hEEh7Ou2TIJYx3TmJmg
9IMsMirP+LW12GoraGo8wmGdYq9NeeztjsoHMqMT7ayEc/1MI/ahTeeY+Xt5SZ0yAxc942KpgbSM
sLSBKsisZgDqHXgc51mBQoYQuWEpgqmzq6KNgcoZJ7uQhQSn2aKlnz2xQT8k0tSl4UsG6ENzUcDC
V1POy/2K2KVyFfOBKDoMuIhAIaGFup/BHfslO6KvQJQBGbWTFGVA+F+KBsL5BnKZ3KQfMpG+a3sJ
hcZF0BHuwVirpYqnS519sQQbtLBLoMdD4ETaxnkfmUc8QN86UlvyjDMxJjgIAlCWE8wbjcnb7QPw
5glcRunElUdebbyoeXWKc6lPu2+jvSCAufH5tbU1FajsGw22Pb3jKbFKakg9G4J6YrZ1mynhu0Nw
R12667BwaMoLCiiCv3m4+mO9YYMZlW1M4UOoExydhockSXFdrsWF931IOx7wxkJUdAIpsOwoQow4
F1ShNPOgYpVzmSML2w/67yOhRjb6+lUm2iJRnYsS2DXkBJwiNgVg6ctpukK8ObvG9i9k0xS4Txlb
pGCeFtsOuoweOvGF73pZOHq35VIObLD/SisM7gRuwvp5uLLw9nlPjw37fcSeMb52J4qHzo8GpvNH
zuNrkHPdwD+Uvaq3LaH9dR6aRE2KgeGCQr/BIbXBFfC0oN00zI5WTSRdu2QNP80wnDQhg950ogd5
K7v4eHPg9qPsSddHerKQFbR0kuo0zCBr+grodUbiW485Bl3nDIIkBqeDvJq5/LP36g7sCp4WbyGe
t5o+Hgwyyphz5Xw/t0U6WQ8iivO2a4Saqu19ApR3K6zZqHjf+nuspNwmg8nmlmdGzag5RbNWICRI
FB581uihUEEqAgzvktaORkhGSMtRsb69OHYwhDT62xDDs5RGVqT3FclJumJmBnxwmXujRNGD3Gux
4IKwfOEGXgbrJg6Tg4nHl1uxA+cGrk6yroVDH0BeI6TLhoNK3aqEiqdwgk/78EuQJ5Nw6LtCWQbj
nHberYQumKhN54G7LdBIqv0CuXcJmvh9memfw0rIT3ijXYncmgupKBYByFIw8a2FUli7s8tt/nc1
hLIBG+p/Mc/Rd17iM25jRk7v9PdsB3SK8MeVQORazQTfC/AWgVLSWaDerrBWT4X/+8F3E2HSbwi2
R1qu9XmlBg+OABX2lEuIw7MHuFQdj01iLtZiNUIkD8bj4HTNtAsIZDYu/1q3plIrDB1iOfWFVXGv
WpgsxlxEhx5IOB6RQS1N3bJdoDr9prkaHWh+RylRYLMaXv3YVz8392lEGHrHR9amvGPfq8h+JuSZ
2k2RJSQ5CMi+DZkxeOiOLfr5wMql5kqltqusYRTeS8U4WiT7RmZv62AwfxV5BQQbyFObwYIVvaUI
d0tw++mKBFMTgjeO49arhA7TmcoS+ndQo0lHyS9a0bfvyOMnaEy8BrQa7edSiK+7cKfLact1RpMe
IO3De6pyee5gzFeNRvFjo6L+pwjiz/Qz+aT9yx8I6NkJsqmwp7nb6cOpkM/JGQB6ionnPJHgoco1
PxX0pcJFWPrHT5oxz0xT+JZR50J1/Mv8cbeTaMDNusatYIA6dJIzAK1M3V+X0hXWWti9WBvrEJ+q
EoXvX1lW6wgRzI+Pmy4gV1NTvai98vCZ4zzuPJWsSCLyh7D9CLHV6VJ/rxIISEj68GJqTINFqSf0
aAV473RcDvUp8lLkm2x6tz/82TyhjMlRNRyGgc+8gmmJpYeHUuV5CcWErQEdzpy89eCWU4JPQTT7
X5lTgPUDvyrDcQsQA7PF90SDyLxuIP/3H/OD3uF0hHHE8+S2WKLIWWoy5qB5GDuR/VfEohP/Vozx
T7209uoxfScCNCrk0o7O18TpRKviMqT3LTUNfhZUVHIcVqXAsxphrHcQ+2ZPcnE6g/lerKGCu5Tj
s6e1fo4+kc4tcTVVzCTGy05ETl7V6hURL1z6zYUsiEWITTW4wjpFPqlZhBj3bPqO6tSUDWxyNtUz
KoqA15u1CRgweSwh4n20k7UlH6OzowctTNVqH26z3VRyI8DWupu6ExXYh1j5lQ9pFn/WLfF6BDIE
spCDhuBd8Uy36ZXlQ1B+fP1JDscQLBUsk1Hp7kI644PyUpvJmOCuu/2k2T1IDnLBuU2dHHu0MJqG
n05H1BH4fxwSgr1Ci77iXg4lpUo/uCmiAl7VtQpPpCYrHQIrlNVbfOLZ5xdwA9CtJ4uIunY+RhiK
n8qAL5iHrElUb+EWEXC4GZ0CLcT9MLkyEJKZXL9tXXK3oXmjiuY51e+G+VZfXBOzwN/cQ9dRwx3b
Zm5JHajXOmeENp+LU/fQZ/BN2VYRMtx1qmr4ayeYU9nuaQqs9KpYAO0v7UFAl6MQhkq+w+oou7OY
x5y2ZCWHZq692K1HqJt8zw3MgcETSWHkHhjgBER3cRM4Qw0NaQs+6dG27cIdL3jAc3+HByZudkPe
oeiddFYQoDuEtBvSKjpXKJsFOMSTuw5zFyZN1CBiSyuaT55jWPGY1DcG5mpdBHxjTlrJ93LiY/I3
NWoToAO1D5ALLTJ7JIJHUbSWCGg8elpWYWU+HFM+SodoMJm+ddZ9B9k/XEwJZqRLQdgCd03wWKS8
EJzacLukrJmT/9vSn5Yc9HCWuOdRDPIZcM6AeWPkBZ12PPxWlj6kHBdZXRaKNrDOlqGEZX6jNubO
A23I1zv69DH62KeEStctC5sMn4c+d48wS4c2R877JaLwE5Pb3KUhWdE0L2W/GPR8z2fZ8oOXzF33
VCD+k48UEQ8nZlMWABQPFMVNGcuqvX82wn05pqDbqhhbaPOi1tVLm/r3+Ifx7AXUbdDocA7XWpDb
2F3I6nxvEGP0TFWsgf+rg93yNuxasreFD5E4hXhvLtlr8FEYswMEYLBSiCwmLFhCb3vByVR59jF4
v44R3B/ZJ/5a4GduwrLO+4qGMV6QpSXux/0Ad+5Aop865lK/acyhuAiTXXwKO/QmS+uXI/ErdM2M
UjITvlZvbMkGOoLSTKaj5iWE5eDmaWW5zPMP/iCFKE7GDSsG6MdvGp+6IQU/3XKdQb/16/5buLlO
a/ccRvq4jLRHt8QUnkLr4jSt2GXulPV53XMzEOfZWRJnUboUAUnj8eDu1uV5rPd+vqZiIzrmwooZ
kWTF2gEcpPmJsLTmNTkPZKWMfqUn1GFXHwslYcYc4SR9/GPkPAEKJbNjD1lmdCJzJ12GZDd3qgEC
5HBu78cWJscOjVLmTQTwAWscKP5qHomKKaGXuOv6aZ794Zq++7Vu4SlFsI2Pi3bb+WnKf4EgG6uZ
CwaU7QUt46WdlgnaqLI5yzfBf2CJEaCtmFbFbA2fwELZgCN6M0EriOeEqKMgmiHIfpfa1h78m9K/
rtmm72aFBmrY0WkSDAsHE65HLKEMgoEvA9pSgisVr3NM3lBlDV+png9G1fSBNb64kzp7uyCwD+ia
bLL41DKP8DMZmjhRNMcbqikQOfytHr+265pI+I5iGZAmVfnxyOOtY/2FNxqFLlRwswg2sjgHbEYk
QasLaL4keX8kKsTtco87Dep+R7QsYROqVLjAFJJ7r3dRcEhIcdg1hxEZsTbfdofRfK18knjdjiOT
l6s0ccrzRUpGHPlxjbe1Mc5oaPy7gcEsa1k2yNfWGsGSzh4QUEQxUDNmU79tVaSgZE2S7KLLOKi7
mReB3UIZNEH+w0w/GMLgV3aMIVkQ3vJxIyvmXPXs6IvQ+tLNz1aIAUw5LrSgK6h8WdAXjKdAbqHa
rE6HPjvkRCqowfwE4kYFnNt4Yc6qn1ZYGXLye93FlUxKPATUWSEMBdmxOIrYWTfjV8aUkad9WwRw
cMsq/GhluC/6ytDkRog3p45HZ4F+dbhQAUMZdWkRiGTusp7ggK7LA9c6lP4fgbv8ZjO5Dmd5W78z
VFpOibFOI/6x4AK+vh6nFZzYG9LcZwNgO6jtmX7/n32xTfhydrNkaVPggloP948W4zIFBDTyQ+ma
t/N4AfB8uuyaQgUST2QSV2P/Jy7ps6i2wqsAzWANCE/uQfOP+xXRRRqlVSO/8dDNj6sLugbenkxu
b7CrtmTaTa2LYYpO4nQf5qIBd4y+gPkZxcY2T+ycNA3gQWI8pAaHmFzMWc8dnUSi5jel2AUM4jyt
3yCpwBy72j92QMYJK/WciFLnkvt5/Epy1ONIY0fypL0tiWwbRWbY3ehVPH7RYzMmUcBNcC6m2i3M
sViZcdvk5pt6hqu7n4xN9u7IphClGq0JxAkdpsanFZ5eEsUv6jC8/SeIJlMsSpd9NJg0S0eIosaJ
XPsqsUpmgDhP1DF0snMtOH2GLwWSGXxd7esMiHLgzz1BPQC6DBLGjsurHpFaq/XTLvq8J2+yszN8
c2nPUt09oqxtUiDe69SJmuQUsWJefMRA4Bsf5xzmvXN/ChwBQzZmam6cXQ2kGS56acoR0eV5kqWi
4lRd1eCVnHFHYOIJ/xe+QZHauD0/gvd+WO5l/fRV2OpBWpkmWAyzPGgNE3hu2DESzoMf6vFWcwve
5JJKfYMCw6unf2w44wl9pwyKdrWKyGZRlrKigmWf1qUVnVszk8ApTkh7chZURLqizKRdW5z2NKKx
QSXu7PO3ySBkW6c3Fnuc7E7WESl2pT1nFb1DjOm+qm1upnnsZgtHPGw1BRV456lCLNLuH4KBYxXh
vw9yrR32GnoGuH1OSCr+zYvwZXH4UdsPzU0DbJDQifULyqEm+7QVQvxAPOXky9fcP5Tm0fmjgBnX
c/s61qbJcjdhv4sRitfyKVGzgqS0i1NrgY61y8lgh2m5KuIiryq8TJHGb3Hbii9Aqx8XXJBO182/
ZwyE4s3XVwGnKyseBLIK7pgesLRlXbHCShVLxtDmSnwdmG8h5POAiMv/HRkfhId/jBPJbL5Ix18i
lOtXF8oiiGrTHWzM+A2lhOWtwNRwJYr+p1OSz8N2cknUTqz7w0vRRSATgy5L6DJUmGD5/kLNpdEF
speC1rF8UrZeklI+WDZUMbSXyt9IzNPA9w/L61wNchb1avTmvcTuB06qV/j0dWVyiPQ+AOgOoy53
OtUjkOoCK10vgpT/tUXBc43dALaKV1yrgfzj39VXQLkrlnx8QsxL6RZc01a36paDGsuZzDFRB2zS
P4YMuECp6c5xX1ML/VhzmYdr6lA1+f3dT9oKdlM6g7aRzTVZapK15k/RxWNHAyAu2G9YgB+xkPFo
tNk87VSD90bkTMsrX4o0bdzwl0wRefa2uVJh6sOQeJDLihhGYDSyiXbWYDcDgST4nzdCZPeuGw5y
5dZ8k2rIZqh1YIcrbEeq9jfEUevbXlzyQgVRHEhHS6NZwLODU/WL1mL3VjVvq7UjOIzUAf24xpNf
1w2NJ7vZ/nhTWMt8YkZ9qVAVS6kHRF2c4qldCWMQoJi/SnsQBrxN9aRMFIKtQOYU//Je804eRQDm
pN5aRu7Jj0DNIHTkBZ9VGNijWfUUevP2dR3HlPm/OoNf6hrqBiugEuvsVeUaLDhY3bn9nwyFRaBS
qR9HfAeVBgXWsEVqSOJY/wKB+OAtQVzX6VYMpVdjHd92VA16PfqR7usysCaMtXHoDuYP5dBKBlpx
BQjk//2BIPv+YAkKUoOhKzvUNwjnrs0NYG2Ye4lF+qR79Jk1HzVcEw5gWEb4MLUWvF41DwvvnMCh
6RKN6l2IqsE48kAIuQiELV+I8qiYQTlNdcszMZRBeuzGFEl0SxpnLibQMZfS5JnmAj3Ei3OH6XmY
x53g29JUGAExvZgMHYz7xtbSNQGxBgfmV1RsGXwAFcWRwybzX9vKYQLoFaQ735OVzywjUQZODzKu
cNZnvuQCDJ7KHltGsZN57f/ijD7ThKX9TmCDL9Kh815oXk2vhpBnZINeVia6dDRm+eXj5d9QWiNY
ysfyFjM8li61jW8ZWqF/Bj4U5RMRtYVsH8ux+XHm+wZpcR7RTk4RlMzgqr2t3svQ5GeTaGp7eRqu
Vh5Rel2QguKWSzYuUgN359wv/6ex6bwScT7FGF8wTE7/XxVlcXinstij3/oehJkgxvGq+iNMjSgW
9o8K6o5aiv9HR0bLmwSoIc+a44GePcm+fl97IOMcl/U+h7nw9SkUXUao2tMSq9s93nf3IqAU9eeo
dRGYAAJ0Z3cOCb/IR3962wSB3yLUFN0tlBXEqU7lnwn4WiOBm0Zu2djkDY0t/a+HcYRdsuoju0F/
HRIfdHjOLIMInCBaP4bC4N43cKHzpi2+TREC2NGpfHSopWPT+Yw+rdIJXv+qUSn2Lm6+zPWk4IzD
iOJ8FPYr+jAnHfTbRpmn1WQehJfAcK+iDo79eL1Ja1e3ZAZ/B6UkfQBHKssAyEokd9Od4TDp5efe
yMctaMRxhpeXF77eld4TB+tus8iWQ5lpacdnF4JxlvSZj3a/+eex8vv+q2CcIKY358f9Xm+tznX3
IjGBX7nqby0Jsfy33SMTUY6jO+/exw3BN8loZr2YwXJA+Kipymzicx7P63i4q3nMH7DghvhVTxqE
5lbEj5wuLCJ1MJ9iq4EBNIlQERCCwwUvmn9muE9aeHRZsQNcpyGR1nLREiNSzljGggIq9we3xuyK
XNb7FwXH2FSnSxltPn7OF7FVp9cSInw7Xq6bWCgDPy4NDWQ3BfqzINvSVgIq5I5RQPH0J4Bwn89x
qdejJZYb/twMwyyJovsCYXwBvzkf0BdDJsaR/qZk3H50fLWMYqtCpyvIuhAQDrRD/nif3/8xVJyS
xypj06UOc552W6PtL+aJe2nHw2tNrf6pQ0pULjKcxKk5px1LiGx7rmVPFcce5V/FE1nhD2wwvfQ/
pDLziFLsAJFn3OutcSiV1cElCMaQmrcDNHviqnFfS1q10SUsCDZFb0+xmiKsaLbOSSnD8VlTaB8s
2DVGQgyKE8hOHmISYA2HuWUYxfHd3uJPKPtLNs7dpSpH2HlvWTzNlp+QYfevweAzVh85V1R4yX5t
qBQ76hu5h9gr/SRuSOrhUf4U1QnKs9E6IUa35lGVS06TfizChHpBpr9fbRifFSAfw7YHqyO+mp6g
NcwRrAmkMuWwRXEkVqFxfp4ciMdffdBbbVfB620ndNU9mCNUJW3za33c5bDEb9qsdAdA5ZH75Jos
TZ4clp9oCZtzbXIK3Q+ISr4liXdpzk7lxqo93gX6KrvFr4hkiaJfeiNL69c1Vuc0Dro2GXfe0JPw
kgLMpd6ybftQA86Ln75o0DR7pUPGVtVTM4MpRKHIj2qfeyWB11A6ZOLp7/Uvs+kfqHExHPMM/duC
13u0WUv1wrtmfCXBXXwNsMUOlMELQKYz55NuYWTPjH6Ac3frf0xFdn/MHjhjoeScGFyyqQkFpAdx
f/qRGin+BzxYRKxGrsPWCPFWuo1ZdHBR4TCIumX5/I+48w+7doj4ygRgg/zlOwHoImHKHar22NpU
f/q95DbWkZk7a9L7ZM1EjsXh2tXafoDxW7RY2Bcn9mG9G02ibyfNH7XtnjYnnh61BVW00Io+liiq
Tc5i3Fn47rr8V43bc2SKs+5ULPGxG1LGiHbjwm3Oro30ibED3ltbqN4rbUrKSgMBOpLGiDoUk4OP
1ISMlVdSXyhOqy4JBg1kIF6mP7i7tj2idGYPw0HX+hy0As4FPrGXdPttKULKJ7M/CzP1CUljBD41
iJQeVUWQBYVoVL6E/AR13lH+gszAsTzXBxr2cgV9O+7i9XKiFlm4OPyZaIco50xmGOaatw+RH4H0
s0wvjlVav3aKuPJjrutSkaLOJzgulubdCTW0aCBuyo/llYRNTNz1HbwXQbhGhi1+/jl7wSrK+uNl
+6WF01WeZg0MXjUePYDAuLWISbR7CqPtOHQRMkJ5I3HugM9sk4Zx49gv3R2exRexWKmeI9HQoWPf
cfXiDMn8W4E6i5c6XmYnH18SeKRg846iVMAyotyLzNV1y2j90R7IsFmF25dhsJGkDbqardZUWhMQ
0y9uNeeUFdw/B74ZZzdmY0MQQ5FqH2xeGrIBzyySCV8+/N3C/vobe+r5TN8gyKl66fnmSaQivFIH
5KzdZjJeXIfGMR1krpo1ieqaeHU8Kwv+5g8quqpdnIAUS6ILF/p0ovgP7B/ebS25SCZ0HGmF308P
kOvdDS2jGJRW8C7/hlk7qYUUNk65EtpHSPuts1Qba/veeNcSyifRqZc+AZiadf6XzkG8q5Zca2W/
YOozZZoBq31ka4KcvcmAwlL14pePezBElsabfiyRvvbyn3CaPbwE6L9yx0rGpBvOcJfzg4vl89BU
SwW/rXiW3ZEcIFIc4ufm6r/b6JqejrJGYEDST8oh3bkLXcPeUifY86Ai7rNmyIPnyLRZrvmsVwiu
plo02eUZzKN2e774aY9R5d+VffUNnHEWUk2gbh/Q7tbA7rZHFRuzvfU1dCwgHKgYn1XdTP8KWBwl
A8q4IQ/rwRkOVXvA2cdWjkpqJw+JkBSCR4S//TvQ7H9sQ4sI3kKXQkIdtf5sZ1qODCqLSuPSVVj7
JSxwwLKaUycTNtUdlhHCEYnKs3Fc46G9pgU1Y9e3rFLCX2Mq1Twygfeb/puF9tdtb4oZluxTokIe
bRvEQcavf2bfKm7Xmp1obNZybDR+SNtBE5iZB0nGRUcVyUSP3xafIo2ZQ5sxNdUP8vUDPxl6tyiB
t2F5Y+NDSJr4PzZO79uyTY18W7DWVudDZ9d0FVzjz1/mgFL4NzxvKVvU0kSbo4FYFkkf7l6a9RXv
eRLNoUXctenzx+jXF3sjKYEhgHSRHVT2sBNgzHm9Fiyl/VPo9zaqMtnMx9nDFmIcRpIXzr+RXeOw
vqGaGFqvzUr4dy5FtCEZV7hhxqHRQ0co1AkK75G7Cpdqallb7TgObSAi96srLI5pmNBdlzyCwUf7
Y1p3XYfwIY81jxzKZhTAn4+wtyobqUmKzkOoKdOXti3lc6jG0SbRXvpNZTAoQYGIsbqU1janyZ/H
/Fz61EyHYJJbQ2RUxGyHEB/2WaFel5H0G3txU+WOsxNubjEGUcS3Pj/veYUXlpH+3D0ksJzqVUlm
i1YDCaEq50pAm+K1KRSfHGbk/gu7OVOwbsGTKsrsvs8LQbYUDOqE0NShfqYxyl3JfpNZBZAM11zC
07dmDwlCcXUNbi613wMjCBQjY0MKs/IS3yjLcKcTiGgjuG86G0qw0bd75wvldXw185AgGBqzNI+p
UkAE4sdlY5YCG9XYJZ7k+PAc+z4WSo4U7bVXp5HR8dyhTQzoIagnjyPERTpyfsOPysYEXAlikfys
FRSqUFtqtHSXbJINIHerPy2cxAB4C/7lsnx/7DF/Ljao07KOPw08fIx+LV+D8Evv+KYGx62PfIB2
4KUczorp/r05bwzusLMFvFXXN0u/fSu4HoegSuTIUX4GX2HSzOZyeNZjOL+yfhEOEoMSvoxftwbW
AEHVhypKjv1PYzmWRsDTdCfLrOIqOvgY0DsYVlr+7qIt5PEbPgwV/3njeM000B8PvuuIGpCk8qKn
7ThHgAfmvqfPUO8wYMAW2nNtykYsCLKhe1fIwB56y1D/FGaRZUZ13jIvcnH6FyRY5KpDqhVnLyNp
uq4gaxLehh6FyQ4uf8j2RxWzPszyp+t19/OIFyFKf8+Pnu+gffu3aK6+j8j0QNS7b+zgxrSKigC2
wPSndrqnoncAO0/uidEAbzuvxwpCE07ImwlVzrRt7xUMOrOlOBMfjVPerdmB65A5ymsmVZbxb/iC
V/nc0xFODgoNO0ryl6YObzsx78/TmSW/Tonptz3j19Vib5gw/qP3djaceO8gjRS2BMLbEDOMFMwy
gCxPr+bisMCZlaizXVLFLDjhe54Fy29TKk2jVtWI+AuWEJ9htLkWrCOV4xUL7o/qA2K7OMvgUcJ8
LA3qRBg3H5xXER0VuWnG3w5n4+vEE3z8Q7nfHmTIaTZT3gd+z/lfdwUOzTMiRM1srWcu4Msg82SM
mnwmG8z9Q6RlZbfVWzx74E+m949goGG7nfDDvUeD2RwJCcD4PNLEQrmItej2nwBIitKh2zj6r79N
cwMw+yqcKt5MLt3jKD8AXueFVSh8aSeyje953Hpsjph5Fth8kuG0xjTomzE1jpUG+wVpZZmTfoQD
cnx6YqPR07vsEWIT1s9dGDHZVvZtMPjhDIMgJv20lPLXV3OMnKajClNLv2nZB+KIzfkVi6UYkCOa
tJxsnDWCfOtHTjXcwS70KhcVXYgksT0VPTTN6JTECKxFIr8OWLScFxJauhcv1Z31G8bH4ExQq2sL
ZXyTXUdq24ukwYRTyCvutExwOG33mem9vWi7NfMcH54JkZAmdmi0T49Fz2kniknOiKhQbX8wiZ8A
a7Y5BbC6e3Mnsd5tctkcYP5GEaKzZQgTArOOvww5sgcgUWnRH6fhwYRnvALytrlEEDtHNzbmO0Yq
V/3qZVI1/0MEgepfukccyUjqYfbQKizi8sA4SvOhuY9WR3TFmY4a3cuGz9pk+7xH3BAd/HXpEPdV
lNeGtR/ocRyJ2Z1CeAVSUZTao4wpR94t41YUAaGGUSErFAduqPaIKzfmAoXYyZrldDVbW+KqiLZI
Wt53dMUywp2fJpT7qhsv+0npEwqV5ExMXLuyRdWN/usU9AFBlqn3s18OXxJsOmRz5ofWuQhH0Way
IWPDm2wWWaRPoHZ8hrVRIiIUxd/n7fsvmHd2BEARdlOOOL4f0qf+Oc0iX1MUjwZdq/xnlHtIsxn4
izqoX4s5DDERb0O66MWbRcYrjPuD1q1Y1lxCvyHtADxfp3OpX0YdOok1YPKFm2CcyeUPQlaDbrQR
JO5wYPm/mEA9N1t4RKprjl5OvNI0JMBzjy3Q3b8ByDU4hiPasuNBRPBhptjxVEEa4uYPIWynvh7b
FfimDBbUst8craBDkW/ziYwR6Zp0lcs4/ntWVHPvST4nbynPa1SYsymIHY4ovOUc/GphV8v7lluB
NhazlN/Gi80BpcAfSee61aLPQ03rQhygdS3XJVBD8mXm9hK7Cz2EEBVxZxaO8yN5NBfIQaNolNuJ
v+A/wNyWfZoJ3tNGjx23BsPW7Bjg1VBbwCCRqYAg1iwv/grTClFRs34ugVIlvuLvPEeGrTWPrijz
zor8IHu5/94Arj65/etzNoumUulslK387z277guufZG2Kg1adQ1eBvp3N7WR4Mg3KnFtwoeEBq1q
ALEe1p7A88AEEAwQJTPkpKTP3tHjN0LW4fwQY2vOAEBnsm12mTaJv0FjaYoLPo+WEvgs1y0xr/+d
OGdCrJO09EnPeXB1pCRhnh6X03RGzTDlpNXzOEf+sibjt/HzIwXx9JG9BUQClv3CVyCIxuP0lHjM
2xflyrqs8Y+yTiBsYSc0lGoiNKa095kzGDgwgF7pZVRh5vjJvEVzbz7qyFyjmyVn/rY9Zey21hwU
iHwDuW2ajYuUBu+oCiSa3mH58JLze0GFdWHWJJO/toM7GZasZ8XPIHE1jCvxkQKtllVHEP+zlblE
fdgaxc1SlR232WmDkOYaM+bugjnAM65T7walCioRud6CroFrE/1LF8vnCyv0ccWtZsRxq1W8R14f
lqbzTjLscGjwzV84uGbXXujVvVidUCc4H/NbqGtFLZyawUfDcIdOGof4pWl6HwLoCCdxFC/o2XBB
4gZuXvoJDPW/hidMxTwI/i9NedLda41wzO9klX6AWNdHUil/9mhgR4S5SCS2ivsOyvRQr8s8J8av
gXmXXnu2xjnlrAB0bZxy5hdlNs3dFLB57t5fgGBan+mzzbqYQj74SgZxTlk7XD/bwWChGRaef3YE
r8AHrHuI2XHk1eMzRaLqwpW9GjE7D86wxwHX2GztPRC7SQ71oOgiSml7HutOPjZhCXOtE6xkApEC
6Tl5TR6QaOBAjbjH//kyT/ChPqte1WEwgbxTMu03lWib+rcBDBWHfh0lNOPqD6EoyB+uNNCRuNKc
VxjnG2M4ZCk7WF41Ro+2jEGwDYOCOXcWACptHDnirT2pv2IpigoFSakaZsG4DWDsdkFOfZQSpJhQ
Gwbw2RgeoqSj5w2Y8AtLQhwPMdcT1TdEbMtE+d1J7kgY2jQNHz+r+RCE/hgLEV+Mv+MsEyOeMu+o
Dapa+WujwThYvQ1nqq366i49pMV+4i7fZJeT06cGEAiY7rgjG9RvX3vc76TF9TpDxfE8u/0fnM/R
jd0wXgj6h5L3Dg8j2gzSdJ7fST0uLn7AZs763HbpM8yIUTHRhcRQBhiGU5u7EEv0N5zuiWLdO/5e
bLiT6p0PVAOA3gmMz+HwOpJyziw0qg69Pxn/xoEJsjUM/dZP8xy4BWN3BXZDJ88IX++Z5UWfDFRF
muYCwLLIv1WnlCNMYxQRZiraLCOzqmdMrzPfyZjTbliQ1w2xRmkkvzHL3ru//bd76RxqRB1YZHVk
wFxC6846COEtVKdgIE7KeYJHR2BVAm/UnnLkwBeXh1NpPYomwAe/UOJX8ptdf5SGmtWVJ1TGKZav
gpmNpcMX++TuXv/IUV4kaV5v9n3o5Pnlh8miPU5oKih7XryPGSdAx8wTuDca8yzPGIeDDfNhlccf
j7iXbSv6fcW5uNO44bpONHGezwk1STkYQ7kuHHx421dxjCDnuGbBfpxvMjaMFUJE0JWUclDGu/pF
C3yz0h1AfDL1Nhd14XT/JBwWk0ykhIYvb/DlAJ6TB08l2uh37O59nOs4G8EuhKnMfNXi8HIjBOKy
Db6linFpH23hMy97asQEj+/OzMz4S67+sMqg7HGxe96G1MvKXtsvBUvKr7Lk3jXqN+MFQJsaHayi
g2Uhx7wJfMoT/CXxMX9Tkjvt+NPSvJ8YF29KoFmbjTohfNvxKV4WAqEWLutHkX0Eq94jgO3zGMqP
yY0+R5klKnBWaAYREWVlf/yet4BCW0IpJJzaDLk4O6oSH9ulPdjaOybVy/yml8DpWFLX55kE2B2k
uN64D9bGN0tF6reBfYxNiynyk2nwjcpcuNMJOdwXdhAzTmGZaRNI+YXSf8H6bACHbKgBZC1InAor
WlSTZGBEYivH2diKKCRrzor/6xV8cho/PBbU+dHTZkcUlMUlkJDSQuCXACyE+FlM32Yn/HBClUHu
PqO2gJIjVTy1dMYDuhDUOBBYqVi8+QYsug6plMUuPDbN6dm9HwSYZ3OI1O3fZczzN4BloR0NadM8
I2doifQRMldNgw6qUmt4rNzqrQX/dVNYcLRIVwgjY+twa28MoQB/+6wjVFgERdAvNxrC+C7fj0as
h7v0nJU7FGTSBhIImyiwCXxMDkou22iecc6/nQgBkaH/Zng1kyNXkCe0QCOmksfVHp3agsuL2z9J
MQ8eeZzIooFCOiTwpfoiIPnHqlD+sdhgSwoKVp4urhXGHgya9eMrOnwKxDVlDoanVowpvKNGoAHr
p5qBWJGhg+PIrM8x4NVSsGd8UyerMIEAMb+iRCKFre+7+2trCQiw0RmdjixK/xX5+4iVpk2qddvM
qIzBEzLo2PUDnPDo84bR8pH16T7crSZjdZz22dRgN0WHX6Uw4/5thpjax8wrp8zhjV3cE91sO+Pb
flbGubXwBU+DA+7/6WBVc+nnjbPa29XiEXf0jsIbQTnwWs9OUf9ohfGdfQ6GBCPIxgUKYTD/QPIk
1bVxwBedMwTKC2iX33SWlttT40O3WqltnLf/FCTQ45WafL5FWr98Z1mQYmUGz8nO0Gl8afzEmDO9
zkrwWVm4TGtQtX3ySFhedaScr7Xio/lxgLM66q0Hd/AekVeH0YzrcK/88kRTDHVOf8a+ulZ/Bhq2
rKPtQ02SCyRahLW7/T8Ppu39uOz0dHEED3lKmncci9704S9P7DjeN1qDRkkcorcGaJqFyamGzd42
BA6awNdy+5NFYXEJKDyVBbDCs9piPZZRDAd7Ea5OqdwFLUzsRmBBKQxvpJqEyf5yONdfsouGbNgV
efuEI0gniFz4cCgRqufVE204k8iT1vi6UJO3mrNJCWWXNhww2NyYdEe9OoYBp1V3SyTFacJHwovO
dPip9hbZssiUhu8ewZ8l7ies4IlgZbmkT2JrpS+5MRWqSSpwCAo3u4Ny2Ayad6AA6ml8gRs2Xy4X
bU5ni5aHSP6xpR2UV3z/dP5FBmiDKgDtr9SZ2LINqzEwlFBdPll7CHri+j9bncphNrRMeayq2v48
3P4djJ/9C70AVVkGZyK69hUPlBjjBfgD7RKHnmMnfy2GIY7nmLkSk0AM/e/c0WFK/bODI0bRs5lR
8ZhHnfCDrTbiGlS5suN2G96fth44DZBV0GBF4UVEZ4095u4qaemvOjFdR3A6XPiGb2gRM+Tj2Su7
vG0aQ6YTU6Lwd2IFswx3wwGeOQZpH6hJLZO0e/e4h3UFd1pfou7IIN7y02b4ewgqMA33nFL8Hd5A
8mvocKLNcnHWJSHsc3lRaVFpclJBc8fKqw5lbksYoaE6ZkB4cOd0oI/SK9B7gya1azNGGdagGMZt
o3b3bZOaXbALRtCmFotc71QAtCAFqxxCI+dPC+reWirx9pA47bIL6ju2RUqF6bykMAdANalpnSl+
iCHWnT9e9B+5lTxLuT+SueXc/3A5pyH6EJyGIcar8oXGqmgRJyJrGb78t64MPjomu1cmKdtaAw8l
qvF7Vf6bGp3DWaPtorjIbbz3uXafyG/KcfVk76WJfidOYsXLysA+roNwmc3RImyr2W/OwWs9mdTP
s+rkjMvuTBck6BPGmMcrXo5QOos/BZkuLeQUUqzyrIEzxFtz1pJr5vcTdR7kpI3zJ6dX6aF5K/MN
K/rfqc3S79Yc88FhPRB8dUEqyhhdlndm2dWShe3hC2cJCwhitwcjqsW7U5TlMyQ3G8Po4PMiR41B
o4KKpG/dePhiDR1canqmi9aOV7GmhhCibwEFPUBjXmk9R5oks9OCDSf/zjBp1tUYUUgZTM+13y0J
d7vP1JGOgwKegyzYrv56QjVfK0Pnec92ogaJQ7Wme0Nc3JKqZcukmbVDYsk8Is+OT3211r7Kcw4I
iT1F4gGeAIg59EPs1UQXMZHd1vQTa9q3QG2CrT9oNsLw8Q/+YHQB1qNInTXhxDlXeJ6p4B/rJdMc
bhsuNOJ7Y5VLj5Ao0s8GETph8m/vqC+jkcpYqgUmQcEr/B20l0jCLtI1jBWoRHq3B1KGH7UGllgW
eBZb4CKl16S+6MrrD4t7o2038oRUF0BztJUgtk/aKC864p1sB9ylYi9cKgRWgBMOukYVdiYLzhrx
xLlYe9vj/dcnLVQslRTCM1sDvt313iNhUZWsOqX3Hxryu0x/3iSPBjBxiDQzCuk8X+zpu/bo3WaD
eC1yN8kIanJNK1UbQMG05jbx2yE/UGwxcKOlnudBA//Ii36P18CIgbwVwVHzdHw5d7UpM3P2w8WE
GXEfpLW0kBauqQSXgnFPBPPl5hNVNjt0OGkss80B2t0NMWD8P6Wt+FkF10Vz9I42k5KIgzJ816XE
sPeTJddnBZFWAuTsgul67krQKGKu/cgFYnesxPHzz8zliQhbyWcWglaE5cENBGaMqJxv74Cwkm2w
EZK+usyEuCWm6A0hHNvZcwxyFxg+Nhb8ay9OTOOLqi2+yGnhJHhw28LT0XqR62sN1tWft3iepTyA
w7rt32li5vvtrYljRn616Dgop1A4RXGysIQoQN9LwyXZZqwx8UNoyZ5bR85B7GU/DkPYtNzbk2y/
fR1yASYf+7A+Or8C168jbPM6y/AEhbUHTLW7UO3+7IBiklRa6UhyKNRWP3VYmCiaK3S2UaiOmqvl
9/4dazZhYhBOqkhli16HD8FfqQ5Is8bb8OHeqoACLok0pQxNek60I/9w7iytzes5FPjL+2ipWIQk
y2oZSBm8CQjX9BSLn3GIOb2JE4LOB5Y8oP6Y7YcFxM5vY6Ck5FnwKHHyHFaRMA1IS6LqWnRqGD0f
rPfYUGPGOeh9wZ7oYlOQPsOav0PJ5uBOlp+km78PDMIkCk0N2K5xVZaXH9nodEsCZfEmGJye1GG+
Kt0dX1ZdrsXP9cbQHJM8uy29F6HHmvjbb9vGprwCKeL9Skj/AhPGzgVg8u2MRHk41k068AOXkvVV
CyHkDmRpaqcDqrkpx9FoViKA6UYudfoi/MHjNXfxoHsT7M+0uvWQKGFUIWuYxhOFFoDImxHEwrEs
tljiXsRGxP+npERCsnfTT9vfpQ9KifqFtsWxSYt/wogal4/lrHUbRrXtakDCqcEHZMmoKQpX43pF
UJ3HnnJoYG9fJdQOS9auTqNm9p73m2W5TjEK9+BpjDM2i1JNW2tmFJQs98dgNGXAtOSwJnNma3OK
ZKtMEZYZ+WKYohM3UfOMZ/oC2vvoc45ZdrMJnTgCW39uHQp06dzFHSK8X7hOft1EOMXQU2h00FSN
rbEC7Xh19xGi9hmSLpYZ0yaOzFyPc6+d6Hw8LUL92dmu8uEealcZsyUk2Hd3FSQW0zSQwqWKfD69
1U14wYdr4WNL74lTKGOCLABf7tAT+GUAITtJqeTgg2Oo5LZ5vjw7kcdgCUQQfIyoB2watolfgPuZ
iXvd9c7VSUauZMdfTIbXQvQpKeWtqgCFUFuMScdYDdwrrzWftF3ZJB1oLAUsco6uf5jNhmwJV1ev
f62Mf7wNQtJcRoA+kEzKf/AzZcZtABBaRKk6a3b71JxTfZuSkpZ3Qxn+pZsIEw+K1ZkIKPQWwFjn
et4TnGSYCC0Nz2NayTKUbXU5lWR9n82l0b609d+dRi4r6xj1OnVW7aVdulr++B8H6E5i271S7/P2
sJ9K+WL4xze1oLBEyBzWIOSIyCLsH7iwVhN6JeM+vzxbqtRVxquQgWJ7jdY1H0+UwOWJ3jvqSUGJ
MeWWXVV7MG+0uY4mgwclpxhLEbtaTWBNJhHPWzFOlfCTHctmskvSuxBhdO8nVmStdtqk6SUio5Ho
hzhJ5uuUloKzMTmI22DhKHP3aTsNHHt6pkOBMNFqDy3Jmc9OZpnjODliqEuDqKhwXAKtTZCBuR/Y
W7TuyN5tZfHEauHP62DFvfyjUfDqDyMl1G8nejkTHCtouCq6sqr65K9OTvziZGQAgWsVoJhGWbYz
t8s/KX5eb8u28efK4K1ASmQdGQvVD8xUH4/2EilLZ56Sa//aiFtuKVoJK0zePFkt/YP3V69jkKz+
l9xg8nuIM7r1QqlytmSqMT8LBHKJx3PXCEZJsKx1jOZgkbMTHrCgNhz1RNVEG4EOT+0XB5xtPDYY
28K9lZeXs8IOC50mhnARC/JLApfKIDhvh5nWP/bt9MmkhckzkWeIO7M3fyMNEfhd27C1ECTaklGC
xgMlNzU6IUfPc2AprLGBLBMqnHjqI3Rg1t19ufRDcURH8eXeu04OV/p/o5y5t122cskeXahhen4n
6C9Bga+ASOBpp3QdQpOkRDVIPpsPuFLWWixfejsAFhqLcULo9ZiMz/W7bGj5r7/M61IGwm2xWtlS
Tndk5mz3O5SCrvs6ftAtMM3V+qhhh7FmpdZ8Xg42okULa3Om2abG9udSrbnR6Peu7Quu0s7/nkzg
uclInPsNOtFu9wqF7FOAsuoozHB8HyEB7BFgzMlxT6DcN2iOLmXABFpLMSEG1QaxCx+57qmQoMu+
CCuB3itKPbWtD5Ayf/duhcyZSnlbFNqpoqgGQPQ6inwTpQAySANchPuz4qNRh5kqLsGSruHNmZ6l
XJoBvm4C0w8UVBLzSsgiY6a14p/uRuoR0RrUuyPQL+Z2MIR7fG5BujMyUBZBzPq/NhABFVyI9VU9
NBAZb3nEiDf6YNdfJ+eoT4aDfwcApeGh8NoSCJcnksfzoRM3Iqqenc7KjOCSriZGPAohUum2XgUu
j9D5YwgYmfWZ7udDN2weA7Z9wySibGI8qjfh5kqHT2NR1pLFKyLymf5VXskKRAaILuNG0tUCZVoR
vyPBLx5R5ZC69vwHDWIjBJaW3p1yeU7wz8jlTUOssvCZjZi1Fvhq1gaW3GGv9pQK0Jlgnx38XuWK
LGuLmTeCuY7jUiwQaDr/o05jiiBgnUgb4nudv+rOCnfW4UFVu0QhSZq/sUBA+3bDD1t6IXmybKyS
X6FL5oEHSXdZ3zEMAVJDxWYBUNqp0CV08xTYdqhfjIYgzMJSCTY72/4tUPJpuSURagoE8a+oERrB
r1j722ABWD96iYpBpLuCP68PYBd+4fqP1lh6Sefw/37vYYOoWr6Q0+t0maXm9MG/9YUtSyxeF/3z
H6RHvXsPJgElhug2B58rahUZ8O09ggU//DXaa8xZUWGJtb9gRtSNG3kWoj+ERyD0Diby8hmFaUJm
kmOxPNXVSy1OLL/OOkmfD8AgjHcbL3/5E2lPyl1US7QWuPIW+5Ed7YSFdg/mk21bL3LbhcEc0f1T
qZ/e4Oo6m/m3Knohz7LcIVOEPl7ieVgp1H9NJbP00VuNQoU12rypYF78YpD4jfGlh+HCpOFid+PM
VSulMb9JUOmEOrWYY1Y1PtYqN1eYOabpYD2BEDVLfcA0kG3tTPlFPwpLC6Yy/hILvLlMAXjrbwDb
waMrlSndwbekUckDEgImpUbzmWE2lsl0nQGZGQMkmUldrYFiO3hBXkEsSyeXe9k0P2y1gWTnKmx3
tadoJB6UnjzESbI4knkadTOglOCq3dgAoq9AFpHYRF4LI8Y2WmRobG4te3/AZm9fBFwGoPN6Dq48
56rMEMj4piEKPuAyCK1Nki+Gk1XJMs3G6m2HPnbjAiaxw5oiOQSk4fMa+LfTsj5GLtCwYQqtKCGe
y1tqnU+L1ZWdpvqs4JG28b3ntgMTdGTj2Mx+rKB+S0sO47HGRe9zHJb1Ge5nHyCbEEJbk3cpEuvR
A/aEEQPGxRGAN8CSzApu9jrUnwnlAgDOKVvPu+inGqPeq7C+xCWgbxyQh7poC9fgk8ZBDulqhZ2i
2/v8tW4X3dzUqI1ODQP/FB0x0qUqoGb5lhuhUN2sV0sP5XH0ZZzDd7vhdseJ+E9NHA0OIqzgS3qp
2ohIM8onRtks7tjFz5AK/N7EMKnVHSDspSl/7yL2KvDHBAakt5+ITo18opYSlETe2+DfqJensJgw
MKs+rANVopVt6oxExNIjjxeoziDZXvE+VbglztzGT17dPQW5slxAfVPbkHptRsITAvSdE8D8L/Jr
4a311nilAVtgiXwTtOyAO2xnbltijHAMMj2oWvAQf6HUql+VrCVNGKkCgbCggtzPS7bEbp8RGV+2
RvfIj0N771coTubg7i38n/zOAE0zPJZ83e9ZcV1wsc23gaGB07EJ3WKBKKxCcSyrubJK4sVRUQFQ
ResZiWg5WPaJi6IGYmgye2E7Fn/ezvNZ3RmqoZP/xwxS26iDLtCJxUIOuDVitufw20hC78D6iom6
YrvfaQPaq/VLUkyPzr0v0JEkzSabBFSROPvlHbzGxuAXXy0wi78rFMT5UVja+htFM0bN9Wex67xC
AGz0RkHiMVTdtxUjegZX4V9KB+9uScMzIGLy2NDzcb/caxPryNwJN62b0/2ByK128JzPXBa7jXx5
xqsj1z+OXrxu3zIt6uehAe2AgsezMKLg9MAggU2T2iJL1jSiDp2NhQ2DR6f+E0IQ0ZpAoP7sRWri
vKmOdv+bhHweMS3RiPdrUAPkNQYClQx1dm3WmDkh+WSdqLsok7q7w3b5FWBIsU/bxs8Qpj9AOD2E
1J4/QtFoxS0E6wzXG4fbz/hQ4SD3x3IHIuia6KmnWH67G8HkHroJo0bpR4HmSpU0zeVx09qxRJVr
tvMUU0DI+wLiebtIVdOSD9DuVKCrMgpNnirJ77Cd5/n1wth3Hptg4OWpKG6e1fg2AjnAVXHSpr/H
0gq0/6eVYext9HTsQotme/iPA0oXgRJfP1iJ8q1TCttTuSBYE/zMp/d2im1TzRUXHWcLO4sN/Dmo
qOBE1ENOiOTu4KL3WLHDvQjnuQm8I8uM2Uj0ZVvdlJaaPAu8Me6dn8uznpgHsl9ooclfhqQi3FzJ
uENkRPilocauI9iGcpAYaJA0UlCzdEc29yB1vW00WGwIs9JFpZO0zzjCxWZIRrvsyp2xXuIH3CWS
/frTBmr+NkygUQ0XAf1PY+01SjvFXVKqeJh6TsHdjtA2VOe07CzLo87LT8HL3TabrORaR901j/hH
SgWt/fKZwb7v46jsnwhEpQIyYKBmLO+ZPOfB3fhftJG1uOdspwsxCNAuOlclYhFEVsghMbk3R7Mm
eKHIgcVamesnzFCJEjwspHm6a5kCDCOoZhd/KaawbmGcUBN55+StJ7VU+Ghr+kvx3GtCyPm9JdPv
pPfGRGzS7NLm43GcpCo8T9WhN69vw35BbaJ09OUaPKeYStja+utSRsYNGd3AXjMJrX99MGG5evv0
RBcaVkQxZg4mC71U7gF4L5iu2OhlTTvamEdINhl5CAUDu6SLeZv/YZ9bl4dSB4s6a5sn8FYGezzC
VWixpBUlkLPMltIEsWNegLTrPGUBlcklz7QRA1ffSI97Eu2U7o8DB6ZRnZP8RN4SVUXtaTJVW8fI
sjP/kuLMvhXFMz670fiCi5oosSOmWfNKSAI9PJgM6FRvlVmFsv2bFYPJCWq17DkeEk3YO7kSEEOi
/l1oRnIguB9kHzp/y7lQ2CQTxixUySSA/+fLrVrzkX5/NUN7Yfl/7xhi4KjbIQuHvHuL0r4v+qHJ
QFsDUH5lWrGgXuMYyV6eMA9QGwtf1yh9ewgc9lyolAkaE4ahfKpXdfB/kfGmpwCL/Vv6sfmKPoKF
kl1fXYSOUdd/gf5dMeNr5kVr/j5ippBJJw4GwwH3LpsQ7yL972rhbreQG7i0NiPUL79EIMN5xbNk
qXuqN6t/V6TFTYQoBZM+zYY97UvtX/s/jSUsca7flcYLu8eSUMEFb257utzSWN0svae8w1QsFkd9
5Bz20RxQbkuaGEyVGFcLaldW6LwAsZ5RKYvNZ5VGbx8WNe1oMTRFISJGkZjajL4LEj+cUDq+Ogmh
hl/gbKIQSIwWiFkHrcHW2wZJdFbFRVeJyUKyB4OBLfaoLb0sIeTqXV3obZ7mbVwok81JETia2yb+
hTO6tKudRoKsEsDbTJNddjIJ526QE/3pMh6MtiP0hNA+Gn4hrLLz/GVtV8lz5L52dn2GnEXNz2kx
vi8anIAEDlfHI7VBShIJC/J5T328gDrkvGPcdsXBwYDYK7fEl12vyuojt+WwoxQ6NQtDFH39XIud
1tlPnn8ylAnDti9UyjgWEujbzOQ6zozjdZWUlr2IO6Q/a7bZw4amp6B0eTKDbBPGmMp/88Fz+GV7
+44Am+9EvGbjLb7Iz+E1RS1brxgFb98NI/rkqFqwWPZ567LLsl4ieQzliG/OkxJY5m+BdfHQAqVK
z7Xph6+48NCtD9ehyvT0NpErtfUgWHAPIGE9wO8VR8bZbGSJ34EyCmpuqcv0nzZ/x9/MigpIA8Pd
em1K40dvycdEjeOM0vtiJPV1Ox65O+cwMA60YKWc79fHwQVe34yhChzaU9/6gIRKm6ngMR1/Iy63
bPrP9ZeM7afrDCA6CNwZ5oh+L7jY/kjC0Q/omaC5k3FYWfx8CQdNWphPHi1rwyYVmxK7zp8pc9qQ
VMflSPja4stvbyLONE+dLzbKz9A8kqF9WoephgXFxXKYkwyZlBD2TgLVfACIupCbPinz8A5HfJ4q
e0NEthUhGLoa3ReQj3logndu6Lq2t3ObJlswh9AEcaY2xFzcF7S0pWiX/mtkl6RAJJd65JoH4KlN
5GiCCSNmQoobMwasbbKexeQFHHmYfVCvsweIe2+BCzuofgO5kqRvdxTKPPGPKgDdnCjSiWI5KtdX
jGjT4fHW8d/y68AeuXiUD0T1f0+bldWSO8YxeWa82lwD4uXA/aOgPSg2ZJDYYTCqlqXfgIy2zBV3
AdiPGsklFqKNi8gQLg0LUkoU+m46RU3Sbxk9X9Gk9q91wKMWfO6Zp1mE867aQL04Vm/L27MaKB2p
Ec3ySG6SHneCVdjWDK4oHx71V5gDSfLLC8oBkJniN4svibxauXNp1xyCAjDrx2lbhl1YCvOYaeAu
5fw6SB7SADoNdDABSNWyh84ER2AurbYs9gNscM9xpLzYdt9dInoRYTGGldpBoOhTcMjSz9plZk1U
4tBmPfHcV3eitpzt9s5XBpe4tgkh2lb1V0p0iTyPcN0hgpmywxvS1fx84LARpkdVKz+68AwWHDXC
iTuaAoKo7Pl3AGTHg9mfh5DgCTUPMYdV6LJFF054Aee27Ym56N6dEl+FAiggLa6JpKUIRGL3AngZ
cEz0oidDEciE6wh+DQ4PUmPqPSx4lXtQmQ4LFLt4tJgOzFpQGffiiRa72U4xHL0KzlPUqF4YHyOM
er+Qa8uI5oFfiU8ykFBWiBAIZ5O4dxCCFDyvPGynuv1ldrXbcVeuO5llGynO6+qeOkCpiNBR6fxE
6GsdAzPGHRlazD6x1AgffN/Fv8mw64wJaHYPcu9XO8yTyb353ctKv0fPKHYDYK06Khk9OiXYgBLh
/LQOqGxo1GzxWHUEQ3+zxl7e/javnHLwJuqnWPYxxb3Sc57AJSI/eTQy2bW2i/sZE+J2TcjYKOiw
X5LwFjXhYTyYM7HNfsri9MGTWJnjVrWpSjPKWsSHtoeWVW/33uHd3e+yddY3t+eBgpNxcpDrUCAf
cM56tYyk9zrvQzYTYCD2l1GKqNPGwdruVgXWkss9tAk0cDIAu60XVkrRZ8dbyJwNmoEV5SRse/83
IDsEzTMwrkZqaUATdcy7BPG/oREDW5VDvrNV43suheiADptpoTlJe+/JvQXjlpXT4wKUPbvEj1g9
BHjt60GNFztlPVvgXYuCrB3ph8PGrUXPLFT6sBzLEu92TZ7nNA2puHO/+MwTq5LSNgDwDcRbrmrB
BCtrVNVArsK8yZI2k/xVQBpRQuZKkdcinuv3gMRHvdjMsjcbrEAuiLhEX6KdzoyjjfAbsuMSeoL4
YC3+bPUw8ueXEPPlfjzjdRMnndpATILnj7HP5E2vOVO9cy9czHiMIKVWabTQBQiyfoVmXIqHoXXk
z6WC5mWRvjFAIjZvoId70DDqKWyk20jWPN/w9Zwq1YW9Ra3OxmxQXNtoT1o67IQvknbRrH6UcT8W
GzY9xaGOHWpxsVsdnd5xFSg2OQEA9oGBNvAqbczjXlnwpjX2RQD6etNdQFwuBcQl9SQRlPkP+F+r
ByS2Sz5qOqyEVopyT1W87HsxwtMEhCUoLe9+aL5kfRDvnj9gLdNDEAvU68f98LaC+dM3jAcz809U
Es/7yLfB54Jrpe9QZtfiTCNhxXVAhK5Dvqv4x5Pd/3kFEvRFIMAL5MSGwBs0OiEPAdyD25UVLuCS
vBvaR5kjjdokepraRu8l3e3a12hQvEcXQddTxcDE7IeoqJSuQfGxbzMK/gUZdzL5ALcMsTU1xaxk
lKfkPNTfifn62ndZkTqca4x80A82ZXSu56+NbbWpC94r4comVVt3+l6zAgDTfpQ2BnvrQHlhE3lH
pTfEB9gR6PeWxs5jqNiQ5Qny8IYmSmvRJbTRNRVoQjCV7iBdWOyr8ngZ9kpBEGfuTojMi32uL3tm
nglV0x2q3QKMPBlTxvsVobMZdVPqhvYGQEg95C4JaounG1rjURJTuOUpuD2y7DmuOcNs4i/9Uhk1
fj5F2za47XRw8Myoa7/cc3zVqNrLel7p/duikG4+ZCpQCPKKItfmkV9pPlBUFvKgnquOFya01QtZ
Uvm849JkqbzSyquLhY5hdWKaoTeTxXG54hd7N9cfLLeWht/xFJzNBJw3NBk74vdaoQYs91IPzJGV
R57WQIiax69vnyOXNQmj+YxQJ3rWznvqKb5AlTswbJjsZHpjOiNrf7N1mXOwMUvqm0b+tzXSCAP9
zW6jUlOMI/DMJ7ZWsYx+XFfn4MnRhRi7oci+2FGNO9Hg59cEeHQdaj4amPUiNm1sB79jlzHBNM3U
A+z8+1iyBewF5UnywzP7n9jQRbjxHZ9o/EItA79BqaO1VD5dbU/7M+ZBTwto9gG5+enZytqoEjwC
x50UjTwi/sz8gY/ur6YXpgJoVNKh5NUnY60L9oS3fsUU5xokrBUQ/6b6QSpjG2K7WV9c8PIrW6jp
5trQuLe8bX8hTndr8/w8Tnx8xSJ37aVjf0JlK1fKL5uvfupiDpBMcE9X+cAIXRb/yk3R/DarTYqp
fNfCBupgRv/V2N8+gyOANjZ/dC9srSNSFmN3YiOLWhW+2Tw31z6kbnaq9hL1LE9x4SMvzMcOi2UQ
kvnxgjcOwvCj9fNX+4het1DNtSuUu6cF+sOouSsI1CFWbTQA/U90RCmyoXhU42grEvAP8vlrKzWH
pU4/IhRfrWwUYNZzj2XQkbZdmgTKrUzMsSqtJv6kwSFUGvtB3IbIVxWFaZ7bBMD9m8zKxsjDzri4
A0JkOf9wBp3xbMs7HqOQD8a2+9as2g2N2GZaHA8rQdEO7c2IaDpEPiLJ+zJF3FPJpMTo79fKqoX+
2YsW8UFRqqjvYpyBw1XO6z3pprTfBuHBIb9mvmpCuB+5o4IpDxN4Ymr4JlABQZOnZWHPatg8n9z0
Sk6sYcMvFLE/P1ALjVo+LAEYvvMrA0yYFG1HfYIG7eJdjHJIPqAo8ZFpyXrGk+bF8ovWAm95fry4
kz5KeG81T2/iijTab1+gKDcsb1xNmVHlDyoEqKzMFNe7DxBg3P/cA/teStsR5YRX3ZRaCisMbCug
6/Y4VKaBSa9zo2ra9hvRdshVIgv4lTeOdn30jy/5pnrWQA4Qe6zCFOAb0PsFmciBQtPD7DcknnqU
EukmRMtJ2k4QnkJB8NZxUTmT/46bhyhC6sLLn2qBvPjQBUDmAARtI1HKbRQUUwrSn67pH12N72fI
cWPWigUUM8/+RY3miF8paVDcs78L55Fuw0vFeSQSZr4RUxRoN0xaL/UDwRJIxz3J5TLB3tRlS4C3
qtxJfLqPA73LINDwZnoMkzc77mb4CEJTdduYQ6GSLoigdzt9j7jI3E7ER3ymT5nM7cn/tyh3pZMI
S6qxp0T4FwuNYUAeDASWOYDSyqVCX9JoELAXyQ6FBXgNALrHQ0ClrTSP3MlT3pamvRS+2BuY+Gau
gwbWfu+wTU1RNxQJJuYHYzzV5NmFqFDuz5S8aml1lxZ13kKreFyiX9A69ZjWxqDQarAcptDNN9LT
ByrYorg55HqC3VgFywDgMymMSr37rq385RAKcE8b5r+CKNdwbFoqLpkvnKlgPmTqyhuPcUxNLRns
Sn5imLkQ2s9lMTEOPaLry7g3NrZR4baUo12woZ3cmZoJhDqEOEfEcOs2lwwwRqJyQtWHxrMJ9o7O
BjFg4mphwyU6/vuMhg2t12BK0N+gC1JXG514y7Zb4O10xge26zpMTb51mQnyFOTzmGVe2HOTS6WA
0waK7yxYOKoQfDdc9R5A/r7TFdwbLTnQCH0rG1oANNypPnWqg7b5oSeP4N390VdIWyDxGDYBZJzC
WiddW29cPP+8KE/kTbbqnYSgv/PIwpJ7CVRlvdiCSjCvmTtXgYDYIQTyD75SlODofE3WUGvQQk+J
uDJrQ7CD5/jc+uWqnHzt96h9WXgpr2qOj0CI3nRyMDQoj83HL4dC5p6d5iOZENqd91wn1wGnufeh
SFjbhJJso+vCpyKSPpOrdDCW9CbVH92EztAzvF7OBt43VOWydVg4losA10SycP2qTRbW4m0esxgd
uHN/4VT3Tb+jyBbkxvMwi2f/HREU0UZbO3tw56HAGEV8yrbGwYsxM0E4op9Scq5XcStbPIkzYHba
J+D7eD/Uzj3THswMyVN2mm4VtOrXB0tE6jFth0jZANTFwjrnXy0lI63G366xjD3NeeBWFzzLfxYx
e5QQNeXBkPcG6vbhWBZFoXGc7A48mXzoa/zm6PY2my5tXzcFEKbGaM5DLmLAzQEZpu7xM9xlb9OJ
4ioSGhShp0GC/sCnI++CFOo9KCdD3BthUwRSPGmGCTfIiK0YEtQjDUc1Xb7ph65pU1SCtuGAFjs8
N8lRZ1KLLztooBrNAvcwodAGA810nDJUVa0jlfh6mZ0oG3vS4csn0sZLp6Pq0kRgmdPD9PSKaSuV
MOl7URkWVR67gPgl5MysjyR6EaQvGHfWiVVdSyV8fz7aAsrmn8DAG7SDYKNrFACRwK+DYZSim7GD
RXgGoPSaMWh/N/1yKI4Dx/tfvnNRFJqn0IHMfuwwwSlweNUNYAcXNcIbvYd461c9+Q1VEW8OIQKE
HhvRExlX5mw10RJjYqrjvzohsVJj7tgIm64loYpioYfgEEsQJ1vGlu6Ly7kxKmjD5rBbXsxuIxtl
RAcTilReIlEv2C2Lc0cV7qdDYii8Ln9S8iamNQL3lyPjXfSFG3IeNgGkjKMJMEX1AiOgyG9JZ7s3
XYLchyrPXAFrtp1zkzr3OvxCYB5PWzMsWYjdYukif0jJ3pZsKtn/i5wQOrIn6jwPEpj44dU1/ZoN
46bkoN72GubJCPM8kJyorv7WYd5Je1ctG+gggaegaR+M7+mXvqUD3kOujbOpvFVAdo6chco8FUK+
8pz8+dkxr3TgrRiHw7lwkx1AFkaM9E3Dn9BphYBh9hQpAtL6kDxliO5m/P9Nshi85byHwScpKHhm
qWEUZKHloZA0is/CJtWh7q4qXnODD60CjIm/mzD9ZsV1pRWXB2hE7o2le+5ri++pbgjemOn4+w2X
JOsDyy/UjT7itcceKF/qJPo4RQmMaKO5tOPP4u7k0B3RyHZxY1XGiBOvkhys+jSCo6CSOKgykD02
Af4EWSP8RjbAUXBs/p+vdBDZK0j90zGDf23I0gT6FbM4znl+mtVyUVXeqWaaHVNaxp6/3IVVxJqd
7XGCR/QroHg7yt4Rx/4bVdrONqW7hrth7cxrusx5ck7rZluWAVZ30LzURHAPSlWv2CCKAEsq7bQp
NfnQR469xY9BwIBkAwsz+7kcM0Jpr4QDgJZA4rhrxlJL3nNidfwHphtXXDuVmofYS1JLtsu3bH4N
r9qybGfRjpIppXHciJn5yT7XyTi1TRQFA4NCHnidpblHBu7HNrgzUZVYNdwd7LtXcVAZzOEHTrAY
z3jlM+mqS/4xnNm9tpRCB4PZuIZBfKTpS2k0e4pEiab7iUQpGYU2r4mSbTiM8Nw8r+WfFLNpbLFH
CuZL5Fuda9syiEbrt1EKvOFWGiguYw4Wr6GAexw9QSrN9CfYebc6Vnsoo+8Uj6KsBSNY0KsbT8+I
M64IDWvyMeBtvec1GkvqUaiPxYArPEownOwXFSKNnMRA+cD7rZZxqNtNdAAmxWdj5mlJ+NSH+36u
w1UGPRgluRBRY9R6fLF7NwWzCC8pKD82bRknU8Ppv/ZscMq99s2LmLJHnGbQkL3yNACVWN+j3H4p
CKY4O24D5M7FvW7SGUQ5EGRuPhhM5cpIkv3r0tpZfwdYWUYcZoozbcwWEwbt6bRMslGPUFVvPaGX
RBFTgFlrDwGY/jElSySpM8rieRt8inG+meXBJxfcjcnAuluRLRSQyLUtxHOh9DxJnxRPtr8hkrfQ
DA6ZnwOuDp5MjxxKtGsdyZ7XS9JhSyw1UC+h89fdvhJ/DnvuSv/gl+ibvrKYISbpGbUaBTX9FB+p
MRFEcKdwu8yBp4DmSuFUGtKeFeUYDa0pYN4jD42Vr2kAw/GanrlmI+TsVm3dMLTlVyyawsZY5QKa
BbpYedaCmkxQbti4QmXq4LZ7N3wDVIay0+pX1x6W0Bmco81U6ITkKXjdowxDRU/FvbDb+Ujdo3AT
0rDYFLLmHTJNQl5s9EcjkfM2s8ANZleYWn+LOMEWMXR8YkVYDbLYcuexiZ0MjiOZWhcoUZPIP7fP
lFhsg4FSge64CQqfAO0dV7swC5zOhKRY70y2a+GtSr8dOJhFtKlOT2qTtVq4M+XZYC2jow8C0hKx
u9UtRSHqZYgW7tfgagQ0IPGnEdaKlbS8r4hJEB2ySU3gJs9cTaSM54WGwD+JBXSFpQGiFfR1GiXF
aLJwSpbwqqtolGtircilRDtkVZXlzxmMPkje2TUtMAbsGMpb2lcsla5IP51PUUp3kdMZy2NsomYE
V0XEsBpOAKyy6v/yHhBVFFVDc9lL6hYumPl9jcBJ/TrLmDajAfIwHdstXyQrGUHgs9WjelVv+TBM
ubAB8OwyuMyhuQnzChj4c26gDpc9z11BVY3098O188quK2DCj9deTvz/YHNms2/qopFW9QHgEiKm
rRIX8Y/dkxFvDeJwAD6BoPleA9TQlHuRoKJSs8xsYG718ajK/qnRUO98kyrDCMZ+scvIaYA4oyIA
qLgvYx59SJ8Bz6TSxTwkkGDWULR59SdkmBoYcvXrqdHpOj+dqqYO+FkpP3SO60AaNyNxyF6lbYyL
KuYAtVI9Gzuthg6qDqhXJwZ7orY42QDr97xqwFLLqOeBdcE6oLFcMB9PnRAL/TlAemBynbkjRGTQ
qDRqSJ04axT/utyYAl3ueDSlp+4DSMiTsVWUWJN2PGnkIm77srJyrSfRZAQEVeRVRepiKDHBfH/r
Yklaz8On6Us7U8RoF7OzbSNshdgJ74YILunUtsGSxl7+gM310y3dkq9wDDn6lpnCxnSliS+5a1r9
f2DeqIKvZLXuJrRBDZJ7rytIvFHhVloSabbtxqbxftkEewKSLPDmHcXq22X1KhiJj9D0fROl64K0
Wcc00+exT0ZcUrOG6WobEcGWjhbnZSwAsLpOisjnuaIFTlE9is1tvzPZiL8PvpxZiRCyj0PoXZw6
s4L2OO5wbVwtyNb5fYsSWkLb5JaAa4A2OG36RowX3pUjERRsPc01gJw70e3eqHUPQMEvl4fxac5f
hrtiMJn5I4UBfVqnSGz4za7jKveifNPGa6Oc+AyTlHiZF/SdOhzHaKZP4BAhfUT+WIfXQEHXvrqj
+tRqt92/NhGjt3zHiAd/y7keQfSRhmDV0RzQwmCu/V07GE4TYpFlc2V7gZr3Cs8pRBkRuHO847bh
HoIgq6hDktqPNDtByfplxLuzS1HZWsBIp47UNY/oKZR9ApwCo+1y5LZxdIW7TxX02qDpHepPMiTH
GNQ1tupVjhjjJIMoudT7G8GEZhJbO1RmOQIBqzgndroMj9+nSLRKRGNRZ47Nk3aMg1h2yyAzSSNs
M0pe590pkO/fpNG4Cjul4Tt4xV9vfinhMplp9VXSeXMmDzPyuJbpw3ezJUFgRgaT/+t/qAGch8th
BMhZEWea3+tUsjo0DIz9sR9OkWBh+X9TWJDdcG8DdDxi5vgbVPHwimKjhkJwXuV3wFjbmHeHpRdN
FF5hTJLkeLwGGqcg2YKT2znxvEUpH9a0L+cg08s6cKBLiCsoW2M4ev7asrn5S22Mjlwq7YTg+G3x
ifhlbU36ZSje1/84gjOzVFUzQyGQCChbRG6orOfglmZ4BjdX6m+J7KEBSg1AZYY62aFzEadcwFDG
f9msR3vG9RZQde11CdYWnCgWZHQPb4HW6uGM1SZ9ALHh3GkAVvnmR/TvjC/nG56+xC9GTIfPR15j
fx23FW0TwEN3oHvIx8536BtJsYATsSphywJmD7Eb4UIj0/FwvSgRQjUW8eswFxFKTgQREM1zJ52L
VtcPIsOhRKDArsdycp4gUUMbf4xaD7fT14HSbQj+Fx618Mam232dtISc9a1obaJAVoL/Uu/DAXdB
idBCeAEIPW5HdGUV2Cc0DVqtFd8HhsYcoyqFFq/eJ5GWxRQ8z8bfhrWRBBMTxvzI11GJDwAoI+Lf
J1WFuuMUl19aXIu+BeHXHa/j/AMKVQ6UAn2Z3A2cpYYF9sxhVuZTzc+r2zweKHxa8yT4GY4fQ/QG
uQPVFXzXtg6TZM8CqHjb8RfRKtdYI7BBue+S8G1xllu4Frsv/H5raFE+CZS58dNy3MHCD8FDFKEn
Rdlgu9xhhWElja9ocfZZPxLs8AS9fqAKgxqYhj6zo4faDqHBbIHVlatQe+w9+cZX7pc8qktjoKMM
OVodsAld5pz5/cdY2R87cytYsw99w5+c0ygfVZmUtcySiEYOzJ/PQMi2DLFWff3taP5f+tFKcHSk
Y+9PzSRoCv+rZdz9Oq92sbq+CAmRCUmO0mRmkivRRouNewwZYfsSZ8WJ6WABNLp4AGXyPWVH3VNv
TEd3daT6gUM1MzbstWpS2T4ij5mCt5R+W6bQaj5zqCy1VvE/FiJu2h/nXm5BAPkpi0IEyuE8ywqK
ZWQMxlsDs+EiMtF2i1mymrts2TVL9cg7OvrcnRYsbsWvwKnGAkotCwcGeKjUE9zX7uNf9Y6SdiwG
mBRIFjEEqBVphPH8lif3KjRMMdof0vsT7Xn1INhz+g8SrVUjBK/FE2xQGF515GRG5v9grJQvezYh
BLoQxWmBF2RTUt5p1dxuVUFpwXXPoJH/EaIVqTFUn7fyaM6sNqJAoVaT6A3mYDWkWEtFnoMEdmK+
I96OHlbIIH50xzXNKTXm1Vn/l+kUigmgjEWSIWFonOB7nuX2P2FnEsP2BWVIMfhWMmVzzPT7cr9k
eTENu8AnDenv0T2o07xEuaR6gDHDW1t/mhOeqpplG3SRcObnn3jcg3O95Bv8VcM4ssMwN/aV43Ju
2t/x5YISCekYbt5X2xi2cM2H/V0kMunLwmu81aRm4MAm4sVUZ4+q7B4OgYViBTSOdUYueXGG86Oq
hQ854EfZ91KBkkMg4PWgA4brTVb/9BEW+6t+LPPvf1h+EqMCxXHTwk5gcNJ0S+ZqKo7FxsdU5myR
DoPJnstUb+OARwzbPnurBdhEtyssDmrn9n78lZXR6w4CMjjVOOomTsmzKvS0pG7cJmEwh27OVt/B
ecSYWw1OnNzLP+QhzneYBV3mQOTlq/2aLKuGwAZtMUU/2JrHJDqWvBE7fuZA4L/SZjWwXnzMIEhA
ar5iseFqAjPZYErOpSN5apD7yKl/xwomTI1PtUfIrC/ldZoAuNgsxeA4BgJwHSyIAx+qHIPGhT1T
ECihJKCYcCt8S9ix9cYYEgrpoPJqvoMn3FrGNPmxIO4UMmP4339AcL91C1LsY+NgMkEheMLUSsdx
i4Ep42T9GnaoxHukNXGd2RCyFuHSwU1VmVg/CHGzpLHJJy1BV7fStMpWrena6RMvKW2h7RcY0r++
MzIjcRo+zKkRENzcj5LxNJxI004EG30kdUJ0KJhH0GHFIiDh7mjMIZyY02tAPGS4HtxkgmRWGt/J
AX02UFxVcMOTRwvd4uCKvNMEdNmEF61P5Ogu41qv5XmNMJSngNWDhR0jfH1Ke2U/54mhcaSvvrrj
wp3AzFyF5KqkHXWeRcwgBEkwiXHwFcQMVDAo5EdF3xGSmf86KAGqkD2HT+GeFQJwNGH80VL7apdK
y/EQr0MMexRSzv8uFFnCzSkDRad75EF4k/je7QLSmu7ihAPWlqyn5sw3jw+kachj4E12Uavj96ZE
sSw9VbGo1+qgIkHjfQC8pzAkQekujxjCOF1faq+/TjCz9izZlOou1nmlPAqvJbEdGW0kzvx0BAbI
mA0j2oc52ixsMfQjsEyrd99R49SxnYf8JNa88d5vn7kDBRGfmF/ll1HfkhuPfVA81S/uwn+ArQYB
g2+elhMjiKPwJIM7DuSxmCRV5ecWbn/UuUuFMuyhIljaKDiCxIwHxPOpElSUfcVkKa9qj+3Qupy0
g+YVe4R3L6jgX6WBco74tXKLtbFPCudjIcr8mHgDyS33tvuqwnfVk9O6ZaJvL/aIBBbJXxWL4gLi
hlQlfk+1x4OYEjIPPKAVgBd9/taC7KV1bRgS6vHY7mCGajdrJGbKTdCiwrYjS7Xxwpiytkc+YTEt
O/2CDfmI7PMRuXgMX2z6WzD+aPdtkTw3PL3AbC66zv3r8YeBmYpq5piAmkFyIJj7NEi8AR3bDwll
+LhzEq6VJrAyxrivxvCac7fMC7Ak2QKr1fVh1vETnEVJV1RlgvhsGMpeF61n3ZuilnGKS/3Ro77D
fYf/ND0mqPz1K6A7vxOUJEroHYATYKvmMnZtuzhN73QtoNzVi9+tJ4Wo/QkIGOPZqcD23MAxkpZa
CorlnG+tdKfo/ZTvZasxo9MTXNzDXrV4tq5iW25euU4SqzFC0ffibW2GuOdmCxw/BxHnaiZrtDw4
foUuaIIS2scjhA1vErr1qrgH514aOQGzkUjXhqC796TVhYRx77USEXf1ulbutuwbyTg7eDlMrInn
Y2HkA9yfcGsohVLZZ90LAh4/S62wal1EaAb9EiitJc6VcazyaXKVWwN0hyUg3zpspLELsg9hqvPt
UdU9lclC2xXIrE8+iXVOVcUD9msiYr99l3M+gRTcmRaboRpS7QOm0E5H+KsbX1lmoZrHz3G4XdFU
nv7rdnkeeJt322qgfvyhwr34HvQkWd8jIFv8zWfJLH5QseinitnmGhxZr4Gzxd49/NMGFIc8VEJF
/Rswp4kjJlFNj3RU60OMtj6NVI60EidyMSIssueGSrR3wDFENh7CsdbNgqwL6eg0DIzYRknO4GjC
h01aKvPppzvdF5CV5Filcfpl8yN1tmHKhS4nIjo+Pnqs/t1nRaSVs963nOilWHWu3eqZ4LF+Rnl7
hsTwovi3vMhetN595DM8APqgw05teM5bTe0KdGssUnhVPFqBTZFb+wk/AG+ARaIaY2m4b9M3joeB
q1FH6uD+zGOlEgxoGLckxKmwGLT8Y3dob/eNjXszHkeLYOMb1IsXb5Dm5VhThc0fOWZHL4gUdiI8
q1BGjyBnOrQQ0DSVR6pCk5ofgRWHvfAiB04L8V++DtPi1Y6JvOfvJgZRr4HGu7ejZ8heb/AIz97G
uXd4KNWhHOhKF6jLGHdn9LFTt9XNo/us4h7Y7+vOKyU4rXenCOFchbIm1wYB6d17x+mAmP3Hzyuc
evXndzV0zqjFiVYzvQnWUF/VrS/uFqb3Ur01bl7EiTLUoLq0wPyEaylwF+aNZenzWfUczs+8a22S
ZFMD5FH11Ios844sJ1TivUVYa7FLhHjPnWa+6KnI1qbZ5qfZv98diK9tJFLUNiU/9M/BkcPjwqma
w1S4A6oJd4dh0UjGBDiyYxKB7RlqgtsZAamTug7v8bqhnZs6QZVpAk361/9U6Sz0vvV2l/5sXu/d
IUDUvN4qJXzPXoh+d632DCRnU4jDOkUZUpEQKRnTvOPi7kmdNjjIM3TISYCEun/BgvhDKM4gb+Qk
JOFcEtBf52aB4l4aKw+2pCffa1BN5efMGo4blkQQqIiGAwsVAvQFXqlEiagTmGaRwldqOQzmqW0l
yKfKcAocenjmYLoZ4zoGhfybsh402oReN5w+tITEePikGr+WdYTrzthsX8lDfF6uJYKnqcU8kvGD
/UaSgeWOIh14J8HgyluBkJAolMMRy5hLeKlYpnecnX7IJyRX435cyQqpOjzbckK+IRzE/hwbQiH3
DCnWQQnjON1GXYSwjrS5pjHqsSLLrzVfrG5c9beNUo88H76DKdjzGU07wpZVPZE/x07sWMDYkv1q
H8gCAULVGjELGdPKFMrM6UXqecJOLFWx9Txf1zpvIotd4y1LrXNq7RUsIDBoqsW7DGQAsHNQ1aZq
d8QLxfMVLGiRw8dcd7pF96DKT4ocIBCniWnBSG/VGAPOwAubbSLG1Azlsk5RmJP0GYERbiIi5r3W
Q9WgelVG/MaYb5v7t26qw+33uWP/jqP34Mn2+eWjDYs+TU8fGvMHabJDJfk4p2J6Odkt+XI50tF6
pBOdu7+WlBw8MYJueZYFwcciCmrheKahII0z95BXJZ7Rw8d4VFj8UtjPtLAwzcrsZ8vipMBhXk1f
51CZSxoj9o3LhAdpK6f2KieFiV+muDItRDBofMXxdNgqXDrQQt7DkaxvOvPYZuC6ryDEzZaf5S5N
NUrJRaLlp+SZuBYKAMoFjVTtdxLRnt1U3X2NeO+UJD/R1zFEpH0b/wJATtpCOVL1dD2LUvaxlN1s
UCCM5eFBXVwsaktU39NH8sesnyeNqjPi4GvJXSYfoOu+k2TPu196FCHi4Rqx29pp1UjaygVhTnG8
7jxYEqD8xBYJBp1B5ZeOJ8gLK4JvIpJvHubeGDbeycE1R9Lc44QwCHxuddYBQnBD/J5Y8t87SxsG
4Q2kvXjMDEQAJ0PHDGag3lSOdnoJ44N9Ht3OdrM/qYhESgHZc//s2tidwSZAHKdgdoDymMwCCx3B
iS28WuCh7MgiRYzIzSJC1TAvcUvPjQYvBk6sZYaxmkAGlCxhc6jzBg39ubTsUvmqzN4SyhHwU8Qb
Jevq0y1bibJITAGlk68DlvTgi7qvquQKEUfZupKUTAMWTe0ENi60sAnc10MjxMwzqriVNVlm3dUN
QnWo5hjrEM3qOc0hmm5XPkfinX89xh5drapVu7BqbW9h3dF0ZatKYqhfqSWGLnRqGxHgRdXpQR0M
GltqoWwjXZFI/MWIB6TyVKoS969G4c//4r7vc1hvd0AGdmWQgrkq/MTDKHpgERowI8655Yuabr55
SoVTFHIJLhcWkoSMHEOYbRUBH/t5hidqfLLEe/4YHLXi/mXjJjF9hccG5exCjXio7yXDxRG7hnx3
YuSoN9VhiA4pRYudRiRpaDM1ZcuqzGytyzOIjJXl3fjMq7aq6TXK73ibInPyf01ucNT3bIAQKCh2
STitm0G7NK/IBcGlikjXU/K0AQCpzueisrFDLrNeA82ef8I9dG8zwhLwgxgzksCPVx8eGp2a+4JS
2g1Ezt92zfvCmsYKrHj13IgimsVltXGOIP0xnHuFUHkgWICbZYcPmjzPQNH1NPm4chwOdIt+qDJp
M87Bp9VH/F1tZKx6LxLbEC9K71MZAt5w5gZ5+Lrhxn0fPU8YI6hgcXOaas0YxWHqQTar0wxEotqA
ETKZcQeKBS+pGeVacGnmy508c1gyTeo57eVGHm7jV1JcFYttw/W/zPntIw9J1wUdef9wB/FIjq9s
tYtkvfzj6O9db1smGjUdChKq0HFvQ655JW3SegNnBNGEv+UJYnxzHNESC0da5VGexdcVyT21xYIW
3khiu3UeFTuroZ9VBY+KHfILfRQu/BoBdhBXMGK9Qjy/vo3S40Dzvridai09hhY56xs8X2p/EtM2
hZud+fo1ZZfTcQLSOnzqm0FtbDX9D5I1Sq3tWMGR+EJk/LndZzAAi7obhGj4rUFYKgQayrnJT/H1
/LgAbo+sc4rVETSsBAxokCoNwss63bWfF2vRiV/FScmwbOUXGIoHkoRnhtz2gtrWv7gSK9xIVumN
Q1llER2d+D6qA82JdDWBWWAj8ph1OSoXEenNRZNrcu2VUes14Yrj2VCbsHRuUGmDGPBuT3tDmSiP
1YsA/wg5dJJWY3A8ulhI2JUX/5xlCuM4ToWm558gHDr+kUiB100dz0U+D4dzl/5mUrISA6Mc8bxQ
JQKQEDu/ZpPBAvVXyMlPIDGUyZnvsZMi/bSPpVL1ikH+Pi0K37eGzfLyvMNtahV2H5pQZfA0ZdwG
4uu9GNT0FnoC90EEdfVIZPkP9miwURlrZVLxZqsy6+w+pXf+oSlOxnjQf34kOPwejYCLbh/LKrf/
wreFghPuYNRrUSybG1/pinjhORLC5OIcbabkxlhiR2N8ybJmSji8yqqDh7BJn5usg+tuxxIMbibz
yWri/6OcEC/Ko+sfe8IO23ud2DfDKfu7e+pL/Q+IyhlGRzkR92wxiZVLJpVcZh6g9Xo+TEnQWWlA
ZTBkjxMwU2/mP6cW8ALy91YHNNBIj2I6M+nFVthZ/uSSpxOY2CKd4FsXRtOYW5v8l2WM7ct5L/7S
lYNyPLe4HyQdNrPfQEfYhHV7UC0SIY9dIOXbnUCll3BN7lpZ68tz17wwX7uS9ZieTuOLW5S5KOx5
y2OobkHlo+TeQyAE0qlfr3nZ+eXsOlX03CK8X1cOWVJBwlycAThLe3c0ZWcSxEhp/clnMDiH2lnI
d6WoTnsdyoRnxxMXlfqsCcVi26gz7QyQura3FOLgrqhA21tfbE8semwm3nT7Z7pr6CWWGR38Eaem
TtQipedIiVfkDo6NDCsp85u1GH43EaSyniDcXtYNGDNRTYIWTJWt5BnNFf2MJ2cHlYNjPe7KEUvD
nPht1qebhvB0GrZoihlvsD/e0Pf0nOlCIo0T2eBs5vKsGsRZEDYM8nv/H+oRl8dnyLyldG0gU3LB
NgZv7hA99DneuYmftVc8/c0lzvVcpw7DzJp8R+sUI78tLzO07945Hu8E0rJ6xK5uF9V+b0pK2bOC
1Tl4jPxOAsJFMF0V2OCLnJvWQ9fF2BqC5pTvgkoIFkd6r15Z/WdZVEi6aCORjD9kBRUMazAZtXCb
N2h4hvxgb/DYWTdfPDQx+Cz4ny+gUJ3IAtjRKXiQGFDv/NIUVeN0RChCcPY5avK6i+iSE0GIqT7D
fZxBqDPEe3aRvycOKzwrK/HLUptfclAszNk3yXujhZfdZFO7rA3Pi01xSFvLQktvMuhzVgWwc8l4
F8joUtxaOxDDZ10ltjt9KlYAa36WwSJhjEMb2yij/sPXxJp8PxXiVvBoE7mwqLLxT66lYw9By2oi
JvC60Si9+o1tLe8/HJuHG+XvCUjJSAjjoODCU0Sqcblub3465Q/TVEqWQ+i5XyatZ0EnEcQ8BYiR
HCGPEvdoGTk8RejvHSNrmHlrq6q5Z2liZyzG3qsQ2CkTmpvBf25K0FH60Lpvdw77lgEnt+6sHTI5
uVpPOSa8VcieuRVJLK1CU6xXyJ7jb3Tn87XfWi42J6RMm0SqxYu4zxCmaily+WAFYe3GTmes/ZsL
ecltIVvyEbO8CP9drqFCv91xqkRdXlKC+b/6z3IHJfmRseMVzCLhb9TwYGWBEowvVM7yL7Eeo6+n
4Yxe6Ur0oATNXTTRBIbmK9zJNJr2f1A7aQnAa2abO/xScpoLy5yd4+XHItnBBRfckFhq3iBYhM7W
DZSTq1/e5jEdSD4G/KNppPCpp0rrUjwwGUPrg4Wjr7ohCSIk5abvDfqvknsRrvMr9JH2ZTuCxdw5
HknGUCm5X6bgyk8TGkvhatoH0AnpuOsir/BXyS/N+NoR8hOmIyAdDJhRn6pUH6rASfArP8LeaGPv
p2sQfBYV9sfKQpZXqKHiRFrStQeP5yZ2iWVb3sdVpiH4Rqowv2w8JSY3prKYPSc3mW/n5V0YwGgC
JB88bUFUnHRqkbf3DNcX3cKsT0FFK9jvOvdHzuymMLIXTj5CeSWiDpT8U/ZaJtqdBCnwOxil+ceW
ulE0fx1Dt4wSCJUFJHmzsyd05VA0dHOLxQGyVvraCFwMwlaedcjgZ+mSdwQ0rvxV66IYJk5CoWSp
mtHdN7o1z+Rw4l0v6cEYekonTo9lrSJ/xTFJ8DDFUbKhPBF45Vq9OJ22U6JtB6k1x3z0+0VbFRlR
juyFiAgyBIQ/gH6N5QPX5sfSuTQL6Gf8/gBoAXzWna+hoxm8oBj1pXPJqi6OkRSkjOnFEnVziDM1
nheIMrrWYUwFYGi2lcE54g38Ll5L4UTBPKp7XtbF2A6prydcsx+Ugi7KlV4b1r9QNpDrinN9vNwn
Kb0NVaVbLY9vZGe0NxXUWay2c/7uo7n/NmlsBP2DnLVg+6kZS7wZi/kB38Dotg/rZuaU3fqQKdkz
R/muZFs399SHfkTwxANTr6qd24eJlkT6hVM1FdrN5HYcTYe+5JNZQsFnBYgCbpzLRldjpH5bk2/G
yhS5J7ihUuIZ4gNRx0m/3K1CdtHZeiOLjrlijANnWZRJr+cC9L3m2OCtM/j5Ama75/AH5C7But21
kaNpx3oPi2k1teO4SdUdxnLNgKy0bKyAY7uw+NfXSe0SEDm81DCSGZMICbb37oC7ZH0ZqtfDlucH
PBz9dIqEJRgFf/q7rtIqAI4BiYbiAPS36ZrmN103/2mXrvNGOdgaADAI9/gDiIkStfuW2fJRYKJB
ZVSu72bz8gpUWSRje4noKzTmgAbiPfR34tswUagELEe1NFR8bo6+SJePh2S3y2Ux8dXCrf8xWA5d
ZZQTEviXFa6XTUu00VrGbkSe0JcpgYX+cGjD60KUujYzEI55Yr5wBiC+nH/UZ7PxDrCjyOJxenGC
mb11oY4EnN0oPh3wmHKW4u9ILcd63clOkTUfNNQP5xxsW4sVCDJ2MfuwK++0vwgdi1pAZF7rBeVy
jOtrjLP5GW4B15TGJgC5SxDdxmKtzKBYp2KZHU9H8ehAIXPvY7q9eSPk6gP5Vd7Oi1OgbCURhkF7
2qIOP5zheFu0C5X+CzdKfKNsywO3BjPqYc0hX5yBNx4MAArN5TT828jcTyi26eEyhT+XuS8paDfj
YklxP3T8enaX7NBIoGxZWdbZCUe/RWxbT7vLQQ0kbeyBnFSwKA/cRJVt9ksrQR4mrM35IQ+FdnJG
FDTV8HVo7T2rcfmDVJNyUI6ZzDgKNTZTJV7rCAYJR9ezhZ8pv8kdGDHPnpTzFVLVzQ5tSxsJhxFN
JVAyYAnW3wPFZLXCzRIzNejYvTEFvmXiwRMWG1YTS5KwT1fzBOnB7MR0ylMG8ZALGduiPFQ9cnBl
s/Ra2mwcliJenqck+iDO5p/YkEO1YigL7PJ5jHwSrv+mgAUdNenYoMWsd6V7OLHSgnPe4tPYn4FA
Rz9oobEFjyHhEUpC/K/L2lsxTazUlA9KfUOi54fwbSGPVwjspr4BxekH6dPVsNQZUdNtI9Nxl8sV
nO+AZY3raaBw1GUbNImFPs1cS9CcLYwjN4OJ5Vm2j7GXDYrEFpbSnvf49u04HhEAesXvMgCoF03p
LDQFFVZOY9x/Dt7p7ESqMitA5ApKMgZYbA2B9stECpYtFKwbfIFes4kKu2Mt1I/+zdyf5kS8b1yw
WZOZNIUL+weqyvuD9JWI0m5oc9cbVkT7H7wXJ9BDqATs8Y4Hyy5db1ixqLnDREQSjHIWjZNxMsEI
+vEThNVdr0zTMtf0185EiiKLytu90YkG7brRheSuKXCzSyLQduxCdDijZ9yFjJ2pmSa7pX6FCDvc
7qxkZGeT5IJI61rtHJtk3xkx4fCE4d+tNFFD4IhnHNevLdQPVAyeXPaRTJxgTTvZPxEiasmFax62
EL7u5t78Zg4iXXY5ydre2OOHu5sY814EFP10Ga9HIuAzlemQnL5xlBmYI2XJpjOCTtQoz3gBPJ/N
eFCc627I2HDNukZBzuoBqWsY3F5giaSEDAcTfIgpgtbmsjaeRMWEzCRcSIL4HXk30OEwffvUor6X
PeyURkDACrZT1C2cLY2hlnhw58c9VDrO5SkKwnwhxm7KMYZfkJG0FZujtyUB+FA8zG7MQIhGnvus
WkkuM2wNd6zFH8vE+gx5M9XX4IKTx/NCT3019kRH4/fGjCEiioTE0A9TO6xbdG+2MGKf8b4j58Lt
xTzL2X9ITEYeThQoRf0qGM8Vq4Rz7HUdKtpF+Ac5Y5ccjnC4y+IYwMkgjFSwZwtVyg818AOb9qs3
cmltehNiEGf5JaW0U70yqWX/sN8U3YfIpxkzkZys4wpuXhONZ0f0uS3zKeTGd6ByqUxtNvXORJaR
byC49p7lBwxPwiRjOZpwYXi9CUbtxXlhnuqhmy4XkcfA5Dhl+aq5/6TUL0L98fgDoNZoT2CuflQT
fV17XnXgDZozzFQqV6KIKVKrqgfCwSD7XypaurDeB222Xl3qrwacbvDfIFARt5XyjiO1ukUmhbz4
J+2AyKoLeXClGbELED78MhuGyH1ofFAJQztYvR87b2mR1FhRYny4VNafekKEi5BqAH9cohvBwYFX
ZWm6yKgjosf/53y/qVAfQUQQJdtTFzgFncglxJWSX1ewuWG/C9+99YfsOkc2hZM6IOoskNwzpFhN
/gdvhwhFTHQBCG7kaQjh9qBVGEKgXi+U1kBke7i4HF9YF02ec3lhjOaJNNOHDBjYG+j82+aCJiAE
Du07TFQ2C5zAgiQkDAlUw0WaGHxhny8CH3krBqzP0w3S6yR4i+7qqtch6HCXHTxJSyEdxhijFwbR
q/q1BKOG1lUWXIAAK9zfmgVDU3rePlVeU7ridr3Wxm0u4Wl4D6xVCk0tR1eR3HTGtXA2/n5DVpI0
kR8fD/1xeFwav1aRM0KdoB4SdpPZKriCWoGzt1Vt+Pj0TSgUb6uz7vsF78gfiTOUFsmxCITfWBEl
Ry8WG+dOG9GxJmgDbaTSc/gaJ5EEW2xsQs8WMZGFsMG4EzCNl7uwcuz0wntoERVGiJK5F/RvmESG
9SZhwrWd14/EPudokFBjVQqBdKhPPKYq0v56A54L7RY3VfJUFSxdkkm14pNIjCedbfUAY88aA5wN
WlTgskUI0vPVViX4BiVY7uGilsFBcwBP1/iD3YZ3FjnuB0NRjvFMYobG4OS3wdvUdseDl7Q1f0Gl
Py5v/vn4dXi1W2bHWHvV/0ZWytY0Cl5Kcncaln4E+pUxP1e1zA4rNEukdksc+xSKS9djeFle/YQo
WA/AMOVtcfqIZT+qBQGPoaljI0k4PrHi83pJoG/d8PwasvRKNlPBcRLNUPLEkdtWpHvQPbiycMXH
BvbJDd98YexuVUZicPkEB+AmqTgxXK8ep1D1FX7pp9HAKv+YpNsnSe6DhVv9gxsgFPKdpaHLUVWJ
ZXktp6GG1xxrMaJX+o8LN0QS+m8GfeYrCHX62RuFvxynJyYtZbkkSWiY02TMVyfi6jHcd2HQ54eu
c+VRrZkqCTA1THJEpATg8bs8eBCRn/gwF7NKuXWZE3uoBMytRPbdfjG6y3yG3j+omSHTBRzCw8VX
PuwlfKOrT1x5cl1M7hIvB/qAQLI8rhRuox89s7lcDuYFu6EPIKETb55OdJOAVSL18LHfhTqMkBcI
WOxgtz1l/vt7xkMO93wb5Ia72hEosw07ccmgqqqByD65FReKLSuUZB3x91uYEYPpOm7Jz5PDSgU1
V6ODoDOzAYWyLbuZiCspXIqGKOVSKo22UCLojSnKUFiZY2qSq0C+bQDRCvu5xoOvT9knpaMxWSMq
bjdXT0EwRrGikP5Sn0u2jut5jMkH9cYP/wMF4jt2PLwV1Ey/c/btBkbnTNuITXw4fRF/eWFkpsOY
+6q2gNzftLYP0hrCLcv6YE5M1B/bebka/MfGh9ifE4lFLxNCOJgO6W0BAF2IDShPJMvfdRCwR6TW
WHDeEvFNyMdsWl4TdSMMvUGluv8KZBX9ukiGzCYMjbEYwozJWxN2YqC989z/+f4wpHBR3/4Xj3Mh
r1n6XOlgerFOfnnBFzgw3C/n6/z+kC9m9trB0ETlcNP50nXdSNFIHlAq9Yd49CsmsIqVCqSqPfnT
g4YHwsHZRuWApKtGRTD/3wENUh1/xbpCqjbaIk1PrO83sCEQm4iwWNgkHJmOt5XoAUmPYNGnqXG6
BH8wMj0U1tdxsi9HnmKRYfap7NEISdDA5XD48jHJ5XQldF8xYU0Hng+SVwD1pTRoVVRKuJJYMVDU
1yCesHxJKN9Bfs8m/DJjS4gP3LEclyKRKBGyZR67iJwXE8X3umQpFWjg8xGHogVkwJ8oNALkUqLE
X+7YWFwU2hmRUUE72a33EiCVlMw4GaTNv/jU5QAPzNmdOu2OZdjhoQnw/ccVceM07c1e4z9jd1ZT
GJqNxiU3+jgVTG1NzNGvcHzNZ9nMMGRE+YKCxFif2k4mRmguk4OLYpHFS4nEEoIFBLJJ7ksnokFO
saBHza90fot+EkDTGSn52SHpXpbCUEc40OYXOamWVBW20FLImD+9I+SsDq9DqJAMmVRfHAk4jUAA
Lc01iL+2hwusMWzDLgOgKHL1vS7FhSDTCBFdVPxTY4h2zZG3lPAlPG78DleBAmIGSyqzcBIaMuPG
zop10GeFfIcilHBVmv59s+8O3wMr4DAbwY4n5NKjoG5QeJlC6FXmBnRcywMSk42QQCm3be/l9Q1o
tVZCxnIUNC6OVfeXSDoEoQj6IupT84d/lVMnRcAfvCoRiVtDi6gwvxjmDsbMzARw5wPbexUlQtHE
zcf0evrv/ueboFdlAiz9nKN87/kClz6bVqeQ1O1C9gPyEhsctaSt6MiaXRisRG+dNBrpiFaJx5kn
R6Fh4ot725NraVNkN3Rue3XjE+kG0olQ367YqdXCmzrLjVwQSJkOKm805UypHSBOcn9NbnL+g5xK
DMTGlifnI5WcfaoJuPyA6HbMX+yIZnnw+Uhm3yMaDBphSfZ1ehdLguNHxdDG+3C2kbjzi1ApP+bb
XmFQgFODHATVz/3idH0oEOoQbjNv+O1xF+vl/yzwbfC3j6cukiFK5L4b4Gp/fFttOL+Ao5HJPRt+
4LKmAkN7D8RVIJ/uVYRmau8VGrDBf0EfGwBFekobpkHiLLltFK1JX9CONVmsXmloG54KnvfQ+jU/
Q1ekMrHfU5PSLenvV4h9jn7tzuzyyirnhFI8bBMOlghORhC7Cs19wbu4z3i5w5ezD4LHeth38FYc
4USbDgaKnMKZaTXbNMdBNGZSDmktqLDKb1ew0WR1bs3DvDO1YZoEUJA3T1ffMt1xyo/zyJA5Navg
osSHfSfIZ7WgVB2nennPZVMqbV7KnM+HJWrwjE7B6OvRiTjF1E5HR4URvvYah7b0mgd1NIQD/+eU
bjWbcUYSgmWIyvR73HJgZ5UL9l1AO1+D9SemCFqoL6GWG8ciQs9AekhUD9ABK3xptCoe3gmfm2yU
ohBL9Hrb6Fo+A5FL2SMYMxv9O+0zXJQn7uedDBXa1AKQeLVfTx0pPuCWYwiXgUia1SoUWMpE7Jnt
Z3fFwR2Ay6/PHsIjzq5hHTTsSEwHcXtNG6JON/i2DSLysYZHeNoswCp0ZafoapSUWG0HzAGAd6c9
XX6+YZqW0xp9w1TLF6jKUnUXy8utIrf7/zVJXbcdcJNXVYMiedakrIiA1G/Hh+5CgadvN7yDC26w
ElPqqJwoF6sxpurAPcu7pIxb6jPMHgpDUbwFP5+TAtM9kcFZBoobTzxHpLBxEYQkZLR0rtSTIe9W
rUuTA79Gmo1kQnpYlLq3VGQpgeYn9e/lSirLky95rh2Sfo88wqlUXRBkklFUSa7tdWsgDz3dW3Qb
COQURUQ+HtMi+eZdJhdKz7risa/he3fgQD9crea+6twwX0B4N+qdGnXvseI2F2N+5XDvBnN0TPUE
BTNUjcSCEbiiDE8oc+pcmug+I1i5kjSBafiqU9/1ddrZfbhG3IphxlJ44atLIPPJNqu93CrBPRop
pQcoP6iFh8mIRIKwVPYrLg/xtfmzeu5yFbXGZ4dIg5PVvsXjfYU7zl7Q1NHScxxt/zPb84VFHMHr
osYryZ2pVewYuDJXjqimXSKWbI0BwSDKYMv6G/xootXM8IY8hWYPIV8bmsXkx6GHoWUQg/QayxG+
K2krtt/88IFVV3MbmaPuiYvBI5SgiNs7mZb9d4xYZCoBROHcVQIlhE5nic9jvEbmk6t34KnAWX/n
tE/Aqyi3G0oj7cyaiYkiOIuTpTCNlgwqKb2yWIDUVHQYj0fbdoa/1hRQlFHOjdcxf9goY6D2+j7c
WQEe1NhfuCPNYu3wxQ1eb3Osuh/HpZoixilDVg2684RDdrhKmvCmEqTxrP2sCXZnyYMDBlYgBvd3
vMM1hVRORXQdBOw2+NxllyMwl/tLRXQU64kF1T/BzNzrGnMTDipbsFRwlvyNqjnNz8aZjhmWJpXq
xdrncVR3XbnobwAIeFh2BLs4pL5ViH3hRKKgruEjyaIJZdRvP8DBgRldT640AJI0R8xWNnFjqbjU
klTMbp9NIzO2qQv/p63Tkvdivr2pvddb6ZoXbyFqiTfqp/AVCoA/r1Qg9S/GamPjoOHyUrSH2b3z
lBTkeI+H2K6SFcigJbpjfOopFUZuM4wHhS2ZuyZTZ9y5i21ltNJACLl3nTk4ZXRbQibZAqbGEPUk
Q6Jsj40rqTW/HAlRpXRjm99WtYyMi8wONeYXks1iSPx8Pa5DA9SjSq4vS6eE5YfYsLAWP76Y+331
Ynu5ngP53gD3S3Bz/VXy+8RMBQxakoGPBljE+EP7GJvLR2tamUDlyx/+VXW2QRuIMHI48yW7ZSGC
U6cz3Ai5PhYveO368+M0iVcw6O6oInsUp069qOZb8MKh7JcT/5P58eBHeWIqbRJNE53AOeKgPtr9
/6vLXB8FZM3kWKFabvjzy/tvEDKaNB+S/fpP6kr9pcxMlSIxpww4UuiBqGetGNMwsz+UW6Ingi+8
wR4El3CSdAcvK/ADRybwUg7gSOf0L2mfdoWYGce4c8S9Ctr+dLNtuEEZ1e+h/vZeH0R8XgqVVA82
JV2ZzUKf7aZB8DSpuoXOqW4GskxSPIYI8rpfugHSsDhhnIc9Tx+VCEoIIKpM+ncDniRbRrQxQ55A
je15MvPFFjtJAp28eYi1GceY7gJX3JDIZmnz4G1Ww9/VR/Vs58/WkS/yiYg6GeX5XRDsc+t6oPgp
wpeHwQBTog4BC7GwTMSEuTAaVXuWb6VFAWVwnrk/A+ciRuR3BxlURbR1uo18xVp2JKqY7EsulsLg
+1A8GkLCp+AMqtgaVaCMBAB1CuOwyCtMKm949siIuHXgycPojBuYJ0HGAie6ekCfhm0nejzh1HEV
vzVB4YfqCdjTEgyemFmoIUOyYL+kcGuDQKKD6AzvQSv64JcKD7ehoig7iwBveXiGcj9WsHq57rr/
/2DhmeCu1FDo9dYojcbzG8Zd8Nei4mhjpMo2RO0lDPaZ5vOPPOEU/ZAP40+akAeLaapGI2cXeg1X
Mmu3sJEh8M3qks4rBA7TGH9Hn9vTfhEPLWjnXS4xGvY3xFjWn2Ax+kk/lvJZVomWQHcbrwcXOYRX
KpWJ8PRDrO94VkJ40Fn1egKntxZabvkqXhZuAJXF7NiQuOhvs9Bs+xIcbQtGVa63AV6hXiZW9nX/
wn11IUC9G6j8RWx6wv1XjuxSnnLLCcHZ1nvaKUEVdSqtxZRwGafNMVqEb6r/oucsQZss5zbJtxL6
qRtbZ2lLQBX1qZsNS9BmavBQPnZ/uzoLmFhJ6xOi1dVG7CG7vWo1scWpgFuD5Pz3W9Cgc4W2evKc
LLkGJxM2uZWNUtFgyVUyKEJZxp06cCaefARsL7oyJb3DINYkis9NVwGtjetHVwezFeMHwipL17rT
vIu+VlZNgfbP6y1/IxJ1QMSM0xtyodUOFHcXlYq7wf/wjZ8h8dgBrLszsKoy9ZVka3IEJy4m8W86
B8mt4u99exaa9oRi5zNBU6Fcvi9bHBwK0W6ByL8bRlKJl5c1ZArQb/MSdTX6JQPnJCcH1I7uifmI
RXH/D3XCLf/w1VWgoN+ujYL2Qjin7yInobkGLbFsxYQxxLrDIMzooMpyPuD4B8ooq42n/YWZPJmB
erUKwBS8ArdGoT45AP8su/ufbTupyacaSzsbmLPZoZce/7KVM7FJVmCZSIrU6zKaNxHKb1DJR5nI
hH2JiMpWQOs7DahBIPrplkddeGLsluOlwjPMmw1mNG98FaNStpENF/J2CuFkCa5lQNDn661AUnDL
604B42UnZ2QNeIIMoJ2pQT4vGWzy3lY6wJnQDrwFtsVBdz7Ve+/4BTjPrmpNab3dcbVDlGhD2vsd
Bvll6s122Ek4QUvaHHAwdIRTj/V4eH/JPLezNKY9XuckrcAN1B+6s+aOJTU/YA4iJqp0ljIyKFxn
sB0RC6ERJ2GJIN0qumt03p3DNIYHS+/t3age4ROqmeUTeeYUqVBEuG8+oCjqoBKxYj1a+StjjmCA
ItnIILT+VDAJvGUAW2nIO9x8yYmMiCmgF4ypgUdSGSfipBEH6KVG6CH3fDOgo2ZIYu/wuPEvkqRA
QD5C8msiFEiWiZTkS3SlY+fzn5LIOJ/0BbSdhILzD27yyndsIkOdHmXIJkPSlLVvlVZFKSbO6AUf
EA3JBN8QUVk+VrWuEeHLsZOOTWjnePHGw6PNsTD/+XwLH859uEmqfJZ0FVGNCzc11zhUNToe6Fcg
jAbltqJ4bidBF2UG1ArOlAdcHUKH0cbKQ2oKXKkkLsqVlaQCwUK7sFull4O0ZEfzI7fZ3CFmqa5q
fJ6I9MC/b6MEmNRP8Qi9efxICdI+zF2ZcHsigiFuKwcumqG9u/xYVfMXcoXolQVPH++oXBEIqM7m
qX2L8GnYJ+T7p/ssb/l2t8JjkQTwZD/PfkxmHo1/oxgcM6hsAHSFJqK0NYxjKIcrCucsT1NqTvc9
WzLwH7hvfKQ5sF6ZmHfKKK3MLMeFNpFyl+Woy5UXaiin/h7n13nDLsGmO5yh2dh7CTfAbL1ZcsgN
0gPXumVd1ru/BFVxDnoXNwZeuJnxuANod82LkzX2pXVtAJeKk2Ympnp0J9QAaAasidJ2dWmVlH/w
Ykaj2S00AVazLoZIdkziUNi9uWBCzU59oSW9sFKPivLuPIwmEJoh5DfkGLnxC5Rd5J/Z9qwf2GXb
EaG2boS7um366iLzb1Z/jljmWI8EjrdwLfHBfq6RHB5PMw6N3DirBV+MSGhPDaxeyJd8SYE2+Sl/
hFgW1MR+mdfDzeBVvQ5EuGrBvWKMyX8k+JVrUDFee5L2kQWTO04s2V3+BrKlBbciF2s+FOwoydlO
1UTptLyYoiQ3vtixPLopNBK9nVVezxqgxvCwra4KmuEbOuVA3edsj9OxyBJ2tkBwVbOdgtbY5yG7
cKt4Mp1r/fohdGX+jV0n0TJULz9eXlrorxSnVpa/euFEt3z9jobxyVRIeOgUBOBHtG5TKfFx8vlj
h+aMeDZPVBEpK0KOpfgwRL3qMrSA6ombXygJ8W6DxR7gT9z8tXX0MPsuU7NxB3pkxf2Vy1QuofGr
EJBYzk0J0RXnjkuaOxWSVtqnrD7HedLLoz4pmTuU2cYlzgX7VgbPjUmHEyJx+RS4mOvxcp02rS8E
oeKa99rUfykLuoeRg0liYh7rD5nNueowvA6fp5vLcndP5aJ3PGcS/6YT28vhDbhtXXkKh1hK+r1w
wNtkmrkCWzwTBRbr+WYrM7wSzaLPjdOIVz/AFKxG5NJuZ5w8LC5i0ntBszj/WEcA5Qr73B4Us6sC
NeYLZGryTgte+Mtg3sJGf7ZFD9gL1/AZZ6nGgIwehE+rT1esyvD6cKrP7iBZGuaVCsxFaSCov4uj
JhNbn5kWCMDHikxS0hw5JNLBe/95Nw4JZrLyJWt8ueipOrokzO2cS0Ej6DWBamyzq2lrVh0AQ8+J
JL8I39DoCoaDf1UBU0mgpRcE8UQIe8HPUe3dh8I4WDIh4GA0kpk/1yZHMeAa3QOxPBBevvcr9639
lHnTAA3DU7kx0FPcDwRW3uVIxVlNKxcenQnKo94ixeUvsg84DYYvqxFgBhxqP95jXxJ1dooEYYSK
f7mEBx8qG+Ic5pk2s8bcaDdDN9dihet5oggYlprgU0Pi0UElZZ6tBqYNB20knQtD6bAKxO0QHF8B
c9fxjEuqnayCLgDcVCHS4JZ9kxIncFCX5euTfrJzLtmDGKCK7DbdbMtCNQTwCBLY8sIdC7KLgVWr
/IqGfkBjTTWbc0hBQfgy086tywvXr/D5/QUL6LdwWcGy3JCSihU93hykDKb1OwpvlJ0e93JSlflM
yeglWZkislPEZPSgnGIjvdz086yphXIxVepZeoX072lT+3IfQJg4QVk+SkGqMVS6Tvp9uh2LRaMk
A/9HSQJNWkvEoS4qtyLEPQ5nNBvHKAXz33ssTh1xNkKoBkgKx/Uo8i/7N8o4XlhnJbTeK0rWJE4u
MqfF4Vc9bSAwulH9ZRbltkViBH3QnPue0XljYFYn3iQCpW+0EgW+W/aGTwblWJXLn7xlopM8+pkC
32amolAZLJ+ByEQQ+OLXfhsLYfOxPTzdrbXaQDXPIyyaoQHk/6x4AHwrvciT5aXymRO3g6NJJIyC
56eVrXREpQB+Mxt81sokNog2X6FjQijK4WGl/WoAIM5Rq5aM+F1YBKSUtx82dN80Zkf5QlSAfgEx
X9mE5bZzT86I4j66Pj1+V59Q8yOws85QJixl7YkEitED6VWn+uK2L1qbp/XysApzPhA6to8babyt
1rCXiKVAjbMKqGWRfQYwB0dZgLZYpkG0qX9HMlXwqlU0EXHhsj9/JZCRzn0UxxCmsc16VqObbOyi
LyXhtSlZD79FvtKPo31n7g+WIJAC9NYraKddRUttZVKuz5oXYkoXY89fQzMQOQrxL2UPecGAQuy9
q6O9IM7t1D3k5pJUysp76rdObPrXmFjlnyilsvI0LCzdWxEM7G8kSnKV12xuDb4hGX4zDPguZzqg
HrXj7scPOZPN5nQmG3BEpUfZEzJt6oC7CI9T9LRZevcqtyUCAw8O2Eoqo71Wfiz5vda6yjWYe0xv
BzwOQVm/1dOMun6c2+svNm03bYQNa7jxjG64aAtow6j6U9ujXIfw07IrNfdCNjogT1VFqpEOC18b
e51LHGPSDG3Wxw+GhJkmos8M87QrOGM4ygawu8oVlMHu+0Q4AQvcmynO7zOnXigaA37KqY/vHYWJ
uS40yNYu+SeZ4QVW/xKU6iN+PtmBigiDQCKBBjWqjWgA9ouQhm+IAexBiF1+nGMtyrf3Uf1mXJtx
zn9T9rDxp2kX8rNbkx0hfUN5S9t9DZSbTS/2KeZA3cybcgMcI4BtWobQn5yb4M0To83DZ0lRy10D
wdJiEIbeCgxDZmyXeUHUNBlmf6tu1AykOJasZvs2YLpVWydMMHRO5mWmvC9qM/R3N1piIt3NPj2C
WbD/f0j2ptV2N4/saxD39NoETu4h83CToBNb+nXSfMMryL88nsVnibP3kEomeTBbv7hY0Ne6EB73
NsT6qHLyUBoMVPNoWdw9bnnYYfxvac/M+Fa2V0Nm/eKSrRY9uFUezuuCeGnsBv/sADc+q8/n51EK
EBTYRh24qy9fSvd99hfbBn9VxVXBKiP+Igon3mPBzQ9JI5aiJEccoi089QNXHpn7C02uWwLOD8kS
vhPSZhGPt3KQ5iApqjKUe9SV/JNRH5XCCdPTxG0xyItGxWjh6bd2HzRWHs5ito0iqi7HAQBWZkwf
Bw4IJFJO9Dr/VjTXk5oD9yu4cA3M0UXDmJQp0EYDYzpLoSMhiP8BZvHq33OfD/bpF5h4mtjt8TxA
FBWsIBLwN8tYPlm5uXgBAHZPBv+f/dNWxx56eCjlc7OoPLk6pVouliE/YK4Pr+opBdcIa3NbI2ie
s+Xb1gk2xa2V234sp7d8jpmKj+af6cJLzQOqM5GuNus6+jnnD8YnkBm3gAf8n8yWOj6nu8rc/RDB
5B9YkRO4MCcF+gmt/0T+or8HwCqhTismt5+UsLxrTBFZ72VRGhu4jbxuWlEeNaNF5AI8Ga7vkBpR
euMYD7HpRbnwQWAtecVQrOJcy+WdmaVMFy4t6RXr6mZsiTYxtMNsdbVCaroZqXiu0CR0Wwj3wLsL
5GN61swCADr1dZr+TgsG46lvQ/7kc5inNNPFQ30kueaIdTmk+eqeDN0s2/E0ovMvx2AY8MClKI9+
6N1bgVl7G0A2o4LZGYF6TuNzCzfBLeUNRchXBFuKPyWS3YnhvEPGjdsdruHM3s2qxzXOG2yLT4Sd
OXp0W+DJe1k163MzZ6zXB3Byd3jfJ8zJiduUk+5QlR77URiZrg9N/bIkR3YH/9wPzZtNEXlV+3su
Dw7j5o3DbW8As0Nkv1yzKBagu+yjjHWLGPN57FKaWnIT6iFbhp644ez/ctEnLyJ5hWcRYqZ5t1Kk
qRoqMwTRoI9pGgqIQerSOfJalDtBFWVnlIw0xTPgAWSRmtjQOODF8hGmEfy6WpR4c6KO+XRSqNBw
hzpQN6RvzCz6fApOPCkCAYPUNBAyxw7bIn6gXhbH1dnc99vb4dvybDe7879ReQz7XhWIh4v82Y1e
jk3aoNbmWJhu8jtfdn4FfKThaNNu7zmIrgygZWF+r2iql46yclT2WKhrAclER3oIIxn1E0agBkg1
3+8AkOPfTAWMEw4HcHTol2/AoJG+igWav+AgabjsqfmF1ha2a6CET7hhhTfvwjCk+Olg066O7EPw
5ebuiZ5Pcm3XkWhbcQSEgJkqZiKpavOugvfIt4gfZ//FV81A0y8JtXUI2yGLtYGI+1wCcqqO7ZBb
sNGfpDPaEdN2kjDBsN5j4FjxllVF+zVcylrhd1Liym7RmSDEcJemwruQi+1nI/C/G6Ubj0MiLxd2
HKjmzYS9QenX2u8j++Tj7H4Zu+8Qu+H56SnDVMZa+/Z9fvU8se945z7LxMV5NC+6VqtZYzEiB9uI
yvkCjSACSGEVJcq3qsDGOw17RgvmxGjccOOjR9D2pc7eRNngKmq+lC+XiFgJjmsDlP2zzWA4ZFnC
Hjw8QO9R5ax6bz7GZykcljHKuO8uhAMCygnc2yMG0YMezvOQM5azdNpdoq/Unh3SuQKBMmmsvv+J
3vJi7GUUAXEFjRYca7xPeFA1QNqxQrWUMpGvi8js0Ot37VoZtwToZ39GB1h7GT+K7+wTKblfPML7
zbrXbdHb8PlCa9BFLnRW8JdAnjLNg9+tl62Y0ydazCBvuRPkaRkizDe/YYQe9EMwLfOnRh6GRELX
kCnLEb5orQ1QosdgA33D3L0Kec1CRB0bsnyT/CE9WyxPVwhKtCzWTHB3jitn5PTgkPX7lVRiF5f/
nD/nsKX2vRT4aytW6T/4vs+pfbgRlZEbFy86/emC96wLngHf+0CCGkbPs2NxNk4h3ZnXuFBvWPJj
7vkPa8UyZ8DsUlwnCvgJL/09eb4j7z65Ksko1TMAskgkbaW09R4rl/NLzfHn7LRIaq++CJksiPFh
mhS0ietyQFLN3eBAMFEmGd/p6DhIt1Hlb+74iufnYYXqtsuYe9W/nOJcQ4OxDj/nZacgivm82uWW
xDuhV22CD1x6esB9RGPbt022naUB5ut718dbkHFnvi2r1B0gKTro4CESyZL7UNF1YllVfuJ28frs
aWvLZeFIkwTRHYh/Nv3xLwAUYm4KbmtSe7NR3HRrUVtBHa0TNXyNpQ7Gybf3ODFcO2asQIHanobA
PAxJ2dLfxaQx9Qhi+qoCyWf2QdofHl9bPGwBkm2BOBIVtUXnCvLl/7LplQwL3vOqAqs8pGD624oo
s6URnjRxzW2PnhIYXO1dESwHU42aBWH9cnG56jJ203ng7ahL2r5IVlKOCFWp9Sb3bMQxqVvqe8Gm
CFGNmdx5VV3WrsNrJYbHNZVDqheWp3ybgCRGoYPjwTUO0bLVegVXcxRloRvN3ZL/rnkZQBsTQq8x
j+cpWbOk1v/+1MMoSuE3T3AGPTGP8MO2vJQG1CujZwF3EDN5wdVuEjWbUwQK7Xb6lGcHn1UgX0KS
pyFFoUYzjrDNLHl4ndZkWaEHjRAT8O+cDP9pqlqXtQDyaPSRULLOTuU2kQe753+TM5aB6poFNg0v
YbkloqeTV2Fgi9cOxEq+8W+cj1H5dijbCKTMdQ33kJKN+ksIuaTmZWJ3GymBhPaHjeFtfaRSokwg
E1c0bCLne7qWvd6bCgBa9Zm3jFUYhheOdRqaNzu6eR3psoJQ8OplXyZzOpYM78bVcUYGx4t/V0cG
FaGYFyMbWcmk3vXEbR+/aUDb0ZzS4v5Pb1pIcNCncrZiDytqxiaILu4DxnU+ZB6uUQE2LEQ7Nh4T
in8g1i2dv6ZN1wLGKCGLQd9n26owEagiYhtf64Xh7JVtzZeOrt5A4H7kazC4BIMoMGA7VTPTtMqH
g3UE8QZDy0LsUmnSK5AH9sJFvvjHoBxupy0Kq+cVIaDnw0A9VXxmWzVs+C4WgXJcCvRNqF9f2HSf
MPTlZW1AQPsyWYf9WBbFxUidPv04TKGPZIDh4t2tJmY5s8roaqRdEL2+lx9XZ5DxMBjKPprz6TBM
zgVeePoRUPJ9SHiOOWGdH194U3SbA3/dO4mHQ7Y1BK+VoPjdhjcWRSD5KHaUrWi2DxzVF/DcneJy
/203sfQFzSYtMkOHTLsyrolCB40af2HnirJ4c7gwdKPUII4EyZ6Jwbz2IOSlbK2koKPnUayddyrX
lzclKt/keLmaH+OWbP7Zpt1lsTy1YESRik0EwlrBWJMwZauNk4U8+4x2EbZscxHcmKXS5UxGOUZS
b7j8ZGrb5XLQIHp6PoElgMby0g2u16wDZXtkQSmECqytqkJMheRbS4OGWLpgjZBufrC5so+z+ekD
naBLNO1m16eIXFFuJ1B/0m4HACnTrw1KuZB7YqjdYyb1ymNPIt8IiXoy48HGmqi2ZuHPOWFK5P+R
lxvpqTjPZFxVwkqEJhxLd5fUX07DRt8/nYR8DO5Eh1wMIPhqDSZ2hHZ+eRh268wWfWszTsun5iYv
5KeV9sbtGYH6q5pIsq+HLh1+f2Cv3Ucv21NrSHO5YjIpMActeFMarHS+p/oI19SYCy1FTf4v6z4r
1gk13zNWT1bLXj2rNpsDmTZjpwzcEbd1GBrZlYhoHwE/KI3258qJlDD2C/MI9ox2zQETx+dSpF1C
fG6PZbwaksiVkYUGNAGFGTZGqxDad4HTkA+IOOzfQhMtK4v+yMYKU74St3xm79rw3jgsGWQfP+g8
lOlxrL5ZCOBW3g/VRVmJjGfy89pHSBjrcsSPR4tPwzxpAd44fPyHWioR0K8OIleaZzlGGo3VdM0q
udaeQiWww+nxGOz7dwfDusrojgCgmSr6aqgBnXZa2VSrprHooJ9o9AKbqUV0HHxbd/HGBMvl+2nn
Qa5NgzaohB+yaIsVWU3ekLdWM5kwBS7ytWTSM8+buM2cHp7BhQd0iKTTBHSNH0RVkmiZTx2RzV3K
Y2ezrjkhzIiZoDvD1xf8Kv8MqjVu2cp5t4/kWsMOYmBOiAltfjoRaFDJha9mJLQzq0kJKkQZ/4Re
LYke0SJk48i2YFdYklLC9Y8QP5U3YCEsyxDSe0eDXpZUvzx216MGi7AQo0mP3Ug8+9U8iMcH2t9K
wfGf2ex87iAGtKC7CHtkYsseSuSPe7/j/+UQMAuBXCMXlCTR5zVbT1td+cVJXyJCajFEBztwE/k8
CvAot+bjeWiapmfksQfMf89OslHEMA8xL2/Drb2P/n/q4RqnGJ60VJqS5GiPHSN50Fy2tf01bqC4
kKQ5aCoZPbVLs72+0fPi9upg1fIlcVyIHHzabuTuAj+5zfDteARSHqP3QUk9X7gOvMohXhJvicx3
/hwayAEpl7G9W6RNzLOPEoiyE7kQ9jXxjHtA7LfkkaPlTbh7D9viMox0eJUZxrlZfM55k+dRJ18J
45IUl+oBUhNwIo/7r8WuzbqRXRL/ByWR0ztidTyNDhlvGU9rLESUKHlCQYrlx+kXCtMMSK9Mkcah
SSH/x/XUr5BuZ2z13TvaPjmo8gcLdsCV2g7mrL24y2hESDqyzW6fYoTRC8oF1xGBZJcFuQwanHmP
0cYXmv9Z5J23as1Auw/ztMgZgTT4dh+GUyx7XP7YKc/DXrFuhiJNQaYMzjR0U+j8lLPLmF/Oex2m
sX6FetwwiIU/uKJv6a//W5kSSB17XwCw8reS6Z9r7r18a+gYEeZZvihcAUKgv9tB1VhzvRXQkRpg
Zt2cTVgfx0uM8ULwENeJI+0dCXGjOlyXZq1YkPBqLwV4MR1zmzh0a3Yn+RjJv0IBbOTRL9TL53IZ
h7F0G9HuEWb6faRlPtxeftortKltSbg4aQuw5vFofc8TUiu/no25IQl58pqLAixfqISDoeaujP2J
rzFUy4ARvf77AIwSZgTIR46BaBKc7GUKTrsXRKNPRO6u1S5QBVIrcxrOQ5DsYZ2AvMwP2M4r6jxQ
Mw3pdGapGmpZdRAZcXGV77/SLOs1VSxlr6NvoyQAvxR2+IORLuruUJIvjkAA2mp/uZxE/lUXsNby
7mMWQAh6c405Tb9Hn3shIjJq+xZAcT5GWPJJh9vFiqTrpjSKOi8lGt7YXrEbozLEkQ+wXgIU7qr6
NR9Tx1TdWwwVS7/XwPjQwEEknP5zJoE5oVGUFY2Vi7/3Rxzbli35LkWIEzH8+MO9JFR0hUjuOc5H
fmj2afZxnacjTNUnZklojVwQS5usogSz1/WSbDkH5WhaLASZIgNUItjnBWiN39CpaWz3BfU/dj5R
HfGjP6MnHV+iCVgnRo8KkGFUcJmeYe77s7bYalwYHXs8ZGsA4y0pC8lx2i2mO16FOd+z2sk1qwCv
tnGnzO0HZVeZJtAdgS2Ycar9Dv/E9Xggt4SJnQ5MvARdmEyZbk9ABWvvVHg+G3LRU7mpoqhD7ABN
Vw1Z8H07Spua9uRLRFA5/0uuDT8qY6nZYDJn72PF2hu3734T/NL1d2xPnn4jNnigkhS4NGFHLwb/
2Ov485qz14PDl8Gru8eXkE5TS8yEY+UHU0mu1YJl/+jriDrfFwVXe/H2Irzmu57EqRfSkR58U1Hr
0ReFWnTFtvB+rYgwxogMy46K6g7VPZdajbeAW1KVxV7QB3izVf/c/enPytiX7qwKyGB6H0iQEWrI
SZGr/aF/WA1EFKrYTrWrz2GlMe0JMQxBBHY3zsMdRGno8pVP6uQfVZvDQnJ38EuuOK7Jt7z9ojVa
B5U4+Ngu6EfRTrZvPLZJiGzi60Fo3uOj9x/f+tCV8owpaJWeV0G+IhoSdaBkqMUm3Nsjv3xp4e1o
Kcqbvsk9e3DdLCHQF2rS94AKYfushmqHtlmmO0rSx0NwbuIDAYtYYHqAv2AQQYt9Q2hQrIXGbgSe
n3pLmb36arPxYE22j3mvmYg1WuhEVal4EtlPrZ3arCTDn/gPJyOSmmBczXkjPV79tpsbOr7XdfGS
UIXPa74BoFq7xozFUGDviEUuDjQ7r4Pp2MGlMn7gQsBg0Uf5fdab7XblNXO8OPNBAcoIxN34D4rp
TOkr7n7AKszAAT45wv6vUZfnruhJCo7AQ1n7PwLgSpJmdw8Ko7AI821UNO1OvRgKwf185RiY2MyG
KtEJbE1aAlEiyDGmcZT7vl5HPQtN3NpnHrdWCGsX1gr9wwNgCf9K46jso9glUly/e54kW3g4B4nW
Bkd86wz+wTRF0/90A/u6C3vhwQLnMaEoakaoNG9J4ssXB4RGri7reF0VA9OYH/BUJGxAvFSl/+Zx
FNOysFfrCFu2hwklTL4YCueAAmFIZcdAPG2FkChQ0zkRqyYImXPph9cLo5gn645NS8DuxWbtIEwd
X+0k6jyTncUZ/9zbLL6TcFe/nf/0bDZCUuiHIBQQykDktlNic3QltZdlldZm3sRlEOX12qK+0WOD
oIjxIdV+DkvPMl15czUlvevPIhtwi+Wt5nLjGgBlQ4qgcJcGwC/pZnWNl5cT6nxsY3ut3d+oPQQi
EpNH+fE/nrl/Gt7InFZ+pW3J8RV8p5WrPoCwFfZk1fCJwfWTLk5TeoSR1kXw9sGiJAgPPD5rX0Ou
0zwgA/ZKzrms9He7SCJSUOjxFYCAk3RepudaYyq6t0DVRe48VxVbSIlAwjs2Jdp7eQUclL2L0Q7m
HF6ISI9YeQ0Ivl37X+oTRErSfNAOmHqqAppC19EQA9W16FSyd5mxSdooBsoPqt0UjmwicZ5m7QZJ
mji9fvlMwFq7P5MEcoZjL7dXHVa3QCRYQNJXkacTONBnL8sMDRFa304PluEJoib7SB4Ka8jA/8FR
F7s2SXBkJbAHKyyGMijXwjIlPdMeMPmPkpgz/UwM8mkGubSl9nirlTHo8OY17AHzCMFHtsdpV0x6
N28eDNAniAdpfYMbrIJt0ADnO9OJ8EQzdYx065Lq5QU/fgx/frx8Gi/wUAk0ssvLeUH7MwUGkLNB
n5VGMSxIAMpX4V8/IqlV4OF7RhinON5NyCSLxxvIz5AHWExEQ/v8++QfxFDBmimIMEHvLLaJHqJv
gdbCRNQ3/zCELFPReXyezw8ywFMAGlgfDTV/90xhxErcYBXm+bd1shOpK+rGbBAF7iSAR16LbxeK
hvSvN69WI6YXehrkifXAqBHq0WC7g3g+QFYWPbv73FcHU/AfNejMenjqGf8Uwh1rVnKPlD6r9Xkc
gN8zarJw3OTWVaezx+dal2SGAFC5fqMJtQQNTswSdYLTwkV/D7nztUKj5B0oBWI3yj9ip8UshcNZ
MhiM//9fa57g/OEsMqiFrKfeLjjsFn3G4hre0Jo/vHIu8JfZ7KPfuo4ysD1XcFWtKzKzaX78J6ru
DhvnTpiM5GNNhPXOX4EaEvgnaiyanKwpznwQ+hfbXNM2vjPgak7KxhXi647cRxl50Ik+hj/pIsHe
kl9AfkDK3A5EPJBjQAEqHaH5tkLKTD9UAnX3Ycg8JvigM5trDQO1AbQmv9fOwe0aDADBQZoPCuT4
J021N8x0jEnApdIVG4OTLvBJqcfeU3KgFHCpp3suTerQUVbYdcqyfyL572h5GEwQmxCSG1bEKivu
hYV8quv8/8k33ikSKQltwdknAB52r/BoaSOXN1847QJXLeC4+TzwmxxO9Ck7GmFKZsa9RQHFekc6
sLerZJmRCodAojgzj9Qjc3xO09+UlTB/GMBqPgDbOcUfRRld5Z+M03Wx+PwbZSeuOFVpJ8CVgeVN
pmD6KlvfWt2sMrNH/mg+QsoDTgRUsnYRFGQrK5fUcr40tf5nAiJR+n4zSYrgQRg4KWe8nsYyOv5X
ljpRMTQjVP2Chn/kG9/UKdxg9FxkHhoV5SvQNpYdOJm7RekVEgIYQ9K6GKVBK4GiDao8k8rOc9FP
9DORlnIJ0k0rFMdl0LWyFkvEql+Flbb9oHWUNzi2hBICdemYGVmbIShj6cT+IrNPDcRl3qWwiQTn
VSe07TnVXCG9zcixxdSWfXAIYmlvijeM46j2SrEqg8MQqPtMZwS/T2GTZranIg1HH/I2s0AiQc7j
Vdw2VTvB6hi7VV5hgJI/x3eEtzFGCYFHQiFN9fBXwoab4AIp/QW40UvIza7rEPMnQgUtWtoTKX+i
czc4S41Pu/WL2rzbJx/PTTzZTxo0DQ297zdiTJMnZ8AgBfoLnrRh7pHKXDMI+91M4sDuEP9FA+EX
ryQX4RFYTwGhHwSzfnlSggTJrNvNsBSgAYPI08c00bfq8zDskNXH7xpkATQLv1s49jF9suH4Yg2g
ENFTJ83H/jeR/P4J+aUDN4ShAkxPa7b0WVYMnDdx3kevpeBR15Ao3o5ep7SX4jQHGBY9reEsFQLb
aoisFIXkdk7JKa4CCF0mVww/6xNhIYqgkrZtQsIzcDyWOhV9qdC9c8vH3FVEjIAA0adtSNa0K2Ac
RW8of/zjMWaIhFZTXbUCQahnvgurU0yvjztxbZsZAc/JA3JCUInb5DHIWAGiVEoEKNuPGSUqPXnT
scCV0otc5h8xfzVFl6FT02LDw5qlwvcOF6eTUsZkVXwMOiQ9N0wjOvmg5rT+VVsRPt3mk0SovoXa
O8LLtniCIizcAoFw6Tn8Gn15QGA8hGXi/A2pFWGJDbvvPyjuYbLHd5mj8PTmV22qsZ9svjcU8otO
CM+bhs5T0PlGeKkKibhseowtuq2DrKlMNb0MPtwa5gQWlpj25jPOyu7dQjez2xlVnvAR/uhkOdR3
U3w7UgisPHV7s/Il1UoafwQ3pMonpkWydpdXdWQIoZblmqcCQFkkS/3i9nN4PsPFyWNHdy+Qsehh
Ru/mSCYLnh4GlJpJqWO4C3/3qjvASd5zSRreol/+So2orAy1niarCMweeVEngAXff7Gs1K5YhIvY
GshPm3ikvnVY4fEI00PlV4iR4bDcsFQKrlcbd/GqyEcMSKZhlgfvzIhwZ5GAzoJ5LWiMmo9zUbM3
CE960uNPe/1XAPW9iKVCXmiTki2JJhdfdBbGVpSUnx7MEsLSfaDB9wSuOxbMhaJTI2hB4b3tmDOZ
aoYC9JLERcsamjZ3hGUXhF+YPqnfMxXBJwYyIKea/bNh43kdeI8+ywdi8pKFwJ4b3J9O5QsyPtWi
JS9BwoPPoI0CJs4jemNFIXdIoFH13v+l5ikUWdmecAMTGkz6QvpwTcJQzyi22xKSQ39tJnusnwzS
qnbSCr2RFLAHjYmOespV23XvQxtuhpUXRB0OIOxPnypXfHY9HsaSsf5JCG8YK8AU+ES15eY487Wl
pxeKFDjfUrSJD0qBpHn/XR8rT+4Zs8BzZjWb35F7fszeY2LYVr9gLvP7ADGWL8qXmZS7QRDAG0ao
YzSDt9pYbQoSqXeVrI/0PHa47SdzSQWYujMZn0kDmr8Oim35EmuVuPG/xjczYUKms1HS7qe+vO+n
rhsrBMCqIU3CYTr3q9nLr0nF3rKn0MKsd6gJu7jpndtUQSEc2Qh3LuaI7YF2TScNNtycnXZehTaa
D2qX6gqa9d2LFQriRBd6mPHwTRJi7IFTw7t0Fm3ThV54yKglX1CKRNMoGN0+WruoxbbhJJvQiJfx
aVCAnwjQVViYpGoT2WOTn05GQ+5UYp7chheXXZZmTt2vcryAklYiz1YYTiq7v0dHPMEtS/SejhPr
cYURfuKRGK4qucPF5nP4YtxoOrRNTDJp8VVM686xWNHlOaCYAuV4x/UfkLwIlJiN6ZXYs1qgIWwe
MQiArrnN6OvCmBtu4ExR9PlIq6L/UKNMXU4dmV5iX15coo+ulRz/a+3KuQyL8hhX3G7yLKElCDz2
Z8NF7bl9C0JwGB9n0LeShQkwjbUFtFQF7iFC7GzZjpCt9Qr99IMEFHqc4bdWy3eRQQuQk+rSOUe1
OV8nC0yFbzb8eqEy4gDJp4uUL+oHP+LjQ8bwsBx5Py/ADTcxXekVKtvLgjTP6tpN/sRgpWGhr1It
ibxwFbtaL3XhN8oWs7ciRNc7wNwyEfb7qWyQz/F9J3zZK06t5tzgPCiPx49kRCOxptcZ+/22ktF3
BEX16xMVCzKfk9m8tppHi1aj3SDCegNnk0Y6itCKLI6X+tWzuD6j+bAnc6AblhGbReyZu5sNEM/G
2MzLSCRh29mjClFC35jHBrdSfaoWAWBYUqgb4fIKkHYEbjMOvM/mi/i+XWEokAHOIugkNg1LkOyu
WxdxqYrsQgYBXgN94wqIfb+eyYrLONVVO/AfF6VLHvnEG1H8TGEiPQVZPtfxIK7+wJNV7vPSCrGy
wjSNFeVl+WK11Nv6RjszkM+fkPL6mnXkp6LteJHjBHPbGES+564DgUmiz1LOF7qbBL+rjsaDmnxV
fO2avgiHeIt4Dyeg0DYp8Mso6qEhsGeDAkdQrW059Bwd3GHsZXxqTqs3xnvH38XWgNFRqGJ30Yu2
veI48+EC2psEUSU8gMcb9V9u7Ul3N1NTT/UWKhJCseuI4Uew/bSY9heW1Gm7EPZ4Y8/LfmJUMBPs
vOn8lIf4arBWWHPoK5Y0iFPUVtyEMGNUmBTP0/AZETtcgsYeNsQ04MevDQmhdqKrn9CZf7gVnWGA
snSmL1ChWickRZTiF+dpzRX5491KJk6d11TdRuu6zdBbuFSHmgiefxpS4CCa0JH6yqCAZZHuzO/L
FmagBwlEPqB1i3Dc9Yod0LyV54y4do6MP3H9vORkf6Q2QspJLKA/Y6COPVEre9D5qbl34+GMTiBg
Nwjhrc87fvgtFJORcFdsNZ6juQYEB1Yk3yxNzHiUu8S+N1XLQuCiVhybFoyatVKZvSMZ6crhBV4s
nsxD3KF22B7O+AztIYs+dDYtdE7I/z721uA7RH/d1o8d1KmJNEhPblUyu2kkBeZWUCC+XNKafvh1
3HQCaUSXtNaDJv3fIGrZBlTea74/YJzwh5u1nJ2FkD77cdfPQs8ZdvXrg/ghGszbpGvHCJK5vzkF
KQgZZx0AI82Ix+Dou74EQpdmnnlH2Gqx0PzAqyuZoyP3FEI0kjizD6m23TOMqWTls2bjKMFmHXRJ
AAydGwhs7TH3HVF0uuE4dLeaon6Bo3Hwz87DYp04bRyNUcrhR6QPqdB+MoVbo0oqtzzTuoWHdJXy
AEaFVRu61JktDqOeCH+XbX1i9IMO+st5TUQMYi7TdAi9fP2ZxGO3fm87N2sisC+7yHW4FHyhJYTP
dzH0H8vOoQY1IyjwPgm8U7T7n+dMiSO99tLG1seOIybra4uT0TOSjmBu5jpfSYr9eTX1UTzoIOFj
E6MNtY5jsLjnF5N32fX3J7ZoM1MsAv3U891dSp0LJ+WXcH5vUE6pH0dJOmdoABTRKAcKclarzui/
z6GZWmAnpQgqZs/+eSQdfRASKhGyc5EigQA3HM1HCLNLmANTkARIsHYiioJN24208kCGqfxpF6CG
Ii/M7vtIFabsjWzZdDFwYdxt50oi47LdJ/TX8CHF7IMgkEsTtaHYEgyqe/QGVHfkPPtfNvtvydWa
phUkI4IIBvnAc8pPUsby70D9PbT/31V7DZqEoL9A62jKRYYWZHqx1dUgs6acG4Ud/DyqO72t06Fz
lqMExin8mNy6X3UTDcR5yrGxej8ao+hca59DJzA1B1YDPgGHur0i/l2vitAcjcvs1/WUMITwDx19
fcivDGPZAPuqOel7L9v7CotN4gcWF89MLHtNwfajaL762oA6+YBUnj8ceZcLC34G5dsslj01AegS
pqs+nTVNW2Ykqq5EiqEsyfxlMTc/UfZ6ybVVjnI49OpZ5ZRU0Y/VgUpwpx5auQCzfBnEhR5I/rGX
PwFrEtcDds+UfpdWnh5/PJtbhYySm3W0/JajDd0rPN0fbHpG2Lu2Hp3qs3PUtZlPQtYvn05iYkQT
X6NPFx3m5wMCVz27+91WAb5e79eHKTgG7erLZ11NCvRuBNOFWKjyYioqYtsgv0fDSV93pd/TKll8
ZgH+yHygssr7hJkF3Q2zR6CxvyKTHcXNg2N7tr2AP1CZHeFLKL8WR2VOLh4MmtR8SdMZKcbqH12V
ygnCCgkty00zgzkqFzbzH1u9G/I3mu7E7/afe1rW2h5BPWDz9xFqx64iqAUqMH3Bbit8yjzJPHVB
26cBDX3dXH6+npNDHOrNvxU5WW9356nmzuOl/RiC9PlLp5cIYLyctxESn65crI4fhBR5Q0MevWG/
xVsMRksb5kSQzezUTtHclSWmDRXCG71zteK+ZbKDkGKnx1+dBmaWuCOuNRKhQFENyzD3NUtnOFkM
iJsXTZDZ7myXmDY0lXqolCMDmPH8dUfhFgn8uLoBcg7NJrgwn5Gz3vHvkiBHU92OzDJr+da0BU79
2zBOCQZF/cm2b1uoaAA7XRv6pk4K4TNK174oJ/tasrKZFh/mDOUNeNWsXZgRfGhq1N5c0WuRYF+K
4iFRT4qirDiJO58ceLs3DWNq05TGkPehdlTiz89owOx+oLrAnq1qs4cBC4enSOqDDmOb/2E1RwBO
hU4kr252BBV8G9qAcTxOH4tv5zx/ZRDS9jKN8IXiMw8bnZVy4NKapMxAMQfxhUsmJE8arOIw2U50
8mCo3GqawTWebJLwRdwFMQUwOeYUnC6lCum5yRhaKPEveCRAMZEh0sAd+7+GlgFDby8bfCb/mEa7
bHflRKMnxIwR0bjj4blXW3MjXyV44ZKsHrcucOpcERS/5kDy3LTMw9rdl4NRQtlBblJ8S38vkzcl
hvVjtBZ/qHal9MPrvCvK1+ObU9Z7dKrmNZez/A1A/2oJQ6fBxkjzGJIMo6e8SKm4BsNCyqym3ehJ
Bzuwxfw+4CEov+PzYLmMd8wS3eORpeXOurqk6E7JFNIcGjv52D6YfSdrOfsdI52siHMmH8XyzGBS
Q9pQAm0d09lGgeSvOCA94LxEbbJzCihl4OFTFIn4z8jTbRd1MtV/sWrIcpJfFyvCIvW7JpJYlLCi
4rqn6PRdFDw3SfCrQAow8m3jN6qCA+AeOiQlubRP2xz1/L2wP+jtciiMF9Kp5W14JXi1Cb+OWydN
P6PhTgBEEJxxLQdn07ArA8xx1ds3+Fy51VjRt5QRRtsK+B2JnW/OAeiuGYsiH7I6CuDncPHQP2Mr
9z06HI42n98QqaGqkKooUxODbaKtuH9K1WLoLzDvNSMk6s55TByHeDx5tSz921GX7BwQy7Fzc2bK
xck/qIfAXrrxpLSWdryrE6z+ABHysWbxw6qoRknYhlLpjXUBPTJnG0kDLFuoD/5fLe9AIbww25e2
70izFNK6F3kHK0v9FpFoc0x9Q0oy9JwCRTMwn0CHzz0ZsGXoWBjEj46k+iQFABQBL+0wSwpo9cHK
tPdUDvw11g5tKzF9jiq/48XlbsCyRT5ctK+gal0432w3zp3SaDIfwS2rHncG6OqoP43IXdgbU7JY
fRbMJOfwe8ogeYY7dkG3qM0Jk+0mxxLcHe4uzSOexTD/u8qjDiMLnqo/1fBj4mvRmuLENk2MlXsP
WmW9Og4Q7U+LaCppg1rAOrg1nCz5mDJt7K0eUly/Oaqs92WPpgTPr/PwENErqN6qMarIlb2C8Bu2
JaSh/ZT25l/V+oX7NEm9F9OCFQgU0HfWQde+kvkm9//9AAp65Hj4Gy4u48yU6w7r46PJkge8C18Z
HeK4AQgsEiXgLIqMYg770o7SN3nnBv7H7LDoLJUOBPec2ItZRnw+N6t7BrW6WjyZIGMum2DV1beP
c9hEPpgMBBbd8DyVrbIyNTShPtDQXCKWkVDZddm0gFytntG8XGreAMb449lBGuSb2CDBJozCnJKT
qe0uAySd8gfQPNbw2GuXzi/aa/vIePMaXbtmDR2joebpfb6kazg8fVLE8Vu2pWTIRAv8Y4lVT+Yg
GgGVUN9UHIUqOktY92M1V4s6QjVd+qQSWykABQ19uPJNjnlPHnyKTNeu32Aix2fPiyI++4MorYsH
gr9Q0nFWE3qu9b13CGS7aiMSA6xTJ+UyM6hHKHdjT6jWuwxBuVvFRemLMbroJE4m618cZbNxjaYN
frwvM8qckBojHqG2ko9GVUfuwbsNw6KJZS23fNxLrIR5T9s0t/zKLoBc4gJjGaOUET4cdkQATZat
jzFrEtdwha5TzHzIElE8VyxyxFita+n4aamZersymOgfRW8TTxfdm1xsDVYnhf1MXFplVKJw6VkZ
2ROT+btPdleSVZ6/QkEyvRKr25sjfzH5KPNAxhIlRm56NTkL5V2TfM1AuxwhypbdL+ulLIRBXcgz
DllMGvzO8THK9NFwJECDdo6hribCaoVDyv8CbzRXZnhx1EgHx4TPQQuSngPgOxZN6P9t9ALAonnM
h3j8tgcSDjppYV146yb2ovEa1zhyNTdLx7aWYp2GKAyzaiLLN0Abs7PNnuglfOExd4RnqfmmqB2r
fdaGvbPKTPFaJMIytUxIa42jtCb43HcjVgHloAtuB25CtzB+v6AWlxayyb0M8HzvOUhyQJuZ2Q12
npYS6/4NLQR1wK3HY0krVXDJEEQjOrB5Rq2pa2B52ezn8zRs8veMpBSZdHFfC4+oPnuvhktVfLJ9
YPC8Uu2uaLh2+5ur8uPl27qsy7MYs44tDh2l3bLCVmdDBAQA30boIuM0a5EaK1yAzcVTr1oQEjWT
QPW4xhPX2YTBlTKa2hRe1zbe1UvFrdDgHsbppymaiWvBYW+RxIEUw7Fm6LW6ICHiHSlBLItJDViI
8WSaMoPFQgqcd851OKBTcy5Oky6G3FBt97Zkq0nJIAOCScpkUWAhp1Cv54JTUSNcoD49da1Tjw+B
/OGzLujGLSaH94tHZdVPbobnhK2YeKg7Hluf7NB/qVf4kUFLMG+PDxhmKxk+1EuvE6g7kK7uTiQ1
ap0PwWat2fIzv/j693eVtNE4pysma6sATKU7As/BQroQ/HXftB3bD7BQLvb7W2YPzt4z9OgTYly9
IS7bDnGCw0FmsOq94djDbb3vHaELQgyse1vchSYkDfOgJwvk4IZrnX1prquj3UIhSYFGFkx3Ezsf
4OwVkc5ttLMJzXibjAFcJ0pK0DFx38P/GWmQuBtyjF+5ywxLO8SrEUBuZamOq+OUrXipQ+vb4B5C
A4oepF5vjdv9y9fa+BFex9k4s8wTnRs/zijzgqmXxo4RdzSvCTX7b/QCy8OFN0algKH5xUeBAGDO
Hnr1lkL49WKWDLGrfBZPmJik+WOP3AOFKR+CvEczCCZ0zH7bEsowVIajwdyPdmLt75oz2727o9/3
kcCH6zimhy9du7CBj/Z+3dF1x6zjoIhpoD01kzkXuqOt+w77hXTwUmJcv0uHnd0gJJ/WOIou5uNS
bMcsTnjYiLvIbySH2onrfGf7T8211nQwhqe2k633UIOnipyF7a0Di0y9I0TIpiLLyUqRKJ0xzNSi
IYJT1Nr+BsIO001uDC8wtXh820ZEoeViYn4liAL5aSRg8MT2RkiQERtCK+Zef5KgO4g+BJBzSVmG
0Ugi0WRhT88ng5aEdti30Pp3Qg4yJAI0aDDZEeFDTx2WrDd/pOoPHiXi6ySXA3oALUeQK2O/gQtD
6apd3WdgkKrWQ88ErqGLzsyUYmP5+jw/Y7qKAR40GYSPrXKxMMiORjJXlRRonYWI7tzkIgKlZJJO
X630uEgIhP1DATmHgpCrBbvZwmhS/F4V4BfdEkSw5QVVtHRLJFK9IisZZn6O658Vhm7aUy9KChRu
meurJ8w63BaJVw9o5VBCCbX+SmZoYJZR8CIZ+N+sUajRRAaxhRhQpV3CN1DqH8RNOLwRC/agjKZr
7FSMEyHe9PI9uAiW8LCQoz25IsqI0CfyL3IJ7FIw0pERe0480uOaoAO8nf0NpnGJdk5eA98eDSJo
rN1QwFVqEKNTBdvldelXwKVtuB9anarpWiiq3d/4sHu/OQy7F4KFIXtBlhPI9j2quc4v7Ie6qrFy
UToYvabsYuysvTW1dHGURYRbCj3taZE1owNnlHh7SzvVmN9d1ZtQl2+zKR7x9GYr08BNUP6XZkYQ
RfWJ2vn/LcdEAR+ZS5mnIs/jAO/WnAIlv1ozFuqgTPb3/WkdB9FkWk0klzyk+w+SiBH2urHntDQe
muHnw6Uk75jljwaToQP/4+V0nPkXvlt4IVSxQspo9jlYv2kQLuB4vPSQ3U3/ovqbElOuVUw1Zq4J
WtGbXMsL8C8RdgS5vS1qJo4Dg8WcUQEdD2RJoDEFBd4nDFubvmZUhLjIhO1oTJbQ4oldgcoJyg7P
rX9UEpKk5ZFk8wT+E6OiKbi/sMIVZQYJeUxq3MU74MICsvfMnoHZ8W2A8QNyXz1UNTFsfhf78xEK
2N4BBCdYOvAjbFgoY4Nn1LMz30IbMjGsSXF2w093MD5NhEgZ9c51l5ZrWJgy2E3zmnWrO5ScuHSt
TD5jNLY7c7cscqyv0sx7mtHGl5F4SX7K2sTJpHegnf8XmvV8Stg4RXsgkmN2myEscbhWFwbPzIGe
LJLoUErwMogmF1IfNnc3c3iRZdfMxGfJ3HrU4PDGu7k0/OipkIaycvZG9SfM6zroSNjHx9R5V3jo
I/di9RTOSatT/1Ym3uAKS+AjZlYVTbqyuesSdAFokY0yDDkWVIBOHSx7tiINsBoDEVPyRnIRp+Yj
8Go//2HQbgl+78n9gbfMXuUunQJ8JFSbOp0g7AYR1At+b4rTgGcBnvdvf8P3TOLZqztbJZCINnoX
wstO4FK3UIPLDYVST5B2X0pcQ9yOHdTaNLB9pQ51Wg47bNAf9jdRbaSwa7AQ4zzlV/T9SSsdmAa9
28U+6YbIH7CYcLebZ3Uk3p6oIbESWLp18Uw0F/hmNV6+i6HlHtUZt0TWIkirYnsW4nEmbOBb2S9E
TcNEqU9nYnh2HZHFCEE2r1V2PBvLO6c4jkXcuF4VGKShukkKIhy8s3qd3MhsJjUE+QG3992gvZ5Y
K7RwQ5q7kAKgBl5IvxccfQJSMEO45o0YCYzIsmSH1i45slxMITDqmVZkpi3TXaKH5cNS07C/Nb6/
WiQ8B/nkBAX5sAQxMsL3aUHXu1kaJisSUQtjhl0EVFwkDOH8Hjiyo2x3Ndk+rbSFd3LGG2F97eBx
QDWVll5aStqfhyjLd0/Y752NF4Pf+nn3TnUfw0ekr0ntpcTkSZjkPOUPeq4+ZaqiYV+vilZ/8zIe
cUWqy84FLCpnansKaYxwVnLZMRcwCW9LDYInk5DhqAUbd3eaoaMjxyJypn5CSbK5xly+V5ZH3qGC
H6dGol32TbLaIHudypOIxibPrVw5QmrMPJl825vSVTbvQYNGIhSi6SQgZJMiA8G/YnX7m/47PBHr
StpXylC7bniESFbFq7OpvRWVc+k4vWh4AOGp1K7C/yaPgKtJ2ygLfyMXDV8XyzgFmJ4C8oamrOAf
78eTFdCLunkvrhhiJ2Ucp8cxDJeIImBnH7GErPtEcA704l7DGmWmmMAsIZdOBthIUKdYMmCvfOyc
4At2ug3R5Dx/0CSRxyTMbiRJvkjR6O3pRXc586g6eZhEEFKLZkYl5RkmDP/leR4Hy6cQWlZU4I5I
So3tO2EKVvWmrAC0WelGwKSjgG8KTiA11BqH0HrLkLF6w4Famn7wZ+dag1zZMVEXLH5mva9z1jqa
h1ZZUrSs18d+4C0p3MEz1ci4qb2ps90XGWSRzdHlSC6JjufRuGhaJqJzcNFc2kZXTHNjsfyX0duD
0V7wKH/mi2EAk92MOHGoHUkPLrSzaJr0Ynl+vhDbV3H+VcIMP2e+DDWItqEvx7UXsT/X9l0kdk/b
SVw00ljt97OI81Ea5oTJ5bIeQ0gllncYInpRXn9ThSsaAtub7E7pkwGXRsKf+AeV7sAz4pvkH5bE
G8rs7hyyv/ZFp1YG5E4+HdX8ygxbW/l2DsIqU8MNDt2W745IG4MOlqGzphgiwCMWwpNrmuILwE4U
xfrC5hDyvcXylJd6HeKkPJhlRM9OWrREKS/w3g9K3GjBd89R36HtXtKE9/xO04fCVEZZvb8IQHPx
jSvuYAUhM6ElRY9CkJt3bZ+FYU0J1zCWLQsHohbDDKLkyQ/uREgmtQg/BJb0EuMFIJEq0mkGBckQ
7tkx+/p7VysrC5cyKwnQ9m3MCd/A+PNXgfQ4Hy/LwVRc7d7839C3i5FFZb5xU8uu8syoMC6/pCFT
n+lwGxkVL1syN3AxFRRg24yoj3Db9PxxxMUl/r+l+/u4KaGjB0HA+79Al82e9AS0wduBnvGbwePu
9QPIQfUsP3kdTLSInqpJYd7kL7rK7ekiWeA1BNt6nhJvtt8CruZmgC1G/qAzA5ms3TUtlq5Y+Rj+
b6P78XthVyGFzAXQgGQUn2uOuvGtSmlpPgceB4RHIGKTPFtcUtfWJ/+SOy3WEpTeHCwAS3jdT5+A
ZdbVTlqh6ZmIieQdqgu/mlWjY809r/bPqhXLZLBpTQlqnKRqPO3yYCBeIih3eWJn3QdlvYonHWTE
31RtmSPg5FfwlCmAPW9BPsD90nJIyBGIzdL/P2apzNtiNWy+2oqUu80Oet7F/kT6N4Bk34Q+2pY3
+13Rggv5CWXwQju+njctk4wMpCWueNOieW3n0ywHyL6WMQnq4WsVmtkuX48zF2zGkBjf59TlI34B
Z6OC3WLfwUVsyQ4fNFxkQ7aNaNZdLqtYYK6q+0ikQPOOC0NkvYHBPd922F8SpUjCk6TXoYSphs8w
p8Bgdlat2JNAX/z8kZNqwUrgoNRt/e8uIyQ1P1paXyXaxbSm/wrB0QSQUZHTR44D8dQmG612SpCD
SZBwvHvOh/94jEyzMotoxAF/06aVLb69/BySbNTscKk9NWOlYa/4wEaoyNVmHDq5KD0tCENnxxOf
gx5NQAMY1SzeO5p+zoCK1N+azmlOjncjzc18jt3Dszo7gsvE03xXX6rOWyFyeXtkL2sG9Iojoxze
X2mq92ZvyUpqgt4DzSydZGYfX4oeDxv5+aKtIWQ+SWKFlUJzndjk5sUEqGDudgvpU2cWE6umMKKm
JFtovzUAQeQd/Tfwrtb878JKTULgDLOP5hY/3a533JuTK9+gHzWiLL/nIm4PwX3BHHtj6EPnMRT2
1bfvvYEl9RHeQ/haJaUsw5/kT9DEk23ztMCFhUr+/0vsLWBDMp8F8Fno7H/IUzbpfZuJIoZIbqsY
LMrPWryF7lspP/TKWHFdTBVzRPbxea8z5pkxgX2XPF1M2UGhzI7yme+6dJgxnkaDPZl61fTi03l7
oMiD0OQD9x4MHT24cG68WgbPk/+tgzELmIXjhKGm60G4TOM9x+coTM7X1u/dUyc2tNuetoQgT3pZ
AoFBISBAi0vTqmclXYapEc+Y4VCndcoGWLipI9LWW0qgNBijcgb5Yj2r9ZRKRftmICQOsdq3SRbe
VbREGGfX0p9pyv9fVBW1g7ecAaarMjFEoN9WwhPyKJoVaKdkDesa/NFxpsF7KLt8r1+CiYkrLfOt
y368H9dAmkCJ1BCgaoE/tS7q51DncBKyiwp5GtKXtyucopruChDO7ch9WRAv8IsG1zRaMO7owNVU
P3TO3EXyGsqbdVapVlNVWVccTxo6HHX2QNDFeDqg+fvabJswGhDWcFg5PvsKvQfZ+T9G/CZGoCwF
0CLtp03c8JZlTyedC9Fye4iJ8OLC1QU8iR1+k2yrkXOHdOsR0rZGIh2nCVC4yGL34HXqmFsd5djM
/2n2pZwso1vAhv/dzbBhfqxGfHWIkCiKfGM/RkbOMjGETphrpUd31MOtGCuMzhgfXaFPN21s0aRL
WiuHB64fc9R25NEmoLPc1dfsRrucRqjPefUv936jPQX9YxiLTlodoXo0hY7wYE5pi/ocp0xLEoLE
XVj8+ThjSVoNit4CewRZIf3SzYREhoni5bSjOtOuOTmaVDuM/LMcLobfXJhirPs6dpEapdugb08V
xKzGCIwuAwNkEnLYSzQ99Njj5Aw5OtJkUab0J/HT+RpqS64an/DTLiwcwLxYfdXuB2LFPqU/oTpg
B52xsBStPG5PNbK0O9wkBfftF+nzR7NBQ7mXb6Ywru/Z+/nOdPcjbGqcaE3x/U8FbgRM2UVXiRBZ
Qy/lJMd3r1SIPgDOxQAnywRwipg9jdsEPzuHz6moe+anbrX370RQrR9GmT9ExVQvS4btyeW4AICW
DaJhBcRG5QcDp91/30yCEWenUX86GgHJPWbh8JDgp0L3KLWsRnZe7WiNv7KG7S9cYpl00Ce7M3dY
8F3t4xDzPzbh2PenIKgRso9dB1EC/iKzZa0S/+IfM6w+xth5uA8fmymbDr4iZg3VkQQ+AbSJcfoZ
WifSH29k4h5PLhp1lMps5r86QDTXu85LbJX5Iw90+IDsH68NzjrAd6jgB21IX82iFsglGTdg7I8s
Yle9JpmvxO422qaRawEU+NmmdIm9kcfkiOxqZpJ/6D8vjvLoOtJ1vxMt0OeV/2FmXFxrtdJqA6be
BL04qLJ7LwMkqjagXEixHp/SOc2mtjCM2JCQ5znLgAikGLPGZCGX8s8KV3dUuGsOblMm4ZgsenQ0
GTNZRYP0ph9bPaMfEwkpsch1/ylCAxnp4nKHBWZCVNDxCvPLtqGbQ2sNnJ5GhbQzAHQR1tKUJ9X8
g53rfQu33RVFs9lTCG1B6Gk5eWFOeo7Aoi94EoDG/0ieur9lrBbrobS/4Rm8JOblenhGsv7W2bHA
Yf+oRtXMGXRbPf5/GxWa277a1fIwo1pugcGUpqKQpi54ByhqC2EfSiGiVoMbOtxy53l6m/3KOXmK
NAP3bcepfG3ofy9Qb+JcaOguNZs2yTGdp9e1c49jCd7TeH7WgP6jXaOTLQWrlZgfaXHCCy3cTs69
7b3Za8PUj/GiMa+M9Ign3y9U5v3lmLqTVolvIWwdlhUyXibkTY4tBm1xm1GfiU6K1WfsvAy1Jhso
ck0JRF0V8uZchERHRZMyUMRtjqJX0QZYV59ud1IrcXl1DXX3aRkjpSXEZpXbtTTpQ7vCwQAr0nrq
89oY2Xc0pRPTAf5MyHeH85Vb5/4d8Rmb18oCGZAAhWcmR4MEhuHdRt5QP3dwlaWyQi/31vGX8vEl
hv+jX5BYX6s0i8a+ToFzERxYb5ay4RHDBZ3Km+ezQ+/NfRY21a0wKyxHEfQnY53eBQR5FB3pRG5g
D/kxX+V/DF6IS8NuNrjWD+0X4SgSM833sSerCRULxlirXTHcGXISvhrvRuRxr8jGRH52wYWzvAo9
cr09IDusRKvXjRr+Zg70/M1J5Eb1cad6GQ1V7zOgbtJNk3E16L4rmmum17tVTbAKhy5xjVUPeVBe
/zQ3zxaG4/wU0HJT50ociJR+Ze/kbL9Be8tViY7qg7+UliAlUIt1Fy3oVYx468dEgzCx19ejiokE
MvaBvnVH0p4t2WTUZL8uxqDTtNvulZcECZi1RKWTCyFC8mX6YvdyinfldqbjL7RlGrziT/MGlKbC
jk5lK6ISGzkHf9KCKaTHoWjN3abC1QUXUHOKkvtZsBS+wsu5GwzGZGGFGG5iTUSPcTQOg7OKGFno
apEC1J4KtoBDOiTlUDPrCVM6KmR5WHu7HwzY/TALP4VuoVuKRj+7pxWImKm+RjBespru+gQScz9o
PCjW7plhjfyMyY1AI31EtRiNEmJZ1gzPGtxYMCKWU6Cepe2qrXDJPdc6F+J8SSI8jKp67u+JMM92
zCzMn5Ly59SGdAAHIX5yLcwdwFAPPY6govKFEXjyNflCSEwXdAhXD3rqwUv+bP4px347dwUDdMDu
wzViRcSKtjQrihJLg6DHepKflgshA/SWYgpwaWcHBurQGT+CWFg1wiSm+8QT2IFjuKRViRP1J+WF
ANk0k9Eq5Uy7BFjSJkREReKNBbw2/DRIlAkMPZMqrbqonv7fV39YzNBXm/m7eS5xzMw6ZfwJidCj
Qv+Iveo0afHJOoMAofCqKdqbDLH1Y1VoxvHLYRyNrnEXXRntETQEp2Csvi/affIIMFZmaNJ4t/RO
bR/e3NBOMFxGtMn9VIRW9RfZ2ERfRe8PUQkzI3Y61tuyrIxntyNsBUHh4uXRJwFLqcny5RIppOwb
Vb33+WJdPa26QAM7Sy2wLY5nYnWL3S06SOk9bqZqBCYVB7k9zeIJSY2eO1epSj5UJCuMctwwPv1s
zQkWbMBvrHPubqXFIdLfLdzEPRQGoGdW2gXXxMI8xMPqH9MYQV4n4LHhwMofGlfOXjPOpGKldDHJ
Mwd+E7F1OLBC4342SWf/Exno5ohhO5OMNfhhiunDxtxJPTVdZWp57pitLrJ6v32dxpacsUN3BymM
RP8nBBPZwUWqwqfFkCU/GPccwQJeLMSM9QlIYaEn0UnxTg+JVZ5NiItUwHhjfhuOaSqrkLx6Xbe/
es3uEz4bviWxgSNUkSCTVdn5DM9bWsq3XlCMMFdCn7M7Kp80mbvBtOd6l9lvWW8piY3RAYQMMkjr
3m4tx0vVqkdWWrZG4gR/EeWHWmDxhrviJYqaOfn5FmsrZ8ezJiAwPdSynfHP6XCJ77d2NdR3s5fL
WffArZzyuwRwV+q76c/ZATBAbclB4Bx0Pc5L6KyWeKyWm7dkbU+puSNgN0IM8w4Uo9GhsFSsxadJ
vWA4ORtFcwDshOJ39wuA+PAxlX7l5ML1h51w6GVGcJVIXmw0zNoU72BWlu8B3kgS6hrNXRfYOZdz
PTkDOdaHYa2542l4JC8Wxk0uwHpMJaXVewVH/Q5hotSKL41NehYmk9zoN92a/dn5nPVndHs8iyZJ
2Hf9RGQH7UrvYk/NM7/31CyhlLrQXJo7c7Rj/Kh3hXKCBNTvJbpYxXdeP61uphC1pZA3MUnuZyfX
jy9WztbVRc5lQz9hc2fwZqbhu38euD/dRcMP7o6S5w87bW96V0FNHEO6i85CXKbOIeGvHxrEsXtK
i6X7S09WxcPat4GBTqJ++gFT0aZi3FvyK2+TCkuVSEOAN7D65/AfAOMr7x9UvLtV1BsOpzhky9EQ
q2n+S/7/6J0sc6r8/gQJjIEwyHe9OVD2jP8Sl0np5qwcnCSWo6H6LkREeHjEw5r6PIQ6cmWEBx9C
GHeoUTHMf9yrl/RY+dpBXBLuPeeoCApUR6/ChjNsKIO4c+vA0ElBEhKtl8jVHlWXms1y7pwiJ636
SxV00XrF1JhVy0hylmCs3ts1LcQVLFK7CRB7hqqiVWggn3EvIeEyeYCaCSEnCOmThki3RwFWsGTM
eNAGHFMoAkFVkIfoDgriacp+rKgM661KW2GDiw8hDvlxDzeNdqEFB8nh1jdJFRNgUDtm9d2BeP6X
rZIMMwLjc1njeDxIas7R0BRYGiMch7A1UiSwabKu9F1bzmFRWq03HaJssPyTenewBQ26v6UemrPM
4+gLV4FXfs9Ab0OFLToEocBlmh+bFlzLF8R2Mz6kIMEuaOPLF571gn4j1G3rsxeP2L2EuIcl9zSJ
hOK3QH/2AwqfLqj0h+dju/54R7kNCJJH5D3Wj6F7kyruEuZe5munfvqPVIJbzNxsBVDTo5Zc/aqA
+cvbZNcU3ehzBjk3mOgrJ9WW2pCsNIpwMOJeIV3v6OQe3SOCVNTVt5L4h2ZbvFmsXPJhHjsw6UPK
qjySJM5G+jqeVugycVibUhwwz+cOyywW8rIldCoYZeZxuwh7MvaH/rdd79wDndu8gLLyTPaKrbcd
WVnKUGxQgLSQja34VyUVFnLY/Bbgvegwwd9FD75mgk4Hfyj3BW72yROYAYEDRD9RID6WRDLditTj
Sg5oYn9yPjBYpa16iGelu0psLbA2y7y0J5sIz8XBzml2yWrb987AKhIvO86qHRmYhTdzPi4hrSnJ
JirWCfgFB3hmD0wTvj1zfoEZqdX0uVYkYHH6RxoFj60aRTqBPtS2SqtpFfXRfRYEjNqgMpMf8vyh
MyWoS9CDRBBmfJdGO6el2GuKLor5hxSwahLyK7Bp9KMKW5u4kausIMo1OrSZzNVYakxueYD1M1Gg
D6UIDUcrWqRNic3fXw+1UYt39H17Bc9+lMxKYSAchIX1t7C8zt6HTj8LHuMw5Zqz0wlL3Zr8zIoK
kSEXhY3rp0MI0K56OnMqNEGI0HvTxy4Srik4xZzYnaqoU/uSauRhxLOvTpPowlDSVXSSJ2ePEC0q
rP/3XsCr5V1pERinFSWQfqT8+yv918XGAoKwm7h5WjmNKXymsDpSKqFbeWti34AnK9kwzTQCjJhA
Cml38A9eRJaranDJqxx5/mbfCiPw97li0gB8sUlgH/wzC3eRobcxI/fpsiiW9Vln5CtRqHO9PF3L
A2aTQ5QuakVwfna5bde/ZC+cZF2biZzXoRxF0v+A1ctjPA4Qf4vWBKqvdBAfXljpR/C9ijmVM8LN
tdH+wXUlKTcSoaKQyX5avc060u8b/Jj/rxYe9SLaVMgPmK2K7xkjWnQGzh2+n4dbKsmw+OYslJbd
Y/C7fdWQRCUuPQIjKg/7EgI0LgSLRwy2a8FWtNRPb8J/bkHC3Z0U1oRCanU7Vh/P7MZrC8MTqpB3
D6wUZtxC4Eg7D23BqjyPKF2QP+0wRUibMj7MeUHX8ASKCTji2khQKkM6gkgKL7cWbD53Ya7LEu11
ROSAvyKdL5aY8rw4rGCyiTccfP+YZoWxEqkG2i9HM57G5mLEOUuRMqNfz+IJIV6lR5PnA6eo2/ir
/plVZz0zDrWgZ0PoY+kTpfnWR5FeUebmy2IrE91Si+0myzXQ/nh5hn8DNQzqyEqv1JWLn6o9DB7O
u+q1Wis14FVsg8fvs+PFajp9CkLtVftEr37BhglZwyWQyGgRTmgPx+FMsYVwzWi7jF3rHPnKbMFV
WJm8c/C3UPtOli3Qe3RkcXwiJ63qaKOL+8ONpZm4zS3A1eeiDth9A4JPEWka3+dNW8YAO3Tw4FyK
wDOkO4VtS77O1huD1otPnpn50TMfhicV69pSyJCdamEp23iGia8viF2WSdkD23ZE4XSjVqwsvTcw
/6tujQ/L36q0D0bsf/i8kkmDDfIbb5Led5I/lYcmXSMnVCADOIhQuyK0IsQo0aWHXBbvTSlkV9/q
42HHNsxZ6lPIhPoTulv65pzr/A0KEaGINa6Pu1ekCjHmUNuyF16EjeRUMw2BuK6AQevw5bbvlj84
XDcYAke40Z8ot7ouhVrxWF5iXl19wcI5IyvPm3Q1eag23wNxeA0UYWYE4NOfvPPHdHsQRKAmpyXP
h6QLzalA+OqfEJ/TRFMUeNLjoZhgAfWiDZTMK9EWboGJv/5U7l1qiIar85hMk2vvJgK7x0wk9goq
nwupasnbi49p1kwtnrwYegHfAfiQRW4rb10QQqpSBXjAMbgiCOe8E5/CcZ8tfkMdYrcyMjsvZLFh
nxjYpksu316eXBVN37pmpJiWxcozN8YtInfga00uMIWkeUMxi5Dk+NJhqtQIHZH4cPGvn5rVXXOy
dWJML5x4W6EKQg/8dwUIACTz77kUKUKVsj1X0iOEy+mkLwvZz5wVE2TBIA4f4k8ckejEmwV3EJhS
cV1Oz9IL7vvlWWGLr3Y7in2UQ/D9ZpAMksFYYHUXeK87t61GLcO6/j2Eh1mjqEmcTvGtYn43FLxX
uvDPObjxExpIE84dR/ciPpRbAztpHAS+XhduAIL1vOZHw9lT8ryLTbulPznt1Tg73mfKPE7hR0+t
YxlGVE7Np4gpQApI/v1FmvJa438+uKIy7vXqLLpsGVmiEddWQZOPottInwaIQUU0Ue78LTt71CyH
Tg62gZwcXUz4VeO+iwXsF2VYVbF1LdCWkUP8Hz//nWmplmMVjStXUFRaD0n06JWzfKY0K+8g2OtS
B5deENYvOdOqAqmTtuI2bwub/iru5EH8RJxpSqICEw2pHcU0ky0ydRTNxFSHibDR/79ySnT89CXe
kkaiExBew/EeqSB+xP1mOdOu/oGl4xAuQRerCe/1dZSjHeKpj8+4evFgoklpWvk/jQF8pVhbNvEH
oo1wbPYYkn/g7fQWrJVhLonc/x316IBMMCwFqzknnoQrujHdYBPHzsScii59ns1XmJP+NuJy7VDU
aRfyOlijLPeTeeeyzY+/uCObQsQVuX9duCn5WZEarghdm/hqUpzZlnK78m114C11p7pxMUYzBHvn
ZNFnpGMGlUOxTdV+9B+Bph27YnFTDI/xooBLFJq5HIn791MaDaspAlmeJ9RBd3GW3QoFg0h1zdjE
6QAeD8YAwGpEv7bekjgUFxENFh/lzm7yEulI0ZpS5Z8YBl/LfzVO6MCmQaSnRaiMvZGtx7ybFDLs
9F934qABu8yt045J7tk63GTaJMq0PZOL3E2mVsMqTNUFebvxaKWBrbvQgSMYCLcbV/+MaspRafbr
XcIT+fl0OZjvsS+W6rWvFTUqeANBxeyW+N4kVnMkwVh7CSY9IEDh2i3pyD3MySpyEAzgR4NQj3bY
krRJppJRLE7F9xZfRG2Q9ZHwBOoObkQhHrcVXX3gOcawMUTtD5cCyVa8qcKmct4fpkFpkGkHGXSs
GiWuJ97WTPb7e4hpBFdrZ9kmtByuyTp4lU7f4L1bsffH/UV70jeKAKTC9ZsemI1LrPTVlSk3uZn0
2KJu14zkStF+atsDuWBfdRo+6n1u03XJzBl62qxk08MFMdYTJZNvNQ0qRyHbwUgsIa5WPS4TNIof
6mhAH+dbP87oks+uijT29dnvezx/aHBj3FhWi6wLvtonAd/B2qvUKJc3ECh+fFEoZifXbB2Ha6Az
ccFgHnOewBNPYasZnqQZR+x67WcXmr8vITf4dreP+WpD1u0GJC1IyHeJkNo0OCxmKYlPmKVeL/vx
6Pj1Hf+od5n3d7gDGBHPxl9E/W2ELgA93FvSXJx1za08VdD/+HLejGZH08I17+gg/K/KNNzcJdxA
JNOxzhQ6qj/wO84+d2EkhdbxvaucaoTba40HKzglJmYmZt2ofK6mfJxX180FPCGBFIJUCFfzGzVE
jjd3fbok8R1dZmjizwjuccsPM219GOFE/Tp8VeqfDsdAnuamOsAK+7YVDav8qaaa08QFAFE3Z/ws
1tLtUI9xniRL6Fdfp7TL/gvLUigyNQ2r+LbmBnB+FuoVbsUK4UYbevuGp1DAuUJ416eB/Nu0v8Xw
1n8CPfCHIwjKK3H2rJY7HUJFMqsSl2utoSsSVb18AWBUUFpZzIbKB0A6B28uplDdb4VjKs9yj/zb
loAFEIbQfYOnzQQY0h0fKGs0i2mR26x9h0yGRCWFg8JylzU0KjxoKoegOnA4ML1r1B6rPi8xsKKe
8qYExF/fqo3HR1B7zbKziLN/DBle1gAOCFUMQa7RCV8H4o0gi2wFpVmUeG//L4APQHt8fKX0MJ7I
l1jq5dfIDuexxr9TWJU7RiBi3dZdVbsjmlSi5wo7hrTPsoo6z4WBUCXmRLIGZnZ5g7fJH6Z6A4pA
SlA2+8qBnQeonBxR8dK9E7nnsSJF+HLXEjV7tURLK1dp99tbpR5ky0v44rndUDBnXvQlJVMbnSLd
yHiHk1D3skxbeT3HsVE9Es+jznh9WgMOxeSTnbvEhrIYzDlBzdaSEO1NOF/dY8stRGAXyPvXbwU3
sYFO3J3goRJZAPKvKOdGfNsdiQyi/yTE8dB8FGW8MYdLrU9TbLN0GO594umNjATo/tmAgqIYQOg5
1iyPMWqVrkn0TWBxKm07v+SeJkf2U7MsXrIRc9JRmNX5McfKDnhvWm4pozqw1wg5CZwQIFvAJacd
QYLNqNoD4xb/WKHeXSfftWnEplJ9FQVJ3IPpTZLSdsc8qqXS1R2GXzSFYd2PfQ71LWaHIe4dmFz+
N5cWgh2jkVwQprlxJ8tJajdkYftNq00oyGrH2VWYcN+kRRcQ3nxGlYxsEa5+/8sYXCwimVfVNZGg
TugvNryWqOas9ZTjbmsA7QdRDB2tySvjOHZGCD70mA6r1cFikTeU+b83KwFzZQ33WH1qYPFL6kOx
KBIRh8cByKhZ4VxhGTRNgCckZrAB+/f8RH5Afb5Nk0l+EfFg9n6ZbStxsuKDmzL/pC0VorV+3MoY
hejfFsBam7zcMdX4hRMvtT9KJBBuuq1N65BBkyzqXEz+DKJCKE/ZsNJ1AjDr/BEgT+kSp28Yt/Tx
ItOdsH629tM3cEyGZE3UZJwYA+pEeS/o88BLCACMvDsGipDAd+w8pQT0N0g3sdYYfS2wjGtNDEuz
siI6Vgcwyl2I2GCi6vr7df280c7zxTWPwnmhnu46YBrasDrUSHm/R0BuYS01TNK1e6u/ZLmOlUbc
FliYnzGWuIBV2YsBfXZQn/CL9Jla01QUZCY6IOez5VYDnckWtclF6RsJf8KuY4x4619ahSCsqKX9
tcPKiXJ2NcjmUHg7zxd/fYD+NGLAS2cffBKD89f1RlwnZE/7tXk0auBmc6UNnTW6vfORXBXyAcAB
4nLQ6bORZwYqQ9Z/3P/oWasGS6wk3Ftz1CYSW7JzvwaWxciR8GFEte2o7qNHBqbRcOUsoyFc1R7Q
YsPDiLoRrf8ncEzwtXsyFFtlg6lh5ILCCEt+IKO1KZ89KeuMhkBKh+PebYAi82jBMRaXFXfBCH+z
IqlrazZlu5XREfrAUGUXilk0heC1UwsDxLC380t2isgVDqVr7qdde8mD/UmwGovOf3UOzMCAJOyz
Fl9i/C2iYnMY36kaA30TDRKT27kpCE8DC9SwRMHoLDAPXAT5O0ih9Wxa+kWeryVisn288mPHOIRZ
aAcO5S2VNgUYKUzFepVik97TX48kKmXgtPYBMC62SkSyJOmrgs6t8C9tY8SNBaZ9qUaQ/zEUkCHL
X5dJJEdi3e2/ZZ4uN9ZdqQDDWtAMqBTfTB4o8n3+mAHwDbc0yM38j5sqGi95ByttlSGbqpbfl/Ag
ykCFvPjQaNLDZkOSN3QdsoZI2FW/X6d1VVIteoGiVNoIQgc/PRRyYR3na51cYTVARFlF28lNDRd/
8b31g8SsNmMaJg3wIbkqMCkiiIyF+19Tqx2oBKjxgXGaOKCH8BiFz3rBfnxngoRPcxpGgox/exYr
ct5OpB3IIsUl40vu5h6IVRwNbI5sKc3vjdsHWyCQ3sgrXFKnCTK+56ZCc12taYLT+uBxHy3lryym
23tN2lZG9d5toWVCu7TdJRr5WotjBXGRLO9MzjQg29r3bUuGDnwCzWU/MKRKok2YYSL80ireR36m
xAvXoSVIdfIsg6RFXevvd81mqCfpvV8/XsNIADtCnILyHwkeXBkpM/TAgIoM7QBW0T2qWcLRZmuU
znXluwCGmAoLILwEMBFrWhLOMx0uJlelWAgP071eCDYh0Jnpu7bhafdM329M6SfD+39dkDj+lJMT
Bhl8RPMPnReTfhxFvkj8ikWafjzCvUTsNzmxAptIf69hSuNbCpjJhi2MmnosjyB/GdN7m9ijtE1O
ClTfeRsZ2KvgIycqln+TztJw5RbwLltS+arWCndbEPRKuz2Ea0wzko0FCptFgtZ0godTRcasSq4l
mamqzhsyOXdqsGfmPhrwmTMdSzrexDSE9P7DeCkwGh0jpGG7VX8vO/EEgxFtvf71sGjWaCZNQITG
BE+yRaxwbNxiEIdSAVpZHXwhptdTdqHdT4e6+e205ffZTYHosq3jsBt9dTibnwn82j4V11PkB7O3
VjU0mUJ5HYSoN+z6RphqPKyj2g8F4fzz6TZgLeRyzy4f2lkNDkBK8gON8Zdo/DFCa9XzB28IDmuW
JJOtFS7eILafFbpixwwEJZD+L6w3NiVU3v4bc4t2t2lFFnucA4sOfxr7Gbgh8+iItnTGSeushBe1
NN765cMvcOGzCkH6MP88/BNawGe/fRBGsP8ZW5O4+dDAektACwUL6FrzsggNMHxAeRGd1qUY4If1
3myA8QILgnsRGb7TfT0I9B0OIKx4uuq/SU65hhzTG9SQOC4D+hfnPS38fjUBSJUAQlIh6i83Tk2t
Ayl01y3kSHE1R6RJNPovAVeCYSTV+eoemqAJh7oONl7fOHtbLtWt/2zNosAbZnPSbjvJ6iza1qLL
eOO8/DwD2Eea0mGHH5sAdmw7zgz/NP9kXaVMiYnHJd8TLC9yTPwHEFdmlS/oSzHRaO2imWtCiE87
jGNemBa/yfB/jp1i4UADK1wCJvv0TgmgC/9FH9Vh8rsbq+zG5dKiEVzqewk7SrxjSwYtrTBJiD4j
BM4wu3PQahi8/YHHp/i6njdoTt5j2h7yx3Pfpr0mhoE2nHCqmOTXLAfflnGI7kOT1e0SOy8fBqpi
bmxvyFp5QOQuG14y75mVgPefTUuPKSXx3naK+Ol8o7bZkeMP26C14p3+fmUZwSp3FDQwNH6m+HTO
CPuGnb6oAWgEBpDb9Zg9dDKwWhMx8KQkJuocq1lKm5D1hvTLv4Zq78pTndZYXnKnGZMXsrhDuYWq
mmfdAl3WglD3JtRUeP7e+VVLSiFS8L/R+j0m28/1VD72RONd/HEAlbyjEBtXjazLXXVSo3TQZzto
rgn4saUOhhbs3ux/3r6PXArST9olJZD6kl4gtby188jEPJ7/xyk1nWMvCn3mZCpV44CyyPTgMb6+
I7ShNEEK8jCQjwsDy/8wcuT+i+ahafjoakpbsYQPWvj1SYGFAIGzKbGZCgGYmimAtvfigeaWOhj+
e69awIP+b5AaSKhRQnsd34X/H2YUqfDauMyIjNcxSJszAk9BXVptIKF/ojGnw8AAztCPAG0c63Vn
KsZgcx0EE3PrDGkSAg9Kfx8L1q4TbdFwUsgy1yIZj0ZN+ey9CS2CHAO6Rm8iBc69XZT7cihHHJNu
nlQYoOme3nA/HSmn4xuD1hoMX7l3U8KXK0CoHSrWVdILv/lcF1j5FKcNNcFPB/LQvomP16Aq12lr
+jhLQXKvyPwkmcnyPUCQ5jjAQbxoRHhLwpDozLIjLZJ4sviu4Qc6ZfeknAXE55qY8C0LAib9g3ap
mpb9rA+g61B+dAs72pZ5xj3i3beyEa9f/Za5YsCgszOUr2u1Yp0u4DE487gV7E60Dp826ZlZLE5s
MZM/AAit4vULNzLOFSpbijwG0fRPIOllN5bqbRtgb6sx2JapnNpB3RWwmaN2mZSfWeZA1YINJdIu
ZNlLIIM+caE8Hx25ineHD9jq68o5Fa6hDmwt3hkN/ELzzUoNDHq2SKOdAAfootljiPsfjMUaCjeY
HWou83ThvFBGTCgoYPSPpHnGYygU8lVEECcIp6POp4j0npkEQ2XZ76VwP3kO3EPmp09FLz2YzW8R
O+VXCA2Hg7JaO+XdQfeSs1V9+76iUvrqTzMxA8Awk0KZ5a08tU8R3E9a5Bt1RmKMMfw/ljwjWopG
gxjps1wNdUy7/EdozgTfOMSMsLLysliLft9ZLGaIr7amLI3Zj4WEkUebrg3UYLyNUdAeRyK84g0x
e1F4iC3CSuM08UdTHm5XSBApy9tb11VVfk64d0HaKEW1tJUOu0NpY3n/HLa4Y3FaaSXh6ZKxHqtC
y9qF7jPjqXJNygG0Qh5NniGiqitZQlv0EpxyY+Q/0hi7nYhMosbXwIZAnw0fnKJC+kq13ARHuFTU
qTcCLRkaYPS7kyyoAbwJ7Cx8OfE4lVv9GRep3iFbk/9WO//aroHzl4VickOF/eSLcaaqVLuLyhoJ
5+bEkR+wR0rgpKFZAAVhwOOHq8bzEWghHIGdc0o8am0l6bMaoHpphSSGXVxPD9ItYzurFpJZVt8B
OsJ1FTfjhMfW0j3ZMSWDnIrEUNx+qY9WS6sNj7dW+T73fzQelln/vL0AwmSjiFwdaMibvMA77Yrk
MTSEqHRpT+l6nvYLQaY80CSA6iYMvdOJNKA0v7hKcYrcsLGkK+1vIPkDdSIB23ecwjI3nW6L+6P0
H1Fsp2qI8snaL9Mb8oX7aeV8Y64rNpqxnIzCFslxZz52EWFsmiW8o6ygY5CoIr+7GIFx7LMYk8Tf
81vt7/a/CISBzOTKB34jHnX0KzRhT1whaeq3YL59rg/n9IllMC7yVqG9HXPCdSX4O/ZxBo6aIAj9
yig4acrGjaCMNKGgZRQYSgjPpRMnYyyp/8WJ0U7eQzW6F9GzJV31HfIXMAiE6mezqJLjCbpTmov7
QyD6Ci/nd9qLdbFxVTl90y+sKITsO7xPFNCvaHQHfANKD/WOrxlfF1ru+5ejNht6uNHlASqpP2bl
J9s+VMPA3/j8Em1aEhv8nZKVJ51CIXoroG/v2dIT3KBf8yTUrbcD38CQrSw79o30+sgRriQfSqhO
45IbzFKj5iZRn8x6wtxEd1l0OMQkzKUVPifboxDzgi8L4qSo4OOYc/xLQB1EdqJ5NBfELOlZhEkg
xBpR8SRm6ORnlB7bLUTv5SfeG/ucodrBOA3mwNHGJ2w2rgg89zSgXGNLA8xtlTsCgijz2xNCScFE
D5zurDrcxAr3njQYS/h3dwP1LL12s6CSFGBAq7+ZR6mMNBQ6grjd4WWiIEgmZG09wUjra/Crd5b6
l6dUhLOSh0WFFBM+Y3qSx2INt4dcomNP7reTFWoEqisArRQygWE0A0thBgxin76S3lgMeVK38sv3
0MAhwsSG5hEFzeCexXG0YdkV1HIRbYgmD4YHt6sRHAEUPUYsifAJTLja7+uWk99/I5P/avTV1k9g
eubLWH145M4kugA4R4nDutw940osvST1BtqqHnD+5ZW7VE/olLG48HJ//I8lqeL8Uug8A5wOKdk0
30hXw7cxvaA3T3jMRtKrSsgjiBmVdUz219iVjifzb5CJv39H3iOdy+gavABbfBEKaJkh1dOC8eBI
1ereT/gtXszOoN5M7Qpv963kxerjvL2Vt9kauR9EgiJEEAB3DTw5MACpY07kcpnL0s/CN08+Mkmk
LYG1soTCioRlAYCi2u1eTDuaueoV8UJJZKwHLgNiEOaozOS46Lh0dBU7DUWOvgY+/Mm3hB+x8c8t
PaH4GXrRX2j5nw9HOS+nfhTuhKM18UE4rRaasHK7S8uaVTgxSZqL6Ermdn2z24B7j9rJDAku6P2A
3MRcEWjFRKlXGoZg4nNKQbNiwykwpWcQZ7HNxc45MP37PTfbZdymkma3bdVB68GC2GVaUWA9hrQb
sQm22DP2NFD07KszvxaNh0+uGlk+MdYR5F9sinpeNCyREDw6pKCo7QpW0hOmvqCi3V2+Uf+hYJb9
0zuVJ0DEEQmtrs1jtdHYQKRvNtMJFf9M5UsKQ0Plcmp1qjulKv8496tOK57yi47pNx5oZtlDvjv7
SkvtWBuWbyuZsz0cc1C8KBcVv/xM99VGwHr+lg84Iswb/8LhB8kZZ/kK+m1In9WRmigrp0IGleUn
VtC/tK1TMFEoZL3yb4/fuTiAK6Nz7q+yTkEiQQROxi/yZbG3NrNUOf9agCn140Lf+dfKuG023spk
HzgEK10jlgfUE8qxDO0BeCJ0w2fvdvDKDrpTtN6Ki0tzd3RFJlb7E2fn/THyHYhGD3eFo7Lqe4Y0
Dw2PHLnt8kbdgLP4LNCX6zKfFh/GVuQ6IGiqX7m8TeofCcoxdCV/tBDtlwwc2l7tInDsIpCqEOMY
YbRVi7+d5M75bhZo8g1xbFXyM1URok3c5HlE+tFzoBMsWx6weW8vzCevvngkzrPj2pYo5O+mc03w
OVSqo7JBHIWoBZviIszyQrDiZ/GCgJjaxnD4ktIQbVH9HDJ8KzJytqiojKFwI7hmQ1wuj4du6/Fz
mu3TBveDOaW9rmvzg4xhdu256ngPic1+1xsPcHAIyxzetvOM2ocXai7Zhxw++9S2UytHh8PvMPkS
BuVpQycmgoB5/TpAuMTj6xa8I7rK7iuhkS5xEk7eaGYfO/BgXHkcJUVAMWpjKvgj8gOaqGDMuw0c
9PIx+PHHMn/UMU8TZPuRoj6vfo9v521Cf684IKqd3jgI5/SwSpkQWlsI4488hol7dYjp1owYcvA9
FjNnh0jLxMfnfVZfj1X3FywTwjJNnUobE/P3Yvkz5LjKkUC1CaRzOIaKN/pjwjDLmlHXPyZPeed9
bHLc/8OMyNHEVlQkrJWI4eILBPGfhax9E4IkDRpRbm8PzaSLMTQ24gP9wwK0NGB55wOF3Xd0zDS6
JBSwjrxN9ciwraf95hWYglvxEJnqaXr1M5VZ6nR99SrpCKoJtkgCS3OfPNmcM2i9y0nn8z1yBltu
wjOH3Zc+yBSAfanGCoNCqiSHOMrcX1+T/mpW+O2xnU35in9k1f2xHo5X3PbnHqnj/JqEcVamig2b
UagM8hxJStUUTJVXKCFGAN2B/TLCyyb16j1eqydJ9pMnndeDeWO8Y8mm60zt+mqWaCTeekJq3QSf
N3OS/9O15xm8RGq5CLQcQGVtO9eYcANJDH67o9yF7HqZme70jy1xMKMLpnxmdb8rz6iHnaahT3oC
rEqYr5m9Hw0QxYoO0ipUqZom1OeF5D+sgOjAfqoT0kx89axsjspe0zEW397LoF2WilJOMTUL5XRd
4RIHsGbYT9fzeYHgzn3XUtlCclsy9k2YkLcjBhVcj5przTnR4hUoYsWbkWOp3FZFm4qoC5bdoolx
AukmljSB0trpGtA198oQ2gpYaA9zacjqZh2EdW4ixds3zZoo4efDw6y6DRsSqIHKUQ4n30P4BBUO
KnmBDR0L1f8d6U5MrG7Op9BKqvcDjlV9FO1k5O63cm9qSGFVqhCc/C4v4DaHXhAMKTmCc8Z5rH9w
8qh7b4sYzXzM17EErjOZGcirdt+DTY/Gg+j56QaU7dbdIVxQQt2DhAlfY7n8A2aKErd1Ttp7bskN
10wNYaLuoqEr7Q2YqjuLI/bh9ecjntxthM9p3ON00Ldyt+NUTFbKhCSHax/l7A6r1a/2qRoO8er/
gjPcsAgBAzbo9VoybDccOkFI/WJIGZXNN8TK3VVm+3bq1Uc0nDVTJMFajvA8dxssCRNyRrtA4vxL
vKjFHNiVTfA3QikTvQQI3zynpCL8tvwNcnd5SjIcBt8Aztnm/vH0qjLMXgadwm4UrJuUB9Bm4UfL
Ba/7UxOVQ2A+iDoFC0cUKEHzeHImSyooHWvuvSHa9GQccio/DikvwtK4w9CC+/QqwR6w5bmrrQAM
ZBr82TGIytXKTQrHcuSSlMl3y+irEtY8aX7QZzcJIDOgaO38m0ElLCCPrbSyUZJRwBuAIwrkKLfV
as96jwU/9DbZoYxr57ddZDGTpyx6Pf81iDIQWTvuwOHY69RwK8HwIwc5XLGdwo+XBR2BFhO1KPKB
GCILbSEXcK4yRLbOjpSBX+GjNW//V82Y81amyFtLaDJCD/j8+PrQ7Bz7+fqBr4MkoToLCz7HuGEr
Bp3jpuXpUKlyjiA/A7pAcAw/hCY5PSLCdSjDBNqilgIZ7crTT1AgK6Az5mUMNnaLD9VPVhA0yI6i
fuSuz6iHWIW1oFEVGzWkyIXaiAwqZNx+PlvqoQUoziDxFKgRh70qLc60BpDKNHMzN5b3QU3R6Tr4
7ksyPkt77kGNsOxhisxQsO37SEgHC9zHs2/8nS1hvxW8B63onv0qVHdpbpyptfurpcw6STT3pg8F
zbA6NzFFlvCqNydgpVVSleIcyWvI3C+DLCl4wcsbC4g/pOuC/eVVJ0p4qY80uJniDeTkdhXwEHYn
b1XCDDU5d4lQxT5j1aNr21I5+YsFGomw7JJ520t+VSo8eHdnNsVzLRg4WftwUb2nkYtyHdDM3RAV
rE7ZhaOAzQ61Gxm7ynSrF+/u1xRPthJsb5Kjl3VO00ZxWK+6ydJXTNY91ZctHrLlWroVyA7AhCb8
/P+mLRq8WIkvxL6fpUlTyemt7m1Z5z/vM1XH/CbPGJr+MrkwEhLb4E10gW+Q+6kcM77u1cBEPXUQ
7C3Cn1fVWpAGqjlMXo7J5vu8ZW8Ah29BFJeUa2/U0infIgVHYbdV9TH7YQ+tPfBvR+EeTR12vJEY
S3CaONVPKEy5hLfF5MHRFRFcjArVEMz8gnbw/8Z0sJX7qm5om7eQZt1qwwuDfwcAxBghGggalKYs
FvUUEBY81X8gZ8CHDfO2IUPwX5nhf1OYHq/OxYxHi7Vm9YBoL2/jgobvIVAGQvZqwu1WxSPAAVKI
tFAH0uzco6DtvOk8xSDmi58k1Mvj5SkJ9I4Q9uXwOtk1Anv3r+ft5IJe7V4ZLqxHrqdgBxBnHNTx
UOr5Hn3MbT/y2wXtyVuYpu2qhrZe8uzDaXgdMj39gNGv01D+gkDgp6+s7tnh/Gn7l6I7Wtubgtks
eN517DwnQA4m+iitwoX8rlzKxQoUlvtJAg/cfJwV1DPBVPwp/vheF7ygHpLrgVa5Y8MgBS/bh2jh
eD6PDVYro9s8P/KirfVmiYqVxeAwr+nTi5DdbZgXT9Pyr9+SgWtkUQk5Vy1OagtjyuQlceuTqCPm
KudBKhkaQ2gBUR1FUjo8cW+T//r41+XgVZfHpnvVASJXff5dL9xBLcI7EstLOB59F5A29XeVi4tN
QAAoNstu4znX001lcaQkX8HBfsPjjjJVc5zPvJ5BkJSwA/2BaN9W3gGMzUDLEU/X22T/3HWJzDPA
/L2QVaFZrqRjrXxso22/+pKFb3wH/EYF8TbtPTlGF21EdgJzvv1I/uTRwQjQ7hALJ9dH3WjBo52G
EPqzjWkpP5Lqcuxx6FovmB2vOnOkKoBPGwgmBjPmTprlkeIikUpL6TI4O505z9VeOXQHsQ/PL+b3
IqAJf+6AT6gWX/B5DZ+wpN5SCcqGaj96VMoXfXlGUjpevQL3DNcKHUnUx80fBQIaM9+AsHjZt2Vu
REGfjBCXTZ9eDBr0FqtkJutV+cwaF/6KB43laazP/D/c+lBZ0DwFLq2lWf1iZyywrcSsif75cv6Y
u8prGWP+VwbN+5uH8/w5Oboa/eM9UtBz4M5OdJwTxqRDuReEtA5m8f8tPAZEQ6ajpAM9NNQjAXw7
Lu0Lvo8YAUoQPtd6oNRsakrGViy5RfDHVTfqWFu+HKBVBvIPqAzDr5X3sXSVNNtvB8JMPytI8MLV
Cb7VQK1hjGX/DIBVJMYDXSmbA8Y0Cpd27ezlblIu7X+uN4Duk9YEy6DU/RB1LIEtrP8nmruzLu8U
y9Mnpvow8fLZVaAX8gRx66X5q/k6gzDbxPCx1HWKcy7kYrN+lig7VKHwCKHy90+lchskNnXK85/U
+0r1DgoGD0E2o+ertPLwR0VJJ/8HyaTerLkivyQxAUaaDBymmFHPAJ6Chr44YmPJUs7NVeT5IOFM
nwtqTsB2L+W9JboFcac+XBVOeD+VYAO5NvV3ZfF3O4Vx050pECNDJeSlnfCuvIXIXozBkXzkLIdT
o6ws2IXulq8aYr3KjVlQBGOs4cwQIR4icIvbE7Grwr2SC/J3EldXKVzhv4a7qWdT2fMEuwMKlCT6
9c4hrBhJRQi+ndCh3w27ZmE/HPi+oK5UuRm9X/Kz9bhEatW+PLVYFo773w20moZmeuXqELwbhyiW
dWyxQ2F8hIw1Tp3piJxmUxuosiYnIvWP7AJhue4USzAQ2n6wt3YMHEh9GHqz09UasdQKQchiWNC+
yGxvmZo5kEWrXMFq0YqGV82+wI6i4JD+d8bpWvxvzf4T+hScR+EwWWuHuqB/golaYgtHoBpZubaq
57aDYtEDwLEMhzGqMxXMK6O4v8n/6LPogZRDy4nYZobL1VQoxJCkvJpbboULvcmm5lVkSjb50OBG
V5+5tViEGlma+EHh3KbsMjznhLyFRXdkEUux6w+loEC+K8pNJXmDpNpm7KkrzAlLeTv6L2PQdsJn
r0nFUHait7CCiRiESjp3jxni2wP57AyCjiCY4ERiHdqFmdnvulyL7tRg2wH0jhL2Y6WzIR9IG7lT
BFV/Ka3NZzzTGhFD240P+24Y+/gaWYqJf76qVqVLm0FevK1qwPDIRHhM+zb1kTQrHV9VeM5Yzl2j
xdJIy9FckGLzoxDPlaCCR89QOlFV9aJIvYTfjWKaLMooIH/V429V6ZePCLUgPA9N912w8YjrCtD+
/i60kfpy7Lh6a91G2MVxAqdyR8B/vfhfc3uBK8XAwWdRLZpo8V4pfY73NAtOYU1YKisgMOpS1tS1
FPIejsQs9xI9udx8U5x5Tz3LyzZHOss0dP7ej58UFpJ7ARuwaMyi4awN31kFRVwpW4tIMixTT6zi
Bl6/BMoOQ9RvXjxcLTpRq7ZDziIjDAAksFxLdsIw2Jnf7RvLqhQ3mMhX8wRZBB1IXgmN53NPzjgl
0c0VrcHFcXwtrTFjAQLKDKEZ5wg6zEfmiA3sqS9JuMe4pApjUb6S6OakmZaFjpnIe3D0cpKybgWc
pHN5q03udswmU6Q56VrSEhWJZR4/Py+KJhtL25HOGnTvMiGLgyJdu+pRbV0nA2zb8jgYLMItghKu
QSwE7ntFScTuDqag5eKymrxaBxqZlJI3yyieT8JMIpKL6JOcAS7dj2tJFAgJL657m6CALel6wzoN
mREXugJQXwp0t4ww6S7Huem9L+7rqF8gOsuHzvQMYcSW2kWZylEe3nfkbZcc3MK150tAOuLh/azj
MpFTNyn+C3qM+6gdQk3jPgECkBZeSljcjpr70hEWNK8/DQwym1yErebEb5SAuz0huOui3TEblluF
WmYJb8qEyBiQIC04dWbzT2ZXicQJWEGfjxqCqzAEu2eOF0VoG1+sDxmJll+ylhh2aYbZ8eGZdz6Z
JYcHnDiGDAV8jUuYczlaydEv97ol8QMu59I/yB++b2uEYYQ7SNEhNXPr1qWYAQmAikv2LYAtRaJG
S/TtpSSskFNzklYpLwqXDEqCuqkZYeso6P6tmo5J4wlgL2hVcyQ/HpSA+JX+0v3H1qpOErFXsd1J
7PE29+P9Gxlwzzn0RW9GfBeE7aO0xILjToVEoCo4LDadhIPatMK84/93k52ABihRedqY5Dy/HcJE
1ZYuJT/7WMfJKEHSAPGBZIYtDWaNYZ2stCZZmBlYh7Ob3T1xW9XpicZG+rJaQpJV22oBFB+b5U53
2YAebznULgKLj4sygvzQF/tfBAUOnkIV/GxAtLT0PCsTooAZEO3s9ILVsrVJMR6d9W2qsqmr2IKx
zAJMDtojVhUZVtAjl4mY5KiNB9htDr8Ez4tAWJ3qqbA2TQ542f03JKjyOMsHPn0/n26wDqE7iFXE
yLMJB6UKM49qDOmHS/CBf1uJDrhDPKszbFe7h8ZfNK1iuYeQ6hmkpQO9k8j4NDeeG7yPWBHENvnG
TT7Jj7kpAKAhBb4d0pdsallaCVA4mNJYlLOjDzCOUtTQf548Hh3qDSz41HuAabnjZs04t0aK6L48
8F9hX5Jmfy1oriG54TPmILjMP22xVI1woDsrUI7Uk8odMUqS0r8oO5roFpuBRI1Ob+z/7u2+pi1O
MhOTQzuvdKIMi5qzO0xD4yYlZh+N/3AuUm60L3A+5O7PHGViUBIKQrlERfSvlJmfl2v18AeSW4mu
bBvGgcGZEgAgJ554b4msFNGASHit+N7KwkkKMuCnI0zUsnZZ6YRHRKTXSU/CkSAG2QslZ6Gpysgh
Tqhfgx46lDy5CnciAa5wvAAOiG56yY8oui2kOuCabjATYzUECPD5RzUiFaL7ZZQHlCqzYcSqgHr7
JV1yCOMz4GgAJe9J2LDVuAvbZDUJvcDe6MCfikolSTP0KuOoYFcz8Jb263yfM0EYdjKukLfoV0z6
IF42BwiY2nGyjdH7apJtEZ6+xeW2QUkWoMrcusgh7bc46uahJ5okHjEQZYYwa9PT4+bJ2/BWK2fP
FnYLAOC5/oQcrUIjnpmCzSumF8ImsifC31pBoXMTiN+YoPJWmRJdvQUDFQSp7TyMqk5itAY5VpAa
hw1RKNDgBkUzIkXJzoA1Af7+qu9VYO4ClpCRTpHGhK4fSPjEiZ4JcDgb/0FjpLf64vte6h7lx3MN
BgNbQQcGz2z5jLOpfOnNKe6SMO0+MhgeLExfZjFORpt7JB8uG4APOUf000nRqySXeM//YkCfDJDO
gDs28JFuOAqMTxqyXt94VyWbK9pybx11gDHk9Pr0UvVcPrjnOVkpsL9ZLUvaRvv/uHvhd9gQhcd7
/2Q4PMU5GFQ01nNZglZuxjjPKw+8Kt4tMpmZ5JugyyHkZVgSP36M8yzxSNJ18MBtC086C2pR+r/A
8ir6Ltvr/2WkyC8g+M4Qv5Em2SncjpWDnkEC8I5BQZxMxDKR+ch3QqnDxaMB4DS1AgpgWzpHRkU0
Bmh4nHnknhYNXV+HMa1QRhS2qXHZre1IDKFQ51vDIawZdBSthId8OYk+PbH9AhLj+KdTGS8PAgDm
FRB/3+oxakgtcnEdtnSM8feXmvVXL0IWFWOZlANISVAj6/GblbsNZx2YR3v98V6Ca+Mo3G66QM9X
aYaJyBHXoyvuGRN0sHSWPs3VRAIZoCuNJeiC4rh6qRJJY/WBoNl8Vi6OFLayTc/19m67WrnbRhJY
0HKAsbsvoUBssBFOIsLybW3fMZLeqoJ/vivo//74Shym5g9GRJY0NXYkuyW5k865GZvAAv2brX9P
36/IOPEmkhnPg+tHDjUKXgae9qDc0Jppn3xSDLozW0xrD9GyUY4R7jO6fiqKC+Rd/cKeF2FwKcmv
1yVIYNiqzFhxcxR+GOjvdFo6AdWvlTZUbRkl1xjrl4ZVePVPlgJdXChz54KUW4u4Ow3a9LrnbLtk
n4HCe3EYUTSgzBahLnt/tr2KojHc7pA9r06iZgesi+GgHlyhYetxteFf1zWgb/EskRZdgfFg15En
mU3L8p/u5VADQfGVAV+BCq7DyqXzNilLStlJL98o6LHii5JXrvj5/dNit9ltG0W8ZdRkUV1Lzu1o
3xjZfWx1mkohmAvSFYiw2NTf6DBSKPTJw8aUzxoEGBXViQ+RE3ypJm4yMZmrIsXINNk3xjZGUwUo
RNUYtr03FFzn+o3y+8iuHG5J74xcJU0ToGK854YJzaMz+/IBJtkd0CqnWHjpcFiAuzAgbRi2aQFf
52K+M2hQhJLQB8+XcbMrznCKEtNTdM94OKnB6CZSXd5bWNNGt6xIqLa+mtNLvtlzinCDYMtiRYF+
edz2kwzt/fBy1lh1f7w9nEUTR7lFR1HDgh+0V7vfXJOlC5VtZl9dYH0K3q2QO5fqDnpt+0s6Nwk7
6AmlOge6PM6Jt/RH3eEKDzYCAvxMn+lIz2ms8+Dz+7edE/WvLlSAgdV+I+Vh1mXJcOxSeLbaTcGj
F10rJH80LRIqsifFGOAX0k/dObidNItbEz9xgA2s6OPkUXYwgsA1jkwOPQjt4IcY9BIw3atEWEZa
ogJF2ujjtzU5obcuPylTI3Ui1X6bqHBq/R8eDd9Lfb0tpZeXAecn2j8xN9d8CLJ64abxQ2emeUkG
Zfp3JS7iPJqZajOsg2LspBWgwnh1FagzxPJ/nR22esl/NNwwz1sZAZLbQiz2Wr5rRjN+ZEvqZkbO
h6CgyAR+iYxOsSl/0j54x/gs+gkMZAD2o5YwMo/XIlcS/1vamtIwtCsl1MaVUc5V8w2Npz+ixAxO
kjA+VrU68Wui6xKrQ4CGADvxbnyxia1FwNDkJROIROVCzkJ1wiOBzh/lIBmMu00Xtt/ceDn7orhZ
LeJRFWcDaAugh0ab6MvllyyYQLCT1dSgtsH8FC5FPk8ruxdGmVp7UnFXGc5LWfy87z+mAg9ddSOS
U6vPuykIR3cftYyeG9lBAaLiPLIgI2uvuUvpYsIQeD9gSY7J8hKrKlHmpueo7yB5EB1CHTk9Y/bR
ZMU9GzbhVZzriuXny3GW5W2ISuxINB++sQM12eQ9PTIhjlFI023bdC17e2Z6OUhiI0svmsYd38gX
VlAOB0qwtyIVODnNjH2OA193PHjDhX50ic3TInB7+CrJ79fQWJqPu+SA4rQMwz8GKK2Ko/ZkeMyO
NcLCGz0qdhajRtR7zBuO30KnbF1RiJiiIA8fTZty8X/beJLZm/jLbQ5krP2SBr9WJ5E0y27q9lc6
ZQdgx/yDSju1A3dm47lXVnA+wonuC69kL1Yi2Hm8Vq919tpqW7yW1IZNw2sFK2ep/ZAdYp+3G/N+
CoEVqft6jzL0OyOLaa3wivri5QqjRKBy/oUXaEO/n3WjSitObx3M/fiJXoGq3WMz71mCIgutMcNe
ctDzMVE/WtkkTYI2dWabljFt/Xw1/pfwscjGLE4A0jPMMX8Beri148ia5EKH184aB6WvSnbNLciH
+vJpx+CElD9qwrxnqaYSvgBtBln7j9W0cvwy22EJnFV4e0p0oEM7TBdPMxamKA5hdpWwQJnxbMLS
50mix2sd8+BBJQfn7Bb0AU6IcRxjbiMNlEQ67R3WR9aiBBYfgBZCIyg57/YLrPWwTVfguXvj0exK
cE2xGuREAPdQXvoWu0Yizh9Nh0gCrPH+aT9feQeVbgBi8vqqgAgFdBWDmtPHST6ejDDCi1Zpak5h
Ca0UZY/KVJ9eMAio6UfWwxyhsGv4Wk0603r5LSwxqOXzfVCzELFeIsVobFKrTXPOT8SeiEQ3T1tC
iBOTKwnhwUbc381uNabt85njyo34buAS0QT+VDXUZUoJsxzZzJlURqnAhCHaAki5SdJSIKzpWB32
Kp0ymJjGSOKTZJNw5bcKt05UOu6EvtQsiEIeMQqIp5HYjrqba8cGmnXR+qWGgFvL8mj8IcOWx2vW
JN1mLd+UAfZwkZgP5O69bUoh6pEA8ttM5NXJv4YxtjitWBhaad/bkMs2MMzoQFNQ/O2ti2qelKZX
m6fe/V83UEwhGBq5iQ07oaXhvIPlFmGqpKbzIEdJ0x7PRPwMTEvbKXjWQ963F+t54iqdXfhAkBsW
b/Hrtq2hE52qrgN7e5wUklwYDc7oWVP+IOEltZg/I6g1M9Qi2QTCxxPl+9ozBoVll3TAs5yie5R5
awuEfv+wiyrPdmoORjudnf5EIvXKdoKZ6gRHP7Iz2YS+Ddv4WBao1lsdBYkv4nWi2NXoBRc1ZWpn
RrncqNSDvhjz8k3K80Ln3oRayWFJw98zIkrR7H+4G7OAk+tr1hklxOqxFok1ztX6L8Mo7oywbLNq
Ek9Y7NBKKXsME9MfS0dgeUilgOGK6EuvGR5MN9Af8igoZPLrB9hWj0YZPBzqdcttQr0Q0W93SI0C
wiaml5fjYwYQZY3G/XD8xpTNMApF8Kurp6hJux0bcrIwhKtL5tmvd27e9knLsjHO4TMruD69oDFg
WNE3jg1yyPU3UacJG+c5PLOo5Vpg57/XzXrt9sphx9iq7gBmE4zFeer/H69vAo9ibdScHvNY9RXu
8eTFgNfGbIlk4AJolMTr/YHTfrgrBqyIibngtnUpsk9n8nc2LjCJY3PHl1GfYp1w2Q0CaxqxcWLs
ZYKoqX+J2fo7VFJJjB9TC3+ka2lJvktbVC7DyQTJDRt1YmcMjVeOfqt4m6B8DkSoe00IMPZRZbmL
K7elbPw7SMkYIoyAz8Qr85QDyC9KV7H4WhRh1L7XVA5jy2pPVxKxNoEj3xfZztdo9SXZ+ZH7ppS8
eq2rzAhsODAdDZ8BLB2HsMItBuKnwOOMFE9E79Nfh2XHqzDoMrdF3Nzw7XiZudeQo8xCfvYFWtIN
9USz2QFVOgaDJQ6fjAyGT8BVRVQfxROKYMICmU7rtzu+CG73rFjIkFP3JzWp369QSFhQI3LigueI
hpnB+IeY1Ym2foaKgYPyjFJTttf6QxzcaYBMLEzdWQpZ1a9NVzX+Hf0udGik11ILaYC11DyNJmA7
XYJNCvh94HBcP2e8zJc1blDNHP70eQ3k8+ulagRgbccFfdM5OyBAWdWC2N+RxYRoAzwIyiFrWTnP
/TSrOl2NPUqGlWI0jHL1qczp8kmYo8+desvOpd7ZRLW3IoSfVScymgDTz5cb26FQOpggu+RfAKkH
bwDEdRzPNpdHsYUsnBH9leIithSutQM2T02YXUqdnxMzL6OGLNO4TJvWgjshZMDXTrFqz9QODHDf
cgmQT2EzK0rMTiWWh3zn5fC8aKpNjCdiN1/raPOy0SBEhhiz0gjGeVpBW01bIkBUoYyUCt/iCrMC
pxFVS95VW/JtZ4Ia4BHBpvUWEnmfHneQHExjUIhui0PRM70OuGAUOilWOBAx1rX/bB+QaXL8IXGO
7nf/1Z7N/tneQ735gfU0ogueYeIyc7Sc3WlSRaMn0x8L55/UubxKaxYM9XGurMKbVukVrrDdQsbq
2PwsOam4CqRNKHFQ3UA95mspC6dQIImxJN968+SrX6H26g9QIq6gGO0qx7y0T8b0x0lBH3Est1PK
WU1DP63p+rdvl15yiQu+b4SYM9jLgZNx2788/UYaBAmLsiEIatLOago5Jp8tQxg9jLiY9D2v86Ws
YtJ5NFtwAy4nEQ8En+eKNHsXz4nPgDCiklTvNKk3abVrdJ3dCAqnsqkwreSXTWPiCMPohQUBIDWY
qoOR3dKEm/I4ioNl/P4ZW+Oy/VJf3Yeg6JDuOXizfjewVInDY99Z3BsFUEtsg37JwfwitkO1df5V
+0SSD5TXzcJRPnjd96LIC25/KyGs9KmvSArZTYMYm7/PV+cYboe/ph9uqDk5MNeUiloKJnJMARBO
4+4r4PnRtxm+c0xve+mQl1AJbQAFxaNplLZLjY/glXNQiEVWp6ynVGIyvR1stn/xAViaZjaBKrDo
YQI04R0DAMEQipOhqfH9ppIXtRu7mqx1qpK36U2FJtu3s0jww3YGOEpoqNJ9SCg+RyWv03skmGcc
LOcdbdpYzCQz4I+CVczl4Gy5m9UHbF5nXmrgInuYBE/xzpqbk6emL/QXYl0NZRFfNHyvapnf02Lq
+CDyMQdNfnqVwPWdIz5HjBxY8V19y8eVOVw38IzV5Uc9H4PNxQD1+0Lo8zhLH0W+rFRBwHxnrXfe
Se2fl9jhHMlnSBLNTrNcfktJdKgWPZ7o3x58BKcIoaoWoXWhsD/f6+NlJHy8OvchQ+vV6ErdYO8D
GTHXrfc6Xv84v5Kh8EZEqA+NntoVYfU/R3uHRcO6oSS5bn5HMtU5dGUn0Jf4iJaom2+TDmxSNfFu
sqOkOvkdHkwS60mOvsGwRd+izl5bBH67hoWm4voXOKNswsY9qv7tyk87hdVtz9eVRrux6er6ztE2
1XSrSSvc3LgPsa4FieHd4+kaYm1XMaX5CWxRfO97m0yWb24lFurDhSn+8n9m7a3MSbp0+TNiPaGK
EKDcjX0mNbctQi2I4FRHbknPrzD1RO92hF5pweuKM1v1BexTpVASyaT/lNL2v1zcr6L+NyWizqLY
UargktXomTlczAHvgMuEeAn8QDInPt18WR2q1HMUhjCFk0/IvuzfDkZSJDO+Try3n3/sGx4f8iU7
P56hSRs+vNVRMAVPmNpu+HTRo5l96DcShkTbmj1BlYSvg+ggpGKold3DF9a+A1xVNwT5mT9hV76s
8y5DNMg4PPrrEKnaFg4RDKVIkpJE8SCUWCp71d+Oj1KWXJaxPLxuXTYOWchveNGvrd1h5flIWOqk
4L+jQMeulJGT/Jl+Ax+KOlZwRKUdRUGgVnX84/VC5o8BM9yOIa7445drFE5M8s6bwbmDob0y6Zxc
pxtHA/6ur7fzIkfv8+E32XHz0+6p2knYTyN43ATOp4F8SdmKoRuxagS+90eV4mz6/w2D2E4NOCsm
P7DHrvuMHaIjZiWkpIsqtEHhkgrVc2rAxyXJ4rqDXTDdVEtMDeqKraMfG0tCBajIsvU7O/AIu4Rk
MhaFrtwy7z9qhcztZBTmxgZ84SbvaAbe4r4m5fPykz4IC1j+MJAVabInVtdKUWgHyaiO8n96hkQJ
6sM5Z7bPqrVfc65N8hGoyxkt7RWuNlnVfKLDoItNyUlatAor8vcjoV8PcuYG47Wu3/kydqDOs34l
2REuF0P/vt1YJZcOPfpFlHejhZ6+mUx93pP2jifrgL7/Xy0TPAN0fH/6kI5DW+1248+ygKo2m0fO
6DNOmdwaM7mBj+AxjH9Eyb0gy7w6vCC0DxYagkdS2SpHTR1QayMHfJdR+1mRaHK4CPOBqGcCpaB/
RxfsvvLhoJH1WViEqVu3LmAnU0+0saui5t1jpcfhDcmqsuigvqYNJkMSQuEYDCmCLU0cJKnWFyyl
cyqbd79EzRKqAj2HeloGjWurpccPmtlAEFWg5YRtofI0fAoEIdsLsC6gyE87hf7xC/KZX5eR1Lf7
lGgiJD6RNWi/KoBwsBFTggDeGVWtqv7zxsBEQ7N9WUa5WD7Ja2pzzpVX0j/W/WH7vwfHF5m7p/o/
9tMKJFxST/aS9OZ/joZRfTKjYRWfYVDV707RVcwrFY6TrLx5ygL2JH0evMg0EIUINzBS0jOR0JMl
O+DESoOydkcPLfGO+MuaOVaiDQNigdYF0h3KWn4DrKdh6AeZVTAmOPdbOt0I+XBVPN6CqCi4Oi4f
Y7YMj25AKQvIu0zhox2wMwg4X0yL8Qj8+G69Zbgvzuso8///blXX84sKrqToDkNce7XGYERXRUK+
/EpsfS/8jztjX1zOAcR2TseHKDG8uiTo5mwPnGxEAVCWj5w1JQEeD6D09SPADVoJPWYth7xq4sP4
YPYeyT1mUjjSw0cMOJol2PwdfBjBiMw7NnTXrMWwM/9ad/JjZt7ACqy+LUWKj+dbFzNRnnwbPBlP
KMetxJbZO0QC4ZV98/QyqdJc41REiyeGjeztWSJVmNMrmtY34quLl3oCGHDeLmCn/esBHOrQpZew
8bj+9zL6wNHkbh3g+dR3RoYCxudvxfuKnLjWzyN28qR0mUKOPJflvdOLP4rAij4jQgTu3jS1hDiG
ufoeZV40zcuviuTaldRaxN3GJ53jDAtxaKeYQgDgw+P2W+2UqbE41CHYALSUdKS9ZrPkjr3ObNx8
0TUnI3ngOwjS9bjYAkMGR+WdkzgzW2OdXWYJqWDVqou8UJj8ep7EPHqILzeecS8xKmFT8Vc1v93V
rVLCj/DhIyl6bIwdp1oMJzS0zAKxCQuE8wndbSF8MY/ahtEaHTJhwdFULSlK0/3aVB2JzgADr3F4
eMCgDyw3HwOh2HnGdSDBHgIn3Tg7D0CsNe+q9aGVeIqOuhqI6jOJzVYXtS37aLg2aCRemzBdF1Ay
lv21W1avfqNtOIUwqnautBZzCmfEl7zASHRZ0IhjIzyjRRFaicfrOaAHuJMhErs3HmwCyYL3dQOQ
TMaE5wTJCD55K7ircuMp+wpofXk8M2hQdJV4adgVtoODxPSlhJz6nC4UiS+xKhWxUPkwgVmp4s5h
HrUSxYBfy0sJjwMrHAiXA56W/ca4OKMThQRvDW9ssIBYv2Lz2yGNisKrVtGU+uJ7uH8qlQvtOlgw
SovR6ZkfQva0b3u0mkODfSTqJDqjqHs16fJB3d87/l8Ew3fM2A7ZiG/ZyI/Z9aOV4jnLwfg3Dbhh
a96Bw9m0+i7ry9wJD8mO0dATLI1HP0B1VMbPO6hf2UoZt+d2yJWk7kKF+EqxGHGhgkCH7eSpAzOv
IaQW6jq3KnUbFjD4Fsb1vbReI/rafilVusvaAGsv+QMxw4OA+n8zwJz2qkF6W20sqgL3yot/4ASh
wOK9GsLeURcKTTwjqioxy5Txhfn1x93hTcZ+DbiVRXfwiU8GC/34KsJVcgSuyEeEhVC0k5exS6Pm
QM/+Ne6XwGDFXQA/E9qfSo9xb7iUUaxZBccrNiAlIdHSwAJFfsRHNKIVgxZFAMF+oX1XjtjY5/tf
fHXjEP1kL6TkzVOjHyUDUv2xrux8oLrJAQJPfccYlJUe01S1hyF5Ha9dRPkfQlKnLt6tpAOTgCUc
fehtd5UOfMX0ci5hYW39ncb0Uh1jdx+AHVbaOA+ChkaymH1G/Pc21JFHDx2/aNeR7GP7LFT+Dj6t
Uycj0Hn0OkB8pmO3H2SLZkkAY95WQZbGnMKfrHMFgdZU2X0TjGQyFo71Ja0IIpDiBBv8ZAoNfsQl
Y0l6qluw4+xZrLIFmeY3E3WiZWOG4hAi5MbQ7xUu7yTxK25W8AckaKpn6Kg02IMTUmT8qcvtobim
pKBkT0DMaGsa/KCzGh/9erJJYzsDEg4o/+djQt+MdGz+EpQY1HzSPg4voq6yksJtCzwQ2W/q0ZfX
oSzU/53xBBy89Qs1KpGJENEvRJ/u8LwbG0ji5fsN3b++nPRy59M3LziAP2gKNVPOejsykkEDjhqn
+nLLOJTWM7Vnea+d84KRvRbKoRe5qmq62dg5UDlFovii8VaLOuzpX3ba3k6nhKfl0UbrIyCfYiR9
2SQgpa9ln1SjCSSm3BSX1zgC528SZFNUmO2RVImaKlXKEQz76t9YHC4ILb8zCOGh2+KzNi7D6DR+
/W4DEwp4tRFCVS3BzOlIbXZe6cOKi9ofrwIf+GGcciMu2R8gOO0qVoOk1v9CJaATBy6xlCIzh4yH
fqHoxWqY+Ak0xetiJqzSEiFyM+/mYLsyiv0VZIxCaqbksB3i1Z0POkVESpUEXz0YopGP3oDE7LRN
gE2g2kZFxyb2QaiZWiIdiOrlQjFXvG+wphAHg0/xU9lyV+3OcACHPXvPm0VYK730wqxyFK5hTig7
ZVp1sjzY8H+zAxTUol+5wqfod/RYvbCaMgS1hjwjRrXKGUUAAlHS7RVx7zSATE5f7rnR7hMvGA0w
frBLLdp3YtcdZFDheLn0HQ755RfaE6ozR/vfBXQ5OPy8uvyEyyJpvgpL+yv6zUR/dQ92U/Nvt6rb
b2XC9u4cGnB3aYRYO4j/qyj8smZo6odP+wow1kD4aYtYmmWR7Jrajtq4+ehcSu7i1d1tklKbppvH
K7rzFDMztdWrBzvnMvG01kT1rRBypUD6Flq5yc7GZInSEz+jfNmb/jbQFcLehSRF84TXaJkWZdBv
dEvfynpekmQm+vPCEDIFUrZHbThHg2IWETgoFOhqpEt6cyheBZDBOPQ+QvUce7vMMOD1k/F30gkc
ZhwXia6rkwSnOA+90tXsRy6F6asayOtTyfXc5e1M0kr4d13HBUjDVNebV2y+q3kEsvKqgsNDh/52
6S0c99zM21pMjuJkGXYkRGEIMQNkpo7Mp6GVfsBb12SRR/i5KX83Zdct5CodYK6KCnS9bQqkYybj
tz6kxO1PVYlfhskDS6+FZjq3Z31rs1S1D1kB2IAeeLu59/Y2z1cVw1GDRywi2XU9zPEy1/n0eLc0
w2R4FiGb+cBdGVSyfo7x+qiQGO9zjyRo4YMG7dDShdqIZpybwFtgoFyt5+o70GyS0XF40cp8DVpq
pwtZHQpk1YoHRIaSL9AIFyzKWjCluME/odg2ZVHsiMj73Jr/E2iY5mN12aX8oxZNK+sGL404BG1u
lmvUqHP182GyZZm5DMXgjSjytNHRPnbodJjtfV6S5bM+EZSLpx2h238QY6l8GoSITSbYplmN/z6j
onSN6vsSfa56nPK5vwrZ83NcaaF7o5+xYHt5V+zllUX151oolFHPew6Kn3N7mhvdkLx6PpkcYuMt
AkQxSseoQasB34Jw5u5LfYd2C997umMiNIn2tlXuDrfsaQyeCyh0f116Btoxb5VnL9wfSS4BhLwj
dLNJVUeRhAZK4C+1KluTGtLAvR0R4d9XA+vd5Aq2zGp6isJm3rmhpaBmk/xoiokVpC9aZz0TVqdZ
yDf8hIBWdIc5SRhoTEZXSdkYAFIM3IhJBBIeGus6hWZaYp7GR9xXIeMgNv+avsPgqu9TTxcNTjbE
R5/EXISUhaQUJmuEhgDvzKIO6xE6EGr3L/Si0+gKC86r9MV+bUVzxUzo3NLmYJIJGA6Ec6vNeqCo
2zrLPMz9ZT/q1KgwBRbGSodh/tEOguMbvvNsFzi4aBmra+IlodtRtpH9wNJ+eL4lCjeSbEDLaNra
t7mzJlo06YP7KviQT7su9wgsJgzO45Qud2aT4nn31OWSl/MTI++cvrpdEZwzI32yBdrz1HT5TbtQ
YTmSIL+Yreu1A84zvu6mBd6U8j5yCNWy3qBMqH11j5SJeDZx8Qtar06OfF+q5vM59YU5gO2yzl3z
GNR3G0/RmzSMJBu2CRRRl4sSvKv+2C6VAyKLZyyeY7QZqTLT4GXdd+F71z3I40kkDofZVpGqI//k
eQakdUsBxjI3zbJXtJG6fucubBqjTsy9HM780b6gJy3vgKijRJY5A2PB2+zpAhO7wxRFneIGn7KZ
YVX5qpwIXlf2MEFjJWg2GKFzaAUYCapRBYK/Zr5msr9BTQzkJ23NBP2KgtAYgF1znqUoA4tSagjd
JfVHplK6k/VAr3lx+S40GdHmmjafUNtvaAlQIpUg61Q8dra1RzyspgF2avrkk+v4g7YsxA7sHzID
HM6imzxJOsYGRyZHDqDVMn3MoJpow3gThZzqfesN4F0KbcjMuqFMPyuwuuPoD/8uS9jQwJHEgI5z
BSlbeeI6TLXqzhztR5sjuSzP+8bJ5bKgQZljumsrxGBp5MYAeB+f56YruAtCWUsSSjaLkte0Vvzx
qQBNqyExo++kS/pucF9uJdwGSYVHXxpZV11uVjAxQ1LK1p/L0bVejimwYNI93YmJIeys67OXTM1Q
aFUUf9zprrr+3VxkYEovdi0fRzxRs0Qod6xpZdDa7usgJCKE3/Jq9Pn4Dt5VjhfNCW9ncmIEVTx+
+bjXtbh5KLOcitMgqt8/M8Bc42D8RngfExKWBMBKvYbWdGoRYq1AcxAURmRS/eozwjvZeELjDt7n
LzqoBtqnWFtRJ/pY0cNsc4EvuN9ZGGLMd9emMEw55fKBLrKElwx6tqOZcgQANktNYPx7Y0NCqXte
aFjcDNpQJ05WL5r54ZKWI/5ENJQ40ec9R81ROtnQrjRs7GfqG4c1L9meXC2U4DXq1Ff4dMpINL+C
KCsXB/qnpIGU9ggtIGlH1FP6zbO1c1kDAKfHNR78aEx09Dbdd2CnwZjkGTqhfWNWt8+izb4TC0eG
uULDHt04DU9VG/A8LxZwQ93CjEZobNgv53XT4gLIAMsdicKjkE/yWkKJGxWm6l0D+BQ8UPngDEve
+41ARrLg5ZNMithfqMi9G3PFMacSXDLcVY9ddbwx/UvfE5lbJNZl6sxWDIyYhSnKKbkn/+1GCgpy
hhSMAfS00y2Ue7r2zypUPWF53Xef1EzG4gCoH97xcB2SDw/Oj5wVBJKmfhQzbX27sAb7G1UrPxOb
oCz+8dkBiTB7KC6ZyJv82JCBmbtSl6iO46wdYQ5FIH0C6hplYMo/oavVLtZBIwIMdj2DMRzcYqNG
lUGdOHCL0XBZJnYLYDLTpWmT3aNZIBp1vHiOnRzHb21CGBHk+KNzgDrLv6JDMjr3SpHFc4NaI6SB
nM0r3dNjxwWRjAmlXwSfCPBQ9F438KbDyjBxxiFtculyehNp89s1JzP+FHzPCvMn1hRgF2h/U0z1
8fL+/bFcYsynXwRz64gM1k3KEHc9KRszipRFW1YOlOPegaxejjKcAbYYXzOZCd7AbFlPvSCJNIr7
CfjeOCLEh7C249AgtqZT9IB3f8jjFqs74ItZyD+myXg+cSzk0mdwORc6Tv7mHS5aGfLDWAspc2Fr
1As12/5f8vBPK9O2ZRKdBN1iqZ6rjvGhW07j4VaHYgNNL/qavc6pR4S5fcUr3t1Ormjm1efdshzW
CanAhIXJfe8RXJheLZkR3Xr7hWuccN3tltOrbj+E6zlR+7taMthYSDANfeO5LzFQUY53aSjdKKr1
GDhRndLIKzflD+0pX0cmQ6f9E6lPmN3pI2F5E09BoalFdz96T9/Y61J7BkTOSaxwOKM/sIgNjxZ4
1yF+Z+206drDzbROmrDYJTtiSHJR7yEkTcfFixWy2BnwCxbqcEW+FpSvByckzUBowb9+E2cXjuQd
97bzqvPL2myr0P/q5W6e5g1+lzh2bYUkJ+7BCbSk7skoktR4zBnQtrej27w52fBiTbZV04TYZyup
nSuZTf9oUtrBu2RE/LrMwgMd+Q5jPPdHGWTjiUk7Lpcyy6gN1XFjRJ6OdrzKmRo/QgZ8iyDok7D/
27ifft6WioETGoMWsxyXHGWgjktbtJD9yZ2catLgr2UiVsQwfiE0KzEKcrb/xDKtBpETXI3Iiey/
Uh/IiQ605tIvsCbNestPfO3/jQMekvMMXCgl17op1tz9hJ+6Escpb2iYQkh2PecQzL+LU+VvfoGk
iWjbiuf2OO0930dyplvnqjUG+G7rjDhVn01d5lI+g2X6U4nxeW1K/JthDlM0TV3IaHY95HsUajb/
lIrSz/GXa14mP6ReewDDO1/3XYqF7gNraWJZRawjRGYggnIeINsCAB0bQf4TElrt7Tj8dU0H6z6j
1fM39tO3naqYcoMmTEVQ/jy4VcKtQqOPvVFvhrBLlg0sRcY+1Ntuqx3E31QJjsY9ftBxeMFOoVGN
ZIEEobotayodtV3vatLpegu4HDxaRPja5Ju+Qkyf/KFS6dHGHnxgnt3MlR/3UkXpyRlB7zEfCWNE
c4reyl6DD7Nv05qDuH07j+BfmNg3SlRNyKY9OFGPfVNOJWS+P9cKrsZj/Z6pJ+cRj5X/yW021/ol
bMT6z47QUM0QeU7JVU0n9FJ1WG9+y2KgnoLXn8Ipsvag5+t7B+uw5e0nJ1KhE0D2IcoEPz03oxAa
xPXpWcA5PXB7v/PYVj+NgXsOeH1lLSgDbw0uztV2O0UIsYSbMvlxly/nnJpSq0OVxDJaNOKPopJK
UYdYvbxo6KxCluPV+UF61mN3VbXooqXzg8RQIuq3iQ0nCeb7F6yYPRRjswsFPHcfrPGvJW9SJRoJ
s4jCM71w4zabTicNIJw3RQ0cDKL6De0X1spuyPfFYkf8G5HpqLKwzAfi1THUoqJbo2z4s6TagKen
ORn+zeuZ3JvG0AeXac3prlaOuCup2vx4avy2/VbunD9jHOQyVX1ZrHHAq4VQEISH2z54maQvmlHK
16u0QHqpeLIlAg8cUeRBpW7QR/P7NO3XGskj4CK9Oykr8YZkkO5hTgfTYuqaTF5pBjwWwKlp2rcX
iy/U5fkveSjHlqMGp216HxUoJKrmTnKR/WM1i1RKH9uUBR2ja1V5N8p/f0CsteuJkAehMeDMcSZ1
ET/1bOc4O41IWxG8qBAD0AjYYVnPrDAKWSioY4ZDQDXRQYA+ERVexxVblSng9+nAtDQyw3u6B+Z0
3n9GTO3i4gTLqgst2JCYM+pykFLrrvuWOxygZ2Hz6h6fy5Lb61lrNu53B49OHdNyI04YkszTGjy0
rF0he+D6E+OJyP8vYB7PR9NNJ5Q0qgTOWm1I5x+pQWSh0mSk2XU2S7N9wn5bTTl+rGj71XqTRc7P
8kOMdO9haoqlEY77VjI+EMn6QIjF+3LmB5mjmneDo4CidQzBQ5A5vStmF5+nVq0R0bZM47YpfDX2
04N5X45wZ76Ek1wPrQcuKTxRtFqHZLynAl9b0Irtx9u5eaquVvR+LUXZ9iomlSU7c/eE2J4eBFRI
ubRut+HtingjM8NWJDUbP35vbskxJFZDcL+kh+0lwWi6q0kqJlm/iA8JkOMFZJ/+7n+nDPvxbchV
zedH5AkMEDKDUeRyArW0b8Ep3OXD4TMYgF38m529g4MVSmNukA7Yd3x386DaPw7kvccEg3FnpnVp
o9nWBk5+zco0e0RMaQ/riGKU96JluUZmA1VyerA6fuIcC8ll5xmUM2F7bbvxu069QQEWqmUrtEvd
g9yd0Me51NEpNFneVGxQHAnNXsmz0V+Rm08RtTR/P1k3OJ3sT6kI2B+OZcZpyacBKlofhWJnAFO9
EPQVumqxIMjqy1nGM91F62uQTbZ1vX/X5b6h7euzag5e2osb73klJCgRp7fiXmSF5sU5/cYp1aki
X9s6YeODT3Gw1Z3mAJ9U+GRqfS4yr2xzfIzyVScpmgWcdwXD+s3vFiuMXucEm9FK2fmVCtFEFxh1
Jr8Kf7uLPiXFuRmdq374hxleQXmXaNCsFOWwm7rAt1C0s50ZBT8qfE5SO/ccAZFqPoz1mv1tf21J
yDola96jLw+A1eAZTt8fqr+XImMfSsPSzLU4eopRvlpnA96RiJk+p9CCleoQrh+GlctjyfM7QvuB
axZvWRvoHd2XO9WsEye/yCb+WJqhHq6GmmSq9VbwLCle8LpgP4Cr4X3/OE637txn9Hz5vX2yoiS3
GZgliAKOBfRLiQfEihSSetDrmdjPWe9eM0cmjJJEwVqC5V63OZOQE08KmmhYOQcvIO6cORSaPrlq
RwPUXFS1UOU9omNBPQ6picJE6PQArs7eVHH8gSE6+32gwKHU9VprN3TQtmf5V3mzLx92wkgvEOgu
Kg75IhhLFd5I5fZ/Pn6J0i6Wr5wmCC8vC34u2qzcjxtuEQuNK5k0I2UbdG0lZLAGmutDHFnhm1O3
wb+ODI06Y7LLLBrOQDPa23AP5Jo9Zp4ahc8AZy2VQw5aB1O4CO/jfqio3WIWWLmysxwcwhY9O/Yn
/ia3uYI9PXKWFjtm/j3HiQ+xtBIqO0mgZLTv29S5XoXD8n51n4sZigydVdvaieOtNqcsSQEWmAOT
ymAbIuBnLCpbJJMPDViXLeI4y6B40/NuKtu8ZaqY+y7UZYu8ScpGhlF6mzoHv8pmAeJBQPapWXKQ
HpyWOOY1uynGeAow3Lv5pdDFjlhocLTVSE8Zu3BjyGmL+wMA/f61VywtBjKLZIDSnKOYGCbQCb0R
LKmTUohIiYr/NhcjLmD0D1cR1S/V2NYWOXqHNX7kideaPtq3NtqXwFqNS6ZuZeQLWR0b09gIFVGj
m/7rQn3+V2FIt9+VlSE9zzxwJycmiKPkotlLfCNQ5EcmYlXaI0g/FXraySpSRsvRxSK9KomogdCZ
Sn8djr4rIau6D2qJkQy7n2dTXhiEM4ma72JPYgsAviSQBums+9iu69j7ZgL4Nsecj/XKGSN2jIXA
kIhYZ7OAZkX28LihSFPikwBgkUHBg+Yiv0n30Fb5T8nR9FyvhhLsJ5IcwaiNm9PqEbwtDlOZTipD
3x5ivSQyf/7C9tTbCfLQXHO8QW9Ji4Q9yYvY7R8Zd3z7KpQDgGbpdzoeIgB8bcKCQieZDzYHzLyZ
2k8idhqjcTPYMmMjLzxOXDj5WYIchwYHlpDaCAJSLDzSRu4cOUH8nZGuH2aAGNc514q9bZpnYCjG
pEHwXDlrBh+H5nojuTRcDTm/S51Ex1W1vF/F08sIM33lxGF2dJds8wXN5sK/X8GM8fpCN47Bak1G
WsLhNjHMDFqCIDB8TUB/sci54Q6lrmFyMYdF5rICzBrAEwweKl6eQDj72eLZ2jmFAgH24RbUxSJW
tYKViA7QdwlDTVx2X7NkRpk3RXk6GdEK2xfepe9z2E5uqbvNXIkwjvSm1102itnjNhgST2IURCLU
KykiLXZUsOkGBVT2MxKZlpTJWYN4WvCBi1SW0P7Y08tf5tfajWJn2OErpJ0rIWx6zlJ3/jucd58z
vyM3T6ggKtkluT8/bgrIicNMPoCQwzu8t9x62aSNrJMMcQR0pdpR5gaorFQlXqhHGzNdN/DZKcXm
S2WzArZBibaj4j/fTn6PFON6wknPe8g0l53G6cOnz89xuUbOuYLN6TZcsp9E+8SYDAdxPLSkDYzU
z/YnQVidVHO69zG5/qiY0/AJofysHgrp7mX4qR1vnly+PneVnJmeJS5F4s+k4ORwI8iEb4X/e7ZM
pqB3uy4GzXkO9hVSLDScnwInsmJdwfay+X1XYIAED+e50azf3vanTUTOIa/el/rQPZcWjdeljfbQ
Lvm/VArUb1ofgelc5KD5zbAlb4fe/Yi5n+RRodAm+js6BKp8LSQ8xLNf5faeaOx7vOS/u/mpvI9B
ChMfHkVkLorYAXqSN9Ib53KIAdnWe4WEY2zYZnrGHsrcxcuaTZ+ePb3/aWbRxAKxg2ewn1yeaH/k
O7rHldyRR7PunmwSg3KSr3Yg79mQ+fLLgJmNMc9w4LT3VO3DdfwEAGNqtreK402lmsRTlCewpXLi
ZE/N+tyj39en6wH7mVaiImhlJnLNvOKheiWLtBNJcL9cpWbjbhRBqrSioT77fDZ/LhhnmMAhoxjR
XQUV3wf3uBiAdue882NnT7sx92W5hpZxhPBQ0sohxvAQi4xNgVzqTPXr9uZeL5BHvbNq1jo01s7I
/Z4xZ1uZ41SP4fxXlNa71+rLof5FOj9+OnYqUyVCp7PgpNAahQBdmuGnw7Ifb1jOZCk3gnPi4im4
Ab944JWDxCuZwZQZFgI5DV18Zr8C8Mrj6B/srAjti0/DJKu5Wou3t7YvWabhVAxH6kRdeTYaXbzy
i0abXWnml0yGmFRxTix5rszcPCa/fzKfswySoh+cEPAzSu0UkMWGxKVfAnFzTFFa+Lxw56M/wQEb
XYM0VIYlnpAwR5IbpnQQTTIo07YtvkNhp6z4YG0MH8rpQN8CIsvb57SPY45w/ST3zRcsb8cnsOwH
+RxneO5I2ybBKzqiSTWAByScMCS8kSeX7BRppftgpClR5opNQpTMVfbzC4MU+AWKbR6svS04KgDl
XX3OHmFva0SRg5NWtC6W7fqJnYC0ivGA/VLgy65doTiy/IPoo1KBmpg6++vs0AuluTMv5daRTelB
2qawA9E1u57gWOkSXNlgtXEiG1TyuxnM6LygTzqOZ/2KUkbfEs9MCMZ33NjIZQuLnRq0JJtxKvBo
ww/N29gg1IlYKzHcohLj6NHl2wzWGWNka5m86BlQxGb/p3uDCnQzohvjq4C6pFImk6Bh/efCByTs
MMUfmjZcWurxunnc1xTRKH/fJHMbaW+RhQJDKiwdKCOsDrZlMTOmx3FqSNe4pyLMVEGrf9btyUQE
+r2svSNFA8uF8XMVyYxFAhBGPTzwhltxLyyONvzfaszu0Bn8huZ+eCDxLfhprqP0EmQ1jZ4qg8hG
P/P2DeuUxE4l4mpCYnzVVsmrPNh9Nu4QreD8AIk1aIARlOLBQrrx2njgVOGALDaWu3F7oXCh6+yG
ptAg8mj3Hk9Kl8RSXjVi8aJ+2sXFKwEj513fs9TUKud2HdV9jZY3R2nvPEbQhoMDOHUYqb0P7qWN
mXk9p1Ti5OkHvVC4mVkwCTd3/nmhsysDkJfhbFkjI+5ARNABuFK8+zKkxqAbH7uoix5ATvKpFbRr
QjALAFjhGrE9ecDK4qJhpf/KyunAUM+Yozy2527LbsSSjeBOImj0KaFtPTYhnJSm4CB9IH5hl/A2
8ih80u/jVKRLY9FnZUrj9irpPBzp5qShXCF7weYDe7QAlgsBlF5qs9UY31A/jP0CV+kPk5I3CO6z
DM5L+2T8/LXGADtWeBpNyEJKWVmlrZJsWA1i1eGPd8rB48HpL9hTsGtbTS4Z8HUAJMRcIchAKWOr
8MNtK11BMXAB0oqHf88n8B3L8tAXrqZUwB9jHm6hQe9i6L38jy3RmKBovdwvfHwkkU/bmrqxdjMF
d7SnPafgaSWlLGw1wOa9oDiBOQUQ0lB+7BXYR8Tay9fu2U1vSbNQa/uNW11veN2KqgQlATUEU/1h
2ounKSOlA+30xoquO6v231Z5lJCV7aLrwLQLvKp7doR36d/2YjmwqvMzHjJrRq7eNyG3+BLgrSDB
ouXOkTFA7RCniVY8z48pMGGOCIeZXLG9xdXA2dA5ktC8WuNF5u3r2wJivudZtl049Jb4j3H8md88
aienES9I52uJsZ2vHnFfnxshZCWlg76VU+fcAtWLHVlAHi7H8xtRVoEacO7Q2giTSAaDhrDNBfZb
RS9+YFzNtgd+dOgJlIoZTKV9yn3HcOiMR8ChZVbjTJEAcdBb3BJiZWXlnM+sUFQKF1lNmirQ/huX
OCZyOmDBqTueikBtnAdhwppomZMMBOJ9tsFhLAaMSv+PbILH6AqpfIqs1MeIdZqz/hT52UProIqt
tVDCZQ1iq9NNsKWe/HVz+gwPyoRSspm0pnaZN2xFqdLUf4KXa2FjgCGct1ZNurHxTs+0C38CLjs+
oU9TKgKsJWWYGwFGO9qWzQcUprAiGRBTdyBEvJvi4ReaV8SHCCMk8Hhh5efobzn6zI7XtE/Mm1EN
kTagKca1UceTOouix6wxyWZ1hf2ruaTOr2aIB1aXXkoGQvlvqwYRlL8/AtsZkxGUWXSB0aog4co0
jJ3it5KMyHq7/R5d44fJz+wUi+LJauRNS5KoMJ2q2YdFC/7cXEGXfWarw7m3shoN4Of4s43LIlZC
0rJAZPy07e9SIt0BIi5cY0LOxttGwwtIOsaE/R52S0eK8m1Bmxg+SSHtrww/7+yqLHWc57zxNTk9
IVwk23Sx814VtDhaHY+EYOle0O47PbiU2mFn5ZpF+Y2PTVxH6vuXfE9UjUA/Pc6EKui6zpx0+sdh
xzMih6Sh/sATerlSbS4+UoLQdS/Jk5X3wo+WnlS6pW1uWHgEwZ63Q5qcRs0y8aznlTjAKN/S+nWD
gR5PWXP9xtQSxAtYw509cWbmjQEfDBTyBt2zD2l3DCn71+BZG491tk/B7oiatVPYstvCpZOcaIuy
drS17MMGmzCSHB5TmwtLd/KB3EqVllgBgzd/2sQLOYpjJR/JTtOgpVJXiaeEk3h/gc2D/ChIgRHS
/C8L/DGQY6/y9XSds2UzBQY9Mmn4z2svLrjFjZusgGcSccRjtWBP0g8WGMHUiTHB3ECHeqcWD3pY
cnJcl5zyGRWJjyr8hY7AFtOFIiIUSGFIVcqHoJxxnvnt2YBZMYGOFTEry8CaynXgplyBBxb03ajG
Q6PkyEwDFOf2JqlI4Mz3DZaWKTWlnvCTgWiU30bCKNChebWCF8trv4qNpKtrO7cTfNvy9tCal96p
4mNRHGgcpQo0cIHE7+bNRkPRZGwMKpIAhzso3/jXoPigH2x7VmR2bSh1ZsV9y0VI6YJU68XjUeyB
bz4WXQSH2InisZk8o5+t3XSpCYFoHT07hiaDvlg9K7NzWg0M5OmfKTFNiy3YEdD5CXRP1DAscZKL
UNYH/D+DFC22nCkUU7+t41FSmwgLUFUyF6vnMEnRJ8EJpXvAUQLadbX6iVX4reFNAIIQISBVpuP9
0pmF7IACkiRvUwKTT8j30KVJBubocimUyucdtp4F8jHH/K6uaOYWno9SBukqwNsK3bZaibYinmmA
2c3fiGSwPtvFsGawrrS3GEKexqzDqJz7SgcDmXwWtsmk36HzcZoNEMINflAfMTk/yVPywjUUw/JU
DcrzkyUQflf7P65iwBYBVL+UD2UfFLo2GSuNZSz26C80ZkWnDfDnRIjFddjklFVOMlwhjNwl8o/J
viqgy8Gt+JfseKXl8LeVKrDnadAmhVAZsRduuCuEfj81YXBarEtPe1fh/fqh+IV3QuxxKHB9SckY
1DwL9SIiWtxcrzncbBkhj0XCj+GzIWXnvYaVMBjOcCMJR2id9wR1dB1+TWqJv6mhIoNDajs4XvI8
13kz36qWr8UTzV2g8NVvIi6YwewYj05yM/tFcm0hvPckrRxON5gdOLLQvd3kwwOurEONwhQCqPIt
IhH5c2nV1ngWPXzml7ydIq7gJO/QkMrfaZJ3+D8O8kkWGfrgpFwacTBSj/y4tUiHf9zGVpsS6F0f
HsA1ISCHlLKWuGJIoBYCMn6YvLTzFFf4cgxuclBEAxdWt9VSPImqX+WdPwhGylLTzUaPXoscQnRe
YRH0uYL33DCthSM2xOS5V//SM75j6cCTwcPeIv3wIg37mAQf8jOcfMX87ymzzwjxepZXSvn/AzpG
jOOc25SvLES4eCV9kXF8lloKX3KML+eITcKNSSlS3O3rpW3Dje+i8qUUSTtblQSb0eTmod/iTYGM
iK4vqZ19a+dgmGqw0PLxnJLsdEN6kMD0dCxNm0MGC5tJCwS84zo5nSj//RV4ZfwrpYb1hGQEd1jp
BYk5/flUhUfYiL56rOpt9q2Vj4YuITeaOiOi9KuIYi0QVxZ+UntqJdE+z9qgli9Q4e2pBF7bnmov
PSXlXr2AIlWA8bawebLlrYKIa7NfQOMljplvd4A45C5+L2zmaJGnZC+H2E8qO/nAY4iMHiuRCS7S
jp6NPlChb7WU3mM+o/ulStyZjcmopi6lySmweCLOzAGl6RUuvHGyVKe860jKXV0bM3wy7nBN1oCh
2TPL+BH5yj91W7WOOa2JiWC7Sb3DaCBDmvNRDxjvS/k5BWhrIjrXQ79DHRFQPB9JIBj3dL870SCa
S0ElRuU+XD1VJwnwuYoBBXJDWpvuDMfbNj03FOLpgou/5Gr5O0guw5hcGHBLaXLSfaCmeeif2/Vs
mqcCFZR73LNdANyrvDliCQgWO0zpV6iyu4TeE5vF/9k6yaXE0vuB9hWhrpF7AfYos2QAjeZioV2y
XEh5EQAVewomwa80hvL5JsymEQzHkhQi2/iUdzJCvKr72YMMp/D32duwJe6NYnIBFK4ye0twRIoM
sms5IscWsMkHizRbtU7cCBN3jb2mHSUSubCIjE6rYtC9+5JYhi+wOgDiYzdUX/bF0aIpZCaIY5z/
gMBBrPWKpWaI2xA6zxKUDD15QxaPxUFi6KJ7IDBFc3ubYQU/nAL4EkXPXHrfTINuNFcDS3AHu2sb
mGPhUdMaVxdOfpqzP/9OcHMdAgLKH0AIivzjiEdFkC1m2ykhagVwFaaAn7VWQdMTcM8E2eYpSFoO
Vs525pzNWrNVjwHN96JwEkQ87F95/SDQDkWCcfMGzX1+jsUuD9e9pveQJkRzVmwEXasmcDQrTPeh
7B2aDCoc6NaysfTASrG/r7QtLmTTlGBp5Nm46FJgvmIBeINCVM/Z3uoAtqfH+wkYuugOTswEi4GF
+t7bspjLXVLGdmHLelNBjqHr3Y9VqvN9uxgQwgi7h0+A+zi/x1r3ajL/x3hU6Vs/TY6cBOqjC3zT
4RQIeB9qMLFtOxw2TeHHJO5ufxmYPZgtoob8kCcYoNEfQsHjPwEiMsIChVwEp96tg8vtDS/dRKuf
rA4MTfKygX4zO1KBNlz7MLiZjbkMNVTVf86JZOsmurG9leh+ZZ7gvHSNqRcOOg/FdAR2g3OOZX9m
bWcMKHG6FUmbs8bJbAzryD65WUvIB5+ElJgqtxVWbh3ynj0zEkFSmh+PYUaVJ1pYvbjJreyNMYBw
9fpL62fFro/qdg5w+BwE2Wx9czm2aHAae1UtF6mp6CEa7SyZr9Ulpi3UsGCwd8cQ62bRQ7hCgwGI
xGe+OM1GAVkZV56dvTttoxADocEzpUPU2iLoV8fSX3Y3kYz981oXO/9vdegboyGOg06UNBE9BrGA
AfA/f8jBDoDj+nANVMqii1egyOrkU2A+tzqIjkbGDl6U3pgHifCmujMEyUxy4EpMOWY9BoLztQIv
4Bz14uwH1DVX8UvxJpB9AgqnC8/U7Q59D2FhRUzV3Pnv5ldcviakyVd8N/6zYXsan1OGZjO7Fn5Q
EoXuUi3O5Ng9wF8Onq4hWd9l/+nbjufRxt5h2RqRSIBJMrdgm2yeB+RPn9zhy4+l8D1jZ/Oc6Nq2
tbOJeCSHadrmGOd68utvK6li37D2IUqK2t83MgPPYJWBz60ahSicnpCC73IznWIQxn8Zo180qfFR
NzQRt2Y8OUNq7VunhOpHsGzwKmolTSDsUUptl7TTZ6laB1E9p3FNjhtoveyVFF/ahYkmOH864O3T
f1Y5P9PUar/mwUggGGzt29f/W0UC23L5XTaCjbSaDtA7lheHx8CrtJxAoQ3B+M5k5mzctSU0jbDw
zkRc32G3W4qpdvTf9uz7ryP9CuU6Of14GGaPM7xZfekoWBLMj42gQK1lbmP9AjX4S0s1vCi6ZNX7
EdBc1woBXpu1wGslDCybssv8wrEYadakmE9ze8pdNfJSwHgoxCYBl2wslfLfXPxB41LCmzVPyD7r
Vd/thau5kj9549gsWJIu6cVux2BtmZAi2zksqrL4oOb2RBLgOSfaZ4hjKJi72kgr2sdtGA5ZjQjm
fmKLT8Kx96SBebb6SIteQgVS03iqdHHZIEDdXD42u3T15LQP6S7HW/+M2xtrx+o9EM3AaZvSy2Rx
6imivwXfNa0VRPgmjSTOwxDGwKtttZmhuXvV0+qJaoq2dHm+gvTWWMPYytb6C4wx3gSkrOjaPnt+
5jpGPurDIDIX4gLJrNA5tdJbTIBgcwuUzkXdiaF7okT6NZFTY2CXHb/AVmUBFwTj/e6kUP82YRD5
cDHZSyLxQscTpMflyB4Veq2u+xJNRIx1ZohV/EO0SsbI9jATNpYlhBYjlJMBhEoqR/8ThQgLMD50
RByA7UDGzmoXVqZ6Red2ckWxwSa1Oz4uKpsqwuUQpDnJTBmU0cxQ2Tyyv+OA4EPBIejYBSvtIJeU
y2H4KuzuEan1TD7fxzoVQU+mAZ9M8DPriZjV5VPrSMY6cqQGqVmYohD63/Dclfx+qFefYVXt3hng
Ry0DBjoYAaqloPh+433GS97Hqh1coyNJxMDuunkWoz+dYjiOr4Pw2UFIFxJOgQDXZ20+iJeR6TRj
RGqUrTqddXxKs70V+lrFUJ1hiB3nXSHZOiTCk2Y41iMAQrCPuFOZw/J6o52lOHPYJjiVGzV9kqrr
olxn48ePKUFtXYjy2AlPFgKa5fjWxyCdf7MQGbYEZyT680kG4JPplbtItnOZHjxdbdYTU05VaUg5
i6W4C72WERDzjwbMna6HIrmAPWHx0JpjCq/XlCBxFBG+Qj6GL02XFgnV1QrdHOzaOF3dGJEVhC63
z3Cxh3pQmEGl2yrxOVNU/suNYixtPt45k3T+ag4zt8/9JTGPJS2rcPCKp8rCFW+J667sNgVo7bHs
q/L1lCIQIwgfSSEXDkY4aYlTRMAvONtfKb14Jt6yzs66055iyU8eershlQV7huXvH/ROE7eCjRvH
TBPPhAK5AQ5jMoEYJdQnsrxbRvBhFJcaUh2nu3VYDggRCF0vpyU7pBvXvb16fOTL/k2gs8uiXcgX
JH1jci5RSpL/uQ7Sg02cqZReW6JIzxBLG8ScsD3DdeTFlDJxqqcA8mz3NfdRcnxNgRjzb0AKiT0v
0lPGE3V9V4TRk8MnmkZmMsdMtnOoVXDUT0eOUDVdXBwSJ9ywcUcVGzoH6RVQEMWO+CNMgZJcbEPd
ePw5QbpYG7JWc0/begIbhofaHq4dQR6QkckoFU1H4NcY5tBq3hGW8ssyOeuT9ikLnoaFV+BTU9wE
1CPpDRE7Ob2PUiiMbibNsG15xi3rQNepTWS//Cl7Zo+BzloSuP3ozFmqylXzGG755Ru56/MxQXYc
o5BgSuAqF8/RPxSUFludGioEJHj/B5XTtl6BYuQFIQbAz0ZNMJrbhzqI3rz6n33/YWnKIbdrvLmy
JmoSzNOctiXLyvFPsjXo9wfIOZZw9ApGzXMOTUANoIe+0lgC6/nZcRn7mYxUUT20htWu44PQz9Cb
RdbbQSg5FtqIHQ0nJZaXoNIxEyD6xXwdBic6fDmRwuMzh8qya3Ls6g1dx5i7TjqHXvPzprq5yIZl
xUQ6dHhpNdByIXsutMp/dSVa+JzY1QNGYzo130Cn9aEbuZo/0warE1Cq+RoayAg54Jz0YDRmOne8
aTVdmMyEczyH6wKT0bMB8A2rNjqSQhqdnMRx5i8OoTTzJ1TZPKHdJv2sZCispxF5LRWRTKg5/Ho5
M+/3JEcLb3tD0VgwuoWS/TiOArOQDU5GiaX+2zcjy2XzWutRWYwno3WqW0SNRw7oAbUzIlk/zAJ7
DnfdI2qvuGwO3bzhEod+KSGLPeGqq0ChXsAIe5ZyvL6rBvvnOoKLERt52Fk1pQnTymhPeeRpBW/r
/LyEsseAZrS920++HgZt+TieKRAShp+Qw9LP+OOy/bZQncXleJpMYu9ZoNh3c01edn1Ropepd+s5
W/qV7TqpkBfEb1pV2WRLW6anBlC4zv65FNi6G66jUbRpf4OvEzgQDuU8yxB/ixcfvEd7V5K/0SCe
D4L8fvisq/ICGSp7vfWhffO3nTQz70Zr5FFpr+IvN42AgJJ/n04VqHzNwpzRMWh3lWDNmBmsIrVU
xFQfgdo9KSIq7ckD6FP9lqu0n8g5hFMKhhVxxPTBZoCVHhXtv/oY8YiXb4RiIbWdz7brOEtL0qj4
HuJ9jQU1pvhet+5kWbxA0vBrCsu+z4GQlEVgQoQMhAjtp6eOeZ1UwkUh+UIcys7CArtRghYQRmsZ
1XCORBiEI8LJE1dcyFsU9TPnMgyYwwqprE0eFJlm3VBHgsOiqwwGftKr002D7mKak7zM0Ao6n1V4
tJ3qQSlw/pUIhJd1Lhe7AAsYFoHFW4sJbzv/PQ6NavzCstcIlCTw5sZamaEizE1INx65ZEaOHJOc
dNsCgig5NAw2nMnb2AL7w0Q3I1f0BggAc/DMZhs4b7Jq1/mEqTEx/kI1BX0gNpw8XhGL7PkCVTnA
/71sgN8IUUcTTQI9o5oK3kKTIz8eVOQU4JbQit4qW52t0Tt9UYnvuoATDVQBTtne6klaDG+hoDtb
GABNm1Sh3nfrg+/h4+on+zTv5R4v9Mb5+a04lECtKtURdmscOxeLO3g1u//3dkv3Oj7FoLQvJAnJ
ymEJSCiSr8kkWT3QFj89QxL4hJLS94UwQFXLqcArnowuwoLzaLFizd6T+wYcrrnuIRmubZ0CCjEg
2xGvswYiVtgd80YXnnfCdaYDj37nQKJVFkqhbG7DwsA4EDpvVa5ojeKs+VZhPhnnEBfql5Bha+jO
TwBrb+Rf/vMHHdn842NqkdsGuI8hpOFuKInpDLoDOL7D3G0Yr/N5nugDUg114Gq9BvnFKcyqgCAM
tueggbj2psrgoLPZGqajdIFHy9E/IahcQ5mTnQLaCNgze9PQUEJiuKA/4euA3m1AA0n3sat73NN8
L53/gWRV2o/zuug3Uq3xpJYYvGv5B5ks2n578w9yWUZFwvL0TGpHTgercsCviiNBcBWD1VqrNeDc
dp8W1qQdimHofWNcQCt3JeFrIbipQHHBgZj+43U0lQGx9q+9mq4und7ejyF6GqABxkssUQJuYVeN
+YMBTAo+g+CzDMAdFNz/vLMxqcDAwGaqjtcJViFAKF+rl3VRjY2LxXcVGKEgsXpTbrhmdN+fRFcl
4Vu6T3jg1HnWtYtXwtHuOGnBRxemRTtyVh6G90B8lLKn0kB0gVlo5K2PDGt1DEI/tp+7KUHHzy87
dcK08H4pLdO9NSXEYYj+h9/+YR37mH454WG0S3Vksd01CzJOjgS3B9BbaI2L5d7VK9pbWU32v8qL
RC9rtiLFc8wJirPaYA6FuZc1i2sulq9xx8hfkrUONuX4QOyQg0Wz2kdlmFOFfsvd8EdfOvP7IqB8
nEHM8hMukEWJkMFcWLeAjJg5cy5cTP/bBlphwos7+GmzZTBReWzhHOwbwSPthPB/K/6GGr6MvNHY
NXzCOP5EnKOKXySUOlwj+mIlncgTBkRIfWXZv2tPIyVQvEge6kTfdVFHupAYAlNCz0U5fx9Y2LAs
NQe6S+GXFvV5YiuDBH/THpRw9fmh82q/p3mP77v7Y1ZTdM3uaL2r8F9HdPijTyDL2iBa5AkcKaIR
JZIf7Fkqw9WUd6SPKP1lkkS6j9Yio2tkNR5gVf0wUIRgxmsKh+MPhC0yJg32Bbs7OGN8lNw8fTdA
YWWAI/nB2aoy0n+CACM6EAvT18gLdb6Gdulphs24aMcOZQ0s6G3asA9NOtITSo8EvB+/p4tBmCQp
xObu/sdPdF34dsIMZaNHQskZrrzyvJbe17aPSlxN0POUCocCOfbvGfITwD2y2SFP3H1nF2GQucFq
lLPWShux2Metbm+kHUUbXEP3cDQjVe4duGuA3C/WFrh9dnPNI8Twev8TO4UKmDrEogwuaub4LUBp
EFRomoBefSO7bq54tMQX6TUOqUGSybZrLc0+yewE8cCrBZjCKdWaDEChkLAWmXIwSLm0aSmmTbP0
GERk6HycL9samgfWTVlBxvam9HKHNNEE7QR3M4GHn4WSh7j9NYuUXKaGJEIoNMc2MEzBijkzsbf1
R3ygjvXySBsQiHWk8tN4y1ZsAhvDRqN3CGqGvgNXMJC1T64+3bY57GzyATyIxRs/SPhfy0X/k6Lj
ipHW8fNwEiLG89zCf7JCKYF7/dTBytGsIxT00RHBKO297MJggs/2xG7KiTd5uUe72chCNkepyl/r
cEykvXDA8nCWQ8oLiCnao6oEipH1ypbqEuTMoNVjhR8RCht+SF2GeuxNZ+549AWDHyyK7oaPieUC
fWSK7sGj9LnpYzyi8AqnrFlMoF/iE/7C+ZLDwA8U9jwBaMkDHDjQsV5qrFujtXPylT7bNs4Jw8Rm
v0ngGYs+Aoyl2ZtKaKkogNSBDJ0gwcHs+oZIFyaw79a0ZT5tlc+zNEmykFoNUQh4bWjYpkh2Nk0B
D9vhUzSrE6jZFsG6keNgJoPsDAPCc1qfif5xFWhpIpCUt6lry/cFLdVpNubEedHLyPsYXcf4hGhm
b4t2nPB9tzwJHMgKmTBp4Urxnzpowd/CKl//qHL7ib3QjIyLFQlXBG/hX4LpBcLBc/ZT7uzP0tAl
0QrZC0FJgPKjE8qQRTM7cNDl0NiwPelnq3rzUQPd/u7fAM16uigGTQQUQAATaqVtKIEjYRUho7Cd
URIwnCEvhSGgdS+6k5xeQN9hQVAfh+31H8xjveI1qcVfofWfoz0OIxEatmj2Wvjnvg4RYtXHltjW
7q5t5Em6vI3I3J9gBhq3Uw+b47qPRYunq9Ks5++DJX0fZM0lz22/WI3gtwENY7rtu/ejREaYo3hE
nCj20dyavgTLyM50itHGPDet+GMcKcVsZZxlF1lP7n2U4WzP8ayBFObTeg0HXd3WNcFPuM4JnAcJ
hjFIWqnP3R7M9HBMcXtXOcyMqy5yeBfmoSK8dVd0TY3Z5d6ZWDbzZaaM8NBsigljFBBEixP32oBb
/e93IFixzuC/ZMF4JxP/bAoanNNStO60WQAJclELDpE+H2fxuQbu9t8QcYXn2rhQliEWC6jLbrEb
YM9WVBmUF333nlaxF4ajvH53j6BDtJnN70Rt7DczpQi5wfs04cHH+8ndt8BAHYB75lPmvXtZNvvd
ff9nsF+cM5VPkRUbKJWmEXfctgmZ61GsC6ufqyfM1ge+ELePjwm1lAZf1JkIhUfR/xBQbMVcWZzV
TvR9XUu1WZIFG29Lwp7VeO5qXtxAnWfQxBhSzcNWh6IblFi8ItHUVtQ72IdUauD8rrARzM6B5WwH
jRfNKcAjeRKahaOnHb05OY444U4XQxg7muQcbIyrBvSICGJUXs1Wy96R3sULI+pQ4a5D/Wx/kYpJ
+cJg2B79BQBEJY1CfHDuZ1uJa2mbPAHMrZQeiY/TjuxvXevph28fvSjtcSBTVeGZbdKZ/tj5jRwX
iO1XfesfW0HiWHStWaRK5nip8y34qGZNUuWml4y/Vbf0WDKKjgptpnUpxXNLmTI8qnqk5QpZXiTw
MiHSB6smSf5zVHbubj6DLCjK20+QPQs2DCZqfEos0sxGS7wU+lYkVmyZxuNzrKKhcxNg2NCUED0U
+/BOVvGyF6+PuNSPax6DU6o6Arn93rb3eemuanQdCluPuKcr4ILSUNG/Fd4wClPZ0TjQnFDGQXwV
T29Dpyd/W1ya2rGqD5QGxvvZ08gO6bKRBlEGF8m7wSHagX6ZWeTs7xSTVbLLW17kXvwylKFhpLtP
TuCgsqaJhCOiSLJ8vP/jK7S9seUESFgPuteRJpIXC6trSF36Ibq9UjYGrhWzdIbLWKjltBezlZff
f4QIoTot1tKfiN8z4kPkBRA+1et3SVqJQdiiT72FSAuveXNcwkpRnila4WG+C0yK1eWPVh3V+Upr
JmMqstkr5m/K6YqJedcNO/i8M5hQizpQxdr8YAPdPZksyDNV23T2trNR9MAFNvluw/oI8ZgaQPOe
NG7DN5ct4ql7XJPna3NUbPdmXnVsLcqQ1uQ1wOaSIIa1BQXjXx7RPXtxLPyc8m8dZb86mk5PARhM
XofKmZCxtKSGzbRFIkzOqXrJQuliAMtZsBiFmP3TLGfK8I5ln30FrT4wONZeE5jVqYRhsmNViTqv
ZA5kc+DH7EZsQ8eYUgKB+2WDIq76oGB+TwDkhnSsc0U4D5uAkGH8LS6nv6lMZWM3JlVbqgvSp422
IIBJYYbbR1QJSayVUqr8Odu3+Y4Zl/D6Y8AksdIfk3OKs79comaLnzD1HexHDADwthFrR2zXL57t
bt8LBU/NpdIYljCeWg+365CmCHKjDgmBwFmttEPGOvO9Aq9eoxBszRmdittX1NapA4XV0qSCNzwz
KEU2N+W5R7RnVV0UDbK2wSwVINywYdvEPc4eAxdsuIqruQK90IF2+LZfVexlwjMdYbn+S/wgSWZi
VopBP+9M5bsg15wne7+ag9/NpwsZCwf2tWU2/NUsGCTCK5wSfT6HQlgr0k3wcIlCY972YmqPKMAC
DEUWBMR2BRcRnx7FWp1v0INKHmH/lGbFXbeIkX4qxTHhyHDM6hTpeVhZaPuzEBY1dAsXiJJqqmrB
aB/C1KudMTCMNF/peFvWXhebTDVsDdp3zfe4dqjYPxZCAG7y7IQ9TUKFKVDlzSMdvNPWGv9o9xFd
eTuVsZ1mwLq1sYLUJ9Ji6yXLa83rQaV/uGyhXPJ33RrikFaYJW8/lXoYTCbxVj1kk26jxoVGKMzt
xROT/PBnRtsCfK4sY0wtgZI1tjTk1IAIG8qhCiMf7t8KdQA7N6Cz+bAO+aCzu/W+wphRcupY3FHg
p16wFzh1JRuJWoabW4vrPuNI4BCuOEIAlbf6lMlHYOV1N2ne1aNQO/XNZYwx79RgYmHDjbzMIVfX
UlT3Mnzf+gFuQe76dRdut0OOx6C0ZzRXtz4reLVMcPggu3OPatoYVde8jntE4b1pXKktlGdAS3CL
FRboMYsFTdJdKmX/uga2NM7HtmAatZZrEEj06Weo8lm6JhOuTqKpdQf5fTKV8Dt+EX0yatNzG71E
2JZ73AbOxeaIvj514mEfTrXH2xZ9b3lSsbRCBEQZLicWcpkqrpPzoVZClzbtf2ncULwmwqoh6aBg
0OIUiQ22mTKUVJnvVfep602jbCkWf+Z+GrZR+Co2tw1D0Jk+rldBNS9JZ3t9xNJZxH4I+2MHgt3t
MI+vQ5Tr+NixTKETHrqCT1z2XiRtlkkt8c7swuiOD38F8saLFfdihN+8hwHzts9IdK/posf/MDK3
XJaThh/nIagwTHa/NUVFLpE3dhAP5grdsBc5EnJeGnJpIQ0G9ibVaj6fIAEIjGbasjlyFS+6H4DF
63Ow1RxQoTTwa/MnuBf3HfQl4fK+OLoL2tmnjDGSxAdMdEUcdOqghmQ6HhZOJWuJWduhDsj5HvPw
TSzUPgVXSB90LEhofDeWoJBVCcFmKqSlEPHEVuofuDZC6wt7jE2EVa3EWjd/TlsWlzMjUAZN9E2D
XnBOfHSfnDLjMmF8fUZNIUbf/woT7tinaWqPHOPzMFBbCu0MRyka5wDsEUgsATHFXUmfN+nmgEju
9AEIrybd7CDA1ygdNVPUiXImIKCO92HLbuhHn1G1Z1iFtqgjbN0s7Nz0xgYfjnc9cxm0WmWhRz3x
gGk6g425Y4ptRrTovBGc2vCh3MSBsMy/3+IjA3XMkq2VtPn95uPPAE0gNsNYCvJ5paB0rDJ9h6pQ
V6T5Ag8KH5whxsxBxLemr9RCAcFGM0OZ2GusaDasS/ZurC47cURwKUYlgB6gHaoVGfLHuCGw9gbf
eD/13lzRiC3EEN1hf3OfCmiTrjLsbFycMbFL1Js0hT2xWQwHz6hq72Sq0WVL5wO7L51FLxAha7CO
KxWTNe5DbDoZnAFUXnCNwaTnsQEu3yxBuBN4A/Ct9T0u9tDKkNBoct3IwMMxA89+4edUjkSwMmUt
hqRUpPrBAoRMvbdFCJ6hzyJgaka4Z84UcmbafdwsYojLzQ85oXBIl5Sa4n04LaDxbKB5I8/0QpiO
oE4w3nNri6MURO6JBkDOjaa5Rr7t9L9yO3EGLMvP+pCLYvF6YdqaCT+FhO2sbbNankUuUkPaBKd/
NdnttUBXzfsoR94HfTPZwUjf3D5n9uSpAb0wPzsWB5ukgmfE0qiTqH6moyyCSO6CbsQx7cnaOnlD
btU1SmqZV81Pe8krLg0UtqMfCWZfHlT8zvUNzrL3Tok4F8xNlJjTd4X3wWdsGiVsyEXEihhhT7t1
rJ6/H9cyAGbnLMeNFBkVNaD7nZ2mHOsYDwoKqvmYO+jKetgbIk8I8MbrmhVhF3fO0PU8qp9H1Ni4
Vq6CxflPWSmLiwnhk2u85ntxPfbX++UPcqfrTwJ/26tIRFcMQvKtUToyqY+cbuwy46DwHeq3sMM9
v2hJBedT6G4F1r6Kz617Y1i7BAI5pN1OCWvuS5JfKAAo6dbLJGGZ7R852NlGgIEwjTGxdQhGqhk7
+Gt07uJebB3Zc89/9jjQd6KKQpF4oI+3Y+HX+MEhI4okoq+5tYMgRwJaqmdNew57QQQJF1fBem5w
MPjvXE+WSXujPJDxmZjjuh/P+2F+jF+QgaYglOfK1o/S6ibXC7SEEqz/sX3c9A+FGF7e9yKj3zzH
h32LzpPiVlf0OER7TmFz06YEskTPduDVQpeXE5ZY17k194IpGzxab8mKDj/2LPshvIfnvHgMAr7j
b0k5gl6S35tJwC9XQsA1pkr6TfLDWCF5UNFP0a2huJuS2Yfg4pZ48Hm9jrakdYDpmDnhoX6kAUmP
t+4B6ZSxpSaK+vYNx/ejb9nRmrrWbk5mp+fBflXpJKTaZ8AamTN+QWBX443e8wZrE1VLGorb6aTv
qZbJpqOeqPK02qzvF41TaYie7iWz2Sgml7XDkm4sIAi6vU/K4J6u+gGiSGjkrtiuUe7JjmgzISga
Xa4yR5RkuSnLsCgZBCGydTVyxGNmaDgDmu0Pl4KpYQ5tOu/BkrYhbpz73grpRNlJBbOoddtPIJIu
sIiwuBbvCkaKnuMV4aMQ5lzsyPbUKpje15rU6OnJ/vv0ib6NBX7RpwBHuww0fvOnrWHROiXlKXPw
5c8rjexPK5iANYgJ5Cm0nEZFpFQ1G8h62McyBrX9TLV4UcV7ZVU37lMc4O6S3WdjxfDIRK8sJngl
7Akn/ARWXFXEAAFZ8KavsX2zIwP9BJpEwdxCc9w/cqv0Ij6aVeco/nzY/CRS+nUztXBkHOpGJqUL
aVNTGVsNMxtOwLF76yhBrjUrnQWKIXMn+G+GMHmbyVyVRBAalwMCI5XDSfNQxD0+PnKgNF+vc/8N
witDIDfiCPcEdf4jCrORtGDX6dvFTcjyaKsy9pPifjpZQr3z35J2e4+9bAev7qxObmzYmN/Q16gF
tYzT6K5/zE6QxJD7aOzPm5Xsn01Z6KvHdnP89GCe5Z8sRwd0LAiQpVf+wY7u/uAEAnr9qc2Fm85m
Zb8IBX2Deg+HFtp8f+hfQP2uxp5BJjP/qdjyzrUTG2Y2Er0WpnLWl+ggacBPderelabPGxfxNibM
+M/snzDtRhdVaZ0OWo3H0Q8DzpEWXtpw+e7qtnXMl8eD8yr6Fcc7yGOlrtBMtzK+X4V53xrDCRiV
KzOzUf88m5Z6nlRwoi9ZZaAtDi8lVdaQ9fFA3TQ7TY8cyX+ElKQ6uc8gBds+CcbAk4WEqe4xyz81
cUtJkO0Lpa77JcdLLu5lo2OyIDjk4xWS71JCh3Kc8VFKAdyqjbnODnrkCHvXx/wK38Iw2fzNXxI9
eP5cZ1o+mQ5Hb75CFAnfFWOA/Qz020H7Lta6Dsc7Fl43J38DiymQH4XLfDmnTj6bMKO9Q2pTOFRZ
cFpDmoSy2LJnGzQKTWrERllqq3SuoAQNjx+s0vNidOHLNOEIc5T5LOakO4ma4E5bebMGT/XoAsb/
WaVdh+PA+LdF7unC/uIFd72BK7iqcvw3HX02HsiRWfcyeDQ80bEVQhJej6qYbDmfFRxn9UmoVr2o
9QZt7vmuegP/ZKUQcYp78zDfAaQyjEE9McssVOAV842+MPVZZKYynU4fHyYKZgUPFOSZo17wOp4N
WfT9AAtNyQcNGhMgKkfSSZc8EsrJdDg6Sw1EYpILF4Mobn5HwUbmNpEyBJUSRQEN0dXVfB57d+vx
9H2OaC5g8SlB3zuGEKDI2gl9EAHk2pcXTkP6bqcffhklaTG0h65wOeG45RRB3t4xzYky21Kaj2+i
FVrr6+F7NW+cDfdTYaJNfFsEHufNeVFljPXI4Nf+ekmLbnTqpKWubuWdmIPVljivsxNr/Mh+yLvr
9cbQptMTI1WdhTtQ7bWFgdEXk+PuadNbQmyJpK/1nfKPMJ8CjTwuOz3Ka2AqcLv48AiJr6H6rl5h
k4H9ywr5MVUJr/waMVaKk8F49m6p/BQYLVQY10LazBKmzIWsk3j+A6HXZefR8WBFtJSK3mkKdAFF
QYnPnzKkjL0+gpnMNiCfIbtbGXEdJmW4I+kuwJ2JSEggbyrZV+R6gfG3SKktGHugwJzU3MmFT4wR
bBwsw3MsRN5yw/HwS2lhk0RmiYKPqaIcbZIlLzh5RHeDl1Qejh2/XELxa09FdmX3SiN3aCz2+ZE7
FM1guKzkRVOqEt2v2RsBSpNgafpPX+j84fhnjm4wm0H+aVDoEcZeAtt23vOOxOQRUCkyIZxIqfVQ
3maA4Qg//Y4HFK/W4q1upX5dJrR0ETRwSYrijnPBaVELpnH3jK1fYpzKlGmkbqX2byk6bU98zVyd
BiedGIjUfWRi3W5s6yRARuKKRk4wvLCeOh8FcgYvRzE2qqdmPo+nScEXxeRDw9h4N+j6mg8nI+bL
XD9tQxY6y6ji18boLVTP3xd6RjkPXCxMkk8JVom/9w5Zf81Ai4oYU4wHeMoq3r+m+PGoNTqJRTRL
1pIfvJZx9U4F9aY9qiUTQBVumsjiVmk5M5kYXmpwuAaI/QgIi+wI92ZQk1iLGEjdl0cfkkxpbN0P
8WBzLJYArHvrqdNyZigejp3nEg1ABam1KbD/F56pGfA173LHj7SGNwGIK6NCrBp7R4uZYeM8HahT
qQ1eRweN61BJXHSZ7JRYcSE1IbzJDvGEM/hsOlgWgg5qLF0f5bARPJQ0msbUI9wot19VMUMIGHdA
3OmyRGjqNnvkqjtR3RYmFZ+nXPRyMDL7nLh13d/07RANIQ18wGBPvFP6G13ZlPgcgIl1p8z7ahTf
6StkZlgOoUYLOJVa7ax7N30LYX17yD+v/8tF1HkCA8RLXrfoTvEWAg5TCESDYoEiZbeDTdAONdCx
F/Ib2CHXbEYwDFDIQ7yCs+zs8Ypt9Hs7r8/GEvbe9IEY/TcXRwM34zm3J8omivVT/6vcn+SA1f30
2GmII/tDz7f/Q2AaoNLl/vBirAAxx7mvJuNk6ChV5eykWG52mpTCzM85QYwOWbz4kcK45rkuf0lD
JD0zN6lj6c9P/9FvJ42S8dMyVbUY/HJ9s3bl8hb3SKO98RNWQRlnYapRDF7qJjGFmijSoZDjY6t3
+oFB5opX94/TyrjIIWjtyX7rfQpOV8Qws1gjQLwTvnlvKt25Do0s6jOHV4KqgCaUn6EFJ3sGMMPx
bbTCITuguj9OQUjAI+QI0SCA8OWGNRQ+ZOssvE8gO3LEqXomBNFVqmE9afZsfgh17XJa09niiAta
wgpPA6ZI72/YzQldODIhQSmV0vegCa+9Aty0+sQ984aBAlaJVtII1MiXg9VRusm40RMcOo1BwZoq
6GHaWU9u+irRC3sKEzE8vUgkYsem3syNPhTc7CuYf7HxEejJSUCqS4OSkhqJ0IjR9Q0oY91jk2e8
8R4yYBaC6DEaXpxB0gKOGUS6MTUW0Q/dUavMen/P+Pq5iRf4aTi6sgKfzTTJ1tdNWxYnUs8xqY9y
WObTMyb4/d31z2TK7YmDdH9gLJyyb0vQxOMrYgJed15BXhQ60T0LQ50VapR5oQHtZUT4snF+0hCA
IY1PZ/YoeIiTj5Ryfzg6dJ/vDbHntDBYf+mfd2q4Mc2q7sizHFyhZNTmDRf0opOTndhFSt8lplq7
OKoguCqPwHFnpChGsQgCRVe64uOOeN0Im9enX9AdLvwSl43B2Y2Az6fytaawPUE/8BOAfLongrVn
ho+NHoT+O6CJEH+V3unghKPzF/zhkoIRKgkZw40JkB9A254r+ZjraU2yObPYfkHqeEdhnPhw9C6v
Mfg71oUk+yyYn4kvyR+F7luYXnpwxHkXNqWL1pzqpk0e6i7fBtxOr2tM9yzU1CE3VJ738wIoEoAu
vM+DRBu28gdFq2wlW/fC6p2BC3Wa0elAz/8SC7P3LrVd/nGSxJv+bdgaM2wtCXfS5noAdOm5HjOA
auNdFZTV0m+lS8h3QQj2s3MC9cnhosSZyShiVFJvKSuHVklTR2L1cH14q2LZouDXB2pqq9wmgroS
O3pqu1+5IwqBXMx6RUc+lVak6rEDZPFGu/slatBw4BxThtzddlMBnVRbrOigyBhEIwq9MN5PO8Ce
HCd9aMvIogqQL56dzHukqxQCmPv34z7EY43KPkplWnrevSqdJSPDzWS80E8GP7/VILH7urSbbPVr
FosY209EXbBvAywWiFH+KY5Un0/FcjKvvq58zzGhk8Re//FcycSMBd0CJiSbsM3B6YwU3DIpFj4s
MFzvgH4W5zPKqsg53xKxcVsfV9Bhosv/zZYOC8Q8+0L0QtnV9Q2vybrzqNC2CWmgz31kbnIXZNB0
LJY07xGGpttADrSEkquW1qdjMD2MPyDr4uCdPfCampBSxmtnHKYijQDTREvHtiob3knIPdqGMPk0
V7A88Z0LOUTFAmhoz4K7xZBOVZgl8vdTxTH9gGo+iidl/XGYx2W3uxyhSCm1hhbfAHGBgmXiYrLY
uF/T8n2XUGcVS+rilnuUDGRaeP3F8Zd7VZkrd817B8VS8FL9j+/Hdz74mvEc5GWz21hL3Rs+lkyQ
ZWQBrpV+DElMWBMGXQ+J/b9pbm+VcHgqALjH+60QNkGUczge3LXjaIBnBvm9OLbiis+NcZ0UGRKN
Sp8UWroemNBNXxjUjFduk0rq9lclFt9vDwpyjcHOsSxcl8RVA0sJzbYRnLYa8708chhofy6DceDo
cIaBstB5ZwaOE1+fx3qC7Vp7NAMfFjqpoNE498Pf5d8s1N5zCGc3OKQn+QPXkKUCgolQdynVgcsU
QphcxyHFYrThWNXgzxW6VNK4+4/02ascaO73naYb3b5nV/msMfwgD0gZWjIB66Yd9dnEis+HcS0q
q/6Oj/z0uIW2DhjzCzsRkbC8FlXt3YP0Kxe3zIKwLd+Um5Zr86ZcYwsabiZ9l4I4DQNLmnNM6wRP
rSdnn3oso21QXOF+MLj18BCvDYoDo/5zGPdOmo/poc76yYnG8wk3cc1AJ/DxKUDHo5FwkxmQ2swu
BxWSUUQJn7KL4GElyj44v4y7UN5t6bgPsXWYh1f2EH8p29CH5zqQB4VDcQM5EeP35jIVodO2yKJs
QHvQY2kAaOEdg48de88ojXF8BUMUrXzG8H4JvZrD55k8GHZnu/NqeTFznaBamLVTxPLRVAugQFaH
Cb2a9ywTssdYzrQITy0G1HPzav/lZpJ4tmDqsXmTihGAnFNnJxm1TCRM/njLTFReoc/sPUJeTQZr
ulXw1VTr9msKwElOlCxJQuSvFJXk7Shmt9OZj8tNhB4mriOb5f74Vpu05zo3BEPy7DWVXgFIbQaW
Lx9m8Bv1vvAHg51oC9r3Uz6z45WwF8rT4jllGPmmRoub7/J68P/wEYpINPbbbpaU5IzWPngLs46D
6r3j6uGi5oHoKifD8n3k3IiubvAcWj05NMQL2OjSs0VMWKuEc+sBZVuoNSOxrtfyJ297EtNoMXCp
AGNbVHtDt+AwqlK9VCXpW/RRl2BiQ6orvBO00HEI9uD/AIaUjnXzNCIRYgQcTQZpu6d/+73vTawA
deBKESEvDKmbUyTePxJTft/eVdat3QKExk1YZ9TwC6/RjYpZRnBRG62C7YSO/JvkvOL9CbW99Cwa
tldindySKfk0NIewEhOqoG6frNBptHG+klEcM1xpOtC+Y0bRKIU8RFpz5nMwBMAKFnTYDi2hs3j1
gpqrcB6Hb7vlX/20Y5Jxo9ltXg2LawF9zOMHQRWcdZbUZo99ifYTGj/B7e3f4NGBKsoGcZ50FZAt
dbLHVGh8MsXTqZL1vMmmTAqL3mt1xJLiKladN5Ck5OaASojkO06oru0gLzsgjnAhDyqqKQ9oT5n4
nV+f4RtdZjfWpWJQvJgYfIm3STqOyzxfhCTQU/nOFND/Ad7Mm/yZgnRfokteqY16mHJjvP6cp2nK
PT1yWii5JmHUzaAB58avMQlSa8NQK7RvMKImS5MNLlNtSMi0sbZqKA0PwFfCRo9+aBC+FvQVJamK
/8nA04Ncd30Y1QLBYE2vROrTbdgO9aGyvWS5UVJ7xhvN+b3Z0IqMMxr85VMleL9CPotX7x7Ufmcw
F5CtIFOIA/reU0oytpiwuCLJxpnsk0cdm6ggWJPmhc/xOTQufCwWXp927v/3zKn2vMKTkyKzCzxa
ETBNNDsEx8Uqn75sq0pDbLYUeieDe7Mt6ghzYNegWsqfxbLl5/Ktmpm66ArodXjBuFt5ppczpN+S
QUdTK+XbHgCmRnkNXtk/3mQrigKlVjnYJU+Mi66ns1jFMOCfpI55V4vjL2WBu4qPhR9mlBw6o+XL
C+Ejt1mKgq8SWgBKkxcTPo4n3K7+rIaUVOIjp9MV4hbuDa3GgStOY9NSo1/MJzwk9RQIfT5K7Xph
rbxHq6Iy2v1+J6SCiyaPotDUXmhNXp5B3WaA2j4dSaaphP0h2QPf3uF5+OvNR+1tBiG4RQSXvoE6
s2Igs17PNvHam0op4TXlt3Q2DZpidotKR85SgDbNu/IizsLZADuDh24X8SycZ3wBhASaR9egEXwv
FSYmp4Fx+4WsMLeMWePmF8RSnwUDl7OHGK0jTHWnga46Bc2D9p1h+jubA9B+m6wF27uFZYqrHpVH
pS4A5wh2b53frXFDywSMk29Swl/6LxnZ/+6kGn/jRuxmiQLp8iOsB7D+WfQ0dnASnNbCTTd0fuOs
7LSX6LAvS9U9SLYGNDMUy8OolWQXj3ai3YajyKSYz6Gp1vUVA9f8PS2JQwW2CMfvK7eIckpb7seY
TByO2GSw0240TNHpSmQr3NrEd9iRhj2rkZUcqgRzpmOF8Zn4/Vu7qvx5BOA1ei3EhQOaDNO83XvI
1QCutclVCvDWJYTCCatL02nnX6R0WKSWNn3Gu2UB2qbZpq+AD2xhrQynFWibQex75JuJKACZHHut
OEJJkwTUT9E6jfpbxNDfkaZScTKdgQMlgnm0PelbUA6EK8446IM7b10420CTShrXlWhnm+laP2mE
WrI72FIMl3joh4b+xV6uxa7g4PtjhHoFE1uPhGCaoSZISDql64SlP1fYCNfi5U0z8OSektVcKRFY
hlRDA5c8zfeiRzSeeevMMaQSAP371rcGNdv91KwSZlcXjpPc9ELOMJLBVx7Lb6zPF8ZY1hIAhaNH
QyIRfF7n0vqXUP1ZDv+c03tKpQfTywPKzA1a6bl1UWJWEAT0oW/K1qvJL0w8uowD/nuV+xCZCI0J
XMQcseH7HOdAab/EC3lYEl8NzcEvEPHUWbl50DqF8MrKYIfJ18bUkyJMulniRBL6hHrPUhFleNzH
QRkuZ/SWbl2igKEOvfVqknq7TC9LI/6g+W3/7RpnSDRY9G4swbrW479oNrlfjTb9zvE72A5wDDxD
UUzgy/FpcPVXYVePoUP/D/TE80x7xbT5/tMV7OUYk/6U5/I/UOuX0ya70UNm6IaS5iMIMRbv+l2B
0zhIXrgvhLFkW9lYV8yDjoVoOp0nGFBQEOB7zzldKoks8Hgt0I4m1gorfbBQ68Laaaq8hI8UbjNk
mbGflLFRVYH6Wm1UV+1vvR9BBXe4SPLV7AV8GaWLG/shbdJGP/RtqE61YA5t68hMs98tjrwZwdJX
O6P338JgK+lCrW/kcCSm3EnCckddsOM10rkddILvsFavMrACs9juWGA0ARfW8W6TohRLvZgwExB+
3WJKELniEvsjyqawz9qwRr86bAtnVg8mJtMmUbnZJ3jC6Nh39MVYJNOz4PAk7GVQR2cq42cgSizE
OWgWsoixkHDCEbtsAXm8Zxxi2UuY6aGDyQkLDZSxh09HN/mNV0ek6FtUirzFRQ1Wrn+q/CZ2Hq9L
br6GNrqJo1nQIysrDoBc2KrAxFd3nKTPJVeRW7CGMbMxCNgvRvw7FCFHc4kpiR/UfVwQI+tU+UHf
ZCXFdaFd2zFLo11YDVRkVFYRZ5Yie7LYEO8zmV+bicb6y3Z8jjdhl7S/pnf+VrAQmqbuKl3fd247
Sxsrn2piIdm36s2ACH6Gdvfd/Ki0upgHLrusdwk38RhQOpMtBWPo9zaG/McNhh8oYYbE8s/99y/N
VQaJIoY3ncyOUChW3D5rt+SequFEcRa5+X1aLH9Kk/Qbk3qrRkxXSvJcCbf6c2fIKTrmJuJm/sut
HTV+DNCmNndasbPo7XxEp1amgwmaKtIl14IrVzdIcopPNd+MFHN2uig+I8pllqZBfQ6WLWtDZdFp
6VS7zfBrbtoMGB96h9EpVYVcE8j8K9b/PP8UuR2UIoCmtcd1ank8/EF9S61W/ic9tt2z7bN6FAPt
OOxwYHckXYEBvEzyTIkDrm+CQhl3ijXZPhAVRaBNbjOroBiWYw8UoOiygAlSX5l5FzwwezPDwQZw
5gZtWOfDuS4iH1dpMQOsTOyUs1a+BvV00sYaxYSgl0xLX1LHZ40F/TJY59y+ohDIvXdMeUU2bjNm
N3zpgI6uOMHCXIPubbAOw9oWDQ7MttSJaw2bfS8BvWRlSzKzeomT6UiL6aJGPBH46KXKG7kp70hM
p6NNi6I32lzCa/IugMv+YHFxfa2YYYSPc1rGO8NeRPv9JYfRNIQFCcCXOiLdfkeO4S3z3mNW2ous
fWkSUJ9QYn9Re2Mh6OfFOfNPygSpJb3Y0KO+1pazu7vqMc3TsKNOrEiTLHN3w4emOxJ+rKkSPIQI
Hhj8ewszRH9d4tP2ijJtSF+2ykwD+QR4z10xRgCKkzJozgrpClBox41hy3URxKUjypOGvkSKRhIj
sexOGgTNhqj7iWa6goycTuCAM2mmYOhHKf5YsB2WUF/W0MKia08Yv34qtFlO9FtmuyrvDvnvIK3a
NPO+hPMeIfFmogLPj00nn8M17/Px/zh0sHmmGG7/V90GQPskjEzsdZzM7bdVHN82QbRHf7liNCMk
XDn0HKJNijy6gGYT6s037rxTi4BWORG04lU/7Xai9gunLkBslZdtTn8mDcBEcBTbTLAuqkBNx6vI
bn0B6BEAXEZS9Ctdx5HDjvHPj+FziKCz/RavNZ3LV11D5+exqIte6aB35rswlZz9X7+VPo/XcK+u
kK5mYpexo5D6gZ/LKObg0t0kPFUJVoa5BIy7IbZ1noh13tlztFDYZHa12aqomuR48PXuGMy7foDW
OIGAG+k2a47EP736+bJhHQGSrsPEbyCGzyh26FBS9jG33JKlC1zPp9GDCRRCOnt2y6u4qiC5ztEd
8tTTGwODlDvtDunEBmsX9mlAKn/EquxlVHlb3IEIbm0NJxYDAKQJwO+KdV/CJsWJPqlUdu7p+nLN
AXtl0dSPnLuFa0w+ernjzWFfMyb4OpZzNAP1ThTejEQA9tALhtEMomw6DXnEhQPN165L2fwWCQwR
Qvaqp4tyCjV5vfhIY/XkWdj4U401ntOacycN0eMnjba3PwMC6xqQWnOWN2cCTgrFUSwzvHXTefzv
dN7KC4t4fI7Y5v6Ea+dqnM2QsyypRhU9pHlny/R65NsQGoWGhzFYC8JiMiHvjoD2ruMCiYyBD0pO
pSa/sGPMmOVmGdB5P1hruUFHNOhCHhPNXDb/O8LV+16IRQfWYiN6LK2ZK0Zq6q/QfIcA1ccxkSXu
k7foEXRYuaUWilyWcK3/565P2pIrfwwWUhthUeFAyJw5l2Q5dlez+RXny5Yy5AepU6RluJmnbP0a
Pf2f29PlNSVha4+NH6H/b5pK7WjQnK5FeX1MdrMVbHvalYFlK4saV1tZTHjQnoVS+fQDEgxCMmGk
nd8mNsos/Z8CL6+sp5g67GxSBmbxxdBIxZnjW25aC0gnExsa4sM+VWvh5Ugtb82CLmGiTzTBMjME
NFAkPYIzVuU71EOpo+5EkhxqjRyl9wndhkstbbcAMUhsPmMRWnjQUGjXKpFuKMffAZR92JDIHeFd
n9iGMRtMvY6Ga+DaEVVHyQdhXlP5Sp26UzKsPrYJzI5RTVOpHvA4ZaOGiyQ8+6Sl4/7B+ter2BGV
v+DZ5NjFX0d7KbwdcgZvVhjQkGCs+APyDrWVz67vhOxXgxcck4eCvlKJbHSEwgQ2gG9c7NlRNrU2
jAfZqhiS6dP5kQBlu4BT/77PnKg4dP9+SUXFbxgcdATcWd1vDT6EuCVnzFC9WAigL1W2XeLGgMc2
6fNCIlan2j8t5ve3AlCEsyE90RTv+llJGX3Qur0Tk5jpPnwk+Zxg3UDu8pg+vw9FztuDM5SRfHZf
bj83q7KdZVqI5PLHLpyjqvRz8N8v4is4yiiTEYtfufwbzLKbEwHVmPoXkaKg/CZr7eOrxvzVumIZ
XYQZTTrGcgz9MybnKF2G6tKbk1/sMLNSgn0JvwI3BgfUlBO8xMpCSK1/qIkALElhqHCP11usvgxD
lFiMJlk8zLJ78lrDwOVy/zjZy48iPunejWAFL7aS3w6rvc7v7z8417TPbLZ6NDeoVetGQkNfAsMh
bN2WPwC21tVSAvuRt6B1izCyJ1NGdYQ38O841Qw+IKTtcZPsKwlvUQE04SJGhCE0yrx8dY4TstqF
8R85UgEKZ7eDnOg+ME9GF838CeaxvYzf3e9gzpDIWCjdKsV52O8h3h9LZZrOq6bdWsWp1QAH0sgC
rdBA0KMsXnyYxiVkLaze8GmSUKp4xbJL48hXAt1r3OP5ejo63E+EiIBYeijMjPrMdus1pR2Q8v0Q
j8BUqIorUZNRAV7AHFx9rz/epcrXeFnsLugjBY2a1MyWpCDboonPFyv1Bk7bjPAnnBa6QOghlaTv
aqNC2MnbdusFSA3kXy9uMCnAzFYNBDZDpH0OV5+hSimIj95z0bwdaZQKc8O5sVy5k6PFtyv9WrmY
67LLGtj7ygzECBLP8fTPoXMiL6ToorqXVwc2pnkvJy/DSzGs2WIaH3oNUSEHFqsmElnHJwYbSLvW
3Fj5iCdJU76RrXfsVSJXE4Jnfrwgqn3HqyS3aPgpaJWc7/llJSW6RRJZbPtrM9Mwq7mWOaNpZxr7
xzod+QDH2LeSWzJpCNrdS++Ml3itqxCvEqqYhlyfEiGawoFbGpa1aWNGGSy9eLSSergnMkuXccH9
+O/dBH30O3/BkZE6uedBeMTEbGe1WodpY2MnaFD2dvue87uUD6Onl2CTAbidAzTo4uR5iDAZ3Gt2
nnWteyjWRy+aRAQLuaTvjlR2t78CJlgUHDKbR312G6IxemoRwJW5piHw6KpyIc4DCz6hYik/tEZv
PMweAg1yMjrdx9blIRsnaVnTmBVXcClJwN3hIUkWiVHyKM20etcmgJYTjGDEE+pvCBXqImdfq/Bt
LknfXRJToMnCuJ98SJRsau70Ztl9Ckl1m2tQgPEaDl/21vUUPGjaHpK/JY3AwTr9e8JUrtdHZ1RK
pHex62M+/oo3FiFkogVbtDqn4/+AeZCKIpbfJ1G3uFC0dHTFN7I+uiQSJcQbHwTX+bC7GVFo9bxc
mWlvn4JFVXL9rJY4ts8GG7M/4heI2BQDYpWRLTkS9IrI1JG49yS5t4tD1dyJ+ygOZtQT68TX+DWE
fQnkdBBUEVNZmVUBxV5OE+/VVQXUCq09FkXBe7jFhSSirG0bw/7mj9Wdi+oa6BD4GF81BgTEIwUY
C5NdEF8v5ktNHjmD1ypLpCSoywVXfbNdPKyaLOkjYk8F/rHYKM+wphEYhI+BlfQLpO1q5y8sz92z
DenFLJAGJ+LqEExGhOYrDBIhDJAehsagiYeAxPTUaO9ZFhlSHX1xkhSajgAxReUpofp70pZajZhL
WqgjMFnTmjXmgm4JXDbt2mYaMcFlW3tOjeLzSEi10W+arMSX89XJzuZKACddkjHKPr6L621hOfTk
2Xz4+dyTkSNx65CKW9JQxqMzUzbNOGruh0f6XZkSc9Z8FPDD6m0d2hxr8KyckZJ/XwufR2MFhJ6T
tEzNrJrWeY14AJHyOMYgfvwcC51TfPKco1K2QJ2r+Qwft+HQxaUBgOGhYHWTlAPQ/XEYq+tr/i/a
NOiF8jeOK1ikqmhW+irBOUQYBs0EbyBTldIRBdrXnxul4S2AG3cb4ApMpgOhiWHvXjP1upvTsQNW
/3mvR/OyBobvv2yLn13tVP43Y2/H3vT59hmzFrGzqnSHWJGRfZpjwZrftQYIUZHkRewfa2QywrbO
va8UfrlaOSRkwyHXy281dNiQ3Z+Kgsc7LYs7ZciJsVfvXllJOOrSA8AkDNpR6xSL05SCXC3NBmEo
JF4JEqDEbfT7QYcJ453LDOLw/9o1ecWaj7sCr6TWj+Jn1leJmv0HetDR2FaiMHLh9azmQUCK1pJm
Az+K2EdTN39mCvIy5fjRjR4jVkEy+ZHXGu/qWV3w+KJe9etoKPeh0ddqok4N5wkOb84+0i3YC8WN
vqcf0OUGRCw2PXHvu9cLBiXbQs8cDi1cbGw8FoojahEUZZ6burfbzQsMR1qqEr5AoP2OFwQLThw+
przXBqJUyZ+2JPj0t6ibLMMXxJNCQNVWuMCJn+nIKNvamhC7D9m/7/GAM7e2nxzDRj5CdNkTCc+/
PMW2F8ez/KyY+TH9VwvuFuOQjupddcjUkYPE/7UkbxcaExetl+zzG/J/BgMxMlf4Q6YSeCdb+icm
xbyrfzWmDQQkLp7ofB9jXNcpzWrhoTqaN9k6QmNSKiQ2sLqI+QcUzLc8LPEnGVG0AlDsaF04tbfO
msTv3i3dyG/cHYGg5VCH+dmWN5bGddV/MIjaaYQpMkuXVGshj6xD6/KIZJeP9GIfRJQtERzhe7EG
lIFov8Pw57ERVXSsUknKTW5PQNyrOgdRZvR7hvN546V8DTmNW0hnN2xtsqRWWQo/r1iV7S5xhq27
rLuH8NRB1/6WztYWwhSClg0iTVRv3xdzro9CuICYAGeyIP2+neFwfkVpjgPYI6dol5s8SuJSzhqX
9GZBrrn8rDI3v5Fsn0ZKUXQl362jfnIIPtwPQxIx04CXM9nvL0M4jidxKaSWfg4Zjq2b21QnKrnB
Aul1FXJdL+bniDThfEYSv3Nw4XjWmA3xttoVAevhDlQzDKcXrFDtT99M2SV2lUG4J2R3Q2753wdE
bNEnYFFCdw88Ua+Noy211LkrNp3j/AHz79CQWOtIqv8diy+B49nZflx4hgwLJvOnMu5bpr0RfWVT
5CKyONgSvSOl07FrU0HYJdqJlQW24BuopuhyKbS7pdZg1pFSoxlWgShgX6qSVEER3hhkl+NbUIAA
kkrHRiAn31inGNQ0+mRwZkWLbyG8iLfxT1jw6cBwXW5pgeqhxA44thjjYL1Mi5RRZkMxw4IRx3AI
YB1cdBgPU1uZFqSvOveHPxjkLMDTL20uMfGgJXTiXrjETbyDp2HRGV7XqqAD7ROrLazfWlZNSOY3
buNbKSZA9qNohPIncjbtPnoMamSywpwspMNa9XuKJ/koHEwhG/6n6GNSrKUCUkIaioS8W69cL2sY
+689/YYfkN07+txLLXdw7cJkW4cEsU/fiqVtw+9QTvdBoewIWu7gx6C+/AGphhtRtGfB/owLMdRE
zbyoYSge54RcLiAFQcdfIjDqyIxwmK9jp88ygwm4p/Ix+NLutXWGh+r0BtY4CdOS354shUuuFMFd
JjcJpB3WSTHS7AzoHGpscrpbpjhcYf9F629KogyWX7eLdEDHcDQXOE32xSqJIf3CJuYC4lQVrG8c
QrkLg1PVit1FXhPDedCsGNaTVwen621XgyIxObz3UjDzfqK3C8AQT6t2ouyRQYtMPArxEPN/BQpL
tT+LOB+NwTRITjdslzB0oX1tZ5XKzvW81bsMOh/5+RKvA2smNipNtzK+ymFioQs+lr8EO9heaTHR
DSH03oHMJ/GUatUEpVLC4g0aAr5UIcu6HHuX+RenrO1hGDauLjzlZqQrsxnPcI/3PR1DlWCrgeKt
v8zVLY8obezTPwLWC23TBGx2FtiGmywK6KRM8aqSf5q83pODF0wKW9FPEhsywrig4+LgNXVOK71n
Kjntp5ECItz/cYKHuuRxcO0/4G9N1uKlDLCpNSxlt1RXMpQB6c81XWH5ZPBQWqsXtMiWX+Cfjd3a
5sdSTs23z+fhh2r/IXCgvnpQoJUQEP8d0HH52BcDUH5LebE4O7gHaypQjY7ESi0ef+mcN9n/dzox
JP1lOmMTxmS35IxK2DAMbdC1Ltx7sDMbPz8cen5fEBSJ2POE7qu1hljPZBYf3Kd5OU529Vl92xwb
rhaxt4FMm9u+q2kYVQA3PHbpglRD0NFjs0tp2W/Ttqv9WJdKir/YZTCBqZLpXcz0ssvdknVfAs4O
jYKg8oFbCRdMKdhkDhqAx4SnNNlESPL+2bqRpzy5fGqxUsoZYS04hODOz7ff++RndZPMJztqBxTl
iqYTt69f/1df/Mbe3bKqC025VnKSXH/euYbCzOV4DdL9uiB/nd5dC9QdGFJhrCE5bpc86Mi3Tpl7
Kvd+xpPYdmC1Mi8D2rv1dYMw46hPTUg0Mc5eFzSsyRwQaOB7oUqolKkLWsdRG+zjdSxN+u06rQSD
JyDjtNjNuTJVeQFtadFV90fdJaxz2iNIm+i7cAbbY9MvCWAJF4smwVLlXWuaRgiwTKU7xH9W8OmS
7Vz15teZ1IqpFgoev6qGnGCJs5928ztNPTErau7Tas6MYmRu0usE+hQ3vk3gcdWJujGsj2DoNNbC
4XS7fABj7KtJvGcp/EptcdcnYupSEg0y8IDfbhwem5VDShHE7Li8Tr1JqE9HSzKDWu0hpP67TO0G
H09rI48/e0vlf/ZasEd3QrkhHKT5NdiTNWocD7TE1pbVKokARSbxX5ShGxL/bAQ/j8o05VUey3Zi
ASr7jzpg5yqeSz3FkgzA/ewz/CfDmxBzJcQh9xlIhcBstQgyke3eveCX3uHnSNpBh/ShJiXAQ4vj
c18CAVCa8y2hBFOu2lB5cIVh7BBPjAQfylM1qEsVj8Zb3WnjRO2BlMzQ4D68YV1qMG2Z9nZI5JW7
THOLMA9oENpXsTjRjK625+bmSa6fT0W35LcqYrWFN9UpMtR3IH2AjoH4U+kLrcmEIlLu15X3yaL9
stLgkdAVjlC5XJE4NCpdBSP+1S+XMwuoRp+RvFQ/xTxWj7GmeJfp3KPvw7cbKqaO+etL+kfolSbG
ChxSLI83oGbVFGeDovYIvKGwDX6EznynLVU/Y/FdwPq8xwLYq+ppuObbQRS9WI2kuUtvTilhrRGr
fEJF1orXZNvo38ep4N5AjARVSu1sK0SeIv7xTtubf1ouBN+O1mdht1oWIX4M2wzZn0yQrrshSb+R
djZkM1dcptK1CNMMfCS4zN4cC+0l/xYzUORiT5xNwTOJymDwhrcsGjOCnjB2pWrK1KuqzJyn9RxF
L1wf/Neqy4jT9PwUWeUie6jz1H+boNLHHZ8UiOWSpiTHZMy+kqo6WSpK5MxMlCqUKUYQATFW5N2T
m8YTX63JIDECmwTglYbsNEbcCYfyBoi9oA7oS0c5Uy5qjaacbSo9gzQFIJDfmcDA1iuJ1H1yUog7
qTR4hM3Nqd+s39MRfsITxuGtLUNCqUbNly2Wmtc2AoCUfrHq5gcl2fQ0JgASPhHXd8c3QmDsvu4D
mDZ9FviCOy5rewaod9OKVBQmTWsPxqNHEHw6PHc3o1mFTQ7lb1RongPl8iNUsUkiwq22K27vayay
96+HXwLgcD8YK892TLNYpDOpANz71d/OSHaZ9h7698xR3QXBkb5/WExQ1iKOwJl6lnSHOg64HP2i
3F3/ZJsNKfcCP9Re5gTEjP9MaqRrXL3MiHovm8sSbnafJOd7aSonWZZsH29d7tLomzOLr1vNs8VQ
F8ci8tBH3w04kjhfpfsJsAoxxwuaiBmRDKA4cu2sNHWCVyUBSVNEEfz4hYyXhXmnu9bjgvQ9qfkM
cO/C4cecnC8QAjYa45NRrPArCPRgdzcw6QVTl7gOgKoJ2Sf11AnVQkPDCHTNhaIX0uQcml7SUTiM
D4aiPsz9v6/QnsMedKaXBNNXxeXLSoctcBQpDQtjyUUOSbKJvmIDkLSqjcXmsznALh5CDuRNkvsb
8AFj3pzb+2dpZRSd6dkQCjZyfhKy7eV1wtxjYqN37rs8PQjS+cqMM2tB7m22iOZYV1xqRcdrnX6M
DmmabtbdIgJJ1HusYrb6YsEE4NyoacP2P/mhy4uMWcGGzZBl1xbOHgQNTO7lP/3cThjmAIuN2WFI
Bq74+5g6SISkaG/TkaS6BxvZ6/Std6UHN6js2+un79eNVMSUbu0F1x0dpbuUFJlT6tD+EAA1mk+k
lxLoLYwPAujgFvv5OWlNAlXk5vzAsYQ8vo/XaFcRHVv5FUJ93bZ89lCMxJ0IRpg3rQl+yHCgW2+M
MAb5WMKDhfvnYX2y+At/b47ldIytsnf6D91LEMqGD/9NC5O0wzlJfRp5D4SBwFLg9Q4kAqydvz0h
pLQqPdhhupdPqanjLYs3CGnz04Qp/WSWWu+lNzhGx8jV5NSOCbYJjhUjR3WGVcdpBmC7n1Hy0ue8
JsNcs+bsUf82I6BKliJhJnNi+fnpHJ54ArcW8GlX7PotsvhqiV4BdB+yn1Z77SdhwT+aqTaTJ/WU
bMsbDceoNfBYq+KEgGI0uXhs0vZ3AO4JhnRPIGmoKZErirIUB4AgQt7fknQjhaUm6N4+hSE4b8Bw
maGajvqKJ9F0KD/05QAwwEgQnQ/oKWqkBNt+JwNTeLgi7HUyk/nHnO4vQ4EkSZfR0B+D+1udeKTv
82obbdCdjrvPybO3ddqnpSxZ2ddKuAO1vkbUd98J5ZDu7lPqRzlwF3E6n2OKlpnKZKyQJMmEXAW5
vz5dZx7GLeitSaLcEFsIsCUPO7VQIzyQkwSPTUbRoTmmEoOpusYgm33/PS69bJZ3qioxJ/VX960J
Lo/Hm95E9q40VX8hO2+oRTlEbchLSDCDrRjnGSqVZUfZZaTLzF5dIQF1NdmTpkv7ylIk/Dq8nPKJ
Yck5Lbl6+UToybtsZGBwY576Xkpoy23uBH9Frkwfa7jXBmUAbAvrag7TEFgZxpRJopRBYdHRmVha
AHegm9T9RS0dlSkyFLx1vaxZSaUejpiMIexBmTm9jdtvtnP7UMQGDQkvfz6hB0PIdKgN7we9BK1t
dDrWukLX4Gy4dpO8CcaD4o15600ezEvErKmpdbqg3DoFgKol+NEbZQbNW2xVSm6VrZbPvrzZTPwq
QJCcO+jDLL1M18tWR4n5nS0gg/Sq3ZiaLfm/3iJ0Jj51zs63KrAvFkmKEvCOA2pqTP/PmB3KkY85
1LrPl05jFF8yzy/iNCySmbO1FTVVIN0Xo7vR87O2/BX2/qgc7suN3Nc5jHMz8m13XrgyhxEegJOy
OgfC2QvnvJ2v6B13pjshY4fIxPVExHbmGh1yb8BaaZpaQfklaWy50oZmb1sIiXjkG1wxedTdyqfR
73G2P4hyhWrpY4HlisSFG4vx1sCElaJR+P91Rkcbke99may1PbxIdEwYl3S8q+3W7/og7+C5+azV
ESLWCWMYCmGb2qHn3UHVKMcEukABuq2E/Xa3QbyOVlbxEyuEpWqNrwGSN72MVx4FvPDhXHxBRxew
TOVxZ0zUn47S8bmfFWSacfo4zizxL3n2msRPxQemfUB+QduTT+lmLKhJLzznSl4yxZ2FNp5qpsQ1
Om7Wlhz5aql1LotA2BmkNc4Tp9Tfl0tf40mloKf/EoJScKF8jVnaLPNP/+f7KFBEPVOGJVQP9u/0
SP1aCcNtEzWaDiMS5MIcRqCx7nQx/HLhnKetSttwZ1KM5loQVM1NSy7Vb6VGM7peuEmrc+Dfrf4M
uZtE8uNu4fGJwvAzt+u1U7NP4ipvXQUgHamyaMw6fJWmV1LYRMs7E3IngGQP5yBf1fU4zrzS1l/i
TpbT4qBlj+XqFj21yzdB06J2PwfqluaEIVPybEfWG1/LNjVWT7+mIADubE1S3E+Vh+yM7fyLPjrS
QgvjqMjcvZ5qWbrBSi2LWJyoJtefCx6JYIHVPxF5Q8o3k2OHFT8GjScb3Cgh+QYmiYp5oCpFA3H7
u/8zKJEYVJ5FLmIhOhx1Da1ETaFuvBlu6KZOKG5yby66z9dTcmp7ms2WDoBPCYYefCBwAKzXyQ3d
AO1QPws3SMU4tI/wUfzjM3lFsCmzx6OMn/aWDKM+6me1QRJWXnZ541asOALNvy/IRXHF6fwyLaN9
dYCTz5jPEuzMSZY8caIiwmtXAjnegfejYG6ZCm7T3rOV38SvUqrO6J9eSYnUV3jVi2WUu35ougw8
wZXeBSOmrzTopZkr1bIb/I8YXMaKmwUDTaOtR3CP9+La+vGHGfpp4aMOoTAWg2ofOLyzuXWv1uQw
KdKNktHfRlr72O1HaQ/9jdZLgUSEXYXubWT5Lg5El6QxDb+eVLz/iXvgJ5u6BCXNQGkHkHq480q+
XNFpZ6gDUMzQbDDYRVgSDOr7GdOZMamnhSjTTD3CMe2UN687amB9XJcAB2mO1cI1LuSjvESMkflJ
IAtLxlWGogJJr9k8WjoeWd9YxDk6HQ5YLipvyyKGhv3ljBrZh8Zpr460jFvpGEeKn949Mj1qXfeA
5qu2KjKFV+afhBiHErN+DcMXmbhcEsWV4Ui2C/sPkGe+0fsu64OxfsES/OlUW8pYtROB1Uwssd2h
zjOnSuPIP71gRGlgoNcf9BgTNRHxT3dnUssrXE5PrBxP/pfrhWkNi542ut6qoKlYEb9gcQuu7fFY
lpNBdXpHgfauMJ44NEDZn32z0oQbnPFAdlRJ+P8781JhZjEXac8vXqmZXNvd5k0DH/M0VoJRBJYd
P/RU6mltVuBHTy8mwr8/oQnbFJfAwWebYAkcrRNG0G9hyJOKWz5/WGbPSq95xLr7cEnT0VndufA1
Y2EqhX1FH80qoxue5BKNRu7nXn9mQKOE1WzKuxiHBF/ky/hVgwQi9kosmFkNNhT/8GvEAGNRD9H0
2ULe8oDxT8ZXXH/b60W+Qp9xBypUqlykW4x/JIDWJa3sDS7/IVhLOTELKBzPsjbrIL0Cp37Os07q
ZQELfAiYkeYy7NilXHto3GN0QIf1jyxwiDIRPgDDXO/q6rwFPAO4u4+GG8gAWN5k2fWLD7rYZSqY
+Tju8lLHOneZ41Wz3BMo9VLNCRRmHKizV+ZN0KLC6VdkP4r5fJNP0mwYpmDr1MapZfXifof+6o1z
/UNGcyyMK9RcaTOoh+diydhdnv7/yDL0V87W2qJc3ADSkqvSb4JG6TkRwIKWkX9bqckrQcze5Hks
BN8EXhwvf2CjHv19n1pA9nBZfI7LfkiH15921t/0t55irWRrQd14HGAE0nqsDeGfRQqhjjG3N+5s
8xkh2s3LXBoO61BS81QJEQ4R3RfNMaSs7kph9XN4OtSnfox+qQGPv+cD/x1Ov+3jDW4c3co3f8YE
RoHlNlUGqsfmwahwYApTVI2qe9NHi5oiD8TQNTRUdjFENIG9o6qKHQCayLSiACA4nys+c8ZCcOF2
SPDdDrkpsUgZIQqcNQAuv1pDBH1K/i/bZWpDGQBCOqzik3JsHKwl1b1q9JimeRvdlqY0oZlgCySo
g/Bx3b6tyAdAHrVi0/NSD+Z0wIl538cPZzE2PBHag6wxjXEwfDI4gDshHUsNAQ0q8R3qfrfXdY+j
1W7SloZ9gExvRNaM8a7QNZboiRxMTkw+D7ZvpiM1PJQV4bkx7+7hB0/HuU8xPkqtXVTT4I+N+9qP
rXy7mIF+EnJevlxWmcdspdKK+iQ+a4K19xNRQwl9G2wMKudiMqZb7UD74kRIYN6vXRtpSkQEJRkP
7rWA5wrwozNDolpP7QnilOQqk0//A7l8zK4/6XQdNJ7SYHWSkIrlvuFjoV55SSAdlSwrPh/tPoZg
dEamm/Xd2cWsa74GbFeEAge/uiWs03UMan1p+V7egWHxnZui+Cq3Gn1gpFmZSVduNahqXilM1mrt
0+v/JQgb3VhmAvHIdzpkR5XwajwvYCEJbjPwIwikE4PkUYm7Y30crFwCArQgED6YPCoCLP7r86le
zZhIexUYvZ/y570nrcsX6CTzHmOu71h+T0fxK2E6gWig8ySiE0gnh3FWaAmrxpSkY0YTvYyHKUKH
781Vj/9Y5OZlme/x766jl0Woh74M1AmTpknuICWj/T2hfUw5QQTNzSDpF252kFgQN6KA892HkVA6
Pyt5v/14boxPilA4ONM5v3rpv7kZqRGmWZZ2Nk6V9jntN5+QVMx9VRIbwdb6rS/bHnjU3hRgb443
LEk2HZeomiQJIH9d0zmatHcDiiX3/UfEVfA7NzW/C7fckMfwb2qaaLmP+G8Kw0Z5z6pZIR6wINaZ
Mec145v36dvJOPOOC69wHusiUII5YDkwyGeqKDPUXZ0H/9/1Vy2pua2I0w1co6TqAJUXpyc9vOqQ
rV0ckqPL7Ctv5n9bDFOsXhgjSI+WBV4sLHR1vK8tJ+7EbPsvuILJNFq9qz3EFj3iyfTSr99YE5kq
NJpcXcY2ezo9YaQ+vqGOTme9bj6zvH0S97RyNK8lIkGdwHg7+khNjAnWk3Vip5eEvkbiNnRbP/Jk
qKVCHlx7blChkRm/jcR1IxHpYG6/vf8EAieYIhh0D2HIZklB/UWuxhFmZSLnuTBLIvf6yq5sz1Dv
3mhZgDzyUTqcIn/FgkDEbyfU0qW/3wdS9MPnxVTrqdPoTVpCt9dzpoeBYzZjblo2fW8UY0Y4kGxl
IkOdseYEJULXV/fnCzODhYnMlWO/NaF1XAZv3JzP8y01bdTZF7GZAOrzQf61iHzfzomBy5rFXuMX
TFwOfz5cZ2Oqdom17c+BBVBD4T926gsN/nAQT1ba0yF0ZSepJ4bhCB7OB/vSsqjm4bkODNQG2yet
BOabSpOm1opvvkxZ+RGTYYOkVwg5wMLA/R6iG4OvVJKKt58gM51n6qUnlIE4vQKrltXcL8P4ZQzy
9E/C3R7JmvvMrNX3HJbFTjcGdfqZo9R2VaUR0xXBK3aUIugN+qwA+5o2RjdP/6xRblbsfR+2q+mx
iD+y2CYe9zJUvtf5EgtJxK3gdB9V2iazcgCCfkQmQSxvdTpmnaEUQ78lxEQA/tNlR2ZtHjhgPGBW
qSOSbb455orbpx3vztLbISXYA5BlpQSwWKw5NPmjVi6M9oSIvhr/bnLmyGRuRXlZsAiCsHPdiyjt
DieUuB+NnO2m0zccE0Z1IZeakEDgMfqUyWKdxnExHpIds9bfUNUb/OrCrOsy/EIYl2L+1Vp3gjIZ
0JdUp0wJBdG+x0lJ6+u6bDHIU4nXKi5GW/vs0C4OZtEMcl1J8VBvVxPVomh74MzWaQOXfksl7aNL
cBLu0A+Ky+xixh4pequZLPdT/pCMhgyr6YFjVTazr7b0l1wwGyyTSJXWJ13j9QYsb+GBcye0ZrkK
8Vw9JYTCpYOtqI6FnlQBigC8fL+y95EsBUB8qhkhBBEy6Zq0UK4u8oUiH5kEI5xkkAS0YhCJy2qT
6RhFH4tyPoMp7auLmGVB3N1YB2A6e68Uq6UcHt2KuguvBJIiblt+8XvQ0niySteNtiIbySU869W4
vkmiwhd6To59nhWOf3Lmovnd6ih+kJgFJRN+K3DDyV6iao8ghq9IzHTAEuXWgCsDjjxZQHNtpAYj
8huCjU97y0xPAc9RNL2OwCtM0iDZgFWtTg4krq+PztcXyZ9YqmkZ8kUK9SYtjA9xqU+j9Gj9sxbk
t/Un55BIFIUa35bVKD0BlplnR3aJ4FCSxzJXUCpjUccXn0xas9+eZE6NhZmn0cTVcbJUpFe6rhp4
l4A72q8JtBHwi5LE95OwvuBKBLcuDzuBrK94OsYqKYprjGJWMytf+EDH0XOhjdyc37/sQGWrOHLp
b8JCiik4KvxWKvmZ06/lmlKO9OvR16V9QA5lKnCF9xTdgJgg35vcIRmycwcc6fpz2vcGoe9a5ZxR
HbxNB3GeOssOxf33pi0SEZ05dBWblqQ08lAEbkh2nQReo5EdJDBum+NByBmQ0TnUVBbooBtTVUoE
ESsWbM8IhxTU/rGEARJguumnXJNISo+CKYiyYqb/8fdaZtyilSdJ4d28uFTavMkYXCw+yVNCZzCb
U1z+JdVM2vsfMxEgR0qG5Iup7HL4sCDh2fLH1o4s5XnBgsr9w55hZ2XC+tLclbxFa27BpC02KOaG
eKhFQkQsMdVlc97RaEXwsv/RjDxqpPHU/1R48LZv/JitFVqFgwU8Mfi4w2aSaHLFL0vTVTfgPMNU
z42RJyt3HTLxxxG1fDLd3CWXFayFISk2XXJphZybq7xqeXlG1hQ84EemSvkW07m9moJamoafDAdk
+iX8fAKYX5gWw3EPmTidg+ZMLDfW16UNgRKwF7x9iYtjMJ8PMwjY/0RIRKMzyn4QIw6XKJnUd9WO
0LJqTXBPIRfv4lPa0oZ5XYKSb/nyhTBs9X0lgQdr5QDugNyiKyPdhIDpFSY1Lv1Ta7i4rvr4yVXg
RGsRB3yV2vFmmgR3APFElBkxEy0Yw0wlBBNRge1s/2wbpGQvOsxNsLYgM3gsYNrQ+NBAv4mKqs+x
6nQD1JKeXcsjW2I1+Ifdx8r3p9IemPl2X5sKkZqN6hDakrdea7FfrrgoeOoqx3tLmYL1QTvM5D+2
J0lO8EHgGFPzQWM6CttLfZjQVyj3TRPVJXJDvpvwYIfD3tJj7O9MCgJaMBfpNU8yVAMfHG9hEh6f
WMfCyLgnmLdhQ5b9nedKgslxE3ppoXC6sWH/NqkjX9FfiBZ3F8jt7Ei8JBXMFbqcFLmduVlzH0Ng
WB3SZoz6huo+fHpkXifTQgQCkKuqwSriKVGmTIqWb//p3iZGJNvdEanpCOQm4NLALm6gvNX9K4N+
/jt2FtC7y3wmcKactxNzaVINt43Fv4JNBx59yuUGNqGAPbsPj5xEkeKmocmBlYsJx/hotZIP9ssZ
z0TgOuMlhysL3nsCGGZDG47KR8vVZ1yrgmbAvzBgT+Ai9MdtNNZI4RU4J6d0hkXMkDJo9OxqS+DZ
SHK5eAMl25fgL+5rP9Oj3ZbHCUtKgRav9PDvfNAbZ5sA+5hQyGtGAGknUCs6+lfD0QE71iV/IFBy
HgJ/m8MpGCJsSUWpop1fdnIztfU0ly2qFXaGC6HzpCGhjJM74N0LOmg24Q7pTfZIp3iZZ3gzdR7m
QGnv9w6UMp8ZxDKlrfe9EmQNHUiV+su9BwW7jOLxLxEbilYSZ8ZbUUPM4jdQbidYb86han7dw1lS
QylgJgeKrP+RugAi+a28Cb/y02nwldlJdHbw4cn8JTfQBFFr8pDZK8Z9JhfnEOC9xe5frx5UMSKB
whmjbxt0/wv4hNk/CMJTEd67jxL5agVSus21XckXs+EIrqsPRVt8HNDrTHb1a1ZYmRlVveLWSfSg
HNH5VIW0wU+HrTsmK36U6hVUW4csYZY54CvOU4Mo9VypuFW5kp+EZ8Hfjp0Yi/5VdNsoEEqyG5Cf
csnZFpHEb6pQ6Bs9Ybh9UEYvzqDMlq6jKAuFpJzgMpyzepUc5zmCSNLAEDcuF/uyDuBthKO3BMTJ
ZUwGJi3Kh/OTCDRi6UvJSsrgQAgvUY+93+S/43VFy0sQOTQDQy7wU1DkuCgF91jHFZqi6t4+ED7R
ceLzj4UE24/JZ1kZ613HnHwtDRwEF7Pvl2rdKHh4pOs9QLWU4K32kFgegMr54GIQrBu4/VgejBuG
Gnmsp2YU9IO3CnFZmBfHHlmqcQek7F62Ok3j/wz0dJwxwx4MazDdHJoWwMLtynAz2/9jYC4YwATB
c28Qgb2Vb9ElRu8wcQflLz1wrn6TUr2r2ts/YN9Ud+TQhCZIIC54PoXRud0wMvNx2I2wUHqywBaQ
w6MJ7djifI08V/kfdgl5AfZwXMOjsWbrL2tWa5xmBp5Z5Fm2S8Dn1RddxNfHE/QwbVTo+BHTRs/j
kLLKBh5bko3rDAR3ZRZzeonecNhDv4D07NgRYel1uPgpzvdF+H+ArVrcDe2t+NV3bFhTBFUJEB3y
aYnT1fYzbZUjUSM3H0HGNe5Jkf29TkMq/r4jAapHSfcw55sboy/kDJBx/FuTMAfzDscP0zpj+Wuy
FiwO4EVsRujTkk+JscXubHpO50jwJo4YsBTy5GjlAYMdKbBlQNqXNy1hRvk5bGuQUKRtNgMccfKt
ZSL34EZoelAg8SzxOL5RNVCh3BbEH77ozYCnVNji9YPwtMJiLWXkjoX0VMuqK7Mk7s/nRN/0DyGn
ou1ve9Eu4zf6cBH/azWn+wBIonb4hFI7UNrM1UBagHUwLu+q38/535subfCuvjPt3u7rBdP0qhz6
zUxLs0vkXYdp427YcLzk/c8x30tS9iDWLzF0NOlhD8+ku68/nHBSEt5aZyaBvE6spHo94aqW3T/z
JXXzRAv1T2AqbGaDzQuZi8Li6oWjR2I0oeUyDmNz3lzlAJYRpIEXLMSt2EIpvpmELyweeYVKYnDF
RBVRk/jJXUv1K1wQ8Lru+GCPnLklgNs6uaUvhkCngGwAhUnxOmFFRW0OFReIVRJ6bM56ja2K1aq/
fMkjlgInvOUfvt4jfXc3a5wnYwjXIiqOcasHqvp3fFaLdlb4o0Bxzgh6oC9DzQ9PaDQoIrCBLEJH
q2YS7IQfdz4bgokXlq8pc14C1SxRmTb74RNxcHux4W26a2LPmwBLdPIJCA5DkI2PYKjjDyoHvGBD
rmNeI+tX16+LEfQUCYujDFJ/MheYnSlVfsvKM/GPr2C2ssM6Q4Er58jcIhuNosh5Cjd6cUljikQS
CN/OPkKExx2Kdgbt3YXYAgOtoWpXqIJ76d8f4LNh81+YvA4M2hHUF4OvT2bJIDwLndzItX+XIdsB
hEKNJIg16Y6xct4CofNzEMyMgD9cUfwjvw3tWsarts88lCasesx7AvDQVeC7Qf0I521yprTmFGvZ
lqVqhwnFsCjkL94oim+yEVByuhT29MMa0gP72rnz7H497aSQMgZg7DPh0uesSTlu11xuOyv1D4Oa
njKs737tQoqQcQND5xiMcweMyiVSBozb/OCgu+4JWaMVBu1dAucVDvi5PG/oo3Gmr+J3LbwNFnGV
5E8CyeOcKN8hn69c+xpuwcjXcm3rrQaLJnoQzCmy1CNJuqO7QqpBUn/pbFm31Z40c3TvtKYiCc7Q
JcxmWgxgPRP517G1FC6eOMYPdVS7nOqZqSYMuK2/G94CTZVzrWR1XcluFtf3IUesur2y01Gj7pfE
NDmWfFiIgxLRKd3EvGnLVQawIlsRX9qxCWEfabmqhZkmUetY91MZX+MNPOB+YetSJ9Sz6JRaW4TI
ZS9AXxo3uC7ARfarMGP0dZ+oOGJZsW7vPb3fFsjdvQy4DN7qnRVj+L5WkNRIT1w+60wWFDR+QIVQ
hYwEbGx1m640MJ0lgqku3aOHvjcSKwSfc+EnAz+ZSOmqYA+jr1sc8Yaw6b6N2sk3S+Vvf2tJxaD4
6Op5EoFYNP46WuSS7nLUgdwWBKvqZmtCHyn6Alqleqm9vc+GJ+fveXIGQaswcde7WKN2lEXQ3D62
KoyNisttvup8SwysNdB80rZyeBLs9yUhRpCUuqHjiMpc2nhmtRpoXNiIOZMQ0CM1y3SbyDO5Jg94
eZqTloJEmgUpCiHCbLOLWCobwAxmvjcr5FnZ5wpK6lFb4vl7dqmpE+QBQoMmJbj+Hx4LGtmQZYCT
+YHCN/GTDnk8/fQ4S/itD3yR37gVm1gIgPnSH/ILbgfCpupU0QNn3XlsYx1GACVC/alIhAmeA95H
ykYAUo5tf6JEQnDU6fYHcS1n0ikHZw0h6Nnc1YoIblt+W0cvybFZgsX84aTGCv7rFOMD/fjD8Pcm
UZf5eQJdjWVQiIkhTbPbCx6qbXMVKLtrCC9TBLDUP0x3ekOClBIWL45nvClKrKMbgbAWVrMlLWDq
JgujO4B091JChlEkX9MharH9oc7eSn7/H0S54juuTKWOpSvlETYK4LoL4xUrom67DcCGlttBlwQV
fwyBwmroJFqlnFntZfKCK+3DoZOM8FQ3ubQKvwkmoe0STEhAIZrGtxOUIY4sqq9k/N9yOfe7+L0j
Dx+Wz0M0rvd0K8BGzEciuervq8SBhHTB/GmlCrkE9yR42rqfts2PF+uPOLJJRFofpRGoc7npbPEy
JF35bYyQPSCEGeB42qzq6in2PnrvAb470/v8LBQWD0pCRYECeITAf4Vf2zZrWKnDWT11kDf+H8b2
fL5XpU/AcfO10zz0u0zIW2SXepQlvWE5v6CuvZ/MnTYr1XTWIm8P5pN6DU80hqhTvsJCbjaBc8ei
NxmizYNoXzyD8V8HVlFq35R5osTxZCgivhoPAsbaU2Xm3SE/CNGBnDD1vp7aqnKTAXrFJgaDwBmn
eQnkelg7XzvTMD/9FH6fdD5jlD/t4kVvIJ4lS7659m8PiWGft0E8/dz7t6TjvwIcs2QiaUpB1Uw2
/YjV1LGqnuDFcp2VlBFu6U4lY6owQpo9B4YkRJvbR4W/L0Ahg2Nutq8jUAplXPcDW3exRb6S5m7G
ChAkKYUx5zxMISHfLZnv6xnpohL0ngyGSyQY78agQQYSR5lxNEmcgymIa5l+eDWsi1plbuL71GQX
XZGnYC02Lz5m5M6a7KI+2oyoV+ex4b+r0n8LgazayDBCJgT0m0M+nOuUHKloGQqhU0PqonAOTCOv
9Tm3Dh1QZLxBmAJmDswYVf8OcgBVtTXupe/Ovta9sbmUabiXbNwPIjjxwIahcIYf32rErCWyccMp
r47m2MfFdveAu0li0X2LQ+BjZtyCKS76AWUO0RY8xFi3dLYlP8vDR8Jon2wMVhgO8sl4LT84vET6
PEMH0vvOBxkWQmqldhTwcW6KvHRyIPmrygDlOv2ARmpNOyNHJj7M1vxm85PzNNrLKIwgts1IpbIs
KztE36LjSU49jlGEgiUiZIH8cfxiXNbXnLL7mJq+aDeBomix2MQ5AZaEhuVP2+HUGNBc21fG5p6Y
ySyhRYTDnS4bHZcIutn0LD9nV+k1crH+VSO5Odkwatp4MCtapiFFZwhTuQfvH33LQehl7hpTGuE5
HKe4WgmeD8peERW7obWWc5dHQwwOhoHDmcgkK3xFSfd6k5ttnwXUdWA6kgf10LSj+mHtjKoNSTYq
E93tm0UGSUc9Yc5f0M4474fbX8AU2d5prc6jIcgnVYF5OveZMzITRSXsm8Tlai06PYhQtLwLu2bi
JPoHXr3Ugo3qLQ0c/5ro/CNqIUAFDH3JOZYWlI3DysN2Dr9Pj7rUdJTc2GqKQ+63P8KxifwKO1xL
rO9doRlcUu3GCDnTfJDWPMNl/Ir4tpKNx8WdW2YNuSHSCXef5h7gl7Q9ol7dVVAbUmY9Av0ulMhZ
DgZC9kw2fqQ1VFu7pRK530rYXYcfMYkfkxpXhLIjot1JQW+14MUsVaMouCqiQbkyUjcEQZN62MfO
ERh/MvlBX/l5gNHNTevrRbuWlv80hS6v516TJQ05YZQYmHOrpu7pIsh//SDNXHFUxMeFYazAH67c
qNhDueQIbNHwcN/IxGPjz6GhE4T0R2BnaXuKkGOlBA/lnOcoxnOGot1BGdrIFfwWJw285kI1Byz4
tqKzarix18aVLNZJOiw1+J0MpsFSsKKlkjjyyYZ7diZgfMGd8wrm9E/FdS45yPBCNWeHCj2CZOw7
5tik5PVCKV0QXjxflY1CqBLEZymET6lZTPrxdEJ7awoJfms1BEuKN8qlrxT0H1StPHjbNCQLZt6q
xnnFe0AuuXxrKGeYnrsjRwTC7FQokAZg50Qor7zHDuNlok1s41sClDYmtk2iB85jwTbpFvraSETx
XVbh8iDiaajq8efAX4XLfAA+ufbFRwRBMoq9PoL50+zS73sUV3CKnePaROqKnn6hOSsjOsosIL+N
qdVLd6EMrbncnYXZuzFWifOzlbMwAdgUgUk1Fu94LZv4r03EVLllSwE8d8dCMZwzm1cFuMrlPFE7
7kHlGq5Msh58BeIHaTYrGzVig1KnQntNLeFS7Ocz0NxEaCTix56yh5th2N8Gjg61Hz9iiXaMSuAN
v0eGXM+kOdZ5KyGq2il5+b8LieKIHN0hoXdaUhQ40d+E43ONGjg5YqNfElK1Z92HbpDmEgepACje
6o3Ye46gS4xH6funIfUuV2KwJOki90B4UEeKbsTub6Mlm+dvyt8CnXIJAxO53y3R4B8uqMHLb1Gn
FeiHER/rIrwhtXBd1DcibRJU3SRuQihGPxWYHCMNhqj0hffkHXvwcl1X/x/NzIetGE8ufiw305lx
ueUB1NkV2+EW+hIPbSKo2ElPtdQ19CgdvOtA0VFzIRiff9kTMqxr4quDMhX736sMutwwzFUhW71x
VQz761J+jQhcFX5dNdRbBL+3PiOTcdkWgCEwZYvF6AWZSjZUTxOncocKT2pB0CGW+Bos52nuxzio
kPeZukrw7WI/GHgtc8Nnn+jI0uCia1LcXQcY/5blxJ+xbZUxf4OTKSLYcKlCBmyMPKqWk0DdcpEY
03SQBlUXRwaCF5gmN39qKx+ndJNTbXJsBr1Fypz36j3kPEP4inYuoh/oKtw+kpqq80MtszKJfdVW
gcNErpJP040CAUTAV/qhz2vvs3YRcMMTRW6XEWLg4lm9hkeZlRXeWgBLPy+BJF6M0zdPohE0a3LM
JAidyGkjKHbFM99A5owh5YaGJrzjsEG3wrqB5IDO+fRJR5KY5KttoshtpQl6gYmiEN3QCMtGYsE2
1xKcNJXw1pTHAbWsDBlRLrgdBqV3ourm4HKBMxFDZsp7lpNVMszjP7Wei51chZvVtaHb3cqZWlVC
ZIPjLOcjsjePW0xp88CNaGWU1++70B2nwIJpKd4AGElt8kYRtPG5+RGNAfgq+wsVn1Vt3GG0aac5
WnINWs4W93BoOWW9HxtE/q4PKi5GAjYhdx5o9x1G/rhw/OJt7YrHWc36yvOVgZImVqCNCIfLZS0J
J2vmqcm0HfjeqRdWlPEj7si2q45Fx0xkMRj2LnE8RX2qWNH0rghdH0j/ft/1M1h0MMzH1Dc05Ixd
MOzTbxBpYtfDv2qu6hjR5GneQJVQSdbBED6Sxmu3ClIMV/g23JSRC7TFDTzGz41XcuSTrfhLWtJN
i8ZG3xWZQfiOw/i7fopHx+yIco2ArBLbHozYEjr+UtrcvKQNrtpgijUT7Eyd5H8dDe6X0qO7hess
mfpHtRB5dr7P0kmGssILKq+naRVcAVIsgWl4EOMJh+LVOC7rLQLRcmtqge3xQGl0sGMpHJIgjKze
Lr9EgIMwQrLYrkIzmOtPzx5oV6beOAP7e6AZ+nzQn2mROpadl+a49nEZyJ0HLgxputi7Kz/Tr3G6
fejOz0HVpXUXtBiObptjmbnsoaIrmAx8MOqpUKUfFkG9PgSX2FP3n3fdPaBWTLe7wq6ZqQhdYK2v
RpE0e2AcrooBPGRKuf+0d6aKlOenMdKY6/Ei7rogmsHROk/90YoQBJeikZ/wguIHXyq2E2XRs049
V7gFvZjMe2XQK0J5lavRGBGq5+xj5tIt1K7Aw2qyA7SqXPi6VJjL0y65rBhPXpg+goJb/kyHc0+s
Lx7lLMgRQBW/CSVLdEkk+JhUR6YJyKH7kxrWkbKDOnhJbt+thxoFFvvCKcGqd0kyH6JGtLacHHA4
w+8IDZQqzeVkIC/c+km5jrqGSmFJGh9uqFhJeQ1++PKd7XQOhOcbERVjJt9Z5z3dSixw5AyM2JO1
hkxgwxgx7qeXxKuSnlFy6C69CgZbBgy58MTWZJGCGL6t8474Eg6Z76cAU0hrWQb8yoRw5RQ8m31w
xmW9Ih9CuQ0tCOSMSRAklf31qYgEpcQ8gs3grxVMnoDmgy8kIua4sHykW5cXxZyzDEXmLIgMbHhm
+E2ho+FA74bP6zhnIIGhVUCgg20lgdBD69UDfQdNUNGG2iu2rkHB61M7XP89vrrKQnyDFVEzLH/T
k//JGwJc1QPvoslDx0QusWC1Mb+EqF/rJyq5DgTVxJ1U0dCpzDnuxP7Doyb9y1DDbyc64ARCJCDb
fJubhY58q1kWomqBUOYsP/Yn91w8TyXsSBkE772qawaHSMQbbybIjxBeT8d5XRLPJrtMCA2fMZlq
VsrAd7hiY+jjJ4IrtSR7qBj/SGKdbzwbmHNHDRzpLo5TmHr/Wxhhi8HsEIzkziIH/MCaoPkG5zBy
CB5DPAR4QuzhnidaaNXI8H7H9kLxaOyNfwisIwF3A9ijq6vCnlSWI/aQ4legdnE4OigfQYA5TbpO
HalOlZEu/HNraCvnutF4iRhpfhpUjJGKKlQLxK4Y6BWnjhK55MmV5RPRw7Th1I48vzsEWy8yhq93
AdhVt4zobv5unNh6AYkvKBD6HUvLMZqKoCoUCcWhlwCNGlKpukk5nfASk9fEtywbZolVu4CIucMO
9+yt4wYZECWPaxI06eLQx3EGpCkqgFLuO8IQqZFqRoBS4xuZhoVOs3W1A5fpZA6IeVIbEYlrRk0Y
3IywxVS3eyPEirNzrTwWzvB4Mo0+lhfDY6zHQlUkdgaogfogyDMdpywbBg6clD5XUb0A/Fdvayq/
Lx9ezarV6LGJiGLn/2odhdtajXFuotM2wvUxj5/0QjiOtWEEbQyq0eM+NWhZ37WhFyEPasXfmUAk
YuWDgXZY3oU+6grcyYrL0djTWcK3SOEY1yR2ROJ9/Cpw1/H1FuJjNkdhbLJeon3YU7uI58QFlt+o
ItDI8+7VeQm1iuK+DGv/MhNso/AeCpNhGIWZK2LjlaFrKDVF20P6AyBqE4BMJJ+t2DIROPbngVUa
EaiIhdciHeVLxnoFYVJsC09m5bIyOMA1GAP2cB6YLeDo0aZw59qKoHU7ZbUTgbd0MxCjCYxcRK/E
GuGSIGrTI/MpSDaA6UVeu1M+RzXE8csi1qVGuxT99zbT1KNDckFSPVd78otN54uo1kSP/6Kfm+P2
28nePSEtxcclcMZchldLfCfBBsCQi56cuJFCd1C94zJvru01urjfEOq9SRqzSCsdtSRm8bsR9/yT
3GnbJbbREP6Z8FPqP4P8C71jpI0sQjU0jxuSyIu+cXcjLOLfjvk7ZErJ0z3k0QMstkxNNQXnM4Wt
fWxoRb2Y30AWoQZ7J2dIJ0qaOJSWNX4witUyFSxnFdNBpdZlKvrkP93xXeUviaNzhSKCXqfMTBtl
V0VaY4PE9U8vwSTd8FJFV2w4Lj+VempKpDvWBxXhfuUvotYOLP3xlnEOlb5zdBd3S9OWyCFZr9up
2m8TK999sTuitJlPX+Qu94Vck59uAky2k8XcJq5FejnCsxC6yd2KfFuVrFppVe3Gb2C+cHErgTzJ
kvkgm8OQpXUIbS3wZ4hK63LUGji+c5VK7HAYp1wBuoTsEKITuKlysFK1Fsm8QVPf9UCLOvVpI3Tj
Br65w4gE2ZVCCN3HeVf52ozvS/Shfl6hxHJVua0bwad0TIBIMhneE44PBvyd/UnGHpPypu6EaTJW
aqYVwD/XLgmb34a67BU3dHeO4d2003m6BTL+oUqM6cM7v/FBSDguFzmgKwEI4OrjR7u+ZEH4ioCX
1AOEBNnVsb7OL/L1io6cM7jfwGJFpFtVj4NGNjCjAoRzpAxIrADSuchc3+pTFc2Qlw0yEPnQG9EC
YRi8r0Y1f+7JSk9TMMkNiyM5nAYo7jG7xli9v+Ff7QeWV5Xdz08KI/pc4mfIWk4Q7wc4AUe8Dh0T
jJzzEvzZ3LGGOzMcrTEldDmsLStADtGZ6PwwxXvmCz3GyjERIYa2BYfxqbre+TnH/9umqRNXCbns
YHRQ6M+jqXGKlSmD/vGSCwJED0UJVdc2Fk4oLAJlRR9ypvR+PpR6OwHkciydJdDcgzClrdibfFVC
cOmQ2bBZtd5qTiTgSoYOMZyyLBAU62Z7aEGgYhrXIrt6U3xaQAWmhIH0DRPR4NY7RD8bIUZmA+wZ
QQQ4GSIU0hIojAPOlAa0zigkbndP7CnN7Pt/S1C2X4WTgM2f8+dIsAZbyQ61ugPzFkT6iEI0e3pk
0TZvq8FyHOCmTL7kcfYlMfXtQUO/S0YJMsXrllG+GHy37scJ0fIuqAQYplQ2PaHGR4xK1UGjQsGG
15hg+LTGnvoj8w1o+EIDato0s346InmUoUQlXBbt3Z6lFkxjrAih1YqoeVP3OBlDpPtOmWFRhXr4
qKDmPb/qNL8rKwXxyfiLtBnpXcWWlxmhWb412KD/+8QhK7aGvLMHr88fvid6ChjmjVlWbbpO/h+y
1Q9SVXv1lCCFEzRmmo4Ogqbz+FRjq9XsWkPxqvk71YCwhQtuuZbfaD0yHZiD59ZECyAX4+t0Skru
WferPNkKC7Er4N6YppWk/os2tnkuxILC0S3pGuq9aBoypWl+0Rvb+Pg3znBuOfjvds9m/MjRoEDq
drSHg5IvRUmqjrGhJ9Z5+ZESktfDUWz1hQi7uS7Y1zcZ1RCrQRQVVzQT4+fuULmXH0jxkpydZxTF
FhjnV6Wm4y0Py+j/g5vuv1hbhMmRljOrmzoaEVUvF3W4zABoKBC2OwbtE8+0E0WUjaFomUgyJp7i
kYhtaTJL3wYqLAVMQ45YaTiWTeKWIfY/45Y17fB3Hez10PC71s6YhUUXkF15hf3ChBQCB6riXI26
IA3KgHomSGaRX4MqackLuJIPn2GS14Ceh2hh1odGSEBu/SiB1WMRr3Zomif20soD15ay2GDn7fdt
6u/q9HPdANmEGpws9TUHnvi8G8OkDrZSdF44GOFlwMy0O98vlW2HJT6OE+JbhG5akdrlYxcfxrk6
hyorpS1WBEkb1fIxQ6H50P1d/yedXbkyp/epaSdxzORkIzFcil+zU4JA2uO09CXn+uWhdg9nkJHx
qdISGJngaz/FnvNT/WHoWdcyLQuyTHd5sqisSoo66ZtTHDU9I3Y2h7vQyAfeEDEcidu0/Xy1tSJj
qHQ7Unr0qAf+9TKxqQe77LDq2YeDT7oju3BcKbDxeKq23TUTf2DKuSjBVxuPXPvi/pMOKvNHxX8g
XRd7Ckao+DMRFUaI+o8DIDVL0pA8VgBOhYqx2M1Rlx5BQ+9QSeFJhpHtDxtm298xzFTJ1CUscwC/
BDBtpYmZrwB0FEihStcA6L5JmP9hdchu9chdrwno9XtfKZrAzpjEOppgAZVH2rrKkDMJM+oZW7Uq
57+TIqHkZCCUkTwndAyCiJXe6d9s//fARP2vt6zK8o1ZXlSgA0s4m7cb/cmoneDcX2jdQcX0iY/0
EsgS4wP4H7C1JfgQpEX5GWdUsbSwZypILySZ5qOFl/fsqL/lgz41PaRDHOVF/Aow44K3/o9+x+Xv
yBpxmn1VzuSuISt6PtnAbJ0yDsM60KzrPY9zt+2sy+IH0Ax1dVEc5kCA7GfJaLWmnAB9qKOi3VAh
jqg30MY8QA1Q/s4zOqCl136hXWh3O2IZW2OChn8eyIYafUE86SVpj8ck6VW3DBbQj7cjN4F7qCB4
h4pwEAdS9wRbq7IUo9zCpFPPrSB4Q5apapkB/dzH0mto0c6j1Y9IMmlXRzIt/3tIqSh9UV6SxN3L
QdD+x8XFaNeiWi70gX+6rqv7uE1ay7wmZ/GXBUi74zhpQXcpYyfrTOY+ep12XachDgI6i1cIVUe8
OLbbj4zuiOQse2HdUizD4J/bVcUGvbf/yFx6ux7PrajBP/FqXE7ErnHMAhbonzf34V6eY0xIUGqT
SYm8G3k8qcn5b2+v0cR3BjBoWPIns0iUonXDn+mVXKW58Ez9BORx2vXYxyoDhc+3tiaaFQB5Bfod
sOfzWuGySCdY3hIcZj98HWZunld34Z6PG9DoHpc3z+bKuBF5nk83T6xKg0wvXUhRNfvAaSMMfGI9
0YQ7aJmR2oNj4yCWiVoaUn5+oz/nB9Tr8SUWK/aGRM/Mf588+csgdva9KdCw6oI2/YwHJpxtAnVn
O+AhSqspacpx9tqsuthbfqppbfRtjkTk8KHvUDON8lXqcuvEHgpLGqXtk1XhCavz5LU6ETPQKj2h
PBiOYXjaH+lJFRt0kyR8C0t9V/b4cFQGi9wKJCDfRuBXd0F7/1ErSQVSFTMXHQYJk4aBPs62mWUo
vgEhEfXrZ2EMMHS5oAtoJofbVOWX3ij7T8szosAbfyexn4FMiLYA+Kwvy+IqIoR4Cz9QPhFrYtHa
W29zrf14aq/kCBq/24MxPpTGRlPsTAKJoseU0eXy0oPCLLpkx4czDJzU4qfjqhDcRliWux7I7wnr
cqGhB75KYLX+rKBz4B8Fn4gvQODI6c9hI0QlBvwOeCOsetHMJTIHPckRzsnX/uOzENsc9/9IL7Zi
cz+wTyWsXB8q4x6YeFV0fbVCqN+/zqS9HTA6FvGaaiUTN+n1DoSfY2oigH5oMLdGxs2OIBAnAouJ
WANMnJspto1xzBCiRQhJng5wgRgwKymvCNzXDkHP8pWtY/BOwbWiEC6icbzgv4B3xbLpTe4DwX3o
o6WeNnh8OH23hW/0ZHxWdV6ibjPgUrLqZBKrnhS4oGCOuwyu3VD/AYda7Ib1LKmOMpylkVrZu7Hq
fYwd6OUNLsh2cIkTmFNb7P8SRpgdmWwFwh5CVeU6ZdemQye5PjrW4WWHZTxG3Tvu5XM9Ir/WsSyR
gkUHc1TE+XrRpZf6EpUWz99+dUkGHBqBSD4Yfa+YSz7d37b4fDawLCEW104chiNMSE5KO9Rsacme
0VQLca3T6SKVgPNSaXhXlfhpZPSDoJhqdzp7ZRjaR+bUNtwp293WP1DBtD786pE1QgiSqR6p4v7O
NsXntgdyTqQ3TplN9baZGmT6w9YBY7YIDS61obr8ksqrA8D22FA84eeF+VaY5S1lE3+eEA3dmhON
1CsD5Y5fzxoi3UWkySF848PvoyTtPA/JR1n9J88dMtT86CGkHGUztMhXrifEGAbg+uFEXgthcgLX
Lbj6nTOVpckIlNztSgI56WqUNCXW0Ah6E5rgIw+hZnxfpLkAM9cofv6Xu4YRegtgg123/cwKROZM
ZWFpDdAXED2sJwqsI/j9kgZHln0cRYcwFgQsw4JPwnl6vEsPOeSC+R62vFlyzh+q7jZHGmcbuW3U
3xjRuN5v0n1CZOH3aDVa/abiE4wuAD0QNJ6dfqlRJgWeQn7Age8cLjV6wLGlvYQBubPYZco6qtfL
8jxipYw/VfakY53B5tKyLIVM/yl6qjv3dXAcURM7tJJzDhPFby8r8ejKPNRyqLozvq/3ZJtDc+aJ
/fQy7oM4f8cDPFvKivmIbJJIT3VeqnGVvY668fn8JN2/29x9UlQuoScft88HfG8q9H2KaUjC9esx
Kuc3IG8rO5D2JrPi8qda4Iboa2gq8NhbW2QAOsNm0F+H7JiqZ/Ghj/oQk0BBiH6KEB5mZ/K0NaH9
iTNF5ym/yu8PLMm0QTKDABZKYYvW16EAaYSTcKRcXWIMTCOmRqmk3RFLfFVR3jJdr6CGUWdO9Tdr
HL7KRdsnUyrli8jPN3XibgUxT6horOYlUTOsQMXG22HLmsaARuIVeQ0ov5qnTYyAt/LBdF0hif5z
DjOAYzfBgBPTlgDEvxm48MIMZ2AYqj5E3cXOP7sbRmkEjapSOyXfgEHYt6EApVecS+dS8Esz/txD
RQt6FrfXYyocuU9L1tdhLTyoLhiNGeXatNUt7Bvb0CUKObF0mXyOorE9Pc97u+ljcea528zxHvo5
cygVR909iawzftso8aS+Q4xYv4Psrxl+fyy5gZwihh2ponS0AVOylMggmUOd7rfYQsPRtCYF2vpe
yCqwCKcT6emW2i+i2ZbrLCDQMZFQ0H63V9s6GPGLzCskMT9mvF+AObpg2W4FxhcW/7t/vJqM/1TA
zFMe0D0nKr1S3OxOiN1JdNm5FmjqUK/QatemasCezalTN5fR1W6jLw/9l0fblHvvVg2Yz5Ua4BXu
26WlaPzzJ4SWsxhlxnM2A9OM2J/P9iK0fEPq3mnq5wR/aXUOB8wSucLSe+E9wV2VunT+xeCEDSRZ
fLuh+p4YKm1koUp7lhBeW+92bGJC6l5a8hUxMAw34OVGgUlJ1kfdAvz00/fszCwJ6Oll1dBrtvr4
Pl6ctRJFu7I0UsJQadjjmoIjUDsh/pDw8zv4GajDaCdJyT4MD4M2Sk+B85t13qF9hpMnbn89GfC6
S2YU9FaXejZLbBa+CuMZb8YWOseL/7EidKwuAoLj16GFWiqtOPg+gvdsoKEiuj6dcE6pwmLBOUh6
BKDWEoth28QfwY+I/rRXNlHMLXkktcyVSU9+5/A6GJnbLDcs0drGfyoTCRPTb08aAxalPXBMvGOH
g/SKSDSjxTNQWBDumkGrfyHMfwjIxqNd50o4JDckTsbsqjGBE3FNtZCwrdzcA0FWhRu9xlBUhDx7
u5HNOVlclL5ZUXg/u5GUKA6Q31cO0+DvlUPOsRl/mr/dmLFq0RTcbQSUMIwN8oaqVJc4ToKmzvqx
axArg3Q4SELO4V7E7gRUWkjyuhapHC3iRXuTXGhN3FudhISLKcRIPaM82rX6GJdnOtxExVb5SLb2
7jvXdCQC6JoB0DDZBaMf7Umm0SKzfxvUGoZsrzwENMM6wtspQv9u0Spk7QfoPPz/QkEu/AyBW5cB
oFow/4YzqhPDYCBjR0ckgulNox0kfGMvqMErfkimWLgYvFLzJVoAe0G48kSOKYcZ1b+1LFUiftsg
2osHYvjGLrl4/ZV60XDif4uv+W8huFzo1tlmuZYgTv0QbcRQA4/01aDNfnnHCYiq34e8u5C4oq+u
voUJ2VyK4Fc5iVmZQtH4DM/BEuUeKY7ZjB8zwFhTqIhBBV9Pva1DBVY+SW31E9lbQ0EiTL1VlZnk
FU+UP4iaVscB5GztRyJIMkdP5uqsi43ng7NrRbXkY7bZWPdMp9IcoFVnSEQK42LcudicjoF9pv7Q
PX/QGJutOvNZVwBHhh0YcQMEkgpm3sIu1IfpNbwv4419tJZduSurAx6UZC4CTKqO2jFACa43esQ3
fpmcXMbv1ZWI0aAhgO/USHEAuwElRb++P0BSEe3P4u2fruwt6TGbKm8kYpg6HL6bzNxbKGzXMvZ5
T4osZ0Vk2g+SExbjJcmsrjSeU4yxePDnvNYX+bAiAWdR2J+8mcYFVoeOL2z35td/W/pCqN70Xj2O
AexD/lcWa8toQce4vHJFvoXqt2XGI/6zistSKIyusDA94b2yQNl+mrFK9aCgrhry833BP+iQwBPZ
9BtYDQFN8g6UIspuxiBu4a2xcCxK5wPhimGhUbPoQTD4N4X6DBDwWmTzpD5of8l9N4aknMbEbVDT
LlBrANhfpV4NnUxTWPpa+ksBJ1rDAcJrrcdzzEFLG3WaKPlexKbC51xd6uRdyf03LHJdxldoFSTU
wHDe005J+olicVUcxVQp1WnnELXN+9xitNf4rCbh7tVLznjS5W00VPEcSBV5gEVvczWBS/5plwrg
xE/qGpZtx9vIz2j78eucoyDvJaaBBdjhpU4ZoVzoudyZRik3T5mkjrPZrurOFezmhiqF0ArSmK9f
2KWKMQWDkfv6dUAP2UN2eq2TX3jAxLWgRiX2KnGHq8dQKE4NNyE7ce2eGbMk6G+N+MQ4yNO7jiMh
afJ0yWV3qwptpsr0IJia0lpmsOyDVwrbe2XUEOFgFiKF/clvCBOMnoySEL9zzbp25NWUz59IKRZJ
5aU3iAequwtOxtnBYLGOZtAUuh1lEBU8yoZmcliyqqN9aTNUMMLqNROcj62cS+xE4S+jUl3b/lsE
e91Sp3AJLnXezAMEf3dIN4ma8ascxQo4MtoDJGXF/mng/xRXLR1Pck+ycIcGCwTM5sOeWmGugbkx
GTwK3+hWPPbt+DD/ETme9Ey10Kpkvj4GnOjrs5BDszVPsmLbTbMgCxYLLSI2sukzrW9vXVFzkbpS
jeWJgczlyNjZ6CDFu20JZYR/Opjm8QTLs1qDkl/4i/JhvgH3cDOGFhpQYzUeaa8kQgxHgrEKai9U
PMxqSMB4cDSE7ZszboKyJ93HgShdaika0np7ttdQPAPGsrtTRArMsr0gNQfTcHchFgKtH79yYwL/
JGAobW/cc/tmAoYjVbmGdSW4BIHAHb+IQdqDjS/EzDqzFkZiNURcSFrMYd/E1/KWkkk2IIv4W3ij
Uo7kbEQyjrs8uGkFXdlT/I0pShNifyPIrWOW9pC+bbady+md9R+kUZ6cZkKNBjMjvJpY5WUQaZP5
U/wdJqGqKZhIWSeCb/7I7KBchMDm1isIBZphgaMXaOma2AGKfzaIH2IwDMbbbie28TERMHdxXhnc
Hw+9/lk21x+7YrGpn21TqgXzJJdMMquObGfVCGdvj0i2k+GLYgTijLhbQKi/mhCluDK51TcWO+1P
xrC5USaCWJLWvEJqrKvow+O9/vB9RuHLpYUebkt4xU+7PvPJeR2mDL+TJhP6Af6w2pJqopnCGJfQ
qFcHdXlkSAMtor6lRR6X9q1AAG2dvI7/2xgBAe78Lag5SBj8FpdtnvKH4WRPI1QbXpZxlXjBBy3I
aSmq7h2fJBacvLInla6LSEUSd68UYQ+w0ZY7XadmVFqlbYyDTWJR1eFwcvETJgipHs8xwz/id6nV
G2KJigEBJUKLdnoTekb3oFJnMDlrLycqVgdKVNcTttqoOnUM3kJ/UV7pnh7aX7ZTon8SX6vSlxFp
iy4NQMt+U/gY2GUXrP8IArNkGnjrEJfF6LoE1PmgymlF1g55NoxAi2hC92ZXbL3CSYB2NJs6BdmR
nRQhSDSQbRSM4oCY4pWzoRKjC3/K0MNt5iXN5yLwKpF71+G960yfwzLwwXX3PcJryBtIdQURS7Vk
lh6sLH/bwpDCIeg9MozYgRdNwVWDYhkjLMAccG/uWsUqaoKzTcw7WORJ+2zI6yT+iuC+yS7DBjvg
rDgwYNv6xHnfQcK62fIvvYbKO5j2Z/14HVNnX04uXmFVar96zE7ttF8m9U5fwKxQ4CzBv3BZ3Ost
4xezQ2UjVd81nHP15T8j0on8H04RTVhicmAs6O/9riYZOZGna2VNraRQCjCQ3Lj4Jq+aLkk8czDi
1GU/1Jb9uOaKPGaENeceDGIgtLQQz8sy/6Bs2l0YP5h/5PhbNrwQEJnNWbxouH2ij+AoBizvwvdh
Gm+urX7zy5wkOwpJSG86OOo3Na81LuABt+9ZjNpN3UuokS2pJ5rmJjlDwRcYcQ7vVPH+ubUdJ7fT
MomMK7uARzSmU1Lf0gDZ4DFvb+ANm3wxRugOvP/PRwqSEUw71tqaFlDM9zCc90N8L8+F8iVy5Q1/
yqlmHzlyVNHffTR0vVBxlSFYETinepb1rJwNPvzxWMFD8tvvoFwJc/ClRnefy+Kmqn0JhHWBt4Pj
cilOZbtrRu8zVQ99dlR8+4cPRlPAo85EIEXDhMKNOxG20KvZSdoXSASsAoM5ljkQTWxgHLy/6kUc
KE/u6qxlwj5I3oY+tDeqW1kcTTY1DJ9bH8wCoUkpyWOl97qhagSlwkA8MrqH7VkzaLd+G12k91ja
UUojd7ln35A2mGgt3JWzzTgin6hVHGZgwet76e5PQ3SHexXRLktDkfOOY8tJv4NYMbQ6E4rgJC30
l68OC00Xmx95oK9nNKAUDgb1sjotK+xE04V8i8iBYaGQZJ+QTW+VpV9k8qvWMmdu9OiVQOpw5GNx
N9M4dgsDNvId/0YXEjv8xt8iPzHPZ6iM14dGU9AHzqRmRtgvGrOEXgVGPrIainvAChPR5yJJnw1g
2aOTsC0wuee5F9o3vvrc/+X4JmyOz4DdD8ClTqd1E2lrcw0H2YXHtJmgO6OTrYtjFiT4d5P+CXP+
Zm6/6c4WgvApHr2RfveuKpgKE29JoQ6noeDG+rD1s66dH9CDz008X3jN8nxn5jmLEzOLs93aE9ZG
DZhj4nidMAEm0n41bZd5fMNNGyjHeZCER4MKBmeSK8J+uwWt7Cq6N7snLZ/ayf7HfZ3H9EPm6PWq
t68xjGsZ3UmzVNuuvMiMtitUIAlAylRgXei6OC8eZe+xvh7vtS0Qsfhx6zDyxzqChUHulqwsODGH
pzNdnVzGhTXZeEh3Ul8n5Pi00Q3jHdFR5WgbtUG854lCrskS/Cq4Z89DT3ogcrCRjlAsXS7ZzSN8
sEYJ4GECaiJ+2q/jmmD9BlwsZuDLdYwgxYJ2pGcIyiKpotyeJ2Ss8ynqP123M2zkMxd/xKOcrR9k
A9F5MHAmZLj1TTTgXCuKoNoSFPeHOPHSNFFH6KBwzGt4PJRCHdkqnb5t1Dxfcl8GxTCB6UJQgcB0
xb/213ByJemb3JZx6XDHxzKR0VuiRYwcWAMS3FTVStSJtiZ7Haw4QzaCqLnXDbjPDpfDDv2ehUER
gpdeYcLj8/juZUTmx/NsP4bdzJ88b5cXz6qlu0Yp2jCj90mUP7iau1julO2MzshbUGq+WD1eTiQT
Kso9NqDn8YLEklDTScT0yNw0fMbkyeGM+G63Bkg0BQ1AZiqZMfVlbZhxkOQawScQfgVtqksVhoAW
ir7l7Rtl0RM2GlYKxoymwIpi73gqkzJSaBeV0XfNZ9KNQglL0v+dXEeU/TMTRUxfzJ3UD/OjlXLK
qmqQ1sTzffu/9Em2JHelxlfM3CGcBmOp52Fp5mXUZRxfqwYnciSYm505QVapN9cMG/ONhIxfaJUB
xkpvDnR8mQAr2IkZPgE3yj5KrIVu8zggEYnNUqieYR958FJOmOsEb4Oq68Gu4lt1oolySwEZOiEz
93yFCWOD2Wm/vlkc/avqqg9iu2qt/ma+wD1O7nvzQ0uGhnSeTPbrBAVaJad/kIE1y4rC0PnzbM3W
UI13NOXtVPqFLIFzUYQmS9Q8CIe62UdXx+azLC4tMHif9R5dfhPoYTlna6Ca08jfmEdfDuZmRmKl
1NxU6FaGZkawaHqCUU4KkKK4mA18GvSR0MrFOd01TP/yjg7k3TXhrAWCPkT0hwNzXQXLFL2KVw/F
JjDq+Duyqc5xOEuCEDci4FsWw3B1GEgFbhSCMGrfpwl0/+NdX+bW0nE1gYbXqVq84n+dPAQZBFzu
tft7zbBcG9USqBDAOHGGqggG6nUmIrRWXsEQ2FKCz/EfyZQadtQZhQadYfVYAdeGX4Or5pbA3x3W
cNY+SGzU32Xnjba7ojTjVIoKN3J49WZPxYivpXMiljQ+5oQPkLgEZ6kERZGfg9ZIdraq5yOyAOl1
iUz5ST9HqjtdzxlJvminbqWOm16Tgqc/ZlCza+Q4ef8cU44QlTZRwW72k33/nvvj2EJeqDMM/i2o
DgvpPgdnZYVICmL9oig1iJRp97lVyom5baDZkjKPuwt5Lgv7Ttxgl99Wiw/d66eeQ23m2e8KDo9f
aOvCL6oOVKlgrTIgyt/zU7QkNVkOZcbvYfhLQjHDuzQ5vZ5SB4WJ/qhi97uhKjh8mQWzlC35FuSq
sbqAqXfI7wBjC5m7MNVj6oIJc9/Qi/UIlLGICcjBpwKQJFFthC+t8aNTjc8KCFjnPzAtNx7iOLmm
Jvfg3xRzMyxeQazlDAKOFY7Xznd/R8Yz507tmF8Hoi1Hskt10+e1ZOtRZUGMJkyXvEspHF7RyTXE
YsZB6Y33rXMxCkNaSYFoLbLQ5rdRchbACV/rm7kyJ7ndFBrmuBXtf3NUzkSy9/K1m702/GG/sxdd
CqFVjDbQ/ONPUS8h4iQb7r3iYsWZjgeAQeG+U1QI8eoXfBmtBoonDtDp3XWB9jdDijD2sd95wQ0h
KrdV1+dCzmA5MXMbGnCaBAomasw5LBqQ/UBwN2JST5Xt1IXLR9h0K6k/vkOpoXKvJwm06ClgFv5n
GcsyYNwrw7G5PtWsdA756Vioa5xjQJS4WJ2sNqndgvF4g0QCgJWn0XaVIhlFskKYW45bOc5saoVg
wSxsuZk6d1BDxfJkT04ApU47Y06C2M/W2hy+YQJl5+SXlm5luG9V5xCelFfO0jMMACGoj+1ZCFGr
chv0uuUrDaHlEZmGcNF2WRbcjXhR7ianBRXBuIQ8mPlPLbdCDNwV8cE2lNgXfiUqBfnWxQeRlxwC
JKv+k0tqSv/IhV5zL7kNu1dLGKx6ObaVtU0LaMWlBi3LtpZl+4/bfNl/hDhEPAcZE1u9CJno8T+1
R9u2FeJTlW+nhHhpZB//yXpX+wt3c+UL+pA4Uc/KTtbl4CP1jsZanrQ8gmhf7G3KALVhSpjuernF
IMgsz+jt5M6aUIMyWSJ/Tx+HBm4lq2qhvq3MWw7qp6VtUDSMn3gfGNF94LRrDQ0BvwuNvqCQ8LAh
oydenvJ5OdL6iUGdntnSjBiGFltLSCwqy7SmeDrgFRKi7mQyXkgkkvj08gpP3bi9dqyDVxhC2aPs
QrKho35gBtpJn0RzZ0HJRcgbqmEt6xj0h/4NstcP7JR0WyRHupbg62qUy0dMImoEsZmBHpxRUpQ2
dvLbg2qKbGNVlwtDr6kdAeNkZAKrw9lIbCzyGfQO0Ih4PPVQFxN8nI8laJTvF9Yw4DBBt3U1HLHM
Gldwrt2TTt2ojK594nqoHANaU+CmpVlSTXmSvVvCgitM57Ag0C9UioFeQT8EPs3XlA90nAmtIe/K
ytR44hJl6hUMGN4iumbkWnC+lvggDzDFjWdFHRJ4aFJrYP21RLBpylMexDe2Z3JAk7t4F7jW7Gix
ZUTQqVql+zR9XvmFoHxT9Ye+1ZUKQhxOqADX97BKrXf8zydG7L1phz1q/UjJJxnXiPXpi75MzZ31
kXAuag2WonSZpIyoXAMn70m1WhJeSjWzYWxLpWfbwt7bow43VH0bXudUDJTVT6W19ExNjyywITic
BFeWeKL+Q/xWE6rmxHBk46ImOfeddpvXwr4vO4xWBihfmw4RIKT8fqvK3vuAy9XRDp/JSUyR8I+F
WsRwtVVXz40uqZfUvgRlr0P4WK9UBVzn2UmG3tlG+JTgIfPxcqsFjq8NlqG67y6s47jTDGdk7T6Y
YiHQlLPyYxMNjhqc1yqiTt5XPtIpdOmCPuq0+8RpvkR9CwVvoo2cKZDNMm8XgeA6a/LZdNgNm++o
srG+GhlgrCxaj3d4afqkHKZeTqd28uzIskjFy6F8TGVwYqfoBiFYvLYcpnbTNsAzXFEyDn6nH415
6QtQJrrR6hy8tfF4gD25BUQrVNtH8MoqY/BBHIrsW7taZ/XVMuF0ckOb6nwIRA2daU3LisnlcBuC
Ns6GTXC1DubaXw8L9+uEMtsPCbZVbJTyscRnglRpZMz0ZqK+FL+mZDCdUR50hP+y0mAwh6AUunRD
MSwLBVP0VG2nEgNDwhsE/FvFoDUwm0o/M8QR3uUVsrde9iMG0FnQAnUYW3qu29fkKCS976jvYxOl
bXNWQU00mny6CZe+MKDVUJGTMOW+Nv+v8LoPfROua3sejiGUvZO7zSK3t61EYhdqynJEkMBOmOZW
5nR2yJfdUPhbZKge/tQa6HoAdB4VCOe2VgriZMLyqdJ5wTqUs7Rp3PQD7wqz02V0tAOoQgrUuvHT
GdnZYHOeJuVeDWdi0gLYJ1lQ44ysvCF1NBYCW4nzrm6dFAqCdOsCO7pVSIBcTHmik9VLwvVz4NSU
pUsMR8yHXIqWyJnObki8gdb0XNJ62zlyl71nycR23d5m/hOjwYjItyYV8Y5b6yMsXnJgRwCLXLia
tUqj2z4vHUDgIAwLaJNfu2OyV4tFhJaXpQKI8uLA3vfqiqk/bWwRrZhhyMcXP4La9zO0FB9WMdiF
gXGWIqGwLfavRVRns7WwYIIAV4+PNNsN7fsjs16l5kEu0GXJMcRjZVxrpIhACcby6IRGlWgLyybt
KTvIYGkf9R8PNLea1mxMzjrDQxhkdhkeg+EKY+84Z9ikpugn/X8d2QlIseRWu1sdgBj5yStVMvbl
533OG/4+kVak06K1CcIlsV2VwOTtnK5znXxwSiVspeyR/ETmx616drx9CcycHqCazTTjbmZVhicA
upSeRNZ07xr1QDBrJPBYf5KRLYlupcgYI7+B5p6j3r/bMgbzCSleoIj2ifcQHPIa2IepZfxx/5S+
5rVRXFj1Nk1v+a4z2rhk6D/Iq3Lh7NJRrkGpJi3ILM08kOwFnUJ5Q/GhMUuoMbqqcjPG7gGHOzPH
oZuWDQnx5L7bikvYIudaCmS1g2pAQw2yiLceUOt/GuRFvosrccn/c5bPD0Omr+2BH2TzXAyiWqZM
26dd2vKfcJF6ZB3aKW+1l6qffoGf6vtxgQum3e3HR+66NpTRio5b1CnFiyYmKZjXCPQkWA7PRjEY
fr1UMnYPbV4z7+Mv1sqRqI9FiPAvkZsb7gzZT8aYuO7iUQ5qshTHMkOd+xDWjNK08WgmcXZAyy24
vA9vo4QbdKnfShES5vyacJKIe7UJlyoJvdFU1Z3Rj0x4H5pTyvJ0JbcP9n5Xv3QLsEsrcbuJt2ZW
DFpi6+RROvygLDT1JjLeYKzDN/nNAozDAamUxR7LdPu2lbU2+Su/P8ZlRORCHWh8mYjKsO9s3amj
3W2kgnyHdxbrfCtl2MQrSFJf4WBMeDF0LDJ97YclwmLDdBf5P6jZzwhTEHNbPwdDBIDAP5ii21Fp
EA0/D7qObryauJRsck9WWnrEOmGvjUHxhkB3letftfqn3mfkuj0e16IGPq9lSS772X93VrJysss6
mGcrJ9V7dGrzboQt+4+0n2Gf/sMdw80dRzTrCrBPI7BO8LG03cGNL8GyguitoXmWUFpjlp9QUo7L
pTKOcs0YCtkzIe5sxrry14+Zvzah8AN+luftAG9SBkzg3QkxOU9KbHyBI8hPjGPkAZ4pilKnTNSr
kHhpkU0UyBVyBq0WRPe/s76qCViv+dcno8Zo8WQUOuQobPaJw9wZ37pmUU0H7bdb+EnqnByAJKaK
YTfbx1ZGmqV2Xghk4TnIe1fWzwIhVDAy7E6Y7uad2hOIn4nf83tOucKd1CYVU9trdLk7giPl2r0V
9vpw0Ve/xMg70+1p+8GhaR0sFHDa8+AtlS4r/nkK0LHzExC6j0+CHZRETb7iIuhvkxSlYSxPEjFh
osqouzvMnsxRIi2jUzXxk1d8iLzQXhANsxmkJvyINfoCRpuvEcmvvQPsdutRM53nf83f+u6L7Kpu
L8jGuAFq+YtI7YVYVHNuibXIcJbPIgISj3mHLPOCakXs+V8es+vRVZIm5BskQFXvyBqIGYxH9CLa
sz3VlHNQ9tYnJDVTbeu/UynSrhmtYG9o4++vFQWQYC595AKu+CgFZmjp+MWI2V55XqbcQm+o07XN
UJ8Jot83ZKbY154VI9drvfGNm/jlliTTqOHSzQYbZC2Zf+g1okXs3XHnnbaIN/7lkvoBv/CAGuBi
zvqoPq5LZqf+BYWJxJmwbhw725lHw9qezL9GpiHAJdzUVn0BCBkD1XOIYRg1R++h1K4NwhcdH6Kv
aDWtM9wjWHGuZ04k/S216Ae+xt0tIWI3uFbI1X9U+l5KWUIUvuAxBJxo0RNoU+JLKLLC6n4fs62a
hj38ZrneVku79lW9Ggt11JqnJbsHr+v8ittEPeTbVuGrMT7jt0vX//Jp91EkSvAaaQ0Ucp7HLx66
u7p+cwVv0SMP8zQC7L5uWSZbK13LKPdK5w9ACraukJxiIWfH3WU0L0/VClPY/VoAPHazqbv0MBn3
gFPwot3aJ/klm1PBUYfYW1H0KSDb+kkIdZFLbPJp/11F0AH9iA0ecJRsoaqyxfdxp8HgI80+EjAQ
Tk2lEKe1dT676xtZ3BwJgkyzbdpmNfEvbyM1C/ttAgQvBr+cIHzX0krQ0jlaGKOjV5sZonRcuPJc
LYO3G8VqQpm+wIC93BbBgD/jnUYOdtO7rJXVao8NnQ8GINp36SsUhXQ17r6jutAGKFd1EVsmHrXm
c/KujsxuKX8kfnN7LQrdqhElNFdXEd+7C7gWbMVpisTa6MVoVzHb4RS6+aVr2xywM3iAHvaErVIK
gMw8Um9txUYAb2l6Z0+PbRk3+WSp2zXfnb64cQI1hKtVDEnEoFBmmdKWyzj85WfTwIW4FpyA/AIm
Vkxl/e9jY0Hop7tDgBBz75MeGS+Ds/snsasSZzucqgauJ3UVj2x2l47U+FB0pwyOXEZeWsO23OwV
sQlV+4e9nvLJxqLUE1OZjLb3A7dca4Lq45c8z15HbrlDmMYG1cWTtrw8vnpdlpHYCjEg8Ta2XuBN
C+kSpMVY0+Y1L9zES/M8Dl5QEWgl/CN7+kBEA/AgMjgkRoPE8nTCdqCAAVXlClzVj+wl+8BybNDL
TF+DzbcGLCzviDabwMru+8N3TgPPsAHSNt3QrW5dyjpelbXoambNfLa+gnmwtcnBwEJeqB9U3Sw9
YTLTjIXpeJTgx8oVtijxwZ1n+wQGEVpLNMZUGn2Hf851OSJHw4BYZ/5XcZULDB4lmS4FOTkhdxD7
SGWILLd9wbDiD5rNeV/nIYM/cJWOxzKacClzGds9Ko1xzBr32Wijx1lak+WNS1VM3VXE96EGsxJe
9OHGyGnfDUw9UoJ1dtJ3Ki3F1qh1ZwJDfVdq0nD2KH2sXvS84O2zBD0Qz14ei4nwXVvO+4pwb0Zv
P1iTMbmMA5+DDVE9ZGIkBcjmiVH7TCoCpX6TktizcTS1xOTCNTtp3nBMDliL5/NxGIyOCTV9HJkN
A19hZ4OrJ4wBKJGqqxWAwkm+GfGkgmmATd6itvw6q+Cpf+mFLeoKEDpRC7PsGPDigfog/IystXuL
Li3TtOoz8c5zxVdJERW/K6DKwZNxXozSk3MieLUC27k9QI07iN/miOwxw290Y4tAwbL43VDVbfH4
LwjAqvacJalm5Gr8yZ/ZnpWupY746Vj5G3kdi4Hbsc64MPbabsSztMNPMTG4a/YUYiSAeLIkSaFk
8x//PIaPYqYlI2AtE2MoFDuLvx7yLh5K0lu8TC6ZSG31VO8XRXDbDZepZcMKdeXKwRupALyKKIm0
rpc1X9/W2mYdTeeRyiifCCJmgxIaRrN3U52m9FbqXL+GCrHM+T6a/C708SpuHWmUpPVQMuRI1d6/
7tnFpp7FRqB6th6UzFDf4sElYRMpaJv2LWccGodr/Il69MHvmZYsRL1pMqsyu++2WEkEtxplOtd0
k8xn+h08OoBAoDleSnqjmjn7wqaavSubTW6Hre1TP784IBuPRsKpcJRjZHN2pIPmy0zBmhooLGgq
s50dqk2QbgdnJWoAatQ6qBs0yuoQQB0bvuYLbt9anc9LCFzap4LYwW8SSv5t+tZDTGe+PZB4X84o
P8nSPuFlPy0CYg1DM3vEEZ35tg0eTUycZW7h9Lr2zYldmB/8C6lEOe2TW22sKJiPj/qaUPIwwxte
ZzTodbTn4RUXJ1GXImwhjiSEsgsP9UsqN/0e1JdeL5GI3ydEhkkh53tSIAM8M6JoDUxz0cdnvqfH
zY1A/j18XOkVGtK9R/VZAR7/6RFyEyL09+9+zm2HNsKwLsU2QP6DRGc52yni4Z7D7BmF9mzqQIRZ
IS1IMW6YXr8oQzOJsSPRYnlPP2OWWiStvBzwrColpfp7aLmQyuXPWBVrDKHmcrEgYBUZVth0WVuS
FO+zLfxzEYEKHTveWYas6O/QHQrrQZ+tr5KoAH6NXnt3yIbIS504TYxSVNRdRJZP3bEZdll0abxd
swI5P3l1wMlHVjL3nif1rfLu353I13pzGs8uwJx4K48/sHTXSt1oGKkCZr1D6fdNDwYeY8fTE5+s
PJFhV2a6PqaF5RFiH1QioKjfnvg1eUEAf9FgGu/3vj9PYh2RYCjWbpncgwy4Cg1nudXIuAmrRWFx
0JqOo1U7KFvjBzwm4t7IK/22D1VIhMwBcjM4N2X44I1aMiXc1EqMUF1ov9H+H5oy5Q9uFp72w1/Q
IB1Y5MJsaO4alWE/uzT8Kj1LIwua5cbzbvt2NakD3r92FPLY6Ue+bPBxwDmmhjlDZTcnHBJRe6x8
Iqe4QTduQLlqU5mIkvzhe+6rvUdHhWEw1ONvhUWinqg4m754TzxACGwKyf+krROLqd2q+bJYUGYC
FUOs4NoRzLaklal0A8Zt/kYp2SeLmh9kw5jc3HJ5R9soCEPMkdST/+dIj8IFK+V2LMBmYfgWdJ48
kJMKbczLsBeV+KiEb4oYoqtaOZqDVP5eB4EH21rsdPMuYLLe21WPmu6gv1iVKl5X0wFmutVDL8i2
uWEZajAvuPFvZ+E9n44QYNI4NzfKw2s8qeNgnlzy8ik/bgVIbq1UAEqlpZhsAMNybL22r3krMG9c
eZImfyrgdvWfQcp4emy4JkQHajtguQJt1TXu3oLAkes1QFR9t8xxVDj+5Y2xNMmZ4HMSPY+p9by7
IRPXCYiKdKZRzIhMXrid4TfUdlaYni6NoNoMdoQMtcJaf6aenUSdusxHfd2L5y99frB5Pp1FptBi
QDjnnlWhR1q30bhMWmRZrSDXbwZoGM4igWyoPkIZF2VV986UyYxS+9l/0g+6cw0N/fxuQLZlX0/e
3hyQeB0K/Qk3HSttbYAYx7D7HzYWcgqMmSgnxUZBxFqfVEQvmqrIBWMYAsUUySePXHu/aX8YXwI+
Hf51wKTqV3N7FxZW/huJg6wstUYG1OtmDIyU+uroUagZHwyrZ8cnq5SbEpo0TEOTbNY8VwpEil2p
ZTxNG8KwEvU2VkS4Ku0rM6E2mq7uNC6JBzdrcTnxGTmIvuGjlgSJFTNQ4MdE7+yNbXHvTC3KZGPq
RwsNyZQseglDmFFfqMtBwyISXXIlm4TR1oINxfeTngcBcJwvo5gWrvINvXdD7WQpDC2j/DRXGB7t
L6jILTz2agFdOdYAfUSM2ZvoG98pO7U9cAOa63eQrAjx7XjzhIuDc71uho4AioD4MOxkVeEgCNqS
Q2EQfH4ChZU5UrI3s50Jx1bULwl004jjpGt1JrxlIJEphUD24CdXQ8nxTbwpqPZwwuVLv0rZbjg4
HFc3rEkld/auqZNM9Y47id5IFWonknRZhWuDhmw10AT0wQpwQCEnVOnUtO+BXjuqoY8I7UOdehRC
pWCigbEzs5dwkUz2OoI58rW7oMWFSyQUus0iHAFbCuRh8L5QcHow0cgZEIExlu1qx6W2tTHc3PPR
qjeOPQof6M6D4YZF0BYp2TsE6ImVNbRffR+AUF7brNeTrgWcfNtPoj/+On8LHFs6Ac4EC0t3EGtS
5weSK9CeGseIbcuzoQ9JeKBBYJmI1W8Co4AbmCvxHGk2xUZaK6f/4Pmz7Dz4wOMpB9S+QJ1lioRD
0A+uyoOUaU91AjzKPI8Evvy0LZOHsAfOyTUYSft7xwJy+DtGvmfKbZy5J8uPBfJx6oDyBFAm9mrF
0q3C+gnuB1unI5+gxDJlLn1+z+nw9sNEZWb9BQGYeQ3fuUcJ1G+iyG4o1rQpTbXfioeZfizeUDHq
Yy1L9FmTjaV/83SB7XxGUfqxHDmy8AU1FaLBE1BUhiBJ5L21+o4UHlz4H5HF1ijY/+czOsvBzlcc
peC1W+2RuHsZvd5A9cb9vvyzWujnr/7s13JL9mEX4iKsQ0y6wZxhZXhxB1LkNO8eXoGfKfQMwU4h
S3Y1HsiaefbLnH6yM2UoBs26qIRQOIEQJQQQRopyHfQaxhLGavwuczJ0HZr47OaaNIpB4iHebPyH
c9hN0RymLcSVgSvYt/kEALwvIiPSEozMtYv8KJ7cDMmXyIrtHByKtACFKlr/eGCsWK+x12JvuOMt
dNzzWlcut4SJiftejpG+TyrzThgp9CnuSXTw2bMKDiwwd9cq8zgi8DzdWXzNN6oXcugXqdpjvvNf
LkHBZA306gNbzbiRzitPZ0G/MG/YSktPWsVxVnH9pQnuR88VptYP+YJVAPhmTm6b1B4UrjH1oTNB
2cLT1GP50CqyN6pBsGDGX2sryZPahPnvYt7K6DHTZgM5air+OkXF4Z4hzXgGrkEbA0QGttpFcb2r
OI8buhLlUUmImTvwY1hZIlHo6ezq5/rrZ8ionzlIMZYoWbkuSHZQpOFTWlZVUbzkIxfkK0pOD8ia
eLMj5kUVSX/Qu05TB+hAVynhFUcN1xjWJduXplzNovP95tnId6mwY/cjOZcpMvV5FK4C6MlILORd
N4CbAeaOAjl2zvKVVo5RgLf+Hff0goWt1NXvR2xYFG/KuMkiz9MLiQK5NR009+YwqPlvnlwmuEhP
sfqnUK+5T6Xubu3difEtfmxJFtPhLAF+WEMK1R8wg7XrMpZ7bjFQcxh8UQMhPJwb1gJlCj85EyhG
Y97NbwmQfB5ABDPVCmV14Fbg6Fsj94i03E5o3091tuH6/sITb7uHd7Y2sPesn03u/E7cesHX8bJk
23jPdUR9T9HI824sozFS39hzc+rG7KT6uEgBeYbMEo8vQklRoNA81K4A7hLyCjtLZt+dEeli1F6E
SNMUzhZb179FUHpYGPr0ELp27CErR03y/uld/Dqepx8oBz0nLdGyWhm0zdeGhxGx61B+/3PjdKls
RA7fJF6h9NwKqEzWeGlkH+Yc5TlWRxj0+UaQr5TGfSqZjuRup0vwaPW+9wQikr8Lyg3gAqlJ8r3K
H8Ze5o6WtBvPzVuJV4LTLw7Stbdgn52yPmn3MZ44ZBXPWMQalCnJW9BeHWbrOG/qBHZydVT6Y7zS
6TfOmW0vsVcr+krX8Tvod+pQNvu3nhh5O8YtNZCuAtT1e54Ns7+g7rzqZvsJaIZxLc5geWB+xp5s
JYjpQnb7C+E1tcxScBW4B0MwxMPuVC5KuBjbcN9jHC7Uv30rz85ji47+tTdoCfd784hSuxTZngjZ
asgmHsDW+m6Sv8e41ay1/6HSyStkewwnbDeBDGt3SVH3s5WDR33Tfondx8EK1WGHp8TDHqH6iNkf
wNDAbYzC7TxxD4v5zUZZm/HBGaLyIFl3LsfP+S+MwTDbkrl0YsGeAHrqXRVMudZH+AkkyGVSLy6e
OLWowDsL1xTqbjM3EUuamBKzvm/pRqHIdjffNPLbpjzzZcEKqUrf/VFPKSIF1y3Uj1b0RF98NDQF
04xLwdLNSVEAt8xUE2UuV4z2n+S5OwE2JXOjlwlOE431BZn1u8Vz0754xH2TZbppshKs3uA/xyOy
JNzYzHzH6WbP6ObcYjt3eUBl14rKcLGF2/7zhPzC8nOzP+SuN6NTVtotc1dIYcfpdilN2QsH7FaM
+aA+jdchw93fgmHd+IWokuuiCxXpqj5ShIi2/yKIahcGdPUcIp7rgbPfZq3iYViliTMhG5fwJeGV
q6RXZMtHvx5D3cAC5RgJHPgkz5egOmFiRRMO6MqAG8jdnpGTfAO/fS8sj3ioSKkd7PU5pn4bzKQg
dEjCsPLjYCNJsz7n5XxqqieE38q5rcwPxgf7wrUDgBWv0amoSX9jnipHYNhfR0JHWE1CaTJGlX9j
WjN/HwKCiMoYGob5czLt8vXfpzlXWwNj9orO+6cVHMkjjQZdQWyQY5q6MZEW5eLyCoN0A1gPWDrR
h4gkGnhnDr/e23EcSoXHFI7WbWVz+8qec2vcaZSsqiwSlMlEChNMMGtWKWpbRfiJzQTLSw0YNQQx
2/gn8HRnZKCRq3/IMy4jKqPSKJy2VnRpBpEP1PcVBhLheFyJ9IJbzMKJ/wjNzoPsMk1g0M1zdNu1
8qwmAJ1yJm4LpQ6T+KQt8wYxpIhQe2GF0coCQfk6qAKV0B2iVBwB75/KBPYo6yDocpUyfEK94Kav
NwhPdP+AwdyZiFgNHberUlCvgGGfemRdDd/h0gD0HEQ0sB5YmXvYX7x/zuYW4mIMEEi2LQc7VMFX
Ap5JgndGeChAmB4Y1rFeGqFZZg70VG9XPenUidMnW2uc0bx/DCBy5axMgT5CrJplewFhkRk05EGw
JBt0crZrEa6aB8HJDBcHuYeSPMAJWAZ+iCzCX4pqkpA2CdoRsz/GiAFAgNzEKl7A6VJAxXN4/dRp
NXwbUQNg4v2A7V+DVl4NGpc+Z1XapZAXQFpgUuv3eSkx2kk09Qvp3WSegzC/f1/qa8QxpSEpY4ph
Va0LWexunqVvZNL3r3lcfb9K5ku4esHSFnfodJpsxUpuHCYbOz/8TtQgVawnCviQ9ioEKRSAzwNt
bPcSut8TghwaYqhoO5lAKiZwJ2xzy3G34QsX/aEQAlizHyAg/sLWqFy8FrRIquk/qzJJLSO75Php
2RuwlSr7kYEdGnsGyNffrO+MeI16WYeHRp18sO9mNWSDuDCvH2r1+/xlWIPaGDbyFNhyxO8yWxRx
z6HLtOj1MKp1CI1lRqMWNmdkCcvnEgdGM7CkDLy5nwv8Shbb119WDWww87lSRL1EUkSJ4BSwWpv+
Rj3mOXtsxr4KPsPR8iK5w0r1SFgH1/wA/y0GI3pEhJFq7NXLifA1dNf3PkqmL1p1jmqgoiHFf7BH
SlH1bH5U6p4nE1W1IlRiwbJ0LowlLiEe66vdFwVbXgxycDG+6Fu2b9hSxVWHZw/4a9ml3AuVEbN1
o3T5lnKKqRhobkc70jMDdqMc+9STm3NnJorsfZLNHvM8XAFJkTnrsvsB8Yqi/mEFhyiyZ/3fC2Be
FB2rZz7N0wgwHG/u9WcFC6j+jJoVjqfinCqBc19JHv+7/1aoyCO08HwrGajp9VSU/qXfKz29yDs7
L+sIgCxqin2PelQy6kMGKFlAFWQWQK8XjkBIKK733C6iBHgK0fq+sh0wMHl6x07biqXPyXqsxlcE
zbUrH+lrUn188QcIqU0unzqvVX3UCVUPoQIiwH2NWuVjJm0iRcDXtKt29GTqQOEIBbYmXmMpxXpR
hezbUR9mYiHj2Ri/0e1eiX17gNC/UAMGjcmiqMy5NwxT9Q2/d7iZHsEyV69yzRXHSL8gmHdFUWV0
VkoWw5/f6evpzjKVWuP9LWp+XtseYfArTcLrlG/0m30F642nBO0AFvDianhBkWm9SgtZhjzWf4E1
EtnJXrpSxc17EdtBt7DUoQ/dYCIlyhwKsmxsVWWObx9gghkoHTe6rAkNTTWwMvp2SCvHhkRDXB0w
qohZfCoWF4+Oqc5HSrVvTOHdbf6A0ofDXm4BjHZ7ikFut/AV4THC1Y6AgfKfnlt9I0byJiyW1tb+
wrvwqBgEWj7d+jNXaVwZj1eZZSD4S0cCe7dPEWohInaCL/umnY9EQN9Lqi6kSi59qbBUAuqNKT9O
UcXXs/O6xBrqOIXnSq5OS4AStvoagylY5ipGTa/tZ6ONSVt+OM2tsddjpWwjwWLg8LutMD/JIenS
TOLwhemkGBT88MJ7lPs3K4zrO+ztN+dhL/eacsY34TTlvAx2lrQk00wbUWtwGXC45ncYJV44vzxz
NGdhuzqL9LEmsWDOYRCMKHz2LcDPhgncqEPT5x1h6H0y9PnzY4AQh/9tiLzF32f0jMvDUTpwpXTf
ghiRdwctIHbQGR8L7Puiury1yYUCFpmOmyl1fmsCeir3dMDo8z480LV4Tdoe+Zw6puQq0NV+ICz6
3ChtnOZjWDmBlLlLN9f6nG6+YC1GYrMyNuGTLZsSWxu1W4vS1hkCR+wehM4avCDkNLhOlWTS95fa
5xh4yLtuK9CTlscr34VxdWKY8K98tqWRyBn4/PwBYh7xyoYokcJ8OzJLZzaDSKfnWL0TCI0zQ2MP
pQBIUWwm2/MK5avsIjAOeRwvWyA2bYQA658mHasHsn+XBooASW3QiSpjDwF0+/DLP6Yz5VVLmUh+
YvEznS1LeNEIr5jF9RCdT9+FZz05dqt+JY+/w6mlN51Wo9+aiQ+c6q1Y3O+rXUgxJ26oxEdArC37
LUgW4PX1NUWtR0IogUm3WrrQEwbGSW46LMcLj8E53dMlxB1xmceo5ce2mmZI6xZC92q6GWo51Mfo
IUj+xKFvRU3uBbB4z48g+YLbclJOy7jSWWNWOLyjttJ83B/eF+YdzdMTvQWl3i+vTIsAAcGOZkjz
UXTtSQzbkuDC4GYHLkBxddPjaQYMYLAqEsbezY7mv1QIObmLOfp5Fy7LqT2MSHabeLMtkd6+gV/O
dKtNy2P66QBKowpbM2B+Q95VjlnZgyEeP6rwxEgLOCT0PviYqH3Jn4DH8NPSvEW/ZEqYfdt5JPX9
urnhX2QduWTCsj0z6FynLepGQdqEvZZVU2v1avLO9ZP5qe3JbzwcIzKSHS1Tdl9Flx3nMPYYyZSM
VOYhqxdD8wJz4vv6/ibljd2/R86DNjrf5I4Bq4UdEvdAGsW6s8BjjFUyKKG9HfrPZlEPXCqf4+V3
YPwjxbniMbTEHThD97CrO3NOCChJ1BWY4Bp0jxffhwNwKNKOklonpWY1yPhC7Eqmh69MIFHfL7MO
//pkBwkNJmkCsO9Y6el/bjBnm5JTmahZx8MuedXAqVyJ10zsCtRhpiTwsy78lxE10JZG/MApguYF
W76bh4HF6c9GvyZsQWlb20Qo7i61j+/BF7rz1CHzR5l9l8kajnjRfAlpjj29G3EHrIEwij8UWzYK
m+N2pYIIGm201iFf22z8WPYtGpKyQNk/tz+VjSSR7/lAe5xeM8OWj/QnwzgKm1PpPNZnUZZtlY9P
sfWGtSiqhTz3SzYgUAE3B0hzSkwqRglCd+yFKx9iN2dG93COXzKJ4ycbe9G2NHZ9gSlHecj0uHFg
k+GBVW3rj58kAVkFxdFGPpUDtMphVE+bkiwcBbDkpLYaUcnjVLQYkVQRzrBAla7rsXELA8/tJa2u
ezExrCMp4oC3FXioyzvaD+Fs4sgcehEgmHeNhU8nZec3uTlpJ+9+k0nTXYr37ibess9MnGWsRnOi
saDdd7BMIWaS3+wdaYF9KmQ4748Or9dn2qk934rxfhy0oL+O5U42M5nMtNj9l/haTODyeiU5o1tb
W9TGR1sXrMPO25gQj09u7lGiZzRyVQghGx7czCCTDLpvt0ZacFc5KF4STDwi7TCrRXAmRE+/hNvA
xM4IrxDbQYvsi/Rsu+ZuVq6qnNnfDzOjNlRnP0WVvdAfF+oeInvbN0ScRmIrXYytp++bRPst+F+x
DzaxHdYYZO1UEy9cisoyiNxk1u0bxUebznJbS6PFPYKBFwLV0u0EF5oKmU6Iwnv6ihdH/HsItK63
SkACTYzW1fKhD3CgALYabGP2qykKp5XCdOg5d3dHtIjMCSZg5CxFifsjCNiTBfHwNvWxlZifoajh
RmlSiqAo7U7xdZPfeFvvWCkBUVFAwM4jrX561C+cP9+naHdWCcJV7dqRw9v1axIzNXuOpKrnsyQN
dgFTynMp/1kEXCBgp9HjiwH1qMBJDPkhnL6RtgpH8eM3k1XbtLLN/eCA/sfDEdr/qoRCcwEetP4E
K+5cqwLACzYmUFIs3Ida9+lTcjzPp5SP2dtc/Dh8+x7+p+PG0VfAF9VJ6n+WF7rpis2jf8TgbKAU
XKjzmcwDfjyOhqEBydWwMXHgm1j+5oQn6Z2Int2CmmYFEzaPKqKQL1X0xl4HsHcqfGUSGNy4sHwD
ZxI/fzsE0m71OZuMzQkRcrDsCQpSUJW64RR3GtaSWHJzvniwBdNhfDMrE1lcexrQcNEF6/iYEaSA
RZXCIdbDWwcONqVgmw2AS5yrn2WZ+33gHj53s1G1+358ko4sY+3APwgvpFMGVEizAxLG3cVKFJIS
vR/NjCEbglz5IRRBWhjJmBZskyCgs/ChnMLTEiNxRVZfd2CfMMpm+Bk4yhRFYh8boO49plEYIiCM
hZ6FMd0YSjUl/0t+RX69AxZy5sOPqWL2VwzsLxBILAMg3yCncSMvIkkg9zwUqcDX00AEdeXOwIQq
M4BlRu7CgKpEkV0T4SGRvArw4q2xUOIlYiJPQUh41Tlb0Z646FAlQMxTwTk2zjbT4s5N6aMT2+Dc
XRxEkcbUqlihWsWVS76kxFfYsEM3C2e8UOxGDtBEC8XF3POY8etq8PYtBDXdFP8CaSnyMKX1j1ri
clFmCkpB+Pgwn8gqTflU8+vmGoLl7mwVZ6L0rTy1LbcD5bi1du8y21mSFtePDMH4Ih2fV8tC1/bt
qa6gxxk3XndQsU6YC3XyL5wzFqYzqBLbbO5VzwvUScFGMx1cGEJhQZ/r3gEaP1Bh3RgqKcWdtu6m
2nTIEMr5IZiS+V0VyUqMU/GYDMg8iMhnaNKowVyossF+E4TVBlNzDWz+khSDr3DVUAm3eSk4fQ+m
jbsT5+O/+jo42VjvYxIIoiA1VYCWsnMoBfMUruNswcLOK73mNQuRe4PfW1G3B//wkWbEp1nwobG9
nd2DjTfMjWgsJa613tb3AkeFuWCF9FVu4XjxDwADnWIzMjR/X8UiLOBG3x79gwmwfbUYKxZbzW8g
nZhZWqAT2ljTZ5Ti0pNYzW36csgHXCQaVY57jjT9SAQc1z0nJ/bZZLxJZXHt+0C86NAD0zVsp4LK
TxktrCwzimPQsFetXDcp+zX7Rkb2BRJ7EDctge1OPJZFuhJwAf1+FUF/nwS0H4IL3a5U77Osr7tU
t2LL9h9G+k+TzOFObB7FHLPmI5IL+1+8q199W0UgNovV6xlBmoVWSLVveGwZjN2GZz4XNLtlakO5
B/ZxRthR2CYWZngsUXmWWGhUEZxrnTmhBjDFgoBaYJtBT9zzWDU95AZhv3V9XYOLiErDbiNcJSci
u4pc01IBef7TI/VrWK8qtgB4TCOe9D9VZVwTfI7TsouODW9fMI6gS03v72bhT+/AaQeG0/qbabbx
GVvO01xsYfw5xkhmjImInjmtmyAc6d/YcWQoP/fOeQRguocrTDc5mLJClfMhaO4sI/KDdPfXyNPV
Ib09AjTA0ab4pof7IaNirL5JZgo/7i7h/mN7Mwr2WKQ7ttHhtwoXCbr+cSMRVKVRnXczDEkFIFGF
4mARRmTqgkwQA7oRHXnRAx5ylseU1phqKGAxbnpSnLR8BZ2+ICXfM9zMkeE00BksQlmGV7AYE+9l
IinzsLH0PFjOD00rz24G7e0h6wGyqtBbazti7hcA5Z6I1KgYkxPnaEGx41gBHDeCPZd/4lzDmlm7
7EdMZgdEbPAMAoUZMwYzqhU5mZBCycXmXAOiRHzoWYAPANznwCntfjlchGDSPefB7IHINSFMaLkD
2YnkRZQLWXsscATGZyVz0NoJRnpz2hSCi0Z1L+LRQXCw+gv+776XrCp+Ql1IGAnOnewiwKxMyWuD
SVfKseuNu13n5zdJiooB+LrWUWiSWPudKJSGkdqn03eNcW7jM8iDbM1KGSiWrb3yUmchZRTPH9Q2
D2UH86QnzlmPUFflNFuk/PM3cfjdKqD9L4aS59uEVTmBWoIoUv2qeTJoQ0ZJYE8trlafkGXZYd3D
zryeAuO0hYoPsU8Jemoc/+2Uj5x5cNGJLXShlgcqvOI9vpfq6tuLhC+AoNU14PHqdHCJuA7dMp0P
UsF2d+mEGzGN1Z3jSlPvInOoxc8c9gFG+5pnkP6Om8NTQ7+oLtmaFG63YSebxNv+xjLr4uE4IJLw
xV+kMwGDPKaEfS4/j41BxqKe+22NIaDq8QsyBthkHmHlRWQhqxWiY8KRxrBtir2A5Lf8a0BgxEdD
s07XH4b/XS3ZhoEcq5TKS7Hl90P18h8C1XGxxMVN51GA3CpIv/T7trqpk0fPQNl2/4nlvd4o9QLG
dgY9k5Ji2ChbnOZ/z3bs3PXegV4BYW7iPcepdfDjRSRtCAFHU3aJd3FOrQsi6E4kHFIdY2hahHpp
8CrgeLBcGcPT74pwvRar3XsP/8FJWpLHxqrpSlWyzPOew8brDzfQDCUX/J8kZ0/0d/CovF4xmzUK
ZnaRUqMCbVsQANcOdGCm2AcJVzzknBz90gZAw2uLWoX5Wehzh2+aN2E9kshVeinruySipfOciFLd
tzJ2Ax3CFANm6uBpjpRoXHeaxyiKz4hG0QuhqZA5q8wVN4R7zlCI5ANeXb/Ux2EkP2gvz6pGxngv
mOBDNwRK0KeB+zaljPaKfgJRfdAzT7HmZ6vZ1QYag+zO7EPRvF+Dau9vscPB3i3yAUiPqsfxQpI2
6hua4TKXyyNYAHamyz5axcwJQJf+4hS3brRL/Ha1BDoU+LIgVmWfzMAyt66kY+TmUVMG6zzefNzw
yGOsYKsId87OP3r7/UrpXJmLYHjdaXDNKDNvfqcz9/OwiNNFtANltA3fofTje0DPkDFFd0d6HnSu
8tuT80srXbFGDmAbcnR6dtuUWQjmMSktZ6hA31Kto0nMkDXNJ2hBBHEFk50TvnjiPq4OrrTxxDhx
daVLoSp6nItQKBaEOOWAYO4d/Ml9IRUJyWHTY2Mqn3STWPVK+nNShm93x2X8Am+3OA6u241fJ54E
McIJu9swtwn+VKNQ15htJznnUKvEH9p5ed8VWUTb0oJAgXrfac0hdu/2241BncwTMZTqUyN8djhU
HEc02rWIl7psGHsHvPse3DexDAtJT8xyM6dPhaYHlaM83YQiWmvcCl0ja0UAyjWsOmnKtxsqXZfu
TLP4bkd8gGFS5muOXYI3+RKGIEbiGe3v3HxXfNsLS0p4QPgqeW2ZpC76nON6bZz0nwFyiGrGZybe
k4RccMcDlbWeMsp7uaLgdTGpp6Hdw6iK8dAooHhD5A7ybit3ARkieQcN6AHUmt5DF9ipdd0dPS/p
sntu0oS8yD7M0byu+WfU17o9gLUCguwFt9xTbps1l++qTUoHWr6AthAzalTva4xKjTi4MnaF5die
B43Y0t8GKLVVmprYHzig2oodbIDEE4rPWp0m39DukDdXn7xAsZ0uigDZw8UWB3JMB20ySDJtIeHR
RNmNPdqsxOcn3u/+weLINtUdu9OTbbCBt01K3tPssKxF6bxR/Uyj83cImMQtYntn63rXFvH9vV1y
ZSs3oELv1EE1iddXL3BITCJ+VFNk13DcmihiqV8dYyQVm7LLc6ZQ75noRH0aLUUHhskrno52eJFc
d1LuE5YbnST+eZi1MHzAWIgStRv/wS4z+uOeHPUB8lRDfroeFpW/RuwoiVEufviqoiVDAvGG4Ev+
1H4/nsTeUdkdB6dsody+IbyW7+dMAmo+ndnu8tmq7uEBuXlGiEtGdN1E3xwini3srNl1Ki2NoiAp
Z2qJasE5p4fi5/A07PKPk3cEQsWoIyduiCf6TGB3DSQQij2VPpAW/JYxUC65ucGKyuTyx+4RwcZn
cxtr0daTVNdMFfcVDQNj1H6qVcEuUiGfAWc2FQi9OJexevmFlaLvIeRZW4TLUbBplU9EW9fokTVT
CedhghvYE9Lgye+omONhidKO0CqDZRP4Leo8Co2a4Lp71ECFVnkEH+5WMnMV8WjMVZDQEVWwlTqP
qQlp22GlL7gxj0O0jfdFgPEEU0zwfEohSFV16iyIdffHY9ei+qQdVapUrnpnno806eGyIw3kZxWh
8qTev1fL7XT+czZQxku3w4rG3Rp/einnA99VzSd03HymmokkBOQ8NdM7FdWaaJeqGaNPRGrwpA7x
cB0yo3V2ZuuZ2mOOOnYNCF8oouR3+6VssXgy8lpvgBg9y3JXtLZtJMfQD7+andfQasEe0vlY2u3I
5J5dO0mERhujWSPZWSeYKyuJcISEGo9vdaL6hukPFSkCAjc5barLJXrMjqHPTQqAdBlBiDa/Qcad
zVj6M5UGC6P3mX63HKOhuLeXmsWCytVHFInhjBBL+cwcmNNhCMuUrdEr89wYau8qCN1HtoiY14hR
MDRP4WizbAUWAeEaY8ZDaLYMfKkrf0K949ggS2W2hQwMVIrhgCQPc5XLhxqloE9rK8f2onMVvSlH
u1NWty89IqWh42/T91ahdEWRPibmwRI+uzGYh49BuZylH89R4H7Q4mTJPJP8Xj2oVmoyTmxAA2HH
RbIeJ3Fgwgvpl404tOCuIIO7ynCcg6iTM8uxU5rZqa+ooH7WTD7k98ITvEfn1+p121Vl3X49Wpfn
ONNJJysOTISQVFr0Q/cppUIwnDIxIYVUTjC2wTqOc/JEgsY7FETvcguDUvRmeDg+Jo6eboHAl3df
qwVK0tC8WdWJCr7YfEZqG//+vroStdmkU8bQGAgc/Gytg/8UiNjTmtoWcubPHMvakTJ454OBBC6x
1ik0dG9NQ0QNRKlOBi2ZdzAtTw+tkIph/EzcvipSsjJ244M4cfRZ2EVaiRgaNrqZoztN0k8IZ5nl
nHvEL50gKK8XsSo4J4nnp1m97MYy0mHEaGj1NQnJEZi6CilztaoRbuzf6ovGJLxTAjr7HAuSj5qR
tABebx3bZ/JJ20Ph9sD3GfJWm+TJOpmRN1WfiBWJMl091xhjoJ2IEmiKUXq+oKN71RPFwczYYWZn
QYR8SgidoiUkcWn7qpHHEzeShPTkPQNYMgQfJiK/KTn8u/jJUsE0zOddqaejUAb5VoxvRMouymYb
bA11brejgo0vlXSNKSjefYJAIslnvh52KE/WflY3TzdabzI9Ec8IyYnk0IZKKfDJBPWQkF9iflzU
MuquUGUxx2xoK+uHRt2B2p2WudEn0HAD+xXXyQnzrMCDrsjdlSTy6Vgd6hG7tg+wVQmbNrg6rbpQ
b+tjUBku56O3vMxNx1qatRny4IJ8/oinnoAAjlPkwqnQBixVp7Y9g33fLKOxtMRJd79PzVr2sBul
UA+0kLNBsJIBuvjVJdO+prhHKGYz+YLCnNQHUy5uWqviyTFG+zQDaBzG7sX5NpMTywazaM0mxQkp
r+g7qeBipqFRZO7qys8fwDflt+az+dfMERxCmnQV+0iAiAcMu+PeCTnSt+RoIOw+H/59Tl2e/9T/
MGBVilbDeRpo3H/BWbVFzPv7ldjT2ZU911gX/sfbjvPZBTaOuc/QH5pp0Rp7O5bt/Lc3On5VRejv
5PY/1gaysQGz82UjbslnW1aoiQSNxxcCB+mR34QF1V6D439TUnPAdJVY3D5E7m3MZgN+xAwzDZFi
l4e5lPwbSDq/EZr+T35RYPB0lg+oHRN//4yrP64+TaO5uUmPx0Lxqzes/kk1RsZsLF26MsuuQ2aM
mku4sSNXYRTzLglm5ooNDVTUO2MasnxhySFZ4w9tKwDORbNV85JdA79Na/gzGJtn46FTJ8zAgrI3
0CKHM2rSlfHoilAdKN3Zw9iZOrJH1fhTneUzifI+L9H+ZnC7Qf8XZB23dQj5ZByWiNXmjtmaanmE
d0MkVrnB5AKpl8gStKr74nr3HlVSWoOrePx/M1UKSLv0W8jtvEWQJ6bW6OZ8Oal/ycd7zwXFMJwn
jV/F0KE/+IsxJYo4X37LfEKf0HwujRC7IyS9NSi2D5exApUYHLdSwHBzauagLwwp+ExzWaW8My8r
CeWxXmS7ueiRae9TVHyQaSAJXWy1K53ObWYOPQVXn39I1W1w3i7Hz5l0V+CFDZItIrgD40+//JCT
T4WRkE08H8jbmFNmis6PFhVN5NFeZ+g4ftBLF2hBVMW+cxo4DSk4LuAlK9aUfkLiqzMNifnOeNA/
z+/ZxFVTSn+K9+wVBe89PrD0/sMeCVtpsppyTdqcH/Tb1mYJnWvQ78QKNIbVgjH9+6PObQdDHNwc
XIdQ9+iitf1NDWxp02yxNC4sHYURomKFZqs+iKeXadYfeZc9b2rU6kcdMvKL4zAoS5JYV5hfzMky
bnkRl0dMlW2pVoct3hLwFYB3Zmh8vG6MF04gu/muMd+Rkp1gz+3cVbZ3+Ux9vx9ptdEi6iRDTI8P
GrtjxRX1zCl0CqOj7hfKXc67UbuJYm6cQm+PM03+jR1XqfBs1OzbJBrxqtxdNT/Q7b1ZkiWwUOcc
8IJZ6j7bGpRlXmfruBBa81WtCn36j+rMQtHuyREGYFR1PjZ0/flfdQQuuPBJMy8oKlnU4nymNxbC
lmiDgBwRlecvybZVmP55A+6wmfb5aJEQVIrVuZGMNn4Sl/IfkCKxB1gwTqqszMIdjnicMi6Jtoqe
gCM7RGrKUCGj2kGMbYoZXMQv0nemYkwxrMZ4dOAGCfWXlEdrtZ1KFBqn1Imf8WCFcGDx+HLvY2/Z
Hb2U4RMpO6qbwwvw4aTmajAWQ3Di/usPA4SwlDZbb3CcYyJJPng+ZSHHHThWtr9oqqemss6elEBB
5IZdIOZNWas3HpWeQaYKGMNKH5KjbH1k3kLAgiy3nHXY9pbVROmq13clonqF/DY3MFQT2YO5kQOJ
q8exVtpDALTR35SDuuwxuPncs3Ssq94a2U+c/aKaCzoA/tHyhMhT1wg/nK6rfbPEOtwnC0cQGyb3
M51NG/5pLCWvg0YEqJhHt27xVfh+vwPrF/8JQ1R+Li1KuOS2wm0LuomZy4Rl3rBfRvVCsgx05oGL
1rTYysYuL/3Qit9lxpR8BpWX7zVR5VyON/znBIhGc23ZQJYEEo6cz4jjc9XcJAyNRcXrDoDII9q7
q4eUvm5Rsjv3dATn6Xlaq7XcxbVkKUkwjl0JMCkTDbjJQ9w3pwmUA2yXUKPNo/3DSsW0Ulx5pQ1V
Rv7XU/Lbt31ZJaZ+F+1G3nZF8UtThhrSXEhCETAkBgRu/nfuCKLCWSgqxN8V2SbDtjNwq2QuUGaQ
PF/H3xL60ag6Q7ftqTbS/z9iFiN/y5wD7XCYlCATlfsuG2NHntk2MifXqqVmXmWbmZOrRN+5kx3Z
NkgxoaBsCKPb8wdPEHe8MUVWeTSk1Nd9nWDtlWthKZvImovL6/Q1YERqbUy+fbiyBGZvzO9MpX7A
ikayTMyiCafdh1EiBA5xGpJ6HZtCtum36EN4u9gDgkmhz2zozDME3sj32tLZwy/D+wOXpaIuiF19
b2E9ibxsI/g0SO2WEqlvw1O5gFiQ8ZlZAiLm+0HJvrSHpX23u/fxxkHDwPK3Ur8o69i8P1dYq7qJ
Agn0Zs+mFys8iU/6ZvFr91+TXULtXKpXRYZ+Jv6RDMuh9/Gs4llqkawvkdKumeJ0pQ6Kn+4uB6nN
/SyO8Aq8MncQ5Wp0P+aDrt5+w16KR/cgo0glJZHYvOjE+YUI/poF8J6O6RpYDj2JR+bojPqVxGHE
39t5Rb37S1D/L6RiZ11yXO6dFwIZ0l14mi7B9xeStKppWWp+2nNHq7Yv90khW19NNFaUIZq0fGPN
AtMlBO32EO8WsswSVFgpakYTSUslo0cw6U8ZK5FUhI/GF507g9rnueyl2cpJ5MwqkIOBcLMKevr7
UhVd0W0N8k09jbKpWl/I6srOUFIhwR7lmizmuGRu4GGpFeNErp3lf73WGBsKkbAdNUD9w/Vttci0
lYC4qWnITcv/m7XML7DTkP2WhzNadZ2DGDLlpWt/b00nfc6VBrapnK8lD4Py1mm+T3XQ4c44T6+u
It6Pd1iQsGZzl916TiU9fUgFrGd5RWq7m4gOGf7mzHs9bpjdaGmppyBf0oa1hd+O20ptyrgPKWrA
3gY1ke/5PPtNzWS8SvOUc25evchcCaz1ZDDpO/O4O/+836xZxT6GSS9IF+BMW6T5Jxidi+Rwp1Qm
6xGbKYvh4RSJ1a7Vf1nc1gczQEeh1NCFEFqZ5kt75UoV3HTbtMhxZWUfp3IElaJh5Rgpjeqxj2PS
eTY3d4uMg3l6F2XmcYxq9NvMhY8hn2YDcgbRQnRDKCAhug1B+73z8QsmF7gtC6IMKRE1dSQSuIre
Fzw3oBmPKJiEJfRdV7uVwApcbLSEhtbSchwNpEotHC6yNwFauSAkjOXNgWaHxBm1729uz98yu4Jp
fh9azA/ac7QKZ8tarqKtJbVSn8uZqpoVcwOw97s9P7Jm5VC0HkXeSJYcTFXf4fNKMuk377SRRKfZ
q9AeuDAUQ+uwSbhZTaj2qFmEipnRuB1kdxudCS4PYzOVQOyGjzzQiyWeLM7W3MMwMaBGMgkOFd9O
tBVa9LHBH2+nX6gUJ6LA0nnilRZxXxvyNAEVh4GylwQydJHU0K/ccqz5plTGg6hkfXTGN9St8k0F
K65h8tPYYT24D2biz4ABdGs5WzUwd1dRl/3exOfcBMFdzTzCUsz6tpPyZkuoZhMQKxp56hXt0W9b
uiJhaheg0bDb+JXcx9gcLda2LmxFnAkboy8QE6OD7TykhsaeDx2GSRUmD407Z3PN/8YYXvdbNrZp
kUDzWUdd4xMu7LEQ17YVZpPd/3DRR9eSG+zwiRs2aITTqloH60LvQpEGXENrL9e40bokSVr2Z8xV
njpzTglE3Z0awf5gKMOlM0SIWJ5NHxw5lj7iCLvpSrTK4zMPl8u/PPThHnnqg+Jj5FQyCBVJRDYm
fuPM+m8SjjW4qyOGf/JKQPrWTAzOAYMHIAnoOBHTPCniLbZ6fgK5N01RQPKkhHKkDEpFPsqVfZmi
dMd/DM0aZt/pAQ5GN0Ao7p4y2Bqme6kb8tPtbKw6qAlSHjHCywWKiybPkEpX/1YGYQ97yqJl9biW
wWFD9fhZxccvvUyfWCfgZDPSGsrqX6Su35XMtfjQ2PvtwVbHyMjmHXERui8q4Rylv2X2WsfrZwmQ
gfGSsPlaQ09VhG7Wl+vyHEMjqUpJwZLAjRNTgGTabtDQDr7sgxNQjHl0h+BMrRDEGFWp44s9mkbG
OIsRO4MeP9ARVI7tmHX7a4GqGcYeUCtkfhUk2fco5E/uEj8hSX0Y9GmZL+uYv7bOSXlfWZR7Pyv5
f1J27WTuKcV3sQ5sSdKNGgoMgKDm8BtVpXn8wBNF1RSBZ8fhEZvm6nZ3WzGR6jNGy3w9BZlB5Cjp
sOhSntAIAPrqT3mNdFC7JXnU0sAkaEtiy0hrWz96iYKLOBcoTB5q7RpAAhLU1vS/VXjUrBbfG/yk
Bi/mGLXn0GfbkWgpetCl/b5U1wlI3i6e9XqvKdhLSEHTSgveMBo00RJFQ6Mwpuf28YGzQOfPzJBz
t9xKNZPPRVbVi4QUWKvg4YJ9R453tvm18df7/DSTF6U2tPmWIQFalw9xye06VtX42L/TQ9AdP4hs
f8umfnSKyc1BTv+8jFGKe9lh3HONsTcodJ6auQGbu7qkZT0+wBYMHkKLl0msOZJi2OGlhFTOyBYo
Vph1Mze1wo0DFzHNFfPSav2Bd9cTrjSs7/NpiPHSIFTm0yV0BzIc/MixdlwiwRIZSqgpMXBK5Bzd
8AQ6IhMvD/fAoiZIlOlhaRpEGWP58+JSsKUNwpWnH7/eqkEuoJjqoVT4uMjy4fj95DKlKnyvng7T
/9SOGKa5brqQ78OnLijepsLMPcsMmr20xrQER43lYta/TBSXLHbKLhfVwMG4c8Kv1LVRXQYApsq3
qZLKAWwmTkDgY9BcM6X1gtFT25rnklGXW5YqOIA2oxkGfEKE1fGUjxlIPoQqEyavuRsXncYW+jYn
vX3jBiqh1W9fC2ULtAQn6LLqvJ9Xi03kMYiLyjH5nZAEcqdajWpWMDRTDOFfe3mPYIwvSbBT1K+i
YmoenVTdq+yNQKbmRdHo8B02TvgWcveXfDIM+ae1LiBN4saSdc5q5YrarV4Md8zzx5CGmjMPAvts
VMM9IErv5KK5uDodd2FNqxA56c8h8o9DuyW63dOA3ETgGeXZvrc/CRssvjqlvM5KMuYx2eeTwiL6
fYq9f9p50ONyG2bcledPUpJrB6GEIb5dY8fuwJyQow/9PcZkhGjgI5xmaCfpFvdGYOenrC8wiXvk
jofyVYUxqE5m1OFJ8C5yBqYEmtHx01sGjlHBzs0P7cdzTMnOrO4K1MFCZlmvKxilRnUd9t+iooU7
868EH3oMM28LlvbG6+8qVKfa7A7EAmQAUfSkvsT4/FXpINP5kFFb0c1MZNsF6+UPLvhefDcWmSxJ
ESH6IPOgb2a5Z39sbkw0Q+f6Y2RwIIStF0fhseMKNq6xU0qBXZYXnZueQbX9iyTpU1OmQ/1ST8+9
RkiXXjGHYcEXWlcgbkFkV7f1PK6ygTn4F+71a9DZsvcw2U0t0o/BfAZNHB6fXHlFZkHylO83hyUR
6wEzoxRQoOR/GMM+4KpajZQyWzhFU1daGSUL4vMZRHlhR4W9ObkrcI9FjZbG0Ky74DN9gCK4/YWd
yYg9LNHuExJ+qpGdZJCcRUdRv0KswEbeMqaKrFN64e7PpMhSaAxNoCCytwoHazr1Mn83hoXCSyUp
VKj17qPpl7KuHLnJaNczsOvmlp4jcy3xcKzkCfxTzS0CgN71S3J02+CO0RrQGEuMTmu9e4oWd7ZP
TA3UpatMole3og86gvhmsJTGBal6W7rcwtOyurt9DPxIlX+MryuX4Zasew2pf66/XQkjeG/P/EO/
YFVmFPNHpWilyeuBGtYKND7EiwpWvBrKEOVBoQIJtyJ47yMt4+2sUBw3E97cdV3Ei3JtElFLQqs6
+d44FF5ExTqBuOgCPBXezk1a/Xixxc4vSFhHEh6krA0Ykjq+vsW7/cxZHyf+pa8NR63yIDHizlek
52PgYXnfdchwnaZJzh2pTcIgYvHZ/wSjmUKpuvAf3ycT7U8NnKiAqzIHhRwZd4scCkaXFtf1Skg1
4X90LRVDcJzT/qkF7XIXTcMKBKXNqzswXz3kNgcjpJpZcUgR3NZI2ucajVQ1fXBY1ALQLQBbWt4y
kKld9ha/BAftpnVtvNqIYmMAVeKnPwFAdWd7BFxuMtFJq2ZXabM9emVrP4FmmTGQ0AS61QNVKb0H
ersk3xMtDDs4nP0iB1YOj+02l5+Wb6zBLs5+zcUSXE3g8q9rniNgcDcSIenm02/yuQEZoSf4dzbP
Wq+Gpd99MsSBmzGWS6uWvRRV6UU74WsHtBLVxRTFJYI9LErIp9eVQcLF7xJ75Cje1jZQ83FabsTd
85PDHaWtKD7zD2EsLf4BlhwlnwCxA5VipS5SIwEG4B3FxVdXvSl23iqx3bu03RQVdYC32RsOnn/n
IJS79Uwsp+NvFcMxiLxU6w/8iBH9K6iAyBtma6J5FFqCcMynuiwDmsv1giT/b6yskV0DZP69ETca
qxJMbD0gOlm7ZWvUTuwtT08LFHhxl4+Jtg8/M01H9SJbLyJHM4oQlIpVaVNC1hktIOE57q1kRhqP
9CtgfnQoP1dNfgvTDvp3xXvl6ihiQ2w4+q9GjYXauT6XuXcynicD7KV1OdASIHv4aP+TeG9536j5
MuKVz1TpjQLIANYtNFqQDxZAGFGcSLPVKycmJrOwZ0PKM8R2Yzj4I96w2ZKozbQ1PeqaPiR19tID
hcLmeOiiC6vnPo4BNuElaqwS+CtxdRQZHCUhctI8HPI27lCXFdqgZnkAVxfJtTGY6vXvlQ87RMii
3qN+G6ICLwEnhfvYNAXUb+fTN4H1wtgv3KBj+TdkvMG2cCDg6hzTmwj0TDHKW9UUZlE1CEVOnMER
hOOn03vWHNOj+Ilgpyj2Uhk8I4cZCl40Rfovl13Ck7np8USt1cQtwbVtSBmK2NN43v2ViomZzQpe
UIeVJowOABbiaVUZ2ihdeYBVQjmao3DM11ajpFuTYeT0MNM4UsWF6tImzaFq08L76hoXek7WUQq/
ySGoS4oiVF5nnkf+CVRx4QHRnBXc/S+VYqWZj5ltuiRm0MgXF4vF+dItkjCnzbM9xsZ8s6qqZX7l
ETRc6/dsZb5U2Jam8mK6JUp4l25hLE5TIHW+ABT+B7uJmfdr9dLtNVE40EEtRkWkAP2wFaciQqUB
3lMButirNLmk5+WsUH6PfEymChlmOXx9zowXR68/UvXEjjVSTbRs9l6nvproN9S+GldKld1iImR3
Pb8nYTvtbZlMvbyy9XgaXtgexUEIxD3o/2UOVakhL53uUUvSHtT1QFsdXv0beaK/pD72aXZZyvHz
hgF50DHjQ2CMgTHRH0Px9hAtnF3n8EnpS9A7C8RIL9qaXAkqWu+P76Lr7u4eiSTg07Pj9Kv/Mylc
zc2VCcKJMYLuLYG9KNQBRGCbfij4NQgjSSGSrEmI25q24grCPBVkhZd1ZDdGZHtZTVBzYMbct6j2
DZmrGi9I1PKjVYqTLvz2H3H+SdKLKrlhOtT0GEYby5gEonrnS8Bg2QfF4a/UOL3ll2DxXCOZiah9
2SnOMfY/pkiOdZfOGtDqGrJ6Sx26/bzNI6vaI4kZvTtwKbYf27Y8Ftx+i0s9XKnSsKlyrlU+K6db
qU1/qMCKuiUgOko/YvsjhqFNghe8Xw2wMgaqCzG7lHsPxbJnAf1pcASWC2NnzCOzjKWq2RL5ZOyi
US4N4P77idtyA4ByFlh77OWr6o1Mo1JKiSZTZfJr0p+cZYnCMFrJ3jftCqcKVjuYnbFvCWrx6Sf0
h1LQ/PY65DMU0ahTaIGgmtJ4B20gHwTkjwJvRnP11crEilm45oCQdIDOzyYpF6bMyF8zHGVwGUd5
hbpIRw+BJVQXF0ovhoHRYv0M8vNV7g5Fz2I3LrDs2MmYcoKmha+LKThXq+GdBq3mEq8QB+3wSbVJ
VCmeyKY5KWcz1yQfcLhaicllUpR5ypB0xtGExwML5lmCpT4XaVMC+6zGMxvGfPluhqxupsdtTFgg
gw05fWIGdfl84yI1oNEpwBJPiYeEoI9Ok6RYLukENdE+dKm4sPt34p7nIyP4r2p+b/xM9O6fBnNG
gReqQQzwtwPBPSb35AgdOYKYxU0l6hiopQnF/1rkTEUqui/ttXpYMvcDZl1lAIJGQHGgXugvVSDj
49M8LE+1CASz05mkabbr1effwQWzWYjQxzq4TKjoRnSV74bcJPLMC1YfObtIJR5iXwFTipGf2cap
B9gwliRAkTZOxl9T4Bvo5Zu48YgoVI2pra1MrvYzMYdV0fKZnVTCEu+gaVSmKI6XvPolE7YVMT/y
Ak7PvK6EiBIeyQGQq5BjuuBMGnfu2Vp0o0wrjxE0MR7Hr/bH99hzrVj/u5rlOMKo4lB1If0JgvGr
QdupUbiMBgt/YzO35VhWJIru+6eAgwZ0BaHOZSVbbVXq7ijdcuQUvB6w1WePO9QGlczAjKvongD+
z6kDzF93kRw6CFg17f5EQMNjDGT/YFKPSCrQr6pt9En8e6MeEY1yC9R/4eaJTMoDgwC1AMu/iovo
ouF3MaDAJJ/Jz/DOq1QaI8NGiIX6M/blkgj8RnAp2O0f1jWSMT01xSJKzHcYNReiUEGB7LZqPv/+
QqkfW89+3A5HBGsM9SNenhClVIwVOlZM3LxVQD+GpnBQlSe7h3gRrjo7A8ad9SC62jXNJvEx4/pf
fYyOfVZCM7s5ctVBXyXn8DnGIX8NOb7K/WJxc5OSP+2hQ/A8y1QUUDnTIQpWvmOtuoCNLIffQIvm
RRWxq5yXs7aSDZYimUhrAdtSAer8HH903w9dGgWtQTE2ZZiTh6jMRCEmkI+tvzWneIGIuOwv2Skd
j2MPnPaQUULfqdc9DqNlMJNYE5fQc+OEhWVEklzdbZDGV6gk9OhnHXFspVPYWGHYxC8ALL2a5UeG
DJVCqZuzU6tjncWS/KcZ6NlRwIQUDNGqHU/T1FBNhpmYnlS+qj5o5YxT6i9N98n2TTatZsoiGNiy
wGoWrBahqIcLyPqeZVwqA/XY/2eRjfti+xyF9a/i8QvYo4AvNsg9lnydtFzE8hqx864nmg62Hf1I
tG02KLYjGsGGhmRV5b+bJQNa/276gJ8I2Z87SJkomhhBa3vpLreH6huCnfscdpilnBYky6wVczcA
6AJV3titBMw017uAdQKS1nQC0oe8RTNcglxV2ip1xp5t3bvrZP4DoMB1tQnJuCsGaxYGBwxYLTE+
43X1vBeis/iPev4K49E9xw54z744JghdU8e4DIF8wOuUl2I+P84beIh/lV2E97YKrE6yrTzeMq9G
BOGuJII9cZAv5OoknWpFSM9LgXUb6P/9IxLupHloDSutbyPxE3+eMco/FgHzyMHXhjXr4uQEXE3l
qOeZAEs9KcGuU1UHXOyBSkD17aeaqoRzMaOmEcd+wNiuEcWaG+D0TKcdjp7JJ+1j7AGid47oQGjK
W++2YbVxgQvrN+ushksNMnjTSgk3QICJNvc+yQtAvCOiDLC9kBcW6i/LhR22672PmgRZ2lVA6twL
iN41xgd9TFsfAGz+l46ocRmMAqbWNsZT03qcFB8OVsFri+zoueMH5pPX0yArZAUXchCzoiYCIn4a
41wg/O844NV6lU+Moa5p47K/9Ua8I45JvU3Kt+4mAHQnltTQKKRPj3KbxNyBGu2adLzHf3xfbgt0
cBWvAAtmbtxNZdxr53T2OpqKTv13gP2/7yL+/Pt1prAHVcfNeisfsjQRCbeKdHxmTCrquWTmzW5Z
1VphvE1kDV0y+6ktpJWzcZC1OAs7PPISrtS8y5FBXNrtl5SIFHb/q/EsbJtzL3toqXYKvj7PI5kB
NlqrizAcGgqcb9b4TCd3Yc7UwOZAQ7/Qi1qOc2zN6bFejH4Y62DOnx2Bp+rg1bIT2llD9rt2TWKj
9AurH1+E+0KjtmN95t+zHAZIR91WLpe6OHW75r5XI5CR+PzQH5H1ZUjLJEK473VFJK/ssKuU6/mp
AQy+lZ3wCUIsUK6KHwKOr/LZRuI2p4IoDCdx6Mx+f793grNz6YJ2oeEL9xarZ/dHUBCgrLT9wbI/
dn1X+0fAZbmELwGD0BlHCpuq0xkrg7Xjg4feZwvIAD0K1Sq2Lp3/+AViInRuINDZ0+udqizJDdbV
NnsPVfmKhZqbFY2yv2+PSXJCDmhLQN3h9JVCzwZheHB8oir+AiZ+HRuSa/rzumKvcsgNBYVHr1ko
EL06nqgk3tgUsxeyAfu93gWHIZLvR+EeLFJg3A1wY05wYKxk7UoFqM+8dR2tJeH9M0CchwiMkrzY
tRzv/5w1S+ckecwej+VjGx6a70WfvTdsq+RTdt2N9Lsv7/dPtzROFpNDCihaoK2YNkHJMTjIWgyo
tTeGbqzRRCT1FXrVa5p3yLeFfNWFa3Xvn4A97e++2VOYR+SnaweKI+hU1oxUO14NbvruALEkNFlK
f6zi+2tgh9F/ZzZd0E5yJAZzGaiGpbQ9IaqLpa+78bZXr2UzD2Qgw2SNb2OZNptxsb08WKVpunRY
RPFUtuUlONlB2acAA55htZD5soAT862gIJCYsDs6cdBgpr3GfrsSWuXQ/BrKJU0AMCdaySyW/ewU
ZWmWRoI30kqOZDVDq1sd/2cm+KJguj0dFTDNjBUXMBJNuBErF27ls9X91/Y3kuqDu94iVTe05qhN
AT/ciToQ84heM/moU4zu+LLjzMn7RWIQ/oOBmbLKfR94tFVqGKOfVoYLwjW8DSanisB05tg7dQeq
0AHxc9UroeZwOaKQUHOgXeBs6XwE8wBZ0vWy6KPUCPcu4sHEA6gUOeKek5XhtFhTmEMd0rn4bvBp
6xnSQxnVdKw6fWBEnCWvaCSwWg8XJkljpoXHaw6wPdNojM/75SYTt75pVyxu50uf1LodeByOpG0d
FdNIUIjb+prqQATdqiBXK48pB9fxfYJu4W2o1ORc7blApHGMKaKTct0Beu6HRhZyosaYoR/ssScc
05weTCTRgE/kLA5aiyE9SmFrDEGyIMO3yiQjh5EcvWk4+cJQmuMSzvoTo1E5xhy0+wWaJtGIaAp+
8skEC3DrxBMaOnD3Lgj8kagm/+qwxrnbg6VZYNxEDnSpcKDWP+D/mb64q/sPFNho1ZQM+9iPKFxV
DRf1n5yS6SyX7Hg3+Bj0dTSD8gdxtZlon3EeXe43Jn2K+gxdCSK2hk11qvr7SJjl+Q0pEWSDPTYU
7KBKsJy/+HiW90k6hbsehyu1cEwap5MB1XFVl8aBtCkY7C6M01gVHqhZ5RnMzrjbsia+prlOhqDt
4KEUM4iNg6mWhPDj8uAFcNtcPv1b7bvoeFijrLNJLIfhbRF+SQN/unwJGFMlw9yM2xylPFtYgG/L
o3XnLJjB3Zei24Fcf6Wn3msmDIXfqrR6o6T3OH/TTVUcUdT6vUkMlpFCN/1ih0iONCxcxIIC+g37
H+rM5+7zuL8Sw/y+uaZkXmAXuxItWkQb5nbcPDE/b8payDO+CPt7lK2LsCV0HVT+GAzX/ZzbxX8t
WDApQk7LOmAKTyG1Q1XDTaYZhaQpHwsP9GbQTU2G0eELZfcpFiyEMbK8HShw4ofyrD5E8Ft27vQ7
0sf126n+EOQuFdZHLmscifBu8eUdpRRp/nGQJn+5FI3p1rwyHHrGN0gmoP5blz3IJwzQkgOZxqs3
y3rSteAHpUklL+9Ha94/AbUNTpAxR7vjGvtmt3u7hv+d0xD9Dmh0JwW5zMb28ibMIKihb2D+MVfi
rr5cxZgPbNLwjujwEaQD+W9WYr8tM6vcLrlRmwb9SMcDnR1SYWbXJNCrevA0/xX/8QKfGNmCbKsg
CMzScmOr97FtOdmFFpDWOFwUqGbs/RTTVTUmw7wCExyQ9gXbUrA9mfRMNgBRol4n6ksg80xMKo7z
Eqzu5ODxy9kkjn6Qzn8T4iX9tGEuTbXy5et4am5Grm3NddcI/J7ZGLsvk75no6cLBQTWD3rAEJ5Y
e+cnAyn8+NuJGAhVBqU3xmJXGffS4d+akgOXCxzs+oKSgpu9n1f6SZ+B/UHJrUNlImUcfkvJHAbM
4HGyiFPVohvGhJ4HyruhMEu3xB96/wafBKwKHuvoX8ACFoxnYEO1cBX8SzXpH9Ma3WJLYFIdkhjA
MMg2jDIyXfapDLXyEbGp6gvoVPhMjEk4RNOhz+zy8NdO1Ro3Dh6IH8BTn1vtrsThWXvGBOA6O6WC
DWsh8+7Z8KdhPeaPnzAzm5ULr29Cn4nrgkLVZ9upPSiF4QgXXuJY/CSPA666U5boazOL8op99Whk
b8MOADvMXXSEMY+fn6abls0oWrXpiPCYQBEZPN0x98UbWH3irzu1XUznnRsw3MS7vpMPp6kL/yLz
p2BRAcjHs2oNGUVbFMmkv7IsgTbcnUmZpAUAEBbeWFUo1rRdEf5d1oLmORkMZCzYyUZErtMxEg9w
T/lSta2maGQyXUp5OG+6pALdjlYhEaDOJ4VaRFYBUq4YhHXnkeo/hwZvHVxcLFDKUEVkwF0YxvEr
2rI6caNGk/GYxuuEmYO3YU4eb5byzdmvv7/h6VFCSYA1w8nnNMQpPJ47iO4r4WpKE8tE0Ep16KbS
NX4a+cxWAUfJlJ1ZaBSkOoTCvwuGCtOnzYW/cpxenlDEZWPQkDNa5REgAGIcy7lsmarNFWmLeHup
XensJj5la3J/z4IyIp3VaDx500uo0EoruRzwGFThdj2Uj73tfr5DHhtottu4BD1s0FcuitoLst7R
q9P8hlWx40LfUXEeIeF0ZcpgMb5S9wm1jeg6efymOEr8HMtiR7ztJp1iSuRhGDhaZwOQKcJWPu4D
MH6rIMDI47gl8lUb9v6gNs1RXKg4fcJsU+O2F+VDpgC/1ut55pNcXNvQgPgfkduBgTSf8XLl7pwV
L5/HxMdUDwObMXNZbd0Hy96J1eU1F/u03/GKHT21tRIiYk3HBUEPdLiDwYYaGcYv17j1j3cfK1Ha
hrmXb0pE94xpJ9eDC7zv8ZmNtKfHa2XxorGaE9XXwzrDz/btPK5usNj1ziZj/U8LRlai9B6NiHiO
6RBLkxceouR25SLN70UvPzdEM9BKbX7arxUuMvzMoGt286SDEHTlco/tDlC0iHT2qz/AkhOrgwTJ
DpW2UwnkptBaosfz9IGZ2s3T+KdR4q8lnQMtnM4z5fJIgyL9wm6uAGdK/3lmkMZGAxBdYYvnVA5H
FSgdWQAGFQpr/TA9Fk9QmGS8ldiog4PAsvDiKyQo+mxhRuG98AarR6O/gVugpzHzLo9TS2w5N1MO
7VadmpDSyfN2M6P8g2KKG4rX3lvshiKVqysGD53ufLfVWySBLzcSWOOPLNeMnC5xIEJaz/RkOaan
bV4e+i8qGoLpQ34Vag9e/sUz5SAFBRb8UArW1pZoiQHf38T1ocJ2Nm1La1f4CnXUvEah8QduXX1H
OGR98k2ZAyXib7oqOOgqjaOMKhY+tSRqOzLGYuzKpiH0nrOEVhebsUQdR+EdR4uEmisrq8nlzHtY
3aumQTGgNUeF5u/P4UaXrmeCV3jH6/gvSAFdxy59y7PXPxl42VxaUtlKcWC0QkgdrQIpEr+c58zp
jV7tejYtlfJ5a7cATtBuE5ptmew1lYImsQJj68IsluiGO4MAH5AaBOemsk67MBfSr1TKqUFhjFi5
abo6eI4om4hB17FR1ZQwgWzdeGjz0RS9CX1U0qHBZ6HIwQxjmHdUzrjd+a/AgruxquHp/YMTnAis
7XILf4atEhLzCqSW1mDKBG1CV3WcyWMF/lDC+AtCElPwoG99pLUdAWVxYEKuyf4dSMJeR5DwuGla
rqHnjha/7l/LLi6Ou8y+6YJZ0lUtdOP9fSkvz/ZaPFx3RJF7e8xN86ry/xulHQzgBbwh6QAgAjC7
3SAGp+CJ3lBRFxIStDYA6urDPxcyIGHQtYE4/YgpTHY4fKQvLvNObuRGHK5Y+SWUcAfvjmqtDCJc
XrNQE3K8+wE8yE+rHVXKI50ib2akk62w8uCxanpu5rrEE4Kp3DDRzqVf0dRZ9Gr+0wwkWcfgTYWk
gkVNwytw8b/nbyvtACeBUkJEEuVmvGeKQZ6yMgiCJE1iVE3b331RCoIayFNbRjdCN5nQeRSvK7za
handZTmW0adc3cUqTCnGN0rs3niQ5Bi9cXpeYtUEaAKo13t07kkZZ2/S91xM4sHyTbKBHHXY5LWo
sQ+vgHNuR3I6vN9uQhUqCCIrgIRJQiPd8uvjL3MiceFkzMeLyssl0mXKOomIBmrYyDYOpNuAnnQ7
DU04vKXCA1neu9zOCgITlg3BYi9/Gbe+dmrKw5d3n3rKHun4UJ2X/u0KoPfo1TrlKNiXcFVgkUkW
EmzdU72Tru4MuYSmcRCzxwSp9pldIBHDO5d5pXdgwKbyrXoNd0pCexy1rMH7f8Ne7YQsgPDvl3LF
4kK9DfeuQ+ucZG/pUyMlEKzwI8Z3BOLfUSCTK09t3WJD9zPksTaQlWom7P3bbJn/fcLrqn4vIBzz
9Foz75jZWd55NuErAA0etnev7lOs1q6SrJ1AMCNK926sdft7JDW2K9SIYZWmZ+eI6Eh85tOSYvPr
mdncVUg9skM8KbjSOATOo6PAzMqo0QjoFf87EteTucD2AAVUNZfsfDrQbqu/N2jM8dmfmxQcfOyv
FvshVVoFCJ1hH2FVOtzSOiltkwKmdJYCYdJoIYVlzhj3dCYVCQ5NVdEQuS7Wt/7d9HhAv/tBNeKa
WgvzOt+HBm1jKixP5WWhH3LBVii7P/pkmccslCLXK/g6ERg25toW5E2qLuJoAlPRq1rRhM8cXAjv
kiwcmpI2d6VpYlYs2BLjHkzsOpXuUrWcAfiO+PKSIQAexrJgL7H+IhoEVlX3HVMZcsyrNe1hWx/t
dYdvz5arInBAM4HIPiOf+GmtGJVrFyUiHkLtawMi7mEA1qIZYcnJnbrPBzqoV586DSfj1stG+QtR
dt5Vsk4Au0O1Vru9v7gJBGtIkQyNqdraoJOdC9P6fSeFXk/etqcHZfIA/j5lAv8AQF/wN0+jll/v
zo0gWWRSXkdLj6I+iyNbohjlk0JnBxu8k63Jk7SKuXN488lKB/Eu6jNz3mrl8uUlQzLImGgNKxEN
8CMBn/8POvbYZ0SCgTs6ZLcW+RlvLBcCigRzw/LYhaOD3YJegwMBRJ0+Q8s98sxDPil1JmxFgP8Q
KA19eNaEEe9z75DRmmN7gOHfJ6Ipc2ES+Xj0KRrxpP9yrSOCCygfX0BKU2yLwia+spL1YhDE0mCz
WAmnv/q1cbM736WKBlQUxr0JAzROTulO85qe4l25q5qzliyuDPQfDpyHRh6Ji3DB6Yga7ZBmR4Fc
zpkfVriNSB3V2t//wp94BdMeCUwkh0N3ccWwTcXorAyNDXqLU4/Gn0Clw2VGmXTfutV6D+Vb6pNU
AIkwCsHoIDPEN90LC7ZDJafyJIGQIii4zAQkeXIlgFPw18etdK1e9Rv8EbMREluLK3gk6gAVhBni
h3NbmvPL0R/2AkRdKeOUqdK6s0ASADf0MaatLOeY1zzysHNy4C7sQWD5Rl4ZK08SrB0SfjWszs1Y
PTvg6yoKkva92iNkx8bt2tP+XxJlvP2ugKxrfHPW9LMbsgdiVLoXveoSJxTmjGVX0vsiWKtR/6f3
TzF73CZFjK2j2hZDA7wXCN5GvBLbWOM3Ks031hS84mU2cbBl7+zgx8LqipAPr0MPCh24BzEJetHM
yTEVsewy8v7z5M4N6H5MwdR3OEirijXc+I5msEUHDgstiUbrcaIQBdJoWD4tNNm75TjDbUqKlb69
r1D5IKzWIrVPq7XTr4TI3pTHlNjc6b3RBZgVwkxDo3C2VR1//hCPduE4iWndOLb1EDjsJpDKmc1X
HV6lODcWpD0m2r0KNVxIieDFxBY0/8hOvbh8SPynpl5qeC1oEmi7G8SmvD3vm48xBLDd+cGTjt/c
Y7C1ZD7K3fRLwRlQG3cQlN+qb9mhuJsONjT5K4B+9TktkMb226s6xwFdTItZIDOAAlxSfoE40FOy
7mj8znz9lqonMsgMNbleDk1qLQKAmybKBEXPDD/HexqgdEfjSHfZQia21iEpNncIuQCdpmOo6eNn
iDcZdmyNV91fjFEOTTr3p/C9Qdr1MdxC9PeNLxXdaq1baadO4QkElXBZgTsMEzvmIjuBGSL9KKYi
a4ZAu1X9x4UDuVeJNQ63wGkf21mqtx7KYwj7kZBPScoPF+68u6fMACqlGcWRnVrSpdL6ABzhlNxC
jWmed7s07LqFCJ7ZeG4QeYmqv5ndhXSph6kfxbf6jkflYLbmkm7YIrHoHix+ziwC+LH1F54AXHik
1oPkn5bWZ0N8np77XQtEKoStmn7q09lFoVjVl0R2RUf863AWWLEGZHTcLhjihXklXjAQJA7U6nGj
qxCNSsDM+eBbgpq6kLFnw0rIrPdgzZWucqMaPT86qxbQ+uhjdW9IMuWUgVCfs/VlcCtFaHpNPArx
2QjpxuqPO6SlaRN9In+T8Mewl1f5D10l6km1y1yPGW4id4MpBeYDkG2V/KhrLHDgEdqzncw7r8iS
gb7UTrXdNRcTRip5+oQGDET3d+XbkEb4NMm9GrAyb5zFHVpg99IYOjY5RCjdrXbJrbVp5O228iun
ODUa7hcrwkzRMbC4YDQHrlFJ6Zj54LggJB9VsioJaskTMhhk4o6dc59ztzQl2vjkd7xErlPUGCyC
2lckRmaqnLnvsborNc5ju12DLIVsyK1wLMmRzF+/Ji3oTERjyrxfxW3Gy2l2uTZXvkd9nQSIOWg8
fKCGXZalRrM0DLzCeg/nHjJCwEUhlz/lNEqCW1K66iXrQZ/Hvcbedt9XxWmG9qXtNXm1NEzqae9p
fA3I3iPid+9FpPxbnDEsjUL4uw1JwcVwSMRukqLzK5Gtix6okXNI1HdMpZE9dIHnxYqfeNxk98Ke
rFneFQ5g9/N2EBH7fDwkXT19QkNZAQJPWWO4PgTHMkHkKn/3KBoW3/Eo0qunVbSMoh7Anc1GY8Na
jMFpvPepKQehR2Vz+8G18RayGr9aTVpBWUqc+fgDjxME0q9qXmF+gDLlyptPhplVb0I6yMv33/kH
/S/osVFc/sUaXxsqhuZQxJs7vlWfGh+uGLq4yq1vltFvtkEzaC7EJzNjhtwuNFjH3dHoxGjGL/X1
nyz2eh4fsSq0FLTOjuOUKJ8Xtdoitfc4tCzXXe979TNTYS+FEI9dBK1o6/eYobo3xzF6HCGWMqpj
+TsCNnxS/5ajm7VK76sP3seAzUYotl/1Qhq8DdgnW9ALeHIWDL+VPa2oCey9+SBjmpUfmWRAhYhr
RxHrifqqxWSxLLiqWTQMJhszO10Js5fQ8DKEaKmmCYAX5dRCNGszFYNMVq6jkyYryVxukj3RpOtH
hVPveWYxH4A2jPd7RJi4qsup1Bb1ZG8iiekLpAbc/6nfpzGoK0jps0lkcvm3ZufoKSTO+/Qpx8x6
PV4q2u+9Lebk6H4wsXpOYHhu4qeHzUx5nKNy4XYOcLZeUUAkC/RZ7MmrDe0zjDs/ZQLgJ7We2sMr
K7sw/3veHO5Aurmu1nfmdVa9f2vLPmONBFCv9TYZRKUW9M+aGlYdGvebpY7CAeuw08Z94T3U7Cg7
lhlPRiRc+Yh5PavsXHNnlJZLJU4vUd30EJpRVVzHfoX6/3BOrl6b5LK4Xw1wWZuEJWxLuBn9suou
mfT/RUS2DN9oajagl2ZqfDZtEP0XzzHZyN4iTxgzsHY8KHoKs9eVHFAezHzyOb3jH6p8/tz789Lq
2X+/xm3oyNBf+YhESX0iRZHmK4RvfKHYpVU55xvLyti+IS3hkyHwVjPUk22WaOrZTR7v8P54b1KK
ZG4eYTqUm+thm5OQ+coQwKwEUs+hime6075AzhDw3ogQn0fvEb9LvGLBi0pmXZqYZuvoxaYfONdY
89H70X+29tXFSRSFArwty4WNPeZ2XJ9SjXZwx1eGpHaGZBAH7j9f8g5QZeIykCTIRWjADLRspqIF
w6v9HLtiNjc9mIu0wdKBPY7gGwSofdRmgjwuXPd2g5j5yV5BxTK2jIddEfS6Pz0cYKtthR1mKrYF
XjRsJpiYxvgZXXOl72VmSZ/plihjC3KAAD1cVsuLIeaYx1uzsuXqifaG0KWE3l2JxDrdmT+n52+9
olahlhS4QUB+jPaOy5nYtx+K6VrPt3W0du8oH+WJane3zzcmD0YTHokmHAEcjr//85L6WO9eNYSw
wRBr2JyS0s3X+nkvY7WRRzy6hiivkY2wTbV7HHzbrX9StcfwjK5Nff2i96DN1pc6n/ckaNRd0ecu
aeoyW04KaL9rDL4ICqzj/8jtkEXN7k6aYXThoLqoQ9uUs6NfQcRq8zHqFUopTqAKD6RHNUkidu8h
HPCQX/UFlnKZTle8AtEaUZP4L88PcyNJbAOkp3KHj3BYisBa1GaqrTvIrevZt4FN1Es6qfitrdfe
YjMiawDyiv+yBA64FbZbKNp5WCOkq1bQEXX7rof8csEzxrQuXVUHfoVR1uN+uYIzeapw+OM9z3VN
tu327j3JwULJdRm3uc/E/R375XcC9gxH8JwkeDkN2Y5c44mJzDwVsYNlQO+eAvaz8xab7Z3FgNWG
2jnWnTD57h+gm4eIj2R0g5aqXM8nC/yNlQ3eyZcLKqi7GWw4uXans9qpDMAA7LBL8uieJWeBpFCP
1N8X1iPnCe5dBmlV6mlIFQ+VJVfndiaOUkOOxTze6PAdceMwXspEj++eDpG4ulbQJVCtjUfJJN+F
bW7yyuVr5p/9csrtH34h2QNGU8t7cPlCCPaxBU0d94E3LsUs+nYF9cn7YjGSdXGgtLZ4l1pQY3hK
uRE4S33BkvqcnbTDw1f58jBJwZF9p+WT8DPag3lNxxiNg4ch3X8gHAJpQU53nVbRPTErHA9jr0QO
aTSvwgXNEtxL0GoVTIauJnERTX8nW04iQ6L3YQmpIgWtD6Fg8StlDQ4Xy8NywK+u6ukVlbCjWRyU
bKKKJ6XUXkWScpGg9l11MpmC6xu+VIC+nU86ubq+uxaF76Cjmtry2vX0XZ8WLS8jCgia2NfIHCm8
nR3GH3BwYwRoJAyvLncnWG3mRo3DwSusHeyVsifcJIQ+d+txL1UNUfWYuHZWAFBKZDd0XkF4BYuC
ntPYbgKYAS6g++MBerzSKviwWAjc0E1BfRX/AvyYwviklWYpQHNcGrhgnVXbW7GsaufkXY8dFgej
1yW2wl9KTlPl3yWWMzOVmrYneDvHNMqcY+dI/EqzOdjdT5096YwNgeiEusntjF2ulQsm76h9sCHV
Xd8z0Bl/TJioB+Dw8pT6ndcZG83hWeQBi2rOdoYZ+xetElri18DGbY48IHrgzCtnQmmcP0lICUvs
Lvnl4iRs5xSPgV2upyZZp3mduTmDgJMxLbIj2spdmBkdERBc6wcs0fZKX/WE+fYF/27uZu9AdT5r
qGpWwFWgbWWWC++nEgCIoExbs4aCHVej+Q4RMsXo7X3lVTckW1RxlyfeXP0lMUQcndsfdXh3c/4g
6Brv5KuGAlxfD0AHIs67I6iQ9H3lz6kAhvHZxJW46TKP7fgFTb1Ti6weXuc3PXeC/MPIYtyLupLg
6mmGmKfz+1tSU6hDRj/AdtT+3l4fZNKeT5MYJDTs4D5punD+cb+r0sfPtFrxOcB1qXA44xXD0b06
i662h1mcnnV1hBGQEW33Y110pS5qZRbRIs2fZyYsSJAr//IydcWq9pThZLbyY9LHGZ6LIBWJkh7c
/fi65UQZrS3g8mH7bXuHb5eSONeo4qzmzBquAKcOHVj+/ISlXFBnPI1rR8nrMyr0smH8jn3esKV6
aGo3StJiytXmO8DgTrMR3eaMG53VfefA2kLP765JLxBq8rjThNCni/jIv9eQrIIjJcRX1PuqBq+C
5GaObR9/HEmffp6nHSsUJxOAd4WQ4qts2Bo+wM69eLJpfYnUDqGK8G8oaGLJrIFpA4RbrcpEzeih
A/yr87rrpaYt9vYg6qaWCtDfUcjS0qei7fL+MXRQOTeDxFS17vA0+/jPVYHcohgyjZBkdVbsBw41
FkEkQXa3MRFkG1ye7HSpnkUG68eu+065QDThLrqhZPo/Dpn+/9+FHdIp3pvsiiOBRj3kW/70QKwD
Mt9StnFCkIWdXGNjFSb8Hg/ZwXzXG208nKSkE2hlU/0xFx/MWoXuh8CaBQx9jiKprwO+t9k4MJa7
QUnSrwU1Kj2HIvyjARJdai52dcvYEr+YccTWw99Gi+GOkFwXkrzB3ovbxU0ASi7dfMZz0fmSTKcl
x74SJvDwvc3fOAio0Tr7dCe63JbOfQ/4hECcyjbopLgsFYWF/coB2h27AQKuNdU6LU5eBL4innzx
ys7IsaFxqgqjsUopAyk+beZVkqR9rq7whNhQ38lQ5IBGdPGxarD0f6q9ZN3PJbahAZcmDLLn3rQ6
1+XVX2ck4RJF3QHAbsBuyOacZelaMM6Eyq0PRbL52aVu2Wx14rv8Dh5gzKX3dKQtiaTuN82FONFw
sWvW8Tlp3/JyxWz9FngczEMIlIG53nRTpP77BANNw0aBrb+E54vBGSVa0Z5cex6bTbtRahS6rdkh
uRUsJnH1qRgqe+nWJqBJmQYUl6us/+3ZvdF+xsifftsg/Pu6fEYWVtHsLM98utPipjWrdofaUu8l
cWA3v9Vtf1FJgL0S1OKAxcnC7R/H+AbesSbPH0C3YEKqADl51UV25ZHsRx22ilmLeMu6AmPR6ktM
qx5Erv1shDNQokTeXiwzqj0VeoeR1T0ApSV8HR91f+gzZNn+ZtNjPtXJ0uhSj2GsWvzeNcEetwjH
5o+i4ivAl9z4YlQM7Y2KNqeQqB34hGJfDS+k3DprFJANG9fNyVKEd/meYNNWbqgbzMMkUIhhyFnj
Ue7fbnf+8k//dU5ofus0kxdEVe6D6/jPPjNt0foQKzaQQ76NHr7Aak8/LTHxt6ElTf76TCd1bnAJ
AhpPPw5+FCVzztLipHnoGsbSH73ac3VXUr540Ytp9wQT09LcCL1CXoDlwsvRFy3qedutwvRyaVD0
EqZFGz+xn0YEbNrxABVGn8Xx6GKDC7Z+RsIk5/M5iIbX121mEI92J7nMzk0FrVBWKTJdUZRWg8UX
GQI3tIROjs35u+eWC85ioQy/x/ltqxxV2k75aFFkiIhMjCsmyNhyZX5bELnXSmea8e7a42IR16lS
EipQEhyHbVjAt8A3SJQG5wMkzZE4SvDnQmAatqo73nIilXG+Mf1LyIrKpzkEBeETpHlHw4NvKm+Z
I6Ug8u7CVL86cHAPR6LuRHisdPnfwFdBSuc3P5IyTV/tjJEwxTZn27E9u05Z9sA6QVhSux25n6ni
Bf/Jlm2gNpTvtOhcxbxEJG3dY3AoWRjRDfugzKN2kBnFLiM/LmPSbUoqrxnhl9bM4uLxbEbR18Pi
zta5BPRMUDP4wV3e1kKAyh5c42rw433e1jeCIhtLHPNHIZU6DWuVAt8kDpqzcsDqk7Y6rxWyr31+
mXEwSWW6gL4EsNubj6YT7ez9+96+6ymUjEI4Z707RJrP2u0dgOGV6pHR4r5KqfzWgPPlHI6IIWYm
Mgk4tNIQ/dXOwm8KhIqdwwy7YP3j2PrKGoKLOunPv8LD2vvk0WneYB1rlKSL1tXjxgksqyqZOlir
anNpE+esqh8dhgkINdYD4yyvaiSR/ib+6OFT0YKa7KBo+Evdq4x/gG4WblHKkoYvG9t+182LcRUO
pXcYBbm+Nx3RzLpFAtsihPtTeoJaWIxO9CMYuz5BIJxZjteqNGliBNXrZQVdZoAO+8rdCVqyt9Ng
mY0KXCFBKZavpOOhmtVSLgawp9cms6o9A8B9HstGRGdnNjjlyy2gpo3ipNDtqV9/2+J3xoaMA/e8
JBhKwhOUpRrFFQaf1N41vx3vSJsNCSZhIPdytYlvOSc7nUSfIe5yx66fiCMb6coy8sq9xfYUqglK
w7e3Q8AdA9fKztAa+jMmd2YGQCqiyZbgsAbZf1a0Enl8zqAfjbrheKBPLWC4gD2/YG56tvsoMOX2
G8xgAY9hCbs2dAKFVabxDlqgbfqz2BHfqRPzN1nM8fJBbtvPMMrpHg6nS+BK+QhqGSomupmD0Gzv
TwSuZjTytmNQvqGbfi1CWXHBBS9cC3DxcbW5RmUFyXq//h22R1+8QRboFhoCuaEaoXO65ee8NwNS
kGlvnakBRx1hikibyJNGTnNUtw7mwZO4yfFf5JI3O5JMud5eUAJZ6pm4Y025rG1DWQqEsQ95MnGj
P0+plGqxlNbnB4eHh4c1FjeLrZtCAPd/LX+vIq9FX0oWpRD5NbUDyeefF8yWCelRGq+wTxCpa28B
AGc/5s4/eaI4e4fmY2hHKcGmIKyV8hsKFxHtdhYdJXqgsmteS5igGTMR78ENclqgvzUCGdFoSRF4
Gyo3XIw1uhHQs7TJdzLEUVX2VKw0wbAMtNJbNNQDGXj29o8THGmvUYb4NhvpE4DUvIfDWgVbr3xZ
r2xqVOF+60SIu9jKi/xOSHoZr4FxCQvIrMcr0FjrefYG9dV+DqODEADSDKo786zdNlPIiZ4kafZf
9l6pvp154xy4TTG1vl0rcHSRttHE6fZ1aQlhnXVtoRlrhd62JtUZMmOlARuoHwOGOfPENfLgIPvU
eDAloK9ZqYIv4tl9jpinwdglJlI1LpcN8LHWNdaQj1M2oGmPIxzvBln1aPYWgML7qRE1DcOy/jk8
Ymk8MyEQdv6a4Af/Gv6K4KYs6Gy/IhBknK/VmKj5EmrU0zfGb/WWtRSQUkfgR62C5WpoZijAqqWb
RbxIHrFZFY+aGqqaPim18u4Zdsn561v0gY38lwynf5GnVZWJCJsmmygJLk3tKi+3phLuvOgO8O8e
zhsw4bC5noCodqhtnBPAMgf9/q8okoOZg81FrBcLnaJgn6sLITQOYKWqHgpyD85gJSlIxZUePexd
DirHKcb2theLEthsPoXjJ3afXVSRhSxA232SpSAL3QJifUKJquFjbvbJDWGO4Wet2cXTrrQkVKjM
2HK4+JMNMNjQ5uuwMkOUBFTN4thYR3HBYu9bHUjNzoioFquWCKbHUrUvymyMuZkhRWIrHPNjsJC0
ppshxjMcCJ0nYj4qbS/qo1KiOaGyMyGzQlYPMYeDJ/AOEeZJ3EBSANNsVVLjHjFrhKOP48Cmpo/O
szq89uLLgux/2lvdY1PoeW3a9XMbPal6wqXEikwy4SNyBZJErRmAqNrsgo7uPRIP2L1guLyc2Vf/
lG4U4H5MVVnbfXMwFlgWNxUgEDoyPx8MMioVRYq+DP6XgnsAy8vnJaht5KGTOPB4rOc2DrSEWjmY
6++E29BGA8fAGkUs4aW5EU8b5NY/IqcOZrYOxgvlx+TdgvgfhKyfeURzcHRtVbKaK22UG0LvYAYa
Z6VetmD6U9mCUvyeADUkX87ClrZBeSEBkc4MP60GFJb/rQewLHyO2UUt4ed1+veeIuvrD0/aR4bT
WCkFbwCqHpBjPjbPRXnP+gt4rzsv30iRWDTppRl7IlI4UZUXG9h+bugRxTpFKVYJUOQL+7aASKsT
UN2Qv3zbEDtzXXQeVNaaAoJEg/0uCrU1zQRQCWa7A0JafLCTyLyezZD9K0ZR5krpWWRGAR8vhlgF
T4ulffWdTgLmvKnuDrHoAvGT3ejw0YwsfFCuo2HguFgzbKLyTT9ZOyGtIBm7P0iFoV5RskSs3zeU
5PvpVhjyo1Xj9XGPeTKuZ4+duK9kp/KGO47u1rVdZ/u8bIUCxTkC9izP0ekYgYeHzjKrGxMUKxuP
Dt1bTpNAq0MaCjp1BOGGLVepnVsek1vhEXjnaluiIEoQFv+JB1w2J+3OOC5/BEhFHNmauJVB2a+m
iXRHyue1EGxVllyr9rsxc8FIa0nAYO+2yksM4yJd5/OtO/7efYkODGArS0eD0VRHGOwk7E13LYws
Gu4brbkkUqAyisPXZO3ldMDlGPrl9XrrCuAfRq9n6sciG67v++FejZqlAg4fwcBT1QtJSnECYoKZ
9dbd4xj6tR8YFR6YX74hr3KK4Mvaka3UKUQ4OW9RrPcm1RZY1l7nlKdeqFkR3zEbg0UeKTNsxDQ0
7ozMYQ8ppNoL0z/xQlOfES5NMSy2QiYiTPwa7zDh1d/tSnocwhUHjoaXjmPc+6FFA0NpERuMTBwf
i0yp2IxBLhox0MztE9jbxJ7ouOtqWhtWCY+C6Bzw4XACj4zFR2AFOawCS5mMTD84ip/wH0FosOg9
26PEIEpvJCWf/dOalxUtEig2bNxz20lcKPoNeIDfzpjf4hnLKnkaMv7Seerl4uFc3CpBqyAamL1+
54PO8z8nJM7UKmZ2IdVUtHdbjoutSRhXBoxOXl0yh/6LkGLEWbxQh3fGR+qAoq7TcBmWDIYrr79T
etuxS2Rdw7K+2N4ltuumgFxjd9VCbceEhDdHu9u/aPZsEnByZTzHdWKjxJhN2G2wHtggZ+uEcSpS
l4N8INUwH55394YSsGWsTG533FUjfM5HgmByFEb5JK2G2t8VrQ78LWFl0FG/JwEuA38rVB7aW6Sq
cys5qCAbQfOgmKbCjj1kA72Mes6qNowitMrD+FBSkPl6M+etWQ7y5D2zcaG7ZwAJloXhSKzJh8bO
w8JQpljqF/X+FVfcg+B/70SynRoX1PRduIE5PxNiwzwuooDDSiwvXvEiSUk/r45pL+2Diio7S7e6
nmSu/unrLD+YFHPji2PKUNJktIvrDFLeFO17IEuOu+LIJwQOF+iqBDbGxtvUvC1vvjouXo/w1GLa
fchIVpJfQ6dhqZW2P6l0rNt0FoxDkrQdtAZC+NWlbHPFwgMx1LpDdpVxivE/XEPMeoIB/mlgLsL3
cyYPEi9nEOYp9Ippx5gh/5VUmqqTfB48ptMO1+S/z7aoV/lYz854MOnNewCGlvHYYWiCUmRw63yH
CK5N3hvc891Y+sEIklgGv5zUB30rlIrSPcqVs3K4HaS4Xqa5LI1LElYw4LHM1l/bkjrjvLq8aBTI
NTgDD/PBlGlcq1OALQP91UlcelLmgIZKMC/XGe/Az9zUydLY18gAJgbV6V1HeZGFb9VDmFVO0k0z
1/68YVD9P9F5TnyPOi9HzgCAncPItNj/m3+ORZOn6UXT8GIrIZR8z+11k3E7hJWexz8fRmBydGtV
4BjiQgAFXH6HaASM5e3fJL2eE2mGp97DrUemDuEFfJJatseRJE7H8Ia4uJSsqSdheYESbI+HIsLl
V/zxyKPYvW0EqvmqNxT/pi3NjezQHUTdNunKonMrJJ9FUXrcZIdVwwtGBQDXgHTTjlQgG4kgF7qG
8NuX6vdFJSgGPeqrnOfbPKhVxiZ4KHBMi4JrQi3JEHU1HuEI4fluzRZ5hSHXMOAYAuit+frVQhCF
dy4CjsvN116MW5zjte3qU/JZ5xVBonYObOiedDEP9M7ufdfbcA9bC71pgeJV3luED8VvnSnDtxYP
xnSkbm623LFhWL3GOWfezzuUcHel5sZNBezZQ2VtS9O51WhxEcUUsF0yyKhoozaDdqP/s40816oi
3h6fOW6Jnh8SIVNHMLOdLJZ2XB1Ws7YhRYNVzRkonHBEmKv3Ro5xD0llqW8bTK95ryBTwsFssAj9
wYjShRk0S1LKxnkn+XWOe3Akz+5qj3yw705006JZQ9tAqP23zoU8cIdVVHUM7eSoTa1yeqdR2T4N
pgKsbRGvjEoozFSxsMfowbN3TOam+ZhHuGSsx71MFWOxsOnDuPoKwbKUwqUwiUYjtstcK8YIa+8V
EAf2KT1LpmeZZ48PBV9bZxHUHoIw51jnLAps/BbL2ND9EHPEvUThgIwyFCg9yOqF6+cZ3wNXsd0Y
CH1u+qZLa+GFRbM1cyS+G2xGlN+hA0G52AcE1hT0jO0rGOs5B3c/+Hf9ebFBZAeWy23DAQeaTSgq
Z+YTWLByad4jKA0o3xKAVPAD+js/7rQxNRLMyIXH+thBIik+pp8qj2OfhmSZZycVf//a75jWD3qn
qM9PBpauUrXYwDbDcC31dKublPsm/QAPpqR9A1gCMNSDzf3tjcbgm8VBTFvjSqpeEX8r9MMhVB9d
AO87QrI+6dV/jF5F463skzgJst9dVBAQ5R2XVrCGkEDxj1hY6m44xAQnv6m8HIQvN0Ab/flq6Pvc
b7h65pA5Lc8fYNFVI5TQfDdtNrOi+k2WQJmcMJcOL95G7qrJdO5cvQ46h3Fbnf1WcANcZTCydKaU
rWSiHNrXQu2fCBeqtUHrgZHcDAppnbVstmxCCUlVNePJ7+PMkE/oK//NPKnglPtUPv98cIMN2BqI
dmimEQgWLKohg0GxCd+n7Qh+rTuSVhSsJUHoqo3VdlsxlPNqAStzLq9cRh13QBkUzZ8LWL6qIPtX
V/XSEY7qi1QHXO6yHLTCpuNvU2R4ssQYmnumHqKoTee+JChSK5cdqlJmSsw9CUkc+gxwzed9pd0N
Wu/aJDE6N9KZXrCsmjRnzLt91Dtbg0xqSSJg6VFhYGVXnP/wcUjNH3AlXM3JtJDhqjB+L0PgixP+
ILRTTFuZ2yqVnbX96KL3p4EJ62MP5MeEAWbT9cVUT7r/C9WUeHT35sOT+JfvDqn5E4K7/Hf52nL0
AjOsv6GlO7Bc+CySQe76jtvy3A2giLAxRr65476vuR68af+hBDspMADi2DeLcQ7Inmbn25/0j3sV
Cb2KAd0bUghaSV+Tdp8Gm+64cMgxHeike2wmZH2CRZx8EN50Lw+IGUcicWFStMDsAzZxILJvu06V
me/WqtVewTyh2aMKaThAmmVEAWS/0rbS/6XAzanPPuB8fGahoi+6RVSrkxqzSqC2IGZtSmmxGsiR
h9qo9lfPQ7De4Sx+mk4jDGW8lPuGisi2cceEoMeQ8d+MuZ4dg/e9IMfy34UxWDDTmJjYnIxPOeS9
HX6FrmIxijMzwuYtHvZFv3d32a/OF22swbbyIvavrxZlRq9/KsS8M9lxGHYQ56A3zNHsNW2N8LKL
BKfDG3M0r6sZ9CCrHWqPuHFV2kapT1B0a2RSJgGByIcK3MXFKhzHMmosyy6offP0AdP2pK5nqiFW
pnv76V6xSVu4qEhd0zP+iwxDTPEBe8v+7NBgy+679K5t/y//0niHB8mapV+bT93uDrO8RdinO9iM
3EncrAMPgxGwdsgvNJSKUWwuXgpbd1L37GjEEK8weptP342dr39nx+gRLLbKxLNj3RzfA6exm+r1
XNkY9/TBc/w7fggkvQQ9aLwWqItOkqbk86ZY1XfQ5OXLVnahJ9GyxJdJ8WGslZY9IfDK7V47hhg2
Ax21VjZvwu+bFRZ9RWKhxzvXjkLt1LSb02cA9qiYWGhhq0AscColaz/OzHfz/qRCqxkzG9X2BwLj
U3QIhCSvKfGZBl1EbGmsnL9unmABTthdKCd1oTj1ncmHbA/nkI9U6bkdPyaxHHaTMHoyTBZ6Th6D
8WSCWF8rTqzQJMxF5bGMdTnd0rEvbj4/sFLsWiq/4Svadl9oOaAf4TVMpqta/zQMewmpjxy4LO1x
Wdq8UNr7/dbCgmPA6Xxc7b1+m+It75acCZ9ou4xJbfonRT6csSrghYsPTtGX5MBUShgir/E731R5
xBSF56GMawb6wE5HfZzIsJZDVLUHusEZlynQTy7tf5aomaMpvLC2n0O4OStJ7qlP1ptDLWfTiaWK
3TOit9PZlFMDK4LhBI2+qbGcBSqfVKUAMirATSrGwCv6ZehwQV78L5YMwaVCspKEJC0RGVoYcjo8
/xXR94AH7rHDRfKNEDn0en87wbxmcTQZmKqxrn4CCDz1x8eSJg3W61NGdgQx+mcDPTeIIv7maVFC
IEYzPyxpjWlx80YGScELos66kOrJvWShQTdocrfxc5cJH9otb+npghszdMdYykfJpscK6F+zfigm
3Hl5YxRundRctaH7vzbgaaaRXtnGLlt2kkqHIIJ25nNLVVbOoXVLT+EzS1c6CQWJlBHzA5ULp+Il
fLSJbIiABVbrC0IwreAjIl3MfpFBe+4L3I/6X7Kl0sLON0q6V7zvKHodmlrMb4vQx+s01GcDoOkm
SGURLJ33fbd03JtHhTxbStW+l5TPoJoniSDeWg1XQmT0AWqG/5GaS4A2wrIm+p0GwRPXIz+0ZKvv
I6WLWHSnQB6UtV2uoHJe5a8jH1lW+XGZ/HBPuCJF1CBeqnqvnAQBBROZ3kpKRObIbnZDmw5YicyS
GCok2PteWcDcTkPYSWdACskJyviT9S1e+JEpvWgI/mg8ZxBGdPUzOZYiqSsikwLFg0FuJzcUumii
H5WfEjTH4fb89PRlS4cedLypqGa3QNqxujngRVV2JSC2d1By0GWpBCbl5BM3bwje/jYaONQrJCJl
WxRz1tajCLS8u17R84CFhoCtj3FLGhkxK/6IJJr9gavMfD/163HxpIMPj66Oru5Zs0aBBndHQMre
5SXUT73Np+MbLaw4Cq7d5CkJzHobSxucd0xFg3e5Sio4xBM8H+HYe9iWFQwyrYhT/0DFaU5+imp5
Qq6jXp/YiCGXU3D3MxuOgMBeVXmsx4veKJnVvGNj2dITjK5l0J6onY8nskpVMe9PxMY1A4EhV6f7
FfCScukX8Xx+4B/kdBYJHVk7Iu4/fu4tspegsYJ+D+cmZ4N6G9AyTyQvOoLxdzQ4yZ2bvgxxVQG9
fbCIMQkNu/+v3yPJyLjSMp+DOYBfL7iLiSQ9dBeZ0ynFmSy67wzQIHxKJh9roW+W7rQ4IrJleubt
aF8trlKtJj6yhEB0+b1xZ56VD9HgyCGpHxVBdkYOfH7vU87YJYzWEBo3jWMvJ/kA0V62zZkOLj77
YyDz+HfMGNnOe0caB7OLdPwtU4DDoguPCfR4O94gmtwG5G8qNJhTuZiB6HKPVbvxND/KAIWIDOuI
CBYeCcU1hAke/tVzqpxkzNqc6yhohJfO1LEYmV35R1ONjXTXpyYLvmfHvKpIVullTxmSbn+FpiLa
ksz0gxT4NnFf5iBC9hW1Jfs3Mv65beh0pPxUaPLh7nWIDZWBmz+jY3lzO3Q7dNlrREBid0IFjskq
wvmTMMFK9XD4zvh2WHWnCwv/b5GIswuQcbfaW6OCHa6+j9/c6FLLVUC/xM1XN/okjZzv6OeRE8jn
/XFBJ8cvzaif62JEESELKL5W7jeaTOqKJXqKEXblCXPTM7Qx9AvEHErcDq9XAsGZT3FXbAA7bNOQ
xYZQ3etT9uJKPvboo45vDU4wxbzOmccTv3nUTUdi+/bf/5yZaTOHqeQTmbA9wveUrN4CUGsctms5
nLmqDftZiR6Fq7YzsPf/u0VoJ7FDFf7moIb6vurs4jftO1Qrxbx9EIopzeKNCMZzfRT4mh38RGlj
HWBg4zsKSz/dryuXkOO9LJv4qelwGdW7ZsLTLskhIdtITjkIFj0OJw7Q2kItU3o8fZssMAS7Gnhf
1Zd3dJiFDUl6nFbvnzBMB1Wu7dZv1qnOVIU9L/ZQuCWIFLSEg37kO9IorCTJldAPF13lcLMI3FSd
NbL7Vtr4mJtMmFKUUM6TgX+zU3RZ80II8FmaXZmGg4/4Re651LYkFGGUg6NL49L5+LpqKfy9jjrh
D1WrOQj00a1sbURdNh2+nnNKfr2IeLMOQodfh26XnRDrnvAiC5cr4AwQszywSLv8iwr0JnepXHH9
q8d2wa4CJW+xAWyiLCC2grgnylfOJ7Inwr87GIXyH5ORBklRJAJFArvCOR4TNcQ9QO6Gk7tUhSdu
ggaxLhrafZYHgBqNr8uC8TsJJ3A0uIsTfPWdP2fI4JfcbSRfd1WMT6zZTW+UjzEWbf8GmD/Sk0iF
JzXw3+Q6lGj93xoNXBKtCztW4idQnwqj9UVUqX6OWGjcmY/KobF21fI7YBEyx7qOG3jCMJRseluz
BDySgCdeeHHU6oQP0ezyNrcZ3UXcrdAvINmjb5p8ili5QlrT9sdW38GIVSlKehmOFso4Pl9iaz6z
crt1FdoeXaiArVt5MqtGUHZy2txQF7v11xF5UCrOHqJzJdzNbO0wg83Dqz6kgAPuh7cSW4sC0tvH
dHGNRWH+010rABYhpLt5zuKxTKoBOfe+L63j9iBL5QCxJM1nooLWQQVuhoqDkFp73Oh05Qt8F4yx
dD9mY4czmje+xiDRO4S8nQPoicosifaNi3EHWvcKFzyvO4pe3R8X8qS+uhtyFbn/Jc2iJ0OBqKA/
8+IvzyX3ViQpTLPLaLmQjr1EXIPOVZ+kANIenc4fNpX2JISciiCSXpUevPU22Tt8xVFZv1RRqt0R
hMqqUv2Om/iZHX5z5vbVLF+AJ6OpU5YBFXSgVVKlcm7/lqWej1+F0yAiz+eSsIoZRI7g3SYw5Rgi
PqTd/GNkP9sk/ER3ZDcLo7WcRftPZRc5HcFjqEJuaEmilBsleqdCyJUVbDhvymwqXMyPssOk3rGV
AZYZ7kef2hgr3UhNjJwodwtAiJUf2s52wOxtCXml9/tyUo37s8joCZc+doVDyO9saFwyhdivbQHn
ktnQhHnRVHFZlY4ih2YCFDq7g4Yw9cdwE2Rt8D41dhNKaN3SOj0mAKgtflQDR0Yquj81WuNnGpZC
ykseqzGAfXolMzfM5HE6t0yvM40roKND4fFVbc8x5eM2SEwfTjvewNhyfkkp3BoXwqxYWAyiYkjs
ftF+bFVTofugYn+opwXMUVFG5rqI99YtTWnsMeN0/1t9bJWI81i9MEAcCFegyEzSvywkFKGvqGq8
PEuhf0/DkrOKSOFVkI2ZTFSx3Qm9JZ7gYxLAPjABp76t1yNd3gJ7jkuh+SgVo7eNo+k0CindCAT4
7yveim2UmPXdF9SQnz2os01ygwOAuSu+gFjh59FSSQmAEQ3ojYec8KPS69C8VfNzytziZb10D6sD
9kgaSAawZKeC3GHdCjrZL6Nso1XunUL9NZjcDdib56NAJwCeq2Vv/RYclgZanMUi762twsOfdq5t
C9pIjsV+imDXLDwoh21dfXgw18S0qzKgUWiHKPTiUFnJ3NRlupUS/16ui8sHBWvdJVr5yHMfjYoL
SOZ6EO/BIacnYq/2t1vlKoe1gCU9STnFINEgqMqCEHWTpdkiDGaG3XVDmMQJYh93IpOP6JE+ZSjz
ON571+7jb9aikCYWbxBiXwXhSEaEWSFDXR72T2m/eWGLJ3vGViXaDVhZYqU8EidH6pI2lJFulMqz
JRBsqEeWjqh7kLIG86/c/zWoeUj1ka0v2G1vG7fTEXi7aUYoionww1UqWLEIttAhRtTRlEq6BG6c
BpzNJhMyhwh4PrhzkPQ0uN7uFfE64lCl57+oS9X4/yGFZsfFL8ezVx/4VjsgN9PGnZC4Z2pHrkfK
M03cd/W8ixPQxLnIpCKdS6jPjIfzZPXqmQPyp4Gbj2VyRte2e8lBb0vxKMKIcG642pVkcBUXiCBa
QFVzaMGORb8VQTUIzHqe+WLvfa6eUO2ltzim1EGdixOayrfGsbr/eRdYtXcTzBA4N4EIz7cslFPq
wpabgPxo9RdYN/P6bAA78T/6uld8NjumftHe1PejTsjlZkyxVypTIcC6LltvVkNo69adD9FgLmr3
uCrUtnoCvVlFzee04L/jokKGmMo6G6r0wyVmHvh/mCA4DwiUVF8d5ZttScnR14aVw1nUlPxr7hLs
nweoP3D2KARSetccl05MJ78/Df5HBUR4qeG9E5ZCQVJfW2OoXp5dwN62faaWBhmu8kAnZ9xFOgOp
pGo614rQPKDnc6QQ/bfRdyq3iPJ8kue5loKK+Tk88cjl5XPDR2QyJ4l7qlkO9KTPZIdCyw7G/7zP
rt8FK6oytIkR3zy5NpkEG0tS0b4AkCQy+mwMqFO9B6DX0v70CVvyfNKNjcWOROx4vlXHeoG84xFK
1DMsDeNHadV4+1RObELGUrYM5FX/xwHbFuHlzjPCXUFCAPruwrPuvF/mTM282ELYMzEsI/hx87AV
7WAuC7M2KIkaThwaWoTrrV6Bw+viTO0LGrLTy4X5WXO6PE21c2MrxLeOGIWHY5XoW4VqWRLMjCC8
POzMyqc/oHOtePyZ60XF6QN7whB6L7WNR4RDmgCSgeyp9ggdvsnLzDIQlw9hwFz3a8lu3Xqc0G18
cpTUOmpD0oeRLoK8gGj43zCBkGT8bU+M4gLjhEKkz1xxfRHUYACApsmjrHpTIwOReHsbsHWbtppb
s6gbYDLPvjqSfkpQZLtyPlJ1OAl3T56gWnSboAZjDngI3NHQv6RgDQA3vr/KMG4KYSKOqL01aEFQ
Yb8Uq4QiOGD0uKyptCujqJxVjxFaRbw18Bk18Bw1qshxurT7Fw5Og6KNYqpDjn5Tp/d9TeXRClMJ
g7ldFBWpfKdOD1ceQh0w17eifSH/BgSzHaEw978uTXbkogiwBsLAc5PjURo2f+1lk3SZWIIG+GTJ
Ovs1T1Xml+7Yi/mdpuN57F/m12MTIQ/NScnfXzalS9mSxUbIVcJNhgcjNYYK4XzRvE4EUrEE7Gzc
zxBHFZhMYMJ31HqNJjtqxEhegxbLPaDi4JpYy2Tz2OJEoZeYuvhRNLSBBlfdJg/wYOnrUVkvYQKj
sbAWF365O06fsQypOgEL8pSzCmidhmyzi+APcB77j/usg9mOisFMROAdAquukWEw8W3GKwQOPiW2
8SNMHDNSXh+GYgpaNXgD5d0UWOYncBXtyC4+QOnvoB+XfteDToJwKwGHSRzNNdSMkV1/mbY2+uyI
pTRkbvyjHmR2A4/jQJ4DkjNUWiyeZhYV5jzyr4SSPMSz7Sj9OPON5GGLMSyaj1VsIdpCz4fNGozS
zaq4eWgbK2gpvUM+/tdylrWVf9t1wzIzAAILeMrVIcdASpuXlH5CblEh8wYnPltC0MbPD+BmOXKk
B+awlDhW4+Ep6zWP7MBf+h7cX7D6Tsn0A+RCChf7X7+6vHZ5jfA+NKUjUDoFWdoNoC37Keetv+VT
i8XruluGhPNZkOJKoGmRT/XLR2NMsKdVcyMhn8qN4XzDUtepyxk5fqhUo7TSqVhPUJLCCuNvtFCZ
kyyqzEaHkwxOnJCeWFma625HAnEMYk6q3bnas7p10f6+Xk5iIElEhDcglsaA9dXS6QPJGYYHFyM4
aY0VnfYT5GwUW7C9e+WDWHo1saD8qk4DulMJ94wOrfF6WAuPGF+RqZhNsZCngw9zyRnxjj2RNGxj
FVPdtdjhQ5SWou4609sX5LCByEw5/uKWRVN0YavltpVH7v3RidvlzXTVT+Gp2QhrPvX0LfvMzWV7
0rashscNKP9dizSkCN7bE6h4xU4MZXeHoPdpAXMixPy7wKxUeVlRpca4h0CaGPItYQbq1c2TBWPh
XdCh+dDNJEmI0FMsZkAcMeVmRH+8Mwdltr7g44N2wH0y0ASULGueEk2vosvLObe0ctal3bXl8pjo
AIMAGC9Iy1RwllqFr/jo0tfOiVTQpcXNNzxyTKfqQqfwqD0DFb3hvuWYApilq9Ivhl9QI9+ufZoR
DU9l8Vcp+W8+TKlrjgOPnP3B+W8u1fr56HuXPViOQiwIf4f1fMIotn6rqJh/+/IyRAp1xRJqrAKk
SfRTlvWjQruJxds0jCgD1b8uSRIF0Oa8x3m2rgslH7wifmhZdEpwmCgAeG/cRNWSjIsrem1K+NJe
aeH52k7PnZm/Ro7NkzysKTc9IV+txbKINr6LvgD1FDLZWLSyqxRQY4EncIMOTI3/vsJlEEBqEJJN
F2+prQhm1+CirZzqJOoljgKF2C5mrIDYQjzV4z0iiYVamLZaN4CJSnCtft86idsi/FFmFgdVApHc
/V53PvGw2sB0xie2eM7+4ZTkXyQJxiNf0hmuA/ZAmAWroseX22t4C4b9qYXr9F/+uDhBeyy8rFp0
2qwgJq804ENt3VIntNIWrlvNwEOvKVTVm1zR9plrQ71I3OIgIhAtXFZ2UN87vV2JZjwt41OXdUct
EdiTLOuoZLLUd/5hzUcAA7aCBGpm8S/3sxwQ8NaSa082NaUGlGrnIFUttjcibKuXNQSGCIirVRPc
zzFEUHqsOX4kxR8NG0COx4LyQU4Q6kAcRyolqQBYNN2ww8i4VRDlPJLk5QR1I5ODGFvBwjzsQVQB
JHgHIg5yWGmcR83l/q3QmkbKZPLtJZcQ9hocFmLKHGuetOUOAdKF2G+tRxQRtt8gvKo7YoKXypsu
3GbqUMrM+ZJAsYcrdi6TwtIIH6Wo6pCSIEtNH3GQC13UWPlMMJt4NrRpLLYJRmv6fEvJXyGbtCQR
PPYWeFOB+MQsa+i3Ab/UDqtrvxKhrYofrYHi6ngg/h2tB3j9gosDoU6hib9d/VycJGIf1x7IZY7z
W4r7PpKceg/7QO/GQihSHRrf0Z2Ed/+yYHAoI2rbIJbyUT40ciO+3xWjx3u6MUSWUaBi7QSsBdWp
CHpoVsoO03mOBQc+2wMC/12YwU9w1nqhBASvfiex1d+WzfZZzLz3nOLgYHUCbhR69/JXmI/hrkRz
wzBfYAGOXJWcjCUGNfAtSg0OY9vMY0XWaiTk4IVEvzKMZuMLbuLbyDhVrlcE6Q7cgbFMJDGvWNbw
cwXXwXSKLb6MNV6SNBPkRcNASXTC7rifLWx/NSJ/OLNHWAdf9CsZ9gwbdbkmPWENJgwFdyul+lo2
AyzJBI0IW2uYzyTl3+8jkJPMMANiuFacgASJkii5wS58buED8tEHJIKMvUFgpH+rW4dNG6tGUofo
eXIajkCL62pXENAi77NUlqy7zUNhuC6LMf7toJDIiFmsRLhWRpR2wM3U3UzPUSS806/G2MbqZs8j
VTyg2EWSS4ZTMcBn+7x42OtHZKckZXllyYqeWP+RXDmpHrpHCfyVH/wcijo9iqG9pmw2fUKCgWwU
Nww/q6P7dPPcokCfC12un+1O3BUf7Spi4B6Vmb9qwKaWKVDAPHQKRvtzZGtjJ5C36yKxgv+BV9/F
xw+kYoJGV/oQsBc3q+x7CfBw/pElPx1pwvuckUExf33rjfR105XPiYC+2cjrFkTp8DX3QWxuVifc
LJrupuM5L0CyBbEMJLnZj4hnabRhi+CQd61VqouCndn4P9Al4K5QjrfPTFSFtheoI+G6ZqIB0BIZ
oztMbb/jIfHLD+mJRXLyOCc7OEYZGIegWMm7p22nFZsHJ1pOphNd0F+ftqnYRu3WWQb+WLfR67Q9
6yqI4Iivnm5wz/4JaUX3HfE9BWISGOe3C+B9jov54NzhLsqSrkjH+qfxJorP9EA7EUeUqKKWujjS
ZpGHpqMkh9KgandBijH1xST1CI4zlqpjRb0bXpir9Fnh114T2OhdJ2WyUd1zLWn39AqPWcRLDlov
21GQBUaaulutXa9fBZkWntjX0fyHTnbp0cBG1KD4wYMdCOJ8ta9Q7oaRD7CG89XrFT5Bu1m2NcWf
ReNDVq0LbS6JAcOZkye8c7wnDEFJMPr1JfDc2u6CdGbZJ4947szXNrZXDwd6h0nofq2x3c0qM4E9
/pm7YymsFu+O2zbVe4/B6qGlvlFmw0JYanj/R3riWAZ4OZUy0QRk8/ex/FtCxIUrBQGSa2M0QHzf
R1njhJR7+laIyTKLUgLF0HFm5128mR9C+MMkb38TMfuzBMQpQlW755z3Wzr9OdMbMVn9ZS2ifV57
P9SAVRe/9/mmffH6m0VRXVHWl2P+vh2dAld2oojlt6fORRHZYnSgjZXgv+8eU5vRFNBloNjbPlN/
me1MfaigKfirQZJjrsQk3/q8HuetnIGuxg5m9Tp3u0a8tqU5vdNWnln62jmcy/sRzBFQ04TrpX/O
BYQJ5PpC/W0qIxgRRyQgg+QrtEKf/jsMrzYxbQhS55Q9w4neSsYicPGT6dYB7UbcnJzPrn8Mdn/s
9vKdE+x74M6ugob+K3F1xIEjzi4F5R0kCtUuJ7bhmktc/bUuG+eoQy4RtN//XWYRO1OvLKlTsCua
lcERvH5CFZ3RGRzESm1V5HaydcCyjBenq8Boih4OGUHU54leY/0TzRUBvZtrweNRr3CGo6aya//3
9RQVmw4S6LEHPKu8UFol+/o1vGBRuL5UrohNITPYGXVPrjw/na+eDttrV5lOdPS4tX+2WZ4Ej5tE
bnnWHoiwsXJyf4VMYQTsjisGqhJeGaDuNNBCEPZexf5+Fu6rRhHC0cFCTOLxhcyqA+2NygYUES5D
O7p1Q/Vc/QLsZSyFOhCHDE9SrgYFA4PIQxO9Ix8rE3mO42EIKbYTJid7/L+6L6ROocH+eY4hyKN/
fmM4p2vaw9DvcgWVVfU5tZ2i9ztlqZIefo2pN+mFahvg3XNVAOrBYm58Idw6ESuTD64inMrNsJVI
eA3KG0STnF8ZtteUrWYbBKotslFsvQOCM9zY2kRH1qT6C2j3aMT7PFpobEh6GjfSPsIyZEcX3VoB
m6ug6lFuhChSRCMzku32jO9hmAm+Hp4z4M2iAwZ7w+H65PWfn4LLxt6uyDpvfMa7juzu/TlV62Jt
VJUP0Evval9MGcjFf0PyS1KcWG2imXgIkaZgDPFs2VLHQJSlrCzXQ15ePeXHhw8Ivsi+7AY1UHrU
vuWtlPjbG//Vmee2zdKS9hZ3Vvz8QrP2VgkxmZ7rauhb3tQiEEEGzBNoPnRo6P5uhtlfUFnTqjoh
bYhmo/8ySHJLVDimc5OobJsuj0mkKuyO3tboKCwvfVPneDlJpsy9gFsrftX2S8HuE8GRgRb3carz
9QK6/hIZk+0BX1FdWKXQZqVghAL86QTVIdBCiXL5XtMDjJoWZEtyu6p2voqkmKeupWg1+jfHVvnK
JxP/aSHRv/9QIT1uCjqRUGLu/HizKdR6u+vEQHZVgemBuiSGLFuAJ90jUYy4R1ND/HqBNUheR+f4
wJs5rOonQMEJgfztMENCP6jWCV3WTzsHLdTt+vuens67qagbLk6aY2WLJ0nIAHJecCOA1uueEwWD
Ta3zF+eyDQEYb8KFZXWa9UKAbiqKngLqAA0cN8PaQh4PFVrqzeQN8nvsqc5aMjoFP2Imp/E0Givl
lCnJiV3H99cccIJbulR1sDathqdzG3No0i0w4xDBaIfXJp7izDwghzFZ6ilpRApsQKsn3ifvLZIh
NCiJUkqtko/iwESDTYC6LYoZdQh0G4z0DxYjzj2rhhWmp0yCS/iu7he2uJATUdHw/jN0MwuCmyLk
qrdtQR+M1HVWWItCxAXDReVOZJSDZlzKrnGtEN+f3yVjgY9rygQyOzSBGSLjSiAQmIZHRsYWpAUa
OaUfhPC6oz2qR8DIWRQ9D7jgvuDhbK9ByCGPGK8Jrqb2k9rChsUe+qsX7xFLr2lxNbNhpeB6SQO+
VIsthi0vtpJU6KSWxcHs14eOzwSst6GnB8MESygzTJh2MtdalkU6uOmswM5GhAIys3W7vAxGZejT
ipy+M6iVZw8xMmtkOnD4Dm7yNnZQLk1iT1hLE3F73G0oyDrrZVYNyp8Cg+iwI9anoN1ZOsBMci7L
O4CcjiP7VzuaDMqljJywKhmasTAi0NCbQ/h9r2SdGN5/dZBolQxvuzkNrEjAbvO/8MYpZ1aV3h8D
7SvSulbrMiDGa3jzNBgNWZh/VxW3NdRsx/M5rQp7LClLInGdnN1vsgGfEUms6JZ136o7zF5GKaZb
fp1pkfLzKajkz8T3PJ3ntqOmu1Z0c+D88f4qA17nZCsnCs4BWUf0aUyFLEuzW42qROlJmMFkRzVr
5ge8RZOLm/Isso/0ik5aiLuPP7wb98AnEuWPsLnxXq+vfVtgYpBVYPPvq3RFuvsQq3k8li+qUu8j
0Lkfb+qQEbtcHq3QFhqiMCqqJGmGm1oDcCZS5ENDbQAPCzh2qaTGGMdcRugbv3+g8XT/bNoVkdyO
LCIrt6LbRCPvz+f8teqR2n9whFDC5BvmypRQFlk8yNW0x0a/tvCpTdMtKdFV1o5RTvh7tW780uPR
qJeJkdZI9S3deeL0WJxHzyrlXY8llHar8+sXpfUX3lJfZoGdUpVHnOAq6y/0Dy6exAB3qCHUiURU
tywFZPR2LAemqNoPz9EFi0ZE/GZkjoJjp0XhAK4DYxyN0xcwmQv/rjWJvUkwDPgI3puq2LN3tALd
Z6UqiINoJFn+TBya2qltnkmJlKYPe3m2ZPXps+ELQzAJ8l7GNGT0v5IRnEFM9jXeTtNOQzNEjx+T
zIuibp2autghLfuAjWhbOYjKxv5E1b9aqD9t6UEeHPNGpK/lmltO6DCr2Rk/Q8EXHoabytT5M9fH
pZ8uQyQVwEFvrk+LjGby0FjQV0flrLdsoOw0OZOTVo1v2Zujdd2c3CTDrhdA0BdGf5o0jTvk4zWG
c9e+VBkyFwbplfxzu1TZJr8jMn+K0k0tTdBYo6eUvhHmND4m/Be2apuwYCCzHBnUizpcrOR09QNu
vwMao/BBzRM52FI/bqqWcBxfx60YT3opDavdb8OsLZemH5uGyzlVq4aWyV3yBpZkHOS40ShGufmC
xIAs+tQpEJVWMkoTYuOUKKS6/NcPYa9XMq2aH6GvNe6VfxdrTSBHJsk2aJFHZB4NpnZ9pK4/b/BT
Zxc7hrzZBdsmCTjg6TpWqonJKfG1lpTI+rUoMpEK3/GZYMdBJwXF6sRlfl1g99R7jaSC81DuUsgm
L1T7MyFBxgrvXC0gZvvQizTiFvHc3peLortOPc0pWDs/Dv5yVMZjTsXAusDnFdZ0d2iiDKSW2fnk
wnjW/fJBP7kmQa/Qabik+62SWIbS7FIobREzDFNZvQuEI3fGv/NJpLiuJ21WMDy10H3OouiuKNS0
Cdy1fE97LZJ2IK/piADSJB4IO1rAnWmisjTQ24CKen6xkdSPGcUk0HfQHDTQuuUxgZYZkT/bttma
eVs25srmTZnMcizn42OxrFMlU3jrtgWt8RoImn8JO2FicpKGX9n3kAgyclM8OC3eKKjRzEfx0ATD
D6CTYjAP0LDU9yti93vYGK/5JaC7roxOaWf1oWu7t7d1cZmvgbYTUJ12EzTvJB4azmoJuVWNdKGO
CaGLkQUNGVjPrudZEBCGAUQ8uOGZ2NwDat8erOHnuMYPmrfNJAY7a3Kz6DbargrERodsiVE6zWjy
blXGf1GfEX7OmrvdGtFzoBcBZatLoy8S/OM+nv2NR7Hwf3cL4z8Cy3mi3V9UttU2EVZksBcpMfT/
bfzk4bLPXYMWG101a+tVW/RwjDKt5n8PTt4wJsbThJvSsGYkAaV8dphOmQKE3AEEhAD6jbga0rGu
pcrsPflrkAfuFd49xYl+SQKsvLexfsjBIsgBzaqM68ht3S1yqnvcmEPY7kdtd+4ABO/q+wUh4pMO
LFRwWwKatKTxNdb8wgrCavKG8mUyBFFoTdqsJQqxjVdcePx6oJJlEjnT1eEHGiJQBj5p6wxPgcHT
tdWyoPTqF6ls1p7MJuyVoRsEZV7Hm7DydEZRVicLzW2zlMxHuIox/s9GKFJnVByUODwbAFmlmLL7
ZuUE8uw/EVjaU+d+9IF02i694K7Q/LH4340qHY+mzGfvLlUzdektPr8ev+pPT8y1rCJ/CD46UY2W
7iHPlmL0oFZd1C8mimjISk/3ZbOhK5/fJq8pWor3IWByhdMon7fNO2creAe7Jwf/zVp9eNdSrPeG
0zfNjT2c7R2g4pDaoSYjhegNui6SPFIoBd85SD9cR6bzO15zShY5LY7X8dK6AHxPUxVBwlVlod2D
Jtb5TZiWYquknIJQ2h1YQHm74QU9mLU4bYP/yNRoN1QVDgwaNkonrZNsDE2HDWM6uQD/PQY+/rOV
Z1/4WdW0Tb6TTwCcmrz+qnD/MIt7j4Gj/vNnQc+fKD/MSkRp9iqc8NIkZD7DTdZxM8n4Yg4pVBKV
glGGk7JMxNdf70XkCWcoVBRfb3vzgR1AK8uJCCzlDMKu9LQQ0fiPYqvQV6Q+T7x/tjO1gXhuYBOJ
5xHb8XmU/hXv1dyYeDsOCHwnHmdDnPoXGm5t4wKc1O3XpmozHow056JrLB6K164+YnqKlKKU9HGa
Qzsun3o+HmGjAEbpncl6DtowsGT91958CLTcgGLqmpvTotPafLDI68TaShqJ7/CvfkheUR111Brm
Dzsji53Qckv6HxO3YrywdGEPrbFmoigZq4iraMPRWvpF2/C+frPtMeeNaoQ1Nb5HOW+esH7hnO/P
/n3SGDOdyV5IxxI0bS+Qo5Km7yfcZgD9PalRRs9uoOQwxqYei/TNKOIDfNTmMRrbvWk9yP63/Pw1
cEfkrbAR+Ac0wzelO3BOw5JAQ3EQ+sg0uI9WW0M87mOMQTZQ7KpWbolA9VMG5VP1Ws8CgmHNU8bE
GdBXs51MAHuRimLJHKJ5pvXZuKTys0zU4F83g3AF1vRaUuIRF9WdFJr62OFkkq+1mfjya8WtWbV+
lGTZPT23bzU638qTk2PzY7F/Cgx+X7ZFMISlSA+gDgo2RreS96zPYzgbM1fbMYVQE7euo4vhpms4
mdjTi2ZY157V9sW5x4jMrIDJzD5ccmL5wVNteAGtk7bKELsJ2UdJnmFfYNQNdbnhJK5yK/a2peSp
Qp3+P3zBf0EGqwL8796qbZZPNbxd0OXyMtSg9wDfer55cWXXAKVcvACs+7nradodAzK4zcGvmUD4
UD5wS/AuLrU5+Q7tkpiMe8p1c1XALBq5nO9Cw7Tkn8OZEKGqpxbqOClRMaHokptJ9PumwRTa+Yhi
jPydAIbMb3I3d54bGJ7tYt5VDnfarVTHQnjY0QnX4/8LE64xcFbfbthHWm22QydODp9ALoN6JNbt
oCbmzFPo6xbmbJlv/PDLrabVA26fPRxECZkB3cIxwxeha3o82wf+OkYSwz5wqoaG6JrzJ0UesKC+
3d3zX/aySIKl02oVCHnYDpsApIAIMEwUpWhJtNo6wkoPoFO7I4kVDLl9GIp+dd3+bKtdhNBSKGGY
JE92kzFOAtMsiaIsoDxDYVIVAuxRjOFTVwhXeJrxmsf2k/Mq/cg8rAzLmlveZkstVrJ1TGBxU0CG
Y5HXYVMruO+xVifI9SFEhoOpD6W5lgnSMSBLcR6gge6CSs8KoLOsFPjZ0NRI+f7TReoiLvtXXdKu
6zq0NTzpOZKZN3XH3qxLXl8Jih73RKEmR9sj7BRwVnCS6BZ2AUenWabNbaDST/n5CWB0dV8IlPKY
jogSA84agdq8HNyAJ+W5PxTtQOLVPG/X2fq0QyA12VhXGlCHx1Gp7jfXdE0MT1NCRmYEM5co9jed
H2FOpx9LZQx1BRcjOn3Lf1qG+evY5ZJh9MdR5K58eYWXlB0aN5CrMBmQE1CQjMSEdT4CEhaxUhqs
enj7BXpSftI9YYC4dzfIYsZUn/p8cJW6pug7kLU3eKfyC0AYwjPLd4So0kU3f6edMmfQvuK4aC+h
khFTa2PJ18pc9LGmggWbLvMTO4DOTM5AlMZ31bZVlof5k3xuU4wjqPurRqluMEyxpFi4WdBA9PxU
9prXEKIKCgHhAP19mVBx7Rbwy7uuGuOtUOtxE1Qj+8p6Pt6I2EePPBaBi2HQpgwFiWEh5ktKxs63
Adc5hyg0R0RMUPH1zvTt6ZVaglfnmWEz0gZc8Pf3AWAu1QeWEw9L3qKWrxXmIQxcqeHmSAqmjhaZ
Cv7uat47lUdMG01D0ICvqGsXvXpqQLAKXqU8z2dBfNhvapY/o/nvaJ5EZHqJTzK3evyWhRaHLAkK
oa1AqH5Birk1xVsirOYWv2w2bdrcRKeV+ul6dUCm4NkrLadkAdyhx8J+GJT7QHP5J0pnYgV+6sq2
+8/n9FGNg0gmA5S4vsqGAz4QWnEtO5w0an5Be+hf8dq66zWS0jVxO66xLFrLcYdG6tjYyijDV9bZ
CT+NujYaX8XAKRYDsFN0NAZa0QHTMoHr8ktK0zO6KbiHv+cZl3e5P9rDUKTqQ9dPmacB8JYzXe1p
T12avMjp2pygSSdJTcsBF0TAWBPJqA8GG5ER8SlDeFb0U4GD71PWMXOTta9xNBmDBHxGhyWJ8w61
oCm6e8t4qzalyV1WrP3BbHZu5kUS2OzrZTOww4GPSjwQC6UUg9bv+Get+RqGYGRPUbtt+DlS2mSe
P1shryjsXXza4b8XOwpAJeB6z4FYUHbPAnS4Y1O7jPEEDhd8is/AK1q5R7L2mIwROl910xd5waul
IovLaYzJY8xivYZhYZOUyhZRHpss0DJfRc/0PxWlZfqa+ZPSjKG6cspzmjuJOCZvJ6cDsTueEVB4
QSQvZXfqKEinM+U4yvOleIqszTEqCAFYNI52obpnQEBVoX+Sqcllo8dWYn6XuA3KXPAuty0Fdbqt
TjMhurfm7jqnppafI8q7Eh7cVGwyFe3zv/JceLDvkwvs2co1xMy+jkC2vcGvn9q6vASafhRpoR1f
Dv9XilSzSUqE+GxSHMWHx/Grb6xC4B/2FotxGR0JkLlveODqzsnC6nOFj3lxmFTSQ1IpsHmVQ7mL
i2coRj5nsuP3nBuLgiZ0lTUgBzpjAl16ue8773Ml1d04lh0fb2PqoTBJVNw49IYT1xCa9mC6N1Gn
H96NVxsG6u2KqeYj+KVwTL+7l7kKfCc+9PI/KSDzv+gsp48N2/nCkIFP5bBw+0c4Kcjb9QQK4Mpz
QU/v/HDOn0jAbHaoryB4ovRWgxo0ByQkO3q0dJ2gWQkMKmt8hWdJp+tvoHTLm3sxFblkIBPSkzXH
IudKMxw5wgHYt1A4ktST0qqNcrHaJ2EjVGA0bwaBL6cDI39td11l1nHWOnTLmSQrjMHhrQfnKAZI
SSi4asgMxeNUmBmRBTT8z3okrESSXiptKaUAXwjsD7PjV64VJM9rJK8MGX2n8wBljwwg1b7t4+D4
204BvEr3Dv73f78/BuU9vnZBmvQonUyUBInkRBSEvkTfzY9uVXd4/mF/0kSJQqJboSDKal6M9ZtI
gwOsSWI5zoBIGqOKRSca9ULKeKODxkkbRNu3TCcC5bStZN3vlW20UFP6ZjAaBskVRUuBLMhkLOPw
wt9gUCSAnwCaMNl38o36kXo2wJvqxbPV9be0WH5JJ1jiPido8b07FvW4AP4NCBjbdD6xHCv86ges
2oth/UhFTEF2pa29ZsBy5cPz4IG6fXXwAbDLEcgcZYBZ0i/HfSZDj7xy0KtDfR94ut4M4w49y6aH
lFij+HMzx5Hmo8jL/+oVQ411z8fdmcLu6fCJTTDHrXVan7rc0KMvvVDsUaazCbt8yKOs2qS/jAqU
M226zDhPz3QNZlJGvK8YZZs/7KJmRWLdt6J6HyOq1LA0lDS1fBUmhTyQt3F47Tu5uOsiwX/N7Djg
r0J135wBr1iMc1DVfU7f2Q0dRjvsykfMhKVyYRt/rMH+1IHVMiUI2Tb43ACqM5V1c7iU0TuZtxjd
62D2saGvDVpDKxEnPe4KZYTioeHs8iNr9l6idGlVOm13+UlUn/a/G0iUrCrstfQmgpxAdq2zMIcU
8aEHxAOamWHrLEDWAPNsGRh9Mhumb5+fGZPtKfsuBL5XZTiWzxT7N5X2Bd0eJGR2EZxbl6ZGSBby
AZ6W6kqYz2r00bMMmDKVZq9p/Gw88AzlKxFdo1lO89L0gsQlpb5rsGI6jwHPzi3ZT8AENlmrHBjx
umxQxVTUBSj73LYd28ybMtsBbqNs9mWT/uZmvGlJcWaSRxrlnM7/9uaqoBUPy9/DZAvvPAaJ5PHZ
sk+o129hJJdKn8odAZSeqGpve4v1jEegSG7ao6/Wc57Q3Ze7hcn0gRWrdGfCg9I/qLyUEWGre/dh
v+w9vsdXHbd13nCzmYYYU5u/VDItUUKvSlDV1zIY6nMfs7ss2USlecMeUoNUxIr9mMQ2QL0xv0AH
brUzCANNO+dQ0iZPzsE3c/XuXeGbPUWY4pHWyR3BaehJk45GYOUhWDKxhPI98IZXqLmTifqA31kb
fsRlhbCeW+2Ev/2h2sfm8eSjUcATXg610sdaSJmaAjEhgPplHjXAqaosgTKT1Hok3Ku/EM08Hj4o
5Dj8eLOHaHIOasdC9D510bgqERQ+NZ+KLdOvwxml/NKlWgS7PB3GtNbPPPv06NiNQDrPIMwdBB2Q
FzK2xazgDuO/oWUO5W3jb2FPE5Ii1rhiz4DIcnh63jgyN7GkLfMc9jxA8WqqDhMgJmvUaKKoxQOo
cuk7AEI7MI3KfWwpzHWopnAg0VzhkSqeUh+J7UmNQ2YxGiNjGHbc10mpEG5tUC5EKHp2QUFFruyl
bZB+ylk6EKBw9fujKImGayn9I3F5k1adU3cubaGqcR76gX+j/VeYbAgyMS5ftdVDCdEOAC/0bEWm
BRZN0+lOp1u03Pbt6qiL0vJFZI3B1QREj0YXh3tOlPTRQ6DEcDwvZxWQ+3LwElo41oXJfq0X4xG4
Sfh0mF9mPlhCst5gMwBIt++/sjk8LkcJ9cBoYsDbtEvsvCJ0QDy2GYKxufcTxpYIJ6vd0uphyn9b
mAD0IEW1d+ujh2uqgdFIkrOtdEqAHeaD2jSmaIOP0MOXHolV3eXp7fJstqhBuCpEwgjuX1k/zqs/
vO5l6KtAO60mcyM5gzsQ/WsQp6B3BN+v1h8KrzfNPdw3Fy/Xtf8qPiwXMOs360RF645dk8kCtotA
gBogQjUOIA5wAXxm7jdkWpMDtr5MQPEYmUqTaAF0epIHQaS3/7/neHDbOQ17I7/USfVUk2D05qPz
Z+6eEbyZkQxrEnyU0k3TOdVezuTTrdbbwKP8PqK+4uGVKIio9XiXioQIEqNXG1bIC0ryi7Tsw1W2
dE/Vr5LLQ5Akd3rTKF5O7SAmFOunPclvPBdvd1bF1fI8z+2gvjLfRuTJ+DyIBsi4nzDngvDCmv+e
icGnDECLsZzWWL6eInI18+ECrMgW7fGoYtG9ULNvQwWXQnH784zRYl7N3/NaCYca5SxbHvfxfxsI
mUkJSLtnIPbEl6b9S9HAmr76KhKNTwJKwWt60MVmcsTF0NZ7g/yrDpxv8ZZ33V8fP0jhoClvq5VS
Jxpg54WnDvBY88GDDawnYvcYwJTz53MtFEkvO671fzdPdR6c4MYPI2HxpRBchVt89zCxHUa0FlEV
AFuw/9O2vD6Kq8fzJJSZVcaymUItY37NR8VmGbemtyUZWEvJt5kjk88k7k2r3cx3yN6RZKWwWl5F
RfKLp8cDhJMvAQRVZCR7R/Eb17v9/b6VNDboME73c/ax989nYpALS9ynIWBVE88Gd5vRTY6otCnZ
Kz+2upXbT4KO/1OJZ1yG6iqyT2BNLV9RbYYN0T9ZKN+leQXYY+Ldn992t59yKgpx8Ln55NHkK0bN
Ud9fXTMA6N9OGW1Un7nDgt7BwFidURZSvdOt3U+jlZJY2QU5u+Ddp3kMzee/0j+Lt0g/tUobYO1N
2IEhYMjPHw8kWK3ZpXGiyMW2XmWynyC5INruF0kE0YWZlvooXVRXySv1FJsL0F6jh9FHp4XvEdYB
lS64sIczJrFuusuEPlFpS8y9SEWOn7ybfpc/5rl93SFUjDaPmXwj6vnbmxCY8Xe4/9H4mK2mGbVd
1w+vh8N6lJkfZK7rPn3IJ1vXwQ94Gs4DL3Y0jBkq4wiNelolYZ+5Loj+uxfPaFuoQfTJnwNBAx3S
OEvnSE03LpXhu/bqvaSwpdIWwweCytju2pw/FDhOPrw8QepelsHCEeNsjcuNujwWzIiJR0NotkiO
HSEJ9Hf2JxMwR3a6ZA2Y6N74zaiuiI9piAXr2i8nkDtnGVj46Er1NTRVxEfM60PCNJfg/OCRcB0Z
h6S4YGfn19sEHDeDUiew4TBb7Zx/9hfQI1zB2RvDa3n6CXjXogjz/zxBA+rviyuIAeCeGtC3zLA4
8RY1xjh2Vmdjk5i59dFZSD6EUfQM63mZIEafX2FkLcdGiY0NTqw96x/dwn1l7/tv/XYXbnZ0Y/bG
CqWwoYyXpcvPt9PyyUDbfIno/9VHXVKL1KxtD9y4ZBNfvXprT0gcRHb2cckP/U7LMFeknUvUCGHY
mb5VdNzmVHHnQPP2kDGXGuWF5h3CbImJakAOS4m0CQdMO0HOpXnNYiG9kdcbNTB8ac5Ttenpd61m
2O2C767OpZCdZzyBm4SYcG/AnIk6ik+kHBzYYUKkGYVIr46cM/HjZXB9J2tpt9QE15bVnenBcZfh
w9u9lyHJMZmunqlSzF3bs2vam7r4mZWqRNfWWfgWWnwITw9jAxtGduQGtKJ+3VsDPFz5RrgYtmu+
IEb2LHG4WfkFWAPCoDfmAHiRpd+8QgcfCZXSGaMsvMv6PH1UnBFKyPGPqZot1tvsZVXa8pBXfN3X
QBBSCMOasdWjBAmAAaP4JUVCEFqv/eNGMwf0HS/v7ESuOWh/5hjmsb9wcEyyt/S69lGXZ8qmXHTu
8iihw5rWfL0DcfcoQEGfmqMiqWKEhDe983CeYoxr6uvbrYmfy2BXvDZEmE+l9MvXlAJe6O4Lzh5/
WBhH6aPncvzG/iDD5qZLleCjjkRJyQoDgsTw79ruTogUtLOiMs2k6fNG2iwHq8Ke5A7e0ENUUn+f
pZ9H4iorqcYB4m2/uOWcx2HYAibYbPdUVGrN5JxTm3ezjeZsa0GnUUyFN5gydJq/6+WKERa5j3zt
zwycLhz+/4bPCXmTRWUiZJIuZ/USzHO9lE7IdNi+d0KTcUBdoUd5Y8qfFborYTa0nQ2DmZ7ZgAx9
qcrhnvt2XznuKP4Tnllt+LIiUbrogWLU9oA1Hkp9QuJ+0AtX3vZVl/FeJbI8otWcy4U9tAHD2zv0
OBhjHLmBa5umRnHw8X3S3lXcxx9wXiOe38OyEZXJuCVcLxIIi1V2/SCyTzFd0JRi/P/AgOU5Vpj4
8NIk6bGNyaB0crla7NxIZOjUjLYVXKIRMy4DfgrvwYmnIlqnGp6R9ISOtBSfA7wcFw0zi+0l9TrP
eElb2izCy/rQwqTzD88DdiKV/awymu7GbNifXjreDzhB+U+3Ywpc7/2yfFAmtVMj2wSMcgkVR3nm
0HfjeBGPXOpMmnCh5SVNjWu+UgVwr7BTXNcYy4a1pVahdOQ+B3BncKhYbjHxlvUVoyngfR+4CCQr
a6+9Z5qFqjfzoBynCWpjSRDVxX6BKklR8FvqfCCR3gJsMI2OQ1wiz6tpx+wShDh3rjpWXlaJdrMJ
bAWAL69xuR1vSCpclnD/fTZ80qU1IL5zdVcdzSTH9gS8D2NS3eluajhzBbDvBTnoOJ3m6sunK56e
5asYDKoBoicLnj2vBgJr8Q5PvohcE7rLQQ9DYL73FSWRLhyqc4oUWn3xSSGjXOEOcu3dVdxAX1Qv
8Ah3YqEPPmGhkDtTW6nCT1FR+CKCCcyX7o8q9t2UR+bGIUQzkUiekoMutSmm77xXYPCjS4BIwiF6
9MBca0U6vccW+aI+Trq+ycdK6yrVUWHrlRUTiztlH/cKrtUGuhxDvE1hR9KKvS4oJb91p/NKZLov
fTUkwzN572PAztd4b8YWzqtP7/+gN62pEQ9xXOUR+M7rFojwYQGz88y4OoeJ9v23YNTw4JOf7wi0
6BwxCm09a7Tee1xEwMDhA1RbgBgrRm55VCN5frd72l57kzr1HCD76h0O2aP60ZkESVe2MFZsQwWr
9Q2u+8ahbSROyfkATwRH/g/pwayE+ynQGOp71HfJQWleGO2An/NcrvyvUtTAlDNJzl8aytID/PMq
1UcOFaMo18f1HcUvy00z4SXlrjiRZXkW7bD3jykIojdyM2Rdxx3gZCvf3x2mWtNVjWBg7rGyHzdL
ODidD64hpQaEXhWVp+eeomD4aRKJWYaSoobJaTjePbg9YU4BFR7LaNKCkKpaWEUxOmXnUlLQiFdf
xxSmPOyppkYPg3E2laBxMCjxwA2TjIk91kI3JAzg/JzteMqRG3BwilS6KDMbM/xDa5CCYqLH30IE
5B63V5Y6R3bSI3aDkJV5M0JUoPPImhmK5ZzWii6VUyYKOgrkeWHLopRLM2rtNcczMk5doseTGp9D
kYNdOjzH2+2KQMr4uPWX9zUbaRJRtjSxnHoBEmOY/ufMygxQ+7jwaKvLhl/YW+UXtzftJEOqqbie
0nqP2mzXnYazQe+R7FrUipQZR6coMPce74aOAruv4aaAxAo6o8ZwD557O7U/gsaI4od3iJUSxo+m
akmzr+EwFqQggvHsbppW1kcAVb6Av5koH0kvkTqT7hmrpkwOn/p+kNJD/v9TFzq8EURbjj9Ft7YD
2J6rBrhdHTqez/ke5PY2wFa7ZQs2WhNK0WBzIJUzIUI0kqGgU9tPI0T8z4d4Dy0puWBzrEcvMba3
XSpw7pWOgZAraFBxAyMle8bdVKBNf+wj9l5dEv/bWG6PIFyimxOaFeKgUE4CLZuA+p7kJFSY8HkC
TXX7RES+RSNHTiCyxYfj8wjLoEGowsTrPVY+t7fHAY1r/UAcpaqzHg2QuqHtcCBJ5u2HP0baQBVp
j1FksQARDyVQqZnq2rLmo80ijHugYZha9mJTbBXtb9xe3a1fo+RtFaJSYEtsxN2UeA10KASrZeuT
CtwV/vP+zV/egakW4hrzb7dQFDuOttMQCzGYeBr9gYHLc2OrKtteDxEpHfB6yGOo/abJwswh3+Vh
Y1/DN3o/U1lMNBiX2lIfrPx+HJI7XB2ioeldgNU6Z9yGPeOEHKbuIgqGWsBMCN9ZFgRD1SkEcDFP
T7yUFNbYbP9c6x2Mk6UPFUqKcdNGbxYE4m5OaaHaMu9NLVEhjcAU/V2XZUtlO8o/CmxVGikpS7Ta
/V8GJbc+scysQzNI+DRpn8vN3Ojw48I6LAWsffzD/9WxdFiB0+/HuZ5C0nQiPNwkMYztTc2CRoPE
iZg8y00ia3pBHaEplfWEK2DPbHeHTlxF1PqRj1FdQYJMeuPAJpBZGMAeda163fbgWj+BHpQ8/fFB
y71NQ7LYAWkdoXl+ki9GqfzXCfpAzP9ngyT0NdA6dz50h8kgWLqFBKunl3aAAXYxGkZdMwOXjN2O
/FiI4/TlgcgGv1Y8nOwsXvzKn0UZxDNVZ5hm2fmdY2a/HgcUSphS1/wSfa1SBmqOXTzjRj3zgy8z
j33uT1QQ1S/v6bbGsLULi4MmmoZBfs0aVkD9GvLZQ1v/t9vGpSeSSYDpVz1pd44K2/E90BKu8NyS
jHhicL+rsThol4aY5BE/KdLbhQ26OHVtrKf+4N+/iUEokP6+/gheqSHuYe8MAiI9L4DM/6sZ70eL
NwK01JvQk72HdDpgVn4DE5LMbuX3vK8Wl4MxSC2/g8Sa4RQERt6aySnZB0EDHSy0ZMHyIfXp3F66
TUrFFawCyNUPRxZJcp/tokZbVW/WknOpbi4cuRw2VScNdfttipT4twCysof9mp8T4W3TqMS66fuo
cyZ86pRXgwH2yzCXr+SmGrX//eg7c+4q+eZ1X4VMWFgAGOqr+r9L0DTvTprLqcdPKu6wM6dpFpRr
hUfFT/u26LkstY/4bIOfXNtqMXi8BrbMwVdPOItGCloYGJw3LEy+rV29clJJD2aGk+iQtgfFKEP1
W2sRz7hZlB4/xTH4MkUHkxLb7R6TyKZhOuviqvZqzKaEHDhBZlRk6iy3NwutnxzT7GJt9xcGTPFu
Eku66p+hwTNdDi/n4Vb3b4fAemcTDiC7+nBA4iN4Qk0yDaPREDnBW9DqHU+CxDINy/ePYkRMAS0Q
DfJ+AdPtZObn585rtxqsI4e6y/bFiMhbcPYu7N46cE7P0FbUCsAjNmEdLDmLWRgq8Yua/AP6BeED
J+xD0rezAaz/+OsNXTugqGpzLyGVb8ioRRR16YZNq6/jBts+nNgEMT7hNgd7cxFIkuZuJAjPHl6O
4BabOWvxr0VHcxwf7f2rwPvhE2jqCXqVEoUra7MGYVIHSNBIMeCBpnB/+ObSKSkEb/HRt4zAObfm
VS52EGMqx+PLyvrurAyVVdK8PGlPnbwPjsCYHGZQAtyaOm7CmU1f4zDLc4lAzbNxTRp23tT/V61e
x7GzcOSRys1l/KqTsR83zjoW+yoEMedF7Q/uXXMsnT2pcXRsiQyUW5Xbv9JDuZ+fEXP8aVIJWrfF
w2OCmRRdxjtNPkQMBik2nsKY+PBxERlimAjs6b3gPh86NcHWqt2q4zl9atXVe05MJGyD0lMIv0Wr
Nu4oTiQgvPndBsg/z7Xkmr8hmzsytJo6UoE6hSY/jFu1wCl8iSOtagepvbkAv0G7bEt7X5lZPThV
NZjW+hbesR22YGACwxSO7HP5ExRTTCmnnXCHzeEzNxFd51qL1H/0JV6xBcrGPc5KxXdOkxgFegCZ
eV9LONimcRmBkjdRSctMyh9T0NSykkalCxfqvmpbHsfLcl0KJHdAzWaCA1FLzulGNerEZCTu9fxx
D1G1rAVHa2gJ3XgF0TervpXaaKYx9iVl/xE2YwDgvRRD1BPJHjApEWENggUutPRfjNySMz/2/3Nr
1X9oxhzj7bxLaH5vR5iasaaq911oRNLfHmfY1XggF2MGkEHq8mFmpsAx4wuIudvfY1P4n/I0sck9
/SptLz/8ipaAYEavY3BWQg4HWl3vnnYjsPLCTSR5mGoUohrZKnXzdd1Y6Y8HNATcLu7uXEfsVUMf
OaWyREysZosJ0+YwQwunpysByW5kwJejGUOfm43r49PTvXeARkBBx6FuPrH3iTtQFCyP0wJ3G/mN
J3N1as8eSmzJCjYyPIv2p/CfI93IbaBOHMp9SEYctk7W4Y3wZjnDr0FWDc4CtqKDkpS3zXv76TkW
CGd127dZ83PUnVtKi0aUCLvDKVcY/B5+bglvqNgu/Mi5zYNt3Qlkmq80co8iQ4/xfHG5X2+Mo9h9
4bnvfaeWRwYgPwfEqQsd6qYa6FIIzY6e7IaypZ9cnTbNd8F60SYuZau+Uxlr62WkclqXPN8T9TEe
kuYfEaj5msww/tWESicWRJRRu6U3RMRxnu/emFVLI1aysXcLHM1EFpb0v9numTRjQa3GhvPf9wwk
LCjZmkYXGEp+nRG9WiqvDu/SMSnu3K9SqN6SXGhSVw/p+UMrLQBak4tIk/WHmpZQgThGcaY/A0Op
XtTPoiErxHVgfMBX4WMCv2I0LWmmaXfdZ3McCjIreqR8fMPACEremhs9qoObE+/qGK5kAALs1HH9
MK0oRM5bcuuMzxoUMRPtKG0bSZAw9mOsZ0dH0rhEQTdOurlk7FTiMO85yiZvFcGpyS40Vr84z4tf
+cOMYRxmEr/L6aqcmad7wt2PJM/oqDUJhPPCb5xxXRTe8LSzEwise2j3Ws/eDhKWQbHG+XaXjXTw
41AeHzjOpaPfHObGDTiR0lBZoifrr/rJXZrSJsKkXilTEyR8Qhbh8ea9VDi2hCsFDgapcKK/4HrN
wB7gchztIXcx5IZ6NsoagOWBfPC/HYwGlgTkyFuUcrDOD54v9/JFvId+69lrWHHoVaKrMgoT+4Sc
SmsAq0nT1+xk6YZDPLPvWWrmxgz+1VcCGQc0RnrS771EdnKb/0wI3naUleII5IJg+QPv87sqbWsY
zeYXv2WrJa8h1I/zsgZak3fU2l8hhNTNT2VR3Io0r9nHl704y6OicokcQF0J1UvZ6SLRbpUDUCHO
SgMQjVJQ/dJu3Mutji2WxD06likuQxs3OmZJ5FXyjOrBm1ko7JcK74qogzxjanzfZ3WyjRb9pmpU
kc9dplGu8pkZMG182A6cUeLsWsdYmQeGXKokdvLkLhId4KBkisRA0HegX3DUoLTG2RIXFrzkgS9e
Cm2f+3nYL4CowBeqSHMcJuM32t+Ip6SSChnEkh0Ss8d7Vi0ynqXRIcyjijLoBtjQnb+jBj4i+ga6
tCZuw7GMU2prA63zPI+gHlxDt4HroBF/klUa1PVuRpjohcCKGdkyvYEOR7h3WiHjkKq/h6wne3LG
fVAX66zre71EPfGsCZiCCXwIoF+oYrMjmQh5tSD3AW/oHH8WLlacfAplBWZYvjaI1rWaFZFU2E7R
Km1eRDIzP+DqIeGfEjpHzE5gbCpD6g2eSiVkF1NVyIbEl7rCbFGGVkYltfq+d0dqkRAAqPzSDW7N
pup0Vx5U/miXlOP99W/7bi2MQaz/UlbHtbCJP+APw8fvGKOdbVo8oZdlvfkDAKXN3wovlTB1TQfE
ebp96DnU4ND33UqEEIGX3NurKgXe11x/9eEued7pDblCeUZj+EdLiscWk8pSk1bt9i/Xea9Ge3kW
FuR7KjDhJirLUnNd4pMPGOf4aaVgA2K7GCeSZa1vzYDnjtyr0YteSfwRxKQi2binTOSD3GHbP9dt
7mLrUfkp9oUbnYJtWJbYX+BN+4a5NHfThk0TbZSeOKfU/qQzDx9ZZNnhYC/DvzruLIvm269az4yv
NbXeLvxvKN6zGALbwCXNHgvf1Ery/aztha/boVUAI9J7vMuM3qUGUfx+l1o7GG1qVGeEvVfOFom3
Sp78bvYkfFTnn9C4ZVAn9Ov8Ep+fAigWFT27uaWXlcpwJSuN6DssRYiOMzs5/utWe34L67LgwclD
lULG1u3jIim9VDzuIvAetp/JcfBUA/NOU2qpr1+H0o/WyNo+cG9C7QJ6UODxhPvpMXr0lpwApxAO
NV1mORlDP7op9qgsnZkhHOdbSRJi7ttc9JOAo+Wq0M2kUuvKAbEh01r1W5QT3afjxk9Fb23TM1D1
nurbMCMNYjCCdNV4Qiqh4BSxvWP+WSIOGyBR8dnXz6DUXwyyZx/yVPa590BDiCqZZt6sJkeLyLp6
4yEIKcd1M9MwKV3qjqoEt9yxJL2I36SEAYgOBQP/R8Ds0Ia89P+vRVz7CI48FztMWbRl6J4T5VAj
nUhiFLSAfGCJ0TIyzW+OhOOEH3TuEQXARVKWhmosZP0gpHAjvF/ee46/4+whwbZ/maik61wosj4C
EMFg5QNhhUrPZPJUA7sBCLIrqC0oW2jYR+7CiTSUioCoo3YS7WUScMrpbTMlJFhPCk8kBPc1K9TV
47nyAo0XMvhmit80lZsJ/XKK0GusEGdcC6W5LEPHAIt35JdpfS+8ZL+y6qVVaircH+OPpkwq18e8
dw8+ImbJNgaFsBim4O7kZMo/Ms1eXE8A5H30JxoTXaH/oSKYDKVXkvrYCPX1M81ByJ47L3Gd8y3W
RILyyVUbjiWPvwjbd9+zx18BsJaXFWYu7ryXLQ2AAdXucdXBg8cfNPZD8BhEWmDL+3N071NjQT5N
pz4pAmcgOG0g9QYYnxx+saD3iOcnIlKmUIXkqsN4FmSGfX3UwyxJI2P2j9A3iorrTyd807dYX+M0
q7vvoWVXekPdmAD9wnRx9hqiAPKkvOu6ev6DtIffV7UPJfyKMUP8JIzBP3T0djvCQ/p/URHT4MdL
e4Pf4nB/5C9SnaL5fqMHDODImMU3ssgZKXKHtZ5wKnh7E/XLV/MRxh5o8bul8czSM9ls2Ow7Qzup
uBX9SpNJhjpiNYkvFRbIKtlFu/tWvneK7y/B4bs1T+PY7sh+ax7o8n6R/TojXmHwr+ArneTptwI1
O7+F7SLbn31uVK/WT6KRPDi/pUyfXohNG/eB9aEk+wA9STolaSPTNUXD4uNuvI6YLeQ4taiELpt4
2Yn03LMFFEFPQjCOqyJCGYo/CE5AMcKSBKyDLvvx3ALMvJ7EzeTW/0JwRBEVdomvEft21M9ZTrJA
6H6nvqRjPRs+uVO+OrI1I5icK3EKvs7tptghGdxqNplD5VXyDd4m3y3OsOHv54dw23SEZsfZQnI6
bdfs3dGwAlmGlNyRHyYzz5aWL+4kyeZcBm/6627dI7dFZQRxIQzl92p6X8d9yyzTmfnEONl5VofU
3EN3Wng9dLeJP0p5oXgzVewUpwY5v7crfk73modIhp+Vsz1IgcwVpF7/2e1Az9wr4qfWSBkeEgX+
Pw5opIil2eq0TSF+7LPEBf6AaxuT1o0rbOmW4TBXPppVx/Vkn8C41MNEtyZBbnqrrg5wm4Zpr2sN
vnhH2rFXJgWBE5vz1BbJIqQoNwjdUSiHn+SUctlZXcBFN1kcgMbqX4rB4nEMSGuP1idIl0wbxc8L
DPhypB6HYjkSww6xbeI23Fqe2F2SX6o9pc5PlXS6FxIhMwcizvZb9jaAHEh3Kuqiu2aHFOKZkbEi
usCvRSC9OFz28RBwcbGz54X0Lx/Gh15dTksZNwiowyU7h2Zb2Qx+ZqL5epvJYonybwzUvywA78yZ
I+MdKPXg1U92FCS5osTE1LpFrVmbuYUIYSzX3wjh4r5o9obgpfk8C56sgvqA1uMN4x0riVzJVyRg
1hfpeSJrjzSofA4dXXVDIsnVNPvJuJgziR6NgJlR6ZcFRgdpxBcznsZjjTc0hEG6Fi8bHxk6bCGy
mGiojcdO0+onyfFrsLdxPMfAJE5qaJTIj6/dUS1XX7IzUGomylI5Ybd9Al8gXcyFaVFVezhBM9Fc
PHxZ6yhE5ef+rRLpzivQCm3mrmCHmPq5L/gCWW/zBq/fNjWJOoQF+vpdOtjb5XzTZh5IseI90KDv
pLsvxcouWmWtGV5QnhWPq3AcQryVs275RycBxf7SJtgG62m14/kFomyZ9RekiWhrGqkVt77/BC5e
BrwVd2awHbOVbjeWjH6tqYRRrOqvTNlXkMLDWBYO+B0bI38F1aaff+N5foKIqTflbtfgyebF9xA1
jg1csoxEUXfaQ36Qd42jJIeplbX0I93JMFOn8iyZVkHzvOMrL/+pE0y38osr12mltvEudEJBb4EN
ARpJnqrmPXyd2KqjuJxp08VYiyVktV2rjrtEWEHP6wcETRAZ2TkuQsbDKM/50pwHz52Cw3I/CRA4
KepzH2F5pOJiYVSUZMqPqAmB/R8owail7dMQ49F5NPYH6XJ8qquE+CnPJmVcmxpV334vfGhhba+J
R9xGTHetELB+NxT/gIjDXDWTofVm+FTNJWMmP21RNhnfluAZdTPM6lziRNgF2Bq89aUO+XYVO3VV
FgOCE1+l3Ih01TpQpGuFkyP8X9i6XM/9pWxkcuMc89iu3vWTVeQespAT4srZP1a8+2mXBfOpcM9u
V/RK+z7qLsobLh9iSuM4D+ZK/0FrkFxUMdDcptmnsV6WiBdkHh9MYozrNPcZwmnhWR2TcKNmjeSK
5mAIr7ytMM4LZCz/kGWQSehAXuZ7ch2DGZLoFXqOmQa/BMhjSDSCDsYnBpk3kKUv+kY4fEfNJ8cP
iGoNndUOikMw/Q3zht5q/zZTDdPlhuRUJeFAeKcr16uZsx/XqU3cP5b0x4ikn37qQsgkU6XhkPH3
jxBzCg37T1EBL1cXiPzV68+Q7oEphQtymKyQaYi4b5CmzGRp2d/hQniPiKyWusGyzaexLaq2hVMM
oVc1knQNC+dxkhGxZC3USgSm/IXc/gzYRKxkOm6qJmt+nmCNZY6VgtrjOW2nitKKJhrvsq3nRGiO
ddSyJerF8eHJO2qhsPcnpCH3QInnWqXYuLx9S0w7emiIGN8NA5uCNxrw9evBW37DSJS+pO8vUivz
nKzyPWvwwHIpX2AXfN7smgFnokuRop49iurcFuSPg6JJhhDD1sYojobMUmFrbswPuCY9W89GkAVa
/XHwG1zzOdoCLHWoWoAQ5NBEmxY7IK2CxbJw2e+JtNufNJNsCpRVQ8wGXIhw7UzvqOtZD6XkzlOg
EXkV189XtpkKYAPKkKmn+/uUimDI+jSpvORvDYNsAsHU4Rl1OWu7zhDxg8/OPTO2riix+x/5wlIc
HgBWVdW3ME2M2GSGwf3ZxiSz4kaInsP4127AAKpmchAyllXC5Pmjt3oy4PjvvbAURxXazVpg+v8N
ebkhUONkileaczaRMgiO/fEExXpf2vP57RqGq8CasXhp1Aw4QvdI7NKXyyzK3vceaRoZL1k9DjHS
Rgw3ipYn3K0GN+7alD31dSEvDt9z3GwYt5ybVPswEYkMsyEdZYP5fg2Aihy+o1XBS3snxPZfoBYB
llwv5Z3TaloYHoQp41oxiHnjOssr/B7PutBmxNPQG0WMz7zZdjNPM+hTx0We1JDor34QBOPASIpN
TjfAMlL5RwC6BfRRjU0WZxfdZ0t7rOYR/8RRF3dZ03EUQDFiSn3etIVESFN3w4e25CtpF0N33qzG
x4xt0JZY9SHXmemDrtDcDQ+4SdnHksprFLeWYUVhK4OBBrMvRr034Mpw21sza5bJKfCsijfbN0e1
Zyh3GVVQ5iRXi+APxyfdbWLj72gAcC+iu5AkIuvJ9BzS63moftoi7RMYrHVBB+eCzX16Vo6kO9E3
PYUj85kjOpoUqRbz5miSiqmm841lacRawZNlfS+Za1e2CE67Jt9Nonx3b66OyTh0BBHdSu0tLchP
jKicO2lMjwiH8a24AZfiWpqHNVZ7TfldsK+LOcJRJK+BDKbAK3qP5nPmgtOSe4biKaPGSVUUMfCD
CgDRAl/3edT4GUJgc4X6za7X2juU8byNXDErJccJ7O1A3InD25eJKuruPuO9mZNMfYI3Jxcm36O7
UII8JoPW66vcpY4N0vXoSQs4023V4a9x7zgRRoa4QHq8IMgiQBTFwxe89FkNj5en+6IVChUXlDIl
3x/ThoSCtIXm4njeyksQk7L9nthFdonaDSnkxdFOrowZVGyFyVKFt2IL4bfiIT33kWMZlbAGhSRt
pVf0MPW1S1xWXF6dTw8SGg9uOhDlNuhcwtXuA7wKRMbYFwHZ8vX835Aagk0Ufc6An3ik61u0NjIy
+LWue9wIE58NqmxWGuXt/psAYhsRG8snd3KNELCuGzaGw84zDIDyIAeyqF8htvgEtQrnra0NhLEH
rx7SjyQzWM5uvHs4pUhzYiGHvJe5dKias3LFfyWEJIPC2H1PGUKMnQREl2iYiiEag7P7JzAAVelh
ZeFJOgv9gQLdlSCTvla5AExs4OyihTSZnKlPoZhQTHPPDbuKLovYpCy45Djs4NirlUPAQWSvdtaY
PJjJUIU+kV6IScPGhM9rC9QWTCDrQxswk5B47cSDoRyRp+JpYpqnT2/13FGnK1h68KlK7A8/2INK
fBX9Hq1DR0WeuWZGYt528kjB0TfYStwX27jQlbpjCprB3E5LcVvxyfOSLGOEyWjBCy1YCSQ6oF81
jxE/+UdwIaqnjU8kINDpaOSKrj93MXbKPaE+Evk9jSlPtE+vu8rn5F9ppTF5wUHciZDwKhg8V02E
WXPpCocYaCHXdwTrwYt/2hUKk2YTd78zr9N++xx+T2pfBNrRg8klDPq7d6syCKaTuPZWm5I7X09D
HGY07+hnosyJ06AZpDZ9x30mURc5eQkd/QgnOy2B4TYK+9PlQ4GzHo810QWrOO5NaOGRydVPRLAa
6N2JHJP1cx/8DtH5FEimDwi7hmc/ZH5iXckPjHCoMYTfTmUhkUtIarTmvcKNmHEflADG+8OcajiP
S/LT1LXPt4LeqFblW+4g/DZzoYf8CXmoJ5jIzYhtykxxaaG4ppG4goheDQNRsfrQ+EllvZcOiiRw
7uZWX3IA7cAg0MaeQoZyRL0CsY8W9dkVX6QLWgg1+kAxhuLygjI9jbOUhlRLZ2IGef56s5+ppbEq
U79DSUdiUUNuvh1GLqYAEjleWfcnqNVGLKUa9RuSQif3moKEYE0Sr06Ke32lCgOjAwBoEv3kX8lb
1AIxgWe8ivAiGrhrWeXMqHMI9YjaKZbnYB4Aox6z0c0NIgdAMfQlAUIiKIpXfzP65Spjnm1PmnCN
MSVSaGcOzEvKm68LvmndO7OY/jndjUBjAzDkramc12QdnDWGfo9VHYHi2CEkjogJnj5gTAVD46lY
Oo06+DBM+aCXFFldAmrkmCxfQPwfgFJ1bQ+sH2PmjIUxZ01QVHI59f83Os0BCuA0nxGew3tObVpD
XrHlvReLEX1dKj+u7J0FPu5HA2Pk6svibc7CB549VBCC6JqgwYH8o+CEtSjLGcGC51S+ROl0VSpm
H849SAuAAi7AWLwlpJeZYgbSEMobIxjHkee/sdJX6zBXbIj4aNuW2DD4XVZsfst3PvIBBFLHKCyc
rZIf9U/Lusz0MsTyBYqO1VChSgZihb7PpQSbX1BvAWWdS/whyEiBHUQ5XeFqSxpTcKZglzcP7kQJ
0NuqhjyklttZk/hjMSif97BMgjOpZNg+ksJboCnjkOz9DdLYLe00FHhZ+BFetX/EbwFcHMhGwyb6
hvHbcJQUdLDNnBO9Y+b+bZh4N3WrjVFuFWSBGuZkA6gOi6CKWPRoXz5mLrm2S1zgv3HbHaVRqtIc
1RQFT/ZU9/GqgOUTA59l4njsieAR2nMPO97nmj5f0hNhiTprlSJg1B1cLXndUoDXvIpaR+0NqSrC
EWV2gV0V5NDJkl3R/QtK7hDOsl7Vsu3NXbSOKy/aYreKXkBYQjK9De8yp2aVIjYRC7hSkR5whD4x
q3t9nITQdTdc+7pGX4MxgWdWZ1t2fGIp5VR9f9EAScqoicH7g5qHMa/wBAHVTzO+mev3weT3N4Fu
GpAb40w/o8PZ/Y9OWCt59UY+UJi3tS7u0NzwDcyV1fpKciCwZZy74og7xmpcntpCqHfLiFG+JK88
V05oRQ8+ZMhU/8SCXqbKvl1uGzn4SbxCIw4/5ycK8GIC/9Pry8sh24wEm7Zy51KHMJOR153qdB28
WaaPjVMgsgbrhUCJMMNcE/+d9UFhTST8H8S8HmC23++OQwC7hamQ9uGGrDuGNaC2bOEBpuwX+3zn
uNSGtB0uPDeJ1qxPHBx1O+V9Yq6DPz0f0qN1kC7T4Y+y+Sc1P3UO1EGSYaqAlp0B+b6zSfb3e836
5d4MNRLSlYiVoc8KvGU8uqifATNRXiHMdA3WpO9VoULcePJ2hJYWP23k13YNw9W6e33FPOxGdg7W
tehUhYRXIRctNA9+D7ko0HkBOpjmIcKPN6kYgdusUYcOa/bPfbcVyc+UeC+0T5tH0FnjF5Ayi+1O
drBBs5jazwk1YpH2K+M0orW4GcYtIE3xj1D/J1JJ+3zVSCefsjB8sQH159cxxF4aPpL89oEkVeYV
yoNovO94Q0GBcCV5eHeLTh6Beq2QHirPft+0ofLqYhPbOm+SVJ1HCsz2nCgjFvuZvRvXmpEr0HtH
/iE5qm8i9XmOpsjv0hQIEVRNqMooXqQQ5o9D6ykb5beU6SLS90CENHBfWGIRFeWpuwICUslT6i5P
LoVVl144ntBgkIEa5iGrZ7nw6ncb8QM5QnCtQgWO6VPUpolZJFoNdZA7wHvGZhkPxne1bSTeYPa1
E4C3yJVUrwtLr5uCyZHV8mCLSigXX/vU3Z4VUsdvbdKpsaUoMxmlv4EEkWk2DchOEZlcNRtuxoIT
vno1d4pG3kYtgRbQkgCTkW8KvybIpZ58WeWEi67MZh//Xg/KUDOKf5o2+dgOc1rOI1Vf8PsaJKWt
rBiWscC1aUV+TiYjD4Vegkag0OyqiCzWWYAKguy3tXQQVTMJ8biLh3LC6xS4UzNwxbEL7STEBkwt
qW6rBKvknGmI//xEmv8Uxhrk/A9N9op5zZABVlQhAiPahpMeK9dbnxqayyluJhfgCSxCfxn4NRjS
fHpX/D6sAreHqBUtchuyx2nxp7Ravam6FOr5taxHxuVVj6kwAinoX13BYpf0ABYE23Xg2CdZNJwT
nqjzWj5X8dHVrGAj78y5xIRHSD8bGxqebpQ/DbPiU53N+Wh3CJdTD9XkE2erl+/Ny84PPZrrVHJT
0yPfSCQQiIgzOdNqh/3mSTITTO1pyuUObcowLLEvQszCewt9MRb+ZtcNovWLlyFGfsjGHXA/GaMB
7BxvPYGjz2sr5VlEZuTdeqLfHny3lQJh5LnKfYoAu1DMeU9OjDzasf5ufmG4x/EnrObvX2bQxxOj
LTYpMZi9fztxh5zawdtDDwD7Nz9Z1f9VdXvsxBA74d7mYk1b3bhw4FYP1vpluMvlBwOophHY+JD+
/LlapaNdJ2iA0AppMSvFoUJ9uCZb2naD6ep/D1TNUop7prnbEt/gwPSD8lBH91mmrAbCBvARUA3h
qMsRinOACbUiZjE5Ca6wR3iLIjzTkhoQEqhnm+aPgJF4VFN6OE4tCITDogmbPrVXwt+PYHD8XXQb
uFsEJmDw0YhE/xBiB8sjZzU0bNLDPOr7JxhTw1WnNcosJnYievVCu7PshB1BnUQa/q0nYEzL/rJm
8Aml90xaNLv27LogAIt/jwKSjgW3r+k2fEeEM88ipUy7LaPJuYDxcuFU/svvTECwg8ueCcLFoShb
x57VbyBwuCeUzH+fcPQAjvpsnf3OsN6vWGYDNJrvtmNaYBZ8Yewh/oKIaCUQpLzeM1jMtINVZPfA
iY+fMkre1GA/Cl3LB/tfEzkJ74brRtkBI+MmTprhyYDw0nzBsv7lFsnRIjudEDXdJ8wI5YQvfA8s
rYV1iwpBd/TdKlgJOvELdLgSORn0nJ8VTPa6X+7PQ59ozdwGpPuLJLcu7HZkN1q0p4xD9SjIDc/g
m0uOoPLUiNdTRCE5W5gihyvvOBQcV4irIfnzBM0rXA2tNLTexfjg+WJ5qvltUPNeV0QBFXN2D79+
JLZKNcfMl2fXV6HmcgRUbL66RPEvj8B0XhKk0sgrLKdfeoYpUQADwbw9+MrauUCAOf7V+RHXsPA9
fpSULtHoga73LlNv2c1et8pAlqirBc7bpC56yIZSelTX79lpUgN+ebgPrMkORoQOgfKCn3S3PY98
01Ssxjp6mHIEaEyT0jQt2BLyOeKhrRBUOdlAYH5nTXYmTXsa56PHb5YC5Dj93L/RMgm0+V/zr04x
4kb9CJrtim07ZzUnlrMd7O9KEcb5vD9yuD8gO9kuLp07gN+lOraF4Sr3p/KUHn4YBG/5CKS1vsI3
Z0OAu+To2XFJmNNw6Q4r0I3AScAYqUX7T7m9GhdsoZpYO0ZzcjIJsGu9eOAiZKm8MAq9Flpbiby5
9IFkjOX06ExnYvdlVm+vzXGhUxsOMuACFczraNGBs4IP19CU3VPph3PTm550kj8pnhS6Rrx8gKWw
WDr2y6BiKkYERw6H3Ior21e1EbGbfQHJQ4wMYVHS3G7S6n+0WRjsS0qxZhrsC7akbIMahniYINBi
/0zufExPLe3t+AcPuT8dmN47lcNdFoc6a+s3WejaaOFjjU93zZ1yAIj1rczWlYejFI1YgvsSuex4
fdXTUOTsFhgrK0/t3yoQ0AP+NQkFgd6GGTjwhN4C5ehTbBEHqFbR/JrMwxj0fPBNss9LxkYyAm+j
coJKJD9mQXtVhhuSgpCpG/A1GSMiBlFH1VxNLDkZM6rhMLUm4CP+3q/0hqevpRNUGHA/SS5kaRi+
JpMJqiG/GmZIK1xzOxGGJQeQrw+SIZoFRoJ2CeFnp4ETWLQF2LUa7cjIVtCurCbBqblho+1Hck+T
xOlC54foaNtCsgbJlSu4kB+XhgpCfH+Pu+TLqfOOYaD4tMZ6dMMiuB2rgUZqLrok0vIXlbo3XVdt
FOE/LHT8Zu0G+zWvUa874iUE+cKVlO2Tk2IxPZUa842e5R5EcLCIvGJ3hj5zSC31+GjL0gx/J1TZ
/nmyuDuQoCwVInYTdIep7wLB4O/g0O8hsAbE9jClnGMXeB/DBfjwsekn8P5wJKjSti8jn+L9cByR
LKHqWGfUV+OsQiwurXwxPWMjl25mmxZTPlB3xfB6eRoAnPU0YIoWMtB1NGqLZdqBUddG14XdVV9N
vCrmOBpIjag6b303kPgrkIh+ficbNS9wB2nLI9lTFqSDDkU34hQkjT/E7OnVQbMZqNlPoH17VtOo
3F/zZacTJSOEe5GGvuWHftJ+kY7IDFkxWSUunU8CAIUUbxcZ6zv2jPOl6ED7aj/lvF8kmpvelt/2
6cS4gaGEWTDJZ3WBMp7fcJc8YSgSHdV4xwZ6XtQZtKnio7npMQqPCVgE3Ug5x2q3wgqAwLNHDEu1
42cdBBlwWcVJFPkPfERUiz87aoyOUjONLl7NjPaOqCHkPRooYSUWDmu9oDRVG49oe7lASOiUK2O4
+Eviyx39qx+zQQgNaSsh01cFg03rS3VHyYn0aFCzCP/HW43PeN6JuTZWdXflBIZpxHk5RWVrUX45
r3T931jdzIfy+DKahpRQ4qO3MbY1ldTXzynP+mU0GBu37UJPrggldnKGipvUuy98ruE2vhopBv42
4cT/7+/Xw7JrAQ9liV6waw1ptJwur5GIEFq03RlbVANj7N3tjO4t1XDwwDKiDl6QB5oP9Yra+G7x
uOOywpumquSkE8JdM/eGZpg9vvHlazF+wcmFhJGtcqfjIKlctMJnAhnmdTd886dBK8e1zWpPOpgv
8d7xSLt/wurcHuuWxDZ492bNFGaPbMZ54UqdEVvDkIcyCxVtnI9D+5dAjvNlpFvY1C/+k0szPR85
sNgkVTGcyC+hvXNhRNV1XdBDSWSrUMeDHlEirpXPuj7C4RFQIFhsjuKww1BIDmlcI6iMfftUm4QI
FfC5rMCExw54eDI5Uo6dI10PhbbJwjMz1RFAyj25ZZ+fdA4cmyy0Oz7+5veihoBvbbHVI705Qrf+
WUPAnlv0Paoy2Eg2JwHHm34ubdkHRoLZgde3ip8bx01BSfUKY9Jlscm3GLIEaAsLnwBXsymsTxhB
DiZ5Yk1+o53DJeh2IND+JG6QCqNqXBbJgR9OVFGMEtZuc1DN/9ik6ENLGA11YRALKA9r6nVyF2n6
Sr7FYvZ+D+0staq7zZezl/0bmQpekCGy/chWlFfFnbS6P2v6i7VffzILsLLR30g12SibnD/WL+9Q
xRxV2oSmPAgFJYTlGaVPIrEYy5QtaAtAp79rrKljjMmMJpdk0JqRSHmxJKWgto7nXtavrae3A9ua
n0lUt65iOO36eMTjX65uNM2B6uHerHBHXNFIdweVXPfWZrFxe1J1syeefdzhZeieOGuDUF9UhHvN
/lEegf+A8GtVOXDPdh/LQXG5RDDXIXuDQ1AtYWULJMf/YyBdL12s/hceW+WlDbkh9nxVjilq+DnV
vhYC3QMMvywAmVzQ7obFd7z3RfpPiWTki6JvUh506zPynsVSeisdlbOoVieouaJWAPnYhXhmrr6w
RXVX1rpzS9n8g40BDJm5MxgxubbfLvdrBGaIvsmG3nBiLzsR/alfCDe2lu9XCzflN1VoDrXmLX9B
N1CHXjgc2ziyf4tCO47qzbBi3GQKnR1YIAKTO79ziDgzSUJXZ3UlB9+yu9st9DxEE6ODgaQ2Zlfl
FPq3r9UwaRoYBBqC+E05LyZZHbESJiytsSiiE5bZnLhmO4nX0x+Iiyf8BLCCFPnH0uYzfbPqgRaY
ZCXe5GCH6MisqWRYA/QiJRWjT8qEY+OUx4nPiOTnj+0gdxpiMqS/tt/RObyaIuSBsNiKZRrQlaEf
6AS3/KcQ5ES8ugJ0XiJC59Xfv6n5rl7Rb8ke8QYtdjzjqwbTPPU+m7zw/bb0Y/lSE3zN+mxNr1rn
3THezFNiQfwTbDemsLyLxzIiFGf0kpI71FXCL7YWRqAnyfI8oSwYDd/lYlQKhEpM2plZA2WJFD78
nrcvLddVYaEySLHBNSmKvor39j4EQae59xwVKov5FBG6MBpWCjU+iyhlKXApr3Tkn3Jbjg+6b81j
pKRIxfPH0nAMZobP14eg7Wzd60rIOXN736XZhIUPt43fpWwZGuH6HvMUA25LglvLJ/SKc6NJUyS5
8w5iE2ijH3jOV0LFg33KWSRRVQdMhlLt4eG4ZTp/TYAXljBpVgoQT/UO717b6DQwBhpHymgofeD8
SZdFDWw6Wn4ujyrqehtS9hrzm4SJH8vWelQ7qPL/TRlv6vti5bwUHjJ2YTaFD5xOEHxxsUAup+Li
k/kNL8f7g8xp5QE2Y8UVzlGYbQOLzkHY8mHVeibA5kHmaIh8RqjVdzmv5ul1iNZfqdElBEzln1Ly
7Z1oh00oKkH2mQCTkIJJlJ5f88LD4ix9RslKZMb/jjPMrFBJ3V5FdkFI2Jx8VCBxkmEIJ4IdES/S
0LKgHqWu9SBmpjL/QmUjFK79q+n/B7NyxKdi3yhkMErSjg9xjwqUl7aCMdoxd1qXAEEHjjT6xZbg
ldzzb+tOsU8luD0Mfp499AUzaJnl44ToqSlYFc3uaJlwXTZ/aLAMa5Ef6Npqb64CZFcv1TvbUtHP
NKUpmUk1ZodNG7F6cQvgx9mkn7E/1RsGwgGBH1AiuAeN6FaMM39b74Ul3g38PED47bjvzUprxW1J
DsNbOMYY8AW3xhNeibmM3p+bvdupzSX7+8bmDrext1WstnaWOeyoEMyZs55RxNkR2EUIiuWVN1g6
UGpuzRsGDTf57hTW1Ci5vIJL+Krvzi5scXacdpnKKR1m7EuZL7vgaj4NqB9tbFnhH9rrZNalvOQ9
2gW5rSMTpWa1fpGXDmjWpTJHl6pLz1S7wgTOlO57Fi4jBOUhrOKBSmxHXcoYECEh9I9YMcDI4vC2
vC4Nwvpi3ph+p4MyMjCy41I0uLtL8FDQjPc0CZAPtn/AEICBPwDMMbne8PGpETiPm1OECL3yBk1t
55MgSn0Y6WmxB+up0fGuAuVMvv592588TUANU3o1icglRRxLGE1xLnl6EN2O/9uOM0IEeGmK998M
CffSRpujIUwHblnudWlbP470Mxg75xt0OJ+ihGYx9+E3gM6gKi0Lf4jN/uAlAvjFn9Zc4AQcyhZa
GSpwbOUBGbAObXfy4I3vQJPoz5UOxymI+CNm6uhAe437YowYZ9vuIms2gotru/vsV8meEC7242aa
UVzNtRuyERXtTbwNgdEg/SkAGokFnA88vICD983H45KrnDkbhTjHarYnZFB41apFevHhtfa8ehWU
iuobif7eri98lsDvv0TK1DTGuXC/XR90DdkKT460LUNIK83yq6lpehK0CFv3qFADRGdoBoFFZT1O
29wiUxv1ltKN2THlzPRnTxFeHiv01fRhuH9KFb/p9AzKZTsqsS+itsT9ko+zpFRlO3fw2hDQoNhx
rr+Ry5QqZ6s9F+lCyS3sSiszjva+kTPxv6bXZP+2aNdg8/6MpK6QKWZnOayjAWWEDsjiGK2Dp3kA
FI4j9IhOG1KFArSt9poyXUyYBwAecIM2Lvz6/4SXM9ZQThCLUkNTBy4//5/c5duKUKfBa2NCJKl8
4NJboZcx+ESggLJyXt2SqrTeiuguNYfcecsYFwV4IgyUT9sghWNvPEy8UwEpWI57eFOoW8R7jvuC
sT8Yt7km5md+bDDZYAFpVIK4Y6adWCJMkxBBQMFwJal8UNdJ6LrlJMxQYdvQcyx9PaiK7xHZCogy
aZdCk7VWE/y1cd8RWhe7bEGoFYrPckhA2rgT+2osqY7ZE4wsSDUGx+sJTN/IKWgQIwmX7HzEeCPz
aTbiEwwUH9k0hhB63Y5D7yO9ZlLTJrIlMdE2GklHwdNJKt1CErAi45T6MpRg8W0zrzFUk7PMVUh4
3oJHLbLItpDEPKg/6y+6+cRcYLGSc2231/VC5kK55IeFenI8d2iH6QHlULUs04AHQkBpYrRv6e6/
NNya3ZeSNt26cwadBOLInWORPsHKNpKwUabDp0czG/5KhztBzb/oP4V3/Qcwdc2YqSCa9X4CzeHU
NhLXMGZhpD/mrTjigryF52s2/BKPBVjVVqMMG0O+Pysn2grl7rVAixG4HMGfSZdV0sUlEFnYJXBA
sgLSdtHw61nvcz9ltTiEBKL2Py/9ZADDK5BSZEF7i7QwKXzLEK4/o6qaJI+jtDOJO9MnRQMRwrvE
AuUTaamLOoXvy/UDYQKLq+e7IHARnvWNxvMAhVDtys5dTNb789ObbbFeFxkrQqnA0hI6X7jGHoTF
3d+VDGty3rkdDkqbf8lnKKP7SDx41P2jZCb6+Ma9baR7wTH+VSfBDmsIlM8QpY6sozBZTxc8ITdo
Iv5goEF541fthuIlK9wa+QWr/W6JiDhiy2l2Gqpaq5j/5hf2PcfQG23zfbAjpyjj1+bQDD0K8mRM
8+Tsxu8IFOHyBb+49OHgMVp59SAhjMpsiL94aLnfqa61mwXHviy9iMglmolf7BS/fwH2Cz1DEhu/
faHVRkKEMifEL7jnpa7tyFkp+vtsQ25g2TAyIN94Kq7jSSAKBV0Fge8RGYG7y7+UjU49TwHdiIvs
3oj0W9yZgQxTRSv236X5LoOVe1YAQR2xh73EuxUx9CP3vdVn9MjCXgD87ooIEQiAsagohIP0BXgi
7J6yvvnipk13kYfH5O/dglMmMJAOKI/2K9OGrJzvkJkjrtXOawkk/TyINyoCnVm5GER7jPpRI5Pv
4t+CtCnYpKKbwnDRXJ/8kSHWHzu2NsfVzgjlA9I0okWa30CsO71rTOJAPYvNFu1SaaLKkwnMYcuQ
uwBmTpdg2cqWTfbz8EK0m4D6rTSbDgqycI4EeT2+qvrRrIqxtwTexpTD6RFaU5s1BvAQ5F0rR+vY
rFTNeViXz51aG9DlIaw2NWoreQ90K4zT4GbnQCSwQ+5CJOGDnFr2udvokWIBJ8aQLb9hLGK48q3a
3zYLfbX2RQBf4azjbrycYbARpQlDjcAGBeUftP9zNSPrVuSUoVLA45EdTeFFKt+Qgv/K5Nit3hY3
vYGQnUwjJ5tb3LJBXk21bfoeS5p0B3XJZ1P6hRMhQAsfIKQy/FFqqSbfdrfNk2rlHt7ggD60+DR3
ilR/Kbn6mXtlbLdWsvVr8tOP4dVvvD2xk/ZGF99hMGwH0qKyBoImB/L4XgAECH+qYKQXQPu5276W
KL7ecXT3tFPvTn15Q0PZJpz2BKvy5IM3u6hAtUDZr43yIOwtEX0pAQ2iTO62beFKqpxM6DS3aGi7
kYXDjxQD5F4vOukWFNiQtJjGfYyy7KPsRd9bp4mJ5fKJhm4rr80hDcFiLkPKaq1/zaTzwG+Sgzy7
fSXDNJxABVfSMt7jPkujQG1DyDAEcmhxxDTddOQZ0BTHv/DTcGWObyNKrAn9mZRgjqF1cH/NadrX
zrZs7LGw3ZltIyJa4UFs4q9czdPjjq6afwWbNMyGVhrgwSpe9DeACYItXOddKg5X5JPmnjATOISm
g797P2E0hDcKENlVF7Ar36uA2pntCFScd+2S7oSeeJ4BEGWyjwB/oU2o2iM1LAnqBzA0pPROixoI
XH/5Z7gueWF886C+qUu3VtvXEkMCAW4rPqdPaYyR3vyxCdMbDtRiW5hbBKVcN2cF2OZ1QToLljqH
Nnj3S/TGN+gy7TPBkosRglYIVJcHkMxeyZPQ8CMtLND8/9cwRy2n31T3MU/gzZW8wR3py4Ur+5F4
XZ+X0BrUBS0g4jj401UmywT+1qwVtUrNH85CD3EX6DgzVIIoAG4HJqNlg94gaqCgEACV30T7Ksvh
PAXu4ff99dk1+EC+dzAFkd+ARpDSQMSBiXkKN4g0wXFQLNylK+Av39GVHu1XeTRZaFJ8MKkTFKS9
SgK5DfCsdCR9q5RP+F+s5sMTBUd31S7nBpQcBSUug8xKCbmpNgD5NZrwk+kFREAj6Ugp1AEzTUgY
xDCE5pDIuJdRk1m5cuU9j0xzx/eNu+e7HNr7h4g9YfnHEN2j9V42jEG+zrPZ9bPbPzRXgznuVGf4
+q0+U9JarLkStW1A9T8EEPH+UsLpPyu2NnkIrZVRR7hYUe6ZTax2UgdzYBoEJkqNeuO+bqTScgKQ
j34wK3UQ97uzmTshN+hu3C8oaNABni2k/OgVqbLW6JT+2pIE0qIXB5K0TiBJE5VI5lZn9UdRw8YO
9tJTsAepZppHVGk20KwjzAHxrnYJHooWx3zi6PGB8XplH4Tbl3L2CItYos+Vg3VqEdxnNsu9ogEW
qe8BtYhAvw+iAZ1jHLgedfClsazVdfPJ1beHHGHifNopbX3tYScQErl2O3uZjZkjVTqU6pRlneRF
nX86Q/w336HBx1Or95g6IRIKt+dnJwc8h5PKrM0EawhZz/Kqekzqo5FVi9Y8pSb3/mgQ+aOr0VKi
JkpvISu8ALt/QdiYAPVXLz48t7RqMu73MWM/CSEqhVDVoXEiYTAtVqD37vQVVOBWJRk3+AcZvepP
B0lLlJ7Zes1La4qBzNVp6uMNez69MpAdhSvGMQw9J+BedNQYKfAHaj8fsh8JICuN06oO6sI1JUwY
+DgC5TM7VZ1/rnYGgKZ0gHfEp9zEyvu4TOIdxeRLct4mZ5FJ50wV6FzQEv8mjB6Q9zODsZDOouSw
0Fn9onmuCfwKvxQKtzHOWpd3gTOABRiTmgyg2EYc70c9rALa+Y7f1HarQ62p+QQin5vq8jxyFjgq
uvTeEeOU0pIOxNETY3QlEZZTj1DOl5G2No7sgsNZgKPa3aS6c9CAzNScSkHQK3L4umoGFgsQMYRW
ldTpYue8xcd3LxH1+Swd2J/XERe0gVB7Ll2AkJV4AxvF5JjPsSmHdvm03PzDmgg0fEHKYsZXky5b
Vf467kFZnEUu5KIaVwrj+JGBvXAqlvzSR3b+5AhHrHMxqOvjeUEAQNOz3M7rBud1YXz51sAA/4Sh
Zqr7ssaTxQ8MBFImI1PvqHm8AQXIJTtvfNFkCDwurHH7Zb812isMWIiM7sqvdDQJCxb9YR6kuulB
HewL4hVWSYEuTesT07AZbBKQQFszH1rireEuC3JYlFLd9qNI2yeA24jsQlfzeckparrxXuktYS2+
Byf8PQqEJescWHlqUfMxglQ7CVi4NktlYkmOhmU1mBA/ojjC6lKSnU2LEaaayYOYdfZqnA9m2wtN
PqFPsWfdpw6l7vGNy1wRnK/z1UNgusYLZfu135H5SK0eSZP8jspwIlxM/ABJhQI/6jzh1Dvbsqf6
5p7UVwL1U8QuTP+rMGXHo5FoO47w4oOzZ92KVmoQMvuU4aQbqfVWU0gnBGKzP3//OmLqzTy/TreR
pZD5Z9IvGvMDGFwG6RELykHoR4MZ+Qd0EEdkPhuBYxwQp95Mlmh0BMkWeBLI+Br0n3THy1RC8rKD
ASIKn4HB+mNjxYcQ3JVZ7P7GTqU6rVt+DqtTYc78braL5rjWqRuI9/onGuPa3hmQmrnJ7Qi1wG0P
LzmD/8Vs22fRHvC8EeDL+QBNmjA/WJVPTBLRFg1fj7p/97Df1M+KppyS+cCBCFqyzPR8hQ26YxOv
feXIXt7ZhVv2kG3ggT/lI7NhVMshDOCTpRrFVkbo2wcPHEczcPjBVR3l4rls4/XSWyKBs5YoXrOI
jImvEJCG26/7o/YObLSw3jB2cWb6IISQMzX3jv4QIdLlliEmZbR4EHBVQFmzFGCQEfH90iLeJ681
fy5h2khSctCfo0T3OezTNosTSp/rq0/sL/aGqaSfxhpg4VHajMKuGMaCekWcRStL2JJ2sPPbtM+V
4WKII7jdISks9SySbw+8USrshepWtmCaFeA3Et9AIZVDMGyYohntrsRqHiSAYV35orWoVeBO8V0F
I+R0BkUru37rnl8HvSWlt3mnS3ooO6xOwrsgyex84LuHe/T+lDI15NNvJx+AZFbPJkUHS1AUeEB5
j8ZmGMtVtooZynOOpF8EoDa1ueZadhvZw2yo3tOPlxI/kIUyn8XVA98tf12z772Ks6PD+nYcjhkl
QOB7D92VL5IS7HcRcJnKmBiBt7CTPnXClV3+KGdY7JioVwpVkYu9WYstEaDbDeMKMJ9peKdfD6VM
AI5wcuj2G+UiNMndao1XveGdDv/akV3nLGTdFyZrIo7IJ0lKn0GaZoV01priWv5Rq+fmmRw8rw05
MlY2/r/YgRglFDAV7BOH76/O/R0RApwaPZa0nvABKlcppEdX/Ea5PPv3KxzPAYu1V+eSBskQDJUv
rLZUS+3iGUiEXy3atblKezuleFjO8ngmBqFOglK6Ex+AfksnQOh3jsN4wb30lYe7ZR1gsAMKLN+U
Kd7uiHtxp3BaVsagG+uStTa0WlZMgfEPTfFntnMyFHz/ctpyD4XJ/CS+IRHBbirn4ZwYnorMFE++
78fjXEmpHmyEjVaYVCh2Xfg9oofLIAjW3/qEHn/dtM3SgQSDnWEallvootZQrp0/tFBnTg/fxlXo
EXUaK9OWiWKh62BUiz2nOU8WDAeR4LUwd1Rvn/gURrrC5o2meT1tP4vost5fpFvtjKO6wzvqq5cc
Z1gFwnYVUwyU4Zx/t3YtOVhm0Ois/W/xXC4zixySsQfn/jqZsSCEn9JWT2nlLOH4VmBJ/cJzXoAa
BD9GaPDSVcFQhW4GzESreSpyCJF9+lgp3PucOqLOyoV/r0sHQXSgI1MxRiQEt+nw3CKn2QHAwbgZ
+2GuwiHEWi/3Ck8X4IL96/ByBfFr5qlWpecmhRHEMnlaMuvhB5qPpRJTrTZIiZDDpqwbKxLelpvC
PhS65S6DpauN/iBDCngrBDIFFKp3BPyvNey+jPyzYefupGlPXaZmTSSyZwiPmT2PO7vp42zGQzDk
FWktKOH7+ZmCQeL/+plmVFB7llRjcyFKmViQ98pLyGttQVpUxtSpJCWnbzAbUxhPsvodEc/P3zfq
jZnKKaE2H4T2kaWTRb7AMXr3iBHIqsiTWCpsEcUS++177uwJacwMt9/ophD6YStKMxcuX9svqHvr
R3tc7BP5YPmxcGgkZbwIl2c575Gib862d/m1mrVI++mzFWZLdMrE8t+Weqw6hbVy5dj/RUdNyXYV
CJt1amHb/DS2FvmFICRtD4nIz29R11C5eTZ3dlzHb/dFewe8YtOt9LOwjafbYv8DBeokZDPVr3ao
lRYg9w/aphOwJdvGoqOwatrdtvsQ9YahAHQxcdFC8ispqU2phgxqYWYPVLpFr/5+V3Y2vNujt82Y
7U42/XUe/1p26dlZggyhleEMDd4aoh8WHDJP5t8V63R6OdeYjzmP21BMULpe3fQ92E1u80AjLQjp
aZw71YAw3DA0E9n+Wz6FRWMoqVPV6s49GvkPr3x+gitDAo3MMXQ6JI2iMnOc5M3vt0bR/Jv5k4lx
+YJ853SUThLoRUcE0qOs8yn4Sjz9Bd7nYwvXLIYjPTNtIHCP6iRIhi8qDdOTO2URBEa0+qOmV+KO
ENXA1gW/OlwsjSWvI5QrJZ5KxyxZqO/Axm4XxeJDq8yt19XYrOFJEPo6GJyhRydn1Ge3gOi9NCCi
4INjcBbO9aakbRGMv274b4E2vUtUSApOqF1U0K2kMybpE4KLRk5h3zNLlDoXpdriRHyCbCxsGAen
5o+fcvV6YvJLTLZCKVMeM8w77X5sMxdmLkrBevUzkMFiW8N8vioPIRqOF0K3WrPZ2CyoSf15U4h5
NNIGZQCm0TZnNsM1zCf9/6yh4LJQQyn8c0m1fRKP7zZeY2Nrbzsf0tlGAyr3eudCNM1rALOD7eNu
9dQhWY/nGQNZr6CRdwov1d2bFARgj3vIuTLyotuZLI9o9490dBx2Q+Aq5Ixtb4FO6kUU0EH4U8Yp
HQII8r2bmPssLbeGsz76Yuafm5NvaNiA19F7XKChT2QKeyJe0mRlGr6THgNSXwofyUfNimCddw7Q
+aNxrxFfQaO0BJbYmNu605lcQuCL/se2brY7pwVnwyjTFkRTIGP4wJtJF695wCVErmbqyGg9jhTK
zt3HOKf38YY2FKmzh0ULhwyaF2iVmvP2zq2DZdCVjnvGNnYsjW3f5AiEOPNqRO2blXFbSXMDMyMD
77bVaabVOhd+OBlWfpVHTR6IP3ZQGh0NNcuJOnf0lvTnNrxxbYeHFGUZWpmJdJsI7r3nR3M63lZJ
z6VLa1Iv7WPSJkF5ZxbY4KpQiQAeh2qvKiBAZ/6wv1KMkiTcW/SNAEsg8VBn3V1cVBOtHgemXEjJ
W8RtXi0RNr1MeskQKpQTxbVk9FM7K/mhLiTgpo7Blj9N/bmxY158IO3bgzj/41uwpKw/9UBvZks0
v0KD77KZXL2DhrQUF36J2aXZRQhzfJG764csqgRCqBwBYeV7calT9emjlILokWs09Qxn8yO0bcfS
GeHBE5PtRIeHQ28JI2VH5EkT9s6aC/0uSx8lKhM/U9T/3r7Hbz3itnO7JHU5GotxUaJDy+pOBbsn
d62kkP+mByaFngZRATOs4N6dg66YyPI43DU4K+Kv0JNgjIpPhtFfJbmvmkwW+RRXF2dlCL5dypb6
eMzxEHFlZGIFWIDjXi3XjlBNk/F4gaUpVM43YdPfgsNN5ETIZBMMtzMKi4lZRcycf8bwYhm6KGFL
UgSq8vvQe6GkHgZ1jUq+bOE/ZfmvHhq+9KDRrDeJl05+0+8dVnEOHRA9BNNSUEg/wvBWgh2MhJcZ
riD57FGBqKUGwx0fL8yuWfgWW4T2dr6DY7298r/y6rWwRFxj+4NcvrYEQQ618z66hFfvb8UT5jn7
TYZ1dHsYBFvv/nFknhZfeq/jAS3rAdBe8LFIF9dLtOufYnvD4eygvw2MhvZMIsyrp6GgkTuN32XW
vBTqbxLtLR2OmBvLKBs9fx+w6t4w8/+soerObIC0CDN33sO9ejv5groZlg714rrFJxPWq2DF1X6V
whFdlD1mxzYiVOw/wmsIkD8iWHc1ciUe61WyVnREbNQPbEhvp9IhnCtTavLEr5n1knSMAPq/bugd
ktZN8eExenE5tSVsF2+PEZSIxKAnnHnk8ebZFh3xbUozYxtqwRmhoK4si2EiiCkUu9X1lCYiSnH4
jOL46t26nWLP3Lbi/a3pzhyqsxWzlvGmpRegGXV/bXVkRIDybARjsiPEXacJN0r05nBWb4vesuh0
rDXN6gtAjYFJZr4MsJaeik0v0d6d26eVrpGHK8D2vXqJgnUOcr2Ge4pQqzxtloKGQ/zHDy6kewyp
gk+WbspUzHDb3fILRtbdmzfjXJepot4uSAIXL7re63Q0wd1bbbLggkmQza3w/ccsKfRX71PiK1SX
rLGLZnnKVQJL16atD7DmVTOmVEElji7vHfduiysbsxAX85oYcGmW9TLe5DE+u5b7xCv2IUH/nRMc
7e0hbeNTUTBj+cBLEdUW41TMUQhKDsvaOVo9fNv3GM6gcqN3di2+PB4IORUqsJta7WYwpetJHc0x
aeRVlGsoGPdHlmoRMZTBNQX3P/OZiGekryUmHeMWLzHdfHuoScQ/NIN4fFUOgQPLdI4nOgWEfc+A
/XFK0x6vP8XvrR+OMrWcylyusQ8ayzFBPesB96IziFaV40BjQ6CXKJlnEojvl/eTFZo3kSIs5PaT
2+2vSIk/ez35JQO+scOjSlWuD5p4zPAbn3DkLqzwT8h9ACKZGq962DcFxhXt3KR7uenPaD/yPF2R
GRj/fuKJxdV89zsParXnhhbDU2tuUSxbtMnd369r1HOiMSzDqyaUh7LELKRncQhoYUEp0YdUkJrl
gFTsTJIw7InZ8P62l2UmGxxgy4mkcWlm7+4agxHtEnmKHa9Spboe5P1R+m9mxbDmm/cQnZWepJSV
tTCW8z1ymwKXpKvSxu9gbNSi3/i+1KIDE1Ll+UaFAvXPmPN/KDNCuihGJkFpBL7y0AsrOZ1g+4yt
vjhoAI2rQ6cGihbhvkrm+YfK1Gi5/PDilFK88k5wSUipzskKBuZJMVRlDGqInLbxBsfjZWBUpMgf
TI0V3rxVoYBFwziayGjeykqcae13BELVEBJVvpp32zZ/A+vhXlATpJTg86sI8sA508kLPL3N096E
5gaBRYdSsDO5YxBNkIacyVk9hizlL0MIRxXUy+YiJ+q9haAKkdzrh26ZCBUMzhZ0Ckaj9HcBlPvv
AeFqdFyz8gpIFq34bfdCKKwgOa6u38sGsW+VP1Ixj/cGtNa7Rqzbs59VEWRew72C3Hh1niR7acoP
Zp6Vw0QPubvDNgP3MLzx18y1zHbfHkD3YNirtWu8WCzryIpNo0AeP56BHho/UYS6VNKwc+LVWPus
uTdYIIx1tp43h6y/8w10GLSDn4ayAc+v7jCkqjQW604ylwpRYKZJCQhLLC+1/CFuFAu9GUqA3/Vh
KFbHUQ+TSiQV2fzx/TBqpf4woXwjC3nOn7WzCH0Y8Oq5KN9xV3XYLH5HBWYaYAuIUb+zlZdfmScl
yygbqJ1fDLht2AL1ssHIsGaFRiE/EXJU3Hz1eTFbpVddivosBSIt/z+1iPdXxzJht94bf0keJTrk
zQXnt7WqW6mhmNH6jhtIzpktX1P1e1MTvH1Zz4krNfpIM4roTPZbxav17qripZL0MtL3oJHqj2o1
71JvVBpJVPW8p+zK1wbP5iVyIe8OS4ydGmwqXGYWQWt2MisP//ttK2UTE6SjEH0691Gjpu5LSLP6
dFW2Mx+GWk50R6014l4E3l48f2ChMtXS1GuP2728R8xZk9LuNe3bxQV+2JU4lv5aC/ukhZZOW6VZ
LQo86OOZKO3q03D98EfcteD+W2Y4taFvWC9b8IjDloFNFOxYa7ChW8L0PcZ099zdre7nGUBTggSk
XldaF6WaOelJ3Rs3mkaBPrrXQUSFPGivMxAOiGE0NsW+IkU82KHfCx643iwvD423iMgcRoZm4TQv
n3I+YlkTIghVMeYmMLOLFdGAULWflUMkTGrgqVuapcPW1MCBPRH1lYvmp0ZupwwvmD5cjlBWmUmS
CJmSO4vRTH3M7FdXdrK5lalf4S8EFHuIPuW5yaz4BR9IO3rruq/9sqvCSr5K1j1TuIrT9Qj7TSUP
Oz1WEfDW+HFBGcgPSkp6Y7VUoPpCvIvKaFnsmk/Cfa5dyl+NU5LYdU3Rh84+XaK681Cda9JF1hHl
yc7obrgWLDRZTswphwBgijfMCa+OZa3/Nb+bigBNC0Yf0Tv/wYLIfeRC6J10ndfvNMFS7rnDa0oH
4wRb6VIOIOM6LHC7vUJ7wm20QK92iG9fSJ7JFUBXrVYIjqTRgJFv54u6/6pMGidT1qmYvuBtXk17
k4nzom22DZNavAMdo1VivECRyTkzGolmkOhpGShcgqhLXJlgLFf/4DEwsH6Lk3fNyYCS1wCQqN66
Sj4qYxh18fXF5/FtyhkMP8ovac2wVEcGd9kUOxZxIhvIP+dqXp5+GH3+9ZX/EJIdsvoOrrZtrPzp
AggGVsuwci6Jr5hHvBqDzcDQdw6T+pT5r3SYYwB8NStE0J2ORXIxRXSJIp9CV9BW71FE8uSMuJOc
KTULnuQk7tkZjaENiGMSoZC2sEbBV1bJwKVByz3383m1GReVhuenvm2YTzQ2v7yNtP5wjtIx/xEM
Yb5H77tIj6W7mn6sS5jnAXZxKChha6yLpinjnSnEmQ0C010qDJeyeeoJTh+1xBd4u7liC0VG//dB
72qgAhSNx7n1zTd4/HVsFD8OktBsXbwtZY2WpuBz/DOTBAsRon0ffbemwiduVXstltUmWVNhCXxM
jOILRhy3gw6gO3rXX/zmyxBCJFvdLlY+XD7t0bamA/tMP6N2iKgMqxHe90NaLeUX05m7GL1EVv09
8tSF9Dng6kjBeDkjLigVYQfdXzfQLbjeuBj7XovHxfzRFl4uwysyVlDjnHAhjI30iZjd/zMRchuU
uBfkqdbRF16SwdmZpVpUZg6RpD+pLXhUogHzvtEnGruEScOLNFUB0kGYFsiXRugvr69e5N1RtByt
JOPZsmNkvFsuxrtR24bHZWWeELUZHP7RbMGr3ZLDQSnAtco96LOnNcAA2xCg27z0572ZqixzrHkw
wvUnAtV5s/D2ZnavJD6GdvCAN+JpyALBwtqi6pOyuZYhZDGP+L15fnASeK3D8iUQ1zavQp+PGNaA
LWP/8f7W2XOjQFgbAFbRakmAKFb7uP2YdUUGL/MHC8NIBdvbPOnCCViQHCljGfLJ2X74U310UCZh
1YwlfV3NIdIprFKcLtYNxqJ5hA+pO+xT5TpW/pnl4uJI4HWRLseoVsp7o13aeJL7p1gc1vOLcnyQ
Vls0QGM1Fb9SJfbrf2ardjBFMQtAN8vVowIM/+0qT1RXuQsiF92oniWYFbAZY+y2sg8pTHf74m+7
v5w/KwbwtMIINTyqetNfIzxHPYHWCnjyCfV4BmePqfZ0NLaNMnU8uu8fTN2E5ep67ofMVhHZ1z+r
qvF0Shk9k+5m1n/5I+AoRjdLMGlWBMJ9lyzHgx6sjarxwhUD/h8w/plOJFALfPXyRdpUeQclKQZ/
Nzn4k229JH08xtkkJHlHpvoN9F9wxYUUNS23+CAuGawmdKMvp01oiZqwp9t71k7ZJwkHrOjg474F
SyU0CXR4cX8jG5LwBqSE6rpmefdpjeOOlNJsFqvwVAOSpVlXfdSeSkdKOcpTkUSHpSQDS8R1xy2Q
G0VzPAu25TFmsTNEGZgk6LpfyYotc5Ss6KaFjxmNJop37p3QbiG5fyjnLT2j8FB5Vobo8mgH4D0y
Qh1FPeA20g6KHAUi3mDyez/zV4oNCc9I4mM+B1QLV74Vzk4TxRuPssCK8+WYXbLa4rSsVKgE2oR5
xvyFu+Z1RM0t0xC0mpdowTN5fgdN4rZM6hpvWjWcsxEgTiEljE/MOv2w3d7bQ/CMpVvFSdNFVH5k
lNYINlTmC7yNh9omRv9dPV3+G5mVUFukyYSxWOoMmiDt5IbsincclzE5xcVZXLBSi4BFUDLN1yxH
hWs5lFf7vS8P/kJ+rY8vaaPjY3axj5XDzPGwBRf8Jdv0/3FhIgOg4mZ20dqFfR1oGEtWaibe5IS4
j8dBgtk+nZx65Lc3wGZkEKsAsRcU0lWIr7krNcw6AqX/8XdWleBRWF9w1GDmXwe2MggJ4/NEisPb
7LQ57oRWVzLQNOeWtB8OhGRfhCzepm1fYvtfY8WlzDUAlhz2D0/JxlLH4yw3jz1Yr9DBlENZtz08
UtPk3nG2c4/iICjqcglb3YY0p7aqHcIcM3h02ZzwDYjsf/je9Yp90jZ6Nsmg9GCk2o52F1dtP+RN
e/E2YezZraFpcFYj7B12CcJZBhDCqd444XxfB+3ZucpSDhjV8+8qsn5j1lsv+9GLEJa54i1aCJ22
Idwp9J+NygQTiewpOpWRs6N9T+hMICA4HZM2/OPVP2A2XlLnwMT/EdOku8VO9UFNea3Wek0gmwyy
sF8txeqUfIt0V6STMKIF7P/q3Zt4yOThjtvKm3AiXRIM5AllUydUYDWLK+61lHM6Ii5uKncT5JD0
zZnpz5Q0GMxZY/k+cpuWsn5BTH3Jo+qy8Y3nNEMv604+t9vKUxZha+xShMTxuA0jXgjklBK2mZT8
k5IAPmyLB/WzEp/VAFdRFydq/MaJ/MdhDC/eQFxWe/X8AGrT1lnwFD57wWnOD5fk3K5dq2Gsdhaj
ORmUPyxRp/jLJLBw/ux/dGGw7EDHiGyxs/hs5fCSJMAVyXo+qUtQEYKhQ2QxLL9gaMnlP97JcJN1
cgD287llDoDHKWdkbM3pTYjj42BsjSvFiJh5ACypJdhbisUZCvnRi0Xopat2BZdaGvu9Dx59/mbK
iyL5yuJWCbwJFY9TXKwjtvxJkpJ4QeJrLkYiDfJv13+bmBZDvx8abPACadXzdJxxWG0OROInoCtH
CfpO2ZfV+QKtPzlu4S/Jfee9CMrwr+MKGV8GIFFyPZnLpLI4Fbyc0YW4AfQZtCbxWC3n0nEmXaHn
+a5aGR10g3qoASvQPdI29yR/GEoJDpOkdi5dz9WRmugmbyV1lhCjOQ0VJLdHY79s/QoeYwocTj43
QsNMTXKvv62l+K+mtkZFcZbdstiopLd7rLlIPClMJJqruM9+VQ1WSZjsss5z2zFIWfTmRBNW//CP
Gv7WYlc9fVYdpYV00dv3RRrjgnUinXl/TRz3Rw40QnGKvNZcEcIl6uac6RXejhM6RiAiH0LgOIV+
wnYN8uRjZQj0j7rduY0IhbexoWPiRjUYPLQUnbM5c99kgYR7Ycnn9ZhKoxkjdhDmWlfWLdCePGfu
Ai4G40RJjjBWA4bSa7r5ItYBXb1jVpD2s/hXY7mxNZ6R9k0lc29cEIi5cxseH4w6dAJlXKtQmzfD
EihinR6xxoEQj1ARmIf7cJwtilDdGFyepwegxCtVbHMnKPUdQ2FS/TDvoNd1ft8haYovXmFEWfVY
hSJU8NP5E8AnfZd6ZjAlw+NxW5PUHfd3eAFr5l2jY1V6s0snI+oq77gQkAjZo06ZpDl51AZYg3Mv
h2mBHtaBrW+LXyPsaY32x0ULMZpMjPqvQIRm+xoVxbebJeHAInXdufTP6+Z4luFudmOFWPtkihzB
szgdAYppJxPD0/CP56lY53zDQidl09Jz5tg7bHc9cp2EPBNKo3jZVg0JcSBF6kKI1XMayvDhrMUZ
oZYinve3/5OdLaXe6mdpUWvOmUXNyROL0ufb2MZj4yCZoUIMR+QLBxC7s5xywc0NrAfsSTMmekwA
XhjZE7tFiUMZLUKclU17ekD80qa0wJ1ANN2RDyahCVFiI9RxRCCeoi9sTacFPcySQDTWjUfCoc7J
kqiRnecC94iEwJO3XVsXRkaQihZl+ZaqG8pLQMDpZU11y9wsV+fXJdKIbLewhq/+rgFOht6IzWuH
gigHKO7Zkyqo/fSgr/nJEwQ7OmfRAiRKNFT19oV6kEVwj2yLBMeEvHKb37BMKXUo4bWNDKdjw68P
m0SZBdB1OWB9YrJW8YT8EWKzm40w1t8MhP0QTI0Budn+pscQ7ujK9/lFx3AtvRiZGQfuHkaU+x+p
iOF0ZX2tC1Wg0gJlgg5yRh5KMrWbMnRNw69rcO5ixsXSLtCYNnLDgaH+PFST96riWOoPutqI0hNJ
Ov+LlFDJ61Eu4t9sPS6VUnB18yB2iicBO/G6EmjfIDxIqWTndkPx4uJkJ+m9Z1Gnaijd4FrvIRe/
jclAhw5IL/3GL4cAgTDC/3SW8Ze+S2UuAN0bcfRVT6d35Ms1QVKkASUHHsGcF6SWtow/iMlmopRo
xEn8TIC+IQ97OmctEVON6bP7TgJegMtZv8AnPxMh06i1ZIm+jo6iZeVoDI1GRTJRFTz4f45x2bIV
akSCpdnU066GX5UiwRXElNmjLrT4bZ/I7TSi5tRr/EirOAPF8ql52X7VWos2XCqDbzVJBh700xA5
cqyAFsBbmzdf8/rqYqWJ85V4Xw7i1YpOlIpYKHO55L8x2HNyDylVQ6tXs7NvrhxybJObd7JB4l35
rjNceiWvUpdWOl4hfjuruJjpHP3kqTnYERp3j88Xm1pFm16PVW4tEZ8NuFW1y/LW6F7TrXXZcYF1
ZZgatagMHJKdv8Wfj8QQWBd7xGAf1DP+EVzzxkZwUBGHVL32kFBxJ/iwowtxqEU5NRnX9NfllTda
OFKsngOqfl4mlhop2JS4Qvl8zcBb7THQEGYXu3XYQsU6kkXir+Vgsj1MYYnIhKO2spT9ex9jidcd
m9g9QOFoLEp3QkIaDbeG3QB1c5c3KMacQwk2TxkayRLyagY2dUtjDvXO2VkQkdWE3JCJ+INnmx4s
JBSuwZ3oJ/uBjB1BwuzsSuzdP+JW4n5yH7w49d75BMzZJ/49zZ4g2/BSmovvv+ZtI3t62fwkpzZI
sqMKz+EQlLtG2pqzGPw93HtPgu3KS388wymF9ShBj3vnzf4sekg1iLiWvwDRHunH7K8UeeQOIYFA
ejLBemVUw6vmjhD+GKR8ADkCNf6MZ6EDNHg3Y1EB11NAiQj33JwAAO+FHMSvmMONEPL6JM+ICsqf
GKYYY61xep8S3CW++dZgZY1hWoYkRlDS5x0zR9ai0QvAgWMK4FlQIUGKaqBd54uUj3CNkKh6HSVX
8+jE0HmgrXFPMcCFYAWJEkpbqEYum4qK6Euy6+qOF8W6gyz0+M++IWJT3qhyvNfUw/SkWW4ZjxrP
hCEQessw01Z0Lc43QjHvUlfc7Olfkt7SiRh7A7RfOh8jd0s07Mt1jjPuTQ4qGGha/utnSNVolkZV
qm3ao9fRsw1WxVy0KUWwNiHI1+ayuURutrsy0UPTcnAkfflCqroXnFCt1Kmwp4eNo8UYwnRfSlAh
WQzPt0+D84AP/1gE765qmdQOVA6pNBf2tXgkDvS6mNcHE8rxqe3IKBOA9Sj4gq8qElVAbUFL3OYp
bg3B9sqVcwNltQhxfH0nniolejN5iAmMRz+JXwuh3yFPMGXKmsFkNUcrrYzOjez2+YyU7Es2wVI1
q5HfD+DB3JUDGEnOT9aU4/3dWgkWTF33n92QgWdmIu1XzScNsems4REQ+3xsR4YxQpComp2Lv5eC
1Ld0ohKfAI87bkCW04/ifklxHL8qEJBbb5QqjupaRdJtJQOJrrzz+2KK7LWmnIafbEHa8NV2/kEC
1bObWMOXQX7m3mZ2ngmxs59l5OvOG/ye8YCXwJ9mDya3I5QkxZf7fd40nJj0PG0w/cbLVYNTzO0k
tFrX+L8ddoP5LF3DuS4jhzaNkpdM+dMNMC/o/CPJhIe9dtQnYPlMISHVwX7pQdkMAbFxLRmnVIkr
eTubnDbh4MYfhlhfViz2etKm/9o/eKJxXDtMzru9B1EI9+nBKtB30T+y3trcQzOcn5uw4kFj6BNa
iMdSgbW/eZl5WUXeqH/Ggj3HWBPn249ylz2yS3aNZJ2l+QIcJWwiOzQJlTDtqdpNZ649HuF7fEJa
CbB8ZfghQOofe5cg2woOZ34kXlHbGFBVjJuFmbpk3Y7/3VXI80qkiA2zIrMHlLpRUWQ3aphJaIwl
9MBfNgweWJPcJNpoBddj0xf3OIBTaowKbBdCeaR34SEWj+NmDQFZ+ZXDXztuqYxdPmE8VWO2lDru
lO5BEBEMAVehfnCrWP7i2sK11MIZEmSqhBjFlaxemTeVobqx1x6ygvgGZQm3XOstvWa5b0VSlhGR
8Z5v5hvaE1/TuVIPCZacavt+vTrDB6rKYEFoXYmmSK0qQNudRdClovlXLhCeQnSpfdg02LLhbP5e
3NLXYf7wS7UQr+yX+h9eT9DOxYc97/Rys9ohWZWMBH+zwwu8GU3aqvYgpZ8CmCZVSoMAEG4vi1/x
5qUPjJHgTUnyk9RnMzE3r/kqKnIZF7ljrfqDZjVc9soR9w5IaHyyl6XzYdDI+yWUROX6vdGLlgOr
QGxw1TJK/QEIVWRb/q3p/xvjUa+bVL7upcgSuIgcJBzH1k/ies7TqESpBHt+IhB13dDb6hWqzl2H
dddGru9dlEpz2z9lbdnRHWCfgJkWYA0lMH1KgeQNsAO7IwmDCAT42ij4kCGUOUrT+ehwCtTtuxkb
ATlkAvOGAwDwR8WN5QoXkK8IUAlat1TYSWFvFs3ByiBXDsXgSpDh5AjE/7vCTwIzfVg8TPtI/iQN
nsFsVCcdecNxFkes9RHL21y4SCzNDoz/z6+tgGLxTTzhJcFHRVoyhUx4rBGe3mbqXqtWGBErGHUb
3JK1vZRXK6fl3knalX4R8XzQvYAyih8nOZqMckFpquWDIzWD4NhZFruH26HetPDdWe7y71TcMWq9
o81X/6ChAz8vpVB9DBARWllTOYKfjUloKJK9OcW60SRBqIuZUrhiD1DgnwYJG6VfYYn54t/cOoCx
pBkbS/zwsngb3QawAqNdwoGuo+ZL+UeC3EI8CB8akDvtaHRFtnJXueqKa0/UZzNUotIUyTcspB1V
Mc4nhdegdcDpvYT7Qw7/5OFiyTnwUVY9+ivg5WuqgiuSwcoP2UMx1xgO5D3Wt6tQzoA4o3evhZV3
qwoN0/3G5iYGBJUw9xo0Gsf8PD27DymW6fTtuAVK/nAIuUOPO60ocOls9n8UrSJWYN0qekIzb7yG
yHoUx3wSI2ga+HDOVt2xREpnLhIz5aL3mXH8noDntYkwnun/B/QlVwcvph+J+KWSB/1oXEtUzEty
I9IokRaQlUkB7SB0TTHHHETMMi/rDTkICyIFOlAloLOfki6iKNUEPEwqt2J5TxrqA0BBCBgVef5l
yCQ9w0/ny/kfwgYIKTBuUVfNHBPIPYJwgVmZVOiuRsa6r8sgLBC0P8vZyMze1MLbO8hsc1oyvaN/
z0WRYubKp5ImkIeudzxYZQHpoYq6XYXAwihharhAv/YDPcjriduWn5dvglC7gBekYVmzow5E73f1
rhECmSe4ktXbC9ROFCQCkwdy2WNLTM8xRgZ+gAmVVuNnupvj7B1C/VC/gBhsSRFzoQepznLiWXAQ
OhHjFY1qYq93SG/89A+O53SStpxvK8pV/Q9f5OuFpb+/WL5s8OziMEWdvB89NC/3m0ExAThAKOhD
YIZHm9slZJwRt4CvpayFJFOJdJIXUaJ0Bup7Dqt30n0hzWIX44b595kRtOvoCmVyWd8JP2H2BMbS
yzBNnrZxx1U4++LBAkCc0Xxwz6MXygE4eB3vLSINZSnTUWN91l+eCywKIme2nGtrkyt7mVF6VdFQ
PYjz6IMl0tyvsdNM5U5snYlA4hpTwMZxkot+0R+4FLcr3kRBWeXhr/ENAr4TmoVqAoKbi1Lok/CU
FbqOKyBVIl82guwjjOWLqkolGT253EHCbftBQ1/Ngfqdr2Vl/QTx1bwWPFmyG3WRaWxw0j+VQFJ/
lYjHfTjoOVBKW4Sz7gcpvC5aNnvsuuK7Yq5wcqFbseHmvT5BDbR17Mg6Df4Ezkl47tjWPN3V5oG0
jEGJ7sdpaNq0TdwLtPd3KtvRatpfBhM0i4qYiPSQlO9jPqYhhFHfEkgq7wuiZmOlvfhVB8QMW/xp
QfY3Ah2Yp1voTZFzRcPeDs2XwMueEeiHXDethQJlcY7bFqRIo9JMotb8WfJbEqf694AFg3iS/Fxg
HiE8hrf+9/+ePrBpGtBv04KSUF3nLNBpXvA5iJ5wrvOM6IyikG8CnRSkMGEZRwyoiW/mqeOm0e+V
8+iYqG4TXQLRnApmYdY/wqdWfpDM1h0MtuOQDjs9N5jzUUKdMBk3Oq6be/w7Y/rC1RgdiSXL+2ll
iGUHk7fsl5omiHA8vvyaMgk//9MhpdROme0/wTJZoA5EeR3PIzWr8PnFka8cKHRRcZDTO2pm/ZA7
PVlLqxRNaPKpzoA7Op7YOKnbsowaV4ILeT/3wJzdPN4fmaNVM4SUuS5hIksoKQTYBA1I6vbDmZFt
2vd708hZcCFo3fuEY4H8T077jqjxl2pU58IqqGVV+0IXePqv5pk291FJRM+SH/gLPheU8YDRtNQ1
WEub1SwWi4RuMAXOta9kmM9QYJt4yzp0uywuCR+9VtR3Bss8vRixE5nfqLc9T556ZUN1Z8VXhEbj
4JfUm98d1EH/CArbLDRVWMIeREj3jmvZPr/tSnjudL48JHMvsnvVqsEf1U4aTWfPPR50jpJU52XD
cC6gmFrk680XuGXoIYpobBj2Py5OyZMdjerNn56NLai4siJ8yyTorNAafDgRdAtyKpIxVT4GQcGr
oIWwJkVEHkfe/3ud7HMhLYcxSiNkatE2Rh7tOTV+p1vupQ+Od5RAZlQuotdYOrKmW4/IRMtha+Jg
XmhrXjj5I6DkqGSz+7wZG/ub8FQiwfk+o25he/tC0iOXFBVYjZ5UUwmzZQMvKxKm/WgL1Vkbgdgm
sNXfyuy9GhX12qk41MWFeHDkTEXa7XRxNvtVb27kIpMLlwWkmviFe6cLVrv1K0i3DHRGl/yI26Vr
e8KmbVJpOb8zFtmVT62M7wG0Q1C50R5Ti+xMVjB/alTbVUBCloAEsPMoJwsPJ9zdRs71dqrjt1op
uj5yOT3gn6jcJCDUM7uuVwjhSz56AXRhEWf67aNIdv7Yap3xtw9lG/mgR9ZIjQ15t2VuGl4sUewq
l/JZHk0ugc/piklxzGuK1iUY03d+EifLqoGhWJJGc7qEePfQQa+ub7sGKpLoPAIn//E0L1A09aWZ
PDYlJ3DCkoM627B01jCmrNTWG8kBrPsDEwTaH3XJe+PrtUDubvsyLI/jviMyo/UCiS8+lfgmgW2l
4Ez3hIR0oxNGi5L2vMHo+D37BgjaHoMbhjpHYV9ks1fTUC4V2kAPMBUVvgygBJibukSqzt/rPqlq
yB9IRfvCSe+bJ29AUa+PFQUSkrsFDpX/RZa5zUnebuCQNFa+IA+4MmXEuFi/bVgch8uePqyvdk7B
4xjW53eaTF3Fv4IE/VEImriy6bCJbPIXuo6tnGEbhEy2WZLE4taG08sA76tFhJqVag2TXgXmfmm6
bcKCYXC/iJRvnQUbhTyWiVYiixgztGqwi8w+ZQo/vlEKb3LPeW1QcpF11Vs60WeCjSQB+p2jdqRc
ZYBlJlZuGtaLWMZrI5mXv66jVjZzxlJxBVrbb60bmv+RhvAvKy5hsPP5t53/x6+8QwaxnkpgYnQg
YQtYhIuXKGjOmcUXFvO0YhiOc/xboGiRn6nlc+4o/69+DeRI0+EuUoj8S0v+9lQRJ3tQOnyXywnv
JThMIrEjHsJvZeL63v6TWCSmylSJDeAs2UFhHOTHvWm0L8XhZ3HqWC2s+6PL2I/OMJeyZIRTMCIl
BlBI/rhfdCCSvxDFd0Yw5AxD/jxvR+8l8yBPUJ1IGLOuP2msYPfukMwEgi3XfPndKLtycVdgZlat
eXqn2Zjo7dGtoVMXe2ugflF9SftMT/rXwrxtzjIuz9tac7GPQZpWZZmuAuMLt3yVC8h1/uvxi9+/
NIjYmyPvgJaDzfrCPydHcAYHI336Q2TDbiezo5QvWQTVKAr9dqrO9RmfIbaVqkquGk2zCwns2r73
+9UvCV4aXBGKXE0P5MQX+dpUAoQniFtb3YmbZcMm4wijwlVb6wKYiJUyqQMf3nITm+6iwEEV1EEj
Eq3Apf/QyuObLNuFo/sSbN+ItvA6ohr0HdW+sQFe5N9CtLNtXsDXo1hxIkCv2Hjo7tAZckUtpxF9
2v4x7Bdtk3XIZV0yW4lvkdQOMmxe/MhyNY0AYhqGeFHiKWhqfvJ5jPi8+UQvK0NqvRay3K2DNtlK
XN64CIfbEJjKz430P/7M/EJdTv349uG57sVA9PHFW1Y5Twr6U+kiiGldn+MouMoZj+D74VasCxQd
xM5qIunqk91U1wg9Xk4Oa/cUf2s8hv5OSQDzzTudaSdY5oie9Wh46s9pPQcIlWj1ZEQUijEHiH4F
ma3tBCVaC5atJ/rqw/yfFBCcHPBlXlxWwy5l2ksKsAdcL8p8hqYB1ziN8S3NIuYiYMkFSm+6IOqS
mcRhLEAylCEdXh19fFM4nMfH3Pv/9xq1i5VbFiHz0zHNzAsRAuK2+maW/QtGCUhS1PB8kpePFYbQ
OvzE47rhOosOhk0FBZEb+DNuIQX+a4t14K3PqmRdUmOSwupyxdSS9c09Q+rm7t/6gFaGyXXiBzcq
RoU6t8i/Hvrp4qp+BCzBrO8GjEy9jB6ty1sCNMKcmnlbMPGlSXCi0jZWqn3TnshwKXDBf3fVP1Ig
AtOd5xdegKZnFdkg+wWArmaSmdRAAacurnA6ZYqnQAhrMRliXw9NdkUlgkBcFCF4kMHxyD3uEANk
FhdI3wr8vZ/i7XLQrdCsJ7lV8B08LfuMmO3xRWki+6X/Aa7MTDF72U2FUXWUm4+TPHqNeK5/ft/p
wumGAg5MWnMXzmclEtKd8WHltMjapR5QqZDz7nrnUzSCVOT6fMFnn2HAPk1SCeQSPHgN+vqdsMKL
/L5R47uVjnA6a6h14xXCYGlZ+flBjbPrNy4NUQdUh98LJCh3bRqTSWWXLhmnZIBvhLk0jGX5hrUk
RZ2xlJHLFWHqm5J5SBzvGYwEbtE8LQuppBViYa1zZnU3xVjTmt1rUZHSvM9/Dh1rBHb9/ikXziH8
GyfxzBlztc7kUN2nUvvz0sOeKXI/xVYIKQUHFJt7gYZGqis/LEOjyGHMNEBWc28z0GMezGrUx9rM
UAMrcUc3hNWQ2PjK2LEN5AMQS9i+/kf51XCXZYBoRXXGKGkKoWL/S53dmwQ8P+AA8XVZ0iPAXQ/U
MZTEfOZ/wdD/1keZMTCcRhWx53NSEoB5NwVv0uOi5w195yyGTLYkf+r5xhI0gb9IJaSH5TIcHqOm
CnFRJlp4MhYcRk0AqXaY7MyAWDszkIs/rZsjlc7a7UwgKHHPIBt1yafRLhPbtenlFeU+W7qe5WG2
6ESc3Gqv9SXZYXgF3eluXjQeXCHkrVzZB/ZLqfzWK73KlI/PjauPQKQl8H1oPk1YKw6D+VaCMBRF
MbfiNTOxitSY7H9QaxaxWBrAqjg5Wuld09Qx8Z/tRK2ysT5zlmpxQ+8fq2hlXLT3krLaxyQKA5u8
zsBLr7b0+OHLmjmOloGY9r5qTJdTIx49budCyZTTC+kcSIDsPRKSWhNjlt/3fb4/+9UeeY4pKq91
Ddun0zVfoCtSHGhBm4yM9gOOc9nB7JvMbSoLye7xogLI2cJt9eSwjj+S0J9QwjQzvETk9xbrQUN/
y+jqI27DkSxMna/qGFAMuXcXu7AECulxphUEa8jU33+t7KTSlK2go1HP0V9ylJmfSYDlRAPeZoVH
AD7sGOPvcGneuvW51d4FFBvCY83opFy06awbYKLxu9avJxVk8JU7Lk1SKtFpnQ+XHIfUm0NBUtUE
GMtpxJaalVGlWgiqrB4GjeYKUzEm0KbYdcctu2OsV2n2dAgY3owUMjhdWiCt0ZQKjy7hjCTKN3JR
PTSVgkyfUoN3Bst0t+U1DYqFVGqRgkvJqKSidy6ZICZQL1pO5LfkkZMjd2Z9fH0KQ8acywvAfsPf
GfvAgHzKMbewibXD6Cmi9QBNABQyVhz8CUHYIHh49aP1GVPthC4QxeTXlxJ50Svdmr1dnG0gjcIq
6enbWcksHXQSMkKHPgkZcYHx2tOfu34zdcyFrwnOPoUPqzyvk0zJlvgDdo7fbbbQDxEdd+VFTW6K
CQaqwJ9esx/5EtUz/bqmOqT+oq1pi2HM3PeCqmchVy1lD6WP9vwEVkA6lFhPxmqKYUZvk2Rszj7d
N4RYpaqpAsqADhzldc8ZzkVKhirfnL7MAX8msR41a82RE3nRFlGOiY8UzfAzi3W3AifVc8vBzUmY
OlvDlbj1WfGLmIYERjEDxzTnVp2oWOUzS6CYi2fLkfUxdMTTVpBh61L0Ie4fku2KK2fq5so5y8+E
vsPh00aWFh/B6G3dbxdbKDDhwa0jrLmN32qCdJG02h0wfWDeR9UKrXE7cdZx6WtgNhVAVqjvOAQW
cTJGQuc7n8a7ZdDdKZOjrUGqCtOLwnvYB33rpy8FjT/Sk4CmyOjFBGVQKN2UMUo3l4xaWYrZ3Bzk
g0v7ReuEOMmRT/LFvl0gZOM+J/P3WtU1s0s5VqOj7WTA+vn4/e4eJwbv+q3m8upBSZcDAQxbzIXO
mY1NVLYh6hLNbSIVXapkdTE6YtzDruOTGTCpLZDqm1xNEOKoVPcWFSwFIE5n7kQoUV1jiW8bQu6w
zVywvwHbZubGMW19R+D/uWZPzf0W7NgdEWOiQtCkSwq1MVHKLbTNfX9rGanrr+yBgUgyawqrqf7u
RigBgpSmfZdZ1lp/o4YF4tC3fb4nLPFuTwP4eIeQYEcO6y0SK/7IO27PVifJvhswkRECvzVcIewG
srFOUOA2Da6nsa+47+C9eYet6d+69fU7hS3rxycduEciyobdpdpd8IMc2W/ApSBU/jTnc0bYQ1ca
chM1oBiWORlF2TVlFPGxlyN6DfOWkV3tWL6m9DQuGb1l+SbtJn87EZxDpFKaSp5kqg0aE1kFKD8v
mEOwQTBSa46+CO8mlTw9xXQv6lkpSHKh9DZ7P+cChF3hXWCE6Pz88CaqSVgPeSxwqMZDUBnqImzX
Y77ht6xjYCi2Jez0e9cJQaPBmZBqSi8dbCtJHcyeapF3PyUunJnSaVn0/FQKfxm8itZx+Mu9fLGz
AIBCYteEz7gXMLUYBmDXIOq+xra8+AkbvaI32+6m+xb/kvZNUttDx4KI8i83OuFjk4GlzRlVikBH
QLlgCeyopt07H1cycl4JkpNOOvdvrH+af2TX/ef++38qnMt+nxgqabZiHY7PWN8El4Mf2koKEZlV
9DU8WfXchaOny2V7Chf42CYylacBYOEtiSb8ymDeqv5Ckt7pzNvDzDD6SWSBAXGRy9inaeZ6Chl+
MlYUBdZioXaWvzOvjvt/305mu6hx72pnsY3K7d/dYD/fh0gK1zmEF52LAEU0VjAnTbVMobLWy2MG
CI7uiJGcyGFV3zRWMnlLl71n3LcR68wCli5ZYLHz8mWNcrvNONoo2I92OAWnwB1sD5Y/JNs/llMi
kafij2wYaqKjNMIy3M+L9PGrmYEa6o6tuib4167/ul7plSL9D1gemz/NSCjAz/6IbaivG/cifq3k
PpNXUvfJuduv/57syrlaJgbnLk29Kf+nnrIMb87TryKMvOxyaRLPyaHVguOT9WEd7XJ8tX7dzG4C
qgbCzlfhaX25LesKPWIGXtmSdwo5tZAy6sNZb+aekpXdUOypWf96tQg1KoypK6CCqrFxSlk9dOOl
8E8ZhIvuWHh5qzuLzqVTLn6yPvZ/wObicQTWz3aKG3/QsK6uStH3bZxKQkluxLx3eXsuLuzwO+g2
Yywu1wG4mMC/ETCUBz4KNKKbQOG+uOpI7hqzVezeOynfoqHvQoQYxxw9IUWw1VN8lJMKKF0iHlxl
Jm7EeNijrM6dk8tF5oTL0DEZvEHXVHxcV77AHrUskDEcEKd0L32LJFqW9ZTzFN0Ccl+mLAhKGPub
/otPMDvwjBq430eLGcuoI+zGbbQNA0THNFP7HDVLt5rZ2CYVqsCZfBa0MZQ7Z+91kysxPWamLXlt
AHSOjG0MV+1sPuj4cwmCr4Mrt/zNyFAYuhVyXUEJ+DnDyC8fzJmEYhtG1rdpDSEHwRD2ajInqSQH
hdpeTql4Sx4IEjm4w7Zc2a8sTueQmcCUsagcDyJtmhGG3+/8TTgpgeWN+YwxeJKGdTyWkGwlV3PN
vYbp7qepqzynaRadDJHKZnRwu7jJ2z4Sw3Uopto+fyxA1Zk1guFADiPfmxwKiO7FGxuzclHieTSY
P7AqHsrVgDWLgK8AttwfUuvnciAmnQCMIT3JHEf9c2mFzkjyT3awGcjZWy96sOLyP22NMQZc7jrf
8UdpiAs9PQaWAInuuIRXm1dR6WL6HHiNl5B0POEEEe7deOmO2/fsSNvo0Ao0UBfL2f9mN5bvGCBP
7dD7CeyzQGhtvq4Mp/c7WjypNiboV2p1aF5yfiNxZJ6dloDzF+TAW5+9kceFuoTySigmSgQK+6np
Td1uQpCZVpaOJ+Qb4MZPBmEdAq+cVPkGfKOG/HdtwLCBVmzTG5icQxxpFo9BMHaxFIlGCW3eEPEL
6Iu8O7onYfTY7y2eVi9e3V+cy3YDU788tRnaTZRXe7o5TS7wtdRfdHXA8hX56eUto0ERCXqFmCw9
xxgES+NUORxM+D844zYmf6CPzV/ZS3NiForkzc1jLzMnAHtYW2/aUmT8eC4WS6oIKxvZ6RVS9SOD
eT6XS31M0rYMx2S23EVUH9B0A8B1hz7+05kIq78eAr2eL4YWUx2kiO5VTpbeU3TH3mBn/4ywtKjo
LXEHLGyy9PgSOPz0ZT7Y+RDd76iX7arPHOY/7d8fiJdXOYmFJS5aQGgT2UqN+85Mgw+qQa2gedxU
yT0iHg3STXvFx3tGpBN7gWUhDo3dzx/YYRKUzd543txGbvnS7F2D1r9+P1YZbV8U6Jc3npymNFWE
oFOLwAt9f2R/7T48BDeSeefCUqUZIWD4xtgsG2mmeBodqyMSdnK254ZAX6OKxfvd+tk67hjTwch7
5+GEnSWIRrYAGtYlRXTmE6PwckIBJ7pdVe9L3zzxIZl5cWNKQIXAa7lNYt5gu6TddyCDpoYXzFxs
9vpe2BEjNXkABbLu4YIcoUM0eF5/whdBFM6A74Tugne2mcRlfsCVcGZG1+KbIRrkU9nhrmv8zQwz
sLEzQjq8oVq8Fvbcm8vDVs5/yz/W9mIqAsKofzFcrFUtcvdxWW2aUQwx9yjhbtvnpaVuwHb7+t2/
e1zDEM2TcmRM42E907xyXKtEPtTqyslf0zvQdTOMvt4MZjAPDUfR1nH7EULRroYizlAbSia/2zgM
BEDuBYlK49v2VTOLLd8x3T2r88PiSjI7YK0yAGrYdnWGd0mjyKVRLoTrMWQE2SFHDBj9QEsZXVsI
xImbhFBatXVq5fJhAM4wxuT7P478cYFn+iOSEOJKr6waje1u4Xkl3XBiTsgK2K5UQrPr6KGAZqte
yR6H7TV7w8QEowKn4KG7KDcp/Scue7jH8el0n8UZYSramnfPmhmRd0maXbF1f37LVtztSrixfbDr
SxKHwBje6dyNbIsq5QHqtOopj0645CNmTFSSnoE5OBnTvJYq7I/suDwwldirx8mtahlfmCtqGGJu
L6qFInnCqz12guxJhAcdVVhaLJlfdeBDiclrIQ7+12nF4Z0rwmRsLWHLBDGYdyp/9fLNn4KJ23q1
2FL7lOl2oRVLEFTtG47rmms05Okyj2b0a2xwtkRYt/RODYPZ96SrMARYeCZJsqlgMgUKIFqg4+Os
TYivT41+QGK7YR87t/jBS+k6nxZx9bIY+RnNij3dxbBd6Lw/YjaNOcXWbhsWDkGAAfRB1ld/roZD
ZW628BS8wUUuCLbJ2Rp6iZ25p7OzNuiJva/9EogEerEF+VbMbqn6/GC3VqgFF0dH50rSoNOzAYIO
xr5skd/H+9Os5WSVhE5Jk7wfa6LIYxxytd/d3tvSHMAB4P0hAD1tAZPKQ+UJrGRro0+glHjFIkN0
OXb8oy36wbm6gqWVfXziFJQFLKsa1Yc/e20r2akeWrW90q+TtrmaawOjtN7xeWNt2HWghhr+Xk82
xPqiqa28RO47AcJ84t/NkcrqbQDqudHkyWATJRjh82KxqTlOJjrAdXSjCHAZnoQxWHmlIcEHmFB5
co+AypkFPAvN1bLZ9QWWIc+9MKFfd9G4wNnY2i3JUFacb0+Ne+7tKGpca12zQ4ZxaGgUUaE3N0q8
atuur5QyziVBI/jrMtmMDT2QyT4CATCpGqdGCloKhIMo9DBjHl6+NLhnwbAY/FqpZkvMTmp5lifN
8mcWX+DzdO7rhpl2BKMgGivGz8G7wF79ycQV+yl67nAkrEyEYtfD/J0SaO0vVMvESzM0vhTLRi1d
tGCVbxWwtbwQPhic59YkCmDyAz1fL8vSYBv28GRx5tCYIC9G85cdxUbN34Rj/C8LNF7CzPwLE+57
kRnomoGN3tbDe1uW/3oZYC7k2qsiVKVlgNoAewRWIrxAoQKq8vHSfKfKy1MNeFodc7mDTeVWKlvm
FY3F+5FIfvsKTVSDROyNVu3dLtVIwVxlJFfXDs/zSiO7Ql8wWowvcPFDTvtaj3B3suwgP4Nupgh3
7iSAYnDxorNlxEYdtfwgIap8HgCiLcHDdfSbUkucF0Y35F17ykwa4WH7u+sLwKe1Lc/xLYp6supX
A7PiUdDId+ZQre22VJteN2fI5UyuGEGE8NsnEO+fQ036FeUfvVDbNLeogeKtco6qaoMtSmcAgX02
DVNcmjvQ/Lj9Wqm5oeQm7pRsnRu5x0uX1zI1KBcq/fDbCBO3d/FLHaTtIrkGhZOY+GAcBanVhYkY
9t0CTeKB1WmhF0y3BIJBAztimz2oLpj0X66S08QG0E7UbJrx40nucDKlfr0NGnL+JKrS6NwXTADr
S8RksM1ZeRFqUyTYh4NmP/7RYQH4jScP/LW6vGbypQOCTEX2adywPgs0uoipRiB45Ejludq78FiB
phy8qA+wstGEamEjQ2MPKZPh4zzSuLmxNWf23t+iHo8Erz9D6L5JqXNBqVL4X2cyJXstZaSpuYTc
Kww75S5/YaQ+PKCotUgTr4lIRbQHHJPxl92q3udMK3ScnwcH61uEuykL98W03wo0CVWwOJfdKH0+
+OYIIURW5HWkx+gCarJnL4C49ZI+wixK0OuxG1rmi3bjRTUz1OdOcd4AH+tdVnu0Evh3lAiraaPi
PYhshfIHeEw6siZCzyHb419DltiDtY34zfMP3DbrN9kYUKxvQ1e8WzbCZoB74mfLL3yGBXMZLYlD
fqC7jMcb3dH81G2l9qVOyVp2Q1IJnTPuV/3DbtSO3BuFXI4tDaUmDZyt6gMs/ZCFvyvSJkqsoqM/
n7CS2Qas/hseF+a0Q/kIV5htBNXYr1MXwHjn1Y32W1huoylGWg9CzDqeCpyHS9aNDDYfnFF1PXxE
eNMj219VdxnZUv/YnpWgiZba3erKR7ZeRmBdojqDbYfmTJ/8KC4xQid4vKi7HuAbrh4aM5S5FX7l
VoXXkZdZktuyS3FdaoTDlHLfSse8K8Flm7DACKeVz01H4Z7Wt1nq8Yw/qQG0yqLrgAUHnXyKLFKQ
eA8V3GDN6qxIuI7FkpAn0POB6SHbMw0tV0pthPpJI01QaHjGFFcANpQhiQ3APoqhsnyH4dJ/CYGG
A7xFUYitS4eWohS2ObUntsi6YFFomlYJMK5XwakgJkUAQzZe0IpCT3WElYrvxcOo9Qn39hNZeXVt
Jy+PUk+202tTCPB1zpxypVClhAjHyNM+ql3OusT/Amo1KBgJEi6wDAKsNad71m+tKYKoYA0lCQIZ
awT3PE74Ck/eoCqOY2+G/1FQIvQXSbyqALfT6ccO7OjxOrlRHug7PVEvs0cHDJ43sfFGbTbIZzNw
N2kLE8iEzPW2bSFyPn+cVx3AXuTSObaRm0VWYZZWsQ/nzUwsGa4lXGHkBmqkQm9U961EwSh+zoLD
PBcngQAEMtrWsbF7fIyxYUoOU9vmIJE3Ag9HvIscklV5Iu0cjc+hLqcOw6w2hnfFKOU/lujFHGTd
yHBZS7RTS2icxirVArrjYagYbXuBJivOcJvOtlXtNB+sEH5L1KXttnkMqecjP9ytP6vmzf5ZVn62
R1rlJ0vWUW46v4zcCHGyDPditmLgaVtwAtYfL6tWCx6DYoUEtPnn7imgraBp7OIpKwgXxJak2CGg
Qk2qG7l85xh11eabq4584zcIPo0DO2plqWdA98wIKav18sdNR3r3IMdtR7Pafmn9rY6ESPb+YBRS
7eZfTD5mIHxZGOAZFwdzyS/AVseQ18f67+bkceQ6PvnmzNWtCXcLtMGGH0cPIveGGbrmad61lAB6
kwDSuGScgYgyiXIiNmDqGbITfv3agdrqt5h0jGdfVO0hq2CYTcLAk3je+IiCWa8ctP6LZuPs95YP
D+hVuwFpbFCjb9CosPEMCTaubqzdGVL4PO1TIjRxSf1Idc/zeSDgiSyS8O5hhhkmPl50eT+G9Yrh
PPs+231z1K1O0KWr3lwW6BmG+ZsyF5z8E8AxzyWmShyrqZixqqrimA4G77ACMu7gxInA4PkVt2uz
o0f5OU2+Iyoq7KX69kTj7jJZO0TWL47BaTvkWdSlhPnBaTDgSlxwknXxZ1xV8aHO6wZXTgXXsX3t
5gi/eVRpJd9c4CQwBhj3wLijIKhjZBW56eogNtw1NzxAVeLp8Odrt5FQBMl3p6ne0MJiWCksaRJB
Zoh3PJnoON/QWp7/hTrtipi27aOgmoIaIU+SQBS2wctc6sr3MdX5tUS1DznvNw92Qx/xoXqeHcTl
zxhNi54Xo83s3v2JcPb7nVjeQfKTjwkUTsBbM81Q/3OIPPhv71yALNoHO2/8kXrwKq+t+pcPWwJH
coQ9WacFTXbSqZ2iw8nI/QqO6rcm0MG9SDUfT3741Eaj5V8H4xnvnCMol33NW5xb7U2SULLEUZgS
V43l8xZ6UQjaW+mf/DbJBU+Hg6bKY3dXLc+WFUpCOGSEbasZ/9sdZDe4AhuISCTB8dSKsbhh7wUV
qzb/lbv6xCa2DTNxtD/1gflqB+Ir8Ah2QO23V1rfFneTci69GdJEBVhg4L+7KwVae1vzK9G4NomK
rEexZmUwoKSUp60YxS1OtOzfgBIHrGN8kaAtUkJLeB4ZKE1TAOgqx9m2lUOinRyRLSyr3PMeLaaN
7bxUi0onNOpEh0J5cN0ffOD50S3L3HUJHPjBA97vr49xDe3tbacMKqt7eEgGfCPTYxTmaffOyCqv
zuccjCybioYJ+DkrKJexwgSkSA1PSqysqNc7lsQ0nVokGSbFFwwf1+TqVzfRHJBFy4NeFgMTyBMz
5YjLoIB/Kxa0B12rq2ykbk0BmfaFaT1mnTdSkoU6Ca/tw0ETT29BCv5hibhHoyMQ33Rr8uNL7H32
gDVOPiUgmMdverP+tFxReqgBoFl2BHUKmlgiascb3DeEZf8wYYkgpdQXj7qnNvrUq6mE9sooRdUO
7A5BpFOwn/O408GT39Q3hoLpAlnDAomAR4SkYc4K85KTjYd4QZ501D6s97m6alZQpAvMdQnPaEgc
fn5kmTksd4vjkTdgNvuRURKjO6zR+nPcxJajXXYpK8/XQVV4W92emwYU0wCrydDvSGnp/ZOfw1l6
CWE0lBV7HxfygQs++3ZvkPs/WiUHUoin4NcCITqiQPscmhIIur/4WjwK2v8re2YKjppK/5tesLZm
9iF9d4ultELZArBmVoNuK56Z3AvlqRcxPViJeIGJ1LkR2XdlhnJZri8/+SaZVcnmXonlLXvXjp0L
+6U236/XoLS5fDHe672mLJ3CBMm6c8Fl5wvznLxOjjZ/XtT3zC7ayPb5+Ic2/LFc3VwFti34P0pK
UXmZ3HZ4ty9+psNTPp+pq0s5H9n/1hMW4Yayd3OxkC0ZtPJJxbZQS4G/NZk64p7Zc/T9AoxgtPC9
R1Q615Opnb5TPXnpHK28kZjHGD8TCfIvr9Qh2z+oZjKfxH4w+6gHBY9rJn/acanCtxQ+xcoZg1Bq
Ib5ePdiRsxPwnvSbRtmGD4Z9zSR+oqzc/ljSXA6NzYmp3sWu6n2LPpdkl8qV86xQiRxWbFoRZfl/
QIgnPKIc0XeNnDicLKOFvDraN21oz/MX+0KwOmh2LJGmfdWoD+1FwceYK0788xdmQ/MxjQVTM3jA
J8aFLBWes5lFK39Af6dyDo1AI4bU4F+Zjy7tOJBQ4pXZh3GVngTtNiIgn2qNxIDy0gCXuETRm5eV
IL1CKzXCuV3PHgvB1Vg3huYnje6mSCeOVvHD9aInTRhGOY8+uCd4zwHzQKPh5wWnDAOdcJ2u9xvy
EXcZ8zP47uFtbkgpi9m+KzVevbS3fuLhm3WlF6YFnStL07OSdXEEtbymTMOGFXBmhjimjp8/Cxy7
mT+69a3me0+eB3uufRLVspLRiioHk2CYLbjgc5XsgE4cc3YcdBu63BWJrrCTOzk2ymPUTWHdbZgQ
QSwz4SAJIlwK+XaA4x7ubL0XYCvks4TwDkBYFHeLAybRtyPQIl/oxESs3TYVUpkJZyfMKdxK5j65
apCs01srIgCQL62MnS505dG8Yl9ei6TSqxshTChaTYYfn8FaahH2N/uq2G4IuwLLb8fP0Hu9IVUm
niaTHAjH/D1Y1clCLdC9qdXO4HrPGQpxG0u2VaVOJpMwycjaUUMOtv9FQMyl6UrQHn9U693FVR//
OfRAwyfT25X9F9d5e8PnkR+qQMJiAZ2QpwY0wyYvCqSvnn+tkb9acbP1Nz1sIrs1iB6nNMeUpKGA
5JGmaf6mNXQ76ylIQDnajPPMm9465NLo4q/h38JVBz+bX+X02nK050G53/dcV0C0RUvunhEuiXyv
V9DzxvRwNlzIPrZuwoZH+7RMsLJ9p5AguxZ0QjQakh8D9kaOuRXpFoIMJB5TH2lumkWv1WeZTQuE
lS/fUlgD5TS10dcxcyHpR0DZsPzjz8FAQGoCvggpbh2E7GwqegwgCKwEZ0VL6eMbQmrJHgfU+/GS
rLt8Qi5WVm+C1ml1PAIGdO+Gic4m1f4mU+WrxpzxikNbF9pD5ltOZ4vdK9nSk8iPhDABh1UHLyfK
WGiaSc73/CR0WG9OUzO8gZAbGtYiF+RU6rki5IFH9+omqWwQ320dJrPX655LpW8U6IKQUkO4ajIw
dhdoPAw9VEzwHEx9JKINHEqM6jU48b+WSma8bgZDP1TjBMAsZA+4sKZuL2W+B+Af7KjXCRJch43z
fEaPByMrzYJ0hg/+4Te7wawQMapudPvP3lGSEPj+MeHgCTg6wGlHoTyjOe4+EZzM/nEnx7D/TQpg
XghbQwyGPBa846nv1yBGKTZlvoMeLAYIsj484S57Q7TEsr5PI9VZiA6CiKv2qxJabeP9ZR7sCtXL
iE7IDzEDHWucimUWNywa/c46ZkHEooiauOM+tHBJZnwgr8eeVXSxBp4NgaIavKaYLsoKxQEK9Xny
8gGJoKR837/yIE53WvfD67Z1SU1MlUaa5rUYJRP28g4B4BjNs7NeVIMQsrFo2zqLVY7MgC6QljJj
z28NO5hQxcaZG6DpCpwOc0WwscSEhDS6aAKoCSMQsi//pgsIT9BgjUXGMdN+5qQ6I7u3ghCF+mkN
9djn42PAZlcesN4LrC0p4w1v5g2UWezA5BlDpAtf3Y02DxLX/AirPxJfYO6qKynuRpYJg8WVuEmW
Q//0EvfCiV0N2BDze7p5TgrX7fcxmC4Er9PUMYJMbxAjCFtqMAG4ALUp76g7G7rqx79eLGdtu/OD
ov6sCCfF/zyW4GdrRWdB3vWK5qoWbSgVGX+hwJOyb+J2/Ug+0zDI7mMEdCN3o7f8pGx6705qldoF
lv0xkXqwqpgigILEZWw4DOpJUG6/2+9T8t2RWbhAebAJljXEFkGeKlt76pwEpcl1nPtNQNV4aIGi
Zk2kI1p9NzEsBvSqMtBzDN/paVdtPxcmEb3L0D8IlP+5em1oXdcXSgl/Zh2JTrU4xy3IuVyLlbL0
YF3KN/1IzHHFaRIZ7IaLUPKY7RyoBiaihkoo/SOhBVPtxK5gbAAuiuUMAVTMdloTXRPrRnRWkb8O
JOgUwPVFefPFCb65QJspn6SrajEdC/NsmbMwAH4phQdbW0t0nZA57JVSlIEtnlieBpKjbX2q5Ihx
+of4rsZ2d2NyEn+XaW6M+2ZoZ7V23XRFx1aBW6/Zw40Fq2RgLCD/88tByYmjRkRKCub0PSN2TOKS
40TA2THgnqIJmaSRwtf/iS7RDUrEec4mZguHeGDhAjQVvVA//cnF3efXbtt85Nr9EZ8+e89Bf9cK
ccxbzet6/G1U6g0Y9Jnok+tUQQV+ULA3fcsUgWMIWADK9buwlwMPlaHZv4osCKasp+HgGaa3Lbfc
47sD3VDLuTGV+rqa4AKDvwFp6tHlLIJESqCA4zUIfb/QedlPVEfg/qPv034CJ43759tiu9wpA2G1
3ywvto6rvQ8V45WPotPOgutPO/olAZW4U71iolRT6C9eVTME2BeSCz5cmwCt3hZBxccAj8VHK41R
bfOIcEYKd7r1ayRNQ8K7wp1NlD5d4EDei4ydKtLwpxPpNfyD5+yMEUITIm5uwSp8DhdoCsPyq4Df
KDP/Lx8F023Y8ovUe5YDwfVv8Zh/X16FDP9kjYOFA5NEQDE2QBy8Qt+ifcm5vme4qGoI0xJuJNZm
gLM2JKEBnYCwbBzgv/tSkYP78Eaao+ZYzztwdQkMUbNtobyEepX+w4QcUuhjUMqrLuLNPL/RwoeN
c9wEytXnwMpZuEonlMNTSF5CdA82isv3JScEtPmBcp33MCznW/8opZlKxh5g9NyuXtQy8m7W8iOI
KPCGtBRQKFdP3STN4xYrbNDtQMRFYUSMB2ZCJ0kno7/xJjATd/CF9IuILLca5ZVet0kQ+Wfbm2OT
uuWdGmzg9Y+Xp4bdAm6hZ3zpZ+zKiBFnaXNfFKkmTW426VsMavXsjXcpfirr878GgW+fqwhbrUjr
/SE1Q0yyQ13pvrlwhgG5sJWz7GzpWh1+ZdyFHGgaRVhcJwZ9Erxh/s3jplUkJ9NazDS/eF9xrcxx
ZwXjRFlEdQGNYOMdje+Ej17i5z5ROYRVl4e5JgA2ezlon/hIDK2byV9ogilsGVsZY5BqZpFP1EhO
Gzt9Dq8He+L8gnPO0KRismURD4MlL6TaVFBXDQlRpbRFDXZVgbrf3+0oYDzx88m5ay0iCslkATG8
G2DzoKGKjp9hnAPLIfoP+WjnyDfXAq6/A8JQ/yY+pRVPzHNIHTpEoTm302ZVBX+zmVq3FsUO5AjA
XBILtOkJB9sW9AB5/W5z5MtBtR9STL13ge06PVA+TCIoALu0Y6VMjJV3RHkfnexv2rbL7ThTsWtY
HJp9rc8D09WjysXvrMoiJSCpTOIQbxYXmLjht5blG0qG+qkBfmz5NCf+yq3x8NkgJPtnVsNErygs
k+DYKMW5K3m+xse9a/1DyXRhbG72OhByWBo5/CjKZxbmwGWkoD6pbcnDVZabaRX73Dgv1yKtsDUy
e+XdjYaMlXfh3Bdg6RNZZEdq5NQCBA/o8HAes6a8ZArHwn7LJaDkx/LgftJoQUal93XdybQJHhQv
kAsmpGAGpjJOiqfU+lqETreKyhCTD9kPqg2QtDnsFiptQHAIdmJ1SPG1Go9IsWXwxZ1GLWatMquO
bNYm1wXraOe48duH1AWihPe9AO3bQ/y1TwFEtc06oHUsSxDP5K9DvETWefgjrYqT78v/yHMH0rib
1Y/w6blNhOjs11WJUs7xAuDhe+wLUo4H7aoQZAN78gwXokQ1XR2qRR4BM/aJPL/MpClEJzdsIEAs
UW3b3xfch9RzS562OhqhAi88GxoWv13+WDdVdQR7GJghqOpS//wExi/8Rf3x8lEgP0XceZbfAqQ5
C/mJ+SAs6TpyAgiFPDMhtmpHZUQCxUvJ9Ews95spzMnh7zF4erESV38RauVG7JR6qeJ/gkocpfaQ
ClNv3lmkmOB8uCfXYOJFuFZvgoW272/3R4mAl008/iFnDWiA6EWkwiQ5fAw3hINwFYkTRKegIlKo
YgCP+VKggLYEiDsd9h6HMAT1spnViZeVkJjVm+Ll4T8vVOHzaR2lDppOY/3CfDi+ed0zEQZpI1vJ
K3AKj4FSfMLC9/h20C15Mwq41SrNuTbPm94z3BnxlKHGK8nybsMHXsz6Gns4U1KPB66NJndw23oV
IhI3f70LoEIP0OkLJ3S994FhEL7WaPjnitPAEXIjiSKXSOKsxoBhprTDDXOHPe646aIBTwlMZNMI
c4i3zRTSrhTeOszuwNafbHFLWYFcPZPpfLONZIlQaTUmhOeS7TQ0Zht1t3w3tqtVGp+CXV0WgJ9+
s7rCkitunTRLWosBgoQFj8GZtG3j5PbH8zanNusdWPdK1wwn4Ah5aKaZPIPzzXTlwMxtX6uTtQrp
m/lJyyD1ScTRzXButK39dubNCWul2t7eW+fINA67ppiJArGhv/eQigRmSxuwDHIKK+MGty0OjZIM
SgPVGrtVp7lRdJz3ZTB6I9sDsK8PLXKmzCzcXuzvGDopjtpLBubNfzs9ILAuOdd2zTQW1JDRAjsh
tFybf8WmNiaNCQZ6tW5EYmgRhTc8OddV6yEbmLCQ8miQnktfKh+ZeiRpQYioBzsNwITdIMwlo+5T
O89wa/robblJENc48sEUQXPmfAXNp5Jpveeg5LbNwDijPVya8Vi4yS4AKqnIDdG/DEYzwnpviops
DGSNhnePbE4LFExqeDk54p6h+BXhJGOBwKNkkv3mQ/eEvvaNg29Na/PCrj5L08sc2oTXCMMTzXZX
Ijewth9RAxmbzEpcKilueJII3Z5ySLpT7y9gw7fxk0W8ZWVWCNLiSuj3lVubCF5/PaaKwKMIy0un
WL65jnH6DoZbprzFOBNwOrVreSPIwpstQ6GKnX0d6ke4RXAihG+ZcC52vLS/0wZ9GX4Mlmv3bsW4
cEByjQ7iu0rkmSjNYliS3Y4tlYM+teX2tfJkdBf9FNWziVeo3XjMs78dHnK+NtCs34Yw00OnUvOF
wmfxipRA4Ge/93wr+WWeNGSHoxyyDvDizdziEFAX8ZQeT9Bws/tPuxp9e/dsX5Bepea9LoLXkPSt
T+5c4LVPdhCySU0Wi3ukh/y+VLA6jQSR+CFZks05ADG9LutqajOLuRmLxhaTIaUbR6nC2DCrBBo7
/mTIPHMk+ocOdpDSIt5loq/AB+ExA1Jc7CEFD+ky6KBgIx+NGHbJYegPOUdGN/VQZhjVQkn0Ll9K
ARiPDOo4VA6da3SB696TwoFwYQjx5Yafc9a3h7onKs7jSh0N81y51Wa55Lm9PRHF9d5FiUmYJq4j
Bf8+s5VsdepZLkwoGqJJ2vaYIgLpalgXKD4W/B6aAUL/+hbhjosuDhGEGZLMEVa/kHsLn2OsRo32
mZ+JL7j8o05YngaoFWB1cccrpisjwF3PlzFJOJxaeex7jBNslKissDj3IPx0bvo3H3DtG0tWJJjl
9f6p0aOXVBtOf0VjbJBpYxkBRuw6Q5IYw1qaVGs+F6FAQsQbkRg6jjhH8GeOP0ayNt/CIGseNuHp
91JtEz/dEZnCDMMFWN2I8kGiK0u22jdfSLOr8l3XC4MPxdoURtzhCLnJWpJ0zp55NB2sw4BNSZHl
N5OFJMmLb4NDoA7GTuEiUV4Oi2B9u48DzBjaKRzC7rbANjahnCcJd5WgCu3PHIQNGLgkeywMUlNi
fE0RdeL3kbpsgE83sCorO/1dX0Tb4FqGW7S51Q9uY2iZj3jd4drtPI0mzPGqiMXq9metxEm5ea85
LYZDzE3BNWPvJg9ItogV4TItuohajVip2um+Pn76yAFPdbF2X/tDdada3MAtxr+w3z6c9FA0a8EI
dt2CVaWT3XDeYgiE18d+iLLsC0Bm8zNsxRecOpYk8h0j4TdIuwsE1yvNaymQOmIPNJOaF3/ZfIP3
cORDbA/G68iHTxQc1H1FFJqIdTyZwUxnYvWCY0r+Aygm/lzB3/2zp6O1aB6VIc42aY1nDIoyVJV0
9HWRUueBXLsdoOrtS7/s80oC4MmoWuZhnFM9OroqoSEbLPaXPorRtM1nRmb6PCOtI61BYRgPM/yR
15TkOWhG3VjMj5Fjt7TnWcCNzKl8m4ACtURDAawcf8OVCXpJcXWnHcUHTvYqYvACBr1kj/HCxuqb
Ne3rD5aLq+09gjFyN6rD2rWvttz4hxxjcuowbmIV/g1MWTHy2MLaNF25492G6D4d4JFAl8zrNJg8
5/Xyv8uvr3cis7v6B3/GTFf7ACzWKjamK2M3OiRyhP7431JZ7oejzxiZNH8ypNSiBzn4i6lPsuZ5
Xj6C+PppGAbrUtvZ889q6nnJmJkFlwvEG0Jo7DNdUKZANC7LeTWYGY4m9sl+7OsB6v85T/NIsDrZ
XeQZztT03TPXOAsCxCFxMbshKOKYpbL9LSvjyBxSVWunkxnP9H8C9i0kbRauEwlL5dOrdAvS7tnw
3/atDREKyB8HmMJ/RGoawdxawZlstq6xy+3vjzkgkZOZMCSi09D+pU/nCF/qwuTgTJCpfYCOjcex
CSO4DwyCVdF/RO5j8X/vMN8+QrCrz5anP2PbsFVx1IYQJXQYsGk4lxTzB0NtKXfYPZfU/exmWfym
RoNACvaQBx2/qr6USie8zBWWnkpckdQElVMLB2oZOnVkXVjmzze9I2l/QE6RkQvItuObY9igltbX
SOZpdgC2fFa/FiMxdiEkvbQWlPGas2dYbRVoRJbcQaZu8Tjhez1n6ty1YpQpJGA7eaIzT9DMyXam
prwDJtc0RMTfqKjHWxP7fDnau/bvdT83gWEoC1jMUg43/JZz1GUusalVAIL8VL/ianWVCaJhRLCJ
KWrpsjTte14IqcTF5Q4AsQkleJe+F93xiZ/wAIeDImNyNd3LB4j8J+nPTnTPTD+KGPMe+9LD02XG
s2XYLfdbqLrnaxBiIgf5MvLI040m/Xm84ox1Y9bLuoO5oSqrOJGLyRnqdsP4dErrK0hBBCP3kr/v
jOROUQXQ/uHxQKNbqo9HWbUepfJS4qDrBdttkW6Lc0YJwDJubcTBDFl8FFnX4QkfWf2SstU32MP+
3G4fQvLMebZIz5C5J53V7J5BuCiWxsaKI3Wr88K7Le+KOM7OWq6jLyrrlPzPCLY4wJNMPKXSdffy
0eT96r/CFWB/haXb1HyUJvrQlASMMsVGKlKkJdmKlXR1sxlmWKpCYs6Jauoj/W9ob6QUOh8TgB/N
Gdr+cYlD+LxiScUGSzlMMDtvtsVGF4/UH3yAHIBwkVd+yx1gdDqcB3JgSnRCPT2MtcgHe/5RGm4B
8IFx6R6z8d5tJH6AZMByqfuxChzOdNUkxhR+RsU05AZOjm/u5jdpwykRiWhOuUxeCFoqXb0ZL0fz
Xhil4pTVVPM4HwP77iKl+Qa5u5dtuojBtaO9o+BDhiRUtmzINLcEIx9Am+hkYmi6qwOCZTcrebfc
QhqVL5H7vo0mtPxq3F3rQlQtJYvhwaUuFOp25rK/XL+/vuiAwo7EAOSBNj5PIgmkswdJ4x/HYpIl
rtmrb+iaOaJShElWOuzTYMgm6os6KXwXUHg3gXJT/hgd25+aCKogcMsHrsez5RGjRJ7TmEb+y6vw
1r62bcsLBNWv/ZCn2R32DRWOLgCdQTsbdPFEPij7ElRMCjUhIpaxJ1ZxRg3kWUJtp7c/sAb+9WQe
+QoWeKgSgmzaCZCJzvIpWhlkGdAKz4lbPbR3tnkSqsgQGeSQzEOsQf6N0JPKoXc/nEtondXXA5gz
OwfX1MIA72HtabzF8sjw1ovYxxTdJPmB7q+g1OKVB+Ovbt4A2/f1+/NZEvnfi3jEP2FqtT14tARR
lhlvUphRKQnff1PHrv5taXauPmIunMWqeXSWZHiNoVDFO1Ls+qi2OMFRjKVETh+hySJxH1NckXji
0k5XIMTL05mEaBysK9McFy62DzqGK6ym5uf7VQ+TgOMXMNuMgzPfc9iuqgdGuWVOd+ci4lJRBoYM
54sZuNLE49ms13qow5O+w3n6vYE7J7sImTU3LLBsxL3Ricow6vRXcnMm7sCIZ3Pe0/qBtPWKeenn
BzGRDzF4ODLjCy+lbCQiV4sE7VEBA+kCjVnyd/mdLTlN0sGTH4p7qykXK9NR5nInICEbwqqJ0Tgd
wg/kvyqYXpKSXUShHlyCxI2VENgMKIjF+QL7+GdmYReHeROz9pdclxuEj5tg7BtiPbXTMk0i6Gfu
OEfF0c73iEsuGZSwEiQbZmrE3wTuytZqkB5hK4GT56oidW37r3LyCiXCZZIHAxt8fj5IVt+FT52X
i7wFtlZl0vUfYNLx5P7uDxGdLQbEPkF87fdmZnPYh82dLV/POU6xHC7guOd8rjXVDnM1OaDRazrP
m0FcDnMfypEWMp5LFJIA7vTbqsEVjtxzWVggHxfO24ozU1Fm17upLYcXW7CYZvQBDUwZW9hPcXW4
Y5CEtWuUmOGVYJcKVJJYtdw5motFNunOH9RX6KvMxShMdetYnozjWGaJTucczk1kjMTLg+3cmrle
+Mcynx+IX15uIYu0LnCMTdFC+K2440DivZRpbcK9Idn6Q88KAf39DMJtnOSAwwuAgTsFQfXbMMFm
uG5pZwOkKu9HPp/64ZfmWwcRbyyl69pFgIbbXNleIL3R7oSpASFCBSy/muyIwjUzh5TMDDG4o67t
u+AX4AFaNEf6QtwDrFh1h9fMZXgMtkcntlIJIcpYbgdPxjLIBB2DzErErNeNktMiqblAUwS3f0O0
tg1nJCXtfegCI6ALjZka0gJ3MS+7ZfTdwj+uqTcIgRObkCvOn97iYw8KXoW3cop6D9g48blZxw5z
B4SnxjK4QZjHpmgtuB3dP6ARtZqT27DAOptSZgYAMGLTP8WLBdZvo9ThFTqR7cVg/+/RZxoVU4Vh
Nr0tJ8U/J9MKtMwbCPSBcFcIIsOPBqHNW2aKOvUfry4JsTQKptvMYbCA1sJ5PEQRLK0kjIaHqA4r
t0O+fB0hXel/sWrmSIawku9HSTX+p2EVns/NNlH4W0YKc5KyJ3uvjaKHJ2j4hgLJeUbI5Gp57BWb
PeMIWiYAVLEhkvMSA7vOw++8ZasuMN+AvjVCnEyMBulVrH1TzJonDzJeG/VmjhZfGZtUnciZGdYv
n3czof+yl6o8/DchPxBphqaEoidh6Zsc1XZtLg+5mlUcMHnfsohcQsyeibVb0klTLnhm1TEY/FRx
hquPkMxe1ea1YtYKcKyLpLkyGrhfVanIV3OmlOVqwMSH79azFZ9VFxtK70s1odqRt6GYV3bBVybw
312IYk65L3OKMWih8zhKKIi3szxR/IiQ5xU1dsK26Uc9xmea0+p3S6O0Yt0I3MxlsrpDBTxf1hsZ
hALbK5+h/nLcXFUuJ1Bx/NFdOdB2hzgF2S02BnXrThrl4SsuSYV/HUqgRnwCDYXbs1KC3wWRgLU/
pPfNrrW794NgEH36t+DhWmi/5uX3niSYEGfWyifseuYDsn095SyUyGTb3GTJTJMxLi3JcJHSUxj5
BrElWJfNBLPLeSw4Xrc+62Q1lfHTMdgRrTaZ+S2S6Bw+NbS02QXMPkiZrFbtqrsWxcuj7Riy0EEr
Nx2NPXPM5iU6YhRbcyXj+VGhsGRSgC6mG91Qba7kiNKEPFdokhqmOsesyD/oNE+YjIhWOxY+kJ0Y
BRMlod2R8GfB94UpfIFXTxsInfcDYODRCJhgWq+QUbp15HRVbj7XW1kynPEz+W5LngXM1AnOKVN5
jT/GIWuqjSAsjDij/EMftLJ6nZFo0kn+LPlIvZ+yjHxDG9R4wbQxFRfMb5JZ6CyEQE2rJeu5Tpg+
6sBfTkqqvXZtxNaGEx2mA6iuZaPCujqa1HTCqls68aU1n6cdVrady4mWpGgKHYNTSlnsyMQ9Sf2G
cEdORRyg4ay6L+WGmv/xUPNOlIazd4/NRbZ3BBNlJ2TMQCDYX+eZTykd3px4Kr2cavVNoF+hU9an
3h5jluCmNuVHtRDbWzVUMqQKaxPb0h+NZg0x4cLVebGd55tgIYFiRFpEYyy0qs2y7A424c8cuTAF
Ow4R0yBnUu5zADofWH4b+m+gXJ8Y4enLuh5OsW4Noq4LbpnGv73P84voH1yP/2z8MnVMAnF0MVTk
cPiCJHtuWEdFf4Gh2m4ZoMCqPQAQajJHVO5Y3sGWViFNbk5MbafkDuOVOiDLrEPqfOEc/5gB3YHr
5zzTiPAgV7VmsohOwsRXxwC7N3Hn7YgUgzPg7NR7t8CegVPdhJVI9mDJtnKY7QJLYZMrYZ28KmqT
yx36rcqzHgDYaVUdZZylxMBeAyDwLvROSgRb20ZR9ckzl0h8YJLfuqo3EpQhKxSwwZ1LEKGDBTCW
tTsxxN+i7rMCUQTIwduangTo21un4w66xnAyIsxE+0NV1HfoL3SL4D2lyfB/LTnQBqXPmBOg5kRp
1a+7gPMsM/QAg4pC45YqWB/rXk9YieaiydGHQ79XPYfP+KYrxindz0u2OtezdP+Gmq+6SG1yGVeO
Zr7jd1zDLfwpV3uJBG878fSOCcRyWhI1jDOm9XwxP5TXI6sBiLZAxmI+3/YtgvksiZoTFtmWn+6S
uRFL1FbdKnMK0luYnMT4WjkRrfV1f3eovYQB/Gaf39ybVK0ZS79EV/H3cHJ0tI4Mg1v0IKgfMGKo
YNMelddNbDVfomxS+uwAtbKQbJxa0DqR3WFZt2WHFl8dztYe1bSgfEi4k/7d9QiCqI+bxcr4IyEf
jVtiAePcKDH2sKYn7op+1eYmc6axoJQCjtTqgO9hYQmmFiEhdmp80XjUg4py6C82OOC3KT+OOhdb
muXdgiNTg+2xZcah3/6qzVdXb+qda0AW2ZLuUCPCCA8DeSgP0sQcg/pHVORZsmXjZJ3sGpPp0TYB
IdzHy50MzmeL9AGkjuhRG8qh3SCcULt6f71fj9IzkOG0WW0S1wCor/aDq3jwbZapMnV/wE+x1Z06
ggL1jkRiMtBTlpVg5Ckd5hAPyc7kSmuFRq/COuLNbY69YeQPhY4bFZLn8gWG+R73Z0MyoJHF85xV
R+PBei9S05Mz3qkNbO3PV+TmpjUCCJgLO8dtgN7SmdutCPDn/qv3aZWlFfjMdBRz5ILjEjHFZNy/
3yQtt4b7IMq7u0uk+8bkImdiAJREerRzFjkqy72uIl8YdggLrLcK2x2LsBEbfWPv739DAiEwnaLw
hJ3T/6nRL3Y1OGfNfQQnSIebMJW/T5UE4ZgGZdotzlMbgqbBm/5oHn1sJzuxBdDD46vn+QD4udyI
oc+g9WxZ0yikNyPG9eMlvx1Hsf0EiqdXvjTM2oyzuMtvAcneb0FeXQNsiwN5ZYA6SsGPHkxVK4gc
h2qQKZJKaFk3htQapFcHlAoo7G3u7g4oDiwRd9M25X1KsnJBign507HL7efqk5B901B51gPUo6oz
sSBj4yB0MzYjVvlNrYsJHMyfecB+PhMiHS+S01sxKmUmSP0ZuHWcX1v44NqqHwYx0E5onsEwyVVy
qZsmAWww+whFUmPJuPWlT7+I9nePUuzcTtQiyg9LpR11e8iGPOWK1m0nAi1rFLYS7L8I0jbDgOVC
f/CKrUr3dccaFXc8ZoPDwjY5UJvF6RI9VDkvmUQ96Y8+gMtQXXALEgYuKOgaTtzh4FX1CNuLd+c+
J/eaaRE54qQhhXVpSkeWyiy+shFEEyMHQJ+IxG5dsTu3kiYX9JmsH13+FWnmrrUi4ioHBKkZIN4p
+S4VsTIFqz/fQKjvwHOfLCVv8GcBVmR8bAsGaa1yMORRv2hLlnO3xHvp36Ho/0cq4gLaQbF9qgxU
JrGV5rayDZCisKkejRWGsqF/1UAVpkuCLaxW/QHMG6A0BNh5mLbuY+Q2RCTN+qbru9FbLj9TM+x1
LJAau5Y6AU1W9V6S8Nza+BPrAbpUR9XsFtF27GfWR8ShmXDt1XT0zhhoJ7uMpKbzPHGEFc6nZDo8
9di72j6q8jKj3RI0wNI14IdKPlzz4LKFcNFPe+4z0VOFNnPqyHKNofUXwkJZBojhbpeYuXlPGk3O
zpGzJxNS8ANGNsDOD8okqkQ2dmh6eGWeF6hUWlH/wgebw+wQjLr8x8nPL/6BuTOLlKztTrplWoEZ
pmQn8fgdDH8TcKxMzl6LjRv6QaOGpO5H4jEUF4pOasES1l5Y5Pyx9eT4MQEswvoiqdqNv+mmh13D
1aIbRpzgKQkIvBbUpHGToK1//o+hxZ5xhFGouM0Phtnkim4dm0jtw2ADcXi2a/6M0iTHsXywiYtu
3MjpFfA5i8/g4yJZOjv9WQYKBayVj71CB1AR5YT5etjQbjFgFU353KBGmTIBkfCqgpoj2jwcuYl4
9duaPUNBsprKNLnnIzIaGTNEtM6eFEmegjV1wIOO9irmdAQoZYYNuej5xqq1kwIoCsVb23J8qB9n
y6z2R/2WLeWNQvIA6Tero2w1rdpLzDKsw7p3cAMNSAqkFG4GGj0mYRsTkiU7KmOpDjvndPqhgjdn
ZtnA/ywbSeunmIgSZZoMhsqYYWdmRVYQCN70ajnOSkgAQiI73lTNwlKH5N+cu1hXnteq4K4iu5tG
CCQsCE5EsE0qwVpFKvP03LSmKlXkeaXQYTKhTRvSmSYPN2pIqDyptH7PAxR04wDJf8kvc2N03WzK
TBr7/aYDw9HNfZt7QDSxK4ajHrQ7rYXMr1eQpc7HXO8LIdrFTHu0x+snmz/k43rzuOLTkNKOqhZC
Kv4uidO7IbEyzQHNA4/NOVYRxR5TPE6HeALCZSwFPgOZEtVS8AQMVTewN3l4nE+MuA4uPaxT+YhF
r0GBOKvfOpacceghLOYKNwWQH+HE5HHfIrihwcVLexo95geuqCiNWzq5SvNCbr4BAlOC0TejUsoo
8MYAljWH8iEJDXGpPJmEGTETM49w1u8ui42BUuWPhmRaKqfz0u/ego7bF1wk6rufyvfR4Nao7Tyl
E/mWEUZ+Dn6VJ1Qj+nqdYsoA/cERqYuC1A9q1ocKJHUeTtmDnmzOolfSJHmVU62Sv/ygQetrfW/O
CwxhxTzg0F7WlEZYbdfFrr4MuFfymqheGWj05qgE0h6+w7ybi5S0cVkagBL42oZX+scSxKYX7QGm
5VeA/BSLyhW3ebPUHlmalOdJRDLN4KEGGEVcXwh5lrrnH1EkQjmruygPDk6y582OaZEyeIurGLUg
IP6ntI81Mwn/O7uPlAARmuBM/pKVcVe5lhXqvfcZZ8t7e7iP3PaQ5Q4TAPTB0sgQRHWbDROBhUcP
9JKToiqV810+4HVWOrxhcFu+1ORg/V/zGHfQLdHntRDRZVWQwoqp3r/wZd8V8H06Fzz/A++5OugO
77qeBoKGUHfU1LkdNRxKSOfu4Jq+YEJEw8xHQH11EjG5sMTF79/f+uIh+KzfFPCvFfmEvt13DpLR
zcrV6EVgpJFkBskqRLZ5OCnhxvXMQdRgsA0PP0m8nEjY57IJ2vvSfRNeP7urdpqy28riUdVgC6ON
rx9E09RimfymBy2rHzuuBipxVP98jY942noosLOCrImGT/+yhunALFrH+GXZ3OhO2RTVLTImswoh
wXm7pxwmPk6NKtq7n7oZ8B0LDMUmzymDCVAgxZiAnnSFhqGCeSzvVLGO/NgIPr4QaIW78oNOGvK8
YhDXiuDnbx8+YEYltPUX2yI/EUrDrxUzMH5PSkicP9lrm+ijbUmlDqCACRwqzL1Z9hBNIl3XnK6k
lwb1O8QPZciO/K7I4uzrUELxDWrbIDzZlg0QDLVtY5NYrCYaNzxY9B+DeOcmRgttWdc4yPnXBD+7
L0OlApMsVLjIvyziVyMynT4hjQpzPFHVH3NVEiBYRoG/LbeWpmAf8uVU484fvtmrMfnFGJKpBLO+
brgCwAOiJAr57+t/fIYDw3coDeHfsTvvXjIchKxKEM0LUU6zQCg9W/aZq/sh3y8RUqAoimYg9cSw
pyfk9JPMRgtcQ31382MFLiQaa9vDQg0t8L8M+vZdVuRWuLEZBfS1BgT2uaQtSZ7q/LJm2Z0Yee6A
lIJkpQCAtz0rZJh+t87BU7awDfPsxP1X5on013DFxQXYTW1vJHCfxBDJJ00Bnohh+XiefTYFW+3d
pNqXta56Mhuxtc2q9vYrqx7ERED/JLnS2OZG9cK1QHkfNGwhYZ9V8B5gv5GitQcMTOAhOrozhckt
kHJprivnVQrDmQwcPP4u4WraCrsSUVnmM73N/IQzIsET4hJYzoZWCXaLKlL29QXZdqpc/LW9zWrZ
CpWkEPtsv+KTmmkHW43JYnfY1UKUs7m9ddo1PlEfhBG1hlZQTMUK0UbHa2kksxCtm9j7qQKi1AyY
mr7nSaodNlfZahMr3tv54QB0fUtaBCEx2UKV8XTnwYtXbAGzCZGpcjTeFFQcpEy5IDHZvbFtqqfI
5oY2T89ybpjUsYJx0EQtGweywh4LUQUbxlYIS6UU5ThsjWQvQsNo9sxl7jnE4/Y7xzSe6M0KsA1s
eI2cGCSpRlX66PoUNgZ9UDY+k2IhRZHHq89EL11r6mRniWzPYd0tAgoTP3g37AICBeTUmCHeFI/3
pBXElwjrZHJ3XLYno5WcY0qtvKPMVN5a/0/P+eLBqbIqFvfIiLgW/kh/Da5kdDD6mgWBEyOSyfB8
0vupjJT8xSLcY9yK28br8AiiX+WtgkYJ5m0rFXjXqfZjufk9mIZz41mFGdRHb9+Js5UhmUjazK6C
Sm52YiixX3KPJB/v4oQ744tii9u45WpBDbQ6LwIo8PKZRzxydvoKTAp76fIUWRno8Gqt4bzNZOJc
ddrmGlWHq05N1rGFHCyyxKvouH6x1U4o+QQQG+9YPbvlPKDuojrrMD6s1W5cs8CUDEGNGHI1O/2B
CxsqbQtIP0WZLfYm+BdwDOMCdZp5VlmJ9FuXAcX/A4shlUJ708fSxEEytLrL1mtu82dhF9LNY2Yy
xDcFEMFlECPgN2poMz6K12taAELs6QKnCni6yAGO81152lQA6yj/w4HQfCHyNDo0tAcZ8X3RjwUh
cPV4/Yw76IC/oVi15JkFzx1950V+6Nqwy9QHOOuUgFzk+07ScZ3t60smYKQgmJpOCdA4Jvw5LNac
VlsUfRavqehZoNiRj/b98Wmtcv8gKIkzXNzsb2kSPP961lXt94OjzqXr5R8xcNRXEhJykLn7Y/f+
sIisrEUj5Vci/J333N948bh48GY2tuNY9e1k3BTWSh2JvCBh3h5amjzhknf2RnQvPa3/lUNKvDNA
KzNxfeP7QovHVMtujc3N67jvj+WzAmSy5Lw2J3bBDg5l3iXlBJAeLAdFnNV5t0NThUEjJ0L6ou7B
iYIg6T0tY332s1j2WPay0gYDgfA6DzzISoIrOCWW8CecAKDKl1lJeXXbPbEGJf51ZQoI7D0LQ0XR
e/QwyQ3DbZS5sYR5oAEtXaqGo8t07hCi2FidzleOM6wUSAbcByVhQIckqL+G1PKjnr61/GIabdL5
IvFJub7UPB9QBF8Ot/8EbZoiLbCMwseD8ZTTr9tN8AzR8q3cTM6m6qS545YK8bR4mXL4QHrVn8B/
hAFIeRmP85iiDrJMSJkdpB7tyiqY3jUnCXhdRyJnZNbK3DqWBxqrT7F1+3/lfTmA69YNG7T6n7Eq
IvU+/JP1sfHEoTzXxmoJVQftWitvtrY6MOcHjR0eJsOA6SyfWALLLKWpg/CoGys6sHXBnRwtCW6/
DRjI/aRyPjC4znce5rmZ+r6e3z1NRflUsvWIdGRwtioPsJwYunXYEnrt7G/si1KYCxBdW0sjud4m
RMJmeNFvL1arLwaMo2HWwHWq1RCEjOCX7wfmuYGGb6Td9vDSC7mA9CsenCJDlFYGUW9OPMI22VxX
CQJhJVdopPpYsVIbjHjwvCQ10g/rKyGik3RfiMrbCRAJC1lLuFEOEP+uKJHG68jHn563/v2mPJ7O
WjxMZUV7JAUSLxs0ubY+vBHObcQRiLopfGiUssok6qE0o7DwG6zTY7DMPInkYeGUNySDZn1J3aXD
CPbXOHLy+Hv42Vm+61VnKdDlfQHYSDISn5tkidfnWG/n1VtGY84VqQa9ga/S+CqhXT0C0TO4cYSK
6jjsR8vU2tDH06EbKX3wbWAlcLFxUqYXjWoB1eQYPeqEBUAj6xnW0SGR8cNQQq94td5GK2qxZY7e
nmcI1ig+wWDPdzVrvIGDiU72sEdbhdwnM1I+vEcc8CV+I9ogbmdFMUnqRDd4EbcObmlq3D+W04Xs
8DofU0LRZdrr4ZruZzS1NMuaRW8n7wkOXu91ilqe8s7dd1u8f0NOKr1F9Lm5/FRTiY0ifYd+bcY5
k81tYriaIR0XWLuFwCX4hDFseeLeZiz856hC65R6/IbVN4QCw9hR+dvtOlrhx45VyiU5IBNAF0cz
UiUfse4+hUg9htEOopODnpgNnhgkq1STPCxbAy5+cQzLbitriESjzuvPSXvYTBkWYy/a1D3zKqKo
zxpfQvxxVX1yjLeR1JYOKiMpRBqPYvc0WFZ7eaNBLXe6v5olH8rJb4q5Be5MblExXBfbju8x/hYF
Mv2voc73MC+ezqdwBvwCA7EEB1Gky5zHg8bCwReHSZRZSKeCRHa/yUm5FbBtwXTcQjXbvkhKIDma
awCsbzwF9x2VBS+eatZioxmLZg6N7M+aITU0vKXpN2suhKKZS/maTqRah1IH9nlbi97bFUorqXPk
NylHDOmc9oRhmqiczcLjiIl5CHLPR6CejIoGqgAr3Ai+d7lYZ8s2JNhkKpS3Oa2ZAjKcavGfFa4j
+WNKhYI8AR9LxH8t7/9Ju8xSvZxj0Ck8b5RDYPsUqCfGd2ku3nbz60bsMv9dAEM4+d6Bm/axvrx2
et1SdWbT1wkpy0ULCpMWRxHcL4im5dLeWKS41Y7Ta2ZZ6FbfSUnwUOkkcTT70/iqS+8EUZvYoZqX
qbdLooWYmx0b+mcUE5J33804sdyxat+2X9YuseAOGTsbOEJ9abFccJKvG5JcGteFTaDnQ7DjpLbw
LTLaapnlyNIdSP/Go2c6KUyLtziwRbquAM0p16drcc1opSj8MwaiaIkvNFTEOyQj7t5dzieWCXze
9rynx3adGR3SYZSZXylmeedb/muZyBrcRXO2gIS3OLiN5e4wOvMdQhL2S5mfTINWuw6CFVxKh6bi
hNLHP/5KyYYKIZe4iD8v2G1NvQ+nLsKcbzavX8sppbwXsTZ4WdR3mUZG+hOe0M3d+y9NBi8SWBM7
bZzcvGy7EgJCT5f6J+C2IX5u1hgFhHDLRnHUOhJTg1W0eNcpQgvGrLsxv3kCDmuQ4W9y7Qzi5Yjy
EKv0J0bEWSMmygnPZ97LJgmLnD8MEfySDZehG2hVMZaHVCScukJLZrjY01amQ5omXWTZ//OOgVFu
eXVFkUMbFRk2y4NG+ML1D8MfkGvuPlXR3qpXlnutaJfFtWhSYmDpPGsYaO7moWudhcUU101O0uTq
PZmEHj7TF5rFJQLSNX3wbG1sq4zxHtUgSiMkbi3M70Wj7iPGRhyfFqkkqB6eBDpfu84/pI5T9O+n
IFUeMmNrZYRYYI+/6ptPqPG6/69Rpo3lB/nTauf33Z5F0jP8ztJtitvY7VbbNbNDbciWH4xx3pBF
cc9/2el7mygTic0PJ+QfON+qZ8CZqWb2zT6R8WKg+KzMahKyXaZvvR9fwohaDG6gDe5rz2wuyPSk
NSGTGROyLoXTIQ7dftwIV0RoHuq5U3/r9MF6cv1q3NqRvTqb387i/GzN4q8FwnJT9ZHKxr6YU1jS
I1c1DT8s9977iDXyRWpsbWiQIxhCj7C/0c3FDD8WHrNrXmPlhUfcY0Q+Wm0X22QEFOrUMHXtAoA5
jaK2BPzl/AeDpvN7m2Q/bIGeyPETI0DVGIpl0JCHiOYU74jXe1aY4GiHK8TnVYuhB1BQTGNvtOJC
MPnE/laSqOWmdwblOvJBi3QmDuTE+dHoUMRkwAFli9Hhkj8jE3myOR6P1nkKrhuFdUG4B72VB2MY
re7J2rYTxYLPs3nDBGlzq1y5Kp+p5fSkNTZqoNWILMtwfS9BfpfFqmorlrSJw/GjjqFfwpg0I96w
Er6/WdR2KnJhGOEFhP19cSLKVe/emuJtu8z/4W7usRra2EqJq7k2IR7Q021V2YXjKTw1K0TOn2Fj
qtrkUbb+tvf6uqJRrh5O7duNDyqipNmftA+7fPLu419qsFssWxUTN316xm4CXfM5VhkkJ0eMNaae
ClywKdvX9mRThhddPU2D84c64Fu/CBX8Ie7SFn6fFyxZg6MiOkdc5f4nvjgJCuZyl3BMVZL1SYC7
XlsVTNf0nv/WdmgctQ2541VVscPHvM3DY1fmEfMpWc2yxlV/gXE8/PWlLAVyyi21loRn/oJwAJWB
pLrsrEnu5fQlVxN0WjkzEDwGYIFcNFHWmanfdNNDIXDkR/jVSNLh0jwqQKVb5mqNNPqup3VYrL3z
ECQ8TkqeqW8FOVsEUSdIMIxmwdPFC2h2TrQaIEFs3fUJHyupnfgBqBA0bc32Dp+A0RouGk8xbuXr
JlU/C60d4uhTcOZOJs37NO5sftnORByjUBfCkqDyx/s1TzMxaIR7qRAJOQzl6heuLGgjUrr43lRn
iLapKAXs6g8xhoCI06udCpk0pIgZ4tPNujTEowO5WInAux+FtjBiCm+qDKflidMBe3Yl/cq4egPN
BslJdquz7aDAXeOFlCnTiTLLzN0UUUxKS03tWfdZrXAV3bN5xT6vi2b1m5LW3TLCtG7u8ia/pEEB
4wMUqT/IQURgb/I+nLvDh2QlsyiJft9vmv3PHTErBPJFOTepq//X6zNMocMJew+97/5vHSX5dlDD
saU/ZX9ermSg4TFmO3ASKYzqBLv0F4SxTxmy5JsptskBm1ZFZs2zyO6trQXg5JvPjcwRfXYdVq0o
XrnotC19CawLzCByFZOw2rbM7muWSXqFouU7fV5T6zLVlzIhRp/DEUf2l/mzYlGF3In0K5wkRJqO
HOLQZzbvnuxow2YLTUoFEO7TUdxWSCsIiOxrrGdO10rCcl6qXiBgMgiy/2TvEadQ9of0w9xU6jcN
1yx+f1h7/wFyYArVS+PKHbKi8A1ISoh9byPL84S1JI1nY+RIkaavLzZoCyk3J7fG1sDzuu4RDrmW
YjFf2Tl+TNY5GfvvWRqDylp0ofNr/bdEITSI0pOJTePwQZStXAHZcocwYZPLZ4k8tkSkWVZy5/z0
8c+gi61jgYja8fYjHeNh+DQKZGEGbbkNMSYN8qngNMOCRsuYbWI3T4HenIbMZQbx/2swIsRhiWub
lWpvCOGclk2+zezlCB90R8tQa5CzbCV+gvq/gjzXv/jCT7c1XZbz8VND5gRL77k0m8nUamlAa8Ih
RB5T6Zt+HXU5dd/1osjO7Pe32kUQExXyYf6jfwbyJkbIRmLDo8itNLlHRAC6UNhj8Nu4NwBbJrRa
Y+ILsNsXgAd21OoVRAU4u6b4GXkPsJ4NHSM2hKr+/u5Gybr2M+YvGbSny2wmX58Ig5WzdM/TOUiN
E1uDURSGAAbE2zwIwdumJ89TZiHS3oIJcGrkc+8g1KnZEOWMwq28RYXaYgG3Mdjz3meBHdpPZ6FP
J0QkIBOIgWCvq5RDDbBl/tQ1GkrR6Atk9N1we4eKI50M/Lrh+rzixs7lfd/yZbUal8AZ8ZlzR096
qxDHoN4L1ElVB2O9Kev8k5yiZwyMwKb09cVLi/j9YNf7S6c+3mXjZ0F3B+I1pn7vqN47J7kA7vwu
mfZU+9Cd7aGpSFDRv4ofTCQB6R7YnEtfRN3XuINTLsVaoNrF2GiAwYgwdCZS6p5lCTm3CiE3HGOo
NCtYtMll0pyUqDQepSuTgnwdY18duiyJ9oEc5tcTeVDrAmjFzfMIboIDKKxFxVuocpy+7bXcEwpE
xnVomKGGAFIXn0JwkLfQ9yBZlZe/fsp8cRF9EK/cveUSVLMkyR7JGL88lxtimcoGjkOTuKQptRep
5nB+kDftzlAK+5epcdT+3PtQWiFzdVHj3pKNzYY18+EEz7RBgXCC4XaAr8bOcCof4023cMCN5VCo
5sCwxeHDyXTLTuvDvT7lQxY7F4sD2OW4UBg5wKbUhPJLBz8rkzanIZnJF5EJZ+tYy37c4RJgJMC6
7pbGXM36zwv6SmDFrCysP/JzEJvDqLoKXeruzxmug8Fb8F0QQyjtU661/hdjkEtgSySJFO8q8BBD
3O3pT2RdgDfN7G2/ZSfHI87ZVpaAlM1A0KQ4dExZljuLQ7qZr9WBn9NN1ZbXCY/ZfGiLYoW1lIPg
wLafkGC8KdqKFwvm1sDwhytIwHsk/AS5wynxhcMcg97fc7zEQmviJ+zhQkiSOvab+qGctNwmaKOo
wSpQ1nEJp+EahDIKcEXYKiytRUjZSv8V7dgpgVyUZTRv0CNRmhNbm+iwfLTWhTQBY72YI2I62+xY
8pQtyrGeinSj8Go7Wplt2dvWaXDc4NkPjx74qzgzzTYzkUbMJS4pP6bYydeehU5u5iib9719UJR3
qZhzUWuxEPv74f1kqUMNLHrMxSJumezLfF2UE50qGCt8lswPa4f9O11c43B/d365syFuG7OyL61l
C/LtW4A1Hkr/vXo32PqkKqZAfvfanxGSRgtLiJavMZg74nAF7kFBAIsu4uj3zkvDoxXuqWZBRbHQ
vj8V4ZQm+NquJ+GrD1jBf6Ys3nPuqMI/JbEtLgT4wse3mGj3AdpssrdcDURGIuLTnblHCG2RvKe2
wNhwIb2Wre0/8G6n14MZz6SdZ6dTCvK2gra2d48YdCouq8Iu/eGO8iiszD1QXybmAxGaUWS5Vz2+
8aEIyroWkbY4ioxEjwK7GzOtHfuuYLn/3AuIFd6wyNRO6s3OoFCXIUAOUFCA8Zw28wO+NO0QsLdi
pLBb4CvVgYe2jY6GGndtIKrcR+SHDie36S8nCQchndbHuNotSf2a3JMlrNO7fXUOQ4hfdFhreIGq
LW0JKkTgzw5GsEqsbpDz44z2gXDRv+61U27hMJ6zSkrxpDYj6VofHGoQev76Kyf36Lwj6+VNbO/T
4FvRRsgymmz9KxPrLGT73ZA/rwOCsGkvLPq2/vo7o7fokyVb4TwHccdCPu6cZ7lblIIURkPz0TNm
eIYw8bqFKc52bWDSq+XR5TS2RXHBmHDoo0yZJ4UIbN7R9r/Cmtuse1MS937Ettjej9iJK8+HpzEP
AIQ1ypUC2zYy+8IbCf66zv9LcDB9qQilaJAGmHfAJNN4s38UwCcytekz95f36hHWACUnVayCE54y
gUsaT6y1lWy90HbiR8la6oEKD+T9jSSXKCYKRlmXZfp9W4hnL3N5AEazsuixKmYEBPb+l0d6iAAK
vrOyCps2usytEwzQIr1d84MTpV+9i60sqGsnNp+Vrt8CJH+P3tkOH6o/QcMej32Dh/7YMZ9BOyjQ
xLwcOr/+lrQLhUeKl+3rs8fdwzHrAJdExPwVNF7FBlFOyOT7ndeY9KR1H/cJtUd3fkdO0yZKKPSH
bmpgWV8mYDKylwe+STHsYg/Xf23S598usjc5qKOOkfsYJnDmRrGe++WsxIJ6dcTATWxfu8gFCyTI
ML4ufGtfKIzsk/Iq7kr/xxtKnzOEHUi7foG+ebC9b+AY4h7MJHt8LjxHs2wMJsjFEoyE1B7SKv/N
xrsW2mu1zawtgOWAjbq78HzlM6ezesFpzaXFHPriMtfGniRnzm7m7Q2GFaABVmeIk+eyBSi342TS
3RRqgY2cDMT990CI9b3w4gD9MHp48MtnnB3fuHx9iFiVDpZpXm2ccLDEk8r9T/SZfBrqRtUaBGx9
BcziGWajqgdZC0Mx+EPtyMuro4z+xoddDq9eyHB/Zq1kcsLCkVC2KOT74RrH8xFjGSfYX++mRFum
ESiLnalgB8OPFprg/C+n/QNGU45OvLlApcdSV8ne7u9s2M7UIAInvQSKB9BR0RVgadmgtIo18646
UdoQtAJ7HjOSoXQm17G3Ajo++Qz/PEbAsioREKwgmNZF4Kn5yLlo5GZ8dTScQ/hTcGBh0j2npKFV
S4PZHsqTGkIUvdMijEkC3bOrL+wnTDUcOXYjxD1Ir8aFAYfyevugizID5P6vMaBcLAbTcJSySDXC
dC+UKCQqd/D8wZXTscP6Z6bmMF48qYoh+TjGKjN2xywVH89eryl/V92Swjl/9Z2Kg26fLu9F0aUS
bqCHCSnOD9Miw4QhvZEt2+iQTbWs78xHdwWYyf0iqNXquF9eoQxWw9iqrAduNeC+St+CEE5Ez77f
iOW+Q4k/Kxe19wZ6BR23ItQ3m/eWCBnmfQb9aJXkltM7kqxGcjWFFBKRIw/Kh7xtf1/xBmGRhYT9
Zrxhg/SIgj6tThiWLf5apwgap5Y9mkdtyqS4taM1ML+MbPGRWX5aOuB78CKFpiXUtpMdQbVXZ9/z
6TBXqR2N+5UJsZeUd8gMoC1o88H/569zx8QWvqTYfwRJKKnZ066moaDwXvD1BLQ9cgxOvPZLIR0T
0nekOkpq/hok2YMCChgaGVE55lKG9LSreA6XnP0A8DqVb7it8Lii0zbqQmVueM+cNhLN6TXeMs6T
A0y/l5TJDMKtGqrZsksc/1PAbWtEVeBJ2GisCeeuWqIo0iEnAOpnjDkPYU7LBtHg9W3U45upTVYT
fUbWSzs5Y046tm5Xt6i6QEi+yyz7vpPb52DULsJ2046a+/1bGR34THsEzBHwfyv0Z8b0ZmqJIcsW
XFcyLRPODKiLcBLYp7fBFggPgkTU+xWvMhWgVhZNInWwvB/JH48/0QhsIyB+BXsP5B7tH3kMi3e7
NZUyCb2iui6fGKrSVxjwL3ZDehVofksoqOlKW5nh/g7fJSdceJp84d+fd4yBhLFIgOK+GYgBPsmy
GBarvE319+cZ50Z/xNDlKO0PFTfcRrI/oZJl3BMSdJHRG09tXKAW5G5PZ4mbUy4ZcJpmvSur83XI
I/K4PfP+E7IvatLYDi0ORDvYMnWUOlt325NgeXwYPoiy8/OIbvHtiVcz4Lu7XllTKoliyKSGE61H
i5zu66AAhzZaIcjsSnMbkIOs8Z/+bQyyrpFbJ8L62uPqVkiHe6iY9O+2M06hAXPvabUaw1tvGjDV
IC+CZfAu7DKtJAmB521j205KBt1OFVg7QlylYM6T2cMgXtvYUuw4ASD9hiflHM45Jh2NqisKdytW
XnQ2VwmmWwCH+URwoFxtzlzuxj4Q0iDgB3IiL6wRhLXOLmQtYa0i13yIQxceWYkx3JAUYnOuW+vJ
iuu+lhyvwoAtaqOsC+UzgygL4BiHptf+SUgBi2lswHyQqlVA/nlv4pxT4nBIkKp40pIoOX0Zt+S9
JTCtn6QCMNIBrigaOt6QCwYB+vV+NWrgDi1wW243o6SpzfTxA0su/tZw/18UgOCVJ7ZqLYzYiGVL
L6lDAd+43Ev0pBkCUCKlP9+vmDNqUihWA/uQ2QdVsg+DTRCalFckkq9j4GVWbvYGm0vAt2aQ9/ag
/4nhFaaIfZ/xFq0UNYdrwVDbQ7Y1TEMP4VOJqN9QX8oz5WTD+x2s0FbyLWoASsnX71U0S/RfWHAD
fJo5z5/TBP9KCJRHSEFUDT8jY7mpscqOHbZ9cBijnRXosTDkSg2LernxB4BCkxbsfrLoUMx/DqcK
hILBIbeXRA8b9dk4Bkx6CwhUVcEwkvqcpW2aGC0iSzWzOApjxoGi4t/PSByrF7yr8d++ymJZXoiP
4zVluiNXd1/g+rtl3Oy047q0zHH94z0qYcgwjD0xh5y5FxzLEZc43h3uPm9160I7P0Xw11vGa26J
tLnHizblpFBPo7bvlh4/weopg227rEXDfykbtx/7M66pUVkc44NMasCL0To8ayhy2cVS4m6hI54I
7CMhEGjZnDlo6e3XyP+jFzHhzCBxVAP5bZedtdkDv0xAQO2IjMnY1OZP9iho5oNo5VYV3qNIcxMh
b/lwYaMJ5pJoltJOep1svnlWkRtfWMfEvEwPFQRpzyzDfrdQdPs8/eU4c4jdrGkN6If3LFM4/exH
w6RkMmpZP4ZQBjkpOvJcXA9lSVMQVsK5XFSQMxxfsDBdZbGBki0HLVXAXFM8dNhX+p3vxbh7EybA
WCZeVZYbyP7WFqmBSot3MSg/gdmUkxVvP/HHdbYKl2iWGBqy/Ru9BCVKWcJ0qX26d9/v3uCXr6il
XEYScS+sIrnOvPU3WCs4Ik1hmwF1+mvcj3xQ/RDHIApGEalAfZKVbfp6njuJNwQnQBz3GgRFzCWo
bPs8l+9+1OEue4T9RZLJg0xlcvAkxi86w1nxNQfkMzsdCvDZ/3TWAOoYzojHfSVSPjkUJC4ZsVHW
b2KlbNfDNmGS26t2TYsvCsxcBzJiEM050laK2h3JAva6Vra4QbgZoGsXjvQ4E8yFPQ/Ja6onZpfZ
TQt7VKuXgaepYNN8f+DxHDuj9QuvzM17mq5Pcxerv5n6UKDHaPXl/drMe73qsU/YGLLyXJrwt1p3
Iy6lIPmgGRT/pTOOvI3wbVzuSkiIYQzTi1QTyEGBeybP5L0RHs4/jvtPe1zyCIhOgt/UvRlxqv5Z
DdG9PKkgWncGn8ehk7Uj9uJ5vBl0J3+uAQVGGlZI91ALYReI0qXbYlIiuuyzopKnA6PYT6WrPCku
6adqQ7Ph1P65fZ1N2to9RVgd7yAxnbXdux795ghtl4PogHDJPinJbYXpGByqgtLH1cVjM0fIONqg
21lKlku3ALnZJtYXGpy6Jv4gTzWoMo5U/VuPc6NLAvIslEYOvJ4+HJAFi6k5ciH0JuDrBC4wBrHH
H9KEcaxmfqSPPlfr9mxvcfrVLH7JxlitXVl6sj7YIMOiHvhed379rX6m/tHx/7Pk5MtEzWwXRWFf
PQIg3Y9WYZAcoLL1wZ405VIH9xzv2ZNlFS9s1qRc8awbPRgsl9mlfOY35pzNdcEHhKJafmRxn8SS
GFhodOOQlcr7spa6sIszbyrOhibOcI8zhpksi+Ik7Ze1fRWw2jkNuGjH46WF+qBKV1sh2UDVPjX9
7UgMKXiQzS5zCkZmojjv1Jwhw0ZU16b32lkz7/9Q7F1v3NpHhasCccNXJx+kAu/u/Mk1HuDNFr6V
3sMmmGJWdOexDkdvmj/mFJavwKzRSyjNZRpT9L80NHgwHKz40NaKvJawCIwOCji8N2t51IHXsoXM
1gMGc1VIfLQ6e8qw39G2Klh8ybJY63IeMb3iJidGMaTex7J1HRKIlBFTVduQOiuISQ701GnMLFbx
ZeBS+IklerOoVqxduJsDG/AehMGT3eoa2gXgb1jm81EQ4NZmUlwbqZvKxiiWRmmDzj0kpqG0TcQ4
Iz1UNnDZsrN3n4khEveE9UwYbzqMCmQo1zdlsVq2hRrq8cRuj4xUaK5GiSka/hbGtWWDo+njcoN6
X5TqfNl99xKopbGrl+cwlhw4ST26cWoMIjZiMuxOeBS37pDZg5krVO7ZwXfqJdBj4sgQUVh3rxsU
NR6i3LQF6dPTUBLC9Jg6XdfsErwAIJFYaUeAb8hk9oPSQctPIGuXOrXTeIIJrRVL/5b48/nNNszf
XYYsz7pyWd2jRJ8cObTwsrFDsBo3J+MTZkLF9XBF8rS4ZG5EWdMe19owrDnx6i6ENn5h6Tmmjdyt
x59kVr3zFEM8fdczB8QqzTdhJH8jyKl7TwJhF321kS12+8SYpl1y1msBNcJQR2xubuQh0eOtt3TW
e8OgVbyMxIkpW1NSXQOIoVbH1WkIn6a+XXnUA8CD4C6kxBfkFFyoEJuSEjJypXvtOOBfwTunyMUz
cfhmrzmognlEsIG+HdGgfU4x/5qogicjezRHOduENMal1jJsH8IdLzUxSouQ4iOqwsPjzRthg3ow
7QlCWNZtsifBfGPMRYsWxj5VNj7PUUfq3Hx3Ci95VhOyHkLZIta8r/MWvk62fdB8vmXrSsFaHREt
203sVFGRHGIb/nwsRVikW8+UF7y+I2BwXJncyinl3DItJ8yKFebBGmn5WleqBptj9q9a1US6n5eK
VulOPL5JJ50fdkMg0ko362eUiIma1cAqe4sga89X6eIG7twE/LtzWj5RHqznKDnwyHRlcX1QOPjy
OUJj/EjiAldA7iRsktNURhpEhuUlR2ATMnYahN0ECD0wUpuSMaqr/h03R0mWOHGe844IXn2lNlNW
Ox4+HQudI2ixx9tdz4YsB8BSP5vt2O4n/IYJBBTgZHKpOL4zyVfX6lHJRkPVw56z6PqslswbtmKq
fBvv49yPXgPzFFJX2cJsPfhdhIAwfl0cy206phiY3FWG71QzE1wgRGSAd8u8SwwsaD4lk/AMhVt8
mwFM0v0Jrpl7CDmJtbSFXkb7g1ERSAGGlCZnHqf/wqhaXVSVzpDQQXsZfl7XzrCvD5MYNRu4RbxW
83OL6Dgq1cFOL2fH8cKl21lGywKHQPQDvjA3W+uwUAC1Wcq97e4jfYCJHO/ztG5TnIomczhUL5Ju
SQ2bP+D0k1B6H8mBxXEJBgdSCv5PoVobT4yE8YhvwtrTxqwkK/SkPYPXuHQxjJgr1IoLQIQHhXRI
i9uZx3yZZ14RB9eX9WsOQHH9kvyaZXjKWReh0Vd/ddp+XXYihAxG6bPWUrjS9CfZeIH5d33/J+eY
oZ7/E478vkNJUI5C2AZ8uJWF8eW16whW8J3d0FGg0bBKZA6/IEyKUS3WfH2k8b1Wm1T/plUvM6au
q5Gw+9m6f6eisq4+wN7DZsoReEFrzb9BJSimWaLfo+k9gLClZkA83LM8YkM8hkZKuAqNOGfhwKwM
M3+zisZ3he0fuEFYrP95b3mOWesda1gahLkVULijcwYdHo0eEsWHt0fUIpESeNu9KD0Lkkl/AqXl
9QM48ZG7jmwPRPo+RH5qEYOf0Tlw7mTmo1R9Jk+DD3TzljK3xczrFJFzC/QI5NenIbaQMxK/6ZLR
5MOTthSPKgX8mZFgoQuRaW95fSJ7U+mnYyUaHQWpYbFmq6gJuVKKBrNH3TgelSUuHlCWBZyzgNEe
nZcmkQ3xIIMPKGcTXoMXb7Bt9xWLjmZsReBXsQm4GnkMNMvaDxaE3JfHc3KLenzOtQyBCTSZnfyI
ZenpKXa/pd3CY3hLkY1Dl6IMFi+xZjSAHbJG2/rfdLHFuHYqAR28+syRWGJtaTvX1heg2PSbxfa8
BM7vwPCNDWoZ8YZRcj0dlBUDRrRCgJQyyCH5QlzkhgwZwdc+JLv+j5QnnDjVWFHR9zmpvdPJx7V5
7BZMAyN2+Zj0iq8dlAfENh+QjtM9+ZicOYLAE1Detgwv77Z27NcUPqIM3XOar7HdxjdWJLJlqA1p
abGtz+zPbU9MrZrsInh4GKoAXLqgq7GmgYqP8fGPISihMVlb80gGiTRFXweqqF2b/oMfTQA7N8ZC
P0iMSlGzPONj/vYw27J2fPOy5NCyyiB72xb73IANr3Ae3m2qtZHnsp+NiYd1VbbfhfqvRz4/GMss
Q3lvU2TKwsAS22yfBjk+lmqw1iOpzo7d3nLccONCfoN8TuyV/wu+Dkyp8n38lrWtPPxn4GcIwnjX
F4H//o9z2IpYX2oNX7r6AMXdodCyWeymeaL6MU6IfDpQnKv6980bbBxY6ilz4bxyQ8a+vjwKigg8
GBZiQyM4eeIiryR70cl/a6R8LyFPKIG2KepQI+LVImOexJJet53TRulcLdfe3ClCUyIUHhJc1EIT
lMYhqrG7qOE3X0H/X687b8fUm+WIDu31++S2uc88rJGIjpJdOfG7QNZIK5Tuj0sR+0GL9rJajOAj
azYAxPcKzNOtIjpnrXQZ2wyjjkze4lbmGeXHhedeVWMcACvXVhJIf7DYbu5nL74RbPuvaoxjz96P
EGZKuApMjWcf5UygVtSWFImRGpUk3mgjfBrg+DDDYu32Uaj7dvWTCAEqfXJv4HKpAEqmRNNB18TI
A7rdM2hKSe2XQN45W4KqCAodxXV3i8USnVKoGz4f/+Us9jA58d1QTbUM5hv4Ebm2/Q1KJBeebmCG
JYM6hyjwJfb5MiCOxuk4ureEdydCseLaliftjjQwDZc9H8Zn7MUG9c6m0+yyBnnqpnFGcVi7V2a3
G+IfAuoyoaZaTPklfvv+Jk+lhFH+h4nr9JqIlMfSn/VxZ+ep2Vzy+/jX/s8FMLfzqSvu53pR6W+c
msTTtXjmZbugymgqNqs3KxLkOjh+SGeQgdHSjiZv/LczSuWHmK1ixh6zqsZGD1nzcYqGjgJ9Imm/
3z3+Nf59QdzpoiyGfB1/XcSG3NgsO84bMWamYqYbQSCkHtiWEoSDnyDhS6bM4QZkwY1oJbh2uaT+
xQi1R+FwY+2bt7AM2aImVpLX7VCbqZTnbQsmatZkO7JoEGdoHQs4U0zGPtopvUGw2X9nkJRr2ebg
U53OtBdrCTrxkd9tht0IqQElutPymMljPzZxkbfbAJKD60kEaD8x2pu4wuqlr2OcgY6hS4seTA5R
9bEeKbwph8OJepQgqYGMcOcsH3FxA+z7j0T+YQlqGErcKQDXDm2mAaTXwlGt894A+IfvZRNJot+3
7IP2KLBbPpxWCh3yw8EhQRC9S5RKJLSZGsvNPBHR9De1+SuL+XxWN4DfOIYYXl/Ld2tRNj0CX/oD
0k4YX3jYjkrgtbAPauZeKGmDuwQbTNngRUUGjvD3xwq8/ffXM+PveMPs94+VRgkXkQxZ5nM72Wix
reEfT3Adj8dKFbgfGmGeVsFPXozhyOecSrPdq7vOqgQ06sSuW4PhSlPa1lI8zYdLd5MzXHLc2CnU
CyAQuimQcNGSTO+Nh2kozyjuNE+K+bnq3e51P4COVGlCxmN9P4UZKLFCE0h0Nr2izndZLH2Ccwly
ocX5KjaTzvqhJQSqx3RQDyRwpiBnQ4xOXyBwyf3wASmt5O+XeKbyXqj61GNNY/min6rKb9Y3cn35
xs2gP8XoJKsTQRWpR3tbxxp+IKgwQPUCYHRb9YDk9zAxohFVINpyMv3KRL0pP/ttPVXz6Zgb52Wm
YojAIUAPBjBK0O5SZzpG+/dZP9itsJ74i1P8q1h/1VSZBqF3f8D/FEnPCjTgftwr8GezeNZhAWzb
Wv7HlINBXJl9Ez7UUGiuCm7thdI2kLs6LFDqH6nN86xMC8lGi7M9iKakpWwohzrGr1NwJd833MaS
jbxPop8py0iZuLnFMM5M9vYzsDRG4CjJ+Ra/0xdg/TZCNxsb86113pL1aNIvEogjgUPRyjikVzwt
DKc/0MwctmKWjOvHmD//bZDjHvdYuwsNcvPr+FU87aF+AnIZg/qEj+qj8o51yCVw9Bd21unejBck
qWySmX15pn1oBjyFCacOBOCjPd5HHEQ95fCIKWuEYOPVEPp5FdnQ4ibkO4jyM/anFu9VqOjkZXLR
4CWpVC/0IpOaWa7gXh7z+SmxycKiJ9McfxZeNz/CQi6be1T+2Ag6kf/Smj/AlX96ujj8i6Ut5MV4
Qmx6+8LU656UqBQfhQl2FEjEnzit6NNBf1L9Rdm0hh3M5zqby6aIeGVk+lb4p/ztkOO7BxM1g+IK
DYbxFZl+F6Rs5/tvMAm+cBORtk+kO69nUzp2T4q96XRoCiUuybvWhlq6qiOA3MdYehaRJAqsLGeJ
34uZgF35GfjakU6f7nS+kz7Amv4BwhIqiF2d6D94hJeAlkwEJV2nRrNqjHgQVFmgeBTkXvotwIX3
j0pPcAi5/CbgBWKvvrB1L2zyK5mtlufjDkvsSr0hPnThmi7YGRex6exlVfsGfWWUnYyxC7wJsQJK
6jNrIbU4+9UnLJO3fiH0wY8SW3BmMGfgqFRPhjZdb6/D12jkVAYUZR+HmJT68VpEoUDb4DJywpN+
lPYQ4BErYgWySJbViq2vojE9CWB2tBuH1ZUrJN2IN03v86zXLFOu1K0fQ1jQp+066reclENN0/nQ
RfFK1FzW1c362eRiXYXY54x2ku+r4P59QoVnNDSmYAI+CrktKaPgFPD1pPSHd2BhWXCL9FpzQ2SW
CosfALHNHvQZNffiF5sSz9Mv7V5ts14oLSmvKPDwYmrwumxDBLnRMzFTHOSs7rP/h+zigyhzU3Bn
j2vDLKWzRnuSxWuxGhlnUdBV8VHEEUh4CGT3cnrVX1F4suZvHtUFk8EJHzqW3hjeooHPjx44mtKo
GVR+6OgeVe2Y0w/RcM40Uqe4nGIfVk0IbzjGkdLfOU2qZ4Np6bl3yMaIqq6potj2eWtd79cFjq23
A9YCzagqVoqbEYDEMMackOyDH65PIlYWlgTvbUz3d5NAowTuorwu57drFTw9ylDcDoVFzKtuR6NN
c1U+sPvHxR6WUNdsQcZSL+C+lvKrJ1dGmsosywud0P39YvFr/twYSPSxNxcc81qTHf3O79lkNGN3
jDiUJuGr8Cb9fFq21LHyHLe13SJNrzW0PWhS+ikkNqHvq88eSownc5sY9Mx4AnYHTKRTJzhYoH24
aLrCY+WAHELzcyi2oUYCYbvJNMFGr/FnvQvWSajX1d6PISTd0hX/q+twyWkxgwfgL8q75Xzksw0N
OJHT+dvGjL5lNUU6geUVf9EQfOpyPovQEwwmOl8kXTzCnmLbgt1T/R0YLTqjPTVM3Ifh5JwYidF/
LxYD3zIDnHwNW0ov2jhQ9O8pO/WiBmf57ScvhOeOJ7GuzypDm7QHwnPVk5vAbPBvKCp+hQMIT5rO
tfC6djDNVlqJG0WOj04qD5pyrrgYxokALaXXN/Brgrxnx9cnQOTHM8+yxbOd7iHBiJgXF8Fb9qGp
JRNhCOE+irG1EoBsF0tmShGwuvavQDHeJ8Uz+5lVDXhYAcD99G6zbs2g9kYzrpUHAULxy0i7bBFV
BvLyPPMup4A8Q79oPBCNeQanF0IWQnk/nuLZnMCXw1+Jegybm3jT9vAycWQJFlycYcvegmtQp6t1
060OK4Ve64ytkbiefThUmGVj5O6z65Yvb6ZALWv9NLMUn/zQxYvMx7uNcffi1brGn+ohIa7wfQnq
njjWws51cWNCk1Kx0OZQtuTLU5hAeXrPBTcQxlwOLphaSy51nFBjGizdFP9rQizEtLLAWRYYxND9
EgkjC6MqW6OoiOWRFGkc3/UjSHlXTnQCNKZAqra6KnTFZsptDldp5SzwU2ZnowNeJWXPMnrfq2/V
1Y+QXCoxhM+bLNq2JMFZIDxDlgs/Mds2SahubCirMCJu23ulz42zGlnnA0AE+JiGdj91nu9Npv9y
AFTQuxK4RMYReO5E37MXXrPBN8/OostrWWBTwBpY2pQL0PVUPziT2Wurnf6e5AYCDvcbwewYIIPH
wgrzi4UE/70Qlm97zBP8ckAbW0jkDKb8UH8d3v5mTPN6m6rBxgwJB8Rkhx5e0QeHBY9zDlEnQOzD
MCRJh+IF0M5sIkayJMf8CQ9oVTtolL0wm99Tu5PaN3nQ3V/Q3nC5gksS0fO7fliZlAzU+T0AvqDQ
GV2/8LDx124bWE5bgDEGPnReOxs/hjq8j4r8PnS2mPmWCZWgb/zxnVJnnQDGUzZqtbPvYtshLN7Q
SWvZSy4AsVnsCHRXFHD0dodNVVL1bRVEWWBx76HKQ2JJuN08yum4T9EXDyzZzck6c3O5Huw2uf/1
n1DdwAMRnb/hiaGHWmZx1DY//6GZhP48bylPNeMd7hmeeyAU4ySp7mXzWeyUTgM+vDSgH+nJeRPa
eybZW+6MlItkeF+otnZOpzBvunyT0S2JG3ScClQL/wgrAGH3PBlklJinw9pc8ywZjZKgd7u1CmvD
v7uQWerMw6d7fo/5ClWvFXdpQ6c0u00A5hMDNEU6wTTHwzrNVc0pKUp6GxZd7WepWdjKtTKiEpuB
Qn9UTIo2IpmL9KRxwlGVfeAaTA6z7kuAcrEXgzBjgiXZBIEZOXgn2iaGmrkoXZnp6IfEO7rKhmSh
i6Guk/3aTcCbUNXqJI7NaGU/ARqbnDxztzDk/naeAhz2skIJC14vuCqvmRLblve7vat72xSPFyxE
LXp09x4nXwj3zI6hBQpIPDiiOo0WbB3GeEPc1GagCuSw6v6ZJ1NF2faCjCCghhwkoo7gm3UTMT2B
6oQtFUYkzf4dVZn8KYfti1iLxOUqPShQM83Jwm8t0eOIFOjO9FIqnJJ2A+KsNlzDjaRCzzz4PTMX
R+BEQfIDCMot/dqqgsminP34tPrj22YecbNobKu/ChkBeDjZ1XbH3c75yfThYuuETQDItEC7fJoW
7+vYwQbQ93zZVI9Bd6Tof9JXOeZ71MIwMgTYKvIhhGetf+iMmhrPK5TyN8gZ+U2AhRhCi8o9QB/r
ODtdPNHIIVfTgq29q+p3wf3HqtwJ2R8DDXSC6/EKI9cl21yeBBsNPrM6hsc1wYWgmu4nkp2VSn0M
OBJslIuRKOvKxL17UK0qHWNKlKeVvEhr5py9mhQqEG2pmVvxhfIPbtTHKAbX8UyNY1u0+DMDNOxa
/YobClC2BnqseMkUvaLgrl4AdluMzAMSHEWwhcCUnnIkWCnZ8muCpIPZwrb0LGLiBvwx/pV6FQmj
/QaIaODoold/7GQHhIbkH9rd3ERgcnXZzzvCBoeNphz3Jzr/xno1dR9ZPnHmEO9zDilBtSCLKwlP
hDGXi8I3ajBo3tyknhVfhDV2V+/gVtN/WnxFg9JI7dZrO0k15vSMrHxnkpvngDACIw/PMc27wjD5
8+ZbQqbXsfolkqSuWTPSBRvnTEIvuttGq5KTfFsGZNNij8nQdHKO2VdI8/E+Dth1O1pwX1Bhop0W
Lox9I1d/xLb1M56SiURVF6zZomZ6jtKs3TSGPeHXXQKzGSeOw4jtrIwNypozD1g7ExMXk5Grs25A
3+s/Ac3cZOtTGQZZuoWvoY8OKp6p0gE8Yii7xKRtxQP6SD/Pth5Weo8/uR37zHsUCTpW3gxGeSBW
2ODTMVhcnIgKFW+VTACmdBTGkWLhv5/lNLkMh0Ejve+tHf3jB8B6wSM67Mxyl93DLygJfhc8jUhp
cLqZrLx77asuGEYetSw6h2rqe5EaAoCJn5CE2p1yJm6haV0Sd32BjxsUebQNbym7FIh76lpCI/x/
zhoGgx6ikrIZefQQaTIWpbtF2JmC+UyIZEGfCwpqJdiGhdJ6ZvTRgEUf6A0R9M8AHDJIJ8fAugm6
ucbBbClzb3w10dmuGWshRjV4FjOrf4KGVSA610Nw8M606Zhg6sxDgQ5EzZtQt0TJTTcYTAg84fOS
pGcGJToZHeFW7QxO/p+oKfF0JcL/IKiukAUJADsCh9fyXSrf7mrd/ChXvC4bOz/iu742/vSkJ9wi
M6ZmiWDo/qxPCti/jdYavRJcN1ts0hdA7AQF7SmANoSyGjTkdaag+jEjzDplcGmu+vidHS9fgTuj
4nLDGFxZ2XXVjmEtsJcPet23V6lFEUH6AVI+bUVdcVfYZekW8+fYeNsHMGv2rKBSukefPTvz1ae9
j8udU0movNH7JdVdB+/ZGAWePzCzYn5N6Qk95yaoAnMjiMg+LDAQsVTrPlSQU8VDMye1g2lS8q8H
OJ2Uz81luzmg6bulC6/2crzDaz7JdGUC9rYtgvrP+qDoWY8LdNEofTbNQPXUxpFEF4rK3zCUkXEu
gGWc5oBTb89TzNqlNzN11cN8diLSgoDtnuHEs94g8CuwpPKcDf2wnwtMfkYaVDlgE4Wg8ojW16ys
kDez+iqG42WtDzaH9M+D+uyFFNOFyZgFbStGkyFmktvxUSMUV2Rsn/siD+ojfv4rJVYGKg/DGGYj
CZLmzHtwCzMYCGXbas8Z9GdIwIvbA4lyqwoHOhGlDhhMG3tePPTJy9z/Umjjxg6olqmjF+RZSFal
CUw1BLfZYha1exGpwH9g4m/3PAE2ezRPY9AeUs2Mz4aZSBeeV0RCne6jQtILoZEnTKKjLDoHST6T
VWPYI5CdEhvTbMdkjtSGG7Olqru7S2LI4DjkZuGTpYtsZL9b5N8qs4nJpOZXhAgiluvoNM6lhnHD
8nckO9qRzwEOybXBJHsQDs0GEMZCzm0OltEFlBMjuQUETDFTBFmbQJhW8/pUX4HUXAiL+X0nhsUM
wUJUTmmLRN5n+IUmSvNZFJeuEOgAlB2EIDgff2EuqQ2/mS4svjuNRe4CzGsldUXn9TUGme1otOeB
6B7lD/C9ehdMy3BUCKd2qNoHM9lHPnj9amLI3UaEHZf/fx3cjgpQkvCBPw66pWvGsEEthcsLhNY+
7gk3ld88CGZLfVcYSURqCV9GBQaNS4FKqwFVAUfhocnnhx89g0cquVfvZfxSK76lkNTcgzLzXgRn
AIqkVNuDh25i3H2VEBbJKWOCDYD/Lce1TAMgyuxYWp7DsIxzIIwi5YkrpUTn5dHI/YP6ZH0shc/C
45XV35vqkLxTkwKhxBumpoPifgf2dLv+T8+aDo+tMBtszRqYfnZfgl38Ka05tnyzLjObx8c81zXC
6qAphWHIYhR7AdaVmbDDUedy+wfHwEwBzVjcuQp2+AK8DwqVRsvjrvVsO1xNwmipyh+6/fMAZawB
TYqeBvlgEhJhDi47ED+KgR/Jika4sze1kwshtl/8Vm8/66peGoppKkXxRnZiKoukMkNuQ2WPFnm+
L+38ZzOqrZQoffaHMRXToU9Mvb4C4db43hVbvHIrEKn9NACD7jmsKuL81OpXn1xxXEw3Lkqu79dt
ZNKJhOnYeVHMW90ub/+n7P88pOM+x8O7Bj8pV0xyKeBD+BzfVyOb7EK2bvnkYBpCD5sW8Uh2g7z1
cfYQs7y90LLjJ5yM3YvUavOaUGXVvzuBLl+xHn+k9HWoOGPGcFgTJTroPZd1qSYDzlc3TmShf0kS
JNgZmMVpuSu+Yjewz9Ru/kywB90xHVIYmG33F/59yfubff+gCVSybWF6x/b10Ik3ccVSnamIKtay
1R6XMZaK5YP9ARx+V/zlK0R2tCyG44hYz8RpgTy29JlWD/c8/hoy1uQOSNXb77fGdLTz73GRP5Vf
+8WAFYorDydT4lBFSV4TheQHoDxc2M2egxB2o8K3Z4zgVjdrohA9cMNAeQXUiBPyKtLOYucM29LP
Hw4K81CdCT9vmvZq8At7S37gPnC4a8MI6CVWF98Xrx0desLAJFePr8DhLm8ABU28nbVbWYwoDgcB
EOGhE8Ey+jDZvDTvYNehvowzwnU15dxE2Q/AtJq0FwbmnnMaGdlxfPbFfjEdWzLi8cTceWPgwYls
N+fCau6Lqvqi4WT9lZtycAmhz9Hxj2tDZKNyuSnvlNyv++604Ls0yYwW+4A+IGcL4WyitYC2/33r
gvObGe+V2W5A3CQDW25/ugMWY+q0N3tlzTojtY8aC8eXYtDijRW480wZC5BRkWoalYUJpEmAgeIE
RBF3P8bkX+d4DEgCOs5k4YEn3v96dS11n5g2Ipia39c3/Gb4W+m84pKdGN0Vouodkdikg2h7c/UD
YByrVjCDlo9n5o+lWYT2MCNwhBWXi5Q6lKqN33xXZjrqIq70PCks1oHPXEgs8Odob50xKa7gVLb7
9fW2NLVMTeA54FKPHfk8zckXAkDphlWXSwzcoQLzFX0O22qd9fvVJHGrCJgovfaZ4a7htSsHN6Rr
iGvrttCY2bB6JxxQ5QalYh8bmQmSAX7qPiiNvD+9rDGy8wys7WBr1Q8L5c35iF1QKCESEp42EwQ4
3xyuD1PrK2MuV7k0mAIsXkgo5WumBq15vhshksZ++OvfV7Q4cmdBeLGtu81NLBPgZaB3C96IYBWw
LbmTAAPNXgHTbMaNfI1jrXnd/pWdpr+5faodNE+bIWHkbUFDqhdt/T1LzeNriQCcTrgF4BGcmkGU
bpH1o5CmUFyKn9ETRNP5MkQPXiuA1xeZobuuVYqMqEi0S7eBtZKhdF2XRMCADiB1iXQ7GjrlFhOV
MULBxFK8cihGGZ4IUzkkKflF2q9df3YSAKD69jxeVQbX0NqDXzQFnGhx5TKRq8v1KrkjAPwcRuIW
a52sA5vx4sxVjSSZSxCv3Vhr/VadqNzVlkbjD6hQ/JhnUTapnDLfRKU4ZhMIlSpdxT2+Xp8m/AQS
GDAsVnMVi+jDH6sj0VYX5G2H3QCw+gSj4jMVkH+1WBTPALT9kw7qjCyxBk7vjG1UFDfh2S0P3Jbc
qV0CbPGbO3OlP898ycSQWJtWC/88GEELBwXW+oSMAY39jfCeOqskBgeZRATynRP2mbMfWWz6dB3l
HGsKG11uOw9OX1cb+wyC1zbFsjr4rTt7El/d6Jh3yYgxh7gQ+roG8TYOJnFn4RCwsyBePfZ0gVJK
WNPfRrIhP4d2p6/U0eAjrBQw4P4Bj8PSpEOrfgz/1SLSC2CU+yLdYI+dtPV4YbvE/k+DnYzdjqIt
HdF4T2lOWK/Gyrl6Dz4EiP9g9N8pphqRHGgpn4PmW+rS7Su/G62fqnLk7mur1Pgyic7Ww0HnKNg3
//NlEGMz8QmUiEJ0bawocLdTBdBkNhT1fSJ24r3Dz4HwaEynIwpehRjByNVwzrouZre6mF9W3mPI
SmcGRGE/ksDrQ0OUqzCYhGw7yhVp42bb6JnJkmc4jtjMnTAErzzXHokSyUpjX5R3YataT9qn6+cV
qYQhv+FZ5eCGyYZM2MSRElnrRaKvsJaOyfhSgOoeKW9+fWtNiwCRBlO90KUdshWP0Tx4ByIkcQmW
KuODm1LO6NMktfOEORU6TNC89kHFT9Peg97X9YZEb56C/cT3lK7P57FmLb/Qqxyb90oUIGIOMbHi
a4EeHrsGbynA2PbZonT4bIfOPJ9vsU4FASUxycp47XGZ97xbmUfRBtutVjjeNtuH04e1nNrPMrLq
DvWr4uI71cWZmDDK34q7t067hUwzXVh+UIZw9FNyydDRy5CJvWP+dN1Q5bFiCM7jhQRlCfEamTB9
BomHBAQBOznheqBNpK3rGAzKL0hZkLerOWgtDUrBNigBnwS+a4rmfEm8lrxiiKFINxBY+pqP94V2
IlXWMJRe2v6EiHja//90YDO8yNQgwdcy7jDq2RXkN9YVFgZMjVtoSaZ9AyuhBWPOgM726zNv8Ia9
ohCrW7grt19Mu/GlgtWrObJpNWSXpywBORTBr9hrpR40xklKeJTibosJGxfdCzcU3GgbARUT0LzI
f3Rt7jwd3A9wSbCL/Vqfh0cO5A0SMf93ioIFJ/n7kQ7aA2rBIdn5Xg0H961VYRhtmTxOW5gf9QZu
u14nI0NZMvkU9BwETiHylVvQ+aqsAHgOLagrDPw4BbR4RBiEDm33uYLFy8k1rmJI7YJd/p3kPg0C
RR+BNJwD57006y+df3ktX9+8ZgYApaFjhPxrfZaaeEq9Ykn0yTRUg4PezfHZO2SGl/sg+9pXdv9Y
wNjr62hhXZmT1Tw45RR9qZwvBW24ZlHeLXFJy1qrkh6OuzhPO+bL9GD+tm2yMJF6AgtGeSFtRb6y
jCUDqe2SftBJHYDN7OIwx1SQGW33Bd67C7hZ8PKgY05R5Cfh4XLv8MjVRANtZh92R5tvPocUb79v
sC+MHfcebgrNTliXdNJRqG/f/6KG/BykB6qD5NASPKE1wTJHZvUFUMljts5c6/JvTH0e6RW+CUex
RkhGQ+/o+yrP0XGH6QiBPuY9S298gy/aNV9gi20ho7G3QKqxiPo6Z6bMaobjF+24XZXsGotzfdGF
rygBfdNcjEDwpjNFIWJxj+BwoTL7EsXx0ZZZRRXzpDCF38/hRZxemA+90qvF0s3U+odJbS4Oahna
fj+G9dcLpXJ1LDBH9Pi3BpVSIdS7FIOaHZpNs87KQihzvf3mankt4G8/NIaCQ6D/SKfrTZI+goPf
3NWG8w5pbgWoGq902P29F3RrYJcLRQwOf22zEIrMUFut8T2BJulDn2JpgOUCZLjJJiu2Bh0XBGkE
vDi4ta+yflhFSYz7Bvr5YvlTiit+Wf10SZyPSJK0dkpDpKMY1Jow4WXRK5EgGaElyeWK19QZlB2O
KcYtJULwEltLEeEGVlmTrxdS8NFpDVchS4iAXmHC8niRAXrVk1DgPGi6b+Xn47NVt9LxkDzbJrFP
MFaZM32XvyA8IKB9Zt4ppUiKRcH3olnMOVkh+BSvJTOato7SrBv86SWri0yRuJXe47dX4Yxg0yun
e1+RR6+Hyi3zueY+JL7lwxz6pffn+1vzLVFRzzpPiWnizLljsgGpkki0TikWP1ESQXF5ZmGnCZP0
48qEduwdS5cu9mZWXRfHbZZnWV+0pDGuDuPdpg6Hv9Rig1TIB5pNH2SwsE7KL/mqhnlFieojxOpU
NhMp6dgslQlj7fBT7117l0/+N34yRM8g8s617u05Sr2UjZdbcFWK+qJi/pLU1wWs+aJNc3GJn2Y0
Fc7T8mHVj4tUrNJT4P76juBsau9qz/QuF0QwarXXyRJwNmCEDKbfUiLLQn4ayuOxcCpukXFi743d
6bEPjq65FjXKHU5MMIJZFJVSLe2lXZ0jHVGQpBEA1BUYRIrUZnVoyyJVgrohMOPLMC0HnRJnzrAR
O1zD0XtiGxEAVI4esMIvADp1Z+KEZn9VQu2obkiW9dDjj87+FVdlenYJ6UA11863mNc8eElO/09I
BBPuZSJkLhVWNTx7xI+WS8pOOItTh2vlfEczUNAm2MUNzOtFkD/BB341Cjmu7vgOfpgr5ZEkvN+7
XGMH+l3L2e8y1IN5MVP3XJ6fmrAwnDRvT1rDvULijJMSPzBxlfSiAi0oD+R8W8QGVTJCjUeFU322
8Av5TnsiFp4Ma0RNbA9r5tQey4BldDYDsruwSKwqJcSqDdHYGv/eQg33o95kaFyK0wXFSmSiJkZ5
Y0Qny/KferMjjucjMpO36c8Qmtfxk/VW4hJzDuazGzPNF9WzwrfYyf6ZlTZKJtVoQz+PlyfiHNhu
LyC6/OGJaBY4IrRPKYNiI7RNumQLepndp3NwsrJVLYDxxRWsnithkLFt+d3DCl6in2sBHwd/M1r3
yKq6duyo/riaIlCujHCeNWiIZagdz9gaF6cvZ7VuYEMEEKKR3rnDOwERoxd6sNv+lrtJi9+3tNSY
DPOiCyBSrl/DdahuT4CQVYFJnvGv3QOWTvM1LL0XV3ytwLDvE2v78sSTCIDbVHvlWuCcvF/ahIDv
wsILYsuLCKMxTSYWRiB1WHHv6cKyOH3VTvmxsxO51UGMze4pvVoW9SF9TxYPxLs/bPTOdnI7JBxn
6NtmYDLYL473TLWPq5+oWJGk5kMcGpTQ1gkpLQ9AVFMTLoEvyl8EDgS4dFe9wDWg+nqMx0tSUAEH
Gdu7t4Z3GHzWTgXQPPfrrFUPT8w13GyMaRxA+/Amv/3K69oU37NTc6PgcqTiO8ip/KNYiMF8xHLX
jyUtfDFGjlbxmdrKxCpBA9H6lwbGTKsAZGGYjJQYZlHWykE6TkUCUZWNZ2G+qV2RCKNdV933ihTO
VEYc+L31PQFzZWTcmY7/NcHmdBaGHhhfX8tuDZ2rV+hw4RXR01kW9WRCwYQ3idHt3CHAgD4TA1h/
HpD1R5ODmq+usGFaRARB7E/ZRe+Ts8I/ehi4lG/aSpX3v1LZ92SP+IxMXVS6rw3WoKV54Em4b6vp
5QHfahKpoOhMxFGZOhWVnTCEsXG6bRsipINBgdC/jgI8frF5wUO6C05IN/Dk6hnoKWvMtuKUVtFR
qubzxqdkRLKYDlsC+wfzp/H04lveJbawpaZlxXqp/lLG/bzvxJMGc7n68cStVUswahgV/Oaj60QV
HTN4UfSapyUHTKDnKxwNgRaRAbWQ7d6KkuFTGC80B+b0I908izbIJY9b3MgTAKBt++lmRcOyXs0A
Jsnus0F7cbBRfIxGjb+TSz37UcWa/Ob1dF34CpZHGlmvocj87SuhosubBsXzW/bf6fSFHmSgXp4u
SUBaLNmSg9Xsi+IeZbU/B5dw+xZyJqwbWLA4vm9ku1z6WgvK0Uu50PMrRPksILzSVWux8IinsQhR
TzX6CJhfUy3pCrstmgfiByiHCL3WnIhfaVMTOVoQCi+eL0wuTo5PKjoFALqWeghGhbM5W0dsyZ5i
rmD1m6lwuO3TEHcGS6UhZEW/M1/yWuXJnMXDBZ/MkVsC1rEr1PpvxoQqIZdZHZCH1CjyekiSMXEm
P+fW3aZFm/AcQD2iehLGj2fKhXSaU6MbsqwXThSCp8wXEydj84lQQFCAb24pfYD37wX3hBamTNa2
MpoqJvCPvXLn94dpoFAWE23oMlJpdCYZNk6uCzSBeZK3cOpGpYDF7x7t9enS2ZqEvjkC2DxAXtLX
n7Ks7O1vRdLRu2Qz8+bUGiA4QDN/U+PvVwr85izHU7DMTrpYTsus0OlJ9Bm6FK+GCQiUukwJaqiU
9W20JsYLuoWT5OFU4WrkOsC1QeJgmuh89wQ8yxU4xKtFNDFLTWv5AVgNL1k/cuaWjChIWy6DEW5G
JsMwzsXrDIrtMvFY/XGYjqs8Z0RwP3TrAiKyL0hNkity4MdI932i0fDZYXu3F8rwU7DJ+wOWIWWZ
sSdigyPXkl2e3md8uhh27SMkZVNP6daSyr9U5nUclOR2ITAs1Mfx2z6jvstuAo9KOlgIg2esYyP4
Wm/9NdWX46DXd00ZpJ0/JuYYNKLaRjfkou9SbvT1SYvQ8U+3L6G83rZqAtv0mOoNaEwXb3+ZozyV
LTwEh+6mRD4uATnhOc2f3Bl+7fKuODQpaWApe5dhhlt8+cE93q/4zrQ6bAkqozh7046ym4UzoyaN
1gYGFvc2IIan4QfQeXxiEy/E+Y1K4GfhlVdf8HOes/nXSQT0haTuIbyx/3RmUU4QyRT9GuLLNe73
Iw6vvYGPnDfWllbFfW2kk2Dy3xU5R8FI79yGcqdAeXqkHJsEPcCpNYpl/YmWtuG7nMuulU9Bz10s
bko3sus9B4e4xhWul3FKfQvi+q0H5CcQ7Du0pJ/HPeltTHSB3eO/oxIkOAU3JjroJG7VkalIeAT4
LYSKQU9BZwlKvp5z6b9ANq14ax10CUOFbJHSVEHdG7XlIuJGrsXNYP1r7nN7AdW6c8egg2ItF1wQ
hbLISYJqPtyBBc6gdGMN9VLs7orlJbL1gWVpPgrVvNSbcyoKovtvSQtCA5O7Xf7k/AvOdfIRD5/P
XMG+IaNDDExLAvYhjiiv7SsdPOkzxgtv4kLQG0P0Cvkhb2iNOxxrw8geaVk8pYt6Q5glUfzOiAE6
lXD+igcLo57KgRpMqnz0EF1a32/X3QgVBZrtaqRE6P2C7lqSH+AMvPPQecVR+cT4tTvzLKuSd/DS
zCHE2BbIQ2PyC0vuoDD1e4oN0EznZDPc7GoONeXVOFxxD5MeW3fnpZRdvNyld252VNA4j/9Xom4L
uXOlYK29oXcz4qOcXAZL5rC84aFJZDY5NvKA8LokoGSGSD8khHPKflMsGTSu/+dgqdjIp5HC8cZz
1IyksFfp9cpvruqBEbsRrmgsQSFc45YybceXAKqUkPY14FlSVBFKDwj4Hzl357SywmxWJe88GM1y
gWhvVoViFBG+7YTcnvY2vVSG+bUSIikvxDNOn4RY8+sX2/KgoXziqrHo/I3HNYfxbmSgNQcj8uDh
hrydrJRl6VOghOEsVzUSyjHICOQQYqVB1IRniGZ52y2+HcwuAOuWBm4Vi0YWRK9axibwtf8Z5Nox
YQa7kzNOZCvEznRZaH7CAoNGPaf7Jcl5aWVSAbI8lR+wpJDSlA5wgses1dLAgZnJygrVZiNmgbbP
O5GVLI8uDdPVZxmt6YfvU348rSeCVbvMlLbAy1NdNIslnSBnMuwtzlj3aRpRMSEZjDaLsviG4KqD
wGwidMWj/Io5linwZ2SFf8lplmyg4A82vjy8ydV3m0/EDZNIju55MxgCfR8oJKtSumoeAnBvvvUS
Fm7L3lUG/EgHA/by+2bc0zts0amlSjow8mp6hu8UjUvL+9d8w8d1ipvgZaXYOJXQOjRrAyKaASgU
c8nGOj0V/LIwn8jHCqHqx7g3Bowbfdp9CC0/ZmYoKdir+Jt/p1osU6BaguZ/pUDcmoob1dsbjkHv
20Gqj4cnA2zfLaOueRxOKXNCTvYsQoRnJUKfvIwgvEMKMnbMYuLhoIhC2FB8Jk5eQphsgMcMJJow
jY84Ck9Tfkafn8nPZA3TxyliI5s2BnEOZgNhF8IhZqlr41YjyE3uM8tNbK8XhE7ZqmHhH+Vh5UgL
MaHIUNwomQo75b4VSWgRf4QiSM3VsUh/XtiawKPCMYTbGY+itEQyDSBSevZOv3AAPyNBSLXhGk6t
dkOzdWqMbZFEeVVcdUEtTD273AvcyQR4gtt4Mvxc1XZhFVlPkR9+2Cc4ykY6gq+DXrw4b9mDaQ//
2LAjXUlA85LViQCSm1bikNV8j+g7B1u+RC06sOV3DYRO3Oa5hvl/mv9XOuCOBKiyS1JFA0qbGPVt
PMu+Xp9Yu3VHo4YC17SzUR+5owegbIvIhTkP7cSGUI//K1a+RylsgbYQIoET5iOm0r1oCggiH/HA
M1eAhMm7R+QrXxO0uD4Ns/NT/JbtKMwKDdss9PWe5as0NCT5G0z1sar8IG5ScELxhRY6Yb+NAm+T
rGnQC2KAdwOVPWJFg/Z9Go1b5JJhWKXbO3Akc1BGBmy/AYSW1AeB1NBE7TetA1H7p5APK9KQpbUh
Ii2s2LVamS5tOU5O7pXU44SlXeSNi4BGShne5ZxyC0duYKMV9ScAeufS+mlolYA4N/qCW/t719x6
GZMfvHOE7gHmh1W02iXLw4srkCl5dnz+s9HPik4KvmVB2tE2Bbd9e0kFMJP7PM0xWjvskwauTiBl
8DXjWbpQ/nSyd3eEDPSsAX4xuPGIjOjMXFBs1vUmelENOE2gDZwd8KSNpjrat2RethpFxsYns0qv
IgnEoI6R4e0g5ugCDXDDUfK12gsPzUcNhvhC5q36AP8ATq9lsIJ+9LMHcNlLt9clAZEXueq/cCFp
B9WWL+tMeq+TauILcvD/xlF+Sfv71OqrR6fryoXBRRqzllI8GlQ/wp31ayL6KhFtMXMaPXD0i62o
hNQjlZZKtXrst8QKovzHnbQiLLg1AD09ynIWabfhnKN8Tlbtqkl9Xy6HPch0odCfnNZPxc+lBmBu
nwJgXxROcR6z68f9GKlL56hOFIkW42SLUn80CSK0htlmJj0HXuvfczpUl936iZW6hCf6B3LQ9YqD
NOwSa3eM5NonofzbdTCN+cg5P2nWvY9EFGvWyNhrg9ASKZ4O5N5U2jj7zlezwYpeO2c44BjNvA1P
qvU4GyOCbspGdJbNbv/8xFAnFvYiU3hu/whvTDyQg3CeGXhLRi6krhn5hTGqA9qOI+aWIpMhf5TQ
TR93QFdb9UHCRyNpyTjadKaqhdas7hnDdqb+ZciQIyYP8DNszY1+AnsQa4/yZUCed9IhBoo9UpWQ
b0i9APf/Z0HNFTYLm4RSax5PXoY0CcILoeG4eoM55Tr6I7fjO1avuB9VnlO5Nziiqq0jKY0Lx+Sd
qBSIwTFyxXDzLYuzfYyKtAItfSAahnZ+j/A5VxbSq924Vh35t8BL6Faj78eBHyXBJthdxPCDIfUg
QQgcGWd/Swplw+iBghxbeVkn4wv8osAXf/cdu8d8G3SEwjeMUy93FpVAPZIo4vnGBNb5b5mheAeZ
c6VIJdoHSi1YGEMxKoIQu6o99tx1InjT6SDB5deOsscA43XHDCqvKpXvcxZ7B6zjjQOcC0NIjsT9
bZbq+rYAPpPgudeKG4m0pP9sSNA4/PwvoBs5nhIATDx0lwP3tp/ttKXAdLRz7rxY7fOcPp2Hj10T
gc9rgeDOtsznFGKD1Q/IF3dEIx1BCAueQtkRynQFp9uKMH4oa7rXLJSbnRT7Kx0p6o4zVbbOPhqM
GiTBgzSay/b46DlAshjSnu6wwNWaGZFC3QvxmAv1z5Z0DGj63W3jjRDqcQYB0/Q9UX/hH8Lj3BG2
c/0QJNdx1tvG9YbQguo0Awp2G+SouJGzoayyJEX4rEdeVirgBCSpJ9xIgfiHoIt4/3O9Y+f6czRR
LsvmDcWCP4Hu51u7X90QXVbd4OeLDENUb3Aya8YVIjKdDyjkGEqFHmeu3UlaM7IPBhPPDgZd5FUP
m90Y5mznHEm0CnaImmLsyMzfKrMB17YfIMSrPcZkvxHOl4c9rmN0N94qZRuxUwHTHRgUOn6YQfK5
N39G8OmNWo51q4atdrjkmpYRgtG2s6rwvXsGuNEB1JjhPcTso2aOZytj7ifB6f7TofdsFYyE99T9
zd+0R7SkOvSQVKt777+8spzVw59x4/JZ26aNuSZgtO3iutw4D/+YAwk3QICi7fUc89Ioz0x7jwYj
pc5RupwlfLykL5qjHDME1twQhtXRHxIqNq9JwYJ8zlPCefHh7CD+3CUhHANjrc+dBOlP764ciEkU
5M30zmXJo4omksgwlA1LrMS305oNzdkk+vA5dAf0jOg31goc4VLaHpdoW082lbX6sQ1oaU5esoJs
BvWgzfGecydYbDYTZ02mk2IoGaJQ0RAZyU69ZUEJT5PkfY9Hqr35k8DmSJvZ7zPXmEHd25szT1go
J5ctKmSYvv4WEYIcdUdER59bhuUdNA0CmmPtOF+nfmts2GBw66cg+fFOkPGFFjVC+odpo1HC+PUL
hXrClkyHALQurcFgwDkjKcnOgYp2IVgZzXtSy2qEG5kdwWKoZz+sK6IK1b99HANas1p0PaKMKM4w
HTcCJJ+mbjuyV3g8tRJkLiKBcsQetW+oChdo2a1o4lCCwqxAHt92AAQ02hqUIbl6SI9wy9/+TtEa
CWoZ88mvqqSjYjNLQKNNCLgRkc82z58nxFmoQyeqhtLotGhsMISGH9et+D3DGhCgXZX34Pzi62DN
X203diNZVvnmg30T2DAzOoCv50lC/DEISr85/dX3g/P8sK/PXK6kiPRagfrtgIJs8Igz8vt+sGJl
8GHlOJvepWtZczVms5WnZr4HLUv5BO86xti5na3HCxPPG/38hW75lemzxec2qd+Fu3IXHLbFVQJz
idn3MNuEniDX/7v0MGuo3dmcZ2SOcaAe3Elc6zr2jf4hQ/i/V/IIh0IsE01K+qOPFNicCh4t8hCM
z476K9kVTJqiEi27LXP7hPU8Byajl4CuA398KA66XHwrNgcXkCZTFAjAzYp/O9tbp10ZMHnZ0Fma
h0vs/sU4/CV87iKVC59kgaBIP+FKii2KfbIU5u4cCcVVp54d/+M4lsaWhHSQOUw0aPKEg8/h3Y2t
9DPTkGsew5HUMJSow5CfNjxe5zVBTcuGj93cW/fSSwkRyJ3WoLsqjQCOATHWu4ixV2Bu6/t3LP+K
kQsxBqa8SzpghpXFu/Cxfp/X8JvutBL79DCG+rJHw508cBTCEDJIGJoVIvXTom8PRCCjeV3BdJZw
sSWSWb/OVEfJVw1a3usOJpfNyX4ms6smiQOEsa9NQitnpkAmZWuub32B7nnB8DqPR7FwqHi8EPHV
JwRhAXMsPjMWbHI4Q/xmsB74IETKVL3Nq2xchVf4r61pdjSZwtgO+BQNLGr697G/3wHWD8HLYaBn
LY2Ydz8G77ginEIzNIHtz2hL0LwiE/xNfBkTx2hCL10iQ9yu60hMuO68Cd0qxwkA2sVLDh1ecA2e
dCEY5klVxU1C4WM9zcdori1aYIp1hQk1vS4cxYkACsXQggJIcK/RzT3myGS2uFKzzVfMyXoF3xeP
8xnfTDIcJj0aoaDm1LR+GCvC80f2eLqRuKd42vtX0BQ5iP9OSKrbBqt0TIc/C79s7SWgdBqfwyVJ
Lxw0DyY08C4HmT7489aQFBWWwc6+zcUDGI5V9WaRnP+xHCixNxtaxi5NNmmNJhcjq8jLbijcOS/S
SwRtUKqbXhhwxImoG+NhIB/tMFT6PjOVEGETa/1wWjQpdgQz82df2PxZxHvSKPJkm+5N8KvwLsL+
wpIdazP8LeIiqEKh1Faka1uJKJjAgGSLs3KkxbuB4RnsbEDDcO2/5wuA8YfOPP9AjNLAd6vfoePy
poBtYZKQi8OkQVwyRkDXgxxPEzuPkUAJudySbknpEe7+EEBWSNSKkyHnkLw4D9lBMv4vyDgMbndP
q7D4iSeyYND2yu0DJqp/kb3egLD13ggFsm6fxOkkjmOhkYhZ/qWso3yyopJEYwZhfLEEz39wm3Pc
UU+jWUbWndU5SjtKufOrQK8oNfmCKtyc6NO7+C7u1TLQa+bw4E8bXiJZncU0kV1kB40bVdEnls6r
f1A3CuGlOAF6NrB2psqS/hP6x5FIKDFhxwqNV50ss+x/xsIa/gK8cvRGG2gK3FrQyNnqY5c87wMO
Sp2jMR+v/G5bzyCVpgm6XkR34TppmsfrwwOC3DOiRBnohUCPg8jK0FCjixoKh7jnIDWMQY/h0P+X
MSjBpVvRbXMitX6P4AxAWeGb4B1lcahUff3uFVNsdlrNUqpzjK1aWmpFMmW5yhBWuqvzHcGycMY/
5TTxvb/euO1GMsKqsAS/+zQIddQL6hAjcqs0u4WS06znnjceazweKfMenXotyLSCM/bjBxwf0P/E
Y47ghKtJIEcdsptfjOWFzQDdEeiZRqybayJasUzZKIzNs8CEMm2WRc6Ol2HxKty91tUF1g0Znjkv
UjhnOkEs6QI5DsOSQlQBoX0AW+tbqDBlCxWMuPzkbCRlxH+ujC40aaTzNMC//kSTku6OHB9eFsbz
vDSEvboXxIqz1NqqsYtwctNml5HpeOzt+kyKvIsK36LxDAkBySxqqiOPUY/GzhG+SH+GIo93ye5s
Llv84tqT4zGg10Jxj/5WPag8mVhfmRp5/vrtviQP+5+7N8epWT0KE7SCNPyoOS4XiE2rVd46gyGG
VcIfaR1EQ/zUpolDsJwpujRnQipoiDnkNfk6GOR6hA/6QAr3hBqwgZJ29tsYa890Q6B1YkYLgukP
MBzwO2u1yS8T1xd/wF+XV4lYw1+/GzgZdFP2S8gOr5e9+SAj1702BXVthHtzEcVYhwtT3ZyCjMpC
IJcUeYedCMBSVE0Zz1oZ6hsJUqUcBX16MPGmFLRSuZlkQi/vpZcPk0oQXt6t83N48eYELc9NDt+p
+ml5Hpz1VM8WwwGPY8xIevdfVCxIqedngjqXfa7k+b+pMMb6aXIMSE81GptYwzn44jHgE1uGAxmz
EXea5xRmNBRF6qWOGuuq3tmfgDXrl0Wn2aVuJU+qWDS4HtzNpHTFb6Bt0e62RYxpULkjHwSXP0Yh
Byzj8lKeTZ8xRq9piaYJNuue5KnQDhwf7WlMj9rfmkPqUGDmLTx9Cdh6fQt/AWsrVTQLebdKsoPy
n9Xe3RULscYWDUF07cFA6uApNriQncqNiq3ZCfQ1ryH52ZFgBqhQ9RsYbg3rdbLghX09yWi4fNQk
y2HBzSpuYatBtirf0T4tr57cH5tWWFzIljgErZy/HY99hVf7f0qgTN1UqkEfmKL4ssii9BJ8nVF1
Fi8Qg4kFKocaepmQIulFvA+eVcp6SWubb3hEL1Xn1rfN5aKy9jlrjZaR5nDQ6pRnZg2hN5/RNnOL
amldwSYmaXeteVx9dlXaZp3TzowbUn2f2rvRx97dO08amtMkiXCs4sGlkc+3ppLiq3nJpqru/n/T
axIZYh8QWZySYyoVQ/oFliuJvcSPvp2OSGoMagDLhdqS8NX77nQfOS60HJ1wnuqDatNnvYRv/IgF
PkODBlq2rkWN6l9oqwtZtbvOv/i+FX1PaJTUYq3JX1ID6ieduer/Q9LE5F9+J990MtdgzkkrLrRm
1dx1xpgZisG6fCYT8sjVjEyMTI3bwDi2NGFXv/gTCP/f5Cvu1C5c33GVyNSUQQ4HzOaPo+P7HvAM
wqG0coC1K6ZWdp+j5KGI9XwV3oIahLoDTCfKDOs28RW5nXNkatSZ3IhvVZ+eRD5dsuQoaAF72jIF
+YRwKPQ1ebLL2INZ7KN+Zz3S/d9RMF9yPEueK1jpeLEloXb02k5A7590K6NwR3h753Jwz4iS7JeX
iHRNc1J3R4XxmXDfRw3c+Nz/T9+YkTu6eTfS3fbHde5on8NWn5RV+D2FASL/sfJG4f7bc1PVEF9u
Jymn/djFBeZ/7vNb8Y729+4+IaTo8Y8Wl1ETCbdOhz2wtYRhOpKYG+9EcbqSBazdik7j2CiaEhD4
byNe41iZEVfu2HrHqG6tvsKJsm8dbo1wqr44xxKxN0T/t5YxVsK9iwgUTQaGC4zNvT7hSNB84Fu/
Vf46874rohl9fIWl1+11IC3JZb84rGKyVKmJFg7oOzgIpDQa2ug1ZMMR9yPrK/V23+fTIsjeJ+dG
rfgBUaUoF/9W3XFZp5DeqnHEsOXKCAmgvL18trnpAvREkza0V86Dol6wiqDDT32sYtET9OzBryNM
l/wNAOWJERujGG/jsUmNj9aL1+vcqDm5Mf0ZyPXRwwdqwalMHMu7pRbJTBuzyERxIZnixlT4miJa
gevNJzKpilssA3F5GiJoh84mjO0v9dT3iq4inpjF8ckdHwdpfXe8DXsxU48GUq2ln6nb1ciwgMLi
sK6409OPwJOuDayo9JbYw54TDCaz9ZUxHazHgbO+gNsOOD2DbQKfz/Ol6+8M4pMrHc140D9Y9eZq
wsHz5Bb3beCB97SMaGmA3/lGq6Q6IXhEWNo0YSu5c87gXHLIroj3IoZj7Eakx1eNXTXOKjbUt/EG
AyCJGUR+8Jo0AD6Ulx5NmPo4USxyOHlqcuxcsD0iF3j5ZA6O0gh72WQXVywV90rhA8SU3KDPFyQO
CD3WclLECCNmBzbITo/6LK9Mc6brmZHEc+nlXexHKDjmP5bw2MBmQquILF3mG2KVQ6lRRXzZbiSO
Z8pHYusBjY4beyh9SWNRACHBXZQyx3ccRMjHYf+ix20deZcIYSzF3pIY7xPWHGOusNYiGnaeQZ7u
uJtE5AiJcYNRftP8FfoVYS5wWoBlkbNgLz7Pohu1XXK8tSBknu1pcxAA8YvEHOVJd2sO9jzH+04E
nL+gzdZXOk4XDrvZYdI7EOhj/cb+K8z3OfniJSecGHhV0rK/XEJeGlCDVk5a9U7fql4obSlWseWT
rrOSZrORKdKxtzbva0G4Z930gkRPEMHF4xmPHjQyj0+ynJStQzLp/wOEuMGnSrZiV5msc+ij4ztn
39f8l0ZR/SRbBsh8pYnhB8hKsbhZF6d0w/ybIAo8/Vs3jnIxF7exEhlfH5MIQDM/pE2autDfn0Ha
o8xCkO6jNBhL4ca0dU+xoz5C5HWVXEIA/MvtmQMSTLUOoLULdcJmMrlWeytqhwPjjtHRhAMRNSqV
2kHUWykDDq/VxojLDtAkrnGLib3Rn+D0qdDVuXgeJLfXAQp7h1vkTfqxWcOvV/ojo96n4zb5e8rr
0O4BkVn8qYtWT/2RIjsAn6P6lK+0GGBGWuV5X5mKqw4MmHcbti4mIFCdMYLfJ87ydNQik2Yuh5zH
i/DCl4018lom5Yqhl0PtPy6UP3VfmKitjq2XsHpfol4b8o9X0DJ4aCApLdDihFw0TzRGngNbyPUW
D/cNwxiY7cobWLdY5Wup3bWYnECy/9cnMTfPKss9UHU64CBXOAOhRkOieb69U2Xjt8Vbh9JWXdmX
6rRjUhhL6U8GA5GPokR480Xs96K87oTXEKpTI65Kr47fEKaEP0zfVIvHK5S530wmdNOHusCt5dQV
c2y7Rzefk5ePVHtYusFDhKTp3gyE//R65NFLBPk39AtKbxCF4GKm1hQHCkNM2+N/qMTvW63qDP7F
xJCHL8YPFeC5BhSEjq7J37FXGuqnr6b4OWwvUyCUfbuIjUI45rGG+qcB/vnBHV1gDB6CtbD++Hht
t/2H84m0vpvGbVxkFP/Oosqw+uzx+Me7C3jjwbM6f1rrD09ZYD36OGptvK0hO0d3ylhKSfkyXDhx
d0lDZMzQMwt09ChG2ZCJwFBH+2vyDEqaE7uGMFBVZiLxCd0PhUDhvoR81NswkzPm8GdO54AI9aJ5
iQyj6BU9EYfFCrcuK3cQdPQdwKc/85pLHSka5qu9V+2eLe8SfGscD79O1Vlo2dlRxiKZUPt+C5RF
/w1gGCW1R4xLYnzl4hfykO/h0HRrGxMy6lqO0isP3+bYZ88LoViy/LXt0Z3zSjWZD/mbeOzk5fha
mUDGxcaTCqdYFFThZIK2TMLCeJnKSP4d67msrEF2waggbJkOhDo5fNGCTmZqa+iZ+y44UihgILee
N765DIUkW99Oe4pJD355UXHnoRrulBrdlDBIaq0syCYVrdrpOjZz4uQSis5npWzyB5ySwMnlMHBE
yp8/H/fVKNG1Q5+DqKjEGqkZmTg7d7Spd3U5Jysz49tux5hsatw2uWSbvPGBV3CtN3T+aABz1omq
dqoqryiTqgATNLeM8oc/SPG6izZ0fFZZyjCnXjWA0Zq2KeI4aLjjzgMLHSV1I0Yzriqjr9M1PA09
6ES4sGM6Aq8DBBt+mZ6PuiKFj4AFrD3fN3z5JadXl87Cd7NfIho8qzd/qli/X+Fblh7bMEm1jKoH
b2ccsJnkWmjWmHw41nHGNUmwSbd7vxBT4jPyArEeAKm6OSyjMoxRZBAoKEt7nbMEDEqmapy8j0yd
W2cz71m9j1JivjND+fMEWOXgJWVfYiM7R/TiTj8IaP6+znGs1BTpSJoPlAjEcKybgq76ZMeAVAYj
QbWonze5BwmmfDutDBR0bugqiC1zZOfSp3uLz+qWhgbtER2Jett3Afou/KIe/l7+UTrZM1Zf3och
1CFDXeZHU1NKHDLfPtVBPpYBjBHUy2OyiTyciQBPywaGum10acQjjlCF348KSPJkv5JNH/73YaTK
VKxs5eEkRfkCnUPeqPCQpVF/2qK8XGhf8yqyg4i8LOxc19bb6hfp9BXIWbMJtKVsBEMMf4KryMlU
yXSUddGRtQBGRALo/FZRWhOazLD4MkX6ULrsrpfZ6ievAM6rN+pBqMY5w4VzIoNnncBdJ8TBs1Mc
bhQmLuxH2x+J5G7V3ofQPARCfuGSbhf7vyqBjSDVIo8S4MtBzVhECCEoPt+F6AYyJYTnOCPSEs7a
M+LIgUGNfMyCHbFwS2+c9EO8PXmKQFDpY5wj1tXahZuC15gtMj/d/URTR4540i2QexsXDA68AuXo
2VsiphKTAzGy7PurbpaarF2N3RyXJZB62ufHpIe/4uExU6k/sDxm8XI1/APUkGgt3+zu63AYMJ7C
yphayD8lkyroTfy5JzYSCxsn1OSSawt8Hnn38H6JRf1AyU2+bIZui3EqJzgPlQ/bjhpT+AAHZcCJ
dkWaBNCu0zMsRhLUmyFcgCeKkcXQxLg/6unLajJSJiCvpcIEfHCz9a6MYfg0m2HXAPhFHz1cAbyo
sCIqdgsUi0OCFBoZSHynfzYYhrC8gu6+bsJWMZFO8PbrrkCCPJrQ2kYLecThF2XAVkh/AYoRBcPm
AH45qUBxhXeEAuDBMzlAcfyAGtz0uizE/X/lI0soIG5yIL/WpaQr11LvKqiKwPCzEmplK+ZGTOet
kvzznmlykF8jFqK8vxdBmV/DHXAf9LETf2HXG/yLxVFAD0wwzD0KlB1Pd3Vvrwe1rnziPkl+yM64
C9Jcip24rKrLelV6LwG15DUhrH6HHnL79hbkH02/VzzaYYpajZpyh637RF4UGIW/tZaQuwOqUQc9
I8nWjmnzzI3r7kqXi87BUdtKA/N8NPRSBeSxKhh2EEh4fUgEm71tjl6Dh7UnjljEU501TGz1y4RA
m6GFGdUQtJhnjpsJdY5mFYfc60zyB7yGwXqGZfRn8JKfYDELRYFcHtF9GzlAQkBjiz0qeu8si2KI
2AM6YOwOxuVV1wdFDPb2rAoPgyxpas7uPpA5L5OPv6ozcpQcIvm5Ba2AkFDMA9v7PBstIB6ffVCu
Kr3fDCGbEuc6Ismo3fywEiMDth/5mmsadnV8nmm3crOubAWURGoK3LiZsHm8PPoQRfA88Mo23yK4
BmXbjfjETxlJ1iRBKYnLtva6X/X825+gC1SMoPFTOX+RJR/3DW3yQLaCP/jpHpVDvqfJHSKiEPWH
cMpu5RrnwZpHXYMlj7clT1hbaUDk4jbkMIig0BBTtQUealft9WPkoA7jikQN53FvU3dPP7DHBsAy
ZWq+nUy1VfYMZ3fGGF6M5vQLiDx+6heywBoWQnb2hdh4Pfa3tg26erCUXWocTnjNlRHyI16Mkd5z
b/furysvDisV0gJux+mI9ht8wvxjKRZxZ+dLoPrJZdXzQy0E8VyC183xYQxKIUAVsGUWe/l08lOD
kV33uR6jWKdwi4LZclGGMHYnQj4Gdj6Mo0Mvp7ydtAwOL1+vjmWkcyk/uLoTKGku3rWzOTYAD98r
yiqNe4e8QmVpw8BRjp5CtyzMyF10eozd7uFs0OPoclk/4Io3MzyAMpABtG1KdozBWm3sHNohn/zM
wa4wcYk3RvZEgvkBgM/DTXYnP/onXITztRdW4Y9pZzmgxaSma5y80BjagrGbf68PLqMXTvBI+Rjc
a99v7k9m2gRekpcpjNpbZKJyATff8BVgs+blsu4mCBCVUHMG75Y7JfbF7a69xoYRZ1+6Iq0OZnyx
gzVYzw9OtYsD0BrWGlpZZgI8V8rwiSY/fcR+YrWgetQH2t7Vlr0WSqwOkiP6e2GXP8RvVCfrvvPM
VhwvzrBPPz/EvHf31jvgIrWISOmfQQr2WM3gcwtwu2t+WLdmepRpwLcyVuTFry33CmBUsRlzl0kF
Njn2tQUovzvnbbGd0Xhz39zp/d/eYfqnktKcVMt8NGN6ppeRhGmwtugWjK0NwgXVFbDn5abqCORw
wnknDjtS0YUZrCJPbjGVE3sf6zt+G09pxlCMcBCUyE/ytEC3QHn+6aMhbuiUmQFrKyfFipyXtu38
hi/6rrSaHWw2U6dRkslsGzkh8li5aXWeZpGglfceU/aGti3hIagaht+4PJnxOYcFXoVt4yHBwJes
2AKsSlY6JtnUPl1YkngNo5iExENXnPR0w4OG9QFYab8EfgWoVEMkth6spNM5FuZnAyKU+1x4n0FM
aI6pS2xWrd20CXHoXpadAtn+0J/VsERmLRCublYu9hJyA8rC5vY3Yeu5NLBzvXQAAcwurbU7pT5z
g8ifz7YKPLVUS24OPpu8VicwWUQcAV3206wRm2+fGBSd7H4/MfKcLp2bL9bhpUAN8/cTpgAYGiYh
i99HhFw5BqSrFdf2o4DmZQFfBofG5LnWyhDfKEJ7izMM33soRZ8FWZTXl3bUxNCDP14LDsTVY8vK
WxnQdyba0XSSWp1sekI8aSTzEnNLwB6ElH6WpEnNeH5wQIVX7eDwUujk8Yi7jUaX26xX8tXYn+bK
7WbxrOQ1huT97DRZlbnEoHZ2ccACCzv8raVfi8Zz276DqQlFJSw13MQk0+xoxweP3QromN/9OpeY
8M0WsUMe94fMv7roWstiIbdcQU2Eq1hX8QWnDHEOoxAc52zuN612tDZw/K7LPDx6ES4r6xSVNx4H
4IY0EHSyjXJOUFBczqbIX+MdN7dvfyngfWPk4uGxJYwzK75YfCctaFZ+Fd2sePywg4f9zu4A6p1R
Cn+uzXdyS3RKdXEzMxGK6MPkPaFpXF00UutAFpgYFMpOEr2+0X5sSdQOJxuDBQSoseeMoiZXSjDD
cLXPpm4LWSITwAZVrs5VgkEmgwqJUAkmc4ExPB7/J1/sSqfuKyeYmcaHd6LDw7WSZhR+uDkvqahq
WSmTBPGUIFxpfmgjC8Sl0dN52qioKXhZ4QrzbNsUzxGT75hxN0fXfUvB5T/raXcTmWC4BDOy0L0H
c0laoES40XtzsPVR28Gk+5ZMABU+vhD/JjJF8CjJ27i3hxFlouUJimOyi8LEuwUpuvEkfAKe6cwc
AMiFY9qqDmRTTfQHrc7XwrrwhosKX+npEaZ03xEJI7qdneLDtYckfJR4/1PXbsR1zhaP7/9bWczp
uH0J3vN613mdfLcTVGeev+f1oFLzB/+pOfBEnRGBWYS0w3p1wF6vVzzanIUK6OGQhc4j7HzsKz00
fae3W9YP/GAm+7+Y43NOF5KVsM+C+I0ElXL24SSy4GcN6TO6ylX5Yb9IuBDMU4yHsLI/YlVb6PFb
49upfAeU8dtPH+SMEqgiy+0Bwd6aPlwSlC47SK8SOuhfPWBwJBm2e/Wu+k9YNdpcNyzolQMs+DNY
qovZntcxTz/1nxS/GsUsV8ZGtbGXiJjHr30MQJSyRUguUOcYA7oimvUWbJxYiYwUChjbxcU1TbJW
jRhCjnmVDgqq+2c/snLuBx72OFt/YtRc0hWNY/94a7SEpZ/JsUeY3z1109i4KCSAUfnTSQHk5Z1/
2bwPgUKMMwDJT4kcPkVsDHubLdCDL58rUFbtWqXCh+RYiL4idp8L/HyZgTn7oO5RxJKWF8leZO4S
xNnMjuVQ67L2V3mvY1hM64ciqiIh52rEdoz0h6DqQrJx6y9LflH0025Y8C58G7IjLqGTQZl6RkE/
vzh1/5T8fdiH6rO9Tcdi3eWVFqynUMOe48csi5PfG5tFuuocbSqhjU2JJ9dBq+WGwotpjywCGp8W
4Z3o8KAMRmuuzvkHYZbaSC6hoIBwb6ZhpDB8e+761FTza3l4lJeIMUcwAVSe3udET6B0mnzPtIOW
gidw9JfbAUyn+KnI2iRdoioUeMyP5sYtMulnR/5k7NShwCjKeYf1G7ODnRLak04lYbS/B8Uzu/s8
pcF/fLlztl/BTofcuKcicihs+xVZ62JSjFcHdA5kv5qGxyuhEi8XukU70FWA0KcpniVT6qAjAdm5
4pmE8wOqd+URs8Q5D9vN/Ijv2eJ1thEnTo6TGP2gZeUXoE/Unxw/+urYMOJovji5zVjr7pfWBMGl
NmR+2a+L1EhSQtlX9It2BhY9MaBeQVgbYG7KmxWl/v9TjYfAUPpBq3PRrRskexPqiK7pNlED6x28
5l/EZZP0OkAgurkE5GE9z3VMaQuUdITkagAxhyGFD1P3qfn4rMBHk6Y55wxjy73pywHCNwmNtRdM
9ayJLWgBDok6JU4IuYrpkZ2JqJgb8PNJCtciYNFbu5B9IhtncwYawq8RUJ3luuXQo4FyGphgccNX
49abJ4xccwElsN/Nyjoe29P387d/aeIuVNezaf2e7ZY0TgqU32ggHcDMKSJOqUGFst7oXDuFqfq3
MEhk+wpjiJxYGxF+bh+aEcEhMJLBzC1ynt0mvLe4CtcC/RcfHkZCC5rUCd+wYluZcXgdK/SkZ5uQ
C6SjJcBFYJBjcy0fop+gicc7WkjGcRBLJj2q4UXylXWdWLwrY9zxNh8LGmCcuLZIrbrh+d06dcvK
JUDRH1Z6h+8TNa2R5mMzwJKsRNRcDww3LsLUtLHHfhIBE+yDrKpdNq4vlzph1MUlEqvRi14yqaAs
zr9uZISo+mD1q6VxbnfahiJ+3FQEwEYjehrNZ+Uh6AEVoP5TOcil3I5hxQfB/EpQ5GczHDXlrG35
TC2QK8qZbnSap7jY9bnTcg+e0cMih2IjPQbPDtlTqdruoIwB5HhVzhwprwz0LcRSL9+SqbCMNnqB
Cd0IjqcYkA7lt1Gx5A1Kj+qUELEh0Jq38sDg/Njqo+qLtCo3yl12c+cv9L8wZ2W+24V3IWu1+eIN
us7qUvYN1R8DYUrhH0SKJx+0dVBgBMNDZp3Isgdout7m1zDV59iMHxnBWpbStu5tLWvFwU8yYedY
C9J44P5/0HkalveOrKm4PcGGYgawji0h6DiL/h6nGxuotZ7dCbnPpke+nb87MyKWdx/K7EQgTa05
FETZStCYADZALy+7LAzGYMi3egzi+Ryr8FYV/XgILkCctYOIYN+Vx54mD3CiWdNE+CqqSmtJYUth
cxPlfuyg8mdxopZRNUCzsuA/qkA8Ds032cfGz2Lrkw+xuTkY4C4sBgP9Clrkzo724sQUWchgtjGM
u38tIKPCo+E3t2mCQBwxtQWUzZtiONFDWNUy4vVP7c1ctx58sXQXw0YuruKVNsHnLOYB5LwupjJT
CrPQ+IrWThz90blsWiX65Prg2M5Id20Z7gXCtWm5eRzAjswThWk92heL4MfRNlBR8JtWqCDPi/IL
qeGKFF7T9ORENCPglbQqyX/MIAstfRx48lMDmHuh4J4KeX3XpGFXrUdwjMnqYQWesSYPZgAUpES1
BGpuYTLCpktqwMX4K7efrJIbQ2dJ7tgD3AkQD0+yH9l1cQwcjSTSM+j/R0t+P/wR8CZ0GO8gcD6/
Fwxa2/+SAas+4NMuN/5+73Oxm57ykeVXZGEkyUCf0fwn1JPKq14Iwwh3s+f2TUhsl7yIyrUPFCYx
mosth5XQKgTqSOscLE2LAs8tLD6AB4V8ckBW2TSWP9yYfi7+1cWSYI4Xe538qzh5E84RUtodWJfi
3DOoj8TmET9IIHsK1HNWdWiQHp3w+5KhRE2dUZFgVCReSixywK5ZitJ6Bwe+FZ/CqXD7Hy7PlQnz
vhl5UR/ydIlOcSPQqOIC5TtM9OUaDL6/OGmj3MKhSWltCOMteaxc6ZnjaSyDX9Z4i3UaN4HYglns
Lz393cGxFyezq2hf7g19PMl9v2MNRAD7yOY3CYqfkOGkzwKrfj2cEcx+hmh4h0S1M9GH7gzGq74u
xufXQtaWxy1MScS2iiqKtK7Zk9kASmm5YeIDlqQgOjrr77/Qf2yRP0kzwc8/18bhZuED3SCXExHf
qVuHuCLGz/H7no5Ap49zlPmgDc4mXi0ETk+TvyFlguSwBofGDmaGMeUDXXDg5DuEKVgzLRgSYqS7
dCXfGbi3ARAF3nnj3sxnjIUrwNUXkhOuEc6zUQWiClfSeez8agsLavqu3JwhwLm+YedTcR7eMlr4
PVvJ4SWjNZOgQUF1Jw7blotPz+9jEojRGSyRM5a9GOwRZrnJumEemIzS1MKFEECM48UhvlCL8+hT
q8agKdUlazVu1dzLZ2PaRXcd9l/SuUMuTz3jWXYczvbnWbn4dufspT8uNg1wVios6B5+nbWZUdT0
+2b/hD34l+nJbTgZbbPpw/wxRpKQJhgqsMp46bkaYuyr3FAgYNHrYqcUnefGZydPnkksdtRKhbwe
iwwbN+PnA+5kuSEfRBvtcEn4YmrpwyRM3nzdQnfExZaWX+oYbGwCqdE7fi52b77jiNsHXNyD0Xtl
8E2RQnSJePUKrh3qw8ZRBKrD9EYtul8o/+S7O7cHwkF4dTHrCRG0Mqaimq8pqNSgQSb324uY8KLY
3+DSLkAM8Y/fdWBKiAsRn1PNYljxZ515cjXuTDDB9OhdRZ8Jtte5C1y/EnmxO0Gyhv8rPMZEcG4+
OLmfI9BQOEwvkqQzijagSiX8ISVScE1cyof4fFhb73c78tEJQsHeDmgZU3zBEVEPARHW3IPBGyjh
pqV1DXhmwT9jqNesef3OmCAzNV5i8lPQOMLYIcNfSsPVBFbVpCywUp5jtNa9Qf8AdffMTrCM8R/2
Z+fhpRl8QVTXbQFELv+IMtVm+6vitGaNRUUgpJHM4JtIcx3+mLiIMQAX5HojFxqz4renS7RKG4It
d0TYLLdjxm+iM99J1spA8xMuG6R2+gJ4IZF6mHrl3YMbnG0P7Opg8zU8uBF3y4WJl0PnHzY6BZg3
9MDs/whtoYyLhQ8NsGotn5kgr0yCEmQj2Gj1qXgfo6eZ0ujImcqi0crPsE5yNLFAIquCigsQFGsu
IoWgk9/y7mKtNv+CeD4lYHDDkKQeeqQN3Z1gaagdnFVdkcFGbJJLz7yD0HEPxs7LGgDapnnUSod2
J6E6IPsjIDPKEhFpCoaR8lZ+kF1lGmmkLLP9ap6oPdW3LJVpyu6xaz8CAyiO4TNAAkQLRzCMWFuD
hB2YE35KYWSy6xCdyY2oVOBopQw74ipWJOqGhX1zRK3uUNXIurtMkneiLgmuz2Tg6F9jCoriDMTa
wuEEBd+FkwcrrKGZhb1nWeTFwrtQdxPOcB6ZBWz8aEANhqsyS4gHj4EHUKICy9yCXNKVD9k5tDbc
OgPRKc4bBeMA1osi4r3P2tyRBCFIbYbgShjRCXxmbDwUvjtNhmBvHF68VYxVrpX8FvYkIK3w6Bxh
zLZ8IzWFFpeEJU32yQvig4wC2+5qwgCTdAoP6+za+09PEqBXqdk2zyKwa5qRih31719gTq7EQMm5
Ay4jVi7yBeI1h8Dpf0m1qCag+9NiR5C8pLSpquKzXooHZ1dkiTXBAK0UTH9aGDvQfmYm973YO1Tb
BY8oBBOcmHsk+EwDdaK25MVyhPjcMkyPJtkkng99fXRcVG97YtvkhmLrZyMPXckAt0GGA28GDF7m
JJ+Azg9ahshqmKJSR0KmbDTXmEgdZOfbQlAWUuPa/1ETafqeCVda0ujSy7utkSUPkywD3AkbJNvU
0WkPgH9ZJMxjz4a3GF7cT5sjmsBywOb0vuSEhOQZcVYST8lBGQcGp1NJ7D4pvXSEtDTDPFjj6gac
gsF1t4sG+/fIWrZml0wEuwKbD/XnzYXoOqUjAtLTZS3ZFjRKkMVBbYNqBKMYsLCdNAEkepzNbft8
sXkXUcAHcw5vElS+erSsVHOkk0K9RLA/OrYcCsNT6mCweQsRg7e8Zoi0Z8vzAbj7GtsRH1WKIG4w
wcK9mpntuerFVfGZqnlq6FbDsVmP2xBqBV2Jmnx/0g6LLnjl/ReVsFoVuFsv9uPVYBHLyle/FUqH
q7qg9ws1L4MWPvNYZVJR5rAjn+l/girBuXEBVZu15H/MGfzCVGb1g8Q97xkQLEZWZ3zSXHJ2m0Rw
NxLFFL5opU0RXL1i19AMMmslk0t2RR/gc3nQvwPmpp+cB7FfWHvkI79csjShkyHeEmiETVEgIrq1
FyL4g6ICA59z8Rq5M62NuMmu219cOEtmnBUdIBeGuxANV3HffIXFAexL+0c40ozXjHBzpbte7yEU
a60DcMdhkX417X3pidgzqCD053TQy99d/XmuLhpzIplXPMVdnp37i5w5sDc2DSD0mI03o2fyeTAZ
OPxFvRDulSrSbGDs1c5y9TrhCtzRm86QTUUOroW5z6NaJBeFrlkYcYWBYJklJGctgataWHQnUI5a
wAPDpIedtaGXSJ16EtPpuJZmkDDy7ylhtTS17HVt2Zc8RFwtOKYDCRXv/BtQuo2nKbH5Gcl5lAcZ
GME2Un1QPIJWiIYRbmUEgKxaqT2jHRcxOAhoJQkydxITqVA3NxV3l4nd4/iZ7aaDR7WMKf0quzAg
Zl5R32aoZfB0J/eOgLtabVbdIH9KTlmdzK+4P3FV4lG5eCyiPJYfSov7+svF9idzs2HZjzGdPjNq
39SGHhbbwLprbxNo7DhdFHJBNgsqyfqZEhLaP79k6RwyYF04/t7CEKpOzvV9XopJS6OKGzlTJsNA
OuZO6b3+bncciGYz+ed5qlnFBp+H3QGrULDTiNE04Bsm6PmR9ge3r1IXu/bArTknJfwzMS7lMNRo
MW0ZpsxuqJfwebbXoqXzj+79U7egQSbkAz7sh6FOnM0Pu/UtOm2SwNg3Rvmsgs/3BgfcOoKpZYiH
eyNVNd0fHU+JMGZ9C1k9L98swTznTt9MSYxHve3NEPN7zh4ihaxq05rCQlB6zF/kTC34FbQBezgf
VhQCPeiGGjcQ3IKusZBn3wxkvC4+uvKoiTU+dtrjay3qy8O1Flv00chpj0e8MvIyuLsrQIfF80G7
5BDC9L8e0N5Ik40CNg9+V7qJyOiqstQe9VaHy05tAidT7SYwbGQqNDVrz9ZUoOr8douWEd5SoKJ+
OStBnb0Y8N20/eElIaQs+efoudT4eLcv/NFk+iZnrN97CaovIk/AZA24m78wDdADqNwfLtEAh5R6
EEWvSQ5PVs0UAYcCnuggZU3KU5kPZX9tAZLaA5Eh6fXMvUeHXxxix5eH0mrW46bNKbO/pj79ZAJn
EKr6PFUlo8yHcmBEBR2lRDXfNRPJCTa45vTwm76PbXz766leY4864pGJsQdH9Asmdlb7QRLNaks+
87hLUjQNjPihP5xE8urdQpU+gnLWktg5kb5UBl8PFW+gHMVtUbw7ieGeLUNrJ72Er7VZpw/VjybF
CdreNGdevZg2VecggvCp+nQ+czqRytSdhYlO8vSELQDqNdBkR8bsDUtPiqnogYqaSNNBk8A/izX2
K4Md/zKLNtfqXiqjnXudQnqDVKF76zBCFqtU6kLDO4UmfzQO3xgCX84H1tUKcwezyRIH4exA9L5t
/BcIz/Ecbknp/98JoZfoaFx06+1MXLVryaWS7EZccrEjbDo8bxn/Fs9zpcO2UMzzr4kQwBuUQV5D
AQJ6/NalFqkAIppOIQlcYleRtEbTn7PUQGir49shx9hpHu3apyhwhb8wtvD/Csp69H9TWbKw1vLS
pbsUHZft6jqCtdjODtVJ3yHo55Gd8VoWekjZ6SOdcC2LdsqIltCHvcCZmnAYK99b4J3AWay9vl3+
okZwjz3rMfK13i6cBaXfbpVi6ofIryKTuv2/0o0/McmOwLO0koU88GQUY3Kaxzdu4e3eAgAcauHp
ulDPS7smWIIq+PNPeHoN6+p6XDGHv6tRnbk3WrxlCqIt3hf1IEXDYWyr+9AHSLGGOvXiH447hiva
bP2aw5dgJ4/cGeKcPKOZ5JKRz+QCpp2HjxM/8oQk6vk1vX9Z7UpU6TngNKBn9kplx4ECQHfpROrm
SMOAnrbNPOo0tH9/Dp4c+Ix9PmhcBJPBD74/GTSTVPs9eUZ9YDn68voQdOUaRDWR4a4tKN+aFJg2
2gGjz8I/LiwCIKIUzCutGa16zlSO3yco5BBkFFLYhRYkRJc2z12BrBsV2abPP9ddd3E1KIP8AvyP
TgDTGz/xS7QuPuajsF5z98MpWAa6yGDrbwPAlDlnAkE9T9F8PnLABAfPGVSc8CIn40O0XGuRRo0k
dXkzWYA47h0u25p34KkQqV7x9dshK1n15Oq0pcNQzxVhFA+StW6AUtClKSJw32WBaSGqymVPoLLh
QVp8mzRPrizIbaH9+UTC7anGoAi6hGEYT7K5d+ScFUnuXyqaRkXqpYBxCUNi8ofC+DZY7+g9oQvN
FNVdZTUW4no/S1u/VLEOS5Ncoa46P4xT1TS4WcJVzx/OqoH8+QE1LgZFizELTKmhTle/z7ur70S0
yhAzhfABzklS8w2W5pp8gr61d/2qXF0cXtrY5tgAddClWoCcGUTYfhDGXQ213l1KCFCeY2GvXrby
Fa3yihjM3inREC71WK1p0TEEEKEP38HmV41CLsiUie6LPKdgAlodasMf0/D5DFkJXL4lOQNCZDDy
p8nogbreV9hG8zpuhCqrQa7/5qRpRO55FHtVyfxqMRX8NaB7Z79BdGpBaYXHWLETc/DRB/wSpvoF
B+cFgLCiWU8ImtXQ1uN5FVcfsZTLPTZOlblUPHbqkXT0BzHNhdPItiN0Z3cBnwf4lTWcEx/8HwSg
W5RJigncAX+HxnE6quFiJ6UM8zzge9YdOGnp0RSksnWI2Tr5D9YtsJQI9HUaYvgV8LlrkAGoWQmH
17iewW3ZyiEONup+64ak2CueQHzeJrCXtrRqk+Ko6Vjj4Keuzn52vjisPIfYEco6St337zDIlqof
6v14tR+XHC0Q8zfUizgMMwtJlofuCw9t17q4F4oz/pKmGW61V3zifOz5aEoY21svginihCQScu3W
FwiqP4yVT6BM2M4AVHwodA98fV+hLe/1gduTqMshOTilZENAeyj46GHBnBKecTagtJCt10N24Aor
4h8mRfFQXh+fSFvuiAY+dPs7hBO1DREkzLFU/TRlbX+ZxwMTxGEmAOry9CgiRpUItukxc1DNL8wc
vvC4Ru4BchlSR8FW7DtKgGdiHegkqdgk+zJv2R852/Yy2iMPjEgZ4Fhf4hojMEJFInlhSFnC5Uli
LiQYMhIr6pvnGo8CUEkK6HMtcdRI/PYmtAgJBWeS/PCLSr8DnG/IH3MP1BW/RyvbfbLdpiNzhmKm
lwRKd33BwCc/0XjAopFlYvTt1z2w9RzmRxzgwqP9zRQNQ56BWkZAL2MjTLruxRZhjhKtw+sGiuwA
VbAfBKntnv3rypv+LxC5LNaJRfpzvrYXb5tfZvghxeSXQMa05jzpBtmzzy+88FIcokUQY0bLSIIa
KaGCT9f7xhqlPbUfOmu6/kTEmIDx2ZxkSxJoKM9nfFxciV5z9zBpqpLHH/e/THaPBcDXYccRzTOU
cEa3vq4bX3zua+hwFHhI52FQEdDs6LMMKvhg/nP7Zp64pZ9LwKFZ3ymsWPeExgt016DLN9wnDjkL
2RtOzWkQiryuf4q9DJJWe+/UTITi1rJhsVwPy7DKAUxo8rWCQt47O3Ef5s5rRRFFRHIlyIS0FlEh
w1pgC0+5Kpgf3Q2JFmH/YV8iH9rC9sid7FyaNNFIuq4/thFfIdb5Uw1USKEibAgA8M1Fd4khLooX
gzMwQCVqMvH141zpZtBxn9RKbKYL+wS34TWxInuGICvameQ7XL9Nymzbi1fa6k+0SsZRKT/3Q53r
oLmxDnFu5584/GOPzC9VYifIYZ0hfYoQmTNFwhmYgzcngUdVnNFYbvocJkL8aJpBYZhSzcDtnZAz
MPzlkQemfvuFmOU2DzKRRcj8Q+f+p0LKiyEBBd7AdkomNyKSiLEChfdrcXdpkMWtvhyCdr9UsnZZ
qQfviiAlJDkEK4CE5gdJNFPZMR/bGVLSAk7cPlhCsgS3VQJR4fcatQyToBBG7L2FoDSXfKiIvQsm
1+J1guW0AzcpQxcgh8WTYW01Cyh//RHGMVhtvngAU093l2kCLJtz0HuIpwQSLivTU8/smLRLnM3z
F1FRnWAPt7J7tn6ARgiT/cqtsgaJ+ILd/Uit4NjY6x1CVebQuTNLtp5qfq7hYEo7usSGnJhWAf29
LZrpNu2bKevsDbTKDsik79n5DJy4Fy4M9u/UM+L6H4Eo8XL9l1JSBwD5T+Irdajaq1DI2FkzLiza
lCTYQfLRTA/xm9Aod0Vj43MbZs1ozetzOwJUHqcYj+lDEeW39P7db5x4qo2eV/6ojDDF542MrQyG
WjiCd2GVGZp2jXLEBWEHEi0Dyly3PBHB29hdFSNS/EoKM7qyhxme+XFZX4mxe86xr5K0KhCmQ9dI
wKnORdxE56dmUt+7ZUKG1cngp4Z0tTj+H6XrNlElybUWYwAtoMaozwnoB5tqqYPf42Fesw6TsV7F
xbVpXK/o4/ylolgctdgocRsQqEVRmtXEzRJtrTejNfCSR0ql7DtqzKEL1rG8RUF6w+PM5J6UJLyV
Q1bYcXiaenUK2JekLlz2KccL5W+NnXa4dlvftdMTYia8eQVKP+56jxvT2rK6lkZts2hogeLPN8jE
tj5tsqlLxTRsNDnNi7Vvirj75Sh9WiQr6eiLYe1j2acIgj7d5adfaQaexVJdukokPoQnC85elxC6
nkEOOkNcP3/QMVX6hQ7Xze6u7lmnGOWfAmvMoUl1hsJ43QTeiTLuQYJ30YmKQxxpoY98NYwkh+sT
jLIRJcgCaO6VXt8B52oitbpvbIGarHcjkHSSryc41KjlSJDZvdpT8C93F4DymjC3q9fwxqWl3Xkr
/4upkwEy/QYgwd7EpgGqSN8fuqwlcUEk9lPkETlfaw7ZwI2CFo7i7ISz7/f1gQDVvNhzpdGZLB8U
YKCNjmCGbuzh/0jxWENim6Hhh3ghVDDcm4ZKpwW7L8q9ZkZdZ2SLPbQNBNbSSGPMZW3X3a1wbEoR
Blma0vXNOJ7cAz9w/FdKDLaHODLmTwGPl5corGRZTqE2RoVMtyoADfYTdrfuP5ZDYOuMkf4mzSB8
+XLa6a8maJtzl0xxRU6evlu9xbOh110+O1OUbnOqx5u0K2zODjNjMkMTjIGlJ76d4kSHMXZ85NTG
cpx4kJCvgZBrn7G1Z+H7pgIWliTEhxDozvmVFRLXEO8hI6garbc2rQ3J4E9ikpXjiHcr/ceCqAVy
Napu95bSuV/03MXecB3leinixH3dB1LRz3AkaPEz/Z7oRWXbFrYMo412tDIMkVXTey0uUboSPZTZ
I0DbmyPtdOez/729HbWWbZRkGmrzDKiXS0CKVTnUgIqxZ06Jy8OUxCBIYD3O0vXYrmK+wXM2A7M1
D9GGW4URuBq9M1ZB9XF/0tE+N1SmP7dmHUq7jh4X3QvaVSE9odwDK6ncYTPutW3Oqxm0IHzwnSkt
CB55RcoIsylyzFUSaeoxYsIMcKaaUtCgnL17ilcX6F2wsk2r+Kku8redU3T211SUZN8+7D27R9m1
lHDMfBEwF+/AotWtQJtIicv0G9kZevJviv/urYE+x8w5wymN8Cu04wAbd6Q91FxuAYPZrE7NNkRR
DEll2+i+mXmUtCrK3FFR0Vo2GO+qRNsUBnzDf97+cDi0JgvBPD5iW6E1AWfMR1q8dB4/Wf2hKEnC
C7aWI0EPDO0EtsfEu6ztEbVdNw+qfjgII7aKrM/Ofq3x8zM+ItjIGdypn5ygzH9/ucf3foLg/cbz
ACam6zdWmHxWV7pSNpLKhA0xg33MAMv7z1KFdGJylClTy2qIT5MrKSWB83HsJC92Z+nSwkBfFCfp
SSC/ke1KQNp3cxGi3ZnBsctzcQDeHfnLpi1PVoQfN7KfDc1vsgGBNMjiW8aFQyHyqw3902Z3jHCq
0TVbLYC755JPknbWzhfIa/eUQy1iwjoQCEVe2pV3HDY6v+QcV4ENhPhARo6OaFPxy/2I8PlM99+C
GiXmFwX+epzoBKCZ9i8kVsez+BtuQAXfZ2gTfG5HZY3FOqj3+9ZPk6h0DuveQmCLQv59Xo0OIk5P
qhORJs+f+UA5IZU+ZGkxvK09E5SqQ57jn33BriByAPYU/QNmkU46OI5TXJtbOUvjyBfYXXDb86Ah
Qp/3t3olO4MCc2cBhcjcHC62AImHDGWnYDyMNVCigpoma0hV4YEjF0NeTF/ywX5IodN7M3JvJwNm
brGIKId96Npc/LjH6CvTkSBuIBoNsAsbUT9PaRXPoq9rZwmETqPJCRRSbbnm/DYA44dF+n41IWPm
rVlFl7LTv6HdykSjH0jaZRI93jUuscT/5azZOmUgiiCk+I2SBx6vWQh95wh0E28nZ+rX9wqSbTws
+K60gn04y7fI6xqsYYQCzfo4zIv5nLjpFjAwCYgjOi8vCMkvkJlosLICYRJKha0d8zSG4OpWo/jU
oDhVopRhOxiPngRbvcHFGKRCtc3x6AkrxjC5sAO/1V54NwwHHCgcxzYeMRRuOmkgOMv/XTNw9BQf
ZP56Z7N5djzBrvvAlAXa9h50SycE5UYvLdZ9TiSStO2UPXtKeLMhi+Tq1BHqnRdMkwbagbFxCRbT
mqy8/AppOHLM+7fyXzWX3ZwC3dOZNl3hkn6gCDBNwbjtzAL9OaOsTUT4hhh67yWDs2jYPXveVVAK
ny1+wlp4wjNJav/284hRzAou1hPcAGT8Zrjqm0tB3N5Cr8HOhEgXjzeRwXlMeb+neP7cAKOzG2UQ
eYvIGHgjwFzA5L9Vn8q+kq7HvDBSA7IlrmPIlKJyYe1qqf+BIn0tRuD5+14+h75KpUeBquZZSMqa
FxgsI5pocyeVQxLV+8pm7ZsMg0pEt2Cjnz/KvjQtKC8Og5chqVPokAIXzjr09aSWdDA/9ySrs3Mk
sAhm6LdNGfjCTrWFmy7unjd2pJG+OJZjYHBg1SPQo4Y4O/oYdoNXzrTch+IOBMWHMVxVmixCeQRG
CD8S1XOqrKD1NaNtf3IwK6x1LRTJhFksdyKuHdtL9TIoHym3H/zcVbKwEGSEUikfYGemIF85Fl47
/DUTvC56Al+FA2PvnQ8Dj2sZ+Yk+wsOf6QvGF6M65S/twKqvfO2tlVKalk5kSh+Cq/VVvStsz1P9
UL+dJG9Ju++pJbRDQH7fyeUf9PXRIQo2FVfBZ36s80NSWJG9gV38cEqnS1iGTqi0vSquXpjIHv5K
RzsRRZidV74yWiV4XlzCh7MO1YTeIlkLFkk9e2auWbVY45Sra2rDcptyZg5tr/aNsYPx4LMauQwZ
9Nf2+dWcWoZFeHwVPbwuuDoEvffNqXrIiFZKTQMldbEiNU/igLwQM3TqqBhfG5qAdU6ryeeKq0N3
IvXvqmhQj7YhVLMNMmIJVw6K0LCLiZ684UCvbSYGnYMIaJkVQ4mq1XcVtLnjGMTk3mqmT4DXWc21
cEtCSI6hGmp8CrzD8tcLuy2JeTnVJ1Ot+dxPfJ2nRImy8kvXTm1WDZaCqY/uIEXFJ6ZDN1wUAdZn
VlSEVOKTJkz7HSvLW4N5Xo1EkW4FbfcwzGrzr8MQcbmhufmOWQSAMICzFsAqTlXyPZCnddnvGQZp
W74994nyO4FRdfCQe6unqlMqKQkhTVL91WkRLBg1/CI0yG18wlUtEWQGNw3n33fkO7gu0+EACmn+
e6Ungv2L5xg2kfl0VfRFmbMy0qRxOBeYKgPvGMzowscq8HiEXJGnASn3kq4Nf8JZ1X3iO/aBvKaN
jIBTyf7IufXpW2C9wnzIehrMCj7wDgN/oVfzeXlIj8L4An/c9tw/rJ8CN1SBzT04IcDHXbVjCp+z
8j93F985XHuoEyqNPn3CR8qOV5PtJ6sSlaiPMpywqrKG+xy/GnHfNBFohP5sm5SmNxS+0XJEB3RS
WQ10Pv+mlJo3NmWVDmD/3hYIn000TpD1sy3Gl3L6cZbF6B+3YNId0XpddT8p4jcGpnbuzV02c0S3
nbqyfR4MFClbKeQkmsLymuqcNrRNZevj1rukTeqKtJVpjHPfaP71+JAaDcpMSlfTHZcm6rIpZtOW
i926s4jk5CGLb0AHjTX4kEK+m+Nk0Q+OWtBUhoFCovrdXTkx9KgM6D1jm/GRBbW6UaJHOI8WmlJv
8d2drRxSfg+YxwJyit6lnqI1r7gl1O937cxnqD66/RFWH2aLxy7czH2tmCXnUlzA5IQOD1wXLIdn
WI6mh236KSUlpVbKkGr3CsemVlB1ZpKbZSTtel+EjdOtmUwnLsZ80bcr5/7vB7/jS1TmKIOF9kYH
C+0u+mBs0AxqMg/cyLG7SN4TCUY1QC9VebUDENU8vtpn6dCkAoIe/kHDCAZhBE2z3iG8fryOTVYl
6wgnJ4LAaQJPlkcBLIsMH8/AuhqEV97j5Sg2kRo8Tfap3ciysBxYV9YkNru3OLKLLt1rv3JrGgN5
xAOP3oxQdcAsgM0mw513/WqfZc7yEnr9SOUY04KpS+YJvFeyzm+EKr3//LE026DDIDTOSBnrZn46
qwskFsGLIeDuqCsuOqBeoU9SKYIU3iYXw/QVGCxOF2abrdX8MszUndMpaFoDOxPC6n1EbQrDFi7A
2/8f05kpFpytME7Dh1s1b6NTqV4FJmKOcOtaeJv2zhOK8SWPz9SkGSAI64OxVMtDypKPTZcMs9Ow
+QWwluXlqcFnHjfkqqfS4s8o7QUOO1IACWM/crKKkDOEs1sDHLUhzgCOJsr0pcFQdoLTbNcKdUlQ
GuZ8QtEHWP3X1BedYddCacAYWWildTHDZfL6f0Bt1uRkzEXh8NfxVHSznwSnbWt3KufUJjRNl5Tz
82T4Yq0+FaO2rVIzBcUqNq3ZqzzXbXW3aJomUhP0xzslHTXxoP6nO51NV4FiKOq01CJxhyahBV+u
afHof6d2wDVZIot1ESGlePVjoyQoH3+GWelD4PvQtnO+RSLcrZCPp70DS+aJkN4bfgeZO5P7N7oO
97atTvOnyHH8XTWYAfsCcKiXMqWMM4n7U/QM+PdNxXO/cQE74cFph9+3gbv8fYB/wOh6FXLavj80
HYHM/ijaDEOQgXaRNej9+utn8XhtP3hEoJHfP6T1+LN5QQwh+2bAdsPPGz0hZ3vL2Ou48YVGOloT
I62SRxWtUoy6gye7A1OJL1IVunNt2CQg9/nHDVPZYEV0c+snzevYjSIjOlZvlI0A1EbeJT8cMKac
5aoAu29NjzpK/0Fe0kBIyl9bEtodfcXuS+IpQ7DaOmPFtd0CuA5yeGxVQngjq862z9L2ZT1bu0Lu
Edt+xE5F1I/0OcxzcwaRrtgtUXfhLMnsXpW6TU+fhuksmHrfircNxR5e2yyQHIPY1tkaNkv0d0Ik
0LKuRifCrtCs/FDk2USAW1e3jiHR4ZANx995V/zHQ/xJJJL3RMRpXcvvoqWxdUk8Q95NcCIuV7Iv
nbCd2OuLx/JImAMI8EKBilTgczbV0F70p1rDBnPk6JQyRem2V9lF20+6fXc9ovhD4b49DIspesN2
PoqbStWJCF7DGkhvJnK1Hz30HS+648UI4kju1JUUIGNxsn67rYmYGd1O245T7loLHDVSLNozrUvK
Jh/p5sKYD4ZBYBTmc/m8kUq1SrtByiXpoHHJxkZ6Q7j7x6WxRtF01R9LfWAoQ7Q1zLRnn/C1nHl9
PJ/kTtCibsh6Z0mMTsiFdNukuC+ilKSciSJ7luBDDHoXBDRdAtkJ26yfxcOGTpHZmAyenRsPpjN/
k18qeWZeYVYCMUXi7t3cms6G46XmhZcBm09tO/df/CO1ZqOrN2FYXKEPake+D5mnAkXjuiAyePjI
s0suZ4/hMex70meSiYeKDy+lg1QOXCDDiJ3kfjjm2gVKdZAx8BIKYxeja//xfe2Osqmp5/qNtWA4
wGjJbeKmRTMH0I+qQuPELPfGNBnLhRRqJRKrBeHj5jOitvouCBCvAw6oV362WZj4dweUSVNQUyA+
BMDleDSRrlKKHRzZHfXOJVG6kgo4m+t94AymA4verYCskAauTiPjH4J0ak7wpv0+jsC1N4jr47UB
CqIUQbwc5wVLto/irkZtPkZq9+rxn8b7YZp/dZbnHV46ULjWZVxbs4AuNzNuEK9uVg3bdopBGmZI
8iMFiXoYW61z615INWTdCwWyeK+Mxa348mCudtyJ6odWpC9PJHG6I0KSujrMKBQzrxaLMMR9xXQl
n7Z6e0smGPsJXTMk2zQ08K5IVfp2NA9uG2WCnumQVb3DSl/TXeGRn2sLxr3eFES1LQousHPPipCG
lDo3YIijuFkPx+VS6cGiUk4FZlJElhkoFc/a/ZvXHA1PaXhBLFZNsEWMHE+reMqsQfYvTm5qYgy8
JHtGV2QPLdHIYMn4RDOI/0r/v6jUEaDIWb4jDjqYKzgAmbuUZG1jgk6kL1+eSJljrX+1OeTLyxt0
6M6e8ckREpx99Mxe8O79M6VlTVEXdlve0rokqwWzsICOTYZZfy+IIUESe+ASXrf/apsK+NQeTR0i
To/n/ZrRejeqgNGwpgYX+pQWWWp5WR/6owqj5p6F95DBcFR5wCLcO7uoMuhC7DbBY6e1vhCRY5tg
zT3HvU8vwCZFlTsQIxXCuTWMzKZXYztGcPBURLLOB6vBZFLXXKVqa9/TB60/W4y/UMMF7329wJJQ
koiDpeq+r40kTj9/Rk96E33K4vROk4YfZaQIaT8UxmKcVun9PpF+Svc9RlScvknhzrB6KRefiw04
g6EsXjF+Th9yPHwijJ6/xrryxmzf1veYfWnCMFR4KqKlBST4puxoa3K+BrnobEulL8YwPRe8OrXw
esXF1hifyj5/7E4thcLuFy8gczHGJc/TG7Bh64IUj8RjBIWpCO94lOv11kQOeZE2a3DIz5Lx9YPa
4oCFFVz0FJuPLNn3TSP8Q+fhhzFtaOH2Ocl0SOb0ycsWcxTyq4E4KYmc/SnGRL/kxEXEXBwJ2hhH
ZhD+hKFLoEvJ0JcyYnx0rgj8Tp3jsOcaJKnkBrtCjg6qlN+5PjzlShSG/yAxECSFGAGtQR2VWG1v
b+nBABNwEyhYfWyu70PW6Si4cP6APgOTfUYXaLpE0n4+DUyTdNl1jXDvE1lPUoAfUd+SdkNSZMX1
cbU/qujA+6EAUZBpiDI14CTzWUYhdV8dxTCSm8u1CBynjIS94XBc622ZtdsNLM5NJuncGD38m+h6
mGn5zx1Je6fYGkZ8pYINMB+sTQuXDwKD0cafC15QD97w+RtwrLMRJ6KAs0CaNfszF8XieYK6s1sS
x/Sb/uH3YCdCfNNCr1eMuNM8xlKwcI5OZZwLpebhA6k99D0D/L2Cb/zGVABGJ7q7lsDPJlQOf48u
i4dLwVurcIEABtxLLkSfdsU3NP8pOBtS1UYLnDoh2RUGkmZxPlyeHk8IUhbtrvQCfYo98E0b9n98
jgKaIVMJuBQjv05GTMXn7mCydtGr8/Q8BcW00iUniLR2gsMGcDPTC7ZuuRsXXRioSAman3fyniG7
WdfVi6JLx4eFlC4wh2yAiqOLovSca015RiC7rpBbXS1bXn6ZdCb5x7M27QGQOCtm5C8W7gpHlL1S
eY2llmvDI6gEwhOWucsL4DZoRGRO51TvRpI2QR4p2oNz6BSD1X5m9oLJiglMnIQNWuz6VwpBCcYB
ydO+KuHFIt50CLijh5PUgU3INc1pPYnvdIs9C9MAQMFF5gzDWF/gxpSnCBvX/VpkqppCfgobE10E
W6LGXFvC4lVFv3h3mgaBgfZ0+PQwbIZv51yzabQ9okEofkAVzhzkcfOxusEkV4iCqQ/o+TXg2mQI
gpOANYi3rCzUMVPYo5AvvQpWYtwAf3kOpJeV6h1I2d2CzXwnrVrSYoexGXtGYqaeCq0JP6ux2qvH
/VlhicB0NoZipPQcvjRfBANg/JEEHh9NNB0NzT+H0NdVkgpCX0Ctu7ZVTea2p3LTc4iKPMT6OM2k
vUo0/+DD1qQxZVNlbzoeWVqLLExSf3cXKF6qCi268LibgI0GJwCYAMpFydL0nNVXEkHe1CxDjKBP
3sNT5bJ+N5WDLrRWE65zd8taDzb75KHD8FGmvc1Wb3FYyaYe1OiN60pupWhS4L+kkwL9AkYKap2y
pWTH1P62cisqo3Pt8zKepZCt5nBPa9/tVUzXhLtLMUjqsFRdzxbwSAyVBevX6JLBSSz2MSeEjelm
Fgi/qhglXNxRc5fbzWvg89787zqIKX7OL+OZwXL4cCapb5krENHTtdggqIlzeaXLfU8MDtWCcpKd
36lUIQJP1eVQspAHTaMaIXKhNOko/OJkYW83EmQzsGMXGQ1H6W/s6ysWZqs0JNsPlibpVHrEbBLn
8pnGCb+wI9nwOQBPSxcHBbzLRfwWHdP6Dv5eQuqiF1Q9jyay82ztKQomrfy0vj6lTHqrc79zXGgR
jhgENthQCZSqew2JwdC2K5mQoi3pHaR7PSmVgCiD3dh5UagBmSDR6HYoohrDEW/2hGSu96U841Pz
xhd62l4reD1lD4fSVqWtRg80ZO7qZ4/yB0oIegy3nFqxHk9oEynhIkR7Ob4ThTJ8KUfX7Nh+/wY0
x2Ljn3WCH5uwPCeL375c20D5WprQq2mfBs7zWkge+8fCE4g+wqzEbZyH6oJxeQkEhNUsM3/aq53j
U8ky7u7zR5L0y4OFe8WUJS34LbeN3gq/bY2e8JY95MjtHn7EJcbbKi+3BS681xZb909EZtcNk6tA
Q7NoFp/wcClSPySBv2gCIy3F1LxDNr9kvha4CivJRQFPUNiP+tvxF70EYVRITOG969qYCBwYEbAc
qGpeKSTWACCKAptViSINPDKV5MxTUoSkB5WoTAGN5qgpLxToHHbNsZggtjM5WAXvqo6nq1ePHsHB
IddlSa0g/GgkfVIdlbRd86+oQCnbl5j6/q3Bcy3SzW5g3Kbdmc6Tbkbu0Brzl+nfyue5n7mb8xVp
wTPnj8JWAcdQasL+LOg25ipPC/J2vtpsUIjfVkkLpb2/AwH+njoO4/ezVKwgIbQDMQ6gDn3/A8H8
dkvf+VG2Xnyl7M6DChZ3ISpOuS558589cuSdCjNfGJke55368S7kzWUtk3UFAEb4H90rLd99u5xq
gKr4X+lSx+a8b+BAq9j/TlTsMo+fqd1fY/nzi1ASRWTS8tVt6JrvxxgtVUmOgJke5aWOpXQ8YtJr
2vFLWI/N11eyoVltkeUuLS7bps2Euw8smpPL5/jgLDHtp7i1voDD2+KSMbOFCRqMv23FB8jDr0Ua
dqJJ0MCdfzHdnYWWcXvJ34FnIb1N+RNp6Zhiu8QY1zpwrr/hiTkIJy3vcmTmtCYvxjfRgjcxBJbP
sosN1R3fGVwmeFtgpaPxYMfapKH0OAjLgXXM1Ho+PbPX+vAfCsd11FTZ0FARvV1t95joM0F8dKqd
atUQ1eDPdsfu1wlcdCStwNJe6zmrb4uKC6cpdWr4B3zf9F0/+Tw9zeEQtnatsX/DUZ/qEFxye/Qw
3z+MznV7Cm2p9uwPXzGyCHRE+9cDG9hMqUwRNogvz5+W3APN7JE1PyiAGZaY+iwQrZ0QIeKslUUA
tnQnERUPD7jWuaIQTwY9UOa440CTiGoffSQZT29MGK0J8K3wxGBjgwdSNyWcAnbjGO/wYJIHQPWh
ywy3Due2OpkKQlt32LXSmQFpX/ZQGLXDRzULR6k5GwWfn0x6YyzkUWsU4Ql4+l9HI0594LwUQ0/s
QtdO/V/4/CstiGemybEH+XKzFZagCV2Cccb9wAUgqfpAVi/EBq/EFsKCd7Nzux5FPgcW5kuyP8tk
EaNfwwcJ8j5KkMx1wqLHRH1yPIOPpDnOVY9JB5yRRgbCUDS89nV20QoY69yGxwfOTIiCx2pmc6Mg
7qDBB2AIqRZDcWnOh7VWweQCiiiqH2caTL5wT1m25DI8HZ0AIlQzndtv9fvYHOMpwV1v9BWQ+uiZ
8OVjZsAdHAidQROQrnzFyXsOOmvqEmvLtNkXiTsunkWly3TXO2vh4aTMQcy3FexG9snjjaWwSr9r
P5mRvkVvBcVz00mDLgH/04fkioHiXJkaz+z4hT58k8QsriGlG9jz9sdJGqlj5WJ6cSJrR4axxx7V
a6d0Au75QON9WZACcyHT9JdDf4R+lCB/f7aXCL1XhCUijHdm5Js3AJsrCpnaNclqcURO3KC0IgvT
j73onDC1Z0BXZ5W5gonANdofFRSv8Q1xDXe9+ASLc2gQQbOEpcwRXwYRmqh3YKn5d0tjAPHLWEH0
J012A/HvaR47lpL2oig8vnOzNELO9SkvY1uqKe0F+FP48BehX5AfwYpiu1rvPDGzrsXowjfcZZ7A
qNp6xNfk5kg2h0ylAXloh8rFt71+czFu8DU5RCPxqgj8MOs5nLxMnxbJzJ1NeYmUoX0djCdQ5K91
loa4ne3etScAYB0B/sOumQXCOIimwfWmR58xu0VZ8G/OSc6+vEVvLcOuFJhuvtVdGG36yboP7ghY
eY+lzwQEU4J2PEyJ+q+0gk143uegBGwWYacY5MddIdo3jvIroLIHHAnNvzFKMwMkHGflAjL3yD7c
ljgcavqZN4mPwWczfPjv1O0bxQXWc6G3R0kvYTFN5W6PVpnvs4q4cozmrTCyxo3Gfq1HxIgn1F2X
rwd/Rgra4YNpC5iufWjXENIr3z8sgCZN1w14Fep6/W92No0QmbeJNUTFs8GMAyyxnylTZS4AXuCs
Hx8iUDLyw464onkS/uGgUP86LKKhY9/l487B646Y7naeI9vCjvBqcIuJHOSZvGZLTm6XKZK6h5Pv
SdNUR42J9KdjlTXEtFSjXj668m3Gh0zIYQGte56qYAHEOaRPwZDuAoTGlzSwFHRVHr06JlPLjtRK
S4g26u1hAsCyIRjkJNtIvKQJ0rUvcJ7yzb88dOme14K7W5i9cyjqFOkWDI11/LR8p0vgJGg/1YK+
5aEBhfMDc4tWxgzzd17uI4kEbI9+Ay6JD5Ofnx+pA+QISQDGYpXxG4NlvbUj7aAsSOabktmUUpnP
9llchgx88i2W34z12pehG/S+VtlnHEwRodLMhG1LaFSkMHxCZXxMY9Cf3ZuyVN02DyZ+mKMzXW4P
3Wnf/4UkZLY+M0D4qtG5+LodabcBLpLpAoEjjXuZUfA0fj8D7jqUupQ3UMIAXtpnVF/PHqRqTe15
Azill8gsweET8SIi9XsgjH3KYXeGV4Hg4uK/J0KHO4zVrIhfeDyUhI/3FZVgXat21WZUInClawcz
TuzlWk0nI2cRQvHzuhu3sTDFKUBDV2hRYj+bsVNURoNn5x++9Hrrs6470LVs/UrM5hOrrogz8Iq3
Klo9SfcMlO/gunpg0p9H4oVowyWMWAGCfhlcrKeg827rGiVB3bq4ob3tDrWauwTgll+7riDM7aRH
qxgnxDxmGe8D8hGidVChlTJ93eWbOQvJAbWwyHM08PY5jFNlQVD44JgUOkPFN9CXloVJUDiL/6NY
5mZ0Wn4qrRYGtC8FBXg54AXIL3HPXf4PWkff5sXiq+L/kqhwCpolmcgtkV2qdBNfZVjyjBO4vjga
Yph0kKp1+vi+Pxw0kRmcHVNZExPZghD81MlpMaHPA0y5b7utTbWV4bFVz5cg4O7YCJm+pymljfWn
MU6kr+mMbJT8jg12PJicnl4eJYEnvDlOcg93eLWieIWvc8bUEyVLXv8apcwjjbyuAL/kBawYl5Wo
lj8uLjuKhPNSRGE4R2yYfCrnGAS8K2tLs+F2GWTaDKpPYYwjFXCsdfh53cy8jYt6OSNWv+sJp3i3
N+iP8WZ7b+cOt3qAcADjp7nMW1eY0Yc4oxiW2QQ3ybA5R4Fdm5GwWi1bs59EUCi92xE12Doir2+7
2i0AzqPQa8//laM7FGw0zfwsmh4JL9LZWdxEfN2Q8p5E38XMxELXrtZXHYLOmjLW8uNRAsVxktn7
ITEqppMj7bHgW0rQx/479eHaL6RKyTs0rLHqub5x6NixOTYRE31NJZzc8SzykDklr5NEB4Hq7NTR
NhJdNJFIPhB1/yyab+ED0zv34UoOLycpmhgXW5OkNOZBx0plVBWfbkeQ+s50ZFvsHvKoE80RYRku
foJ+FvqNy/BCFFFqsfL3//lcnZABvbVYsB+pQ5JsZ5PjcReg4UQPG9pFrgVggDDAAWqcRxzbzADE
juHpqp/XMfs5b1j7+Zrs+vs+NTEvpVnC9myyM1EbL3yHw8w70lj42wkCxhSinrJySmTxw5/0e5Hi
B4WwTQPCyVKqY5iU4KwFeZNBUh20Sy6bvQpqOEUyV6xCXN2d6thFkUybhq89g3ks3qP5HtjQaGPn
252QV1iPR5zxQ2Mdlxim5jW+1ajR0nJYCfMxawWNZLRc4XI8IJ11ZoAXl/URQQiCF1dbe4tSe4fx
eE8ICmtIR7skGOvCSHy8uAHblZgWJPNEA66PEwUA5OhoVclGdoSkwnB4dh947KPdUJZyeN5iigyV
TM+nWDSua4cUtvElexsWs3BEo8ocB/gioVjiI4fMQXMxhy3ZNkuZug1DKTZKm8IOdgSEGwigX/bP
5gB85e32bc8EdOKEJ134npbUoZi7vzQcMl0nhlgBSnFArOEd4BeI1PCHGnWsV8cXWi1SzdNq3Zq2
Am0gzzHt5FbQEfD7FT1cRpo+R8NsReH1NJwCZ0X9gRrqE/OftlNu2KIhYXGo3MGNXLxawANXkK21
V0QB/FcogRdBLEq0jeXYIP/EgvjYz/qqhGMAdGOlc1o0VIBR+RjPpDcq1OjI+DtyuEncyQNuGpI+
doMnYtXcxAHIgp+Uhl6rc7mNXLvBlcYH0xnkpCuNzAOHNpJw7JCb8jIAZNBrkS/kxed6TT9kLFxk
F/ZEqgUkqcvoeNLFyF6mQ0bB5rbZ1klR0uFd0HiUCAsBqePEOJVpvGIYSDl3lUdTGxxMdE9ejsLL
MmMEtn3dSJ5+2ZTCV3ZHxBbeN+v2yrcvZFisqA1mYcBb2GNXCSr8XwuYq8rExklDm8Wt+2sALUNe
nKMTwX1a6HwJPrynUP7RMPnvy8yQj/rz6nprEfxH8JIXCSC1B+9nnGpnkIfELXfiBcVHDA50WOpv
z6iLFIJE+fieSRcGowfQBMLMEze9JP/xXQiNH8592PcQo835kUgN6Z9VKXJUSQNF3aBRF4r+W8kM
uKHyPaN35Pa8WTUItivwcWwk++PPjY5yr4gITjzJPpcFLGYqiTBEnkf3l/u4lTJlPHGWdbg9mV/N
9bqN+3pZMGgl5TVl8mMQSKEiVRr+oGC1e9ekpyryKllgKls2v2mcE9r9GTP2QU1fI22TVYBa67Wq
qNEc7+xkcpu/u7zwevjZXW/uuf1kHaD7pVeEPGJGBoEG7ilsr0nI1Ol++E76KHMQujXN841odFWT
b+50jPxjw3luDbRmQ6E8d+X+OQLUJIH8IOI7q/qXAgiO1bgeKKfWTcUqwiubJ99un7tSzJ3nnPXc
yikvm4D3oFEicWnbQK8pkw7gmA17tWIQ0G7AE7gc3nGvgGjpVk9tCfODkaA5FxHGZM15YlpQGdPk
b8+cxjIUa3WL/6SXfNDZxd7qtHIB8DjrMQLYoEE6IBIplTI6u0iS95SPtKPZqdTbKLvQECRgNEKy
IbnmIjY3Wwb3SZk9JZijfjRX6iYtJ4rXeRWR275EdbGRbR0tqtodpNB0erA6ahA1BOt1GnjvcRbL
iyM6eoddQkZ5J8SLj+3M1IUGa+MTsmgebggWgmNsAJuFviSehfKZVY7QAw3FyPXcydEg/vQK7LVD
C93XgVTXDFXne3+6xWSeYu2jKsS/RdXK0x51UNDsphgrSEZdNwfGaiEEmxDDf3VR4aX7yQkAxbQ+
+WuGGCek3I1qyUy43Ei08x/xb+IVoqUHgqy/kQNBjU/kIFZ3oUPUTUSxiUqYgua3iABj31Z+Bbsg
qe0Q9LMkE9eps4nBHftXgQJ+a9lmM9rTWaXjdLijqQ/XPWEBXUr+WY1jqUaMr7QXNLBI0Nc/3ADZ
LwsnSie3Mldjdue1i73nMaHHkZLuGmzuzzXiQg3e6GqxPeXA8cDkl/AdHNloXwgS+ATNnZvQvYhv
xS7vnaajI2QLFQ2TE3aQagkg3suwUbjmtJykAr1v6Qtnw1e2kHzWuRn/Pqvs+Autud851+Q0SbsK
a/dyTLMsqo0KBr2XttzdV4WkUc6oWAbSK7s6bbqXDoKZ1oj9Q6yzx2sNQbYWrGTsofFBiQv6xWPp
3LsMo3TKepdqe8wCtspw7XXvCZ+zulgYn5YLvPgDjij1SKcmXbGQMY+AwFLh06r7EAQ8FEDmTSjR
r9REKjMhFEfwV1L73Sfgo6KJv+/icR9vCtMMisDvtM2Ya49DeWzioAZ0o0NjZU2dkuwQwQp2G+gJ
nABE1nkCB54dBTWu2VQYREc72BGsA7vE+Wm9r83HrVgdViauCN+vcfYWGVLD9gI5rxxYFNw24HZq
9WCahtJFgw3qWEgugD1/+EuMyCzjOcGKcDgD9JKCyAcAhjcMGzSuRQCOTEn6CILp9qMYkyrmGAjN
c3HGgqAtu4lxCn/BFyEIwpiLSRx+DYDMDk8+0NldIsf7es14bFrgwfF9rZ+gYqaAy4eWwxMt1AYc
2Ck99M1eTZHraSEnACvtK05hm88WmQZIvwH4VSyDpwT/eGArPDi+Szv1Vt9Bf9ArJo7gYOwwjkR3
9zSG9ebDnxyVHel6jzmCdkcgCYOvC7vBs/QUnmpTQC6W+EOL9Woxacmw7ZdUTGDunD7TwHKju19h
7lBJqjlSllB2PLsHlCbZMIQn3dpsahW/V67aONuUo8CYGYPCusitSWX+8SmcBmpQGgKpUHe1RePV
BI3rmdJjMfdLssmXZF9WpFYx/+SgdRkZJhxKaIBiVy9HUhJOVIrxRjAK5L1EeHXLqTywmgPhZJp8
0dmUCxrmLlI/g2T5/79/mwk6p0nEv7ty8VPrJacZuWRZvN2sKSt19gaWKQdA6t//OTcP3zJ7I5Xz
Xrxydig/9YyA+BVJOz7ClRzhLlls6QJHD8xe+JYz1lF4dJAgPpr9lzz4updQTbp3x7H6wVNuTJ2z
hNbpaK4VVVtsgIt9e8rT+vI7wY3j4gcK0MBTfPa5y2vx0vjkiXr2u9ZRjAlcFEyZ+RTNm/NzbYaA
RqbMGMxVuosp9XYG2YMS3Xdnz8HDYi/WONtoTC5wu9QZuMxEnZkWDRo0tezVklXpfT9pMvnbdK6z
9nc2R7iIRFY0naMLf/4QfQvMCLdc16e3KX6eJXfG2sfHajoO2opf/RGV9hwPGz96HC2lbDg7vNUv
0O04gJ0lM2ymPsNmPlgCybKXdsNoeTQNnQBY/kAN45rx/VNKsrjd1xF1oEJPv/lv0Cx7Tz0KI661
J1IO6x/HQsHnagp4y+8j9OYNNC1XfN2XcMw1e0TXp80P2W8OjMH7jaCyDpiaBxCxSgXYdjb/ioiR
g2a5oCJHt/S2Sja1f1cZ7KcAE/euGTQP6V1M73Mfy7ZLu+6pS+BMQ7HFH056fjV/XO8FnY3Uoa/Y
iqelkVjX50BlE8HMlsZck4ciqqdrTduaOfa3TRAyYDYlMiTqcFc5Zerzjo9OW1y59his7u4gyDB9
ogYrNRiFo/Tes+t4noAnm6kfFoX5L0KivdXOsjImN30TYB1kQhfLne2UlU2yNf4vQb+47mlCKpKR
Y5WxXWAjaFBhGnJ9FLjdkNR1sWqOr/zj2dGdO4j+LlVzVNB2X/qt1EjTj7iwl8ROE7hyLCaL7ORM
pJ+3RuKB6QB8y0AoirPHQ5fdy9p1sMUwgWtbGwGt6UcEj0SM4GAVV5XyO2erHRu5GbDcD7HhAOCI
8e0PxcPqpoheKsT1uVZOM5JFyUOasqWFyPjUqII7cAx/iFDuCPRSkLKaNZdMWNi7bdoGyC9hmAy8
K9Yls/BQYCPfDl5XJAr8YE31Kt1ZLiHn7SvBlH32CeV889Xbr37GwPT2VdOzBliDpeTzI+ZGUiP7
S+RJN+7xf6gO75Gb+Qy7489b5tXMhun1NEetRDv0VMjipZoY4N6i5eehtn+993+3UWuyDLSx0oZF
fvfHRsGE4/eNQoc8asLV6bQDFGLKJWrqWc+uF61DCiaiFa+b3gUKKS56GwFgEvL/2eW6/3evaGUO
vJ3gz/EPCMaEIfQbGeqhV07HVPSkO86V4E5PoEgLY9BlhYpwiD56VqFVGgSCsEOBnTbNjI1GcvP5
m7KCvJdOw5MmRY6STh3tROlao+/28wX3+ydmQITdDxVZlMWvuhytmZJ5b300JWf/lZs0/Oli5zSk
O2rUkrFAr+ZC9yPbtJwUa+y+3eXW4YxB5cnhwdc+tDY6Dxz4Yz6e2vX79j/rJ9l3XnHi+vewrenG
AHTn+O1eEVMy0sjkY5vDj8gIB8NACsmILFBV38m04QzsdDu6KlaCOy+cK4N+gdXE1gphtD8NmZsX
H3uPtQX2um8olNxpoqCdK1pJqq7ttnMeDgAIrDxu936jUSbdWfIzMTnO7B4kvkdL5pGXo5VwEM1v
cOBZSfnjym6mkNLYjwjTWw4uk1yWQsnTqiABpwPYJ7kffKoHVEO3qLezVO9EPuHJjhWpF+r4jD5i
xl4AFlA2XNC74jgQqpRno+S55K1PnR4bmRQWPd0P8Sjzvaem3UqJwLVL/hSBzfJxFsdtjLL7/yhF
HyBrJGdbzK1UEDaGtrbySWA+3HWy0moWaI6r9FxtkzGX3nivwlYw/SG/YHrViAFLJLSDxkNzpdFO
vMWa/w8W3Wdd8vbXyHvIi6msw+k22sdE0Dwa4OjvRtlWnd9yn/frhBS75G6pVmvVXc8VsQVw5hg3
Crh/NshEBgAtgZ9r1/LdsN8ojLBU5FRxBm2GBMvm3ksSU9pSv83E1nbxVvZUKH6p11tKQtCulGPN
ahNJu3r2or8N0f+O/xPL9MP/KYGgjZjy83fzIs/PiCDnopvFV1fbL89NZN3QvMWGrgoeHs+paWv9
jN42nZ/ZWiQE1QB7xsNvmGkHwhk0q1KWgvjgPvbmJ6coMHuexyR8HdqYT9Pldq0fYbDpCUfRbKj0
3Z0w3SYQqzTuDSe1ergCwjJL28G3L+fRpqN6brKqvvZBpYI5S2ReKBSKZIpKF+NArspuUP5DpG3p
0UOozjb4UuXG7SX63YyI9/gyeQrVeXBtw5B+jHWrCRkSmRgOjojwl03WHP6/1nXBW8Y+Twg1RlBm
ZdFZkGHlEty/y0KSlFeDzftPTeqJGuUjZMaHTcckPNodMZIzWZxV0ClPkA6OEUMSE3EVjCbG3MQz
PoLnA4KqhSUx5FYEX9e8H3ueFdcd7qQpP0R5viNgj3GysSijoQfM4PyKw0SsZL0lEsj9SZDs9Hna
F79eQ1sgX6nzRCb4BJZ+qjUtnCjZS9P2NnIw6Pg8p5E/wFQNYodvjcL77BSoEuFnFImki7U2O4Un
k5izQ2NMpGt13vxfLuc0DqW3HfcvPM4VCdp/59sPj/dvmOq6VdI3FYd+mqkcPLIxoOYn9ekZWgy1
x152jZX+HoPHNba6uIqcH/0fFrchON90jQwK5eJ41QqMBzl84vrwg+4FF0S6KmuaqFB9Yxl7/w/1
6zVkL0WSWQpAo9qk/P1eLafBT3ZZdWIxj8vESijzuklQrAWiTbLqwg/5GD9hMrZLuOtgcVHK8rDc
Vo5s1AWFweARjmlkEgXfJ/51ruOVdsKhfbcwrJvo8dh/sOmArqccqeM+M6IhBQ3WYxo8mT2XkwJq
+AMRKOBztMP4Gqp87kZ6KdcZFjff1h/pVtqKWxjygLdlk2TYNz4K76zoCVc1jeHIJ/xLtOa70ktl
alKC1bKw9DcaK8eelo7nfOOGZY7SI0vf8KJ/zROkeL6cTdA0AzdlTkIW7rHNgMfMrYD2P+aRKUIu
jaZEs6R9hOik2Rs1+XDn1ZROWuUyAC6Dkz2D3RuHyG4MVh9/pRiQoW4/MPuunDmFc/+2PYCICp8P
Zux2sou0z4wiOye6qb4V2Tsuhr9TWe0y0WWDJhd917TlHsKzNR+CkOupN2Pr0McyP5vDbo/MomMs
dyf5MWt8Hkog3gNamxsa9ufIt8Jjyu8nu3qYN91s6R/NPD5AInq8ef+EQcvvsiz4m19w3m2n19pS
kMx7E/s+N2ejHfyeEwfqEpnrKlXD309+a4GSpVzbr/inX5fDAP007XBhvVRixPGt6P2TQ9wNHG3q
fw7I/8iiYXIho1vmf+sePmB7U6vTdeB8ngh0PgWvq5hpCEM7KRCaiVmKOIBsND5p7rrPTc9HixXH
qWx7YPypkwfnQWlwGZk1NQuGjD7qRVgaRIi83kaqgvDHclLp0PT4KCOYx4XepUgVu4biv/BsbrGf
AWEuXmiaXXXs8VgI8v415/VBQ9mN5A2FnrTC2CmejMrBsxsiywhcZpI+hIugFqUKy2wW6GW+z+7g
A9dp4bRZKzPdGaypqwUjZU2jUk6Yxm9+ciO9RnpeLzUkITwnh4SBTdHSN163WL/ON4kkIBRa6Jh+
pn9spBX+ED25UyyBY97/RLn6F0EGOV+59hpl1HKaJRcDdOj55TWb+GZwHX4jFtxG/VjuilIEn8Ku
sw6D2fo3wRY+ji4nJABDxzkCJ5AO9C3+kTUDL88xHo95u945JJ0znNG+m4cXfr+c0G/0zVAbkRm1
U+UWV98H/N0i7Pl7NaZOguqs5SpQgg9OCbLqjPNg0ifTlF/JvKd5iDWvFBAFyt85IDaF3t8hKIOm
CwXCMtvg+OVV/wNDNxH9NSIN+58xb7s1aEm7WMuwZiwW66fE9N6a4ETekIeo3EA5t1IDk6xnX6+O
zDbXgnLnUUPXl+LNK8w0uCr6BTpCqHtntiUYti/KFlwYO/C3EjDgsFYHntEuEpPHaPZzueYYkqbe
3jmEa0bB4yRALT1iFvCZoFQhPR4RahiT8ch60dglvG9XCYhKcXcVkcYTuHfeOp30eeMCV0qI44HI
Cz/oUOn1kjC/O+9XjavkFIWziNKFHbUMnhWm+CExeKH6XuTKp7a1yxwYATIPxxeUsCjgKhldqnq+
zL7V7uF86j6PanqoSOLpMQBpLkMiZEdPhhQaGJWNrReQNrAGtEWQvEixAd1K9NP53mV1FbqPSJUt
IegARBKVHlMrB8UFHzeBSJ+ypuv2HeptjAYL6GNq5Aqmg8XZQfeWjrwGoRsTj6outQ6HCX64Gddg
0a+edmqU2tUYZCGOEf92mRNawUVcp3+5QXZMwGNB+L6pqWNbB3RzPTde5T/KnS1iz49FBUCfSqi5
yud7itZdf0ybQKN+2/Ka9h0O1KGYzlzf+zyjTPRS1fnp3me6D5yh+nq7CXnxScB5ufA0YqNSxcGm
To7xq9MHUfcP+ngyZEoscUEforvdhLG7ioSWkgneN1WnxOnkoFzAxdxqmWPdrdPzzYB8Rj5HQMGn
2n0xtk4YDSK4gKFhTWI9VBLB0WgqfP5IT+OAI1GTSYz2dP0lBU1M4Bk7VmC143vh8qGdUaNsC7Ks
OQhCLjYyy434WMBWZ9QBOkyiVuqKX/dqzfIzMSs8Li4xCirHTzTtmBBdctKu5PqGoff5u7GA5mO4
Ejzk34WksckP13prlFF7jWYsbIm3rwy1EPfwrZmJhgMixILun4BY9UMuM3IfEsGcD1fQ8iGhAHW2
IykgQo1rrtjlKuPN1sjLxVa147AcG7ezX8V++P9tJcjOde/2/s/z3P5xrMue8ezvj/yfm4IXUGf2
hIO3wYDsnSREEjOprzsbfH++767dfGpE0Re541bWN/Mua1oma6Ysid8FVXAwxYEVkbjnmPIgI/CQ
Wah6qJ/4DZ3mZTX5cEevac3j7f9kw/2eCU5rxwUq17wStb92RHVTELDbEOTLy65FoRsuh2CfxoYK
uyErku0ukucQv0HsouJZokOAkSsd9/sYyyLxwWPU8WjJCFHPoXAtqWbHueIQ7OBd6scqKlPq3QSs
vlt2jq5WqIFbEaPg/lpjCAHGvvePRoGZJra+WlLIzP5+PkzN67mAVjFWxku5Gnfz4gq2KM8l+Qcn
1Mq9BlsIlwMxm/IabEW8HlQeREpBFSiQRb5kKZP7H474kkyALw999jdVN1+6kVYAknB2JZTCdNoa
5co8VJ5JTYrvjs2NFBSrTglqQLtdxqXx3Y5cJjSRyRxJIG1bmfJ1MGFHStNxUnSTmEetqpVL2g/L
uLT2VG5ub2wJ5NQPEwfkf7qsb93qxtlkP+WKdZG5N7A60K6hxt7kSZWyARo9R6msBpKKOnIqRJH2
HtVS7E0sFQygTm0kkbvvOwFlNqIPCfda36ti8aDHuaiPue8ZLrqqNXCe+/lDH8xoyjLdKcSFb9Xv
fAnPjr04QQhIxra7EQy9QU3tRwST8Dpa8Uw6wZRA2cOJqKZ3hU9Ip34y/mfg+r/veNM3W38zlCrl
bATKLQBg2iSIcEoAqRBIkTl2b0oDZz3tmprrWyZYbBJElAb9ajMBRCCywWDBzoWzo+OlDM28GdLG
AsDboUhNeRjsnlKu/wJP2oumyGkclH45N/BDenWm25iCnYooOqEaxUuDGE06M3HkNpeku0WW37o+
sbk89xOEE243svubSAEljC1rYFYKeul7bWR+ESLLjilT9MCUO472Ka0xJ6Aqr1aPZoGe9drSf6po
CkkNOk8kk6Q3ruJLB6ZlDeRQ/F1gPpbA8gAPcao/BA0nXjoHCwQe+/Vc1FkD7RKs7l32CxZ7kcQU
IXpsz6CFdEa1Ow+W1TSCwrvatt3i0S7gUpLOsCHfWO5sHg0UR8guhAIXBYgKmWFnTlKu+2nPWCKQ
5JDCI9g7weaCWyq0N20yFWI4bIwakwx5JY7lOxdckvZpo3gQJJvfpnMt2NgTAgLzoA8Lma/h3Fmr
09ggOtIw/ifPb6tkqUn50NvBK3hA2bpGc+GSLv17xNVLAUeWPUAatvhf22BMvti0TCx4GDjv1BDt
j2MHfQ+xLyv2w3CILnpNwoUIrcqRTQHgHB8z6n8uKGngi8ZeH+BH/GqxkZdLB1hKMHBaJ5kiv2si
TsisZoBzyFkOSf1bob2LFGQInDivQTsD7lGRczNh0gK2Ja6RX0BqD7GTeMlQsoMDIXejwNH+vL9V
pd5vM0AMHtswsGU3KXh6iNsQjOl5q6NteaYA70BjLXVOR9RXxS7OEwjNp+Sg0p474z3lHEorD5Xb
0eymj97+/ArucQl8/Dfpc8km+RhEEJh3WsJsHw4pF15FU7eR82fZ//Mf35D6S4DZclztht8oh5Yg
nKvu9bjlFsfqP1ij0Zge1BESp/MfxupzQY6ATQfVHiw+JBOmwy+1h579sHuYdyh8eaVPkhODliMY
tsaYhvyM5nsA12D6DuEp6yprEXkajeUeSAwPlmp5iYt4lLmmxv1USxYihh7AnIw5brEulfbybGQ7
jr/V6fFXz1FEkYPRp9HqudpvqMKIeKeYWg12uRyjyKNh7cGSPYulG4cttPESBqALqV5Guwj2y/Kv
hR57kvAs9T72lJNuCBlEQqplZwmQhNmSnkD+yuSTOTnGG48GPVsTWn4rzJFB0KT2ornHAMRtp45g
zg+nEhcn276Yu+DmTjc4O9+MJQ9R8lNm77QOwAF/XJv+ymuBFVUNSEasfO/tUo2BqmlGp/Vj25A1
EBoLtuUXAEnoace1d7M+gjljnbA0xSR6Wi5tkrq8n2ttLVR4PxbWBXnK7u20SmiKbO5OPj79dKZG
tp3nkuN8dTn9dUaHOo+jbWuWZPu8AeHz1oUHa4BuWJ8MMsI7VoHgWCH5o2/+EbjToIAfal/WXr+c
ZWCWdM+i0xhjjV6mdRfFZSco+qykCcd2Tj4X0gEYBkp60cS63YR8RhS093NHBYD10GPyJiOvsNQ/
QecHMSwPJ0Vt5G7If8JQW4k68ip2Dc1lXScsp5aO8fQEJ8pMcpPeDWtu4j6xS4tWN/0EPWILJqUf
pknUoPivYiPGmL9N+zJ3yIBxDbysvVh9FjFnpKL77pxWGCm3LyolZNCx81cBeZLymlcd2HzE/c8A
L0IXdiAP2a7NOb5GWwbNvR0xXVY8e0xD9Ml7va3F1PF8cDm3is8hdayaD3ayh0Qj1KVTrJLVm6xB
wkCVoHeYED3CKj2YUJiQnMS6VmF8oxkT++MPJmr58SPVVnsQpyobLCwYhXuUOgbK1+i+ZM3Ak2Xy
K8dZlVW4nvffuNbhxt0itnD6uUIDgxOGAdJPla0h8Nbd/pLLSWTo6Dx5TbXZcWcgkSk4WcibuCWS
UVVWSlPmYcp7TYMjfLp1M4q6pPi/jCBmmJkX4G0ALrXplf1EfrfsCiGDqYEorZUwO3ghSEOv/cI4
b/SkK7FwBtfzzc1AXRxhCdVMQJKJgAVpZSSuGYdxDP7586Bu3lJ7AwvbMs1y/9n+o8U5vM1jAg2l
+iA9SYcnnCg6nwul1oAtPmEmhO88zCe+K4R+rtf3k5kLpZyvJb23ucwELgXUtikzIyYNo+4YE5FR
/CNNkdrusYcQeHmUN3/rOXRE9VxE/MT5qgdbsv26IJxizJ3i5CTTZ1CBLtNJTmljC7H7h38l/Nsu
AaBRUjJpVePQ8ocwEBbJJWpLUsIyiXIzvNzxDeky1J6Cgpj2gzuphvXNCWlCPIhsBADS4ADCy7UM
XOKlNV7bjalyeeO4uux0h2rrMP7ZwLPAj/6uDbBQ1VdH+TfMrywQwfwAhSGbYcSNplMt0efRgFsS
0V6FIScXYFXll/T736IK479GiBGvecz2mEUs2DNCsXCjRe6lNypL+n3T7DnhphezwFnIrdlmHdvx
5pGu4JxI8QU5PRR12mpbpf1RA4RgD1W54uy70gY+mm+LLeOash8ItxMl7kPkgCQDeNSYbHVCvjFu
p6Pkf2t+Begl/8tYAE5VC61CNtp7Wzp5Ub9oW4UH3R6T1pFi5OcblvbnBtz5s7eOVOB6PlmY2x+P
HS4H7Lg9lFqUnbkGUpQAHmjtfS4RpEezixALw8rBQLsXwAiQtsDOMjBgYbErMV6l/LnvdmBypX6C
LWOimfmltIOzaGEOHB1Wav1veNCui6dSRbMmgD0IZ9wBV83kVW0+glJunP51Jl/ZsPEbPXQaDxev
aI6XizetSqNOZDOvixeG7mAZ1bbhe9+3YUI4TRH8UtKCBOJGWfC0ei4gYzWaAWlIgPDHBbN7c2m3
kKzOqZwNMmyON2VFNCxAbZ8NkoIm2veprkio932I8GqFuLaTZz1uUabcCLNeSqDk6sM0dhPpEXpy
eg8gjoDsiKbeBs62CrPvFL87yVJp1ZoFcuWFerJKeuFs5b03+BaW4YkphybYVYb/zveV+ay7XCcE
KtZWzW2ODZcO5UjztNfLopGlieqbCa/lLCPdxsYSy2Xval6Sr6r89LcABrcgg4SrU0Z19+T0Nziu
scmhrZ6mv58LI4VhT0WWojmEaHwVslOvnajXVnmDihoUYth3D6u1dhOC4nT4FUIHbmXGhdDtnhKR
uxcTMozAZVplAEHuDAJ7R6jhlHYsmApQLyN0fRi6ArQWkvxXb1BpVCNdYDM/RZUhbtaIJJwgjh9W
cqDiQiypBguteUt36B9sfMJCr9mgBVT7pZ6y48CqgFxlD2L6G3fc3b8fmLkGbwn/tU2OLUbOTbE9
gL+yjMLorYMDMuPYGcZiM8vnjP6MgDJngMEkIgmOWeWvncaBq2+XKYt3oT9BwZbhmD4aB8DytZZu
6hGl2zKcoSBZBEZ3duPvz1N/ix+H7oPap/7aBWQeIeNw7Wt3BnXAYf12TiKw3eVKnZ+rc/sJT6Ou
iuTMoZMrPv12LrS8qz/3rGwgEzW04onI1vb6pNdrM3SEtyGLA37jsGW9cyYKQhDe8JsVqL6hrGA3
9n8yjOh0HBQH1T0qZMoRtSCjXAQQ02yE/JxhqmKkVlBF9NDVqcKIkE8HQ/MRxlFlME5Iq64j9lwC
GOkL0yJdiNxJJZHxZVymqgbVDWL3ue+oAbqlrTVLIeoGsYcA7vsvbza68n6S3v7771gXbZ12Qjis
yKIcdkBpHIxTGW3OoK/qHFPeGA4uDd2S8pMlyDzik9xMdhBzvacwTE8P+MaJ+ERo+3Y9VAgtljJj
+REII+/ZNiCauVq/TClnDxRwygJu0QaSG1Y/6GNakq/fyD487n8QOKy0hPwQYtW+uov0hBY+CLT8
HeDEu8h4umAlpt0mWQWPJLA/90Kn5BOQ6+fFhOpPxRWd+uQzO9uLjdoN6WrJRRI4Wj/N+r//2LUA
LUVHO5+1FkZfRB5N4mE/qlditsQ51xdcww5Ahj6EZ1CUpsvpei+1fo91ewkZuNAxOr2eXQV+BWSJ
DqkVSXZR2NWbtyis5p2Gso90KPKoMMish0Yv9xfiMflFJQrA8d+9i/PLUyTfLCoVZkCEN/hRdgQK
GaSD3qwNgvny3zYb5OooVRqLZCYuoMO7RuO2iS+ch12jaiIWz3Jzh+734vXG3tocOPg5WbprouQi
q/7kC/IQv7NBh3vNzXmKqAPXBe7GdoD7IcnJHCAR/Oxvmpb9sysFFxGmKsdcXBXmuD6Ra8HHqmFP
2b0tLU+PmYwt5R8A3VNiFUbQJIiVNQT+2nx8MxetS6AO0NGPZSUoLTRI8V2g1lhYId9OdRqpj8YR
0VotF9ozMctm2Vo3ZIga+r2ngCNbGuMMF13WwFPaRDnbpB7j5UtqsN6UzV0/0Kr+KVd8TIIggyZ8
LmjkkssVv2MqW8Ri9437eZMUYhDJkJOlLs6UE7qij5Dmza3IRUi5FdP+/dB2y2oN3wy17TLaQJEG
LJ9apzWGmObKiZwcj5RUNINi4OT/pC+mPhavQ6R4RmvNdc3bjZBvOnWhQ6hKX0CV1zNqCNQVhZkN
9QTswFU1zxY/O2DvMGu8eVvd+upxGaDwHqJoCDoreFH9+dyxgTp7N5eT0bd66gg01JHxRsTDcXRw
di+OsECMsCiVWjFOXQwIs/+GLRhnoO/WfXWqFY7Edgcr3p+gWXUbW/RH0DalVTdiCMJxofYjLyuZ
dH9NNUprs6cUx7978EYK5iylpQt1METPPLnQuVAzhE481OsqLErCqKZXTSulD/xJDkkiFMJlCiVx
vNym0liarnuAeXwQlizjGlywbfWcO/0eSxd1vXnhzT6hNtiNOztjsNh3m1Wu4wRyiie/w604apeH
1hEeyk2mn/FsBhfJr4NXmzKxhCDh2btCMFuYkMaBkWPtjiEUdokLLHGtEVBf+Uk3J7yvSkcjuDuv
ISapuyNI6XpYrKnK2+t8LAQf4yTa0J9o1rx7/FQQzh075Or7jNlMFgoRiZ6l+egSbMQn0Z+vha7x
9Xpc2NBTLvX7kv581QSIdJW/Sok3Ou98FVMyQtrBkModSP49f4aAiFvY/Q3OgB1XWor/1OBjXdU6
pCRFfq4nhiFhtpun9iDf/CwBVdD3iltEeoHK/xxoT8/fSPRiwmV3RgZcQQdEruHq9uMwX1UX4H3X
Mm4GifYo9DzoSAaekMcl6J69Yd7lK7x9CrBYCNNlX3u9aoKOA68Aau7eycrhOpbbb42iZRmP+pR8
ILqamUgPvZxyx3e2XooRQMLYSe8DZEMAI04VPFkmKyN2HmISGMjFCT6g28WNx+aIpcciXIZ7CS5N
kNbZzLYYF4urPA29xzuWo/92LVMvQeHdYEfjGq/1rcYM1qI3LutIkuJt5C/IBt0xu+zlgOOMjwUf
P75NacfqgvgTFki01QAEklTlwZP5kvSIaaoIbGKoaCQpnJqmJWFz5QjEkGSva4APohz3WzDhLDIn
LAX5B+xEvQ0R2i3xUmSN024Ru/sIZMOak0malkAb7q88SWdyFYvNmDOHK2OHLZ2C0wnN83+Ipzcv
70GT+WkvGyQvrWBIX1zoWL/rksOCeK7BJDfhS4pYWmGd7tVzT0DxvhOu4LTL2Z9lmglxtj5aaNBl
gUbJqyLYve10OYkuYs1jh57jaaBjqK0VRkeWUvnn69eOkJOLCJzoiTPMvfT3aEqU3aMs2Twq/N0O
5xaoeKKOJBIXswzfCnt/OiSmvvPheCRCY2iF9rM4Io95OxwDZKExidJiDhdwOiVdBTuPvCK16410
/K5hbZIkxt2DtNkIg/3iEpMfc+s/BoPHrExRsRtTTNaVgCggkwTw8ro1GO83RQxRUPzEizbHYYli
EsVdulWsSgTgfrfmb6XQkU4bQ/KeZQxZdFGA3GnqBl1RxQxFSPERC9zMMu/BTdgUhkYnCdgmmncM
i2OUtLkcsSkyvTzemsuV/BjaoRpWW310WfppCPoJc1NpCJNi/VNi5gGjY2XtJ5Il3TgBr4XbgRbg
3qSZ6HKkuVG6aSfwS7nTdoHMEQfW6hPsQ/WKmAu+2hN8lH3qNWFaNmSaz6KIZdZ2BYoUBCETVeKK
ihD1W9x10s3nMgmoUF6FWbkaEDk6YFL1vdF7uB99s5o2195O/dAzR2aZ6RQdU1oRr0ntmlAICQRt
ddBm12cLLFgRv57pWsCBNKgyYMAl1Tcto57JPZSrS4MyMncCssL4t4V/JPNdBX0izC8X8rjlI3TC
upwklmeY5NizDclfU1t+2ShvmRPUDOp5zhdOatNiLu970HVBOGXo3HEPfpWaaAkzVXKcV/MNbWKY
KV+yWIiWuTGmsiAbfujSPzkKQ0BhxFf7vbGX7/vNm4+PSkQ87BanT9NlSopz0hM7EqyRJXYDuetN
5gyjGKrw+W33LcSepL5wKJ0J2exQeeyEWjaI1eJJAE78mynTCf+d9tbK+O7qx1IbBPa6Hqd8phkd
s6kq/ILURx4/b6uSrhLkmO9Q0XjL98qvDmmSEuRvH0nKxEp5JPiEC4AyCbhltwYwYTWLetVD/2CW
oPmYZS2GU/dH7ao1fXCrVbL5tVup3TsumqwZPxuyUJTt/oCgwiFRRwH7Xk/Hc8TPVVGpkoazLoXN
wtxDVniWjyV5V3N+e5jS0vE+4MvzNPgUSa19Yc3v8KcIwt3dLhOzka7Jb457KM6BwKWCEn2Ws/hS
0D/AZxguHXAGELwYDW9GKYuwfi9fwxGnbsxQUuu84ZFRBRJ7yPIWEzKCdftuNBrZLBl7UXRYapgq
Dk2SZQGTU+xMM0nXlI9Mg+ouj0uKC2aBh+gFLoAZjV4lfOWcQ7KEyPIX5tu2koQupKgETLcUFm5e
Lh0t1/k3euP/knO7gKEm+vrk2xXnIcsAP+OQuOZ/6zeeuu9NDMAdeqDcOdwEWLpZtBp1uzqrF3gY
D/ln5DW45qepVhfescdqVHoFf2qRAR7qbG+m1dbSAtwrI3EOWb8FtbQXA02zQu5mZ8dPtS4yR4Or
QlAnMAYQWoiS/SV9hR4tXGONdsXS64zriCYCCttbz9eO/Yis5mW7R9IWByDDhQw9pQwY2bpqy3LI
PbhRMX/TSvlSGPont0+HjCH82s68Co60TB1XEbkv/NNT93wxI2U5JaXOZWgohekvsQff8Z0nUifC
LoG/ALn6KRlp0bvDFm+dXE59YXwBnjI0C+2Ed41woADvvhPrwX7KB2GY+NincXqiVvUvTWBUvSbY
0iGgCIxLQ1jZKSbTs6+vF4Al8KBj2ejo9AMN/RGvTm2lg+S/dKw+ezoAfEVykX6kWYWIzXdWV3Ra
9QJ1x6xvbxamg9Tu7PgvV/gvxHFuPYYmF1W8O40mJydC9Aq9N++dpuiV5eQesxE2zatERPnf1g4Z
FSD558NU8QtGVHKTnf0NGEDpXG5O3iRUDxolCOZSpLq/SOBM4Ot3VPQ4y7T1WVSn6GDDaao0X3CW
0IBulRZhFgbBHJNel/h2FjgWzo0A/8LM9KM9J9LC3oFqpGctLbh0Dibp3AqzjPgvLpv4YnHvzaFD
G+JdPVwksI/Gg2aU+EEtgQ+LwGwPsJGDP6m89GUyZnO7rkglWBseEVrz05vML2i/zQgy6L/HsqDJ
r6SQD/UAVvi4/2Jt9dBRLQsSCz2TJxyGMLWax5qEoIyNof7i6el5dO/TUTWT7Cxtzf5nTjU/9w/6
PU7+WEWV0dnqT5LPnQG2ib6Mf2WDszSJeS6nY/JWqYH+tYdXWy9WtbZ/K7hc1fb/AcHzppkgGNRG
qH8uThUp4pOytZ181IZsue0EXTuTcuiwoWtmbQUc4KuBkQvVVZGYagPHjBnCJ/zZiSXFj24I8jW1
Onm+6dBgB2UBIlb9Kc8upWlgwRQK9irMYRPsBVHqhWJEqebAvkS9I2YX/MRrsT/EJhi2ogZj2xrE
nhvWb4y/Styl9lkqORnoDuokZgZdD8zvHgk820YnlWDKB3aUoLACdidblbAOycFq9IbAYx55ePMy
dsX49H6DH+AaWwKoV8giGwJddtUCBDei/AW7X2A3Nnw/lAsDB/mJFiZiKKD4NITT2+euyJWmYK5M
/V9H2vj5bvtj44EuIclmZ9d795cU6/EWIZZ5k3Td2Gw7e9czNxi3WXnSNkj4ywDO+4grJhn5fVoN
tvNKmMwyTvMnI6YbC72vsACKmDdy7Sfy8O0Wa296g+tMQ2kMuUuWBWBKz1f3QidMmXzCgyHQYx06
VtkPEK4x9Bws3HRQs9fxyG6rr4MFbOuH5OwPpyf9ay0ZY9CWKN9JbdWCufDiH0Dt/4OBH24rHKJa
Ro1QequaZyaMzAxQoTFI/OVbEeCm7HfelQj4e7my4ZoFg9neRwZ6T/lfcItcQvRxkb2bNkJi5dj3
C7/90CVE7dPyTSOPWAJ7km0Hj+adMofQnZZqJIWt73bVNcWglP1f4PsdGuvjTuEw6SUH0Pd160ZN
vf99XF+7fp3z+DOPrhu7lI+kjB0yhDV2q7wPj0bsBOwTigvzx6Ny8x3igwKMhczbr9t8Y8gdowyt
NyTA7Ci95mhr26sqVE+SzFK3ly+XD8IuHn1WWwQ6Ph6RiOnxhEG5uNkxIUr4GEFJQXsromVzSE4L
H/6sIq/06nkgb5hvJcIVuONFiBOgtdXEK0+X0qI8DjI8HGH0qQ4IuCSdS9nzRPaKFZmDgC84bWEC
X7bY13KqRtItpQKtufjG4X5s7gdHCkFuFpCcKYusgIjdkBmCgK+fNr0hqyCDnqRXhVdGaJp3fduV
uZwwnaR6MB1oSnpwJsYK9lxPU304yV17dIVZ+J13m58XX9FOvNQFMm53IvDbeY2lXAiQucjaQHdP
922gJEhNZziMuUv44ITv1hWOzHhcJv7g/7I7VUjeNJ4eZpXy6lrSSslMkH3RUxtyaRxdBVyKFTJ4
Ad3QCHlMvGs/9aQAsRYVR0iBDcqYwyus69isEdBsm7qlqXTZjxhFwhysxFohnkR52Vm62oEyQdu1
vNmN1O6EJ0skzKTs1Z5EWVRyX9m+i9Y7aai0kpuGjg8VAG0yOdG8ELY8HdQgtDxh7IMQCfCQKPe7
FQfRB46JRUzPB3fykJBoU5N9YxSXbnOcabxkyxSTnAIbyL8Wqr3qVFavvytAEccX7qVHtIFLUX0S
8tbSyIWPtxTh7w+dxmk7KE9PjiID8mZAauQM18vqw83S+k8m98v7LTaiShCbIn/ruKdDttfKpZc7
A4JpAh+eDjTahJ0UcUZN5wxVNLWTR1PcVlEHG18iAK6O+DtyxZNz/34Hs4tmwkXWENPgRKDWjKHw
CzUgNoyOU9RfTiav0afX1qVV4LVJoDV3wmuIblR5Dd6gXuypZIlN90ob8fgXl27jiWAir/RweRon
oPW5/ljjC9O+kQhWxDV0+cE1DvPqELOF0DNWlcgyr0CUzCpQayty+1m3TG/nepU9Mt661TecCo5l
hLEBlCi3HWy5LRyV1JZLbNNRvx+OIk52TdDzQ+TXbdhfyAouA/k0/Cme4su/DHCdG6QzkMBk3xFs
XuyVVLp5nd8rjFUe2pDFntQt4dsReJAivgsdSXDD1fzb+P0IfrFrHZgeCGEoMPVeCd3W3Oq1ifBb
LNQd7tH5LEaTSNURGjXvqJLF9V13pWbKRjD/vbwWQXHpAbOaGgpqHt/UxFmeqXB90GCQ8G1eJbvv
81Ktm8YNHuZb0HeqQSATd3AqinDka8YnbzQLWwOwrVXfnk7P4Y5YNyCKFoN6QCVYepcedXK/4AB+
MhsZI9QudhjKbEOTcyfOwU75qDZ/zjJGFkKLhh7tWL4J5Jew3nhxdKUCXbh/KLIMPF8yqrRcxckk
iktbt0ibncx/+R8GKp/cYrT+CJ2qMw21T+kMUa7Se+xUbJJilowY5tDMRQlnNA4g1v4FTPeRPFc4
7/y6+jDrJ4pvR37TkfZRxtGcmBgKx2aWoNehrvGZUmBiLYPyufD4lFd4Y2NV9Gn9PxcfUIyr6d9l
qEHCcvtcLdszdS6y/RL8FIufuob6TqAXMDnuz/Nar+acxD7D7h9E0KOfBVtc/MYAmKMv6IwHrgPe
6duvV7bBRrFYxlvMX2sj+HyHPgnlmJd4RU813nAgDE/rUWx6APrru1Q5VulA5NHFCqMyOeVkg5Jg
syXpAnfuBEXUwknFV/yNcSwhGIvC2p77cIXOERiLAK3QW0whVx9apqpOTkdOWm5QpUchwsH6wEPI
HGnRG+jEOnK8r1Zkv5csZ7RsUJVhh9QumexdMfpEQlOPzJOnS0lBNcbywQfLDKZyOxlya0eQ5xce
meNcEGB15SOg/Rky7V+tfvAKYgRKGczkPCOrlmdVnkaD6jW6jqoO4lR7OOIMq9lmO94R+bhlg1um
2GMTG05iCMiJy2aM446Swh0OLCPI6nyMb6WSNGpdKIq4xd4UhlnN3369u55vNjAkKaNF3Z/DLknQ
qKdmbgx7b1p9jBhXExRWeIhHVoLOGY+rQYIg7yerAc6FvUjvoItovR2dYfkUzBUYYzYYUJwMHCpg
kq4dTLoOflM3Krpe/1rIc7+NL6nOD4lKztr3fdwu799K5847IopnIP28CW1iHng9DgsGRldKJUO9
OKU8jwRW8Qp/J9mAMTVi3/Hkf/7mFsodXMg+KR2OAxudClvyj/B31TZGqClFOx9lMbZIlOiNirZy
96v7LKQqXUopbntC1TQmEA8VbCt3a0ih8nq5jhzS+KZrnAOjBmG3aTcEzwsyPxnmRYx5Zh1l0Pu/
urjDT3lM0d51G4aTjqO1UuXMapTvcAAB0B5XgzXUyTZaTEJTfcChts5g1ZWBNU3tWa4q+mrJAXy8
xLwjQAsSh9ESQDvp/egvxZTE4f+TfHqbd8t8UuA6A0uQfQTa7xdUcDDq3u4hUQ1+wNLznnk6EtnN
RhirP9+CTtuG3xE0iwlU3/hBqanACo3M39Z85fzzNYPgM5rmaI0z67/Eno/JwMdjq9uAFSrayZnt
fJLksM6CmDTqA6HRWoeaCabIt2UMi+vu1UB+NohV5KGrkKg4PmideDTbMYqpn7sQ3fWgm53q1CEv
xE8VGAzEzt3YHMaryEfS9uB5mmlfWJlobHbh+cvQzUrY70j71nWPOZDRbZT5SqUSFjqAMfcmsoxl
m4fpmkftBq0kh4IZGciuHwZOjmE8NCVHP9XYFTMkWlthDf/RC+M1l+h/7M+/1f95zOwWFdIA7v47
hyNHaIk2zVjqkpNhWE+/Tm9ZomTViKsTSzuxKjBvI/2iPZrn3t6ZjU5BRkjiN5vR52+rQ1NwX5vu
dWA0enSuBNbHuW5mbwPHKPlDE2Myzgt3yIp66rcR/0lb4meTmrkjyX714hS5nXzhSnGTzTdYJZx/
kC0WLYOcVnxWYjIdVzIqcQI4xVsBoat+OI/ESs8zir6gklBUWg0sdNBIq3ip1iTG+iTMZz8fw+NI
RrAaYrV17VQhzLW+xbfplRpk1xYOacZsZL/v4Bp+gmeWrfl3sgbdphYQHVqchMDmuxB9Jfif7BiC
TxXRkf5pcWjezSxcpisUtXU6E+82rY/Yi9pp9PbRfgsTEjvjz8l04jF976YRG+rdP0NFXEUBltU9
Kw9da7nhgP8MEjGxCFbJs9cHbl5tIARHeA00xGVYsWVIJCTiuiTbYe0j7zNvF9t1G52ZmC21PSqW
+z8X8OV/X7Ikmz3x+PO4uWCkwlEHHWf3ZSJrf1mUdx1SbmDM6JHWQfnQrg1YCfA7EzCbWXz6AaAK
x4HCpSEkxx24TYwMqkFtavs61emfIgmrszPRTOsgXwkvFrhQW5oluCVbGp7gt0ShQeWdlJAOWKsC
5m6sYekYX9d0RdXcmAaeHBtA4T6ivNp+buvji2xPffwkcWZ6FmT59ne3jm2FaW7kNo0ohIfmNn0C
0D8lnF4MplSsvC3sGF+YBVKg0x401HaV25pfnegOtWAPH2tQePQnTuP+egHKj02nOtE4U8t81Wwo
9XVJDvjSVc0WtzyjOUwJSFSSvmtETfvuAQ3iybZqfzh6m9NFyxcEnA4WUVmsIS+LHAlUekU3h1C3
/Y3uMVDl4xOi2s/dpk7NEZafGJo5FuIR6yfVyeTTVkRIP6llTyIkyN/zt500I669Gf9skP1/xgua
hozBdpJ983Q/NRKCQfo/Ne4vutlW+2kb43zXPMVIwjLBMRQyzLp1czPrEeUi2B+0rUU8UujLpXZ3
YiMowOa9SvDJLFdwTaOPvzFqYy3yRNK39OGiJrajyVMqBFfxczjFPdyaNK5EFYZweG+t50aabAWm
SXcRzffUXN26b+Jkoi7Nj4xpmWLLR/7uEWofKKSScWGoiZyu0g9UhSmrgNNRohtQAWFrpHSZ2mFL
8+J3BozKyD7VR4NXyMY1zZaNH6BJW8p3kIN/HDNdYNXegPIaxXwmZ93yVNXk8Zrwteb9EmrmZDtt
4FGIKWrIRKR348ZL9brnGEqYp0lUR6ukZe0FAE2yC7F1uwYpGhhTiBEZ8cqwjzeawlgs54Ln+ZjE
g+7OHrufmwJ6Id8XCrMi1FDcxMo5pqyZUKFFY1UWyNcP9K8kLa0mmbjkPGV3kKOUnd44S5jMxJZO
fxA6OwmqSMSa+VQIWk2pydiUUlH/N9FZbyR8wQcFOFHcHJQRzhCnzLpmqfbh1hSEbbAkm+MVTMqf
uO/cKcnKCUM53KySTJjCDwWdzkv8lIJj7LaPmu8Xpr3KOXmcx3w3/fVpysFi2sJsD/SeNjwSkbqF
5hLSmeE2qqXQSGa+t0vR3OPL0yshvcbUPXx1F72MKayYWaYMblEGu22FJ5Bz3F5mkCxbCPF0NQMl
Vfmpejo2DYe97c3GMh5/8ubwvWae6Y3a6gRnMliWOZvVgm5G2rAkiG5ccYmBsU5VUENP9KG2rz05
zmKXn/hc5KNhbcIB0ZR6wkcRnxtSCRRu4sLJTFmIO8ejeSdNPHqdbJTPlMzqAiFb5QUGSjDwBn5K
tk9BBuv7VqJA627q4UdhfVMdL8GBm8x7aA8/Yivr59qaDPJeEkpHQIbVozuWFwV1sVsWfqVEMO4j
L0mpx9aoLZboOCDSN8thJKG/hBhlHvpdEitGgx8yq83C2ClZFkv8Am4242qbTJBZx5QO+EyANLOf
ZHYWQscC2jkWUcxR2gvfpZP0hO6aYC+GMe7N0eXstypJZB9BwtBViak9Xd3PasrwxDJNzaeGWVCl
ql520JG411U3o/rK/TKutw9kDuxX8Zsdxmg/Ahhv6L8XDCPiTwOzNQLbRQgd72qZojw6qfFGlnRZ
1CgtsmNdcjcI+tSMFrQwBgejiSBy1mYP6kWoQVVSUxq2oG9JNl/TggFifv67Bpyu9O1MJilpHdya
vpFI8BCAfkDLwvwQlyQo837n0pdEJ9ERVzoCEMrcYtHO7DVv1cr1RhOAfkvfmpBHO0Q9mk0svKKy
Sx3oJT8G+1OqoRoXHwr0QPwGOOKwx8Gnf90t/j5MQPtOJBBf3P13uCSYJ2C1FIuV8mvcoCF+f+od
mNzyH24p68vy4GGy+gYUJOpyjCm3IMidFmM7MnwBpK4f2y7S0R4n2jQiTXJDDZEYUlJro15S8v9u
UCOK5xz1Od5y4MOziwlmckvALTWOwyAekBFwZJDZdb52Z1O3FLsXaX3+C6/ZlF4ibMXmJLIIEMNF
WCeaDvOUEpX73jB91tW1UA2+IYdcTfgKwhK+h9PUJpQnNV+F+qFl0SjxhEISSr0cRxsSqDDJufSZ
S/ATi2PSFw8mwt5zcLGnf4yox8hFhZYk7a1+TwzXjHaej2nePhCAq8m1OT8UHoGVHGo450G1b/U8
bH7SU0Ptfv94d/ck4JM9cfCfVR8vqfq/Ke5RH0vn7fTGRzcXGTgkUHYcWS3jRkKS0y9EG1FsUYW3
XJkioo8ykoKtflTd/aSvgoKpJ1dyIwGh63I72BN8XK3DKEMNmg8VxAk+yqVtCIJwEL3Eg1gjyPUL
KVBB18BirtYlI0vKDLnSL5ylI2/eC03bxEjcQWbmcvXU5yj/EDQqK13QKCOiukdoUGCiLh/d3nmH
CgAYBhgZO9gXAFAWYr1FvP2xcaUrCpyTDuRiNPWs/RRPB1ymOjFRuT0CUioMUnO469TDcuCEZCzj
Jj841HPJ3u3QcHtyr7fWYDaW/SjprlYtCkzs5DXmqg4hv4DZvpe4ga21AmUSC5NOV8xYpPRUEIhl
2FYjwGWF/enLSecHstgTq3fuJsWcQDoTfIIzlLe9LPKt0w5SCAPcaP82g+fJz9aTLe6Ypit9TjqI
Ej4E5uzSgFPx4TJtK3tJ2NxgNdcfwW5+d8Fg3vhvIpFt36wW9rvsJucx3ns5IxHRcDEIOP2N9Pt9
DsQTUjEx+7K06m9gWqtMO51bSBoEUYVIGzS6ek+0/ZvfUhjtpz/X3gvnatKiE/E+UoTWleX20mye
Yq7djiQA3JMuQ5PE18q0lv8p+PZTP2518yV+h7+y8MJ29WPrhcLKQ8oj0kFYC5GA1xVq/oQQsvTK
cHaBw5nPgDddnR8S2jNw2tsZx6M6GyJHyIsBA7Ui48JYjzwTsfcvYvMsKGl1uiH7aDcY1jiWYXPq
exiVNsgE8UIUIQ8Dq4+AJaRRPWq5tb+/uy2iYtwlcbograDB4OIFU1xxM5Y7HuPJvGKaDv8zeb40
te8dkwrffQBst6nEnEAdHnBi3gJ+4pR2mP82iQsO+C5mnoT0Tjr0BYs80pruN+mnYkVG8PxMJON0
DXmo9q2POe5d4l1E0NBBunGgJ9kL17jsH4AkPv6IC2vH963ib02rMfRuix4Q+VdhR7oWpvAtP1ZP
42okWR/Kk761gSSl3iePLTqGzdjY461KgFJxHZgqOkhmsuGlbI2F5N/AwVCSAEre8+FjduTiBqmp
leQnW6GYZS6Bu9EErmnPA67V91y1niCUnHg1K03jYgyc1YJMPtDGe0AK7NEkKmPIdishB21BLkSR
08mj3o2Kxytt2tSeRmKYmh5BEfRi+gnbxeMOOGVJwyNhmGIvP+iwHcUW0CqvyCU1avI62gUwpnLv
gQdmH5c9ZwJh70Kc2g6hnGR0qhV463biR0LP0rDigkKhDCtQrWw5016Iq7G6/xkaterL5T/IopSJ
szR4JVftbOOCkPq8fRhApt+wtnvmyG4v8G1kM35OQsC4oQG0kkO1YCt3phyvOA6xJSgQZH+mSadw
/yaS+my4ZgSfvIykeH3pY5pGbM9ux8UgyjQr4VZG+cMGUyj76uKYGPr7Ng1zbCq7yekfA9Y7U4xt
9Kd72wNSceZqK+bso1HkfE6x+qDmMJSaJTlHJXVfFga98cWbZEY4VfXqLxnc00oP8GN+1Nadc/Yc
/wyaAbxaZuIi9M9YOTIzLgXMSJprw+u5obzHlI82dMwHaU3XBVy6H9M/8roma5NgKxwmoKijm9iU
vPb58wEkaR9DsWaRJlr95En1l9N/NH3HbRUrwNL7cT/bY/m5Mdy1DgOwssFnIGqERyzA/MxekXJC
izdaDtfRKxdGyRb+E8mbqpXpzr94dzyCdCKtVaiEd5X2/V87cPryeQKT7vZafv5fMpZc8/OClRGx
UNCJmN1P+pYTCSddBKKP4FN8WHSRpZGL7lOlOZa1jnYKm91x4Ax1m7Z4ufq428GQLxguXsOSRj8q
feRdeqXznhj6I11fhFxVE3KdOYrb7vk+cGzVKk6QPjVuiyn9K8QVJpivOEYweMZeYQpqqb7u1ulw
H1fWlVp0m+9CMVrbdSYXdeZ/PlBAd4L9RfsNO7cH9c0Z+CGyyzEBaZAncoRxvXzPHYbAkHV2TtNI
VOhw+0jRaeadqAov2ZmsNnNmexzvGZodnkmbGxbUTlpHp2gMXbksTSavlr8XVSNtmgoZwDaOKfmj
/r+14d/ICEIwngFzdYVXGbP1Lvn/4oxk7YJsg2IWefKSQm6MqE/vsqhHjiwJLMqQCNguuqzQrcZ4
rfjGJMjTxVcbXlYkS6TmusWHiMhGgit/BcLO8wqEBxfjyYqJqOSDRDHqCk6uYXSMdhYktMmKobvE
rpxSa1jb5NPGoOeuLSC/t0HMC5QjpXS5N9wBpPQ1Qf8gi638yWcSIuT0S7gDDGCYUPzW+DcrJ3Ns
55o6+oH5KZTtr/ZQ4KqhC28QjSeIqqp1TCa7DvfOP2C86SAEwU1h5tu881rd6/JbCZlnJ6DPOipn
Nelqz0SWVcGFpxfljqWV1C+ouEavoJ2ndDVYi+Pkw8cdeqwzKaFKDRU2EonLdx4Ti/kaMXIyh5sI
/Pyet932zZlz5KuH899bu7jmphieRU/Ly79YB4LXfqxWau9P9FqU3+PdziPrh0eHPVa04OZIGsWY
AtSnx9NCXVY7CUg9xR3FLO+EG+eFRQaXWsC2hCifAvRqXVni5CpvvPm/de5Aym4g9ahKtCuNdJFu
aVjiJKHe/Ln1xpAm4AcWvF/ejSnR28V4iqY7/gxGKvTC50vULdpK929c29g9PSaIPCeInDhVXObO
0hEKq+BEJj9YWZlhpOukY5/lQA9V+xibNdmq2Djkey51DBy6js01QijbizggDyC21Ot81mkXRXzz
EqpzOYkBuBVBH8iprhAbTg3lXVpSsGG4TlSZYDZqhSOraPPddJ4TVZZYJWW0XFWwk6p/wwgkrjow
9RnOK5GE5386lwpoEHiCKhE5fKsi7vfub1+bYC8zIHpcZVSRHVjhgUV3mJvJ1XAbM5Oy4beucvW/
Ve8OSLynFDONwZtwSQQY6+OUvGrTPiMf5ShHQzT/Epuf4/IVi4/iBMavGuTsLAULXIG1Yo/wTJuq
AjDG3bvYc3MTx/cUsr91ezNfDNk+38vUbTcuXBxGsOSoxL/X0c5Zn6956UeQpUnxXFvvr2InH+m4
frjoqHJh8AjAebI9C4YJvbxscVvLE9wdJveUrSZ5cYI6APIDrCEqTk4ehIwFQVtF3Cv75cM+J3yU
trbPXPs8FHK26wsOGjjT9KbeZBgUqNlQD5aNqR3dybwfyVlYF82d/BbfgD22aiM4n+CVxe5Rnw8F
U14DOCSijdEkb2EKLtLbWbNjfZprG5r0In9qi72L+xqyo+aa6NVy9Xt1ph+Z/O0ANU4Zhtnc8s2L
mMNmjnp4qrsMv6EK4CLQJPJlS4AhoEvmoolbx78osc+GnuEHaxmpcksHARxFM52a/L4r8tbiAgnC
ACmFqwO7eSh2+HQpwEju5ixyrIgTkNcrngEHZgg+XfWzYf9wTsFN2vrYPJ3avPPXp26c0y0dXx9J
yIjDkeEFfVZIJIuXlqqi5M1ytsM2cE8+mpFzS6HiA38Krhhr6QtbRqfMNvZ8P7vrmeyFD+r8imDw
BS3PQxxuB8mAQH1mbPF9z8Igl+L0v0TT2OsgWR3VeI8fFKwNrSn6kVOHObFQGZvSmle8k0SpPkeF
0cnw6c3LxwI0ZdoCFbPpGFEFbI7rummdVjrEsZu013XIv1pKwMSXItzU0WorwGKDIiBx4DJNYaHk
a89BcFiwA6ce1rLbgSVCrKi25AJ65XZw4c/ddA9EMIRidwD0ORDUnDu8uShz7hV8qmERyZ/1HspN
9uIhRnhD0y/Rfi5to5qI6Hik8XqPW6eKACEB4V3AIQsth/id23tPWhsja+ljhpjC29q2DGBuLoBQ
IzbdiGtXu9MR1iZCJvRu7YbqVXRLvpy1PuUIXf5HHoyTxq/NZhyt3Xkj+AGDoduFnW1d4MdB5yWk
vltTQpWIKO9tzPhNTgZCuIF0JzgjO0kAp+dkjv3//IQ2MCbkUD8U2tb3lkyIKnXkZnlc8Dt7vCBV
02/EXHzBug8nOOZHyoII6i44iMT4FldvzwDUW/MXm3Ngf4EOtreON8PnX8/opP7BP9okOGwzIyk1
TxMUJg/kJ+pG2ahoF9skuuBbCPynDeCbuTj/HQGV7YrinU9yxWbGEsE56c1wO3dIPBjBkgk8fKFF
dQ+okTi1qP+PeS/z1DrFeQogow8Nukx7Iz/OiaLjZNTh2VN8VAeWDVxZMGxh5P2KKu3/OoYXPXEN
kt7KvqAjKQ9DDMIKXURbf2boKzCL1d+vrbs4/eN6CdGj3too0uchbwfm55hlo6k5QnKWN+A8xXIV
ItzYCyIk+0Oe7IsbcsP3Yfd/rp7Db7JQTwYbaB5ixDUdby+0n/mmQ+/lRpqM9fFwt6hoEEmJmHQx
4AB6LsdIOsmUH6eioUpu+RuCujJ0QXA4p3dgK8bYlC/nTsH80s+/z0hRZYklWTvV4e6RUTplb4ye
c1lWQj7IhUIKXMNYh6M5E5fAISGnpEdxRb1mGmGgONByakea6wMOB25T6X7gq8W3iPl9ujsI/lsl
zbJS7YL/OxhrAP42Lsu4uPAq/zK8N/7/XZfUYuwvvsVlERCVyMiWGkjGGWUnNqJbQTu99OMjCzoJ
Ez2Tr/+9HgM7ayrMztGU2TCBsTz1MLkfqWTgVP9OaKadid8Qws/Mmev3zVrFJq/OY9hGlBlM/NUu
u7QdRyxdn68XXsMaFLPQwxlYzbC9RfNr/c6+Qgxc1/if/8ECNXKEhpgvsly6C+O4fQO1qAm3mys5
i8yh3vAYsG9QAiHUIJSe4CMhe9idprTsJrMa4jsW4R8pXNJ99Xarss8Lkt8M87XL164Qwmg9O/nB
h4Ne5kpHgP7uPOYWxrQEnBm81OCUPVte/L+tkOhbGzyvcT+7xF20hpd1dOKIEHJh4Wi+HI77NeIa
YAZlGT0NzKxq+68CrEk9+lKo1sYkTVFmC1Wg7HAkidqGt/o3xapB9DbvdQ7yJU5ZvPFQMoNXgm5E
rs8R37g3lAboW3wdyNYknJBhPKaYAC7G8LXMiQtzs/ThKfqVA1aS26EhGWIvJw+Tk+C4HbPS59k8
U5aE5nTFlcKeKckdxA98FzvJOPhecb554bfmwzUd9Q4OiErKkIIOhPLtqGbawmizfIHUm39eXJZw
pLLSVL1X5RHBJTUtRAe0F4vCJdAWUREx7/XLlfreoimcNyubWqVkMJoy3Cr03ummMSv+KzYCQazE
Ky3PGTlXJiPZf31gwwGpeCG3X4MsTZLK+4hcO5R5vW0GOZ0WJ3qbPTSpE1kjN9mUT6ahKoHz5pcS
SvYIuURjywmc72Qelyiux3/klysxiYnBjB6OIhXPMjasdAJXRXDOXsqzGifDdW1dIjrge5R62t1b
omZwTL/SpCWTsWbhoh8HuHp0xZUc3X65pJPHAjaImg8pipVdYKOt89F1V6sv0DZ+HKEKbnr49ezh
HOLAw7NPsggzn+UvgG2+jg8jh40NIWhq2LprRTTBD1e3pyMymOEhL9NO44eXuqN2ggNrS63qMXLG
vIdXuYNduo1QSwp6a0lHDeZYrx8sKkU8yGUb+9IoCHh+gaOCO/Z3GlvGU5o7MTGUJ1PRZSnIBdVc
qFf/38j5m+YVWi7ftYDnbJUiCWpTO0H4I/QT2OfwPzSq+KJjU9SgxW8wPC23f/MqEIJKYy4NlK5G
XVq+xyrQE8+g1A9NYy/ROz09cksNFeHEpLRgLOrhqPZCkr2S2NaBmlHsEsCN4K27vDi9rIvuA5aV
6KZKUnBOh5m+I0biAdZ4d/zPSR1H7VrEmnZKvmDp69WGH2TC+/cKNZ9lULPNjj0oij0bvNtAw8v7
T5HkA8O4fZRYq+stUf5JwbiXHjDsDvZPbBAWBtGdZ7TxW9duDTMNW3Ae1wFe+HLigJHAZdvmm6sI
fQOTKNOvyXFaQfU/z8FOIAXNqhCQkucl1UyJs4NIYUPsA8yvrBm9My1OWVslsSIqxtg6B1yvZwaf
sp805vWt0wMTiqUYnm/iiVdJc3ZnYqnyHsifWJ70cVRwTRe1kGVituC+Whbq5/WGklBIQQYG4v77
yYrcCzP9HnMu12/M8m1uNeTLSE5ceHMQf9vhWSdr/h7Ef62Si4AQi1Juc1t/GrO17xsOkyjypFG/
MWc0018JQY/OABuuD+TmBdF80mON2nrx9Pl3RtdoUImBHzX2GfAka6YXJeUIy9vEgxim4Zs7cO4d
PuEbQndTiERsJyQxBLtEDmPW46XGq0e31NOjHDZdWbXeI16CgSKyjXHJBSgpJ5YwDC0cYY9K7F2u
LqmiS+2aJgoU3g7winEZDgBId+jLAvxdCq4r2r3n42TaeFQy1Ys3PjycXKABbzMVdpgRzUf5ObjA
1OMBzCTW4Gx9B/K00NzumMBr1paLs+UumWhFw9PjWTdqkiGeEo7/q5brHR7FlRqKb9Kr5npsUqwf
5Qx/4vp0uERzg4vDZh+Qn1XFB1VuH58CMZQL6kqrRGxzV1/sdw7/pySYy8MSazocFFVVQlcC1SCp
z2mDq4XioD37Su/qn+UW16v3V5ICIsMgr1vh48HSKvVHPvkh0GWGvE2KXOCnRY1LBKuX7sct3G+q
+pQg+NqDVWEPY5aUNbFqtORyZEzZR1VFRgGv5A3fcDANPk7GC8pA4c3utZ+G3zzdW/kFtDtBmhn4
Q/8Vk99NVrxZyDwo6INDQYJ8yCKwGXieOMpCBnJ2b6yZbdqGoKLaZ/WrMDPr+Pg7ePiyKCVaqvRZ
4zdZp5KT35Ypa1OvDOmo/PnRiKA5MqEO6bfTkK2Gy+M5TQTf9Ql3qZolq+coDUyQbKPa84f6aED0
r20QUO88HSIrO6Eqy09L1a4kxH7EtH1HMV7PmHjVcDXM7CZZFpv6M6PbOKSSrieyO9zFRHntGTt+
L/de1ro3Afk0aceWHUNJwZ6wY4q/KNqCKrqfG0ITHJ57g7BaryjeKbXbxVMpUsMrOTuiDV1LhJ7N
c1/N/9Rex/QDeKmw9GfalKCNbJaMC49kVAoqTWh1TIZ34dfefSCO4DskInarNUM9msnMYpGD7Z9a
g55mPeClRCI9MLmENDLCp4vKztyZqxajJ+xOntMUKV7+eG9E0vL2Tfu1CS5cXXFBNxEPAORJH1ep
PyjcvQYronByTea/cHwcqmWst8ioKHiXoZbIV5pR2WM9rmvuYDtdj8Fqws+9ZS0ctwUlFYLWY9eW
jjLLS6Ruoue+oPtxkiAE2fcR1EdKiHen+zlUn4bQqOK4ycL3xAjSXjWksAnioDmPKsW7GvO0Vc4q
UObAp3g5mAWeaS0xtlj5+5iEtf1Vy+mYO14PBrM+BgGkRxbVCwc0Edt6vkmag2y5AXKe+R/+Rh9o
uThr8cVASwAG+36MhZPlf+199LljYTtnyAspiVoblWnVr0Tb1+oQ6T38DswTYvqS6nPOM0N9lRV8
ZrRRXD4pP0DYTkPdljNIwngHgc+3zv+WFKTe/7GBrx1mPiVC3+HXjmM8nZxUTgcb5wGQoM5+40X8
MB6dMcxWYnfpRv6DkOkxAIFvY5cXJ4Mtwq2vEvSHwVrYrYKUJrOUCglpfgxMuJJYD93kO8o2pDyG
1AtjGku68zIY9j3OwtMV1F5tTvjse/9Xafy75T4ucw1wd6KHfi/VJRC6hCVlTQe6o/DW6/rZks0p
yUPUvvoIrTDNjVAjePPT2U2M/GWZEE/Hd5yhQpjTM48V1+VuxAhuy9D8QkUdHNlR+jGmW4I8wMAL
IIZSx2f1n/UYDnShK9bxUHx8L7FrPXOQeYSl0FCAmjrlEq/Dsb832QpyzXU0s4z+qk1F6Vl04U+H
tjhR3i+JdPSVjNn60+sYYINCWQVNqDDj2/9JvEfh0AM7IKjxrfY7CATVr86TqsAZITq5qhAqQVPF
2I2gTwciruu8zkJ51N+rAg3jHb654zRXc7+mBQo9Y0skSzXyzPLJzh+roZMx2UbW7LhQwJ4jaevc
WK7kfzIE/5b6eh3s+WDYW4JJCPW1dT6Zf62oOYOLhbnmpCKQOsv+kvyA/4Woc1s5NGxSvSr9PVSj
SdHEA5WfENKOo4E2ByoNJqoJ9QadjsU8EOUFrh422QXdCJvEaSJoC5oWZ/SYmVy+McDrIDMlZorA
UFL3YjJeg5SZhuqK5+/KdkZIOApjJM/OlASKx/XfkdrgWU8OZ4v9U6Pf0vbwX4+TRQNLZ6RoXsf1
5aABmxQgA6Hb8ZVOLo8+MxvPIemCcr8Uk/3dKe9msYxxv56MFzszCKFGl+PAgqmVx1YUuWJbrvwR
ZcOp12ynK/BSdIJFIRtvLQk0qH97rXHgPTIPfHNWl7QAWFFX6pnv4fjKIcjP4Hx75/XRjR/zWsDj
Q44WcoyNPNoDi0/bRf9Va7wQuuzu/BWowfAnC7Mix08uZYHmkN6BJZZrau7MQ5nLt5mujxI8ikRY
LyScbae/bNd+nEqEo+bKkJQkWet6G2i9BP4ymU30kjeLdz85eozTYfm7DCuRLCMVPG0LIKIJCQS0
dgsIgH84X/89u1+ok8/wNBr3tSoVkIqzreK2FgvtYzqt0+UeTt+0phIaUrF52uS1h1vGu2p7v2mU
y6Y+2ve3wgcV5zjDm+6/1VYQAxdvTNm//I7K05cKOsc9eI7S4HREpOiY18rMPXQUnXzuIlaP19Z/
TBzopp6X4GWzB3blli5thc2k6jOWi7JabRvbspds/LhQZ4g5SlDKjrlDk0SXbCtYThbwVtmSJ01v
RNVVUotQEQtqMZEzDulOjq3mLBAlGBOfjIiRi7oNJUjgVbl5rC2tYCsY+5etWzLc2Jqhay/gwTDK
GAzk+AwEgBOpg0qtySPm00Eb2nAl30umr2R3Md2UM0dbccE2g8qbkFloQ4l2jfw7po/LBBdspQ+P
kSuzaa+l2XaRmeU/T1Lh1AX87T8xEe86HYq6NYWEp5BKQ2FnL5+gh1K/i0D8sbQsUMuQ+biasJM3
2420uEYMCTUJ1JCoVvdqdUKedqqU7kSAKX0UcZ1yDg9OcFFmQa+RadeIKv2hMgnHWvShSFQ/FInK
wkLtLfr2jpRpkBQZNlmxKIfYoEkhM38fPfZuoAEyF9XmqJd45bwKAfyg935Zzx+vnZPDI7A8XPp3
+tu5vlktK/NwOqaNg+PAZXqNlhqRrCTD6EnrHhWBInmIABvSCMCmDd91SDJfeuRrin0KlqlkkU5C
KTrLdmuSFldZpE2OEhHfJ/3zKBYD57bULzBptK1DCN+5Usu/Hfo++oOKP7dyN65sSFyp7hRd3XoH
1L6nejx8R+TSqXSsw0PDxcvjN3T975yz8ChIp9J75EjdXMmLJvkFkud/aGYAkrKOnn0nPsR+1rpH
kSfKS+xUuY6mbuWEKCzeol9MASJHZio1hRGb7YEfkmGImFYnF6jebEGv1OxWgc3JcZDOP9GLjqpo
F5Dvh3Fd0+/1u7QEGKw8x/w7TUg817IXd//WCuUJcb9bjGkRbxsNmA1CdCidMJspL+BAAJ4YQjpe
N9alzvAfTN4xBGa4+vxdZRAb7oX+4xLWxwECTaDNrIE6PndOE/0KCeT6qp2mdOpH4h6/CX6ySRS9
lC1dhMWwEmnB7BvFf6VQxlVE5p+ruFViM5qnd3Fb5ANnz8RgZpQVpJtdGViL2xPlwD+jYkade7rG
LIUJVqD2IqQ1ae00UzNyQnKW0MdnMZmGlMbiLmAWalxGDblkQwnR8IyFvsy57+H6w2oCvkQWpkBk
LsChsiF8eXRmcxnjfWE06ptLuy0C3n7trJl34N2GjhQZxMV9/Io9auBBE7QIUE7iy3UWMWBrir87
qCJTAUyF8cd8zgGLPRBvZzhcHHGwxBAXpDFCHVouVJHIW5MkN4ywqUPKKGMpjKot9MyKsGjnL/09
nnsySyVjU1kPq0z5xP63plEGHTBrW7Cf8wW44pCE//5Irx3kMjSbtg1ay/Y35VcjlQdN+yXXzRe0
oFkKbToInLTq1RGwVehXA6FrtzQ9qc1kdYLdaeAolxUN5itpfrVYQhGQjruCQGqyOlqEc4YnWSOM
biW7eowS3PB9ALbEgdy2trMzQuLUao19r6FSYKbLDGS/m9jGEyYCZf2refKXNY0cDrZdLcuuqNAw
7fyrA9mFWveyaxw+tGBFW/ceWOunIoNAZQcwQJFN5ZGAxqggfHgPguxkFU0ikXqErEsI88EqdBBM
aJS8ybsOF/+MVpmovO/DcyvNk8KyxmuCazFSKeZa63RbeCUOQMZQtHpUJYr4IPWLErka7tQ1GB0j
HDdyv7OlHRO5qQp/0ufA7ceAEM2Q5JwaSwTEbh9yQ0+bIVtXmDqpPK4ahK1G6WhsmytjLHIceLme
xZkyUjtpkOqo1LmmXUx/MgluhfIEAVIZpWD2Tr/YWVOcvX7i2jVJ4RCDrVdVMtML0qnlAJrqSofT
ZXomUHCRM/DQmb6K7D+iSjqmSUqyT/YgMwgRr2nhH8le35UqFqmUs/0Qi64Mj5g+S8eQJzaolBkl
8H9Ybwmtq8/c664O4XhDunG+9EN3ygTj0Xau6cbmAUvGj/P7+srUFNU3LjoDP3cr8sHcycvZiXxw
SWbnqXFprRo6KKBW0H0ESclUsWr5J+3qdmmQrPhQ7tvfjYxwzkHsolFnjY+SEaXe/qpSvMeIMAoe
8fGhMhNlp2oaBSPapQxU4pfVCPj8X43goAuS9C31BH7k7jhcwBT9a8w0npKuCh4u+u4nin0ISbMp
pi7VIXPi5ksD49QcWo1mVBFz7fmJk4m0NDhVjNBWdlpgk1DQzdsmz/zfjopVk6R96pZ3jJaCfGJY
lqHy4WdaSjjPUNppIrNBbHbtsW4ybO1zxMvigbPdzgT+7CtfhBr6KGdb+nB9tWdzPchSqbZ/8Rxi
T0YGuqUdbTSojT0+L2TJ9NBft8SNgtZ3luu7Ce+oAnx1WnXEdTDossRjYSLkQ1CowbWsdIw0bLXZ
pnL+XLuc+0jKxmyCVZxdCRxryxusVOkuIDkEvqE7b1RIBqIOSA8KYbeCd85Yey/A3oOp6BmpiKmL
vgjBhX1AOA5P2CsAZ8APDG0gaMPlIlAVblDcPkE1xC22BGWxJznR1WULlnAAsgHsp60SPmB4pFyk
dNKltUHhtB4/1EMyC2EBCTtkDnfMdRiZz8SJMFohxDjjQkNQ2nkiPIC6r9RNVHcpGgNYcYnmxWg4
VgoLZbv+W0ERxa73bds4fW7I2IohpBsQpKUGLBQA5a1EdEjrBQrOTyZ7jwun9tgk1P0dC8SQNZUa
ErPd8ZLDnGcJJ06yy7hIYl3Zu+qnGjVJwMjr/2JxwY4iMxoBDpfWKotR3N8aQpUwrwoMq8EPwm95
g31Sz0bUNFOUHvakgeYDsqWV/1kNx90qSayQf1g1e7HwGawnDKDPf9oJLz7jP916gfIAKdX3FLjx
CID4cqgQjeIOfecqvxfndLBRogwE2wuauIjhcyjZL654SffyYQt/9C0rxOpxtxYbEzlum8RfUnh6
VihiJeJ/og8iU0kPvN9E8b01U1Ug1hvqyRGUBKlN8lH1YpxqNYJVCpl7zhGg1MUll7ewBaT8gKDF
+BpcdL9L+ieYmBddIHeE4QNH5d/aRSop5n+76+Y9/dkJYNR/YHJp/IMBS4vgMsyESXWtSYlDEOp0
R5WcRg+2pXKEJxlAq6Tztbrh9VCQO1j7GekzBNkf0oR/HYofHIVrLGNfIuzinvezk7G5//1EK5Vq
SU41WZxWDjcveopwSPeF2FvcX4+jZgY4hEMGOert4MyBataGx+2JSZA5IqeeGLhEnBxyFr3dZZIn
IQ91S+rslLpq7b0a+Dwhg1JFAIX8rbNVernO7df7P+VVQ/+L9k3+umSx+3QcBV/ksQ++2xt6HVOg
q+tYwwdLqYaDP1tQ5bqkzj1EbrR5h25Ve8wIV45fgH8vwnyVxXu0cXVfSB/ml2mcHMOIEev7yS2i
mHTkR3xl/8THDHlvbrcRxZ/KvIp2BvqYFEG1EJu7IZiMjsrPfgNO54/NyNewZjtbFztViyOTDBpG
K3w6nE/pQmLd4unD2A0ghd3hr0+0TJ3Z5c+Kz8MdjYv1sZViEhZyvKfzOlfWLZzrUaamuOqooeFN
5DsUEBe3XxjoZI9WMCgOwah53d6Vw4LCFIdJK+0Sb93oM0/NKXW71SB2TEXGMA06oKewnRqFmeN7
dBooMstz/E+8KAN5n7m2h/kq6UQ6H4cY0JqAdEJQIAZsWBweC/R0vSqy46rwft1f/X9mw3poyvAK
MUJbmQgOnmJsMU3tsBjoUvaXr0Sj+1Qu+vdMpyUaMoEtgVNKZK+8M4iO9+BzYz9P+adBLgaRHkR6
0bee9Zr/MU1tJ5hQ8lkqC/mQgc7S8VByla7ixizT8Q/rwC5ErKXfteuzc9rn0SxSM0DpTFSQ+diV
P8kaFeqspwjZ2cP1RWUV05UTWM1YIbqC02bDxDNMhaI0xI4ceTTdDEOgbVITUqpd9djVideJkyeW
YzXx6FETAQGJ8RhfQ7Q/jXMzhmAZZHe7ReNohHzxxJlKrflLKD2sD8qy0GvWc3m/BYJ9G9TblrCS
NdmZ0Wv0M1Vye/gjG2BnQ7BoXmyj3HBYzpBjF2EseXk2Lq1kAWeTqKFSH9FUVFbO7AJsMtwDd587
c+g5WvqOdnriTtBhZsb7ip6rzeFOJC+Ro2fxDkVO78UlMk/68r92XqC6pcWGFzl9qA4mKu4dmj0X
32POzC4kPm/UPIouHHYjsuOL30YS2cF1CIt2l3St6XoLz2GT0g9hZGkGgOqQjEqj9XEj00e+0p7T
kk/LlbRf67BnxFgunZMScSfHvHdZxFUynS8GcVSevZ9eRThj8J15DziirWKi0Hehic/1o0T7D4dj
ZzPwRIrkZBMrNfIIiRMLkpYnTGc8CJ0vzuygU0wrRHZ03MLm50D0n/mCbpAGvvuTiHp0BegvZNOy
auI561j7BBWFg3fh8Qro2bhJPomw2R3dEXZK1WnMnv/tYo9QN+XftppQgjo+z7R1A2Jru71WBt+t
OZ/a9lBF+Qex+ou00FKR3iFWh9rfUv/5BZLNP3cKNm0a/H50Cn5CU5oARCoCMQ83Y93EZMWgt9FT
z+OPCKP3RH+ZoGFSL2OG/0YVvPkW02xLBO2lrB+/hRz0amlC8eMZBZWv3vXtHCR50NDw5Af6vAGD
6r6sbDu1ONgDlejo2b2euOJqaKXzmvKaEeUv3RMQe2g0tyqHM3wc8bN7MkV2DADzk0EPuyjoEGtL
6nC6C7ae4CorCCygZhQesEh9LhESgkZ+eSyQVvA4erFZbOlgmKrTV6Vsp4IhusDz7/0rbK+c3DmD
RMRWLd5yHSNoRtbRgvL5FdTd7ouYKKoX1GGgcP0FG0GBcAtsmPDt8S4Jg4eDgP1ysy5pLQXyRKHq
U8x8XiQZMN6VqeV0c7Mc1dzm+b7g8Z+wCTQPzBvg+42gMWeK9fQGnclepbHQnIWsXwHD7NMdhu0b
tQaBuOXhq66tpNvCdM5cbOjTfjDhVZMwWKjlA55vvjsjfyiY44sUbfJtgZZQaq6G2NyGFIVY7eQC
JCHz9u5W9SkLOC4bzqs12rRj6x5+nBijP6ZVwHb/Vl2UnrZ6EqPNdKncUlOEDKB45P2PILgjrj/U
eeBs9hWYiGsquwgLNBgNQPTeSW0UMEItTjriN5kUwDkHU/Ih8UToWfWWrow1xoK/XoHCFklzAorV
LqXyhN6SMCmbKhg3tuYhJKt7tzE0gUNfjrAOjAwe3UxhIZMKX+XGH++4/cgB0nhGCDpWuqfhRZey
gePgIQ0oxrIPBvjyuX4SpQKH338soNiNHVpqLJB7BfxLoqp4CymyYJqMQI7YGve/+lpIIV1W8PJh
aowub/vPf0dgY15lPpLUz6m88YGMO6cVOaOZLY8t2Q6NLe+pgU0GETr8BVdO3BlZtz3mOP1KZ+27
wIiW/Z7z+0oV7Okbgp2kzba+4HcK3jE8pTtihe4D8kQLqP9zVBMClN3zVDjc5ONWxpkpH5bVeuXL
sk/fpnQzpOi0rAYU7+o9EcJo0mxzDS760TylXr/VyPRKqhUfz1LYl/nzq+mI+yTKRmBHvvM5DI8v
m1cOBdhpKu7wpQ+SQduCYIKP4aSAi/GHJt6ozZNSZJuAZgNpDwPIF8RejiBts1QAdZPU8MKcwEx7
Q60rNPvTB8j4Wploj2c7KGnxEImhAIe4IWcnPC04L3zJPPvOdHjb/wRLofIaATOnWm/JL+E6JLQ/
uzgjNEM9RIO3k7b72Db3QwXe7E7NmoBeTi7AU+IYE8xzHqjZg/2jzqBzvw4Iem4MhUakRsKkF3YP
JT1g35PoXr3NO5n9SaLMf7FQflMnbzMcivJJclIWBtUhAvM5d85g1Qf3+N7LdfDa9ORUWxy/iowJ
2RAmT6j/FwQglr2+s0gkt+mcm4y/hLSzT/bbsYaeInCyAV7pHkL18eVvfXqEfNrnuEDaC37ycuVw
eoSKp8dOVBWEZPX1Uy/3ouOyPrA+32QffsR6j9SQokxZV5Y+KKveL6zGgJfmcCwWpqm/ipYzxa6x
lLe9srZdoEk1d4Xc5B3n0gvT7C5c8cyWLABmd3nw/xQj/jCwXcHjIC4howv4Qb80l88KUVFqb/Ky
1C+kYmujdJYfYrt6cq7BXuwG9+dsQq4OtkjY75c9PLBIhxLQ3AZaZBPvK4eu/JttpPHiI+FdZDDY
grwhyzH4vRmdmz5Rma9zbksdw+neWGLPUKMDvuNYTAE8VkP4rX223BXQgSTXvIbulyA58GFfCuWT
65X+fNE8UQd/WR4Nxx+lyvISPf502HO1+Zv4HEvnkT3eHGUptg4ZJELxON3aWF6ZQsCHQbowUE4K
P4WAitWts8T3mS+DUOazt9zrPvvIr2Z0k9g4GKC3PPzUWT9lugY35bLM6OzaSY9tcRmZtrL2773E
32taqiSMNWJ75DZLOVJwLMTgLJBCUeR/TPPmsU7jFoUbexbyFdOajEAgMZABirBPM+8ReyRKGmH2
s/zDFR6JwL+UsemgDa0gzRhn6t5yiGSPn+QOx/vnkTjXZwgSTzbmUlszdjGZSEuxOJ3qjCQJfWLl
69LiHohV9h2uIxbCMCHjOuQPoYBYvS7eG8jDG9lXcYs3lfK6GumRBofbU5Q1VAIfuuqmIdclZPuD
5bcyVIuJ0mceeVjwdmCrrNbfOwqxDWxEkOlccU+xQoMNxyBd4ZB5juB8NUgxI9AHEW6NlwQtULqb
e7eNqH6MFS3/RFC8qgM4NRgzq6g8w2WrzUvu/dMe0oAbC05RNubBVPePlbFC143P0GqcFHwFaXsx
y6LEnw6XDOhw9StYpDtIVCZaSWw2utR4Y5G+nTg5iw4XeXhK0rZ8IQmFO4Uq5nD+weKg6TXZckP5
JlLJh9vmtonTmIyxZwoNbXDHH4/sKZLhO0IBqLzUrvVhW+2cPL354dF0v2+vcz0UQF+ojE4GcjMs
Gym/mOxbw0GJrP3Dxd2+aq6JRvgWUkKN2vgIpxwHep7gwUdhjgyEEDJfPlh7j7Z6W+WZg1zJlzal
bv60ZNs0WPs5S/8J2iaC8OqQzqw7dFIWIycwGZq5+HnAHYSLnn/BsBrzA31QckOx/OrAdP9YN5Ve
W7v1dhL5XBlI6hdThgywXX4QsoAty9DKAGeWQrXU+ACxgrMclPqj8Qhq80t3f0XlkYPizy9Pgtd9
zN1hObPTXnCaJ2puNkHbv3Gtk46FQqDFiMRla/ldfQ2buoCqVDb9Nlg+zogLrSdETn7zWIlbhbuY
m8NPOkkI9EpgdHUr0LtvaOsr2lDvbWn+g54OYMUSdbGLqBc3I2mIhjA2FBhSuV5bzap94AaDOQ+M
Fbrjnt7N6dRId+RLoI557zUtSZaSsI7mQ1V0o/lxiJ9UcrBZJbizgHCDgVHKjQ/43Ai6oFeC0Bft
FPW7vR7qzuhkQbBYujp+xAtItgbfWMIadbSPSDqrt4p5Yyy8ORr7m0NQfUIB9Q7v2jdPV+0+0xtM
ld/X+rLzh/1Jhlfh5jjaJlv/58O9v7PTOzfxS73kbzjLJs/81aR25iD3234iTp99tvr0NoTAc2dS
1JmsjnmD837DmHVMSh+BqCOyghcw8O2+NAz9N8E7C8NffH2u6LhreAMSnJavPs87AiI9IJM1HIn3
NHa/XoqmFgKHS/SPHvZK1SF4fEMMwsXVEtxzODFAwaD/fsgLWHaS5TKrgjBx8EUGVdy2TWJswlL2
OMV7m7PILp3OiKlVsg+2Kp1F/IqMYvCeRSE7l41NZMxQColbpEIF8hGcOpRkk/G2n+2pWu2zo3K6
hPkRReJUSeUPIXglXQd2x0RPCykXZad3ZyWfZadtBrBY8o1zpurgwMNdSmxwMkD5+vg3jvbEciAB
gxXUNSboMVKpPI8KInX0Xy1Gvd/vmw8HL6irvjyl3+wSjdHBGmM9cxSGIvrB09KPsbBfzkF9vFiZ
kmhlaEVjXEuYS/ywd/kfNrKLfqfaKLWYAaMShqV7VctWOzT56bnQuBxjgCeDxfzq2znKkemceZfj
Xw6DtvC3bjU99QreIsX6XHlVY+/txNeZ5Z2lI1LSs7/fqKVAr2S0XePz8y3YQIzTASyLc+ZTRaXX
YxPD1i3m/Bv7NlINIJPIYtrTc3mj9kdijZSBm5s7k7ZdgZLOZzAKV07T0APLveBTOLxHhk9Oi0RM
p7Ll334Q6nAEBS/fwEwt3VRFVdPRunt9zDyh7mMs7X0eB9U1FQucBujWJn7coE6M3SCmyGIfF8zt
X6X5KzP9BHNCCfnv1ptinUODJniuWrIxyPqANtOVC0va2DZ77Q0AAEGd0jGabhc91+1IUaqSY07z
W068UgE90S4B1fQ9TnrFce5D2um5b7Kh8IpdZ+Qc4Bbm2IptFDLBSSoLK7n/v8D3p+afPUlZzOBT
thot+lob2/M2G1DNqzyLo10BK6YWgD3LCxMx8kucA6IIgXak7AqWwmXg2sr9hTW9/AJSZR8pjh07
M+cmuAJpfLqZo6SXcoDucRm/MnbF0Qrf8oJNp/S5yUmCMbrRN826caWw5xmyEQ2Ov+FKhjHHCt4s
OVepkELoej+3ERJP+Nb1Hn+0iA9phrL4ns5eMjr7NahSqfU7fPWKVRZaGdDPRMCHZKbppka074uP
6PbXuWS8wGOOKbvXYvewBGk59YN4B7x+NQqmr7yJrSptWeYlptJmYPnLxTJwkAHa7x2N18De2P57
eOMf822vDAX84dh2Mgd5nRz6KIIQreQjKHY0kh7Iv6LvbdvHwz0Gu7fuYj/vts1kxZkwZOXEwala
AxsxdfdwJxa/m7Qo7ZG9l0szO5O7Vtpx57kboMD5vaunfFlEtvuAveMQncL+rcyLojsKMMxJEFSn
lxB9BWUXj28suRxbPORmv/6CJcZVjBcYJKkarjmZ57mWs/k52HfqI+9HCq7oiM659UsWflwc7KVi
g3UukNrftgj4S2bt1G1xfqkijfr/EbCGOwvsBp8Wp2o2tRG/JgFXOimBxq8AEo+a06YThWoNaMBD
zUrMGtVk64S4D/J24rzuTlRF8fq2TjbJqKD7o8Ovbu4GbwzNhcZhNwoq2F4x2U+tjX5BEaA+gYTT
2AFud9yt/o7U7TJd3db2LCGOKiH6P3XlTev5oxZ/E9jANXws6UIETnm30WCKBbdLLVj6as455yXV
4+OMdo+HPHf5ZEqVPGig9bjv2gPNLM9x6+2UhsxFm4NbXdTIRyjT6aDY1mze6GCS/2DG+lZzh9MM
8uKjEiQhLveKJ8IIYDcZWKl+QXw8S95OY75HnXfmk84mOm1rYEklFrzW+Glwoot+fKYaHjSz00H4
ILjy2mLWSMG5qmqBEKErxIEr1d/4/Ot40pxH2gGsbwrxoDG3UTZdDMvaY6OCm+lyyEQeo8713FNH
7VEbxzO2ZeqGhspGdQTshYIdZ/RI+7Ky9YgXRkSj9x6b0V84QYz/EDnuwr+d454cU7aBtm5W1k3m
rymgB7Qz1ewf01fz7m++4U7Ye0WEjIzHRRSM+wKS9q67dbQattObVaAvO9ucHvrQ2HhCwD4fGXKg
Cgr7mSZ+WJSRVZAjyriNIpqprHRDH7zVenEK4vAxQFXLPh9rgt5xe3xfYAdf9D2r5NQfo1HwWwg/
0MPqE5izx+POw69e60Qu7PTxF4eDCcl99fZti+oqF+3CIO+JvtjqIg99gbpZUiy29Hn8RRXhwIiG
Y3FaNmraErWRLdT4tC3gfZ6M2UCZ6QRYbahVVcKB72Mpo8fEKXIMqGRP6lB4aVtwS2JembvqIYk5
4fq5RabXQmLzFo9vIfyTxpPW4obflha1I9GGl2d0Jmvatimw1DaUiQ9NzYWBRFfI9urAv/X5G03v
Bad31IhzYN3LRGjjPdYOJ4iXZwydVrS8+gD4rvoe+jSHjzLmw0bhNWcVhGYqRD8VKXzjpZrUoAFb
TSFKd+GyEl8wjzVbI4IKi6HzLcoij4lIKlEmIexjbz8uatmnsOikQLOZLEG8W8zNW6j55jS6U6Z7
ZhMkG6b1KDWXtNPCIrhVe57JlF0VryC9s71NmPlWy+IfWIukBGGBcmqo7H/m3EqpXOvSmLqsEipH
+RrOm3kuk3DCgkMKMfoL/3Ouf8c2+hf8oWcMLwlYtYJHHI1ZfAmvpqB9F+zLhUs4tbGvfLbj+fIB
ss39mpgRoIANF5OPghcSaKmhBdXyPC1m+59VSxvqFbjfZII+9lCNQiRgvPZtlljSNkxWpkC7bTeU
6SBUv5nlwKZxGagr7ii63B9x7OnLs7SzKVWACw4TeFa4Q1hVQacUjsd3xZdYJod9G5fPGEKq8/1I
vW4l18jCr4e2BXJrXc5SeeuY9Rx6fXS1oAIJkAvXGIwhiU0zrjGbEbAT+pj9+KAANwtd+H89woHL
365sDD3W1118aZodLM+AhAYoiLQViTkQMO6lbRf6rXQ7tFAwyqLzPISgU5ntF0FmjokmTsO5HhMt
aShSnWdy8wMFLToicyz0CY6GwgVXNIsrimVoZCBxJ6+A6iTa4+dbzvkQMNnPH1haCnteqd6VpSh2
RzOv9Qh3b+EV9KxHVdnhhbbqO3ctoVgbkHlPzNDJ4QrxAGAoempd+GK+LT08BZVdgqsdA/Hr0LY1
s5phRA4hSUIm5Bv/Kr5uU/tQ6K6NTI6ZRC1jAikzfavFZf3XT1xk5G5RmSCE/lfQfnykzycV03g1
Ki/o0zn/3a/tkndnnkS2mYukRKc6G73MkAT6bTE/sCqowMfXzOkzhtQhK4ZRMT3QnQQoKCvEf6aH
fAwsUwHof2XfQLG/pNm4xvtQZ2kpGYxi+410sI9LpOxWiqQWDllsx+mgRE4DGOezH+4IlTtkw4rL
n4ooCCiBgj9FVZ61rIwQl1SN4bHRzGL+RkSxnECB0if10RCt2lgwX/FB9EGTRK5HJX0TrMNhCzpI
Mjt5sw8Lh7VgRTiZbkdtcTaSXQReSmju6468BYxUs5Q4XZdWiGgdQjcIXy4e/bLzubk/d6iCDHmL
7BMxVx9yyW8t/uuqF9vIR+C/+GRkfvmqCM8rI3jGSbKyZURh5u5JTLnLSYI03sVXrafjFL4yWuVe
ORgxwpUvzwbOMv6EGPZEPvmGUffDyMsMk2FHbpYMJOA/dIEIakdWsQ2HLQgV8J0k1t6gTK9PbBW7
PVTssE7296uCQnzxjF8mKQK/HchReeDnS5FybuYRr+Rtt4d12BhdKooNgUShiIB0OrNgZcoLVqk6
A+tUJyd+MxMvvldArBxOl61rKTulo/EGxky/Je391JBSB8bUIW1T59q0GXDKXOBYkate2FuLm/Hw
zyIN7kRjzH2zTOWnXIjHf0+MwWOrD2c7HtsJnLE8KeYaaJld4CNMfOO3B5YMGPPFX8jdCFck6oHC
Qb9DEi883mtJHyUkhNEncjrPs2hObTSkK1G1ZwS87rKrqwvSTM9VgGPxfAZUwZPjVakpNhb7+XZs
NHYU52OVNW0rmH0a9jW5dWJH57x2XWk25b45mubPls9tG4qC9/6OycW1fY2j3L3cePWp4w6/qz0z
NWSQ3w4kRhi7SKUH/9vkwCqt8x2zI59ewdIR+Iag3BvcaQLMQbt6B6rs95MdRxu3CgAxfvItNuUJ
5u4pHksNY5wDvN01tWB0WHfdHpibm7NGvbUNl473veNB3M2JnNIK4wt69UfzamkW+MXwp/uvWBO6
KE/s9sx6q0K4iqJP26qOiG6YjyTA6vYk52E3up8Wnl8D3sW8Zl3lnBBnhZaNz+GtDbzYLZbHNWAY
AAfsAI3XKQqRrgv3u5wgwNDoN8wVoV02SfOX5qSSlbiAZNfiMbo16JTmk7w7bJw1TpAdOGNWJADY
7upIrtPYCY4BYZf1ofMVi6I0hiywtWaiqt0i+rM+T3pubhqmzGsMNYt0nEA0+c12a9oXtdb4igee
y2TVYacTmpGdXgQx1dheh8nkbATVCpGfA+8rxD9nYiWda331NWsmh8+hBgiTcPz82SLBwFeAErCP
X3keJQkbPbgDFo8fQf6w2YhPa8VUBQREYlds2HgtkkyiJOmU3tS5OLmVsO0pUw2iEFT06Exyv8YX
uJJ/HGApZjspCvJoZTnnttwmh1JmQypoNzxlJAvGOfNCC2ep2OAjtM9mMNreIQ18uPt6XScoW9V0
T1S38mP8PLKqvjVcJoGpaEpx9l+kjE/79gbTLG0c6DmXorEIeOEmvK22pCZMzvQEw82HWQTDcmVo
xDMRuXp+gH2TDDam1YB/lFb3Cmn2sxxMsufJL2Hkr+Ec9ZhhrfsYS2LjtsXLEr4c04c1BLBldFBk
mpYodlNIIKF0FLwihUKHd9H/83xHzA89UYaAdqvRctvDlm4HlxeE8v6gG5ANr/mBcublObyJiPu0
ee8AJzwNG1d9ucr5g4Woub1xjjkMqJON5KUOKvDFia1ZkG0yJwEPvWLUQH0sNy4ov5LchjvwOHZW
y2bdbP58tgB89N+Oadc3YATvaozJmPb/RAMyumzdKhg6YoLljYiVHmJf81OjJmQnEo+51hpTItet
bXWCirrwb6RgXxAYYAGUx6XIACZjt4+dQdbbsKpXFE3Vs2pcVfQav9ISFvCLG/J7yxQLNzOwD+sQ
+GiCeS82jocIvQpOglIHUfJ91j7hL6DIDzThfD/Ql0mcFS12+89AEXVdHz2Alge0a6Fbn96kBHAM
6DGMvtlAclP7tRI8pt/1HHqCk+0sKfZ752qqouNgguXTi91EN6JQ3gGX68njg6K8umF5K5Uv8x6M
/+LxonFzxvSOSlOIvYvzwOrphp3lhxjzEzGIDqyrW1Yig92ezpWAQ+G9Vm540py7s984u2zhpq4C
4Zq01YAhANeJ8Z32dcsecUE0d5sdD3YxjkO93Pc3lBba/V40SEy/Yw8nQePMrxlx6Dbza2u5eHsn
kvDL3UmYZQPBFjEKGZHEkyIo6voWcmfW32EutkVIjd0sF1p7ikilKCRZGatqMH+YThl2cln98ynh
8ZU1yab9uZWHjiR10j4q81Gl4Bsu91BrR/QnhQkDHh2cSXX+3fHrNIcm1iYq7ePjRZRhvan5sxYD
XfxztUMAMFx6r+OrjMn2y2e+hssAqb6D8oHBcrG5QzYZe1aFtxsjbNn6VPjuqWoZ517sfqY0dmsD
ueQTf/Shca2IMGZTVi7agdUEevG7TYwcb8yeBKRj969jnrRxR9ah71UrenbbLGQNAAqizm8HHCL/
D3XwDde9cs3kvf9eNrR6XCzHtE3HOBDmXyJLMYUTECzXVoIQBpWjeDihq3O71/R9/8BeOtEw4jmV
qARXzq69NhfuH52m5r2qQ7ZxBoOeFBIlE9SySrhYkHkPkA3L0UyDXTMPG0tyBUrIuErjW2bzhJIw
PdaBAYaUaguHaQ/ZcN2PNNS2CNRJXhLbgB2d8tpCv9L+d9DEkQZM99Kfjvu+b6kqihN2upk9wRz5
9zXiRD/gmuDtyNZqLiKYnckEadSWA2H5x7CjgP4XydC0VYFIN1lD2itk2Sts7yex2kUO91J6XaIP
CwEuk5GvGDFX9qsasQ8XvpLdW0yWwuguTeI9LkNC+xyKZ2B6acdnPzIv03TFK5Fsn/fiQU9wLJUN
nZ5CiZouU/QfvJtKlH81kvcLtamFnz2f9EZxTcHSdPf4kdBkr//gJFmXf4PSsEbL7zprvUAXqZbE
RJl5oaWw4utEBvSCNpUXjlTetQizhx0uThSIJsovfaTs505+z54BM7z1EInVGCB11rtjZk7ORcLP
7qSLYe8oOFs9fFvr9RFlgAEBnWCRWJSmqBSCnSPfDmZHrAwLGgaX5s7kkD5cavKynpu0OicR+0UH
pmttIkeTqbAOXGQXEmrMBrQVN/sNgSlljH5gFUwxa91a6npoCeqyRG4rRmEzcSscZyAqsgbozi2Z
xYGUrHLYL98ZBHTue+O0MfqaqnnK2ecUHlhtNgBRtcTn9y4N5mF2WwH0hgq48coBP0V3Ntm1cMip
w6fCRsK3x6TYN6gdgr5eZqcTAqX608ykunHfJjDpYA4O2ydUWph8w0Cp6e+QkYFZpRFuLUn4xN8G
H3TQmtcL05o3UFRxNsYZaJ06tN1PahIm9290RqLl7sqJvbw+wmt5jyYwSmf05sv2f6HiWyxygDbw
stPS6utAHufd1sHTNmZT6t+6w3J1MZw6IShYSveU2fdyH3wc5RjVt3kb7Tl3TvxfeTD+qFhDIrNL
Ba0fP+yg48QUSwv9O8FH0JgiQDiwbiDoWAWSUc8bJ5g0fZwTqhbuHU/Zpk0meAaUEnDdKSNHqWX7
NXlhhDi3pBaI/4fMW14iOoN+GmbsTzBIEJt+gLUQWmeQpY23PD9O2WfuwqrJbX8Mxp9MFmXY0eGV
Xola9PtEbfP6swJAYw0qeSKmvoDqcc6RAah/L9dNg6Y5zQ/MqeH3MAJun8cf2eRF4Tl3bMFbw1Tm
PEN8UXpN+jkw8JYnGB61s/KDSod0CV2E79nUHTEzsALfteP68eMD2vKIQ0bh/4/fwt12RWMV+SvW
YXeA6cDP9O8gm889AqLRI04BDXe10Vq2DRfXZoKO7owX5qXFHoTZPYwt2hzVu3ZQgr18i+4u17z/
1GojxnsBEp11zUJxYBEdNX/6IQq3PXTM9exYwT8RkCgjmbjb9oor2TzXfLRuolHnZJ0QQEEhmPl+
Kmix9W5F77Tae1UwRPLMaEBo/3go5Zot6q/4kKECFEquJNfztbjv+UQPGJ/ijQMOk9EVoKIIkaj3
6T6dMLAqvMpCFf0SaHmqrp7SyQfKe5FwkT2vDn6XcZ/Ctr6LZZpkA42je6Mugg4/Bs/kR1wfZXZJ
aWuGtuPr4xff2a/Qo0A1/0hO6qb24DtczxHfp51NcDUryLMTgOjgiax22C8ZU0xtN3fdFdXbB1NU
1P/gp73udkRxpVroFHjziEWW5MzrUd/lG5AJozDP+BXFEWyyYTjPLv6MmIEfvjU7vOFzJyYuddjO
QVOtVk0N9Du6B302E1MoEIbPP87R1TBk5w2YqsFu+35vadu71FKmPbS/yZ4dslAUqohI+Nj8wbVS
ID0Tg527RD/HhPoOWYi9ilM4I0My4eUNPwLaPn5wIavN12q6Y+Dn1gB73m5aVlsw7v5lK91tz0yO
GtFgieM4yCyjhbd7B3W/49YAnOTGiZGJLLcpq6yW+K5w+Lhh19EWHZvroUnYXFRvkP+3zHlLQxkx
VPj7nviGP+dW6oNYtTnle0Oy3tLKJu74TwX29sbFUROn/rGkYFW+2Vhxql2AiEOFn8Q6F7wrJZ50
vhDDTDnPfaM3++NfcPoFe0KXYIpNAO8EqmjU4mr2E7FMLj6sqC6KSVAO2lrg42Ch2E42gKjnQ19i
+ebDqiQpEVUTuVdfCB/co2hM8sjlZK2Tzx78eskt4gvny/EUMvsDCN168eEYx9ZPyTA5DEMDTaJq
jFVhA9FKYZ3PmB6n6AuNrmvmm0HtnD/4UG3E5qOql2ofM+QceHwfK8emH/SlgJWijIV8uUDgYnYq
SVxyjrrRzo4heDGriinvjHewYxirbRWWDmV+fdFDESsYSxH4WLkY/92xACmAjdkbHDfkUS8RfNPc
yf/qVY5Y7sygYw+yV5MOXj/Irbt62MBYE1M2fy+zR6JQBPzTKv7q1k2VKAkUUDzpmkCZwxD6F6FH
ylk8aHTNDL8hPcOvdrl0HI1VcLJrkey6Vc8tDD9YX32Sz0LhqZYLyNy/4VCtL0+vj4Yiw9LNpEgU
RaI+Lty4F+MI/dFufjTOkjScxwn9XII92H/4qobbirb72Q51qXx+TUO7fbqa1A5M/6M1t7b8FDIH
iL1vG+qI6lReEAiBV279NqBd38cTmWpjJxQEfOgviZhs/7he+Rdkfz32izqvlTshjobYsOsXpZM3
nCbKSHYCLwHfM+ywUBbTNw9jChEaeYcoSMZr2CAmqyj6K7LmYp0ows8l3UG8IbvdEu1FCJ8xAyzG
D+j86NVYHGeqsANmtpGomdHKUrv1MxapTiuYRPPCL+GhcO0aKUulx3hyr4DEvqRXvu84d7mOMnTH
IsmPgxOo6xhBfIrbrP5q5fQCBErMAPXknIkhjzUFHu3lkWq5QCJ7xQlF0BO8/siVEFC/qbrwW8Q5
2ERdciBh8XrOkeyczeUZDqvsJvFDJRtgURTf850p48uhi1rTN8qepE1FGEDWjblaPyoI//xeeqq9
6O4bKfxMaFBL9oIhR38qULceK43yHcBu8hkjgwvLYOkaWd6qbi5nacELLEi52UDeblt9EUJ5rkLP
XNYL30BUrxQVbvRz9Arjt0cxdEosLyd7je19/312vxmknhcZcdZPYKc9k5ZXWDcR6Bz5ioPKtNaU
5GBN75DFRltXSLicoC7yiME71+gxAiWy1qpvWu+CdKfl6YPIf8OLRYRv+X91vhI0iTFC4yy8XI+3
Jl6ERr39yQJ/f0Vqlq6EeT9oUXiKmhu146hFiE8uqSys7cTDyYyWIRVb3sydzTabuADsCOU8IhJw
NtVJ1IONs6+zU+0kpJ2V2mZUH5/TpOv883hHSC+s/wPpTonI6K0g4hFV5GX8eAoxSM/PNBtvi8Q+
zxZi+JTanliNdxEx/RSPZ2OYY4dXBnkAHwmXUAsdNryS8BqBabIaD61QXzSkOPbHy27gqLq55Opy
63sUB2Hzr/sxJASW4WmKx+O947MSmZmS7DRkVj6bxcry+yNHn2BH0qtFy0TKhG6GaC07oUhtgIqR
ii48EDeNAvg2Uq4ZHacKtPDIxSthL0tTLZAvMkQCCoNXdOVD0shm8kgHkDV2tAeSZ0VS6QC7zYF0
hxHBxvOSMkvH/D4d/2DS/I7CUbgD4Gw81qjNy9uKUz68XEMttDED9FbansaEAICoR7tzz1if7uUB
8BgPd3GdlkcJIHKRU6SSIdxQ2+2SKFQVdRt3Vqsh714bXzGiFcPEn8dUuAqScC6F2POjUeEBBg+d
t/N8LM1V+EwiruMJk99siBpAwcOtsUQNPpwjpOK2pL7FpnKjmgUnuUA3kx7BiGIQ5RYk15YvYf0f
Bc2XB7TJFNjyuArKByOsX5K8eSU3UsfEUgr7Bvd2jECGdu6NtKTGe8EnwjumG61GdCbxLtPs/rKI
0JR3XUKBS85XcA7IGihh0Gx+jaKMvQANg+69LTxUotgbxJMEGb5W96/W7ECNgluOQxrG1V8tm30C
L+qAOfyLzJVkW+KI7Dt0r0bbleemEpDWq3hcgYKoYOpA3LCOSW3Zz4VhrwWfoR3FIIgUrbE2c4L/
D4fzbUaoYJx+yPbKBfNPRZXRn1f/Ik4ASuN4f3hFGN/gc6rNENFOsGbygE8+wWa4PGCFita+zvZX
8gUVPxPDkSSo5XooRCnoQXeLhCPOuwHX9ghK5Qe1U3ERgueDhp/1BkaowrhEDnNlmeGeX9/TywjP
BvGCRqB60EL8GKsm+DZAAZYbkznzqdp+JryP7gdu4Ylp9J2w6Nxm5cUELaiXT8O+NyppMLrI83R4
Ra/CiR5q/Sqrz1puQswXA5y08wmwuYw/3C8CJHXArwJFjD+3Jo5+aUSq4nrMbhKTFxL4/pgmUBL3
jQwd1fGraDnXNNMPsc7yWdYAhFasNETmyYsNig6+7NAWLJH9bymIdGkZQlfqOItzFrqIDEEyg7ic
xgCg6yNPPGPAuseC4KvsaNaOyVpl+28TbyCbJnP7HAmcnfM+YteLU+avL0A7PXEUu5/be0WWnD6M
FLWQZ+gwNiEraRZQ9dHruR4kh/ATGeTqibyDlgB60S4+YDmgYwdRQb1RTRRo7bztmMHez0b0vyx6
9m57sDgbNLDPYNyyu3qXkazR9tewX+9D6CIxalVJMWrKCipolB3c38gftYrYufXg/qxCt2BVQuRQ
yaXCSliIp82YXy8PGz2o0oMUS3U6hsEf5wHoq4dkGGtMVDBlk4zlml8D9XRs4DIr4CXmbsdeyixr
jPrN01I4DA7ZU1tpjYLa2wxaeVKcSoNayCw8eMF004l0s619UGUryobEu5hz61xaqqHaJX1VnqkO
fSTi7T8N3pRsMa5Vz1Idsc43QarOMhdXVOtVKR6KPzTJX1EhU/wqY08HlepWow1zULVJmMfaSmu9
FgzTa7OC1/gUGuoIo97tmOBOEIw3YzxZyxqv2JjreWpI5F6ob1SI+6YzrS4TfxddVZ00VLf5B8qz
1KmdHtISOPx7BlQZRkERtLNP8wei/SAJF1wedLSxbtkUj+ScTA4FITsfwysqon66zaCFsfvb6Ab4
044jO6e+3ISzhJ+IauqhpmiUf4ZBgDQcV3QH99T3wfkxb+JnZD1UAp2CfeeNclyZL33LglnaeAyl
JA1I9UPo1zb7cPA+Ufa5HdVCK0Nw+ohVeWLK8S748egg2swWFXCjhUof9C4hDId4JP7mBJytEsO7
v8qqXtHeyf5HpCEoEqH4pETozz90kCJcvltizUtgev5Z0fv9enAy16muEPhm704VKcRscRU5X2p1
EdkQ6RjK041Fkj22CH+2duqh/RrVNubwPmFF0zTlMLBklj3q2ZufdbBfdVQKgMIJbX8PhAhjBicl
6F5oGXlZr+A8m3A5n0Z41eE9jiKyzJN3eE9FG1zFrAXKCPeZtjMBBzKAsW9MfTFTcW61TodemS4V
JAq9v7gMv11CH3fjbnUwpgc36y7qKOe0gQMdcaPBn5jTzw9S8RbdSSmCPp7SJggwF20xDok8LwAY
sHVttf9ctKV1YrjWfVoL0GDRHAfmXBH3zKMoq56GoCgW8KDEZQwe7vKuBo2rErSkO/GqVSFwteiY
+AVCUpKIvHnYs3kCiV6jLHBrNAcCSi9T8G1Un8sdFNOF6qubFH2ZcAlVZ0+zegWggmQreEEAfsxn
E0lHsJlBvRmbtODQR7kiz6xVArLhLfgLSzGkZ8Dt+iubj1TSTocwUOfZqklox505OLPr3mLF4H6l
9uMbyD9kwFhVIbdpro3WF/LnbT2owGQzESstFoufZRCwG0FuqTjVxMnl6MiwUFE5yzdAdh+drcxh
irBgd/rGNHaLFNaOGGcivXUDRYNRBqexDq44acciU3XI2+mo1An2DQwjQ/GXuRj+Odh7AOlFnkce
P+h42tlUyJK4cg8ORM1qwT7r6l7u5Hi/MhbJFqgR0tV5fLvX1xSDESeaC6sJK0I/rTc2wEk334H4
2dUdVeWCWyWcwNJScguV53uBIm3Q6Oxb2hmAAtmWYioW6I45ERgGu4fQXswG6ojQpeFrQjKS2X0d
rsE8x7vOTJXORunpU2f+3qJGy17yRSAy2WFCGRVa03HdihHHpXl8mvL0ekiqQgX0vgsAcYlqW0iJ
ppB91EvBHouI7C3h/pgjhznht8xtppuZE7ovOTvLOLyVB0oulMf/8wlunQfvT8OW6pdUJP9iBekm
Cc0RM8oxYzE42nhi2aG3t/SIKIt7NadaSSTl3pbWgNSldiZKJHJcqd+nruJegQlHT4QZqWq6dfAl
DRpvtBOTDs+1D+iI2A+K8CF16qDktP0wtsa1Rb9zrgwbOJ1epKC8Wjwkcc4SbOVwPZrwZO4SgJPo
vYHTkkA2I1GqC1KN+lkr8vsp3CLrtc1/qpiqOlVOOtoMY/ZM1qI103h/zyqH4sPETorskR84/wuX
ZvOI06CiKimhWXaoMEBTkDAAMe1b7hNhbdi8sknIAwadY6z2+uK/QXc3H/8pAfvv0aQlbIixn0PG
r3SjDWok/flVx7/sKsR1e2fW+jp8ooGE3WIFJQ455owKFORAeqC5J9WIczmXNNYWF0fhKhVM536c
ZJ84V2xAcBfcYvWEXOTqesUHXSLoiBDkDDsHqTVdO9N+pOCFNNpUw1ddM+LUgQA+n4Zoo2xzmLOi
j/rt7vqKylDXdcy3R8a2bRKwQc0gdAvxqnoOpUL9tiCTNQBOcxTmLGs0waouc0K6wY+Fg8jkvdjI
uSOV+hrLo1SySYud3cfpMLlQoI4AbhJu0Gl1huGcNSr83UoJHCccUHmqjolMfHtL5m1nqNPe0uB+
rGSWDCErtDo/5vFZtZKc34ev5iT61+dhGusnZ822CbDZsZFHyegr9EizfO0+0r+knJkmELJ12m8x
bFrtzF2pejVAuZ5HEra+alblTDh0UHuWu6brUXCUxRu7IiGzKbfQLdTT9td3D+jJRBomfnP8stXa
Gpo4E7udjwL5iQ8fHMPh3mRaSF/AF9FXzFv5KiExSUSvgj1iQz51xGWs/xzCHLtrrOIHFAyk1id0
Q40fZ0MBnQeDPRTYT95/NRZgC2yxmFtoNxpBdEYXy3yPpsFxmCQzpzqVuTJA1cLiep6w8cuJhBif
M+xDtQKqN4p60eA79g3r5hSnv1kZYCYlm/yRWybgDe5orBYKW9lJBrJPvkWExV3mC5O80p9K5/c+
kySIZ0WMol3Yvc3CFKzfWf3EljN9tky7XiqXgbPRzPUVLringGMcEr7IHIOt6XLZNXd9SXlWS8Ba
3YBXCh0EFiTSEDEW8yeRL9Gt4dObBVsYnsKN+Wmopa3t46hBWfKXibrr4kcXlhocOxCsaiae7PIf
sXPPQHQnY9om6Cn8f7fmnqeniUfhJgDwFAer6JMOCX5zFJumm1sIoY+dRY4xXoLEpp9riDV19+sp
9Q8hZ18eAswKhMhw9kU4sx/7ioKrKgf+LAiXLyQru0Vqo7M8EcM4Jpc5dP1dfLvzioJ3uFbi6VlJ
6L0cfd47mhVaLQzdS9UHBqMGMLHczjlYEuhrFrQRb1NbPBy6tl5JX2rNwYN8hH9ybvwtK361Fqrr
gJdGu9jNuR98zHYBHa0Ne3JCnCn5BYEsuGPJrt/X19bwYPh4WRTW6ZsrL/Rc0yyER/9ETGpPV1yA
tyrx54E3LO5AKncvbxk8/eX65OLuUvSnh5didqQFrTVgwy3GPK7jE+526XfxlVPI0u83/uRMteVx
GcPM9m+id62Yz0283yklV99Mj3QxK1p+k8IG12ywbOelYCxotPjFC5gFl2YjVTqfgLU4f0e4eSEZ
6MkFQehgjDm10SmDwUPfoQPrNb/sDExYUua31pi9UiEA0R05zRO8eNCpzuwQHnWEF2SagOr6D0q0
CqgGlQDxmmiZIdyJyTr0EobjCBRPXoMbMc0rVVKc7Kvd+vALjrLoNnilmEucYWGSjONjmyfzyUbr
Xsq09es7DleR26gS50s2Y7t6tVP/YEgF1e2NSBNhZpJyyS4UVBni/eslEPz7EZAmZWeSYiA/qMSG
ASn+GqrGo6Py9IyPgdMPyf6ER2HZw134/K8jkML2yufir3WB56bQ+2mThpUnSnxeyslZ0hYhYTPQ
J44nNC3jz+7W6K9LJYBH4o41tRi0Kn4JUi+czn8HtLc5Q8023M5pubV8qmD2VQCu0YW96gio5+Fg
7goOzZ5w/xef8US/XdbTiTsuCo6bx0lx7dkOex8mFLlSBXBC59QDjTUM5TANRY+kCrWnVJ2faA4i
e8wMSFsvJax0QY3mDq8LKVSL4ACp1NyaA8pho/WUZ/HOLhUSVmqqn+cFGJZWctB92JLTEpi5ibub
K0SVf5AMWd8aS6G0j3Sv1tH2gXjKeV6qefuFKdrJ8GWXTJnEK1hEHOjoQLrhP2BZIhKT4mf1n/km
GSN8y7AR0PkgYB+e+7xXpyDlITzTrQmF+UTWkhMzkOgat3kKF4Sn2YApzy+BhA9QI1yQqoYovuZ2
S1ZJJoorA6kHolMH2BgDPJ/gk4DZMSV8PIuAXvdTvLng1nkl8mT72i71diNMAvwRvP+n9emMnVNf
m6W0CNheOd2mfwxfke8wSczDvSpUBF6TwDHapD6Lt91EpovgpHoROmO51YFotkQUmJov6y2J48Da
yFSUDpXmrTsolGX24ZvF6K6ZMXkPz5EmIQgtVYFUj2zOTuQ3yJ3VryIqIqpEk54Cxy+5+iBDA4Cp
VE6H1Un3HIH5y0QRXeXJij5mOX5shdgREcmL4zndPXssNGxnTHmzSyPoI3x8E/egkXIE2V8KMiwW
AbIz9Sj3KiFgXZ+vCGEL8p/cb1oYnSzpfT440aRaSECSykkrHJMNXGSjb2WfRsqradxIm9RoH1qU
8eZV6fKnPWyf9ACPfk1vOmKC4jqPLPgD/fnF1ulS774/tMHrRldRaeA4VzLathVRzqYxMhkejE0j
e5gcMP0qmohJVLjt483oKehIUYGr+HM2al2gzXjhl6r8SUJDjJSycbOMUva8qpKuZc9/r78AI7In
o07AsMxA3jBqhOcO5kHnPKLyEab+cQLC2Dz9uCvYO3byvIJQQPfli4+ckQ4hy9Yli0/zn4T9DOg4
6rbkaYB5+BnI4y0ooeT2JSXaWdJW1nTJDIG+XXHOMye0W+R17yUkih1GWIvWWVodZu3PtfghmYsf
3SRSrk6q6Z75FZxjTVKqW4U5k985TP/g91YMecp06Fka8Uf2K8ls/xSg+n1fXjgfD/Evq2PQRh2J
oVs19qvhKp8mS3QPrF8zwTE5V4f9/IeEvhrYNI1rpWNC1m/PaMxD8d6ZhqbYO1vU+6epvcFnNrhx
bwhZNkQPKwH6LiklNapxmpaztIqHdLBrfcArzgkKyoGeiAHOJdpe5dWNl3llrt6xM34BNglTYc4e
egW5j7/e7TFPbH9jTuGzK85L26LfILIAg84NUegJHNNAWycqyeRMOQKyZ25Tv3uCPlZlcJ5SVaZU
XLQYwxZW5vnZSGjpE3fan6Q7gOZ5g3Pv6G0wp5lay0rkdPq3tj7nmDxEYX6QcDeyaGdPwr4iHJRt
or/cD4QE/RM9QwZZOcyndSPkH5vz7Z6yY/BoWWIUFcsro5M46vvZ8zvuI/IVKnt719DFqhIz0LsK
OgiOCbf4kOkudsYolrcVX7tGljL47dpiS9OC4BAO401APOCSphIkQFJQ4H4ET4pqltr+KOTt57c3
rNy+ONMXEhQ/FYphwixHYu+1uJGyouGAjuVmjA16PVtyGvosdq9BXf4YgHfiMplwA0G+1TldgG4s
omrmSSOLemDxS9Or4QVhe+oDdTwoRAxvD4U5qou+ceWCz7rrznOVolWDaGBPwqOmpVCPqrsxLZu4
dQgxDGMZptp3VU0tX4qNEqIhPlSj0TcwVMqHccQJeNdAce/jXSc3VZ8P2Xi0cLY6wQvOdd2xhqJN
NIGUBPvbl0BVZWLdZpafGT/kgNSg1EVvDXIx+vbnAQ8DGuR2hUno8GjVqy/sLHhNsxZPf1ZJDnyv
p5o5xtMPehrbVD5/fUlv660AptUS8pB55BKu80+d04oFDtQmBl0FPgrhoqKvV4l8tyS4zxZAHlG5
Qcjy+YYRKr0ffVwMDNTKtowcXlvj7b5uyO2zAkDmVGLWRSFfUezyOcbJ7OBFyAFkEPoBSQNwhuCQ
vIgvabHc1YsU/XrLAWiAhf8fv0yqsEkLkNxAYq3YNuBLGu/AXmNf4a/k5+/RGpCgZYgxcjpz35/q
Dj2CPz9IiJbAD3xoh3lHEBTCHowjbYBkmylk5nAAMVIOSwgZSNsz10ldCzvQ4Bbwvt+mbOUt+Ry/
Ias8t7lno4lhkD0h/lbHEJNxP1lmTFPMJ7x+eA2gG9PKR8aUpBYyMZS1OtuOfjVxUBeuH34iiR7j
vIeIwEwDgUE0CLjathnYKTffeoLnTh3ifs+GTkBmbJkXrZTNgNcSLenFvyBbb+I6PaAEqPOewdxC
o+gXTmjUqFx9s+IHrb024EzVCrtNO0HFGGPzl0a1W+kpAzR+ZBEdtfq6BcvKJRKW5TORdOhMq+Tu
dJTwprHGqkG/vqj8vt7TiDSDi51GoorwtBh68XyySKRbBA0eglYofkuh8jwmVY8iZ921W5HoOfkz
shRVP5GdNEvU/47l0L/COJZmoH2T2R285rrNdjmJyIq2HOWR4ZmX+I2zzdvhTG6aJO6dxvLf6MTn
KlcZAkAwzTjwU5MJVUPSWSY5Gz4lK3CJqGpRgTvVWtlpWfLohrxhEwR1ckLkKUNE6q1YUdXzzJ8D
YzBNxI9qsResWvgMZnvxd10jFzpp8S/wwqTcZ5i2zD5sGcqdNdSV/+7gUIWk3MlgBxQy7qDzgqYO
ugra859t8VgHbMaQ/W9aCwZ9LOhUeDaFc8r8j/S/Fq3KxnwCPIOqS/jN3EO8snxpo2cK3pEL8Hrm
znLRMG83WMTR7qr5s6VgbSybUxvOuL6d5CntG/MaUo81DMKoptoBHp6C3BR+2wVD0wix3AGF+qOQ
cJOidqO22UqTkpl1PJrIdFwUQQVlnqDnLBuoP00shYPxtuV1sIqYNOanq7Wm9c4BZ2X8e/GRIjsq
hDEAFvT29UetIOCZ2lpKEafvtHffD6RuZMyxgqwOvqNIr77t1W5eqFIfDc8Vr5O5Q2n3UiARVOJr
YbCy9doFgsdMo01lfqODfYGjoC7KRtJbv8HfeNSUKVGCE3iSF2hkrSduZvEsTXxIzGsaZF5oLd1c
ympWurqxdv9x7ULLmEN4Lf/HfesOahdYu1HdzBmrdP3PANFmjPsiFhIhTMfS+e0xy5rEhiVBuQ+5
0yXUH+u0dyAhdIpBRMBHTfUj5d52tEj0s0vFEA/Sv6WV1qY0AmBC4UUCfb8ZD+POERgFsoFe4aJt
wrdO4AUP+Ys6zQLyQxtLWHaFGnWEwN/J5eGicJZq7HOiLz78YoulfQ8iZd8GE4jQvWZUHAX5Ba/o
qMRW/xi4U9odZ2uulX2EykVzm9iDf/waN2+QCTa53Gm3gfbAQqY7AOVKlOuactvRku2nKVdOoAsH
hIvTeebSyxInUOHeaq5NWQTZBzcLxKQtn5g5PubvXgpyVtBTcT5DAvKp+8m4Q/6/5KHKr4sHWgX9
FY54UogKNpmFv//1t1+LJGmN7zR5x31Gq8zsgV9Id6pUnmgRsBs3aS36Tf0ZEm1CbhuQJMel17wD
okX23CVvEL2bQXrspx8elNL8G6qkRlch3D7Q/2b5NLSjKsIuHoRVSij41aAymd29KKQ8H5p3v/zm
BPEPWtyVujcpQ44v5BajNImgEQJDMtxBuUuX8Qvw3Po6+wLB1NBn0zPU75I94n4dxlDdlXc3B3Wv
IqX5q4HfYi3Mx9FOF/dnIL7IQy+E8O3tPgk6ZPfaErSn14xMPhc1zjdiKcUs6SDRFcC65pNT6EDo
0uQBGj/Ic8Bz9MYrtcyxLP9Vra4TVgW75XOMiNzeeHcegUP0vPyOpu7kjaajhxmrdi0zPMoOY9ND
LdlxxhPa5f8kaaufA+Cix7Pdmk3bEP+skm0VAjevoMXNgbdsG/8tAmWbrsMIeoPwT2fJSvVl0Oys
Bt2+XzRk/mlFxfmVFaNs8QrY6TDbgSAScOSB8foT9rTuOReF5LfYGexC5gDfsxW0yXoaVEk2db1g
Un/y/LpWs6Lo69gN/klM6d2lqRwASmYAjQPzAdWLHpS0UcBwFXm9MINGjYQ4yrBOPO1ZZOHYEDcq
sLRsT5ZTz94x8U9ANU+/F5jvT7MO15iMMJrBMuEYXrqHMFqnCqMYhTNTNh59bYedaRWZgCuQuK9d
1iFNg1kfUeMyJdfkASBX8LZMWFO/5em6Y0TjXrePWdNP3Tsr5Fg3xJq8geUJeKrHdFmqk4pj4yo9
QOo2tYhdTgCM1oYxc6hFpTeBzLI7FXcC/f8OAHkYEq3eGk68AON5eTAaQM5gYdHGxFvJVX4u3XC7
9nbT7T4u1z5Vw57ecmUYz1ZrWWfOPjz05oSywze5x/YpcKudTO7OW/XNtnmEIOF1nSGkyuxM+KLF
WGdbDf694m7iDW4947ffFOVODVlBBcrKNe+WkVCpmjy1lZThHcnRJXl7OiJdy2ieN9rV4OpIOnbk
r02C3ZzH/yBzsxjGAxragYIVt9BfKeXQlynf0AWKRNJn94RXzWz3srDTDYaLHfMk6Jbc0FfyPR+N
XPSQeCIB22i+vmLDbEfJ5LWlTU2Cya1LC7t+QD5DDCeuHFa6cYc2E7SdMomHjRucDhcjYVHP89kv
2fGYRWe1swvqoh3+JXzPZc+hLJf8VNqNMYbu3MqM5zwzzjcjvJbjk2unBKr2+YjumF5br18MU5QS
Hh7gOzQNX5tdl+DM2rAY31J8y6ns5frhKUc5Pv0tT9BEDPEU394TZ88ULGO1sjWyckxn2cf+n/42
M2bSo40Ofo5oQnZR0Mokt+uHUmq9Xh4WSD+ckTwPeS1qbHT3EYZZcaGsgTH3fNaGWZRwiSgMcZ8K
RVx+qVU6xc/o3FCif7sz3wI4+CPmQEzajIFodFncCCNcMpe/4b2od0us0fb8t6tFUZLgEPMZWn1a
Lal83rLAX01OndVJbV3yznMalRR6ttazQ7q1q4XGn/faWDSQb5miQaQSQzdwbht8OL071hgp3PTb
2QvWRwz/3uIGmOY1RW/3caeF9iLLDlYOxwlCCMwA5xIK/IjCZzGUQZRWMOQI4nlvnwoQKtGSFZfX
bvNjpEYH9Ice6xe03ZrkroJ/CEtp+TcZCWG+EC40IeVDzPNZ0tC3FDZNWuWZoDMjdDbsyearyUk3
UvW3C5J8jBbeXBvpPl0SpUlg/TLetq+7K14I9lSArl8WoSkucXjX71ulQ4U4pJVZL+tCiQBZl7Km
9CSWAtjRzcVqLcbilpKBWa0xXxg9IPVgT7CeJrKi1JzCYLIi/UT53bJHEFllls++qBY2Xv4sZwDb
vGjwv33oWo7wzJefUBsEc216wpBYpClrFeBlhOFNnbtukR7vBSaxO/4mx0Ph9IDofDWZlPDdcgK5
7TdBM5j8zJhgtdrXKrZLc+yqVS/6tppKFgp1SEFuPL68NXUq5Y5D50V400f8ipiqILVODlpLnf2x
5BSJ1NVQQC791Dc4HOFFFekAw/h1a0fEgQ5QeT8+VuCi1SPPeycZBqSogccObrk4VNi9CwMKDbQr
nR6+sMUrOdAbK1Pn6POxfjc/tcsrfnv9i0Ci5NzafV03WdQDYJOOqp8qqV6TdCnDxWB9SKyLtO+S
MQI8Mktn9XdGsusGkkjB67NP9Ef+FSR9/i5Bxa3a1j4+TpnczSC63wpzJAsDKaBQO4nYafqJMleq
O7+RA9FUN8xBvy89F6D4l4RQgCJuVfePu5p9JkJMuybPKEriQvp+6UCxyypTzZVCy48z87M4ATKS
wQJDXi52hfJ1KhqCYSOBo45orqoyd6cnIWP2sDl/RwgBI0YGtFLyNmmUJbEqoKhGNxsaJwbLpiGR
hL8KsUCGUkVvkyOPPrfCc5k8uPctTCeWcm1eWW0W9wjcT2ASzqVMchnHsjMU0EgvnUJebnZAXU50
a8kgdcRF9Ff6XNrmr3kgXpG+UIyek3a6ncF1RTrFj/vNQX+xA7SqUtY90rtK3Z5RlsS3lB3G/X3q
VT1IcwTsy5vhP/H7FqZN8WEla7OfAHrMVNTttM5dw261lUI5vjN0NDxq6HGONBax5xPIDuk6A/LY
3pec2pIRWhX6nK3RW/hlpY5D/0bNZ91dhbi4by8fg2eKfNlFU0nj0r/0a2r2inG/O/d9devNIN53
2tIg+DqTC71zZQG2raEfgw/iZ2LSAihqdQXbdgX0Qe22ESkbRf4Ppcdd1eM3usVqXwPZL2FQLIZI
WQKhsBf8BayHbzXvgfeumYqaVPzwIq7e5FehzLZ/0Fy0imaUpVuUULJelUBFUUKershNp6Uwf4AX
rpLXAzGt1R3vihrTOgyiOBRgL3iVJdtYAYzRri+rvxG6Y2TDWi2X8rNwMtKfEUCDxUdON6ZID/As
ZmhUtaVX+rLOmzrOE2DId4NB89wTU0/rkH8NFwW9EZn/5NhjN5D31DrFuNfJC5S/jC9frWl+ZK/J
k4lfoGjPdX9JlGkgH4MQ1cyNHWtqSQ2adMGoNjdxjtyrNl9zW8plNdUo/VsqiiqYywPjcEtC3GQu
inl++5CLuYIQJMhItceXOLEM197rlsi3mEchD8GZBQH1bzypDkZPJhDvR5NLaVH6I6wFO0WUeyFE
puLbr4ypgct+59zLMmcU0jcXz/8FHxBbqBIFlhK6Ijc7xaUh0+h3bY7Ps3b+2+uTEJ0O3eFMaXE3
kqCE+4YHuQCZ6jmxugurvpUz1LMNlCk2RYvLnR2aKW22Ll6Kb9JDmqiYXDRJJdIhxhlWbNc6jT1N
/GtWpEDlMxeGOkmhUcCNleI5YxhFygd1GKQEd39senJ5H5jwyZvomPyZA3XS2ifT/Oc6cQlqXQLK
Tb29ZN5fAUK8KZk6XReUYUMS106tL6/5/6IXIHwLRj4rEbatOU6PLg+LWexYXOtlzG/CbI0hP+6M
9FWDnG3jCwNj8A2G7CIb3uTFcysoC4vwL+kMVF+KcF5PtlqcRVMQiP9oBtVJTFNWsxUTGLlpJBqv
6J7S7sXa2aYA3ldC518qtenn/j8Pp1YjKCBOGk6PjYrdR36pSfY9VuMVKjC/zHjxz0ylG/N7WRNL
AUj7fdn0LVzZEIhaPtv0hGfjGtZnNylGTX+5QJUHWrjr1++iYp9CE0jFC3J4Q+CpqaSIr2liCA75
S764WoLIsgMZbTjHrdz965m0m0OqtlqIIw2nXMD2SZiOzY9lKglBsZA18nzlR3v3K3sygxZT5HJR
K2iTTmi173yDj3Sp//0TUjPC4PGDOakgLiBswIMsqGcfNusnHn+ttXhPwFse/4it07BTTC6NMkxp
h3YFv0KygAhBAKRrIYFDCSLDKuTtlpmQyLAHladZevKirxRdUOz94oIu7jv3FEUXKz6TiNrScku0
QYjFtbC6xQKocBWdZ93my4cU0tJVLWb61mfL9Ho9kybOxtaUpza1k4EtyFOyCHRf5+gj1/JNyAP+
ld8lGmnZXPI73bRLAvF+8+SxH2YWdmEw+eEdjZoIEQGjsEr0/WMQUOIWSuU8TnwIGVTEGwl6GvlO
0x+1X7cbBPP3iHDydr0fT2MceAUNvonGNS3zBJopIPy/EUcuELNyq72OR+7TlQ37deGgaO4403jG
4hDBzgWmXgKUgqKAugSC0recnGscNX2y0D5bVHeuKMOUeXQYb4IzL3ZH051CPpCM5aZyh5GoNevO
4xkZrgsx1UiIFrz0k+WVoDO4zmPdhzHgGhzGQIoTTxc8LnHGL1cEH36ZCdUp95NeaqxirpuXPRV9
SgYFlDMAAjL3FZF2y0HcE1UrqXxK2fh5qRLRZLQrKJjTMWH+Nt2aHMbjxhH5ONi3KRkoHF3R5MZj
fOpSvL/JVmqiwGLvE26Hxo5s4qvK6kLpvjaSuOu7uE8Fj8C/89zh5NhJsB7uOyOdiqldrtlllXWq
8NdcvzjnObpMBc/2RQ3nMK8uJ9aGu2cJbA8BpzAgjVwyVYvY8m5dz7/QuPCBKYtID11PrLtSItiH
F8wan1YC0WDx8tiAZoBG5ailqJhhKSn5v6Peffh60osGFo+9lh7sa/ydZAhB9qaG8IE5BYy4Lw/+
2rXSNYDE+MuZGYLQ04F3msVHPAsjNrbRR9uSydwQPBMvxoodK+DoBweF+lN4PueN47S1MarxErMu
vUW4SCxarimALsnv2EO9U8Fev3zxrC2WZ3dUPAJBl/PdulWXniBnL+/ksF79cuRB3TSwsa5d8E2g
KoUYshpmaOM59W0qjUELL1pnm6Ssy4kfDGMuxgcxCYMYRMz9VCBRsHcROGx1Wy6Svd1GYbM5XHxg
id0ZrQ0iC/uZvfHvqiGNmk5fxiOGHSx3XPD7/eOt5ECcyMUm6SvP6+2FkQbhWa6hM5u/K7fV0OQB
ba3lgxwF/6V8YxFsw84++E+wBpISvJY2Q0SZM01t0/F662X5Ng9UVjSnd9FoqRcnZVt5cmAOhb+s
KLmSkIZZZuJ8pDECTcvGQ8WFCy2RF4w68SL92rkLrcu6HZHkqMBWa3gjM/JghiCVKVXxtesRiG0q
WU8EVY3oi5IFm3Sr6yURHzvji1mY2C2i0XtNLQ+SupEbuWKF112ylprNDGKSIez4eUA02q2wMx9u
IzIvRJ8RIwNMj3zvnubEXM4iZ3avJzMXWeIWWbJiVwfqXbKDuUnC/dT6JEtfdrYSzx7vV6L5cuik
0KUUjB3CEKOUeQhJaWeg9lkTt+iwC/rBq6Z5KBRppk/4NoHNsYOHi7N79DyMkQww9D4KZ1opVNbR
VQ16cilaw5lSo3I4K6DNDrCl6ulbiFb39Za1VdsjpztS5w9zPPkUCLW8IhC6P0kUNtWXwZ3Y4/zN
P7N0I5hDyK3Szi5f0lbzk1d3gc3mHy1AatfAhzESAeBrTdbciArg2O9q4vMPcaDjXNlXHswMaCkv
SS6eM7nSWL50+vwfYsy5C9hg1JFFWHtYM2Aekf5s4/VO4nubQkxwEOap3U8OmRumz8HGZJXWeAFI
AnBFYhK35M2Zsaw6LDx6AXn+l0n5cC9xbFbVDPwo5d37fWaP0a3yoDmi+ZxFp0rADlPOxK6QJJeb
gOGIQm7fOFvAp8ew2C5fB3uJi18Vs8TqM9DdyB7MgEIAzv1TvNRNrEKb5fUXxC7RgCeegGe1Up/p
V+E2cBFnNwB7U4M1YwTMo1Bgcl+gtZF7fLZ+JO3vie0szpZNR5w19IRURc+rGqERFOSe5KpCXCvL
ig37Onkjt1ibSPi81d/9m9JRIN0GhrZzuQ3Avi4/GhAF29nsIzUPW0NGQ6Oc9T+arPiI2IE4pTIQ
XIBOW/+ViTxIjuhzQ1fwg8JzT3PG4GczWqV+4WcU8WYCGllxdoUMDghy/BLy5ympIBg6oybz5jW4
aHyU0L4Vxxbs/hUSycH3mBHL8I0sE1EwWX5/YfzxMj1wXncaQWuDjjgj7ezftnY9anBnm8RHL8xt
bwRjcW9RrludTlP8xE4x8PWinCP0hA1hGMMzKeI8MDg9/681UaMphYxZ7Cwrs0lSpu2ieYIA18+N
1olBeYLVyMVl8QSMF0BFTs5pR1YgWrUjA7ei/S9RMk5e0LrUTfn42oqj25I4uVznwmpjikBVWiI8
0plcZNoZ0kCOQ8Pv8IHvwnsYqjIpdvCps1shZTe92HX+uPvYE0t6lq4/7Jfp0Nzu2h8nrHiWrBoL
BBW4DlkcsZEIFAr5qFsQ7SBVEYRn1Bk2kz83tjUcdYd5tZ57vbszNNWG3Hzgqq81jrqibZ+t+64T
d3Emm6JWIPLWarM7hLWvvkhJG1oxYwzNcM0crijiL2nbIKKfLguYl3XWfOf4pEx4peOPuZ8NpxOH
mG58TVaMjYQaZbrOK2d5lsR56YcyNA6P9iY895LvL0QJ9GBnEsq8ZgAI08aXWR80CNZelWRjmEeA
2btVyr6Fok3QHg21jRyFS0cxNovt0rLSoakH4Y1aZKgOLVDrvLN+S9EwZ6UcnTBwzWCCLRLRJAFR
CuYBnar+bGgkkRMyDfssGcfTOZriB1XzSDgkfJNJEb2I+s5HTqU3QsmYb7UG5DghfZRZvL07spAo
ij8NCO2MJqt5+57POlyJGYDyi/Q9fdfQ+s2Pm7pDpSqwNJ/bbuarVSbOA6wwfX5+TCavRXkgu61S
RIQGmL4NDgIj1ZYPaH4sUc9K//rDKQGhAOws41AJbPyMqriqyHYBq++KOc9dqVjbsjCVpNyluprm
NXoZAUAKw7wS3WJjp8xIkrsWlp82p51rjOio3VBXhbBgUFJgutJ5p483ublqk4DclbKIY9CXMktO
TCJM+1Jd1aTijgZBIYU/AT/I3YazkSBRS6qaUyNwdCVDybkIzFjBkiSaB6025Td85H4cL1two+Bd
Y7vCts4NsbwWEIi5bRaeAI4dHyu0IrOAPvCReNYuWjh8V1Yqsv720YEFqHdmnHNWT6n3C5dKMK2d
D4Np9puvItGwrl1RmaYY9c+x2IRM4/RPnDEADDgKXibSRCsZg4FdJ3NhNH9TB0mCpZJLmGTUJJO5
pibP4ErseP7JpzratfjJhL+aue9HgyLPPftS+CEu1p10joUYLIGdE2SOM4q39G5Z7hTkVS4fltsR
IXi07LCbvMcgzE7TmV0+DsbsRZ5c4EuKydlGyWRh0CSFKulUbW5xuHlYjZ5Ls/OVaeKKP+4LydWd
XWIr9sA6oK7UK7peZ3kVq6q9mILKD6u0z9TL6NHWazTRgRZe0A3Gx68/LVTcLn0XwaptH3m/2YlR
6OJmYJ7luPEP+OBv3D7ULKKV4/suR2OUohjV6mb/adeGh5qVlJuPAPw2wf45ePNNfVflCqI9kAic
jfyPviQK7yYJM9fUKTpjYWE04G7GUjhZMLJ2acmR5ltFjHDEZGwNyLF/jQQfeTRK3341B5BnBcNb
pvkVFzv6QWW4rx1XI6jPsop035hFzboO/qthh5QrG8OFawrF9sst8Q+uWAaGaWDvQdW9g2VDYIto
ntQe/FKULX+h80G/hlHIN9d6KO0WrAqoKsodaQ3+XFgit14igVkEn3A1cxyJONtuN+VA6b/bHxD9
Pa33qdtVXYUz0MXUzPBYqDcFkizRNkKS1MUJS85ECt8jFGu9qirvXLx6OeTvRiTIaNfbPdt4yYQf
4tkvOrP2oKcoOy0hcoc9fMopLoPGFEcIS0kOvYwF0DHidsOCJaiKAjDJ1oNbiDu5xROyMM+4AEEI
+tcEnfOXrd1VstqX2hbcMWa5IU3Mzo7BgoBZ3PpJGABJn6R7FEPRMjBIvBYNtGtbjE4ABXyT805w
kTaoUp3R58aL55HVt782z7yHnfWsYN4dydZPa3mhqNHuQ7lB7Kd5W0kazh8653Mk6SRsnHNvwMTx
og6AT5fagBjFO2O6nhyKnPJgcMIypT4mTQvR1hG9m4H7UuONk7yJiF9458+CWM9gEYz62+a5IiIu
hpPuyfNFk52OQkUutWumDQQosxNkJ3WVRsKris0f/ecRAE/ZlxPzfRKLVIN0h25YGC6GVSbYwhbD
uz5brze3xBzshqd9lV2A/vlNXymiKGAWBdo2l7SXnzd+gQ0gxXLXl9JSmudkFicDEGzemelfkGj9
bY13BAYVjdX38vHduWjlL2+UgHDnzzRTA8caBSLUIQj8YQZMIgREjmjZmdjZQegC3qd/en1Ti2li
t6MaQub3Xcj0dKkYy/VTDbRVmV65HbhLh8ZWbjKfuw4bD/sqio7EK6wKPopREHC0ob6U+vXBXc8H
MnWHW4NX5wttndRfiRHn50u2DFHrnXav/rUXcQRUjtIit5hCrszo9KhPli4wJ3rv7QbhGM3Sqvco
tPZBCSw6uu2XsFSKf013Zv0h7INwU6w62gfbDEariGvQUBT+dHs9flby+6ByF0CCP8i07zIUT/ea
WFwt0VQ16not4vCRnSnYWk4LtFj1kejlUfecsRlOFu7LLzWTS/kNrxO3+jkWGbm8MLIbRXVD+fgJ
BgusVEHIAOmVJzbuQnEPV5hlWIf2KInuXvVa8n7IE6gBpFivBGHZEKb2pvdeie+ND/AqqxjjXZrc
Zmluytz7Rai5R4jgRw0aIQedsA8rfgOHpEGBXqk85X5uSwnQHyLr/IBUCtxpRIWMbuM8NTNgsSWH
j+x477+UZ/kMZ3nJ3eH9e9oizjQvsx0IHmaW1u2nsyDAVf4qHS8gJZyvumu/1Pw1YdPZUTh8YyUH
L8AFhXUpdyAjKwJpOF4n3U7v4WVNEAtE6SeoYrAHL1lETtt0K+m7LMv8AXfkYCGSA5NGgpPe/njO
FFoLXavP1aPH7UihxfdKjyuS+YgAYrZ3WUDh8NGdpYoHXMSEAIOyBVyuKbFz7fq6QfYy/9SMTkxv
n31l7jRIPNG645dPducWPEGmY8OI6WwMzOFFwYweAfX8rBmniALGKgRILKvXkxpQkPXCQMCNTexR
9dvSJO9D8WycRXqMk1859Yezc7EcaUBT5RqjnQ3Cz2A28HQc9WgelklTbl66ke0C/6TgOOxYkSf9
lL3J5ulNIdE58DZmgFh3Q5B6H1EOOtUlcA5RmTIMVL3f0xOpgumBVwxuZePiVfTqeCc/oPdxX+NT
KlXWHmbPkpjmVAP1k67CbmELa7fS/JUDkHlLyX1n8AHumA6vQovkGF/X9OhgfXWcUMz/z763VIES
TP/F5Xw+cFHh1cRuM8hf7N3w4IRb1+q1TpUsqPQstYO53UHlJXKurQ8tSRBl/MfoOpP4NjUFz8ZA
xhb7St/0Ur3ACI67eTxf0ZzEYPhahufI6vVGj+hsXw2MzZnwfmb35woa/jCUu9TQ/IGSjrFbMtzJ
niql3pNIg/mBsarGdT2vz616XvOKBoLmygUGUULWNa1OvNRExyQNQ9IVwuAArJ5aH8/1m+wXQrDn
9rmX6Ki7JIOGtV1koPdD4PMiwfClXhRyGP3eMiFICBLmWS0KpYAXZPJGgw2cSPFf3PUZ7lF8lhyI
BKPA6iCWDIT1ZMFHn9kqI1SWtDpohPEP+9OlE8KFi1LHZ+EO07sONvv9HlK6pDszaXDza0ectwoM
XNv9DjYwcZWRQIiS+KeifbUDS8YXwweZROIRb4PsNG5zlPsUU2TgqYcAAPCLDbKlR9HUvoEg/JtB
CUOofBSMuznNtWHB+IeSU92sf9zN0brNbTth6MfJsCCyafFv1altF9YwBReSpVdjJq3CCWb9SCxC
DVZWc/XGMOeWpINudlEq9Q/qeMP3CrNK03jK0BSt7Fxbn6DGrqC+aqeiR1ezM4nHhlxFMosaA6U6
V1ftfzrcd8c9iWhIFQD8WNrYdgPY9i6+C/0nJWZmUwsanKQerXV9GVdjGDg/YId60MdE/u8Q4QDC
K2eyos7CFPi7HODtN1VcTvM/JgtH9MPRHpgQ5EbGEJ8uZIqEkVIWnK0XVYKAlP+mTuXe50Qgd3y6
CHtenc7FB33kMNR1pgYlRPzOoMtVnHfZWLScydWs/gq8xJzekjzJzrwm32iBebTvPgwk9m0yQR+k
7wvudBMXd2XK3ypCTF6Rey/UZrI5Ah6UmEOERK/3qI8uoVLO0zYmnjB5bP9K2EK6iGdVMbp5hYCP
BOxYS2ORhkh7SMGE68BJOoNMwrmC+8tg7L4+EKjRx+ObwU1ZdN9cTB3pnlaGv9tT8MMQazzmrLBv
WDav0fILJ2dtyLIrCuMiCYF5dkpu5m+mFhO0MCC0p7HjIPVppNlXv8DZ4ocTjERKPIqGsV6kZ3ms
b/9Mw5ljKtJ/49Jo8NIeNFAmGLIbCO1QsPy5C6RaT8F//ditykfxPxK/DqZdKSvyWAdfvVNMl/hS
i/TX6RvzbT5TMqoi7icujVn+MnSJ3fAfM6/kYj2tuXKo9OQzdS6AI3R+tVfeXThTF7qDC2vfI3k2
7Rq4W0tB3iOs3B8nwTa1JXNw2d8O5/3KlBiC3T3BGHysTwJFCQ8VqXJn+LZh7DL4KCinOop8PphQ
YMvMUTDsU0lsv725Zbd7Bqn9K5k5auDt4jik7LKNHTWlOLHXlyrpaJA6OS5IpWCfMT+EMqMELZbV
CF/qXZGpOSdqOtJEgsaYfgJjsEMrLZl4ZiTUbTpI3YfSOxdWS9uTyD0wBHF5vZLVdZg46UP/IbXZ
EdPjDoCps24d2345Aq7xsJjQTbP/j7xiT/5ABrjJLLThJ9v/WDExskb3isaKbFJAJMMqpp873Mkg
9RXd+TcaFgn+qf91wgbsdAQnP4oXqwW5Ok8U4QUhVQGswlvtpb4MBa3kvQEBGtY7HM7cvgX2LbS9
gEbmv87PW+u/pfq8jBF5AFza1oTvPSKH8zf5RhjOuJDc01DhXpgenNMGzbCqFO+8WOjxV6+Z8LTx
rMYa0YONU96jxy3H1xOQjChJct6FjC4wZhv9zNryvW1eVgV5BQxwsOH+fXSUfQy529kBWkOrBX0Y
BQnC66mbHtKeq1el3dbdZhpj7NGhWTRof4fR4jpsWhCCLcIDHAX7lQZ2Rw9SdQCzQjekSj1GoMVg
7ixUw0kFfgcULu1IJL5kO/DO0AkRr5RYxWIYrobEkI5H/txI2MlYE1XmerQPQHKzsIT3ku3ddfuD
gMqgm3OiKDX3wHkIS3FlNrpfgtkBY7d1JjHN+IggHXgOK4nDnNQVyqduDNMk8lUvyJ2waMv3exfS
HSUNpS4aOjTeLZO/eUWCesT49WiygGuh3rqxxthekyKd69aRItErzKPU7+Qockh1gw8i4I0wJAzZ
isncqVPECXnUcDA83il4HctQNij/VKAJmw/CUjC/RkRWZfjZ7JDJ7qj2wYsHx8FwN/NnVYw4Fh/v
8U5XLVuusywPLQpj+tQuzKH3uz0tqJBHNGTkZCkPLJPHi6JR9HJN8uWgmS3Ou/q7nussEVcRwbsA
LaP56okcJxtspTuGNqfoGM5e9+kakCCn+LEcsNmyxiZvNkcbgLDg174DuzcAVOMvyrjx4h8VV1kL
lNe4JVU3SQG2Vp/k6wRF76UUzKND6jtBr1tYO5yMoNTarvXGWtS/rQBr2Tl98VlhXpspZV4kdDRh
O0mvuHpjHvP1AwxVOsbJ+VUEyKlLumGd6V0xwe9lKSKXp3tOAe/1g0Z829ByuK4EGO9M5V+ETtzJ
P0chABvsy9mkgzdM5sydd+SwQHzC501mPu+TdDJjYssLf/DQuRMrnD4uZd/HWsmrNZevexZMVGXL
UHVBBIEGNaPEoKQ8mMrKXoPG3NImloC/Z97PbaMqGyvZhmMZ4kE2LqlzSzoNukfjtx5YlgcN/g2B
3aweNX5vOWh8GSQYpzwGTPjWua1rA9KchXC8EDMxCvYezsadFbkSNE7d1JcQ8fJ852Nes5T5/R0V
9nXih0tXwKdlkQ0R6C7SdrQ9S54KoiMNb0HQfng1sILk3xWDegnuTUjEy4WkZYdUeg6PGvCu/F1T
+fI9eXL/xLdJA/ICd3jm4oo5z7YaSBGc0SM9Q/Gjq0VdIzWvoPJfXDTO7NGidSCcVt+DplzNGMPO
m4Ndg9jaPBrmriNNn8VujWf8ZcnerOFYg7zuturzZx9j5hBAVqEyOVznkNLNGxBiApga7PKrMfE/
YVAM7WwOP4IX7Z5VbsMY8tlnDlTZWJxG1YPZ+0tf09ZQxH41GcmOs0jr2IlMHfOjHWAhlDfMaXTe
qqAkxNYQvpJ27Dbjtf8PE69QzrSFnIkyRpxpDthuuSaKOHKOO7WQ2B0yKYNn04RVpmCPEdxEw3nK
gfiUIXuKqjX9xqVwGb73jD9jpbAa68bL+EAJRnrWwQHmPxrus+WjBHDgJrei9LJjg/cmgvwKiHEF
EOtsEgpr3kx0kFL7rzvoaTTZtad6kFvVfe2hbZzPTYENQIPD4MS2K0CTyZ0ZS7Y99aHC01cQhRq9
rDJxExxvHzaFYd94+g7idxwV4VyxgbQXluH14mTliaYBRAj4plIrha8TTY/qQSHW+xbJsaFzjD/+
xcLJyGyAwnFx0EjdjN4F/skIxZXcEiCQL8JrEgsSDh+iyHAoRMKvPBrKzqga/taHTXqowvve+YQu
hvEbgAA2vT434yUvlWQNgWPJ/zySlM+EtflnrKQXbTqebD7RSPehSqYuaqcq0qE4vQ4/4I8V3Z6m
LvniIjDvoSZA7rlJHfoP4Ku4D2A0c7/q5o9fgXv9/BEdsQ58kqdK6bReSntykGbCpEHteAdIwrla
jhdKLv5tCpwVsDVQmeyKq7picPyJgc04q/v5adAXTLeM4dq6fu8jxcc2b6v7yYP6Z+960AWULRO5
oZ4OGSFZf6GvTLAx30kkK5DkR6+vD1r9KR0mWSENDChu9jW7rXB6YSlZoDPQ97YTgD4puu+NnyKH
kwcsTS504MPRhCJh30XNcJaQVMSgEj7sP94Geboe8CFipylpj1yzrP4nvjoiOJ+z79dRByhfC2+U
xwwMaLAatO7ho4utLisPbs+HSJluC2HMZY4dS/8eW14jr4WhsSC4iMF8YREh7odPzIg+3NGwjcbL
GjUECAYaiCXCfEhh73xxVBXh9j8Jn4QMHMzj7b6Ew8S3Fm+FSHD0RLCgMb+N/XpXS3jFfd5FyPiW
7ncuC7OYSUUHst/CYlWPeEpS/Qq7EXuLY3focjxoecwddjt0IOzdvZQK3FoTeRD4RAUCkRAC9CKP
is2tIE3N8VioAnoV3wAp2rlkybB5dqwJPdjN7cKVXVEdpzBiM0Gps6arik9Wl3v/7MmV2gBekK3K
OJFy1/VL0ZbjfHl/0kg6DIgHth9evXanLl3M857jP2zqK8fW6mnys//GNtvWyCRWBoPtj1Kc9a1m
iVJphEX8nXaOEg962Hk+zwaxOcsAdD5xMU7PUDx45Vu47F/80SKl6ztgW4cvHScHEUbFPBiJMdMZ
y80c36di6/tVMT7MAUuL3aWJk1hpr4AUD3T3TF6pdWJJz6ySD+X1Pp+2zefZ6P/LR7NjliB9zqDB
Hc4cemOsU8sVNSQGJz5EF5f7rgltfgfUNbIfUOkjtKei7Tt7Pg/WlR3eQ9meCcVD+/RuOIYAc9D3
HLvEZNkg0haVmAvh6sOg8BeOWY1smocYDtaqZFDjIxfTrPrYM8iI70lVU4/ZpSzAlQT2DKqdUwLK
upTjoqxU0c5xeMyiozeFTCAn63ajdufZKIeDSxQRAcyinN8uhsu/k2LInGbkLV2b24CAtmfBCZ5j
iPkjzQRd2jnMUOBS1RDQAZkrGxlhbI2YFNAKIGVKgIlFeswuZZ5UqRhqTN5dPMIDakvU0mbVC0uY
NB3D/nQImhxE463IcGeLxDxvLcCqNugB7N1BZKNaE+e+N/KxjrnULgBAcIvk8ad7x6hkRP+MmDCU
7VVoQIo6QkBmdxY3xfYsCxbQUdhjvAe2zZNnPrHVXd0uF/YHpc/96OzAPH8YC6WszGVz/sLAHhla
UJTapTWSaeEHWD1aRXUaR0BrgLYMz671pS9hcuyJC4YVNuOIQcDptNfh+0EbPizPg/rOfRMu5pVw
Td+a8qE92K9JysVJ5CX11wWyFqAQUl0IouxcGE54w3dojVngcQk36NIPAEdZfL8TdW2oKtyAHkOg
LAllE2Hv1zUebBX8Pnod+b0gA6POexTL70ATbc41u7VGX8ejRagDXZhVYrn80kPkNa9qqjBXPsEL
7nULsDs1U10sq+EHYNpzEDz77ahD3oL9tNdxl39J3UUqG3VbOMl/hfhmL/+55OtdgZnbjzrkYgWf
UgMjO87SVvs/B0zdkqBS84Ci2zV50D2K5zJbrazOYHZFSIiUJ1pdihfh947cz3ojetr4QCoYDjoA
r/AHGvmZWzBWsXMD3K0K8KBzT3qfsvseYKUqtzQZZQplHWAUGQzhoD/jvxX5BXGHgDFmefJnRV4F
fZg7CgHRNgEBcEhb9IYbdlLDNoq+pIRwwvDsgpELXwZ/RZnnmQ5VMWG9JBHa2j0jhxRf3sXkHMKJ
SC7VOCU4y0RRl3EiwlEikA/KIXbki7cH8aQy3yJpgQ0qp8QuS2QC4YviluqXb1siN+NHr+9do7KU
89MpFqGgQ+11eX/KHn8B8XUbbt0BH2Z3ysGPgXE30TZYDmrqr6muZAQPZRf86lxGAdeZ8MkCP54t
+MGopnV0zvaSfFMIM+Pq5m5+Q1JvdDa6IzdT2/OirNeZR1eX5yuJPStH8vQK3Njgv8S4C4gnXe7s
xbQKyJfm6mJYuoGLllo6wmO0NMjcAXq+PA7InjXq+N567s1JLT/apawbmG7EF6L1LdcYu7VCYoXC
NF5X7TGezV2KCdyefqHuoMT+a1u48G7Q9r1od4Xk/0cWwPuI63jUdy72V85ttDs7BvIyKX7nNrQz
pfMDiFKe06/CMN3rbOhAbVCCzdBXgGmJFQsKQYxqQcSXtoggLCoDSsYr0b7vLTSay5VwdrIBphy/
LJwL3a25pExJlPLLdRzT89KrmfyOYcWCBhzgOO192n4j0EGsOHKV4HeUqRfdblXbarx7UdF667Lx
EdwvBG76lOpNEFg/gB1Zo4iHUdPNpc/dp65z6INPHvR86onjZap2QXkSbJBt2ObKxzZlLPsM+cF6
bb1s4lkZotnQVOfkWDLNWj5/P14XbxYqD3TUTb75+pcTc9vcYTfcOgcZ7FCIWKh9EleUT/rZmDAZ
OJVPv64NGhiDFKokZ+n3a89gSCKeJjW2QxM9WJAbR6kjryBlRKmdR6Xo2b6HQS+G6eXPY/3wN2rO
ybabeoC8VQ+5h8ZVDIXFQ18Tpp97Loaej1Zpvjd1s+xE/j0JiqLEgk0umB1QuFM5aAVD/K+St47V
gaAYOnLu5GJ+tMLCJEpg2oQNGzBTWiOyxdXebZHigERmQmQVsgZl95CfsD17RJA+TYAKu6Zn6rWW
JGPufJXxYh83LO03RUBGWyDLuHVDv46eqtIBxUZJCK9AqDYzwVPIktciXjjP0bupEz4Fu0aD3NuP
+3SD8mIMYrkjm3H0eMMSzeP8HPBnlsXkl1XYtIUyIj8xO2suCQLEEeAm7WAj+uvUev0/KLdDfg2U
6NqqTlhmN68suhHhmD1gAfvKcA9uUaUDBrxH0/n2V4HJkvsmX4g/2R/zmTb5QCNkgDmKK3rSCZuB
VsqAS02cT21/6tW79Gp+s5uu4CAFni596hkUr6Q64XeXTU95Q/y1qfF+A91/HJumIZ74gNt4qqaK
CEhBCG8OAW1QQ6sxtOeHnofHOt1Y/XIyyI02jbOWcyx2f0I1/JNYz+3POGiYnzZj7LRIelhjC8Wf
EVz/s8HdCpbAh2czG5bRwhEpniFkLPQxmi7wjfhJmhZ8KYG8cjALxXKcyLifp/yXivd9L8zsG9wy
4nL1sX3H6L8G7Bnm+BfHaScozRgnRyXsYK7hNFXvTCXSCDROliAHssJIFI3G6MpFpE2IJnRpkNJk
p9kWfISn6Fur7KXmRqlGexj/O3q36IHb+tumpv/z/1qa/SRiSTnT6RFocLaJcdwYcAOKN24noaPf
oldFKpVjwkn8aMbHCeUsGyZjMK4NFENLod4N7XARzkyAfIlQ/iaBGvNTGV7/cowcrbMvCo6q5eBP
U88jqwh9/GpSJSXt7TsrZxh/NhAVbUcpmXfG+Ma4W8vE51zOYjlLKIzHPbUzLQVadJ7tXSaSTwXv
jC2jZwQPHZcgRfnZk73W3RdMxh14uVvvYbskmPY8Ns7h2de74qb3uP6X2j5SrZ7oKJQgaoQBz4UJ
QXwpUZFKUM1alaZssm599OWHVy5UMla5/4zwE6c8Da1zkxABFAOHRplVQlGg+hJhJ1Rb2y9biPX5
YrNycCdK2A5rMrR/4G5ZQbJDVSjoVwU4vmtSA9uXgmLnwEoRlcp5bleqd1ijLmWqS8JtqKZ+ogW8
fPln4rE+GhWmm1+O5cCfzJz/GKmWbNfwM50cccX+XEm6S1dCJc0IvGWOKT6yR89g2PblymDk4Y8j
J7uAlIdUEg8VEdwR4hUUsxZgBm3V4V4xomTsOuMjywlQQQm+ZTH9qMivG9E77EKsuO4gL3gaQdWT
3tdHGlcH6crVIQxzKKpyY29kZhOYVdD3rzpuE1RxM36Fx8umH3WkC2D5Fwa+l90b5bZxfx+UmZZO
xU6mBl1mw3WbCGj6ynak+KZsVlshs0FZEbkin8FDMpwPN1nHXj8ToKnCdeDEEdeLsGnmTMUAKawH
sKjTQnko7obJS5PkX137U8ZE5tTpr9AHpq4QCYVWA+Wxz7lDCCBTw0LXSbWh45RohR5mJmprLxNg
kUHFfgnWwOhCz73+YA3QYLt47KpkVoYVzDBoVPOL9iYx4RL02W2ORORaSA/vb3B9e71y6exXxBGm
XRk3H9xpTblYfCo0lv19A2/T6Tc2UOil5mPJ7f2q+TivGRl6yzVqR0Mrh2qaUYgOqbwaA0y70lTl
U+1UTvF9kkVXV3x65rfJXawEwgoNc/AHUW6k33tn6MwxlVusHWoEisSJfBp7NC581jlUhT8Pl/k3
1QRsmrBaeRB7RU+J4f1cet9UFr66hSJ1Wy9DQQclryJBnTpMZPArOg4tdoyhiJIPKRClguptWel2
ec8Fe0wVaN7SBLeNOwyGFtyG2lShHI1GoPqcMZpb8L+uAbHdMqNfdAXXx4appL/OcIitNdRLOK8o
IwDPw9SiwH7bStvIwPhlHuELFnyL40WolPYEVaq6joMknZuSs7Cn+0+/10nei6z0H5tK2NL8F89c
vdVaWhicQy6C0rww87kI6pYxR9GpfbYI/p9tcfRgGv0fSevX4LW9LbvRsGZXFwA+eF32YybS9wVc
GnFJD207vPaaFZFU9uOVmLi7ljoId9hbdwNGH0AfTod+7oPV2N88J/QqPwlDwkYIb46vUm/eglCl
2PqAdpOidGh+h+o5RJiBgWvzfJ5fLNznyWIJGtfRO142uqKdr5m8oY/CX6nodFvzijVjXJvyqJNH
/3W7LVF0415x4JvDCS/js9ZAuvxBLFtYQ717vGaSvV/MN9rHj4qI8ry7VDimu8Es2P/i7Wqejtv7
ReQ4Py976x5nVa6q508g8bvhYpFGpICpucdo3n/gZJDbfJQMqopUUmNDylLRGpNgKpYb5rczNY4X
VCLuielEdz5JrH2yQrkg09VAeYjrwNkpWBRtXwIbbEDAm4LjJHRzfigm2hnOau9P1AcMd/ctHnvp
Fj4rqQqsLExsV7atbuZmA0S04XfvKnBf7rVfymK8uJsaTZFF5KuxJyj1UxnR5pOsYjUjpIsCoHnp
pshmZblTtYeis5c8TgJqpxlZpLJ7JQ4YliCUj/2728M1x3poXXbYs4qSn4eFMdUmiIY3Rm2pDdtE
0lKwc6rCqC5C/kU2O0dzaofqTQAoA2QSRDiCbNOXcRq1uyaJibQD+QQzd795VqCgTgtbHQ3u7f4J
HMSZRi9l+HPy+HCa/Qjd8g1nyZPea85L+058KtS9fCzPg/+RLWDu0LwMHYhbNPQxWVuCudHLyBYj
yhdw6XrWJAUlOApagh8eflECexwHZTLQ8/d+0z9DJ0jry4OXNxdYwnPOVvkcU27NnNfxKkcQq5DJ
7juDmeu+ZYxBGJLAedMdgspca7xhKZbE37wDzQ94MLu8aOgU4Db5e1qcDo/Dg9HpGpZLQpEVsTzT
9ueL30tmvKHIH1felY7OTWxDcLTAyXipRtuL04GPSjriWI1/nVucxwCzw45iQxp3HXkafL1xjY3l
1RtNCc5agNnInFrkicqsfiL1L3RhD8sleg3Vfq0OHC07hLR+iQqcD5d0sBv22wMbByToCcxfOGyp
XMLshuKNj2eP46c6Kw9YzZdnFMuSQd8h6QEkegfPB1rQEul+ZSRzbfKDDZNYz/AS4sDozcreIDr5
XU4f/7NonUBV4NJN6ONsHiJSQyq4MVe+mpQhzzS0ex+zLGKpwkd0Xkt2+uK56UqamYX4etj+OvVY
PiD0AN5SQYsjn9y7kBAyCJOqiy4FN6V82mbh7N7tInjVHg2U6AqjDtiYQOdckBxj0pifLcEiq4Tv
n4hO3Cj1yboZhoc4qw90lciUR3LHE51thKTPrvHI5UFOjVNwl0d2lI3v6G5jzUdTxazp+iDujdqy
tBSX1HduQKb+Kg64TZGRQrEU2RFDtZaA7UER35IcMqYW3dBch6CnEgwrqtoPZ7qovoTZbPdLmUu3
t47rX8X0Ged8qlRXJVlPVClnXwKBJmQv5fDmB3PzZbTMLBHlllw+IH/59MRhT1lbsylR1FXkUrtv
7zEdDea0dcv4KCfoEE/YeJE/KgmTef2Js8al2PBOGQcBBpLChDJeWrAnqWXLwyksiNp7zczTgFMG
e0Aau8z0l76lTEq2/+sJqLmnWko8gNbs75ILLjy3WI3EmwbkrFgOsWYzuujbPr9IDeNyB/S2ctng
coFZIs5QE/pmG7Eo5LPrY7pRr1i9Et6cHSirZ09P2V5x+3ymPHLy22Z7rvSpor+VpK49zj3f8XFa
ut7MT7Qu9/M0ajclquSR3Yn5yYkNVapKt6cE57exBNmuQCwv3kzk/5i/kwb9GnSvvbDnEZKQ2xXP
JsDdr34toDQxiE3opvkBqQJaO1ovqyUOA5Kt+dcJOxPIfkJ+/adI6UGDEA6v74Cqg/gx6Xm603MQ
BAyLd4ldLkGgLpEkSrSJ72kXQYrHHbZcHJNU9E1U/JsM3y97XlbfZJ88OryFJ+ekkaxM6JHYhBSP
/Em0fxp/4FFUDhiIuYWIKpEIHJt9nL0YMj8/ysJ7Jn9NDxbTKwJN3idPPx5CcWP54QTaahMdBoOo
8TTmxkVErHCyQjM/zGbZGPKg3IHz7gpAetwfEkgK+5y9AzSA8Njj/JVPPS/GhLkD1p2UVpRQetnY
hwcs1DLncLA+wFOuGbnH0bRLqiE2VSz+yZk0EqJJOSbVYCnCwSOKLf5+c3CqwRF91PgBuwUWeiDP
TWvYuBp6Erfsys/UXXrJZm+fuxgtWezvOCTUZY6PrTRnrhkd0vztaEN5ALZ1cV1OyqZl/5Tii0VX
mxGWsS1BoFfqYedO7746jNOmJ4ZPGrji0nvqbeynpIcdMhkrPQk+YLpSwoJ7E9g4LHu5206emgqT
xBSlftcEm+dYQI8u+QHccXj+s2O/94UTiNKWqASiOSinJdh88UEWZ6xTM0tejOKpuELqw06X/0Us
fDqi27eqkJqRgCFyPFA8l7dUubOcqCi05gI1TvijL2oqS5J3xBEQ57siysi2YrT56TkcuWB+rBpf
zT3+HWFnhlj3Yam7Ljv968t9mNVyVPT7ST+r/EZz3rLt5T2AQyHyDEv+hES/muUl6k/7ZNC/iXoH
pPcvq2wYBgBYJY3joKzn4dRapgfMmpln82MoMUvTcpcp0pWks32Xd1RkCWYhYNGjUP3xNhMD0KYH
7ttVz5Cxn/KaQpVpsfiIrVnpQK+Kldrbof7Ic+1fIiChKEQT4SkBBKR6f4JDSBjw/F5FRWFBUByo
qEJMF3GWdr7T/MTM9KjGvv/DSh9bOMtp8pOIn9KIphw9rXkAijigbR2Be6bppV6hHu4mg0rMoqob
RsgwgMGUHvRIr6FInIrP+sDCCRFpovdAMR7+QtwmnTSKPEmp18PFMmj4R58XZpIlZYmtIWeVDr29
Ve2il3gV++BvXhepwyZZtgdYjTOLOYpGQbXvmrkKUbGfcyJMQcI8c3E6DNtSWTw54z0fq77P2Hbt
9BG48J52c9zfH+stoyvN/btDoqaXmZgVlNsi8VBQAgmOMj0a2izaujmdklymLg4rw97WxuzOYPKv
gmOGNwFaOKzIfKK0MXhgmh5Z7dLOrkUY5VBbCWU5UYHH7aiOLz2kWT9CRNTnJsWBJqL7t8WkJ7z0
BqaR9eFfkjhwIYYqLWTTyMGpeLe4sLyVxkzVIPghpQIsEGVv7Sjby+qgrfdjFfhQ6+oKUfAGnB4P
qSAhiuLxQ+RRxkwDYbEPZmzFhjkB2GPlM+g+NOhoj84lyYVnINdJh9KsuY3q4ijswU2mjFfz0aVG
ChfheZKEfO6NQ1xzTEVaNAi7ndKpcIa8Jxa3cbsfgfa15a1e75etkjYc916EDy1Yahyf1XUGncLn
i3xM/u6wSCK9uR6KExeckMOiniTaNBZfd3N3/6T+EgzN6AIHzNT/M63wTrkXo+ROaVXHSFKJyqmB
IgjALA0aT4nwh4AWNsAKMENU9XyziO8bDFCS6hglUDFRPGOIA7pLYJz4y9EwM/GHO8ijyFafM9FW
mVfcFib4Kebq1PGIpdGjgKI9/qGiYzDW8VNyCCdGT5R88XQrEhK56DL87H2aM4+zJKKnMrvOXYQB
JzYlQW3UZU8OdH4bSJ66tWiwuWEb60Fhcpt+ajtpFgcRtGJPrypYzM6vvOwsG1OBVLxHSRIYrLZD
dJ3f6mJ2psxEOtHHieMemFc3wY41d1hofbi1CoPepLUr/gT84EYeYfn5JpqNQ9ypUuZvNbr/BhMx
Eh7QZXfu7AeT2OVkMtkniZT+KknrkFJJx3AUkitiHmYiweHDhSXx8RgCJ4/bnT0cvEp1vE4v1kX4
OU5luLf2OwjhzJ23XxrWdhyVBRDkeEAu8V2UxQ61wPOvqXrVfWc+zfsMaaN8TgRwNARNOOZkUdzD
v2ATjB+a1TeyqyhS4S5w8DU5aUjPdtaAaS5GDzuGZADmdNNcMztb//J8vRtIh32YHu5Hdlz3Zgs4
nEAymeipDIIMkLvYz8siIDt07YPTeA6vWmOgVxc/XAAZrTGoQLb7H/P8FC989doUrG9XEAOw3jIY
rhYCe4A43oA7KIMaYjdnPC2VwxP3iAyVY5zKej+lA2B9hwZj/2l9eBuHzFWx2ullVwt9Y49uhmmE
qK+o0ydEK4pZe5EjQNPQteZvB0/kCfjXXofvSuxwnFp3wAhHZoujaO/hD/J/Ysr+8/5cBp9+1lco
kVcHVpyzuwgdlkvt1dG1aP6ghDLOMjw/uc3mta2aYCV9B61pY9UjWI4kWirseSbmpQSFXkLWbN7B
6P3nPQTIcB38qDCjm8DjJ0741R0zL9L1SfvqxIjQlfqSSCmn7s1u0SajYXq3yhTE0wNtSzlA9F8H
cCBceV5emgM3SJ4U/0jbXi1INN1LAzJMeLZpVDH8GzQu1oC/AooIHBpktDWiJshSCMdugG8CZ4IE
+BPqtXfW4oRo8jXbcq/3sMwr805NOkpu+ZQz8oqNFM79BKuo70tEDSp7VBira/LHoWCyI2av1CMe
BSoT6LD317RgJFt6zmtliFIjOuD7xSXmaBoS3CSxivuEWT/3JJUhVVHly5hfpzQG2YH7WjOB59na
oT/lDOios03WLJKnOFMWJEkOP5nR74tecIftpwTUg83b8I0XDgw0UV41X7nXzcZ2ey1OH0a8rBFP
GUuy199LIvCEwYDKOLNu3gi+N2oGrCJrJD8GGBot93A3uf+y4b5XCMtgjA667LfvNt/UB7qfFiuy
LreTNc3RPO07ZKv7CYS0ukno/A7yKv4ooI1cQ4RQHZAFms7SC08F6/QyVwzPXG5F+VVkfKJb7Pz9
nPFHffHcf/C5g3j+gJgIhhuIunH5hR9LuYPFL9Y+DV5EP0g99TgFFrvenDUjg0Yb864Qv7+XO36W
DSUM8s8M5/L/BMzNwBxrxhVuE6kTcQ5hCuM8sXG6/ruwLBtBL59UjsBfpKVhxFn/NSP9bnXAT7XS
Ap8B8ojC8XjbRif8ZDkkYm++P6HEFN+p4ttQl2KWWxDaetdQm/x6PYl924caLiDwuzc6D+QPw6Rn
0JIVKPDgMBrWiV99Ety0ewbxmWxtyRkjPD+swD8NAKCkFIiPGFFf4Sd8bvrp47lrVzejDVabr/bN
G5F5MXh/n6caMt6jCw7tZQ7Lqv6M+xNaZIHZ7VaIpJfhsGBT6tXm9DP3kRyqg0x8krBNKHF0HyEv
gPvwkk6rPe2JjTtiYSBQJBg52sVaeeDAWMYvSjfI/RAQyRK2T7F3gYN3sl96i2Rl3t6jSELI8bYW
IquqAEVTFA7WJj92N+DPwQ/NLMwl5lGdx3hA879Ep2FX9u3Jn5jZ4p1bESpDTXSrbr5IjTkfu3wN
b48Xw+qJpCn1N7l3HPdXH9kHoIEza/nm/WPxDcIi8ef+4CPZBND9qzbMq7LTY0LyhbX+K/0UJfFI
mc1X4h7h3Fd2S4IMSSkUvdOssOso87cD2PAowzDNfVh1oJoUI67Fq+miT3jI0d2Jvt6KJiLicDfU
+m+8bT0fsPILy9PDfCG2qxUAiMXwXO7l1iczeTE32B6vUfXDtPTTbXSDU6Es8EGRx5WFvem0CFcO
xkHikaFcqQfHHpzSIvRevdYjHZD27J10UI+/VEDmYAmoNymTXxEhEWMUIN0EWKOU/A1yTyk4NMop
A3pq7MYhcRTGJmuxxLvCPZxQ+mUKebJVvpfdAZJLmf3OjWb1skhhmYzoJZMfb4nIEPsyYis8hAEV
Xlt5LF3qv23KRn6quuS45EofMmPF5TetzWgm67BBDEIbJH+1ESTYPIP5WtgYdseHhFZSJQygI63l
dsoBU57MPWDoioY56JRk0U71KHczhD98U7TUYy7iRUT60jFd2CzFw7zpgVSn4GT2QaZPqd1L3DOR
T3QfwWfR3SFE//CkLB4mgZVbQMr4aE/CGX8W5scE2dC2M63A2H1DjNGinOebIeIk2ovvXv+/4Wpu
AT06ndqtKWQxFNJHBRpccs58VO3yKAgLK6SyzuFota8oN4DH6Ndh23yoib0+KftqGRyqYVY7q4ah
SaMFAafMHmjcyPgSVqAxtvJf3tenAAZFDM7hbxjtBZRKynOiCRW7G8N/F6UrsbavXesgwPH3sUDc
G+ulXSSv28N3ZKTHSBsDWjb1WDO0yA85mtU2CZ0wTj/bTD2CsYXuDdyz0Ow45eafPLfDcv/YYbfS
kgrNEVns19X9NG9vOzVMcXBZn4BPs7M2kebf/lVtA8CjQvAsap6WKr7/Q81lB3H7Akw9R6O/a0EW
H/ElKxABxn3KFY/oyyIXkGSSYoKuaYmdpG1aiEKlccIK57FDHErHKgHzWOpzplXinPQ//Eo3BtQs
XI3Gs7GciiC92/a6IiZS36kVme71uGreWaB/d84H20fLhw68JMpUeFuC5REZlu31Dp8uozDfVv3o
pj5KVyABIuNWSGLbO/MWkWK+Ht33j54Y23xSWfVd+cRfyfcs2yynVeGhciXvtYZU5VPAerrjanlx
BzO/YtbUVAKgP39JQe58+I1Go5v7Be52rFeS7jSaDJ/ufdN2exdom8/ctnQy6n5KfAJq/g4QCNcs
0OFtW7xTwE1aKKav882b16RH23UhcNNxveBKs1RKBczhpBSlmoC2JitsSM0KoSWohQKy9M2/C4Lt
37BEqAbuwGZ5sbWd5wCrxow9ZP3z1r/R1EOwFJq9fda3CyWoxMJUBNBNANXbutNGc7WY8W0ev8Px
oAtFM62Lr4+ER/hnNsaWegYNaaoWnWlPR31tu9Uu4Vmq22iV60nh4bpNH+aio7Rzy5zaK1wTredq
1q3Dcto8oqJLYb7d+lSUCpqOWkvN2Nz8aAvZYITLqwayi1uzQtl8lOH3o3gaGvzr3wgEl+6p4YHm
As6ZmJpKqhnBqtPtz1pLq2wDTrtQzNXQHd190Va2qktsOwXRMO+zq/5LfQLiHHlFgCva7CSR5wpT
C6V2hLO9kCABgT/mdgWNu/Cyr/KStR2NBADm42e56m5noYTJXT7RAUebD2EJ+6C5XbUYrIxjHJxy
Q2kiJiLx/2M6oNZc8X4kZVPYBnroH/u3tj4Xq703VFP7lOnD4w2uVd3+eFuyDev2LwE++RcZdXl/
fVuV3JhOwgEFmW1fXIblvBrcDcrnAhIhmTFaSrXTi5wXdUH2puJA+XZjxQVJgQ6L3gMJ2459XuW1
BpbdObnN5ihu2d8p7bsQBCsm28Wm8dqfFw7lbXyGpNWvT6vEPr1FbgwzWYZkSMUVVuoSfF1rf8UI
HBiekOZ0Sd3Zk1gqocl5wydKMzQgeIqxQ9yTwlh2ZfJhPhIp/cRWti32l5XtZ/ccTHq8YTqdYmvD
ass9aNLN/mUOtbPOszoFodz1AC2097TWgQ0yPWCv+r+1L0N8q+fdTB6a2u0L1I85yd5T/jHb3Bxb
+HuZ7Ze4SrCUgU3tB/D3IqEPK201NBAqSQX5nRZ+D///0RToGzBAKAeqQkKSyBlK2Q5uF37whxoB
CpNG+hieDVex3MkxNvQqehDg5hzazrwWsxrF3JBXzfsmpQ6cIXX/2d9C5B7Q8tHjZGydKN4mrBCZ
QpjyEysaXKBib6cHK18k+7D8DgDaKvSgwdzxr4RiUp/N5aGvhYKfQhr8f6AU7FziN2SLWIQPXEhn
uNteMEFMTheOLAVgb3/EsU507ILM9kMv3T40eSq9YO81dVL6rEE+X+ZcfWiJutUbGahx9uerL53p
6Q4kJ56mGZIeHBC1VHUp08Nfjv17ynvk2GUJKOOxqmNqQ5Sn+r+rHu5WTBLwg0dTGAVdowrpv/hK
pZ0knL+SqkjmbWBzqYPMNEE5AdNLmbQwUgfrGE9TeWBPh1YBXEp0dl8VLeqKp30jIHQhSlY0MPsu
m41qkNmqrHCQepVYyS4YLBnMU+drSQqB0BN3CKyyTNV3ue1zUX2jc+opgPcuNgEYR6/jsiaY1cCG
0utlONA2imMbMLYosAerqpk/a6wYZkVBktUCX/lBsRs4CHGCQ2h9TDT2CwJ2jUtB3jCxAcfN2aEL
9jp8zKhlDWKMucCsQLknhsBdB8242GhHFlBMFd2OgexoknSJ+PdNSpO1N+YREsxwO3RVZ9fvvSE+
2lfD4CvQJL/Mj5Q1k6snG0ciIgVTv0y8SM8KI8TxpAx3GeVWQM8ev+EYssR+O0SksZUMCs/rspUf
lXgoVu07UKdYHfqHIg5uhWzT3vui6bCj56XzkIhXaD33l6CtI2H6RmlcHaQfXsVpvwCSqmPZ7mj0
xiBgVrEM4HDohwU2Nelnpm+LCSZkLEPV9a7B35PcEOIxOOo7GnNSbu8xYqPIpL3W/Lrwhdi5Irqu
ftBIu1qbW9khISOC4QqQv3TqGhCOJhTzJiBjBCMNRrvpXZjOM13wFDAOo+hoGFJP5z8uPKSAOp4I
e5OZGXT7ARfLFFulMOmWmd9Ko0G+gc/r6np/gae1CCuGBo0dCj+eMzwkOJ68Phut7KF0kGNw4doT
Hmh8z2HmF0fLz9O9VWwxSyR+MglIX3m7IzTQImjyxaDdLWuLxZy9BKw+rBYfKc0cTjJgUPXqwPgQ
v/+zPFBIRDaMHkplfki/lsyoxrNub9vgOrgUb6XLdRDmQcopKZCUP/dNFKgm4ebiocnGEX/oc1Is
nGkuipAjrbIZDfQvNmZ/uN21wtZj2CVYBQL4AYASF4O57bPzZt5IVhx53EHrE7FiovqJA9TtFm68
K5tobWSz/rb6GGAMsuBfvNfrgOlsmJO28E/UJDV+VrNvFiezG64fklIOQcwCPNKSRCkD6lC1dvPL
2FA8JfRLoQcLX2fkgBEZ7DLGsW4KaH2mtJKMQ1AMVOKw3HJlYW8TQVAPZ9uM679WaytuYr0QnhTb
J2AtZLYhvRRsIsaQLNkke7hfwaEw5UWoseVUIraBy84n8mGEhGnxU706QTmgU7anwYougiJtr2ao
m/gEQ+pGIz5reKtiy3WbYViZMkEKs+2i6Y4Jc+NsyAWZyi1cscZwW324iyePjwrCuFQNx5oWV1wB
BsekHn3mHz9Whdrk9z+R7N1K9gIKKSwgBZu6L7D8hdVh8oDnubCfnKBPGNBrwGRMM9KYRlsGIsWD
qgcQhibB7mDIBYoaulyQ7uSj/vRKxxFnfDjsYkniQ9bxk9vlstssfnpfQFKkvZWaiVAHK54YLnrW
FkUneP3x1IDVuoJyMJx+Vl1iKChNpXl2NACzaaNvx+ODN806ed+qGThBYkCOZTwjQXS6IgyGZRhF
dZNq3gkxIAVlpRl3gjSVd24Q1g5eXom1SVUeRiKCjQGpxfn4cWhORRn2z9AaN1Yut7A3slXdgAFe
cNrjlWSjT8IeS7RMj9jIpdRAhqGHB9CM+7vYcF0mAjxdIQbOvZ/Qpdop8nnlOxF5NDUwY1blynRX
OYCkXacP50crgQNyQGWgTQHSHYFPIXxWrDZ3tMDYuiP4hSuSmrgQLWPkshS2KUehPXGzLyL+ifbj
zG9IvNx+ZkxY831ft4Skvi0EeRMigQC+6A63I+xDs8oMHEIL/63R/fG2x+CvLaVQ5xTwLd91yJSg
9sORomhvzo2Bq7ykA4RtmXyoFzA2zoNXfzcU8YFeX6ByEr3qf+e9XQgmx0tfaxmUxia4cBOqwTCJ
b3VnZbHUuRPBl5+xdaY3D9Dt0U4a7qnZlA0l1OLHzU+gg1tDdROMjpvZKShj/j2fFQF1gmmyQyf6
h2Xd1Sw0JLNReKcbDqKu+i+WhUm898RPeQo2mUY9tm1VMi/2R2H//0/KA3C9FD7nhU/NLLFU4YEl
kARyyU5EEgN+f2RAnWSHhQzVGpgYvxeReweYTbYGMfPWGc4Cy0SfCYE7MyY4e7I+Nkql164mU+b+
JOXIgxaMI56xHHJStyCfKSlCovNZCxWluzKVAwExseOJnG55ybPW+D2A3usvqQ7LThBUaa5ZUNDz
HYAbZb445LlmMx+jgSz1OmaS2EWqaSBRXlYe9JNuvIJfTho1TGUWI0bxqhe74t7PG6SJTXPVa7jg
bb1+1+hw6FPUtvSQQktbE1+ZbdsFnO5DqjrrtdZYKzmwo1BhD9zrrxSdEJYChn025FFgroNwVIQq
yj96p75XC+Rd6UCtc8pvgnWk9qnTuZj6pMQ4rR7O8L0dQkannZ0Yb1+4WpAHpH6J2OXNnlrrGglB
ojbeda3rm/aAfxq4kwCK0nO9lUZFDMd03nIe0R907IVsFrLQFZ4ChA7+BDmVlXC3ehJ9+REUUNtt
xfpaNCSWGlp5adTXcWJzC1hoOD4gwged4DBvU9ekAnlw4gk40EvptZcGxqD931gifz3L70ThI1rI
o/9946U5s3JmyfFyCYRWjdxd9cV6xq+6Hmva6kB71v9jsXjcUiHzkx4u/4ww+iuB9h+TSiFeRlAw
o4AEkeEGmuRFsatPnhoWAAxLWtUM0J0ReENCNv+00AF7PJT7k4/yrOS0pooGik9Snc7H0vkfIft9
mL8d/4JC7zIVdDzBXLXvQ7GQdurrosiDxq+tpFKd87pcKphqG3gwF8Y/eFW2xOBnX1MjDye7YQUJ
E0vzIpDnV6xuj3P7eJpsl0VxcuP0edlV5uu/vKUbeKt/34HY+k3KToPgNc4RbieKfeMhLWOJ6xyv
oIc+iHwQIDKEUooQWLb5qzCl1+7CqlCc4go8yiP4OhRLln4qEZ1zrd4ETgI2E0XHw8k9SlMXF2ZS
7dAdJK/h6SAvJIy8r64qwqTIGrrjjgPd3Moz4sQSXPw4UVlmPk1gJSBUAqmpr6duLDabwZjKJgov
zLtE90peX2Vn/TgGEe6T6cw3AW3k7LVh1I4cyTHgrZX9oUxqdqt01ix1g+X6oYf+BGiBGH7EMopY
nyFYCkU9xnc/5OTeR69ZjV+f4hf2n9u4nlPQRdPSsqQBgSfkTPBYRsyvNH+9bBiSQwAUSjwg9CHM
6RTcfL2JrIai/bG59bVsEzgnahpj1iQOdoyWIRH5xr077bIM2UYFXJQ0jtqLlao5VqYxiC6LDbXe
crlS96zSRzwGBv6kCwXMzGmWq2ISg0TvWy6lr1XXyvHDi0uGbxTRfwqAkxIM4XiCuQbreNePCyvB
/ZMkxWOnZThHUjVGis1L40rbnbJN12sCsV6lxz8qVzkzXbQpMJiJv+uyS0uSLrs15tcxJQFYsf+3
Xk0PRkk5LjDkoRSsJmGWHgsGRPsaubupkDsJm27QrRoAblMLDb1ujGbJ+g8lJSmKddSmcBadpeiB
NMPr5VOmLY5nX4gY3/d15J+6yeXXE0iH5r99zpVCLlZ5eoNe3MHQ9nNoVtqF5rnTY7yBM462scHx
XgHQCXoX9IHgK9SZakFmjzHWt2lVIZesaZoDwAUqX46s8EMH309WJ58JzYOe7ZMXlZY8J92HwFFG
hwEazGq50K2Gow8JBg1a0vHuRDP7xedTOp17v/CaKQ8uezBQYUb1GgxbiOyZO53ALac1BZPbOfNF
3l6hWljVasSULXZ7mk6wTZhnZbb4a7yyMKdEbjU+iIRPVBC70iGWL265uhhn8sIi6NOt45rGq396
maXzoCH6JeWaT7Sypz3De/1NT8MKatEsdzA2lt1RJS2SG4ZR2nhoOZyLQs/LYlp39C1H8DNFo96d
AIIxHic2PhlpdSlFpKXB6hEPsB9oQxiddnIZ/Ho0atbmRZCxutj4NwzeIPQNrwlDYcELUeaZG0sD
yVwjTOGbuPnx0vQzUDXC144ldsZSFzI5x3xlH8RHh9RA2J9+9Ab3dkl48kO5ssh0NU5Ac4GESuYs
yKsbXvCtvj0O+sZ/g/xWlFjmQzq0ZvYyo81BfoZGdrsJjU1NRgvD1JWjIM63+Wjnk5hWRkBgVrs/
WNZI9ByFy3lXr3rmLvuDUovKbC8P9kQkTUmZF7Fu+GRQuMJEgRd+2xacaTuEm5PIhfbZ8vCa76uE
MOCjBP3N5gdOTBB3QNnU1GBmK6yh23Pan6VY4MuVWCnwpI3n9rWmws/IgQqw/mvBz5VGSTP3/vm4
/3FATV+uyO1+r/sw7mcy2DbrM4XKKxcTIo6KCaXozOdFEl0oP1r8UJSNSsDb08xXbLQ0OULA6sV1
fCvCl9xFJy0WYkKYZI492Z8cEFDODAJx0Xj3LnlPGVwhPR+u4wm4s7rkRuDZlGVnJ56oeyZiuHxD
iArLdqEktFttKM4oIEe5Zp4JAQkb/HqmlEOU8WYxULOf7IezHNHZgAl2dMNgPyN3oRuikwM5DdCx
NJwUs0icnvJ+TnuCGnwAJVSJ+/zj+/7YQna9I8GaY2gl3mJlCJOxj0Z1YwqdzgxJMOHpRTqQgaDb
mn21QdmbRPPPMUDasqr5f1yMvQ5lwSw3kbEg4T2h1K8WMBHxNAmLCZ27JveM4vD5P03X6U6bpmor
Q0IzMYAAOSy588J9D8qoxsL6rGQvG+LCKprKQMOhazRgkBoS0MiB0SZcjxVqVwIED+tG6NriY5G3
OgTpWsBpQdFNIMVt9FSRjVdTsOXIAmQoIjPrm/ksu5Iz+lex8Sf7tXeRmUtxdDLic8mmjAVEItS6
l7jA2kepV5FWXgWTEz/hgTIC+2CpGDnIWtH0DdrtakroXRFVKOAGjRHZjiqOCVLrD0iwxWUtGKi5
mC5r50qRnXqY4scDn+N4/oGKJ81enSGJ4bKgVnwc9DKhqreC7EUlHOf/YTN2M2ouiW8Kok7vVJGI
Hg+iA3khEWD3HFhVP9qO+7mPdFeZ0RxwC4WCSuFIYt+mDZ3CM0wzPN5nF3niE2MzuMIQxolQXREV
X7fryoJmExJcm2BeokA3fwLVmoh7GZcgcz4YD4KlZCE/BbTYFg+NWTPWY6w7McUi6X4xZzfgfIDz
5AD0xU3scwOvvaXQ8WjKfcoaT2a3hMvWTKq57Cr+ZBcE+jt6r2gtwpKtnqyKb61FzNeTVuV7MX2S
mR59IXvTNcu4opCMLawyYrLWVGm4JVDsUooB1EOIXv4Ib/tRD/tymhGuWJYF14MNP0/8NvEOt7/4
3oaZnJNaaAFB5FM9/VCauMTULyY/5xk4qxtPuC85jfEI7bB4NBWdVI4+74qDgc/zBGzE9yWDH92M
dqea5WMGUlaxXmCL93xPFiQusNHmuPYVt9tE/eK1huoA40viimKTI/bHqh+gi0jfvYYtxdwtibUy
MwVK/YOM36g5oEh8E51wsk3oJs2TIWblwc32EkD0dPTtRcbMpgC7Vw8xTgBl3FqiNYtoeAp6gKOR
IJwlQN0D4wgPvgvWi4/Ii5Mgcc5RWD93R8GZVKHitTyzn1AaHR5LjCb1cfmj1Wm8m3MUmoIqLVmF
B5WM+q/Ovl3XglVGdl9Uay0+qDDgGeOOJyQIUi7itGmpyYF5PGhB42ZyE3IRin86h5mxH/9GxWbV
+PXzL45yAd2T/wpTK20kvA3ppfVQs563o5XgrpCkN0LM4NWPDXBMWwl13M0ZGTcOi5CTi/kNQXV0
3VoH65G/y35EgPpZ8Zti8TRO43z9jrZf1OLrldI2IWFuYMHDK8g1D1fk+d9ypSQTdxfOdKDcSzC4
aSn4e5flanGhXC3KLD2hbrWJYRMChjy2QURdopU1E55l7D/lQUU1GiGy8hN6kKKyngxUcJKZmTfZ
PVsW+uDER7S55PWgzpVl2YqKy2b805Qd3m4dv2m2waWs06afrIkGj+F1YIeWBE8z+Q83x1bjxpl4
yC3fIfVHRi+myhASo2jjqGe8pBcbMpZlxle7QF3VdiQGPLvgCdloBkMGTB3OlVbThL0QsnmHO2WF
BpW/9w2SUUwnFjfVAS7tE3xtfl3JZ3plo/cY0JhQHf6MM5FsQncCT2f+VyELqshPq5hRzVS9t4hQ
dwCiDZG52wqzRx63Qj43F5rdNjUN0mEccHKB9iJUTiGL8i4bkG3F8tS2sBH05eaoMEta8bkaH+Ed
nNEOT+SM63tTdjJ2U3VDWd6IadtBbqaKbPo6BGdg9PnRkES+3RCC78uSvt9Qp7kdVJfBbKDbPYSb
aytdfRi1itY/kGlSw/hyIsdCmlOl5n+eZaO6yRGS7dfN71NuopAS3XroRdmtOMPML733aRNW0CV1
eEC9tgq+D3RPjH2xXjfV9B6XDrYLVCVW/BX6z+0+WdkIimN0hQ0eZQCcK3vZvfWdGfXJ1QmYVSR7
cqES1yWjMSF9Bc8mB0lS0OkriTNBY0y5DuuZirvsOOFyFuCbD3f4iZR6s4odqLmQJAuWVIDiahq0
a05IVri8h3iDit4GfvVFnqHHqrNLQr6dn5rloWkcq88Zz1jGO2MFRBGuIoCZQL7fFwkqybC75K4/
4saJ+FbCfwZ+wQIHB2k2Q9sLG3iEQPKy6riBK80yXk6wEmZQgaI0x6msFO6zigDKv13GxfAcnY9/
nV7bAx/STbUBi5qbjaBxPKyPyboQISe6jPTki1W/A9ky9shB52bUlU7QeTXoMlHGfrx6rYmP2QA1
S4kF4DBtlG4mrdriMIwxxfdKEnvNsAFrJkO4L4KgzrrVjWeatVBckrcOKolCjZ3P/qjoBwyZDeZy
SATGqUKVZKW3EMgdSTmsfvg4iD1XdC7XQ6p5Mjt4UQf4sHJcb67VsWbwiPF3AmouXqAK6T3TFEp9
KBQIm6HLdBn234D4Ehe+wxUzCUQuqfvIc3JerxHqWI/FcPihQ9Ls8kKYYGHDsNra2AbUO3QIq8FY
6gwUCeLy5imoGh+eTeXtrI+jVZnlac7vWpMhWP25Ev9l6V/LYgB/myvbVxoviXCt84/JvAZzIDAj
As2C4pgP4NvVUIK+j2yvJrSXy5QouEkCff9m/E6FWa8+NpfSx3SnV5t0ocYCYNTuELZwVZ4XQjfk
BAFC3vFK2woHXyJq0N7k+O8dqEzu0DBDZ69mBjO/fgofNMxrqtyqTr+LR+bIYFFC009a+UDs2MJX
dnoq3988JfRwZAtoYU32c8wh5VVyJcWFF6cV69pQmGQOLODFxp2k0yamC4mcRwEjXnD6fKjKDgke
YDlSHGR12uBD81tcZEqhLjX6LsQPn7J31HQiEME3TCvS67Rm5y0fqfeod5FkjQa9Fy6SOGAAiOfo
XdJsd/7z31CczUoTdNVZYhx/RE3dkoZ0kHb6Wk/H11fbrs9a28XbF7yw2PX1+/i9mA5T5O4+T5RD
+msKyTyixELFWiYuEqLvGOrVsC6AFuabyS5ySwdhxnq8YS9n59GL3dQd63ktrsbzn4eEb236XoJq
1kuw5yFknkuU2Z/VqJNRmy2WsLSx6q57OCgECK5nCHaTPDB1MfbdqfQcELIvUvqm0cF/ci3RemOR
38MTcpa1zTADf9y1dfVPV91pjQHpOcG1F1C0zx0rhTfwUf/mYEJieTM/9MkYth1ubl6z3XeKJRk9
ELNsRM/ea0EJSksYg3h9NJHDGf91E4VNQbx8GzC4/FD5G6QeB5LymUiHm/6mTpvp9nuvimsIIDxW
zTv7sMf12OWphwu0kjRNGcti7oEeULr6+BjDNIFXVSp9kZqw5HGh1V46gUjqcXhS+YdVVLXJIxxm
v6Z7taYgyMj9/07mpRNEXQpaTlagFsIIkSu8dwvRqROFLY6pXCzRhi2i7/7aWsLlJHFuWlY5Bsar
wNSFdl2W8XZk5mH8EGBMIYc3Is2RCho+rMoXOJlVyXrCXgT4hkivyE0IbVQWmc3a02lf66wFl16Q
0VlHUEZacPVIbSJHMAD4VkQZFmu88kKbbs/SyP6JEJYLpz8W+AAGwnrGSrjq1+7bHVRx/d5wgacp
+6OPhnVAVOoniCPTwcE/ahxmGp6hQ/RN4kZyrLaJAaTlWorP8Zr0cwMs09SDIqEagrp7Qoyobs0M
Pl3DEjjWwyPliq4oyZP6wMoEKNMIMf0cwmRaIZ6CfvXMwdOf9Y7ba2ClbJDw/+GMO8ZDnYifxKes
7KSOSNm6SYOELKZYPIyagUruUfQBNlf+G6QOPryPVl6E3KuiF/a6wQ4U9OwzUoNfvoFPPMimAtYZ
ZzVobsO55cLawruUI/4IxK3YVA/q/BXaY4L39yiQh/C+eDXr8oorQPabx2ZjHF3PI/njOXdLK+CB
DVWmCX+x5GZB3ER6npdwlzUB/0aanRE+29BaVwbMo8AoAVPJ2RFuFwndcgY2E55/0n3dCCaSmcaH
eaxFaHnQv6o1K9bqpNO4sx+EwHqrDVkm/BQMpktYvIDe1enknLrAb/3UzsNu4VL8JmJtHTq/FEaK
5ykRbWC1ohVVxEa4p5eSZUcAagLEJj7JAdm1aC4KhqeYfiRRdYu8NnJE2WD3jc66TEDuo2C880NC
+x/NUZokAg8BOHqwQKDOuaz78tz1GWlUBm/p9kbSL4Bdl4rgRpFGMMUJVaWUxjrwIf7OMuQYJhwe
KkuFLlor17gFdI74BMLiCRlVMz9zU+3zNUhAHzg66hVtFOYcNruVjwLXC0BOsAV2Vqkz6D0+6gNJ
2QHHLVhfggEn1RKxSceYKMGjkDVgx8EQ8Tov2jvT2MAF6YYsXuSUqhaE2S64pz4EVs3D3aT13PPb
uD+weyMY2Uq5zgjS0b3YvryFUJyO58AeDrZ6pfEZ+O1iu21begY7sHOqPpp7SxnsY2Bb4c6iUErR
IrLO1bGJzsTN3JS6yrYnVF/dU3A+McAIzzmN6BiRmrtlHvOeNdthnbposQbrGTai9/rtayYwC10+
JcTkMJI8eUqhIX683DELu6wTITg4RwygPw40OeASoWLOZh1aghSQCecv+u7w/146yyI3UzLQFgfZ
KoEapZJyai9fMFYFNxdhdD563iQf2oe4T5mTgL3w+ZxwoUcw/LL4bTY4T2h6E/+YvjMIIv9Wl8d+
VnrVzf/u9Gm/nlt2SPNYxECHIG6aLnghRWnsYlt7BfC/7uFySdytWZ5QFtb6xyoxF+1eVO3ANF1F
Nk4Z5fR25Zqxr5amA+7+HEl94cATiPAKJk6hziLwnKrQP0lOFsxC4EoMulje1FxNQgschRp5PMj7
xneiAnB3k6A6a82u5YU+sDEUwyy/4rUCF6N4wicWUibb9XxtAlM5MKoUmefCyepCTIzjWF+yRS2e
WVHiroqsDLKPJ2XKm40jb1bonmEIPaQ6D47ONPiRdI2Cu9EsFxomPlY9OklcxJgNxHbamp8qUqcs
E+p2d7l+EDlM/jw9lqMvLSGgONZfjFEmhOkMNU8fltqhrkSF8G/tWfFEWaMBNGzCKgyPzbjrYqO5
qCULxn5J6hVMy8/rfj31nnZM+TpTmU4fn4I6Sca3J+bmgEKjaPREpLBe437L3CVd6MBJznyqs5AW
z03tPhmsn1JotBBMOMBywjkQF0+0m7s7nQx5awoOQ36C0Bobeyd2AxVTfS8RBNkRIt4qTzfrv5VW
Gea9UD7tkHQ7Ld9BWHJAiV3AyFf55ekBPIt2AcWYpB7Y6llyXpfA2zXrVIGPYiM3JOenAUJZjjyP
YZLDoWyXeX1Yac4BJA77luQH0V4UflIddxQqV/vzn7dbxSu9ZmdlCfXYtaBaMlUPYM9Y3IwTHjhE
7FxkglCk8qm5TJ7c0W+EF7JZGnb0fQ5FgXHTnkQZXN35NiNaANTwWVBOlDidwfdGql7smCHPA0ji
vMWAES0qoIQLSWlgXhwyCNumwp05UmxJJOnB5wRNUVBjuc0kghPvOcPGO0r3M09NW100w7mp9uWa
paH6DR/1xybLvv+5MJxaEKBPD4LxIYTCs6UPXVs795+xXTPFNZMAIem6nwevGD/ynNbvZz9nYlLv
b2KitaNMScMbNdC0QjjoapRmYmpLK26MpyzoerxDgAdpY8MenWEC+8vf3LvkogOsNhakr5lNrnU3
0fs2QrvdTxKARNIdBhInlu9Cs5Cv6h0XJYR6xl3xAKY9TXXM6yxRadfgyC03jPV5bLFAG5O0AB7a
NlbqJSgg6KV+Sv/9sqwKgWORmHxA1AevbFUY98ZbRGSUU1XNooO7+ey/luOqTvC47U8XyzUQ8da2
pnuf8rNzuBHV/h2hbb/kZkIh8nXwy+v2aOK+fjDQo08/AeRGH5m4k9KfBParNR/kO3osxe0BZZSO
SEAjjPJhTfKu+LCFqA2oyWWSbd7aEu19ffcs4nqo45LPL1x4BuHlbRPqh9U4qCdovsamqPdv13Ul
WNyGtMHjwCvBN+05VsMcbkgru3YRirCvpwR7XxS/NjDBJR+XQ1GtrSLs1HaKIbp8/ndE/cQ9GHkL
l/dBeuvxC6gyIinHQkFaJlQntjYLoj/B35EXV8qQxJKV0X6kDVC3EkwfJ9lSZP3/LUUZ8haWP2X1
NoNzGNPN9bHPdglmPMDGrzrQ4pvuV9/awenms/KV6QZ3Hrjs+MBP1KVlFm3RaaMWVC+0X6kZItEL
G/ZcW+/t5/Pg40tMq3xte0aFGFltyZLQ7PGX0vOR4ILtZMAq0w5n99JUE9UwwiVMm5xdgTuj3k8k
0583F5UnBW0a9a2hsrKc7nr3CoULqV+5x/ElDNYSDVvsxO9mMrCVQrnb0v3XMIgB3F2XEyBpPUMj
OLwDXeDfAZyusQT7GxCJRW77wPmolkg/dVfwEdwN+aQO5B51/THfYhW/Vx2YDZ8llOpK81CPOcgO
CtJ5nIqLMr/VZxY3AueQJ/InI+jZ159VNGfp+tFuziJQiuzOXcQS1izCoUH0amAu9h6lzDULFkb0
yqh716hSunjDWR1SQGktliTtLn3f1RtUmWuBdL/9r1p6S/Db8QHBT4kVZmaNChsmyJ7pSAT7j1B5
T52RPCM3rtdFT24sQPrCAFvgMYh2OUxB7v4up/Ym0D8TezYjxgybIKm6++pAK4bCZSxECqtKkpb/
FEjXar4fVq0KuhfASzb6nTdMGryp4RrKhXgU6Dqc+BLo5w3V9RmBHHUJEY1y6i08rLcjZtLyJoiA
WlOkvEYln4MTSuRM/xwzQb3IAwXnGci3EnSpKlZRQQS6HfiVON2VfcVi+tILhIt+nwoMKEDzw+rN
K5TO3gQQmz9VW/HnluilXB29cWULyjahR0UCqaEMgNgyyIqqyQC4XD5cn6uMsz5Xhi5sBWCx1TtW
fiUky67Sgzg8klQ/bvC602YrvAI7ag9T+ZwPgqJuIgx706I5gLx9dfRJlRqAdKAduAigIhgCkrK7
UvlXi4/UEL8/WQvCFyyhlTT3YyCReDBU9HZhk3hDK0rHgW9/NM1jZLJCrdBor+TJ44HHFQdJ6s0W
lt9bZoY593hHuq3U4kX4RgtHmsGml0hwrvIS09/XJnSwgaFBY06X+Xui9fq3L153vKomtDqVAZTA
nLj9X2jhvQvgLMV/T3mfuIaSDDSTl8OjlDWkSaHrbcgYwKnLHmFPEFMrAvDcgyt1RvOrlmKBc7B0
AeeJBUGFwLxcJwhZ8QaOIs5Ra1uJVmalA4Lt6er2pSULPBo06IpcbdiVZXbqOPtHZYycPrPivjGK
gYr7DBhnitFOUxyrdWqJR+Mx5Wgo9Ir59wCmK2TTGwCfym4nCAjCOg5Olth3MG+J0kvFPaY0Qlbd
vzrYuMO8tXPwus29AzXWuHxa4Zb3KsbeROnWFzts9BU3iTBt5SxHFiGjPzqFcFcLO0xF7y2dmyTZ
ctONvMxrQoOs/TrP9kBJyqBiF3RuV8VxkDhcq0VfygIH2lPL/goGhK+4hbdvLglbqbNK9H+Gs4n2
KxW2TCxHbPq/773XpD6v78SsL8rClvf8Ccirw6vr9kUgzHdUaVDctyiZXPN0WT8zTcNDI5NTpQx3
LJT3eYMRmldO6523NbSQa/oRWy49Zx4eH5VoI5GAHp74Hy7jHm3GRyL+ZXJONQn0D/HGDdhcJLEJ
yWON69kvAVKf4V9mvYGGh+ehhiPLQJj0fJ+PybePPXPm/xq2GhYZGYl86desok51up4UBACu8Sel
ECe0iJMPo7hmfD0QBIhbZhB3aMBzZneeMDiRpdsub/avcR2Y5Atdh7WMplrLc+12zA5EqeC/EUIQ
KnuQJ4hZX1Q6cvkqLh4Yx8w/XmgZh5UAdtNcd430H3lm8VAQVDoPP7jVG5Yia/x86QUm0+XpAKDS
08sfjdjcUtmVu0wRNgpUzsSvyr+A9rmLPQYcqp11QckdY/UBi34Oc+B9voe6VcHLwpQlUA+tPDyU
rUV/vSK3nIlSPSq/1ckJ/l3FYjKJJPZX+qDy+2HMyOUWIvoGgbZ4wFCA6bWzgWx+4p9Ci6i2/CV3
Y+N31hs2O1cTdh8giXBi4FDCF64GciR1v98qIC1e4SUCIe4kmRmqBpfBtFOOg9hDqxNx48SxdvgV
wNUloP936yV7sCXcVC7nDryqBoG+OzA5U2cPV3ymNpM+h1GlKY6OW/XnBZ7posOKOpcQC0o6KhX0
RBhQc5pTuqmaicaqcx+WhrfDvjzM7hKdpd9FCieYILaKc1AXUSmKTdMYLFAJu1zg10ItTgSQWN77
nW26k0Uka3BqGnDrIx1m0xEQGY/ShKlOaC9+eXn2jGw0u1yr5VcW8n+kGTnFUkyuOy0LC8FH0Ugi
V6e3D0fGhQ6Hb+a/dUqjO8dE9AsW1SBxdGAfq4dogxnK+kav5KomvCMXH9KpYRbhLsIcu7PEDvXM
hhI5i0NTBijXbMlxupq2WDapCW3l71W8oflZXtAEg5IpYrC9YkBM8txYJ9ClM1uCetGoF62odwLS
cWaEFE9xpC16P796/JFZJKaxXbtBM7HsFJEky+nQng6IP2CYW8V13aDNLBpCHMnah1K+4f7YHZ4h
T0j+DNBWJiAdpCnmKUYwJQTBNE5UHNNLOjE0g44qjmKUKw2llIaeCZfX/sDsCA+EvnCVdqeOA2p5
aj9Wm5oQzAQ0uqX+17OttMeoK/eIM5m28HZmUTJArpmlyIEi9sJpx6g00dKgbZhOZ0lEp1u/Ip6Q
85tIStUq7Rtw7vj7hAzPoVQyMkOQIoP9FPxMP3Fer8x4NdNLX0Kz2KwC9TlWGQEjbno6/COL7X2L
KsvBrsbqdaKWRw8Ru1yPG7qcg0J+qeve55cYOtzRZXtKogtHpAv0abrL+vA9mJbOJ8HevT3fvvGI
SwSo5rfnQM71BK6Lmxw08Kaid8bCrFdd/NmUY+AhadGzRuidtof0vlQ6x/G0onL8x+u7ZDz/LVcV
QApRgphzJRL+odfexQkEBIKc7dIxOH9LFeksZNZ/PJrpGIwPBlzA0YwiX5E4n/AIarZsKpZkcQyA
F7/75LtX5c2/OIhFXDYtw17FuIgGBSHYm9DoMRDZQttYMElAIgWirJajiECitDFApw8YYRclIvos
2OMfbqOHVKmO0hudD2EAnEykFFt/+gZkhKkPugswaUVJi/7hz3Br71/NsTIgWySs1BMkd/Ds+ROJ
37rsuqrYlfaGVXObTVwG1sz+yjNZ7dpsxxAXHkAQHaD1LZspryt3Q6aoZQ/UHHg1GDrwYw2ouLOF
/bfLGoMf1UTdbBh1HY9wip6Ui94AC2uYFiu8FnF/Ml2hBc8hD0vT2+0TudZXy8qtttmBmvTECXUk
OmlX9FsA/5IHtNk2eER3GK8HqwTFbe0NzvfAMiq5msd772Gh9vfpGyadD2HrZDCNsvSyns+g2uss
gDcyC/XnO4OVSs6AMTnrkzX6UlDeWKpqSU/MP/6/vKy5inr8JQUvfco1xmdhv3EUAcnUCYXKmoOk
KvBW65RhqkSNZYaZprJeLGtbxmvcbYuXjFj+atwZQmrBIiWIS/j1+Qzu4cwagBniRAU1sU8HrAUC
wGnmCL7xeqzuoLc85CjIuO/pNBBlgaM6q2o5b7LA7IEesh+mtS1fZrZ0tbADr4A3LvbXoSSeZM0L
bh/91ueLxIiIS4CJ10FadarnUJQDbzHQCHMbRmqwoP0gJ+liAe36plMy7OJIefoCiFMN538BIEXo
ToKTfKT0EfEmWfumSqSqUkgo5SvTxPosLd+Qfks0gwQ7j1p54tQ/FWaDSSAJv5azozbHpLA3nwhL
MWct/1oV+GvpTL4PCkq4jLVp3i60rR1oGvJHsGOOgu7y0aiX2mdzfzS7dBkGJXqCaEhVVVUPYJt+
oSpCFoC1LIcoAVInRfNYEQmcX682I0NYdV7Q7iEQeoqnDZlu5Sd58xd+f2oVBLNtzY4P7c8Gu5Bh
2P4mVOuWN4E3jkHzdIL0YMGk6Ff1AYwCkeLLvPAu1cV71wFSUWdA0X2FOuYhPVrfLWkbSJ7akaF8
iS0mOXuXxfMDAjOg41Yjh9hGevn+AeQGtrnn8S6z+J2XwZbR8k/ZaoJf4bj8nSPjdYXVg/VdR0kj
mTkxNHJhyMnLLu79QqYSvaKaZ4iP6qa1kn3GJy/7NDDgFAi1CAmhs6EF/t2siascBmwxpvXbC8C4
I6A7UD9s6YphvNKZzOk4DHq3lORopORK3iD7ssLGp7tdMBVxneg3J1sjwixRdyB169+x1/py7B+/
xQ8qtvxU7DB/QgUIYzV/ZDruXarZGNdx1BDhk7b2lSLr8i1qDBIFlsfhPRX06xBkWdOlPYqVMuz3
bnbkDWrz4huyx7YuK4Oa1f4TXLxMux+FahltzPVMSEMYbknc6B6qvE+btvtufdTluxt0uwc/VJl2
qa9EuRTI8So2QW7y6aD9K6tuNKhRd7nuYWfLkvorF+kNc5vRuElsOgiA4Z3yS2Nv1s02gdSRrI+c
jyU88kTT4TREsgcjUnhSJ7SP9isD8boS+yRviLdakMIHhCFwmp7TuHfQs3BSEsd2gWeJ5g/KyQcr
6ULtxH7SOcW6I5cTZtnSDYvWOS53d1PhZPMdFMBRs4a9BPi6t48J6/URRfhJx8j0x240xXU3rzPi
+2LJxcLm+ORnOOx5PXVaBGUgMrzVgjcn9OXipm/aMVNTdvp1XLWcVZXh07+AQ79mN6FGSMI0gKXq
JvCZ0ymAwBGaIYtgFilgkGuuYBXW35cgy2EQiLdcOJJKspm4kotlyN/eWrV4ENLXU3oPmXfIaxWO
ACOzq7CjpOIlq9XYECQlV/kTv5LjYy/2kAgImlYurZsMa8/8ZUaGYZ7uJKBTpOKwMu5bfO3vQeaX
kkcoRFSF2qPVh4eFTmsKgRIVp0TDR9S85VoWgQMLK1Pc4oyFTAFzXW/HZ0aZtWJamR0IsFTRr25D
CJNj1p3lbUml8Ji2dHk0bYF9dkkWTbXOs89q9i0qBH/U/JVTakp9p7hc0a4rJlqfZ8ZIUQWQudFV
VBCmJ6cGBrkqLog8CQN7PtSWymHdpM0LosylD+05vvf1oldHv5I9/CpZXyD+HxUwKZcHm6+7MSuJ
Ggld+55C5175s47vH6om+VMCFbv7CUtboSvEZt8OK2D8qZq4Z8qWoU+kBC+RbjE42wHsSRJaNKq0
ieKsh0I+nlRWekmXz1D2s4OOkjJvy8rtFcxuwy7A4vH+zo8oCx7wfdvU/z1nQrWyFyjhBEp0gney
CDMwMbbNdgrHBoNWt8a7CwblaJgJBaVRNjzpbzfoKSThWrOwDtwx+eUUBfkHxrRdBUPiNmoIgZAH
MPSmom13GjErIdkJuGKIlkRMSchuxoQ1OJsKlZ0bS4ZiUWYoU6RSp8z0ctfe98OCrCcLgQiLuV41
Oxc9s4labSnxV5l3O5eWj2aYJXxl7vGgWTxnw+NqlBFshSQB1dklf76tKNvwrB02+sFvrj3GBaGy
8JQY0IVSM3B6Vbm2s5rhuWQIzq6tYAgU0t0dWeY6Rj81pfuStcE+EviPiGK1HbiKboRejRUXZFmb
NSXyYbSrQK23ZQJOHBNWh8DSXo0uwTUiYZ1MpyKg5djxwES4eYC2Q8Qo6jwgINGC1lOmq7/NZI1X
rhHz55G37KuLv+CqAxG2D3EXd5cPJOtmSxYT63b//NE9VSDTVZ+uoDswueTo76lrVEsygmR+FX2b
Iy7+tkDu9hH+wTT6pv4MbzCTLAuB3psdaTjT38dnK/QVQvnPHvYVt3M3XmORpP16bQ37QZIKsR9+
oHwm8vl3ZE6tYw/LnQE4gWD7AyNvl4NMXr49o3VRfFOq8BPVuQezyxJFg3ToJ+nPyU/Y1vUl1NEp
KaqiBugPodIrpRRZUOhNDyMdNOeYTMp6iYa3PXpSmScejP3uqM1a9wU/q0p8QOKiTT/AozcPdagr
RqyyY218bL+2XujA/YnLE/SvrmCxyqVfJTlatIgqwaLoVGnWpBIfYZDfifxjkcF00H1mULtHMcbF
5yN0ev4XMfhCj1lK5/p0DmWc4zuSMPdGMhTibkQLCzS06wlqqPX4Rof/H5ZTtvnCsM8hpUbuLVJO
o71yQnaEDIEMNayZuRx+WDQ4QwEdgggWclmVCAu/CC4DT3shWCC5rA3jWMZuJEPd0jyrpBTo0fIj
XVIEjD2N9TUE/c4qiv6xgvCaSKQedA4+WKm2mOjZ5GdihZZzpzzgQ6W/NNTuJoTiOcgJXebRyR9C
blrxd7or0cHlnJ+0hJQo47/wJ8Fae0/qtWO/ZmCcGuMuBG76GkmiuCLJBMTiFMSRyHL1S5eqG+EB
EwjbjfwNv/9YORn2ENVycjXSUwlNSQafFSUVPMHq8NVc1Ls4ymtCJA25DBJaRpC9MW6YWwiLQ0FP
79UYfH8A7s5qGo7o9J3Pt2wfo+bV9duQwxkrah3TQlM8gHoDW2tGDnQqUTkf8rbWl9RWNyoZ5nlP
ATNRZi5WI20reQVjGRS6kHtx9BC2rLs4TUWxNf1N853VEpvrRZcOE+6jBdPiB32sDTCUBdQIrpMB
FILR1r/UB4jdUP1g0XkD9SC1nb1XXm9ACP9PHUmV/ViJmyv+TVLd7/OGZZDyRo/ODDsbcrENHH0u
atj745fzxRZMFNWiIw7Zk0yn9top6tePDnVdHsxvQHU7RkAptmR1OP7qKSIinuiq9khTghBnY7Ny
NR6sSIZgGlNmewfvoNz7noGQh/51M8ELIRGBBVsbfpLL4EldpqFuQ0WGe8dXMzXI+x6kru/tL9M/
s218XeSfWAqi1ogZRYcYmsSHBrqs3DPuGpqcep1nY9XGqmAV0Rf+NWz5mxZ7fkUO3m/jolRq/IUd
ijni5KkgjbDbUZLX0nrChHB2asXGownZrzr317VRxFoGJYXidheY9KkIZigWa8vlgQRROdy0kkb5
fwg9vrY943apg91q4waElbFj62d2ZpT7ZzUlV67f3/PgqLApGHeJZGZ4vLZxiGL3oTaAFZLvgaW+
clTevuD0xquP2rbOsLW3WjF4/DE5li3FYiocloDmKf4h3ItxG8IRG6yTAHsZIrQBFC94zXKvZsLe
S0TUtovK8RzXbK1dwkeiBVFhXzwbPsMXwrAH2y3OSsFGV0PpPaDp4EENQTebKEN35nix6GLrS/tu
QhUMEBA66toCSscZwg/byiIbuQkPcueB80ybBe63Gkiczj3/sWrIXXzX62X2ciYwpOK7LWnUzfQZ
eWWXzCpjkdsN/5kAGAMqnb/tnHuoep4hTTX9Erf69OA0UtIXXoBP0D3IVqQj2gl0oh9m9u7mhGC6
liTBo8VZfyWRhwysDwfo9FhHNvHPOKHQeH06XpD8+FavcH+ukU1wsII1GG1gP08p/cFIvCzCBfJM
si7uwCM+NZBS3rR3Jc6dwK5UAZLcS7JDpNxGWZPCkWCIr7E6zdLqPOYQk1rSd1Sb8HXjH9ieN0f4
qp4VzHqobY+WPKDguXlQP4EiIkZez6YH6KYnr34NPVTL4GoYeUVTcFLhQRpHpRH7PCc0XXAxjMRA
EbqacisXNt14jVaVr6O+TG4i6SQ9k3+xLHxrtIbuJbZZ5+XAdqUWO4sYF5Tu5XPLc+2krOqNGIzA
6CSIwISR1CE+G2av2+Jei9SuPFhPVCRlF/B131C6hE4jK3tw7fKAKK4Y/ULz6t/o6EJPex9i1QsT
2YIeWOt/ydjCpI0+ItHI3Qmea7erRmWxsv1TJDA5x3kcLLAdxZfDW0Bff3VkWAO/+RJYTJMysUhV
Xci6HG9Ehs8mQFxVWw1z84YXtebCzR7jHb58RQl52L0q3o3dSGYeLjidA/VYxJBUXDzevSxL8yl5
GYX17G8du2AUy9wz1ttR87sdLU9kkW5xaVzzqBnKXMZbzETvBhtjrgSiWN82+qM+fR9UrrB5lPXQ
Mm+DZhrbI/rKj7FkJncCRXRZEXZqjU12IvcFBUR9Hf5lo0pfpwO9GY5SCTcOfajSMMllWOOSNWs5
q565/Y82ENG8Oj1+RYT6a3YCV46/BjOL3EzvqAkOe1nyjFq7nM46VQ9gSHvP6i2XoapcYTzweCJy
UJlB+eWpQN+QSWVOvBtt+NNtt2Cudqf7kgDJv0H3fcw6FugkNQ8RtANp2pMoimNwtvJEVDLXr+3u
PpNSZGQkvw4w5H2OvYnuB1YGIDPmM9Kp5uV3FGlJXJiW1LYugk6TV7Zn5n0UaD8532LtdDnKotvw
nxy4VR1jY9nVfdHLRfBdRUtIHwjXY8GEPkyy1ad3/GhW7j1R7oYyDrx3Kfe/tHiLPNjgvi5cbOle
gaSFhHPsWo38pmqATcH6ucC3l9BcIk15VKuZzMEzWFnt6uUqTIQSKWGQacJXvxL2lH6i96o/cQ3h
nI0UNdmyemT6jF9UKcR8tUI6TjTFrRToyJeU6ATvnoE8Efcr2XMhPMKi3Eq/4aMpuT1/Xm5RtLjh
RmMMzThO06cOY4tJbM8TnBI7DkamZWbdFIeazBgEPqRZ6VWr2R5AneFs+yBt77x16oqstg5+bSg0
oTuX+UEqqaN/cO64Yblz2PllBeK5Nl7jeuznCrUpwugM/+lhaxOZx6tgydbH0NAtDeWsUIA+g2gy
VutUZvP8Ee4zpWl256uzMWJLzYQUf47XA5MgTpF3l36KHoAUHQ+by0vDIyzW/XX9i6Qb8YHho72O
u7d6K2kciwIygLp+rZYF/5VvsnwGMPRkgqWP6FSE5ORFcFe2/jxwBZyCc7osLyoJiPYuCN5T9oVZ
Je4aPNvzkydYdU0+qQzdyJU/81fozNXRcnRQ8Wm/LLh+HAdIPW2NpvdhFPsOwomyX6dHvScug67k
Ntbm3rgOMFzfmRnxP2FN3ZwXrvtakPiYjWueHEByJcw7DMp0hJxp+D8Mdl96dA/XohcYnPH0JZIg
TWBs847AjZQmG9+YTF+34MJDCnb0REL9HsZQ/wu7ZTHnfPWBH9W2gXUaPArNnefMxHXAx+926lMp
NI9qT4i44FDCQLA5whQYR+rixwDDl36If3OAhd9aNxDFhnFNcGkM6JrU7iwYO+S7glBkMuiZasni
ZpDzV7EqlkJh8oDwavOe5jso0C48lbQK7X/TBeq8zkc+8li+35LOy3EL5ksto06ZRBV0jrXyDZcN
+mRlh7+jO7F0ijeROUSvECUPT1CqghEIAdiaIwzmNg5m/Hg8BBHHGy6mZxafk0C2MAKxfaWogiNn
aPVrJ5HYuMbNVAsbXcrIgGQNkRTU7pf3RVY6L5pkuK2MjAbz8NcJMjpZaI99KQ31sI4NZgcubgo7
wu++PE9uTZA/W1V1kZ3LHcsbz45OB8RJ2aPSBYlsHVnwgNwh6jMrZOGCbMVr7y9s8OtW9gsw+3Fv
6hxIuVzq/MOSu4yNiyhP0Qaf88CqEGF9ysaZ3zSndD/aofEgjvuv3C95XP4B1FEwdH7qrQyzfxN1
9eKd1TRGLW9QqNzjFoQ3Mx91cy9/UuYxQ2uhuOtyeEs2IUKgEMFeGgWx+iq5sn4LGMSMkZls4JOv
3t68EoT+0hp5ik7Va8ruWrp0NQdelY+wAlPFsxS0/gs9MNauomFuh/6twoqV3pnWL41ioMax4483
42RqmB9ohM5qjSdp8rt26kcwyjyee+7s+AWipGi8OxCuIMv+4V9fE37vApCfWPpzmonDuttPuV5g
yY60dtt052sB8AKCGgI1KSUWcg46F0uLSb3PlbBq8mkQE3V5rigNsRiAs5j/9KIVQThdFs5wCcz7
Kb+NO0yzj1oX0VQltXOe/HY71Ziahq33m896FgcXkzYr7xxBBJUwSMswtMnB4m5V5NDJ+5GZqVD9
in7SnWgMQXfKv+HcgdwFKFqJxwAtf9OF7o2n7HTvG90HaReTGfIRU5Q0MOBlN0cOnhiPLY8mlo8o
TPcONzrEoQkRCBR2+WzAjV/KlVsCaXQH5DQly7154MrLWzzdR0oVGdrMM9Qhf+VuZYpjkyQgrOjH
lWRFf+PbSVWOYfqxPCOKUbLKxr1Vc0WqiQ1kz7KoDDanoyiJC5M8Gb2ad6lLfCDYKUTE/VV8lOMR
EMn58X2is00BDpIF7oDb/VXz/c0KnHFUBKpkE4MYpUWBXJNcE+O4z8dA1cConCud1Fe2J85l+33M
30yc0r9tVTvt/CmzvXhiOgE1BUXy/rDk7S9IxQEDnowbt8oYedPW0X+gMhdUa1SsiAvCsQ8Bx5xv
xTIXz/WFITrLf37/iwOVOtUJP3QywuRT9PMR1skBgpMNpPh0DA1qaEpkj6xZd0qvg4D+8dZtAh2E
58H0pAtuY1PcWjq/zmiyVYnfidSoa4mCcpZcHAgAcsFtyoi8WjmdIzeWsfd95VGsg4KHcKsv6qv9
A+HosQa7XYVdiof/fN0x7bkB+nkQW3tVF8MmAsi9WKVtJ0lnjKR5vfm/dPPC6o47wZHlSEX9gzEa
2avbSSb+3XEqywnbyMVZzDMr7fDO/hx/+/mw9iivSF0uPncFv4CY62sKZ50MWQQbFOF/BmnubsJD
b1SKLWselwzmtJYwFw8mLdlPlXTvPF1TEJsSzLyezsVU66MxSqri/ZmihwxdZRubSxETKbXFVWUe
qDNdycGVeV4GqGBPIfR+1CL28atwWIGWSY0m9TWYGXBq9o33q5zl67qZn7fmMn4g185FjidfIcPA
pSC3YC2STWvddCf8YRxfUfbVGwg1qPsAZLrcA35Ed2jjPYj98ax608L/kA71RPwhKhuLYADeGpMt
BTK3gN5y5jcVL1cPiV21SwTX5VNkbwObTtQkN8leM1t4Q2FI9heEWB9wbYIEPpW0/01CpUPQqMHs
0d2FIeVIkaESdJKwgLHMAUOWffWKAcU7GA0kyWOtnIkI3xnN07pgp5azm6Xv6/HCoLwLhngzbK/A
Imk0DhY8eIDuFIhH8yewukeuT2kntP7Xv/ThoZ5j4vEu14TS3xze5y7RjhUPhaT0rzZ32dD+uHRA
S+madhI6TxdPlMJ+CFA5GaShwwK6+qzB7hNB+f4A636q+mbc4QpQRrudrLi/clp6Hko1l+EigrvI
TDhkn3HF4VUBW0+CW9MNluKIeyhX5FV+Vjp+k+2ppBBqXXO3vb/FgWZx1y5Ykn3F8zx0OobF9FJU
LM87pmkonwzN1OYSOFM/yJxo9ofWkGhymd3DAhoBL+bPPkWUwGsZQAaOgOtKgplDqdfOf7I9itD/
uGhPtopV40kXGNO+FnTM0Ws3OgRg3ixW1l4ZHN3fsXagY4TnzVzMymGSF4ixeHrWSQh7cJH4zgzK
a2On3Oni9R5sfKWJ4N7Rvi9TsxzpT/mjYtfrg5Y0ByiJ6WVbJtMIFfgeZKPIFK5wysbMiUIh8xHq
dqpAY35zpzp7pYjvYDZ46IN1zV42nZdjlLlW2aAw4iKYyd/dSNjZiWxcH496NCPEYvv6nanrIvUT
9xcIu/8EclAqBMu1wF1NVUsfL+neoaKsNUjipPlrjsfOuAmQE+RjpOOZPltbsyiRpeGhDLhTNU07
0hcTjIrffCoKSx/5y0V89NsJMQDk5mJgBy+xmmW1/cctC/79VMYGIa2YSUD39OfE2qcDi0aoe49L
l0aoL6TBVgec2CIibog8duKgfeGaExp/w5ZOm51k/4WWJ2JJ+OzhyIvlJ/Krs3ngyCY4HR5zPSvx
n+9OLAyzxLv4NP+7bi/QJV4tpNGzAnijgOMzMM5ZhyM6RYCdti10P5ZaeTxNfMfOwDPpTJFywUdO
P+2g9NrbCgP6XRUmChPYYZkh+f28DxeNM/G8EDc/AbVPS1/BN2WsI9+MQ91gMga8e/x+m1NrtZrA
1sdiOjrX44zVnYl1qeRduF81Esd/7pvI+HD6VjEgT+6YZ9vsnjuuKcKNtlZT4YCCjxVfbDUqgFyb
L7u6U2I3SPa7Xl+ie9NqcJPKiG5KXcZGUX6sz8ouyea1lhJsVi+Rr9JuwWIDkelAtiPDaJllZEMl
bJedkt7nHOG0HuaWnKqgg0RGJWuCOx2GQyrS3Lh2Sa3HfkMHhCf+ec891Xdqu1yh1TcK0mbRnMFk
ss8wyQf1dQP8gs2t1K0zA7Qu3ezXtBHMFWa5KnBWiqI4IPQdPWwA/T/Fo+NHr5SDJnOCIhxXC84l
ylXg2OFaEr7FT5xNDLn4D3hk5av5EfREZEzxl+adWlUD3R9h3xol5nYmZB4XVwKtUhji2XHIUBvL
eAw9waOaMQzcg8XE+rjIg7bK6YtjrIy8x1Qsbb8nYhDGVuOkqtva34gxwY/k328a5ReovZS6OboW
dUFB9hxwBY1+qi028JnNevVayzOB+9JByQjGkkOiU0EFMzYitEeNdeXxGhp5vqieMPaG9QueYQnP
+ee56EsqsBikdE0TJheBPNfNJHQjjrcNKA2qk8OX2cFPYcwiY8wnpLAzAP3030W/kmCwWJjMy9Cl
9MbQk03BcwXxWOycnIjT3gI9ngPPBVKcw9yu84fBFlRJelW3LB+TiUztgoW+dK3RhAVjXKIRkzC+
EC3NSnOqTCort5InPqjKO7DYchACGvr4ElwpRYiMDjU6gp83eFPP2zi6iFeMOU06JBw00kas7GtA
G0jbU8ZxABTSuguL1lg62+ZJEcjuxsWxymtw2iA2oXuzg2Q+XsZSTq5nnlP2XAId3hwVJlaBf6Hw
kWpMpdPHYO/cNdVZHARFhHzemYa82ppzCwZFbb0kbJ1cUgMJ+ExH2R0BF9XZi+JRtzWWekxCEmAB
oZIDg+7a2WgjfxCAhdLg0bA8uZAaDs59gym0kY7xttzDvr+ZX1Y0V3+JaqV3pDMB5YIpEP+/T4bm
oxVJdYD9ieEyHjisTi62gAB8DwCtDTbv4ybdJlhqQYdRL3jknAO1Aee/g32DepPoBTMDpL7q76BM
vb00lUOq7oUnQqCArckoDZONCPCdG2LzfMn8sCDp18NeXSSr52JG9XoDnGorrQDgNqOUTxLE4aOz
sIALf8i+3k8rUOR43HFcrCcrihTY3FQaORufdtkNMn84EwmZLovP4aKcw9D9AVJsNTre2eT3ZkQz
sJ5KK5wk5baqSz1we1H6mJvxtS35NLfgZ5y4NUERXPaUsY98I7GenEMkWPNns75GDEk7U+Xwabak
XQP2Y+KmzCUi5HlGXcp98NkKDN7lX3E6G2bOh6WVQkVvO9pKwed1RgC9GhFH2KSVF0x+m2o1mHUx
UdZ8PFwG+gR37x/jDIJ3Ad57KHR87JSytvS3v9hwoNCj3LAenqngwg7Kw0t6Q8dtzQVgIOATmr3n
N4AudhhT0s8Zem/Xw5u4oiUto4wzOp/d5sjw6LDCFVMMMLldYUHSMZAhQAmmJfpMPFnIhDb6VBkc
a/h8mKDrZkdUds2ENGoPJD59CrZQlY76N4ICssYRMe0NvOh4c6XNjkL3o0FPYugFoLCdZ48SVZAl
1X+Wo+aOaW0c8kwegij9djDzsvPeDblKUc5+gnQ7nzmQ01uPx/BhU0ApLvIBdKKaWJzRQSZJWm0m
5YwEsnNWPeP7V2lPrXvApgPVrxvM9+J99ln2CcqBSYyqESqI3d0v705oz1spGCJGWY1rmZtJ7Prq
k4x+MJ3CXFZlfs1Em/HILxa8aXkrw0qt+10W+tvDKmb9SZzdOSFJD47LD+EFXTJI5bF0TOWrzoMZ
dRiygAYpoFu4IQDvbMN/kdZdpvmjaC0mpKIFA8Oa5L8oK+3DXeXNmxj/IniE3hkpKuU1YbPEGPij
4EBOmmQBpZSVVZWLMwrAs9lqeRIAn+3vjC3IZZKKCEMGLJGpoXkVSg8P/y65qYK8sw/CHOpXF3nW
H0heVBJ9iaximle5BLP5mscszrW+eiZcKHyVcA7pYgW23qJOOpdUf298zJzsqmJQ4w2eO0CrkD6d
zeX/DodJ6baoOb/ZjNYvUAVXSFfQm1h/jERFNswplwBAnIKeTj1w4CoIQPAXIxcI43LTMQ6N9I/L
kM0SPTROrrPMYJ8vJrHuc9Y0zBjCPN9sfk7DV0SqFs4zoamehvI0GCEtEup8rFzUECmuGiC1o5FC
yzuu07JLGXtjCk8CX0BpfibFw4UIcxAIqZZcMl2MdzIVKWJWYvaySMAVcmPF2r3tVmXOYTeSjAmG
b+A3MNmciLzDrEbXAXJuxmXjl6egliAThB7R8R+6qjzGp63grdME7lgvEkvRFulXccxqZB6IaCY3
bRvAuIThkzX68DPvaBJlJlUBRN4d3sqC97hUW1uZdFRJBGfBISj+w6OtZgFgVEPkGtVzyHs2hTVw
KNoO1GQHQUMZd418QtrztrlM8lAVQeRb2f1PGndFCXXpRclSDkZgA32RWE6Dx58IX8e9tGNhps3k
ltOCJvnRsbd50u+KFnjLNi1fJAZusZQI6bOIWFNuO4MbI5LmTabFP1Zk+smltfjsvmSGkEQOKRKY
eWBTeCSeIo6VhzN7Bpa0Ni4KT6E429wWoZCg1akZuzPlJT+UefwIik05UsTPgTth9vDyB9vD3VDA
ZFO8fuG+at6rx/qOrbJieITbC5OnEgGUMJU1odHFvEKn9ylngSgDTv4aGuh0LL7iCEjtBXYwiBmS
TYCGXD6lKZbqxcfPlO/sY5uSwM5Rgj7D4wz6uMvwI0C/01fuQibTE53hgTB3kGmE+9/uF+u6Cubk
TpnWU55EI07waI2JGftwB7hhGRcuuOWTyTlnFestDk4qoa6reYaRf3rBaEuNX5UIPIeC8Urgu6p8
nzuJshTXM+UkB6GPvVI2bWszEwgR9oUQeJCrgk6niVUswq3kw5ZMPahsg6hnw9U4Cwy1WoVM44mS
UJM06rxzRpy2Y/7cY0IZD3Sjxvde7oYWy5lQ9DzU8q4n0ijjcHiNFjKcMgIrKavvg04JHkbC52zy
a+LIiKGQmh6ErY5N6dlSKCoghKDNWAYaXqB7uSZ5x6J201iIX8JqOgEp9byLwKGbuJmeEYTLCFPz
u/aVo2Tk20MUqQug6XFeYwLfNnfHoes0z/a6gV462iYefDq1R2SOKuz3sJzYNSGhcaA9rImlFh1C
dsK5lGykvqjbPvAf+D2XvgO2SWgFP0mMh75lyV+zd6nM+NGZ9cFtOmeRq4c6umNwB5dfozilJiT+
6AeDubPMHF8cAX2XIZ0bj0h2p6Mz9kYtS6SA6/dyu6IS9HosrMExD5UxEqbCEaKxEh1FEuwetmiM
4Iap/SMeZIMeEll4FhZvdEk3/K4HcNwGX9a3I0cvjPAoa0J6TILRuKXTDOXn0gpznuOwVmmSYcFu
6NsaMTh2axhALi2LWfbmD62cobQwD2gOg+7Bt3sxUCXPuEI762ny5ReES7usl73LF3M93zsaEcav
dbsukJYDt+zbI4OmYAzCFsmGug6aSGyuQ/COZAnGoaIYiLMLv6qVDzXW3Hw15hdxDwu1JF9zQSAT
dsfmKR576bs3jRNrKiFn2h2gCD5LuVDkuGIabNaQ8G1GX2hKFj2StlRSgGDwOlCmcxsW7bBM2ALG
Zpf/V+9I5A0HZG+7uF8RUph8xeTD+b8j0oFrbuCgOTxklYJvp7c7Rb1D/GD8yPizfnFADmpNN2KY
wAQYl7YGuPVk/7YQ36rY9VZcBv2J5b5IF7EQTvrYYb21VziF+08lIKCTYNv9NGBrXgNLsjswqmBY
qB9GLH+lqY7PG+oGCw+YGUy4dUd9RIRYDExFqaTW7d9iCmgX5UEeCcvZVlab1bhJYmSgSq6ohW+j
QjSmf7hRDA9MFpu7nUdiUy6YoLE23fIQ9zcLC6F3geLa1TSI2QcTxaBcozVnmit3NacME9sA6Sth
utkNKq4G+WZzCp+u6feLKHEOdNZmrF28/FDZbWiCM88RE7UtMKEvoZCYHxjpPNEyXOrk4+i8XCEm
/8I54MB0jifH27X+8G9o35UrXT7k85QJO3paO9I0is5OMJdG8YcTh256Xptp/hN4WrSdBuQ3BHvW
gynT+3+DpXkvkUEOwe3kHWTXRCgsr4ywPQXkM692Bg1k1VzgcsUy3CeI+H9qv7kjKfnCGP/MKLAP
T0DBKj2GyndVp4D/O/zf1WnBuleBSndcTcMIeYyEuCGrtMpUC1y/W9yPTu/yvueuTuK5I6OHNerh
F+cEWN5JSGuZGh0CWsGoMApiy3eDrHoDz8b4Qo6WgWnK0GnrasorF1fknIRorha0pHUu/sjHe+Ao
QXL2yXaTp0IvcDGDhrRAd/1J3jgV9Od6zOeWHTaZkjl5ciMJCXl8I536mAUFQWIHY5+SocGhZR0o
hR16w53DsxMFCyEwqJhfxXBmtA4a+UAo2lr4MtWy4BFrcHJmWznBcyHxKYNHWuy1EKWOyzCSeyfl
ERyaBTPIaUo/vJZXrxn4m/H10+9N2jIVWxAgOTHWM8oGeZ2KiHkqkqCgFVBjXJlBq56A8QlAjyDL
0Cx+OvQANBpN3UWj0zxdQFHkc/kcj7oBmPRiQEiJSdf6PXNmoViDDXsIKXrtczAh1N3/kiw2Lh5S
reRXiKXDDvYu6V3+c9eUdngFzABod6jmA2Qa8NTGsXqbTzkiSqzfM3sofHx1LJGECWUiafOz//j2
sSzs/o5wi7x/8W/Jumm/sdCHiGm2ravfrs4Qmz51xXv3IvVHoukk2kMEnzOm34T0nRNXDtjUxiwW
zprCLOxgl0gl6ZIHZWlYvcups+9eBmVlreF0ApvOVhVfDjxFxFpTurOYWMOGI5bD5Wb1ixTNG5gv
QmgI1Leu5s8XWawhpPpPMda7UdqpcAORXwqHslw//MFVgijrkOzGisKBnYEsRKQmO9VQlMe+FGcr
qDaItERqzQ7gdTf5gBN3ALVR5rILhwKKtcIkkG2I8IdGFCx4AE8cRf7z1N3bEFIB+oPhB8ggU9Ij
zILCr5W7WMSH7e7HIhPXNDV5fMzIEpLqY03P0D/vJohfWHWE9tW6ft6xBQNwQMFLjSIQIISIuGiJ
G0li9H21ZShtvjSdtsWqbdQrJdZAfn/iF9l0azi2TrlvKGNDtCWUa/WJYTWa6A5nvuODjqVQ2QVo
MQSewGHk3LiYwHZRZjfNDcfElKKJ0P5oLCk1X3tv6DhsPjdVBYxNWe5JtDCHfcVm0zNqyV/yn4I6
lIDw2L93ZVGtvzzi+EU+s95dNGU+6l5Q2DlTX3VkvIN3dqowLvtznH2/KwIimYNdykxNhAvmFb9G
UXK40JrOFw8SZcJbaU7I1+z7PsScHHiALzdd7RQc09mGKZzcR4LJCmywkZUd7mU85ejIx2Sr294U
cJwM1dIN2Y4/DjyPzmko2BYAsKAwRUBLRs6mcdvCfTdveCXR209WF2zgWVq3tV/Nfk547WZQNM6w
gW5NRFPA4kgO8xileub1vQqgRIFd2KEm4z3BdgiG0BQLgeDA5oQI3K6J1BANHTaBNq24guyPUQWR
KZnz+WIT7wRs/Ne7FgCREA7k9HjIsqX8k6Z70eTUL2uV/Cl3iK7+eCJjlPYrsprDJg6QtBfaEOi2
PzahMC/ujvTN2Oh45ePz97L0H7/VvLaobTVygxylBRjevWnUGkyP4gqwUT3z+LKhI/CBHqPONlPd
p+8+YCgUPDcI2ZK0+tZBQd8BD80ktRmGy1sBDOL1Vg89IKtiRKsvOhcF9j59JIeAR9ZTsxj3kF9D
t1Fjnbz/6Ngtw4/8gKeQibmoVTiZbzVrFP/Z4Gpghk7ABB4lXyiwqKuvYRyk1EMecrHmsUqyevHy
d1J6fjgzFOj7bcVbXyo+dy7v5cCOYQ8tzGqMsfZYdTZ5SZZHqLMwE3IVRyKOZiQrMoiA8L6WDN01
YCFpKXbBBusnWoEDxRoar+xbcjUEJesJZ4tgg+/aI4NTOT1luM5ceJgmK9CCuMbZduzxZSTBbcFW
KbqECSm83TIacyux+URVHGb+PAIGTiue6idzr8NcPcOf5ESCuT8tCYSqPwjF8oWByi1BNBmRE8hj
mzmKNg8Fwu8YOnZXCXZdQOwQ2me/FXeDf6r8aKwTxdtch7Yfw37JEQwlfESonaB7eHPc02OmNSac
fbrpjopVA1FTvzLjW3R97zzupUQe+kQvqAihpFnu3Lyd1/kyxwj/CC81sYCUXvctWHDmL9QORubS
bYOEGQPfZIb3Wb5QdZYp8OZM0by7x0QzLleJTjqHnawlozA6GiHgq6EmVfeeUi7pzLrLWolCGYJ9
Gdtv/ZNPHfaPNjfuC3Ki8s8iYhbYNS8JY92OtKnlAO9Sdks4UVzLwfBp5o7tunk+uY43FANZFvhj
Pt/1R9rQ74bh/2CXpM4DXBdE16oJQhstEd7gGPYwFlhCL1wE8xlaVUQX54u1XpVNnemnpqkQCAWW
b9fT4ZYsr6fgfp5wGhaI0hVBbcchGjds/tCeMXuH1Mlh4/pX5Y6/LxWsBdEpxFAJXnq6A+ty6d5p
Qj8d5YXGtftwJ8e6jDopiY63w6lR7/ijBnNSSteZu+ALiX94Qw1ybxT18EwDRLVScPt9jHsl/ldO
r1X7IhfHzXsc2+F0EP0bOCPu+bAlkMKnXvyaiUCQVHKdHc9j+/DwMKYYeuyRCcB32zvFFnTtmBsT
bB/alSaOdjVk/ol7VNCyh81+uK+wHGBX5HNFtc0y+mAp+qR+6L071r5Te9YBHlupuEr5KFtrBe9z
JmyZG25AftD0aStIsvP45Ys1HJ4eutln4bxJY0+2v+8H0wgim9xueDOOUh8LtWelHOWEYdpPCreW
kXTGbbecpUVIne+YSC0b4jxQaehLPZtavwXqMkoB7WphW1KQFob5qofaTLk3smI/crF2QhixbgKR
Q0GNMWjYMhU2PEw3hce60/10Xoa4l9P25Rvm1Vi4l5Irl4VgrfebDfgjQqNFbvgc+zS9vXREYpcw
iLoISiiHZQe+I+1b/PVvGa0BFu4NUnZSL32FUhPJSWfzcfb8p+mmfBRp1ofx8JmP8FT1F64CtX9K
nKsDW1nmzhUfyAjjN6YBLmPp9VdcKTheE1CXMuFqFI3R9ex4lPSILXpF16xQpymcOAzEtG+POw0P
f51S4mFbddFGxK3rWmiuoo1h4Fr7RfZBm9BEdv6TibFBl7hZ/MkZOYfwmS7AbdGJl+XAFE+ifmY2
ufwa7UHF5mo9/1zPrWLugx4iRWfM3pTqPGPZh0+al0PxC7pQVa8iK0gUY4oMEWgLlTg66AMy6KiG
IZLcsx/EQ+zC5yiasp3csPXrZ6ojMEWIKBlLOf7zvuMGrUQEWDqPi+37KbZtXwSR3W+I3xFXMtAd
oufAE58nzJ1zplOOEMKVw38PcNUIDzpznUa4gZxnBrD9MPq+NoHG4iSj8G1vd1xmzPvydPXiZ1vN
chdqBv9+fMtYjqoCzppycB75MkFCYZDR4pfECyOzIym33x6T5P37GxKDjqD8KIppLJju+lRhc9SL
Um53KVsQpc3gsssSfCdbol8PnSKZfT6Q+w0xDItxQx6GNobhC17xBbYGlu5Z726cMT9BGBHmjLtJ
u/hiYDwvaf8Ye6oewt5mX+MxgT6LIIJHa96cMgmCTCvraUthwz2hy0SoITh9W9593PBzgkk84knA
2aCI2Qawjt20R85EOkNaU/SO48+27F+m5QWlkt/W/0HjRPS/yXBijD4++CGzdvhojYR1F5P+hWoC
4CYOLpvmvxQdYQYimfb2ITsrHCvSIxBRqc6sUHMezolaMGr+mNos/vrwbp2RWHlnwUc7HIx4ZlPo
G1Igx1Hn3Wz4A1WMEuat5mfFSvbTJkb9gj7iUqnYrI4G/bRTvIM6LljK8cby+K/My6NseKJMexMw
Mq4MKP+Pxfk+KsYGw1ik+31xrn77DUGIFF5om0otxropQNnZL1wSzO74vUPaCCpuZbYaHkNRDdBE
B+9axmWNBww/R8GVaq39nxDc7VHK8b1Q2UDTP2LeuJIWp2cjBGW+YdrUgN4sy9XkmWazYhk7ClFq
f+vLUH3tEepErTVnBKghQSVpahg8KwD3gBHrQgCnIYk2XcMwdiXg2h6KHeri5rzWs03NH0Xct5V6
3VidBIcTcQGrtWmH6AYTUn9T+jE3WNiV+DYucMCCeDHGJjNdFAPxCilOjzqdEAkLdbf3AwtawPx2
ZY8/VtrcRurLbh7uqcgXXtQQth8AF7sXsUACL3jIfVIovqYoAXbR9VNcgYyWYbvYfRN8t3gCdaGx
vwVHUMzdkLl+BOf+z/wP9RdZATuypmITq54lT5YmE2HYZjYDPSZsDioo5pAohdhlVk6RL+MY9Oh4
1ut1UCKeVDd9i2c5DujBSiw7Xn9hbNC9aeyTnCC3lX4XmZdEt8UvMGUTEHcpAzsGGOWBsBs8798V
McVR7BfzNbDrgr2CLBWhjXJzd8ltz3itv1yoP/V8DWLbWm/0vC+TuR1FkLQgGpWE5g4JqwuIZnEu
X5+l8BIw2gKgQe3uzbFzJ7ZC8u8iDsI8DlF5sV4lpWk+zFkIDSYL0XpGJub0in3IpBWIe3di+v78
Vl9mPEpdkIAW8jTuBxVDqD1WSP7VsDCE9LWyLo5WLz5tN8CahWjYFneGu5QQZrOlIhQygySqE8aU
Y+V/Dn4K1Rwd+VZ8NQt2brnEaAUxhGON5r/fHnn7doPVtammB2JMrCmkIXJMCFEbMCdBN+yHTsUF
jcRyZyuxGmKoIq3wYsKsomwJn2UGDg9vdjtOEdy4Y4tvb/6AlpXy43VQeYcDMwpkoA2IrA0hlsMX
2Rzaj6ML9fpPh3zkZ9MapTM/0UCueKznhBZJWnnBYFfRGEe34NbGEbLeG6gZ2SMoD+GQL1yHHCkL
LUYH9zEX0DiJv7Gdypg+D3dHHZR7CkG0OnDECI5ug2kCgd8VNSrlXfMqa39hSuKwX7n1P9DKV8oU
6Lko+VXtz4seVKY5fHgK+TNjFfMOmgU6i6rAtiYmAArbt2B90YOrtsb5mpfKVU7X65lmkqbUCxkN
U6bXL4yOx+a+ZqZOI/O0p8vauolD1nHjlZdtx7GXJ3j65ZULgt5pt4DHf15XkXWHS0hXelyspkzt
n8/u/i0VjkDO50OG/fpGS1YPyqjB+HhbvUbsoXjC2TCXd4C8yaXbb93VJOak9Ylce3XIUdZXDByZ
FCX/zfgkjZExjSRx/T+8OMK03NY3CBjBuUNeBSo6fyjPHSqsdWLLgBXyl60oajW8r5EKaEuGonIt
BOddV0O8Jc0AgB26P1tPZD0bK+xbyTcCv+3kBL0Jknb/0TNo6YYk1J9YgC6KOuU/dhr6+/VmfAWg
me9qYCI/5Og7usqO+k8Py+IV+Z+7fVIagXXqJ8FOeGVEt5+owHlSd0USdRiSmUttsLWrX0Qd/be0
d8BVdySrORMx4gi1uX2FsgWjjePePja0hNOKpX5WIKlfLJy0tsDWlLD59MhR8KCHzzzAJyVdCoqa
KLtlJlTN+ialuB+cXe6/RIGq5Wp8AxqXiMCPW5bqTlgjcssMTQ0bEKxNTPOeGoRZGlPhdsiTCh2f
je60UtZ2KyMzk7C8LHx5VNUJ/IT3h/OgMBpqrZHGsIU3yHkAKCnfkhlLlKnHsIYV1DU7xVq7sWY7
+VR04KCuYykiYSkAwz1v2cnrRahUUCPLFBsRrlwWuNywjvw/7ncMhH7H/xbSBSvvfHDoVeJkHyth
K+LgBS0pxqC91w1oBI0abSH2ZktrRz5VU50QAo3fRR6iE50pGr6SQUXwIqgK4sN2IjjAwomdnjqD
eqOFlmdMqNU15HZW4Dv7PNMnMf1w8cWKgU3JRPg6HMugcaiCr2oisQ72SFm+/M27VzpwvVKVwnHS
OY2L1dHrAwkR7iw38MsMclXAjPVjbk+ZpRZ3nBu/Rim8GKV7gOPtHjp1euW0FVfllaznWCUGOy+v
+NkYY97p/fnLAM7l687gJb6tQHbNPJd5lZ9n5HlBJAdU2KR9gi7IZZQ7ylwi3zXdaO4gLp2bu7To
ETzduorbJup3Avk3oSpKWE3akHTJcYqC51aoSsQYFqEEmbDk6is004tzzmF4xAqJjUQfld2LXXGz
yDCu1UtQqP3KPYIsSRHjLiEnJnAEcxgTl7ZLC+7iosCXUIN/F5l8BxHNBduUBYT0f7B+9cgup6z5
Peg5sSwT3Qiq+fJgEJhZJiwPjAGKEMjGFv84BgafUVWvRtUOUuUIOeLsPnZ4JLSgLYrgfxrTZvV9
qrvlmkU0H2Teyz17+d+/NgFxVcEX6R3mKtk5teux/+JJfgNOVtSYO+ybCHqGcLTa6l88slPOysiO
tRzQ4Xby+l9F8aNqEwfsGRxpFAVNkAtThcqAxDd6gPOhsJJB5Uup4XlnwVG4s8PsCo+4QWZUzH9+
ZM692PiiSGiaWp+TliAVIiiuEy+334nWIf8hj92icP8iyNxMUwpT6FSVz18R/SGl/Lp01MpoeQVN
PePSyrFfoP6zkLfWGB94VlF9F43/DziGTtrfr2//gxZyHeC6bl42epit7ARnqcsvFIbQPixfCPS6
musDio5npvc+hYEL4dD/bAdZgksrUfhJ/uRuM75C4WuwSF73CkNKyKyLs8BcJWB1JfSAOlpb6qm/
ZSvfhraaitvk6kEulfxEYpH+4/vFbdZ9Giy+EVK/dpk9cZRwz99SEBlxKoYDrry/jia/Dn8eGd1N
S66OCz77/ssSdabBVdD4mukWRc+Pa9zEiaCK+BJ58BaugHm4ADtjMZIeQgqwoLWULgFRZos9Kpln
AGeHaBFnvClg7aSLdQnLDNxl6m82rrISKCoqjtmTGuyYtWknphaMrSstGY79m5TrUs41tvuzE7i8
4wdxkmtadoXfZT/rcpx1I2wMYdAKP7YaKnYIY7MHAcu0Ezm4NZZc9JUjK8P/xZ5VAMv/gNqJVG/h
CyEzevGSImFGbFjIgsKKOrGbz0RSQ2umFQC0qTR2uzKOqJYqCO1ugg7MOTuhE9Cvb1PVnUtKbOrg
B5R9G27jtzApSQwiw9d51taWNy8ugrUlbBPBXfMYvQvfIe/pKBaiOYpgW+RVnCTECyJCVsAEoXNT
3G70R4gBp8eLvMSy3xDThr48JmWvnH2FXOGS4VcBGmKpW/yw0JmTPuQsEgrM1XEOx4e/mcUQk52S
HwviGuj2BIYY9+ll3HMAY70i1IHIwUzFAHzRBTo2dbPR1xC81krkifuEY3NqNBWjcW3YVXHJV9qg
EWvuhwoMVFM/ViI/jfApHeOwaAGsXSt4hcm2TfBu6VzOB5up8BAqPG3gapY/EmAmHvvijtdtntBV
o47dP2T8BAOfQYvvbCyexxzad+I8Z+VXfKQC5H4TUWaJVziCtmkpu6wQXPTF/0fLoTMaldqyxrNm
4ccDTiAsfo9ika3CXGG89mxelA1zgKlWkStbiCjWAHEmsJ/5O5MJ7Hdg7LPERAgWlHCLLA5Ftnjs
6PyDUstE9TF3J2JYpAVZxqjnN7Lmp7cZya84I8PF7IWxI54/EnH72aYo0M1HqygsU0XFbpFInEfa
NJYw6WPWqKEfkRbdUlJcBlkq+eRg6opbwToZ+6K6lgfIsnY8k7WX/Js5RaY0X5z2OMMRTSHmWRSJ
sg6xBWMA5kf4mZvfqJWOCj2dAUWLKrtWMm20+rODgQOn+TkpaR8fZVNZ/lOr6R2bMIhLLKMMN9+h
RfWQqACRvtMvbwu29PjcWLxCLKlKgg4Noc8QrM89psy/K6cG2/GQALa9YyYqyg2PAtbWCIuTQuxU
riGXrTStLRfRpr+LyvPux6E5DdKZ9aFIGJZ3uCvTE+o+UATAqYU0iSx2nSG5mNHw/cffV+sP94c0
tVTAZrfMnZ55/sVPRslaa4Idkx0TOwg+FRifIAkjMTg980evKES3lwXQlI80PsqstnYCJhU7xUYv
1N8OMlHN5k8tPkNAi08WY7TGXwg23eF9gQbxQZyx3ycyzwq6MqrSCGwWZjxWXAR19S1H9jMzLyUm
UNB2pKAMU8egpNwCgARtJxA8B97v6r8SjqfML0nahfQtaSLT4fctcUbyR8pwqncQi8t6vGYK3RX6
XRf7Lmhqg0b9LYw7shbo3bnPa6iEPyuNHoYm6mKwKvUXnOz+NBe+qkQrV3TyedRRY6sSk74H+OuT
m5YyORO9t10AYVjJnyvBj1TBcMofbItiDR3A5uWrBWLJaz5XoyFt9u0IMJm3NMfMxPmx8uG4OCHY
PCOfVxY1GuHp+n+/wz2DuHOoFuZQp9ySgBijay2uiJ6UcpDqYKf5SsqoNTvQzDD9D3UIST1Z+GPb
VWmWf3y9EzJtt0T1GzWr4Nxto2+UW1plPWPvJOVwY4zaJYW60G1SD1nsRcgMdHNIfAn8U/G3/xcZ
K+dYhRJ4OjRK7gPObI/dcXgYT8TVH6SjZYm4qNZM0EqNPJF1DfZVxBoIujJcOEnLKWz/mnGxxWgd
n3hMxDNsLVUW+SIR7tx+E5CHrOLDFxG+acbBKYTBWHcYViY7Xs8x8rcetkrZlZtHI+kCQCGGCtRj
AyBF6J8ZaecJcImlOV3ZTVojAJnjOGh2YNAMPlIMWe8EVdr3/caTdzMm8x2BH2fMoN5K71eR0Jcy
pY9EcAqrzsnewxZmiPCDxWXJ7otfa+d2Gn+q5nJ33bspjv8Mnvnm21zRAeaPeSS5Hl6n8TuS7jUY
jupoWsn7mnUjPOQfoZdZYhOqgrAgXHjEApoMYf2Wolt2nPsgTzwUzm2NBWEOe1h+nnXagDgrUkrd
fmfXjwEOFvNIDDAdIz4oK6+S4v3Q9DsHBmnFpc3H7s8XbN9HJVtPPJayIYGYYVH/vwFlNPWKtvZF
l6Hsv9qheBKMJQ7JkiojcBujcMPBZNy683JwxZovGqwFY+AmvgAlF553G+JqW4T4OxfISh4swCsD
JW9HUnitm+5RfccJxbig97ZNWz6bXKD8PJyfR136b4ZL4TD6gdx7w7Soo1E/6CDRQ0EqkGZXtrQu
Ez65AiYncUtThP1e8QbXMkffLg14RrUK9c8vKLB5IlJS5RMRs4xkxZo2qVsIRMz76broa0ePHvJg
KgeDQ9ulaTPGiFIZsHz/tjkaKhnCMQQFvdydMCCuHmnP3D+2J1Aer0TU2hNuXfbrQ9Ehy82iKsuS
DInXculjJANBs8c6qsNoCl+TtgWOrgz6Xo9VdF2aHlPRCPGDxFbKKiyurIitFnZ8JGT1eBOHEohC
/jX1VVX4F8lJyq3QyndyFG2V7HNPCFCVhCr205MRKA4xEsjBtwHZ+AyU21A7dK5JTDF4H/96gKuV
JoK2d2RRcSDF1b6PMDX3jxdzEjg6M1ucnB8SEmADY8iRR3DDgo+EZoVdICP0Xax5pMvv3St3jE0n
9ECa/Klt1HYo9aYZSQPJCFeCI6zoZr2QhUEKrahsl9D1Ate6y9AE8F/hN5T/mnxFOwlMN6kvhGkK
t9qgRblSRRn4fTXV8glamCFjVXpu0bmcYL4IhwEI/GDRvPWJb0aLnbJKPP+xzr1H5tZL3xOSb/XN
87kyQ1LxjDWPSQ2KERH09Espga9i81QCDy2HvTwvwVdPKcgCqkXHKiIVhq/IQEQpmZQ91G+lmodt
E7bhFviH1fmdQWGCNfhwG0FrAXA4Fz/4gZUnv8t/OKc32T7EE3uk8Xvgv6elNxAZ5gGqJQUVS27h
7Ye0VX4ADG0/X4jKtOeo+VxfBUDDuRSXtjaNmjcQQo6ClDl2SSz2cm+M0XKtMTUjzUHu4WfaycE5
Un2fS7lygjjjmw6hl4/Uw/qDsLD6eteaxPiEOSs5zWS00uw+ljl/FC5d+vp+CoHolPq3t2VLLBdN
5gDZArvf0Tzpk6EzK5aN7GFN1z14s0N7e7DZBMLwX+RJkDwqCs6q06E87NBw5epvMIo2uylvbTPQ
vFUDasn+U9tut4q+53UnKPrXC1Hbwsc6yN77vP0c4mVqMIpxvFIQMM2JR/URX91jxw0R4rRdQsPq
84dQxvlA0yQwPMtA124xqVCpBV4QZIjOfMG2NPdLkoNiR41e6g/9PViDZtbW/PSArGUWz8Da3u0S
+Ff7UqMu9Q2DG8eeezFprV4vbBMJsJU01367LohYUwAHYZSNY5RGiUmL0PXlbSNL3tYdyRFRz0wi
xzJrCDH9r90R8F7g0knsU2Y8oRtvVY7q4lAuY46fhg9LRix+eeStbDdmF6hgzjIXSZBAgVB4CrL1
4mHkywr4bjuZIGYYCFPDgiqWVFT95z/6lRXJITOh+dnDid0q7G1NbZ/gdt3hEaZFYunbam+tfBbz
T7YT+h7U9B5/z/ny5DwOqtm8hL3KMVqRbiimxjZvA62qC9IuG48u3HZNR1eplbJi//Q3jpc5YPlj
pupSWDU/VP7DIKSzteUOyw6qzvQ324nsE/O8ngyrMkuOahVRgflp7kdzfgiar8oT9MbCGCG3DVA3
yxo1v+t+cV1g807Xp2WstQGJ+vCOzjBbyeWfXMi98286dCUet+dAhexOotHjHHNirqt6ppspaFd4
oNwM4nVtRdG7shX5e2w6qlssBypG2x6GVYtdB32WVZHikXpji925odB133L81HY7av6eYSeAQTsa
1rReGW17r7QDfu4xe5nZ1KE3BzR+76QHzvUmzXfYN9KIa90fzRikvvlIzrq/UtKfR96hhcflcSe/
Mop0M0tr4SFh/pxKaSz1dXTGjMOG3tgGnmV2LBLUNj6oVBGeYtOblz7RzxTxh9CPOrYOJJKQUQDd
vhomB1xPuMUQqIVPiuum3rLttUp1EIvdhJy4YqNSxwoAh2filL6yVgGKWcpWwNcwcYTzXbFfx+Z9
6qGVgcqOYzrEdgiGfRMofOTe550532ha4g0XGp3LEwVwNLyuu1yy5i88yNtDJi2bonXWS6c5dWVv
kX7nQtcyBA8L3g3DXYLPNBPnkiOgFRwzAuvh3E6sh5PoqxY/1XmMvXuGInh2Jji2LKXosP6NuBG2
ddTzDEuO61Wk8kx8HziiGMcMjLhzjLrwr71dqHW7eU6aXX2EwDwajBxW/vxr8G2p+oNeef4ulaS3
wNBhmo0agMbaawt8D30sfsHBw90x2CsT9eeURpVifWQoEIfre458kugEKEa7qA0So3vt+sJ5VF+M
oLJk5CGwwhg0YbJ1sAOpb5bfCAbOUdcDnHhApESs3IpBTlgnv4vnG9zlt7dpaUY5I0gG6WErSM2Y
scPAgD/KBU6ultDmH3jBt2IAI2ASDDnE8UxWtnGIB+yvtYnNo7izbSwZLuBGz4Fcupkg53BVtBK8
xIoiadAZabTRz+aASuzG7Toeq2oTzKf/Ds657gFeuB8BRv1VskzfKAKaKJBLT5eMKJ443TI7wSJb
tmGZ5KLYU12Mn6TqQuyugvebOno7JKubLkm5DUU7Zs6si4uCYe5dgZROyv21q/WLJmBBZSQRJgC9
/wnvbLNDRvACW4e7KiUwus5pqVPkjilLKbPJBcMAJ+WZY/2s3/ufKZUVpdChZtQwQYAq4uqAxWrE
83f4FC/D1ZTsoWk+A1XTT6Vw3iaYa7kpwrwOGGv+4lx7JAlflsm+5w84EeUgrUXFVi6vy+eWykMg
1nyW0wW0Rc7USsfjLYmmPjF0+gNP+yacp78X0adPL+cJGXaaeKoRg25gvgyZK33S/E4G0iceEIne
brjdTwVocielYa3L6bhv63EXwesmGtMFl90TZsKoBlwwybn6JuDcrJVJaZYXZLvZYpa2bd3eSLwo
0W73T8NVKTTwcponkvrCFQr2plLkRefBJfo+vjMAwRLS7VEZtDcL1iG1FJ4TmSbSn1iv7utcttVX
ch0yCCU3HFHlRZ4fSngRgHFjcynUN2WNEoBUwc4T133UdctwGMHpq1JHxrPVi1fn3QwQ6DOo+DiQ
zswuLBnucAL3w5IErPJQYsB/1Ak6GQgKK8GDvlDq8EgJQG+iISRlpdb0RNHG2NRTMGVwEYGJM9q7
AZ9AsIp+JK4eqxK5ybVkrMMeDAzgTyWl/woGr9xxlkHC22AsADUyrHY43Dd6RPAQ6YYV2LpxYsFc
HpxUamlPutecZw8grOapxsYjYCKc7/v3MmMWNTiWZmcW5d+SCV3p8DZGPOjk3bvdvArmQ4O5sC8c
wa0Yukwj+Pk3cYX9veauhKkvDzq4G9dhI74avOw70Ebwqcos6aYD3VqAJ6I+aRFWjdPopjdkt19z
3i73z7bEkhjlEKZ4lNLpNJo9HLPlWauDpv3CQfsFGBzU8HsymNXuuZjxNNgCRmxY7KCYCKbq4Tdm
4kKMool8uyHwyyY4tkKbXItKr+iN6CHKmkAr0wDEOZNk2xlm9fL2wHm2vd2l3rmxDU5/iN6rBTwm
ZPK7DE0SQb4VmxSXmWMlQi5MeCwlQVocv37s2P0vzDNrhpVFURyrhym1pneBsfEQpzEjHA4I7WrM
lFwFI/FYKPt4ZLXOfbLYOsmh/abHAAOHrfz0yNVjlteVEsWPOoqrwBWDOyaX2zOauWYj36TsIORF
2daWlem8xs7OV3GoxC1zk3CEWRqLaw5NaVpp8SQlNVWD1Zb/2uJhTU4/Bf1kV/i57lwP8Qitk+At
Dkwa5tZbuNlZ7cSlxso7VWDr4/PZcaNEVPEW1dufHaFLtHXS5okB4345/1oCddMc1oAENOBXq2sy
4OMdGB+iyehP3vZyuv84LDCtZAUs712DlZVlkXbogDuSexjdRtqWEb0IB30ZBUTG3dO5/YY2Nw/Q
QQrWAgOzRJpFqLEMlFz4ifMyEr5NWQ85mp4LyoP9xkwXjfcAtdRa6dWxb+Bp79ppL8C7BAs6xiBO
toN9SDd++quP78h+nj3TLNTSArrEfmEllBYvp3/CaMkV143Cxqoso3OMVQuvjvxrm0UtRnqaGGPJ
IrVZJo4tsjF6+Fc1HeGuuYv5L+KAo4MNgGhM00zkx0PhmNDEbCJTY77R23+aUk3P6u68OajY5ILX
2xScd1BMRQRNvdVI1CruNPAgHXD+MwlNzVijG443sWNlGji7rujLSRhc40r8fkshRxBpOLs/8mcU
E0FF8ArS3eoGUVJCFzWQ65U8vK7BJya1qLJAfCYJTBOxu95sLBOalrg8N2GzLKsC5iOKSkkJi5kV
J1zFL5geqRW8zMQU76Q8ox1T4s/mdulWHDKr90PLv/8y9Rf6GrDe9aQjS1zyihHm9mzi1EFVBXI6
P2gcVLMBadgJrqz5IUkTErAlmi+bxGmJ9phgBhd07Zljm5o7eNsFfW2KaoAtXXa1N9cEJug/lG3O
Cp63SvT0EzcvS9CW/MSVfDoJ3Wqr8JulJfaq0rELJJrqSQDK3LEzkB73BHpJBe2c4pqDMbZggi6T
y3PKGm1umAuDzkkV1S1Sh9ooTLFgTTx8VORXdKBk7jFkpNgpljRlnN6Qsgwz19YTKjURUtb2AqH4
IXwF3aTXG23OFXFiMlITjISWL1Q8K6BuychrtTB5tUGq6ZRki7X9Z33+ghcEi19h8X46/66j3kC/
LMzKZRqkNpieoeBaYQOfiEzvAjfnmzQUCQDfL733RW1wXWe5WDvDMiIfakhYhXN6W9EvRj3g+1g4
SYuZFY9WU022lLvM3JnRBv/S13203m8kM7KDZVWKKLWLgNatwOMrlIV0SVqMM3tIEbBsFLQES6Tp
qTFB3ltk2ekX6gcYm+s7goeEY2BtjiNi+PEMyG91Mx/BbV88taSipHO6aLXBlt2wtNSXBHZsKTXN
UOZMPuZ0WTUgpoSZ3ooMI43rTbLmBnz2x7PmGLpx4NtkbzXAD7HJOxAuBuv9ICuP7yCzTu88aALG
GjOHA5r0ey2OZGTHJjkoc1zkh9QzlCE9LssF8vcyjyBjAmpacdEEf32Tw7rqvTy8V7vde3aWWGBm
uRMxySusbZiGmfS90kAb37hR4MVzherffN3Jf3w7RwNaq5gdB/GAyXYHJTnVGP6Ki4f/USv2SR8I
2bdlXZ88TIRo0v+BrpUoZNA7M3J9zGEG9FVtiTdlalLMrJ4/IecV4n7un7H4xRg3coh7xBUe2qlW
c82XsuKK+CXEQ8rB9Q3fu0XmVVENEBve9QFksllD9FO5rwvlkpePTOJfqK6gS3n/wLk2LRCUhpBI
53fRAGTY4CWIEjNXAZP5d6E7PZrLFiKNbmV+mRYqc9VXal8FAFB1sdX/DddqZjquO92Rdo4C2H1v
mLHysBYI73HuPa2xSVNXQJa+OAj0kUtm/S0QINvIbfH+ICsdH15Du8CddRQi58ULqwA43QZgR700
BMaAkyAMDDSjHHOCryPsOnKW+f7cxx7vVm5N02EZ4XDafpvHDgEMKHY/pgz6P4SclXoPspuzbhyF
9Obg0JHtq1o98a0ZueCv9WlUkLsxo3cuFOR8WSVHF92nZFsyI8EzcbGIZwJ0TvEPj8XKolKAv6n2
tyHtfxf+SPw3WmHGw4yy7Zp2GxT7oKpyO7xJmsdGM1qS8ob1mGLS1TpxbvR5iTo4mE0NsS7AbLdB
YO8JU6DdC58ho8uIXZ7BxrDArZXbzM/+Mup9zkTtZrfUK6YNyHxH+baDS4p4O/NuePYGTJk7XaQC
S9wGZnloF5u3OqyjYfoW6h5ABLAfVhHP+NOhyPUYsclmDHGhrtU7TkGgwLtPm6FwfwIV5/ZrX07q
O8mxm393JcyQWuZORJ73hJoFyiXKZLA7lOUQi48YTcBieafP9K4S0+saJx6uVSxFoMBsNDizNX82
kKX+RXI7PFxUktbQvpA8niwHasfPMSrstD2ZBLdWDTr3LRO+BkxO0G1jmLCpfW1koWoqZ+p+uBIT
65BZMoOxxoJA/UJRalZ32nRDM1nzhyCYXp6MzHUeA9puSGEB26ByE/3p7HWStmxHnFq3mtAAtdJM
ur4aX62uCY0JY/cRUjG3HTYB/4sjfj4q4mFnftat71lFktEHYRZ9tOcSOJPhI/Yt1N8smWMWnsXd
EFDGLBzF/7f9tv+ETPq+rP3oNgUsxTc7Thw66q0SZGHzzTvEV29gYbh9J5mhlTwX0QXtex8fTpEG
++ZYBYTETArw5qMCyvCOZ+hKxvT8pKBCQMBnz+MfjxTQgNn1i2vEeudhSrKUyJKM01OXHawbBjlz
LjrGfs4Urq5X/uMWKarFGMWGR4sMrUm7ufWXvfUH2aky7rIdsmjgqQTFO+mR3UY9qqg5Av6tHLP0
q3+3/QTxj+EcPYDIfv3uFIiajefn8+5W1HGCOG4I10tdtlMiA0vJFc9lFa8KxEcMZdptoiNwSvhn
2u0O+Iwa9tCCYuI/a8NBKi/XLODmWu5v5xeKmWfzyWhEjk5sBIOheEfMN39u3rkUQkJYpDf2ABlY
S2b18PZbCBNk7X1zWXrjpzNl3XCiReDePsdDxR4JfqRMOsh84xLxkQ4Zq+54WPgB2xoASSO6y8bI
5C005rpVJADM0Il2jSMUsvW2fht704GnA9Wg85kFC4faRIlx4JXUMmK0XXi9577PRj4yZq8GSGWF
hLtuaWJ4EuoVfzUOAEuI7x0AKsXOw9aOMCd2wpY75izbHrrlli6PSiVqT9dB6Nv6fHWsTLs4FNiZ
8RVAHDuelRFo6uZOyXCfjqj5KDHnFwkx82Gje8wWY01Gn54fpDaxLZbX+lhPvmlF1vFHAVdMWAU7
2p//Qc96DBQG27rs161ibsWgZ7HyyH4Pq1XJ6tkR7cWwPNaBQTQxIBmctiQpelaR78Yr80lcUHX+
V93Ftl00Bv9koZkVlxCQ+Gl0asfmOS0dtNCqtETMKgP25Zmn8tSPHyKCR7kesDHhl5wYArflqtjb
cXkQsofEZzxC0tx9CLw9jMFaVaBJhrGwAw0/MA61qE45JVLiV9A9nrGaRQ/bHyceOGeSN9CLn3Yx
tz2ZqG+8M2nHV25xkxmyEHxSaPjJdDiKDs6li4hgSyC7/EsSVGASQzCI8v47Lzz+ZFDvG4POGpqC
sMB2AwJn4hcHVh7VnLAf+QTMOWnE1ZqHcLK2OHhTtn3BiGlmGqS8LUgwCybNuus2fnlvZtXTIiES
Gwoesp1o2ZNYlVYzlr+ECzBRUZdGWiNyNVHMaiWBV01i2nI33+/xWtD9maCljd83bFnLuZb2zSxl
N5mKe0w/RHYpJKvql2QDkpYkPczyJk7pGPI8Hw9/u39nNkuIO/bYQ+DxC8cA3G4zeqdvW0q//ZBO
zVynOqu92ThLGONcNzi2LT5cVlCSK40fLq58T/KZnV3IYQSZCsozyzlk1qJT6k3osJJfwFXoltzx
46yf9FOc1S08xJNBI3eBzh3n05KsxRDtN1BHrWp8QLwgDgjKyDt6GsZ6VJFhepycB0SJ9VvWIOUf
PLVNZSghM6HMZ9BaRoLw0FVd4kAzU+ZUAvgK/+r2LqC8cWQJCoXpqoW2kMez+ZSkZaRAgH0cFEaU
QnPv2J+GwmWnLQzy5RHhwbMOrZYoJ3SEy+mYo5qHEg4ZDqKSSfcwjrg5t25nnb9HS94VFk09JZw6
7/doEMQoeUwwy/dxs7eicUgh8aA8e1arYptgvjHUmxxlEJSyYpO5fvkAJ4tVz8X7hkU+o7sKldbu
dTEeDIeCUmVJCRKQlYCP82EUGNPHRGIETzgM1MnXQ3vmg2unXw2WhgozFARgUuXoiJQYFyMWPo7A
ljIdoBlaYYiScVzK3Rkuf5q64YiQMYQ69ka+wKK0UY3gnlzrPg1oRzwnHXrbW2uIjt5e5pDOzG5w
0oYnbwlSrOdo/NFT6N5pPNIgHw9Bo9J1589XmhmBW4S2ZHsVL3iYzjg0hKfBcLpiiXwxg+IiRwt3
PGTzmsaZVCSx+f8wXKiN8tkWptgPZ44FfB1XZq8t1ByyZMEqWCPCl5K01qfwMt6XatcXj6xsn6X1
2ZZ3tOYgvx98IL+kV0cPdgrzmKCW+o1DJb5QFUDz1fCic1pHEKQpa25CnixCAFmF9WS47GvSTzCt
slhCOD9jzgbwWGLtITnLYDAchv7kHP7+y7Rt6dE0kvv+mwZQW03e23OsKPQx9o//I3Cdomk3pMsW
8hBDxUuW0nN6U8OWOtbWBhYCSZqwGir5B54I16Y36q6GXnHb6fs/GHtVhgg9QU+xVvXqDcfj+VEI
jRR28+7yUaMO9Doeut0luiOR2g9YHrPXhjwEFM7inQtN0EzrTOvum3LV3qx6ZnzdQWP67WIZA0eA
S/p0FuQqz1tqFd9aY9I+g7skmNg/s+Zy3gcGnpZqVkDH3LaLIU/ONyj4F9pmXUe+RiePRe7QL3l9
d1qJ/wfYqSj91+5HPnbBeIIsdN2+BrlIpYB73VgB9p7b8pcBoBKmNrppmJkwxbCv9dqShq7Mc6lc
xStLsV+77zvzxWahbltIf1Dm5YynjJa+3P6Bc+wl9ZHGaaLMeafkq95dMeqkUzffFLcjQBoFsbYl
jmD1e0in2lmNy+BE2Pex5R3hbJlwZ+9Q5Bz+T2XL+HzNj9058RVUNT2n6XcigGcvPbB0wV3HXBuj
lxCQ740wu/Sli3nQvKro57rsdQx/aDE6jv4fSVDMbKhHwbVXAeC6T1PdZT/Hf9qj8Q2JbUOm2LQu
5l5YMr6xeVMsOe+SgQ51YfPbPd9VlDU5wDRM5GQWM8mDNhwpz9lJcZYvEblghgh11Wgp72802Ebq
M2tPiLkp5bnfwWrzmqJhHzoKjaTKNIKQvmeBVnMShKPlVlIj8kSTaizWizBIRXy0AfnstGZWMciX
SqPLOrz6jmq9jBlJrta9+asD/SrKsUrTX8wB2WVZnV7LIVh+9qCPdY/INx8UOT+9L8rgD99a38Tp
YtUAgKO7lonM9nJZsYYqJHG2c827ZXg4bjU6C6o4nYkq3dp4f5/mkY3dSSY8tRMl8p+9nPXL8kFK
I4JPd8z654Flmkmx4TekYMY+jInWwbeqOeJZlT4zkeD/1mtMfaG90j6UYSp0jN9k2snfgl5k32RN
DEIqDUsfgje2gKub9ko/EGs4zptKGeeYu72dDcg44/kQ2QFlDSjIlfrBBf5zm/aSjw4AkLgLmJoY
+0JIj/F+Lh5Ab+WzMBLd3PERVuELEgSRoX4/6gRnM2O8V7DgAiAdf50suzeC1k0pm3iChY6PIYj0
uaO+QTSiX3oVgZuncudi1cWquUaWBkd0sUXLzyMeUxv4ChU1+tRW3dgG3+OkR+vju6SO1IcZFzdz
Vuniw1O2x0xnplCRMHEX6KYXcvZBTZ23GpNLGkakqzhjcikSAYSATtjlKSUtFET9C8FE4Cv75iy0
MpKWTYSoFm4ccKhnUfz1gCYnAuh8kAmlyg6jJjUrJ99w/5BzG+jRFUQjCrKoU8pl+5mvDRdf5u5H
2M7zhEjx6agNsirAi70Ahz9WGtE7knvBdydvQwjhlL90xi//sLIHWszuN3yb3r1IZFK4Ek8+8FUW
QuBKoZnufBJ//JBMeJJBPhdq8JJ2wUyBqNlrPI1nKSAnKkwdiX54oJf9v0WIbZ+ehTattb8Z4KAG
stIQ4Z+R1SgtyOLbqWufk35Pnk33n4gHOwzjQgj08+rHAwdAbmQtvEJ9+zcoBYqcfrh04Q/wnsxM
Jw+Xm+x/LmG75tenM+qBBsYeQ1GGA0N+VNKMI4wEA0IjTLOaq2s2G862hY/+A9FykAGUuftyu9J+
QeDcbmfSUjFQRjEAkPn3orH4wyed0PXvvCYfwecf1xPikKdLiqLm65c8YZ2LDdfwvnaAAsTfYfVY
viYjapF1Qwjp3Znaky17Cq/O81jePYEnWxsPcK2DzTQPJKY0e1MY409MeREv+tHAyQBiGvaUIwdu
HKFObOa9twSIzBi4Me/KPXz9UEmqCXUK/uTrHjuX9BwvDrX8U/jPUrGESu74NwDThsYI4IU/MPE5
ynUel2gjiSvkp+EvcGvt86ZlmggxLIeLApbm12IeHC8V3TMA1F18JPBGedpt+N6Fo8Kbv/5UdXEn
eoUSlfGR9WbmtBWm/dCGvGPtDu0HigZRR7GvT36fhgYSAWBSrox4QUQZjnzYLwIW+L5us/xkyOTA
vbmoFgKvmhKopQBSP8HvLfRHCBs+j7GCyPpnTm+WZ+/9epv/tSo6g/+cz0a2rxSdPQdBWLy47URU
DDTWjXUUIYik93L0qIezGMErtFg6NMtV2l0GHRFsZwFbO/9AXz/N2KD3CAZrUk8S9Een1AJ0vuL6
PUVpSGaeZKHHhRCYxDY61jKeFLF9dGBuMQdJfNORAiF6oMgm4hCM9lJmFDijz+Hs5zwWDDTAvtdJ
mOYW4l4LwJ69f5lTcEDDxI7WtFgpriOz9r8VrctCXDWAqudW0U3Qj5alTJWUfWBHdcculLyXoslg
n+KeqbmUih76ohwYx+ayvzLTccTXJHJ0JjNHnkIHKSnLAI9OPJP8xKxJP6227LYlMZcqOuE+/l+b
z0z6js916Q/FqCZfHdwcVXrl1Ne5Fe7L7/VYnPuINkZ/5ZdZwdtWqrHto+sbbZoYMSEPRg9hfccs
g5FzfmmU1yyi7Dbrz210t4NyKVBdb9CRFPFyHia6USxg+MYfgN30MgNj/tMbpmM6YNl5Ed8049FV
9uyQLVl+Ad4JIHB0MqXQuX+P2K0I8YJNXETZyD/oTlpsdegKVhFHcjJ5k2IJvEjd9EsG/ZR+X0gs
J0GvobMJuOyYdJ5q7NizgEY2lmk9Z8RcmWOsEIXTcpbd9pdgSmADmU3r/6K20qNk/thlN226SJ4D
jL0dtc3mZQqJcMxb2Z0cogF8DLCpK8Ot/sKVB761Cag1TiSRBkJmW1YuhwTCzLtSukX0fHjtil+M
5cIW3adBKkOhUkBuI3+aezAGMVWihup+V5T6oHSSVRwNk1PeCTDZ1EbuOmiFI2fRPUkfCWgriLoz
Qny23ZH8ZqePXrOAehlNNqAbqW+PUvw3uWaDyhUaiZBmLh4dmh+OLzkfrAmFtMMFnY0j4Ml8Ntoa
w8J181An6KmXnYwolZvozBQLk+b1YKdC3KOBWEeOdWCaxHS+ZNgfA92xN7Sx44pPVed2i5cYdIdw
bnhwxgde7iWVCCO6CZyVoSozFTStbLYwwMa85JwT5fFkY722f8Qif6EJM9YjYGUnKeHDA0DgSdJ4
rk5KTraRmjsATcrMK0kDzdDnn+wwyy4hAnwJ1MIs1z62lnQzI6V4Gs8sL8lelnwsJ2005hXVsmS8
y5vI+JEDBtyzz6Zmn/5kGWEa4iMJaSFWt2P5d2ia1L8rhtodlCRmgEv2doxxOCKydoGIpooHj3bh
Gn5g3BoliM1XMiAXI1rYyiPjl93/BZL/VwPi8BsdHcMjOuoPD+khZzFQ+SV87I+96d7/zQAMTX4Y
q+UhriFj1uhPfljS3kx8CKxQCpUAzvWLqzIPn2LnwW9uWQQwytm1YIUTZ3Cnk7kQKIj2Xyvmv/9J
7SJ0mvSodPR4N0Glg4W12zbdHcDr+97Gs+TEibAP5dGNQAsJLm43h4PyFeJvIV/s6Ugc9qmWije8
wEHKonEeMAP9Nr4029dHjE3UfWHCDm35akkF1qhzwtbwyoDkFIBrZYrwDPd4pTN8pzg3SY50Ogrl
WAu3BgVwktcC2hm02PgMm4G5BsTApxECDLDyJdsk+ZuD8iQpvNw2lf/C79JuvLKfip+UCA6BFoZz
E34hrgwilNsAJ9F3P+6OTxRs3K1reRxDUxEr1PCtOGuuQoO3mdYwn31LvKrXYI1KDzGZQL+Zv2wF
329mvmxREaR9NhU/I0N8IpY97ToylSvkFHU+J+Pd8owAkojneNJ8EBEOjMvpw3NQ2D9rWyhEemjz
2aZuQo/kJE4Z1Lui7nDtvC6AdzhQlEFy8nPLEByGTvGexYqAQPYTz1zgcaQnSzk7+e5wT3sIO6/q
NLTwFwahjwCTpC/jKc1jqpcFFtkFW45/ezvCc5jeeve5uofqIJ2JgZgY5iOfeFDTaPDIOv4C2s2U
KhU7UuJsyz95KxkwOC6qjJ9uFMyX95P7ClyMELZMOBz3pNGiUNTv6qNPnRR6E3+XCstG3Mf4nD+9
JQkLRrnVtO4kEfgXSqsG1f8X2unmFMvpBlwuy3C6O+S6ZYGnl+eBpLxLpiQ/P1UeBXtYBsHeFZrT
Arnsef6sqPa1vCgHheg1/fvLoH2yVjC5M11R3iwkwjW0LmYbmlVXJnsWD2gjQt1JnIz3f0EjHx0E
GTtq5NiKgguyOUwbt+MUyqD5NGcyr8Qgm7DEiF/hjx1p7ux+BdsPc4lgSduVyuqFDu8p5iInZAtf
TYaN+/dnqRRV1ooRhyOBESM01XL9ywVE3U+6rBIrBBQkvzjVzhTCHRgyYz7XFiLnan1v9bIVpS9o
Dxu220tktR7sRIVSfkP2iwcUGKXZiolQDMZNukSIL0GbrcYGVLmZvNjTvS8VXf+NCZfl2poUqJQO
dnaD29CjmeDMKqEjkjqmomBmTePCgtbRqEc8nM2wczpP7rOqoiG2MFhYmfxaWmj8Gt2Z/dSZc649
3iCwTbu6Aho29JbkDlo7v5JB5kcix0BHGB6il6bZdaQQHEpIaCjdC04krNdsRcY5ooOFPsRFV/nE
8ySssjrmJl1Ef61OXtluJCnqS328xnCDo33i3IsYlNZq3FBibGZfNhl4esBjXZHVko02Fi2Ffxlm
jQwsB65INxMV5LJnmw2VCR3LUWiHuBskWBN1geyow56VoVrVYKjTPdM86DSiTCtF6uK7hjXHuZ3v
r/4PAh3+xYvmDLYWFhnyAd5602V1oD0BAb4nj/FeQjUOh7HIJUpMpGHlMIfzKB5WnGJaWN25In1V
epjnf6oGtXYrNcRbHkjCl8L6/qTdd7ewaCxYyp0Ze7hNzEwqixLEUb0guo+MwqccmHtQim+BOGF7
WiXlNCXWxtdDphlKymBulG4J12Eilil8bk78DDmPQNWKIL8Z1wrDmhCDyo8kgWl1UGVq9EeS3tCe
A1NRv+aSEr5yDjoa9ebbk/aVZDdE2RFbewcdHkgB4n6dRnghq8KB4PQ3V/5YUXMSbxVraPIetROz
Cq5ljvHV2ci+GCHbOQ95ZpHI+xbvF/Bhx1A0uPffCHV8wNdLDHpbm4PSR5t+atE7KQ7EPkU8bgie
q405ejSykdiwbN7zMMqB/vK4fq29MPVoj+brghmKHI22VQKQhw2HhC3lzUjExOgxk7Vazu6WS9aW
TeS/SLhI4buFLy2X/vqXqrYlMHasnP+NOJvpj2dCWg3OYhA42NML9QPkt1U0Z/W+JZin8xtx3p/w
hrIwoGLOuqNweq/BaINZKvxG2e6Uj/4+4eOEyKLxujTGMTVe6YBe7D2APjQbEWqLArRqMqCU8930
u8+z/Z94k2bKMl3I3ezfLrllQEhLc/owciCHPqw11nKmy4Y0Sab+8ArOBaeYAQE0SVWuSE4OEqxq
nl8uh/Wqkkdy/oCOFRKZkmJUYoDHqIGt1m4V4zEmVottGlNIyed85kxE4+qsRv22uZ5biGxkupqI
i4MjwYoZVvPoRVw1ZL42gz4zPIHs+i94sNiRvODzUL/GRU7qHYBwk4vAbCrvrU3M/PLNSeZgEyH1
nkOIo2H8NPbYGTPEUkeebFLKz+xqc2oYSpC7h6wywpRQ4OVterTJdMen5TqMaVF5zYN1BkPE2a0q
yqbXH+A++fEMfJiLAf7u4htRy3YDMgvZB+P2uXehkol9h1kOzbrarufdgyaNcnOH9VvCI/RZ8UtO
0X9g1aytfyCHVHx9xC06XRJNMdw6LTNH3Upr75V+uEx35hrCtKMSPCU6n14mVorIRfh/rhw2rQYy
hi5Gl3rc+L3BEgPxCXtCbRCCaUlfs+Xot2bVrFOfv2XbrG7c6gGenAnLGPhK2VW/5MZCu/7Wjvo7
P08Z/5DzRcIm0ehTxgCzsrouBg2rpsAlmOpd+urFqRuxT/T+nQiaonwqojnygfussyl1x8R3nUer
uEk/TWcct1nG678f4s2t/KDq46LyLHBW4nVv2Yw5D48WZ8vhtcDAn1c2JPUgjsSpLt5Hjkx/JjOo
xQ5/WETdmFRNErrBJMcTmKrmX0Nw5Xy7osPGa2+qmcQFUGIFrj/XHZbiWRru+ikjfSFf0y7AviNu
EwAArPGJsVur4lTbT+SgWcq6SgWhqlrvPvA+dJp5D8/ahQbaLl5UOAtNr+xySXzjIADiH6t1jILc
8jlKL1FVNYt22DSiv5MrzCogQDk0jrbWUB8QUmeEiJkATrlwbaThU6Eu5j3e/9ao7L3BqgKvYReF
S8UdPjOl49zEofpGgDshdDx8X+pAsocFCAPiqHtqPEk6NUtAmBZVihwwdONNr7oRQ17xBlDbwSGF
7WxjSBEEX1FXA2Vo+JWJlpQTzjypskWSoNgIDlOVhp7Aald9LE/SLTvGy/s/iimUpPxRsg6jyGIf
hm2y+t3XNzngShRdtXnGH8o2bvb/PQielSdoQGZZxI6XFtKCwTCWl/nI4fRuHJYprcOXNzcx8XlU
qCpRRwcOE4eXvISvbeS8KSvZQn8QZxQcbLpS9brXHa8dkkXRMHNrTsogY//veLX3IyLe1G0CnVfT
yjFDJy1v8AKmNSjkzt0XahcXlzo9CtgizgWxfYbh0cyMUnh0AJbs5Rf/yHCB/790vBsCCHd/wfMP
DPAQAPhMT0HxlPoWDjN0Had7K2vkuqyUBLosWqmomH4retTO947jCBewgofQdKjylgIJSzfqDC9l
p0FuZusf+nSNSi1VtwKKBD+q0qlrT9x+AJscAnUYqhnQtmUiT6gC5Br5dz026O1qWRCGaVEvwnqR
XFCDU7WcKZk1HpwWUfvpeWnX1Omx86+DJFpJH2KvICtRngcvSpWc4XHhaYZIDyBbXnkrLQ6G17mM
FwCdDc6AmwJ8XLVAeAMDIgbOYdgk0rciJZaIWMSFAyALklavGCm1fsn92Z+r8VYHkcP6y8oNL+MO
ECPk993amAbDJHFE0CrbrY1nEySxQrfDseqUV7ArjjCXLkiBmOariIF/eCCqyhfOjp4Q1ySUm8xZ
ckxS/2M1b+GByqVDYK4KPYo24y3NBv3KXUJug61NInm5ji/zuZ534RiBa7vOo0J9onAGdMqM5xGa
aq8OvA3lFBxEYaSoC68NZ3nZ3f54LyjaInWzHLf8y+vmHv5EdDWpoYePK0osE72Jl8AChaGkuWWK
KLvDCboK0CYu53tCmRiP14oJH+5SuxbZ2pYlynV6KDj61E1PftgdxTR1Cz7/nzqqrkDOJyHjey54
pxKk9iiOJZgIn/4g9raAmVaOWv8ic7t6x+iSiAmXxY5rImgCOGvt0rY5K2TuwlOk4Z6kTOdRCSXa
GrKJjpYWaoY3AGF6sFz5QoWfTomT44bU9lh8EaWPB/zI5MVlHtX4QMnq1mH4QCZTAzsaQu05weSM
72t4bTRwj7hWsI5WYYGivIUbXGMZf0aNK/B75H9beOZ+bwKC/eVjrjRSYngZmsYfReATYAkhjMIJ
sLoNtDjX4CJ8KqA/+xe/HGi+HqZhIt3LUXyORo00DQ7ky/a8XcBbXFmVZ6P5R9W0E05O+XAU+RTN
NP91B8xYjXCuucWa2LrWgUmu0C5o2pv3QSS23SBf24EgcmVY9c5g7LJYO5H54saKOSGfaDUzvWvk
KeYeIiCdApX3StWjlUpIqfSoqhA/v1ZgnMvzffC6gl5Iz0FlgvVS4mA1EPWlsc1yxHul9ilazni3
D1P246Zjt7jeTzSzbbu2vvA+EzB7Zhc7Z58UppPnBzCCmcPzXuC5UBXLrBzvNCnTVJ1rQNRDbrKE
Xxs5Ri6m+swZt02Unmd7hlJ7MQfdHjI/w7E6j9UQV/OHcy4JOgzaHksQIDojLM/JwcxYHnMf9ULL
2D/GAbVyzt90aAD4UjH2UCWZ71S5DHTW2OytVX238xpZVr/Gh4R3YQV4yECxGh0B3w/8WSqNhtc5
aHne3H3V7pB3bKX2QX2sp6emzCgh3xU1KtXefxyCIEPhr/kQGn7KGPYAWSSJgZ73hsOx/a0gw3dz
/RafiZdACIKf19V4okQFKKA6fEfDCqs77f50fZd0oLSs3fZAmzWI9gNWX07iCA0+X6dP6MsefxsY
BTOINFN8wEjkvUhtLGzOt+g5QhItjoYuc46WQp8gpgYO2Lv27rrZZMN5OvZ4r1pRXxXkn/gYucOa
WSEFtkzk4ptWxtOQBnLW0GbUtb+cskdH9d0nQTYJ5p37xCz74W7/dXPwOimN20tR9pjYc2KpNQga
2NuglUaXOwE4wlBkOQTHNGkyScBSMbO2DTlUdrBeZiSI0NwHojo+cZ2Ry1sIapeDAJwRB/Kkrn6V
AxEad46N4jVTElAjKuqLHPFHjyGEZtJfiA2L3f4tHFrQ8RxR2DtdHW8dIns3cvsex1hZcd3TILc1
/dy8m0fBZATeDEqpxjQqvyMTHnQl4SpFfWV8SXY56kgo++22kabWTgAgXUv2U9Bmh+3TCw24afdy
3EZNirGxy/YfrIjbRoW9DwIIEsdm2dhVjGklrghUMs4ols8G6z/LnHLokJZ7sI9B06tnIKdxRDTa
wtFnPOrhSlI2F40fRbC5rkni4gVqvvo/uJ/ubZ+NOKzvXw/RkinPR8cCMqlAoJxg8wQHXFCUuda8
cjPy9IPp9UiVdqn/dwIZccjX70JH1VieYFFDAu00eajgcL9OoFKjGDP8ErO08o3P7/dwf7qPn/Cz
9WkL0Ro9hiNaxpbmSeZXu3UQDSJEty0/bzjfzX4dVx/CgfR2BV/3SFYOHKgFOyQYDigcQfN061Lx
Ebl/BuqmUL5AfSF/8NMOawtLtX8yJHBxU1OWTQ9nuHGmVKlSptPI4f40VrezNrvtJJ3R3ty4OUIi
XTbGDARaEJBSRMjerdnsjGm3pI+Q3z0o+y3mCwFcXypOY4xqyi0qROyluHb57AN+owya4wqMnExr
CQoCZRgU2Mpd/GlWzcfV8Vo5+UWyRcJS1rbqArPfANE292YLstC17d8CIqXzMzTUY2DBVQ2Vg+PZ
20uXBeJPo0m4b1AedFmpAxOb8SBTrNlkMDLKAOyLStCcVuoGzru6nFlNrnPycFnO6s9o8WGU/wl2
z9uWqUPEpGIQ2axNZJalgnOs2jNV7lZp9lR2OO00CinrBJ8ZvkU9uTC46c4aldMZP2oFiY1TvBcS
E+QxYVq6HZ6ZOu5oyJQMpQRbb85oTh4w/WRIvCO95DHuXhjL2Se3DJ5yjMLkh5wJTXxm+XPB6BM5
1ox+3CB4E8jNYfvriJDixe1MYgeTwdAJ9SQbYG8gjX1W4xRD3t9FzoVvMJOMKdoZQRio/n8wdBEv
Xq+gt8tLE5fOGAUW5JDymwHHCMHfUDv0Zhq+y689HN0LLAwhtGKwkcz8VQwzdZ9VeZf946Cp/B6u
ZDcAVBMJzO+SLV/puirzVqjvlvZv40kP46gP6Bc+Fq3eZieQ0TySgtDVl5OkiOeL4fznqtcEgzHl
q4295syE5pI7GKr35E5vSqwGt4gkBxXpzPiNnpdgSPel931wNw2tf4+Khu9NaQjp6eUYu0tCdgat
pUetq9Hkec7hRkEmEzBEu6FLzmp6I1/ZrFn5zXS0cf6ugwGX+OSWDHXlqMgoNSyvcR5YpsapdWpf
fCAaGVXQUMJfzzluiI9KEz626sRMqConm+lIQzQG+fB5deBBRlH32LsupUBPU0Re9goHpJlgFpkW
kw3naqeC1kuuDOeF6Pgnyw/FImOztc5TScxkTcJspjQqsPThA6vYjq6nbrhJXWKx8oKhjRfpEGf/
U74d5Cd67fLHBr0aNIsyyglIKLSeqf6vl6NhOCt/fY4ZxpsymE5cw7bErakrQRrcZjMXguqQ9sTK
ZCjApA9Y9tfjB55WTly+4MVNycLZqLxnwkUJoLxoCrFb8XbkMUeTd6Gl7NJLHQ5fJbMy+NwydmhJ
OZ4LBkwrNOXVJgYEF7WImnTj7Nn7aRvMZpbKtilViQYzjTDU3ntWwH/QLhQelqJ2/kw3qPIhWZGa
FHo26r8ilc6JZWV0UP2So/Xhgmxqwnf10qKUVk/BA/pjRzkoH+3LQlW4JoHW5svlyX7G6Q7Bt6cs
jaHVfcjtGGe45r9KR/K4Uom+1UZNprp5QANOr2U6BEqUMv85/QzLTdpnj7CwSI7lUzielgtcx0pW
DHTIaiA+PB/KXN96HMo/avMX2a6IU8BwYQItWyjO0JYccQGTFMZQwi+8XI95NIsP3lYxDbuNW/yW
fI2Wk6madjMdsw3A8TZaDWklwgK2MQTPXZ4ug0QqI9Ogo+OzZR8AlA1BKUm1dEaK0yc2D6XNgP8I
Ywd4GraVV9gnaHre7MGCYvnHV2Zn7+Mbh6dU2kAuedOc2eW1wJTbuXExthIHx1GS0ZdruIJXiayO
nJyp7UWzURuS1mp7jbYyTlEUKNSqs/cItFnwmuwRy76wk8nceUKGf41eOqv3dGsso5oRC8NcxHbO
XMxNu6q8XFvyRc5d2Z3eLVNK1E9BUzu8bMXnwBLYRkFcQv4MP/nBhwsNMiw49ZiMuNSGBlroCDWJ
NrZTA68Pa+mKz1Q/kNGQlFb3QKccMUr7WRm6Cn8Uy06pO/biL488SaOJ4qWuDAK/8OnSZP04+wd3
wjp3P6bZMqUHGAybUlsMnQnxQtYnv5LY4dldcZpof1KIdKrqwxXT8T/x2j73y1Wu+bHaWzpOFjb4
Wy9TFH3RrPVKMz6eNDr696YoQ2XFD/npZYE5mJdT2/DInN3Dgstue1GczMp2mfy0UfGnuJUrL1rV
7WA3dMw+48E42xoq4G/+FIltzxVKdSK+RGxxCX9mUJCDt997D54cZ9+2CcXEp4HzPnhBToB/OQri
m4cNZsjL1TnWoBphenwKXIBr2ali02jRM4M586lp87zDSuYkhCloGrmEOFXSSBsqLAlk9ge5GxNo
CqmOOQtQSPnBIFCOi6uKvzgkWqJ2FbBdWy4ZOuDJsdS1t3Ni5pXDIs/u8ngvDAKSppqo880dOWKB
spc98/NHDmQMKgYtThIwa33Y+p2NoSi2jKmkKDLWUwcJzTPyJFwgEo2iZnjEPMLUgk7Ury2cC3sA
a+rE4CkADPoXIpMeGvFQp44buFw38m6mmSqumnRR86cZsvy7bbN7OaGdHlE/GVGXPKvm5/WOP+cf
ZYPKBLkE9AUUf8AtjfJcS7L1zfp0AIADKRNcuODyTWP6PT9Z/kXlLNPgh1S0D/QFo009yVxyiYXV
7J/JtDop/WfXgRkvTKpExJKlPd7cVVuW60Fxm2a9ZkF0tY1yAJXUq2MboWXVi1GCg1dEkxisPjZg
i054guTXQBLzYSeQLHPnODp/Soh60eH0GwOS41dMQhYgoqpWRqpa9Xtp1tSt+ST5Mmjx0Z2Lt7Qn
g8B64pwiKvbGDErPlN/H8TZXzZ8cSQojVdv8CxQM4CDzn8QPbevu9OHUiRr2sKqdT5Rfn09eU1FL
L71hRFkrMgcrqndxAWj6xjRCgRfVd10HU8NB6DxZgR4UM+5W+7EVQG8iEuHF5XjGq+PaSY6E5e00
17+UxYYBh8WY03klvHzbNgdoHqYhF8UU7uhRvoA9hpMlS6t7TAf0YVlNNoC09gMUJmI2otYvGQfm
Tn04P8WWtZE0kudT48/MGjpuHsAXAZ8n3yREnMjLLkdIkizuesDZNQ4S9r2YT1la2Bet/Fha2wnN
I/7xNVP0fTs7ZxWXqI59D5Qfoy/YFyN401CVwYpCWDbhYfDtK4ObE/jHKkh3znOebUaK/YJr8GQz
tHgCbYEhlx2pTq7bUOhW5w75CmZ7Lr7OgaGvYc1HQikIwENmWOpuaQUI2kid0QAeQGc/lHgzvSaF
XZZzrkclbqdFp8ljT/ngufgKs1vbeCK8a5zeO1Jz6/QsELgaQKDxgvfoYrobCBbO8q1FOSv3foPV
LVrLwtldLVbKoCGv6IeYcfFSmy7f/qAc9Asl9AxI6ryipeHURsa0avl+sH87zgMNf+50N7iQRDUv
41HQuFP3K1ZVbEOptlyFQHbOkrkz2pgCLj80qc+EDLMc5m3UAs1hyfZhKEpn/J3OHv4Vi9+uCgUF
KswtnjLYz1fttNPg4RlxWHeYZYxOEvipgB1VRw2EJipJ8CgdgYg6n+2Ix7Fpv8BHX9Tkw7XLq3+A
Zwqb2ue0itS2vs3XapEiuFQjBa4YOLj74Zaw3Z7ZzL/NRbr7xlZ/S2pncenSxX1siBfklZT7In8w
s3g0lrv/njPPDRu/39/rPO48TRXrT4hWWhKnC9mE6T2/QD/x3iuZCmcgKvjZusUo3j61h1TedyO7
Qhltb8IBHe1+TmR19tzUEHnHuFPgr1zlwAGJfGo43O30QSqjTG24k9AWdfBwXOt00/ufZBmj2Y8T
jAM6Zy5QpafScRnsagRkFPg8BVWk6m+vCGZF9bi+ObVGeXmw8NDgdVceUgwQzEvJEB2BOEvID27W
F2SotZ2YEbY4ijULSkIS2GQREK4k+bAeBd5dICu40Bodo11BBOgkr6DWM+NGlxUkDxHkJJKxRbth
exoZyAfLXWIJZWFKKINepmbRrUIrIv7evry8u8ZXbOtAgBmA6jrVz1GR+Z4b11d6MoY1lTmt1p5S
eLFgm7wy+Qg6eGM/F14OUqr/Y8NX2nFQYMCQ74OP5nimsDMpXvhghLfgoK4ySVIwxy+DpKwGlx6j
PduzJNAOFklCFiLEbC2BWEyZOYKmkNfS9ZgNv1fW7KCvo5rKorGh4ovsVk7zjj+812qXI2RFoTKF
ovAyPivOPVgFps4rALWObdpVLuAdAv8O16p9UqUylLOv3dChzS+iFJE0hQb+XRPdWFspCKfq1nU0
ZvJrBAsUOZo8U2TSL4b3t1uofAWMzF6OotNPJAq2R66w4i+s/0RV20w5saGq9fd9ejztxDeswhhs
+XA1xP+OCZZjg8XEtS+3uc78O/HQFxXTJdQmNa/BC9S04sOcgebA7HMm1FYnG5BVJ6p6WQ1GYkoj
0NPx3ldrUFTND9+kIkMb4FpXJJtyXy1R8bnbcTHRUKo7wyNojk9b4EImi6bDoa1pfSTvrploXjwG
E2tjxxM84evpWhoslSiq7qXC0CFa85Dy9ntfTQCKDA0r+67ZgpeOLV6BgVC06le+vb2xZwSRcDqr
6NohSxtL20O3kUEH15OekJpLgtrxmtcSWQibq9O4zU7Yd8LY1j0hN3nCYIGP1Fn4xJF8nm92RULt
JoXVZcGQAPP/2NHxKKhyQr9PwVTisC49BtHZTmq12CzX+cM+BJz1ROEJk2RdZmzoJKKAxRYzuwS+
ZU3jvKowONa+Dz/AT2K5ysISdv0u+swQRx0hcqOArbIIasXzUmH7Slle4gJg+87imWfzY+R3rGMU
BH2gZ+9ut8ODveb6ilkVExpnAfjtTPg76cePuiKBd4Dh1WcVvrLZKSalT1jUao/Q/mA6hTR+eCHy
FfL3U8hni3YRq0zB8tDbbh54IKagtEbIC3of98LJgruqzRO6eh0I9HjamDceMIUyxAxwM05wiRkC
MuvrS6x48DfL03oS6EX2etQPAM4tcADc/JRNyUm58ktNJ49hDswF2no77Ymq+UGAuLPUDfEht5kN
ORIMGrUeZceQT3fjeBPyk2eQ8FKsWPCvvHNGk0b1iVvI4iHBud+/7/rwcIA7qaqVpyFcN2/rkCTS
dn1aoEBCUVUfMpp3S+oRsdRwV5+lkwEf/N9dWWsyucct0DZAOtuW4Du9XYobXLsUIFRI4w5nFokh
Kdfs1HL1qs/hslA65wMKkG99OMfy6x4umgT0A1EBT3FlYAUOfwdK9OX/DalQGUxoFmJm2OPSrCdT
qodY0/33TCdQU3B1r7K+hM3xUusHFPej8cLaL6ks2FD2tYuR8WN+PHJrxOMQOOdu8TrCQMuT28Lo
sxzM0GfiOjx7Ew4J/HkYRVe86WbKcBQSBTOWQQMgccxIHsrwQWqvyEdtwXvCi5VydfS5M1Wgg2Ac
GvfbKWuOczBwo8+/IfIbyZhnXWeA1Kk8JfxRjaYRmnX3n7ENJo30Qt3KTWACVi1T3AT2lTJtH+tM
QwoPSQ3p9lOJfs5jkEr/jUgWVCw1i3Q3WL0FENFA/DhVr+2fe+VeIO+Yum58KGFPdbDKSfGolu2V
VHipfefYcQGnwGcjo0SSFtEtyq9s3woFfrZEhhE+m3x+EsH5r3AMxAQM4oKrDyGVmD73R7VrH7qA
hDxZ/DQueH/20xSicMUSvEjZqKyU+CWQu2/A+yVxkbiP0jEW9oygy21ZXrkC83rUvNUysCEyoopg
uwFBasTwlRApriTbpD+6UEIVigCEfmc+68XQ+Du5O+g0d2ORSB3FgOBkMUZvVtTpGxqeHuVD4OnM
keLXWXQooNUzOmrvhBhMxn4Qn5n1yy+N0aWIAStvUDiaav7pPephSwnoBUhcTbagVIP3Gw/08D9E
FnyOlZ1h1vvz6JjXjzjNeCx36P1PD7qZXBZNuexvTH8kpmQLkxyixsWGx0nW+eC8P7v4O4s4neiy
J2nNj+/y6SBfLHTgIEvpbkMXfhTA65hfO7ADT05foqnuKWc2hA12vsk4jNAxj3+LzhRR63rkSOY3
OUmmFSpwbk7jMszcDpgErGRqXT1PKQ/X0ehSaO1Cl0cyMoOveMCChW018fSWGTjk8Nmv8UOyLJZp
dfTM6mZODpeH6kM1zsF0/oWl2QP9CiIOj8QeAEltXMhh25qaw5S5OjFiEUtLga2K1FYF2UpE85mA
KHpAmUSjMiwnrZnbqONchNTAS34gWCD3zOaMMAPhlbNTIP0KV//Xkk8nq4iYrFspn43AkaVvIw2i
2UWgajhrUJ0Y5sFNtYgxR4Ol9A9rPUUutscWjBVrZjG/+ZEJ4ZMPc/r6dYB5lP2H8u7+Gib+JvEO
1M8oE+eBAn+sbqh8Hd/4OcLqiRW8cpvQu0uGLkWUxB4A/5+M6z94tQe6nHQifnJU/Xr65YxLHPX5
mE+U7ufHO7pXgDQwZ7K2LiIn7uWc/RrS6xav0Qylr6KGvJhIyJtq1YSFGDybP55gjqH6J6WDmf8k
FA6rjTINGhrYfXHUAb44UFvda4E+gRl+owZfKBFcQA0bXqO7Ie3M99ucQSR0U8EJDbfi/XA52kmx
eotyAIYwtv6kM+xRyA9+1WGMJuQlgA+zYn476WWedqfqFM9J8FejTqOdqAztaDryupu9Tl3fWogV
vTiImxEMSFgitSpP2S8/ai5LsQ2eL4JfWGPz097Qa/BCQU9Kf6iYiRr6IWJwfaTwd1ulLqSOmH3T
tK/sZzLOLlmuzGG+YCM9zzEm8zWupb3iu3Ud+T2vDR5xZJdkofhzRbPW1g3DoWl5g9x+lh1zaJNY
szLpDzs4hrAd+/cF64yyTuC1Z+31FU2zG3nEG2fDlKIWQULAG/Wsy3dZ8bY1By7hDO1YBv2GW1a4
gcIJJB/sD+7gUqZ7TD26vZ74USTsaspgfFDn2szT6kGhPFosMfK5+5B2WIo7OePuwfQb4HeCPQcJ
OHQ8hKow4cc1Jq/2FPXnYxfqJX7L5cfyZkWCbAiS542qzAhh2Ttz6hh7wkCHfCA1lOgp/LkeCl3A
mtK6G8h+Z3Z0hxhu9AwPJkMzarCkwln/BA6mzyAsUmH98daALcAmFgfYCF3JKjesB1klM7ec18ND
L2eRCXdT/v3xog/kLmhlIeAR19nih1bKLeXc6Ly+7Q25TXdLpNzoo1oJ9tX1bf9GYw5PipVZ/i2Y
HDvNicMS7QSX5rwGFFuP3Xg4rvTi9ee6enfuCvc5lXG9TsTfcQZi6u07dbWu6UKTsHcH8OFAvQkS
Xhr4mfZmi9XFLjmqGl6eRvmcG65TR28nbQTnYBwXYMvF8c/f+/0mh1Z9+Zxi/xxtjWqQ8tlCcSy6
BIp8gU3f4ATaOzIXXrKdisFbaylZmqDPyfbDMCoPRkqSEW/gPXsuDcAk30RE3WFFQJ6u4UsbBcX7
13Tp5cP+orJiqf6mAQCcAaBBaFw7dW6qP99wIwDX+2KwvDKPrE0MTRT2fj4m1A+G1a2q/EiN39QM
1Zqm7oR1tBpLrSVDoOrbarJc1XQGlspYddfmZ/NllIMmlsVXABP4Qm0ZiM//P8xgPYCue/nyQ+mc
rmfdDRplNsp+RSSImghmeuLeCU76oBVgtrPkSeu0mOAiSkmRuwiSzZnIsN6zfRM+q96RtddX5CDn
U16ICQeZC4sYI1xdY6a1eUsHlYqPLUOzrGRXxHYyYsGEJ6Ynfb43fbCr8mVV9921lMjEBeQslJq9
53h+Ygz8W1/YXzF+sNhY6qvICPaxfgnq1mCgT8LJhLQIQ35fxQu0CUJxlDoymcTsAlXEp3LUPx6n
GxppBQMcyYfoiRp6+KN/T0XbNTc8nGSOEEQ1BDPb13G/Ub2eqtIMC+34NsMLntJ15QgJSNy9kAPL
89KxSouM8AxvEe4et5bg519P86wSjDq+WXzcYyxZgMX/aOPBqZEPc3NfEGEt1e6spcZDn25uGTEZ
typM5BAzZZQtirjsMkXhcOaEWESwAbK5SQPc/+++ZgDTdVpNehRhAf9zq/LqyPAtzG3hMIiLheuH
soRd5tXF4bJHPYjPGbE0dlLsf+PXD5N2zQYYBXQaD+HDbU5cPoCptbVZimt4HTb4w6KPXv14KAT7
5HpVmwOOCYdGbyEykhC1ripKuE1gRFhdeq8Qrdms+MkfeKI5lOVxnH9B04IBcapYmkeumZcdEOoC
m6Ge/ZFqJ2zo4su3bTwhwsfNq66g51ZBLJvzZPeyOqzbmTLutuB4OD8E9JkCQr3S3iMhFcYv3yIv
U2IWCdbTITwC2D27d1TC85LCM4v0tPQD22PehF1uGDDof+znlUaF5uJuBJLiqr3s4Zt5YctLNMpi
N5xRjUmF+DxTY/06ZtQgAmcHyn8bulbAtlEnSSYq/s+FDUUTOTvJfD7wCfzSJf/71vnpSamJEYjA
RWT09F0HpwHEW7mz0S9xGhzvElmywO7bfLfRUdh/bOpy86+buc1LIK8SpxUh8t99xyNVZM2PmXoe
qOOGMOfPp6YbaEMbXIL9FUnEGlYrtM6v/F9jZBe0ZYkLZWXPhYITig7kYe+0xU/ZUwyWC+hQG/MB
oXs+3GcYrHkDb6lx54QdUWyqeVWcm7ouTnGTBY67EAzu0xAigC3syH11WawLKieZ8jbPoTVZxTtC
PDjvz8VC+7iwEqvTSJ4/xlWmM72fldcyslqUqJaCCef/+IBZO/hkmzCWzvKsWsDyOroyn5ctWF/N
eD2msqw0MLgp379JJhoD0iPHwKdZKNux4H/7wrvDKL7LyH3CCECF9GRqM7icT123M/f7C1smI7YP
jJBbhGKwtbg907XKLm5GmO8Tds6UQrcT8P0+RDplFsX3eJFJPf3EF7rHCZYjd0wvm8Fc81Un+iwS
jwi+OevQa49wel11v8Bnv7u+M2yNJy9Fzvcn1sJYvKKy+bFzcjc9f8Pmqdcj+QqaRW/Fk+8sI/l1
V7oL7fTZ/N256+QWh8RGELfac5H/efFi7Sr4/PwFvGNC+g57inETFIk9DBdgquSClqq2YVxClSeU
ZopMEDgJXIgA3ShlFb9KHg1txzL9jN/Hq4FpDMSFmYxZRj0sUbAfxxKtZOCLyrLM6cG7miXiqbo8
wrpwV05E9wQ3OHoWHtWE+NT4tZZ8IPV+yfSz22eCFPI7NERvO4C5zjnBR/wGAZoQk0VwI6O4ZfPd
+lsc2z9r5cwSPNCtQIRVGMGBHQ1IRy3Za82eFYUepG0g4WizhvLR/fhL5T0O6MKdrdk4ldHwgNWm
c8e7NgntxSquUN8Mwic+5Jn7peOgfGgtJ8ISimkmj5gH3vCjbRTkMUdGEaWzZatZh1kk8iD1mniR
T+U/ZoJ6GbfZ5ijExQ79JvTZdQTteghUvBkGrJtcavh8/Tn7nl0TMFpQkY+4eIdawHDC7uw71MxX
sZmHTzx3WmJj9x2rvQ34BpLaJ1JvxrkIuVLTtqIIJrZ4pypZg6Hcdq6vfSeoWchScg2+49tlJblE
4L9slwb5Od5vXW1eph0hi1hwSPVM0dzV+s8/1xC68QHDROMF0+i6IhJuWLPWbmv+Z+MVrJ5huz95
QTQ81R/oBHOinD66LzA8DTmcciYHRkLgscULOqDdQiwtDvz4ZGaxhcsYax4zk7p+V0imgByrI2LG
AAvaxr927YlwYrL2fiUI3dSzRofcen5E5L41D9vcTg09b+/nxF5EONfCZ71BysbFtJVOygnZ3uNG
9USzBqBUI+Arch1qap1xdGRYo+3jpnXNiyG9fCreHkPAD/3RWjUppKLxCK9Nz19Ej4FxkCTWbK+N
FEIGiYIbSbGOgL3B3XYJZ6r2HbogUexpC7+Bi6GMkk+S1G2mS0rEJHeEZsafuml7yirLrR+6lcnz
DaZgU5Rzq1izgZ5SpKEkSWxrTXEu3kANlPk+WIImbFLdkiJejzGsB1/oZBm0pJi+SrWWC+BrLnb9
oEWoVdh1hLisaUi2j0Rqn9heFvSmi76JAfe0fp5XRxFrJkykLeFO8zwWmPZ61o5htTHZzqHOUvEw
Hay/ozUrR58JrQcUG9k6JJ+dTZ7YepqJCFhSF8ba+0iIguZk9fvujak1N+BRhXXLiEBhsYc0PEGe
pEhCk1+l4L7PcwfrHSU0IuK+50L4jcWa46CnLDoZMSldtx244WJ7wuFPZkcueXeRZnaOhZOtc0Y6
cmzIwpN+8/aQCc86wHarjAyRy9X72u79FBKId9d5CASijSPNp4ubyk08i2GJSMLz+hJmhHsWz0Pt
nvsaiDb9BBVHTdaxx5fesL6TY3va9gFUdBCNatwGIri0BnkknDTi5zxDtEIvZYN7qIruJ7Xk32kd
8DwPQfCvlPA9LQkeEPICahdhqkZEXU4xAM9o0Fu/te/nEdVkOhYmjw9wrYUDaZ93z4Lu6D+dOuXo
S+PuwUlPllptnuoblmmbtV5K4uIm8b/QIsVsRDRX8X4sAI4PMpw/0dwJpQAFJyZt28Ho+JJB92oJ
yloLlJHcfhAXE5aIG9n4sf51szWdNd2KbAU9PFncngEF42m4yHzZFEWjQtSJEZ/wBt4XXPqPUMsh
XHPafzvRZJZ+weWbzv2P0XbDooalbtpnHQDmhCZxVsuHDD2fgz6tyIQXxdQ7k+sPWEy3n/j8gCPG
/Z+HBWCQ/5asCwct4FcQC1YM2OfzPwsWCWr3QZ/5TRVSlkoasRoHQBUvUoQs3JE4sKSBArtRezXS
/uLXCapeqIIUB1BfRlxnflOU5gH386RT4WBM6oV2dk+2kz4uIYQwZDS6zvOq/L2ab34ZYWKqTJHl
QcOyZGOxOH4OQcZUosO/Gx1NT5VEoPJJ5z2Pm2dJbH+3EaA5xbbIaHSxS1ZuH9LSQjR8YY4wdBpN
mbhX3hKxZg1fgvGHeUpXuDstN0AmhK3k+QO6htF4f2lc3qlKqwFzQz3e+D8Zh5mS7V/3q4jTORRJ
kiAeA/caW+V1uUZPEL1IeQbhqNcr8UQIEbgfT2qobwY6pyM+6q9PsR4fARJWAw+VLoFKXK1NXHNY
ycQmUpL0lcs5RKCmJ0StAXbmV7saowxKyjDfB06WIavxcY2SAbvv8Kvt1uEuDoeZrpMLqidKMIhT
btKAHruJkb7F027OZ1gRKp/Han6P5Wg3DPZ3Ck5cQppW4/ZiJWl9vBDWbg37wHwr6kFu6O11J/M2
fUu32HN3wm/730HH64h+ht/Jw0s6p9OvgUFbPTrdcGpx94cc2BC/3jGGElpc5XVjrK//tQoCJ70r
ZTbngp7XfKb80Fk96KwI9oOgQbDa0pY7babpW3lHe+HKXJL/doEjNqggag5Us1xiHn9iVzppmVo2
HatiGIkIHHWRDYrUrYPaA56ABsHciQCMstVMDlTvBBTCkdu2aeOqhZyjoKfMobg1bnAl1qY+8ep6
kWk1RIjd4/IdFFtRgd0ozCM6pU3C1jrsSV5R5AjhNzPfjnP0u75/3SmvWckYt1tkDv5CZGcjfCwh
7QBJpcVmrDmM1vit3SlVegdoM6wDVh+yr/BDevm+YP0apxlbxoYfSfoF+t6c8uMUKOCXuGPFQwJb
jEm6NdL5WqJuEhncdL+r+MPoAjoXzHf6iLb+Hpjm3XZOIND+XNMAizWA1VSrn/GJSeUWcEEqqcrV
WHXNQo1Dihp+1rI+WeH3gfIgQiVcdKElui0bWiVWNYMeLsJCeFdlIA5Mq0mCXwFa/0Su0YCXAe5T
iH1VNgYDIcaOTkrUk43U9ElM9SQ+TLB6xN4R4ZlnOQRtX3OezfSWf34tJ3zMMh9mXGdJvZIaIyIj
rwkaJoinuwHkdtF1787baEYUczoAgZflAlQPZNHRHP7Jx3caXSWxf40RXHK0OZ21Wz5gq/t8+j0R
PIIxNVIbyByZ7Tn1ZPUbV0AzQLD8xw0A2Bg34cI4DYJKmOOAzVDQA/vYh2aeYrSz35c2eFzBUC/n
ObnGDdZCgu3q0NEzC4dTqIpvvclYkffsrb/rtTgRfamjo2WPeXtvwXRg8N/B48VMz/CTLCT+Yl4g
a7e0ek6kEZuinNIAKBhEJtLoM/AJN1shZS3YF+JYqzUcEfWaOCw/d4skIb394+mW0ZwcTsJnZLjp
WUzPGPrgnKalvYmnLZ7khwzEeV+KtyK/k6DJ5yQ0XbpgQMux0lzcSIJ3+PCCs4sGFyEFArCTok+9
GoMZ2cz/L67S/etAs47tcni9zTmiRilFOfw7+KmTT5K/E+95gjMSm2jOe/v3OuQZP64iubDcogKR
xivy3nbO0KSvYqG7VgkQytZqKDwQjKFm0fnEYmOcByG/oZg9rzT1N+wL1V8IRgszaTW0P8v9p7GV
9VlFzI1OiLMVh5hl7SSnx7+HUuzOOf/MTO2OVAYR9NlDAnDNYNRYnHO74wH9UqH2HUAxXBMWMF1P
OTz4hvXL8h4Q5Fb4Oky1YCXZ1nRaUk0uvfUsP5x2qCn29ONFrpC+bDsDwqaorAfCe68n4odmnQpl
Bx4vd/sVbyZfiyjfq2ksZEyt9Y3HntXzDYfBWh8m9BQ7qVNo0zwEYIyfSAWlE6bN53hF11qsdgZ7
izQHDH0awBb1H3uEwbxnP/DIKHAw3tCQOpuVjz9QYMAcxaRIGSewde/PC9QvdgN54IW4GBMWwLKh
JuYWR9PwCKwGaFHx55dEDrj9+X1xHPREr3v8k9Z6ul4XqOwHHmRggomeYRte56JpFydTJBplpVU5
RnQj/EnjtbkLb0MU/xGdvFN4ILm/VOvCHnWN9XYZ/qJxCrkVoWWNSkY2Hc+KbkweerLQE3R2z+n3
yY0qaFOtYaVwAb6k2mxe0f1ALjHzlVDIw1wJvakFxKVuGB6tTYafI5yGOyBdXmE6BQ/RUIp4cqRR
0V5Qf7zKFKI4LWHH7XTl4qUwksQDlwDiOeU/jGJw+eGBBhBTQzw401ln6nNGKaSrbJ8czUdaejZQ
X0xyLPvYUbp2++pQ6ALK17Hpw7LMNjg//jrnxE3tpmbqFOErrZlQMnIKg4daR1k5uipuB4g+YUxM
MWP+qn4DJmADiprRfu9/4Fw/4rVlTi/CISopD2Wu6FbS4hkDSbrKYwNuRAmdID3RifpusADbYSyG
xL82G0sd5xcDNdOH4CbxJ3T9kZ1s1r8L1wmYERAb/ZWPJFAm0Y5v5xlWdTmqDqUk+eceQkYYG2gx
sC5wpm3YMAZqwsMi3jHxBaAO4eJTYWoO+LsbzWt2s5M429hn/eL03hKBrtzj4YSNqCytnW8k7HgF
U71fpih5LUpqYoRkMTc8OBP4EZDy0KJFNboMfWPeEUZgxRidjhp+8l+TK8TIqNnwPvQbvF8TWWX7
G1OzrTU1nwr6+Acp2EZKFIJlbAK1wIaYZG+gdwZKGYuC4Bm/EAOTiJXD+nF/PgECvoAhXjxmwrV4
cMnjqs0y+HVzRZQtckN7SZ+h1p48o4MDlbhAuW8wv25YFb0wXxKgny76ZJCYU71Zu+bC1uOlhWf/
KiMRi/M4YNnXzdMuevxJ1D5sFkoSBNN2/R4k61Wd93X+un2irr+efxYKXDwZw0zG+8RI9Tia8T5J
QXzYJwQMdcMJoEIS55BraDSyIjRI7QunPpKq+lSbFlkXkFqCfhZ22Pp57H+9BB3r2zsojlZyw573
PwoyBsI6T0fmiSU2qmCKt2mKVEiYSHaNvzGMti06ya9N6YNbBLCCrWyvkvcIkLdcmGSuVCvcnHLW
HKHuph/bVY/spN8zx0cz40rEAN7DsndoeuzeNIQf+S1Gd3/brRHWE0ByBYGBo/I94LwpTFPDYZoj
RjDd+HaM69njTTAOyA2Ca35CPKrP/R3YwmyrMF5+InXgLr/UNrdSh4ZH/KTeMGtlLrrGcDGVf+6Z
VVLabKN9aXvgVvX18vA8b1i1v++VB4cCGWPL+dTGfx/BWkT71tL0m1vZIL5YFUMSv81yhnc1bPEt
lsrWESpX9wWnebdhfJzXvy0nMXh4/9RS9YZU47dDJ4ycfBI3k0DNJjLqYoU3Bwi3oupxJi09rnvY
Tl/44/C56TTZ2Kq8SSviOJf2RbVnyOzOxCmdfrHALi2C1+ScJi1yLRhjlzfAsW6BNrH5R7+wZgMY
Rslx7tUsjBBu7cMUVaqV50hhcpUD8OINFEsMadJcslXa/u0bKNSspefEQbiB4u6gKOUDFqjcrTy6
fvkgjY9irUXU3bwjho4iyU24fL1anUhjEsV2VKpiicU2sjdj5YwNDMPAcXDXHfNg8zt9vvqlPYna
I4yBH0CyIS9FqbS8YjD2wr7RAE7NT3g1UQ5cKoXue5NkDhBYzWU3YL7ilAdh4Zec7yESWJN1I/TU
dkZnwqYyFnRALPso45p3Lwartes89wVflE7PaC/dcwwpfJZ3O3/cT6b0v1PMxLaY4j6U53pgSbOW
7Lkdwc6xDrYwWPmX8ieFT//jMoEgeDIgv26m7XV451zVHtKroqqggzaR8etGxtjhJKVH4mDvYPlk
UcP4+WHQnGRLQgyi3o5PSTLgO964hhU3XX5S/qEwwEu8u9o1Z96cBEDwCMM93jUhm/4+w1q8oAwx
8qph30rRNjaItmz8CFJiAWZ8ArCIRlGpAgFd313VLZ5eABQXwuhZ2sYWLLKavszn2KFIej8JUWaR
54LBxpb/Gxd26DVcKwPMnjEaIsBUH/giJlI8ubM09YDcM9cEtpQbPHBxAVVj9TiO7XGJgqUgYo32
IXb0rhSeyIGQ9qIg7jVCOQXjgNn1hmjow0MHABkKd8mzVsT2zEemVYy+8x1bf5XE0u6rJavLE6vb
r0IiVmrqbkJcic1qUOXNAgJ3mBK7NAqRm2vJMkqSCSZKH1Hl+n0rFP6Ls4LGk0QAz80rK71M2Itf
FtV67ezG+aCEhq0p52Qxnjxes5IKLT6/9ePV8ydLkNBaN9UySNayoJXIxdNMyRNRAv1imV21LxrJ
Jd8IfUYCSZeGFAX8/rlno5cgpKapSc9NkLZncw5Q6jv52Pd9YD+UX0hxBOEeMZzO3IlLNObUDDv9
5d16h2tdtsGjUuj8SXeLPZdMnjmAbHAxC9Mt/ai0KlO0g4gKqUXZrf2yujfqIU7Vc05ycEGtQNl5
b+GdROOJTIlGKJhAI7+5jbYElBU9YVigD5F2Z3oem6h2FvqEDua4XeFGI+EfrBSUSd/yFNEPNS/z
p7u19E8Rr10FhjjjKFMSo5oCh6lTFDYGv/Mz5VCqZgH0DMzmLptpwmtzpNAbJE39RxHIV6/kLtlE
IzODUzyns7UA5M5yLo4NiXjOtLngW+kvUJHbYrUyDxD1fAbks3vN1r0bI1KNyYJEDCDV7d1whTyU
t8GRlPIegtnUdmWQpT5b6IrvB9GGYLQmplif/vkP44KwfQfgZFGKZir9R9/n4c8iTaAOdglUUt6C
yrGuSuReX8skkR19//a68t9e9Dvog2E52DcKKtgbWmwLMx3sYcq7WEHABQrhKroiD8lCwZOlWMRy
e9rYM+A0+cDAvZU+ZiwqhAGwJPBd1UfE6jGL6Uwt42AuB7IYSDH92bmkWCMERt9Wrcsq9oiJO/IJ
lpVRiaXYN0wdgnLraAv3RbmaZ5WCE/UzJlr4u/PC1Zhjado0+Y963vypWYC7cnXtqQjZoPA/N8nq
7Qxd7Dy7MZfs4sz6n6cQ2f2dq3WHsYl6vgGzx/M4vlA0n+plwzgYi8vqP12LIsZDf3lHyaB8YnC7
XIOCQ3tO5bVejNrXQ2q8uwn012PtkE3aMrVcqCWrIULIrfFOm44r9iKUOy8htwZ4F9EYBOtPSWE8
c3XLp7YCqNsCsRdXdSeoLUF2Gg3PfUrnk9eAhXfZYJoSSxxK1QDHPzTDs5nYmuH/+eVuJ/L29jIA
msunsUG/9CH4gXhza4v8/f2ox8sdyvVhWvhOi7PF+ilZLp+ajtZyWPMndW+08w92QURmvdAxEGj5
6h2UWkVi5YrPdeziGPIdcWbSdpf2Yym8HsSjnw9f9jmrMJOXPdj4EbpOi3heIueKRewDzxJf+oHC
hgXm83bNpIm0Wj4Gyp9doJ/NC5A5LCK+vIbsdGtlMILXTmZ9YS4hP3Zr4G/Ksw4LN22GvcgCq9Ed
9g8DisyepGCtIm/rGzKctyW6V/0AdhpoOHVtHsnnOmJAeVNEi7C+lIn0CY0Jg/sQmJ25ZHxgQyGp
WNVfdme+pXQ7RGTmSAX1lClDRpcO+fy/QAeDfcJDxZrWygd3VRqbaEYVxMd54Bt8xt4KsTOzB6qf
klSh7Lya2J9SvwU1fRinPIm2rkD5T1g2v3Ise5dlEoUQdu+QC0HAx5gN319eWT/02r0JuRRpKPAn
CXYyYVulEgP9n2FzNhI9cYrmhMAAeNAEpLA+dvR8+aPjd7iJFvysNwdQWa4720z05mAbVgWLsID7
hc2wzm3Vwbdfx6kPm8C7Mj76B5l7v6zlTXeefRn57eQtIZaWLMyamWtWzzShIJYLp97SG0KSMb+J
tEblY2MPtuIpYfRmNjwSSKG5D8/h6OFupWqf/jvjuPlebah1XfwfeKH3ZMu+XHXdNjKE2092vh6F
ggE/nckwM6i/iFnytfp25e7HtLDftx/WAklte61eghsrWTpA2eSmjzQ9N7SDB55t1F+dROVu1g86
lovAoA3I+IiUJXVCEPFwthC60HuldB1LYYu3fZS2+Mf0U1qQPsU3SPsTt6sI3d3ZCnySDh43W0AS
kG6CNAZ6oYU2+ULp/YEMtAN7/dvGYt4iWkC+Q1dJxpMs12i/GBXTdKCfbcgVxI+GAw+DgaxvMcmw
3tI6oNRkKefNDy0a22nfzG0gANKoOdtA7pEmc9vdytRToXkDKFlinHzxyA1vwioK+SzTUdrFgX/A
KavH5AfYFudUrve20wZewl/ZSNmNTntKCjLElVrnhBm5k+e1Kw3nRy0XvtOt+LBOZxTdTx6qGrP2
znY88JoT6TfH8HiE42kXT/nUGV3/GfpZ5rEIJ11JJzXVnuK3x4nZChk2LVwEk3Npr5FiULT5Uii8
P12Sfx4r9qD8Fzi3hUzOB29dpIS6KK6JFx1imJoVuTnJlrWXi6oU61r0TGJBOrdcjmLRBctNBLIp
rWxfg3XCHgS7+m/krIcHI7n6mkFQYIqJTuqHVf8lAptZ5N9b+LP1CyyE1djfc5GxV/8I5IQTviY7
ALl/CAt+yNNLx57LhJ84TlVBf2jcs1ZJNqCRqHepY9a8ULg444FR4vberlNQjhlDUdTYgY8aLUtH
uLoRxFgh9aXYuAifaxKfGttxAh9vHRVqDiqmTeLV1raTLjpwIgT8yEyK/CRdkE7h2uU5v/t9Ft6/
TAsd500v21zlgQpY2tz85ItfnBp48ICTzjJIPLOz1Fa3+nWGlMUYkDNufeQC3U7FRloahk1hL3vS
U2uE32U6idkq7BZYHGCoEXlKMac37Fwp9J5XWmGsLF1Ip0HcCnxcGAEqUHJ7IqNecEvWcyRU5SAd
Q6KR2ALIorEdDed6ieiWkMPUlxYbdCZH9M7zNjhok8W14zEBzjd54M8na4xjJU7+QixyYBrG37Ek
GgRiWg1QBs8VZvjYDZDVMWRo2qffaVaYbaWEhYryJsSrE037QaWuiheVKmL40RC+H0IHMOhVVim9
BWOoMlFA0wPqS/5XQiAON15Ld/t2/5BEV+dGdgGdngrG6KIOKh/EEZbfbyRomVxYPJP5GewO/1tB
z0Y6oWpkO9IBugZBp3i4O4ZKy1sEFlTYAPN8Dhv50Y+Dp3UpbJ4mvc7RAdIjEsr2jpCtPea4vmD7
w8SMDzbUgLwNvwkXX7DLS4oCkMxpqhWiagcw89b19c/PBfXEpefbbCIbOQqkWbYFZLIT88BuGX8O
dQ+lsRfcEbl1MqIT7zzAHl31THMZtMIU5zp8OmJy5KyVrHnUvzhco9paaMdZMFG2qmjvOfHfxstL
E25LX9r6VAd6XQxoIfovMgI013VhYHcY3zbCGY667tbCO0Dh7P8fDT91nAncO6IVySJlybWLy9St
KVTArthg0wtDQ7IbmF72xn5XNH9dXrmJtQI4PzlLIeRIyICNV+hIxSjoxuKUiyLO0YsnNjWNghPZ
DTtnVSf9bw+k2ZLb9W2Tn1hihgVrp3iPOrM1M5j30f3qFr4RHLFmgTPbqq1lGGAnwckt2YuijRZY
s5x6ZDLBWyFoAFXXwke+iOmRErfY2guh/sFCPsM+LjCQFtnfMWIPxXFupmommf/ukl4AV1dyZIen
AunN/IKu99FXzq88vumaetWxAX+zwgKrNlYPtIaK7vkY4YylFk9RSSKwuCbI0MvRSWrTZuFneKcl
bL+95fgYE9hcWeY4s5pOeDAYph1dFjNIPVgY/D2hz3cJyitpDMEF4vZPHCarB+TOYgFnTIzHro1v
tjEAu+gH5VmibLcrxdDLbWVPC/So7Rd1uTRV/hgfBmPjzpARvcXXxuBtBvim8swpXnylzE5m5J8n
U4XhDrLOY+C44K1Z06JftmFKVI+NCbqDKRWhwRhkMIMmYR+HVPBA8TnDJ+hZF+KsVBxD4iZUktHD
8SDLuJqjGsMOmmvMecZZc0/xiPzhwu10hgT+l2byBWoSbfddw/0kbgzkLjCNElaSnKjpdFYd2Q+I
HAv9uavMcR/c84OskRqpTs5h0sfa943q3JN10m5gRIfg/A59/gw09hqr5rHAfIDFE9SjwRZVAA0y
r8HM/CKTXTDVPKwfaMLDudNLFW3AWxX8XPZVcBIxyeG2ba9V0tEqvzlGbrleQqWHBoQoPTvpjCke
NiyR9IGCulryG4tD5NiWxLqskUFx93jMTpTqSv+LE9sO37K3kHvQ+MBiPjI9UyKqk3JeXs9+p71v
J61eH0waIytlbccHyFJwU8YqI1B2iK1WtRYj6qyG7krnzFe2FLMd29vnyItrGc55VawKY6bkAngG
+gaV4YiIpkCJ1N27aF8ucAJO+/J8ok0eth2BJCZjUT8+AWhE0xYQiXduL/roXQRjSPqBuHjSHfuH
EZWSDyDnvQRsN3fFix4i0oPETREBQwb08iSzA7D4BZavUZIb0nbS0QZ1yDZR7BCwcauxde3Q4lCa
jKNEnRNyl6zpGqzKuSlx+4I5cA0TOvycq5LGoLF/3TSk5woh3uYQ9S0t3bpjen3EF8jWOEzsJaDs
d+udJFxipqRMvBvdpLUPLYCrwqWFnuJzn1IW1QVuzWKBXE68mHuufdTxjAsilXt/2ba1PVix/3R8
zZj1kQBWfyZeJGbHSBIZJY49bEM3gTashi5GvswBw9H211FuCfC9EY7f20iTQbiniFjyOBjw9fKZ
WBWwmS9TNHaJbcoyGHHpATf9lnI/uuSXY1XsIy78zNXMeBZ4tFJDqRedYI/7A/4ZArM6Hi5ZGd/s
ST20YXpWHvP+QJxE3XnKv2//fY7lBLM0mmD9H7lgJr5GmI/xSSg30OjpjkZsoxL+vaWcJg7xt+Xe
pBk9tmbPxMn3cp49Wu8dgTvNXvo2DD/ulmK0AiDMDizZMdTA9clkm8zxZfLgQG6Bf6zQgMohzBv5
n7q5W0bVLTRqWEJlSvyifwSvIwGC9+k2I77TcRN5vE5yURD4YxYQ57Cb/DK1yq7IAo0nqVd2sV38
iGIrrxvQTcxsKBoNKAC53WzFiHC//CxNyYHuqVFYsbFn2whsDi1S9JQAG3Yoh0kO71ubfxTukSGr
BD24Y4werPJVvTo7Ap9T4E/kQL4DfwHWsxmlAOU/Ha5YcJQVrCk+XGtT7o/L0hk4bBHWd5N31Aa2
cPQ5zntNnlClKgqgQIo6T4WG6UkJIlZWXKbt8UR9NJxyMrIXdpaOn6pWLdCQX50mtkQxGMRMK0iM
02BUkrKRWdAaVlIvXbf6bOgbMjkckpue2qqdVIJjKV2ktL5yd3SlFHe/Jwi72+OZWkolITdKtpJ+
nFhgrpeOokuMFdHsF3KRiTJem595M4mcoIeaXwOTJvPqbYYoEY3WJWO61k0LmG9Hq0MPrvI+iagG
u0R2fYd5TfBQfhBHGrDAoZHV1PO+fagSf/N0QLpPEQ6YWXMJCKuTkCmsuyQZM4vy71GEsOufNTRb
+3U7N0nAWI/FIwsriG5Nbf2KNYUyU7KfOzMp+q8OkFI56ZzI5/XtGdKakkC7hv2F64R2uwpNMUvQ
wPkPzeen4VhAf1cRE+PNZFdegsUy0pDRvHWPJGNsNpjelHOatrbWP90SLL4LMc+Jo8Md1RjJnpay
74g8Wa9v2PaOq7I2rlHeus035XlwNvAipa4h/M0Mvili19Pv6v3uBh4fi3vAHHk1BuTuIMFdGKxX
zGEqK4rYX5VlF/G8wDDV65dzZVe+yAR+gNWiBR7fEtHSPPbmJ81zeA06HSofR2Z7+hPncH2d1f0v
ww38PlXlK0pCl8dwfIGsaKSNi+s1QL9hQEckHJXH9AOfaqs897xeQ1/cDHMEdMbOTKzAkBs8sSFs
eYVuvqM132pn9VkgMoOv8Qv4x6YcX3f+24c8RyA+Bjq6/Ly7BKnhri2a+BsyLqoU08y5brv7d8rf
s4pt9KtMujssJPM1lAHr1P4WF3ve396K0X1CLo5H5OIys266uhl65vCXBoMv4QEY279WHSXu117P
9V2mA/F/pltMkYAKults7VzEmcoj7oQp69QeYpEDEwMiaknss54G6yGFA0Cl2b6MXouKbZ6XhAKw
ZeJFu4S0Q8XKLRgU7mcCIcXo61EMAhdjh+wgurd/VKW0xsRAxLS6M5XMsJJu+sjh2Ei7dNVtOpEG
j/zBHeDXjRceE5UXHe9ulj0pKZpohclxJsV9p6cnmPfQoFOrDrdoG2gmfo7PsEab+fcfDAdj0SXP
2VKfMb7kuQIl+/lgt/iY3xyce9UB61TNiCfSw6Z12aQofmEdnLSyPqQWVsr1lyDKKCk08jd3J+MB
TPEeaPZIi6n70NoXZA48LpWOwO1yovB1r6fB6X2RUu5N811vVnIvHEGUY12D+q9m5L0TYfuTbbQX
xpjl4NMgHr+lBfeUjDJT1DNbylBG460RV58ScSkUdbPMKY+W8yp2GExL42iwWLqF6bb4SUpjWnfL
P8x0XNtt5UN1ktL+Jo0z8k1jf7reN53K4cO+9lCDbcrdtMshNdjQScZv00MzmLsVAGUpn9BiaGJV
n3c284+r1FUaku8ydsvO8dNdCERqM7ON74tayZOF04PsepbJ+4ZYHGX8pwDAvUiycAecVsR6qXsm
ul0oiEC2yHdOy3sCNHb2nxKuxBE7XIxKD4hRMDYqoaSloC63EQjhQ2FW03GYZ+Q89Xiyg5TbCqDj
SMS7FsxWbNRqWc33OXSR69B11xCl8BBN60DqlcAnUUAJWtKoBuxgd4L275VBgZUm5ZQ3Idzymf+G
AYPpieKrBGm0kIyXAxccRxsK+9Xcbl1BF0DwYpQ2O8NVkSEn+aRiYNQgmAkG61id9tk5qzmDklDL
pSfy1V+PBPNYLiY8ku8rrInJn+XbSRYC9QRf8+FKi5YcQHj1bbwt9wJTo57sQnPkpsRjG8FjcvNz
s4jRKnG14ZnQqu8j5V1zx8J/A3vkp+u9Ei5vJ7ReB7l8WnBpJyOxE3SBuszmjOS41O1b7PHasCPz
bO0gNxl2CuRVUa3zawjOYem9B3isLMxK07Y5QAQEhoqaytnjmhTNWbj4kSa6yGh6PIoDavUBnExU
T5KzxPAyTqmX8ZRwNfncE33QIW4eoJHhoiy9Ts2s2baRWIyE9hDnVOR+8SFhXePBEFnAdvkn2/IL
Osw97cms2RRHQRdWapCB7FZeWtlmFb9zVq/1wuWwpFIlwcUZZg2Q8HiuoSwKKIJcJpF3AiAuQxG3
6njXsIPnFi+gFVXNiu62gPOIU4CeayTIPlSUp/FH5ieVb7zJ9MtvKtQNHIEd1td9epSObOPr3sAi
LLdiEier+/K7bll4InlCkPCRW62mAFj9tDUafFpat1GHvKpQeuSDR7sBd4cMhNC7fbNT3SaabizI
g5VcibWVS6KYtdEf8zvkhrQmi48c/tPLzx5WSsAjCdX6vGbnwaTqnb9omxe0G7fqF4TG/l+mK9w0
fBFkVXmDUKxmoyMJ8At/kZAtX+SHI7rbyUetodA6RqYxGczrK8oxNGxNmFbToXqY/ayrXFRfaEIV
i6GEPiEWSehATNWqx6mhz25oVwnm8LV9+c/JMNH+0Xoo5cMGaB7NBUv1RFhYE3MOJbQOddSd2O9a
RMU1PANGObQiLBLc0kZq/tIy70qi0RqiK0UPNyKQj50FMFqh6JqDNUcyKR58lCtghuj507HyEYin
oGV3vw1As+ccx63aVLlPyR0Mr3Rn1/NBPrbYbxhkkktq81Ma65VfYzcp81wImoUhxgPCh9nVmOIL
vC0TqgVSai7m9cuiPzr18iS7m6s+AhgqibZjKslpUey8b8jD3Vwv5UpAYg1OoSc0SINmNUzpC8qA
6u/Wd4a5af9EF0w812S05ZyhDIv6c8hqNNa6fuYJUSARhRHpc1G+GKNBBZbH62wGGRX+VXbXF+gY
RW5cSxJfXO3zeLehpviEMIliyTSQw2KG5WwgUDvRBf7fV5dS04K3CR0g2iTg1JthgiehKVNz87yo
RSTPYQ8dt4xesIzysYKrZDQblSl0cT4pKI8/n/Y4QGDB+ojsyJkoNiFO69J0UJrgVTyO7h+ddA7u
lhR4WfhW+Z0gcRy6SKnqJL4EDZqr11mFRiPM6FDvYWtktYK7kcGU9K73hepfwgu3/j6N25Mf1eHp
rDGb/TmroDaSE4YRvdXDuNThTZchOjBCjKoIW2RlD23DR5bfSKC0US5Nbl+vgV2MwDQaMb3Yngrt
S505QF141PognZhPlmoCKAWYlQ5MQYrePKvs/qhJHqJKQ4fYnwQQjWE44RiVt/QuS+QjBMdP3TWL
ck+TnyGISidMSNZS80C1Me1vvdv3sM5RO0VAIcUGTf8gisVAYikJ1w53RM11Nni8AtALm0eSo0WR
5r02UcY76LJL2IdZ/vAoN/zniYh4OKmDVND8W0pNJ/c2Ed6Pu6BrjM1w5fuyKTep1RPm01W5KPRe
wwwkHBFiSs/8LzNC0xf5raejHSYO2Drqk9fM2n2fZ4cYN0jNb+vmCJ+1IrdbhlUcR265atjqq2Ig
AhIFqXyhu7hdqKMn51pjtOpXLz71UHcJLLvPDXUxJVSbPtJkfFNat5uME3EfJaXfYrAMnOOj/kkp
vhPijDjVXgfOBkQMeE9+oBM+gFKTXdBSbPTSRzqHIhkOBD/ET5sjtiGksXCB3b0iFcGlzD5eTLjv
qzdqyvpn/ohlxPDybWDStvWK6zOCAdnjEDFjckVqvrWiW3cSglvN8hZWTDnw5yxgQP73Lw8BDuI+
CfZF03lPD2NRj9lZ+G9RTGzqhIjk/a303pSTGwV5EDqrTl2NlOL39wnWmHHOnK/c+ZxGUSVGrTLd
bxcy4uL0P5z/p1rXLJEb0X/BJB+rMyeAvz4cw7W80oQf4fCqXdkk77VLDzngWTiSwkDBKhOlBQuu
+dH97IFx/hj7g9aWBpAcmynSaGDlw6tI0H/27aId4ChFr9WHDW697nVCS9qgrmZhQO0vD1BDmUpt
YWFQaA+RiSMjz/0cmw1KZZ6Hzs7DkBBnbCWnpX0OuNTgetREaY0CO/ypvwlkvRUH4zxx5pxZMjOZ
oCuREywF6keZbD9VCNqubTSNYWA2lnMK2YDzyWzo7XGEkoK+0yBzK8EadBWXjhSO1KsS1a5lSV5q
A7Yy0U+dHmGliKGoH2hHChtUgf25T8hxKHS8G8fFmQC0O0r+DoyX8x1ImeBuSgTm4wdNVYIMfLGK
RR8XoSta5ZKG6LbjniOXxLJev+Td10Y+jiC5jDYUkplqFboRDxUtfR+HumfYK4qr9JK5WiwnUNQD
m3SLNqNCIv3UcQKHdwegp5Wj+3tyFoeh3RIgpWDIWlNm4QE2agIF0ZtUgizOsI+c4cv/5KCfvGGf
w1e6Y/2bl35nvLVlz0NPS5LjNSEvLiEh8LJHZj00TENSD3tUjZh2lFO4Pktir8/g2wQsutMqBmvQ
z6gpAftZhhEsFq84IUVOpamDzJiALvvDvEIkJoTHYwG8Gh4J3zc7PqOCBKVkwHkyLtwQNCoqckFD
/Bm6ySwKXuJiif/5jsynutrMBiBm3RFPYd+CfFlpmO9vf56RTKL1/vgAerr5guAE7k71kFN4fjth
Vfemg89EGj5HWbrshw8rVRWY/bVBGWrZs+rcV6h6VB+j47s3C6UULzWYkluKotQVaK3qzFSWp1p+
fKwV/xlwL6oX8C4D5c48i63keoWXoQzu3l0R4f2+6uD7JlwYj5ZsNEdcjOUHUjdyUYypbmjOpX/S
Da+vyhPqLptc+D+B7ZDSlcKctzg168C/Ow0MBZT4wkkWDVfZNhAmJOuZp4VI8+72Z2P7nwSdPuWQ
HqCNfArUaHcLyZmMLVd63KY9qLcQyhffQk+N4iu/6aKdnYbihYnhzQnT5dBg6v4jr4Ki7ui07KxI
DHhXnrTTyFfINqoRTamM9j0uL2/esK+dWGhnUaP7X95yshg2IjAEQ1+KI1+gyQPZyAuMICShEKZF
vQFrvO253LTbf6xfqlFRTBGlZLwcY5wtygtkiJLFt3Hpfv57GN1PQ7N1FVseuIfyoip3NtWL6+uJ
NCn0bSXHtg4uGRF1mHczvJBu6oEUh8S+jJhjeH9Lu0tU0MefrVORbjoXhhpJKuYSauyiM7b834pD
dqfzmSLpl0rrXD+tSPlYc8j3xf4D8ohinY+tTSxlINLP49TViMjpFnMQfvAPDQBK7ksbxP2xpoEH
DC2+1Dp3lg134rdO2DohBKMMfr/eP7dOiK715ipwPCmlksoTI58/wRhvHC3VlVwL29YZVdXoIeMV
lBXsiwFb1HOVQ3OWzdur8abnOKR2+51wb5x4yScuM/oFwlh0KkCUEk5We/xQu1weJBxcWqh/m1eT
iVPeHDMCyNfrHq6t09sEqST6czVN8cxaiiyOR/VqtziCLC3Q4B1BK6EmgzFliyCMZVRoczIYxrPI
48bT7XjWZ+Em8qYOtvTIex94UPtiivNgdyBqPXek7Egyefgfot9Dh1b9HmzSS9SgirzEgZQw6qHb
9sX8885AfqtR6XEXhiyOd1e8a+t1FM0rN3BqS0JRQ6uDVKrIbk/fZWPVN8aCWjiYyjq1CM59Xf2T
DS3TXkMVaZ8+VHjLKhegHnAS5agXIcWSeYCreNn6ogvZZrE67Krx37dx9sdH2vB/iR3aB0yIN4jH
hq5Ufs8exYRR/C/eT4Gt47hVKAVhdOa2zGVSYhoQHco/0nVo3A2RuWRZ7ezdkEBxJg3Nqof3svzt
WXuC6YoCk9S6ETCr9ZvFB2pMAYQ+rfT8s3WQEz47Uln5VLVMiA0LYRyxqIdVakk0Db/8aygTbaUA
qaL1/v/OFRDokV8FH/fAuB3lPD/kOmRV5tK3T3H/QflmQT83LSdhVznPBF7wLgqQb56rbJnBwccc
Jc/JBIb3ZyqLODRKwViOGFxHoxM9q3MJE0/9OCWv6PGdaRwOPfMYPLuRQCsY8Jzw7O/l4eQrHKBd
5mTj1AIS0+QmecS/5lRR0zaARJ/OhhubDr4VhmC5iiN/coQY3RsMnKCesjQJjZb/BjkCbzhbqHXn
EvAu7cFDCZ7LLWnH0KHZcAxgQJJbfiE5TJZ3+gul0vOCojO5mEYcaCcvhn+kLxSVZ6iHnUNUnw5U
Zm65k1jH1kMVmKwB1ZOJveT7mGuPvRQL0lA4FwjlBzd1u8MVkCw7a6jVhHNPU7hm0MNx24nZcNDK
y5+5WpRwcAHnyDDUqVNaFccT061DdRap9JLLCauIP7KwHwrD1MFlHv0lXubgiBHhu0TjHev1yKgt
qxm5vv+QSpWqwLHUGAAYsWkPLPIQnjsjbwbo9/7mF1lptC9igen1uh8SJDwZdP8Swpxz0ROJvMiB
qAEByzek0KtUu4g69EV3GSv+qIKNZSLvYpw6RQzae9/KEwwEX7rQMYzta1aubi9zQbKNCiIVmV+Q
/p2n4kccTDdYCw7DM6AFiY3FPbvyN2xpTnLjR5duxNtIcy3slvy6FKSblMNHmgtaW/tyG+ZGU7bC
gjsjtBPHYcsz26ujnSPlARYBfdrxafPi6gzotdJ699cJBGNkfJieUj3xdjgtj3AIKIN3hyMDdkNA
3rM753YuQflaWVbu4gHhQHXGmsOh8UJCPXUGnU3AcXiFdQbCuTPf0SsM7sqawQCUvhYi8jyEREu7
ebEfnFVmbo9FYR9WqDwwwA5+u3PIm2gjoMT47xU4jC9JfLzt7n9E4FFmH0/7QN2AcIrogZQzmWSv
jZdbt5RpV/D5yEFFtEGkxa1R6dks7ncJ2/gUPyExkt3QvEWWUWGaA4Shg0qQ7Vex56XfERIlh68l
Urb1O6u8M5sX0P1+d0z+bKaI0DRHClAv5+snxGSdOsXOgqX/OhjOjKIdZcF4f/cfYoslca+TquK3
2dZ3kKBQLY/BN1NwPWr34HA3MArTh5oQJLbVXhwU/IGAGvyzdIdu6i3qk34MvAyZHeP2mNyhZU4O
fZCDzuKTg8Odigk73Z0oOcDqJZKhNnYK6Pcgh7LY8hjR59PprXHZ5I8HFQSjYHZs4DYjlaQ2Ilin
Jkuhp4s6If/jbYrtiWhpfZEuMpCvKqm7giu1f0enGMBF4+fGfO5kiyt/pGMsrYIOzQvXeAsh4CFS
sS5ys7mQsvRX8PrXlkT+ReO0JSXCUU9dIxhGkif9dWW96qa1Zt8uLc4TRRDZHbBrH/EFrvzjnils
+/v6V18jEwByPuQHCefdyZCNSmFQVhVpuc3UmRGnfKsPX3ai6yGOKrAGowZF0qbgJbnu/mm9PzpI
bwbUI9sv7CPfMIcGc8vHAvqTESJ/8yhfpGYHPKll9jJmQy9J674Y6ZwfsMa9gOW6vx+J7gIGmj3Y
eXYw7bjxxtUz44SdwoIkQTnnR7puHJI8/SQ/Q55tEczJy0aCzfgiRUWm3yQ1hGd918ISjWNaEPuB
L/YFxyYoRediZq/mXAlWuZWY+g5dgKkczmMXSR9ZKjj96JQeUMxyqLNTTPyn5s+aYMqsjdLvmcOM
audc1R+oq3htjzl4qo8V9o9q1xrfUL/tO569sOZurfQ9xO+yt7Qar/CY4yUnmUghJv5tfL7Siohq
+YtBc8ypVcNOUtJ6L0rD8w86bjuO4tK51TtROzGmzvoqdPl9liwx018k8Hm4jtnAdc3CuVFSDoOC
nDoGENw9iZE+CqlSYqDuCZa1Igg/MsSIISr0de2teZl6tI7dvCKI26zE20cWn0cfnQlXtuorI3Oy
w/PxIzOlwAFtvpkxm3neXMt82U9r7yDnPkE3EZSpWCerZhNg669kl079WG0AID3tVgyej3+G4BqY
QOKV7//BaShvH1O9cEBkENVpCmlE9P2Z5xTEu82Hh3eDBCSunHBHZ0FYywJvoB7tfZrXy6Hqi7Xa
obaGWC6RMwzlEZGNxOiBdIhTjOpesrH2LdofDwvGjH1HFqIT9L/UQUR5hRrwouXtyTNPMoNEyr/g
XvO6V2trxsLGZrjye6r5Gtfl5sL/nJ2oNbtoVVBD+i5aFtGQP/BQTubFQRoi3owrG5K0zfpkMgHG
au/I3GlI8NWit0SsqBMOX+mavhwuAzCuZVXsmEVB/ls6QOvwhkMtiOUDtPcat16Fgl4+spirdg4V
EONj/Y+WxG3KBLPJ8TG705Y1FWxA1yErK7BNf2GxCeSAEzMyghBcOgoEigIJpJ7L4bEQiy5wwVkI
W0NPBZCLk/LO2Z/m6KlVWOIhVKav+IWmx+AHP1H2a/cEyDJIxIWNpXIkeSiIvuCRC7b1u8KJIqOK
AWJ80N+I/UgMQLjjJac4prMe76l7h+qlhsxgJsfzAWcAsIlBG4Js+9Vz/Lx+QztcpGI+WR/iMqNl
+GeTXIK/pRf5J7Fq9Hw0iIP2V1SwwqYtw/G0uzD+/sLWgg2NhCjdE72LwBTqVqy2CiHxp+uZmYHN
OFZu5cGQ7+9MRBsNysNjvdze3lSU/FbF3mQxS4AdWRlof09TU/3Uw5FhVYdJJjLxPQObvazppoOc
0KlZ+bfWOcHFJ6XvGl5AF0gFFEWE0rpuuhet1s6Jlx2ZdJQCIRYyIZzJ2+Z5y9WL9U1AT+5Kqvx3
YvzK/TAo5dg9wTWpkEYT92IW9wt+qwWVYNLZvQ8lp4iH+zXMoP2yI3dGHCqkwr6jbg9dk6LmXhkL
psXcsH4gX7pMFSC+wcheYh8C0Ecov6fdM0dcyq12ru8OwBjUBPqtWHoDAUbTtXtfgbJEOECZQmow
OI2TY8KEi5EhACYhNClD71NRqa32VAgsLMdzisx+8xxBcZPqmg1BRMti46UT5NumbZS4sqP3WwfZ
0x0mPXhKDxgA3tfoT2SQIz0cINfiMr2UxyDf6A5YOKebHrjtWHRjM2S12b+bFNV8lGTC7HFtdtc2
f0fwX0+x2Qz9MNPtUw9yfjvXI4kUueWKC73hJkctHaszZ+0veNScuynbfssPnx3BG662BA/IzubY
p+tzrmnr0TxZQc16GseafhmB53RRvQwoySWzcsal6/4+6k4X/0MV4v/hA7cukO6TB4o/C8NgSvLO
yZq/9r+bQt1z/ZLLbaaam2QkV/rrplkvxdWSpzouyx53vY4xAWsMRXaoJfEQzEJgW2LNgVeyMwLi
VpJhAHcCSASLWtNGJybeEH2hjtTP6MWkg4tQyql18yZJq+93qsnUnOcDxzR2NolJw4728zWGE0Rw
0Pel0mimRBrOeNVDsd7AVuGqVBfXmz2DfoF+v06lDD7/RqMQzUQ3FMYPTjuVBi/aByANphrRTuU6
l167xsLvRPiiVHWOdc/rVyhnO1vldxmRiB+GvA/iq40Z++gtncngZ87cabyp17ZVq6EUURVlG4yS
dyioPOBiaR+6FHiHhPcXIayox4o+szi90b13/AumT7LLTXhcDXEMsQpZ3WaPvzOYJiogGwh9VBML
P3FaWS+u1jxFHIxOcVYRH+Kj/ASio47+Uaaz9ZE/NhDC1hyKOTN13y23qpBJknNmlVEvStDJ/dMh
z6ln9kOAvhmGA3igEJwvRMS/iK5lQNDZCBS0hcWFSJi5oyh6hcrmOoeFj1cKyYb8dpZrkSsnmuOi
mD2WjPbkj1DMXUPqR8WfmmEdrSbfrgBBokaw0vqFjoCXLM1Llb59fKZMbgN7rOUgf/ac/OZb+xwT
46ijWGyme+z/y6PXcE0NIpBQH3Kjp8qUmh2Vual0+N/BGQLV8QZp6b8b/tNhLqQBPWEjIil2LqFv
6U7mc8A7Vng7DT44ZK8BBt7V1Z0wrFJmsKjsXhlCxG56QlZadAuSi8D0j3PVvNicc78my6lwgwyz
ILHpC0Oq2YrhkvFkg2qHO9vGoG5DuhtepjteoDihsLNmckVkV1gxQNnDG4jvBWKD7vKWbY6XkbhI
cwWwxwQlDx0vxB+k/rR2QvgXhgcAazMtbyadqmWrgPmzL4Hn1gGdrqa7TXmwgl/byLaXSdN6cAl4
gXiROUeUA/SGOuGBQ87TnpnCPsTc4tpfxMuBMnf/lEh0ji3hzYxdDI7LdWvowT6qfa7+7WhcjBh+
bVfJscRPaiQAsUe0cLU/2+84fKM2o9Bzc827NF7X695yMIFApdP5jnCMKMPO90TgWWlwtIctZwi9
ihX0xSfTZUWfdym8VHl3TCB1BtJB+cWPNH+8a17lDuVwZKI0jtcVGfOxk7LQf4axhIwGzCklWOeh
zgQwnXEa1j0yiGxtutqhFy03I+YFcVoAsmqIftpjKibPAvPBMB2JKcdBMOYMCJ9UPvy9UvoWGglA
Pw5JrEeZh5fmYn/+kpXx7BUmmY+VeaUFEXLF6Hr85MPAj134Yx75bMPMMGXNfjZ0ynQZj95Cmx5a
PJhpk+cfD3s5P8DMVQ8OIctih0wz0/mEExdRf3HM+CBBMxkOLvCHzNOVqmLHVTCfa3ZTMHBh0sR+
7OFf90JtG/epi2iSAGNlwlPkk4wqH7ePBQFTeREWPFECXNwHgXl5wgfpMJlW3lbwpMWIdq9e+CUS
sqsHvhHAGMn+5gDlmMEjFefWdWpW4vdZFT6qpG+2bpSFV8ShkUXzH66BEQP3WjpZ4BfYwdCOV41f
7XChlaGuMxoAeHAxdsKzxBkcBB7rPVrOAjchIlE/ZVXAnyhajlqns0PSeHrOj0qyouyv0CJgh9ce
VVpq1bT5lEEu5vMAWdXTeqsQ1P6IMxjHqqfCTiwfqzSyF01dgTbaw/v8WKQ8YtKKhiMXTJxUufkz
KKWCGtqDXlw9p7KzUGIYnq6PxWaeJqyov2DHjifkg9r6Ld6RbSbe9mYaG774bUY7XIP3VjRXXLzG
MbVON8h2eicY51F/5YJXY40O2c33jUNxWX7k8VN9a7yiv4DrTNMSNoangO/I/o6zjfIFnMHr1snn
Efd1AEDvH2Anab/PEtfZNxRm1lQfdr36oZOr6NOU9uHNey3hSBgTSF6ALAkt7vZ3wsZJX1fzGgFp
SV99r6N9AW4TxR1xNg1gJA2ltLDWphWwQCmzmRUnqIeCqJWqODvJxw/3yXclvj/lzxsOlx7t7y5/
eTCCSlDYSM4e80sMDFKBSRc5zDW9dN+U6KDzU1RwXKocuNVesqDAXUqijGd0a8Ycv5Ci7WQSxxbJ
kXmMGgxoNN1nM0ZOO4cgQhFYxP0z8GP6F6C+/uS/yw4SzpfWekRai6F/xAvabvj6F4L5v5SuBCAn
2hQ0BtZe3I5Lx1l+j1RB5UkvQzQR/fw586FZlnnUXRT0pxEmUbxFzC6ahTwZsjNE6KpyuE+Hi3Lq
aI9AIVvMxFB+dnmp3wgD8M45BOpXMJS0O0q7/mpsg4R99kbIlwytCczqK5+DD9yDKDSfupJEkkB/
V1rIi1vYswA8ROqYc4H+4StkkUFfkCVAs9DBKS5yvXhdJINE5IPgg0RR2ACa9KYadLabda9ZKNPU
PlFsNU3Fhd4r7CO7kq0h2nsxjxs6BLR7/cswb+uGB180OZiGeG9MN6cStry8MGZ50RiNYUB6G1ht
V3vZf7wCiYcWja2CSBx9fiI7L4s9+4bKl4Qw6Lb3ErNHO81fgbA0wc0jXES8pRJYw3Z9OmsFuLdk
mCaCzZw9P+t5bCGTyKDfzCdecPZYKPLVYjzCZCsphR10pqeFZd9s8QkQOTJAdKHyn7db7xFnizwe
OQjuG/WalMaaB8BYl0XXIkLhUpNorZ0l7fP/IvHHjBitRfSI7koDrNymgw0EkkosBLJn5W3F6cqy
Fep9J6/P0uHNsMhvlsZjx6QkKMsONQPwCtU8ivOkgTWhyz6A3cz76i9UCgx26rdsDsVJa7Spyswk
uZH8KcomMQFq1y88WPr+ZaSffaMGcuFVUCMD4OErWwbY7nrKi+INxJwi8IMGDiuPWEN9HiwwjSL4
GxRLhLLMuPE81jwpBf2lCGL43okBGU9lN+1A3nYkcOVT7rL475neegDKj3G7ZA7dY0RAbamQM6c3
vTOi0FPF8goEz0Y39F2Lp1HFd+paeKF6RyjuoDW2LBdjgMlm7fWGyZ0LGAz+Ugs26w9xafJNp8pL
cIaOg1GV1hAG2wiOuDnxXpVko69D5p3xVDNYBpjyXp8SahPOnw8iJJ946bl/nylJB6RLYHHFh9r5
e06IQSKvy6uEH24LuLSeuOm+BCsUw6z6YItAkI3RKw/3qn9DbiPlnuDePGCuGn+nokawsSzOZycR
FMKDoaddObLBk60aU/VeghymUq+m+RrcP/hAnQsxxNGxoItMv88PGyFVw+NFX0cdaK7YyWA1uezl
Xyawi62fsncUUS4hhORcuPHvU7LF15f08v72bEON3kdGfwyrPYM0tZt+oCyG2W4IRTwUW7Ns1sjD
3J1ealfBtG4YIDaydeSswj1HSdHfsd4EX2HgR26g4Pxe7aM2bh//crP/QzZaO/VI3s5WzBKoPl0x
YVS6JoN3vOog5djNXJUt/ZINa/edhByEoKnSFo6yhEX85+UyJYj58kQ4LqrjKdN/Y4SnDQvdnxAU
DAEB+lZgGogO+RXu4AP3lOvkjznAYqN2H/0c30mv5gVI+nSWRh0d7Wq4viGo+HTgQuwT/eJFcFU6
88NuL/3VzKmFDWS4VZuUmo3YpBBy3pXJXiAmwsgP+AgLvOoEszjickuivLQYeKrqBaU5Vpab2bt2
XRQ+B6rGFXwLuWVOpt0wrpOkjKE8ETvPD4ZysKcHZwHTaTrPmBbndKZjnbgcOOhndsptQvcxWZoS
TywlFGQY6CmGEweOewlFYdwhsK9gHaMKguE85JfOAWU1zXcZU50zX7NHOCxk5uyf7RHMAtRMeucd
GbGXNp4Z1kZ0bFUcAw9qBRSdx2QIOQbirWK7jtec8U7CLUN3+9Aw8ncBnQc1JqWpmDTVGcijhcnq
mhRMPoIo21TglCFLyutijKbUKcZGyhnIX9K67ZDVIrQzgfvWKLANlxqPkszmrtTK1McOqee/D2sV
YEiUMrvF+hPCUspNnRggFUgcjLRKtKvS/dh2thKIDPFyKpgFb+DlV3hi+agDJDncxL+x65R1Gy30
jTLlD0twqVySDmt/BXOMD5hQpWgPQb9TZVGQe5VH+2Y6o/2EuOx79ElIrxry+4wnVoTJZvvjtIfQ
Y8jxSi831qJqfVscye/ZlEdUzl0t1x2M/pkRQfJUrCGQzI9ywBcLzutPsSX6KQ9h+Xcf4L2np9jg
9FH406NUurHMtDC5g+CHPKgyEyK/kvGvPzgljNA72X2aT6weW91v6CFb083S+ZJKrzKqQnNqPVPt
p4K9STb4hAtR2nHjo8ZXmPKRl03zCBQuDMggX1u66dO9yCn2GVeCEoOi2nLxjHL1ycfNotJYSgPx
1Ms624mrLQAMarcbEV6NSLZwTiDjUTJ3fabd7twwucp3mJ2FIuirPv32gqBZXmeBXbO7FxceE6jS
5obknUp0dOdK19hQjHGrL92UZvEztRWfOSUAV5tXRUra3zZM9tJ6fqeNGr8YzCyibDp5NemP/poo
pxrsiDSK9OZ/exDwZja4PEhgJepvdr6/eyUX4J3ltyuHQJPBSumUMtTJnnn6hI1lQIQi0IVtESM1
fzZYdH2/P+xfHDJpSx8WYJe8oVsYBRyRkOOykZY4LRZ32urgVjIg0uoO0fPwaaJWEkocZi/jQ+fz
cK0/pveDeQJKOLlfRg6JxOQWAyIdscWAt8NA0N7RZ8Ds/RRYRIxCTyyGvOEk/e9KKpakV3PmgKWI
sbyRa828pSFt4sdpMJJkPK041Hu5lND9wrG7U3EUx+j+NAGG1r3FTsOTqlTiRNphSy6oDNinUaGT
D5rvmbNzOC1N3ONwHE1cmTt8u8cuvgqj4avdsNzaa11qD/1WOKkFJUkjTBrp6X9R4rFQgdp34jgJ
hxff9gkngfcVfLbfKAQeSgZ8gteEWrArDCDEwpgm4lX3I4FivgUdu83s/HouZv8vdIPFjpxjtqPb
JZBKzpSfaWo4wqCtZV+maTbj7Ggw6djZuPmFMipewP/UGCV04k4jZeKSGvR3phNIiRxuolK5wi16
MQ4HluY7l/UJ5Prddj+Jj9PkV2UGyzCpQ5uMQv7oR+R7oI0eAKcAIN61IhUX5jGzZBivRTfdkKmW
G+vBkLrqzRBopFpQ3yESo8xQXc4KBrJ3DhsHk3Gp41ZTSz/knR7iuiaXgsN1jH9kW3gO4wOMo+/4
5N0bpp6paR1Nm8HKQBF/v8+StX59/kd6UiNg/l0tYMCBrMJs7GoHIC4csLOyux1MEPmkh8VvRFKZ
WoxBNEulRLyQMLgRsxxd7V2tDAT7bCoHuRMzHk0KYRwwA64bHpaXlsC77pf3bEekK9JPtbW0zF5m
xEoi6rQQ+YQ7DbFUADpsEJLPGtp+AitBV2+tFiE9q8ggNn5lGjlOMGkTzvH6gKbZ9zIV/CUtMGre
5HDEqCmzolqkoUH/xsEfaG1XeR1cLdXdTQAgA2znB+zY4b8gUx5byi7NFMlV+TNy0wda9r9mzQCP
FY1ZrSGylVv1b9QA1mp4BXuLFhsLwPtHQcqpxPeijoOBWFjGfH4FuNQdxcxgsbljRU3ivgX7uIZu
han6hK7CEz49u9X6BhsPLz8UsIQQQnPRom0bsu/surmPyBR5wQVC1meWdTLsXv/dDlI9tmvmywSV
H41qU106t1p994rhNX2giDgywRH1YThDly5sbmOf5kmrS9bn/tMKyDWUyNoukxKDQmuQcRGbOUBP
rSxx+TcakdVHInsqOg2k5H2hGBGeJ0zfTryIGqphRqXjg9WfB2nkRFkNj/MmcOd1Vs1X4TDJ6nB2
yr5aPXQY5eQPKttQGiPNMrFpqNTtPteVaFDZW/d5VjAnLll/h7AZrQEO2w8XzaK1n19koXzkQeNq
Ms41bV/JrmJdWclO44Sx7iprmGlWnxr3TqbHE7dm51HJXsxRJmXEJ/XInhHdZ/6fz8FZeO72D9Py
XgcdoNsg0MaUGNapbRyBOj820seCDeqsDo1oJOTVl0bdu27b+PrGdx79evctXbY3gp6vMiEBP+vF
yYLoWAUsZtKirEh35iZCm1cyuHInnrCIYvAKtee8F5M8XzHar4+gb/MnBox4L7I3Duf13jy4Go2V
BkNVUQbDmOqfEcOcNJgfSP0xSpV0BHiyjfBSCtWSB4imIumg/g4F2FwU4TrGAV9r339GDQlhHyRd
51GI09kFyVMeKCZoHO+4EmEUfd2kx4Sfd/7QI2jYrulwQ2ifByMQrO4cdU4jtaatGWTuNst6GZFh
RmWEtnHJnDo1kpY21o49is4ofaI/2VFpb1ocYtB+aLi+NnJ8oyT3gP5R0gmUcmOx86d3rhCcbKSq
/xYqR7dcKaQsIQDwUVR6m4P+2O3kobjMmL3LlGYbV63qU2Sjadmkpuu4hvMfxeOYH0msI00CrKO7
4DZo6mhZVq1TcmFCZj6KVp61aU2f8B8cH3V4WFB6MAxkzV+NzqSz6u/ihhhvBytQdSwHQYnXcGyZ
NmsPk/blR4OWA+bKm6hoIHm2ih6z40eu4HyOSwYJfwP95XUBIMOBEOQQmgjbhxBrSIF0So81AfPT
Ti8Undc3VY9nrvrxNnPqzh5qIKiOUNYYpAj3odGcGl135HlbcFKXffDxLJ93ER4vmPj7w/yKomi+
WPaLmqYauqTELbPhefVL3Ed36+9nv90wouyMyawzSacuRDAxbAkTaHrLomiNywKnwwH66oOKkxeh
tV8kqdgoS2JZ1FjYlJyXjWKsz1rBENppCaiAy3AvE7T7VSceSaRx8h/wezpwzlQX15/o6SAgVMir
0freS7IMF/WxiQqXxQAdOZYGX6Z/fJyUh6dtVDWbSBCK3yV6v6ljKBXrpRBptax73ggQAk22oD4V
JoCXZt9/vrxxMiHi61Yb+bstzac0pQZLh3SzDumqUUCXmVSlrLIA8WgM1i28xFB6/OScB85sqc6V
PcqJxzoKpApB2QguqNERisGt/6if8fuRGCjfbvMnWhLAmt8Eyhox57q4+VZ/ejcwbv/YHuY9RkqO
MktTZHAqZzrKO/iwcTomgbPsIyApTalffiwibjD/RNJbDyMa0qxAc7rlDYtvm5Qfq71Pzer84TlH
XZyTm5Riuc52zPhVfousjynTPnLbYiT5qRE06YiL2mVmV5M6RZO/iHGAk5CRZm2DAWjH2sOfhMbS
2V2Yu3f5+KJM5KDRRyBSUEcNEJbHX8ELW+q1D9uMGAodPt6hI+ZTeQGSGFU1K+8BgwoPHrglJuE/
uzv9/iT8p2MmfC+J7ep19Uvr6lO+gzJgVMFvEj4a1sFvuMBHaAfTkWqAgggUUUxLL1flYbFN6NLx
HxyjCo6QcJr1X2Efv/l+Tp+Qyqj0L6bHsg6fmz1DiDOlWUEyJ4gM7aj2q6eUuL3KJ6m5g6FO2bGM
Gt8Ea3QrPP6jgUSONW6LIbpRHO6Xs0uaZdlZZTcYHfc/Npt/RWYHRaK2B41RCzvTrHidlEtw+3WX
uQxrVC/w/E7ps40N1hnsgH2qKTftmQyiWV6tE9UdpuUKKZEFk9jS3hzNrdxSspanrXzfoVbMtPva
ddVCC+NBG32YQAQoGtWLS5CHtYvpP/EhYuiBPd6d95Cymf00Glurb/Sg/MQa4WZMg7l0zOFl/+bS
kQM7BK8F2dFLPArnQ7qUgUJ6ccEVI/vOAc4ypYC/dEa/1RMYSdMFOIUBzeL8OpN2o9OnkOw1Waru
bJi71auuWHoUptge+kEVO64RfUNdLNfmzvKBEpdZtm7Ei0jbGcJqnQnw/I7hTVobBzVmBzCbI72n
1e+h+kEKU831jTYt9ilwBI6XOI4lfxYXCGUH+Hb5lpOzaCfcyCA8XDj9G8tF3/aUQRgKSg/e0DUT
hgI39/n+Wx3McUWE43jL/3w5KNnpAGQAy7wg5Rw5D5UN3QkAU0/zjdcSKhZgYMVqZ3+p/1NU9uJ7
/Tp+4kfwtjRqBCoIFDyxW5rdEuJeqdJyB2LC9J0TlxLWespsRPjgU0XIs3g23zjaqtvBNIJmkyRp
e9rQcotcYaCUrrlUvdajlJPIvOZr6n3FTbZTNd/XmyMUPW7vpkxvoql/CM2yiln1/ZJ8WLBvUHcS
Ix5sYj51g0wcu2QXW1P5Jz9EjW6s9Y4lmaGIkIC6PHMnSKtNMIE39bFrfgTFnrZT+u1aDd0CTd6N
IUgAGaprDxPFORw0GgbzwAX6x/Vlj/0c+Mm+G0xXOxYoPVdVhKcx7FWmq6TOB1Z2iKoJSYN+rOui
9hRl/WuIaPR4ea+1K0cpQyKR7Lm4hzS36zt38wG/obptoAg3zsWki0hhD2Dl4myHAzP1aKsiigU9
d4zqS7iRzeJVXvDcEfFIemwby4mu8+aq9lKcDQ4TpwaxPDmpuBXk1+3H6ns0RzYmFk998GiaafyX
ZM+GExmhSg3mCN3sEd7Z6mEuD5RxF/rNtG1rCoU8sDrtGcn+wnEAYL7eIk+wf0okWiq/u9AWNZZi
vZzLpiwP64ZrNQNqjvAGd/HzwecHIrHCdtOghp8A+YKgavIerubLAw6kJbYRH4Wgl5iKKudgtM4A
waIJ8uz5n3LuiSNAcPPjQYY+ZjMi+LzsMXtk+LG6YAYOXz8/Vi0aj4R8IpogvsTamPxN9ivoV4Bw
CmJ36SrodLQTY/JWdJm6m6mtW6jR+OeiXfrbE7zUBVVa+alZ5u7rtZn8SsYnvHbXsgxiWFpGu9Ub
WKOfijbQAK8rinBI1lXzY8GZpsvwPzqvA2T77xaPrqWHzeZ4CyxlhOLfQeU6g0GgtDl1IHrh1JLF
Yl3dQJ1vWlqTnpaEBqMkJwtn8QJ6170joTTHHrpe1/D/xsE69aO1ideuun4K5AOwyItOIyGLvj6z
FmFUgbwlxb+qtG9aZt9jEtd6Y9nQ0FCsmOG5uWEA5HW2nC9o1xSvCq5qS6PWR7xdjV9CiDxZ8Ge0
x6pPqbCIenHeAhm3AOH6j87j61r70k68ODyS4vbfe+jGFrlgrLdfgzHa6kug/MC7GECl/JFOQV7F
nwEw/NFM6FiZVY16McVtPzllsi2MV1mct44JQl49YKm2oOnvipEXmovJ+1+opASM1b64caY2MsW7
eyY4uqEMibdwoF2KOnLYN1Eoz3Y1t0LBu7Aj3X/XZnsqoKZuk9oTbMVJvLOPvA+xseFNrpjfeui+
QGDEHrq6suNjxPFl7JITs1zpyq0Qh1a8eJbtF6QULXsUzEYr2uuqHgMjyXihiQa4cc5p/wcoZ4dV
ig2Ousrnzr35MiFn5aBzGn34jDP+BKwrXowjimxp7jgcNr+uAJdgvs7cDakiIvHsJfPO6EToobw4
Il7tfSBG+FQOlboSYDfGkjw5smjnsPDs6We6h0OYcXGfpMhyQ1KCTsmIKdieSCS7VuchhvY3dvO/
jzxf/vz40HvLRgybubkGv09xAvMhT2K8kkBR6jteApuJ6vaPng6kzSViuV+KVHOMJ1DcmJK0axGO
iBLczbgJ5IxpqftJMFdfqQgLvNq9PW6VpMJZu75Pm5jbKgINmHJIhIc2zC8OpROugkeXaOPPyyiq
ExFtYYWu2vhze34tO1fLM0iGGo3MuGcVA2je94wTWu59yAAH5iSAz3oFhRLIQEjIRWYbvYx+TkPs
x84UQSfrfRDWK2SZV8yvxDvyAhoYeoC5uffc77zUx2e1DHWIxGocy8kqxuzLbhH+gHaz7ZF/wpbC
UyWK8zRSgoMvBRV8uwTtxwjjpp+MBDxNMJFtz9P5egxdF4KqNzPW90dkSjA98edJMWYZFEQ916k8
rVv9UZmIM4yWFu53eM1Y1ZVD2uZSOZ8YFHXlGewCRB+pDGYtC1A6BcTJ4JGUgRjsnbJfDUEBNITA
DTjmJNeDGt6QZVy/T1DMtEmCng6G9sj0y9k/RATqL80YEvIFq6lfniwj7axAR0jzrqMVd17d2Qoq
7cP0lheZIcH52QqR8fBUXzaRSs3EQxbYPjANezQs9Tb8LXnNDGbYiJdhsJbTAW5K96bLIVUUt1Xi
ersbFOlHxOSzJUkhX8nlmRDv+TPkUlspL9+mC2qLSRHAS+0ZFdnqSh/fdXTAhnsguGhfTd1NpO4u
LEyIayC8O4V37XVlRUVlktMpUC4WVoUbPOYf9s9OthQImF1WgPVsXgjLOyJcNnKZK3bJuk5olWzg
/9a91yEYuBInMrOmeF2njfGxu/p19mX3A0Z40qX3beTo4L2gYgl5mviSbrf/xVlc/yOiWhRi5qlF
CjXjBVKD+jiHAG6+SEcXjEBicPXyLk/zB17IsrNyuNWh00so5+X45/V61PhDSdfveiNRYhxcRm6Q
BGm1ngu2W+b31uOn2P1+KxaYv/R8svafwJtpQU84HOTWs6BpS2dnPuVc0UOa/aRP9eyOSco0iBcc
L/EaXZSmcXHdIkQQmCy39apjZCJF/0+WibyT3j2EYFkuYcUCz81zghIIspAjh1MIB7veSkLwefV6
nqrw1/l8rLplD9GzeqRPItjwX5MDEHc6bwOnJcw9Cnk55kJ6bBqcMCgRGBJvaLiT19HEfn6Vbjro
JYcqJD34z9m9zculz4KcMJ5mPNtQ27jK82JdiwGGydVhcgAVZNk7D70ArZlpa4SGbTDcuAoCqnfV
h3pmaut6W4ejHkxfttFyu1YARnN5xouW0Yq3QXgiCIFWQQNGsoZaijjpxcRvVBAErYqIfJI1vdHr
0t/KTdZo/5EQ0ow/xkCZYgHy3VnPXDEue8DHDBcNjYLAxeGBMYASzMLtqqxRO1eHkWHTBJG2Lzr4
9hVozllBK+2hruHrglLLrWRX63HRshSSEA1fPWpncFW9EOd4OhI9qx4vYc0wCuNKKYbS2OhGMQFq
nDMxiENKWvsSOS1FwiHACgqJVhP9N5Pp8/OgIbJavVlZNEtri8NOdKi6PkylHz1GjZfgDYjW9Ja2
jb43xYbIsTb3qMggoy7UtwCcCIdQ+C1sv2J2N16DQ6bRA/Sx7tOAxkcZm0T9NCmoZp9FXw3VYP/M
SCT8WdphmgPzZ1eyhRIX8j/S1D8fWqpzGJKkxzJDgnSg6pjaS+72GLU8z1uj351Y8RqiUIbUTgos
+/v/vZIeduBmaLdFdA+oQBSB464mA1pMYaKlvMxiaQwQyMMcr8PDtRi7hiTVoMIHTzL8GD715p6I
Mj2nufhmYnSxs9Fua4XUwjio7FxKbWIXZ5oUUZWeUqezcvK2jl1mVeEbMod6IPtrbBNi1WAFL/cT
2VnCdQZwsD/8AWy8Pmmu4rvHRWY28IPJnXe6jZbgNJWbn/M7SbooJ4avRELARMhonSQAi6Q4nNXi
uy7WGTpWLx4tOl1saBhBdgVc/150by/iTMswQqN3a0xTKCBB1pQS7RRWDM77bbP02J5Wd8BpuHV0
RZodTQwy8v/zI7kRoPwOHh6B3WpHZGgMRDDbOI0XL7rgbFmorhdykdgoPkhcBbrbkV/2arDbybvf
08vozUhP7ykCGtIyPMhx2z8/+D1F4sx4zblf/aXSR70VGTNM9aRPJtNdyzvjgSrutje4ngU0C5aS
hpslhhb9FYoD6NYOPQXr1cEQzl0XR3lRoqpkRTOMnln9sAeY1Q8bVYhyI6PoKMsJnpNCO7kBDJyi
903mDzF9+Fh8BvoLRS1dzK9yiNa3OjQdjuUCu4mNHzSPD/L/9uiShddn+xOL/t9Nzmic4sjlA5S/
d1hj2SROrt1ReX5OQfZZUqXZzoByWyjtDzYP1VibB0iqAdNrMAd9cdbbqljISLl/rDAd0stRcuZw
PV7DF8Q2oEjHVsmmnPOi7I9dIZrcnbva1TFrgBsKmDunAY5B5G8+mte1NxfauCPn7qezFmUlWvA2
S8PHakEwsLiYR1Uhy37FpoB8kpxaemFOGmSpodATZJp15jdN/JkiMkkVuqtJR45QLsmQzT+mpovz
EkEx3dZ7y4pKJ2PuQoNrPWHc9xSYa8KW1NSH9QxoFxiZkvcBrr79KKDz9GvLZy5NYQecWB/0NTux
iAL4USIZaKgbclRT3xQbtv/e9mlxRsoyXxSqckuQPWKNtWTaQSdNN0q1sTqGCJPc/vM6kV1LhgxJ
5rFlhS+Jq4PVP8nrIxstQqUAWgiDO2dElj8T2jvosQzb5dFafBM4qXP4dnkLor6w1wQqVJFwmJbT
FO6wNX3tWOY0vqQeLa7slD/yP8+AkU5JBFmxsQuwi5GsEfa3xZ4vDcWkXsKYBRnBXFbq0MOkxrl4
zlI+LCTHaKifhfZ/xSlCHwjbAc4GQxvXUngTomdhMbd+JjpsYOTA/l65Y0sbj1tQZu69eVtUF0hS
WRJgfNMQXfFhw9719KXc0pas08kWpyZiVjKyCi3mjyBxw5j5qKi07QAxtKEq0jxHlVf/6VxqIViO
jz9eWebspk+JBkQ4VAwoK8z5GGrc0JWkQj+4OVgQwZcZirxjKBEya+z7HLTcMGKae7ZYDw2ABA42
RlYSsXTIDmPbi/+jdK6fAYEDh3DtJiKIb2jc+HArhar1jyN4YWnX5G8iErffrYhsTbdrOYXWaUuK
QOob9Lo/t4O1VsCQxSkzlCsPHrZR4qVlrx3/Ky4QvxP2F4kVOfv8hLKrDFqksdwc6ZiAxvxf2vTo
rk/qU6ZqC4GEpAGBXCzFY6ZJWzWLorRRj5g2UsfuFSGA+XslxonT1i8M8bHVq0+KwREl89Ezu5Xo
m/U/8HLT5nDoqOyGxwmOoT+iR3d2GzUrt2sIuTmXNMbSbeCEH8JCWQ//QnrqbToEIFNSEwl02E10
5ioqiT0pyTNZUYPSmIVIXrhxhJyld+K/8jMer6KMiuJnfTVrWdowdzjTw0voIpfoQmJBZLFczNhq
KCX1/nIYuJSWUfrvaOla2OfagncUQMoEEy/SRKz8FtROhilc2CyZ2M3Iy/9AtzQXLsNj8D6Swz5I
YStMvVXXJCYHuD8dQO7ueby0wiYMu0XlTGhAKet3Wml7GNIOa094M1xPxAYuLzjtYzMvY6xk5Q3G
Ypo6mY195rfbWxs0QBGgEY9l5ijMcJOiN6IzryzHR/KWyLV4L6T6omW5wQZ68ocp9YVE7HUtVT6N
tsPO37SWTPKBN5JyJ1p9FN3xQAiVM6H8OgG60vYrXQtul+4xRecmvtNWoYSL3u39PH6e619JPqZZ
zQpHYQSsjXlsYcDLPLYcTFK+jlTBgp7iut4ERjGY7y8OI3u80Sg6S+C6GJagYwYHS44ZETBZWb42
Qvjcsy3pTwVfRsUSOP3OuHDeyjaa6+gXf2w+kheQ6Pj4EWUvinIYkq1xKCYV9/uE1KL3i7u/lOt8
ffKCNjJE918q3ZOAqhvoPoTtUqP85Q5qIzktheHnYhOYuOkfFWoC978NORdsXlrgGhG1ajDioH7N
Yf/q1596bzXXh7g/4vl8jsfp7UI6wGE5zJv+Hb+i33WogveJhRDGXApM3tGFZmHsTM0xgVk4YM1A
dLlFXSja30lw6lwrmvtcglPMznU3vZYJSVGabgK6B3L/p1HVQQ+c6Lhb/r+4DjrqHvUSSPDCqWIL
8f5R+1Nh1uviKachW0dVpvAakVFan3LGWGleYl/RJSwsgefkRPvSODVMY0OXs2BeggI7jPK//h5P
OG4I6E51PtVLYTnmajE5YC/RoS/Nbcm7rJtlgT6ByWE6Ozh+krGQ2c/9946449mXB3ExDQcY7eg0
HXiVz7UtfHGz1ntWsZdRQyMz3TvnyJh8X7rFPmggoPdxa0SXzXUVD8xnDUy+bjLK4blXOyOdw20x
6bbJFrvQuBjTt4SO73pAZBIge5V0obAshce2suqFiMok2UGVCnixhY2b84JH9MIcvgVNQQeTPvuF
FCBb6GgYo5ylTulc18pDwo5WBFpm86ijd0rgX15K9Byv6GXH9rgJGd9oCeWqnqCyhm6bjcd/Yl2B
/NIPZd7jVEEm4rj6p0b9wWLeAphqv5LZm+ANbSG72DBPCRI3PLWRMiZ6srnyEDiDj+f9STwNrSPd
N5qT7l38QIV2i4+MoVFqr0ytjJ5fzNOG3O3YJAbZWo6S/m1M/uQHUc8G7MO3uD/nohnMlZEyaGP1
hK4hrHRzQCGWNMxH3gznJ3OjttXxqOSK0eBVOofghoe2fPW5NudfBjjnt3ZVMof9IRRjNTAvZ4dN
vcI3eDnaPy7SoVjxTBxkgNKHTfZyyJi2jptp3m8f4HBmnIEnob1CtA19ARnqtZwf80ERkBMD3Aml
Hn6b4KKA/2h2SHEQkly0F7vZy5nvuE+kuFkOBZDpUUI9Ph4jj+WlJKf+HucHrjmnVDZINNjYAPkz
Arl44b8kvxzLv+jlsSbcwzeq8xCgd/dznDl1ccHCygcl+zwQOJ83d8rGuHVJl2xzIuUPepDQaExM
y9D4mNc3BadsgK2qpBjm27FXVSPcg34qdC9UvHEaSBcM4Z529QxSQA+kV+t3TLMSudJrhzdI5Nag
ShhPC9Bkxw9WdnP9XOnydR2Aj6HLiA52WYoh9+l3O3rXOk13w5qOVHIrqPZ8iRtXgFRTlP3KrlcZ
qNAPcbFG4Yf9b1EQahks7TVuBiF3RPDuhjjRELCqyABqjaPhOOSIkaRO8Qb/Uqp5lMd38FndXJGS
6Y0gPsrx1Xo6t1ylD7A/M9AdMwapCb8zhTdbWYucN03BcQgnlgvH7uGKksuIijdgnhGt4D3+pzIT
a65PkuMorPuPII4kfiha2FyWu3fcK3OKxf6lfxn/Ia4Qj+M9whLPbYAPdc2eDzXrEhR9ObENMMTc
WIKklc63mAlas9DSLrLRAKZcYY8mpIdGHDsmfJEsHfOp3NtH8AA0qyHFP61OqAs1QpIgBpHpYJjY
8P9NBO/ucytgF1Gda0l5f0mWxiHXBa4AuHz5y4ZrBYYVo72E08G/UW/UmAO3UdUrAio0642+NDIt
BsLi/oKjEB8GXPELKm3ogO5Ot1QWmFVXLIwJpVu/Si8uBqVoCVNnvevjDnftBfbDuIS8Lk/0hK40
y+uwzzxK4e4VBEq5zlqXY3bKQCuiqVYLbMz/sykqXj14lQAxVWwQTHFyBfSPqHJ1qrawLk7Zf/CO
ERpmS6b0y3YFYXef5H5PYdhzZKhzFD9cvE7b2PoAUA4HZbHaqna+okDtdBgGxH3CVOb90aoM+MG6
y+A+CPiil8MmqSiGfz6k+V8lgFwRPNqZKRfuv7K+IRcS2eqF5EggWBKZptSIO/VDYx8Vk80XfFFw
f1ElDRUg8RZF/6iCuqVYcKo/JTi6EGW+sJqkJcdRxGQBgR94oiN2Qi06lALEqXib7/jn/tqpyxD7
8zqbFDczOCYyU22q/IkwuZNHLZ+8YtQxzYtLBN5Gh7NeQxb5MfAsQIiMjV9IHGKxHYMYL0J9rIFD
KnvI+0PrjNUJEV89uSwWmBnSWw1ao3Ki3jpzTzXm8Nl2yhFzRyZgm8k51Tu7aO65++zBFPk+ZZoy
yEFQPbAy3m+wiN27vI9yV2vwvs3Vc2KXaIS4TztGkJO9WsCNr4hAaYi+V1RxC+acG0/d772YXRRY
L9P10wx2qo/ogvX2HBBZccmA3Xsgvz8w37CcENq1ud9Bj1SxXmvOzrm/MPCuR8axjHmX1d8RID3p
Wen8A/l8SGga2oucv+ksSnKrr56jUhXpY4mVqarP9BFaqYgYkIOwGhwIVgWBUeCsEPofp1q90c9p
KeiNlpuE2c/HiXAzr+nJE792PIj1fi0mbDx3xKv3kokwOfwDsj7s7ZYZMLmh6hBQcZnOv7NvcBJW
nLqhNIkXtSkpwWFIKFmAwfA/zaZAbNouIWpjSqwOANg8LiexwLxBxgPjvUCmhUvRBDRJfodi+tec
Dlzcx+F/yOFkJRvp82gKpuovOEeYBdZtvwHmfffmy0LPm0hNYmy01cWmh+OPd4uAqG6TtdgL4PYw
ebdx4h3501xwqp+IT+ne2JIC1soZR95K6zLwoi1Mizk/Nj+aHmlbO1odCsACdm9JB/ESJEwS39Qx
p7wbEeo7Y7YeVJj1EczbKcKvFRvnfczJmF6kLV22Oc7xt1XaAc1bEEIBtQyZ7Z7rIMJS/x1l4M4h
IyryZy0Ng6o0foBatKv+K8lQzlO0jT4V2EqSk9Tg5Cvcc5aAHDD0u7es8BmecguRGsqKbYYGXeMg
5fMkLjSPxjSvBag35pOa6wJ9FbY3yBZ48q7ZGET2Q94qhL7oGaWJpFFJfOCbMgULI8SGtjV8C7vW
tFf5/PZPYLd/zoVIMeq4jee4CV5jE6LgR3KmiC07y1nWCSqLAlf+77vcd0P6Pi3yPI/pljEGWGPF
/GHhBomfOtd0LCUdjgmQXLB/SN89NBQcAMwsZTRpyAIl0EcXt4Qh8qQ6A/vilKgLTlZdPh0eTq1e
yIvgtG3cdL9jOhiO1uW/LQCuJfHE5oPfsKHQrLNbE3cawb42hy4KfzczK669Ok+zn1qIdoaTTYPX
6gz0q+ad2Akpoj8gJTOtmlNisZYihfk1mpYR3PV/RnkBp5VJwDcWpqsY2jjiPPixNJu4WRm9hft+
zLT23YY88KDVaThWzneJ80cR1BockDiqbdfiiDAw2eGnccHTYBuaoR8Sx1q789uTgmKYXCjJmpTc
agXK999ezGkRsL3+JFUepCjJuOrqKqFOJyWiEfffESukGX7Rx1MzgCd1lSjgyCmwZDEzfusbk292
ZOomXGA/28tsfpOMamR1sX9l2Tb7Hgfgxok3zDZxULSHsE4fSxkKgH8pNkb6kLRWgvzrI+RQ+WRZ
cddOoYPxquXLD6D9BIBIS8bXGdR04GnbMf2N1k9xrQeTO7Uv1ezy9c+KPCku32W4E47FePc+5Pms
jovk6Jn1Mr1PFdE003GOsMOnsPvFEB4I3IXjRQUv20p0yIRmspZrkXLiP3EdTjrb15jxAUO/g7Ni
FxAzjwXLJvmsnfZX/TYljw5ZCUpYUijJ1YDybEG5YyNIkTWrRREuUZrtBTFi/caw9R+4QGKKvmTt
B8xDmXPRDJ6Q6FlB1csCCOQQpTSe8h1xtmOUzCGttfz9oQpc27NOvz+o3Zr08rFVbG4YPxS/0xSX
Ad7sbwtqVzePUxVIyYpMLpMCJvs8zBZisLjS8Jeh1mb2vTGvXFJlA1vMC1Ei7a05mhpi8pFZExlc
7DMHbmIGQVuAhuIV9SWDa6HwpeBqqDLH/bpieqJ03/ruxpOXltXOfz6upro60kXy+yZyJVbM4USw
u4vr8z1QQj37fXKD2ZIDb1XeJlyvPz8O9NC09phhOSRss3OigC7plWBt2SZ7/WdRAo+XSkEfxybd
vI8zYQd5j6u309a2jL0fITa2xIejnP+Ll5UBXtsbLReGi7BcvQ0LqKo9Kb19IgAwpU+6DjFwKINZ
okMuABMOap4Ec3YSxmeFPRnWPH7y9S95FJwX4R6AeeadREU4rBBiVDTHuWT8OFpEWi55uqK/QmlR
0V3M3ekLjuyX50C6SHirT3t/qmxRX/u7pUfd1t/vGj3C1HvHNQypfOjGK6UnBRnbcSxHvZ7CCfGT
SIswfFAxk0jwM5oNLcE7EmXrYwWPJakC2Ebw2wu5hhCTf0tpS/6NPEr5Ljd7+ficYLbaUttt62Ak
7wAmSCnNGT2TBoBG7ov4gsL6VJQNBJYSxlVe5pGdeXzHt2TS+aQMjbmYgTXIW1HJe1KapnoxZ1Om
NvejkeKkQE0HZ6XCnt9sl4UQMYrKqWhwfeJpc3Ojn62sRS18/4XKpNdPYz8OhuikVM/GG0RSSsUK
mmgpvzawbAEl0JakFCccq9jRr9iIjlzF0CLnjslwuYgCPG53pMPVri62c8zrPn1BNEbz6rYoR6Ae
PSwfMOvlMG1p9EdnneydsO3K8SFpqwQNSNkFa1DD51T2ioE2CxbWHZE2weS9Nc+ip48R6euwEvc5
EV7KJlwGFFiA/k5geuuopWe1S/En3FHTR+A+GGVpVchJlCydPP0FutWQbzGdJzH25vF4sc0rP2OV
7X1ACjRURADm5uydyy9BJFTNHNk+yZou1If5YHSAUt3mFPgN2hfstQmhWRwUPZ7TxppBvKJHFc/0
JuJ6cbwfIW1zk+4p9Eorqf5c9xaeqU23RSOghbRc/glkT0Li/B2H9kguZYm5cH9+6ycSSremd8GE
Sx4RfCmwqgMYhS6/bp+vezB9yfaXjj9tUFSfhQliBTgr8Q3N5dtsphdF2aaeFOqFcMA0CAv03zTd
NzJcEZmKscyqZh5YksVk8okY0iAl/au0Zy+fgt9dEeukXfUHQslrfwLe4kv3854d26BQNMsegVJW
QbyNxl3E5QInjmsd+YzC2hVOgUlY3pcqP0KcZdxGuvB2HovXPZTWdiEKpqIWRC+U2EI+xySA3DJd
2iO6uEsGpN4Aw9NBEv5uB/qOZtzj54NMoXq2BTYwo3ELEctkPwBrVVZswPeXrfy5jON77sQX4GpM
rm0bTQ7E+ZWJwnp9bIzEdTwBk9wtJOt76ql51NqeIDGl+sKF7opQq1HkUOZWpC8Z1PDmmGumnFjH
HLFTG4Z18eFkk1VqA3dt9atDi8BR6f+RG3wWq5lDv6dXm9oxdKaaauwnwussK9U/fRVHG0+WHi0d
LgFJ7kQkjllLzTxMUu02h6X32qLctgQ1poVb5kOLIEsmXxLec4EbrtIOjmxFoikoFxHVWy3Uyvf0
TWBAiowZ6s9ex5vML8CA7lQ+rQyA8ER/xhpGftmA1NBsmwmGGUg0N/9i07Df5kQIjilAhFYazdFE
HQ6UNTt2T6GP3CLMx8/qEPCh9NV1f+PLGIcn3Q3omepZW3KJYrfikNFX0ItI/xV371yUSeQ4nBN1
UChlXKh0wVZ6pLWLCRzAz+6qwpF2CwssajMQdvves3jv1np2tuNXXqeFQ+rykqSX5fqXyB8GxUOW
rixOZKJdrV3uZHTW004zSeSHywhX9UxDaAt9OFrJmwTD7aXduIiHZrJZyhJs0eNZfXi+bVfz/cER
g0sWb1qWyoHigtP4eqdCyhnFC+Hkivnk4uWywLCxFXodsC8folzWxYNJblbjQHU05jgcbXr3jL2C
wGr66XM77okR47xGVViR7gNjnADk8VCd/A/v27JKwSbfha2bCwe+pCh/1gqUwuJvZFMb5c3bvq5T
uYXccIiiCw1Im/nOBUwdyHY/4jn8XW1dCbR0gp34tpVYxWcP5dDAsaG0eBj2a09SRLbDpusrlz90
3GSwNx2CDA3zb5nLC5viluZMdqsV6OIhQs6p7YZx1hQGu7WUQWd0Me3H675fPUFWufdbJkUK2Thj
+8TA9aJwRKZYSTztQtCkx5nbUMPmweD3xO8wBqfG8dGMcQrA7CqM51OFJ4oHVz4dLVKixWQA2Ach
U40zRdoYu7HxJ1EXJZ9r69PyhbmhkivOdPHF9C9BH/21T5D/blbmvEWMPI5aSzzt4KYF+WEx4iOL
8JtGK/8mxu7U0CofIW+aVSDcnr0rS4AaHi6O/2mFH2bD9AJA4Grp4L9fig/rbkp6RBe8YkcjSsR4
BDo06HEuZ4WPZMrzQGTT9iV98zh7XHleAZ6l0lgTag4+87aKTnuj6yYalOUSfcECmmOp7OpKgOYe
hFLlfPNosUVCCzgga9986hz2ZJ+JjJ4DbpU96Qj2ubgfVtpLR365bSf7SUD5kLOiqHuTyQO2LRCo
a3hnFyernlMJfhl9q3lExQl7agCWpu3liTH0DAPe/LVZFK/zmQtcpcgidq4lLNCI+kHDYEvvypQC
IGBpOm/aS0gynAdG+UNYoI8598DZruma/3RYjqGSuupeIbN25LPDsltnASSt7qwGE5xp5dGZtm7a
D3wOIy4MFCNjI7GucEBClMHk0qXAMkoYrq+0nTN0ryi1eBZQMmBALle0lxPwB3qVvng6h0oyZUbz
JxzvKSSK2AAoy2czHfhiFAkk4shTN40puRnG/aeEfkB6e4/e1jP9QOCwb8P8NU0TExxoJulrigzw
Qeg8oQc8Hd6XiX344lQeyLWRUnYy28iWr34yt3AeaJ4yFmgKdfb6BgEka5mxoIOsMgVwM7ch5ODw
7bjRrZonM7xdgAhvnLhw1rndvBVnThR2huP/psaj0h05hU+ttuPxz5rfzLCodbGq/U6EVKMTA27X
gErYg6i/et7S0z84h/aHF5zm3LAy8tJw7AaGly6YVoKD8rZM1JJeyonz/8xNPW6spDNcUSDYXpa+
EQI5Yewbl2si0YC+vk19FZBVGQ3jz4hltu0Fw4dhVKqzToBsnWgIU3oXv0q5QJ6GSLRVGwG1nNIy
BVVa8DmfMQFJp8aatPZNn7RuPfDVp1dMfWS70FpgvOgBKsDgEkntJbvnxNGT+S8r4OJaCz+3RVvh
lkop7lEf5ZVnoOnvKzlx7xSee7gByF3y8L+kEOzbVcMz/Jr88FGbcLl9MsnSlxPVMZwpWY/IN00e
TrfHaz+008+bDaj8NqFNCEJO/ahseUVzUP++RdJVojXHCJ2r2LP0aCZACGCHu5KLr9XYzQmis/DX
pya0w1+UlpZ7jpNouAUQw6M532Q7wmNJU7M3SwWXRh0Ywt/T6MGnBqTfDMzLvPd4xw29s9gJFxjZ
fwKsvyABsj/yCpAO8WE1HzQ97r2oVFxwVsQZxQ2VVlFfmVQpPCHpmDO9kTsNq84cqRQn4kCrewC0
jZvKSGIohhJ5vn0nFtBxUAnvxLghLdqpDXXda2GpohdrUrSeU5qe0VRsgZivnhJxHGCXkgPCimXj
m5iDtQhgBLjjR86EndL+Yrl5oFxST/u0ZX/b/MvRDhkBI5H6LmNS68H0Km7jw/qyGy24sG7vOSlM
XvvkX4mAA2t2hGipmW8KO+6sm2cj4sYSHM6PoQSp28AtjeUNie5RhchES9xU9iBvvmgMF0+XVW0I
j2upzMOk65svktW/dxc/Es4l5W/ZC2SH4XdlVSORVd6sKtTwxQF80r5YuYMIOJo668MVuz5xBGL2
XoE0WlrB1+vTz6crFvouM/klpZvN6jXV7QbCAx0BZ3R0qI9ANMNlvGX0sqbLSjlWSNxwVxiF2zLV
NZsjPotyHqBu7l+U1shXgbtC7Ae5fugNfiHTS3TR91X+/fZsRHVIwOfsHjd0t3/mITfGYJOROaI0
mlQ5jyhIzbZd/pSNMOXldbnIOUrpLjQZ35yEfE5/f6RFlIGRAw01B04rOD+CFKrgfG8+ZnMRT76x
XGTTOm95+axJjJsCrM0OQBFYc2+O3xrMVbjeyziMoN95Iiq9j4Pdq42dGEpi0exDAGPDcSDQyqy4
0basrqIhHQBATsyeSscbMt9j/0YROnojjIUQFZfSw5o2tD5OVWNlNAZU+yhL6m6eaiHNepXHYQVE
nkAmPUhovigckA9kj0orkKUKi2B09qhG9tb/ovNvaEtXsbVZlwPEpzfsMuOKR4Bp4wfkjBSJWcST
k6hlQUjZ+fcuEJt+lPqKmGTPow9PVpKKY+NILsIDtGojglxH4xJdC8sP07OR8M/bW1W6pAbvhsN2
u/lRN2B2pUqDgSgZMqSxVKvIxrUFbLahPU5qkuLtDxGNWeLfAikS0EetC1y4CFkxUOXeRcPRZK+Z
xx3rwyz6cdbdLVU1+ShDpEawxh0YDN6fcc6+74ANbvJgNIOa65xNHDmsFru/8yBgdfURbuMXbodQ
ON+5NSJbM6ljv2q2+UpSA2d1cuAzhAHUgNAce47GihbyePsbnndm0DoXRHMorHUDD5OqyMn6GJQp
/GCiMRaCMjpyIXZO7iPIphFMCdnFsTzl0bTXniHSP0B6mPMhrJ4vKJNrG5hUb4/V8ZYCpKhr0ovK
uBOr935TMyCy+vcrSvYoMAKGIIEdrRrsCOP4GRfybOar4GuxexrAiGvDrTPhcNMNB/k0RX+r3HOV
KRAPx0su8rW7GjhZ3XhgTqC9Um9QDEUhEX+7eqxfdFFMOd28nGl+VgRx9LTS/l8WGZqc8cokAoWA
P+qv59SG446EtS5LUjmCyco5Xr9Ak8tsBCK0WEuQeo3h3w38EC4xC8eSm7q/w77ZA2kTMGZCw42B
+rYjQNCNsWQIRX3+Uv/hYRdRX3OP3SalU6/17GLuS7nrEuBo4X/f7IrGObgLdfccMOf8nGQ2P4NS
I/HPOW4Rq5prSz+kJ/mvc85r3jfRR7azplCf3nCxieAOBXDPepmHVHIFlt68UGaRThZtLQgjGBaS
JoAl0wkbSQFj6V5IOV9Xm1ITxOM+2LdVMf8ixV9aYdgV1uElkDI1Y8y9HeoxaE+8UJrNz8AExPAM
jVs2gsvn05BC1HgzxRGdfuhira+d5UmQL52HN7lEjRdwiGzC7ytrnCKx/aVOI8AvZQOrMElYCexu
JOTHPB/PE25CInrIy0oxv7NoW61Gpk9sk+2HxLlYgzvo82jF9pNFETUIZ55W7wbXWKZY7dhlsNyV
36bAKrpOxPUoeiTXMN6rBd+kSkDgB8ZgC/ysI4ew4S3KTozTPUmQ14CWkvxzrKoIpz8/8EbuMqET
AxHy9HfMe7CsarKuCNxWTo059QVZVFdkBCYMtpWWIPOuG98qv2obYEGcqM63dd7GUDUSyO+VHQ9l
OrZFWgwjHw2sOgbLMPo1WR0q4CVPzWsYkJl6wYUUviL1zVJvx8GaTRMjZrnOq2eTu7E0YBzC5a7z
z1arDKKyCyZUK+Bokbsmh4cOue+6TKyMi49FQmnwm9LfktwMvMRbptq1OfH3j28Eh0HCPX+50FwD
bxRU8ZUr5LzpE9b32MNi1pQaXKt1YD3ytrakOYnMyUO8ulUtn95NomkcJj601LFDVpbpdFAplhwc
Dul/cKzh4zo/RqNRs5npmkJTWWzSoIopMoJXPZXlEPd3UEA0HQIvaN8KqZ2200jl7J3uq3lzl0T4
ij/9troHIg5RdWUaIvsPqBE3Hhf8SshJJrRSucP189qsYcsnC1krxvnKiAYzhcmjfX2xNsKznSHw
bS17rEIJfAXYud3RipWJR4LEsrWWiI3SOv4kU/LZvWXZgtq87k1GycNCOKB8FeD8Pt8N0htsz7Nd
APHXJGjvz1PUVFwsGKOokuy46ND4O/vBwVhLM1gvyqaJsFunPobZO9y15W49h4v0N4PgKXrB1Oah
E10aO9ATc8k9VPVhMuKa5Acmo/I/6P9kfhIJiV6UkiC2xM2Kjr/wCeavJ7Zfxe0vBpK/Zu4ucw4l
9v0cozQQnWJGwO/Y4XUgiwhnJ+rr0zjStY60CWaEap1QLtHeYpluE6Ken4y4GKtF8fvzsitrJskJ
4x589VW0ihKUhiJx5goUfsaOMWYQ0SyYaF57/+x4SGlpJxnU41CrUQiNbA/t7rFg2g9SL3TWmWak
VF0txNAaA+Uf2GGJ7PCj3X6gENWHzy0cDp9k2L+GvClMn8AW9k7oFgQnQI2kKP4sdi37feP6tYLI
cABIbUFNo2J7RpsxTZ7By7S5Mt494zE9hjo0Sg0xudbWLFV8IM0CyZ/NCZfhncB6EG+dgMubfSfs
ySvr8zFd2L7uug4i9OVl4UN1/9GLpSIf0oIF/cXVY/cookMb6TeTL8Y1Pxjz0Ubsp8Qn8XOU4oti
qHhW2RvcBsr/IbSLi7+LBP0rSEwGQbqgKEMuR3ecg4GoPbs4vWY+t81lKjWY5hfANT7O2Kj6SWvD
OWSiL0Pz9uD0JJKkvCenWVBbklFuDO8STJMynRtzH14axsYfuJ1J+nW8V6UknCFCasvw9YoPvQn/
Yzjvg7BqSjMp7d/k8Nk/rXrojdfkFIBDyMjdEpx77I5DLC0XxOmf98dAJZu0ozQj0HebEZMZUy0u
wGEU87plp5/mgAsy3CaYCgUe4WR54Ehjw+cVlpXljmuPHzo/Fg+iGbsHTULwk8O/IfyZQddg9mu3
0df8ZJ9AMqPQjiQxisxtW0YLcH73HOrqhoe7oEONyDTwOb5KrvKKO68m6gy+RS5feGqHzkBqv+4J
CX6kymsjAM+TMzScq91xwLaXSeI4ZAynQ1391gQQgpvjM2rXupO+q57ikoh0GLP1kzjrt4ywYpln
nXBaoANdCnLjiQZ2v+Q33w0p/wezlfbUZpAkEVEf0XDIP6rVkn7UvuAx619ZsP66NYWnmnluOr/v
D+RT1LTKgt8E7pHwwhb4TJBaNS2rkT+kqRmQtGtPBi0+iY56UgD3dgcUcCQTg9gM6+p5sKOqTciQ
xhjRxj05rbzvD3gs8fQaAiocPWTBPN9IaqPIs8gkfdRMHwCUy7WHwXB1fcQOcY2iXaMPilaEi2bG
JjddkDMcvyLZAKI/x4A6Y7pjTLOarq0P1T750xTm1sdSomUDaec/yYBORxxEkn94jYIHe+RC0hpc
gJp/RdLk0ZgX1SxcrLqjoX3nolY4HCBb1wrHmNj6Be9g7hrU/sUeTxAbcQ+qSw1bFELycBkLJqPP
NSblDYyIipHvVdPjja1z2xCMsgshcX4HQk0vfb53p94/ny6c6L6yXMD3U9mT/MFT+2CmuAz68ZiD
89NcfiXY2BWDrE2bKddZfTNIuRoaIPjy4550DG3gWbzhnUeZLJ5IouAKT6ztjGgcrzBIPVj5V0xK
lJDL58j/sP5suPE0fA38KuBc0qaRzdV7IoMWQdis4GGdWbtKpkgPKhESDdP9ENp4HgDiOSun051Y
OdpyDtpslE08zjpP2uSxBZem8K+sxGIsJb8tPVs866XwZwtRMfcaku/yW41P9H8GhR5SGGG+itep
6flATpkCFC81vVqhYA+3aizyxjjU9et/6hdVcogUcoTk60aa8XUmw9rB3yI5tgAu3IlxWWxfxZrR
MCR5hLFkdm4Hq1ejBVIqui5LjcgIwnkO1hFlV6tQTzoTKEfroRrjitDJ1jKpFeU62jcdGfi2jkdX
+MP4yRzBYJ3KHRT2269bMEJpLAxqGh1JWMyUjPNIfWDwNMJYBDYv/8vlDkA9PlCElTYbqEBZ96OY
ry/rhFEYL6WrLUi0ocmswTNWBGY2c4IhCCwMbfx8amdEz9PCGuSPAEeBKMEzzM3oYdSuSJIapK7E
AYmk7SaxDnn9myHTigjNjt1/Z63peiPYyfLEP3hyXIfXycQwcfqMsTX/M9wkFEYyZl96ch3wCp0/
2nd+WpcKhR9FycfDd9WvhAkM43Qs0RyToPeI4uyrlVISuzuXcAdy2VS5BT9IKi6ekIZFNRkhawYd
wDi/OE7ZHWAD5/WyoTY8Fxs6S2LSRB4TPiJTpGDmn5Z3SL/VTHOzMo/rYwVwdzU4tJ/ALfIOSlvq
s2NUGXjLERFLBjzM9bnv2aOwxrEXis9VAPEsHQza5wUsOzlL7VAZ34wH1FqErmjBO9IwFPXIn8/Q
+EU5vWlXDjHwZO7HjmPmuT2QMT8S7H/5UvCBdtc1eHKp2QoOOIRlmzwVWNBgKK9TQG8x7jU6xy3Y
f7B5EZwA0GI1wIXqja4NP1V+L03gfbhHHhEYwuP/mucWX0a5c6J3NY2F9v4yPqBcEum4t2A29SLf
E6wxeqnDOaVFD33vCa7kRZRJRAQHpxQednKK/4e52d/PfdpdLojOyLXCvG8gCldK89PmSWQHv+XP
qyeGs9RZl2qkkuGa554lr2h8UrgDWiCh4JQWgvGz9Ampwl0o956nf2wSpXi3wR5dSMHldvDCFnlj
Pn89QUJrMQyK9krqPSXyTu4GOuqPKpK77QDt420XLVJwDjJUBnU1cg2Skme5J3T4b35BKkrHyVuT
Vk5c00TsqwtmrLu0dXuNIKwDn3XcoKimROAeR2lioC8AKNysbRu7ECA7Il/jmWpERYuYW2SLJD1h
KKAaf7nG2KNn0Pdkb3JROM3n1W/oQy2KOwt/V5mWS2bo/LvIeLVVswjhtoPdUaxyn4PlMU1IbFXD
tPYQA6LRWwkEslfepSBXJfbPdVPKJ8FMGTMhJonmaauFBcdbGYPNaYHnkNTQRZsmgX4zZd5WnNcx
7vPvjwi6E9uUVsdWQ/zzMdqiNsTDo6fz9SQ6l3WfpFyLnHcV7Zm9BDXcyXMugOGndwIjwrwdv14o
1+kaszdN4tlKUxEztBvEwZQuzAYKk15dq9NUbzj8qgtfEfVe9Kg25+JXx7oaE/UC7NIs2WHMXCsY
iAClMFfAHkVs27P/LufAvo9ADDVRIldf1c39YGBdTWfYsjIZd8bouq9DvIiXpVPrXN01RNftTmhE
45ChHCFiBZ62XwNxLaZLvDm6fyLX8of6cKDXe8HRg/y7YNCZM940kMJMGQx+gnZbRBQunK0M7wK4
64ccbpCOpsShXw/wm3WzWO2H5n1j/a8snbPPxTkCKJ+uZNZAAUjspEf+abfAhPK64pQSC0FaM9iP
LywtOzVjYHM0EW2i/egEctDUG6pB7wgr8HueErhvuSVPhzBpZlL7baFzWt4wB4qPTNmvAElwRWpA
/798FiPjLMyA++adUhaaMAKhp7/SbrXc2mFhdcknMUzQFiZ9Qw3KqcM9J/05C7IEzPvzDY2mdOVA
8P2+VuYKPgzn/l2nXtpAqkne0YtksdwICuQtV2guWAwvaLDfAmT0D7TOVs2/swfQNz67u/GphNsy
vNlqBiHT45soTXyl7VTeagsYuXdQ0DfCOGu5OrIpBXyYcjrSZp3/n+baPyEWFBN+QNFcpK1dhGhT
HAKMvqOWadZUEnV00thAoiH+mAB0S0eL4sB45MDZq9wMdGlCvz3G8A3PFZ9m/GuZB3d5DO8ec66V
e7JxckSL+p7KXVi7xXFMaqsVB9A8V6ZB+dkBw7s/hy9JYcLp/XtBTRZCPGHnU7OyTKc9akaA7nu0
NtxHYnwKgshujosbBWlOw7RIQTEeD+HxkoUIfVmnx2LDcyDwQnDrJbJ5NjyTHf4M3aQtOsw3MF3z
4T0pBv3YHxGKm+SqPwrS7kWnj780kkqrgc7S6qk8X8NfN+RJhm7MF8S6nfOn+NQ/UJKWYQ/UYoUs
jMvT3V6IOOPMHTB2aTg7iu9ykSccZlly8886mduYPBSPMZMj9S30yRPvu19/lmBMPx358uHuXRru
3P1Uxv4rxT+Irb8J2IWw8GFZMS8k0PQOY0Ki/HfA8WIZ2dUUCIAL06SM60M9RBCa2FLaAu9Avjwi
l2wJGb4BjHP7KuN3Gqymta76wU6iCt0Ao1f7kFpiOVDmmu/F7T4/8GITzcqzjOiVQ1g+q48hKQem
M1vwsebnBkfTF9kuThF0/AFAujYZmJ14AWDybCAiqSXmkcnZYQGVpdtgq4mua2aN3pPOjy+Z7kM9
5c6Y+IR8pGev8TNHkb+UtzCDphwd5lcfHhjelZE6MlUXP4FMrZzBsQ8fAI4tDcVx2ZEzNEK0Qikh
5c28tCRb+iYEzDLLQ+557gPKsd3n7p2KC7OvbACWTZrBJFHsbAJroQLgJihUua9jCTZeNhsNepri
xjq4n0jAKeCNhlm/Ee87W+Ldotf70wF60+cuqH22Io61U6Oy3AqT3yftxJ1PJy99MBC7TLcyw2fO
rh3VjuVinoDTP4+xtLRqaXE9C0FuboN98Olmosqdm7X2Wtn7TNNNnv1ulL/bj7HUptGyysJuyLoo
M/4MCxsIUhZBsH7sKx//9cqGDL1dLfTUUcI4K9sZZhQFKAIMfHRURia4TRH5POWOjx5CMPLXyy3P
qYUeAvXpzuY/RYz8z3/UQC9IBtN7hFjqcD8vcyKfwkpRAkyJ1xFWjmWK5f/+8EQSyLhuHQaImcYI
H+i9qrkkWG8pGeig+2gPx4hr5WvDG4EFSEJko2wp1250zZl4/hmGIOlN3YNmSvmi2bwbhKCFEuu/
yiBh/pTDaLw09aCtRb83pM6SfTM0UknnG52Iqmi0ORYh21Y7XIGCCeL1hjFBbtBnkDB6cR3Xwfke
ZiIOCPY0o4yl7JC16uyri+cBDl0KmVQ2B9R7vaJW2+Tt9X5OhfXyh0reTMfzTnAEJWri+eM34cu6
XGyGrf0QxqnuRuwyuOjt9vI4eBFt0Sj/vEnvjAhEWbTMqo4rk3oq7Cl7sRaYXZ95mYAfsa8XmX98
2mIMm4JqSezJ8sc/2Fy08YhhXwvAhEAhuuYIco1FvAc0MKTSfcsFzY+I6/8EJW6qwdzL05LTIqB+
GQ91E4f7dr7CWt7l5RmfVhV8lny33egdfocyZ/3AMOAGD8jsTu5yetiXFOMrNGzsdwUvmzjAXI/R
TeqClsb3n9JiPEwz9wTZH7sx5UaOzEWPrzJ/zl7Zm35jYB982esn/Zn/wI9FybBNbtJFcA/Rzokw
hqdL63iW1jrp2o69zVnz51NiSyrPM5AH2CfXqT/5asQs3aO/iRgLZyzzWVkKVsbZn7kpLmAN0vJg
XM2leGACEFhjbLSvL6Vf8Rrq0c1QMzg9M4x1rGVDt+r+53AM3eOSj6LUqa3syc3yYsshKPKr4Rw6
XOeTSchldjILjBO47Hk6Gl5CoDJegHTxqeeZ9xj96GWVfV9GssL7gu+/b/EjUvfnC1CkF9YksDTR
af6kfvdV0RlZDUz+FGHip3ZycgTUFF0XNqTT2TNbPLpjzQQD6K/jv00HmCievZhuxa6KLWzrfWb6
0nJeef/luc72eijHf2WlWxSCdMheEkyL2gVTPZP1gGIpLcJzFt2Ajcit0pWNH7thDuSc7Jl6/Lno
9C/gvYVgd9Ut5nEfHlR4K+djDGYv0lIkFjAt3/xwkVMDgXuh79/RQsDv9FPZDhXrbTPtP2wRz7oP
+eIHLODMlvm6rURODJZ4RIU3uo1rupKHSHV27HWJl4jHzHpHyR6rf1ozA3owe1qvmd6alVEJNiYV
Q0AG9Rpa5JdTQrIOWLMwyq4Uf+8c1pRMIfSZcDd6d7ps3mUet/K1Pa6WJ6lRAXC7BUUcQ6cR6kSR
x6r5r2c+P09VVIYtjfbr20P4gBCVWZDvqMOX33smp+V2EUaYAZ4L0061B1UoqH2M6csTnohYIvK2
OZiAy1OV2mfYDC8F7Z3/1Eorr+qBQo/haPLMSS5MHLCU3rovpwsIaFlrC6MVtWbBv7Bf/3jJHQ8a
X1NTcGLakGjNdlzDwwPC1YA5JpjRwyKsest3ARXqxfrLJCkIXnUC4ZR996zMThXa81XF2X4z7wGQ
B99jwqmlw6/nBmvDGvzvg3MYMITSN+xfV3SC/jfxNmzIWsAfejmkl9OUXgiufG8idq6doyty/pGU
BoFA6nfxAIbpahy/A+JLvzJiarSU64fC/P+R3GUeUs3SEIVIB25hJUnZsG+ieQUtLC1BGTtXLWLk
HfgHYMOMRls/JS79eyn8BZ9JS9bB5zRcOH0WME4DNvxS0X8eCXakk0F3/dY3KjPoQyjJRIdW1BL/
lgt3GDD5kCC68QFic6A9FbM/Gxltzo3YT8n45S8GYMChBluJbANG7PvOJjh7bf+W3FnQ8nFbQP8J
/IPdRAhcuruagx90eNEWiWgkbtfDXgIYVYJSbnHVSgkjXRDwN6w94sosswZOFvY/5k1DGtG/M/58
B8npkb79svPgIT3Gia6h71gAJtVZBEWI0FfD3m7DneCiYKpDfWmOEobMjVZDqbPUUBHEgx7IL68r
ZRncI7IQ0D9Eo3A2yKAZPnBR319Zy2CeS9Vi+583+8T4S/wpjaAGkwbvPamObcibw36Bzwv3et3e
MSaz+eYtHyn21S+CgHVW39uwvfPxOR8rj8E3D0Ut6pK/hWjypRToH+OkTKeQDz1SQVVECJ5lRqp6
7vxsp4DsOejNtG1MKbo9k1X4uUblwcTtNVbl6lin82QzjQwtGJRPXu9UmLBw1Wq5h/oqa3CBBBsM
Q8nQ5Kt6/KM4Ds4XcOBQzsd4FI7R6JBtnnG6cogHyJEfkl04rsTgHJaeEouN/AkIg5GVMCkdBv7b
GglutuNqrZm65htI2DIk5G0KanKXFy4I9N5iUN/OEs0uKtBk42sf6borZke1l087XQJ/jVEozMX7
8fff1vbZmN4IUD55h/818DzHM+ADem5PH1gz60v3FlZnCcXXGxPJOvaQDs/mMGvfi0XiW9VByOPs
2Rra1ciC+V3TrHFoL5+GIf2TeVbbn9cbQ1ElAYcN6bJrNEIoSPBbwIFxZwPCe9DS2rd0TX9nF5MS
Mqvk3zk4hNJ+5zeXr8D9hnpqH6s5Oyd0vyZXI5Qgk6D49Khmye7y5H1gl9nJXC4PP7+IG/girSDd
xsz2KHGq3z8e30UZXry2WTSvIWcOkxLy4voaURrr9XdZpiYMlJFWLM8KgQhkG90HOb0rvHH6M1eX
qvUc0mfaLvYR4d+3mzh1Bl3eTE7Mn4BMcrl6c7WsCzdvsZo5ayz7E9CBQ7IRXYGBIuiX9JWndmKw
fQOA0BLLMHxEwrY6Ic8LfBQD+Bx4mV82cP5av3OLd9+plFwqIr1yKYon0O97pwW8Wgef1DTyXRlo
3pBcVxdq/XV7+r/Sy5RYnLo+N9z6E9ADTmbrthRcHxCYbT4Mzs5jzoEX78+aN+EkX3tS99NWJdeU
4csakAy0t4QURPqqG1X9wbc+EaVHi+5CkixFvANa/1hmG77pHjfeLF62DHfkSRTy0KgjFE/d09CV
4nK0tbB4M5clRvDvyDnD6qRgdcpVgwyFG6If4egX+3ccvptMFUlTXC8sVfQuRqKLy4SNiJD6ZRU/
uIwYDc3xuZUWp4MVbDTItvBQrvHv0KvN8tqXYlTgtG0ObsZQ1I3fplMMYUj6ATgF3eHw6U2QE6qy
1GtBnpnL91IIXzCOiuz5E2Vk06fqLzXgmWO02BLI+gzptaGpgIFWV1+1hcL5BpHvB2TKGSZUkubl
c8qOca+mIp354RPvv+KouYjIkqOj1uV2P9cRrLkvQ/+UFwJCW+jk90oSrgtPay81WU9mFpk/nZgm
WN29kVReJ7hnmI31LbkyktO5pwAnfAwZLejX8NQ8cPr6i9QQD8oY/Hi3OQuTvsmMyLPXYpu5a8Ux
FlIwluK2a0plHxx/r+Mj7suLFfp8ohuU5NVmjy99JrBMT0L2O3oVyyruEKgAehmsKvDyqtgY6BR+
UGoIpf0S+zo1FsL9K8xc97DtC5AnuCwggr53Jz8iOUgZzzPjLeimMhgwtG4QocPVbKbMRAK1BtvW
XkFzuPHwZQul/RwsdYyV3GwKUd/j0Gw8UjpxknLm/+dNiFmYtv0y09vKQMY3lCyi12FBj8FTBvMv
J4IgXXFQvxIKRRBIus6KhXN8OrYA9X/ff1WAPgajkRC4NgK954gJejCBrg1EkTxlzwE/adgpSnY3
3lISRXQPnzdyOl2pJXZ7O1TcMx4xqTsasg/CxM2Ri0O7QsdRagvavr1qt2Bn3J9wuU6fiHuALqxU
73hCIyL/UwWgR4jdtZ9DVy4kyRN539LsmRfGa1u1dnmtJeNSoKbhrryxofl/96lSj872OTnZXIBR
3TZOUXIpOrbJV5LQLpKkRBYdxj3cFB3EE9pgQHMVrgCPB0YWTOfsQVguLN3HAXRMzjv31nWhpBd0
7WY60VImJ0YEJh0/Vh6UfPIzp66YG/+H0VQ7OD2hSiOcis4PF7AmaSjgaiXPE4fql89I9oLHu5zc
TUYHthz6V6CFQeIK7/REOOfIqNG+I9E1U8MARec1JkExLwcDDR6druP9AU38SsF9DE/GoPz5a493
NLRP1JG6hggifJwyikDRhC+wDarBPaoq+eS95QYgRA45D5LUngiK+i173ntPVMlqLrFBIeVCm/pl
PmHW07VEaLW8LfsUCQvGyfZakoiVgl/+K+Dk4CIStwsRYYfkmKA8bg10qfaSK7G01i5LsBHDLeDG
PL48l8l4jAcEgoJIi0IbD51EC+ikrbT+r0sh2/GocMN8R5RumkmHtIMHanw3LSZiw6VTUTWjrWWX
RlIxlLun5DPFVIX++fnEkNigXIdwI94BTwoiAE3KOcQOcZ2KCwmVTM+i0YtBbf7EhRGVaU9IYF3Y
VY4WndAipuCKy/g6HoQ9bB7RDSqKz6VG3Y4ZUsx5AqrKlOMsfOY6p5gasX0Dcgq1iMf94XBi0er5
qHR75IJoxG3f+l1gcHZFx5M93MehtdiNi7cLPAdRxZWNkqC9i9JX1Jld3Cv8J/TzoTP+vcLK2k7F
5uwlxveZ2k/CA5Y02zJwpHBmy/HwcnoNkL9U2fsiN+U+MfqpdD/MxZaXMGGx/63Pb0In4t7zzXfQ
7jhHNVdZ+lYsJsF1SY0S4GNNjoi+UiJ9PEyN33fxTK5y0pGYjPu6tOsGlegs6B2NTZHECgLtAwSk
yKUkJP4jpYy2k6PJU7b+8XYKjkYX5bCgPJkfKX4ipyfg4dvLhTS/Vr6gFOckU+1+xnTXUHA1Uy6Z
PGmSrP6Db/GOMK0pgW4Ejay3hhNMcN2P0O7/52uOfG0j+93P5tgxWSxUXZ/Bdx+yu8hwcfHsCYiR
K+MAhUU28Woruu+6fEgzxhlbJkdwvTvbhUs8HPXAobWqMwVpQf8p3VXEGuh6UIQwLl4U1EQpb73P
2k8mA1j4Q50FwRJym9MutFe6mde5v9bbm904a6akgUKQkIi5hacwtJsfD1GPqzk4EcCsvcddGf5b
nI8fVUMhq/tsk7MYaxLd1znJL+tFvPtKFDvP8DBAKUZA2aPfYjTBayj8BzaRhNP3X2VNPT5rNN6e
m6mANhoZXo3SKSS+Pbdnt1SGadM6dbj+BZqBkLhxHmN6RfNgMC62h7P2nHGH0oYw00OQtYI0Nfm9
C+iQFPiGNIAGspYtQK6c358hjF3VCNGjCQedsVM5uxjn7KNt21FH8fQySDO4zWyrLR0w6r1D0AWs
dUNlbHzyoBv6hik655LzfWg6zUtmr0G5cweQ4ia4SneAZQExU1Bpe3K7CMXvNhtPqS0crsLkUNvs
hySBvaKEpYREppCQUd+vzBteAHSwX6s43ZYNxvz3PBE9iooJWHuP4a5jE2qpkW/sKcvODZBtTl1g
AXooUV3JFREYxK/r01qZWXde6QxLgBA+k4ruYgGJNmQtMWEsWf9fZoE/92JGBbfwLc1gF+LZSp3+
Kij45+thyr4rzjEACZtfU9Pr+grY5rXNkmvSKI+1nhy/139ajVRJTDIXyJ6g/kLStwZ1bfg4hjeD
AgoNyb8IRXbT+kKhiJwFCbZW2WgopgdxblKNpbWjx0t3MxCrEmDy6vqSheHwh3EcZHhTXZ1Se6KY
2Z057n5sUG6H72hZoY8ozak2760iCMS9z2zrEpN6AEEmuiIVG4+rFoJ9Bcx3t0etzILeoh0FL5DE
n10agFr4aoeLlu06Esaoi16xl9C6xvtfUUQYAfMrvNS451wjF5L8QwOKFMED0tNaQ1P28lMLr5/1
qYAL0ISRsFaT2GIkk2nPO3u06PaXeDSUs0xzmCks1GqKM9B2bZkqEXkZo8t/uZt1KonXWMfSe9/n
tEgssP2HBATcn2CPmlIolx7hDqTbUvymWu8WW3ONZRcxH38+N+iosQcJu1pQwSBVosK2wJVF4/ba
CuFhxZo1PUtFbLtLbcW4DE2x6AE+da0RckMlkOniUgAX1M8Ep4d4s8iiDjB0unwc1MtYy3nNgWcL
rjuda1+tjJoN1iMqJzCXSENvekUsdmDubTbl7dYcdZkbdpJ/GZS2TgGK5mgeuHFFMfIz5z8vBkGE
ucBDnZ23wjcC9Yxn0AGcysYDfHrZlVlgoJaQBk1Yc/VrLrhqxEgXaSVRo8B2lMS9uJA3G3d/5rDa
0HiUjZ/706qweINvaRXG5fuWEJnCkwNKML4f0lbkvlx9okn1gasPjL3kiAaiVmaQlXuF/BNu3CYT
jfXvWcM2ljQciPU3SZQLXcNafvM5kRnZMILLZl2dGPEtmYRyx93YVt4QcYytc58ou4wf934SedDX
DvMhBKnzFBeEoi6apBNWuQxr/HHh0MYLaZHw3PxgCT5+BlpWbgbRNEB7CVQBifMwWfuYZzDSaF1K
f5GIW5XxxocARKlNr5hJIMVZfv16tmnKJKGXaCQSWxaYQx7znebMh9DCbLudq8SLt4JIBiwgAWqs
B7NcVz/GOFDRWD5wdtnrOTZrVCIX5k7/f/04/ukB8HhIF9HVQMjdE1inCBReo8NuuHrsUVlhgNA5
TJjEsg+bApn+Bt01rQsEyymFuufVI/MNffTLmGN7dmUr/GSmk1Jwzc4+O37DmwLBZQcfnd8hebm9
ByqFISJzyFFwxj9UTvt3NlJzgXpGQgY9+ovC7JigzxSHaaN22VQ4Ex/DZRvjkAW9n3Voo1Ii7lAs
NDcePXJ21KsjglRNMXiDsRl66J9nLIwE/dGqHhGY5dQ3WE91Le2HRu3ih7CQJqPWSZlIeQFaRzXj
re6DvbSdYam0rd66Le9kdXfTkmIJc/8Y/r0P6S308BWckTYL2bKjYH3KrPviTzAqviXP3gttfgts
0m1vc8nF38gQC1qiqn+9wSlPviv5MPIHF7Fi1svJvaNCAiNo36EZv+OgST6id0s5BrBhSB6tdG9c
xQEDfATAE6yYttOLUpGsFYcwRoti47aC4ShGARb7mlvHl5G1NzI0w/JsYzrol1gRnKeXmHIvzavN
/BPQY6Ee6lDEx2cQ6U7zVFGofmNP9Dy5dR+5rA0Nn/UrS2JjnglotS7uF/FflYmcxWlIBdW5OZXR
qzNPDRYF/hYEP1FyKpjULCwOw89y9L5nY/e/xjJ+/KAhCYX7hcspod8NFcWBlioO96VaaXEpYOwH
cWLEsaSJTqC68M8Zup39tldmgD2rDihkf/7tLrS+r1b65JagLHH+6v7IrG94685Bg7yadhzzZxPf
62H/DvuK5S9AlYWRlYoY1LogYTbaBRzSmEn8j+oAaUZ8k5dDjKX58LIXSbtLKMLujR+bI3f70z4O
IUsB5rRZESm2Gk5ibNiaqGNGWspaBTvpqHouQ0PLQQmioqQxhg1aDNZxpzbamr+SP0wO4rSxMSnf
pQ//KsaT4rCEtFH2hcxtASr80KQfAZkSVsRFwoMTHzf4lSeHCBY5z3JZ4lTOYFTn+y3Yt67+AOJ4
v3MELWzTnUB+5Zxs6y7J5JE7g8gFL+hBJcTsj9xBiYENKm/xFOxeV0g2VoeDFsNE96orx9c9i/C8
4Je7BZyDPfakM4Ocp1y0MQ93lXJ+FV+jdHoADkGKgMR4GGKiQFLkkBIQBmKfmQjSCXRecpIw7cXJ
OpcNbh1k/PzllFFUtVLP9wVakn8xf+NVnXWyCNlkFYgjT9yn+/MXwmE4+vS5SGFiDp23a2D4R54G
hH8emoOSaHsOy94mVY0BCq7hb1FnqEo+8+L+gONTD8FbJYsnmy9UoKoJU0EoKCLPYzfJiaSk6v2C
TLtL2x5V3gufBTrSGbue3zwG0iDanPPivlIuI30DPz72bvHEB3c9Rc4iIgX0Cg/VCJbgCJW0DWWk
t0d1pftRtywetK8uN/8p98+0E8za4yXHJ5O2egsPlNO4A8RdnbtRKe2npFamhdW0mS7yk3bv2LpK
UJdq5hRctixEdSSD8DzoTWTM3BiT8AwLVw2kOC5ki225F6spq1DcunoXD6FpaMeVOjp7Ek8hTtzS
qg/wSyBHKNLPFnC4s4P8sORzyW13WnSJzDoD7exZWZb2A7ZYMxjf7qntXrFlSKEqHvVy3owObVp2
r9QS/Ix/pEu4hJKL7hqsYtco4DDa+OY4FrKV+HKMzq4d7KHuZt83C8idKIs1Kpkq28Mxlpwk7XiU
OD65Bl2hwedABJCi33/k/WE7+U4HC/BUzjrfdRWg2RBpLeCkKamHThmrVM9ucVVEKe/nKT4lheWU
4GEJomuCw6E8zjYuyDZXXOss+ZBnDddZnD2Um68wjpgb/awIuJzJlOscrSLwqL7rFAtxM+D0Z074
F1RBpZWGjxxgtEEEeg6gQiGB8638HABVtdqoW6HNQe+EueABOImXkIiY5oioEM1OWrGccrFtAa19
BDiXeeWqT8tFw1Aoq5uwjVeQ13rzfDfWEJbIF0NMnizPiARUeUEsH7Hw+kWGN47TVhVxyosTYKOe
qkpbjmc4B5EftyjGFFAgfr2nWGxeJZK1hIIqHNM5s5NVlLRlFcSOnIY0BQT8oZ+D8Kt6+2yjx8w3
1uRJg8uCfk5eNGqkAV8y4R7bUTPq2m43QFSv11oo44xB5fiH1+xqO7eSZLFyl35HrO9zo/zw6+Uc
nH0UHyzgndhKQn5DClP/2rxKOgz4dEUT18XCpPfZZvxTFncswBv+1BidmIC/IXYyaUvu4lJ2JIPg
cNLQdnWTnc2og9t3XHGvT9S50iM1YSKlz1WpxbitFXN7wm3GgHZesizdcMJwDiar8PaVILr2LPHm
tUSW5Je5OnQlHrwPP1Fmb38LtrAsX5budb+jo4Apm2/BBK6PNbSS1xrv5LjDP13KgJUg/23iXHaY
59b73oD+HmLIgR+w/0WdEP3dcA1+oCGEuxbHefdgaShxBO+9sNGkS/ccggXK2Eww5gzHpPTT0iNV
mfq5+mUiBbh/6IFrHiZTiPmntLQsZt9DhPyE95rkgZm1Ab7XEWxjwL8gze2upUcSZCFrcLnBX8Jv
+5ORlu0vGTE/TX0EK9IVJ2akRoop1GWtafESwEhAYiMMxz6658BEwwHTIDr439i03tp/L2yci3pX
CTc9UF/B1IXJ9sC6AM4jAUQOMEc7ofIMBXnQzlxMNzMok6Vq1j/9MDJ8l9fEjCW9onciBeFMwcpf
JJK8c1BYLwqkF4Lpq4FPJKb0ehudG6IiLGMg9l69Nwlw9Uz41XQ0bpqG0y2DxeU+oia42S9m+9JI
4VDjwITDp2Cm1C91sdw7sUBEmlgI62cIXIIhUriAcHhGLs0IAtLzTedrhna9MDNoeAc5x6Q0+IYx
UeWjwcgAZ9iNmLhp1G9+mqUmGGNNSghvDRfg4L2kOt4Ql8/74A+GcBoKLF2XKbp9D7V2Fr7506tP
+hDlnyOZTjlyBem4tF9z69IvG9YJUKFQWFiG2CFc4P/luRb5phEw3+zYHcnDhqaXjxEQh41xqKhy
HsFdd/a2zpF7GefCy9aVrnP2cH+xWJDdhneo56oRKgmmdzk+fOn13N4hDwEcUDHvQNEMJ+a7DC7H
cporaVL3JKRNp6bIeU0oCbXNHb1xNPh8O8I26JgV8kdPvOYANmDQ2osRSA9zVZXO3oflt4SPwNuz
/zNx4zh1dw+U51S2uv5c8Ko6ahVNnsSyqLjKM+8K+GIAKFhRQFl3slurp+FIi2/0dxKlEwTXz1Sw
ZqgaAPwMlBfwHCmKl3r99LxOfpRk635eS2Xhg7s/uDfaE1Pn0Y7TlF1WG2RHZi9HQ24gzGYhpMdD
sL0BsbyuJGFIRkFDkOOoiDbRiCwCeCPgtyLWmuEzCjhxrSjQEbO6Tw1nUigKemBmwL6Loz7L2laE
sAYsBi4tDiZi+gwa3G8wv0VAD789fI9s2LJBppu7Wy3M7VEDJ9qwCmj4VF3z6uSPVMd18jr9oRJg
3cDPvSQhOvcF5HBWJkCe9NpWjpzfjyHKT72ElAFFx7l0x42YvzR4TmTcSH9cwmiBd7qxfXbsZr+C
Nw/VksDPWjKgAT0GjKTUTPFBMAdeTn6kc5di/dqnTEZ2ezrou0060Gq/drFIJBk7P7E/S8XeEKjM
6yYmWIp3cwhWVIRf8bAK1CNWi6FYe7+MhE/ysHp7NaGbsAuhIH+E7xuSClnxxVycXYapimTrlFm6
tvMXB642QVlk2s9695pMu60KuS5CO67OI0uLscUAGokVPR1n5UGBTFs8VwPhPS00NEMBTCz8tP/p
pntaLSuHN8p5AFqBe3yeMmj+EO0c6Z0+J6MXhLUsXoBaYk9geDiV3aMlyf8C+9wKVlY8fsNn0HGs
OoJ6FXCmhKfU0tlviOR+hEj8Qc+IJrHm6A3/xEpF4bQYK/pnRcBOeogtiddFVzM4aHwOyuNgzj0T
wioWlJ6LFn7LxtYgRdXvnO03SHxXHssxc/45rkDYYZTFo/cDNeRZ7sHoJp5w67XY8GjG5gaRmRDg
iis3sIT/4MZgZP031Pil4IGUpcASBIXflPrybSoll3AwCtXJxMM2BWy1F0TtnbD99s9XB3ycwdBu
bNWx8TWRjVLd/D3GJwwbiaXsHpvo7TI6VXiY5kiB/k5qiclKe7P64nuetRlpPBAa919qGpjS5SOV
A2vsgoOpE30HjYcx/lwwuVUA+h3/SjrOSRm06VULhE6Yd2s8qIg/Iirnoj7daV0gP2wFgrjw+bBj
7CGv1vJSOronA/LU++kdHgJ7Ul+BJ4DOFZngBgwxfQVSJ/SH6VUDVtFYBiGQJY/X0cfHhSEceaXb
NrBPh1JT9gqgnMqqz1oy8NmGYJy5anaLsgHO3JJ9PDLOC3w3Q1zIdnohCi9VI+KrtDK4mBdYwgql
YpuZzdwvWK418s6ayUkf3vHKEssHQbuv5Zma2Awiyqnj+UXNQKzD21CBg5lMV93387yi+h/jjKU9
2O5JJXSiU1LoVjhuY+KHPfPr6jakrKT008hsMegVrz7ttwSGiAqxHQgnRqG6K+dfAnSnSyLr9bl6
gV/M5cteZ+JvQYBP0c5+Z3gNXBfw+adM53niprTwPD1Vk7pmzLHHjOuGdDz1DQEkCrv/WNOMy7us
xigIdZY9KRRnmr6vJyaNK6890dWA1gpUvUdd7rKUadBRkwV/9JgH3I8nrCHwE48n67XU5QKa1Yuq
YAZPFvXrmmgfaVKBwZFBYzfHpZej28xOF+G3PnnoQtjEebrxDYDKmbLnziCMj2A1u6M7IKNvcplZ
YHsTb6pCYJz3TveOjfpKhwpCL2kMQ7u9n9lxbczQEk6CRpGlePuvSVe1Wtq0HVokBzsAhcu5HICA
4dbMFkvV/s8DK/nPNgFTXCLNt8W6CNsy5bvihQQHpQ3BWTTIXi3BaL6s9tNYthC9pg4XJmuAgyFP
uGuFNGEnJunonIt50/Wlzx16r9Oed8BW2ptft2xL3f/3eC6D/C5E89/f/6SXhRqCcasnBvjInZP8
L7kM/O4H3Xjtd88uTxNjfBLhdlW26zrLT2L4DVx/nqf8+rjHA2redPgp7hznE86tYNi4mNtactOa
SqrVzVVbZoOLXAjjL10WTnRTtlODZBpDkigiqlzw0q+wnfPn7Rq01MPjDYb1gfUfWdbD5PYLgqiz
rJ9qFX2x68VKs/mgOOduPhVXd7GCFoxIlvwpgiQH/aOs6YOxbjQMtEcsisvf4mioMEgtDD3oAo7M
dYLY7yQXicgbuKJotIgFep3ZqBRvPvoiw/EO7iQTumMPErbSxCOufu4CrH8CL/K2VkQ1c9+3uSup
tbUW2VSXFz8beCoaP794cpNu1kC/RSg3ELqiiQdYjZt72Lnu3E+tnMCFG6I3DKK3d2Nacvgw3Vv8
jB2FuqUmk4Xovfqd40WyHU/VGS/CR+VRDFTIy7rDbICuvgqh8DpyS2OxlsJ6spEEkxV7g9sklFUN
pc9UMaE7bWXZM+BTVzo2E2MkeSklH30gXXz6O5Z3VCiTZRaIzg76l3m7xveS4imnwv4YBeDx2OUh
Z8HjYDDmFXpe2SU3p/HlxRCHN+LhTF6PiHIN3ZAgUjrtx9H9uabHgFjtozVRpLzeQv4COIVCnxDW
VY+VLAl1YcHouAsl7Fd60/H7sHV4yZw67FXJKN5VvWUuODIW+7721a40YjzeuO/7+QjbE58eol9r
UheKKu7bqbQKM0wr6xL5lEkXhJZhkezEFFo1NrMofwNivSWUsbay5+EYk9CxZOxfQv3rW9d9Ajxq
/BZ+Z2kW9IDsIN4l0byInZhqrp+6udABwq4hJNbyukXod+N12j7Gntrj074rT5paoKq6XL7WZsvT
HlSRiOfPPueXlR2zNdPRfL9Pk1aih6LHPaCDxxfalGJsSOMOOBprckcpC0jbisRtKJNM2OdwhsQ8
06a5cY78a7kj3VNJhm5QXG0b+PfVYU2RfrVy3X85NUZq5wKCpAGEg80Q2ORCBja2peXbFv9urKJQ
zaZeAvkDlKEmgMfb3Wc2+emXWna09wBTLXbfUXBBS9fBRGkNaLc+t8x9WLJ+iekX9pqmdFx22oyt
vcttrr0r3jd1qwPd934Fvtw4gCCk0XAKl0gC3ATaQYq/t/mMTEURII6am7JCBXZXw0OEBkHb1PgT
3sdQZg4nkf2is/ZbsKQeNLEDnIo8TSzODzwGUTDrTvuyEYhGbBMEPXF+EeC6fAIOu0rdZLjylWY8
iyPd8bc9Pm/BKSkHAMl2K8xqe7TS61sozGdZXRRLoqXASoc9xMsmgZiZ9rvLeUsUO+AStdml9tJ/
Ykth+gPEZ2xd5jY1qRTVAyEesFhip3qDMcDY0cvHhFbZkcJUAcBt35HL/FYH2cecQUhZhmioBYRd
ANLnesPuJvaNCpJqQibSDminGt7kJfiEhAHimhwKKrkAtyELlpU84Sgc72CYhcRbEl2jenwB/uyw
q64tyuPpkeEa56b+psvlsvhKpeoHgOn7kAHnF3xlcLxTOwQVbrWgCXYe6WLpe42CoNjfls6UOKFw
FYWAz41EGqaV2r9kvqWSNy+6IuRp5gRrvHvo2Z0S16/IEnNwWoXGJSKmljD6eI/OkGLhNYTDCCno
N2r0SeM/pToVLUiLJ/fDKuqvFXbgkEpdJP6/Jj5VdzPfNv0oIVPe49h1P9fWGD+VsPPOGwOPJUmE
mjQCB+VR/qjJXFgc/D5w65l9LvKKHasAQBeRv/x/NJcfKqgf58tzzzC3C8Z59HpmD36NX0eSogUz
fdQLF5tEOPYewjz5PhF7rLTX7soh3h9MBj6OkZ9lg8nxqMNArCT8pPFr1IPj+doQXLmNogYgILDL
IslKDh8q2r++EYaa8USVFHItaCCzy2boMqj811cEfUcJfLAdafNajn2dv8iucj9B6flyRR4a46tx
2OPSzP1x3aHntTZeZTEeQoUCLKp1wpRpzSUfFZpFgkWxEdPqn2eUog4BSV/tHU9IF9gUnmmDckYM
0/lFatxudTMaL2gxUR+WJtu3XxgwiJ4i3pI8cdlZiifg3qdxWkJO7srlJw4vteXRek7CM2bBD9Lh
M3IOylXDNvcVTcbeVwT8l7zu8QWh3SiExKstiNP3bAk5JWdsBmepMOqktX0XqfVLklUklOp67eVV
NKQp1p9ILSSiionL9nUBlq3pOfvhnhyEYt51cEWMIz8D8a2a0YNxhOnzkRajUtQ/Jsf36o75vYbX
DGq0Wa+yGl4MkBzfRyqbOuXj6vzHKkzoMQ3yUfzgwNgTWk/7rnzmQpVmOUYTknO6RwFRKrj3Kjuu
6r6iHlp8EtE9YeYrYLNsdROn/+pjG9c/m5E6bJwYbvyVwOSzhjnr8CVl1IdjrrEpeGePCyOjzkxp
1PeJcGtlMYRDbN0kyBKiWQ3qDAt/xqC1K6V/YNo3JQTRSkqmaAcrwpKZocW2rTwK4MGDcH2ankjM
9GXbQHU8c/k67ms7fyLq6tN+Hu/q/aitHdQF1jBYAxuJaitkfb4v2RI8sk5r8i2baTlpKrU2MphY
WV/owKqmMVIQh92IkEPbg9PuJtP+klB9SEnGLUAKURdiVoFtQBsyb6l+8TNrKh5qejXScuJEZtyR
vasKOMAnxUCHdXtqfuxbvPHZNEsQMXfjqJHzu+7s6tYJIuGcisE/NyOo/o90fG6pxyv56WloZpCN
e36gi9kq2tEAMWC+fXNgzo5f7/JCeCoV3EzI6CbEeLEUtrDYc7CgqiiN0DlsyYBjNHgY51lCE75b
1dvcdnaqOOxbOVyMpvOtxgLW6UqWYsFiJhGsUaullMG+O2glIvxx91C4NWR6zKAGBUMgdpeJphE9
RF3dVelX+4S8LnxRLaXh2THyrgAhyZbimIKXU12LcnkOlGak38tzumT+TX6wV62wsIMZERhkC578
jO7Tqutzji+oq32VSYSjI2A0FwZGqhOMyU8zQT2kjzsDtbGLTNVLTQeCd7zfEGphxZajFKhMZ1jI
0uoC/ALQqnxN+AivBm4fyeOJS3FwxsSnyHI201Q2svBx/GVsuJOzAXKWqhuWCga8vS7qnPWYHPUe
HG1K0XwmO50V4DbPVgS5REcTUliDIZKLIxgK3MoWP1HvXGrqjAgvF6ZcT+dtE3LXKEnMh1E7TeJx
bstMw7OvDGGC2uOhCtrVVjiQSEgUj+WqDeDeLKgasix/0Os6YEF9Rk/rzGMqWa+yPMHoYwdLneY2
sMVt04azTt7ySnWFYPGJ2tq/w/EmNH/R5kSAP2/YhFn7ZwFf+fsqqnDXqzkW3wK5QgsQYFwd71r+
NFXlSh4QKtmzbSnUWJTdLzwrjsphjoL5gG13oyDMw03OWIK8NWADbEybYvvcSZz7FJKZ7kPd9We4
qqNdUaVEiXtjuEGG8HwnRp1SOT4kKbsAGigYKLbW++FqRJC0Mz7Vjj/MO0MqzC6gbP9HIPwSyzSX
B7JgvD3fdrWsJBtS6qI9SuwJhttIOXFVYp0+qXhIfvzFrI/e4w7yuuvg58RJ8WQLlthsnboP2bJo
gNbGq/6RaCP+gl/Foqz7NiUsVUDxL7esHLBZlEYL0k4NlZiU6BMalwOztVY/DMTl89ym1B7TSubq
tWwh8AgDaFGlFUtMBB9bMAwo5+vk3KTLP6iXS1MFzPx7pzxp5XdddpVlxol6YM4ormmdV5AZBzOB
qly2CLp0qHQDKjU9mjGmHidoVPjT6gresPXi/99IvZFr1PHLwAFcjYNchL5pP0yZYCU2NwadBsah
zT920XlTRNz4Q6+V7AHdVEVYnP2ww1nXRO6RZuI8H4HeTOifz3GRCj43gBoNbMNVALSDalOlDUGW
j+gKjgwEbSapYIRiZGtsZgv9tdhfr9JKdlxV4BO7zR3L5bp3Xb44aaoeXhXCDkN2PWt0QOuhGpbc
g9SSVgWVk5gcdV316KneCKuzg7AkKTOuFsBRSLo7w2c9PQ+bER4Eol3CTBa2lyWgSnEifMK31HDC
uYEK+GZx4yBmn5fQuoNqivdck/8o6FvFjGGMg9w/VDYcWjv2Vgm28892f58mE9xyb52lvtJfUShn
P+rw1Xx02V56zsUWMJNA7WGIlivoa2j0vnk2IAZFEcUfzKqQ1sFZBwVp+GtF/q7y8kFyMXDzDzFC
RddDs7XRANK7afnO2kC6SbC9qzN6kpCl1kPzUjRtO2YNBDnWZPJX8/Qcv78bbSKGR3qh8DGXv8Fn
Lm420inlE4fl0uOuWkOZ/GAF2CBVDq0qBu3e1dGbpJAQcOuCeZEiD92yws3kR7k5ewjV4WhjFJ3F
4TFjvgFOa9rF2gTnEPDAy2UqIYJYxi4xoS0uLr4RRrlQsRKsXge5RpmmMWBRI39rjNhNtNxvhL7W
MdSjchrFGvo8GpoSEpU0s69cMWn2nOaAtBCujwCclqSfn1X6rDt1zIpU3WkzK2tmhJTJbaO4MUAo
uM7B83MxlMvmhGoDk2bCks+LAhCBXbwUqQK3r2NCAmcM1TLfRaAIP1aGxBeuBYRE9JZzv9sDgO+z
3X6KmceMQVOk9yrc/J67X1mlsVWwwOsSeFg5XzASk1V5Ut4UGPSJxa7lxqBHpEExkcooZZKKsjIM
NzxVtN7Uq3ItU7XrCIdzrNY4yIFFljDW9Ro1ZtBqsSd1VbjszQVf48CFvCm+GuFc6kIxAIW0Vktd
wgtcLncxFs6+vaesBib0NxZoulpSAQqPpYSVbNds4ZvIdIQHEkyXEWn8uyISS1hgXHQcd1RDig4W
kI+yt2OencLCgcFIzccPm/muQ1sLDQZmZpD/c/1S9o8HTYRymo05TE4wLIxGSQu0OyllaMnqihXp
l5j1ixfrAdyninwANVlH/l8aSWMM9PCAnA7Vl3Y7ikKHN0OTIujdnWrATETIKIUKoUCa8SjvDt2x
1YAl2Uy3w8Bn65caRFA6LYBOTCLIG41yx1GBOZVgVcqxZa2dk/5QQvjkOpLmX1XtOAwTX115DbCB
UILY4uN88zbJAohlIVQYRzIYhiU3V9prsEbF4lz1vcatW/gX1s1zHH9gMtTxkUSgdiWooxXeycru
xZVUcAt6RviX6mYnO35MOXeWjMu9yS/t6+P4+XCNy3mEkPX2/VOTzzKmigKuvSpFS4JKDbPTLZ5S
mS1r63cNNDeUZVJY3tflTspyBhH/G0AW2ALWaAEtwrepAVxDDaiChhu9LxNml3tXvST+vhjXNIht
6ZZ6tbfxp+gOjR/kbHFARy0AsaTa1cmPoeLCbCSiMWM0+09YcGzt0mxDdXbik+BWEX7lVYpl1hor
S3Xw6sU2811sR/cuZvRnzqBB+ypZkrq68+5qpCtG2P+XkHJWnqnjb6UTofxdS5NUSTj2YnlZCeBA
BFPG6MyLQVXcldbdz9jHeRATYfkGJ6ZZiBLLSDA/4sHGUJlZfb9jyhLAa4Q6q5ElETqnwQkkQGh4
DhQ4QP6W6UkjguVWM9zaLt1xM8oHQCOyTPpQ9haX9DDTP8R7RE+neRBMxoH2vyZHPnN3/z4EEYgz
hGtmWcxmliWZCzImS2ImpTN9SBUy7EAU9ERztovfKBSWlv7YcQLLTBzxrdjDegesr8YjiyiRRO3z
FaKAhYwf8D9O8C3JvpcwnCxcP7i3HyYkF6pG5k72h1FMF2UrRMDMxhGQQ217E6Z7WP8NSDdEMiIQ
aaeKqHnlyjE0xQXjqXtXcZyxj/XRFZATUyZCnWDqz5iibpT2V1Qozy1VUPVUU9CRIZcRoQUMgxWH
lnAR0PjLsUbEZGSa6TTdpBBT/Qt56cd1NnJItgtQnDOQo3QQQsZ0hlle/RnbY34jjsrY2ggXhw4g
spfZKN1D53wFggr9oUIh9qiB/GbOczhp7+Qv1fbPjUyEmcesbZLKGggnEQNL+luJe933L5HibVh3
BEwUWpG66o3OINO8hJpyi54+neyRMvMgYpw7/i/GjhgJB05L/OzxVY+mViNVdMkxiaqQ0Y4I2VxX
ALBngP3kAOMjPxm/s5nvtxZO/4Rky2ltkrOAUOAA2yKmx3txwywQ9kaxTmoR7Rr2Hl3aIvOuLoYA
t96Nhh6kogRdn5Pj6p1ys8xF6Kw7P+eISTXGUZGenX0wzar2LEAk/+Hklj5+XRZABueuE+ndznQ6
nzCbC03uIKZiHykwgZ4vMyysM0RoiALlcR/7eaAD9lcB0kYhgjqw6Ydr+C/j5RLMnP065e/cr1Sa
4ufgdZJzXPTkKjqW/6Nfj7ZdmKMEeYsuxiBqH6uMKT9I32UCZxeuVpV3mMmMNhWVR3rzWUw5NxIH
jM68JTyoDXvfXg94HgdNG0XLrH3b/em1Ky1VvvT590p1fpoIMV/lP3mmU2PwXmHFunMy2aggr1Dk
nmqiajXr53A7JChJYLnXtKxYQ6XooK3vgpOYyCtn/ovSCE4AoFnHW8yQ51qt4i1E5d2nNhYZ7lpa
iuMLTQ3ozIrHHYPlHOcDrodvF+JSWyXQUsk2vbCfyS994wFUQbcMrvUNujlGe0sf9M0w2beCWn0F
mjUFQ/pksr2SDBQgr1ioCFnKar06w72BM5KSHZFzSXqvfBup77Sl0Z5NV456hR4pUgeKuaXNN/qY
sOs08WYeO0AVMjK+2W5MfXCOG88zakQd9bis4rd7nkRJgrThqQY8E7DMcriDndBvI/kR+lZEwUSD
KZ7OUr8eI/EKueou1Q20AqAk/aDo7tDPcbr0E/gH+q6csIAhvyETxYh6a5cmw7Lb5dXCUNb5oKMP
4cKFS8lXwwGEiELxxR3cdlMc56ko8cC7AQ5odc2tFtD9cWVe+adBc+gupDZafNtTiKRWGAwdxu3Z
JHdfqTCQksWMr538RFQp0sE3oJ37BCD0Vjxs7Is6oEq8u1ICCeUIxaD6N8mfT9JzaxiqIOeYh6bF
fWxal9zMSIC5rExNroapQ47RoxF9cuxqewLwteYzBICcmBmR+EPmteSMXF01fRBWTGbtVmXM430K
GKidbNDFCf5aLePGCcLAgl8vTQQbLebpKi3dwCclo1lUrGvbhUoMNxZZI72+Z8NNb0lDB8N7TN7d
ZM4Yk6gr3vchO775FQfLdxR/Ic9SO24R6tamHXn8Tyt7DESNnaU4GlKlg7+6xFPEJG8UjWFYZjmk
KBTClQn4BlNgY9fvqEQzXYJhtokpigCw1GpZHJ2CyBoXFfexyXzkUIEfJXKO1W59O0oDggi5Qt2Q
Dx0WZWY3cYJELNnvA08/f7dY+PTFoc9tGAu//A+I4N1uppUs+HMmWQrDs4VYh+Zqe73KzJX5M8gg
O1hvHIUyl2Oq4tra3NJ06VDdHzX+OWR3w/yT5/CU9wVWXKrpTwpmpylVwkr9EKnjaZnAjQ94jQdp
iidrCbpkXJT5ynfZTQGEQ7WhKtC/o9u0D0FCCnhT2CjDD88Qvq+I09yNcZlWotoCzyKmRJeiqc24
LoIra+PhNY7ineDI3t4rtj6bbIGtAgqXLG7LDVT7PIcqp+mMldCHaYBYb6GtkujNCK2eH0SPL9dM
a9T0cFA6gesUZTd1WjpeFTrS6VEuISMl/QQYKzIMX/tJ6jTIWwHXKB3D9dwLloOE/E42yPFnNcLq
7Fb4QCqkZbMxX2lTkObTPGh7p+G8TlARKdg43nI5rXlxRwGXzIgrPMzVYL0J4zlMlh58wBblsmCN
9NBqZg+sUP2AMneNVsRytoGU7ii0lRohYyYeBnG7Ps8d+0+wj734He497v2w4WZi2m8KHCDTNXja
tBB1qONCx0ZKsfjEa573AONC9cOBONwOLDHuiBDI9vWJEKHSyRVNWwh6Qvz/u8Ie0bMsgXoGjJcT
dcuZ7UY6nWd7KfecIx9lZmmcex++ytji86+tRktYgN1XDQIYuxK4Wz32aMaBV5TMDe2TCTNJOlcv
1/OPeMVCTkYv66WslDvV+aOf8JBGZAboH1Z3mwRhn30c17hWoXY2obr2IooPXm3hgSv15rLJx+10
vM960TkJLrYBQTofDqO8U5+IwcKEQ6J7AFSOznS/9VKXI8aSX9UnKdq7ryhV/0zjBNCJUA0QOUvz
eFZV6aWe+UFHymArIbYqxqLI2UIalP0tFq3gLcPl9cuLqlsRcXDOzyfHDpcMZ+UxmrJe7D8fXA04
rQdYsCZ02DAq8wzJrkYzsD4IYPayCxrNnXkV4abMYYxLx95XzvX+rVuIJZYW5TjMtqEX7AH5oqPf
xe69we3x9iRNei5BrtA/u+EPo6GmwEvibkN+oHdjqjctSwhEhsO4K6BS54WhKRHuj7kIb2GQHG82
nW8mxxiCghfchU0/mb+iO6MMJX0jN6iuiIBRoCMCns/q/wFfKbSa4iB/u/hcJmt+NSAK/GVtQiF8
2iqJj19IkftpD7Ib1pDieNz2x3dAXEHCEBUbqNRi+9jMi6v5AKPC+V3v26lXdZeSqNFnrH5MwqB5
ka6JWhhoHOIG6gS6WeLorgFB/f6FLpb9VZyIZJL7ZPU6V1F4Zd9TIh59Q9vsjbSm0JOPEuCwQydV
z7pBZZLQ63LY4Z4ZIpLO2y7sSDsPGGGh44rZ8gl5XI2djcy1A1Xhh1soPHKnNYARJ9d02KfpKTaG
Dv9AASjDLz2oc2xMnJC5rRSrW5khdsCTJ+Kq7O66IhlTcu6pbP5MRBC7hBv8h+n1J0eeJ0LNKt8/
c7jHKkl5Qjv65f+0ScFmX37RRnrJUFzx3t8in2dttFi4aFchUfW4+5GcSh3JREkBTnp/gtFGF8vI
aMTWEpvws4UnfXMZOpaAr8ynmDs0CuDuMhmR55DJrfsXj5EBVgC3GeHXUgoZeQ/3oJjiuL64kEAZ
ksouVrGSR4METf+uZW/J8rzC3UXSbl+ksclXo2nV6wsFH7BLBkLMbhSE56J3hI8XM7ka1ZxHnGxZ
ua3xvYxRa8OUHlskymktTD9bEjsr7U0E80pRa59tZMHK3W4FQlF6GEd6YzFbmLKF2+6f9TqIxU98
YnUvYVC/+8rgCFfIk6iKmpWgWv2twqBu/WTedrWIpN+u9YJybsQeDNW05f7Z8gV2VA6vMIt1hvyU
L4v8p1KuEY5aqb7zjd9UsN7pyMF5bYW8fJMWGUZ0nDLdowVcy4Wi3e+J+4PQdCgXI64mfX3486rr
rFdmyetQ1ML+wD8c9IULJT7VF44GuTuMptZIEYRO979g//XW3Fk2pyTIhk8+aLD7nksp1zFEZubP
3k8LgR38bSighcZgC7cNtGGihSO4f864Tmw49r/YCSDlGUWptbiazDnzepSmYp/cYaMo1r5g/LsA
1m3VZ+7otyg1YKxN46eDOuXMwL4wrwU1C+7GlQ8zKLVQrf0SitLkUbuTj3NkRGYp+Jx19RmZImyA
9/0JQvZrfPSrK74+xSUoaYat9oLbR6Y/JYcEMrdHEZGpj4IuQat6hNKVBQzOp2mH9je0IIpVt9X/
yxKqcXXivatepg2PXoH9A7YLhrFf+FVwNLTm+rka1qFSNw5CCKtw+czfd/VTDfQYC1LuOMtFZS7G
/FnF1DaNHHyYYyRBUyshuM6FdWcHZlP8sLQlK4E4tqXa6unNK82xx9lFJ9JMgNg3bhlihf00vJm9
yGzW52esYIohhi33Mq72vFXOkGMid9rEWnnBX5fziU2RlaEDV539x4UkSF7xDDaj45cUQqdhTCVU
rDqbm//V6Kf3UT7Rcv9l6XIUDO5xGL/6biywdZV7JQ314KjXAh+JOiJnEC0pNIQfzbK4If+2CVQu
/WqbWY+cE3q3GRNTBx+DkxdieV9u7L9TPTZRpm6xlQjVlwvh9MbEe2awYNIkXKKByuAYJm4kZ6nY
c0oEuN5dF4wHLlGDVkf0IwbizqLQLfNISIq9cVxicN+px8we81e8YiD+hf9VNKwcT+jt6ALQrI2p
1mVi8CAuUnXlcUm523tkTwvMwhOWjVR6ruk8PWYABufspokif6CPwhgKYhPh2qKptyQG1jOeOGyu
BQUmj33FB6PM4XAJHYY9nD7meKImT9unM2gru5mrro6x8EyTvGQjl3a3KHOBRkOv0RGOqVrR3YBJ
v0y4oVwaDPpDTaFYe9YnavYn+d7rnvrFfvprNSRve0Kqys7dC+tE6RPlwmjT0cnx8FYsFNcnvMBK
MB0GpiRdholRVW6qa6gotsmHTDbBTeJtSaVpu2PYKs8WWG8Ml72FpXHYBRmSE7ehZYb3gSElPj1r
1mUihSU0icCY/xJ3QrsJ1sw1MTIluv1pD0ubawtjEa5Q+PiktPsYyOVXiPVR1P2JPs923pzzSdfW
qUrm8KlqsaetDy9CmzUtqrtgygEjGODK2n6dDDHfs+NVZuTY9I6hAqcOpUqnygZc6rTaHHGgPFdx
nSSOTl/zSBjmBunjEC+Hxl9StRPPZGF0z6e7f3z0SfLZY3IqzMx4CBOch79KkIzMDHaUCo5c5EbB
Q2YfTCPEudcUJGyjG/KgvvG2DoXwuJnPVsR9bXfDpizj2n3sBxfiWFcdgZKlRw/LqUKQIrXD/lfb
OEH2IwLCK67j1gJn/QHSdYjsyom8YjtzP+/MDFzVdt5/LXFdVaKlxw8PW4VPAU7gMpUy5qx0f4P/
+CKF/aArLdFl26hZ2rZi/Z0Scf44SZL5bLWor08+qKuTwAgdFoL977MLyHpzo7yeUNcsGR4gwm96
6mdv+44v3/ypSpGhjXOlCT4J2TWf4eK/baGVN5P8u7euAlBhBBwHB3UCMPN9kqkmLmYCSUOl1Bti
uQJFyw58WXNGXCwBP++ZEELC8ErA2CjW4U+lzhi78iMRFmjMF2zdb0ldil01WwvVAsYaTb5quS03
T8tEEJlCsK5RHx6vIg1JfWhLncfqnM4qgG/GbchuRSQGE+cTki6Ij09ctldlxAxUDPZ7aWfbyall
zVg62iVsd563/XJyd5HGQuuRqrMRDBBm/R44plMB/Wge1IO2rCul8LrLY7yjBzJPNz8lL+2xMRUs
E6vZHDGzSq4qR9U5dZqZm1uzs7nqcKXnzbiszUZAYzHqvSScIuYOIh23gA5isq57dlpBFP05w6Uy
dFjE69Ud4CkPFiwjagLfOv/ypoZapk0Ctlbvcn/aGJV7+UOT5wOVeMS3615+Y811vTB+OF/wcxTq
Wx7Hg6lOcMtqd/GYb2g8koJUXJHv3RArbxS0iPDXdz/L+Jv8YUM9gdyX2YRGzfOdCdMjdcW6eVcz
nCURCgSSk5y/kDMesFW+9yF+SGnP1HuoQ0MVnAxnFoxZcSsZEoi8oP3Cc7MF6AGhjOFhkSZMEtaU
DkvDFSlWYo7OCYP53qa3ys6yPxUO/KHhXADQLPP83tmbH/gCE9t0H+9vcULcQz28caPYi6OTMQ3l
mKe2jOQz9wvt1QKXUVdDND/4Is2oxge0C0UJNqHWCqT7f9M70FPa+fZbEvGjTCtvIn0PTVaGBYzW
Mt8ibuC3QxePX7eMdB/R+V+tEp+dodH5cEmXw2E74cUsoKSUWLcNwFDIfXw4TjqiKjL8b+HtxxD4
RM5MdW8Q9XtXEJYQERAHtC7+seS+AkpwaUwHnkq44BUISQOx/7b9vcAOrQ2EvZylQmjOFO0mLbEz
STJwdSc6Xnp7bi3U/nUPCV/Omc3eaZjPxY3NVa2PelcBsy6WnpZrRo+Q2jDe8GU7+gEcJz1ktyvz
R66w0mw/9u4qrcn0td8PuYI0Xfx9zUYEz8N1/x19mTmGdSkJnY3ymF773U5R7fr3vqDImd30vfgS
eKUVFTbIR1QqVqmSRh1DUDXhsQ1Ezduh+RncBOTa+pVBQL9SPZDpDmJPV3pLpDsY0VcYWSj1Udh+
gtpMwsIXgJzb965H4F1x44Th2HABlzaC4bsjMkYBS/iCAALqqsJunHt25J2fV3p93WZeCdWhMGZf
43omAnKa3NPTP4j0KtvSp9d23wQy/aVkhwf6yCmGPk9Bn3gfc0qEkYcx7h3Q4iBgefeu3mTwyBPp
JJGMeyybT01QCBJhfG+iAJH5M0IvQEK9T7+PBKYvj2sZsXINQCqeDVktrt/UUij482T1xsyWZPl2
aWj7Y8BWHspcpaQt2O895Qkf/ee+12NNgDLYCkNs60EBLMKUp+VgxWXqhZdPEJjKGKBgdjs3O1yk
iWIbsQ8oyCNqVMSOv061/d4CcPAUEHwxu2OJ2E09zaAINsb2o5+M0ImXXyRcng/HlQC03xFMfp7k
+x+vJPFyHaGBfY9CGDIsvIVf13PAkqPEIUVNeQM+QVmvLllUU+BnBdoBav80s0sRM+/tgqhDfmSz
EzQolN34DESOoU1oaQMwGkj9tDvI2QomVnPHUBzP6NCO4qlijEukEEvkXxR1S4C2OM6iSOhdF95e
M/0/18lrOaIttuKLc5P2hAY04pb1gabXAoP9nTjyiy+4zfclF9nFk6v6CS7RsBgccisrpKV6Am8p
rgXNO3zozckBFFZ+PEN6zfhzb5Cey7lCCImcZbeHGt+KVAgGXD1gYmjpckP2BzcWjVAMfgbBBK1o
igC7VU3mtqGGJoDknLSZiK2RX+wMmTI3eZed/bk3rEn6OeJcBOyk9gM9WUlgECOei+2d/3QD2bHO
ULhHNKXlhhojnID2vQwLXPrEQ1iNhwsGw21avLEekYlxxnCrtCe2+BiJI+PnFnGxndSeSIj5yBAS
urvEXm1DW0kMWc7SenuefF4fdGC7PC0z31xwK1mzQrVCAjs03hlslOaLnZrVxJUfI4z7rtNm4Bva
m/1Lp5FN+JDHaBULdUtPrdZO1BRP3jsHY8fjDmbcm0plYxDKv7+tdG27qk0r1OloKgQhBtXu7V/o
slbZyGMzd3tpLwoeANQin6g3FDG9nDpm6GwOHb/4QjfV/YZk/ugALN1BH94QsCZrN+9PD4U0nBbE
fng+6E7SGd/WSd5IyouGqhiMUcxCmxJ/vTJ+a7zRmIMo7dWva4WUlsjdCjCW8oK5OG6ccyCPoBco
T5veg3x3l54WYS+MYio+0VB+rZFnApYA1WeRN5Sm8u1PzUHwJFxllWhyDGBoLfaVh9ixQBKQdK2o
Kh1sxmRYsjkdQkfa7ySzufKy5Ue4RwQknJLgQA7dwMS9gEDEWliYVb7us64YC0RMpXydxkOgys+P
9dHu/JAENYrT4vohnCqqpCgZF+ezd9C6PugmmnsAhvBPFvhWokT7yAsg9vvbuqW2vSSD2xJXNIfs
I0tbTwvnDqSDn+G6l9JqheVh336TX3uaDWV54nI0DYHJQm6ZPITCSbQcpmzzVcQSPL92mhrQ1LqW
wOzCbfYM8Jt1dzy6a46k/n+DYTEWQm6QKrwoXBobszlj2ls1FlzwoqlyRguYuPZGFxVldRzuJIqe
0NDvpP9bkptM07fncf+IMr+wYHr7u8jjr4djoCJw9GdGfWJI2s9GuulnH5VpcoD9urPQwo6IhtCa
RlIx+dXkn3E3lkGpTRKfb8PI7TvCmMrnFj98qzfrps1FowINQ8upuF8M9G+chHAlYJwMksk07ZQ4
sWASI5LdvxE3uLEr+OgsYeRVlFYVDPFoR2U8anYgDfgcot0ODFycneuzAzf1WRzvk3aZm9O5dzkk
PLd2JdHvf7k1cZetLM5sXQF7TiQsALXmLGqwuWfAHf1FnPO6twd0SCNIgJDhdEErxF6sCHIY0Rq4
8jlWBASdgCNlUmva86PLiTZ9bISA19jrA2WIwpcSrq64oNcfwJcAHsLVFbEae5zDOJR0Ug3g4SPJ
AyJGpvoVhR49PwmtdIwd+8PEY14dXg7loXGFPmO4Fu3T96jl2jRP54g4eAF+XGHTNuq98vsxla+l
XE/lBchO95wZYeGpUwcjbGbqcE6MXatQ4L5v2oZU6l5ADgkuIqzxY/vtIqbEqAhWT7G9DH0/RsBO
JwL+pJ0OQ3iVX+cbbFb+2BTpOQQCpB1pc//DXnOd1LX6s5yb1CeG8UtJwJrkxhCQSt/nNU7G2PXH
KIA3JoXDptpbhw6Wa3lq5oiP+yTfp2NuAyoVPmsIwKI/ClfAjS2IedZ3pyVnw9n8gGwR/Y46/UUo
RlMXJ+JR81q5OX0qSwwS+0woansbTe2TBTTheq96vTDlYoLsKFPOsCnGX9hPmXrqTfp1B5I5LqY3
b8YgnK/tZd0iEOwiSYPCj9o0zKVJtA7c30yx9OhBIP7e6lQoZqG8UM1KUenD+QLVHc6TiLlFXpC9
qm4Vyp3mYQpiqZ4nS3e62Vjsh7NHARbfWWQIPD0OGizJ8UDetfc65CvxZHvI7/f1Ps4gk2msmQac
tOf+mVkwFI0YZX+jtRqW9Lqpu03zqS7dvlrcjJctYo3N/4Ugd89pkNbKWC+qQ8wDgWvYeeKPS4BL
PyzR+0qSVnXdGhsMVWk2UnC6ZhKsE6yQM1RJLgstPOEu4VBLyezAmRMCXppLH6aHaD1Z5cjPoHr0
BJFolbTSUrbtDr8PeQFdGm4tD4ZO/BFc7TEZJo0TPz8HQITrFYHeLeparawUznp0Y4bsbh6QG7LU
gYN0IF9Rys03N7HFdkeiVoPd79S8L5N1g0H/ltz0q9aQLiteWQL2IpOPiUjKK7oDsbf0NcQZp8nJ
44/RYA2fteUHjPYGqTFEDdE5FYcKyyCkQ16+cn3bjWKUW/fy3tHe/TQj8WfVg22FE/NQXupLICgP
V9sF0LrsO9Au1ZxEwcLLVZu/xBG3Yr2L5jX/NKQm6Rb0zd932NAnu3ekS6BHB+bUB4Uz5jpomTxm
2+BGUTZ/Xw+2YA4WPxLKWfi+wMZKWWj+FZe4zHd1LupYSTNvVkm546ivBmcVUX18iDh0AeVpP3dW
yhQcMez2Ev29j9tzYPx0iZ3b1x+7PBQIKcKUVNh43Id153FXn4BZttONie1Wv8/TJ9AHsbe0aKAY
YuO/G3VszwTXlgfSsO8peqxBmiT56qjp8grJWmFLy364EQcct9rn/mXjR0NEj/U4dPTDtBdqwRqw
//p013jByWDhhFiAv/GDeTEtauA1/25LYR0d4JrmFBgumszWPwFE3rsMJ1wqVWPvUbaVJEe9UD81
eItE4usuHZVvsoTryDnLLm7301iYD/NNGIyBwexK4cHH0sCtiS2eCkm4t4eLR0yYsCaNicYg/8eq
/H5wW5OpxxvEaeeqzpG4Zg+ww/mef6WM7DpFnw1rXySGJzrRj0SsfuNLnoZZxJeU+e0zpSAiCIpQ
KoMDUjinMptj/hvUW2cnXznF6tl6I6hJC3r4n48byPJoF/Ga2xKkAECxbJMm7ENow7NVjn3PvHAk
zv4NeVNMfsbOT/hPlacApyRH1FMY9+CTsuJOD4mP2PYZMgwDSmK1pijp+eJ71Lt9Pwae4EF5qTAE
MvV/S9cPWmUcaqdYyRfDzlGcVv7OKDTPhuBZJs68CHPDpkVHaQ6Ec7rTNQj5//GKYfeVQCK5cz2o
yWtiV1MMId0uSMQwOZxVTzEYr1VIwaSe/blN8KtRISqKgt7hjucaH7nyqQod4I9Cb31eYvn6xG/R
ryL7ffR+g+Ql3/HNhWufqkF/kZ1lA9X7q0GkSVumx1QLQkXZ+NNtKeQdtcGgLsv0I/PD+CRZLPup
cMuLmp+K+RoFURxq8b1jZHBG1DD4z0LI2I6g3Jwcp3p2N+4wMPvUiC21YlJIPVtSjCF8B3TGWigm
Vkuekcta80AEE9XWZQ4ijy6Wcrn+TEPjPv75WhsnggU4YNPSfuMursySjDBmcF/bswpx4qLiGxNK
HPCROuLkfvbZskVu11Oh1BvfnrH4LLEgOg2Cu83Gjg2vqDuDenvH0G0QWLb6A1VMWboxOnMGAQrC
eN/55TtLO9ljj7ydth+LG3QVflyRIqrSYuYxiXV3/O/ITEuMz0Um4aNB2HL8q0tNY1XrRIHAhKV/
9myk1+83AqyjL8Vd8JUESZlkKVwayJpxqQI6TWoCYCmTCI6HOkChKjQutJUryMc+W2mxGfyUkdL7
Kariiy99Vu5/u2wdgP7R+IGsFh8LvZz++wmi91toogU+AjIPL4DGoSTp8CClJhtc0FuYEoKaqqke
uLDumk5eYmGC2jshSzB90alTLnH56chlMUGkkQzY/+twlPJZKHfwYRzWLMjY47XGcr7/HmN8gBx7
iQhBxX9EM/BGvEfKLU9O6elFVdZjAD8MIpodmxj4jZP7D5h0AErx+SBhwj7SZrB27eKamWNuE+rL
8IBDhQ6TnT4/b7mF1rD7xp8C66aab5dhzaTFOL5ha9PT3D3S5NQFvXT6wo8Wblh5avtyIpr+HIrb
fiGt1ocAaLkhWJb097Ku3SksE4TzO/g69MveX9gKPvuv0c151hQzj4t+HSjleuk6CllaPlsi0751
JsMmN1IBzsJR2lN9KWAKsYmelHLK8jUru4YdzMfG5v4Y7bFPRtia3iSHh1llCRFP+Ewaw2MVecQf
suNbVr5NQ1xPd8JHRv73wEG9/rFFz/2gG/2kfV5qSH0LWpZd/qc2PrQ6CI3PoUxEGDkasNR/UD/X
m+ajm3lyLIPTp1eUuthp36zIpuUKcg7Yo7OhNSeT131SQvCXJ8BfKI6jQ39J7xdSy2M27ovHfeQe
XfssmE0hASkZ+/JR5JmffPojx7zaPBmmzzygn2CSh7lUe1SCHJMC13wCIwkzr7/JIuD5thWZpIrk
Ik7SkPDHoArd+yFFIYNV8E5UW0aKIXDL/CBUDPCBTA5k8qDFckjYwsYkVJ6SRrqH1PT73UT6RJu8
q1u+RpvXfhzMIGntlMq2HsKt5u9xsTDc+Aw9LouMbOVinyKs9tGb9dfwZclAs9yZjXUcBQnI75Ni
EexwWA3UEV+wjVXlHSK46pz4HodX+8+/8GUgEG9e4x6Dab8RRhLnPpsFJMgeLiTm7SmvaiQiUBKr
Sg4Kgj2UTEwj/3pQXExzFjsI0Z50jfRaSCROJ7k6OGwWt1dPS/v70Y6eHrjKtHAackF4OjXFwnPn
y6eeBHllL00gKIXDQ9nro2fKqjhM6Ts5dvQg4MBomgzSeGpLHPjm13SgccyXbd5Sv9BSu3LnQQjn
z8RTF7AODZ/j7HSfDCgGs73/0JgAqGY+pKPlnE5H0hJfyr5uyuD27fjBt4TlvNJE/hgOoWq4s2hA
lVbWiZcfTA7Ll7/oDUM7cBmRiKv3EY6PEIZel8kH5qN61lxOIe01BznfxQvu1IDkCZbxMIOWSncn
ytOOvLOyT2fieT1xt4AD3tYsVxSyfqFki3+QZTjTw+FCbfIOnWScABE05XF/SeTvS5k1zdPKAgtQ
xTa+bI34GEHBMOTRMFxfK8NV0Mc9MTAxoNBTCpwJBjymeu1rWDZBjKQC1GxL0dj1hBDwK6NwJxNv
yHWB5qXPUF9plrcItVzfCPNfDP07XyJl75dXdrhJxZUYeOhV5ilAak0idfiKlD3hsMKUb6/Py4l9
xrhm/Rry5OGBnLK2+mXdMdpcLqzrj9R0IQjL40l+/aurIbYySQN0cWD2QI4uF72+6qvUnikvVMdA
fsQjufZmREW0A2Gxp2szLmPTTaP6m5XDhi1g/h/Weo7/mAL9kL6Dvt89kDQOaiWm0ES8L73g/sza
ootkywZjtJQWuEmgjuxw5UHkVu/hIc8LPBgI9iJqd3O/wiRvpXl4lODb7pjiWvvrZFTKLwMT0AF+
yowt/BXLb7oQXqrM0+ge3UAzuuxNReJmhmCnxwRJgdkoTIzV181ImckvFNJt9th3zsiWEUrbf8ol
1dQ9SGjEim7fwrEDZnsrT/RLsb/qD68NG4ig0qnp00KccgnnMWh99ohr0WvnVxHTZb4Iti4JRgnV
DX2JThV1bkkSiDxVz1yHfxHLo7j2BUWj6WdnlU9tMwsAPMqd/EiPhdcwIS6W52f36YXaTqH1u1sj
l9pUoLarh+YH+VemBTRuqzPhUJEpdJIVVTJ6B9Uj2YrnVnEdukKkQ98nPZsASs3/TS1+HkQm2PTQ
8L1O9uzcLMSe+EXK7QUpYfoHkSCaliDlGQm1JeeBz/yppI4OTUr7zWT/lTJEhYy62036KFSXlNZ8
EUPWEYutGUTJKqkDNE1pv/GrAW+CYC7e5y/FY9OoRNOuBzG+jfmPhNMHp9542/yso/ALK5AMU/TT
mcvUm3I+KnoMvT4ay6J1Oa2MIMlDzETdH5uJi/2HxQBDZwAEcsaBv8YO04gM125aliV6DI1dQnwB
LqALWk+jwG2ztA+o0gEYbc0Pkoxj9pvVL+HrUzcyi5ZxM1UYjg3D2ZugZwrRK0DHZ9VFT99sd5hO
G+0jHYWfdde940kbRHvfJHv4LRuCjhhFoHChpo6MfQu4HhZmSnmFMbT5UXxO4VmaBQcByzr5pFZD
SRasvoFnWRtY7MpU/SarYdiWNvdaIKR+Hp0I7DJC+1SHXlR2AEQYG85GtofG1LFrDqkr3b7Co1Jh
fcIUfm8s5PXASXs/c2xP35R+wX1KPRAeJ+If/0DniDymc23CeDQQ66qhdeNP0am38gtZhWqWyq3Q
iBaa8QNYY9eX+PkqI0/hDDQtSNWETlS/HdQXbXLGqzjrxYwJfqdaj4x+ecXCmuOXqLb8w3ERo2IV
g726Y2BC/oqY2w4fJnzemUfz9ozCMn4adDtSWCvZUUyPepAUGorUmqsoHObkLDg2ksV1Pk8hRRfE
sFRBTmZ0t32jEV4ZU/BNpUkLvrUGFTlA+0QYaLuHeSLBXupUYx6HNtRmZsX7PSHifQ+rMm6anXn3
OqbHx0eMPf2KnMMLaOAPMstBbCn+Zj2iQLNDO6O9nVB8EuCoQpbobEPDWuQ8MmbNj7IncWajR9m7
IPnzUCn7BsiOcinvxnOKCDiQxd7h9PHjaWq5UXN3O7Mp9RB5Cm3L0A29o6C0B1O+CbCQLJIIes7I
RXA2L5UCK2DY0hcFied1og8DPT/9s1C0cbSZdxHvQRyICctdj7u9vyNd8QXjdeoX639S18exYwWM
oDogeaz67R6NrbDTAyUWrMlkloQ4+N8nLi4VsvzXYtcnj00bFNIHd5D8rrEuUWOEM1J0Ivm0Q9zR
XH+l+7c6OIxl+DYn3/LVaTh+oXk3EEAVvQZRh87/gxTiBqJc2qx4hGG7tXAK+ip7UiZXn8KE7MRg
BO+Rso/H7vTvac7JI4Kisevs+Igcz6ASCSfdrVuTxgx4vJXWqGXzjk/U6zs1EZGaCipAFdzOyIMM
i3mVvTkR01NEAm6oJHBHdzmVRxr7oYJZnmYZPa1bjwU93w/4j7mwNMBDv1ZzvjPsKUAasLV8AvrJ
2TvGK3ujrfCysIibII2D0OIzUGUF30hDWCeb00lkPbqBw+ek8arVllL0xqiU27t3vDMbFE8gXi66
LM9U8oLYZXD5JsMZrZzcuUXA1JzSklyPJ0Pi3GysPupynGwhPyx3egO2OUr4W+7DSQ4wVCbmKi8s
hIzSgh5LnhG2vaa4v/bK5froROJDTV2fCcq5EWbkBPI7rjcaZyn+o/IL9C1tlzd1dPOZz1McU1+F
1gcvReeyP2gp3ierDpXjup2L4dtgAdcgqY2tsJuII3aYAq8EFTmGJ7XjQuCyLpznY26qH/xWrnWB
q8DLfOgkTfY2tyar21zNloKrn2pPDcXGJ1kCYyz5Jrj2k4G/JWX3j4UtF4f1TOzJs5dalwR+JO+i
mB0K0lxCrtPyCDOyW8Mmm4femvw/t2/VvOtT7hXUXycQPC6bKlX20vlBSXxCWcuUP/M5U9egrZ37
btxEiDYo2yV/H0tQHflYkVveUlrxl1QeBDjiUdFb++uGKjqZa3d4hukl4vdr5k83c23uG62WOIfL
tvSaus6Q8hdkTy3EIJU+j76uSOsT3MBRzq0pucDjqfb7tDxzm3jWmIm1nnNyXTFzgOIoBQuA48TP
zZYfflU7QryCX+Ic+wNfNNxXs8rQNjVfB4tzU/bZz+6d0W+Koqy0mroEqB+duqpNMIX0riKUD/mj
L3O/6Kg6hejGl7ahVWRNiepDmaUF3TfFuJO9fHjUCyAxSljRNo4EdkBK4VrUuxsjvNfVj+MvbGw7
Fd4YQEMJc/v6x2n2fRT7y9QQqEH1EusDtFfQosOUVFRbgOTDLyC0rNtTXn0V5LxWPrdSCzIU5Gy+
E71Kq5p7CsuGazQfV+Oto/DlgEJ3WpuV55Jwgjhhu0MTq5gh08NCi/BF9yt7+npnmx2j1mjsf2x2
NISlBA0gHfVKkO9oHnFqplNn3S48c6rW6JDBsEV/VNRpnA5Qhc431Q6mNSL6n5feeJteIbhlN2jM
ipaNke/Gn9hd4Uk1qf+PHjojEGgfMgu5e63tK5TFHj855iCXkxkA6LlikuP5RdkP7zI6AS2quAn6
fQHtmTqL8Be4/DhZUeq458yhXVEGxo5P+9ehxpGt3TLNqjWs/VIqZLs5YzuZgaRHRBiAogOL1Rix
yO7HNe9qw2P6m5cNodDieGBV7eEXBfY346QC6OoQ0kMdwJc4trRF5kCRswCUeGdGwNg7BMJN7P6w
pyWABeR3ZJaF5WMXU4k+kLgCyTDzkcJ8J19j3m7P8JqBHlH3iUHljUXqB12e9eJxtqdC96IqQK1L
LfeHPFyJZwBAl6qGUGT5z2YWmTdTLWnbwVTj4GQScKXYKJLpZt9p6wo49wQmK4oeDI0/4Yz3HrOp
bzKeYcUea8Ewb6dFGUfUkzM0TNwRAH+urNxnb+RXGo2GFW8OoBtH+d0uy1LC07R5CvlMFc2Dexlv
7schHAN0Kst9xMMx6EXSu0hpDbutBcARJ/6ie4xZTV4dhigualVhgBvw9Gt27r7dK3L4Ud6/1WpV
fqcuCRXr1pOqSga73n3BHBzq4kw6Y+rgnUXnKl5TVgI8W2ffLhrdK3nV6P7bCMOiC1Z+PhU4Rtlk
6O/WkPExuJwh8Y1OxPoRSFHNI69vgB/SR4jImkqr9VXzIn8XubTY2TVXfFEq9mOSWS2+ePSECLpS
OliKLZJGUKPSQA8Qm5tHcfwEx+eBAREaeCi/oC3vUDOcvNQMPpitiNqCVERZYpTyYSGiNORs3PSa
cui+pWRezrwTClL0ZjqxcqeDAb2cHW69rEVwM80iWrq1SKh9tboqALn9hTVvkqpO8mKipVxx1+pJ
gUYVJv1FtLkgzB42bfN/5/uhcPOWixXTTQYRBRra/viRLMCMX2p9FCKLF9aEnCGIwx5P/SOb8sHc
GpLHwiOrpvpeAeB+Vryj4yE/z82Yiz2/iCEiiJjjdDOKkpv07dQa6da7xcaeWtFKod6+l+RbXWx+
iI9vYl5nqiWAL5JLbB5E9R9rdqxCsOYFtj8PVhfYZp1treFGpPYX6a3Uivtd5/svIPyb1IzKIFH/
bfY/7xPjflUQn+lI3mCYqSEtSuRhyExHMsgBPHjoQQ8rZaxcUU2/lujc32r0E1l58FC9oWvQzs8D
Kl+QUq8DqtawvViFNvJEkkXZlEu8IbsPmjdzFc3ETXgdRED7jmAqy4LwY/bp+l38seO+c4t2ULqh
DfvuJFVNLaVjt55ZGHIGQkLuWt921R+CmGXo2EjoSj7nwf+NFLiPK7cE+JdP8SqpEL2r9ji8frto
qpW7nwjkjm97veP8gDj+AsGrBM8x65n6nWKSbiolZFdZ2j192GCKCto36yTLdlGSMAFWvLtm1RnD
dtXiXKVQvwQKHyxSqahJdAu+QUU8fo8tydj0rFkcOnwW+z6Y6H1gDYxOv2XKo5OczrMbIlQAPX9v
e3UiG6vjkqGFgLqo1N/ZxJd1VGCz0eyO5DjTEJNfa+fkr491+YiaRFYISLTZpLapslp25RFL0ZVQ
S20IQ0lpa0x/6eZyge+n2O6t0j5xapfkd9zOg93JjQRAUWo2rrLKpX5O9DGlaGz1Ml4QLygSwwmh
x3Ol1T/yWZAXBfkfqj0Jm+wkym8MBr/47pdk+Bnx6s8/tFZKl55a/7+q5u9OmE1fFL+ukOciUraS
1TdONT3vIMzx4lcFFAYY1EI/5/TtP35x1D9aZrE8MWN9UXya3gCaJm8H+RLEBespzOHI6GCGxSC7
rGRk8DoSl/7qwsLribYO0eA9uA4OI5hqQPudh66Hky5OVi9iO5yoHcPvkU3D0dfjSZabhtQ99ZAC
7bMV0ecr/s93FGkPp4AHGVKVG1O9oHIj5Z9KrhpDk7DUZKFlVLYJyO4LLKjR+JzQPSddp+uxzw0x
KJEQipb+Kgj1Fmr5R0x6RQ1pWkW2dpU6etCjBcShNJQeHSMXttT+vvliQmdZhtX2BViCdsV7ptlt
pg0pavwhrNM6INue7LUhhzaO/VnxYA9TYO0DNaCcq84bV11UH6zLgH8KgltXlgz/QE0oCNmsEpEm
VRnCKii/DAjgVLjXEgv2BasT+00UER//hzFYD6gXuM89qABQMNc43Ia9bSMbjfoegBdRw15EnVCH
xAe9YbPjFFf0b76TI+T8K/shgfNvIRVyBn/5eakcjweY6hkkAfsXKbTR/HtfN3LyUgY5B/XzCJ5H
oFyzpEnq3wWsJrWS5rL4nCq2asLP7QfobG7oZ0pziF9PjbDuyOOvFxoD61yfmPX5Qyz92VEQ0/Pv
wwpw0eQX5GuDENHvmFSFnVTqZd6/1y56nVqKhVxgJ/32u9Yf4YTNAefns5qu5yqZSGmG+Plv5MLQ
RdRThmxCdCjKJx92EcQAtROq5bxgdH3riUuMVjRCy/0ceBE31c7l+/7XE4t3pqgCK130784T50q7
S57a2LIvErThrFTcGjX7NyvtZfnjBUsjG49aOx5Nd6NY0h7yJPqxR9KrUYWTv6/q5T0fNHkOEcRN
HbrywGWbEYW3vF0vrGuu387n8scTs4nHVGGMU20kKNC6+Uw5Y5OFNpBe1bAMdARfKmGQMOGcXK9U
P6xwS4Kld+4mHXGSd+bPf68oXzL5vMDYZH/P5NNJNkg+3Gav/746S6jWoMs3zgz6UAr3GBwpuJgB
CSpXA0xlusY5yiODR4wQpZztkC/cqEQkVJCXWf45FtI8SUof+qgfgVZbUIGSpp2YIVNJZq71fFU1
0BXbQuJcQzphhCBJvpnQiuyJytFcISzgKg9SXJlrWPf9JH2MSI58qJEEI/kgy+euwgaZexiraSBZ
unxb2sHHvg+ontaJK+9KzeA9isFS5cTkzPx+VPXc7EwyGBARK67TOpcq17WbntiVGOdRfY5fXapn
I7EXHG4S/q53f5M+m7JopZg4lXHn+x2UQ/VMcNeiwZWJWmtg5NtYdvi+ibbxlLz7+1BI8kW3G0J1
lccMgkGsBdEpYBRDvAHYLQ3EKF89bYqkJHFtJ7exXepdqu17cxkQxpftkMvqFyNtaX6yoknHNyJ6
J70ZdAw5edyXqagHoSdRLPWfOTOwN/0GOcV2V0JpElyfrd40MvQlmair2IUHJCS/vPTJsOyRKIKA
TOQ+tpzqUI44jWYekPq4dxjvuqB2/86rXNIHpREOLgZi8MID3dzRnJvyvvX6ScvzNCd0h+kCe5Qe
4irL2gokkccGmJkkI0ai+VzcAvrWbGF3z8XKnsCBTaO9oo8xY/FGBfbDJIjUH/mNyOgVwJvUpuJo
vzLO7GO6eALM5c7Vu0AEV01LdTljSVKG1cbQr02xTM73/PPlAkHiLktx5GJS5cb4DGKF93vz6/4O
eHLNEa8zVc3W1T/7OXz4pACVqmNDDsfNwZM2zGTEFzuT8aseNq0fDBzGDoydLeUaoV0ULmXHkYFd
LW6tvmFmK97+RRCeu54w1w+bB8uevS39EdVNBSiF4Vpl/PVBSdaGhY+kzORm/2lcHAJwi9XS0VMW
2vpeqVIZLAdUwuNMvx88xjt9MdJkqwhSYATNXMmCea0zmLjWG7Zj80NjffaRz67pMh43A+iNSKWD
bqDi/Hi1LJVosrcaJZp1h19R4sAuCzGOC4iztsS4LZLD4+vFaY418Rr7/hD1Tjx+jOJ5czUovyEX
ud8p69emA55oHCQZ3H+OjkXB6ToWu3uBXDTgIjehm+EO0XwksjcoZsPybrxsdZe5Ad+0bIGWXwCg
bQwSAL+N3PIGg0lQhwHWNo0O39sL3UAzgKyUzB/iH1LvBPaVtvwEsOGzg3XuWuyJREKXwFaokg9l
yAHF7lNzTX1RThkv/SvjNW4/D+CtkXCPqzV3ATg+QFCzEKOphhCPdGRQ/3q7JthNVQjKRGG43kMa
/G5HDZn/EaA5XYivWg1Yv04jaA2m/Xuh/aSx2lFmByacSHuTqmWer8ZVvoJMF87n0Hqxv3pU5T75
/VgwZ2oCeZAyWtOQ0Pd82NaL0jNeVohJwrk8ZFkQ5rF7ZEzyuRRIRYBc4QY8V3X84ja2LlKpxmN6
ndL9Xm0RprhKH15uW/VdV7IIkkPhWgdu+GbHSpILXMrA8eloIVX2Z2sL23uwr04/yeauWZT1mz77
i86pdT/wf08cyKH/PLodjErTs2mON6PB213OrurUD8GK1nWIZNXb9MTyNM0jvWL/mGQfMvKsEM26
F5yMI+NfEeOWppISMBW7nMnY3k0QWDx/o/hQ9dl8nLenI7AcAvVzrzO1Lv3e2lwQzV53oEniEj06
26feIvD4/x8Jn9iEw/HI0kfx+IBnSH7Kc0ZDLg6NLiu1PBPnXjUiei0rhYqlZapc+y5dD7MK7upo
DgTs0Qpsl3TPqBl81NJptbYl2MCYHcEf1ri0ZaLFEuT5/kKkwG6QeJiccQBstUuw9xfRahhNh0n2
zFaKScHA76OgpoiF1y9jR8EN3lypzHvJ/Bc8xLLTp3rIJiPrXB7Ke/zdpeItkiHU+LAePvMmOHJ8
2vhzi6Fp+ZXjZ7sQ8y8Bv+fXT2A8A9bUlxMcki2CmlCw+drqa71nH1IDeGnOT4q8ZhqVq2CLwjeL
MF76WkRo/HJugBh1TvaEfM/X+HC/jnMAdTrGBq+MHk/sh0jcoWHnvKGuA8wfvWfvAmxatNyWhvW6
g2XsTLCoIfHaJ1RaaE7H0OTDOMd9o+WjDegkudASrLW8YvH1oo0qBecWCCe+Js76cXNNygXvnlyQ
pIYjeg938QpsZmkqunh5Tb30JcFH5UQj1ZT0HaTNj3F/199YNEo3qpgA3RRqwVmIA4x9oP/fk7gn
lnHXJwFVAzEUMCsL+ry0N1E4Zq5k9Fatc1hvcLBp7kdwNxHJXUNkyypy2A12KJ0//XS7PupdhQjt
V+jEl56QB3ViZVKjSMD3YmB1+VzcRejvPG1BU7mFUun82Pnuou8kF4/F2aR9TjT6L6BL4YS+gfVH
RHhsdmBxDe0MVZt09efJCJTIflNU5WEvpURhCj+qBVQoDnkG5+llXJxMuLmd05K+liFW9X3TjizV
P2gzzuEgc2v4h7akD8rVZFuw9PrwZBMJwn4fPCchB7tiiUK9CwZ6Jo4h54/LEH9t2W2TSLXLMO3z
BkcJhcvaJngd3s5FtcqOGkmhzT7XDpG50qBCMuKliJOxBTm3OMFOr6MH+DuUzOcBtG1Vqigy340Z
tzm2A/IjvnjP4bMVKt098CE6Y93X8HkBsT7htf5zILLqQqXSIOWiwTlp1BdqWJuZnvHN19h+zvgg
yhXX5adVDqW20n70LiSc/jMKbl5us00Kjul6bH5nRcL85XunJG7gHlWzNZ2Zd5Xh+m1fmQQVdu5V
s+CQBmPmYvMRdblOoG7owj/7vmWa+VUi2y254shKRuzC+zYmenSuQo/2RbMWC0quZe4vgBEAySD2
nsQM/GkKNyEp68TbH8jQa5I7YA3701gL9jjxk0Z7fEa5illlEZI1xcGUEM3iJGioReSTgRH58zFL
35ItrTrVsqICEYru2gIptBx7sYYuzAel0gsGQ6pa/L1oFK59ekwTg61FjfTooirb0SKwlcesTkyn
jn9tl7rlKrXDR3X9Qauq96eTLgZIPChAliHoZyNSIxrVKRGIzV20rxdgUL7UwkOTAh6BPhwDDtD3
hYFnjhg1sq+n+buA3zSeZKGBqLVm8PSBlVB0CXAMB32J81KR8SiEOfzhSJJn0/ag3f9h+XXr3ZVG
DyqKSdl95LNO2dCp6BodLFG4TBa2BKb7jyZqWqf4BKQ7y3uu7l34ot18yBwJEODRH3ItmGZ2KfNS
oHTi8XjuXdtQPvTJTJ4xzUPpxE6iyRQq9+dxewj2jbF7gEp00NZkdp5cfUYqmalhnTr9LnpJiZFr
McZb2sffVmcw1IfAtxUgJsF68mjeMlCc+CudD+Y9UNQwahvFf7xwlHRvlMRybefRkgpL3Ve9shwV
2SbQV1Thshm36AIkULKYfTR/P7suyQ2e81SS5T2JdpUu0y3u4H6c0YZQeBTa/WpPZi/eKkxXoA++
o0M/HRu5PvzFup7B0im8oemVhYgimkp+kKSgsva17u4hxY2uph2knGNjk0gd+7wABEiTmJ4n7mLw
kG05yl9dkK7WIdiqkoxUzk0rQpDWPdMd4sik8/IeVduJMRuQBs4HWKVPHv6ToGQYrPLOCQqqabx2
o707crH9v460aMUgK3OL57tUo7BpHOxXCwF+/cOkZGbsc1rWNumvVLwN+bN3z13ctTRoKDdSNLwV
Bg+B8STVGJR9XPQ78v5eMTwKMsatIQUDw84n47G8xeqbOI2ISk4EjxZGfrvuUlZ8D2m6PKXRfDWz
Q5d7w0OXD7FWvrrN8vB3TEnSreClBt895yp9uSl8icsnyg347OthTQIOLn0RWz5BmYmt/D43h2up
DPUPcy6RUpuFFuMdzjGyEXqTy+gPaqQp/GecXT8UxQQrW2PD2ej6EcDMRJecYTwEKpFvJNzKe6vK
PSH/AtePzakv1ukq8uCWVk4g8/1DH+itJ3UUxqEkuxotF6EkZA+plW6EvaNocFN46Ey2I7CMY+bh
8jaydVVmn7jzvBSxm9G7b0rgMWyRxzuIoNQ+0wLe3PMZkr5lwrofV2yMqerr4aQcbufxdmj3L6WS
wbbtmj+gxQSQFQRtMdihDSP7dpO/VPwPTaeJIp5zkY6tAzr/xDZbZEKHDN1nyVsVgQxYYiGiUZxB
dVOhQXR2dkGDVVEObMTKjWDeK9hTo3u+TouknNRCHXcrfrFPmBFz2h8fTjTX2tOISXBWTa3SSNTX
e3IhQc5Hg6vr2n5OVyLKpEcdNWGauc0lYfWcGmlsMQg69XdJGL6NeMtPPiRERJZgkkSzL0rv0W20
7DAnmGgL8RyxMmPjnJolb0fwCPakeYIdwwLMk8Lu1fG5PS7relkIfjNU95R411biAQIs9PCfOL2z
3T8E84ajHqqXPDxQE7PnOwBawJKon1QrqofN9pwm7qCvplXKxj3Y4zRcRyXLS2YOiCbrm+GUfWLg
kb/XdpK0Y4TAkYXyGu7yq/7Ps938BpwiJQxsqUvrDzbqaGpgLQWzapaYHh/70KVfFfihwjjxkJRv
8J3qR+OMY7S91Mrz+VdP66LkaFt85IKb6VUBHDB7FPEeNLJT8RsU4hnQp4T6xEfrxtSQVO8kJdHi
WxH4aJ43Z6tdI+cBijJOjwGUy1Cgzdehf5PAtW7/Gw7Jw7R4rzAlq3dUrVSialxV7pdCIfMVND6K
gpn9+l3jUAjBGaPNY46uRVF1Lwj6VscikEEcClXnOm08IeNamycvK+Mw+MwarIqdbwwwwRj72qWp
FjnuM3EKgJlK5GhSrP4v+XmhCEsbbK9CQiX6FC+K+VsvjC7RdekxdAdlQCGEMbNYsKPWWSe1URTS
fdYSiKmjg80vFvND4XBE9nh+pnQBQ+cO+fi0Vy4X2vLiqaBlxlH3gIrSiJimEy8H9BoUhJBy43H0
V8IZZ2rgaIQtEx+7/slP2kls9eKM4kk3l1cCRddbaOchl1VcPUgPXuh3FKRYekxgj1BmYr+7TfoE
5gfm17/2fIJ34n9gX6/pkY5XG9VYAhM57LH8zP/Znpbj2wGAAYY3RLD4I0N1oldeDFalaL1mF6Lp
gi2WKmiZc6WbHMynWaN4XVkPAhVLbV43Rc2QrJ1zRK1nPxZMVfUrob0V9OYWKagNFt2vBRb63ugK
SVwm2ADLjVSx8Z1CeBU+guFJmzMVFIdr8/vgAAR9Nyfc7/6jpjUpe30ASBEecY+QArVcfDfYe2wJ
5nxBe6ralYsJpNsgbWtHqzL2nprgarPcL1bSXWaPE5Xd3dge/05Y4d+u8cHtfVHrYoO8rXLxH3fv
Ib415kCnn/6582eWa6TrO22OErf3Wy7uKPhp3dz3LdN3ZpiQrj5T423mU1Ilv4ykCCnLy9f73Bc/
ggFTajaU6XVZtikcX0Rj4kmiEVTHBgaV8inltN52RCOxxupHqrYb/Uwj9LEY8BaWwJ9STOz2z+XX
u5oa4YTgwJkZTNXTIH46ll9s3PCT6h5ycIMPg/X4/mvn040jK1GWobdzmaVPpqFSMHRxVohmKFA5
Ff423g8UbzPGzWhgZXGQz3mr0JMXnEvxmMXcvK0TmRkiIrIkhOSNpdn3M1yCNtKfJu0lBZ6WFrJG
BveunNyBg9hW+es7CGh94/roju+rjVYuhKAgv6/UVfyejU25kwiY32CFVCtrBJraOyJauKuenQeI
3wNyDzsCwnzE6pXpF9wndYD7u53LH9YYg9oZBvtngpVjk+eonAIouIuA6db0o2Auzsiz+SvktgQB
ydfZ//4vsdmQrqrlSaheIwrSR7LOenhw1YlhdAYI1Joco0vcfqHCg5fYyfsFBW83NeCepg3hAbY7
lkoAOP1qlY0cYw7FA0PXbQDeFcUeVl5oOI1cyjrsTTH7d5bldqs6nRDeQtcINHFmV/MyjLdLT642
dfMi4dkQ/AVqPMaTKJ6N6KUY7ztUiDRqG0E6yTVEpbnB5fS4MYoSxH3+4Wziu5FZrv6gQpB5VbV6
KtOqTR8qqyYpJ4h8K/uQl2zErJzoPTf7IVXt/6Y/xU2m2vfI9dCS0Mp1nJ4zmtH6liSZ3VKYwhMy
gkduibOoPGchguLwpzoTsSoK2grfg44tMZ6x/Od+onZ5N2eaIAghXcGQQ101GoWRzPz8zlPPvAcc
blSfBOVDO9b5D78GE8EFrTrc8a5GjZ2IY23GWFJJRIhA730Ux+8x6TbiqDtuB+0UQJa+jajSBeVa
BFBfI8T0+MQz/orknYWelxcM3kPCIH8Hohp4PhPF1EBbnIKoqrt6UwaB1MHBlNiSLDdqzFYOpYve
z3ROR7/hSuEE+ZytKM8GYs5eOTmfGd7JUXdicfSWWpjLLYYREFgwW5gMxQribQ62cdRQUqZclHd6
Cu5x2lPXethe2Yxuh4LiX+3FwROqjcQS0917MBQddW29/REuZ10dAxrHThHf8O7wLI46Bwtm2CY6
wzgQLvqAPsAzMg/l/vXgz0SLwWHVqERem7k9hBPnFCF5uxiReyMAgWurAMQDc+WmeqKNWiCWwKjV
kiY2IExMapSnfo/qYMiSgY+spz/t2Yn/EVFlWegL4JsZLcCpAVSA3hx0J04DXjUzzXhh8L+Uc1Qf
BZ70Ayt2eub6XKtmjKtGyIfXJv2tJmsGcyijuFPI2IV7Q6TlQOby/ivIwEy4bsfISM0Z9lY4jpOz
oU/y4WFM6v7DHHr4iiYkeQuP9BBox4oHrPlelPmv88XTaoCcX1x+q9QtJszx78hjHHV+novgsM5v
cuKHudVn1bjYy1c5vSRAWAZjjQ9IsPXmdX34gZpMYQZQp/4gFgS6rFHGGy8G7wfp4Y2NeyhvSESd
vya0kpwBEi5zNylGUWiVofhHUz5PPs0ABQSNdjkXOHmGIPZEH3XCbSlEnvu3PQfycbwTxMKdWG9n
IzvimvqEFcS2GxsCLGOzglmcKtXG7rQxVkS5m5IcUpt1/frentnu4L0ed3pE/G8A2cTBPE5EG+4H
Q32fV9nDUi9ESnVJ24fL5MrBb8tvR0ZhAAvfW+NgzRNg5lH+1PFfW4YfUo3McA1rDSuzRYJKXSRC
UB86krVlIesNArgHQEG4SUzMiCW6i4INwyfh33efDHVIf26qAVBuj79jxo5QqAlr5byTZ6kM3Y5m
Qc5MaId+gXy0ZlZwsrG7e9bsdjg7wHiXEIMwd8pLku4LK16RH49pJsB6rDkbErdrVsheC7T4EX2j
1i7lqiZZPYrHOP5PZKzQaSxkbc9Bo6xl9D+ewV0HgWGVORvlVQ966Jzbn4xd4fMoh4BEdSvxM9sK
fctTh2uPGAxB/M+zFPRjnf063+L4ydZaNu6YW7O/CfNEWrECw43TC3bh+o58WhF/NMOhQ1tDHa0X
EjBLOExv9lFXZdh4GaptDUCqWVGInhM3UvlGUzm4OwQKTO5G1Ie3yzLh6Igm7f+/HcAviXWNJl/q
Pf3lO0M5J6DAOJ7QVCeTmfTiW5XzWNqwoYQAokEWEUKOUEIeMTZQxBury1pKyc7wjxQTItXVPQUr
ZwD/BvItBOfaPIqaslv4QOSo/2CDrHqlroc4F12U62Ctd4j9LvFFFFtRlqsfAvMslyjvFihf3kmD
Qvx5zNzbA0u66KbjFj/6oQX+/QWs460X8jkFHXxVQ8Yy/04neT9rkcrOkdK/SVcfUW+YXXBHf0Lm
kDaw5Lgj2b+is6VmhoXLyI5JHGeSrZi3ZMQaWCWGDzH/AUTaFHE3R+2JSh4FPWPRjXG/nqKEaG2H
IhHSiKun5uxGBqAxUmyQrCA84U0/8UuLEPo5tyOypjVZXETzFm2pXDjLPSomsZYXEokxT23abzL1
g73BcD5OtjKhialGXuzzOwvztTVkOWhbrolb3ERFoHbWSKcLOGdlggrgitfyg7zCVxF5syGhacAC
7WyiWH/tzel2yiLTg+iHDErEPWPNXk8T/fcjx0Yl8iz99fu3OWJEe92JuMikn5QznQABXiLYTjDi
IgHyZ7JPgSyH7NuzzjHuOUxFFDLr7c/aTFY//MofSD6Uj6nWPc3WllpnakJaiMlcBY89/4bnUWYC
iTGRv+hXa85oUTe9r09Vd8kOjk9tRZr4weNUMKydZO2gj2S+YUxJJT7ViGfq7xGA6CV459Vop8OA
0diAPVnBllC9Iz7sI6lSuJlbxL704TADYK+O+E3FhD+NO3CXw/hZDUXlI00pvPdURI3cbSDgNJUS
/gFU1YzGEByy5saYzYdrnDXKjCEynjuce327N/V5knXELJj90Ys8TWse5xmydlbHVuURlFjDmmtb
vYLrXWUz4EB/u8YXDSJ+tWOismn8un8fs0GXkFN4uOFssNoR4wjV5Fd75v9u5NAYswA0c+zbTDiG
WLtWDx5t1hFC0coMceYBQEIUHCClZgQg3eUwoGRNjRJOxJzmXiPE5HCfieS/yKQ5xJWYGLOZE9Xr
68vbHhmxpalGWqevLbyLVMCIhOCeYHeGKN1NjfCjhpEClKPrGVKSWpYDYreYxx08fmATvNQuhpE7
wQGGVASiFHwrSD9RBNS1K6rn0HC/vEetZrvUlv5txOcLLSNY/VyqGG3ok4CpzzGI+Yf8qGF4EMQl
OR50wd3xOQxc/IMZE/C8tZ/4mUkRttbPU7IufB8DLUac+mmxrICTrEgkbztumF7kaUNHORFsRQxV
CKDt3I9dDl6I91KGeU3KwpPsHi4do17N4u3MGU56AAIP7hA4fIXlxgUGoyB7Q2IsW+m7yunx9+4X
YYIa3kBjzCBhRAAG+WxJ00fgTShwiO34Tec4ITz+4XeIz18Zbnsvx0ZE3kvEb9NSX3hfHMBjvMUP
fyb4A7rrAFRWwgx5DVtr1KAIvAnkmGZ8nufO3McV+uyzP0dY1VCmBegD3spJ+JgXGQbGiV1GdX71
JAWfcqR8Bvu9uZ4pwvBnUcATYCGFjFjcnb/euCC8kycuF/401YbTD483YNvZXMs/nW9zv2lsFNsD
OH2rv7Au8MFBRuMnw/K3jByI+jhLGtdh/iyyNYOCARtxAhkvx9JBKogJvSsnh7wlcu0B6XNm2hMF
1hjP8DDRVaVgANc/HcUZHZw9h8FqUNZvINU0+bJpAcxK4YncBZtJQsbFPtkJULK4uq/GKPBQmTIh
VH/Vf/Rb5DN90rTc6Z59vXtBXv9QSwYmugGZ1aljbISCeQ6DpnNRmp1S9YD7fyZvdB1dTmgFoDf4
shiBwRnNc21k7kZBbawfRLuCO52A38HtMYj87lVrEmsEGX8p8UezChm925Q/FssIlF9Quryxdq3T
5MeL2Sz7Xsu6w767kUY/XebH4kjhkFUnM/STUn/ruNnoepW2aXQIYgsvUyWhTUPJCf84cuTyV+pb
TGZDzYXyD0pruKeu+DbK7Lh4oHu3JR69Lyb1w5LzJx+YfuhVK5OJOdxA3FIy+hfV3Bu2lACUK/5d
1+4kzEQg7V8NzQ+XL0BsNWGQbcMU9MQvKdRspjoYkb84/RftPR9ee69rSkYO9fMJ5kMqNqVtb59K
D/Fs83FZtOoigmk08ycTVYjCCPcD4wPUz0TcrASGVl7XVPgVUYv9o7n8I9TtzszZqrYxJSnMURNl
LXPdEDWkXPbjNkJqyd3Zuzcg29QeSHzqR32oO426WM/CeuJo/ORIQNiGbes8Ki0ym947MeX0e3Pe
qDeCmEC0RH7pr33ELENH08sjyyrtQ6Mxh3N3clRuU5rw4iqqHvf6s2zxwll/OgYOL3iCEnqUmpdQ
v8j954/8WffdT9an5BISz38InT2EXxJwLxmlmvbPb1GwwvqOna6oDueLCbaeCXklqfvfsFcfFyxq
e3NoTyXgp/A2y8fCF4+e0VcUmpRmReLcyce24VkHJ+EW/MLHwd9YiYV2zUVKafon7xYECpfaDV2l
6mtnuTM7t5xMb1gc7C5kJCKDuk+ymhVp3Y5e7LqESxKmuux/Vsr+AijfJLemsuRSQNI8XZtr1CKz
yd1z4mU7vv1iKyKOhVYguhp1lAYiX4T7G2sVUxVhQmPYiqYytd/hIKD7VucQFKzTE/WZ8kybzUVO
Z6ssTlWMiyhTzoZFczPnmDHF+xOqeld0ApaOQt4IxCIYy5y217fXNbJwBiafyiliD8Ovei60G1E/
dHg6/D+rD7Ci0zfMiXjLmQWqpH2zH9J28CAJVob/+YabBeUCxgJULVugIZm+6Tpew56jZaQshdGl
OikSAwVETlFZYckonMh0mQ/V0w+nj5tuqq2INpCj+fHVt483NFy7ALF4KShgc6mdRmGphkxgjbHF
xZ4EMrYAEu/qrKGhlP/t8V5dTcXH6QKX6I6YxXcqCB34lHXSYIm74K1FEiElsm/p5SZIQsAZ99Dy
yI2EAScrQX40UOw8Db35e1klcCrs2khM+w/4KVA2xEkT6tTaN6ND7qPa4OumbfmmE2dgqrjZv/cx
xBsr1bDpf/I/CbVPcbV0GGoiPFzjvjTRSieCduDFbzKCya8Fd95VlTBe1NTackObxGAM5J/ljm6K
76fJ9O9Alhkdo46Nh4z89aZzbM2ujyW5RCc5ADgkVl8ztqUooCPYGKWYUPD0FEb+BDIKFY9CKXGf
0Gcok683LjyWx7ks1qwKRk47MmR/1XK+/wPdDAGBXi1f+IuT2rumO5efO4c4Vt+AtQBwBxRFWbzb
XT66iRaxAQscSmdzKz1DPl4RIHUMjcrIcF69hDQ3Ut6yYfAkNLdbm9HqMX9CjMDmHYvt7mvzEAyt
Cick1AuEmSEF2RPF2ZlvjFFOzGVKw4P37vhSlVpix6sjBigMfpXVF2DQkMmowcnYVu8TUNLsDg7N
acdCjp9bZN3wDUetdlDmX57GrtVl2lylsuvoi7b1PLGbdYSt66n9QEXWq/BZY/6ObItOdfV72VZm
zHgIvCSVsZuFyCH+oQ7gKNLKgIwKw3dz5Z1YPvhOdCEufnxwtTP5qdogSUZieDsLLmeOtde36Omx
u0B6L4vEqHH4ldDl1W0Ux1cZ9ygEgEhhVlIrSnd88krOLtx57nBjY1kzr6skgbjrKzx1My1kwEdL
AWqYmOWJ/n404M0H3IO88HYpYI1qC7Jl9lAAQqdyK6n5wl974VTX1O0MetPxf+EOqAdqVFFqlAG7
6r3BkrizPPmWPcaGWAbZ3yZoq1vGM0fMSbCfY+LoKP/smro5olhUszGwcqEnlq+i5QjRB3fwzmZe
HaEBfSALim++5kVONQbed+kh0hkO6/FE0BMlAviFy8rY6fjowaZTqcaANSny/Lo5fqaRlDOzj0v3
extmRa0/81oV9vRu0n1rg+khUWkGoHN+zZy02KKtULCFDq/BMCuqrvE7V2ftCB5xd799VZo6kuhq
peGBsftc6R5GWJ5+uay7ZwOyd7w0nmNgbn9yGtAeY6rwudWZBXIiLB7EI0OuOteCkMkHRv6QHK7U
4CuWFME9pq0/3+SDYYE9hQDYjFiYxcMlYTzOJ5UNIvLhS0rBySZeot4AbqN3M/fsy2l/ZTz0telo
OhPKXuHeLs92MNfKea92jx5d6bRczUi+fmsTdQUBkercH9x0yKDe/O0dyd/LyTbZdSUHMa4OLhGi
UFemmwHSUbOyjyP+p6ROwYmhFNoyqGMaMK0bVdnL76uXN6+cbML/4uXjPwEnI8G2sSTKGP944Fkn
s5xPHK7jQnxLkTMpzOaHSK/uIMLMgT72pMQuB0YKoJVDFdvyeH38bOPqnwq7YYxI1RydFVa8oqXq
dWV47pyGaFMMxE+OnyFJKtVxfYpaVEWS6zx2Bs83uEyIdxKgFF4FziN2VNm8i3jTkaLK6xS2tJif
0Fjejg/VWGFbHDEkRnK1vQpZhV+BSdIO0391/I9jIi/Tf6JAVQy0FhJokZG8Sb+B4NRDOa4HwFrO
9x5/iLTZJ/9l2tysFrPhiWCTEuGEfi+kM4VECnLJvRsBsT33QHr1EVDeN41Tshyh2g7bLuBcENTv
dVpygGmfVkukzR4Nkrw4xYBarP2iQqfEMcKgBXbstWvuM/zpOXFi1G2+VYjMZwo2oOaA5cdlXmfR
0T/XW42VdA77nvhTLGaVJOiQi4lZ6Nu9zIE3MsgGMhbMEtfk1qHIY0bGbEFpaQxVP4s31rnF32Sn
DV1bKS/WKE9ZQ5EJ76ZjrYIVn0cA2L4t5F/znqbQDzywsNjlxSTcs+4fWegvsIYiY5qD/optRHIk
RpRyyFS9hweLyRFow9Xw6GHY2nHsVtx2L1QRoi9wH8CwktBLAKdF5Jpal4E4mUK2obpyq0riKcs8
qmj6nz8hcdY20dI+UjJKrw7x1nI/yBhWjZiLVlEYCndyxO30olo+d+EKaVVs0VXIuXTJmikFgYYP
n3mzRjbTJ2tXsovxZ0Bv1zHkwadK5pqqsJYXlFcNII2BKwNfL2XAlmb6/KDdHPQp42u/bFyoDS/p
+bSukS5POJb7VAg2dr78NGg3k9UNZChjDJyCQynrbWF6wvX2BgdPApRSXXJynxjNFDdBtwafe326
6Uq/la+cjV4qNdOD2m3B258t+yeeu/VmTFKvM7ys/OolLB5bqS8/TfHqaT19m7BaqKjOes8DlMH7
Tj9dp7XGikPPdeRIN6gvY4sjStppuYnmWNW3A2ffrvVREE73JqQI/zqpRXsXqPJ3ExO5pmPhVhNd
4jCRo+4WU8uCr3snYm0IFjegVtwKSIroCP2dx3Amit1Cxxy4Plwqke3Uu8RJqyUap8XeOFA28J2s
12aeqJ7RRKq4s5CDkmHmmOEaf3b8yQsmfSYmgGAXygz5JSjZQ+aBC9d3ff72DgxOjqK0m3vHG1AX
cyjuuqF2egZAez3W9u8vPnrY1aldSCeAq3/RWULqsBLRVsbBJAU9LuAB3+pfm/fhhflC5j9UiWWF
MT4rTqukfo0zEDaWNMnrATKo0gZSHU43M139MgCaZ5JuhKVXrxdiEUZNuJwpeIcxR1C57wPAlySW
ArBWADWxeAWas5XGFX34oOjQs7ytczDNGp5Vk5NWi5BPvG/PDPhEwVvFwsuFOF/bHoqw9hUIwvGJ
+l7bd1TRx3BZFWWnjvoDJRf0I9R69N7q9hhWVQTFoq3P7OStD9SrCG7v226S7b5on2UW/4766LK/
eYwp4mt2cGm+JVy65S8dpmZWyQtpUGjpAadhgNia5HvR5ey6f9C54qx8dWXusrNSfHtFRCZPgefB
r5jDuL5n7E12MYen5DuB0Shfac1miCU3pV4EoP/2kwdDYIlBbrwpX8YMYHYjpnpYxnnau861BICF
JlKj8GZjheFShUGsPcC1Mst9GkIxS3eKcFA6+/e/hF7Uj+475Ih8UBRSwF+pCqsgMejIKxZFrC3m
CfD+05vTN2fCa3xASGo+uIJhx0MVEPbhmQVjLOwSrcayJW+VJbNnde2PovxkBf77PVdQmsHZufC2
rOz+dyVwMkmmNJp6b68L0oiFClhdzNFIwNrdsiXtMIrOHOZ4lSNSBzqHp1FZhQWtd+1YJmpiIHYL
EWhXK9Rndl+JKDN3ZhXBdJu6ORpVNQ1j+ChMBxHipZQg7gXUO7SwMO7pm7O1cgy1nLQgh59WVLu/
28oKH+qkZvl+JmX9Xd6ExRWaLx98fP0q1KvmeVgO48tACY7Y/VqDY6S08MrORQ7DunS0FZL/xJop
ltK4Jmt0inrey9V8urIuUV28jGjHcv2mHeCQRJBquWKkKz4QV3w5/T24pxrYsFGBBRcXdLY2g1m6
uBdgetlynjJAyjTcPIp1gG8vf6TYn9yQXKgtYaPgpeTLf2+1dY6GCRjX0aBafRu39BivwBrAX+Xp
AcJGakWwrVhWlBxYOeabRRRKS+RehQIMFkGYgd+R5LvNaawEpIZIQV9Hw0WoogYEgAmLj8RsrA+Z
ct8J+Omn5G8yA5b13YmjlaT+SJyUzMTK1TgselCo10AnPThz5QWATXKN9y5E5CMjX0qabd23MSfP
EXqiPCBTNDBBO28SsONCKiT2/YprdICA79d/bjZB2NR//zW3xIOobo6vq8uTtaAh5lb+SthzmRsK
EgifA5F2H36X5EyZUeAbWn743RYX3LE3GQXmn6z0rCOKKgO8cKs11AYtkI3oP81BuS/e+K/3loah
TdxBJCoEXS0hyhyxuiLECqqgY41mEvPaKzM49g5B0nZt+/hU3dWlqdXqrzsiHFaLy65St6orSOtS
DQ41FgJiHFM3L/sEIJJD/EUQF2GHk8W0NQ80adR3bFcf2x077HtXxM+f2IPfApV7wTuoCzo0SfJ7
9a3EN4uUwBq0r5LagVrpk/+nzUsP04Cj3U9Re8DFXAoEJtJ5TglsWB5P6wcaJBkPOAd82wfYuhaN
fJsoVh2dquRLNoIjwqOJ5VZwOMmSca9gNZMy/ykB3HDVBUlVGnmOKg/ZJu8fUpQkKTZwwe/3WeYR
bgB1h4KaZEE5CGOznzUooEyBVW7ligi5tu5Y1XLkTiVCYnPtcHsCSbtWe2KMprD6uQbD28yHpLq+
8MmmsKUOXutgLJLMvvOa8uBqMXPoYugmbmaMuJKdV9BjbrJocVi5tzkOLhrObq5zPb8xMYhaK9Hb
nuFZ9VTci6NYBQDQ1fGSY+bm8nrxh2hvs0FZdkbTPu1hqzZ1gQgTgt34jA2G/AA0Vcq3PJKKN3mi
c4hqcOlID4cxuDMbVjYldi0WT9hVdjqHwxn98H8thqUE2Uv1rKKZCqQYBpvu3c2MREAQFpmBcezs
FYHStNtr0DUuyHHdZemwkVOny9PYRvqAD7D3LYe6wrkEEmMBI39G8cGBl5+bsUwoDJ/VBEEKk5Wa
ztHGPrHP2CkgEecI1SqJ9bfvwLbPB/I5h2htRaoH78DyEGLJVE8enij8E0FhZXyX0Xr36TahtYlo
9kwVqSPkYpJln6oey8GlNaB+mr1a4OxBsJgvd/038LkCU3Fvt1nOHu+zcTWhET9GVo55ijZij8nz
o1oy7ZlztwidfL3FRR4HwDJ9tPoLslqX4wJuJFJu2F3Wzozd++M3+iFA46goDgVqcBtBoaEWuOJ+
JNxM1WXhLX1wCbmx2cHfyVhLrakWjoMY3lND4HRK0psTT4YgX8feVDoZ7zKLX6mSb+MidI3joFBZ
joI481rtGJvdmgnZBZH5zgff1EPtgaoiOSvWLnt9jzzzdHzV6NInJ2zOcT04tva866541zIsmByj
A3RbY8kbfn4woUCIcS4UCYGAuxBMGGwrzjB76EIHVWxHXl7X41SBBAg0+JmkqPD8bEpiNfFjmPJ9
q6Vkm8fCWfn8Cv7JzuTyr1l8YUCGAxBImGlzB7yDYLKgvrRJx/KQmR3HcYiZbOUJ0MFAhW5+GC0R
IQonYRvO5EHfrVSl7G8doASD/o9qa8SQjS3vKjClSFylMsGeKsjKdtFKatrVpvsLcNRIPkJqbGd5
TO9oTg6V4Mhn+iiELiPiYV1ud9pJUgMHrVZcSzye549PvnZeYAsF65RFtcOz1rzUMkKQwi0oYX95
a9V9YZ/75CqKQXKqh2asB/dwcYIA6IeavUVr3tA9M1YQNQV/c5Ztt6V6VMUHEUxX8iyiY/Z81C1I
GlSkrW15S/Ope1QJ6CPbpWzBr6xQKZDW/5AOTltzKbkT853riNP/+5O54upRn8vV/4h3hVRapzxl
kklA65oi9FGkBXUcgFBTnAso469NuKYIQWSUtLavNSsZ+vAgyrv5fHTIhaiuvc3hHgWuSOPnyq9l
JUqXjegLVgWEX+u9I8ikG1bzx7DcXMEKeU8BgUHOqZxPMM5WJqIjsU2jbtIlKqb4zOMhX9ASlW0A
LqQlw2qEvqcGMS2N7PL3OANAfyCsWkQEF095ee0ezuGCRXnejUg2cS5SmPgKUoS7GOWe6Km138J+
r91S9JOola6KIv+QaENWt4JmqJFUSMvVDmvmv+kf4K6imci77MXJoIJAyzqnbyJo0V+2QyyEdkPz
rbCURHk1Q9K6IsP/hNAF9MT0HCIVbOwEy8SnJtjd05ap0YhY9BOYv61H/mqEuK4k58XTvaV62tEx
iLG6PMW6bhGn+YS8TsLh9VbVO0gfFQmbWcNpfLt+e98p44mpSaFUxWXBGp7f8hiQ37xNBIZJvNcx
F9+mt5YgROooO8wG9wgLNDFt0Zdfe+r7Zfjl2vPF92Iw+jUj1p4UMHpYNtiQy0yj2/QiLwh3a/q3
DXLzDmmlEh/JdgV78l+i3ZqBhWwhfhXHWgJgS7mxjx33j8kzquBYyh5693ct77lghJzTfasuBtI4
C/SnVETDokk3IWJNzJGb5JtDAHEa9jCSdY7Q1VC1l21y0sne0j6b7ApAZ4jmlz9QWf3Fvq+rpQlf
1XditoqBYfkiNCG7scjNzbRHQx+9TVk/pFLG+tMbQAmL3rkso8PUTuQskuol8PI3dzHXM64pe0Si
ZJzq8XHha+StmwyERte77LGCro97bAxrHcnIxrtBa7GlHhovlCNOfdmgWRFOFxnIJJWsIF+bYuvo
ebggV9J/3PLC0R21Edb4KIgdrsD/GldR3u6fDY0+3gpypD/PsR/3bN/8YBht2TR7jZpdP8uTvr3s
8ORfCWW5UWHuS1lR/50WGK+MOz4LezEdry8EFJp17DZB5uWaZqob5O1s/LiMH3I+oJnVQZlZ4zMd
+dwu79dlNq0B091rmFH4EhtTxrMLkyEc2MOrP6l8KlSfHb3GkXD8ogE+Y6OUAR7cVa/wMftYDX0Q
Bpbyr68D3jK4mOT/8c2uHiTucG3yBfgd3zmw6TI0Qo4IEaWMIGpDNfBEeCckUG8zrY2kFdUBH5UD
AEG1Da7m5d2yiL6xJq9UuCQQYkSjBJR8auq/9tka9vaj2WN1MYHR4E5JqKclljZSlRNNWMhD3ldX
WfGBD6SdX7uTXI+YRKMb4dOno9oGRUOTykvNm5vzZ+nhJGbATKVdqotvCKDucHQJnQHuPetoc6WQ
CDhNJmet2DVSBnn3fFRMIRKfUSMFvO/+4xdEID3F8r67/FwHur7jVJ+SlxmFNmyIMn4hS4PBQhWK
EgXVr//AMo1r3R5v55guOAr/HLlXPsiojnNn47zl+gGDJ5L7MHmd9hatabZ+hFmYcwMtrb0ucMdu
lXNUtVRwjSrMmUAiiuelBPkokvd+T08nAa0rgnNYxH5s/yXB+cXiVT4R/OhXv0kp6NjCDJIitADe
q/8lqMEGGd6sJfkSN9t6mFyidCneK0glNoROzdsx2Tm1LxMytxYBPf8iRpymuORhCIJRHlK5GUKz
3wMJ67lSyyxg/nyZ8OMWPcNintXU6AJlo0p+cQ2vTPjrXTEMajF6r28mrkjJSh0Smi88ZGZC1RG0
wx22bLIwOvxvP2Ur7Bqrc1YUGm8U7dPpXxA0JbpQRpyxR1XHJFdoxjwoUNR3WRDnCmx7f1gW4pa1
NBuZz2rBbKY49oj3uPxCB3Scs9bFps79q11PjzUyFEB1Ffu+T7UPgBOjpSOU91yuxG+78ZwB/2Rx
5XpBOpzZP1ruKPUmh75sOMGKI1Q7xvxNv0+MbvKz/I0C5jgDiMUHPk/rnHF7AzYuZg7kau8o+gbH
yD6h4m8V64TvM+ZjdHUwsqsb3uDu62geEhfhChiNgFxa59iU+vVfU2QHxr8DrMdpBueZGfZQ9r3z
5H/IvQIQJxy2rAL+rwYV1zu7fMUtgAiVYTRQYcBsib/VunhpLeCHrA3bIcx+Djdzi4OGMhHfE9vI
pyO2vlfdLuvPW7lA6XGvjB9HFnsWGO2QBxIER+iZxrkqyuqWrBN04FPqXrL8FdnfecFavsIF5rKK
Lb5UG5cz2mPiZROHpwFb/isc9h6dnzwlE7nD/btmPVR3f/OMJ1d42ggoSjTay4QddDdpUY9b2xJ3
kjRYySgo7FyVBrq0DvM/a3adS0rRi1vQoXKzJcys0mC2lzocwGqiCI/45wtagTdky+dbuo8yEwZG
yj8aSgXl1BN10uvSLUI3DERdZ7L0g7/8w1WJ+Bc40OS5ljj8U7b8ACyB7vj4IKhBj7IybN00dvEa
jaN8XeRfYooiALw0xdwD7Yb4kqk5ZslvM0GM7WRDZj044DhWTX86XXpkGSxTFGkhDP5FGsHRWfMO
KP3RXWOR0C3dtvL0NPPA0WZGxgAw/jR+/hsY7gnGCAtASK0rrJ1o67wYkPqC4gygiiK6oVvrthZj
DfciUCVykhAF0Ni/MFK0DGQzad3QUALTaig99GE5xU9G99nHva1fYMtAGx82CJ6sxu41zneVKKej
ZnwMUdL/B6ebBbMKvHNk6VkKc1LBqMAf10l9jKKbnOw+EHJe7a9NvkNV82YpM4I+q1DWugFP1tdQ
X2HYb/YQ1KLCUvQn/F5xfJDzKddXWzXXZLDuJbncH/FlJ6lTbpJc0GZ+tFoPBBz0SNZXuix0REz1
6bx/K4c91ki4Ky+ZN/+swpH+YmPuM8ZZeXvKXNktsGjhixVKOQ2MXH2Ts4b0d6lDWek/BRbMwdKo
L/qWVF70m++a2AakRlB4u7WypZKEXPOevddbznzjHhk2Oir1q5a8MQEvOwVWTS3bDzjkRMzIShFc
8wl0vwKfI+hhGO4UbIXAe+jAjpsLKw8Hs8LdZ+UZZxDJqLfi+2wdomRj4JLzD6yoGSccJtDAEdFK
WKmuvDM4rj2fDoEMomdBUlpPR7YhEpdaFP0S6SKMIzc7HpHn0Ax6mB67rcRgAA0qwdk2fGldtwAx
2+Hd0Tik2j6lUWS5QhSLsi6vSDBE6PmKuVfVDni/2zWbua2aVHiiqJLZng70yjVPVf86Br9cx8BS
3I1ahTMi9uONfSmyhqanqWsrMLjai4qqLCxQ0b1Et4oqHbdh0az3C5xrnLSoZsKwUGojvKehoSdN
j6rJxqchJU5B7dqQ6i1k1PjoTOs9tK8FyYizcZ/OENRQnR0sBFJLIX9lT8Uk+EZZ4Tb3sy02eL3s
MQtKJbubOfN6BgJpdYazeNO1lnoeIPmptpDp82u+t+0dyQTLlJj19uRxM5S6imM5Q6UyKpVXGE5+
fubxhGM/Z9UxMAUUU/50mBHbNPp7ULGuhIDBvFYU4hIk2Jtea0nBIYVUH/drsg8PQF0RXraGS5sQ
6T5s4CJ+orMjF5OWauyZVU8IDbfiqy9zcVb9VEZ/i8Bsh5cgq5GA8BMaOSKL9wC2/YbAlkpcdlZf
1NV+JW6xytnHmKC1K2vj3nEjcSrgme8+ngoqqHkUCd1myip9RZWvjWA7V4TiUg8DDkVsBbAdKRxT
DUw+3hvxmQ3sva96v/mEHXWOqsvq02jpUQVqv5qeABIWcUmu07nxklbjeFcpuotXA8X/yVpOXO5D
Uxy9XLxUC9v74jOyTDN3DDQuuKtqfYtcJ13MBaYWJi+tgmnhxsjvP8knSsKN7H3kmXnC+ZMp563C
GLngQjmuRuezVL8jtHaRbBNlQ46jpqGDzQBBDlnOraFxjMEZwqYAxBeIyduVZDtcTQcymmk3W8Vx
zFzLZIS7SM0kPfaE5BXfK/LWgTHQEkFFc+caKsGW2DeFfNQxhCX083Q273zIAkxMn4JEIgZGJgtW
g024kjrLSJDHGEunLgfnemF4HGsxTVRAl0eLwwLCNKFUR8wGZc6VNzklIRy74tzf1CBpf4C3ZJ3z
O6QMHp+iyVV3s3prAiGPcB4fQxlRk7EcT4ycvNGOwqD094Md1R9laTonwjOIILbnNc4OO/Znb9Ps
C2errKY5ETZ/sMiukcdnFSAZMiay1qQoyCi3DOPOxurrUpQK1Cm9gxkYtAC8dFvCCubsv0Mey187
NIq4dqo+XnI16prQJvAEgPw1smt4zgm75R+NRqbG3IHzdSX+wZWJEKYoDltDOps3wx9encsOOGlE
bdGHslsF/H8K6IYWpfPzVH8pHW0ssilQ1LhqO6R6cmhdJPrl71rh3Ip0ZNSFpgOdrKWBNIa2ZC/N
EZjMNMwStIl65aePZXNxk+C+BJl1FgWUgu80S7Uz3kB99jiP6988R0YfZ/yUQP5zJuZZZ7wXQJoX
sOkZgRN2e1VF9QLOa2h2B17YpxNwzTm0LQtfCW6vh54Z+pu+ElO3bSQDzB+1vL25UzX3kg0LPkAD
1EYUydXrMXPasjnsFmwVkThSgdMTutMnvY94AQWxLhxjW8QW+p53qf7ZUlXi81BKHVwJuf7gHUes
bXsPbEWJAjuLVyutiIgX7fohpG0VFx/1ZnINxPoimlkn60uordEYm4d5iMOmg/wx+fL58poQ0f6V
DLQNemQaZAHZpha/+Ezr0ZrzrGM6pnZIscWM2ls9uIXDmyRZxg1DeY3T3s6ifwfNY6sDT2d6m501
mt1VEKb0EGTKY153Dbl9Ln+beGDcVOSVKgl8VHCdCSsDoQ2guKLZc+r+jxUPw4gPgHxBlTdA8zVn
JzZQgk2Zw56ClgVbrdZwIrCJV+7h8MzNQpafqVIwhA59C1eH3RIxrtUJz40O6ueKIIgZNSbqdkVe
aG5qkvVbIC8MrUGsrG6E94z085at0OF5Q80D0T6/ZUKn2Pwda6u56jpKIi+SRpRMcQlSDssvZwPw
CiGD2BCeeE3h0gsPNS+oV/p7YPOStnLuflemyM7bcccf3Sn85WaP1rJQ8yRXmoziC0e/6ytXHNbs
bc6MJKwRyAhrKccdzZvG5/z2+EewcQX3cf1n83ejc6zpLugVRHISZigg2h+TSFLZKXc0f+I+tDUW
xA8jQ7dZid2oh4pZXAky6uGZ2tE3yWf0k4s5duuOll5XzzkDIoSc7au3KhhvQaJypEgN5SNzM+oc
84eF8YD7jvdQDPFbN9e1iNLl+w+o5upyLc/1eg5IJRny2ZaFEaj18RIObPR4V+faPSmVgNsYhovz
NENn6L1FuJHhfIiDy1VXWsUKYSTihzzGOj9LC1Bj+Ha83JuSC8KKzkElobpytO4byzURHer6sIuX
wNutTlJUchz5FmXPxepBP9jZyYyrhivhvRJUq6vcpxKih2mk0gOBGPdtVH1E+mcazaFyeB3ACEzE
mmxerkl6yuk35sgtZaOqqLcYvIY8h+YMLySiol/6vrl9kZUEIWqWT1Qo7Eu7l121pFq5Nf4nTtBe
fbQYdkhdgKO5R6qibICzW9nyhcJF0L+wt9OPqFssdyX95a33KRU91d4T4vZETgUzv8buJV+BQHCv
AmDrkIJn+wxc3tNRslVa60Tm8NDmYZVNbo3CvEdUcjMQwAE3D8cOvfo29mE6xbJyfwna64Ejr+it
CuA27tbTPH3SykOxq/SL+rbVIG8LMVCHVatg9box4KdnVpOnQOhjlfKjK6J49BdO7e0P/ZmSvlaw
MCYqV9J1Qzr4qKiamZCFl5FiJnc6xmo4fN+KDacA0euNX6OKqw+odi/uREWlNzE/5LuDhVO02bM4
TGilWeTCtOm8r/5vUorWdQ5NL6DquY3feeX/x/77e3nMLK4XO0veYsdD3xZ+IQ1J5kZBlS7MgyJj
zwE7KEakofWw6p0ch7dbD2o4ACLAzhmjv21/KKArgg2Gps8dTMGITaWxEX6UWiDIKO9FRFHcs8sc
5hBBQVEK84IQXGvbpg1YZso+0qW8Kj8kPDdY+4ZqOb89w/4x0zXN1NE+skEGYaOIJjRjeD3b/+wK
qPgNXikim9K6Bza2Gid0VhJTCFk/hE71ozuuKqbrkE5EQZJ+pZgkd0JbgUpsC3EPulusuLj36P7m
SikCaFECfgDS8Z4GxpAgZZngxo1poOQhbi+xqyrN+sna7CFSRuES3BSHZK+yXr3zJrAZI66pFaH9
y8mRMka9Pu3YY+a+LYUhGULTHQ5I4OsJ2F8tWaeMrRljwhGystzunKPfV62F6s8PqMB8+IXInbNd
/hXTEqIvxFsqVhgz5YQXk5clk6pbeCQU/QpgccN76+VjP0Vi4gqMLg7qYaBdU4PxpbK0LarlAXPU
vNrNrd6wDNMLqMDRZDDoHqpqSp7xXD76ZP5nYSvX4EVQx8C2R0JwcWm0yF7uYKFPG6F/BVGbvUy+
DqMBNNyiC1gs+R2jmUWQv8skgrunzp2luSYoC0QZOw+L/CYw9fyy9kULU0zsu8eSt6mVgcDuZmLV
VuVWmulP07jmMaP8h+y7HaGaHlkWoLEhCB3RjBzP8NQEzH1QBQYBONALLUYZBcZHlbEa7KpdFjff
3x4LctaAmiNBdokuZfrybJ0hVBzCpOWqNAL+5ICnx65H6qCIK6rt/nLkGlJk6tOzfFPlpRqmMmV+
gWAEDDtNf3mUnZjwSXUQJ8sScH3IKSY7jizBjQQnr9rggakckzI5YhdN8hiCPcGWnSO4JWMebVPs
b3RH/MVBojcg3y9enz8o92qKWsXOsUZ/bFq73fw5RkB6hemna6x1jm5VxTmY8uM7p5MzkCchNMhx
iz0g2s/VQUzgtKiKVh/d8EsnI4vjNBkE/4DNTGolYSDueb8fMdNuYrfKgiBzhTs8AK1g2UMhJLGa
+UmtHl2ExWGgPn2lUWcl46FVO70SazB1jY5JDfCdnRntSqVBZTfsgGq1AJtSrvletD1YnIakalXy
+77O9D2ajlKeGcbHtmPZqCACRJz+xuggyW4BVIqUIuKskhAwTZW7rraRMt9BrrSjRvfMk7iRnFLo
TnVid4S8LXO25efrmL8Vlj8UXeXET0sZOe7ntYULfHo2C+Pg3PwW6tc4LXCY8iVttztK2Mk73yv+
dIbyZuGnn9d+OplRdKIbKokfq8HVsJFsdIHWp4DE1eWB9nOT6r8kAzlsJ8oIaxu0rBrXvMf2slaM
PHdODRfB/EDDSI8BRAer7yvKSt2iZIz691dZdQYDyxt+Ojbym0mg8SPV6qbkH+4NwX+5rmH4nC8Y
aeo64ArcEOO1f7NVqg8d8iacV+7b0dwBp+LlFO+SlFPalxf/FP/0nxYexN9q6JfgnY9UXxD0WVfD
WUjUjnMRIndsuWnYfF4xmXN89XvzJBxisRAqZFRtcpCFaRKZ+I59cV+LuVukAM8e2yjWBEYbx5lg
3Ci5LbDeEJDMI1SL36oyos1q2H/pIefuOmH5cCMSFyBbQ/vcnDpvE+q3GS5OaMNL7M+Oh+/cIVi0
iq5pHBQ5sN9RdYc5wHz1olfp7Hxh3dP4mlH60JzYauBvBGLNMyDF5DS+6JZ/XlSAylwIqLX49+GP
SGbzQnJL/KKIU5PYrmv9SKkeOtwVebIEiQsobzzYeUsKfFRJ3x2GjdEthjuofXGcWqZKmqNVrctq
Q7IlqG+wS/LPwBB70KlKTRt3H46/ShB3yfnxvh8KubE84FtmEO6lic6T/235QeTG0gqcVw4bn3UE
HhOJn5N1ePnjEhMPAPfo79vShuxILhuTT5uA+rOsRcrBNa5CHqeN/GhZ5Z1R04p2I9Jk6F8ot+8s
vxTOARwb0MaztZ00pvqd6MI9WfMSZR2IKLRmSSHHj6FjJIPEGLrKpWJ7+8IiSDXcjdKNQsIsA2/j
pA55cMY9u9uZhiDAPsp/cXz+iLIRJg0Bpv947QM1IZuAat95arEPvSvM3raQcNtzcxwmFGT5Oota
PJ+sRz9hcMVtKHllFUG4e0LxGl5rZMqThCDjhxmm5/lfspuvDCZwssBZ9g7TlESTt9bdrdrwg7gR
aXc241X31Bf9pf+n4TTNg87dgfye6gt4EqJEeN3mGTniMw18QvV74GhiVhBL3wecCe5vJ1YoP8Mq
B3hH95YAt3ISdp3QqvSp2PdS78ckHX+M62rM0xYYivH+7sSCaDHFCF6zuXWz4O8IhN/VrCKp+KYO
x51ncmVrsDhZOaWMlIm+SiPyNwWjMhj/pqIcOSzswsyrorYRwpEaELLDYuwOqBkIyBhTrY4KiMNW
r/xgoKvblqbzJUgwMpnXMT/LZeIvJK7+XXCAqUuOGCrDH/1A1QvZDo7l2c17XCBiUbQsrwSs2lIw
DWxaSagk5dePKPM8To6oD9EjbfwBjbab5Fb+zbIWBkTfSuRzuFLqBeH4bffkddyXY9Fl6f6nnZKG
72rnUjCHxwPkmzHk3of4JbmcAl7ndURw2q6QSs/ltlhXuJO52X/6cWkE6t9InH3rxBA/gDLkf+Bh
x0rkxBhuze7q4TYuh14gJxLs4OjpY0zH2a5YoZzR2cXG3+Gu5GQpYapMeWtRYpzsutklwlj5yVsy
gByZ/2IX9/6IuI0Xt76ej414omF2SBu7KG1xd/8TtgQYDOhi0GHGFKvh4nVundeCZlhtU7KCCXt/
9GdMY+Wt+4geTuLYHytjTAtx082sLmsIAssFAOwlxRGWlf/KdQ7oxOQN/5q25/dqQOYnNkfMNOd8
L5onvFdVHdK3wdpr6vLRrtJxDMtTt2oBOZTczJdjVe6wA3iaQKlw5SC+45eFxWHmFJxc0xFeYAba
iNLtn8c5lkHVkR6IQXxrQy15Hlcc7cOZpbZYQyR723lQqlPMiSTHwsvzZSOjewOb8C4pEA4ioZke
pK3pJqVE8qYjF7npCpAN8Uygs12PGT1vfDBMN5dzJq/FI57h+ebDAtQg6ANo8z7sPfX6RvwjOBZh
2J87Mxd1wLe3I01EoKbFdAqcNQ5E0+bOh6dnFutOql1MtQsRPTPKrkIr35jZOMLisIe4Rpps6Gf/
p24rcDHH11NTHDiwN4HqQA3xztwUBd48HINReoAR6B95Hu37KWtPIJPChhHhcB9K3Eluiscma8H1
Zc48Brd61YEKVWWTkh13bRb1ymiMrGY4vqWOBmfXjDXN7o1Z4jhDmwxNEfI71AfYuFjkMqZgxSi4
yDBDSLCXUILFyna0jG9BZDMMxynFgiBNbMw2xD5dx/WmDMr0CbtDDi6j9kkrpsZQFnxCTT7xIFAe
YOcreU1Vja15pmdO8Gr6DzJVjrTqr++CWNm2PY170yxFZptmcWB2naoaOioG5pXy16i0Sddc1clW
w48T7bzdvMPSakS5VQ61x7yZJJoRXX4Wec4WB4inJM69+0kxwW/o9LWdJtqI1+2lVLokB1KlFqdF
kAuuHTIsQDumHSV5SPzkKt5vrXDGceHylKeCIhcdwINd6ovSQcscWSEQYRaM7rRUORoURRruIgfd
4RUBburDFFu9BbDqj66To3rNuz5BWbZu9j9Y50Ikm6hB5Qj5ZAL4QRAuhDewGYOR3txWb7PuXXZM
oiE6MLb96AkguWPSVsc44WwmBLMN5bp0At2BYHTOY1RRmuleCcZTLgZssZBsTVQdrgv/dXjGd/sb
iTkRh1y6DiR3auorMf8bqaJQ58sci5zONrQmhBBpRfP35qMPvrGCufBS60CcTPn83N1o8Vu/KdVK
sHWT++UMNcqzeRRIWgdf6Xy1GYmZ/wzNa2vsLjf//OtpMq1gOAk/QbfoY/8lxGH7Ou9D4maWaRzt
39i8dpDwhZ5jIVWoNNEjEZ2phD3DyO2EAVYRvUCA0+xpW56jCmg8gr5DXP1BUQHp2VdftnhGOTul
TzJMM78ToQ0e65VyYqxvMdrN+f8EvoifaREZGfby9tQYpDH3qfiTqsvDCFXSbe3kwxS7zLuJvcAC
x8uexKig1+1R9qhyMAjrZq1hwhQj+bkTf86nmY8vbFzzRZi0oianTEGgUMealCx5ZL7ZGZCErSuN
w2amTaBmJowA/77gqCbehSPhyoQNhjw3SGc1JCWyypv28f7WrmwDuAYqlE8A3XvNZOLVXctRW9Tr
kaxu1LhDFBNrORlhizcHEiRz1bLR8vqSE5T3aSXSDzfh4vKwgDj4lcwqF/qxAE3YowYJs8Ar4WRR
IPThZwdYLjxndGReNH3pk1y+2n9U0OmdHyQHHmka1OeYfWh75AcHNbX63oXPKSz1P1NVWLx1AhzG
5Gk9qvRp0FlJqgzrvc1lzS0bQTAjkvkWBpu2dRNNcppEHUzJZMas6OwXwSNxgC08GHGd/cMkNQOA
hc9rhsKW+OfESjFLcX2f6nOxxcpkmHDZlWDTJWprd8wYmKTnyokI741NykUD6mH16Cp2URh1BiAp
+tjKyZkvq5Brrdh9UyljpVGdOr0r3eq/SzhIaQ6khbLmcXQW/a6tcPVRADm2LriuG2/Stkcj8tkT
QlxEMaxxH7XJGvUrVTZOMO6iG9FQH8043bhg6fYMRkMiHUhGyZTq2SxrmpVNWf5HCGdd14FsDDU7
SCmNx80ykZAL+LEmHrmtUvWQbf1WFxzpsNw19QWb7QsJwpmT+dY5gMGu2Aj1yYP1bzeN3kvYk+bp
qW7bDklW/zpjLBU4sYZkJ4+ZX2C7FuO3FHEwA3+OwbXAp1cZe/PbXocsUMxaiILMnN6AyAEaQFV4
19s/eAZmPSjg9d2RgFOdbENlSpPEPVrMYJRXlFpAHd4FeA3J2TeFNfzs7wMbFrjGExCujFXrpQ+Q
bhh91C0hvTdJM9Ei1mqpxHEQz5xvEAdEsHz3MBKX0AerXoXVhG0XL2vx1Noiq1a7kmnGkY+N1asM
LduZpQgrErDj5JI/KzZvy7zqFPhFpJCbjlTFrMVtCfiGX3huXdqc9cqmyB4jgXoWRUiZn8y47L2K
wW43OYvxDjnQjzwC3Zn9TYD9Bb5Yo/LGDdt3amlw9UiwFxD0in0kL0SMEt3BCk1N+kPYBcHkckbz
slhcULwrmoIfkiTQrsKcFLq15VPRWM6TaZSg/0JGwa5c6tn0Y61jAq9qTREinSoUPBfgf/WZnl01
Hnsj+VYEmJzjpSd+QhG052Lha5AJ2SJErFbRZbvenGOzfk/irU46xOSzrDwjovP/USyM7vyRDw/q
YWUCCMTkoRHnwwIvzeZkoKgo5Vr2XF0rhhZHXuOX+SqaoImaFELNqDkVLo3PFQC9V7L2oKZnEswy
0x+k8Ccgrp9fwfODkd4+KcwdFLKuS2wf5WC/m4Wa4Ce3PInT2OueFlsykcDbsifUa+duoUexcik2
N733jV9y8gtpNdsDXjrfaJp+LUEghxHjp2f6VczAnwiNu6dt4eu8mnVmKkYOjzFiyUl2HU8oitVe
MDtctc6nsDjizaj8J2BpNB5O/4+vqEqOqsnBXEbkZEIcGrCBfMuJ3dH7UnON/S8112wdheNqITVa
4M/Pn6xqLIc/TMzByZ889IA12sFx0NgbWaVvrfQd4kkRVGCYYP2OtqXPswaMw8OCRpJa7Dn+YRrD
e8LyBIVQB/+QYPFI9+AzUPBPskpsi2CaIK23NHFJb65r36e12PjDdPMwEJUHM7IJb9IcOUiL8LIx
MJuC9OfUY4yuN34UuWdnboUQ+DLizAnua+JkDMr834vTM7Jwqo+4pCbkm8guQ5wyIyvMHT14JsSm
E87kLOOzsV1wk0jBllJ1pBxw/YJXwJpgUD9IuhClefMMJQvhrIYs9W/sMU1VWH9TSOIBTK2sP6Yi
cROTxg8at057jY7EfgNSL0+qAF+kAvQFEooPuIiRC+edBC6TYLPVAoYeWHinmTgrDOMKh0ZLfOKY
/FFgfW8llCRNujkLoxcaQoZejY42kUNegn7RvxP7qZ1GQIHO1wMDDElQfHOvnWOkJuUHzP0kklhB
/LfQ6JD1Rm9wGDMhXa3nAlItZOwWIHGqMvAttY28EL+qWG62bjIRaUFfI+ttwSHsIMSykl7iidcK
1xm0I5SekdzdwK0KqB0z7lBY1TaIBIAvfIPbPZi6as3yh0v/zQNSbI876iodh1nkFlX1Su5nV/2l
HvrGPBI4QFAXu2Oo+P53OFsY7aaz2TQocpPFe3NT3l/351NUWnf9E5tVCmR2kB5EaqpkrDdLRZuQ
HlEGIyonkZRJkW5vPXOJfe9k99sPT5GAErPTmjexnCfjtcMzVk6KBgK+v3ZUGVuc1CNLvKP/rW4B
uaMNYVBrU4G0mFk8bMbzSC5mF/Y3LMeZAjjz9iMS/6VqmrHyYsMsGwQMiZgwKCSQgA/MHrdd3o2n
WimuhD2HqtSCV6LRExMfiQCLaEBb8HnKu4GFIhJARCN428iMoIVFfG4qHUENltMdn9oPjMxSq8cF
uiLrFySuT7/4i9xJ74yUcYV9Eq+7M9in8WlrllXMBxMaNP4oKk8tUgBQWPpA866DoAX6PF8MsLDM
TAaViWGo3JQyticXrhQe/qkUKTSzfy/mzYI0rSlYq0kK+jMTyWH2NiDS1DkhPosegMPRFCilOWla
ERe4ddPzgNhkvgNbWaAxL2QIP4KYK+AjXuUQpBYwJt7/MA9D+g1vtHGqYRngJw5pwevsNWJ/KrbU
C8rmYYfIQvj34p+aKGqCIgS9qcghkz4FKcrAttE6xq4CLCcqlBfMjxIROslXDIFquh/9QXQ6mzDh
LkdalohlzNVkoTx4oAQbnYWleYpCPZv+FP/R+cERSq0VVnjZtr94xhpCYQNcw9gKaw0RWHtumDmL
iZwms0fI9IH3dst3Le5AoPMXrUuWJznZgyAiH29bHR5MZfzRNeldxDBu7tL3lKuObPLRkM/ny9Wj
bb+CJshmgHKFXK6040XI1n9ssJVYH+rOTCEvLqhOuodET6IEHtQEB9NgiqZOSM3Or3YwlxyR2mDC
7cXewrdbwUCke8QNoCCTXno7vIusMU7mrgdRPOZAlrlv/W+S+J1yvFPD4RYOIOH6ZcimZ9TwjxFd
V3MkXUXql+v1iTSWv5Ji90hLW3kNGtVgPjywbLyqB/omaK9OFbbuJAi7oyfl6Bw2fdOo8gz3PedL
o6VUI37UT1UxkF6NbP0/IltBVxAgRIJqXHRp+XlZOFH4DP5AP1OUkeE1zEaymqFD2H2v2oUJD5uZ
wZTACjwA2deC8dyH/gLKgmh8Py7lYBLVKXVRsOalOzO2aL6LR5cvvuI5g9G3aGDY/yLFFlDMFuGW
cRDgV6Uz9oUd9/e2ut/0Y2ERhhwI1oXtlNiBxBwk608UJETIaffTB4fucOgNWhWlNNspBpW7Fcyc
3Ob4V0KTU1hb3KJb/y8BIWYP1Nr55hHGe7YlcpMBI1BDE4B5op0oO1VDkPeslJghi5tdD/ju/3jD
aknGWl7XxXALvyuUdNwYPecA23s/pjG34hP5gwpcVaScwz5W7bk8iho0jPYHsDKq2rEADApzPRSf
3FISray99X3M7ACfSFXLWQaHQxC9btuP9/1BB9E6rPQhgP4ULyoHBBEvrl26cuLNewRn1i+ByOZS
cemqeSgZXo5edIKaEktWb/Y2q/EuKmjCC5VcaOgSdBMTx7fU1mmpZhV4ZRZYt/3w2x4tB1hO2Gva
riaqhOenbyIjRaWvv79VHf1L/3oEAl62WbbrA6WX45rAL0cmt5CpjusMfsDnW/PWo6HPd2Fhi/TT
aNummBUblKi52HQL8VZuOfJXxt1hwVeu/6S1nXkRTzzFNFWeXwF3twM0iEXfFMJcwJ09SNxpTdvV
CbhY7jVWz5PZ99anxCOgx4xaxPb2a/kS6N9Xoh0GyNdWLyWT1EOx5wffE/whWTial5RaUZTQVJKi
TiKla9yn7fS/KQIDG0dJjaYSQ3IHoccnWe21bONaahAsk4TJfTH9BB8YnF58j8EeAUqzC3mLq/q0
mr4FjE2gMjNAuxmTliH2NhTAzdpEZQ6fBvrw/2h2Nv8e3EnQ6liQcGc+XxpRNrhZHPiMsxY9C5bI
zPcoCTOAmFbNG5tQlwH1qguQq8VWsz7myPtqErwgPL0DnYjTcgs0oznlcfvTSwdaHUaUB4jrDnDP
5q2HCUzMH6sPCz5zINj14X/ifBoKap+488+NWVMJ9s3fkNv4SOQKn3OwBE91nMtE0H5lqQaUpiBh
hyeUB00VIpJ8cpEgtOPqBK936cVT/DshEfSpPoy1jf6AjsaX9+AhVvY+XjcTrFxAlJ/6mo9zpA/c
ZzzLrqlAkxEbjWl06/tQtu3yUFyrJGayoWZgTvJJfNBPTJuHQm6FTsjCqCY4w7BfgxW7kCwmkWMV
/QPVl+iK460H0QwQyCuNR82Me2jrjWD9ufSDtuhdJzx9Ebf+y6diVQCUWDjVinxxBKRqRCiISTJt
jmVVHMXMsyhOsPeX0fFiOjulz3I0i2yYwX5e3qMj3BkEGuf9MYhynHWuTJNYI/iCZeFQuVXh7rAS
d+AsEQSnVYMks/jTDYKksr0Bp4Xw3uNTBTVAIEWpbg9yYqImLfULIe6nTjHaH4jJ789sXhWcUa7A
dywzHN/tCWcT8AsV5sfQW8FmA3s8QdUBBySRrx6mGf3O2g2QNPqrQ5vUU68mIyOy32E2TTIqd9Cw
YU963rSiVeH+RMym7GLLVSzk9knzHBneyAthnAbfbtNg+iF6+BpLNFlmw7RRin8EuFu7kiwUY3qc
9mMWzRfHuJ3aaTvq29tDu2v5b8c262ja6W3hnQXL6nfjyLiEk7j9VSPuAzvgrAi08bnYU6FPwlah
DkGls0yBqEkH6oLIQRCjL3vcTOJwO3QFcdYMn3bWZq54Cd1jlT2tpT+4b6Uzgqc3NZVhjVkCS2Wr
Lhex40U7SJ6tip83nrY2z8s8kRFT4gOlNA9DbIZlllBe2MmxhyjO6WOFkIl3XqLxpBTbZ6khY9Hc
+DMynrr7sc+QGROH6dDPLoD20oHRlyiKUSpJ0/4+GxAjeBrJt2icM6tWoWN7nHdKoJjwrz+UIoBT
PuZKWz6SecJteCPwoJukktPucjsrosnYJvIaclByuo/ZfyWX4+0nYHgnJ8rP3DfFSByYsfbotd2Z
LnyNxKnpZLzcobze+zlYpgkHdewXwhMUvf2JsdMpvXb12U5KulE7OXbcAD00yRfNE+BnfKvd3/Vi
zIdXmmtjIC9EBgZI3xFQ+I657UO4LyeECSNzXxWEqYLgZCk6GEPwq3NSCrg2alNM4hiWbjoDUoCP
7cHdRQMLxJUbnS/t8lVif8D8LRunGFrc4lelo4vVcXQ/p4ttnGF7MUzJjj4+0wwll+pIIc6yboNI
yK28EAccdUykmbqabY4gUMoU44fSkqd9U0zNnRNcvAikESOov1gRESyAiS+iVfSX5W7QsDaJq01K
PaSzD/hpIf4EWhSWDWtAopMTqod+YqvxLti2PansSK1ebuALiyWGa0lGDayb5uGw4tD760hgjdvD
lAMSBGD6w0zODy/s7cRI+VTRzHeR4Txx4gbQN1SaJOo4LiG5s4mxWrC4oznys4s1GM/F6ZJaYjPU
Ej26yswVKx4zaB2LtAVMOgelhOimTAzDjoiv6jilCRw240f5pr/rBq0+TMRgoYjCHA6z40wbQzhM
zSykm6UDlT5tv4ogBYDvQ8yDVG5YfbXVklQwsZHKOjpQ31rcgDdzfa7zgYbCFFGWWjblo1oPi9io
IVS/BG2mPFxzPzkCJbKv456wYwCQ8MB83uOAfc8wLBhppUP3k+m7EXlsqSZRffk9MaN1ZyRb4v5L
RcFPnajrq0wEkyLt33ncpI4V1f4tueqt0uW2mhWMXL/x68Ul6kizVRoJUxQn7sXwe2AWa9jL+1R1
OBxAWLSytyWqnG+CrfOSBJZGXT1ywO6/mYVRPPk5IvPb+PJnzkruMHL67eYjvA8s5q/U9j26iSkc
nOcreZ09KtybqZSW7WbQmMkcZPAZwvDQlC/DGcUfA8NRJOug32paM4iheyS397/qX2ulg6/2sUeM
sN8IjRYkg9pk5eK0aUFoV3hhtop9s1pxg93xEN2JDWayUNAf/iatU0A1tFrV0poGtpZti4Za6IEL
Bgf4c3P6T3CWhr3lhYWNaYcbQXczZHfZiesjHxtMG2f2aW5vbfKYCcrOTKtoY2j8cP+i1CMa02Xd
GXwYbRC7qME7dBAEx2rr2QghzlK2xgsJCu5khPJBR122MjS/n7dNYbaChdnLTHt2OsXmivLwnX+s
kK05Z2jSRj2QMqPTUGbLCXRW3hryxi5/SZqWvTyC0sohf8GoYQjlLDOGYCIKdkOQNYMYy1wQ9Gqx
AfOwkt21H4F/qUHPSQWabd+MScexEQYNKVOgDUXcCCv2w9v2yfov/E3G5o+9gV5wraIPZm6p2xVF
cwEWgprS7E58dZKG6g8D0pfYviwwdd0BayJ1aGtmEPo4AFrA3Eikc8l4A6e28AN+yJWN9aiJJcFb
UPaLcKpb3AjMD9kRSvSPxBaBY36tBzpk2qx3XRSeo78Y7Zi1KR8sCwb2AXfFdCWDANWGtmsjbMzJ
dw2hzx0bxGTe6NnyJ3mNy0Wyb5d8eptvwv9N7wZVLaQ6deJWgLWO8mhDudWCgyjVQOQOBTWo1sbr
/ZcUxXA/oWjqxK65LvTqN8xzjc9NjGE8fwlJhfFU+YOupT7yXGN+tH0AzrDQb4MsfdM+ryCaZzNk
Kl2DixdMwGpthoNGsryFlJ/indm++lxSJCluDkGju8S3wkf0HYGMqarp3Tntz3x7VVxynrf+D0KJ
4lbYD0leigwE5gDIXlhiExksf+rQ2Z9+ZW5/EMQKtumObRDnd0mRYRRy59O4jiaP6jMBD8P8LWV0
bIzBLcsVccHLNB6Pd6RRnuLuke4Joco5CVGL3Yiis6Lhl5eyKHuuU5v4LfiuQczCE8TGIVm3bdKQ
AWC1jRycUQO21HIk9Onqei+DgewfA6iV/zFkopL5y6tmFDxatjHG02Svp71anWJoLUwraAfOqYdP
EXHx73cdnZlXvaduxFsFLavZ78zTcmGQd0bLjpnr77TQcy+NqG9h0mctHoH9eGwotdcngdX2nDNp
jUYDgm7QlDxOqgJq3hucbBnO7OKU4zcYEYa72Hvx3RUY6AsgHc1BVPklXr4d403SnMueDJXGqI+p
fcRZFNDHeWOABbrRBmAcy4D2zPLfZ9ddJ5u7tQc+EGYWQ4xUb86m1gREpiEYG5nZ4QvKiXXDNfWU
rxgBiPxh3BjiQ3+sTMASCYEQpbxbv2IOpWj685Vh8RSZF83EWPSVZqON8RaR8KdLY9dqn0n0LIm7
6tifpOm7O7FNqlTUoVi3yZAA5h7xACIyqErxLn6IBWlK554x0UDgvWBjnMuqgn3vhMBPjwZc2Ppg
rbFBnq6C7tAVWEHGS70CFhLE4JhWJOjs6W+qSENPyc3PNDiWaASFps0w8JwIM8dR0mlPT0SvcclW
XSAO4ysrXqnQhYPXgLTVaLONfuTKydo82MwLoe4w/fklQDmNNuS70ErtEYnkKtTdTvOPZ2PzAxgS
n+7t3HhvbQki5rewkQ269VUAH1QaIoOxfTuFdmkeDgJ8GoSyFsnEoTxz5gMhfgvk5qk8fETqufKL
ictJMePs8pM3w1fp6k60m9NiuJ0Zd32QsTlgF72JjDX0/ginAv86tzis1GhpISWPWPB9fCeHUe89
5hoOF9XCJjODFKjmr7WjxXcUYrQIUCfyp/BXnIz0NER8YKwEUPawh2SeX0VVdHvIrPXt2LO4BsO4
oJeNLlu4ptHiolEEVWt36PQTw7/4FQAJjIE4Yixt2FqvfQ1hmo1xxXcOj0aji6/jHWK9tn2UV8hD
TlIXI95ryCAcFJ+JByM37ddc9O4Ste/b8xAh4ZyxxeuSrK4pXn/p+hTjgpQbBn9aemUbOFDn6Qlt
x4pnOYHgKi9UCQe4n/vvoGbi2tMJAAQX1wkT/xvvwDdMRAejJht8Z1lD5/o9zvvFw7CUk+aObwbV
vGPNQRAPy6AYEfxZcojCLkjvhql+Qm/OG/sp5BVPWMj9vhDgC7TT/W1MSKLZBWVmBGqhAf9Anv/k
F+X3fv2zuhFlNXmPFnrAnrMPBYSC2v2X5VW1eSTDBcVa5BMSiNKlSOmwoXb5+gAf+pQOm+qu3qaD
mS80Xc1ikZoixj/I1VkkAoc6oq5cCwxhT28fDbeVmEQj8Mzome0DW+Vlq4bRodrea7Ibwjxrk4Tr
v+kLAupoAoUjDW8JSwrpZLZUC9mLX8yY/1A2iO8yUrfDitiBiVa9nu1WlT+SrhaxCwrdKjvAENXS
Z4T2y1Q6/o7pYeQ260f8SGsUs37XZZwOJ2nSHE+ug+lZ18h4xVBMdcuVKgFn7i1O2prBHKKjS9wv
wvVU3oC9UC16Vn7jOL4svzFjesN9rmJo9LPUBS8fQKBrBAHOIgzpaGZB+3xB49yAQxqHmV4TKd62
Dc0yDxxmOJ8R+ZWHMSykAcXK8KTNshFZ1zFci0nBBRngQZw9LWP5SHdiSH807VC1lL/zlaJa+FaS
VU51NWNdIUr4+YgCv5fnJ1py5jczLIcX+YLNr+tNK7MoeOnrsqMit37xOQ4kTZth+MK3ojYz2AhL
M7hfVoc+/ioAwsVaoHYCFxrDXQ2Z5BhDBIXTtYxOLpfouu8NUPwG9C55uBtzJyFhqpahda/4LbWZ
FtZr18Xm/5OjtmIpAAOhIZLIAlkrh88OgUPHhC2vWeEtfJPJ0h6HkxH7+gTUfdqFGt6cVcRW5/cF
QZVu9ncr/78KVdiqCVzT9PljMQM7rRxCVWEcANllDAVx1w7QfwhCsLOT7ADpEj7vHOnkOjwr9FW/
31nQSSf2nhbaeTjR+lsOAVFFghdcJRWtFWbcT2Vb7B2MnucVEuv+ntVrNDa7t9IRjpBc7CyyztfU
Y3xh5FpxKGCRwt8bqttpJG0exkrTVArmUFt7mR01nh+RcDa9aOJ65Dwy75S4JTooOVeS/U6P8j2Y
2MrnmcI+MLWfq63iq3UfutagQejz1Cn8PIUFJdIaB+0fQFnSXAAhBTyYt1WIoQNgkMh3TfnxQMmN
af09mtjCxa4XscDghGU5SNFy2abVtH42ya0dnSng7ACSWQedjIlxPmPjbBCB2Hc/mXrCSOtAc1vH
ABQsqMDE11GIodZDXPAfLT1YhcWk1anmnLIMb9fUB3/LC51Jh8kXYgCVj9XTd4Lbdu9Mxtszho9T
x9W4FOh0ITBYvjO3kuSSs6g+tC3s3BCUPUGn8FDpaBQiKfk/8X+McsccfIKp8Rk2ZFkOVYsf0cJA
qrSL3v9U9h7mdwUSM5HXkvseTJL6g8Bzr4x4rwmPfM4Mc9jVqas8yf8C5zpwQ57WqrPPWhFNgGKp
ywC9aD+ykRN5/PwR1g7fBu7SP41xFAxi/jUHSw6dl/XKjyXzJjyrF+E8TE/hNq2Uo6mMs7rW77or
5rFG5shGM6kLvYzvyU/px7figURgCfO79xqo1+ZSiV0lhOy9oGQkAdbPnKbuVJI1I8f5RCWErMI7
q3sLly/KxBwSZGPRB0lX5z8nI9YEHzObp/qLOMKbZ2UlbejJ1RAjMJGTFgMNaovVUr2JHUXUZUsf
5kya4TW8sLf8ahiLruM0zFEs+sZZyFJ/9MmeyVSKh+HKwF0woZVXVZzy4UsXpgg4gdiilecDvY/5
yFj0JJstAi5kfbOBG5oSMlj6g4Xla7+8IJWWn1Hj94hEXU3+5hz8kIUA1TCm5fMWiubveADTUyMe
DWQYIxUXL4hwtFjePwpU/jS3dzYje0SX6GZEThcM1zrgF9gPBh0DxsNMVJw5bt3NVkufjHysOBIA
mvOmedsdmFOJ9C7HqqKNmxzRww7EsCIroH2UqPXJgdDkc6lwUyIj62mTtjAmqfbcczjr9yq0cyrL
QrT3DdsCphMjTjWSCvN2yEpbe3k69JXqSy7wAGqEl8vt5d5yNwd1cdbzGmszGf0uFVye5PDo0r3k
0RnaKLXDuBxeAS8/CYT8Vo1nPg3Mwfd6wLUeEu7G6P7cKLM2lS2n3F6t/eF+ascEsutNr7UpqjgY
kxR7zBUs7aNLYYZ33omcLtRuPJpwU+ol4o4+qIoqRJZcDqHsLi72t5l6s8TkVIdjaEfSDp3Gwm6Y
ywobRa+WqlWt4Sixa05iyyR08bLsU+F1Ve5W+fLW/O+pte98dvnG7bfc1TRqrRmfTQ9O9k9C0P+R
+9nRKbcssKGNRbchJXl1dq1DKH73dXSywmvuDQIf9S1dfsUO/U25H5GYWA/t0v9hUA5HMSYHxL/8
8OMggnRfSdj3LDO9qU6mP7JNWrcpt6myVOvo/jfATw9Da5ubXUqNXn12aRRqy1S47JtZ5E0wmInm
bc8nWOokDESH61uBltw8VY6BLVPtRLxBlmuXdhXvJgP6HYrJEZpyp0l7MmRZZDSkGICoBxf/beGE
//CXmbf2Nw9CJjPxJtZAqKjtnAJAIaoFBTcSW+18lIojmWYjTgfjpvibVoqu5d5QbfzC8dKhJtit
LTHs8A3Scgy8Bkfw9jfw/hmQ3yHPa1aT4vhyzpNE++g732B/UQOTumC0NKCbihX9ZkHhhnTaPQmp
jbJAWy5ueydmV23oWZJgL1xUuVnB8obYfofCTAk2/DHoM8v3YZp7d+vKGlrAVCawOPXxsFQ5B3Q/
Wmg//foGGcTa9SBNzEr8gnRBH9N1jPzF+l5iM3m8UCqgAfvYyLwT7SODVjYmFN/Wz00vzIl8tVle
bqkZnsWyTdm+duWDoPTuMua0kJvKh7hennVwYirCUIE5LzuWqn/3gGqPwLagP0RR8pOjiSU4i163
P8zqQ5NWuAlh/LQ/nql5DKbHtoler0xTxYR9Itwgj1QV9qUB9EIXux/dzc7/EvI4dJUHcIqmWKWk
eg2jqX92Lhwfd0fJSw8cJkEphts0h4eKynnNGhEZSF50N/edwFduTRrsmMvHfzr1VEmqur02fxF4
xum43P3BBNGN5f3eshK423UEuNZ8Hs1CuI92lUpOTDFb11/1GGOwDuOgJl4daTgRKMgNyB+yDi/H
Ee4oHwtuhftMVVLCp4r3DE2vPcQwE/B9CEUiAiLWt/U6xYYF5eR491Ut7waChBoq956smQJ5Aw4c
hweB3se5PV6Bs2V+dtPOQ918iav4AzEbhHUSDb72nIP0mjrKpnAxeAUHsC6ldVWcND/sB0Awc8dW
YL8VHsm+L+sXckIsoam6iRqLViJF57kzMKKNcX9WDULqEPcTFbmdL5EY0a84n4ZS/jJy8LCtczWr
l0HOA9WastU3LSTJlvCZNGzfiVgFKhoQ90wtdMegK8PtT9a4xk/cUiZzseFp03Ka4OVOqPDZNVU1
MraGYvJZf0S56ZUHVbdCOERU/Go++xxnkhbJIqdRWCmFnMNmFUHOxxtqTXe3qORjBdVx4HfA3r3q
G7lV/ORrUnO4WbZpTzCjnpfjRlvyyXDsOuKWXAZjQp0wVTICuAf4GjfmGLMc9dT6012xvk3o/VeC
lCWJTmjc5n6ck15oA9Iw8iQ8ECNQOg5ivsMh6etZG84fCbuQ7SOtobnc3vR9DNYeM/UgN0k8MNyX
CSxp+qHZsxyC8NnQiLHf6Ybq2xT7tH2ECExJExZren7/spjsgn0H7C6qietAHLIMsQJdvYkmJnZV
lTuGv+Cy7nBJ0eFdabtctbrv0vjehpBl/7nm6wXydDG824AfPPQsbCNM3W0jrnjWmTBL/IHqCNfm
v5KEMgipiTR5KnLDvsMLfkTd5mmmo7ned36cXjBKrPOwQbbhk1JcjRzMETBkanj3NL5raapWoXgi
YT9RPxcsn59XDKOmoNeolB17Lqw4+mlJ6xYnPcNH8nA2/AyE3BpPnQy8Kp+LZMRwM6x3EeC7/Kf+
1AL6ay0E87erWt1TjgTRSw4rg5UVMqQUHt511nOHQN0rpg/vWm0NwYtleP66AyzdvSYAopAfe78F
HSOqgCUwS9zC6MQLU2B71mGlKd+Or+RX0ad37vGhehi7yPWvRtsXrXvHQpwZuqBKcqJBzVa/Y+wl
Uzmk4E+FHUz2W+5c5yLLreMl2+wLL9Nn9smJzEZkTHTCOy4oaW5ffKifA0k6zg8PHKxzjwxDhbM4
jWjM9Pq3mEBZshDeJqkTCEJ70F2JxiGf/Fr29xlR1uTuIBdzIWRESYlTsIJXe3hS0QFOXOr4lu6r
0ID3gbzWaCWWiZCwY7fpnAkglrUZVfWhgKpr4DDVxWZQSm1527VulNK4Q2i77ghAh+s6LF+hp/A/
G3eifaZScymKqsomtC60C9RPY6l9MF9SkxiIdVG0RRjSpRgv3prOQmHbu0OgpXMUZqGNWAezn/hH
rMBLiyWNyC27fjiGGDWkZua/ykCu9PfOoFdrofrrMIMRD6WVxPDne3zXcKo4iCffGN36VOXQ/T6q
c2HLQ/JbLAQu4XKSi+FPWLTt2ioNDz4xyshyMUZMbzKaYjJIQUIVCQfhRf9eADL7UFFwZO523msH
r13OotnCWS2FSDY81dctI7sjeFFy2ZHEDMne980zMsYL9u23S9hAIik8q9+VYCpqrxYqoPGst+GT
fGJ1fW07g81Zo1qe54ovRgFCcVVbk6XfDRyzGmEW9jfJlHoLlE7ViaKnBbwuBPVKkCoaG7bhGo3G
QCvKHBdVzZuiTD4VZDG00Xhw8zeP1CBThoNW6X4hX3jep0NRmshKtcL3JSi4JTkFsQcbMUc8k1RK
pq4WJTQ4n/OTCxjCZ1SKwiqo1amUqty+wLkLjDT0qxSQIcwE3/T3Kglk3SiZ9eVIv1USiqtkae8I
CWFUfGWxmXttKWVHUmCtrzEA3UUvWQ7Q7zInUyXvxsybJ/fgoDSsjnOPQDo+YWB7mYZtWL996+tM
dBH8zQgPbNyAOZS0aV9CNdD5iwRdPWoqF2efhsxHhGoLQMVB/wqsdtHZej9n5BUBY2ldFD68WNxT
6UrloN2zI6vwZmMvuDmroL/OctZqujT/8M9ngg+lnGtT68deVRuM1/wK665iBCe6itXkqqt3ikUc
QKseV0phGLegRcypl3cQSJ+fCDKhZYiSVHC0mADYdvtU1rhHVOg/S2XtHdR5KWbNnY+Ky8IDq2as
epE1vWjBeR7oxMyiYtIp+zr1Hg0RfMOzpfIPPToIOmXpJVCdYmzF1lm8behGr54exTMoKy+OPg24
+6h7GK/mg1m2phdCmSoXgA5FbX0FjaEkKpeBAlTQqNQdsCV4xb7MRVToiYZECaNe8JpTtgXF6v/i
IQ/U6EdvEIcZB2Vr8MduK6XIJ9vLcvWNZfhJtJxBDxnd1QJQeg37/9faBdqm7Mk9lCXQbvQiROFG
27nqsus6/C2qNPCgx/N7DW660NTZijOJHhlzSz+01flXOon13kYEPFGqZc0jdevs3lAudA6fK9fl
eg956/sV6p66FZFOv8GbMqfk6+K1Mu9qRLPAosffXGgVIZR3p2Ziuu02KNgHjok7xO3flZTfAn5N
hT7denl6PMnt4u7R/oIP17kpskuAeuW3+XVUnQWUqFklSHdEeWEAx6m0d75yjtYcqXK2oTNL7G0q
iBBPHUYPSaSo2JKqxLThtp4SwmeQG55JdTP4G/WE8LE0MlHUs3HCcFQYZ9XOfrXQhL3Z0ylt8Gvl
nFII4uF+we1TbgNs7SBh7ZkG4n1u9qvsH2qQxu0SBf82ED+i8wsr54zkm6KI47LjVVrzSXO16NjA
0mnVNwcoKsVDdV1q8JigdiWG3fkfiF5OmphEfqrH75nQ2ZVU3dhQtywCsQ9PlnaOO9qO+fkFjIxj
YENh5f998sasRXQB/V7HRx9xJS2ipudGCuvXwf9SHC1rYQX7CX/JJTCAU7wYjjuwBkgz9rXpB9fn
qY897KOwAj1w5eDZ6oVdaQM/FHlTPdDL+M5iS06LqXGU1ZYd4GanjLj9NhpxpK3L6Bq6ZgRw4xl3
Z9bCjUzjV8z8pj9MM5h7ktF5qiS+9dK/0bd1aKlEeYoRgX0Cmm+JQPL1kxeyeC6Q1MbdFQQ/FlX7
jDEyws1PIhRswMO7pGpiwz0Ik3JSSqaXtVv8Zk0L91f98zJhrfpZonN1+Nje3Dq08ALRAhfmlNwg
fRC603haOZHB3djS0lmRBuAIsLV1Ub4TNohE9jLPu/CCyhIXmS5a/iYbAFoT1ONTJ8BbveAXCygi
YljLhCqClehV8i9b5Q4Un/Lhkhf2gRPtrBGpASjQntkHSWMMaSf+ghCR5NfryU4DWDQ+23r/s4rh
1SdeSesraOi5ZPTHInbhHXNYuHc65Ii+QXlHdUUVbPZBPODFFUMWTOIG+a8MMNYKC3v8PLKv/Ale
DI9LDDKm5vzbCiSeT/Cveo/yJUlZIg/YzTABxeVcmHFL22wG2NKfFbnRa9jiUluBHgyV46xOWEaa
qjhwGlwwZd1OtpotmxoB8PqDSDUk2mGUmOffVvyUaRADCYJjWRhwYY0676lLRo+YMJUH2KacCkdU
Nv3be81Zm0KXJqXQ0cbkRaLXzKsdTuBqr+siiWPg04gRAgK+AorVePPhSahhp7Zmeefw6gLJBSam
vpb51r2+7asANqVfcPhHKUir86ZYD5YuB+F0LYY7X5rP5Be9FUudE+YFVa3ZCKjBYPcNePBbgOFe
nB6EBB5eGAKw5mg5Wgm2RHFRJztzFXU9vWP9wndO/uSJApzOckQR7nWwpikf14R4iONFP6h2FeCD
IBoHUYt3Fy9y6pTCQXba7fUeJRYY+8g1ZDOJxksvWrXyE3YY4t2/n9xe7ltPvl14jHG5DFL0GlyS
iHXDW03ewE95R5Ypwfp8m+nGBQQiabdWOlZzXeLJfBpZicANQZDMvXhoW7y4B2l/syy8Zppumu18
TFmSvkHO5HDEKJSjN6p7S+vzoQ2lWXCofdpL19lKEDBtgxZzoRY3aC+LR+CP5u37GTtE6piSYLsL
JX8fikvnBn92lLjSrrIQJLDnYKEVcZT5KUZTbILw9lv6pP2fSMJD+jVwlmm3OG+mJ0abNZTJ/Hx6
rzhEYEtI4wJb5jbAQTYMR+ezG1frTTYmGUkAxK21uspUlsHZe0qximCb1J1LTj+n9v/O1xdbkBHF
dBmSham31J+yAvXYW26r8KU1gUQxIskRegp3pLyrWDCeH5TQsfMnMeR2sbotNyPq8kj1iqQalskC
lZY630MkGWsy3p2KG6hblHBDcviJ0/ulM29Q0w74057unc1HQRvf3zTLdhtHOWMZpWh+fbDIC4aD
oDlPuOupHq14yTQDNtFY8UwbiBvzZ9PZK0Fc3C2hfBjJ1xUCSQpFwk+Yk6pAsnACm60UrVp2bInM
YdmbKg4JswVBTi8KWGEe0/maudzPLbYPdc7n7AcroZXz5c9uyVaJjU6tcmCbVDtcYB1Tspcxzvro
wwpkhw84WEFZ6wJB6S+l129qcV0wdPt61MkQ1ylUNHv4jrkQS9wO4ihzYOnSWpd3miFpeEAp/jkL
b/ZTHlOBw5Rysjl/lMGs8S7w37F8Vl0WAbI69yScfYvUHnCLqGrw6+7v5fUjoOpKbIR349LIBiTP
kw7qEyLBXs1TioqFrdABClmP5/aUGfHfJ91kpS8YtJaQh6fyBRkJgvZDO0Wd36qQZNoEHjacFgCh
aBiTwPeO3/nGlcL65V2buMYzVJ2D+GtcBpgAceHVgdjC+lOFU47tr4zLO7qtxEMZBqcjHa/AW1ui
X1tSGxmNlW+YtPdpkKKkK14eKJ8eqwp9tGfjUQamOBdxS06On6RSAN+5UIdCqD+/G0xBD5tVZSF4
kN7Q+8DB5TWvzQwRFiFguO/cVy+RZbOMQOqxYomTEbLlqcjVA27KH3wn51K55vW6i1HQVrTy1hFT
K0P6sUW7lsgsCz5flOEv0383pP1AKVoq/WMIDxfo3C0LI61rfaUOK95uD7L60u8gBR2mqhGws4AF
px11x+eowVMYJINkTXn9PXUD6GA4PxcCOVFtPj6d4aEys4FCxLEQ6vuNxBBgztX3gOwN7hP+jNQd
jee9S0JJDxAwKzryZ8qXeZgy2pzS7Y+MrOBVleEEvEjsNGbhrPvwQKlvRsDzkxC/aDMRQ7Ak2zke
aPte18wRxwXqVrhdwrx0xamgl07ysK49XcXjUXpqcM+rciqIMlILCG5Y8Gdj+xl5ja0qVvwA/WTK
m1HQIKKtpt5WXzMBaS4lylEfmKhUdPW0XH20dfi8Jt6BcWfNNdI/yOJXZ6vG0qD/UZsVk08rbtex
lOJO7x/eqf0EWfWTuBFaKBEv8m5/GcbDCVaf6o93RMZ8H+JupiRRmZpTeEwJL9iIe0F7Xjo5839X
pKC4hiogXIasgD+YlBrufpG7dvd3tR7ayBUnly2/dvL1s0u/ysH3UNbB0YQn1b4PsJ18p6+Hi7Wv
ANdl9mAlQvlIviGLrcmztiB9NvGxlRdCAlCetW29nVDFr5Lt8yH+yZCOKkcvPawyqTBmdCWSpU4i
SaD1HFXjlJh/GiYfw8TMt+7FNZmzMHe+KRKJqoo3jbKHSxj1lKiWo1uPOJdjxbkwpuq2E3VRCvJY
EcIKNmmm7gC72wxoKfp8wG/b3/mU09S8A3VI9efDNQXAHo7Olg72/PAUPF5E8H6l60+PrEMxO4Pe
JC6aqsdKNe1H/fasvxo2PP8RLr43fmnkCi5id8LVlVXaYuPHRJf4PmLd8OjKvJe63VzjVQAVn9dw
9nCGYKvBfG6/KmTyO3b3Aczj1cyhaxsolNjGfuT3pPFEd4a/GWQGCxpU7rz4Il1He8klWZI6TCzq
R19d8Qd3NUb+tHg7OLK6Pxlh+iIQW1E8Amq3GZft4U2V1uHGsR0NhEufLYIHU6/KtgyzaEpXTTeX
3SZlkY150azeGne7AX6KVJ7PH8uEvD9bSqjNonSiEJeol0kSOybZMd9AThcBB2aWDkepJ1jmzFyh
iGGxLsse4DNGbe0pPsG6dbONIKLZ99+dl/EzYOdVy+JfknYL4dkdkbQgPG2zptfoTJ0eSv01TVpv
8QBLOx8d/r4tzRXrGFc0sks3aiSStS4VMckvs2mpb38wSPXnlFOcu5eu+knGy+4UnsTr6eXPNCHe
C70yrdsfl106svciZtzM9/++1yFg7mmpqbnzhiQg7R0nShxMU8X4dHVIwQq+1L+8tzihyUFcM9iV
coPu8tiyQkpQijPBoJ5mwL1K/CNC3r5pCYcDP6VKeQJbkxo/b3JTWhwlUfdZ9iF/wysoSfEPEa0B
VefcDQoZPc1BFC01H505nRT0lJcfl0l3Nouf+dk3dgNiymvvMh5TqQ1yawPTNOmJmq5RZQPGFweE
pxTZIPTuZIviYLrzSYmm3cfsq72fBZ1nsGBQn9QJ8nmdU0+u4Yqs6QLKaBzfHAiP3yUVl7vA0/GA
ATRtMTTDIjmlS/L8tLm0QbVKcDKxkYnUyMIgBJceXfkh6uC0sZkVLTWnOQJ4ceom2MGuz9EtnCDQ
WadgZHQTKtj0sb/YpYJXsMub/PHyZNY9iFs3Gg4eIjFTYnKzD6K/r7/OB8z86UkP2Ak2pAjEkLI5
smtWvk+cBnOJ6T5TNI5HTerjNCRn8vDep5gj2TU5CbKxIu7eA/FqbYBOxEnSrZKf2jd+0lAH/o3a
5MeN1Fa7darAEtwCr9orgxcnS3KNcpQCUNOooWXuuMo/MFIkjwukA1DCFrZK3QBrB6H1k2dok89J
q+BlBdLPw2uulmVHYHbo3uttR5dVfj/z+2UkPCMgyaK1eQArTS5Gwy1xPcqQ7m71s4EPNnwnQSYp
1yYwtTrfdqFB8FwNHZI3chnoetpwejhctN7sXEEQTEzufrdMN9FahdTZ3SzIkxOOJ/AhkgpTQDMc
10Jfl9AWVfh5axcF43U4YWZOS9/aH3Ba3cP+W7VN+8JnIDsz8p81XozEHtu4FWreFVI+JUAF4PaL
//NlVb65+ogRwWfZB8jmwhVU9vECLsY+cmuHrsuxAhiSq1b4DCHjh03GUl1TpJyHgo8OpMJqLu8P
WuksrjVwqsYf/0zSn6ATzKgq9o2gkUl2tQMrpr4gqB3E/iQUT9Aq1nZUCuk5hgA8FuaOJeZZN9Lk
nflp/fIvA3DVdk0bhVtps7Xy/WZNDISVOEjW3H0jo9Wtr+M0CuJFXe96qRC+Ok5bSvgq4rVP6C8R
Fee+mbEa2qfA/3jWB8H+UDF6xDScV59dpJGhsnYBQx8Rcj43yNypZMsZM9SrlN56Pi+Z14bK4H1b
UEWmNdjEYLESE/q2EmdOVhhqAZ6xraMCVUgpKnjzyjcRmqz/AZ5Ogvw83m8nWNrwEXAoBeApAbN0
ZCO/i840XWKUFgIdwYLqNhNMVYaJF0yjYloBvi06kGLri8JbGy77sb3+RwAQbcSJFl8GpZdN4L0F
o2afD4WFeQCcEjzk707qexBuF+86OYi9uP+6HH7xJnsXsGtSuE38qJAz/mE3ewyzIs2XbI+wdIEm
G+KVU8vm5+pOU8EP37miI8dj/zwL3dAkPwuXAjhlRK/SYismrcXM5qgcNhwKoDhqt1dsoynJRija
LzdbYskCZKztew0RruQ9l7DEI31jm8Sf4htqIpRzIZZP6YaVZjRsSl0KWlESffOJSyztQxcWoUgd
Hzwx4eibSH9LVFEuQpBhVHjKca5qlSYhbqCHJ6w0IR8PXRjMRUrFPXtTkoItZQhJVcATMtb06slz
QO+aAp4Fd9gb3dWZbPMBiXxVn15FI6y1RwNDatWZ6Asllnpkkx71/sf71vLUNpcryFtbdSxL7iZq
71wcdt0hh8mVmewkLMTt4xodPB1QazNnbuYkDFxWX7zixNwOR0wDuiQCc2+YV4JzmrIJHWglkHFu
/fDYjxsupWtIbQinZRh5qL+f018siHruGjqZxseb1PY3Agy8Mb+KX20wmXjBLWB4h1t6ywxvNfqg
igttRSzZXJ9IJMc3JpfCKRFR74jzNTO3RmnCQQpdWsIzKQ5ipNgdAVf2JFkes72wR5+dJHrnmeSv
B6H4nC905dFLYP6ALt5j6WQ0v37cz6GQYL7oxKAvYU785/FuqUEN7uaaCBE0nl4jf3TueBkG9yWL
ne/0iqUTje037GoWaJnZXbh3T3YvEj52QCxdWDjyZ0N+OD2znH0kUBCbiCgzfMII7vp8g1qDiHan
Gg+ao7NOFAmscHF+axK6YoUfxkAD+FIcIgtbw3zVODb23W8A8ZLBv9jhQpv0p3fLnrR3lql2KD2a
2i/GY/Gk3mHEJPNuNxRbVqqGYToAAAXru3azBIbIsWESXRSmhb3VnRn0b5Jnd4n9NfO2+6pS1MCH
ow40yBM0D44HONnCPJyhw49Z8FHapj5aUlpWIveL/n34EsHakl1mpNmjN4wqLQsa5a362VET9uyH
A/5Kt7V5HIfwxpN7GJ6r8mOlUZyW9MBa3f9qVqMrA+JXmHcrb59liuFzxVoqlqM36t2L1G+3HQaw
YY7+NeMWqWJ+nQpY9ITIpW4YGf5yPPOyRmr66gTWnQJn23xAcZCHBtxGN/fK3PtgFkPgQ6PpYSTl
POhydAF69LtWOkcA3LBmntk8Fg9RTUrd7+Oa55mBT638YpAX+D8TtUlt3MpbKB5A4kQsIIG97Tya
YkOsEw0aGZ9sx4fBvbZid/YgC2ygG1SyXAf/mH0uIHU7xeqJP3DY25S0AX3EoaVUPpPWgziTgPay
LwhwnyzCJuCwqsEpDZXb2LczwEBlLddZRnIXwfQe4Mh3weozqFvKEa9wQ5QQP/0CZrUs4vTNS5pJ
WLUetEqhIkL1dlF79iKPLrAk6e8rtIbfyqJItYT4IiRo02Bz5BOx3Ao5G6PQTsuaQPxmFwrVbO90
avcX1cMAxHgv1USgV0D9l6EA/Fev6FKevRozg+uPHPeNxXxN/i7PWqxpLtk2QZOkOI0VdQJLulIn
SKXO6JePVMM9aHNUlRfiFpfyUgfDndUAB3PSWeFtgd9oUxECtD1trDvnt03PCpaVdXgMF2D1BYr+
s/YE4C5z8lOc4FIjlQKeQNbJQGcAvcxHle1gbMzFCaZ48bETVvHIys3VU3rGCVN6bYeFKDQcWUUC
SR+aKHHE0LHYA20Ksqk7ZmBmcq1sTG/WmWXhDCPEuyFDmgJtFzUTEDqFM3gw/WZUKvE2ruN0RQHh
Nb/YxRJ8ZOuDwxfn2S9w9n7BrOMmTEjoBAvWnX7jpX/QySI8v1QEXLfbGJQDBdQg8FX8hT3n2TH9
eTerW+eM/OX1iTsoHZx5ccCxXvwv72/InYnGHsxfLn6bGOIgiq9beb+JkWZuq++HuJyINHLs4Vxr
saTMpZAzFnMdTMc+qsaVKXF/8XS+HTijzqMizfvgEpoOYu+Z1aplQuJD+HpUZbUgBg0Cw4oyKGZM
hgj52OBtbNZ/h59UFUg4RerUIKJf3BqfH7kvW5sFwvmapQXUYoUiHM8WRgngE4r6Miq/9ZhPZ/uC
rkQlQ6FLzrdtTtewHJfKVtlzsImCPt8I6MoJmrQuynUTdnyeRBFGhUhgPtatIJTsmV0ssmCeciNs
YI/nZWME5u2kGFxAetuFRgGMdHpBP1FT0MNdFaLXwSRecZZN2kgL9hmNSOsDaHfHrcBtN62VSXim
qOv/T50wvku0GrgyyV+azQNDQKRQTnAux8m7bpeeMDmKYWYQc+hhu0wtG/Zik1rLg1BH50TPM4vJ
dK5ZNN3rX9YLb9820CEM/37ZYYuO8L/QXlPJrKi1vrbLlgcMq9I7OIsOUKQIYvU/xyu9WXazhrOd
RvePhQdp5YsV98cOPhV9cEsZXzexCsD7MPM5tTTtO4lDAQNXvMVmBgzRqpjh6qNs2KMoRwpWDGik
St3Iqw3uc6P20JTOZgDijRFjKTDl5+lmjtZ6kLfBBhrWjfK5dksRAOaet2Fb8DFmF0y5GsEnDtzG
tOc9gTQdn2+11/6aVFbTmInExHm7Qkb9IJikXb/+cxRMOHN1wLaFN8YU2SNuMug5Vi5avt70oBay
rcwZRqfpKSMMqrEzPQRablXl0Pv+eRTyvRZRUtNEpTqNVsMkDWTA7mHANLJ9W0/7YPSm2gwCJ02y
lqXdw5zYwrkWns/Um75soi3aZAf/rC1JwJU8m7i0MDeMHyepWabF7Plksrv0EGh6COu/vJXogv7k
E7myfeAwW3NMYznl+6XI8g3mMhw46GyljBGLFyafAHkfHHlDtd2wyEnYxRL4G3dGnM6UorEue+Db
E7crJpc3kx1US+nqB7Ig9SDy4ZpGUM/l34eenHIIFF8ixIWzEikoqU8wzKw5XbVfPg+v25hWlKsR
1wk6S0APMejrhOyNvbxupIvqNvlK+AU+WaCxqw3DTemoA4hSQAPfz0IRNrpU3h2uFd1l/g1iCOgc
q8Y5YRM+KKHm26SXnxK8LKjexyUo7evh4tKIDx+K92t6io8F1a0Cwj/96KIlGzAhLkHok3GlNQvT
i1PqyDQHHKpcWowV+HcHbU2o+7VDXc67HOasCDERcu8txFAAEfhepPdBVwIUrshBY84lk1Vjob6y
bIm1iz/AT4RGrS1vGUyytD/mSH3UIpGaZZN1GZUyfo0es6xF5FJZ8PHoO9/QihuOIkaPzu0GgLIA
gd6QU7tBbvulZ2wosYoX0+/dv14ZbYNIrPzOPR8INTWDf67Oda+sS1Bj8ynaCnU+mc32eVpb9dFA
YxVvGGBBMmU4HIJxZnP5u1fMcOFWxkDVEtgI+s5OjrflMdWb+pqo1qnBMF9SEqMkF3utUVAaHFjY
3DrrsNNtAVhAJiorfrInMUS7YOIMLk5ztwCob8Cw1v61xJgKWV0Q7cHCGp/s4687gcxkT6QoUpB/
TN/jDURaZrfZW1EItNDMgcLh9bXbm9DLP6PIeqFUJG/xrAV/XspYoqtW1EU6PvbR563HXGYyni/W
eSi7y9E+sXxSh2YCckwiMAktF0oIX59s204RBXSjCQyec5+A3H3Xjb8/0Re24zjjrGpbt8OOZnJG
CBHu8FnH/eyadbDXbW9QIkiQYupO+IRF2/zHfwS0GByKPb6Rb29pRVUtS6rh/rYzIEVLqSb6W5CP
yHbHEPhTWMQT/+nD4UhKboGJvzfSY2AmoiM3xXH/EimM8VD1JgJ/suhwYEblwD9NAM/X0ZmaV2su
MxO+A/sgr8I4vgiEp0lp6sU/gGMG2aKMIlc+gYYybFrOP3+EL1CqLjnEhydpLTuS69IolIV+3aMd
zJNHTlbYv/SljzFbzVeLPFMVq48EJ+i6cC1ynvLFp3Myq1z+SwVmm57scqy09xII23JPWRbq9sDL
UWzM/wUirpEIpFtk96VE5F0Tf6g07fp2tx58mijHtjSqFG9F9/r6s4P8cmlIluZoa7+4HOMv9rJM
shXP2k2RUHg2j8yI4PPU+d3YfmrlES5qL358f9CWjmUIt/V2Dgqx4qI6cv27o/MMsB2/0Vf3XFAQ
AVzpRQeZ5bKfSwSLQRWwLNdXm6TgF1FBrtF18YkNQcNHIu+C601aijndfNAlTXBi4nZjMXl2GpF5
A+c8LTqKMxdKgwxvEtmKcWSovhHTib0EaZRh+dszFkugnidBBhgxnZJ/0Ny7CScT3X5ZFJ8Mx9xy
5Gidg3axGdChORwKRpoeU61cm9THv/n+jYGhin3JrFJCKl5iVHdA77h3c9VoMOV5P0/0cK/pmG7g
kVXox0maWh60qtTOWBOyR0cZA+mGyMXVRPjQb/BHCZxNvUS1KlvdV1Co6ADvSzFgamW9+6PHRktu
MGrrdqy1U+tHk+Elgg8HJb9Enr8RB8YpOzJlNJD9YNiyRuDa05xWTBq5gM73t/IIyhdJA2c6koT+
wl1tWHW/hiCfIyDMON5fXRsE0Uoif+UoSHPkfh7bpOHAbA9cuCAcUrjj/1JEv0OdFodeCVr9mzuO
t2PbGP8d8hlK/j4GUxMdTLmMsBfIfpUWWkEBlP5KpJrbIN7XZWGSUDvw0D103ycLOw+2jSykVolS
gZokrZm8ewMpKHDSNwOdkXQXJrjIW3FYaMwYah90ZXnw+1Oem4AwBnFOUMtGSVJvlLp5E8HKDbA7
GbqNaScrE2kVyWosNtPszbvs+oH0eGPYHHYbNtQQV1QwHvvpUc+K181xEc8wddfpEa+2R+qWo0p8
cRK9zx+72nBZ1UN1VjjY8DcD5HIafHaTvdrIp8/wOIzsDMss85CYwOQNljmetRQlzSw5a18waTvK
sCFXPNcH+7iv94uik7dwjDF6QF3W06nksWr4HtDOVv0iY+e7MJDi0a9xmJraHohVlzyz1cqgyQ22
FTA5a8TBmQAf4QnHK3uRTHxasgEKCRHMB6UTxWPYKUS+l/KJKzbZYSdH13DypsOYuLXlo+6dm4B8
Gk88sE7w6bLz35gl3n+u9/DKbL99+/orGMcUBmt63ni/EbH2F00mxJ0LjTKW28ZJrfDdOjxsO8gw
a8moTQrS/vX2N5dctRY0kamJKU1KhfArBfnWSSRunw6uo5XpFMQfjPr6fvy7MCEDSSz7zZ4k4y8s
/JOkQ+oN6YoXVmFNFSzb+p+Nu8hyN6aAZ83sMMdnx1NWawTTjixa7Mda6IZsvEtwpEid/MHNeiTu
chRL09ykS4bf/+mgLnNygqw/pfeOc7boL5lqTO/icl4h5LXF4qAU8TsK1xNW5d4Pqad0XOrEcYpp
XQA73O7IpeIe7YTbOLS+CVsG8LIqZcDlsQ0BsAnv0h/O1XpGU55QGl2KeGaUQO2NuZzU89Pgd/lI
bCChZ3c+7V1Nr0GtDMrM6X/VtvFX1QzggFU90HnM6PngtGtc6eqsQw/bh1+G4jeQBAYbx6Wx7AXA
9W7QQ0pw8oQ/EMcM4J3ghtNtNgdicBG0/zKvhPG+WTOAEQSRtAfGLQKAEf0sWZswLCfE619FM/NU
u+ONyu5xemqSe9aBjsJjHCeqiexkQ1UsYIAGSzf4AI1Me1JzSpm1Z9iYOBcCuX0KKLitPfvc0GKs
FoBnsT93du1biklbFPCNObcAG+W++bUAefDE05CvR/e2Nn6JM4pNVnBRVdFE4PHOBNUAAx3Pbj17
jIOVRMsKVpphvjeRrC5qGOGPJ8dBUj50bBQ9qwZ4onN8GSo2ktsN6c1jLyy+qNGZlIFPY55SjJsc
2HOI0tTWnY0pGBKgs29sRqTiz8fvxRRI86e1IsTmvIktuFTiTkbA6/DM/Fz/A0XWF/pFclmKZEid
9S1VKJzCRfA1Ds3EWzVTsiTELFjZOIB4DFaRqJt6/l1RYhjJjhzuAGx7cnFBbusYwWMA6LoUiDKM
udBVaevCJ9OoCQ4lDHqrqs6l+YZCQzfDE2dg5SBV0dmW+xlLhrEGDjGlC1nxOp6Fxa9TW9tBmRvE
txwCopk2w2aCcH14/TBQ6wf23raktC7F1KRz1rEGymAqQbbZPA4Q5ZJ754ozaeliZH47SRosPh2p
UdE15Q3rmHThPVeljlin7XJlkpt7HVLiyNj6mZj/rqv30cwOIOXWIAcAfTmfCyp5JPjR1qXKP0pB
VnGzYU9iUh6ffAR5Mk6hZ76VG2jIagZ5l/KIMSkt6UkxBJFgb5FZp5vBk3zYRHBIFXOB4uZY2rJp
sqsOvODN34TnnqFttbmyHgwMivCvUs4dcXmrpQyxaVK5PA6mgqV6/nH+w82Mrpee+QmnccKwInYU
/8LwPpFsWvufrErjpgHk5H6IJN0LO3aWgPLG0rl9q4s80tFuohuiXdY0kACRoLPyXuDMIZHuOuNz
C93d3+hbrmxpH8wOCzFp+HyItBfGzPNrhy+4xH/4RUVvL/aCwqXc9f7+XeVW6gk4JtQwpRf+ucri
CkY0UeF5A6SkSez1aZKVeqFD9Mh6z7yGXSJqKyQ6VgIDYI4336PSRWjI9BDUFJRQS7hGXubn1ZPx
1e9+YK/afxf8hoYWok4QJMPEqHDSAzvHNaU8HbD0Fjh7HZPx3ozMjikQT7th0xBB5NrKjPNC9591
0z7cSuIxihF2EWVwOhYBtxguGE12n2AHRtv3vvqHcB5qTN+0qK4/ei4msrAt8k8etZGgIiVpoE7P
TRB0w64RUONgj1utqq/TxwmR+a7ijgsNy2HBXKaLFHSt6x3ThIP9nyyXRe/e65eLybjoWalslAeQ
k6FW3iaz2XVXu/7LjOVVDzwsNLTUsCoSdqFiQ0q14Hw3HWgOan0sjbizKUiqSX4BG81hAwVIsMsw
6nz4bXSqZLvyQtjIp42lEh00Ns9A2fvo9Ewl2rRLhdqnGxFsoBzKZNtEdF+Lq2kfQcnCtJDCrBzY
/X4I/5KggOl5VydxLaBkelSxs66/ayHrKYQJxlmcd6s7pAPUMWBzcN+Xj5Xt5BNF2Je9RqOjzxwj
0AOj7s1tproHWnvn64eU4Wim3egDTcVboBnFIEiU14xkjSG9i46n+7WSXiDDzTvI14C5yGtgRnlG
tl/b8SCT9WNv6NgMM0J29o4bT2fCIWfB+RU4KJOPGCG318VCAvK/xLGA5nqZiTysBOzIOt3WsMPf
eJPWSwm9TtNburvFobXmrxaw2/lM9ywjgl9GuYsAySDg1yLJ252L4QCJNLNK/ovkH4906qYG6H5J
gDfbRre0+v03sqXOAyb42Q73ZAVl2LcPLHBg9tmZr2IYbWi2FvJV94hThikfMJo3mk5qkwdniA7f
JfbH/Q9u1OCeWxSyR+FWvmmn8OqIDfVLjMZfUHQvE2SuDCoqDkhr4TmWLz3zrWJPh/FSqm/WW0fn
DDEbZ0/knAxiotHAy7vS4734liWkpicnRpK8pPyC4P/4+oxbd85SWzqgMrUlr8GvhYTEkfIH1P7C
HehdKbIafqME1Srup6mNNfra1/PdDETVcISVLzMMMNKdtZ6Sorezl5JzvRxNa5Fg7bMCay9L4RRr
Stk8K2ltq+1LQTGNuP4+OVWgSFmBjBsT4dEfAKBMslOMRyG9zw+AF2uEgKQgmaijuE/OTIFuLmGH
TEKqAwjqFSYGQp1xGjHudcrRFoRXauVTBFuYpcIcctf1Pnww0Hx6QtE3BMu/kgvBN0nHRBfvjrbb
WfFvbN07zF09dXPTwtvTtEjgybCkVrjk1/CKGxOvifc0jkunm8Z6PRhmDXdmFX8UgtTByEAFXod1
B+Car860ld+9kpDXKztj2klP8Cg7RxLgKptUjGHRMLLlJUgsqueLjFMKQpYCeiuIBdbiZRTWpOYc
XZW50mAbgJpHNcFilcSUIhE3Onm/K2OfEN/1LkAx+7sa6CXijcx9N1fS8mCrCU26wtR1nIkbrqXd
zEcXtie6nY/8w95d9+mV5JuyGrgL8piVRtHZccf8ds1KlisVhKpX91AEasarptheT8E+ZnVw7eEu
SJrTC9kO5yUkc5FZYC33U02bsAmTfrFVVgNmgchoDYvLNMUzz1tF4X28idWC4qa0cmOFPGqE2y8r
nKdGG1T2aW2GDnY5YFVKVq5roFDIPa6k5qmJzOKZLG4GPYFbVekOKWkTTLHdsut6Lhb26Ov4uPAk
O1ZXBHEnyljIPEjWI7ki3KZcRm8EHwSRMFd6UuPfm3+JH+gH7zniSNUBv0ZzmVb5SMP3jkMLFnEl
/uo580+jmfq59DGegOosco7MEjTPOFcu2wyw+q22LhYUN+LYKFmGh8n7R2kZr5P43NRVh+0ULikZ
t6gqCy16pE7py7471qPp/xwDYt52ku2aK6/SdFcoqWdXTLg2Rj7ggm5L7gBCLlB3fOW+cRJ1LpI9
4skyUFut7gT04kRhTIoHtDR2+Z5BPBGY4wNU1EQLg15H1QEK6lhCBHDBz80m+DPYVikC1nLxBZUB
433BrtD/TDO0GktPP48zZvedvx/qeYTlzBf2mEvjeNTWGnAW+WBuJS0Of5sS+PtfN8y7piKtIeCn
JscKVxBs+Whbpw1I+WzWDDyxeQCrWlNUxZGxlXl0s4c98MKmNnR9zg0Bd6fg2RNRIoNnQ15jAjxf
ZvbNdbgUu48j9unK5U0fC8OKVNNLEVoxux56yYonFQBysZKMrghZIqUR76GnAUtFD526KI4sfUie
3bO61SKIQ518dpBi65hsBGEkPITGin5cCC8C+gw1ZIFozYybJJipl/rpCSCXMsLpHJfWyOLnx+tC
xfi5++4WHkyMcWDjBfUElHU9iLKGEXoDqkppd17KgxGi/MVbNMuW9UXW0aGbLZayh5uRzkH59Nr8
UnN2XTA+3ACwgqZO0yQUjgkb6hBfGxz/etFXKL85/PK3fZ4Yv9kayN4I1ELjbjd3RBlOrmYQ8r5l
uFWA+Ajy0wiB6I64Vqfy11M2lmhSTUnmwfc9Qr0g1WkFH5OO7pzatK2PZ7XwizA3eWGCLbwNheLr
Kv/sE5fV39UFzy2dNf/GsiGketNiUtutacnADtyusCwOd9CGGG3YodpZwKqYbdPZUu5ZG+AjoX4g
U7WKYo7wWqvDWheJjBZnvp1lc8IN0yN0hwAXdjg99rOzHqoqleZAq6Hc33ySYX+ZvBBg6Mmjhdq2
G5Eoj+rp1p2SPdN86M7ovWuRh/pxk0lbuyoOw9FfUtKDzoPs5x8McwlhXKGIeM3xp8J/nHHGA2jf
qlFqmyQoUK/QGTTojblJmzVtjJCvF0V8QL8sCN2XAvbOW53B9emvfcvNSZDQD+KAOz+T+uWhbsEJ
FklgyRdrf8kwRg20lpklKHkfSJbzW/SmBZmN81i99rfcVRd3l4PUVoy1TIa7jXp1yGDTM3sW3Huh
hpwCu/bJggokJvl+ZF2heH3oI70H/sRyCWPghfMgZCUo4wLESfGKRuY1KRnEoVKL3s0IMLMSW84B
7wgbEGrumRIJaTSIQUwDCBiPrYWs4fbRqKgG925fK2Ac0Uh+w1Q8g2thn15T8CgM4EESwB7u9FRe
P+o2Mpvc3oax58Q0L7vAfHL+jPdfMR/VtqyIpAFhxafxhZXyieieciMzHEFx358caFfb03WpZ0CW
dFAMJbYlviMcm14ojxdDBHJpFNAbkQW4qICpsNnxCY476iHVl5E3b05KFtCPGwnsAYR2qGgn2Hsg
OzpcTRnwkxkwynGlfusICx+Noxoy6iOrqfY/cQubJpjzJvXnS1RhttIYAPFZHuvhdM8f7ZXIj1SA
zMjsCKqrDKbNErxkesbcl/MDkrXZObkBeEwEltOySvmo3S130DZg5UMVfTJMEW1CGboPvpwbG/3p
wkvL4uN0X0nTvXmbLwPYqzXOHgZqSNKcFAlCBReZ0SZueXu99tJCGskJaRqO2AkaSILkD9bzuSPC
uGRTBU3jHPicuy7ddUj+uWTbkjyJM6G6qHVdxZplC36wro4Qs5CXVH0JI3XarRjnB9YuJXhGKeDS
5m7zCXiwBQBGMvsAV0orJjokyiTZt8xeLreDr93+OoKxEq7AQ0UbjS7umfvyCEvPmrnfFiFpjdZp
lAgRtRLGd7T+lza/ccsEmyQMCq46DUKC0lb6pjH7r+MgY/xVtOSrfoNIeKMHQS5gJ9M4vbsp9yZf
F5gW/lJn/Eyqo8JEhYaaNuuQD+TfOvShjDHyMtWFoC86bVV1cAfFwtD23jqCRbK3p0TMZ+Z5VENe
7kgsAHXw43yiZkhXm5af0pvxYToRPDIC9OhMdS4v0k3Q/jZfnSJ3s51ZTJmjex2QrC8Fc/cC2Q5S
UUA+/TSND21geCTqp5KYLXqyGavC8L+M9wNRxLIK5aZK/9SACvoXUo3FxLiQ7ocRPsD+tokkqyI3
aLDZ+J6dqu4p9kua9n2EE/QOAdnikaFYbMEyxD8k9GbEo4lHwO87ikY/AiQ788rrXRiLUQzEUSRf
l8I2cekh0cyabW0s+TGucBUkUE+Ow4y7jhX/1dGuFKM+K900KAd1PwUWG5NHKEladLKRPsqSCfpU
qtZLZBgZQUoJ2fUUzuT236sKjGsYI7QcFFKuO/XQ8v3dTpWGGHRo+4otSazb/xvBFOuVJLTk/pNS
DazQHwlMvxMXvpjkTLpXKJsIF5V68TSP551iXlTkJxIjA+FFhOB/yYJafiK9KlY7kfNaqmkWplDV
q55tHN1KK6WpXMuENDgaE6sK1d6ZrfviC3ldSRCSy+R5MoEtPeL5vDHdmdy7SyETPGAIMi8NBTRx
u1xrvvWhopud4zW54dA4Nt+M/9rOvVkDLlhf0c/8I5haq4AuoDbsETcMGQzvsamYrsNVqy5+6JZp
sHK7f28n4Xwhvo21sZbXmmfiaYAHpUHsdudLxJcrLPpkT0/CloqZil6eZoj74Bcy1aXSi2/+SyhH
gnfhEoMyPf/c6j2aGAz1Xs1fgaySEsIN4p5+83LxBziKOr9Nlwenx/AVOxn98mPHNaC26/Sk5RzZ
aa6wu34IjzcBJLgwUdwJmEJMOGsaYCSAFrRT5JlMUg58G1M9yA/VzM0k7PAOtKcNrO3HDF7l3Z0H
WkBN5EjJt08T8AWmQ1YYq06CmhS3TUwYTCVfMWmINPOAaTTcfmmbWNv6A7DN1WnRfBvb7Yo1l2vR
SqpVXF8gvYitkBBNSSBa6V2wKHePpnlsc/tLgK+IgVlI63gQfN/tDhja0Q6LB1oBSYXm4C3bgyK1
00VdfiX5O1EWwvwLSaya2h645o10rjNm7IoUFUVEZkSj9ZPOc+wbtPdekqmSii3QYc3mYt3twy/9
n8U801i4AVvvcjvchpEy/U7Ff1kOh4fZHVPYQhzwYucaftwe9TNUkWvSYdfrOs1YrDlq3dn1+yMS
DUL6MEIRDPDnlMKhB3oSRFhNYRVH8nwkkFEEwqBpX8n3VQKSzo9aH/cJsgtfn6reTqlr/r8VhtJ9
pFJygtLEl029iR+To47dc+BQ/O4Etm/mpdBWt+Xa2TN18/SHPup2c1RhY0VjodPPWsDdqxamwaUP
9GcVQwDb2EtyAUR4u8SRqLob16fzpZ/ISt7s+jjWpAhs5cqZ4VBS4csWkFvycZcFwdNitHohEkzs
L5mEplj4nLNJNu8nL8EYGpC7CtOjwpfyqGNqWiE4DkrfWu0Gqfm4/Z2MZLnlVjqKSHd601iw0KUT
1+eeh7JlQw6bbWB3d81Q93EzWnpZsSy507go1EBkSajv0P9InROeWc7GFlFJnb8mPegrK8T0AwlV
3xp4g30j6DNc4pVBJlHS4ITD7EHT5/3nrTp9QQEaMFxw6hiMz2x/MKmcSe9Abz3QwaHOzg4Hk02o
UtXISrYmfzCgo3+EdJ/WFtxX8IsY8TVKLKK3+XNs4S8iR4hT1WWxCq1Q1VwnPvPkgzbE6uGW4l1c
ZSROd9HFCnZ0Ih48TcuVVw1jGh8X3NEwC7gf8uS+2aWPTkvPDbXpbjtf1wD3NpT/AOm9t2VWO3fV
V3YQd8DWmsYpg10GaZJc4j4Iukhe055FJLXnOnILOy8QrxjILIbbvndwA3FnjgclofVR/H+jhPG2
KCORM5kRxcchE9P+fj+cDguNqgDF2HMMcWFxQRY+178IH6xgAogueRkYaTLLyc84oyrAE75ReUoz
GDGG2jMUAiguAmamJ/2MFZUZdmOqjSSOR1InCHwcRKtJcQI+6/8FVHPbW4eArpOyIJ7S700BzONf
SIC/X9FlDR2jZuhZGKAALNXsWzujutdBqVl1WODoNty69aUoefVtjXfVksSXR7L9zARx6bs9wwzd
K1qFum28rNNvZrp71j4qvwGrb+3sb+yp/jyapjQSeYUXFcGBq9M4/Sw7VXDpC+KROHdbsfTdBhjk
4X1kEDpNXQ1z9g5Gwl3MrrCuo5bDIQoSVrtV2suBWAL05UzsBp4EsKIPwkKuHVVMpKw2tjoUNrT2
dk1Uk9h6Cibzv7plfSdCj6yBvFD/ayh/mNMGhtXyXV7FgmdPmjUBrh0OcLkXIajP0bKfnMyiCuzP
b/5N73NLFBD5NhLTQ7YlnHmZmXQ4J7/5rX3pRyMFvO8i4uLLUcQ4NP1+CklgiDTOZq8Me/tm0MCj
wdS5Ps3jLpgZq7lgk8FFNhHLiH3E14J4priptAHLVinaoONYXHQRgsca5W2CuAQpMlo5AkLE/jS0
Cmokk65zNmfrVgJwVo39qUUYHceP2JPNbl16OmeNOlnl1pb7w1sp+QdEY3PcyrtvpGK9jdzOo9dp
TlBjfQ07xDkbMxP6Ruqh68D9oZ9bM5S1y7lw7UDv8tTsBSvlKVFJXt9CJcUl68b0U/0nzVA8muio
/1kDRYy45KBpM/GC5aoG34eIUhFPre1juq5WCe65G6Syh+1PTUMV3jPCZZZCiVsJbaD96L3GzO89
RtGVRrigWXTQK4SP6ooe4aKnj3b9qo5f/8UsOFu6u9Sd2lsxUt5KiRNnfT8HvcBJuc9SgVEgfjPP
khMAEnwWRqwleNYqedoidrhJu+4BfLUGRROP5TbQT3PffI+yRCViou68Y0W9Eh4gerOzBtale1lZ
NNCbdQbn4prFei5KLRQ2hTI6gYOhYPz6eq1Pjo3lzbyAkvatL69TYwIbfZYDGVcePVlLrG2HQoHk
O6C6Bd2+lLwAli4WE/wtye5yXmezKNV4L9j9ZjGAuHFG4za8q6H9XhzABm+dQ6IEp1CccY8ecqWG
d9lhy9R5qS5/1YWRqjTNQn0232l4CytTVIBTBpEcT6LJF2GNUkbLZcDcFozrzIjCD3TASfY3MDAJ
GW/fscV4YBFzUxMZGaWQBsI9z7XerF+EJYtXclwsX6N7IKto/TtJ9Ch9g/3bjuKcm4R3VF/HWeEX
M48TeneslJaTnsL3EOnVKbmxqU5usvyXHnbF1SmY2hnCcMeSXU/hloHhB9gm9P85LYTj9ugFORWL
peRA1XVNOnVtSH2Uk3I7TeAvyviw9d1+P5XIhydC1lj+Q86sQYMLCzHhUuE2jz+RhbRLqUvXGCvr
7yjqX2gnCCzZKUeAwNz4q06uVgplZYcQSG63ufV06AMN++3jr/D+1b5G+G70tBCu9M3SrMN07Qpe
FIYDuMPt6d01YA9V250dJiQ6zOrRQzinuhD0jHFsdxPNgWvLyDHRO3ddnSYLATRdseA98HUkenZ1
Ao3SqsKCn5w6k5tNc6GYPjmfcRVgrUjDFSKWBXBlLf1Tt9z4mfjPvqvgxi21jeuCOoQnXO5sawkv
T078PMmdf03aKyC1aerzwiKMhuZH7jSiFGq6cgCEbbJ/60lhC1eClVMbHD+TYwrFXABce/PzaDdC
jJND+YFz3oPPyvS6BJ4W/V84a+c/oxXDOPwj2AmPbItBuHXbI3e40IPgI//AkiCRy2Qz/TPLbuX/
Z97cKceViodUEe9lkYOD3xjCEIK6jFnz+bexY6TiRG+ZXc0CeT3d7BmSgPfbfm/uWERA6qfdSMgi
ej86PXqTNq6RoSkYRE4sSYFnhcdZPjrSd1ntAQ/b+xM2E/anZ09TeWjksfL0sAmWacKkf+9n0bEp
iJHo6tBKgakt+fHqn+//USltWVqH7pJZVU9TlGLYUb7vXEAHiDnAbuFcwKRvr3rZs0o/6EBFrETh
XIIlz1xVuPNWHTvwG7Dj+h8DYcc4m3Kd7iG00+Yi+89a3wbhrSdcl977Dx//ow/7E0nY5NhGtSYb
pw2dcYtxYc1AfwMH8VB8Vp6JHKNIcWbVVpgjo1cAdEmF9nT8YghCQv1YsQwBxAFXvy62G6hRQgk0
X9CfzzWHAeM8eev9SUMDAbOMr1bcuuCROwU198o/IAvR1a2o5dE5KLz7cluR/o+CGa6xxTwk1gKG
1efwQHppR84dUaWjRGI/PbJnVwUJD9vme3bTTT+4KmdApUDp3Y625GwZWTdP3+wt3kK+UpsAAPhY
HdS7EhhSSIw8slTd1dVF/RNwuthS3sEE4ZuitOeNlik0VA5mYwfcq63gkZ8MP5Lu9nlx2jfzcSdN
pXQlEWbsNjzKDH9LqWrMcIUQMCxdNLDPhW2zmgzQeQbqYqAr/lO+tFgJJdUkNvdvT8ehz6jIuLML
37iMc7Rz+bUMwLmxX63VtlKACqGAc+Nfr5LLDQhbrS9B+BhSMMlhVSkpg1zl+5dWpUlGT2YlheLN
RZZb/WOWc7esdOE+iOWl/Ogci3Qy4IQz1PCOpxhGM6O26PQn4Mh3OH7pqEu9c/WLsa2/XuomdeK2
xlNAQWSkKW9bKN+mnK6Yu5JpfEmiRnB7yTmkCDj3K0vWeh9TSQFahffcn1zSW1coydajrCzgP2nF
i85UrGn2S4f+vRpG9PJvO/Gtl5yfjJJDQGtlMCTyyWWAi59D48L7Q8jhJh4vH/B5YqGs1CLNlq8P
pFjuA/9jDzZdiQv1cqi/UEJHqCt1PmxYfoLtcPpw1KYbOZGwR/J4Yn6POB+iPArtI75pL5P0bgh+
NcOy+mO6ElY42SQaBigri1Ts1g9w2lQavPHdqKfCEx/mTUp5t/pGOVbhK4ou827DJ3ofpqKvJZSx
4TNpZNvCpJG8i9lU9iBgk0/u630JRB8+35dZ0xz+g0VqiOPfTzaBpCVPfhIxULw7sHJ9juqMYUs5
4kZIjRo+9YWMHXFynNMTCZ4M51wh6XhYJEmT/hfi06nSZh0QqOqlhPcsmVJHtxEtFh56B2UrgB2/
a6GO6fLGJT8UV9frxU12SNSTy/LuRsvNkyzn9tEX2gzrdX0nDKV2dxNnulDvu4+wu1f0TKp0KqMM
KEAQOUsJyss/lYn4AVdtoJ5a9yBDDZlfnYvLBQz6/Rlso9uxxVAgcMyl2y7Zo9KtnSLZU7WlrFA4
9FhLomoVXDxqZuvqI9xNSwg0PGMeeexheDfdzQKCRR5ri610N9Z32pSNKZoDejaFgUn3JfdurkVB
wUekqLE9VjVGpBgo+v9jgFoeLp0Dw/CR8eDaSswi3CfvAyMoFxClJbyupG46oirNGZGUxpFwLHCy
6E+v7obGsc8HdkMliGW6xt3zyL7Cisr6gWLZB/JZ2rRrYq+stby1yIh/gjDKR1qeBrcMwJNTNTPz
N+jOFC4DLzSQ1PbioEP41AZkDNNYSvH8svA3m4xErJJLI3EqW+MPspuLw7gWXBW0igBtZGz2+d3/
ne37wvX8d9A0vsZTPYKGDcjwdQkpWwTssNbK2G6qJHnODj7/dX02LfEnAIW57x5Zg53kpgxLmOgs
wAgJ3jQAjU5QlIlgGQCsovo/3ixF0y4k6VhJw3Ned8wAbmOCUGtVUpmiFQ0ZPP02Sh0EARW68fVf
IK5bOoynoSuR8R2/p2XiqVrlzQ/3vgtRKf/d9Vdn3iHcpF9wdH30g6U4DeU51tFBXfuZ3k5iEcIF
nE3DDVTG8+A1OPjKCKVwlBmt2wc/Pkc6cBfK4UTABpXnZGX+PXBtwG0qnj9GNpw36PRoVhYJ1QDA
zV+tqc/qf3b5B33EwGtv9W/Vqgr1bhlupQ5gJdgWNdUeqKHe2L/fesxkW+fTBJzR531CgpnQ+X0e
sz6deY1e7TheGbI7Ixm+LKe7itb7P8tqavBpN5AlppMGIKeBS9cfSn8+n62EsU4gBTsXEK2RaJTu
N9ZJMlhaKmF7tlBn1xYo4u3YRJOqIPXdAqhFQ7el21PoDA1p8V7u7ANeBJQjuvTSUTn5PS/9dRE3
NuYs9iMVDKegDlQRAiQlF3djixakCkpf7CTugRgIUi4GYiwO7akFmS+cJdO9VfaVntfYmqg7hWKT
at/7iKpvNDmhYJ38UbMTUX7xa3ZRDASuFvpk0sQp8awsPKnSH/HErtqCOX/DIjQPfuQ2IooRGLkC
KX8DHxxeuuENpIsfWQ/AwYF21SCJjaF/DEi8z653syIK1z2d+fRAy2thpv28kujKkT1DMUlBSGqY
i8H1QO/Ct4Of5gQVpaV1KGuIerahLUIBrhaP6VuH5K1inEfadTXwvFsmRwbmw5dvtKZA0LIzKQ0P
sRMgEC+ijcGQdM3PNyl/MAUrHwBEiKelVINOVIl9MYzXZjhv3Xu+/rwh4geJqhDx04XoSDDP0Yz1
1GGXClPpelES0RqvnjJNHvP6RECvSqFmDYytEBVdMUSZM9OQf/SEvvNBZBCuYWLLj30he2T8kUjO
JEIf3jU1tgE+x+VyG90Zm+vz09rsgQlfBG3P072x6r7yv0xZIzRZp3P1EVNVA1VrD8PaRS7w0dqM
K0y2JPY6uhwI366MlumfKJu5Zis4n4lK+KbeCx+rAoDQnots9WaYEX2cBMJ61GzvAXxfMVqYgOIx
J4UF+lUL74/ZK909i6J/FVhRhMycqwhB2//Je+mzjleMBW+eyXJ6FENz1S1r8yqWiwhsmM/Js/B/
XMVwJBO8/K0oAqVfoQU8ABzzBgb/SoO+JaXL3sUiSYjxpUWamul/V8jNos2w3WUltM+SeOtJhfhJ
+P8pAlO/PwfKTHXthP7tLQT9ZHtiWAvFlRR9QLxinmTQHYM8ZON3Du0B+jKdejZCIl08+Gx+cKpd
wDSyw6Q1xnZLwdgGSyeQ4DoI+0WfjOq4lnKOQAXUg0L9bIHLFOUkPl3o+pJQtf+w5WiwK7DxQrw4
uVznj5+WvzwS+rI2JNTQWWcJsLn7jNO1ggGDOuyj+d8T4eJ0vBJFvS9qlWClczU/MGM6PLHcnhR6
8+aIz2gd+UDgthihBS1+/6h6mI68WeyMeVZZeQAKvcfGYbopny+fE+UG8Wjl6SW3ElX86CspLjXW
l547OrGIZZdxmrt4+Qmz/SvkAXxZb2aRajuH/0aoMFkRmLyhdfL03eryzLobCVkyynuCFWGyQES0
QqQcAIXCmY+3ttmrl8NxFyvSWj5v/rKYV1O4JjK6UPcT0YVs8vUykAUVuMaJwwc9ee4LB7Tf5VKd
evWb5i33KW8xD0uTpAXjyQsWSBo7wf3aD9dkUAoEgrbcX3EIaIFsik4zinhp+vSX2pz87w/jxgny
ME0PwWqCDAXlfQLQsqf/rdk3NaVr30/G6XJGfBLCMV9Qas81y88+53s8/gnM7K9Q9Cc1JEPFVIz+
NvFMIb/vALTgJsAZbXI8GY5iLV7PFTK51N/hk9m5Gj30X0cWVVVakTzHZZvoefulYYcNW2tRt/k1
E9DmCBz9NL0dDMRPIsOjthJQenwd2fZvGAuj4kTMnsb5zORMUFq8EQlzcBIazDqXxnPd93Dd+Tfu
Z1jCh8/EarrHAIPKvSe/RxAo+OtrJpbuRyobkYsnGNiP2cofMGMMBRORBR3stb73G/95EDMjliID
ijBYAWiV5LnghIJkxATBEXOWDebK9aIcCvLP3x4Z47Dzj8bQFIVf0MMiOVUZYIe5WU28XfBc/I2L
Y1pOJpgSjQ3bHFXfig8eMj1BiOPZiVbCdu+wBKbeY/MHkwtdKfUiWOJMGz8Ilqhx0+HirE3rxcQC
lwyfW9/11UBkyzAvKYhp3hz6wqbr1iAJ3lqfMNYJFdf40u2/j8pms10QrDjEScHHcKDf3LjDnegz
Wd4xzeJedSvJivPkQtz43Tj+899nM4cZgRDZv1VbXX+v4HFkIWwF3J/oGuZUt7B84hLwocEj+7Dt
j5cXfypEktjNXXB2SAlpyfBQFQUYkk3ElyMQolIU1v82nbyn/8XnuQzmS/UqQPg/ZSoNWuH0DJer
Xi/jXN/DklaGXl8KHTQZa3Jaxgy968MWzODSNWOnvLUPUs7/3owMTa+4D7iV70CIMuEqr6Lk3Dl7
r3KGMQclyZQQ/0cH8LyiamMchQe3J0k4noBsXAB7RgxouupHAvLhbzryk4C5TVdB1iRKFZA/Zws1
FxW98LkWNHTIynYa1mo1LUHsM8DETmtGo9vUCiWBV+BC/DJCZJtNiZ9kbS4FjlGKbRNBw6AsueYJ
wLk/axr1Pws0hZXzY8YP7RhurER6U/fg4m3nmCi8jU2vUbRCExoAfvsb9Cnzd+g9cUJvJFkTwf2q
tqpkj2KXxx1/5BItuXCak70Z5Stwqgxk03H0lBSVoan04tKQIYxBI7SEziANkenn0ZXMgAimvkCp
n294T5Rb55Q/vGovXix8n/p4JmWyMJBGKZtZF+aF9N42PWtHwEZZutY4OO4IAzBrb1HyFhNBM9tH
MhQTEj6HV2IUPikBuJO/h4c+MW1eresZkzyV/ZwymcxgVMK4jtpC/hRrkKXb6j/2ZLlHk9CopyME
lzb5N1JCgYTuu7s6LxVOrAkA/l91fiQDH7nl15CK3TcmUHIcqbV+rRn/oTMB3bzfJnHr5AbSoAzw
5YQ5V8/rCKME8RuyXnSsQQysQRfatnYIJDo7HjPJU0DAH7KOua68VXjktOUvaiGPXDd7A27WOf9e
dVL4p6ouAOGPv7bBWL9vJjKMYBQXj1ZGZA8IwI0HyeRiHH4b2ONGqHGoZbwk3R9tUeS/Q6TQvR2E
TnhBcTF4hq17XjQuB3BkscL23Y4rcuecsHR1HslVmoty+vAfHJv++faobQX2KbwwydpJ8hCQOXdE
bxmuUkrkZ4r1RgMQt+FoxZDi0d2Om1qxF7OYEb3hGRoAd3Prop0F4l+WCXDvRC+KgF7Ghd4EXM18
dbW/cke+1JhGXJx/17Q5HyKuK9mLQLEbrkGJUsmXUIS9UqG2XkABcTkoXXd2TAHTVeKfYsmgX2UX
Lra6f2rouiU1/m10fHDe0sQUNHCyNCm4EYEmjDjQrX84p/sox/wyHisqHAU+HIyGb0ePex1+F1FU
Xf3iOCfiFSoNqwd05EVbYi2qdX7YiqyGAfZBwWWduSjnZ/o/TTIiAUWNBQ++YUnvdPOGCXGjfK9Y
4CUbVcGkBneLTxDndnzd7UuGp5ybWJgjJrMwiVO2DSB84YC6OxjFnrlRw6+7fPWhvF+MKQILUGRq
+6Pp7f5bYzyrNimoXRG4cq3heI9FKkBb4TN7lJTvlDbJriTDd6KNXOiacdx/tXZdRlB1mBFXsPqc
7VbiW14wg/DzxLfXNR6Ru3xlQxxJWwV6GpPXmZqtsg1ig3d5RVjoIYKVZ20TaZXIDkhPPEDbWnBj
jyQKuWddtwUzD2smc4RRSWWDQWELERivwmBKDYrHHNAW3SILPqlQLqC/FtK8NHuv/mbx6aI8wd79
z093XwrUI1QYuKcDMDHuyBNnvp6kB6/nfmSQKD3n8B3r7xi8+pK2OjVE9bTvbsS685mm7PG/nYh4
8wpA8gDV48Nam2f4KE0lEB/SuCFaKFo2/zQKu8u2egDcw4Yn4eWvgqzW/LDzNDmwN+RDYqCYn8ct
o7TmtiCXI+6owzq7zFPYSH/VQVZ5zmsUcAozkoIIKUkLQOfRXId6H+GPOaxAxZJZJ7ZkhFAxoIpx
YaYwviYVdPTJNjZ/9UyFqxNKQyeNXyVYVEgyGZRN8xtxsJGxh0n63r/A3M+vjgEh13WvSXKCu52O
BcEIZV5CPosxAAsuI9/zwD55+kuwm0C/uS3fR9nQlQFc+ZX3XhAKsYzs11BgSoCTB79myIAXmbiR
1SpVAZmOInHf6eqLSHKaXMHpbZebrNV0CibJhVjmq+EFZJDHR+ftiLaf4//vQz/tgBlRZn5TfUN9
HnqNvQ8y/55MJgGQxg9IMvxCNUnE2oVKqw4v/SLxGnDoGyaA+vpn5ELW2DAaAJ8m7dg6IphihfAX
DLOvplvdDw4gw9/kqr5X13oUvHa5HKKkG66XuYXen5QgQkkAkqI8M/+uksrXHpFWKa4/nbPQ0KU8
MCYo7ZtfRswqzsBRer/3hhF0vYLIPdnNHVIFmRRKso1dnVuVZjKKU5B3csxNWV8hL1NlQ/kqBKok
rqusudM+s9qfZt0D+ItgRgpuJUu9EoYGkQ/sRmp1VYs3cOCXb53c0P4QC3izD/FPUnHT9/ypKNgU
jazYC8CtArq3ML5aGSJQuBcdQc9OVXnesB7XGWELTVR+e0a/xVwdeBC1wWv/TZ7SdE1M1TqNHK1d
pkJ9IaLifAU5Q1iLDHTMpAeNoMzB3ISpex52kosqx0RnTcoP/SHTV0X0/xSimP2URUksZtyCpiPq
gEx6O5y0+XrORzSXDh7Lj9AjTSWD+k8X4df2ZYmGvY35A7OrddxF3A//+YS6zMbcp/U6KMUi9wlZ
a8ljpBy6imb0ANoMEBySEuPRpYaBgKSwRL2Rbl0gqdp9ScB9fVEch8im4zefLro9xkWdKwInEaVZ
CUHoLD7UUsPVJIxH8/lNKmG6uw0trSu706T1n2EcDaJguCNB+1Vp8E/jLYA++NcjYipXprFbGqCW
+DZhXDimEPc8IKvH5bEmstdH6QJRB7mEOGrkwPcclH3FkuOQy4p7zSgdfYYWfFPxz5IV66oQLfxX
HNKO77l1CEpwqn7ipe2on0E9QMkNTJUbbhCnTJUVjXRTmnGAM9nKznaR+4QT9MjWMFCH09nxNLox
CRm+Eff4YzLPIY8nijjvmKQWe4umcANfAX71pca+NoeSyV5YsF6aZFkuoWYwwit3wi+gAiItx/1j
y7X3PoeQCHI+2t2wz0ArNopAuv4iyh/JnjKB6JYUcwcHa9KT5QuCpHpk0qpzz+gZW1JDxBePBPpI
at8f5o2RFv6hu7r8DWFVURspe/xvnupLVpvknoWHnDDh2Wnl2tI0SDPq/srZwlwFPV3iGikbfnMr
sqP7yqiO+QPbuHnjtZhZx5XH5Z3MXwwLg3tJz7F4Wa2SLJ8Ec+itnlh3RZ1ljVRlQsRk7A7bJWgE
onDuw5AOkjvI3WvaZgclp1FAESZzZ92UnIKKuj687mYYGEfyOigatyAERcK7W1joW7NnEQ6r+iSr
BGzFUy+MA6eTB6HL9DpX5KZxAq7OW+vMoM83csbWc04e0Z46ZX4jdsq+He883dqFQB4qGW5K8IrB
DRRTnRp5Ap0WY2UkDgzmExemqf68Nya9rUd2nYg75NoHepEl8zwORl9Ez36Zlc+jNUyod0S2SY2W
hW/QCwxcGuxVCGmyRaLd3XaoCSpdR0e/XvDBRfl0Ewh2nlkMCoqW9xn0U+X7Wlwh+rejTqPairwg
anIuXG1YUdvYFlZjaZvzvRr0LTb0Uyl0jh7uYbJQ3nJaKhUaW4XaV/DLmDPKdnmyXiZDUJ/bgluX
IE3GBJJ0G/xytDVCgALtPplAWJ4tmeh6vhXhvuj3oRGQVw2Wr1aorVmDBnZ6qYrr4hkFZa8shXlL
nte3bKbV7YPaODDeiA7YYrkUtAVahH+00qQVg+H5f4XWMiwhS6hbr1txsl1hNMWdEGV+asxTFMHJ
LNyqJ0l25tAgrNFMS2C9mfR0h6JOfSW4Df04tuW/PZaH1VQ0ivjw97ivUoqYsNvFCrR+X2+GAulD
YU5IxYXosU0moN0xXkHjxKwjxW9cGu0O3sJrwSrcz3PKQJ97x2dfLb46GaaWyg3XfJ17fyiArM2r
MiNW6tT2DkxgPZ7vEdTf0ICDs6eYM2eTYfe7wHda2OEtaCyLoLNmFf1E6mnEwTvW0QN1WWXcbWbc
b4w9fuo8zIoycnH4UVpjyrsaCMiNcEO43SQS4y+DnQ1bsU+DoW+kyWUrmPPIP+xOdsnf6GlhK3UB
OpeKhaz5FnBKWHo1sqBjoKTATdE195IwiWhIsAWPahJ2SmEZs1Ckcudf/qHY2+aQWI0Es224CuiL
nfiYFdXFRKuZn5oPb2tyIVC84nIY3r62KpB+c0JDNhU0g+VM/X73QVSXczHuAecYyd3WFgLcfpnE
IxO+BeRtsPMU3UQYYhVKprjtMuoeN5nQUSR+eHuBxAL1nFP4B1q4ctdVX7536dLiXGfElWQ9qwjp
sW5qKqoXmnoQfpO28IqoPrFATreppWP+4GAzT6edkw3+kKvCg1Df79jW8RTydwATyobQutjE2497
SzGD5lScFXeDXHtwIM4zUZBu6si78iZwSzkIboGA31lbGmLhvxUgCoQNI7pVHjyVG70o+lE0nWtO
icM3pc3/mkCnlDEx2+6WGvt53mZOYx+wNz92/wE/Cf0GChMdpu45qO97/P+1VUvVK9c8+PzGtH39
wGQTFJONkEYMUS0gavYg5gUZfQtAORjrJ+7QLGZUDwt3Qe60RgjqxEpPGyNSA5JiUX5h0ytOS01Z
bqcTBatHJOZvL+ArTkBVFbCw0VeW7yrZoe6GVTK+9kHd9XfgmCywLsaiURyBPRqx6YJpYLFBpx55
lpmM21jVRq9WwpU1ZBjO0Hv2mqssF12veMKQ37xOVKpZhx9CS74Op4o9vFTRX0XUHEBekHo8oXIS
u2e5tlYBVwLq0x8vHYc09zUHGkzDU0SRaURG7UnnaY98nK5EgD+a7hy424riVc2WIjSLX+9cJa+4
7gKd4eMF85yYFEp7+i6o7sxZHihZGJr2ItOLnSwtrVnbWyaYdel0YLevUMwIertofMTy9GhfK6N/
l2uWU6iN15AFXuP5sJEkbUG9/1d5KaZZOdcBa7SKLgjrPEgVZzLrtPftGC32iXODnV3nNK0cwG9O
t0rb8G1UP0HrfIa0wt7NeAZ0tYJVo+TdPkfl+7e6NxqALXjtgoYlZxRQZv/FHR0NLJre3gE2dHIU
ELJmGzPSORGpTSLayLNkALAlERtN5zN5gFFR9nentqj4KEELQoXWPiPQKbVLLR7/JrtCTYRh7a9W
Ne6m6INmjY6XkGcm/tSeg4MVr5wP3MsAT4Trdru3jwlRv3aM5NtZQ/Kw95UK/ttaf6+dICh65znH
Yz9ZMT067AjbQwpZmkC+W4U75vPya7zXaNe/ZcCn6bg9/xZQ8Y8oxwhKEjWHFEMRm4WIFA8YNaXR
/zWIGwyAhI4tvVItJnSyoHMJ15dUWXWn6thnj22omewyUMOaC44PFIyiu+9SJh+Ty8r7hBeJzciL
WVlMKiNBHhkAIZcUgnI0idnxXS76LUzwmpNfij1O+RyhaGtMsfjoGYZTqzXq8J6swmVZBa4CRqic
1EcQ3iIB/fTcQ3zKJa3fVi4gNhjt5zQD8Vv6uDALpZsJkfCF82Y2whF3OjjQWqX/Mee0n/wNe8eJ
IORgnk4S25cjVm+ksPQCX6cEuDr8lV0/GVhR2hnKHGIqf445Vl8mQwYUjZ6CadiAVGqZVwxccEGe
amo1MGxnC/n81MUtwPR/EqLTjg40UyBOh9Id2IFn7zNrGzzqOyrHLlnnzbdCiIEAGYIBjE+zIvzg
JbMb20cep9+B3WcBcb396cJH4G/m+TPjkWEqK4Spi6MvorlE1nq7lXAKrieZAQDR4KU4RDbetAN4
kLY26gas2HIT9PqQKbG50A7dLeK3lh7/EtQcq2RUjpS//0bDiJRxlpvc1kjTIuFZsPv9R7d80kPq
X4rKQH3BzxfAgKW09sCGGFnwjbFnlTeq+tT0ll73inz8tlDqAa73tqrN8ywmVvDn/doGkgJL35EV
MC8I0iR/P5FwthE/D2ldwr1uqsAQRc0EE4B8Ka1WmXRaDjNiByG8qVgM204ObniQZLpJ5BHeSdaZ
ParAoNuMiDDpBQQDkIdH/C5bTwbSw223I4RqAvV5+yVDNwCW013lVcmA7QTuxJ0o3cPZb89lzqBc
NbUxUJisIE0/yL/ZKu3wK+oSrkd9NuBpTtp92fWgxtJmGxXc2QvGj/lADh8opOa/oVEcelRFMgMf
2D4G/YWjqOrJSXlouPru/7d4bs7OrERtZk8yyDifRd5HeMLELP9WqCfGaUuLf+9QGq6q76Sv4NVX
oBcnDeiXNnF7jAN8bdyKZGjvtObLpmfHyLGrKY2icTYuSGNFk+Sgj8Ehs0GuQWfqigj+NPWERxVv
g3CHY9TZyMNE5P4iQPVuOTwUzq0UBbV1ajVI/4Ryzq+3fdp7N/pc7T1wJrUVJF9D1ZHAJBZLsVuV
wDxv2300kkVdO3bpB7tfLzQGmkmLEdS/LzBi5/n4Ldy8EM5qQ7rGjJDb1H3R65dY1oh3Ic+WhX4F
9wODcmqMMFO3FmoQcVf0tlli3rbHNFFCQXCrTBvvMaNO85i4cdm8BQnZnN/BkInqov3wamSjVkkl
S3V7FVjsGFdtX7To+tkxF4zjlqhi29Nnejsfdr1IJTon2zxRsIeRCUGLptU7jkAMv2Klho2a7qj/
dw0ZLjtUJl7bW21TWn7LMyY4Wp2+j1W9iMjs8Dd7+P9ovYXtJwKW/dhBDfjYlXRP4ZRWyJ0aLjwQ
3+j5KbJdnAC/o5ie3r8qgSgZxIg6zF0SWd963o/qp+79JFV/bb/unP6nU3W29PbDBdv7PT04MXwQ
mvIOs5OSM9NkWfE3c5VbGqvAtLNXmC4p8hGn9I0rtAq2KHKZsjYl+DW2PAO4QlWKGUB7FtHsOxHu
H9qCsswTS6MIgmWXhIMcHSbzNlg9TBdwWb2fTH7WAPzgqhqsepfPo3st9qlhXolwkOVlbgXrdBdt
506eSFr45VuVt2Po05hh7X9sH8yTbgZWNvbn5wFIRSYwCPRM2tJLwA4szclbgpnf49a27IFF6GeF
/C6BzxYLBBhpoKK9K4dbdBpaLe5zp8eGpjsmce1lCz/E37EvsatVglJeiJ+fNAPARtc7al44ROTg
XLQiAzuGEacRMRmySsle+lLjThgQqQcOmzM4lcMf8Q0W1oeWX1ExeuXbZIiVptamf3g/nV6wkXUY
ZUF+BIqU7fiGlMkoofTymWRnBMOcj0OPcz+/PJlVFssAmEfh5v5mO3ra6stutHByrvWLlY10MrHN
zrRMqflFwzniRutt1FM/x66FgQ3EpWdjmrg3m30SmacGXL4zzS6CIO4niHPm8MQ0TzHihELHL0Gg
E7DDUGbCSdQWm9zPHuQWqxQp35TtRftwyGgUIs1ita4bV4X55JtR/PiD8NGbi1lHeKw3cAjt9UCB
rPHeQ0IL38GjtUqQhjjNl5d0hRrnS9nZGfuaZPp9gr17NFHR7K5QnjiMw7g3RX8hW+6cECLU/3Pk
A9QvR6aC9R5qOw7t/bgqqLKqfmdU+eXNReGumWLzRcZy9b0+XqcOmxr+butxOxKNKOZTmrRvGwCg
jq9d1+fH6U9uYQeyeovkJpJTbmU2qPmavkxS6VHHhag4GDvxgqeLgfjRXyD6/j813yLiTn4IaPpV
Plm4hA6afgt/pVY5/UIxp8U1jHidqYODMfadqdDqGlLIuG90WpgoVWLS1e5+tEVpZ2DFu7/5+Z0F
bBEnFNxoYS2BtvIAyQju5Ve2jwr1AUzPGotllV2iKw/ewMTZlKNf+OzljTYSOePc9P1GCF0GH+PL
FEQGYn3vC6hRl0S229bKiDngi0NB0ls5GCkwIhv11I2bH/pl5kGNjnqrsRukWpSMkRzFAcwp+L8/
phFJkuaO6RaRQ2zpKYIAG07IzUIiWUt2v5PGibz1klF0v2P9sgqvQnEzStFnppZsqJw9I7F6SZmw
SVrYw1W7TRiSzN4HYgWwvNXyLo2NAur4113S95VeWuVXVRm55Tj9xay7yoXnrjIlXc8pEr7SwcWX
TOCq3gPsaFYNn+lhwTCPgkRFIWqsnWzN9UU9Os0U3Lq9E2/wLtAJyho/CstzK2LE5RbEs2dS/ns0
fkei5o0Ggcv76um5T2wXA4CNSGxWkp3aqto01QfKYQ/5Hs+Cnxljr3ZRX/bMzIxzoiiUkR/BRabV
IZ/VI46B90QtOlcMfFMP+QZPlmsAdJxaFlrKzUgFoqTkUp0WGk74RVwm/XuJFVtJmzrmgbf4Lwlv
XO/kjWB/seEWojgMig3rl+08SpGZ9uOnqjnjZh1HxfUVLyPAoKZDgUHqnmNid1P4PKkouNC27S1K
yMUZSASTPAPpfG/ROdKKOEG9oUtcP15mQ+2E+bIo+ZSzPdo1vO86rc9C5KlqrNOoMG0VyhRGo+wp
W8YTQ7Y7g7qkD3S0yBE68VR4Yioyfz4yJgUlo7ZG7SoOWtz6oM8MnqS9Jt6CYo/Ve4vrO6LXkH4/
Rz2YsSoQRAYf3lX6HEuwAh6sW9sFcqlB3qpMzmty6siD1DvMNtrKq9IhvrkL9gEPCfFTAIgNiN51
eMbEtFeii8uSEOaNsqt7VnP5qxwrR4RNinKcz9Innyj1t4E0t8K+/xwf66B5jLxXEktoSM4ZW1vA
SCzR09E1YtvZORxl78JkooJmIhRXZCYEr1KsN928ehMASatK7pZmcJfW6+cgzCFUpji03ii+L4TI
JeTyLo0xBvlPzaN5OqLoqGHy19H5142+IdppxpO1prz2H2CZFAWRwUWA61sONeF/KYXEmkSzRRP6
w2m+kRCBTxd3oheRKl4kEWnXac0ViOaVwfRsLkTVggSuUkxWao8PwUW2AdFoMVijKoMrC5HYqfqa
o5Jy8OIQV1w/lZqrgz2OYVgdjEE7wtAofdGeNDyh7g5Oz2qYw8GjNcKZWjeKt2EAizQOcWi10HNK
DLUifimj74Ti5cYsCXN1WJ535X5pW2VTINp2nICIhej/PHuPja9ZFfTtFtNx5PbOHFU1t0jCgCpM
KOZQh26irIJcNFhsFDALks84BTiJ4JrB34ZYT1+iUO+KVuVNb9E3WtFuGW1kITJY+QqMIqZgJvSz
exF6zqsBG1Zc78fB05GhJGCGLcTf3QHcYZE27QLyOrZ0PtlsiDUhmTktKAkrm6BN6wlgrr35Zldv
3Iuko1ixSBtt6bfChbxEwox3o88V1sMWgelJ/ke8S3l8M7RGCOkwhnYc9ShZgpOXmxM4H6uvuTrc
xxCU0uU6ekGcLZQFv0nC43cWqPlXy5xig2w0ONJHZ2gbMBoGHGIK8khXBKXv5eWYbJz7HXfw4dZL
60aTDYR3A9ykC+kRzL9Sou5Bs69hHujlgfUG8RZlBg+CYK7X1Zas0DbpXBiMVezc4RALUoYRhxan
ndlj1zrqjNdNP2WMH/JUsvR15dZN7K7O3TKw6JvauCZsNwQsVJclo4xhAJfRpFNesU+TSpnXePyy
IJ2JUUkK4TtELeaO2B362cLJCjq5qpgQt6Ptv15lGenLsV+IwYSPnMpR1ZL5vIGt5SgGiAn3AUeb
4qHnoYmj2GPRzHl4WWq0Kc32kufrNK1XQ0LfFITR6SlqdS4HmbWS0ckPKRXc4fRbLWXz6n49bGNy
CxyfDF564q6mthZJSkbZwQw3yjKyFvpBo6lliq9zB87RIaTLElcVu97nAMNMYtNZ1Fvs0TPS+JSe
SI6RqYRtw7vbGOFfVw+DQWZsrpywWtmifJK5vnqDvsIk1gh7ExUrgdLsAoH72dO8GnxgaoongAhD
eDrtcAWTASjvqQNwFQXLe6XhBKn6zwgWr3w0wygZktfCjNwVrc0uuqO+eJ56pAy1GJSxVz4bvtLv
rslRbue7qEd8HoOz85NM0fVfope2akVVPuuzgz3H6bhWquorsoMXl1NjP4vw89uiJK0xDrlpAzTH
nKeJi1adzp9ok8k8oMU0arH7xEaWDntuVCirh7dxYcZgoRV7saMgjjSC5iN+kCONiTFZhzCZdwg/
7WwJavns++M9rlaD6YzYySG15m2AOoVgEmvD44zJ+9MsUzoBdq854XPMKN+CVV4vqBdGPwyC35JB
xQW0uRT18lnpli9OKug3g/0HsUwPh93EZlhLq4Uc5EgTGggdZwex8FITa8sUFKH+dexda/qIiymS
Z4QQy72hVWIP2XOyXkK6ZAP4fv/H1pNc1QK6hMbrcupFcP6FMV1kBJ53LfdPw82gknJFqdTrzoxr
51rdLXhysrjJbnQeUc/snGNS08rmdZeLJSPesho0qBlMWFbMyauFT3wxPiJbnoo+h+kHCinxd3T9
ypkVwuyz5E9qy02CAuLjfFZ6qwKGMxuE3HIv+ldYimTnZtrOC7mNHnNLBHOtc5GnO/5XqabvuFU+
BxpU+05GS25hoizkH25x3PW7PXfwanYqijc2QjZegl7HELmJESTuRJ545TvmESAJXy0JaYGAP53G
UuXpogxtbOZ87Jsk/E0rvvPpQkyjDdaqviLxE1gQXJvJCedCpluchR+Q7iLeMsIoHcvla+9nFBAP
3eBj7A7nrXF+A/ebkpKdOb6w9bzWYLwUGG4dUjmRX1uKaPFeaaJYWhmiNoBEu6Hnxjj3l7hFtgAU
JeT1+AyC0QCeEWvn9QwNjzKEO2Gn9BHE+Zs/cO4stib22XiX0XLDZGbHh/eXHsgkV6lf3V5XHfsb
ZFYjXGiJHdn4TtHYK8nFyG9CbPAnKXwSz2BXy2bzA1F/aLTHL4bzHpdo7tMkeILhZVacHkKk7gAn
+Jcmyh6WkQKRSXS1mETF39b2lO5+akk0Rr5cjeERD8uqpKmCH8dDu559SfQn4zOJ8BZ6AmjNsXcq
4yGThLviRWGWGQyu93+aq5iwikBxcRAf6muGqDptcYIQgGKibf6SHkhssjeopAB3ga19CAbsaLUR
+0uZuFTImtXtcSMG2r0+DihNM/2XYhpC6AuH6Um5XyWO+rxTud1s70wruv0bb5qRxwwBSlAAaleV
QC2G/TQRNneoVhxycwxClun2keVCDyUnUm8DEiMdWqRqLDmLDApgteBgyMVulGYKK/RJYORdrYCj
rlyvrREARCG8fDkY8vcDLCH1XmZdiOtqn095HS9StW9Ya+xqBqyX2cilU+9iNf9d4Y74FWO7LqhS
CbZFOGvnW21l8uTgxNGjZvcEDv6lgEq5V3GkD5I65Ln7BzHuB/ex/+q9R3gZJgGRkCDzNj0DO1B7
Hxc5gGSSzLvA7QgyZLpamWvCINWwz4TbaziP2zVr0iGZpfdoUypwgkrOseg3dd1ca367zNW8W1SP
naLIr2/h9VUSFjK11i8i1sMRcW/Ietq4qE+DVlbwmUony4AS2lwcAOY45TBPeP3cQzdRk0jbcwiR
bbp7KOb8ukM4pcj7mzskKKpwHdU1xWPyz8b9LmVewBqa9XFQ7nTYAIP8SwcEug6BaNn2uXPnA0ba
hqZBtDRKsUEcwCu2XxDCsrhYH7/9ra3K7SJi0zas3AYghj18EHIZ+MlowzzbyeYa4KwnfQgVJ21U
hjJDrfH4vuGlHrkvZGfWMJspWsxAV5kWLRgXComnzmFI9GIxiUkGmUA/J8iYWQBqQx3N/mk0ymHk
pRfvEl2h01NyoOXPHP39HX+o1tm7bjyMeI21Vcjpq+l7ibaE4J3ppbai4rx6DylvhDq+h1BTgDks
pTUQzxO/xFwK/R//vyTqQAhY1x/etNsfyCGfpL7NkRak6DSQFPZ/juyXVhph8Sl1ygC44K3jKfK0
FpG1Vs51SMeCYDAosV32qwn0zy7EL1C4s3M3ZzkQl1V+yFnb8pkz468vcdSdok5JGVPTUDnvhkdo
DAiF6GJM1lC26WvdNH4k38lah4VxBU/Z682CyDvx2EF6bH1E5i/Fc5KZJbAvPNN7zZY67DNXf5Se
gP8ASzu1ecysGrgS/iaAPRjyjHSAOToMrIVku+zC4bU34RMOYSZIumdvcEM2ghM39UIWQXOLOX/D
I9C6997OmYh+yaC2XiwWbIyciiWzcnZAKqkyrCRcxft2O/EnHh+zg9/ySO8dedah0EZbpQXZGy3X
OoqHHMqMGXy8zSElkN74cCMxg804B307LbcpT5lkqryui7PdQ6hV1wc8TrCIYnEbB4vq6kYyu8i7
yViRxTK3oX3sO6TeT0Rlp2WKRJftcVMY01ndbNHMOb0wPSuc8WjzIP81sJCfsjnY50swF/5U8xii
4BdIvY48AzTdKDCBtGOmhDIO+50WpyIa9WmUwziyM/A/BEMss8Msic2mTA6PnZTZ1UvBBmiGpzUx
iFTNaPK3KzfZ/xn1c96JkZYz8fiR/gjcxgm/Af/EvXr2ydBQiq5o8cmqXLIW9UC/2Wic3dnABerT
afSyofDMfbRwvJCX8HKTUKLe6kxdQF+2hBa37aIrvDej0i0S32ZDkoXaqwlfZcksv+wOXum2d9aN
O1tEJA5tKG1iuRyHT3KoieIx4ni3pYGWCNjsDUfDUpmL0TyrrT88KYSagJvdyuY+OF7GczBajb3J
7joxBDBaSaJ0t8nrWSxbTgJI5UVRos/THF2GtBy7i6DN3+/QZcdWgAVuvlNjOR6MEeNyXFTIcdtP
QFw2axai/zXunC1FKWGvWJEeSCtXFAi1GEmUhPho4vUT+ric0vuJ2Xo0AbaFOfLWrVV2qleNFMtl
BzXGPZkmu1IUA7FKln2xbRXi9XxmumU+m2WaLIV+CaKYNz6y7MYiGp5RN7XH/cboRNExW2bBAg92
urCzs1mGPdWYK9A0nWZEr/oYlJej7tBarAtsstVjIqEmCKhGCZrZdVyESWRzf6UZp001qTnDowoW
SDLa/zYVNSqp6tn6lBdX4N0kQPogbICjCzp25zkSwcDV8v7hEqwUk2JY8dDHqoEC2Lc1PkUbJ2FX
lzyDgR5QQxF+QBBRbiiUdZbMheyyjU7GgEjUbXGUFC10unSC5U6LAWQ7Y+6LzZnbEYMJ2axYoaR2
g2oQ8Y4z8FwmhB3AR856bYdG4NhxAqDmHD7m+wfHsgP3N/E+rc8oYTgpu+yJ03oq0YNm7Kz7geSS
6/YHNncf7nMb8DBFPX5RqhAJN1KKe7D1HHGYgSrX4aLyxOr74BlBiGR2anZx84m8ARe6EnCHPV19
bY5zKBmNnR9qQFnk4arFybSx9rkejgWolSZ38Wsfh00AwJIFyf+FXxgXHrONfIGed++2QxXx2O2/
o6pl+OYQv9u472dD2NSQ8CoZViTGgwdL3Jv60Nb2DUXbZkZ0CGc/24RbdWUSl6fewQoGhwHgD0fc
R+A9QWcmFW2d+3BcYiOUY403Qvgot1vszgzumqVK2+acb/rZiV6B8rje137TCEnd4gGSAR2Ylf8y
lGeuJS4czP26E+9P4xwgwgn+Vsw70Fi2swNRVwDyLUcmajdmIfUfy0y9bX6ljwMBZqg3NFLtisi8
8B6qIxVEg31ntIRvjfPnanpSECH33qtk0ZHmT+MKPoFJL9pXAr5ObAxMlYnofhPLRmasFCZeLDgZ
Ga/yWblG9BCQm55hGKxx23NGe6fCqB/xDdO+J3/lZMn/hTivN2gjAgR9QT+e0lkykpfUCxkgHK+f
gD2pWeV6eylq8XfzmI0C9KiolfmCEch1GSU4sbay6AOjhECmCaXxMYFEhvo7d84ilzRUh6mpDc+9
tL6uSQmpNii7Ia5k+D4pLIyvPGrsIAw/zjD3a5QpmXlsDAlxqfb4BpOPaVyyqY+zEvACXRZl1IZB
rvh8ORYOVFqeHNezTI7Jj1JaCqVBSTzlTetwEftOyXu3Tlmeh+4BUhYaUykAWwHqHFRX9AqwUQO2
jSf8M8ygLWtPaRo1s5chL+XzrC3xbiFGQkK+eznWY9ykdiJpQTNguFA+88/strLGjMX1nvYoad81
/fJr8JX1F6voVmMTKm4Sd0CzyTLZIc6lVeRp6eWSQdEKOu1elue+8UfHmgimJAkglhaT0qMz1AZT
4u2zzHev+sC5QgESaSrwj9bBteSQIraGADM/bdlYiSh4gdYRF6HbPfHvGRJQaQdKcuBBe3BwXvLC
nwSBtPxompCUdRNIHtHW9+cnZq2KKH0nQw+lF/2eX1XNr5MLA1UgqxuVFpfPMIDPKWbzLkhPqbk4
g9ZYLBuToZtNUCN+4ZRThKzR6HIufUnwksnrb9qvj7BlQ7mP3dQeMrwkfg3geA8XUYjhQGXuDsCn
PcxmQeW86JgIpn3LirowZUmpiCfsigOyehwFIaiBqIWdrC9k4WKo9rIhha0c4i15PRfkD653cNt8
I5yJwYXMfC8XfOk9OkrUpPXqJxudth85j3910vUFlish70DWbh0n6u4NZEgWgHU0Ae4JUi5TmvN3
MwuK3AfYETeISbwgQ5z2kjHfldNM2ZHDCMYZFFmD8dYbH4+93qbrz778uD/Hu3rL/+jmnfcZi9R8
WDJrGO7vs79GovHS391TiSihzfh+qDDcpxU0ZqTi9IUFutawszPODmLOhvQ3kZUueCPnYk1YkYlx
nSszQ3VRet+z5NMUJm7SZw/KM1zK7TFZUTlaRMYgrJ+Oqjqj0b7zmi3UxQrloZ2NvHiKL2+0JT+W
FB5ZaLhGAlW9T23sdO1yT/JHC5tj/rU6oNk/M8d1ZKBUFrxIudIlY73PFpbjRLfnnTtY2JsZl53w
SvWxQ8ujO/pv3kt+HFQKcCmY4ItwgbUppn43uo7wuTai6AbXLFBQ2cXO2XI4UKtWQfW24Uy8g/Io
Xy5XKWULsulq8JBNXDO811HwFobVSD62OI4VOk/k+Uvy6i3idZZligSFBcsiIjHWFBlwIMh0/N8s
eOlnNhSFz24akrs/VX8ofUK/aa0HsRRonD9KsVDDpwogkA6mnybehqP+llZIX0tc6YyqzmThuZys
sWWlXbJEE8P3WRORGATdfIAK5b/2LqJDTpU6rF2ch1Xatn2HoxO9cluGzAKak+YNXcD3/EuUyZcq
kn74cjhHsmvTuJE6IppuoPCSTodAJhWKWsdf4s6Jj1f1cEfT4p6FlXZ39nV2a73sKRGdJDwb/tlm
HJjYI1DKVt5ydUz8RCah6Wq8mck1YEmGCNSHCjWX0YjqtxaJcVXAcPlqyx5IxSGL4L+bPLmlCgho
NqTis3iLL8serPfSmxCRi/BlnLawYILphPhoqxaFyWTF4V7t+9ggDPj9+MpBlB9tL6z9WszYP8Ux
Z3YcppsrLdfIe1q12mAxBxwH8CUBr9VBnfzc1TpH42JjX9lXrroBloeA8PwfvnVLRXCo0odEwwNo
HjUpk3VDrj7812H+ehqiaatp7e6YfU/mw0Bee6E/INQxIZHaSqKKDTVmby8x359nyH1XTvqG25V7
MPB6atOunzKu1lRtAQcrSiworTBGYVTPhR5PMLtAq7tbmoGoyiuLjX87YitqpQu+u/Irmv/T0Wr1
a701nX3+j90TQ3pN8kCQI3Ok+6KpUekeJ8NeTFp2wG5meK5B+P+sE8iEbKFtlyUXJS8FHUgbZCVA
rQPCOdLZ6NruO8PQ9T3P9yh7RlcbBJLFqObK8vTWdE3v09hy3ZkBKvSjl6qhvVq1bLtOSIZATT1I
Q+KtDjf5/GjiDP5wSlA57odwnwpCm3ENQjQJu4hnFvqf54LGj60qg7BK5EOIdgQyPDrGu/6WJ2ow
TDttpinbt/l6VA+//C2k1xLe4+py1ar6UX0NlqjdFi4OiQmKr4u5qj0xbakv1kbYZBvL7ftzr5vm
uVxpClc4phn/fX84LzykVg+zpkRCSV+X/zWZmvtEQ1Cnx2K1xQGrl3jZ/Mbf/VQMIV+dbOOW8nf7
A7lAbjuivFZyrOFX6s4DjGv//1T2aNtAkB49NRBtJr9ECRuJj1gq5Qc2EMyuhkJRyL/5YiVzIAJj
+0WHOqkpKq9GLtBqi9N69ihoyUhsEXdT0oUxLlfzXJQori5FURVfiVmroUAnPWq7yHqrsFg5POaH
HYV8X8OSB2gnzs2o5612Jxwop95WDGDuQkEHX+JsS6H/0mHa0e2WUG+qlNMdH7NsQ/j2ItP4NXD0
9gcdopSq0qv7o+5pkRpkK9q7MLqQ2dlznnQaWTvbZyMCeRkGuHdR4yRHj7DjG4FSZGsWXhzXj/Df
gHb/o1S+jAmhGkXUgmhVhg+tzbozzjBaYvslFZBN+eZsQE+p/SUN6slK/NSKWjbhrXIjR4gBieru
OO0vwsO2LczOj0b56UbCjXHsUpMTjf1xrLzCd3ldlyIEGJQXf0oMKfjlaF/E3IqtjR9OE67NtCCj
WEY0QaGD7s7ElbypmwykJKGfcK31ipZHxDBedSSL6e3iDYBsWHG2Xqn20XWxf8CnPgRf7EiQFngC
KpOvjxxranwCBxvijs8WtbS7TrChf7rN9A5NHhfm6MsDcL75o1nYzBrCnEduooHFLaoOJZLxgxEW
ImVpV5OXsdPHd3rc8xkJXV6d8VV9O8T347COltP6vB5jxUL0YRJgGFma+DIIiYzz+53ofSi1cHoB
G6aS8sB4vNoIJAaHKWuk47zymwFI0nCNksRiOZA6hAQrLC3OXmmKi5669QUeCbJtV6ntBgCgYdr3
n9+YsmAAjStL36pq1ohMV9lHoIvcP6QIA8HVxd73x2S+fbx/rLT7xuibqvFwtRWt/PP3ZA+5bYze
ATZEItJSG9Tf2yISyDne6CG329awym+CC7rR5XV5qr5yHS/2DXrMf6b4HwtM3ww2exy4bxz+n+Hc
YAhhkdadfsXqqdbAzXEMUcNREDuMV7TZ9tPTDYk8d3gb3jGRchqRSY5uyE7rsL1cAhFAn/CoTafJ
PDISJ4v6FFGclA8w4t68eemNvUQRHvW0PS/EAfF5mlXUOwG0kMmII5ZbN7rzHcrOiILoXpJxWIX0
MTIRPnizGFjGEaFeoOkckioPXB8rZ8V1bODa62GmtJTtRQT8dZo083jAVjQfq8cpXscTg+2XODXD
zZxNdMjVNtt9eOVGWiP4FRZpAg9swV/whu0p+RETfXsiIsGuqdnfDTn9lpwEygYYYsKdY2NDkfNt
WDTAdzB9/DqSpKjnK/AKZKFbqGD7FkNPbMj2xGIO7K5zOMlHqxuNFOXmfWquV/71N/keoowMrECf
QE94m3Jl9YX3Wen8bSquwP56rEcuzFzrSsC48jpq0INZzJ2tRP3NoD4Biw4LrBxPDLAf2bKZrF4m
dweYv+HH0g91XtnIODLdY0SSTozhNjQW4ZNtqXF3SIhBeD03skjU8+GJiVSsuCGO2gtqGXHpC6Jf
bI0465p+xO6OeFetC1VMooITe8w8RJAcAdq23MjM5LKc8koNeFpA5Xsvb9ydK6MKxewcjCfw39Wz
8OwRln0HsSR/MNTJVGADctrDrhgitVXolRghp20Fs0Y/dF50skPVPdqVBSbsuhLbM0cXZMZjVXTh
SFp8HceHg8UjlV5zpJY20rndIZGf6EpK5QZOmfKMRsB4nJq695sqvq8k0DrWDcFY2f+1NXP32o5m
si/vxqy1+CLTtFwiQ8WyMXyGlRChrSz3uFmgxiLi5q/D2YzBpcqO37Pasee1qvvXJ4imqGiIOJtO
P0OygYnpQSzcCq6J4dfmOhQpxiB/umsRznkoYcKfzvZMDczSnC3usItWEhIxo38isbRMKCQnU47/
lL+b/46Rx5e28btTyqdv7Z9MP2ns5V4CjAl7oYzZLe+ycKeE9eCTyAADam4HLYE/zCN7ImwVgXvI
hgKeZL/qMzgsX2v6ToCmAE4zMZ4EzS00zdBlATOFocJK9DDOD80XYM6Ylrlwc3LWKNri9PUcCFVm
qX8uqPCa+lRYXg3NJS28QjOy4RsmgXQOI/NgvdbSHZXeOsnVM1ivgdqzK3B9Rqo8+CENRLVRFC8e
m3NMcA/PnXSn2XOy/4hpJ4vUUoQXBY6TDX0HIuRExM6JNbYdwGXsv66HSRVFidlrxEPDGDaAjwxC
Rq40mdID/9Of85AVRqv45zIO6DTQeI/okDK32rAzebnZiLGVWZ4iEaks3QbDNkr8a9LNLoSU3kbv
Rn2/KPKNqiuzbr2Xfaa7WI1pDAYiUS3O5sddSlZic+EPbI57HCl7+NYU2bYv1yYQ+3T7zrP2AXfp
l58W2dJaEYHpBqTq4IaN5TuxnWWZPIGShRtyw9c/a1tdP3MwaZTsggFXjVrHEcgIWhleRWFN8VwQ
vMIiuwynVHUVs3yE/cy/h5nfNAK7vR/7u4DySyS4o3Lkucz4JLFicngh3AjpSIGGgq2VaVdBDg0t
mwDB2gbBM32DXJseTTWT/U7+SnH6a20apk/9xz2SDQ1MEOi1yjWnVzaeuGEKpJcHWk9klsbHRxKf
ZrraiDuD1/KWbITdmdsYkJ/0jH+Spv0pjlGGm/8srbzcdAGEGwYBJ6DwUVDOrS9Meq7HUAeN86ls
aw+U6at1un6Ci9KYGsLFoCwidi3Xb5y2QcMzooKLdUMEUFykc864JtyE2dxocVP62aXyCse1f/Cq
cWyThN3SWsINqC2f/GgIVWw3qfuqgvVy93LW55JtC35W4H9mAZ4d4gI+EsqNiuZmv/5B8b2QzPlK
M4IzJ5tzG7t0ANIxi2jyLBjZI0/UCqmN4XiRgFnIXpgHQJ2CUIiELoI5CIC+svumpEYLyjRaWODp
AXv3oyS31cAtvPDbOpLD2Ctn5cqLK/DFhKGJMbNMbxZrQZ2GBTdMSWMfpfFtAicpN4dG09lPIoF8
5FXjilq5pABC0INLmrNziEYdxBvvpCukQP/OYcXyjKncZuAnJHtlxwYntw2mY8i7KdWiaNusVIdq
EdSYSB4Ht5YcDXx7u8vCQgdS5KTmofRAucmA4D+jCFVQ9cMZO1nPSWVNAvQ6yxPTsfK4fVj6fHNX
FvhiREN8QI2/ZwTYW6Bqwg2HXhr64ADXF+hHgf6iKH8YBBlbT5t2Fh/bOR+UX/X9ApqvZkPBrf0+
xhb89bcVCxyPDgS/7SGpGY9Cw3tFjl348WV2FQJv+3dT3o5Hgo80PuMWeqDgQWaVlpjKEITNA0yM
1/ERVEMMPwJQsA472CWRbQppLS5+QxEER/dEEdb0WnP3eYUILr7Rs6EYlXCoppqEEg/4G24BDIhV
nbs3hrIRrQJN2qFBxo1le3PeOQ5iCJZF8NUMeB4xS9GlBQnyTRFgxF2r5lb38SPNI68EAhyBq4PW
lSdF4SSNbv3hkehKFnMsxPF2GpKyDnFBhg82tPpWa2rNInhPAwdFwh54Pc+2WF5faXumE9lDylN0
4LCnJY2KgbIVnR+jL4ivfNkqq3YuNV1/jtn+7ZPn+KOiOR3GUBKa4pQLp607KwuqUD+tmyj0V9X+
8zaA9dasjeZXEB8F/69dN5XHVNQ8LwA1VVUQrhL1nr+8q8vnvrxgExAxV1SSuBqDWOFcWJsQmci0
be1QpUhmLTRpqP55HtLEKuYbfmCCb8NL6g0O/rS0QX3Bqmo0A4iGIxR0OosMmHFtT5sEVdqa39rb
BuQMbkpago+c9qrlqxUcoBP2MDV7FXeJMg/mGAh2/d8vcbQbsC3WU6W5t4SBt0qNb9106M+EQ4hl
TUgKHPKwcHMzvHcGsrX407KPyuQCTCYzP3vuz6RtL5rVbJsEjybSpzuGfVwCCO3tLWXvsDAZITkM
UJh3iMOULPMyn57Pzytk/fe0ltrr+B8e3h6oMp+g4AXuakHGx5ylppiBMQBlbVcWl9bIUgAQ9K+F
mi4fPI6HoGNP69IyUquykRUSqlVPbi0QdhLLF1h52YsvI5mUF6wCujqgygQ+i4kj2AAufgowWPmP
q+tuNzL7FWfOVhShQbWIoOb7P/yUu5A6vghzmtMFaaBPmO480hqVIrTIH006Qp5impeyzmMz0J6v
CYvgIHjeVTdTRFwF4eMl4g9In2pPQSGMPOm/80psPO71fhwWioe/1oBAKi/BjPkZ2MGBB1pGFmpT
I5K1Ub6PtozGQBuaFmSHbzGmG1WvvdG32CdN3zK51/kVUb4zbI5jQ9s2WwWkXbYrex6/1eLcRFHx
UrwwRijn3JFVtnWNkiRsw1B3DwluirgBz2h2HamWPjWKlwfHENJ3kurIuVRoQukyrd1F+ESdcxBf
k2xFZpLA840ZStOtPDTt+FARjxEjcqkrMeEO8zW1TAR4bfB05xZdq44OEa6tODYiesWTwvy6CnnW
kYp5X70ibYc+ww1soJkrwEa6LqaR7dWz1TEfMg8Sq7y27WMMs4UKpvHsKl9cJlynioOSomYatbEe
2pjTvHdVqpysiuVQgalCGEuEWQo0mDndwryTAvlVoPUW7QWlebbv/3qsuLsDZviaiUUVNLuYtxkS
aVlXyhM2sLBFOB6VrrMrTjjJ8iVJv96RboA91uRXEFwn6WsXYdnMJSO2AeFxByhQ6xmy3Dv0Rm2J
NIqnoEqjKhVg0LEZY3z20+6hbOJpEkgsvAv/zNyu8+2qzi4VCf58LXvAbPPWOZEZEnVBsjorzunZ
exVOeCVDfoiPrzjT83HFj0/KuKVHUXO3cFKQVzMZmleBE+pl3yMeMO73LB8Z8SpwA0g4mm8Bs0fb
p0+5P3r3CcqIFC/w/LbvZGd2QexqTFgazmihhfihwojHU7VjhOs4UMuKAZ9M0AuOwg0rojRiP3vi
TT0nvqvhzRgy9vVJfm8xgaUhUldgOWSGddIMB8JXEOwaaHOTlAmoRkqMX6bsU+f/nZtz2s4ISqDr
l42BoeXGkqrSsgBkOJ5+alRG+evlBU18sqBUXgY5vT3MhszUnYY1F2KGVF8lVJKfbNQGCfRtOUEo
fqAOqrBveaY1TQVMuRNBsM3oa44XxBaoz086DsVRpIo0vUgpzNjeOKXJxd6ZY7aYrtS4CoHBsgN5
Za53Tpl/Ud0R+392z75Hmu90VKV3GlbJtyYCUJxkvkLIbb9UP6hMBw0EG3VBtzKEGo8hPtAQb4Dc
YTydQeCHN2XhK2gxIe2OWLqWGVAxFp5Cprc/J5/AqWqb1GPtOgFTN/upYDZhrX87wljS6VXrAX+j
6ld9z3xvA+6KM2x6EpoIMMjnPkdm0cg0UxDmjCpG1g5jJ1I5cn2DmqXgo8FoBZ9DHTq1NHkCRQDE
VO0vJpbnAkvlscb/M6R/XRAjjmUcDdZiVrZlX+rWlpDKO2VlLSa5D5Xo1po13BwMb//l7q+a5aNN
CyM05fp1SxsD1udEPve/0XFsCTJFRzUJdHp6Bx8DjIbZh2z8j8n7NPOql3DQA8s9AWs0f1cAGuPP
rMFiVofSz7SSApOCHHxPet7ftl+IoIVn69qBZfs2E/qa2oNt4J5/IhAMRZGVL5pj75kcONpUv/Cq
KC7Pui5CqzTCLPyrQRlhkctL2wTPCV8C2ni+Se2j+W/zixZfYvTpD5n2r7MD5ZbYLl4cJro5f4WU
2ghr8Set7VttmcnpEeXkHS0K8HUFxITwptefCWrp0or0zl3fJiL7B2nORXZXiytaambjQ5V6p62U
Rxx05EtemfhGc1XItnWFwxJSL0EgY8oFU4jaeELoz8FAJY4zqr9CayklRuQM/uNQ6D58LJbL/scx
A2hmGnKEfghxvs1s6JRNYtAI3FmgZasVqiWYgDo9hHCMO4JdiFdEDqowVoyktdh6vqQEPKmEeMe6
/t62U64faog9s17+R7JsZJFg/s9YDc5XLeYpA31zOIVlbYyp8YgeOCALTBbrLuk//VpWFpE2oxVa
0bsrT73FUsG51kxm8ghbt+GB34b9QfzgZ2uJze86laIoaVW6rD5NypqGzvGm1OXXitY/fPzQGcww
IvLfwRt6iCFcnM7/YQzRnrizac/WjaY3Ro0OECA/EYcYjb0cuwaYDbdoOlvtdyg0tJLe2zu7GhVf
GKynPEZNHq1Eiw8S4fD6KCz+FYEHoywkq3M77QFfrWfgdblcwfNemgjlHYayEtwoPBseN1ZCIkYJ
KpQl/3nK0uLOPf9ea9sOc2cRSnyYdM2I1A4L8G84+yYuTNaMhLdnKNHQeGZh/yET3/X5UruqSA9f
VUSRRVtN7nzuxcCsaNN9Z7wcwBSCcVJ569seFjoFVX0Wn64r9cJebz+XQnd1xhqkVrh3K3quc+py
Ho3Q4VmL4YcR91kyvphYlaTf9ZbBsmaqtqlx8/g7Jd8LfLhVIevmMsP8UMncacJ3ZOZwzm1zlUHY
ml1tYF1PoxYwOlwGn1rdNq0Ys7LH2YoB/8MiwxL9YZc3u4DiABetXkYUWZRF1O2izhC4oOUTOknO
/iZAXgp3lPGsk+xCaR9Yk9TmXFs3rpjubMjRiIAFoum5f7ueWdRCPnzISXmkilXw6PdFSk7VCcQO
hFkf5uEGm4F9c8iQtbtRVKsGGJXqYw+uOBaF3yWQn3gb5FYKczdmWTyTCU2QYrZmjO1R3zytcfKz
koWx34490LY0K4sUr+0aWwCZoxgPZ+zT/TT0e/1AMDHSsDZaRCQw2n65kf9nhYYlMskIHnY3CKvx
UE5RQemM5V9NeyzSmsNHVE/ChDeTX0z47bW/yG9KtVXQv/Yrp15kPrRn5m0Zxb+UxXLiLKXJR+wb
mnvAaeldFGKi/fQ5lrL0jtwhDcBE9nB4g8+iJSTgDd6sm7dsQwjlfJFRFXNTq9uVf9SRIzhTRRI8
iTWTD9IJ24Ay+1HJ6RLmedUPqRoEIvvUCx1PPWff7PwmjUj9yfl735dlXoOfYRSJRUo037N1EFvj
9hbayDB1MNQDzqnAp410ZNd33NWrbElLPLS+5Ntv3ZAYkdLX6Ve+pzj6WXs861/qwNAaq9FAX68O
woM4shDqRMBEziwzw42b+btL8guCEZe1jZiioGotkVdmnqbIkIEiWmN/KKoR/Wiral4vXwEY4VrR
DcINy1E0EChP9P7XkL1Vj6MJMld89O2G0OOcGFGgJ61ZQXLQWbhF8roGdj48bMX8qPMLDVfjinME
2xM8NGBxBU2GDXx9X+IS0us3FN2b5EzeuCKwe1/D4BJDlWtv0tqUPg43I8zksfuXTK/W4pN/+cLW
LNZBxGqsRuM1GHowKr7YxWlxIFp1Grxf8wmfKe/461wCWinj35BYotEwhQbLBnAXf8T3JkS1irPL
heglrjvFwdxBDGoT5vX+DtT5zqfKKy17CncMm615RV510QXgsH4mxbvwiQplTx9njCeinsuBqPac
tfyoUjSrzS5qtslQX8YmuiU6/rvEHTd/zSy9dSqLOdPfjwhHt9sV1JKtOeNQFgIvbyho2LZwttXD
KryDrb4c8A3rcZZP3IXDE1cWz2qTpqZuyf6BwWrcvofb7QVqYZlteTzNJvWuOnhk8CMGdXb/Js/P
pqFJhfd4NBujK4CsZ/MlVwfc5/2ATlRYfa/PU9QD38wkadY8BF43F7Kfws1IjyFkwcwfoHkpQHew
XLrz8MffBOLRLmh5f0gR09m/rtQceZ26qRaqYVtXJkwy/uKdI6eF6vcnTp/DYoupbgbH+zSyv6f9
mAJ8ZOo79N0UCIFBQuTG5IjnGrq1/TqPoSAAWXHrsC93Sni3Y+XWMFyp3klrM3sQGIkjjpBj+R0d
78z/a2lY9I8RT9pSMJUN0EYYBJwk0u+af0BqBoSyA2I01KBOFW8xmQPnFxpKmbk++Khj8G4tbQ8q
hgFJ28AvmglJCZMVPrm/l93Irr1LjbykMgR76gEFVv5JVKnY2sNvoPEwl3OZKwXI0budr7X274D+
r9/36zCtC4btxHu2ZymKvvrzz8g5tMnrjiZNJS+Ujhji58u3hkJo8tOiIC1DlNvUdmThowdK2apc
9+guXSLtJu9MSHRlNvENxv0ALrKTBPp1HJ5mOzHSPfZ7y1D395P36hZR6aBOvB2JjGDQK1Vq3TG+
fHBxgkqT6x3XpGBDlbd3qeJcnwyZewRkgvCxi/7oPyX8T7mWmfJkTNlz/UzskXokKkVpBoV1OZ3h
ma+rGcULWwB1SEjZJ9f0XFlfwyTV1saJDyihyDGwmV/20yYM9tcKmpEVdI/N1Tg7EQmgCxebjsGf
DHUMkrFI4MEsXUasIILyoqChM9ZqXNUWY/EeB+lYrr/vIWARfDgk/ElU/Axaj+mULdsxNGihGGIR
NsBTjCjOEzPoKJuLPiqVpyceyoB/FTLuX6g+/mkmp0mKV0WX+5i6W/UMpibCBb10EWjo/sl98NDd
ip1Bo1gWpspj317ulcYupy511NhJki5fo14UUiKJNSDeWPSVeuF3z33VBqdWHMNzk3Qe0+Rrk4X+
ucmUd55tGa5SBs6088AuT5Acrd8MNvWk7XRrc28kEJC2awM1fs40lIQLm57SeY8ugrXI0srymzjF
+/4JRiKQ2meFFtxfeWAkQOYXDvA8Tz1sWSuSemcs15GKkGceFOxWozC9LMCjyh2bGm4b8HPMNrnM
OssEesXbP7/D/3eA379WRY6XilD8jbLyXyfXuhLEf4QIP9ZvK1ULTPtQ0hqhgLJ/OCjx+aNK8rdg
jhGW4Z3jdXxgEGXJX3ZnmAC+TsYaHd4AGRnFiOhw0TR6FbOvb0hOsubq+Z+pyReuZtnRVJ/becqz
DLwN2kADSBXotpmZg6FOOuqxCsAIGXETR6saBcSiWsquMJTuz26NecxMsIqexqCT0Ezm5miOdVOo
nSVu9GEEhkbO6j1TDwnsneF5MNO1Ohl+BayKaB0k1N/aJwjMazMVw3x6IsdUdcBEndFTjrSqcoSw
oG8jDglSIrZQpCnZ9NzLfPBE6hk14Z4Brq+2ae9+KkMnaxFks6DrJqkdUZ0oShp2ZmlcGQH5PWPk
fjlupy6KURvN6NessxKTgMSXkDgWMVOju3+0MZYw30480AMlk/K/Jo9YMW4fvmn6KlbYoD/QPrZL
T+FQYUtTiEct9cEfKjgOjX9lawaK9SNrb1kBSHHv8I0u5lSYIG668Sk6HRe9Ls6PiuecIcoycmZ9
e/6S8pv0IgQ4v+iC4pztwwg0K/gLuIphV5R7Kv+wWvTuH5x/mTh6TzT8tZYap3Frzh2bDsFVQ+DE
AjEa/FPKVvy5+TyBmnQ6HKhKBKyh1pPI5nPk009qyKnQ0G0vc0gOCtHaYWKzpO2/eXuSYwwz4/E4
WKErlLNfp88cqVoSDwlsygb/dkxeW6mNVq0ow6tIout7/kmzCDQ7HU4N5TtNmmh+5ibRSqkXwtJZ
dexl2xZdSGVEXnPASlzwSKKND0CJssqiGO53myRy/tvhvS4+IHosDiIoze8oLSHYu1bDl4bkVZ1i
DuClKZiT0ErQiLwpFzTQj4uuZnO72BmtjW74pgUUhU9O1EsV+1AQdm8N20vd7oQ2hSG0dMXdQX3M
L4nBVxGM8D+lMTAUQjhAPGNtcPZe7kzairI3Ml1b8dCcalbDgNR28MPqu5jvAoaTMJyYivRv3JMi
jV+xs1Bi8iYyEXQ7ulSF9Xv8tJgcaDqEXdvRpr5CNcdtAlWrQj3JGIvjIQ976Gtt7Wgv/KARbAw3
ie4Hy2ceBb9ZCQISQw0pqyZy11pCbZzC4ctRL4U/lTdoNVeeBCAE5xRTPInQ6nOwrpczu8OfVDu6
snrK5ntloTOEnmcP455Efb2Kt4XvvW0q0kSggToirM8C7ytCcG1k1H9ioEnTVHkOGZlOUXa1m9B4
BhlNeYdUMSqguPLTDr2LdSovt7c2Y0360SFJZDJ4tew0uJ3LljtCKqBwLXPGdnussey0ou14MHyB
TlAVtC62qn6eQq3QWn+Gy+nDZaOFLbFI1yunob0g2lYgOASWaCMLuffY134RhCvchSBlfDpey60m
vYTKJl0ZsHRZ78YlPbOjYmplkg25nzkhP2D6gVfavZ1s66pDcctLfzyZx39MftXnEB7HCweYnd7a
Z4XyghOKaCqtT0C8X530SGjOzYNQmYrqR3gzvN7ml8vjC1H3w34pWn9YFrZIZuHVhpOeB7LiNgkA
EK5YbPBNk7VeZ+xJZriqN/sNXeIznoo+QeURcOr0BmDKrNV5Rdvns0wdpRejIRDkmdMLXZHCKMfl
hMnPDoUE6K6drwEmVFq7n+keBPyCVUS4PR6Dc3g3vVwnTLvwzIKKmrY25i8pNaBYLRUvRrwjFZYW
hlyqRLMbrEEdeHcEXCe8RE3mNg2RSCh328xIc9NDVfTFhgqFk09GIqCvcHDcigJI2ZRnGzq4pRZN
ppKfFfo7a8uDYoFySCGqS0maIKZS/ZdAC7Kebzj91QGsK4ycySHNtbhlo6gBaarALHoaMKLr8VGQ
RXunugyzNQnrbpUuSTrQN29RcCyGYJ1aQb3frRkkC2bDDi6eSgC0B9qxOUJi3AUHgCLdbQzmktgE
Y9OyNoCVexhsEM4XFbnF6P4n+gSP7hy5/b4+qNVWJ4vEq0YCHzWloBCp0M88LFon6DMxLsaK3pS5
mO8hpdZpuhnPdoV/++jSeKQid3xWrazgI0BW9ll+V/UKGFiEyrY0N0tZvrIbnhw2xeAVFsZ3cJKd
e280MriGaqzX/mXF6hqIwpyWjnL3pp7VQvfeC4ffgkbzjyNlDCMqMCaezK7XzOHIRieLoml5xcKJ
jdgjYvH+WYhbLFgAMO9ALG1hdNPb82DKQDjDv843WjPT1k1rsL5lEs/V5azD3/gELxptQDvhdl/f
GzmV4Uj1rcLMlMP10pNrpyI2wre+WB2EYuxXMvQtdj8OagEaCFdt4Dx864EzoJOOoPVk9tcO9lGm
uxcOVxSRvNkccqD3LzaROdbHBqNQv/kMqg7WVmhk3GUPfHdygz0kn2Ez7qkV09l954AYP/Vo/mYl
QI2TmF1dth7UHgbtV5NxdHxmL+iB4nMmoiVLPmAZ8egBCWfH2NnUi24L+X+wbH5YbhAuZw61YpM/
Ac7GXs2NJsFYuoqpepX8RjL1VO/lI66swk7NCgR5v+LdH8B2PKnrYnlsyWEL5msKtky6cbcSfzCx
mTIi8gJPyC24dnggUByJkxtLkyleeBj2FHQx922TRN7LO8xxRStWsYt/l6ncYX+TYqAVo7twOFT/
ybmzFfvj2kRS1XsPOffgqQOqkD4KCQsZYoiuvk452tJvd80erWwfKYHvbwPNyYUpmfivzZa9J/mP
JzUTUSt0/QTyvPgr+Yo08MHjS3JPVLNmq+ATE4BU6waYiQKj4nZ4FKh2sotVmTwH63fGPCv2dSOj
nFKglGtVgeNUuTEsjuTLmyml0jMYwR4q/MJDbnMO5VEvXmVIzNBQMxie47GvkO1fWvREnxFS1wNf
OfmHnzpzYswBN3BYSFai9OEIrucRu419wZmkaxm3eMNUcGyDlRuL6nnixinuRiAWwcz+bbZFYg2g
AOb3+zpbs+lN6kobhXmvTjLcjuzSr2eEH1D+oevTIUsf/ogqO3aLwkcESaIYc1vIRRMtnIPRkLv8
x8TnkUpvzKeYqd/YU8Ab1tLYJYGdTWpucBs5M4G/fGQzhrMgXpiryUR4NTZdWaYi1PuveiGmhYxA
VIj3ehQbyuIaKLbSK7RMyMUJVT9+SrZ+1YOtPMBfmeMpCSKCXEecw21ULeO6kZqE4uj3aHVSIBAe
FFwg3gUhcFufxO/AAB8lly/6uBuxA5n+OvvoCuZnzlYpQt6ePZhu9H/qsd9FoySdADK1cpT7Sp0w
Ye0SrmMQ9oC4nsAy8kCtCEQnVi1Ely5E/zv2s+slDgyna8SgXod+UivDmNCdvF7pkxNWmydzBZC1
CQPWtKoLCmLRbLxC0qcle0Ztzc8tkSoSEtmD5VZVpdn55hZwigV6sR0TabUUDmnU1gXcHv9gtRUO
XhCqL+t8mgSG5N0Nsbkt5DuEEBp1Rz+3Znz3LK4F0iR9QB90wUkk9mF6BeDJFGfP3gg0CzaAiKxb
h6oqW8zOERwgYvmeDHHdCw6dBmkxIjXE6SevRvZ0+qrmeZHHo5o9n18qOMKhKhy3WSJcUpOwpWsP
wC662nNQjrKuenkEXj29c+Lc++SN27afk4Vn95FjJITrQa9J8NO4r5r1jovJU5GE6uj41vStJWRW
eNYxhzHS6aTve/JGylOTOjN+aVfIHiM04RWs/6g0WjQHq9HPDeS5XdbF68jhDl6R7IdmAyAt35JN
d0LpmSvWz9To3V+K9mYuvtjHZdAJ0zzf/t6eFYblIhEUvNIshY4kUtsGOKPySWQjLxy5USBie91x
o86SiqNey9gACOv+rkCS8zP3tqp9mEFcvqhJT7k4/gzTMGTZ4kaAnLvvB1ztIIDHJKx4LLZJ5RoM
nRp22nMFYoJ5La9CYGdmYVr815NTfmNaFWug+Mcd7SKTEnUR5eCW+4OuOHag87icEQfbMKKwNGmn
19Soij05gd2XcvHlKLdNyB0bjZvxECl3t9xFazhfmIVyZga3AMYM8WBvGM7tGzjGlMfeWryAaiLC
1nmdBTYgrFCYTANuW9yxMG4VpahHUITJvEXB3DRtpJWayYKwaMD5oMzsj94FmAplCkoKFvH6qJL4
siblqFak6plbZ/iH/NpJhZfx97UGDAFN5r6a7QTw47gSOvJTtPZVuuD2Uln9agxeQIyMRfjWu87S
ixiUryFVj9qjGJoBn4rpf25eY03pOKlsF3qtdy7g5x2hIfa0yY4Ns57gi81FRiIOXJ3qUUsU/QGK
Dy+rc2QQ6y2xi7nUXnjM+QCcg8fgwrXXBYmZ0oDc/7brher0RA3/RoXsifDKhApqCETyboGHGZYs
COidFiSDtiV1t6pZ2bSojBGYdk48iutveH0DLjp4MG17kmlcGLbmwotCHzybF7DYwuHqGN2pQQgP
krmGVgCJtYDDBBkUVlgUlwRr06fWdil48zJbO2puEBUMTlizHmOGhcu+gLEAZAX/R5lvS3lCtclC
6932LmsomQzCeK+QGpGyVPaQ5bUUM6i11Q3Oy7MBQcS9tDLXydBxAuxsHkoGX1B7g753dex4Amfn
JMkwJo/cgpSnL33tJ6GeKsOl58VXSbO+TRB1oWe1Zu07pgTCaPsHxMOok7fHS74AK1dO72pE1txT
2KwIUi5/mxv1BgcuslZIwJM6tbvlA53NIW3ejQ/4JDkldpDbrzFrTirbVolHYkVROy5nUE8BI36y
OYY6zBZk8xp6GZYCPTp4I3AlsVez0q9+LG5Digf4MAyOH6Wu+VN+Ob8UWhwBVJZLtJZbLhNixbYm
vZEEQrrbTNFUtx4GhFYSpg7eSncpvcSa90GTbvOaBpUp6BsWu90SvJdl6NcrJsSHjwo6JF6kmnpB
Pm5MwxMbEqpfngcm6B1WmOvTNcu2TOJO6ZbmpWQxG9IBptfEfPxwPvcGgtYLYfeOskLrochMbrXR
9FMCqjtsnagsPSpQahgk6hZ36mcIAx37kHqB8VK5M9bLWk0hKAuT+XGHlry3gw8wo5JUrtWGGZAZ
4S+2KQngIt5jVdCfnp6K/BEmB3Cg869/m6JTD2wU4FwVJ0zxXvhVKO7EkKDQ0kvYVlaNOrtj5lrd
fnuPxHjCPjK70JTPxgfQ4zAE7WeKeBT13nb8fjmmA1U1Btpb3vUSOVJD3kIjklfBJmVbJTIkFYGU
4WjJ3krg9YKXzlHDal1/1mA0JbrZIkgeTi1sOSk855LN1OWN0Qk6/AiYXdXEVrinGvCSieokuzK1
loRxOh2sJ0AURp3OjxxRhJWXBYxNhX8qKOMq1UgGa+dUJjPhijSMpGQCFTAiJE3Z03COnTkPs0bD
+6anCiEC1Mzb/9cAg4MqO7zHHJPh0BGASH4wDDFQZzlyxC+apDxnfPJNnliFjBGIZAFciztBoaWJ
u0jMUR8SuUZNu+9IKaTNht6mDQQ0iyVMa7RStdFiTPKwpggIkQE04qejOw3g/hBh1eQ0B9aOcHva
ZNEoUZjSyelHrnoEb4usaSJzQ4RhRgSpWia4TyRxyKx+EZ+UfeKVE8fnGoO5d95q7ggOd3fGt8uq
9TW0cGu+Z4ljVNtLju4LzYlcksuMyn/4ytqbzEEs5pxsn8y65xISa9FNEI2rPPXiZJxLusExduLM
wY///TLKTKKu9+cYqE7beLfWl2aWxuNwoLVFbTfjp8V4FVD674EcGwKI1YsXFglCCRAlKfGyRCE+
UfcBJZVzv6eyoYetYDPN9Xh9xz97+/FrLvBJZ8ujjnMriZUyA3VLgwf8JKgFMu+L7X6jBci8S2Ze
bLhPh5u/8FPp12KfhcMYMJuwf6CG7zGdduOi4KnP/7hbjLxwTj23FsS2SXk5EzBgcYtbHU+sk7fS
EZG7BfK3BdOoG/I9/dB4SbRjWN93ZJfQDkiSoS6UD+MXpotZ63I/78d7QBZ8Na/ZhkD/mbpj06WM
ZBddaxCm0v7kS2DA0B2Fp9/qiqD1gdV2I6sHeA+s5g/Zw7eYUDyIyH4Ek+9aiJwpzgcapKYI9vXG
EZAqJ4yV6G1N244o3QhpwK83FUUsYa6GqO5ialzbUUTlBc7cYqU+vo50j4Punmz2vOyGVsLabfqA
94b16x4mvRCYppEskph6pbsg3AwoSGqUopWd4c38Q1P1pfYuJ65T2TlRhRoOdpNzuuhY0OP6VowF
M90AAf0ShVRZuuFlRVoki+WDSbd4yR+spxrJWQ+J/KhFScw5LkQct5XkDkxoPl0a2Yu/ii7JE1Go
GnGgIZD4G45+HxywQaBIJMp+ODuxjxNmZnH84+T1MZ4eSEdS8i5CWBpGETH9vHAIflNKbJ38VrPh
WfPNIFcntY/c9oWOTLj3Zl/29aa9m0PGNDcpUV7CpxU3QEnoUJ43Lw4C1xDqfWSdkM6mUpO20mJm
lR7Up/kUCbdhy7I1cu9U28X6+VORLSxvlZD/rB41Q24hq0kuqEnfuncW2CkyYTFXt5wl071DaZ4K
jMPbTb8LRDpCBARjITslf115E55hmAFolFYmgsxSJvqXarlB/8oF4ecSETJkUYOW8a7qpA2XOws1
Ch9g5astx8zWcaMDg/JegUYySZoPQBySkiTOvsKfCK0f2olwh0cDHyZG05JQLDqKHXQrcYuOpWp3
cS+oww11Brv/wMWuyp4mKzuFPlT115RFJs9IuI7iAI35d1Yth8ZiiM2SzH7XzRBjlzIrOAo3p3XD
SNyhmos9reQ5WgWOAkGwSv6fW8Wt43eFKxsIXZE3RHvMsIFO/ddYle5MUqHgiVT9Ii4IAFpfURbN
HtY0MPQKlvgE8+H/MX+xjyFuKWjrC+kCkHkGPpwwSaAjmFY78cny8qKl7B644bSurM01sM8nGIFM
eMGqcV3MBA+poXrhEeC2oYHqMNU40R4wLc3sDBJfy3cf7OqQ0f5nXllkxuwvdw9YUiJMzeOEcVNz
c77EQiyZm6MfBJ5cYGaeATZLHL6j07cNjMWuxyCfFTYl/a1aCEIywrk1Jd0adT0Z06J+aA+ZUy1O
dSc7eL9IE5LGTRTLVdCR69NOp0UtGKpotJubP9ZgeAzMqHcNle3tPtsFtXHTjwDFB55xU37nSe+4
bYXMiltn2FcAkMOmuuSFLObx9Vcjz6YBGvc1JdEMDdNZ6mJdSHApRpXnmZgZuUldRd1tJPsNt3l5
G+LIXVHoP/m+/gsrhc4SmmbA+EFBp8h0gdA7Y/7CvxeCBp1PsNsPYlIaVxBbQZFdM8sxm/Ohtmdi
gjTSVDCmvVSx1JTOZoXN+Ce1LaBLPKd0oik5W30eI5ytiZXHWC4nU8J94LzfjDEf6QmuT6yneSWk
B0YDmSeF4wfVKX4rBg6Q/BCP7LlrRdOuxx4YYzgM4WMptpkOMpH5RGnA43vxrV7K3xgaC+8xuFnF
C2TvSSQ+AkJ++NXkc51AtMzY9YvvfIfVaGBI1T8BsM3TnZS1f5mg30NkPBSPNVuPyS3n1jC6LQS0
yqBeA369cpOTP0J3pRurASXfECC0f0UGew0dSX+TOyx4wWBJ75doy3liOmOLtgYte9kZ12cSCRrv
O9ks/PQ3EDe17fP9J/5VvFQj2jTspbEoW4gyXwUFlagKI/6+lbWnTXD2wSFuKt0BPemeXoRKtLJ2
KNRwqpLMr/fRY7IfMlTD84lbljcJ+YUZjZSzyUexnjIbs3+2lXMm62T8gvVre2Yu9EU+vtGopoqY
ZpHvPg4v5emIcm6KHH2bwu4MD+ctCWnbO/aA7rSVI+U7rqfGFMdOytLNkA+iZ8GZMYUM8+lw+0Hc
OheCgCFZbPlLvKUmukZvZ0XDeJs/KT2V6t4HX5cWp7py960BXLOJ/M4+WtS9D4mpbWwDWUikSqmj
xk/4kky/S5twXrv8OX0W2dZCDtc+qGqkE3Q6wJbPoNJMe/2J+mDTnqUSkUq9gjcvz8KyWDkPLezc
TaTTKviik9+wV8esiQww/DqaC5G4UuM4nqTxUP15oSJJgmeywZk/NJisMR+CTMzh0FF6bFutS7Ys
H41tG9a3jLECajxjU2V9uIuUzdVXnStWE/GmUeVOG9ZXJjNLaApWceeMSEv8wCzOT6aYNU64hw4c
Myn1uTR4pxpUsjZpCLABt4Fpi2cT01O8QDkOXUpVhzWlBho88x4pxsaHhrdGCW9UbKs9gAfjIwUy
6g2c/mLNuvQXEXhKqdyKROGmB73Gwv4pDCJukAmjSo3tfrFAUXcKmPIjJ4P45/XMoTuVuZPYTXyX
COt4jsTLGjqPy9ZwnU+VuDceaAO7MZj+rfWOEYuABDKbWbxDv1/Wbdqr/UeGEIuq38gLPkC3wLfw
8PIVUnNBluRCFmACvCEp6KEaBcHnptMcc7NzdAioQL3ynsY5Xo+VFWGGamP9v4P39Ayt+ASgBqrg
tnF2SKFL7jrRrMkgXztUoKuvTF4A0MbH8fxSNdx2HIWo6gQmHRT8FlQvU0s3v1bd4qdWK5MP/88Y
fOo2C0CXQX9kXPCb25A6Vk61fNAPsyNcFhzCWa1+j8lbRz01+A6TbILd4RGMqBRW3tquKSk836n2
BaUcRs1Vb7I69LXilTZzlAyZH1gfXVkYhhc2vP4d+0T7Hk2QUt/wAOTlIbgHcd7f0sV5VDo4A7cN
iM9nGWjo+/gGXl/cUavAUfAFJGw2PgQseW4S0AqOA3xx3tFddbxEaKNx/XIcxWLiZnlqD9A+ME2B
D9c9e8s2XeKGAY2MchsOfi0/k1juxtONpa14Mw7JcO5PWT/mKKkSkeIhLzuf1xhsFv9WPlbK5TE6
7zqxo3SqF8lJfY4ofCcfZcMfgS2pFjnBMCm6EuQPD6LqcoALnJgWS3k6KAlNusz/I//tP9EyhbJQ
jp9aqXk8y5Pri9Qzop0t18H/3lrlcQ6jc/idZ8ZT9e7dPioQZIBb0ZGdUU7j/VAar82Vv51hheUM
FKcwqebyCHF4Z8Zu4AbSB0QoP+5ZMgY/V6ti7A/1C+Hi5l6vDLxdmjSyNJ6KjASY1PaAwtvenZ6P
MztdvleAIylxykYNzXrfsq6uNocwNxoi6Xu1huATjj8w422QS/oraFu1ZVbBjP9FcG4bGz65Vrzw
ZEp35wqiFtjf22Ha+Q3AIqqyfMs+gP12VjwfNZ/g7fwMXnG6LF1W0pAnNpVuGVFoPP/rm1Ur+Prd
jHPOp8h52JSXmBJHJfy4PaHWXzcAKfha8ZpUJ/zSv8wIk+MfSGpAyRqYnoI2UbYboFu5naxhV/z1
N5oOaZJE7ZIaG2uhi9HoFHs8GbCCE5r2sH6MGF0/aXBwAemN5xfPcnBCeij43inhRPwklUsQRWhd
8f/thf5jmyJX6c4CdpJcAfZXcMhzFUm4UCBGsyK2OcXSu7hkaHb8tbPZ5NWDW/9BZ2TirJuufW1Y
ivr2Kn8DBRhY14zFrTueSHN2M8EO1VzC2VKjxgo/C3OeQ4tgbw5AkbXu8bPEZxIxGzUUinrfD1wK
km6RmgIn7jdrU/admLfRx6vZqOOjYHaIWCCsuL7v8M62C5mimX2KNMDfoRWlY6GMKibje+fvW/AJ
fPvzpPC4FBwciTRnr0mBS4QYElbESN6g1L4I8/HaI8X7BiNu/jZHlmGqlP1sWwr2ccLM1DFLilxG
b0v3mJ3zmPTsCrybIpBhmQpqCKpfa+CDSEsE6DqaGpr54i4DMBBK/LLmb++yFQmvQWHiJndO3wbr
QQou/CNzOaZkngotGCaf5BKaqda/2y8jfSFGNsERjOf2NPV9kvKdPU2fxH98ugGwsozc4SwioPCv
dHuL+VwVsiF+EKn9HdOEmMevTkofSy4FkWXpwWb2cnEBxy0agqNT2cTTpWlM35cJNfVOS2sBPNXU
mSCIaJ4lL2JnqPRO4jQoXtW6IafDJ0YlEF+LQeYQbw2AuXuxAFMwpE2bJNaW47ETfy2UWLcqxPaG
8uspt/sIQGbe3pHMG7AwBF4dHJIZM1i+JBDMyUvTIJlcPIDyzpnmkI/sjIT4/IVtOzIsgzQs9rh+
RV9qJfp9n+Pynoyap+RBS3/ZZPjsUwaytu9ER18VV+BpI2kAKcJVYX2D/rTjYPQKT2nJJWjtS+0I
Mtrj8UN2T2m082s01bqUSBuHOtY0RVG2HgwN+t2acLsX6YHpb5xhMoQXf/pOMknNthdYoyYQYDbO
PMeR5zf917gak7zQxNsijJHE60RglW+3T81UYI/OWxCX5XA5DIIfG4Mmp/SG1cRNyu0QeY+s6Wnf
1FdknT4lQp4NCna0C/wbvZbYNOy+sT7uafTi1LIzBOgPCGkX2AXC0mfvuz7FC6v6pI8jdQ7tgOku
XGFXpHljaalkP1SbibGai2OsEahYXLelSSJQaw/xFoJCJlFZqnL0+CP1vD9M7JNWkZXUSCgEvyVy
4uk75Icwkq7cbNOrF1ZzexE6ZSDNgxYJcGsYJ56OmCmpupLf0W3yT/ihtd9Wt23hM9CfTcSe2eW+
7NtIGjVG8svNKsxblbD7D7DxzN2VchZ8S4ljVEHlUWJ4nru9hEb7PLJmp5Ng/YnM/KEt/LTm82Rd
keyny2ZPBkUCzVAjpVWxzImKJlpLLSFakL6xwEiOw5fpHBwXSUKQk/l1P0OGqTu/I29gAWu8YdCq
X/EQI4TLqHUDoLah1h8yl6XzKubbvH6Fsg5LrUT63NWn5WnZCJr6Iksu9q/C0CpYrmIwCpfvEIcv
WJNrwy7n19EJz07SlbezEG4ncRVxEuSOuTK2HU4s5SjEAguW4MA8J0Er2hlB54jegSFCU+HJACfT
8/VrFC1wmar7JkzFM0q4nSDEXAidfhmWMlvaghdv+6ReOgVF5FcJSEL7kfUyOFGoCtzB+TvUKsKd
CaW5nibDcCU4pdkfOT3h9DYaP58HxJECnW7GXGbp7VIv/OX0G1DgvRngOwhqORQ2cn79ZHKtw46e
noSDMA9xsvzwFbH8fgk4PdpGK5KaY29+mzCw3yGb6ChI+ZGZUSkseJq/low/K9gDJPs+IKxOczcO
gGR4QGLqXY0K67HYJFE3Ok0/Xu5rRrLntetxOIZZ5Kn1/3OMxC9sFafOqqsNODuMRDci1zyDwkc9
v9QTzkZervlmrD2QOlHHWiUO/J8vBaIXb3cjCwADCFEwQ61TGcZ+MptqVdj6E4cGMpqsjbJ5OOx+
MKXxgImSwsy1BaxSbADzLb2U0eLWzdZuz3K1K5OKk8K7XzYmXKuG33lR9pXYZL0FpteAu1gigi8t
BhrPxxMPXCtUN9Ziubk7As239CqR67TjxR/runQhPGmrmfpWtTww2UfzpUSC4Bd145m5U+uFdD7x
cZEW6BvIGEy+FW9PLldrmH+165usik51G6dC1b71nLWqe4x1TlWYPFqQdq4wCcH7l1LEA4C4AjFG
dzS8yvc7PBXj0wGNh6Ae/cRA/b+MDTzmQwKAK6qPI1Zj0C+0F09xHANTk3OjIEHCznFmJIFoZGMa
NuDjHIdQ5GDbabdV1JrHWoMsmGhW84kwb4ZVkyrzG0k5GNMtaSZp+iP1NIisSGkMOZaFxRz+O2I2
QXFUr3zOaanIeCaQwFOlQn7YHbTqFzPlkP3qDW/GrIOU2hpE7KlL5k7w8vmk8MWpG+nCFjtfQxYM
C4HhZjQvxvwqA8Gkaq0jh5MuWXgDAcBoaibU9oRvsi5b6Vp9RIWcvjv6R0N0kikheqsFFYDiPZ8g
zqGChqdMP3jVcbdbRvs4a77P5zIS3CA8xg4Jj5caHEb6jWdnwqmMrpGpQrvr6/pva4wlA6JxX+VO
x50pGYB0C6TNhiiV6wekAlAbN15QgwDvnDRQfxHq4soOlUR/AjLTNv/vIuBBBYstrf4JP89cgwr5
DWnbV4MGqFdCA9WvhEtJurzoSUGemFogq3F22HZ9qHaIrlGCQzqw5k0b5e4CQ8MyDuMzOQSqe6gq
0wnckYnRqiydo28v4y3ST+soKjttUlqzrv2QyV5JO9taw1kyjC40X11DwVwR2S6ySsVLXBEnpeAC
jyAjOZpLBPxtxsw3OIoLy6Kq3Pc2noUOx68yLJZ7YUxM1NTsdF+UGXIsbRC/YMtHyg4pev/ZkoUI
HInagsefxA92vaomYJRZMW0zI+xjBxHl9WhrJeJGyvndVkUmm26asUZan8TOnuJt9ui41OlhC2X1
lrlLaECCV2NHuemuhJqVjGaBhkgWtYE0i6yRxWB6weCeVQRElipanvIw3t2yvM53FCWMIW8N8O3O
7Q5SKzy0cflNgPgiZi+vyDfZ86uV0E4G+XgDHZArzhOBcar06+/KosyuQWI1HSTMMBJVjO5FoHHw
ss1KR7UZY16Ne4OaEqk7uobZ5mvaOF/fpmKoB7OHGVq7wNIFKIDpyzXAj6fUbpHPgKw/tvG0SN3y
7ejcdt+qKx+yFqauVt+MPrfiEk3WwLZDT59BHXbUzMIKQFf+FuHjox7yZm30dtLvIf53s4RsuykI
vsb/bM+TSIEv6MG5/kDM+bDb9jgs3/gKUyO0A1lSUAUQUuuP6/HIe5UtWtqjOnmBF4Rka5JwXZCP
LvT8/M9ewNYoxH9VS7wEoj02C9AJ1SSrMa25lIj72EjXfRywiChJSflgxtSYFRjZDhpcqeFONtAr
1gI0sBTm0/r/R63RNsyL9xkRtvsestvVter642LubGhwV0bMaH94rZwxaqaZqMciR5KXfKBTkx3R
8+F+fzgn8OTxkV3vayUs4LMkN+9fliJlexa3k4XPrbRNSVOS+S28Tk6aT1R+Zi5Znw98D27fyaAp
ECAKzwa6KD/LOJul8JcVIRuz9UuxDy3ceLunx2IZBludpILeIVXwS/6z16dWagZt5xzTCJbVn37m
9CVt08mDdvYrxPXEWf/EiTlBUOeHrA+A7Cs78Fg87SO+AzIahi8JGzR/NmbY82Nh9IoTKVGTdLfh
1hgPRsUIMk98frR9pTa7SvK5U39x6KBc0h1fnAMo0D71GJAeQztXLi4jL832h+4FjVPs4kcUYGrv
3Iyh/VbsH/L0l0ZSjSPh0nbkgO40eFEkB5BUCqkAs/ouj5Fp5Yhr7qZDCLzu1AKZSBgh8TFSWxyx
Upu0NTh5eEffGDa4eYBVGMEynh8iMEQKl/accnCzIYx8Gifa0olNU+V2rXG7UudbxNMk2dDwBEIe
3D8ah9vrVQvh5yVBK8QN0vk8EYogNki1ZghAjdPLjDqcgoVJGNzbP8tPi90unG4Km7VBVhW3fQ/F
m8BJ7s2vLcmao+kGF3/gbL8e6HnzS15n1sQzyhEzkXcBRoGvJdTHvOWSYXZDYfpzJZkyrql793bT
k2Hk2eVE92RR+e8XtBhUfUZz+w1HC9UORGF041adsBrq/C1+7xm6QJN/Xs0qWnHtr3qcwyOPtPKR
DWdqUlVCqKLcqNpB/P0o4IOY2GfLj3ILtouhQgKmMJrJY8lB/IS6Xm5X9yKx0nALZSMZqklzFiOU
ihMYjHkkkbEpQJq6vT9jj/4XRgyqh5kFEX8pR5Bc6rUQ3UnJZviUvRVPId9h+b4TpM1a0gR5Ku+d
8OpY1u72HT3uDgSHQbR9Lxkuthx7wNORWe29Frka4AYrBu06St9AMzndRKDZAq28VaF388nW0nVX
6JKwYSVjJWvATeaen5H6upWe0LTp+G1/DoZ+W0Bn5r/WIsLHrZuUyFbG1VepdKQOlfCVD4naKOKm
gjj+HDNSr2hOgO8EMVPencvNqr+oAW/9Swc6HXBkql3lo0Z6G6AenUTPzi+x+0c9gFpx3aAYsxL4
pTP+59svE2tZV5rRjbfi6qMupfHFXl8J73YHLdEOJZjTTNJNTnmQcSFRRJm46rzEMKCYEq+Kw+j2
bpYdeq/QeLbP9Hqmr+pR8FsvwHn9mKUrDv/BCLUMZAD9wIIE6nF4+6ukCV2HodXa/jxB8dAWRJ/g
FCjz+6cEKFtbfKGOYjIr5cp6Hc2eEEnmmRlGUrxZZtM2CrthomEo4w2w4b1XlHhdbbDlUgE7An3I
zeKhmKkChGhIOdPBN43uY3vsSWnIjr+qhqm+UOn7O19XbEdJFhaHIpksWh0tQuw+DUhwlJ1WBpT9
rMmGlCgWcoiD15eRjWgoKv3gLlRsbZcGvYyRPtoSrQj2h6tlvmxXLNR7ZNWcr2R8it7r5KcM1Onn
BoNrt9DgQxi4+jTTp+qysnUaoYJuaU/mL/glhHMWiSPZp33Hctwd7TnBY3G+EJdMcgOAVK/EDzCu
3asIRq8WRzVzsCT9r7K26ZOpkfhMp3gl5iLgBDT+F7wNl4xoMB/zEJBP4TGOMRzxvFLSLwgalzbQ
sWcHVx3kfRzLjvQxP02J4IsV0w9yebgSF6FWToN30/dUNnQgAjWhLk7YIUwz+8vcaYjstZyjJfFn
j9WSG1qiZQFUuCd0NZkfIU4tWRsuEMvM2iYJweM4qQ4OGvW5TQEtOu+laO7JaiaGfLjrD1DygRIA
lCdyzQIbSMxBLqj2JxlGLZ3akFeuOfxE5E+xOH8GcaqrELKmVk/Z9YNrUAQfQyMgcla9Bgj93x4M
7vlEh0nJojDKBNVRbh2xgsaz31b9ZbSMT1jf41Ep8UG5N/lm1d5H5IJpJtsc70YS91FMMRoZ2zxk
91HtqSij2PR/I8MxorgFN1N6Rq/x0GPX809uT7tRvR0wRNdFAuh1Ypuxc1Ix/D8kWahdLcFalLPB
D9U/46sBqJg3y5HJgXrn1FCozQ10Zd1Hh72FFf5+l1b6uHcQIqpkO4LjmLOQxbqqXl+RO1/dJkaC
2DFkmscmRymL13Th1/jyNA5QqSwwdtmH4gOw55TEEwEsFdekurz+JYfn4oaP9wbvSentonvJBSwE
RNZI23IcN0kT4PZHxtccVjerLKBAyIVdXvDNdtw8szwf1cuxdPqLTUubMuZLcWVStJwCsVyK3huk
D21/6gyKa1cuzBB7dmZsLkFgJx76VeeeGaIvtxmiusphZzNqlDFW8Zv/S/BFtp4WcR/L1oKxCv2J
81Tr4RKoLl6Uv0/tzp8Um2yajPbitlz5rLEbLc1TE8oCYQXYP0KH0gfRgIG0h8uVumzNfdcddhcq
08EPx5zPqrIWxZ7GCeCi79XMTCi5V8/5KtH8OIW/7IOrcp/RLquLPODjhG5D6VbN5UTK89+bhGuV
3Gz/SKGCLI5uBZ97gfGPh3j8N5Jqt+SvF5gXUC9mlKsuK9pw6wKYbXzjvF9BxRMDbS5Le1iT4WKb
uhFkxSL9OraUO/JGgOEb0ivSgAx68DCXrsHCMMrDNmLXbWoDhWiU1R507M+yi/TR4zsF0EbqvOdo
zqvzTENOFhSB6Rbqe+olQn1LoQq6hOsz1ttGuN86YhYpYRLUMRkHQcJmFK+TB77N7A6Nk8uDJMX+
1VTEXqvgwAyTiWzDwocPI3I2rQhcnc5LXSGdJ7dNDby9RL6fP/qQ8VjfEmCgiExoCYn9v6rNjNet
jwpfCw+1Rsez+wYvNGKke/1hJlf9EwyXBaSNfBj9BQBKLZJnF9pV5RHqxjbmSr80dhM+MJRJYXFu
Owhevxdqx8MDYh2BTBrXmdFDtKUnT+VPgC6d5meRMAmBQilPWJL417U3dNjB1kzS1qU4EFxX5B1Q
nPQgspQ+uJ9rxsZFaeIUgc690gbAKqoZBTcAIfFkpN64rnamkPtqKaN+c76ubhawRoXU8tFuIlkc
9V+3asJKkcanexUTl0qAgKXSOdoaaH2E1OybjsagFC+d/4DeOz36nsbn+cAt1eeKew86qI73Vnh0
8l1DJGuboMleQena3kh/ZSeUsDXUX7ComOBG0Fw2ulR2YrvNaXsWWLuRZg+3OBOX2xOO/sbbyB6n
+OoPllEkv4kNQO0eN3rmtIrSKNS5M6k6PxYzj5rP0rVS6sZH0eVnu8THGSRABKxVawLfwEdZ/3jM
ol5OrjMhIi0cb6/3rhCXaWfyGHP7IfYIEbM9NsSx4dK0hkWYET0/AnKsacTBiBJ+xKYZtEyhvUY4
oWnS4HDwdevNrKioeEKlQEMIvogrMby8Yt0tG/GTdUu4EoAMyyRj2GSj0jMOv8wdGfrCsCZTsk02
ctlpi+zGi5tkPBSMpuCnZygG6GNW3Xbavd/RQtr69UNgywL33eIrxSmE1udIOmWUfQX4hl+Tno0o
JkCcJLQxs1o9nq3ENJN0xvqf+eVITp6rNA+qOAgiZ4QzRkLfwI3mVqaRpBmSZlGpNo5cM+q0eL7m
1Ovl6MEcEZjCTA1Ax/frDGgGyHzsURTOshPR9PT1IxFExyQtY7RCn47ZD7ByReIX+lHs0W97kWg0
3/hYK6REHVXGda0FDhdyih1VOUmot1q+F4dTFTrVyHzOjLM0ezBemPv/nWxmwDsjOGYgP3DCfdCE
wMSzE5KPXmd1MzSGgL20PDu2avho8WwanijEVeVlgzIxW+HYUthJxLS48PJmfwV0iSz8bLlket36
QOAfqnHQGAm0bAU/SUypfEwk5FTmgevUsyRAPI/fybqkNB/1ZQyjVVo6VytdW/KTSAMktndzbcUk
lC4Qxp7LpIgJYBejBEfyX/AucmMGf9KlBjSJyujSmHFZNhLavR7Ik236qyICgnrBQAlt1QMUrBxV
ngVYOlqghyi/UuvpfMEkCZi4FcUdBCcGt0QzsCL1TcHsI/qy0fnxpYpVWHAOBIjFwy2GcZEsgdAk
NYZkhhEx5i3TwWwXdFNlCoQNQVT4fSi7v+p17mg2fmgCvDidb6YY/+Wid259Wm+WqpL+x3qz2Y0u
1utPsRi38Ss47ofuVv6zgGRa1n6fGkiDRCDI0V7e2Lw5yeQOXmePIUwcJeK2E6pEhLXuEPSQLlb3
5cguW5a2fWnKejOw+7rNryWd8ULhffavcDXQ4Yjf1LFBXZYBs6OJ/7MnyzrLjaGXRcv/wa1SKI0M
n5EnVlFySMxbKAUYIM1l+havqPZvHPfUxzdG9HXojoYkW6NE7Hrmf09ORDMbcNbr04xGDBSqQatk
vL8b/COZJ26Ab1K9mu+vAf5eGUx9oB7L9sREiydBm1MFNjw7w0tsLOYdlct5kyPNlHKjMHCT2eIc
s6dK5L6Q8/OjNh5jmHm62GDiaOF49QHwVel9PEDz5/3HFHjyWys8zDwdKEpI0aZOmQ2TBCfVnXff
eoJkrEkcyG3J/1xybq5Sqfx4SZBNrZxVzNQxktq63VWBPPZINnAuDfDlZ5DHCHMIEbLmeFng9rT6
V0bQfG2x1PHIMh3jLsayIRGs75fkRkjl0bRO2T+PlDqCqpUcnhkp4SLt4h/yqqid8AyN7kx6k1Ao
1JA5aY0QwgB5L2pvt48XT5O7pEUsr+AQ6SHmsqqFwR22TCMUC3ORUV1kxTm+QTEopkUsGa4a+QMb
tb9S3FFmkd2AsMebYc/WvIAu/22aoYbHsO78gUIGjZTkXmvaEliVgfp9/KaZcWIdxux9Cq376jQn
BFJyBtOISALCJC/5uTx3Ce4R+rrSmQeKvsKewtfgm+90zOYcy2XzRK1VHBI1enblnNOBmYlAwsR2
1nct9hk+QsQCaTkHEkzNV5XjGzC4YRBAF/SoVF5oHiMvPY5T+Q19Tb8jBcwuyeb3qhvbrZrp+xvT
ENULut8FvXHyeXV4ngIuX3CX5/dTdeoOl5HmmhQ10PMyK00Eb92lNzesIPi+dN7OWq0LvsPEfN5o
Dc3QhuPYHOeh0C3NHSySdaaSHBdDgD3DIBgNOQSNKD7cuhslJklHSmBi5Zo1d9t8cYrTlhR2grYs
2GUhluuPULOjqiQM1hCvmM5g/UOO0yNJ2KHz2gMZhJ5GbGcIwwiaamBV3pk7x3QUtznwG464waSX
fHiAg2yAttwVOK+U8xqW8VnTTfUJ49oYSk8CF6H++yaNZWFmYUVB1UnlyMgKGDNqcaOWxyyZCPq+
+Y1Q8oKoC1umS5k6eAKpip0Pb+6kmNgQTAn+k5NrUGkJc3wrIg65JE2OdcigtgVsIrpFW0XWLI0a
rF0UPlHYxBRJmzN8x4SUWnxX7bJ3NbxVWCK3KFT/+Ka/rPkqPGOoKrpFrfES3/Pb+Yn9doDUZND8
BfCQcGSKTJKmcCZqYkBWmIzd5eHx5JCrPZgZinqknP5C3MB5Q1O3gH5CfdFNOmeORh3HEMMo+XWY
5hVoJ1ZIMV381Kl/HYcgxBSFscTr3qKnxDWjJ2Zu048afgP+z7dDj20riG/ltdyrHwrU9r7Gcahi
tRBRE2UhKNzpX2LCRItFhz7s9HVfKE37663Mkv0tb1Cp4ziNRiI6aNdQeV8ohtt4nHUVUs+63U8s
AtuA32jjwhPz5LaraetSah5VBV4vqFIWRO6ehXFaUSc+If8C+w9jPWxm1F34dH3KU7Wy1Rduk1nU
bp1EZQq63ORwsrb6kQqoShgVu3h0uB7Cwd7fwl16CAnFckQC6GaS15ykJfd5bheGxRtP9+RMRP9m
uRm3aM9OIXJAiN44EJz59gJWF55ifCTol0CaS4tupnyZsvRda3UjEJynuxgQHwj0uU86MSZ4Qp4r
iGoRR80dtO2cvRilexdvapaadsBmIOXiPps2fm62JW89i+0vkjFgHZC7MhyyuAsHozN6G65QMhsE
DsJMyEKkurS0IXh1zCXJ6eBcq69RlbTN5ecvPMEk5ommsi+PR9GsjC6xu9VUzQEE2Y4y6ZTKzDOg
vizHLVS66ZLoHOW2DiWzqbtLzgB4MVXSWHNXBPiw7+BTZeFLPnpNWECd2d2JeohtIjW4aBsJ7Vax
Zj2ECtxaPkge75y/x/bX1hOVs8nVkwfpc7+VJH4PCd+0wFghCLr2varDmrqQ31CUcDWHylv29dp7
3RAzCqIIF+GvZ8i2f2D4T9phc5gkxcqMhy6gZAn3J9pWxyV8BAZoljDn7D/5/i5xCU+Dzi2ZNNBO
Iq9udMejsDKXYmZfSwquTEyFpQTegUB/rISpMzBOgorE9fjia19hbNniSOXLHEVN9SbupBajo24V
SJw2jTjF6aywC2g/Ju93REIMgp9vgOYVZRKeLVfLUtqbd4wEmsWPQWvjDCLwlkN79ApwDghIvMc3
P1Wwpl+Bou2ySFqvaz3NiN4ZbzC3KeiR9Yx+gffZWUdGn0iaC9Xyoua2RCzfT9TCSqoNQ8RTE0kV
z5yPxdMtgwUfYIcf8A+AkdLjHKbcouh8nc6u1uK0uu4JPwZh1RzS4GCt3Q53uKn8HwBtdU2zmlVL
L2sDA8GYixp8iDP7MsoyajNeZ4EGtReGHOjtutVgWlxCWdilCSmj6syFIjjo5jMFut1Tt6PInzLs
BnUEW7vNM95GH04ygezzukJdzCTsV1eeEho/gL09UwzWPx9Jn9PiMq89DXfko8+RWoBiITfAXxMw
IfcTrx3sExp98N4rgVaWbu1AAoNipS9P6AkUs3dnFqA0MEmPdjHCUXuEWItP7CKYdSuT4zQIeGQu
aTfP50yAOc28ijG4TNnruBd+Pjm+VODAtCRuSbfiyLj2Y7CY484+kx8o+aQaEm43gy1LjlnNMYUh
DDws13qTXV8HVkrTLsd97Qjz3bNl6NG1UJLX52VXf5S97RIFCx0nwaVR0vT6+fwdcNGJMUWGScgF
84T9oc2+M92LBnw4iX37wo5SvrIkHtV/qwjwEZbyxjiSp+ZQ8lvVIMoUshgEjNtSbUt7XXRJA4hd
kYj9NwmhxYKfb/Df8ohOU7VyCGovLDgceKt9nKYdZMPaRVLSjXv/BysxlXRFEqvgCMDY4r97bKmF
hM1/sADIfBr5582+WpscIJvBC6CeJ/6YF3khfIk9+cH2WtwQkf98a3yi8e7kfAI7BE6x6+n1fxhN
r4wKSWuu3UjPy4s7CtSVQhRFojMFO9X3FrQMR+1uf3/x/0Ym4CEE2ST6qgFsgdZLFQKAj5y7wq6R
G1W5LhmPhwn+ujRBKtpWx6iHIJ1A+McF93MFsgd5b7Yvcp9S1yWDJM/bYhSJ6WbcR6CHE1Eo2E9o
r68GxDkq6va9wDLD43S9CsAuRs6gBGE2nSQxAnHyy6UxwugURbKv5xWYbAquvoMhA9nfyY5LjnW3
68v5sdcyt966GoCUefZsYsRhi9/bsXwXFinbAacJUqRbXzum3ilQXODeVGOKGJgARW8YdhDiv3kV
sM/q1PtCRIWZ2P+FiehujjTrLeArWNou7dpyEBMpOvnHq7Ze3+0/qDU4s4iaMl2wbk47LjuFbNEh
3ehaz8PeQbsb1i00gxIPRZFN6tlL3d94UpnBT9wTh15WHoIy46cb6ZlhwL2rKnhqjqOVklSSrFNQ
OdVHVZzS7EiOIhZ3+R0A9059J1fLm5fZvXZeW/yrkGC1wh8K+/7rbuOweF2brP7Yi944Gh5xeGiv
NkdsBn/e781iwBcz4uomE9lnmYm0kS/Hzgw+IS8gI3JKqJaJwb3uXfoeBMlJ8x+mKvdRLXO9H0N/
vk1olrj1/C87wJBON62wEywQejMhU3jUAdyZzUmcjH1HEf4/++J+4R7HTBxXAlYaG4GDCkuJM0Gn
UglSbgTVCxIIDpTvg7ZqQhHQppKR6QH9JpK9GEr9JOuMPPAwtCsBaKWsu7hz6M4odNWuIsQnrrQZ
MhSKHI/PdGJrEzDMBd8uJ/Oyw1NitMkGLzfr5qxB83LGLNUyfT+BrAKDeVqVeTBufs3ZvSgrPGl+
426omeMZAotOn9wghH9K0mkxaq6cZP8IDSvgn3CQd+YUJz5sF98FLXu8ABUtvUKwKkTzsZFm9F+O
vvLDOdlg0c7Xr4x8aNodpGZRJf/r7ExDS1PC1bSQpzQtW5VTXNGhgL78ILNq+9awHrzWV+F8aVTm
TLNSPBWhTLK2flSI+2vkDQY1UOGd6Jd1nITFgL+BMwqbDPaF/YcXwSqVjAtrko5S5JrsH4nunTns
vzWpgo3g6cXNb1FNydEvpicSwwKJ3n/2rDgXpXM3SJrw2uFO+oHuklwiTSRPyGssbUOdFpDORyGU
q0W03D3iAvmvcnPU7DUE1DbL7Ovk31/1h8dO10tlLG5wVOywYjHcsA7lsyjG68PzSMXDBqKcuV+I
Szmjd6XTqdtRCVYQdO8eAqUECEv3N34JmV2yjr91Bjesb7lWQDbOI4i59tTvefvD6LWX6lcN+Th+
0fLJJcI50VFF2SZaA0y2dEHXV7q6/PdJuBcpNpcohfZRNW2RIlk0EwhYcByRLZk9K2qc3NMS9zNG
PafiNeJDo0uPwdpoguyO3YfBkjIY+/oLIdtHS95fuRW3wUyAeRMVoN7eLQyDBYvXAWvt1luqIIDz
RRkdRZasrlRP+xu+9AiyF4ZjMgy1jZ53r/9CfqR0I2CDUORJTAsFAEnuhdLogsgveF1FCb4NXEVT
iMFOtXjSkzt01RHqH6Tf1W2/98mz6xPKBuTAojp4zrbibxgKIBkczem9RN8Nu7yUCiDS74LCLpFI
V3eywE9heOfc6k1tNkfzIDFpTChUmA6t6iS8qKdg3WYVjL/Z4qrpprUzfnVoRknUF8NsGrxnr53R
s3hEP0arL6KZMOaw2cyJ7vbRj3P6RWXun1dc1C0oVnsIxb37VcsKU3QyrXvj7iI1E5at8goquElP
4RxlX4ReKoJiXGoO899HL0X9/T1ZVkMFa3tjQzDu9Zoh7j8DoVjYpUXYBRWntl+7xhd1/73rtDGq
tLGYMI6V+nZFxMc8MUNSgiOmO7UvVZ4y5T+08yXsoJUjVBqgWVrNuT+yS29Gu0OOzdrO4JSJHDoa
z5d92aMN3ojGwu1SUwxqBWLb/cv6oUYcfzOmCBA5klyRsA2ZQTYk7CUjFjJ1Z2VgNreFRz9AypuA
Yo2e4HwxsL1jgL2C05r4mgUvolZzMGg/yvDVi3dFPlv0f6oJMpPMcvYg6M3rvCbJBrG57q0Rz3nm
CbTcCIWEAv5S+Ljxbmcn2DRJZKUNDDSeOATZFVbV2G5yuCTP3wlWjoNCuZiKmPDLiwXc/JJBh3oN
nlMlMCriL9yUTNmQkiKXzSsXXi3lCKc3wT46d+fuc06xl8on/HRiDgcpkC16fsEG2c7H8JHEi49p
1+0zns+JBy3M1pBzYWdgnpM9AucpfWdQg1ISKc6OjXjIi5D0GFcIT4pb0eq3fIVX5jxUULfT06vI
hfulmhjwzkvTMCa99ghI6lcD6iEmYKPpqc/XJ6QB6frvnA81+NGeD+vXHg9tWMUxJw2sp1Vgh4h0
vURDGtt2oGKRnSCRD0Heg8DOBhjfYUcXOx2f0Db+BeJTz0ozk5ylKVu4IwCgzRFx8YCG0rrWJlh7
UR8W4zeuI8MbqDeZCLimMCZDC8v3ZfxnSgLerTqGbjs+/JkGDnTq4oMwWg66LAAvFFWrvsjY4xaO
Cph2FA4k7eexXncAKC3S2tfgUGBXQLdyS3OSQKuW7aCEMt62ZIqb+dlYuEkJpNrqB2RoDMfmz+tU
sdW1V0FyYHFEVgha3aASJlAQzUO1rd6+3w5lq+PV6+HE0HiKzjDdZZWyWhzNJ7gcMU1lq76DP6xv
lcG94RsRYaY9qbhSe/V1sz8De9V9XkXEG2SkgepQMSOHs0b7es/JkoXud6UFAqVo+42FGlP6Rqxl
DD46kWkRMYKoC2Cz9DRqS+RRbv8mqTHJZjzqpYfAX6rJg67d2/hyLwh8BVQI7Y+KHvhzOIH1rjQi
oTpzT8FM7w9IhYW4CPVZIbu29sbOiyYmEm84A8CW5Tn6ivNT6qpabO7zN5Wos6xKU3jMLjjswWNt
m9pPfK9B6M9VrSdiiZd1Ik1QeU1kRHci3ttbVWe1YaWILZqaoxufWPajHlJfGU2iv7ttRgsLHBlE
cgN3vaZ5YK6c0QHi7TpnyoYDywVmpNWmvbs+VpH+xlEoKk5t5mrkGw0NZKI1KblBz82aIvrLJhlO
zQU583r1ac4JFsv9Kn//ddoyskO5HtkpOFP5GSFOKODEw2+nMTwaQeSSe8slWzlikhpgjJ1hiGjl
0qUobY/dd+o3BB5TBS6b1q6FXUl/UMa4FZXHv4a0F8v1iIDhiyKRZBenRsUwIK0nMeF3I0ur9jd2
ft0jU+tI/u1OIDvsxiILZ62F9zmR/u7lqR8a1ymlOryoX/Nyt2NLnV5cGMnDKZ0ABE64fMvL9c4U
0RDVKvwHxAIg2SVG9t9+eWcpx5t1RW1jm6AUA/lqk3sM/DhXbOwdsYIslwIfNhHzjStlIpXF1VM1
Nn6cG6GXXTtKEjznMfHrxmCLU9YXBH8shR0gqtDZ6y+vDkqq+u24mKuhbgT21iChk46iskQ6Ou8g
kuSIPIbpNqtMVzpkl/6kGtV41JzJ+52qQ5SpolJUgSSBIzC/FEgDQwgBr8ZjTTKtvXzkF/SEUAek
7DfkmLFM5n9CDr3oOxYBlt+IiKjIPo/y5UueEolxYBt+IN1g3UFb8F/ewSTZc2TxckLuZjacUMoE
xzQx8axMutnQAKJmbPfu7Si+1imcZQ0jnwtGyDy3oud/rdWUVUFipkEPv9ASgBu87gr7gh/sWzT2
vVxTT4WOvRXQn/IOuXDjPnHMOZQGwtMNcgMaSuNFZqKCcpOZzfRKjggxJ9B++htv2bVSCyBI82B8
4CIksJDIklQw5PAbmM2hN1EEPw2F58VJSuVjY+ANCdJoINuz5lemU3ISfFSM5UQA/UVD6CkvxMtR
EDf3HoIN8s7GVjH39J0RzpT/mSVqQeJSsLNndppyzpU/nBkq9815aunJ2LgOcbXF5+s1Av3XLcx8
BgqPIUlxtASw6j/gpdEmysGxEt/lbYC4+745Ear++bsXo7NYCVDtxPZAs8N0LUCdlhLcLshP8YSg
BhQYWYZGsIfzh4Xb67KnUVBSZlUqOdDRJ6TrQ5Oww5d7PbwZc+U7j/l1n9+850RPbmvLwPLi7HjX
vYfT9LiU8cYYpZj2v5kMWgLMmb8mdk8pOHU/R2N/6jiden6XamoHNGtAfNkGnFEtC9vydtNAz0Pw
iLIm3O1dJQtGNb3HfiwZPxtfEy3N2krLIuDqg2owIg3FPGVovDxw/pdbCsM0LUnD+7rLbLA14/w6
IXPy/cP8u71KIX/AZNld2V3UfTf+1eJWr5NNEPxB+rVmWE9HgmPQ7JTrxxwJgv0yh4ChedSkoyJW
/dWYsGg7amcjjJ1NOAptBIoi4aP8nA/YnXVrKfKLPM9p1z04BrA3jiyuuVCT+K+PoQjBE+CR2OX7
LpbfULiGaC0CBAdwcnYi5dZyrBx6hgb4CwK3AkJfL1ZCY71Yv/y0GLszAuABmV3vY8I+A0mQkQ64
SKiuc+4C6aoMKBAo+T6wJIGPyUTb5ryqUCGTNQ6ldemUTOj59pvIyj0o2aVLosZnKWG1YRxsyJsY
hWvpN8GNuD6MWQVlfVyXXB9Ur3MvxwJnrWzFBOHGshoSVl4xph0rvKyzrGK3AOU4I05giCcoPT6Z
anz1/LFrlFa2QkUnWvhUbHyNTIM9Vmy4d0YPlx964b+D1mBIDnOZBs0E+wTXERWA7DuoX+E3VVXF
VFCd//6V3bJR8NJaXRp98v/zWqf5h7qhIgQxwAaUc39CsFu+/BrvNzyBPPnP/52EF9huGuvq2DJY
GqcQXLnWsR5z8Yjrb9CPPFUao1opM0Vzy7djjIFTwyTb9tiQOhaJD4LobbEgP0QGurBlFg3/4KdB
zMQZUCEYBNwQb0mx1rGLPi0xXtu6fTJArTgCGO6DDKzAF1EeNkRjqg0qrh4tODg3RaPg676dSucx
vVnj0Lcv3Kxw8qADtwbZ6UP13nUvl/xFfmbEnSR7xb+7vr8aGlQUjSMquxoujKZ+8MUdZpiUVlbo
X4p4nYh8Bb9k6uqA2OOaAjMj2xHfQelAOqPgSAbGw64LDRqp5jHIBqCKtYW5yGbPEyz24OGQQgk/
g9W9gQFXg6L7lsjqYaJASra5FojavpNnqbZIP3amgO+DKxhS+YfzF7ftJlSg0pi3+iMgmaaVD9tR
uSo5204YOvqywXapYP83PyyRK86OnFxeD2rdp9cCD40CJTGKMvVhgYBGCxMy7bBBZtyQG5yz/SQ3
1oHHANkvl5oleS+AXamlbTRAcOlF85OsHz0Yjk2ghxBT5c9yWCQtH+vvEW+8jm4wtQqX9uzl4wyU
RxahtAnGvkczAtIFXIjUPlQghsIg3+NbLwCS5rP0VHEMNvxG/Tnfc/tfCQ2Fknile7ZAqRABkIoa
3AS/PwEgomoazqn14x7ost0xOrE+D/z0iP12fACbrQ1Fz8pGG95LM4lq9/0UhtnG/Lpai/M/PAgp
h3waiQFCBsrjw5ZF6B9kbGBInlpJBGZBaASCqrojvZclCcCdGhJOCDcx8v9/5+Nl8tL455CvmM+e
0FXO0sUt5932h+cZPmXBs0PFEagcVdDupvgJ75/yH0Jh2VYDptlNmXArzFZmGDrbOLd2/J37stRa
6XJSNjrvSAfzqssWIZ9oIcuXXRgHuq+FdxQwIV+KzLBQ4OtPewTBihvjrypQaby9QiOfjOG3PAv5
1NEYDcB7R6i9cc2AKedPMpWjkSlYTfDGwqgcyFG8dC68zoC4ZwFlj6jelDdndikbweyLY5Za6mi5
z7cRZ9V3h80OXnLo6pOvyIBR5VYy+djXNnhGTZvrijZIHCFYMTVyymQTxo1sidOeNQiTPBuQQMma
ZRaoJRkBPpKWR9Rc3idRVs7KaexCka9G/lBIE/uoo6BGRCFeErCZIPO+TDdRMHJJ1arxTTHF6KAC
X/N/VudMsDzk/AP/Y46Red3CqZmrGZDXLdmZ0l4enfauBxy48pUvbclC5xHhgX/GrDUUQfiZmJPz
pvgP5CoBP0F+fD18NpjcfQGgprRqy8eltSEey6fFCMkR8uiw2mPVjfHqFTNU6DI5+oKeysM28+t+
CqEiyjq0Y4XASqqxAB15QxSL/28pb05A573c2172mIaUmPj2Up5ghHqkpbFG2klRKmGGOJaJT99Q
PeInvqZN0DOsY03rGGgilwgIzwWkk74mKa4VcgknyNsl7iBy6hoyyjm+1FQ8U2/HH/RHAanSnhz3
91I9rzNc4WVWE6xOMaT677R1Rdd/BL4x6i6bEZDxBlhl5RQk8LulOvj5rAY6JATT4wwvh3kzlctn
yKA4wFx0gEB+nzWg5OSLY8FXYb2Sy0pNSmAT7YLNB3WjIld5nZSF/mpQnEMSQrCW9OhDAVxsn1xe
0rYPPSb0x+HDLiVdunllAXgYFsRZfcboQ5OWPecnK9uuiqh34hXpQgozlNw+luhalb05Qz5B0qbV
mUdu/PlJvO20mHT9Qhl15PHsvJN3WzIgNICaUIau1zBvkOIp7IqAIocG5irPe40ZaGZEMYNEoxt1
/+Gstsrs79xFfm3k7+pOnaWiEg+7GGNun8hqed0kp8Ncr/Ttv16YDGPXObUJOE+G/qM3eXwgsl9e
QEkw7tvYikNIUwdKguHXFruq4KMnrauHeydTYJhP/3zAJzW4hirUkFsw2/MqCF/2craBgQgB9XgK
3bIpDU8GEvwgcFP7/JK3gy9OYqlKtuMjPq1HH9Uxw7DGWtP9+tYqbK+QbOJtW5hSOh2EwFSrY9D4
BWe9QjYnxKCefYNhy2Cm1cHkI56Z3v4eXgpZ50TMUx7nltMY0yF5WpIY0U+5VtIHtt6EzWTwO8hz
H8FrFH5vh32zP0+v2W9gmpT4deqq1Mr8W7dCwDW0XQAm9nHPO8g2/D4T/h8V2GcxQuwkzYSo4IOc
Zp59q8uB5Px6hmECd5OdrA+1efKFtdfprPsk5JgKzEuRY7DV5MpyVojLPlhua03DWLgA3fmv4iSc
G3lkf2M72YPAyMBj54a6nNK4K4YpZ5zwZm0aWRAKcazqCBiH3yoJ4gqZ/VINAeUroJcaf6q0t6z3
cAFRmiGrqhtceIV69uLYlbUi0WPWx2U9x9g8BBtj605uPEFtxfZ8odqFnWRQjH95u6EaqQTMJJ63
+zxjJFVQZ7dAxzEac6FDmHKc0cc3QgkFatiSUGGAQxtzasEgfbl2If0iugZW2qqYkMlnC69BdZyl
VUD1k0HroPh3e0gtcZ4QgUWznazWGif3Zzy5Ax7DhgY/f3CNMKblPKqYX+0qkbr2YmU2WumQPk6k
KDyNGcEWyZ1ic2Vxg6N2row/JVrkZExjEGQQ028vtxd4+H3C2fLeTn2gQRsM9msbpT8JiyQk23U4
I1n3ayvouuTGHPTAXZ3Pb6elGWzkxyWRJT9mgh+LEg4Vsbx8bUGYqJLnJXjphvqmQXcxWOdK0mbg
o8O4fV59aNKl9wL281ZHvqcXRssuP6vHTisVW0+xCIh6q31UrNkyHaJB98T/R9cfblcXcbn8bHK9
20Xc69cQWIYIE0CIW8nadAoORCZQalwnae+zQwxxMqeISkQk9DfOrKaPLshE6LEHijRgBGkOIYgQ
dXfwD1Wvks/yU/yTwMsz7jmA7bCR3j43sNonJbhDMDP9I3eY4obuSXlekr2+Mho4ypcvVO4UtcMA
R83Gv328jMoJiAuEY1zZttkvLg0lwFGZo+PTE0vWeaUa/vKLagelhgzlX8N2sz2HMeSEIxhVrJ1y
a5skg3VxLlR7oV0PiU6zwlOw3Y/HMp/v6Rubyk74/BpZKhdB+xHEPxxaPSjTPmxRZCaWmbIGeyEj
AGuCiIA8JpQzZFoCfBlR8qVP5qFPGa7RT9FIbyqsxBUbgOoN5VWDBOayU43p8MRoC44qZw2cQD7B
HoEK7Yw1yuSWDTzF1uyw7Visd+Gv3xCNsHqnRx6JwGmomWeSU3dou+aD1I3UugcurDybSn1PTEVm
2Qr1Zh+6z9aJML3KxcuKr/0HEWE1kfOEhf5XNWjID1dMS5GM6FOYTgy4pjVOYxjssEtT7iJ7yF09
ZM72f1+OJXd16dE2nUaQefRcJcmznO/xidu0dbBW1fVzND0uOBjRM6sDRHn6h/kjWamd00x8UcSY
MXEhPKmPCvbEJ/0rFm1bJSCP8tVq3hI3bM8GylsdNqgmJqZIXgMZoFqwelbKtke6QBW1p0H8A3TE
RhxakwDJIEz7vWiNqECDM/S9YHC5nHkrfgx/3S3TUrwB4Ei9o7B/5qqV/4sFBh0MeStNYSjjcGez
ldnRjitdMOaOmKWEt+689y6fu+d+ruYFvQtYEfx/0RR7VyR0Mpia3T1ngBRHvEOktzs1hn8ZPE+Z
xkWWShGL0bQdXuPHk9lqvObJknq+USE3ikHB7b8IPGOQQ5I9ycb+TZPe2n7X++6eUxNrRDIhWVxF
J7G8l8wSUU8N89ArieAO7GPLXijwMJI+yABmrsC6RTHGqP120IgL2zdpemAi8ADh5Cn2KnrS6Tba
LKHmnHU2U/NPB9jMtYSxCpSA8SJDTfB6WkYKeiw9ABFJ6vJ/tjgMAQ1jTO+Snr0424oFC4mqkfMC
Pr/GdFYM9GgEirTSwraH47MhV2090YgfHY8Mc4RJM6aW0a5M9jx4CpP0l7sJ5H1GT7PtKiEKJCwb
v0ei1rT+NrzKXXYKZGWkJVVZ6lcxQ5Z06DkokVo339OMxhymMqp8aHcvUJV/oM4zlJ+peP10WZMs
Li35jGd9n2/CySuCr82vIoH4ZJRrx7sPd3rjod2bIBpR6vJduZAA5ehjFmZ+NQCE8DAfx/9GvNaw
UVG34V4EruxKw6g+LlGviPBCcMnoCNcXfjbNTtoc+/1ZlNosFauQvivJQOMxBxsEps0UwpvvNHEl
F4DyYZsbI0rK52D5J6hv1mNm9cejLddIUi7w9EamaQJB6XqC5kouGl5iWZ8DIBRVtLhrZmQKDSnR
K6RLOUtr/HIWvdWf81Oh5lC6oMpidl+HVqaVekNGys9ZUC7DxUElgiOFua0T/7YjGIrsokOJk+hz
iQZJd7p9unJAx/g33Zwl4Mma3t16gkDXFWdwJUt2DgxNi3SFFexYN4LLzYRoYSZQjAbkhyQ8WcMq
pulsPMjMdsPD0vcljNzWJrXoKFYWVk2EQbJpqTwXzsEvWtUI+D9GJZVso5pBHqui9vr4oMxbm+R9
5VjsC1qZ2Wd6QW77dGXVDqr9cg/HPHMZ58texVQOoW7PhNg4zqCwyStbZbwPjUwYDpjqCybkqYl4
7uE5YCxhOhpXFJEb3XrLwrWnD07cxHQ+/8FPdV4mq2rDvFwnm7CXQcRFhVAimod8IQZ5aq4j2e+q
JofpauI/lld0+DCK1TMnRrMckAeEfoKQEn2OtsK1cSJxlaRmshEmPv+3YfoR8ZdFRLtol64fjaoW
mmO2wxZyhiFGjz9RRIDH7bhiRzd0kjRRAAYMd4Mpr6CpIUTQ7mJJpLt1xLDVQxGmQPUwmWjl3Ykt
4a7B7+dPh/GfJeOr+mP4xQuNQDzYSiurg71Mb62EWUD3s36/WGEX/evXN6W0IZ9m4RdmPBc3fZcY
Cxkmz7Q+JhftMxeLPkUJ4pYV0OVMW4yFH3OHbudZCxiYc9RVz9J9roxj8Z1ydN1CZV1dOkikxUqP
qDnQHy0AtbwhM3OjGVqCmtJ1+x+eVhKp5ZuvJ2XtcoqZHxzY2Z4rJO5cF2FMq6WOAuGgqDfQZbh1
S9hIe5a4lHCmT29RmV7lAykS/uK3C0TgeR67/yCUKFlAGiqZXXy52HPdjQp2XOys291qeOmOMSQi
RG3mndIMh+snLkGK02KAH8uRlCvOh7fDb8jIaRJAamV5W8lIwQ+uBrEndPHyqPKi3Ubj1DwwP28+
LgJSN4sUjiI5SNyrK0l8PtMKrV+3PTrcLZNWVMNr5/LYWHSS9aJgk9p2p37IHwBFE5Mm66ewQChm
ABnjIt5OoVqxd1XNX8OaSt3M5GqL3650o1/kZUO4t50li22MzqF/6pbEO0XWzYk8JBiXQsbWvM1o
Rwl7GyVyNktwL/7V9DRMFTMag3qN7RIIm36qHYraG1p497cl0Ngo9ep2gDbJ7PabqxrD3KnUpghz
Eg846YTSL+oyo8K9TcUlEoiurjYx9v+N2aByrhZU6C9P6Bm7KWVCBiLxO2dtoP4RGT8gkN4SxY2s
ghafCulKZBLmlQb67Uc5PJpeGTBmNFw0OrLLvv0z1mdzkPOxZ4605MsiEiBmsyjnNHVvLTuXKJkl
aSOY/XPsSgXBfYAffCGNcEA338B+9rHyu6k8xQZYkX/T+NFhp3Aim02fG0JVcGPR7PNRJ/dr4v5d
3u6nUntGi0jH47mpxjIBr/EOFEjtbhDLELkP8FyJrcduW+nfuInohuGpDUjgXsDt/4eigaqB2zfz
dQ+DNEFDVTzSgTNeXEV4GaJ7wQ5bDnc7GnsKfwgXEhRJDdlonIFGyPBQl98HZmZ3womxhKOpKgdW
7KyTmznq1CqQ14ichOUBUk5AyD0ic3EdU4vQKz2WeCKloRlMXJwl+zhIlwSKvEdrRGyPyYhaga09
n/ASz3wVqHHl/4gcEeZ4gvU50Xs4HM5x6t8seWAg/9i++5RZ9iT3QjxLDx/dlC/aLZFxaQ8MNzLC
EM1jw2WFjmCRdgWSB2E+MbWUcASvYFgeIxY9vWTtpbF+Ops7+PyE2HFKSttv4/etJv0HkTuyNrqN
LiQGEx+Wvv/rlq/0qPvornVggL/hENy6JPegkPPmwhXCmpJpfFMcrdCOTK7DskURRexyyRovcE3B
D2SBBPRSvEO6dPHjFpV/KALoxEqFfmLY7oDmPTxFy8uLQCRzqX5b+disaAUxF3sFmute9pCZW46E
usFgO1/A/I+tJ4XpK3wyKvEb7inXo25hDFtvls0TpFVmgMk+lraLEUJn8oYlKMgCHog4pvikhpk+
tOOUfpWcr1uL9BMAnI++Xtdm2qosqUuAHXYqJpfkeYjcM57UJu+8GT6IVAyVWKOb+e2J6jC1Cb4s
i/ZCCPXgD5D8/pLTVbZ6mjYrjRPcCkHgDy34eqdfluLKLbpBoBa7eN8a3tY5169KGxqM/fFeN+na
MoWKMBJZMTs9LAoOTqUy/mJWhlLR1a6YgEZRsMXPfYhOsXBevTFqSrr0/nD3I1//34ui53MdVUN+
h9dDyIdDYeJLj9K7Hp7OedfsAX5HALFr9fi7ubcUynLuV99yvYIQI1oq72gQQlmkx4i7VW9OgcVg
v0GEQ/siTKLD1PrNMsjQrktaCcgC0tAr1F1Gvbu+fE5Uf6P6HiNpyWvQ9vi7JxEiItKE75ioMinb
DJ+ZN9XI69/GI5LrMwI/MB2jOhAblMlHlyD9LuQValdU+Td+H3Rv3RTEQYmKsTmiCzCS1xe+OeJc
eUpZN6lzMw3GTzWcmALffpvzJd1WEVbNjsQAxWt4K/ofl8Rx3JctLUDWVZau/E8vOSTZGppO6JMM
cQK12qbxu1aSAV1casdazZyTwk1mFbwx5zfI0dI6/EugmV29N1kpd/XsmxNZRQqPQZzZB956t2Bt
jTL1E9XSq75JDS9b8I7cwELv1rb85vSXzHQwoX+gzTR75pkI/uIYv08wGgOTahGfHyv2eDfXlsgP
H2VPrZ7eCVnSFbg64S+66V/2BQOD6UtVz2rlGSypw3PM95Uyv5J+fwdI6Vb6/V0LYNupLi6c0y3Q
cX8AMVOA1hYFNOLc7kMMvSEQplMIUJplVbNhBf/ZtsbF1JFYLjlC+T4GbYrSetCSU1o22D75eYQ0
AoPRXLV+7KkuUY2eUS8IvUhBsiD+zJGjuq/vZ3LbmHa+skHNo4b+FayZOj1xX7siROBXmj430hz5
E/WdMqbs0xbjHToMY7hl61yZ/2fu7L5jV+qSmKgYRDfOX/Yxa0bJIjUK3sV8EKOaRIB+0AOhvslk
OJQuSNapfsaRorYyo6K9h7yQRHzHcU7qAuLpVctfDGMykBhlleRzKzBme2dNiRsxbVGgFIuJf4Gr
m2jiRSYxr16yIoxfagLXdFVDia+/7IrURjgaqmVHMRGoJO2gIvijeRVj+PtjtR+xjp8545lEimLy
5RsFe7hWlgrRzTPzawjk0jZ5TSdHvJhA0YM5qP7y43zuuj0MGFgK0+ZmMhVY6ehbdxTkJzsdGyiQ
8WTnjG5c0Ff7eVpnEFWQazoP3UdO/o4NGKHrYsu6GyJsgYEcBytBCAkIXp6teUWYfpSpD+Ey4gql
rGB3tmMVpPBlDWr/AO0GS0DUs4rRHx+tVxR7kpzjlXyUOVo4g75o7pvNSuGAcXMbSgGnrVIEpFe6
yz4NkRLeYOSA6Bc8nL9rAfFb6AeXrWy+R5MZoCnEbqPTaosHSBf6/ytYkdX6bRglnTcYidAs34D7
8MbN0Pef33H1+fdBGvXyhH+KD0B6VCzENp3bP/op8m9nrM+OSyLoFQW5c05htIZjrzSKeUbCGio4
Lx+mr0jO49iuQzLretxBHojiUsPK7TeyQhsClNCgLvvegVV1cVjjh6jtW46P529hz5CqmroGXU/x
H/+EMLyZEzMtxGazXw/SJT2XI0gRN4HRXqGIeRNBkzlyfuqNLQSTM8y7Bf50uFzG2IPxc27P2xHx
6jNqBeC42kxiGdsiGOPVPpJm3/OVKOlthE/g5Iv6aYFFe5axTMeSUF/ggKn+yXGfvkRk7ck4LCOl
dpHGltB5PovtgSpcHJee8EtsLfF7fEbPb9qV0wMQ1DoxXCnUe7cZUS5U+BWPR1by5DKOe+6qQFSN
/Wf8Gks3Y5zgNKYZ5Iwae4/NkW8ZP/UuEF+fwPVPxz19HdsWICzF8vNydkJiTkj+9V0cLIHzoOp2
ZfuV9FU+BVoXN8jMMzikEZK4RuWXYKUYhIZElYTp8ZN1b4enHK+Ml6la5S4dK3Pjl492wnjBfNzB
K3/cpgnSnQ7kkyksmgVRn0UpG082+IlYsfABiKmp/QjAcmboZkl9cwG5zRLdON7RAYUpxcZfs29z
fdNwtfb5OVCShveTaJBfdgSnEdOCJCYt38E9KlAgv//9IHSW3LAZM/JEjZKPdD6SJkwPuVk3aeaZ
m/0rg7g4MePaIZRvfSfHJuoAKeIxgXGLCDYW2J6VjkJTKoSQJTUyHzG4xR4q4+gb6RgK/kGw9B2a
Vpv4GEMDL0O5Sg37kMm/oWi6m2u0E8wX5GWPKyFCv5LRqe90JkkzBJ0mxehehIerVIZ7dABW3oQq
X2Wqmbojijq0p2OLB7DzucJYhuw76tLHqEuex9UNS7UlLqGUi86NxcdNZ9rz4F3NcuNnWFXJHy6g
aErtCqUTxvWlYWhJDi8uIYJOj5qLojcsBk2nX0iEo239QeXXNcpdU90ahSoBMgwG6123wCfqYtwQ
Cz3RqOpDjxSr5E3j/8hOIDSUZTC70sYK1vWO8i4sp5aHY0fv1eUkVNEnQfMpSXlZqPVTwUAJsNjZ
8090gsXRNnWyK/go55V7OE9jexcrCo6Eov/1klMHqJ0jRIobmJLkwuo19xE7GLTp+jmbDiukOGNK
/81cVtCogGmsR7zvrcKw0Ozq+vM6RiOaEccIdEeIivYJZV/lhivOzRY4GeeRScA6RWLpChmecRYH
HXI1IuX/CT4E2BB2Q615WnFsExIh/A2+Qt6cuIbSK7dPLDidz2EZ6slxXLRR6CHU+ud60Bae4IOT
awm7J39fsgWDxvnIev45XRJeWlcOU9skJFXJGUn07s3tHBbJi2kDM5uQgNXFpzLEACfQ7swWH7lV
t8I6VzFF7GNiTrsrn7FNtdq49UQDvyATOByLlEAk2sYn8jeJ6u4AzDJachikXNWeO/xIcdNSf57Z
alhYXCkehdhpqH31QoJwdwsNen/FZv0txtqcaR9IedAbaNZRB62eCPLb8lIuIxnQv16Sihx2snNZ
J38sq5miytFF81bbCCWHEv2sj498JkfTJTOPnxxqZYKxB1ClXyweL0y1d19P1dG7Uy9xlEWtbFXt
fo0IH6L6Qagcg8tcM6soK6NzJ9ro/ZMpM/osn1XS1RNvl2KpXDP9fvJ6t1qAa7DG6tHJp71zOiz7
/C1dikgUYSSBSMJHaVb51MrZGjFJbnEY9OuZYXyCm7o0GpN2+MGPfskmmas/WoHf7REbncA/D3/m
vdRMxFocghH0vGeuNzURqGBrr9dXf8/ow39nyQ0XNUHnf5/ghJcge1J5yIdHrbCZY8NnU56AmGIi
Z+EBstZuA5/fqgjQdG2zGTbv32PbMasc1clqQTNRezC9VVfzHHh2okWS1g/JsnZMZYDXUeTX5u6r
6Pm95Aj3rPsrfZPdl9Bp1NzYlZBCUzpnxSa+9CFpl7Q520PY70noPZBxmuqjS1MpwQrSqG9R/glt
aoY9ee/M5Y5GZJ2McgvoHNnh5n+pEM7HL5KmxjoZA8EIWgj5F91jTSaBhOaFzvcOk/uKNSvW4C7u
k28GVv5v+c+o8cYZg2pKcyXN+KOfhwYgEjRRufw4Y7OMukQCCIjuibnuDGZznt1HRYYRwxMGI0/s
lPtJ8rHgEWulVg5z5BNGRQ8mKvd5QCo4cJLyIefs1GrDqwdD9UWlsePfIpGHZFYfv9hAubJeId90
uM7zo7Fb7y7h2DjC2L7r02WprHGVckryBwbjp476E0GZ0Dc/3PyO66y5zdfX6wFZgt8GtmNTCy5+
/1pFRqJDSe4GOLLgTO/NhJcIURI9iQIdcPLojniCgYLIQZOHTsyHGN8wA0KBiVkzCB5xwOtvpbeY
ZpEkFELQLfkT/LF6yayX2WOZOZq8rfxeGLOg+1i4fB8ame6td1CvZ+DmNdpGthBJMsAa43e/YHyN
CqQU7JlJOjOX2Pn9vHQ184+U7rxTzJK2qAzRGVTG6UTaEEpCYnNQ40rNHcokePFIfiEdVZIGwQvv
PS3QjHKtQTS7JEZ00B+Vq8rumFg2vcnh28fyEAxNHJqFWtd8Pcl+1dwzLPvsAt4oE/e2qmX6GTDf
nuzb5YRj38GyUQzRr6bMg2nm2fHRELEZR56ERkA5br3x8Ronm7WG4tfhctFMgGlcYwMPfJQorUPL
CSiSis7VXsiL1DGxoKfg+WoznNkD+8lPMkPl3HCL8VDr7kux0BL7rHY9LtAD5/VM/EH4TYfSCxFj
jlVxdHJByvVMy0I/pYYvxXOhnG5kOzyFvDoQl4MIDsskIu5bbC/i8NA6xcEUp3MfeMt+j118kTch
sNMj1oLdT+Cn6fTz1YbiUHm4QwVkZ3iXVfLy7L1CYQyYBdtmXHAqWN/Su18xUoLMqrSulptTwDlW
eWdEZfRVo1LOVRJNGmsbv+BszimA1ZwNZmoWgh4FG8k5ovWqBxD8kaFhhSVsmnHX1SFUbeFjN5cc
aU3ItpW040MhOetgX3NBpjTsrOPXBX75F08TeE4p53GK8weziVOR96LO0x0AEzEU9Jc1fcpP9Hde
llDRhsvAhjOUdxVzwYtkJs4GfOOHsfv3kQ4oXhJOa4G1ZPfkz2PDtGB45nZBYApbs6U2wJbaXEiG
r7oEhavccvuixJN6TMysY5wSlqz1xNSJ1X+WPorxngm3XsT0/zLzj1TGW8mBx8n2GDq8h7W5Zpt4
jdypSRsMTxQ/AZ0ZLJf8HQIeqCSgiwsxUt1YtfDSegR/EosB/L4N/N8OqspaCc7bhHUjE4K2sq0F
uEX7bSEwFfEK8tBM3vpt+Un9YHcnXKEyU4IlNbjJToDlJcHj3AI7BufcdT708dToAgIyvabSZI4J
4qIiK0Th9gsk+UGYUqqcu7v8TvCk5AKpHf0O2I9pjo6QXcjsmu9DoskeysIMUKjaF2di8eGfYz/y
RERrZ5NSNjFdJPucx2xx/M4t61+RBe1fxsO0C7Lw5mcmwE26Qpp4/OTERKLHJR6pAGcsCjS9Zpxx
peZYSIMJ/HrCs4wPYW+k68RqaAIBpEFLgb780uQZdMwj2H4Kfm//BirRUcXV6avpxc1n3ojSryru
dAyQFWvS5rWd86/OF5eEBRE7ORaP50z6/DPOE/szNdJHemocTnAjAUjTrY7R+1zLQkIvfvCpfK+p
eFkq+W2cmKVjYEc5E7yQw7H8f65UStTfOLmYTIel/alB4creeQpPt4IPd9nSU1ZAJpQP7vpaS79u
gpHlYJZzi8StDNuwSgBhlSoo1+C1lTpXQvkiR5PTFcmJacdaSxSCIwoQTgt0snxVcSm/kpVsQuAp
L80N+RGIVewIVs3d4aRwsOl6b3BF+PY9/EYV3v7Jxdusy4EV3LCS0VqLZzPXT3ULiYkPCiVsSHj8
czGUpljoF0REAEfk4A2oshx682mT9XOuXPeZNvO3Iq8xmukQ4F/riL0MY/gfEZOPcxSWz+sPaTPM
B8MI9fpBAS+a8mAvoMspQxNbzfn/IhYXnE1UZh2bIjSA8FNAlvRDp/7OlMRJJwS1e4+ylxiKAPub
GxCVk1K5bVvZfkb/lWLGhgLxRV5EwGvKty9iYfnqXKZiaavLTnplBL0W1Q8m1hVzvm/l00igRXIH
6KmhFh9xylKtE/pV5jgtiDg/qkhySThp0H+uFyS7hn7YZeAyUDXcHjK9A79oZDxPjelrCycw0rxW
5UxHQua1nxXMyDXUTc0s1vmgekZFMJTXbnjTf+85/et7xQDBpxf0+eLgbN77ex4t9lze8WLaDW+F
55rV8a2eeo022lAJgPRz32pxY1EisNYbj8vDNB4IKx+V2mOhzD51q7OdNUKEQtywkjXe1GrXUoKg
I+6HWXrKZx87a76iR0IJeWWKBRB7fURLJJqjKlIN92yRtVRR0YrFGZBWb8McmwiHbZKz9RqEbKxb
wAbmK7VS5mtwrr8kipegsO2kbJu9zJizo8IfMNRTiflwmpwYbjEYSgVdwxOdS6cfD0ICb0Os1UNK
BVGaWpwwSm333u/Yw7oto92yybCX7UkZsAiRq6e6Gj8MHNj2A/xWsOETxVIAoiy6pPZ5Plq77JK3
RlNmevhLtMzVTh9ZXsVxYK9jd/IuCW0Tvf4ZvNn7ensRnKnsqmcoYAxIG56IRGHYcyDfE5Gt1UmU
oScKRgShVrpOlTEdbdvwPbhCys4H/9reHcrKlf7XIorTaST1nvGOPIarYDyOMagni7WPc9UK74yx
LNyCk2IP3NZVVUKkipB0PGJyCTrf5cQHqhm6mYZP0fCOFCq6JHRBdtRbphBDX2wWKtojjDahxSW6
JTaSKbmls7Hdb0h97hEYRQ8/rawvYXCZvXTCa2H2d83vdboI2bNSb+YgD/SMpWoJ4zDDRwjgDtqq
lcyW4vR/bwOAt/f5MGaKm2etbzES24KZG8U48wOuu6Ms7vvf+yXgTbWdsdcnhtNqXf4pqSSKGL9W
o+eVxyuYqxVaW68LVV77V3rySZ0gN2MVNaz7eWfGlCPwgsqgEpY0OjdMQmSTD556uqLseEd3dZjH
7/3aX+ynJ/BOhwG9TS8Gj4FhxWhT8zDqYFy81cmGXUs7NJPlDcHfFMZ5R0dbkdivTTKLLpuVkkPG
b0/QiuQHv5crVMYYAa3TNjyE2FWLA4BfmMmFeWPCIaH0MlLogFpcyfOb+78cjz+49QFjn+HPvahv
6T5dKqo6GB7w8g/GamG3fr3GjfbJnXiSuRCd2T1hYw6AnXfnZDC+a/7sgpWQxLcn8yyGN0D/xaEV
2z55HTJaquLgiBsW7AsKp96OiXIl2RGqpyJu+PP4tT5RkralC2OKaOJPP7BjYHzExuXMloWUlOT6
odelcxohpNxVVGJ7E57iRu+OiGzpKuvymB66dY/Hr/qLP0allcXZ8aUZUXKJPHrluLNs46E+AgXn
CuIu4P6HF/h8r2VWFeyTyFygMaEcEavltvmAZHlWH0fUtWilg5PNZ22tjJWxXgIvTRN0gKOU0eWa
kZkJ/tmJu9MJOA0VG9LWQEwIZYTTsmWX7Oqb/zew1bBLoTG2yM7n7bP041j/kpZkGWFgS2fIVfHW
cnuLU/vH555uLmAC+IkULvFzipNsMANtBuYapGWsnxAa+mH157XyXZnA8vPiRswdWGUjqpmlbU0o
jd3BWLJyzw1zNXspgkwhhcAQi67iB1c1+UX+zjPkGCTRIqyl4jTLplYTIUh2yHer4K7ecrrjNX9r
wH9t5NzVaaGjQWNw3DXhKSqF+WlAUnSgnWIpRmOPcPpv6Ee72ZNrjDdqqhRa84tDZoecafNWEfx2
ZO18oGClhqeoE/mrOEYGCR5plEXvVWVEGDm2dbnm2iLyIjlaGMgtP8CI0iOwJCExIGQUta3Kq8KZ
VUkLpYg6YdDIMV8dMbdxKGVt4eD/He4MEa5/2mrKURp//CV7cjjQEgIEgKezvkQf8r9RGFGoNKNX
wPag0DVG1tADXpzkzx4yP73VUl2WV7g2Xdtj5G+Gn7gAx6o+gctoTX7q8v6EHYQTkhQ2hm6HQ7BO
IcKdN5Hngvo/9Nb52x7FpQPPxNi5Y7FoWdHQ8S3+dtOC5kLj9FCTen0vzZ6Ls9Xc0G1vEFq6Q0uQ
aMqAIm7QuQ934DIgWGHms+qp3veai6H6IuWeprStwE8Ejshj3baJvEGa5GzIVlNuPuBEiozVMuYq
CyZWU2d5VrlbHZR6aLi2LevUq5wFdLIi3CZoQi/XvzFgFoL48AsEdMgRyiktRjFEeDpldoUfRH6r
GGlHJ3lIyizivQJzxNC8FnWvtigEx4HP1UbaIo1FFDaMMCgzVe5iuZGn9+u1Epe1vZEaDRh6G4mK
aO58qA8zzlfZI0tDEBVo2+PSXEb/9rqW5SJya23p0nGFezq0Qltt/LIsN7wi1wdy9HThozaKFa1d
Jws12lKjzKDZxBkDSqdC9CM+Z+mluSHfxr64L1zJDbB4EcYRJoZ09doHi7m6rFlrA50a26y0EeLt
o3uQpf/O9r4ihHhQdssnaIBX9boFEb7kze3h9Ro0JUzYAl9KBYHfMa2Tr6JbcR0DnypztW8vnIOW
7WXykKQ+Hp20vwey0crE9aCLDPm3P+LWfmmNNSjrsAHoVZLaDZQk2iOLepYhiCmYEu82krNWPOcw
OFC1SG7hgBmJZ1l988JOFrKM89N8q6dDJCQdNby3Qi3EEmx+wcbDzvfmdlWJYxNGK6xW7arwLytP
KgK6UZQuKJINYSwnkVwf5ja3M7i0v20Nn6lPBg3P+0W1YwOixpWRZisqLOZEAuogY0CcQdHwxdny
xLx7rge0/sjoZLidjbMqhKVQc+YaS+CcvyAT5J+xgGLthCW2HHDBnP/FrGiXAWBQuLegQF0zkVfj
FhKP6Fnfw4DWmJeECaolAQ1KX+GkhrGDppBhbrjedOWV3//VOtYo9W0gPn/Fz9WvJcRW/1yvxOF6
zZMyQ8f+7f3oa6fFRdAlEFdehULlGxOpi18U88ysUkyb0QZxbx5ROelQkDwBJYh1RWlS3qlCGg2K
pEddR3tekDG+Aqcnw7Tuw8sumd8Tb0RSMC9CCm4FVNc4Ng/dWPhwj+GEqvuuOBfkIDUndnhlysOp
6wHzca2ATK1wicncrQLGi2tB+Kuk072tLFEVh1DV7Ch15zd5++iqXELp4SqFKwVyIAJSaq8nUPH9
rqaW5I779kC6pKrgIfjTXn2yTiiTpEKqZlcHylcXgaR4PbxfqOXwQauOcuCt9RIURMubqS1XL/HH
RhutEJXPh+Jf1Y7KazgA5HhN2X88vS1I1NWs69O6M/gti+0jl3Kyl8uCXD7dNKA2EFHnJ6syphBL
geDy59aoobwdtsMkPzBeg8la3XJ3Ntlp3/WoubIVvlzxUVTQ6atKVy1t08aolqKr2h0+dRATr5RP
zjF7T5XNTQ8hW08vFjbQdPxwmChIQ1V9sES7FLgcPyLf/cVU2CfIflkI3ifA+l7k3Eggg7BXZRN6
zQxZJLxvPuJSK+yKqzz+kc9J+uihcG41s9nH1SMVuOFES9Q5J2+NkIlAAlFgIOJ4pbhOZAGCGmQf
kMz38cNngThDUmJ3IKIx1CWXZXJ7Ek2LjJggwe5v0l+ARJTkLfaF7fENkOpotTXdpiXR9JW95XH2
ZX/xUwoEuUoeu5m5KPNuQpmGEav1qb8PVLOZYuuZcqYB/6YzlktDHX9ywoJyV1+Z2lN9yHdnFiBn
cGt5/bAc481jbdmCnMvrkkcAc4WxQT8j59usU3lpF+RTKYs1NRolmRjk5nEe/Vf0+HDRea768R4e
clPq0slRwOV9C9gK9W9LxFZie8DQZUS1kMPjre0WORbkleE8C5YeMFOb4wjzIYo5y9X51iRf65lH
eVk82YR4QNR5hgRwVkCPoWiZAZE+QYk01qarAKZOjfFvoatPBZogmevzGLcdfk4PoR59VQXSo5E0
/MlhCnJ4+vqtMOCGWEGHGG8qC6Zn13wW7LjQEgKzQkYbA9dltzb8Ykaic6WKghGSaeMemquVwTq3
4jNCAkYjk9l2NzzgPIZJzcfLwJqFqDAzEkvmJdssqNnMtL0z7Pxq4Wac78SAvOO8kpMRNmwCldcP
W+vq6He6vPmHHKp6CovD9JqjwmJOMaQ50GUD4MKaRDWS0FeBg3e1PC+NYhxnNK8haiftA8hLdX4S
LlJ8gPX4ktMeXNcq36WwNtcTCgdusu62N3a1DKdX/arCIPeNN/VuOg9kjFqELpbKRzB2orAIPa8H
9AKWySyqAVs2agzzNL6Ukzfq+i7vxbF+GKETXdMrAKFYUDSxLY9/jfvcNAPltXYDrwe7iXGA42uP
lgY0IZEXs41MUxQWjKmcitwouJKjzuPBqYSobdERbnrtlKITjIfqlKWIxDzBbjBOGB0qr8ErOIzz
9Bj/KweUGdPbPR+qfEWrfXO3zDIFrQ784n6En3cmRrhZ6pei2c+etsNdGnvfIsDtSba8+5E6O6dO
Vf3W6gAb0mweIepjvIEx+nrbHvIZXFL23b9BWV3uguZdnHdtQLU+oqk6hVJvzNSr4QV0EjlJyRs1
sAv8YS/LF63kdKwMEGDQqMM7gGYKNW2NuO9cIsFDRWP/QEKBTbWyG9MNRCvFdargxYEtAaJBa5an
hjeroonrtaXKFk5lQil0DS8IfPp0YSUqyzZUBcYWcK0SIm9NWwMzHUWXYCF48gTWIRkRR4UBtTjv
UIr85aPJHBW5IA6GTkbdPTEBliRTe0yR7MBxfGAmslX7dr9FGe3zGvxfPEJ4VnAh//OLOr9e7ucY
d35jGPebKGs+sisziRCdlO3slgrVlCDn27P1k0vOTCjjLUr72coq+YJkbFUMnUVcXBuBLoW66kB2
DSOphrHV+qxe/PcOrS2vjx7iA/HmiaUp5i0qe3L+xyc8y+/iWP1sIn+EiBTG1Xo4hHFUXnI00mHv
ydmdrciai/gV/XA+LCJIwk/9R7JHVk71CKCELKH08ReRM90EnVznocy6hJnR1BF93pIZj3/w1tZD
k86T1FZXVUimaI2qxmDnir7d12T3YNzuaCD3LzAPvio8cNKgKXWoNJaxiaNeC9dNZca7hPZ1XMNs
ii3fTygl2aDyJ/mgu8UGzPsSNscjs8G98uAFB6AXcyeK4sLERgbz0d5LisLLGvP6DPFnx85m6zv7
oGqOWaOrmoYqDDEuS+63BhSE8qIrrkbpIumHgvHKGfTUEGZH+n9pp2aMFjWNODUixemVyuIvtPoJ
NjUoEbWONNC+kz/RvCMKTD0IJfkI1vTuJzi5V37e8aYiNqexRX0kqvHYUB60uIt4+x+TFHt5Y34V
/oAEVygf5Vyx9l4uZ7jmQoBVlmnRqoVnFP6V3Uls4qVul2cPYIYWJCKeVL3mgMaV0fd4ZoPcP6Ol
KBPywEAlikuR8hU4l3qOPhyJJTHGpo1U//6J3R1QUeovFbnlmWygz0JdJwyfLrP574OfWN9R3TOe
ReOb0IM7Z0Rqh4AaludCZMZYNWJ+gmCwp/AZCs7736W2RYGHD7VU6pJ9VVQmqEdAIEVFkPnDN/t9
4OlUEVHOBaUTyZPvnEHmIUvnVoPkgxWiK2qcjEQLUxNPIMyCRaN07iJIoQDhtA3LJLYRR2F/yt3V
VD0Fg/7Fqr34G51JAB/+xhK6LjZ3H9VRr4tNM8U/hICRB5B5EGbkT/xcagHcPZ3mWraeZ+5ydDVk
P7T3GaYOGpr4LofuQxqHhzhEmKWXxTSuQcsNUdBzGII0xIB7B2a/zDtdKkcE3m3hqNm5aQDFpdtR
vU4dH6QNNH7b6siW14n+FO1dx9lgwookNpLPd0vjrh9V9GDwjXwh3hisgvb+Hub2uIGxxfGJL55g
EgqsFVch20cL2UM4vx7VDpX+jiJypCk1Hd8milldAHfR2ytc/a0NNHpRN6v7LmWjN6PLibtgR5sA
q1ab71NrjrEDh395MRdgYBSOBYYf8IXiBSSyuAN8Yt3Be1Ep4GYPOfurQeb6zjuikdLHfpXseFmm
Z+F3o2WmlZ3DXHi+hFxk1tsXztqxJJF4LqVyH2djV8AKz03jhuA73IUNbaTj0BnZm8WZ8+NWGP5O
G7TE0+dUWs/s6CXNHhMEiwqdQGUozQcMeKTpxrkdAPTYJ160+J7q5nigdUCiamkV1vy0wyOv3nDR
oI76Rbk10VFjGiVCcMVI49YE/qKW7e6tzrlz729YYwnPm6N4PZ1EZIJ505bsulLgIDMVPkR3poZb
PWkeqPbkCfH2z/gDABlx5H2OyJvky5cfesLtJZFZNt72atskhnZ7iIAMhQrKaMswL3IlDhfLIR6T
B16oYSGBKPqMFEZfNueSeuRikGBy5FHzycG9rg8R0NQQHA65h0PGGmV1STp0kM2qv8zvlA+1NVLC
yPWGf/ZoaroM1OPbG8fgXpnmcFqM/Iyzg4h93/FTln/5DBAkGoYmLi198iheLOiIewWSgr/pERX+
R3/4Qvj3HO+XagZ1VRpsE37AnTHjxx8nJWp7zgayMMnQkMDSDbHMDtxksE6XzSUzzLQoTbRn0ZJd
Tm5AJk3bO+AUtuHoPx4PXxF/V/uGJ1f+AkpOMG3aQLFLoVnAUSxPLB2oqb83SUS2d0eJNmBaDiOt
Vn1w6qC6CtzpUPt4Fwe2ZXG7PEheCsYkZHJyKpxxSky0GSEK+GtFk7PhTJpubEixw96hJSW0n9hZ
spcG+VuotJ7fpqyu9RDHYKTSyjLYpn8uk7KzPqnV8P9ormO/73OSIQB1DXL3QNGVtYLoiVmwUwtB
JJTDwRGW3+CKszoxYNhwigugqNg2H77wxk961epNyi/uogB6B0sjAFlbbUtlTw3NV49lPS0m1DIu
7hrmNb/aZhKneDCqAfOiqyMth41wTXLV8RlmCmfV/yMufyjoHrOTjQOYFaiLQsCjsDQCPmUR6peI
rR/z/zDeVPit3iIZCSlsVywk9hBp+DQ6EXyf8CE06DiYjgeNEyn8Pxaddb/bRlyFdDmjce8raebe
m2cdx/5bNnO/BMHBS8rmlg701s4qZy+Oc507llUwRoh7JUYfrEYJZeCLaK5WRZEpMBBH2gB4dtMa
2LQ6AvaS0daGn2WZnT6Nc/D8TPV25ayymxKpvRQCd7SAQM+oV7hd8BwzzNDlk6+pAf5oKeTOexgp
5zo8BYCBV5NBVOP3gzoSloV4aOt2cBKl8dEv/EB+BSQe5eUpTlihRGmbj4s3Bj+d94gllxMP1ij5
oUUXoDBStwA7kQEh4CZR06gFSe6VAIC4dXqd3sRWegXk3naWa5GIBnhQD15UoRDQysU3f9aFHpO4
JNAuJwdRwPAGtktRbqTDWBqDU/DkihHT2JtfzJXaT4jHB7ZZIpcwxc19AwDAYRBrRlkIrYoOinnw
+4MDZ88fKVXZlcDnU30xhOdSYChbSBbOaOzz2/NjpZJFUKZk4fA+RIEeZ6ltnCNHW3tTZO2MoDLR
b2xElu9jkjPOO9wbVkWHe9Hi2r161T6AfkUzxNYaU+RrkkEcXkjNWwdqi5ul531DE7eh2c6V5IST
RGD5IGPhLlbmBCPO8dZKwtG2RA+gDKTU8NdNE2t0UqRYrJrACdt8skLqhYs4WoI1Zdef7vHpWyff
/iKVkmODhXtJzrP3iN0FbJiKhO/KdQE/ZYTHxt54uCHT3W0/IcXzJdQDkFe2A+BZfOwh5VPcX+Q8
9Zkw9KahNC+3x3jBBwaGC/LT/Oz+XvwhZmowEfDSr05heZI4AxrkgXFWsyDkOSrhAU2f3tatJLpd
C8LaOpfu26X3G/5sV5Ayn78Ys5qHWM1V/uMDSX7LwJXrgs7pNkjiUOVeJCGywm9jNzr0rXDE8Paw
j3zeBkFg6Zkghn5ZZVvXP4cvys5+vI+9hM2gtWoQCQFwBGrHBVF5/RvHfVAS8OzyhmTvGgvD6zxu
857HNniWDiefXP2BmnHNAEM30yrKAgsu21a2ZE2rZ3k1EijhizsafCDejaZ12GnlsKpu1Sk4jcax
X0RJzll7CdRQY5VSus9rCr2oPf+bP/RG+jMzNSWcGL8vQT/pwbA315CEUbMlNg0P/j1sPfuVh512
nqpp+RMhmnXHuX19xCAQDmQdNmqalkWh6HxS1q73iu/Agl4yaY01zc+gQRbV7iM+EzwdQ7iu3E+0
8h5qyy3XoxAOwL+U4+cRMsF/u+UM55odjPGPl1Omlgy+qAUms3Q+8tjHH7+WQvnCrTp8+9cjGhUY
C/Gg64VrMjq1u4wWd/sk9tzQs9NEZtIHqrPRknnZ9LEDYo82JKCYHPBtvn0xFydMSitSg7zBgYCI
2hILpI8qAUztCwXKWtKvGAjpR+7nLhd6IucZYsV+zOpL1a1sfubun/VWn1CSfMH4dNKNMMOezjgU
eW9Mci0BdJ+k427tAdzQfNzqXicwe1Ry/dA0KrIKhn4zlOIP5XZ+XmCkneTvM3om/51ypLWlJSpB
hHIWrkhyIUGPYqsOPdVDavkLeWywXUqN9287mXLd4boJuN4Ti0Go1A/5Z1ezs6b6wSHQwM3BATpw
/gMjBuUtnbmEGgPPjaVkq0aReHmZkRlFha/T9fcu6WEUacpLpQRHJfbcg1c2XtVgkwGBqDM26M9I
5sCaMwFiYzpeh63iosBFMXQFVaCg+67isabL5BsXtuL7+he1qlFbO6wEKM3t6kPzPmUHXG19LvbD
tKqXtPchi9vHWtqXTW5wmVqTGywAyrl+2WWHCBaEiiQCPPF2ZEw2ccfqva9lscgZKhO2aroEfwLO
BaW5zHmqWY96bhQOU82SZnCJUzVxHBLHD2m8lt9ppkOQMzsPSbR57jUcfQAFxJaBdfx77StkbeIu
XukoAGWHDOLw0Q8LeVvbZXeRiSH48Apm42KJ77gdrdDjHzHyx05g9xUw42dWgTKae0lRRiuHd/+h
zvH1Zzmvt3FBjUlQJQj6E5Woso0QsKFMEMoM9PSvbpL1XxuWX4wWj5VbtIKVQskvu8MCBUpJdWts
ubkg2AwbEPQ9K1Wyjn4Udf5mDVCfQr5V1dsp/6htZ3fpLHtkoAt4TZfWUwsNnr6Q7/KtPm4z2qYi
k42UkfjZTzmLCrOwmcOW6sPsR7mJYV0mZNdAaQZGIX95nWEZpzdy01py5SYFRqTcSzoYM/9QiTrA
LohRrosJMdOgk3g9yNoWID/NAMUXnKlNLsbW5Hc8DHA2oXsIaaN8sNtWN6lqhvtNNNclfNwiMwqi
lpf+RRk6ofK+125MPe+/JpS09n98r2ORPJHXQhXNO9Wwt++Q6PTjEj0TpXJcr+waPg2th0H3pUrn
u99AfqT6NWa/4WJsq4MGI4EFvzOLf1dlPHAts+cb5MrDoGdnVkQ3RmzdPlSf8qkHid3bPxNDFcNv
J4W+fQZO8hHez81BinCxAyVHmQ2/LjCry1hn1Zeaa630Y2njFBmnbS2M+Wxj6H9dW+ep+DPZjkJD
ZwFMGqPEsGpu4Tn9CPpCF+2KtcTq9AMozysaPlENcAYQzw/RVx7Pea8tlk54NdkCvoPmNW5OA823
k/P6vB+B3ieEHzxyRFoG1qYB5Qg1EA5LriD99Oq5TrpUPRajGDyqeOrxmt9ujsWyPXci2xxZSp4d
/bW32Cfptyo8u7n91c+lUyTRhNiaLS0pA+gxxH/wtP1T1XzVyzekM4kVgNhzZ59+loB7HV557YKv
G0foziM9XegwG8xgtxG7eYrm+BbFbVeNgg0JIgtWnEaKUPRe/KF9htunlZsqLqZrFXdBQlnKsgm2
0QFh2+KbnlwqwmWDTLUy/rQ4irkDGZeBZ3VU8pBGgrEFaRaUp1DCyp1j2KP/RzNleNmyeZSzZdGC
Myv8ABe3k9WSYIYoDTScNSKpLdfdofyla/p2Zx+Zyk3tCCjIgw9fD8P3o4fsbgfeSvoiv+KTw+a8
EArG30rmbuOaFYmcbG1IiKuzmSc6addZL6h1Gdevd+j00/fkpjYCaGrMeN6fKUnsCiOxIINFlxFT
UVEcCOCZ/sklWULerVmehmsoWQEmULCVA4PBwSbD04NmpDq52Zi/E6rxOeh0IcmsKToMmHxHD3m+
98YmcAa7HNONQhAdVIso1tT9omE3jx2qM8iAw7t8YDduLe0xQpNOmTkIPN/HGxC1Mi8V2YvTRc5S
Pxrle8BOmYvQJcCND16Z9P7GxyH7J+BimVq9RTDrMVjreZIoiPAgrhrk5cHBrVaQ+YKnJDIIziI7
YhKziCoBF+FEPqGnPdrYGaomECNpNQE2/t7oYPMO1DOO+DPQcwNV9JfWIn84Z+/AlspbhIKQCuK4
X7rGNtgEeFxNA6JMyGaWkYscIvz1RsPcKC28z7Q+nHS73o5LxTsCu65r3NrslFApNYYege04D9zg
a+a3WwiWt4rS0mxaYMFZ+N8QZzdczXLIGbF+SBUiE3vmU9HSfPnhV2eo0ZKXxdjCKcOV3prBWHMv
hU+8yhtRMImeTlh1RW8Tv8O2axh0aosCUvjuY465tX06Y/48S4MuSdOONGhEV75vgu+1UXfnDLwl
rkD/PS7YSQJQDh8nAHlknc3R9IZd/aZ90QT9cySZ8UaSG3cJd28Ggujaq+/APlam/gOsa4n/BAcj
VeFJyUJZqg5+hfU2LRnfgt/EM0k99GufN/EwktnN2fDg4OCu1QTcS5F7+INBFRGwYC4EkngniLil
M50ER3BExaImZCNaIyMFNFfiltiOwtZY7RmIAG6lYQmqlYyG+7rOjIHYXHjk8M3KUXmMX1m++hxQ
f4sNAkVioixA9A+jcxrSTFpukfHSGGsVSMpvQH0VH8U9Rxiuw8Otk3fmUGeZXgOsgeMz9wt39Nwv
8n18pcWecBGs8iHLEojzyVocOnW+iFAcc8baPE0vo1qWCWzSAXsq6K6MqqumGr9Xv/tCA6bhvjU7
F0RAiLu2W8KAIc83Dp86gyaVDBpSaDXhi3oHS39mjKuKY525X9sOevIM+FOtWQvRrj5RbGVVqjZH
vFD/nj6eMEQSZ9opja+LFzzpGdGuxM6aZjS5IIuay5RFJiQy5qzxj5rT8gedJJSvAA43zm8dMmyZ
dPg8tTYxH6xqYApjo+khBzIw+3pBPOOiEYleP5g86EhNs5WPJSclU9d/L/wtLPgbm9/7lJwa5KuG
xhJQOnZJ/sCuMtRDhFtaAayHikEXy0GXu04VP83vQbCgLzRhNYSZZJUugzvvr3HFoigB7WuYBErm
OqjUbPJnzXEMzCV355LpwHfTWNkyVVGPHh3Jd5GNxlGHf4C541JXtZvNiyfd4mDx9slppeUOVRDw
0Ms5LkdqtDiBbg/+HZBYjhQoMHYkGNMrhv3xSkuXmdSg9v0tVVzoZTlh2Sm+2DFgRQB5YVYtEqOB
4KGQjeztDvWaA4TJxNc++Ot3AALwQn602cA9xOqNdKGTeesSECPA+ibBhVRqASAPIFAZ9MNV1Abl
L9+Skt4z6vR/is2/87EnglJIgJSnO56w1pFJoG5XhAnscqKMOU0GkxVnVUIsC1QNkAfamD3WCGGv
K5JchjMWnjbRiNr0tY3dOo1ei596WvB3daiovIRQCMfM4i4Ry75TLrEXMDL79hgikJm7pCwj5q2+
C68Iveh6f/4e4QXQUvP/DVEr2QZN/PUlMwJ8Dk5++czWzhDd/socdQNrXPzc5aOvaTHZU2lCoNZ4
CH3kw1iZ5+vHVgLr1hxgLbKVhy2LpsoxbMesnCPFyyfsTFBxgFy6S9fX1xsp0hui09niyppOlUvW
6P93IS2K5uPIyJeLgdOWioF3FTzpcMCqUZDQ5lMQtwidDoA2pC1My2X6jaEPub+qzDU9VDiF7J60
eQw22y7pYu/cEOmTP/EyPQB7as3tqHHSWUePOHFZEJeKTePH0FYdzgfEb2FLmBvVg1G5cnoePKIJ
3uBIAPVjW6kHhZLToRUDKLq90wIX9arbdAaRf1UlcOFUwborfPGdoWHYw8OtBz4BjzwhAxrHibJ8
nxu8OpAkxONDbx/Q34AmD4yJD2Ee6bc6NP6qRn8Cbyqy+3p07j4O3Aofn6Ti/XiGdKLGqmFA7Q7b
ew30muF8Rq6QUJWhSvHSMX03xktn02XmgvbEJTHf3XMmAxVl6TPvBKqUBeNNis0dSLRDMspYZusk
fIHVHYGNe9TFy4kU54jmfrQJxXHLWkE+E/KkRmHPmbDSoySvjGmNidQ6xsagzt/FuWHFIcjhetud
3JtWztet3lLCkz24Xya2fZFzSdjEHskK3tODQoG3+F3eten9YeS54RQMLaPnppfVJH6DXaqcN2Yc
Gyw9Le5m0zhGV+aVoYeILiTRddKLXpCY+qnm+JWmJ3mt9P2N4vvLkNcNDeV15gyJN3bHR6bG215d
RgcN/M6XdiEXvd9CPLKZ7aHFo5reBUDQeFk4GFQZnw3YRwHVAj2n2tu1rnkQehoY3/rcaz8i+iR6
s9qp3gtVzGphHnCU122eenFHOp4yY2PX2hIFYzQw6zlAIJseJezpNzvO6hUT6BJDxE+8PastpkbH
o5qXTuvHe7i3jX03kkPnD+s274XUyn7/Mn5hUQnpAyDgGLCe8jP/JIhvyOuVHh74rbQEd+aETXJa
43z1DMZrBe9tTl1MjS+JwPsRh1j/kkkx1u9gHjYmpHQyZGF1pA1ToAYApPOPNiKtJBATas+tcZ9K
uO8DX6V7xcJQ45D+X4we06DSAYg2Xkyt/+mUWa1130bJVzUDVB3aCfLJRi3/r+lsarxFBMqFWIh+
JGjOM4PoMhlIjqXGICi255uz4iwYMFV+L002geKD6V/jP3nUUdL5+o7Yjluo5mAKSR/H1aKp265B
Bt+Lx7TAQrnwHyJF7yUpNQlGxc5sEqOTSYAoRItbuaHxHOiRiIrOc2FUfQStbWpOnbowpxwuxVzS
qjE0KLhTS7WQfeHFcn14s7JeNCFpEzDU/OYaunu7DP2Yqy+ih0zkwtZ3cc10LRQ5ec32rG9mpfBC
npUbc9CMYK1lcOQIi5jlrUQDwKIHH+8iWm/z1NkLFvtK/L9rKauazfSd0bcpsX+0o5fJP4DMPGT3
sJmN6K8eRr6K/OQ3aJPrrVHWyCG4ca3upLv23ACJUmnXEzjZNb6+OH8A6u0nIHKD9gxXMTVRxXvY
b+0cbTSPfJmCQWNByh/fHOPa5jqd9NNL6kRmSASCZFJMC4W90Q5lmx4ZEyXuXu4zEG2X3WTeKR2w
KCD4z2/nBabcntNTGTu146Zy8Zyt6E+Ctf2i3aHY4iHpWGn2NxzaK8U5UwYQPVO1afXtCrgF7A6e
JNyxD5DeVKe4Bh53jMk2FTdeadOKa32JU8PlX/hht97LB1lMGbRBLseuxTw1j3WEmOrJCfTMAhKK
GDdbgRH41iRTO0tB56SkDNKOAFwrJ8dHqAQMb2bjZ3ocVsT1cn+xNlVyVVBPS6Rlgv2WavuJyM6H
PSTjwWp3buX5bVbyS6Jd+9l8Ur9moxUIx7Ha0Tvi2ELNkA6gPGBtA1udm+nNuP+4K1P1Lvt4SnSQ
RiKJYjFtJ7e6nSl357cDZv1RVRZI1IFmUbCXaZAIf3s1bIjf9iEJnOZHrDPGSzggfetR9Ni+jmok
wJfZwDGLVYeAaD00PJexeC2V6MYX7NwHpX1XzYgI0XKcQX7CCBp7N1u4vrLWtBkcw+hSgNbcbKaK
9U6VnbpBO7Q6UAYpNd9C06fc1d5c2SMFQ/bRnHrJDVBAUP6OVPubhhgYaewBxA0C1QGW2cHh5BcP
Cw/XkmGfkq7+BGjOfmqT7us/hWu1U8YGmtjoiCHBACna5NNm4VVv5gm5pvrYuQ/akw1XJLrQBvl7
bLlZWUXoBXF7OShzDC1ye73LWXuzGQ7PFe0EUSnBrjJqfWBWed2Zr3f8O8fqc9Vt5gYIWPmlOXNq
Cd82+cyhriQw0/eN2hLu1WhD4n0CO/NAFYj4tcuMgyxHIdyxueE54s70O1Cr+uaXz4Ez8mNg7AM3
YlKKEzqKSUEe9iknw9zPovIrhD8FlTmSZIgL7PwuvPcCOGUHVfBtkqA5pXzZxp57G0HveT1NA/1G
TODRwxxPd1MRy6W7v9W0rAgMEYl0NBxtJpcL1CdqGn2TUMhfSbqfnHbu1TLP2gseWBlSlbQaUz5u
kxrwVn1YjMmqOTLAMJ6bZzxcdOc7W0YFWZQfuCICQdFPsaB94zdoAf3Ufssy4LJ8zGpwid1dG0e9
wpYCn1q7sdFvf+DFDIbjJB7/hNgUhiMFUCpkinMBAazHJKb4pvJN9pHZBc/Gk0V6Qa9qV1jf6XEf
P7qQpiKuN3Z9AucogPdlsSokMY76hOXa8+49y6S6xRonhlL5QmGaZQavYfd4eV/89OBRfeeOfVdc
0B3zFwD4fYsjGuKp4sML+/NQjO4DlHlOXlAni3wMhXoXDkvEogvan7VXHN/Hs3mh4q72/k+RCrHn
yyZZUUThnI6msxKgS0VDJTUMfHMiqzNAVj7Tz6O33HucGaZsmalgk8FcernHWktM4X12Acpi+x/c
N7dBfvvIZT7PMG+10oX0qkBiH8BjpSDKbNKcy51d0tecbAXSpus3Ij0k85zbHs8OClj0r6TrpQeq
ZGxDKxbpyjFWpyMrX7EkpESu+y1YY/hyv8XiHfsElPaPOnlO9LVY5pF7VxLB2aXjsdwPyq5eWSwp
aIaG9WTri41qAtYtMRWyB0Ie9UeAcqy3+AyFlEYB0OGemIyIq3V1RoUhOl0R00dZWojsw3oD0w+r
yz3Zil6Yo3p+FBJbJ9ftg03ysRU6bPrGsbCd4fTOCk2xcV5+X+pjtnRQOly9pBiRX7RKecVGLfJO
NanMzCHO7kVKSjhxEDO7hyttrmeZRaqbkbyOGiOtF4Wv8bwOEZX4yyZ681V9tw/sIDiR1HTOlHXP
2id+WeFP7XXxUvEjV3rtvPmxRJFH4XT+MBv8/ptxYE7jiUPG+Lx5WFOG9p2qT6WJulIWgE46nA2b
kCOduhWQFwX+Eb9aTM8O20gc49C5nDM5npISDusfg3CMQpWAr5CEa3Aat+cUeyMwsa+1SW4oksA0
vT0CT/rM2AYO3B9ol1SpyBgilZB82AkT9Fa9IijB7HjPSs0B5xYwm9W22EZhleHQSOzxAfc59Ecj
4QRO/gZEfvFPzyg+9YMYmV7p/aX/QVh+n19eWxjm8jK2bNnFivrM+vBADZ6Hnp1cPYTsSYf9ZKWH
bHTTpHpTR6Utwf/A174/oOT1rpnYYqQkyDueId2dZMFcqRJJkt2K2PmwjNRJTtON5d9lti+NPwot
+o/GhWzCsNzG/y5UyY5DLzICOQPEjlzhhT5NNQAIS15Q13lZQDlXAY5xLjxuqa/2gI/KiGgF1hvm
5l435zLytQtjUapKM99FtCj5psUggwk+NAOIB9eK4G8xCmz+RwjYDd0uNPxZpiBmVD69lAlNcI3P
p9pgYFIcx6bc3fRtGpn4iK/LPSD4ELPZ/Bzb0pTijWmIOETjIqj7qDyCdimeDwiWdS3eWNmqeE3i
SJ3hVSpxhJwHWA7JrfNYEiV76PqHWskpgb69PfEX+M7YnSBiBLunrfyWWyV/yhBuIksLEUGseHSL
ZXOVCYhUbVIWy9wrihjkSEQPQ0TE6H6dWjNxOtgjysI1DLyustOG+n0emHvCpU+/dT2MgnnMhj+1
vG/fk0AiYNzk2kcyxLDI55ha9B4C68F7RMtw5KQiipI0uKkVxHVJ13CjwZqoEtbRs94cZwBzo9Zf
cm5yYDGhM6dTECfzRnRkhAkoW34i1aiNrOcpyVy0Uckv4r4Mvd5iJbRgQ7NgC0eQ11rw4xwxHavn
dM/SZMvFEkLvDakl6MJOqjfZW8747EYn2RpdBvOk+SYGzoov46zrOwmK7g7bwXar0hrqimqJeI+3
dWU4eN79+2iicQqc/lxM/afmrigTHiavB8ATy8UjIDh1tMPlXVGCo+PlTv9qIiK/MUluuKahTtva
bFfClEJyxHB4lKRzemIAKGCTWfc+BXjFc/cYLnJzOEqiVFrL279DYOmbkFkCOzqAPnzysmmtrxC6
bFSqGI9Qq+sTiPNObm5QdrEa8LuZnW+jkYNICgueF9lk1BKxnX8k9vZ54B5NrdKWPMYPH92Cs/ze
qlL/CdkQiXXVIa9jIAJqe/tlGEicpMT+7xQwtz9DrjgpfRwsNz2AAia9/uolY1vcM4csn4wl/ic0
nSQ2UmdOMYKjIEas6Y8QL3H8BVnrOm1X1AmHZC4Lm7rcsXYtWN5sowrDNbwwC+vnRJFiEDdbnZPF
2WIqadLJO4LSjEgQvjdnsHMcq3D8GBacVF0PlRoOWLjSUNaUzmNg37PX4Uf241Wbl7smrYnZz2jN
RobLZZZC++5XB7kb1Sq90plB+e9ca5ahrHRyRZcfpIuVyucbodgJLNh9aMOWISfj4vAqyv4lyUl+
eVpdLMKRetop5lGsLLhfYubr5ks8/6751PGSwWVxAXmJ84/501q8VPaxCerj/HqbfCDlopbNagw6
zUBvu/gX+mvKXVPx3kJBX5FerRK1U7avKszlvarZmwOlGqUjIXxl8LAE8HLVFsnkrPdVe8qj0lcZ
+YlXEcogC8rBahdnUFDLIcbkM0xNZgkrugHxhOLKum070YGJG5yIM1yyfUCxWCbM6fewbC2/wmnX
G/QTfejSsD5BU8lS94CG6CsIeMzVSZqen3QkZIm1EB2Jt0cjt/UD19MbXVzxM+9zLFCrQWrQOsLD
fc7tJbx5iNJ/qhLwa0yUahmCEXXwwa8C84BIPHG9Xkd2/mJzEGam8Jq48UpQ6xSSt9D4i0UvYWDa
pjbZqJSXvISUkq+w7nrolgzDeVoG+pU3sOVcmKSZMvUr+LSUsUGwtqbdYs+hMJdGSO1Qul73/DZW
vfXrh52SG+EbyykbBrnvE9XbpH4gSJ+xdGGzttCJT+g8cDKMs9lnn9GjMwOTKIL6ARv8ovXBckjc
EEP0+MST+VvuKknyvHzea2SmKoJAjUyC2Dsm1fg/ewO+0nljOEK+nMlqLSXN0LTn+W1moAqxlkwA
wy9XCV5QEE5lviJ8yfynZto0kITq3EEhozSIRal/oYSM1svC6mKh+5NnhSHwdI/Ct5u+IOat5kwx
f17vqRM9iheYASNdntgXaX93v2uwie3I8EiDnuXklEhd24Fqen9iTw/KtId6xMDzqKWquMyhnhgu
WykvzVcJOE3ruiYAiblPsljLfPbEqKV0VlOS8a/vYUNeVsKciCAHgGzhUNdEvlbghLdF7PFh1KOE
Bka/1WxUsRI67GXI2sOqNSXpfOLlp97rGdzrijS9vmyLrMtYjyItJTFRB0L40ks2mTi62yxwrd8E
7Q0tXTHrLchxA9HFOqGrTu/IynQkAGzqUU5qx0pH2CH1TdpFxrma8W9WisseQrEg6h9JEDWgNpay
LlnwpcKJ9fzeGkf1UEQ4fc9kInbFzr2RdwHML9+e8C/kLq+bOuAomS+dhzMF4mR8A0c6MeQteDoY
8rnystTaRPYUVjOo7+/OPaV0IY0NOCXjhv5L2ZBDtHs93CfTzH8UeC4GfGPh3Hlri49CHjB1ZUxp
EnCsQkq8ZinrAXl0Q7iiOdQkoyflYxN40niEMKyun9yWm17jGz/8JrnYDgioMaE4U8Jo0oRJ6Few
pvYrkP3ijJZlLsBk3W2dNx8/IyGqBWwCJnCXUTlwLlUzBLSKeW6i1t2UDX6bVeZ5xNzwlwL6IRDr
4XdShBiiubBzHStRHltDYVqhoubb9W1MlqSuPaqWx/H9mv/b7EnGk5Om/lbb0lYGxlV4VgrfddS9
j0mSMi0vLlMNCUVdbAbZvKhlEjdt0GL98JS5aTswHIJF+mlqlpAhJj9+GqbjrXUECOBXwE8Yxwmm
Cr5x9Cw7+0/WS79RgsBg/Yx+z9Dzx/cKGKNVUVunHcgMa1ks6jqUaT2JjMUn6ZMxwlUXSsFzOFqN
qv2xlIyBRUulS4b/hBJ4HlagSPEpzpKB5YTr9gerPbWkiAXB/J2wReMT8BJ7Xeew68l8YRLuXPkk
BQq72MbOQpTqGvMA1cdwEkRapqqvONwqohjCRmn3a/oSnGLdnrye2c+QmcM1nWDRSXCmZ8lF8zV+
YchIl2WUQBcHklaZoJIG7a1zXra2rzussfgJDIFHAa3/FFLMm+a+Lx1stW/tpvi7YNkmYvFCZG2E
Oz8JfEgfo6L4l6ciDIi25woWuVbFzVElSVrBWsWkF7KKJTRoWyMrJhSn7eCvScTwig3sSXO16JOs
mfzkPpw852oij0LdzIT+KxsWJdBPVxXQcTHa1AKu7lG1YGPtWr3CpByq+n1Zy5YgXENqj6aMgiHQ
kHdA4bOmFLgSGK+pqKMblzjhrZkB8gusnmfPWBqL+BizziTT1j5OfchBFKdemxZanFdTtvndmn3w
RTXRFZlEMbEAfLCM0BWvkUgYTwd21MG80HEyfwX2XxRFlGkSLqMwt+s+yQcwqr4F62+RGRAY7sNw
QnAWvYOQX4JFbx+FzH16rw4/f3GluGV9DfGUN/aRulwIibO/zil3QE+Vh3kLBtvqxDJyq2A7e48U
HaYMP3J7koysUVZ+qXxZ7jAgWKhhglqhCWSxmy+Dps+4+fvDML261Zm9+AOKwXu5DFSUU2lGN3eW
46o0nFiad+C+HUmXuK5hD4voZobY6pFRWQZyQeOeTqc5ua7HnSLR3hwzngzoLvyjNKmAB7VyOXBR
1Y6o4p5qd8rqfekMUkEDqrWFI4LN4Tdt1OWjCoIpY96QcDVcu5FUWT8VJuBsVHkB2DqoF21mpmbD
fS00R3JSTGb1QG0a/gzysTJqTq8oMCr3Az7SvMLZqvryUFsixje9DQeeVg24HSSE2sQw3g6KnPYn
DHXz8V9+051smbG2Lt3h8+Pte1OD2OPInS+I43Etw8vxrqKzaq1Y1tYUAM2f9tYQ/8OM24AiTciT
d0UHI6hT+YLiou3dzgyuLtoCTTCQwFb3tFXwO1D/EzRJxPp6hlcKgV/twQthlM7ND4igSaB4J2Ph
/2wRhNyhtxSrkXyQmEm8BBodCGti+JAGFKlZqnNrnEDo11awck4KPf1kRFSXSmu0iwTrOVqAc/5j
zmjEZB6AQe8Ukahm3+CVodJIdsyMp1M3dmdc/Qo4zULtySjNTFlVGl3Kb/B9jY0FLOfwl0AZlk04
Fd7cc6/N5tGe0kJjI0fD5RdYMiA2WisP4W6aMUN0TTrYgYZJoXTa66pE/yUTwUANuefqnTjmMlaM
d4bDQipTgVBseJ6Zzd0MeQquUtF+Vb68zPK/e+bWk5q9x5od6FvYWLSYJz1VPS4r0/i09um+YwFk
o5FQMKB9s0A4JwZyEI4nZzif9+AiszXcARHNvvESjdv/sieKwb0PyThIF+o/hA/ycRGfpSSgZ3WN
T4uyMT6T2CY7ywxP5XBZil42Fy8bdpfhuofb05EG/FC9varuFPVJ0VoiRf/zH1GAgiedtO5qfKDm
U89yJt2Z786ziahfzHxqpJvYApFyHpJru56aVGbAH++kdvDF6MX1UtLspZoZcTfjWoPuXuoyQZCx
Cp+kPASEH2Fd1SuMx61Py6ThuxqxOtXaPsLO7QDAhC+K3J1k41UtM8UD6d9SJAb5symiafyJhyk7
ZsUZ3LKbRG2E1ZB5+dJcpvtERajz/fpMuP5cEEUZX8ozTQEqi2RMzddymQ0pIwdupY5eqaRk1Nrn
RYuyfWwN+NKg4mVCz437SvjrqrlETMdsFcjo4AEipRtmFuVKyPCcJevrUDKX9xJCeo5H6aLA/d7x
dnfombUFC88iFcTy76vYhOjD0IbbtQKl+zEfGhW3ZsN/IYyFmEa9Uw+vMXlQpC6UFhMAuLaHkJPL
VwNtYebt1wtEx0OVLlZOidUBSPCKfFSEAafezZwNVE8ChoZJHJUhUDBoOAsomXIgWfKpAs6FPB88
LHg96y5mmrpdXac1PjToC2aDH4U1pZcn7DkToHxaY0aGWcYNPlMeNVFSOjCgUJzWBd+VtPtxuy/s
Mc7KzTLclGzh2c0/UqilHVBSFGVTxNpwp1ToN4QN6RSOcRZTeCI1DO2wZ6tqVgjGiiAddAKM/jo5
Xjt56kStEKB6JeTD8eVvxSLVPb/NUgzaunbXuQVd/OC3yRlwHy0jj8JaW+PpN5dgxo//KQFZCqZN
AizXxknBrv3KG9szK/l/Ff3yVAQi3n5Aj1tgXj/E7PIBCK9sLLN59ICIyZ/kzb5qeSR9AGdbiMPR
ubxH0AoGvCc2jX52VXxglHqM/7Dl3Gjvk6FusGdFl5q97MWwWOFAQbbuyReNe4aeLWaeL7E04lwG
x/IRqyDw2c18KATUoKfw1ln+uY+NBQRHdpmo79hZNPxSg9UC3M1lxxbN1Yh5iVvla1MIRYGjo3YQ
oKMZZoQ3ZX+0GZgvWkZG280MpNKy6eADNtpeTz6seKxmXM0niJMlHnTP+1lplA1Mq3QgNrc+oDUZ
f9xGeWAuTyo9vrgJqEGoZI3vP2iF9dGaYnF/V6m5bQ1+NtQ+4Rnwh3oe6V1f+SfLmqv1vq8yDb0b
F3cIzt6f3E/7NQpomltt89RZYDu5h5SuSk7ogib8hZUzYE8nJH6tdoIl5YCcyRe8rE2Kl9QTPjhP
qFvxP7y2FB9X0J6MsuUYW5kXuWlCSHsPrJXPPhQSyd++AS31DvVb4p+O6tqDvZTZT+n58R9N/wfS
knBykgO4P8z5OYASeDbO/VnFCggqu8fVtWuob9KJa7M+EP5GeX3UHgqjTA1m7Ddc56P7JCQCMPng
35MXdfHf3cYPIEX7kdTnmJvEgL0HEnEa1u/EL92M6CNQiceBzWYhJKEY3sPUD9xDCJytvsyRQI3x
OzNAwwPzsFd7/9ZvpA8W/+bm5Xc7UVNCCUVbgswBy2lMVbHnHbIXTOfGsHYmN19EquHzNsFuvHur
1hVEEwGboVqRZZ/E1UIRcyEQSq90cQFthVI0qfVjMtUKjQ6KwTbNFDCl5d2w+hlFlbgV3gPibIVD
/0iQwSVC11BNENQIaihrRlfDZAeBdNG+/1onWXfe+QmF6cUBwNyGcTllKNAl3WIyRXheAUOu13sb
5IKmeb16jmmqV9qkYdCAIQO9tZkLLJZOram83wrUeX+sX/YAAOukYc5JkwhF0jkmviLckpJomRRl
XmKjHB1XEtFgJYVWZo4vZhF6f7pibLmIkRJrEw8t5lEOXim7zoOumdyPpBv+TLaOOY81j4ovpX3T
iKz/VNIFhoVs1aoq5BfWpWsX5UdEHBjKnYRg7uzeHxeSjKAql2PeIqdZCQa2iaAmhWnsTpTJ/faL
UWQ9akxLx+Ueg1mKh5RDU2fRoWzc2mFlfFE7efrYsvo/Cu+w+d8JWgs2Eet4em0OT2vQGo5Ium6D
0kplBtxSD0zGmalxNtxKJsAmNDJmDOJEwQl+aIptknhswir83RIYyENtax1z4ZmpqvXmzopuZe2l
0vsa2QncpPCYEm4DyoqvFm+XKLexqM0sSUnTVqbRD/IFw9VT2yqUm1SO2HYa3t+4Fo4STj2eORpW
xgTG1oTkFvKtnNjHvAHoenByXaiBpCvdZKGT0D77PyVPC5Q9O2VLcdPjfMckKArn56tpgirIN5Bv
MfJD7ChiR/HsMReObgKt7BDBulfEDqvifXSuLDL1DmD3lADVh2PCRQ3wGRz+7UY2OLzhEwUGgQrb
haMXUKotN+lbMQh+866AJGQxfoku7pNnSmC2pSY3J8u7gN6PwGm6NChttQKj3m5moExfnm9uvEUM
eqemxJnyURvz3tooUH731QNS5tW6ZV24M5NgjBoSihpFxdyVNRlMt8WUKOJVTS+vZxXbC/dtml7H
IlfThIiVV0ZWlQHyqekISuEjOwp6S+BQhYnCn+sGglUCfTX9jlKAA/V41NN1UVVRQZeH6eSI/izX
fbp8X6FW/TcxH+D80zPyXZYtplwXqsCNwSWRbf8jmdZ3ggbphMnqz9aol0X/11b7ePwMFcMAvda0
4rh5P4sWp96RR/9fZ6sxeLd5FytBaL6YFtEq2E5N46LCEneZRNUUB40WhSqIATlG2PFGSixOtI2i
H1mpr3au3YAc8Ha1OQrdLJkeGYMEA0g++VJIwACt/5EjDnkzLpEAsaSET9U4AFr3GRlJxYM+bTmB
cTKUq23tMrVSVDt46qVPLW4KHBRTLre7HPtAyduCljl/CJUTZDFXgsaOPfDY2X6XfIAs244zZRRU
o44UJTYJ7YQfmeIsUOVjIwkfArx1CAN9LP/zy0i8RxgqjYZIdzbzHhfOKObmA57hpU2/SWjBwpgM
dRs6oliCZEJSSc8DkQHRHgNpGPdYEQp2zfA/WqPDXZftKs/JNFlMvZvBr9YOoz29o/ok8kZ/BaNm
BM/0GI6384MG7fu6JOpm5VAyRR+tD77yt7zLD6s4EiKECX9l1Tgh4XDr8Kechs4VsQrfrmGFFDOC
SB1D2CU/QhZ9aW1pKNleD27BpX3YNPazuSirS/UyuT0sirAIHG6q0Dp7b4MSxEEtcCriW4o8oYqN
f6hOcsYzSZcJW/0aMDWJvEs854Ca+8va7qv/SDFdPu9jdFg+qoOjG9D75VbrWapm2q2ajADfz1Bl
OYAQFmbJPY8I0Lq7J8R5CSo8yqZZXX9omc3/EsAVlRTs1Htm/i+CJvUw/b1FLy34lOsQqiHTP4T5
3IyKZnwOoTOJ1GwV8YfsEmR4OZzuD+UvVfT74X6vk2nFa8Hhri55GhyPGYcc1Dbp5Y4i+b48VKGE
qw/ByE3c4hptpZoHREU6xXsYJsyHNMc+nfgt4kQtaSv+YJvvGXKsIRpen7sxR1Zx5z6nJyl/OKzH
sWo79hPnu4bXWeNUX/x0x90xY/3q9wKgkJ881KXQbRW2brH+DZesoiR3VvuTCvVPlU007pC+ZcpN
bsik1cSmWTx0db7qUWqIV6TJMHdbHq+WNtR6cc2Ynu3Z3aQ3k2ksMs1Yre/iqY6u2i53H1awrJFe
reI9v/NPCRiaN3gQvNvwIXu+UOvRbz9yjRs/+B+8O/dLrv7EH4+7h17m2NwOrb8FMzmYaa3XpO04
mIKZxY5TWplk8yQH6X2Y4JlUzxlxcRfaL6iyxLWaLLr+sTrjs04O1yAFI/zw5g6F0QUsvd/2V6og
mPXzmLhxDGG55xsozfyfyN06qkhsynV4g8LDK3OcyygWUrgvWm+QaooXeAUqrGGy/oQBdkFcB/wn
gwavvrqGN6JEohILoutfRL9zp7v4G/i/y6XAav7GQmrsfA5QBjnXeZOcCO2gd+TZD7RljaZm6PiX
cGWCE2EYcD4Zc5Otu/zlkZx1IwxE7HSfE3vf3OkkDopHNKuxtY8U8t/65D1mTe+K1dXYlL7dijue
M5/QTWYTb1NR2BDtjw29kr9eEiLjdjIhwRRIU8b7bVAWdGvNqD/AUN3M2bD7bS7bwAuwkSQK9kBh
cfF6lw+9/E1asXOt3ToZPv5Mtyu7CKjBXuh6DjdAlosKnHd1etRn2MH+w7GeGFvo20h2iH0Z466U
kGeH9ZF58l1BHg1MdnI9IPvg2mlw+nNKjf2w4IZN9lK6V0VraK29r7vZNQPrE9L6Lv8xLO5zqfW9
7C2i4QMzBkyfrd3LRkB0kBsli8s3745HxtmLmLsJ8E5l2UaWX9L6xpItMV0oZs5Ej4gQ1zOsqHOu
7a0gdjXsGoxEMqaSsvHpXBiWTdUkt7z+1PAHVA/XnyCziKaEp/TpzTuOvfKY9yk21l6+ElMptCS6
xCKHGbG7QgAVeU58tpz2uGHuywg5fB9d2pB/5Dl+gc37AhpVPVcrQLjrz0vvw1ik4lwq1I5PIpQY
XyTrfJlLiNT2gEnEjQccYcNY4G2VYqvHAlxok6znxjseTM+RSeqAvsuhIcsGWyxRKq+52JL4YP4p
5km3iz+ID9POQCkF+E9BhlHUA/6hLEUN5UWsynw2anxPPrPQqCCiCRET4aTiMIoANNLSjMkv5vO7
M/WizSrguNYXoT8ITT5vRuMeAuuUyJjjfaqPZTIEhVaYib0SKxBKTGaqTiI503S23OKurlsEJpty
FKMhVfdAKELB7o+PWTGYvv/Bxc+0II+bQStVFNW0Pm5qXHIqCS74jpBtepC9P7du/oDvzzKmdLff
GFQUcxw4cHIpxUaiUotgDjYmvldH0aY5V9sK0C88eEiG0PAG4G2PQZNUkmSroielNpI7SCAWX/Fe
XFBw8cL2vCpLtqpmhla6o0jlhF++N8ZaBxzhYx+RYt0cnycZEO2Bn8JD0sTMCZN8gyZBrJEH3/CL
ks7QTBjd3hJcNdEWWWWMMsG6Pv6kow08hssoOkcmmSyYoIB8pLa6x8m8T1s4efy9+vvD0c5Fs6pH
TAoOxKKLpMl5B0v+61Y7XGBdAqidsmcyDJ0zqnrbq02fiXtU0X5j4YnFGlVGBDuo8LOM8q4cjy8E
+NOTtJzeV64PVqEWHxuiVgvTrQjux8GAmeMOKldpYM/KZYkVEjgCBQRIWyXFZZEmoteAtGiwU4z+
r5UgDJqM06BpOfYU+CjH47sc/JXW2VvuPp2sTtU3DqGS7cjOXpZblUDaMkDqFF1WZ3KzfzHzFZJa
AUiDg8pfj3s4kN2XCKbw4OA5OUqXt26OSxMRJTv4FhgtlvzCqjvzNBXjs8vqTi3GN+cT5/CW+Dv1
QReeemZJk/dCPdssyIl/f0qUDUdkANRg0VKeFwt/e4i0Drg+L8qiyULEIyjMVqkyXD22LKNNO7SS
1DvP/4emTcS8YLB9FCJFXd2t8oVwVjgGzHpi+K6DI+VZcB3S5EYKYtyyPnqPUxx2nA9qqbcoUO+j
lXlBF2N051vEiabx+EHz5ebFAclOhCDMB4+8N9y4d+RWuKCoVw9oTnRdCXr16udoF2Iui06CEFZz
j3wvmSOZQq6BRZBikzlR5wegU6t4gQ3rrykNK4Ccm8HewRXCzIN0885HKLE9bjqiGPFl/4a2t/9u
gonFtwz9W3y3olcXja2HeIdxA5FwhnGuoLYLiGcjV+3NtDTTTTO5+yGuY3mGWvRgWGzLMhhCWa3e
jLlgKaxfWZkU5T/hhokvnnXo1m911opQF6Kt6i13OqIz33aU9zsx1TmExVTF5nKkfqx9dS5sMupI
5oN7O2GYxLyDT7wlKqRtPDehFb3FH/YJyYswlX8Ym9+PIKSvkhghRDAKtsbsFQkC5kBOnyt2ZN5y
UqFitzWYLKej6TtwojSp3kzQsM9suaceoCFUaaBtowwF9d6MpgMj7plaS+QJlDDDxr4zoCfcOHwI
UJ6AII7MVqLBhs3A4e+7ce0q0MgCi0tRGqluGL+IkV9Ot23Ls469qXW1jRuUb36QAH1k58MDyDy9
Vr6GvCyfD9GPDCicO0iJaiQMsptqmPiLG2sb6y8/HMiIXy0Ixa7fUxNeUKGu4czpYi7FzvJp0WAL
AUgXy0kXTHKWBqMLODEstzrMrLlVCc1J0QSHaOftgZC2R76HelnhCMwPkkkOiY9F92WP2UHGYXQV
wxAbGN6pw4E1l5//6uR6UF71feGph964lucuXM9GNEqOIptqjqUWILaAyR0iKEzipPA7A9deYQhN
qvdbYqBfaWc7vDgV5S95TsTcT82DmfXh2bdqlVutA/O//vprecj/K/PT2iM0ab7C0tc+I9S6y9m3
9JF7jFLJB/8jtPmGA/4BglEcAQjiPwLKSzmbZJzUbuRRpL2M8MxyMSpfxKOGLdweu73AUMr2QuA5
2rk2k6efyZU87FWlg9U0zWgwUqmuZvrkM7CRULeQKdDgs7nYUjmKUSWQmzj72xkZRKjxFRhZF1mk
51dEEZCqR7LIMlM0e1EGKfM3GZ9HmtlPTrSwC9d78Cym+csylH2V6CjklhvKE1VOD5+a08vrkS21
SUnnGiw8PW/uDfHkElD/EIPV+ZjYkvKcadfc9NxHKs97LAd5S31co9H8QqwrHvUE29KmgMFfWrw6
KrzKDtPnvl5GXAeKQNd+IKmpFBUpPY/LYIDaKti0HVuREJl9q1ezoKI3eVp5AUOjpZwG0R23+MZS
DDAkW9LaEIwNox7D5AH3ocVOsbBLgdUA3rArxaemINtyG126SpXarNW0g8nbr+2eT/J7hDjszZjP
7USbW53k8Y9vPgIaLYpwWzi0I93NKhPglFlUh6w4e0DNpL25Ps6m91HmKSTzNJAl4TX49P/Hq7t3
OlPrKq5QI3ynhz9R7eNPZoVvYvj9edgRMhlHDiUWmurZrLglLKaSsBHDxrnJRkC18s7iP/7AB3s5
CLHeCpEyTTd0srTvOgjQfmTQRg5jNA/hHHddBL3HpRrGSGejjXIQxjraShKfArcNud3YMHPe44Ip
5xtMl9MSU1WmuwvMKST1WE/ajKaweZ45WCwipMN3l/zc8FQJJpNt5BUOXTHtDL+8/HV6i2LiKgEp
III5MPV8HIi71ZW4w36ay551SFt6TqNzK3W5ffpC8tloE7SB2kel13BGUgBDRIkVoLQ7qyGqdDPL
sSIWwlEVsBCcKrzceCnpQ/nSxmGfhwajSkMN8hF76wtynX2jv2MwwPEA59RSBk/KfQiu+XlBFn5v
mTBMsdebvE5ppM1g9OZg2cxSBpDIF9Sk+sxLoNT+kFVlKv+iuAUk194yA3SVw+Cuo4W1yGcvQOn4
j1sQovaHLP3SH6MylKzAgPvmlacnfICAMh5CkPI092uLDHSwC5h5giKTR8RgTyfIx4hCM9Vg7aUV
byJY4y00IUY/00vm0qn1MP47JjhopT3F9b9jqVfkIjVx5b1+HMhT78Fo0Bvqs6y6QBGfhzEtvy6f
TtNYCIYPC8I0heR+evqL7b1T6wbExwJXZc+ihium6duepfFyPpzooWzanC4qmfrM2TtLPZJ8Qi3R
OyDxCLd9gzrWbGBvpQSQ1Z/u+LR3MphPOhg4PDG/VvtaUduW5K+++gkEoCTV35CfFFjN4gVSH61u
lWXdkuB5kX3TX83dW8Gn4C/qaPiXGpBr7jwz3MAY6p4+FmZO5eMYIwUmBg67cQ6W3dWe8ARuQjSh
YULdZqqgvwh99Yd4/doZaGsfa3kiQsg4AXF3V8/O3xCkfQAjauPEGOc20WHdYUihsvMXmQU+YfRj
uX/uXPnfLjVTaXjFm9i8UtTsq4klk36j8HhrNj/sl5/LcQPhKEhHpgWv82vu8gT8gjt79+SK6sDo
jhieC7N1VlzoiG6umM32pWF8N+IQsUoobtnRn+BeqVDUTaXLnx5YvGRKVnXLoOXDHtU4PxSBwkM+
fY33YXXUZ2idV/CK0uKwKiKogRgp2uksoRYlTUObHR2zQNphzha9h2WVSgc5f7PctRHZAGKq6veE
+Z9MiiRH0WhsqdL1wheBMDRxCqTva/8cHKxh35kg0MwL/7BrTdUywLqEaX4/B9qUCcj9pRCozO0z
9z5SyJnE181FRNhaEMAtnWWHXkdbS15Konyzg9j6PgeqN74nh6z0Qvzrj5Tv1Nvam/LI6QX9K9fT
hUrmUjyfCzCS1qK8KOQTo5lhyCylAZ0Xt6aBFtsNChoKZIuGOuSECUlrTUEma1/SUiF6+oPXjd2T
Gd8YOdizw2ECnD3iVwRpUBWzY8906EIbaWbmB57+Kfaal84dHITVyfY46XD5Xw4QWC0ajl3fu+tg
nZ/zjFM2T+pStFNzFsOyMzv6sraN/8lT07dXn9NgpsqcBJsNSS0skczbVDubz3E5yyiyLxICHHm4
7+C+PNRUDNDrIEkFaiRM7qQsRBMNr6MfxMu31L0PXTMnnPRSm7HKr4UzgBQaUzz/02xNLVaiMh3q
SIZZnFTLFBX/a8VuIyrhIcoJgHF/8JbdcWqjVzE47Jk/WlVgo1hYjB+RqeE4ELsjXLid6BuNVfid
OUDHgOibgUtFRnYlmz+EEC/PFDsGVxW/zVQegOL86xB1LMPjtBkA27FL465Wwk3cDwjixHfsuZHL
r0pAY+2LI1rANzCkgzfIJ9CReiRtpIrQOP10LAjeNwplBcIvqm44swaYveNmmvzX/B188xosdcZN
fl9A3tyzxj3v7C97K0UpyhFzgIjphkjTH1a/9/PoeeI0x0W2vT5ASqQBrPUl4Isogrk6jlXpXYY7
7COdiwzSSW5sxTVxSEswbUE6PYZyKdPT2S25q0EIu9KrJsVx6FmR52S0U7dxKq6WGLlRU3w8Wl1x
qWMwe3QMesEYBrhfPfx2YxspGyFAVy8CTNmDWclW1r5qlJHeKAlYPCn44tL6B2G8R8dt91bRTX9S
d4O2AvIxcc0zD1AEFhYc3ThR1qQxnkLmQIBwuVSSkpYEAT7beEpJ/x/FGc33LeaOQPLoQzggXPRK
55Li4K22HlwI5sWHEDG3+4312Mhy2vQV1S+UOQmgQvnlOo51CpFSJhTkmYlCI/XoxoIV/gossDp+
Sjmqn460mROLGjLJHngEpFpB7MUKF0W+CLdASI0+Of1ikmtrvHQ8I1h51K642YKd1IFrodA0SI/L
JwAc1hdlThCY9CUKDwTY5p0WaeH7BclQXilVFdOsNfo0LqSBZUOIycVI4NwoDXgoiw/AOrwyt1Qm
wxIWZguc9PW1v7IJLAZ8X4h9ySOdNnuJk1Ohxqkr2tsq+JDStCcZHd5hq7zgZuM33blQNrrXUXlc
Tl2iJEW/wdFMMSwNWzeE+84iCzdho/6EaRTnLNpiD5EA/zYug6OEK0SUnkar7tIYEg+5hvg4qOd5
psgRJdjIxks1pYV6UkyNlajP9al4pY+270YtrlBnwfOfnYWNbteDEFh6WGYo+O4cQALxpO93K9Rg
Vv4c0+9sxJf9PUAA4IsXy6gveFS1WkZFLl1MxbJIjIdrThWZ28sRfCPJEPY3U37ktk/tW/JwIKGC
/PFYwBKqn6pnAHT7q+ewDR1DnNKvboLTF1UWA0sQOWpSjsqJ5yObhwPa/q2tEPlGvOfWvAMyAQIm
08x20H0lWivr9zNI/RsIklySUz2PzVNND1RPmuvcJPf6/UJPx61sl1sufif0u+RTua8TOVP8mvNJ
icgmGkuLNZB3jrVFNilixuddvmY4UZ9iO+AvFUpQDWApgHhN/wUcPiwOQFSGImEAlQV3Tb98Kaws
OvFlJHeQ78j9ZAKr4IPHtoHDAOTRZiuxhQ+RDUVT8meYXrLCMYwqSeAckKWu05TcHAzFB7AdFTHq
5FFGGRRoFWvmYL8VaSxMxevikzg69YO9Guu0I7VSwvfNNwxyHFEBZLHtuEWOJekHxbaPG56DJldy
P27D9vJFwDa/gtHvDWsEBAmAqepI98wi7X0pai3jUJNHZKUYPWK6a8LaO5yBkwJpuOVsckL08WoD
IUVPCKMxQBemdCMeQ4PVslbm5cZn3DsCXrRx0+jiW2I6NXPLQFBAMsgM51kRkz1AmjumZGh3bx7F
EEDwJLq51M4PyejFJ4ddX5lXW/uDC9GmR34FV6XVmEQ5zSjxOS5hzHwDr+4tTw4MEH+7jNbLCsVt
836Pn8uKKk83Fa4nxI8QVJ4XPrbIN5e5ci0LE3+vG0w+uVVv9rGlsVRjiM1FIWALxvBT8UMOfFHQ
euEpg99KwWpjfD6DMkeiJDY2PY7WugQ1NDQ7u6guz4qS/RIkuHzmLi+rd9Ji1oWBiTll7vCTkXuE
mV3caW7Olr9T3Gsj4TqKi/qKn2caRRR7e20RkUJuxtTD/n9bot0eszT4nnYnERwXPYAH79Es1jdC
eCVlg5ewCHfLC4pAK/sRr5O3IOA6qvgygr6XC2Pi3sIaGEIL1ka2gFb6k5fvbU9HieE/tA0s/CeF
4/vaQUqFiHcP4eshTKt4y9RXu2axLf8qVpLJeGJyTDC1bGS62jgQXnvZrvoZMXHInBRIgi3vHwBJ
CjAXm0I0uj/nnSg2ez8YnbqDLJETU8ykVF6uAnnP5udk+nVlYA+YhdWFV4LJaoeyS6g73/iLU6G/
1I923dZIFVvrz634NXjJaV327o7CW8AENMzwLk7kIHsIfdR15eZyuD8gwxzVu8kqJj4bBt67w92t
L2mknXpFypsTdDE714iZWC9/1bmxHSN8HuEZfiuoliz/yta8WTS+6rmfECvLP4JDJwToF8aKEN5N
aR7nwF5UP1LtZ+f9c50c2oY/c4ldSC8Hj4T3h/pgq91RPV7mX3mmYX2Sy6s0lQJjVzl0Vmpo+cZ8
cMJIaVlaps2b45b8jO4c2v/FyUOOKglWINmk+kU8ebZ/KMD8rJqe3AN0xJG99SJey4zUA1E//beA
w5ooKwR7xKPmdFwn6T0EukorfIhhFojcRqSkp6pZC0SfRdGfTbovOHYFa69q2Evm11yEMpxzL13/
sJQVj6gts/eLl/ocr7v0I/U4blSo/E/PQ0X38W0Q3bpRzQ1+hqQpgZ4kmYE6rTsxGZLbLbqlGcFb
x8z9jSCYCpVFiXJxWmf0hAXbt0BczTm1k2u+U8MzM+Boh+8kUPMZO6jt4Y6LtsqUayIzkKWK6V56
xVuX36MBxU8mGqWYzeUzP7qoWW1nwAzqcWoKnGL91L6IyXsAZ+6uRZqGByQgNQAPggmfPoO9kNJy
q2oPnuvsL2VouBCvXfrwIrg9WdUCdReXdsU8fqSY2WXlCtpes83Oz95+Hgiqz68/C4DROYkoKy1O
yjujg1UeGzuVPCGJNqA1HtdhF1i1Bz0B9pfOk/wimbAFqt+b7gVlxU5bjfvazCOKzfwOYlzgl9UT
jZj/9yg/ObA4DrILo2oZuqwF0l29N327SOkXkl1v4udWVq7gSF02JaCG0D/orH+/lIX8WP31l8kU
Jui+2p4LBgWtsOXqOFqhRVWQ4wuVYt5HO47PbNE33EC2OmDmhytHqg44uKU22TuRa2tGoSDNhmdA
N6W0VkuzlL5xlg29LKlEjMWm7/h+Vmeh93rDjaFyHI3vKCcYDiB/9omdE+22fL4/wDbaKIi1FpML
sTRvBiThI732nxxJfSqn2ByPwzflnILJYQvZeHnyA84flpc0ds4W7beDTC7gWLuTrhOoQemorRiq
cRpAPmL3y22h3hCEwVd58xOrUrchfaeaomXNhnG7rbrxKdYRwI1acOTzdcI90TxjfVfvPdi/iTQ+
mX7RcmwrNjXO1Ok5FbBnaH3YqniM/i1toEsnTe/cUNBIyUSILdI0c2zPFfOEBH/D6eI3rlaxRCki
Z3pHtA306OHc1O1LLphLa2grYhwvivh5yBhQkgBvSfovVJMtnWanUgu8ZtSnvNybkwEVro3jTOYz
2M6oPetAxViMTm3u1vGPSDNMh7aSD4UnDnHOSLimEEgxOwDASN+SQxNj0oh2YiMjilcncVv65diC
FxKiLOTD7F89HyE+ZctUEqJ4jDA37cha1mGjr9bkbtAnXysDLIoS4L0HwdzqhBh4vdaa/Xd6rQ69
pJtW1UR2vvq3KKOEEXm5XrG7HfalM0BUYsICnwKiWJtKQclGGhu5HHtPsDWZF3LVIwx8kPsgwNZf
mbVDCnUgOqES5IThybQ4M1y4k5Kaikl3v1zzI2HaCtYweQuxyafDoLDRnryDZ/xyc3u7+nvTtYRh
7AaReIksdNUsf0iJSNxD99za7UAeeIoMldmKuXn4ON0tA/RAV6oPcwN+RUpjVgasZrFn4adB6uIN
5QXnyK1asLLRxUo9QpPWxV8qM0MkHrIdWegFbQDo4dqERwcgRLEHh2Zndq91Cju1NW9qappxUV2e
VzExMBSqYmFPM20SkaWEQsX9MwWijcg5ZTrv+Z9j6RRN429DS6scw9DWMzHzgLQxXeFAvxoGPwOZ
djqDBEr+1zUXAn6ezpctaXlwifmhNpFj3j99ProePq4S2pzEE5pbUOj6qngVbw+lhFn9Tugt71MX
AHgkuQkgPmhedjgW3oJ62DGQh4USeSr4HQvxtNy0pQbTjKYrBiJGq7YCW3Ooahm7q/rpVKO1aHJR
wHX5oHmw1N1NroDJEQ17webA3KI1d8KTaThmZ3iuxl5JJwgbKBJBVyS6s4rDZqZwJAH6OwiY+4V9
IysW3KY8rogMZo5JQpj0t0D795rpO5PcjmCP7pyLZkZe0VNH37edGfwdAqsChjX5Zcu2UFJf5AU+
Y/QLouG2SkPjHLHrktewwmxnmlyBYyWXZuUySRlab+UbK51QyZhHDHxLtFw94LCVqDq4jQ+lv9nK
Tt86hYe7562jbveekbXPciIPvsHnTR8fb20mQRYISiq5M1plpRvvWaVONKuQNcuQ+CMsJQXkbLGJ
CM2DTY/xFVWlBq2vQUTe630H6si7WZvEPQIt/0tBTGzJlBXdHKNpdh9MlOI38/9LqPn0g2A+QHFh
OeV8SakQ3QUyfxAple+uLGKu3FlosklZe3rHwaAwnx4s9Szp0DJCg+h4griErM9Q2OdgBu6WzV8W
bVXjg7ITKcy2S9C4f03VzFISFTPgX7gAoSctLnjxSlcEPOarNOugKRdMf3gJUusPOhyUq/gTOGr6
uUnBzqGeICccsuoJAE/G2AXtJk3WZTgCEYOUgwHcq0R41j+9IPGzgE8BWFO6O5x/nHyOlwEcxsxS
Yg1Yk9l3cayPdYoPwwgF7loH9m+TypmhI7CPevnOwelZ5f/YU2+cH/baK7CWuDuBVNHpLcnyaHmo
C3GSGiHGsV8kiCquSOhUF4YsnE02coUpqnfm9f1/tB5qEOh1DMSYYAD3BKQcjsfadt+K1VgG+lvb
iDjZ9PIDZWpC4cwKR+1ZugGvOGpPy6Xw1vM5HQggL3EwqEc4H9FV+0i/Ykg17nVSMkcI5wEBEEv6
RYlLuaZcnEdBtFRtQI0vnBl/lJdBHC7jtyaFrFQqtG14U4d61eqzRkKa8WNniBPx/YtwHmBO522i
9LcAJ41ErZMx4eRKdLkO0I0gsmgzFsZh/CtL9yP6HARMWD8WI7kkTd7NCRFw6UZWdJvxQSK5pNfT
DH2y8fSJ8+D4L5waTnnejkNLU9Ri76UPip2wcIsnCs10wzUJYahHryXGLRo07a/kPdBiIw2vmT4l
jrbWvGLulQzlylErkje/tpzffRyjcIMEvPUXp8ImJ4ktK4Iby6cZVC0S9praxmFlaEpaHLUhn9pY
9jQ43KRKGHMrVZl3FaSzMGUb5zzNBKDPidhn+8WQ391MuAV8+Pyvf8+D63fdK76goxDLKgK1QB1X
2JPI5cVIlCs1YysN9lOxiI/2RNbtVlXWFfqnO01V7Tn1VFBTMA7VT7Hn8IgEFHQBDI1hOQ1uFUIa
EJMss/Bz708n4I19C8ocsugLOPj8jYqi+1TCbNZkjvyeJsFb/Qknd6qMT4lfA9sTjyyyFxoWSdFm
jj8hzDv1Ak5yZHUMbZUc7yUyP6CUA4zmu6H4KekYwshMViLrrffBY55WY8hVeICGQvnozhUtg43t
scOJA3R9hx0usdW02PpAAV448h7/bnj2+u62dAjeiyaZ5LcUka+bthxM4uI5bg8+giqiRiATgrxu
PqvH6uIo5OrvMfZFDxU7r46KSa8akLaBdjGTv7Pp0L0VCNaiqKsXNgeBVDMEgI865VCjVhXW0uAg
Ps/bSKtj7oRImVjB1GlGamlw8V0MuxVXtEpzYpSchKRG3g1ChAH62gbox2UYL1vboj0a/pmc6U7S
SXPn8PhnPiGqy99KYjfrIXUh6aj/ndofSkw34V4BtHAS7l3F41pm4C8WvjAMdH81bSyOdEe/HOmY
Q2L5Vi++y5XjThTxvayuGqnua+hME3aqUxQxGh5ZKWx+yofkpI5PWYoPCaqELyP5WhpCpaZCHqMI
5grJ4DUYUe3onuXiZtZ07RIvqqafQZSrgZcsbE7Pns+PrAa38VVT5XnKbX7SrV6VozrN0mNpxHLO
DhPujTCK0zB14CQLWmVkCITBsB9ED4trFM5amcDcCSkfeWe5pyrocNTF97gicNsPat5YLnPkOM3r
YxwSCmEPpIhIqgdFNS0jZ1SWrSh3trxq0Ofex0DwS8Hs668sbyBPqTv3sEVhJw5nzoUS3DZpKypb
AhiuYdCWdsNQ32M9HG9T50WWUZ5csr6RocIxjJnGMo8Czof9Tg9TtStXZBAAa1/nf/CptP+F1oKP
FmOyfgoNFD2zMVKz+NJsahjuyNsHqUVbrLf2qwv/Nu+n415E/CBdMfRoTEjSXqo9ruYiEgz3rFiI
pdwZGG14iE5fyJ4R9pfwiMPKGCOqKk8PTPQplNq8b8U6xv1nwzsVU4cT2hLaAZ5GKf/BfLLkTVmA
hGrHoXa3Fci/Tl1b9ZhdTJmcs4YxGhaXtCMWmBO6oCDv5ZXWhrJRpnbsu114AGPfdca4Q0PpfoI2
fo7abVg/Weydeyka5gj2L/6q9JTGDRiCFrad8/Zhv2p8sjGPse9Z5/RFXLUGd6bA37mNgU3DuNu6
ih3D0jkHqQFoEjzHZyvCpo2UC3bcGvcwBAr5tiN5xWXeLi0taV01shJ7jvEeDc1tXgUwI1p7gv90
PVLZMV3LY7ScS/IofHAyS6YYAf9amY5wxVImqYYjCfckVI4sPdX0TdP5UDqOC1t8P4tQ/q4lhgv4
Q+Fi8oK3XynJgtW7x8gnXRwvTxDdmfXyrjg17R9CD9KEG2WjNQyWcEJEX4yoYjYtrT26IAfVUCqt
f/MmfJjhWVIZWonLRlc8qAn0OFs0lin1qY+is4BeFj6kjPrzxInqjtTxclzO2ze1hUDwta3mnJF5
VhcLTTuX75mz0WeiBWFhMUxsCoz//ikwgDBFomIndXCBdvPBIDoiAeAuvsaNdGz4qI9GfGP9LHzX
CuWiUfOVOHR2iXexi8PnipeZGucuY/iWjoIw6MyAYjA9XdhfRyLQi4gdO2Gu5IHAi1iASgtWWvMA
cpmvti6p4io3nFnQTU5GvHbkGixkVlGWxFBmRFYqd/kft52aofq/t02i1HAR1RIJycGmtz/kzWsN
4OKVZ2S+mArKh0Uy+ttl0xj8OmLOe2TpguPERIfuxb3FQFMCgeg4TROoYwWFJciGuTqD0tSKm4+o
L0sriepsBpHMnb+NsCa3yOtAgz/QREDb+IukbJ72JwwF8d2VKis54Bmry7nMOoXp7Lg8uvhN1LnK
3oC38lG8lkyNjeFCAU9BTnIRVrYLLaZGJNWuWpuIU45wrBRERhzuMj2PCsXNcIzgPm+UeQlxLcd0
Hb25iEeS9qx8Gy1Wqwue9JCxkx2GhzonnnXJCmhfrEMpPGoVzEYwj4HY8fHcY6I8cDPDBlALv9si
sOp2iVbzZM3+hQxhg0+GzDtRi18HxWpWe6fUWszbD0yL6sCOzjVFRB+GucFDJEYJS8DlcE9w2Xse
h4Smk/Cr0kpJRNk7RmBKMK2UkZjdooU9AYOG6x7apbsMfIUWqrC9x9of9SNohF+eU4p/oSppciYu
xjlIBIfoYxCQUu9VtGdH5FZ2Yc8lzffmF0Bxg49rPt88bx6etbaC/YBvtWYTFoE3yXbXTVX+eY3b
vDlvB0QEcOJqj62Cfb8GDsp6Qx53f8fA/htaDimnKnVdTXDAKs/56Cnse3Xez4vt7jOwQWjxqCx9
AHiaMepjgfdITEfH0EPaXi2R/Mfriv/pyz8sI21/8tj0P+7gD5A0dVFJcNfVdzjY+2V1Fx0oaaRo
73Dx4J3h1uJuHR/ifAxmysAdXYJ5opnPcRNDOVDmOfVFKFnkapOGDLSoSa2ZTuSYXqQlOHxN/B5p
QrInyzpx47voDkGEnv4oW4HfpKiRJlWH7Q/KDhaErm1RCgtyPPWdQ7w1ieV6WqkcdaW/syQMwCjP
EIUaECjy2XQnGgL95HYlEDKWBmZtxvcRm6wVWBXbMFya1ptMcYQfl463btLFzxMP3tlbGDK7/VTx
MUgSo+6oWZKfoHS9OfAgt3INkeeKjpMHNYOHjy1eyMQmZgst+stihnM1vW/vpr+efvAeU6xqFrRD
Ix2OJ37OUeNCDXrlQjIS1Gpg+WEeyfVghDkQgrqBJkS/3lvIIl+8TX971EM0i8F4nyPVoiKLd1FQ
yvqvEtqUzJqeOUALwP9qo4FvbRrCrjeQoLRXRQsGz6bmXHhyffz1EdRAL4z8b5OtE2aeX/BLDnEH
Cs+g2GrrGlu3pqlgR4LXMXNdExftGLXtOnpXINYRiCy8Sb+JagENYVj/3H08nzrD6HPrWhopDwwV
U54udXnK/k0AEveyL8EUNOoVbmIew/XeIfRQGNDBM/fodu1EEPc757zRYHESMtQUsh76z9dSwFZA
WbGbEg5sZb9hHtp/AwL0/jH2wdqbfPdC/oSyCL+DClmeoerrlaHdhTldTdF9x0sPQYjLkBoIiRqI
Mf/8mpraNe4Y016HUhrayu6XwRuF8GLUSScSNTOvlLR6W1uPOJBcloxcPNgWl0xi2+o0RxBSRK8Y
2a1dL3UW4e9rGOdB3Gn00tICbe5OJHIAtX9gTgWs6Vqg55XSfG4Xo8h6wfTgLfXN1gaSl6r63rOV
/7AZzSqZ46XTu5qBeeDEiW8ZYYgy4EPPPSEjB2pLycieTOnVad26suswmqecHnEMhdE+gjJLEiyy
eU4CY/Hd7Q+C5C+GKKJcFRAaAejDXhe1I0NapuWrx75pa+PM1BYiwpxSKps+oJIuV9sOz4DI+IZ4
IQvxk3bgUJlohfRiOEFUnRn5f/FfkHw7qVPIVLrejT1NazFbsG3hhJaaKoTPqR/n6OnyX+KwRSeh
PCUQLrH7e0uGvZcWS1KC3JJZXXgUBm0LHKXlNeFJXBnorbLIJ96IGsRB8fjPGnmkAgqWUCNbwdEz
CWQsJvdeLBBp5750Ber+mYEWpOSGidLjC7zHvG45wtgCU2mXNClbyFiqAisv3l3sHbxjm4p8ksTo
2nomX81Oqiknw7EiKZjqnrfFjH1kBnH3zsEKbARUIMwYTuUM05I2m2c3wkNf+jn1J+IRD8AsGNZQ
K9ysJEUmVTnez3P/PIT9m30UxQZLSObC3cYz3TDMBsYh6YYt4oOE/3NJd6+s2wP+BRJY2junwxeG
nTDGULy5trvbpvz7JbRarqKzRxmEoB9PMw4zMmFI5BW+8sTFY8KlUsQUlRJMvN4BoLbn92Hwbko2
uEa1SxMARxs37WBFo1/lSnly8hX+wv4Wt4G3QNGfcRfkrns0qWD44z6gfzQAAXWYUBMpYgV3lQ6J
+IrVHg4DANzqdF6EAw4VhFrTR72j/RYPJMAIOHs39m9vALITChruacflxSqM5QnbljY9RkabAeb2
j6izOCbfsqw04Se7fmPWtxQzYayBYnqLykJnqIibjsh4vfqCR7RZ77TD0iK6N7iw6aqMxvJ1758o
J9shVmW3lAtbCJ6SQiEeZ764hhFpztgscdw8ajEosizEk7KoLH+mWEdTw7ojeH2bJRiql3bFB+v3
7YuZSkYVjVuiIaOglwejYCkujFkIN5MiAYYl9Z1wDmrUIOL/AkY/j9t/YX+aS/RMcdSRvMPScB9Z
/MIJrz/faBzsoorIvla8v383v8Dt1yKPmZi2o5sZvNWP4wdELsQ+5ZQQhCHec9oEJyc3GO1A/Xv4
ky2C7f+S3HXBwBENQyv8byoPv1bQI1CfxLMBEHxD5OVv6jy7gB8uBn7Y3Wh4VM4sxqGbox+91W1G
m7l6Bzfj5/r81vp2oynrHZzi31QEU34swLR/422QsmUhq9nWGatYc4oU3EIhoVuM5USeHsDiK5q1
Jyb0MPKwHJ0nr8M466Jucd1z95ASEY93e0UWbfGc9Eh/I0KXVakj9V0NK37tRk8JC3PFpmfykc/H
dDyNEudYd2ytPqh+WcR6IBYomfWUk6AhjMcvTz1AmMu1743gtpsPG33JrjL7ghgH6GlFEBn3gvQC
SDoJWoolcQFy9VpXsklkxPAy17rYImCWBFEiLNjrYIrfl/2aZNvELZwu75f5iF6JP+8eDGfDvWjS
+qj7nM1IZnyVLvIAdhx7hckWQw/qdoK+LwckGZCPepNjuFsOcmWZgTUzQU8qluuOEl9DxGvWyAc/
DrGIgcQtRlKpNsQqomkaZqpY7nFGBhL23vgydSta81z0zATCAcxpIEDSOeLyLt8FYsjRFdW8aAaB
AwIVtBn75P1CWcrMk5+KFqHK8dj+PRUEJ2BzKBDslU1HFsGu3x/K8kQw3DTUzhFvNIJ9/huKPKAk
JXx9dkvGCVxhrUu4XzkQXgfYkMgcv6lNERWhXuN1QprsT41pizSz3sVRTZvh5TZlUFPUcoU2otq+
YVsbwr1xGWXf6GMXvtSt8gEDjSIrQgPouSidhOkK33OXLCGVGJ7VPqMT26N8V1dXQ22dXjLkbOzL
5DNMVeKzPgTw8sXvRyZhG3bqfrFoHzNA94KMyPWGfwKUTasVCXxRGJCM3ZKjHhmwz+zLLJLbbhhA
lCymGLjYI7iFWAQMuYrqN5v9cxnuRxMVGyp7rLkqHBZ4PQMrqyKkoCKgjd5E8/c9p/5/CmtOK99Y
Rfyl+X1GxRDEtEK3PLz9D/XQAiEEW+L4LJp+Y/vbLQgedk713ruYhKv5F8/JEnGUohPphlWzcpf3
w4C0tE5dYAYbkoOQN7pjmzYFA7B++qCv80ZQd6y/xz2grmXKQhbPjOICVM+Pogz2Q5t6XZN1J8UB
C8faALXCVnVuJlwfwwwxkTexkxK8QSj3g+2iYTFFevywMDpGiqvzzjD5Va6e3iFREmfjsHxb1qRN
k+sCRJdCVCoyARNFBoSVI4wgkmTGZLZW989nX3itpPCgiMNseuZ5OEJsU64Y4hp8dPwG+faIwP87
Ib4dTVHSuSHY8INS09n7ag8JF/hpEzOpa0UBIvJviOtmkgetkqr8Rq+8ikxdbSCLYVNpFkxYyvLk
lD4SRCIy2iaKHMdUS1W+fIUYj84kdJRuNa7QZdKFfa5m2DRWNpYl5/wfclt8U9yta0UyXhO76dje
cr2URB6M50G3nzdz7tx+7+BpfQ032JujBJOkm1Es3AnM65qNcNggGPqErnQRTUJCCe/wXcHZktJy
k2a6bnLP7fgAZRqaWmCzAyjbMJJ5vCOLKBjT8BtOzRQ3/oIrR9hcpA65KTCK3ZsX2LWWi4issewv
2oJ0xnzHIo1GE0ogXrWIAFM3mKIuNJGczCzuIuV/LSfbyO+FKoFRJUP909yExV8JFLybx739xyWg
TZ9j93v/T7GaFhPjFRD+pqITVjZbWFmZ0s3PlzSzB2Yy+n3VGC/cHDQ0Uw4Lroro8d37FiujD1/x
kKtoqbJUNnnvJ9x+hmKzIW4SjoPaDP7Yv7E+sfy9/Zhtf/mGFO0DseV+0bQKIibHXpGiVFb5q+ec
0KYbQUEodGJvWSz/dx4WOTtPjrDC3NWK/QumKBxmQSLQ9Ic37+Iw0pwyb0vpV8bIO4HVdevB++qb
PCKVftAhB7GtRQEuHX4yDIWBA0dxs1iHDo7QoxVgipQcIkjC3ZGwSxbsLkhI6ppe9QbbHeABegQd
kdzftjV6RDeQYFNogqnbusMHFnb8LJMCJrRam1czcsHAg/c2YUjCRx+0VhYJYvxF0a3jWgTDNP5J
gRjoxoWkzE5ZSXhWK0lUcnWCwYyPihT0z+VMHOI74qC+A8YOTl3G8vZglj6eqMx0qc+3wP6LAVtx
lDK1Pr1woGq5ydPLSwTNSU758pCPL9LZFJJ/RvstXzHCtVC6K33GPUV9NZ0vzNXHUXUxq2BHsJp5
4bfFwOcbhoupVPzz1Uv31pduECbTq4o/wNQRa/O53MP9NYdB5ABqJXm2wYhcWamQOjJ3kfexgpgB
kWHbC7F07Q39hN9muT5ra3aPAZgcqzpIn4WJUgRL/Oj97xDKnNzwis0vCaGwwG3goX54QAmbgrsi
4V6MmIB/ahATqtIx5G/fz0hTJwpDpNMUAeBWLCamJonBmmSUT1Merf9E3QI89hnpTnmAv7iy3h8s
zb43k1Bz2sL9z8yQLBW2jZd3wBYVqD8I8J6kdo2MGlAjeesoZ0qp2WzRD/ImoeEi1A0SUWs+UzBv
pJyH1Z/YX4i0IBgn4csmlvHCouL/k/8vgJhAboL2awmW3YvWNxOAxOeGF1v27nCxUQL7u0ihlIJv
ppYJSUoVer7lENkA51FfkbD0/kMXtwiE0UMS+JLo7XcEoWCkliwv24ILhYdxSDz1jWlWn6P9qsn5
BWLFv3TaB4yPs3nh6WF8EWgZtZLDmN2cXnTEmcYLaQmpdRW9Gi9ZuD/c8n/qYPrTf5pgzcq/EbYB
9lIWB/kwp7299aD0xOFH1NYEATN+axkdEUO/sFoTkXVZ0bSmKbihs79p92hafGrtKJzNXx76K/iv
m0a9kmvyxGCJl9REAQPnfndrWh6/Dy/iB8ADhhv4txG+/1w9RnS6yuibeRkt7VbNckIpar7Vh5DB
KHowA0s3J5d9UQQAgckFu6WQ/tGHqe5dHSjNCHPnMb7Uv7wtN3mfQ42HaQAMbS0A6dr8BvnimEGu
aa9Li1grPgAQHR9ZXkJPeARNaVa5Gkw9+4+IlMhXuR1OIXkdfU++iNey/EP0K7+N5nx0u+HDFQ+v
iDQb9AosNYL6yuHFfZyJ1QB0TeJqHwNiPgwQpFOOBpx2Av8CGk3I52fUhJxMAwVxOTEU2n2NwTqT
GRFNbrh+vCVaUtpPSPSVs57yGqroDkT2KCIJ3DUpoGA8R63NyQbYtmNS9Qsz+DLpapsjb1xhzxIZ
eTSOaqkGFCMD0G8ndw9xrJyj6MIXXKdtXIJh3vaeXoe5dzHWGMSgN3m8MD/LApOdCtFxcQ5p7ASU
UOHb+3epbXG2jc6u71Y1C7n90Snd13Ofq9G2PSSlldQKYQuWphv9xBbmjmcWMKnG1I8dPBFQTtQs
AR6KxluLchb0le2htZKblpkWleZLgI3+Z9o6+YMSQDK0nCapv2tI71pOw8TfZWL0hY5Jx90NlVXu
EDQF/RnmOzwCqn67AGQUkQgS++jCxciFgCMWSXnyg7R58eN3K5XP4hBBJJ1vrd2J7I4Fod1ejOZE
W1HeN+2TjbTcS4vOYGq8SUgfzok78U/G6IUv/XOi0jWz6V1J27VgUXS1qNuwGBbAFa5CUOVX9oit
vxj88QHVPc5SmYpidgFHPT2BtvgwQGpIqsUZ5EWCki7jx/Mbb7/pf+kBO+KScX0PwyTUblpvfnGI
8wlXVhj593hFTHfbsMXnWRczBWYUq427/275e6UuQJcCEZQ6jLOi0/IjjHmTVWFx5eGiEtw+2BIT
y7mgqI5daBhqf1VS30ak5PatI3riGUq6rQb5buiZ0+eVFHMyRotG+9/RO/mBQLiz3JXty8zARo+e
GfBbb+KBWv97Oy6Y/bTy/PKhqVkxkKfY3vmwCWHyN8HaQoP9Kq4JViGR6JWyN907skdG0sDd8j1s
EWEaBfYnhRbRbF/sMjcGwP2AN1LMwABn58eqZLd0DTO/111VsvHiMvGN++cJxHMfzZfn4aYFQcjX
qSj8PZuCwWa4GLGGQ61B2E1/X4XLWa4phvsD+7i/EICpqz5rlXc6XWE0fYGEPeijK8c0plnM/C3g
9nnuwU9EacUVP4yCL46WKmws6V6sSC2ZFKzsdzY512u+H9PVLvDFJqr248x4AnM3mF/9Wxsfquj5
rAz+M7wav0Ap/Bg+Xj3Sj+z0//DrWsLnl1cUVTtB24vLU9KHEUqWM5cLVHHQ8V9p/48G4MFbtAPf
nP8DrucZh/zms1l+alwiKcS7fQOLc1gH43JEcgAolmO0yJTVRi+taKhRI32e7Lv+Q6qGWSz14AxG
/WGxl5rUKblq7+fYhPMKsiqCEJy+gbd00TCKrU/w7IQVvvk0z2ha8LSWaofSB9pCRMzaeEdXd62F
6tLBCkaTrU2CXvhqB5s+MEJoJ7Rb3JH5goJm7CcnD4b6WBFjh7gbSbEGfMVHDXDvK+wZfC3H2ZQR
S5Xu69iLSYOU5f/RuaqxEJcapNXAq9CV63ftfoq5HaBIfCkDAGEHs/hRtpnTer9NUiX6z8/kj6gm
WaKhUzc8QeawIqSmwSN2XgX/FHQrMcP3D4bOTKgsliE1Y8wGhq7UAFXkvRgsV00kZ8yxMCKZVF42
AMz1jITL2xvJDBGUglnKL0erISRKUnFRpZiYEzSNpZoUkUN+f15x3H2sn6Sj1MDAKevHnW9ZcR8/
Ph1bi+Et4PWXag8S4cY1Uxwjc27Ot7RZb8qCPsuC2Il3CLF1KrW8Wadyxm7dSl3gy1sio2TU55UD
YP1LzkG6mxbxfljGC6jcV5NFFdGsn0KYBiO8Y19yZ9Lu+k6BTdmV7n9UZ+utZh0calWC2yt0TdqJ
estIIT/MvN1j/eJMSisOuANWoOVpQAtnjomFnSf2W2/zxf354CcU53181PVFeuOUfd41lwAIURod
Ut0DaplR7tVdt1PeIhwUkG5jxqHq481Qq1px3HFHddqyenzz+Kn2XAKyZ18yE0JQLko2QkgBLyDq
QeHDRok1ndywvx7vjhh8AlLdi+sYpeAOeOXm/vowHe3S7q2EsFc49ddhtd7MhJCFZougfQsmNEbT
PMdsWALirDyIGvkCGCOpHV2X+dnja0KgX1rOk6qFNNCkwSyIk5Eza08A6HKY06j/FJC/sRSNs9El
e5i6MacptDNDeeBA2u524LpIN+OTxJcLze+wWGeER7hYgDCT7dVs8UyupcQm7EfjlUjmf46KCNZO
teTqnZyNjNqzurM2IaSFWKZ3GUSzcU1qF+OH9VGMXIpEWit6mRjYnPC0VjujSd4dPiOqWGbF68Ko
ggaBW1i7fjB2fDKFX/NuGDEe2jn8QzwToqUH30pl5KCmxEp1fIVPqqoWF3hRzpNwUZRFx1+pHe5+
DzOnxB4GeWtxsZvcOhvN7lbjTWfh6uqzb9dDCj6DD67ISyMB7Wtn09Lf8cv71zBJwrO6WYjFkQCs
u623V+6gSndfcOv8jQ/w+20VudGasFMrf1/wB/KCnaStYJAyWr5RUWhMXTwvsjkpSXp6VtiGGdF+
neBdio1s1mnJG6kEztwU+5YutGS4RSOXvncKSr392yPSq83Wa060eCyQXCOhU/xJA4ftTDyhmc9P
JFc1aq6AY7KiyUL43BiUAyJXTiHVm/Y4wZPzo1G04//vNBwdEyR0iqiXG4Y5M+pB9uMjHL7gZ2mR
bw7GyZiYxZQTa8MfStd03rR/ZUw2Sz37d/npPz9nqgWRMuqYjIbEQp6p98wEQ6c+rXUcMVb64sX9
Zp2j2aw+UxIZCm7VIKpsCmm/wngESVM7+PkK0SorVgr5RYFm1DZfhQW9hekRcSTKfgcSnxwzGgfd
b0+vkG1sXA/elWhdRHLpyItmxDlkyVuWixB6p/wKN43Jur/lM+4jNqeNtbnwgsHWm/BgxegNDtZV
wKaRPwsd9sCEk2jC8FcqtMVHG0GD/zxfrDS9xcaHQd4BEtoAerDF/Zm0fZbukltsh6tCmLtR+OBv
LTVdKoc8LIXrSW27FrfEW6C6P8dnhVid4rzK0eXShVqGbTlyYX70SdUwS6o5KOUxiULLrQ+kWmgI
BRYUTBP0Yfe0mhsxXcf84FPPT9lbp55vaAK0VG9Lm2dsQ5EYs1Zh6HKL7W9KwpnXDa8lps65wnD7
JHE/RlcX8mSgh/pw9ZAhQj1J0pNanaAOExdhn5Q5ornND+Seyk6yvJCWe8Qq8VnoAWdaFWLu/2LW
B5xXVDjnWHUXlvdosZrx/gsUVpWo24E2saQryCoJ5ltkQDO8j7gTjnzyOD6sUB78hooW0oLqeoog
Nh3jHRn2z5fonHpJju1qOZ2MfYK+SRHr5D0/jVgZGKKITcL/2MNXxL0L0/Wv3QUu5Tl7Fvjvf5Vh
NIwHgshuRH7uiKZu1Tois9lL7ABuZlQAaeRyRmo52XG/mI/gUPMTHAzUGapIfBr5AyWDCQhQS183
rxd2FXau/4I0TZiVA8goUFNucyTS5RjDR10VgEZHvpBbetsVCKzacQfiLsGCc10Zrg7gllMqgG79
G8iZeS1YOIo9Abq9h2U2KKyXijLTPyKzdNdspQHKa9y3SHdIUqfA+afIJK0vEoMOF60Vw8bw4E/M
H9NCEqTbttGPPk863tsAsocTK3h8YQTE7W/HiKI6l82WJJV17bhIcRHWbEKv07YBnUu2aKrmxSPQ
11eaRvnPWbkzrW3fr6piuSoR7hFs80xvR2jyf+rQj8Q82v98okBrIykW9JfhgVETECI/4o2iL4RB
dkdsJoMYq4KGI+vjcc8e8zbAAQHtGH2ayUmyW/ZpoXnGqMutGg56uZUiHEIqSjY/f/SWbh3gAt2h
LbNaRRnFWurGX7BGiC5sWpeIelZYWhpkN6L0uLZr87KHjd3zu9x/YRFGhGR6RzRv32VLO0fKVxdD
BOQxygEbjGDj4GLJzA79+jEqyiWUIPHlJYHMk2wTxMRAgwy5v1RriAcF2rReYrA6oVWDQO5t4NXW
e8UFaPeMXgV3kCGh2ry3KDYTCLMdUh6gW4gwTF704zPmatRH0o6H+hNxv0N2vQMyQy+wCBBeNl9a
OjFHmnae7roe9siLGxbVsIAvOiXKlwDTWEEg39gzV96RcCKO0gFwfelA6lnwu69guWPHitSFBUjz
GVXtg8ia2IKG3TPBzP/GpcnLrs5UiKgMTFBuAWjmq9gXixIqT//9HOXnfCACFxl/msPSAJJAqVJA
qWWxIlKD5ZRwDup3uOuJQdc/9+iFA6a2vytfHN0modAWtN/JscJaVftFiHWArZntHwIGftSHtQ/r
mam6Sa/604htEUtMsfDBqPTJgn6wu9rK3ZiRgZcSYQyD6pxIwLeb9veVioEzh1kRfAEWEkmXqJqJ
5Rn15jVMHjEkiEP6JG7KN08GreKIp92UJDo++586rYfF8rd+sCC4CwjutgTH4mVdfgC9iFlrc4/0
jmQeJmXemhr1+S3yhP9Yw8fsWTXk0VM/GIRmnkRxGiGRyETK3i0oqOJoAZeFK6YA03+DN5HgxATv
VC2xMbDyFWEtRLo0PdiXQ8Gb1J8rOGi4Qv7Y9wLqT+4cBAj3mOYEMmbXWDdRZqltjdnj2vKUHCwx
NYlxDhlxLWzTEDuXO5b4yf8Nmiac85S/JsXjY6nUJOOLHdktW6mmGRDlaZhWSr/sIuGiX2hIoc2o
Vo7ZX8ucUD/e+Di58xiDGY+c1VqhgI2s74oB6qJLywBbk4RmxEulL+xssp2jQomUY8iYea56l1SS
q/wobKJsgpDzNa3ncyFx0bxIHzWUcSEmJnAVl74YFk86hMnlJDt4pkO+KYIjnfQK6UhzVPzyN/N3
Ez/62k6pyHYDxnk8Na/MOivUfAfIdl3zTq3vL/aq7uVpJ/9p4BJCaMI2DL4hs7RexfxY0unrfnVS
Jya2nK0VzDqQ9TLhGhGfkiz1SiCnnIoM3yiFz2GA8FA3RN8UJWQwUZQRJC8OPrQ6waXUN2KuiseK
RXTgEM4NMyx1R5AWHZ2C2VVJNfsH76ibqLl0IlBqZHj0JZejUbConzcn1C5WA3ZW4KY/ePhX35Mu
tAA0myYyB3w6Crbyz0M6hn9TSr+O2pxNgwe9AiHCltqzxvcR5KHo2kf2nuyxhOgJNJy7j5/oYgut
KKe2PAsF/UvvHVGPFq31sCITrauSRqktKBuDg1X/0/lphaOwZGCzlABYLFMvuwkjhtup6O7fqoSK
WP4Hh84k4trTYvpGfuiQWDjXimpkZ8WRtk5rI4adBwXu0uzQpaZge7HU7fj5ZIvoj6sHLNDyrlF2
2y/9X8R82+uwpTRHYX1NpKoVzZKj+uZ8L3dW/D3xNCy/8mmlRzby3i+oS+4ADB4hRrzC2UDZV2Vv
95/JkC+ES53hVerZbTllxufKzBdAG5CVTvrjz2L2Mdifr/qhxQNm8XbshRA9ZIKH2N9Hx6JlliSm
HzPrDXdOyPFT0EY0KkoeY8jFIrLBLE0sWih6CVTnkqQVx2ZZq36zeFcnMhByb+bjrfb7WhRaFWly
Ahu8Izq1UmeXJHU98bz1OqsWtACvMxE7gGig3BEs6QHFsN8gyZFZ4U/sfzsZM61aD3kZcEPFmAJy
axCiErvHWw4xT9aIhcebDP5gwqvZBHbtECI+XEUajcYdxDl3L27afNHcDagughxMmPTqzLCDmGER
3OwBKaMIrMAGeiLRFyiMZ2l9d/tqpt87c+VrMoPE1VfB3APJ8g/Bkms79hac6qU4YKYf1XHQPlls
3k/YxPUZ0Z8KOMTiLNBi6xNlazmrQ+7VWu/0dy+s2vPcCusldeZvgaOI+U7f1JSJk0QRL1kRX//Y
evb09mdyraNSGh8kK9Q9T/EEn8EZAGfpDSr7jSPkdjleznFPWNLB44383yTITxTeGRL0L5UNjidh
boCJUF99uNE8np3oSuXMG4NYWY9EM+gHzSwFdcqWkN1Mz5np69QRGRuevMwh7DO8kFpacwKI/sEV
0Y2bDSAlE+qAjaeBZ614Lz9tgVf3DhUQgCteE5blpLLiSrrXxSuMek4sfG7cjUsZ4AXpBlp2j7b9
xKTIgxrAXBsk45MG661QMoKx0tzKvz9BXb2Aazhf8eFdvpTqVc1j9xwTJTRrQ6huHSoM4XaBJ8n2
imayeIHt6MytEPpvi+p1MGFpWpG7Xo97jXQch6ZVwsdVvYycV7t+dy3Hw6H6sa1ec6wff6kc/fUj
UtP9LgFMStbATQ/+kgXEZ106JxP7+K5Axj2QeKfsmOLYmXpac0kI37sTNybCIWmOTFoR+N2CZLSy
gKwSY0M4uj3+lGwNIJHCjWr/WIAh/gqwnH0zwSbc4HgxF3AEX3H92xiJExgAyGcBgfrucxuu5sAl
igHZ/KdLFd/fZIcgB0PVbmr0BDfDsqsyju8Dbr6dWrFyZHbc9G4cAnlSUtSWX4NSuV6yVfq3Rl9K
tt32mmUbXN/Rv6savod4KxG7JycyOc+EGpubVjwvyDVx2mLgHQ/8X2jj5oiAX7EmzJpzF0vbQ3Yj
MgmFMnu1EV/DnFrVvvMwUlJGH/9obD72+rl7Kw99b0VQQKMuHAB0N3y4+V4pPd2rcwJbJqTvUhhb
/jIFerZVbsPC/dRsQHOwiWQwu5jn7cHMSmHj0rf9zJRe07u6+lepon5FDNl2JYCMFHJnq3buwTlm
OzRuhUXPpvJagEjMOx1TIGtimkYtmNU3AcBDug4eLyp4kGI2mzrVSeE84to+vWsvklUKXdVPK4Lw
E+H25Ufxs+nlmG4+UH13J/ZBk9YY5fKnSu39hvaSW4MyX4/EJCaigYfeyC8RwfxKK5wbJasrvD4r
rdyjzypIlPkHl3/sMiVkgLLk/gY4H/mOZsRNjjrjSzOsM5rxDF+IOXQnKN+AdDxFYmGMY2l78vtk
npei3oyyC3ck/EVqV6yLKQ3PvPTCbGF8AT3HfWvT2Emvlz3hyyAUl3NG4W7VzvPwlcsIVneFLWdz
eXTzTMrMDlwDP2ioycqSitgB4h7uYoHXESHs3jfCzaXWIKEwaSvJGRdef9V+fCzZFuqjP5ah7c8o
d8jmid7HiKVpkMjFMSeGjRj/TldFCZnEOtAvOQTmyLj+ukH96NsewBImbgWS8+ixlnzSIvB60sTi
U6y+u7p8CZtuKidV1f7BJYp3il6jAu64wQdxvLDdZ96o1ymyjHQFuGwI/gYGJJCPPIUgbr/o79V4
H+PCsd8E7CJm1P6wjPzy/C4jMs/CvtKnLa4JwrRRuCdOPuewJBtk+X5uEXMLyLYV8tBPHJqTpDzI
JytQqgCd//ArEG7kXkoOPAMmYhHMa/34IWNXpPHiOv5KvBTLTIPr8tqi2ttjdd+BJVSN8qWjYLqK
lB9uLXH4PgK1bqhFbkVLqbaXhiEfdmEBZzQyNnoi3Jpu82OKEbsf9hJGwLRO0eND4W91Nc5YqS83
OdpIkoWHifMaqP/ofcGW7/t62je5QWZz+ApA8yPGiFjsIWx1FdpDrOwRXVFmvbw9OcQbx/rqAb7x
NOiBknpnk3auJrb5LWh8iX6aFPGH7cr9P9hBYbmAMOqWWx9MA/ilH8koZAGuJabzeJNMtUST3jIJ
inPK88jGpLkE5j6Vs3CRgyW14xybUeqpa+X0Hga+M9DsL0VQNuGCTcrwLMk5s78b20eZqlm+LhoM
dAIA9pMlPTJalTc4PhjnwY1YUjv1VupLM5cSfCgXMSfXWlwUht6elkvyuYZplPlzvku8Oei82iBK
o6bxMeE7iyTqcQYLxgharAsgnZu1gaZMMZ/Kz2SSy9fAviPb4upZUV2akfrrWpeKAXfCNAdm7r33
bjH4Dg8zqhRyUxWuoUYjOk2Q5IrVKnxE3QGx5VTa2m48rGKnaLwCC8drc+PVwHB6iOiHtRc7Il3x
RjDRVVDHWCtS3NIkxVnAG1hraYQdImJ1i5L05oAOhviOpCgG/Vk0092juFQk1nWo95tBL5QX29xr
mBuiLeAfgjTL+qoDypQS+q3j02j9T1dPmRsWUjhmknGqhf51FqZH8QwNEzOnKcF8X/U6GRscrmGj
RTZI61PN49Jji687LCpIf6urj0ZPOover9lYjDkVRxwrL6bIo1QnPjztc/ma2XO6UVt84q0IUJgU
Yx3FJytpsE3IhtxkW9jJMhXcMAycMzwOjbSyh7NvlgKDjJyjvRBk2A4MKab1udND9XNK8ltTpRSR
8mvRmlKckD3mOeE7T0r7adPMXre8pyNKzUVsCYQJ48tj2vnk/JWoJuirBMZFpjoXojUPXmCeFEG6
S8ssBiXw3AZFk+STA5qareHzfgwQQBIafaRsSvnQJZqdRJnK/cTaN4eVEqlDVp1x50VieQxGNEAp
SApJ980jDkQziba1lBl2P51F8e8eUsmD1SBrzlyPT53vb56CdYbbLxQifBOJquujjVH5KDFz3tPo
36bG548J9qz8c57cKwlwU7+EoRZja91EQ0wPX83X2TVA4RTtVqxdfca/kpanIsDl8QZLdBWoYYv0
Ah4MCH2HiveZEFHKg+QzY0vWzGzNxxXNWkEHo9GBgWPmQeuajGAp/UARAh/dingSVbD6lSVaDbgb
rg1XUyMpYz+adRcRuE35XQX0CXSZKhlDWt/7cY48XJj2OAETH6XitwWCJOAq9Rahh6214n7KxdL+
loIN6OWoORekGDfJ7ThBfvFE0+PRwdvuUawJfRIVE/GxN+u5EM3uVz6ui0TM9s3C17vRGun6K0oU
WjFiH5GSJcrzMXnDyptfAkOhKFqLjaLfi0eGPwVnkfIZ7WXlLdLXKdKT6jIDn3n6rgmLyvk9jjDb
1Di6jib5PsfYw7Lm8FlV2C4/KAPGPKPWnLc0gE/QA5CBbCHxx1BYVwH7XanjjB/GoSVaj5hNyknH
I90f9rxJObIpbJssFaYgvaBaOmYwKUmpXB584cvOkn/h7ZGbjrMgPiJo4c8lIAxslINJBRXafE/L
KPkvjeda+whglwoJlbXkEeFaz+Qed/pyiClJD1AF2qUp6jx/FZHYrT3mCdH1Bnyn1e5nAYKPWAQS
BeiGGBX8rhuD4bNlLsLu+rrosjjM+hl4p24i98ZH8tkzGTtohMG3geUHFY3HVp//d/EW06hQYlq1
kFiV2Mnp6Y0uRPIjxuuH4H6Pf9fXexZPMQQ3+BK5g+2tEf3JpCfGCgHt7tG6yf/Ch9GBLDKMevn8
Qomx6CNQkEZd5wrKb5C6i1hqnqopk8S+xWOv4Q7rUy3BTOavLkbWZIyqzlvVfvkY+0116CbvO0vS
MMdydndo0LUL+/sjBSa96k9C6ZPMCYwmh0Av3CEmvb15jBHt1GPzMeOtq/bZGJdMsEFT8OjkH+mX
lEMxtWRtYBmRVb75xPFXO/b2rlf2kiDft0cT5vPIGyikOOykjhliNMTNa4Be8WNX5sBOBBiPcIdw
ZSJlhfXbzNAlRByutzn/xXpvH2y1RHsKp64l4aT8cHOsztRzmZr3FqXbbGDuo54qVqhKOxpB8Gl2
ouI6bySFJUukAzGRCGkDXFtgpnRrjSMXOXRO/21Y4lj/ohEJi1mPPS++ldU00fPOMbrD2OVFv/TG
inSBJe2M+07EtlvEjPx06gMSyoCgEeWce1WyrmR9G41jehjgvvYI41faOedDXNLxU48wRVuFC6bZ
8hwOx3Tcx+6FYgd9b6FedfhIcfgEE0OHnE6tyfHZ6S+bYhmhzrT3izjzqwGEn6XuOCHJ0yFL8q9o
Q/NVaOpdGm9lUnZx4jySYP4taXkSGS7E5xgiojlpsHx7U6ztF87tJiB6LKvChQUA94CfGwdirnEy
PbmE4roWSiIXQIt8lVNpZ1kM/53wK34h4qXyQv3kIeWJGgLAoXNlYTpfBXxwFPSzImaHXtMofj1Z
DyVbcoRi8QBlwOW38Cs0zxLizUpoZksga2bIIMgZPK1BK06jqJOuBy++TJbCGS9zGpX31LOaue/g
s/FVZbt/5hzixro+6HnYTeectmX3rNOGoYjwpBY9QOqHiQ+ojLC/C1RS5fKjNjXd7QbQE3YHM2gW
z6HjkwJ7zhQcYdXvZBkBRP3SgpjoMHR/KDnTgzps33Saq/JCgXsr/oE1rNRI0ki7pzy7vH1BtPcN
npFotG5con3fj02fnIssMmD1cVMzZT5yz809sSGXSIDbmnbjQmNrkarPFTdnxDwHema98ulRpcWG
8ZjzGOzUCEya0s02G7Xai8rrUMA3fdqbgfGi2MeUB6b9hGiOZKStM3dkCxt7CPxgnCl0yHKFONRl
ay1s8J91BFKLOG3mT+zjU68T75XqUgEEX5Q09OZTAuyf/ZkfiBuG4sjnK+joaNL96YkLBiog+pel
Ijq4kldzq2zPjQE6zuIeFohbyElLlS/azb7LXq8i9I/We5urq5ud6EHOI4V03qlMwA63O/5oK3HE
/RTFJeaxADM65GQDY0pPDFH6ZhWX65gNLkkvFGNaobpVRpPdtFTZE6IKJZP6+3gGb39TLI8Eax2N
iWqgRd1LnrXj8XzLa45wqSsx1z8zKs/XE0o9T8APRH8cuu0jSB4z1qwBuFfrEzjybCB7msDxEWVE
smhDbYILJXaZoSqcJWaJHPivxpd+93d0Q0kLJUhSgodftK0D3Cp18IQFtoDZ85Lg8Zj0ZLH71dMK
qKJnS6H03mUrfU6VWq6j+hA8xz/eFez3C13/VSJYhJdnaBDFYMl0X0y7DCAtoAmMV9CaK5kDyhQ7
ALFlaqQoDllIX0ZebpJx+RXNps/hkfYJ91sSUQ13pbmUqttyr7iH2IM5U7dbvtAZhskwq6NHxxoT
i9jmmAO4aQeE0wf+xesAFToWpvAiARu6M9p4pwN5Fsh25JkrVd4DS9MJti38LrL1gHwpafupZd43
KDPrE+sMfwqBAtEVsGOANI8R3vUiItzQGKyofrGNY1QsXbuwf+HLjuXZzgXTgUHz9txca7ozQLJo
th+Njyq1Rzane5q9FtvuSASZwQDiRBadtgvRoDc9NpdNIJTbl5KFc5qAc4FVoYgv0W4gN9MzQhEz
2gEUsI36cG0ZssUwJn9RZKFIQRBc649ogVt9UGesPlPCZSJt+rmqlksGXNtgBE5IXTN+SEZAputV
ismSYvGr5wt0x1etlPrJN/FkatPhSrVYDTSmGXItVlodH+sXfKdgQshRgnCFxxeyJe7VpDywEXvJ
quwdOSRn2P9ss9u43A+NgATHP7wUM1ih0KaIk0IoL+UjwVMg4zXZvb1IbatxpxZdc41nQOS2oea+
WsqCK5TMD8rstEMnwTXR/KeTlKCBDyv8IELrpYcfUanO8A9YT6O9LIZg+gtTnUxHRwRSH/mLYOPB
/fo7Z0iHLSi1GEboOELIt1hXnMBmAWURLaWqoibDwZQetxEr/sGOq1UrvxNwtNs2KCjrl4cdqdiq
TZzDw/2jtuKVLq5X0IvqGHLiBFmu7pdGfMkfErvWe8AIIbglGFzqLSDGvBCu6Zv3SQ6lQHRpHMp2
mEIRXv56uFuyZaRUKIYIVManf54cqOdfsWlN+X//OjuhlxIHOWFHjBjREI0b/4uGLuC6GB9xYJPE
B1bMOjN5u++M4ukUVDLQdZ3zipvJc44mey3yFCjjkZ8L7JTFnZVSQr0ZZcVBHq7syG4iH0s6L61J
VdSt8YA4+QTmzR/Lbj4fPBri99pdxYiaBLHQ70AIxyfaHvdxLkIx4ZArPndmHp1GhnAtib2ocq6U
3heTrF1o4PFFBJWSKquEBmOukU21vjNh/0n9ikxvDwt+puJeVHnjrvdUELl1r0COeQkXzyDCZzJn
z25zG7RqZ7TGnjbnFJRm9T6H+IQ1oqf5yC/GKp2xkgFl+vGpvogi4rabxoBL/e2CHKP9XlnukKzL
r+8Hjh09aFgiwxy+6ph5KSqMxPKMDWretxDDrdQXhaOSvHqBz7LptrDIMCYTikeILZx1cDAK35xg
V+SKdqWB/+evvvfehloaRhyjFFwR6Ag7dtp//fyIdTQ26f4pZ49SLr8bDmbcq/Rz+OvekhmD7+w+
112GIjBHYHHjAPT7Yaz7AI3OV9BLwyvrBv4VJghcyXYW4aYNO/8NTYIjrbrArmK/Bq9/OcA9YzPf
RpEoFspktDY9SX0Yb663UK0DGtIIaK8nhVH0Utm/aiOLNUJira89YU7fM8IX9xMvuSoyk6xWoUZM
fSvJuMBMzTUF4YQbe2PkRNkGPRMwU9YzSl3+m5R+qucWD6b3E0qM4G7HnjzL/8ipC3ubdURoCDBJ
C3lxEv4fmFhSWPoO/He0MNJ3uZu7Bl6wpgdRs4bkvSOBvPSZYrs4zWwk/hovif+BDSub4CbUG/12
Gs3VyoHFN7yiHvJR5yTHMIP33iido2XA/uSyQFoUsF0XiuMNs4iKfvHmIDu+kB2ZOoc4FD0uzMJs
Sdoti+6D8uAXAoMWjRK7HcUrFjOp1GdzW6OREIzSJORA0e6AnZ20THcdXIcKC0sCJj5IbsqBMTOI
z3otfSpJ5+I3Iheab4Pq30xoBQODR/FalYTInpfYUtRzVJwdJ/yQhEGlI6dEDiNj1CDgkjh49VYf
4IEibepIMNC+H2tGFz9bNGVqTUYqvUI0RKuHbqFfilVvKOHTBZIlk14dgpaRi5dimtmtnqX66k37
qjvPVJpQxZddyJwxgprPyI2nZ1TeXlZA2uwbwEuP8+9rg4RW1P3tAgXoL30guXdN0yoZmoWGta/A
A1aiYsCtC5txc8LKyVtCzu5KT+xmhxg6NcBjZgEgeT6fLvejq7su3VoiGbrsGkFBOXqGWzH37bD+
dHrvqlZBU25sHbfxDM2dYZ3Gza9PKM6kK9e2TMjCghkjGqb8Byb7cC1eFxPYd2ev8yfC84jxt/cm
5Vw8zTPBDF3lX8xmWN8somthZ3rY3fMbT20WU2JF+sFWfFHeBVNtML1bAhz96/OkZpTLa3fCVYOH
OyYl93nzdgRGbzqQJXt8v2IgSVYgOs2fi65tEP9543MObrZuQeGr1igBr4FbKUjfjGE65/mWx9Rz
wrjGvZmeHb3/ZQp54gJLS+QL3aOdXzNHPUPAK4atXhmArvk2RB6idU3Rn7FOEXn+FPE2OS2wa8yZ
2JeU8xEHHwCxWcK+AOdYL4Mq1lR+QswlJc3LEXkE8Ng5wQ2XPw/3L4wCOZvS9OkyjmAHUeXYY+GO
3DPkPGnTrcY0kSTyozGWDuzwFGPIfVfOIW+LByENvLkOw75S2ujo4MlPYlXo2wBFJMaTK1IjHo3+
3mM0t9TzfbkKkVQa8cc1gh0jXdjLpPt/LxANzBvEsOQ84m6Hee1EBFL/E4r1brA4x+m9xhdcAiIE
kMn9hnDtdhVeCOPxWjVjVS0rs2l332zHXg7x704LY30A+Pnwx3YZNIA0YbUGO7AdzuEOkPAVCqaP
L37XuS/MeDIXNHiyVbXAks3BW8540F3JpstAW1BRMSM+sgMuBAObyqKBEZdU/1g8oJe4pI5uIqwb
6tYXwxMpZDMBdtib6sEuiAF0GBfs8PnmbZZXDGORMHsKkcm/mSdJQ3NsYK5Mlli+sTcTbuJMSggf
3eguTG58eZ3RjMdUmj6X7mysv2KFX9pADTaGS7bdPFIxMB4Xu1wSr8KSEhaobh9YVj/5HB4M3O3t
JEr6/u6ld8p0MJsbVQnbJbGIjrpAdSI40vkWtCkyhyxrSnGWJceWXvZ5AadZhK33siULCHDpAuK+
KRXP2q0gIRFf293er+5M8yQUSfhy8EfYkiwkNXSS+dXk5lczjWWAKyONeKt7slHpmI4DTt8fLc6W
iVAPFrBJFSroxfLKOLAKpiKbyVGZgle2M0EAV0MWTIAzhknzIXqe4/sDbTGrKIAjn7LvtFckPSPx
a6dYZcZUKtPkSUrxblQdrpWLUV9rWKM/t5MIaDQO5cOmOyIpf7JfpL3HXfX1IDNXaaTWjKkEJLQz
GRucnnDAuWluSIZq8r3m0G0OKBaAOOHVxRaR1uBI9bTJ9eJ6MH0wJbPZ1Y5c2OkJAzgrmi2hpRrC
UgoF49LdsKy3dBqe6Cqy/5GD4O2ybOcoy3v2mfIQp2DBDCvgZ+lRZ13MtQF/aEvlzQBiQd4Saqx9
305eX9r6yJOi3uMU5zLJSKA5RHRfhIPEQJltsr75MGNLDmr9AC5e1nPobBjM5cNZQwsOupa8W4Mz
HYiP0/HT5JQF1eitrkJ3SaMPcm0E84081Rwx8WgtCTcn9kySThxuVXxZPDqcGGRBYkYzKX+iT++r
BL1SHMEgYbxxpmOhwXVLZ3muvjbi6aiNnFqTXyakYLo1aFRiMIMvrA8yxHcjRCa2Fb1xS6hQnV3Q
uZ9803Ed+t7gZPwQesv+uHBH+h/L5atYlOYnQl5B0rdHe+ia1is6U6p9ZH/FNL/b1DmxfG3uk2tf
/p0s+f6lZivFHxOGaGR4oF5AbI7X5ZfTUG/fhiSdsffvM9igC8daK8LD+YElOUBixMZRpDEixyjq
SrGAknyc3/UXArOxbLXBQRaP2r6sUV1qtds+EYyyJYImnMVVjv5/9rEP/WxTegBz565R7ReY7VRh
i8mdwSADw4aM7g5RZKVjM3lDIefjBMXUQ/S4OUMBXt1P6Hwn31A5b9+Ow1kesayqBRNuRjulwutK
DtHEg1xWVQe7luP9OfdPz0nsv1SICxoPy9qnRyrdLTa3WaKM89fOsHJVhc91EySGUV99gpXW8gxL
4HHsWVPiPqWgKoSw2O62oRb0bjp62MLzs2ZgZ2rj6aq94y8UlXwYv16TM6+N/6QSzer0xcn+RK/c
LOn4grnV/J4LRfVApo9QzqyvGkv1but+DnIYxaON8qwa7QiTZ6f0BzrS20JAXIv8pm1xO1sbUqAl
A00pd0BfW8ddO6yEUf+0SmCl/ow4Fae1sqJJz9HSYDMOXDE9fcdHFUakMNjEqDkOotdVKk7xkID2
jMhEHATvFWa9Oc1svr+2X7aOwx8hlAmHU5nzb6HDQstlBM/GI2vwO0jsn0/5yBip6t4V5DyXwOVx
jJHyHLX/5aqFAW6WqwlJtkpkJDBqz8cYmjLL+X7q1Zs+TrwJSfC9kY+ZHZ1CU9h5OLXUKb3CgjCs
RNhVyvgx4LBkD4Thbh7eqL//cDy8ENNIP7Vun/FD/I/RsMr+umk3K6oto7qmVmW1k+0/d67V116M
8FtVtXILV0p6J1Jx71ROfatwKzH4HcR6+O4rczPJeE8xGIi9yP2TqgwNOs+MY8U7lWEdduG6/4Dt
th0StADoG+UuLx6/VUGGyJWZ0tofIrVCvRLuUG8XqOGKO/uMhl4gpPbhWEOQ/Pjy6dOQ2oijUWtB
r21oF4abKCwH+dmLze6cYIiE/bN3QGOOGn05DqKEXAx2bo/1vJmixTcDPmi9Vtys1F1VGvazmq6s
N/aE9/4GffmUKLAmebsspYve4YRgN8GeY4qLnWudrbkF/4YTZ4eJi/MsdyYF09Co22bDMcE1cyyu
qOQOovEF6Ox5J5znua52xSvkvl6hQ66GglzY6Z7JXcjr+/8MjxDvODPgEmuUiwzUHwTymGlet383
TMlVIQPmqR036tQLtHcRHkBTNPTMjbI3fjkTTCiw3BTnuy52L5n4pzC1COJLJeFWwQV7pBZctBIU
zdko7eaX0h8/HJdrA/pbCDZkKS0UbZgJ/8rLjidwEPpbjnugOa/DCjrkpx8OZ4eprB2KuxSbq+cM
0lFEVdMYEz30IvEfMuaN+27yxtA/Lu/uFax5OANtxkYI4NLA65uCsmnOwXIJVwkgYZuPsuah56wj
8CEOHmaoO/nHKKPx13rklOWvMKVVRebYvDsCCiRaHkYYrJFQ2GTI8rGNBCNKiOXafzSxKDnErSOI
9FScybqeGShEc8Fps0Y00YybBH4z2UesAB5NFrR1Xe06OEat1RZ85mq2T2DDiv8RIxtABBeevPW6
CUK9Or9yiPha2ctg6/tkqnAC/t0qNusp9om8LlmwIRrGBuWcO+F0vsreN4XcEXyeuNOSZ0zPBP/o
Fd0mgRt/s7iUhY0+ouAMQhyu+YHVdmaW1AfU4OhwhNKJESz/0OcDuirZmX/JPmL2YhBIkQejDMe+
3aXhWpa40bp2JaCwvOHQuR4jK7zOjgoy5I/J8ukTpQzPHEF6skyIYf2CHVCZ+BQAyrbKRy6TzSNz
viQ0homYnyRmaPHhEUQZNxkxZarhuAudxytlTn1/1G/IKkhG9a/p8mk5e1ePHZ2MY4r2F1YFScWl
4LwlcqoELXvz7s5mwi82akrUYptn6olHMvMxK573C63M5Z1y/scr+FDiEDxb6o7px5Jb/gDN6vad
IuHdVvxtnbGXMMCQ0kngLTxvn/V2YDjWq4sZRHw+sQ1SclBsvl5X2+YRBKAGBDDpHDO2veEE/Fva
RK0/r6Oq6/j5ZxnH0Azh7/tpBSZx9ApuqiTZruNQSk+eidFdxPyAeIkm4zaLigcNEIl7OgRMZpfS
OvO35HgT3N49DjyYA4wX9InfXTdp1o4lfUcsHop0XSHqwoLls1Fn6H57lbi6OKWfuyPYfZO2d1Uv
8gAOUDsxSL/Zplak7F6+z8IqXps0fR1qjG0B6ABKX+ibcky+3WNy5g2e33gkDOGkKf6xPhCeQXuO
JyZ5d4IFpRmLiLUsiHcYOD1Jb6QsTzOrOgEL+Vfm8R7w3wmirXD1FWIiGUSBUj1PMrZHPsgLKV6A
VsYQCOschaR6KxxwXYfJasj3Y7UaUqwjQTZ7pjmbmm9xN/d1C+hWtW/T9FO8O4AQv8xbihSKhAHG
98L8srEewlmwt0tReeehQHRsceqke+VVTJ79Y2wYNyakPBsicNEUo6fsUN9qfSjk63LVHKoVu0ga
vvaIwbP3YDC5mrUzSEWnJRNDXRaCZ5peB0XAslMxxueIzqS4b9dUAUqmKmaXNFMhN5hzEFzVXWXW
YGkA+uzZNw5jPkCf4KyP944CB/PuEi1nZN7HIXztEPiA91PtyV2D/STVyICtA21BWrerUu5dguZ5
Ynt7QjawSYSRHnVu4D1I52q5EqtQR8Y2/i7Kps+zjidooAUG8/mjwvwKBmiWVNxL+oTVOmyvA2Ii
cxhJK0iCpn9Z6FAvvHDXHlgRQCmnXF5vbHGnlQ14qgZ+/Nn3fkfVG80Pp+pF7aMxPi73QAV/k1Bw
L1pX/ilLMj/pagQ+XIZ4k6D4X4PitFEByvGOZjtYM20p35/99Vxk1ojn6htCfwh+oBumHOWpVmJg
KAt+2ZztyOiIEa6U6Inl8hViPjBOm5akpgRBPEnnzFA9qsNu6XHojcosCbLl/hCzwUIRv1O76e/t
jc9LPy3jHJEKAvKiK+d3ro36v+duzxFEkniEWHRsLrqyf5QKkA1zha62to31atx6XIc6r1CfnQTU
QdJQIDpF+MkfY4YvQzeZmM06lwh5Ct9zRxr9JbqhjS32RQfCQUC+L0SeJcSBZODQtv+MBgk31MdX
j9bNiHudraVXAG+eaq318gFrygCiy36cBCSNmJotXENyTC9232Uu7NSlwIk0FXOwIODvcDAbLXJ+
T+A1foxIyoC0XUOWqeSDyTm/izJUQaLKyaXyfepmxYC/11R7TvRxqjacJmng+fzOnSuXiOSsdmL5
59A1A/raDvgiAwPd8I9Urp3ORhKcsZo6LVnofmWYBGXrO8hatJjvNKH9AA8XIo5AgBk0bNreqFq4
+KhHpxckqLh9MpTR4tPUmV+qT72pB62ENU7ClDj6VYG3M1u8ypZH7Yi3KPZpVIGnlJW716sjhPXW
2OV5yOY2wpFWr3GikN7TIivp32fH3LMu30MSZatBjzX3bmRgbSzeyZ9CJ3KoHDQbFBwdFoi8MePh
FpTUdaeIKmdEf4oJKqC9b+6wPyO+S9Ieg/Sf+RfxiqydTxkiWs0nWCxfBKVcAWx21QKGdq9K8IHe
xsEOY741yGMUvWTFr0ts2dF3XqcWJQzfw/20URQNeFgqFmdzysfrPocFPmhS4lmNgAqmv5lWMSN1
RZ29WqBgH1AkQBwt5H5kKtONAzdJKLTXxJkk6agjbXytV9U7PakFuIMdhBm7iXp5PA4vpPNNVqw+
Ve9+E2omUTxUXcTr2BnUH2Sy5mjrdQpNrz0Iy8F8sr8PJB6MtdtmvjyV2X51yA4HSpfonEBdZ0W7
/FV1kMht99u0rJZkannGbheXsOczTZlZpQ9TsisetM4DVhJVphjje0hw6lB0tL+fxjuCEG8yZuu6
imD8DJk98lOkejVoGlPLNNNyIbQQP1ALwCpsVWaI8+041PijdOLsRU70TneE/HXSpapjRpx+yhM0
RdJN02LjHuWual9mRigc3KJzcg9sdURlZpa+JTNbF0VB3gIkqTIBBU559EHpmpQW8bWdePXLblNq
sHRaQJhwcy4SxKpstO/p+3gaTKBgznM5X8friQUqxPiU3OUgdhJpjhIDRItH4zDaUtWtXyjXgeEu
2NRnelvheRyWYnzPitd6ktIF8Dl9GiP6rRfAkAGajIYuHjz93gECAuPk1jdT5QY8Pmn1F+7WegC+
G+wgR5bcZ6xYiasssxoFmeK0flmcgKsM5H8rRU2zlHAHoQG1qWVMBdNGs7Gy3yGeUl1J3Bde2JJg
zW1sxqnpXjiOctd+2yzwwNfKC7LrAdQyvSq/vH3GYmpofc0cbrMZn6VGAR8+Jfi2LybwGEPiiRmx
+bZRcpByeZid68XPRFOyqO1C4WddgvWtffNbeo3T1WVcHfU8zG24WTx2t4VDNUmgmuocCEp8K6by
+iixXLeAKNN2dhSXBebjpAmPM9ZiaUKIf+8Tv2mc57at5GxPZFgM7N5v0avgX/HXbvowoT3qVkT4
ZBImu7puC2yjYBjvVOiC/LppQnMeqIebBFvdIo9WauvWc3ikx/9aHATqsDdyObET/1/Mqs3ZWfCR
7Fztf7zltadd7cPhohWZetB6BjRSSYc0XVTT9Ts1j3Y93CngLwlgM/wey+EK/X9ANUHTQEG/4FCa
bWZidjpRGTYjKcdb4khUQ8ZarbDNBhxPORLWf0C9Pgz/ALUlloGj97ecJIL5iwGaW/zJec0oCvuk
DxtbxobOwmo4pWS3s7QrRcYDhICAtooyNpYoaXiOdJmist0zeysD9bI/LgSybAbqniZwPHd8Prlo
4ytN2ke2OV5IYd57zhdScK4MruS+nGBpjuGlhWhRpIgRXVybtVIczMXJVRU96mrw/w/XgLnhIRdn
GaBA2Ce9tDTOVdbHgCDvHBldRx+TQ2YWXujSR9Mc6UcpNBAskwuxewZtexJT0GOOdCccV2ySwRr6
EF0knRrOEvknMYx3sCXhpdSQ0foOC7nitu97zJZ8tlLa+ShKB/Z91bG3cOVikSLzHBG1f2FV7OkJ
FUOxemtJfWrcsOnoIvus26+SB1+CfY2p54YVksnOSPmIca1CCT25wDfo+UNgGeU3oCeTNRZiZVMI
C+IeMZNdXZcvLbbsJsMViQJrgLYjIV+atEgsheJpalardSvhExocrHS5h2ofpjnWXcFLqwqexUkT
d62HyVQlo+f8GXJQvhN/GD1bxvHDuaBdaYI0qze6wSgEAqMKa+SxZ02n1v3U4DPcpZMLmSIUn0PB
bzp2Mg7986Dc98m0hSE94dOTAGSYFq0CjO0yZQwoNPv2I7R+rXXH4ArC+/gSkSk9OGhAU9aiOnSe
T21F6F/vSJAP6RaGUyvAy40IRwSkC/gFvdryfKAikdwPIsQwbTJ4TGWs3M2St+dhwP1p4XZJNHVv
3l+vOVplbzwEbJA20PqVayw/CrZHkSbPQo68TE2yhWLvxtHViKOkNAuH/nIvOS+uSetGfm9B59cU
DAG9gJSpvGFP+RTlcRZHpTbYiuGWTO/sOy/H776RRb4PVot49ygZ1xpXULolQobtSHn1UI6YS8Vk
HsHxtf30VkrRL429OEud2uCpEQpmeY17bJGMIWdsqXENl4XDBZXQVwhfBHG8+N0MoFffzu08EYjR
oMG60CHFt3qABMlT71pTu5aEYXhpqK/9wAlYxePTj4O5Ib0V2eo9DTVHll5mB87dxRTxNKj4/PAK
5WkF4GtvZw/VFLJDsP3roC6oH4vpVCP6Od8pYQMukW2ipVtXUWKU7SsBXzqZhaKB1zK/Y9Sae4Zi
VT5v7/Y42RvuLCwKZkJIL9GoZGa8obj3/1sSaWDrtem7V5Pc4Q8MKdyCO0D8X6YWZhPVVPv99jv5
m7AOWWFYYQbVc4QJ4Nx4jtu3twTs9D9NUXc/DfEGJzLFXczVB6c4gm+lyPdzr+/dUHmovh/evr59
vmDA/QBI5vjjqsW2GSkRovjml+YbrRENfrBL2pbQL4J2Ep+rBcemJIzQuMoybce1LOzK8+nGS6OW
XBCctSi65lnZz1VXlSQoJWDd114Qf2QfyhCEy7O6Mw6ozkXKn/uTihnmQ9n8dIpCk0TS2LmkC+nU
TJmmAaegN5luHLzuCSJXm8fRJ+IBMQyuXv7SAPDYSWDMU6jKW20QfmrWEhBtVYdPYKqh/X56nNQ1
tqLDwWUqHDCK5rtTCXSJ2MlbgvRT/ZPRmuUgzG5Hr9mVXolECfbFtbltkGDDSgr7Q9VamGKQLMFn
FLH6xH7+iJm1u3Zwxw9INXAL6DY9ArW+0ltq2/gB/Hp1MSUJrO9+XyY2ii4X7rD0WhXzsxWmUn/8
j4NuFWeaLjpSqsC4GQxaNN6ehEFTDUuxOvfH/OcpfFKcHwwLdfqAXVOh6ukZQmxHToC1M2E7MWvY
gmHF5XCSNFhfe16adx+9rUO20AfCpKeIZn4QxDs7X+SbHMOj/YWgHtu2RSs29KO57PDR/zzNhr2C
FJWwxFCa+pbngNK++F7+A7I4yEHvKDJHTBGLw99G3M8V3VFdpZ83Uob37hlqGBgXqDEK8dXvfPHz
Y0x4UMHCIi7WNIH22VmEySPFj2yal+ccZ1bbpM2KaTWOK0932lxqoiMVJMrNzrFZvzuVyz3Eu+8N
r6G44F+t4GWOavFpHxpRmWjnHVmKpiMn5hVXw/1QNC4W2Sgc7OQZuBrosVgx5VuDIK4hwIuypiTK
5jwAs/avCzCYCz9QiXKoM8+/nUPR2feRYSRlsRtWjMxh5Slgs6y1ViT68RTRsRNFa07nNktzEPoW
EniJ+rSj17+cukOhoxDzRB+492FMyf12LEWq/yUjtLevd3lwvwgx1JOLWIZqGftTEtHH3QPCoq5/
rrKn35Qcgc5zIwvNc9NRDzAiXY5CwrTszspMtGwHE9anTaPfl/49Bpkz9V70U3D5+Lnyd/x2OrJq
7pXmEfD7frBitbcs8Aa+CWrYSQf26oBg+hmyyOt+6TeXH+B9tzz+zRFwXCP9UHTJ2B+k55iTFtDG
1Np0tXvacYlqqYrsBH2WYJzlrNkLdHmjrsv7PMtsuTsf1FTBnoxdsVlb7m1Vi6g6b1eAwbXNkx4C
IPbzw6n/xWvozyQHxHyTPuapWIVvWjIv/LVZdWMHOYklPDXG/Egwh6MYwEr6N5UUUicSTs5g7LEj
5AiGvGqDr1Vk4BF6IGQ0dzW+sC+6Hd3cnyAv9otQTk0Fcjf5nY3vWnTGy2Tmp9+P04PNEQNaI0Vc
77nNl8ut7YHsUUmV6P5lVIomHHb0r5/0jCVfeNQGm2ApExIpL8smg3PabOCqAXitp5orKP8xRDnY
crAs2sXL0pSLAQqIcC0B1j8et7qJggcluTUoyn7XrCUq7uHH4dRULwtxI/cJvBI1Cx1CYXrRpXbY
J39YyC3JH/FYuSnkrbY326JvfhwVi5EzEOhdyAOsKE0/2b5AugtzFc1osj/bUCjMgawxkhPveRGP
zilgPAc+bJECd9cml9xCPTN/Vhw4KRX2SISV1nYwuwZCX65yL9eObXOzG/BA68sXIvtqNH+pupR9
qr9tSM+aua6GZU2nhzqzT62KFmNQgJUwaR4WZ6Nc1w1E3oI4UHhepz7SeIVUyTMcUSPNTlstnU6s
2Vk9OLD6CKVTnTbXaxyP+OsDrlNKMUYgcr2rteZyRKcTzyiRuZP3FURTT3anrnhdJaez//DPQuLj
xTlnsH7j2zea/59Bj4lTLqtVeurKJ9Qyvzs2/Y2P5YakFyeCJ/nTuKUNi0HwavSokY8uEUd0/Ie9
ipBLUJNAB7ml+flTaL45vkW33aK/RqU+SgEx9AGVY2GCv1I3WmtmayjGazqEx/WQKg5IjOeuvplV
+e1/GLptFXXWTaFP4deWaJJWTIZckSUvLFFiXC3s5mWBBb0VEuQ8NPD/q6GoZEjO/lGtQzY5Xhff
RZR31y6o3phtET5E4etaAAdOxxTid9FHnaPTbbO/ZQSiskE8QuqCMfvl70eAc/bNE61VBUKorkNB
MgiYPqVFw8aJY9M8gl0SPclYAQv1cfkOzYebE1DYthRPCgrxaMIOerozcabgJQR2hUD+90zkOyYq
ObzgjcLWefuZgYmcn8n64BCZno70hXckP8ZMUv48BHnxVNjSoq4AniU3iU1Op8iVpEEq9ASKGFD3
+ZSow3fCHXobBIipES4RZ4D68cjaK3CCj3Af+6a4sk8+qN0nGBHvlNJi8dBjlVojaCVR6CxC9uAO
/PBvfcuIpAirlPPdpqta0iPYrGJ6iEeEsl3Yqy7fqmFKIe0BcWvyBrC+t5/d8r/IE2j1iz/jy/zA
C6i+1hFxgJUqUDWfklnuUEdhkm67wBW67Dd96ssEeLHXwJNb0G3oj/jYtqwtDSdtDnzsZiWotphw
gXHHwQIXDD+yx6f0E4cZvz8OGXH8pXFgrYu4D0Cg2QFtZsOmi4FILcn5hfAIm7yVIrKkUoAUYU/Q
fJwMuhmy3wTw3zmnlq8aCQYm15sBCDDIOEMOXJQUcB/G04w7kfPq6AqwH3fcMxIPppHdfHvjs/fL
0SjS84b+LpbTyisSaZGhG42VqIZnkI6jLWJcsu25xcgcf58UKmHoqb5zVICsbIv+xGGgacvq7Xf4
gj1nMsS8U1sQju8Br8uEcw3cFZCrFPG3a0ZD3lpXwa+YV1ATQzF4L1twnaerkA9DunalZEc4qMZl
PmSGpk71/w7djAbj5du+WJzkMU3UUC+DDIe6j3daliMWx/ipSQu0TZ2AThfvprTDQl8GwEc4Hjww
VlHpwoO3ihpQ6KI0YFKC9ErfYTihVuauhgW4HKjAYoB3SrPDTfA33Q/+nuPlneKboyR9hDnZoH1D
Ku6ChGloMyxUn6gzfGTIoPJuAhQ31Vgh4q9HDwVK898hApJ565ONQ9zAegu4YBhU7V8FDwISMtDD
nwlaaNso+Qkv+pR7BJ0lHJ76r82zdn7QjrqNJl+oR6h7fPm4ZXey0Z6ZTOIKLDPepTAMb7PzFjzf
4j2CRE9pUxIUBNXNaoKFvHCQhM4hWXh5r+kdUah4y47wvwIIpwFXU7OkPKT1OnnndQ/A2bLFwZH+
DQsgfrdnlbidSjiv4GZxKdkDWwcA/ejtLD6fp1KQLLlr59RJ+ECnw7cKeGFdEL9FtV08vi30qufz
qCuHlyks1HRfusmdUSzkF9rWwuk2P1a1ZzDLy31Hzp1wuUtodrrVFTWtESC4een4hDGnbee/IqV3
PFKgvcOE0aOlRJOiJhgp+o3reudjBGljin0uPv7tjZHVD0uLyv8zjmzVSatEbmKIlIgaicdkhA16
+NtmzSyvdKPEQPRjOY2KtlI8v3DzKb6pgqPDYfYbLjc3vqBDeiqYHoS3hXKwnLwdnct/CjC48OEk
dGRqMQeeXqxLEq4W3oI+mbX8YqxKy7F6IKbL2SXYHZbkM+blR95QxQaiegUInPrCxYaRw9iKVO7c
hk2o9Gk7c2X1fEs0AZwQGRwl0+eguajQ0cTvWOQc4xtfowTKgOcJaOJnGUujcM8K+Ngi2RTfRgNy
v3ziT8qR/Jyl7P1z+36j0UJO77uURH6ymySjBeduJvi9Sn/zlEanxwy/S9MfbrngGz0/pWN4u9xd
hUrnN411TlXC7tIOqerdWgtPhXz1SLTD0xbuKt5uLBeDGB3wlXRvDY6Fgx6eqY6Xxn9mt8beMgkl
kSyfEN9cCNPcG9KFzHxprxDVpMDSdMZHA9cj78YlzXV1HXtgGYGuDTWHdAqwWZgyQ68PjXchA9yY
fCWbMCKkY/fKYUpZRQLqo7QRdkaxiK8ZaJPbiqB9Xh2r6iMs8YmqhKt/5QCd0VCnaMJMFy7T27Tw
g2sBQ3BmvX8NkvLU05uGyb3mOZk5SeXVe0rntIshoj+MG9o6nzPLeBKilR1bQPcQydsknvYRvQPb
2Zp7qjsYijaBKniEybsQMT0ZIa2UxoxhXZmvG12X974Ze1CaP0JK5yZfqI/uHp7TUMSnpHjE98VH
yfu8b662iCWY7hrhPv4jp1DpIuH4+yI7HQs6UslmxZD2jwoaS/f+Muq4j1HX8PQLExxau7THvUIJ
bsmn9ObRqhPsQ7nywyAp6UocvFvAjwBy0UVQj///qr2RDUFl2z/nm4gr4JK1sy2weYdwCSlhUbcW
o/+RcLfDpuTOq9t3oPpVhqYNbP4uTOVzxCanfZ2kz6OoAnerabZw8PB0hP8z84C4/WEVBon40sh5
8X49/yl8N2qUDskLY+h5XvSMFMv7FkzdVJWfm/feSytK9TCqnYCr9TKfiLipNrTUxYNw9uuLgADM
fG03MnyXEmSryLDOvsl+tsaFTzaIuQGnk344xINw8QzVsI8g6bVih3zN60BvVdlp5zSIN5DoKO8j
04RGFcaxdxWuCt9ST2bGr2SAFthS51sU5W59jitnAxChQTskEx+p2mw1PFMTjaKVSBMyQvm76Bkw
x3zGpSdzPBoqhWRNbBj1LB2ZW8X8P9YIvgsmvu+1iHmOb7YT/qM2R/AMS2RGwCRV04RGap5h8qGD
96SNmkjdhEpxsTx39fCySwWYJ+WdgKqqVGAXjoY/xaFDiV9cf/EskBTAd3r00U7U1aK/TmSClwSO
1QAHTL+aRy6JnA336PHiDDMkpT7PRMo5+A6P2mnyTqW8LQQpQAobaq8RrlDMqzMJWjxaRuSP7URy
IPNoEzvo7rnEqJMY5pHu1NIa/mw89oKzBc3CgdkQFNVOjSq740wTMc8YLYb801fbViRj4air+4Ll
wVpsQY/BPAJ8D3vN9kSTtmWo9xkQ4LJHiw//+dHF1KYHkNTGtvoQoFh2J/34ZamkE6Vp5gAQ46Vy
8Rtn0q+zGCOzrdQ3hHRV5noJNR2EaZT4xBogYjPdeDQm/hNEbJmda9WExLlWrHno90th15gQcfnh
J2moNF/G1TIrSJskiow92+4KvtMwcxoDrHHRB1Z1Eewo/cIn39BgbVLyL5jYgNhTQ9pyezJ7JQCX
Nb+u7Y/j2NLVMt2+TrnmrPcACzNJkoOCjzayXijmIQu6W8nbsuc2bOK6Hb62BXJxilzJAfM9S5lo
yoIqmZ8vgPXPQPl22yZKmbgg1aVYhf/0nlk2leyHUug49j6ZUbtPl6tCDsyw0VMX/I/Y/AFLxz7+
W2yMAjw9GQDSD0BU1JcJOFQVURNnOkBuwAyCdYDqVlJSmHEuwLSeG+iZcnaz1Bzo6CTsjhxWJeus
A/QjCz5iYrscQe1Wuf+jnKOW2Et4FBOxq+R5ioq4gQXfpudUOJ0NniDtNj6+S6ZQ5qTk2bj8Visj
+dw6O/8t7X1JY9JiW4BKT2gzs16jrGHMXFhgq90ZYPzovalsnluZCmjZZzeQ/aTlBBOkrqyqVJjZ
7kij972WYhr1D6TVFTODmpoYkUugIPLh4jToL7/OUnH2PKNEifEfYxQTLEqB1ZNT9vtDfvQsvP/Z
lx3yuMBVYHjvaKg1uwlFCr4M3GSmXhdugrzXiy83ulyJFLV7IU+/RNOhXdUKzh/IFxXhi/JC6DmG
iMf/egeH5UMXQeSnAF/iqf1cohH/98dIZnCav5c9v/dPkMvAjZa7eYZwnWJmZji4FRjTUbOensu8
q7nV4E3pOBedMucYXtawkBddiaEK+n3C+J9pEX5M7muS5y4QRevEL4KvpxTT5V3YNSSnwPg+lCRy
NGgF5Bdpb3axrtKVW5RV0szsIm7L8FKAJlJaR8GTP+hWZcBG9NHPNCnqJQjHpGYO3WWtmPXeNLiL
cMEehR4jjFpno4MKmZHRaP4Ibvm4qbB7VkSbHda0En+6jcRYkrI7gy6IXQKqBOOUFIvbKfBuOIWp
A7m+uPsR6ljxMxJUadV1sWEY3jQ/8+JS0XF0nH0Ce8KSALdgOqnyDVSnpWOnlao3wNCTX93wZ9Rr
YwLbGrBzzmyTgNsCawY+E/oHD8ApG2Z5nc9hcl8TWuY38IiFlE90VdNI23r2/AQB2ftuQJOXVT3s
MoODk4ARJqGW8stWiygbJD+RiSmgM6qltCRTz9Kz7BVGzh/2bGsu6Q3B23BEbUlj7nNfCdT5197I
kv1B+WG123zMgp2MfQDDueP3eoNaGGj0OgMDMtXcviih3w5iQI8l0voheH4RuUP/GS4yWcXegmii
oYYEqKVE/MTp+xZ4yCeiGnE4TyR2AKK7P+fTuc5sZw/6IDD+dU9RNcJnuWeTtBAHrb4KEpgrYDj7
e64bCQ7JuH5M32rtf7ihrpANZkToWWqyt3V90tFW9mONZc7O3LTEAmAoGqFqYRUe3m5PryUM2byI
0DbB/MADI6Po3BG1VAJnAVekwCHiSV+lmZEUG0WW9b+leNjKCRg8Pb8oDa9dNYW63Br8uYm1o8pY
JDyGsR6M23lMjI8RVginzBZsw48CNWfF+DoWt4F8M6hQ8I1ddAUqyG9nifoGyq2mKPYlQUIh7Xpc
eUZYhMQVbOp/cwpmcpReihA0QtVE/Vcs3SAXN4y3Z/hLyjIu0fV088mL53rgS/rCH8Z12ZCSYeJ2
CakDUeVZOc2fq1HpcIe/UaG6Z22jbZLmzaLk/1IM2ekCaH9qb/h8zd8YD5DPkI6swmM9TsES1MxR
PQxY5JzLJCy5R88zXaw+gQ63Jexm5ODLfgx3QtE85B8NEOET1MzzoEQ0NNnWi+SOYz0QDUOHZTJ1
YNac79/R1ovq6EXuEXm8TXEAJtjmPs0vo9iO/sssbLbYEgQDBa55482qye399OJlh+RLTV4LKVBW
j+3ZAR1ZVS4Ejzz9omgrIaCKN4gwH5XP7+9z7fb5N2mm51iKZDKnvTV7VqlW3lc3Z1+iLLqJh2gS
IfIjyrdwRKinA7WmNDGuLjyxLP2tG8sEpasZm1oLGUhdeZlgu5wgSYhLNPXEt+MWZrDNnun/mebH
nmbgCwOkNStfyn8HFSzDKsBlFICt3pBmD1AKqso+d59enw7Nc9gqgdogdNh9hd0erNUT6sR+oAd5
nCMsW5mJkToN/u14aqDBWVTmxHPi8T/XMITWHnRdMRxebNyEiGYR8xoKJAg0GcUko9KDKxXmU9YH
bCC3eeeYOVHxOnMMyIui3O2RpOBd+KfL/lVKIXOHvinesiHMf/MN2zC/CjF1b6nebe6WOX49O2Ud
FhkyxmfxAsY50MUsh8upGXxAIIg+3+IsW3Ez2israrCV17m5xyb8UWJNZvtxCHiQ2nK5gdBIptaf
MmsbNzBVSSvbsuTJXstDIWJDkfPv06SjaPjtrYpgmn/8NudqkNbCvPQOxI9lIThqikuWA2BjUJNK
AJODiiYbyNj83la2pWFHSx3WSWuZ3NMRryCMK2GP5Y23A2lRVunkY/dchqVO1JR0KjT/cZ4C1wHF
JCTFvQdScf/wJ6VNzPgncWcVIzxV7GejbqwoLzYtQslRm7cZv7mCtnFqWy8r3NZVzO6ZCKdAYvFW
NrI4pzvTgMP3dFw5gAWwmiiP1yTRLYv3XlMZ/v1BOUoMDegsgC70VFkL0sFOATNhVFZMFktMCO9h
0BEDFzz4iVfWBmmXiHUP6guAMRLf0VSMLLplaxZl0uGoZ9wK1GDP3hylrvkf3EmlABpcHP/GcLDY
5URt4eVAqFBPoRTMPiCYzp+C+NCz3EW6oDuc3c0eDjlz8zeUYQyQLPPALE6Z+IDG2O0Hs+x17a4b
eIcXv6uAbNZ3Q0yr7vjIvynIwYTm9REJDgChCUZYWcoS1xKnSho1rPkQJSEaZxENtn3wEvqQk6yZ
WkaqjAJgUi8tIyD3z70PStGyC0+Fma/yBxw96wNGW/YlfG1z03e2qXF32ZusfepyhVhCl0VzOS9G
iqXXiKGrlIQiNIZVlJBxD4DXCax//09AkXONgeNbDvKeZlXdR8TcJxdTQXXXRAmLiRZ2wDqv9PXD
oGwpqD9vYCDRcIcOsSprnRbtUZmLiv6ikroHDxPHLgiWRbtZu/Yjsno1rcC2fRa03i/l6gjmpmxm
i45LTUzz1h8jrVrh4xl35So5NYb6adRpay5jxoFy4Pe76P4ouPrEQfC+zIX6l/TUDDsP1Bl7qiTf
QSf0aZBgDM4IWkm34qVg4WNjIZPq2rmbSIL0a3yQxMx7X7oH9pWd462yHfFtSDi+nboMtHUEdhLX
tBTLJGIRajBLYk1kfN3lzY7JVNVUlfvg2gxfVMQWj9kgtubIG6eXoWsIfeueQZID9r9DkR8MyZzq
QawANSFDTF0anavVGF5K5V0TU8tRC/I5YX+4zAGz25trR8LOe1yGdQrkJugQNl+au8aySVrpFTO5
brTT4AaU/60vW983wTHB880h+xb9eTVP0QMrHMcSJYBezscw2M1bmAD0+e9+/gb0LKQTDdUjUdZK
s843RttEJPDlm7zhh73EaDR32XMZAfWVWO/KJTt5kVh25VySzzNGJfa37VQ0Wq1kwQoTu0zc9v/6
vD6kIyztiBOGZ4q9/28BBtkYLgKzf5Gpv+Vjf3+op5GO42IAn5zyL7MgseztMJwaPSj2WpPSXco7
SnXSWIGIhtLqyPPQjho2lJ2LqdIZWCPsJTYuQ+GEEGRbXrIVFpyJM5vVDwAdks59GO3sF76RpvLx
T2AAGEeJ6saCllRLkKmqqmMWdtCUwVruirXA+nLxKMp0rd3Oz44S6WgmZduMVWfxPA4dU9d8sAHe
SOhOz/BOrlAsM1LXn43YL6s7K0Qzqz3J9AYRCY32LHhJ+blq7VmjIgLeSJ+TgBzNcDjxbNTU5XX8
3d3dIH3QZV8IuOry/IR/trsnh4YIR2xz4FSycs7ER7OC3v7DurBGCpcg0Q5gqWIYGGeVVsz5MjF5
KRnaQK83eTntIaI5s7Jx3UJGdNpnVItg7iS7bXvnHCnI5HAKKKDkQR6G2GR4if+gMWZJkCVNKh+8
uHTYE8WuqQR4ck0Ne1T9tcJgO4OZJH4dfsZj44pCfOoHbPokhFCfrAaodqNXFFXwTty97yZMpjS9
578v7CWNlNuy74d9/msYPvC+0vkXE8pPki+A9XlFFoqLB2OLVmaGQDpkxghc9aWltYZWTfEKGMs+
n0RbI8gvUiv7l2PsN1X3yRursznURf7r688ceQb2JTgz/mHmhJll+SD8DENfdmgZVzzwbWUtzh6D
dkNuc5LSI6ppjFrPP52pdFu+lSWmsmAEIXxXPXXjT91wcW6cWXWjwltGm2lEb17z1bh6OW+JNEIP
P9qoBDD5GYJuJqhSBRiKLs2OIVDrs3YaqKRG3vwCfhXYv0UPsKiXmUfv3Ij2ORLkSx01G6ME9Q4W
C5W/eMWQMBKCF6gY0R41cweI1NhoJdHdkGcXQ9+MQiM2eBKeiZhiQsZsnlbca3P99DEzXtEcrmBv
Nw+3EOKfeH4AjGabHThxSwQUbHz96fNTx2ojsEwQdI1A2/BCy9rnIdFT52RhewrSLstka7E2KFs5
MOkFideGJ/P5AUzrZqfNdfBtUXZ3Wr29/W9NvoAP1fjkkR+opfvvtfneUdLhz+XkT6JUrtagfHP1
VL54I7KSprW8HPvzdFDOzHJqkBigNwGnudQB6rlzTr+LVcq3aNGBq1+zyzhpZFvm2dMnnvN5rnKR
5K65UZ3dJldaVy8SwyEjFMy3+gLAAy7eCYG3s6vZzHbUtBzLIpMNEn0ZZDxQro7fLVd2Voy6lfME
cGPMzbTmeg5OwtCn9VR2ocm5N9l4Si2DmUAkUm0CU9eAvEXwfp1Px/rU+FnaelirNURlBMl3TkOp
MQ7SgfULKaozjfZsZucF5zBMxcWEp74V6Yj5BryA6jxFq9CJXepYKYd7d/txqCDcoehBSsdBmeEC
U1lBmmgf1WIG5Vi11zEZsTpSYfnTPAItRLwmX3lubzG0tGmyWPFd6f42BWOpKRiQFTxZ2pIyk0+c
Kv1HybU0IWLEckN83KMprv6n2CIxNDP/eFAGuzYNBkUVQogckks91+33iBJ65tktOUMZ81i8Ao2W
yU9DeX2hfGLC9GuyVIH3ekDVTFw6nGL7ayGOrausav4faguUUcchrtv5sFrtH/4U6VFAcjF8K2/e
U+/tOr7L3dkbLIcy4qBJeWRwt4nS3qle6kvcivGeIpciQHEXllxPcbSxdmBfLIvXxXO4/TcCLgHS
M5bHBkvkAU3m/xUacSTPnqObPP6r/dOCBDxmjMI17gzdxRdNe6trRJGGzHUZhpi/qHyIMhTI85Io
uxA1zEIMG9O1eAc7tgLf5+g0wFitRO8RiJlRaA8k6xDCtiCesraPSn728kYeT5LIzWFjeLPG3myO
4y0f73Vxu82l1Ps80SVLKwaIMn7TJtwm1OycyjgzO5RInvld204iW6rR+bS6t8o7+qLTWYtgWnUc
k5yV+8Qav8aj7nqAon+lNa7HIhr5shVYkz5jf5fgxvXuzaBP1HeAOm871q5DJ14uJuSIE0527VSF
jkUNWAnnzuoCIQGFv8i4W08yJ40Ps/Fj2o30dbbjY3qAtBD6Qwky0oBpNBxBXm9IY/ocpP2LQ9n6
QRkSSfi/G3WpTfV8yRms7S6iRSG5spwTqiz8Jz+G84ypXfTasEeeJajitZVSIJDg3dLn6Vq9hFfE
FQPqiBJHABXy1X7G4y/OGfPGcX7EGQBvoZy05ZcBFNZy8h+Um/+zT1QikWR1GNetCxbEOXISvAPP
xsNwKk0UsTDG82Q7Te/0hQxyO9FtF9XeWASuO8KscDO/PA0c0LSDlW7SJQ4nS3z4drXSsRYaONd8
nODWa3/4O2BTZAmYZrwcMr03iy8hOhypYO0aPsupQ/FnUhZW15LhkbkPDWQWZkOGtIIyXLmI97Rq
hY/ooarkiqAbGWbwuirSUCMMsp46XpMuLPhO55TWe1PJ7OkHPxnWwd8WHsnSHjYtk0XKXBYS7hD0
olid+iSaAigyPDZq6lA5DTsWK3RA7PjDn55NB6cgFiozLjhavQ/AHkodDRviznmlqBaIuSoVbkiF
JoCDZleQX25wHryfphriGv6osGad1YeCsmjw9oYmSKw1IukYSZVprF89gc9Aw4rAffZZ9WWC/gGT
XaVpdzx2t9xZl1jce5cvrcGOhR8RKd4SCCMzO01PiBcc5YoAqlncxS8SJlqFI9FUjPAuHqxFHBRC
aKqZzAq1YGrTGU/JSa2sktmWyQqWL+PYc4LYB0ZT7aAvTqDJoHKqAijnn72BG+IopkaOkNubGFSx
FRP34Oww94poaG/6m6BzpYNGlSKTf6dYjYYNbbmIIQIQA1JQYLqilSlETmKpJXRvsX5vpWgV0/F3
FLIK+oP1iwM1RIdxTPE8XSiPm8d49gbUHnII8kbede/W3RTbrknQV54L/jFshOl9UcRTi4BkQnfo
yI2DbtP5/F0kyUGYmHquEP/z/aOSc9TWgp8j3cbYTmmfFwDYErLhMR1AN7zbb4bgsfV9bfwyF+bI
VygXc2+xNNaWuzoFrRQkQlnJhY1Rn/yU3xu/jBi9A2WSZc/WCVOvL4d7/EV2Q9vKZH+uRwkr7HMh
wH3iiOTEhYbbKsCIKXA6pGpJtNqf1wnyMwZAMM9ZhXW9xqqKMlxyk6uKYTsE/3Ikg/meIFTjYfhs
l+gm1gzULXZe/CuCnzO1yOlSMtZwdc0w3PIITYFogTWuHKEVoHPRTfPPbgnGHHe/qmB/e+j3mlCA
ZL2aYc06P7EJlFZr442G7Yno7YY0/G7mwwANGOT14qt9UtiHUby4fp4Bin88gQ+rkTODx7zDzy10
tCOBsW3zLvPNYgQPMJDyo1dold7Xg91YOGq5YYWFzbYNLG1uWfXuvxKuSiyqpkdcdK3WHl80vwRw
/xGpEXQ5lxs5ewwP0qfDCB1C/5ju6Zgl1MJvaTmPVVJLuDi6yBGBf/qtJHlFKNx8p/DvnpPgE8wq
1RAYHyY9/sJxlXXqnkkCGwfjpO0c27X6D8wxhgxx1BX/BUMWUbM4i4qSJ9GkQC79ZoLZlPfBlGxP
VPvOspzqYMRw3n60QWpl7T3LX/TKq3fBAMGMjwjc/csJ/9jQLG+uSR+ZNt8GbCNE3ivHKaiikkdq
UtXNjZN7M9W9N174wJcCUtN2d+LVugAbLoxLasGCFIKNU8aNLUIxOwcBcVHu0I3/x3RmmKB9Zr8p
FtyduFoZMQDRK9RX3USS2ovC5zPPt5w5pkUOLSL8z5bbt34UVbIuuN2HN/9y7591YRyG9XVXfR6M
TxKqlBp1qskmzX8CQFMHjLliogv+n9NnMOnmt2Nx5fcDV7QK2nHct4a8KSrGNI9zZwdOAp14C9ZN
BRkYOQZbCOUV3Oe44V3MvRTV1/kR7HWF2ggBYe6IgXdNPJX2q9cCSvrYdde0iRgmmBuEu86xkY2a
jGYc57Ms5cb5sDY5QYwzn/1HCS2OrcM5kBvUbc5ZsLrts59cZRyWehc2H6W+YJ+WUIgFCkznKoHm
aJIGBxuilUA0bI8uk/jYOP7vffXEqaKW41JcJGaaF+UU/OYsVyralWN9PeoZ4dfGx21NYPaFKHJB
ZBgwD32vVb/CQrXVlN/bXapt4xqAH/rgL4IUtxXNomAhlMW1ZUgcLlG3u67nKQc2lmqTfhVVEo1u
w6TAysdGlHRLiMP71OekImNmODixcL5TmQZZN4pNlsSyEDo5naoeym61KI6U/IyYEwylyXe7C+Hq
Z2PYXHf8GBEj3EUrXQ9mYIYOwP/1axYIq8YnnUZqpu72UhyNqaT2ijtN3yXrZ+5JGSPZepvM+xm7
NnFJtOECv2ATvr7E0XK1+lJhzIf26qGGgCgwyP83FAWY70IXMXQhiI/kNHyVKOi4DMSAgeiDhTjY
cDMK1Zk7skJm4U/cLdorJfVHldXcBVE+S+WzM9tunOiFql/SKaVpdhHt0/eFAx64r6zjzxnMcjVG
0+H5k86IQEQiIZLaUUjvzUxsHq9n8GluyR+ECh2pgmFTkJ6yFG0mn3OVhToBeXRkc7MJ0IxQ2g9C
oUifVlUMPJ2QL4rxN8Y8M23l7ttYYBl6hyeWt+IGSVcwDbvDKjltW8koUYCxTlPUxMnAnlpbfyRx
PvSg6HQRmUIz8p5GCC7R8xb7MwryVpKK/wYpG/Y0vTZ92QUeahMBhJhXafjT58pxoi08t5HMjSjG
pxyW54nIj4d+XClRQ9bkQOttWRrBhExQcVi5Fnrxd4T+5IdHQqYy8hsKR6b2ZrWyISGF5c+IZutE
HoEEeyurebVyXZ6cL5w9bKX0fvsna/zcx6kBRdrUZotcwhFM1RoAYfPubYkDgzBZnxKtUZOYnT95
sgSiR2TVEw/TTH9NR5n45zJZq48802ZSlMPtBh6ftofXgvaLGtqpREqPbOOViA9e+R1xO8yJO6ED
BnpSz+0Wfr2kM+yu5a+w5A0dDXC4mNlPG8xs4N29TvgQAmARfTEL6QzPyKp3cl3Y//7Ar5wiTmax
LRsEVaLcsExeqxH2/aUnElQkPADjBb9Bf+tcodqTCGzPgdvCDNxdi/qHqrmH+2ND/7/RBVLsuHvd
KfWf0nTnjuMXO3u3szyj6zy+o3yqLFMyvBhFO/wbocCmLKttZg3Ufj5BsHhgHK9KU/tRr7jrtVod
sSZLCSjFCu1a3IxUW/Dnpvc5asjRTMePf7uD7Owu5zHgG8MLbUndzLB4e8aQjPMxF+ZIXoQN4TtJ
LCERHSMJqU2rWxfhcJwGswlv0rqsOyyQOnmgmVz2z1YKEcPHNOWGFlBT2xXZRD3Nh2HrgyOVx4ca
yZILBS051Dg5wuG20o6vlcyJ/xG5XrzgLSFeVqyjZP+/dduv11tK7KgLvpdBd8xWVucoc17CxApS
rJP7j8zNUB+E6L9iWQ9WQqFR7yJJLtddDXK67/DVlDMsTIbxSGrgIZNzBlKXkv2gPtMlo8FmSv/j
qa/qKmssu8kswLqE3vYJahOxulj+C5ilAxniHXBtOMoX9DkLpPBVJ42GqepqOI50yHNr2+9k88eO
sPpjnlVByk07zUXFhqkCejGnM0u6RJ4Q3Kio28kCM8IFnY3MFdVj8d4LWLWrDkhsCs80Ka8A48yR
ART4M+AAxr+dkrcK40LKEVXRR9YVXoR5zV8HzdI63vXojfclsYIoDWz3G+P4nQS86bffCuxQDbXT
1arTkr+jnBvM0cAOq7N0ly/wzFmSRfVdEPEdH+4UVBg6tL6TD6qpHnueXdGcOtHr8z/ev6DQZIRu
+F8jshMvebG8kF7MW+5eCsG3J65e/yQqHgJRTPK3GOPEpAHShESSPYAwq/ZMhylHycIIkIGcRGeI
MfjUDbuOm7izNOWF10CSw5nmOmQ+NOgec5ENky/ONFi4XDZllipapd+Qhf7Q2WLkYg0UVcBU5Apz
46BgD0HTWhap3dexJp5q87qKYLz9q1vr3pV2K9jU79VZEWElANWaFB2zGw5aodqql9fUG1IRFKKC
0Uqby6rsJaxSgFpq3BagUugNiQmkB2a4WEu9eTqDHo96/eR04d6j7y0nNQUq0/f7c2Xs/yusSP2W
LL7Wr58iTbYNlSvMDx7OkjV0hEUYpWEU9AECdVnlZ/e+rvHPhsK8PlF3H283TIJD6Ya1ohPimbdx
8UO4v7jYTCO1yj9z3XzDd22gUpBt66gAKCljEG+7AwEEt+Pd1UEQOf8X1HLX9qusk9SAkPaXl/9l
/2diN6DOM3KhO4WXVU1v4e3l55FTTQHvhLSI2UIz41kMEtzvrUBlWc7k3HXoFAB2xdECMjSvVJJF
Nzajt6uwjDll7GGpgyDETxM9ch4eEqwkPmpsX+M3fqfyrVrJ/yRkA/XQGUFR3rhUcNN42zvGfq/c
Z90wq9L1EITjONQLY+zAGcsTRuDmzkmZNA34ZH4d9Yz5i2Dz1iJnahCtq4L6z6GR4aH2ix+a4SvP
2L6IU64vxKpjaj6uEcPiR2bYRwn9mOW7IO5M9RC7pkgqOClMUtN6Gaw+tEs9m9CWdWToL05Qv+du
9JGI/m2mftHPHtwC51GideIGffo0jFXdDWQPB6qyM9YHmBUtFK63fuCaQ0bSq9PMbo1IdphDK7K+
DFCY/Ov6ub8UgQJ3XP/I7Dgeqw6JiEn1tsTf1IoWZ3UthuyodRtHIBHCFZqaKUBteYUU28gTl2H/
Bv3Cw9+uJbJCfjqz+fQa+ZgyO/U3Krmwlokeyfv8ASZtW3FQmxZAHmBNC/Bn5qylDse7QmgvInFq
tNweLxvvABF+OCE4v17eoWEbJtyK7mQBJLUtlykV73fHEAajzPUvQmXlitftkeMNSuc3Ze+koWl3
9Gves1PDlhBqmPuCY+yuVxTNiX9N0wi0K2KFRwkdWwL7okFXc6KIX0B5sVCZvDgBx1ngr2Uwkhp0
l8TSuQ4ZDKaZXb+ADc3PQZDIgRd2vBrvo+Ucia599e5L5ofCn9W5HrZyb0iWvtOkGZHfVuh5dr32
SEtH7ATkPrqDel9R5ir6khUIy43Vf/22nGezHl5D/Fq/JCnEozEu1sX/KZEXmQEXDxjo5ou2wuAc
t52ZBkqtGLv+XXm5ZJrIQJAXzqgqQSfkOxJO4htT0c4FNKhHXw8/j43uUI44m02UT3Wut0cqs8BU
277Y6N7BZfZmco7chQs26QXLdlWcyDypI3mNMnErBLIRptw59d3e7jtbTxInHx0/7LK3/QGTRT/L
O+ZbmPcvh7UMjvu6EGhi/jWPFR54/fXGa6SKBtP2zXoGmuNdDZoopIzEq8Y5Dtfnf1tyG5ZVdwLa
JPQqRvERgzQkix48cUjNVQ5Tb1iVOkt3ZQOT6hB3jHyl7Zj6IDTeYqBaaDqWMbM/xXT1JKdNxRvW
zWcSL2O8olf/clnwqbWAlfsjd+jEO3mgtD4JIdJC74U9/qhnWVxeNbZ1qTfPp/4SmjRX74CivO+9
mm2RHCm8SeZ69hi2tOsycFBWQtHHdVdHq4ZFzh/u+n/BiwcFT4me2D9FGFlpEL6V3TrHZ1cxH0Lh
lexZNMAwTyamRuCBusFYKLcRR8zNscda796e5nXoWbzx8HN6hnQsMl/b75tAFKtzmLcrnqwW6Zyq
TcWHCJ/YmJPnaBVFA15iY/ioHLOdmsdsu6B+IYzY/361KzChCiWb4NARcjfW/nWxq2BDQujSVUWm
/zVTg2PSWveW4MUSvwEuVyTiX8OkVZ/WMELXe5P7gB1dFR9WJDnvRnunE6bCFsWHf+ubeyd0YYMg
aUEWR0xjy6iLkB/UpicfPDHwu/ZWcGBexqqIhk9tWQNrvUO5nwFx0lCfRyTJkQbaPZdctWNZ0M1R
QWbYyZOvSO3fnqKXDYxJ3sZUb8Kl4uXEU903X3nwKkkHkUjbIrvLDYi+OTZ/5vvQwwVAKKCh8hMF
gTOXNROPgcBG9bI3y0GODUslAX/HT280Rf49kCuRwbX7aO11GoIHuyFkOm6QCMDxV8wYe9o17JFW
9lhy6M0jE9YsobvHVEX6i1HL7rak9KHQNwXSERfVQchgKLV8oxQXAqmrhLSNoDnfpxxD/S/VJZPE
Bl3sNzxNuuoN723WJKbBZ27y01m2EPMwYnqEniAsEQLV0t9HieXSTW7bVCtccwEFwin+R1tcHWyd
U+BmIK7YUXmmpe4f4HClIXzIu2zgfMTaq89XsidwKsIxmDu9v6kdpAZlGZM9w4T6DWCa35iyckUQ
6oaX2/62gpSRjcfo9nslyj4qIAsZ1UBtzm/cqeod+E+4QwIk76mRaExfw2w/fET9+PzDqxPlgqJm
Oh4XN6reU6x8NbkJ7jNIKUVOZbGcEFSk/ASWV+OVpjLyCXpKjD1/JkWYHYKy+PQH9yaps04uABoE
irIGfnytxYrSKY9XAJcyc1cuu/SSrdy8n/vhXJ9m12mDv09sKp2zROE0HOm1ApIBaKr/6iJtg5Uc
WFGSgmNbWruSe6O0dv0t/Apx5TahXwhQ8/SUARIJYhbK6BMOm7lxnoapHM3qE7LJxTePBqRjUy0Z
tmzujxXF6uRPiXBc/VBgT9GCIxCNYqeE5esuOUveruhRVpC8AKGSUWhAopmHfHLf5b5pMf+Pq1tN
S4EciW3T1iHJSlX+YF8Wkw1DxWPm1JvvSDK4zVkkefIA6lhFuirm00+lf9A8seDWYxfqwIGKE7kw
kzeVC+7JeIx3OW+k4s9NJmQ1mAIM88kh/x8/221N7BHGS4kcrl0WvxtNHUefoUyrSNr3S6Eudvgq
iObLEFzYFKxGLMtpXrYHWzhQGHjGoTudISpxM+nD3uJDHCqPHNdzxe67Yi5hm1FxTCOwQUFUwmOT
pJpdJLgPkkP3ywOc+6Po404TGVgdXNpwZLqaEiKtfcinXcy92mDKz1ENm9GVRnceP7LXLJRfmHPf
lFLYdyZJOlJ8slOU9owax+PpiqFqmMdphEQFtptug3Vs8LoL7vQILyU6nPS+A0LOiUFPQDJQ0EfR
ep6ZGCnALOen02G43ZIvoP/++CRZudF8pY4dZgCxWIdlt0GdJmgF9ixuCvCbjz/dwa6f/bsb82NI
83xRR8mFSM2EpmQ3sLggAdPQ/tpEgy+r4YMEdIRoGuO7WqA+U1byn70ZTgx4PtrOf1W/RhAPrqWt
00MjpreVdsA542TxBeWDQUARAgH9d+xzuTjpSoCtg/H2s7xLU82RusNSq/nizMQAEM3e0E+EkX8t
pNwCrhYxtNuJ/POw2N5i9R7Bg6uodMUpK7ZdR8e9DWVK7KuE1dcl+UYhpXaSz6iPBZvlF6d1HCZf
INs9lk3dsSC1jbMa2r+mK3rQiedpJS5l4OmXQIWHyhTKpYmy6VA0T/wGrndiKQPBlrUeU0uf3ZVU
AVdOeYyV8wEbSFyCvXDKeLUTrlzSznFgA9i6FGC4mUH++dcf3HcUIYzaPqE2oVbCvNNGDgiquu8E
ryrVaD/f8MJT7aOgIRdL0uWUq8uu03DfWBuEFz8HaPdUujL+zZobtGPnyRVwoUOSrybYCjx6OM7a
/x0qqjugjQWtXVbEigRBgcIQXkKY+pPtLqkRUL+QjbLU0c8caIsJOu1kqMg4mnI3kyNaz8zb+QFB
y9LXq/xZtMsjWiyp1VuI+AgsCjVzhkG6l5Ky23Qo7+Ooft0jNjDebVbLqpXG1n1F8sWqcEN+Vo13
/ionAVOEJRxQirCp757pLpuL9KeJhDdLhf781MGoA1I5NHOkSIWiuOBbLDVBV9l1VIOeaFgFDzwD
qD56c73j/SwVM1AOyfW5h6uUKhBO51ek1ivBuq2p45MDGpHcml+A+zR0feHqUCo/oQ2RDQ9cY9vC
WPLFdxgMqg224B1+a4Z6C3ZaRHPbHq1FBsJy6G4D3d4fqP9F19pDUOeXxJPDjc1qk+KrSIOtZQDu
0yyLsnhrRrCvA0H7DWwcvakMkwmpnTXC8Z6sQmL0xpDYi+xawLbh04OoN8xy3z8jgxUbTeD7haVG
PDUgE9T5/KWqaIXtJOFYXyNw4/wvrneBizk45I4hLfdovkADmD49gOm4adEi9x5VsRLIZaC1V8sz
JrSRpa60pnlsn/dHX75/HwSURutROZy1k+l/0LtKjEKmSljWIT/D6eMXQoTgLxH7oibt65f+7So0
kEzQuUabngK+TgLl1QkBHblG6H0NaMm51UHBh26YnVfBw2Z++H1IkG99BytnXarjvC0h6/usEp+Q
6QeyfJsZVlEsnAICDxRdpvsRyWrT4j5KVpEHTVRmeqXAUiKoVi72XAwh47xNHTf7FxYE5zIDl2l7
TBTpPVC+BXxxP3EjnOhrFA9UaV9EGWmkLyWx26OWXvUdFpsURZMalhcnBefal7QhPUqhxUQVmToW
FcKaAUUjH66ZjC4vAHO3ulTLFDPJ1Ai/CyGzmCuRvZkmAsGth6DKg3GXpiu3DKtiBpHOO9Zrtnl7
BeUpmt8GrbuSHnX/3sx9XnYcGJF/hh7B/vk3OMnjFuNxTA0We4D/Wy8Z//ARzLF6ZzUOLC1nZQSz
5dXWGHL3Ap4A6gGKDaUV4pHTlD+lCgh4RM/NLNTSrzWCFeFTpQx00O/0YUAF/xUdJtRovF44Apoz
30q/rCGn2PRuRJXyAZnDe3mZ0w2VjEjgfWa/zb6UoChR7qQd3GRyodJciee/7JDAWa5osjqyEIP/
wr1+5uLyxo4Q97Vtj4ATI/ba06yLH8FOPXf6sN75oG51cX8gLvQEdNSa/wW6arGKy9XuGhh6Go5B
4mDdV7O1DO2geQ1SsjNeJNrffRb0qT52OvR96VTuuYoNnpRpefaKXCk4K3ohPDCL8ip8rl/VR5SB
JrUFpSTlupDbfxCWmC2t0TMZ5yFtflimvTwafHU88xh7vKPr7gLatk17VZ2H1VURzZKk78r9qX8v
tHNuXF94doiCAyfT0c1F7J+E3QqYxI2+r5ed6EJLZ/jlQcWrNMzItgdca5m0voE1H9F549VtWKHx
Wq+pMF+z/NbN9jNqoKxrFQilzm891hkqQlC3OOQv2UougPMrRS84j9WqUAFbSQkGfMDSUbz2/0s6
MXyGcB1U+dlX7uuahMNpFVJQC8+89s5+cNal4U0Rnj7o8P/+hJtOOR1xYcx8aFmlz+s+xOx0qDW1
G3zr9PtIfzFMC9PCko9iYLsxPmSOGJOcNiwhPbFF9FIoScEUXBwrk6J7EETdTpDgyk+Bqna8uRvS
q8GSUeJyAOPTrHeYeSLZIDJHZ6SCM2gKAr3HFMs10LhDvA7xS5CalqLgqZICP7pAHzHV1lAQi1Xp
mZ+D5M8qk9stE7lXDyi3IC6aq5LynPIMtwKsAhGOt2zHnGBOCjeraVezMewmsz50Geu0sJLi5lg4
6y6PjHqCrlnC6EZ7umfyG49xA3p5Faq8693KiF1x0g3vbwQJVtWI1L85n4bDD8VhtNLCPGFPQfQu
32m1CD/5kII74tERXsWVL31xZs4AS0tY79yie/e8mcEBqlJsZK+f/25L9qx/BLBk6xRFIvdb+MQl
FImna94aQDzbxQabXiHnnxLr7u6U5PUToUnKv2uro2EOV9kiQRsdEYc1MbogdxJIJY+uD4ISjFW/
AQ6or3bc8Bawa6KNQULdg4PxGhD6k8a6zzT4vBNtIbUvPMQ9h2YBVsCfxiVL3koLS1ASmHc8ELti
fMxmfoyWXTYkDYbw5HV3nd56tHWhPk40dWiWMJxMWBWJ1iSSG9i5sjd5ZItxr4tKvnsHjcagnP0F
G7j5VV2pkd2tsOxZZ0aunCBmRXP+FYRfnvTjCmb5Fad+ZNRuU15nJEC/bTPGMEl4fB09gw314Pgp
nmxOO8iwHCyZSpwZe3by7/2ZOJ2RSNcwpt3mqO+gRSsaHnzjg2sMxsnzxihwO4YL+MJ2vJWjMHrX
Sw5fFTxgjntfnCDzZIZuRnGCDwfyTNzY1lpfhgGyfykDESd9bVxOP2r8LXlBI6BQkK/8rPi7/o41
0UXJUzXpUeCEoGm8FK2zwt6nDqQoxz1dZO3SWx/7p3yYCbAFM0WrIPBxahg3grgRz7YN3TgGDEk7
qQ0NNZ5IxfFHJvIBR+lsL0GQXpONWAjNy3KRnspxYUbWkrVN2YbGss3oMCNKicN4+uyPuzalCB8N
oVM/hgUMfJNZJpwheTwk25msZdezFOVyctmTSQ6UJgux0UvSCP9gExySVng/cS5Z+wHTDUm9verI
QSDLNbSmLit3zjEbzAELNjhmyr7S4qPxX/qcXLzY/eSNy2AZGA8ExtRhpsO2i0Wb35YFSRDUaIrr
V1FU3dHbM2BuIeplX+beD5lzywg7qiVadcLorVyf8/0dNqSLGr/pPlXeSLbmJUYnkaIIDCNCVVNy
A322UbWSTYflqBMbOA3NZ+MlgoKyy2XBBvu45md3fsblRzsEqwgBKIXOmfduqUP3TWYk0J/hpT+8
kedk6YNCcXaX8myIHamGdGwbsTPwfrVSFKHHzYen2EGxNs52mxisFBsx2Mq/iB6dSp46y1GVeuaf
Zu+hNf3NiBEUB3ccl+MtGFANSgDLVOfw8AHLo/m23gAbSPpAD8CNuWf8d3+d0ff5eCvHNBWkD1//
m9aGHdQA4IGOSic4N4A2TJAB4dqo6Js8FYGmmWx3viR6qVVuiFUfBUqP8oH8pRq6MFXJgDq0sk5H
TrsfNdmj4Ds0V/gCu2F/VVWUbiw02ON5PnNCOgNUMcKIpcfS3E6RyyWZwEO56koJCtLYIQSzkKmf
7xUNuGINs2AJUjjUQ6Qms6or109A83SAk6gm9h40wjYwvSxDcLqUi5yNtFKAubt6gUX7XOjykXm8
JY8p8vrQeeSSl6odpiAigy2nJWWix+LW4VaIRtBIPEGUi8ks31VG8TuPb2D1G7lNGiYWXrJ0S8fG
eHJm4YJfKVc4KJtk4XuXNE/13lmutted0ttNeN/9N8QO+tkX+X5xaiSh/trN8nIodWGWbIiiGzeK
4fSQk2v7BOFeq7kvjvCbGj1WRMb5zFw+KFnPfsy5Sce8HTa0ensvadgF4Z3cJPAVTJ0CSA89r8k4
wfQHPW5DcgqweMGVFXYqxtek14zF70R93dQVfAvTL/zHjzShq4RJGIXmLEkWJ016n/i5Im7g4fQu
AjSiPLJBi9HjIqveD2zl40CCOorWrbKLhbCkWIjyjEW3ur5mFcaFlSJ1wbvZ4SD91QHSlyFPZWTz
e2bN9JfIHFq2UnHLpT7nKRxsYSrOW4KKe4O/KVC+ZHoTgYAmimVP5FO5hH7jdo6yXR1MBlsprceh
yt+3XQRf7UVDMy2tO5hNOel90uxSqgTh2gEqozBp6Twyq92RCRnyMH5WKFyqqCTMR3kOU8cycy3I
BRpkAFQPQsPFA/evyWX09K0mEAOK4JirWTiNlLqC6egR+925re1NjFWzoIW17ZGNvzEiCgfUUTkZ
oyN0adsdHEA6IM9yEUK9rpVLt5QlyNK98FgpnMr1zpiUA3SFJUGQE6EB1frtmaznnd/ddHH6u4ru
K6Fqo5kHAvf9dgcQUIVwomNb8Bek7PxQojntlVoltSFEXKkYhBPh2VnkntTSbwXlg/akrJrBhw6S
A7TroyojuiFIAjg9L+JDAvdY3MPQyCYSkWBeGmomZ9Mr+BowgdUTtbaeuEv8S8Gu6wpRF8C5x0He
g8bu+XQsGx9E+9EKDouNYt3Ebze3xHafrO0bgKjnlrIrEeJCZ3QEWxY1Gx7eMnyM1nw8kB2n2vez
FwR/6ESxSoU0jvpDaT7nCIGZIedww7sOzyN0jTsV8Q3Eab8q9pW3FxWcAVxcUffxqTMT5Y2QM8iZ
ge81h646w53hLvqcKZg8mgP32rckwQv9l5LxLwJoBxtM1YBU7/EieBqUlIifaT5lF8WH1oXHm5eP
8/IEphc9vnjh+4WRZFaB2hTDoUtUSky83Mrct1tIDX2lhCnKLIyHV+OF+WqiWtcGeMKqyb4LiT8H
e/RBrXCDdpT2O9Ar8JIRpEAFNfIWY/8Ga24WJVqo+07VscDNBwb9F4ddx0UJlRPh18TRU+98Fz23
aZjQ14fomPifpQ19dFcy9iY+Q5shKJ845Vc7HkbrcRq4VamSoGUHY3NLsHsPGy7M7OCOR/4EO8mm
1Bxh51MCPKqwWpE6b9/e841lBqyhFQmJKJz1SIZLFIer8XrebWC3PlAnYaFRo9L+V7OCFYV1Y8Ys
a3NVPZfbhTEG3wK9nel/1U9a+XWVbg8EwehSvXZsrbqbJQQnYNag/y4Xo4BgfRiVlins5IP4aeAU
DqJdfAP4Ne+0PZyiW3lusvR8qkkhzksPSfX6ZZUYGBLgtW7XF5i+ytQ+TydUUaf4nVlExBXpi/zP
mf/ZbBtbJntKUKhIIsda6oe9BWpFmTLfUzm+Js48AqljNILS+bYLQAxiCzD8XEoK6BIvwA+6lQ28
taM9NTRPClCh/AJ5URbFGR4Q8Idmiqw9ONkaazm4NnlN6Eipsu6JuYHh2HAhjQcDHMqZP3fefitr
mTxIqVvrUTJ8cgzTaelUWcldI96JO5ko+7ugCQfwMrf3PEVHc82dpl7fSo1y8oonuwFZMwwHqTNy
cvCYmQDuz+e54UP2HUq/tS4VE8sFGxkBh6VC4qamCKSdkIjCQeIKoRHxNVfShhnl8LPSsJNwi5D5
G+2v8c208ljVEdA0EEOkCtJMn7KmOvtnk+oGXBPqy9jIOEzh/StVNDEmgu2WwXTElHliWvWTPu93
zSO7i8aF7wuekWHhp5Rg3JyZWetWvdkYNqi2rLBuS75wjRBmzLWKRDU4n4jNCiQk6ksI2yA8XFJX
nb0n4dHX+t6zGNMySQiGjFvtD9YE0gHU0/ysyEYxxOdpY9ttxOjGlbxO8i6vkImJtjV8JW+CvEfX
DtXn6NN6S/JtUEvC+88w6UWLZjhEXXVomJQlckcOn8tCD73SSVwN4R/9L08Hd+rRVWbGuLI64J9s
1+sEdri03eXA++1mDifiqUBOlmT0Isefd29GbyRG7bigEdjQwqd9Iwz5DzK+5rAWfBPcx1reqWvA
rHC1IR5Nya1HkfDv5rYy3Uk5037FFSs2Qip59cbVO+uOUcStpAmacdjsim+WQyIIM/Zy7/iJ1noN
erbs045YhJaoNzcrRkgQSoUsP2QwQRJ+d5/dD9UmKnM0fv2a+UWJO8rNbVVVCQp8e5K7SGXjxOwg
6lgPh5fPHZK6i50MksDv+scB1Jubh5dLjYfjmEJBs1yERCB7P5nf3jQCEu0hYHjpTvZXZhL+TrqX
Pb/6tPCQ/bJ6VE26ODiC6DIkHgdrFfi6j3cW+WMaTVd+5LWYqcXurD9qGe5hiT44wLvws4ohLnLa
ypewSYiSywG/Qa30Pvk2NXOhMaAeeWmcw0hkj1lKBanFA6k7s+1bLpTVPPYSTRSaNm8Akj9iWgv1
QmjQJvFmMAUx7px1GCtIzFnw8U+inUCE4VXA4veXsMOlxuEZBlOjBxooIWWUi4U+/xD/XOAtq96u
uZJtZ2PClD/NoTAQ9/QZu+l92GmWo+oxGnDPM2r/NV5ni9NxnU5jdSRtzCukdTKkbEvD21x1SPGa
vuFgVIymCNne0cUyATa/oeetXMJI7OrX69fhRlsFV+NPuNDcDurKYfm6ToYpo282ua1f9Zryo4Q6
jfxlC8YVQ1+Vz5136Co4Wt2tXzBuNZxsRogsHIxvVo0fgmpjaU4jjosIH3QBh07S5XZxKaZtPuzT
Mnh8DjG9MCVAhQB69WdJyAz6sjGja3bY4et6oCziJtMlavLf5CieviFL/U4eZfZrjpWqVftquOMF
GMm2rQyZ1q09U1eKcNtYjSQg1g6Q3At6wV7jB02jcC1Q9ba/pTmE/SmgVtsxmSzMGOrfRj2+np9N
gVSqLZFqVjo/vM0IwEdQ/9V8GWka/UErDVzle29aiO/mk+qhml5Z9eMEdF2u9tcuMPEOMU3/IIis
g1anZ7QLV+WcLtuQe02S93pQI2+5EexUwx+80Gszok26oe9dhSd5aFteMla/rkFvhFKi95flY9wM
T4tnGZsaHMloGaMPtP7AjzSbcAc3fvl0aXW7Lp9FYOgVfBY0YyUZWws9JNEB7QACDiBntQLFoDQy
AYyRhSTjOvkrkWbqK8UY3aw9lQzJVt0XUDdFSANSTXA3zJfF2caiVYBJ49XzU4OS5Th1kwPZeZ7U
x7oonTp/y3tFkcyNtHGa8/dsV6QYiUKT49eWp4dGyJAXnCjamitQpQrQfyyNfrm+Y8+9OSy6KbVl
+5F1DtjxlPD1SJK/lPXgnknqy/Cv9N8wP1WgzBcZ3sYe0pStX4PUchoiW3m+L586LXxy9lePm5Nq
m3+Wvq8QxC0w/G8kdEGl/FGVhGft1WDTxVpdbtA3SycobPCxVNjzr28iSIMpKjQZlbRStHxeNhc/
TtA/cQtfwPaPF4YNDZQO9kZfKu1x5MHtTfcnw46VXLVJS6WIgab5vCNbUnRvv8yqtvXCIUaW68KE
JvSqGvQ9IIAiHUYDG3c9PR4yO9ETUFjZRIqK5r9pFg/LQlH9DP9ZyXk+d6AJCzGRkUPFnmAZibQH
oJKTgHV4IuzCF1O2R2n6qW21T8yiMjjxoDd/Sy56EGTs310WSFByGpCbAqGMbqePWuHxJctvhcdw
3D5UTRd2QBhIwQS/XWoRCUxV/g4XKaYXs3E1jEAdbYOBF3Lb7d/YjCfrIP15PvpAuZ2UZZCe3g5a
uUSmkC7+vx42N49mmfCQxND2jlwmzZ3CwNRf5XSu5mdAeobmDW77232/mIHa1tPG48ecYq76w53s
sE2qB9Tni5pAvRzDn2UKdwbnZ91bp+ePqEXT3Cz3AjTLddt5paUTPfxYryCsOh414GKuNnL8GEHS
ku3MY8gIc+JROHoTwRoxAg/hsUkWAUWrxOTyoHG5Q2WbOpYJ6hLxcNzsHSPD26Z41P5VwGcNFakU
3qWILPmJ13ISE9KylDwufqjg9vEU8LOeci8bhrltgbjhhH4iUUFXN25cpVSiVBLJa4+xBj1Y6QpU
nLKlDb+z3rO3nHK/08NhjqiUSiadDVMSC4hIJo3BOc6hN2wYAhciju8wCS75G3M3UuHRTl8Ub8G9
F9/qV2Rho9e1QFFc9m8nRnKA2Q0dgCUqCs+G5uuWUl8fWx6DhaNDD/pAaMxEmdYRQvcNeQgonppd
sCRfFH4uhFKz/bpQylYsVrU6NNaKjGHtrJU+NldFzumzPtkxmOcrc83sNRl7PjGUHys7E7zPp2b6
CDo6TMMsvJyjjkWuG64CHxjumC74DCRXtuf/n+Fv5uvK48oNf+pbgyXnowwqovtCc8j3luHBgJOA
FnwrjbH92lbbkY8fNICJxB7cuAqf6bGeLolFkS2OgqgMZNhgwpYqRLvsN0VhLg0GADtLGcroOSXe
Chnb5mvDUADVXOc/OWSU8WlDNB6mAVyebeSpjyHPF1fjtUZ9hEbEWMNcEMlJM0BiYf+2AysySZtx
taOD4MYfHvBqhcxDqeeX7Bib/MWwIFVsTyvgE9IkRhBcjU9ItNIAQbLGLkDamjwpAWdG9qwWjg3B
GYIZA0rCUx4thZXRSWjuPOMU+CUt4k9I43UYLukpxZvrbRTOEKkSy41X9iX6SnI3g34PLAqjqZSk
6zUHnj1BP/pJux2YMolcdae7FVv7rmF+eQgAG9l110q0WbkI/rEZ7vxqoa1dzRvfFCg6w/YMoYk/
csVYpnVVbqI24wd4O4nMAe4JcXvK6YmHV0MZ1Db4v032WQWTggn65qNqETTLRRi+Qe0ooZp6B/2N
pu4eg/lSii+bpkxy8ll9uKd164dwB5UdvPw+rGXWR0OJU3qoe2vujYJ7QbCOv25gmrNRxn2SFArx
DMWd/AiBseK7R5Cz08IkwX4a3qOHoJN3rck469C/Urp1PaEZsqgsRdZ4LMgvN1Jl3xanMrfoovrA
iCyKGBBXaTdRzGRM2jkk8vsws9qUQjFi0TKiepieQck4CS7zilG/UxGA8Tu3oMpct6m4w8cbYg/B
EwjyIFsv7GGr3YZUDg4OKDK1I899bf9JCGXKwytoFveaUlELbTfAGZyJi2oq/oMR8rQItFQ7F+eu
3Y93FCzlln4ZWDccBW6M0ovaSaJtxgO9hcP+4XSDNvCSvXX4nAPUEphwFg3709oD41d1jt8kgYsq
gXB+BsXs4Dr4FcKJkAtO+yEpAWwfXWnVNAJ6dMOMm4o7wjxcwzYVkEIin7t2NLVkKX1b45zuk57/
dMIS7NfcR9/7E3meDdrXniSjQuY6RsywOXBpwIXJxCARt3nLghPg7uncF9i++HPpRxeUWgOEuc0M
R/xleasGj5gcbjjYX4dKcHBAyFuSSp9q058kiG5g2TDBiD1RwWFFRIebpSZPrhFcVR7Vy5A8YX8f
LFBJ1ZVOe3v9uahuBYany9Xfd5pCZHmkjoAMmktKIjVx5lGsb2xSkqIYfC0Z4AJQ6tGGuwRe6Y/g
o2PWMOwdNhC6kLtJHWd2IeHJewWVAoF7qssfyMCb4xW8arQfM3NXhQcCwoOq08/VaPtPDmpkwP60
kx8lSd30wMqDYkk1kDZMEBOR/vdq2ynmkEiNWT7ySUZBALB/J6pfFP0zc87fc2k/XbpF5+XnGMk0
39lJd+xIMMb1Vhcoh3eWkMA4eQMWs7rTGx3jpD+1rFC3Dc7wmNRqkmIMrHoh9et7PZvG3IcHDsGs
ycU2a3y1mvcrBlfIBQA6kyzP4IaegulfWGqiZdTIvTel+cF6GvT77i5G39DdLIknA+CcNPYXJ4Od
W/pHjAWW68tswoc/Y5YP6hgcLF10Ta694F2MPBKRDOw9WYMsUlUQbI6nWNmaE+kytXmUPhf/kUXy
4bQdXwuU7oJiii5n3eNYTnNaBO2uilkA4FBo7wzXIZrWYSjEfPIvoy+nKfxSSYFPQHdfVbfkLylt
gdLlpy/MUcse9z5SUrc67H1COSDKJNt0INXEd7NTTZrtPWN0lfYBHGBujWSQX4l3h2t0tEKDb8lK
Qe+T3E5ppA47BZor6x2JXdqti7MbFnZQga/aYmL3zumHnASqJQ6460k5COu7xbF8q5UgnzZO82kz
a+Dd77CXlU7w57tT+HF5NTrv1ibs3jl31gLm5m8unagi0sR+bbcr8lYcLfk5zDuZwefs9KGCu7DF
oLE1Nt0iVErUenQj5fzQJ9JSaT5Wk0zPKIjj8gpQKkXdaUrfwKjAWbkUl0i6zXUi1foJzFKg2sJK
zedNPUh8+1TMVKeeIVwvtxQRCIcTqlJ3f9wYMLtCVSvz+szyMUZMFyhpxdvgWqhn0VNFJgIZreqC
YtYlxfuoTWRoThL1MIEMwpOurO0+/MAVOQ9eQeAS2wot0mZGdAHyikcFmi48kL87XGHof4pEI9RR
5+C0N3wmy77HiMO3XSVPEyPOpiq650dmNNkxwy+CRPwv66ClEYO8dACYkAN79+PG7GEDHm7Lhw/5
B57oV3tFEvbs0SoWu6nkLa5jeA4khTa6/2PY03KhaxhbJVm9+2ByU32QbdgrkAf3jOwtzP0NEsGW
+q1OyYwkSs6TdVF4I35SAGKMgAeRm7+DVOetcY1cNEyM5KNY2VKXdTL77yZfVgEz2Ab29aFURZxf
VUf18rdOCddKnusCsyjr2N06ed5BFcbeE0ykUTok6C0ozblAHPqxLzFJu62wN6SxCYnZ03N+Nclp
D7qKU1K6/Qd+ux6Er9odEXX5F98PxrsCxRuWcfFKzgBEa6PXDuJsLDv8ZuKtm57qVRQAZh9+Sl2w
CUbPQPxeMfqueGMIE5CnAGwDh8sEz+/PLzcb/BLSvyShUw3NNTW0mbBAZubmMud8mIn6OBSB9Oz5
C6mPfq4KHr59Pf2xtTZYTsF2Xjr2TDzFR8xNHZzsBJgy+DlWHSujah/SqHwZSjl3+3URF37rPSyB
j7qteBhT1VA1A840d7WIEuSK2gWbcrJeRleVOz6EzecHXlGhb9+bpaXJ9SgGkB8zdHskTIxu7Epx
45jmG0TLOot2/kdwIil3AnfRLvAaaefoLFaVQzKgyut83ufqbMtfTxSfLWRHFXbDXR3y0qNEIobV
slAb2JwRKR1J3jY7ZoM9TIV9naVxm8wC8Ksasg0STCyElwSa1QGaeFfPnZx+X96QzG+ywJ/z4FPl
L2kTfkdbEOnldEx/h5XdEzhqQes/DTPRGVw5gQZYSnefEHhgfeHnkyDxwuyvy6U6NadHC0/jUkjN
i+gDUDOz0oe0dTErBphbXep4MuDWFibRYVOsqTzxjb3+zdt8Vh5/jcq49sT3tjYQID2y8UWf8Wfz
9RSOFzJDsvlAZQAQLAYA6e8Z866avEmVdah7UBmhvx8UbYujjP+fmbelo9yoKA8XILuQmwm0XdLl
zLiK4QbvsUhqNHq+bIPl0HWBnmU71cHJMxYpggRNzfW7wUuvL8+nHLpU9h3oSlD2MsTjathnKeBl
RnnTArE8ai761S8dcvt9eyGgr15QXo0lGquuXchbeEzQqrt6/XlzR5wgi3UKiCcX6w4JVTqZAdrP
dT6i3Ze83SZ28L5bFYuQWdrpH1v8yBTQijzXqjTNf2PW6qRvLrmJ0HaCNM5/JEIDH/aE/xsCjrIh
CrKBKtmWairAgjr10vMWZXYAhLT1RWZ56qpj0EJTLZR6M1LOenGGurwe//Jr8aaK0MK0i/KU4h6k
5xfOvxwVZa64y8P0mzNeAsIvUBbUMNTtkVsa5serRCoFVY2uCgefRr32FRAyhRSjrN332FdweUo+
erfu/5Iy1fu/DPdXiWwjfZCdYaf1hW3Sa1vQRO+4daqnQcydv63lNtpJHzv0KE6lf+LRyIdzMn9q
hJ9Nr9StSovR5EGq3bjzw2Smo9HVcZlWaBWc1QLH+4IqPRmzfZGR9BylMj0myXkIu5zcrKS3no/c
dmEA28kIG3DF9SsuWQ+wSzhAnOLQmhlAuloTghK4d+JXp7AeKRjw+R2++MhP4GTUW2t4/k4Tot8m
23pasmRYPscgiJFIvLlKf2PNcQkgLTNdEt7/ZfUcYDsMykbJAU9F87vZwaEMLqCmOJWCtgT/StIb
ofc7LjCuG4ygU7zp3Ew4pi8mWNDauV1j/BJLIXEbTuMPODf8om8lJ0kXVcjy8OWQpZk+glqcBhxu
tajfKZ7i6qfFXTOnrvr+/DVL+x79j/uWTlRq3vwQYj4+mOgh22eU+mz8ArE6wJm0Cwrzlcx6PU5S
1vBK2aNOTSLjJU8RqMTAEBkd110dnbYkW76jaywd4QmkpdIOCtVRt1oKW7jtzh4n6HGesUHF1LxA
J50I1bsniMGED7uhw2PN9l6iOeMz7egYOrCioKPSsEAlgTwXdDOz1G/UuAF44sRRDqCcJeT5N0bT
+4CFuXQcOQLho355Hz8AGjjjARy9DPvQB5GKINZF59EP+zfvukmkdTzXzDJZSJxABZ/RNMzvQ7oM
49txUv30hisn9dMvfkXDglX1XTdkUSFiaXEQOj6JiyiGw6m+VT2SZ++KZyjaZzBTomEDGL7J50y2
wq2AzulX1kRovZYgWoKIKnGc9q6ogqVogJKxr3W+Ac1iWXfopDjW7dlxFIayhO+CaRrx0+9iKTFm
8QtHM09+7TSyzGBmqUWfxznzY/h+hYncVbh50yR249YHraLQpEh+IMev6naYbm35Z33IJL2fEEn/
3PvrdAcZXbhe3cBynuR29a+m9DZODc0rbT5tnzFvFgwVeSu9Jy8KbdlJlXHAHbcXrmYoxx5rBnLs
THWRbnGnPd2PyAo1DJNeq9IgPaFGMGShGMieyw/aYNmPuMyCj2vOFK9568IkROpmmKfOufUcrV4c
vQoUxNg4V+6j2hvoT3q8pDYJbENaX9JX3m71n3HsxWyy+nx7bL0r+ivhUvhtIpUVOaxuwr8TL3xi
qB2wZBzoW8tDz+c9HtFV0pZmbqtf7RTi01q2k+E7qx4eywlbsILR8A3ndvxPVjeZHNgXU5kaoyhF
RrUfaZMXnb4zcgZYPbd5ZAqDOqcCDjrKtEGM2RO89B/Mn4JY+FW7U3Nwfkw92FrDR58QE4lvyEkj
x88vXyIfAK166yZeW18i4xWjc/N1SQ1+P7FnAw/NC0GFtxWOUcWaNqgzjr/zPtRm/0/LzRmh+roo
Sy/Mw2VN/BaqqE0tAztcmmRI7YPgOuQ6zG0jdnJCkpLxUqtDVEj++PsB8sldDvAAPABnqzH3Xog7
PKdtAIu70WoSjnQWG3viGyjQvU3ystqUlceQC1V9EtURz60auqK6Sw+Ju0A1e+pRn+4lwt/ICY2n
TWoHyYr3TLazX0k3pudGsGr3hSpfqsO/K49cZD0LZSuF/PGaWNBymvnDrNneZh1EqqcgsKH1Zrmh
Y2lqAwa9FTKW1U+J9PM71eysjCmwk+BHP0GDnwHDARUpwgA6LeGfnRI0dqeDvrvahTSZkqoI529U
1E8ZG6Szy0jyMX05zjc1k3JHX541T4+92nvhGPmbfiPQZZJzU7OWwPISlukWbGJYVqT84zEz5GW6
ZwN/U3Vt+S5HwTZMLfq+uDBsVCHTSTF4cwt9yzziOS+tQcrvQjFuvz44h9AO3k89CKlcj+1CeV1D
3j5PKB1p6djsz5vZxS5LkaXVttGywUKZ9s47dk4dkyHmmCdCax3EyPWUc/MBN780dk4IvQcZbXbU
QkYlhKHvMo8vkBW0YoyTz2bBhI93TY07FGrNv09ZzLDuj2o3b/2c95LQ9TJgcG7jDxOUBwN9RG+L
ayTQQla77e2PX8E4+6w1wEVzptbtcXTr739xQPe1oUOQN5lcoHTL8T4x/ugdmNW/C+NCDQpSFbiB
kc4VQSyUBmWe+N6CooraPBcaWB+sW2Mao6R+dj370XqzTgthcTArQfb81KQofaR0U3kk7Tsjhhv7
GhKOZd1F4cTqrnA1nLaQ6L+363VopRsznFqvvbDYG2dllDK2a9PXBnkIJ+50VXLMadq+I8KW78/Q
s7Pc6xZP9XYCHerx0lImr0yXJfR1K/XBfSgkiZZ0zLDykiLLkdcVUBvuBLIzYCT4M7qahwINU32K
t+YZ0Gzac4p6sba4vBJJyzZCLftpa47dLHIGxi49eVIVoSGF/05+24r9WSZgatXJ2hcnPPWy+9Tv
XaRcts6xd2KQbSZV+fPbxaJ/bhX+Qt+WAWxt1EjdX/OyzehSyqfM7FUFfvL23KZLf70XEsN1370B
Iugs/EXgYMVnXidFDJW/xtTn7aHFOtDDT3iwiUomkFnofrYu0xXqSPPtD/4TgQOTmBqam2mA/q5P
ZpQxT8I7swTokaBMJU+27tbsyzN6dLJJf7hOyQGCI/GOJpN0Ns+jz9oQnrKZCwOlW0oTFwLXWyep
ydcma5wwwpok2fbW2ULyXSsIEKONAmpo9Jh27+RtJIf/cyEmkaZLzzUmcXsn5+AQOqaFnOG9YI3y
XexZR3c7ayosHe5MkgIc9WnTRxtKHnHDv9zwHWyT1GZnyr+a5d2w6mA1bC2zWhsZ8VRBgzg8u55q
cN/E/t4tB3kge7nfiC5nMFaB5CUwseBaFSQH5F5SXZjBS/IzLgv7qZEiTM6pPkrO4GuohLdkP/fH
zM/zXYDpyDKGNM5EzgSPg7uj7tszF+I57nV4wl8fHFRO1G+6Bxfm1AEjLNUN9gow/TfEJYja8AX6
Rqa35o01NY5x2qo50ZepewIVEPzWdn1H/yc9hK9+A0XrywrRT6wHvdtHPNeMwvhJpZp5T/5TT6hs
00lYpJaio2Q3XDOZj8jM9BJHLcyfcDkYD6RHqovPNjhOaB8EO+2ztmt87crodPdE8tgh+SVXVH80
sVpvGmLd7v97flScqQvOJHmVLPfFAJVnFPcBx2yn1lTgSHewDIQKHs15Kjr+bUuGf/PwPbbW4/na
u9R4RatkN13Iv9+QsXkBPT7YxrRllrBIbRKsqbLLcWLbxOxHryrk7PuEkzwpfQ+jNZ0OOMZFNbIO
LKqg2DKU72s4+mgUuU5OCvqx2wjQRwcgDsTEKqJjpygsdbTjFXcbfM1U6jKoMFvihEualwl0wO5t
cLC4CRrCSCZEXpN7xqtTKzC2lXULnaXV3RKZ/Z0PNcIDx5woddtIzG5qr2RzxHh1bd6/yZ8ZSSIt
FxCgwJ0y8GNKbE1CbG6dkW6IRXCrHRGGGQYkU+wF+r4JeJyo45ST+/n58owPDTpyr6wdLYTfsncm
auaHT1/4R5tzs7u4DSP0a+XL8E+RqklPJGkvdoGKtBo+Mro7JzewQWsiNciq3gCbBdxgpQRsGsxp
TgR/xIXI2e5nB39ZKOfiL2QX9IIEjK9hKjF+/A+mW1gzHDQ9cKYFV4ZiXwvMbYZS8Uf0fhAdjcgi
+gjRueLqnz4uMlxc2YEWfP8qZwoH9HdXOhzeG7Bt3h2qvuoLoBz6hkKL02mVkgVc+5Hk/6y5TISj
T9LIlGRVgfmnM6VqdhWP20fIV3f+wwIPTz0+4V4zwGx+A+dPd4Xhno2ZNN0bdNAEDPbtHpmUZnb7
ODIxVZJm1AyHVgsoea+ohxqfWAojYHXdwe/RTPUYfxlgzs2qZRjQoxhx7fKV8UpLshHXjW2B2Qq8
6FgvLPtb2B3XcsDnmKXGK5w1er1D0Gfz0yhlet44kSp05zcB8oN4I71DLWvFW9yu6zA5vitA5DlG
mghoTz6xlUrg1nGZAsKMe4fTXx8HhaWdFOV7nUYad1MIJib5Uxd0B3aijuRmWPYJpoIDzt4LnOTx
KIMrynVuvB5xBSzkQ7gFv9r77hDBh7DufHQ+Kh14F7gM9hWo9C4aAgbAOCIWqAevhTO3zRXjuZA5
dpL9DxmqXFw3tXQ3T/VDjAJsj7hQrih2qRpSa42xveXqSWd5bMtiHgGxTfo2/PfLXCptUOAB2FwF
eWIR9wy8QIPXJC68WbOy0HzB6pB80yvb+VFU7ugyf6Y+yJRoohM6wrQCR2+fvQ5NJOlMAR/HL72E
vOYG0CJO4j7mTzZzuIUzQmzM9O3qKjOiXu7zvTNNo1ZDo6Iewl/yIDoSP3DJNqEncmu3go+K6TWJ
HraUeOkVL+ErabqZIRYCpmiPhFufzXXjwzBYGEAMFN3839Dih+MzUV1ddUb0G52EPTEkKrOjiQyd
3dERGkJPm5pDI+bFF0ZsOdQqiGeSfxDVef92e3v+rYO7c9Y6t0PSRhrcroftnTjLcgTzkjmyFu4v
8SagQO9L0jPM9Y94868YrFseKF/Jm0ropXrACU4rabl1iYX7i6snL4tR18fAG3sWb63kNDifiNP9
D3AK1NiTdFGI4W7iunjeJyMns55gEO/g0caxEfJ0ykX8nz8TiC/t+7dUmYXVRsCn8i/7YYdsMQa0
5UJBElnHPTjUPF/tww2YNHw4wNJkn6YGB8a+m/hhlG/SldUXu7tRI4HYSpH36liO+TGmQ6+tHBuz
/ERajYXlsBxretn34AaLw9yhL+ZCAqolfwKhnIWK14v+LKEAfRnxa+bh3Ca/EUnSHedLGodZYdty
GkZq0gnrUkalWfrnbqP+wJtrk+OAMLVQaThhK0jIWTQugQMjufGwvYvq5l9ui7g0chPZOavQwvZC
ZPVSv1foh0gjg4voa7FRugLfW81V1X2EukZkKEPc0n1WSUVq3iPuYDyn1iCsbgQF5xRlpNNaEY07
Wx5ZOjMatnh/KlWws7dMHCvCY9VVJ8CFVai86exlmrfinOoOe7+44wtNta6k4nCbLWa57G8s1MsR
I4mOL5P5nxBu/12fxfhDqRl7IZPYOf/9fZkKuz4Yu4CRsv+EbDH8+tYQ39srqq6NSEx1jBXhzMpZ
1+ARo2j8Ru4bHaAQHTVxVodhSbXuuT3lSjuk8RQ2iU82Z4O/4AS0amqdsyWWXscnQ0pnROC1Zulm
rbUqwzyxJDcdAqGEbagRlWnesHiBRUptsPDkIYFFkqQFXsllFzX95aL43Snb2KBcGnJyVMTErb9u
c5tTh5xvOSC84WEIPWo9Z0NkpcZlcyJyeGGcNKPFH/VO+stwPNxnQ3/EBENnznvHPQ7EoIw63mE1
J0WuOLsUlYy1TBYD8+o1ErVVB+nrBrB1W2MmASEi55QgD3TboTB6IWFJAuUExJaM216EdktqwOyg
N927jwtaymmW2QUvdXuK6QynDio/QvuiTW8wMi/JE8FGACx03MH42vR8WzhUqsiJqYXYGTcw4mA7
QCoDK42KP/OwlNbaSYeyN4hx5VzxmkBH34prlM4qFTrIVpKz19mYAMDjlxOFChCID5l1796EhfxY
2Ki3zomelM1YiVxKkyzmR44kudK440plp/DHW/cmXe3EueFVLBh7/+NbpXoTFLHlZ7Y5bsioGNqZ
HJKHl/rv9V4homwQSlZ/2hEY7KGC8/+sY3LlTO2B51h8dKk7aT+Ci6WSaWHHkzeBUByugB/6Y8BJ
UlsyzPFEf8mNOYmoVOb4Qf/Lk+YvCVSvxnMdGX/3qzHluLtScmAT3nyZq08tFVHkHcGPpuNYfw54
yUFBYvdY3K/RBbbo7EthoTSNirPvTxzUQBfPt0mmlsW0ExQxTX9cy/RL9yHuqVGBChY852Q+JkkB
HcDO2XfjXyhBGNEBzIVakjHQrLJilamlA5/IDcBbxGPq1GpWwhhCl3SFyUYZ9mwzb4hMfREat1Ij
j1Cn6iPYeKO1GZjqh2V+wE+qJjaSj5XpHHHiB7eJqXXz2bPh2eVlomwl7pn2wPAtzPpdPOZh3P+x
hicxHgyE1PNQBwRxkQygNfWmhrFkzEVixWLlVZGKLF/aD2+0I9LpHYpP/wTTtSd+C2I0hkQViJAj
qnI8IJpfrZ3vcO1npnrFLJyIEg7yKwL+joKxNsy2T/fMUrwmt27j4d3Ya95FdzCX3xrL4YrUYyos
hf+gu04uLthFEwySCwZ2yPt5c1zZIH8at9L2+3pXT0u+A7Vxd4BvJO4QDUH/iZzwSdugphTHJEaC
vGH7HE8JmLcXIrMMm2PHbTUvsqdWhNA+ADBO/+K4JgOtT7FpAWzyVYrIW2/t1aeoQtdjjgg7BL/F
KG/U4cLLapIN+W7dB3+pn+FGcFxKBSLM6hKN++JPgz412wMtr+SQWowbiQX+ILy2EBaZzDLrj/Ji
jtkVsmoTRdgfEcdh6YUj5neN9zxNu+7amOABbi5vM5Sc+tmvxslPXWN9EnZ6NOYnWxgL46oTI98T
f9LDnKLOgN80kIQTRtWqxUm5XbA+qS5d2M4sm38rLvEbJBYS2yufeivEWv18mOs2UCRli63eBYDW
PCKjds7ldmIPA5ahAlroyu1ExwN53VuFpovlP5LBF6oN/QxjWLIzVUnNiJqrXAv5smAjlZVg9u/z
t5aKT02lrrO/zSa4gSgKj6/d758melIcdx9HZfUwTg99xzcHAubB9DXpgBVcuwM4S6nAy9maaQqn
FC84MaI8uwpu6A4GH3xfLRIPpvxe4laiM5Cw+Y3RMlJNtuRXgBYXk7bXFB0gLN9lmSG+bwISabVv
gt9e6kIQkkAKjDjTEAlCW5BRq5MFZ1PZXfthTjTKU6JfvU6Ao11w8J5XJG9uSYmRPwGXe5b+Jsnb
U57y2M7ieRmeB70PyDp4Ut8uDgDuEsRfCyqWKLCzzZSDTY5HMhlo9tYKxRIKamlWGTKGbq5RY6ni
6imAmSJuHSSZtsG4XW++BjpdP0fNAX8PIxyd4tVmqIRN+dLVW1oUt33kVExpAJqYABkmFJsLUQiI
whmyi/t4c2xsapcSdi0ftWgriET0ndJa9IcGKDDxkPUKDolIvv0+a/WsBfUmBXvi2bxuCE4vbwH1
bpwswl02GgeT369BiuEknHn1vE9HWyla8JvLwI4RUDRYoh3Z4+cXwFRLoTguPwcOBzTJ38xI7Q7T
5uBnlhsIIAETaR9CckpVDzV4SLg5a9cT1QKICLFRuFbgW8jjyfb0bIlU3EDekuh7psrwPWAUtF8X
3gMo1YboSvJPUvUnU592eq1/PXAhQgxnXpSqYtqEKlClf/vWVGorZ9tNUhW0vyg4QU6LeVct1WmQ
oWbGgWjaR9oNVXcsPmkKXhmb1wc9+CVgXOCqqtGc5mdh9Xm/JI0c6ucmMXoMMCbKgDd/suoDOYWo
vAvXKCjDf6dQQQh+MD2hW0P4m3QfG2dp1wnOpxkDvfvlIhePbAHXge7RVBsGDlAcCd1APsvg2UnN
M0970rt0csu0aJryP58f0lK/LXaBsb7VcTXEQVXhK9rshGEso+RlGvn6ennA6sxlKdEeHsCH4/wH
cwWjuA8XefvucBsILssH9mDGL3YBMZsz5z70SScf9wMS6mn0AmwkBewDe8z0LuBMON6mlxLO1JUR
b58VsLwjledi+wZk9CuTDMJS31+ei3eqz3xYVOyrrrI29li8Pjwp8yhNXpwPpgs/i6LPT3SrwU6z
TMB9aRGBsBMi+4RX021qCyWceve94VT6jKXzIYapjH7SJbq/TRPx7ABUemZi9lfBPipO6PYRM7hk
ZLyhGFiT91CI3YHCg9xGlqUvvZ1ACPdzZuQMqMa7Q3x0850SOWLFYwa4xvJGu2/+lp2nDNdbb6JY
OZ3FGHO3kFMsNsYWqFwHXAIqsSETTsNQK1Qcy36fYngOLLQHO/Fv/AlD9SYMRvIEDMuxt736M0h9
DgiAsCxg1YjX/ITEUU1DKWki0QHKsHGlkQf3dkxZQVxXJcVSCnEqNKMkkXoQll2iPMQbql9DfT78
dB+xNLLW2+1XzMsLFz74Gtn6+tYcnBhA61aAEPo5DKSNtsEYolZrhfrmrxtN804++u0hVEuvZYmk
vTdLuqV3wPPKVlJpX/uPPRfZPbW4u3jCOO1naNx8P4OjQyvrQCaKg9NZWq15CLjqnqc25oorbo8b
BPe+TFG/TGZBHuI9bQGMDr/DTcNsrXLlfwTHZGAFlwpQuyhnUlfQo97YDNg+YLdYOTmKkhePNbjY
BHxhF6JlvTG7WBe54CDkYEOv9McSJfOecs32CmgtaLjImzLdHdGZ/AK35+WwXAtASAHMi+lixUAV
d0BkHpLEQMSnhc7Z5g9CoeHjXbgEsGalo3R6VVqJFQRbzo1rgIROZZfv5OipHH9tzfpvMmqyE/Ot
OvP362SMandsDMxPdyKXpFtO1XOg4J8Vctqr0KhBsFSLLoxb1fDY7x12f47dwjKfRhecNYkXK+Xh
lcrkZjOzcwjIEsLaQdCsjTVVk7+m2wBUUzvitkFHoiXPcFEYsfft/ncMcj7NeUfr7QKAUEniS4/d
ui3A49KnkQGRwTqG4N7BPVnaCg6/ue1rIhj1K4Hq18yQ5y7Fv7ypUt9nT3JAvVxy7AZEOVnco7Mm
EhHQR1lb4LgWG+SHw+5jDSVT24nhHZus0UNk3umPWKzUrSZ4Y8mtz9Q9fI23XDH/9MpxE8hlej0e
vPWpZFzEH/I9qnwrvg0VsU2MPZY91/1PehBbi1nPkcqrg+AZB3W8RHfd2xGGigaUPpctRYDNfiha
Y4i37M5DvWjjMPmqP5kT08gjAs/fRgt5jh7hSRlLjWvFSVEaf2R5zIA6agLZQyAnOh1L0/RJbHEc
0sXrFZzufjWhlhSNQkmGtPzbEMFGVSRQbmDjHxNDf20IBKKJlDbCbY35mbqxEYIx/KpGLwPHzJYb
JWFSDmTSe8bjOv7iyEr+lY83RiD6oGa4DmvXbxGIQJ/UvjWiaQ1VFC2ZuY9msolBTHFjVUazOEFx
z9Q1OdixHwZXYElrtnXPxtFGmLnu6w/IaoqOoc7t4w6Ies8j+vFHefm9KvHmZYfL0L98fSSa9ajc
FZ4Yt5gFVXqqf12bXcZFdapvnvg+wCeHRSeHHdFp67RDiZKT60VRu/zdH8GJiKhNWgxr7/IFmziY
aAn8I87mi5RN61wbb3qGXKn74fjoxavWpACxli55yPPVJIyxlmpqvy7O60bDPARL4o4iqTOjvdOZ
/m/gPnzmr3Vg/uMOKCHSxpQLH9+S9bYTISFYIaNgkXgOPXOPEPQJUcP+LWHHn0ehhYbN1i86DD0E
4/BrGXLzchIWrqgVebjYBgbeMPxdDQXVYJeJcApUw4pBvz4TP1GUWRCdInHbVp5txT0jBOUKd+iz
+No9KwN7BwAmt/VA5I6TVealMc0trGjBZy0vKug6NB0nLbPClOvnfL+VR109R0UoWugXlmWfN26k
ptdRmeymVamlZa3tUHAfXBVJdj9Sdk6ERFqmh1ORGdnNcg3VzaScW1z+siT9jySf0hH9zpVsmYi6
EcE/rG5oSnoPD8xvNd21nLUozrg3wixUVHdsCk4Iv4yCvcXEMgmBGNOYB71IiImAyoaMVV18NvAR
/UhODMwM3Gd8lWp2Ifj2fXzpe2+A96K4E2f97vWWjjKO/B0nQpQYpgnOogEfKpKc5piZPBq0Bv1P
ZYFVe+66JPcaJ3sPqGB4r6bWgRZZTY+lYBvXfyetBbKISIrThIJmaBUvTC63FgA42/+DEm4GDVKY
fUxzQ4gDxJB+bS/+vIwIzDCZ4fUQagmhbZpcdQoPAvheX8T1cZgwn2QLkMyQitmG2RDOOQ1vZQyc
KKYZvQ1sHebxeWDc21L/Tu8pYupL2r4EOar5RrtEJDN3vVmqF5nRJyT3pDaG3/TYxd0rtKTkxhS3
LI4sGAKSqi3pW1BSaaj81p1c2nwzqf97aPTNTjuYOOicGyYWozEL2hx1W6BnSTvxFA+sxpsOL0zB
DxZYYK8EniXH0rHsPRfWqaJF7lsJU5oG+q1mSP9gsCFxZDof6/6jGzsrm/vfqqBUjXa/rLDJZH1k
kpOlmukxAYsZd4oaWUAiwdpQR/OwpCTPgf5P0nCODgf5ZFubc6JVH+4hLy1f5wdiSzYHz0DUKGTD
XQ+t928qZiL2MNE9QPHwijZ9Bw0sLYkIWa6WqhZ3ryVv7F34f1kxbze6ylAU1H7+8TynxxCaqOof
xIwdH2S4QQGHpcAJCBZu7JzDXPbRPwk531c7ob6ZM7BhaxXbsZHiCcxpuyVmo/EW86ym1ZGiNGg8
kcQNG6EBENR4xF7zOeBFMuY8dttfur+MwCRvBiA687bZBMDU6gGKyzx/KXT4w60ZGLJqiiIEU92P
jemNPIJToZkGWBkwvo4Rs73epiX15ioP06vQfWM5QTX+KyvF8kJ7yF6bkajOSHBvCd5M8CbbL2Qz
18bTtE5mT8e5CADoB/Ibqy1VdbtvNpPfeK8CSdOcFSUK3S36uiIjXrdZet84yHyTbzB9NHDgd5to
eytVNHzZO+gv9xXk1hPo1mhMhLQB3VSpZw87y/a+BvcpT0suk5Pg/O53SvAwQzRpUgqJpu7xIcG1
8AxTZ2urKXbfpTePc8AGJKUZmpoYPNtzXg5Lr6rvVplnzjRl8Rsw1HmSH9UcyMy4u5/uUjlcnNiK
6YBRL2BN4X1EjSZqxOCG9f0e44v7/pPAZCpXrO+jZ03a8SuiSDuypdLbIQXmIHzSHDRXRveLzlta
65LnFCqmRTeKvKWDKuWXqcWFlcVy9hDmf6UoejRJ4AFdPVU9gCCybvWauof1VchNsOMGUi1KXx6t
PLPvVVfni+KHtHVULPU+2wEN654fiDABfT6DZrFFMDoAmHhFG0Bly1ZFyRb1oQ+I/KtiV9xtssjH
t6tCToLW0AlzJfRnEVcP/JtHc3DmuAjlM7MWMquywFLeoxWHu8PWoTntgcn3oRqicur1XR9m3+BT
KNTcFCEz9PVk8ZRcmRQedNUqtdoxTqSOr2pcc+2F/KovzzsfDEYgZiRE1ZqYSuj0HkY0Q9DGgiL4
Un1vU+MDdYUsF6+4q90vX8kHERw+eVjVKNyiRLqfX81yZXEpYrIZ8OTMazCdu1JwftJAbbmtxofn
81+L8zjklO8vyOi1C0+qfvsOc45M9k/xTziuLc/DBoau3kYKGUb3h7HeL8HnYckVOeJFHQaMLZwq
DxW35vRgVLz/lW533vawcSedoDDdd+NpHFzQezglGAGvq14hzUwCi/rVKfGRCAJNj4zRGR8IV31S
anK9cbgcPBc8fkKoxDeQaD80v7FmEL21W2PchB0DI8Vm71qhov39yY5/BghCtNUb28b+JXwF/i98
q6AUrZao77ZIxzzxovJiWOEOvvsIv+4cpptxCBlN2dStmlbdelJajJUkBIeCWxeaK+oyZPsMlN57
9gNZwirn0sGDoYC2zIiMgyKc6TwSgy3u2L7wt8/sZrQxU1TfPweA1JaBX/8HDB5ptRmdWogMvBUS
g2IquMS0ZeUo/hqkkX60UJIL2p1uO9r0MHejKX4wc7u4VxvmJ93oPa/tIxYwioZyqlLjruGQcSIY
ZR+ClNW7UZ8Am/3fUG9Sx3lCQfmDOB85e2naHnRmP/mpZzP5M5thdQawGapj6fPVdvz45AWUBOF6
24awYmy6Zy68hCjRFrCCcfdNIEQULdjUNwGFzapOGMQonWhFk8zLTosIXmwHZCIWdpsFX0pLarPu
opHWjYrk2Qusdn3WHf76jRPwJq/t0aYRQaGsF3tdNS5AposVdlquv3//qK1mzcKxl6p83DwJLWMt
UuIAJOXfjiokY102OdqgBgLZbLfL1YJvgCexTv/RIXirG58h60TvsSuSNSPJcCUXB6kaTa83nkwr
rXtAK47mp90b32Fhur7pOcdCXImZGCmW/Rz6j8pTnELHE9jc+Wt0J+bbNjlN0qKmkOKn/jBpTNXO
dJkDiBuSP5eYtsJZaqym19jS9lnVD2DG6T0jl2BTClZipfxN83dDDtohGyFSUzuL1Ngg3Woi4ebf
VJGekfe1ORdocX3c/6lykSN8ht6pSPMlIH9IfMPYm5rV17z2HyfB/PWw5s/OYGNWr56H4A89qDNY
L6Ap8BjQEB01O0s+TFxQD4VRmMjOxzYLSmc5pDmwbGIF/X8uNSaGyjdK34k/1AYSZIyGQpU8hFNI
v8owgXvf30ZrX9/6vnMe/9TPskls81xVLSbluK2J3dgzju27j4hnOBDPY6LcfIl/U00JkEXWu3D/
TvbBahNU9g4NQBcLr12CwG7Swrf5PvfCv+Un6F7HmdpBJt1RYt+xLShkpC5aG16R9nuSRxxt4HzJ
/5QY5mflRIE0ghVE537/EcF02Z3Eb8DFBCqL2C7ooiWUzK7InJasDoxpXLspokNfdVHTtJpQ+roC
UOERr1ll6/nD9iQn4/jpZuCMfCTk9U0twHAffznf5Xdqckf2/6MfcxUFAIvxBXHUyrWcYTawmhIA
4s7pSE3/PmS/viWmLevEtmc8s4pnajoPPNM+9sc19C9QtxpsCMEv3t7WBY9NwWn4FG8QSv+pHs7E
D2P1Tkqt8E3fxRF2JtHSbIq228cZEyy9p5HO50x13MhzszrzXhjft0RWloSl7cSkw5NoPtMe5Yo4
nxCpuyzBz1rI7kSCyt2qehqrpAneMbd+cH1bQKFzkFVpBa2AU3lzvi1bsW97o/GpyvwM69tuY7uW
WZZumF4GtERAYRfiKLTbWl8xtva5OV1mqgqsKJc8npIOLuxplO2axR7Ao2dUmpKluMLrQH1QY9s8
eeetgLv4ld77DP7Rt1JCOb8+RueVqQRIO2mdiynAQUR+PkBVWHn0zAzjLnGSkM5w1/cG0uvwwhJX
OkNSNB8XE8oQw8y/IjutRRY+TB78oqa/EkQOIEMiJ0v0LEyvhZmQE4MixGRVPfNCH/uQbMyndRPr
3AFPfUNbNHyNjdR+jykjAOgdnyT5QFdBpAvGo+pZu+b/EKQtbgt47zJxwAi47Ewqq31muodoIv4J
QuR8cgRRy6w0xqJFky51yyvIum9TtrDvB0uFSncUWID9xjFd/u8jOKiGsilqn5VlekoxQ3mg6f3L
Ukb9LPTPsdE3r9fZDxXFAFQB09Q/BDfGOBKyAL7arIbuGBN39WRmP+X4N8jKHu0Ajhxg9WwtSKiz
zofoDzIyLioK1kVnPhW9yztUGViwQ+LgUvHa8nsSiGoazpDXIskYNCyz6J9kZESRn3G3AYRpLz6L
+NWVWf0/YKaSoDrApd1FkTDx7+4/w/5x7NT619LAU8BqvrCSAqVlCqkv5LdifXjbUehA+m+z0ygY
82i65SrH332TwIKqmNZkvqZhbSTKY6DJpq65AN5mNNFgeIcSKVNkEhI/GWl3b+I0uuHPFTWDKLrx
zvjRgldDCzE8RSsXonNX1clrrxjNAXrqIvKfLKjPzMY3t2g0XZuuZnj7Zx6Qhx9wSaU4xzpGU+0D
2Ah4MavJMYVignU8xwRhL49br0nEqS6+O2e2Xt+T0QDHXWZYVDomWGRMnY4UXWtOafhh4CkTj5Dp
LN9XNuOYHa7+p3uHJ009+aiGy5s/cPtkNx0pwtbYEoto6czDTB4t53RbZZSYBZclt/fBhuYdaGJL
ipJW9MXhCS0BwxcZ+zXIivFiZfKjhz1LbeyIjdcOiQUaCzpDsTyg0Y+LSgyqoEgFvK/KlMtSo5EQ
v7IjJND69XaSSZdoMv6e+LanDyHtDt9lN1r81TxmJ2lx1HVj1aoV3j4KDzz1+G0Lmk2DiFF7nhKW
roUjxI9Cd8DVlTeeOU/D9feGjmrEO9YxZLetkiPk8uqRlWabi1qfVrPMDY/Vd2AlpB45G1ah+avm
yvdNQBrQDxZcjuXE7gEFYzN+Fx0sLtn9PfaGIC0PDBYn4V2V2iHFOLB78+BqluUDPmp1bdn9z7WU
sw9sVPSjH2EphvjI4OOWuIudyUogNDv5Aj1fk6nk8rdlHofKTiBeNpmLTtzV6XxVjI6/bnNK8I7Z
fRcHLzHlmYCvzBPdgXd8D5qDINY6BOpZt3gx3VpaFj1hgHqejIz9cND+XRyntrwJOgQ5oDnCzn0r
+fVAdGQpiOYSR63FVvo+T8FWqyiVoscAMZa+4OHBxPUYHml3pfu1/+Hgeg9MEviK6OdvZU5/B2qs
sQKNBjrkGfSMo2K2lKF5uI872itWDVcq5sjcqnox3B43DWRRL07YLIrilAUT2OE6nXQ/e7Fuxzn9
6bAUfD2ox+ysh5Sh7CwCFRcgHkovnirzc6YCt7ipSzc8pBs3ya+4CqRn/hk1T7A5pn4swGe7p/SO
ViAU28pa0ds9MCTs/pXAhm2vKrErYmYqZY81AyQ7xoAftKWSAk8ywc6Hus751A9h9FHxNn/+e3TS
9WQNVcelNmMaptXD2M0HeOX8YLs7GR1Z9Wd8/U2ynJdZGI4hrXjFDh5HuvW529lt/qbKiEJ52tdH
tfypxqOpLMGkklPzJsRTQwwOeSZo79o8cOqZc7LeB5UiaQ+xqQSj3CkcCmDvTEfmF6G9ReBOoREw
GRscm2W+lTl+aI9Xw8aFGvG9REZoaW31G+ZvY1CfvkRUz7JV1WEXWULmbkFZTY4CGbYgNn2Ac+XL
h2XdZykbWG9+H2wq8KKTWHfJPhAf1qTvZOjme9Uzvt2v/dVA0/g9sx743YZPDolowKoC3IcDamZp
3TWpq9ioWqRpalP3FVHntuqmMZyQ0dRLay79dycp+xAgYeXcd7+7N7P1Xu0Os/QwmfBvhFfDtq7p
EGkqsdRwm7bqmUy0RjvJozs6I6RR018Cn3WyAi8D8KAtCjlgs34t0CkpgkShJF/oy3FohlH8oOrl
SPtWLQIFP0zhC8VRzCGG1qbygXoAJQMQFoylTWaqMOFLSu9VD5Rp94GhBzcHkBJMeo8YIYzuQ0N5
sdYqitDMEsvMVvBeugeTfbFFHtnvlTSNV61AAZGKeNdmHkDTnlXKj+GfUNwLT2mbsnynhHIhEZv2
0FTxbuLi/jFURchfGs5vBo5ZrHP5PTdNz7KN1hZg2vT3tl1ecOId08aK5uus32TdenAzSiuepgOU
bFdaakrRvPxvXLb5E3x0AQ72m0QyvopWG6gPELswsfF3A7LkcCujbQ/cUGXs5PUMbaiY4UseLdca
F0KqeKHNmnpmw8dEvA/h+ve68Ny/SAcpbOgTQm92gGkDje+qLAQCYapfyls7t59oMlHkLkOqZZlh
W3Mj3SUC/hKO1w/dXXTVWSotrio+4DdUaSpKY0mpKad+xCPEN3gIU6hVOkrdQYCCJ92Wwul84to8
VcVQmIrr3mn6w6ykIJJ1gV+rvgJIKBn8e5PCBpLZkuF4I1ztxaJfGLltY3Ut2SQFbNF6pq2RI3P5
6BOasm5hNNsdfPzHc/cWaCvZl6hvrpIVPBPoXwYyV2sMCC7GDj2ybklnyDCzefQ7p7eLgODm8OtT
Mbj0oDBp9OGprFC5x4P1zZ/avuHlj7NtfOTSum4+CM+epoFeDBJnhY/DjRn90XhzdRoYAwRampH1
UNypQMGUPEMhRI1shrVh7QVzlYqNOlX2t3D6OWpRDQKmrqyf4Iqj+DzWcC/nWVjiAtXvUiYAmUII
DTunEefIm+Q+Qr2TITs9kLcW0lIEEo416U/Sn2XKFQiMsoAcNvNT8NDrYRs5gIVAmVMhwBK4IH2m
dS/g+nG1CVtAs1dSVOqIWtvEDID7PkrhKq9QKQJfSNpm+u7DnSjdsAvlfs06WILZOrufE/2TJLjL
RbW6v2KPO8dCNX877CEGN8ITsQuwdbxbfR4awdI96CVzjMU+1wZZzvbuaLn5OyRMdENHvG/wcVRq
SSiqw92/wumE6HefqEi+piksM5e1qPA/1tAbQ7gO9J0D87TIkJ4yYg/XcfvgbpOcP3BBJ73Ehe0/
+eyp/Pip9E3eoVRjlO5mcTludVPDAvb6J5uldyeqfufgLALdhKXPmh27qceGhBdRCGqF5Pd8Z4wx
nFxONoMZxh+DDvU7P/uGLNyeu97gdwx40YYk36nD3QR2Tw+s2nCknWPBJxkLD0X92wqviLpWlW9z
fHwg3z4UzJRznzWIWQoErRgtm/jj5YJfDpWHpQ3/tGMq0CBMJzODM89r6GI/PFGodz9gqJN7kopd
NByQx6q+YszN+5GWCtU07y0PKltqSPmfFZKviyPqA5Uu2WM7r0hORtBCQM/5l5T02g4OzDnF+Akp
hxP7NNmfaReIpqr34/dNk3enfZuYMJP4isHtSey1CxG3xxzgQ8HG+avIlrpOa8tr98yu7dvchAgR
bVEIInuKKXShOITXvgFRPM2VJ1mtA2LwT59MUF7qbIiy2arcSMxuuzTRjpod1+htR/x3PZ2xWduE
Iw51XB3FZrmAGH3SIs38j9Sc+/xxmLf2T+E1/7iGn5guu/FyOsZB2NPVoSDibSD139DKWkRIJfFr
cqrJUP7w4ZaL3SM5pU/Vy2lvsQK8YkixAg5nGdtUYc7BCP2BVoUJFEms1xtI0vDgoRG4B8GFglOF
2XOg1fUT5WlSP80+4E7/XLz5N3YyVGkI8m3PtrqsFYYoIbY0Nua3MMnbAyMtHc4l35HIm5g1tI+W
vgMNfpm2pBpEH/1uLVQv7YKxHm+cVDCjUslqedX3J6wf2aATFo1ACEGGuD0zOyQlAM89//MoBZ3H
FS85nqj5YjE4YRgp/wH5+ZIAqugUWZxraEUlaIoFa7qaihX0U3P0uMZIGXkkTaeTxXXgZ8vmQ70U
Wf+umbSOj75D+W2E5LsFPC0UHabqrnAjm/YmHn5jFzSFmNWD/zaHmio9zqc2itKVZlUdnI3QASDE
aXYXtI7XG2UXe0nBThDHFoCNix0PiF87hUVQFTLDHyMWIVZFuqH/3kCENyBt0x0e0FdlWH4moVkw
Rh3DcBl/AEM9tGdtXtPsPwvP4vAGvKCgrvFsz/kc7J5qD393W6P0N5vX3mvssxNLYaAHvwudJNP+
j4b4MfuP04YdNaIaPdRAm+QxRg7XDrqHAC0diLywQkgQuKOXpf+713lwQkNwIBMJDF8C4Zc+SHNG
gv3I8Rdou3v5LdgmO/ppSrkzFqQfpMM0gima38NriHIYgciGBH5vL6pXKAYDewkEbpSkCmZ3OH4b
g+hAHx4jwSEti788dnUkWlAV54fYChqJliyHQRUyecZoOM08FzDEh7P9gckjTVOioyEWoMICs7Dz
8x2qDzuoGJUNmBS05MUw/rgGmQRPpWVwuwwgtBVYanMTLmaahevosCvxfURJRJR1+0hT7b8I3n76
QVvfxNeq6zpzzkbYNZfevZO35woayiqGsd50kq3Mg3pdPx3Wq//byJFZJJPMTSjgHt/+v5PYWHw+
k/L9rwbU+PoRzq3tZ6bIKZwkVXHk9VTwrfKuvjOKFyuZIC4QY9u6XNuuAUIqytvXMSvxzHgrZiCH
42GkhqjbBeSO8/ZkGhFJJJeW/eXSGKULBFdbI0aRCVeZZoE79rP7F2HJ1wDexMiXSh5Os9bvLJNL
l8Pi+bEignDwMQoflh40kePZxCNbpTgSyeU5QYFq75LNYBbIJPQPT9DTcuiuL6ltAfqStUTKuEW9
jzdB7xcX9UwgNzImctZhye0phLAsyvrOq0t2DMZA1jOt7f2CGcItFBIChHzymZjR/snGNVH5Gkp6
cu3xA5d5yfcwUiPD0/pYYwEMhPWcEAMjlJ7r1AenNjBK9Cc5RttUhexao7WIAojOuZCCvt7rV7yI
XUdlBXHIuB6rMxI3ZwWFkdVwNaCAw2ze+/VsZyBiBRteJJA3WbMRHv4FzrA796wUif2TlL3cRNcz
8FrMQzr6R8c5dt8q1S+kvekELpN9RlEhna7F44m7an6xktf/I+D49s0xE5qmNTa1n0vp9G6vJ6iq
d8lv0DOrHzSUB/G0TpC4n4QregRbZCo2XdnXbNqSDlgwk0SgZKFnBJbzMSiHXQjOYOd7PP1ZE44q
Qlyj/pshQmQzl2z3f2Sz6GMdUR/HhjNQHIV/kxjMPNkW85w9JGAQ3hu3SssKMJK8Hv8AudeNHAG8
9tY6BHDl7FxHlEQcB9+EUtmTIlKkoUSNMRUqYDxZ0vCwH1wgPT59qoYX5jNpyizQxIH8X1sEH8nC
CrVuiBskKegTxr4nC6mr8Pmjg6r7PQ7IxcIsp6szwXHutvtvPpWjiJJw0PfXy3QJVZ5g4kZ7h8M/
L6prNFinTPculfi0stOMMyuEdwdpGBZiJx5On8KkDJ5cm6c5bfIOf/BEgD59aSsxaBYIG4dv215p
rxstZDhUiHojwqwsgo1Lz84zQQd2HkV9269L7qTrMlpI0qjiLy/oY1bGDY/CdVAnbFMpBR4EH8+0
b83uQTacdqdKDGlo8KL89h92yZKE/prxfvPsJQPp+Iaal0oYSHWxVPclVmfx9PpjuOht1QZKOgfD
8vQC0z3+lFwIO9/tftpUwz4cmVRNyh2LEec66+fjuI/oct7zELMXkxDMYrkMMKCp6dDzOJjsP179
pvD+2ExvXzDOpsTSqxjkjMtOOx50hipV4lUheu25ogTpM7NUOsnvXr8sEisdSyuIZhL2dh91cJyi
xsKokPrd+YoxUTAeMOx3xkrl2xXyN/6KnOcrE6qGr2qj0oz7QUGNEJkoEbtBNnY2xCDNvVLWcwHQ
RTCiX72xC8hs5bPes2YJbNcUpU3Vn2IZG+DS3zbnC9Pk+FYmLV8xPhdSritBTQ4LhTc7EJJCLdAW
wNrnnBV5Q7kzZxKPETpN2hMYJqOxD42kjuBJ90NDaU9HO3lqXZVtis6jfK14d1CY4kBfZsqAXCab
NA3ZZc5tyVcdymL2hslKc6tTTQpYbXI3VEB3ctexNHf/3TK4dKqSLdrHX5aG8+r4wjGgwiLGwt7m
L1Up6gbRo1fHcOMZF2ziZB+aARCCKGYiqdi4IFXwRhAlYInZfXOmeHRHds6mpQbYNIyzKFbjgee3
0TIrkvgN+psMFslRwOFuIntag68bOqCbwPFuWQdNfmZIlBBrIkc40jbW2mTOH0pPVKWqoAJjlkCy
1nGVJs7KQGPefVZkUYfpzqEfLBUSVvikV2Gf3zL0ZgF2OCqe5qEBPFGlGytEftb3YFFewYuXdmiA
GOylM0rCeiUr6ocvZ6uRIBd6jX4sYR/QzHp1AHeji0y71G0/VWp6gyEhao8WDGdml7gM1z7OI1HB
ADJp1FLYj9dNDKYF9L37vDxTmUvUdz23hNZaZ+56FCBcFXUmrorBBQz2ZhmmUGaIFCU6adV1PlWc
fgntA9q2Zz1W22m8js1YGfsYjBpeGZ39ODmBpS7BfudkGFCRUL2rgcrKpnHA0oYweaZi1CG5BnYy
S0t442xqprJ3xDhmK4QcHFeEv/iWKhq2OAHephJzSq1bM9wIw1a/lC9W2L6/Xr+tRfUUv+gTnG+/
Tn/WjIAWY24OYkPUe782yx0ikQKvkObTqj1O3XGnfblU/FJIxEoXrf08FBFjVpc3XRqt945OFmB8
dZFA+4UlKXQOzKEgXY4hZyFF4uAWPuRP66K2dzYSOEifQOEBl+nwS1jA4KDsvr3v5mP/mwCFup3n
nNAVnV/tL/3MRHyw17wFgmkKek0cPrl9VNUInvICxVmaLJyxVdPPVCxIfGcFz5ZqRgkqkQJAoThx
VIoV2Q13UegSimWl6yi2grM4gjr4OCuwozi+n4XO2nn8nYnCb8KSd3bhoinwM+DVCkM7UIgklsUJ
wIEZPAVYrEKm2PQTr8ahySO2z1JBdkRffR4l3QvaY+2VgumOFVmKsjeCThTL2++WgVaj7PQaJgqV
1tIE6mqeapTyXEWvddVuF7brXvwEDkYNf6uH31n2Yu/GPbcn7bLiDC4ATxdwhPEeyu2NR8eN1BNM
UBNfyghe2orqsZlaKejixLVK/HUTJCaGg432ai1k0jAbQID5jmp4JFOShFqyeW1Ex6QG9S0Y0+RU
QmmQdF3JRbS6M6MN+ZGsOSTyipHlCXjCmDL0Hs6Mpf4v186qpYWkj1Wjr/3K4g72eUoJZHnjrS2E
LZhyERhtSEafATt45IuMsvYkK67IydYctgjHFTG3T+7TVR8yLsQz0GdxryufYXGe6Sn8RT0VIe3z
cU+U+qknyoVDm4Hw8IWKAKWRZjIlpdQynH7YJ7mibTFqt4TJh9ewCtf4wxNbwldD8ZfU0XKniaLU
jkvU4Mtye8eEvvOkZ/LSQpeZC0l/PCfz4AuwbbwbFxeLi2IIpXBfb1+rS+WrrsSuGDtb3VFXibUj
Xs2xVWDTxRfsFHxasTAcfJDJ/cja4d+iRugicNaCf/91Eu21ExU+EbcV5Q9+fSvXDeEzuFw4ZNyc
EpVEV8JxugWC9XeC45+DbDUR/N7ofTtsFUqUVmDsdlLxvJGNE6RiaM0NXeg9n3sJTRVo2/oTu/y2
g3DQlq04PkBZewSzNmT0IUYESDqsMrdx3qBuIufnvN1IT4BLONaHdqQDYOF7VU3vJjkaj75R+SP4
W7kzOPsyTF1ZS8m9QIluwE0FCfiYyfghXkESueQbtknWxDu45UqGdWxuyGcanP8NyR/4xiLEBlpO
AQdjxJmfJpZL75aUJNQIIdiuR09K+Cj8EmB2U5x0K1HOWVvv9dz4uc4gBZA4XlMmywbmkeKorTJo
jP0TXEv+gpKDmE+fXZSpzw93zC4pZhEDBJHITbKN+oN9bXCSxjV5YwKrNMRV4zxZ3l2nEc5Z7r0Q
xe0+H8/SCNB4fcfagiD5AnZo5jdGHzeB2lVfV3Hg/F/1bQeEsOMTEhWi++Y2GokhZWbO44a2PCwd
n1HPplngE9WH0aHiLBNgC+KATVbSTl5TtbRNMbLJuyPaOQQbyBQW0Snzu64l0Ie2kRbfOUHeZr7r
5pcFmugwmcNr/VrMlWJ54H4jlcUmZ/YvZDqZxF5hg0nRw7Ctel/kOjowY1hIFXx5rQW1o5BSsIKc
huhbvH5Yb/JU+7ATFGKX7vAvq7fqC4sA+sQ4waS9KLxzUG1DIPSp2zwBrSGdsgv2IL/j8RuMeBGM
RVmz0ubgAtUp+L0BddaSssu/Oqw0Rtgg5elWVieSrIHUkFL+58TqgNKKSKbf7EMHBRxODF5FqH4C
MvICfrdzFH7rxcQQKOHobtpueCLAQ/aX7w+QDFrRCzkPCa1aRwCIrwFa1MlC4fc0MisolX0I9EJH
pMoUTAcDysRM+WVtGTJm/s95CWZ/2wyD2KBsb2dwtcdcMADk2RYOTG1mvhyRoQwesvAnmROOPgYh
MzRQyPTDruM2hSy/T4/LFApmWpJgdz35+InfFDjWGlvW3zIcINJ53jE04OxHlbeXAgkh27qBNc4F
+UH/mJyRkPYy/Tx43JX0cgFreFo44iDc+tyz4KEQ6nDTnaWAHkAih2bABvucc0YhHIOrkqYwNvpR
WFADKRDHJybUODpu5XnzsXNXFFPndubihb3OE98C4eMvpFp+nAk4hYK6k0daaGSPxdD0oPCDZH7b
Zm6r/D0OmIBD+LRf5Yzy+jYppB/GJhpdbivfOWmLgJDKSdbr0PpXpmNSuTsTN2wd5sdmtveehQPh
HgQB1Ws3X1lniKz4dgnSbyCONcX/g4yyPxog3UppKP2eJ7BLhv5QYkca4oz5YNxAYiTd8tW9RFue
eO15Ur4QyXFdmmcA9vWJP43hgpIG1MlXHxRaiWaQAhIaoeKQUFvb0LAo9rdiDk3i43ojJOQdvg4x
wlVZkkEUa+JPeZDZzomutIbqjGDUgFLMGKfOaMEbnLh6MwjqRI7J7C0LwL3FP+LV7WIiWmnVGkqO
PanDKTL7Ndc0bMQxuVg2xXBhQF0daiVFPtIAaJdwuzsQHAAWSbE9hmaRXliO/sV1GI6hv1Gz4iz6
zYh6Fcswz0B5Yo61qNTfXYm9Kgix16Nt5HTTChw6wQMrwJXxNTgwxZF5F782VTYq7IZG3nmOwPTd
/NlqBuQxKe7HtaVwn6nak9IAEqQ1kHRpTAVn5M6JRd4e31oFArekdpbaODznMOVHECt3JU95Iu6o
XicCCS4wyJHsmacOkKjVedptpSQ3ZpuJznAkiLy8i+NFlH5Vg+i6tyGgEyDNqtaW1IFAXNMErbtT
VUe0rAfBobq7p6y4Oaod4l1EBzCHg1nF4kZXSIRn3dDLu+kGrqNUSgc44syZgMStY7xmX+cPeZlz
fr3vAtspGIj9k5fuvdiYeCYA78YQWUqd52SyTAfARiFHCfd5R9mAiRqIrb9ca5iDY/fiBWRsICkY
pxFCTsVoQn/vWYabzUPftrLbeXqc+SW3xmtchzsCVcFEapva2T2Mofw5trUBmTxjqtXBtjAMrDBr
vPsyp9g7aVIqPmCEQbTE1BUjeYH9OiIGeVExDxavs1lclETwWj/JjUp3W/dBQk9YFNfydUPdx1A1
XWg6YeLdVufMlRCaKOnQTVqej3bipaQSVnmywVlPIwxeneiBd4jQsNAjQuOEIvj5Pt1ke0GmkMrA
zT0XC7L3UyJDsJ58DRupHHnFNBn703e52GeFSlTwmH7RUO2iNbFwxYVkhqPonOunotCKo117nHj3
9UrTKA8/RdOLIC93oqZiZmhqhKZQWvHijaRAEtr1QARQzHMhasF4bfTOJIAxibPrjlAjh8n1xctK
rq0Nyam8yMhIEpM2QY4ZN3rxOO5TflSpaYCZhKosrNgDYULgZ8thzmgZa5QEUWheLPRumOKWW1JO
5LFYuOdMKWwww04+qrQFyYvmcIdTcIJe/P53iUnfKdViNh7hgi+HIQG0UoWTBXDfzSK+77QfS67x
zsAoZR3woxpIdIojqSL/5CDlWUU0FYaDHimWQ16PXiX4FCxqf6lHJ1ssF3kcYuex/IaZY3iBfVc9
+7ZqvgB1xQzzzcDN3cLrujtfKSoyZdwMirm2TXOQ+0hZZmYvIU2SfQ5Gkw8X/qGyErMVXgb1SIO4
cUqNY4xBgH2TV3B1ESblQxr0CEEG2py3+O91bYSqTs5oi7Fra+yZH9k6PhbbeY1ixw9ln3swxzts
6pQABH/bEafC9WyUGgy7adsyGaxPVnX81FxKF5uQ8SkFjSdjHTgMvQ1pMgzoFDISmbG2I7UaFNjv
EeeiEwtDUgbnVYqy29uzRtR/Q8zvpvGKzio4OxVwQmn5DyUgKbob1FRvq5s78hj/2Nrp3eAG5FCt
3t/i9ZdroDKyM3ubBKP7EuqSQCVX6CE2+4MitM8ttJuVRfbzL2T4fGMvaXGT9VmDwDyj6KwCyGDa
rmbjIMte4CuYg2V52gPNWzYL9i7SCC739uTSubh3z/0Ch8dmJATnevhUhhOEAxIP72uIxJZ6JGY6
v92j20t998JdPVg3vhOpxRMI8jTOF3HieaD2bgDV2/ytMXg3zhFJQxvKykKqBiF4/ISjCQdJeM5Q
QUGqd/SipWIf8TbGaQJTpxyavPPRMbtjQtpStyWimBJj93K956Ud9O5Dq2AMD0gFs3Y6Ib/eseiS
TCveb5fg34j4lpqHP7BBPhPx5j+cmEB++B7Y3yCmsyggu8Mtr+MBYBxHQSraOWFJ5NTSPb0RoJQq
eXbWnsEsYeCGka6vKMzj4oxzrfG3+D/S3xQSN+u5KhL4Eao2ht3Gj6/wog0FpA/RGUfmS+yPRbgD
534gWgHnvVXQlYaNVsF3BYg/xdecgC7IMuwu7QeUZuornN94ojkTt4ap1M8LFIV7v2a0rt+V6WSq
cH5slfMuKQ2wtGs1sl6ePWDuD7iwCTtvyas+E9Vd43jVph89E6NUF87UKCqhsWbXYNTBDC2lD32q
Xdeck8wsKOdSU6uM/uwXibEZuxKB+9LIJd7QtB4IbVAGQ/tknB4EmsaGEIJuKCNmgAoEZWk3oEjK
bZpz+pbU4ik1DKWqoDg9Ur34wmA9TES5LrvhNnuSNmjhvwKR5Ut7YEv44AhzfbgpYSuPYz4CHz5z
qUFP+4lf/X8wbICOEbUix2HaNabYvCGau1yE/JcpLglqXF2Fs39p/6/Zp6JGX2eiYydNpzsGByae
gVeZlRmBPikJVsWGLttuFxA64FZY6uuaLs4+kulYeIXvUk8BE7HQprkGQmm2QVzp9ctpwXXGotH7
PX+5crplEC0MvrDmmbD+Hetu+ysESN3wN4di3I9jzvAibDvuK05vbGAJr6jc6LfCHFGHyBTunzz5
msfaVj0u/gDGl5lybzqtvawmHgCxPzpZaqOqgKqENXndc+Kl1YsGcaahZdA2PvckNaBQPH0eJJLU
SAXPv7GSKCTr3UkQHf4dbEfZwlpYFZpBkpgtYxXwe+a/qApudK6mVxGfCH40LyRA55bgG00FUGW6
xWHVv1LR8tUZXlVcnx14YEpO7qAqPXjuo7pCm4T8tdn7ouc3W7vI+Rf69Q3UBMOkkA9JJjVzBt4U
UpFz/wqniFtpS2I29uWl/VkDo0AxFI+cGhh9KmH3jbqbc7CsulgG2Fm33gYn8Q83orqyOBWEFM6Q
8ZOsUOXkxyeLM3Ab3N8PpjReIToXze3GzhjqYJtWdDWE7uzQjbcK1eNL6tyj8tMloIZjZW937Qsu
pcrIKZvKGkbm35FDbIEkOCzmQrPBaTvcPk6azEuKaUwYUVGqYqFX3VVP243zH5Q9+uU+w4r9ZZkW
iZHOoQi48IxhLvUbM3jlV45MHPJ0t5TmqhxWazAz0usLgeWwSDi0TcCUoIxmu8kcxzEF7mSsl5n5
peIpLqDPjDvQxqmAz0x80x8ZAg5OcC10mrF3Gh+OBAL4Sj2a2z+gPPHEZt7yYWUrk/9AGTIfpSCP
Pime2nhdRWJtKMPQsI9lOZK+5PSuBMY+N2nNE7Au2hd4aAF5anQWoomYIFhCPO7PfZgD9fduhS+h
nGFhVk/WGECD2HIAmuVnFHTkxDznbGahwddG0/i4r7ggm8MB6iF66w0r1WkoBIXDy3Gx2CwRJC6+
H2qQnIvxijqyLaJR5ZAoxRT0zpN91Is9jqN2v7XuTmDIKw03gYDhhp6KWGEMwhEQEZ19eE4kDTj0
atlasfW2fzCFD2vOCPCw/NB5LQSEcEaNTgNnWmhsBbGwzJG0SnRSHOvqUye6TEY0EIl/gTf2yMPG
t5CZbF6VemFA0SQ16/+mE9VzJPBBI2pyAg7PxN3y/dZ2sCdmBlkIqfErL75+WCfMQhld2+N80xq3
DVWQOHraUdGdlhjz4LA7VLrOEYAkMcSXTT2KJ9XtUOucBwv7hx9FyEYrwHuEBXWmWrngUoT8ISRx
3ZgJZfQy3s2JTrUKOReB2SUyQQSO7sQSGu9kfOp57XQSorAn7RSwXUBz2t5QhthG0Ne0WUMXBbSd
y/fofNJR1TdclEZz6ta9yty3sPZSZk+u4L+XfK1CdzBWkztOwwQuWFx0FTSgESqjRMjgLPlOJOvA
uZQatB24SvLLbVBQmZzIjCVvJMcKpTV5rMdRdKbugmYt4Xk8SdZnIlDbORCrd4cQcWHG1dpWvtCh
TTZvEgq8IjtMa5KqdA5cHUvE2tyIM3aHkxwseZMwN2UzHaQTd4Adj5E9Aq+oEAoVvqa5eEAXCSuD
rqtFCQ3l3BlNxN9En9OtxRxdKSs+Sgz9y1SOm6/0w/wRlNOKWlGixtttfwWZHa+6eF7kEfGP9v2v
Vp3J1pFhyhgzaEGyBKwbKancSjONtYxbfg47+hBl6E9sEh62cHuGstN121vLyH96ZSAyNJonKASh
/a50qgZyJYvLLvu4jO+3IGfEWqYTNEyzaSsp34ilS0H7NHPsbrsmiu8FcFNdEfFKkG0D/F6bIaFW
JfrII1lgdT5/rMhzvdQS1lgdhRAB6N5k61Tj6RfK5aIZ6iQQFyGEIO+kORTCyOvOeSaeCEN72+X1
byofMFlfM9PAgFL85VqkcNkdI1Z13f6RKtbu+5mXcIf10O+OCmu6KmXJi7+oz3jVi/Mw8ZIaCHbu
SvRYmDSS8492ZVOZd8ja7OwaAaSF93h3dKVHx89kwKWRXTjxF+aQF+lhZdjulaB18nuym5e7QCjI
f92Bn4xpBNcjCRMZfoPYM0ZTGwhRvlTe2G25pwQcsnytFAXA8zJwe8B7AOQixleMw0Q0jFVpedWl
8tsroQ/e8aFVn1w2/+DKJ3KkN8eB2Qew1bfXaEBxSRFmeRHR1vmMdGVWma1f33aRGWbasoP6sA4h
Rx5VR7iVAoCHy7kgcVRuxtQNOIO/KP4248YA0Up/3ZcAdRQeULqcHyazkY4uJFqifhPB2I2Khb0P
2DPYHgHDFWKnIeP5JObGIyWoP9BCxodZ//uP6cMnMlUNtXRnx1NrlHma38INthheu9kCD1p9/c8F
AejU7TykbD7QFiKscECJTanYqfPgOOOI9HE9JExY7XpiqtbEwRkGYk8SHIPVaNmk/6gW4DtraIu8
3upETMRxgpMp6bYYIoF4KeRbI7119L6YG73l26RXqYberggyhvM7PdaCXRnLwbAQkBY1ty7vdRAU
SiP7Llb+AuZDIYFHFK1ziuCf3hej6YMjW/gllKlvAHzwsKmSY3gydvlkN2Np7Bkck3MbAUXIGl2G
xWCTOSoV5DswARFf7mxtCJ9+urBLa5HaxHw1eF890cwCFb1mSSrpqxE+V58jcvVbKAhLPn0FSGhh
8xHmMZkPWqQSUOiPnUhFF/YkCVcUm9xFmZubhKcWBaoVUnE/IqVkHHA/9t0rRIoaHxF6jQLooo5t
/xiBCoeZMw9uv3x6rjm1Ol7zmaQoRyV2xeqDosz5P501cC9USdPWaESleTYIeK/ONa0e7W0SFCzG
sFbFf7OZ7T1ddxHuS7Ytl7Skzt9djNRm/yuJqUrJ1N0otG7r8jmuW7dnpSnIlMdQy0f2fjs2waBw
lMUDxMboG/3f3T1fvtM6KAux332KScebdHiblXRe1hBjdj69KvXAmfX/G/nkyRhIbilpe/mpy0w2
FmS+a4eZ22A/ZFRv5vUnhx2qNUOg2Ceun77DjrL6kqFw6jmN3xFCNAfy9fRxAqL9O0vt6nXF6K8j
ygqgoLuprVXGQMdtP8uIrax5WZpMHew+i9efqJ1oluwwH2DOI7PrIRqIs9IILRu8D00Eo8n0Vl77
TF2og3iwLa5pmgRj3udL5dbg3aRpsGqoDHy+Zi2iaWG02PvHcw+avNZdfZlrPkX7eqRFVFX/OckA
nHn2FP1YBvCz9rnYD2SQttmU71ICbEzwGTFfO6rcPiIhtiih2hdQhKFlqKMkLdB4JjYYpp/+YGxr
dnewl+F2Ppo2YL4cTirCYBc4dIaxGk2IshPWn/5XtDlBesP/hUISp8RHfGd/a51QS1S8bVgqlIhJ
xPPcK6z71Mp6jmszLmzF2aLzbzMvTqVoAR29GGEOo7D0UfshjDeiV6OV1nBrKD2srbp4VLQ8Luwl
dW2SbjO+LAITFuMF0RkhRDFLSSFguuEbr6zi3x5KwUymVR2VksQNrExtzHlBSEkoOkPDKBjqcFeG
Fq4g4n4GEijUv/0nwaLvv4cgGyhf34QhZdfbCVCZSUb1oWsXiiUmy2F4SST41X2Z36/0ZaHDB1Zt
Q8hLkw7PYCF8KLmoQ/QayPJSbZtmqpREyQTJqPKPjL91R8S9g5M7MGo5JmtweaS+WtIWiBoFobwe
165A29fGWpy0X/mWWiwW1KWOmrkOGvVOjs/LKvN0Ee0PLC2tMuePXB1YJ7+2CwRh+8adgS7pBcK5
VHE+LXO19J4WFnP137lGZIcPPhvT+TLDKQMUWU4jSfEWv+pXLTO3wxlbAPJiYV9Rl65h5kJNgPOC
hboaqE+GhmctACLicFsXt+waLNscAJGKOYHx0dWfb3VjLb9lmzPcs1BN4KubAAQuNWe46rF0YGUz
9K2CISe6PTYM1KpYhC2MumMuX9O5fshcP6mS3pyVEWNsC9VtqsVaYaPl0x3BRL0s6u1kPXgGmi89
V4J8R0I+JJSkIGY/EWyrKJh+LeGVqmh4KkC8B5Ow1zpAxwVc6nf4JSbiZp7YO53a0bKRk0gpt9cw
86c9sSzaU1jtefCGYoBeWlfK96eX6q/lVvWA8wVEJR5TLuJFyuiq1U8e4prOamorZ8cVl0fUoTQV
Ddo3TGqBJ64LLCirLpNFEPLROTCV+iRL6aDFYMdBSPn+MCXx+2dIxEDPI7/wlkgKa2E2iDHjnVVD
14LwgXlhE/yMXpDyzdrdatmNQLEdPPnOQQByLwQyA9UJzOhO2U7EtRxI4e8NA5aChm6fEGFnwoL2
WqEDi/X6QjnvYClcTe3cs23Qvl3e9LXiV18TBrY48ko5mi7vQe0suYZWIpwzdueQOkI12hD+XqCP
3jsZgB5o1LWrwwkS320cIfTfeU9++IU1GxkL66M1urNe/GAEg3ZfvEsrVzMFfqsNobpn4Ua1rWBd
y7MWzM9FNBpjnpVIAIlILOkBDcfUqoc6hU0a+VIQWX5fqXt29P73s5wWh5ZqYCODvrywNofcsCTD
ADIsexnZXUeppxm1IOuBo7Lj7+GN5VP2A5mJqNgG1eEFNTsubEcCTTk/ST4nXASHgD0hZeVBrzln
kmxYKofwNH+J3/7Uw4AUjDV2AW6iH54xG20XLLs2m5ZUlyF2NhgVHXUqPb74w/yukvIBezSKveAb
P5kwgwwYruO8RsOTt7Jc0oAYRhWPhlHqhnl9c8o6DT7/dfesIwcr2f4lfC1TljMTzqFxCoyzwW4k
SOS9EVtmM16lEn/Ve0V+QTMFlFCU7s9mexri0WC4gdpn3zoqRV58g1qatiUqBc0+kBm94rW7l/ho
PQvtr462GFwoKPkcFo8ctJOJYs4Uycri8W2dmJgsIEfQi38SxkcjWIhu3lj1NG8BY+qQnVjGYetK
QnVnD6m6vQb/ZsDHrrhEgV5CTtsPxzfRZpOr3JWpMLPpXIx0NZrqzStQ/L3iUwEWYtxEXb3a+Sjc
wMmGqR86NRXNTKjxP39A2HhTfvDsOd5hrA3BtQJCl9ZFmppYQ5WmoLr/bd6ZlXfB905HXf3w0Rwv
AXnpkfE+HM2tpQVwCbZ0rN4/Qu2PEM/V8OA9mkI0OAei2XVXAjjNqhNjAcNVFfPmcPWsGVvvtgEP
sKtxxyMeSLcUApTBwXQmbDff46GSRWhQUukTc6Fly7em8choLfwsbYs1lg2u/v0521+y48znaaPW
c2Lpsds3yFJ898ntheyyxtnWiZxmniXpNDp6lz+KtJvY1b4ygNK34xLSZcUBUZQvNYrwASGrA3Gl
O6D3LAEA4ZQSI2mnV+jjyerMXMllXbyCNf0e7G8Wuz1xyvuN0VKaoyLx1YZwSg/la2JF2ERzaKBM
N+L5pdMDvPqzl+h9fC0NZwI4oP1s4CyxJOepq8HX0kjAc4Oq2JunYnTeUpWI2z6ihObUGdI1lo/o
6dx1VJxTQU6YPSLnGHwoNpwZkRiZK8PSSutUZca6IUvM/TY8iuU11kijOmgmAulZp1jHTyim3U4i
SmLbG9cc2eix2FQLUVFNfA23H4q02blSJl0JeIyFKUdAyZHObIhc7+x3XA4NCrVkDJ4eVPiR1/zY
8ZvJ9/Q6k+wyAMgSg4GbLHPhXk53/Z/fKcAzrcGlLmwg377B035KWTIk2U7DrR5Rr/Ml16KZPD2B
KwlSJ/xB+ueGBKDh11h8rqNgN+byJKqyYYb1SicWQ6fbw9vYCYmfYaLZK6MGiNWCAk++SQP0eUIe
16zmn19vcnepWfEa10ZKHzJEuSn6cdeEWNLVXBmPINkhIbXZOyG11YcVORzspwPRSSh6Sz0+xiP7
wZsQtQ5paQKwrvc2/By6Wygr6T6mc87iQ+w32kFJlOnCfx6FyQa3/YDTBKTaFtGMH82Pi+JTvkyT
NGSG2/TCqspjNuAIjhM8kms7hH/W5lvHAMnYth+voZrGAu/l1Vxrnaj9LjRS9rrq4hp0UTL6Luir
zKzbi3lYzEDNvebEQn6tFgdJ0yQFwOv8iYiP7z3xhmrArDWhxDO+ouiyVuYqI9/DN8zTwsF95cq+
qu+/MrtTzGqOm+nvkVO8UPVlKasvdHclQ3cuQbB8fWTRqpT9NK/lRd+1MGzrtvTBQuz1jgvlWvjJ
QEUthGWCtokwkopESs8gjtw3qSCTJKA17xmCpwVxbkB3LecMkPfhvBAO8iTja0ulFMz1WGR0XkAa
Zg7wmdMzQKKOMLC26+h5ebxue1401iQ7viDZjJ/HQMikMjcKPSj1dq1iKSgUMJB/8Xs+Mu170WXr
xCZApNqmru0WiAhP8eQOS5rFWp+mFGLRHXMo9JOYOystRKiMEwY3dd581NsSm3AYAh+8Sw5dgOQn
1EAQLdAfscoDBpMd5K9jioO2gVCq6Qx2H0APbK8Q1vomFpVUtbWNYWpTnM5WpPeLT7vLnn4MVfVX
z1hwRCwS6sniA252TZMJ8v2fXxvi0H7l/zn5hm8bO/8LO8GCavEZYzb2VNXb83SIf+2OB7WkZx5l
nrAH9A71JzXztxoJLjvJ5JIdux1/VfH3LiPM7tb4WtBsytBqpKcaGUubQAcauxFuMeBwsKHq0lYj
oxZRZUS/CnAhVh5CqA5Qp5F0QCj9UbFjHmTFSlpFAkAR749U06S9FbB/ifC+HVG2qHg0NQZ8b/4U
RByJteljqbSVN9bKxdSnMm/XDcu6yKsmJeu31X2lhZNbeuJxBBbz8l9mEJsRsPeXiFMLRvTwc/iS
uQcerGY7jwPqVY8Gl8LySdH/cMZ6dfitXhhL0uKk/5xQC6T0OG2HVSkT4woB9fRFxjRx3MatUDVP
Ci44aq4TWHCVAoPOH0QIn/1IU0jqHF7J2o33pVdedrseLJcLEZAtmsrzJrytn7VUgD4HQbTwEhXN
IzGImfly093+iIbUGUKkrxdzdgIWlssLtgrD60132lFMX9M7vLrvBOvfWXUpwA9hBCVLbE6pHlVM
diqwvWhG0RjOtYgReSIIgfSonDBYx6N2DHem3m7nW+x7LuwtGcidyA0d8OjI13xzt9qU+Wc+EN2y
U797L6BF1O9kgRjehamn7s7bT88VVcbJkzUhBJeG9EI/cgyDXSP9jc16OWv1Jq57nwCEdpAEEgmi
HgQJChHKrVaTVwnPYlXzywp2xHVZaOcwBNvbHYHyl448LozVRupTmzv4qazRYb4J/JUAabkRc7qc
8jSMrOVZ1ZaSSogs4n2jYl2R6tO2ThBTapvGXEtZsPh3b0XlO4s1iq/dehksUIROAyQkoGGgAsgV
Bn30qz1pUXNfEbTrmLIurI6GJWD1sxZGtl4WS7oQ5ZILp7w9SuIvqzXUsUmju9yZgOByKXkmGawt
2IRYNsvV5IsSewHbacSs2GD1ElVJDC+2ulrTu0YERrDSD0bbcy8EUVC1nbtG0CpbPznY+qNMacNc
RT+qhVO0OJPbCN/qMwNCQnsgZF8vOwPxHyVY/qKPDabipio8O9ABqlLDYfwRBqAj1GYiFuczArHR
wCRivB1gwffL6PEN0uFNVpEzgFzRy7flZ67+bnqOhCJcykrYeQ+wEhj6nxCcm91uefFCyR5M8e3L
WYnBBFR+yFqBZ940QjpxffY7MXQ1uFxYFSw+5mbAiAS5FmZzKEe2Owaru4Yi+SiToPdJ+kU4ai5h
9SAIXqRwWSEPathVG1JWkaZwXr0B1vlg4u42zxBt0boTM5IuHZMRmQqMP9GYfgzJJBpYwrpSB6se
mkQC6dzfBYHgld3a6AwGMdUM2/LzLOVEp97xDYFQ+HTevwwX8N0vqhQ/HXRNjdp9rsX3XhVuWFZu
EaWQF8K+y9MpoftqVFKtqf8TjkJC19Z9wPAb1OQEgKeqvLlykGIsszLm5Z9bHhLRqd1F6lDwMJ+0
VvbsZh5tiQCK9bLlTV2IgerxJ7PItvt/LGCihvgcXhK0qg+p+uVpxIsrkCXDoQxC7p83p/U04q2C
5talHCqsfoi/Tb6zQoWrEuIrHNhvPzPqonZJJdT7pyPLui1gRM+QuifjGvCckJiqIyfFDOde+Ibe
QcIO7pKQKvzFCptfCG2+aasP3J3jNg6Df2+Xj/ibyQ8CSnAK+0Lam1aHtp4gg+bqHnMONK1jJ/sW
Mb4SUfuUfAnOOAMR8MGJCOcOu7ur1uyKofaWodHP4E54vvcRify+3qWANLZ8a4TPjmibeNvjv7fx
qSFzgkspfo4SB4hnIPZPMh/W1HB026S4+xXBn+0XXhEwdyKsY2l0Kq/8SVzW7ZydvxvzDhtaoenz
XwoeYtK3fgBfO9R9ay3hW3PYG+l2WvTrV/HSKmUWL3xLXBeODPkkilXqfmLwxpW92xOi7TkjOq6f
q5krcSEVvMqif3vqsX/rHCu+1rsGlL9ZWBsI0BRhNUa8LT971NgHz5qYfhxVScuZguLgIq00e2qj
izQHG07ahH1/49ePN7var4uK8MHUxy4gSjLLVTswbkklIJh3ylGQ4QPKn6QQr2WA/kz9vRDTYLZr
kRROC6crk1tbS0YU1hzikCtu8UdI73/ZYQNRShpA2SEt1tRHLlGdsPzCYxY8iyLUN/vwmJ+5CA4o
IOEvkDaX9YIzpq2tmxlUSOOlgMw7WnLNE3eTI2E3dDjyvwGWQobmkb6B/VkMIHEAe1SXpgXh/ILi
D0lqLu8W8kHC2bRVU1zrR6YNyGApvnx6+fR6046Rfnw12MmVTiXzrdMFdi4H/WkHtEr2GCVfjQtc
x4sE/3OH2MW+J3dikcGsW28jpqensOAW/NqrwURh7ZFmeeK3RksoLAt9HoYF2bhW/IK5RUQJhPxj
FToWNpnbhBRpOuJLPPYX6Svok/3SqJVtDqzXmDUojT9b84PEuVZhWf/M/p0FnwfXRA6fkm1vo6Od
ktQqppLVoZrsrWfoaXbqIQSvev7SLv48tTxyPbjrEm+A42fCQk8Yu4DyEtAcuLvSw0BchZF0K4cu
qNVxfLZ6XXsOmvQYouEyKz0+fjQoOVMBTHOWoJrkWD3fz8r4J9kgK+XluFG9Ck3SCKKgHArKUJpj
iigLLi/j5J9eRPp7lLl/3k/mFAEvIPtTcFduuixt/m/ojEbk68TNQEg01G98/cd5lc5OKx7GlSUQ
YT1cRpT8NjZUwKONeNtj17Se3VdBvzdMU08Nxmq2Ju7tmcdqwGYmW5wd0x+OOC+0UNJVqxATQSip
RUNOYz2tRqr1P+YWOUWFJnI1y3eJ4zEdSrFPEk0F/che2i2Yt4K+7mpoe73WfIghXyBjjtx3UA8v
xmf5EDsLmhcdLou8dwT3wrWY4ifJjayGROTQ76dL3i2kVEzxZC4r8cwtOJif5IUFFfZk1F+0Z+4F
AdFmiUcSr7Bm/dh2GdCGT5qLM5MJb01O15tIn5IyagpGqUJjHUmk8xTWeKWYbcsjygki0/iscz8x
V0wisw9VFdvVLJjhAiMVrQre/BuQhcKEhH+o5VFZNw+syQvoMUxguRW0EAbhGoSw8SitZG87cN6q
np/4HpIeg4jVBm2ZRPYcWBz9s9+9y2t9PCyFmpF+ABfMWQJvt5dOCOpO4A3JrFO1BnKcRcMs7Mfb
ZQi/dqFeDMz3pb52l9VSG5Gs7D0SZY3Npga99b460xEGo2MGNspJogs7EWC7gonTkE9pJ6/awVBm
xUP4WHp2cyujb4wMdYc6QfuX40m1Jn08uAzb0hmmvrx3ZmB5ahz89iiR7+GVAFHupRQIx5Yq0ARD
wjozUp0R74IbYLuZ/cU+k93qupI03kuDWZQ0naP8Uj07l3QwaXsjTBFfcI/+ZnTyoJXO+QVoSVu8
1TMrqetoiZ69YCg3CHURYEpExZ5yDiwaXxbMEXy4QBnNkthlOngtLTPiXqa3+kM+hARvDpVWHfEc
h6lw6AaIjxm7zZQjZM/b788a8SIDTIgDfJWtUTUZTHdw9lbPB4GSALwdKeiVzltXWxbMCK56z+j9
jgAwE2z4UB2T6i4KgE7VnnGLMVMY/UCoPdS+sBkkAA2OY1QcRRelBILqDNaE6rVebNYYkfWvXEjW
LuCUqHwezplG0ItLlpj8WwPnYbMRBYoXGhSzvX5K0jkX/CffQkAgiXA+5UX1h0kZoosu0q7RYnOA
H51CQv88dtxnPQJZ5mzTNuoaNwManChcDocRCAnXbfOPtuAKwvNVmljCkvcTjJ4ZfrOvgx3KC7WL
YDil8nSi/XjPdfT0aAtTjPaT/mkH9Pxd9i8/nkNc0juuymMlNwQpLCO4tTXYmsHNe1j042NPg7Zw
CJhuwp2LH7DoN8q86bKaCzYxocy4wErTk/VVV7w7wZt+jne6XlvafwC3rf1FyWgc2j1/x9D++m6E
RrjZbztu+5tHdBOmwwqOjPVR2ovHkRBwNkssxtkkQ3ohMnmq3Uu7iHe6eu9qmf23Sb8t3dzdmA6V
eiXdi+3SGhVNmYv59XqXlrTu8G0/QGJN3PXdnaVagd3F1TIlJIQg023aLCfPXBpL1gs2FBQawBDI
U4B/d+iM7z38AEnjaVO4ktgEHasWqd2Y+rBfkFkNgy2Uc1PgyeTjnsLKUfh9jV8ok8fMja1F8Si7
gqHUCJcvgsfM8vZ48SLB0ztxyKqzrXK5SkcWiaQEyQrofsc5ryNCJpRPrM2+DuVwxNpkZG5ZECji
30Nty7anjzvhykM2l5TAWHWZc/RCm0KLaC5UoaKSsOtXDpxw4sil3KsIGubWaAPqQP1zzEC1iQV3
r1Nac4shLEovuwEd2zDtseW7osM/DMO1fS/Nih223TgBN+NzA4ORlLFJe4Q6NCiFmlL+jgUkRF6w
aImwt/Z6yhp4+JvDgX9PVj3o/QKR241yvrOwcr9LhnIdbrE16d5rnbpiLCLTQF0QNL4g2rDk+LCn
q0bYkbgWhM729vOY00vfCZGHzBqkR1QFN8Kt7R6nqjiZBX5FLDFS0kg1ca1vKwr/W7yNS2+5gZrQ
dliGzBLqv4o0W51EyxuooRConUbdflB7Ne8mGH3VxIiHpCxKlYG8fUy3uRpMGXhxJw7g3f06PYZV
wUAHBjhvS1aakQFiwd3DpqNXAJFE1ch/wGgNGqCkeW3sq1x3m/98Dbxn8EJtm/oPeYXE79qJn+DK
jyKjUvyNNuosrTodfaAPC1cNCI7YlmkQ1Wuni9XFb2FzNIOnNwG9S/WZkruDHptd5WDJ04uNNdo6
g9jYaDrarwj25yMmeg3cmJU9n4C/uFOwbQGZlQU6dgpmrOLpEeNVv1uyjQM6gc9rSI+6RLGyR0ab
yyEbtW9yIc3nW6U7OuGKy2YtF/ehFDfjQOlpAEvwr5FUMQXD1KmD5ecHU5Nq3ZGA4T6IxyP8n58w
BOhtkyMw+TJXeBLIFdbYIC5bFVPziuTQEM/6wN6xdeNUK44TrHzY3/nYCo6wbIPD4fsZQg+zGSfr
uBI6UFTKa7bpyDwUiGasCSmhynOCi1PF9VgbK+9YQSoUfYGOegK3wDBC5rvo11zuKF2zd1x5Y/zD
RNqxOdCElzE4rEr7ITaMAOgnJqbA8as+Tf0AwMHTqPUzJwg+evbDXSKHP++mfkRiMRq7xDKTf+GP
vSNak4OvptP9fg1npIWqolBoz75N9A7Hw7lW44Lef2cVetNbHZyGzfGA5l9Cao4V9q8xiev1T+AJ
fWpNbMmCBB57RBsHzEMicbN79jg/PBOqtwxveZe/Vpcra5udEHBdyiXYZWn6FOt+TDxFFvNQT8LN
f/valGCsaOa4AgLBqz4ptBGWt4kJLibX4XAiMwDsJatFKBHml2meLEjkR1sYencEtlKq6g6G9rS6
q9D3XutWCgWEQMQmhZmRli8wZ1zBpIxIjYFCclsqvGPz7lWzfXFocOpMrekznhpZq50GAb0bhqVB
IWVhDTwOOVtvEauXrV7CrJ40J1GXbZhTHjiOpjm+KbiZfIL5Ye3ge1WDWz3Be/N2RFmg2NJ9N8zF
dnPexMcepOwk8STQ08VNpqroJtG9pR3ClIkiw4xk+mu4CvME2A+Ho/uX0kxlxFfETbigRZ0XeafV
EgXVMydtWkuJvN9zKZqvnEx4YqvujWBwJ2Tz1OZkGqxGRUVp1Ns/3DFIYoldDYyqgTspe++Sec+i
yN7+VGkpDsakANyibWLHuUWDcEqfWuVEazOwfWvfgCNqGtGPc15tVxoNybHnu5s1FizkZE8mEtJc
RJfupBtEesL5dYsLJDiqTyl2Q4JtQ1U9t6ngbNKPeyGeyhvkPYzEPe8cw5yEDSYvoexd7xYTS50f
LyLdH++t+35kYI5Rvv3CyIHRmZVnMBji9XyqXsprTOI3FPOijNM0TKqRD8d7tVM3j1DYjwZ9zO9h
E53fO9mGaABwN4HczFZoN6cCm/vVCFU0zE/Vl60WsavPo7R93qtu4zznkZ6ffxSrSZUDhtGy8uji
6lvX0wY2LUFQILwpxUg5qH1X4OgX5ptEtrvvsS38joBvSgMLGbL2UKkr4KeGsE7w1LwPkowExaRq
FwcdOGQFIG4F325iXTCu5uML62LS8IcVEgxhVKMgV/2PTKQvpwPp1tS1yXzg/GamutX2weJ5LA1F
LnUS2LsCpAj/QUq386MF9caAVGet0UDyKAfT8pj5Yu2A2pwPo1/HwkzIcdJQxDT5MoUdiXWS5PPk
x8imsdIjmTfNb++P2vEBnoYPgyOoIJIfDgiBSqAJfHn/7Ofwxf3mrvf+3Lktl459iuSwkRvU8msY
6zqQxhKO2pPR1h8gacqMYueucz3zvr93BjFfhoDiz64swSoI8sZzpcSnwVBOpkqPVt2jl0e1vSo5
St3F3mbpLsuHLum9Ie+MtFEw8phDcxG7zNu22WJPx+aSj2bTvwS+rMm9an8nY14VwYNfcQ47fDO4
bnreAIr4saTAE3PC1D+fYqLtpV+RFh4a0KzY0AjeK+6ViOeuwtOnVDaHB4Cf287b02WStnCw54YT
48IIpZ3WAiWG3PF7t/2iyp9GEP3l9OP00zcwLMnhf48PFaCS4GRyhCW8CjUAw/e3qshC+6c5i0wm
5b4nUUSk+XpNPKaI1dIha/CsqDYGqjuT2yda8up6JCqYnHqfLpusZOMxsOx1u0OurU+obJpbcFyw
RGZsLVj/SdEiAP6guHHulsOY++S2tlBEQRl9LGQRmkd0SbfK4N4zdHoV6byePdMmRELMGVgm8Xyf
Bt/z5p4NRTwIPIqqWsthr0y2lRLlHBa9KDK8tGHSZAyVqciiM0DK8PF5CwQxmX+P5KUygsEZV3jm
adjGLC1WjY+1CV9Mnq0glxC+KS6zJcxFsE0xi+AQqUO9LAGTLByUZy/huiv08HHIaCMc3H3b2r/V
8cIjKStCFly/eIAVznrmNWgn7hS+wveU3ujTrpE+AbWje3OLE/oauJ12w8dFJ38QODdCq/5eWsKR
b1WMGztKtHZq6YZjheqng8OVy/6Jmzn+DNAKKvvdk3MTpc5Du6t3aIWGg9VAGQ0Xi0nt8F0nsGFs
RvGUWBNgU+ToWeCEJUieUlGr9VGh9LbJqcpANx+kjg84JAfVFq3sElvxuoPgJ0a66Bw7OjXu3gWX
AyAkBTCTJVBmgrLv0Ffy8JfK43EFKGbqY0Kgig8JiaUjV6R8Op1hCXYcwaAbJLOH+Bk7JfXs6+bd
Qa3AcFq/jnG9z98a4ie42YPAjwKiE+hP+dZko0VjNzECys0jrz2kf9f9z0viz3PIHeuFxqc9nKkY
3gmwGNVu0+lyIdHXxdZgO8+CYyVVJfw7uCq1IjQYGoTkE/A1LSA+Wwu8yT/Ln9iBOhZQfKKSj+UR
lfuWVggyGsnC7shHQ/+S5SxTvYXKlUyW9OSbD/jb6H+v3haEqlF/Hzc4sRbWxtAxnDATDujoT43G
o4qNy13M5N9rgzdjOhhfJAfM0qRJA8ZC9a0HugA+oC91BL4bNfvFsk7sGWjBoP9qxex1KpoeeZ7d
hLRr/x4BPKfneIkVoz1TbSlZ5jES4rx0YT8LIemHDfmLinS1Lf5kpxOrpFS5/1GsaD080UrkWR7G
rLzksmxwIGMuqNj3nF1woDPgC4rPade05Fno/6PUQ1515FBW1fDiWQyNBqQoA4rxlK24xfqTd3jG
upySVwYq6pAMpd4WytqMpgng1/P/U1YpOLiyiBjBwWSmRvS0qqDtNz33hx0r2rgyhgvMBs1hZMe8
jWauH5Njr9D3ee4L9puB+F0eL7/F8PLUKGI1MNzVYMlkmSs5GPHnrOhE2jEUB3VaGDW1Kvtgb261
0JAwm7fgNtcwRkcyHfLNoYmJ+gz+dxibNaS++sLjFmztjt7ez1OSBFOr6Om9eyZjqcuYl87kmrg0
gjvF5fTh+SdzfJm21Jev23Xx6a4uQvzP8FrqeuXwdcm8tCs+yxOkIluXuKkmSf7OAl6OPLz7kBeG
U+QWKaXtBHEbGNMCHxK0yb5HvxNr/Q8SlM4fgvxjpjV0bJohuUqeXmstGslvXf0jibWzrt4s4hgn
0Sf2pXD3csydsr3alCIVhPk+t7jcuZoMh367vtfO7r7HGPHA4dH2IK9hiseCoHNdWH5HcdMKv9Mk
FhlIYzW05Nng8F9mvDtebjDFzz42Zde+1Jl+baP73HS4OpedNf0ahe401hTci2mA7dtk6w24lG6j
srmbjmLSk4SWB6fZDj1ttX6pQsD1wWHTlEwOnHlFiTzRbGU/7Fn0g4Bm6BDBLeLqawzmUyESNFOM
loyJQWnbdWrUJ9klrx22K/eAJLh0vLZxUm+3y3qj884gJ96CBQg6qAjf2RAs+K/J5RW61NSbL5/w
Uw0tw1CzuLeCmOJR2Ajz/BcbIqPeq9Zo2L52vargseEOuNGrTyHQKG4eweTLi4jZCMn8f8bvGZVz
la1STc7ojyQ2SIfKQe9yBP41S5J0hXevao4pW/za/WMC1GSv5RAHfk30Lhfk7F8p1JTQjuSkie02
/uXItOOqX6CeI4sQXUkDzp0UCM/nBq4uixOel17KUkUE7jsPMOYE5PrplxFGaXh2VgqKpTMeTXZ0
Rra79pb3dbdJIo4HcRSZ3aTU722gJ5w+v4zXHR7pJJVVeGzxnP1T1s0/hzh7oqMJaJCGpGIOm2SI
WeJOIUw1v5Vga/EBWnklBqLR2C8jFLgsOFODo7lsYeuoQ7EzhXJ1kVVGprqn0BIbt8kLsE838t+1
IsnrDphsp/ClwNm3+G9q7VTAzCR+6h2TlkbewTpC8gj2vJ80By00Re6tr6AScVWVvODPZPo+3myl
RvmTxp41jYcryeUhlwgcmpmklbiDn5Lw3bJ7Kde0HSlb75CHL6oDMRdwR3jpW435Oj32zngReuCI
uAj173VA1eEL2g1S1GA7Ih52g4xblZLnL+ouY1Ex+wIYZCYVsB/GSIn7si07N3c96Z7ciz6snh5u
Olp7V6Ix52dGr2eZtbzAeV/OIEL8s/fISal92p44Kqs0Eqle3MuoY9ZJ5cwIO+lfqh4/fCRBsi9w
CXoGdlkM91MvocXa9vwf6hCCuabGWRH/BAgQi6mVjACc3iL1xfYNoR9waohHVf2LlR75keshFsMt
UH7/zsEgwlUUOM/+xeIDaEAUH22JWMTWyDQiIhR5eRBTbceIoFvdO9zmzs1MnJt79aq4o46wcp4g
nG8pVIgyDR72VTVMxvSjhC76deb85GhN13tDoTf0EKc4Fv+kywdwo7CUpy1LF9Z1D/+ghKTHEiMC
TecUy7e42oWetnKaiO42KA8tULDw+y1ZdniEcSz+naK1OFp00cBVQ89JDiqVRQEyoYyPoE/I8Vjw
2VBN28NFLbTZF91JGamoOgP4adLaXhhbBBc+WLaczI2VGnsDWG2NOtQ5En1ISAbx0RaVbcnKDfFM
awXCjeF/kZfVhDKqtdb4ll/cyQa/FI6+M4JhIQj8u++q1Yq9ZdXGgJwH937SORkBaC4KLBcKSsEl
JYJsKlrth71X/a/wuJ8Sb7YKLadaiz9MpD205ddraoPyQ4dXOWanefyEtprv162Yh7qinX+ChTAO
I/Y6ViKy9jyUrC5F06C575r0yXihzCtG0NfmeOsXn7hFozfzTX3mHcubaYTn4ztKLiXvrkj2Jbny
+RQtT+ek8XM0pK8tEn6o4nUBXrKNPOTR7JNMnfMPcfyLPGj3rX9DFk2X2af0vqWSTLWXmNOdT6s5
afvMMOtyT8Jn2srbI3M8A8njBY2biMwIua9G2JW/GxZFdH/I/Raqypch3fYESquGZKC2N0sWOaNR
6hB2hsd4p7Krb+Bbi9goHOKtvYjYv0NcsaMq5XVxkj/91iIiqBPC5/fklUofSKY+J+fR8eNTgTTV
lMSJNBdRwPGXlfxxuHkeAU1BRGAjW7gPEUzLi8R/QjnYUh6A78pTeqNNQTLWFXp01qBX4ksqMk++
X+VYfzVAnxljmQbT9K5bOcc8MGdbWPO2SpXsF/fbx2tA5UgOIQapT26R4tY7RVcvJR2lKtRGZwpO
EPdYeCQs92cjoQ4+V+KtgKxKlCv50bWnKl515nGk/mhNxRKGzFfh2fWFS8vQFf378j+N8+MnAyPx
AMKS4g29Dc2ijUWsTitr4HjShITPS6lhbAPW2TrrqKDgf3KjSdGH0QepZKig4fhrp6yK2thj4BnB
P8AZBOjgfkh/+kk36Cu2tM38hd3V6aagPhjh/3LK+CMB8QAuuU+mVGaah+fpW70hN1rzjMK+FSwV
6Y3OzpXsW+JToxUT6jcL3L0FMl+HtS+ZpCIp6320LwOaGYnE78GbDvYCIXeCHzlGm5xkz/ZlQ2oG
Z1rqXhh80cdUPTaSJYqNk5JcOzCzep1AyfDyL0+zswl2iPEc+kBND5zj4N192qk7g/JUNPXkMKHY
uto4ZxANalutmM6iW99pDrULPzi+UN8yQ9r3NFklyTd2NeugVIV/G4bGWca1DYsNIExqJ/kwTEE6
ZDB6KPN+R/uYHpTvm+4HheeC+xsqBBKqFRtYarZZUwIRTCdc/RbPFr1p2lo8CRkFqmcM6RmM72j/
z7S//sSi6yt0y/mj6yR0uXAfyiPRqB1grxBuo79y7lr3RhbsV8KDY3MQUAyYDgHKkPJVJ2uWvS7z
5GmO7pEccGsIWx3GPaawFUM0WSz5MMO3mR26hD26voXzZfMFipfhJWUogfD7+dtqpabsDemkW7Cq
u48gwYGfWUNfV8vTnWfd8dFOUGobAD4QHgZdOj7/BY9MQ3xN6r4hTgD5CqvqLdfX2EB0ytilOJ59
emgFIInyVkEs88xeqPV50m5Kxwirhg69WqSmyArHZ3VKwwuIaldBFUjQb/OADeYbMcoNFrtEV65H
9IZ9VW7Q8WdsAV+MgJAuIImaZ4OB+h1l6FaaLv6ShdbXiAM1Xs+vRn6cbph7UxGb+tK2kSpH8tMG
TPEGuGrplLKE3A0lScypfxilxded5L2vAi6QTTMgioE/CCSmNW1Q8c9SbOwo/lBrRH/V1LNPx7P6
if0PqcaRoV5+hyDobivaYGEl40rawDQdFAZw23CfGycN5zpzmx3oHWRnIqmFMObSUeJBp0wi9UqC
Pbdr8wcxWiL4txY4Mpgeexxea2AM8uhiBAh7HvLlJPNFE+1aKDswvfP01RoUiF474ac8vxRiVgEJ
LFaGQKfXD5FH8KykkI5E9866b7CjSPDLguA07iWoc0G4GM2ShumRpF4AUKa98U6Nk4lI0OBhiO03
+msone9JQm2Amv320bM6uZ7IeOHB87SPXoXL2iOHFDvGmIClWjOj3WMjnCH3B9mi02Hviu+f015Y
zsVRojPNirSltZR4hjAQN0t0M0O5m6lgFHGovjeEZbmkQlis/99DmTU3v6/VToRBYXJcG9RitUt4
si0wgBhYManjnOx0S3sqwEmkx+2m2RVvQtePvkvWVUXkjdkIv6vzi/S0Qfl487bKdZzeonaeX7SM
JgwUUkqUG0qQFJtUEfl/AFiqo+6bN4mxKzHmxEPLqxUsj8mlh3P9A2DIJPxyqW+X3rlNM5WPg8jS
vNNI2DsIVAgkeGQBmGOn3t7SzrzGjU2nbI7h+PRU/BNuslZYd0SomegxqcJbMPo0IKSw4fkXoq0R
f47HylyBma6tMu1xueTqAif5NQEc6lKxb74sVmx4g1PHNHyEslwq1+8G9kLNGoroSb4SQrTMyHsr
fc2Oh6cfYZYj2OHXvf7/FUQyQVK6pZk7rvbFEOnnSEzybsgkoaFm2I/zpKEvKu6GKTuPHBgCZgvU
nEdZtYoXfociWrGe4Pru2JZJjXl+BY+n5s6d2GvSDhTKWflirkuEvCZvG7n4WLbiM48jtVDyQFGB
/y0M+oZjt65z8VMWD2WOdVyIjJrOodJF/YDjUHXUif+sur1nRAlbvRmXXU3bbdSv9qyzrFFxYZDT
USzZSja835eGalQ7Wd8rvehgsfk2Yf3cU1FsOXUJhYcjoJgGc7MwlzijK/gyNIAMav2C1aQQmGlt
C10IpuDuA7JxFPaWqPcrfk1J+UiVAAuGsaVt2JEgM2Vh+csuA8bDMlWFI8wlLwjIb8nF7azOkHMK
EZ8KhMmNKJ2L0dxpavVaIDV8qB+v09z+x0lENTkoq+2QY2CBCC3CeBC6hx2/KWVwEEJF2LDcD+C+
tnOSb4jPt7IPA3vIR/1vqqbuX4Sl6WwyFgdIA0gzebEAVRAb+ibcsBxO7ehRk6tfIBUdfJqy8fh5
CVbj7fEji/VYu6TG0rvNtORHuuivibbmz73wVBuQLj7ZtLniHBUqI5d6re8fSZDXvmyrQevPrOqc
ayuoghlZv2ebuNjN6vlovU4CkgldO+GfezjERLBKsKhwyvPrU8V3R0jlANCr709oKlMpm6CwUaAd
OejwrQXKzZTPP3nkGHDRVV5zJyWvhCtByaYi1fiazi7mR/ERaX1i3xc+ZGyub1brGBq4bP5N9PlT
hlAf+jQLuzaJQfzkb9ccfpE0YHLbyZEImIUtLhPSM17p/ZN0K9gglXISzASCpZMsBbbwHmIcr47I
dMOFaGY+0v0aiKT1FnFI8eZuBD/iiB4PUFBisoKRMk22NWWZPJemVpuPqQIrEKjG5u/5tGprg6p/
5pRxw09S7ULZcVcdL/Z+vuFXAyZY0IgXXBONmriow1zAsJQYyQJ9V34Wq3DBnqibzkZbYjKfVIEm
GSSz8m8+pThZ2ZKwZFxej87zt3OTfunEkNN3/R+L84zNBIXra+SPn9H2SOR5KUs/UqvogEyp/V9S
x/kovSb8c2T30XaGvKCudXFIzHuxSsyDn06omNpTjLccOSH3NN3ZSBzHnBswosuRVQVowyBiUII0
EYgAshN0BAvhk/FRkuSRztEhcl+XsoEdFlbpS0Rpu/zJYcGCIUlaouX2S3vptwl24276NVADJ+mx
2izYRxBTtd2yVZduQaS2IB2fRjGB03u8YJc1Y6PveclIHVG36Ws5T/9JJi/2zkVtJLNXvLOH91CE
CtiAIOLMM9rGMemwIb3CAbldhyY/qSKlYPRBkx6wrrhsIL/Cncf+y/3yPd1UzL/DU/brAr0sGsT8
ZVb5QOAFIv4e3al+P/9cikoAORfxcgYag2WSkaBku8hxfNAkvb53ZJB0wBlLBwy2JI+JyFxMG8Ij
LRAG84pN6HENM4JERGihDWDVbw2uYfic6eqmZUbWsWJlr3bz3izbCLJZrmm9JIhYpAN1/dEnZ52u
0xCxzimjA46VgKW/mJ58llX4vIDz7yhnAOPePbPzzA4r/CZihQycipbpfqGFUTjSwAqNpzdEzALw
5d6W6Ibv4s24HeKtRFVxByJ2cQCPXQKeCJ4sKpW56mysIkzcM+C1354zFwxm09gwQd2p9yjvrmGk
ScwWr2ctIdEYDE+z+p2PkSm7/XL5mUFCC2MLvfbxfZq/8JgoB7O2q7CU62FjMjL02Ds40g9+ZiPq
y82Ivzy3/3BIDUHpCqxiF2I+HtMfyZ5Ry0peH3mV0C2BYdaaLCqmT4LV9Qx2gmwxU2bSqAWb5wsU
ySkMaP8fxA7eYss4jyBdL1ZLwwGbi1LS0NjgzollSenB7oSfwbVLmIGNV8ZgXUdAowqGYcbdQgnr
8OT33u0TjIFID2uqYaQgPYYE26UVE4w4bBCvTS4932pF9gmS+TqEWL7lEb8ZcxCJNi0wrI5Ckm4z
dnddofAMOj9cWh2nrVzc7ekoJVy4dcafOyeFTgtrLLP6KO649BAZjjKjbbjqlk/Y/CLge/4Mg6ye
jXAcSefJZmqnjPnYp9xjclRBSImGes688xT7qOlNfPcMZfoYa21FIUN3Lk/8rlQm1p2ywlQmJeQB
9nyKexbjKEktM46H0Fb0CfC3e4l4Yaki1EzadMxbEbsGV5F7fUaU2VRKKLTOfJSpEsVeOZso63LW
5O+BGhOkKoKJokV5Y2pGm+PqdKiR0CxkIk4JuN86AFRtsrDdvKphOhx3Mwl3RH5vsuurXVys9lL7
RgtZAQfjteQ62+wJ65bOcJY2JgiSN+aqcJmTBAV7PAuVV+d0KoAeeCFoBHPBy3iHqxw2nJWJO8uD
oND/g4EJ5qpnTPjQnXI8beEmvbvvjAnExA2CPx9lP7BmSlpRSwd/mr86ORks4OeOmsOYJc0QaoNy
ogdc+kQ0ArRAThqUdHsiibDl1OFIkkA/L7XYY2FrD1x//6q0OFBlWSLiDAYLqK5NZTto/HX+TB1q
CjCi/RB6flnDnFdpghPQmQbpbfHSyOZKiE8D1VJZw+F/6XixmWw1oSR2qdH/rNgXYiemng/79VSi
BqdaghQQj5Z2q37UqHrXetYjNXzCQ8eugO53B+9dbRVzOhJPKtF7DXtLSJl5XnTd5fyvS+YI9bSX
MUKHlAKQMQTXfx7LD2kQ/eZWRc4EugFuRCQ8M26tKMDhtPVck0pUvvEvUdzIQMjTIEe+sqonO5Hq
19tsYLvgBXvCzqVTJJGVEddqAKys7UpYKIMx560uX9FxdMZT5LiibQUT4EUYsk1SZjizEnoP/b3I
L+MtnPq0jrIA1i1i+M9dbV/20TFNV5VofPinESzeYzKTuo+NERkINQHic1VCIlrNxIlXjmPEr8+Q
1nQ7GxK86kFODcCRU8VuuzJJwwCBSzVmypsaTy1WnA+ilPNJLATcWQR6NG1JNgE+Jaq80+xqs5Ey
TAVerLNchj4DXt6tbcMQ5PJKTh919yxxT/eVOp2oN2KC2Sjq+BI0bpB/kcjAgDzSXDnBElYPzN25
eSjMPJorGMmgoVWDjII0bp0NtSayq/5+uqSL6JKZwryvMKnuGCaqnU5ELEgEk/lujz6pyAAOZX5R
HbrlHaIpw1CqPTyuv5t6UD5a35QFW3pfL+aRjUg/2vpduXnbQs/yZ9Rgi04tFd+qCmavhSGxuT/4
T6p8vhhcrCh256/lilZDCNn6WP0LyHD0w1FFimI/RkrRKkvom4/EK8xm9d3gdQs26ZDKfMJq3PNU
ooZv/Jc8B2hLCTJerw/ms9b6WYkoLdvydXdCl2oiv3aE/tExw4I7X0hEALMvBCvxKeUfdeFgdOh/
T0voNp2kq5Fm2kl3snpT9r3aZrJm2slqp8Z1kjymCoMSO596RMBgOTZs5yBJ/FwbL76Nhfx6OwMU
sulnnvlA/TSSau5VPef/kK8BM5WqNxPnE2OhJW/6AQz9sA+875k9ReikrITzqM4yHUPiYzff8c9E
7YilIhYFDbmPce6HYwG0vwGqKbFlJDI5YiwBRa+FApfJAAjE5+gVmEr/W9O6Cj7gbBEh908b8Q+g
SYoRHV8A2Foqppig0H06OzxQZ1+8rHNZDbSF+BQDLZHWfwk7jVMOLPIJlwKCqoDp23AUFcf4iEFu
ezvkop+cYgGZdJCba+0dB/eOhZ3Mpg9tb3HroYuVeOjxi8EQBDNKqUwIgqbxz2OFZoyx/WljUNWN
Qe5BBHu87mtHoYBQGftOtZCDcaZpwHissI92Ra41k+aqIwDri2UYDa7NhNhAB097vtAF7d/k4wcD
K6Ga1PfmHXDFb15/MoRUopppFC4ReJrjsT0+KqHSfsMYivDnkHh+FOzU2LhX5NdG/vjvMyDe3ZdB
I2hQySrqZFYS9bWDUmI7zJyiXERV9PvwFGZBh5mXiTnY1bAiMNobUpOyfg7eFTax28QvHz6jO2Gw
hR9X2sHAtQiEucr0rplrzPwzzAX2QJ9XTDTyS3Gv1mpakePJEORwgTXRaN6kG18IG5D3pfN96tDi
VSvNgbpjEJVb14gxyhD7nqnOm8KpaKscBwyMVxzl5m8d3TaRp3SMA+oPXAJXwv2MSh6PIeZjb3Qi
sCP6mbdI9pMJLwM2GVwKypIdWf9yMMZwDu9Vph/E0mB84QPpqbKughf9p9btGimCuvkd2r/rbOWk
TO1dKuRPOnQk2s32w/h4weMT1nWgffrdbM1jQ9NiI8CgWobBaUGxHcFSQv8g+0mPs9Np3wBLI/+Z
Jsi/idL2qObgb4/moAAIdSUs5ZiulR9da/YH1ZY46QsqCMi2/NIOyvI9JSW5phjw9hQJV9Hr76X1
0l2knUcfetyujFEXNgNZNJQpTa6bL8cEyaXqEOBbLj40W8f+NsTc3Zed/6AZXZLETnwYXmN51BZs
3mr+RB8yCW4+nk1+q02ZarzPwRzzC/Bmb83gw8ncLyGIgBKJfOx63QvjIqndBRzvvZl8cojsowtW
+ccfSXfCLvzTC/JKamkxbmdlkESI7HpNnVVABWpu5hxL/DYlYJyjGVZNWwIVHyKtfNVmwWR+dHRY
bnuobvqzrSRdxhcHYYDfiEXjyFI3Ihbu9xLPtSMUKc38C9OjkjoAsNTQ4pHbqbz3okTAzmoInABL
1tViB3FMK8YpzM7yQB+qpq49h38mF6157vcV2oDl6CE+ncoPdDKMkTxDnOsDTkfH4vh8gGoP+Zn+
t2R0z+2KgLPW7fr4j4zXrspnIeIhLpFZ8KtikCnQAy8Q6HlTnZ+PSlUBGrD89qBX5zsJ9SRxmhWe
X4xZ4Z+rrT8G0xkjxcZrevuuETRm5t7iR6v8miP21OouYYCafKFBbmFXNJPPwoEg64iQyUgb5AHS
Ws2kfq0F1Jx4A5UYMGm+ENRsKFGm22w9TvnwcKuLBF1fcVM6QWHd+T5npudS+xpYH/oynMJ3bLjE
MqfvTW9SmaSB0p+UeUO/qyHn07dhFvZWZPUWBd2mmEhB9Id+VH/RVLbAZnGNzmwsVHQgUJ6TvJpH
1oBB/WKK9YaLXPq5Di8vXmJ3aUSs2l0dZEFS/jnmd3KmZ91XCylIreNwXZdqNO3gi0MBmbGuH6/W
QcuRcvhGir+zfxF6uspiu0aWoLjF+TjNnwDhV1LN/nN6Byp2hmOuLM6wTSBhD3O2YjZ4LP6iRRPi
yzBqYRe1q9KKXcJSyZUUNU9HyqBiDg8HbE/ywJFZxqZmWy5/qHnqjhHq5+wYcucw4XaPvY1xT5OV
5qqTNaJVBU7OAsBMrUeaJPXbGR+KbV/Wwd6f0pfHesLwR24gBJ/JbH3CWC7kveDhpilbPp3y8Gfy
EzNnB4ASPCHdd8Bhq/9f3y5THTJYBjR66I/PGewCLZn0YzFSSqlRMe+/IJ26aNtpDO3dcAPXMibJ
oGouF2h1TB1P+broE4jIzu+bCwMpHUkbZvSvhkTq03YToAeYtiR+Wdz63KDFijq23UxQok9Wt1de
oqMgx1BTBefyiQ3MZG+PPVb/4wqc4Xiz1Clh8YoTDIYjeSIAl3j2LVNqbKkukIOpRAQAdvYMI5nH
Iz+Nudkau0Yn008U/ER6dl8V/Po8fYLjw3AlX/JR1r2QBPiP3j2agABSi/oSlv/bFWvNCls5yL3Z
J0zwvz2gC5yE1NqZQ0aNORT+M8gbxPd8o57WJdTx0fyxYpalVvcGsguej31Z2knQd0hlBiUiabYe
5lpghSoY6xdK3TNcRPb/LsSL0rOC5gr+Yg+p1GQndt5qiRsLHFDgzLK4EPNrofXEANIfexkqGJQW
BYebsMm5vTgNRJ5MB4TaHfWkoC1fouJwVpUkO98IRR41y5jUxxxH4dPWq7LXFgBceLGtulbzuD6K
27ImomKnQGvvFxztnE8e+ZgB2wVurKRB1tpGxfm2LIrEZYVJUnFISTuzAf+HbbpHi4B6tTcCTzM+
DofaI34uLkxvHor5p99iQlxSmhGADkse6tqCl6bMncSfUGcwbAIIHAt6Tl4sNSmY5lkTXAPl3vuk
xspMHj2LDPzkNCOWNSdfOX/75JaEFTm+Gw/4zTuFgkJDyzGX+RsKYwDZbETJKqX0lVUo196Qtcoj
jNhg4Q7KnVRGmuAJhqqoSlvtWInyJjWDccTbcTGuGls8QkNeKwoudg+O6DUL2uXp8PvmcpA6CrR+
9hG/14rSFEEH7HHXMpikkb4SNzCwpW4fhBXqjUu3IWGGxaKx7Eg+RQ/NCNSbm55Q4aLuBS43lwRL
kOHV52KU9E+bFGtbxrb4vm4GkDEr6gARXkes3Zi6TKpSxPOp+NS197KXEvZcjqPFzQVuKIrWUVF8
FLMuw2Hyidskr/uByV1tjXLjxYn0JEQ3xGWHkr3yOgF0l9UlVN/OkAuwNFnmN7M5RhWEy7LwQv1t
dXlHPuJiUgBuMxECZupInxWB7SB3XBNEiDa/PgamYXsgWj+BKQWFpxjNrKQfbLlJ4HHXG/f+yEqO
9udBtV3RpfxkrJcaO4bD6mHE7mFdF2gAafiB6V+HxuJAVYgZ3503q68HrfucGKS4R42U6K5evG07
SxV0Frtm2EnS7accJEw7Jj1/TyOgy3Eivrc0ANCWjNYbLxoX68/qqcN1ZP6/PQ11KGDbzUMsGnZH
apXIQSVTcXexIBaV54tf4D1lBGs2oU1xnFbOdd/M2LEAO+R5ufbJ/6A+og/VoerVZ9YhV4z1ZIvJ
Rsao3mBaCsWhUo0MpndrNf0Uvodosp+pG0kxS2nkrv3u8xE3hb2w5y74qR9Z/8KOymYxrHwalgxg
GVL13HBjQw7jizfDSQmsSh2GC1ivRqAx4LfTwDEn7hfy/hlv7KXhHFTskB91Cx2cVtcOOHpNGUbS
nMZl7TfTbNagvKiki8ik/1QEhTTWpv7TgAbCVVsWfJ/r16fkbdU5vz02wsjH64Lfm1pb/oFWGD24
gJxWSLk3lwZRX/MZIQJHzSmV2CoZ4BWzgyp3vcFvwhbHs+uRcX49LrELAoCkSRuXnZ0HCVnO4TVh
Ur1AWoGcNOqxMh/vWSNJGwW7NoeeEcHv/spojqfyiA4upeJkpcnfo2gwQ1oO10FrerrXxDeoHyu4
71wVn8n0c+qHJXygLCj+RpUAhgg6bzZap7Ti2HRDDD0IJ0RMKqSLjGDDF1D6I4GsyK2r1c0hY0YR
+FM+3qWPsuVL9/FefhBcapQrpYbvtPqbrwi+rfsijJjX8Xhmpwsa87C1IEaLqs8tQdgSCmZMtPlO
igD3Bjs/lSx6C5JOOB2fjHPSvTj+R5/RpuHdwhvLkC9aZ9AiQUGyLUvIoBvBhZSMwksAaGhz87N0
tULSOXVZkHuQnwFPoZTNlY7O5JF9i2tZ1SOkcQfszgVl5UBOaENYuTFc0/eLzl/RYa2sywT8in6F
x5bHgtW3aQipDuwTkzkj6QxKYbXEQY5Xe5723hi/fTpc9VaqZhgQtl+qVGnaXq3ylCu7Q4mNmksQ
USAR2AKRyEHTxSwDrxblKxuvCRseUIwxGqyydcfPSUIEeHfG5jiHdXS2r7aQlqXn29XubKf++dMa
WqnvFXH//kbpLLgBgtbI3eoaeoVKZuCmzuxH+wgcm3EK+SUDv5jmLo5caCuZ+Fe24uN3vKBBONQk
fczn5GWfCljcln4ar6+ZOvNFNr00Ft3lUj//4HXyd498/9XU2S63l/lr3pMNYxIrNt2USt1bnV6x
xdaekbyvG2ZQN4NcDYcvMSfIyld9Q6w6TXKNwyoP2Yh+aWulSXG2/aPUsEj1BfhwngIGRQ6ChY5R
6VByGOvNONPDq8MEelX0WbQqFWB7Ad8VRxyDG9w9ITzFhUwL0wf9Db12alTltZqoQyX+vTl9yuSt
X3bWgblU48qb2+7vZyUDL29A1qkV0HV+YJHXt53Xp46P1cKBbI1kxxDf3+IXZv7AknFHxv0G/AoC
kA0N0WgTAAb6HK8P9NE+08or0VaQ2P1TFVhPN+7zSH7q2oSlSe/Cdo99Orf5CB9xYwWWUrBoC9R4
OkkS4LxprBfxTxgDucl49v3AQYLO5jvjVOXMN127ecIoIEk8G8enUHQFEG4Dqz4aQ1/ssq0xQ/V3
rsTfFPhx013dufO5d3IUfN15F/6qhucGCMkYDpCE0WYGe1h+c7PphH+UGrkO+UGqv3/mI24tXbbu
o8/2letQsbJacEDzzgkLlJnIvPVJ2moXfS7k7cuZdljnY69iHQp+v4XaYb47vdIp8CIDfkrgTg7X
Ic/wTKp1nrQa08jwhBPqhIpESpg2+8FZeYvnARDiCf+fsCcJaaqs5mmfezW3FcZrwUrkL+JJHMi2
qp6htsh1hPZq2LZ2riSFQn4r8I45WOcy5C8BiFtTG+Mm4Z25ii6wrwDfs43yNfO/8L3oi6yMfZoK
QTqPksPXvZOgV+3M7bnK7pDAyyFA9uSMjxkOOzavtgPReXXe+J4btrabAGsde87sXMQrFud4RVUo
hMHdC93xpcvIIJ0SmaJg+SHMQzuzuGgGgluwsItHBrWV2Wm/LyUAL0fdKH0C6jebbBxUKpw3KOq3
QLjBaeooEGOCBoQoMlPRTLqB8qaQV41LLfK3iNNu1ubhOmRjVOqGkbv1y5PPVHuA52zxcowN2Y4t
4H2nz5CBXEKMR09EKVlBooCNfvglEufqrLa4sl/KouMwfO3wuWg4vh1FNcKVa1x4ISItQoJvmuUl
X1naUnA0NqS4PimFrNun2svWavQqIYr13KATO1U+/qm9urght14fuoo0YAUw5zhkaN8+fHwW8dst
iBrTM7fu/K0CneN79BO6EEQIPqKNbB2QMQ2M+mgccPO4j9qUIVa6PfATUtxg/LsBBl8Vi2r5p/eB
DGMjUZ5ahD3fAm1Q2yVVXxeYCgyHj/nXvbc0B2I+ngPplsDkq2drg2swh49VeodcX7FLj3G2F/Kq
ecVYijwh6SOpBMSDRkU1MHvu5F0MgrIzoddl1wzInGGjMs43bSByhnRAR5JIwQ4nVNVWrvRHaJJj
68RJrOGxR2sYJkALomc+SiOipbkItlyReId6DyOhoNwCVNYr1N51rzBBk6es9WPmAvWG5x1uZVJI
igeAojrcFdHHCzmlOUR6vtqUvZdDjSt+xHnanx09t+h1tiG6qTmWxbC3NkqBzy6fvsW6Q2rJPOT5
GcSke/9TE9ONfAi/zC7IrMzCQPDr2UVn2p8k8y8PETlpszzg29sIDhkit2eMvU9/oRBsY1S5vURE
kJOZeZYM5EAp3+LI/iRuMc5LIYQTyC3aY1Iz7EstV401nNLR5t15iwet+54qfaM6TYKgbK/fWV4R
sq8/ALUj0OoR5Crgd9rSHAnQz7vpD3UPwgyjKo+jfyNvY72HhXfLeOGyUsgDTgSkc/IQ1hlj3rwX
sQpv55V9nVDolgr4UmuoNoxRyduUvjmAu+RZg7K7iA15FsNww5xbwnXQwYPLEaPc9STwo9sht2K0
XtVNWojT7Ubts/ch2LXJwE/UIW0BWU7uBIm5jpl4yImcqSfDcnmTK2DnEb/otiWwhIugO86y0liq
Dmpl4lAVdVaD0bdjZpU80H03W9RR4+3K2EXh/zsXn2BWVBgy+gIBGB9g/Kj1Xn8ICx6gYy37UVoz
OZewP2MFlyYT9IFafublqON4z7d7Fzj5CVAA6/Yt6tnvqg1zH38Vx4oDyW1AbBgUoKqeT9Z6eolf
lVdJHTffuu8D07Yh/g649kAB/9t3nPXZOgvv6X7kz0F7VyA/iGj/Fx5jjH6Y3TX+mdRX0qjA+UiG
xFzk4eXaQHfcAiqFW603Xu7KiZhtVpGOt12RMj9S9M6yUwUBG2ZT2c4qM0SFu6gkTrBS0EXYNnmo
Cn6ULH8APtOGTODqebwGqHOYSAUEbLyY9xxzXON2IsQlayOSMs5J27YufrF2zlNSHjp4/Tc5S5eN
A6cwDbRvmOMRSco27JvMUtNWeFoPCGuYwW0YbMPbKZ3//6gz+YM+MMR8ANNkYg5FozZQ1GNQyfrR
KAEQNoZUZTLukemD0MyqyKqPBdUdrHUdPK954IwOLIlfsMG5Zv+rJiEfL599EU8PdDABsAxyEhID
EQr6VEnsvlHe2wISnaOe27FEJs13S/F9lV1htLKjYmehniYnM0m2s2PGUmB+MGQKtmSX9F/3CfDS
vKpJKUpFZHyMZESOtmey5R1wIHtGBB1ziAm0+yXwA4cGuUoRsv4XLD2mJ8cXHdXMvsx7UtNfULzB
2OkxJCY42DdrojNIdwfoxdLAZvsqpyFPexk+pf1IC01f3QKEYcshdXrW0c2q/t1Ixi/wdzo3Ri5O
AM3hiJaaubOCExt9mvNQJbvouvExk6AzRafd684u48eXlrjECqeCSZLCQ0jTS4MLmD0yACmE67Zp
LBEFqeXp2PFNwK0YOk5/fouUqu09ptqh9JvTA1tIGCdyzSC0l/G8HOv8Zggu6U43Qaf360+Y8h0L
pT6qPk2wz/pWrFiKl1YiR83OaYZSKWddVMBj5dEo32AJsnWdBG0f+QGbuoYGfxVkayZkL6Lu8qtZ
cUTSvU+o9vfaz9xXb3yO5wKysTrd4dg3TJ/jt21Ki2Zh/KHpt754hlzcWpPmbxCScstDgcei56aQ
n7Ant9I9tpU2ZKa1yT+jgMMNWrPMGKwwlDMZsJHKkjE4KnUaRSdF7xG5M+dJ4wHwHlFMU57/2umC
HSd6cfKAISid58aZXEbUAGgbfi0ukWHdZSlsk05XiveP92KzX3PBgiCzIrI5x80nzesgpSP/EcTr
jBTotKBHzT75M0ibfWPKhDck2luDFMEa923/lV8w5f+OWUdVA5FygC4TcJaqr/lT2LK80eo0d+rT
4traiGDCQ201KzQCumWeCKZ4lMFWRR9h0G/gvYps941kVpJmR8KmfR30Bk3LagkkupNpQpJhMLUY
hAHXOohiu3mChsPvbeFHP+g6Oibk5aUq3zY5od0j2fZGVm1q9DpWae/BfjD7Q36vhXixs6x6/bsc
3Zzfp1BFH24SMR7Mhs4jSeorjViBMGQ9ef+eAM8hIwV9cOdj2YQm/J/PI4wjjZpDAAhEGY2yN+RI
p1twRITcoJveRmSnFNYvzTlGvV9y/j+Q54ATqlo7+LTAHH4bkexZPEDLXBNf9Cypl3FeN+M41eFM
SGd3TejjolL3ZC5pVihshhxV5Vnn/5jf2X+mYDCg2MAob6K2vUYbXCurLrXW0dwWSoviGErjIRXH
KmmVNkCh1wW+u5vKxo8KifauIYoUOUZXkZrZ4jQqYGXq1bGnIRYX52QJ/7C3SWG72RrTwDy+N1eQ
wVgT3fM27eAbGJOMgi++iZyq1ZoDGUJNWNX5PXQoV2pUfFrf3WFjoDNdvrcmfvFgGmTLsaILe8Ra
X0VbkSAfeepuF+ExR9VkPfJ5IvPoRXXulDAgyDOBKdUMjgST/cqJ1rUAlWU/2wKeKNgTXgYcfWTe
W9vn3VSdQ+wZ8QpHnabfrfZbS0FHh1SqpBPxb+1NC0MoLXzI9oZLSHy0sZ+YSREKqV0QXIJW4Pe0
8RpgMz5sSwtBjpWEQrmt84Rk6Yu/MtvslzVMR/DHjDCPyj/dlVyj3WZLFtJpvue+INk/KdJ/lzLr
1OmTeui7Vc3CZW9YVHfILapYAcwh8ewmYUllD9iwg4Znb7Pb7on+TrmswHSoO5LB9908TMu9KLVt
y9AhK2z9WTGPFbBMg2t/BqKAL6QUxtO22+PtjPGPFIrSL03Smv7P7BnCL6rfftRA2jY3aIBRO/bU
M5+gKpHXjSWlkoW0rWgdSQmP5gygiR0fT3fG5MW8BY0wDCczH48U1arpyIBxjV8MpmrzY2gxOzCs
1jxj1z4bdxscNOynE7+MWRonJiKSYc4e8PGbIkZM+HQr2JA1JiX0nsv6BpEq6gLE00YldwoVwGTK
NIkL5okwOmbRrLuEfB4jVWEE4VfiATdJqttwVW7Z2BnzNbRv+EDb3FVOM8MD089teWsp6Gno0/34
G/CBMi24fy/bXRobq6IrRoEdTk15a2vT3rvrzIR4nGGyxi5HTEPKaCKMx5QF/Bp5MLQnoYCgsXvD
dICJ1GDX11s/4UXmwdLhrd6CzQ5trOiX29iVh3pN8uV/OoC6GwS+1DPTBlAI2WXsob7f6hTJcAnW
FgJYVg3XNmqv0gYwtIm5GGFUZu4LS5iE717F6PKRumaM7XEiqTH5s7J/9heM8Eed1bd8VapY+y69
rxq56/plFizqW92Qym09c7Wu8LhqRorzWwDvGED6AJJNsDkgw4wOV6McWMacoMCd9O+WAJ5hgWAZ
8sQIZeZ8dYGZIcv2TACO3XWnGXAEGBXeC6QBRg42FLVR/3ZMx1J5OrOCq4KMe2iIcMZJWK+o/Q4l
RjTZaH852foAQLY3JNU4Ixa3i/1HrV+jlyLkUOCcvPLaSh8uhyGnqlx9SvqT/3U5nxElUzQru13w
CpC46t99spiyKqUYwu7mXVj9rASaSlH/zzmykOtXDNjwkhgm5H0qQVl6lafKK4BsaNIuCZKjxMI2
rP3hsKPp+fhZC0LVL7J1ZIIhoBxUSrarmKZJBJ6haJA2RmK6WAAM4ZaSXTv0bpStX2qIgDILKcxt
difDHPhQlXn7QITKMyLmVBq3V+cmysbueHldWWuOiOPruW2kZrubVQlGxs5eUsDJg36SKkkOV3OF
RD3oyJpMT+2Fj2ex1REcL3a6VfZCzH2d872tqW8CJr0RldLlJTf7fo6UeL/Q7G7gYGHboiM4zomT
J8H615Te1ugXe3kAd/eD37szRMU8B7fKB3Edh2P3XhkXwHQx/Nrk/DXmyswOQtr7v/nSKaRE8CTT
cnH2nEKmDLG3sQrtxyc3slBvf2IGxHAO6gFzgO80ZgFbaiMLVzGk143Vxx97B/UlxhjHJMooKJnI
siti4R9Af4nMDZ6GzkAK6TgmyqBB1MWP/5I/X2AWz9L0PZTXOqZqsQEunXJjKRlvNjmEm1DOBbin
PgIMnAvjBxGR1DXsdp5v75LMtryMcRWseUTWFRystsJ5/Lei0RSH371a6unjAh7iBw0vzaJO9DVQ
S5/B4ioI286+7xUcBU5nz8Z1CzKWNM1jAIAUAMA/If0rdVGxbS58gG9Ibo+SDseh2oTKauOkNfHI
bC3VROw50DLbgixXzGRyjtsmLdXRsMKhQPGAVEE50KospSDmBCq5Lnb6+fqsfcLzlvxWr6yfkOy5
SMPcG3owhtXX6OjWgJowOOnAxiYE8AtYysNCkPFhus5ECXe7EcNfxF6U3frP5Kc6BuAHqMlpXzID
AaB7fxDKSey9lvYngmYIxP9Nx5bwsSobiCXXPW5sUkzYpdKQJIVsY3SjfA5NRXogpf3ZJ6Irkve3
BJYGstzlaY3JJLK/tC0EO/7thZLXgjFNa73sCnYNj5mdGLhgiBFsPceUroLIdo5BZuOluazeWqs+
EQkH+HGGBtM4HCMdwgefD+QRE4A+QVPxmwUY3jzviTUlXBT0rv/T2+rZeVQ7nn1T51EBZtiPUzuc
uZRR6UZoRa1WcbRVNbpk2C+QhJk16r/lSB8Z47ul4JTASPMI9J0iYPRyAjFDT3l6yq2JJ2zQ4p30
/z5IzN2qPpQHPAsGBSV8aFWeECwvp6aG4jgzqddGNaf6Ec9lNMTmwzKIrVdFgSQPLbrCtmI11uQ6
ZioTYKsrxkaVXg9ct0VEjkIZSZ4jd51r9DgsdDeqFzRAdP3Lztwv5reS19LH9RE9kyFeFFQeF1wy
wyrv+lzjliRldy144yiRrfQ6jEC6sM8ISxrWiqpCuDTBwW11Ve+JsOMuAuYkq84b2dnmiKMoN/iq
5eV3FAKzddFbltXD34F/gBXWlNA55H11gWbBbMgYb75MuWUvJ7kYW2cw+QZumNiUsnvwk32gIhh8
Ql9QUKuizNlvoNbWeUabgGA3FkZwwFDHdMGOqU+cVU+vqdDqp+klmJqnRrTY0EiF3mRJuIcpLetm
H1Tg7SSEVd5K6YOqivjQZPpIY86P44YYTPo+89Id1FPLReiNgyoIXz3nSG5E6bY+/M1z3+TdqXNG
lgGCKiYosOd9L8PqFtPD8ixu+4g15tDJSBfTMucTvPswNccRY/bgF3upoN4JgmZOegSuB075ZEPr
dncSkgCep6liLecEYXx2aM725IhoUT4GMIvnUFOzmHHvhndvgo9hgN/GBZYGk69zjAtYycO93Szw
+Tg/icc09Fj/v4vdFwPIxvIBfJb13LnnnnIb7BIGseLlv5b5383C+xvrWqC6so0Quy58gaBgTayC
DdLUbLfTC8VWDjA+WuPZrZk15ms4aYtCEUuG6sNOAqhg+ScXYixY9+X5GhA1J5n7tffEZS5MIIAL
saiZFzPs/sbIZNK3uXHsHyNS31yQSVFy2ATxmBvem9rYbC0oN06lXrziwXbQIWdjZqpnO3It7hlK
NwQpvS9L9/CL1N7QsWqfY0GMRXHWzS9/f79URkOkTPRegU0XB1r83Yme7+Ge3heRYxMklZsOUNft
AH0qUz9jk1rpDaMU8jyAzeAbExyzT4UKhqFSd6ex6c51WY7D0nGdefr/wFK9Y8TTbw0HsN5fC2j9
jg0q18qyne5DwFWLBuvjJD8O6ydm66e0Zqp69tycJR44zfuU6yjr4JNWADp4JAVwXhx5UoJrQ1fW
VRvsgesyt476BWnxj7DC7rKwJ9PBDAmfsiw8xoBs23L8Bc9KuRR+BYfQe2vEkIJcD5RI8dMkdDD9
xwdX2WVOYAK9V7rlu6NwZ9UwWyppzLzBTpkD7+9Yh1P2qttWuR83AvJQMVRA/oxscuY89/dTVqqH
tWShChiGJsfBI+sZyzzty7/RgiWGDh6qZer3yT7dCYRy0TuBP0n35a1rn3ZkFTRaq9T1Tbr1qvkk
Rq61fM19JYu27Iv5GPpXx+yppbpWsOTxpGjc10pnWdWLYZ5dJxybUMgI/3unr/eK5Rt9sugG6fTx
7sJK+OKL0rkWAdqFMvW00v1GjK3+J9QvxmUq9JdPCUAD+8GgC+N/3XqDL8wuyRWNX6jxNEpRqWRJ
k7/08fUMw/BlEAs2JIhvwPSEA9wJxo+yBaHvKYZfTFyY36xVlTDFIK+oS9IOuJrdll5HgWw43gQX
SScWHBahplaGYyddUqDDzNbheAXnG5m9K66R9MTvx7/kLjqgL+MmKm8UvTjFMFpOEoDA3BJhMlqx
apl6c9NjqrEcPIjfZ8X8Ev90pOy3Ob0Z1FYBbYLNtySolrYQTGpjCGo7iyQt0ThdLPVXk0YvFPwG
SvLINLE90psI/amSZkm7j89IiqeTjGmF7UMVH51IX52FzwVfv8ZMRYVtQulQ7+uvlKd7LcEWMdwZ
NRHXp6j5nr3TJXllpNFsLTmBOKS3xLMuDLHXveuds2AAmE6us1m31QSlntbwSfUvibIrH+ucmps/
hiuGJOkcGdxTybet+1sD5ziKIxniANywYEORIPA97o/n1yf3cdQspF35bKL5XyaNgTwLMQx2BgWj
VVr0XQxcfIBpfmCKCjRGom9vG3G0XzXIOdZZ5BJbpzUWol/PtPDqa63XnTCBgJRmDA847yKNpIjx
Jsi+TKOoDzQgdA2XAqIUDFxGaMZIoc3uHzXZTYWGixj6d1cUWSxEgsoMhAsEDWpPTVm2mT/Y1fwi
WvGIeFf4y29wOaLISpuWl2Vxfa6mdnvFTJFvOxRNOHbdgA0B9isunZgcVlffwe6vQGPFFtMV4BMy
ZP/g0wwoNLMN2+UEUuMJGv6ayx7kJIWV12NOlYXOnu3iPUbsBreE87xIwCZL65oVQj23CMLlPvXG
nNAZhg9dZCncxNP+ewbHJfx3fS9FIX2D5wCqPY2nDcXi6eDEcqTDKuGvAcA+VGy3i8ZwWvu81yeA
yOmVvT2kQmYIpucGSzBG2Srd0JRz+JEUSyMReH6qqfddA2VshjcExN0jG2/FELIQ1R4pZOsJjeRT
ej87xJtWJ2pxd+q240NsXOvRGNhVOagGL7rVKW/2Zbo6rYjYJylX6i9H8haTRqZ1ZegkPz6ukiWh
bSNIpMi8kyor1sBq6ZCASGqTz/eneENSnxASC7FJxu0bCfZvKRFpcupfYsOXhOPrpZVvwynht2tn
SnUXjgWIVJ4TA1DvFZ/k4puxR9xv179RvBbGxfQFLg3cXvDvtmpjjni8ftZQxPSX7dwIvmmCETqj
e1atNdiz0v1FZc5o9rO71c7YRwvNQWKoihXT5WpofIV/ZlkUWiuwD7QU2lHK8L1W7CnGVyWJnt0N
/stZO6NOZNrvriplyaeMEJoY5gyqBsOT3RVXN54hAiye2yUbYHNon483JgrNBbYvb8qwCI/fXpJ0
u6fwbJb2FGF/V49DZbDBiJHE8AOcytdRkpcIca2EmC06u5pJDmmLgWPgiix++V8X4bwnkacJAbYZ
dNfIl50JTk3ektXU819Zz7R56HvkSGscRS/ObolZda2/C8cjHcTdXKt3EPCzAV8k7V84k3jWOF4h
rHXSWud5GuH4XwTaahmpmtAHXNSDYcz9nhM+2hSRp6BAlFKNWjDRH6GBAAx40yJmc6t8ZFtXH7o9
DQxKJMvojgsw1gSnO3SGEipVM1F69mdCirFwh3/7VuL6HdrOUQiFGtJ0MF0xlwicMoxb7k9pJI0L
Px5W/w3Lc0PfDzxOxelYBhkTVbDYcQlNTzhaSQdHFMcwbOY4q8Ow2DAThLAXrseLvRbyjT88fdtO
Ea9vjPDrgMtYhpS9oUyK12cNbJkCi6ytbxOqWs1Px9H3khjSbKfarb6vmrKuFuTVlUUswkrRnLoi
qL1BW+sku1pSV7iQrqymqG3ZAU9VvqwpzlX0NgU7GU2gNdCWLBA6u+uoudZppTMFK6RMb05piqif
O0WMm6N0/52jeyewYJ5mlvSAVva0Pgh78XsmtaTmWj2K+Abs/p0XAF/QXSJSDYgCx51nFoRJx9sV
f3kjmgRDIw56c6N7QqdPP1bymWUaCQb6GYV4h6QbP5zAU6QII3udS/8ECJ9QWLxLnOtjKt88wwIa
ix9uY8FTGKqLqqVFmoLxZm630rDOrTmhp52WM7LxzZ/9Tb38NMHmwxtAmJtQcSkesqGRyuK5TNYZ
DhwLyPg/Jqq6Nv+ltPln2Cemj5idhjmeLKv5V28lJSJgQmMJNoWFAVDwTEeBmJlYfATo0K0G4LgG
eAeE3R1qzRbQBEO3KNn9EqSTuDids2GCe6ds2PmVcEgvKC4T0GSMNCr9xxAzT54DBofTQ/OpDV6z
55LyEoJ8RHRYxOmtyyk6m9F9TdMw9AflWx/Om2BrXPDEW2Ul7Wu76UC/Auj1KNlSGdzmbwc3mlVo
ZBmaOube3GnLqKDTzladBD8CmwKWEX1cJOasYrLV7tUUTLLIU4bgTnWQxya2p4TIJP5em8VKSPs3
djiJU61FfQxCttXVxN3xs9rg58kEjVwr30/F5cc+KVgkEIg44Ft6ocklh4Vse0TSOtugq6IQRVIx
DvxMbRpsOFtNw9yV3vmrPD3CAxmVg6FsG9iBHB8CSV7z1w7d4+zWfUR/CedLqP5k5eMuZ9ZNYRRA
RHn+Bp2nDMikCjmL7SjmQDMtrpuEip/3R4Oq857K33BLtlZfGG/5rPVtLVU4ejOk0wc69HDjRU5F
6c1SmWxdcyj8cjpPCC7oiRmarBZdHUtQCWluvKzCzBuMdp08/TtVxr6d3DFtGBEXohVFeEqLqZqr
KSr7o3za1BOAbM1sLKJXQVJlFb05cxjJZPBUJU2ofYB8jrormFE/Ifz/ZNP1kIPej2IBYZoDPQcq
9zr1SNjeUPQJcHjndkSLSNwHnR9cuEowu901ffB+jP2ST2R914VHqcAWuSSRoplaqGbDvNMqlXDZ
wB6Fly5YOJxjszWVvRKkdi43edJ9rV+pW9atP8ABIvBpxaSbWWRXe/Vc1Lvcmrvux4/EC4Q4Af87
rCD90fwvjYqqE8JestDK2B8WeKPPcDhoxs5UOLBW9YpjJRHWzURq1KXowLEQ0CPhG98yv8yxBECB
rq/Ntu5ddrmtuvBrsL1YAXnpoGUGYt41XWk+MBHmQn68dniuw7zEodU/7erz4pz3K4e/LaKQpqiw
bSdHGDaEGK10IgBOSw4vNyTu7+gFLPfg1L3qIhVM3queCv19mhiiyd6M8q1Mva80UEsS1q1CY3jt
Xeb5kn2LZGKPbVg064G8eHRdm4g6Xc8W+MN2l6j05ay8QrmjcupLJIv1mQLeFmnLMo+aYQhnDNwv
TDvbH+UtEJ6NAH0YC1kJ8ccvv77HXg7eiWIe353u7dDVF8+DM7AIQTdP/SnLCJAjnvNGUwDU/QWq
Q7qU1ZwvY/bostO63Al0eoP9IUnYw3YXQabdVRbGzyDv++JRlxpNZyhrwTz5LVOM1HwTdwu6ZjF5
K+RcGLRLyORLKrO43M7tvkzwisbuWJinCiEt6OEvL3QPfQZzK7GwFU6Mxp4TsNQ/hRxeDaKUNSTU
JpgEo5oyD8f297VctmFjtk225qo3UQKQD9EZIxZXL0CDFclAwQz8qKL1/ZlGlH1VFc/Lf3+Cchx9
8ZXg85JZxqu6gUEXqJNgpXihcu8O2Lf/iRD1bqMh3iyBs8kDQRPqIEvULzfEvtXKcD37ZvV0p/Mi
F/TN6iLL4uXJbVBRXqu+yBvgP+BFmTKXqssk7w6koIPn20vh1YiejfVVWba/wzoibl3bx+oah4X5
di8kKzJxP3oLPMSpAXvCekzTCK8Z+ui30FzMhgdHbkMTXvPhnukQBOT+Uj0EA910VgSZJJXYO37v
dC8G+OLfbVA7tiBz3JR54Rj8AGlR5EEX8bTJHZlmNCC5Q8xbxch+oaZ4ON3SKx8n4zUKrrJms7Io
AnM3qFee3+KQwn8Y5OO/2jOIjzRc8ML53AEd403WJix1rUXHL7xY+taO+Fm7FbxYaQrsNifMWaGF
trjSIwjJxJ2KbimPZJafDjioAWTRJlMa0IGjySSETZJKlVbOukPm7+hxOAf8T2c3Hcmv6F4kNucD
C35VYSJ1HDQdNdrvKX22aHABoWkwFJ19RYbv0dFrxJxS0P3KSrSoy/Hk3GrjXAcf6WJKd122XyS2
3GwGPPRGwxKD2k3jqSgH66cYTcWB4YyRDeMUZtPZS5CE087gvLLQrAmaLh51qBmoLWHkTIhpZd7A
J0KSJyfZhuufhvrRLm7giWPJ566v0LWU1ZRBQqIhC790szbKnZKEWkJNXRL5eiTGxZycWDApGPcq
42PnYN1WxHFaYUigjo99fes3b9hIntNmKqYKb2UlGavyg5OqsiflneB/aft7BKm2jyoj+tIPIPpu
4Yuq/GJ/eru14HUSDjc/OF2JtaOwU+P7REtqzGWFmxsckRmo1R4A7/u6TKlIshCDUwey14IZe3UM
rgcliewJynpsg+3/xoulrL/LJ8un/Iw5JBNro7Lwbr3mXP/njmcbW1SJj3lUQYRCQ8MR0LbszBUc
grW2Llu/OM3F4G2NVe6CZf6sNLcCj4hQyMyJmnR3qi9C8ZsEu2g8zqU4Wim91rLZPb4R/HMgNSNq
1iMarJFP2Y6k/GxFGtcheenmipfTRKoFm9f3/Mbs0Fv2hwK1gouyorMni+Kzo3LV3EjN483+P/EH
geAPZdRbpMVzYyT27uZ6wToDsyx5Qss27ciRZD5oUvy3vlzjjj87ZXFjFXTnMk/mkbm5x+TajgOV
6F2FClj7Y1Ebex+iT3zAndbfzGLLisXU4eT1PVsbAN0pRDRfMywwbn2rFtwR1gvh0VzZqHfx4D3i
G9dsGA4MVwUVgOMLlNwAEL8cIFZKw+D1wGJ8PXdzOEmMHEQ344L8PAHQ/VdAlkjdhcwE7+jwb/Cf
Dj6TPX3eNGmlF+MxrklVOuEksPa+bRAWrXwyg40f4/VjgI1pB8Ggzt0ghZ/XDUsIWXhJ+jV8UQGr
sBmi7bKftlNPMFqcS97AP8+fOMsa1ZPUI28+N7Tp8wjc8ohESzUBwhj0o6pcbaLzn1YAR/rz0c+3
2cuFuqU9f1pgF7XDRnbWsH9xNPan4YBMi2oXUyAuoXwBj0TcNTjaWLlrU1r3YRtklV1lcVMToB+4
Weaj3CHd+eKCtbjtz1Jk50SYVDoZo0PDMWzuZjlM2dsC0Zn1Cv1E56g3DLQ9RukBnPH7NJpX8KZY
RNzHAPPx3iD2HSTKRZONckrLKVVR/EFUnhm+yMinDAZJZyRv8kSJVQ0PiPn9UA1tE9kvsO77aQ31
mVjUKai9hBK02DYaAcifKrtyoIwx8rJ15Eu+ulVILOZvBDMl6dP/rmGVuA9oTNcUYY26ZpkY7e/z
JtifK4sQDIKzVkEMidCeBjuzxjuXbMDa7wlztcCv7P+y8+y0tyhvq5tLdUvQNLJg0uQMESWfbAts
l9YUG2I3ohbltb7M40gAdQ4W14k89U0o0wjANwMAVLstOJuoc6I/HB7khnCRyZku5aI3HagYgMAg
iatQkkGiGKmYTy5Fw4I6vuNG+ZBPKduy5+pFQQidhRJwQIolBhFzlflYTZSHTSqwqpAcbtzglU/Q
LcGB82NWytYSQJtvy1yTGJmSwe7a9DvXQQ5QXaFH8Mrflwts70dXzxnDmd7QsqSLRhSRWE3r9Mo1
x1Fz349Tur2Bn86tCWcFY350ZbzmS6IuSaWe8PBJ2ZX2EK0betnMpzk+NhYXfQZ5YKJM4qpHxCFB
rvYTlQ9m9b2E8XvqlGYQifVSvxks8/rccoHZOtmxhR9X5eWCwmIaNAxANRwLvNb6bq6+P3YkGYp+
ppLAYiRhoaisQSKXe4ZqInvuY2k1SGC4d82WMk1cryeqslGH5wYXIxuLByYLtSsQmmkotzoM9bVn
0LWxLqAcsCq9bi5eGQhWPbSUq1QzuOvHq11sFbrcvwAKWqGXTUXiQzhFnlbutDbpw/VWPJPMuwkC
lf0q+535d92PVAyVePTYW6vgQXw/3lRv3Ng0QPDR3o/3S1Yk0ot6g778yikKEARrn10HWFzyIPSU
wSE5kZKPSmUy9d+wQOy7BcY0CseaG4iaQxaOR7Gt1qk4jc7zeZnIWyEZbu8bkXg4rVuFoNV5Wgap
5upHhfrz1V/pZpXrFXB2mhWgyh1zYcOhuVjSCuDocfmS1Q2O+WPcKRnHEq+FYFLoegFenfnNRogx
UF4VmdiPaQw8kRDORX01EhgMIdNJUbcvfyFhnJH2aJmQZaFRAl5LPLIOITX6B/w8YI9q2jq+C6Ho
Mzt7uXdh4yz1L+IE1fa0vUMxU13XThNTu5r6UUOWzW1w3c0mnE8KLgpjPFiTfZzlZ+y+197H8piT
kFkYzSZJebc9+nX2ZE2xq82+ZtPxv98BBc62RJmH6F7A0rIibLwO83DdVqP5SCTWMuaTXRf35hLV
W/j0IFLxcboYM+f8QFwhXmfXdjd5YfUhNSsacEsgCCDNye5HcAmYTVr/ZU6sM5Yj3IuNdo/jjgO5
3gkS8zn4m8T5Y6uZMfu/9kts1RV7rmAJ1ZpFLLaMF+agemY0G1GoJtd21FuPnMW+oolPbcGPtm69
7lt2A1GFTFuss/swy/WChYLj41RMXD9bkFfOHCuMKI6ttOtPyvHXohQ2HVJYdFdnpEwZHHd4Ie1y
Z+HsWZHxzCOle8yovHfPVxYAAg/QB6AHI3CdgHfYcXc37gzHSlCDXNBg9eDc760AYXdAGpOjA4Lg
De+LGA44Nl/zyIkxo+uB3F1vwHf6s4ySzbh7qIOiKrZErR4LuRa+jq+MKwNpPT1d7zFenaZ2hDAG
xbzx5p6uXMoskGYUdtzQcVtESuAlAo8MVMRP/7f21OcTqA8l0/0xPyX8ySm9ltNR7+E6Zi/s4D0z
IrSnH0Yr21WxcQhW7tweFAtkSgRoyMgkrdrjtsXXtE0up9l1aAdZRjxDXgaMwf9dvuMO2G7HpScP
0WGsM1JhOjNSIhPTo/CR/VQBkZA4vgAmnHYC7gXbGrA8ddpeHTPHQgx0BPDvz/ApmmE7jGNknYUM
iRcP9ZnH4aSp8YwhqR4D7SWsFP72Oiw2Irt35MudOPXFE9shYLqU8jiMkkqqqqPUi2KuOfqZoKM6
OYJ8Cf0sfPA05AUOCXopWevjdsgTkiUJoRxUdCwGj24TltQUCsuRjWu4nZFah1f/P2CRW1A5xvoo
zBcPkUGBU22DuWhwONDW7M43bzvOAa0RTz2iY4pIBzaOCr9LtvrhFVC+ymQX7FAmXqfNDBbkMhoo
/gUNmO4tDewQOFaTl4uTsc/aoHyl5jXCk83o9Qw3nP7QhbPfJMR9ZXfSnbpJgJxkZ3emf+Uys+0V
ZUxSOQx6+btICLTlFf6ULr0qZgD+XQ5iRfUXh0AI/KqhfsgIpeJD9r5xoYlNYU8zhICebGAfX0RL
bticW58gFaZyqdlrOlwS1ckp5wHIfk1I4xVDMGLZXHR0aruvcZn0MjycYtKpJDg5SG2ocbP+DOsh
FY6JmuEfT7BIRuVT8i1EeetnL2xQWtH8aN0k6d0iALE7P1NgwKvE0rOScglkh272oE0D/QJJNgNI
IqkcfXUNU4AXB3NeTnwHHd6P+JH5U58F3H8CPa8RLaG+KA54HUTn3q7cjGI25/ktQoEDGCaw4QC0
QTr+blzz3l2SdFq1bmrUCZeUlIwEB2EOTCmCj2OvAE8q+wiza7b3tPFtjsDSUjsBUOVonQiTj3Kj
DCuNG5SYwN/a52b+F5hFP6urvSWPNfG4qXzSDRv5SoT6SGjRgqz93j+iW6ZS+eUJYo1TP2nzs6V1
FpSpb2rgWwvaHn3zUJgZCYujoi0jnmb4kIsgjxwQvNdohvJlNwrIu8APbHLTugXSFF/yk9Pi9maI
AruQLOPC3ry7jAzwheU2vlqrQwQG+H+3OQqKnfp+sMmLLysfhQ9KaF5IJ8kE4SSa+fKefcPNrpMk
g4BSfoHl6gezE3NUVF8B6qhY4VZPIlvep2ZJ1lEwwUIs1wLJDb3JqwenguT2oc12yMCTEHCAnAmh
PqUkM/mM6GhkVVy2SnBII+xkFcTTj5hiwIb4ZdG4TR08yyKx5Z1fEKPXVbTdx5wF5glj9XDtIh5O
3m2rasXrB7Jaut5TIfQtHs0bmOiHDH8G/Y/zv/3WI0xXaJ06mwfqfKi+YIcy+Vxm4ctZf4TaCHyW
ZgGeTztJIt2e1Y1ALTTn01Iy4U0Wuijs7C686JcGQasakIFgo/h8wsT9CM92JyhjTsX1Lde2keao
CDvI8uwtCkIV8nP5Ue0s+g2g5OEmhpb78Nj56U6G80LyjWQISN7EWzp0MFJlVtWGIraW2NBjD5kw
IcY6ZJiMhlF8xNT3ILZxGeth902FH6e/QJf2Kjm8Y5KXIlfnT4KuCZ9Lob8rNMx5G1H/My2HxHLB
crKLIcGz02uXOq2tJ/Py0Sg6tcG3tES/SaQuDYSIjmC35YtDmlLH1t6G/x0IDYamevwxswv/AWpo
9VaVVNKvYDbf0KmkEfVcfkF74JL5EbJBTQHoiR6ghLT7biQH/6w+iU+p/Y64fCJvIGtQAd81lUDJ
usSgmrYvx6j200hTtX/Sb3+zy/a9q+DZLopJo6Y910LvQK6/jSR6KntjjYSLPCGMiEeU+9D6zH2d
PoaEwe1qdW761Xqw8hKCPOiR3XBWxqkDQCvhDiXboIpbBpu1ZYEsDTpxQwDcycM0VY54MTCR7nWa
d7Rbi1Ab5+QxTTemAsuDCPJ5NX0bR2Y8z20dbgit/F4cU1HghzvUdzKwBk/uKzp1CwbGsvjIzGf7
873SpQhRjJznLEjosB9eWTYUIyyBnvgF1WZ0g3cFui2fK9M3bDybCOubUGOrQe6WjiG19XJwsoU8
wcdORupJ9VEHOwrcCOEZfZTmRJ61HZtXR3xBSogbw24xUjeI5xH14X1eY3EXeB8b3+4ULyKaUVmr
ejcCiXDuS3PgqdfXTzpodVCq2WZGaRy1ZgX6Sp9GvSivuBnwI00R6VHfKSi1mIBjIumjxfSVWVQN
z6VbBksNKvIlZI0a5rjPOqIVmRipQ5060SjRzF90lUClM9w4RiRTxf46M6OrTgFfTcEe4pVALQ8K
0l8oA2+tN8AsiKag/MOVZ8nfI+JF+K34ARf3d9w1SCsQ4qHSUzdu9IOXUXWMFt6HaxyTxUjS8Cd1
C+xRIpwjqPQH7SVECG2OSrJnis9ZnymjZ8YkCe7VbvJIKm9xf7LmTH3IPP6Hi2puF0nACIwsBNFL
d1BW8fsWJVMvFxF2IqyCkHOVBiwkMWb0R9tbJMoSM1YVS3g/a7gsIlN9/pDUSKck1wblRkJ2Z8PT
kBcAWRFyjuMqhGo6pUS2Pg+4BBGS4KCEh6l9eDRBcupXYv2IFlHyLN7kEYb4Tm/GAjuF24vTIbiX
PClq2acLy4fDzyHo+OZNjh5YEiuLAcEIWQgWCdAh/SQI9tGQyP6j9nCPd1KwOPb5otZIMp8cEB3t
TvDluirD7Vu31UyxRy3OpHeOcgTPjnkFQ7XOIcGcgqE4a8usVo5RqRzJWYP15yeA7uH3MDIyvnP/
vC0SxddKfo4yDQP38BsZJJzkECFt/yhRx48fV+WpQhZQToDPuf7CllT0ovdI3FGBrHtnUevECX/9
9dIdPlPgiRt2AOSnPvagMwsUdaR1JtzK1QVUgamlKa7tjnhzyCNsZyCyBMfPOw4NTa3Qk9cwSqM3
VAmciRbNMKqVGixlxHZnNw5oSjYss2m17vU/gX6c1nGYu2N1HmuC2lZ69wXM6CBDejKgtIeejRs3
gRCKnXo4IJLqxAkuKKhAzQKFJqC89wbDqUBWFUssefOOvB5BHmWxBDZRfhmz9Hg4xSA+BYOpE8E7
urxKWl0AJelNr9ueGZS1nC/vUcEHCcP5E57xzkMRmKyGP004/cNI5x+YSzMlE+NyvKfB05q8JglJ
GVMiDbbqilR419fUc+ZEoiy28Sm1HtZb0ciAeKMKeqSmSOX0sb8bquPkXsjnRklKOhCJWY8E73/l
lN0Ypp/f3hwxTIEqSnEv8Pn5ANPK0qo8Qe5Owon8Ail45mdwHGS1uxJFq7yOB7WvC1SVtoOLiwrM
9UicXH4LGDEdSd0lP1HAZ8ymBZei7Uzj/KPEGhmdWwB21usiE9XxJs8Kr0KnXcqfYK1n4gYDSHxY
0B0bsuLFFl9NvBEqL84CCdcm1nZ4qbqO9OXIk62sTopJbbzq5aREWcBlIMOFuEXYdcvLpKARtwOl
iK9J4MglI6XuFTmKT3iRfyJYV+Z5ojGjqkmGIgS2dY57gWzieK0ADM82RQqwOpYFpsJJf8LHu4yQ
ZXjnw/vIFBa+GMfT9BvJn5m88Wp+zmDLMYGS6L7Y12QBrBD+xorAhC/YnI0moBnzfMPdWUUakgWO
s7R5TAS3PonLvJZIgk4mmUhiGzkQMT7h2lCFUqSlBT/MoXPMhwTsYcN4bhADeFImPtMy89uHjDa8
YIJ4ZoaEmDX3b+5dZvehYSZX2/xBfd2MQSBNHJgx9P8nPhBFOm3NqTljNVzWszQjRjhmNoYo1fb+
CFfOwyAyGBfzKlyNvw2wbHlQfUYIOrq8KVgXH7gJMQK7hucnqGQDtJRXdO/FUhlZjKsMuiqRPavi
Vgi7r+49lgUruTiYdiKomgWGGHH/7kjJzPIPFUY8hUIMRzGAHaQCE0T/DqQErpPVUmRP3K4khHfY
qwm3Mh8eXaIFw2wtsIYoLlz/5WJ/3JSN28kbPOwXOJl4XsNT5Oh1/RV5Ik7fUJ7Mj7aESrbsIykw
XWAPJYbP5ps1pdYxNZxt6YhirS6+0xfvs89DonVDlmpyN7Ao0rUMR0IgHt+BbU4B37VsxJdgX3k+
gT64AF1TjYd8nvp5alOUz4ClLsT8HXihH9Z4+l4CsuDCqA86hVVWUgeGDbhQec/yDubJbwQSdX0w
M/dNUW7y+5xZREoIwERC6joqBfGm9dBrwKXXzQIm2w2hHMhqirc47Z2edyfCVzJCif9mLezUhSpU
y82kqlafSuaV5DdrJDtPMUI7a9mVJO0VtaPXMBgAgxgRSmxNa4eFTyAdZBl+FGUCRyD834L3e9eR
+veDYzRj3AMV05FqMQA2st8wYBhWnXSnY+4A9SaHL697gQpx6+azY4FDFbs0Dn4D6lBiH96UJ+WT
vxa4v7LZ/4U4akEsBBYIny1cvAXT65UaQJm4VEm/5TeGMCHzFE6lZ2IKQWoImCj0OM+43CJcFCiK
E694TCyHJCgQZoHee4CxN0/3DplDhyyAVxuUKcs68JTNgGq6f26StrHgxEqdizWJAU1GUoWYXLZM
3sLQDh9aZBrwf7nhvWSLnWw2OCROLSQLGD6mRBO5nLyPd7j+m02FEg1GBDwK+pHyrl9WEPpWjgfr
Yw1zpRXGg55MIGOhjZB3hSO4xcxJcfcIIgDzTNcZm0Dx8oBgMbLppkGgloNKSz6PC9eXwR38iSzD
XU/AJZGxldJm4n6+e4B7DTKyi/rX27pK0B0tSOiP0vqJUAZDkDNYgwq9teeSew7LcuwyerA4lAoz
qCvQPymplRS8TDOl2phFj3DQsgfHnaL9fGq2cw/GAe37qj2wmCGPY4kSfrvI8vGqRpdb1eGh6NK8
eaqO8+l1s+WkH48mrp4rfKWWGrCdua087sDixH+LQEUPBpKgm4YevgIay+WAysqBrSOd7cvAGWOL
VDV95O6xbitkgo9dRumZdiHe+9b6kvdVVmbS8fCkaBtfWfRJz2mPRN88aSwMo8iPavfbDcTFfbrW
eiyxgOXwlX2Z/FuzjILyJ3ATHVyLE7ejJQVJMKVvT0bRgu3K7qyPZy5QjSZZ2OkYVqr8i6UbSfYo
Y/xaRuCtIqEA1c+tMrbWSc3hkLP56oLn8v8TmbJigdOMyJCQgbuXT+OTUGv5k8MIOk8UgX3Nw1Uq
0DCg3fxE9EaV756rUlFiIkATd6di2Y/j+reZVorJ46TD47bMj8ocG45gJmxy4+FPpjVqR/rhA6hU
DCcqfP5ZgW7MiCgxC9gbQdd0tgS/Zx/BCznNLX2y63AvvSpkySEJ+mzgvOzCfhYnDo3FNI9mJTyE
dtvopx3gAfRKZ72nHLacpbvDCHp+EjZUfrP/LBo+8jbZcw5uM6uBAhf6QHJ0Ts6OnrRGrRhoHZkb
/99rBXGPdXVCRLSZmmBE2Ke3mrcj0qoDugyN26QCo3NTKT108KJSJfO0lYlIJBKMNBV9UEl734YQ
z/kB3rO1600y0tNRyASG/X1LFTtyHmB2zuWuAunLx8VwAdsnxYGVF0Mx2xSMD6/B6Xbhq/Eg3tUS
M7cqZTGKjRZOqw+9auvsejNtvEI+XY/uLk0TE6Ch6zMy3CdmdiRZ9PfpR0D396NI2+NVwHru/dCU
O+xkCacKW+muUj/vO+032ycI5HNOpPJQ2zOHxMIhUh+dRcDQWfiKYhR451342tETt5g9gObOKJhN
Lc/wz6UbJZOSH/YDD+TXSSXBMTPdK4VD9u1m+bCmPs2ThUMwrjXxxUTPQeseJ3OTTetep2ownGsN
gIo/8IlPMJonplEl3eBn3SN7HrFoXrtJWyFlWmBfKcsklyBjxAD8osoyQPVxMi/nVlbKtJzmayCi
DkuqhWYGMSw+gQJ7Nx9PJ5zRnV4GkQdRbUFyiy51/8KQLa+mz1pfBCP0ABoIOkI27iJ6zL0YaXJK
hMAvhs8ucZFJxg4AH7vgzqS4ACTrdt0hn7qRTqqfzokZLtiZOtNjkl0SSKMMyrrGMcTtfaQckxuX
xdZ3qgV6d8QXx3A5VfuHl513238DiYeQasv9suSzY3x+ziHt7hKpL7EB2hcqDhdjQswmrMHyVnIq
Oa2zRzbo1onqb0NcSDdvv00oHotJhK/+e8V3GfsNNdzaoO8y0RRuVvXtvp/q7k4/FxF+Aw5+mIDH
cUCsOOR+kPzBJI8+vuhYecV6emUGE5ccBOh8vNGyjuCg3s2ei1L2TaWLZR9HzimoxIWQjCVIlnG1
XI5CAmQ97t/zIGW/XZK+pJlIv6dJhPiiOVoWbvp9Y5ZOggSZNcAWKJf5ase6gm1DyptrUnhnqiiC
5HwipNUMLSzHN4TzQCshGhkdp1fsl9HF0qmErE4BZ+9ONNGNfk65vHYyC9V3YQwEgaudfhK7KuBU
yDRQ57iQkeLGRsU36d6Mm64MLuHntuETYCIUsXqJ5y0+mL72ezL7TqO1j4NGb4BTbVbVfpDhGzK8
byQWvhlJF/BI8TinQ+mai/RfbHwY/o3o3r7h0FQRAmDsC2xIDIeKa8ZFP5mjXFwp2kvQdaNVNxuu
phJjXz6LPTHcyRMzMeq7SY44Gg1ciZf4zWjMW18626ecn8APpbUnIzkcFtUgZhS6qHYDFN1+v9ml
XESQPiV7hDY4/WOPAgeWa2X8En7TpF3lhi3BQSC637rQZUl6pDI+eQ43UmtE7JyIpfIw2oy1bcUv
4ew8bhJw/KLaKmIUakY36OsnBrhhQ0UPGhz2+CC3q4JXqChNOuADgD7BFyqZXQfTswRhbeaIeR0b
jHw2KHsvA4b6upsVw/ymzRQhGmxAC7i4sFaTeA6jsuDJ2SipohA2Q1HnY7hYaEftmyBPD4dx/bLl
ASpcpKR/mL3I+i0uJM17EGrJDtlT+JawF2lspwV1v3KmpJv95tyEZZxoT8F+uTzVH9iBKWvLBFOY
17mOUhKITBjG/vnHzAAWfgnn+VklsMt1P47QDor20z3bo/VrbVQgTBiFZBVcunSCfgwTGW4MSbxB
RwHrQjq6kzuGyy0pmtHLMVlzR1rIQDkBI8faPgTG1dSfZ4CVxAdI8sOhLcYhkeN+WlGipQ5DGLFr
Xlc6TiK7op9b5/yHzn3fOUJIb/4A5ufBe4C4FOh6xrqVrxwb8wNIkjpMLKdIFFkqt2ncpC/ubKzf
hvnWamHoYscxDamj6d9zjYDKbd4WigPKoVIp9LvIlVAbk1/EBaSkuo5WMpQ1FC4o9Ld2fQCz7Ibo
hadT401RWbvJpTevpkScoBBUZMksyt3nSxUGxC09BTUC7HipK+VfjuL4RdPmzhE21cUok4v6M690
j/g7uRUbEcxifDWXOO9nK4wBhfJHrrzlB/zJvKfts+OYBvGpZJB22fWhG6zKNpgGM0zI7q36r7qd
xNag1OQAU2iePTuoz4AE+Br/vO6wzcC+/i4biLR3x3dXG15C8107SRaSzV1xiziCV8J7lKcKCYLP
zTw8sSy4an08Il9hyuuhHRX8m+XcQLKy6/tG1YVM+g0oP08cEfspcOS9hbNR6Hu01Mboz7gQsdqV
ofZXejWA/sD9jLYBu0Gmgj5PpIhwe0sp49cwss7ERJj/9lm0a78iiDG9HRKDoE7tnbYD+ayivw49
2MsDb9QqEgTo6exs12nclT6OCnYu3qw3SxKokp1rkxxjMxBXhuPXN4439hbu/xhKYWtqiPHA26ee
xyyDElUpIYJ5vdHlEB9O0eqUKBYqOeRTsGFrFfjWvUqI9pn+PeHC2H74gAmitAYgjXgW8MtLRxzf
9Jo/rcdnFGiLvvzg50/5Iz2V/qxCo4FahSmoWIG1XhiE69iIijh8aoUWsxxfMHD9Qe15fQ1R6xMf
763deJifEMrTLC6Q19O0lWPdnm+pAfya3ar1tPTbcL0+wJycCICfjC6ZmXXwooWkfxlEeTomeM+H
3tZLDe1GMoHV7QKxkmY+hy3AADKmHiVzj0Qf2KJnmZRUp3sL1Q/TG7jf/vUymEbvEQd4FUDLlsua
XJPDUKpdINS5Jp/2e+9DxpLWLzfbLEq8n+G4nawXcyG3tbzbhPtysJACwhVxWtjz6zf1+4aQhyTh
evxXSYyoED94SJqjUepX0nchZ6YStOH9y+5uUklRfvIEC5P7PeNhapHYxj9gjE402ujN5gCkE/du
hXL2E+iTQiAnfBhj3SZA342QFnMNjw/ZFy8YZ4TXu6ovpKk5IyTenN7oknhXq9vuVoOp0pwDZBcx
uwkD0JUwSVYUzRYRQwUqEWlHm3EEnr6GjZWULSaXCKTE1EGMUaTswDiJuaxRnFKhO9zk2i+9UDBK
C2oeCGiSZQMGXHvMeQU8WjE+BYxZ/7+ViyTjY2v/IlCoAZTG4sqpf7TwNbV9pO5TrR4TkCZL1C3V
g85OA4uhZqpiVaFNLL9wgajAQ/wHEcVwrv3ELHt9tfeiCMV5m3EiCGPanLxAe2dHY0oawVbkmiuX
jjVN5qr7ajqUMpTjf6I9ahAKQ4wXuaB3fsFcP7BqCVOcusmElyM/stBiMxLxhOd0Mugr5eHfOJHA
3vZXsdbcDRZ1C8NIos60Y1yXW27nEEgvvYnmuaUXCZA6ac8nJ2D9EO0Sbpz8ET7zYdh++tcB2KZ2
9GbU5V1gwC7VeqvZh4klWs5RK0VDlFiyRyco8187qIEUT0yWpz9DjpTnrrj5kc3Yvp7qC2IiRm3k
mhnSDiSsCI6x54+sl+uAOZXOgtGaRbLmbF4NEF5jby34MXJBSBBTCEuUKse7TAtk/e1KHRQ55UfZ
evsOCJ8OF99djcba31gSOUjlLMyOJvoZoEtwkuSAZuwgWGX0OO6SaoFH0Lj5QCn6c/Xz6iZu+ifI
ZUV6SjtaLZWay30vsj4X/LMHIYSARqljiiLdkzBSfp9c856VzneiU6yiUSXYJRrPXyawYnDau8Tr
f1fJRZ6LkzEgQIl4KHPbAtA+M5QIfvv+X4wkqLJcQV/H3s8pUZH6RjWm4CTSD5w4c4aIfi57znyf
JAYOsOpeWsXX6pCLigBrX1JNH4+B3D99ys4koB5FUIZl7xL6grY6uJ/iXYdYev5TNlPXCth0L+nc
hxAbxCb0uz9ALD11HX9T/HwX0F8bASWkHsTEih3mbJX4O7GvNfkkCgyLnYn83aXGGPIcVioSMXT4
g6utHezYp1dXg59IXWJrbOyPGWuOhtg8wq9mwERn1vmaE2V+XwSueM5iA0iWMvYEqS5mxcvzb5s5
RtePwdk7Hd7Ab1+CbadEkl6GaMUKJXQHrlmGoKfkxPb992XtLQ2vG8jPm7k0z/l7o0fBUMAs49xQ
0if4cuipYqRyJPQnd5R3RkQtTiExRVdRyDYZNDBz0Xp/TwHIN+9R+dLyJ7E0Mn93x5v4kuLrtjgR
Av97kR4y/hMvHf6uVdBLM4SH/9LVMAVTC/yLQTaCfP65hfDHwD09btGJzLELu6GQBdpap3XcE7Hm
mOlwdw3D5+NO5nb6ZtAmaZLXua1HWHBa+LdBgJ2r8p0dGrd42k6kdQ4+qW0sP8aYTAEMdEzvsbxE
mB9UpwwAqxkgAGoH5h5N7kpu789XM+V/EcHMMLzOdWX/r12WJ+dwX26DqlibS9shNd7LPd7De1TQ
SN29eJxlHp86USLRC2fRPMjomZx457GlZK4ho4FLpjsXV55ceDYCzs99CS8Hg3purWTHTifv23QR
JsZ5+gY9gan7FY/PqI+hVqRM+V17bDxeP0srS600keP5q3mEa1VRYo4Xm12tzq/2xThgEtS8gDVo
THl68EGO0v5mqj5w/F9VVHCfrQCyYqZjSnsfHboIpfdsr2TZQhpcVLz6AGQ/S77gLjCATHUpnePx
+3Mkz4mds3y5yotEozBq9d/cQCQqgiIKu308kKzlYRAuQewK3NWW0rRcmpDL8v/NruAvaYgGpHVO
01SwDDIvNGGsmRIc4CMvnoPf8mN3nOE0r21wyvXMZvyKSCsWIa1nrnTa4RbTlnqAK/8yEqsOpjnU
XOhoDpd0l5afm5wZZJaH+pFSQ0ChN/dGa1kLUfk3lpXxxTB8ljiYHRP3jmBt28+7xHsDz41nssrD
ER++02KMC50ywIA3wG75gE320gHi4CedukmCyLR9CFHiZ726xQMCYU8mrh5Gwor4i7zKkR93q7YG
fm79lpaDuaOIBBb2bVmz/l2uw+ZmYC//8kX2MDXhuYZ0S9NWsx1GKyHwkCj0HiPy9CNeF3DY2sPF
rkrYVUq38WyHUxpr2WiX8gHGN0TC38mS4K6yb3NwVcaKXF6UlfZPPo+D47Wp9U1Gd4iLnEP7khsu
WazPIjeUm6g3aaZo3xIXErCm0BWNRUsQH5Fhh7UaBP7vubTevLnS0T1wTeUJpX1pWJVdPp4UqP/S
fiWV/pYPe9ey0OpNgPQZrzqidoyoeXCvRI0eR2esKtXc2i1AiLpL/gKDzQZc19Ppf8P31Rz4/uB4
vF5FsnNNMkAYJeFH7jA+eJ4QCDdkFoV6raI6I/61eGiaHl16djrPI11Spi+8s/VXIJ4fCkwUnbsU
+GrwbOGAsd6sfCsjcJ4t+9BMKq1/AfjDL+nM6wZ3VME+9yXT8aiCh90ArNkC01uTnb9GfNvLyfOl
fxImnLeYFUKglzQFKzKk/mPsKpG9e56dJxnek5D7hHr2yWlg+etU5OUubZ/laoNI2AFIqZotG08H
ObQ2hbDCJ7/CHTsu3YfkmPB+ardv8Opt8sSXU6+Gl6uRNISfk1ZDpzb/DAdD7dy1+W3jVRJ53uXH
CxexxkoHECKJ1VB1LZItmJY0Vn9SN5lMk7CdAFz6065813mDm6XbcK1hzcG4vQTFpCs5MQ3uXfiH
YLImwhpNyAqBGMD3GdIWdcvvNuxuvvLSZQmYikIPGA0zscZRdqIZ8t8IoYzo23UYxKBKtiYdfWvt
S3VRqHhhKxQmK+asfTs8nljert0dtBerlU8/d0jeapLDGT0bSlLKeN3ME5W7NM9fpKVLDfZVCb3W
7vm159SaIPdXPaNzWP1+4wOnGU13CIb3J5xQC80s59zCHGqXp41u3uis2h9YcZDGrwXEjw73G7c5
PyUWJYewrdXuAuUJ/OOabLRegLwtpfl8diTTKxbG6wRnhkpmjNOVtmpTAl8uu7YHHmzRH4uAi0Io
+kV8SDG2qFDNX0z20IsT6b68x8fhtMkRYVPiyu04Bn27yaj86nfSzeFahUm/6hX2ezrSqQ+/KWOU
u+8uiEDG71ZkFRd51+LDh3igzlsiHuJdPzIgSf/YYzVImiCX+rkx7Q4mYBbSGnkNE4rUMpWvcSLw
yTd/yDQpwzVElK8cHEEkp0/7oOimap3X7jSpeeXuEPWxovB8iahjR8tou7dt7/GvFXMIkEZfphVz
kETQn9cE9qk1N/zZEMJAoH0xBCwqbLEHCIkLpOUXd50G3ip9vghbDrezy/Pg67R508sqB/nFaJRH
/TN0pPhiSJo8k0+yK/YYuSfp2a/L9z+NtRXTRIl4fiXbFDu/O5tupLPmMhjYFZawFZxCsYn/CC99
oc8Kvthq/WJg09y6pKHmuJ5lcIdAtwah4IJG6l03gg9PigXzEm2y2FYWtNTRcT8dRyU8m/xV1Sh+
RaApvpl74NgikyygK5nGovzHc5TJODFPWwO5IVeeTGNlVXIqBBHYa8JPrX7zk/3HtZjApSZF8VAl
/BFrDkhMCClyBhLh/VM4jAYGr+Wui267lDgaiv/jfhpXyIjYtbcHrie4ZgeO0pJ60hYuMPH6e5iA
WGBg9Lyr5QTlbC2xsrZNj6gbRMhLDWokJw7ex9UEWLi/JYzKW8tzpkVm27ZuPMu2hS1rlaVJFFXG
0XmMzwgiRNygdZWhqgjmZo5TOK5LYOuEimnwKa1McJwS+IXUqRzq/qKTeRM8XskCLfQu9WfJuIhe
P5xdqyM068+MWsf2Zh7DUR3jkXzC/bV7yMCq43vYbO3Gus5DFbaBYoJVzB8acWvO+m82EgfXQRu1
p8zfJPvmer9LG42MQbFfLrDJA3o1nnqFj4LTNdpimD5SwlJjucM7Wg9SpyxN2esVLZ3Pdi0biEQO
qroeBnu32NP3I5U4DuzuflvO8MJ9JpYX0G6WghGL8R9KV1R4venDLHlIwuzXk68K9N1VgSOHp6rz
hfSV9xeIC9Hz87Lf0mmiObRsUw1UPRmU/M6ARJEMNJckL8SDTXQdAxGNr/4uD4YiJfaRgn2WXnwX
VnZLUPGFntefa9d4+/AFWu/QT/iNn3unR5cX/7DAv0K4UxMA5vQPHXGF6gxmynhi1nNBw62j03Fj
iA29QkxgcwZ9CyXA/UrZ2TrmGo9lEjKVT5F+NfFutjMzM0tu6IGHtXJEEb4jjiW6gm0O47CG2EMS
k7E17EmKjbNFsXhOweegRzUmNrbLgkOydbFmWtNwO62RpOlXBnTvpgYAO9Nc3wwZ/0G+e/+XsRZL
lquv8w2t24bjckTKn7wcrwiZdHvZqVXwF3im2tpnxYFBoJO/3vTVwzwBEADnmJ/xXMawLQZf2wZN
gURRNGeoJbB8fM19VVrQHRZclI9wJKnmpzLRy4wmnty308stEnS5sLe6FBpvg9jGHbZWP5mdo0l3
yKaHBn/HD8tcpWzg2EIXNX3c0H1qkYqXhB5Nh/oLzv8eG0sdOlTqiBgpkiEWrGXrirJ++DJ+AO2e
5p/asRa32vxX71JH7txfRKbdUPvbNSnsXfc7Gw/yAEFTDlGOKMSM7gBqSKBVvfN/+SA3BwQrhWPa
NR215CglrX3ABnkoVjkNgaacTI9a9K+dLQdujqLiavkiFgEApMZmSKCyfirhuWzifwGlZfkCQPr1
BUnyRgQP6yqpLeNGBh0Rdwuya54tNGx1kwQEKibnrKx6lYou2kt5vuuzibE7rvsV+NhbdME79UoJ
dNJ+AUvbfZwgUwX2gCMVTHLKvakQogfW7Y9yd8ahhQpcOuAJfAuzUmBUAG6A+tHBIqyk7ciW9/kO
G4HQ8RJOKAcu7gPgJ8oLHJsJc1r3G3QtKGK6kKJYund1D5lISHQUfCs3qaCYNYFyc/G3AF7UVM1g
uhRZs8Ag4bYtefQLba1ZIjakZgRAnX7LI/6HaiwO/AqgHK3db86Z3XVf51NdFDc1rcKuoUVE+p3x
97DfxjsMIxhyyZ7H1aEjtu51IoRhS0S42j1gW7MHgH0AXwZse8xvaHhg2eQ7Dz1gTpuvSYOmZh7m
y+CdhWwxIH8nqLQxr1GnkKfmsB67DlSy1uoMrgalnoKa5/tLGSN9rpf94RqiJGvvKGLiXj5d82Se
yzHwLEN/JHnZYHAKO7dXBBtBy5wpfuMxJuw5O5cQBHXD5gIuhKB0Oo6CNvoLj823EpQheVTY5vxf
J1nPUzxtHqDDNQdakXPLOa4xRnpoUa+VxkOJ6GRL87kNIBpvYEcv8TfaRr5i5zWqIZ+r6fJvgKMI
/E2bKbEJ6F+xCeYrWcdtYQjPq5TGMhVbSmDOh2nvx3bp7lATUhGRk9zXuMBBXGgGlpDfxu07JBRB
DyICZ0MFmP2YaSh9N9+ElWXAdSRArZYjGE0KdWKiJTVhLU4/XraFK759x+7s21yicDWev2WOddUq
2INuAWgsF8icdffza6W9TTEBR1P4ycfjMCVA7CD8XgXWu5SFM+mg7S0R+pYEMhuf5rkTjANvJSHO
F4P2r0nYSRVJUZ9la7MiDaW4TLjnvsO940YgMgCObPJVJD8P8SzVwODt6zuyNZbkhhzrkJjTmK4V
bFOUniqUCx1SJi+lVxNLnnnd92R2cLpmkE9gE+JKRXxajCwxAzopfgfru1SHLo5h38Syg5/RnFzF
PSWXvN6ZbtH9nAU1byIawmrrrO4MONB2IxJTpjVFhKmyAl06TqaeR0dF5Ydrxkhofi3NE3KtJPmE
7bIMo5kj4dJEyzv+et0rLm3IINeICMO4N9t2Ra26zTT0K8HM6wo3cuyDlznA7b+wfnsrtEWrh0lY
pv/ljpyPyWJt9Qdkc3tHuVP0DUznq3HNFkgNoQGfRzn+yi0WX7cBi+e7PNDaUszR/bjxgDS1sodb
O09ybcMQkqIhv1XHc1bVmPHlB+8Qdl544nmokURntq+Ucugt5tSZDBe3TBT591/WxvfB1mvNn/kz
6KglCL/DF29SLVbo6zyWAjYGDLh969v2sLdWR0r1VHFJm/92Jfq+McIPqmj6WrkBDffamt7ZLI9H
44mH2Xok9bDYE1UjJvm4QbGC7CFrDj/TYq2hykH4RLsHejfIkrYSPcJej7oRR4R8LdgcrPK7m5wo
3gITi4AfWiOgixbfni3rueaCEfZqq7+5LW9cmcK5u1zfjhGZh/xLkNLaP9bfaZCLA8F8NUNEJ8fd
HfjWES/4eVY41j4Rve7TPwpMEo7tsOc7UUa2LpCzM7IsS+N4pZe6GllRdaVsWXhltKvhRr21N32L
IWOoM9RzjqlCii8j9dRZmjySdapD8dLHY7W+EJre+dkb6H7jDoZgEM5UNR73QAN6Wg8efWJwPWK1
Eg3uLxgL8UgndwLfB5Sn4m+ntdECIJJu5uTQ7Pw3L62dpIxXDk5FKwmZz4BOSpIv/TwRKeFiYTAe
SRpLeu4Elcg0d5iaDHFRZ/4gvq3F65HLRwUo9+yS7Yel9gddgiy3VhGfmIl0jfRfOzNQv0vGaO6o
JSVSdFWjl5c+oPi46pa7lGzMIcGigTPP2Bgx7C9Yu+Cm5807baFw71D6bt3uEhvsa4vcT3kBkBTs
m2JpY4M5vJK+hbyfGBu15So40ZGs6z10r3qneWJRiJnX4ODzitJiYNHptSNEm7w4j/x5YkrEmSdI
o5xPQZJ5JqQrUrDV6o5Bjrq6NdvvoaL99envwRLTejC1ILkIplV1sVfJzwdCeIHNMpUloDHklQi3
6tIq5iUas7nNyZqTwI368y/Uu/Nz4kzkE5VHz5uHurz/eAQhQcz6f2GVWIPpiS5U42r10Gdtimqs
x3lMg2ZMdJdzl8uuWpfH1/rdF2Pcb6tYQuSxFRaPr5FEp7epUamOQMAtNLh4dXyvn3p/3/JRRqWy
jo04Y2WdZZbpyRLGTtn4tTSO3TRZ3SnEm+1ENC3aHaZ0//U9Rl0HiAbotBkEbhSz89o2a0k4crV1
eW7CG1t4IOLXvLpxE4d0x1X6udWkHZQmHhiLRSkfRk8jYnO+2aTlAJhMVB3FvfdG/QdfsG/P3O7o
CffuQU/E/NdOqLHCtT+gvkHSFRPPG5dDb4VuWmXPuA2+Z90p0sI112WOElt8qWk14FuWO/q4znJm
+zKlMt7mZ3VwSf5hpxWg4Lh8D5f9vKvMWfy4StZ1GZ/7IIdibQ7BM77nkGBHTEJsbM1WQbbQeoOC
DkGBvazVjJxV5JR8XUA5dgb+l4cJPKz9mIi31VGJYC1dEiGjgDyTGFBcNCJdQ78cXNPy+c+GSdZu
Km26Pi3xmMCiCTXf69gMz6WFe4AaVUnRxtZmrWAVr7shDXH536PtTupRceQgIY38ikCrkXitpTGx
Yz412vvE5Z8whph4Tl4TinJA+Dm1iEnIhxWMO6c8QCuAcUVvCwd2dteKQ7SqONxMw6VU8ByE0pn5
I6jjjGVnnalBDVwlQtDHtKRTtxTL5uTAShun7Twn4nmiD51hjxcnXmZ1s/yWj6R5q2x1kgC9LStt
VYC7yX92lmalXtB6Yza+Gp/NTiuOYGhixRFQjDccbXRRI7+O6eE4VRHkQ4JS29mf35bfQcZcmL94
njkOMmy4qt96XeA/ry+qAGH1wMPA+yZP/suBY7XfZslDR3xhU4zmC1pV/SAs/Tv/57DYbemSUwCI
QQ0bVyNtOxYvyjfR1IlJf8cT5js9Zi0mrh53a9bEvyoqAZzOUkikgbXqmHpjn03/vLIPBU3Wz2wq
sF+KHGOTMidsPj4hPKVwFck9zlK+tzlN3LO0tCJn60L+1wR/PCbhnjF4HsSR6yXeqnbJDiZjRfa/
pemPjW6uqbKZlp28AQerXFlxszXdG33htk4A7QAck/b7kbJo0Fd2yY/MoZiYVO7eEdHGWE6Fmth/
mqixDdLArMlKupLqKeacaFKAi592Z1N1z/s9I2bbzQLMUslCpwUoveO3+q9iufDgo4BNkuwCixLe
HIN/tZtAHHDxak2OsoqU/52OF0KpnTIJgwllf3xt78hSZ/aFzvBJz5oAjNuKasHb+4cL4GrmDq84
0FpqiTw6XZGPWuUIS1Hig//K0QJ6nV0MAbOsUCGn9FcoRsQKTlfBzuUi+M4S7LdOYK3vbOyGgkfH
UaCT+b7gcxKZ8jgPued4bJRzLQtdok1hzE9kcMpmFi4dhXAD67NXEsQWAvLHI7tJu/0oePHKbQEm
MX9BA6Dn/b81A8V1qZmjoMqaqJ6vOzDsYxw1r61dlCsTObB+5ZCVJPtZ+JKobmWMs2AVyJMSM8xQ
g0aUaTV4zr6wU+DVw1ScpfLyWb9HdXBLlzbZf4x2wHSJO4ttcOcoSibZvGIpOGigHAWfNUYcUtyp
c5ZBFbvGWC/heyihz6up0UbLg5xOO0a0YQ4SCN3MqoUtAEBqCeWi0dj6tsuu34xFEYNP0EyAixZR
5Q1S0XRMkfXc5vquiI2Gzqmc1Be7wQWLR07+aChzzjI5kqT0Bc27JKZVRKVQzQytIyS7GhuQbu3s
1CqVwthlGasL54n/vCU6nExvg4kRGGEWHvj7nw44PHlmnVJElx0s8q3Duixwo6HHdP0bkLdI3ngG
CQknul59SauoWee269YRcJ/c2ahCJCrVcdd3kian6cYDsrW1vj6U4+bbuOTnu638oqVBqXMk841v
HBGpT78RMNl23wG1bNyB+iwb7ChfQ3xx97YO8WWML56xipffzW1CrAff5xiIkUTdMrOcnTogCU5J
RiYYFxBPbPPCboBoOSrtZ2jrHK/X5CxL5/2Jop9bIThAQkaxDnpKY1KbBIvutEJ6CSR8NaIO6aJt
Qdo6fYMAljLNSvsr1wk16mzxsQCF/RAETHkeXfRTfLmy2fXHttjWkj0/SkTW4K133XGTURMk5Nw6
/R5BHdho6JDMwkadrZ7OtjHTswgcwOCiJL7Iv1G3/xYeLNt2WVYrNMZMzt+X2gZJ9cEg9wHinR+L
9QOVKUWBlJztkRUrPnba2MDOU/UKw0W8fG1aosgVQliFgmJ5MPF1LlY8gfxrDu1TDIYdro0mt9mD
bAPQp+zMqYkeQeFp5pYMkweNa66LubbXC8i1Jx9oF03w7Ogm+FUSqDyp6OO+i6SKzDj5Nh6UnbYE
Xw6MpZN/De8vPUguprR98Bio0d3xqjgM4yi8pmR/TxulDvmjksW/X2pSCLe8DEz5nx3MXnlXUG+f
49vrWNxJAm9/2Yy+/YR/ozz4xAV45jzPW/28s2wg5sCdkI4QrUuTlVWbELRHFiLG0j1+XJiLK8JL
5maI/qqNjPuVNRZ2v3pbPdzqgj4dvNidDZwjnAYGA9JokYMAocUzvE3hShw9PFw4vRmx6it8Due0
a17WggxFKCEgaHObV8DE/aqcDuA3EUZr9TvrBFF6bKKTeGsRRdke0mPSNsl7a1/PtFwED9FMNpM8
R+5R8TeGvMVX9ImuwzPOIy6qxQUigqgRWO5z6swe//ufZv/+WnBQPHPKu+UEJXcaqf07i+eEaBzM
WoOeqNzMqjHhTmNjJ1G8aOqCJf+GjIceCKmc9WsG8DPn3on0o+Kbhk1ljKJJxZOvy/oQA4Il2nkf
MQJtYXUML9na59n1rrsTjpIsxikrteJkVpvoIzlZYbB++QgUFdfJyKbKGPizUJcjKxqtLjFWyjyp
SvjUHka8zNuVafFxkQMKix08o9Sq28RO3mpB0T6hME/27wb7pAKmu7TAaE+Pi4Md4ewMWZHuFD3u
6UEPHVEeOYOD/meGYGsz+4WN0Fo0YwskJ6kXwHJyre3QhnUHeQ6FAiTt9NzbABcTrKSsVTkleoOH
0lvnZ7yt6T/zT8RCtyDNVLKvxDvgDteJ3WMMEwK6H/59iQCWL3qjRUQiF3mkcwVj00OaQb4KvoZR
4ivp1yqaRJK+n0Y/giomqJ84xZf+vQCaJ1YIey+RIiAEB6B642nDY7g6/XVbJYhb/tRdIT36k9/w
TZ8xxtIVai53JR5PD4I7Up4+lcSuMYGfadtatMhc+EB4sdl9vJw1Si1q4JoH5Uhia5r4styPap7j
RsDQr2Ky+dZ6VlslWV08CM/3WiateLnm1GG3g6i3tWKqXLF4Xbep9MOjX0WsyszeWyevg2YvvmfN
Ub6nyXnhLF8rpMsEKUL/SuZoXbiIU/nxz6QDrZTQJB/ontx11hHRuL1q8hblvZZjIOGxFkLlOE6x
nHiQpcO6x5y7FXuyBjG2jyJ+kxsRPE/2rZX2ogxo/c5TardVLobmwYKDR915dpTwghleGmk3QcoF
Ua9gTTdhOMPUJ4eOTNBQ2T+yhaw53fcA4czf7T9XW7e4+ZO6MY3/XdM/F2AwN9jrhEwd+zMjBiWu
AKbor84CvaXSsNT/9yqSQ3Tz/1Y/kKwg7vkkAa2sKYdPXFxm2jH1WpN2k7bqw6F/Opiy5d9DmMjf
JTIBKQns3xH2HdClL8UYdyrtJgvT0I1TRC7/cNOoS34jRsK/SDOBjbMWbrr0KrLPkKov/GC/RgSh
LeeHfmAB7vcxtEkQh2OLaITxHXmTA9+XJr4cD4e7iqSU4RWqbX5KNMhiCguU6CwqflP9teAKYGoC
0TQe1xjlnWBpH1ZGDlXOnDk+1eDACR/Z9GMwWXaKNhfTuymqtFcIPKD/nwtguCit2UcF4mKg/AhS
QwsdF6Z3GPuEimL62O3fhV5NQ2I0an8lClF6I6Hx2ADU/5cnZZZY6lvBYhMIt6osA88DQ9REZyr0
AHqLwt7wBQr2Y/yjbgr42E2rVcENXQ5UL0MFKQhbCsBwUpIafTqkfdUxe9pkKAU/JS2K7XC4vaX/
tVZId4rXiyuUk5+yoKrLKZ4J/R6SGKskDqZKrVGOmnIrxEnaMvngRmVq/MKScYyaqvwdEnUTXAe6
r0b2n9f1Pot6LFIJi5MFmFWZkM4Ur0brGvaTs3euczZ0S7c07Tumrbv/4odcYmKRXqLQI310s3vJ
XbtVIfEzTtj6VmKpG85sfkyBP/wv39cnstgG1unx2hUH2Q0qqdkZEVZhUT+zGm1z45LfHBU0erOb
7X980dc9G7MhiSd3qWQ4HClgRrGGSEqpsIvBPum5XVdUFdJ2AjwU0iyUogEpDUHl/aI6btMJFpVP
N8teXkq7FCXtlZI38DTzBxDyEI4dO1JO39tYHscAIfcni+IKcqllz0XUXop/Agmdsq7zxQ1DN6nE
lIcFw6RQ7NZ9P7D3tnB+ivSBVhPbVYsFK3mP7TPGUlGKIG/K2Dn2KPfUnIB1DlqPdalbgVgdn83g
GKJ7OeO2J16+KlhlgcQVAOTCEkSwJ7to8wVOrhlK5mCk7MtaoLtRpWlhB7Hn0vyeXsnufYlzpomO
6PRsQfk53l3GDg+E9pVCN7LFEH+lq8VnOcOxqAiZCCcZiibzkLWNFRPIaPd9kTYvycQ5j9dLlK9t
w86MT5lStGy/OFPkfRYA8bq/v5UL3XwXMpu09rQEn/xCPMvt+X7gNsX9U3P5oBVL4MkuWQ2lXspP
V4tCvnkcl/fNqqjfJQcoaZHCvtsigMltfN4++ykLP+lD546g6uCeVAwGi0ejUeh1tJ73u86hyEKR
tfDBN5IjnaETv8EWXfZ19C76sXcvd7/toh0ZPo7LHfeQhT/5NUY96Ol5OUVwDhEvfuFEszd4AH0P
JgVQ0VIuJNQuhh+dDoed50zsOP/XWL4tTUzLYOVVfZNk21zQIKyzS4lJsgyXxx5prXnTmdHIA8SH
4JosuquzIawHGXpRk8/n6IM9L2/9eguZq9FIDX+1CSFu94LCND2zvi6CkzQiAbV7CEXcsKpCqm5p
fKz14uGgj5mcG///RHncr79IkMgsqio/6vdZFkxLkQRcvgunalJRC1eBO7yzjeYIrw/hmb+TmSSd
McOzouo1qBp2G8EkOvpQXsvyuexl5HQmTRAIXfT+uZ0ZsGHFB3MY5waR83YvyoP5RCgpb6um+3ch
0lWBa0lss8o3CQ4SwCKc/CCjkg+xFCxi5CCc8+C9X4KNh+BoUyl2JgXPxXqLGQ9Wzfs7ZlqR305p
bhr/QcluVcX09kTQ3xdcykKNDtR6+ypWNlZhnISJidfei9sgAlLV0fR5seXY9g3u3ToO/uPTHx5P
2tbAKMmaQpO1YF7AnrpYi8EgW8NJH4N6UtfIxqoc6Ucmk6RiPfqyr0U6VFycYr1QvD213UE7UquX
vZ41S61djyDkc34/5LadedS7BX++Vhkj8++cMbvvnZNt6YeGCeLm+IbuEInWeiMIjE3BI4r4Ioc+
hhlffDQ7oFL5qSFeEjq8X5oy0oaNAh+hUnA9SjlYxlBlUyDoyy/V5g0G1vCifxi6vn0xYSweWGxJ
9PC44WKLODyr/E99i89hxcGN5KchWPz0Vw54FRUW3BEW95KZav7K74xQ1R0mH0PFx334sG8CCmFG
bYEeY6sqsflUNnvlXEA8gTfuttdt7giXjkB64tGLQs4S+kN+HAArzbGeZPmOyDAzjWLyb0Fua+Q/
TW6CpchLDpf0WfsZn4Jkdu6/bYxo64HWQ1U45paq67qsXZQ0K+GVPCWLqu+gxqjqIMD/pW/ftHkh
uEHCFv+ETgjgaLWhPb4Cbit3L5Pgbgx7SYbcELn00ExgBKhO1UgDIXnsVDu4vrnfdJUziIobWyqV
2/70EWMwYwWgF9GPoXOpBiq6R4GU5xupK2wgzxglSExDtHQ2j4H1mi3Yox2FQmA7dsYa7uqLyK4p
9DForksUedp2WjqL87idh/vRre70zsYi/U+PSTDhczkDDnncVjG2UsyGYmA6PhcCYsKiRlXyYQI2
XPDM+tRkqnSDAQ4wYtTot3E1h/6bcWMygESHwVS0WGlY1noMV3VVQrVn0c/fkbSS9ogbMT4CDmK3
HQxQlSXb4Zlci9MVRlgTeT8VDk5MkyLWNMXHLe1gp+hW8yoht2uq0QHMARJMu1bvxKZYDW42bB5E
9xS725mPk1RdWmfpzCq/kYND8AENXp5kIEuN62UJ7fzISCWm0Q8uveXaSWAfkU1rgf9rWSZOwX2r
NxwwHEmfojsNwSE4z5yIPUVUheU1y6B0NlEwOWTHDjvGAW3buAW0e2bZLrgVtZTZoS69Uw3aFIR1
qknCsiETfXz4ygWtdWidXnOxhgkLF4phFLXsJgY6lgTsMZD3oy5J7MZRhHYlS2AiNdH7Q523p+Zb
oP6oMbRSe1Wv4wNlgrJ2PbJcDR1SsIWbQG8gEJhWVsFr3yRPVMygqKgwpCpgbEtG2JJ4Z1r7p4Ew
Q3Brrzn6HbsiVn3K6tloV14WHEl2FlWBHoq0PuJ3bkYd3Ie77QhGETQ8BLgU+09dj5JF7/oqiGpH
Zr/XgnMnAmg5z/lWqsZVG4edpz8JPC1C0KBbHWLoYzAucLViAd9AQewVFviZkBuZufU0eusBWO1g
H3os7vhVO5A8Lrzd/Hu8EVAgedQlAV0MNEEL+etpEPd/LA6UXUXS0H0dCe9z/7lioADwrCxuAAdi
xgACYM2V+Si+ZyWWaTXcRwzZmBZHLndADs4bMjuD9hOeIeRqHtWWJddRaDvBC3HwihSsRDf7N5qK
hUairPINBVxKweTHwq/lbOpDNCPAGtsxxJpIUQi3zIIG1u1buxjNVCS0h+aFlKsCBRLv4W7RVgqs
B9RaPkKJpD8w4EdCic1S02egJErY7kGzJQAczJPBVTWm9i6JYevI327GtSWqvzW/RGVz3sHR73Gt
lh/r5pqVNSqiw6SsUr3wWrkuggo6ITutVLWQIfzRx6Pyghok4BXHCB0g5ybFtTromcXeUUXRKJfu
LnjRUwLhrvJg34CcpUHkEjRRe7HtAicpvr0dnzvl83RyQsakM5xGgdc7lUnVCNaSUo/ceKCPntFR
HE2si75KmnLulKinPbrB+het5cjapm5Yt53Z/n5uQwF2U503TBn6HIsrspfJwjrNIkqhX3rDN8rE
tUTRMhoHeGFdj7SeNQFoWYduKXPf1OwDyEyOfQ9lgYNKMH2b1JM35W70rRS5g29ulfhcRT1cO1dt
7RYrBv4zdWPvzO4WWIQ/1KCG/DUxtP8jQinVIN2GYdaG/CmAxCM1BY3MySBnjPSAISds11kEEhJW
C0EMRwk6wEqfhK9/v/vZexorKKZRnT+paXWy23phsiigfVBZc6ziznbj07fxGUkiw/1LDWCwytCg
8pwUuAEOFNdS6qdJyKEQDmY0VVWHocXt25A4mxmzySG1O4qTqUqvaB4C6AUVWaNXsqt3Y3BoUZMy
6nDSy5rcjFi4Xgd93rBM2My+Sd+URJ0IGyzmQpAH2hwxnX4HvxskVvjvuFdJSyYJYunCNX8Pw87N
1Qh9ICRSbXSv+op6gDJI8kfUhnnTXsHpyjl8LjnY79gT1thMx+XrugN7NN6rOasGezwWsjJTGp1e
ZNRODmmqcr88FqnwGCl2FNnwH7sPli8/DJn4BsCwDO1JRVT637KFEGC8mAstRDYlL/+SceO/onvW
NFdnJYZgBO8z8JeAGGXNKpiHuxvcVvkoEL6o+9pS2nwgEcduaHOVE495DEZTwexwBcQhNjN7Vy3R
rrTKZjrpxuKG7DYlO9sHTfBPrvQLMa1g2LVhKx3XR7++ncJ1HLQzap8Ga+4md7k/j6P3ZHbVu/xz
GZrYAUvjauFGAyQxEbqBFWbpGycHiWBy4wjCOzkLQAabIAoBNkjAUDbkfW3cPXrz17Vdf1caOyLD
uBgWEax0w6aAxbkbg3HA8xxyfjB+bqdJemDn612sBdQ4IxrZ/MjHoqVMC+NShIa35YgjELExkFOP
4R2SjYHSvihxJrBVhFWBF5DtZIEeuLEXgsus0XWppmntkLycjN2Eg/vDFHRtpGpz8hLf2wo7WxuF
PFeSXMYjmUqWCVXDoN2+71OXhOUbJ1A/0dhgKVfRFrAQoMXkeOoq+XbOOcVGvPmZQDthg2lH/PE6
XJAR0cFZYnaWATgV0Aee15Vxcv6WpVJWgc9EJb6AS1z98hSO2E8UcirHoksGVNNw4kz6Bw/sU6AE
Y8D1MDtuyQwiVNL/YyT3dYGUoz1RCPUWthuOHUfqZ4Uru5+H7bLfsy8y6NOw60BfrF/KpZNb5Aa1
qjM8oJTu8KLerkVBT50NGz+qdc3IfZIbu/H30nZ1usvIOSosEQuQw40aJpw1Nlh/8gI0No34UaSM
QXqHzGRN7zXEY/ttnabmowtMap0rx/OPnmTLdfOKTtVEQUD1Bu5JR2YLxBB9J+FebnyLqmV5wwoV
B5JJpFRy3XQtAzOwyt02upUBeEcdZKw29OtltSXdqQmSujGSKcca/rYfU/5hCynoflrctRg8pevD
7lnkCeS9hBF/2ouVOlJKPD6mR045p2Wp/j0v81kIZ+LAQ3XSfFuS3t6Lv6mGVQ1RXJ6W3DNTpkzI
oegQrbTMwicDShzbc595ZhpU+s+7jACz+wzLGiTc1hXAIvnQBgHnXnvfpW72yaccqzTpZlyNaXsC
lfre9QlgcnPycdEVGoBSj6yBie0VZppkNYo8zLlXFmH1phh0g5sdt5gtewBxQqKV2Ocx54mTwP+U
BicfRqgKLLKTcPbwScCIVsnuU5ts9ot31XHEbhg/rHKHCVsuULCS0TiINQO1sV/kNOFHLoLBtuHi
k8RNUUAXL3wu+VPjuqd5g08XmPsEx9MDhjVRcA9BM3kAXxE5rH/+ZRnlhqFlRgTAPuaGhLJkD5pp
t7N8eZflPypioCqOlRYmFcmWD8w+Sf1cf6C/g19ilDc4K6/tCEtWZe5yGHopiO+r5h0e5f1c8vSK
Hv3TD0Z6G1Zdr9dvHN1psJ+OEhyKkPJbRpE2UqXV17CFkJe6jnfwJc0yhqx/TuHO+NfPh9B9dEOZ
H26qP5UfrERcIYkMqO1mzKlp9ya+6koJyahl9QUitXjGcEfTnBRmA5zM3dB57GW0/4iykSbXNswq
3YCxl0rmoJLY95Gu6xt+Iu7rXLA8Pg62XDD3F1Gup8YF4ZTWc5QNTfKl9w29ZehTnGssDRDthkHb
qk8ZNBuKBkrStGaIDpt0MbuhfQ6qr31NhbniQ/ynCeN/ULQ8jLzCZqQyivFbSW0dllXIdlFY8Uxx
krI734AIHuMOvWpbfwC+eat5MEUf24qoFgALmeiri1QsxFeaYP5yDw3l8M6l0iWSh0KhVbiJUUtD
kN+nFXt3PwJtpzfge7ySvUWq5e3pi5/vRRyK8QoMo1S87h+y4etCF14SDASEHixP+O2hEGdeq6M8
/fK4cu67I5BvCLgofYDCrQ7M1wh/ZTMeD68zkkrq3wxJOYnkCUOIc/URqNfl9CFuELspsFt4VjeN
jS3kzmrpb3Fp4Xy1qmRMc/mVyqFUok+vDF3NTtGn36OTfcmsQnEUfKAGGpZ3D9PhKkrxE008gcDx
BuSUSMAerwjswZtGmog2I9PfsVoOX2dd3QaNt68sN9PMJn+sOxwzKLz+GTwGo9Uy7vJ6xTWYwvgS
gLhDzBHj17E2nMuT+EWfjK7yS7+3nKKTOfJ2BevUQ0B1nOZl37fv9SMwlG6AeMsMsYyDP9dYwf1l
O1QFs695v5pkes4qHEnXtSm2ImQbXXmyAF3V3Qg84JMSVrAY2MnP3xZz9onNfjLlbdn7unEiPrWT
kskxx+wNBzgWSCVt/OvhI6003EKjC4kMxl3YO+BBZ9CINvzd+8+G7sOG6ghXronYHlokxQpyvP6t
dOR56yli8RZ6PA5FEuMy2dlItLvWW7OhJw0HP+jqOgYwqHCZIe3UGIpPv1NLt3Vrc6YEYuErmXnP
NFf9sLIL7Ax6hPwo0f4ZsLNj02fA1JmL6nEzdMCYHsIwAm3eB3v1j4kwiPubWKBcs93wNapFUH+Z
4ogOmSbNEyj13P4ue1dJwh0Jzfk7uji5/tunrX4S5OpDf98MLal53BOT+/rJuiKJCFeJ60Arwb5g
rlTcpgTvq9GnCVE2ZDY2nis36r2HF09WSFG3ovd/BV+3fpTrIEuzS599vcLGMaybcQOohXxmDGdo
yEi1G0X4TmGsGyfY3G192Z1cZiYIcCrO8JV/wNHNmONaDb425ZRMcRuQkLH5ZztaYbC48wH/B0me
a1YXAIMNDa37IVEJiQr3UhOwjeEJU/Rr+hmo9OFIAs2G2HFbNGHEd80hBOIV2x1ewSNUL7qAzkMN
RggxqFLN0WXIbBNGP8Xv6/K/LOgomvR2Kh3w5tk4ylM6bXL32NbRTiQSUTdBtoJas6LaL1hwGuph
VKdHPVFaKVIoh7Vo3Gp3J0QrBRokz3uLt+U80vpx3g0HcV320r8sTJBT1KGgNHBzGEPImcmhxTAk
yLi8yRVF27/6Xti5x/Hk38Oyw+Y9A+RtVMvtfBkBVorjhWp1uqgMjZwR8X7bJ4ebsyiyX1EQ62sV
NGimdy8Zj1NOETGu0W1tQIDBU9SkvOO+sQEyPGkEDnyt4oNeU3nfOpCQhPh6jStfHyqYds6v++T5
eGuIO6o2wF4ORj74zSYYNzWWNT0iDGxz6EoijsDK7LsRo3EB7uls4jIIblQIW627LCcEEpID8ITK
9OdVkBAp/OnW6NDEXM9IW7VvGhFvg5G0UrcwrbR7H9YWkE0pZRvuBOb8PPuNROXf6eLneZxrMeQX
a3IqVg2ik4z2ABET82+LxAIE2ggo5T4zB2/krCd9wanbMKfaYT/GNHxD+f8dxmpMzw76qvE6XW8G
nV14T8lN4dgminkquV+/Y+PVYsSpGAwfUL8t35A06FReWtkaKBcsvQu94HR5SLYnlnmSNaFEpIbm
vwEpRpS2NFQzwSN6ymAQ4s6VfRolVOP2VwnAjlGEuPsw1EkPRJYxJPDSY7j96dakM8p5es9/SBmH
gMQ/RAAn/65ferIzykcxmxQ09v02mXiCOLdGYLkgwnN/gEBcmZ8Qmqeq1EuoGBgzYeRvXBQu9vQw
Uok/YLrKub72ewFegzJfZi1K7CHGLD0hMiaEzVFm3ZIRFF0jaR3hOCnxfadObxWFzN0jpjJoKusL
pp1Q9t7Ndj9DNEXKvVJO3KOX1iAQmUiSQGMYlbh+S7vcePojN/89QMOkHGV1faHJpQj2K8hGg2GK
wMkfaZBSSardRlc/z+VcVlk9uRlTiDsQ0gzNoEc9tGffLo2tzJfzVJ3H392KNkYeByV4hNA10Vf3
kGp3UAa941nSjPwf2ieU3yYhrRkT0kdWCSUe0f1C+R1Vj1r8ngvj0Q5ZdIR/kNSx+ODhw3E7dQJ+
wX5BIun7ZqX1sH2uzwhurlxc85jPIsFAfbODGDA8fCnVRFzNAqzb/8ArTKWeNvbyJVd8Cr+422t9
41T6CbmvwpTZSb0p98M6SBwSk+/s1DDzDYxOhg9ZT9vSVWA/8HoE0jFj4Nh9Uin5lnKnnWKgvFoT
RmAC34BheIPc1PScKUNua0zGPeuKyWyifX0nBwKe9kbg3QIVOfwIFevLCM1szEzntb6g/VNuECwr
E6IF2FUpNqCdtFOa17XoAOk7S2LIkbLPdRAvTrJ80b6lnExxM6MXJ8/pfKpyj3OBvA9mXqRgEQK7
ELsmTAG1DnC1grAGqZzeG6TtzmWojocKaFzUJuL7dnw1TWOBVJviJxHihpvDBptScuUqGQWR/qPy
irZREuBrQxapRF/PJftdU46/gpNctug+JRRJCwiG+ZiIDrMZWtpOnrM1N+jAQjqs6miRc0quTLmt
zHBfHwwXOs2AMMbMvOgkIVJMniexO3NDQfcSXat3kcXZTbO4tbydhxtuiHa5qby6ygi0I36IImBn
cBrtGYYN7znE/2Vw1e029XNx0lhetfgkYUgqdOSitdBmJ+9cpbPXQat6s3XG0M/7GI992UAuTTVU
ribhhi/4PuWUZSfFoMXnIKIZJ5/H7T2zN/YCboaDhZt09X/sjLbRywfa3KaKl69gzNTTpgcdxbA5
QTFom4mYTfrajxYFt4yws7xQvQ2EWyfO8MPqqGoVUJY2AmQvJzL43+VPvEkbPveC1Q8xWue5q2X9
JffqT2rmqHjwTXCugiDo4Y2Gnf35c6pMFgqpZ2fLbpckig3wIlEeOe4wVx3nef1/PzEuWdhNt1Fd
TwHP5oB1AWfB6mRdFrTUTeF9OXUqHuEKJIhfNibm6w0fHI+RK4LA5kzCtOBAdlBPp3gfybYXjI6j
g/e0ZK0I8cCBtue76Yd1qC2y4SIAvPTgDy9V+2ZtR7TgC6oNeO77fApTDWVaaOGVNfztjQ7/TyXt
yyDku42m2qQnzoSlmCeMgqif6DxE1GclJrUylhxheXTrzisOjKDeA2IcHJCogoTwX1KMRoQi/1Tt
UCNA9QgOEDAy61V5TQM1WcSDWMvXoFd1nPrVsd09H4TVnNbpXs4G0mxBhI1ELNEEaHN6BbkUebFs
02etgceYeai3lUOzaVjsa5xU/R1OotuNtuywiclF6UmxH6iJGCypefsFan2NknSzA4iz27eR3TzJ
gVJIyOPjc0+beZpNaZZhc+S30v88K7xy9NA0ewpT7GfVUSb42bcDsUbf/jnwxGAs1QTvwkts3tsM
lu4SdSbQAickWKZQuUCCQ0xz+aOffU0Ptdhq1z6fRdiiNtu29J4oTeTZg0Cndvn30Azj5Sk+4s3B
5GSTeRyt/XejL8OFlHaNoXBq/XVduRF4TIXozZMWkOzpzWnn10w23VWjo7vcWd8koyWl80xqEhLb
aqnUI3SvGu2U96Gs3G0Wp7v8er51LvL1Pc306exWoUGQdKFE477+AVlONvO9nffajFskCZcWpEJX
B9KjiQZc7RwvE01LUkgyLx6oJU/eSWND2ku3VN/l/ecsxe8gZcJ34VLkTlCmwSRUrXBdTEr7Aa2w
Iet0aWRglZKNm4pwFwwckq1nncTsv4pg7r6KtcBnS/hAnl+SfddtUycKl9Jj4MSgrctgwwhUIbI0
dMMukJLg6dKWl3p6+R3IH0fsf66v54wEGzUV5WpDiaNw9QXunxRjo0UUpmEYoIoelXnkh/OkUdjr
Tw4js7KOcq9tANw2ZQDC1EvfVq3V8oxrlUBfT1o8dFwIQ2tRLb2vJSoak6noWNza47xDMQPvjoam
RcAzuY7kya2qCyEVVASQKbMyW+VMYsPYx2N1NhebeV260i4iWmu+LZnUdCuVVevRHWc14iU9r1eF
mF4MrQ3YxHTrN5ugEa7euRDoKSq/+7/KnJBuE+AIa0gZGjCzajF9XDLlU2iyUpYpqucdcf25ShMu
/ZTo9JjkTitH2QFTlVGg77v58DQK4YTMAh5HJ8v6xH47Ur04dH3viRwm9AGoSIQFimJi7woRLmyj
KHXF6+KndNFsHtUs8Qyfem7VSgFQWHiqoxBH4zWPK9MSx6l6iQ9jSt3jPMPl8bjQMEc7AnFh3hJ/
qO025x9ZBaJE7R75I43TtJOoaplrSNmtkiV3REeHaSALXB9F6oMQyE2CR0lPvr9Zqgf/55LH89p9
sGhmU49rkJHMC4LMJEOvTT7d1IRmk76fS8DFg7tMtEzYRCBiRgIBfn4SurVrbjYjxrfVZwA5/eo3
Wvwch0i6TF1nSDyRVCmOMwgxww6P7xovxOHVLsmbYM43qPqdGoH/ErsvibFDcWzS/B+qbj3dKGDm
u/nwDYOuAjBjyqRSuGOv3hq9wYgSZ94uHTx3P4Q6t4SoPiwx8pqJCjJwwt5dmMdWGBfAoPwofj9n
6FiN7DpriRos07Do3zsnYYsi1ymUBOyPFKW7KWpaIUMDW8pt7NcEfE16IWuiKiR+gGeqcXN82wro
PB0hwY0uixnbtiBD4RBrjbwpOl/65lC00UaphGNyqQemIYWmN59CWZjJS9y5y6xMDSlTe1MgebdP
CpA56v9Q/NZ5IflnkNHeTHhXVIFLnSw86LSs++jshl+jhfOrCpfXuoYMDVqRVphowfktoABKkrV0
aisZzHsBdQYjAMD39Rsrsf0KiTKPWGaPNglhqCcLVN9fwmsawpw/eFami2fjkKCvmpajOnlkSIof
OnVAJqDtYsuVLNRMdvvlR0FJAXf8qncWl8NfM3nnDWQ3Uw8UYtN3qoclnvUFAkDQy+MSE/5Q86Az
mkEI9InoGJOfLwavdjT89KEaelFlP/0rhbEiHQDsu2aF65mfKI1L/6IaDDuacHDywbdel7Ee/ie2
lDJLFCTMmSvZOHGHhT3KwFXFD6h4Ow8b7nVjQDBW40Jcc7Bumudi+zI8WvUvbAqb3KYtUlPG761n
AnXcVG2Yk4cI26gJ5qx80dfMtsTCddEQnDqiaaby8jgBz9wGQK3TU+wQ12VmlEe/7lifFgr8US+u
MerlOkigjXzJ4mCcb1u/k2OPaeZloUdVsQ4uwSkW7PLV8ba7iMEZjQi9nQdlgN6Y22wfaPU3If+1
SAkqI4rR/60FGstdBbG99Z+hgckQNJGpgqyZUckgoKytDdNlwjaDb0g7a92h1vTxbgpYh2LNMIQ8
u4+x5ym7Rx72ZqI5GzYdgK5S3YEWYcVab6ALYqBg5Avv5nJcrefyuv9oBsJPdOEQhs/AhwK7nKO8
qe9u+blE+tWF+8QE8d40j8824wwARnaCzmEvWtKvmGsgRfsk9awT5fKb/yuuENpnGEXBYnV2LZXI
P3d/wFQTGc7HIIgZB6vGPdeNTQRd5uL1uDNQbD/M49/SQg/3mmDGCfjIkLwalYDrnjbHbcE7tQdx
PDGUGSCgJyv8E+1kTrxcfNcRN/5Sghr3ALtmZr0PZ9MS/V6XM1WcTti/KxJP/MrCJeuzAlP6qOqD
d38KDWO2Mas5dLFW2eh96S8zPRlYvp1dtWbdVj5avAv5J7sDFblgMC1JR2v05e6C1ZDHM9w0PesJ
qzpal4OYHmmeLYohBGndVTdHXxRSXKmAzF/VlSFzxGIUSo0zuxKW4kmJXehlXvM3AH7RTme+KrYS
O5x/Qg3I7Im+5zaucX5+pakOLJ9Pan4MnT0f5CEfR4bhkyx8Ty7SaxJKN3a6pHOwHnN5JYgKdUj+
iFTkW9sMmlMp67ADOwBrAfzGGY/5nE1UCX1uBJtUs9ODnzii3NwC6g+LiDOyasFFupIWu6F3/4Xq
sv1czyX9sGozpCT43ClZ99Iqv58cxieSm8Z5G82jm/osP/bKCOZwdiRPX9cz5WQtYMLOteCzhCpp
JTPem7xerT1kKE63JWtNAPnmKkEBDYyZIyZ7tQkjOYzS1QtHKgQlzQ+9b8YjhLcC5+O+GsejZ40o
q8Lkcd3ohr3sOoumJlTrX2m7OBvIlloevKB/qFHOuseE5iVhJelQHLPM68BYQJuxy+vsiHgneCEM
ZoWvyDW3kugEYyedO+ounPza0xny/HUSyyFR2954txro+KMDo2V2YVDMJ74gI9NIQ1GP7TaQahW8
tQIi58jD0F/mivcmhd98j4UVLI16Xl/Q8PQOp2VBS/agN6owTyvqyDUsNEjj6BvQ2PZAx2Bq6CKw
l9Hjf1Z2xvk0sL83mdRZqGpvPHEaosoYJZpm/SIYxXiI9RmZCJTT5adP7I7mteat46Aetty7Fhec
JBKMPQ0XhO9eJYKdPONbdEx3nYsBezpqp1ACfu/2RDQrjbsAVaNcLKqXA882wX9TDyQ/47PVxpgf
4hGAIKOi/D08lT/fjwTK4nm5tZd4oJ1AOuhnI2uTESmnkntxr9supRzbGtBNhOyj42aaE7WWFm25
4C3PmsWJ+NyNmOMMVUowxkK65j5YJhmVgY3fh/U4mN0+C8bxJUYe2OXfrsPivgi7ldDCRn3AqcFS
dwrlB4zPsNsVX++2cdGWQJlT241J0OPFR9f3wdqwmdqQiCKGN6lLtVh4JIBYQwI4ozmvIyfpo+0p
Q/dkAvI5oWq3LZZ+eN/ovxJl+kp5ACmhPNbI/8S/6Ms+XatFC/kMe5eG+h827zAG8pb4+Y7ZU4/v
CpEzH/+cc6TjxpUHNEF1lRkHdy60yJPAfXX9StE1RQdJefXhcdTj2xZ++ZvoUIGJXvp2HypxmQ5n
8uL7peoHDQ7Jliigxj1/T4If87aBKPOL5RIgyzFMEoa784AKGfczkYIZkSI7UCjHnxAEY51lh67R
vr5WWbU/ru+SuNFdLFNswT20bHRcymp6rzQUuuxdtaxQs48DWTyIwMVx2J24t9FxQg7z4TKWLbgo
APmh4Bj7uO9qjgy4CkDcGHFsK41HUDeOhMHKqIos7mMOcQJJp4dIJlKd6y5Gf5buL5FRRWnuT2qJ
trswVaNu0GVira3eMldGeTCrLrzFC1U/c6i5oo4M/goJLpe3vaT4GT87Mi6hlkBBigDPXlHBqNZs
O+DJKYyolVv8Vv+GwA0a9mu26I+YT6eFa/3Iz4UT9qFYgtMyl2KHoGpJ3f6JizBKqQy9jxLHN3s4
K/zrdMUMKErL1kpuPRRP3yoj8BO6YjIx04nsVjH+ppbUPToCV39zBejWo3Tzc+zIIdHA2MoW37Li
S0+mz8J/gKVNr2pHtHa+ymFkskJg+9JId3JAetmKV/4TV+/0XvJF1EpbE5VNh6GAVzIZ0Hi3Cn1w
JSihshC84bZGWlmatvkF1MkpVQtZBc5+E1VjssnKT8avGbl6fAlbzSZEQ6nYGgkDh+uqozsIvqrX
ss/JhP7OVKfQ4nw0eubyWexHlp4BGXncNDxTyR9No/urwnoad6pNtYEiSDe10nSpFOHzt2osmZKT
MpvujUk7c9Q34aKo1JIyZKFne4WWAs30q1J50enrUxux+yyTUSq1z7wA+OnepaZ8MUWMzbkNjmGZ
H674x8RUQEOWJYg0jzQj1Q6Se08XXQz2dTvKZHeofPf9YKoIIeuPki+g0LnOnkhmMmWDwrJVKXtr
5YRfYC0HxHQaP60IVdQsKkzAXBaLy7ITv8JHyfG3+qYhWWyuSiM+Xyj/CdzVLJ2bF15Xs5/KAmYC
/PAlEerjIj47+yaOMnCkN1YUDLRsb+Z47nENwf7FzFamo7RssXdeSvAQ90HA71xjhFbBJFNE2LDq
rpI22RFU6YY4gtjclsBjzNlfz65H1YSTMiTiDJRWbWDaYVrWwanogKrqERfgRK/CA1ZjUDVz842z
S5d+z1Kp7KDjTPJtzwRAru0R5uyB92UACnTqnWgLFt5fjWt55+wy8AkIMf3jgcGXoUILyObJDqRA
f6FwVfuXeNoTp6wKC6efBG2Jep0mBSNS2PgDsk3hoqDgh+jifTbQ9sE6Gj0zVoFNOXM3VCQ2LOVR
jUiZM0hcYZ3rvLX+9Uol3t/Ad5SuGcHYTloYJ74Zw4AzVJXBS3Q1jz6EsKe4/ISCbnCtdmx9Bhyd
Xr9OW+Z6RM9VcknaQPmgXVUrER+x+gdpS1thi/MLFCk4tj3z0eJuSTHFCqPFscu7E8ozpmISJEMS
DPvNiD8J/cT3E6sQ4DNhPiuzJLaEGEpXQGh4ky3gtz1+O6CyCgkGbXuNXumiEY1cleMtvzQZEWpk
AabUndqcDRQ3/lMVAKf3gHL7fM7gR9WuIj+Nuz8xXRpCd7EnxnEomQIpHcsPO376tHZWj6Ms84FR
hxbC54/Gzca2B8h1uK1Pk95GnKoQY22kXN8ahJXr7t6w0YlINSZsrqNNvtM7pNcvIu/CVLD15HLq
wGop2prVfWsRb6A9q1qwxPjDjgUoVYgXxVt3LLxNrPYyYweio01Jh1/qnv+uMkoQVmo1nqHxJYjc
HshM1gVaTTiUzVeTfIj+Pl4tp/nIv1qII9nMOG9Wl9biZd/MMQ7ZdFsD8wAdZy2+DVbX+Jw3F3zm
x1fQlRh4JN+KdmUMEbVeYew/jQdwk5jlmEN5U+8z60K+7VoXtYMMcqMUddLSf7T9WGT57oq4NZM8
4szpK4tUCoSEEOiZyRVgoj80itifl2b3UAYG9pzLmY256KTw+b9o38hcUjusc48rACS82c+9w209
B7rhxUnOYeuUdsHVudY/sVHFTRM2A9YW5h7v5twWcr/QRw/RLb/QDTYQxDR1m7eOEMUM74OiDzIy
AFVtVNrpxtb8HClPzEKSIuP1cqXMf7v6Ec7dxnUnBZMrQfP0vjp2UXyt++dittoIPELjfAiu5HFK
FUG7u7BQXqEe/rQNhTM6y5IZFBtix9Bz74GeQafW2urTAlGHKOvJP+jMhmShf8HLxqMTVGQxB8CG
5wHMFuJgOPsw7TMI1ikIUgu2q82lAZP4Nd0Eay++XSA3yU3P5NPVjh/n6Ccirv7fz4s2TntfDm5H
KbSnhYswjscMGa0WiX/Fs8yH4/i5IPRjnmuzYM/SHM5MinNBGIDP3lCDjbBndXv01bzcTAoM8cjj
4NEhLXptNjjeIxaXKCYf+cEaeKbsYR3SnvNFtXWE7u9ebU852+J2hHZYxspt/gMO1pcIVBnVieuT
JB2WFmzjWvbEdFinPAVkzDnlYH3N6anesKwtqQfN7lYPuOv+4stJ4M0K8H19qLa6YBGjUfH//Aqb
mjeScpjimBYVdhSJbSQ+d6VKnPbYp65icevEOO72qCk2onxezNpnZQ+av/4PiBgjFTCW07KZYZyL
1UTPRIThP0hon/l8+WuzIJMHgHvpSnBpMMf7iZZBT+L/bFkrV5jVTYN2hogsaFv7IkUHIEz1rveX
v5hT0MLwdP08mDyB4SFqRNrR9VDScCBnjYt8zwNwIrDQI+jWno9nKipKfOSy+x5L41v1pm67/BXn
R2/1q/9Qp7E6qIhPKnkRGsuZAapMi2hEB1UG0YZEsiOng5CtQ+TbpQKKcc54wHAV8Voyu+pIrF+A
AiDuYsBOEmbIfI/oFbOdiyV68IiKQkLEVAWJMdngrTjE9k6arMV6XYu9jsbK+akglnU75vf7wJ5z
bN5vlF7WeCdSEPbrPn8Mt+V395jtpzcJnpGi+ajNTrJfAPMY4euj8tc5hs4lmseuoL9Tm/vZxyRO
eXBm9PH1+5sDN6htdZaaJP5D4eX4w9Z/77p7ykcoQT89Vva7E35JiaMD+UYp7OpQ99SQz4GjX7Kx
jHrlvH60kV993q6W8MHH+1+El3erzWEkUsPeeTEx7CPU9UfUHVBKcIwkVI9dxJyxumnBeKkQOvCa
lcCFosSZd3rKfPPY0+mLgKQ3Oy/GWXNYziYSirHmpe9cbYID7N3Po9MVgod2BneaobyTZWfGTN0R
jFQmvGbY2eCBbt8+Jf/4fIQeJTfdWAHgg/DgLwU583/aUgN112Ln0GU/MFRvx+65fseTFPA1Lbp+
WOrgzqDb/XlkXq+3YC3SM1X8F1QevBIAY1KS1/Q7ddNrTHqAZoNP0w/CcwjZZ230cQFefRXfu3gy
R34RrB1nSU20nlMMw0BJUvaRD1+tXHBt5Z74TTTsQCMRpjM2lSMTOHfm4UShMkY3i2X6u28nExvT
D/mWt+dy+QXWL+3pGePrLqyMJlWgoHd5LpsK7WJzR6PzDpg5ClaX2m8oIVd1VNmRfx+go7YnvkAW
mzARIEr0w89tfwalY2rB5SNE0JNjfaVISUDB8nzHFMzjI0TiPBFKjWRqB3P+OzsbGA0BgZx5nM+p
pekJRuURS1rl4F+SURFl5ulTIHxsHsiSX0RaQTFvb/QAECyZioaLp+fNYrii+AiN/IjQOnR1Wsi4
eLfbF9DT/kkoJWLZWdiprziColJCK95an8RbMATkQwyq9gQr5kh64BYvWx/yaXMk/XgzvdXy32dp
/JqAW3u4BA2MxSY20zObxjfk00qd7KMwwfD2G2LgsYkx8Uk8FvsgyvnVwbORdrrKpqYeZyfJxMlk
NWRsE3AE9Du2N0biXffPATLTf0uWlPsKyufgZD9ZHTxsPkAuLZhlfmNxBBLm8Km4on652X2ac68+
AKRYBwnTzxXgNt5IUdIO8zSvjt7byuAH47D6WLZ3OD5V87sTkCu1gnBvBPEtiORZ4HqNk6hrztuz
3OrRHDXTYl+FhVfbQW87rJvWmOnJ23zdzbzFdOKAw8Sb03w5MlGCdjWzdqSmQlhbIJr+MECw1j17
7B5M+ia7LqbrwJCmtU6heyEATTqB71Ip0BLFixFKyRQ9VZtHIGnpCTee8AHDQsXXZIiCuTKK7cBH
7zt7Wkw4UH8MTlXW5P8ozRrly0xF7EKGZXOR8vnisSWzc2xaj70GnBIMQF6GhRbe0mhpoxJZcfbP
Jru0difybLi9H+E0Qi9fskfDXoHWfzCl9MMiUfIKu9LmPn67a8VvyYFbz4dK6GgCLkCVjrZty8KV
K6LrCAlkdbM0OaduBeCDCQ1iOb/6RMgWxMMptrzlXdQgjnvtpEMVum7bnpqijmdqvajO9U1NUiUs
RvlDfxhZwWB8eWiCiTkQW9npLrkWILKp+A9WMC2SH1hSjK5ax7of6StSR+ySgxz3vYKZemAQ8lyt
T9g/Q04qJW2EzxUnxFPeTk23EU6zlwd7oHHk7l47zUTsVpmn68U124zfr9BK9WzmwnldOabiZz8D
sAaH+91Z/QLS6ZTvS9XY70vAgOt77IT16k8OUfYGnEdxkHU9Hy7l+U84wttZlQVbeRnQpxymYdxO
IBBKpp301cLoXuWmgrsJdvss82miRVGiSOQ/7YyXvswB9lc3zgxJGjwvBoElZipch/G3HM9sxaTM
yC2VeQxXMgZgEiZZX/LrAaxnp14Cz/mECL8VzqyiQI2Mgy1Uq/hGE0V3EgF2AX9WmGcHRU1kq8sd
iJGsUmr2TWEzB0nsPcTXv0rp4+23qDou0daxoJbrItvGLB5OnIofwrX2sg0jh+Koa0EIqYa/sTJT
PdHNwcuEli4r7M1Vp6VtTfKkCZHP6egkSXYerDiZjR2LgsrbsZfSzwrpN4npgn3Drtk9qbCk5lJ0
C+LzeBEyxLxYNURFzXzGuq8anM8jzDO13TKMRchLrPKFHmvMV2eyWaaZJr32hw5ZBuC1c3eWzCyc
qbZgeEG+NWowNgy2jDW0HJoD7rpOwFaXgB2tINOv4Km3uiKBIdyvBjayoMrmXxP0ngmxEFOvLCBy
9vsSlwLG0pG48uTKAQD9VM27Ws+BY9uFy4mcjDvnsCk/2JT95ylBMMmvRAqQl7Xrf4PpDTcC7iog
ZxeeI+QaiBqvAyfxzcHO8PbmFAAPJRqTARtLzYt2685t1XReJ8oVLdsj0o46dQABZQzLImrH0lM/
Hc3OiErWI0YgC71mjj7MNjX++EiNb2UappiAXzyRroNA1ajoXg3KPbGKXISCpXgQ32zxCiI5YTI3
D5xumu4o8okSOnIiQBxnni2JADrlnnQMWbgDpsCD2m1GRdGJNbqDxO2QpfMAIegPWrvW9kgXlQB7
HkL6aRkI0bNLenXr0a4DwnE3k+HZWAzhK/a/Pn/S4KFb1J8TEKr5mHY7CGUcyhhMZL29jmgOwUJW
AjxNU6BGtZft+6JjKC7Yt/QehK/SK1dJ+gUEwptkA/ffStLXPZNIj/lmZ90bt7fvVnWzINAcJRqy
52HewjRHpbHn3+0P1ILJ5s3pnWDaTTtlMXKSKg+V1Xw/WGGXU2i64pNlS082PMzn8mdfwm3W8g6o
Y79AgE8tFnEfgOHI8Tcn+RbkgS0Dk7yP3gJiA+gUSv9uiksDs/BXCu5N0D9dZWIPwmgACSAp7X87
nhx6TEcfarOhGm6OWu6ym6WgjbtQNVy7Kf0wgg4zSz+iBWkNU8yNxjx++VFqITWsrJCBMWCsOnoh
85BXoWo6MgCNmApVNHpdPRcNs/bBJthiOHIh851ByQZgCwkBk8G2e2rY8svTH9MhlMRMWtOfyP2V
YTcFnUHlSWtxaeA/RTY2eb3am6FsJU4Lg0n36LiUuGxbnaGzniZDys6VGPS0YnDT9wPR9OAHsKtL
AKoyH0WES7ukr0re3WjrSWb0+JSXND181//DPk8Yy/yuk2udi79enPH4SPiaN3/rAq6wUoALz1LC
JK8oH/P7p8JRdik/BwHvBjScFvxJyxL9eM2Yo+AOcp/Alb02cuyg91xLdpH8PS7N+JY404aisjkP
s94qJLPcyuqyKLxx9Oh7BqXH8X7nXLcWFAiN0nq+Y2yYhNKXyEv4Fw347q5IDKUomCP4L/VVMVnw
ytNbUC0DZg0xf/UVePyacLRAoDGU/u1n3hjIs8GbRFNlezNx4Q74fQmyq3blcLQZZJm17K41mHnL
Mrt+pdnlnEZTaIvLP6fcXUzHdRuS7UhEibgv+CvBAg5phYgy4vWgkmwVuJGQcWULHdgsnZ9GAl+Z
J6M50WW83ofBCMYfFJskPKrWs1MAZ/P3ZDxtmfmqdEJR3VKLzMWjuXkAEQGwsEBUumYYT/3wabTr
quiGAgcQmw5jAY5BvMkX3IClJMUtotVVL9SCz14tWvzSk5SJswnOfV1qzKoCx9pkRIfHHW/NBNDj
ywzYq+FRtzDQ4WRl5oXwZNAARuB5fBS7X19l8yv1EjPAV9sHKqJRNSM9Evo9YCYm++S3r4qLDqC2
rh/Suc20656Zt+UXbTWFelUM2XfQY1kEq3AOIIMWP7hHbBbNHyy6jh+L2qJVXjYZD3iRjnkYPoYr
fxnfBBVS8dPlVuMEemqVh9VyHA/gKkzuV0hJI5Oa0WVqKgwLmx+8ee8VOYVV4Vt6Tx4Hj1wG7ps9
Bb1nePvI4XGUW1HyHEOuUV5yrBf9sBuOEokcl7dz9bXgq8UBgV6qAxZuBodAx/IiamMfrH/+AMzH
Ww3irQXDpwQ1LghEu9RrLsQ1xu5iSf9wxAlE6n12kQ0VQrlVGClJIK7bojg16NieXQ86vAprYsP0
EwF9OD/Y7T1LdZWWxhxm71Dmu8BYpOilYcGSbiMhmrnMCLdAhxIQTpSQuHRADtq+BNU4qjVUghk2
+vkDcFvBOR1J5Z98XxaXmmQNgPAy1GxQATub5dam+FQOcUPyP0DftzOjunKPV7Wzh1oC4u+FLK1x
L8tYlo4vd26kqGToOA/MRW8DJk2Hm5hafpeU8Kqb+/iwOSX2Zql5wpUAtmzb9FMD8pqjR/gFVqAg
hnzDtE2PY0LH3557uKmWWJQazBmcIIGohj9aLxk4BxtOkhpCcl9YIl+bF2cQ8f8Pp72RB6JpNKZZ
EDXNyqt24H1zqTrHgSSWDHcWbLI3E27+LRZ8BQWppjWpnhl7cIN1RCc6WIoGCiWD9EMPKAGi8KE3
pYXzbtvqDCv0PsMTSJ1pqbvM9EZOCo0aAy/yKJsc0is0neKGcxgNe7OX7JGb5ze7enW8ypYDr0F7
tGlkz8cg8Ypdd71pxl46U34zppY00TLE1dduc/k9aH4OuLs6+5qBAn6PtuTi9+5PlQX9C1hsioCz
flLPpSqhbC8EA1AUf9i4Ha9FfskIYao62IP21oSDgKlldCS568ILj1Oef4102VXNe0LXmLrk5JLS
4b9Xt3ltQnPJLG1oeYJ2iqtJYcbFcBRyHWneAZ2FEnQHvexoUyLcWnPeUcPRe5H5ceLGX6gTC9u4
90fjqNPP5N+1DCDIhD/Xv/0U6OI/8/+CU0PzcdYGwETxrSScjkaEmKrlS33LR5tb1BqWeEDCmo9e
Nmrfe1UryPP3XGNwgqGHJLfmN4H7IbHIImGFPBV6y5PUj8pz8ROUjv2l+Z7NBQu2EZaDYI1JMVJz
cNknIgBAso9ocwurHue9ApfFODsDL6GzO3bDrLazVNINqtWNBxuiKRvr+tK2XfkWnOdVYwYDPo0U
TKvnp5sirKv8cRKw+dCY8uNmpLiKph/QaIft69gEQ+8gpxVcVX75vRU9jNphBuPo2bRAiERqlSvN
6dEgpPocaZ3r2U4jK37PmExR+zDFuvPwGQw+XRYVS3ORaTFfSEZbOiXGFvWRSTHWnKFd2Uwf24Y5
kVFPkqIv6fmJ9Xk2nez4cnAPLCs/4IE6P6pJ3o8XfPAl9rWuhj6dGy+cphyTWZwRST6r5L1UtQR1
+GtEDnPVU8PoKA5kI/GaeXcFxOwfvG6nq8NPwbKQjhgGW0/XS1Y8tfg88MPyJFHgKf7kAf265r99
8ma28JvBaF6czqPmUvfHs020H30qvNEt6PoTedTPuHapT7GaIlpdCpD1MUnAE8HCJjY9Qwn0xYBG
WrL0iommG9Tga4j98MStr3UW/N6xsiLxEfsYQYJbO3yFJPf61J7kO7RgKN3IQJi1QriuIS5lkWKL
q3eF0B9kdL0bSyy+BCZMZJtcE10hWs2upXsu1nQSnu7hqJFOfyXTPDzch5qKhIS8/sIIt00jsikj
iuQsWJ0gysTcilq9TrV6A4yw5LQHB2HMnA1BBymSOtutJcBDe4I03dkuxt5ceG4MJQaMGLaRpk3u
Ub8zJKXc5eoXbWYxECA/JMAVjLzeinlzyLy8AN066UEMjRCd6Zm/mkO7Lx8do027zyoEqLxAOGyn
zD5aABSGl/xQooRw+Hjs8Q9eDKnQMc8226SkIeDtW7olQQHHljN8vEWphLdkiFJg115pl9w8EArK
r020mkcBjSWAFQfFMHh0U6/L0CfUPH6Yihkt30ueGpP0Pbd6RyklLp/RizAg0TuYMwlsstA3Liaf
X6eb+1rZd8fREuWr+IMtsCNNiZnPxOW1bkoQEEDH2kbaV6z6ChoSlS+0912+drYyJ5c2UDsBS7LQ
+cixMdyCtxq7oQ+wlOexI8zO7WVAZP31bwZwIa2uXHMoUMfXvaiTe/Srnq2wM/omb1h7jGOaYZYO
0z74fHLtFLY63BmYaVZll6IJe3OS5h974ZqhzS/4Su9SjusWVe/sFrF3D2Q/p7uoMqTJlBwDMToK
KMLg9AeWgGVyDhx5BrV2JaHheVe6xr7sVpn7/bYWWF/OrL+7T/xBzPHtCF6K5eZkDVCBOo/WaEzW
3gFGO7LAdvJUxdG8Rl63o40QTZCjvoghkUZFDR1c9BaEb1jiYAMfWLBJ4JQN84vmdWFfXMMEZ/lw
3ZrVaOSpHwmUFTQ3iRN4uqBoDkAfgBzsZwhRHtsrkIcTvpnplmca35rpeo39XXrJNKzNb9zfAHD0
ydpmtUWCWdFS2nckkTguVh4ippGGF2dhVGYS53+LgZPuMBNQGnJJSjWN9I2Ef/9AlCW6e8C8GTRO
niY7b7+ChMgtmUSWmjJQNBaHmWn4+IawIvB1c8ab75LM3QOSEnrOzVnEPJYBOtJN4Ap13yQ9nNHP
8xqYs09jQhNLrdPmekRGI9ThgbqJr8xkxdHaE44t6UBMhuQ4B8npZ96A5f91bZqY7SSNQ3L6/pcP
ZnCqcpYto2hudaxxvXV4IF7oxKb7q6caj1joaelRageNikifvcnXT/dxoPlrappVJRE7Ida25Nl/
SjjMptPUFc9uGaFlY/oLWOvG/Aamm/7OkxayULscI5TzAGcKIrgtoqMwc5dMe3qMC4wLfxQLA/f5
XJc1lu7wE9ZHKbC2PKC9lo3ddsMzX7ROoB7xObHeOc+AUNX0lMMHDjuXNXJc2wl3p1ErFqeSI5KP
pb5r2kXLtsDNActf+a7+xzXk0g/JO06Rg3nVbLwYynXetDt0p7p2gjLnrzQaU7fcWAStDj4l32QO
KgZcQEICzL29CI45lkJmz+3W9KJ6nL2BRT+rU0/caoC8imO2bs7acNNz5T32ta/lFVIi8408rvm9
b+/cuOgRxshB3s3yRC1vb0wT+sFZovmZ+VajmhEDId96We5tpSUsfkyBPCSOdxII2whkk/VNhnlq
frpYvKjomVuQDW5aTvhgYhC/SrftC/a4HijHlU0pyCeKOMKEo2R+WZ+KgUaKo3YZCnvcOrwhEi7m
rP5VU7mohyU0KteqNeMpIDSdwwSxiR/jgRRirHrQCAFKHtKawyfoDBcYTe6vaKrqbI0/9JHwsvyA
wI+iLy34147+vvFGGZch5DQ8oT46jV23EetB5H/6wcrnIhdArOFJG+FFmyHfF2Q+M3eP7wgMxxmJ
Oa/XkSJeknnHF/NLx2V2V4sKnPlz5rHZri2RlmDODIXh0Id2N+T/4kZTSoOn0hFH7V6vJarVj4Aw
Nn+mX6aqaQMDG+tCwSDPeK7UHyES7FS0PgOxj0eFPK2myF0BI0RVCnGi2ECV/Mesox28fhpr9S/f
HWUuqTjr7IXcwTbJyaXu5sFu8DscU3AaZMaRIo2RtUTA/7BHjlp/0ghKn5F9pgMPOsLMlg/oMd8z
zaYE9sMQnAcj5F/i04zkPd4SEFJqejOwEV2KYJSvZfFlEPDRVJF6mhRdiZbuUrLO6K3/YteV6/P6
NaksT8nJZ8QmnIJlgVHXYDIiC0H/cDgHgMs1dbmwuOIgcW0fQWvT7y1JHbRPStqJrL4W+Zy6PgUT
/RMl1Hf7syRAFymtIOy/xersKmcfDIqqbhuu5x3fRPfqpduuCDY81xD2qAd3D545ApOzDRYPgDfF
9m6jIL5osC19u0cqwba654upDf/KIbd5wy6xEdVsNj5LjLpAUtINUwVD6sN5J1JNhtDKIVnY72De
d0OpgFAc2S3fZtpuWi8gScrr3ufGl6D0Nd/8D8Kev6UXT7qKvh4EXPYq87gCumUMRjXwP9H4MT4y
orhGQWq+9Mc4jxAxlcS5PZZVWqTYKFXLwtA4pRSCG2AB/reOQYB33TxpD3GRxTkNJD7k/xB23ytg
ZW6+25fzJ5TXXLkdT3nkTE/Jc+zS/xIZZD4XSkQBPJm5boNrHPSyzE/4To3DEU/PBuTxFpY8V4N5
FXcb+pRe0MTre85teYmQ69NSqPJvsGAM5ubJpRVY0aTHg+PvSVPOwHGuc6KQw4X7pKgX2lsYKkXg
qLFZse3WJhhnetOfum7ManSycL5rBPt9gKPqe7BWakneGsFlGD5XUcksr0S5YRRr/Gdz/0tt/h1u
59Kv8OAXkCag5xHUQB4Pal6JSNk3zUa0dOcUa96RlK82l+UyEtFDCUngfsfDDgmPGJqQsgOJpgPF
Medzyf0xzgucEeJ1aIbDL5nLR6WihW+iPssGTKdYF1Uh9dqqKpbmSA6GYdDO07mwyI4zkd/voIkL
BRHaZ2xnoqdb2y4yoeHRSA/KIBEJn2tOY8EvgeCDkU4W++LFOBERSeVSQucMbShFI2BXhRncQfND
x3i94tjTl3iJa45TlCMKNQZDIdnyR/73xXBl+5KSfupunj9XdXDsIr5J3+biKoghd6HWEevgEj7N
bp6Gr0kJ6NXz4x+w2UoGGG/Zfon60zXlxVSZiACZ8mULu1mPu9BeTlQ+qFaIUpySeWGxJTvnvnln
F1cQ9x70B9itZN0JQfUZ61mptQ2/OgsDpfot+INqq6uTFYTNFppu9Zlx++aIIbdhJIWuwk3hVljF
2wtgbOEOQFmxCiRl6ly2W8FNjbwrHgOGep4/tvDC1MbOftZU324nycnHlZPVt0U9M6BLlYQWdOUp
JHSWT2ftht4XZF7RU/0i3n84MN0Fn7ge/MV5O0a8EhukuMO2NQVocZn3YWXbVqSagGJ2zLq3H2X6
C6IyzB9/961SAmDGNEM5EV/VjcTXM428eMXRc4IIJsaaQSpucQflWBZcFKsrH4VcV7en+uNq90G7
o7izWFkvAGJEGmIjL2h+DYMc/w1y7WG73dei1BiLh6rBx3flJhQZ/u0607TgXW5sUW0s1BCDmFPh
EtSpQrkhBCUv2ziE358x2D7wSNehHUQdd1YDUo8xj1bUNfzIMjXkOm21hZYLnFfx3dJf52cGa7mB
zPqYb/XPX4VPyYRIXLZUsZLPcNW/cCjRFZZPNp3LxCXBmb9yY33SrsxBAgm5gPtFOW7CbpaCmuub
jlZ3X07/2Zle7ZOnuAqZoKUsy8c9od07MbbYIhmsQ8CaLlP4drzUMvh93eR7KwxGbsTjGfrClFbQ
0e3Dk83Jwmt6PM1L4lureSgwujoXCZXAL+6RSMWYLV+mD9+U91fCXU9OLaLwudriImo/rCAoU6vG
NKcUP4s1pfBOw6nSREuR6IyOY7GSZ5gSTBoUiEwE+pzY7uhSvIl3ik4okIVqvo0Apu0zMVoRyQwO
3PPg+0v87NCLSrD49u0ONueOM5X+SXIkZHEuklVrEbMtnB4PB3BZKFQZ1k89kLaYgmIfiMJtp6XJ
rxc/pOHgwmRZJCwsbGl+d6JQqrljP2VBP4ere2RJNH6Hop1AfzyJS+/CxCiZfNb/ohpGGP9nWubc
KHidw0vFsK7gi7vJd4XOrtUDsN3lEZLcdv2gDPgYF4Iv7kj8O7yEVv1m+gE7so8NGNT+xMNcUdex
dnO3NAylDQljTPQx6eiCs5XKO4dPb76iWqoFSJ74KqCCYVj/C8H7cVL8WRUplzp0r40ZAIkF/JFT
oflZhp/642L5AlI88YMRlyF5u//jSzL/Vo265gu5EOhQHOrH3+4qjw+VKrnIEUDuYL+kUwOD7+li
BgkohPuKoJ43qczBywg8FzOvR91b4rmuf3gb2wZLwNccmQxgBKGh3ZqNO0OEJLaBRZIk1IRvDJLV
G7UzCt5nNpuiHKwWgRf9YdumQ5ZipB++eQ3rM5GFB6Vcq8U2NmtdbPpDtBi284OFdcugeNMhpabW
awtkpgwaq28wUnDK1aQLEJx0GAWmxialfkx4Oi+Z3nEP5quqWEoXzID35Fq2HB+0mRnVY8gHrE4o
BxAyI0YWG+gfj8a4PRDVqbj8kzQBVWia+P7TTJcoBu6zafX1HstB1mvDLvlNieviLTLn+mT7Pm6I
nh2fTV1xD0kOAYoxm4+ogw76HA71dXuehuUFd+ZL40LrcTrHD4cL8Dqh1Kb+VX6Sk3Wq2ey+VDG2
uK0ZnYWtUxijUZctHY0wERt1NvAUe9bRdGYB5VyWWEfPBmbcMWf4JwblLlrQnTX8G+wT71MsDCIF
bjrkTXNDFwGZQ18r6HFvXPwwNcqicrg/zL5//FvkZQXpF88kje0tw3qAu53MvKDpCvLixw9jZRux
LinJHMFr4T76iNkFSSISXnzPxr8oDeISLqm1dEHxNEAb9ezytt2pb1inc4o9lRUFj6K2h1fAYgAa
ENlY4KhPCDCBU1FstCPOAFskmWddHDjV4hCa+TqoOpNrBoZhqPYUeo5Rs7TVGpDv0rEDjFACHE2t
PQLl+3DkPZHFPnz+BGfXtfQInBIn8iS64B0Skho3Hqg2WHxkQgc3CWC1+CUc4Zz5M3ly/bqqx/7j
CBDU32AGK4MWtXXTPOYEv7T6FrEGGWbu7fxRZTIV7XNs0Yv1DBn4LDF5KuZh93M7ELsZ2uHXoAYR
397/AUb34DWr3YITe3Er5XrEC4Z2vufGf5JcmLdMgeN64dQIPstQtAX5sf0mjY69izL1d2+b8yjn
vAg7R0FuzFzb7FMHjYC0DR8OY91r7s45AyENZbQac9gWFXMzWDJpSo/UGFx/H9ZrK2Uo7pwIxydh
ASTwUnH0pX3OCPZKAmjHdd/mybCZrnsXzBEVUp6pODedFk04Vnb0kMHLXklvPzOEb7jObFWTku/j
ITOAA2ulDvwDzCFQZG/AF3v9Wsw+PBckiDL0PmK7ywgZrMy2gQ2UT7AKpcAUv2QvLdHvuLgyCU3z
27eJJNaXXglYtEnoTkoiZFcL48NUiwov9ijZQToUt7by6N37o5ODyeXsEa7CUUY8gTem1tk7/BQL
u08QYwYGtOYjKOCanJNQ5+iBiIKOb7iAS+m9J/WRUffv6IvmzxaCQPXqrlVGZZwWDqyLHOmKr9bX
XvXqQflemzgTl5X32Fgk4LG0P3Ai96/H7mQVdWXAjOlwQ/Ghg+wOIk+c9cbaW0Yct1YimxfL3QwO
F+jsctpajddm6++AgsqS9sDk8gi5Y+Ul2I5PbK7Ur5fkMMLEdLHMPeUcB5g3IyKa7DAuQD1OiCF6
xwLLhe4iawA+cxGRFYr+tJWiBhieKUneaajx3Aptwl7EE16/Ojw70D52FdaIC2XFGVX1TJNn4bzo
tqu4mtHG4mPze8Sd0r2umZE/yWq99Ev+ova2DjxgmNP1tyJHUL3rMyrKx01jdhcHE8tVV5d/36KW
Yw40tIPT4zIAIwyDgGJW5dIa2GoLZHKyQ+J34L5+NJSmlZgSKFBB3hinfMl1s9F+JlJyUKHPffvH
u1+C/drYV8mR0m/YOtO8p0VK0c2uMh4RjGxpTGDftQ467HjR8f++A1DyJ12poxuyZ0uVUoQqPa06
au7AeyJt7KEAEyDYr+FRb3mHjl/OsrYoWBFHjJMr4GRa+omG/VwYyCAdaWtAvyceyzEQGQb52R4x
MPC7pbsO1p/fGLTDuWcHGcNLj03+lzNivxpUyavJg/kyKy4XkYnuFJMtMewDIo0YV+fC6GL2ArMO
gRN3rrRe5X1VgssklC/AEcdyImZUxMys42nFBdhJMlVhUkVMsqOBe9d+Wzym+trVgqCohtSi3lpB
qSTq3wIWUncd5/Ly5LcpmJtqV9dUua8M4VbcF/dvn7fEaK7uaA8rC+k2lAmkGytfAZ5TK25/zOu8
sc+rldKpj1sIUTovW9s1X1IBm5k8iR0DIatPVib7Yk/mZi5tLGAM3fHpln88S1OURW7xglA79B6x
EN2i/eUNr5lhuBTstQD9Upmgl15QrZpF7FW7ZMU7wPN6WNud6WeL0TwK/GP2DwHBXmd7aJxgEyh1
a952U/BdKH+4y35k33/UFmTJtZLbm2dPzacFYzCyKereMAag0wGCFbP+dquLMNIGkMnmtRNVLqCh
0FtrSIHmrQi9kSkX1Ae7GMHIQxTrx6taX6IZ+fi3Yqln64RFDpwxmXPoQbqcmWBUCJLylhkDw7UY
kOHWRk9QAj23U928OnMw85ZfgM699OEs0+dodv2kLioa3N32xVEtzba91q5glMK5CxT4/930yGfX
/ly9PLvZkIwPlwmbFgdtBcGTGid5iwo8WMjXr80D4StGKdcy0/lDLEh+R9jo/lrZid4pTh05lPGm
fqd15JWZ667xyqXuuiEYP9qFxsBlDmz3748AvpIKLggRdLtovDQdttInJS5/2vzUAyVHlCIXkFv3
iOLf2+DxYds1joihAcKC7N+RYrUI3BSCPgLh5FHITSfxe/5qogCvP87WF0+7TA5t83mxEjHuYYU2
2tl6BtDtgBmiuxZ6U74dUBEoxXoTvBovHD3/CNviw0oriEEBpRIJyCk7EG+1TrwDBtNDgtzARw5T
Hq3lwPHFjXtA59I2uLo1J0tv6ZaJ7Z5iktJFx6uvHTDhKvqPTl4XySwM84+ZKITJ9d1/8av8jggD
LUya/Px7kYgYZWCBlNGEYbDv62ZhB7cTdZ60xkABcrj2b1LIgcQF2o1Xcfq5c/uuJIYEsie3n1fy
tlwwitu3bCfSJc67ELTAdQV7ErnilHM5X+CLw31JVCPf+vvrblgPJfiGzoL9I0sFJpKhwcGwdClV
zLc0kaRHvrQvj84vDPoQb2xR8KEc2XbV8GB2RMDevZlUbIvBD9v1V9H+eZYsKrOps74QrjAZlXWJ
cpnSAxmn9oWkQVh/lWnEky8oAaPxWfk+naahEef3oYUeXwU4aKPBV/bixw9tItlmR00DltUG+3/q
StkXkLhfbqHDBDEV3CWKSJxJOFqpP045q8pfoMnEfr+J9o9bdKcobJ74nGfNkyjjPMjQde+f0Mfy
xlXWa3gZQ505wXXIxfZMf+6RgtW3b5F2dBLoooyE1jtTe3MzMlbkmtbM8ImVJNN+rXIpz+FZIXAq
N3KY4nTkciZhbD4tUxAFYfdqC/LijyrIW+2Kve9BepfkKq3JjM7DGOmQwbAswXMbxdGawRESDcxb
tB/ACh+STwFrHgKkXj5i+2s7MPGHo0+nX5/WB2fsP+uUoWS0ertp8YFtI/90qhs3UwsCpVAdLId4
FPK8PB+UYzWPaffwnG8IJmrA1XpEqUetcyE2ntQVqcd1Spv2dC7AcUWeL73pyfjEBae0WJU47rIX
RTOlMupCVl42bptoXsx/KsWzCtRBzpQfZnEsGQ4N9U3++wn1iSQ6HwouploWomLYqXoIO7HsXFiB
I3WEP2JpEydcdOlQcXQs+5K5GW3o8DCzeu5/CrzrVdV6Ttf6jgs7ASo9crcX6t/P7mjDDPLM9kGB
+mxcICOI3akt9oF3kBo2I+g/LzXnxxnbpyVCPJ4cA24gHVCe2DS8/fMgB+rE1HjvhTLyGhqECLn+
j/VsEOXprxAaiAVQx0PYmO3PxLbCfEiO3iHursVBqSp4j5XF8Um2bh0bKMHU2m6kcgNp1X2cctWA
gci7mvnRGQLx9e8M5xmqiuMzwSKLppjAN8s1hHc70pc/S7ti34TpK0OyIzRH9WqLOEvY4B7t41QH
wN3ZDO12/GOyAUwdfguPFQWyvddGX8LWvzciRA9Sylo/bkNf0au9oV57l9nv6hEZXeGNQJqamFrh
FdtAJqaZDZCKblagGQl7lOka3easwR8T5R7QS5oNOeoNe/JH6vcV/9giH4ri4hwEd9ww/kjMfavu
m2o8asQChJtRMteSUcr5JvKXc3jP4PbJvkqCUxnHVonTXXn5qw1P9JbsdVMiEDVuQqZsJS9u0bLh
Vn+TgMb8mw9ZziazedYmzS3CpXfHohEYqsyFjhwfcdm0/oAUUgbfbsMh5W02t0fm68hacNxnLq4I
0/7/lQfuiHtH464Zvnmi7I8m8mrZHzOXssUHBNHOWhHOKhqHq2rVMFJHXRwwYFGiy+nrOas2bH+/
r0Y5qR5o0zncC3MhWjC0Iq5cqVNDj+2gmVju5UF80GNcjGMRPa3uBzEars36SVUeaN0at5eTCPZR
mZoO3maZS5dqZcMOh/Vjl4SyrQemML4Ju21OWqhNKDKtrGZZZE48tMgOkvl2obFUdynA0y4GTd/0
b5rEeaBWJs+VNVPbYKgc70TdoKc6BwAqQ0UH0Rv3yZBNMbzKSiQUgB3fqFvx0KNojttizipw8aD8
Meh8U7nhgDI9rqRFc0my5qncy3lrqhU/sU4yxOP8zl7LQ1PDtvUKjPlQyT8d/lp1w4TY0PuisQr/
babzVldjkhjr+Zw/CNHJZbfib5bzqfsCgfmv+FDKV8IZKGjSy1KJHvm7jRJjQ6qYuMJY9nuKnesn
VKuImyKT+MNInbsON39KPMBjT0XBc80p3ULzkUjeQ3B22+QPzdiyyAjBLwJz/gSHFX/wI0t0kYs4
Ht8MY0ksXuF8CLsz3NbosUemXfyEam4K6E/b8sBhohJba+oQ54AMCyoU4gPcJbi/VUEr2mxrSMBh
cU+NcoKinRIBLEdWbMX2cwW7C4rCEunK+yVu/WZ8ZSchk4FaZkr+WMtQUzR/taKmkL8I3TBTecgj
jMbHIqJuD25h6Nq69d8wZx8DtVv0Kmuvt2WuKyPHOG3g07bhW1M5MMXKf/t1RPbUFaSMDDSlhukl
yvClkKiPY0OH9De7VMRQgqGdQHV2GiLZOLTm65H07zN7cxajbP7v1wtA6hT7fm8Hh5q8SNkOSWTI
KU/5k5rni9TSn05MqZY0UJSruEFMtiiCptBEDO8sMyigBnHoIuFCALCq3z9AhvCwxFG7m/h3TIkr
b4NXOhrJRtkHGkp+zxv09QXYN7sBng+d9GaCNDfJA+wqeAwfI7/ptTcimwYd9c57Lkj1Y+Sgt0jg
29FfTSeHsqrPC/rk9mpnmCmZRhoEq9PwydIOhC29gHjUV39ryGPzMO5bBNlmRGRmYh/ziKuUc364
j+w3xoNEXBtFrZj1wrIhlARt0mBLaqMUhsiUolGkJR3KjnI+e1XFvdJr1GUgjLDCEWJDqv9LYYhD
Yn2c4GZYS8uinvRjKBCWScxR1BZNzOhe9ERfuW3SbBSh40KVL4T9XuNVyd7ZxNAKVeDYch1Kwacu
Px+FnekIqwGq9sXHOWYRDG9ReijozKUccMES3RgFj9VpQDmVCfrBS1WZWoDsoVA14z+JFUxEyjqn
xasF1ac46uR0I1a/Rza/H8c2xAt8DmJ5QPNrK/D/NPFuJfyXT37bqxnhmwA3SEHgWK5aiOwrrdzL
B6VIXE6orhc74q7d4uCKQHm/alxmlbml4ZPTzSHrrgTPiGE/32PPm2CJ31fq5LXFCpj1GPuMTBWy
Utvr9nnOKZTsVwtVE5KXuXI91JNl4vODdvNDjTyfpRt8siIPQOOV9//Fgfy4qqDHoFZ1gFiXMZcQ
znqUov0rn9q64ntU4CHYOnKyp45HeT1lmbjqBltCj8JJjsO8ODzVT/LXcoBeGtqJ5hYd6t79hj8i
ZWxpcOz30fARJG7Udn5rsXFNO7vmZg5w5kyKubS/fyDC0UbVmoWha+CXpcU8MKut3vw4IJlEHPmc
/cdwJaF7i79YgSIU2D+RUsmwfGv8FGUeF8KflqWlYG6Ymg6Ljgd/iLt+GaNcJHHSO+x0d5Zs+9+4
iYZIrq93gpUT2/ET6wHF14iSQhQmCX5Cskrv1eA/h1AW2blnV0Hx3v9TyNBeYxyPxkZraknR0QIA
u+iM2zbhKtmnTYVy8I/dw4TQnMg11W0p/7S5uZQkq+pM0w9bp9Sz6UBIZTxi1H3EPBqpJh1oKn4J
L4+sd70JLsY5MD+IUsJDwHiNUh+53EhE4wUWZTfZ8RladXPm2GjzR49vKdqbCxGB3Q/7H0RNhruy
ZxurGin+ynxnMRJTH7fB9975YUX6Qot7JKQaYsr62QU9cUq+3HbPc5V7uZFkGhGm+7A1AdHYYT8e
LLQAJQlzx84sTHjw5XrkoIhH6WSZ8suEtLgKd//bFKjFfrrf/She9fgOScSy8N12P+a5g10J0UxO
leyBpYbLI4ZkcT3Uwko+ctmTF++6FYXs34JLx8lUJYW0Z5P4gsC+cAAGuquMbaHNu/CFj4SWvFRz
Zpb7kbqAn1cYnGdDd0nUKAnLTwbZmtGF/alI+2cAW4Lw0OZvpLqBuSdmVHcD1C86zm9CAI87YljA
jNww/6Wft3gYx8fOFlNET6DrlDHzfEeumedRWQ2fKTnhg7CVfhnOdW9nyDYqe/saPR5/bnWRbYjj
P3fMKuA+Yps28GJHd0ket0CmlgZrZLQPP3SsRyhAb/1SaMBO9240gLb6fx0U9JPStKLg1vufn+9J
sfdaNY4jJnkOVdauGREhDwDT78T3Ywb/GBA3ENWQw5Fbij8SD72hZoliZ4Ladw1/W3OSp/GCyTDH
2QtgMR0NqTX8ouPmWNRWfUrFvJkDb/lCEt3xtAQXDDN3aexxyO3NbnWIHgV8dAZc1Y4+Ic7etNqD
R22rGOYQ7ll5CQptxATnmiWTiDZzM03ayOreIOSJP4ss6fVRgqzj+x/C+pxir/lGA43T97J1AUGr
dJ0wvDxNKJbrN1OzqUTmXyZfD+zysMNTOdIjThkmCOXtj9o0GXJRuexxtRXMjsexsWUFvz2dLAIR
xPddnamnsYqY5S07MTh1c30KUXWvvjMyigTQP1BffhXxlQJnZECWK03LOaM+N7sCwvmFi5ubpJ6N
uIJttk3b3daNaKP0iHSKV5yWztErTZilyYgagYkxNuUuYUE5hI7jseVtf385asE6TDeU1MtSqf10
OlGslSEem2oMxGpFDfmDMtUIeh18838guEeKefCS4BOx2AExBFtg4kN2xwrteGNoriQddIl9IY4F
136XbIH8Vg29DQMIvtUhA4Uy2z4dZwoQ0XymfZtDAhIA7jQ9SXr0WD2e0Y5RX4cdwmWtjC5Q+etY
IYpeFQP0nEbHs7OJ/PL37JEifZ0Q3nXWUhL4I+THL7kbbWe7yiimLCtlIcuiO1//RCiYAlCfBhOh
SVxhJVJqc3qwz9nHMlK6wH4NyldMSSLpeCQIErX02pU24zECjD4+iTcrI+Lc5czExgUWu19yx+xm
ITWJSOrxJLkrRbNvOu/j6MgFDcw57enAHKlOHyebZo1bkFkf/eVHfxo0C47cduV5MnbDMhglEHch
lZt0/zGYCVyX5Z9xnZCjvJ3mfF921m1GWnylrHc3R+K5T+x0aXRewf7gMMZY9zdzSt7VqTQEPDtX
5DOJM7plaLPH+L6jCEMuqEVR/rVSPVFePF9lRcd+dkK1pizT0bF/6ShayVeDveLq4TBnFP2VIg6f
MVHMvxyK6ig/dlTR/uOnnm3x7SNfvsIVEcFgRq2u8hRQZdupgS90bLkaj2PxKad6fDrf42PDVsM3
dqEELSa3vF57XFN3GjF9b838NVNCJdB7zvqcIn6ZqXB8beyxbEbDybvSL2ZfZeqkC6T4ZNrdz+JC
hInKWPaI/HnFSTkJ3UsswIg2wIm4Wwi0TBvi1YjOCU4ja4s7cRe/y7+FxHd7rgfo11gS8eQocFZB
k7d6IQwj+Z0LyIilrhtahUM5M+pNlMEQwUt978ZLXQt/WtKfH2eeP8cKENstJofWUlaISZvAcI5i
i1pwMosg9SHyrGIpLO0KLB2LfO+nGfya3bj8Dgo9k4oL+H5WUGBF1qpWPM5XjUbWss+1TOhMU/kU
cmM2kch6NqtnSntaYRGF+7DqdnEBKaLtErbgfm4prfkT0rlR7paggPP/hIazNEA5IADWNB25bK+/
sEB5lVA5rbNaIPcYFLS77y8C3iqkzZJ9shMS2vVmbxv9OR1goKYM4127iFskWJVpOq4iuAjqQqGL
iXPcS5kotPL5AwioVPw16qNM3Qw6Vj+FFVM/3ZSWtGSIsnPlZ8ihnR57/+MCfW6CJoDblhEu9nxB
NSJBhPN7pf2LGFwQ7UDdzoj1k4ETtcRTpTpbCAh5qWbAA4Rti2xijCTOyPB2lQxJdIhj3LwqQKaA
uOpzc/CDCf/nONeUrI3+XsB8Qgnqp4fswsF7hIbIvG9enuoNPkVPR9aUtinGHqgire9glesmel8C
kCrtKe+eSRYwtdq8wzCcJSekxacJk5wh+RK1JtykdNp3UnhvMDer3kV8qKs0vvjHUfBKsWyItz9z
GROejkoKHAxw3t7zZWZ5l9P64il8STRz1VzkH+IyUwIBBS60CpaTVDZP5bZBD/AjoogQWe/s7KsX
at7jeVeP6xUjcD3SneP35+kBAxJ8qr6Vck4O/9lV6kMp0GZCF9W0auCg4q+4EsWqSGbivDgw2lXK
DK2cfijmqh1bfHxecFzL5U5FD9FQe1kqqciKKbN0/R+d7892lVeE+XaQh15x7ifHrmuMljcrrqGX
2aIZFzOBCQHFd3NTiAGfrL2tZuZG1zh+bT2SQJv5ObNZ+0rpVuNvH4lSp2+gNWtuGYxWWuiCCT9w
BTWSfHPoYflykIwZy+eEhaJMWFX+yoTqzXliUEJS6iUbZ+fp5pqirV2rHxZ/U5H5uxkSLFjfrtnc
srDuqm2CQnHDJkFj92FhwWmjmROpBDu+Wn4KBn0RiPXloYOxiuVqpt6Pb6NWsueWUKDVtMn7QS3/
K36nn4CRVRj7hzcFYbfQknUyYeoZxadoeaavKanA6RW44Gh8kZftOWyQMX+1YDmKKvW1HwnnX0ZD
EgB3G3Yr/Ns/ltLi8dRYgYgCcicSvORZZJ/u4uBILHQ+PPLcPfOTtM3TvGxcb3oogqxgYBtAfZiq
YfZAA5xxbhtwwU9fOITDTetZoy3EvsodD2IsilI7gKI/LBIX0ehCee2b5GXn7Q1kJq9KHI+b2drG
ABEpZwaoVgkdLDKqWwAmhqvNVfx8WfDq0t2HSSYZgmN5m3djtwPHnwwVmUpoNPzJES2pPvIoO+H8
2T3isZyIr+Whzmy++fzVPEQsO1/Mc1/aY3lsm/bGeeP4N6jTSXgTChtYsjAaf1qF6GH4363dcU1S
hdG7aqhCKnwfzqYCq/8s4UEfhswiimQ3eW+v0MvrWipMiYpU4lBP7tsG5qmwcZF39BRW2fuOpzso
4/z/f+5InD7gLjjhLCMv9BY6iRbPoVMymJ4brJihxxQe99kOiHxn/MztncOqadwqpR7nZe1Pg+OV
VO4yi4WopLd9enBLlTsDB2DEFsknJ55pigMu/L9wCmIE/Ti0JtnYmSXGFtwpV53VQpaVz6gVkIfL
Ujg0xsxG7481foMrbrks+gCIUBMmxXVBGYcOjJPqmckhGaRSgI0PalSQPtKXuNfpzeTKiW09UY4j
/nzjI5lTIRMiTsCiCKlnHb9keYgdvzeJJkUNHmAjy6P649xqmpGKsREtLdU5xs6rwBGV6mXnmQ0q
zr0sq5ns4D5Pk/qt7ZnR/EY2bQjShjQrEqAZ1WYMVBXyh4YXgQwTe3dx5dyjMzSI9InPgJKac9v5
oU9+4n0J302oc1YqBL9L0tb5xJ1b8v4/fjdJyncnfEJN/vDkW30NIG8IBDO7xWJqyrVQYDKJBgak
RvcBc44BwRGsRpumKOf469TsJCy3r6VPeSypYKFJHttgWyy8gFrdbaZe7JBfOlxhkVf9S4zUOOpO
kPtkBY2uO+jwluFxysdGZORi0vGKTjesUk2fuPm0CIwHJhqUFMt18QqkQ+A1ztk2hWYGaMxUAHOw
aAbhrJVLijha/+PgZCp0ul1YgKWByyVRO094M3aAuiuNgq4meLGRibgF8Y4i2OvDxNSZAV2yFdn2
invx0EX671fY75X+/BbmVEMydRhRGaFZVEdJqRt8tCnySfa2lma5NiO3Q++yaechVorEvyLXPMjf
F8hxL8L0zrC1lo5ta8fcl5SaI9C+dSUw6ODNL35vK4MTymGPhKH2YICV1vEvTQhiGDI6xAoV/JeN
VZ018h27nV1mDGp4dIb8Yel9AEQCOBQb+6aNe2DvXPR6hITB8QVpIIG98F9nd+IZbnBU6ZL6IBNb
/S7Yvr6w+EZt7DePMUcDXsJdDpTy4ijCI8D5pLiHpJ1A7qJSNNAIIxaZHRGBrd4qEBp1RA5zEPhk
Tkzreg5h2usoWcKikUpAH4Ve/U0PEtBRZmxm/YllZeLoXcJlsuHLaYVuP7XVebWB6WR6gFbbvK/i
stM2ut99qKOnZsI7HVBx9hlZJiqAUf9jC/+8yuqWpxnilwEaY1EIgvXBYiBfLYjLhVPPCqcAlpz6
pYmWpMaYFlBk35MoovcEcxLeoJKIPJSLHDdW6JmH+bLnMPODW7i3XPaaT7/2HwRH6dJCKQrAA9dY
6goVAdXMam7Io6WawL3vuNuMcfeY7R52rjbsexLXOmLcGUgo51DLbSydyA9NtCY27jNnAi0BcCDF
sjm+pW3syrUKEN20l1/4rjLAgyfYOIFokCTLOjmpTvONWUwB28JBjjoxUkjrVBnzwSiL6l6PZS1d
CS+4fSRRL0nwQMraZVyPOcPvhTnZ2JZ4uKnOkhnNEUHDPujda80ppVKTpVMI88Pn1MDHH3o4JUst
A7KpXD4ciRga25er81t/n1kNaV3Sl3MeoGeokGez0i4GoPfYjlJZ09Wz3f74KqrpLKwVJkkWBTEy
VpJwVt5EafXbFARSVv4HouHVOXs97uEd8D7r5fUf51IllzruOVhK9n9Tk8Ax2HWZacLGaH0jMIlM
pxM40UlqEJR7W65hGmHp4JJhvKnjuLjENU6XqKm9XJckslkYUgmeJRS08nDFYcMX9/ktPs0JUeen
+HSwFJE9xjric5LrJmm3FGpeCcShvxLrvr17eJB3aKdqjQTnbUChbknAu9rZTr7AVNuBYN6VvTyb
sHLFgIkjD/c3L7uXpofXQkT7e1YwqgZPIhX7KTEaVuY7HqQ7vjsWPYjeVkvBiV3G9aF9UnTg5gkB
Ne0Roz67wH5LHmDOjAgx17hQ4MMOspzhJ29i566ujHAaG1w12Bhth7ECipZFPWZX4Lm7ilCZ8+u9
swChaqhmnYSJlEsJzb9rU0XmFv+EZMqi1ENzllvz/7PrMc+atpyOFGCW6zVuoCjFAinUIAlDFXBG
4BsA5UBUwY0c0hzhn97duDt0Ybq8sNWTbX0Vz9H+N8UZwXvf/sbpHD+i51/AFuQ/DSVU8+BO8WeA
iKZBQdosLh/fz0QvV0epHLbP/XNggOhtG6uccHo3wA0AZQ0r3jcE35I0+S1dqDGEdAWu0xPpmQQu
ENaL0At4tEMVfbz85FL3CjMmQ3f5K70nFtZ+Qmd0EKPurV9TBQBDNXfBjaqstL60dAC+YDM0aa0U
cT5gk4hk7jLbp7VDNtdnAUc6DM6WhI24MgjQeqQ/EL3d7CQNbbs4iixB2Raqr50+/J9Hs0TMg+FF
PHbeyZ0/tS2eEDgU7cDwx7GKmqnQwGeyMEDbX7qCwr8xAe7dQMbh5+Bxa/9XaswhdgRZNsrI/E49
boCSq37a7Rr9I892o4r4IGB6RB0I2HrAellQvl3FbafK7s3hKlft8kOujWQFcFc+8u3S46mvBWKm
RiuFF/RJhPRM4CvzotV+f8ol03yf6Tmt4Lla87P6/YOz2pyG/9KlDFFLFRfk4DkW1SLDJtaJj64n
qUQd9by05IbMUsxAsFi4W0STrgXYu3bu8eV4l+7soQVG0oq0MVP6ecIcRRGaTuZ65v8jgIj3nucy
lIDo8qgxzBEu4S5O1KMEQls1rSNt/hG47XSyN1jqEsMvB9mW+URlzb0qf/ARDepQNIxzgNBYnti7
baVNz8txoTFg5f4gGoxr+ySo1y8Vdfzy4Qt95AOcp2qV7c7p33eHveVtH0ygi8aKSF5Ijods/j9f
myGjYyfbBmwEIyojk8HNHQERGWJhjVS7PXV5rp5yfEVyavBikj04511cAC8BgOJUhXssrERbVHBL
DNuKiI7OMrGH8Vho9oKRnGQ7FAVJlDcx49Sj9Of+ZamwavBczhl0XyP+F29Grfix0YPHO4ZZ4XtQ
Ap2E5CZL8I4Ak92bUZJgz69D/Tz9XrkJBPlsMoa/QK7Qt7aME1/It5o9M8F7Jwdx7pBJHvoXT+Or
BOojyLUamP/LdgyKnI4/r4DWpYndWC8rfR1w/JAe3cHvO6TV5LaGMn9Mye0WP2g23btcKuWerIFj
5JBnSax+RNyz0d8HYsNNthBcLkiZcVPNOoAX9jU2qNRrT0+mVA4oxmg6POiIkFnBttA6Aj5uTgsQ
UJR8vgGnFI2u37dLD4ECXSQiqPdUxW5kWJ7Oms+oODbB8IYvovynav6WXbuz9G56+7J1FIzoaBHg
5DNHl/WmtbYNduLw0aUWf77V8TOnVIbI1689m0vRuxvi7GOwRteGIqyoS0MVxV8CMAo2C7IvSSTW
nq5u8q+sAEUZ0fcz/5GL4OEm2Zqde7LbIyUPF2ol13zyD6eym4IEC+UNKei9D75rNknlH7LKPDYh
tJiCS3hlxdpiZhJbeUkHBeQo/pOUN9gawWlxqyC2lugyDxhK2l0Famz+7oq4vACr6RJtsHlsU+87
u3ZLvMaiWSOpLSrepuha8lVpoBa2wf7cY1E3QVJ5X0MClf43zH6+VGiV5H2q6typjC1iTixakLKZ
nJ2CScqlobJc5rUHIR4NdroHf+pbmwQVJx6Jd+EH9uHW6AsRe+2SlvkBaiiQYyOSlkuqX9bcBXxC
RBGd52yQHIZFiZZfA/HvjI17QrtiZSGMZC7Gp6+I1QKoLbEHr6MtwV9/0R+ek/z9jf9wgoZ58bNQ
EHwKh8RZpscMHCwyEeU6RlcL+xy2HlbmKLcJbRcmbnroYheDjndJfCom0Nen2zDbLmCx6POtQU0n
eqrvgHMp8GkplCTONvO0HpF6Tz27RcCTv27BOiluF/WFPlzO++zkWmiRh4Y61p9Yw/xjLLGCZV3P
t491afw2eQrCFpaA84MVEZAyWBzOH/EGkiMzkrQCQmCv6nA6jhpzgmjdUOSS73jeFQNRALkJKBUY
X+wTPgUaYD+0PoRMuN4Ep90HwQBZ78zqJ/qOFklnaUu+77w+m9D47YbmI59YuwNbMw5PfQQroXKZ
PHqzdhp3oVd4gcEHfPg5EovSLH9SgXbZ4Ml/LSoW4YuqjrMKNBQ/9wELc00wkFsgbGHtNPxcfpPg
z2aXBhfRcj0QCNIJhMPSMkgCXaORfZWqZM40Lpt4Q++9WctpW5/F2em6o8EskaaSXLmcF3OyGG9e
mhqO7DpfGa+EmbQdR6crvOeaq1ei6Nj3Kp24qABNupJoOTixNz0ub6A9O6DtIUfl/wtQlxURsHrs
U+xOmWfFa7po98x9xDYjJ7yxyt+JTTptdPUaMs/jRvT88QbkwsQrJ/29PcnOsVGtq4INmuLLMGWk
QeKV3A25NTosHQQYgU9VSxtPxdFDrif0PKb1sQ9Y0tGQf/Ci9TzoHw35Xjf7YzeVIOPp+QhPHpxN
cQDb/Hn2JiASzQKrTuxTZCVk/FsqVuctApaCT5ED6XppRFuoxBeOwWl+EWz+BMS2HZPr/rmx5l7y
m0N4OHcwKCL7Uqc7oehdGEtobFjoS9yIcJ//1zlFEbpt2mCzNM+VvV2zDA/WMRre68kVIcLBzTqp
JtHOzhQBUl1yx1G3Ztczluf0xg/E8wAgZhNi6d6t4osW5dUxUuoIqxOJDrqycZSATqpHKmjbrHZ7
8ffmIfnWvhsIW8yys25CEIz40id8k9VZa3BDB+1v85ZAjPQHSqi2O67LyT7tyGoz9DYy4KmLJbrx
i1htmq19j6ACCdC41X3YNzwxaY6wSmYCs2J+o5vgd5sw1bNsjT+pi7pvPAYEM/VEdsjJYmwg1Dt/
j2Z2cazaVptnkI4jLhVh/Az5bNvJKC0G+R8hg6pb6ePMYpDlRxUWF/9bidOMwok6nCGln1mhEtR8
29EkVe4yQRmilhrcBB7LwivRxP48r/M+w17AxcoiputM2M9RqL4NsiEMQ9T5JnGBsbHga36VCUl/
Zzu0XuQJ29eGHM98y4IwUMHg+MNbszXU5UGjH2Q9BiCza8hbx/Gu4RLKGK+BmhNMkr9+u1ovBaoh
ZJFD4frwgd7T7y/AowZMjvJYzz2jAvDsf+UkO82tRZxDHh3VX0Wwlrryk1Dva6cktITCS+T4+W5d
JFA67rJvT7QP9mHIe15GQd7YKEkmf+Wj95FROj5DCF5FicTgX6ummhRtJ+b9bnU2rsjYpgrbBoC5
1prdd9GQPxLT5v/8nIDMYV6M9inrMs4jsnwouVFK8zHgOabAb9LeY8JB/m1BZyaJ1Z1kS/N5PMa8
kPgmb2HIR+TnHEGbR8U5GVIfwZTmU4AORPGBMYBRfaHEZKfCgNpKAAR2cSEZW5bQcOzwJwqqYTaE
jFmWgFppkP3HYBPOFnEsw2Mr1CXBHRqdfXul5MHKD0KxHreYKtDYIlg5lPRtIWndApOorhCM/hOE
tSBORk062etTCeOteSy3OW8HsxbQbGidNWDM3Jh1UaZrW9LHjt4Xd6XXU9lp67/g3R8H0rXfQISo
w0VYLCDX511YE/ZPIcm7oQN89KpRNGNtWeGPWbtHZEyLOBV8SJg6Et31zL77+Dub8Fj4x3V+8FeK
+DMb6hy8VyzPpvh54RUPGm+zH2c3B97zKY8dLDeRYkov2dnE319Ce74LxpttPBG+nf4ax/WIPWGH
qgcwTn54nMr0vinuSY/2W53fGjdknnWYyAe0ptlIqveJ0iMcJiQC7mVAygzyKojimQVwXYenZemi
FhuDAoUa66ebUq9bSrrJUPfN5U6jZSDzD2KJKOm5zUERQ7ZPrjGlGDv7ca9tAscNCGk8N5zwtBMc
/lhMyyXbl/fjZZvT3DEII1uo0EamCXSkntmYejd4GnqjA1DzCPmvRr9nZW4DGBegivftDzigzbJu
EkKdv0Lhi32sNDVIWdOkpqag5SH17CTyKpYcSL3zLDTILaihVkSx9YxJ6dZZdIsghDfegTVzbCxZ
V5vbHxV8zhNqyyX0ayXZuxp50TnsE/q/Kh0NQmv3518eul3BtQrgR1dLaKnrV6wuW9KWMGsvQ4x0
8P9JN+psp7eLUAS+SpOyldclUFi/GKzYZDHVuO8sk6I4FwCsHRTaI0JHuJeVJAXvPfJuXkv0owzI
ULHzR78EtBt4York/yCaQBtEmQVWkCsloVEkypPHuo+aOVw+tL9sOv5YX8zs3r+ze1FwPoVME3Gw
R/aUi3WtViqkX7Y2uwtrBRKh7z5d1APZEO3dIEnj+Ok+v44+Qu/Bj/QcPnV6ngGi3UgZGvzbSCqR
icQfINRJEtaoKB+SCMExCyTU8SnbkUhCpCJ/xeeI3iirxylcXMXK0Z2lJDTlFoIaRVolEFrhJ7A9
/O1MyeLWvYdTmU0OqOVUuctomv96hkyEaIyeSKC71C1BYEChoG/6l5OOifWaDMeVWIpG5GYTDoAl
4soBQf+2wzOhj91ROP0EabgtR/82WJHR0yvktcXNJEJSyZ4bBYhdatO/IqeIKxAPvMqiVsKCtJDa
qRmnptDuoGf/UNgdRyGewPKYMsMzyqClTAoh8KgrpazAYdWBfpeHK3sY5/wyvpm6DU/Bh7o/if8p
QW+VTEeZAv8JPFXnrFh/CAOlgWNpjR7EFgVoSTer+uyjedzr/2dy3svndf6MHNot59cs02jw5+fu
7O97Ej3C1NOqXSB6dN5qaihg6ExG33tU488MqH74xnwSbTQlxNjmbS5PbrgIM0DrmRxUZJOX1KH4
l4fIKArxABj+3ryxP9KxbMSGmqy3dWp710SeyI1I+f19fRUnpr15/vVfyM+kZN+8v6Q8vWD1tx21
dDakN941Ghr4aZZMpGZ30aaroh76rb3fppOsFV486IidP36oN16jZargY5g1EYO5X0JJhvTanKUY
VmdcwYBU6WvWZfIJ/CDB8LNoFiq8JGHKRZHuLa2oxvajy1P9T9YYWOsHmvcAvymUdd2bgGp6Xj/9
/BMuPJNGc5g/qiB+GpuV0Z2Y1zkNERybYqYjdGXEih/vEF/ARSm8yQg+n2b0AtB6ACwjWKtodyXJ
Q1jbJB8qWIDRZ6VCCpCNgJkA6Wc8lYtYpk82mUkATu6GsVZ0ERpsjPwC2Zu7Scf5Hl5BdcXbIYe1
UofYNCCZiVGFIDcJ1ArJ8M1q1J5Gv/5CISVyy3lDjWdoLMnV1uYTQm8E2Jm4k34VUmkDK84G+Y1c
mT/ivhf+T7es16bBqoG1iGrjfFuyZy2oTix0W+BB/K5EcobWqEz5VLTOlSgy9ubbulaW2Ncgrvc+
hkBRLWGpAji7b2x4Mj6H6v/lpLqkHa0e0DltyEO8lRH/CWMESoUAtyDfvLT6T2Up9XrxWcICI7qc
3LQ5zhemHN84VnqO3cVqUezL3mJDIoIz2v2EfHBK9x1tkiwQfuPuW9I6JrGVsm07baWx37DU+jrA
JnUJa72qb6kcZrAyy03j6kzD+2oEhP5nI/MD5aHv/LiD0NAmKLX2kKQwZV7zVnQ5lsYJm/irSiJF
TtEDarst1/nr7Ra/GN5QLTSqt5H/1EgQU1EuvT2GOiiDTAr667T7jQqYOM64M8pQ3TW6RY3jPCXx
znf/Mgr+o8wGjJKvUhcoZlDC32GLDxX8+f7oB09Cd09scPqRUfvHI+OzbcIrv3vVWnkINunsXd6F
7OIZPdZlUSsxfOh5IdGkiVxqIRnwX4CPoK87tSoIYNBgWyPYDFIHlU3XL5WMjimD+6+UCWRuppAT
iYj2Uc5nzpR6qH2NOP99zZ3EyRXYWO1Kq7tkNB3oWiOp7FI2zOMClaRUB+l0C5coK7EeUI41m8HK
ZADFjryjM14HQeJ0u5OHs3c9Tv2w8yxhXlBaRT5aDqSBALRoP+chkvPWyFjEkCWpEFG5eLud0bat
2mYgrt4jg1vCd+B5wNykFumYRb+mLZlku6nI962YHnTJRQY8mAPNAHtMarAnJkAxTeAYB3kbf2rg
NqcIMhYZXy1Kp2qMrs7/CDGdjVaVeQtsXfbBmNsTTVq0/zWXrc4X7TcS+zoUZbJ+VCvoyjnzNikO
za3WEeiEueATZSqvlaVk7zo4OK2fvirOqMdylDUROOz/YBhnKYC+fkYfx1owkDPEQTj2CeyGtC9H
MM2U8Up8HIJ7oPcLhlFbJxyec4JcDDR1M29PiI8K7yUMXb5i8gH2oWzFnfsbTDWjjmEQs9svnTIj
Nfs/hea8Itqov1SisHxm0FLzM4CDXPw+0+Jhl3gjKGobtP3OWNkVisy5/463pjYtLf3qR83bBThv
Iaxtk4RpTxAbyEmgFoMY5cNu3Ek8v13f4aLs39je8Al0XMBN7ktfH2+l5qS4rzqg7TcC+ngC1t8w
K+9ELvh5yRwf3FPQtR2ABoPcYkoY2oTXDHuaGBOAkKA6ECwwOtSp59tyliAOeJ1JRx/4wQMjfUJG
yTWK4VqbaPuhV0MiFF/LrQoS5SBxaYi6VyEhG9jo92q3c04BDPBccPXyJggj92AM281tusmKWwqP
D39VCxK2YXAGB8GbWiCgRc97RtcyCXtpRmobur6hXiwgWy6AhfvvdKNN9hSPZWnRjm4mvApM4/0g
3BIF0bZrMb9EcFnspPB52FXV0RwQwpBLhoyhJSHGlmd4Iup5NHgvxxQgdDZedOV3eDVhhsxYDer8
Ar/DQk1mgRTj1/H0aXnQ764GyRVVYApMgkG5GPGkxkLFvGvS8V/BMIgNsqqokog8jbPFw4tF+npx
3vH8cqTlFsf5r5a4vdFc7dtsHpGBibBCLbUAnnExJu5IsMwITpjX1MTgIP9bHlEaJ1w8j/Uoyaut
slSqAxwEaKEDzdAVo/bUdFDF7EskUgq+p0Inb72ry9Z2PMJ3KY57VNq6PKczv4edY29GRlPYwN4D
dYYvjVK0lTrBBhU1VvrajF83GH02JHL3to2MBt4hdzBb3DRKUOMapk78PrciwaohNUTOWtDw9o48
YRHjfaT+BEeQUcuwiza/PFQ3y4gY+97nNYe77i1h8F00TwN8bTVvoAy3F7dsSa5l3hqKuSw24z93
sShKJt7vgcyJ+Y0QtxJFzwRvwzKwTKSyzRVsBJpKZd5PSRdTxMm/Ew1/p124RAihliky8YmYdm/j
o2vOoXLyd0WcVA8jMAqhYVPOcQFIi3v2Iv0MqsRfFvpcB7P8r50shWJ/Gi1C0+LiwybJJcbgkAYm
KY/j8G9ZIt5Ckcm1e2a7GCn52UJGOlqmsiMDt8JkoSrtOTU/WagtUzBOrl5fMTSe2XROHaJOwZGP
yxI/06W7bWPpvO8XcURjwm2O1wVwQYTkDPIIqAORiUMtjULwbI40o0Me93OszgH7eCGJGo5dnWEU
jLWZp6ABUVa7/J2fG73Ku5JfT8YuFh5k08JoJFD9cInB0P78GipiBLGnYGMjgjx0GBs3Tm9LNQto
V9gVMUF0OiOjhFtuIxWYS8Ku3BTIz1P/zH/iAPql46HalWevNh/xqWdmUSXhtwels+T6mPEQ+Lxe
Pub1ftqw+EinThk9Nms53GKWArgxcRbAwIEpRqseVcFOCAjyQEfRrhFD2NiLXJr7z46D2FHT0IHe
izr3EAJYwzy9DZC+dPPccPnZDvsN8I9uxSj2ykTn64kSFYBrJOFnEP9e0sN1jFrzU1NEfermA3hQ
9z1JFXoVpoL4U/pUYS44ekn+K7/bLsKEUJ4TiFQd74y9ct+kgjL/1Wpt3n5ovocWSrGtAr3foqTS
m3m4QIAvrPJVVKgIWn3gTIs2k5EpZXS2u+N+Fzv+cqyUEXuIukigWkHpVSbyFi969gVVSvch2EPF
14hOiJ+BYS/FFTtsPWHGP4s+5rxoAaxFz/qEBQkeUd33c4+kYnOafkyY8LELE+9djzjItjzkGT9Y
osdjEQxcxdrTGKAdTsMD8P1RjwHS83sAsd/ET5y2woH5LmQ+KOnMb+TmG95hXn1Pjd/OaC9kkBTj
2GV3hegu2LcJ5YOEgqFDtSBwPUPI2B2cmvrq1GuYmAReN4bcXgY+yM1dC0im/nypu+lP0zYTFewu
wdNVx897fXdhJfRKET4AuS8cIq3GwRESwWT3PPa4mFQdoTWkwTNtkydczGzdOJR0SjkhzOu4+bkn
/0PiOdyHj8iuZOP4HhmrLHQH6lTts1pbUHhrcar0cgMvu1gvWGqw1/sqFXoyc8sGH6DMrs8GDyPF
ygiEITtjmSAydvret4fX14zYsTwDPuDd7bvYUIGTOIU23LL7BisymL4xpdOCKVkiGhRRySxLcPp6
dupw6I19mg1VjlfOIU9yYhFmSXi1q5FNhy8mST7TyFFPg4hfHRPNZYSubPTo9Skj3ZfYbgosmNkh
Yf5X/4gWcMgKEiM+93oxboEwTccOS4xMh8Rmm6bu9JVMjR5ijd598VYM12EJQWzne+zJodoey6bF
hyJ7BJkJUMEKko+BHcZPwI+ofobwbTdvmPk6RMTdO/e/ps71lBfb/jN0bWGp5xdC3gtqJM5XenrQ
a16oDVp0rb3ysGUIcqAglDl4SIq7xKvQV9aPA8N6yPtxHSksxCQta8RmcamEW3kkV2159Dsu/yLb
uJcatrK1Tx/zXGG/ZZgtBQSKff1oLnyJ/p7L26oYPEHBNbPEl90TMq2wtza7zS+KmLUQTH8wos8c
ZZFrmymGHt2fJoQf1HSAjZ9QuUuq1azKTTygYP2OHMu5ZxO0tthWq1EYV0B9xRBkVkcK0BWopmKJ
3OEy9E3xRGPhFoibKEfZmKvN3/W+7a++wpAbkSuMj265iUQGlyu3EQnvuIthBpfUjoJcd+1DXVXE
SoYTfIrj4lIO5I0LtWiYT+ESnP1lhyncVRHKXOERyD6pqfCO91zc1tTJsKrtC/M53hD0KrjBrObp
4yUhhGN8iBWxo++bcfTwK3KCHTS2PjdbBuoMJrTezqD7k/fFQHXM12CpluddLKeInzQnZg15ot0b
U2tsQyxyDYpFzqAnjQOTePwPW/rMwrxLHds4tBwG9qU5wgTDTetx6P3JPYvQ+K9QAmaXOrwWbJPY
utr7rrJ1FDtg6vo2AQkOp3wpw7M4f2Trjj4v2wSHXgCUMEBDFueHE1cMC/EUjNL+m0mbeNVT2+A+
Za488IaCm9IEVpsrsn1GXCGXy18kkE7nT1OKLnw5r6FSTw3asBVR3kjEPFpq9rpCCI832IDjxrsc
7c9EmO+zZIchjh2WQpQtsOtw9oESw1oFgizAroWTTdXRmhGA++PWZ3syAgmGSAbifrxQBKkV9w7U
ME+93HCM5+hW1HbAykmBKVDllIgNN3I8lIRELSSU4WTCsIBVGfROxm4rK062jE3tFsZY627Za2Bm
ehJzZjOb3t637e1m4zKMWDK7tDI8xJ4xwPewP06YJu52xNLSoYisaN0tPTCmhAa0iN0hbO/KIUoF
T8YZFh3NqNqgD7ftIrOKo42YWW7pP70u0PgtGeve/pYhSilLnxdLqFd2gTDWOzvj4P4fldi/PGcn
Ok+comv2xBgePawqXFEHSd3FIAapblLZ7DbfxRfaSE1TDAj1/vYwYgh9TqHrwCcwAohMzZRKlccJ
UCD4VrWPlt4B+pwGaLHxyCANxOPspQ3bosZAE0LThGKUMlB4WK8xFBsOBi7Y78OApSIF1NwkI9lF
c5rAIaPhdD692HjEkDXk1ccBO+3Y7trX4XYP48Z81T/CCNmmeaPfP40XTDpWO7YwK7vml2M7pxxj
Q+EzMr5Nr1aJg9eroXYwlSmLqla5Qag2P1EZyynsua2e1FYZ3iwKXlgePpR1azrnwCEdrUusP6/2
ZIOuRX79lEZE6mFjIO6rjMIzqQ+Jj8xPef/p26kRXgFE54LxQjl5f477f040saTw3WJ2kVbBmFLd
QAYjkocOiW+I2L2ZyrfYsxDCtx7Kkt/WTdZZ+fOEPc2sTsdfq1AUxk+3uAH/Ae6n52vPiu9rHqRx
GfPuX7ISK7LJ/VFrKQFZpwsZxxZHIo33pGyUBlNyJhyz9JU41NKTazAgvkMAvvm0aSRBeEjHvJ0Y
5sf8SeDsVAK8Okb/01CrHU6SWW1mASSyg1l+uEWFxIMqdpNGSXkXm9AZcAXRuR7mOTRU3R8FfUFM
z5y2ghS7xBr/VtLWXf16px+K6bsRtnnlThC7E04ERGXnOdeNatT9cDoQFyMtH3fYtHcYhtLXH34D
ECpmp6XRUa32CaI6vPIUe1WHq5HhUIcVMoPGPDm2iwe1HXEEPTC3bw0HFVY3389LeEyh2cYXAiJo
CMIGJaS65BaMzxqMPR1beqiM4PyQSOAtGHZXTvk6r6hAHfQlM7nFTgl1aR0e1WfKc4g9T3k6MT1u
Z3EOClgQB5VZbehMrAr/MoW8cSXWuAisV0pdbcAnJkMHOcsVEcp1H/FCYXwpvR8eb3g4WVKqVClO
4d1NmVonIvT6695gEG/Ng8WJ8h2kFKDpRoplEIKg784ebZdVNjwSY3bDe36DOoaVwtoZ1zaZrG4a
6dA/N03OVBWAt4EgVa369xLB2R9lXbf9IncRxbFBXk4Hfj6SJqN36E2MTccdtUO3wEuc2axoTgsX
Cl/JLKgb6xXZ1gjyLNTe4tnyvV3opdhN0nuOkikoG1UNzHCofTvx5qn9rmWe1JmDhHEc3paDH5/b
MuTV7my2o61I7z3AP3K/3q7UZDlSCNgrRvJMIxm8bOeBzHvtLEQ/lTOFl8FDPa4ix5x1lMHVZPMF
A0xPxUbNOQjEzTpTLdBx/4MHQnPvE9kw/Mb8fxb4bnaWbKlRU2iFByD+5zrXZ9vD9nAxbh5r3GLM
rotCggl0wF/iw2SNqVs8rUtvaQAyBunM/gU/ypBI4IjkwAVhBj3X+2HjmD6v+dJXyaYuTT5GZwhI
reBOf2RdP/CZLV2ftJ+/gVd9vdQvilAVqVDIPQhtJ1z1Bq9jY65+5nLA6Bf6QbXdtXly5qjWL+PF
Eu2RQzbuTHwqmQz6d3da6uL4OIBPMcJuZT9S29aFLmZdStpW2jH0n7rNabIaEYqaIlTAhoTlvgFX
g4zUlAYfVzzdCUfVMt11AaubrzL9GPUE9huOpvcKKOOVnsc4VNqSf7dL5fVuUSa+riVXHbps4mIr
AJfniYQNLL/vHldMCQj3a0OFIkKM01XhWoRgJWKzUsw0fpm4m9Jj2yQzdhKOYGtQpIv8T2C3nJUV
15aZd2nmaFL9IKSNP993MPb88rLwK3e1/5VpAo0AYCZooBxOQVDm1NEFRUYvLTxng0ShKlWzBTwh
8uHWA6l8pjYD+dFRmhahYg0R1ELpPqPxSQtudSn05L72VeMOqbbwO0MUwuLtkulYKVuT5aWXilQg
b7Xxzjuy9YSB2tMdPdlZz7SYk7Gl2E9dobuNZa1KFZUmnLQTFPs9D7GVXTPpWMQ48YjQQ/DHRQg3
P5TXZ19YbI9TabecjuWmWgyDuqwCdj0ghSXxTh/PaKvp323mRC1Wxew3eBQ9MA5TA8q0yPWchujU
ZopgRXWAUTn6tZ9k/ojuepAV2kkGGKgyJhS7FvvPRN+Xn/nhPTiUzBE6iWc0xPQbl45Qe7H7fnbO
sMMDT1YgRsk4jKvpCYI3N8BDp9I7qHdO1RGsIrhIm1f2eff+TNPAlwk3bR7qDvJhUBGn0pDIIDEP
MZ72ItK41qxiY1oPBO2P8i8ZcovldJOvsCAEMt+2qkjU2qcVyC02DdqW+cFEA9FJqzaAXb4eP3pG
px1+7E7VZj4oCfSgeNivYtVLQHFxzHj6iCjuI52njm8duGqOq1U3Pi8Y6Wbt3nbH73Ue3BXKAOxn
I37Qr8K1tCLx485BbRgP7tsxeNIGG/jxelXUYIFS01qmxxRpuwhVCkcC8iRzfux6JTZ9sIDs9dUH
8A4h32BUB5QyZ2UQ8HEeEgkN98fu8G80Fq9HOzLKZe5n9p4+R1XOBR5pbDsYsICo7pN+nUPHDvpO
N866eT8Sv1mH84jtxvY8k8L/SJ98ymNKb4mRsVQ4BTDJ03bq7XX3KiHv1dw8ow/gdvhPlHipWjyf
2Aek2GZ24CUs/0TTM12h+m73uyHve2VcF3RQDajrBVt8+V6IbkDzem/1KUfCWfnWpxQ/B3mL5BdS
7ITcxrmrZzPGwXinScYNiBeKjmxw4WTmOcfnPJqf4XKH+4W7tLUOpdTvPiGUovxC8f48RzO7LWl+
2C9inUtjnsvyM5C/+0NltTPhWeBhsR/JtKTAUJAVfeETMs6Xjy0fQs9LFqnF2roQMU+tzqxtSVP7
zI7JRSC4rGoBK7fAVwyAWjEx2ACPMNlSgT5jE6/7kogShx1QrqoylGJUbE31gwiyPXmy253MsbwT
Ssm4uA9CG8GjXP8wYWXmQkc6vY9SxdKdDAMIIuB3M/LUxEe0DmtnMHrtGheayQdxAPqqBrzrVLCh
BtCTlgxICQtCVxQZldHBWyjWZXBZvarGxeCcdCBHYM+8QqSZjeQ6eL490OKsKkejsicwKdbvJHrk
jAarHwxFs3ny2s2adkqTRiWYc7y3tynR8gi2Q84w5jlY47sdFiomxs61NX6nJA+J0FZjEStnt0WW
KffvlWo9tyufegAKPPJ48NVwVkM98qIa6cTGyAq2r5vmsSWXuPnNxDB3Ptd701SB2eIjJJVkcrvK
O0YonYKiN/OtRcoSwXouG1ZpaylJoUd8eFXuXvuwgBfc4h00lVWp1fmfDyzC476zPjlaT3wF/Noc
9fsNs9YGxxehdMA2Y8jSwB9CshW1JVMyW61P5edPQSyVAua6Rr96YP88piUN5bJurOevKh9E+bVN
hdcdWAI2FVUQtXqutsBJMZBo+v4/rS73xbCT2mkThgR4GNX0p6jFGbXNNg8YsIqcT2zldwvtElze
wqGl1RHN+vPa/a3l/MrvitBpQr5NnLdfV+bWjsUh/8pK/A/pIczg3zNXZgmSwCNKi8x9VhjFGthY
hAq89euBgzkbOFagKpq9sl/MRQ/aj5gpGEkru+svigGV8jWSQmRPaqmqc+SF8Cm+qskf7EsVTNSQ
dNyVnq15AgGXQLy9HM3a/EviTIuoNdYBhOn4bxcll2S2GUPEhcMSV4YRygcxOBmDrCwVqg21wlT6
lG1fzC0jbb9HEc271O+aaH6CL7YL900GVE/thPhdnsfW/09JYlqfLOtNjxqBSumpUCZr2z7UYqXj
hxnF7wtnoSpXqiIaR1WT1EkTuzrZYzASKbTX6sOoR13+OWiuaysBStMThCWpukFqXztPLenm91ag
6liLcnaOZ0NLPX8f9LsJOaYVm0kF05NRsThmGl1K9qwsAHj3jpeOFKgu1n9rfN4jkwOVZpHByIjf
UXUxqHpfgX2fPwWlb8P+j50/I7YKEDdflPQ5WN7Xh9O/VyUX1Il/wV6dyoHJPRL6jeFElK9FC8QD
KTA4kkku+cMC5E9z7QHp16/ceYLYgOHkoVuus3MZg81arUYL+peJX3dp2Vi8pc5s+oOJcNstA1ED
tYDuFe+ZsIKr8UVGmKczQ9qg9AObKhgrX2DsaGi1RVSJ1IH7wUZr6JIvJh/ad+2BgK5MqMtdaCHo
lFFVnVolrozxZDYBFT119oyje9g/31O2fQzzsC801svkzqrmmJJmgqUHWfnvV7XhdoUusKwXQeHX
weIUyHl3S3Lnjc8pSQLTjjuL5fTKK6JiA9cvgJuknIIld8TIaTP+FUMNmXKirdq69pHPbC8U/sBZ
UAA+qJi1GxZq5S5oQ+2iYud51mylZKiNSYJ2MU9OPFRD5uQj2A5Hu0zapdD0Y8lMJL0FWk9KR/9g
+H7f2Me1uN1EGSFJe+cM5gYRa3ngMLsdgd8+ih5Og4TH6EwJT9e8TlVOSojjPJRrs5+Lr1tNBDP5
ahwiCNiAFr53RvJZR1tBTXPPMsU8VGe78Nv7n1hgKU3gyipKqAoS6xJpklZuTB+86lCeAqw+dgju
Xo/6tcXuyejRL5K1/8kgXCOmn2vjSYeZ1VsUDD3iscjA46KELXEFrxu4sMtEEreggmbtvr86zkoJ
x0mUJDwmED6Ay6537xRtlzFQ/z17FdBIYYuFKAwQqG4mipe43rGN4NppMhDlPpIq1ND4viFwLNvy
OgQRaHcsmW+fcFqDRce14wgOi6cHm3Zfv2zfEzveSTVqnUSawud+6BiD3puhYfLcu9JukLkp9Ifp
P2BIDwHkKKhZ267/ATRrvZclvySWLSwhwM4oHUXBW6eHt18aJzuiRHXjW9HM+flLwfcuZCWH0XKH
VHWmN/F1QTmolSscYcCQWhQ8oqYOqN1BPh75A4t3e4pbW8l40WQ29LVtzo20iPhRbVI9SOHCC6qY
AIGEPB4kS+/WdJYfEUYZC1b9r1BxNOpSxyf3IHPuRw7oNOT+ZoJMdukQISpRwMkyk0KniH2dyAr/
GRnbVZvEa6GnYQ9MCtRuEZVpRBxGrQ8SMo/h9Fqymm7VM2SXxI/U4gkup87R03ZTbrGdvLNU7E5C
KImFv69749j2nnIPuzzzvtMVMvM4ZSER+Lz7h6diJR0ugAD/g+qrNKvcYHmTTqBmp4bqWjmQKqCL
OZa913L89kwRxdsC1svauczmxkbc20LoUeNGiLHGMsunvBdFJSJsA14Y5dGgWDCmgXDKd3WpZgX1
apKSQfJLsBRwyTp/fMUIRouIkMxl5OHSJfHvhV+/HbuZeKn5M5AbHU2OATYskAKVGaKCMQwWVUXD
TL4l6gsTxPU4FuKvSK8egiFiVn0MOfBFuprjIlux4gULnmMuRI+aRWi7qwiiwZ0f4GngTkfzaO25
9FUJTd0AsU1tRvaxGKKcsJXTHRV18oCeHxO+X/A01D6lfI/Ts8rn+cLYK1N/xFd1Ej+Zv4EgWCIl
N7qJXHDYrJenrgT0iB7Ygk4aTxLS+tXqb5M1/rzYohHWKk5JK1aQYVJfqWtA8SFYbWWYUT/cKf8O
TQfx87SOyROFOmPzoDsFxsoUFyVJpkVBRqgST4ck3Sy68sz5/+TXYYWReUmTeKHSscwGhd23wAp3
3bNxiimbbVTY7gzp/3LVrY470KHmh/T01GEOqPMpTe9x7teg0Maf2dtOLHbRH/YxTTpGpaFHPvcv
U6JtoJN3Ax1p+8Q3gX8fJXzR19y5oAN6H08GNGlYPJGCRpNgscGPRa5zXLoQ3SM5sB4UW02qmkjB
gGrA4wB3toez+2MrTtwanO5vpO62IeErcXptnJ5DEMSaL/yjUHZlKVxnKfUQbTKG4XIsJTgl3MB/
+9kj7Da9zQaLpm7vvkH+IcDaf91YpqBAO47KS1YQGRtj0Ja0EpxEL3u5i2xRseiicRpb/BX+nUmd
Y9AORNpCvFtNtdba6H0fQpgyItF0FPvns7bHjg9dmKW1Nm/+2h9p3t3TZeahZ1jYYfJDWYiqPrAp
cDX63dl98niJd1r+OTJgfbjCfWNn61y8oQn9TlDt1VSXXr77yeJg4v78lCFLWPowTbcu0sdrzfgV
0ZvkYL1E5RAYESs7ertnRrTpyHPaZMrYOqgzecgTkij9AQad31G6IQb+otvTN/mLnOzxrg/4ppZf
kqiU1WHD5IKYwS52+nCX5pbCb4wolpa+0iXX6GOgxpQ6Rd1gYkJwbwz7Wkoj6uXvH7K2FlEPgeZr
5trzDtvDPdjvhnUZ3XVTm9f1qyiK2J7fEtNpeiDtIgIaW1K4v6vDNQYTQwAetIt7QH6btZMEBMGY
KQ6nOKZBSagnnQMJw+E1wJ0fEz7QXh376ZF30kfe+8rmTlLTtSAATmzkJV3YSZ7FLu0mvVgeENA+
pkpzxIxhFnFZXIrHO00wQhU0O5aoYa16WCsgs0xndo1hrJxMNgslKAKLQ73CuoOM8V7BhcK2t2p3
4mSROXYu2m3M27TLC426cLxjkNPvRb79Kg5HCVIAQNKeQhKmiBMVWIaZMzZPdeV4t1JXzqgDxzxl
AY9HhzuCiu33je15M6UHI2hAKasQzhNJ53xWTyecJcP/ZebYJDMG7RZNwBsZeIgFXuq1Suz4ffLd
n5SdRCex3aYhu5LDI7nxodLZPaxAl6xZVpCCSCjxMl0V/wv3Uh82GBI6yeSNOhssdV2SPcL32Y6O
PeWrDoVk1jnhhLHqxJGa4u78F5XE8p3R2TfyaBGpqLt31W5ta20HQN3fkoP04wBNUUZHMvSoRWAX
Fw93soazq2phRZRbvqB7qg4XoAkzfu+n1yhqXAb3Yys+EUFmwJOeEKYa2t8tXwrmHjL2A0Qw5hnL
Jn/5bON3m8kXjgn6lBxCCyqTSRX6q+3lKZT38VgNtD0Og/lcY+Cg731pthdMiPSntv7oxtgmR7ai
yWJHy7cIjkBtpLupI0D17hgbI5YdZfH6YAYzT6Q/M3n/nZbuwxlEFpUbS6Yk15Vn4XnE3K99mfbx
9ls0mx/kaIWLIu4LcwJcw1pn+3q19HrTbVIFPlohh0vfJZ6aHeMnC1QAjPE+ux88B8V4UtMdkV4G
wXiBkMMTAqbinwd9WLv9lYQNysp5LonfqEIf+IY71v55i4rxF7mx+PPwjIbYZ532jYdbjxzFSHns
OkPYnzfYh7LpJmx8EirvgBx545XTsBMe7oAHTJzGa8w4MMHP7TQrmg1NFjmH8+GU05i9+XfYVtOb
tzhENIOPZo5GHOVXN8Z/zGg1k/BGhgdNTCKcVTr4GvQQuAlmtPx3J8HF8Ti3JYrw811AadkQl3AI
v+rEPpRJj/fIerfYb5uKTEb8SiATK820xNU9M+2xJ4AWzZX1y3J6QXnimR9xU+VJbkIwfcZAlp1X
r1IFa3KaM/Exa4TTI7Tn8JT6urbpbFgfvAagIWy8Xh4M2gmoeJBv2ozZ2TCw+lqTrWXikg/JBU+U
iTbltjzAegT1UMcn8bkU4LMdXbyQGRBrn8Jd3uuw7DUIRdm7QhUz0tdrD0zXK7P3WCLcgFBlipZI
/Yj/XJZFvW0gjx44qwvqbKpar7tiOtLfR8n+cEtvptq7ivmP0Dbm3STCA6nlgj1getnXFwGHKJ6a
sktz+mY6AbuhbDpD7gx9Xh3NuqcvOB3lCLtecS0AACBZW1xSTgr0PywjFj/DplHTpgNFGeACpxhJ
/7kKJfxJgQgI71Ou+cblKV373iSZ6z6ddlhHa7YI5laBGtMRV5huiwKpWBOko39p3LnT0DUQHCB2
mjP6fS+XQEHfazAvF0Ke+FaTXHBYjS12OiZjCK3GLWTnMd9i26TZLHWIDRhmkLXykptdMNvDzHdh
MeEy6DuS7mOqf9B1YmmpfD+RfqMA7YuQD1G7lhpKtpGIbghaIteB0aBTviOjp9fcj9SkAImf3ar1
Z0PQ4g/kRpvMlpdvD/OE98B5qkKrctIQ0kbd2HJrQlno/GP0HFKHxhnZc5OtEBqLikoFsWxJipoh
UsOHH9gNjnw/SRR66RaPn5cidwEirJP76Can5TQ6ns7dHq9rKTtIxLMPXfW3Hxu5fP7ywMZEjkEf
b31Aqtvc38ubik8vs28YSwefvbvKFBDkU8DRFrE/33Dxia3A1ZnOnFJMF7nYMCPHhReIObpnYac5
Ny6enOpK+9z9jnkbf0YsbEWlqsn9nDUYY4JX4AnvnFFPthYKPSa8l1LGzGEs8lulKEoIzSet5kQ0
VnPDj6Ux+NO0SDkZ/wDzwCu4VmiBQRseK9580HPJHoTD83XiHM5jFf522xaJsDEKPhVRH8Nx+K1P
/SHioWAEFmDyvo8eTvfn0BojubO2Cyfoy4QrucH9S9/4+AXWkiHiGbOOMaiV+GkHchCqzVuoa+Pf
ECCgwaxsiJapI2QVzNylbZBzDq+e8VJB4gyu22mPZsEOy552Cjy+xhL1ijp/9DAHEHqPEl6EXsOF
YHJ/cly+XNx63qIbA4KVVwEJS36ePrGlSgOG/LGXNzcgbKfTvgGJLjwXYwCjd1dqm+tBytC9kx+1
keutGq6mm+h57ltv/buNIm+fiF1AG2ht36pBNmOrgEI452ZjAJiXhTYUU8/4vf/r3k2M9J7GNRrb
KGmyW4OwiXQWLU9vf/ERQL5sMawSoY+m5HIRxth8NwLq5uRP4x5tqEHl+AL+GSqU4isqDR02F1ok
63ZeSAq2lV9JPduqH3MI2sOREoiiXg5uN4rkoZMy2S8rPtrD+YUICVqto3HJMSXcVtIkSEJ7CIO3
zQfU9x13QUw2EeQhtNMiKjve7DJf2vgM50/s1+igUBRaaIKjwO5SkrJEtrtoRi993bobfRbum8aN
3P6mKbW76K2JiNER7/3Zo6OWqMBhSRhDVRkxUjDsybTTiUoXmpolGbzbXlKBxzzc1pokvKX3hKHA
8xAAwlozSyIVxLB0unX3wy8nrqYmHJbrGm+CKfMmEQ2q4ZuZ+j+9VgxV9ETpuetmxi9MkGYB/INf
smC1wOnuunZqSoFjG7tEur3v7eomxJbSRzQ1/6d3nqiGjgaf7/Q0ZyO+l1etUNuZwPxyO5xpKLme
CofTd5BuUIhP58hKWp/0MGTTEdnWh8YES61ZL4mokarrJX7AaKyFadBhIT3cxQqgPIwVRYC5WVty
FxJt2Qr7tvxXRnE9y2o4+FTSWMmUT883bCcoYoXcCVpoONUrIW2hcFVDQ/3bp32Vwr50BGXSLyKN
BpHEsIRYePdNQtc0vhaWHbKc1egIZ1x2G5SCZtL6/C71HPrrFO0nAajoBcaB5beRC0ydAbBcBCnW
owm92/uRx8+cZnI6uPSvcSJrxCfAWtEJ8K6vp0n+ztVWj1T0MG1yqzo8QdCkMAg9tRAdfUDGmH+e
z5Qq0jgXFzCQjOL672fjsGOPjkXucKmyabGZy42zhc6A+9JrTXznbCknuM57emYPH9GWgNQRLWla
sPNaGQgZiNuoyF6+925+aLhr0am/xqeI4SGIPLYgmh8dpCzqM/7tbNAJ9sAo7c2Zf0hJWgtuD6D3
0J6poc1/Z6LwLsW14TBfHlJmTJ0tlYBdZ/YkX1g4N7iGZ0N0mkkyEJ+U/iqtXmesKy+z1ojJcSBb
jjn76+0okDEjc7yxvpEOzVADQc0kTRUEBkIPlz0JDIBYptjvKGB08bjpBGuholErODe2fLUzf4qn
HA1RVFlm+5TIPvrm1oACct5PkAONnbzmncx3HwiRg2fOaxxyegv7EUZqDciGWqQZOVPrZvsY7pAq
h6i8cG9Rafw4imA+SBScLhwKGcM85gyy159U3Z0/1+L3yR9PckVDag1Gw1BiqRpE9hzRs8aLG/V4
wQgczInp+B2KpSiBIaJ/54x8+v1Ycr5BWuDF9eHCQO+R97zpAwWWIGTDgpQiry7pmI1TE8apS2TP
+lEeG0pmtGYWhM3TZ3Za/sXx8476gK/Y1cHz+fyXvkcgRj2elr+/vHwumDpSoHsFOK3JktzdqGKc
dZfD7WisibLEDGquTf+I4fZwwer9TllxZHEnTsexYShqaIGnuHDAjou3XtP2l/n0LnppwBo5hKIh
hANuwGK1OZszTLF1+2xt5V/wZhsRw6yBIcEypXoB2Dp9fXzk/rIVdUJz+HVfC/h4jaNpWjAsFpV/
SWpsKqptoPtYnGxLgCX8TYGc2hnpM0hCDNF4Fx2g86riEmnyHB2APCrzhe4notaajT+RcaLmO4CB
xgg5iRfQikcLKD7FxbeWAUgTrcn/k5pvkfX25wcfrtRsicsZ8lqdgeEyp/kQFeaFaKDEsTB0rOMS
PwQi/w6sQIh3cNSuQmcsYb5pP6NG7ig+XwxANRc4eTj6yohw7K3ItGvotB190Y9HEXfkbMGbQ2CS
6bNPu98Y8utGGF9owjukY0YXs88Kuqmu1EdCSc3hBjcWuDgWe3syKUqZEKGaIU9eUDH6qSSMB1ds
XiMyQvhcyn20VYkNwMvLikuYXpq+p/+ST6grj5o0IdwwoNhZ0gfAKjSjCv55l3mOYNGfr4qK99Ul
kiXe1rwTvt4YuWxTs6RbQec56/RIfEwKLhrndUROgNrTzca96dzhwtYUHjJz7VND1JRoKPZlpDGX
KIDK8rd4AASESTWIL9zI+IwZihlJabWqZj7Mfw5WioNVOxlwiyJcKIMifk1gcywuEq+af72aJoWX
EPKVpKSiqcc66VC3z7Rzakhueu2+sUElJvS8WWUyQJ2OEnuQiQSK7MHiFiGkM2YNx6z/kd5eAfEf
jI6H6wPCW6qXFVT+vDPJn06oEF4Ibrh+UGd+TnwhokzU+Z6XZllui1EP60Xr9kpYDOr1Lr/PlKxq
R7+OWUaarkGRRi5YdRLS8tPT3xdc1Cxu7z5bDyS6XhE0lIpPd1EphP5kmtR8WDbdda3horYw3AID
gQG1iqxim8Bxzxu9F8yKD2mMYRs7/fR1L3iuYGj/rRDYSl3jkpwOCA1ikxpwdlIV46sC7Omvvmc6
/0Es4EwSluT7s3V1gJXbElidvjkGPieaGO0SgmRRnI7AH5z31RMqRfpvSNJkD7UMjUKvM2fsvlvA
BBrDw5KQsaY4V9l7Zr4+OgmFdqxRBmOoHDrfmVw8U6IoMuvUj1Mw/bheXbSwCx9Yi/hJdp+vEZ6I
8CgafN9851IwwL7XQKdqNQfzL5/TUotJ7oJ6MpaZGvhsay+dCB+Ufc2N+DIKlh2NfG00F3Hw0VJc
JaGPBAxT/wEpdRgYCDGJc31BrQzFuqRoeCcOQ94DIg7QBv6zESGbAIGq+GiwBHEJiEf41Eo/tf7S
ILslWDYNYVbWiRolgXAuuuIpjs6aUetpJznxVYa4vyTG6X2FAvTv7RORJzYutJYcZVNZEsM6zRQG
ZuXvKQWnRct3BHJgsR8glyvVSrzj/n/9x5xOoLNdNfxkGpP4714FploRgwSF2UqCa9KEKUuHphov
k00bf91nPN69fyhWBSOYC2zO5beZutw14uv+7QlHGN85IO/GBEyYMvyNuPivSeoFTOVl4n6Twbbx
0dss9xhsCqaj5BgXm9JWTkaW8k2sg4ELxIpP105+4Kze4Yf4opj0kygAAMoH6g1bQQPGPkjJszPQ
SmIuVC7MfZZAnsdLl2c7OJPs3sYzUfV4kvHDfNA89ffb7utq9a4vr3K+vJljrMYOeH5SeuTt1O6C
jAVrF37zYviUhOdX6CHPd/ZgBMERn0x2nRC5Z8BgCJsdZ0agve2fREaDAkbED8r6PyaEWECKWp4/
0msiqHlslGnaIPd/U2hOIijOnGYxFJGzBhzXJIdjmUPzn/NZeWiy57T+AJ1fvfT2erSGQKOUI86V
WCFgmUXl8NiUml9PesLJopzuhmdLFtDSRi9HVDoBJQIdxey45fd4bpZ9oGxh7Kjr12fdPbYF0ulv
xFXj11poLYqtutiWwU4k4/rii50/02H1SjYz+kFotLqolwR1Za5sylrn5eZUTL0KBnwjcC45taOc
Gb7eEf/ryl+rF9AWkNhURNk/FetR+9U6Dfi1nhLMa1XK25BUOMlsLad74jvKju1TeqnvPcc6mOld
FtZcTWI+J/eZbPCJX2YlkKNIYpgo03HCq66TnB0aPLkqTW1AaKtuBShbgtxpTNurThFW/+q6wvOs
f5LHyydhMbD0l4A9lHqofSZMMIpadaXTc8pWtJzeFXabr8h8Jdk5C9gzQKT6W+EF8i/MBWHf07V3
5FYStWudemI2t18pPRATMSRYHDCGdAG/vJ94U7MGyvNjZhS8pYA3L6nsuTAQiEGiYm4DKyTi5DZu
0kMfd8tNXPWhJQzgCdNC/0RnL9zVXebtd/9dcMTrjX1DZ0yKNovNGfnP7itk3Li9DBAxiSUuExAY
a2X7CdI5tlm5lP2fnTFV9818tB1G2KZvqbsRR2FoU5FHznWr8VF4TmRjllLJXm+2srJtg6KdMHiK
OpEZCVOaM62b0nNco3CUEx4RHpgpMk6QIMukneZEicnH2UtEAT43Hdxb/EFaEuR3Zi1W5danzsCD
FJDewR1zmOfZPWNrEZE1iNjfy1XZ4LY0XU2DgwC2UERgfgPvLxx7ja4G//77MaK0Zb4SG7aPUgXL
Lh68d9HZffioKdB/1TnXU1MR+Nbd+B/pz+TxVASXas8wUWWc/rtPwPy40eutna5v/CcVbetyDBa5
x5mLrzCD39BP724/xw5SchZtWV+H9mX2c0IqPV7juF1g0WoVCbpN3vvhgbdcMPKdLjlMTIMBXzZu
hbw17BwnlYi13ObZFZPoFJ+nn3M4U9s6ISyS4YuvrAkfHbx6kSXbsHnNTCH0h52rSPFyWqKFgQ7t
NlqwIuYkY+ZKYgqH+AwuwD8s4pbs6X7a+S3+FOZiHEI0po+5Vp84KcHh3kbzWu7FUXz4Yci/psXY
h5+lmNJe1FKvYOxn91MNlkAW60lTlmGGoRQ6N/R7MaCIpKt5yRMQJO5Ah5Z1DQPC4LKIxnCj63jo
PgB0GgpBubZkZnO7ea66jrY2LPVs0O0gnyZfWZIBf+5IG39BeaJALVmCq48OH93zR29+z+NJEFcD
O9UEe65dcSYUcBES8ZH9MguL6qI/KYgTF7V814dlkzeDOLkQkwjrXUUevPX+BfssYuCJIKAq7R20
x7P7YmuiagrPdKf/lYBNk0L7wxc5C4LZTZWJSKkMMZPDsrpt/nuXemnjb3xhG6SqPFCtktMhMk3J
eZBSNBpsIM9H1gzMhrvOMOGe/f5xE8McyIZZ4/Hh0YBAsx8kjHU+Q9TO3AFYQMg/xpC8Ux0pOGgc
C2S9aFZ/p3zrlbZ0pmC7dpPaUuwvi/OIAk0M+I4vhwiuEyOt+8x+2A4t5yxG+LtwJGgfSvw8vrIT
GsE3hoYp8unFia5kXLgvpvT6vtoffvtOHEGdx9KvLdI+TbuaIUdopDBJHwHTyjiGj+iC4t+4ndnc
X3xObZuJCqLaKQ0HSLbAVFk3qnFV2hmhvxea5CpT+d1LCChV9vZpjghuHqBeup5znvKn1SUb0/4u
J8m0Nr7/Rbjun3Lz17StUHdfy0iIAKGz29yxKkJUGxVkCC5m6fxJStBt5eH9nGhI6EWIu3IB7aEO
19yP0ofOqlfES4VqfMXQJ97kDfN9FTVyMsiqCsCslIc+vFrWo9SQP8yCdP/wKpnfdPNrxfpzJoW6
1IxbQ1BnygKhxlnq0qu9KGQhLDxgwzmjz7hW/ZX0qHF6e+WdX7eDnwFmMFqLTQapXlIaKOh4CUSd
kcxPqA7sPYkDUt/yj9zt2E0iUwk8iec0pRjyZWvZv3cqaMh7qq9u6GtbOcGuj0mq3eILS+NpPM3t
rJqV5lP+mFOUZsQaNU/gAC1cUm8owAguXCkDtRAx280uptksew/T7wWKvWj6ubEfZYLDN8L8FfJZ
l4RVNkIo8dPFmpQv5OmfoVupcrBun3Hk6xnTosyLX8N49gWxROaPyQuntwrFxmzLi7AbAk6fQd1D
kbJFCMHmqvseATvHcoB/rnRY11KZLYf4e1arnGvCpNyxTU5YSiVkwfwcK4SKVnWI7KAuMsCgncBR
C/y7vNoJq2yoEMUVD9oeQFYRmCP+DcQWiPwToHkGgFwPBf1iv18DBoj3+5jNdlpwh8HiVAhLYgdV
CPqZ227Ps7tv75myzlzwm9+KvabwqguB9JGnZFvt90yyz/rRBIARUB17Kp9NLMXmRBZU3YnGrKkV
YNIYCv3B27zJuigOo1ZeNzTrNeI7TGYLMPGy3n8fUI1zFPI+uYuVEO37ARXImStYte3QzUox0x9V
tBrOkYBiz88txTmQ+TM9MuQzFEbLFSv8ZqYU8SE467IAYoOebAEnpmfvFwkrwYeS8on+IuV0WF3R
A4VbuuDNVxEoY3lS0/DckP3W+KBcUx/SOWFQrtc/j9CFwCdzRGcw0uuUeouv7UmWxJUVOP13gv+/
VRciESpJ6fSAXtsppO9pP5wAmHeADzYyz5y8bihbu7DkcPp1mShebndYr8/3KT9oS8NhhUiFwlPi
5Ulfj5BPv3wZMMpmm3yBfwY1b6KIszUaN6Jc8Jz+g8My0WsVlzdna7dE4ySZ4ClwT1RiVZJHiP2Q
/iG2TRfzaZiH0/TNpSfi/35GJPChENjlG5KeM55ygTYbZhoEGm+PaAcYsTh2anjfx7zHFNxxNdbQ
acc8inuJjTSphM9lhpUQzxuoR4snx5J1uZ/dKtR82i1ucdli6qWvl1TWMphjy2MK7Ri1bVPTFWB5
WoPfzHsqm5C69UCb2XrJ38X3L9RWG13n/b2gDwTtE/DgltIfYPQAJyMxbxsqf8MyzJ8z0VsmBpH5
GaHkVWoYDH+8UjEvCiiOTaBvrk/rzHY/YDEkSf1gQ2YLtcZbWqQoWaum3ItNImdXvng953OMQxK+
doBpk/bJUOvJiquu5k4Zfv+gFRNFoKULF1rOglMeM418PbDfBrBh0dGhjN09kwEBXH7vFrzbIm4C
Lnnbf1ql1pMP4MgqJSQ6oHH2sfqquohVNfgelOAsJAG+OUYLAYNrQzE3l5ej8H/WH2duXqpIuWFA
XdVqV+xaphHaQnPsKVGMgsb98waBfvaPSlaj2kkTOgzwuTYKzvM78A2UWp6KtAWx90f5A6tX+2fF
1mbZYZCC3hSgqWjtzAIXti7TPq2pOkjcdmYAeB0f5ZeLM+oOJNOLskyHCJTUoX01bnKBImYQSrZU
wLsmqL7ECe4980axSUmPoPSXJaQKSCJEArdp14s486YnZX/Li45xIH3vTI3pde0smTQ//mOqAB1y
nfm4QbjK0zhRW0xLrxFj1E2Lzbr7rVW+tyn2vmahP6GhxEL0K8J3YqgaZXWrGW3fMe0ck63spc/W
P3Wavt8pE86mXGedXXhA3O+oQs9ie5bGUzQ3BNdv05Q36K5fkz5iEEefMymkNmB+9+RZ3P2wxT3O
w3DNvE7gfbwGnTZWAO4/ODX8UEsxxCybHcSKhPDAfMXkKcXamnHYi7DNCxMfLbsFBLbjCkI0fLYN
Izh/wos2Grcj52r5CI2SboYQwh7J5p2+nPSVtMglgV7R2WnnGdF6p27l0VvlNr0m3yyBd2NKqoVP
lPV2Frtg9at1x8sy/XxHbBuoPDmVCFb+6qV8Un823f5WCKKKuNY93Qb30bRFFgVKmADTcOU6w5Pn
vA7f4MzYGteeMGBPD3NJKL5hS25CXyZX0B8B1LjUeRdjZCfbVRe5tXwuxUxi3CItCQFejtihQt/A
xh8ktOvGrM/PLk/CvoBwZCHWb+Ji02g/7waaZpV0MNppKzvFtXG7AyqSs9UpHzYEeYK54YxpN6W3
l3gCpmRfzUb+DiSaoB6gGbqscNUe7WoNT0T2w4rJ2ofB5J9DNbqtOI0JxnBqiaOh8lkOHAAL+7a8
qFo1sLdmdcvqGVN7JJH5VsWQRLY/49UDfNyBl7+ILKtDXdfesb4mocKZqPHwWx4ANCholpnt+w5T
RoD4GP7wt8cU6yQs9mtUKU6U2VNPwLO686/5cDa5xDQE/XU2fAlWVeAsBK7LdPWvGu8Y0oY+sdpP
kT+0e1pnNLbVGmlVk830Br5XE/hTHWuipgiJfwaKmF3JSWe3FRShJdk0s7cSX7uOalLyLhVtfLuD
Vn1xChbsOU6+M1KKJ7iQUanfSySj0r3M+eX4Q0ki1ohBtj/M+1K5alGw8vmbVl5EUhJdMSO64WyC
5YzQHkrXnvx4sPf5NNsIDfVfn7ZpAmufd2tUPfFUjeLn9YiknBO0M7CeynvTjDu1QcWShwKFE1IC
a2dzI9WPlUveWKMfLvi1FGWdyr10Nv4ySRee5Gj9WFjGZllt4yxEwqR/+dLWIdY1lxQ4pIrqrbuQ
TomfwvqI3zPfFBvQEt2XIgNbYd5GCSWLx4ge3iT5dQejlO33ElhZQdFbiH3g1JBXQlVmpol0jBiV
1IopKky7aKYxSd2xhiB23ljtLpgSK7bBgLue+CB0IY1GmbWrVWlsEvbIxvGlNrAeoCYbUgtWM2fw
8ETt5OVapZm6K4hvm62m/obkID1gTrdSryCNpZZn42u/qzdFlKxhWvxr/5wKgaJUl9l4H8qTmmq+
NkFtdyUx16bsd1ol7dxTLker19ZnwKqDuUkqGSS7mYHJiieg1s9ZeVT6RRZ95ODTMlyr8cx80MFH
ssJWbUi+thipeZA0Zm0+p2U+39ICD9gfPKiopW1lJYLoniYicg4Wwg/+kMHF+Or8xwAOdScqF2I3
wcC+qCB9Eia0MIUhN5NOgBoquuXpW2Uz3fuXssT4kWlbwHHTCR0yaRdodh/gog2VlJ0fgYZ8whjr
IRe/6sMA88QLzAZ0ACVNNxMpDM70GuNk9xviMdih/93Xdg0H66FCLn+Sc/u6JVG5cH6znU1omHLq
tqhyY2S6PLZVUXzntYpoIKda7WKW96F1fvn+aecFOYL5zk/axn0KAhKexlA5Ac2vflhWra9QSbtd
BSis/QQ4Vm+d89FA9XggbRM4vMCBhFlxuSW3Qjtms9Yf+I2C4lveHjJKlgS+LjlYFksMTFEw0vAK
Di/8sAuzeBc2DQsiKFRWD94zQHWDzFc3yqFTK6PfibHmQIT+BgpZTobMVvOyDu3YOH5w1bnitH/B
ETw18CRBaJBrztNjkHSD6SAEMk8xfKvO7OZOZYRVPBFRt3c5rJeYKrShy3OX/qqmco51RpQFxkTV
iz0FFeCnThyrwz1kbakAqO21SzntwGsC13awvsyPZPplF1pIAnlD5I9tMF0wu61rlOu1cVNzUrhd
1lvSFZ8+13XoZnlyhVP4XXXWlD8wlTe4yDOWSXbLNW7dfR+M4gHwPN6RTcaL8nsGopxayqUEThx5
ZUl7WaJ5RbhNJa5FXA8i6LL9BpF9gjFBVo6Vl9wK2Eqx5Dy7tQymh+7bhqgqJ8nTKB6DUa8IlULT
iokAGJi2Lj6NajbQmlvD32Th1t5SJIHDvHHsoEuWh++ulayvj7j621yvemxvyemV8JNQm4dRzDQb
U5LDvgyncKK1dr5NiMVY/AL69hR5Ltf3lbt3HNSnIbNSI3KBlKBE2vBPkdc/8V7RFfniwx52Xo55
ox5cYrPUZxvlRmENpCS3EBkYdTxBwF1eQFfVXXEjxxl8QRXuBtWuPaRwP3JJ0V7r1G1us2cOt0/y
h4ZuMA+3iKnWbxlVnc5bhmCWrDwXcN45qyD39IJXdpvqECZZsiQYbLM7LySzQgvGVSBUMhdoxWZh
+hA9zmGBsBr56q9MeOEJL7sLKgk3hy0qakEfNJ1QBbb2TkAVT10bvEgS18kjLVtcuzvr87nlfW2V
RKJfOTa7TbZ1w1lzAr+baM1TuDBQt/N17WWPge4uJRWt5hgxCktiZUCI8yz+Y7w9UFORwWT1UIOQ
TKi6ccAjFR7vg9tL0tsZN2ctbRFrhyXBNrLw5YQYmEIjxMBPmfV3JUqIatig6UlMIBFnJZ7KQJ9t
Or/G/Tw92icdXEsZQSFsE1wpASjzuY6XyfgXsxBxyeLtUR55ucRIf1zuCbjbYtEcoGpOhV/9G9Ne
bqhkJ0xn67eUDQUWcRimmecdow6vbW6LRA0lVU5R8xTdriSSTSgy5DVSZX8OgzD6TDlYG47a+heY
ZRdNH1va7LByWjr9g9m87TkYD1CyMus5hEjv1fcyYOZraj4Po7Z2/vzvRWOzKSbMKdRvvYpjyvV/
S6BTM8tnnd8NCoc8r5Vf4TuhQSQDVJvPeGBp31CTdxN4oMnsTrEc44C/uZIxxJ7bfgeNhgU3lgsb
l6Xq2rIthQQRBafmciWaKR4Oj5WOwcQ4O2PCHFFHh9tekgDPVpEqtqejlz+eRTdGNoGjh8o2geWw
A5/uSPNnupepM2JeUlpataSWgO6NlxkJMVAGcHTGowj5/FtQ4hGVBfrc2z6Pr/yiojb6Fl55dOUF
C4I98a7/nxjcX3Y8p6b6aJWkqKYVK+ZbqSdfpNzn/pTnY2DmStVLSdbN+AFwSwdpdxd6/ZqlOhfz
a6pxDJ32QP/IGf0o+ZFsQjXIUJ4Cps56mywgFU842Pjw96KwT6VFDxfuC3nAkjtaPROETMwSewnW
96e1BDlskm/egYvX5Wlkph93KAjZ76nYryCboj7hO2lEpl9WIq5D4rgs/uMFeG/SmTfHDcVCTzkN
CuaUFq5K0YF2SfhWPtPHLTCUSoviNjh+LPCcuVsKWGqtoR0RoSLbSOfLOoIY9pccBMVx9V+Zsw/7
gNzQPs00D0T4h3YpVJxifwvvZPTS5Ni0p9g8Vibx/In81BwMKjUF9JEO3WqMMEVlCPC6a3I240wW
v38ucQtypxMVXC7k+ZGjC+b18grm2ZUs+VPFK4dLnA3RCLwUYCppGu3yePBoIeUEsZuJZepQkSfI
1wwLNApGDHRx1RBSi1TfaSk4qGDQ9NDEWtKYOx5b3scegkE+jZ0zIvV2CjSoHzGmd/Unlbl+nDoh
hDL+QIfaARU2EfQ+Zm1jME3rqS5QnC/IDaiyWtNBLMuvA6bbgotWiA0ccQinl76OlryUGNZQMrCn
ZREeg6/CU9zEipVKXF9qjMrr0iAg/wEucmjpDLprf9LcFinTb+RqrHf/uesWTJxq06n2nIOIZYCA
IGIF5MRc+It/D8Kd0B/Lvw4kqWzwY5WvTi5E89zFShM7+piELKURLfyiGulROXn9Prlp7c3QnL93
kOUb71niwt+MHb9bbGuWl3KuV/V8Q5lqT+rCkaTw1BHDcTGBLprrBxcWuni2DukJNcXUWgSMUtib
BZA86/O0YOLus2lPK2BVflKz96CuT51vo4euydeouSHIVaq+AJZzGg9VTr0ykU41C97WgdozBDgx
EhVv7sCYlKk2r3pJyZCE9hBd+nHZwyCijTPDkWFdmC2XeCLpms95InPiL8fEv4sIAUgTMQPs/E5A
Wir2iAo0kvym5QtBqUYZEG2jJgw1OpkLHD7/IugCuZN/i8ZCOtztqL3KZQynrmuSiltZEPS39rNE
6F/uJHSuOnGLEf/fjo7I8Omz+MKuMJjFM8BkWRddSzahO/lAfM8UdS0wK0MosW8ZluSTWsGTsOwH
ECTimtyJQzAwwY5QSqfVBSRFF7O3gLeUFmFjMUQ5O81iCkHMH+B52cOS6wx1Va2Q9yzLPM9f4OP+
q+8f+y3Xw/YRA3h+tS7BojQe9Ib+7asTTCqKp1goalbGtst8puoQ7IhOeha1wwtPRPLphVVE2CXT
G2wLGFtk+6do2nBmVNlFX1NiD6v6zObDMn3DJt9nv21IpuzJL+joAi5Kst4Q9TDgSHFn7EE+SjWZ
2gVLIdnS3j8PQfqs36kIXaWh1u3OiDAWWKqSMCCPhH10vLqckhiuKviyPliD1or86etfPiUhY1w6
avVLSpjKxlBT3zL8xFqlsAY8ZaAa9N3EeehEL+v4EywxhccamT40GvSwYF0ZgwJoC9IHCAGj7pGm
1w63TIS71ORxE/WrQf8U6vsunqa8lY8jFQIwRMV1rcK+s+mEoywZISyQkv6MYzaO80mfYSEMdS99
7CvN6C1ZgYv9oFaapyyKif1VyY0A/JtGkCYXRcgFomu7WtkgiX+pxqUKuO4NCwePrs8FQwOPi44Y
B0VHX+LzXcW3Fwo8NoeUAvSRoTnc4v1VUjbqvuvELgDdI56FBStYBCJPn7nN7ASxEqzbduW4B+YP
7SsDxTpVlSUOGLXeVERZ4glXV/AjIjgfIZFECmR0BlLqocSDWDQ6NkTDobFm5UGG9aBxnv8f6Ufy
GhT8dvrBb/9DNfFMNsIdhHVOb8f0L2fDAqmyAChUfz5PFkUY42GOv/5/q7cwfpzFaE1866AYMuCm
JWfd3VGzg2cjDEAqQDAZkD77SgqGnBWbFfcAD8eSLUuO2+s41sRvxcHd9qh4PHjXDdWA16BqzaBs
ogO30xTsxgo0+NGmsYtBNV6toz9rTahR82GHoGBdQk+O0ZnyemBeDn/nVIzE5Qt49A6KX9k3pds4
iKgAiXtMordC+/MUp8ocNbfZPEgZ6N2HyI3LEY/UTdkutMd0LnJmS8QPKM0IECqrLU0xX5EsnQ/s
SjVLbypkRQwFCUY08fbBOWPwJUnwFBO/y0/6hmsPLK5u0buEbSiDZT+8t4ZnpsiWNrzvFY1qn0hT
CebVa2/e4GDomi5bEoNbQizFAdxHqdAUNbK4W7mPHWjmv+UlGtFhfh+V7rVMSPk/CBtyQekM0dzh
zpIIpPZ4Cx5f4GAzMp/UahDRh3aHUMgUJkAH1EIfqk0k1g1aTZQN9N/o9lc21B91+WMQuJW79/cF
EREREwcPQ/W8f///YpthR8Iz7+ei8Gy/+AYIQFgl1E9t0caQ2CypHkiQHxZcNUem7QkACR/Vs60v
yIKE7D5mIGsp+en7ODDuqfvizA+ZV5wj8R4gfcHpDUeGvd3PrgUcsIcGS70rdvcmr3Rb+Ha6wFFi
bx9/CeUrwTKbvbpaRio/akC/UbjmLVmnBeMbC/qx7xj4fuU3AQybEnE4e97InpLjTeDeZLhm+j4r
RNOabS+EtifN0qf9c/l9CI+MMb3ac/375+CpMAc6x5is5N6e3ZKTM15V2CdcEIyZC2OCUBcDyvj9
62rDLlhyNJM+NYYIR719Lt2hxnhU0zXPHvEjH90qfnETQwvRLUPWoMp4PqG8BizWbMZGhasE2g7Y
E3DcWZpVlb4WzW2zn1SVunxP9ujnSSCqOySuZp4o1T8Krbiwt3Qk3+cspN1QIQk7PWLrTK39oDIS
oo0WuDyQqZE6bX7UEBmfdX8Q+bnAY3C6fN4c48Xww5gfP5a5p3S9Q9WpKUuimicMPv8jobEmaG37
l+QEsFDqE06Ga1VPJoqRqDBDO/muVMWslOctB258Qs9aRx3qY8rq0alHvkVL2uN1vwNpSy3jUHRq
eJQfll8hvFyPdgiFuObv8w8moUjBVfi/2d1MiqjiAKhMBP5UKgtDLOXYb24lIgWT7AggVUFLawWV
+39WY0MucgIWG2pL2FQpxprjaIeZZ4wHXgANRr5ylXI7MBh8nu5GKaPvzMSoVzWFAAnTdubMu8kK
USifJEas+rLj26UE/thBM8z0P3JEOfc7oeShne4wSQymXe8qxs9bfS/xnNv1RHo2G9MKSTqka6ho
qZiLMtglBwlXxrKOQmB7w53hLZB7c2VnpZaGrZH+DUZt/tLokra0D/bJ1ssHtsB1qRo6A1vFg/Sc
QqSF90oO2lNZdomH9gTNrjOP80bb9wJ3Xfr7Zv7mrB8/vPYEGWJx6x7uxLfSfjvAnXnjiWt6n7hH
VVCBLTRaLmCsqNtqOg97lz8c7NWyDCkA9olC2wxkq9Ue1scKHqx2b1rdZGdkna/nv81MxFK9Zy68
hXpaRp6a8/n/reqbjvSfOX6masPGIuQLmH0zYj/D6zbgOoP7Qy3G5VTKyUGdf7qrKuGv/ruffpLD
m3Scvz/oGwWiVJ2X7T3VyLM51u5PMoF5ZlQzdI4T/Gt+aRg2noWkwnjqiceIF65gqQZvsWhNn3f+
I0B5hAnd75Z4Cm+5V7twIDNNdi/ZnpV44HYvaQcokGaDm/I3jEqISFvcyGjCIAD7zNfUMGDuuwNM
bT95MOCcYIAOOEBFtdlfelGf8y0jBytNt7hoqdTMPUq6C3AexYYi4ACvY5TIv1upkUhclxgj9lM7
B4Naoa+TX9ChaSzpntiplFJwIN5KS/i30hBCVf3E3kKLj3IttHfcvlIjIU6U1nWJBY/mdrHjoarL
9su1HYDFuGLuUm/vmQthxJqP58T5pIrYggMK9doRU6Ob1XyPgCKMJJQD71UAnXIKkt+Or3p6xwLE
P3gnXx+VF4K4R0GniJyGIWE+reQ5Lez5hQ+evfBEj5kZKmB+MeAwkC8hqzwdnpokqGbopW/Y0C/T
JBckQKDzu/g6OMYvd1oKZdddOm4wowBZGtqKq0ngWnJ6HGjYtpg6igPLAJEqm8opaCiRuIOvd+hP
eUwp/t4Qs+so03e02u5PLoqJijjeOdlYeUYrLXsGJGzribkuG0WWa/Dg5eCxw71GYHB8jxHayOG3
M1v31JE63imxkcEcVnsVW2ATIvsvF/YwV1/9jqoZTxR9ylrx13ACgs8WiccqCQ3F7fy1UmlUCxKR
7ZpFXAUIAOg10QUuL2zzYFB1ubgLSR5CxaPqf1hsy1Kv0SvCH0rml0WgT0x2ghZEOd/12a8x33o0
nZMD7/vehzbDJ2aERYFgcE5FGIn4oe6aB17GOuUNVHey/ZmCrhAiGNbBD85zrpXrVAtGOifu47ox
lDPefKKpl2+WP9iWQe0QJ4Xar+yy5mFlNgn0FhnqfLUS6BNltoeHiW6l5AJeMZ/vo2xC8Hh7giGr
2hghw87BJNO/zP/orjdDswigVrwLb4gxDHv1WClvO/GqRbJQueu3r9YITJJItciONdh4Q4kbTa9M
uG55w3auCP0HNidowwhpVLVGGdM8WVbGZOaAYOCciR81ru5wE5ekHXkXzqrhIVUvDZomxN19NOVv
F6CzyxqaEQ6d38EGt8xU0JSgytO8XFU70p5jpaZAQNkPLelV9sKs1riqfR52XVAiQ63/qs0904Fx
UW1j3eNMwruVqjk6lt2WdckcuSq5kt903fcX9okv8+LlVcZFSqfd4NIKhYyPOKew61psiBrIRS46
0qU/4bKoA3E6fzB3qXmQndmqvJn5XuFxa/7n3lw2OXl4VcM24qhH0rxYKUNu3r6bgij7hZpcaVmu
pzUfNTW5O+us15ghX+/umj3OQ3JpMRmShBvX7FTWcD8sA2cu6yk2G2j+PR7j5TjbmSXt5hImvKHN
umGq9PepqIowhUQ1uApVFyNsA5jU0BKqrACfwoVcsr1d1BPzadhwfvIDlgEtwoqPjE6qBj7/WOLh
k7qXI3olpVTPdoJ8wUBxwzYqKS/y5+YnHeGb6RsUZfJRsLQIikKgmRPdOPSAnd/vQMSIaV9suZY1
NNDI6nYPGTZpLty6gHHj2vQy7vuVV6z2NsOK0g1lREgWIiMabDBkimDDrI1r79WCa0dz8oFArT/w
GNSknrItIYHa+9fgK/MWBmlI+ueUw9lbB7VpMCkUNnFqYriE2h1rmEog0LjvfazbbPwbaK3LW1xL
FYrOSqa8wky4IStm2pR2wCwuyDWw3PdwXaxK58prfc9Fx4mueIYqxsp8Pvf5XPw1w+eJfnS9wVLT
TjPar0U8dJM+o/mpLxIHKa4YTpG79vxyEdH2cXESNHPnDgAO+G3zCkJRyP7uRTExnvMwmncMXdpv
MNLsvnDRi5Xbt6buJmIZW9IcJSLllGeD1CyHTgFxHr+yHBKqbAb6Y/5Ewt9aV8VixP8nSsCUQHNo
+l4bNhsK173L/OS8zKA/v4mpOgwNpoX4oh+IOgfYRmGvZheEsmfvwXBCvnBtm5YGeDkqMKMQc90S
QG+n1e9XdiwfQVSGSPDnxRF0z4q0JiB0ac2Rl/0BaoM5iHWyHO9xMGPeZm+JWcFZ3MhJg/zdpeaA
PR7cw5+BadsWSwDmjmdm37qe48XyEq7sFkp93K8ZMEvX0vJkv3PL4iGfENBbuDUZWTCNd1H52NHp
xtPjPPUUhHT5wkhvThs967Yfz4qTIe4/VZL2nlixo7ahI8antHk3nBqITTbFpMh2E6e48yJFKNyq
4BV87VTTeqNPiRn7Ua43OiP117NtWM0ox7SC+Ikl/f4CsE/8cme3RpnlwyBt8xoz4hWSEK4PJ+om
GpDTSPlLkDexA12U14/+5HxT4Jb1+rkPyhQOaivf8eS0ThTuHR6Ck27GqOb8w2PIRSdEl0zyeZJK
RHqL6IHWnL6EMBvCnUmNVfT1GopiHuGQxvg/umQRXtif4G40W8doO0G5NWX9UI2VWvrzf42NMZIL
/gqJRJi/fyyD9uCc3bvRrpQAtephUyx5fH+TS4UUxmkr9TW4yjIzeczbnY27qa65iSUkibHxSyHW
1ZWI20tQYUQJCC6blUs1uBejQjmNn0Gu9JHZecUMGKZA8eVdQgikJgzJAU/gtGbsI20dJ7JM1JzT
YBWUPifhGVv41Fo/K4ZMsgKvUx0dfmjDRsG7tW6h+9SQWdGjPYDI59JtLp+tLLtm7SjQrB745L+K
Pm5NfpzmkL2LECNFp/dG4Xrs1rVj7Mtopt4LMuIjxGGLEgn2b/6eGzcjpz3fcMc1XDyTRD67POKH
6JLL5CSybD2iSCLUn9RSSVUrmCUzV64CuQHLGAVqtdfzp3rUXwhR4Lj2vs0Oh37GHCk4xgkAbzFd
J0pd96keVX0fK8lj3fXUfwaaKoSAFfO570JB5d2LAVAYPzZwnLvJ3/PRUN14EFX66Ik0dMEl5uuN
kwAP6fSTTXhUH3IXzixHSx0ADGxPzE6X7Sx1ucIgQmcw2ovjTvoEJfVlAHGDV4sJ8epI6NnkclV2
kN8Csw3zS3d8xI/Mq1a9ow+dB+fjg9uzml444wNRVp25j/h8wJOR9EwulgWw20sNcaE6Vcn4UTmr
k2N+Pw/eDbbN28jiy0B4aylst+jurEgIbvX9GxGkU+gcjVtqgBtAZ8654MV/KTXigY+jdk81EoXj
iySewlmmXNFN8ZX/A3zWArnABxVt72KCKGckrGtOL7AMlXqgcHtgDKqF3/2BkvbFQhtUDbZVnyuV
zOcbi198WQkyqbGwmrsJayCW5FkVbyzPPtQ8oBju+V0I9lfXW4RUAlrrWL0vauf6Gr++xwRWmZx1
RZ5cO7W+cdeFrSLb+w+1NX+ovDXAMSnVGmlxSlAwI1GTLvcqzfG1Eliq9tYy2KMqVIneqPblSL1R
BqAylH4uRIdoZMV2X/rjxPr+cpAliScYPkHhG/F+QnQY96k0cd0ZvFVakraDdLHrUVeT1j9eCclD
8+TwZWtn8ntA0yKvEvW//dmRhQr+dQCZjLHRv498NiFZBNfJV2LrLu9+3o6E0cCshvaONOnGY/md
W8vKOlUuS0qN4eCN7yquKnyQGufbA55IjAk8azRXrt7KoWTUj8mLEJg189iUz6tm2GN0va1lXjTU
P9GWmWlxVPC8+AFjT1ILPtnoLpVFMn7S73W/3o8TPBukrailiryadRX+FlPtX7Svjg2ug+fNQocs
r0RZ1jaBap7po6no0vA9Ub4+SWyaZ9Bm5+bu0snhl3NwCPPz10ogdflbke5a42xAC5h7cceW1UsS
tD/DfAN6lORGDMQzhkCssKsLCfAJ9kXP9NoMkLHI+Yrd4Z/5VByDP08wWA0d+9RqNMMP6/hGjZp7
+ilpjEbVIf75uaBPIvmH8knJVRbbblrDQsHFE83gcLJKBMqsJj4OkKk8wy3QhTlcPE5fyIqjIFTj
jyViXQUbMDRb0sNC94BfEQm3vOeN0fypBx16v0KFgdlVSG9Nil4By6x0DcRN/zFQyP269A7rJC3i
VWqDr6492o72JMZyr4FRBry/FZoxF1/wbAz3nxYbaAMFZAkI0lwmkLlnicUlt1rm0FCs9RuR6Gyg
TwN4WanwWNo0m2FGhvb+Hk6zsXcNbeK75z00BNZ9rP8sltQkSYPzV3iXgsvYKWcbh7LDXm6QJRwp
npji3g4TCr7BfqkhSYdTuAli7qvNPuJJCtZDBZev6I6HkOu6QUM2X2jxVr+TEYNWw2/d4OMcCZfv
FXlGZvy5wCDLMAbAHRv7iHorHDR5pYoLs8+Zq7qlu7Dr/JSigSSNh53jUcKty2xp/pNAB6g2e+5I
ia1cpOPIU1n4hlI/FLEUAe9VMYDf8KWN9U/WhoXwZOa4b0b0wTMECuI0vdw6QLfZ6perF3UByT0W
+8QrDTDyYDes6gofr5LTDz2kP9AauBvJclcD+S9YgXqkHxLNN5nx/26SCx5nbGPazj2y9v9E++Kg
DPXuE3SI5Vc7wfhy4pSWMIzr04nRhnramZZF+mVUTg/LlrzujlQ14nS85tgIl0NY9tR/R9GmnaBl
lMfwCh1g++X5WfPm+mZWEgyK+Zyfxjea4dZ+UPqhAfNZ90SjthDo7cY+3rDs549qG2D7pbCHssMo
Z853L3JihZOr9C8CUxc876shnR+NAq2v/yaFAVZXsh6A0ns8FFSnKWTGO5yxGbs07evLZjupRpMy
/smEey+aviyiw9ucfOh5XGyVJwM+1je20l8ggE9L6NPTKzHe0y1RaYG99cMo667M0KcrD1l2pzMz
Gl0j5Go2ZHJBHzQgOk2OsPIl3HNGPi8h36JFCXUZrWhQX8CdkvfxHSK83OrgXeuw+XYdfd2Mr3EF
vrq6rmqwmEXzFxNBPGmu18Z+7kOIogaTmV1QC8geUJACpMWU9Htxz4O/+j1SiYPBibMraR+5lOJI
q/NKhbE85qL+AfvnBwv6/5aUINyOIxPVRnGyD9t+ZrmUWoDtUIy0cLwt7Ku7abfGd++ljkxwmqqA
vnkUGO2b93LvwOz7MBLH1EkkSH3mWwbpOQAt3SZX3aIF7HoeuhMQof1y16ALfp4gcZ53d1vwxOl3
sbr46NwTRF6rI3VASJpPy+h/GGYbr7mQ3OMu7qQZIXtD4e4JXcsv+lO7iuPFcdS4ptkkMb7GwO6d
aSPvmsSZqvHPBZIPKOpPc58DH4nUIADPjjhp5YjAzuwsYBSBt9D4QuB8m1db5fQU9DqGOX0BXROE
qSJZBkO0dAsM/zhLDhgjpRRdspTxsy34osgWIrz2rJ9PkVGOwmFctcFPe5QWKj9wYkMm+smDIBnw
I5BiTSEqrdEXxaRPHqwOfh1zYFi7JdySLbFb7GGkS7lnMKjwTI258hPTidcrP/ojgjL2ejjgkpvf
P2XdtM6cyFj2JxDwW0+gbcotJo7NQTgSTLCmI6JAa2dOInk3nZK0kzeYzklzTOW62JaaHaAeKNs6
HWF3AunMaPcKrP6sG4ndoFyW9RqWcdn5YiwEmd9qe8uo548s5EKIDbJkkvBhQIlT3JCuhIU4iLvk
8y4l23VjKmm9N+CvaGJBqfkl8G80D7QZMqkIlGkNALEK/BZe7+GyoEl6/+3HtT55DKdLQPbbCM9Q
XzbJjk50YVxKcJmW5oshyP7NNeJStIOEHJKRwNLFEZmxgTiTW0d83+2Z9qYL0zZqSZVOsa47/VFB
p1d+cMf07NTUf7Eo7FIKXJ9FIeabBwEV6YgPjPrSBBCXyNBhO+a1HDne187wYXP6tS4RHGGMKuQ+
0qo0wiapUGO0huibALcfujkoX5MsCXy8lKonho8IzseXwMQOmhD45LlEZxX18B1hz7gsXPUzKCot
X9fo/Z76b/TS8Xi1wrKDdZh8V5H5OJoMwsu9j7CShsHbeCrbgUfMHM0U1miyKEBHMuvKpRr0ORlR
iHgyELevvhlMErUjxxvabzzhLY/ayyqj3TGbcesFW2Uoz68wAHaSxGJ250j37x8IFiQFgKimNeln
1wVHtcnM5BRZpO2wG6OzAJAfVG4z9qB3MGDq8rcTeJ/m1UM12/5juiDHSWgaCDElp86e2y0NQQvp
UMKBKbKJxgPZicSIBthx5mWIZG/HppavRGC/h9dVIffTkVTYkPqnVqwyhw9nquljf9Ua6WyIvqUH
22m1mDY5HD9StMNxFXM/d/QWwpHobrdllhRjr24dm/LGPsv8VbQjblNWbqGJOdQCVRKSu9uZHy88
g6HD6uALkAyDM2S7pVN1+37IjbTOP3puXuM2REvHc9s/sKKIQItD0aYvuH1tHD13PXLrlhPzjsyr
MyYZbhmUZ4VGp0LSGDh4Uy1YUOpQmntPEWsXuWvjgnrqFwqiEQh1i/8nbTrCM/Cwyyw2tKngJhyF
p2+7Y/PCbM0ckRX9qH/a6gpmobZtE5v+LL+D1tbB5T/ZbJ3MvmOIdi4geJeQ+qbZg+cm73fgAnUK
4200Ccu8RWh/3FlhpVRaGTkWIbii/QjrsYTxcoaHQjyZmxmnDuXSdW10AZx4uY63TFG8tqCLu8pl
9pB6FVbuYnqhMim+aA7mCLcsG9Tn+jUtmjmV9VXqF9AoVYsfdcDdhFeUwOehP0o+5KwUnVwVOsUM
gwJYjFhJh1VGebM0D9QAl7B1ox2c6d1WM3RUbkv6wG5Ckec6yhM4J1fpSbhQ/zUwXCGRUrETBcjw
qPxJ+RPnk/q8QSct2e8Lxo3yyEF5gBZMmGIJ2wBGtZ/OpeS/OJxsF90h8KBO8LUDFTkxUOrOHr5N
9BOl2DRDX9NYxEzz1bo+ZTjmx1YVgZyWnasj+AjMQ/hprMqZ9PWoBHTJOKQAz1sr8d+u0Ol3KaOO
LFns5H6NoozR30QyjH7cD2ZBguzDGN9DBK2Jem24yJmI06DQ5ajEh7WEXL/RbnSiCT73mdAw6Moy
gh4/gXbH1/KqBtY4DKjOOFGSc5MmWVRHNoLeTfw5QaPZkZMR/geBCWeB/1tuBVQ4A5qbjpsVwmHP
LyPzGS+XxjkiyaQ8dPux3XwovYn2oRG6SFi3PwNZL2A7kL4FKE1T3qKsF1O04qRgkMeYqTj3YUrU
T9bHbYUsRrxPS60AzxXO/0PNqEvHbL5uzf5m4+cVy3RO0EAAJ7NsbaSQrRxj2Rr442VC+HgwGzMz
gEn9OTJeNaOAYrtATMggFbg7XjQVGv7zCePsYNc4/1s8ltmc+m4SNAR8+QG0qJLhYaNL0x62Bp9I
TIQgBwU7NQztjZeyPXTJwiBB1kiJZ91NLLHNFrzTnYkVsH7If/L2GxH3P/dZjiz+ocako/Z+jSDF
7Wa2Tskygg2a48+5MOP44sFSE5ETu3UCGa3n5sQcfZKg8D87JENEUN5sG6ppmf+lOyeeyNFdJbyT
mSag2KFOhm1DL9GxP+FuUoCAyny+L45D+pKOpYyTxz+9vS++njwp/RDbeS129raC3IQmyrivfh9j
g5pXUE+jFEJ75qor0mg9vQFrmDxQWpHbLS6usfD24ijSOfuvJEQQpceOJv1W4b9Rwx0jBH1WIdc8
r1FvjDNKivwIva4TEYZv82kFzxblsgzxuxFwbQ10VoNczE/gxsuIkEZfHrmRYw+O8oED/2s5ygb2
FgxJxpXwMhY0NxsCQYePsP9v76rhX2/8hPAmcPogicAWW/yP5PH2xjxpo3HDNTvp5RGFtIdy3By3
hk/luXzcY7yJ6Bxx+sq9G55YlEGxCHFAD19IBYzInlSzP+FYG+pylE3dnlFF/fWXbnBEaLAJyVtL
wSW7Fvj5qS7FFZfrbL1bbFTWizIXaWNEv/sXRldq0tSmg2bo7uCUOfaRHGhr21eKrnCiGf+wVZ5o
CGLf6pMkdEmDCjmZ1rVaF+3jP0575pV7ioMHl1/3ZgxaHNgFvU8v7KXJHh+st3laE8nQnR/4abA5
dfO1NcBtDn7PXXIEaIOWGl1Qn0XjUGfGednsOQYxr5CyKDINvEW6HuhG3gRkkG+uTtDON1pnaxPN
hyTXxsnN95qsdX/VVNZQcEzAS5rZqeRxW46yS4dwzJshELJVQGEiJYp/h1bJwR3kJJxz8MMOLMdS
fPcPm8MEgoE0CAeGZ6ZkhrFtM4S1y1EpFXDWXImDlXVEyviXj4RzmsueL0v0llgn95kmh+whmNW+
miAmnM+H+kwXQ66sOA6PSgx3hbEPvybCQmo5E5RO+r/YJ6ZAOgYVtpAHgF6znMkZ1JGcARLNTZmi
e30mrHa9cBhCiz0J2lhR1T7vsRYBlVTfhjwzmPkGUJNb/aqOMtPQDzbXOrjdPwVwuSVfzIFGF+h9
zAu58Fz+VnM6xlNprVnh0oa9EMB4hhrkKNZPfQysewYYvRb/sqTRzfZVgEmGnK3sAUKYJY0tT3iZ
k+bv6uTQdawLcxA6SYz3Hmqc5o9I+SpamlTHRUwZYqb1SNOfQLlNFzjsQ9/0gvM4+evZk19+9ajc
t3xN7pzyxIHBJ8+4Wm89uOS5krCOX81WW1OHZZmjPY0S+ghN0Demi3TZEoXhmvXI2XWiaz7YUpXZ
RT/drHDYGVZ3HFVvG3lSp1gCoPqHTQMzubc9esZF1+7uZp5jESGHRA/fh1f7j/K9oQ4WFCG/m9Br
SyJ9KHwmozgzI0XVrFNGKo2rU2sowkJXo+dKiBCNehRGWNUj5OFkL29CX27BE75HfXtY5iT7/zsS
tuS+Iv83LQnFFXeDGsW7eLYtOSIPjaOs4MTxC/rzxa9khZRwFFyZCIFJFg2ousasmPAn7qiOwSeN
YvJKALhX7eJEoHv6Tr6YHL9vRP08nUe4062oetrd8ktnFREdMgy1Tp79vs9b7vBH6HAFDI6+nb1n
RACnFLNr15TTy2TXFl0CJN46RGpyP7VBIasTaGPvHQZfc/KGmlNNW7VY7Ge081UrQlTS8No3X8Ln
fkFEQFxdS4d0YIeWrdyYSIqKzRoPlDiAUoYAuo1eqwzdkbcW5MCoJDmO5PkuYoBvNAGN7lswE0/j
bsYOg2oF90lsDinE1wE5LJKGQDvBBm45Eek1e+LTruITCtjYVaz/mnKa6MfnqOaf43qjgSvDzsDS
itJHJjEIA/16yjqFJp/OfOHBXIlUG9+uZwZym08+5IT2apgxWvIg0ex5QmwZtazLRZddoIFpaDJj
pUfk9FWUOSMhzYOBXWwFPjI4HOi7gpKKTpHxHnEDbeHlEF9bDWBL3LEDr9ZzlMHGaGVz3VmAJ1V3
ZZBq+EU2G8fGZ+6sDeFC589rggPumSy7Ir7vxxUz44IdYYRHVNp6rvQxaSwOmVIBMiCmF7a1KtpG
/kZkkn91vDIGheGQ/k0LJjZHvPcBiFdcVglpERUThzu6Ty4KS1WF2qY+LJaPDyjk4WaCvYyT/MQp
GtFQXJyNBf4MqOAGm1SjJ4C5FQhNm367YIlQBYYqK0ecvhS4bGVkEHvYKZQjYNr+DElzyP0cUDP8
WvGXiy0wexEKPIkCOnqcXUAf3ryuI1E6LeY+xJv0DP45CqlOzPNXSQlbGzKC+Svngt2ySpagVoU3
GdG42gMXuASEdNqyf2IN/o4p69+fy3ly/ssWFdoyMcYtWx1JejWlU3lx6hWqH9UTRMmhfjDp7Gpo
bNrfq9cJMXdzg6sd4nCAIxqmIj0VENe3HPgr4/pJwWZQmkooMfCdUNvVsSaxj+93q7xmjHE/EBeu
Dsvwqw2sztUGycOnF8sw0t6CjclcJWnFpDBqXP34hsBK09d/S5+lXC5pGeVL7o7DSz14E0s5/2er
UxgNdMVerXKUQzTTj7uvSfSWUpSRTMQgY2TTOl5yQVcb23drZVgl82emOE6eiAjPC1JhMlCyWRdf
GFtdaU67gxgSmd0uxjf6lYMKTCDzoTDEwdqQnvRH2qXvVBhnOmNFm+XYh2C3gY7NYV7NrThRTh7K
YRLANZigqOFUiEReLNPe1NobsMaaJDhkJokyWRiv895g0VUuHKU/vK+CrVszcqrS8sagOhgq5grb
qU1phk9hYg2xnnJHE5FIrRCzS2i+vfVelNBmIPsiIsEsLvDFvxL8qiZRKnr1ZIV/x4I8LWfPzf1t
PIh8wslkStgdN0sCagzlhxQuW+KZCmHjIW6JIVaUblMAhTAr1sCHhoT7bY8YTWXqwCgBFbbQDZ21
NC0K0YTE7C8PinTyVin9lkO5HmQ0jBDxJ/2W3k8k2hFmFj/Lhw5a3e0uX7Yn7W38736r7J66Lxd3
a4xbYOrCpZMMGQa86OgGCv8VzFhyeHFtdXURiTwTOE9shKsHZaF9kbIKvS5R/3d77lIEycAokMfW
DyXzGxsqVKLF8yTcMuhqZEa5KNSdSy0bmEADF8ig14BK7DCRjfN3HmnjlnhNpUtiqAzuI3vOBnyv
cUxqtosAP5KfDVhXPDeIUFT0mITbfYysx8jpGeJoctqASpjIVk0Y3DkEiPSXjSCr63VuOA4nmKEo
FqzJlLqEETEgwGtEn9acDjgQ+5wXbvzi4ogB0ZZNcggamlInSZbaEqY5iA8jhr2Zbf0qbnMc0kZ2
qRCqXKk6T8XglAJMiSa/Na3U+4VzFPGGW/iR6T9Mia0yKer7pm9avibO70sC8b68FaY0l1RIZ1Nl
Gs1OqDRgzc5NB/K0aH7WiYiFeLdm3YL4/N4VRSPm9/1ZuuCIImjywssnWiYjh/v2yoMIeP9EA+Ne
fPoMbctrQ9tdOBDcIT73H/Gl8mP4VFBy3BV9L149XMenS81soLpoS6qxB+lp81qJ2gCHLcxPXeE8
9VPAFkCO62UNh9I7uC3qKhg5xr1Vc/LtF5Hgy4MhU6XBNn5JDKAFWC97JYhctKXFooNPzXCqACqW
m4hP1dkk+Hf54yX7lJJRqnymj0x+PSn1vRT/FrAz1e2NhWMvNFxr/VVxmDZnsVU4TsHfl4LxXe+l
xe/NLnlR8MPf98wF87CKAR0OSuQWVKv4ahAPDmwSldDuuXOedqjHaGu2VJzGm0+a1gPksfUboyRn
3DR2TwyK7HnT4kS0mBYampTltpL13cMzQjG/9uQqw+Od+mGOl+I5TBodLQUq1KxZq288Xo+TB8gA
+3StYxRrKZrxHX7Ik3wFljZE78urlEn64OFcUKW3GwTLMJZbKGpfTSa0likOYHlQNNwBGHG8TXZo
J6/VxZiByqnCNpq1bnqZbV7qtsBN3akU9kiPN2PEo+KG+ACGebBGmSEgAMDuC5utI3fQ7RSkrBEw
bYVyxtWkgenFflXcZuEFoK3zhqW0Nx5oZ6rjfn+m7L6Aml4zzFlzQUt8dBS9g1952q7xlEJ8OYoG
WNRwJVgN/XBsn2K7sjBHRsu9Vmd68nagOel73G9Pb88s0xra3VYCF1kzG2DeNkWbz1uc+6amIn/i
EMSaelMiECnzEoP8EUSvSXXpkA9ztbWlN7k8ewchmIfASE98DGMWw1P3klQYZcEabB7u/POy+imq
KVbeQaiVirJQt8stUu8Gd6v0L8594Vz5RqVv1lFhWLQAdpYS15EZCFqUkITDhVgf79ZuLK9LI6R5
JZ7xyUa39h8YTVIiuIRuB8WNZYGOICqelTtmH0E/lPJ6P+VwfE+LD+SSwSrytHqyO8tO2QFiGDxt
pY6+bnPX1jjgnXq7WMxVqSDnzjyXk+aXtSJcr7Q74DaI+fo3snb4uqo1eZAIcWMdNGrIc5IDdiZ7
M9O1WZixLAI3ItDte/CLUGEgfPH+EQCVpkzURDoUGIkb2NW6wRz+DV1Zk6MeRJGdD1hqYfPMyrKO
kQfLKuMD4QMK8SlHx8C1jOVJIoTu0D2k2wtauJOND5ICfILIKTKWLsb60YaZ+wssRxJGtSYNHf+7
XrQa8WdyawA4PQLHL68XKR81CIX2wSUj0FW0juZ7bKUEspSDjSQ1U/wCDYYEblGmWykaQBUHKhZj
OmN+gYdJApppR0cSuyDtARyYMo/N5UmUU01kT8lFvd8XfNqyaEzNa7k12qRZl2svJrv9f23RfpVK
nzFbUf3JLTMbUiFkwQv5gQAh7CfXcb/bLK2V9zdDIjUJbh6iKacx35L5QukxaFlHoQ9lhjU2z4DJ
Rw6IRmAh1SXY+bfbMVZC7LQBqC40gnpWX5KW73AfTsz9dQ8/PSr+oU3twvcI94KUWRFPI7nBk+jf
cEFRXafoRiH4ezl52bTB4ivSaI/POzWFisdd1+aYoun51IyxgeqbDWXsNlEgYMx8MC1CPpLXp5Sq
F01cCNEXXJgLpR6BQwc02u8gXphie5weYX6ugf4lBmpQF/RLt/LI2NAQPEAFSZZe29Mhfvebx5wg
mk8jMq3knoxH57qh4oKQIZ4WERGKeo1xs53dDor3X9PiKCh83BaSegDlIP9bCOuAM+xuCJZnG/1I
uWbwjXCmi15VjFagOZPVgS2ujQ/v56eZihT3tOtSJH5xLbD2x/Vt6jjIcq8/q7X0OWBjlOa+pRN8
qvlhYbMTge0Fjv+VEtN645YhR2Lji3qr8wGSGoScauKfCB5K4mTSzIQRPojPX+yp1fs+PRSwg+qT
syHzs8uxJjAOxmPe9oaowg0sljwQsEOFhOGS9PCW4Hrt/CH7W3RKLJ9qy0CN3Rh8pxb1pA3lF+a6
v3kPmwTIq9aNIn9qLhQ+VqBR3Jt1zj47PYynAFqGj8t//QK/4GlRSfN4fIVyYUYcjFuiAJJrW5s/
n7hrlED+xnWd9lX6xZ9S6/zUBiRWC31D+4yL0Id+W1jXhkfZSBy/9+CcEZCcJ7gOCWmJFrggN6qj
KuHnPZ9TeLR8IQTC8lk/cXj2AtJZ27hgthD/DdegClJmyWmA8UChaHa5oO7s+i3rVww2gY8QTe4u
VVnNmhMFPFJUDKWpAHADIr4sI999z381AtvcGp/bUP6m6Zw6/aL27X/tLhlmRzgtFR9e8A7rRW8t
mfmzNOnZ4VADlPtyiYvfs+W2hzM6+UVEWcqEye6jNByIfO5ZOovcMar03+YBYYn2HS37AzdxAZpN
4AyYovsR9Vvpb1Wsnla8lw9CpAoZjKorovBjY6MzbvGiAsf478rPOmvLOw0LlaBh0Sd8ouCZOPXD
vtVLH+biE60FoNk/YV9oxD/atRcMLFg+/wJsxl0NtG/rOJ14ezOyi3joCnXU2cpEe9srhzg/4XvJ
if7YvU7e1aS9swrU6kQHNRdUn2JmTFpfQSECLYQXhGWWb447qWffA4D4FWO6aw7EoEUCJOAL/Wmj
EKcuiLjSffC1Uksnq2KSs5MWfGE0H9IS371U0c78y9R2vyhWm+DF/QIREmi+A7pHjqR0qiowzU4b
AmFPzQZzZL0/XF+nTrBDD+yQkY004XK1tweLxq5P1dmJxOIiimkyJ3ANRml9DbVe6vjW9dWWU9UW
Q/+99r7i9YyLe1O2sHFfmZ0hLH94YLW0BoZP25pDIVx2Iy/aZo9CxmP7nl0GhfX/+CBkj/JJ7FwD
POmI74YO9q9gsDvswKc1YPCG/C/2JJQW7Loj6cZoLDgWL6+vxQKGCpELhI8Wq5/ZVq5bqp2xTWoe
V6joxEXdwO0GzvcezCynOAc0gScCHJlwVekOXyvFppyCdGdQWhpriD/w5L/Pb+pxdDS4JuXxzhQm
5+hWRz8a2gdEb2xCXVHQJkq4GcFVNMNQdJ+ke01x/yiSH2HtdlhQsTAdqT2xCsbPHepsjCmDQyvk
u1CFnM6qcj7J2RBGjvkA2nhxDdCMQ1NrV+Kq0z9VzM4ctw3bQEIVJb9liWJaX3FysLN7bXbW4Yyy
9yA1M3RBSQuEqyrl0d+74Lt38nkCP+2euCYzbHCiEoUbwDqhkeiIPcP7HjzgiBFDNRkhXNsd3iBK
hs2EeTB+SIieBkE2LPvn1VkVd6/9fvzygsPTEbWMRYq0QPo9aZRdexav8Wj8+asoXfwPvBMI0QsS
rtSK4FAwQCYak8IU5Apw7W056JyGF6pdr0L3lvd3gI1QHXDI0SdJ/PmAVggZd6h8d8E5gGPQhatn
aAvNnyLZRnEC6VZvcQwT9oq5BAcj6OOEb4iAbSXlANQgGXJtBjyUdrD04JAlreh2FTbI4vJp42WG
GevQbf+unwIFBt+3RFhcl9yFIiGWzE+yIZS4T1wGlWbe9kKfiwk+VnZB3FYHm7mxoQZZokBxYJP3
vVfwcY+VUyXN5re9Dbpl98rimFRAWAMorJ4aLeiNMJGAQJ3lmJIeNADNsz/a1CBTPbxy08ovxR8K
aTuESZY+9oetA6jdMaKCeM9IY1Dbryd1rBfmOVr3n0CYqFK3GDCiHz3AGBJ9Hpbu2F8zXia2Ryu1
vB1CS9XnyhbZo+fdrG1IrAfIKeAAJMfLKsuj4NgPAZEpCrDtbW/LgomcE19tGHHE4tGOZNjNlclP
cEP7JKpz6pszb7cgy04FP/AlLS94uG9SkMl5ZT6ATkFvfJBViQRXgOg9f/8OWCtahNQyYoCjPU90
a0zUuKlU/NFBskdL3vglFzCHVxyIc/H4Py7JtIeCajoE0GSxdFIxjWNNUUMgRFBXkqxHr8FQrPPF
GxrGK2l3+huBtGQs+7bMgEuP9rNTTvanI5/AQEW7Yf/Gej1tsQpNBrRecCaNYRxZk7cPE+8Inp3d
76xqxyXRWqGgLKlDAqiogP+5keMwIqDJqyKfEfx9R2AjvmBNQDMppflhSSSj/MfHGTXHVKsafs7r
MdMj/4aqxuAGeD2/suHZnSobyqO3rOm9LXLFZMnd96kbhkt8W/q0crXnh/jevayHaPat8TlgUFeB
N+tp03iKzS6RbcjdNiAtFgAqf3eoIxH5dHNFthY0E/AgbWUpyDAvaKxUWoLNIJPX8L7pKysBj0dH
+YPQazTuMJATIVPXUXuLkSFUDfQYUZmRO31P3kNqG6A3Nwawy3v2VqvlnbIuFozjSSbO1lfNPwG4
W0jiitGt3rDOKxZ/1AaVyue79doSMQJgoMj6FjjnOnOaRPLHzj6ou4UIUcUmTkVOVVcZ4kyqoqTk
NYBW1N47aTm8VFqrDr9Lv8YZVH3WS/YxqoO2vZgmNUJMpANiB16dQHxN/geeuob7cPqguD/CwAlY
zjr110oSXjffaH0mMHxGC1P/P9Fe6SkKY9P/OCFfW+phKMSPvTU+ShtxeEAPFWcfHs7jFxHE2P2H
OsffJR7G7x9T3IpLFrnrFrWlKyQu+lgNUgMlPyzg+JxFrRTAc4gaLyr6mv0Nw9Vi9BgT73l2URjK
KlKrxCS1KSHpvU+NUYYnoYca5PJrHyWTACkeUV6elBS2qVdhDk746HBG8XlYMmgtfjBHIUxCXY9V
F5eMg/bwyJHVezKJKiwdsir/EGGjSFWf3XXHuAJU1HG5z9vq5cyYBUwNeBWunFmo0DltzmCcVBaZ
9LifZ3VYusgy3C2pOrBdtHznhgPQD1y46hfgFAAnC3J5FtRvIJR9Q1NgFvrxPaySGyYwMofaXUv5
ArkYHAukRNxBd7Mb6JNf8/AOLxGqfqpxsjCCR+VI2JSceU0M/8GDbk2Q96mrEoH3Y8kyDpS4KUcO
xl4tGn+uj0au0z/W1/9g7ihDFr0oHQ+TFuOmSZcSybMrLG0oeuWLbTuTE8tryhPVBKItCqnJkszT
6bJ3Llu+NKniEtQpPbT8fVvUsX0Fm/QWIQHwtUb4Lw+nLyJpsKmX89gGRYDxXOomONT4xKxKbexr
dTjy3RgDMKxy1USQTdtDnbem3RujdvmMU3zFgytiJYXVPez6wVXUqsdHQgbVtDOii2eFhX7ibvgH
2ePNv4B1IPyfcLSNO9pMyl/7p8xuvXvMMOpFqaIbC21IORSgRwYxOdkS7vyB7p/mkiVl0w+U8Mft
+N2kpUR+OMo5cPkmhGsdTO0/Ix2aXiJUwSho+3EMOZg3+t1h200RcK5/2pN5zLiaCbxThN+FoR7K
2UerBqQaI3htInS2CDsRACTXyr97FlBk6tdFpODA3ZdT7npFuDRTVk8ZLCqsHnMtwZ+dQpSbma+v
K8CCq/5KobN7aABmTkUCpQmQKVuDj4l+1h/8BgxSiFo2+Ixaf20LJ744exRM/Zhyti2sRHY/8AaZ
mXxj90HGJ3bg3WoOQiIpaEaweiZcl1IZSuS9HLIoVYGO/Yzwk98mChfOa3JrnjrBjMmwc/aFRHD+
Zicf22k9IRwgcqFv6ypc8TopJheuYezmDdDou6klBocyShsmB2ryc/OxlPwfevyz+D8a+i/08auF
faU2czispO4Zlq0nLI591hD5eDr4qI3NT7yyRlAWEBPSnH270+W0F+xb7eOSNv6W2iRs738XvWv6
zH2TX4cbs7zbYrSzDCdzaLzS5G9Ei8y6yYQlDp5EpNQ40EdQsOB0/xX/bccgHomI0DhT1e4j5dNz
7TPls5gY818N9VHlEjQOXkxqVCW1glizLIO4/OYDuBnocbrganueHB3O/G4TrOeeL7wg7bxER/Mm
lJ0kV13tn4PzT8ridhFjoZDjqQTmC1dpD0+o6PMnWMAb1TuOCAP3oIHGpYDggHmsFC3Es07M9S1R
W+nTk8fLPwb7zpl39mXO6R1J/L3Xabg/p0jUodQDTGDaRAgk6/5DF8TG9mbzENofPpEq8Sd7lM59
W+j2a1qGgYSqqIKAesuyETr9ZFKwSOJEEagwy9v8jq6+ik5CfCln3x3FqhMEBiPT2QgL/ZaPV7/U
cllSskS7BphaUlnOXq1VnbWb2hd7KUsfH6YQr1V3V1I2SNQ8ylpj2+JOWEXD0JogQm3IocM63Bs3
syIBCT37da5g5MQ+qoznHxZMjfXAFiUVOwN++8VFR3VymMPKtdZshsKoe3FoytBtPPawsj2LgeYm
M9tq+wBsM3dF8aund4KoeRIyA61YfRxwOxh5GZGwF+FcdXvvRUlQTc/KwSjVzUoyZEh7UMBAr+DH
pGOSSGPnOZyjOoKnSzNh7pEqFbfaP/tPvk+/w0fBLHXMbDoCfCpsylFXNQW1o7oSDufXS5pzYs7R
hHP5to3wD8z+i32p2JB27XpjLPqDZejcXuHVQCfhQtXlzKGdUxwxhaJ5hvMzUKXctwIhjZJn7pG3
e6NDt+r4cGMyHUqbFf7d7tSdGCVEA8pynzWN+cpDvtVxVGiQBmZqqJk1W3e4FtklV0VR1UI3QsRa
ExHS7GsK1olB2U8n8S7PtoJMY5zvQ4hNnZMZROA2vG6DF+wauWmCCmMSZ8QOFPb02eN9skHgFZdh
Y9DEmECGNxg7qNDlnPWJqMkV7QnWOJj0r0sXL2Jf3jfBP7b8JLjNNwVQz7FlI2ofyloCDtB/mc3L
+1/xKoBktu20H0ZExwe22l9ZHgGI6kV3y7YCApD49l+/AQejccpvNC8T1LGBxXm9tsHPpQwcAliC
LHdh82c4NZNPr7ip0krje8mdXoTupOzoZlYfXDkOQMpaoDoTeW/MwTTWbLGn5wURUR9K3Ig4JimI
zGim5DNszfcZCPoRbvwiTgrIlwwGSV057LnkA4bPGa/Wsgd12aAFd+he4DeQH4ehK0KHJTQRB2yk
0asVClG1DkuRZtHNpu8TWlGPQeAiwQU9K3eVfU/zFZCy94l55pS2K6F3T3/mSNKfm30I8DsumaHc
0WH/QtIlH7l8DhJF8hhwjpYHlU2dGwuM9viKzvIpVCeXt4sw/CVSCgS9CP8N++A259/ktY48kXfr
F7t/cNa5AR230WG5nJadH9LLWrabJQRul3JgflbmNpl9MsAB+WUEBv1omWp5jqPvkxTdfaQk/R8O
7W4LsBnuozmoKNuDwtuTvlRSAEo1bsF3zB6uDp0f/6CirIMJc4RG/iabVEbbnE+78xdX2gSyxZEi
2ZGxiMuVkjfO8v3dlPPbZLRx+PxC1+exkz0X3MoZGnRDvwWu+6hdBsGIK3aEtReRkDfUSZeqe33G
rFOsWOxCDMHwAr8CtFsXfMH7xOxTmfth/XP80cV/CmTIeNsO5081oSnVoMH8lCcffmw7lgAlgGRw
WBokGl9rGfGlXMVhOdtqYZ5YJPLzRxClphL7hfHFNB7GradaHvTRlBHxbybM/PLadi92V1tvk8Zs
93TMUyv0HGcr6Epox88cPT8iTBGCUxCCvIww1isX0D5AEgK/8hlTE5dhsnRUwYVSTzVqdji1rVIi
0b4cRt/NNbaxN+A+KgF374232x7nY5zieUBxxbYpwCjrSKUbNeDxYosj6GQOzdLH8dbS+SlHFmbi
MZxVDn3674ewgDr7j0DZ75+z+JDofZ1R+uHIXUPYH1hVw7YJweFhqflkaXQPVG/ZB+3ZryJJuiMv
YtmtE9Rthk3yHedSgc+VW/P9PWwWCOb78f0kveC8NQ6Lyf9vH/DvnHFtFmww+mLkPd/OA0CIwaAT
1ZxAJdCqkz+XPZXakRPVeSeIxilWbjmR/VhnoCdLGbSr9GKbg/ftkGYMNBzMl1J6q6oI57v8pOfi
/4TJVnf4cShODA0J0vEDleqdbR55JIlCopbTU6XFvud2zHE6ZCd3r3QGv2t6YRJXDGEbX8vPIbud
Cjd2L2HUMjx7DKhdlFf9D/YSIS7hvO0wqtInk7RTITrJZpB7HLF6WLkyUzATTDwFKCicGZlHXpb2
qRsvgRSZ+/ObXpSwmCr4udjaN7ZtxO3ccP8o8vOrdy7o4ZZzTr7JZwou7sT/BTXvMWcw5mxHQryH
DkTpSBdwdfg4izipHhCtDkQkDQU0lOBN45Y0Xc3iJiMknTLgcpTc9qgFeQqM+vDaH/qw5DpOg1kn
bojYTfnbn28wjPOL5gIOOu6zQ9rKO/6ms5UhGTTsNMfnlpYOqIiCa2CrYnCsdqEUDwdcbz4cjXbv
TV4Cgo47QAejjVfI7FGn9TgdK6ejbwP3vvO4OiD+uYa72Xo3RzVwOiauS2aBaVZTioUGAJDO+RTM
kplv6hbUdpP8haN9R8u389oC9k+fnnVHjMVJF5jlkKKxS9aeHDKpIwrw/x1Shz6tJCrZsWoevTPE
BuzYL+WKuMpBstpX//Nssr58n01WIO+ZHA+M0z8bfE5q2XOvq6J0Qlowb2SE9InzmTcmC2+UVG6d
iWjvk05bNilVmrL5ReBh5X4d4I+BwsDmwSqSUgN2yAEbZFJtPvg/NaSYn9EVTkgJLhprq7ISc+op
riP/Vbhi3bvP/H47VJbggioG3F78Zh2ShmhsmWkPdb04f155XfzOjeF4TbXvdSxzpzYirGTg/ldl
2WRcLuWc5sAk1Lp0U6MnU/T2vpyb3iRw96CxFz4COEn9vdNxdn2Fnc2SXnCJ815xylNhwraMeFMz
f90dhmmewe8zmrar6RCjjXCAil3MtEXJWe/hZB4bGHQMJ4ZNEL3WKkzA95JRZoViHu/nrE9Ra7Ul
U5oeyRfMhx+OeIoLXe7G7+NTjRZyc0sD3c1d7+iYpkUuxjnlD4DsxNL8KHbaKZomG/oSX115e7UB
nJyK1oq/eeHVVR9XB/lZFV1vw4IwFnTn8a/UucJL2K8geSExcqAuo90AVeqMK8rBCdP5sv+hjlDu
UIQOnA4Z/5tFRO4NCbkUDYRdWokiLgHV5dbXMncZ/HUseKqkxRNO5gRrjL+yRaNNfwlbfSnTKWbX
5NQo9PYRyYdvkHRWoazkH88erc0dj7T2FsjiOchwRzKcMEt2X/+DN12tTIWlIoQJwVrDezJQkEEB
/qutpbJ9tETDnQ+0CcTZEht/VLnFidxf6efYKXQfG6EzNb2UUvBuAoYgjDqV2amYQrQreIb1ZEmP
6ZXVEMijlmZP9VGxxzXdEe/tUGRBVa/4tBj9F3S+uo5cZ0BPUaID77wDUwUslo6ibTk8ktAlDpgM
QlT0uokHglSj/VMj2pamYagnjHHqGkXTgL/BTO3onE6BSl2Cc0V32zSbumekB2wUrPBDIc9GcckI
tATxfUlup4vimPjOnPhy7zTNAFlVy459BmTqzE5bVjuTiTYKtK3mWMdamKAheqZkHjFgYHsWghSA
tzC2Z4BoNdQqucrn16W2GifD7M48PHoQNT3hql7JE32hu4JLxN/Ox3Gj7U6XqPZkN3+Rbc9F6YvI
Vfw3Z9astdbXr35YnTfjGxCd8G0aux9O5RrVVkB50H9+0EKVYPm0Do9T+qphTtAlIFXEpI3I8uks
YslsQEPtkj5HMbWu8QB8pJq7Q9B+f02ME3ikzzMv40l/LcdAaKXHXGRR2EtBfgfOC0o97j/c5uxQ
PuprSRS1pco8DQWmA8bebJHHj/zBixJeCITdWFVQu6+oGjptnAnG0MMzLZ+nyYu7Y9GO0FVpQEyM
WSwcoQEr7d2j4Ikb452/Qdr9fa7XdIYCk378hFxQyD5kKD7SUmsShbcAhc1EKmNjINFCqAIHQHq4
v7/vFB8BpzRRdx8TEbRVKwTv8xSL3qpsSzfXa8pPwV+ZjDz5zkS6A17KiABMHBcDkKSKa2Ob0bld
iDtlswJikgS8FxcOd7L598wuLjKbViZAX/sA5Ady5A2xK3g5BnVl5+DKThTTg/uEs8KGpmQ4kHQ9
5p3gcGy80tRqBeOZs9gKRiUHtCQ6dhmCV8QLopmdhSrPC/GxXc5QwVNp19ETfQCjllLOCss4ct62
rRoVq0aYaFMCon0mF143V6rr6ckT54oEyMJpmuGVl1J+NP/cG0iVqN8eWxdoEGznY5bBI8AxE9yl
MgI0V8RhE3D3CLyh+ppE+05S6sWkd/aQJZdll7Q7UwNRa2+BqjflNZ1c0Hfqei+w1u+aHlsHTcRu
wF21NokhwNhsO5TF7HIlfpwJyob0rNBmZ1YdjbBykYkX78abBPItFwerfln5KXcI2gLY8aMaUmRh
ACG70oM2LpC9vfRo5XSP+ur9AAn1bRC3SETBadT9S4cUJwXb4W4kcOSbbnB9KXvM0cbrSYej4a3x
kMkpRHjoUuJvhcboFeJZ3WxM7UhGrGsi80cwwqv/N5wrr0mJz1u++56z6XK3Qq03opE9n1v9q7Kn
kRJXQe+sqd6L2Ig3J0mmhaFLMyWyCnmXctN7hHG93M3SjcTEYGRXATULvHZCxotSjqE/SbG6/lFa
aqliEp9TW7DKW1UAtaGq8ZItnnVZr67ar/6b5ruWhLFfNUJ/kjSDl/TXhDYau/dof3rJDxaCVghY
KHkHNvWj6XaTfdxF4MPh8K3ckE34lE7PupndDRUVLof65sRoUAfmC6XWGmX4hgUPyAljyiVIMFjU
zlRt069DDYxHUmChbz84uQLhHSlmqHvPQYoZbFwrrvieB01VQCT6UKM/RZ3z5yykgi1hQOucVUd4
QcSqBRoyDJhwg9/MRxa5tTs3lDemPFW8ZnpRbWCWSXzyLfDP5F9KsNfgGjYYmqzMyhypBwRjxpDP
lR6EgmG0vr/ZJuySxnRd2iVXLtpK1qvaY+eM8G/WmUv67drFqMa0ohM1wutlOhkTOczfOjSNneAg
llHFg4iVbeVNJENFg955nJEeOyFBAFcqm35Yz4SqDMQ6gGv5IsafY06GjzLW1kN2yJxWZCdfn9HN
PNN0ZKmrC5UkpioNJxlPZxQlDPW6erHyL1avwxGVaSM4qyyTqj4RYa++xRKAHdwctEiPDph1V9Ik
LdfOeyGhwr2RWHFAFo0LE3q6n4jOXLX4ASSDK3LWv0Ry2ksqWfOFCFUuab2riMGElQ1UQu0yy8uS
r+mSFDx9oulqyjwh+/O4KJ+BIrTbzTe1/VCktO7NojcnnAzUwWNtm5StV1+7c/H+6I9XJgfY3Xre
cqhdzn6+KwU+MdmQ9AJIAFZDYUfynRumZ0uQvLzCP3KtFaLZ+iCvC2GaJuqN/jPrkfeeHXZHB0yl
H4knFhS+axtzQqaKO/buFuAWw/BfO2/qVO2kTF5sOEWbq61KU1PPPQt0j6Il1lxQ3yoIlwvSmuhM
q5BO1K9gsCku83UwPc08yKgd03WdXKhk3ikmZ2avxCIVH70rH8VEGNTpPnoBZr0K29Cp3tVcuC2v
YFdwdlDjBZU8+sd6GObYT5qTxxsKvlZdk0OE3bBafiFlW3UnOy6J3olC46mleSH6j/YUzkpvqOe6
+9Ch4Yg5k5ABGHhTeNV1EOs1RdOp1a8QMqdFJpf26OcHEwXUBufudpRUh9OUSSv2ygkGI5ZiH/rh
O5RwwfgaR3dDa+b6ZFXjNsuk3udQxVn3Bukq7w/EsMVgqIH1vcZ0FmScWp1QGkhyRcspsuLdlpi7
GmZyzfL6Knn5VUgmowileJKFaFSqHfCtymbpex3wp7ww5KQk9oK0HBt6xwxtuH8OrSiGkYYYIu+z
hyCVeXwa/prtZtQPmjEVqWF200TGDT+PG0uqkNHin7uLt8IOJ6PtrhhGRRjgylBTD0zA0Xsa1Evp
xPhY4YP61ke2b9vjsd9rkosrRbrD0f3219AS9/2Fjyur17vp8h2BnrhfcocNf0LwgvOnCa6B5f+O
9Y+mij6RO289GOtTAwM6zqEd5340VsoeoY1OzBLy+lwIzv/TKqq6LcDjpTyqn+gaafWMuJ7jv3W/
fHHnieTgBuPaiYAX9u5fFoz4OIX6ofdd4mMrMKMYcfvbCSxMvrMRilz0ET7L5Oij7EOviSzwEYPs
qqMiiBBXzfpNijHiFLsR+3J6+wm3mPuDDdF9ryQ2bBBRtMlKZzEehrAcqHmJqNl10ngsRqisSbV+
VmN/WdAjbxRpVz2WOm9o9EJIG3BhIQQrPBflti+teCLVkG/cx3nz3jOE5PUC41d3bIAtWSLDqLtg
2yL5aQSpBbNwtZoMgyb3P9piHbz0OUBCFwr3Czuqg26S/ZorwIv1NDmzZQNcwn2E65iI7DQ9EhaH
ASANqHDvDzF0MFobw43kMPII8moac33yn/88V6UVFpVVR324Sqg5L7A0Iky4PPX9yNciemZ2MSJf
smFBhjx5o2sgg83daNOX+J361OiyXMGbWtPCdHPEmJ8Y9P6O46JY5vk6CdC3j391/qIh2No+z/CM
8CzFIiIyzf/cnZa7iuOku6r+z8uFks+CB+Y7IEWPryLC4nNNeWWflSC1Qp7l98BchyJ6Z9Aqob9A
JAG1T7CPzRlfXJ16zBwSl0X7H66ezO4+J+MVEIVn1mi3ieg53cgTX1jDwdcCPYLD3N0PfcWQDGD+
JhcZDcBmZ16JM6v1WahgQtzyWvBN7rgmVKkL75N/QxWvY0FZQ64wykYu/HjFPCY6wGSCje2fQDLa
4AezyfYODzpupvxl2jXo0KOYycLWstVRpk1HjlC2y4ntr/1Vj52ryX4TzK8G89ej12PIR3M2aa4e
jvIFY2L5p/ajvdb9sKL01WE5hJCcC2U1Pkk1yLTUx/2bx9WPOrGZudUdZLi0LShULZuqUGcj8YAR
GsWjB6c2non8qAekyh8Kd0rymZb5NE+iK0O33tjiOTmvcL8n3OWfh823ii01NmoG8Jjt1ZHKDoL5
nH/IB9AEgw35TTyEjyp+vhzUmHgDpGJddUuDnWpMGr3RuSy/CqxZ6iX2p03PPSUlXwK6dKKzyRB2
DFnD+UDyQiOqSzkGBekJpFWOT9wi39aFe8XPpzcesza8+1Qjjg4VVaZEScjQOZUvVjr8QjbkLDJ1
FiMrlIQc9gPlPtrCREL3vHjQghDtfJIHIC1toLe6qbwOXM1a4g018TNmCMOKieojo/pfBsaGxCr9
gC4YgFeRDJtIf3NYDWSPrCNZSlAnfrmivkL1gWIZ9IgJcr6I3HCiyYcrcMougFdUpzV4Hmt4eXjQ
qctED16KasQGOizAEOHLZw83aAmnzytN8jwPy3l7TSrGsLMYWcfWXDzjw5v4uAvODL4msdCCh6gs
uFSHX5EdoyXpU87KDThARdDRQbuIUagvNMOMNViOMIfzsO9CC7b+CgOJBlEhqKVLzehDEpChUvg2
LD8ZPDQold5SiXq8CZwW60wmp1eE2OSpNGcEQMmEcvGKMX0JmZOblGHqgjjBy1ow8uU6HtRppLcC
EynqfV/X+m9Po4bo1BCPSJsSU+GwkRBxPNDyWnlDK/VTJZNMzsXJd5gfLJUp5mfTm1YVNIFLmJR0
mLy2xEyue1v5UrSdYPtXVIeBt69nqjisuMJJSxYI8VP2IOo2KI3BsxWfGzcpPi711Ilf99x0xdmK
awJ1Cu/iYlpHSRphNJWVcNqusWci1NeeDOOGnxm+tXu5YpA3ZQNbPeH84KL63277Mj6TYX+EG3Ca
ThBvBgxweJ2WLdwz+BNfOdbFlibmrS1vUD6/VZhIy6Q8i5M5qyHfn5IwFZk8Vgxvmobpd2T1Hdbl
ZUi/J7HGw50wYaeCbrp2sINsjYJRcrcOEWF4Eqmn+sQDBSlLZYfPjjJJLKWp0415EFplbKkbCFFw
iX+uhbt9eVEPC9N7oaoBe5NlwkKvWa6Ua6yGlV29Q7pBxx6H915/02PvRh1haupLq3D8r2VChTfZ
9t/A5BL/SEGwfipTeDyXr3nMGAhYUqmqIJpacl2UNPA9yxQD/EWYxBunPSiyVhkXUD7odKP+2zlQ
eMrv7nlrLgHv9GdwoeFROzS3PeKgV/kcUK4SVULej2Ohg0X3dXMnnVZedwJPmjcESJ4K4FpGzhSc
/R1wQRH6vT0kkwlVOwii+hZcT1fXnPml1huntgK+9H2FuAbzCtXJtfHwCwkQF3yfzVVS/OZp8I+4
43U7ewRyKAzCdAJ1mpsQA6gsIO7vbTIV0ZaJAP35Dz2IdYh0yOM2weV1wnZdZoV3TR0ZG5lo2LUZ
Jg0q/BJFb5jJGOM1obCvqM2auDYjr8qwMfgI2Fewja/qmLSV+MESTsglfvMkfW/xC0IFCvvVOo95
jj3Ib4H5z2UCl9SfbPUonNrcn+r4FKc1XaE6kj0Y8q5xJC/fFe+CaVm8rm4ke/Vw5EMpEoKAG5BQ
lUX3f/akvdFyE+UZDjE5dWGc8skQXkKRRLTTB2HR8vMvDKEohphPjePZoqE5f9SZOWgMR3oC0m1A
XynL4TGZaSjM3lkaigcunZymIWf1Fm5dgT7KNMXX7p6AdEbprY/OldhAgOIiMXY5qAO+Ae1EfgMz
qJv/fnKnbn9rCWPl34OxZB3uI+axefRaxOw8KrrHlNf7Yn6zAy4xgDILDJcL4DcKSdRSSBCuxeX5
bxOP4tXdbIZ8GVnQ50DinzyKyCaBlNI8RXmM91cSjnfbvIJTbYiTMbm2N3UguF6XOZIiRH2avxc2
pVDYG7VmdqWGenoQg35Z8LEwUxO/zOXLll+/x5xheBibK6hJd5mIN32taOZvwXMyniA8YkXZ7VdJ
HALirtKvhvkQHVjkBCiMtLOZcBgeNI3dZWTAq5CTmbJUbzSkZ3HoXBVvQD0Pg+6gVn/ihPReZMaW
wPlKJHvRaWYi1/aU222Cld3kQGeULyDM7q8WawKNYWO6G1QC/DVM0aCs5pmLfzKP4mlbgIlT6wcS
sWjbIIB84jI3ygZVFft17/MiRJyaggX88zi33iJfxwLONNpnfIIOz9/9sR2GJceB45a6HfTwjx0n
39Dap8ch1HXqgT+KNiiiuQy9xBWj15JNUY/N3izKFSsGl/bPeWDKZp3n2Uy9QRG938aqoC8p4XWC
J0UPEJj+axJDKaIY54oek1LNFHqGGCbND9pxTyvYuCYB39ZNF+x1ZEPdTku7iKJBGT/PHoih8Mfz
PSc/IblKn3kRo+EscBT3RFTP0rjEbuBHFiIcD3JSKiyHK7ry4McDVjACg0h0pmF318/TGXnyr7lV
HonEjvwgCSfHZ/veqoclQDxvYkvs2NiGdht40YRJh4anjlc5Usnmo4dDd+2hH0F+1hLPCSLKxWJX
M/qWe9oS5c8rWwmny1mlNcpO1l/rQ4FBiThfvnAk1yd2IcaG6+wurULFJNPzATJQqojmd18gYXJi
tLpINaIAuvt1Ysmx2e/PWw3tj43alr9QRT5250g2lNVxVcnOBATbFJgTMiSC0HzCg711aTDxkqlY
mrQ+frLvIyBQRBcw2yE6eX+v+4GSYkWu3bxC7FV7iA+kkiVqN87WREnUaKu+Vvq0sL2q0SSQ6RC8
u5aP0UBegMZb8kUIWGUmkPeDHzRdH3mE+oQRmKMePYhy6fWbJDuSXJXYivJ4P2pi4JbsbUrhX4Re
04ASzaavBG7FF4Fw8E/gYGafrdTprf4EwAPr1PPlwII4QNz3ff1mWXmhGup8yxYH2y/jJmRQatgY
QrwI3SNuwxnCvRZF0RSrDdqOxT0Q7b784QDvYAk+1IZrQlUaq4wbcW23xiCzccjHWKYeyF7fVvo+
9oWMPMi0B2HoiSY8KIWnHTkDUQlB51IjF6lU09vPMY7VZNdAIX9j2SmKRVY+2EJtW/WSNT+vwMXe
FPviCX36jmaWFY4kHW3Kcs581SeaevkbmSRXI4Jru+rUAbogGmq55Pjz8nDppJhXeuNJUtCkSKiF
7rrt8ZsB90ZcXS2D/+3Fc9tup951CNMplEHV6z5ys6Y2lJXJIL9D0n7hUQHag4sKC8nK6eI48hIU
Sit48rAJQD09f8cZxJS7m+8oCqVH2V8dWhruqsbxFhkVkhNFyIQg+JOv9yfHkCCJOXMJFJvvPLnr
n8HSfPdogrjUWJriTiau4PM/IChlD6MB0qz4lKBQjcY0qqSj6vNHMWnbbd++Zx8v4tKhTAp6a1xQ
h/RnryJ7ETOtDGbNbC90AQotovasngIADex41mKHDT9g9Y3zzCRFLhLB4OBkE7tWuamj7HaZSDh4
mvfnTXIuoek1CYjEt9iX4bx3SBPRW6md3qjrxnV+5OAkOmIO0SV5tN1yx/2lHKunsaOzT/v4alTQ
YxeXx1LTlv/PmGlkxstVSEqstQTDq9eGfU9HYgpARXm8mZRxjA9XF4JvkNn661Lv0JDuL79mJZce
SEAAuIlGx+GX3Ye6f5TqZjZwhHX0GLQtAHPozBAuB7cSZ8G69qDXqMsv+E+YDR7dWJ7bIDIXoJXk
a1bbRM+c/XIOfLaP636An97Aw+wH40s5jO4NWqoQ456Et2DmkHk7iclE1FPwIb4ncnsCdsflYTFe
Iboe75eZ+0NbSNyIbkbOjwZwgoMR0F6axBRCl4EqXKkLoTBa34ZLEiKsYfuCMb+mR2m6v2H3DzK8
yRSXZnz4s3+SdNPl/NvKv6k0w0zd/xnoJe6MUl2BJ9jAVsL7ot2HeWbSJAhEeRL1xCG7hxtwJA98
7x3d/Oa/lzLVjO/SSkCyjxkFuMjCv7a/jllFlZX1wbkdsMIRP1pgck1d4FEFr5lejJHCYP+gkPBc
9N07X4oUBQb0GHTC/iLI8Vsz7Ds/mXDiu8sEYKetGeRYhew04uF5IYazRrcQII+2OgljaZia0xJy
fHI76yrVe9kd96BcwnozWUIFFzWdhUmi5on0XbtgL4BKkx2WA0dEw8C2Qrxs3RJ4wunbgPZNZ8oJ
lSCCkXrMrmdz/dG3nz3ag6/iunIAz771Y09A0/ObW9Gslu+SgsmlOt/ciFoJ5y0Mw2hXefTZeIC7
YzKCzl0gv9+nxbhk/FQTbXkCNOgmEg8m79z4FFZTLVbT+tOFjTI6rU/9El2re7AiDK5yPNEYnoFe
9hIynp2FSf+tHACZvXiBQB4XNNx1PgFJPryUWnCumJl4dldCjAvUx2jX96flnJoMNx8fJni/k/5D
KWLHMfzundWZh0n6uSlabd8w7Gxat1fae2l9u79lT62ptkCoooarrMvuKGQ5Ymcmm0aRhhuxlpRD
7U5XKE100F5FllZRrrujlsi1ZnAc1POn9r3ajoIXkkp5CwTOLSt1HDjE9LiYz76oUhDDnkJGoM5R
E11qxxo1nLn1QTOoEGdyoc6yUeZ5xtls2BuBPeCXF3mPT2ZARo6JITOzPkLP6HXYtGMI0Ds5t1GK
4O7IfluRu7MC5NhFXVYshOZX0WHCb0m61ls8eHykWdzMhCgM1ALW4NjRsjUAcvIrNofTG4ZeuwPu
oeCfJ0eQfRDI3Sg2tOCfJE6oVtcza9xawuxkrS9Jc0p/PW2fPTXojJpb1Dbqo/1VZYTpj2SMbmeE
ppt+u326KjZB14Nn1XrG5JmIvL5/i+rio9btSJ1t2IGsbU7Qb1Vvcnd+zbnLWCgQA5vVjSayU1aU
j8aa0LZI7NZ9fdck8XEGMh10LrgjKxY7WLzukg/sGXoxS1/yMtOhdyPwCvrFZvvZV4aKNzJdYG/r
3XIIdvr8lvvopP2sr5bAuzuwRg+pTSfwRROeZef1mI/sEXIRoFszWjIs9xF6Oy1sweH/At5oGCj3
Ly4thKm9mnI/KaQqGYcUONBijCuORpfuzf1ERussHyKeThqhlyhDsMQCuGDcNc7sGTNPqpJqrZBJ
X/iNVoXAh5Ko49kVQlGfrW/mccGxXMOsuMyByDjr1KAU6LWDn68zguAXqZ1MJPbLyExNdaNoDwfh
M+mTXio7kLO1EeOUPfA6NADSi3i3G4Lul+Fuz7AEM/5A4NtWZ+zllHIPPQwhNFxkGBb2dsNpJ2Qm
ooAUFHYqbEaq6ef6Z7OFxf5sAFoLVIh57OiE1K5dfrLGO88+1XlfLi9gy1G8NIOrf+Pzxc5VkRbC
9cR+j6S6u4mKadPC3H1gCGi9sg2mSOp5VoTXGRk0dVEpbPGhlVMlj5ufdAXFd+7R7+MZpxpyizeP
K1ZVIYc5WsTgXSg88wcuYzN+akC02CJnt5/zk7XCqlVCOvXBWfXGXHn90isi7Ss4BQeplFn0yjCP
c6FMAgYMnd5ocJbpQe8Rl2phJCmlrdk+0yak8WL1Ey1liQDv7p33ppHef1tupz3I7mNM/8l4EMyo
d1YfTkP8DAYDocuUg3refGn0Wqu0gfdQ3MMAtVdTHNQotyvJASaIOi2Pb2w7Z7G/JCAVnoMCXxxn
w9q55JKy2Ki+YdRAAewEup5lagTMKHauOKlkNLq3semEQUiSck13uZymcFVaZkJOZJzTJrcXvnkn
PY4x3Rbj0eyZBvDEVjIaHRQvI4cgK3eBc9j7zIi8QriSLlEKEraV6gzlJrnj30cUqoKDoYGov1Dv
w2+s2Mi5lJv8zRqT1NSzsokBM8BgUi7aBZdU38Q4TBMn6LG0uAkBfy/dKfGOqkxzHmDvNm9dYpEu
dzcfFGBOYAeT1HbKZSahf73TRNYed9saen24UBnlxqaLHyeQ/nQOv96NAGEig+vdJ+puF26N5aFI
dt+RIeCBCD1sYHsqL9JHz6aeoQAlyZp2anninod9GucNdmJ0HzranQLjczoB6cWCxwFulE5P/+35
+dsqu5HK23cxvIVjXCuDbJCpv3t8W3chjp/WcbxyioF9bGcvPKv91JVSxKjgOXgz1/kDnAibNr4J
5gtJQGge56sGrPDoYPtyb2Qdy+z8wnJdh6/lGDwxyPjXs5gjkalkNYjRV0c+GnD/3WoHYSplw2Pa
P8amG1lryC0LsqkjAGfpzXGL9fZ2Jv3PLHgbydjkE700ICovJh6EjuN4kaNsdX7udVrXYt6eDCCo
UNDB8KxB0l18eXc2WbIXY5sbTvnR6vgZ8WCmbzAxJnnErO57v2TSJqdf4D703X0gbJ2osndiT8ro
DOKSwVk4c+FXQx17DMbFH70gf8VYyB+/0HyxqTz9+GXCi49WDvszhAX8Rhw40IytslCNxq4UJrYe
jV6vWyUVBcQB8+1AiZ2p1Rw80lG24VnB6+ZN0+iWwMr2g2KiG+Mq91OxsJp5RMOySDKBosiP3vZX
Q04ajM2Cik9yr9ji2KhOd3msuMXnhdNjqoxszUhDsD7G97Z55umoqXhvEQUV+uZOL1UhM+vcMRIE
PfI2da31y67lbSK6MYXPnblOXD3ra0H8+Ye1YJ0ddoTeCGRGEzf/mQEHn35gYjjF4no16wCCDZrN
R/d8ZIKk6UeFr5+7rFPEXEF+rGrw7ScuNfbTioB5ozWwZRM6MO2iM2WETMM5I6fKk/WUyuy/diVa
f35myAf8tfKMap6g4WH6hopErqXiIrp4mDrQta8c5fv4CsExIehn23jmcbPdyuwHljjOJTDS08b/
V5Aa4jg4uXhbi4Yyjf+Q5WnSRki0iOeDXHjXZLO2nX4B+C19vTGjhhTIL7TrLUkgBKpE8GNQoopV
CxTcMgIOWnWcvWmnaCIlQP3aLP/UQY3pr7570+kzAOm61k7ry8lNy4Nil4VL9m7QkVH+v5EoTeJ4
G4zfHkPTnRmsHaj18+m/nZmrjzdRhNtNULRdt/8jJtu5zS2xNB2tUKtgY4hO4ppXByUM+QuXL5o/
wzlCXWdGQWbs3HjgUSPozCbMxo/9RpKGx6Pn+4O93aLRUVzicLl1WUM78RDtu00bLOzEA8RBA6Hy
XYYbwc5Yd42FTC6IxFAZxxC7aqZcKKnFhFCSUclvJodpI5yCcphcK5Lzxly+B4OzqNXzXOYihLjB
nOXEIYGy4CtbznPKpbgmxgxKzTTYtUizlORGBNXZqe7KoUdk5ArIZIRg1g5vd9rggkDaNuhzVKnN
f5HbutQRwIgbo2rzDOY9BsHpV/DM2bcOb2CYUh+81jo7YX/PRw3lZoean8sZ6dWsTKe6UpHOh2Qm
b3KWT6QpsXyc2KKUQ4526r2/8Vus0eYrAncc9H9YtmjgZhVUOI74wzF+uW2ObR7nNOkIEuj3cxDg
4mCl/MbnjqE1VZvm9yFThHdHTEP2pXCHA48sv7UKaY7tmvMfNRLL3tWvpGcZ953rb9hi+6uKbK0R
1buQIfJhoPEbIQsjKkzViiOcAeRuUfiC1IRqPi8cMspkYvRXfQRMHke5Xy+at7lTh4YRKx9wATJl
0A33sBqEgjbNZh4tbJEeC9UasKAXFty7rOy+cejQyRFXDV18HZg2hwignnK42076Lz5j+SclYUp7
zRgtQVJiYlKxSAorLwp7kDY4F8WXY0qBMY/bj5Bz2C2+qIpj/U0xaz/kkQavKoaRVFC8i62CxS2A
FcjR1qSqEV+JRiPjtG2acz4R1fjxrZk42u5dGHJZafGNggcHLt6WadO0GolQ3TOLU4qyOwfsvPZ7
OfuPo2PiVxRllXZPW36W9lR7hTGspsL/3eHAvu0HpvxlFyeMhLyKIsSLoav6FUjf9aPnXld4P6vZ
EWL4V9yW48JtDMuADcbgySR8QLAkVMw4CBjavzopSPbrvFFzz4g9TgnqfB+iwNyC3ePxx47ZMUCS
Ss7hInuEwDExoagIGQo7J6YbWa/oWSJWeIz7+hWa3T2Q4ChVqdx2VWc8iehhAGUZazitjd7BVs20
EyXuA6PUGPlNsnGVOFlKpttvzETOZi1XyNODMug6z+HWAAxgAl1DEdQbW51Dp0/jXz6pCvDQR7MZ
200/+WY7aCzWRvCfmWnJkcNrhIgsQWeMkw3bSbMCmvEKz3NxcROPZ4j9q7o32GnapRXkXOhRNbXb
bHBrrxeyfSustAJ9jMB3ybdZB4PnUhBVQXOzqtPfXSFS+bVecAPKMe1Bqpk5wnzZAxmYVPT5vPjr
7HSuSXJbxIB6fvXg+cr9T77IpGoPQHUgJzZ9d2KJE8ZXZdZhKsVXnQpZFD6jd9e8gijmS2jvBSjD
1T4XPhbYvxcGSCnKG5UocQwcdwLl5rYQt/f7o2oxTAq0F18UT6j8PJe3Q/V/4j+toNzlpOJql8+P
thYmDKziwOUgJiHw5zbBgA2CwzK7rHPgouiQ/4KAd4MwSzojWRBFBlIy04uL8J9fUngomQiTnomL
SgsdNPAd9aWI9Dw52lVhMajxv36cRIbuN2rWjviqNqFuHzlZDlKvMIa+bTBRxFuQpWqCB2RdrAtw
9lDS6Aa+77JA2L2IGbhd8g11v9HehLzKg0gE4ARTgeCw8Yu5cxeWkZCNLAUl0rSYX+W+39rtj/Zu
NRNTrluA33lWJTy1HI+xLoKtqsVqvjgoXmtzMdrhfQOaUZ9PrbodJGsBNj1Ijx9zKbbrHmqp2Skn
XtQsGJ2o9ILdIyySa21g+L3VPBdR2YnsMmirc80lZ7+hXNEBcD3CMYc3MNeAKSTMahHBfN68EEYM
medngC37xG7ksHuJ9pb5iQD+ORzKdsQBGid/mKETYou0T15vtqzzlxyfRDFZZ1gCzWvHmHYKQyz+
FJZSdwtpzdcdl1tdon+YBuM13CHjoFe87LGujeLIL2PxdJ4LkuRV5GWllZeNiNrCylYWWQglrXT+
Gx2Bxqqr/0SCcpKlreGk8sj9EDIcledo3rr3MLRYpZzYkFiGWmRsFyV9dHMx+ySyTrJJSQXbboTB
5P0coNTBjlYyUfjGT4o7P4On6QJQxrGy4Bw5+GYSq6nw9iTsAYIXjJDflB+PPri2EtAa5QYQVwss
rEZfmbJBweLgzjgguDUxrjIW/M6XUDFVK8rKDyNov3wcxvGSfxJbc0dXQ0gs4pyK24pi5cz09TWk
AFI8tNZHYffJELfWmEgkKEETek55uByCRbq3E7B7pAsZmfC3qbbBMQbMmhj05DzeGAoowQ29m7Xw
/DH7G1/fOzLjokkDScpOs2hhys7DtCoEcpkyNhmS6wGalvioXG/rgEqElA8bL+ARh8SL2DVWyR1s
SmBbR43CO08V+slu7ch/9oLL2KKfOuTR3Ts9TqqdWTm866Rv/o6aKgqDjwMx5goVn30msY8rPRCT
6I45DL7Ka7bjxDf25h7yJ7QkH9MVWu26Gcy5Ne0uMcE6TctMvzZDPdf5pHJn2Fw9jdrxRi08mJb6
uZe2H49IcO7hKc2fcyh3UfVPvjGlgkizPbokFBm0TJwxj7nHCcwcArvqkwHkoXKhWbdm+7wXFZeD
xjTnd+NuQEqo0157lvFx5illLaOFylripVQEzto7TRH8hXW4jWl0CqY1bPhKruMhBu4wFD0CPwDc
pS28N3MtOMQClNtDsDzspXl6R9F+hSuHSTPfADD89RTCJBZoQ2JHGHWyckUPsE2nA+7NNcqo7mLx
QHd/sKpx228u5j2al3/8AzvT17ARmvaBLHwc9VWEwUaVAh6ijSo7h6oSCKWEjzxM7Ywl0Mum/wRc
oByoiCeoreEBZv+ho1Iw5iSVLbPbynYRi3bDvs4gPO4jJrHGWuy92mJTnzJuvaDScBA4iiS1NS8a
21XIe+KjiL8gqxOuBCZa4/GAoNkjOJGbrwbGcwRseVuTLAM8fER/VHeTQ7Wosn0BWaZfgSREG1FT
jbPm0McFU3jBsP7CKLeL2hJwgOYN4TeA9Ho6dkdQx+9PYUzLUexBm/oL2PaIh8KFFC7aYZIXe0vK
oxy03S6Yw1+PdZSshX940KBpKBTI9W39Cq0ZTkWjDQQrjMqjdTu04G4H06wDLV8hKC5KbTous484
Pj2mYP1tuih8u+FwZ/lWm2aG5Fm5z4zBQV985TyZubtjoGZVdjdwjAchvG8f7mHUj1ny2Rh3h7BZ
7rKq1Cr1SptaPVppldx/aX18D4ahzMUAlRaKOT6gfdxoiH4vCOqtDNAjyYeRrWWRNFs51Z5NI9XJ
bUE2GVcjoA8UrNNJgeTPS41S8mVCEP0llz7FDMSQVWdNiQd28RP25h0s1e2X+dvz/npVDccTXVQj
Wamm5lV5Hb29ZmloccVAityWmQr6fyZCj1jjtBveBSgt+9o3r/CcCqVKOQCRzEy/kknROrRNJNuN
B2q/KD148SQ1IAuGiAOrSNjiMf08eheblFTJA7yRBOlCCadq9kdMvNo5eFNbhHZWYlotYJbdPRVt
5kdpi8zPW1NU/R+srCiuDSsmCemPQHFNPfNDy25Dvy8sOIQh+Mmat/+fVVWYjHyRQP2TKOcDLgEL
urY86BUTQ7LI/5nNcorzsPIsLdx22sg3KW96nPvXka1Ys55qCnnKvJQBUFzT9GBnD8Wey9La4fy4
Mq0Ic4N18+ypgr8vgN5zz8kGHmNhEVAwTkr1+FRvSur6fyzd/xb3EzbSITGUWm5yYEo/42LLLS+J
TaJNEHMxZlaVHLfHjxLmHKQh5Po/lWJWc/y4LwbEQNIMVRebpqeA0DuT+fo7uhhyfA6zYmKdrRYR
KvUV9GGEZ/JoGDXTNnumPS/Z6PrpwkL7Yq8Kiz2T1jGrf0oqk9ZkV2SpTbg6wcyd0J/dUELU8VHc
iTaSu70VwEMzSfxXKhXHX7c+pUV90hnxJwOXCPWO1Ihm4LGhxzW79FkXcXV+joJKSwgJZ/o0iXVJ
flbD7xNmcsEJ9EBpxGEy5S+M7ZppYphJy1BTKeIQfRidL6aQoZqGOOd5siaWsxeDC2r70grMNg5F
XR+Vqsf/LsINo9LITq0cTx1y1goxbg7eD8OrTflrjzseqRGc61XAAmJCpP77hFhLbvoubF+2u1We
Qbcfsd3+P5w1wXiFD8+ROSWyEMXyc18SFCEJ5tT6NY0UEfdyYcXO4gmI/6noEoKiUrQEW3ZUC0hE
+jY6EELbjpks3WcDrsBEamc9zKsQT0cE1jQZw1UByOBdL9XZTMeXO0+GEQR4/rUlJt4AS8TxXH/0
3GdAfDKPAgU+Eek2ZWyZ8BApBxYQ40bIq8TJICXyWDddS2xC/Dz6Kt80Vu9vQd+0ofb1NtgVfIUb
J7Ns1xze/qMNBoJ587z2k5NnRLY7GodG3Z4edvMyts5v6+Lm6DapljMLZDBl/trU3M0Rfgn0GqYA
xkfORiZqAhkShsvPSonR0r6YDegIdMSwg/FCKOtzFi5xHwPpHpQ4dd0R7dXsRUuKaoEkSBpu5C4v
LI2LoZgDw/Z+zUtRTAkeDCZxZoa/0BN6XyeA/CXsZc5Kis/IlubSOMBSLstXz0qoTuZpROAv37D2
KUd/q74t9J3yiKKqg5llsinvRQHUzv6Wknzt0N11NWT0qhdiJsqhArPO6vjAIzEWa6ObVx7jLls3
hNQPaFwbulxdX1goV3npJ5HvP4kFhzI4LrwVEAV/O75Miu8aAYAhifCYb69p2tEvjbOIIMt+vy2I
6HGjHV7RUIbZoxcHJ10lK6QubbPbk5HZrsf7AgxxTa2CTujS38Tcs1gS8YLyY/awVKjZ6zgsGdNQ
w9JZ710FXCKgYo6EIunVa1Q/Wa1BHyVcxbsARlNLmhC3Rk31tIZG057eXQBEbpBKUNalSg/9ZVrK
EsYcQRHoFIZXRxbvv6RgmfeedBj41lOucwGhIowlqp5D2PmGvyDRD9Pf57ya0y89sZVTlyS7kGnY
KlL6EXbSxUAIQH9C4ETtHmn64Si6WGjaug6kvGBzONjauHtlcRWBoaOm7RAJFpv685/xGiTSpiFN
XYaPqgXiXw7H35pAUTtbMHdro5a9dblqnSgZDDgwozQDnOP5xpN0VssxJygyC9oNSnfQLpHNYHdZ
lExVLAnEPgu+xdMWxALeb+w8MhVuFjeT4qvyDCWF13ZpmdET7WmI4MVYpGC7dsYwG73RFSMtdS6c
f/Y7fQina/JIOOES9PaHYVKP/bqjFWvxcaiA1LE/QYsshMLPSiP3fgeCXV7iuKQwxb8KEcmwARwA
Go1+X8S9avKokG6K6dCfcFhQ581FIpLiyBFBa47Vbw+esKin+96OxFh0870rPwMaDC9SRXlGQUXy
fmekqv0VHbaPSnfyFezvoQs55rno/n5i26OQxtlCzr953R4Efw9mpBpHYxemdNzsbKPaFjqlp+X6
WKcPaUryy8/+WSDvVyrCI0gxR5JZ7UttRfNWOgktJ8c/+XY73TOWCjhWyNbJZInpM9UP+iKMjG/J
zwGDvRmU3Zffp5CVlRPnAwY44aElC+IV7D+YGPXLyTrEnkkbUxc9TQsab/sAzIcDVN0k1ZaxCmre
cR1aXDm3UTJxeQTWFu/7MqsExvWt6VlVAurIjky6MXJJ+KNDjxyO0ksvHD6qDEdn7tEnKYNXWVqQ
JLfppHIknHvSuSoeAuJHvv0ED80wy5ED/yuWF73Vyf9hIYPcnBgnShDOobEQvV0jNqOmKrSjjGXv
cULEBz8jNjhPv5pAF5PyBaMKgWGL3SrtVq//QfA4NJ9yglPFmMVFPG7mbSFj6HMfzICNHm5AgX4x
ATOT80tDrJoMwZ62NIFQHdkptXZNAGC//iHph2MugdiI+Uv9+h6SVJVWBhXugHWxi7omddPlVuhf
eL839gGh4641bk3+BtQsgNn7CpBSUVL2JTOac4cwFyh8wA1D+tzPkZssbC1u+yVoq52uSvBe9BwR
MCBtS5Tv7YpJ5Q3GyOEo2QQ3XQvLvLuyyqDLfAlAJfOMQcItVrFLeJleECCRKDuDVfRQNqOCVf29
hG6ANIYgMmVw1LFKz6a5VmJoiIgc3Z8ApvJAtb6Dz1GNe6GRC9iHRI1jbAZC/7BMEmED33cloAPG
HcGcpIbuvGpJQtUlMx6HQaPBdMNaF3EQcdFj4iF4rdbmNYrVOPiaQrhP1AvzncqyuQoED5jCFkAI
qSZU96sTG4WtQ3kIC5403utLJ9BQdW3Lnf6ZlMvqfEnjvlVaUlNE8fTFMdyqAGq6zJkViUln9MNj
Y1c4Auo5X1KFBa8konubnB7Kd7/0iOH4H5gos6hsjZCQmyGOW1xneD5E0R7stUTsXv9Ta7qkqItu
wI3jfl5h2Otf8EdUOvE630gKS8ki+Y93i9/6cKGaGhr0g+1VqrsB5K1LsbpzvJnt64nEn8C/ENGw
w3KWSuZwTZiWCLoSGHXsg0EN/TbtRwN2IAENFFPo97wyB0GdyGjfV8DXKICGAmANggBjCT/O8Cmo
IXp6raVTvRJD6bqqQs61Nu4akw2/DZ1ohw3GGKgUk/cuvKWSmoArOAqyIxhTiJmXOh3bw9p/7B9n
4fHHTI9lk/1OR2MT0ur9iL/iUifTqcnbJgythx8VdDbxHUVnnZlATAaKKQcz2zupDh8z7WlToQAB
8YAMPClRVwlNGiBxw3qmwGW5GOmXhH1VvNNOn/4SfZPXn3Fa4N+rvhdG+B7btr0YBx2So5qOSs+I
4Vk9pu7wqBfnIaS/hz8BaM2WJejHSxT3QmPcuHJQLiuOXYHqUAGwMSyJs5U7SZP6unvJhdRdeg5q
SmPtV+WqrH5tFPk7wcq67KOehG8adqRJUaJ7BDjOWg1PG7uIaXqwag/0GRSZDn9VIbCfrL2l1K5W
zH/qrsgyzHzZNdSVP2S+x09hjn4Vm5zHjACU4ptgWXLoMNx5nw6gi6Ym4w+9ZPnoDi17sp+c/947
Zm98XND80EF4W96dNGKbmqeMbAnkksBAPjiwx9smInEJFwhvcwfgp/VONDx3Vr4CYqQmb87YBdlQ
tULdvYuMaSWA9QspXxoHuplJnn1thLwxGhNxVbpPZcNJWd9rvfwKtxACieP2SCcdlof7nsPvOJdi
s6OSW90p2JRIHdS6knFTwbw1Kid8b9aQjOK7rRGWucQBaiUneLMUDZ3k2Gdt5h4AQIFq0k/eA5II
aqwDjFT5kZFLy60ZQ1Cz++MDLhMwlTG//XgSYnTFEOqgaD8FF5QdvOyomju+QxdeBjfN0pJONMYn
s+zz/ueQUskg733PqnXktncESNBfT/3/Ut0cQfsUnXxebkX2GqB+cKXUUo3UiwiiYJuRYJAEwLhJ
LGUUG96pR8fpHQph27NkDZ3DWK/4rmCe3ALppkxjUHWcFd4211TVjrezTa2E8K9zynS7+izVm6qG
uD/o2pzlNIymrGQ3WxLgl1mcsnvfp4BXGUvDGiHyf3XwKdqveZjibGQBqwiMPnLXpg9bHU8kXopo
rUpzl12Ja9kD+y3kGUD5B2S8r5w2ccpcWhUoDrZfcH8wRYV+NKRaX7tZ2aX570SUbebrI4MA/O97
aih2LJkjH0rpRUvlCIlTZvoNbRiDkth5c6JKIJ+enWHFY1qJuKi6c/1VFx4gM0mHmZJ/UYnJn+q2
OAOkS4XePLdbDJjcNMGTJMQwUtAk54SmX4cldKi1KBjWl01cIGblRy8K3mxGEC0O7XZjVtU/gsFl
10y2lsG+IBSn7jOZ2ecwxFLqObwued3H1xctVCxR7F3LaUiqqYvXsl4AHOEB/himqfT4mH/P4pz3
wnzI2UzuhTH3XjOyOmAxqhnnCm/el+NoAkoPcGl1K/CK9spkmzMn4X4TfzwveA3n71LkMeNoDMA3
oyt01UzbtgPJ4WQ6Iv3se/ZFvsADddOM6bTVCDImY0gJKvniWLlPrrRTV1HyAwfELbNbCqFCenXk
w6IviQg4tTxIkwlrE+6alPLeyn1diqBvbHObkSPwcOzLCrzJR+zwju9dFMwafPkEWeqwLYzCF9n3
ChaB4eMEF9CqXjOzlIJjAKgQAmRbPyOvGfXeJ60ix4ufbp9+hhL5LJT8KxYt/6Y3oZgTGd1wHeJi
TjeFo7yFzJeg9GcuClO5uC++spSE19Ta+hs4/4hvlO7RKAGpGb7sLd4hAN5YydGX2AvCMULujbKR
CbpeyVnq7m/VXKwonay1c1Yv9q+sylieVJxolv7fC1zn6wnmcuTlYjgY/WFQVivSXzjJpewmdUHr
jvjGErdUPkGAp2k9lMogUyTGv/fPeOGSeyA9Maux5m61WlGpIlxoBiyh2250HXv7MN3gHIm0Cjjy
QK8gBofCDtdoPr7+FXfnN8DJORwgU0RiFoZxNS+IubOyNa2QoTTEIFPKbhAvXcPAlsDYOca0jFLz
fpoDfnXOKfvXZHNmRhSyqi7ImmXD8u6tQDr/vCedxGfzQwPZpMZPgBKYAdj2zuLqcAA/k4Mtm4Uq
smyLSh8dQqnRth3bQD/VhJA2LSJfjdwXn82wc/qyYYIPoAf9dpIZ/OnBvEyxa8W2KG6E9aUjw+0l
iIA7vhhx2/piUe3JBsfQFrOLoO43sTaZEp1wgPH1yI4kvi5rMXGOXsHVFSr4OdaTI9jpwUaAECz4
ZU2TfvMgeBVmW2E7uCA8uuzhgA1kZfi+RVn+icrWPwJfyp2+b4AuMlH3O0UNF7gDq65efchIfCM+
aBy1m4cB/08+jc5MzoybvtcmYDN2r6oDSlBbXZLF8VhE5bTnqZFiS5UnzrCEkKO3LcQkZpTuVRFR
9TkEmicHRy5FTVGnUDGq/4DwB3ytQTqmJih+ymvl13vwIJVa8N/g27kO0Yhp2w2JRZU8bHwM1kEI
5VdLsHXKCmD7AGIBCImkcCK/vuWS4csF0weyuuJXRJQkLdzD7BnaXjtVUySD9EKZdMD2e7PAdydH
yuFA49j9lcligkdTpJ11ztqQJhByk3pL8vw5tt7hErK9Uq3c7cQhtzV6nKS1cZ9SovoCwGXJ6CZm
GjDpwxsLwK7H0k3wUulv/uZYQ+92FoegJrmNlVO2Co2SdUYjciu0oJyezd8+RXIa/cp1ZgdImQ+O
+teysVUqftOmdgD+NBTWUo3uuS6LG37QmTe5Iww6ETJTo0viE0MHB78mO3TtXSn2e/tpZpBMikNO
bsDiU+bbjqXHQfK769eq4suMTCSxKnmMiye6mbgIGZ9yUGSffBtewz9AW9a/qY12vLRUejG7CwwB
mjtE6Yg3Lqp/E4RQpUpYjIVDa9KiynlmyzmrlK0FXXKXDtk2FITYzaHsS9Q9RPVtaepYhM9eSjrm
ris8yo0AahYkzch6DDwzOcALG6iHJcxKIyJ9gxdMj37Xa7dLvdDaUPxc6rmEhe35WcH5OTp9Y/l9
91RMCs6QdiAWl+mK6oUToYCtBsUZPxpDx6Ww6k+CJUNBwF6QduNAJPwf4Wqh1ALP7K/2o3Mvj5WL
VHrfiFbBRn4Sj1r65iKNSKmyYjXpAEiKA2dnCSbbCDofqBGhd7lgvMg1heKv7FT5wqk/EMs1vNpS
Azb3vlIfVE8RBL3TXo9hfyGZaXDZo/8MnAy6xVBGcdu8hZLcexBhm5xHbRlxAwMMpWTsz5X2/Woh
pHzyWymLG6MFmV74muwF4rTay2S/lKuzol99viwYAsmc5uUuKL3UW1AdHz5YRpj4A94ZfNjVmK51
iv9OQJPR2k7A1x4VekgVYhRLWh84dUzsfVZEyiYS+FZlYM+3UamSYA0BU3WR+37qg07MQBkjkl0z
5UNF/mF4EmGOOBZN2ne5TgE0fy0Xdx6IMH95cW8yrgAAmcrOOBD0jkl1T5JACtmGsB0YBDSgEU/a
71ayp63HIz52WnCTw8ToFMLmtpIVVeXmjFlQBeyjti6YUih30KQe5OzDeJ65FT0qsQLX8ro3lTHu
rNwhw2ce4Z0c6sPTrVHf5fxGi0sr7oNer4zVjTloACQP9mp7rhOxyW4q98gV6gb3D4coMgiHmmYy
YyU0mTec0myI6VIzRl+l/7jm4OGdhxq8qWFoFFwx/6JyuvYeWmXokXEyNhOPP71agGxt06ucuLZ3
qm6WvQovLxNKilLJ8z+pHIlhXgnWwxbzCidou7LSNWiQzJXuQoszeBDglKRxpCdzxyqvywK3/WIT
53bAy48V8LMjtXEcy3Nny0dokzrO6L6fR3J94lXtfnsmDHBcspTyGhOgnDjV28/ezwxBGcwBPC15
TqxSAuxwb2ILEcB/QMNuB98KO+lN2YqrMVI5Tv8/IGLb31I3AZ43euhRA3hIrp7CEH2+lSH3J1/f
w6ekeYQ/nDZ2yzl/eaG5cbkTun+F1W4+lwFO4eHjZxj6896x5ILn2/SpfdJjscDLMp/0/8qmShyZ
t7wyxF9bGouQzpqijmbwVRJfz+8jImSSgCDJBZN3RFyGYJv8inEhj1BJGjJbZoTkJ4mbJGYiykeT
fXxrRGP0eCpWXTWPE1t0Ns8vG4RoIrTNiA8wmfobZC7q2k3+YI+T+ZVfQTHFQBfFsdaxkjnGorJO
vBfw1FmJ3+qpicjB0bk/0JzA24uZ0+TK2SE8ox4QQGeoQho4rwxUjnoTPwWEcnTWj2wKkBmS1bX+
LI9vGBawbXfhvd/7yUw4zWB3/W5MsfIWb8542t+SGaDLtQ2DbQP+SjseWmwtHQ2CrplW3RQ9Q3HN
fHR44T3e4Op1vvN5ZryuB4mvrO+wMHJox3PyVf6cRsI01+DxXOFBm40imcVEORXR27L2PIqUafZL
QZj2mToPBeIU6WbkkR3IVvR+6YV38TNvHjnVmfU67RdSvQkQkmW6cz6SVNtQTemMDazgnHBwqsbe
HQmQMBzldyvL5SG/wggjs5fKhGdqDgUq/KXLl/idhTF2JTxJmc2TJ9Sf1ERamigmSU8ALV2p2Zs1
QM7JUjbyaCe3UGJtKO1LznXcnfH01RT8N33uD1DOI8M3gE07H9zr+hNy/n6KydHwMDwwVmoASNLQ
VgZZaf/IuHWNnY6jbuYvKEAJNFi35TOdX2+oYZyeyacYbG5NYqOkEGx22Okw1DpxdCj993Y5WoQJ
cmHu4Rgr0yEhF3pDu+bMmWWeXS37bDt6EEPvPom9e/arPL7VDkSRI1Y5Myr5uXfTHMoqge3R9W0m
TZrzCvmQctuXr29yDn8Cf0GKqtyGbTr4F3NleKAV160mzz2YBaKWpAUcqmPyEVrJKk1IkBAvqViM
mWoFWhw5M5UliWPeBhD1BhfCGLbXa9gotx8Nrn4tzRIde6tULZguJxKmtEm2WPcdgGY45fVAtYDN
VasM104H6iHIQRkC6J3XLrWbURh4LQxXWW9rbR4v1oDKVRxMfLLIHF26bDdLW3bb084euiP5E3HK
PNLQThrgBz+6+CeDSijmtwJYTGCSl3f+hLq2LCcG4T0VtKXGsuBWInh/PZOdYbNsJNHEO2nfOCdz
f2I0umwS2/X17cf3rranJQ186coUjx6LczNz+LQcLdIPS/6fun9xbvWwbjSSiVAMNcoqn8CzR5SW
0qMsWsYs0SX5EbApTB6D1gWTCO0atf2DB58RpH17J4YwaDNScN1fol8CgJDTKDtzIZkqFbHSeUB1
ZxWVckMRuMsWqY84WRZz2DLOlxt0dU+xYzJNaygRzD+mF6h8TVjejDt/pQXBhGDU8jhyQ9GU9aKK
8OUkVZHsA10trXDSGRO+gmgrkBmNdVdpQ2S9BA3hF929F/4zaLoDSqQYE0/v2u3Qll90iwh3F7EV
IUAwtO8TkhwRy2CPs3klRawa4B5xL1yYfKohimO8k9sL7rFqeAcqLxiVIxl2BsxPuh+Ywt1KzqQ1
oWPShlj11tIxqpZTMWgE490k7l/ERFMJBbLXxc3rbjMGd77sNc3L7QTspVbCG0CapUQkeEyXCdTd
8cNCCZl+LSwvoNQnhGhL1kmzJ8xf48aM8nbnkRyfjy6SDMLKfyp96f8Y4CHNyL47i2lbf2LfIE07
QSqCoyQIBQhXncEq1D4f781vcien2J2YknXjiAyZqTSQDtlS0rqQQJPyYwYXi5/HR4LcOKfSBWlX
nRCOZWqsu1Gjxt2wUhdGSxv5ghBmiSxs8qBQ/Ul7v3RhXxowMSkQ9NPKtCvTrOvhQgaIZuEqLo+q
OnN7SxtCCCKj3zPRDbzhRqSRspd/Foe30Omf1Oi3hc85L0YlYOGdHX8/AjU0BNIfGkfqeM8inj1q
KtcGa01ZJ3iHe4Vuya/mfiQ0HE5jyk4ewheRodOVY5YrD6HsxTw6fUfUjeQlsdftI3m6adFugPUl
DuGyV22pYmm6/HbsG3ksFQr0/Jb8B545Ei+5oOtEDn864t/NUJfXKkKNF+Q705wUGoXulQYE17T5
zuGKlhfO5Ta0GGv+oubyx/VbegUz0+ZLiP3vVVf+HiD3KPBS6J3IFHR80OEGLLwL9BUDQ6QnySzo
ogZk5kuV50zN/By/ATRCeWjZFmY2NXUKtqN2boWMjCjaasc8tZ12YyYWgPa1vsk9fLRIGzBDWU/6
8SP/ynWJVHfHxPUJynEumE3O+kKIn7N0LSlsUXcnoJBG78oqaXPCqtGBKD9nd+E2/uFeYLCnlPSm
sQZeUFW9N1llyJN2hv63FnfVZNedX39PByNzz3ngEMTG0DtICfkdw65lfYSzjPRxszmFS4uT6kuY
wGn4gaOhpqK6rmk+zWBAFItPFPaNMhN2Nn4IyzxpzpjH8OVxp7YPKiPEMTt1k06oTvroQYJ7W8o7
nZ9MMS65Nnuf8Zhgx31fe+Gqgm9rVv6ms0r1g3hg/pABhje1fBuDNbXVT7ZoEX1/e+RMTQmoQD8r
BY3whN5bCbroXQczKAAjo4pshpYMiqzj6TJHbGH3nNODib4iqi1XJT5l9CRkrd3VUexpt9TDEzZo
f8Y2jS83Qbl/CHMs0VJs8ZSLFstWxwI9nXkIjjS75pzSXp+Xkc3xM3HTRk9CkT0mAX1//ZmkaZWf
kWn0kGYKuYtuaXzePIs4oD2nZVNbZNgSljysf5TKGk7osIUnfMV2vxE3kuGkfZ/wDL62ahH2/MKL
eoMsu0Ov+Spwx1/v1+sGAJ12MnxWE96KFDuAcET2T5w7hA4s+wlg6cwWOiScTgLkMGj26yfQX1t6
YbNMe8FEBeFLjsD5wrGTkrUT6B+UV/ityBZAmJC+0+HtTmRi6Hg+6aG6D4jw2jfO+xcTxLW6qyCh
Um+pbQvi4y7rjnBY1Qlvl31hFHMIDqoGNK4uOxOOYGTU960uR+gwhXSh01JJqo4icFxtYhDSWUXK
ZaB6vtkLufwtDq5sc923xlZhISQBhlKVsPiPRGJiK4nEj/G8Ykbbg6WHsHfp6l6EKzWe+7f+p9E6
S4kemf1d9GYZ9kXodgQfgp0OBxN3mRKBXKeMCvAcURB+wGpqOZ0DJCV7h2ngpllhYYaHDW9r9UVy
92o9bx94ChuU+/hMUPBe4+7pGlSMJhPBDkZsIh7kOlK6DiHTrojtl6b4cZzGThznyjBIxQI3qaLi
yDFUh7nBhhDBB1KdYcj5q9JQb4z0CjFme0H7CvdsNZmMvIsfNmohKYKZKaCYeuCXbDx1ZxOjlEQb
nR9bw9IgtFqZZWrZfscutGFeQ64iuty+v7tuaEGKsjh+NbsGTSzjyaAE8jXTfGZgV7ekaJzWrAQY
IxSPCNMDSVTHaFgeaC9BFnpwxbba1Mb3UTiZxf9leEPztA/JfK8IZ1ePeUapPFYe4GaJKjEAmhtm
OFfvtUu7W6GAGBNQb9J2xoFY5FcvjtKgjwT/fxdY2+zFDpvV8FJ33ZOIxtup5BlGlMH83xWAdNcj
7jvJMJw6wKggdKMaLUtfzGErBvGdSHhuWv1ieBKUJ+4IPg9uikgcWMqcvN8X0JbHpopApWRafXgG
KDP1T8W6Oxi0reimVh4aqsHQ3tjhyk69QgQoKt0P7GVPeIGwDio/k+ggt3vwxCVu1xKMO+Yu/zn/
wv7Ohd386f4Oy50VOQwmcJIHg93cyA7zyCuetAJlklC1DE5uGzsI06E1Fpop9IcJzJmKPPtlO+fC
snVFMOMNlQc3QsBb0VRlgcYDitTn1bkxg/6KPQSl2nUwgHuyE3A2ot63lY6r0MLRDkx2nHZKrAaJ
FR8SVc4+89GmIRPJ0nElhcVpuQt9tbiLC8u6gihJl/mn6YdD7fOc0KYE7Mld4tMmZYSFnFnEYX6F
/gMiUeosaEIiSbCIPZb3qKzsP4v/qEtvGSTtvaBoIIRgGn5LqAFyW+jWCKB3dSLOqk7qy77hwNlu
V5OluV9cIf7NI4nfzLuZvbvD3T1POseLQmFp1ZTmpYaMV2wzuWP6QDhtR6l6E6f/jYJvvL/BTVMM
y13xWPHJxDYf30pX+wVyt9hs2CaFuV1AlRgulSphqw2d6NcJ3jcE/M/93ZaFcxZD5cAs27C3/auB
eeOrNrgBN9Zl0ni99MhCjuUq1ZgCN2oGeGq60LiakzaztEk7k4TYVL4mj50Aoa0xzKbD4nvAK2V/
4JTvJb5PFhQjg/ffhPMlnPgVRitRO1yJQQ31fGyP2nlLW2vNkqDTvZ0kI7BfShF+gI6VaCZj61iD
86v3iFq5EOgGjYaqXMUB97av88DRpposg/d4pJ1c/yxE/JV6PoXJwmsWU6npd3OZLO1IxtDsVPGl
DprQ4k0rhdDWYPz70dojiVcUC8Ewe9jRWYPc6H9t5RzbzKFd2sE3rf+PKp/IACN/fxsWicEuJ5d0
nolIi4XY7qT3oTeOqNNLRoltvCzuTts5k0Bwsy40CTiArfNQ4V4vcV9Ov35ZTaHUbJYCVQOaLrMI
cn+4CX+fJCAibPnbLsfNa0jsxJoXnGGpRh8JmcP+u3w9OiouonW2XhOg/HSrZrCE4dTkurrJAfhh
o+s6A7gacMaf21mEelVdhzkcNroAKrq3+stemdK5Oqv5HU+2T0G4DTTW6bknqcXScYstAdoYf2iF
7uk0Hcp4FoXQGwPwqmbjT7gJNxSPTPrqqaDgF/7YZWFeeupfr4gxACYwYRAKM3M+ttH8+IwtMSes
WmDb9XubgzZ837a4r4bpgFX12Chj6wEcP0fUQlxbTWKfceemneY7eWlei7+8IHuYTXTzozdlG/j1
01hWzgVDC9QXxzOFQY6D7N4Kj/eJOQDKVBEYGcX+lz3yqyKX1IDGLx9hFMqmxn5gksXWsLOquQzA
2NQ5yn0fibF9AfpAZ27Xl3gD4AG5/6Mr1G3p2E6M4+QMClT3C/Wsx9DkUgvHMvuu9SEAybg0sAZd
/8G1R0Y6b50xsFuth8oxAMdvSRR1AA6ukKxqKFZZyWB26/nWMSAzCFrjhcSbHxAi2fMDf/MEyrpo
8BDLPn7EZ9chMDHIBQE9duKb0i5o4+mkIQ4qM9xmj7zAjLLs+nVlVkbn+RLc+N9lXCBXyKtH4p1Z
I1K4jUaofFJYGJ8cgsWuUJp8LB75FoaAFiFny5h0F6FaS2dEtMsL5UQBzGI/Qo+kWKWlj5ZZwUPp
KriqsH4X6qUDWOoqx+i5ky+gvFbQa9MuLlk8osCAF7WbS//iqzqEz1bQNeGptWL7reE54+l9fkm3
lKXWPSihMOkZdKgawZgpG7jnu+EsAkOXO243p6NxxYLA8fdaKkwGta7/gDeDkhRUNKruWh6wAiOC
nfZlc68DjSS86Fffix0RcN5kUK/NYfHgJCUmk3OdUf2npnVQPvDlOhl+uDSdi3t2tBEQRqLnFysR
hZk4WNABSzfKTqpi7FSIlRkrHfeM90yKOUvQXRWFBvtCzrDFBgvoCH/i9ajGJm0FQIQ6mrUhUcRT
f0A6IknP+q9O25WpLR3sGJbQMFx1aS/Z0SBOyb149RttQogu6LBIHbZG1gQeijBb6bfSUW7Z3Bkr
yXHfzwNn1Y/jf43xb676707J1xMeDsRdmS98kWYGmHUmQLYUbulugyfzVz4XKYjmd8NmJq8hfkUr
o1IkVJjvN08pylVyrzVDeoTjsZdEKB136Ce/lqvBC0Ri6JkJNvJ0N8IhCyWoi+wGdQbZkxGCEN1M
k6dUTg4UqHnguDa9roO4p7zCRayZZSGSWWo3f985sB9gI03v8TPORHkE8vSJULfs7FsgJIrYGntH
Fdq/v1cWkXjSu6TV9svno7ULWXDoFZ1XO1JeoJAmCtfPLtus4057k11+tMEF29xrIs6wNOdoOPq5
a5mZ5GRGf+bRBMPudDogUphc6oMmbdYptQ5A/NfMCN8AEqOp85LhX1F6AmPQY2h1YmbEVdCxk2X0
P8UseR/f7B3ZMFE/TAfbCjQPV3zQarS+YpM7L+lxbjn0UvfXmwcBP2bjNp7oKHwQdkw7W3CgvTue
4SRtfmhfUel6V2zQ7GU2Lv4qCpY4kMkrLypXgYvEooggv1Vn+fzJPAr0OE+MHTxGV9FMJkvcpz6J
4W6x89wBJQqp7EeJT5DqyPAGhWfiNKgfG/HjQhZTqKcZaB9zjyLD3oJgo0tuxxGU9P2LAErv/plO
8X2kgZlyVzoFyishIsp9LTgPVEhUGooi6ca9rXnNBz5LAr9pWksmNskXfUEoJ8xgZFU8ZaK9KFcw
LjBHofgF5R5pti+B3FCxJFixiP2Nfm6wTHM+ALUDxCy9504CTAS0rvn2jjvN9eixTZr1xBCieRaT
SxM0L6Mllo8oHbq2VKHDQ4khi1P7nBPZasG1J6dUOWdyAi2rWTp+DRTjEsC2Fx3O769ugpv7R9ZE
QmPrYaqJ6s1JFH4pNBgPvhExXxA6U8cHZXC1A4dmRCTmvAUq97c7oDDxIF1/gArQliTaJzSAzmqO
jnOAaXaQKHFcS8pp3OT550gv7foIfTnPrc6eHQGh9j8qvoPlwGKRYgzw3mhmMDMK2f9+nBhgifUe
Vebn5HsHyCRK3weTSSrkZgLTM/Hc+FhSGTcm1uCaZGMNtFxoPW4JAC2syaD3Hnqx74KZdNpF4J/r
as6/ANA7QxZyATyw1bEaEp6TQByZdjIxcAjDHRFTu7ISdFfcOYEB8U34vgYTn6Zs6E82K8GaSi+V
uZni6BSL95V4iXICwefS3uIigNk3CMY7Ygx8WrwhXuwiYVzYrpnhbNNcf9/OTMA1ouc9/vSWE6Gn
SnEBvt1mzpABBib2P2UOfT6GmIUwa938MYNGxbf3T0TS8NYo674ezvX6hrIRaEExezX3cQLttqiT
whSSKh5RtxG2SXefo0bRKZLEugX8ehMolU39f2NcEhwAM15t66/0PwHqB0eOgpSa+gQCOWusMW/t
mOtSyXJruhYAEATJ237AR82595O1Y+SNCEDJbUOi273QWzaQU/hDmUS0M2vzbs2tT9x6UxaCONkn
Z1ajlG0fw0YFbkmQhtcuZUVk0ebsXRSNJEsY7IYkPosLcQKwmw18tB4qwL31Pm5QA+EenhsImfvn
1uSjjqPuJwkipCmNUZE6LWz4zPgNfX0mezShL4bnM8N6FkO0B1Vf91m6RmDhql6q9jO4CnW5umif
SVFtuBr/6Z0oCr6EILMKzrGcitbZ8wi251JhEfip4/C13AnlmRGs023nIdciw0/NRYFyIaoe8Pol
Zg37PqfniSV9DJqbQ2w6TkTOO3MI+GTtY7bH5i6ULF+Re4o3JGfx49s5eNhuxPS2/Kh3pVJJnhDN
wAbQyl7UMhHxrX5MdHwXNGKR/0/o3oxTqVA4zZ/oi1ZEGdTWszMXr353CSJmFesoklXDVchIxGBk
Tic1uDTkH830w7ODvECGWboJEVJlegJW1sdEhJ9T52el0UXLZRg/HTO13XDebaalRpwJnuqlQ/UT
4IbPUsvdW7XDCHVDlJloFvGB/ZyA2ueC99HtkfM76HHTvzoAH+o4ShHo/EutX3qt/cs1Wqa23jXB
R7fMsoTUrr1SgI8h6mpCiq7jM8iNQZ+AzuMMLwKGyUQ51vAizc9Inrc4idY1hwyilCCi/OqSNCNx
H1Npja3StGfhHaraBs8f9I7huqsGfpmcPKdemDTLFRTYDhYINOAOipb8yd/5PBMRT73DCbA1Mm6C
w/7Y/fHgsN2BfPqGDjqLeAwA9o1c4/ro4hwdbxV3kV0yWPhkC82GsjpSaKNXfhPV0G5v0UxFITiy
ieJZAUnmQCvXqB6jlTZmwWtaEf73gWHLyMw4nEGm3FvBXUGPmkiD8uZtpPSWn6Xok+k3c7XiSso1
qtD2RaMwATe56AmC9xigttY+9zlLdhU2C1oY6XebA/vhDPpBm/ov+VqXzmueHporaKts7gSD3qae
TGr/XGcLVQaXy55rzujEEcQgfziETzaatB6+OzDBL/aHrXVE/ZYXksMnUq1L6A8r+Px4M7ZlP9kx
ctnk1Il+tlcccOj1/RqMO9acRUMGnP0w9ZAXpQT8uaZxRL+TESJPrhGN1ztRAoi+fFR1C+mnSY5Y
9HVrSID7KpiXoBGN2rDNSMqabOgoE22aU4PiNeFlMAS0rcVuam3vdMAsXqOFsDJm0Cj5Aa0QfUZJ
k+/QtdrP0I7XEX7TSKtLF0y2FpzdDV9iIgLMpXTC6bLAaSn5ytIW1vvBiYUqHJOVd9AU/Rd/lqZl
L+q1flSJr18NvF1kE1r3utU6WyG63Aw4ifDntvP9FHMlH4Z3+chmpxayvXFRK8PUIhWqV6Bgdesr
N0xNOlelROITg5FlinYbGx9yWu7YOG4GfrcmEqMn6mLja+O2EFQFHXMWtRx22sPqREFXkHhuDTUx
/1DNTWIuqTK4i1Aog6bgTjxEE5UM3IuPSEXOxmGN+kr4r7FHK7+Odhs7jQlEV3OG8H5CHXDHqvFr
h08IhBEJYFxJPfD4GtxPnHGD9T3KwcF1EjuWkuAl96S24Id0x6sYRnWpn0t0udzES1kTz4PAVy11
TgiDSHQ9mcH7GSyyoqAAUKFyBFK5U8JjXqYR8rRUTWAKI7OtTyTAIlLJEwKcil9k8y5Na6mM35wY
s0l4p3Oi9EqXqxj4jQg4NycKAW6eoLZ6qCYxRar/r4SzvwYuoZli6X13DnJMGA3F8VyoQ+XBZfPa
4pYCMdrs9RLFsUtSiCzpJ+V7hiNM/0eZSUrOMWuOucIHBFQsXVFEbl4wBoAayBfuQWCoDBdIlYtu
v/SodM9J6d0UaG/BrVOs+2EQv0MY/1jcuFIFfn7JPOm/uO5wRsxpmvAaw69F41Bn7cmPmDM1MDTj
PbutyKDJ1SXIHF6ZAwJRki5ODHhVaL7zH8T0BIUXmMu4pNhfXMmAzNo0Gi1xxdXtZ4COmiDZ0vGV
ED1bHOOQrgkhkYihCvZNwgxGsvGeV2uOCuHSGOuP01f2L3O3BPx/5WDMNMmuIlUG3ihnVXyJMShn
S4Ndh9anyh35fhCiJ1xFY3cOnCs5BgBUWj1hSWfSqtzimHG3/M7wfOO3Ui/y9USqwq+wUeEpnda9
JQDFF2E0rIlVcSV/vpLeqwJfEpIZ4wYLnJcvqlApb+Pp6ezh9+XYeHHUuRh5w7OBzu0z0K+zY+Vu
I4InUcL/cBDaLbyF2fKIO6GfprOibncUy1GdbsJyyLeC7nPgpYCf1rP3VzWZEwrlmXBplLPR0w2v
FJygaK7i+oWYauG4oMxDjOPdULpvQ+MTp4ayGZ7S/I4z24YoK0ERSWEe43/hUQPiM1WIQJ3IYJKF
Bu/cQWW7HTZDGEEkSqiYnSyZZhkocQRgo6IvppTdJQM1MVvSYvRqUeAFWZTVSBxT7iieE+1QhJdV
3pn7FktcCKpSsLy8nv3pXfseGRk3dRD5IC4N98xHQXqmnxzGqSsquDWwv7nmqskXoTVaVZ564XxT
NjwHHmxBYeLsmodi7HFUsPFkMNMXAWMOFfCaAnkHBzDtvAvdWIx186at2Y5Udwrlu28JWKslFSzL
dffjQsdtqct8SImflWMuNw+dc1R90reG3tClQl1uF3kz9aAsAzhHrxpy2o/cyDKdwUFuDhu7xT6g
+cDWGnnlgIekYMXzEzPW/zUV6sZtEIITvfJ3LUZSQeIizebLEeS5cuBsVUO1gCtEcnY1dxWcUcQ2
6FEfBazC5vqcX8Yt5rClXUnCNC/KT1EhaG+L6NQ7W2pM3kC+rv4rluEpSQNXae63jTVmyo6uM6CI
SX4Dn1SVaWwoMHgqLOfau7/6/0ArLQZhYsKxdKQQeUCPXQgKGoEloUBFSVcU5eONcH2vh3QKZr2j
/S9lcbZMf9HAKhy+M4s1RSisjbTWfzMzzjEBFmrJ6YhQpzRaqCiieRN7rhjfW3SD9vJX0Mnsrpjb
WoQcKNz3z3q5OlYqVC3Jvdq1HoLCz/eKeN+sh9KebKd1ooYA2EI5cidnKDy7s+XO4Qie81hR/91z
f2A82nOGPILzmRhfLu4pjiQGexthEKtvL7d1S7ROR6E3nUW0ToU/TPSOSoKk3e+53DEWreoeUHNs
BSnYBIDoZYheAiKSQSdeC/riSpM9y+Vqj/qEcKCEuEnhTlKMEU7+lIfS6uHegB44r46U3XUH3HD7
hn9asivpM76GIy5EdAGRSqDMaEzs1RhOw+GgLO8ZI8/rHjP92IGNHhNZfKAZH54Tb7nJ2r44hIxQ
FltfbIUH0epZiVHqarwWfnQyu9JEHrVWQHHkJiktAYP+VXzwWsbz/+3f1R2PJ2Lwew1QpqZi3ZN+
pqvYK6sXDxy2BfCh2TuEqbf2hyNwISm+Q7IDjRgcZg4gjbuFso6j0aL9SgX9mIcPCDl9SBRnGeXq
jyDlMvO4FOOTDiNhWBFUjbCnnR6u88BLQfOKxzkHfyEBHmHbFIhiq7+NtlaTJhLlqGDoDpPWkRQA
Cbr5ZymEAJvqAk383h7kPzupZL48g4QKxtLbHfocy9gRzC+vwq4HsC1SsbU5cpCzBcAaIGeAvFYU
BHAJAbjS7Ujp4exN0gDu98vCim/wPPEeJj87o5rYMjZEp+ar24yuVZKMWgcE1RdnLmujInbm/q+R
/D2ahd/EsHYU9LXsaXie3iJMnnOTGyseXBvJiSRN1n4pqDJMg1KLdHUpfU6FapHyO3aOxnD0KtOX
+O9Hxngwvn1bZh33rGy/6/s8vcPrTjBG4u2+oK6Gkm8FQZ9ujYFX7U6sF40AaWn4eGONNdDkzv0B
aPqVkzMsTVKJWFEVt/rzvhUjZnqiCJXP906d+WWLUYczWbfu8+0d8kb4BbkTlkMV6OovtOBy2cTu
tBgKPtePG1ffffEKCNslW7yjeYYhCzfoHcnGYl7o5IJhnTrNaF7IFJ46ejKOqwrdNoftaAVS/Uw/
nZWpt/aa1YK2vD5Z0slRtpKjy3wEE35+KfS906po9psxECuTw4a5DPXV90xFcHRFVpzXkzzlesee
AE7i8h34JqFIE/e/gJf8FvxOUGqWPcMh8NO/GD386GBICylH9VuZzo4NA+mqJCkYUzVHKkIfejKd
4cbCxCATssbxBukiAAvVHll9QVAl5O6vlsqSU8hIopV8HLIGv+whgvO47zvb11EEmtM1kmSbwta3
DQdvVgC/E7grZ7PlTZvDko78DSt3ImxlQKeY6cPrLkXj0u3mJZH8cR94QnaXZiOHrXxpFr7vCIJm
VvlbOIoZ0kUis3Irz6av02uyjtvGeCFpEu/Ek6pbpWLxjf50PveN4x1TrxGlS27J1Ci5/bgN3LYW
SyFB/2/4s6A3bmaM4xpc5UDAYXBTiJY/hHkDdwxRB2sK6TAJmObITpDYP03tt7IIXeNzqJEkjDiY
pen6b0Fn7Co0LonBgotR2ydtLa4x6yu015t2oNMRqKSkCS7MNsjqWIFH5K5q+8q6NoQ8MMUGMwpe
23DbnSvmU4lT2Zn+F5WbIz09w4uaH/xrlpa1HOBtnZ9hC2FbfQPZusfHG2bHtcW1hELvR11OOkNd
GsDm2K/8aYQB52/litek8tAP23eCyk/NK1NUuilNKVFxif1OMY+kI4uxISc21zsxL1njQDVVPfWU
i7LrBYd4xanAGuzZEBQhaKR8CIP5fnwz4x2WPKEr2Q0XzLYVwa5OnCLsVdeOvvwe+wmTGCRWSkX5
TIGfFxwsm1MDqtgAC1MzwVr+QfAP/6R1tGz60QECnK6Z8i4s36/coSh/TErZkImXbodNJ9Pq3l1j
G8exaU7RP/ME+8oUcqrZXbvmEBXLprd9X3ktolRWCFRcqNMd3ndHcyClkVqFMERzel30yep8Gj2+
qhqvghRFpNPQ8F1NFSEXWuZIRMOvTZslJbEZF6Nry2QBdlkQWLe/8J/9vBmDOd9MlrACsAF49ycl
S+lofbRJLH/G6lRmUOJR8xB7+yWcDstgyw4W6ZAonVqBjtCWWegO/0gyfbXFYUStBZOShVhQ9Q0U
taqJQNAOq84CzBF44a6Ilb779UaadogJNVeYTBavhDsdMRz5aZv+q/bUfMPt88oFlwXlXoV+yK+u
8Sd2MBPTrvGxKmbGT2De+9eUEBoqDL61EgL9qk6pc2cN/p562WCT9iv7qTUgiotrbpp7O6DREKeh
zpwYaOf/gpN0TzWN0RDtgoY9Nbp2PecZYTY/G8hdHxY/xbiY93l+rM8SPc9/njlITGlDf6H13gFH
v5cDwF66nxKaXq0zHQz2hYs2NmKoRDdM/Q94irZy3KFspJbZ93g4WcRAw4sItxiobhXD14biRM6U
8lZfBiBshsvbtyhqwn8IkKiuCgGUOBMh6vzoRPFOKxnB6Fucu4b97nevKWzs56huFOLUPh4y9qNf
zd9g8zLnfzF3pcAZZ1l0PZQs80033AFFmY1u1qBnhwI8RF8OKpPA02m9K6j79R93KZTFCEhYX3OQ
4OZ49SMmTGULeuPn6svCtAjlfsZEbN0CtakXjpm+lj4SbRYnmyvI/Ak9yZTJVjnSU9vmPXaP6hbs
wmUySwiRWU/CtexUdYbeUa2oDrHW8EimADOTU84pYvUx0EokJOpUYeqQoIZXuzUnQDF76PWlDrVy
t2CguszxKe2uqgPBDH7CzO59bystr98VUy/WR+LC0V6tsVRCMC6uuIm2Bp7HoZEcHdvkTCK2Y1Fb
CK9X3dwxPc8XsbjW2arlNX9RTbHMiPXKJehjyASKENsEHZFydB6gPx5pK76xvb5S79jCvhFeyc2w
f7mVrXDBL+Dnw3eqmgy5nQbplKnT47Z3rYn3yRv/4ysP1qkGluVuA/MUElq3218QyOFbBAP43tS8
4yzkGDp6gxt194KzcphASCSf1stBBGouvBiCFzG39pb4fH/ym+c1qMDJxccsCYCQs6MMyHC1UOpn
9z2o1CulLj349eTzaLTQu8fza3mGz54yZ5Cbbjj+VxfvyhV5NjTiHayxfKFbK6zR4IGGnkPQrIOH
tgoA8YPsyLJ98HEHmCXEg+890mXOqIabVygRjcGmGLZpaFab3R0Svy9doaZoIBfLVNOfpt9ZLOJG
piWbuSpfHiT5DRGK1vZVGko0koHtolYTFBeEODOb2ZqDSvlDX2zwgnJ/mWec/dP5+NjOlV/rTQn1
ulQ6Uup470h8Uim9rNkaefTyJ4rlohrXRx05mmOQKruoSWhnwU4pdpFfGDUN5KNzNWSLpoIWB7Oq
3obpsjs+wy8CZLN123eSRdxfl35CrerGrWut6CyUCfc3DdaDM43v3Pgd300ilcJveAxG/IlOKec6
hSmMOd75h+6d84SRB0ghJldUuLNZPe4gcPG8cQ4kyIlEa/XAVYFTd157LYFW7laTDHhkejkY/iDf
9xn9fkrE5ef6XyTY4rPBKlXzBC67mU2q0pdH+aGUKqSJgunYtQ7vxdQRVdGLZAey3APHh8TCti4h
LH8R+bMYuqXS/CEuz48N+TzBLZAZVodxfwQxHqsS4oZLj2TzU4guiIaFTtV0HPhReMZYXaGbvPLU
zV4RfSusnhKDgnS51HNBlpVkPWPw0tJBUp/cHFt9nbco2XJqaT0CmO3VBFWMwcZauvcWWji6+Hfa
I/Nec4iODqpmwTTk+issClV4NNyQQyCAgzjfRkEE89apv/Mpxu0dlDJ6jO7pvxr/LTUlFJCx7v/M
28LB3CN9K+ANxwHdcc5PwR7R00/85JyhhU2PSzEYCLz7EBt+X8uIh3Lk+MqBuB0qh2YMZ53lqtZN
BA7/joi3jtuGi2ZxBcOiet6omuQrtywvv1SKzOT8LHgZYTk9PZnbLU+OLt7UirJQ7l5JkQJA/qTp
YR9Si5hKoGCJ2+F7Hu0FaeW/wxZ3rhuiKvkVQgz3x9eGWsMugiyWKPTLEyA0ETjg4wTDzeuUqcb+
e7Dicfd38HcLKV9xCdAs9tvoG8prfVMDLs+GMf71kkih2X7X0WMRasDWPJGphPAjMvhHYPU/xGTa
EOYbEn4JZk3qHeAhuqPku/5TVPE+Hw39XZ7DfMXqQ3gfr/efCJwTPl+kSMLy3zVOWb3KKkevUgm8
i6WdBZ/Fqrw7FdF/viZtDoA0ctw0bTBt6sE8fAMe9LCtGKdHLNmcFWcipOVvrBOFXsk2eElINYWd
iPi3zqFg9Kog7WOI4vhShPnZZAmQh2LZpxVxx/d+diAcEdyUVh1ioiA1S5JZ4tpAWW/lFdRokqI9
NGPzgQlAau+SOJC3to23hozve7FAJ0hyZMhBwYjSdXXiRc+r84Nz3NTanRzMnW3qNBNY4je6GYvu
aRHNLI3js0qw9WJ+essYI8MIPFVXj+4173tJL7kuIfMn5FojjYWiyTLk0HjtR2TqhUbd8SxHyqbI
Fgaltwv8ogKR9dLFff366cXtsQhB67YgM8mi0c2yXtbRqZJNUWh3gWZIZ0Vbt0nLzqJitTz+Thtc
MNJVuJu1LHGBNpzkR7bi2B7MrOq7OqwDwG7oXC9GMMfEmxddj3N1/vlaJUOE9mffwWJy9Y1SiG6a
6PrrNNs1l1W5lXx61VNqEokF/H7T+29z6dQQkNw3gfLIckTzCclpew/u/kBS91GJEAosbVkUwzJs
bzqCvsORP4IIiLkSCD9RDAWw+mC3D9do+MTskekhL3GNkiC2E8ax7dB7WNe0P1fx18UMkKBxucZD
L5hFgDXcrM1IEP7oyqAixO+bbpJBVJnveypVIAY9Dta/ABwfMaT7isjOkV8M2rxx6AV08B0lIICf
T8NfordPRsn6ZXE4kktucCLpTMZ5g18UHZA+PTXOWzA4EtmpbSu86XmeUaRZN6Ixh56gfbf1Rirm
gnSBUfWCnoU+sk/Bt0Yp27CHjE/9VFiZU30lLrhPNCeZvFPA4jr19B/fqPLYlmQJMUegVll0xjeU
E9GbnBDUQ2FSUqTm0oDuyKtXj2f1FsC1Ftn6hIbNXSh42xL7Mo+cMx12q9g3OmrYHNVIM3Ep9e6p
XjByuvQYdjXWe5sGMn3/GiD+dxAtLVvAimTnVXx/WV26zhgTIQ8frwo29MrLip0vWhvMZHTlkuOK
V6AcROXrEOoV9flhWR+9s7XyUd7bMnxJRu4jyJtWSYr2czwJp320nzRoTYiPPDv2AByLEx2bWcW+
hrLEtlIapjs9kKwdEaWczMtqJBnD+HZma8+4ad84YqOJopDELvekTxnC5jHg/Z8X4gkK7Jssn/6c
Zp0+QSDhqoesitAm+epgx5kDXxqAnFIpfVM0JsY7zvBg9zXQDsXXBcIjZJBIw+wIV9iuswesFJwn
dSneuzYbLyVbFQq75UaLCh2o/iGl2JSoFOO9U69Qexvn8VQ7wY+Sy/wDnnHU0PBqHtE2lb9YV5Zw
s3wFKlrpt8+3M26G8ms67rdHfotCIgdavtkcenYQ8Ipmcum3FTIzWfvTwghevMJqZnH8bBzdWwIg
6XCrYdKtSWnrVmYKxx1VohOtKuWY+zIjpnL3/Z/fbWHY+pCvCUysig2TgS8qQtiio4IFB9RvR2vX
7IYiXBOtS2WO31kj5uXjyRSvl2NUKWMnOefNQXOfqXExjQh0FeaSVletYzrI5SFf4BG2O89OAPsK
09F6X74SjN9/mKn+vL+B3mRbsQcpCPEeQy014CPpZfy5bZqEk/97AvA54wiW8UyzwniKp2tFQjV0
O1WfJxMHueTeZjbOheY5+Mb8/+LiOlqgVv0sTXcql/j/4DJYPpGc/pAWkPre0OWgwnRZgvedRhXs
P7xPyCwE1fXw0zeKeOtoW2SXIHGqTNZDooJQX0KfY1OHDlokmB4PaVccRc26k1ddgYTlXcYSlNUQ
Fu9QoxN+eIUVxuuQrtAwGU6oKWoVfQX3m56RYAyHXE5zjuCEyCyXi5ByA+6FT1jQXUAKUkH6KABG
zoQwebsLaz7jhCFs2QS5uN/eEe4Pi3vwwWdEjlKayrZ36RGkSIwWDJdnVSx62GygjIpgdMw0QPNN
2rH7QdmP3KvsE6upLI5vJuKvJJjLD3rEJ8qnjAQcL6omWTSgk1mS+QHG1DER6dT6m+TQlAoQJdoA
k8MRPltgs+P4Q5a/MIUNXAeP2JhTU/y8tVM5h9+Xd/ekBu427QS3cpjimoMMpYZAFHae6F6QHWhX
3s2mVIefkRC4yM7Gk4zqTTRvh0O4TMMbRD2Oq5G2XXKAcQIEcihD6Qo/4RYuc8CaxWIjhVE023iP
n895fiM54At7Hg8+cLBT6ND5cKZcQsEEUZRVWUB7Flm3MO8zn1f6iThyHVuKfX9KsoPJ2XBwtH3X
bkl1OwxUR79KGrRfd4aoZLSIwwgonz626NYBwRVCBYVEUI0kqHxj5yTeR1JPkEn4FRQJUjmcEfLi
rb+Ic+WfqiOeYDP9nrp+MtyCOBaL8E+RQz5ji7cqzayAXLehEXT/TipOrYRm/axYxE0Kot+khm5B
LjmAWAdMXOHQOLBL5hoKYkVON/Z5alwQIVKntettALHEmrtITTemXVTFEgMjcMGGxmKEuq10BXvQ
SihXTh06GDAhXenZPwriuzFGRX8wCoAdNLvmoYg/TkabCjRODQQe+9a+Qchlt0+p5V25P1l/rLZq
MpcoCkhEic9GTDeyuYLy7ktTgfWjbH6/YPYAGhEjcnHIej5hHGhFa3zNkZtD0Ny7gU2dtxIb0pDo
3a42vY0WoVwBCmE9w1mYdUFy2GdXF62XzawY9Ihze5hzYXO8rZ3pmeaNIb+P/NHUGWZEUnS/tpIk
YAurwQ/KxUrTprrNcKFpKbAPNEjHHq/xIkI6/m/vzpXuZS4xz7ESry8/RLp+KT9yhWFUrUjFhNNl
7vr19vH214KpmMincobfQGX5dXdrdWK7o7B1xKNfGoqiqZYycoTv6gyzyipT/lut21vqbPF7HD+P
p8wKaAZsoLF6kvv78PpmF5xNglAO0Qhp1nckSzUnvEaUqSXFHIC3BwXSvkdyRExaAJ5GWjhCHN0i
cqXpMHtljnpQnrSzNoQGwHnNc56u5LsJGqneDSCrILh6GbXY8c9Uyv9k1fQ8hh/2joIpu4Ebl0hX
3qUeADAigbuQshrqFsTELdVIemRBFx085WscyIMNRTOZ03dedl7rkIujMPi0Tbqke+5/t/pVLQu2
aTblskmoIc4qArae8JuPnTQh18TlJKbBF6lKbdhXO4KfVKc0IMwZnXoJlNuxXrg/MmosN8ec35Wy
YIyE0Cs98qgwn18hQMS0VITysynws25CU1D/N4lSjp9fdZK5jgyMHMerujkgzFTgmtg6eOxOQjE+
a14RJ+cgnG0IZL5eVRnhQEuke2boq97/oCvxfMucR6nXExRe+n93dw5GQf3jQFVwKLk4fiyeJKGB
b+0gdyy0YgHrd0BlOjLTstwTHXIW8ZsopP1PZZOj72YaE0IPovM7Cp6h0LEPbgBPm357vJ4lUZgE
TYAXiGrC2F4AqT00w5SdKhnFoWipSZT+aRyVkzt2j9D8y1OeBT/G/htfbz52rsqGLjqHNVC9b9My
iS+feKlBXOalpA0g8lKL5AXQ/MK049S+p6OSptnM7+K0/9ayrTEPk/ZTeJ4v/p1Sy6ecr+/4mF17
J6N08VJ2nli5tnN169v8r1wy+SfOnYDdmpc2WNcfKEqkopg1fT8e6vbNg2YL6fPLUjUTvD60LpqD
Vh9Bwk1xXsEwfKzv6o/mGZjNfDhesw0Jx6YvQiyRIyOKt6gMF3hGQTyGJsLbRx7pSHLcsXwlDa5Y
BOEEredYLl3hIFIUVJCHMpfPjLbNITDCR9N0M2m0uW8mzJq3SpHWb4miF22xXhKd1kKEahEIXejY
KfvaRBCXAe2nE2zBYybPxv+5ogbf0nhKlvuu1TWzWkR1i37nga/RnALWtXoEOywnumI9kDnw/iEU
zpmP7RdYLysC88ar6jYzABDBHw1Qej9FpbDwZzLBIR0wy12sFeGwDp9VbEt8Q73cStbE3MLkDOdn
Xga3EezXWgXWCWCkDAnejtrlKKWfb8FSvfWNSyM+xd26qzpfWLkxJUuaDaYQvJpTHW/PSOWIIyAX
o2wspOV6/YPA4qS6seQYGecJyD/v8r/r+fJDQywSCKK+pRN9MTXle6j7i4nzz0JCexADsfRGAEnD
jLbe8j+lA7mrCTRtYP0YHxDuQLa3A4eKWBXluX0byDieyLh4TRDyU1oSCbl4C/rzoM5O7WVOy9L9
tFRnsmxGpP1brgEb4vror2N0cQw5pjhz+G7kLRUvnwa7BwIZNaU2Tlzz4lrWCIUZXCYd5veh1U61
+oF5Jb9FwmZsachTH6E3mtVxE2ogb3G0JgfKsL/2UkR6OgNHpHNiaOh9omVuQc6dJls70RFEtZWm
UXUxFMU9Jneynh8rl8c5bLw0oV4m3beJGVfv84Jeke5xBTXG1bCFAMlF0+R61mqqWMZGUr3utlOM
dnziJJknk62xxugeWDKuTehy0omlZ2Vb+nDoEcNsJNCCqmcJqlP5CBUgYMyMIvu+6RnK+NDILw8S
OiaVCnTDZtaWGmZGXd4yUBz2Zfl+QKUWqnbJK1tKMQYryomo+uB8zGJeCh5WGBEZXC3Z4QE6Z9Kp
qb/6au1GkgsujTbmjjpTaF+2bsDKQn/pOYylIwrxXWXSSIUHBG+52JwZ/W5BucSDtTRUnlPGYR4E
rucf52iHr5oA/Hib8Mfi2EJFtXNpnSiDOfyXItZMdKwlYilvpqenejx2n3D98SMwGl9Yx7dGO593
MUMdPAerrENidGI6h6yzTP/QNIZpiNFgzcrcfDNxkkVngc/BTy+Y23SGZlrlrU9oY0oLFWerzlFV
d8zwvMI17QIKKnYAosYdHUGWi0A4Eg2MwWpsC2s1D0b4rR4h/u6oMk4MD590JGdp4cxEeHH3QyGH
cIiiW2vGsxQHmCPYG1hKs4S+mcp1NKSctwGY8MqMkoSbohg2PRNfQkGQKhKDB+R6hxlxEvQEGWWX
utiYE11I2w0e0t9QCCl29chjKzgwfd31H5QPjMAmCkfp0hGBWSh3uYjKRuwsFAKMIGFOIrWYvri1
pDorY3b3EDzdOg8itrZtl8jQqAIgI4aPL78PrvIoN9MmF8tqNv6blbuPFz3ziSqCTRGiR7G3gKNO
3CxsqdY/VHBYYWdYC0EI3lTXb+1NSs8E4viLywKN/r3HAlxT0mplJI4bWjrLJe6KDuoDFpbqpAcS
LyKRTUMI99qPM7bjzA6Tuwuxv7kt2gTV2Rf4cGqlJe1fILo694kX6WY1ueTXStbUyopypMYVRENE
SNQ9UfrDFVPaaGNBpJkPmMtThyF4BuMhlbg3Wbctc1BSy4wv9FHXrvgdz7ehwsxbmZvf7OtewJBX
EzLss2kgHh6xBwAt4Vz+4gxS1AfFtayfWxhzhVb5pQtVM3oulBvXomslsfMgBWT6mCbPmbQzFsiv
yMslB/QXXyCqPUw49a/JKmY/eoJsljMS/7dVncVoyalvgzINpPOaK9SQRU90XmO6VpWdOv7pTjZt
kv0FJR6JW4g7baguDur7Ednyn30iRs7RS+XhVn95hp2QTRHSxMb0Z4pukYAyHmrdEv2zB5d93abo
GzwIuse8+u6//ZcXoKb/1hVL66ibzyoBprv2k7pFZNDvQ9RY3wJ2oFTw2IEvkjO850pFvy6T6eTe
ofK4e5Wh/IXRbMqtQp+MdBA/3KLiTeWAEQIi4MXXx9faO7fo9HgC0Cu1vCaM8m0Fy5EMTEfiAeJD
8jaL8EgoyvJ6ioyMz61HVfW4ygBGM/yoGNvG1GNBOksEE/u/5kn9RBYYO2d69Q1/bZ8afolrzHiH
JT9dALEUzLMgWgBW8SmcipjDYS1fGxr7VIQAUpWB1xC5UOcvTxAsFDNFFWfM5HiAvViWMLt5pykY
4DNGeEgzJBak1vWPKJQThTIZqEPcv0b1Lb/KdVf0aCeuyKVHMfdtEtbpz78V1VK7Y4cyplbehJK5
QFktIKKP717qUdOEFyZadAoecB4TBbC79d90zjSslT9c38sClflT88yyJ9sKRTiNOEq+2DHs1nkx
xKEVcO61uT21cHS4nzFU0IEJoBi4jj2nAjh7p0MYrAjKgr3jKfd46pFAK3vSX9SsQnC135LVul8q
VG5tv748mCEnMScXNwTEQx7HmjLiyCOkC/MRdIqrd5rrdZhBcgfIU5cynQKGteVo/UuJoWPoLcXd
99U6w/uFhNx0BAXlWtNIUrueJk7h1CRBrNairlnu/8UsCkjD+dwvX5yqNOevbK8chuZ6B70G/uFk
PwqySmkbxyuZlJwA9705H76p4yinlWypBu1XDeTANetQGLla8UnIUFShltfBa0CEd5GSFnvxINdu
AHNUYNpQrAERLhY6RKID31NLSW2Cg5/+WpewbEYBpPNi5yyQOtWME/P66bkYw29Y7fcd3idWtY5t
JfagoLronS4CX2oABexSWfbHZ8xo9vtieJ3gGPbQ/2Hg9NQK/CRZK2JqETMfV+gXkY5gw1vUlG8m
6BoKmQfA+QFOPOCbULr/W51BV6kaWdp5waxH3S8AUNswiEtUyV+OW/jhRHPCMuDiBE0hkfUT0oId
d/31H3KlSVWrm5fERHFTRvflR2NrVAQRSxyCuas7ln5PwCLcY+pcMbOxx1AiQjBmffNKhJ3MA9oV
Ffw8Qt7PnIdlVRE2FE6OOkQY65/xAFZzlDRSQHCltpzLlnX80eNcHq9YmWYMpEw4D9qDXqmclxDf
Rw6f9/+GjIszMOV/7b7mJAcvbXzPPy+252PCbF+Dw1Znk0TZD23jPnJuTXD1oP6BXW6j2vkXdjEl
Y+rF9F5B2zD1Q7FFllRkkVCuLqofTwaRZXeQM4NWB7rWbgILjBa6dR3Z3h1pQ1ryTcoM8ss4W6RF
uXLowZITS0Lk21+7bebntGP9l4yQ4vAA8qQ38mmUHfVD8ztsBMcue8ntbUyjbyxvjczAfzFp3Q0Y
a8f17UsurpEWxo/D7hOJMFs/bfleeW2YjBAYCtigq+VaZcDo1ucuer0YEwsnWtTbXyjW9VDERpvu
mBzclwaTBU4ZEEw3QBfVZoiyiOgQDooqA0DGMZ27iVf8cPLGjFJgHBhvCymGOsfSqorKlrcBSFNC
UgN9rH3Vkh0M+Ls3yrckGWLPoCAhzb5ZddGgC2SIyZb0WXiw3nAAf0zlcQ51X95GzniHBW0LUqPC
DC8IvJEzfhMU8UycPlLJVV5JdmBCo7Pzh//ARDq2GQGUDNo6O0rRfwrEgM3FUK8dVqcZVOC4qhYS
0J9+2yH64UB6FyxpAeo9gjtUS8VeaPwbZI5MKg5M+Z3FWiYMAT27nwlffKzWY+HslSckOOK3vXlb
v8RIzwbaue9z+69CYhQQz3Gwzvg9bNCuDGF3w/ujRb311ptBKV3mzIbzwNJ9ft0lK/EOWcAfputE
Tgp8qSk8OVnBIgwe1/fDcNA+XvRMPo9CQCYI6WB06NGrkyhs7qPS8rc/jpTrlNpzmWsocmsgx5M8
HDi1lK2JPWflGP6edhtdA6Lmfa3VLQO7XeJ/s8/F4DSOtfVyG2xaIS3LgkSQc2pyAEzjruxUH+3A
q96hBwKmNc+/opUghAyJj951L1qp9rs8u1zt5cTAp92AxtSZHeILTEXqqVnE4SycCZOqm2ZvL29x
+xyD7bb6VNW+E1dsQzDGmkZ4yPAMCPFDMbllSm/g5IhGGNPc5lsL/4FM1BIdXQEkrj2R9Avk2nuk
RWQ3+uM8m7SFpRJmSeMuWRhxHMuPLNMkmg1ysx4kuYyBmjOe5BUBzNPZdLYOe77wvuN4+PQsUKKB
mmGIpCUkmMb2TS791A6JYCh5l2HCaTmmSDIL/1wNc4AJIFBJtNZv5yTMKpyF2Jtf8yjbfOFSUznA
PQUG8yXgUuxEn7KACVmzvrNYJZ/ovGIwdfyIa9TDJuxvV/+B1fOx2EkyWizz8a7dV2sJTrxI4SCz
EbJLVPBR3tBu+nmUj5hUhFvObrDoVo9jwyrZgBV4DOgCYZlc8GPuG0tl8Z37mKiWtl3eI+oZpGLe
dTVWqd2wKgytvxqey3KKwrUM5yM6ObxWRi1c4SbNYzochlcuF2tDRhPl7gJegku3dGW/Yomfsl4t
mX0cpX+KaTAZpYpr5wUzTZkW39ToEYUUFfKSDamiI+mR7ueOfauE4LuB6X337V2UrV0ZBMsrW6wI
GtXwBamNAIXHVLfYGBGwWrgTbrcdVR1sDvhfzmhv5n6ZLPkUJdNJxowReOLlDdmovTmChRlHtegi
nxi377R2BfBezv+qlclt/OumCz1EZ+ZkaS/spqfpitKEGBWF4kdC6QKowfPSHUU8KUwOI8VukZO6
g9mGV/prsVTEMX1ymNG6ojc6CH5Yvxroh7Z07Vw2FrjYDOhd5126GMD/uyyC25dv6v0ELFUFCgPA
8ZdTeZ8Lly5EK8QgRMEjXTBNa8mhbHATFUoA7rl6M/PUQvBz+lezOxikcPaSL+RxWCGTe3vP3vaa
/lfHhf0HWnuqhv/v9gbC4BmwMCLzl1gT9HglDdDECgwYS6Yf4yok8qVzH+X7ZqdyMeY75yma277s
XsfW+kKcGDAEOfgdaEO0wn+kcMmzBx1cF1HNEglDcq9U/Yt6aJ15Ca0rOOcEA4XRoqpo/ZQfhEjb
z85EJylQirsKPs6oODnQPPXWIgkcp0hzpflEgZ03zZmdtOlys/aV1KmU9PvDIT87bFyrBntlL58x
4MFUfkngJb3XS9rfe3GHME95sD03JIIDGs5DANgQ1iX7shYYa/ZlA0O9kDDMIlyqlgb6g6YwepJE
enSuMdTscEZQFqq+eJ35JyjsFXbtSttgLDqCP1gEyGjv4/WHNKDWDQt/6wol7Y41yIBrUH1l8VlG
Cmc5NWm0A/X5D0el02PAK/uXyOrpwSg9yBnnKUIpBqp+PdU7C2rq00XIsUZDCOeK1WFdkl8kHn6e
cIIWAtLj6g4ch+k6bLQ2bkUAY3EUy3AJAtVrzMfG4XyprEMfjn5vNXl9Oicpzd/RtI/vcC6pX58k
XkQHslPwsi0JwIulWC/voghgcmmfk+6/HLerjfAo3VLv8TIL5EzVSrByNvd1A1umb8zEvPtWBa1/
21K97i+2J+A+rQqJTkS8EIrNjH54Kc5tR7pfm9PAumSF/PVhuGmgRwDuzvCllk+3DpscbxqEaXS4
CCmXbU47ndrC9DvlWUtQvUEWKjE4hzolTQPUNRNrS/qbBZRsysziRUqITq4cNCw7MIpTv0olmOCf
Rrt0xTl9LMlFHdlIR72FipdFw/AbW5vyM5m2Gaf7Xg1L60Yy/AJXnQl0XX68sj0jgZnp8upB43bi
o1fbacOUQkZGekTVz7bGf6x/9HZ6gVtNkcLanaS0KduG8N+2faQEg5uu627IKz7Kry1lXu7n+STb
m7QnrNTPaHpYq14roIrXUh5wPiF+egfwlDwNzMS+UDNRbd9KxuAshCP1S7FS+6NK4079o99Tg1gm
WJrAlQ9tXVji8c4ffLn5iejkAOvVA4w7GYwaUJZjVKEFg6C+ksQv66lDa9P1oZzC8jlr4WCRWRcI
xEh2hpUJ1haRu1tDYfK/Mpn5s3rJYJNTa/pS6whaStH8TYhM6e2gQnMocp+S5n1pf2DC0BzVSBdU
eMCy2DPeMmLMdJmqAoko5S6t6OlabnQnyoEBNf8JSdgyIt9/D5K3B105ui4Kb4FOO+iSDFsMqUZE
wdCKvlTDyTpfZtXaVVdVzMqoW9SidGktR53KH7rlD68L7OoV9AtA/+NS2F55/M92Eq6Ksl18c28w
AlbCwYR7IG5LP/ZnPSLS3uVj6lEMmCx+wgLP5v5XfKNnuO0lG0R4I8+F57IW/n2zeLApLYBNmm8j
xZ/U2z84+PK2v4KQDljZmvxwR1J3fJUwVExl7Ih2RM4LwBQ7T7HRt3+8qG+IfFQfG01QqQoNSyrh
zgoNJ849kSv+g0/MPseBiWqDU4xCHRieyUWIlxcwUim6DIRtfyAAf0WK3i4jeZm6C5mdmwwymk8e
TtN1HX0HzdbUeOEbc3hAskfBhD85BSftA8cGqRpwm+ho17EZvZf0I5SUPSlSe0s7gBuLBLNtKxQ8
TmsjMfKZI3mNVRpFptmkwJDuPigFTlNW+vx7QZzOO+fSSsDtyAkbLqx74UlYi2Ybs80TMUhANery
nZQS8T8XlD3hB9WEWzU3NQrN4Et+LLFbuD3403GQh5VfOahAT55OPomxUoonG4fWyE5QmUyQLPbg
z8L9pSYDidBPaAbUt+isr0W5dnWWKZ14oXkRzVyMNWSAjrVGBqYyQEHwU1k2eN/k9Q0CN5GWVZO7
4RxPWUQhGGHBPRjpsNH0xKdo9yAzknbszjoqg59dkxtTnvMUBh+4CK2hjeoLf09Mc8WNEA2kIJ0/
9b1T2etl2ZDmOljThqIBY0xBlpnHkUsrLNOE575D577nPNHtNYjHpU3jie/7Ainpd8rS7TCJKhUK
vux5efpQ80cwzPtwYptwIkAW/iJfm8YkEHnmEzs9ecv4/tFcqNwSCbBO0alJSUuYsuz7aV3EHZ6j
FKjaYHHuU0sxOE4Uu0hCIv6Ihbb5RRa2Cqx5cnEeER8qfCC7tDA+PWEqej8wK6VRf4v7Me77WhxC
34JtauR73PDNjtYdRxuCVgWy4F8ESMbFaumcHjIZ4Sd45aM1Ys6Humo12LfY+5TuzVu0NXIaxieg
p39xRIjGpA2nIlUQrKb5Oj9vSN/HVMVV7e3voWXB0F5xkHgC/UQ7vGwMEcC4pasiD/PcdTWEjTIF
/dXwlAqmDD36Acu5bHlyB4TmOZyKTM8HT9lMxRy4tOdfwKJyZdFP8gWxuftLNIgBs15iKmjVZwJQ
Q22ubRwTvzkc5XyUYOFKJvg1giZIXZRKQ25uhGkRTL5W79fwqmGYgO0bldiHZZlP2m3XkGspKJKs
viITGjK2u8HGC69HdIwzWMYhOx516PtODCd4mekFR6wSiD8IOnxpP+/yJgJLJ16AsC6jM4lPuQld
HgwhaLPhgueCSL2nxGEJuhpdhhMhDiTy1/upNNHPrGUwX+2orP40kyqu0jYeb3pISbf/GJiQIxlM
0QPvOkjPJE8ADKkW8Q2cQrgO+yOXyMWkIOcSll3FHCBd2a43pVCnRUCY6fLZj3OJF+2ufqe4PQh5
fcORAhLoFTFy0nefDJRhJAXlDUIBEoR16d62OO7ptxr5CLEQmFgiFUTlX6MChKiJa98yDAvS7aKN
912d6nRnSzEoiTttYhemzlgewjejw89GeJz7WSoSbuWVTsTPAW5ypAqSc36y1vz4Udg6++Yd4Cei
R60uJyaHmryCnQpvSWBhNcIHov7QYoKJQA0hwWSV1V8UEY8sp1mdSguafzm1HyJVaw4J2/dKzHJ8
7gSq4q4FLDXNLfqb4ZA5ojHoFPUfniHjJZgxSTnU5FvMTm23BLCvlk7lxIfnUPI84Dxolzj/kx7S
UeLsdNrN2hVk/mJclHH7oFyX0C6xtvgiAESd0Vzab/8hlcIHgzhov67fqmWsX6nLU4kdVebBc1sI
GoRPu7R/vDv1QV3qq+bZ/WONhmbXjOSxQyQsbs7wDIZMz/Vosq60lcX5fRpstw37o9Ph+BwKGXXS
PuwMppfuinMjXv1MIjV1WrWg9/OWZVZCuYpzU1JISUNm2RvuKt+VzuVog+vmfXMljsA4wyrN3WOt
X4Gp9YNAwTQ5vZzNf84plZCq/wSIFCvVDOciPCuBsdz7nrruXhbYuQHGdc/L/RGbsbXz74Qx+lbg
MhLtkQtByhIfHZtRmaVf4ujiL49+/5LAzuYjKAHTHM20OHFfWzvvpQL0zZv5KT8HaFa7FF40jcYI
AwS5AVs2ifqyyzfYsYv0dPSYO2KvhqQrXX5BX7CuOoRnLM8n/V8G9/wHcJDUI/Mw4krRABXCR1DO
preuzpAo6YuVCHcfFrfTDQzIEOgBeZhEQgr5VKgYX1/sNvQ2d4h2l67XPj/MZzgRqDwWqvrMZ5XQ
sKdX+xEYBxjyAMgGxnouXr9c6XWtWD3+xkPgq+ITK+gLzESldE5+Q7QvMiUvsWsc8lsFIXMyoXJ7
ypELqyZUIvhDRiIxanharkmJQT1M3FTNjU5k3H1YlV+SAByfGuAn0slzfh4tdnNNvydkx0AoMw2W
E3EwxMFIwsPl+oOLpaNkVwaAq7z/N9P1cgb/qj+mcbAYObZCfBHp+AdxQtBtOIxDLWvnpPoIO3gz
OdCgLMvHnl/JKHPZd1NmDCFguPCuXU+bd36FtQm5eYQkshyR7VFd5h/b+O9GYoccppu08KVaWY8i
0hH+aUoxSA7NgBMhtFTTB/HyqCNmbZvUEMqmVHssAZkuK6o6Bo5DITLO+9BqgR0Lc/IkDmNfNUw6
aKSATOTSbweJAxjzMs2SU6PW+3dojmSHEubIwrmOf540T5MLf/7UrejxiIFcaBK0C/TeyUdrSjLD
sv9GtUIFuroaY9NLtyz2ULrz4THbQwA6NMcoDUEWEC5PC27TMB3jZdcPCn1BtGwMVIZzyYXgiN23
o935m/CtbzjFq0qr+zi+HwhA6g/OGjGQUayV8SABILBqmVmpMzCnq3S8pDvPB4f4X2PvvaABOTP9
fyQ0qqyfJT/1tjwNG42RryupkaB64W6QdVoldzJDNWcfBF8K1OwmgFoRg7QsK+KqdJJEbt9FGeSm
NHtG4NltP+zLCUYY9ejdKH5ywB3CO6kAIhzmwA4PFhWgWZ6w8S/PmloCUGiudtPvZ3alPNhgTvld
gNHfv9ZxThy4P1ObnkKrFJzLTozmu6kH9JyzmYlawj4qRKI7P4HOjLgu5LKrTRhrRZniIQw+hWrA
Il+o0DS1Qol1fVZNvstWUMAOIu3VzkEllY2TuF/iDbcgnriF4WKkRu/rruI1bYUOF17oqkVEXwAo
MqLF2vsdRvWDUrCInV4XgBw3P2zvbNXmimlPeec0ijqtw0P14uh2ks5/2zPknIeYnRhcA2ixcDVd
kHHBpNJjQrqZPBF0Arvhi8768JA8kc5m4DrbGt1SMrMkQ2lK8WuBGxhoT04703+8Q4qfkbx9SOWz
Xd9x0j9VtrlGJr8LaSQPElrJf9DaSe8EPj3C6JahRArQ7rOonhH2HVYQe5w8OhDlBYa9Pe6W3HjN
Pb1QXOP20ODfEscLdGFZnvNuRLPj8JYdydwpQiQDxXJVEbzHLl3zqwsEPljoO7+0H4+58N+D5DSh
Q+jZThhPDwUXt1XQadEMRj09V2cNgvTdhSPZYtVDDsxuBGqiuaHQdfbOxfmoPsb1vveatusgbcxt
HHFBAgRYspF9xjV8QtvI3tKIfCccJml0IG4/qqGrHoFOSQ3oHF4wjqbJPSW/Mb+ikKDA66tk9kkS
dE9qiydcB/I/31kDNXMCksi/F1daTN2QTQZeVVFar4NmKUe6762fYZMAPfRFdgl6K9g0k5OPmwy/
Z55nuHQvWadRzprzLh9rFGayeTUVDH1L7HaZZ9wQrDV+iamgK8uMVRpXNptXBk6CQCk14lRyGuDY
a1iyu80rh3KXMWSqk4dEOc/kEf3F60VL6BciifoVuyg8tuiZpxbqdCTtw7yE6foDkbx+tGAORmVm
UhlU4w/24ZySQlZnXPUheSHeytiSBDYRWQyw3xKPbf8qTe+m1XFRmDDS3jFwcgZSyHessMRTXgOV
esZjHf7WG5shbaoeahmbwi/x3bP35R2gdYGp/5CqGs9DbQdbnZRCBqq1yJTQcFsUixoxdXV+gp9G
8lfZ48TLS1BCK/FbW77fpgM2tywyDJYR8Id3sChqqU0PRJhIdTzbY8WWVLXu5iL08agwz9T1br23
hpsbfK43+zxyxQB498hDAzacl12se0+pnE7bcUJfx7IixpmEqyT/HZ8rjQp7GMPzGPadWVH43vWJ
ex4i1pxATpHUKup0KeZQf1PODlSSc1bJlmDa7fP8wR5uYZQs5NJ6c5eow4u/zXYunwpuq08flSnI
0OS0HJYv4xG0k4fiQO2n1rCLbFpfllCCDRBQXg7tCBrUz3Cbodx2Kv6jVjPV22WXOkLpSBe3QsW3
cZApiqddXsyaYEm2EjzcUHH1tyRwaGyE4CZmyekYmM+Z20aSQBo8hcBxuw5oGcsesa7KF7QpzPCw
yNEmCYRkt6ZOcxI+XYMmkBCorJnAhB32XOqkByQhudhAA1OW2ruci2YDEi2LMHXBkUFQJz6JGcGD
7wpkftQMeaXW1PcU8g9ABe+o4/tLq40QTSDDTdofUxSJYOjEMOtDcGLzh74cud/9vsaT+eVJew0i
MOr/jP4GrWur8k2W0M1KGImtjBvRQ4+aDWn+WcbYt6LJTIH+BnseWnTC2EwFsV0hexeUvIGMriHQ
qg6Zuc88dQrkG+wurfOtmD2xjooLUdB3hpN75IcnFNYGh4uYOKCaq7OsCGW0/fHNrDKg6zOlb5QO
PtSd7Yhiut5aGkujVXA1Xne06nv3S3GRHKuSQKLXtpXyF0xSj6o0Hz36ysLk9XyjWRfGiepPGZBQ
EEKnIWQRgSZEUUeHxF0ZZU1DBfvb1oLpr0sWZJOKZgJJ3jLclAgx2ZqDlp8WqqzxV4CRBaMGkYMs
7oaqvMcOt67O+tobduxCJnyUZQYPC5OL3gnHHE/ExF8aaD6A+/78mN6ozt9V4R9Jj61G8Kf1fQmZ
3PalywoKPe2qqHQbjFqWdpiV/NjeJABBEnne2gn4xU+YVRtZlPQnqY1Auc2Y6a4rgsq/w8AQZ7UX
ufGuJIfxSwZRxUGs/CvxLjlFX+f+fmhwityQe4r+XH72AK0rAY/hMNZ42n4Lm4lcFAMGNHsAhkuu
vk9znnAIRhLTPV3NQWzIoDcYOSOGZfYCwaYzWlssVWWO5y0sQyi6dJn7A24xtFgeGhYs5KA56izD
m4R4b8DTf2O5LijE+dSNnFvyejHLA2d3WhlyD7gErjLKdYhZ6QtsFYHNRDMI6JIUpnBHkP8UuArF
p2ykolV50whKpl+w/oFB1WyhTyPDqNcj3E1vuP51l6c8tsx3UV0EYGDjWGnXlkx5lawgZV2jXDqE
hPByG3I3CmSOpxWNX/D6B+MWOWiOqAFXvwOkYfF8zY4z+B+ix1zGxLcO6lZ49eYpnrO3syEEjjff
TbIJG2vf+xaMHZAH4cmu9XzMe0/wgBsk+L7eIYGb7XpJu4LwW82zRFwL/7I3rF9Pc6UZoDbTvE+n
Of5CtYJQl2KQTsyiwV5Q2h7iZWYvvmwIdwkfjl9hK74m7yVe2JgV3TQNzVn1UDUXFtPZTvxpsgTH
Lwktyrn3vavDJ4LkAtMBrSzAfNfsr9ZAkHLVQEQdPbpjndDx0SCZRmHjIlP4UEgyqwBzJlLlKULb
su3mjEf+HqXmT4GQSKWIK3C8xa5mVD2nEkYrqhHtPRT8XqU+hvCgmKgavTerHlgOeGOk0WMLemhk
+SN9wmKzUcqT5wKdVPaHIlr5nN5tBJIGYCUVQxzxBW5vLz9X2Pgthhw0/aJ/3itV/Pf9jmKjAeZm
teXEKseRZhTUWy3jV2m6+zoKrHjGDqWYxZgeMrWXiqNuKsvpbRYCVVVfwcViypEhv0d249HXCoKD
30/LKaBYMF6P2de34skFXKovloOUPSNkCPRHprAM/9bH0BfYbV0qM9/MWfS5RKsnVM0SBuTAR7AO
8/zVLNpNgfBHqCZBzMTbRVv4yOW6e84ToL0Te2VeaJpxLHoAA2yIuLApVJn8Byi7sEprDm8gBnGQ
2SqKNGXSU/bub8lWiFW2l924QUIGaXbkNLVZ7XX4kh1Or4baJ6xwHb1hFzDDhRGAKWWXWjvPElRm
onXhLOiEQvQBbyw28tNzoD7Tl3x081drBHaBA11LIphr6IasetBmbR14doRz3metPTn+4VLJsPyt
7cNISah1xgh3eiPMT+PiP3xBpgWzr1OwMM7C3L7CYjoNtMMOz2sySAOAqXSlhZKHdIO1Hc3kR/CN
IflQBext9ez8u6iywWCzZ42vECocjzEbLf/XcACPWjwhR51itKrvi0NJXlgOB5XeeKRaqT+c3XLo
phSKgSbmIgEeZTjhmHBjcbLOb4DBzg1V/C72G4lvrJuwS64D92aHoRsDz0NcPB2jsBxeiB8qHgR+
bDb0CS0HAExogSHUFiTx1CifSf6ySnpOBmdC29qhhv3pk613dcFmYxUAwzo9LPhRmwJh1X2jp36/
JJkjQCPjqe+SryNZ82e0kvr3uP7V3SCbzYHhaGZMAZuuWVJYVpfDVUqtSnF0IaePNuXMBHZ9tz4l
coBsA29zE+ra3bwjoeKyNWj222Y9+WxSIq6mYgTTn5jlv//cp/WkZEB1zjY1NU6/PeX8DK8iY/W9
xQGhtgihNERmwBDlpnSltzB1HcvqatmBdwSwQ2pdoqlCdWpey9k8aUf2BiFxSgHqFCpTM4rXl34m
WC5QfdNFultHd7I3lbKXmCv/8bYsnqB4R/qoxNh4kbvqvoMRavfbDVGJvStjxWk8Yax6UBM0Y4/9
ffONaNVkiQJw/HEgLA5X7KFYyUaE4S94uNLyME42l1d7EwCRLqG591gTNfmHHrRCCnvClhFonVpM
Jbwt6ews4/R1k6T9AUHbJTdwF33riWe/IxhdoBIJuKjXrpB4pl/hFQWAO6fpuyMQsLAIZTVySvVw
5UWRB8Gk1yoh/x0PuQIkltf2R6aaGb1C5o4kQiZqmzr0W2pPzuy+BUwGaLABmzC7zOnZlhlU5fWZ
T6bkctWoruEoYmPM4ToQRecPvef4d9B9fUyNkFgNgHKi/iW0IlAIwlAhKHrf28zDsuQ+e4JgZxPQ
JCQ+7PsR//QEaig7jYdVTcKPTy9UhxsysNVYNvLfp1KCRwvBUdE/vva1QvYKxyy2obfI4c8Wzsy+
ixPDELIQqcHdoojM939nDZeU8rPwDO6e5WfjIbRlUrywVfS4cBZ40witwbODKvA1y+7Rd3l60OlJ
fLc28EY7zMAqZM26oWwrh3LWgzyMcvXOfep95sRmGvZyn+PHGU88p4VwMBIshf+yaNWUkH6D49y9
1zTE/Glu3EdyOlkcL9OwuXjDBJJu1JvXU0ynW6GSsJP29+B5q8oeotd6SuHbIAoRSaZEVq2D9FQ+
2gVhpOOyIIBEuymYgQNDX5HGz3IhkjwF62hTqAGK7+qgF5R6SbVfIjmKbJ/NIjW93+8RjBbXJbHW
8z25dgxWIUoun2m3utHl3XUJ+uqbTrmsTu67WSnJ9FikM35EktQh2J+cQK6md3sy8RJe7jCCJB/Q
X79FCxcuZ/9gbyoTf2/DZ1/mjopzEMpoKsrgUNZsACwHq5u5+AiZBzEYL8gUSnR7tVzorh4pztaV
jesj+1mMCgtff0GH4yE84g89MT73bN7buzp3SIBiWo7WIefABUnFjwalI9Wl6TDo48Yr/F8wZT1m
aNifwgr7j5A/YDHoohwZqmT0Wfvfdi11kQnjUaECZ9MowE5cvV7L4LFIgsy6A9e1XBJdxSioVLhu
5KjBxev7J0l1QQ2Mkc5QW9hRdzIsH6MKK6ZnskJdFKFJCVBobgy4t6/FG7kHJr3bOFHP9u1z/MRq
/1wK6KhEO6Mo1g5GGymJ1h4QYg0fTg97w2gU0YNQs4VY6k+KQB9JGCAYD6FA5bzoSWz3oCbCMUva
ra1KuQtX2PNKvjQzvLW7Mc7mQ2rrxyvqCLh/bVZzMx27iu4pBWfMcmP36QA+OVUiksGEqWFCWp/A
QX+WUVQdaaZgI3RypEO9z20sLXoFGP8g1fKprdEWMVP5fNVqt3PLVddkomWFew1ZTJ8kAJZ5a8mg
G3LWufTrGa4M5UzMSbbqLVXPI4afZuvd16oQhTZCZPsQyux152I5O1WVJCMg1dlxNIq/AFkYPXiF
JZUsTqo8fHgohutQJAu3195g6+Rqn1LpRubUHU+LKaVigyECUZtSeBm9uqokWwn54uwIO58bqA6a
EkFKPJupX+gztGAeYNpsJZP339OO6IPtiWwZg1fksExeVSyT8h24BRGimMlj6j0i0zeSCN/MKKCa
AhHiWHKlZi01480qQZTpLM7o6vcgsyJr5E2g06uJN3QSjD/iF3YcyTlqzWBvHKU/gi6q/e4vdUxP
z2zkvVmYeT6N29E3iPA3hRCbQjxSNQpnO8ELnzp8vghyBnTREi8L1AULKxqV6DU8byLxScAwkZbH
LLcvoEFLdposlOvW6XZjwMjK/vapkTiUwicvZcZWP/j9a2lykimGi/1TSPusFz3tPG/cE+iTp5OH
Yw+eDcPz54Mcd7pvNI7jbv43/f7bhm5s3poxnPfO7lLubNy1J+ngiGTBxB6RRdE7TKXf41Z3c/KN
Uks8RzHPc8wIa9DmKCGtgaqxbZxqi0zRTSBgO2cKWqevtefjgFHgGcAYr2f6PyuYALIpmMKWEuPb
N4Y4KbyeRpksg51v9rerX0DvX1dUcWHg4wQdtH9zQjhcTUES5YrsYw+7xZajUCQ1SuL7Kz5x8dbv
ZjQlGQRZ9abnlatrHxpjMT/ecIWMql7U/D+caeLoQQwTikWmKSp02sV/4t+kWQ72N66WhBpjrmYL
yuMFEof+cvQswjhBJSI1rtS/EIUFoRsgn+fGyrwuBG6lT0Ng42+TjSdGn+dLP8Ym3kX3obPO4HLJ
qrQZq6rILbhQVT/E/kgtkbJoM43D+L2HHtAKMqbekk3PY8gZWIitvmSYczokY6DuUMo3uSbZJ/gR
NlIGd6/HB5vdiRw8KpZKGxseeRqHs5wpW5IsGk+LQ0B/iXv4u9YBYC0J0Mq+7zu3Y8NL1zin9aj9
GrqGJMQc3fY0BTodvLGWmTRaVRH3UDN4RAC+Q2ipYu1zv29TnALKPc+lRoeUIXI7cdonvcdRXNLV
fYnmspvP7blYuyc3JYA3OAfiC122kiYhbtzGQ+4QfjNAeFmpNh5B8KxIF4x2DADxnFoKjNr+ZvIk
bQhzuaKdxYsRDJXG/nQTMZJc/JU9j+4nxuq7/VjBejPzYFhunaFuQJxFxEiYYhEi1IbYuZKL0kg6
coOaUpOBUkl8WozO6n0BhxcpPwaBSXZG4D7EI9/EDpukrAmb/KZ50MIh9LYgunefyCSCkV0anS0l
v1DO5UtraHjSLpEX7bk/UbwDJwL5uv4FcFO0ctn2XH1dApqPh5iJEvZ5YbicYuXrJkNnptZXRtuP
dQlPVA2bsTebNfovY8s/qM7hH4/S1+QwPilD/xEPAVkPzAe/R7wr0kpMKsyEQ2SXRUqZRmKQqWcd
yB1AByWiSf7SR1vi+z/iD8GvUS8WlwzxdBVoDqLti9xoHougXkTxYrArKt0us8QExrzbjYf5YIVB
HCFVv1japGAZlRtKHcYlVS7LEnsKsqHN+M/h4zln0ndh9iinb5mwYERI0J/+nPexA3wAbWUGQbt7
yOK8eH6RliBgRDZu1QOoDQDTL7w6PoRfBQwyq9KKwV+hRUioiihh7s0T8D6lMok8Lf0k6KJ645If
obTO26FVmyVFYOABTjDkp7Bn72Sb7/OkaBT8SKyBgPUzbb9BaNg6ZfTbA9YxZT8aSKlR2xEbpxxY
E3Wgp/q3AE/SDBDqGBRdzDpVPsyGUQa0QhaAb3XSVevndCrEZAxA1/xF8uSNW5WicNtEoEhNYI6w
nKtRj7T3zLAeYz0K2Ad/T8+bGJXjJhY9RaB2XQOv3tCCw1XqtUYY98RQaNPRAvhE3mFcr12YNqRA
WTev4uxLNDgHf6UsJ0eq30rDfejEaD0RccPPHuza0ITY5fp9RxykEJVqyiIdq0ACmgWeyEy/7zzE
hkNTgdw/dC0py0LUwgWgGbVjtDgxfjVtg1RXSByMfIq/CRb3EEUcHT/7QVInuDTBb0COzMTrIfqN
zLQ4J4of7WBT6PjN9crFFCaqQ0EHs8Zw8BgjUcXFR5KMvqPtS0MT202Qsm9RjM1ibbfuCwuqq3Jc
fIQEKYyrSU9m0RrBgIecwhicIsTwfKboNY9xVDJXnG5mrneZ4QAlO3ssUais9NDt6hte/bS+GM+y
lJxQzdmT+pyGTX/AGOWq+CGbopqixk47OO2U5FeL0FCXDWj7T4sG4Vmn3uhVqB2z9/8v37gB3eEw
QiEkvN2JHKCtZEs0SRPivgKE24aTkmZ401HgB4E7O2NUYibwxioEYs/2sM2YsMY4t9IUZ3e+qzKb
9RaNdIiRpqiIsJgzj+wY0kGreg8KPlrA2UdTKprR4HAvUfHEQV57fZ/hwKt21sVBTKXt3SuppqHP
eEjyQXFpqN8IUihnpmF2+85G9kW9+QyFKKdehyXtbpOyzhws7arctGEJQE7LmN58RqEndjQRlZD/
nEf07lI+6yRMDNkeGdpcU5kyJvA7XcdWMraZaubUatzL43Aiw0AWIwmIA8Uy1YtH/xxMK6ZNxhAt
vuQd/bk9RGQxt2mRkdGI99t9BrZA4xq3dGbq0wqn3WtrNFnIFo60rxXKYAF//HqbSHv1r2zlEEav
xQ5Q/2ri6w2pSbs+ASnPUjOIYa6Z8kAPEvbCDLEu/+bitRXSHQuMnYHF5l2GRnoS1LY6bdevqcAD
pGFRrpHX+s/5GZIqgrL229W0NwFH4ax8+fn7RbeVDJtfbYROKdfBFM6wNd74EazAdfL6xiOtytnQ
tow/o4KsfHw6Ir0hKO7edswp7z9rLnosxlWNshVB4QdMqE6EUyebdkN8KlaEmg0GEwCP06KAQm8y
OxwMdsY74xkwQlks0plQ/fLCq+F03kI2TSm8UqTO2QRtyIbjXmFBb+6iMYQBZlsDnAweURh2bP+3
0R8ydx0XE5DW9oqdpN4sHBKaX3OmTZJ8+LDQYVhZCGksfuXiWgYSDgZRj8LMyTKFSH6PjRSUD6ac
ZfYzVrkge+TxduCZMRDWwg3WagQHmwV0twxwiq4+Y9jMWkDEqN6A3GCvm9RZST7r8qSfNqcQeqI3
yydvy7jcvTss2lya4kJYOzSy0e1OzZ/vRKZ1q/RCD5UgZpuiPVqTJMscxLbCysXfAdrY0f4+u73G
Ww7jVWlkmtjWSoNgd4Ie7Uu64eFHSe/s4Okz8YwkaLQCf5hucx3i1oV1hTecTrdVLJhEzxP7qWeq
nr3cwE1umg3H79+9ZMin8iBIorJSo04k7CZ/+A8bjLt4ut25LHZ0Z7sOOQk0T6z6EZ5Zzi4J3t51
DsKyLvol0HbBD48HZiekaF/Nn3dmS4VeLr9n4wFhrLt2SVINZi06FYOD/B+Sc7qgYjhIk4rhHKUQ
18FczgnmPmdJeFS6hiiPnASww5c8xrmY1tlc6Q+wekVIk2kz3QQKzVeZUVGEAPxMIQtjnKv+Myje
Bt9mzdGZ+N7vXfDgQB6o4uMvBT0k3Kh9q3UGFx5a/aM8xEokVOhkgCAepw5QA7cC893HehiGNdUf
hPFlpR68CZUT8ubKa/3zcemUeV/26t6BkB7cl+CqzT7lfJJIafL6N7jsNEWz2+zDMdrUL2ShY1wX
qoZkaebxjgRDxsFH8hWG6Yej8iHYrvJg6gDVkYF1GoLaij4eTU0zxMkLsJuOaMJEBAEEPLbp6MaZ
uak/kLPcN0fhO0bxBbFMH8BUv8f3chGttHKNoV4AvcjUQSq5gZ9eBsDWTJNgOIiFXPu3MMXdZZxD
Q4PYkaxXqwWoIs6O8uQrKOydb64Qk4PMyK9bsCLlMWzJRWaH1RwnBvYwTFpfQgIxPD+jrqOxzMk3
rUFFbZ0lWain3LW2SYFqHxILrRxIDdkyckfp9VqcmB6WkJeS/Do66TGNsoJzG3oqb0wqy0A8tOIk
SFZt03ppLOZfm5P2nWz4t0DNVwCHMtBKk6P5A3UF4rV5Jm9YrKTnFArtJ9zC0FjygMWJ8NlbTd7C
JUgNafN0eLE6ujBwr7AN7ksfsOactYodRZWvl165ezC+j43bN5p653Kae6PJ+D2y45qoeh6D7Tse
TzLbBWVJ0qC7xaxJjzRI9MVQqhFQxDmWs7QyN6mLlsG39EBjtZAgDL1nDli0lgzXdN2G9Sd8+wBW
0+9NauWU9IonQ8fq1u7Cz7dgTK5r59KsE2UB2P7lRR9Q6HD6IYeXCG6E8gZuKYbPJ4pUXefM1gCw
nCVNDBpL/WreiCS0GzaQUHxnb21cRjXDgWQr2vKO3/T3UfRFpcvlbYuDaaQgM6HMvGZEk48HCPZG
9i/88OfLDBHr1vYvv2Vz2GyYVw0mucTSZe3DQOOdjwCKXSBNkDTMhsl3N013dhAfODlaLhrrVvOB
cSRFmV0OS1qFrDA/OGMAqJ9jsjyLC+qSow88wHMElUIkvo0HLDhp0RPTNUDJg2f5r/Dbpic4nN7Z
BSj/ZK8VHIF9IZAMM64NJ++499s6Q+O8JCLqGW8lfwjupBjruR3dSyvO7VTXAf6qKYevgq07wkEr
B10cmF2fDggFEKxeNiWJ0Bqd83a7yHMDV1QPjSC9wU+aY5DmT3x8V3eA3v+xXzL8Xd9cpgEXBlX7
vDsElXbMH5m75ladaW1dYL8kG6Akcc3qFOjSGEQWaP21/7Okhd8gsyumV4fKq0u9ovOuE7XcIf8Y
Pb4ksmHA0e5IVNFx6RChu8slLWeQyntTtNYO4fKubvgxxPBADyfwC9VAFOiGqHFyC0Gk/ErYwzvg
DcnftH6le6QTKjWHJdEYvIJCXxKAaGMMqPuo8o/RSvsicgpL23Qjul299zJSqd2xTYNow/VGlbWL
WVYHYLFWXEHGIL5nSgrcujQUc3gIxZ9lo73Q5r9SE2xvtVy6HL5S9s6dne2PaO3K4OWh3XlIjVks
mBcmq5Wy+BwN7ihSCHqjzLivXIo3TTILdEuimMGEMONM098kYn6q8B1mLNvlbzFPF66vuyqkFUnj
d+SWmLssnK/G1pykOPEwiToX6aefuo5dA0OhL5ZrMB8+ci2ZkiZQ6ct0y4taoTgS1/GWJldW5fQm
x9ynrLLkqNWw35gmZbw4Ftydkvk4sr8JoH2D0XGvO56rzndep6N7PdCEITKvxcz23lszw6gmOe8m
UQ+YMq6gRmqGv9C1r1REmtPk/323vptFr8wtfqb2ZO3TwozrR5pPQLedqRkWnesR8gEbkfh83tYE
blIJUeHlS0ST11lE+edGUWtZlqHr8Zp7i6Efiajz/YlOMrYe4W9GQNVhkV3ANaB9tLK9di4oMjvL
BIYjs3WPMnZ7by4r1BcBQwCVIvb/RKfrcl3gNZZyyqlZhYKCHRSNDqKdFhFzwfN+rQ5a2TMx+z8p
/wbTavLgvO+BwF0xa/ZXmdXkrJRztudkpjBUeoFOhfw8kJWpkwwpJs6Wp9hsi3ZsD7R4HKWMaN6k
oSLRynWPgLpJ7O64lFMVr8x2+SlbSZbZ3ne+XHlM7iwdxtqLXYLU7zw+YGciz34aLzJ+BZtHLkbm
qC1F6ZTfht8XM0tlVg+R+4oEhDhgi+/iHWyq5gRDhipMgPblOWBB+YBe7beYogJ1jTUzEvpe84VS
uFq40HEwI86vll5D26jy16wN2S42HYqL8GtnQ+9D6QQY6aaA6jmHBKgyg0PPblxZPlbvh2SVohtB
Csv9gMMv4inoXQ+AUBwfeRHzhY7WKmHJ5VGKadpsmJYXpFGR7LD0dwyTlgU5fSupG2QS+8vg0cdr
SNeKNRpGr3lnqzhiCT7pfCFAfmUUqO4tVF95pLswl9gq2o7HhgOT6j6dZsviT6ifO08xsBy2F717
7Z5iNRKf1+q5doryuSv2afV0/Qf6DCmfAwpq/M09vdyDelDDSpTSDybcgmtH4y35UqvBPnftSowe
YCvVMEbPMwngReI4YmZBqo1X5dViT5WpNr8bYidsp7zDiQdEo4ql8h3gbclFUGc/sUdSRu0XZHkD
F6rhj3m8odC71iyh1Mj6UOROP+rw6B53x9we95RTnXFID7pjX3jgqEy9SxdmTvuKha1ykYOL3arH
g92RRHLiEAw4YFdFm0t5JjGwACI5On8k8/XsHq4Kb4R2o7IdV5kHm8p0HI2bx1at6syNbf5Ma0yh
bnK9SgHKM4J4iP3sjqIbOMzknaQ4r6Fe6R0Eqnbk1U8H3Nl0j7Br8e5Htf9wlREwCzT9ntxevCFV
/pQC2yVovLRwiHDc4Fc7J6qZ0gXGpiWkWuJSITxI/YhsZh0Lv+Xp+tCI2ppVF06DOLlrONoOkloP
9oemL7Wzz0tPotdHszIiY2znCsrGN5zBKq2/ljx98mG6erCk6XTiVFdRNY+/CKJsv7oqmS6eGHAO
XYNlq6fE06rJ/n8cy7Dpybn4V7mpLcUd700vVLrZT2XyOW7otKtk2GO5QWtfADglUS9fltCFB/wC
7lp3lTWNFc3FBTGGxDQazBWFoHp72vM+cJRgwoXKEQg72ByRY6/nh3yrxzHezxxMLkCLqDPkol0i
5XjnptBPhjXC/ViH5Y32xJHJAGcQb/fhD8ITWOJ/o3gUc8h9TIVn0jwfztmIb1FlULY+o/2VE9ak
XJjGi2eRjc98vlxzPpt1mwp9Koldiv+n7wSHAxFFXGCMF7l0BOkDL7PluW5hltEs3leCnQ3C4XDO
vItOVheQKHMJucZX6dBWdgI1eEtaPw3zdKSouq4MOyO3U4HkngqttBBHF8N6mb4J/3Bm43Vw67oP
47XEw5nKJYxDTv7CjbdG0oMA+aFCZX/l5qAhs8Cn+Diq7rqOBS2q1Fq4At5wSIysO0HF45Ue7ujQ
Eo/wIR8896500h9FQaMOnsai3o/Wwz/WxtTXac9G4p3BCct3hQfuHTnIwmoUXLO0/2uYZEDPzx7Z
K/GLeb+1U4/sCsAMxt4H9isosiQUa6c8gNUuYJvRlCmLJKu2Ahz9zFQEWGwiLgPKALADPZKiGI8t
68nuD0wdFTBq4yWyokcfCrzVCk2ojT0wn0xlna34osfjDUHg/GOLMR94SoyFEeCW3wqwt7WbGc9s
9Jl+n0pRnWCah1VZmzmst7rVRlgESbGtf3VOA/M6Mjqq+bF0+KV/7hv/tFzkrOAMRt1mvcFsaAoZ
FHqBGa2tiwR58TckfeQtVQUA9qk+k7xClD8OdfSSfjubc9lGGQNlF9hvWN/rtwBAMACYSpJjzukl
IevcCWRgDolA05N36oeKsv45fx9cmSPKir7d82Gxhz7Xfq1JOvaEQMRPGP5nAyWByAPGPG0asfno
sM0hKZOgR/IkgxJD9yaUqhGFs7jSjPsJXQ0UlJChjJie0RbOWyCGtFaT7fKaC5INplJb3monXE+K
CrJQQG+Tt60AhDCxoCtKczzjR62sg+atNmLbw/2IO58W/obTvlrGVrNG5JKdd3wqfwOwlkxxJ+z1
d2YypErdEVouUChjN5wZApyzp61tw64JMJsMqqFijHVnzpetlRqApNYuL5rlVkxyeP4GeLIcfc3+
/EdhXKvbDoohOgEJmsL0BVm+6tnoWRFylOabePWX26HVG29JC7Oa0c0P0P4t3KxBB1TvM6oKO93N
a30Z6BYqTAiYrok18y6SjgeQpMtqPnxop8YzRmXhPoqDQz2A4npzVJiltFcDcXR/H29hXRaMR4hg
LMrwH45BJJpRXGLJuM2OSR101681odAJ3PjqilGZ5tYs80RuyjQLqd1FY6GeFDDvGPoVAjK3GRQz
7HhBeGovq1oD3KPgW5XlkLqF+HDl/1nzUF+3Cs4PYyzdmZttFlzsaZ3Dt596GdoKmqIru2Dksvmq
gRwOJYkZtHxYh1ofsPDNwdydp7X7OpiqfvpGvvl/J94k79HiIMb+Oh3Orxuq5rTFn3ekDtsKHqtK
92phBHOYLm67vd6HxZ8BxXf90NtkJQzyfdtkmEu7QCNasWzIEV1U6sEQYU6pnKKpA8SARVyISGXi
F4WIAmoUy32vP0Ftg0qmNjRUePGBQMUXj1Fy0KG3G19cdbnEvecbwmIEyVG+MEiyG3h8jQLWKra6
Pi01rczncGmMriHWLL+Om1catqTOjdBe+t6zI+zEIaszQTqM69Ipyhp1jzPdOg83sXToyl8C2M3Y
oUAAOvR5fgw2wwzXrEdJoMUuw/T3tM24FAbksN2lMd3Ju1YT+ZoTqqtanWXsdhtvQKtkRua5w4xG
ST0VVVEtUXBvuSR2YN8IPjMDB0Er2VoaPoPDw9eeaJKWA31wDm2DONxnCq2Txf4s2BHUkivZJ9sQ
iAd2p5WUMEQfw6ZBpZXzv1xCqF2aSSjZV28BeUXIciFdjLa2pzaYwguZMDgk4gw9Ky68GjMnrKiW
Y+pPTH/FapPNn0oiwMjSX5ycZ//TV/X348ekfN6N0MVSvCbaePGkXu+5cJnOU3rfs+/e7b4F/oQn
ET/yYPmlUafbhTfA/ju4n6wiAchXqhZ4bAgrRAVhZmCqSfyaXMB0c8WkCxcAInE5u9+lFPwY01kM
XIAj3p/MU1ZcX+KwDvz7rd2JeY1B2noRLzrBlRLAtJfUJQWsxeFB8ew+3l3xSebhyNGFNRBbJyz0
OC5a/6GEOUXnKdTnQVts2GTBlUJO8kBSYg5k1UUnj3I5GbENbMiu1twPkhsVqYwmmEoflaXrcV0P
QnN6wm4xA+gTk+qrIaoKwwZLT1vM3WMi0/WvRZV1xG5ATvL9TsdtWNbA1eUdL18ZZvf+HU3lMw64
0/rq5nMNXoUiSWtfTSeslJaxiIcnq7/Hd7kFATKo7vX65qyie2va+Luj4Pn0Pa8AHwxmWSkhXPSW
rb5wdf09f4Uf7+g+oHMxsRSG38jcqEmBPG0QQ8RFptmfYm1LEILqzhDZp2uB6ZjIb4c9u40sr0j2
SNpRi3iLtKF8V8p7w+SFyrB0O2+b9auQNrhxDUb8zFcCZocWxYBGlpCUIXrEwXHi2jRZMSKE9jmr
6UGNWvpBrpycwRcYSAxTU0yqT5Rm7t/147yCM6ctmh7kedoRVZMPgf7SebOeME45Sv3VrtzS8rl/
Dqwk/Ci4SFEZ0f8K+MZhaAM3VOPLtEziAZdP1mvOauLaZ3F6ybB/h/8B6H8Ncs49unRZq+wYNd+p
HQetIOUTQ+LyX5a094zRehajivbcXTi5/d/+gnI9PIKxYiI6T+tSL7T+MDW3PMhlgvO0VWes8oij
RdBHPQPqD21I9ES2UqofWtQczwqPj3Kkh6qSW0lRirQ1xJEYFMvE0JVlCOipGtHSjYoiWn75RpKm
fE8eVVEOKgc+yNsmrxWHRRDNg3h373cg22p73Ek1FUeS1itZbzzela5NZQKaR/iZxYHOqfVgUAZ/
jz6ayk3kqLECjl3vZnjbeTkdGEXH4sByJPSTPeS1w/W7VwKqwSN7lKpOPJMNUNXJBuR9RPkcUIrq
avfvFcos69d/oQHFp0EOk3c6HBE8VEvLo3qVqTYoXJjZQY+jEJ5boxy1v6H+PaQ5IJrju/OZ1Rjp
qgxPUpEuXYhaQ5SUfkHVepTN9T6IjNovLZzqWfqLYbI1JtZAcQERR0t3BQWtZOO8gmlhRgzC2V6T
QPE/IyJy4yvdolxYrBmr2sghq5E2r+FM/U1Tq3POUwImGA0dFGCcQCl60fV/hFpntuTCOtmx2qT4
C4nkfloXpwbRsVFaQIRT8FJyzM6G3eCUsj8b1/xYfmh7MinPcq60AZ+8sNHZbNedHTM7+o7Ks1cP
aBitSSqLgfcZecNjJCLeglkHRxkx0OML4t3nXA5lYofMvXZ1stAntqZUsqft41jpVlgjzvxU4aou
x+fFmpDmd8akrO2rGWNmGmm/WNEhyBY5D1Vkj63tkAVAj8zbD0oXDSaqsUeO8G/LSt7x+18AQKB9
OpPNvkC6LuzpCrusy3nJ1Zp5ipR4LiSwA6rfdFCAWpYXiUruytI2WJ+zb2FkXjV43Ec32LVKYAmY
MKRLx+5Kbs3l4LCsh49xAh/V1DR1jye28lBn2QMzLqcEECFzWz9LN86Vw0eq4Pjmxa5jfIBk5w+3
j+CsjxlxsTVs98T+FPtfOw+8Q5YKgYIRhplIYOa1FADzYJcrd7qVRLC3WHKGSnaQTdfJBZ8iomL1
TIDsMlmADVJajVV81152/OkNOnrOCD9hh5REA7/+MuLiC8+wZ6oX7zuyByIgLccviCnOyhHswy+v
Z/EKwyscQT/IrdNdO+tpXbIbm7wW9m1GcSvn5ddTwIuMebtUVh2MBUmywHc+9WvuNDos+l+Tvh+A
Xg2nIXab3yzl+zkLdgRZBCNga9IbCWHtEE96CxPWLOMXXEBZveus4h4m6uN0FEfHywwIn/NjKJ1h
+3Sm2T7HYFJga5IrQy85OHjcMBX8CeSMMjt0C/abVqSAK1rZDobWrPq1x8B8wuxqcxDrUBlMDl8F
dPhXEGSz2mqS43T/PflDViG2TMEo+U/qlPWQ8ggQ3R+OS/c/t+sPRtOULDOWa1UQI/tgK1GzKHSn
QVyeGzvURj0+IVUSlx++cgg+duD4mkEFKWb0xnicyCpV33cV/DXCyALTloJFqaDVGev4nx2NQEfF
CJhwpGx6zoyqUoQ9T00Fb5ob6+goNkn0wrcefWz/zLeY26hlap8TBPfy7yHRCj+XD3qa9DzX0pwb
8QnHzGxnVHnrwCzIDDfhjf7pSgwNh6EQigoZqP9suEqnP/xb1ZP9XKoSoXpWypltO+zoMv2A9/4f
8cH+4XOqFg76pVuErvrT8O4xNKkjipjs11XL8uZN3MAZXgr5CRk8jnCg1ZYVl6f4BU619b5/SsJr
8qe2MdhZ6VNL+bpFPfZWjxZfXp4jg90seFZzNhz+kjpvHzD0NSKlmHBuMVN70bUxf9teocByhzp5
irHguAtPDWkUHkt4aR5Sf98fm+bbo6H3OGfY1kjwZiddzqRjqcoBudAa3U+iCrTKYIQlftpnD1WX
smTGIJwgGXr/nloXeYCX7IG4BGfkR7LJUH6M1aDD8AKmYty1tilQkjSU/nyiXZsliSvSSD+gy33x
UvXz9MIsO+M6zZDhIEf66AKKHE/CKy5bjce1h2rNmXoJcZ0MBHMW508MZl4PnlMQ2/E1hX1f9Gca
iLRbhANqzWy1oyffNYZsJxr/IJaStuegOLMMUtKZeXkv+CV1ZCYYLwlAeeGhMutxnqTv48GkcR8W
AX23Gkv3IcvEVhwCC0brSZz6dDfLgGCxS9KvdcGuZBxT0zslLEqBz5opa2m02KU2Un4x0syIsHYn
/+9Sp74alAgy6TUwC3eu+qfkFY6Xv6tI/Jp+89j/y8S4KFeSjqODOba7F7vCjM0PsJllvO9213tk
1JgVDek9MqhGHtmapkxNFNZJqSRJTD+HJD6GyDcq5L1h2L5s0mcwilRJZ2muD5va0xG70xXTyIfn
I1Xxe37FDNQZAXKWXLoCHN/lrdzSHsdq8iyCKXr9ZgqKkZ9mj4bSdy9F4wbAFFZIwaSA3R6ta/I5
C0mTXPCAxxrCAtwcpqbfjLp6Nj2qMWaeZO3NTB7pMlUJ2EKMMb9VMyuUHSrfUmnbivyc26zEZ3Ce
EXRzDY/buocDUT9souuDLEHGoLEAww0xPS+wLDWcLTaWFb4giGnsfAjSI8N12iWIFQQgAMD1aHSD
U9Dweo9MzRRFTNJeKmII5IP9zTsa/Jrj7TjXmsEbhD/5ID+t4/fflOtXauk8pvE7k3aCukfXlANZ
AIoMK1CXfvjRdcoNxxwy1UakBigov6zGuIMfjvD2A8Pilq5YlJN+BqQG3tTMvFEYJb7Oyww8uK1a
6FyoCufkoHAcAVsZcQCUcZ4/YDt9h+fPKza1dy7WWV1RSfeROwrn6wHBtqPYgkMexqaWlCLvqNPJ
WDwAdOrbY97EeB7b0UdKoXuQyCj8TaD5zmSx4HEwEw1kO80ljNcW4JQi2eek1jn17lRlCyHlGcqT
gF+i2yZtoP6qM7QIUc1nCvpAo51jNFDfDGCOMHuGDwgfZz/taHrelKIYMA2i5oKxJBndcDaGd26Q
At99g8P3GwYD+FUDXTrMPR6GLVJwSYx6CtkO1L+VbfKmMWsFU6MnbX4WRAZLDIoQbsFpGYbtRXWz
0EtzcPvMwcd834TYnAriEJE0VsFoWi+x/33iA4xpZ+yOsexmEjNAOsJtPJ3dQMmSkOMx09u17GQl
snuLRFJ5BMpoMNKc0QIyiLCWdR7hpeuqWJLWP9IipWzspRDdepwPICXG14lsXt+3yfRNIC2I4Ub0
ZKpMojpEyW3jtJnH57bH/ZRcmRcIwxd2yPFqtVJZP+MjqNdUFPTEcclugPqO/R2pHW8xmHDlDVCW
WrLqxvKI4Nb5RaawUzPfOm50KkR6xPozrX5K6V72w9CFkSplDWQwJ0Cu7e3FzwzZPdK8H6N8Dolu
Bn7rWa2Eeh0NnyAM9pHVxllgkWAkqkXsYslwb7eom3BRedwBaGMEfoLztQAyIi/emRtBafYx7+Da
RgyeeE1CjMoWQZk2nEOv2swDpSZZcEW7O7z+4pNULCforXziVSDXf8KeJfOfgdMEX8RInHT/vfnk
brQDC97Wp6AAnND+vMXxEy13GawWwh97JWm8ASxADxHjb7+n5Ql6gVKbMXojC8G5NGMiFWA6pWwT
6qYbt70TOtAYTLmtWnwrT0QQJ9MN3PZCAuEzIA6CuOXpmEEvACknMvkXACtvr8CY+YIc1NiDw+10
0rinUlnjaRTopQL+bR+LdjiR8q/AhFDMK4RgqYxVlRXcHjCILab06VYNh3JWjF+BdSJwe6kRUmI2
1cyuBXOU5oDt10NqNaEYinfPXyydPHPiBDsP3uK7/M5VjH8Qys5jEBEfZz++JMpsi9v8GGmBBsq8
q3YfPzlng4Ge09KhdE5W+5rRVA/jsqT9EjTdQuesk82j+TLvZ4/WsiaYVb0zCp60LSwz7glo6Eic
lB2PE+lsbCgFqQLBovRvfTV48R4Ren82Ccq2up34ZL+em6NU83v8rg2mP4evIjGbWvcOcSGb6Ef+
yoARckzwZd6lnDOZRVNnnhfzpuMOWPfcIo9JvSoRHMDqGnHtUdrbqO9RykQQiXO2cRRvIezmhO/g
wq7uJxeVKQnedqtiO0pK4wnLGpgvWAtX3sSq8gAUemYywu4naHUfkosE/ylkMYWKMY1WaHtrvL70
4ZRnVVMmPUJ8/boIJXMSB+AGr+4OyeHs5oVOwQfw7XiuAuwcw/5qnIlhIcvElMBAO6NhLQUNbuNd
wgfJt3feC2IH/NDr0nkNh86YV6rPDWOVBWayPG2YpSuft6XpKuJ8HErMPvQ9b0lckVOe3zxxiTLK
oMEOwCEFK0akBdDXDm3caWFMnKTzZGMQH24U+t6NG0iPD5NS9uE7lsOlv6r/xb9rVTvYeNVHkfX0
NqoNDpyT4OyCpB/RIZgx/VDJEsI64L5BpfFrk9I83AbJCk7CGZVl6YNOgfYZ3vMSObH8ArFCIFeP
18dLdwiS6eFjEgwSwjVRJvbqlinEDba+21Zfl2eRfYX5AO/krQWZrs+Qz7WeGBFSWbrMpOnZIoQd
+X+YFUlMEKFK70ngD5tcbwFkfwZ39LgrPqfX4zzIarIbUK0J3gSUlDRuZvHW+Ia7Qj2bZ9z91iHZ
GMrg9eG4vXk+QlmyKN6EvQ7AGdXYw3ObgWCpH9cGuWyhK54Ivl8O0KhEUaM55UCtkXZ3tyYJM7YX
aIjq9ml3rSbNUTjJWGFJ30w9xHAJ489XBb2CHXXjb4vlr+K4L53l+vsNpQsdqKYHNIOTBj0IuCp3
XcrrmlhTvqbmKosGtEjTeWxnA3Uixx4qjeqAfnr42cuZhObMfM39BMDnWZMrqfeq5O4m7Zdh8WLf
Oko8uMZ4dbAsmXcqJ1RsEynhEtLSZ7cMM8wPkpm+e7G82eAD5mqf6o1rPPGd/hW+J5rLqJRDbvKF
kR2/36QuzpoPDXgeq9aDh0Lyu30Kk3LzwY7Ph6SMkalGhnKONwKeydcjtt/Vx9d/5Ak11NZ4V5s5
HUEKhgkMk/sfRQPY0yeLncYdbS32FpSzVZamlIiK0A6LV8r5sC983S22YdLpB0I4BcoFZcfMq9OI
xgakmDFdG2dDrETTpmCE31c8ILaWy9lV2U6eJb1AN9ebhdBszqyuaS6IZ+NyIpni9xkifIx6erLw
Uq0MzbscJNtZ6XnsnUmwY4U1rtc2GLlh+kH9AafvWpqX6ZcAr/HqiyBt6godNt4BEEV18FjjAfNn
iIKEPmmOMoimOQw29OhVQgnLLUccJpnbD/fW+pDIdx6HKpyUSkC6wVzxhGmIhEkS6NTOx74+/2XG
PSpscbpNu69cVwcmblIXI1T84PUIUqkK8vii6PbV62DSwN1CbYYxbRwv0K6N3GfcVx9ccBHBSXqp
lnIwZeMXOCT/uOLapYXYoRQkmT+B9UkukLmlNNF4Kz6kwcGmvh9IuloQ8qWZavf9VlnUWfmOThzP
4Lu7c7DiSt4srSeAwqx/BsR9ZwZg0Ov7xLHPDOS+BENSU5utBATIzDTipoN+pXKKJUJj+N9AGp+K
3TEd0rvZuE8+KZFccYSh2hMe/mjIc9ubnE9ATOKsSOnYiEm9fmzJG+RL1oPiq+5U/M8yFb8d5SO2
t67RCPIA0dIoH8qlmq8KmBL32krF1yXXtgvvgcCw5mo48oZQLurweiZE1JT8b5npKKGcE3KdR28g
mrEBxmoc+cJ6hXrONcA6Hkp4ofjnSIZntC3pbcAaChw4b8DKTpBwyIlIaG+wXCLlZhleDiDf1YO5
axQd39hqaTltRFQhqOWrLKUK/WMizox4kdP/n7CTm8fc67iu71XXgO35OvFQSUBTIbLMtoOeaJ8r
d3x/zho04tRo/vXAKaSU8k4TWM7eizS0fhuHkpCa1ef+YkTBkrRoW9h1RM3SNTbmhJePOG0fjvUZ
f28ahu20fMzDggbdfkULDDCY6MwVR3VNhygDgMRXaswc6ArDKJpJTFxJEfz4bMVnbm1mPNaZ0ZCf
0WV/UKPeYQQ+mCkwvgrwWmspXVD+wc3gOq9x8JtnFc04oxNk9Xbc4hXT8LdIiH9kclQtKOORkqIe
eAnMYsBblVsXJACtSdbl2FJeyyf4029O5ZhQAKsEp03PqCIOxmVF+uuWd/+qt4V0JoxCyh8c3ojk
MmKoDz5gIDj0clz+QDjJWwxO2qUM9KBkxGzOwzQvPKCQhckJfQvMmbb8iY5qbKI5Zseief6wANU5
J+zgs5NiI4516qKNn8HfAfMU1eeRPSldu1fpdSpymSyiklWtCqW56G3RzwtjVr+/I+6tPNdz8uOL
pu4Z9Q7LvrgH7bYhhRhFEl1pRS/76dWGOniEJgNZzMGLo9ozpDKbcFJMKJXpAbd/fMhgiZe5e3ET
7B0Kb9BJLsCeSDn4Kh4oHGG0SY8KhZW9Hq5E2nHsUIG5O7TjpFNue0lIMnBeOWuKQvywQeJJopTS
47KuvkIAAF+crWerUA7uJg6qm/+SVjFKFyCsKgYOYj9a51eO5ieIK7cu6GJXK7D/iH4poHK/l03a
+qgh8sREs5StvbJTIs6/XynkC28zHw/Tt3Aj/v+Hb08o8kHYPBUQ952A94kfCAzBIiJ2e6PYgj9V
h/Di1cgABZd4XB3cOgRJotehXMr6QZcJtg8/3zPcQPOOPaakDdQ3lF7czz4NVNNrV9lEWmlEdrin
BkPhc8vkb5s8O2My6rYH2z1WT1tjv+L8294KhY2sspYCYfwedDViH52yAXEw/9bMsrVQTfOX5UfG
9NSXP55dJN50FH7H4YDCt+Jrkl9fKrmZiXCw0Z/RV81MHkH7MkztenPUGYiHpMLSRq7+2MGUYP+Z
TLt20dekiFHw3jokr1RfK15tFdcZZyGvzk3bScYJa6ejf1hvyCZTt4GH7vqwi4N49B3dpR/RgP4u
YI2bQkCd5cfwBx6QEwMvocQ7rIxXkQ5+qXEkPQo/PEDZxjBCuAkKtZ+FM903uG/Q8UavRt3ie5sc
LdX2YyLkeo7zNmTkGcg1vvHFol9HCPGJkVAwWOy+T5dUwCRGjbXWQ7MV8ND5Fx+D48f/TdVI/g3n
LAIopfFIQCX0sTNSGMM62BiedbLINvJQJLbGoL9wiTJnKhCXcQ+XAHJZad+pUueCmwt0i2I/3N0e
7MRPsKZHofjCSCCQc4rvEgqjoOJ95kDFIC5uMWkt88ufdTRTGyBr4y+SqR+cJDBI0rYj3L64CC14
enPqSuSj0iUyofjZrnwXHmF/KoNja71r9u38S+0Pyw0KkOosjdP1esG+76jh6WPtlT5wruQnHbia
9qHrcNtTdKq+jbvM2lAyvW/RlJpj24MGCKqEd7DatUvmswqlg+J/vsLLQTsTxgvjToZbE0bQ6Cny
36fJzPSISpdQikEPuBLMC3sjLLAEgggjegKDJB1iYpqPwUkvcMK74e9EhKwkJiZ0jP+dBn6SbHK8
7TENgGCTqIfDXuGUp4Hgmhe3ctQGbOLLFaHO6haEJtXM4Z4VKhDRIfF4FcjwxmXkazPWFHWDA+2C
JVxhNytTQqm9XV4z6wS5bnyuj47kY3MqvPbNMy7pDfVL8d7O8IeNX6WG6p+zvd+ytYLOnzqtRSzc
Aktf1JC3zqihMc4SCB5NpW/JRV8cwwdGNd02DHPbQswPKvfAbBkKVLAvtLi/WHrbkBKz0wH6Zlp3
eD0Hqh1NAy2Agr/tUtTYIkN9XTmOL38wB07Cw+8pWxcYrPw7K3WPSLFxt2O/NtPWqXv1Y9K1sHsN
3cXQWNjlaMppV2dUK2mk17ZuUIg33VYtvEUsj4sQXZjdgcb4iehZR9IE5PUqcRNoxSSYVrQbwswo
4SaH4TBVuKvRlpYL/7tSxkQ/U+y1QKq52kQD+OWOJcm9/7WztNFz10/LW/v1C71tLrzrBEVilsu0
A2+FnD5t1l4kcsBCYMcTkmniGUWgn0kwn48Qc5w51NI6gTzL8lCkX3mSfVl4bYomfcALUK9omPTJ
Gua89JVmOEftCYNWHhYBLGm5t9ltUIjC5NFLAj6lqVcH3Ucrwfe0gXrkRslt/zJnVtCCP6JpZ4Eo
SoZtN6WpusKUCEOWPN0mY79gfn79LW/zy4SIQXhppMVdI1D9fHzIN1yaIFzn23milE2cD5wRkC4x
TtQkb/il13uYECnczT2EyvTyZ/3gBjzmPbzmtV1/pbpA0XPdCLapR9CGTjWXuSqSVtyt0cnDuwSH
BcDD1T4Mwj3KePGV4G/uo0S1nRwEVjBeX0DLgGbHjHDV1kn0ZyJeEEpQsPzd4hTBy3atQFsvqA+g
0MS+cwj9DhEz0ZhRLI+HY3bKd1hpsYoqAh6ZZ2pPLHqVZMlJWs4wmaVn3C5NKGGbuhC5bR7kjJWj
dwxO2423XCUJbyqv1ta6MCNyaRZI78FSehsy1X3jGiCo138/naetcoBoQrvTJawtg+SK2cuY9uCk
dSN1UPG0PYllPHWGdn/KUa6CEd+UjgEcpjynvLmWTnfb0j3bXidMmSSKpJO0vB8JGmKhkgTMFMQZ
PBZrWD0szvET3GNuxRPRUd7snJYXy1QtbC6SQT0TOjbNe9jJugTxkPbVkbZ/gl6E00LzBsyS4x6/
5NBF7M+RDEl+mkjMspMuVrlIM7FRlFakPOshCy+D63r+dtHzutPcQl2Ye1wRyjDddMDNRovyM521
l/3xSm8fUC1Zrfadea4M5VOQ27vbVWvvjiXcXpy9p4CPgUHOgPX+3aIrCtZ5utEkii6ThiHGO9F7
TrW3o2Nc7kT3f1afl6SpEmRYPBWCcDE8rwlH9wDDoRWtmJyujE4CgYxtWbhPVnlJUJiUx7Id9E/x
HJ2zlatQ6TkpMV3VTlLTBdI99ACt0+nsX0g2qGgNGrNMvdyRZMOThKGHIIMsHvyD1RXVlMIrRuyv
ILH56BH/JaxJac0raL6v2nvI0oKfGpQpCM4sOhjLBb/y9ZEqsgcTj47Ec+FPoIUupf5StISui+7G
6NxQZhKebWgB9VTp2DR/tMOvQeEBYdcXKAmLbFYZbXCMF56WONJ4JUC+qmc+hgSRQJJE1meP8cG8
ghMTLdX9Q1wC+3Jp1IkkDAQgnHyOlB5jt4cFsoR64/F2Tz0FLkhUNWCc11GAt/1S1UKIVxqa3Vj7
+MtBCaUFZykK/WiglnxBOKsHFvE2BIICPxCaFdxo/dd9VewT2acLLo48oN8P5iixsuX0Ou0Ujphg
IlYqIQvXqKEoeMmMmjDLElNjpQDlLMALTwoln0Rh1c79OdBxa+qRAgJE1IW9Ge0IXblaFvn1yMKq
oaWxeL+oZOdyVffAxI81ojG008yenakt4qvZxtRH3cbQwthvNAhTLEbIJAFrYWYWDUkP2efYubQO
/W1HGCwmiN+MseWWAQwc+7vK0uOrxoHSvCxwy1Qi7VpOI1mKe3V/cldfiH+YMHVdMw6sCWfPuL+S
2Vf4R4WFfdYjxNtYTJNLK3v9if04sdWhLDbRqH4mSWO2dotP7JyAaUNrdcxeeHmmlfv1SEZth3rV
dQPScpLTCRfhIdfmLXpNdZdAyRkLhFxECeAI9OerNqaly1CcGm17FsW6xU1X4IAiUPK2h5frogtv
S+DYUAWhXFVzf8PJtCA3u92w9xwl0knMF7h4R81e0yeUA1rRjTL/Djp549yeWKuKO///0PntP1Qo
f/CXx14bZNgNWQOLtkHsJ66RK1Q4Hs9lpFFJib+0Tsy+cLU8lUyFcP4qOHzj24ju7ydzDUuouDCt
bnlOYLwbwWb5lsReqyjDceOWBW/8cslowEKUtiCJ+3UIcmbdhj3JlfqX/I3kS8oCmbBPrNieOVFh
KsREVPOZ8yKkKY37Hq3geojYjWft9jeq2+30ME7m18d8xgEmWckIJe7UELjdurqvX6plOFcq/i8i
NVkxQy/rfuenPW38J8AjtQMBGKOrytwBSSIsse+3yb+eOeyAo+t4JOpEZCoXw9o2/85wIZja+Bqg
re/eAEiwGmT0yvfdnNTYGhRxE42rgbmb5E/tNuivGMoHAVNnfulWnz0MQcwQRFgu6byILQjhId6L
bCx2qFRZRRl0sUtPTUip9WfVDOYsa+59uBlGBluyjOIsomL9oSRznfXq9jr7z3Ext7yFVKgSQ7IJ
KwQ9XEFBCw4SRRnbWajYgslibIsTqZpBzJXhnpxQQ9/zHnxQUxiHIvZBSzSvcmL8Bpu8uczFoNOv
JhPh10gVK0gqsqJHKK/42Xdj2aMEGaX4DOKGDfWkkDJzn87n2J/sBG7NZvGgLoYpbefFZbgwarzU
ufkZxfhc9W8S90yFOdJXn+d3qVvASmeMTTH0MsDiy3qrLHvaHJl9yoqHlPjwg7c7fzpzX+1NSTDS
3nEi3siMZE5/CooJhNUUbxLub/cCMV+DXWuYBjPGlIlLIO3kKIXAAR0tl93EK0Fy7n37+/NSD2S/
dqLnozsH472WF4T/dPNd0kZVer1RL4oAAIGIIaZ8impqKMPubPgLzYlKRi3XrA4/nTa37fO5M5DB
xkM3XL7rQC1lQcD0A2EkwT1K7ZcMXVS0xAops0RQwIueMLu2VqR4thUe/N0FCy2oJL/lplSg8tCS
g62RDj06mpbfSNQhr6zUDx7dd/aNSdM7iFkF1IHGYlVXpEW8OPleJmwOQHkR3UDhEVdHUhYeZT7K
95TYfHJigiluSLrUcad/EYrK1S07DyW82NFdfqc5ksU6SntLhsCo/I563i3piPFJPUSebjtMq8RM
4VhETifDo3Tj0ZgxrNFpa76JuXswIMKbK9e1I6K2/eZgaXjNUK4ZXIiw6ZdZfhlXXi1krqkiByy3
pxvemkEh3it5tOFcEwN81WlBYj8DZYgI9WUTSrSCNBqsT7dFtFtAe5wDI1gTKqZa0KTaJaBrLGjN
m+vlzgCjM+E3IMgabXf/N61MO40ZN/2GoAnsc211XePkGFxfbsSNn10oAKruybFfejQ92sRteKYT
HH9ZDE/SHU9lKiGaX7CNj2kVw5UsVsQ2lVcV2r6C3U4hFcIJLspdrfIJLDtO/aNIrURS4MU7j9QH
G1gCEoqXGRGMqSsJ+QAgk/7pmRFoyEsq8lomviYBLyJj+A6yv5hnti9wYFIsA6mC3+xvoFCcvySp
Pbs71i5VgyO+jPlB3EJRDBgt+rRa5pfTR/IhWrC09HYu9GR8aPjoYB4K0lNyYh3VAvFtrZW1rVtq
TqwwQhooaiSI6Y34BiaEeapjVSQear+yGKQWrk0mChIyNljOX42J/0QvOOTaVxHiXFggo7LbThrp
ac1cdEdyugblEJIDlJiVVzDNXwsKk7pyQ4GhGWxtoZvNbq8nQUlEatUQTklzdc9tOo1ARkX+jwhk
s56LfDukeJI9M92LG7gqh9yzqjVETBkuNdc1kRSpK3AN/6vijYA4HHBsHXneEBYP1rUjh+AKcK1t
rR42XLFnTD2bFEgAvGPLXr2ui+Z/NpvobkEoB86Ot3Fkf/TsoOEzlYIMEw9Av0DWG+2otvIrM6fe
8qndrIJtS/b+IhRdpk9mAEXdEgGgGz8mcdoJH7ZQHYba8ht4IjzqkP8uDJkVqacHs6m4EW7z3F3M
1WX/IQKvzx+2hoMm+i01jU61M3UdcW2Ufkol2DMYQ0Euf8xf+UGMSGTQaY/+0chN7+9RdjiK+Ij2
I79qIhvaNL5P8mzlcyvaB1/L57BkdjbFqrpi6SJYB49Kl2rvOWFR2EiV41i/iC5CeReLZKK+aX0P
wYCRhro8extpx9ZwyQrfxBG/qZLO5Nk9u/IZsQIZC7OLl1IDXyjJXeoNJnMfLji/ztaI6GCqs4aP
VOWeiWP24geKuq8SzodFiAn9gYHD6tx0Kp56cEt+NS00/vJW43Ch/YVeusRy8dZxMuLUEz6bkult
c8JPh5Zo9IJKwTUHacNW8rLIbTKIfyCA4rrxwbEB86HnCb9rItP+xsKo915YrSAuAySOOC+QsTMt
r5hIahLw9uaeGKO3WkIZhmVdL9U826RItwizpAGY+nLhCRrBl4sHvQe/PGFRKDjw2TS1PhaUn2jI
gQqss9hoizPdqYVufROajZdQ33VbzGayiXb5vL9WrZV4RIYVFFr30Qm/mCuW0l0Y4daQ/dx/L9pv
lKDgzgVIwyz5nQeLNR2OfXUBwgRjlD4Ex45Xg9kYESQPj3xBj3sisZwCmVgFm9PayQFFmm9QIvm7
OBRDTLecIqykzM6UquZb9ymSuzTkSpWPSqfOor2PFpnMK0JzPPHzFxK8VTHLQM1kRkqKpUo5eDGU
QXTIzDB5+/nvW9/ClKwaH1U/UUSMdEceN/5YBf67Hg0DmUTOpbp+n5uy0UI4hoWVF7w0WabJQWMl
rCjs6Ed8RdDHI/JuCMnEb6upHuXFqH6dvDQx060FM84/keo7Ildwp9EHufM8o1qmsE0Ckv8tJYdT
/Q1T0fM2d04jixKsasa7WGRtYq8nQtPcApwtpke38Sz5TWOnlRV1dRuUAIIlM8KPQNFMrzTgO/Es
RNo005fvqAJEtmLhb/6MYAWwKfwOjIpF/HaJtDJdpLbEMQLep8qIeDTMSOYfq8YjipaZOarawhs+
loGgIIGDmPdw6TkVptrmoKscJPyjynIM5ewoH4oYrFqlUW0kXSF1jIPM8z9gvSUk+Vxv5dMxisvS
B+h+9U/GcziwPUoWwfki7+ubUd0W1PaMkOy0WnSf35OomK52nvPo7ZhgI6PzY0GAKfA27zlb8McB
sBn3J+h+exiU6r10LVI0EccYmUm74KwrEMvKAaQDPttLPf3iCt1vN76AmMUz9RFVe0iMQNPYypSu
6uJ1Ewl4gwhCsTo6XCn/HUYrTiQ9ccljknwfs2Iqiesx/M64PEFxmD7pKqR9TRIbj95i9C25KGM1
PERLfbaxIfrT2j4gFHc0w0/P+tNakKnZZiWOmKRbZgUQEq9EBg7MCjkVihMudMLXAzNJV1AS+kwX
MNbtwaZ9OLybtK4dHug95JdwdoWV/6k8FPYET2Y5muuFSZEOLV5lPiZYIHKHG280fjxpPW18BXy+
TkU2vHjLHfK2VagMpulgjpnNmfCKRinLIFX9yqPOi6OXOMoU/JM2jnzUMw67vnHvtJsYYZxgCNB+
QfxdJOFnQRNRclkaonR9j9KT6+4zqRRlRO0TqH/JoKcdmzMfD26L2psfbeokRpmVyPLhLUnFSy9G
ruwoxL0NZWh06PBm5HxlPyyUYBqm4RNdW3zCogf9xrm2XoLN+a3MPP3Qembp4+7n/jhthiPI8g1D
mFZj0joDR90eUbMhbOPCgIEZbrU7m3MNYwSbdj18pZ6AFhbERTK99rF4taHvnxflATGgh+rpO1hU
pX9hXt/dbJQsZGwmXkB3GQEV40iTyXDeU+3bpYp7OPL01NP988nlxWUNvWTNWzHqUQsFOQD65648
WpyW6obmJu8dFrYti216mwkpwVhKtt6dbfP2o7JddeZDTWIpNWJ2Npk/7LzbP45lRLq16NYOuO4Y
38sRQduPoNgDO+ughiiGA5ZRXJ37ve6DQBUymwWTqicRbeuv5O2Pu4G/b+q0bsCSNWrhF63Yee3x
moe2nEgbwIZyPvws7J6KsgghVXQL4uBuRcto49G6V1CaVxYiJ+9YALnFe0XCi6Jl1fgTCfZzQtjq
h0VoYgt1qIdqV0dd5N6LPpMmABrAyyFO82gGBzqFcGuh4HfM8i8ExkCoJYyBLAHdlApGeXpedwxh
2Ykml6T6D02beFWs0qruGDUPEO3qZwnUdBTq16QuX3cmH9zZ4hGQ9TGL+iEC1EHu/FZ1Y66+C5An
GkMXVxkLD0MfVh8YHCKLra/pt0wY4xEsp1TrsAuFQJnFXwoWFe7ou8DDMdydcKqlZut8ezHoCIbb
22X3eFFHpUufasYj8NYkosjV2TQoMU5EeYwB8lWFsZUUOgFXbR6+61VnJF7Y3yx3ejNeM7O9GVt/
/ZT7jzzyPq91BHiTzaPNKrdLbaS+5Cf6VdSO5TPb+6ifPSn396rIs5/mHghVdOuUb1HNWI1rdY+k
hSOhIuoD33g1fz3tpyFF5ft1prIzFTqC/DJuTtQR0WfrLvTagt+sFOn/su8Wg4iYjGmURlYmqV6J
Hp/tDMwVSw/tP47J75twjfX3iFVHYe3ukvYZ2m1AvlCfIhLnD4YJ5ACV20weSOLZXNe9T9LafMZK
jTy6Htsv8qCVAd/RMK55ocZKv8Wm8Vic8/sNeGD3IZjuPA/wMIaz6IGj+kQZ/oH6fVaGmyjRxjsQ
e1D1vq1fGi9VeMODUFLdktds1fXOBq7UaRKdmbkeVBpSeL4NUjG0Pwbn/+NtxUOmlqx6EfV9h6a9
eUmM789MrOsDFcVTKB/yGQjzLp2PAPH1JWBD5i6dhWLYuhU3V2VXkU18eQLatNzrRF5lB/aUJSX/
ejq2EGCvm22Y5cpe2dYqxiuEsayXoTpWFldtqTN4pXO/kfgg+VdNBT633XDOCbBMk3AmD12uPIBR
gemkG8fwji7M7EXPfAxP7EeaQ2QnQxsJq+s4QtUHNsoFQPDIqiY49eBg737zlM9eNXYKtXcJsMV8
MtjFw1LtPoq/GN7itY2Khei9kx2OtbVrucD0dZ4150FsUcNc+9KeilmjNAxxCcUDnDSqs/R/x/3Y
sUvkKDJA21OWF/EiJCzuCeRPhyKybDz1AkdmedezQZjYBJz09sxdC1UmoPHO57veYWMNdf8keytr
GsmTNoHxnToUHVxV8ppR9y8nG2tvb2dJqlkQFKQbogE/EKUn1+JEilkcGDEdr8UYPnP2Zr3jdVH5
QmjzLEw4iGF6RIvBp0pIeZCPB/YfcpSbLqghRSGe6PmCynVzwF7/BN7FsdtattyG4iDb9vxjT0HO
HSbHEavfuxGd+CH8M9JTl7Gw92C3ZtmDOyN9b4zHSGtNE1CK/MnkLHZgD3QkWnENd9T7V9Bkr/lf
3s+e9PkJU97dHTrQTfidA4PtbYVJicuB4HCC6ZnR45ypdYxJGKME17wKZdPQGs/p3XJ114kOXk2I
Dx8CMcekjtq7H9Fiy7wxetAUKj1jKdfYD5bPv0b430q7ghrwdMP+Qpe/p7tv2WTeII1ZnF2wCbon
3rOJQJI7hLj0sGeVb6Hy8uizjNFeCyi3mCi5Lmpln+cT5pJ+2wq0QSWtygl4gvAekFU/pEJHYm5g
Xq/m8qoemkfnuzhoC4JjdhhWUuhveL4zeO+/CVps1Q2/vexWl/DVin4RMNbVjOAOuYtNI46kvfC/
NfboQNMuXUzwJ8EFpdb+akxRl14Eb+d2MnIe29rHvKuZcWROLzWY+y146ZWznzhhxpcPbrCCHoWm
DynDlPz0swfRoWeInbC5qm7FBCv6oM4JCqGk5twjb60q54JzrwqxUVm6XQIcJOsAMyVV8NBQfAMd
SdPWWvzXxSnoqx2wfZwYEg8WPGgvaFZ0zMIwhKTvNMLanohqZw7XO9sEdrqVN4Pn5XYn7Qi71J/P
j+Qc10qpjJHv1LaxTN7H3gaCQ38ge36fYH9oyAHS4ChYZH/Y5N/ZPfiIniBXP5moFp7LTajR7h7b
p+wPuPAc1K8uG0WMi+wxrhY6GCCPoiYJFIr9dQNuDKK6O5r4CfNx6+Fchd3ZNHBu+A1kCiODLtv/
ZbJt6KdZibVnanH9A11RCi5czCYjehzbw+Jpy6BI7nbWeo5DVU2NJ9QQense3SE6yI3E+71XnvOn
3C0/UHN6e60f6gSZuGqlmfYdvOjO+mkK7NaROeBjaKCA/bvl5c0yvb3Z5NIPIrIsfqNvLguUfFK4
ednPCr/PxbpUSpld4augFmdKrh1j1i+EbE6yA+FlHgrumoU7XQQgtBxY9vlVfPBe5lIAqRrPtGx1
1JqVxKRgNk4UhKMhWRmwJbBSjGXfvP7W7yfLvtlsp+6wwMysjczVdHcRgLnm/c7R2wdXaEoLiSdA
4HjSI/jfCqgwCcSJAh88JOKl9iHg6Pf0uaLuD1dVg0a0Dsh41a9/GImAu9UqkaeoPh8jjZx+r28W
2m4unsqVnDR5sMRw30B0h+XUOJMeK+KVxu4g6Ky6XVjAaHiMoLE73w7ryVUO16VzfpNrWB3q3V5p
zsICsFTxhxiX34nXA5oLk2MlxRSvziQE7jXprA1J2MK8XXIYyqHcQUANJaotFsr1VomWGaWIvedg
A8khXNFmfqMpy5c7+XZChYV5n14XCvjQZRlNFJkcITBcJF7oQO9hqPPJomyX2YUkqenPo5Z1/Idg
dlgUAWewK+0yMhUiZ6RAxrng8PcubDMIksNocteTaT8P/bT949q/C0dPuC4R/ncOmSohZKtdxA9u
NeVz/8lRDN7BsXk75ZgbmMBdvDs9qYYcxDjedurolYo08vzBXJ27OYWW+ZNAnZr5kWDX/n7+ZVe2
WxqyOLHqxfp9tJcaKN1jbS25ObqC7YHTj4CDAC/6hSwuPmXEc3Go8EmVkHgE3unoPyouViUqDvBH
P9ovBHwkGdaN+UvJyiUiB++mvHUpL2dFLW8/rJqdSsDKSBEVhcbjlYQJnx4bFTxELKHn5X4EzjZP
liZ8FIjCT1hqLAz2TzqXb/p/U01qxMtBC7wPH/aFPSWo5ROTIeuee+MpvfZEXdLuMDpklKROwDXT
CZCGXYk70VLJzTXSJai5jCp6r/0A3+J6cML19pomLMpfFqnB8OUczeTa4WOopb4cXmJc116Bk+Ke
J7vodMYkYqoIMEe808k0Z3K8L/nOtisW0PHZn/LAPsxElpl/PxsJSAjS7cqX5ONu2s4q6fFluoNC
OfuKboCQSY/PuXq9MKlxU2XrSgxr8EdV3KW/No7ocxFHTBygEzrFMKHDbKEBuo+IxTO7zJFcIDm+
ijVI2agPhgMrWcmUUj0Lh88OIslzTDlmAWOimPwgLwSlsgQgZZi7ufvmyciD+dOphh9j9Sws9hKO
J00eFMRwt1a6+qOJI7HKY0oSjy1yycsTXg8eTiVPlr26wKW7vA11CtNSBW+7JrDs5iNQQPaA1IcZ
I6PJvGJc/bbZS7lrGdT8bN0uTXENsyjAbGW1pqB95KPyenqFhjpzgdfoIeqdCIulNutOoCsPk9kN
LJ3cxGLCHxcfjBLpkLqDy85DdhNK3+rUdo/QMMZWk05JOuOUo/J4ePaHgFuLCe3lBqiQhWv2AGkK
gf4yjxxJvnUhqWSofG0iBo8psoUKI9rhYgoqUd4vq2YUbJ1cxEX/IhCquPIjHG06jrgWM0jfptFw
O5SvUCj0J9/emJzPPdBNdVHJjPq2eRlJRWK3xldhE5RX1qGI12jgIMm2g9rBniOMqyL+DticVuEk
QdU08u7EXqN2bDpmuZjG+oioLXC63zt1dH+8vsYFHHYm4g7sJrptAziSet8QFc8HRAAn4Yt3eOBX
IM5Ee4ZkiLOVgQRferQzWotKG73VmIVcd1zPxbByAfJdSGTrVtaqRyEbMDtR92JLoGqKNbnI/nvf
hNO73mvt15N+DqYzMpT5dE7WwDqyq/KtgSxx04/zhYhpUzA8akPhUJeGwZYEh88PIW6j7GFCjHLp
HDlbKOr93HYsj+ee9L9eG9W6txh2r4UzfwPdC7gnDAirxj2AINts/Ce7Fx+shDYq0wnyrFemdTaF
Y6vOqjSt96YoRqhZOsYgz2Ufon9nuD1ihaD6ElbJynXf1F8P/2rN6vJ5d/YTR3xESK59Wu5RAl0B
sxYbjzeCgJdO0O3gnm56TOYOyqz78rjO5Ehk/cCAr6R8ArXa9vcqJG4XfiBs84nsYv9HdJls4C0m
mg1dpuHfT1KPD2+LlGk9/W/QOiIdi3UJ4DibQRynfbddgY0rmVvUYqRfmDbdcFvIrTzB4haUOMyI
pYv77uoXM49jrFj5kFQlQgzClneeQxwCe8tqK8mMQVt5q8U63YuwqiM8ZAYG0qOIWfTkGDMijC/z
Uv15vk0WfFsxgWAClFtu0XfUqJHEtsmvZeOvPCHL+NHzBwr+2FaJN6GpVX7064t+B6fiZvGmSSD8
eSdGRfRs49/RrJW5RRVuhIgyE4PWTfCKty2AvIGZFPy39HQFlZRDlDKWYJcpG0jjpTUlMfMArG9e
jqUeRM0hVjW/mnlcT27R1FUhapMa+dNYZfyHWubDYTsrt1yyRqb2uNMGESIylgKnGSq9tDIgUVQZ
qOdkqQkqcics1b4IQsxew0tE+Z1+UjO1xcbV01xibZtH11KyVB9hdBM4M7IRaATNSE4zbtZq8RIe
+IwcyvH1HqHnZS2JhDERW+sYT9hoi8DexvGUF5WBcT5SsyL8mGAZbcb3lNUF/Ueeq8Il8HVOEidP
q80XNHd0zKowV/mQ/2rbBJxZ820CVINAjSoWMTCNThwk1ipQLS6DlLf2DgNtrFruBrxj8UBKUBnt
j880wWKnOcoBZ1m0GcgGLYeMcniuDj8CKB5recLV1ScRVIYo4l16srkjmdp6mQRdERm68jt8YT6L
gy6QN7tiz77e859/aw9kEAbZtx0svF59wR/rRtGYPZ9hlkvmsoBpsJ+d9F3MO25g4Gwcoat4wTEv
zsRUW+8a/LvGoJUCG0SNiUeatsUwDhLq1HQK3jTOpxXacS2Qsv5e4DcH+MbGSGDbrU30zHD6VNnj
kS65XNmeE7ZcaFsVxE1BHzQlmHOQLR/P8JAz5cpymJ9+xtY53WpPkiW4a4ZkRkTgYVD4PSa5yPJ7
OsDqtRdT2CoOxoC2ZVVOhLC5jhXSwVkruBZsN7v3Kl/LHWV+4h0LkWbvhkBrA25Dj7R2RTkX7van
x/X0RTTnzKf/ez0yDGBh/NUHBXe8QGR42fE/BRkkkD2itpsCnIS4S7li5ZyL1mH3aKjncd0x7BcI
Lxd7h5M6vtUJEruqKbWqsS+wQplgFEXNnfjJ6aywBgJPtu444G0oiq8hFID0P/cDMSXcPeqTLy48
tPez62//qxWWX/DlwTX9IlAJI5bSuh+O7vvBSYc2vm7d1h7grV2PcFX1XEFvKtjtt+xLqDURE1TV
ylMxsomYo6vx/86eaC+z2rf0HMx2gblMSaj9qESxlwlQjTuMWb1o/0lp8xYAB1s25TKqHKUr5Xs+
6jQEgPHFLaBe9lqJ6ihaBYGPaj440d04475prqH4/QwuZbm8wQxc+jBm5S4KCQr0A0oF1PG1+a7Y
okGk68EG8NVnMMQsb/J9uh2BOXZLlW5xAZJfpoWqzKtxQwPgmLAcQ+oOzrcJdFczTTwOgi4i/t+k
WzsIzfzPUENsNETN3u7fmM7MJJaXVZ8iQXZqRoWivbR2yWHh1UAQHxcQLu4B8DlVI+dN3y4T6Vm3
vLGgkeud/w2XS8SyiFnE2qX33yuAzBV36qnQsaUU5hguYp3td2y8cjVvYmQ+o8wZ3Lb9EqHig0fJ
mKmFp0DrIbjboRPurTGNCnkGAb1CVAZqZcxs8PfDzT9SRpOCTR03/aEqYikus9vyvQ/nWxSvACrF
p29t89DEz2oC7/PorwJztV/6+zuwYEBOrhQJGEiT8+7V7NqenEzcRPVy32iKriTqg8SV3ULi5bi0
2LmWiIx/QJ/zcgjDYVjKH4Ggnm2TzKNVb1HLtW+lwDI02aKtOKqBIiWVbIMw6KotKs0JvTcTzNS3
Ec6Vv0tkA9oO1hj7KF/qE0XQUvualkn2euRhCg/xaOUbkmXr54Azj0lLWdGscG+6f7cjVQq/xoL9
tkFCn8ffeBgPFThfvf7K8dPkwX8JcqTURIqO2bj4ZZQa3HuMlx/K2n4zGJoet0bzYZ87azXEiOvM
tWWKDV9gPBKcByuIhQI9n7R4tgt7ORE58S09EOmcStimaY9f96fqs4I0jNJFS9CQLffmFOta6bFK
JFZSbFkW2lgLwwAdqRrxU8M8/VujZ1KLmuAyFTPtTLCYavefbv/PXMyDrcULw2jaUomIX0NGOkc2
5VErXnugEQ/Uq9jXnkJQMeQGmnljm9hEpa87GHv6yKzrPYk9jkBhyU8NlI+hho1Xir1uNXyDW1fp
RJw1yTOHRNG81+Gv5HxwVpDdD4Is0FT2HSj5pVAxmNNHK3mgaRTylgkaNbU1gBd6AGCbd7b0ucBC
jI32jIsUfCm26/aq6ezjmi+G2GVKRUKqyErpa5+7uAoclKzBgyzUPTg6JO8pSWsS+VgzGiLa7HJU
r/2TOxJSp0P6Q0zlcz41ixsxTRFZNK/OwZPyDOHd1xyRzhEUA6s+5nF35VVzsT51zjB3XicgeqJV
jImc92hiXgzHBzLGXA2TBB8HQpILx1k7uHcHl4tLX5Do05OiPkv4D7WPZ5ot4VpAF/yNEMBLq01f
+tPDt3LCsyAIxFs/+h8zkfLVbgSPtmLdk7XHOuVfPeS09eUPib6LkY9tvBDEW1pGXrqRD0Amll/s
tMA325j8WYsdqe8Z79Im4nOxlDlfqJGrF+6cRKt1btoHEqaNFpTFTUFbUGX1nirJNJYxTjatK15b
xEdP+KUIhxxPTJWLM+14SQdYFuzkBv0M9N1UbwNSBxjXXEwlZGTyiwH+h96MUkKlSud/L4IFuHFD
EP236KE5F0sOBsDOwRZhpMxFjxzPxx7QN+PZOiqBcfTPP6OYCLZLZyHGfX/Kut+fhQXMBNr5QRzh
QaVjaaIDkvo0QFIWBnXtZ1201udMwbtv4OiRXzrMvKtNlszhO98wIbJsQwYA14ThMIs7nnPXgsDI
X6RffHp6GvohI+QMJLjpww++auuZHTUBp7VUd0wYOxFGHPBLw4f2s+5KIrUVViwvM/IW6LMh5ruq
eML9lRoiOF+StTzcJxORYF6mdYWd2Y0wtj5YU4Kq71CDWr0MQBvORnUGMy87WAiKgOF/N+8ONGWs
sH02SvtxUomQzWlwCc55pMemdcNE5zuScXceZScDK7Jkpx0hm+7VhiH6BMpkzk9w2/GB8+Z/F98J
9hIEUG6ROTTkDb4f55dUdAfpjT59R7LMhUL1D5GUGmxpuuInm9Iqm36dK/opR8n4SH+5VprDPvXq
CkAqd8lVZQ77Qjsd9ViCSv8p93KpdbN7QaWlopZngp1v9QPWoRr3eF0m3iM+Qx54J0RZKeCtcOTg
CV5ydR4r1nIejgJb8pgYKEZWcMMvTURcnI2Ko77VlNF+7qKA1369vvE+cHTdtc37dqFB5YCwlB+p
rO4tZ7NNE99uSnJ6anak4tyMeUtOTIePtn2oUOmTMHF9PJVDvkn19Js4r35s5cSQBTcFo1de2kyw
EvYet/btX/J7ERkquWaF1qNPFkQs8G9M0R1I4FNV6DIfUSP+EDVTMmlKYsIia39kbbxBEDeyWgTj
g6XLbr4ZeTtX353USyrgGY9038znP/0ZrZVttCSx+9vP+0zA4smVkBeJiDgJcThSulbj1vnIP39L
ESfb2kqx5E/45zIJGHEgdmO1n/IXY4yyl9amMxhX7JC9yp1F4W1H0/jrlqPsj6RhdWCRPcOE4r7N
F8anJYTyju4A6K3aFrFVdfiY5OQBbJ63e75Q5eFqi/HxopUfR5EPjM8MCcXLJjNvizy0NOmNZhAs
L8LCLe+RTXFJGItUf9jimcbkORnzcsVWX7f7fPA6hv6EB1PXkOhhpu4ION0x978rNIGUS+MgATuB
eRdmoNVxa9sU6LTkLC3+e0AbpxYgJNFslQKeXhL/KVEkmnqK38M77mhVuK3hDuYas7qkbUPwz6ws
bMxPcvqyinz6ZLYE342GdwFt+I8pTDb7f1ZGBHzjqqDg9v1tL3SRuK2QYBdHXz6gZ2vaBEr/IIwy
Cc0+EZWoko361FY8GztG0L28CZhIDmgI++r7onNXh3zbPpnb8xlVBQszNlWU6DFLpszYDhrj8cC0
WpXjzIq3GZYT43wqN3ts34lSLoGCyfdYxFUAysT+nJdK3YPK6pj7qMoMv9sHbByHCm7m4FSQ71HN
WRHPQ9u5tGESWPPv39e9Nu18fsJa+8Gn6TLNV1ybjJuSek0bRUhZby7eUgq/vo4Fhpx8mpq+Q1AS
m/NHmGqosoIC9+EbG575WLbwRkTx5G85fQCSAfRxJxzSwad/EK++ls3SirzKmLH0zk4q+z2kOqrR
26HGH/JIWZ/0rNGR+LLITc+b8hcO2LOzp991EQ6o8UUO0u38p8+g/UzyJX/USeuKULdejhxq74K7
Y+/Zu2oW444Oq0ub1u+dv0ubTyUZZiHVeSFmt4DuNFOWVt0JHPnpjgEnrbIXrJC37kwTN1Zjaehq
m/JVwV9xyKJhEPtCPKxn55Vxur7N1BpeF1N+1a9bFdcwJw1GKs1mYukwFT8Z2auyz5+6+2YXfocK
VlG8EaExzsWaXW0m9e/0oRF6jIsCTPybk0TiB/NBk4HVzZmnVjCP5/chwwbfH3cLoPowTEoBsmHB
Hz4ulBb6VZRPHipVRkTbckVuHb6eBRD5XsRYzO4G/oBhukSFoYRDolmpSwh94iARXsDzJ9DxfvIL
FnnsCtCq5gaZMZTWct51dKYaL/c297iibQRiPmA5I+YcCI1BmaXamY0kx2cxC4o4gszEZz4yDivZ
UdKM7BUdS5MZc4ZcnIOuiCbZkcjGnEBcRF0PglUm430sLnCWd1D9XliTtWvhd/RYo4lgCYgxz2SH
fGBa7+soJe/kk93FOFH2pgriP4gnb731TT4NUUlvlkjOsFyunulnB2Jk63wAyyuonoQRgKNo94Uh
pLibkMR6roW3qiitwvJlFYin18Cp0IxEWjiOmWaUSfb7jkoMaUkgkQ7QfQcBA7ZVtbENvYdS4fqr
0eSYYU9vQYlBHllctRyTBQoNT/gibNNat+NP4Wd7cKTYTYc7GKsJJLN4+94N5tColE9nT1Jy83/S
ikAD8RGS06T6lZe6fnBTd45Cd5Vg30NSzxpJ6oJcqmdGH2HACXIjZK1paPCZ4A48u7JBBBKgsGCp
1VvHY+PD/Z+WobX66wVl5sx9c+3vEw5Qf3oMn4PyCFgwBjz5idsN0jWb5/5htg80caWBELVB/yTz
lESJ060IdraqQ+eWvR87kcF3Id9RzMEowiYEJciykWURNsDb6erhLUP0tVaOnG/TdwA8lqjnSxL/
XUc44a7QEk104ohqj14OOAFTL0xKSITs8WPmwzuhoWe6WU1Uprqp5kI+wAyZRjLvNehEfI7FqT4y
FXxAiidSNWckEsi+nArOmK4au6mTfdSquasZFYgPKkmI/FR4xNyvRNXo6n7tlwJBvKnLIdeLrvzz
+zGPtNCdb7QgT5Bj3QbpGh6dBBzyz3fxBX5/jLtCOT/BZuylE20uaXufptjCYMXDQgaAof4FBi4L
8iLtJYW/4rPTa1GwMTWeO5hqcxiU/ASNgUPo9vfljtSCQvnObziYiXmntBj3Wc1hH+VgwM/sYBxk
MJsQoQo8B89HIPyuA19VZkLGTk2nt9gDE9/UexmuqRmQwan0Ofq9v0YV78UnQ7NzNclxkbFddAXF
L21ziyRIW8W6OyntHmdR975oQe8ZlnoVXg86edOIC8g8vWhAalRYDMgvwrTOSvT93kFmR0LLwjg/
qjyszmfdjCnyiq5JH28gXuotuZG/LL4L3Li2c6sJlJbZKL1h+syYbCCi2Y3WCoWhZ4xawnc3WiJC
8hMb5oywqo6T4VHvcLccXOC50Ts69sM6AI/4D5TF7WyPvVmPWmGyRT1xuSqWFv0aFEbBk/L4XtgM
RKKpMVjNhUeHuS1YQQGjwSyYevmoaVpgbSY6pf/QDYQZrIKIwV2EqODDINVo2PAZ/Io+e9BG31nE
Z99qFgCAGWSMahxcuW1ObhjK1C2vavqQOsqO6+j0eVG8Y+REBKeRBoR4ZRgRdt7rDHPPakt6YO1G
jskaMRBwU643OVFIj88h+SYHgRWSlGJ1Rq0SmP8hGNqoUOnxK2nP+7jzsZiaff/8nQlzopxBG54f
iyFejlQxeGau1x9++XpgD46p4RvW6792+KBkDKdX/PcfFdwbg0yItDYStbtOTVeLkepK5eblW25R
0Ecak0I+uCjyJ9i1x4rlOjb2UX31rYX7MNfWWl1ZvcgQ+j/wDd5S0xvOn+9vt8TREaFaM8pfLd2l
YZQz+kwBYUR35R2eYcTNiM3fO3qScuMbEdQ8IhVOclWuKDebBUsnIxA4YTz2kbygizVezJGpl76m
wIh780XDUvfQKrBDcCIj1Ab/5w0Sa6ekXHf2Ntt7xWIxpPLlmxgIIANf+hgxuH73bJytab/t6FlV
SbK6UATLaDjlbP7Lr77lAKK1Lot3LL19C6FZzrWh4rv/RwgW+LkM9Xytob/bMaAAejYFDGWb7+7N
4g1BIA8wm9PzHtfH53QnQT2Ot8/xHlqRVZoAsd0eHzeiKFMu7eqxmGb9CAULuwP5dDXSR2gzRN9a
/HVZvXbtNf5qB0AeAQUD/NMx6vDOhX5d+FuWcQlqbJXsQ5YmGq5Xpr+sLa/epeXh3xZngxECqZW7
S0uE5PXsz3XtOFMQpx80RyMMAnHHDdrLwzcLtt/J4TbXeJetEweA2V8AO1Lp9VSjgfniMCCBQBek
wBXBWNpV9CCy84W/2a7VSHYZrQ6QnrkCYUhilaQYIL3U3Yilp3qXY9aTRAcFcutxcSaDqv5Hkwzv
Vx3HFCbNkxzDeS295ctcMV+Wa6/DPn1AUholRj9nE2K/skmyYsjrJEjWF7SnA5q9oKlBSy7nL0e6
Qp03XFNCRuTY4Yj4pu9x/EEO9z9a4Emm4PGmWiJCyEoXd+FkTmiU79Imcnew8ujCCYBcj1JLqqjA
utJ92aJvb4JMOHpaVxfCVzfKP0tz6wYWHpn5GkFwoZpTJQN2JhaJ7BID8Nb/zjAZV51xvkg49Z0g
7hA3fIXrRpAZveXFROb0ACLYLQGZBd7qiqXvlcU+g8O7oOumw568DSlGtzQqbx73fEbeJd8sYWB5
44MCC4Bb7Rli4gBQ08tV5rGwZT1VTL54zZSpwn6Qi11KZ4ulHO7+jHeuu2l+WEkNTYuQn/wCksVH
Y0IMUhojXvlsismvd0UXms0t0fpSvnyddcGAU9YRSsVrMGoaeLBfeBw2JmAsLxZl6fWtCMwAmX5I
br/+z93RnNWCbVHD68H6tyF3/382xKxZEFcSpJzdhTiycqaEigno+3071QA8+p1r5Cn7wQWbbt5g
dQos7Ikh/VqooEdRszQb4HTI9q1AaTkYaSM3VNVE/+ZIXrUAiofgCNgDmGA+l8wggMJXNh7GIM6o
nda31YJjlg4vRLZkFLFvNI8l42mzrES9FJtwkpU505DkzsBtSgfg0Swa3HU3LvaNyEi0z3TFMtvT
PaekI9FdXVEhJwdvToRAP0fZ6CCignKGhxywW23kFO4d72J7yRqSqdrdYrmqI8XsT3bZLy8QqGQI
qBbHtQTs/lbT4GOz2NNCSb6VWGlX5D5bteD8M/DKF1OwNpATCGiD2j1k2RYvLgKWOUaU1wnAJRI9
Umpqm/UmIDYX6Xm6bqhur6UW3S16hcbVg6zKc8D6cwCQxDXOAn/Nb0rrbun/zK1WRmGqnKbmZ49L
dpdMtoiRZRjkcjqAOCDoNko5/fZrtLhPJZnPlKXLlo0uDWto/+vEN6Xmr14i9GDOHCu6ZWNmGZwo
Pl6Ureh9iRLCiGSMbOQYVZlok4WH0FR8WHySA/ZZ6HKaDm1e4dxXxxMA1qdeq+GZLYJLrJ3LWGKY
ksrDBHLAbmjnr1AUder2VrMDkQt9WgHTCJ4nDG/oKtu8sq7qQeS3qJQtUnCSNyVdym9gGGA2gZ8v
uQSX4SH//lvFdUkjLSE1IeOHuerUh3zl9TcIlRWZY9wUFSGCNtwdvYdHSsRo8jJb5KlfQ8p/iFWq
Mr6icUpreXzRzFdUsOe9ZmLGZvc2N1nRIlTlISP+0GS3Rg2eVUZFrd25KKdI7aeg7wE8PO7bntPC
oxqlXy9MhAVAWBuOjMwO2sQneXax4HrspqV9yDivcgtMU2RBWEqHHMBYuyDVX4kIOtO1xsBeYKIx
BIY9p1M2c1kkIHFDQiIrpzfZzuYk2prGylmu/XTEtkSjCcb7FUp/w/v1uLTqQ/ydHyM3Ne/7EpCY
4YOEtVXadni5yiUontbX8jUwn3EGe0qm6rvaGiUawMX4azIRQoPxhQYj0KPZz5FwNaG0levwAR7g
hw9jCugmVtZegNYnXrZBVOUbFKG71AOLfUBc02qeVNYMAZDX0upSi/ZXnRofjy+eTsaRQ1d2fo0l
rU0RHKM4bugChu/xoz4B6o+TiqFkwyyfgRCH0ruagL7pBMlPscRp4HD2G2zIszhXTtM8DWmIOygf
PrvXpt01loRuleHmOiUhpprxIKod5yhGREFGDzwXMgt1Lx7rvR+Igorrqha+AZ8YNKwvFNibR4lX
yI3Gekm8z3UHxo5wen2DETAodZWBr/4tjamVbgbwJtj+4yA7sdudiK2LGW9QNihTMAUbQp5D/mhu
vbfzsU+41k4WgsiRTsdBe02Slipa+IM26jTYR+FLvHdfz083jkhvFT5dROH6qOrild4RsQ1KFnSv
GSzmQFEcOMtBlV4faSLMtZMUXTU+FU52U1XepVbeli5PZKtK8QpLKPnAn8pnXmOWHZrzuONNCQoB
i1kiDknQJEMUxbi+a/vmQtl4+6HMJMgEVxvXPsXYwNYHWO6Z2auejn1nNO7dj33BW8Q1T4YJuCSJ
dy4c4gSEjE/PT7r8bDvzSBGyV0OupZJxvCPZc1KPbYWoQ9ctt5Z9UNvgOngjszkwYo0VcE+Q1fYU
oVfSIKk4fz2rhrPB1Q5ZFXT78JesYc3H1G3U+3AZT47p4PqZffidihrm5pmMkORDym1prAi/v+S+
ZRJuAAOpzDlJrG7B3Suxwtuo7Sv0d9lwexo3Nt2t04OJIkoq4M5EYhiolBe/6uHBVPi7rY67I6gi
TZ4Ek4jcMVutul/HHQeAjweQ9kxJ1M3j1NaMztX2mAc/q3ZXahBU/WgyD+ez8W4E4eGJp5C7uKUh
dKvGVUsNQsG+PuWc7Qq84Cl5MSlVaP0YzO4rkmyZQ/JwWo+LpQpQ3BtZ/h9RJdLKxmg/9CuAOqkf
MnXSgqq1F/axkMzcZLjxltILaKZrM6JD9crCKabt+EyJOdgjeCcEfif3tx7kwX1gEsZlOj1zPBLL
JmFd8GUvtD33Kc1aPRq27zVVz4qG+RnRVtil9oqLgfImcwX0M5C/Ee0fo/D5/Cdbz8DydcPKY2sH
Imxd318UfQZRtV7xsnWoOauOaXCSCTvoU5AZwiRyA9riL57ivXnqWqvPgU0jVvXBgaAa6VwHfQEm
mNThqAKMkfwApYryBWeuJ0q5liCnf5f8ODQKD5WqLW6NTjzfVwJ43LyJu2/5n1occRZ7Md/QuNUi
BOfFRWVy6ZqP/6TdD3yz18TgWNDJos/b718jY/oQN5ZJnOuozA5L91iA/oMXdUpt0w8ALS7rGgZ/
QbHKk4Poc2dGjr5GgBUFu6I58Yy2Df6sr9+QofieK26dYmIbXGoSHTICSAMaexbW3rJl7boK6PD+
o2qlPiUylwSsSC1Oh7OQ29L2pX58VnGwA3FEmJMw/vBZRW7l8VCCZ3X0/9PFMRlhETO4u24t3d2N
9R3lLaRL89Ry5uoOtg1VfES7YNoOBZWCTqYgpVXmxsDRYAKMHqVdP+9LAQTelyGHENqQQrM5E8lg
8klYIG/Lcr+mAn6dNoPgPDVez2IdqxMzi3xUo0mYc//4e4sclkVs77nk8PdwsLGWwL3vq2T37Y7v
HCqb1Sk9gz/tM8ajofKJ0o8OhoE8bIBWD7U/XByEhtmBt06eqfgmf9lIvUJLTQXTtDwUaU1DZXgP
y8O77GyPBFs5iwYRFUok09UwTxbmCH2zrycydAxEGUKx0ySO6CgdQnaoZw13eH2CVkIs7YdNGlw2
Z/K4bHOv0JDN0v9rXshdDHttOdFYNITu+qh2S54rjH0UqTFMh2Q0srtQsdOtoZGe3+G+NaHhbfQe
aDIIX+oiKfHj4bZeNNXyk13R2+xsrVy8S/JnN4pRdxZRyazDi7EdQST+ytM6hZtgUdKcM0RGjqHz
66s4KlgJeXNt/fyvYbm1yW5LXGsHM4D8Me4uuh8JP47+m5ite8dlkO4HMU1ZPIMy7Emy7qqknfbk
d3q6fp2C5xAh5j0klBxFZM7hW0M8zrL89Y2p88cTNQ6dwRPPYmqSn3iR3lpPyAy4HcnfNR/qIIAp
6KkJeG7VQKhY3+hzl3TnHqJE3NH/6/RsCd19GFMF9fa5ZB6XbgrTpYni1fyu9Ofn/09PLWCW60au
feszjW6Ja5WafaPSkLmAMOKEcZnxADmVegsGbKwOMUySq6XY2hpTG57LYJrYVpcwpFnzlw9OzrK+
9GdKkccvMAT97njfQ3rTlViHBybwgBYT/Wo+SMeRBTRWmUesXY86gGkgl/fVLx8+ky5oJxCnRFtp
Pq9qgUfarpjKnk0c2yPh/U1vb9tp94BcnMtet2PnhTgPWwDXGVqxKj1tfFD5fUOTTPs/r9V/1V2m
Borecq0prMnBC9MObzUjaYlTxxT33MaiGqFKkqYr9IyCY1eL46u+WgoYZ0QTz5kXZyBAyk/E24Vg
YQQR2dBMmDoqSnbG4Y5P3ivcN66aXmGYeMQrP/2fhR0jv+G7pQx7WKD76rLAvK7DN9yODmt0vS8f
AnMwtDa7xFgzfH475FZoiW1W91fWwGmrwEsJFn+qi5kNNwrtgM5aggLnOanjbTJ+1qoFq/PtDY+L
hejCoad8K5dJgHCz1OD/o01onNC3neCyq9IXc1zJblzF82vynLsD7KryqPAt1/RswRg8Nu6+C/61
tPhGO/0MeF/9bYttDKjPyDz2sXNQpYVPoNOnqqicN1eLNrnuA8larCkbVbOG4cdEsue3Xsr0oub5
JlJ8h8fltdrjmKCdkDrb4OpiA8Yq95JXpip0x19CkWpjAhtozz+PZUQZeKP8Alum1ytkfm0mt/ec
IIX9IwlkkDFWjCWN1OQKmupgnB+z2agH/nGXb9s/r6b3t7IkPn2bl3UATw/VxrRUZWpJZCHz226w
nqB08JX+KHqbeoAqG4CEYHU/4dBR+USiP2Litzyaex1cO/Ft45Rp+xWfVNg4J6KNnqrVzqqJod//
SOSVCVRyz8SkMhULniWCd5cSrziUOFh0g1W2eajkGWh+dypvrhKbtmFDCpAJ70jWuSQ7d7DW1xKK
0wJ/jiZolJOjBKNfX0G+J9uOjBEwXXXrE7Ta0CEt39K4XANIBo8lk8e4OixCfqKwoC+eVWzTfAVL
bJpYPz0T03QFqt41Ov/umob13wC1YhJ97fupC6ARzQCdIPLJKTVPQVJXtf0jICPkK5JFPULdwu17
bDhpCloXoMP8bBjhEx0Y6mVqgyFfdzbLoEAfZ9urhKxX5PJi81Z0cKGIUUtxR8d+QpqY1lYpojdf
L/5k4/qQUndeCOgIJiPkLP/DrrPYz6ECB/LGl1RbY+yxSqFwrlDL20M8Lu4FbNpGMAB+Sc8HvevM
NKdSjniuR7AE4YZ98YhSEuEUlXuAlO2mb5fSzdElxjQVPiOBcWRuimtJlYTQX2FRUNf3A7Rnob60
/ofgz2gdQ7UjvyA0GZV0a5DYqJeg2+Nba8o+fWxP+wYiNoWG11DxHZkMrvsBoXyYdxBJf8c1873E
hyM4hoerJeG0qJMqbVsMFR9JtJwaxtjINNScUd4T84Ge8lSBBm4eks+qMw/3e5qpicvCdC4XcsR4
MkdfLRmDHNu6UDWBiqFbui/LBWdXpS++UUtshayFLTK6RBc68C2DPdViNneLNSnuVxp7kyimJyAE
P45WOmbl5doEVPZ1W1zXy+asbmu0AcCz87pkXHARoYTyXxpexZPNEG6cpx9mAdJoZIHMkFzNCZdS
80Yn8RECNGt7M73sRbWlEOrkjjkfl4yT22y7N57k4BCL77BWbb8d/2cTMMwgyusxALxqccyaf0pR
pJKfl4e2r3MaOd+d22cUGh2Jw6VHIYaX36/+QuKupxk6bLT1o4kgv4iCd/19wGUJkBDfp297vRJ+
q0Fiu+ZQ1GCOZs9ox1xk+SO9DYaFC61MDJ0FEzKsKcLsNqckTsyxaY/gVTpjrUBZi/tcz0KduUvY
JzPTiTd8tHsI6Oefl9LVCc4I+RNtm4EVvNCzxUatuQI8zf0bCieNtEBbbpwjAAHrgHRtu9Hv2XMo
/lZ+Ov//VinMW9bjf57FB48Gpz4gK2f24XNVKMGTv2ZGfPiFiIF2C28GtV+96tdwXrkMuplrS308
lYXKv/Y5t1Ktx3ezc68M+FLojRW+F92pdYSbKlTkFo9FabW0+oBCF5e3OXC/fD15loQ9JOw89DTo
Rmcw7BpYEkNrgGZS2Vr4Psec46Xo8eTnCQMZQCLk5YeSYq66VA1nQj4YvFhp5260jc9QaXbqRvyF
kBlIa4v+AAlUIEvoNFtRJltQk4yBBmvQuvmawmbvoNTbcsUzbxFYUeej4AXk8Fpe4qDk1JiSgbi1
zeHG87SvxN7cpTDu2zH7r/X/WbPUULaA1fhspNm5CTVXf5FATduDjoD4XqYb+9Zh/7el2KuGwyLV
vhE2UT+6RIj+AeqRPDEhlGXQSr1ZaEFkZb8d4hUlFTzuQqmHg437MXEwzFf2iIa3cCLxlVZyz2KQ
FM5mMTwtlEIXZRbbf7u2mlJOit8g6EX6Y/uKq9vqfF3+LDXEV/hgdPbg7bw+I3twKxWI3QJdNqBm
tBTDA8X/ovL4GN+AhPrO2sg+1Wb3HY+1Ys+D7OL3obe+dqHeMMfMoGwCTEpvgVsWsgZvSyZw4qyc
ZTyqLD8gRyOQ8T1HzGADelbhj0p7m0UpKuUJvOI20CXuVAx0+vHfgrL1QCu+DB11pqLP8BlqDb1M
8FX8rMrcGDLc95AwFMgQBY+elbvdoZFxfwieuOhEK49bLnJf6+VJMAgZMIxIt4hkWYdT8f2Pr/sJ
1OuMZo9RLl4PTBJN0F1CrdOjLkhzJmdN0Z6eUichAd0zrT13J2F4/6kMKyYChJHSbhtzsKxIwrls
E+LBhbu1sJ8cUisQFfokdIoEFPhpRta6s+v68WyXhdFvjfVdI1K84rdCShYtRUuu2uP9B1TSBocu
RjY60c/Db7hPQv4ZqWbPknZ8GAxA5uWg/ojZzfAJLxzE2UdW0Bs3ElaPfkL3F6PrXy8B9dLgFJQq
YuMx7G70+FYlYHYWspxvR8O9l+CrqxXYWlkZcDHDhU1RN2IjNzAAkVAwNvQx5U6T05+d5z9/uTEs
HdC1r6OGbKe0xMg0S1nr+mr30byvOV/gFJcUQXpxvr46liddYjiimhLCVStLu5j1lrIOKwRGF+hk
aX6cDv5ajZXxiD42ou2ouaq6Jt7lyPitN6RDdubrSdvi01hFvK98ZXkDdMzBtj0EXSkb8DNmVCTp
j5JZNx6PFdP/dt8NSst0z1u8TXSS4GuyLp+JSPeCJg/tR+S5DSnGRNXRHOvxHSsbvLEMvtXITAjy
R/aeJv99aBda4TlDxbBmTO71kaylYqtIE7TD/+Nt/pmNg2EaJD3b99lOPRihaGNGc0+rZL4gX5GF
Vp0r4Up8tQyaBqs8O43aLOzlTO8MxEZepTNgVRQjKDYAAS2Jlchi/dc1NvZAkJLsyq36nKOkRUVR
S7tdpJlRak86JlYWQZ/omwQv0qI7QmiVyAYgauqsu8zDMUJrPdNUShAPOeR6VLx6x1015QwJ2mZY
IyrFS/15aR1CZrwlyv9KxXKYZJ9sqZ6/3s6rDp84giBSM4y85xqc3QEYUZNa/k2B6F3JHCCyXdbQ
mlVjsKg1jmU9oGbJRfsEHuhDq2McS9js2kUVnYwOml5xSkYqKhF5XjeXKrtk9JgRzbOMWL3wiTM/
E+YVfhcnQDIgq8OP2o4MdFFbXqG9g7xXGFRZOUhJ3OumvJaRndSP/poh9MJPp9QZVt1pjn4Tq39K
f9Aw58keygAtPWWdVKoK6+HNrIXNO1qKJfF+5YxjKGVKHllkRqIfxdGb7+RUEX2ELUFs+zDTg6vf
d1MocpcWc5RjkouLqXRf8fN7nW5kKnIdbwHIA1mii2R/D6fFPn3RDgnbgF11g2pPdVZoTO5TC5Hv
Lqp9Zkon5e8z/JeU/r9y0LQ41SdqBewaNiAv/ZwZmHlk+dM+qcYd1TI8MUq7CugAKgLW5ZK6+8yh
/pV5VSYhB1wKOshRTvisb+59+u/qpVDxlSKIXYxEEcaDJ65Yt+ZC4wuv3ZRNtpQ9tKiOPNDN67FG
IfHEJ8GJ0JryV9da24i8z88WoilkILhJKSj9Pc9wVZ2uH5gZHyPgba1+wYdBIC2JRXLuAQpKevfw
MduExlNfTsssFAiORAn+W08EZwJ5++d7w7S1OeS7xLg5y1f6mW7qTtdivvgt/aJZi4JGov3LMNTl
W8+Wr6mzwuJcroXqbdOJv/rxo3g2jtBgt3ZiIYViK2d0Q0FXti0mCVPzWWoOsWaukI+D66kyYd1U
rNWYxrq6xFQzli+6oewJGoZ78b6962lPbnK96xvlB2/Cx6E+EREHLvTo1skFotu+5Yd4TmaP/oZR
0UceuHlhBztOZA05c5XjcGy6viG/9GkiEpIwLwU2x58raWhwtXnxqO6o6Fq6UYd6xtvpt3K+m8gj
NwaZNlxImGaBkNcdGgc+kkOwheyuAzuYBxoa2JeJ5qt9/Br6fDc8zNuAYQ1BiRWlD4cAJGiuvyAl
yg3eECcjlT+3cZZFY+7jntuj2wWH1QWnqVov4+dM7DtTfR6ABwKwVb5hXSQgC+uOIfY+/WtO62fP
rrI9AK2G2VUz+ugao4zFzhS6dAqQOcMIGLbXJSp8uvoAM4muLcTXJo6pgqNYe8nvdTm/9wScKXFF
jpDdXFYCjg8u7ttUmTyhmtgvlGYSlpiXP9H1ehOddp2+0vph7CAFtu+IAD3MtUJWWFE+RgZeqEfo
hA7DGGd+gemFr15QPbVjDYzl+p4yRW0EFr1Z5FTrZbLsLCXjBqd9WGBMETqHe34Q65jM4y6XpRh7
xgzpBLaFnvta7JwtfKcqQdDeCG0mrzlbTPjWEbMDyDaMsr3OEWPFUTu0PREmufWE4EF06/boGqtw
MCkOL6VlMOBjnQ6hyt8C6e5zzuCNjYhfjS7aJTaYvOIMeZ5ZUSDOEGuHLIiGtc8+wrJu3A0zRUpG
uqDn/RhwLcTw7dtqFgPcqyVLErok7wqCc0dZtL3Um/6UoQBzYQuxfVsHZw2AtQKArW5qadINOkvp
NNojjRO6/k6RG21vsLYSFv0fQRM4Z8mryOn2ekzaqMoAOTjWJtsbwECMCSi5nguSnEzH8QCvewuX
GJdb+E8N8Bp3cO3PPJ1ya+ThvPh/1DjaDliOz4T2sDC78MSBrOnheVL7yN5TR1UmTG9rEZie4Ccr
OEURyafbyWhJiWyAhRzdFGAQpVP9Y1Ectyt2SViDystLNHkfYT3qj5cNdWAskN52eSxuDtJ8vtLp
y0Y91SePfh6mAHrkaOtqFFhwt8NEHf5h76z6K//LZrdMENS81eH9lKFB4PvgUN+rZ2FaxO993FPB
yoA1S0ueIhe000ZKDR3zb/mOhDR62DCxKlxx9uwgsgR0Hh8varWnaMdco3dPAZThXASVW8lapoNm
0W+eu5VejJbANUgbOO5I4d5Nlc52EeZGceGeg5jyxdOzFD+5IG5DUkftepWdsvGFS/9hKXNo5KdF
9e053Gnsl31w+N8dIBZoJOEfwA4gtLxyfB6CVLHa7RPk5hnnoHURzwAQGdbS5Y3eq5563mLG30d6
VarskKX/nlcV3stHcSSC+FfRxrhRIRuyrzJi8mpIh5Hw8yt7wM1UTEH3/jN32ScUSsIYfQeRohBD
aZK4j53UDqtvQlJ5loY7MIUIzZANr9ZS241fMqEq67zqUZVqkWQwXFUj3ODvS4HRmJF7Ov4Lg7v8
XhnJKBimw+BKvcCfGTpn5kJzFhVPdtuR8Re+lFZRR7DHAS7+FwaAeI2otwPzcRat27Q6t0bjjwhp
yLZaW7nd4d5hia+XMfUJv5KB0YJo5ikFWpjGdc/m0W7shrWkdmt4zPmdiXrtlin9v+2/qXHaeZM2
CkyIA7H5gKnTdphIessTc4WH6l/kfCoqMsHb4G39HZZk9Q2EvMfu49qcnb7obmKOIbNro3Iz5dTi
Vy/coDe1cmv4OasLbC3U0546CU0OVMkRko46wyjQLnteLM2IQrJncMV0MtPNQbqePMkRsc6NdH2+
JkHmgMsBXWJYac1bp7Acaeea2ZghCHHGOLR1bkptNNT+c21s+kfC4eVL8hezE+2oN0kuvHKAcbkg
suN11GKBV0LTy2pnKIMKsFz6Pcu2Xzasf3G7NL43ULjUBKHItHcBvGQoGpIr07G9j3alrAEFwZA3
Zr6bzzaLAx1yiGc+ZHZANrZhJbMMf3JYNzbA61RjI0dVWZws8TkpkXKLNqHeMV+Wbrm0iwHL0bvq
F0NLbMiDuc/hGV4EBXO0f8dw87H0f58RLwO816ODgUdcO5xO6QxaDOz9vZsf5tjq+nUvlNka6HjI
R9kQD/efUy+VwvsoE8R8tVX2U0/98hBXZlwabId1rWsDTiITYD4smAAisYXng1EgNuhc50kgBC89
g7CF9DxykJGw+PX0S9EL6vufhAxqrU480PKZEh+Pj0Vp6o3a3wpEoEf3BURdObIo2D+zTfzD0t88
tPO0+nHQXFVFi1fmGka08heV9i2puNxIGm1seKc0ERq215HqLdQooTDrbkmVT6bwfedPMxt7/GT7
PE+R2SayKjbNpxqLjx6zND43vhbOpQxUYssgKxlq5ZHtRQyZs8lyvxfim/dsdkgTQ1MrfCtz23ym
MTkv6gMp7VwG/Vzhw6gJ+KXDuoRKTvEUwVysvKzyX7cKAoB9RDNz+5iujiSJeaO/cWnQszpHAR6Z
xHnbQIlr+8zyxi5eRVu8PyR1Fcq8SCQ3RQjj9ZElz9GI6BSP9O3kYQaIwBY/FLGQR04iK4uy8qq0
aPjuU1usUXFT1KPewj3ElaIo/ITyOrCGHS32GGY1+kgCGvo83zBCMOtHGJvvvLFFIWziQpCWDHnK
NYssE4f9ZBtzRX9SxZwxC1i2yUY/62l0CG8e5QR5eqDQ/T3Ku+/OJqBTz+U/GDO3YSQT6RE1EL8F
0g93d9BIQjwTkWIEwku+hGxsM3ctePzu+F7G6o5XblYcZ77W/ftNIlZqYbsQR38ROZJ6HaHaUJ3F
e9Qo/go3GqTDVtWyUxF+DBukvI0XYxtOGz/5VhIqqzJu89W2yTsKNdh2HiJO/TiXKlWLMdLUtpIx
ZRyPFwBQ6w3OkQX83rsZDTTc2psCgXrubPKnfQkhZrxOjxwW20xQsKa2SpwTnZ6fm7426RzG4747
QJjLqq3atgtH+j4ZlsI7gNNzDFUAw/Y9oVABLSrD4e9gvIjMx03nZA/KbU61+f6IKD+AZYDmClvy
vO9lr7P46WAwaj+NS7X9xftirO+JL10NDwX+Agdhgck2I6uhK8JSfSoWCe6BW6fKHbh21Cf2wcVk
o5Be3b//jCRqS4hwLISpEvaq5yueDtDFF2YzO+K8N9sgB2JXrF7xWMoIt5Cm7mesCaBBF0CT3jxB
kKnziTtyll+NqcnDWxNL6sXZBy4REGbHlY3RlhoQGlQtQJfdYZIpvJzvQHj+jo0aS3kyUJjvj29+
bdciiXN0wH7sM6XmTJoCNow9QG4FPyUsPdiRO9P7LHnr1mDDr9pEVHhQsElurJum9d9V1xFrIDGh
cmxraxeMKtqkQpCN3Il8yiCCPyWMYcVu7qWe1cqJydrLd5+VbXWNCX8C6MyNj1VFpTcEXuYXcJ3q
FyNfsU2Acup7B9L0O0zlZ32U3UlCbCWCPHZYZGEZmQptn9librIxRAoPPMP/JiuZETJBVRBa8Mu+
M4tKU/cGjO5K5qYUJ1snCCDW+EBZBJrMYvxRdMPMkDmQLbeDelOsXiYnU3rKn2yN7yVuGXSVUjT3
NeQW5Kq+sM7g9F9LVl/tdMh68E+Swp6QQAk16eE2AJL/hnMgRrO3h5yzJGukncnWa0Q6ACCsTX5S
56NKh31it67UEzMURqufhAnKBmvtgSqe8flxIAPyUZZjvosq9lOgSRcu0rqxCJHnLTmYaA2DycSt
wvZKJMlPsocJGlt3CzgrmMiV8IhKrbzli3beleDFQ4KN7sEZCRyXw+/Y44/otqW95d70GhPSrSHX
yzvx6dGZfvYeOenziF5ckXkK6yqnJKkGeCEl+HcIiKREHcEoGunaE315k8thMH5e0jep0rGCxk5M
7i+7WGPGsRRo547ACbLalJ86Zqw+SLtxTOSLZ6+eqaB3Ss+EQ2EyDIYjX9RAowHnXCG6yaqPLZbM
KftN4YXyUoFZD3NLPZbh/bg34nJ3bH1iXuDOQQBghlpQX6guprtbIBmltx2zQ5Pgn+QjX7FViyzD
x5s6PsUtcIYvwvJP7nNhf/KxcLKO5VV4nbDPC2t3UR47YdrAW1DxTlH3ZykoK+Jd1rwlTfzMV+Yu
DwxECw1ROhSBGtA3CljMuXKWfcTF3BwuVZ+j0nLAj5AdDCJJ551NssH//2uUtq3kbjwv2D1cd+F1
LT0YiiPYSgTTu2GwyrsCh9uBYc8dlGTqQ3s8o4bZNyPhdYX3VSJWKoM8iB0+IBQ5wBWyUBtl/+MS
KZWQWXKuIjv5NnTxYUaiXPYJg/AbwtI355NV50/abDqHnRT61qb5zwaviWmfrYkVz9p+bx7ubl9e
i2otX2Og4q93ftKs10Yvylx8/vsK+aGxPpfKKRMQKhKFnxU/C2SUbiZR5tglWf3I9wROeLl1H0Fx
1oF0t7yIDRtRVaZZsgUCgJpOlWBANVHEN5kIozEasKqMTxBMxZMStqVS9xnGagVUcN6HUDL6dqeW
FZe7Gh5prkET/9IJD/3USl7SRybrsjyLc9Ma2trnbba8BsnZmT9XBB5lEZfLqB5AXdPsMKbLlVf/
Hb77Lxi6m2fZkxYUfsqt681HR1LCwFzUJWcYKJvnI+sqScD90RZXC+4XAlye4hfkVy87tr4mKNLj
ZTInHJ/ZQ/Irmuf/QrrZ5YTH6miXnXn4sHKOjo5ieFV6IyHACmYrP5xVIH+0pVV6ErqIcZADl0/8
p0n79bsczGJL9Pbn4nJ9d4kPwG5aUQ5+S/GJeDxHmwS9glcQS7iKhW35j7akbWipyJvlEMixAP42
KC7nPzM0Geblgq4dITEqSVnfGrQbhAI3WOk1DERL4RC68YOrbwd+uY6+FNRkX3xoYypKwgphmi5j
padASEw/rFKEBgZ+MU+NJx3hIIwiqpwcN9zCtc3cbZ463J7wcX4t8Dp2FFp+Tcrh9fIaFOWdu4wu
CNi6ZxPxULuQhcJYpMRVE2HgJIGJNoTmULN0WHmWET+4g0TnIWby6ic/wGqI+AzmjJpkXeJsuGIr
j0cKgXqezxQ+Rae0PdYvoc4q018xG2jO/qMgIbukHpzCL9U1f3T+xfGt8wGJOpnA2fpNvQP9Y7RU
YPRrzQ+snK4FbD/vQm2y2v3J8lIfqGQKfB5DaPTrlsGc6Chk1r3RlU9xSgXUR2Lu0HZrjFIvtyaA
MpmEvwBeiFKcQhSw0U3aTvV4YhlcOl6LRj/bNxAuYvyP0A5QpC9Z9yINOLTcNSbL5Jsg8MhTXRxc
FHW4HX8LClv76kbolFfsBaGC9bNsxxXEk9/yF33xT66NlKF8iAkuUjXkPMRbcL3xMCaBCNLl9rwc
Rw5299QsdH9Nxapmc0VdOU1JRRMuVUjvLDsQmvtHFrkQj09NEZfTemK4NPydO92k0b3MzmgmtF9B
VB+UyRdFkTvNmdbxUgvqZ+ZGIRYKzRSjatIoUDt0er2qa6n+G3wG4vJ0jz3S53Avgr+P3TqpNKtR
Pv7Oa3EZAHH4hzSddNyYS2t5clhgb1moOhdaoyQDogzehoKPUcVouN5d9sd4uy25lFTj5xWS+I7s
4rmJ+P1SBbwSSnc+im0bFm2oLj/UucFRzyLKqsulydt6ZfNkv6qrbmKL3Y1VJ2QWOBr06ddwFE3E
gLh8sdNMg+qXOr30hSwD17zVUNVOGfUzGVNqTcHI1Bj114QY6KW972VRPw29FDZ8mhKl4ZDAHSQL
K9N6Vs2KsTaAQlKgbVYg9b0NQly8MrLbXiNYJiEzHqW42OvjoD3/TS1xoEza9qtt7SOObGxrY7PO
oY/HTIuPjxc2d1BoTh0MKmc69bXt8cTLostdpLtovD+63cg0P6Fr8Zg1lr4mLU3vtcF1FAUpS2Dz
1vNqpFjOhzc4aCrZ2A1lBKprbw07M8Xk4/pKp4KaCQARAOw5JE6RkdeyEvPxF3nfJ3PezGRYBvpY
UOlDe8Yo29Xf0RqPvRwbRGW6Zl76o6ZwJQ69KGWqGKnw62BRYC92npeHO06RewZLdNob3qeaK8p6
Ep8ABdDzkYSK1XfOmF3OBcMA9Vehb61p2hjH75UlGRYRx2bfVSdRnkK8WxUe6+sHiktEUZ+ELq+w
6f8Fc0VT5law5vIIq9Qd5OUz5wYJd1EN5bQ1mma91DEktYpRdRxflViMpV7GIJ0tstVcVazes52j
Imy+PfL73ySOCF6cF6dMyoHVclpl0wn7hHbdzxwWBM2+pRt455+I1TT9pb7YfPA76yFEriub4u20
ONXFk198cDYUTB7PfV4v+lAj3jd69/oNCxxk6Ac35OmPeRMa6RgXmDjmvrn7GeswuCNpVRuQb6Vo
b6QLf+QmBEwe0W8tkfG0X+U20CmuYORLsCfc7bYDABrLV6OjP6ZE+f7i3qD4TM0/nLFIgipj6JO5
IaX0wPV8AG88gN14Q0XnpbRqVJzhk8YVeR0KcgxFEjcYI73lzusj0vLSSGv0nBCY3bLIo/PnTfcN
HSVWrfIEw1ccJvOl8mdD5VEWR8W/bd9eO7fXF0Sm88n38uztNVYJjJGu1EMLWDIdI3TKVnzHjPcA
nBiF3MLCVVdiDccNgqxBsfL/3/KUE32PRardlojezzc1VsdLnud4qfC+PBfihnPRBkDmRtJBcSxs
L3dR+FsVUrKyMcXkzzSG5vA8qtiLtjCFwdwmqiH5CEEJyQVIbdGOqqSNOtgz5mNkPa2WZxe4gI/+
Stu3hxhH/unqlMStU8/PXME7YIIwRga1PwDsZ0YATdUdd2esLEU25CsJ18c0Vi3O5t2+jJezLM2w
8ZyR1FbtmP4CCfosu+7McAfCG7t4CqVDhwwn/lgre2Y0uLHQMpg4caYI/wuX6Q2JWIAISilJGGjz
/9TYCSmuOW5OGx9q2kuHHirV77DlO+uTDVZGX7mimTzQ8nt8yl3miq22NVd3GXiQ7n2w2oLCPaD6
qfjgCUmpprvNDvSiCmdsSVFO0RiHs2vFaxv4VwvI5sJDcxtS4rbES20lWvaGQpgeZYl7WdjNJgde
a9QAn5TPtP1OGWkz5bG56HquHl+oeggxcrLw3teHubc42/wVketnzE4GXxADNk0PamcFBxqV4/ti
vNkp1XBxnpKvY0pQ5a9RCTv9I8p/FA5u4cKtbUYsBUjejXYNIL/znNxrFLwCKeZ0pboOCkkSFSsd
6XHk0NgH3uw8SqRMqDzQa4In1s6WaF12KBMJyTyfuTgBjQBu39dgU4/Ub1O6me6FR8PPU7HxC+zX
DTO89y0TkbtrsH2SLM2zN26gaDEkk8XBhhjPAJps8N2Q8N44gUI91M6WpN0pPMoN5eHHG9nBv3Ca
QnLjNb6RwctCRp17bLbkHOiK+8AIrZ8OXdqdxNeXtK9M+PIGnE06O0C5fEn4CM2b8Ntr/WrebpeR
Erbyvci/WlL2Nl+//sm7NAWO+AXP/zfpzEijPedHF/nWfs4TrLsRs79nIntu8TuRgFZC2iLztzoL
ulVnM8Jtm83q06XfBjKcBtjTkyt+JNWoyeY47w3vpD7xLAhCLIkQEdnapm5mTjnJDEGn1XD+r9IK
2GyVmKt24G7SVBsQ20yALtYnD4VbvzEV/1N/Omy+OVXSOco9T1Z7m7Qt6OkXVRC4rGydFheYjfPb
U9gllADqCavAxegarLmXOWtTAVK1p4aUAmFWhIdA6iBlWvachWgKA4kAYlSSJ78qTbosYE3TPGW4
6/RbvswWi2zVwIzSAaS7/jVJT9Q8/ONPfEIunNaeT/z7SAPnC8VW6kuXcAoix+8uO376GfYQ7v6+
A0f112lIIspXGzuvSbjBZQcA8+45yOi0QFI8cGaza5s5ANUC6LLz1dDMCu4ovX670k64vMkVHH2G
RZvXMB5fCFPOZZskOESpkCl2vGPSW9kPBGF6wZHceotZzaX68tJxC68CRx+WQqC/TgspMcIMyKpu
9JJFcaWuNEXP8Uo/3tPGE9DJglGlwX11h4pe3T/KkhN/2tbF41r7HQTOBlhRf4yPzO/JSyTMDolz
H1aXAxXX2wsw303u3MGnsnupvWWzm8HnFPWQc2FzPmUENY9+UMVDBb2U/xBMSiQ4CQ8cstsKpl4o
XymQl6fy6BlQdK+oJrj03QD/smx0bdsTNW7F5V7cdS9BMzRkaKec0yHN7MmViBi5P/Pjn3AYgLKC
mA6pc9HpnNBXXEwv3o67XESkl5Yi7UyH+BFpa8F3Fku0BENx6evNuOJgXPxXa3BAOlD+sUJfP0/m
seEzGEqlGf0jBVNBcX8pY9zcYmi+j/tpjS1sbCrH0rmCJDLo/gpZtPFiuNc2VKuQoPxx9BSAz71J
oFeE9wngPlhRsaLzGp/9qPEyKp+ElO6Ov4olgChfwC2dHailXa7o9LHqu6SlHhDMu8iGM6gcqh0g
QwP26+LnGGc5QbNxH74OX2qKwEDBBtSWMsFWr4Qfa7E/4u04wVYwgEYPiv513dzh8W80fTdI4Cxk
jYSS2nbOujD4lrvE5S0eQRQMywfVD3kubpHqo6JiYTcyFJttFQWxSBtcMZGOHiwdy0JJl3Efv5v9
09DjCa81jisaJrHFdeRUwMY6JLaO7J+8Je98pWQd1KsB1V9CjdtqDUam0KisljXcpEHITRVZ/LFC
xbFy6AkTUKuTfiOB/RODhHsDb+9JN6bUSX1bK3Gb6PwmWBc7qiWHpzPEMPhTGwKdCJ5Q65Vad9a6
tN16Q4QV2ZGDv7y3ZXIDB1aHK5tx4t15Woxt6RG4RDHcT2pDZdMfkwSf7lqrCu3MH3uMKfpde0pM
e2MX//Y5BT5HD10fL6rxBR6ahbhKW01V8wvQyPKD1x4NsPAanRPbcHBdYY8q8M0APdQq4u8RDPQF
tlM/0qvTDSyMMOdmc2oIG5CaeON4YebI3hdrG3AkPkIroYDJI+wnvwL9cfwqtTK67l1HXv1iec+/
9jYYQ8hmQXTC/styTInzmZ3ZWVMystEoHZD2TDSY8c4yS9rY+5EN2idoPsgvRGWHPLY937aZo/dV
F8t+sexKWpcng+Oenp6TbzPsCkUkFeMvJhyezgEWh6F4R+rfAljsGK5+ICPxFugeoHC6VDM9KCaA
6TQRvZ3mIHmE4OGT2LCyhuYvYtRdPBh5tOYpfFMyhCWOb6Gzh6h1UANSMwgNLg6YeHHixuip5zaI
U/+iOpevs/0ys/07gMMgSD7fsqko6qj/NsVcyu2NljEcNbvJtL8i6/+Kw7eEYIrpW0pLUXigMoGq
P+JGy+EHDHgFAb3e20iXfuqVgfvCIP+uGwOmdEQzrHClXP9d3dKL+IMrZ/fece0fe7ECr/+ar9Yf
03n91seowiZG751GSlTOSRBDZksF6d3+5pKGOzapvhkPjmzrwyEESRQCeHrb+op/4zb/EL1k9Rqx
357SVz6qcwoB55lAG3dE9oidGDuw94AUFgGX5iLKd0oIkaQ7KkfMMpCtacRrbxVfacL/Hyy6NqUN
nhQc/pY0H92rUk2FL5g3N9EFVc7Yoz693ExA27t5kP/twR/FizbwXIEPBSy74M6M1auSLfyIZaOd
CCs9UAXmVcZCa301943JNMpKfEe1ayPYI4khMH4AVVk5rm5iSLhEScwOtQXjfsVI66WNAVwg+lxE
OA28tKairc9o+3Q3Vyxkx3VGGhWpqVVernmJBScocT5/Qoy0MpkdK/DnQoWU5EfDAj/+dj17LQcy
n+v6POcUiPZqDdYNspXze/UhrZ4TiUDSb44HtCKNbdAOpUv6Flhz/gbKPWyE4R0ei1726b5NxQdU
Q0A3mXSycex3TZWhgQAVVi+svqb8Gy/mMYvSDlJb/Oa4rSPWdjqmPxgTqmJTbaouBc5//thpve1U
dWg6I/z/PQCIptrRm1HCCCN0B1OofFC353B9CK7ZioI1q0M7cmik/oAPnTbBYKh8l+9mW8aiy83O
0K7G7iVTq8q2s4m3mOVPfdV9SeObXCRzZJRonU9ysHpqUr8fL/8Kf5H9FDjducGTyJBBEcaUROsj
aw4AF7RyN91FPRgGNws0d4dSgeLBbsKLA9Re2GPvDWcmuNJPFYHv0JxEmvqx+Y2HTQ0EyWfHa7m4
Rgoitwt9UlKp42S8MA4UjF3qZuX93pm/yigwrmHSSEI6C6PrnoT+rIfJvkJAsHHN9/Df2DiN+ASR
w/A/+6WYqq0lRp04IPyQm1g8AG/touEL8WZM/I/d8LuM2Yu/3yOTbbsZPGCo3BXINw8doJ3LGhdp
OXMNPKSrWcBszZM+SHbW+9xrxBRpo4FbnwVV//2MSj8NwDouYfAgGtkj/83rsJIpijqDK3PG3/f3
aI/OrbqxVVcEPHhT1XSMTUSwxb7U+c8R/k1HAL0VlMWlCe76Mutd9oXD1IHHhq8NYkqrZ2b48Sgn
aZ75ZHNhDS1v2qec1WlyvCLkrupuAbMF9wjdt3razwoUiw9DG4FZ6DFBLhFrYhlVA/uoGs5GVV7X
veuXuzK+Bs8grRdOYDCcNuoAk2hHa0gG8QG/+Pr2NG6U8gE9x2RPL8lRF69p6AfgmPDkQ7Q2TkA/
pGCuGtHb2Z4tIzViWTZwM9rrfWRHa4poV4orf6vOmuoCbSRod1arpmjZ6hfJwI8hcpTbC2lYMBRN
UcQEAmAlvvKJlap15F1iUzT8ZB/O9CipySvdTClXjonSs3ED7DUAlF2Urz0cL73p4Er7Yj8LoUPX
wkePwfJsuvoGl6GtydiiubZfB4UxXSwCR3EXGmq6V06j4AzFaMSrlNKzOYTM94ZRgAAYDRdRlLBf
WK44ybHsLnP06Ap0bwB95+5FL7Dx16U0Sp249GDNommU5dYBI7uh2CK50iFhj51If87xR3rMamzH
GUqjHDSO8JdDVmtfFHm2YsBjnns/BeODXCkfkQuQDYXuB2cNoqV28yNoaLvTy0ooM+o6d5qZ0nJ1
OQOR6OG/3a1wBDj5lNdCAZtc1vNdIwXz9Qcy2ageJ8sajuvR4Kj6SbpL6MkZ47O7PzIcw9mJXyfa
HUNQOzeb8cu/2YvAi7mxdN/7DbyLAztGcvhgCkG2JdEBZEeFsSfIVKHfnUC+28SuUMnl9mkP/wHp
hKZ/Y6+a8GSfoTkYXtmMSzpjjbJfypPG51zM2hoYFbk/QTyVH1Nr1y9dRXEBgZ5ZLv3tj/Zn1Rf0
HkaACvSJtxxXf0Nde89avqp24ThLyveKP6ZjPmY9zWwBHGlbD95rLNjQpy6bDxxzDEBmqv+BhSIQ
3AhQVYC62wacexaP2HeyrZqDbDizM3ONMtPrLGnQ/nyRx7jqQ44CpW3OHf4qrQy+TMbDcoac2lii
wzEovHpy4QyP6Nh7zcBJyR8nsNfGBOBeWJWq7ufe3lP1QGEkVN/ZLzF+xODcdHZngRevGN9cHm1+
kFHRJcOR95B8QWyYmollsOMIS2wiuaGzuJDmgGG/nlBMZkXaZ1SAyIwCYkrRSR9p4kg5f56Wl7ra
LsBibyaozrU4s/KzAuY38naZrLim4/bu7+U3gBiSTZr6quFzPTGIJicN+mFQpI/9fFYcsnfxtdRo
swSdSVyfUn6d8eJKI4VpC3N+DEKFgUjZckDrDOxs0lBQP0S0PVZJG55GrGll01estVBwTzwJXEmk
JRcubHVFzSIrSd14X2JrHgq0Ab3l1cZDpnKZhoL/aqxNitHLLICo5czDV1yItxVA8YtD1A53S4CU
JmYOsgGg4mWbg2AQVXhpz99AiP4u/Sf2i8X4lVFeAFuyHIWUnjBBXh9b3yG1cP/VP2CODquzOQYS
pJc7ZHsDKeO9Oq4HegmHOzJbyY1XAotzlYy6DOvxrrFAvuf/N9t61Kv+6eSSgO35mV8eFEVfdDmS
jhFAOf0BG+avjJZJwOBi7AJ7pCcwBpCvh4DeCsxJsdO80GS0v6pvcAFHeLkMuLC7MmPw4B17szdZ
iY6r7CdCNyQvFXC8mLhLHk0eC/PLYVPvzMf14mTRl1iXwer1t53QZeIgcZAkuAQfTkYL7T3APdys
I9ERrHTeaRKjSfqaRbuIMJ0rMUht+FO7fGWcNOeM6ievhXcWBLzhDWpJm93c31nE29iIHii1FpfK
bBVyee6QbEAdBVSYvvDR3r/HfhiWLWfVkc0x7JBGJYjnOBZV1tt6obxmuuohwcDFCITDyN0iEm+u
59bgVyPuFVav2rk3UaPRB1evrrMa1pbmlC66ltKEPR+y35CDuJRqb9hDKeZwpZKEZUFBdhobaFZ3
nzJtItM93aDTkDfJLIPKLWWknTzpjlveU1cNK297TUJNY8FHM2JChqYIIIP/j0MD++WKw6ifouo2
mG4P3W/gT74UOSBARbGOfN0dvWD2rtSG9K3KA5DibwFSPtXb3CwixkMSRurFVVRNh6hnTxkeA2KW
ogeAWTAOOssj5NjPWwlIO4oKQ8r8X85gJUW717fwhDdQTI5Uy6wU/bperv0KIpmHwL9lsx+5chcP
2jX9uD8z6jkopuYWMupkY8Aj7KlYm8OzoSTnwNqdR7x9qqEKoS0WRxdQLohXlYpAHKfeLbG6sOi1
+kYtsRbqP8wvgoIQpsVU/cSXpiCgglx0MsHO5Ha3YBYBIO5kKhJzKhwnTtYSQCR1ARDk/bKrBylk
5K0pa8IsD7VPi1J8pkzJZtf4tQ86g/G2dHH+Loqq6SQkEpghm8rMIdbXwLck90BVZmyVSRL/TObY
rsbI0yt/zUn643j6xfBHYrcILUtOyoVBKfPdvKjfQjyHHHru1MTerxVz/hbhOt8oLQe8Uyk35LV1
onnIhuIclDXJERWHhYxrG+em0daeZL9DLufIx6hoLxhW7bFtqi4vNfljCzLDHu8FhYqMJ9AYIt7Q
gAruE7uWBAQm6WHeoDPR6W1D+wX5l6Zy+GcXD7++Y6sF+NywJ+dOTxRJsgq9k56TAz+eMvFdaBRh
fbDg50DF0EIz/j2yfm0Kn2bJjY/DBp5tON8VE4/lkEaUt7kRSglEW9+2HpfXAGPPkS9Xv2xEG6ry
Vpm+kM6HPfLkw7S2LuhZVHVGKQPUuWylb+f/5wQ/lKj3I0d1H26tvFc1WGFVXxGXyDxg0qDIP9jr
D9S7LOGlZeEpZSyR22suQKnuaQKwAgtjPgkbWEGPgjC0ua8xaotJHdPFPycRF+rN8t1YRSKqVEMz
jmV+ztRqgTpS9rDBQD+0bUSpUDwblLgXVvM6sjkjnOkaLedjcfojL67im+jsS4MQrAAynVW8EsjZ
sNLxssR0E75oHrrfPR9jXEs0Nj5yWAiCoNICDuA4Etg71MjQZazT4HKa6TjWHXhimvxio2DE0muR
AqlU04suSRpJH7rPd8m/nfOWyHklDumI646JgZAQFzZjUEPOGhErDrwcGScEVnAMBzhQsIhqpZty
sOB/YbHGy8V0QqMPFVjMUF+tlKEWRCWOalfU774+46/++MYyGC++yScxhyewN+tu6WgIybOQ0vIv
XIcrTYVEgum44kbE8a4MICrEeafvLYGeuWCU+EsBq5dbMFe9FqnfUUFz5ZrihAuDdL33FTqaFWdp
1mRDnatYPHMSHGM8ybDr6K9FzpCHu7f49Vnh/cFi8ARkKJdW8T5Q0lPKrYg2zfIsjL0UNdG2Go1E
BBJ9xnvj3xpsggpAwimhzy5jxQDiHc8cMGUMygUiWKpURLi0yWSd7aInfyXbG7bVN+wKsSPhrzQF
k9vMjB+WFioSV5PufVJ559Dnas7Iv4mBN9hmZXdkIIiQFmqGAbOrXa3gwHuGSWLoSUMSw09AQowV
SMDxWGaRXIMwRd7Z+t+Cmu9oFP5TE7u6zh/evRY/6nzQZx/LGRyb56s7vE9Ebx8iyRXMx6PncWM7
8hwxVNhb/goU79oZWy9UkMi3v7KjkrZJY0q2SE6pE2ExIjmVfdwJ13vFSPnPEyYtj81JGFKOwXbW
Bd7/qJy2bAd081OkMmGuXoOgEy+uD6mr4efBTKWMR7cIN/MUQQRzXKlDpkV8iVSVr5ZQhHDBnEWU
6NhKca/hPTj78+611rBTrMJsYIc3ry91tXl/FIX1sZloC1WpHULyAGen8diRrpSptZA460DQSapW
y7D2WXmUs8UusG/ldCswhBUhYvvMUvmRMgiYiA20gHmdY/Bf8dp4gaQFHmyisxTg7I/xO/cE6Dnr
6YrZTEl0bpsv+aJRjEylvKWhw7ZY7W2SgH5glDwVH00OOW1JEBLLD64RIAQIlCglWwf38FP1Pn10
MXPua9nhJlJMxEq2QQsyzfYvr/1+A6aC67ChzVmyKCPb7ySaEk5TRWpdLe7ey4xs4w9GdOk0NjSf
Or2nz7xqqoIe7RI9ZFQT/GZ11zT+9X3GalTLsMXaOpJDkk3YxoJq8YrkGePcuHzsHUZ9zZW5m10F
TwmOaULTNWIkV5l+xfAbF2qSZP1lFpauej+Vy157bKMzvfiPbtmVHfoVYWhyitJvxJCjMd9RCUrw
ywlCrnyt4NPPWY0UK8Yjm7uSaNInokmE3M52PMPPtokcpHttkHMy+X01fN5ReoPAc8Z8OIRKcL86
0m7cNV83kmrc7aHKcht+IzhEdZylWYnngrE/5Z7otb7Yfhm59W/kkcT8yQpjEv+3gEZ7hfLZmvub
/lZJuOs1CGMXq2h2HQFRmppgxta4yJLLwmzzJfITRIK92y9fqpYZBbx9lGw4sHPUM6GnD+MLmMPN
nAA4/f6XjQdWwgdOnI7zaPYBeVS5Z9Rat0hi22gKQF8WdYgX3IvvK6eKfP4/2ZoBVhm+xUsa1xiH
sRuSVaiTGcKLlWfIlscwvdD0hqVL4jR1Fd0W2iZ4JIYech6AnTrZlWAgNpYdsh5Y6Ev2yF9wl5Cm
31PvJIARASB4sQryKRI7mygNqWshsa2Zxt+V43d6kCPwe/fZkSwD5DIzQQ/DD3Sg6EBgBdSadohO
zm7tEsF1bBabr65h5Gxu+80TJ7Sc8efCpM2T/E5cPoKM1PL9p8TrQMINZJZoll3QsT9Xmz6znFQc
C8w3j3MB6AM8JK+OR66awuYUQAMxQi/KijooTLCqpVQdgS3sgAXtyNnBsUFeSL2GSnBd71s3guTu
+Qqu+RwuMhEH13gOAPk7F43aVXD94WPVrsvnd+zMGZAuQ98lbeM8erWTH/FUqPMI5dM0Hc9CBVv2
DX3+rfFy0Wa7E1WHyN/+/EnxomkcQchp28etYOJWggsDsV1iLdsJRXBETM1Py7MNtwdoxMZvKyDm
pF0ZWgsPPwXwsSBnuxH83CPoyfyru+kPZULq1NptQPZMiwH+Gz43AlrPcu3+hEp434+fOFsH0Yjz
ULMiv5XO+VLmIc+G+cF5QTMB4WcDEtXRzY8msGCbFwU1VV2nyIHFXOLY7OGe2pn+tkGBahS9NEzX
83lS7RJenEPQSC6l+SNVizQowzhZiD1B3rh6dK7eCLyyFqALFR3pNbP+zdHQEJB8D/4KoTYOup80
RPPy/7ZW6pDN4fzRF1iYgrd4R3lWVtJWKedVc1mKeQZEz323DYJcJ+t46oXyV4AKui5VOf3Xieo4
386vnRdV90zge1U9DF1B6wvEKAQPesyT+wAFMXmGGhXHWTdcFuK0Te8dqOC9z0cBvkDAuuO6GyZG
+RCBHEemwVw0qaqVVUp3Ywl1UXSRo2CVRPjJ0u3r+nEAPNaStiMseA635hwNOCxoA+L7jZE6u2PB
ltqjoO2dmg5fQEz8Al0IxjiAMNRjqgNRNVruW3Zp+6YmzOATquAvSZk8bo5QN+cYcKX46SCXgTzE
1+51mjClv4NHh+lyESBKmHPEScPw8fSW8p+re6So0XEoQCwBWnFksOJXB6eJSmP7yf4LulxCrB41
ZDDdHipiHIeDbH/qzMNcJ605H9ucUAQurbz01UheoVnR0+VsOitERgHLhpKGovXcw7UYFnP3e+SE
6PGahsASTYNzZFRICUnBdx2rs/IAAGwezHRhkWrijF4J0vHG1fEoAqq/C/aWCTn21LnyNWvteT//
EHBTd8OTAg6bVKWGFyvkA0VNTgxqORjYmokQsCNv9AaHDgIyzrS64fnKmrTURm7U8U4/zVEfwDVC
GwT1bfuwIOeKbePjLs4A3ngoJoJq0SUemn00UsVB6PdcLb/dnzB6ruhoWYaJId9d11Ag+TsNrC4d
U6tI3fyqL3t+pe2zWZ3LnR07d8PsYV8ZK1Eas5XTKSiyuvLdkYbVCuR6Wvn/2mtYp/7mJIW9j/f1
swhbFWmzWkHT+Tvsp0vNTF5nCzZYcJvcObEJB1vyl99AqFkKJtdJSVpS2BDUCZc/Y10aQwazM2mk
HgKXbaMI0Y1ZialyTFFQwvChH4zDAjFWVkx98k24yomIIarXGsVjjxSIHLoVBlRtGzA24epZSywu
zKDuECchhL2zcvjkTvoOVGgKNTf5kCbMiZAAeqyxljYSbnl9FPwhB1TRL/8vTQC8E1in+XWoNrvA
Yqkewel2OrCDtNdmmnomhoDgGXH4x68JMnkgWPZszXwmCVQ2UJLm3nH5EVI1i42dYvmrdPpWLMP3
69noCFVIieC6N/dch7u/HlKxsOjqDg9tFu5U8alefOOu9WYg/falURL99UKyp5zMLK7bcjKQUdQL
+YaFu5go4lpbMBOoYETjH0kjF4VyIrEtTOT1h11mL8iEM3L4DH2mLW68KIbxDPLjKrx9+fBq/u7e
QFwPlOPPiULzsRzdOB2X+TmmiN4GGqHREjy+u/rVGiJ7llb89exk2Th0o8n4b/FzkhmZAne9BADR
ImXGy5XTXmDdhMoP4vGVa4Z13f7BCFjG988dAr4VWvJL17chvWVJOPY93x5HghseBFG9X50H7jYU
WEtUFeWFPd44cSMQUvrEVv6WuFkxbtVLkiyakZqa/+mSJA9zyBC5zeLGrugeLVRc4KJ55TlJasyo
B3g5nEyzyJKgyT0LF6xiLG24Hvv8caeDilqbf1RuuTmO2r8CoKjYdvjzYLbpb3s84SYK7zHv2LcE
kuC/0u03lWAokvXJnwCqYmlUfLKuCvcMXuP4+ZActU4QPXGVt51MuAAJteSZXYFeXVrG+h+0K4nV
0sqbTm6YsK26UvyOnodN6ndZyJQlFRl0ZkXvXECQOEA72NWssKhLEpJwgfywHqo82jPbdYXLYaVz
lPlzQzZf+UJGFOgQBaVsE4QgYcZr1UVEngRNiFZgk77KfbCfAUZ0imIw7MPCYe/XT8W/5ZiXnHfh
NHjIIK9r2SvpMT6vVEbwBjcLhe2XQEkZ8RMDmIsSL4bYYcr9++LLHtBy6ThS5LFyDfHVCPd2LCee
jufv6JhDn+seuCOkjJ5izxYfwBf7JQ4QfurqusLCiy/gcRrFq4qb2zAxMkRBzG4Xcs89p9EJ/OFz
bfavCkklrn9b4CoQkuoBDEE8txIQzY4ea5ZKKS57o8/0qfDl2Md1kOV2WeGXMbB6iv6sp7HhEKe3
mEOtbEqnklCtORd5fXJTKzCmX66ElyJ7Q0w8Qt5z1QS9j2Ozw7vWlZdfi1/poiuM3Q/zuIXNFRsc
zIEelj2l6fUjPZLDgF1EH9dYvReNxffplX4yqTrj3LyGm+4m+TdUZigqBtSPlgH89FmZEHoINf8m
279ZkF0dxAYInnSDEdypevNolse71PvjKT92iO5PZuElVwNXzGYX3+rnYcLkvBHbkiSL4h9BCmt4
640F5/Kdboc7WYr3W2NAjwZtFsZ7jwigw4Xzq53QCrb0sscsy5ZvovtwDfKWIjZkDtFXWZlCkuNj
1ABCD6TicWPIV5phWVQut9cRfxig4NgqkK+cTcdYcTCRhCu6dNuW6h7zJC8UN5cAmma9gzF15NFB
mcwMOz4bezYqj7GZfyGckevX1CnSoZPouuW1rkKP6Q0CdfBnRuYnllJQIUsy1vj4i2wMxqj/ifUv
058HHqOybREx7Ql/phmQW8J1zAasJRSyVPOjV4SG6oGBr5Eyv+/jgBWAsoPrv5ZoZ0fNs770ghja
iGGwMRGdlItjSFoq4KamNc/IE1WYpPshR1klfFAZGv0HFMCdHd/cUD0Jv3gfZ/MJiNB/ar3tQHrV
VnhcVuU4SzZgn1Ev/+RnVyCEhY8hKDCSvHqjmTdNal3T9aLzGZ6Abw2GXgYeZM9uWGvlR0u2qHy0
RwTMQtrfxzNDD0o7VnAM3tK/9sUyZabAkExA4qAjma0mprlCO8/WLRkpjAZRaYNgr/kI7ihZJFkc
U+pfn3LQZ5jK/wkUdQy3kSTK5R1JKmvP0b/gmnf4boy8UW1IBQkEl9wh3cvGvZu6g02SyPmjxPqx
evmLWIrmERT7Jbo8Ybj4kDAepK0Jv/lVx6WaeHFtr64DWUhmKVVFUYhMxAI9qnumEUeTSdUwrNSA
z23Mhl56WGAvGHgsF3h+0M0dLiTv0KO1doBz2GcBlBJ1SO1kYWXt8ebu12R4Z0/23AFR99B2VfB7
saTH6mnsWJ2kjH6uV1b7xnIGMHzV2XFgd0zJnTsom1RlFiSbmVf/QaHWRr5+j8GzFefKWO4xjXCj
f/0iP7BD/zTa/DreAoCrr223+RxxN0CbfbC7jM0MDSBpaNLUxcUh2NxOVOebmUwyioCn5XH1gBJ8
ZIeay6q6/N8uQxeg3vDQ1bYvCBqyMu69/eWiGtpFpc62qeTeF2Hk7F2J4xQTaCN63k8OWjTSRgm+
SEO6/XY/6EttXL+gKkhze4FTCMZdSHnhPwDRBcYhS058qFgKn3fO76CAOdTIdkPKBbFPXNNpNVEZ
bCrO7RSkvPcwh5PMzddajJpdHSJZqMdZp8S+tTK9S3QvzAnRxi8hjz8+90RjoJ9Q5kAtSWt3o3hi
nv5if6gn5fkJfinZKJNcCbDaz7rFiVOFFvkLkTOGdvxJGJh9ahWXwTXYut0RRygJ8bH5+bimoJPH
ajbEseqdUOjkW7SbYHCSLjzNEop1lKwkWEdTCoDGPMGSIE8ZnmfrcMT6ba1jdQbP1/VFdciR/Dbk
iT+gfHsdekwTHQ66Le1Ds708G7KinnBGm7ePAlmdgfgt/ug7pVjxpAKvA7V/afy/aiN+Fgm6NyGa
3AwMXY3uMD3kvT2eGi79eUUiQjeXyPz4jsCXWaDqWAHpExVGTAc/crT3y+vfMM8OqHx68oXibBRg
c/zt0VgkF2MPn2ei12Lx70pG4T3bEPdkY8ZjuFZcgDK9wfoVf3LM9+IKMBJJO6rGPpJcMaDZNdwF
7UPu1OMHR1jfEB0IdJdG8KtRphh4FuDDr0dIOKrkudH7UuxTr81eH/7j0H8w3hDwjLY0oFPy4QXq
Hwj7c4ZtJM+LYuLy3O09ECdYE6nI3AUwxoauxTl3KJbvsSmGoBmlqsp+OqojmDZufAGSIqa66baG
GANlBMRf9y1de8+X8liwO/IuVr/6Xi6Z4YOTP2jACb6grhq42U3zW6EDC9SWhIExvHvNW9S+BO9l
yYm/S6vefDnjuuWni0T2WpxB2Tfp4CFX6MfRklz4gMXivKHFBGUUdB+4JmINv33c4l23VRjjWMdF
aC5XsRQOOWnD71a7U/ElnpaqHCgagwbzMbOLZJn3XmBCwrL34heR1yNCciXE+FCkoxw+GH37pcgB
8thQViK8Tf9F0p6GB8V//7W+j90MrCyx2np2PlQNx1maq6can+XYZBg/2PtdMlUd2AqrWLmBU4pg
Zq8iY0YjZk+xx85CacUvUvlUUyWE1RqwZEBu9hsfWfAMp2JoF1+Ii2F0qv6Mci+IjvVPeJn+c1jE
nX5KJFSRs92Gmco82X/ZmPGyCzy50RsD+WjatQ7JRtn/GrdZRxNgtpMkbbWghtFJiUcNZgGuP0D5
mWZg1X2ifr0Kg7F1G6NOQJ5bxU1F/MHnha7kXXjAFk6hxz7cK68ClG8K6EEi5fVqxzAMj5vLiMDH
finyoQp0vz/4uAnczgwdvWytqq2oRw9v9NZSxesj+Xs0jlYWRjZfzSBXysWu6IwFniig7iUZQpKg
XJeBg+U+XL6Vq6RzX3KbRPEUbfTV3MwWEYBEsfsrBNmpSk+2CxjtzHL8QrkAaKJTSucTOv41G3bk
tHczVZqMN4iZEgUV1SRQTB59FAdqZaYuxxQHPy3i7HGY6IEhMtZHU0p9JhBdu/hukyzd72zu+8eY
iBGxvDUGJ0tmrH09A8KV0RDnvXFavg5nTy3TAbkCLLT0Y1EeUg1bEfCR8mZkQBPUuHHMVD7qIszL
IQ0P2RLUV6Ja8dF/UYX5Y8QeRIxBaI1g57FF8LRJRtB3SOFGdjhygU4Gb+WwfG5+sWxVgvPJalVL
SnVVu/ARvXdZutI9ax2JFtYNs30NDqVelONDsL8Ner+3q9E3Tf4FHugXgH0hpsCom7cT/EYyCDst
4W579aUdZS1T7x7lSGM/4fzrdmsB/CY/cDNutPd2lYS0IOkc9KBqWj09vNqBnxD2qfQ79HE1YpFF
EACVEvG4R5skNr/16ClPy1cN7+R6mk18tYOSJfAbihyAgAl6Q5BGe7R6rLkhZW5Tk09bcbYMlfDK
zWG8SAHWqBNUWBks9WFJGFnTFmPtCtuUm7dCRN4sUhYB56BXLrDCHV4XCT+lciIm6XlHIy2hjF1e
aBSFWLp0a/nEwL2kXR29ldDHW9hK1A==
`protect end_protected

