

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rLWvNa4xmaUmUmTsHaZZpmf+vdo1ZTZAwtQ7nnw7ufjv5GWZXhLdNQy5Q06lrQkoXFZkjYTdRiP3
F6m6R2KGJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hpohmRSyxraB2TfGOSuLyUSGGabJEMublC4fhU+HZ7LC068YGUgk2aE7EHkl1WtDE9Bb6v5v3Qg9
2I0FD8nMKFfSIsem6wrqx6FPpal5aJB28sq90dkao5/Iru4xYelKhv5oyEvq5w9fsErMuciA6N4Y
mVn0CtqFHil9PLQizOk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e2qQeTSxab1fevbjz90nhYXx0vSvMvWBAXsx6NPtcQGmGbeJ/S+FZG17TXPSmNs8pJl+7MKHcPRl
s4fPkRF2q+UUqzkqGrUfIOlc9iDcSV3G1jvuqC/KwL75+As0dV2zHDw3g6spyRgrF/QyMSev2EDX
wNjTOD0D7tDHqk1b7PsRTM/m5LabqbFbAoaZk3OIm0Vx4hjx1H+Kj+5LKlzym1OWRKYofd9Pxrcb
EMUCk84oHB+E99UNC1xkjUMB3ggxmGGz+tj2pQbz0ixGcWE5awa9i3czC6zJ21Sph72Xl+p+aRC5
JcGtcY8i/+JbJchaWispPX8x4NW4FjK9r8JxKw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vltTKSM8a/zRJ1QJ/9B9ijVL2/YbgBrtsRTG74WarkSfaW1TYFA90LAMjfijw4Dh6V3t9bzMVLiX
18WW94nb3vnRj+WAyEjiDaLRKxJmoyxgwsVe3baoS8c9YLsCvI4C+2FRQmKh6kD8j1o6xfJUhYAE
QHwYAw6Gh1Fc1rWYuMM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jeozeC2hZr+0l/LK5n/W7u82KI9P5tCxn4L5QInLhVBS1ZXkJv19EUcHMrHeYhgivoQ0MQ86TEXP
Iah9T/vQMV+h0mk/ZiG6XOYby7qUUR5Ipu6A3NdkCDCZw1M+w2At4X13RPUlLeERzh2uCLeznee9
UbtfGUHB0e0CGrBNEj1LzA1bbcGeOcLXMz/DrWLUmi+Iv7nTaL15UXhNNoh+XY7m46jwFf+dQiLA
SkppMG/4vt/EhyL+TyDlc4FcuyPEIIJCq1gQ6KO1U+4QL61Qp9FOEA7sAw8XZEnuD8uyPmi6wlXt
gqJWUq4qR9zExL8yZmy88nYYAn2YB3+3OVd4ug==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 123472)
`protect data_block
n7wXYgK0v8+Mt5IYLb1fv3zFX6Yh25lYNydkbl8l49wEqIbwnn5pYsdRppOXUM4KTkJyYe0JdoLe
v80H0UOnaAjYRMxI7RMqveJkcKJqzVP9vCVykN0z+2x64u0vn3kLvnvFA6Ae3StxRIF0rSON25LU
1RML/FoJvWtqnkg1A19rBWzMivABXhYtgg0ws9O+F7k28YYitYIOrerkeE2a/deFVjEaCmM8CQxa
GKKflUHw2Qmt20uXJgspKJJ+F09Wl3flsDu/I6X/dbDsU5S+ld7tJz3PBC2J1v8qjMMlueMayd1f
y4CLYQvF4f0SCfFbVl7ft8zU34YTS2Ekwt2GITiyBhOZTnZAK3hY4bKu1QyPVlsXrNfFB8ryV470
iNZvO8TeaEX7z7LDpbXSaYIGQrWT88t9kyE0PaN5DEB+a3uxKhYp+8gqM+m5xAfaj7ZS2nJy5Vha
rrhEYeaESHdSjB4WLgR8J9/1F6VZnh/BnfgLqbXdeRJOKRX4Qp2JoqymmkPEgIpk8Ac4kS/zrtxW
PpjHYFJgi3WB+kyE6MIYCxMzG4rwCQzT5DyAUoZ5BAABzCjtIy97ltv/wzfGh8DL+Wg/lNptQfbl
D8JayF8VY5F2MHtqJjcEKoSfOECpo9tp+K9PYCwaaBFVt/WS8wTj0zXc3Jdqkq5qve01wXaJmXw8
MmSpLF8Vj29wNQEkokbvR03Wft4DEBQfLPQGbdbZowiWansl+ndjwBH8l12NzzUgH9FI3u58f5Cx
WjZFtZly24VJNQpDS/dfv1rJvOKLWtNtqtWFjB+q+VPI1hxon0ylnXN3ESzjntIiriHeiD08R7sl
OgJbBPFyWDLfss5ymf6zrSVDiAe/VaVVTHTzXJMYNz2zssyT/abmIFX3Eh9Do285Br/ZqaqCM3u2
aHko3VD78AaJwmOjJQU2ZHcw0KrhVzAwtGkobfI4YohN40mgyQKusbokV0RfkUmddLvPgyTqQwYu
A34WNGK64y4linN9txDpIFGLa4vUXb5DMf+xH5byIvSji8hMWDpJPWSD/SP9qecIQ6b3rC7pn0sd
fgnU3xjZ4cYydxD2q9oXWudJc5s5xY2SMoBjtqlAfCQ52N2G3GREHGB0D11vdO/nt+bfIJMekSx8
Or7x793yy2osa2LmnoiLTGGMwf9VANcA66hLuLodM27R/FyQ4CwhujgkU9uvvLuKpWb2/mdJ30ik
uqy4etJQMislfqe1jBLjOQ/+E8b57IF3np75bnD3USiAxGjTKjKKt3tB1Q/kLubArtaGa/EYT+dd
BbEJ1ostz18pAK3hTi20/QG1jfNGhIRCRGy7ALmiMyA2HB9yQn2onEqJtCFnL9txLZssw2ABRaxL
2FVjqNX9llXXe4iewjdLt3UiRJ61rvzjNl8uskPlKfkGIpTS4wf+EqyMRXtA1bcewfIlsPJRiSmd
Z1cOY88+tmc65Ypdtp6tDtJkvBq3Benr925OOGLEmgF0QEja7UQPJPbby91JXvRPjKnKWx9nv3+R
+hpjcmMR7wbE0lMYTpMaOjOXdeMM5VdJAnKJv13+YncXAeew1YHz5VxdC/nPnQ/rQGgBn/YaQh5m
PuD9CLe5rG+DO2CyAZ4hnRsNaGFxdZWq4chgdAaL1mQBk/jnQP/2ffYlJg/I4yPrESpKBp/CSuE9
+RVs2BYW4MwoY/TetUY9N4a97W2jP4JKQ4ZkHlIe0PRDdC/LsQ784eadm6KgKwH1CuehyFVZtReC
o0XHlay1qZ4vrmCRPZawdcPeq7ech916TrYkJ0Pq+CrjqOrwMdYsut6qArx9uGFedkhscy+dI7uu
K02WsObZRG82KW+2uxPFF9Udq5t486ttFAIVnUrQueMDrC+HJD/YJNCoP5/iFDohWvKg2hFe6Iz6
OSBmeTXLgPIymZdWUiCpD5OtL/SGXjK+wwJFrF9XieCSncIeWsGeUQGE5sfBGvQXNtak5zFHF1aG
8fI0Xkjkz+pk2Mt+Z/J/megvpBFH1KIp2m0IA1zQfQADU9XM15EqtWywOXjs2PhBORMIB0FIAk+W
sSPBHnrr4xto0nvkPzXvIa6z3Q9QqsxXQ123NkwJ3suFhbtVThy5H0N7Se05eZdJIbMHz9Ihw8Eg
gIbTehDSC1Ra23HMY1IqxBWDoDI5sSCGmyu83KzopaornS8zDkPXXFDdcBoeFw19HGB85utyG1Qz
W1P+JvkL5WWnV0TcU2TqHgrloM7c+zxWtxcvd4eMc6dkXXIqNUxkRQsJHYpryxUVoqT/u/PIsjNg
gLtIj1DAtEEsDdZoe/43Aiic27T3TMfZD8euFgBTS6X67XGJb+SgNhZporB4szRTVNqtHE/uu1Jq
pmnEcaKfXnA7nwE7Ax5OVyASJtrCThoDcj9TWNHnAP6oI5sRbaSNnn1t0W3i3AtULso2TMNkECeI
O3hgAQ3SQLewGYdT30okPHKMMGMGnsP+YDjKTlgGLk6giSIOy6TuEOl2K1OMwIkcoW6W7EQDhPUT
/+BGTmoZZL+gnXEfwoiYLFaxt8Ut+9pxofGYYSlLUnRrYdpxfIWafNUGV4aHkYnEFSx9JbNUeHKO
okf93QSiqbpt5f8ZiG54jXtWyuep/yBaHfaJq/3cXdarpT0T1S3OaUlRBZqQfMe628W2u7NMDL3Z
Ijr9dK8NnHEvx8qw4wcp0M5SAI3TIpC6Pedwv4ThDKsoMKxmOf4HrUjyWrWCZIeW/EUoFNT+RnLO
5zdFVa3KKtFZHpSwR4xEVzYiICm00I2nZGyygavspLGoZ61kfmuNZep8Yj7s7+c66vMsy/8/4TJN
IgdQxzaOxzFFZueMhWxj2wXQDvWejA1U2W7gmP7XU1aB6g0NqGor38MKK8pP9y/zQksUkdrAC/ZM
sl1x1UMaOFUYy83n3/s80fbCC1k84Ig6HOxQIqqiBwX7Z4oYXe1olxjMHhMTwO1RmVepvFbguZbM
tjk0WXBozBExeMZn15xPRO2DCn2VyBa365t++tonsi0TkVW3vzscx4g+YFLo5phOa4FRAuNPI1lJ
s8xxocZeIU5Emjp2jd+5vADXOMsUwu3tXdAtEfoK2sjsnIl/Jjv5sPW+0G7xwkKPRJdrYqeBdVo6
U3qjUx/UFZBay4p1aXWAoDA+HEND6/gTDN88yid7hh2sAhViSGBIJFougrrh5dlq0AdFr9QFuny+
euZYGp/n8R/TDWHEwTnKl0Wa/7otxoT52mtnTSeL57iABx8PAu9SFfRY5SEBQQGOt6YHXOjO/weB
1I2dCjjaFEbJMVKargE806MpMgq6xufZUSD7FK2Q+tyOPpVbiCCmu3L1IbcmyajpkIo0Uiw3UmSx
sSXjuzqHbouioH+5WfVd8jrQXMbNzp3Lc9t6Mlccw1cvwTdcJAlteSh8kfg19BlMh51ksolmBUQA
Ob8+dWnD0kdPjCYTGLg0hTp/68tcwRcjyyhfhh/qrs8AO7RcpIujpVoDxXJ86bKaJMf21XV/ykwH
awwgjz2jpV80SO0qmIANFZfACvQQnmUc/OfGyKcWktziq/SZhMTHgk5SpjXMczdxS6UtKm4KDwX3
IpWUZkY62fAm/bZEa9RrDi23PiU8a6l0Pi67kI2csxRzv5GsQNKzRuKe36F0hzbZbycHUPm6qusy
btBNAzTPYuBfVFqhbMSY5NygbVjaXuKVFiJFUXzWPbt73rSuvzQlHxAUBFSuW1xdHcxXMcPN8Cyu
I8vkpH78dj0OFRSzeFNUYIFrJ9YuyN5YA2I2NdZVIAkSRwFttLrdrlCR0os7ZDsDKLYpC5mSoms2
HJrv7vxmOBG6ozqp1V44ixBNbksWjsThS6ej5AFZ+nMcK9Ww3kQcufZGrkfqO1FTIIIToIupH5ms
qQObQ3D6J5CU8z8GClB5L1oMeXwPe8o0F6EVIjYT3Ipr4ryFLY+AsuPS+zbrYVYpobPyxkpfhtrX
oppX1DemhovrtN5Ic0usq0aoTIipNvYi0s6VQesI97Y4e+4wACEo6BXFoS8q/UbgmC4FrM7BYR4Y
pF4ZRwqesIKljXr1RQ31g+0DQWfh/G4a4R0UHoVt643+dbln0hA9Rv1mJDmbO3AULnXlQ17QX2fC
CRUqWIjdWsAxSzaqQ65youcWzO2QOVd6RgEPI4NrDkYEZh0v4v2E/y6rIM9GGstNR6Zt2/Q0bgPu
Jxh80yuGVlVSs9zrB7JRaOALfCxgV9PVIlmp/naWLgoF+qL0QM8z2NjFbENqGT5lh12CdbCT076x
NVW7PDOEcCGJ26hTik7lYS9Z3ThIX9HMxaLuuUdZtzkDmkDgAjLPAFV32SKlT0NYk2jCBXQLzg4L
OQYUquYv5nRjwafHT09dSqjw53ZF27fPWeDYzAVkLMwLwkBfIEI3G+j90oDxzl4Ar1YqDx1FWE1G
swBRruh3aEuJd1YOJdcsfH3AsmrqsjR9rphO5/kuZSUYgpRl0pzGnx0hrtVM0nuCcsyq9kvAxte6
RGMJunN+5AykGsomM+IrG6MRUh5ssO6C1GPusLIIhjS9OtzHjoKHClcWNo3AelAhevQ/kcbG82oA
abaDAQpkXYGWBJQVZ6W87AiI4OVzaOhS0SPET3gr5h3XEccP2pkHVN/PQCfTlLFRpm4RLeuOmRtg
AjDXXYgSDHQ27eClhkg2ScOdhR6Wv7zpOUkHMDqEiBhuIq29MXBuoEh8/v9qgzLSzwqhWLLk2Cy4
djLRyJIsM+B4FSFC/QKTnoloP5F3ZpRhyO53MwUXT5/yLckA87hml2CIgffJSwt0rsFKmUy10oY2
TxfWp5DHrxrQODENBX8RFGhbZtxiE+OKE8r69LJ6h8ZFrGfDkhnLo/+w8SrfdYw4ismeoJlpxOP3
e0gn1pm28lCk48AzhJPEdpDtRxnWaGQre5ebgZdXw4U0ZBpMdu5+7Rx6nOp1lipkEdv7uhHervSe
0fp0m4AVMX6Npy5Lp80tgPIKJbYB6/H7SGbrlhs0v73hOhE1vpRjKsQa/5lmxEkrDXT5jNUXLyeN
NnN8FTwr9m+Qn7S6mRLZ9GWadVqGWQLbtSyXmbGKrnXdCyYcgeecQMbENCmY6b6mu3PXQPP3HlgE
3sKVVZ3aOIstGRhZpE441GhuMEOHyjhq9TlaKa72zAXFeUbcM/dqhDpKXo3VsvpCqMm5hG5Ux552
6oiYLzWqZLHww11KBfSOUmlvQiaV3Z9zIhUZ6G3LsGp54UyGi42FcYQwrZ3fnr0fEEcKZJKyu/SP
GkZl/Co/YoxCCmupJ6bJvH0U6xN1D0AjXV7buQcD7tDDzd3IJkjmEwvWqV/9muA40CQQAm5OqhiK
eewYOWwTXBEkEo8mAeHegywxuj6j6t7LSBWQ3cAYLMgRypvNepT5I9arPXGCB7eAw28YY8jg93iv
JjmmGEdC8aHQEA5b9Dy20XPGjcCzhSK/967elOzuM16Xp+DZgGi7gtUQEpRZxbTWg0o4FMyvtFlh
nIvSf9oedlskHXdoek7lPEpyas/E6Z7cJ3lN1ZiQWTGKa7htz7OGmIQxYk/WpblECLReqKGNMyR/
hn7XKB7bzKSN0XygL2HxW8nJ2JTCKfgnTGsU1IXdYNTdxBl6OHG70LqU/qLabZVVNS2LQCxLx+09
wqPjLqQlc4ZoyJ6qavbcNnwi2ybCMcMhO3BbwrUkl13/QV30C9jYlF8RjO3t8kEzSIsfCo0MKmt+
2WWESKMaLzcgDh9EGlKqwNP13SQ53Up7gcOtyAz5SECz+gr4Q36XI7Gn6sRLGwFCMf3dFh4sBvFi
O+4sPEP9ZgAJndH++hCrVN87eQY+w0rDt5lGiIL/nv/gx6m3KXp+TzZvC9F5OZSwPOeY4tz25OHb
dVV4GushMpdmEwP6ee+3egLdqbV54J83+LAQRo+wwtVKDLMYsoemk0LIWqR9awMKAKUVR/TRTSCh
CDN0CWDeyXUBF0SBoqA6WB/8pDUUGxuXEHyHXBHwx4nM2GYQylKuj+t9uOd4/IQ/iSZAWUkdnshQ
t6KRBwiXGwDri5O6s1B+x957Pduk1Xwh1AHJBORvUHJdDwMea8rFxou3WvKIvpXh7HrGVeeHyCBS
IuRyIUz0EFYZB2iewGepM2UDVDirEQ92RcJ73DDaU0GldgCKYwmXQLh350h7UdZyRYmH2rHGPXoH
qhAWHQNYCP4fGSg3zHDDi5Sby2uiYli35eiuB2ppLlvUMHreg2FGTnb1202W9YvD1u69HRaohWGz
Tze2XX47Dlz6Gv/j710NehyLosSlkMUepc74shwX85K3XVNnPKCFzhbMCYiWuFrOmGbEuhBKyHbk
f4IlFN1oiSEvTgumR8uipYrJ/xrN/Z3mkoPhVmjmtQdABIwfqNQ07KadExZqi7aAxGnnM2eQ9XDR
NXM44HX5QOcnITgRkDrFDTirPgVlw8Q0bjZxDdNjFWo2TW2dKlNoAr71Pw5QRPfaigtgn7kvcd8h
OR5S+NrxNvutqdD+gpswidmnYeRVKot9KtzmSR9cAFTcLDEObzcX0PXPDXp4ZCKpTS80NdIFZOaz
NfxyVUKeZQIeb8dKzFnAOqcDY+GD1BmtnnlnKVi6nFYHcR3xx/ikxZYNQYhg27LxPf7fb08cNUkY
YcUSxh6l1XrTLR3DNl8b3/1qEkNDJlMh8Cs4mkI48j3fcxxH69JQHC4zhqpPAJSJeVz9OwvZkD1i
6/6eDUS1lmM987bXMtgZFKXEyQYYvbB9LSvKqoW5ueA3gZEifDzz8gNnSL7xxLx+OX7n/b27LAAy
anzGjHZuKZpZPtA0yM2kIWVqaxIKmqe9cIIQYMGEs1l7lXBZpMiLFxhS7IsxxdL4x0Lw4UHgFuhl
jZ4NtcN3vx6hP5c2h3jmJXfxVd6VPckoJJ5P8F2aF2X+iQP3xoyoVOJ8768r8sy3wWfwlZoSnNqR
eQJQr6gnCgYbl+hCKRvv+PWXd74mCx1jzkUDqqR6mbTeT9LurH3O38S49FI4WeuYgpF5KtabyVyD
9Iq7g58WPDAEzhOsnHFCvkgku6M5BRb62XRStqZYgjsxAhgSmqgWCaC2+Mm1VAcD9Oah4q69urP9
MW2jNXGECRf46qx7H0/Ftq5OXacG/vMKw8H8DEdClZqqTyOntay0y3aQcGRy/66fTQIWBZVqX7ig
21JCtjcUD+92xq/jGHPDQQzERbBpJ4HO96V1Xdl34wBDGFzvAtQ59+GOaZwtc7SY0pD6plImFm5K
wtbvVq7tLnXzy3UU32jafVVgWIzES3a6xEROJlBYrhJcyiaDiIcxbkzdRzPPccF/AGlgdg9PdNuG
Ii9sd0JIcYX+80EaMjSkkL6hxbbg5EL4Wcrfyi/qgU2h6+A1oe8qygMU/Y6DfgJQRiBaOFVeg+YF
nsQ322g/NcebypSpMOVt6qVf5oZ/w4uYIAthW08pd4+QvMU53hqVXvgQEaog5SaE/MIDAIfL+u8L
6OgGaJqyNhU03mEleDGz1Kc+L+1O79RbHgh8SlQ21d1ppHqBxyUvETLYwvYif3RqZBBAK/55ylUq
s4yakVyNAB0zno3+7F7GummlYwp+4H18x4FWOVXMH9f5uyHat4ObaOPaqQ5dgMP66KqlUTxLcuwT
c71GknfdXmOBMkginlV4+yIK5wxIfwYWBURYZ7wVjIeuUgVYrXLvGzYIOI3PYyG82f2wr340J7hv
IJFvG6vKYlvzVfq3BJ0OuRTOi6p+73YvYJpR8goAsAWj2rLKQ+EWRvPXsa7v/5VZzZMF4WMRGD4K
L4EgYD3kl1njtrIaJO4vhP3DQzTd3VXj0WDK/HCkXSzIdJnaiv/AQA2EQ5JHtEhFpBjpGbwqNJdI
8ZxUxa4ucSiufuhcv9qBWMTwKv9sY7wb/fHcX9gmfumu5S4BnTvBdu2TXCCu6pH+6buKGY9K8hhT
pGICErI2xRbynNogBMVge3VFiz1y+uNVWIBbR7D03F1g6ZcxFBioSoqImbCc8paCitwoKzCGW8zf
A0jXI/HkejgPoT9M/0NRdb4XRTCX/M6GW9BG5KDscqaqYA4GMmrSUmObqURG9864v4snkxW7Q3ev
Wq3W+vipMNy7fg8c8cTSZA2X5XXfGnzI6tRFTtswdQYIxvK9SNGvLFsnWDK8jpZCK4u1nN2cu+vX
xnxT7g6Ip+T/gT0bTeuB5RhRa7Qhe893GX20D+AFQKoBi5YipVI6nw90H6wHTfgcmkip8/P8NA01
ehnkWYISM/J/5Co2dCs0j4PTeiROws3b7kxqFFRKZ7r95++apKPjHOMi/+QwHXQpgeGj3piuMrBk
fNndLbgpg8fThUtkbOgf9sPSRteN/BnXznt6QhTPXZz4u6qGw4GTrw3GRmxZjV7/vV/OdaxPeaNX
88nl/nYRAPtKLGDg8GjYDSV2D/6duTVSi5G9HOCz959laUJIVam5zR1m6Kd0/3ePK6fRqrHnzAyz
KvTkvXk3lt3KDO/ftebPYtHFVPh1wwAyNrluFsG9B6LuW/jR3ly66DKwhrLjAzCn1CHiel16ra68
WKnpSnkzIOAGrz0LLBvops3AWOntq+NeqY4sRbu/M6u0rkwhK5e1Zz7qM5e8PYHaFcpdHkR7J/gx
BJaNs45yiwn4H9ywPRW1cymmBqwLCvwvtehMeEvbx9mB2btmY/p3fJ5xyHq8CtihLzEWaUXLVU+A
QhxnrtcEUEBFD0mRAwLeRADv4OfhIMiU5JppLKlTGh4z3kJ4UyqvV965lGQnAztjcVaV5MkjslLA
dc3krBquUZsbVYJYltJU/JB6URdwUyuB1//a1uhYxj3zXfMbl3z6nf0uhbdip38ZVTgKe/o1qhmj
WQ2aVNj7sXeh9+sIBi/YFkI6DzMOqIEk1cQ2DuXHgNtuvFn3FqYM6+mAmTjA4HspCpjEl1IuUKjH
bHgJ99xS0Atsxxr1jlKCkzH+YMKiXCRnhbjM9eS1XXfVCTWAAsLcfHgjwfn/VICXtW8OrorboLPl
u5J74555jKhu165ZWr4HRd3Z6xxSESm7wBX31tZuIvO4INHkTODFOtanchh8wxDHwMep1oXyAVPi
6WFmTxUJo62vNjDR0b3fAn9SROKwStUqyX8uhM5Buz7MkbSFE98t0n7IJQ9qUNSrC+eU6sOM7cv2
ybzLhsFl8AHdmgf93xl8dOiY1Q9L8IxBkOU87pgXa7naGeLTiYIiWX7iEN1pWXj70vmWZQ8WfK7m
OV/1DzA7fUmKcyPPMLkllqHjtEdAlNNqYcufyXIHm/cgfLSPdTkff5A+5FIU7B+XrepgY+HDUsNO
s4BdQ1k5SYZ1AvfwPMEv/uCKXFlEIFi7ZY/wONSsy+n1I4aekZjM2r2IVu3KUhi6GsuSnhsKU+2L
FGZJFIYBxZ1UMoR2L6MTSXtqWvLhVV/O3jJGhJiGeBl1K9vvbheykO+pVO1CXsiTiG7SnsJfvkFs
X6tw0Uc3hN4mWXAoRWuqezfMw/jx+BrVywDItL0+7GWe513bx5DkJHz1Vuk/25aCrvQM/wgnBxkg
7Z/lijuMn/8Nvu3riENwsCKMDYmt/5mFtb/B0foqgyhcyvNBlSl5d4pATO/cQbqH27S8YNNPO52a
aPYfgpB4r7EQU7oJBxEuxC6k25g/nOQzoTV+FnZywArY+DonhmF74+Cy76EsGgnquGExIAdDBlHt
5PTP5TT+bpHeKOtm6eh7hieOjGMZJmvNqY2uIjc7BSx7xBHbnGN6XyulrHVFl1aysmNYoLf8271l
MIwSx1qf5Pd9l3rjFZZWhqUqJtY1XliJGon7gj76rIgZrKycG4RC8C9nANZTvK2ox1x8eTvwEzEA
CjJ8hs8/yCaE9hNyDYZiWEbeIjeb+0VtgHqsgAJz7l6uLacANPYz7VmrlwyWaHHrHoKv1v1dgcAE
IUsCuDJb23YRieaL40tBYCQ2TJrGr2IydZUUzdM9yF0yuInDvSlHPB2iQ/YHrdlv0ptlVMLRRGSB
8QKCzFX9F/WqVtKa7RjNk2o80xtgHJp6ZRWOab4hlTcT1zciJNZAyO51WBjnXTty0/p7mgSY/6e/
46RsmQTMiKae/j7EnjBAc/V+eBJM4s+nwmC9NH8mKtW8VDua933IhoepHsrTuQQgq5PAfs01ZRzL
3zSjkw5L+rZz8OblsQRac0Zc2nYa/tYLfNB/7+NNLfa2ARC2aT2bWc07dMRHOpdux+CyKSWzKbn4
nZ1EFE1FPBZ+igNB+HCW45BHpbtDcqzQ/3AxeNss90zFFMi+MAx+xwk4gTISCyffpjH+l9ReP00E
M8IH44VWQw6cI7S/hhoFEadFf/h6JkwcSrG7Znc2p80QTWD66SXRij4vYANEq2DwdvbE9FMeckWK
siOP5we2VjZ6uA7BhNt5dHac/byzuomLTBmgEMVA3Ay6vTpTIeb3X35pq1BQYVv3IZ+wMLU1jV/8
ogMM5MftkJqe/nqovQzJdp++j47xBg0E/x2i6SJ9mE98iqKDL8YekpdNDuaumSJvkINdGsW+8mX2
LESozklo5HzA5uav36lIVltOG9Z/NeZw3e9oEc+qTMCLwV03FpRGBxovhnV6gtay/+WE1F/vxETg
PaTzFlXuHZzjN/FThqwS1lKnX/HlNDp+DZF4o3oPN/x1Ccch0PuxAKyJH/q3XnWWVXeSxc2+r9DD
6M5w5F0vHopyxSXrbjiKBTd1/x9N/5kbmaIPQTr7q4B/YWRLR4lTx6p48bdNiOIU95ZnFAiVDM/N
BeBuMqsbemxKrMafoXx26erfn4aAdg+ruR7lcsB5AtFhuQ2QP1SLY0zTlGyhq6LPdUMw07mabvIi
bKlkoapqP6AdJ7/SXpe4F3Ih/PzuYe6ToLbIn2+YX7KgU4sUZlNsD57iVWP/0qysI6qRUbbcl79b
AvlilYFb6jE+KhOwu0MQP0qCxfJuRroROSvg98xEcomBtdDNLpOM4xK/WZKI+IffZ4nLWJchheek
5ta7+tgjouBz0KjLGfXcej4q4kxzUfC41OiBVzK3x42wiGiO1Rd9QKWmADUOZov0rlru/NVxZtj5
b9ZZOSCCCHui1o89bBIn0SQDscV4wYQ9ev4Bd/8OQYO2e7YXiKvPdqMabYiuhgzSqsZGIRlRRoGP
ANArJYwtUJZxjpJJyYcnhb3I9fw7Lpxiw+HSUG4LB+FghWIeGPfWun3mBhf1hv190GUbZ4vNuvkD
BIvoKBvs8vt3VA/WdP4hw950EkbTnM1XHXk07+StFQZfy02yJxBbwwTydIgU1YwayGwipmWyvJMw
wQhFGRuHwS+1fVwv6Va1C8w1R3cKz8Vc4PAqDEg1fvBZ3y2TMF5m7ewNpshje6fHD53fVecoQOyk
j3KqpE03eXD0ErVflCJ5L/BhhYwlfKRIJFVvNnDYiNKj6/imQTclhkRjV4iHXMQWPEaqgN+a8YsI
ymrs66+4K5H91/yYgUeqq9m2bqz/1qwtmRDGA0SZnup5dtBLkAOqTZtaSauTvi5uD6vAFR3fpVMc
Nk26OJpy3to+09bPHX26Lqdus2rPGMQQKJjkuuwm8bYF7QsAJW4Z9KJJX/IZWCCR6b81WXDET4V3
B/AuStXZaANswDeCmnly6KBDEfyHCxH20oYhd4x66G45mRW18LjhcFlpi0jxhi0TI3+LTKkSc/kZ
i6czI16lSoRUushDlvnYKq72k+2yB2C2wC33SAeEVR89huYE3oB43JmAyEzH/tqMQ/7u5wNETmiK
hd89VUnNgjAy3AuMpkRC0nm1VPgbsFJ4CAy9DGrZ6cAn0NdutFH4wzCogwySPXNPHS25iTVux0KB
X8FtGy8rwQ/nbb+LN7p7BmNZEW+VPKZ2SiLzHC8Rjg/fWAb1lW5a7OrpK2BX7LJGCxeFaXzZ0a/6
XrQcJV7rPrG6v+po+IYIBovBHQl9HULpQJD71glAhQmv4wNxc0Df7FmQp+7UOwXu1mFa5KW3ut+l
1W0xEoWgA3vjplY4jhENa5Xtbr4DNy53MHNYSbQQa1rkOQDCsv9dkNhzZTqipgKv8v46j9Rwkd3Y
ryWgSNEvTF8/AEOitO74Zb8Pc6d9Czisc4u6GcXU6BB4cLYj2mMdBp4YboxjSdErMmSoh/Ch2xJB
YjixU0LPhMZHv5459AfjBpoCfr6wns4cedFmtQOrDKM9L2+skzX7Wwpitra5J1/zl0A9CbDCZhai
wxXb6do3Vqryt/epzdeDDihHgLqqoCeqMyVQr3BXHsyvtstHwfXL0yOX75neu4W6GIITiyS01lJ6
/aaCEOPIYjVBLtKU7b1cmy2o0JiwzbQFa8o1OsKw56545gbjj4x2hlQMV+nvJkNgCcTdJReTCQ0y
7mLpI6c0TsvYfA3/Vm2yJ8zS+WvU+SeC2FgO7XJymVxEl3/TpqWkKx9pzZEqSP5p7ethxqpSEy8D
qj4+kxSomjqdJbPsoalLOV2Q1k9jPhIvm6YmSKrtvDBK3jUmIAEaG1yDFdxvoyvo8sPnGTkCDcdX
DNQpF9BCP08aIy9pAL02116nr947Wq1FuQJUx0EVEI182j8p+Je4oooWaL/jQknsEVObmvsDXdUg
kHa0uluKIjYTnwBP82RuTq0Cjj3s9eECP9awBE6tCdFqbLoTkGgdSitbP12ucPJWwtiqg9nzql1Y
ny7LyWn9CAsSHO5fDpHRFduzppSciu1g4j91riZ+85sJfxknz/1hRv/MGmJkWx4GDiGMyvSS/WWu
Xf/EEHrvHs0HJ47rentVGJWypRx14n1HDvPTca+FQ/N3H/21RP8GiGnd/SHcWglJgKErjbhlFoG+
1kg+WxhOKnD293PfMdR/eRb0XKGbY5m1wO6CNQ190A5F31lfkg+qY7eRk7KJyIySpA5oUOOdcEPt
CzXBysfn3+JwZxo2QJKJaXPdIOuN5jT839zbdS/OPL/op2sw1lNPxDhUw9LW1RbBprcUDIyKAhIK
UcLs1FSMFA/DtNwKwQcaOj7DTkEjt/P3/jT1080I6RU8w0S+h3PGe+IE2EZQS59WNH0geoYHO6Bp
7mBalEw7hdx3wORpfKl9Fg8oXP/Qa+hYnfxnrVW6wYknI/GSfUNSaB603j0zweWlC6pexSUyz9nG
vMnNjnDeU1vOsly1x4t34TpU9l+XggwCodRTUM7+ukscPLoFScMyV7yHjQL/M5bmY0+cNIX68uHz
+7nKIg5U5fWibzio7J3LoTNRw9aNsc67xaSbwQY5kh6dXOIzljdcqOH+0xhIRCbzhjHRPdj3Mvwx
6YlMaLrsqFmDjISjeoS+ThW7WA2nwy1U+4umdUBD1TctfgPtHlh+CFR2y1pjfOh+HaUuGofZDAlm
2E8ZwKYywksdShDr6ZB08m98BiGpWIaUhhTXTEixyXHHNx+fqMtDn/TX5WSkojeK+VwZYMMNtH44
9QfW5HGpF+aCP3nGB5nmZf2Oy05XtmO+g70spsSLGg+RoWg5/Csf8/9CdPAhT1biMOFjT6XJ+lGF
dVkj/hKNuoOH2XLEUR7PQlWqjpsAerXzFuQfOnuaS5HQ5mB0Dv/U6o7PXCKocKTAHsEbqaPDWYJV
Po00mSeGZt2iXd3G3F64AERqYg8pEhdH/wk1ZiKmdDx5KrIEE/RPNWagDHt7aoOn6L0y296RwEdU
c250w+DkOqO93ADd+5VgC6oZlu3l2YF5BufQBqSckuWUmmx1SpypukE8P1TOiGmzfrUFTfthtswg
VcIxJ6cXlPGEMj/e0OUjJjuKsj395eJNtJrtTivEMDyUu+ZQsvk7McT7D64Uci/fru+LuYhYId8l
UFcoPddEISrpwl7iGMPogxgQAwG4hqopbBB0NPZGY4hGnqQ74xynaTAT1T1n1i5FldlJCc5LB16H
re05g77fecxtOMqkKp8Dz4NsPEjIc6rwdHXW+x0NO3jxj+CFpjGkuGpG88anZNoUWgGV0j9qJmCd
C9Y17h7H9i4YIT26xA6xUyNyCS0D1/X2KwoqRqUUxntsmGLPBlM6MVADFW0na30yLwjC9bg5W3c2
Dz9CAfV+k9hbcZO64lfQHROvXiERE8WZFad2atANJwTATVpXRwKoyg6xsk7BEUee+ruXt/MkKP7S
jdYYPPjUh5oR1Xhq9wF030TKYq7mbUmNHsM/V/ms5tIDIfHwP/xWtmwgVBZCOHMC7gDFO6y2ek9R
cc8X4NIlJlOa/KDjR0Nl0YC1MsDOtbx63ssw1wMraM4r9Pqg9BIfLzoV6cLc1Br0SFxMR8yGE2nv
bPCPkQxw8RkfPvMBkJnq0Y/WsBRbPbuHDRLODp34Pc/Nhdscvv3mvUZe9mGmttxGs7JgfjTnv59r
2AezMDkKs+kdkZPz0qGIICkPhgdkTbCL3YdCcvT74I7i4xlBKdzmefN0GIiWcLpTMCBpnHCzGdZK
7zfXr+TNhYqMsqhcP//xD+29VCFu8GdXk/+K+aad1bYR3XSkfhIi9cmFb2+yRSSAXSdfHR7/tXfK
YIF+q/MBVKvNfdmETZw8mctM2msC35YLPGiGv48AtFeVhhKWMp1pLhoJ7wJs/h3O3HLaxyeaSq6D
uKyonwA9I/AgHgr/3iR7BpazGz3Omf9CMuWeNCmDH8TY8cH+W8pquhu5e3i4rFLwzC50ExJ7UYC/
Qwdub0Ae4DD6mPsvKA6lNpdapPYdK3WsHx/ZzY6lIs5azIuVX4W3nwlvfaAJSI320uJCupSzMkE8
Ri6LVZ+f/FNmPrS7SgtWZIr4FRhHPq3FNUbWHqEY0H/yoRDIBCUhZotBk/cmlD/9OWUsyOI6Bhna
Ci/QL7z6Qs6YtFy+WHJGyB8RSRsVdA55+L7ORq11h3Xq1SmY1aRhnFUPE0LagMr9AD7dX75tw+7i
i6NhSsW3a4spAS6HUZAJJtSJ1hj8WQeUfb5QwIcJCx5fEyu1bQtj1Mj9I2+iBCVbr6VIWGkuKDut
ukz4YCwtaEpjgk68svhInwGyXePTGRljagKhpXlrV9GdJyW2kHuH6zE0EDnZmAVl/wDj2qSp7+yd
/B4PBW91Uii0zf6V6Fw3ZK6u6ruPG7QqWG3NAML3fV7vaXZoWEWDr3p2OtgofaRgcLihH1J1I9gQ
SYtjJeAeuEvB01NZxI4fcCvpVrUHOjqqtGGxL2rTltCDMQ+W7RZT+OecHH/AhlN+GZGctX8bKFJC
vcxrxtjwjA5mK/bcIcfHrpap3lgZSE1fD98Cm7xfN8vCoYXPC60MPnSt+Rh/yXOz+/lUT5Qg8q+Q
cvRcc4L37HLhNAUb8hmN1b0zFpG7ZsvqMeRelhjX9/WtnVuPZMMWz1NQhKUmnpwCaVKEB9kHAlUN
51zKMuPDIBgyC641PS0m6e4Bo88273GcEGdMLojhL5sALpr3N0sjFXwgeJwZVwQJ2SpusiZJY4zf
hrzDWd5k+H2FTtEWzg9jB4RNEPKEZUUbLA9zn02G09QMZbdNt5Z/YG/DxOq45zvsUJN4UvrudrR4
3CwhEWs1rxnQsYHcNi0qmwPrIhGR6AyMowl59OPzmFeVnuDbUbCVhbOmPsplPG9k4Bi6bUU2jQXZ
t+1ujHTSy3ofkKQpGTYRhdEcVLRtuEi8M4MKEwvzDi74nfWPfZh/8WUHo6JXCQ+X9tZDDaM626my
qVa95cSDhfPKpi/yZ9LLpCl1icnrcFLkWn+NZdPvlH0XvC0Mu0VfczWcn+OGkju5NY3OU9y1FkIO
M/nt/hw+1xCqSH+0WhCAJB4sGATrVkMP0IVqSkAtBzi75qP+AnFCHJyn2KxcZV/s7peszZ3GJRmu
LV3+NHjsffJpK+k2bJUp7oOXQ5dIsYDsU92ibuVLBmu/ULRrhQ2eiwUiEB7bprfVxMrYGZLbHYS/
vqzeiXsQ8bXDEsF75bJuXcuWEPR7TDKc80WfwQl/hOh+KVQ3vimZ/3XTJHt7UUIxs56fAwYf9FPf
9w/aTTLvZgc8n/qPKxIkUVjazxPD8/KVe371d7vfDWmKllzWSplKwqIxlAX5w1/FqUA/Y+tq26jE
zzpoC1Sk0UISRta5c0aCbhrJ0DNdCjab0Sc8sFjzElab0r7iYYSxAZTQnE0ABHsS7jpUXsvg43UQ
WDOG7hvtuykWjdSN85xaGFjAIg4SUEE0hrnT6Bw//JxAIlB9ztqd7WoCWpBvkMlaNFhu/ANNlOL3
0mdfs7VY9MU3zLToxZZDqO9957/E1yki9Mnx9dvGsoIxcfJGdxnpEBG+v4I2QKBthZLiTdxB92fz
rXlmjB0nbYXRk5xtI3gCk2hNyVqDMzPrrHCLRcvqET4eRSs0pEazWLBffjq2TksmYgNNPzf9oh9+
IKJZRrR3thDw8SmYt6REz1C6NeuClmsuFd+ALB0S0BHs4f5TUlkC6tTcmlyZjbDhkvDKAO42ko1L
HAc+im81Rrb5BoZd6H7gSLbYAER1/tc3lUt/jlhMVKpcjbDIWnV/Es27rCyq9eqD/NIscJIjqCHh
N0PBSZqmr/NeEODO0sw3EwOuXsyH9t99WWr50CfaGDRiXXY13ZnDKB2xw7T0Df9JEag4pkJfHHTZ
43bIWHvaMG/+GXmpuXeDfF2SGQqDpjpVMs5RTt+N+PJPo913kqIxPmx49HzXgbt/wRNnHvZxqT2o
kiHxlduBErTFMfcKrRiZIVmNQS5PcmLh/I8GbTYSszjqjQH0TErx46ybmmrlA9pRj6jxLzFdztfK
uqnFAS7GLkFH5WEHZAopjqsTTTygo87ZJsjkxKO68DZqlCndQ/xCjnUyDuBdBdKxuTQ5Sd+s7fF2
LWRcvgyCGEODQgIuYemAVQP/689QB3XtiNNv6M924j2GOPN5DawvLTbcD4fJvM9NEHRfPbqT3uNG
gRkGYU7tVt/gF+KjwfWOg/yalpU4A4hvEYHMR0R+smBiN9a3G1YXC9nYEWiCDYU4QyeP+nbIWnoa
WqHWaMe7bKthvbgcIcV6BNba99ZUockdUlAYILQ5mWQqJKlvL0zGsDmHnSLKkwPbXCD6yfSo43U5
KNfRr7va63nMrVaDRG7EZV8hhhikf57qE6ZC/IuSOe6ONOsz5akBSBvyc9VK5VxN+vG8mP21DI2e
kuUGBTKoqZ580fL/JX5kPCWmjEUlBYuAyuvki1YC5clOFf5NsScva0IGUxpZilI80CqnGEVEIJpL
B8nAFlQRgbiae7Y2LV2Y04dIjvfD6RwG57X1EF1m0rjhCy6hcj+AyE4VH48uOFGBHqZg3Agu+7O5
CQCWsbMBV7Xv6LkpGqGJouq894ck6hg4xMkf7Vh5u94kiHY+ujkYHrjaMXt1RJRBcvapxplyMiim
xwzeYf/8sygawsCIOE95xhX7ZzuLpGWs2Vn/bMKct9wwocp4O50e6jySShQ08G/4uYHkrRbDn8ky
eVG/GXS0bCIZPiu8xyc2/Dh09xubq+SL97B9nXTG1fdYSXNpJHH12jUl6gz8XN8gp8rVxmMAiy3z
E5jtPHnhbFjX3YG/RrrZnSwrqvcNs4/G64f2tAiplDHv+wqtHcsoMAE41RWRKPF3UPdQRu/MBf40
3IGZw7g5HYQvsrVmMJrcjAWwjTbcO/w5dlZIOq2z5cEsPoRitLRCARd122zFcPqlBrRWyZnM6khT
ywbuzVl4xhJDtF6JbsZxCzGPpR6C17BHSe57voLPqXh7KZV4DuQIw0lMWWA0gE5wUThNmCh7ifc3
z4IlTP2guHLoCrlUwv5pHKRiPjwl4wmf3kBcNYOnbbu914Y+HtE4kGB0vnif1kFCetHSBBVNAhz6
RiPLhUxhW/mUsbgRGq8nSDv081n2OkoLgbR1snZq7Du8jWMZG777JNIKVS47zhKqMIKAYM2yiCoI
JClq7Pg3OWGhUzli1Qm43bVfRz7k65C7y5pIXR7mOm6ZdRs6vssW47xvN1XUBn/s3GNoDxH5VDnf
0vRm5f8riQ2Gz/mEfah5RYfJ/vmBM0fbTAzplViwyAWZ9aqjJ8ZvLffst17A53yK0maGU451pZhw
BKP10JAWAOvLUAP4HVGUImGGF2a6wPFj7OFRO9Tya9FK+bJWGBLOw/4EIqh7uT/FSFdpCVhCjvjo
IzqofDgx7HpTf6Wq4deBJtsZtLgm3RdhYZzIHgdr3w+DqYib0kBVWx4cHIhau1kQolHftOEt7ohR
H+tXhEhOZzew5rDEvaQy07hPoBgcCzXefBvNzFn4Dpb2vVuRg1VuPIPXiL+qjp9jHEgId0OixlUa
LjV/kh4mX9VLYR8hxglazHoWePIL4pQs6Grf6hq/StU8SQUz+xm8kcBu7IP6KRhSQKHCoZLMndUq
TqzKceODTOlbqNOSSuAc31ybakxAAL6JKkYUL09Jq7kJ2nLmbSCLib6oo4ku++Wg/t60/pcgpwaz
RhZyk5yTcqXEvi92+yWp/aSzD+3hyDc5GfCvSZdNjpD8Cqs2KGd29DFZKvM7hcCiyNHFtIqQqfhj
1fyB0ZLNrTUxoKT48a/y8iZgNmbn8xvOdptkN53i/WSkelM85FAi6J+OuHONzhMIXGRuRAEmFpJS
E+dNto7Aq3WceY2S5MX4mKlMq4E09Brc8rfSyaJCt8xekOkzq1vtP5Nj3fFdALhxkGfYFhzQWsla
uwyfGs8ioVp887zHJ54h2yfdzzCG3RLKumZ4F2wsa3Y9ic5U0Z9IjH415jUAE5809+fnWfJaLzSX
V7jALVsiITpOpli0ZoKh9V/eH8pCM67QS0WWLri1RuHS/ojMx/LXLH7yo0h2WT4yX7C7YZCJd3zy
Oge3u5/KLK1yGbcuNpUaX1qU4T5RSeGJF8nO+nVb5tb8qb5si1OuRT+vJjeUzhiokiPs2oHtN4pR
kdtD0JVP9rAF5EAsxqqd6+VQhZeWynfA9M65jkOCRj/ey+fbyMPUIur20Guo0mxUsz9RJfE2oaap
17XoPd8db5FyNqmx/yuzVmX5rDFJEDhhLBuYpwLlOjklbjQWYjzTzyzECvwy+IO1j/mKm7EpfV1F
iMvj6tx9O4LEvx7AWrTrL/UsMRpzKRkoKdq22Icr6VbOUVJNKx3BueV46hevBaNuHF+41TZwPKbK
TQknWbrq3ICfArk7C32ccUncTrNTVQqSAtg8z91qBdBh0iU/lQ1utTOvbN9iF5XocqxoeYjUaoRj
M1PZRTxnc0o1IK5byEo9GSubt1grTOW9PrdIUvUu2qfC8ofJ4TKgRVGP9ZjAYrc8HjRxZgOvZ8rC
g6dJNAsd2MACBy/k5hTTYJdpdLayp/R/kXxZ5P7SsRqLEvpdyEjEhZBWRmPKNfrWsd8ALOaDXKBt
pJiDSWXrwJUgz0wmxRGP5wGdTf+ogMY4wbB1dKBNAlOu37I+phUdePG7RWV5fVZ7jC32/Zi3E0dX
0Az/3guKkXc3wxz/w422mnJgIeETMIb1LoCUzpyejw0lgUSerbNAIL8zfer/q6q+lTKINSimNr7Q
1ngO0OGRdMgnFnkopg46KQAJMTNgqJ17Bm4JnCzDOlyfdot0Cr7vPkdrRRmG/DtSaXpmm70DDdAN
FlKiGVm4lHJxcT1zSy8kiOEnPoqhoVCPC7Y1utcGmEEJgwXY7109DAfPBRVmhRbtXRV+CYUONOVV
nSVp0PuB1mplil3Wou01tGkCGCCQWgNHrPCkmDDMOXR4VxXzT+R5ntZxvqTVpAPtqdkUdKyzAejf
kYI9QNyRn0soGrABHSBp7dUwmdlk0fjKv68KrmPOsLffAjx2MzqhRXzPCFYRSU8yOqX8NtoV9GWQ
W+XbAZmMrT/8jA6lFb7Ow5vwEijpZ7i/JjTDGsq0rDrlpoR16lbtasRoRcdOn55uPMsDpf0vjegv
vWSXlZStK/gc8PsImJzSx83/ZtVajvtTGhYN6kodPpt0hOvD1nUqEYyyljjEnCpQ4xpM1Do3+kcc
63uSY20dYcYFtqgRcnPbJMSWOUvE7Hwf+x3UCWvNuoX1K1rYHOalsqCq3UVOBurteTHBgv5ZHb1g
XQ3RCyjlSqPlN0aKVCMHCq6sN7oT/qfFq/Bm7G8KLnVTKYyKr57wQsaxfE+K6D+x4Y/OTlnnAtzJ
TJ/pHWvbOGh/j53bn883No0VwA98DGXqiSNdRJinNF4IwI/ORqx3WW5IS5K3BLTt1asTXavMyCQc
jqTWcgLgFrvWOncnms6d84Aa4vvPHHhBeHUZfgHKfK+erklnhIHe/ClYJF6z4/HvTMTBK8ygbX2j
Bv5K4zShAq0+DkkaB2OHmLChmv1e9U/3+g5XJ/0UptcW2xdCQbNPyn2TjPKZ84Qad+58Bjyvx80F
bi15uBGJOqusRZrN2kPUKV6GOctcESTAZJPY+E9bQ35MsWAmu/n0pavQHHMYoZ5x6pJGZ396lZOR
a2wZwq9xUWeeGEDAP6yKXPTPgehfg0ZnA7243r8FPm8k2qUm0HQ2BRapBPEN5iTfoeD0D4IUS5WH
2sCdSSPdlGqauNcLqve3CBOMIcJgixp6Ngm+cFeTwmV7WoMdoEsCTvV84Rd6cGbpDqB5wtcjdq7l
QCRdorfXoUFhE8iV09pNojwk6tKW0T2pXuJ/kclDS1M9+lrm+tTnARzTFH05txJvAKjhZjMJ5Yyv
IxQloIKxxkSJYapCutjC0mEy3lPMnkEqG5yzkzIHii++uKU1V1P3MQb7mMlcF2Z5LqzC2uQnYwuh
mdxUqVaFe7PV8OwTh9WvpXMHTVQzbFVpsQjAwrDz8XSD8jvK6V5SSByrYIW+HVhfuTMPt5NKR4xY
RrlLhZRb9V3OY4jqmwfcm4+xPc5lEmnjlJxS8z+wI6tpq/JWlDFR/nOvHlWBqA4BZuRARL/P1ct0
Itfr6BtSjLtoLw0Agim14FcCylvs3AVKf/kIpeXt9fkYYfFmJ2dHlQ+tsdKcBy/5RU7LhHFNmbsC
mTmVNFLNj0jMTE8BI7a+BNrtzYSgpJ1uPEJZmglaXFb9z/Rm7KkV3hHM8x4Ew246yGuqfmAwlmaH
dSOPuGp5Tgx0cyTCXAEGv3HvKxayOFfvrc+MHN4gnrUnWo+WuhU0cirr/dEOBc+3p/w3XBzv1MOM
XR0cBM4U/9GhJepETG9OmIi5lpVZbc1U/MTxvnjC5v0XGhM/QpyAlQJXhJ76Zsllr4WJhgH0eJel
E3YYrpBs4DL6XZlymctEqCGsx8tORtJhSeFPFAQWDYDQ9/HlUI9kMXbfZVUTzPli6sbIrhRxYGLP
L3ufluGHFT09Vl+1RJv62tklp9foimlDtrX5orT5xarpNWJU70K5SBxmucIhkvKSxk7LS1El88MA
Gx4eV4QglNAI/0JkIrG1uhJDs4JBu44mBvIr5cT+twcAALPLkKGr9CL2GWa9UdPAtmhfzUMKvW/A
UBu0NSdtrV4l70DIok40Zyhpnzf6zKlM0eqRFGwXL+qkS8BRz1haCZWNZfpJ7BqUXd88mRhm4kTi
0bQ9PEAvTuvisC/59efuZEQ0/B9pcqwu+Kv+hStH5+8C7bo1OUsqYSFPvsoTUH1c7hUH+Ulx0g9S
Eu8svWDlwRbvAtLoRs/mNOWmUvjZnXpHf/dAnCvQPN+1+0aQiaTItUc4gFAANOrK0zG6qK0+RcYa
cH5aDyUJMiC4AcfuN2YVQfwn1yo7IjLyvvIygCqUtzQG9uJi9hFskmiAxyOieZAWpUK4H3/1GR/l
eJMZtSMe65NYSABh8cSE8Gu83fFGiqaxTD4f7fWGa0oGTw7TaOqQn9bjIOTicg0UI5hauHG2m0WL
CMTPVbXaDXe2O2Up2cyJeKGjSCfrvM56hP2E1j9/qR4WoHhglqSrSYQr7E6Jz/VJQtk+05dJgqxk
9qwnU078PUxiPLFctVh5tHh9mIW/4Qq6r2egiwTS9uTZ7AX6a5UQuGPaKFLD11p6k8z/zmh6rt+C
ZWLB4SoV+7YOfEc2uzRUMl7616AQNNVR10ieBiJsm0gQxJQJ/s0VlYkkew9RNHpPWEh66jbsz4ny
glvIM2kZo7s4/MbYcXQaDv0N8P3Ey0/QZeFFn4XUae3GfhDkHvpRZMjgzbu9sCL580plMUxNZKFK
fm0UGs25H6BBk2g1iGEIzed9sumpCJ+++NbU0RpvetAb8CoiPtzQeVdhHv9ZHVx71wLaIghTZBPE
+o2OfLy1uLs/CRoHuZPMRYMSg0jqzUyit643ChJNraWhmY4wfVCZp35CPZh/3svsZgukMinxEu1R
08DwIsNdQBHuPNJP1z9I63iYPOwhi8CFtH8t/JuNUAihEd86jG7y3msVDJ0UBE/umVk8aFCMMlGS
9kSktzyeo+c0pwrnRl8X8b/SggQZecwy4FqKZkcTqSebIOm6Y67jOycDAmeymFdCwxkpNHwTBCvt
WMXbw5XIkPmZhBCtyOlfQ6bczQVAd0l25ELAeOZZ3KS1RXyfu4FxdB4NIB+ZnAGAKLjNfMLZDmpV
v5/5Mt+ZXwrYE6N4/q5qf7hy54FM6HNI9/sPI0IRSScHre9n8hVJ4Cmj+WLALcwDuHRnbQwwyhot
bXrHfVH1PZKRgdfgaedudiMvISplgU5eAiltOcDSyZBQ0UvWwz41KiGDZ+o7c/+8T6jhZycqiPwG
um0eDF1KMRv62s7OX3RTYTKGkwE7MqKSJN6krq1A/TeGs4orrNCqVS2mxscXYZghMc4IgUrKoYR1
FJfPj1klRlo7iglyvlab3nxS9BTv0pJGvH/RAtPAJv2ZiU632KE6PoW4XWdPDbAGh65RmeZIGDV6
L0BvrKLhyYWqW93oYe6ari2XcH+bQkiyB3R7gzLcrVAd6YY0iPi9HTj51Na40JrcI84Bwf4yDDS+
PZ7v4K03NvOl70nJjtSrIumVgBgqYwisRB23drdmrTdlQEifUE0CKviPzIT1BKhyNiKXm3OM68+B
YV0X1S1QEG5sWbmbpMBfiPtfHrltnQLK964lZeaqdYfVdSaQrPusBjv8dQqtrar9wobSDK5VqUGV
oC06wJcXXgg9Zv2oeeHwrmWyaKCb7agM3ioviXFi2yiftMAbE5ZvUMiaEn7i2Z01o6kR53CY4X9W
5/hXCHgtYQFih3bHfomDZeU8HCvCLOi3+0R2dK7gFfA29FZMPtGXmGmRXXTgJ4JB/OvEY2V9Ykdw
5EUMSCP0y92A8qpdClKHNcpgL1DUh7okISMYrpTjYvRBzQU2GPjX2S1dsPCRfr6mlG8+dGbkbnrP
I66RnRT1tLPISiQcWumlA14ALmaK/XEnZHU7E/WaXsyX/R3i7l27UtM12gnnZ42oyy2vwK6JIEdr
eTski8yKhvzSnWERVqY8oAC8N4ac4LIpn/T14Es+PlRdnEEU5BOc6u66uDGfSRvO59fTGVco5Waq
UcGA28xP4/dp0sJj9ef30dUVarJwlGV6r6aQ/lz/5d7ptYs0e8emCTUUhyMofX9oLwzYkBmNcfvV
4aSoX2prOfMlC3MsH77aMX3fXGVsZaSTvMErKOvG/muEa0YgK6BBzaTGUBN66zsML4dbEe+zoNp8
w2eIwA6FZ/JOJSGHa1iStg2x+nDbfWcHiWiT8NEVBWtDX8nd4SDN+06IxYsAxNiiSFYLlbhOAxo6
I3v2LU6U9B6Vj0JTWLU8vSoVDK1Rxwt9MEeD8+6VBvC4g92P5lTb9mmQTxEqyxFVv5F2KOor8OpO
XCeeGfggzN7CgIXQgElKQNYgkSjPCAoLHU+6rq52XGnjBn8adOdmek16Ex/JbJ1RwR+97suYpP0e
CBfN6OJirjujHSvTraqRedb5BG+Wwn1YmLNhmbBbF+ZEzK5VYQbr78WWwnRQFTGuzJh5qbTISZRu
RQtpC/O0C8lTyXy9PvamnFX1EAH/CgSAT/aO16WEcPkrPS0npfmKXEoQ7GTDZdpxcgeATy5U8E4P
zh8IHaFo2hpKe+hytWCiKiSfZ9dNzpngaMWc/NEV3z/2TnvALtVGjQwKH+gQHwMKmJhCdUO6Dhzx
vBF68oRytZysloOvSXtn0L9fEV67ozNTj41Dvg2C373j+7lz6cpYWAV7wQRx8Sv8xXdQSDq8yLve
rVnoctTDTey/WhErJbq0cbd7I6itPgqfV8R4Hz6Cm7QPnB1qzUKmt+SZYME6hXMu0ABj8vwGzv92
3ylrhD63x2smIo+jyO8039iMionqhx/4HQvQ7071WnuEDtsmWR1dQJEcg0GpHLrRXEbFhtXdYlyP
okFeOsbCHcgDy8JYdGC3jYwmvwLM0G6YZGPltMrr/ZjHCrLRVVOKAk6uIEz6vQPUw4h0FIj8p0nC
teLCJA79pNtWCsnGhXlTLiH577IzoCSjtKPBee1YCqhVbXAGb+l5SH46SpqwLUE9l+xyxUXS8Mp3
UPPdh4gZ5OqTXxmINbdsyTO4ZVDKK7YWNkanl25qmgpQhrHbWXRnHZcApSbobPd0deQL2FQkHRiB
r8fzwlzLxtyGVaHkAQrOslat1DXFl1lybYALW9Uyag60dNYk/p7yKgWxOH1IhXHsEuCg0u3tcLKV
6ySGiqFheo1QLIDAsgiqc39VfJeRJKRF1GyTM4AeboP0tsrhs6l8mDlo7gpqcrgKGlVMyrfSx8Qb
OnJSemoZtNgAHGfHnzsYoZ53HclqN0pqlhdkh8XcaEvTUz7X742TOaEclgfGQbydoXZhdLiJU0HS
l4McbaCVtpH2KPUsiBns1+rZSAcwVWvA56IBNPojeZTFFdmjxnexGm60macU1b3DDMwdhoz6EEnz
4aI4eoNtfE06qqacznjDNx/g4rY7eStrfDPtvb0qLROfJeezOgyN5SiHHFIDsyewjDdVppqe0+4l
Q7+OYVJOc2pzIiLmZmHzwN3gEiWUFENUGVRhQNnovKn28cDgY04koqAsRpXZRwvnYg0kVOjYYuP6
H+c0S2eQehpcZeQr8stK4aVsVVGuc4peu3UhtC79WSj3t3IZPEY6v2TyBYUPVQuOFN6JJwhtGseJ
Xritqdoux4KwKywkjanTQCw1oRgcJsIxF0SUDggJeMjunBKczPN4+M5bV2uHsX2J5k+zeQWY72U5
ESoPSAzYeYzmgGckklF5duTdM2sZgZHST3rBs10mLbx0lZdBg+Mb+IiwzYRcxbEbcJ/kdXlzPCwh
XFzFuyZqILSaWy8VD9v+hR4byTxYm+nMol6v0MLa5vT8rfH61HmHMrqqZyhSEMUdbx8R0ylPsaQM
B9MiqyHu2mDMf9ZeY8knao5hX3i/VvXHW2H6fJl6YHYVmQ/N8j9wXN36NmXkwwXlMbwW+KPOwr2k
bBN+KZm0cbpYd0MT4aTDJ1HLbYOFgJ586BzGCfkRllTQe7dOcLEruIlhk5Z9mN2dx4+GjZcWIDJG
REgNg87KKZptDttaNwq/GdmfQcRauJ45JIfdKO8fBfh7R3nYqmzPNbDcGzlcBzjOejNSTbglLgkx
5TiX/yF9M3k9Bjh4LE62oVnaon1wEFIhO3KxTp8blpsIZox3v+170wkUsUSnjYRG94UBTwftaC1/
J4baYdKwdp0uGBFarx4M+0twva+wOeAVWVvqROmdwM2YTQ2uwgq1EoyEY8ZjLRhliXaZoCZxMutc
MesnJY/IWqHXfApDhMuUauZ3+bpW5w07kac9jlOreqMrYbbZkUijtrqAKaP6L7UN3kjPJ8HmGTno
uN1bteQ+VrUmIarZbhdIHVhvErjehgcEpDRx7SR1p7dFL9sqOsSpf8cB0AzoFrVPZp+qMPQHMw+4
V3k1xWDBUmsN7wPkNCMNe/XRKAEAlNJoBlDu42n4u1XTaP5OWzkxuZFhF3WwQBfobVc4rUOXmcbY
qM9RMOw7YF7IILsM9ntkZ6ZEgUvxfOD/dr5UNXrWYqCR8qL8x7r73XtTxljD75R4l8ECLkygVJmM
6BFcsqrKw+ZEGZ2gTKOZUJGEr4JGI1no4r5+7/HiwyitEG9sPoON0KxZMmFEP4a1iTM0IEmwhqnq
rWRREmE3gqWYXO1s5hWAvqUBl4CKyBbjPz3NLoqvp22v66DK39V2GD86cZ+HrkT5ZBYZHc4oPBmI
3jWibWp9Lt/s7hgD4fI1KsNa2+nZF1kqM5vdvExSS656Xvfr2AsOglqf2bxKlcl32yogMEK6GXau
XasK21zY4X10oPhZE4NuwUrEEh4z+f/T8cdWRrMhQ7KedF6UP7TYi6RK0kXEvEJLQNpHmqeXLu74
SspRjP7Q4MfTeCW9VpuKbboGT8l+06mv3AI8hVkArc4UcPK7qwUvfDshmHEE9BCwitIm0+EOYg9U
RE0sNmbF+rlSWTaz26z1x2GGuUpfj/9PRkx3vCzkoymskCIEK3jSYKUC7RptlE17MQf0KsWIedr2
HdDhlFSWd/G8KjglDBmctOgNDN4tcw6/M4y1aWmVxw06m60Y311+I0RzcEaGwJ91LlYlYHJgJOKm
d07TmH4JwVaWeoEuykJIhryWcTgc75bEznqUfD1wyf0oRRNJ2qaeMgH2fHq2lK7lnY8mnCatHDjn
kBIPbzRVWb06UJKLZc2yLdrP4dGoCjOjHJuCs26zzMOYJ4DR5zDJeArdV2tLA3C81AFogWm+qQbk
OEU7i0ISH9JlEG6OuYxnxicO6nKhjcJ2HgeIbFoTUwsWvP6rEJ6pCvnmeNdBOnbDF/sOgWSEwX9+
F1X0M7HK9LAJeQwX2l8p65r8esc7iNYlHn0J7scwPrFKVuZu/rg51WheuU4yixCmEC65rUSsAPUu
On84MRdRpvf9S5w0+L/4ZTXvZa6WYEHHV4ZpfMubKpGlMrm4uYSM9Ajd5ULPHlEL8UVIIpZCP9uk
NG8fNEi9naNiT9olo/f0Ki3JR4IqjRQWQV7CfJ8E1foKG47a4KaBCDjzk2oZy4h6ae04nH3EeN6D
Lv1wEln6XgT93T8G+eEMen+gBSK5h8S8d/sWQRChWsF0fbsG1gZ4bVF4jcsv37LaAO+Bdr+FPIVz
VveIq9fewY6+SzUSktlkNsBKSiwVMyxbXo7devUM5hB93P/F/7UaA+QIsvzLAvBaTR/8xuIbk/xv
+Yw1FSQ6JjS1YkINNl8Auhqo2+RMXQapo/WB/SkZbG0V8QaQMBDx/t+0Ss863ShKNFZHIAg2B3Y9
KV8l9DINypXeUrW/pvS9wlSJLSHQUW3VmN6xWta9mWyueTSl9RaqW4utvNHnyVKnq4SrQ4dXQhDh
SpGZCa66kDGlw9gjMPzuCaqxGckhZxcR2KWernAA0Q2AERQdZh+tLfdwfaFiwSJ8tl486hHxZAcW
IZNM3QygMalEkEfDjw6kK3rZXSdiIgaIlJRuFlqtDeL+rceJMbAfjzfhRa8BknDBf9QwVGmD4Egm
f8dsZdmJ7aBmcFqyuR8UiahuMY4EpRbsoSDEdu0pdPhynDf8VZrXRJ1uFL+e+bNi0IcnwH4xzODM
EkQ1TmCWqT0AAYDD0VesQ6KWe+T6tTFRu/jA7uHxk5SdJvC52GUT5g0Iynk3ivWbkQNj/edSpjZl
ycdV908t57tiHrW/NwTQoVG6KY6eL1ysQ6haxVUJu47a3oMYRpx7Y0ZO5Ck752urHkvkjEJ7aW52
whT+WutXxacDFdiu0hZBg+3qlitVv5HurlmyFME3Md7KdD4qIUwNgXxZVVfo9mC60TgkfF+Eda82
dcRSFk3/Bpnec47H03XSPNOClILs38rnAuAf66be9eOMUj8JBs/POpyZwOshFWtEE1BZ/of+gozR
met6G/hOFa5YnvMJdvLzPkrSG+KVWbYpvxnjp/jsJho5QIA8cQtB2S84gWc+OLMnGQIz3yztji41
da+Z5Vyjo72sh3/kEfdaRSTX15e8Vt7P0mAmMiEbZN1kxXCcCJ/t/0dzeyCViMX+gu90S+5TkDJo
tjNav+gavUI//wXUVzUk0vdzBZdPrfk9TLeDoY7mZHljtQvqCpi1rD6bpiAGh8p21qI31bJhIeXM
7FPtwYIXsiPnTM9VmT34JRYPH3LseAgCpuhn5aqCpBmUN6tEKx+R6jYLR9xlNEBnPr/ZSfLgBZdR
zyY+UCbvgYznYL3x5pCzrtklo36ixjyMsULJeMi1LJiRsnfFd1bA6YNQ7hTV5L+dFgMxLBkXzp68
UgkwC7+HbNRzD3DysTFatgvnk3fQOY0QvGw0qXdMRMBPlI9rrOKHeceCdhfFoXQ/7Vt0Ocll1778
BkLdab0qsw7ZDSlzuSjFEtF5l05U+Rg1stY4Wa8DRiSfSozaqCLzLPgb2O6LpT6nFBZbjhFSjnfn
fp60zdHNOt3t+L4bHrKXHbE0p+JBL1aX284ewSTBAUveTdhkejzYCrrDjyq8JGXhE9Qfp4sRIu4E
QssDqER93IyUlMD+MtETQYXXanYDXv/veJyAEXBOftPSSFBnD0+FH3Fidja8srtrHalHsCtPxiW/
DgK+nmwKEITr6j4ZgaIWeDl6QMQxnG0IEm3YrircOhi0s8KZYXenLS+fBRGrSKn6eg16QHJsq1yi
usB0QQJg4XB4eKDueht0CHGtnLBYjeeBC3xA4zK+0QgsEZIlgMoBsIV9SCX6aEoKFm6oa/7wz4Tr
V+n4j5KeLDE/Fq5dz3fsp1D6uKELZxZbVqQiYzukEj5dpnPnLiCjnG3dvKSpjhvNBgaRyI/Q7zSX
chA+wxLtRFmmsC4AsY8cbTpVIGMhBoaysTdZegNj8zJv7JXif8EhEihdLOJySEvehrMjE+/SE4Qm
6jvSZIGARSGu0esz+eUOIOEct7p4tIWbsme+zo/XIDK9OkkrAV7gNWg0/Gpdc5Dnr4jewpM9JRfr
ro3ESGYcSnaMG0I0Hco9SKKpUp7BXXkmG+HQ2k/OESxMfxw/EE15q6V15UxqI2zByEKQvSyRwm1N
9LvkUeshInMS+P4RB6qytUAg8sZozioXmQz/oCeh4Wf0s/b1NfDGSTK6Enxoi+NPUw1pPt5fbknI
+1FraBpBwUPsvr5GGPtO6dKqzbeWbX6Up6vHPw1VlrYVUevtLtMnCyeYFprIEQmt8xeZqMSjhxQb
Kodd/sDOka88iLs9loN/T7eUEvNJqDIG8bMIZDM49cGvcsDHWv+tOLQpEVzdzDYcsA4S8GLJa7oj
+a+QVaxrZrAHEZgJlwc+bJSQrPp3a1qFMFyr23QdTX2NxgMoocml0+eDjL4ZrwHdjLKYT1Ad/SLL
+xViUACzke3V6nqMfM4AnhIhuDupZFEn3JLamZ0MnoVp026YXCRelhaFANdajpWdBBjrE0E21Ff2
gtpt6wQMZ7I2FJu5RLxDfCBbpHnwl3wN9eZgswBqRbBgRpiZvKGMwDNGneRBPWhjX98d63C5v8Q7
D0DT7x2MbF0bXW8WFV+k0adJCeyowDAyu5Rocvo97dIprhm+4CxhtZ8nqPPsYPduANTvSmCne5hz
/nA3R5iv5YqH3oanM9QqKQCRJQcqDOAFfY3hP/LP8KgMk2oNxiN8x3NxxIsfM3ulQj0x1uXVcBeF
mPrOL3HZ7pHQuIzOw3JSafmCe7MMdZYBCm4HAXNz5npyM0FbYqeKbVWCKYXzD1LP7SaM1lnQsV3l
rtdEAwwrmFFNA3V77fYkccpyq5Q4oMQsDg5QJrvukOpVCRW3gN/8wdYzyAdmQb82JJwNC49W+FKX
FAObDIpVZ2fq13FEU6aYapWv2R80XL5igLdA9AIkfIfQTX+hTh5aXhg6YT0mfN+aNPVuRj0Y1iRV
iTC8MmHFd5wRysT/eWlLKnPODlAQqCeh84DM/ITMgxTl3L8p1TFOPyoKed1WjW01SOTU7k0Uw3Ah
ALOoUXe4/Jhu3i7jqu7O9K08zTNfUbavIzDOSnVUPSg5A4wauDBuho2C2DFvKehrxFM7ehNEr8Cv
/Rfhy1RXpzfy1Q0geylwpALE5aQNAWxyjE7H3oAiJVaX+BVVHSK1QFK0zfznD7KjDhl0RJvVwQB3
T0+1qsBe3I/CSXITSzTfV8fnzhcHny2hGQZn6E10MlGpyAEPHrzCrPp4zzSkvtQj39RcnMOGI9Dw
FmK9dn+wSFM/3WdXt+6zsgjCi7IrC8pOXhGSLvxchl27ivXzpzDPdSju7NdW3c6KZOwc9oIgPTQ0
j8L3D6aCDaekdRwUYx1Tizsuuz71b+l7uk/ESuACxnsNfHVstZA2ADpBnEzKy+2QqU5UbmAGWKrg
bwNopDJ4weC08zJNd9VXz2M9D+UGAE4sF1GvZj1L8ccauNWF8WPTcAix01YiHHRnCQrz5G3Y0B87
AYlt0TDilTPjr/3Eu4CIohO1U0yAz4C24pzbxHZsKDNHNtW77QWHldqS5wZemd74kBBusEAbpd88
U0Nftg0lN+GvR6Ol19weJPKlrghNuHTjY3F25uqNWYGltKtRyacXndPLbz5eDbnlZIjCXMnmuN89
sHhtWZjMy4M0cO9B4az3lJWs5lxbe3MDH30N304kWvhFIAH+8MdNRBHODRh2HtHStgFd+NjK6tMt
wRqvHCJ3kt7WehVGn9enJv1IpJAQ+HtRsGsSXQ0BDGP65xsVwy8j385VBAn6/IoyiHRxVFqlD0O2
BhJ/9N7GBhebevnDGtf9XBXmNoerin+uohS8KU1WuMEZaD/bfZM6jHnnumsGBeInYOeGS43e3rwh
5goBhUUVoVWDNcDUfFRyYelCWUtO9GrRf8l0Y/LtwMuV2FX1pOwB6aMIF83HhGPwZQbMWtGZnq/z
oE6vRWY2bfeJGlqvp13i9SQ1v5OcLqtwtyMCxqFL6H77AEOen/4gbMt3yAnmPnL7xBTY2m/CPD9/
qrrlr4jdFBm1XAr6vaXzYBzEaQdNhT7YfSuoQrqpZsQlvk99bu63p/ubIKqXOid3Nk5j0oCMxT0y
E/H3waDRudcpkOqTzUrtERqvfaX8iLfkLgI8MoeaNErAxa/hXnW2NVqCxHazN8YixZfw6iZCPR90
Micu5jHa0JiXzjRz/TnEmT0qKGuFHOqAS+hqAEU9kGLW/zgK0q1NhmKQCG2cuYS2+mgv7JLFNfOD
lEe78nizD1GVJCO3SvyLEc8hBuICp+RFgqKmDWrd2KE+8tQAc3vGMtPQMtjKL9UlkIepVe7c7jIQ
tTQjIUEN3pK3XiOIXuBhxdmZK1+paycZhq3zM5I0l1wiEiA2n9TAKESleGDmUNuw6zaz4ymmhO5S
66Sqx1f1NcS37mTqCV9MraXAPI4GQlZ51sdnkJ3h3B8cFQjiLLH+pM6zUZHefGtbfsnJHTrX+851
wMsWpKsHKbSwi9OMvqEQA2Ar2Gt6/2z4KT6Vx7IiLPpelVt/IdhHDAWe0bXIipTIUBJcE7CDcZ8N
VEdoAqQaMFhLfwmrYIGsfGWiFEbKjts1MnRCT3nMT1yUpJCKknW8fV7EAXySA4wS0SDjg14nWsEQ
ig9OdzKciRQBsuN9fVq9W2axGd2Y2+0CW/8KYpbSg7TwMMz0WLODfsTUouQUIciiUpBQU92G7sgL
K5M10S31lJRqWtEJGKkD4BpcVzDSl9kwCC8O8IObIVzAcRSXcKv7LBGZpBR8JBUd7S4mViNQM3TN
2FnnqmsXr8UqPf7RTa/Offv/mfaXZbmzMj+4RnTwPAv34Uz92Wb4w+mwqCx7z9oh431lyPTZQKDK
mCEEnWz3BA0XFhF0fybTY5aHgIPCc6P6NjBs7XmMGJJqtoLOMdjlk8jjdSd1Zz4QZR7u5HlViEvs
Ou7oLmKV5KDqMWuUyJK8OY2VA/M6wGsm0ZHbj1YTinObusZAars9hkv72MpKFAWuGfAGO59VX1bJ
IjarJFI7YJ9i8lwzlifHH2hIAV73fZgzykAR+nyuXYEIJXJL+//aeRdaIFHWQaUOEkcECMB0uMhr
mgFzsAz176O/lcRT8U9IrXNp8UCMXkE+8NMkxjVxf3uGuPhQpmjnSi7RiyhTi733U/PjsKeqXTVi
28RtCz9ygWGzYw2hBBTuAgpp6HFQHKzB0S8aXydnpXxctFOJrAh68FUxN974OIPOlXXtKIWVc1Ue
RXPk0RTqk52fN4afU3OFLdmEeFC4iXCXwf7cDsJucSHUZeFb/LTtO9n6iVTATy3VJdhUEJ3aYJ6s
x76yLSjIt/X/e48hM9n4hIgup86oTgH3bzaN3yvK3hoSVK/7JP1Vr+8Ka8DrLor1TpGsujRSa41U
4jBr6hd5twWyty4xbDq+axqC9sVFSlilCZE6XgZRs1YWQ9CCBl6E0N+Ug9Kqn+RlzOe3oW8RCPHd
GCGxW07ptqdkY9SJUHeCSoW+ojJQu5+3OwGtSrU6UrFeGjzBwG+93gd3L46sk/MIOnKw/fz1Mmv/
QMtH6zYxbtv1ilZK7DFoHgpO3bmSHAOq8Kur5VD1DIWdMoQfXuJ1qWhxJqMR3xOc/IbfyGIGRa5y
OiaZsW6Ks2bsYdSnISrlg5Xb/Ek3TuwDM27t4wqeSAISpPahDwA+JPuuqpx3Fc8Cpih03s9h1/T5
H5wnjPoHHAwIhr13+l3sEQyu7YTWbM3fIQHmmfeJXW8Z06vQPn7kVLLWk+BxVH0q1RPOzA6FykfA
gqXzeeVxkZg8C11yRbUDydogrHnyHTB6vaFJB4Z+hdhkOwtukeODv8UrJwJrABt2+H9ZWCCR0BcK
gT1XjG4nPaABh0Ig3y/3py5E57va2g+hga6lv7WfcnQaZzakOEfa2thQyQGCtti9pxp8miaR7mUt
GjN8DWYnlrYHNT2mmCfa9ND5G24MACYpov2xe+uo9E0pMhcQmROVrC4IIdX3vHCQ7zzm4wjZt59a
en3eAJwAai5YIMDC1t4+19b4erG9bo5o1BTa2jbPyPbQ1chc0mjUqQykA92fJIlQmXWNyxAOJ5Vr
H2KWyqWva2gW3/R784yVnWO6h5wUM1u37ridtT2WL3W6g4hacHo4ybnh7fU+Wb3CYDNrVDSVtpo5
L57qsFeqzznzXUo3eRlN0gyPd8srUl8lj/bYt/RWeJLEJth5FFJwPL9hYqCOnqA/JzLjGcCuA2RL
bOgP3K8+ERQAczvXM6XJDw0pUyX58m8/26rdk3LDKAAmW+iLyfU/rNjN6Pp51tAdIhbZOPMSbWF/
7FX1IkXuoTR8hV1rtCTmXGpQpbDo9+nDm44/+7xpZF27wp6FeHI2iF+4+efRmd9nHmolZ/OuqjPn
WBnFFLBty8nUATlOaU+t33edsUfmNcggXYl0r1vwkFsClt6doUAlhet9yEFArLr5qZ69KnMDrU2Z
V/UXmwE5uug+etp2i0yS+FSULEngOrccQtDEbMJnLYSkbNg/szdeFR0YZ4k47iXcxsZpdyxWIAfX
nqWacqq86ZKlX5CihGf/SWdvTGc7LI96qS3bwBbp5RW3ezev0luqJln4DJL55R5YnepgX9rU8DJd
P663uJQDjRGHzNxdfipq6Dm9NzRA6oBhKkBM2SWfHgNnf+eHJAXPjeFoYLd3kgdO2HLkxRF9xgF8
/WNdBhiPWd7jy0isA7sWNxZpWvfxmxLTd0Qfb0oFQSq/3BRv3/Ll48r7vu1US6upAxQ/TrczoFyV
zDKRd4QUVzvXfR6RMAMGW86nCALQEGZVDvT9nB/YRyDdvCNAehvVq0vffTjaMoFZ6569WX7cswpW
bval/GFe7ra0SzLsKs9OAj7ewX2EZkTzx4FPoS8q0YQjLJTMsyQn2fxtkYXwt5CqG5RQur+shxOB
D1/cfaiEwGLnVDbLBchjiSOltUrulGYawKGeDiWQweipVm3E1UiLYEzbXU9sOlFimFjDEFuKbzSj
yPGMuoY0lQsbMduO9/JQZVxsQLCaHOy8PkKB1YVqjPnpzaQ+vjwmmAK0hJYsEaiRScQogXtGbhqR
ZpHLufoZE8If3qUC+e/Jkg9F2km2tLqKTSSyE6rWtPrjKRJCV4VMITJk+Uc1AYyquL6riRyq5Es1
x8ssdhJfRH0Y/lkGhJWPiigWjqEOJ9TZIBaBahQYsATdcgAC1meiINATZzLYc19ATTxIo7MTlwdD
6cJkM0o3vE/6muUIlPtXJhlHkrHHIVbkLJe+vUDUBqZS9+2hEksoh8+/fE2w8MbUhAE11ieJCOLL
UebUNtFtBu1w0usnUHLZ3D7lVL5KyjOM0lrHZrL/STLipBNnJdpqIg1xPaWtaxKxRTK7VCOnTl3Y
+/04pZWOeuEUO346trqbo/nOfrnctXfAuWz+fBPDN/3lYb0NodxGpmFBAUP+WK4QGfScvXzAhLln
0iHsMfl0SiA50pSQsklqoqFAAiF11G/o98PBoL4lX5MkyApPSJkRrQ5a9BY8a5VIAM/zBh+Z50/8
1/Z9MF5W7kFk4ENJWvQKBlttZ2QEJQMfAibzjJZHdnwkORBvC0l4r0s4Um1vcHUs7BAqPk+AHMgR
kkfmDjLy63ZArGnK15kq4puk1+TAJT/QRnFNoNyJPAFS8t/e1CUH4ECE2heF8xk2xfd6mB3+R0aN
vU8Zzgw9ty5DU56KynyHdJI8C5K9LuJVD+N7jkBbwyLkplyB8oi9/wUyd27qJzxdqHFaAIbP+UmU
dlarSVXJVFT7RXbtLYWk3qdvXvGe+aiYhhpPvN7zwWJWR3lMXL01s14+hUpc2H42E+DjK+QepNWT
4IaqCpSKIfgb67ns88KreoqwT+9KPlUmDCpSk18UTXGdFhPGWplWg5ABSSEXghA1Ld8y8jFMYke5
Egn4ZdDBetMJCQgYvNL17FaDgJ5frAUWZeIEKpcWWrjKR2R2Gxpd3F/+NH2BqbnvCwLmiA1Am5wy
ot+vTD9AAa1C7115s6Eai1osLOh4Q3MhxHyqElJubDhOEqY1XTN+rqSlNuCO4EAFHWe9tGHt12GC
QFCaYIrYm8hqRq9P/Gl4CImH0R1E17ojrczeTOSzNtkUdZwUGsJrnD4DkNZ9EbPIaD5hP5N4v7z/
jEsMEFOBdr4thYgROI0J8iRVdSVvi5W1/VUpVUj5z5tM3AXLZghoT1sXvexyzQbxdHqeHh4jvt+V
3zD13P7OBaxG1bZeR1lQwFQfuGz7W5lxBAH+iidwze2ewkTqfw+NJe9I9C4PcPFh96hrWeFulDM2
B0v9KGMwfOJ017Gmah8OorBXiUViu3HcXQ8YcVKtrt2oLXX/266P4prjZKceFH+GZIz++pRbqAD5
k3ChLniBwg4iWpDn3wH5jbg8i9Sgc8OGr5Q5CcfaQhSeOzvcC6+2QTGFYtZZalo6h+fXyZCrL/Aq
PwiGJmSdzz4X4h+DGOawRxveK1PvnnZg/LUUBhhW+g/9ORm74KG/I+g/YV4mwDOo7AUtl3HH+uaF
XOS2bYXLBnLnQ+6wwr24Xj+FXXWMxA9VjJLMU75tae1DgHIf2Q6wwgYt5BnELlcHieRMw7WbBkxd
VHxBOWj4qfCD0sVstaUDoKcKP8IrQ/GdXpAbHTwu6ziStgkHpyv6u5/tqqFGKoMpqwZnB9hvdzFq
0BEr0Eb30+hZWhiI5Zz9EDGVNLxATcqxAT7bNWmwTtAg9yo8Mj3MLcwBnUT0SCiKmDwyFehefCJo
FIiUGknpzoXhEhQtjLu5tkuAmlVR5VhAV5P3ozI+mA9YHYzB7NU58PXeUuXld0l8ZdH4cK+6RaUI
JhZQduXZQ0v88gfJuuJ/a/6wOHCUNAPc9C7y7MEOCwR4JN/UmbKg5UXmeHKAfN+FWRtNJVZlNYRt
82YEpred+46sYWyRJeR3+Ce6nGeMpITHNdv1Fn13hPmh5zvByQKy+HJAP5uFf0gq6fgBTLe7qVB7
E0DAPtRrRhmMq9NtZO7AeNdkIv5sFnQB8C+rV6IlfvP7c7GuTlnq6MFoDrK7UCCyNQ8qxD4Yiwau
c+FPKhnij5ID0Q+xLqeU6TNQcHxf0mLjgqzAVf6zWlaFGjmXBYaoCcIbxCkv0LNhzgjKXU8vlv4m
iBN7zOkHF8vOthxkugRwKC9M9O+fQDSkq7jW01rIgPebGs5eeLY5MlUaRG+4XS+7vV+4GBSJVVXJ
Lux0MUbIG14IxxT/BCL6J6RodxGIbLauydUkfx1Ulnpj2qmBwdX7/85Y3v2rOzhGwO+OYG0q0WiP
SBY/za2TwiSMv8bCe+zzyTXrsjtUF+JIDb27j0RVH7MrpdbfYEetpzpzAHVqfEL5zvNYEkW8TH5n
9J/K+8sHAhcAATLphOw9MsSJXWBwiDlDWFvdBSbEO7smuaOTY3BvRUmRmWGAQ7UKl3LoaAmqCNOw
mqiWHvK7WjfjVpaOMSMQ3xyrPNLxsRUNvmfZUrKcKNiOeXl5kC/B7V7feJu9pcGLs6eYaKIh18xQ
Zsh7sEa+TLx/NYcGibCZoUJt4ZfnMHc/gRqPAgLAnZqiB+DrDusuKsJ624n+d/XsAGnfiD+ym8pS
/QnPvsAp9U7LJMWwH8Z5RACo1PJXkGTtPbkVA9NummTj7tYNyblBInA/GzCXJeHrXNXt/oAuuUZj
8F7nJeXIScNp5aTXSZzetvID1U69Ync6DRgTMcx933HE75sEE6+e7iEGtEnpE8Mv4uKZ+JTi1xR+
keNz3IFpLiSTIATOkgtt532htLqz1SUsaXDfMsL25we5y9VHojpMnwhP2XcJgVOOMj+JeXpc3Kb8
e6M9T2i6pmER8LfqL9avF7dPaSGfmiFZmeV3N9yAhJ0rllYBNPG+dMwgtXAPeNRKXRFGryQC4vFO
SpKn0xAGDFkuciXH/ZOk2QKq/RH/I7TrPqJNsl+LR+T9+SfRDTHxmqhXWDN/znDK1zJwpFJvEej9
5YBuBlNfZp9vUTl2O5hLbuHAj5Q6IM/cvASmzBDUMB5FHbdD1wo7t1Bzca7snfuycktxnKbYf8kr
GGqFrk7xRIqgHekj04okuTqCGDoEd8Zif6EEuleH1DvroPfKM5fhwIBEhsvuHlyx+KPk6YHn3eLt
FTF6KfqBfjM+mFNNe6uFM2ecRs2vZDjlRLoKCENI5QV5L4t01A/U3eC7rcnJclLO4FT8WSRezyMX
67VftxBiSGnrM3O4TIxGSB7JM6uVgCukhIwjEYlW008p7/XaqiYSrLpConj9NdMGnWH3+Th8lRyg
/1fzIUpzcFZIfEYkfdZHKsfsFJslgGJEJU/F4wbAC1SmcDjzmWUBuTfXw7geVYfSksapuzCB2YtG
ajSsQa8/exbclp+r6XMo+rGn3X2JuQ5utCH1XsWSj2If8iiEevi/InzkOLg1PyCik1vnwvaA2o1c
8Xu+h/wNNgbX04bjndDnukCugMSYu5W5XIkjrHbH3bGFcKInvqyrdNtFHTOD2EM4OnX3ts3gHCqd
PBYZakAIAlYVAFtdlRNk/PvswyrA3bYu3vywPi4skfjnxfBFnco80RmERSoKb8miTPkH40zAX623
CsbypnXH9a+aY/nKFposs8joV83YfTGMyTPpBPnW0WNFg1mo+kt5hGs4ACyS4Oz9tp5xWlBV+gZr
9Ryq15oAsYZR2F66A/xYJIVs0KG3eqde4uXXy3GInnqH8kmkY6w/az4sLDy0FIx0SThAFb0RkaCe
imBPS7NdBiV7CmF4rCp5ohSG8hydU5lBy5VATtZRhh0TqeUe61y6wF8shVcxYDU5FaDnrlEYEhxi
iiJdENh+oD281LhlGqUPR1Y6wr/xf6Rv0AfLz5tbT3d5Ca3KftuRoj3pIIMfC7SW9rDhGjy0BOe8
y/WGhfUu/u9FDF+Ksn2pc/HeTMptmjSyRauunPxtb1dMs6/pcaGPj19Sd3v7nC74FPWGY7TMH9Qg
O3uM7k02jtDXbZEmT21vzCqdpfCm29mhzTANFiEAPtSeR60qmLmKDPLUc3O3t2Zyxbu0fiFC3xA4
i6pgA/xpe1EIjHLQek7hKrnSD08/fBivRanTtLvEUakrXaqe7iO0wYvlSS5wPkPpZ4w5iIKPLPV8
ulw+88XpKreBT/Cb/43hj63ARRnoOqUId2jZjZLA8mdzv60F8ZFKbKdAxxQqhwSSRXy4rGwBmcUr
lEpcwbvuq/QmzgV7u19Vtb+Y13Q8nhHqNnzNImO+CtWhgtZDI24rq92yvN/QR8Uq2neMEX0yqq8A
rDdy3Jq20qgTqx8QcFk717KTqKMJz7U6AAQGdXIm+ICJfvrKllouQGR5Vu5uv/72wV2xg4kR310C
R23ozkJoT1yy7FtpjrV9a6x/5a+8GbQ/MMWGtzXGkMdhh90vXH3w+5+9mrSoUFY1HG1Tri9ax+Fg
ecf5iJAWROLKuJfqGLo0T8rmWz4+F2eJ79FVcsiJkOwjOOp1zErC3d6Z69Edj1cBA2mLNBJKe0k/
DRlTfuhztB6OYYBRBWSJXFk458n/hiOb+zAOo7OwIPW5tq2AxXXK9qX/t6hvWjt/Y6LzRX+kGTet
BKJcyUXXwTz30ywpgt43yVMVJA6MxefdFpTRna0cH3VqmXeK6I2ml1iz3np+IxWVaM6uQaqgyyB5
K7sLVm8OsZo2l90BPm77uTdiXq6PhWISHX5u0l4E/rLgxU8g7aFHGiFOFikBjmyjlXyYjmgg/EY6
ts1OhaYQ62oHABUmjT+yO8jSjuQAMexV0TP79o/g4TYI+qoP+dhSSo+hizkfgugjYAB9jzp97w9I
EPwWlXXBpbVDzGSpTiB7PUBeHFdnntvfcUOcTzkRwVFEjXY9sYtpznJRwad0HKMYNKbqUyIqfvqF
vOEsB28czrHidJF9F5jomqyeL05gKOSSpiYIQ2e5psJFRgcNJxTxaSAWdej3hgG0a3QRuwXfpjef
SvkRyO7OMcdEVawHCidPWGYLElt8B/sQGdXWG9H/WLjSRZdWLc9aMCmHsSxAKWy3Ez00c8TiLWZY
T+yOLmcxJIL6vgcraPZ+ziy8jPvjO/ROctzU6fEkrcE0kcrwkc1XKn0Sz8s+gcvWm5xW2q9JRBu7
jF8ccjeOuaK9tug2YhrpfqdANcnyekVW3bgMKgtjKdkf/M5klKc0KVFOCovPbM9HddbRedTH2MG3
mdUYZKoRatxlNJMwOAMkj95VuH5EBHIgKynw4FeDLFPAQ8o1xAk5nzi9uOEc1+zGz5b0OmdOWjrL
J9VWbDKodKtUdzACkvVFjYfhttpZ9SRhwOMZYc9Tqatvw0d1zzbCnw+4kE7gDJqWjzcTtY217YIA
YqT0/IdBV6Z6LxfG0v6t7mflrPZqJMvx1ms0RQxgaekT7BzH2iawHdrS7cI7nT3aCKCRJF2wx7di
tiZyZ4fjc2IojF0nCfE3MAjNLEzRUaSWQLeZgXG9eDPGyCMaEOD1Wpi02Bc6qSKi2PY8rz9O9/uV
n/r5xzQ1rEyPV7eSGhGG4KHCnzCznhIh3mil8XqjSmqc8u92uBm/zHYvN4PfKqM0saw87yNbtyKS
hdq4YV/0/kUw4Xr+vPwlvq66lBxAKjzdLSdJZpnXkgDtpNghCGNCPNWjN5IGjRQo+1xEKoDu8CE8
NkOgy3IcCGZiNLmLkS1tEvTfWvh96ldjhKW19zVjhPsmrX/opVkbr+xMIewGgC5HN8etYdLNGwnt
ypF7TiksfDR/IOgSqEUkr36FAAyOhqXD/120jIms1jW61ykwjlRKtT+6L0E7kh2zdDaRMFfbOQ/E
Ld2u/1JWfiiwl7kTGWtwYxuNqgXAgAzposbfq0IWtUR+11RFQRiZLB2WuM+ir3WMl0YXHPxvDs9J
zeDQdRwt6oj5bXVH636j/v5Fpegcfckf+Uq6hpYNZxTKs3HRLLfW29rhppg/WEqA0Sq+DBCO+p+/
M7pFV2KDc29D/SBaPvjGiYb/b8ot5NycHkTUaPTZEgYTEL8gavU97jsjSCZLbAim+Y0eEvdGouQE
/9pp0lYsGTZ3YDS6e3oBcnmLexgIWmGMHNIK9waUl4YPH3+nBXN+FBmkUGtLpmlCxvM7OzJeDKYC
BT7EOE6/YzjoLnaZOQAtfQexnHnjX8WY+zt3+E/kBbOVI2Vpxe2kqNbnVtMIuMvUT6O87K6VmXn/
hjTHAo2f6LMqplUC4WrhJcobwfAd/acugcwNVQlwmwtKbCw4ioVsU4jYwdgkEeyM+fFhjT29oiyi
LM/Eb2n4N0msYvQAV+m0Y28Ilt70Q2r9yeMPcC/ynntQYvC5EmtxZ0rrqZ6pM020oj8MUjbQX9xk
Heixi/RtpXWMvXvGDWhmmEXxWUjv6Vhz521UrK2/ytenkKiiHsBJqRI6lW942eI54JohyOq+C9bo
w/QW571uGzMfCeIcMMgYJ4jqwAawxAVWRmBjX+96ZhxMenlpEstapdIzku8desdrML3pCUPL+RRH
aQgP4rzi+Fq3ScGctYs4E6t34zXKlEKC7poh5dQfKbJ00UOUjSH6RGINr126CrGzl6/yiCy/cDT5
ACWHw9PQGBBVObIQ0PuRtMsM0AFQO14PlR7juBR3KtiU+kIXBcI7cOD26CiOXqsfa+yxeURz/ofX
PDjyY0QEK8kt+s25F/ORRIpSlI/jxpsQV3DpM7dvhs4N6ozLhKGBjpanu6caRGBRZ+/qOjgUd2Qe
UQ3TznbixG/jQVGS7DRIFpvKglbLom1PC5hrBekYd7ul0Y15NN0SMP7UUyB9T1/5rZz1f3bnXpCV
aywVBWoJb1zTZMii6uPAtbYmym1urqjkFvxBxD/TPCcJMcxWBJSB0twWCU/sPycCBrXGRJgc82/3
A6wvZBGWj6+ChSBq7AYyzMoQ8d/ul4kY0vT/KKyiM3NajB+CM2ItfM3fz5TdL5rcquMj+zmm6mqL
GRAEvDvaZ6sMn2xxjjqVCAKF9Up/7d+Ao1EJcT1vZGsRtV5K9Lyyj4lci8uBL7S4iM3GPFU8T+7y
+L13n0pMhUivQOgKUVI/PttsONUfgqb2GWa1t46pXcNxYGS+ClbBMfKt8EAcxB+xxreNIiSmM1EU
bL+JF5wz5UKf6wAKCp7Vg9/G9kFg5pD+23ox9auPuxDw2+T2CPUSHjlBNA62+0Q7sRxvTIiT47GK
8D//wI8gh+K7s8VYTiJpKk1DR0zfsgha9Pz7x91oRGN/B8ZLpQyvsFtCIieymDdnnsYNqHWporsd
wRVoCmUU9cR8iDVRI3AV8s224BpJL1z4yQ3ZvpBVHLaBHLuqJftmtn6pmlqk30Q30UYpiscQHRJV
wFIkXAqKQF5CHCy2reGvQM3+iRFyaDSLDgbMsT7ykXysUtYEZnLAcPpjY7osZLzUMaJCDyZq+KIA
bl64796tRygJeg+C1OB9FkkMhVp7XHZEJ89jmcnRlmoumzF/W2uJm+ONpMhuM+AcJto+jK3sdmvd
sQhSarxCQwLxJepW8ZBe4qk4i5el3AaEZBxLnWn6DikP8xK50qnVTpFknEw3IA2LHPLcCek4qxX7
7rGRfM6k8GVdS7lQNuuAYjN04HITLEwGqL9tzKfgt1Qzs/ijD1g2BBeUTIaQbND8H9jCtgRo9k1K
xoc8zVivg0OZmdK0UTBeMPa+ZdgPqvjrYIOcw62xDfapjJZjJvWLcUmkCFrmeH+6o+ym2qwsfJhw
+RyMnEvFJeQq/qzJSci/mZnUb0xY6IwPH9u2NGDdyA0tWyLAe9OfeT//BVwEPJz8nWhDlambrgJx
YGj/SaOF9ksoXZcnZpZb5ydjtQMuAoPaGvYYx0zpQfRaOTkKhJVQQWjnzqocpwEo6lJDgjQ91ui3
IL7mP/Aab7skbU25frD+QcxARU9WmJfwx+5Ji0JIUrVw/94PmnSy1cv71edFfbxfjWoAnVck8bBu
t8iLS3KdjOcuXXoNlJywM5PWbr2WTw6L3DqqOc0ak5O8q9E74/EjII5IiErAIg5QoFRXWCXMJEBC
VV/1eQ7dfMManaimYpAfFoDU+0VWkrOY20aQRy5RsVjd7Z2oaO5Ez4CulnWsihd/Y+rye0GysAK/
FJEkuebXlDmCQYLoX++ttt+1AW03zvnPDlf2VPbv5zxaJq69k9jBXfEKY9Ve+KD3blqDMiX21CYe
XkQXC8ZiEhEQqiYR1YAwJLKHoPej92sSqwWd3MxkLfhuFcraEpAm5qvfMh03yHYdbNpgjBSRtmRG
sxqw8NLUjVo0CseqNurwUmZwrnO5tSPGdLOYkvNfGF6m9JKwkxUlPO7pSjX1mN5i59AU2chMKmm9
YAYjQ39zc3CxmEdR6weBgLPbOdnOQpbsjcc67SpHgMDQNU4axVVbNOR+VwPGhkyJd/NQ9gBbVD3I
WdsJr5EKsj4RSMvqHX2DnZuWWy/KAlBi0gXRSvNbgNy984O1AFgMFwLc9/ITOt/S6XvxYI0P1Xow
nuHoSG1zJIjjN0cMyh/OULJo4RazCuuzWQeqP2ealjUdcbb2MpqIL68SK73QesPLNSJizVuQM69a
4KPg1AxpedsZBDFwulEB5bd2h72m5T/sGMwOpu7Io9YuwnvAN/4Y0p6fJAC9z4xIYXKkEMO8gxnG
sTLThYFdgyR3RAJMxh/CSzJRmS6++h26qqJpWuyPC3GG1IbKeS1nNm3597uL4o6haBH3n+W7EpRg
z6jDv/yghqFhxy6+yXp+gsw4Mlcfpnfs6lYOb20VZnYp6eCU1WuYnfmauOAlsceKJRR6yq0OyUXO
rtLVSyKoLyRtcKJTUuV/wKs2WxH9mK0sZVpQt8izJ4MjpDCSvL07vdmhjIiPBChMhk11sOpkTfm4
VdBItrfXTgdUlSiY7a9w43za528kQ9WtzlXz4vhukfqUYkWfHY7kATJ6T63N0fOksqtJDB6Yl94g
kxGuftntQJ3qdFuNGPXszc2uAomA0RIyrvM5sxDCRvMe0zojh82TY+lSRu+l0xkuCqHAq1/cXQiO
F/DOHmMxag4JxzzqR3ERNHPVKmNmyztZ2Cx4u1sbWvQIphJdASxK5Ik/WIfNccA2ESQqLrf3LUpn
h/OcIgal1MuHzwVAAjfvgQNfeddFTavYuaia5Y5NJIdorqxD3hLz1BxzTbrmN3DOvqaBh9HOt7ye
lfjMukQ0fugQQwrGrw4/MdhyXyhJejiBZsMW+hSdVyxUpyJRj13UjumZMJaAIhA3H8XaP94n4amV
Mxb6OYQLCoRPjUG7EcRm79mhkXXbPUVC+aEWod21aZZZLK+0BWYGvBzsPFPbVaPbnHAF0vteOCki
nDase+8EnLmNus7JmnwkgW83kMeO9H033GF9D91vUfBQ5YhnGMpARKrSbUVVlXqWfCupUH/Ou32m
sBGXGUh1zA3gqKp/S8gmL3kcSnxHlrHofTstSqssKLp8BbsLN/o4Jrs+bv+bgQWuAyHPBuvq1x3f
ZhA0xHHVtfhpcfUXtfHcyYUjXgtPMDRYEs6W4CqfaeLcRoI9Wm73ds6pPN5oDWA08eSjZ0UZTIpc
dijjyUe67bTDqDr0FbZJ+QG55Co8+aJ9DiHyaL3wRhrS745A429b90LzG+sXx5maEj4MqMNAk+2c
sGbBkz8LHX/JsMFNYHleICXxQgPfd6JF1z2h8DJ9TOoMuQ7h7ZOziheamQ58hV51qBP18FVkWUO4
/1I2S3an9fLYlSbINNT6C0qkiq4dUrYaAULm09UabpA0QmU4crYyEFQxwjf30/z8QJc1IyWXpxnb
tef8BKkY6nWs3KtCsY0s9bXT+aBLCcuKb/QdCVce7dUZdMeULbErbtp+prOMyqlR3TDbrmj916/F
2HiQulp8pOjWxy1HcZM5/WGPsEI+BsJd/s4MrTTZ/kzbeMDb3TnjGGYocxF4A2Ym07EXiWheuNFQ
egeEVPZr3pdoh0VWibMPFGjTF0koVFARIgRbh6fet5bfbbEyHCBRg9ONDd/lRsoE35pQxEiVeGXx
juAbZqDtI7B7pg6N6iLU1ALd87OR2I0T0PUzN0/WH59DRfbNUTRCTaVZw44lbXkNRDkcefsGwykS
U/daA2SSk/LjNeJtm+Bm+NGIJezREGWKqS9dCjcjr7d9ga2Yv0cP8fmeYtDEKuKkxwgM+O+fvBhF
VhmOXkQTnxURH6pF9uSxAvWrpERzDqArUwOkpuIprgzDxv3Ke3Rr4LkQZYf3myuwU5JqFUFcgpNw
CBA3wvlsUoRzD+ni2h41Ei1nbsgbu1JtM4204lKMZ55WE0MRK6p1V6q46z1oDdZiBMTYjTsl7zLi
4EZpeYmHUNGg2F0R+sLH70W+71AmN/5gC2vDtR5lGq6PjO9J17qiuzSde/0wQ2q4fu9SRwaXeq2W
jPZhOswl7OAu9K6Li8kubyI/1slXbS6nngye2+tSAQ2rx6PydlIO+Zr+57QHu351Q51prFX+3Mpm
V0TbplkkSHPnmESzh9ra1DYnY5dFfYUW5qtcjdZWP0RVxAzJpiTap12NRdWaP1MwAwJY+yTPgEJ/
H/QAilzfSY+JSR5aFuPKk4ZROdDMKKELFeFokO/VlFqvSr0gBSbPJ5cshaqCVASM8EClOA9FItgB
q5OYMSEqkHHN4uUee98z+VcJCtZZW2jZLjLhYuWXX9AmHzEx6tK/sg9oECFp0b6gHixL2/8hJ4DW
CpuR8InvrLKx1u4/ZvTnNacKiotMNfjfCPRSr846nNxi2ZxATprkqjC9EHsUZEDyjTZMRFW4hXus
w8iyzJ3ko8dfifkWRi5ciSUXQ9sf/ra8v0kW6QwE2kKVLKfm0dLlyNRztaqvP+LteFFmiZs9R0hW
iX9Z9jznrL20KL3b8R0IrrZhEoxBS6akACp8HQk0TSWMVcZ7lk36oJp6cEWE5fPB/MI3o1deu4QG
7t0mk6hwdQiub4stesM4K+9lz3TdvENSM9gjyCCSVocxRW7ZNS41JtC1m07k9lm+nnUBkUJp5k8A
McfYDOpCn/udtwUlq3UhWSRmbwzu/ygMJBwBkOCqhYRmIiSM0LgEIlkSZB4XxQHwh009+y8GaJ6p
3kFpl0l5zP+2ABq8TZdwyyzkqu6AbO8hHWX+SASiCKTCVqqlc1GuD9ekDRxRfXSf13ekHKdqjH5R
Dqs8tWIFKHxkHElknKPO5DIduXOkNOk1ZO4TjCLeL7WwgykWIIvmWYN9+pa3UgwstFjDqHeBxqeF
hxWcgTTfPWEOuhNM85yNnxSkDOKUa0tnsJCOZmwf2rl2R+/c7ekK8SgglJu5fe0uPWDucXhOs524
h4r0fcG46/GyE9vx22w3Nfkb48hkXfFPh5AY1T4c1wwZr2yE0aXZm32/Mc7s9vaKjBrdSmyla4ag
rMosdgbWe2tm39ADGVmCOQxvIi8fqmLt+UaDXpwrskbPl0jGuxl3uFY/A5J7AlE1YlPNyGcJqgeP
TfD+tAUqghZ+7vUkX5llNZnAQiX1ALSIvwWeGLh4nlIMU4M/8NXNHNqcg7Kn/Dv1vzs4HBHvBPUS
Hxj8SQVKGKO9IMwZ7fTX8PoBm/NBj/RN7AwtX+cq9mOVHyK1j5N1xnFyLshP/hjYpb/lccisN7Nl
2tx2fhRFTRl/QQsZ4QCs38SsR9gxR2MBU2H4BjzzOvCkaXA6AUlRqk2FwPvJ8VSu5TNd6Ngz+pyH
mcwxLaZ+QwN5GDEqq1llTF4t48SO9PVhKtUfGGNwfvzHqIkzaxADWp7Kc1FAG5aZMQz3ze83CZlK
fUufvmxHZVtcNPYqiZ9PU0IjPIq+rCMgjyxv13wyffQxjJ/ij2agv6BLqrbRc9hUprcuaN9z8juN
lJPEIpzPMa5nA9d5qOB5L2tKJueByRudkCKsxja2mUoaZqIfzOy4sI5TTIdV6FU/E/WFHT7xWKje
cPQcI1LQ/5n94cs1P6AljalLnsvHG9SWfYmAyp8wJrtBCx4Y9RgurG231eZ1RZlz8PnkCylVQNSR
EM9r32/TzmG2Ce1uPoAFWFE0bGBgzNCH4Z9nu05R+IElbmw+egvnzekpn6Vo8YBVufE5/n314THw
kg7uCvDrkHUGb27kRk2tbSa/RLB+drVqkLG+zhg9yruCuEMLvqYcxHLLH/rlmTlLjS+3wLxAdrWR
DCXG6a0DPREDLzXb1GBT6jowkM02EPrRD+kILebFR8kXuBHPtPVPoMhZZABi/OqURNRflcyurPiZ
IDlPQ8Tnk6aCsWXgC+C04+iXedmZl8/XULz6Yv81wx704fsZedobSLJprLI0BlIaEzPbsnu5JHMK
OFjbu/ujJvHz+IgcrmOFsyDkZOtI2bvvELw0yhTVAVbFL2b/wC79kocu87PZu7YlYKZQip7zw+4j
m6TSGOwlFkaARpjYTgyCN74GZPXNeAES9n/w4L8ScMOkQHJvih4s977qnCR5NRN0dnEAiNzEXRI2
aUE0Np/25CfxTTp1QtmhUi51w3k7ELcaROD+gdhXvjFIBo8B/8apU9vFkPdm3n16NAe1ucbFx9hR
Dqlvj5mh9yd11Pe45s11P2EIhiEJiuIG3fNSTm3fByg6MPGMnRVuidpcMNapJrYNCNaHoxhOC38T
5xXXo/Eeiq+GLfixJJ9Ih4OJVzUBzmARa/fE+FaCO2OpNeLMhBoVyuq2PeKNxBpUOc12ELbjJ31x
N+HpFICnyrr1WEwfnhdmR0K+dyvxweDzZWCpBgoljDdOKBMw9EWnvZjEj7bf7NfnVngqYMrg9c5O
kX29d53ur0uYyW5QOwck7yH94UbCK72O95KMu9vRpR3K8+ZTcu9a3TQ/4dEc1HUxSs8JcxXKEnEo
LHdnIxplsdTqnJ9C3EpWrQ067Ch6PZC3sQd9BrGPJadwk8dBGSoTs1gYe/q8nwIbgpczYdU8oc6Z
KF3fgHhu6y5Uutout4dqYfM3EEa8lP30kn7o1VtkQimtsttNbWZQtHCWR2hCGyhOYmvn0U7TT14S
J0HocllIVnFe+4amra3FoJA8jddGaglevw/z8aEZjB+8AUn+ODFoQXfo+6dxaecSzeAOI4eD7rab
ax3Mx5nREyFe+upeeq6QWCz+A0f8J15sO/7Umb1rYsi8wbdvzBMJ6Qr6YI+ZF4NGfsyphDjL516T
iDaCWeTCryrVCYObOx/3d2vINQV8u18cp+DLnvloD6VFDKVXbA7yoosgZ4jl6QX54PYxPo23vooY
ol6YgxXt6PMxtigTUjXc/APGKNvD66DYYv/9AzH8v5NUX3ueLyFFvAk2tZJJ5ga40kUrEhRJoFb+
0SyIeYnZaKXFmnw1ds4vgLM/p+eDR1xQxwkYCguNi2xLRpF3wwsNUKRFPOzeiX4EaNoVGK6V1hYi
+O4gjlMMpPUPWKI5WD5SNOegRK3SzsnrNWF/enQJ6R4K6jITgalqOfo2Hq5xMP86yfZidxNQmSTZ
cJLU33STg9sX4FOXKG5fHZadxhLPtttCmt4xNQe3skPkNzsWJfAtTTi7SzQtXuOvRtOmXUPVYFhJ
KLbreI+VQCrOBRnj90LxdJu0cTBi18ED2fuOrms54Uz+lw3WGbHEwGXbb9MhCHH5ZAe2itQ5q7hf
TKqk9CKwzqqYRVH3tAxIybMiyX/CZP/yf8xgq0Sgz0pfkBVHK3vM8Px2RX5aFeX6ej3q2gwRm121
4XMiRsxLLXziRGfpda3wToGeNuMrPqmUefgYjclSh1VIZCyVRTky+ANli8GqzkTnya6G+v21gK5h
x4WbTAkXs6nl/MPwPDWNnfwOI+hG4tJEPirIoK5KSG1i/7POwc8lNVavplO8sU+79lzlqrGwKTj6
In6SbAzrb1mbPo70tDZM9ZIinDBWejPEbwuCgcrlGnJaL8MQlP5EkRRWCe8mcJELrZj5mSpGkQYu
+usEifs0SkJuMEonIbEanlsrDayWppNYCAlqBCVnYxXr/yxYgsy5Ru0jfYn8sVmA7DTluSrQfPs1
A3wwWRRzDApBVV7RyTEv+o7wCOLWFhs5GRYYAv+1wgdJVwMaZVLNwZaYxxYBJXjHQXEWuXeGcQIW
fj6VW3TUlA9mBx9SJIQ4/6W9qzbUioO7PFNayPL4AdJ6YRo1AP5NY9vQLhk/pY1Exjzen/ptS8z4
09mp8yub/CsI0Fl88hJDRTRbRhJtP6W0l+VI39z4doGbKYhQNjeMd5xn9lYT60cWckebd1LE7HKD
n4RpGIngNbGhl3YzM9nFtA/ffmMFBdSpmPVhwbWc2smBvrm9zKroqx4TTDK2RaGQHrs1V3m5vieX
lecvhnK/VjPeRLIsGJGlRB+wreSeyBWmRs/m2/UOCEV68e4WQaklFceM5u/+iCz5gZCWdHAn+Q5k
VGbb5KVp+cWkv5lg1mv5p6oldyM7fKT6f93nFpNfjdZpMdgIVpmT1vnxE+Mh6vwxUUHPAs1aoP7z
YogrKS9Yku9GzoL4lg5SXBkQIKbMH0nCjQyO3G3qP5961rCWKPogeY0fYwupbAs5mfxYAUaZruTz
+YSn/MMjFGWAEE5I2gQmPDwrXATbEJ0F/uS79CbIr9ww3M8Hrq0/7lieyWFc9pC2do/4gt32UjwL
pGoOKINyOz3nZ7PtnDxUfrty6j7vfOAcJ0wDZ9OaEsGdnHmMpWQoFm2xEMODENoC1UlGs326EKO7
b35AlzL3Z9D36dkggT9c4WZWBhklMIjR/f3qbVudY6S0X9gIjFR/9zTC81nFLMoiC63BwDYW2sVu
6muIz6L8i551bxVNVRGetMwiAUVzDnapxCaTDfeDYC/yyy7tl7euuD7+bFKIYyrtLfrcw4anal7H
JTNOjnk874N1Q7cE6QzMh7RfDSN4HCkk3Kb2mCudwYGB6iIa4dbcOerV4zOFhxXQzHh04XX1904F
mpy4xYJ69s9j1pM/an/jg5HjduIRIzBGKdZC7kEA2uLbEkvf1/lxFoYG35JId0OiEQp/FnXMT2dF
u8k3a3D2EkFUTf936eLHST1kAakVdcxEIwc3L1P/aF0hs87MNhlp3SxCS9nLCL5pk+FI12WJj595
sfP9hruyncQqjSN9Lou0LtFCQaZY445X8GcibROtT012TAt6as33mLC7sXAmbaEBN+1cwHEYEDKI
arctr6hQmV9NrVplSzvlrl/MYpeid93noA6g+S+JcGErawc2DpbUVjF/zG/0GhqX81pGNqL1D6wd
afUs56LCr+5Q4kn4PVqtq027VPPpMzy71GJIrQe23wEu1S9iLGBPgNYUXpF4tsrggBOU76kCuom5
qF44PCF4HpOqDXgNUpYjI4dMt4T61sQRCmcVVtOuF+dhsSmdEaCvN86TGN5yVk8JN1NFg1TsNZe+
ITsvoD4mzsodaUMzenI5nFxSiWEijSGEvtjiZV2F7/a6trLGxfgJZ/ACDj3fnSmIM0PdNTCLTAt2
q3HvPnZ0FMy40/k/xIy8gjC7uy6eHpB3uqiMWHXp+T4WBGOdSZv5BdYtSYYwXPWO7/Q16bPeWVxE
qy3DTHveFZU+es7q7kTyn9LutZtN/sbNspypPx3KvFs/ftWMTCzKcSAOmslh2Sji5o/L+pMfj42O
pSYnFIG2aUmPNzsAgi4VyrPHsAl8Ogx1WJWWiwQLo2Zip2gGZgh+RljrHVnzgnMxr8i60l+ROSMy
Jcz+ncxw9utYwDVops9wJ7WXUlkr075rSwlWGbMQgcZ750V01Ler0SxqaWEgJ39rXsAI6gVUmhrH
NJuZ4PjFWusfvxG+uvDRVLAjTvM6Nxb0DqOsucWjelHgoQk1F7vS/pe2QdFcAMYbUmCVySTNYXlu
QBC1TC9zZHgab+smRZiVRKTCsQUNy9Svg9zbPn9qBJcv3TVSUj4H//+crNDHl5aNUZXh8790xjOo
AzHhdRVMoAq4DpNZQnQzfTUzlX2d6ObYI1hhzH/cD+lqdtGdW7oFtpXqN8Imud8THcHox2q/z2m+
+QHJAorFR3hW+dmT3G0lMA2+dVghkHTUpONLMMA7vScBIV+1teTvb8ZC4c6Hi8PSo1j8z5yLSZO7
8/KgRocaKvEgpzfBYYqXKUi2Jqy8d1MrvMnS+rXsFBKgjsgau1KXNhU/BZSHHkX4Z/c4xO0sdQRG
T2tnUeAvdzvbI51maNj+NjODYOgJVnSsX3zhsaVGilUtuTfp2y9dRsQn6oQiZgsfA26nlRRVyugf
8WBt8Uhn3oRgySlhpIcZGVpW0pUJvGy8dfNJHZG4IJJZfzHGqm6rb3czVV5+Aj9ce143pkwUO8fu
tanlSWb/99bOa66exsYP5p6GufMFcPGY02yCns7zuHKwzX2EdWkpSukkWPdohjZsmZO1gUYQs2we
WtA7BjERW2Rn8BSDETX+HTkpz2kU3K72fFmkCwt1ObH0SLVQq+r0ILFg2tvkRCys7vNiyAdB25Go
XWL1GnwnA993/Th5lwIhiQnxQwfp9eIZkVW09wDXS+diBki9u37VNunOi70mGXawazJMVB10Dvwx
XGt9i2voepyE+2EB8lOcKis0sAZqvSTnZoCpoFh3/EjnIFonxtp0qqxSoLUYqzk2EUnKGpI+WhIF
7a2QmX8JAnxBEX/kpmZnDdVGk9Q7k40+mGRX6Bkc/GqcSH9sX8E6j3Z6jZ/y1l2c4EZSyiCI6veG
UOK77Zff7ribubojMcm9ehGzPrZdDIzBB6PNFCeZwpj66TnDHwyaI6tSw53Q/y50+k6To7J6Yh9R
rKBxhHNyvgOuLBB2qjdcrUqZ7CGHoDBEa93UWQi2dOWkuwGNV5K8G5UKJg2BiP0AcxWn1vMUVUO7
zkuWvwNivXE+Nndu/ZuhpFA3P3JG8DKBKFZDmiBbgcYvEDO1cHHSGLyo7LxRohU8xGhdjYIJ+Y4k
kWkkqvXn04FOvXZLl3pET/I+NCLGMFTYdaGCQJLPIOck9bRCFZ2S45Jk8DNHENlx9mAde/s46u15
K0Yr0oN9q19HhH5RwT8YUAl1PaLiCuH9ZNtAXsPhesw1dGU7buw2gk+XpyhRkKPMQit782SioSDH
d9is9T4zSuZOOQAWMa5nxofmt24IO/B2M+nDLuvkuf/Tbm/5V4ctNrXqpfwz+S/AOZIvvXDAuECC
qS2X6zfzgmlec8MVuuHIs8ORm/tEg48dbs/owmYkKVndHIuwL4EwiE5tkFF9B6ZfiJvASAup2dck
mlAPGHkL4Lpi3GP8Lx89L+DVlVA474My0AdEYtIRar0ef3cCqSyTXy+9ZysywYGgQmMZlk8tAvZq
ITojU4Y0/NwoCXKqLozaDJwBpHNu/6m6kgrcbjao7nGbueT38gPpOUlS5jsh5wgEctXYGdU1U2TF
uIrUP0pJ3IU0sZLEtOjmjyNBmbjmuWNHu2txslHY4j4bYkE9KQ4n+MzjPJdRI/LO5RYV6dzSk5wx
GHZD6qI7lc+BB4Xg10VIBp9m60VQFVoNrPBozVKBokTG9rE+XYc0JaySkGe4raFjwTpUnoxfwqfy
7QuN9cZenbyRyxedXctBPlnoOVJd+eq3I2CzTeLPOX/nT2lEWL+yU7Amt9E0ikWJY60tPQs2vLkj
9NXsQ9K3j3fNWKRv7fQh+wOWVopZDU6ohQbJT5jnOGYW2RMXrh+zO/0y6tH2xsNMBAigx4jrSquc
S/X+BfPOnL5Xw0mg98rMF350bC2IniUrKprAMhJ0O51EdF/0CD4v8iNiS6yo5oJ4J34VtNui0p2u
OCzz4p5zPeDe31f5PbgBC8KiOaFV1Ct5U6Yoi99+ccdXwYJagA7w+mr4zrCRRJKfnAotnTFFSDyM
gzZEu2aXVYsdCzW+S47VlEEFOfKHCKXDSj/SZAOuQ8UwR+pUeZM3kFdPTp08fLveTSwBKsEJzMt4
2rZTZ9RifQpEOPHpvIl3tBbfos391U8ZZmtOBp8gd1UN6t6PJpZE5/PZQt41O8raaqNZ0+zV5ds1
+blf8+b558mZV9voMyyguWCUvHMU8BbOQfWrXQmda8i3Z3d2Njo+D/g/gG3vWo2WwKt+hCZnL31p
zntBfRH2Q9qcugsTYF8x42MoKjOmmBrEtsm9hZiObscDMe+Y/skm5X64F07o0LdxvSwbCud+fRlK
dsctnlsY8sjjhjEnn/7HB/TkrMQlg39lSCBrYK5swwKoILcLcM7SyD1f/4/ulECPB91SEeB6zfv1
GzxDv5bphIw/UC0eynChq0K6N8prlw7hlAfifXpD6+4fC8Lsh/HhYU5xaob24/r/imv0TJykK1Qo
7viEKTX8ic5hIX4P+9tpEMSR0uqfE3gRtqmS98P+A2//04QbxKlwwftAHmYpnjSHeVoo3B2XaHAi
WOIYFMdSgusGVNtar9FHm+wug3w5iHAhpEwaFHsiTBsvpH8f2Vqj1n7+XbW1rWAzxTQnioqHApiT
ImvwBki7fPM5Ot1OZI5MPd4eGbKEE7VOYy4dQNu8WLxeCl32VUu/KlV3Z0Xc1bYs3E2eBTt4zIMc
EiyYH0tdILG/VI2KQPQoIBTMh78p+v0L6WjGPWakJYCA4enROIkCoN9GduXbR7HdfHFSvU5kOJ+M
ySo/klSpjuRxCWF5ifw4ZVFgjOxQvJbxp5hQYJFDkfxe7874gbb/1wiRh40jkPdWl4M+pdIOkhwn
qdpJIvIUvAPzx2+UQCec+a6hyTiq9WisMYzB62pcm78XeeTFpsTEranFeVdHOCORB4PlJAOawKtP
eUCKLCwq0YB1467RR2Cwm2fCrrXLYRv+XE42hJfEkzxSic2H8rxSaaV107eg3ZjVK7eL9fL4gc3d
GJs9xGB3SbCmPqkF2k8duElfGorjaSACTZ1hlilnQzByw0B+X5qXA+TZTNktTpePNHo+EQ8KImyp
Yls/8ElhsPWjrKZfnRPZ8/ErPM4Ltbg2n4hVt1PMAgFa8ueRO+a2p0XFJJVuAES2T/bWq0KioUe6
MVJka6O0X+tY2M7z7hHTB7y05SmxTD5FfPZL+a9IjbD5QcCnOsXtN2HFXw1Sp39ptYvpUU+Gnasg
W7BJO6CWPqHQS6G+DXgYY76vDN+SGifA9HQYqEUJ9y/q2uCW4PmzPI5ZHTZDcdksqZFXii8FZWSU
icwmEMv+eVLryrLNvgkJaLkgvBfpQ2r3DDRn4Bu/5dkLqLb+ZzJceDdIM4Av87XlQdSz/1RHz/Nx
JFZB3T1JzQFccnWyCsEoPy11sxtOS32Soqi4DwQN8PIdiTQyDgItz7/tj5NIFhOypwpGtaO6xDcv
HnQpPItKH8083IhB1XXYr8MAvWjaUUQzCQXRNnKqM8Fpte8itcFkxkLPkas3Qh+yUSwA+lYTABW1
dtWAmn4foKn1s0Dv0PbURoQgTmP5XsnHkpsWjNS+qJfYr/ccaVJ8dKAmMHWIKfM4TkzIE+9w3imb
psNma0bSNy4+bbvzL2oxbbL/IHDnOif7XLfySwrk5/qPaAeujz7041tUJ0nmi4R0ocHw7CnJkV/t
nYj9ObNYOEr/zJjqEjsG6x54SneqaMXJE2zEu8tRd1JsXgkVO1vVWOMXzoHZfVkpMEWGJAoWbbVJ
qk5SbK5WzZ+Iz0YRkVp5UhSJJ/7mm0gEKijanDZ0fZ70b9WWDrSnulGWYd0gUJCXctJHTQjicF21
epxmMF5czg8cJ9pPholE2feCKHpkPkcdTorLWkHATGaNqH6CcDoIjuUHrDSwOgRyXJx25x5+WB2Y
Pnm406EQ++JiMJh8OxCgUK7GqWtM4OT5d47ooomzxbnvughGWFTOuLYwpjh41qW5DYo1EVoi+twX
tDbdn5sdpWko9okVhhsw46E2Xtk2vCyIk35AK7ApnIo7v55RwS4I7e8iNP6sg4Tw4P80ltNyWxhn
ic/iLVkFqqVbgIfkVSfp8vulqJutDnX3AN2BsmQ4A4SoB3mFo/DVoCV9zl/tB5YilEe2kCyCpjSv
ZltvfV+LsRom06JJuZaOIaZJyk+aBXAgv8d55tLXohXFS1tNN6Nuf9FH+yM68Qo8SQEOATHLt6Fs
N+GA01h6GsgrurjQXcK3FA//2tEL7xJBrPqBoJN0F4hNWVzRl/SG3+7aLzMTRuH0pM/gyV5kmF17
vEWmMo8Z2uVOqDqR/JBseWulpfSDtfR3aYlZHbFUMahOADBW9sheuApGazLlzPcLhxzs0HnpdwFF
6KnsMN2+UyUdqnx1rn63XMOvqSr56r0V2FF4ypaSto8hDBDoFJfaz4hXwIStYo315qNT9TOzHdLB
mN+/ZyhVc8QEN82HGPGhT1TbCo5fptshaFhSd8RPeYoVS/XC1yerZ5VQw7QXauZoWQ3W1eaAONiB
bGIfjbMcT4Hhp78xJo54xjehxbksDkEcBszt2hGhW2PAFp+NZejMbwfvYgd6rHuKe42bMadAEwAd
l4U8CVkaPJ3EE0RwoTaihjl0gKs8wOZlkc9P69+fGEfbS6czVKahem5rJD9xPO822ETXGRn7s0PG
6Y7zt2hybZ5bKcqkauzlizPRzez7NyaQvSsKhGieccito2RbQ2h2Z+/EsK2LIJtObseyOGbRy8g3
AvCXcElwikgo55/vJT3gYoGZILmsOLik68oaae99lkMX8wlAdWc8dvaFHeiFkG1ac1uqRTmw8Y5d
prwjskcI7fSNEcGmQr/isGU5vkYKSCWN2CveqpHoSPDsMWxUlYNw3jxKB3ka7a5H1YCqw3i5f7z9
6ZMFPF+jnazyrXqjvJe6ASOAJpXzJ4p1nb+ar0gbHGZgZm+TgSQpK3siVhs+ix5XzQw2MSEDTnrx
RgPTT7ZIkz2R2ghKmibVoncdnKS4gVIpWWAC/lDhVgZwTME/UkWRA/nDzTT0nOJvvBvVRryd9Ei9
lVB+6JVOjFOG0vKcOGHf0OrnBhgywaTzbnas0UHFnPBrCXKEV1GoVN4HZJmLNr8Aa923sWnDpCaF
/Reha4t+o8vx4rhwBgQAOOrUEY3xWshXSNvHKtWyrM47K8C8GSQxRie3L0preH43XUa1hYezkpCy
C4+6Wy2WvLBkWl3ReEdIx4EC5IpXfsJZ+9g3EAmV6xIbnYGOwsKNEiIkp8rfw7sjvo3g/yLwl5Ae
QzwbE3xPbDGV4RNpUZfz7b7tuioEh8BcqBczcGo03xwpWAjnu6Sqhc2M1jlh/Ah5C1l7IZ+os9Qo
DqTZz7EWT4bCqUbCNnKM+OEKi51KxeYb+fXtwQtdFeZSuAcUKG9zOjTfnrBRsG5M5WspNGrsRdVi
U5NjWwO3LYYdSMhd3TiB7L5Rg3aZ6yo+yp9WJCza+LiMtnimCp6FPkXKLx85nCNTQwuWOMFlQ4IN
1JV/6+/VOcohLe8TJ0T4kFmq4McMLg3IUGt3EIf/z2pf4QMX2tBjLVdMie+m/GL5OzF8vl+5SbAM
WeHGLuMOjDVu1YAoFg3U8im4g4JMByvEHAyDHR7zSomDErNQszd4JwHGb+TJ4NXe1zkx27BZZ9nS
0p1Atgtx6gwp1Re4TTcJyJFiAM/zSaei2CvUaaPcy2uRVY0nfaEObZJP1LdKYx/oIexc814rOlDr
Kr+5c0VbF2EMlCO4M3feVpLCMecBJuxi5bp7BhcLxLtX35FBef5SAdCkFDbRkjdvgZyoGG2P35B1
qqxg6ajXhfTpeXJsY/Eezh0g5tRvhCGLvXDCy4lpSyJXbOxz0rrdGQ6aOfjqd9O3h6KNFoZoRGXL
Dj8IOyY42sUn+GADn4gaAJOLIWVhHgWGuElR/wbvYVaZTDhL3T2YUmg+YQ8hGP6H93p3/T7eVvop
55bN6pDXLolUDs4jg5aYvTVNsaI7A6LrTGFTsMsQtFt9GwJaqvIbQp1OdNSx2j6gC0JlxPQbezy8
tdvucyTtku2z7795/4KAaTP4inpW5Cik41TdO7ENeqxZz3SkrNRF8BagjMq2FD8CptUmCEs31iWm
+6bE8FTMs7sJTk8gaEc0NhgluMIZEZ8QBzjcNvBB5aL8awCYHB1i0nTbBNNQa0EENa+2A850kYQ2
Bvc7E899iqrFRSMUD4SESIWDxmVvtwHmzv1r+CX+KEtO47YJF17LBgADysUM3TrXVLozTNeiMLy1
fk+bkEnSK3juj7evB6YDmydSlPBOlal23Yf59c2/NMX36vMMCTSyXhkCIPLjY6lhLEX6SjpogTXO
vuoqu0I1d3JKYxCrJnDwvoKUI1VLQCTkCL4TXvbK5UBCosUHyPTZU1UHsvojTKBywKV3f3CbcBzR
U2fpF1fjOvm8A+Fb6iiPPrtqpvGhbwcHO4//rxIm6W043dAgg7BGebHj5lvOgxxLsQa5TvpM9hpT
MKPTT91Ixn//tKiLIWs82d+fatMqGj5kFOSre1Wz/F5xEnx2XTHtWiPdIvZB9KBCi532D/H/B3Y8
40EjD27WAN+/fwKihDY8pJuMuyzPb8YkLa6fm07wQPvG6Qxop9fbGZP9rZrrs8qqg+e+U27gWGLp
SVGJtyoAOAcyoHLwMJkQjJIn/jFFhGt1frHoBXB4G3tSvPou79va3wEIETELb84KTacB+XtS7j9m
BBDqPIRWH9P5kRPyp13hTuL3q7sHBjn58JHsDIyT9p6c+HGazKcwTP1C/XuMQ53vZ5AaLKX/rMUZ
RsgK5hjpFW0PaOCPwcrfwcJsEA4ON8J6B488FWNHyJCJO+6UjDmk5Di4JUQ93uItoZLXvwTGMfc4
hmmUOlaGNAjEE6nxAVJD7FYRe5zQp/yuInYUc2Qai2AodMe/BGu1fBSijWnEhtaAMqbLnUuzgk+Y
b12VC+4rb02sVHt8bONzO0SH/tobVb3P+fpW30ZLNwx5PibyvZAXA3eM/X5kEDEAxVPL2YH5yO+T
CHY7r4VIFZRbvANBAVgtAwh16rZ0yN5uOvefpqqyM5qR5mtS6yGdaE8g2kYp+B2OUvQipfJPmtey
teQD0TBfpwun1J9mB4PfMriE3azmBLkDTd/1MIJGiLEeuAnjOMAP1N/R+BAZ4S9Sv+fXnmKBSeaI
udOvv2uHfmN1mjeOlmrP+AT8I3/3puw1nzsuA8XDCBcJ1w24JDIeYf655Zs4xxCpJNySl6FU1/lh
q+8hWJV49ELHo2nkEOa5GUEJ0e1D+VpusYMNFv20w1pNfBQMw8v98eBfFfMkJN1CeWm1Qk5G3DZh
p1LxuPveqAlj4UsSuRyULjfzEc4wqr1TO5ehM/58kWf/F4phALd6VrWUab608tnN3evBIE9fIWzf
5jX89laXYjXBxYGVNllgrlC20jnRHdOwTgjJrNVk0x++uitELY46LHtvt4du7aFaLpl3rYlbxFK2
GwoB8jAA2PQ9VZunMJchh+LE5JFEmLm2n/wJ6jucGKf7q+6SeuGumWwzWHkGMrSqweqZpIVo2TrQ
IH/Y91otL7HoWpugooXAYUt1lhOj8R2fHm03w2MdKE2iiyJF4wXBN6SH20893aCzkiK6cQ/O3L4o
HBINqs4rYzNbXMXHsXxNlKXrjc+tps47JYFrXnYovwHFUSwkEO/iz4mDwrihAQ4LLreAzKFc4DeC
/CpsKCgh6EUUzNQx4Gz0yh0/OXF1WoH8tDZDNvet77S4FKGaKXhad5z3zV78E3kmJqGM2Tn2lyDU
31b+VNGKol2yEX2vbtkIw43kqqp4/8QgXUd7Ac1Xnd0GQE9MnzJ1x+4k25Glu3XxnCIDPaypB3JG
6A3xo7lQ19Iyi5x92VGPXiuUpc4ii8DevMgMXJxZ7n77bQSSD6O5TpAAo9QIW6mTaRvhZd3NS2X2
xZRAJrfz5jOEz7kpN5KwC8cyDkctiAgEUPF2tXXSIKiXLP7rGmP6ERUdQzicXEuZ4wEZ9LB/xJNY
TnwJPYrot64Wtc3Kvy0JGmBEL10PNeeGZJiXcG02csx42ZstWQU9c1qs7mp0tOaHEal+zgt9R00H
sWu+2xU01obF7zCycetLp8+LikAVkAoC0Id5aLnqPO5jCnCOl0lb048xvOwvUWeTvvdMD0SIwdvv
yvPHUnEwxFfSLAWG70in5qXyeJNYhO4G8pNpB3kBoKoxb7POz2jZvjiNWJqESykMZD4i0LKtKXsB
KguR3610rAX3A2j4qbMS6JdHWlBhzivNrOyOYdISdMDKz8UySmENjMZlhE8udDeeIyvkxcyNBcC8
b6pRPFkFdrTWU/5zYwIxBx/B0Y1LoknkBP+vOKkkdZp/CuQp8P2w0McOtOnPGeWdx69Cw0WJNP75
4BmrLHCxKgA6oN6JMnZNks0F8QvD8rpI89Lp743/OEOoSmJP+NFarFtKEL76Pbl++jMTfOjNEO1T
SGlz15wp/1ayvURcS1Yfu7IUOTqseBj0j/Vt+K1wrr/c+LIpxC2SVGjSbU/orj4BR4ONFgTpoY7n
CP1hcZLrIM43mmOguKeyt3NwPX37T/i/mKWsiRVBavpv18pmhIbmSyupHnNbm9zd1Alrc1fC/Bor
MsTORYrYNcwD/WrsOQNscM4YUCWmw5qSBvztwYBjLdpD/ht5bK3KJ2FwL09Y8vuhDQpMU5ulb2k7
WCLxkJkhnE04y483lPX2mSDCdFrkkDzGIJ296SFMfCWadAyz+VxDfOA+assCgpzU8XOKvv/2IQyJ
/xG4L5NAqnCnQXZ+h3ChU4gXnbAsjCSZtayM+yf0RC/RA12mhuv9xslefnjoHyOqsfw8czmdspdF
x3P5GEvWG86bAL6wzos3m/EXG/7q+mMCaRh4l+N2R8h/ghEgJ0ajV3Z3TCtXStO52czrqhn+Nvop
YY28PFI3DP2iF1wxtFAzVnW9cM0qSjBRvN6go0X92Er8ZddeWmWiXnRstc4j2cY0Hks0Rz+zMq7O
7JSeRQtCBbJO/b//VRuzRBV5wLmsjl3+vOuc+/4BMjO0vmCneGKRNBM837XY/x4kzSNjDnrH88id
Dw5DcyNBzmzKQdCkSIe1e1kQ0Y0eX97f4sCG5EknDEWx/hjNOdJK5bzh/z7zDx3o9aDNDNCdvqjL
LHuTijN/XFSTIEwXwby4uRlls7hlG8dp783nsB4pFLkeOFLEaVciWLAyEbzfpsBlH5mNiZgyNHEh
w9nBwe1eLvCZAGscYWrlhO9LK0CcRF/Z/yIg/5cxTXGPXQLW4t3FbsdBGXcOwKAXELW+yJU2ytva
2WMZh2p0MWDPJFCryDwUER5d71NmX22apdYOVL/2GDTa9lEjCArpxSf2Bd1YGtKH9yxzwI2TsOy1
XCCZKMAlxeC2mM5lbrzxiizlx2j/dMVZGeNZGy7WDABdP7sepAN2xMKBOh+8k02gnXrr1MYJFDIC
fGPEarYnPS4PzHogat6zENbEQUrgQgR6PLgMGrAJhEfRtFZSPn613mKUf6xd6Fuh2S7Xl2ZfM3yl
I7HXfQglEuFSOjdgThn42V0IGJLETLPP9WC0kgHVsBMHcb/q5sso2X4CxOnq0c2B8IfKTGKj0s9G
odcdLTpECvSEzjAxG+Rwq6s82azukGgR7gfyKhQf7LKXDDXYrdKBSYmbajeiGlx/JHfhHETeSKGS
eKcwzmeKX+UTGmKUfyZGbq0s/I+oTtO+MrrZRT/CwY/x1grHoyleCsdpYjsvyxIQPA2qM7ddU4zb
a9gRtZh1Ek2SelIZ/mEhJzG/ZzYhpkZ7HCs95wzEuptY7vjSFXki24wRSeXffAttBW1NqxHrt3eu
YJiIkuwhv6Kp1VSqSD4XWnPoIg1/LfbTujsch2vLelHt7R3ax8mrm91bpHXtUnRu2ux6C3d6u4gu
vwxBVISNZUZEPkweh4SH+f2xRcgYYl5ztEJD5vrPnx/k80BbEirkpgWISFHnPERhurf/WsHcDyka
gAQ0W8CKGVoEL8fQWDmU7b1/7n43FBtiuAKOl4W4H16d4kwg55kvvArkK1+1YEA3Dz0BY91/4yXA
QXvKvAb9FQAMbbK4occepv2b4TfcvMiGI0quW/3oH31WyLK3NHpk/6rCPyoX1iOnrgmFYDxRnnKV
wcs7DY5UobBPud7LYNzLiFBp9LI6lY7eWnf1Sr9jgMxACUtjj6/mQp6Xas+cUbapEBiSs1fN0DdC
6YUK1KLX2MJShc7I0gvNo8R8ewbZz9hI+AsZZP42XaK4+XfxUczxRTH3aF+xEIJzLl8awC6xEFRh
n7p6v9unUwt5dmoE6RdiMMrDC0d1gYBy2An+meZz588u7qDbrQByMk/6lRE2u9DBXmvi/RysoTHB
Ub/wtpuXHau+AGRiHTcdKH/3g+n+oFlEExjAFuscwrjbxOKEciMOccNFBW6ZA9B91fl+tJuOQGlm
2QZT1qZTk0iopM16Zswx5lBhQZqWkr90iB1/7fqzK9GJoVsBySlqrY1HU44/GGQCbjitHoaiSLni
1hQkTiKI9ZqOyusYfl7R5AXU6oM8ljLANWk29avY693hyyJuDwNO7jJYcbQPHJEg+mCuZSQTnkYG
GnRLcZjEdrEFu129uc2eZBtLvIKC5KA9r7OWq8DzaMjO5zr7tM92Ge0H+yY9mwwjSJTH607k9342
OhDeVHjFt+dd+aHaZzlZ3NBQsFDJFJpSFcOqm0zD8Osipefx0BWctaWzbA1lsHHGGRXHRoZm8ZMN
LtuVm3HWMsbU3j4eqy/NfyhvEeMgjVVVfgvHlZ/p740DzgP5eaj2kErxi1Is+yAhiCUBGss2h17g
wIgV8BA+of029buv7N5OCthdTqAv6jYa59oDHlYCNp6R5XmFdyTJ/ngAmILqgnA7zZahFet12lEm
Um22xY4jmEJsc4mUil50WkzWLcphSd3iydAJYb81bdNER+VJS/Z9QD+NLZFCuiN8VrfY8+M+BVDc
zny+9Kva8bSYb8ZAI+h7QB1M8I14WUyzF3krdf9uV3+p/5d7A5MgECeSWZg+u/n34coBGTzJ7ZPj
zDftTA4sC3HSz2KZ40x568eZyxCNniQCOMr4Yn0PE1dLFuAyJo1SOUQZPrbhJUnPC6+88piSX3P7
Nn1tMkirNpgDu789p91OaBpaxRfe8Cm3Zp8n/8PTrr7SX7qYECN2vmc+hp+Ck1qXfzucLGEr1Ath
aB9kqhdrvUJ5pfc+03WCFn9a/4bU5fI8OP1lvCGwP5C0jknwyXIoUeGeaOy6vqabPUjlVIUAW6eJ
139bQzbXW5O8FLKNae9DPIzLLcxOC80PxrnlSCcS8/y8uBo0TsEcpArGkipX10Sa2TZKkcqPrilO
K3puE7EtfKf38BMP1IG60XQBUr8p507c5YcCnBZsPMnykpuCZC+GOF8IJCSJDOYqyzvGVAwNOzap
VRQdh58uuAZV+cNUZkBT7erIHlQO1fsRFmxTqyH6twkKGmjhrhSIu8Q0aWfq2hJ96rjm0a8a1tPZ
W9E9febtp+6BDb1rqU7qWOk+tC01TyyqqmW8iY0SevQUZ3/wtPtdgtaWp0cVLoOBo3XsPaOaX+z+
0G6+C4uqo8X4ouXZkUr4xPWL4YWpDzT51rVLIy/f7OC0g6YV6s8VOJg+WJRlc6f4+/jvr66oK9ed
H12bpcmHVo0ocbuX3JlVaRT+IoQaElY+cu4gVnw7neKDHrFEBq7HI51VFL5XyoVtGW+O9nkA2n9E
iSKHoGxCNMF2MfrZX+1emn9l4l5xLdQKy1IDyVrYRIOxcOi37p/dxUMlbCUhZPgNn5Ja+h8/7zzZ
dyQU+K5OwxzSkcHik9buk2aX+5I131StgHhWkVrjIBCBqAaJ4hbLZRUCZ8/z0HmCTrCokKcz9TcN
QaC8/eiwdSUMHsBFUJH8WT96iXDgnxfPKZLI4pjVbc2dghP854gCvSKxeIBimWzZPDGd7thoyUAr
pktvBMGkYaKt6knUTi5lFNZkDKxDV6K0tdmq/dXJiU448HvIOhxWeJVaHA9CgMTCJvlRMMbQy+Aw
fI3XyEI2ZMkNRWx3EaXMmonpescT0TpRfN6eGBMYhfR4jrZM3TGY9JtUKZ7lRuUkQIgIiO3IblNf
MxtkACMbqovsXWNJXbdOJY6y4w3YpY3QY8FtrRDyKQaw3EChGEQyRMnsQTtlvhZ0u5y6Qo0HUJQX
S0qRCQ3qz4BQ6TF5H7NBnWLUkLtc/dihcHbXV7awOBkE4RQyIYR19FzouwptaMHyu/RwHfqKCSQj
AuxEUcPWJG/03ruPPycu1g8jLMZnhgYl4jt3zgobZHvhX6EiWFK9lLJo6z1ZVI4RU2DIgl+m7ZZq
yCSniA+Coxc1g8oL7GDQGv8PyRHVu6ePJhTYrrDs5N/fHjVAOytOQb9e5HNpDwLUJWsEGaRAytjW
pecBY7cl1rCFMyNpOnWeZdu9cI5lYtCBP/MrMXj2Gh4h6nPMxGZd0Kq91H3KcfrDx9yC6qvvQcsX
h626lv3b/kLW7Z3mB93vgtgBoJRaPLqcQ9XuEzfc5k4wWFIr9pXFdycW6Z+3acgkTLzWB6uqjY2F
UAonCzhFTRMTD3/KaWkYxLkMXtL14FSx09xu9UhARUfRORNMorX3QDJXG8ERqXxVjHhjXs3A7LI/
7fEhS3DS4B9ZwTyHS91kvpC1jy6B0IpbwF6jZgLBIXdbOsKxvjCFTGzSDiLSzc/O4bod6aSQ7N4t
kwCXnDGltWxV+k47v3PQOx7P5ERipSh50H8OCPxtme/eFcm97GoBGqV07UdpcfI//ftdn7s6ZLcz
eXnUey77Saumz7BgN9irjzTiVeHtMz/+lg3kTnQmleC5/PkqVjwsoO+PNXQPx07P3PL47AJBRzna
3M1xPGBAEzDX/43klW5rn2eqMNzDxeLGiXYsh2wWk2C/mAcTVk/rNgk2EJDwBZw5gHUmK5V8wrJ7
Jk92RZj1ry9GNmRPEbNHyYvgJbxFLIo1MEvuOuy1+MmDQQ6aNTIZZLlwaCcDPc3+Ez1ks6QYa10j
qCE5x9DYWMOA7z+aRSrcfx71wz9HxiqGIBfRPG5skAiso05bsl2K9oNoXWd1Bx5isUBBQdg+m0dN
oZCzmdh4elKucCj91wbJl+jP+IhzUmnCUDm+wH6p6dLXYXZ1BgCyuLLNFb+LXAUgCXA7heKNB4Ry
8YEEdcw0+ZYbzTyZ1OHVhhMRLNVWiIVNl89zQGhandS6VFbmFlEJTrePzBYwGqEsDz4CNxcgYG3m
KFHmYCyyJhfljKKahX9AjPqLOh7Ok/qhc2Dw06LmbHPxj0TVKJRkzrvvrbPuQSpF6ts2/RuhVCGc
4EORqffiXNsmvTCq0XtGRTUVK6CM/4smKuZjC7XZ8wAMwnG6kD95balsWnL7uQNgCtWtNaR/Lruo
fWiZsShrw/INO1+OkkxM91S8e5OvmzUrHdTXglp/+GhrsrmWziP9Es4XZIJDFXO9fQFH+42Lwy2O
2cuAxSndnyQ6ICRQF6vquAlix/KQ0L+i2izYKjjQjWL1ZOUI5K09ne7/h9QHNfteUk00UdMPdojk
4Gbm81Oj3rFnbOKhhKdqMHzEwPvj63tF9THfgM0Gj7C94EeqFgKtVXfVq5sSO60imwifn5etid5t
pakOjMRQkLwTlOlRHs+3PwRWQUiRJoshXQFNCj2P65AbOrgwUkCZ2Og0oaDdmNVm+CTvlqvebnqz
pek/3P4kAn14kMG9cHeMUb/V8S6iHcFr+SaAKxkWXTLmRwq9yEXHEU+nzFCt7WG+ToLR2H+uc+C8
OHPB5ldTNza2HonsWQKB0AhP5aVtDXp3oWwDkg9NmwMagGyBUezbDq43ZXljQl/rRBUfuPi6OATQ
rBtewaGJ4o4m43TU+6dYOYvHgrd2YddN5iRzj1vSOEOS+05QKqj8PcwClmmsj6AGJZo+9lhMYedV
WWSa2TKWdwPvr5CD+elpeCSpofFEhF2/tC6Js2zPVdt/jHr7GSXnqoo6sVLBAtGtAhElgZChJqOJ
PKeCBuuKZUrLTWsO1kT1F7tA5eIhMViLWBOvhbxx7phKoM8UZL2F44bRNnqGavNXDMWRKSDYfV4+
4NZwGJxLcDiMk4ioHLVM9QfRrSKPAIfy9dukKLXCEXFKDM7+CodA7BuZ80No7l++ytnol1edcXbv
Nu098SkaPL7m8Ez9wmWMWDvud6Ose3cawmdMMUDi2OmXYHxDo79c5U7eMuJ9Sdw9dyV/ZtOirrH8
a+LjcJPa+/VGUaHPlDb48mHNkP13rLoDGyFJr9Fz/x39bFh/6VxW3yw9rOxXjC+cU8ehE5IyaNxk
JKBAKjiTRHhLkDb3KSb+wpzegwUDgYmlEDqTce7OPfdokeK73xGT9bgcJaxTijv2DaJPRtupOZl6
+pgToiLPHTIeqKB74N9CG7b/e7Q8F51PzcuV4QsIXmAJrnqeyRs0jIpM0jfWDEQu1OAgGElIJSWs
wS+h4cwnw1wJlABrKddfbtMmUK/uu/QYUz6s+tGDtsHm0w+ChalGPyu735D64iAj9imU0xqRQOrQ
aQUcmn0EWVdS8JmBSUV1eDruHD5VZUEYE5LwUOqGRy7PQho/P6Bodu6Wg2PPxjlVnqMWfD//Rmg8
pNibVbcHTHvOMjBmd5Dj6Vg4bEccVfnpsP3bNvJeSUc0uoUBg+X6f3ZJrSPtICaS8Z5APbbBf2ow
szVzb1qobrA5jGLZVD04kZMb6JM1hNAo6usioYcJiX8svOFJzLipFpzzs8Y9Vf0dAcFYENsspUMz
G3bTnNieoV1s86V9DIVFSXCxZtUhkMgEZymqR1aS9MB+MJGhsceg6HhCZYumx942+o2B7hbxDi+n
d6FoA6tTgSVAqZNjHL6lkeQVhrFVFKBOWjDOhhNPIxsP2V5o8w2auRxW4/tma91H9e6JPo3CupnP
tVHjD5SgTGLTQTc06GODgx6En8VdphjbY3m9njqDPqo2FZG6qw5ZxfYvR6QS/P/WyRrIssmDby2U
tPU1LBgN4SQOxZOTWbV6P2no6uJaLdZlvPGU07BPgCjT1lHHTz5neuGzlrEkvwkey/o0uSAHRmj0
iEgJtK4nE51oaj5B1F2E+ucN6tbwJif7boI8K4TBwB8h+aebAZpVOURTTG65Urj0xE7xY1cK7YmM
Y7d+KX6cuAeaXnWygcu1fXRqArResFyWBMrqrMboEbXoJiaZIVBUixtbxALtSmZyZUaGhJoPPk7v
K/qI7u0vDnmbI12CNOEx8wqNi3odMXGPwNrXc068f2dYq4eJh6enNlEHExCqRFxX+AhCKkBcQB/H
Th9GUL+z2c5ZcSxxxyWj1iDGnXr8ha0uye93/NQ8+wiUqKCQ5knwarIL5vsiC5i5Old8sVrkEYtB
DbcQWNNsEcIjyNtgP7OKysVJ259tn1/weZCrGnzfCcfKSyh16hOf/VR7yX/nRdcykR2KMrD/OYXq
VJ96DLkkQ265VU6T4NYOLxqVnd+6LaJV9xiXaO3P7BHub37/FT65lzeWO4DNrknYNhY62Hc2PvCz
OJcM8p3X3qrdyDIP+oiVD22eD8uv1XXMgsEBRTN7wxvZ+z5Zj7yHTfgCJ8721HrBXpScFeXyRhWb
xIq8c+8G/2PBTUwm347DVX3IsNvnDaVZoCOvoWHmveq3cHQ16nb9zKqXDCk+B1Zo+o1H8tKMDjK5
e4ooT7DhMRNtv1GwmvI+Q2z4pLeJIYkIrNDsl/gDM7RVGN8OSzEgCdOm2M4GXEnArtRlW54chy3w
wJVd6JbUydiYRMy44ejQeUWSx1retCrz/7bDd2Yz/ddy4Xkh9z/Vn7A8MvJdHWu9L7a2XPi7Ccu0
0qyMYo/XBFVYheBzEKvsdVesRqFn8ZihDZy1F0tfh8rm+YR6wXnDwLfArD3fnm2jBdLD5/2nA79d
/sodvoU1zxr4qyCMYrQq7KLpkIucJQjQCj3u7H4EJqbZtQ3jO4dqZVe47/6+bOGGorFYAkgF6590
9783XP1D40dF50BX8lLxBGllKNdUsMk7DRSasDUTC3gT7WrDphHJwYvsCDBuxkdpQQwUawMcBqoy
TJ+GYVuuaJ2/zYcm23igjlkc19TIAo5OsJ4SuGui3wRKOrU4i9nsrlQ44DXPIwe1B/VoNsZmOazA
+joSBH34iXXAYFclkFUZE8J1wiT4FZCxRKNcRWKJM68jwa+9eDLZFSoYru7sEv2ESIHf7CQDZSz4
Ip3DwhR7ce831qa8AhVT/uDcI5gIn1+BG/l1E2mmiUSk7BmJFvYKPa7D5L8bua4xjsAHhq98EiRL
gcCI9LVjz+dEa1PDvWBBUS7Q0Xy5dE8WNiydFHj5k0kDk1iYT/KiwEXbyz81ZF00YT4euJj4+IL0
3mSSpdvUHCLwkgmeBnpug/tUCC84cmI8HjlsRxtdc/0qzczZYj8dxcvVVJWNN1q5Z5hPHVQzoIzD
8t3M5eCq9BqBPUCrEHvQgw4d9zfRUd3WgIYYu3SrlBm4aVRkOA6LqeM2o3LsP8RueDXI5OoIEwJx
4ag4TSu7pEiN7FWodiUate05Lulli7UjTNJC/q6/ezE8L78s+ZDZLy6+R9Jv0XkSKE1cUEWPPj6s
a0Fl1IbdLGocOnI4rdEFIDSolJTQ7Yn6Mb/Xcuk83GxYTkufqB72XWAI3cOMiXL47DgOupMD5tVa
Tj3XZzz8mYe5HmsA4DozD4bSjDJvR5uRzGVNRJwGjIhpDA0tYogmvcn2PlGT3pn//AI0R7ZFbFtQ
9pFGMwhh9Byfw4DZVihG2iZJuB7bzx4n3JFrXQd9ZAHABeMkV+PrZ+kZkWcuOIfv9Z0to5qBkaxt
Ky71R7TM5N5YlV3T/Je/n1ROiGRWf/htHxD9/LH66vsoF4bi4mDqOA7jwB2r8HUo+HmQaBr+VGVW
Lv+FGeFidD+QS39JsPJZIi8FZ344P+HpmNI9d7vZkdh4PyhOnW8OVDiTpyKUlN7Id8flTMENCG55
PFbjFmypp8CjsMUuoivJ/IF+Kfjl31RsAl7c3rgGOYkZQ6kfRt4g15i4mhdal+Xyv/Jf2IP5kHW9
SK+9B6kbJ/rzt7+heTGdc+AwzehpfZXO2ARbs7rayxc8K2w1ZEsyb1PzBVM5pAvwHZCytK+xpCLh
O9SF43/Yepbg2IedtoXIxg8a+v000BI84EjjW2QnycoAhfZRIu2Hg72CuTj3CuWp0GFJGLtKtDmX
D4PSafkZdR51Wi/hG8/PDIQJluJo9Trkvpg/JAW++WZEHRxTF8F7gHE1Y/rOafYn1zImD/E1zLmI
nJUF53pWow/QtBWH57xdMyHFl1ntztvIDQUSydzCYvpwkJX1Tgr2qpPA4/iRSq0ni86MB4Nk15od
ZRHqY/otpLKoaEooJeSSQ0Md1EmMsRfvwQib6hnFW+RfL//xKiMs7VffkvmTUyco3KgQxuYN13xZ
Wr/j1GluA3DfdzugQKTo/lNckNMmEFYxqah/wrn+Z23s+5L0VAEO+uCld1j+ZqtHbTMXuUudyA03
MZ5UR10ePmDp3JDX6cTbMei8uZeOX774ZHnI8IrLY4VBqCpL5NZ2bhq1zEeG5AgWXNe9bK0ACLgP
fEQgShnwlBzIGKks6LadKZpO96tIEru3dxI/mgAbLb4xwm15c4BGqk1xz7SpcDhV/oJWHWWRmaCf
EDBs17noHviQRQxB13i/M2MPfkccH9PcJc5SelneDCbRYIsTFmpjw/VYhNxJsZEG/tA7YaV93KLf
subbNNaTvtHxW7rfQTPZvr+CXTZwrMXQDqkVxKasVTH2vpUUKS/CyBcTDB2s4f77VHdDEJK4MyVw
KmDY6Gp20qK7pIVLJy0j8h6uQX9H+XEjdLhU47pHdW3cUHVx1UzqmI4ZVe/xtY5k8BPEBNID4biL
0krxasZ+pHcTfsdB/XAndOnh2XJfIxFA77ol3xwSf/mwvuDWYt5xt/SbijqR4bkC78dnjym6ijq1
DSe6bK+Q2eCPlvhts+FW7n34yFrKdwnqGFle7uVqWhBVXrhVH2w5i9DfCdYxoKjWsf1I4P8VmYij
+uhRTR89OH6ATWlXpZpmsBhxamZu+XEtA30SNkjJ3JUkeNolKPVnCeu/6VV6ppWwcmsZoVrAO6I5
2S+9dXOnuZ2Lo8MCr1SdHwBBlqya/hRyDLNvRBzT3HOTMt8FG05TlrI7Bd8hzGoFQ4y0RUAH48L/
2fctWkUugAXXyeDf8p/dT0Iaya7+lY63BT18pIM6OxZHePg8WPJwpNH0HFkaDoveKaqLLCkamySB
iH4tjWBndLlrXNyhBm7fhXU6wg0jPf+xKJWes/1jzB+cPkp5loNicHnvcSVcVbwJRtOPoN8k0TC1
jYlgqZ1xyP9xSdZ1W8HvbJxKv0XKpalZdRUt8MMhsfYf0YO5ZTmvqNqWBDU2ge0uUV4CFbQcH62K
2WlCg6UaZPRQwvnzdHnpjEwwjz/LQcDQrsSGmSltSH4GrEQVAvjB5F1r5iRkI+Pn6DtdcNsRCvNm
twqYsassNWtryHBsNaZnDaWo67pmxM2YxFADqck0ZoP1LF3Tdq5+1s2HVmAlniudpyz4u4Zwxjq2
RV15Y7YwWFli+8QBH+MtP46plKUQLpSSbKFYYNNJqGEKhmR6/pR7zua2gxdwclhIwH0IJEQzzcf9
+OJyuWPjfhmslWh9159CEvETs1EfBp/gR/GAGUGqjsNsvUT4m5eV2uIphQuEcFsyM8rSk47Cb+GQ
NbMS3WooWulfGQq8dywAT0Y4F3hWYs45BQCPUJPWuV7SQw6Tzr5ELgQi629f+N7I4yYzEhyjx2Jw
W4WQaPvNo4WYv5bcwT09TmagvuUam5i1hpZTPiDK6dXkUw7qVQHvYzcTp8SwvGzwDY/LrYUdNRaq
Mm+EerQpANbM+ItEE39KbMgetosOj7Tb+ZySkZTV0GQeHSWYGbAxHL5jFao7/gl090VpdTb+DqCx
HrN3gj8lg+RGKcLdXJZ0Gwb/aBR+TyGNaTHTtDNU8EDOELVvje7fwfBdaMiMmKQuqlicwkt3n66d
DfjQjNe5JoIGoi4W0//ydtX4TZasrXlSi7KbP+nUc6qZnAWoxz2h9HCN4SbpjynPc5x8txppYWW2
WBttFTbZlE4uAJ46U1zN0AiC975ywENgGEA+zSCRx6u+CT3e9Z5Z8F6DJHi44Ws9+gyWRWEZfgs9
blECPPrVBdumptBoQrcPy+YtC1NiBM1s+dcSa5aqfAfXruiBz3CMr/lzOTKvzr+O9XUPTNvMwUIL
N6WKDH3ee3a1ftqRbeCZEIXY69PaA1rPdhT7Wmgi1QhvnAsYvLYlqLmSC6w8jCXc767/j1RGizIo
EKgI3episUu+ulwyLaX3ljSdqoa5x0T0iL8s3N6+mCIwOs2uvA+JpfBtqC3qeTDNKW1f0xD/T8zA
z/ENr6dhzx2X7zZZ36q2NLXkAROoUOiKQWdIrv4gRnJTkjhAiLKP0+Unenz+ooDqfpBmNUeHIbhx
UuipDmyAHJtknUfwEPSowVsyAdjtnzAEvl4SFeRgz8iy8Bj7KOKNczQQju1GE4yo9amvWRVKBX40
IqO+Hn+uvW7gzGywB+na3jaZtSO+M8bxu80wl/r1w35kwp2L3ZUNWLdY5nYgC6KGNLvOQAo5jEZJ
Uqrg+G06s88WlWXu8Jr6WbFHi0eYmjGEwPrFSZeXIO2a3UKorXhWgSLf6xlcao1SpTcxOwkGwHOz
bq/9k1Xks292PZrFTs9URuy3H6Vhof6RnAL+ZDXYB/+EwymhaFnmvFU4+VxSQdxvEPzKu2hP+oeB
5EZEiPB22WJesxpw9hOavsxv/iM+XNBBs2df66hjlOLkf2jgLlzjmpwK2C9HeQN6VGDvIka7KG+u
/Xtxxyg6A8HXWgbQzYZI5RClw4feeyTPwBrzFAHZaCMGCzCPmLKZ/tdFZ+1oMVNLWF1WPQue4c53
rh20zRs2GvC/5jYZe5d2daAXxWptrhhDJPWL+7FEjO3evECkD8LOfYiGvwV7kWbBRjhtXL8DuzoX
TsxtxeRoceEyLMeiGJeG1YbSf4BZ/rKVD+Zp+Y1+ejeMCpVjT8W9clAJF+esRYKfusr/H+jIM5rx
w5Jrngztx/PCzZ3NF0OOt6oFVHBVzxXhQAfY0pyIt1S/SpdjNj0Mx6ab4jzV0bRFTil3Is/jy3i3
HvwUqjHI6EIKn7+946T7dWLDy/aBuTNo8jpuwZuGskyUfgW+tUsszcrLqY/ppndobn3uIc8dxU+0
0iUmQVf+qOu/EiK19HpqQBxK/biiQ+vxN45NhgCNH4FZjSPrGFgRjzR87/713YNimkBBt6UmswPr
c++ZxGGXWgjneeJKfyyQeGIu+5AfwvsOCiTSzHcpiNovd2b2SD+4qwaAjJiR1s9Kp5dT3Xsubqsu
ZQvADRN8IOm9Qprou+uLyh1c00gAH5kXvE3zfSJzHU4YvH0I8bAjn5f7V9Iyn1VV/eHbmZitOR44
KsiXW6klxkiA3ACBYzcmpVyKlIDRKKcLLFP6L4giQrVjg9QHpIaN6pQ6JNsPAXv9fFbFNT3v89pM
o8llmjnzIC6szoNTvjxAzNDaGu3pVMPpzFPFdqzySYk+lnOwmoZSP8SbwnwHXFOzVzdiSrLt9WxA
hA2awBBPczaxy3v02jDgxB0nKLNcrQhdKfxgobSho3gYT3Uq9AFwBBlOISm39NyK34P21JqHrooS
cD8t1nOqtVtvvgQwFP72ivSzUBbqOjnkG2qzfRO1dYNOwilcUf/MWVPMuIgRz3U9QUDcgmDCuFRp
XfRvvWuwqA8HmFtAUUsazyen4HNWkZHJRXeZzVYXdiIF8RlJsDzA4duUzYEI8vSM+MfD8gjGfzQu
dBCbgZrmPGFrWIFoEOhbtv1MCfuJ0fpWPgghr7OoH0O/HoMZtR6URxFPxIcK28bkyGdGcnyi7ISM
EnhT/6ustlGnOFk9SI9TEwD23NdDG+2QrLZqsPHrIi0ShCKyJe9uGnj5jSFSrV2oAv4//xr87lX3
UocLr4qly0B34cH/4v9QLFZuuw3sCUjKI2pfFYoV86wgyXUL7sZujYLVdkUqn4JwKWrPJ2LOXQM5
ewOTd87FoBaJKeZ5mlRZEYhRBfdVqxZFJ/QF/uFq8qub3NeHt1HOE6TYpmIXVNeHRlVRPvmF7eGM
nZJaS9I9LokONQBnfeYbWANwvAqIoNYbJLsS4L3oWiRXi8PhO6bK9XPRvLU16nffigjsdQyk+h5t
12Gso2EFvp5eyK9ZErLO5pPoo9eYSKroAF7KFakZcv31UpoF6RoBbkPDAoK3/AYWRz8W+xOOxMBa
NBlFeb20xTn+NcleXJ3bwcPhG+3F+nryyXuCSbkPl2hyIEaDLyXoW+ovj3V6+uqhdkSeAgj3eubW
LidfTYNYWwYxL7ddbmLA1+U7sSNwuq3kFFz4zNd+xJKeYLQKcuUAslGzbkDH8ti5WJyKh2kAsZO1
94Pqd85iIfn3rgfJ4hiDhEVsv4OVQ4E0lvrpeBmWi4YVAEuf9+0TU17cCTXkpFjjYnzhO61i6w37
/axTQl1CcDsr5yjnwjIASDwecwZhumYZlSlsjs2AhEpuX2/gzU+9ZwA/x5VQVWvyoZ5ZTjhkSIQr
RLG/OB/UOP5+5zWjRm4n8B+PfhkDymon6sy0gjUsFV2ty6Mmj1NB4AlSOuWIRlebbr7jCAfMh9BS
iZP+4npE8RwRz4oo6oxOPVrhK8bFIMvLC2vOEog3Olctdi/nwpj764UKw7kMQ9htfVSL67C7WAaB
eoQpf9MQ2RaiwInBYatHuxiEOYZk/8G+HXFzUg0BmfSPfAYBXjL4TSYi6LuubOn7UH++Y0LirXKW
VG1fkmRqeO2Mt+5pdleejPEJsiQWQmCqdzer75CUNWlwTzdD2YWVIVP5SF7JFpVvCCscgErIE8a4
XIslRuwcuHXG8NkQKddUlcd9sjGw6wZmwTY7T76BejF2PCDqQWXf7B7tzHZiFtnhACUOkZRB4Rjk
1+itAxZz6l7lY1Ad+6jx0ugiS5PlcOtAtD6UjSJQ5QXX6q0xNAxozjuj0OvpkZa2Emo7S26mMbBh
nAyKRAVYMIRCIcrTbbxBZU0otjWmdKBm9vHAA8H+zlqxM5jzPiuBb1Ovd52twfVdMsZ1+mQbjokM
lQJ4JZEA5JS1FiteCZVp7dA2PUpo6k7GGZzHLUTtsvtxRPaimiQsHBaqeSJPDdZlh0UyK4W7h3L2
912ScpOJSDHJAt6CLYgKJV8ZiS4JRpFtkh6FgWt+DwDpyk0Sp/GG3gVemqqprvNCVaNx4lI30ghd
y3TYYdMXCvXoA1GJUYZu/oRf7tETm24Tf8+6dBPP9FOmcttYGXx8jQ4r44yyvLRsWEI82vhjX8Eb
zxcdaHmLTxRtKFnY4cqInbtgPpL3AxD/mu+5kAGc10HLmbAm03dXuwM656kcIpUFfRSdvuBi6gF2
geRVGvnCPDbD8xh25KyvFjNBsj0M8938rV0Wguk2KKb5urwk+JdSt/NB46zDZnvcTEzHcEXeYSfj
GuHgHAAlHa391lDFBcUex+pVyQ80G4B9yDX2c3gS8NARrMfwe9bbD006Yx72E1228ua3qjVjEnEt
MHPDtQWx/xOZ/hzGj1HEkzsEZ2T0Vo4cO+s6SEPOTrr8RoMrhyK5d5ISkV9tlgMGMGBIyi2e93H4
/Rqyr715hhvnVrCWCPTLa5ORg6bpfuL2/DcGr5e+/ezRJiNMCdBzZ16U/0hN7/b5pDJqfjVZh1tp
bTAo3DjT6fbLJZtfmzlzl4ALmmUNgfNWgkSMUx4ZrBIHIeUgk7Up98NbKmqI+RReiozB8mfscwTj
8gPKHViIpOssrIKqPUWuywmY3susC+JESOmU3uJPQhlqdcxzQXz7fmNT+t23zleuLxoPzZdv5us5
eG59UJMaEjRvPj0UyJDFQgDUn5ryL1+ZqCNtE2Lr90CG845HkiQq4oflWMEBIDkTUOyw0oEXEine
Qg6V3ZdVSKMxiHODDlT4WhCrol7PPOt4K4fs64A5N46vuM8IqPb1LXyCgsEeLtxpN6YcSsbMCTYk
CoqrDo+6Rjo7UKWOjBDwOpJn0PBxX+hdhbmSrbDkhaV7wFTAfR9sMce0AOyIqOSbYsXk4bA0eoqW
sHqIPZtgqMmLDNGNO9ZxPQ1TLu9kavV8sI1W/1KLRNZ9F/8Wv4GKsopmw0xS80wexoFvgvKfVwyI
S0Q5XmlJLp007mWGAS8zbqrtFnihRJEwmrJEZ8SqLwMKGp7xzAG5Ibc+ZsVxJyGxjGfq2xkwN2VZ
c6/qQ5t/637Rhjo9P2Q81pHdF15rklF5l3N03N7wGphI0vTGc/BQwznVOTzngNG/PQJxFc5zSnVh
Fc2yTHShiowC9ztRs1OSw6gBxCrNt2hKrnpB+q5/7olfBY8gonnSlCS7O88FD39urlMyHIQqtF5c
PxUnrSbYM0QUjlw2/4WJoeNB/yRV1O/gniF6/Y1JMqZMna6VwFF4vfbX4ysdg08TttzuhopA2SG7
8gd5FLQKUROhNwF4tfBFlA8ep9HysDMovDbdrYNG9Rf+hHgWvtBQAxqWJYlq/BrRm/q7rX+5nrrz
ecpnERNeZDm2ai7nKo+xqU5W+hFC/yrjgxCAiuFBbuVrR/tmQADg+9V/THQf6b3moF6oNE+PBBrz
W+5PcQqhhd+X7Ceszcf2lBXklLzdRpaXL+Q7v9lb0G5iU8f+r+/0Rr4AFreHo7VUBFciVFBUGIGi
E0VIlw/SXEosb/iypggkLd5imUb0pz/0eRysePYnsgJgFh94Xpo78B9ycZ+0O4OVGMkmgXxUpq8P
F17TjPDfvkc52YUO8cIFh2yydjDfw4Ve2noTOOafWRkCjVfffJj2FQYVGKTb7cmZEvlZSYNvkt66
WpYxGJNRqKR18pIc3MiDXAP9Sm81MJPsppngBQT+tK7IVXQMcnG20fr6r3V+/xgACQffb5dgjdaA
SohnKzd4owh87RqWb2OpFGQxTzEFMMaNg9mok7n3eNByLI3FOl5wJp3Eq85KcvZ2937qcm0vA8e7
+tKqHdCDG8Ws+MihYL0+LnnQ5rYhos0HNQ/nuc/M/2B3JRO5lTwmt8H6/pXsOHe6bI9VMW3yMOsI
N6DuguY0NwKGTrF9jGJpROjyQTom9mvrvyZR5PpVgKelpGG8vHaoWUfp8V12KyC1PCg6ODWd6gET
xnZz55nQuMi9My0o4HUCsV5F0Stj5n2L4hc6N/2a1o7V5LKk48PelC4zzbf8xDBxZbjibOO7HJbL
zuAOqxY3MmwfyrD6RNm9lDjPriM3wWABEBihFuR8SmTy4VK6jMH23mZjCjUbSeAuWoHudTME+Yqi
jBxE+c5T6xk6Y1vxuGh3hgvjUWbzE9uQ52lrTgw9Hw2pNbQ29Ez0KE2BpWGwItd5PxKVYHhAU19t
Sx4d+GZ8kV2rYDyvSA86ulTCziMcBjDArMEFMMnwNtdaLYIwv8IB9H3Pf7giJog6yUtuEvVvZ1XC
aUwiWdOjR9nByI2pgIq2HDRoQEYe+ikxcOZHZIwQXa/sQpDSqLRWJnLNtLcszojlaY42DQ5mP+6e
gH9jPawpyD71LcS/YxaddBczoMKD2IQ9arZQSAMJ8OlldTebGmhwBgLEbxfnNchdXIV6D2mW052h
sIA5wG/H/M+glGNRE1C4qxfU6RdTok3PuOZIGj/6dOh0cIoMUWeDXG3030DgRywuySk8YAWMYT1D
MwXk2osent3hsXRDs+7wHNIHTFJfXhHJRAdeFMG8l6/LASP+ribMpekO0CRB3tWRAwA8y2Nhugw/
mBhpeaeORHzaQQmk63VG0tHOzziUeK5GGtetBIqLCBeo7zVD+NUZsIY2WoJUqxqCn3z9KrniI1Qg
g19HeMwiTEs6sd7YJaGlQde3zSxqhSuWl8dU7N30VnKfCNyqFJSZuXHar1bd4RWFgA1vYHiQgK+J
R0thCisU6VA/Rw7r0HjgB9gTeN5ON5/1wYvjP9FM4XBzQcO/swEathzR4kuOIYyPuql1RtRUChbg
4CYRG/MCA6+jVkdFGXFTWBVzmmZKKYU0c9G6cufpVHJbGMwiJdtHRaY60415z8odTA6AvfrI/++9
7cpNTd1iDgsgpLT9YyLMdzh9znh0nyGHIx1Lr/mGL0oQuKdBBZOh4NisY6N2F/KeWfp0wIkYCdHf
RKFB3VrZVc3ERT6ISwCcUrh16M8NQsxoEsSJ22MoMwUrRlnFWdp4/sxLEoocTfFCSkM00nzzZc9F
AeKB9ChKEa4DajLm7AWR3oj9IX8iVe7ig9Lsz2rMYVfWrFr0QeHDr5JzRu+X90YHO3ibbj0vIBy2
5+6fKGV8w/kTYad03HArzhOcCMnzJYikz6eyEjNbke400aSiTe/irnsmin8SzO2UnvOv9J6qmJxY
4UiQw2bkAAwr6QoIlBDkYGm+FUUzljMZrhLya5xzvyOLVbnDVtsn32XG70n5rFIU+zOfNVy05sDc
5ztfg1P1bvwy6cZtv2U1U6lOfzsu800rE6GEeplADp5/T7MkLl9kQ4zhZMEnyGOptNHIabtMApbE
FRiF7EkRUgjTTfV7jyYuTxGPyYfuVXfjhepztwd5ETi62GapJWXKf4CHhyi3hFCI7yhz2eLsMzjq
eJ+ow6AeP5tP7HemMgshSoevYMw5XyGZRrNQh4RT838uVHQjzrl1Q+H8rRj4G5MhD7zElmEld7Se
8uUY/Pb0WYi1loFQaps6L1RO98U+IwMIOu0nlbApvr6xdrYqPyW/paIl9N4H/ghXkHZVPxJLpWRe
DMa78OLk5kIsBYaCAhwE1jNxZs4CBEk29vuhfChv9azApEtUHhVs9L63T06xZvkT/jLksqcslZQ9
9qyCn8JV3Smv/U7wTr0sHmF4WyM3j1gQNGqI/qum6x7Uu0B2XkEfavljHoYNyH/fiXoLkQHpIEXX
B7TLlu8FIaBbptmVtN0Ff+nUb6dHZJW/636QRC5Ki3WuoDGrOnYnlFJFGHE8/uX1Drj1glWlZxDO
gQyhwpgHBgbCRUWISXjBBXGzJKItLKryuY9n3U/4lUMkNi4j/FkNyavNp0chZxFP35X82yG6rDgB
gHKaeADFnLs44wBwWD56R+cJO8MYWIuql8Lg6i3vJOlV+iCBkxAYixwFpNYsdrQwh62iYbH4sRpe
oGRzZQOje2BjsGkbVCM0mSc44JsxJsvDO5yF0NPOy4jUuvRUtsQDhgqOAYsRK6uWgeC1v4PJQC27
sR7o+H1FKI6Uk0sK7LC6v+Xj1z80rWKg3CeoNVOy1xQQcMh8eJyDJKSeYo3UtDWZJBnFbYJFdEpT
MLaq3Jyu5ylx+LjrIGY8VjsbavuOuL3I32czvh8TTP57HwRtsESp2aPfp3CWFg9fCIQyr/bI1t4I
30e2DIGm24Svk26T9/yskpkGkoJvj9yL0PJ/ifUnV1NP+Zr3V38RE0ErkCWAdAPOM6ix9D37u2y1
nHW9aVBTsjZv475ijA+lexRA57iIfRCTrWQMDi00Mek8DUonXfmPzOR+QvwVq+ffbwev+8LLAnVV
xVHJfOjXL5wz1gjgwYNvM0qX21KyR34SnkETbtUWaQJohVccT5FiGYFqN6SA7K4BKdPv0rsMVekZ
EKn8YPXVfkuI2YQFdmJ6J0Mna6g6OfjfaLZpCdOQwhDmSdeJdrj6yAB/sDlXFgFuDSdK+FGhHIPy
yPr91R+B8sojgvqSdEqKrmdCdFyEt2caJM3gI8tIZm7c1dbpAYpcZ7X2nneAeiw5XUXfGXMilQnA
2kWjZxJ9JgvnZeI7eVRRHtilizv9D6okT+sJ2N+vJQoTEajaiIbYhOtKdleZlZt3tfePCKF7w/vO
5MqOCSGymBZk2k9jvUXD55zzxZQSJL6ZdYMPkYp+9n4CcLKurdauGmB1uDyenearvD2MZ+s9XJdf
2PcNQajTipZJ7/9OkM+qYz9A7Jzlxevv0CFEH4swaLAxaHEqZQ4Y6yr19cKRUt4WDIEXMie3nLsS
w856OyDRKYiB8ZakToMt6oG40hgTUeTtnDzO6CmuAQoDCIGBZ+Hl8M3PBpsk6eYpeE2sFcWXMCJr
Dfxjpl7wX25yFxudDEON74MjyqxsRFdGAiDdRFJLqH8TpSHCmZC/y29JezsRbirmHueao1huwWIN
QIM+hzBY6+/Xna6EveJORLLG3BYpTYGakvnch3hDBXYA/L+/4ihDJnyGPIBew4dkYBhk5O00zAHS
TSYN/I6pubGZa4M1cJSKGKuiHbC+7cdQwGLK/z0zhc34KrYEfkLzaPYnFy9nLoYnvx7omMzpS1OG
CzW/jtXESpUq1/ii0Td4xhHV79mUwXHKuW4kEZxzEXrXqYG6WY3Hyfspc2wRFbcK3I8sznWCUOme
7+zHWngUAVUsHbmk1TO/IqgwZpMhcqLd1WHY3E05aRN5+/pISNtYWOFgC99HKk57TCapjyVAj1++
QhtLqlOf93zudyGl0sNJTdT9I8rF38J3vRNMseVr/Ov8OgWNNZk+1MOEA4Zcv2+OkTINymh2VSKM
q5YvbUUfeDH5jUoWmhy8X/tbmQxUlPT72cXdnVXxh/5sZr51yJNmP/3DVPB2J6dtTf3H3LEBBAIy
/5Sk/1POsu6LIlGuX9Es8wcxWwKY6NDxML0Xbl4RvWp8wfFjUz4qpFETfB4vfAKsi2zTgPyUzUqb
FvtA/DDM+XC1RUeWnqD+Dylvy7pKVytjnymwDtp0cP9vHnskpX0c0b71J+bKmQWSKUIdt1+nLYpw
6ULT73tiLz/uJzPpzZ4ZqEzu1JYnehFlzQwyvgeSyNwoH0wNG7b1y2MVbZDxSWq+n2ZkPtRs3MBd
MBhDYzfzXUpd/GrLaIHGSlJXV7VN/Cad5bpJWBNW2wMcw2yUG55R3rETBIIP8ekZ6VmahjO7DN9m
j7jY2cKGEeTnMPEL7gEvJAUtaN4gGhQwl2s1AtnAXTZO5Dr+jkDTjSkXsC14EkmgWgGN0YGog8lH
KewEWwhZKp0eq/rk++iIEHBXMzBeNc44RKW84MZRvFp5kcR0xcWwnyHCXlpnXsr+GqS81zU5xzol
q2qXCECOSK6JqUbgzOps2UayW6zRnGq4VmZMQA6agvjztzzqB7yLHWYRPxxMnWUxek8JouE0uc0k
Irma+EuwpaOg6k1wWa1HpEX8yWVFTsBvdf0qfL+RoUzKyE4nAuTL0yROcoCoZfvQT2y1w8gESQqO
Zcr2isijpu5DvjqTfuvjC2Neft+20DRLVnppIDt33WQ4tPXxTjSNGATDV+/aqZI9XEnBp3Z21uge
lh94+m1hqltVuWFLx9/d3ghFMiZwfvbSJj6kFNGuniCFhaxUuFyNHt/pHzw2/XcYq0N2JKBvg6A+
iRopcsMDgdM0ngCPriyF9OgylPlDD8xBngc+pGq+qXTXPaQcS6UJFqf3T3bXMp7SNvVTIYjmhti9
7IzJHGL4yXnTJ80ZYD2858Wiu9Gq96HihSp8B4GLV+DOEWX1Nm3z5ldqJS/YsE/VyGxCKK+3IwBf
5mVVAphHMmRn5gIn8yt0nLDW4Psq1DLmRl8vT5kyB2wE9pk34ayniB1stZPYJS5WD7PLtXCAoJXg
e7JYuR+Nc5xXMyekPVMUHnsnp/HtM4LBfjJYI68lEjWNitX0jEBhFcHvUh7dDvXnBwoWqwmLqjaw
wZhTVlkHFizhNzjVmnDnPCvcrXyfvaHAggNw2zSOQX1DaBL6Q5hHb7yicRFqWYpatTrGL/QxDSvu
TglG1a8X25F8cLRL5EBoeVhGWe6uA6MVLShJGNOEQoH1CyGxf2Un2DSCoH/yLmF9s6Afa0Cwxzs2
6m8f5VaVucLR1VtX6JANBew1A+iePLYCJymUNVvWMmlLMnWvzMOwZRDG1HPFENPz+ClkqKxjJzsG
i/6ZBqb+UNwoiEKrs2yz+d1cwhPfuFjvccMun1lW7JHh+0BOaNIP739a1zdw5ok24qVKrFL9WSKU
kCRsuRmrh2hoJFipJG4lWNaUaJtl4rsbp1oIR8iyLaPBBe/LnO55U9wX0Qb28fw8e8zLCrAVFRf7
6iH/iAbzSop4h9FdPleET3PCEuh8CVMJL47Z2xO2uFqIpNmBM+EySiDFnreBu+7BuaxjNwcD9VYu
DHbuS5I8oKS7odpJCVHtYfy0+CzmudHqC37UloIcY44CsCuo9z2mcLfy+Kwt9sFGVS/2LB44KM6A
+srP+obNTsPK3YLFFRvfkLLktDLJ8TPJA6SuuNprJfLd2bEFlZFCAQxSK5206FR1nOprL8Vkt0eO
qJ6ZFxhzgV637a5Y+WZ2W/WViBVxRzFtq+0V5bkDfv+wIIJiIE4L/a93I1hyJk75BrunGzxb5iDS
7jmAgszPQWWDV46plK64SyFfNBBMysqwfPyRhZr1TjQamfWi5rJ8kN2h9xG6mYr7/Kb95CXyA3zC
hQoYTeuJYQwCVU/NBmeS43sDmpe/japYyzQnd8tdCsRgmf/IvkddQ5P6jfBZFLklrkavNIOw0Zwo
k7ouKzrc/NXs7OYqvna02VB5sBS966VJ5cwUuG6bxnsgDkFCJHa9ciqyzfQ9VLCBN7jD6fghOl0D
ZmKUCFyYssp+m176J6xYGFIJHNAJdhdyXe9pZs6XoTpN0MravvxX0yQms4Q3XHMKVC0mZ0I791Nc
Hn4prO7EgAmmdErsYH8OuPQjc8wh4xml7HSzuCahfkc6DrVdP2f30Pq+OIxI9bfZrT4FqFgzv0Lg
P74Wrr1ydTqRQv7vJlaBZ3SVhmHOO77D97Gm6FsjaMOjW5Vs3nBEpF9Vma7H7oPGfCXRopS8yayf
yY6dR4h24xLzrtPdnsP7tlNyOOpwc5rraEEkMrLw9TmmiUJtvNzRTh2yjVLaSgxBWtGKccpj8Vz8
oFcARsgPFFsTPHt7tYkRhcOMXS4cm4OZDh42wrrIFsUMoyugFmzKMyxmPxncnurD9JOtvuN51rJD
buferOOO6cZ4vh2GvTtOaSSdTOZ2d9YgVKTDIxFaG2jFzWTtfmVG9Da3wXe7mMUk4Mnv/QfInKNY
23UQPfX99GuN6Sb0g2jzt9VIbR/J98ordjncK6wu+Edx3kMRCUkRo3U10IJlePa6uuy2mgUwCFzR
fLq+7WQfo62K4EZmGsW8W1Fkkx+FW8BBmsE5b97WwWTMd6edEWIq9zGH7f09ScxEJJ6uhrcaXHEx
wbkDED6v208F75ff/5jYopjnMlTzYer/ZXPNvu5S40ds8LgSIYRkgvNbACkzEDUDiApz0Me3/sD+
nes6G4r0mT378mAW+peLagS6wb+quTH0n7lCy6Q76IBFUvvymGi0YfBYg9Bp5pLqVozBnkLT9Ok2
vwO13UwxZUxaSkqhIOnARzWa2VFq1uFbLa2ntbK79duwDz7Q/Yvc6fXEuLxzmnLICiYeGCpxk6ln
fHaA5bLTXPE3RN5dHIdHXimYx2OeE3Mr3HaPmddnlk2JOmjj4VX/EJcescpKQte63/qSCHrPF74s
sLlihmHpDtNdTdTNyRI09QGM25VUeyX+enxKZifxoFz5xINQw47cGKhzmJZWj6IG5Lbsx31KwDBr
9ZqvPfTQ7HRZbpd/u+zcGslWWMXmsF+w7AcBmH8myNFY12P0bu4/X9tjh8f1R/SlYIy86C/xPzb/
U6e/lE/lOqACrGhaagbJXXWcPkIWyQcXZd/R66T02AR6CDqInUPdGlvme39W+z0woX0/3KDgmt6m
OZ2H0CJmrdu4xBJAEX/V5OTP2lkIYWQ/KDG9L/rzFysBmu4dmSRM3CUfLMFqXTPpi9cbink9QmWa
Tt4z6z6+Ek7+QmpVAF1IGu2MK2XAJ4yNrVTeY92zFK1aDkh+fbBiRQXb8HELH3IBvIHM3ruuT5V8
TUK/Z1Uq4z7GeDyiBirGQvPAAy9Is2W1ISdzVxhvN2J0Z/XZg4mYRYLESat/9zHwwd96goVTlLNJ
OZU3Cv9BLRQOHhx6RbcgxeG1j6A2Ha5NmzsbypNnHjm2tn1Pf4+yvOZKjTZlTKo86OUoJSUuUK8i
BDvFaU8IZwLf1dKBxVk7S+chTBXtF8oMmajgbFBPSa2GjArd9VKZCwbK/TqXszbpbVd/wOd7O3jT
ml1rHyn06hV+bCpyeteolH3/CTkCV611eLzubcrrqz88v65KyQ627WDyBoJLRgiSqJ+wGtgPtTdP
oVueZVzgh527u7IyQ0YT2s2NS7KDbU26vvIVaGnFeHSeVSnllnZ+esMQnxzgqKZYcgDOE4Ch6i6B
6h5Qzu0Nt56INPHnpXyqv/lJO55sH3eGRXuixVvisOcd1Nz16dMXE2li5A7qx22DhylDZhtAHakf
yES0UVVc1fFYpsDVZPpESNZiNQI8g/4uBZvXukf3CPAL8XCN95K7mxCGy5bZkbU92sGnXy4eTwmg
FmP+Duid0h0Zgz9Y0GNXs6Ddgky/qhzrnJ93ztkKQS6++oX0p628a7O3ydxIDmPoNBDDQAx0LkiW
GIqhmnpPGnORPiPVo2B+l7Q+zKTOyhshlWO9U//aDYK0MByfCDC+e64Mt4eZdNNRey4Nc7/7DNed
vNGM4PGhoSdgSLCrve5baOTk0xQYe3Lht1Subn84sbcfVmUOcCHjt2sK9mFdmH2yePJed3ASIwW2
QZ/4406TyiTM2C47lFJhSb8zeaF6UNfprHV4KSYWnUybue/ct5LGPMuF8SsR7GgaCqcsVJFWM4+k
Dbbm6KmHZ+Y8YheDZvdohW3WmPkFV1Gu1M5AzSpQ0VpXUVI4XQpv7enEBwAY2QixfqhdlFIE5yCv
sO2updf1/300aeOJ4cKKkdDV9/rRbaImoOJwKuH/R4/Nrj5LzELkAAtjcLSt1SwO7xwmifNopecF
fkaM5yB3fpQwX4RGZnsvQG3o5LPivybylfzIzf+o7myPS9V7ClTk5H6sHAQ/f+i0h1bC8X9QxHO3
XLnkRtl6Yqk0rorvT6qYDRL1xDW3kE8mSmis9g4lUsyiEImaEEfOP1MKB023dKjvjKSOUQh/DPSh
HknMP7A1PCWtxAxByu3+6ppn/Bo+wQrAJP+wYRc6P7WjrZnKUk/NzsR7Nt7atDk4lQRSgSngtAaC
6zrBIDywUZmNSR5qNpXw7cUzeWdze9C7U9i4JDsf+bJVoKwkAq29+6RYSZHKPd3yO665q+8sYyu2
iZeaZMcDm6r28AO731UJwHusYW4voYh2dYzFXlLmoaibKubHMySImffbOJbEbAgpXU/FlfY6OMe5
390hdX/cZV6wPIrFKUNtIO+kKMJGz/4oz1u7WC8Nu5nEMnuBsTxxajY+Ph8b6wnQVv4Ea+/zvf72
bfaCpPYFxrEgH7Ulm+xGlMk7KtK1xG5lugHFXFN0F4Ds1KIBiGLPQBsq/bl/xfmYvIeumM2zn86e
GrcPqNdSoUK+2tHIFuP+qfCSxgGnBP7rWVkOPM1H3vIX9Tk9Vn141UN1CXU3LTiInetZP7PhQds+
uv2bZuu4hJ1VMrXJZCJlNhKw6+8GElLRp0QSyzQxYeV5N1oKdq15IKTQDURZNTQ1leo0St44+0+J
53pbJ/RoBM2qnIZc3Dxc1y0uR+mtLtoU0GoYa+anoswdjqKXo9+wgsreSIjnIoFi1b9zb4hvI2z3
oYOCjxENu+dwdjXhFx3Yrz4nQYEXjnkvSSypv/DBem8+zdgzvDBkFIXUTqBkr5JNA8PAVygPcsCP
XkCDPQv5RLahs4gCASmtL0TirBjVozDDGJ4dkuNfbEdGrCDqVQRMjsh95q2GEiudZnrYcGH+vEKO
CwsReFcjE9XwDivR6gaGdRTujm8H4Mv1wVu+cZ/h8kWhsSM5w407DdTqp+1Ht0Lhe+Qg8WYhE5Vy
f23PZZlm1YHXC9FiFi/uI2qKJQYF/cxtdPPpM3JoZVwETDI6ZBSny1ZNdmMGkKRKYyJ0FDrTxg+Y
pA7SCzym8zIjFr3SowEb6yuq6PkCCMbDQ/m2twak2WEdqwmfx114utQdEJN7hPkek+sX8CA9PtZC
w+YGLKI/oywYt6ugy6zewhvWNkUZCWOCPsL95vcm70y5jXT9Mo7dtOQjJ2UrcaTj3sMh85nBQuUh
y4Rx671OtXd5OiiMAevJALEZooTJhNo3Qc4kX6SE6A9DFGfOHjDyM4aEIsLHiJbxbA8zhgl6IEBv
VXPH62WlVmarXtWJ2w6J8q6kqtCNCPrswxmr0AdbFa0sfLejidpXDvhNn1gMjDq69sOm5cebqv+M
akKFI0zWSEvnGaNpwXTh6eZx1x5kykMxEgRaY/ezEnJas2Rcdl1i85W1n3c7gnQ6LPUzat0pwLrI
WhGP4AHnqcTPnU6wYuSHR3SQMTmkfHTsLCG7YmJuGsNF3KjMbf+r+Rovvy5a2dRUv4KFzMjB1Z31
wYSO2lF9jzhITrH8vRIs3mFdOxy7vXCkOSpTIVQyMj2J4ZEjbGMbXfhj8q/xFibzC7DX612PfmKF
VOn1IzdEVv2vCLMSHBx50Uo4KWWYu89LuEDEso/LUnB8mNrG7IpEgrp+83hLJ7+y5W6FaRpzQimi
/3fQyKKYHsCIjxgAAthiJWjqAginAeMjt+M1AV94tkZJlsdN7H+/G3jBQu2nue3rtzMPiwUd3PuI
xtIDnKCNzeNQ6EcvxdGbsuzcOOytkl2hPLZsJIOaQqzEhSzH6OqNs4BcI7KUyBIY75vlG5oXF3kJ
XvgCwxOdoLazGpKNI9JvJOKnfeK9nsIX6yEqF6aFOacACScABCMaHL6zeNZJJ/JAgvM6Sb9hB5ij
6W+CRCrUbFtwceUcV47sOIDBw7V05gb+9BpV5DHtykrsqlj7UGqjJjILfpnloF1i0YqfNQjxO9nT
BfckPKFNZdBBK0aQ1kxpSxqdnn19Quoelg8gCACxNMNo8h3gr3iPSgKUFiBVMjHtcJbAI5xebsol
rMeV7n3M1qgkUWV9YAux/5a1QvHAVAZYMFDdA0F3fQKvpiKD+osIdJBUo3dQ2xmrG+PVeL77tZcv
lmOIZEoT7og7ce8eretLegJ8L1+mCFImovdpCegwMm0pBUgdjKtLrjFu3G6cs8uQlU60mtFIHR+W
apcep4G015PqyOnzl3AeH6MtsyOICSi3X7RhlHaFdhPOsx/+FpcecJFbQLHGAY3OynV+WxTZbTU9
U69r+XvTAejtmt+60tb5BKCbzkjbgES+/FNk3AfeSmkURgu+lmOANUSqMyEz4AOv3kQltXLYE2qk
WBX1Z0DjqGDQMHh5u6VDnvw6IfIVtV8iOYu+DML5Kdj2aBEEowcKyNV40K7QJfXnrVR5S0PK3eDi
nVG0tA9SE3xOZCZlfkkF2VrmUp0mfWQS3m5x7O9KkTHC9RP1SXdoo4cYvSLGe9TMgixAclhojvSO
DYtJgKjrSwsEEcdKumLbGCw8hwYpLpXH4OCo/NOMXbtzOBtygbAqKAGz23th1yBAoUdapGwsCeM5
JZtUS2MztmM6Z6O8IlnOW4nCg/XIvliRqpNT60mX5Ob2AtN4B2UpQ9gBpeV5GymltBxKFDRhXS5Z
zzVabBuil49caY6FEIiRquXXSFpFYXTXmuU8KDIbxNL32BbBBNINAoLWZVswxTkoTTetIWNoIBkN
jL4lYVnO6OXfotjMK/XL8jM+vgLL/f7UaYlpwNQCxEMVo6AmHPsga2cDVMp6jQFZKSUgdMd3+JG6
okaf7kcsyM50vHmtzq7Vb4N+oP3e9ivTyckjNT0g7wdN9TCzesQPcuNJDbltKwhZxJ79si2gQGWl
goaAKcU4JyegY23YilgBx4DqSiOvti3odb5rix+Rvguauo4MBBTWNY6OK83vUN+pwGYk1j9hVd/d
Z6wA5ZhJHpAjf+2rW7R8MFtkuQ9Vc1g/HqwKfP2D4Y6PgA8gt5HpEn7tc7OXS53RAfdmUAd5YbaM
lcmToEnWg45Ur+5ZiVPgkZAiS9TJ96KiflJLMLMNTy/fjVlHVwpQk0RuMHyLyatYIZZINAqzMff/
Kd0kRDUuvq6TqM+/H/jpxe4BIQAvRsSzf0aiMuyJMluGBLuinFeMSmTTTWALJpk7O7cd7vHyos70
zbK44+uGAN1w9nsT4DWftnHIBlyo1A2Sh4SzzPwEUk67fiDT+eNozS7ZCTsBJrciFhqmArhfnLEM
Co8t2/lNUblXHtPF/w2YoDB3Y8Lrc2mHMKDQO5JhbWjP1Tl4euk/EYdxcRwThFswhawgNuA9GMYn
USMkAGIkJ2FyCblPAcaFCr/Ns9LYEBoaebuyQD42Shj0CW1L0cKr40X4YdZYOnABoKT+tW27WmA/
gaIOKhLMJgCURqrZGzYDD5tZrqqPXL4Q+WdMcCXHtkqEQ/gUltnrxZDNxYTlrF9BHUJdqSMFfaQB
bonD0gZrDquKkPSzavVElkH6eVfNCGj3gRVW8EAd5xyeX7Ke+TVt9SXnDs9APfnJjUWcazS/sTzB
EixPjMzMUJqeAPYiuJqKHKAtzJmMNVJeulh2Hh/ul9wneDUItdBEzyKErJglKunf18tAO2ZADTft
zQfuLD4v9FQUFdNC06R849FVuPaGmWsW67m9bpjxxHRwt1m5S4H8EoiuQrZrP+ugWSurS/AImmf9
fAKQqlliG0iTzXSRNlKIWNvzVoagNU7jyr3jlTSl5vwR4sD6wZWnV5zatEN8uRbzzA4tzJSWDN4T
vNWE/buRITFjqnfQXVCnNuvoCtJbM1EQceFBv913hjGOsY/Skrx2QhAuTKGSPB8sN486QXlxFSil
DnGPPLFbFoonE0OuPgwOrg7qXhSfF8V/6F6epv0SrNs9g4FCOqDcS74ioIMmARyYgjxXWNp5Xx3d
50w7IU0vBq7QBJZ0l9xpxsXgoUslq9Ry5zU5WZyVM5kMgv+pmvqEtyxp98k40GEVlFzK6Qmw13GG
tznBKXFFQdiV7sOe19pRaYRIRgv502SIY3LPNhMizTkVttEwjb9VaffCfCYlLbJp37rwWQC+Wjk1
D/jjGnV806WfhsLwRO3lDcok7gL1073KK66t+d78sN8dVUe51u0xqIZlp9VXg3UV05gMRYdIjAk3
UfYN3hdbdkAzJyB45iOgN9kCUKkrAdPJciCBIvJ5teFtHrBuLyFuLv2XMzzduQi4i89AiIWXQeDq
spSqvg4btuclpNaHiBlpV11MqFMp6LTWsVeLa2/mEf2LUHUQ7Kgz33Rp95cNgCqIr8/eiBf2Aghp
G6B3kBlRztbvv4gDCl+yreGZ7NK05Vn2uCsb15+TpsXNouKSO3JPl1QcrmARnFySPBf2MaL0xkVs
4yi8LtJZNrY5K1mizRpENj6SCwYX5r/LBWFfWGAnBSF8XtZUD/LXWoLkVS9gllA8lHgB8JGBRAQP
ZN87dzDuskEGJ8usgDOCf+qJI0QFJ7TZs/S0QYUVYvvx85mBQpx5l5KO9Mmqxwoo548Q+sjIhVmY
W+pWVqGWv6nrEmYvEUSTes+liArD070WD4P1EOnq07AJ/mG+6/Rn2WBJRlpLUlhmOmtRPFyC85Ww
iXFISXvUCHYrsRdUGEiIAxvjHcb0wGXwKKetIndP8IoqaT5wRfAe4sFpQAayiW3wAdCFY0rqi+xV
FrnfusGDjDKqiPPgNK5DEkIGQgxSajsYudoEa9jWjcPzxe/E5LWOIIeL2eolWyoUwVFox5IrsoSa
gHihRumCPfe/1Qom4a3AYKhMuVjgZTbQf7L8NnA+79mGsRMEq6XL2yxlX0i7zEwgYeMlFTRcgAhy
a269WPh78VhxTgEBD6boVhZ14wSuEX48mbmDMP+s0PZqLYtNx/HVuHcsWc3b3Csry1GvWHaw8e9H
h5ayjPQretuzjet2l7fMqH7O/qDpExW4lsgd1VfH502O28m1pHlb/FMZj1VXz8QPTUkq2CpVGmYG
NziDbLDFseCnqA36sVUC0W32vxsCOQvm4somxTnCOtsMf3/fXUnizJOEtFqLMfBaIj63MQg4h1is
4oU+bsPtettuOvoKKGj8EElaDSWjP/elyv2ePqAOlyoeKoiPK+3pyRR9/w47DnXKWLF49RCm4BP1
UwnF5cHokkpViSxlZQ0lEm/U9QSGOTWHj+SDgdjy311dAW+C10P0YLu/keSzR590kqileMiwnVNW
pXoa69S1d7Ziotpk64sWW7D20y4U3GecwuXxpOMV5mCQEkqZZ5K+8WLkFjaQZ0n3ERwZYORkBERx
GWAXHXgu3pxOgM8uhGKJY6ncBrFBR150+kBBzSDG/DtOYORgOCM8Pk+HeNjCPRuBaMbfSDofZUyb
ju4elWgNuckxmzG+vqlUZq+FWzH3emNJBQm/TpRnVBrWjepEcJu15lPZ6qXNiCkG9GCV7ANoFPqo
LisyhOc54jhVpS4OimnkVUL/qxZaFN0/eGObz2ZJiYBZvmXVHgXyV5rnQiM4EzDvkaFNUaI1htmx
W4PmhBm+MlKAshP39HXHnEje4YVBNsxj9XCGDqnAwLn9YmsaNatktsZtnQ+xWjUWtMyt6QuNWeCq
JZsy7G89Bgn3faIkrxu4rtJMk2wRtrTGL8ulJFViCXjnumtmvWVnkf8Qf44tDmzUyjpopo6V7rbh
+2E6rcS97kjpUOLB3eR6xY6WlCL38+7Qp8CnL0ab17RDORg2Z8g36m683iWCbUG7tXnVAI++AwSZ
j9YDsD5dv+OHbmhhz5ui1d30umlD7dOHq7HghQw1fAoGnielwINCGX0bYvz74W3NPYfg4aheNFhP
KA0ZKCp5RKT6dCZjGMafO2OKKhvL2IFlEVkkT0h8rY4hDUY11xVC3m/fCqRbgynsFu0jLhNuEYgY
xfinOlDHhsu66V9u/ppWxZB7OntIqbdvw0hAslTY33Cdf6o8T1aKLpssPQUcb0uZmtaKWKfs78qH
Oo+nF7oHUyCIPVe1C4eRB/yBNkb4Jtv6/jbi10FVk7r60fkfl35v83GbTIWPZOcs1y9Q43orGlZh
9ObcS7M2CEF74JJgiUJESwqEYtFZUczWtILn+4GZvgmxPAnjLgUPNTUB+UmgpsA8TMpWuDAAufCT
C+gCxRU/B0rfOT8StkkWes84ZMBRP2X5uQiCF6RIMp2aRR5W+GElJos4st+2So7B62/uwfks65D8
55P8q6lWjQKlrOddHfb/bg7haebOvGgotCPLuy/cXyVN64pehXbhvYjdxaDzvZX2D/9XY1lQGJyE
KZfJlV1W6yuvD6J1PWyV9o2P822C7zhdZkz20Csumauwa/1rCHeusjEvGfLXy2sqBPWxVk/K8iHp
KM2PINkOPKEiEuaHoetzcVxPYEUi9jSY7CGswhoIznQ0AcaiiTN/mjUAEgxor24GJUKQ32FoOe1a
b7g1z8kGx2TNqX6Xz45m3oWgxExMnmDW2JH979PyZOMOWd1edHtr+tkKXsKQbYJSiPve/Xfu/LGZ
F0bjUY1afVAFx6TXTINaurxEM9qoxZMOg+VS5Bt7j206I7zACmRmzpA+/HVrYFxs1DmQnQAQLt29
ftGYoHVpGILDeJdCxc9XV7sjbYc/5SFbSE31BzUTSh3PWh6komIe1a1lnsSF7csEMdBoLdIv7wqv
W2k1zRptI8cgUjebzJ2qo69Ll5OL6svowBikCaOvW7B9GkRWf30wEN4NTUkD/GjABc23ex/xLwrT
i0wr3XTgTUxuY+2vRTyCWXZ2gixQS2IducJE2NMtDRQn/OKhceKb27QCKP19fDcXvggJOFEN8XKn
XA8L77Z8AJNV2R5NCcQYa+i3ZhC1DGZr5KQeqF+ll8D11ntojaSvD7P74ux2FMBrrVfdxFkAmOBz
00CtprH1R1hqdpmpiR5YgAAz43G1MOQ0vb2TPMaRz8NdmWHPHCMpWz4/N27m6Zy2GBIgbHYmRUV3
0TC5EN1COyuh426WCFsXGmmXsHF6s7reEwRF0uouNygyP/GJxTuKXXIxdJY94mfzjnnGQm/PCblY
/X25aLaUwp0BUZjWMx/fLNUpxBuUUurEzVDdRkCKCTvHgLSnnf093XAlZDXvK3M1yNz2J1R9G4fb
x0hkEnusHcnaLgxry2wIE93+/NgaZMEOUYptUJDs0mkqPSIn9AxqKxi0oLvaDEsSWkfijcEvo6XQ
xMfHeoqhwQzD2pkFTtaiy+ATnDk5efL9vgH3mqvuNibqkeXEZ1QnHK7YWs2A8WvfXBSRjKnEhuK7
mC4w7sGRx9d396VlEmAgb/L1lREwA+Zpp/oHinQKKzAqqzLWbun4kDoWRa1A9EyeBzDeGFpbIwGx
DDg6ni+hYv/yR/BmX7yR1RCQJsTOjkK+ylAfk5GpSZtTzpeoNq3dNRL8hjM1XHJ6+yzyKi/87zX6
DADL9LiFtsN5oQyLxFte79S4rFN7/DslVuXTMTMqG/1Dudmi8j8Y0Ct1fImoW4QXoeyp/TOl6D0n
c1QmVKYpC2TPqQEtyG5wFr9zWO9va4GXAezAgfdmtwycYMIaynFKQWlPbat1DrJ+OBeUVFGaZ4/B
RGz5q87CogjDa374AjtzbK8IyqVgTK2PxZAPHfxmyXfOJfRCkhl+9Yq7MqnNQhT7+cLl0ThDtwRM
n7s/qtlBPNvM4TYU+XRtPYkw/H6b//60yMNwpapNHnJs2Ak03pjs9t+u4q6HoW9Rk4uHh1MFnRvU
0NLbH6eAkxk1HiqmdHzlXRnoxuXt4Ny9CY8O5TsxydGla8bwBpU6QyMfY/agDA8GqxtZ5iOIOpGJ
1fHljqGAZdp3L1amflfjxLGWe+QSADVrDzmjR4L6W30HjZfBS47bHh6BpClEoXrN6fL3RLbDeiGT
TgcdYWSIdJfWrHo6UJMP6uoystZffhOkHY1RLCwQQJ70TJeBnIkXjCwhBY4DMtdKDY7bdH1sVj4P
OpqKJAYG5wBk+qUDL5TlsIag+MmrFIiraRr18UrUxjlJCJijV9sUeReR8xByk8k2IqmIXaq2OZHw
ymT/sD0oIKxSUE2953JT9LNxEHom9aXn+yBzY6FwcJkwEiIx/621ASNL6ZP5lXl6Pk7o4vvh1w2J
SdvIVMqQt3nme7TpdkCHfbWyXakx96Rblbh2U4/hq2vgGr3UxdpzfXmAJykDbfXl/O1YfGPpO2ES
CRszi+cMnzl+uORBBRHSCoKAz4vIU9ekRVrnmWgOCIQruZycbLkQMrgvmSTb+rNtPPalwPDIs4iH
xZqOZGOwfNMVZkbK5UCJaZqt5oo80zoMT+KN0A7laRrvxM3/4z7nHYIC2OifK1CXTpRJhY8xWz9V
NjmkE0muf7NssDtV5TjpYxh/UgJuKBkt/XSNArd+Kp7MtDDWQjTbP/0SFuDMdGRowhzhNRa4iftO
y9mEzNYL/NoB3y1yUK90tIm0THeNX+UuGTSBjMQbRdK4+tdyGADZPfL8EGKXBGo2+ZHIWs7sHZfK
2g/sTjW7zjdImMvmBwclhyq8m+wZEArrbZjJoNKfxI6arwMXrghrrsIokFC8H/HpnMY24XPMwIcJ
Pl63HATEKDVWo3EDymuDGh6AKa3ExEdsKNE7JMrF71J064Q/gwxKmwYhYhtQMI94tT5myceNjQBP
OPxV3fOSIJKge0+f6PwGPGR9NFXoSEpqB9tWSNh1kV70aXFR4/nW9ZOWnngyzk7rD4qG0tJ7DNft
h5tj7IF5mQ6juras7V2fzWvyrNmuh3CZy3uPdWaI9vKMJF1Mmz0aytYI0mosbrkeYIsC+ZmeDJ3z
urvpbq4tHSLsTELKbofEI2CeiThIdc6ggTi/XJFWWJLwIsGYKht7j4uMPrxaao7RshSIAJzCPrpN
mdFtYEKfMBqEYuwPNyVLCyrVN3OzkeRC7tXGIVPHJfUuCSzmQ80NStqhq4bh88C2hjOMAul2Qhtm
KqMFyLHiG9wDU/PLA4xLxWHd5b+0i+u4dNqnGVCa46EwbV/hDC7bj3/sXThNmjzaGHsIL6hki3Nt
TXTF7sIVBoOeGQzF6r7RWwCS/1mUPJPiHgWwYI6eA/++sig9fB4JJiOtFnihXLNxS6BgxFfnmOvl
+PkwF+8YeqmNfl0CZ9Qd6eUjMVAs4ruGOxlumSXqQ3xpXlZuGVFmFCxkLOn4k0fqtrqgAq5HB3PV
QDGNkvg2qwAwTRf+YbGyb1d2gYqu1sHzoa84WjkhpmyVd6lB285o9EJ1A29UJzk7xZYBb/+AsIlR
x5TRfgAeh+1+c9i/1UdBKV7e39AHiY3/qHjLoUBEENilxPeT33d2scVGrItvTpWT26FVXzyF5/x3
sYIELJxP84ma4nKVD63K5brBwuHMJ2H5ktPIndYYQ7C/4jl1AaEUyBwmiRNj7pX2KTe9iAHh+rA5
EeoeKCLRYRSTBqKCfWXaVbYwKUDwx40zoklNZ1kfteQd7fBVRTYZnD/brN/iwy0KLxg98pfXxtPC
2k62mI+lIX0wnpU5jHwpi0IOrLkuT3Br3+Cq90eAaRfCQ31Y0CdPMEVjqKeYuKzEHSogObbLlt6c
yvhyVYoc7RBKPmAFqA1wQ6pS7wywglxoTc4gQs4r1OvC0vlS61goBlN8nwWHb1ZXxvuwcbhrqMNa
dCA7JKw3s5MZxEoxEQzbvV9Z9rUh1GkErmXRu3Yu9phtAEqdEO73y45FiKyO1v4MCKpG2otWIcnD
8rmk3yVYZ10j5z31JDE9gC51odXwEuuySTIgtH7ESPEAyJcsDlxPtIhlhCBP/oOKUpsZb0e7CX5i
0hxdH+8+L4nalS9nNBofSjzswAPqf0/Ms7mlJ5gTDp1s6QNEerv1d1cnXGLdhZq45heMaPpp9Zqo
1pAp9BmPDp3JzXyMzH130OVZvYWhSgE+/Fdn95fYaC4qHPAgY5LjIKYQrywT6P72cfvm6xM3pSsA
vTFjyGGxXhdT4pVyrXpCvoL6yXm0RfjGsaCkEBMMusgm9cOCAX0EaRM118TTKLw1qM4COPDGh7F8
cdD3WXsD+Qe9ILKmyuB7+llMnKUhfh0xx6qo3RoFLTSpu23t9VyQSX14DthH4mDNGhaXUlVhr3WA
vISldd3Stpxtv9Bo0ZzOIa03uXfV95v4QN5ss2+ulh2Igrc9cNIkqm/OU1GD1eQIzyq9BWLqfjXC
Yav5o4tocIf0Ts7W5EdYrkPH5YVsYSoEXTMBuzf3pzuYTLI2YvpHzbxbp3Npe1MCOol1I57DPbUf
OpCw4qfcdvdbkqnmfkc/MLukuLYKJxoba++cm+q/EGjHNGFAk1/gnp3KckOJw+izLjko1nmLVRac
GEM9jlgi9MtPtJuhWc6Pkch83DEq7u2LNWxdBTioqPRY4fqjvx/ZmnqkSF9UlkbFxkxRVyjC4DbA
BvS1sKi0lHpycAKnJrA+T7USVpalKxAP1ScqD3DXTK5bPGWkUUuk+V9KLDf38xPIgiiPip/BgMhT
QBV3YlcbQhknpluRE94JqYtGCq0JVcq5+FXMxm/V+0IMoITmMi2EZeJ+mLbA5YnCoBm3cUIPv89T
a/tJ91kQZb7jLM6HFvkp3bqYkaKp+RD28fXEDMECt7WUmX4aqRbHZAsHUuCFpBv6XTEn8EoTDQns
C4T1MLQwcCTrLWW9aauubepAUSraCD3hKAkXlqqdh3LchdrAe6vhZQpuKnvxFxy63J58XagPHUnE
F4vbdpdypAYRaZSbT31/jBHY/TiMe8cwL7eoTK8DN+H/Y4EIGmzMpHRBojd8IufQ9ztAmNsnvkC5
poWfmX3rlQwTZdgYwoimK2f+7H8V68B1WzVzPGup5WP1Eaes0zcybTy20nUmX0GA/ZA4gfTuimUg
TCzWnNXcGko5HseBGR2Rauv20Qkc0yPoX6Xz4sxczdat+mUA6ZolEv2aeaIz1PXI1GlIH3k/RqXR
q4OPBV2v3ckM2bcfoz4Sv5f55LX+3OzoGfOAmArvOB18sgydSOFQAZEYFJD1iCfIt0bHf+DCOEFS
M1uWaMuSSJQC6j2hlnej3UpaOegm+s8q0pD6tBZsTLBpafHSC2mJMP35u8CsK+o7XkzOOvmjtt/E
C5A9I/Jvft8UionOBPSRsbTuHK34ycbucs7mNGi8kZ6HqT/6JCLyYjdPZ9PgEJVdHwkXJghqyvup
HwquYEuC6BiKhyZFPPrvn+T8+xqC/Z100tjLAlH7D5b0vRfQ8Uw5cBxFGPyrqby9P4EE4R34eXyd
4/cBcIy1tQSvlAXVH1E4Ii4SREZKO0TKz1qb1UUecGLveXu3L2cp1fbd+boXhWBH8r4jMFQvdfIm
Jcg+aU4PBAdJpk8+1QUgnOjTuigVCDuVOPTxhovSR2hU/mADbhCR5vYtubEBYZ2Lb5FqSfViri0/
25Omy1MbT/IN/gG76DglHEUi2RexVngGf4q/mq2QdMJQGL8AXYRXu/1dUwdkBQsRDjxFH9Sr+/Xc
cPHBnWuXwPy2kyssElXBP2yCW7Rs+H5Nw5JbrWkZUvc//n6LWI4NYVRAl4IKP0i2ZwfJLYUd+oe/
s2e8rkeEnO2aSEJI61bhex9U3aKe/vNjMQX8c3r+cQcsmsOqCsE0DTdKUcULiCnJ3hvLdvQYp/4k
RadfEXec0OC5uM7iocy4/JJIfbVxcK328ZrCAgqs/dsuOf/6nC4MDKMgoUFYo0cGKtUkIwKzsD0J
YIJJbZqQKzxlzLSmOmffL9D/WfWr/31SxxsDscUTqCQHRtRr3w3pH+GmPej0/zphnt+31t+81rwv
jCBaJFvgxYOUImUkAqbVpu8VhV/N2+qXQVFiaXDuNuLyQ1ua8dVtd7kUPxfARegfaUMJZ1xXCAmA
bsWAn3/V7MKCjYLRqC+K49ghdFVrrcOfcfFTtXFOHXRrGLAvo7Uup57A2TzsM7E/qUBQsrezXE5i
xtQCwZt25ra7CpeQGz9aO/7l7gTvTJeow43Eg/iKX/bzUQqwYxP+FyxPHUCyshI5Nrvw7Ur0fh78
BOjn/smpd6+EdkP0KoFZhB14yJBsA02Tnznsa+nTvjztjAgFX4kbrjNF89RoGIy1QPKCsyt8EqwL
qAdz9vEIZ1OIPV1+Xk68VeM1yk5EoYHTbmKbioSi9fGEZEDSZwOr2f0JCb2pODuySSdaVNPNsC35
8Lw85mqpF9p+QYH4sJ4sqpYUKD5qSptNuK+wlz/yay6bfDDemy8T36rjfT9lADF8H4ut/Gv4nJ05
0JkRj1sLCX1DtoDLZbS0wKPTIfLVRAtdhAoS6YhyAziiSO3SWs/5I0m5cjKT7F0VXNNrL4Hqh3zh
sYeuQg994HOtuloFHDQxIuAPW7Yv2K180BoYuqM1QW9nBUExDs7bCZy03rAwDM6DRM1PvaJ/Av4c
8rXwq/1SSvQZ3VkMQRjdpKWzIZlbAK2klGLLLT8eoGZFb7P7/VGF0cwnrMrKXOsa0HA0tA2d5bfj
gUw0LLJbmZOTzahAP5CoXTP8Y0l3hvK2/saY+SP1Tz+xA1lHGvmutIPcSl1NDpPInGSWeyyXryBj
qF+JvYab30z2qsC12KhevkzirUL3+AJXJxXwxEIQYw7mVxNeaXHnn+Y679BR6Ch+Pjp60LQzxqh+
YKWUIOPSJ3nhRCLRgOcUYbX6opunTqTBcpAviNQAX+6UKPnMqZbNq4dVFlDrcTjbKjVjcqHR/vvO
efxJhVs5m2BpawaYj+dL7cHoyURVbRMtDw4kUYX74N/PTS7wfR/SUzcgFT57EdhphsLxqQhdCmpD
EmDf6mxENa/FtNZ59T/ot0GOCoR0F3f+KfQviPvAl/zJtYKDao1WHb6HvrYiu4n1+vOuWtEbmfAa
lXtIKmpMzweky/cW8coASeva8qNYw8hs7KCeAY7fw2YvpQ3Vo/yXqHwX5MW8qu9w70k7W50JW/7i
yC8/qn6o7RwSROLksilyfr0q7dsfgH6Q9Drx+2g+03dNnxCSCfuQzZkDRVQ6e29nq67gVt7p4P0Q
Ec//t9yzexPKadR6MhWjM9+7LhZppD6mmzhiUrxPNjxgx9HGM4HQV2Rqugn2osN90aTSW3MQkA1M
cBLR6JDBmYN2zIuG74tmug6CUKjcR3Yokh5+jfZ6dy+jbftCQTa82Bf4kr49HnbXcTKF+FEf13YX
dQCAz6xfUsLAgB/QNLiyl3TfFcU375V5rlSE9LjGwVpwquRNnGo+qmfWg0XgHgKfbRehHw0OcQHX
6yEwLdvImGsISsxqzi2pP32x1qMwAnpADvj3Y+xNdomFCq7ev4OzR4XZBp/7hOSTGxaeAjGnrWg8
54X0Z8IHcpMqyDzFBH4pcCx1fO5ivjMIGAmo9sbvPJpIcT1P2et1rW3O55zBq/TnFkZvGoKNN7z7
vdNSYx/LNJs6OkHoGMHSnCq+axOt4mK8JqpY+6WfcHhpaaJEEKfMXvDYaCXJC8Jy2FBqS74qIWWi
1tDKB0ZRvTBWIMn57uXWfuiQHSLDRYSpYYF/TH6Gm2dyJX+ggcY6tsUlmvsrDGQNSxdTrvB7+tGw
XTr2TBrh2Sf8CN/j487gq4kAFbcXDcWmmhW1GFiKfYTzHQutjCb74pbXQbW6jhrX493dR5ko9zyA
tpuOHtl+kOlW+yG2C/nXgrfHbWNVzsfdJhf2mvKyvweNRdIHc7D3cYb+HdBetPtijWUS5j6wTcO/
KSmXRiXtzgpai2g6fqMidbltHtpj7Z9Sq5mN6KMOvLDp3KkTlm2Xzjyk8iCEyGyXB6O/jcHlrDiE
tvZQ8KxFHOIsvVOuoTe7aF4qNIJY+/puOsnDEqGdwy7uaV6BNSqGPBuJON9LjH//eGlPWLtNV3CH
LsSuZ//JfmQaIiu41CSY1G4Tc+rC4Nvys2GsnAG2LUFRY0xemhdavKktY8Lsvz9KMXAk6Z6/L0m9
yDs/mh5GeeCwSQA5lVN0mVICKDgJxNi/nMmnwhesXJ7CqdtcDBjAq7flS888gcM6iDYXrxhSigpC
nZyW4YeTJ8eHAeTS/OEjPDk3gVMSu4u4xYMAJ1+JXWRwWln8jM5EL7k3fL/9RCPjj6cc5kKenIBq
oVIKZLT+9JmCc6seHfuNZacDOdwhjz+iCrxn7TSWEppgd8Ji5yM3SKYHrw1fecQ4SZiC75OZou6T
tEmKbkvtdqLTp4xeNvCIgKBzTbUdSFet42tblyduy7mKDDbfmc0vI+gC3pNMnReWmCl9URDL832o
QWthtgeeEkR0Wk4HqUkwrZ7J1NkaY61w+By5aZQG/DwAa1ZIX6Rs/woCPRxvwLnKGQwGetPDm04h
YL8xsWhkC6/+ZBSbXnNFLccif3DDBxiEIauLUkMM7Vt6xwqIls0OoLcp5256yLnf5UINW92esbNe
Ymv/gn/1V+U5YOhuIm9T4Rry9cLUxsCi+PX/tMrHmLyRsFMs76mp4C3FVsNdVjCNYeFbHIsxkAdk
5UuKS0HWjowt/FvcYozFO3qZO/CsZCLhXhvFTDSrYRV7cXhmT3vCJRi0PjumxqVKAOn1T0OO3JkE
0hVHbU+JdNHYCdc0j31YBXRJPjj5/XnBthGBdw0O/8EGHdzU5WOEC598pZr4rUCHcIai4+q4Gz+g
nC8C0cQ//kfhQMjpJhuZOXarDj+FRWymL86iljEo83TGERdpbc2gMOZ8O2jDT2S9+R9Z7/IDFxDX
sQG5cNKvojQw8piPenHAqghlRXD7pNhBSrWH2UEcHFOzMgea57O3CW5Zk2wp9skv388GJOcpRQcn
wp2dAml9bWHlKRKwTbDlmicRYgQgEHp1XpNoMxQzNX645sWcrmkv+97hSvcCMOvVQGdIlwIPVmOC
cSLytOzCZpdHU5icIhbaqtII9K0C9wPLzVDGzVA4BTdoeJXGMD7+luyIQRB7kUC9nXaQiT7yb5fa
/2+a3GkrEaHxwtS7MI0IP7So7hjpKrvwOg00MiK192yBXSRoPCWrUhI4vv5ZnzyPaP4tWVrRB7rE
d0KvKyBaorbMkbFXxBQwJTuMLxjUnMXDbmRGE6E/e9E2bT8hbvMMRAV6O7jG3ZV0rcjcR2A6ezse
8c0TD4XLmh66Lfqcg4yRNIBrQ+L77vRFtq9MCHm11KxR0me9//pBzUQxl/EasADOYzfeHypyNbU5
ZWaM5DjwHG3+3XDNN4Fik6fwYKqDkPpcHT3wGy68QMZNW4FgKDBVXyfN87DYPT5Ds20kFHs5Hf8A
h2KI8cLywqYUDeTpLS2Ka9CbIcTESpVser0upp0AhWo2s/w+FXOTSsd9engcfaEvOS6ok4r7fxGV
xbcL31I42iKsgtbfpBSCptcCs3WqZ1fTfGW1FQoaZhuG2SOyAo//8e4FasVUg+B173tVXLu9Z4IQ
mYl27+GZ12uNATdldW8fNQMiWk60LKxJu64BW9Ehh1fQC2xGn+J/u8aqOmFtQnWYZEtHWerx2sK4
vtgEaVuAtBkd4TdJnafki+qKOKjOXc5VhdJ5htJh76IsJdOhRVvpg7pVf179ACGus5F85GR6MgcZ
VUNk215Wcz3bxwI2vAa3RObyHaO65jMUSIwDXws8LFskDEfN3Bt1BwsK3HvWXt4DogH6fpMuolFP
zpfT40tOrkONr0kQ3ZWAFYxqMO8KNAqx58Sd+K73lUDVGQU4a1oVw96tUbDnoTIusjH0RKqjPNfm
I+xnkRDYkWkmszYgFTn2Jb+cuLSJ8ryvLn9OwO2EukhMH5d6w+Kmhkn5q5G3kWXsj5QiCcVWA6Re
7W/+4tSPFb6iXFC9tPakPb8niNSECHfY0JJNj1P5O558wmJkQVJ17QTOyck3XTtSm5MH+SSPBwmI
amI4JmAqy4OZHAGjxnLh1/gd1XIae144THjxZbicxALeISxgQhDDYzK4RUD8z74SCoH9YgY+Q9Hl
uii6hmZ11ZSlF7JxS4ef7SlOEr5Gb7uU3yhtskVlqKUiLWvR1wt4Kme/leGn8Iuxsj93AiV/mBow
qSTOvCJdn/mPmWYRBS2+A2ieXWvOg7d0+gPjbT/wjVoIBCn7/1Xbbt+ULMz9lB31pdViP6twwgSx
CvJt3R80XSdDrGH5YAMT1bJZ7/ul3j3hnR6e1jQzHLetEAdZgn7dIW1HaBe74QEjbQRhqYJpjXdr
KQ7BqsxIRyLUyOXz+WIEJW8zbqPhCXyVvFLSRTwK1vwauoLtM6Wr2tUCz4eRu+m39doYvdonIjA7
auEqJtwItI17EhGcFSJv4heEwT1Z/W+195tvPCV5gMK+b3aE04zU/lpHYDKZO/70sfCrtExuU6i+
Il1EOhtlrWBxdR69pEWhbRtxpi5Xf04fY+L4uKfyeMkqdwP+2GDQ4OBUPrEo2gOilKE4P7hcIt0h
fEtu43kS7tjAaOnJ/yNdhGe4QQOjys4L/kP0VR2gEUs76a9GFwUvSy4QClznbFFc46j8Jn6Q1DYa
stAp5ninSyU0c3s0+18PkH9bhR0SNxlqFv7tKFGvlk9I1xVcOCpLXH313ardz6uICeqQVOP8h7HA
Nkeg+rFd3ITJmt6/7Le6F/Elj+XCWewfGi6sdeGNbF0Aqvywvq3eyH2bgxem87LHbOer1OpHlP4c
xVe5YAhoCONTxS+r5IYhSPCDK7N/cZGeVNccfNi6jUvyCEYIEbrJAZ+r8mFEn4jRwhjiL9G8+4AL
0m/zJ2sa/xHTDqGjq1o3Cs2/lgYp0mSrbFCzsiosOSyoB19qpLjo41HWfru9Ek7hhHSNiBkN2LHs
wkyf+RC60zWMk4Yoms5f1CQmCY8XDSIeNVmi1PNQq+tnkBTZwkdUlnzUhypauPsZ2EKZ76V66M90
kiQmSz00M2FQsdXtS3IPVp79vialBO0/sjegx3xBKVZspx/OmboqrXcNDdZspJLsfe5gyusD1tVQ
GkPpuQGqQDPTujTUHHuJAoKU7qtc+F4ZkwL0Hj8+LrrVUwDQhwyQBo8l1X/mYatVg30Mycao9CIh
FmRDF4pzbPGaQkNCZ3YaqsoiyTbp/SJkRiJ2DDbjd/uDFarMAlHTC2apE0JbcC8e4AN25CDm/4Vo
nSanxd1aTABfBcFVN6umlq3rbZduuZbDthXwLARQiZTCUVwnK1IeEfLEYcUWYy8eVL+m15RNEEjS
SIFk6qs+F326QUOCiBe9QZOTwhOZlqKkXG4v8wXwGFzSTqLVmb4u43/iws1gPV7j3VSi+YW/i1Ax
lg801fpyLvW7aIGa7IQkajsZTrxIHzAfs9Xwtfstzsu+qIQ3YTtBkyJ1UrQrjW/z+i0oSFUPVmGd
07IttrwuKbSWu5lFBt8e5emQCFoq4DD2EIGbxIEA2SrFWbszbNfacAEjM7JRculnIIqz+6NF+zz4
zYy6cB4Ln2+HSQIKtmcRZrJHBebKqw2sJZFUKrXLT4mIHPQrB4fE3jpMG+I5NNayAwYXnxkvJcJ8
WQA6FMHJy3a04/9FgYKKfa2jpbg49ulOxb6knzsWyvmJmghU/FDrCZU4TW10mDT8sZKwJXGK9euH
uV29zSI/jqz2BYnYDsKwomc+RlQjYEZgvu69KEterIbKNMjeyDf2br/wFX99pD/8xsXkEYADYFMI
hwEi/7CKuSHMQAyoadnCGdEOxJVM63yPLn6bioWrDApbc2fyBOnvMG4GXZUWVgRLiQwnmgUJCJ/S
ActAoYKox/SpJXksMzetg2dX0v32RnQ7zZ65s+2Ctfh0uznk4GRt5Q1NRbMgHjulKSCqcx1jqhuT
akeWo+/jRbnke8+xdfosnX7cEPaC1O6VoeY1Oiw1xDU+BovIE1If5AMf/nQOQ/4dUNXTlqBkRd7V
sAk6xfHiF7YNUQ3TL93HTjws2P0k6BRgRLnNiJ5LK/OKIIhn3mQWgT5hqu9woF6TwgyZR2ch+FWI
dRc2KQkHMyWaN4EU8i/ha4OSbefn9ffdsKGGCxYkQIK49dZtlm2GXyAqV4fnQVQqUH3eys029uRf
TgZ2hrxdeJuDpD/EQPjZZl0IrniJKlje7ZsAKmm/4ATnpccCjA7xmknkFu9aD9iNwccuQLPVqK+e
qT/91BLNtci6289TWP1jj0OiU9OrOxE7AE6j+TtQGy2PtGxu8YkDFyBlLKY47bPYzVzTokeX/KLB
U0OXEkuWNqGqlCM6LJg1ljSb6QjM2tpNEcONDN5WpKiemBwgpadYgn4TUgr5TpYeoUFrz9Alkd6l
iKFeQao5QowSipwxcCn9b8L4/2laq+3kzRaYNlcnmxluoUmx8yQvr8jgm3mHUu0ilRbrdiTH3sA5
rcKu3DU7F0/DNQgwPm0uKhqe7i/GdtPXyBkuX5eYYBirWQ+WSIrQizzqkxXipQDE4MZBhZgjLp+P
gGyOw0EXv6847bag5tzFQN2HWEmQMBA8T213o4Cpt3s7y7pqSW0hjjYzLJAZNrUjfdVORNlZOboF
MLu6Rjh/6Yguo/SjSEboJizA+2wDpgjCM/xiQBOM6FqT4n3gHTEGqJgBHGXnxe+B8AWnip3ktreH
F6fkZFagr1h7xQMS9Aw/+yCxRKGkrxc2jpoLO6yUIQW12akf8k3v7x9M1E1xXkFIlalBsIFZfBQ+
MNtekc1PLGB7GCqeny7ROR9E63+YfE8bWMezuvq3TOzDPQEdmVNjFJaJCfWihXPumHqrjWSuEy4O
7acdQG5PzO65ZOeKdQkJcBTX61/HVwPGdWC0olBdcqXOu+2cvnsg4AKDtEOHYO90qP3PEF0RdhCI
AHHJbL5llEWxycm43uAqrSna3McfTiu+JbG3WPmbGSndJkjl2JfC6+8+LBMgAl3w2wsxTjFhGMTr
yxB4sEbtOzVB0cepuQG1BU3zFFQW+eiswxEaqFmjji5NX8G2fWp73sMC17dpDut1eSJ3MQeIiBwY
CvOiJ837rVz/GaDKhxrJcca/wFUzb3mOknMGfWnLcW/kNiqr9X3cbt8pbEbkwbschcXjZ6s2Jqy6
h9Rk9iFi2i2e4xCTWrIUhl6/ZiLUhAZnBAurApN44iPB+e+/pWsIqmzD1DY5lK4lWPGMRMBIrM3C
V2YsjvT5EsyrHw1U5gjMe1U5DpUVpVjbWQLqhFF0bP451IvOYZQfqaDGjqeYcVPghTmc9UigM4Dy
0x7hrS/WKYwiw02b9Xo9gNiIZQYIZOHJ6QW8qVI7h3+kg6ndIuB46UsS2kpv8znlFpEvsjhtGIXb
Sl07DGmn+AwQFPw9HTNwIawkK3r98Y2/6XX5vt81U44SoCp0Khp9zA3o7QgVmRT9VIG9Q1IKk9ZW
IBLyx6XufYaoMUmimHqa1QdKwgdcVhcfkN/lcWdCg0qkjZhxsqpQFg+Pq7ZkaD5pLfP+7o+VoeQU
RqzjWXvVMMf9JLqSbu3gixtQmQ0CMzoiRkOGg47R0/xKBOjCVgFt3/2L2FGcf50GL7QkuewQWLAQ
SQ5D4blQOaJFFuCUz1LY7frOfVcCqjseNtWgx2/kzmid8oDSoHUj00FXH4Ztv29dDAPYqFrl/2q5
7rAfZkKw7Us+RZlH8k2LYeia4xiNxKnfpgfit5nvJYxFJ2xXvOa6o5YMW8gmnUTo7xIPel2s7hNi
r5kKIa5oJ3zpHQYb+WpXKYWOzxJ5GM9jz2V5Nce45y+uBS1GA7iRcvn3lJ0B+OovSAYwTcqhVFpk
YjupR/dzJXeoNtXUH8pf+1d0qKXcQlWpb1034tesbaw3rE+u2m8cHelRVjF0q/I6gVE6hErbkegN
PSUM/BQL3Fet2bPP09cAAb12+dFKHZ32A/msXsQfJ+Ly35izHfOmxENQS9ERIW6erwkwH/vnATBb
wo4jxVHuw59gU/GZ3snIkMDIFo8zy0gHYOp5exNqMwwyqrnT8AdfaPsqYXjZElPfI4y+TZqckMqW
BqwtyMaDHE3k/t1+Ex+TD+CWOoaqHKFM2cPNOaAYrrtiHYHHx0MPIBILumTBL+5S2Sv7LsdDp3Sl
/at/X+XL/ISzebxm6oQFDctFVJjBysM+6NLjPpqhWheIH09vdBKwgzQQIXLgt3LJkqUyqiLz3uwX
i1JUdQ7Byf3wiMNInmGoe+hGNTjEFZTfNdWbajd9sP0WDJBeVnFdxPtkRTJdKuyhGP5tf6TfnhOS
eqyT77IvjCdYDlnTfqmgDBrkB3UqL1eR0hAuCiCl3E3Zjb2I6pwSpGewh4lbfvnwHG49n+/tqBGa
tzX5B+fsYC9QKs3/q8dcazTO224kbA02DRewHTaItma00DzasglGAj3ROrRqBiGUkxkgDLu6acNo
UWEJNYYiOWU51Gn1MkSIu098ONW5BFbj5StK5QrEpJwVUozD5KD+6GWKq4894lMy4NfWSrlShokP
ZJgccAZFlTChOZRLjOvmq6Gm3sMn6aK6t/b254dDVmrFwiFNM8N5r80xHxsUJq99uW8Ye4Pi79hl
ZGRti4ZdELXVCfC7CpPjyEqdBr2mEe8ZeLY8vVe9kZ95yDE4XitNf+D8+TWwHJOzUug8e93iThmx
UoD63WQjQuB3ySy9uhQuoFwaVYQO6avjlSRaLz+bHfxlUnmyj7GVIq6vGsA30jba+F+hGL8FU6w4
MLRzrubiSY+GXnGWNwORDalr0MBcU++Pa80wInVTXGMGCW08r8vI8wfXTUApAOdUwQY792+h/Sk9
qSBCzQvMl5qmcuzVU64HcQ87kcCbFg+Vib0RMEuWhBfDIpjiAWR7cb/vb8so5CSt8QzUUDDmPjcI
uNnljbb2C4HPLC6zp0Eu1CLzG+dy6VtGi5tTJ9IAKOlxOwdjjdf5aQ0h7nNqjauHj/Pea3PuWQjU
FeFpfg9jT7oNGPiCAawlvKOHYVaOXGjjAX49na5o1ku4kxhRLfdG89+8UGdE7k35uMtVev2+qq7v
47DAs4y9zy/sp2dGCArnX77y/b9BlyX/HzWiXF5wYhmjHVtaXONrwNdRaxmaWK4ovY48GtrJUHQo
UGUVV2frayFX2vH8atMTn+Tx3AEjTaYZ72sgQEEvBw6/yhPrTQuA3jIsO6w2rKhiDW1R5rZhxDj/
8ozfl8okBE2zYoECrZCCp4qUi36lcZOGAMRCuAjCPAIihQznE4b5akpRHwgshchX9vNsd1mz+CBc
PcpJpHni2XZnxDObif/o1IUQfgyvHLva6GgTLlCdmlSlMVwOGzc8HZYD6/hH2Gz4iPMfNKXoj4e+
WR3ds66n6VVgUDrp9GR40uhSdt2o+Z+elOBoSXgHu+DrIg8ISwar5PTqj5TE0taOiUmC9Ky+Z50M
tN679W9azdw7R54lSRysaYf14EqpSx4N9Sj837UoAiI+HK+MagPICI6G8zUi/AnwhTCtv2BqZKTw
jI1cvV116b4kP0MIvo9ZPTyw001+n/HK492XgjWiXxkSblETiAWAZL7kLbKteQu496PNN1/qnO8I
ox/YvotxPZYULpIFNdvDZVlHfiYQ77Zyrct7KYfg+eJ5c/iDkxoGrxOd1c/eVlMaT8z9yy1zSC3f
jZBMrpJPvSZaDV74FvsFURgJXotUGNadjp259xHFDTs8JMyD4YhwXcCMBM/DjM6qmSc8ZdqmLHjc
MLIWCNbkcTH5/zZZkXFSkPrR4WISxNhxqNnfGy7baxAGTHyGjTqipTNQYQ3OU4zRo9sAp8Ns+w5w
/vLtlIi2WzjjTM4l3dkltW3a3ViaMI4Gh0NbWQvbkdUJBqnJMIOfWHW2GnWYaNIBITFG/njPgQLN
nIYv9Vm2WlxAvQzHtYb6pHBq0pPOUiAdj1F8byH0835CoapZgS+HBZxkcbZ0pZcEZt512ZyXMWUy
J3oDwPmpx9ycigOF0Hwn2GBIZcu3AMOofS4rpk9M1Ul9AoOZ1bNu3MEBPNOmtoMLlk2DGtuZz1eM
vZ8B8cdWPKYj/pwLfrbbKg5Q1S3CHLMaSpMnO57ee0aCZ6VcWC7Wpfq44R0L2cMVZjouh7YrgFyt
tB6Os+l1oSEXlEkJJdE+DtbFKywwvYuhruYcVXL2PhvD38WZZnVmQwqH1wEaRaPs+1E110pU4d9j
rx/NMzRRy/op1REP3CkCyxb9FT1xp9DPCmQdfwhwSZNcEItw02idOqpojX7zzFYnS3u3DU8eeFth
wchKfOdjaZytbGc/Y7Z3iedu+0YmW2ji0eDfKVpk4/JIc3SUCXo5h+dqZrFBpSMcgQN3K9+Iaxup
xnY+6h+HQpILrqt//gvAFyLC9LZn48OZKgy2Xw7GkaJMWBuQYuBbFEC39H49yCTBbK230TY8TIRb
N/3SsAXAFnsvteNKNPqjlnhC1i/OUe9aNw0Qhr185fR5MVRmphBTcXu4M4Pj0i8VRt0l/XCnRai/
ue23tz09IWhwqha9pbk2IFYWplO2Mruug1LZ77wHTNMwm+sk4X34+lOs2MamvXYgKFvOJPKrac6P
if3+ZSxV9PAMTldrZluEcliCC0iZ37p/a98rY4c9GLgp7oWSxy11aN4YHEHppnIuB07RCuqp9kJv
bZ1EF7WHVmCpN6i7cMalyz/p2XvTLcL7ZJYfhAxNmsIkWpQblze6Ere4hIJTRVr3gxm5Zkrsz15b
ujrs3eli3QGCg+RYJnZ5qzxO18BelgpbtzVfKndeNHBnGOXOY0sV94I4/WzLk+Sdny9m1w5O7K/O
iLFDxZVo5S/ZUJvsnlcpfnOEferakVlQKzW3n8u4XkhCcxaWGadspiBQ/4FKsdEqH2+is43hKtZ6
o5xyhP5XGyFjJnzEocq6ShP0oi2ufRzFXs8JH28oKVtk/2YpL9udqisemXVffxI4S+wmF28vGfLW
KvCSwNppMVpV4mLgU8G90iCD1wYQ2spFcnH7tOPA8lhGOoG7aUMsGLjr+7dgstT0jBqhhY0aE/Rp
ns87hJg/CIO7T9+a7yz90RRIpnJsA0nykp5ClJENy7IKDytP6sgVmP3NqMc1fUPDXAy0ajdEeFYx
i8I8UZzWynkEtKG1Qe1tOUKmLQ/MGCGFQv3U/tqHYLCVxEBQOuaHRTB+I3tac4T/n9TF+diZjENd
yHicxcS26GiRm5Egta3E1j98Em+Rhjp6cbR3+VsnnkAjlkgTT/C6fhAwWotPbfEOzTdRjD4mEQgA
rijehsrR+JO8aEp9BaKbRe+G0wugFISvV2U65k+IpMq/IzUMbxv5mHOJEqfSKxqSh3bFQujaFqnZ
aO8fAswkKzrKTqKTZXMR0yYd8ZhadBD2+TwhCmCqgloH2BFzdTocU2VJ4cbLg1FRN9BpFUIor+E3
xMlSk0uogbA+G+XRUEEcqhQun1BI0jL/CUuJMxEJRN77WlqOuwoSafv413hfLeG/5BV6r5mC2GUW
aNDE6VsLPKwFTT15sRCQTOZJOCRvv7uqVV7OXFMVdTqNNtZ8melypMdNeYHedMUqgmvrvlBBcxuE
zVbnn5YmVAAMFtNjCFWBWiTrPqnPEc50BOgaHDnGSNS/Qd9rURKQZEobdAHYw2kdXmx15dhWvhwE
IZYf8GOWU/U4Sb+BmYiQRuA++jTF6dfHLh5m4xQxc/gZbDlxpCEYB9cPPCbvN8QH4XTdNwmR3Zi/
cMv558jWUrvq5/WP6dmiCjcBbwzQlPgXUWukaErxaKkDjaTjvsouUPaOaQR/0yzXFfXNYQvX6R9I
yrdwvLffaBBKqKPazzmB5xqNohhEYabILShTDdaG4oBN7TN/hkngFoda5bzyzneGX5wG/w4QOTpk
l+uW8bE3IG2CNC6wDc++Km9+LwgrrvPtsM3yPJCysNxNDQ3p3Wm2J6YGAwh/nTypSeFtVjJUH9q4
liwVeNwUGI70xycuLCLI842MTsieO5U9Vrx7hyd4BKtDQdTwTWDGZ63n7dZikQvNIspJOES8+fCB
TPaT3iYGNlnDptk35zSRxYmnoS+Th6UPbTichDVcWtNrYEY7f2mTUDg5MHQ9HOA5+PlvbaDe5Z1Q
9m9n28kAk95H/digQkGN5EEFaYqQduKJylFW8hCydDtRhFuanhjwna+bcB3v6Rx11aQiaYCG/2Rn
/NUNfT+vbXWerDSoQ2Js8vvns2zT0LBpSZKaq6SETmtExfYXDFjavjcOcwcTtbnmUxRbTmNk2Iml
DLmUHmVxIVc0GguqAGs4cZPfE65/Kqpg7bpJRV7cWdKbwqzXmr9fjhkh8rVUzkKy+VvB2CZ9H6KA
ny8Q2cSB8VUyTueD5w2GwdtnzJwqW79AzXgnXPJJdWam2KaMZCLzg6lnIFNGe08GPz56KWx0PS1x
bKT8gKetV8n3Lt8vUqO9hYBVRkOSMih+5gF6RkqFgr4EtD1W6uQhuB6lgCx5kLeQMdlIcjojcNEY
9nbb8iWoFiayotKiatpyt+KONMsaKUTzmTUiA9nx1mfi0ZKVc8xheZn3RpUfvAxj1FuDjOGFXPlK
k/IpfD7uKqFzHDwiuMweK21fDCvVYenMtYyPKoYAUJiWj2BQgKGKUIH04nT8oavM5T7XCd3oZimP
YoZe0sv4PeBKhoP9MjO2LkM4gqkbA7EdEr78UgtEEzLz0oCoDEnHvqWO7Gf+fDiyTqoqIodhTA35
WZrhLnvwvDhyClurnqhpWp0gT3+3OeJy4/A2OE8Z3QvZFAsTAoiTzlT6mRBYQUSzves9oKOr74cU
o90kqARLe66xiZBIqHCroiYQG7d08Avfa6LABKchqH4uT699hXKL02puvfSJnDxlLoPmbzFI9Igp
ZDDavGBejj14wg8WYVAFQkVE0UCvs1FSreVUV8vfJkesTP6hfW1LWSAdNEJq9vnjKHNcOR2tGfc0
CabLou2fjKC1F56EWfx+VNIPUbpbKCzqV0zdukTR25XKT/TgUvM6KtdS6FJlKK3YArB7xqfLh/GI
zoNDiM9AOETu1aWipshFvxENkfxijKeZZ5oluyLbcXH5zfQTIlbBJObI5D0jddndDJ/UrZy0goJS
C4b3DAodNPYyvMhqKGhKcXAsa2rmGuHPdi4yNaQRRi2tE02A6vsRHGTNG5uG16T82/UDDH8+dBRp
eI3EbDALii+YOQpRxyRpJSA5BVyrCzEmnQpypTvzwuqOhipuKFdR8gqGPqIocr0u3e4f6oCrBSeI
V84pOxT2VOBBQBmnyvirzh31rZsjCmk000nQtAV1yBcqtcf4hn64nM847IvU5cT9YYUbAD4G7tAN
veejdUE1SzADPkRZCAZr9inhM5Ybiw6zTcU7M1wijpYr9epy5m8d3+XWlDp6lG09klRN8clovzXb
YkDlSrmNWAhr0E8TZwlmf1jK6VF1ThDvlE7N9MCYO9w/Ioxm99fc/+WJi9VTAjH9ah3N+SCjQqDH
EOvlr91jPZXPiQAVU1ce+UwBRgPKIFqvN1y3kz5ed0xtlLlak4CzD2xars8tMgZHDMphwxJj+CfC
nLsh7cEZ2qm8VU0cB0+skNp9zk7UnN+cCtZepD0F+SDNiYu302bN1S8SaaNW0jAIlMnxfgG4Wyud
AURxGlh8Qa3jEXN5OFT+pFqWKdL7fmtyFouLTyuqJMLXsz4S2ndZ4ZTIiq3AgUCEoeyhcjlGd8rd
UmQyMU2dgaNplyuOirEWuh5xo8bmgtLGjwOrv75EphxiOoPGib8Tn5wRQu2P+Kcb6vkD2HjVhCiA
D3XIrznwdC/UbnBbhuAVkIhvAsSU8g4oLPeV3r0CFWKMckGt8nK2DCBTxr3M7vHJ6qzqDejkbtP3
ljUGD1XN05KihiZAoGv3PRqZKVvaTCPmI0f2D6Kig/B/0JuFJmeZeCo1C/yr8/EfjBceDS9hKvux
uptai/bLAEBXE7BMnvko3AQENvf9QlFmz8ANvrip6k1x6iPMyv85srrQW6JtCx2ZHujhb+qrT1E4
rYfxvi2OV8S5rC6uQF7CJhi3PwwmuuMgW+LJeV4LkukFvDgm/BkluYvVgbUkqT1zqFI2fd6WoM0P
OcSX20C4Y0FlowxdF5UvED9mbQIjO9V6mKoGV+VsSWTzhLIdus/zfLmQqZxbkn00qwPZhVpajygZ
fOjNoQHXsJAcguByLt1gIZKtNo6Nn7dwyvox/f0Gd44kWVdlH1CRXf+ZuxjTge5vHwMkcQzzwlfI
efYg6CKxJQm40lxM6b+kgNnzVQKR2uYy06Av4w6GjdkZma1I2/z3giivofltP//q0WG2tw5UGmNm
YSCAHA8PKQ47HdFf48jypYWnJ0lvlkZMUibXpgqhFPOzuaum4AdAYr3Ht82fXzqs8nPXpanS7WYX
TlFdZjejxIHCni72NxHeM5UGQMKW2fQZ+FLLhnfWiLkqpLKrO4jaGe7HpX80AfEz+j74MAkFSWEg
D9xggXi4sQPvqUjJyPkKVJheH+mTmY5Upg5coEoiXi6pRJnlppp+Zy57V7LbFYkTeyQRJocehBhX
14AesV1ajapgIysDkSmBPqYOlSp/jBLqNVjLqjbIzVxb0QxxdHzB2Jby7NMVBgcJ9fqezYonoCMo
HaXKGEbVyX/ZSFtU7p6S5u8jRJieEQ8IBi9wvOG/qaUkdIsMpK22+Jh6xhbiELq7C17pv/FWF8jG
6Q/QZv4GLa6sBy7AjSW8qkp+W7jexsGFLBcQWqosSRGi9yLFxJecQVPRfJjr6a76IwXXu01almsC
+gmkVOFWsbm3wDfk2Bmnq0NbCwjqTEwxh5BrN8NJqhRo8Ughn8a463k9Ng3jxQBAHLJiejr2cNv5
b0174EPL9jR7T6Ct3pggChFy5EPqgOX+8HxqZuTf8kq316xJRl0IniKqzy4oCA5X8m6oC+OCsZzR
ObyOBPYGqvmpDZ1uil5cJZbmFkl27zGzw4xybbMTN+3mWqTY920HPuhjF2JdB3Oc7ijZpcHRr32W
guTYhwjBM6gDjPpuZ+zzLbES/m0PgbggqDG8QhDr3Wal/EOko33C0ml0tf0utDlyzM3EvXc60Hlr
2pbbW8nsDXBn7HYiwmtR6QMXJZDhEMhtqlauDocNE1GhCA07Ztgp2zHYhsD7omabUHKghdg2bWU6
IWo8T+8fSI4/uG7+Q9KpamQT/N10zpn0qiGno+NwkquzRskMTvxVAoOfjb7K+Hit3LISnEAe0rOJ
NulIaYSPzvERlx0XvbAP/59NDZMfzuxj3xfit+mrBLPKZ0ldgZ5cIGjjlqHp5N+AdgHyrF1ea6eO
RcwstlydnIW5yS5rYe89qi1i6XFX2S74mfzc21TTbF43VycgQDTwcujbpoQEYJPs1QWXFAKY9tht
/ALc1xg3jJAsnoMv942T1NYAqs2rpVVrvHWMp/oD7yPvAWyLLkvF1YHSuoJu8AUxgwo7uP3soYgF
YIvybpom/M7vfZzH0tNCgSvCsKPTFz/W+b+uzg2dhV/zZAJ73E0lNV6w8+qx/6YwQLt2B08ZFNue
1+AOUKU4u3aiFbZ0Ot5ardwwXu7DVd73et3qEIoL73zQNJtVzILs4MB9dqijqwwrKvrGIfnIY24N
+dizwUwAmjpATRv5S32KzjeBcnSRQ2uvjN07PzW/ZyArvALS7sC/Czbs5Xd2f0ntSi7y73htPqk1
vAznhJO4qmbG7LnXJ+q610QK5fnUEUDpkd+Bu0MykPw4zKxaPDzM60qEZleOuLhB67f5yg4sStSe
wgHr42EixsLze6DJF616MFiJZVGCLUf2/5zWGyOHIK8RqgKK8SWoBcuzUoYqT9jG1SzdwlpxDy1Y
2k0JRzfeI71zWHDFt72LanYDvOz9DZy2TAA0WNkRvRFhi4gcO4gtlf9pwsxEhpHQvYVj0E9xwTCz
wCvw4COc01116Uh5CrlU3g2w/FaC5uA8AhnadJOENMjD8m6nteRlyg2vey/LLDmBVBjsWbOTyhZy
LIh69eK0GJE5XRxekSUU/hyiT5KTtVs+tKHIRod95D1an2Nhi8IpgZLm3nrJwJDCQSZ5kSGUbEpK
vk0DkbYp0fW3i/r0GdJ+apkQB2Q/eGByS6Q9wwqTqgcwnQVdRIC+ikxk4UbWljOyJt6xSE0i3w8A
M3RsV2QLDJvVRT6xYXcMQ30JXUL/EY85lvgt1n5AYT/qDnrtRj/GtrTrz1JhwyGLk7tNnx3mepD0
zCe6DHtZeJ26pFjtYLxh9cnlx4PeAthrRAPaGahIU36f+Wwjdo0UyjlMyAKi040NME90YRMAHfs0
4mwCNY+XkpX7P13Xjozw95QWnqU/wHVfoPTV/KUkpSIBVrUCPCo7FWM0lyfniHg/Gn3Av0kTIZ4s
FxJKSH0ao8zmPuUaa7k3KC8/Vd88rVzlKtzZQDEmieuRstl/ocbFELxW8EEFCQkhz9DAiPvUCqTo
EMQ6NKovoaCaknIqQq2zIjG0EkB2CS1WGxcqRPHvP2+xPxeOTxTfGFIU38jm6B5NHSUbPOw5/xWW
Tk6rzFUTC2QwwJjIFp11vvWX3xa9A4c1ujUcMbHLgVOslTgPmgOAIpX6rRjoVubRj6BEjnC80jK8
1PRU4UuNhm7fBbk1GVFawPeJAjAQSX6Jc/aoiGBrs4v5/IYHqLdsHXNapeBn1/cbeZK9QgHoy0C/
YJL2RkBOi7OXhqWsaXXRgfiYdLpHMDs+WLMmYg3xXP8eRK6Bsl4txn/8u8f9PzRpjk2XAUUUIWgg
gzsiY8fJkd6o1kV/ev992RUxuCirs/+BtCEcX9xEV2RQMGajkjUwyNQjDrCcOWfs1FAyDMoEmHrJ
qrRCHPt321U3pRMOG5Dlo5hCFEVAXHsejnPNuxrOe2GBzKoOmEC8cWAbSNNb+1bgd0XSFDtwsgTo
u3auR4MQXLzKxJp3qFrqDMut2Qlt/emWghTTonL3+Gafu44vAOPFSg963Kc78SlBlMCVy3ymB/6H
YQXc2MtJKYsiVFpTjqysrCPOKChjedIKKPwt22Z1FCu1iX6yKB92DBjHpbj38yx+6vRat638D96A
KIPaYfJXlKfsIhp9JTw4M4Iy7z7IH5ClzAaMYxDbsI/13j73RvrgXEBBjVlt0Ac7RnmNUpvhQfBd
H80GLzxrNPRvo9gVe6+u1+tG2AeK2h3KSkNX81hB+F6BEJ5fOOx8hpywpVBwXFBJpu0uOIGaL0fU
wro8OOrEwjn4L7ons9cvRljpK6kf2trsryTpN7URy4OOEZ6L7I9eDE1j2F/vuoLYOR1vSu+rvgEb
rh+o7E142bG3gTTi2bUBiAI0bH5A0IJAgr/jUNAWE4gkLYlUqK1RdcND0hRAyJMXTf+gCuVg1QSc
DixD6lxY0vHtso1tdq6bl0/iNj4TaYn7U6UtHqZDnB5wbumMDemhkAGt5pHalu38rThUgq87yhlj
bBy7VRynMdmDA0FpPPRQxAGKQB0ckdKSK/xFNXPpqI+bsH+2LPZ1+80xJQOIpoUIfX3twJWDlrkK
1Tr//04uWhT/09P8cOwp22SeETAL1xPh6lHXvXLbARrlASexSouwkBXkGhhEmAGcgGTnZ3VT8vxO
SdwPxZukadIZbN0LL5j4KonqPbq+CfL1vs4X2vHgvfTgDNwoH0c/RsHbgHDTL+XQvhGdcOQtg2u0
as1++uCKu+rhM/CYX7aTTj2CnhDxkRgZw8n+FrOZ6oQvUZhjRxc8ODc/7+M/nDDSzQfXpB+xrMTG
708pXG6Fk+7c+jlZ//ZAMVmcAfdZsLhpXFwqv0oyGHj1EEpZdRrvP+OfuhJoVNa0GXi3IirA8QGb
8b9huydOPfXa/6IYW7KboQukjNq9PLTTzaxekY7ZRArh76M9uLDReheLwEhnhZ0X1xjbgnkftJgo
3ZI6tNfUoo+zMEtQgvTy5eXmd4eLec54eG2JOIEvgDBPoxErhmPHOePcnWrqv+nmozimC6KFBHhg
OaSTiALpnPOQXZTfFjkjgb4ckTiAd7hV4kfcRY0mYugI0YwL8Gm/K7UiE0kc3EEWAUfZVag5s7tO
KLTFdFXz+YCc3DdnweBhfcvG+KyyoCmgGL3kqfqngb/ltw2NlIirLPUfymxM/zwrVh6pv1/mfk9z
U/XjwlFChSVHPMz77Ne5IgDW3WXGNBUweP/r0DeX/Vmn/fLH6Ad/OzlFSASVAFQg4B7X+TYQBVQr
r6EQx0t+qIEhlVpOLLI9n8gjsnaDzQGQUHZP8Fr9pXQD/qxAvIN3PGtRbPUSvagWoWK9uFqcSd0K
drZbyC0YkgzTqvjn1lQw0BdAb6kEi2O2DGYKMLnBCfLwrje+fdOq5dWsF+aneccBgYKDEM/5Rps/
w2gD2tpvycCRK42Msw71CWG1cBF2fWijXoaqhg1IFV19PEbn3UsnN32Q2pZihpU5qjJyduhHQSPD
6eui1IBgIuL9j1UItEVf4gA5Hr/owEmIi4yRn480udRPjBPTKu+xKOXENhsgNAGb9YRhcEgxJrEI
sYktR1z7o3zTLzw6oMRlzSwT14L3RcXbsRtfFM7HFn3PbGZOFJSoFccCIkrYe2G8dm5laKLGBoxx
WxBttpXv1Q0OmtfwkGPeePj69REmC4CuMtkiW29DTIBT84LqqQ7Mq2PSBzQiDRrrPA3r4rnvTEE9
Ez2GcmcsFshyVBUOlrKvWq8PV1gXJHd2j1OuALz892lALTmoNkiiTEzCBsq+Yd92ZlTOTVeoKvUh
YagTMl3U5BWPa0wZm3pDVzD/j9zwSdxMRcwTQ7JvEgbUB7/FO/PlUaR2zt6VET+Y9+2Bl9WgUvt+
serVKORfuP4w16timtyAJs+AGVFhEf5FAC5Jw33L4oq42ndK9wp8ml/clsMLfrQeA5UB6dXpYwWB
Kjl8GkpSqWgS/KEjBREV75mjUW//VUgVzmTbdwvxieypU45rpH5qv8xm3k9Ac7fG0WL8d4yyoTOX
Yl1obxAUOoHUWpAT+dW+JUv3Bs/U75d9O7e6v0YSkzFAiNzebRO8IAbL5CrQtV+K80M0wtkkjuyX
aFy6LzHDVkZBTMYjZuZfq3xqE9j5xU3o74UtEhaGPxQJoGE3PhcwowlLLKa0BgSqkMP4fezpK1ks
n2hT3iea21njXIxkr0rI2MBDtmIllGqhNqb18T9Dn2wcB7FnB3h1BTykrBO85RX1+KX7a/fSM/3K
S2UxmNYx8fVZ8xlLx6SAqvbn63edUyF1jjGN7qy857TBW0X4LAOotaH8i0hv1o9zk2xahc6TjO9n
nfhGfSetD1cE8ODbfeVbwSF9cdl0c48kMZs+fnzb/LDnysI0TJjJ6FjiI3uBrqUHHJAPHLmkXJjV
McUQdPN9Evrly/Tv0XJcxMAjFjjOnZt0x2NVP7WRWbD+BZcKM9DmWdkDMIquMYZpMu7tR6NA1GFm
BwrdqtZHM1uBld+8aAtF8ZfQ+4iTyCQdH5pzyrlz97GX27lCL0KfiQO1XpzhPE8QNmWJWXUvlOHp
kEAmR+Pda2wBASmbBnezyeD8/wHSp6NNOXmLYyJQoFhb8HU28oCGWZERTg8Js03VOZRTZrvKvQFN
fifLklGT9OpVp/a0Qc26PUITc6LZSONwNFVg74ZofpIrMIvKe8gMQ78K6h/nokeXKfsknV5sQ5NB
xY+XyDSgS8c6dhmLAMxYuRMKJOOjktmDe6npeqKdbN0enbQ7jC8v+NlRv4A3x14sbZGaT7YtN3rf
22+bT4X9Enu+S2brwHbqJf8sKF15R3qmBivGtfScL9v01DIbEc62d+aBURpDFhXF1VeYKFBlV4A/
pt5/IEExz+H1elzmy1bxhGfJsMLLNPmFy+gGLhKt9xKF/SAUscnTE6nSac4bQ/LLsmaKztoCQuKn
DRdLrD6gdwDA9hcp6p1DyXpX6yxpVRWwnJvzyvsKkiFwSS9jNtmc5Awq7jLRrmixQKZ9ZRRTxJWv
2jWaHDlPl6gWRbnvdVGoet7BdIlzma6YFzHdtJhcR4CTfDACJ12wGGTQm9ym2pwyRKqryomTNtJy
mkoHeRBzZzb85fwpvnp2A0ob8sR+et+DNvc+ZoqAJc41tiNw8J5XQd6XE+r3IungDxxzQ/3XCuVI
voMyd2w5WYFCMQPZvha6HBB9NSUF3fMkGABNxg+PkmMzBLhx83hSxXPgZmxv+7E8ntoZUsACOS1Y
oNSI45esPDXALW5VRoxw/OA0j4Eexrao9Xau8+Yt8PzLxZJD8o12G+wo2vtbtnSItknWQDjKfSKP
VRtxnzfOB3cFfwEKz86qwQkIAknR1jJc6Wc8qlqT0NyWaZz4On2K+3x4ffNPS+cJrVTdQB870kYz
CO6i3EnOEFknkTTztfO5seoTyV3umdQ9hU+yHgo1/QuEOtT8jTrQrSjW8NcV+Yuez0uR1QBugu16
0e/fHpNooqLFMdgJYQ2/3ze2tt+i1jeYjJ12zK6T3TwPk1hA9r+shfE6SGUnr+Cl7j2MBB8b/qYy
7fwP9S6Hphvk36tMVMACHqLkURqW389YtpT8brUArp7U6auUemHWfbmKB5ogvFTUUCueXSugNamV
frfrX3sTNLv9PQXQUgceGXUWSIvbAZshZScM9Vi5dyDXvyEESBayhLwNC34dw9zPDClseLJefoqt
h75TbVjBMHYaRgChIWigjDEavbarTvtqezT5kvrnMRPaPH4d5gSf2SYdG/zHqZwXnpVE3z2V9zkp
CRamcu7z7mQJlkZ1JR1wKREP2LqY8TdlqehUxp5d8oM5XhE+FGW+X+u8wIj2PJNIROSDUUFGEvtw
6N58GHKsHwEzdQOLpedhX/iCMOMP0yze+euyQ7zBmBp8pak/5s195BN1rEBZw5kMd0NwZPnHu+Ut
5RpK8YulO7R8iUXyPtAb80wtnZG8Hcw1v7orUFnbVjvGprdbfCXTOhRC0xPsZbAE5vR6uMtj7aPs
AWa0jk/t6kt/TjdnlZ8CB0QluThLRaGNbxdFP5OH8dinvubrl3X0Pf8i1XeRh3d5jwGnYJElVAN8
r484UK40I9kzh4ZEjCHC0ZN6txnn/xS9Fct2vHm5WQ1QzTJdbSa3lrt61vZAg9nDqVJxZ0Lfz4Ok
+Ygk7AQQgdv8+P58D4G3Of63G0G27NJA5nSz7QoCE6Dbzwv84SS254O/Zmgw+mvkETBb/OnRA0dp
+Afmr67Ehbi8Y4Ar5EdEYJHniP5vfdc1NwYCrYhU0O4cWwBf8EAN2AXEAoIlg14sOuQZi0XabW0+
TDO3X+x3j8h0HPD9GqLv7sNahkH/ZwkrIluAr77qx/btz0VQWqP98HekXL1qrOlyBnLC5dAWIaAo
bX/fMeW1C6BhzeFaGR6LeTHx16BZg8yXuycAAwhe9j0TrI5UglhVRiQjqFSenOWVUXStYERsTF2j
9dmpLa30vwrIfhCLQV78RLGEk2vIHirO7SZbEgALlZva4g8jeyeF7bnEOqUigLbXvJ3iv0SHWQoA
IBi90B3RYJoW64cHBkwbz/A8HQT3gXNCykoDiufzIDwIKGkJA1kbDbfLAsGYi0ShWHTxshFKEB8/
qTLUhVx+QCzUVm2555ljRlkagx6tP9e4HsbLKLrSMefd+MIbK31MzDCe3+fccYQ7APHb2h8ULgoZ
OSjP+AENoiDLBd/5NcJ+IfJl0E0ThMhEwlsIdf104f2tkCTXjIf3TSOWKHjQU9nvGQ8W4m1J0hVL
S2wz8huowy+ZzoE2bpGzsToPot1gMlX4eXeT9xPYRJeyzBBSLRepEmFr3g+Ym9vJaViVad1WmmCe
WiVzV2RNQlKPzBF57Ns3WaF6sSKqR5SP8vHU5d1tcKSQ057303NorwjrN6B4+bY4AypADwvEHii8
0IOZ0n+0XTdnbguB4Gi3cbYtt8WqGfZsYrciOCI8l1TiW7a9AdPPT9TfpJAHyQqTYpRqHsdnM8Xl
77xM8+/vEpEkwpGhN5PeszSqqRtCY9tpO6zR8N4WXPmMvbWwAj1uFlwJ3Pyt50kc13mZM0JK+eV9
cF4Fq82Uxgf7twuCIx0W1jmX0dfIpyVFy4KeC6Xcj2sdRPxqxqpP0KpaQFX+N0nkElEiIXa3TSzg
0fP49cE9iHXtLnWFNqL9e9nwi+peIt/Sg9vRmAclOk4PfpGnmOcMkDH1jZuw6oyHVXBSodO81r4M
X/gOj3cEtrxuwJ4sF6EcKLox+MKBJRI7Wtsez2YWRyZr/+4qbDPvnhlfF0TZleDgsxGucLNuzwuH
Jtw3cb6qD8cmHQuRZtiB7RXMNc451p79YZX1vJJ1gajDPYcTflhYLfrdjLGtJBb9eZWQYgrSK+6c
/Sofi9avlEG7ZzfliujCERRcmwgVOjRJ1WQyaARhyoyzlyrFJD+0W+poEUoqYe42zMTZO3CfvZme
Tuve/C8x1EICrxe7c1K/EpoC1XzcC2Dg1g79v5hJJUnDuG+w4A+gzJY2RVarcYm8cVjpGdTV2kFz
zDqi6D6XjetYeTs56yMlIVFhCLrQdF5oWkw37uA1CEwjX964jwCarRUKRM7IpgDq1aF4piglab5v
9RbjFlArP0SD5jFkTwRms+UFcM0NBMKdLTsIs2P4PlGEI32CTRrtnR3e4qpa5tnEC9JLca4wvVUQ
VhhNS2kcgn71aMtkqoRTD0KuN8STjxT71yRWsLpT33ljBjEyegTZdblJJxccWfZfyzQlddU1Y7zX
YKd0E0fNtya+0CDIBh70/xlJNacaZASysGkvnOYBbZIZcS4POjzBcYvVZe3U2Mm376QJ1iS8FqEP
GOgTm+XZrzOfPp9K+8j5hV/ogZByuQxYnid5GIqYHRosfObi8ihBWyKUX75xBmgfPgTU9CVJZPI4
OBWnsMyzLIj1zYwoR6cwzEfLvNsSiDrSrbj//jRslGmPCUIpF65Tyv3O1B/wO3nGwKr/gGhHELyQ
OfOamGDsBy7FSwujPDI2KrYwm12KHckeKcRCgHnAs4mxXOVmEXeRWj6nRKjxRzfwsvkB2mYTvUSD
aOdxzBpjawr0Catw7Rbz/WJpv228vShYAG93WaMLpL4joqw5vFqU5eTrhNY0KpTUZ19ykCPYubtC
qgtNZocaWCNkCJNNVmLG6AsCDwdePbSlg+SwUIgYvXd5gtDczKTycSiXB7Qd9JrDSDcqbMMvsHbW
uMk8K9fospogk1zpPCK9lz7nQ176B2sts50HZbra7yTNvfy6m55/pheXv+UMIlulvUJAZt+cMwGh
IqyZ+Izm/KsuzPgzQtbH/P80+62ae4fdl3Y1ho+0Y/RyBubt+KqQ4NRSLVMOlXnSWBx0u6mRZcUo
YY4uQsV8um8+XC+TwxvbYboGgyhoZ1fc/hFlAVy4EhfIW0eIzhdOCujWOoGuQhrLK6owT5pNPxg8
uikDatgPQcvVau9qhGksrTXc9Qg75fuyeLvbjmr9Xznj4JTiybF+ac6WBqBLW+Bi1gylO1ViLwiL
vOUeEF7WGvY20cZNTnL/5pnZndp8YN5y6cxm0qDvciZJVAgFfX7Uyb8VjTGYhNoqrxVUi8xmO23R
1zWe7f4TsNuBnosAPwdY2QO4pMGn6T9OCdkLU+oUiwxcTLzE3NuhfoMDUZz213g81B1NguwAEs/p
LXmd1mjW9Bpd+irk/7N3uncLJZ4WfVGxgwLV0q6nrzeEx7xmH/gxZrkv/MRMuNj/iyfeNPqumH+F
GyP8A4pXPWgVo3iKzWLyd+ZGTa/u4u5NZ9d7l+AOgTfdTbNvkiZZuhCKpsKEVPjEBAwFLkDT60ef
9oa/5+92hh+OLNjCBooNvk8w4ZD0EoJw8pV4gaxZo1liRebDdV91Ur/Awa4BpiZPycVHHDQOlWna
v7nEqK16EASCrSykyXT778ZaQIh1f7TfDs7S9M0U9peWPKT6nA4qm8gfp+vzSJytisLSqIHlYLH0
4ty7YR8szYTFL5GVp4aRSxkeTLiWBAZ+gpBLYhA128a9WrZ9yz8ks3Lh2g9C1/jYAVbLUacgoEB2
FolBwkVeD3B5wiy66BlIfNfOXNLXqmZAcmM3uoC8+7HwCH+u81+5faFFRuPbGySD/AcWVxNyVCQs
+MqMZ0XRMzqSVqqZwIJo7G/U+E7npBa1382eILKWKF3v0SalKA2hgh98zSgMXrPc7yiChYVlBDIY
2gxBERtjUadd+q3q3m4sb5YQzFKWGPoqDEAEkQt+W7nQ+40TJMbVUFfXNIE0+cNHuqHHNFd6XqU3
Zb0CS2pfSNOmA9d4+pgbKNd12pOSNIOMBh1yo7hJEtdfQf6xP6s/V/OBodgD5JCwm+DDTLNTZAOW
ONyXm94ORVaQbPqt6kH06aEvp//OjD+WW/bLgbhxOHd84GFPmASkQVRgPwCQmtQhUD+77SqoJ227
cib6fixKOL66gh8Mn8JX6obi0b6YhM8PWVeEYVsNNsfMLRyVB207xgOCsbjVUpDFnVnHsdDZtdHZ
zTdYJfkTt5ukbgD3Rxp4+C2WhaJORwuk5zEuif9tN8OkgfZGXCvaFR/qjyPShDo8zz12lKb3fZFM
xywPlcnSKll1tlkslQVT0cDfwgdrpfY6geGjnkEjsg9AWo9MRuaVeF9nFtT7yJcdeG7li0zb4rSP
JLeik2fMFltbLGtp1MriJnaLKuSBwBAmGQp6EmhzxV2ghhpC7Dm8Jpx1olUIfRDOoZwDu9kSuNXT
X1iyhws3DHJrVw/2UbawM9ot2M2pldaw4xXUDC8oUFIoTPdPx8onlU9ylGfjAnKbIxQEoSZ+7c+y
Qit5zuaspNzdbpJzlA6YpBBReSZeHqXq3JyjOA2iTGW+UJ/i9ZERWzkDTq95TyIXa9rRw0YFqwKw
YQybhy99S67/8jvrJq4MEg2WIcX+iU0DcNtYvlgSEG8JhJCNf8iPPLTMrd3iyJS6fsUDVF79kpl+
5bZIitk9qM7Pj9uKWJm8fzRJVlHUkCVMHJXjVDHJm4duT8hT0PIxR9QfL0wvKUWBHX9XxSwCCHOC
8GHFsHf9CMRFHrmPx3l8U9GSS0DE/WpxFWw8u+mBIYT2DYb/VbvOrnlqRuvBqB3QniAEvdkyUicH
XD2bVDKNpykkePvNkNQcvlqvFAjxiQgpTevJARBAGY5t1u4y7tSlcZ3c7Jte/34vTmtdNSXyfw3o
3yumNr9MgK/ck28ckLPOzAYkxz1naokLl/hC/0exyeiqTqO+aE03IJZA5X76fciDQ1mrOzpmqhGu
/tBfXnpY4DTbQQ9RY+g+ULxNLAi+qB4QivdJgQhSALqDjG7BaCwe3YsAk//Q1QNly6TCBae9F9tu
zpW64RWVA0+a1BcYzoNMjzMNgdfJyW7FQdjRccJjipRDgXG3p4X9mOLQyaOjR0kjn60uC3jP9CjX
ewpqYZUsviRafc+lOV+AviHuDIm6XOnI3J/5xrTcprb3/WZfxVFw4qfLDPeGZrmohY/tLmFQOjUr
HBifyvRZ3gsfZA0lTrYpNDZ882s0fHG+h05BpXXgO/VCa25PURuzpv9ZJzNaDkdRYwhnCvq6mvrD
aThmoM/q9bWvuzwNDS+B2sPmcn/FGFi41fat6LYVna8BLXG6A8JOqgkF6guRPg9Fse8yntfNcwDz
Hei1jZljNKtH/6m7yAg4wbUm4c2pyz+eJbPqGcsQW+BxMAIo9FrgqyZcFi+POwgyN8Hto2CFU8T9
mPEIBwMi0UOW0gjCaCyCUUzS7L/Y9zx64QiQ4B+lrwxBRCfq8HHN+5U9be6rqdA0Qj+RkQoe/NGg
1SCE4CvcVx4QRC2G2Vd+HxoP33AlTk78FE2JDDyrn/8IamVOHS0f+F9k6AijQQ1yqFiy28j6T6zh
ICVgWC3bAOB1XYjnNdqqxX6hQVeyO2ufWC9Yn9bmRV/lD6WkRnDBtXfcgJTeUuSOpYWDwc6ICo9m
DHaoj4+IuK96qeYMMXis8Q/abJW/nbqcJAX9x4MKiBJTLupWRCVJC+9geAuMMP1HMFxD9yKJcMV/
nKC87JgCVvVIC+UR8gw+r7way2dLwdmwA7YePU0dn9V59PB4gKbn2wUHIRC3hir0waI3zcWi31YL
JcP89XtDULV+DQKZVD1YB/vMJ7G3Q8DU1pWuEDKdSrNaBWdHElGe/mF9a1knsYGi1tkkcx4bwIs1
gHPqcWpZBlU7UZdAvYVzdwP9Lt+VWCn8+uMa7b1VlTffjpP+alKf+GBfDNkjQ+JTjPUd2a3AVVsJ
vP7Ue5CxKpSFETtk9y21H3aLx2IeHoSfUi8uXIY14iMYB9IBxV2N/1FyuCav598Fre9vnAs6N7bU
/IMcXlA7LHQEgJt/+gNQ1130Ak9P1v0h2ZmTriWoiTFnt9GC3Mq3kak2XoC+1aCWnJE7SLny6fK3
kAwhYrql1aKwVxrS7G6QZFAKgbM0hJ7O9vnbz6YTld/kKG5Hi0fzIORcGBFM/dt2wHpmuNnKM2GC
fcpFVv8ohql+32JHSxkMGOXpCGbOwl2OwlgD5Bc35Gr7s2+Eg79qaYSR8n/HWmB3S1IwnDYd2ZgI
NyxzDSu0USNFZcYMl+e+9E27fahc7huVoy/XrsRE+JQ6cQJRcxQnY60MYuGc8m76vFJN9Vy21Lwx
pENsUltdSjBDeR6siH5PGUu6Vn8PkcYCBlYnUT+Oer4suJf8fqR33/dHCJw4k+KvFCWyUUHV8jtZ
+Tbj4qaUm/nj+JdMQo9Sz3zbn6f70GupJGxh+y7uQnytHf69ebMAXuYRZYG3/hVLZXKRci9ChxP8
X1nhx+LAlZvPOGG7RuHak/hT+1ymChGW2XuBW4SlDKwShLx95a2iFUQ5aFgxxkQxvddzJ25qIhpn
wTQ9LnS76hlzp6Padtgr9+570RhWqC9AXPCqE7ZZbWPlO/95CpPs/+jOdJk3OHr6ZTR0pDj8qW5d
Q4W1wmNDXsKpqsr9oPIdm3U5ixUtLftNnYfT3XFFAeRIi4xvSlxz4fZ5FBzWFLteiWqvCpkHcgQK
+0q3zLqn2CRbgzIyVcPtbkbD9BoXyyR1suADEDp2/WLL/ceLUC+Jz/5+0hc06eBq2sgQpRC2ui07
8TLfDwFuU4x+ZKwOAet6uzBi3KUP59zwv0rCQ4TeUElUR3uAy8TREVdJNQxdD1x1tsE3Qh0aRf3P
foD9WudqrbK5YoH0Sw6C3bn7W0SrSaGsFLhp7V0YwxZRlLbEl14vbFSzAUnKYKgGxYfirZ9YY63y
mVn4ftbaji/5JP3YJ+LSer+qPtCrxQG0rxIt9C4VDdbB8Inrhv5L5dwxo5uArSqmT0nY1e5l2aWo
sRWk6lznfFYj/6fy4e3NtZTyMW0J4yZkDmS0U1B9QijDKELcY9eF4Te4lB7+EY3QsLnlib3lWSAW
QUKJqDy55GE3hqu2k/cQLtZOkzbnq/6zpcj6Y8EPZ9mr9RS2Ru4F4Rd0R0rx38OSo3ApKOdvI0di
TqBkm4hdYNOYQ2YC+lZINk3N/fokR9HGPTES8Ixa04kAsc/O7M9ok8FHqPBxwe4T5mfDrKJNqSGb
v0xxYSy113eMR9UntQbV9kGjO4Veui9f52/SY+4Tpmd91jGuABjX9ril8fBw1LJF7G6g6ANxxOGk
uWsFEgBvJjJd6eacAI6hhK+hlNBcFh8U6mjY1uUOEqhpmG63YBvrWxRpWrJaY1CgXSgLz9SnxpHu
1b4FO8gS5ZhHmBhLuk1Y9FnxcJBxPSSSpDKw2V1p5dOs2WmsrYs5CylJvLyAl/EU5/dUNIBBSYET
pF4UXC8//0PdmCetuQFfrFh/he0eXl52GDcXkrxK7BiMF1a/enFfkuYQuqpEbzEKn6KHYN5aUYnT
68s0LcHJcmbyenJpXerXXWkLxHIsDQXhaMbgAXbanrIKZgSHWAYujZ69DfNXEYuu6yGDU2HoQg8o
b2RBnY7Anipg+ufbkyJJLuQafdr3UGkvuCFbwDbN6Mg0vViet7PnXIKwo+LLVPIDOyGZgz0RzeiD
dIhgw//GnpbYFHddF6S5UQhuWemJUZIYGmbc8X5Rq8XgJQf7Gdo7LXffhO9TMENI3XSRk11fbGMC
SyQ/hc7vUXoVWzkCL5YEDy2KterAAH3Zsr44HMRvMmLteeu2KtJLWn2U0oHTU4nIqv0eq8LxwOYY
FyueD9K7weArppBH75Y4zax5mfPmPvqJRdpVExYC6ehCfmuI4ON3o03BDrmOpduEwbmpTfk/NxU4
Bi5lgMXrUBmjoYMHDrJYfbg6+1OmjSjUlugL5rA9epdHXCN+kBqK1PK333j8nHOK+QJExpxQpntt
rHAtxz6UjECGlW5qwiZyqiMAdZ9/ccTGBe/IIjyLcWDEvgMgsTn25Zu/cLJA2Ze8s3XY2OWODDFm
UAeKPKsc9nXTRNav6JwNDtLRQKYwK01bLDAAAhNIja6KCYOxJxsLJpKwnopj5O8kr8ZuywpFLm1u
swjfMRBgIA4zof5rVz6eV61o53VsrnWGj+YWmC2MnvbpHqIcGs3OkawG4DUSoauhUlYuubm/t3DN
tT9sH9rP/JakTmMTwFd6lkEVNcg7R9iQdMUN7L+Fj2h7fePEi+nMLjanJA770S6/E8nWmwkMPFCK
Ygs4bSAmezzIOGeOHJLPNspnhi2aGNvUziACzjOB/2T4fHHY1Y4j/6pfey7CZs9iwJ2t5ebxlxZh
dofI78XrN5VRYO+v6qCdO9JcHaTZbS6Cv+vkI6s/Oq5iPrIky403SvSgvflGOLFO4Fsb7GU1M2YS
Au7fk4wf7Am7mK5+t0aKtHppPnD5mtrDrobCGjBUqIS1bi32CsinP0icWcXExjS9RZBHidsfr+Qo
gt+Knp1BEql1/pFHq6hqCBr5Wvu/pXQjobKDD/CNbTJLOBXHC+QF1eIsU+MrWAD3SPHlZ7kT9IXt
KVW6yi78BElBxUbd5xOxCsYH8r8z23gGKX5aJEtMz0YdwqVoqn177+A03/0f0JdtzloTOhywK+nd
LbvnB2Hgi5vOdk2ii8pE0INMmc8ZtrfHHTdT19jgr2HJ9c/MPrxvzZ334vKLwG6VAuyNOgxeOajG
0hlu/0df+1Yz8RavOSzG9chRvmpYaTv9zZ8l6Wbp0wdIy+JsPioWQP0HtwzxikltPViRzSB3/5kU
5gwdxdjy9xt54uIitdYNZAV4HHABpjeYtBT6F/XBY5Cp1GIjzNPZ8X/A18Bzo1B9OprXuG55lPCu
QyDEqxVAlAuoXAnMgAOrdojYbilfNFJ/V0GcxLb6s1uFT+VFxU4fh+qplaymnQ4tOdre3Yl6rgrk
kjhBjTBqfbv7l7kwKZCkpHHA18rg7RHXZW0HDUerP6O7l0bZTtXmuBG+kouNpFuZ4gIpp9q23NIU
pWM+zXYUxfxjqu/GVVo80+8MDxdnNrceQtSQ5gkqTgAzmwd3QuuaeiJc51cYtW5RubBWf+POch0X
AeCaRGLWa3Go/zgPFC/Lkh+0JAWzVzq/q5eJPGqjbGKDexmZl4fdx6E3vJxACiVnxrTeWZlDojJ9
SkJYqvlAjaGEDJUyCf4XuY/N8H9ESMHXgBQryRoP10pj+6bRazZ8bfO07xB0a5Zfg+1Gh2S3ZYqz
JX1FjIokCpVvNWkscJECiiiiNznhFixaIq3IHdti1XDvO2peXRDxHpd3HgXhX1KLX+NEU4I4nc2P
hx7wMrFYvjLXKg5Ah1h1PFPQDDkd1YcYXmmlCVsfboKR8o2KFuK20Aql2k/IYsDUKFzipW+PrrmO
N7TcQ1+WBoK7xilPVIvT/Ay1/kOJgAP68PqJv5/rba7ZGXzq+ZYBZkSsPOjOUTgGYgbWlBWzYNNf
9rV+Fsnx5qHlUA4Yxt0nkXkfF9TioJn0oOabtQzNCG8CpjvSd9OqW/W97swl29bn8bPvu1lBnrkd
hgEcckvI8XJZm2kYhf2BU47s0aOakSFzkyoqMYVAsowv1DHC3TjnmX0wiW7G79YzA6vK3USbJuvR
sn9EN7a7uhim0XwrHt3wD5E2jT4KeziAgJKaorFI1DGTv/wvCgOJQiIK1Xi4Fo6/2vbacmUjftAg
QCYFMum7lccOHc0g7V2v4J1dvGqUobCA8apm0nLPN6n1+EOPaaFsaTRBZ4nqNx+fBznMaCILMrqn
70dZfupt+wui/JeTDvca9v94y3j7VSK4HJoQjBL9dX9EtYj3+oVZPM+XoD5hXw7ug1SnB8Sdk1Dh
NHWDjs1sFQULIyoEac31APekbMd/HnFbO3nibhjabThMGtL9SHDEBN4f69mhrMTi0ea3V1UvzKrG
2vTjCigf3EkWJLUJPWQo/+HMcEjxa9GROgLkwfJIkv7kW4sfcwTz6KnUWgjqNgfQmuaarMKhRmxz
4YVQabcmHFwX/i9D8Hmr1DjAdE35o+xSSR47ghx1EqBQnmSRamCejEd4e8tGqPENhxEeNfTwlPYg
DkS+9feLrhnX2IULjYEma1KhzqRHeqBKwhelDDs9l2tnGdYM7s1jmMOiCvmdFTqbGFtROgY70m9x
6JEgRV5IGqYuD2Gk3LUzDbjgHl6hES4a/Q90sW+xqEyuiLpbGIkNdPW+1KfLqU8VkVHD73cuhjXZ
6CJCksiE9aw4xPvHCyHizgAlrvtoz61OLmmt6EuuLMigPLFznq0suFPeplFRZQYCNjVeR8E/Qwt8
FY1RpsETF5KEAymBw9CyrDGEbbOi0Yu0ml6OXqLjbw8YgZ/RFr6aesV1W7F2xFUL4Zbegg972vBT
LRfumaJUIMbj/VIA1syvw+eSHGOs0t5DSfSFyemfE/VuQwUVPS0yXxLQL1XoSblV6S1fnzAyCW8g
Wmi7NRArIrIJvUhZn87ofc058X4UqO1tYBZOZokOrzk4gCxxTw91IuBVy7SurR5+s90zDsXYRzqa
adBysvaK1HyE6Hej9C3W74OxIipQf6HI3D9Ge6s0oeervqVywlDG4TQtYOTjibMzwvohfiDjYOZJ
k7ie6Q+sC53hr0fP9rfZCz2Oe4WVxIp1hELP1VqOFg2bc6vOX8ZARj4woHZMim3JF2W+zyWA/q+b
IzISB5Q+w7Zr+TnYQxVtH/IydDJ5hE3H4xaEDA2REt3zcs1m2tN5VUJEay1DLfFDVHD/fl2TjZ0I
e59MRcVsON1QOCejxLrok9JSHQrIJw1rTooQmM7zPkTtwIRXttH5K2hczrmm0sxr96VEcfQAKDPD
sa6rSXXPi/y/umOoD2GWew9RkaRI/Z471rXCdUQIhePflKT4HpUJnUZmigcQtn5Axie2zKzJirbr
fasP3ULqMS3cMSdEIHe7l3fC0Jx9ixtvFzjYXr1Wa53epivmhZmV+NvutBi8LiLpaC2XY+78FarQ
UGyEiaBTeUaoqkbc593h758rNpP/LS+RFJAracpC9MQs+3QSwe/oEjGSIcC/l9nyxBDidMO+H2pk
mV/cqL5U6SJkfGbA1ZHBUUm2nuSKZyPPwSuiJPidgahFiShbxt5X2D3BoZgsxzt4AoRN1mydZbp+
IRvT30DKkh2GF0qT8IAM7q2lvCK64/HG6RQC33n8tpZOhlf1B8FY/veexLjM9DXSKrRpjQF4w8j/
e+p7CaRljGwKV+kGcv5QqPeE5SHPqzA74FUHEfiM5TmzKWWeHIOauYvqEJ1MlKrXVma2fTdFwiad
8Ow8xaYYd7qioSW/5bVnnPgzPBWOOnUXbHCIdiTZFDnuNXthCTf4I7FyqgCFbEaE0iosFnIP4JZ5
v7PLR5foga9+8WFoRDUYE5OtJ0KyVr+Wxb6N70MIuADP9OpgwL/ZhQFPlsx54fAFgPgwiqxr0vuz
NhND3yJL3QV6WAYZEUcYApCg3dS5MsnK0pxFQtevVB0F3UNvtrOz8Kivk8BqreqXJ9Kc3kq83m13
O4/sjoZdUSdQ5TEgCZT6U/OPtN6mdrUOdchxWkX/o8qBfreY8Fdb0zscRip2PyDhIJSgL/svcLEd
YDRKMBYtLKEtObyFhj+4OWaKMGx2Zl6UHIEEZrxIdwFETJm6esg5jn/hx/Kh31b7KirWPU9wibAs
qMRqsHEBM9sjJVpiMN1dTsdgwJBcSPES4hkgb9Lr1jvri9vxu51kYBdKl1F11Y6rTgyEkc9Pe6ii
WX/zGIoQoJW9nu5GH0NziY48K1yVtk3pRcsCcbd0AXw7hOEB4ClCiD5F9y8jO35uCfu+BlB7oRY+
GB6olKYxpHN87KuFx5QnJHsxODOXmY6CbAjdvpcCmBNbXD/rZ9J7ngCr/Afn0Q39Jju3jsrxhD4L
r92ogX7XjNtHySux3pDDwjJGkNpLX+JSyBJLQcuuySIEChvWqOaqHGZtdpnzOS4YOofbLql4GinV
DyklVhgIIc5++SE5s3AtzXPaSW60nGzPevg10SWWO+4RkbIxeNgnIkyZfInC+XDDdvfQqsRYSalu
X2FRo3DUh3XqPET1JuY2ko1R4sRVso+Xxwpb6bg7ylohybYDPEYLySe+nVF3O04hiJ6mSXJiUdir
5fp1wjoKehYicaGVwcmnCIX2xqxA064nrQMN1MTx5wZwO2dRiVzwFTFWXBZm1qYim/gJGxe2wuf1
K8+2iIEm0ywUUQeBgVhY3EzQWpiA2LHBKHk5I9MhXRcOHjq/GQeERB6oFtBC3h0trq4aF+mnEtBz
eV3cBTBC3eeS1t4gJ7bkEcWpG6Ei0AA+A5hZMtnlwSEaHMiLjtO1f4YJxG5vL8e8KHoldxGb+k16
rS7/DLQPvPSx123nWjW7xy/z1mFt0TCHDq+88Cs5mcEaGMMjGIkUcRhGJy3nwZWua4nppf9oxif4
zPFVU/oEl3tlvguqK5QFf/HoeaqzxzeeH9n/rzj70kxgqLclhK6dF/LOCdpUTsMsJT9bCv5RmdTZ
N8tNkW052cyAS87Ogfo3v74UXV3e9S8yGvW3g6ks+MPYcGhtvZHNFcj1CMffl4abuCdpESPK3C+K
ojsPqR0VvTp4nD+AhD5BBdLKxxyKsCTTpZiJo2mMxvX7flY1a/ux8FHGjCSnNodeHGpuC5BGQ1A1
ZzVgSK3yHxrg/HxcAYaIHSMOxvFEQQGpFc0v1kYVwfc7jT3yM5Cx4fbEQdxj3lWFx2+v65+RdrGs
09PKosdmlgk+M3ANHxmW799K1TxQeXjPdKUI2nfLCr6Q3gtsEoDFlOVnG7JUxrJByEBuDxomT3o3
hevgK0nqkiR4kqJR1forwC9xFKKOpItMNS6wA8qjDK9s0a+pe6QnZ9sKrM5Xfv1ZhCrC96WAEKvW
VH7YUPVgY8guabpKgW4+kIf0Hn818IYtpcylcqqeoqSps2RpTCpW0wm1s2d6ibz1KC4lAiqQ/Eow
3b+0m195eaAVD1ij8JYzUseOThqw+erieyaFUbzbpS6iHn50YddlMLFqb4AdGAt7My9a0XQR779W
F0UXVsTVJi1l8JAprEYmG5p4iI0c/yRXnW2L7GaSDwArHaXTkJzmxcd/oogt1XQ7ykVH9uHM6dRr
Pr1ciwsYn/AIpFENxJ19wGz0/JpNuwkKLqYTsbMpWQWwBzh10QA0d1LAogAr+b3GcDJKDMSBBrzg
mMorpIwOuuSwsZbUvHvLgS7GJSlPL6UhFwWQybMZ1sdt0m1wQ+mxuiOPhiCW9kVqcLp98Q3wEZi9
6x7WS6Rdg2ps/cdY+dxLSPxV9ODP/t8L45R9PHHhKZQl9Cvuy74d3O7IDVyQevOZtN6OLBhRgBCD
SareEDqyGsME01wfdVr15Cc+OlGzDUmnV/6LBgkLd44oddlfPW/shFCj++GTYKHEri9z/BF5FLRn
Q32PAnyBL3rVFtqw4E7bcdbu2tiRjtGSWsNlAclF33yOAt1cnlW+wRlsUCmW77AWyf06XZt5sa1S
+oLd4fu3nDhbEvvyd4j0BneRQrJgF/L174Fbjq3G3s+xFRijf94fZ/Ansge7p/AHsHTFthjzraJf
3XH/iEL9ZXoxNOEe1vEC+/xTcKKDl4Ucso4FBn/t43m2Fww3Ng0Vx7YuJpOXv3xcH8H2Ku/FbZWl
raHc3+LIhercYYrCnJQ0CzuObGY4uF0WlFoIrPddqwWs3GFetucvRsCTV1OZ2Ivd12I4d8iNXfRR
IhA3wladYDd1ALbvfA76yxuzrFzBZdQwMxUtc/fbFHhT0JucTiSQwSyGBmRVUMDGgD9scgjCPhtI
w8snx0tXs+UdwvilI0myGOOfK9oj3EOzhgJiUUPedC6E9Y2iRMH8V0zRDiaVLbbZO2h6Xljh+hNV
a8MalGJ8ACGO0y8OQMNJk7LXbGM3U+rtbvtOP+x+K45uBSvXwjZbAkQGve0113xwK3VrQ02ICwFx
XPQpR3Brknklf1uYDwQMCEd/ib5wzddyL8ssQeKabHim28yW7pg+kw2sU1Ejclcu3D+R2tw5Cst/
dWZy680r69krTjdj0KhBqX/h8BqPVTh/fmo/og8Bk03ntCgYZFJuqPRr11v5/eheO3aXeN/MzjhQ
5avvwY/TusGXR7t/3Mswcd1EGgy66lrLdxRTGI86Qp2IDJ+KSWjLByCKbRthJK1FTjUtWwD50M9J
0Cwz1bMStjT/jSg0u97sYY9Y/c9Qv9pKioQ9+GW8+hcfyYUVYhniV1LMyHhixwbSt8GL56fdZKWp
quCR3PHhiTwIbuvS8a7VKBt9H9dND1VdYpgZZuIsCrXyKr78VTC7p8joGYfLvCJKzlFE1yg30W5B
EASzwqus9Tp1/mPgQ6cvP6OcxN78uH2FOoeu/Zbz2P4GyiZYcuBJeOKTpHaZvkVW3Jd64e0vFJzm
kdis2//8//UBp4YJ6rYVpWF5211ztRYaTMo+LNT8OiiMYNdJajuCNMDWlySjfdu38BdE+4y/UM4j
62LrcqFiaNOmNR33kptvUlevpUVetYp4qG725Fq5K+f+MzpuCR1HD79cg+TznQsjO7cpo9cNb6YD
PfIwCccVLC7NuJELVlw44xTEHlohj/pJ7cHYhgDb5NMC9A+ecGLtFZF4N0qSwZZChpY9PW80xRR8
RUbCKC2y2IbmZ99eIiZIyibUMro/S/aS2l3YcmYtY6LfR7NU5gLzeBGypcUuNjpb5MqWFEX82zt/
KUvQOfjz94ERIkcojtg6aUMTqIku0bZ/O6Cu/yi21n/tdHcATHQlXW70U2tJqEu/uLV8rwD+8WoX
npL7m3nlZG7FNI6c/n6qu84NIos1BsFeqXleNs4KR/tC4y5Ddwmh3K0WDDOM8vNCUB+Qj8KCLLY1
33Qnkwk7EB4PwV2WHDvDJPTQ1PQ4c0VBKXgFtu97Mx/3wfI5Zx0I/V5iQ2T29jJplrzYkSssbkv4
79bhl8LQOOxrms8Ubix48W8yI9Dd6cpVDDXuwR1LKzZDreFE3wIyvFKm+TvL6yTd/AXZEfr5vG/B
jEnDPE/HvaTyrbM/cBGo5/HxPpE2ZtXpnvWfb7RbIRbs8etv0xwjA+cXJ/OEfBFu9SdQl5adq9eI
N99UMRXh6RKqJropLw9zhSIemLaa95maw5Wqvv5xVk70NDXzZN+sNtw7KEbmHHZhfq8KMb6ZaVdq
vvMw+U5KuwQenclRq3/G8VVWSPlJ9Wsnp6EjQAtphuAreDaqdngFXNGctfevpHL1YUThtnWtCLXB
s9GsAkSJ6UJEzNXvby9s8t0TZ1hC5yZSgq+W2tvBacqnzG49uQA2w5XGDtMqs05GTDi9TmRLDq/8
zVNCMw/HlJhPr+ebalYki4t3JDrOjVYpDUA9Z2zX3kkAAKXkpfEprFdI8IRoYp4JXdUFC68NqRLZ
1TmZ3qI3wNeNdt3H/zs2W2m13PcG3HVjE8SEPlEKGsF8MREXHaL77+F4HSiKfGMnGsDggLgvph8p
OlGyXm0SbnVa5+iNQo81xQpt3gpm+qm6YTgXrZ4lH6stdMIDq8t5HS+NJmuFea+J5VCluW0At4Is
78SAhppW175/ZZ5Zn9gAIJnf784K5zWdBYxrBIR1Pwf2AK1mGD6h5uR3bWP3+WVdqSZg1RAE281E
2C2XskqYF4jVZz9RSwT728/7V3IcdPe0Sodr0SDmCsvedUpsz0ltZ8xOMPkFpoiWPcpVCKXlWYxe
QL2FkePb4rnwYcWv5Ih8Uwx3cH29qaI9pVwdn2B0DdyouvJe/57lg8Xs8qSttSwiFrFNqjuE0GRC
yaMdrLwwXxGchYZmexwWTnGZaHeliPpAaHWDmY8tNJU+q6MRu5jSoLIkd3wVmTJ9V6uvql69QQCW
khOceZ3I3n9Ugy0QqUpGXwRM7/kh6b8ACIhSuJRE9oqBiev+XBm2tDjdXgw7mLj6bfGQFVwHe/mQ
fb9OJ5GKKfo7aNO0SqCvz++9UznS94JHLuAsZuLVUgGzYofpDREVNOgZn5L4RbnnwAG4ze3AXtDo
EAcX9W17F2YdaFuOTrN/jtpH868XobuPA3b8QRXt2Uw+WMRw9K2ry2uikulCh4XieWSON65LQQoB
dbxb9m2L4IV5CNKLgjoeYbFwIEAQ37fwxyY3UNRb0Vwm3fedaZHrZzXwJhQ27kOjTQKGnxr5YE7W
43h0w4QmxI2zXAvf82g38l/titDqMTmIys3fkudVRgisMS+GUZYAk2alNRXxNCFy81PyT7X+RwSW
H8AbJI764TFNdOWei987/SDE6pjp3KUCasJhxIWcZT1FPswfsSEh0X9zJHg86ZTcch5fktCGsMxE
RvWzCuJa+ej9wEDtoDnSveilsztM+CnjiYYj+nfAEfM1aQeGl3PAXKJw0bKqe/+jQOTsOYB+VDTt
0KlZRxA9zhd1qaWGq/CnptRSmKCX9/lkw6MkupvNi+tPXOjbZqnyorNYsb1ftYeixisCJ7ssMprA
ROaRt2BlxB7zYzXCD8rtri4WFpuQgJiNX9TlPf8WM0w6M3tFgh0uQGzwhD26IfH1sQrXQJ78HXQW
DlqihIr09SpEkIBFMpIOOfOIxxMVCLOLrtTUcZ0GNDbLi9F102nmLZ1GkLjcbRst0mz52ADHFP6J
uQ/wd1Mc66K/wUPP9k6pMH2iZY5JdsUypwOGCNetuwYXylarRVAARtKW8qrMcSSVw1mqCNMxtPlU
a40mMvO5EkTY7yUpe/WBLgTuUgqpPh8TXco8JDBLqR9R80SkqUj5wki9X7R+SqG2YCDW/su7Idzs
vVKs6G6HTutA8pWgFLpRrll4ehwIiYljXiaumGHMQqYGR0qQn1B9sinvkoXsrqaJNmvnH1eOU6k7
pvEHIu+2sXbWWA19w14sMWoHfiVv0VfwTePpxrfkEfj02LQUUD6K1ZRzsyKcawFGTj9NZRCKrqyq
rsstmeh15EGdiy12PROYNBqneysgsudG0MMN3jDFpWPeypkp3yHYNJbsA70hSeysgLzvLgQV/Yeq
lvVGS1iWmeDz/nLW0eN5t5fGy2KHoRauS7jB5e+0r5Sr2BZCaEyifcQ0MZltwMH6baQwYBYCQhcp
TUqz5mu99WIEJ/smSULKUaziWYuNhw9J2lnBjuWM02s3ryq9pBddmbXnjJe+l77xC2tadsv9FEgK
H0d6LpeDF0WLHddqQg3FMHTEH3JyLJk7kv/Tw6dccazJcQSQbX80OM6Uj9hvTQ6WrbE+V+xwhPXM
uUbvNlu7yaqUeiNmRLtosVzWvXMgQX1Oxoof9/+z2rP5e/ZWQDcCWtvVZzkWdWu7wIO/7zJcoluj
dL4nTMWwFWknvRO6OYG4spXgkTsgB856muNGAk7uV6rX41dwLSsB0DmPGsfPHgKrMZjaVc0GbJB8
PVQB1eGp+S92kz2d0WGSXJsscwXJVe7MsnVsIQdhN9R4djp5n7b1F6kNhWx2Oc1a0Wy4ux4VYi/Y
ykxsdgMDfmBO02iH/1tMvEAxbQPDsRwp+o4XICyf62DobR0IW+/ZOZYWxpfdAvC7Dl7fI8bhQMv7
AWkX7jFh6PFyiSVCJfcirsW1+trGK9IFQ8EEHtJZhc54no6Q6e2BYHFKfjnySja1RYiBBEQhdgQ2
Up6YGPVcczCBuvxoRGFevY+iT9pcCyutTmWjqYg7UI6M3QP6EwPSy2okm2vTTxzuvzuG3zr5QDyS
/7ZRaAuh93STUXJikWXyK3a65yVGlAURak1APi/Om7jdSdBdpz9txLZlk7pF6pyIJBIkh/hJ8hfI
7u1f27QxLNwU+o5hgKCfVGSBpmCHe5qWYDora0zHrvGZUzDhmUnipJdB0Sg+bSAWwqkYcq66DSsX
+ZM4/iF2bNpnLJIS1LitOdVelmkEmwhn2cAH5NOV1HB8jEpD7SeQckxExRnTxC7HpvplDHZQJQXP
XH3Hf4G///r/IMFNFvOlaKZDokX4MBldbQu58mmEUsDsubDZ4+eaxc94zIv2wZvNE8iGWouLGOCu
3TumCdNj1iwlw5BbpRfTJp7+48fJqn0N27mmPsMZoiDK5+IerfRwWawdI8H+Ovrr7uhnZMn1IVNE
6z/ZpqPFVAr6tH53TOh4HwdKQKp5BRJwDGJbvpJBeWjJ0R3W2wL2ldFBJ8hJJKVWNWG9hDU0ssMp
x+HZ9cOK7OP43UKW6P40SS6WBghb2ifts9GVXWWDve77OC45evozkdaeaV6gsfjrGjEc1/Twt2xa
ynNjpKL9cN5jwAkpj1d4RO8XZMc09qN+16wLyfRgP6N04ISwb3OshWNzrFXgE7BBiG7TrQsjM0n0
JqpcOXGYH44ZHE82ez1+o8ONhFmYQ3Wm6ty12gnxtplbmOdxgnl98rcm6aldnB0O6mrecxRe5k5W
g1oPB9KV+JbhuwHsYCcGn/PEk6iQ0IoCL5vp2Z6g0BgECzjgcpyZi0FDvt/xX/WjZ5gQ5dfa1X9V
7C7YIWHR/YkZcaDTRAKfgHtJFvlhELtEZGmVfzoDwsWwC3K53K/r44cFq/Zim46yqb68kkxDIWzJ
C5sMTV7ZWFwK5oVspdhWR7ie7Ang6d2lXybI15qV5rBOgtx3S1SzbyKduQJ8mYrHRPyCN5xXVtr6
5Tz+qD2+9AtjhwtDoDHoLxzLcKBC1NhHrMB5fSGtfpv3rHOoLL6yexb2J7vfBlXSKNkVmjBgBFDP
EopMtI5iwPcb0bVtRqbLIG2hLTuddvr8+2E8+zfxwNDyEZY/YWSyaSSjxCt/OFJI8ki4GgX1QC5/
BK1SqK9UlLmWdrtzcTMTtN+RWOKmpSPd8E3RW4IhHzrApKhV3/5Ca598IcDxfCqDby6xZa/WuzIZ
QuBgTmLJhGIxUqGe6GmQnGzB199O4VnoJ5qLnYPAIaQ41h9s62q1VMbiZQKGByqACKhky+wjX0o4
oDvz8vKSvJlEa94nVwoYf7hZXPdpbxYgdbebrOrDdm7vlsfYVCxaXLyMuGuYoA4EI1fGQsbfQIJl
8CxYzAmzaQsYaATXldtY+L4+ajTHJsqJ+jOR0ldR8fLu11Yk0H1400trczbvVf1HqBlmjlu93hp9
Gsmb/6ymR5670LC7Qakeag7N5FKrjx8F0YurE7d87ISUXTjL7rw+4SfPfiQblfeIsQjJRb4EEEFd
61PgpSnuVQVHMZmmd8H/1gUwneNmIRTi7IPLhfjWwNdoir9FOek90kWVP4LH9KNfsC9ZZl8sLy/w
cqJShGjT5qSHqCIBKXoIgwrZOrYL20WaBazWT+rmt91FQ0cxVXtuV/jTo6TrVZW7MoC/Nj07icvA
mOsZaxBSBPXU9gpLFko6mq1WPy0sw3LpyyjHZWD0u6YxDzI/mrjTlyPgRo1+/o/MUhsRZNQPUkif
XyTvMtJDzgBpueVacJWjiSkiqCWFyRF81MndXSAHnw6IWLalkkE4hWwiuRzRaeYxUB3qC8cc+MOE
Dy9ABDHzmgXwiDXypCqdNcBMQml/+C4SaDU8rtG3sxOlRXU3939aM/1Gl/veb725GWDF27EMbiE8
aZTIvub0HeqKMTmlqx6z8z7r2NPB3HyQUZq7uI9uM1DRBgpgO5Jriliz2XMsG1UH5QN/ZiZIIIu6
5VLAvW+hrJcMAG160kS6QnlLLNhJWpLdRQ0XLkZXVNA6x0KvTzPb4I9jT7VoSEZWBvHZgANG4dgA
pcHI/XOC0Hj5UDQQBRNFocZOrO+JrD6TP9ek7FDh/4rKPvl9TRK+vBA8qnlHYq4sAoi77bdjrdvL
EZ1RG/QWqxxl0YMisXQQylwKhI86K9s0PP9zYSnz/MMZfahhJ4NQV3KN0nj0UETL/nhQiWkHdF/i
YAhLbaF8di2DA3OVvsdWZvM5WCp7zq/xBE7a9Gm7Lq6SJvorgncP0IEisgIDXo46BvKXr8WY0X99
GxwPOiP10xQgOgNn7kan9zxdQYAOi6BipJGfQXdXD5YP1h+ex9k+bfbv8w2jkadur/paJ60tGQjX
xUIa2rbkXkUCf8TtMjslzBax2aE0K0lV0EUet/QsYrm5D2To0SN8Cjk2ri7PSo622b/9VlmgN4f4
U6WznXMd6ddu7LxdvlbfHrVCPffmnjPuMxlq+dPdqM4mcLC5a1rkz2MX10ew0ZEHIQ5ZGS4IqgAw
fsal0edAwH9ELvRREXuly6+vmUI0s+P0Xvy31TGHOoYMU7E0WjQnKR+ACF52ogesAWcFMmhQwRT9
pFsW2I0MGuHJ/6iU1bIweQVk4D3W6UbZKxFdpaG0jBynxkpdXNZxdzDkan3DYytFtZFwt9Q+jUmz
sB/hUX4QGS+bsPh6APVd2ncWYjOABZaSq1O15J1rfWBnLmzp+q3YHrfINIhZc6FDP8fZALO3Y7oz
pLdH5X8U5X7X7vxaRObugNvU4ZojGn1iky2OvyjukFf+w16zC6dersaZZSAXdwDsXs3EpKUBQSKB
e2NNKzaxZM0P6P7Kl4RIx//fyBwi4c8QmIznK70RXH6AwA9aiU47OwBPsUou9hn7kkvRJOgGBdSi
T6buw7kGJ1jFEUM564iP8lgrI2Qc809+zs3exS6noKmnEMWR/jvO+ffuGIzsHUA+xk0+C0RH6xd1
W7+hn2Dn7gtO2W7FPMAyJEyrA3mSFD3TASJNrEbFgkfBLvS7L5WUl/4qumSiPb9tIl4ob3Q6yea9
bw3Rwi6MaQN+Q8gt1iyKc80X51Ts5BiA3r+xQeP0St+S394cllaQ3bgbpyI+6u34gDDcwaSl3TGL
OUt4Q4L6Obx7U+DiHujw7juFiqToSf+BIzBq+S8MMY2sTzeodjJ1HRG59P5idT+ena4YzNxBk2RR
kCIFOhef8upRpvpJDz8N6s2ft9G6aGCYv9c22+Cvv5cD/10sbqNwIhZfmjW92WdjQXjmBs7Ct86/
3+GKb/PlAfjd5Jucr4B8F29zegNxuhmZ8q1a1hiIp6HgOEQ2TlIaFUfB6tyZaaVKMYKC1n9m2zJS
5yc8MTPiZD5WgSZYTQdRrw73dE5GpDi7DW/GDPJDcTAvCNZX3JMGcLi/9WAqK/ep5c/wqWB9HKEG
lVQM4y+wGpnVqH9cuoZUCx6vOLwwUTZPpDOgHiHNEZC7Phj3fBMieLVXsQScASMwxssj/AIy8+hM
EI9DvLn8HrWeENA62Y1gqOv+moMKG2vettLVJxAQfGpA8NNYB38W/wLbvZaDN9r/dYL0h6AzNAgx
ELJ8d/fx4rvkYt3yNbjOTeLoXJuy+U9FuACSNhvDGTAdBHAwX6rmLgLWj5FHucvi5VD+dkBG7ksU
bFFKx0PTtNmrWIXOQF/hu5P9aFq3XgA+7OnOWR5OEKIlledvKE61yORwuURrmEjyq0FHjYivqLDH
AZkD+1q4N6PFX7LrtjJrIr/4JCukRjHl9Mpyqk208xfSiE8Hz2EDMAy9nP9TRCVqQcCe5v/o/Yvd
7ZLtWecMqrHYypxOmtNtjtbYm3np5uDrL3jR+4aBPn6S7G3CoAc0ZnIurSIKoL7q9dL+OCdNDUIX
6et0KfhTQs3p1Od1nBzm7UK+iqDulQtCWf1D3XL/18q1keqrrbaSMzs6rtJxny1EZnuGXuP2dv6+
QJJn4Kvl96qY9OqV6R9l7gMymXb1/IY7rezBSTfDDpUHY4c8KqfmyKMSiDWnNPdAb/KARd1Ry2Re
nopy5ywffY3jzI66W6u/Dxa5sO4uGkAMDa7zVqjeXMhaC6u5FGWm/G2+a3OjWLiVcZt3m4BR4TWe
eWDYr7dBg+JhXRXQr1yuveX9Bd+8x6HoHu7rqaU0BRS1OETceYJBERFUU1VNpZEuRoWCnu78vuRe
AUkeqfuZjPJ3T+LYqNaDdGP2sBEAXL0NMldse4GJckuOXs6roGyOPcxRC+lwKmK7FM8vPDYyTUSP
+Vau5tnIIcgif0dL7a+o/tEknYOLUpltbFIEFEn0kyg7DwYIF/1Jrmqw+0JR73sfQDdK37VB2LYx
O4T6QrafefeIIYbXAcEpXLdWlHeMQbJs8iG5kDMj6EUq3VnD2TBmxmTdOVrhFxAnXIffWyIk+IGa
s7SpaJUco/SJO80R0T3XUMH9fkmfO78hRq2DGq6r7CJwSVuHWCXH0FflxUyiPBVEwQTXHlL+Olt6
m018yrbeZk7y5BL6jgimFU9xMd8z9B3twqawRDd1uvmoe0/bilAi4ykVKyy5ghlJglQnwQqmQpwi
EQlPwgDIq9fwloo6dERe0rxjNuIje3LgT8WcyBUP3kgfQeZtf0tItivT5I2wyctIUM8mHi48tlcv
fkLlD/r3jshoTe4yLc5j3ko04A+9KuDy8zmc+mdxToWtAANvvMNo415TmWwvHs7hrisyXExYVZg5
6Iwh6j+KzbYa7A0UadOvYeM6WtiALduAwz7MX8R10v5qb8SvIUj2HewQjRPwPCgV8oWkPpSARu7f
dTTj0C9JOvaflXe1s3j0stI/0tvuBdA3QvhO+BpP1KMwOS4Nu47A+41362wB2GYmR6KUOpByIrlS
6nmJF6PmVXfVQYjnh6s1oV8iazrc0Z3emQBfphyznBM9AGsBfY+d8QrNe/KTWhxtz2FTmDozLMnt
jExwt7bcf/RcPnaY7aJxJnADq/sffCwX1uma6SBkofkCRn7lH1N5RyrDcXtaAaZrWmFkfp0Vqbh4
sMRfK00Wg/ND18imQL56sK5dFQqjJ+iV3j1UMd1RdcFve71dFwyTd6ms9o6AQUzrGjSyJQGOk9tj
pMtXdXUW7EFNPtqfqw/cUybyX8G/yBDCgSF7j56Hhsy3gDtzaOIyb65yy+B7wV6LqBhqS6O03zl9
pZKUigmi1a6ucSFzug+ec/icc+tgbiAGCEkKPWIBNMAE71GClPZ3LRCRtGPpD4elZClnZe73+hx/
z84VvSl1KSMRpbWa7TXzzPjg9yWb3wFrT55aTLqD2j9i+x4gJbOAIYfC7FWj4RFhMjIqWsW1iXHn
cC4UePlfPx3JDPKSo1e99YG9ujrvDNDJmmprjfpdJdba6nlxE/6CHTf6fj6SC0JzZUqB/xyLASnL
yWGYX/aIqxqG817fCZ+jsqoSz+/zX391eGcYAz04OQO0nJifnXvGdtCjUP9UnRJGMUWg2/FNK+Ej
QtVbwU1BnUOL1HdjzKKcaMTySTHuX0OaIlBmDEbhK5orEgx2QThqorv6TtZpy4sxvyBmFKxsU5yA
6zH2jYMVd2GjYAiW0wq9THdnhSwJLlR6mqjCb+cQUgqBtpCqR775r+aaim3Zkuwpwo0g+n+B/vTz
G1KE54nBtwFmZDFmqJLZ4O6e49E9x70k09rYJhxnSWK4O8UC5AjsDnMRjF8LpeOuTaSyNx9R5OiY
6sNA81gUOs5jOkyOEWMEVOtFcB5guVpH4JKhgaEr3BSwY7ilk6fDV2NWkFRctfnSnY9WiDFKF5wO
nwSNAd+cD/HE5jfXxJshp28qV9heACDWEUVQbNZwJffAh0AzQNjlR3sTv0cQC71KlGVdf7CQTPAq
K4oepxRWI/QqDTnk+AUg8y00oq6rogUpz0X6kUorQRRFpqS4uGOQrG17Xjnbn0+EOQjO3AfVA9cK
dlZ/KZu4CchTrKXMjsDAScle0s2Ik12NTqlEGFM/DiefKqvvkXQfRtBoSRsNnHHA0q+AIcGTIe2X
OtE/lOGTVrr+LBJQcqPT/llAMn8PBjo/xmQQsV7SqAGluGoqXpWYksF1n0CZ3XcFYJkM3U7iIG95
4V7vrHGPc/tejtkm+AvgoAqMSx1wpqNJIm+duISQ7OAXL3l+QTwY2Atl4XJtU113v3xDxMYYegzy
cgP8adK0U67KIRw2khi3K5LT3FABt5+7DHP8zqhQiFrRa2I+q86xVVR2WcgkzW4ofn06RCDhn2lN
eLKnWm6WtQeU4Sl1VKUZbfKbXOOgeocu8BlP0lSuZ6E8aw0eauZlFb7Ejmy7dWjjl4VWnLVgOcAy
Wqw+SgYsAtMGCGSs3CCwDMoutjG5qie6qJWRMS5rihGDIOWWZAs9bNKrfngD7b4POuYT/7v5GWL6
YmZMDZSVVhlD6LYWWfSsdG2JELiI4JgzAiT08dD5fCLKYhbau208WbNxCqJUn3qiUQHNjkDVTuB0
KTXhru8yXhJx61yryGrRWxlOMbVeLQllIGpBF5Luo01/TwwAcGxalL7CaYGgsMxFgX6fiYz2OYIr
B+zX/Qpb4J9BIiDtOllUxAt4ibCsb2m/aCeE5WgvHyhmHavJQCTW3MR/zHLHm4A5Ju1WEDd+lLpN
OqFDjxEr5WIoE1SBnDg+6pJv9VCQ7LTebQumgfbYRRNoT2R30S3HAl0oj86VA44b5ftubFQ1xn1O
9C7BERtuNJGi8RuJGe+HqF2Y7ctfJC5a75mBqAbrxDeIl+bmgCYYwPvV0rhwN5BuGrUV8HMjREeW
gQ2NoAZG7HpgkQRLWW9a9nA88xBN1BU2OqQ1BDPFKGKnExVwRZpB9wRCZ0skvru7XMwpw7NAWbOQ
FlMV1kvnN7hsscvoHE9kRQ9iLLc+RBw97PIO/tJ+HlcfIwtw43T+oRCkEXqnG6uC8NYQDKZM13hV
C+IbA80+W7CS79Gb9TJG3wGF8xe5cS/cM8MjS09vRZVSMqvH2pNmpxXv2bXZYtFq872nDJ9X9f4U
TmxCwPwLq7rnHHeOvPzza2KQH5XawbTlZObAmM05UDXcVOPMq0oR/1ad13OQhZI8igoRFtOxHp6a
Lod0wz6N1EQUHKsm4tUdI8LRTxP4T0VNuQV67S4pFprVwaQOf6J2XVeni6Uj30s2LkfXB5TZjNEi
RWAZ1gE5FcsbXp80EDD79gv02tF5/UIcCxEtYd0UKup8NdgP6O8hWulXcH8XRglM1GcnLXcSWGx9
TnIE1D0y4h79DCcWMc26tL937OzhpOLjCCWLyobC4FpJGhCc86ZbZr3P/jxtwSxpbSnbbfoFv+3D
q0ssM4nB3agTujFfmd818QOey1A0BLdX6O4z2Ke+ZykZsYTi//ay7Yckv/hXGYyWkdsUYq9hiNnW
4y5D/KKKOGpGNGOOyAcx9tLq+Ntkyl0N1PBKb6Nf0MOn3cttXE7tldoforFmtn1DX8BSc5wZIQiU
SK3jhjMa9I/jhtFI8wPhfDzPd6NCN/zGeiwxzZxH3+0o6ONeHZCs4SEbol7ZP9TXQZPqr+i/TcPI
MsI/W5axUYY3GX/24v/0Y8g6n5mH4kSyZPDN5595M1OfQCjvMiHmBQshGcq2Q/ElhPhdqUw7rD8B
bxevHiysRVb7Def5r181Z96CKToabIvlLBG3Knf9D+ZrecwQ1j7F3RKnzARzq/TlONYOww1Z43wQ
CnuNJVmU2mAlX3YoYTyIqPGsW6SAgrV9uZ9V6tLyTRbnUsgAwAfamkzlf7Bj9oD8Xb0xc7TCd55Z
HkUZ5axcBXWXu8NkdyKVP+BUbU0rAM+wRA9eAJ7mRBONl9odQcPuJjy0Nfc/JIJEhwFLIE0twzqy
ZsfQ+m/st54fKFxwVcZGI16YQeP0cVZSHTlAn4GXN+3TSsF8YrLLdYIKuUu/3TI7m1pqJ7D0wODl
TXvL4YLP6wjXIdmlaxMdtGvfoCmL6jBRoP7MFnK79MVOW1n2vuuxNxwQ4Rnf9cxChs8DmMtZDe3T
jF4sCkvo3+Q0NV1+y5v/KQDgjtnlJbSV87O4B4hP7NjV2O7r/Rg0+rzlbNH5bar9AC6P69fDUfEs
v7rwnjJeICAppgyBZelU1kUwAgBy/TuzD5OwzgMiutfQwFTEGvTIgQaP44AtTg/YoYDB7UX9cAVr
358XAPq7ii+zACj414CocRM9gxN+kmLdOpeh1tgT1LwfhPkr9X2PQzxix0rkYR9wefwjdi5MQ6iS
d0GaataSXcMrJN2PyJwkJ0gQ1krG/Wvnj0ww3PhiCFqbsBk31rrGw9W9r1CXG8b7UeLVf88kjdMj
MT8dc2dK1iHB4mGuEG3Cv48alAOGv7p2VIfVfWN/r168CSY2RpVd/XvN58/jnqhKNJYC+Krol0LE
ia22QQ1Zk8baoRp7+t3Jpb0YZ5pslntOiFfGbsvXiEhDhUA/Fu6ynSijOtwDKNJpSTPf5pebIVn0
Xj97DCRSmwvhqX6xkQxGKR4jiX9C9a/fGgf1sCX5lD07DZ4A1FO/pkQ+14LAlTfVcnY5ZCG3pDjf
iJ9TOwv1tc6dzAfJjbEa3vMjG0lcUalkMhuuLt3qUhA7c+FY0SYAhwSWx+OSV+/ScN4AMSGnu8AI
N/qn/wxoR8JF8kFfyqY0HIVy+2pf4xMI3s0YSQOL3kK2gT2IdlV9oAqqhVBVIjmXYUDq+tq7By5v
6Czt4ztu/KfrOqfb5r2yFcjkQCgGZO7utwrk7HGpqVV+3iXr/NJZJA8BOqw794V4v5BvAPSxuj4U
2m1Xo60FzmRTKSfpoknOiez5UbnhJpXhrM6iTKxFquCkuqndodKoq7mGJAouJV+JKerE8DUReLSS
eEw8ni6IukmqgrPmshpIXd+D70dBBSzXpfOJVvoeg6zNrJQPqutNQ6mfSfVjfnu907G4OnCBUVbE
1bQ3E4+ZpzXTz9ZcptCoJI/UDHTJNT1tAu9sZJw0Fn9SVoSs5NxzG5JrwDoWw0YrBea9IdPAJY1Y
l1S+uUdzFOm1oUELOiigaXS82dbPIU0hV6X5Ozjmh9zY1Epqcfp+NIow3Zio37PNBa5cNgR//OC4
zipQq1nxW4SMjzpYiz49Rgbxnx4I+aOs0iDePHRW/Mxw3z6j67mKIgwNfOYq1NdaSXWGM1ICe0Oj
62IzIeL2uD5lx7QE3ab4/fN+sFh9s/OAbL6ps99fGN0vT3p9Mr7EKqQ/tRaB31D3eqjHP/Du+t7N
jKsumRPVYusNLIbm0V8F3vnRitA2arsdo8WRCdM78tutg4x+nkwmKtGwk+xidF5B4Ei9Mps+aqkG
sGfriPN/2CticLKWXykOsAdYdGMT6R272ut125AENK6K/KDemTUejTpC6I/IvylC501KtlPi5iNC
5l5mJjXqS/vXB4s24zKulAFmDrmataY1mit+s41lzShyuAzidp8rPdrqL8y5yJhmuwDEkBnLVwS0
qlXmEoRB95lD4H6snqY9oh5NS2cHxT+i/CY174eEtvfT3QW4ihhlag1agee01tmg6PS0CZVmecTW
ETLCc+1e2QYzdR7LemwhiJ3FwB/6sGdo2S+U1vIb5+nmh9uRZNKpPsg97AhvGq/lsBPZV5qTiZrg
f7RcgknIQb/9nSibftJubhCmoiSHCBUnT2x77PASqwHai0lnzsxZFCzAiBqRBynfbXbAiEsEg6Va
t0Sij9ScxTQmFKrTo4sMUgkfkygG9moW54HOfa+XOhVxcwBoob2Z6sDNcpqqd5SzGEKqsB2RVsPT
m0n2YTx36rDAFxFNNeZ0vdGjX1NcZJfetcgYYxtkZj1Zz0JnGGILc4/IwRwyZRbMuCoz55k9azP5
ylSDVCh+HiqZwoYhEU3KBbDrF6N6I+6EJIRvS7sbWoxgmJnK0DQTCj3b3OTDFQp/Zx0vxSilB9Z0
qWU7qLGw63dmnDE4c/GtKIKAlo9JUg9rt12lLTX3yPh2KI58Fhspyqvve1l6n2LS8L0Nvrmga1u8
HZfz63Nx+zHrc+Czbz28YjlNGmwKkygmdzxVAgSffhG352Gcq6hDZ9H8kUIs/JwWcTR6muoIAgIz
xEXP1j1RZnOb/DMui4u5CBcKdv/mjMcDdvaI93A1d3gxS2ovvIg+pnykYp9YsW24ZmI4xd7kA7A/
N6bFEdKA8N/jUab2mXHRdLUNPyswl0eA+o4xbkhtRNRgbidZ75GCCzI14wi4LjNmNtxbnYaFNJhU
JrBHSb5RSI0rT76bwjNL777+ler3M8YyYHY39ZJ8EsJrDxUeHfZUeoKShlY9Foyi2h/SqCiRmgYs
Aatbh2OxV1we26WXp0D5zvxdkxfUH8JrDRb395j+xmVIpxexAATaas7RqwaFjyV/JrTU6S0EgtRg
W77ywWNlo3/Pg3MRYBBOjCMg4z4yGJSkxY8Sr+coGiVkgYLRDmncYLrgDVsZjV6HTNuX3QOKnmTJ
RyF7X44N/9M6kKnxtiw4gU/nurqp2DhIJQfXfv3acSNcQ3rUEWW737+grQQPEg3MF+Oeu4vwA4UA
zQhR1BtxrQp3SvRMiA12Lwj9qMs188tYWOxJY6s2+91aGJ/I2VroL14phS2Axn4dSRUQ7nl8/ZFR
i7h4taqMf1mmgM9ZrGiY040KJQmTLCWnDCDu9FVa1Pfu4djFPvfBuZSj4CguqfHl7Vb+ZK+atdr3
gBg4s7vtQiLFttgrIbOUgNab8zWZHbrUxZFyhg5Kblf6XU2aMONmzA4hbExUVGx9Fi9Az+sUqRm9
gf1N+RM7qSeou5egXaTPG2zR5oZsoNbsdbtg9qSXMF4yrASkmDROnQAXNffPSki5V1V76AoJ1anJ
dx3M0f8spfrkmcIJAxM5uyii8jBqBfxjzBVAEaB1+cnfLfxRHr4cShxr3IryUVV3pdHe781D2Ps9
Bts7y0Ds5vLtHqmXmVCjNZ8ZBKEPTaDbFiFRfjMckh3JpTIoC421gIbRQQSq+gIOrxaNMqIuCDHE
u/U/p8M7757RZRnX2Hy24gcDICbQw8p0sx6HQ+8PWQcf2qdtB4fVGeWyP9sguB1NIQKwtuNBfP/d
LLMVrQQMxEM8sP7+uhZdKa5Y8TgljjIty5aFcrYmJ4DraUYlzddj3qoncf9/8y8zD1jksnO8HKAy
sXv1X6QsTH+9nzD6kHbbJ0iMuw1SP4WwBEek/+UL5TOI0uO/4PJEX95uSZ7vcTwwB0Uzgp/wBljj
knrDL/2Sf20qGgzeqGWSjRBei6ft6y941VU3UgLY89QUAkS8I0n7+h77EHtFV5zi5+/zg1nh82c9
CvZ9K4E4FXorA8Kka3/KnU80fwfjn4k+MZwgV/mqEdSsQZ9Y9SAd5RuJcn+20tOFi/7qc9GI/6sJ
BLIQSxRs9870x54gwXU76UhDjE9ZumMtVp6JFuWjFSmHNL+F+YXPfnkyft2VrWjwQ9+Tvyk24Vr0
hkfOd4fMxKJgtzwRhpw9GEeU80HQE3JhlQYN4g3XMA4sccasigLGOFuPAA7J2/KZ5gl/Ki/GCGsc
ZcoMEJNTqvHUu88lvJeGP1cihQ4BhL3hUiQwgj8n/fEgc9f6KQ3zCYUiqFH9xcZB8gmwYqZ6SU5q
PkVdyYT4o2kgBtSYpcxk7oTfDCUdlXLaKyhh4wgpYPaekft3aVOa7S2HUzFVa/xxMlxC6bqjZGcV
qULZMsI4deo1tv3yoUCxllFa8W12KLomBbDFCz62BZcURAXpxxjXrypEL56gNyekDML/qFxI++ys
z/OYrQIX1s0fEAwgTjsiVqMI9LX6Wtf7RHAf+U0A/2MsqJvjDDwPq1NPjLchiP4DmKxpxWQnF5zu
xDhKW+Cuo36lIj+HuDzdeqe9xkISMhpbxTry4mrbDxx/E+9tZl1Fga4Sdpbuzhyl/UTMuD6dwRaN
jasVkH1OfqXPfbAToXmptjXw2lj++POQmDwDPz5IH8amE+6JnqCl1dkML990Ni/JHQ05KgOTOmn5
EE3GnFaA5Gjqj+JRs9aaNYUBJ+11F0eLmaUdXl2zQwz+QD7j/pH0zY/2/07/WApv8Tx5tjCBDPwm
H7e/VXANhPx/7rHhvN5u/lN4UA/EsG9usSrXuDDC1dl6SoD8cJZekLw8qFHCGsv/DcnJ5etB/xGt
UR/y994ZeeQRs+ujMFUIp8ok4ON8wqw7Jqv7ZWFrQJ6pX5FI61Kie1K2EjKTlaxo6+ujkvkRFYCl
NHek9UADGVDgG6X9SGuOrnctX0DrwBNK7DArmB0+gszzf8z1Y2EWg4Mrp1kynUMbDDSxIjh7fIjE
/stbuXM/GMKNe4bxoJqpRFhdQBn6orQX8HwCpKWkWlw/2PjCtjqFW1VCslGZtXzLyKOf5CI7J96t
x4zj9YMTdxZP2mNJZqmQqpfWMX/hxabPwoghgMoBeqy88En4ovYMHx4CSndu5vglx/PujZVg7yre
l+2dWJV07poZiQpqWnWUQj1jdQx34igS8ATTnlMncnaq179wiC0sL07B8iKX4TaUIsSLlCSaM3ZO
AKJCfi9j6yoIE0VFr3ybVdhJc8ITzgkq+yroqTqmZbTSKvADkEm6yJquO+4EQav3zDCGJ96a3218
J+s10KY1M+OLx6sgw+xkCge7rDlabdEiXmqHCs+rq1kIzBtFz2b9LLCHl2EHMfba3N+D0srgtQq6
of/z3PbD19A4fsN3+eW1CTpEkaDJa/cs8qZityst4VO/mEFcJotxNJI//oZUHsLOrEGgg3miaSTc
qz8XZ/4sror9RCVO81bSvADtKtyMAAQ55+QHe+0P8IJy0+Cx4XB5PTHkdwJi4ZGwFLy6FI5a0QDZ
uN7CEz2OriLfHlagy2Gbvl4qXk698MntSmJ53wY0ODepeTMiZiAsg+mtVqrN/DR6fivW+gb6NjDJ
58gbkj3czNoWS27XvJ+Lfq5sZfMDj1XKhsrVcqaJJwHGDYd4Hf8BYWWn/Ax0b/DIx6Zqts1VRYfC
mNU2lU22bNvFQroJ9+joQ68fdubq7SqovSRS8ceMw506twALVG9GtnZWaUYOq5Npe3YdjkPM9v6h
vk1s2bIMnIBXy4/hPC3zbySj9l5Bj5CaEzeobXaFsBnjCqPAOOF8m9v02XKnCS0rxpub8KCR1j4G
BdN3/oIayTl6GbPBmIjKWRizTsl3cGfjBQHhZglqk99Psjcxxdi32e1zKxYoR+19TF2i6trVd5sZ
isB/W01OenmppdinX/lR8+gEAFTQ0D06W2J5s8LoZ1HtQ2UQ0JF9KzihrPjhPVQTqcX2V52e2JKe
1PbtKZjTL7gKmSfaLo+qF2xdManfLI0oOq0Dum5IZkXwYZLYNQjIx6WK/pZtmLeyuGxxXlTHFIrL
bXgHfo3xQfAFk78b1ET0j+5l9w8QtQZeYEhJirEjLAQ7yz55BL1in1WiSqu8StvfTF77Pz6awDKi
kK+aMx+nbpj/LO8MtYrTF+7V1IMIEeVt+z51XjGrgXEydiPrObh/3rn2Wbg2A7CXnjjO6yAMa79L
vt5DdPiOxwarlw2CofxIny53PG/G93kos+NofTNpl3LU9UJ8T4A54yBSDfUXZ39NHC6147rDZ1IT
KkSdJVhcMwFwWnF6SIWy5e0SeTJH0ILbfo1TjxkkfRukNf6ZPShd6DF1ttISsYzeEXToe7GFBpVt
8wnUnC9eeFt+y7CE8mRaa9VwpsZLUpEtWcqXxWZkiMGNP3oE09JV8rFfc/HOR+Y57RJPKBY3mB7U
uRLSm1FUB/3xvQy7m1bxBqF7MfV+XOJA9JCOvckZWbCTUbVct030qlZkJdIjhdDuJvPNfdLGsFWw
8dDv7n/SwIdfuBOUuE+K/guBLwCd3sisPiehPkAblyfIfoPakHNotPAnL4MgAOArcWnL7pxR2smY
XGWXy2xRBZTs2qj3UCjSi5gdQWeDlrHRS1mCxMwYSyf5TDCxODKLofcFl+Uj9S7+42uEvXJK6fGC
ngjmCiberAjTzA0ofCyRHyCSJMuS241MOTfipkADxJWULkACP3LoL9vXUtek04Ds1+T7jLg1207H
9kx5sHmyVwpGeKTa9DPZk4MUp7AVD6V5HjSs83M3JZQBvPBpq3aR2XUEr4qceg0FqHrvgyqNDckz
S8b3qb5O/8ZtYZ215KktRfIJpzKqcTYk3MtZpVBUfadzcg3hNMUkH7w6WDa05EqOtBd5x2OIZuxS
Kzb+Qv2AQXCqiX4IJSVvFJg0dSlvQ6/XHpCcdwmpktnvnr2HR9S7/vBYGoMdtUqim6R8YCSIqPvg
z1EX2vZD9ca6Toow/Mk/g5e66RggoOcpYPtAifsBLsksCUeu2seT9RMaqmShUnJW3r1g+t7jMCua
Ewm4EGbvOSgyAEME1JUGz7k1Tzv6qwphYDcmM4lU0hMkb14y3K+0QuunXGLBQ93Wn8mAJg8j9U43
aYoGGMs0erzkl7Z8n2dyGA0J6gRsvzPxX3jIrVR/WMBCLTaYzDjrroG0Oc7kBDv1hsAznVtktNg7
wFUm8BpAf7jjp5HdVp4oDCdcDJdnaNIspluvJ2drBT8I8Uh9YvB0aIc2VlIjDB4P0nvcVz2yvYjY
m9PD2pFYnPCbRJFk0KrL6ng4xFRJKtV9Ekb7k7LhJn0TxRmswP5hKYNZ2x6t6wYbgBg7u/sH5ile
fI3uvUb2Xm5ZJlngPOSCq31jSlQERUhn+UefdULWpET1Dgx/vmscgAReqnJbKGhWWmhOUOCeetJr
Ss/xFr2mMNsdRR0ERuql+jGUslhmWmgUJ2XEVeBI6LYpkVAeu4oYsCfZTacnwAPF7M1JEHiryWFy
aimzXmEAnt83MePtMlNKvq70mH+4iBLeYfD43ULGIWA+6rPTsdJ7dtnYvAqykeQ6+pe3zbD9KI6t
NYwbHk/XK9jNc9TtUoPlYcKzR+73QibhugRJiJoeSKwrTwPtpGgT6I5/yRogViQ1NU0+rjCoW/uG
NXG2Ca2BkB9PH2rqma181qR+CYg1UtZvI48ACKh/sZgiWy8HWXdUU3SeOTFsH2HC7EGoevu6BkgC
QSErRgCEEJ+6w6FYjr/GadELZDxxGdlvhV5AuRnQx1eTQe7mqaTxPwqdIF9CDzjfG1Glp0ERaepn
wECKO60XXYqRUwlKQ0AQxFx/WZC5hiiMiNd7ALmWY9zFHhIs4XE1TeIXgd8Ikp/WQtgyDhJAFeVB
PhjDXKo2X4BXHI+/AS4dOtsO3B5t76jLLrBXO0ma2FfDwdLX9754r9t9emZ29hIjVOFsMq1x682G
nuUGZJJhgncdpy8tgoRWB+/chQ172j57tLHo+yt9pOGu+D4Zb7i/k0gJSDYAx+vzEVHDCZeOkyMp
FoUQG/5d7pCsNT4UJXyuGrrsaKUlan9rgDjHwk9syy3br9iSRPYmEWLB6i9eKpATq/akj5hdpI5w
4LiEIlqI5J6Oubsm0kyDbYzWF3ABxAE+DUTdjo/RZ38YViRtwXiCfJAxWOdbIaPL3eUWTwFxj2YW
aVqucBYOMXdxv6cXp7aCeQmbHPaCz5nFRRSyjVvlEDJ1UuSsQQ8fJER1N8OBh0B2I6Zt/HGF5Fdh
1/I1quVX3pA2zN3wgLbHm00uUeB/SpaVBXqPwMcZnd6ceetKecp13WbzzsFh54Vds61JIf7RH1n4
wMobFFEQRR+P6/OV3zYV704eEaAJHMziRKeMkG1uIodEWHBNnQt3Yhy2SAx6vBtWL92+GiS0bO4Q
gdOy7MsZox2xtrryqiL3o+F//ue/YhhPbmmObq+CRlfrRxK3al39H5HtAGfMuJzwg+sUBya9jWF6
m4n4R1Q7v1bkaq3DmivjKyHyHP0GB3pQTI5EbtcJcpSjiPozmuCOgUlCRp/Q6u5E8zFGBkgbXc0F
8AQ05MBRmFcolqQ10ZoWiGMIpyCCKQHp+LzQ3TAQuSnSkGGdwqk+S7t62ybrNUO/NaK9SoDH/9Wm
meQ/CI8+PhKqjWj1J3gYJIhfhUkm+npY0RfTICs8m2zd7iXBi4ubyQTdEum0KUG+y9Uwx/cDjUn5
ddYC4XRbfQVWyXreZlwqgQYd3ZYp9eWf1m9lo1xfEKIeGAms84JxYImV0vSeXD6PojOq0ClRkkTc
FzBhU32kottAZnjX5d4CvOPH86xAVJcMgxhBqvVcV3PrDKIUlvRue5T24uF2r7rBGOiBcT7dMfWx
7RMcjvbmLatTBpw/TNOXybMtUWqAdWh5NIZ/QjRS369aVqVt2n2RB3PVb+pPCRkzqEZ0XPuRTvnQ
vuj/Hjxz0Wdr7PWpp1Qs9S1zornFCFFJx7OTtvHDAsc48c29es7K1cSkVjKBig77nmmWTqMYMq3y
4tPCVHi7G7ReRbpaoQ95oZkZuq0ydElKldzwIauUpvm8ZOZxrYhjBRC0pTt52+5xhJvkBpVMNprq
UqbM81LhY6dJQ7XSlEVAh0I3YVUaQgMtFV1BACGcQJ+TrHQYq6IVgdfDC/NfqBl7PgrBc7HsysBO
ztHJnJAWu4ZjRqKp4uDLKY0visOuFVppQF5H+A1gMQI1rZgWLxwnS0X9iAKaUZxiqZJ6u4LbwnMm
6pG7Me/abMehr4+1TrR7BnIdsLc3Rkqy3K99OUl9sNzC2kV1fKi5OUp4gZ1cgcUYFUXAdOPtGN8V
f/q0FZfggtB1Vbz3elgwc+KkQ/uIBHmuM7+WXdH6VQrZ6pmgWvN9rlLZgWVa1Jg1cELpDzmrBKOK
+caxCDF6T2n8JnSkqgR1q1Us7R095NWL0AC9v2nnfcrrkjvBaAxJ7DMOWqqHeqA6x2W5BwKNxPJB
H10eIFqVdIVKubzgEyK8BQHRWavvjo7PSf1UChcnp5KXD0DENsSKKec37EGqwgN5ydqW3Ytllt4v
Jol3HMSlgQ7PQG18sUrxDgqX8HSkdOARycqPcQ0C/p8gAxMzF6x8ZzjiWcule0+N4hxG7mvXcix3
xZud3f9KZ1rjIxt/sgB2qjXflAAG1yER+Dr2xiPlK3VljtdJzQRirPZDZhW7cnD7qMbmkZi82Ul6
nbfV78R3vkhTFnvWJE0i0aXoTY1gQ7tj1pv7VAFVQvrMxhusmdTz4PRDy1SDYe7VkGee69tkbMVi
BWo0+g3prTfZuuBOP1BG2pw7+uMY2IqPSnfXe7NFT3eru91AelC+ChOosPBVw/C+QwmpIWNbnKjQ
LF2YrpgbRJq4v0hLokjca0kdH6H0ISsg6yPjjCG7ltMJjL0y5Nxi5632NAHyQdb4qcE/t80e5nbV
+fnVQd0TNK2h2OeVSVwGgAJvlGiaZE4e+HSIpYdC51RgfNizCWiOXrpuM+UyaUg6hNlWzOUzbza2
ripLW5KTZyKbb7jT0Ppji/d97oek+ZJ3t40iAyTX/2cppuepobhB1Ty/t5Ze48ynihB9RHo9uFo/
I6vTbUyaPthCgLvlzBw7CWkBw89SzzNcuLwwGMV0Vf/glxU2epmJ/60v9vOhfNyhwSNu8hi+7vlJ
ybR9SE5Kr03vaL4Iz+RVfojsCylnEz09MWW9TcIjeU9Qy8UpZqmI2lNNQTu+xSjSBUIvlcA/jFLE
rxWrnx/mWsC33y3J0ZYRzdVVroSi9eZSOF5zPhwmGu9vMFa9l8TGl4IotCp/tOT46d+nIY9h34ld
Y+u4+zQYNwvqLgEQuD01p+TX3N/HMjfZxWVuA7NN+vQLmQiDaAX6aUWkFc0T2ycestxgI+HcWFY4
LK9GyxH/5/zdryN5k9q2DDOquY4rYgcn71co1ZO7DAbK1K8XhICCPyPNjowip5KB32nM7GXDDHmy
3CgMmqSYY/NwqCJUBm3hZwEVevBwPRFgjaQL7Jta7hiY4eL1NcRpNfslpY7rPMM5ABKkZS4WKu0/
QV+yaPbj30Pgz9O8dX+lj5hGtioJT+rJPP31KTy/OJk55buAVpqWKf5v5bUYw0bvkO86JNyFYv4N
koQivRu0/GsY1M2ySgSBwuE8bAep5w/9bL5WMKWH8Sf9ExHjdkLWVTjMfui4GCti/A6xFs5K+Q5J
LRFOe0eH0ptPmYo0rQpsQx2ydkyMmeaduqaRhXZvgreAJiqEahDwSI0vnL/LclKI4Qiep0hXr4uR
zsvXE65wB9sKxWcpMDmXu9cVpukocY4McOZgW5FXt1BllT73yiZ9PrguSbsnlMP8eu+TaFp6LozS
Z5wvaYlU+dK6kcQMbrelMnHo7xwe4O0Qw6RCyXvL8F2kNj4Ua2cfgGqbEzWL7BnO3tQ5XjMpvP6V
Kv3SKVhyLPhCaeUkCSns+MnUHseeW4c/JKxBkhUs69f0ISnwcuf2RnZcLjWm3aD+eLoaiW3DHGID
925sc84GAjzNEZgKf+WxxESwLDUKUDNX3806BPp3iPzXczEHegePvCY7B4KMP3xJQqdHwmOPNgPn
n3CsFbEtYuVmV9wpAEYoLHznnRl+H77kREKHhxlnIE3Gdxlc3oEnJSb+Fmq1bJO3Wu+p5XbawCGi
U0bMc/131P9yyYcnSEbbPrk4D3furQcGBgdEuHuqXaGscKfgtRKAMQZX0MCDY1DXrzTeFm/khnEw
dsf2sm3kOGham7sMMqpjCW7RQgzX5ynrwxRDxGdqA+hjPkbglUVsLP0ydhs3stweKQkPEXCbon7e
dHBVqgqvhRRL0UMWHOW2x6ZIYFeRoHlRFBrme1FOMBc3IRSVg3Jys5TdbQu2FvE/CXZSrCehFdvT
MgGPw5OrzuYnIiFxm14Exd2FnPilf/r2fsAnd/zGaQZQ6/qmwp04JfuZPuvipClKVGTWFCTcQ3o2
R+3cQvL5XJGRzVIE7XxnSf+ASEEZnh3CH6rvv3yPwpbKcKsVCUaHGzfYmHkP9zkgWBfZp7ezikmR
YN2vfSCIGN9PO/NZ4xQfR8cS6SksJm2j79DbafKX1gyuX9sh4b0cW1NZgr24nS/nOYAPQpKvCBAm
kZDOupWQtE3jn85ForeMW9xLdjJl1/5bvEfiioqndkToAjE/7ZIb1p/iSEO/+Mfx+2WPgRHVQLbf
S57pUXqokgLuCNJXQ1zE7al+RBCNg87qwK8O9Md0WaHsO/DK+936PtF8FyXJl4YNrjMWQbAtJQtH
xH3tcIfH6u5W/OVliKnGdW4IRavij3KrsQsznvEwp6VfREzHbMvI8dLLHnXNelzAnbnwt7yKpWfZ
vDrMTCfeun/SrKq3YwPbiJz7QPg3DKd+0mxKxfyKWI+uNU1CWv7tsdOeZqgzNHjbVGXn4i3dVCHC
QkbuE24LQ1FQMqcvLfRdsn9N5pamUYJ52F0KJaY5txkBxsogo7Jt6jiIYA7wBJ9HFrzBeOrwHAjo
8hHCzHdNRLVsNxn66lYbk1XDcCKUyX3+YSFwT8BwbxIhZrED4OIPPFoiXYoAx2f0sdj0kO7KeaZq
EA00hfChSRpH3xoSfipYIeEA3y7QsmsxuL8a8GBpQ3gJb0S6bfsI3s65lTzxlE5fqwOexyMLGsdl
t6gW3Y1/TLCiqW99SMysjQA35yJbgwSxmYKXOOgDeqOc3KZNNkCWg4X9bJdrgZ4mH3r3PRr0DCid
lYl5wKJAYbiiC+aJ1lwlqobTAD1a0AvpJV47Lo8g9e2G1blb6sE9z7unHArPjCyoGH5P3/vtmLWP
WzqPTy6mHBhjGy6JHxVlx7AcDQ6Qg7ZQcZh+qnO+pk94M2cFAF2iJyT6y4YUHtvTHwDCMtXLDnPT
tTI6xYTSANqn6CeEi1viAgogcRVIRn9AZjH9KtbKu7Nf5RYVcAk01EOGBgFZA/4l/IdChgFOIEPO
/IvdcOQVcdeVSKWn9UNrqrhSRlNRO4yw9zcW3ki89SnjH2g02yvWgB7vfVbgZOv1YNUFkbXgZQ3+
sxN76bzi9vb4AFoU+dPLzyXYPNCY8IGlyktvTc/y2KmHQymALSqJSCjkyrZ6RGI3+7vqggeSjM0F
Kt+xM0SzJHQej1u2hdy44oxZakiipzALFqacRXK0vOzmqkS9Aei6vt5UxjCpNZc82dKXRykPMN0w
e8eXe3UT5fK01U6KhDE5hL+IxA/9VmiYomSxJBXJCv53dLocPZwd6H2RgHeH2CvousSOzknhIi9R
P0k043b74jdEywaQDxV+4Hi7OfnU1HDGkXZOEBehmOPaWXD2iupHgf+WIu4TJBXg61eFKphXGPdy
XRYLc9qWYvx03yBJad99DyslJyFnQlgHFOjvMUSz9dxOq+gzUdsURnRX8m/ronnPXWic0MhbqJRg
yFEAPgp3E+tBrZ87gFCLRue/5kpBYR6BAYUaBKrgcpitwKnEhV+PIN4iuYmQFEysLXyxytdBlY9P
6xiiCidsj4+Mm0CU/OEzksw8QtLlkVc3DLtQQdzyddrA2TS99vLcQ36l0eZqQC3na70agODM3rZ5
viUzwhcTFtbqEZtDW0csP526M5CRK08KLFiUFwtqFuHHgcTQ3aj8lnfGIt6z3bPjGk98ejz5khrm
BPn3qb3VH4qRCfwgTgedmp789jQUMMs8wIZPKWGER0qBckpU6qu2kQhBB3wviTeSPtb0bpDkC3fG
5T0a8qNHwDXXHzNI0JmDPt+54Ww3Ix7TsQUMP94rt4ik/yJgfGyMxYYK0vQTJc6VmQrY9waGBjgR
PFFIiKbVW+rSPZZrVjXuquKwiGrcCiZuecS7dmcq04uZqhT2rWM+RHEnJhkjUkm8NCkQQsQEVxMd
uGhSZolb91Zznu1nMulbmrNJlVDrzgVWMFJFWSao2FApadJpDHzinWBvlQJt5vfoO96rKOZBgRFj
mgtbkj+hgZfYU9cdVGTo1uOrvFFZD06LvuFat0LwAFFEGIIMqapJ0widGjGJNFl5tUh56qVut6VE
w0LFSst5+DFqi+ibPh5ICZupBjypVXAyrnnpO1FAysH3/137b6JY4NK8A8dPMfgkaMs9QyeNi/Gt
ZeU4umPFVr7kdGacs2Q8a7OIzb+Rnv8SU4oQ4bNFEBCDppLkKdlfDEZiPM2EtrftCZGUZgKgbHkk
N1D3UozhKFJ5iKrUZ9lqPoRYLdSftBT2BlSw6YnTizZcmc/Il+8aW5L1XjqoO0Ay+qMoqfdAFszz
akcTPcIuGx0ckCl8SIzJHzuwHuQSpMzdPksqeeThtiKErDp8H8Gj9MsqF9LzZti7O+jxFvuW+oNf
nPJ+cr0JJ7ZOyySxGQpg06wQJWu/E3jgVn0ys6gYzC4WHbwhsTgvK3KFJMhB8zfE6Nq0a0kV9ncZ
47/PhSe2BVCTw4ubBWxLLYr+6lx3JD0YSemMb6tA8e9n6+2MWtGiuZGOdGw1BCIOW99vjlQFhIMX
KvGBHwKgDAtelEx+ctQ8hwhqgwmHPOA0/TirgRM6JJrEciLScYj4dHv45kvJAqnVjGu0Jc++pueg
C/W2o0C1c7cwjbgPeyZolYTgo2TFVnvra1wKo+P/TyqoYADFk+SyjyI0jTRWRXfNYlOIkBCsWuZ2
zxXjPyDAYCoYydfKJ1nWj/9CKCctGw+Al4n0doyebUWWRxW0cJaCo4Q6rNEVUZnZZBCzND5v0mnt
gj0wMUSi17MF2guYOf0UEgRS5G3RBCFz0dS6HihkynjMDXLgAJjxF4+L97pce4W7oVGR12oYOmmh
+xcXU19iQONKB6jKxEPx+POk5ssmiUgCAixq/+0mMcf6cmuz4XoESnZw+bFkUXSazso7BFX/0V7h
5Snb/hSfs6bJjJWJDD56A+9fOeRCVfr+9W4Zdpq8Lhwixt0ylhPtzGQuckC7L5xtxMlSDDEIKlrD
Mqt8WIsA/IyrwMkeJkkIa/nmCiPeST3cK+qOj39jUWJ0aiWJ4IxtHJUsV0UG4an3Lo7Gj2IT5dxP
RYfNDAaD6d3DCQKbZrl7gkfPXrx8Sja5N9d/Y6joASbwZ/FSoP5CJbXqsnc5R5KuNiBiz2ajfLo+
zJkp+NYXvLI0uQ1maWt/StRBfNNUczOlFEDjWHoqNuXNZ2w47utkTuJxDX7QB8Cgo5boJJ+Y4WxA
T6wJPLLBLxOy2Zcqe09tl4fGthYPpExaDLekCMenEj9+fCaAjLLqWkWj7TjzzN0euVHsLmosS6hD
MlstXpt4JKOCEd6dcD/fherFIJ1SF0V/EGvpRZgnKpJg8sUkzunVUOe5lnX+Jw7mZ+zEDKFNRxYA
uQuew1UfD9mLJuJBX8227HMUJ8Gtd90/p9vRsBOq3SfmxpcRYfKpXxy4tL9Wk34R1+Lt/aobAkoO
7btOn5tFJ24sbQ623W7ubdZYd3xy3gLSL/8ClNKcs0H5JV6Hii9wfaICU25B8B9NKYEEqFbD2YtR
dU9NwtX+Qf7cJuLNwF2XSE+n6nbSm0E1HUH6aYMhsm/09SVtxOpETQPPiNWWEfb0eziDK3y3GG6e
Qoku062kN6t0rOIPovo83Dr9DFNcMfcDi4eU9W6n2mQJ8goMalQ/pebZL/PB+E/IigmMeEonVUJe
NxW3CrZRsF6hjTUOcVsk9ks9D47po6+bLSsTB+5JUKzSGurEipPTbZEvMB2jxXXM5GgdSLycdGpp
w7qIEWrO2wZplmqpqOZzpsIbgp3r1ty6VBwMFkXD01viB9GqfbwyAgjejyNrC/z1k2XlrJBkKT+H
aBZrvbzSwUcFUnUi4njQ4omN3/57OIbHzIW5+VNf3kg/TTMAiTNeucmeyDUFkv7K8UNEuf/gGbsq
931bkRUCn9jEe5y+90EQyxBe9B7oRxW8XE2+Uv4Xy4wHy3mj+1DW6LVM6jHQ8H7A/EeuYicWx8+9
OuCZK7Ju0B7xIi7OzFTslBPsgEEdo762MM867qXOcLrPPhoQ1mWE2Gj7NquWREhvM8iSPoqavUSh
/o2U3FoO07lgU5+Vm6YNcLiCzvZcHApzYxTVmQbINi9SNHs/0zRzzPV5PXXjoGAw4jgrbWLZHphN
4ESJUocX9ox70v/kPxeAcJRCXOBPZBEHihJsbVSAbBwm/5s4TevKykzdGMmJxpxHf84fA2RIlVtL
9Pt5C2url47pRR2bNiXUwX0qQK36G5yWesu7MAufsJsEmOeFz/VBzwkmoLEIvMtj26Cs3KnY8Ect
+FIpJ+X9XM7/PpDMjRqI6/PTR+UzgxwCp9KaeT3IK+xJuxoekbbpqnA7bdJAbG10w2yxHlDhquyB
PIg8VTBBseDPZ/44QjuG7WkfN62Knxs7TiCv/OtpstN5TpuORRAdU2jZrEuIwUtXgHtkBhCg5kHY
ElZT23hDeRtxUcENRxbvxnMsE/puFwF5cTdGKc+23o8hwo1cBmn73cPPepYwmYJ+HBDSsN3i+gHN
6CpMGvXAcU0e3pjVFB56a7MtSbOyeSO1AOWGUkYczpHa+gPxW/kthkGYaysVgUmnmW6MTkddacZc
fm+sFE42m8dSmSbVx+a4kmnOsOdz1xjjkpQiSQTmtljy2auQcWcK/vj654LwzCcvSDOkdnNW8ZKo
JAOoqE6eIWatZYh3LjRTCOMSIZBD5bTaqkT85Nwx9mWr7dsk7tvJWA8r+2VYLoiPS+kviuq7d51P
rMNPibzOBiEuDcPaYhQaYg4yMgPIAd2quG6n5YiMYHnRZgSkQt5k2FYEYHGwc0iBDemCOs1q1Uio
Ck74W1hj6JimJacjNZW6IKvjBKRQn4saUUPceb9E8S90X9kM+eAG8olCuvrAsG80OlJJYGhXQePY
kK03xsctJlBYTLLicNG4HxZWjYps0hhmJXXNAc6389bc29orE7h6IXAD+oVQwCTTRMzyHgnUHGZ2
pEd8CzyQiHdB++beGfFlqqwob6z46jv7RfMvwwXQVlrYM1FA5a8tirszWzHI/IhJlImIu0WstFk2
xoDGi+DJbxZBswkDAutEx3CMYpDVL/1YYQKhgG9Gg6v8ZCR+uz+d6XyREyPeMWi/4AnrieD4i+jO
sbdhDtZThRxSiBeNzEp/KiSk9V4vTyNxFCRjdiSY5AfuBtkVX4uM4P8reVRj20Pjo5WvDbJD6LS+
bTTFLygjy1xV7KJDcHgC+jsrl5nphsN5csceKYNfx0qyEpnQo3H2EAs7EPUM0E2iTE8plY2N/9oe
GAZwXMM5cEq4CX524N3gg9D09BYWNjpIpceMOm/gvWtyr7JKVfXU1mR7TgzpmMwTa8cvj5FfuRMR
lfCmEbOJiVP7FwO2KuoXfzwQuc0ExPKFw0euCjBnkMIFDR4PrpUu5Ls39rL46b39Bhm259SitWco
JdGbYNXpbhly/0SAmgUmCdKxKm1lKV4g1fx1Vhj7XK7TDtESj19Z4S8Y4KDA9YCa5QQGy5iSlNlJ
+E1TeeNEyciPP6N/cWI7xlK+xrK91sfGeRG7rivET/MIT6F4TLujQSGec1lL4gxZlopiUPFT7p6j
b+Y5eOpBxkHRTDdSsM0cpw/jjEloIsU7ZSxQLOer0iVANb4h+IHHCqjJ0xuZ3Km1XFtOQz9fM9fB
y2XpalHwCNFC4BNq8WOXVmZOjn6QsHDCDWdilpjNI8UDr6PsbyHTo+Ya+l6TZkwAhzqq1YDTjl3f
A4rD8Uec6nZ6M2EldvxmP3QZroXUF0+iwy9hcLwEehnQea1Uw3eMSXaLuAyuMfmvBhzj7hXKs4Yj
/R6KC+/8YS+URTeEibzZzEsx5vGJRIB3xaEvAAY89GZp+DUu1B/ayOX4BHsTE6VB/1NzgvkujjPa
ShnRcZjNhiWXDW7nriKeeqnEJBJKTCwAHDDEfNewg9zlB6GM0wrwAisdwM5iej+290fFbc2OjmVo
Xnn1KKgopOJyT+78hyEiUf+qaKZPagu6UZg/kczv6sIRFwA91aIzprUEZ5uAJ/N64JHiCGbW2Hqy
wWboLdlMBCCRiZHtOjv/dNeoFo54ufseXZqLCk7HTGWJjpaVlQWxW7aPyaxkH1xzjMgjmUkQnTpJ
kvtfIZcD5vtfa5e/YEHMN5yNQLGbL3pHpf3mCsoBoU0HheMPmHXgiIpTwFVYsva3O6fwHhmtPAR0
LePzWCqUzwt4PBIIPHOQnBjZjrjRpIbqWfNgDzacvItrZPYplnGqFY6nKHm8u6hVjtdvmLK2ochJ
onC9SuMldQLz5f72Z5VBt//jK0Mla+mExEf0X/HkO77FSo5R0yrWWjFte2OM4rn6dHpd9ZAebFVD
tE6vVF+uax6G/N6qI8kwpjoGkbwmOpYQ1rTYQ20Gxd53YhUtSR0NQXPGRpqP+lZAT6JYeF9gFzno
L9lWraVcBv6NK0vJ1ARxzOO+SBjYjaCszpcuU4toh3BltSA/7d7C4n0e6gUhRvZquSIRLH8bok5V
zNbsM2M7IBwI+PqNb53rceoUmdK8I+uXb7+Z1wVt1EQ7a6h9crTqcuizeqULDw6OdZ/Sy/hVjwW5
fEXVque9iwk3wwj2mqzHys4kiNOUyC527+wAo7LbDIqkmgPVKtj0JOSSayLsvvN/OajqFjuaNR3o
PWHknoKYBXDM1+kltCU1n17jbq43VwwWWr1f5BVdnPiMBAsED1StrhU1dR4ry9pc7sW7dWH7ZuDq
BnF3++6pHDTKiigdj+iI0O7UfTuZ/UhbTiU28MgKa9iCk08gMq5MGO+wSseR/qaRnlQJ0KSW1+9v
+lyfpFdm+gkZG9B7xUTd4IRAVwijN+AhhR/SjgJ+JPRHCNifWey5S7gtK7jEJtmL5XNHMirv7iJ7
9cw+YCWSL0u9z8LWQXFhdwoDJcVd9MatsRudd5zRSMTzrUBgvX9v/CFwKe+qVbUyyxfcdClqaiy5
EeIdXan17E51mnKfClgiAveJdhENV2iR659knO5IQ897nkkDXNnQn7VbOkdTf5qBWJ5kCuTtjIto
rbOGDYvONLmcO1qOBrl01B34xr2ZBB2xObTMml2WCFf+5nlG5NwI/Rz4OtkOwjr7Vqx0+8k+uJRh
stZlU/Hv3EbUY/63epoOJyvQ/9kQUrKlJf1y1fJp9rCFURo6iXQaJHScTftRgwf1U22L10C6tgGx
iVTZeWZmV64p6gA2rbfGsUEZ5dWvn+oU2Isic1nhqzVcY6NClV52T87uigZLVCup12pKq1Zgz3gx
/9BmyrsjenRZ1i9Y2mOroPSLND/t3JCn2Sdm4jUFjQC/r16/indGJPIhbRJLdxls2jDilm5qCfBb
GwCuhkkVAbtY4hIWWKQiuXHBB5yrHxqeEo/fySfrsii78dlqOX+Kn1TZws/sSZD4AcZ5ZDTewQbm
9NZ22rYN/+YWdcAnzNX6Jndwhix1WSmGjl064DYTTEOX5okMcyq1QXBrC00S1qQ7BqSXZxZLJB+y
RZmfx1qrDtfjSBG3tTxI9YJ14f3v3RJytgjMJTOAcW+2NmFAgl1TBUQfbw+76CR7H7ne+LGa9P3o
tCribMsAaMBnZgXUXP6e9Bn31hkk8b/T4Ya9hn5ppFsSP6q8ChhvCiPxeFFA08mUSQiTPEvzuXBG
nX4u6sl16gtBfb5qorHu7WTkErOfOCWvs00vy+0tEE4jQzim/wNaMjaS8VqF+liFf+B4js92w/DZ
RwlRbsCZz7Ek88HufEkUF6gXrHgSF31XgyW3qKitPO20G0J8+IXQLYGWFK2xQimuR1Wma2k2M09V
IMq0l5b58UXjSmLQKOZBZ5clXRd8y9QIGucUtDZL/zFHJ7FiCMRBJPXyc60TPWXcaezV3SxskU/p
FOBM6xrSjAAEFQc20/AeD5PxaVC6FsuWjyvBWCWRJ6do5t3asr72Eb17MP62neEMZwmM8vqunsO6
t6MzlRXspNg44ehpg2Ycn7vxnVVm2Ue0DDatEKoDO6Co3g+v0I4uUx6jN9ex/db6mbPYZGiJrMtC
wXgfgqUZ7sooeHJntNHzaV3NSugYQU4jUlMeaiqyGKTwqeJfU3Gn72wE3LO7IDE3bQgiuOqFD4X1
04A8dA71N+GLmLNBXrk/RAfz906PD0lS5VClO3AcbH7xr2R7F6vC7Ct0v30i31v9pfhzvmOJXjmm
EPYhqXtqq0bBnmZOrzt1RPV0Tzi1qSDYIj4QdluRJogh2HLM5fVvfKgxNJ00d9zVV17sdIIBfW4u
0vWN3q8zOfaNz+Wse/wXFgcCdmVjRi6lBbOnL1fzqQEWVt6fntpSHUbYIFFErc/5k22vLO9slq23
BivYJ/5SfcV2CeUpGm0Ji7/p1HpdhP+ujQLcgsZt9g8df94EXHTjKqkNhnsIteAVi0GRRpbwrvXN
Hht3inJdE1Ju1B+YzwhF8jVg5TMbcTC+p5IztW7UXZutv4ttmRuc5HTydD2NdQ6mgnAYlyANQtND
QZAj2V39kt7c8Pb71tZMIY584hOO0LWXP1LC2VJBmmf4C4Zqb5nL6vw7H/cRwwKL3GlQwoz83zFQ
xGW7N/35BrKf/mvnmKDaiPPRjdj7w9BOjoA3DTQONvKzPY8uEJq/jAWUB+solvG63mTm5BTTZu0i
sZbB/v32US8xCtcaM+QiwtTXmeTegPEehjGuZPtlZF7GA845ohaenb3Oe88gwUBvkWKa0ltmTz5N
THM9j3vp/90NTvl8S6Q8UmdW7mi5bFopg6giqdcI3IKO+zRNY8LAPABlgxSGYCM1NT3Y026EJ6A3
PgPqqtHbmLIRsYQNVJS+lb4xsD2D7bPq+6Riu46oVToWfTvU65avddoyHTCZcl8PoCRZECk4dmnr
Lng0jeTC+vN5MRbv7oQ2JAgu6x+/3afrX4A7PtmY2dUhSQBGbNgnlFxNcG6jaPTUEibE+grU/fY4
M+pjd7mSED7zndhzdroW7kq7EDAiSWrBBAZnOEn46u3b1lbNtMCjygcl++o+xX6KWf63Pc8smmG1
E+XNDFY+i07qSKu4hcGFW/mGY+DBrbntfhJa4cPaHlXVUiEJpRJunuuzVHgva7YJAmUoEiqYAfbb
Yl0zlqEtoYMquHOTsDc3bm3qJ34FNlG4tHmDPY5e8PEn0DPSfdTbZNIDdzXJJAyk9LzrEOXBo0Yq
DNp8hNdT+1ci2UIJiJYkDPDnZjqr4ZIFu3/BHXnEs0752FbIXyP8nOmAMflxW9ekY4jd4DVhTktL
T2UQBgs3R04u19wnUiISgSuilv7vZjge6zVndn9nyMMs8xDvB2Onh+Jb7hndu452qRAvw54ob1mR
bCiWTZ/wQQZNCTTId+sQcQuFwZcplniVwXOY7gm7v7TdUxJBfyMpWqalzAWmxhRZDo6IkE+Yh0pn
DeDn8a4cA94/cDh5/p128R04SRNlhidv/51jP04yPshhebdn/5gXPx1Z3HAhbWurLl3QI2HbpEPD
kIouGAAJra1nrtn8p9n0BW6QEIUkp3vh8IoYQj1emj1RqrZXM6R0jSSmXojA4YiyUWpbxTpTxnqH
QzbTS7HufMURMmXLPfyiqisQsdj3tp70p5ungiKAc/UqDO1jShyO7N1ZhOWOUglW8lIKNOitRMQ1
g8tqTNLR/vbgEk4wB+i3LUAXmcPrgId011gOr3xbbcD94g7hX76nXE0A30cWkvhc7J1Rw4hj1hb+
CyX6aCk979P457FLGFXH3MDS1AuyCpEu1pWVmyJrUF6sn4PFINRA9OXct1oxiDpOUvd9srTJ+vGd
MQlUghJnLKX27yv04HVEiJMzVADzxllFmvA9atJAkywicr4j6JKscHUtTmJama4YC3G9EuQDXT4V
IR+uc1pzHgTsW2NvrOycU+8d4UUJ+rOErKjIT7Y+A64vl4srZCyiDDPArjLhErqc8dLQ6mgdnuvx
RT5ewwBHHyoXLp2ujUomLMottZBFccHDzDEBGPUQ/Fv6mMtu877W6ZeEerCV6pQ0ejin6sx+xgdq
ScD+O/zR21OoxbQYsa8EjtmRUL7o704/KRBIbOyxDV2A29m7omam92K1fKhGoQhJB1o1NXJHJY0W
3AthGwi3yN3LjUUuccrkipTfO00tdrSXKLqEqPVyC1YrqUlVMb0DaX2wWC4uPqXVSv5rJRedjTbc
EPnn0lGnpzjmLj8U4LLuNkyVEm2ZYeoS2X+WmoWk8Z6OAZm5mcOSotslkU8gsajWe8mODDUKJMFD
lMb2wo54UIvpiplY1TYepBeyeHXvDHruGKBMBC3pXLismkgdgXViQVj6YpROlgh6yPiRHoKnx9IQ
ljzPIRn2rUGqtXY1EOWiY8DY7d2lPXNVknCWCMcBA10aeZkXOPNrhXldmxay3niqpNxh551slvrh
pg60gSP02qZNlqr7rHARjWAVHMY1kuwTypA5vdifJcT3CryMbHF4KlNtqing0slxauAkorERPCoC
hvCW8/DklzzNKvjIvOOo+05ZsW0gW/q+is+f/E0sknwBmCmsiojWRX8XO1l0PHnEGSOP24DiWs6g
gwdKE6UT0G55H/yBO+8bEg2YYKNnje+Kl52HfF9efy4SJhRXyOpAO3bsEpA3cdchjG0JKpJd1iz+
lqZU58OK9oG0A1HeqH5esm+aLH4jlb1rSSFCLrsbSc98OAqmoNTBX/SiG6FXoOnyNhvVpGGmQJ+X
IIdXXmSfG9VvsbxeEM/v+xtJNUzZcpmRabzg1gm9VlIFpRCVfAgtXUKw9D3Gbohbe2e072M6Sh6J
fjscJ7bYaRlK6jLUsOGYJ7UwRyARqc8tcucpm5wHSMXLGINOEqresNvkt2CLRoZsJkLP8fvQUWOU
/7Uvvyf4DpK+pDOk/ilcOIKkBEij7Kx5/EpEyNmx9WgyqEBRNe2/7fJiD1092KaY5SVvFllKHniR
Pm11TZQkyc4R7OjkHk93XfLr/bEj0Qa8FGSKgh8hWOxeGR93FPke4dTp7FmzNp2JKh4PgxAo3KEt
AsQgIb2k5r8Hv/F7n5H4gja8k6uWYEwrAPAw22SiTpT1NJY+Mns1W+9gU3RWHkSR0HMt3va9Q1Kr
zzbc5ObyTHMVrUW/v10uJbfQrIcoqmQZ7i05sjyreLz/N05J4GUkczotLYiiGUw9SQjMAbbvx20Q
H34vXU3cOnxLekUCImArnIfI/FQvgJqAPJm5gFiZayL8QVmNvzZmCVXq7jTMiYWM0IAEZ73zRVm0
sl1SS9BdeguRbURHYSkcVbIQDTnquSt2lWXFKtBuLNh0rvHwFTn5QShdAJWxLEg0Yff+9VYCA5n0
8CLMTQp4AmPs2m1ElpeGaCLj8q2WuEfcEz8xurRfMIdH7NpWcaSEslbCYwPG2JngwJFQ32ytFT49
8Z0PIbckIHUIlEP3rw3+PLCfQIG+WXSRHHkI4LIsTt10N0M9/Q5rSBabcPhVTDqn1j6rOko/Oedz
z0MLIIx+O2dnj0FXpguUwfaAOE1+A+IANPxUv4kagN60ocJADckI+UwTnnVenxsekr5ml9HOcQCj
g3ZiAaFEcKwDVMgRo3mqHTPPOiitJv8xJ2YM+aquMfyAidU+z045P2X/bDWVNgkjjVVXTxuf5Yl5
vUXGmgEe9x4qYKEEkv2pZgNWGVLcp1IhTw6oDjaqig5aVFPN+skNA44pWBDpn3a8zCvQsW49PSIM
XS5EgyQEq5hYx/hvY4vEzNG8ygp2PUrSQ5Huv2zoIRfc9+TgDaBS5CQaWviflwnyATyjMMKoyo+X
2lRSERIcLH9CjD2h8UBuL9r/fX3FSKQOUaZwokofytsXdO6actXkFLRURc2hfgKvYr1QCJ3H7Jgm
7QFt+1MAOvbmHApsdKD8izWFCi5f2TukPr20Xc2xQatnrMOilmzmN8+54AVTeK8JIFkEpCJ7S+2u
48lUC5c80Df+2yFhJcltSPSSITNWkQX2ENxabnPMlr6FM/f36RuNnG4+mCF7DNrTAOBqgLE8t73I
5BVRcOUhjdlcvwTsy34WDfM/xgC+d2ZU5ohSdZKPINZSYBSfaMvADTuo2WDHi4ZPY7Q080Xgvqga
VHg0pzcLD8jYmUGfqF/daHURZjmhWQLYCtLXOVWmQKgMnChPVpYNYiU87aFMbxrYZDY4wq4hKiBU
BzRKrC6yNKXgNoJJNeU284aWUlbmvue+IYGgoWrGz1CuqWdAuMKC6ZCBO6046yNn7iS7QCpoOnGw
BHhtVUdZAmzd6H5n5Uf/IAWD/1e33C+6K13kD/YPYdn7pKubG6BP6qqRz2/MXO+ZbU9SJr1VMxdq
r+ixedXCOKD9+uyWgGH5DTfYvz4sWN8gDvuApMRD7cvhsrWtT092pB8ukOMsmpAUIUxm+9RmbrF3
/8pKh8FSWPXMpAmB9zfQrbqT8nRFj/oNd4mGRMvlqVGea1rL1gTE+EIEQ5no+Kdd23uQSd72t5ye
SoWM3sJ2md7UarNqc6FkBRNKatmhhTUtteXOZjFJh48knB7xVPMJY7PrdemT3fTrX7xrako0KGLO
b8Q6vTlVE7SIOHSE4w/o/qiKIMxepCG8hBmF7iYpu5y4vlDklQfCcVcOzV9YmeIETOuNIZxf6VVc
4n3YquSnGd/411u2h/zHDU/j5M2hhSVWE/Y9Znea4YeqCHxOwwE+5YxbV87P2/0XvxIHdgy+Hx4r
WgPE57Em9T1JiLHWQNJylDYT4yi4cKYnG1e1STK6nHlxu18kAzUVVwyAYUF6M3oTzyWu62/m1JRD
i7jPnxkDyORXYHQVzOQf62aVEEhtQDfgh7tDRnV8hbd2DAW8CyGzPwTJ4SHHJ6hazw3/G4SOjHvu
0lCCrPkU116W1F/MxwGOPu5vwnU139fYszYqw6FhUrlP46ZPpe/HOQc4ZORUD/AZwwt/t4dTxQhx
afvTFJ+s4G/8OgWXRHGgPnePhfspN2AfRiNsm+Wo3geaEoixuwOdYk3dcD9WBeCPslNWh60q3oif
2Cz27oGtrDicvYeDxBkXrK7juNYJ7EOyfd5uPpJb8K2Vmk6aVeqXTnEP99yg7CR4JK6p+GN2s7u+
cOtl+R8IUWN0zfZfHI6dyV0U2Sosbwc4gsbdFYgW9tw393bvuxrzp1QeUXcF81j4SRh3LRMyQqAZ
Nxet6rhMKZLzIl1KrWsYAosX2DcFLH6nB85t76tOG9+YqEaBlghPVQjlsUGMCtEqlX78DUXbqzGd
0p/NbsTGmSb50iqEButwTiVztB4C7vPdSgdW3NQnEneZIKq0bpAGWJfOcLwgZ/x5zOscUQ26sAGD
SfsxMVRMsbmy78O75P6Q/Eu/YxhMFt/cdgH1pTa74KL6BjWVkt+rk+pvMOScoNaw1SOST+MePoYJ
asfCDjF87iOh1LCeOl90z9cfwEmApzAHTKSnLaWTV41dnstnGCFgPTDJT8gr8d6/x7/wxLIfpJRA
cHy91YZ7S1bFtd4MUNtrl5PD4PX7a5iH6TOOdEVX0ZFqtvbFvdRJPDCObLYuaGUjeAYjurxmhz2S
tcLVoXmmM4qEEK2U3pnuZ+sWsmDCapvBG9M6pOe8HLR47Y8TepRxTBLrmoq+kKC9bv+rieNsqYpW
BmvzUWBxkdgujEEJKh3YhroJuFzgitSjYgbU4GXtoo4ThtjtEPFd8VG6loo6/3uCa8w1KaGreKJQ
BRuwry1wtF0biMMJDGRPHadt7wF6wiNZt7HVq/0qg51At7nI3KT6p32CJGNGknBQvumXtdy7jB0/
Menfy6szqPF2tR0lNbj1b3XIxe9fDSW/QfXwtECHjA97e/Nh0sWZ/GE4VxcmuAIoHU950c0Tb3C/
xkip1e7OamhUAEgQ7t+036qqjfZjJKiAP2v7BUybI4UCfB20Qt5/YrD30sp/L9042Msju4YbJ8Tw
yBK6D1HlGa2iG4AWOTVUrCtktc1gFy9Amy9vXLsANN4t+4PO4akn7Y/WBoC4pnR1kgP0rJrtE//U
dBjtiNN6jCyBShjTD4T4nYJ12BAshlJli+mzlqL9sgHoOiDQOgWhcDcrZMILtm0lXzJyt+nnscC/
iSArgZBYlOeg8LbSy4kslLNqXwRkhRElWGaW6D4uVh7LhxlwLoqQzpNVgKB2lZWin4XkDrNbDNN1
Y6PRIqk5w1MMVYrgKf4Qy+XcvSam18RBc/qNjyDDO6aorIhIZefHbDJE1QBibPyMUw+7GICZ9FIO
fyfgChtV+KXbBBZATdK06NN9NLRlc5ewz6FoSwFtCpX5wT0lTTKFj3kMAPemln9XD8/73f0mIcIK
pBSBKta9oQChALoNtw7n3LYJ0j9bM9nZLB+Wu1F06Yn3kNJuzHNm1lZht41voGE6sezD6QrQw/e3
CGmSalwoluZEzcc4vCpug5grpKaKpZSk0/Hy2AyED1SukG6/ZTW7bYNY3GkvpMjaHVYzCtq+qOvk
ZN1riovqy3gfAdxhUEv5vmGbn/1Df/w+cZc1prxXknHYTb8dPoxyGRf3iZpF8yGv+PVfMs+w+W/s
IuSN28HpVsKjx+7LdHIk4sy4fz+onfWMKIqwcekbsVR+NWJaz6kV4EOJm0I0uGqxqFpxPOWG4dyi
tGF30803BVn0estTLubInsy0/bFh0H/McDkk4bxCxjnmjSSNb8RD45K1Gt02q69+AXqwqCMbfHIQ
yiJD7mTD5/zNS5pF4Xdnhz1HYS5+eKf5GCBFtIrqxhzI1y9jQyDSCAzgcsEPe603VlAZrriQXMVC
MgnXQJ0aFuJBrL1uiZVJKWnOroh2uWYn4WZ4bHJryRvgGxhmIaSsLJQW2pp+l++kG3fktW6ytflX
LH4gdKpFN8khW3k4TbeRFzIPUWvZofVT034G0hPl+TuUthfNUWrFjBGevDzgNlYCIMkzkndGT8H7
YEm/O7MQlanmxfR1GLhYE8+464fV7KHZ++xU4PTq2LL7JJs6he6f98JD4CIrjap0PQX+hYwWK92I
BcZ29Z5pRVXkeJyExTfeu+mRkHQqEQyuLm4JarpuWAoBIFVfZFJ8XidyhBGArQuopoDfLQfNobXF
PP4rB8UDxujZLX9987DjSuEHB+B6ZZqoaIm2niGqePef9j47wUwOYxTlbgTcdSl1p/p9wPpJHVQs
KXrKwvehUuV4RJiH3ZrlrL0JM7u53Lb4zoQnMYRictwS0+9Ty7gakbIm2+IOUM4ptmfenX/yvLTD
D9/06Q/nujWZHA==
`protect end_protected

