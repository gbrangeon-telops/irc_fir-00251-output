

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XHCjR0nUvMBgM1clzO9mSr8YEx9qhDtoXdaphp+J1JlsC9lSFtsV1/eTy/jaNsyBimTHmHB4CLra
VqfCr1I3uA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ebEJK3bmI2t+WsBGbhWIt2XB+F+QW56z7Xo7/vGiNjxPbaq48cjkY2KIIwhppzuYFDUdRDxp9Iva
RlWujqNPGUrxJ1F5Pa0zN6dEMkhKPrWWxZpAFto5e5cB6DM88tJus2O1hLy9PRfKWKn8u2fBqIhs
zvXwIEX3Rz7kU3GI+Wg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oZLpbXnbPC0EfiuqzOyPqmT4FdlvB20VtdO3P1fZux3uAWynrmGeEUk81RKG8dIjeHdSPnugG+6c
jKeGIJZZbH6MRScqnz2QBuupQkeYWE+dCLOq6/P5LV7F5481QZZ3bx28u0vHGlRYhLiMW8KnJ8Xs
JLZ2IP5YULE4cFTCCV3WAM+IdulnwSP3p8oyM0uQffeAJkOTKR9dl0lslKFBplzuTZ7EnXSmYYXA
x4iYEfwbmUZvdla6dJXCCjtKnKqL5vI4L1nHOaep2f0bW/K78py/TJVV+vsvE7+Fi81aNwDFBE3d
V+IzN5VNKD8wM+OpLL9AD+xsAbJ5JCLz2sqFWg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YaruXmtmo/2yQOaZLp6UQc/TTak5F2uchK3/c4SsORqNnQQMwFmjpORZM2++MrgqzkHH5KHH+0SE
PP+ha/JFKIuufLvaAIVDYgMKSDFaxIIvD/8aIAhw7TgTE10+TXTruuPFiw9U65VaBnD/nSEGkP+6
2M+aqBTG/2UNkEELi0I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SWJkuOmi8gVneMbAS0rfK4gI+24fr/0jQv+b5sUWbuvKyCco423EdTDwW7ROH+M/MaGP2QTzNz1B
sh1p0mypy290KKaGmvaZfJU7NOmSNGAsA7Eq3zQGPHDW45/4GXnri5xLLNnybO7r0Ndv34V/fxH0
f64f4NRroCys3EmRDJeCh0D+WDA98E/EHP+OtfmYOGeO+CDzxS2m3FIcGKs7pkeR5dgt+S6srqxz
96yb5/UwV2cpnC9ULYZHZVQa9WYc/XM+Dk71YUYpaEFd7osc9zT0azChQq+XAkJsqukhufRg3dQK
YVPZotO8blEly5GYlPFGnRW13eEh9DRYsb0pSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13296)
`protect data_block
2ih9LyCJuTDcDydOwf+bBp2Z1zutv8fZsViGQd5jI7OJeRrget0fZ50zyUyzyu6NH/oCn7Ub9GLK
sCOMmU8WuKaZgw0fTT8HuJ79wOEqVYw4II7WVIsT5kYN31BLffScyQBgF4BUGs4Q88sqoYpsvYaz
BFdfV5cn6YJkkZc8VK1t+tV4AGSr3KtuJYE8PrmkQlgVhexOlgiOgSbsDhiuEzWqZHaxuJ1eiHxa
4hlH3UhCO4N1y1e8JQvX3LjO0n9CmPO8QKC99vY/Wsr+l+a33wVOLlrb2GWJ+uXXGzBCc8VaxjD0
Z6dyyrjuBVUs4exRG3CNZ76QPZrdaRrqL3KITiZGNVqS7+YiVuJgcflG/1XOFnAJN6JmObORJE0I
GB6gqZaNg9xgtlX+yT79vrqfIEQPKmQeCewAZWFMNDYS/jfCCohz2yUq4cWnDlYOcZa/3j7p53b3
LchMzKFVO6CyWf0C+tU2+w2UU57ycIy+c3sGId/84Ee+cPQh3LunSlZwzzoBiS2qy3ZI/AWzwmcG
ntEGNbUvziZeQr50QNAeSS617nCC5oK4mPeUh9OmLmhW68XCyOMU3l35WSXeWN16q4wR4aW5wS3K
7H5u/J9ZJnTKmOMLD125StFxmQMFcC52guN8HvTTk0ncz0b0+fj1PmnE34a1o4Mp5RnGdPy0mBFW
ZveifLaBnkxcQICrPMyvfw5oh7GTVjHYJHW114FnBVZJCXGqBSWKClUURHyQt0QVGVLsXCkQ60LE
8LP0QIrbUFRZ0SveoQJ474FfBtJUThpYIbRU6LLIfpVv5nu5KYcwHBpWB/S9GoYYX4+ZZAilvNZn
vOhQ95uWG9KMWKj32jUzyl/SYjaSx6l5KqRek9LzIwDcFFXKMUvA1R8sgvUrV+wgBRUsA4tY1j0u
ctPxi3zm+FmVkUsl4BfpTIDnObTdjqB+nO0dCz4kVVMLSvVmsiqhaP5s4r/G3JZdbJ+VffpeTifd
XVc3PXTSOQZIEhMDebwtWBZR13DmgJ3CtdE/Zd82O8ReXrKtV+zjkEgiYVcZp76fi2T0eRSjeJWC
ywr7ETolhsiZE4kfUzVPfpPr/DbcbzzgupVtrJ/a1J+mcrynRxYX3Qy+/Q54gWf8q4HU8peOcRAE
XkxvXkgnw3stPSATgq0adC6qIXualdcOTozLiKgDsqJbFp5A9DoeAdBa2yHuQoNoXL3b/HKa7qsH
twJ2vU8Q4do6kyZosIdFyjzu5zKQWFu+DHRQtI8QE+ZqGAfaJ6YOaOIBtV8W1ew0GgqC/R+iIduB
CD9N21VIhyK5hW4I60LtwwGMNKfJysgwusk6FCCRz0M/UX48TzzuvjsY2X3WTxknXYtTOFL6mmM1
5p3RrU88gTnPN85Z1KWmXK3eX4cAuY7g65hmHTdhuxCfy9z+x6t7PlnE5/dAmskG0hZGKHixz/mh
aSbf6fqLZxgpIAdu6hWFnYT0VIG9N950AXFuPz0J18r0ecmS/zchnOrXKCkVzG8gZ/Ld0KrOJfQV
WeK3SBcx1HMySfMbbKp0U/pM8dx0qCjOY+ZFYL71eFp5fjokGgjjI24wXnnK1SM9Lk3zqbDykUdJ
8cVqyJ31V5w+05iFZNCzxhB7pOIHADZTlbZSq/eDznsHx09hUlCnIcJ9FLEMP+Z0AtqERBpCe/rS
/RsaCDquanM9iXOr6npgOh/1Eu3IjEvJtmEGmo2c2Sgn0v0bS3ak1ilcrpjoRUS747I9A5hzYuIT
ARU7/LorRa4HDbIN+Va8HdMOqfKPiYzL0UayR31tjY6z2AcVowztfAZo64GS1mqPLuAlS/r6Oh68
EQkAu9lAjlpAZKRGL4uQ3jhr6ghaXzwT1Gzuj3OPN8ux/nbvhYIXS6lQGtIEx9QSNzdqSQu2/GVH
Xfa9CQerEaPOQuzz0GOs9gStcRbXGoc8Bv6gNHXPpyW3YfN6TzWN3E/mHsjAWS+GB0TwxUXaSxrS
VuBNDoKKi+VJAWeZjI7JrzyBXuz7RWidh5YX1itlsfuyzgJD+NsCrNbMagX3Mp4L1EwQxNmEvi6d
qAGeQ8BdT2BWjLS4J7bJdkKhH2P2evlUr8M2+kEVkUWZHxGrsFS43aT9TeuBDmCxOXIwalvlNJiK
awPiU5AxU/n7HiIxMUh1eJPXVlaIjRTqRoO0WFKXjSr2MGySis6sZGTLVt/3qcALxmVndpTMI4/r
+GVHJ9lPsUiA7euw+OzmDxcWfN0vrHKibpXYTOhbpQrXR3X8UG3TD/Ew6rnTlAv/wU8PNCx79xgT
CJ74rAZ8JUUVp2HBxJrQ2FcCxUC/cs1nVVsdaUrpXz16Tf76MJpx5w3U/wyeFJfwIkmNYwYSU7Q8
01ixh9V8QtWVmAuot4upjqOHvj1tgNkHMGCQmrcox6iu2k7TWYCbNY3CiVRm2fn6k6AsSY6NSyV3
eqgdFv8lb9tYCXs9ACxd6nRwydqsr2MqkOaxDIeZvFcAXAxEBB9jkqKYsaU0QpMsm5tRYiIpzE5r
9qzJUsrSoyA82fiYnJC7LK8kJBgN8TcWzA1s+6+F4ryKGGVH+xysHcbXWNg/kUixowbSqdGwCgca
nmWl7g7Iie8qxNaL5O4Fp4DCFw77vtYPgcMccdE5N7FHDxMbBxAyihDjnhufVShgg0SxFsPvJSru
3QGkk75SdvyIxPDha+bDhV2j5UZ7coF/9m/ArHanfa1H1MiyJUE8yvVyDZ+lfsuZLH7GEVK6lZcv
UVA0ktrP6zFAOh5PrmCfCQVU/y93mKSrraiqduB5HVEiCS3tyVoSKRbIrjd1/KHajP3Vx+RI/Glm
YU+a2GygilNhtIXMWYwk49PDO3elO/rY+ICosiw0EHvzOW5rE+AODKEZWc4lJPP66LXnJ9o/pGKG
6uRdgivh50BU6H6s31tGhAVcVYB/BcjO86l7ElN5+KZKOESrOu+3hQ9kPlMEKuk/YRZi3eSggON2
SZbYr2XMifzbbjc9qXqdZtAbhou3UQ026HGZ2hCj57cWJeX2P50dIe5GE3yH6q6F2Aa7drDjGaQL
d+HscJKYCB305Dko/0jz9/Qs5OGi9xq0dkIPEvNjPM0s4yZ9gcELjg6h6WtEFNCzg5KTfijbuptd
nvoTCXOEST2dT0bpDgfnHuPp/PeDHV9n5vdJFYcawhDjf5wgtvduYV6PtLiovGLQcGkwS9bdJi7h
D1ZQbjj9Cv6JhMirg7xTY24AQZcvDs9mT8LgG4FbDkubtm8JCvvOqakbbzzYqUlf3Eik8VK/FUgj
cC9EFZa6340X6xwAt1k3MVk4hkxhwKCbcorkJGmG88dro8jl+AOByZAHRY6Oln1YTyemICOa233s
b5JH8GLGQbq+/jjhvMEbbsqzPtUOj+b7bFtfVUDrGxi8Y8fbO0KQj8LRFZEwW5gCxvbnnoVpOkoK
TAWOzeTT97Ocj3w06Lt/IxfN+1+/Nvc9G7kRp9AxFEW4cdIBC7NYenmT+jNwyMSxBTvgEbg9xJM0
EP6S2iTC9gZPF4sEcT4apPOw9ziSh8B/5YhN4A/RSUex8Awit0AdxbOdAMoXBnSY6wLIipxGyStf
qZOqnCUDV9XhBtliSNviF07W6o36fWfuUy5e+4zJKyFfpv8/fGoXQPINpoQaYdfmNRR7irBcPfyZ
ct3vVdg43ZsXqHtVJhyxlhEL8OmU/Qcr3oSOVT9kufChPeqdxDpWg1qbh22GEW5+TO7pDrsZBe5u
dxntFolcLT/wjU7suri50AUb8rn4qKzoi+MRIbN/vOF7CaYT14fzOB6/LPepcwCDtwBk9OE+/lzB
nll6lXRQycKnNAQ+8uNO52BHSWlgrFKwWaKsOs7v2HTd/UkVv20WFDJ492S7+QI8SUHYg0Z9u3kc
Gs4vjqc6TNOC0+rJQlciP/6hJV/1ErkOaL9YJIauirjY+KsfNwLBuSyoukDPJS0r9Bq5ty3+dxL1
/YGq7dcFTjTvzj11V/qjG+FsefWOj4hC+MlhuEZUQMfJySJ8jAINzb/FbzXEQu4YFxAMr3Qzi7aT
zj/IqlVasfT1Ql84wcWzcsNxKdmmzidOKvDZg/TsX6b4DTOVoBGJ8AHPDAwfZ5HhoBxp7K/J2h/v
SipM5rwHWB8vQQEJMFcZsACIYkPyTT+cTEDwOGLXZ71nY06dV8/DnrlEsQ+Jp7zoSXhLlgQhZovn
9xoxWR+5JpTCDW32ns3SWfvcO7UzZGrAPHTLGAKeLowvalAj48f1WPNXHVjPLOCPvoXthRjglNH/
Z6IbUTBfp7w8ioftK2Kk3TBdQS4cZhvNo6I/478zAwy46E67tFNGzd0qbvkNlzhkhe/FTelJ8IoJ
pdf7ZcVUUZzx5d/WATUN1ek3L0AE6FCQNMWmkgq/QSMJyy+dr4hth+Vp5cuSNjRFbRVFT8WQsH7P
b/3iXZ1uh+SPGxiSMlGjYIoVjXBfF+AQvSRfhN8cJCXPvcpp0Jkd/cdm7/VvhOXwkxcHKvQHy8Jf
WDg8Kchz9SOvxii7+zXwy5A/z9t/44WnV40jFJxtEdUlQlpbwm4aVecfp1PEMk2cuAd6wSG6bDwg
a8aO0S5+LxDP3GfMWlzYzsxjQKtI0WksASZniDcfOwNMWh5hRaBn2KRQMhvzXv1imKGqO95D+woY
YTwAkNpwFahhp1VmX2259LEit6bJ5Smk4d7DGo6dKpMA35sSEoxxK73Aa1m0OuVWQ/sPTl3BUIh2
GK2S76/0FBJ5x0HpbTwC38MtcYhBI2wiO0fqm0U+WG7cQ7jYw9s74+Z6b8tj2w7KP8zDLH6AuQeY
pDYLP3vvAhZGIb/oTO3DrdKWxrJ3WzftiJMvFbxyO5qGbzT4Wikcf2YaCPZSyMIzdLbVSWuOXzR0
Y5zIUfzqZwgzArydFkhQr01fbDkUORkCW8JIbr6Qk2vCNEwbxndYG2aT63KObcrp5AbMBYzBWu+O
DqoxnRXY/02DySsPJkwlRN2ZIgV4N8IF80b34M3SnKexzX/IBUmAHVkslF5dtO0CeoIjzPEQdNWi
rTSzh11l84veshqDGeJgoXy6dMU++Dstta40sLLkrGCvwd8TidoI2iew0/kKZITPdpF6b6rGD4IN
KDSH5rctX9SoOSYTsRYIoDjvFBoVpFJ5ycG5wXYrMYlu4DDzewcz6QE0tEcMdbeMpx73OI4boa9q
8YnSAef/48OeuGx/RXlpkMN2FHPmPt4JqMTxF8i5nLU3Oh0tjRHgWc6zX1EK/ElQBgVLQCkU7St6
ofmKgO2A3L3B69GOQeIKglJdItgN6vyOXGaV6LrVVIhKXboYWQ9AeVDb8LJfGi7MScz+kxPwcWzZ
O4VoGFxSN7Uyw94IQ4LrqHQjKgk54tonN/slAII4nkJFi+Hre5qlIxehtULviOpG+WNLxxHIr6+w
B5l7tNiDehyLzkjERAKT2ErjCthDqMp9puXrUUE821vagyDZXo6u1n3yMBACXQhJExffdK5qRKCT
XLLpDk2m4ZjQxm8AJxoCBK/KpceY5AdiPuUrGVxc6MLjtegY7MzCFj++0rJuYgTYsi1i9/wg1p4Z
KRpugAVOpUqKJ0e7P33B3lLgvr9LDtJAfIzIGIWtJlcQS6SFtXc4iM/yvz73BWW70mC23cHhbQfR
/QN5eOKGvrCG6u+mQlLzU4/eHiD8fobIa8h00331xbWQ4+Py0gaFHEYei1mgHBnlgMZMpOuzaKLb
YbIzDyKXJ/r5h3mID74BBeLG2/h024A1Eg9Pn2kFXXSZ0SwW82Y0XcdY7l7iI6vh8wPC+c7PKe46
rPeuFzYPNKWE7UcTgLycLkKYs5jMoRlo3XSy2F1lBuqIf4RSMTnpmIp9EPo54KKBexYCQ3xF5ka6
P8dEnPhOIIRHYNNf65IGLCbglYNMsJ2AoxxPXdG+9KY6Wt014ygmSjeP9OIpE1DVKN9Gx6TKHkQ8
s6EInN/PBbMMHlqQzfqBnZGCIxw/Cem23i6UtUU4fBKMAEFsZwgvDUlxLJgmoSrcZSSoPmpw+VqL
VKKA3NJpcHpJ2e5NacHhmf7ulYWfTK0BViPzUWvtrGIUdfTXsxnoZ72j4bVwOEKCO8Si2FRkQZo7
FVEttiYK1YriIk1o3ghduLdsB4k0W7E5XY6m/FM16setzORd1zp933J7j0hslJ36smoZYL4jolvl
Gef1UO6QlwRjY8nKMzYEvaIboMcK5+Y7Hka/a5QejpQBJQTneTuGzedFwripJ1aNtDingTYkAf0a
+FJwjjaC1mpiyR/2DtidVjWQBnQvRplSj8ysKo6uADvAtaNXouvUYTTcKY4/lAlnQ5t/xwBPbcQG
fXmgo+Mz8mbokwQG8WbkL/JI2O1cSfWRUWxHqH2kvVf067l7FPzdhXo3Dl1yPcfl7TihBcgwTP1U
8yR5hkPKMshhRq89jgoc9uCX2739uuhg+0twkMzm7xb0c7dzY8jul0pHIhH6tKHQoeFTHm8Bi4m4
ooHKBXR4x6K+y3+Yud0K29T2h5ed9NJK0eCTObtjdB75YrDdZofcjUm/P+cL964h4acZe5iPD77k
3k7v/wdlllUyo5IrzS1o53b9Cb587q4XqtUgLEBd9CZl+On6W46s3kYy90kVd5W5tU+uOZfWHABa
dfo54LxesxHFwB/eQPQ0eirC7SF0PGP9Kshlp+g07vyoQgkvMaq0DkPoutp9Xnn8L2IWp1+JIWoi
VWOjEvV6orO2S0Sm0UMfYkfskMSTP8t75Ce3DcTGDOLT8MxcPmewXsJKe1mvF9YajxhsFYOLMWXG
RA1SZsuzLvtwY9FS1Cr1WV3yPxfKeMPXqNEpbKTEXVUDDO+rTN+kLVHTU0cD0YDiDidGLrcxUkxk
Vjr3JtwiNwbudrd2wQ8nLidXaFYQ9YxiYk/yo9UQx8GAxtKIaRpuf7W/cNKXQPn+ACN2ooS08ZCR
LyCjECFtlAmbDxTdg9D9LzePHYAEbc14e+aD1vVkkgRf987IfaEmsmtsJxTrjzuNezY8YjgPVBCn
nBcvNcUOEO36od+9dcl3LUZG2MWCNjyQpLnoPdTHKHtD7XPu2xJKem1eUQyTKJDDRbMElqED5WuV
TworPdQtq8rkFj6au4RvcHutZC2fhY08rW4bqmVXwJZTkPPMUS+NrmQICukDk7hj+Dzy3OauSV3K
AFEbtVYKCvGkTAnGkpJ2ZtDyafod4OcYBccjJSEyKCk/YByzvakH7HvZut5+uejCFDHLmy8w0LFi
ShZmL8tBhhTZYxYBBpiRK4ZC4piXXbU3zCYeGJlKtPsUfT7Ts/701VGzAvWRas/lXUGofaDSk5RA
3CCAzKKEOe6JYaZPL/IkmIeayktM7uKJ34ZyJKYPg5K0+MYu5ZgsYRAfGRBaFZPlbDlZalf0Tjfs
m2RfPqY50peqYHy3obFqUkstSKpsEUdg3rGA1RrQ2jZX02jMozNrFvEDxrHUNhYLJn/pHv6TkkT7
362RHQa65owrINvtjXOs+CkB19O5ojXmLON72ipY179848EqTldt8//n6kM0V9G3BjuRAJTaWmY4
LY1ahWlo5lUhdIqcbzcG+OkoQLedvhgDHTl23Cf29QS46bPCOp+QHMPBc/bnyFl/1R4hYwJ6B2vl
VgmNt5q1YCPDIkCWMq1fRFpZNTRBmHypXSc57rPT+Bom5z6b4MSWwvJTBi4PhUoomZzYuSIzCevV
yoj+FzHVdfMNxxm2+GXpjE9EJMNLD2Ei0ihQKsP2sidS8OCcK8KOnzRQxNS51j3016ZInfclVQxk
q4X216Hd5h4zl5eh3E3zQbF3ZnVRY9lApT6umI2pgGzUeGOKEQ5reMw+mbJqZFNY8DaSyx5JMq4O
4G5yAU/Oirb9JjYpKdYqWKQ826yqMqMZEtwGelx8Fk22uq3fPda0kRYv/eLXJASpjdHexFwuCRbf
V+CLJaCabrXX4fsJMSlVJ/pcDixwKdKqG2XWEa7VoVj/Ej/NBCdKaytP3sFGKfO2jKqdVcXcLQ32
R1I6eT3w1LMikwEk6EsRrajOCeMbFjkMRdfC7HwrIe1+zo7w/NSDKgCE8TqEaEbfLj9oebqyygHx
GPn6138+B37FqQbHrP+uBTFruD1iKpLjQc/7aUY+GVZLfz852KESaDLR9kukFQa/AZeXxRfDz224
OxCvgEH+WQqOvRw/TKcTnXBdeGy/b3KqOem/KhsGj827ub+Cuor/wnQgr7piAtxtE3lAjB7X/9qw
GUjNSll/o/G18wr9bLdk0QJtWSbUs+X+Pfi+P/hmfd0wSh6FnJCY+VF613JWu7GaySDKU+bd+R7T
A1dqOB4YNNiCVqEDTxTEHIE+qg1B+ZuzHjX4Xk0WEvZIX7CHCL3IbjUo6i1eAAsROoTOTYKTQuvb
hQdPxZXMDGY/t8Mk4UKsWdhVNCOGF/pm6nhUZE8IF0dSapEWJ8Eu3TOfRomluNrHXvY19j5DACpH
n5DEEEf/KxmWcg6IMnb1SeNVJwLKBK877DDONDKhHXz5jUZ17+AeL3hItplcoJ9GEXRkQCTC9u6E
YvJPfl4HpoojlMP7z9CshmCZmnpffbKoZsnOutxcbQUv7Pvkbm8Uo1lFfCbXfuSGTQb2680OudY2
0xPmf/dJevte161OrVedUDXXyUnCOkWqV4Tnn69DIRJ1wGjoDkaxWC2lZSm3fzy9iXQTzWQTff2h
rdGkWQHuzAu76y6wp2/iQqy4pSnYduMnyit6j1WPVCwTDcO6nFQX91xuqEWKdaPgc8P0xy+dDOrW
Qqr4Szl2VVihEMOS+oKajhV58H7Lh00ubfRLnhCUOtindN1aemq344YGSchIc0WLX9wBpg0TC7o9
afsRHXXHCh+dmKOLFxVKlrlyjkv14AtrAhfJqQJo7LBLbf6cSS4jvVfr0Fmi9d5H8ycY+JChdWCG
DuDD02UTiCndprjMaN12xXfqF8EO43STZ4ciqKuStYvdl2THH/Xze1771zWxJvXkmdadi1s3H6ZI
eKVTGYSJrRuNJeoArI9WCY/X4Qn5GMQnk8YmgS/ikXWni4wKyzzxgU2n48e2jQHPiTUd9NS7ejZd
1YqiKyh15KSmzRh45/XFJMOnHvVCN75p8tKw783jPsac2Lgi2a/avfe9YNjBKWg7ImajDmT/celd
N+gnovDrh7sJ0rzd+qbMmIDqBONAkmUAv1AW9YxSjwddBIxgr0i7KZ0RiRn7Nhekrl3rmf/dVfes
a/rh7MkPBtETe0tz/1/EUzSKDWfU0fM7X9DhLiJlXU/VJy3vTwYXdr4knc0MSl9FmUtfJ5f2yjkz
9zrYsiAusbdbrFAf+FuiZwX1WvlzhzoXYnySzEhzx4GCJc1OwodoAo0lbJosfooQn9xoRQVhfiV3
lgayiyMtMAkIxmBdKH9S9DXaJ7AFjVC3302Ae2Qa9QTTrYtetB94+YEJDOXNv9dl+HSx6P49hvr1
/xg0LsuNRNUvvb13JE0jFZALtjt0p84mFGN+TOq/fE3BmVCejjUB1RT8JE0un/v7yowRG+oYPjR1
cwP9Q7+Wfcv0vjl1CMKkVnhtjTHVxJ/UgE7akv67L9EmTHuHRC8PnS6PJ+alZ/2/10IhBbwPDCUg
pb86JssWhmipwWuELxTNS95YTTF3eSfvgBCbRmFThUNa8Oo3+lO4uqxjCjT+xwVAP/7alzfIzqQC
CpBXtzNI1KzibrihfWwD5yI5fcOszFUfncahqWkeanMlZDc14wNWcBlxogF5rhBzHhRv9trs7+rN
hdEvhCgUSroOXSZqEKNzx/VyASag2xaN4++0kpEYREy98I0GiLXjxpCo/gSGXXgc+PeHbe783wnG
XlF6sOPS0ZD5BCkf4KZrYJqt+BRUDgqvuasUwCKyDDAcgBQYUI6t9LK+hRmp7ct/VACrSulqNWvS
4IqIsLPNui+t9jR1HPhuJQzxPFP5XZsGRpCw9yy+/UpVKrqtkOOx6LGJQ3WSVQ7cTXJtPWFTxE6u
jNO9Ig3yBklRKnhUFD2PDdOryR+WaEgFpoVeimgzz0a78mqKraAEL8hDwz0zUM0ggQb8yKgcVXbY
42sB2GTX1ZXLsxuXDEKxi1a4P5gcH8gTjZoTkMLaQ2JWksCzHlhI5h0Dm9k6tqza6LiSmOJjYOVC
ejFMd6KglYZYQn5oGHkxwz1FAWDYlEY8Ny2pmcCKbDdJ3hb7380ATYDx91Eiy0X7e3qHvxgNDQDS
uOfz3X7LBaEFfI3bRrgIOXRLjsh5hYn5M46r3MSkdltOSdMNrzKT21ZGpWG303d3xetxT/WlFQT6
x8Pn3+oS+mB6vIypcVI6irpRxqB6N3u5+DhXdnfz0mFASNSnRkrWjfBbyOWIvEQFYI2mPpiQkmI1
uC7qKDFISZvO0BiRN6ODHw1rondzdWCk88RZ40F1nLkFbvG6vhKEYHcG7Kjk52OmxXrpwwewzIBB
paegL92X9TxWtir0A+ImjJIccZkfbuTvVkinW7Vxa4C4wMUCfuyzh/fiM4IfmALs0B2nFRYJJM+m
2sILlQOMt93+2q6QVHydZ4WdcH96y6e/c2/FZTXgVoSY0x/bvSjZBiAoRpqEnXuSkhLut94XgYQx
1W7KoRJiqMMDXefs3lyw4To2AYmFfhaS9/EIjwoeYGPtXkcAHQLLLlXmv9Scfceg3QRD+P6yjfC5
iVRy/XIpsA1baNB80gI+ynd9m6UhZZkkA3tJEAOMjruaqSTbWu0GGFmrkR/itovpnzpdVu+LHOo3
WlCCx/fyofuLtLjYt+KvJFs7JJVVTMCYu6SFxGhT+cvUyJ5lFy5Eq3vgoBxCMJdvsIh+yvxvbLfI
hRurkQ07gyEsjDuYM1LG9/+/Mt3brZ5b9VFtE649uDw6YmURs1wLyxv71IaAIi3y6FB6vBfSOagM
EqkzcKAwpiSVp7QNqKKAQIKPqVwU2Ibw1gyHvlRnYdLJgoh1CRLu2cIVHiF28qOYLCJTpEyugjGa
gmSOo14FU29PE4dFBNZQXRkvXJGZWNdXXhs0SUhFL35rdo7K+pimb5IUb1LEeYTu1JoIDGHPZOw2
mGSrd4u05+//I03feIXxY+NlCXgG6dMUbJ2sOjHv7YnZ6EQpywHGLRpqu8i3uud74Xc8YL6LJZ7r
iLITnbNSNPpnSI7eIWAbPa7jyGLTVFjYdVDhIHp1q+T3sjHOn4k3nt5+MfCaGlHSK/G1VKR0Frkp
uWyM9sVDsOh/KD+bY3IaR70jjfgAY4SuDBJEGK68Ss7OJhniaWDM0/e/YBEPKqPCHDEcRaldvXwU
8IYT6clArXmppKmS05rMzPknpkfN22rLKEb23gWPpmW6L8HlIdRuxtjOkiZwKiWyNvWL8FNsusa7
IgPCEfJXFks1ftv4ENzF5hffc4sZnbDxKoSd5PWaHkf0N7BNpE2SEJ8Kjcf/Mh/3BM9AzTPHAHKV
/GJt8RJhjV4wnEbvPWigXR5Lf3SbkHafKbz+A1mKbuKYg9M2ifoYqcT8tbVBWWu+2QAfmR/PYQaO
HpDNjXp+b/G9Jmsht4rsy+6luhiiSemQX2lhKWQqkMuvsYJkGecO/DxmonU5n8kt5ovUnJuCxUtq
xvF5piIlsyajKxUKyyg4WVDO98N8BhYUwfb1JQQpaEDp1WuRqD0tt7C3ly9rBJvFZrd3xwlqmiWH
Xd2YBxLEgxXcobVTmKMeZjOTOfnElZ3WSVTtDRxHH2iPBxQo/2X5zYjYuPQ6CZ+5VtwdaSqK+NdH
LHWn0rrN5qJ2tKYsP8+BdY1tnZbU5RurkMdZEA2THzwgEMmufC3D0UwcU8ZKSau5q7NSuMwCuuob
X0KRbIzk58xZJpElbcXs0L+cCNJzgRD6WHLxHhDXR7QovlR6Q+VObzvfFa8H4YbH7Xuz2fqEtkU+
wOQlNif5facUaOjvL/4OrREa1X1lmjadjNH37a30T4ryKPhfxgYtdfqo8N8U0O4gHqu6Tm0tUkW8
ma5JkFolPY8lKtx/oFBbE+LW/gzlpf9AAyaLF8Q5pA9Igt2QA/z1RUjOSJRgQ+yyNRzL/E9xiyWD
NzCfVb7GbDfsXMOo4ZfMN29Unzdp/UOlUa6Q9B4HdwCFePJLLMGyk2A3AJUwaDUNhI5WUlrRuMcS
W7QtIpjK0Xg1s0+vnOw7R9VFq2TCFvUzTztE3+C7S/R7URwsLjKLLy8gqXhik+fEvR1M01ZiuUgw
JSaoUpfvsOpxsMgesVbf8uz61EHjKPepBmSgGCI7ZM8Ny3oxzq8rRBn/JN7V/TPUu5FxOSooqGBm
Dm6nt7RZlFbQsmIF4B+B+cP+Zogoru5gF+hLCPVZ+5XsI2S8wFWi3vfgOf+YLdrD59IXh5bsfT3R
NHAJnWZlnY4VTqdhaPUKFf9f2IpN8uxlQTV6QiXOUFP00vlJGUCfknp41s1DDx5kg+4TsdRqMF/S
YKUN35FOeJLg8bBKZPuzibis08cCfWBZIuJHjrY67cWq4jEAs0PMc9MDfS4F3k4mSRjTmHk6P/SQ
nVxqI3TheOK3DxvMzhkK9vhbFDAsJVM4J3DJiIZ5ZXk6cVy18JgSc/phEkkSHLIX//5r5kl/4xDk
G44HuAVz1VBt48YlKKNDRSZU4k9j60W7rvse6nFOgrSM3Iy//Xsfv/2WmmxuQq66dmRqULKW80xY
Rjf7XDMOkRIkXpOlt3Hs1SGMgfW0JavlgAH0pbGTOQZgMrcCWdrudd8K0x70TmQTsLwUVb5C5b22
dElbH4SwjVGLkkP1HWOUDYXG3zFSFvZMBWAodkbH1W/QouQs4ParNyHamQBTjqNRoQ65dbo7sjm6
R7gMIw3wEeDtK1clAO2GsmKGZIujjaklCSWbXBgTYf7p38Yr0sohveznWKmxA4g5b4Q6EPdI4qY9
Kf8q42azbJTvtZ9/Sa7O34CeIjX/BQiz2qBvXEO3cwIpna1NMcW+LUMeZHw5tGeKGeWJX0TEulm0
IospykceTcUPn+DIvpFhQn9uyCzunyby1NqVWqv/i4DoBrL1dGiDIP5d1dU7+8aOAF4tAeExmNHg
z0z/GCEKxvgIwAl581vRin6OBVCV7n56fzvfdBfA2Eh0cF6MQK6z04IPQVY2lIVaD7kpA16zXhqW
7xSSlDwwSt6ATLi2zhbzsqC9lDAkqTNiOcmXaUpB3n/hXrJVGdZrPsAKHYfMe1bm8C6F5GV88cVR
XwdJY4UySG4l011i1JGxNWDdUI+Ytzbd+lL5OpvvpvJQoy0B9EhkxuFX7efDkbRqYtx9Dcu9ogxz
qb6Y0TOwtCyqogwWWjdc7xNdHoUFixtNE5elJ1b7/HzXGUZSUPx8/h91UclpZ28vvGYsqCT6nA0F
BXaGXq0hO/l/WecpKTYCSqvgOzF01DZ78jq6rf3W1ESIeRPeLp4rEOs7Axh2hc4CFLj5f8csFtcL
mKrOZnRpDXWxVpokeVJKVN6MKnMDoTc+gGzE0xde02Zd+LEL+QbK92TMimIlaZ5iE2fAe1Jknn7h
6QHaySFGCdUfbNYAHgR/Lra5PQuLY1tVyxME25lTnB1aWIwmqVKqom5O8nPNTMtbhundmxEAerA7
A1MYjMgXdtj4g4wWwuwmkMjPymXFbgH3U2fXtqXdtcIFKEYcvZibwhumynHzauycuuxxcZS6Gm8u
eknQtt9ZxO6zbmBVGh0tWb25BCFxJTJjele7sqBCJRGN7HzLf84/fjAHWPqlELoty17tjGWMXH/h
r90mxldNzV2KSzQK3OmFZSBSLRo3qVftvr+hJTVXKHd+JhZYV4yx4XHSPJwA6bj39HWU81GBvHZs
rRIbttK+kn3EIWDIqvRdpcDsTSTC6ifCBV2VGllQdkOC0UPwhaZ1J0ZDa7Mx74oJDHz2Vf30AeiN
WRHdWJHfg7xlPBS7+KTwm5mf6KlRkY+xY4Jtn771BeFjn7puxxQB+IqyzL9OBybzXAzgWcIsQmJc
y+jjZkHa6T15vNfcCdTOzlcFkdthabvC55wFiVoraKDdhpQaiM7bcMb6ZmRz/x/DCGjkCzVEqA/B
9c+HkWX6rnpYZ4GSmWv+7cmOCv/VfMpfLojc3B+MhdKe+CSwc3sBWFTnMx/s5yplmgyepnroQAga
ZU0LHNR0fTRgB23wAIwXr1eAjEMLg6voJFqop4quzV5FKWflJPKNslaV75wr/3OvaD96ZyPiq8sw
Bid4VBpDFR/k117NI5/uFTHFXbGiCU3hcOj658/1/DpfYflFbQjL///D8gjRh9G4Fsfs0TpwBpRy
hkCcw+pq+8uTCpLXC0P59tyKsgd/qLkgSvLAqNLPWqW1jcyZsaep6MYNgEVKzNVoGMH3qe7/dizp
xBlndOBiEqn4VWelvsiW7gMrq2OR79SSBY+n+qU3OnLnFXqVy4Z+qTZmXhZOTovlu4lKPuoiqBWv
+SVRMOPaxEox2YCzayT6xD3vJdNxLRkQzO5EpDAC9wYYQ+npV0LUf3liSiNWUmWugvfk6ZuE66yG
wOVbnL2/iVKk7T5vXYWospqjR0j0CeS77yoPFdF//HtkR+KUf+v/iImK7pKbkcU5gp4TWNvAcudc
mFKTxqjCWuTN8EO3Nn7KTPIf2W/ppNP3bIznLZf5vzkx+Hm4WNJdkX3068+r2s2rLO2FklTDgkJt
Cma2tWXRyPaPSKFSxqdsg1Q6ra2cSXWeiHU2jAbAEJP+eh5xovtSbTkVeQLnYikBEyvKV8X1jZ40
lRD+V04Doa+mf1WMY7csThIEdjDpStwBhnzoMBGSxA9GjhsmC4CyQco7DwUh0g1e+1G13irQ9x9o
sNkH5cSW8J/tNAvXaqXiamKJLuz8UUPcWkJIL3XHt6mXArOkItKxN0BikEBYSl+lf0DqP1+rjA2j
wFr9O8VtKaPWYft0YPeoxPY5NSbmxYb2dvvFbRpqIRaty3VuoS87foz2a46Dox41Yhxg41EMIcb0
qDK5892eIJTXUquf87OphJtdyWMIF43qVdoTIrEfMuRPw6IZi2o1SRn3bRioK8o9vSn/OFPi8CeF
2ljrtzDnwHEYrDOB6y+4KBd7XEVgggv5tpnUpbxw2gJtGzv/r4SIe2iuWJBy4oRA8cUjE0+3LwkW
YFre2CsCyfGTkmJspRc+bhJBUU9nO5Ym3U1+dqJeFW2Q4Lb68nnAEGdPxOASKXQPpR7lS+D9HXhP
92stuau0yeP73PTDwNlnzNwiT7qMEW2/df0B71pFgaYgS1dKWs6OsDfvWUdNnva2cN6EGPVwo31d
hf+vWXJwyl6gBuw1rL3wVt4VK95TWC7blIzfHXVSInXXTMzD23dV4iHIxbIavbyT3My0+3TVFMZN
QQJJwg5j8EWI+myj/fAier/1Ft5HE7UBvo0/A6wICcb7ZGwt2HdnxGqcG0AcafEZ4f5kGgk746mO
zL8YOdcjuIuMBOmovHA/wKtghJ79k/Q3rggT/C8Z1vkUHFggRv19mHgyCaZfHuemiFzesk47jafM
MQEWynBAsp1lkNIwTcWyqMxEjhL8HQn0WbCvdNPN51onIIxBubmIDj645PDmO86izUpZ3CyCbTan
Ntg6sK2Zcowp+ScAvC78hOeKVGHbDtWXMj99SUQTG8iH2fwHJ8mSi0kSyIY6zJT7vDalIDrcQymb
D/Me/eKBpLj6J3X1BGJs7V74vBHSXE+cAfglJBOikZsXHu233f5FsW/q684TBzkaOQIicp/20fA9
eda5Sg+9I6BXIPBT2zZTnCKfNCSGB4ROZxkCMyj9idY2m6UUAjyyD356zAxgXRe3Mm4fRb/assr8
hEdGcHXLnyrq1gSm6GMRpATjT6smxHfX6MJeqlL/WNKyDxrresb91LI5iYUVFycTFAO1T440rtxm
l+AKAad8FrRjYdlGkh0rdcEs4MBFAIOAbjH3WGJ9sAeyWGvEVkpEVUFVn2JSub4sZXroyaRbgEE0
P1oWP+e0DljEupSWpOz7rnK6VilfV4R0gf3pho9KdlXe4QAJonv1VmQujg1/jrlSMQTS3O/C16wZ
G0YOP74lDiled6S7R6FP34EaDPFU2NlvoEX8GxuT0Nn18vUSqs8z4fMYMXAX81O1xfBiXPLT5b+A
RMEr3utD4rRr+EDCvkeM6+aOpf6DBKSYaYDAGD6vtTEDcO0ArJwvZ7oFUyckxaQ8T9yiLk2DrbTT
CFBxa+hjFF3IRyOXBxNewyV5KzYNRkcZ0MYFBGPcI6NeorzlqxbsS/ghQjVqhE02bpXYSgIoGo9q
FVmtDZt0x3632JBMD94Dj70A4QepSuvdLGh2+e0DPttGYdYyaGTi2XUU7Ef6iWfSPQ+J8lJO05UD
iiSIiqmxZLKt1EJDk8TNqBaTNFN+pN8CydWVUelSq7bNpIgCvA27LuQ4QF6M07MbuXq5J/TXQrpw
x8g3w8fh+39gGyoz3xSjmXOzcIN4FBCYHHderxeLdQ7q23is6zWS//2SFEzKoyCHrQNAwHdxI+Am
2jbaGlr82cN9BFZVx53zmIPpH9ooI5sAOvVdUngonHcpn7o6eCGXb8H/p/KooUUIqiWz1IFT6TuE
bcnG05XPJNM11exVT/7wrPeRlzWxhIFKCc+BfAtTieqIm227y1q+V6BlaL5/q8n3aYCeKFrkoUZd
zCCNMgS0+Y2d/snqyGW6buQjLn9TrK8ni7dCyc30jEnRolMCRPnvhkYDzFZmbFpwDkgvaoU2MpuJ
qCuzJY3V6GPb5XYatkPoD/apFDxiP6jXHdQCLIzojdBOXJzAmUegXWnfC0ICHQ0D2CHpWdkJPWZ8
CUpwiZ4TNAJURbNm8ZWJMqRXoGVq1Q7cKfzz1HbSXJ917ilyRmn/rXC5jhsxZXGP/6bxjL5XDqdf
zFNbpilI6cbTWy1DXhD8aKLZxJmMNMGjD4PzN/U+9JnzuD0zoCwyWjJd0aRC20YhEtEMxEhbzSn1
TVtKEUcvQcVamyWUmFYbMIh1hWdYLhwkvaROmx0RGRdulphjScC4VkiOxX40XO1domC2qykbS2Zn
YKnBmOok/04ctwDiCFGvfZAOu+D1zKkNIt7DA/lPHqPp5SSBJRJAzYDf/WSChBr4/ZyWbWn/LSmo
C682xugE3CkT1jM1NR3r2RJAmx++EYQI02x2BocHV2Wsa8K0cbQ4QIO58uHCAW+tk2b3mGhjeSfF
Fq6QPwxfmzOmT21cExjAqHeSpAIlHJydF25d2FkgjgjOt/QmWSrQUPRcWvSol2SoKloEVX3djrA7
HCmDibT2Aw/ReWWONDIgEdVrTk9G2S+3cQG/o1XZUVhSEQmuO/cmbo8dxwrYlkEmOmpDo+E+a5nF
OW9xCoHE5PgbL9h+JzqFd0RG8+6t33YCqaHEyAAXorgeAUmh0cazuujQz6upflSGFHbei8eKL7rJ
eKzf4L7j+kSg+WG8YGM2xrqPoRF1QhWC07QjPQq6DUrbxUP7hV0DALI11zyRVhmNCsFKR4+tCsBA
hFtCLkwlCDkJ9hpEpS+urEkJkvG+/N1rvz2oblyRMbOP5Sm9DPX3FQd6jGKAYjz0MftfGhXTfHj9
tiTS8QOPC5JHhHIqX2kYQjTt9tfVpqPH7ArIlL892zM3lYMtdcsU83oiS97trkI9LugVFddblP/t
5hEdInW5TchjaHXJL1OOUAxzKCrbLfAuXzSpLhXpBlceP33nKYHn483zee9f5lMMst9puLFtqW3k
5DAwFYW+UUS9GDKYpPltmlgQ0xhZ9wzMEsKL9IOuUfiOdGObRK+Sh6TB6dyZme11SQhbUxEXSF83
UuIiJFXpsoTmzlyk+VJI
`protect end_protected

