

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FAkw7gRmEwDx0cT0lLfFXgH94E+u7pXWs5ahSt/pzljIAtlVd5PhOu9ztNGUELVfoO4Gol+zPLUh
TN9yRctY4Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OsI56UKE4Z4O4++RpLw+Gr7y1Sd3eUkdDGmGZYBu0aWjoj+iDwzKGBcBG0rF5D+4LwCAgnpAGiys
xLyYTz/ObATK7L0zNe+Mx/H+/j5j5SXpNvpcXkGCWx3Mtg6EpqxneRyrD34svh6fn9QBg9AkFvdb
eTcam3dZU+Gacfm2Ivg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qc1VB803xD7sVBXVT5KuCy+daGAjeSNtMgViDKH2bpJoW4aexvjdVOFa9Cn3ZQUudsfzbRtbOfND
3qwRkfwGKGa/rWJp/b4u168LG7R497q3mKgxz4wZrw5VVWth06zATVCPkvVwwcP1aVCYV0wxe3+F
BcZo/LoE5dzRftELWM1hbxUlZMlSl/apI9c5DLD1ZPtssPXqyfH8yGBCJ6IwpqThHkCcKlxPWOFY
XBErOYYrcO+fou4DBovYWIgQB0ZKOhCR4cvN3q6rg5XOYT99xP70Y8jdZqXKRq3PuDDZEya4uwav
9zgp9xA7sRjUN5/fcIvFMcfDutvNPIc7IvkzWQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xeydwtnivo2IBZhciZFfy3r1qoKk43zuwlyfDAWr7E6QmSwqVQF5VHmc7oNu8/L6oqsi8CW2guof
n3LQZ6J8fPLN7CBNStOEImWoOU09vnECk8Bwe5gJEo2CSwnqojJJlM/jtH5jKtWnMb5YecjpsAkT
3bnS2U0oIgAvNLFItdk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QglgmN/aSMz0M17AlWb9oRKStkdBh5nVOwe4/WnjlbCHuTNXWcMIzqLlv5JcAmIdzL/13EAMS4W+
LbXaFXFMcWHAzC/5AZxX+CZbwE46qfB6uGUmUBTFEckk+Ba1aO38uKX6EDual9TqDkiz6OPrjmC5
MifvdDzh7mlaB+rYqb5sjxUWUfJCpXIOgO6lavL3535AS2e2hAYpmi1PB/ejGTuva2r1NRmDkiUk
Uq0oiyBI4sQwmU7gFF9pADJRyzpgRQuSICfI5NAGRTR3by64/5TeOArBdjuY9arezL4gMGXoOIu4
E5vrAQOLZikLF7X3/wpaihrUarYdJnuPPVXNaA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48992)
`protect data_block
+oCoghsass9p8lV/xmMPo6MtSWghX/Pgwt4FRg6ieJERLkBIgwGyaRSZ/Kz+1Bnq2WFvPcCahvfs
e15JqNIsBtRSfT/DTknmyWik1xiB/D2/BPXS9XLqQS8aIqGfk8W4CmaVMyEP5pSf55NGKbOv/cn3
av+UmOpHN6DbdqJkU55n+GOrZxxQIICF36M0aiFUqlAU2QnD8QDebNnjJOMW0Fx+Gga3Opi9aON7
JOHeYJsCPSbts5TYPAk6C8SIGWWENpTl3+RQMwPlqHtS+F7HDG2UxkowvNerinobxHsvRGb9/UaO
/aTJ+3/ZHPEWferHZasypJj992/7Q5AU7JPlnsUYOcvE7DTAOWIlmKqFuaie03DSqyMvUgZFcrv7
XsI0K5w9HBkZpjX/rRrpty8xYXXATwtGGeQ4PLRSot1nQjJDylkukIDulOidDhFL7wRSuduC/H32
lMpE9bHIptO1LiQhDRleRZHZSI8urKZsXg74+C/d7fzCDT6gTfho/j/fO3qI+MXy1ILxk/UH1ncc
VaDsQox/mNrJncGyMhFbg/11GgvM2O9JC+fMeBcDhjyXBGlaiS6yvfkW2ATICEUcugcBbuoSD3sF
rM65HNyiIYssoWXeNZ8/vMEz1zFMC+uQ8z5W1fKD800CNqXPa/CuZJAztD7SGW0eas7hEwRTniB4
lj32qGCjy9f7pwrxMhiR/5+mWUmQca2ZhBIWzWHdZ/DfW2bfNZrL/xGaGecV5NgOEqFZ7meA8q+0
d98lFKJjBeQw0VhMnJPqt+jzgAEAXHb1BF0TQ/244WaD8iWBBDcQN9dvDS73kR+CiZ0Dyh1jPdj8
pRewdkePS/tSEq8xxnNMlyDwi7BpCO5xH2zPYWaeroM9lImweyuDWGdxqdC8ejk3gHMuirpek1re
mYW3jqKati3w9HEi9rbgHVr7/NjEFDClLXnDi1WSpVZIeIe/xNYjO/+2we8hIwoRI9z4cGch4uLH
og3qAlduc8sbXc6qk68M2aJECX1yUGTI/yOBhQlI4W48KL2Uv0j3Otjy4dG8stfzfQagr+BtKKcD
uWvaDlkQ3MvtkU9AcwiFVSZtFO/I9O1W9uak3LOv5G8UrZm8UPfra5l8cf6YmR+dZtHyX6f3TicW
1rGkND4aXF7dZ4Juq9dY5N1gn1gZvwslWf87Qsj1P3sLp2ObzUD4KbsDmhQEJgBvBifcqj1MReFa
GWTgp3ADhT/zi3fJZmGvqtOcRWyPujQwWbIDRD8YlucnToQTR00UV+m2M3nN6qEnN+NKn55KHLAR
a+opGAl06hKOWJrm45mb91B+3IUO5B96F/gp/Zxjb5gXjluOy61ucPrBpMCRVA4kZIUoJgfiWNsj
G8P4TifXn3lGN2W2Sgp+lx0aXeWzeCe2fbyDgoUirCJUdv/lCrEFgR5R9mH+wa+medOM2jFtiGP+
SVDxTHZXgKgCxMOgQYb7wddBscWhM+SsW5o50r86pbeS+gY+41IgW3AW4VrEN9O6gIFBQOYLZiVj
HPtB4dKw3wHy0Cu5aJSW7cna/d73WGSxfty9k4YIgVkBCbpl23Lcu4xLgBxQURj35oxZvGHOKGPj
/zF3iXZHgyPHxnDinQkoG12vSIWhN8fT3NCsLbywfOxq2lFMldaEksn2knc0FoM7bjZaLgfIJUyU
6DXR3i/A2LCVOqW6zo3EDEbJEVZusYfY9YDbEK8sZ7KqHvHQvERzxhG0zBF8pU1mOkpbMdOc31Lj
qb43UuDKh1Ml0VQpwqLL95uRTePZf2q61LKjR4j+1zYXOwuI/jA2v3/IrKKO+TKeAJGE3KqlbjXB
3GRzaDpo7EnKtx/AUNB5FEucG2N7qyNSqiAVHaPQ6nyBI7IfoAj7hQJBfUy0yQ/FLYgfc7jgAo3J
hWNI3Xl/LGf8CV2PhZ/SEWhXexCvoYXK1oySXAMHJ/D2w5Vw69dgDyNf0Vb3Y6EJkHgUcpKTjqAm
2P617iYZCjdtvI3XT2bH/gtjmHbA95ORyennGsfltjGxUWojJ+9rZcMYEyPWGeuxGDtezQhzEKdt
HYoJynKiZ6Ya9niGRVYsjDX6i+aK3Bx+eCgAbWhA/AEOedGkLCJJHnCnaMyCmwv8B1Gqp1gx2ean
lvyGbbHJD99RSQyvX1sG3QPYNg5weNzPN2/sg+4QODoai7wU3KgHwdjKMnKYcGKA539cFTLR4B5k
sHyi4YMyzjKmuWBYiIkf8UJofLicwRBy/pFn8RUdoDTrxx8SFShw7j6DKotVuyuTqm3EdtcQMtLo
E1FdZ5pW9v/zKSXgOQqlSxKCX4lZ90HvXvsx4ggqgqVpKVk0+50RPqfeF3h0vFlVA0c8W9r1HHlA
buFx6dJn3oCWMfiF2uW18b5br1AQSKwlDhoIVzsySJ2bhO905+jVhNmkddmAnwQXfo1rtTDs3VGX
Jkz8pa0cC5VKjuWIwDe747++BC9IKFjMLugqmLe450lhow29cDrrMZ40hCqBrnDHeCy3l0634b4V
JxtVlp18bEpkj1YiyXZe+vjOR5n+2WCu1sGMS4OqpfDxednBFPyd0G/LmHSzmb58iep16fgIFzNW
A4cpH+qowUkezxE0YES1dD7tG19tL/bqn82PweyVK5GOH/eoTNP3u2OupPyZbgPpzoDHMdYsLT+t
xsuHTlIVfyinJw9Ky00LcBrnkEVBrz0oyMj5BbByDBmPY9IEoaupxLwThTyCgibPBQ4iCGlHXn/H
j/318/Zr6WbGXxtjQE9hwNfAeKSgZk3X1fX3N591mzqCojFVQe0hc7XVTB4880RVfUft8XYyvBRM
VhyOsx02CGhT3RinB0vYKuRuo/8Oz3z0+1Oll1q0ofGucjYOjL/dLTWCdF2y4Y6YNpryhG783Spw
2lVevld/+TCNmZjiAwbtyZSFQgsWAPc274m18HMFpQzfujbJEpti1qXvUGvp/idHSiAY1LvzBGir
ozM/CeVl9TvPp93Hvr/TJ/xvRJYkbB8jFl9xM8n6MryYqFXb9oP3iYHmP6I7bdGuryUiGhQeSHT6
Xm+sLWAyxx9JR9lBlQIrptqM3bb1zzTrwsH58F0/Ck9/q94Y7axV/OWLUrHgtmpXjVTSNrlBEAxT
UzabC7+N2o3Ktmd6Fx89Pa6a3Vt2ZFUpN5ppMFhy346NyNRsowbzLUsYOPrO/Ivm49rsP0/UtlMc
89TdFdzgkNv3B8VL9Sf30BffYRHlxW15Klaeb1UUajHU4/cg/m1IjTBWul6Ecx4qnCOwEdgbvti4
crOtrgDz0TgwnLuRvrZCahqc4tfwqN+29TXK6wkxhV7qKtbMyJXshndxOE96HwEBwC7tpKYiCd/2
YYessZVr4B6GvWzD4UW4D9mdtTtoBE15a8L5j3yZhDGqqRmiX9EFHgf3rgi9a16ObnLdC8y0M3as
fNVczVKzRHgQc7LcNUIjcMCq2wJD6rQlT9TjtMzl6GdjlUdOe6pjW0OdgD+bL0YZrHFp5/Awyg5H
VA51G3/LBi2PygADMYJcblWMLasXr5UT/gpPN+mOE0f4EY3+q4hi4YwJM7SVnhfHudb7XM7IkNmi
j0bM1RU3ktDXanKwM+QKTSwZDTfiEY5DjItkRxPBmz0pnOKjpMcqOAqpM02i8JNMtf3C/p5aV+Dx
yLSPAUxCC+b1GN45o7ZxOJZEpEaaSrWgr1YAnIwqjKny+g8/Nq+O/ULiAuUQgcqEU/0gwG/j+19x
83NrDEIYE6EEym7AODIAs/ErQX978LTZ0MfQBW98FZPONL9Es5C69QC1pcG3o61tajUoxx7fRWv8
+sL7criZfBw3keKTtRNX9IPe7poFyv7a/8eTt9Qys7W9y7GOBINMqAGAdiZ9o/wB9EepiuIb9scF
RxolHsJX/RASjFIHLHO7HqYkjJmrPROtI4peNi2qOW8wDE/9QXRPeUYw9vzUdY+aG1U/3sRn4qmS
GpOQlCm/LrfVE0PAoxa4cRd8eEWuWYM7jhiGXSwV4KvL/bo5Bv8HHxbqKGhmOxduUN5eEMZeW05i
wvFQyZnbfKx9+gVzuSM1SOoq5JIwr38oAJMKf7VoX3FfjeLJFbTODb1FjhPzyNALhQE5wZlnM8T2
NEdIjVqaIHYMzfP4dQ9VGX3TQRWrP6xCqBbYSjOFHg5Dbak6QPkt9V0sdt42tEJXYBuB7KQl/in9
BBgkrCcNA0Dv9rW8bofL6r14LE2VYJ97Kl1R0xXvorsBLlyjCIF8yY8ak/OxQBJKRyFFvYWloa7d
6IOUV0QYCVlr2GiYIk5xRtaH1jq5abDcCevZuQzNBHrcmQSeRlZO3mqoIV6rX4TyFbsVMwSdp53V
rf+9qYEcrXrLt7jKpVU+t1aC9UeVceThiVfIf4sjCvGz1KXacG+7ufLFG1NOW3Xc9IzysHk5eDYI
8LjRSDgEzYwnU7fJkY7EBQjFeT0kHZ+pr7sIdLjl7x2YQCyAgZNiJV+LmoZZvpz8+Px/2N66+g/7
ADUfpyiHR0EnOLEmDgxVsUxRWFtgFWYrQ8GaDF/iEyMx+SeWtbEIhuQTA8sorTplHYnS++vOTUJL
K4q4u0HB8ihxki/B2lFRxHHM7sZ4bWbTZBzXeprGMTiYRftvUzUPcAulC7el7BlPGR+T3FoulACP
/IiaCt3uGAAKSbW1TBb8IdcDWzHWLB0Flh6ZpMbNdrSG/ogd0tE+UvjPXjQ2uQ1oakvMWVWcmepS
bvYbX0Os+dI4ynyYx9fvuCKMrPX0U8vZuZ39MWYgEhpT1WjJU+0lN8qxUsaqs2SL2wvBWB95lqL/
y18zSsENAILV8CA+RvgWSK0eUGZCQw5rpacLgi/h0lOseDKRve3QL8QzeeUqxIeUgdZW9ZASfiik
2F2FwKUuZ24a2MEE4GEyIaAiv8/jkPMFlOMzqOSGfN3WuzwIE5EJ/XrC8ED/Sr8W0yNZxpAvKj0S
wMF7/2hSM0P9Etqd/zEOUikAiF88LYnSVGTFSLhUVg1keEuNJHiOCQcLV6hFo14KctGKx9Dge43V
726kYXiQ9vdN44omMhynQrQDnrragEdEpgwtPcaPaDGhliET5YcMkbiN/6KIXfV4VTyLiFyd1Yer
dJFy4RRhw/DbQBdj+gE3EOrxKkPNl+DDsZuKfKM1OPNvbSEDyaB/yyf1qAqbzl/OfCMHw1RDEuSw
M+JMjPRzMugda7a757K3m8n9K+zZROQqVdljjS30S3+KImF7phTHPDD+Dr5rsGSEd2Ac3BWIAwS/
hnIvrifk8OxAZtC4ymrtBT9OuOK8hz+IMP/CF2jwhxMd/+VcSnsh4lXG73nO5zrdMJ2ObY3JGFDf
71M0wP57MZ78/QAb0C/kb2KmnlmFy8KSrdAytAnShhqU2LiwFffUd9WsRtwG5W+1iOuCgNpkcqVr
e8hhyDhLIj8EXaONbL7uUFzsjygo3ZGiCmGS3p+Ac148k2fUgDMHnTnvM+MsO2fzA3nAa9aj1YM0
aPYUV02NBD6wNmBG2qSkOXBb7xKHy6IxxwBjo3Gz4Zwwd1kQ4ab2oEkUISPt3Ahsq1ye59o9Vrou
8thBIpWxtuS60157iBhT+nbEWO2fQFwqF8mLlOblCEKO4Dl2cb7mkeaGMzuaPhQIvBsL3+1t+XYX
+68DTI20Gj7T+e4HySuhPo5L4H45LR3n0MZJvA2E0x+3wRtBR9xt2TNgn4ciFJFHejh6AezY1D5A
Uk+I+UNIOkYqeEp7tOtGdG7M07QssQHXRIDTuhmRAPcbkAkNSqa9o/znbcGIpkggBnLQNxCvNJhx
Gms+cmZar2r8VePe3lS+GD0UDYlY6Ehh+ufsJjm4F9t8nRgR5FVRHWd6md727InJXZKKsaAJSZiT
QCxJBF/Hi3hJH9xYpw7NF4RyMFQRMK74zlsVB4k/eGG0tqwGCaABALgsllXvDCKIKIFjlTS2KDFy
t7uYuf7gVtHJoFLOxo7ooXSW8GWunQb9pKyl92Z/TlqNQwrB3UtqjmtYI0gjgTW9mvfNQnWB1DEU
ISAwwI/8GeHxkci+ZtN/U2HSSwFvvOvPHeMiOiSjpzgqYcvwTlBxCEPBctlxiJBuHfW566ej612X
a81WfmrLvVPenQakoOk/KpCg/fJM1pyUXN2nB1KaL2DbB0akppGoeumdkvdmaD1T0i7h+wDLwdvH
vDdOXOxzE7DeS+qlO6M4qmyRfeUTgo4YlSL6Ka81c7MiqzIOUChO2rlB7jN7yMgdAp6iMooz2BJr
NS1b9Nol7O+bYUPQzOyyvmG2tUIAknG/xmuUDb3iZvRrBKsFi1KUnl8dtH4g+aTDjTM6GFWivXSH
N7/kxakdm2VStKKkGMSP8VSdBsk7FvmYImV036wAaoxBSPPoh2CYKsi08pCZxCVjuSCKv8SBvQY5
1LMNxB7g/dcHCUyff70xQhUqTr1QRbBOlq8F2vxGfjgihGjOl1DH+pewmNYPftmPkHLj8Fm6rahx
aOSM1kgv1vyCaNQ+kM16/C/ASgMHpCeci/1XZ3dVuluB4EzOU2kptxY7hBoeF4F/5km98Ooznu+S
ndAhnfOR02A49cwxLOLZh2adW8+1NYoGD+ujGJgh9WN544odzjhL7rwl2CMEwlGwngXUHzZo190H
NXtucAbpDHB4nukXD6qYeI3jiS/QH3pcvlsaPXDU/gHcOIJ1+Eziwubg4KxCeRbsW+Qtf4NxUGqN
ZYTj4ZNwbKvhMc2tju0oGYc5UTCyxm/JzU5ZmUhII+Eqk28gZOCqC22pr4Bt/3w0PnPNnFqb1R57
qU6FfTbDEYQ8eb6GtBczSy6gTSHlSTBD/UydfDK6VKQIx/678YawBEHDFo7t2b9jNJ3dRBNyA5p8
nAJlnlXpLVtE2zT1qQos5ZhuDKniZo6PSQcIZ7t4XC89OGGei8JpodEIfO/HKZelsEzZMQu8mD1R
VQhiRVBX9JxJC6BFGk+QMhf/5GvTP93O9Cxiih8IsOd17XK1spiusvPccvFLYXwIcezFmGKGQNak
8K0lJte32RnwE3P97LT7iPidBeTwgBC1dhSdlm8ITQwPRNvjbT0v05b9CwfwALpFl4fbZCvOe+en
ZLoLoo9IBkRn/Ram0J6IhoQr4ZAk/e6ol2mvV1Tj3ZJvmg5HJfh3crPzhrd5493UIraDw1bVvZhO
SBFWLuJ3XYc7vcdQLDmd+CKEM97hXAxE7d3ioutd88icCQlxpOBBiyZ3k9u3YZaBFFdLm0UvsC15
TUNeG9BDXpBfS1t8KtpTI0wDdTXqa3Hy29vk5c+A2FXLqwHZpyKqzQSuGXz0sSSpr28fhoIyl8Oo
m65uEcOqQZKZS9WfBuJ1KbCR11eZp92uojJnaQS0U2IhcIicIkqsik48MuFoVo+n7ofPYTypv73x
Nq11KuvUYc5PAggauj6qhn6hQyCJT7DuMFxxVtmdJGJss9Wgi2GuQioCpxhTQ3voQygvgzOZOsc4
/WRUdmldXpbLxipsP7eCpQ9TcqecGUUVddg49mknBmMNmBPcoNlQBdAS5Q5fsYjEUlnWI4TUaGyW
216jTM2XSRcBi0QbRqDp5cKqkAbbwZI6VqaryRg7ykAGg3DRNk3pTeBeQN4JOFddZlvnYxK5Tne8
6SixeBeCo06hmzACdl/smW22Xit+Tbl6O5JChDISmmZcnj8olsV9yMWoFyy/MUWWagKH0pMj3M7s
EWqbyKy/nYbor6681MoJKQXwzo/e9duwNJsd8dDAg4DL00xiB2SBGiUIzv1rvyjEOOZr7OgqxXL+
kA+QYqNVhdMjthva6LwI6SWSltnE2NpYERF6Yp4QNW6L1U+PWA2WrR6ush1Ywiq52AxAHhqMEOzq
qu8VWpl+0Fm+w+65Eu2jlLJVadUEimIFmgmAzcn7fl5cq0L2ISUZS9C5CVhPsUz9cA7u4MEJdpUE
H/YUCNgaYGWDP6Rs0Qv/tkGwQaoctKeqkHptX8piPB8MUgGhSTdOcgZZzTjKIVD0Ykz+hAehwPSC
qi+r9xyJaBWIvDJpGhkDsKlaR33hrTuvNekruDi++TS5cKq9WZOXQd+Zm3ew/AcOy0nmTjQhEN49
3cISVAKodyOK+a0yvNFJytwqKy5mSU8YOujWRXf15ElgxBiTgcpX31FlyCvxQgP7u9Uu73kXSIw9
PH643hAx4sM6FnMUOUtEKq+J1a6wHaT3+0zJ8VB1iScPS74+bwp6RLzIbMIEtYWRXVVZMAYLAjlI
Ruh2DRtVPAEyfoOckpQM2rAKv/9MBeCI9sh7kuR0KvjLiGkI0y651bpdGcmB+PI6uBYHl/Un5Rio
PClVSkf00edqg1Ez87cf9LKnt1KSjmNion4g+A8UbgacXIx+PWETrLQy2DqHG5fiC7q5Rfb1FTx3
P9EtE5r2h8OHtvd9l2z9K/ou+V01VQxg9z8LCzf6hPWBwWKCV3sSiH3lS6a/PgZEa9aSv6RLO+dT
SNBorwbUL3D/3X7npYGtBBirL6LDVEfhYgf4fcJs0clSPOro1J4hqqVn9hiUJGy1v7YfSQLXx726
9AHUhbnr3oGMhOstItCk3CX5Fl0LMYgkfB7UafWfXV5hPQxhpyGyWiBiUCX+HNTRTNJCW/u65DAL
x8kGtS1BeLsN0gUAnj5PBb7EVppYgWETEhAKiGwIidyuxbkN429LotGN6yh7Fb/s2ft9ngonSnjB
arvoBbXjI4a5DdFxGpYZS8vOw8PSrOuOsLb5dNbHPnycgwgghDGrgO5SHqToxMGlDDA5Goo4w/yO
PLJcL8MSs3DCxqJapUzJCdH0kRVldHy3V5eMfqY6Jsi8YJrw4SsMwN4C52X2htQZ6rWbTQcjyHIU
fts80mmPDhBDMsGTnc/k22fKfppkdHW7O5fv4n9vTt5pFIuWhqjRGBUPu6F3ie8o8Vg1jDlFmHVF
iHOXYeiY9e0xeEQU0PYgue/eK5bQmjQlnukiZsjQ/hKQgHPJMILDtrXes0YcOK//WT0FxNQkVQYQ
coehIKnBaEMHVHA3/oooY6B39a2E2blhBuACryJE25PvfR9g+7Pb7SmYp3zbFM46w6XFyuowsSsd
GDOUNhLZzpJz0E6lQfoLu9Iukks4KuNimC0jV9owonAQSM3F8JhGnt8NBEQAbT20dLx2CUxHoY1N
PSwBndwoHUAHVrE5f2ag2kAMIHziZ9DO79r6I155Oew6B4q0x4RVFqFx8IGV4q6gRdgAGaB/7vkL
wOVFFi0r+jy0tDWSXulNXPgZfxGR7EiexjYO/T0Vpmx07olttnxfrRa6J9iWqM9SIgOxutmu8eyf
/2BN+2z839Z67M0Q+AdMALgfm7XLqm0aCesJfFCTD+bZJKlx0JJ4s4KurUoJH01jMNiRcTJ0LxWq
Q2yH8A+gYjAd+tVsg042aGhKTMq75HAC42cCcJQJ3d+hoRzWZC4DWQ1tu7Eai3/5bLWZvPCNe+bv
EcJY1SjUyne501OhuXIIQdByljQZ5b9SWFx8SU+EA9kbQDcv/hEY/aHrTStXnkwv9o8jEkyJHTXf
MAnLaOenP3TYck7/V+ZaGPhXcklCSh8BhxXs6l+ysLM2qHmvjiRIz4PkYXewpVx4G1zUGgTd1qlX
qwoxlgweUoxAV7A3M40V8ch4K02n7PYoiJNYZUsjugn0CIa386hO7X7dEMMShaibrvfg+Lv3aG0e
tXUTDx+U/30OklYe3sL820I4Fpcmi2Ki4d8k13mykWQ7o6tTG19WCHWS5Y6qepKxo44MOkHYrqVz
zaKLy2gTR2h5gTlwoAwnWvB0bBh/6fNhhSkGFKTiO10nC+uFe+jHjtn77v/V2jhLC1J9ggV4R8QR
JbCDOl0AukPLFzF3HDuV35tY5t5jhb0uK83tbFPs408g0BDqUnzBjuKKzSXXYGW0uhWwRi76i8YF
zLc+STZuCYEwPzGUjcgO3Nrpct/zDtkupTYyAGBt4l+AwYTxYo82w2cYK7AGXA6x34drlix9iS1z
uV4UpZHaJnwX8JfotvRGGAKaApwdNsUu2YbAo53z0Nj2+qHBtw3Q5dMBfPLCkc83cPAIhzgT+Gf2
DKlB7lG9LqDu9Dn69ffb2tL6eABwqsHiPwnY5CYJQ3LH7rJSsK4xz5LQ0hFVnxxHPM/cbglxwQSN
zeJVtteVbruDmv9Qfxp+y9Dd/7XrKaIgN71BF//0eJH01lTVGKC/SItZgyqvrDdOsWnuIFIGfrvo
8FdVDI35X0URmaTeAYJjRK8AflKaJoybH90eSmoOAu29XvOPd1LTi9rk7dZRGZ5OYRkzzMxtzuca
NdUIe9iaVoD+KQQH+DjM/ZFa93SF2Da/TyLs4PVKd4nG/o7twSXt5McT5qB9fuVpU3I3Aujg88+O
15vhkILwex8ao/CzRLYc1qRIy/GvV/ZBmQtFsu21GNcgEtVzN0apAcnWOmjxEzraTgLM7cj1b4sY
LxbaVFL68h53kjjqkX/qMb3l+KUmGKRK7I9M3h2yYOISHgiBHffGsZB4JrYe4wN0nR0HS2O66+H/
U4lot21aU6umfRBlRrvFVi16lOm+VCc+Zj2sh9zIM1L9GuicNgb/nTPRfv6UnqNIm2BiWhOxHyyh
inQMrMfebUUigoC5vOzohWfpGUqAh+rNQHxKGc8vIzybHJs0/A5w90Ks9yXz6J27NiVVIED7Rr2Y
obICfBSLXvjqJOdezhncZYrRoTSz9uEZ4XUBLQetU04UWxI6MTu9fn7HC7ziiDQEtLXpC4oKknIa
BSCKQb/BiXaUdS9VXGQf75+FVYrowhODozzABZ383llpiRpm4yAlWQEO2pa2rzECYolzHYiKc9Pg
MUAAGrbLYtm/OqMwbmdW9mO94dLyM29dlz6o75vBy3KqhXgtMZwmm+ZZESpDpDGleBO/X17QnRWf
lzoMNGXRmUbkSpV+SUBbKXitxL5zFUYyJsdgHQ6PBOqz1RLbW5EicnAVTmzrPtxKo30I/hqRp0r6
Au2owc4xKP9PIjxitInCLoNru8tKOyqVTgXUwR7V7Sjs8tQ7+P3Zb5Lw2uSCoBIbbNN65nOUMewh
p6onX0rXEJC5mW0h6i3UDHVPVGQ1QcyMFZK1vw6yf8B8SW3TISM2h1DaSO5vcnmYKpgSeUfSff5/
uPdAFDmOLaDBSUuIFv5FAK9Y5ZL83ytyp5JFD7H0+tRnB0QkkOoZ0Ly4b66BBjlZVkQuHr70arDi
ZWmj4R/kXqiLN+5l4T85u3adDHYGBFX5x+n+FinMRnLX9QuRv19mzyr95JDuBpOFLfGIDI+lrl3Z
6xVH5kTikeuref5XiKIbHvEIApPH71DnUn3AshY/l27qTHFjQfBgc3ViEb+967FT+ZAswpfUnWIb
d177qM2naBsKMw9g/S3g9CF+HEeJu6EDw0Np4+mBf66Rx9JRLhJuVR17WqjCEkQYZ8H+gxC6QGly
Y4C1NPnoNVc/RWfsMXhFA/dkD4QtV0tmLGpCA+fsDDqSQUpx82k/c7rkSn13KpporXhUu77qR8ya
lML3QUcAm6b8os2aSG1cg5NdhIF5ja+fpKEIPU95pZLIwQ5xpbtjZfbXc6hSV+Wv7S1Zw1PQ3SRx
QPcRNzwt5V1nJDkqaqUwz9SrPmzlilmAZHxDzOxAx+Zcddw0LcdZKTwyPZP49jRre8bKkRRgCpma
8+ZmJFSyjNh00+HqCxDP5h+kdmUpcNUR04d4G3jzBttgLy6ZJcIjkgE3NUv4+FLQYjKgiFtFjDk2
ntZb7Oy4+3m1kPgcK1I1e0YQ4ZPEm5opsZcIoArp2FQqEvVVto0q4tBidTOL94zWa/AnR05vr54G
OWyxaCwc2A0acsFmPHG0zb5xrWoEf/WU69uP307nqSVRUxmTT/taceZQmSGuTRps+6MnY2uigTVX
Azdxj0clsz8J4DR4sVYch+VycdfgS/yZ46Ra1+fiTGv5UjWdxhgjIaXpck1/EFtIOVtMlgHYefT2
F2eoUADw6wRxGnqKivBLZf/RxtgtrtKYgzK0kcuOwHyY2diE07sd0wCoduscoFsDTBxRvHfz5P71
1K/WMOjSqLnfYVLqnq2UlnckT43P3YMgK++/7lP882kJ1RDqPQPnUml7cZcST04bF/v80MpTB1d+
JhGvj5Fxb5GPsvgbfgCVQegqfUN3Y+P4IUnwcfQkiC6Cdc6d8V2JAT+ZvldlFiy3l/uiILmh8EjO
r53hWoIU3x1uDDy37A3jYAGktnFsgrcDQ/GZIROPlq7XsIO0RU7OitFDRwh8mpAa2YQWKkqvjXMd
KvGFahTaJPNOXlKyrMjeXy9GI6S09ddkaAMF0Z2FP+iH5Vg+1jVhekaUxOmMybzwcp1CTAMiAOuQ
RaHff7lhUGbeclQqYuUmlXyNGXlNy51uG7iurRyKkZosZZoq/2QatOTvArGkaoW+EjMjCpu4gaE1
MHPy6KNtncEBff7ZmIekFs7ATW4/zrKrwBTcPncuq40sFo7YOP12bdw613N2/HPRIJJQ1rt1VTI7
2Bmhm3R4TVmApnNy+tX0x9aNIruUWEUqWzEmR3jkY9JbeqDDy/QijBByry2qhyKkEXwz/elj97Ly
fPShQtv3nBL8baSt1Ah3SA2UrIBSHFIpE6N5bEnz0QpEOvHw7sYCMC7kiVAXImqDb2YO/5FO3LBN
95D8uzN485M5j5DKSWFZWcFgBZiHFaclXZa/izp4gfbQ78I75c91IOf6Czq/9wtnJkOd6Jc+zYpi
86kfN5tf/h7HgM7RJY3CppU9PhQa4jJNFVeSxaPlVU47K3Bv87Orno3m6VfslL4svoAOvFhagSAU
yxjibaeLtfkDLm1hFZ/Y9ifVqEYeKZe/sWsxnkxb2DYw4rwNwRxgvgcEvMsHxBKDvko654ZTfFyX
Cye9Wu1C0wRVxRhZImD3UgPIEb4YYsMDwwcs0ZbEOftcPWpMjnphJLJjau/uzBaF7CPP5QkzjejL
fete2PAcYuFeQL05hivbdXijOmSvnvGTwYqozYk2NAwIa0MCljEHzMNTY4UVgUOdAQLly6OE6+et
bNBMeujOP6DxIwm6skjLqc65c3h6Px9dCNDpKJso/NFNOYDTUJsIwiiUi7PxTRS7b//reJZUwdO+
4LLJdZn3XvsmgUDKhPLHLJtH/hQxwd9h+rp2bc+cKESBIbO1bljbL6OItb6LzvS0CIY8tE+7S0ub
yJ6yMQ2lwPetlRwAqt/669tzVOr7EuN4/h6k0xHEtmJQAH+ZleFi2LrMbAhzVkU4H5zO2FRWSVYY
q6EsH8WjPYV7JnEY9kN+hI7MeCuN57uHiFg/FzjnuBKRfWIvDyxmV003aTHfSmDHlzrFCcgoKmdx
u+nMuLapy5W4WRS68k4PDFxC7oet9fFsrmgbTM7HPxPVa/zYhlaEB5iUHfTNl/ABtXKkChU7JjQq
mJ1RrmRwXrj70Jw00vTbLlNzrLVvNiR9pglDV0FMy5Au7R4fc6LzkVyRHUSB28eF8yKwoLnRKlwL
FcMDzH6wFj7JEnFMU6BNXanMSLNeIpShrT0Az8VWwpYXJsbEQ33HcaIaFLMqnNNgCv13KER/3Uyl
K6dJCyfk7CDnEavLYEPVMzDls5w8OodSBlZf72kD9APu75N4QGJL5S3AccSr7Lv9JbdbMBCtvAPA
d1RLalZ+TcfXg6GnQ1p1Xyno5mz5aKr0dVhQ7faD4zPjKtxDbg6munarVY6ULzqD2CWBFra5l54t
MSUBxJ/9gzkaZyQWaudngYM4Lsq6/8A2ZbD8A49LT30bhwrkNE4ikSNptwZmN4pP8Vj8nwVoP+U4
Sw9EzytWdBZqmnxxs2PsdeLTR5VvEBdLSBSw59SqwMx2/p+yDsQj4YJc5RGMNGEusktmwtLe4V0E
nyqN3SKV9V97g6NK75MzWli6nafLt+rtqWECkFMvTI6R3yGgQhUc9I/4u1bAjxvb9Q8o1ZPkRrsd
C95OpTI26WL62foraI0TiSpXNT47Ff9SYlmn163EIbIuG5orvkRHxWu6dS00UuF1JjbzJFRYLwGn
UVpQrJyw43rl2Z6ZJYTCV0x7dUGsd+m4tlC8K0OJgsCmyPFJrxhwRFZTzbYzBzDvy1RlwbCO1wK6
Z8Zy2+3FP3EjDoVQOj7yOPDVZr82JBII+e2LkvpfqTs/qhTLwHUJCDYUSq0y+nV2UUcrqctxwgES
56AjBmkPvusrHmYecoc42o1eMMrFu/hRN+yFQUl9TvfeKK97f3Eeg8eM4DmIDrQkMdV+68cimfcd
aGdPQ14Elp4Oq6DkreuxcQZE0Q36NsfdLa03s+2f0tLeyIB7gNOBVDqZWbc37TpRiF/Cxe3ml+wA
Ca0P1YD2x2f93Eng5n6veAmpnU8Gm3yBTny+Pv8tBY3hm7nSXXSNNX7+ONZKuVlkX23R4d63wN4U
ypXZffhl0Luu/yJz3ZQ+/DyRfY3X00qgxK/4FYE7AcpiB1U05XUXKWgf9MZTKuCddQyq6FEvA5MM
NPRSrOC905VbDIxGNXV1TohqOuLWXZHXdwKxYtqIFJ1g1EW11ZeLksHmL43/8JUfmpO9PZVfRCEJ
df9LQN+O+Jj4nMeLXdqK+f4LtljWosLNl04DMCkGYb50pAsYIc3xxGlburTuHfk1acahas8WoUKJ
3LDybJls+cH9LJ3lqO54FCH10K3rut8SQNrcHKKeMJPFZGsJk+ahHyJDHfOJsdwLpxg1JeOwIf4c
EgYyBh3u4AMBWwzaL/XcAONiXWr9ifQL3alY+JssG4iBRy8+y4hQf68OxaRZfjee9Na4+ArE2Pm1
T1eM6NYbQkQJsiZgx/3kNcVrPw3vf13XRKQox3djOZ1t5LtBdFun7NsZ485JZt2hOKFQ0MEg8NlD
36RAE+WJ8wfoB5MS57lOVUWVsMZrxv6JbhKqinXT9xZSH8liKcvlDQcMFvVtQAlJ5sghdEVYf2Gz
qmXbW1s7bJic8Ksl0zk0xDLgTuUGLcXR7lgvJ36cKYw8WAxchGtSNurGIAM0p6CDmP2BfAeHDGUl
1GNODczmXudjg7TPceW9/O1WHa/T9sjCEZBRmq3djMZvH73bxCssReEkRD98an+YJ+7P5qyeO9f7
Sr2TjrS2Siw647W2gtPALqninsCdLXODPvt0h2n++pKsE+nemOUybvhTDFmU7Siz9rbpm4b0y7A6
ei2Gxt2RxmSSLBv9S9SrTrgbDzbmLpGdd76+xJkk8UeKFLoVhc3PVYd0TRU0nTJNfzWy1km2HKZ3
ayklIvjarnK1XvZf/MaJw3/9cF6xHnUqs4zOuu6cdDacRizB0KgQd+8U4Tu1hLO7Gc5UWbq4n11O
+b+mwEG0QaZ37QE4tQf8U11zG3Vd1mizVMQJh5AJY/VZh/lDsuESkFrNA7nPPVqpoVcsDOOPz3X+
xYacLBytKYkkrNpNtZKrJxYOKNfvKDJjSmK68pCHUY9kkh7Ld2bX/6G/XGq3WHgv7rUVSXLNSa5q
AONCoQtkCZOL5C07gBeYPEZLE0lMKcgXQ3ypYaTIJ12H+V2smMjZDtM6A/qWAORxdoAdrdjwG4TG
cqKezlsBbldz16g0VBLtjYz4y5IcmOwHEIRtPdcl1qdd7VT4dIafFlicwQ/hLrZRaaLpg0GahJxI
tfHSTmaG/v4Z899dGQuzn7wrGnwagpXhXJsSM2QYCcJYv2/jk5iJ+newnmZZQF+aeNUlbHY8yAZr
uTu0cEQTKyS+l5uVsiUAyyN/9D08Tj3UBYz3vZnuxx0wDfxIDmUUBMABY/xKz+vJSTscIpE4iwQe
n4P5ZIn+xxJ/Ldbiow56pqiDroxDHaiUQ3WdghybIxcZVrY+pTBVkV4nqezY1p+QoCLSBB7M9Tgc
oH611GNbYACRzVYrhREz4WMz6GLPFykUXBB/HibsR/5nAD+zBXYUIX679vLoq+yWKIoJqHjgpb3v
h0qnmzkTU8E8+ejfuS41m0YjwFtnk8XXp/J5xjpvntBPV7mIuFROmlZAEjdEQCt3azWIYwTC6/Zz
r30YQ4A1xEY8+6AXOsBX25yok64kpJiByYnPF9XCMFN6XVuwPOylfaCxmjVPOc9gvxXd/RoTQxQV
dlxH7nPLOey5P5maVZmEdYCdUmyYJQGTRu0ErFX2DF9dWyWVQ4llmm4VpQX0ktCnqIRsC+y3OAGZ
57u9ip41RN1bqSNv7sSx82fJo6SEyYXTCMaY6mj8kPdwbAKpupOqDaDKlxVkEbPet6aBw+HlGKZx
K+pgT2VPeFeizhMK4RQ5jIxDddsYSW708QcFXzsZlFKboNOE09nYQc2r1G+h2PZqG2Wq1nSp70iO
zGL9BfNDFjVAPobZ5k+UoTgCFXg5iEZMc1S/z/VM2ZGbZpOhghR8JrInTMkceAwczljjgej9PvWh
P1zxcitw4CCPEyFFNwpFUgQkuVTR0V7tvgZtM83K5nGg/gkO0JPzrR2k1/0mhtEgL4YfNrt6u/ji
d0xGTn+e6+Num0FB5uFo8kQVrf8UtKg2NofTTKbdg9OnfpOrIX2ND6zsDIFUum04BNLyBjD6bsdE
9UVQ3t0daiPGNxzjHIrXf/cOBqcHlmR9/hf/wBxvW6X5KYpMbHDhX2x5eRvNDFAl+Mrq7DoQY0dc
X6fzcrpnFIjx3Z7LETVipqjRV28JN59U++4V/2PtlSthCSFZwsk9auAkBdA+fnuCkbqDjT8eaAXj
VYIOhh1McUi4UoJZfVUmnyXd6PsBrcsKOlk57x/bW/x79fjA8LWqDGSuV6pY2ta3OZmielcMOHnc
fujw9URr2BysKJRJLQx+yJjNz/f5/euf64aF77VUTo77imqcfoDdG+pr++QDd+ZbDCaVJusvLqf5
oJPRtVxJTcw5pUm6xCoutIJ5flrRJWA+d4q6s3rCMUXh8U8rqgiOmdSilZEw5tywD7VN97YNOWp3
NQlPiUH8GsgBP5AwjHb+oufxujpLFpFTk/b1owp4sJqhzOyJTRUwbt/wUYlm2AG/7I6QEHSSs4bh
LkONaX6LsgELd1iGnN+cNCG5ScNxW4O0wRRvBybAErNNaKiBn2uy3huuLmkd9YgB3QFUV66o3c6O
dFsj8/XiDwYoDnphEbfIMm683Du8rmDkYAnL2/8J0zfywm3jMd9gs2B6e62gkYxTdJrRqPl7Tk8s
IwzdGWgK7XBkRUsXSlpmJeG7LHt6LVPKl7yHG6HlX485WgR4RX7Q0XpYR4AGWy9g6UZ9pn6szGWa
gp0hrSxORULXNAWYg9xzGVGGabHaOXRwIVZloKmRWtFKogA5XgI9BxHIdpbd9tOqRHhhirbXyTlD
FKffNHrNZ2+1X362kDfg975wjWJJTUDsYbpFHoUgRXwqGeQVS6to05xcJ3okjWivbyOtlj57TT6P
v4aFyTRvhj6EDFnEiUe4r2edWJ483J4D7nqGEHmQaY353f6PxO/HCoX7Vt9TQJLoWztqpHXKlyEH
WR3956KlltclHGkO0UUshF0FZ5RcBMCSosOS1AE12VU4QzWjbIq7/KT1uSLmoF+mPIFZnE2CBTq4
CxadnMSEwrQosEXj1Wu7y5xSzTfMiNFSV0WsWOzDgrVnQ+4PsA6uDNz4jRRMb9uqjIpZb56PswpY
yHKXrwzFdChu4GwRuwKIyqzTTm6FJmetOEY5juPdYjFw4i+F6PXXSt9dBPqyvfYq9g5TWC0fbFou
8TKAbUjuXzZN4f0izraL1k9gsk+pog1v+RElHS/ZVl5bEoyZZ52vG1OqBZq/Z/fSTYjRIDCx4OOF
88AFrsaBBy0BFWGri2J4SRIGWWbFfOe+CoBHAngs3AaMY3xXvfodBbvHmgU/eo46Rq9YEC6HQczk
aTsG/k0zWJpu11HFZi3poFvmCOHPraa6WsQE+Fysp9NFMQQY1+dPNlGVL9W4k7GBdiW5NV3awZ9L
fRTD8c2zV3TjIPAPA1evQMN+NCD+Oz7rJU7Um+Pnsc8fAtuRofbpRkxhGqyoIsU3Y0rBzjLElQ1O
owuKGQinI4yN1p6BQA4kfgeNHz/tNNeCii738DfGscO6nrs6nplTy5zLydgXzodpPT9inC6zTGwW
EXeBTPO/XVdpu4uSVBmlQA3l0CPWwnmbRFc3R8mHzXMdZUdb0f4kY2VbX3xMvALYxOY2IAQemadv
BYShDILAE/rc0Pira+/IRy1ttdTn52Dh6by3BrzC6Li5Qx6dhSu5h18vIjPzsUJhIwhDJlt+KweO
V9AsXPmQy4IYMw5aYNwnOykeV8zO9mto+Zv4Z69hOGS05xYksaNkFbrusWQAF+8i44fqtMnOfZy5
FacvWUzcPPwRnZeE/ST9xEvCTxraOBFt13Oka3UGkSjbLwwKv3OuZaNJbOJ/pphOufqu922+c16c
pVXPffTKZ/TByxE2QxBocMUJMWXYFY59aaDE+8TDN7zm8S6qi+WryskwyfqwnN+kojZodQwYyzeu
f0Rpa7RvsYxGB0vPEsD5FOcHatBj/MJoDplAWZDwncWoEkTTWj2oCsO1Q74IlBbCpVh2WMsCQEec
5xK53kcnNfQi2eQFmFQAACGlxF1KBz5tj+b0AcDF76BBPgrDIkhJTr0zqoT1Gs+cwQf5fyYA4VmE
TVpFUQmzK2aQgfjrufna52DroYd6v2cranPDulQBmOikI5e37gVDv5gQdG13/EfYOUPNLxo4rvh2
aqcO84NUYRyhVbGGw4/OBXQlmfLAK5sS17n+gp9cs6vYyeAeY+4hz5RhyjZjp/OPXauyT5DzgIco
EVcGVvAn6AdNMCTsjtTlnX4BwvOdwmAIuHAXuwRANOW6VlFT4rmOXFQsZIFagcu/1vd8gcg0KG/H
8AA5MhLm7u5+XsZY3TyBxMI7VT55gT/ZSL3QRHSbi2NSiwOmdlFTlEd/lj2Lg5A/C24tfWlonh2z
QR0wGypTJU0QQ2kzIM9R4bXed16s85Zk5VtsTIzWUHZ/KVBdkyXf+pP3wE88B1JIlTAsVtCtfWFX
QDchFcAplXmEOKeSkkXOdM6WzlrwkWz/qXqICk8JYIA/oLzL+TMWk1EioX/dHJMXWIBaA445SRaI
xPvx5LuUefvJQj+Rn9SnPHhVn+EwUe8hHSeDGIxsKPVP9mZwwMk08Vb74iCr2yvCwUhwFc7UAn9c
lYoTAhgnTAVqIBPrnaEdkxv/NJqzhrEMrsIpxXnM+YMc1eC8Le9k/LfwnnrfGeVH6L0egjDtng6j
Luk1aQHxmKw8gtjeIpCWbtc42SAtAwWCHKFWsmD9zlG+3Un/d1AKIApYudZzQr5nh6ZkcjroBv9X
S0v5kYB8PFkS+kKurJ7p8X3YdrEvb7fCSGoeIlHuaoTrvmODiUAyDWOiUl9DRG5hbxQsPhu89pA2
RwaHOMl4wlvZQ9lpk63vWUO5xsXhOvbtELi4vHXLlaOMqPAXWLuqz/aaFLpb1WnpIB2s1EoUS81S
cR2uNPSvmZm403fzist3A+SpZ1iXsTyEtEPhWmzeNT3CrFe5D1PdudUXfjPLPjxYLuQCSP8w4R0o
aggSrXYpS34FYI3bvkRc5E+yb7vdp1QiouQBtDYQJX01qU9L/VhgyP0UjsLj9Imkd2MHKq4DS9e8
4kCVeL7go8yJh77/pm3k/aXp9Rv6LlVx1oHVWNKpHJmyBtF595mhr7xbpFD0e2yNZOaBwMg/DZFx
foCvsZJAqOdi8rR8J8SwNkyxQ52quf43wuaqiKkiEDE3OTMeaAIthfbDArYprjBZUIWQ5AY4rdKp
AuHHBaGBIG5h338/QRUecnQ1a24o0TX+QcIoWItVz/2dE1XKms7/wyikAkWHlfpnPgEvcnqzkb2R
q3+olFQ3Ch/dShmRAtWaVc9nOU80A8MoB+ek7RnNlCJJRG2d1GJixgc0eUtaabv0RNwWmmAMXs5I
i+jVrM3JzvnyfoR+B/UmLf+csERin62s1Vfw2TnN5Fuo2HOsLl2swhyWbZmthuM6JGn3ujKGvXd4
7ggCsyg/M53L9GE4e0vks/rbqk6+H/DGesPnjxt1+SIe1djhWQ/Wkp3vh0z95VTkgXL96l+svcbl
w+CRqTDtQ8/GrA4uBL5U81YDb25XBTRND0kPoFk3TK6O56YbkUTFbhWLnhjzkik8hLB0zZk2zdJ+
5ZIGdnckvYT1JrfVSbpTQhPX/iOBagb/+pCIY2muSIvOAineGi7kgcxgPEHf2xTVPuKl89tkoY5w
UhIyGhwZHr1fPT4cNqFBhJe0jJSZjU4JJd89wga5wpLkZr3FcXV9dJgrdBor5NQ/Y1IfsLmyQ4xj
RVoQdXRuHj+IpGC1akluRMUPcuP6kfUTXoqeG/Ggh1fF+0JRI/+jcsZyxxqu3Y2n5TmkYcpVYx6o
JvjREipMRyHAIO4u2iPdVbtnylozaZwV7H04iRztQy5EGQjQ7mYfq4LITRcPLVHdHTlwhyn4grEw
7ced5d3l97fsnAuRxptf9fWp3zeXncRpCOoH1t1Twig1wtqC4Tpy/69ELy8lvUuxQQZAZz52soOB
MsNMFaoCac/46ImZVWOqotCNgeMRefzMYV5dU9QlINYBukOs2M1zlr61ozhjU0ebxTWrYdHycqjO
jHlC/CaWV3q/B+uOkA3J3bEub8n5JH0CnhtsQZyG5qa15lJLKLRogeYoB/uGoB/87Id7IAMPL8+9
UophDnB8Dm6KLA7ds7LKVqCzRsDSfZCwyzQlViun2y7FxtOOAfrbYlAELXpsFzSttiAfs05noFwm
PVkueKxpIiYrWFRviXCJKJgIKDd2mAo9keLiiMUwRYqMWAoUkVnl2qAEaeXs/QETSUdUxA/q2alp
7nNDoY0Wtm95jt0XpK62DPfPUFVcRQvfFK1PqnaKylV5K/csnBmuJ+LV0fYORaeRV1ADe9pYuqX8
blsU6320v2HkIL1fFV6H9BwSk7NWXnySzW5XL5vIzSCp5bmvSGyY46ZdsTJYwX74QQiyUuJF2XtN
Sx9KnbqiUoUhZ0yTi2i+kLfa//wljIIzapMDfkJVrLWc40mrohIbLNIb60igRl88iR+IqPO+7o6T
0Dj5OPw1YOfH6W76/Y2piJ+hqlYQmAFmpL7ubgB+V49qTtfIgusFdCpGHcZ0xTG/xB6mT8N74OMU
qys1XDSLwVvAGBI2HsBzR8plbiTI50o23GeGwDa5KpJPPr7A5OGH2G/4lrKU1Os64LTokf5W7D2f
gJ7kXHxY0bYhJ+i/aKg+XP49XdEB+2h9d4QPsCB6RAHjrMnFKjMMEG0DhjFWKgzchyNTJcRY0JFy
WuC7KuURGW3VF89K0kyo42V2ldGF6ydWi46eDc2HM5hIw75EigUFTfc3oTtB1MmjdRgnkmrKdls2
h7nF34rJVJ1Ng9ixFfFcYh6vEULWWQcgZOATD1puN4KqoBNlsUycArlYMaSzOGpd8du3F2rB1lkj
wk2GJVGzdR41Kh3cpEke2WdmysAyWE1qsNtHJL8D9LCNkEGEucYcM5dr4c8UkhDnQPjlXHXK/1Sq
AFVLhR035WeswWRuywuAbHuRqMDksNO9oEk+eyG02zuGBtC+sPiO1XsCkqBFAKehmuvgfIxQ8DCm
0ve40iyDEQzbXrCaKxafZ01QMhID30EsMxzOcKGipdsJs9tPCZMz0CetQzDGWCLF90cGVUdE7eZM
hA1kF2dDrzVdWcGcCQumWZBXE3FH+vi25N35ovr6+IccfSq7evk+hlv8//LDrroDZvnUo2v1WG9J
wjBZJQLldFEvKPsAjodoxC4l9aJ8eZlIjphmmyZgTmUAgvrfaZhvVqukVaJndGMXPb8SIKMR8oec
UCz/xLRZ700z+QUiqDOoPW7oUgt6MoPP1GxzFomuvcSW2CoY54pwmld0sNFhyIxEsGtY2DIIb1W+
BsDKIUwFKuGOE1TtExSxvpF0tSUQhKFHlJngnfCrwG2HP7Tjp2hNL5G68cQrEDz5CcasywWHTuNZ
NImngIfBissq6n08eXCNW4I7nU4rdoWcHuSdJGHUn3JwcNgmz2SzRi7SieRryUM0agjCz209ww62
nzX8Tskne+dbjIxQIr8wZ0alJwQia6UN1bJA6qL1JyozseOSuRGar83zE9MjFelR3LjY1TDdn5t2
ObPWg/aNveMOJZX3ennhv09Ebe0iXGKw9U+lvF/NEPbdvvlq8NVE7apOSKcvnU5RymS8WDkRvec8
SkzqdTL5EJxMuyILhrlkUQ0WEkaMXm4lhqfDweKzP7Q9zzttfRInNPiDkJtGakn/PRyoftqkGYUO
xBfzauQmcKNoPc/e2gq5uO5dQHIkbCW67fORMOkzzWmQLnq2vGASSkCofmZ3uU1Fxeyt+vj6oqvN
gk2Dw28yVUUgn2neTyi6StqdvDTnPbz5ARHCe/nxLka8+ibGBtMgWLNzUVLo9jynA9o8LPX3C+6v
ddhJWzXog9TBM+c1ZrkKvOL0xRqeeEATOsYVDKSDKGKKtqSxZGBCPL07MoB/RG31KIRRdFjPmcPU
+VCPinEVzgCzFU0FvjiisO2qTRNVojtuyYQ286hRKccgie40pr7Od3adTa5ggCEQcpuQLBWFYA8X
Aq4JyHerln/oChzIghRf9W2jzIRB7Rtw51zVWuDloK+mbWQb46ZRM1/tTIuaxxYO7KhzcOMtMqtK
dnog2L801XZNLEI+szqeY4mI7NFhNximIdYTmfeKuSZF+0ZIL6Y5A65sM+77OroBmLFWTIUGO6Ly
AKBqHJDd6jt7fbtvZSuAYRJuVb4pLyJ2X4Hu2Kc4Sgh0nP7GqnkjBSKk2I9o4kBVy8gpiFR085fE
fZPOvqlJe3sgOcwoFPfsZm1/GzvX7pcKSDUMyIRwfIz/wMgnHIGiZATXb7sldm3VB3/oCdPagAcg
EyUF5/+mHTlwVNswzs4BZ8OKiknYpyENgYSdHKv+5lrD8eMrm8Z23h3IUtx7p3A8HZ5kYwu0lxLb
lxdMV9U/UR/0qHAgDjov9TMDAPg3WIbIwMeXQESCMfo5lOGRHFvw/aTBdhw9HzOb+8nImea4RXa3
h889YmJYSeqkSy2zNvm9SqyiGgCYV233m8tHIYuzfdgp3uyzmm1eiq6Yt26vRlzPydpcnYzpprjt
RVXw/PhpuDcqd/Grd8daj0Vs6HS4cKgEaER45J4+HGGH+fQ98NhHCfAKqg4yqy3cipuXPVGv+zoT
ukrjNlv28UoJqRUjaexaG7U+/M6POoEyNOeUcDKk+1CN122sDJ4IYy8Ei8UWOsTh0RiO3uupF85n
QyAOH8n96MDlFFsqLwi2Iu4V/N4YVlFeOT9E2RxgFBl3R64f1pt2iaHL7e1NXT0S7YoMYKc0nIaC
SC3HhakNukZOQnzZ6aIqej7m2syWp+Y2BTevIaJB6PUyf9AtrmESq765/ekZrErkxRARNW4/UFYk
Fisnk/6iM4xjJkpwenLaoiW7W4xYPOaqD3vxWyPOThBMKr8tGz+YPyPaXfxg9j8msxhhkVfRekf3
MK1NHTKT+XIRZ/hPytcpA/Xw28XV0+JDGawcnoSF0CtejDQHDa79UdiSCNIRyN5a8qc/IwSqIxt3
78D5TH6h5iMsEwLVHkQ+YPSOcZFigWQCF1YjJXJDCVQ0b1E8VB6y+19s885PTEUbnzzYrhOQCsB4
jlc+2aHsHlC5WhPeH1NiUwSMNCKI2SH9w/e/8MqisRMWfWQ0mZJcJCSd8qeJBY93cb4j9kmNF0QN
LqH/bR8wi7o/n+B+teZa5T/QHpItXZl0OJ/ALuqFYtYgw2O3kQP4sxQN/tTCBCpHZRwqjdqkpMZV
kLzVTMlt71yXSw6eZVSuiMUXU8jq9VO3XFOw9AXT2ulfdwbe8VJEwmKWcQ08Yhzwc2eqQ6LxMPRp
W7tlxZBJsu+z+qsoEkm49+8b4MkG5diMQdE1m7SuYF4HqgV0Muy6uoFrhHbix4rj/Gi+UTeSwoAx
eY039xCQ1PDGHB45pg1q1+xt9PGgL6RCHLK9GvMcAk3eX8jZeGyTMaWJoVF+mgvRx+oCj97aAq9t
bVLR0t9xdWTAhIymH93EXGRXEgvdmLknu1gONpLfmNSBnjqZhMseJbDYFxKpVNtq95ZBp6iAw7DZ
3gis66asLm1TWXsk6vqNQDelZTfdNbH2PSTwTOfVOrKtUE4lyLrHJF3ee1xapV2kRxznuUuT2wWQ
bwr+amNUVGPNQ1rY9D4kQ1fsrCtcP5FtmaooGvCHPUNJZW+X8CMIwwgAnntS0pKrvdzDPwre+oLc
8FrEHeRL35ykEa58oPFOJH3+vVg2q7BslCk8vpRE86wduJqMwRFlw+8LnP1ZP1XXUp+KLW9JdjaO
AL7HmKQvQPg1e4MVPgfRTPG7jnE0m8k7Gy+Hq2pHBneIdp8t5bBbdy6/B5AxV23fL1vuWQgUtmOh
dCse84FeaVpZ9zr+QqI7/gVcfK3JQTb/CeAEoSDtWQ3qArKxPmiUUH86+uYXXOxQBobsaikOjggj
Vk1xSEjQ84lxEQYyMeylS6vvTUp/grll8+XXfknSTP1zqMdKQAbf6rAMq/CFXujlWXc9C6oKHBgA
av4CagjZ6j4T8qoTu+SrJmKEmpdL5Bnhnpja5Ftow6PCa5YaX0S0AMK3aS597oMHSY6v5bZvVrAf
jlKNzkcFT6Mq2LubtqJC/CcHyBIo8AY0wAZvt1uTQQiLaRDZBVWk81zdP5aFOnen+uJLrhndP6ki
wkGvO6iHSmryOZemsfgFq56q7ATltz+gi0zF80rzyssqp1qB4ujMf5qoI1291hHXfZpPqlE4KdkW
eMNhH/teri2x2ecuWdBe14wqsKIIojnfsfzP4GcjVqmpqMPQwCiX+qU0MkScz2jv3Oa8J/vtsTuq
f5SVrdZYZlnbWlM3X81cfjzm6ueDmL4c3JULhDYyac8CzDnhHev1EVwXgvuMC4ah2LqKow3gTw46
iQ2GvtxbPK0epoRDLtbN58oxCbQxmKae8TnTXnbBlz06qoA6Ci/EUAFf+kC2nagmuiRHnAeMwyRA
+wcUvw708JuO/NrXnefzQ6mjV8i7Dv+jnfnzu9jGIw6XP/R+1HHv15hrUfUKOyJ4Hf+4g8vAWHhR
UozFBFnO1Y0N9YNA9nkwQTl5wGV4XHrR3UodVro4O1RVFY45LnrCxzBTLF76aymo6CNyr8Sv9IdM
jDuEfSBTxxP1FAVCasizuOWspfvCxeijpi20fzbqsvvH+Su5a1QNG+eAKqw72tLM629AMF6oKEV2
QhPEi+skMpmz8Uw+fJt2pw2BGx/sCKEGWsrwFPvJGQ6M5/5h7CpRA/IrADFVfuD9lnGF8nggSUmD
E8htNJTk0K60RRD9bqZKJwY78fI9mBMekQKYiQeI/4oRWqC+KdKBo46N0joFVFLOczgOzviuIBWq
iyVcajtl56eUQFpAB3LStU0fGC23frZvniIMobodHHZ9ZI7RhfoTAD6sy7ThqlpA8c5/x9h5N+lW
9qBVxahwjSXGGyKXS97kxszWg3waBE1G56bwydAmce+PvyyxO8uQMhrKO1fTKIe+kYTV5kLAxZX0
QPjFn0v5CqEMy82YQHzfNCnd0nhCIF0/COJN6wiNdsp0sVjAjYM351/fxD8zxg8Q42TCypOxyWTJ
Ohjth9P3BpHfiaUgE0nXUC8qMM+oDZvEe9kytb3lcra0G7aZEfOC/DUtpkzNjDtS/pwiD977Y/Hm
TTMklItv9ZL+jnI4cBEajARPx4TpllpZt4Asfu69XFS6NNOVvCvwlnffXLusrbZRA7Llb0YHtHdb
cflpuysq165KGuVttoM3wQK5S0TPSFjTj8/mv0Hdum9/XbEnxqx0Ol6ZXob2AWaZ/uJW3nVYlZ6j
bhrCZmt7UX7rue3/b9OO/zL2tUrZDc5unr5p/lRoJdwPMaGb09m1YCYpaj9IrClXFOZFHborSmAh
hRIHXzcjD/zO3Fb4S7yahMTjuzSZfaN2WmctcJhn0n9rHXBOCvMb60XoAXoAC1RARoBbRHvkKpnx
Fufy7zmen8BSAdxVsbSfQpl8Pqw2ZalQOCnhi4dccDnu1Gco5mIyEudxW5rpF61wShuVgsK+vQqV
u3RVWgk0CtMTKHuQjMeJkia5rvOk/zwjfy1vV4pGwIPsl1MzIryRO8mbAc82EPmO8U2rOo164FqG
YF+0X0kmuVIGFTs32YT23mpVWdD3JnTy2TzWQ5ByMJjcosd509HN6oOBZAB6rkfUXcvczoy03YYO
3a47Ap6DaN3txe+BGwnBPpm8BQ5gxUd/gbwslJyj2csF9rFeh3L3BOWimGcYlP9d0PiZyuQ2++CE
qOQGKgGdP5DV0Ce/kezcWXLsdQexzHEbyWGhV1RO+vkaX+PCCIAAMVjM6sqhQeoHzoPUrT2EQJTi
uI6dNn582Y629yr8nDGCJDhJym0JrIJW+dYh8fX7ShMHRelQh70R7/iovD/un42ChTagMaSfZ1I4
OiX6UChg8Wju7WhKKIXye4YOASZeoEcs904H0E82cDLs9Ttmmi4RabaL7fZXoEvF8K+N6l/tLPq2
nF8WJWPnIZgyymGX5eZys9/e2fatn0ETdyqV84ljhZlQdFNN+Jzh1lpodExCosgv5g2fxu78MlY7
KLyVHQCOiwmtye3/TClFDjCP0lXGClMBz4yppHnRPenpjnsFw2nfyw7guQqyoYpL7pSJzAOqwopt
QUK/jMh2hshvzy3sBWBTAHS9gVgDgY+cirQXyxunJnusVBHUjIBCa7nuzXz5c9LMAhmbcJSI/iHO
+oYneQ5/eCbhCubVBkO7nE/gGG971K4CiU3TZHZtH0bBvGzR0BFX/srBXSy82lnVPQYASU2VZCNP
PHl559It2bGN9aAKY6uIlZALoUv9GPLw9oudID867GWSjryzagemNVHZbzeW8k4f6SVRmloJsuSf
Y+vp+8xUSlJ6eclNj11pxOCRANh5A83mwKKCTvVKmpX/7avegO/mnam4eNJvNyaymBaY0kojIGqs
GKnlowusV7joRj7/LafA1JIh2xq6R9Q1WE7y5eSQzi3RnZBYd4a9dZg/9MN/oD9XruXDgbaJ1LLJ
//N94PeHZxQYPEg3f404Xft4mr+j4jQusyz2sci8/HIAziYAU0Kwc4iqLHY8yeyno0xgsj/p9B/R
wGsvSsINB0ChSHlgk20YNXnsy+pTme7XRkFmrRpEnOYbu9kWzex97LqmxiYnFcEyYqmZlkyoI6Xv
30hW4x440aIESwvWVadhHt1gyelImrnCaPs3W4nP57SZNsqZnTDSXMNrNpJvC6blslrUysaxhWCc
+UvP4bdhCkpbZgI7COrme9J1b6kMArhqDBV4E+8QZSz5ztEObQ11z8s/kethbm8W4ZDrbptTSQqQ
w+zeJexug19fRCGhmUs3/KwCoyLFzRao6okmBothDbIKPQzhYALvYHFZqILQcsj6vXb8v7Lf54UA
u3QDc9FEMBQgH659VMVORdTXuUo7BQMa6Ga4zzCyoimwIA5iBPV0j2pcFoJBhB87QK4wCvPxT2QC
nyBgg7ZnYLl719APPcKNPzQvby9J1KKtg/JmiI6ekSwel/GR3Ulb4sxfEyHG3LxjIRUmjscSfhLE
OeYcnd/cHv0ZtgD832vqLebdBRLVWK7n/4YQJfgD8on8YJhyKNutow95CutYhMq5aG8QYhFxgO2X
xwwwvypCXSSgLgSUbCaTgcvG/haUssJfOh1O6QzaFMEW6fUuw4cgCKa+1qiFmn7GTKfbLj9Sr6u8
YVb1dxYwYpLid1f13Ldo2BgwB+P3FJYi7UwjnZGo231pQZE1OdjOlujX+zt9CeEdhMpl/EmMpSsm
plxaWCw9l8P18Rvopxs7ugZEY6Wvjgs1PpEHRVdXYOuzH7LSP5r4FdCjqEXQwGX1IJ3BCrZsBCz6
yiO+JxmD0VB2Njd4fFqus9ro9IViDp5n+pTCs4bBBLyv4AKIG1BqEqd6h9W0YurlFCn7eiBJId5x
11Oz5m4Ph9FsrQwLLv+aGJclQxNYlDCXPBd/1vmMqSmSMQctinEF+qcyW31KzLovEVbvJ5ZQs3yS
2NnQR03tQMkW9xPf8CJUy69SllAyjClIZ8ZN1DKz0rrNPM1GaTgvSMM7dYTjKjronMbg5Wu/4DFK
v9/3IVVeI1opMGxDFaD/Rmx43H8Onsc/fgEx7B06RoOveg8pBhpAdTnsBchK7eI+Fw0kxrGhPkoU
L+hHxwdC7vDv80J7B3nOGKcMGlUeDAgmuI0Of4rG2q2oB30VuUhuO8alWEK0nM8o5qdg8SBEK/JX
++6l8S0UsJWccVx8UIcm8doEZwcL6dr0P88mlcXCTrKGLlNGoQXJJICfgsJwN7K03JM/vjLVwM5t
0P7Vq3azVkeXXbDe8CSHVnaPfDRbgFYJMXRerUe2IXmYCEsPgXPCVyHt3r4k4PYuht+CpK9bLxVM
Cu+o3vgsdx/hdYf3stFhviFRQVemggRja9MAMklFY0fnGvK6TYkYhNgcytcXTLFIpRJ92/hTKsa2
yEaocaZj+L9WlG+T/YHgu5ASJaUKrtKPdjMBUb0KfaxxaoxZrttn+NYocCJMD5+wzgD4ir2XSDLY
K024tYNCi9T4MHU62+XM+V4wcQpX6gtTLb9EGmOzzSxbqhNMU26F0RSr1sBaR972bzB1al0+CPam
O/v+hDfeoRpeyjz5YxCk8Rv/RP+uW5JGpzouy8NrPqBzon4xsgIom9Yg/CHUoKP/QamwX7pgTF4W
w9V0kHMcP1tjz9Hcs3z4YrqSrdaY3VvF9jV10Qv+pXQOBSGobEeATTyGMJreGMvSro4f4xoQtduj
1nJql8p/vE8rO/UTnEFDiZHjHgERfGJDGsLEwnuORVlCG8lCvhajlVr4TNr1TtCJ3ow01f/ySlIP
cKqLxsAYlxdBSqXl2htgYVvdWH5bPaHUoFbVI2emvKahDt29q+6Bsdu4KSXQlEHGkzyHb2wA1apv
10dY9VYkrZOhlBmwxQ2aXEUuFb27mfTrnrdhnuPNo4XLykpg4HNr8LzJTgWuAyfibzkOCmjfCoAH
JJYLf0xyu+98KvVTpG/3HysIuvOwkhop9WmYeh7vl+M1yCbBop2GIxDei4fUw1Fc2e7V4sKLK6+Z
jTIqgUXYGB1Lqq+yBp7Q4YUvLUnqJ/yGT6y6axuRhBF8sSgF8BthuNdYTjLHg990MgYz87QJTGGq
DoDJRo58wlckdUQ8cEBfkVz7LJAiWbGnlec4UocKJbCDfnk7irfw8WO5nnUPPa1DLMDHgEutuIdo
93F7B+I4qKB0rTCvHFHm9ku6+ojaQfePsinck0/EEC+8nGRO7IQeMo0K1Qdj3Hm6Q/UB95FhOdSJ
S6aOQgo7AnvJqWBYvzLtte0/kU/G9Mnw3sD3B+gwypi+HLogC7ZDTs9mW9Ns5shzJNuiz4c6TqH5
LiJB3Y+uYZMzZCrVGmi99B9WC3yheNcZJ9OaxaSqPpi1h+G3ABcNg9pLIxYUMTJFucJdeIxXDWqw
SDGIsg6A+WTgWCvgbTIRqPnsxHpVqp5rMA2hcP6wRoXDBpAdJonqj7zgmZhD5ty8/iJU24j5ls2O
iLLNF/eikwK34BO4QQJZjJg82KXq4DFRhCrjaeC63uHB0srtrJkF+f3e9/HVDowt4L9kdOqkVgVc
4Q78b++V0EkE46ErxDPjoWaHAG9iM01mTV2FVhALgstKZM/kBEFQ24xASRLdMzNKQc+o36xgAaee
oj3lFn+hJvXx7EvBvxfCmvNmL8bg90cGmfxWGsAY19RxCDIO04sB984HkPealwCOh3D0nqhsfmha
1h44ihbLCZXI/lhFxuB2de9ScDy/8Ws6t+mNkgUpJuhR7qpGyJc+LxlGcclu4DULxgWsVVL2YK+i
AqbVwnsC6Y1/dycxytlQwWhFAiGKDyZG0A4X7E/cHTgQIZ6rxfjXp1mAaIg9SgDKWJ6vdoJEaz5u
pkg/YHFP2cnZ/nIxEol/ftPYLWA31ZIXHTQptbq+V+Q7E7AiAymmCZNR3tc5b/09317tbziAR0Ni
MD6Ws6UMBzTJfWeGPrbZ2Kga/SfYJILVUyfF2FqZAxPK90y9qt7W7V4wt1Pjts8Sm4qFr/x1ssDo
isGWHwprUPuGMn2gCzjy2n8Tsb6+xziGDcBHVRXBaZq5jFen60u8HNOfMComKjxhWmPBXuSoxJcT
KQg4d+m1jDsrKFPp2WENZPRX1dfARqA/wbmRN8MPgOF0+UP0RFU7k1OoMtMOVNqVE0YpVW/5QHNO
uopHCMU6swnS7x3NKRgFeUHJ33DG2uTwUSUMMz3JTvqmvn1XMAE2zYRRyZqll+5jdgrZPXGSPBI+
hupjTvtULkJqdxWb8U5fBH68G9m6kdq1vzNO4pYF7+U4VFQNI7jP4hKW6VsYx6QnUOGdm2VD06r1
tZ8QwmILvEm207/Zl83PXsbxpv8mggrEZnm82s4Ck1D+RBdjowODkyVvmxWcRNrNCEwx/Yl3qnIK
6DF08d8qOF+SRYQvjkeYN5fjpt5SNNA3n7oxZtAZODudZiuQQA121axv+fZ73zPG/4/qK918wpTq
Ur/6KVobutkRL49O2vFlcmZXsJFipzKX/olZQTYuuo/IA3Njc5BPdj+IVryPTNAfQ0yg5W/bzRyj
T7hBidRfznj9QcFHx6/Z0RdJoffkQCpvzfn1BY/gOxMyAjsO/zv6SJOH32fWNWmU6lpSNdYX7Gjf
i/4+6VFQVAisIrL318OfMxKNxjvblB9hARJxfy1XK3FPo43WxAq4SFybulGjUT10k2zMrBFG1ruR
woXpobpXoO49TfE2DE7A8Ra1HwUQdK69MMFHh463K72DurkRqKcPZXZY7bpYgLezX7Ce3hUpYqYR
fChPOtW5p1/lE8nAJE2Q5zjG7aoYZX3Tms73b4ZDWx0B4QK3svpHRD10B70Wr66KSdocxQntZkNW
9PnTwl8TFex0dvfvTdMBRxHYR/V5UrOsPJ+RX9yFPxbg9rRdGjJ07cgVL+vexUrRodm1uQwDoBp8
BS5chRR9RkEOuibQOPkst+K+oy2enxQoig1XH2RKPZjXavczvTxrp6y33IHIevRJWF8Cf4traABF
EXSqsJ76opMUpTd/cCdvkQjk0h6kj5Mptso7/vdzBiBOkop/7PsKcDJeKUy78V45FghwbnAAzsvk
9Sgo0coI+7WMUyUDZ2K1wmIARqegdFBjV0eNPOObBnmMgcQIcYzH6lwpTrUL+kqXNYyX0/u5IXk4
GtOxTDSy/GdlzTFXboM/UY6/QjXlppLVzwH9lKNBlu4HwfhH0KxImKv2W59coyPFBfbxytLXJG0m
4QBbWRYiq9VdsMyGCMjN6YGwHEzmhRFkFOOEQ3VAKKFlQU2CSZxnSt4U1m4xRDAx0od0emnBQ2RP
Y4QxAegK5febM63mMWs0hjTGw7ZxhCo6Rq0ykcqaHxr17C1VWRbp7CjENrcR4L7SyFq2pTfF/FCL
SAkJTWRMTMK1fWJBxAUMBGPF/NuOtdP/LfH6zmhmZS64L6glFcMOGGeMCQkeYRQrEUjP5CAyJKbC
GKYwAZL+Dr1ZsJZHaAHqkwFu0PWjSAInMQy+YSoom+jly5wbxO8dBJ3Z6YnhDdOhGgQl21uGXdt1
Pe0Bu2hFz7q5KR+yy9Hv3PFcyeJD8PVyTlFoYpJQqfD6uwkNWTZGwnsc9ynNmfmwH1Aqe0yAVaUS
XAcqhF+oRbl74je2vcms0ZA8jopfP4m1DXPX5Iltc7nd6UbHkbLggYS6e/yVJpgxlJd6ZPY4MWbG
PXOsrfwK3SC6xZCkM7FwR+4wD2P7NO83QbTRTYF8X/oLU/Nak4bVu4ayBXKLwlhT6wpp6G0B+B/1
ff4S+pkHaUNKvsuGAvLGoPN2XVJpug4Gg90JoWrweUF2eMiKr3115/ROKid1yrm22PaXgDnJjmPz
OCmWOvcC0o2AIXOdvJ6j0TByoF7t66udSovxNTM1JcIRnlgx/GgwoV2/5mUDdrny8Rn/yy3caj7v
D8JDW/8JShMNKR2PFMuCx0K6nFPc62GqHDlvxBOxplRB8cFMptR3rYyxC2c/ODl7VxCElEZ/GWtP
kD1FkcVoWwQ2nZaS/7AsqtUaTIQVG27n6VPWJSu5KF8oN/czZQPIL/qnvnxD2vEytZw27voBiLUQ
6ahrcZXsD43qqDLD9kXCeDoDeYEH86tzE14SSjDMzqTaK17xxGTYJvIfxhEyWvSorv6OshFNvAkm
z7aMgO2v/6Pjt3Ke/VLzekYpzxzmgPw1GNRLIDb94Mz/LdLJJp3tl7psEyOXhTlCC8oNZoV9QLRQ
1x7UJdiQMsM3DNsGRCPBoe4+8LatMv6/m55B5eenHcs/Is3NFCaqtpYq2kHAtl85pIib4CCdbHUp
fEk+d48KSinjBVPiRsPFnccmyJEkerkzd93CD+HxhKYsUiaA/cOQ4yP+FkgoAcns2VxHYtInIfcC
ab3357wu3DCrwYZyY/VrTJ4Wgv/ALCgLBQw2nNVmXURxgoLFDQPb60Qex9PTkrU72lKfV6BHwGyw
CM+IX72wTsheyU39arTmKt3topK1GgbxSti4ObtMpnygVKG2l70d/LHclfzEcRfzIHj57yGkOpD8
rQxjOdMSeJxmxcia+iAXyclf78+n5jIjoxrwqdAE8A2neE/I5l4BxVZTpJDxJOUvs6qYiF/uBE2L
XYpDDeoueNPyOFRGg2RSUljhfJ5uM23dXtfLWzO/QbManwtCuQujcfCxoe9FQ0PUUQlIV81Tc9Mx
XigU71naLpsenUKKG1mXK18DKTgffMs5ezo/9TsbTPSEq5ASy9Y/L+NWl0+yL8LeVWHORGiaoP1i
xBb5QI8z1J5ejWsYSQYDNVVgcN/WA0CZ8G71HEC3ZiuVBtsM5AOyJxhq54deeHh1UXwAhX2AR+pR
Olyase8lMdu/ABtB01/BLBrsbAid8GSh3GBXjtVdeqqOFqcpZ8CS5RpJAzqtPMlwGwq/e2nWx3fz
afKbZBlMIa17HZ94RPj4b4jqJRr0ywAApSImsXdaXPK05Sq3NruobhiLHX0EgS3zZzHkjdFfCnOe
6X750VmZI2Ms14XkKw6jezn+pzbOQ2Jtr5VE7zN/eVQWZraACZWNMSTQVhIn2IHLCfC6xJk/cTbE
ZbZ/jd55e4xdBYA8SUDRGKzJzj9R0T2pLqZG7Rg6h9IB8VmeGuSRjYvqUaOaOM6Ol9yxrEcz0LsC
9CLGZ0NlvWAJ/DCUNZlOOXsxyf/fgvupOZFksqPe7kgsNun9GFFgcBLSJGDGjPHwAMwvx+v+OsBy
fF4qXKQUu/9rQ3twm1TXA5Q89f7dpVmsNtPegrp5tY0oH15Iu74EqxxAYxjjMhDmO7sXyrZGwWAY
bFv0GpfMXonRcOgm7Yolmi4Wkl2ImoGtla2ckk6fsXc/8Q7+0yS2ZsSovyop/woJUvaGS5MJWBfo
KWBueXe2YYKyYCJtLpk6ckSIL7Daw62ubbSq67BlD6nnWh0xUa7D5KUiQG4gHDVLCAfnRIrcV2ud
uomGrFaJFLP/LmOwcQxOGq0UT5coEuuJWGrwH3rkD+Nzk/8clOkW5tk81lfkoRi63ukxV5xgZMnE
ElIJQlT3WKU/KT5G2RjCIQzAsJacfd5kOrW7DIXnSvFatCvwIMdPwkaOMXNBP/9bcWMwxAc/+5cw
Ob7VjgJN54p0xUmcELbSlWasmFcKY8ALTlEW6zZvbS/0jqDC+P2I2u/B1I9NLIszsKeN3XaSS1J5
PUUCBZ7ofxE36etZfpaTVNCbdDcsriWZbYgGMshEvrBfR0NjGc2SOG3BVDmFTpPdTRS9RjbmYo9a
kri4FehRSYvmyAgo6eKXz0a5k6BZEgixUh8IOJAh64pw9viAaAVQKCc/zXJl9MNlB7CNhAVxuarc
QGSVf7JanljHDiTqzL/4pCncOrnLmUCUj1m0phWcclK8obOxPfLtCY61Glt0CNT6nnKvQqj2tXOw
3yzqkRROWwg5RhgeWAqzqj69+8A0VVxaa6DBSXUJ6kwR7mrrGzDrOENm4AeWUKNrDS0QGEzOJ+oF
1LTN1pewl15ra1vInuwaye80Lh5el+m1BHd+gYpjXJLOEtucaJ9PwOQroipCkhgz7MOSSKeWPmuN
bXu26lyaSl6sp/D09v8zkRUJVaSOAJM7XJx4vKN9zyMSPpiSbSQoMi7SyulsskAMq6xerCFEwkcS
tBAWoY7W9YcBvmGe3iE9tqxJlojp13BDv283SS4BAHMq2wjZAA8IciM5R+reHyP31jSziUxbGQ9h
PrWYxrfdM69BHz1R/N3sA7w3r0Mk4bc7ooa2I/aRHcgNCmhLJlERs0v88GX93bjO9bZf1SuHFgsT
BKAl12SF+qHUDnPj1hPBNqGTkD1SqAm8KwLO2katXwuyOmXeFsky+TEG/v67BkvKAO+FjA7kTAPF
kEPP0gZNDy5U9YdpDOBn1/WtAedjDnhGmPtInuovTlEfDzNLLBABOVUJPYoMQ7GtMThe/N4qWAP9
6Jo0yupxLoolu/7QFmfv2PYwKjnHzI2Cb+fLIAjPhTbV94fDmzYkdIYxqGqSUpv944ORC/RR3Eif
S4SN8nG5WY4EFDEDu5HvN5HF6gK2lEnOhJkfr3CCdUPc7k31Dv6mJJXbNTjRdC2vFmFlo+uF5XPw
vgYvmlwQ5cYxYL/hc/m9NaBa5+KGQvp+XvILI6eG7zfjYPiDOOBEK6OJJDqrpjL6gm6qYucn6eCR
i/Gf1tEi8Me0Qhib7D8M+aqBBayOLyIXUJhBQb+dlvCgJZJV+OukgcztWxbpF+m4/s0G7EBR1qCA
Z8OGeWMyED+gsdVVRkUf8v4ziurNJ7FBNfV8ZD0kzG/cOIelHnKGDUpjj36gDDmPEP8tVP3hteAU
pW1Mvd+jV4RaYWtTHVuOSE3g7JOxd2BEfI7G4KFpJA4WqVaUNe8k9N1AYD3w/P+5tiI9ibZRhNfh
Zbhrk/jFI/5RtqX72YfjmHzXu/PliSfwX1dNtWgsL+BvyjJfu7MrI33HSb2ZhWZhpxO9y1ubn2Dh
G1XXMAewrOLTSJDWc1voU4JaSJ3YXdodcfF7svVU+jDV+nNhVn5xhxwD3c4ifS9S81K9Kl/vZTOC
kKRUJlmYG2aTFlcIIc9HSus3IW6jeaYP7mClBcVscNkjlolpAYNYhZUhYf7X3eTLE4G6FYDBUZTD
lhWfRpn70cCspU9Ruv+SUx/DoOsGcYUr3XxzmSkkVxhLjMJRSCwGkZxD5SEmRi9AQEF7+9hkEnRM
sx9FVO4+lP2irhkAes/Z3bC7L3wcopAn0G0Q8/Xx1dXtNTkj0GTDQbZFOenfWYWCLSbJ5E7DHQFj
VQFX0UKuyz8Hx5M1Z+r8kmhehVohdNBq1A5cDhJ4VnCGi7ELU6THIgdb6aQEeoyttyyE+Fn4a0CW
r8WtHP+YkyAd59Gs6/AhO9AVhEjL7VkKUBFBmwL0gUh5TzN+VyOd8v8hGi/UrEaILr3OTrXgXg2C
ACFeGUZ52kaHmgJlt7U5dZ3t6Zr9XucERuPjREFKDdJD1BeWjK5lsktQ5JhiIKGaAGuwBtTGJH2i
uKe9Q7qMKxR/++ps7FhV8wNnUXmSftO8zGN+d2bYW2kgaz6vfwqawL8bO6Idvk5YHs8aItyxQdCk
CDvVO9Y229JiUI6D7F+JAaiBLuFqmvNKZn53GeQiISk94pcNlLPLBr5MReZ0GsmEMuUYXn6MwJZA
KUH8yzrwk+Z7uNhmAkbxZ+qH0ssjs4S56OOVvuP6tDauzrGYAq2hzmMOwICx/ncXTJL19IdjLJ8J
4ewCbfQGPGu1YbOgJWHYKS8/IwsdsuWcQQevVJxtTk2tzSrZftyNkLyVh6FcjtBhwTQcuVzuU3qw
13pnGzsHzdOt6uKBmbYcoxXW9/doQCsJaMPOvyvfE1ImFGDrMIlQ8kY9Ty47w3QJqUwfHgJxBWEZ
Rm/0q/rzxnAnJ7SshGVCxeqhVtLgmJqSeSv3N3+3q/JYZ9cGUWX8o4yQ5DwOkPywB29cMp3E+9Mm
5qvammmJRCsxDX5ptfxSq3Z1hjOP/FSgLph1SRbkxN/W0pXFvohyBToDnkWVdYPCbXeiWe6BTbpm
uKln57XMbHF/1cY3WJAIbtNn689wxBwm8T+kNmePQT5FRiYugk4lTPQuh3qOGHQHTIeCIZXplDHZ
Rjf2iFhAn0ucPuuuVy7V94bdV7WVBkFnxyDT/RhvpUjdRvAecFf3MyV1RLyi3QgipOKP16YnlUby
1lAN83440VJoNoztmvPSt+1ErubaiUPuRBsj5r25Y4YfetnnMy1H9IpQToPEmnxRgLM1h4ilKFSn
o0nD+0rXsaAjV+r0u8O6d1H+1F4/vLZnURxZQxOyMZKJ6PhLsCwSR6cw0FWiFc17ojAWjY2ETyQ2
VPxjVrzIIpBwG37Y8GCV7Rvlks1hlKKn0t/S2tciQTmpWaWZw4NMcwBjIy0Lrw34PKMFH5d6Wcdm
jbGFiKDgXesSbs+nEgmR+6o5zB6+LxE6dX1zFskIYyxSOnqDuCH8OjYLo+Ngn0//6oD3c+O4Jxc1
J7/wq3kPEk4z+Drvf7vKcwMOj9wNMk6j/YNUWYz+7W1AMIf8wvXKWeoFawYugk4vi5guoufthSOd
wdxCTAD4e4YL73M1lrEvszpAZ1dfV8FzW84pi5bTiuYhlTWV9kTsiEheL+eoTJeivQ8dS0c5A7C9
855vOL3assG4TDyJUosVlPEFCa5c9kjdXk0ycoGa6dsDThIufMqiC7M8YvuFXLxkCqE2u/V+z//F
gRX/KMPfdrxugk3V/vPHSGyjCcpRdE2G9iNeSbqJZcKuXBMUssWLvAoGTnCPnKwu6dnI3zzuDUTO
HqdEneYonz+qG1Ifp+R4LHrB0bIS5cJzU2uYNwn0nQ+XmcHLzdnNB9aydMw83s1qNQ5xmwneV/ka
zz7j6FWQZPN/sZyIhIpKTAzOaamLYQ5yLUMAc5O/+A6lXw9QQWkDH0kg+JOF8IxXGz/TFLWF6uyP
67Rx9N5zOcC/VJRbii/z/9rAgAOHMOmQbXTdeGYYprccyyySYbLyZusG3gLbWVzTD3AEgPoXEOyN
W+ycw3+QMnQuCrzce9/GhSLS1a6kDaNoZaCmsxVyOAQz4PA6SFJDp9XB1goAwxl6yKbr50gTwquS
xVDC1C/5D/8APp0nmlM4DnQmAafy+ANdSBYOW/dKY0tMbNGFEpROIxsYWwygOxDJgNmf8w1N3IK+
H65GVf6E/xp21/GH767PNIdxucVKElWTRGvAq2f/QmveWHXFLX6zPk95L1xG5+9Idf/91vR22svK
xJ5ijOFsdkfyd7EYg8n4NMNc55vmsyDsuW/Solby9YcP4a389oG0zk3P3WZZNm07EpRXy3c7+TXQ
mYdb6oPmuTr6BMB2pFeikqOWZMNrfFjLwjGpZ3NSqGiWFf+UrplzCvtbOwKftvdMVMX4SNb1xRQd
IQti0BTFbAmi9Cf+RSWakly221Af9QfRPp4+6pjfq6HK6eyiJwmC7ugNvVazf+dMHHOMNS9AARul
kE+Fvc2JAYMWUJ5TG/VnFn+os9jrnafBVjYhWjvE5G6zJ74t+er8Hdfb/CfgKt2f2o+Y6GRDUQfe
1ZO4bhLJb5TCe4WjMGjcHXcqgrRHCbM6d5dvtdMpwfubm0BQnqc6+yhlUdLmOckHJChWYJjEllb+
4waMMYPuLaYn+AltzMwLie3R5S1KLiryP2RIcWoIc7YiyUxyiKa7fxN3Cm1myPO42NdX8VLdksRy
cgqxDonCO252Z8t7DnVTbOQZjvqDbTUw9pLdSRpqk6SUxY+veRxwER1trMGAPH4njDwYH4MsvZ3P
sIAcnpkjVzodukMDujOOBAMPrbuMKvYBxrmcfF1w/D99i9OPQ2kkux3CK1DnFb4IXF3YUA/6481R
CiNw0/ltyiKDSzyQO1vd+DGGMjGDeV3L8hD21SpHUS3HHTOTg6mc+MHkMedaH7M9+6qzgLb+WLRS
iQMqX9MVkUXaHvSuXsfMCOMgysVjaK2A8v8VB9mgEJoF0RVh1Hhe+Q+MtUK3Yn4VqrAsb0T2KmV+
kJBJM7LoMr/FvvouGObgp2u5XivM2qc2MluFDg7RefEdQIaZnOTfirn75IV/d84jIA6nmnpylB+D
KjQDUQZETEb031/o8AHPqoPvQ0PSzQgXBgo0WG/NhOwv33HkQnssNL5VTC+A5FnHt3UNxWSWwNsr
q/yXnSzboFxwjSX0wLRAVzUtgEReDD0gpobIafigbXy6/ZXTypd5PkdG/TZPHEIWCSH43ZSPICcN
UXpSYJ2YcvwnZ2O66BV9TapCEj4jI2ULZmeKEbQfxBD1jrLoYtdi2U9Tfw5yZ3gEbOr14eyQKFB7
BQsYHeZTgnY8OnvfD2FugWAIk7SDYMs7j7rWcX7f/sBmEh00i4Fcythtv7VF586pq5S6kMoujlVs
HATupkE1Kv7jjaV+c//7EIVnWCtaryjMH8H1RcFLRaOsQLD6eGEKkU/8pl10IqQVbxkWkVWCse2j
UHwkTYzVVELkF00+7iF20IADmXBxg5tayDG4lzfdiwGeYsJ4rDe+Ab3jO9zbAOgwn6P5ocTmkHGw
4n/UL0WGBeO63e3p0wsI54/Fn41vJHHOhtWj9J4jq4RKpdmUv6ZAcnSu/nGB1x5i5uoCEwM1JH2i
dPXx/11TtBl59g/TVFhgl9zXcI++ujPI39cbF5s4v6CN0u5K/1zcWgE0YWqnKZf+BN+hBa2g6qSm
r5yRJfjcYG0XtQbAU+54eVjTnwya3kNHhBdoaLq2vmvTlTlV5hHjgRVGbu8anPkUw9f0Vc5w5UT6
n8yfgGMktDahowYOdveqWQUq3q9/1Um8Bz7txSh1RPs1Xi5/39Ny6KYQEigRd4mTwsSvG3PCp+AE
mbETzvZa0sgxVBtQjC6UtjUVifB/ICGe9LuD6Fupfus2+JGh5IlDa1RKCXeQ+NDyiABd6sp+sGrJ
FS2RXIbXY8w1l8rn9pkCJ4vztGaxZ/t8lwVpC666mKQrxTlR7YccnnGk5deO9fr20RbFfp8RyoSs
kUPEMLsN03IUNh64IzyiRD4fwcIfL8VrRe26cKsQXjREoATQ3IlN5AfcffkM4qK2pXv1vKRF6VJ3
tc/bxVJyGZqTDmvlgr9gYe3qNyTBqKQBLZwqszdLxEjTIJZ8HGxbKpx2TtEvMsOd8/3ny36k7oDR
2tNda3Mhz627czENBq9hCgWgnI+iyi5XCEWlaTAkBZ5LQ7iOdXbvNpDj1BA2sGFV098AvkmIpGYc
a1jkaugFvLWKxxU/u2iQxi8YcChBAVZv311NYQNV86nySlxC5QAfgjCJDzVWQT8ysDM84tCAjwvs
/5CSKGXKmEn6/EXSmqM+Buzq2QwGMA/rMbT+4yoZvX7HY8UuoGTWwurxRAPs9u/pZlt0/hZ5euom
E6j++j3gNlZYxfrYvVr8eFvKVyVcdqVMdzlUZ/KPAzWygFUBJ42J7nZyXH9KN9MzCPtmMhtypRZg
rCUvxxZuRL1QtwWxqbeXrJO7MThFZ83DNspw5B5MDoO4CeSCOXfVNwhsx522gFR3PZdB8xqzTs19
pa6ql6kGCCQjwCtvTMvoos9+lPWcEWOKkua2ndvjVHqQ+m/d/ZJ/jO9OveAcPX7Rmlxq3rnDYyDc
S8ApD9zC9/5hTHhr+z5UPrUM4tspJQvtl31COC/L+banl2vdO8EWF6L8ihLTDuqn2ZZEa3G1BiHU
dKD3nho/1gak6jkBAt8QK3O12VVr1Gzc5KWHnedRQ6aZTlNywRGwSnTS457TO15mCDfiti1ouRF3
xJQAITOzpc6P7fxKDtuvQpllNPLKLPjyTZi8qL9CWBdMecm7WrKL1gM+BauCPFeWn/Bza56g8CFY
LMTuiS7uV8T/w6Vhcu0V2Dm75HDb3NroRx7CFfMc2fNYn4ttx57czejyi16FlTSL9moQWqXRPE/R
Otg/tpBX/J5GcaT6c76cZYeMWZJ/pj5j919ga8OvLSs3yJtFIZPOocb27SEZ2m9E1E5KSxuEDHdQ
vrocv4Gikb9/PVBVcND9aCOjavgj61KQfKSkgQmzyc/uMUU5uVwOYJb7G1SNFBqxT/tWD7foSdPT
5nSnTSN/befNteVT23WPXOTj6vzovHRwYWPSfD9IPPdxLlk9o8XEmQUoAnasiRPzfVl/DQQkg6ZP
4GvlMLZoUpz2B4aAhx/Ui2AA7EBkmtH8iCCKFyKGMFJwdq7ahuEX4mVQJ0EXgrW/ZmWW50DSILEh
tBQ/TiMGrSRo5NK8NIRS4X33VahdlzJMujktezLLUbpbcktjHqRYZQoLgzH0BBM7KMMbE7sUSmLS
KSK8uVCv5aglUEK02gu2DTA/qG4eEfeSMq/EXsiBURke4HpF1MCo9MddG4ZCRaZcPqQ3Tbp9Nlqc
ZJE6HF+Q9XlTW980TH54A1zvxrkkGDZvT1YM6sfGsl+/gO2ErRmkYktb/TP77+nEON9BIwav6ZAu
NS2h6wZroj6NzBV2mfiPUgCU2567pjWI8LC308+9lAT1UC42qEYN8ds3W49M1ISvlYGbZAUGDtU3
Lae9V7tmsJMC7rVTTh/pMxIi/2C65W30el10yVGVILhmUW+uVOr6XliOSgBSZxmBOF6AuRf+IIfb
AZDB76ziAhJhCStyu2Tue0VSOAn/WDq8cKIrGGh7TxfkXgTsL+qLl7SiZsHyM8T24YKniH0Mru7Q
tbKLRs5eoUXdKN0I+RwofST6/DJvW8AcMG3Z+cbQM2qH1UiXTUtc39T+G1QHsJO4BMQbhSwT1saZ
wMhRgaog3Sk2ZK4hYYVuOsBCBKhsN+hFYgtTQsbKo7bDYTy6/M/QcaM8DT19y1zBT/E6a9DV1ya6
u+wL9959/GNk9dUpeCksmTGSlh2xmh5wQlozCU7t7sRADbBG6oQrPW3s0ZecYbhC+4xgz+loTeIC
gartZDr9vSe033pzVqQ19fg1ed5xnxuD3kuqQGPItABzO9No8FIS9UQ/t59t8n4DvrpDwvt+TGZR
pHoCzcd0mdAVdj5cqL8wWt0NMwnq6NFgx3qIMkdWi3aU1kVacd7jykt3deoANBQZaNfJAkXtE2L6
Qouz7YdThOrt+mf+jKxNv/6vhFJ01GYnQ5x5GLVfZgDTnObSm5+BhCU/5AaPcTfhJ/qhDCjmqYMp
rCU0OOmOpH0/9MnfXXnk1+humz4hjbgusc8Zl6ETSWNrEY62qQTvtitCgvup3rPaxQcSC1CCaTjh
0Ar7ACAIDi9aDZu7eGErtIdBxJ1WlFDSJLCsEQMP5qWQvHFcjbcQEM2ceVzyD0EmBX8jmlW926Fx
dQsSWubVIHlOoPLJVNM7kD/HrlagqdsWtY2t8eBcQTO8KW77spboiIbh6MZSPVTX4zvien8h0q6/
0cSwUVQaZHTEJpX1J/9GloYN35j7NAf0I81TFI/nh9B/ClZPa6GArXaooyTp69rx+gZ64yrEYeXy
FbJrhDgFSiHftVXaIaBBGYzNHKCLBcBxfikrStVt8+iWo6DdTag0Iu1bagXqocQcitKQ2RmHfCc5
zXrGQ6jJl8Zq3k2QOhtSjiBceZBbGha1MBJV1QFw7kKrcSvsscTtrGBEe+UVhF6pQHaJo78czdVr
lEwLd33GwWaogCqDCUb2reFhqlbS8Afe1GXTDdfwdPKI3rGfFQ/mAFdfNYjhLwrQ8NmfVBgf5P+K
vCbdc6D4a/RN6/6JWAVXZTLy2flnPJScueP6MKQslytohKadQGBVB4OERBp/FZ4eSX9gO+stZgkf
fiNHbBe/ZV/dwIwie+Ll0uT8jM7p3QUD5A+hMtF39yk96L7n4hZ+3flznsIhILDjUcQxQH05LRPN
NLL8O2kUp88d4vslInkAvsH6PefPHw7fXhWggRZ6KndgRnnSH6w8QooVDwJtxl+gVncRiXWmCqoz
G3fhh3FoxHuctHj3zdAc9Cow60FRvpg9mEjXtxkxLfOBpAe2YEJWBztKIAud+D8lJKFu/hGdNSHG
YDygD6KafqqvQlxMGp1IiYpnvACrmIq8KGS8hqhxgE1FeG+uHrNculZVS4vieHF/dvw0IkGZDtnq
DtyeL8RI26SRcVEr2i2gBTmzkXMuSH6e9SMnoLnvQWllC/8CjzFak+rtT6p8NFL/eFzD7johrna+
iuj3c5LQaRO7oeTbWqz50SJ5F8vBoH3fnFrM4z0QXmz2TbqIfCO2yoVxq6K2cNlFjgVM8xATUoS9
q0xR/huJFTG4irU8REEjXtfBIemGJ6ZqvlwuFlgSG5reSs6doHtJjVSATu6zWDhAKWAYr3mlslRE
pbkfUQXr0lnFrD2F+5WEw5Nv12sFgeLvutEdz1gM+vy3XWQrLpPi42A2I51Tac/MieRGW90cnkFf
xUTBS9GoTabHsj3K1UDpXZQzgwA034RvDopCzeZvSrcAtIK3sz3sGDjQBRcphc8zqT7wkudYvYfH
t3YdC1ZY+yCG17KsoM1vCapIDng91t75bSpCsHmSfixBkQugxZKwcoiubPnvqK/bdRFzMxmesQjA
nhAkeZ5afT6v+9BfZNvn5pxkW68HyLrk8pheXM992DaFWjjYZ0Y77btP/olniiYQhuSFqXgPf4YG
vgSo2QwDFhDRwemGTOSb7Iug9EVHswYZpP/CN1HrIS6NsoFxoCz+MW3HjMf8xMDHJSdpRBByGDFX
Awr8FhAIZKYN2SjPxL6oB7tdvdVkVsDHh52NLEkOu6Yqjt+dU+kE6W5nAj34H5JZglXkClf1vFKi
dG3wvnnB7v800OWC+c9KROBZXuHpk1a7eZBZ17QlENRLr59FPo4HykU/EdhhgwRSdbLbl9vZoDJ3
3A5x6Gw2r8KfJG3d+qukVfD443sXaIjdm4HlSeGeGHLYsHsKPm4HN4bkKcMfx1t5M7hGxPiozY0i
G3u1iUQphw7WKurYmdvmMs6qavvwAe5dmfG3g2sEuZybJx2Hyva6smDcmEOiiQ7e5mU/HJV/0i4T
TYgUxDYRprvXv97l9Zdv+ib9rxxE+Pm52+vskAfF+AswsTjxkYMomkA1ES+XqD5TNNINzE/kiYeE
ot93Bwky0JtRlhlafrf+K8NLwZK0s3k3frt4Pma/JHWy79gRXzQF41Igu7697j7lfhpKCL4AfxBV
VhfYQp0tqNeERv9hT/3LYVDM0ce5nvCJT+gvVdULGablwFWd7BKgAYF+pnZzHRJk92BYGXSpdbrh
TwDXS2tG1pMXi9GOuj0XQDWHwg7DQEL3D/x6jPHNw9MDvy68sMTkF1dvr7/BR2jwLLBBcZNr1Zvb
/iKlxR3Vse+Xk8t+8XmjAe954KwumnJf04E071eku/9bwq9dtfR1z3VIZRSlSLRfRBPa3C2q4/TN
yhhKmh2bRcEalO+xnyWOhdJXEWZGP3LLvOrrn09/6UAot6FtLPl/5fF4VHLLKfaAJ1vIT3gVuME0
dXDc/NMdBwgcE03w5Esqx4lHb/Ckegfxa8xktZ9iDOpBmyVnxrUT61K46WSaD4NSlXxhaWh6W4dw
0KIq019xUnlDyQIn34uCK1Ax+C6UOlSix5Z0PuSMg/noHpO9d/URzZoucYRmDmuINLlAF4T22LVl
0PwK/SQB4HR0V3V4cUdQ7rBm9MvXSbFSLNlsm0LDCz8+oZUN8vs5bXqLIrPVoNfoeemYvahfrqa7
FDGc6UZvl6AdLM9PHFwmi6NF3Ii7jbFZZ7nh6Yus53JVJtVOuu2QeOp/KGm8oR7n5bydXNuCVVwm
l5ufNXtBSWxi3+WWcG5A739hnOXu0j5Hl6IkxyygrxBubRyLfQk5wXNDLGR+G/RVEQKkHaQzM6yq
FjjTLgRWF+NwHgX5j2hZDNVF0ReY3ffuKbJJ8Lnp0AzpaHXgUd26hAjfKydUbNT2aWpIYjCjCcTs
VQpUglJ7AZyENFGCFTg8BDLWphaMoZ0fyv1UjnQZOrbr95sgUD7isAP+9qifCNjW9l2ZLuaOwlVQ
8d9+YeyoqzXza6+7GxdKhMiHxQ3E2HNL6JE+5ZlEI9FLFo4apIycpb3A/8kA3YIchJLZyCRUOgEi
QWhM4VJNyLWdBJApEZXzspsS7U77aUQNdepn2/7/F742l778KsjuZvoPSa5bRuTvqByttT0DkE6d
B81EVygu9EP7V4vJCzudod0EPP3SovgV1ALmOSaDreOJ/SoXrCNEQbjGlhSp1jrVyAKCl0mr1e02
g4g7rezrRIBYbpoy5TsFXETTqv3vArouPUu4xU3tznmtO3Jhx4d3EALwi4k7/rqDUtfUcNoPOdat
Qo0i/yrHWCX51/V6GHJDPeLJap7hlu6xLH46GZQ5EoFn12BkYUfxuFJcgz9VothA5+PLZbVjX5qA
yPjx7RlCCXgIsp8eveb6Kw5656LEFXwLR+KbwdquR7LAyzXl3K6AuHrOwdRFYsr8uD48kftwcZNT
qbwYLz7s3/mh6LYJLvjjLB8yL11MKLgFJWQfWb21aoCxyZaR+13hdwYqG9S8lNDrzaO8ZBOJ9Rin
caJ/jACkXFTlyhtO3lRCS/ZaZPufXsNl8qWM4wj/M8sLxGF1t8lQiZUThq1kZEVoLIwqE6NuyJb3
QHmRgcNIQwaMlFD3BclSeuyf7D620eqkEkBzpOJA0KSHLOPNkXpgAu2/A/shEqhi83nfexH2wwyq
nPBfo2kq2sBt9Ids079L3tlkRb1BTjqSj0Mm39TffUQSItPgsk/5m6UuQO8CPl0fCgETiHk+UY2B
e9gpwUzGiQcr2aMUfibjEYQl23vMZnIHdoXHdpy6f7h8OXhPRppHmKjuu3RMT8NlG7/flItXJzN2
yq8Gs2vJGi6NmhlAWMKadFNjapLVx8Bd4qduF+rHOCDBIiwu8kspAACFaJ4XUtRt3rzK3JaPPJlT
DcUSFHKae2Jm/6UzpvPRJF79G0jrTmLd6SJhAomL1n0FzWdp8BaogkpSKv624jssPLtKaGtI/GHG
TU4ngE1kuze4wykDZgtUlivhWSo/94IXmW+cBVo+VeCmx3IPUPZ7Z1GLwAgeSJMMRaYZEA4kR8ha
B3Z1q6Ytd+0ayuifIGnAjR/FA8KZz0q9OH6kqkd+AG/q294TbrNaVkk34QQG60kjW1gIFYUrc23v
PsHPl4TxML+rrrQvaqBIwL+JNL1LmgOr7PUYsSWo3PbfcfL5bWdCZTXFKzR3wh9dRsC/JQsajcwt
tOaA5wN5nXNLA2IIg+KLJxFusDkiUsKiz8tJIk3zMnmmV54cpEGxYLeGwFhv7P3Mc96Z450JVpRU
R/YROPaim8PrEajQl+FO8SeuHzAaDIb2PC7LdQc40Q9IPT3Dj03PeDXYoGF+gaYW/qvCVPG1LmC9
prNuc17dJbtGOclOYoqhaAdn6Dy/MRFIpb/x6Z5LavGl9WVBcBEsMxSvtep+78Xi38YoH1jGlP/I
kKNLVoEekoXnDXA/3yHjx49E4pH+AH3Gi17rm4oladobDJXBdKBpAzMlXPEXBZ5F8a07xvdYChzq
HF+RvW2LvG7GnjrtV2toIA9LCuRPJUJIH48CWSCunm++W/U1PH2xCXZsY8G1CsZuPIpPqoZqnct+
UXOsxi7mU3go0Db6PXMYOnS/oHR/muO2ZSwOmcDvoPIqljvT/J8z4+Wcn+uWV63en+AJrWjwNYHa
iOby50XiVtcTOSAnCzQ8ET4uAsJ7h00qZJdBe6MRwGY/Jfv3atuZLsS+bB4Iz20ktR0PkXGlvs5l
03vg/mUReiLeIe7sDlWKETvlvYpr+2EBtPrHyljbSTa6K2MPWSSOCHQH+4jTUDKWKjyMF1xC7vm+
Q7esES8ZFbBhP31vzxI5M2yy3Fu6ldQzUA98Ozii3MMBK4kRlzoFKouB75mN0gSOslpWLSyN6f5x
GnqB/qU6yoegnDyuDNRo4aIQrTmOLLdQ2XK9uB0zLgnJtLntoEslPP7WidBI8k8wi/eWHja8A3w+
A5bFzKaMXIfIpyDN5VH+1d8kImmlFx+X7d9xbHvXftHaMPEgXmHgsqom1rrbF5XwBA6YuKUL7Qnk
chwixmzzuUMhxWeDDG0FNZ6zNbURi7p06F84EeLqsSWWEZ7HrxHSUYSz+MyuT/MwAJfUftOK3Nmu
WQYGi0hY66TzgSe/NyDje5BKnO5s4lR7Dv80hlM+P2xKRwowDEFnLcO4xDzR1HIOfBlSXnUE+OkC
cbadxRLcZKP0fmNv2IsnwHnElFMHLO6SOvcds4g6/YgLFT38I3BiF6kcnl/so3KXASm5wch3uNYn
huhuLMCoSl/Wpo2zw95POEuxbvxi3Oq/3WzZQg9pYOGhBBcp/gj+VC1QZ4/xQgPZ9O+3qdyizM1d
rV7IcAokBCeKT8hLCK9CIWWjlh2fJHRyOGT4ulI4PkgVqLEXV+q94HS4CoJeUDql9t+2fgWYA9Iw
skzRh+hKF7n2kDyzXaaddmv7+6uoHRdDJGPOOr/u2hMSFyqqfi/PEGREN29DYODKNU2UxMrnP/20
247nbTjF2PBw+RCH+PXhvr5X3eL6cBbtS4obbuwNi0ZIbXZOhIzZZE7qJoKVuJqojvaYEtI6IMmT
oAVNGjnt4XUGzQG2BdAmb4GzrIV8D8SRDE2+mH5A8/UQ91584oDIKUcX7J2NtKzf9eI9phTgsXk6
eOdWqmmoqDwSLSWK9WkadMNb4JLO9NiToBxNSKRUlREWJkgam5dDWjrbnIOrd6rtWKBNbJ+ydDMf
XOgEhHtIzzSaXe8uH+cGNM8pYj+pYbQ2ak0ANZWlJWJF0UiDd8fq4CokF+ClXnVKJZh9SFdu+yK1
ZtOo2g2gACqVGEZrR5JuerYcjzRoGLuWvgIchRYg/3faxN7mbxe2XyoM/+fkSXlfG5wXo369DZm8
/frhyFCSeCxti60PJaR5bDiPa0PGzSE3JCj40qA7jH+x8yOEvXisLaCvwBbiZ7mE/dLIgUASjTXL
Emulg4qYdRfIIZcg+LmtBGKdv6qajP60iSBq8g7mN0VZr7fEtEUXVT1jgcRxqnpiDJUC0/Q3qFBF
9dyom8XW7a+TlZoyMFh2Er8uMUSHf9j8Aw4gc9gWlPYDdq/TOOHTo2UpQo6Ay1pPCglJgpQ/IeDn
89Adh0P1ReWRNNHbB14RQ+txcFHlhcTCdSL+5LgIX/cAcLXn+cPleUxgy4ssmG29kKB63BaQfnsd
3zWvqh98jZ3uvrbYU3cTcEY6P9bA3hBzVVdkjKfdZcVRTB0PG6DGMXHeL5i9Xjwz7jwk8vRNYWqn
RQDfLtSgRjmt26COPqLnmVtEg9YMNYyuIzS8TWJk6XimA4RYvfzJSBHA59mAaV9hKzZMLFxz1XhD
Gai38MNo4W7qRQrk+L/NTkO3Df557SqyxuC1SUFwB4SxaPwPquMUnluC1svNBe5n50jSlnv/wpaK
ef7BdU9C+Fqujqqz0xHZGQ8ewGIUA6KQH18tKCah4Xc8md5bLg1nKqcku8xQ6ZV7KuzKxogSfVRb
Ai9O2+EfCxhGPJRLWRhXq91U1KHG2jldN3XTQW2mVJKH75NL89SKgq0/DmYsXcBTpw8z0arK0pZ3
n6c4rdIT5WTek6BCrAwF3XY7K2oTotks/pVJ3CpoQmmZtw6CgwZ4wzXcJHi7wbJ9fl18M3E4AcrO
6r6pN2gTCD298IcbjJa0Uakw4C57FXAOWMledgGLo9ZoInx2em2mqom4+OVXy9bhrptw4Nx1KcVS
MqbNS+Te4/8i85iA6tQIJ/IaNiqfBx/LLCYM01wbTd1GZ+qiOazUahA0Gb4m6ukXmuPcI9VUHyI8
8/V5GQXbsjlxWMNFGDuqIRdZrxh4jXCc/lnXx6yZTYKNz04Kj7pKRqieQV6sjYCZVTRu0N+2+WlL
YhaeJDD0nUfN2MuZVB6nriPcNl+05/h3PkNKWncEXvDl2e5qzRDOrByBMVtPLUn4mPmWe5GZClWI
hzjBp9tw85ov06Iz3ErE3yjDouiQgbOZbhwLjnw4lEnIm17xhEF26ISVGkzRXpmy3mEy+TeVO9zE
8NNl7Pdc6V8bAIR04pl9+SVXZgAu9vGL6Q1w+BdjpJmx2u+QPuM98SsdgJe1llMQbm7H3uIQXLim
OcGB2v22vGFmrxUq1TwT+QuU4dvrliENwQCriihpeO8IoyG/a+hxixyDWFZfQg6CopbcHjaCL3IN
ZJwhvQ/uQFv2KKnYgrrrMp7fOd4HXcbfvhHFBOxsFicBWYSHLX/S+L75Zk+MGBEzxEvIAWFabikg
vEQq6wOmsyG91uds3TLU7HI7qGomJChOmT8bsoWD5BBE3Qs4XdySXObXiPuIEcoW6tvxf9+gd9um
XZyrUP2L1UNfc2Hv9xCBkSGWlWOV+bSh09swa9MckVJu2UGRUrz4zlub/4HfdfDzVe5iN83G/6I5
/mjLiVaRQjccQN5/0yI27M74kcdJG8xJylUe53Zxe4pTxBWqKi4x55c1NpsWq6VukF/UVWKULb3e
ggN9akkVERucEPs4Lve27TwaKUtc7df56AyzzlFlJnMxV56r73QYy2vFMc3/ywam1Jyj5lEql2oy
B4RRInkjtNCnWVyCrPNChoyg87keW35h3hXdNzxkLAb1pn0ZrkSXLXDgK8Zi1yrCmdwM5LBNlbCy
pDBL/p12cNYbxlqjdiNKJTs63k6xgfUbjKPLmHqI08auhbPJQfvzqa+4RC9NfykkcQCJLZ/zyJT0
muPahTTs7meFTHDyMybgPhlEzp6Ve8aBIiFxewM6w7rCLa3grjWCwlyivvbi8ACqQWKp629trCoR
fBHAvQH2uuZPA18cEvAIKdYZqAZpMm1AsfZFn3ozZ/pSbFc+xsHVtM3ygT4fasNOzOaIRU2L4g1W
fjPj2gP7JZVyP+tEXGr2nHgCNezTJz4/nm04gk+v5kWRDNbqSSoYq8PlbYvPj+yH0ZAuSQo6v+sZ
JVIX0NJMVOOZlpd4dwupdl69DUgX5at7fekZmW23zCNH7vm+BlOsyEf6xJufiyyHBZfoTlXBVgRY
5kpK/HEd+bfG2gNQT5E/oNRL7mflhmZKJndXAWdmWSqgw1+R7HhWJ9h2DhheEHMsJVYvL5gn6eKq
YOHxTqjyMDQ92S5CfnGHAQwy582TRDMrdO7MLGoFbYqD2E+ybI0KDvrC/NrZOjGGbqQuJEMuww2p
ymsvHjydkrdrDHWRynj2Ga+FXWRi5NcJ1b3bEv7EKSoLD+SdRTDodTTRYdplM2aOOSFK/N6fEUo7
7gT/uyNCgjmoe5EsG+yD18HWpKf0WG+Wx7bl/fsZamBaBqyDWso2UkURuw6MeaLUHCT4qOJIKY9Y
LgAdjZRZk5/iZXBuW+0Y+sovzHRzBoOYFDQ1G6MSiifhDxrEUyB9/4WIn4fkKqBEsYqF35d6qLom
X/ho7yXvV8gpd3S0x0Bm03nAfpFHwc03kaY1FZOHji+3Doo/UYNbQThZrH6ZrFJRwcDmCK3gDX+P
qN2UBIHlTxwaKP0j823srTnFjF+bDpocYLHarSVGAAxajFibM4qTNDvgUOk+1/ogHpEhu7PLOtXx
GuxPyySvrVOWny4sF78VhMj/3+JCvdoDPpF8S4dswfYD/Ti+KAbwhVOtLkOVYya17sZxebmhhgdJ
VcE2nDmBi0xBd+11meZRQkfHuzslUfoyYPZv/lrLKML68eT78Sc015BOT9JGVRUl8XzYulijnwi5
dXp1d0p+V4cOCPGWSkof+syVmeGk5qHeUQNgzygREO3XiNnBFD8jGfwlCGQWIoXuclAYclaCJge4
MAzfm1Ie4IDqN9k/uACCsO2unKxnOLZOkfPxNdkaNtsmQRo0MEfuA7EOsXuPN+qKUmmR+c9Wm1Yf
hHjF9nFjQpVpOTv880z07VA0Ou/jGX/1N7MKlNL5E63Sd6u0EbcF83GMm7xOF+NtQjXocPMykQ0I
79BZQWHe3YXdQaPk0OCWah6BdBRQImxdVWVO7JrtaqfCm0T0Oh+uMffeyds7EPjHCAsKJb8qgw7I
0tIO48Uuq89PoTJDDeClzOPjg0RdLR3X0WVbylLg+X1Ky6uwQapxi4lO8XPqZlTI+s/eHtKwnmmr
pOKezGOXa6QnTpAc2j3ETkVtE8R/t0XhTXUJUco2V1ygZM2T534QYoi8Xq9rwPBqEyHRxlQqDTwP
l05oYmTrDGOu0M2ur4kXISAxgpg6dIpWYmJeSfgFPJXkV3ejT7haRsKaeGPQ9+vPUmvGa8Te0Qr3
8vLSGr4QPlM/vI2Ot7oHe9t83GCIc8hXZrVDhcG3lsNsFu2aFKulGcOAWlZ2Tn+Ivv1UGOn0fhQQ
FrP7/srfJu7J/6EcH+pUiqZmx9t4ob0adfZNZlBJKZyD4VB/MM7n01Xu5TEQHsTDzVKyK5UO8aKD
JtF6F6KgW/pXn6B9WglFkklRF5vPqUssUY2V3om7FqaZKXSfi61t6iKvsgFa9VJEmv3k0yOl9f17
fjNrtzMD61bI3ZVedVPQqcKwnRoJw+WvfOilHANfbxlxWo9cs3R9+7BaSeodSC1UcpEnsrpo1cMA
iswdjQmRB7geUMx/I7Ncneqn1o3Akj7epVHdl52nRspyQdDITB1PQYXH92jt3HxswXvY+YVzaAAU
JQuw9Ie+Azjdv6xY18Hhy+xTFYTwZe4V8wrOGcZE8P7X3WJi1YPVo1NfCADRKz3UB2S7EUzDXUZq
FhtDDT65CSmsdP630cns7QORPYQODP3mkA2p7SVxztliuIezS7iVu46GzRIIk+JOOCGPyf/71dnU
CLrpLkPjykq9nSO8psj3VZwtQpQOBIQ2oNF8E6krqfYjCJkls6NcKZTWWOwWVF5LZGJkiPihlNP1
unQ2l7G2/sx+DEKz9PphRNoZfhTYVFFKKF2o8AQPxRLcfPkOTbuLf4g/zyeJjXtqnVuiUL0DD9+b
cKX79kAPxSQEl7sRh9xHiHCZ/gOFeXDq2pw2T2CYRqflpFvmb0TMKJVUeL5lP2AmBLQ18b8bmz44
WkIpjw2VANbtsl6HBGIdGOWCcz5HCTBohi2fd2lkrxB//fVugE1Tngf0pcNV9IBLYmJSNu4gijC5
r4FG5g1sYlUDKOripYVLgUL4fIrga08y9pc3+6bYAnfOkWUnB+2AfeQqxT6ZKYCUQazV4Vxud+3L
pifnZnrZ2NLEpUTKGx43HvmXApeh2l9Y9ErLHZJSC9v3buDNBKlLwPku8x2W0ZsW8K+vYwtWt6G3
2XUJ+duqgBD8DpxtgKxUtCjaYtD7wP/O1tKcb39UT8lB9rbKvz7fg7ogxJZqt7Bwoqwg39So2ceM
v5c5gsJ5uMEHQ6wLaoL64Ht9QBQixVwnMDZB4IdwZRGB5ZcR+eAMeUQUG0YOQeMGpEjAizF/6uTa
L/uUORqAiAxUbgYTCD+EPhPA0TH2rIyaLfxvH2ExW8XEbOaG0cjcfX6WB5DCV4Hcz2glazHfQN3C
sdqA/lJsbM5djOuezOET+4eYc1Ef60i8yyrIYGN4iMuA85lFLAiIzbRF66wlc2trgCQfyzDWqnCZ
9v2TeVITwekUQVmi421XRypgEuuaq6bQPZsNelw599Qd5erOXwJylMaSaqONznljahbzAkIzTSbr
w8PgAIPq6J30cKFbPguPSuNAxVihOninfRIohE1Rdaj+bEu1iG2lD/3TyZGYfmg0qk3Dg2q6QkTC
+9d1Raa71h5zkix7cSN09x9E3+cChbX6jRwsovwiohR5Vv4Lssg5jV3woKVP7EZsnfscQTGJyKAF
VL5ln+OZYSSDQxLXre1ICPVZHdunPLpXIJfyD03s5Mx9T++MtiYVuTSSdZmn6MqfnK5j3qhGvfnb
O2mxuza3fnNDTYXdFJauh5tTU/iR2AVc+wzTt6JW0vPLnB9WQ+g4zkGoP0tNBn+UCkvGZsmfZ1fp
+wShQ1I5MjjuxN72j10rNW3HfxOGGZVsxKn2DEHAykUydaoWJo7IJdViXO4Nv0LsoaUKaoRdcDu/
AoeyQOSW4X6HKkXtMlOGqyab9oCPXKQa7x4KIeVoIK+vBZYRUM9Zv80V7sdzTEytujlRE1IPoSCE
cvgvNKJcwh5cTzLNVe1r5RNWG1hgujs0Wo/MlE11xACQAvNOpOUHQuNeqeDqexyA3YgEwnDvAzQf
Z7YUelXGzDEMRt8yRDSWoomK7jOyKx17+QHauK78lAL7+oo1IvFwOrM2odmePsj1EGL+VtdGD0OK
BQbOIpL1rdcuZihkSsIpcz1gP9LVltOLDik463+pYSEyejwrlvT8uwh6CK4RcW1dHXJuv+zQDFLK
AEYXGZ32+hdPbiDRGxKkosS/xrGN/XmotlL0zpbtTRS2upWd2rNenlDbZr5xPNMxMA9K/diXzCKw
IN2lKsElvXZBfCAC0htiRwbJh1bJ+bGr+7ojXSNIyJuT15BaftIngc1Y2jcQsQuaad4GitrXQVlT
aDvriOvIdi/Gcxp345jD7ohJIDbEchZCl0oKlUwpipSTF+DcCjAkVmph6oNrgmseQC+KBSydae07
AULLrTgkbd+/0H7p1Fvscc3rRYPjFBFYaMrZr+QcRSBMG66Xg4Iwj/Bt5eHzAWA+BbaAdRbupS/l
2/e8T6vd4Geebtw7qt9RMTRbV1ZreBR2sR4fvd46ipLXSvpSCUKLlJKJ5ljcld8QXRcbRcujnOYx
kESMhIGWy4R4lM31TnDUbIkCqJjXdF6xLwtgmZrQjip9laJxgk3gO2FLaU/GYCdkTqoJvHiBl6Rn
sx0Ns+qCtxXTORT/VACaZ9/VX1Zj0oRupCY0rudJIJqIxcd829dMCDte3o3npdNqoPcFpsgoJe4f
a4adHCjf/9pnn6w8J75c4q4L6CtYv8qERAtE9Wf/DZw4YKtG8fGLfWD4t1C3k7Rvb8xprKxNIPZv
bOXtbslm52lLgRnvdeqWuAKCpV11vbQRM4c5EsT7JmCgICfvk4BXY4CBU6NjJkUXSFjgtZfMfkSY
O6eIQurcNeRgXCWR5nLwyLJ21ZOhKmHlZweWKJnWzRPELmiiPNtDn9nFdscVOCehLi78+EmPrTFd
QGtSbOqEZ29S6LRhZD9ZItniKFs5NUPxhRKChH5nQahwjnT7uz4jwWyxHsmvizYg/m+C82ZlL64W
qYMG/ahAIRzifj4d5VF0AvHE9gydquiU/M2l6K40uxlcItYvPyx+zrJiuniayMc0jxo6eAS5mOAk
esFVYu4W+rAjAhl1PSWlLaHw891DCxZbb2BV5zN8TIoph9fWUZ4Und6prJAK7rLlvffDPbPxjN9g
EiFro7e66pZrULKsIZWUJ/2W0cmPukc0Hp9c/MDyeJ/Gwl+6STEk+mtrWXdO4kYkKc1XCR2y6FWG
B7rShAVsouadLvOo6WDWa5YLDr3wSv3mj9R5RZf8DDsHYqSGNbEXM4UCBcw48N1d5mW0hLbBUoQi
oJqbVzaHkqeolzfUCSElELK+jMT9+MDLox41FE2iR3MnC9A7UWE4EQ1yF4F32pbA1N8o8fCUK886
ougY6+LG6EcVnzBZ4r6Vs71he/xRQF5QnwWBfxOu6CDPqKf+t5/tm5fH+FyFVvGSBTalhFSxLhGp
YGE6PvsE7rwSfu77V+hdXABjW1qe7KUf7HI7c/aAmo3OfPGVjThOk5vret0ts9EOwefb+7wIWu64
jCCWVdfrB5oQE/X6XO1m714BphCQI/hQUM3C2VPYV/D6MhnXojWLT5m9BqfUYxsusYuEJZ9Pnpzw
aGOaXHteBKgtGytpkIh2+TTS6ZXk+VXwConM29ceQ926AK+nPS2VhEk+29AGUPLdUdLTZFoVrL+V
8FGmndB8pSgpbjTjBiXVqT6l2pDpTg9ksIjNTRrO7X4xbwhN6F8pHd/QXM4MqdS/atlWTOtgi9AS
gyXs1aKbhZ7FNnghL5G+YFts+bEETg+G9iIsDQkrg0AHCg7NV2r5X0eh8y+1OHLZge6Bn8FQrLhL
fYrizcBzlkzt5EVMjacRNpXe49YdDLpBM1H+sUJImjyBBypzMhB5yOmH1Qxm7Fau0c0/erUMAyAU
pX8FGoIiuRlOSUStGiaQ3sexNdxpLZsBn4//YQwllKmxbszODS50hXsPMsp5EQ6DCzMwvRmYHX/H
wBHao82Y2pImuW6QRmzSi7cm/js7ZbQKl+ZNbozbY1+Sum23EVogb+qgvu8CWxr5Q2ZPQF5eYEmM
CeT6Sp8PX6yS+43x+I3w46Oja4x0Ufo1Hb2m+y8niMWJbgwdmMA4QJbQCbZm8spQxSQDLF4RquMx
48dr35ELzCyi/nyxjGi78LFyl3iIwpK6+YSbP4/I7/vlge8PGKpv2ynKjNUxT10chOQAwWWTB/TU
5AGVnyLRnGcAGw49HqwiUU9sCYKtOevJslEKJcRMm7VWuID8e9pW9wvMZYJKBrF5s7GAnbAclxmk
iI09fyNNU5EPxHL3Ev3mUIj1whR1qScUD/ENMsH464bwEV2WWR+O/kgXUP1V4w6qil7/T/pDvptQ
WgvivktmkKyLCSO6+2+Uixl/n17Pcdo+CpL+m0tZ1xdMsE7Qrw1Me/tAARIVcJ9ds+Ar4YO2b0Uv
9CLSUaoCsnBgAV9XHOIvHtxDIHaMedJd4tLNVNQox6bGaoRVRreIYQgRj8Os5GjCJBWJfHS/EVog
Nvx2/Yvyn3In5kDxo1HjQ1teTznSiexCr/6OrAajsGgYqUEOYkfLO56mrpE4vqb8JtFFvwAqZSqD
HFgUaki7aUho/l+GTInlK7BHnVUvOgWYHYuS4XZpjxZSqiYYhwDMSbmAjqZUBCW2CuSsgpgij2kx
u+7UjGYY5PLXXr7BIyhBSEcpF37tmeLZAjQiHWV4EuSpl9jb9CfGGhmpgvme4CrOBoZ60t5aD+M3
nTCHC6jswgFibY6az1X4CrNeWkJKygbkPX6Vh1L8lzMh4zLROw/OZAFkhwbur3GCbip1btj7a+Jt
7z71WxXAoGVkjXPkkllEUyxZXglrrebnsj4ToypouqP9SOB481wA0zOyxvMZdTMybVrFINEyhRBU
yx/3bRjzaAK06CD3iDWTnwX6cpuEQnaIJCuPceBU0QcZuJQEyRPgkyoC6Ofs7HH1k3ZOEIVJIDMn
sqwDioJH9VzzBkIB0EbpYapUb9AEAjESpadjAYFQWXzWHDzD2lxeuI4nAScTfxNnBq0dwlvToiq5
K4TxnC4Clay2HcyGqerTo+j0VdM9aArklvmqWpMh85dXZ5DC2KZePyhWJhJq4ooL9aHQBMQu53nH
g/A8QJRjaaG9Ed44nIr57bJv8RPAoalCQh8ilfE8cUYAfSTx44fZh933jA6O4HQGkrVR0a+5NExz
LhmeD/MxP8ltXDc83c+dKrRJXXQCE34QctH0X/SEwhcysprsrPXTCrgab+9gDCTlLrP1gI37UkHj
2S+kL79Cgg1+cV0JNjUpGz+sd1pHTH10RLKLMqSqSFc8X2sAgQayNdqGdJkRSIoajgWNAqgQyTMk
O6OnBL+w3sIzPlfE3yilnNI4WrrzFHWjN3DVn0Kda5IFFKgIsWmQBPeo+FFjUtUukvcHOcZthJ7x
M9n7yGA0RzMPXzb7FlMkEh76SLv1Z2Xkvcze0K8U5Rwrah/Sf7LdIk2zYeHeDOyjixqo72RD7/JL
5OvYGu+oovTu4hjEtRUrxJa42dopSh2/E6H7OObH5XSIB2GwfXI150edDJfmW3u06Yl80ksXuDOT
GQQpu9RlgOa0ma0tZGWY+3Sz2U3njzM5x30UmIP7y+UHncq9nbkchUDT9Lpbh+Nw3R5Qh4gaO+1p
zkC3IsYNx/E5BfQjyxFdyDwPSIQGzcNR9vIPfUC3GNVxIRdQaYy2Ahn7rMgoBWSZpcUPCsoNwFcf
b/0ZNmVm3yaEfgIh3ymb1J2TREGkWY5bCpmh6apMvvIf1YJBaWx5sQfjE47J8aw/OjFdwCN8OPXG
v+p+7GDZULzx7SN5oiQuiPeR0aAKktsHGYIQ6+P7798761WfJh36ky/bX1yoGF2QbHooAyF2JTbw
hvbPnK7j5kaLB7rTAww8//LkomBBL1woN5uaClQtwtF93HsG2DfL9MavJ9Amnwzus7GkqeQ9lsVe
xcezY8o+IbUOsw/ENPnJCdtugS3Y4wEoVSC3krLruE1wqTlN4x6DyHwBbpRz5fdIL+pC9GD919QT
oK982Zl2PHUhThsLyxPLB0IK64rVX2GLocw8QE4KU484fvuavqxjJGu+/z3lvUkdy+7mO9lA4Fms
7BahZS5kgT2vM4rTyIgIVhrB+PJ8NOCI2PDMbiWcEcvQ2OTq9tUhHzTMKwHqa4PuoSWaK7ARKbsv
EM9E0N0e7K7cdxk5EmqfnXrFvflW4xK6DdenL/21uNBp7YACyPhNk4URU2AK8csgB4vq0MHibC9x
JrGT26Ssa4STD0KJx6ZKlvG8uycKdQ2+AxK/KTSsLa+hKT2HeIiHEVKBIYaZfoyrZCUh2KnsDBQP
1IsdF5n+Zb0znEW5kiY+pAcYhazH5XlBAJkEObG89cojKGvxfBTcDy0RDa/qspvuaVKl0Py/1Avr
sMnt5QKaacOIWjen01ID6RUX6ZvKcZAW0moAZzFvslBdZybVXbypfx9Eq2XgwpEC4voUIbQNrJFV
PyRoI3zpsC+aPwXRNuLTkp/RLy3JtOuNcUvy2+SqBBvSk+EftqCPrx+HiQgEIkTR242ztCI0JI03
cN3RTQ5G1QM9EYrS/pYnzeIG6OtvZk/s4M3MIBygyvH7MENuo8rovt75fk5T01H0I40VZjZe3/+t
ZagsFoZ5jgDWJ63ZtGnxcFKXjeFcLuQUtiPP0GqaKsu48iHXJncycJrR8m1hK4pP+L81/0gQBIfZ
FwoSm4rSrRVeH98RnC9S1yKxZZVMk4kPoFYXivsbfD1zQsxyZCnvdgirvM33gZuqMnnF3OjZnecl
M320EQ6m7fOFmkEpyrekvg8BDatjadmTRhlh2Ofjejwz7vwvHcAkZ9Wv+2JjjkvVd9Qj2KBvBa5f
S+ISMzcyF7El7U4CUEBUVx13diKi1EObBeZ89/cpunTcBtdhFEWHXgrsABMPM+jn2qBv2cb8S8+L
rfmfXKFGyfZfKfkQtje79WjhuvFksRYZFGr1BGvqJuayS0jHqQfe963CY1uDlxBtYyFxwLuNzcQQ
3A/kXWxl6M7XPNEaFxi5hjvvj7mWyGN+aIIKG+rdrg5BjlnrwzlPn7F2GMBtBvW8r1O2A6ghu0zP
sOpYlGSkEioejbYkNR/G2C8lF/+1g1hWwKjl//V1ikdKxliNayWy8qP8y9EsHCgXv7+QNjFUG3eJ
ruWSUKZiZZIdG9qQ2DzcTA84qD9nJc4SylM9u+fugx+d/bxUuESxstLMI0KIT/OW8Hwcabp6h+T/
vTg8N2A+X2w+ENdfApORl02qnCPFSBuwhPpMnjrVP9w+moiOBs0pI9dhVKsan5X9TmYiK2VNdbxk
M/vTWM7NC7agONqLsRMMuY3DDtTPOkdEHpXauX2HJ9cYSq2vHYKzJ7k8E7/TXySvVlB3H8XuE8Uz
U7pC+Do5Cyel9TDEjb3mdHQ3+Utl5alje3wfyS+K9mhjbvcWm+qWbvZO51TDRiFr2uvIcnrG3akP
a2v7+zTIMVtIsL1K935l3QHGpJsExUq6x7u3AlpBYy1jZABLc+QVEXYPcqmYDGdyZRZ+oZoFXGJo
RJabhaE5sFYuboGmWwPJnp0J1cPh+TkKpdJQSReG1ldFH4bwRJInkxDThn6z3WJzOI8fMur3aIoy
8VXJSDZZa48n2k36Mrb3HV3W8540fYj4AyFjM51mg7myd/wBqq24huNCgj5Y28tBcDf9leQruFzZ
1sXGJVBH/cIpDo5ZzUjQvSNnywl/OGt5XqbhWk2cNpuX8NkEhujU2Jlx+nHF4XqhmPf5sZX2Wny7
qWNJkCkaoQaepwinDP/bMKavK8NiKRVLV4HTkmpfk76YKblVRwQzrpYNEzQU4216UOs+Tl6gGtEC
BtZiMta13rveFNrEmchpnx6kW6kiD7wGVASbRVdkAs4szb8aaJwF+QJg/CYxeNYbX14guvKMaHzr
PpO4+UoALmdtW7/F7Ooop+GXP00v33HP6kY2K4tqvCO91VtJXXku9z1MCf5prqTxq6TyDPFzfIRa
t+Su2SrctttD04HjNUNpLp8A0R31gY6DV5lkSqcNlmDtI0u88wTF36cFdaCGrzlrEtzY6IfsMBdu
E+byCIEGB8WK2oRxL/BIksyQKgDA0+uk6S+1OHq7HuQHM/qoRspW7V1Ovw5OdOgGZqVcjmKy6wyI
EcT7nPrUth0OLqIRWk+m0AG1I9F2U8VOmx4EtChZZNDd5++qZcP/DUuXlVn9YZIX9GjMXtzL1CJu
gpm79wB9L9Ovz9sOd/U0AB+0KykgdrV9RGWxCRB4eAxfCmnexo10J0xJdeTdgUtgJpXXlkXQPRYw
x1Gscas1EktiGhVFZHLn7rZ4Wc/soQubXsHCflafMfiwqre7Di6fm2OKi5d3Ex1JIt/zaNTvqKY8
bMNArL+4+RLvVr/gKBkAuqruCnDEOjiPxXAUBsdaq6V0FSeILZpI9Zflb7XbdwPY82we+8mtbMiH
V3yFG+Lc0qm8RYBQT4RmRrKPvPMwqVU3SPl3nEQH05/aSPt4hEpBjCH7JWbbz//VbR9SLH9M2DXM
RIthubWzx1n6+uN4RCeUetB9lD9dmaoRhRAiqNBxOLiEEhNsO1yoXWqf0XNO1lSAIvfXVceR3VYV
cvnLE6fzJSnwH178kuR5wOsSrJUhPo77mv/fupIxBLafyeXHT6VciaLC1Pw3pd3SbsKU+La7XLJu
LlXdc4HSNTUgm8zqLmrew4d6DadpXcWaBX26U5pKJIkLBokow9YgjaUwJ/ulRvMntulZ1C2/vEMU
yLk5HOBSaoBJ44bamwXlWdEqOJf1g6Wu5gtL45g6HzDfONYV1rmtf170FNnEypE208sQjpQSkS/A
IxNLZ2jFlkcSp0CDGsIdmeJYoCGQs/rQC05vPK4BkyWZwGIE9J1++ap8vOUeUYHbHsPNpdcaIDoP
CaAbHTylgIqRRdoG8/xPmaj3KAiRWhv0ijoHKxU7rHuGW8s1OQB8DHShLKb4p0UDM7gohK2MMnOK
UO3b2fPWc/qsMiP3c48Jh2Z1ZX4PY8IsB4Yn3tgV6dszNAe3EvxlzCsXdFR2Cj7uZoEFwVJ2YbvP
0WWWlaAiw2iQrmgwlv3udOQlGgcQFwQi38F0kwH3CJ0p977ye5Z1UCBipCvRZYdg5e7qglD108Bf
KFI1FYk5gRX+bZH9xhp4zmxJRDBg6UwEwGjPyfZUI3mYUUdIRtwhRoZXgjjAvGVmILgAPznyTX18
WcQuVmv6byNatEiHZg3Pl2EZv8C0bKXZkxi8sBU0sC2txazx6C0F/VS7/FRtGLE+ugenxDb1Xsyp
0MlLjRjMKs3PZ0HxeGgyL3sxHiCx+QZz5hDN7K4+UmMaV70+vF/tey5eGN14Cia+DrrnQXe/iaJo
zefFWvT8lliDZwwkivkscmadlXbvxOBcCv82vOH7wYQyGKAmluI8hPSiRB1fn4GRFpMteCgTPhS9
qBVEmx9FD91BGiJRICAm/cZAZH9sjuoiWemniEjCGS+u4vQwdrP5Tc2NN4n4ah4WpUUEOKMxl638
ubtgFAdFpd8XIiLLU4viPaqBpKp86leEtwNnpfVlFVLE8KJlVMMLPWgJdfaCLlaxmspeE0KAI2sC
oiksbvRV/IzuUw3SK97P0JUz1fOW10YD8EL2Rb5vAq5JGZ/7BV2iL+Ntip/swRycGHXnvbK0d8aK
I5embSoRYMjZ587tHqn+zOwhEl9i4fEB9wM96vGfVncc5/pHXb4jz1w7CQMZQVb/1GCY8/RlcCW2
VbzG+XaWaBZexBgT9tNe/z9YvbJorNWSERnFp5aqFl4BLtkTAL9izOjCwZaew89J5npCTpNIz9DZ
Ru0a+1b++S1aiByzbpGA60keC/pBrRRI9jzkG08OpoO2eyeuL0zjHGuk4u5wfZC6becFdjrp0rOr
8jDOrkdXAVb6Qc7wmrNJeicsH04wvXmWR/Var+4dvsBClNJDdYKV6sORoXwUUfFLolWkxr73kSBc
qvlKYdFSpbOxFkRoMg4OmC3o6MK8JaG3dvShMb9cfRp7iHKnpEP33qXw9lDpvQJIK+gbacR+VkqK
/8gZ/Kn8UZzBtTvP07VCuuJDGqyX3emnPNEwn6wzkvqfRCg+PGS/tzAd7fg9YA+WMyMHRDfCNvB6
cl8A2RfPfHlz2fqD/eRZFOVSg7zs9ouV5HxY/uQ6029d48n/NnyFJznlKsrXxfNfR1A36JrVo4pE
pbmloXb6WVjcc4qXNRD5mEo+1rb0Zp03rYa8bporPPa3qrzf5rlonRJCpLSae/B8RSZJJ+HcTPhM
SXyy+ylxpXyDo0HlH5RGW2/0uKjG+KaKdAsQEn/ikIrJ6id3DB84KEwM5bbhkw25i0JKPeVSGVaq
m+4sLRM5S0jvj4VKr6pO0LrKQUwq5qak1UsvIukiqBYtlIy4WtWlyb7Sfq+UG6TyoHgE5WId9Rpy
pxAX38TiaYXgNJ4EOGfeG+jVf7MFmj2IdKRIxwssOvNFeJTuILdeYGs/Ge1BOdywgv5rdmTGsGm/
lGR5dYuyiEUq7MuEnHICjek5R5XLiF8yyCVXaR+J3UjGqGz7F6A+k1A8/Y7RBFKwgfg1FczM14M5
S1sQD4sSFWbkm186vzMEyMctbifbSnEXB/bjwkG8PHSXV/FvtfAIgABbRLUq13JsYM+w2+0HPua6
Pbo3rw5X2hGnkIkP5ymGx8ELV2MOQ5bEfimoGdqO0kn/UL6XXTPGaGWhPDiebm1toVvunCYPmfSe
mzCrZOkX1mjs+Oaq1/Iikvhz3RlXIRc8/mEIvoA0mKzRUM9mdqiLbVn9YbARs/OE/BbzvntuQozW
sJIGaL2gFAfvrAMxdQjA5JjctJ4u6eCJid08YColIzZ9h2SapjC7LEHMZjGTgmQBYDhzUJXKcIxJ
DtN+3JecR/QT79ysb77bzW0ar3cg2X1fwGGeKCJkCBoDIgA3S1e6cvc2VS+h7zoXRfGQWNfc2PyQ
KskWtfa7sLuKBCsA+eC1aSOd8lP20JgwPLSah9AERixLW99HepmTOPpjoNeM4fXXqz4uriwPu037
RFyAqEKXiDWUtHjXNmKnuJvf+tYM5upVe0qPIOpwB/fhbZ87rXHDeixbzshd56FBHGJb3AT8kV34
CAtxSteSJAvVlU3hGSHS0H0WT/TC4wyxh+HWiO2WuaXOIfywcSO4XNEjzRE+ThlT2pYYsiAodFt5
X9WKUTrg/NHy0pbcd4hsu+pN3xvpJVy131GqyBkbX/qtWywGg6RTKNlxrVbMQElRftcnzsOCSf7m
zYllt7sDR4xVQSHtjDVj9+OMd2rQjFZ/6JQ6cdJWXbJt2snCjSkzymbm9hc6XIoPA/y8VhFSvfqS
G08qbRBkq/onspkAaGONfRtfbCBWloEur5C09A+MUa2QQFnS7zsWdf7ZUzBISHjWoPZpO8jB8Jiu
6KwCQiZ3t+iHoiLccVoGFYvn1J/vIkQDRZjLLycHRcSQuFgoa3nVMAnHEH5x/TQthfc0Y3TC0OKi
BlgV0EFZ+HGreZ90OVDPVwN4D2RUGhZaqvw0LSKOGy5lC3TraGz8xpNvatTV4VVfJDn/ahQDfdTK
5HtcJeaANhHnU8D46BgWu1P45fPBKZHHODzC4qtk1qbEbK4o556Tz80GZ4/KPhbL7RJewTLUl4dI
GZrBAQyOMUHAfLqdusSIY4JM5h6bKATtk+AGw1ZR9cKxEN0YrTIO2wgNEMhJ9xWSI4HWYuRI7znB
3U0VrOeke71I9id8iojagmWOeKckzCncyM5sz2mhD+o1eF2dBJJDY0NKJBCkHkbbuXXQndkngt/k
TSJQo8/jMQHnf0PR1sIhOmqwPubbTD2POYWD892wnqEXMtRqay9o4RwIFK3Ho7bM5a2AY+tlJOlS
sL8z+ChNzq1alRN7SMVnpBm+92QNPeZfjE0B7s6a5D5LIIXMhIi12byoqVANxHEp62vLLk6cZaU/
SMPkJojIH4yVt9HgqLxpGTZaSVAYWx13rcZicb6fxn/2lQpJb6DnRROPHgw3BkNHHjeasCrOVvtT
ZI3H7ne012C8Id7wzADNwpi2BrGEyOGlvSDbdurHNOXwP5Uz5cb9YI0oIGzOUjv8KLDJKpHgxtna
hsuXBXCKFvpmwOhFwT7Uvb9kaZXYhbPPBj2lKr6fJGsO4o5HcdyLG2Be3saTJdR0+kGqFrWZbnPw
apVeYUqASU/L0X/pz3KgZ/y1t5uR/oe1XpFzv1J4SBSquZIV7vU5OnKLJyHxpleit++S9JhIXC9a
87l2AtJbcRM51L0BytsdhkNuEg+DW6YX2/Y2ELH/Apu6hA6fLSzyusr2COtnRxDzMBIWY+XN7/kI
c70MqyRLsqIIOwmllxHC5NukpNYOO7eKNkisD9oAbmvITBDgPhmwBKYxwk4QjGRmicxakXfC8qSz
xfpE0ynEgnZ/b5SBud9D2r6PQUs3YPSm0lm5xlTRCio1kDl22On1HrefOnWeeqlhTyVdfyJENoNd
8APQZ1gnQFJDoD3VqHt0pSkUhoTz6v8nuMJ3CWDfuG4+5kOmnmxuVCfc4eVnnmgBSmhfPKLrVYN8
622e3WZblMyPQngHSF5EpSrMtbKFg0ePfU7qhT2VmcVAUVbt/QjHmDR/XoBMS3s/xF6K0CEPKOih
HZUcHwsU2d1yQvlXd5RmCE+LRUK5hjR4Hr6x1EHv/0JSILh5+DO+XMzpCCNWEz9w/V42lTD7o8XX
h7pgmkXW3wN8JbNrQXQZk5yqSrG7S04K4EH50407jR3xjDYgI6dmY1KsLu0Ahb0BfQmVB8NgM4oJ
d/KN+/QY9cIYvMUPvetdLgWj8v/+3riWfrSN7aEz9s9JG55/l73yy+7aj0DNRtqVwlAt+4On30jo
0vawiy7otCf/AssVLiQ6IG3DlQwBgx5WbBonikuWIyZdGwl7fGL/bTmMCqUw4GkRhXFfSBfraUSm
bmz9G4sNk5JpcI7lTVdWvs2SkEQOZcU1HVTJnhPHXZGzSvHt1wGPkCfqJ3zt5FHVkD93jAESa3YQ
if0m0emGL6P9KtSw2D4hd2pM+DboWbhFPqO4fZpCanR8JkTkuzswXZweCI5Deb+30tTEoYoG26f0
J1aZwZ5YTTOtnIa5jfC5zoj+U/BnUY7VDr9r9kRf6Nj9tdC8LVv4hyMyvvYpn63vDL1kKYzPzNPw
BFSNslHtO+ZY0UO+onAamZwdb0VUXAdJHNYjOwxG5wpy7Jm0s6dV+RT6JTJn5Kk2xmHXBbi9MbZA
GpE4kFcaiS5Npi2galhw4urR6/rUT9tk7lOzfGxP82LCJ1SAzc37bgtaqgiKTxxJ+75rpGUALeva
+TS8iGeVHForMrhknxl4dndhkDhoOQSStzeIQSK9XtMiQ6HD1wUWZ2t3wgEgk2CaW9m2eXhqv5Em
oCWsEDvW2aFO9fHhIP81hXpzlgE1VE/cX2jRe+a4rQHsFUH1JK3i0lVxVBZrVyGBLe0AZQqn1GXq
ATnzaLM0C8JEQK+Ld6/YD0YsB5DeNKmi2ivgJZagZ90SPm1/2GGweaNiPQ/Yjvr+yF/SQEeCV6Ko
poNY0dXr/GMykFjlwTwUOzb2dOD1/jA41JK9svgRJXUCyLBKljXupERIS67oHGTr5xrGvsAwv1eN
67SYL6LrtS1fe8vNu9wcv2kfJ4q1kFkwClCelBLx/2B5x33BDJ7WDspBD/FGnNs4FSRAOrfm7wQY
NEOnzVIb1mXB3vv5rzV8TKkZL8leJStHKZrHt89qv+9/K/R3Ax9XTFLW5P7mCLBWd3eVC18wYbs4
roTyag6JTM9ebhNgRC8r+TLrx+IyXk7DmPM/ZPngPiWrVMQJKg/URH6HV/qrcYJOTmVGD+D4f+S1
jFCmNCzaAaCzXOYHhuHLt+FEG+sZkWs3ZCzMAmI8HRv3PCcByhXWx3C6088mdSOPUwB+xm4JWFX4
/0+kM1alhiThxTC9r/y5ed8tjeqLQzAa9npfsAvbfDWo9O1rA74/AXpBnF07pW2XrvOAm8NMS7vh
QpDsGvvMSdJUov46RrwO3JEB1JV24XSDobR57xI25HtUGewxxZT/LsbK19WHEg7Klon2DoeEbvDh
ysAorBolg655MOMoRwmV5iJG6zc/Z6FTg+6S3U0266GuEsqtl/5QU8eMcIsCyVAKjlHTrYSv3Qsm
Wh9bgcQOqjBsVlzKpasB3ihcrTt4FhJqCF32J1+8/xVNUHAtHpCHd7OWO/bPT6vzeH11DqUj+FdL
urLBedCoDB2PBsKDHk1H+hGmzXVWjrW6p7ht+lDLOb7b0ZYMmOnKnAS6ASJS6JFsIr8L1/stXbfJ
nIcEP6FCWhl52VIIbjBu/7s9vuZgMmRZzPWlOS0CEx099V1RPH8iqByRPk+JVl2BOZ2EBv/jLgVJ
H3D6vJHGQ70ZEidNrjOM83mt6RQP/W741Zd+JbK73mLz/Sc+a/kKsNi1Dsi0NVlOxlTz3dMywW6j
S4KpvDGIyrnXOrL5aUkcveVnDeDDVIJYRtQ5CYlPdHwENvMInF7Qy4+6bztpTgggfu7b7Cwz3jwv
pOp4MfS/ktIdiKnVsK/Gv5mIk5iOQrFYm7cXE8wzPKVUttMkQKMs+ZghMBoi3FNzZ+d7ck6RmpRK
m52fWHiZKbR8+7xrsFW1R/INiFR9h7Lg47DDU1B0tW6qryzRwrtnvw3axgVGyQEwUTcquQkRVj8y
uuh/R03AjDyUNBEqLx6EAYi91veTPHWdJk7lQw5cLDt8lrng2WlyGJr1ThkFbNkADGNa9EcHP6wm
BA3rdhJgef2kiHcFt0YjBt58K8UOijo8B3MWLebGoTYmjAyoxQfEQSCMyNtenwbCSSohWMa3s1Cw
DtlLQsGpyJzGCwuvJdyTtl0Jz0TFeFBEOM2P8s+EMCO7GOSudizuqWlizXrU8XAQEVmr1L0i9aMe
ArVKVpvTgGXgcfZZIHiS9TCGdS/H4VJ2G5iGEM5mn7Osg2neo2nlV3jWH8qvSaiQjwzccv5d0s/h
MKZEgtZHMZCYrCw+vetyqJ9qQytRi6WIs/Za+MpbllgVviOFTARZ3ycgGfeMkl67rXY8zoQX3+6D
tplKE2LvuGIH82mL1oqH6Ix8S778oUuCxuci5KQQ/jdzgOZxC4VX9AudgD62a08q1Aois4kfuUDr
LBp3vWyKvDtQWjHAolF+yNwqVWCR/VEBQI7/DB97zIcgXgeCS8+O6ZdG0ADneo3Id+V50nu9p0Ne
F3bOBQ4yvmrXxGI66KuKaITHsba54/dJ6OoFVxo=
`protect end_protected

