

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PpoeUczC12+YQ6zcBW/hk7KVg+x7UTioMUTG7QSkaE8DKLm5OzMFnRnSP2RdM8C+WL55mLvLDYfA
5lOC4Ruqpw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K3yZ7/h8XZC4VnxKqSX+X1dWQEKELq4EziAIjvSKKzex+MM5ch0NyAGabLWybM0VZcnyA2IuBQRw
LXtEZmU52Vw900CqGAC8j1ob1JJokunlfDgROKOp9VekmhrNu0zlywHl+eh6CQ/t5W76EWfCnLXS
TKcvUxKzMPqBkiVg3Y8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NSAGB2MTAPfuv2AfQtQrWIP89UNTneL4Bk6/B2TdOO+6mmG5j3iveazvIvg7qIHwAqHfCGACbbAp
fGS79Be+x6ilLMPgwgbPlwYl5oARsjb29GILZJJbq65kaBdWWJCFrRmIDIFHXq65c5qChGV/7EF5
BRY2p2sjUe67cd7MFOLVO0mKHurU5wiieT+wdpbGs9uEgt/pGFeQKlj4ch2XzN03R8Lg3KmqOC6w
j6pa6lYe8j+sQMdh+WMN3EmYurAN2aA01NOtdnD7EoaLrP3ByXrwCKFB06hQfAMKudCun+42nXbW
17uiY727vjm9PIB2xOmQazUdPEZbwz2Eeua7KQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NPiHNhu2YI6wz7attBCDx15tEqFL81ie9/7cRUJzlr+aO842fU7+GGF/JOlqWsuQg2RB92onmIR9
gKmj6xIVPN77wRnezyej9aQsYy3bBfOSvbf7a7d2lZQT1pTZcYMfp3xveVQ5gTGk/1BN6rnnT8J4
QRALHC2oqPHhQZ427wg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aHttOHUQP+m+tZmSEhqIMk3Jbc86fWQ1/2LKPbbHBoOHb+XyETCjDqnDo9IWfpo+m+LC80obW4Zd
cXgM5NoQ9F1AYdG2ggcdGNXeaparpheOz+XWEe8nirOAN+Ks5VYo+yRWYwO3R0Y+0V6Yw8r7cd48
CXttfKVhu2QOlKTiKegYDKMRGhVyrdNkx/KDldRFk70rkBceBbiSjdBniOrozyhG2imBoMkKkCmI
8TwlLhPf5Ra+r8wceN6j4BjOnyQ3EtzJgw91ujnHo20MZFiaPiqLQIavDgBT1y7leXT7TIK9Z2uu
L3Oj5XHzPc1v3FMsMkjnu8xWqC9pP05Ha8xR1w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26736)
`protect data_block
mLZb2L+0wnXsQLsTjelIVlofuBcKO8VUU4T4kw54CDvDDha4u0ly3VGji8bLvoSqHdVsD9cQZuzt
WnEhYb2GXrJdRlugGqrBkHK53j1zsBhFGS+8cI/E8fNiXXoIUjMwoK5WwZMomTu4a9fqN1AnW/6r
iquRDa8jhtQNakmktpTKEU5aY4i4MInkVaHuG9Nfrg+dwRaiPazynTknU3NRJoTCqZ/yK43UfrQP
bV5Y5wYcx63FrWN7iWwmGsni3GvpJBvN3y8qtDcoWG01Cj0oxHbidRO8anBC0il/olEliZd/ePwD
zw7MyKB2eaG30iUZyi0OjpTzi1XZCb+4ja7kV6fA/RMyHt7QRVbX9EOWb33WC6zclMOdkQgdnvX0
Pjd/Qa4kid05qe06EqiT9Z6SX2c5pAtAVRpD+CfGkx7hf0z3FrB5drLZr1MfH0HaGqLjvJnQq3EL
m9VuP81c+igWcvsao+DUSKGV69evBeYoSJlQjVolt7gqjkCxS+4jAAyVButfUcES87fBJsuQqfwj
8EcjGlctWjS6QilU4w+skwcFMFU4SHwSXE2x5iOY2rPCP3tJbBI+Nouku0GoG8TdWRAoisJfHRwr
ifV49nFtmLhwre6x+X4ghibwyPSB/dvfCxcL/CsKqJECtxWhEKgAzsFa2EyhyRgLu4v5xTsuGkYs
ytPHO9DvZe2uxdSGSNGkU1vljAuZQgcoywFZz3EY//t5tYiHEhiykVNFV6mKABMbLhEzeI+NW797
QHq88iseY2vuwHTUy4VPuRO/5a3Pxzf1fKNAL27T1k4Uw5xcZ2+lmLC5H3heW4rSgK2Eid+0Or5l
z0zERD8hyicfUSFecG6CWcz/U8Xsu550wmkOE0/Y1F9rR90Yx9Xopg724FTuFvBmVn1ptw2hUil8
rWXUuNrP5pFfiSPu2NPYzsubbaCnmR+xw471FmRDvH8lgES9MGp9Bv/5BCmof2GPAAwg3cH+rWkN
gv9+bL9xQ5UQwsQNt5gIbBY4rvrE1TebxO6CUuYMG0PEmQtO2Bd+i5grkX7zjEiqHenluGVC74d/
sNSoaOwkTOVQckrfx4dmVNzaTp96TylQosFbtiKtExCemUyj20fc1mI3dPT45gW/AhcBcakTwkrr
QQhGZdv6fjDIP1dMdlFRgTc7RWC55WXlIvFvnlwbgQpnnZiqCgtC5sjqvEGTErRMXzYose7Ocqem
kqhW3akyvTcuoLOJKkjzUtA4DMAwXNDIqzn20obTrR6/JlUWCucMIoSCVg+VsSsBYCF3+PyWxkRP
Nm9QwfNgPwb2pS1ScIKSeUd4eBSH7gaP/fGvyKLHMPGPaQjDBNdhYeAyFqDMXdcfPvja1iC0l0/A
1ZOMwPQsER3nwrzdguLcOsRjnpe+rFfwqda9AhHrayXdEFMQfa4EvNI0scCXwlvkEBqob44PuG+c
3VGEBIUAS8y9kmHSoakiwbzvM5NAAdITtensZAC+5k2qv4+jyO4spJDtPtd+C/LL5X288Z9lD211
lHhHPafDewz1Mn9J0JYKjUqwaqyDnmI7bbeX4bKxwDzL398FAEtoW7qDf36uW2TCNseu5E5sCLSx
6Tskjtk8+yn/fUa2m/eWL2aKTeHkb75Y4bzCpz+eIGMsF34CCEnBDLtvC9g0kDuGo9qyNMywP/eN
lvn86TQ5hTxj30C3mkP1bBkAHnRgAiMdvAqsbhnLsi6vyc9t8rKAeF7mMtVoaDV9L2IFFem+YFOH
rJXEkCAg8kDaR5BJEKtu8C3l/VccvVbbabvN/nxWuZWnARFTW2xved195yc0K4FpBQNWxSkcxEWH
bK8uCc3Fb8Xei6Jwl7NWB5McW/NG7gF/or7y4t2yJuTaBPsPPdmR/munAMpBbe4/e8GkyF2003gR
0Gdc+ls7INx/nOclXB5zYEec7PLrUKV9xSqPGNwD4lMYlK0rvhD75OBOzz4WnjJ9aoDaIYeaRBaZ
gaOOhKxNFuaVHHoJQDQ+eoGGf/eVUclOgjzS7cQdHE7Eq/yhDjz8AcWvhCwy7BvkUvHEVNGR+0Hb
Wg2aYNzPgpY91upTyc9WJjI4VFzgKdbfeqM2vVhHNIDkjKm8NlYlwQhcex/4hdtg0qxRYbdJuv3N
Gt2uP3KRdjzw2z2+fW1oyQefetDBkMMlbve2U+o1bh0A9DVRkMMFcotZG9eiMOG0NwNcSvMQ+oB7
odJbGpN3vJ+F1U9Z5kLF1iFBJMj2L2LMfI0qVnHGh1WWUflqZIw9tPfjQnjDer+zfWz+oxYSfKZa
Cx5i6gOpqmvEFWb59VPDVDJkcDBXCIDCBqNj6W2ec/ururyn+JgpGMdwhNycs8ey1vbzykVbCLNa
Hb1Q1ZpL4WnX2YAIxzDye/ZcM2FEs2L1LT75zoqUI6ipzz8I4L7rN5k4aDHo5o1/cKuXmN79EJI5
RG9f9gIxIrRZTRurGR5/ptq8DKTZV8PXst7J5aRkzBM2HMHpS4DjF7UjaGpUAkVtB1OStUrBho8d
Aemv+JEdQPpiVUjxZBbZiKKH5O6uT8XYSq7N8Y/GKt6lHLS10XZ9E9jqGhVsYRzvYDMRoPWtaOGp
jXkL93bUpk26818eSRguXXDXAHpfQ8t7euwuyBPNPGbalF6u1AjRF8RtiUn+k/2qBxqdsFwrPCxp
jtkmY9veeZUXG/oJ4qMBzDdk0ll5g7Gx0iRDGNvPFlhCu4l6f7Ez5pdOLnFKR+xsIvMQtbSfHVHN
aajYfgIG0Ez5lnnAc4sTWlfuMe4p7h2jOJL3QI6L2WawNc0uIm2p+qsCetakmRGzOg123PGM04SV
kauHTD7HgHxOghxhLWEIyHYYILRbG2m3Os1pmRTqcAbOWmjATHpzbcum7oNCj6slJtBAFcaHFQ9N
emTmCe0BZ1FJrlyIgAkyGJzdK+p9unilG+Bey9rweAX/pTLQXhEwfUIbUiP2oMJoWBmj66rUO2uR
ahJ8C4STpCMRCXgD6uS1Wzh8XJbD+irRqVrgRotcS0IrP1DZ6O0Pu6IuMG4QPF1drGPz/oPY/uex
LCKe74nnYndc2bppvzJOwpyFmnP3C8RdI02ePuovCCEFEgXO4LdjkRPPi0lzCgrULen8V03iVzoZ
X4rBXvPfdcRdhWtKWlm5gIFWn8FV4YHQadLCvQkmtu67y7uMKTM/6OUbgqULpq+98iDXujvxvNj9
EQ27m+QNwtBMSOC3HLWf7J+/7AFlNGdaTn3vT05eSlKFURNoYIdfr3RbzAF9kFdhtRwTvnjoswbZ
ws1RUrWrRpcuDIIZIJTkOxbyhR6y5UZOOmjI1Qc03HREnPrz8MPELSJ2Hb+ioGUM6RJdfZlJpVSI
2ThRSirFAxuq2RdSVhpQxf/WyduhkwW7Wbx6m3bM7rJRFGHTZaOUX0EtfEzvaYvAAmtDhe5Bf6e4
7lNGhHpMkLQ6E5aWCqtYQFZH2zjAxB7X+E0SJ6RkyohllVmRyecy4CT2X+pphBPJklypGOnWhmzz
5RpyGdyr/BEHpOBjNaCmnMm2O8zQ+1DIFzNaggAypG6ftpFV6qhdiEg2epIjTQxGIwXN1l3GfZPX
dJ/HpB2jBE/BCkgQ+kt1spSkSWPC7IY0rxSE38qlsqYEVHQZss0yzK03rLLm8G1jMMdhHLBWnHkK
aaDI9CULOtuswmUvVyCmzHLPTkSMHFcxP+MznSdj/pr+QsHZz4jxalNU94Fn5w7gkx3vlPuHG9Xb
fxSNDGsFKgf5SlMtMn2YkqITNgtBqlxFYP3/gw+o7e9iEthLHeVuN6tSdn1uIVBYoaxkwmbSWLfQ
xwVi05aMidBBv0+Gj4Od+CZUqImsTDimKf9ypYaQNeOuJ6T21ThTCtRVFxJlg6ZQNqIwxCISQdlQ
gzqENJerlY+jX3X6vZAfVL28Ra5f4qq1VkPtTFbWw/W4Rfqof1oQhmqg+hzUImJA7+aBGcnQmwNn
ggJhvJ4zgyR6ayCA+mFnnb4+5ktZy/1M2jA0jcGkbmYjT2Xt/TxLtFyZa71Sj5tYPetmhUcT4osZ
PY9+t7iN/2xfmwruSfe80oucV0PNqf/JZ6+3cLOg9TRs8R/sDsiFwKmquFfHO44gX8Qe1z+4Xcnz
Ne4YAwbD0Uzj++kyGXaO95dpZdY4UO0oduIvmxcwNRLIfaCAOWrrG+6flwyst1+THJza1I9zUuP8
zbCjG9UFnrowSJs4khXWR+72Clx3R+9nUAReiMGqtbAadOmcu1OUiB7fYZQO8bneIwAC2U5dSQU8
1Uy/XKR0JOdwASFpzGqBK0YI6Rkrig+W6qmfH/SNzpkNa1Wi9B7Vcven/9FqOws3WC7njoiuqPBJ
V01oht6PmlEK52AXa+4AXIvVYsJBjVcFJG3WOkJWrB6KReLmdKNWBhLUgTY/5bbdRsAbEpuqT1y7
iLMPXUoBj6vREDG8Y/f6Ej26rCM/oFsT0SZ3Lu4h/wYv523ybvA5vGj8VuodzKmb8Dq5/vRER8Sn
gaVsBoVrvmfl5ZYAV5/fkJDSK56Dcoo/oIolI/JKtPFPaH37Ow5DPn+AekJUL7OZR6U5r56msVxp
P5R4vlWdcEd7e6KK+mVHOZxDeKtY+AQCQZ2MCqvvR42RiY4XD1SoUv6C/A9KcKFIaKcgIY7Ds6W8
Ej2VKawheOqs/xHixi7/eE0vzFhrSQ/o1HRqk+4bxXDBq33wjsgi7flQUiUuxRFVkRHdyzHYFQ9/
U6+Pe+8310pZQbPcABPHpoeJ/3TON3sfgSvXGhIY/hKqKOzLkiIrwuD//L7HEiy9vYG+I46zLkE/
d00UNAtUd8MVH5cjqwOY1rumKS7A0ki31UxUVCzdOJrnJbK98D7U+j6duYD9ySjUDmWah/3gGn/O
vG28ejoPDsD3A01OQGfaRIKAkIA2XldHzBlSJ6qPlV7vZRTUDl9cA402FGhE/TR7umtpvWdTJzrH
MdZFD+tXPdaGWbyYXAuI+NtNcuwkwmzJzLVX+5Es4YE/Mt4y6uQHDihfSM+jGPE320Hz9Nus6kMr
3ByQeHEr10xmRZnBUBBml0ZOjnfWMEySY/ZCI9r2yj0i4pFfvL6b3tHLlMUzrMUVeOgkcQrpiOuk
nzCIZ+DCVHhGgOdC6wj8zXy6DR39h3r5gCsiqfN2SeWjqKmHMJpD+rv7o0fWCmvA0Jkv2Uwpefmh
Yrz5F+QBciU4BG0xvE6l9OIg1MwfoDqLCLZ/Oos0NV653uQ/rA1ITTPrcIjFYMZR4iQ8601Pol/z
4raQFJLe8oQo45uHRPUCrlncQBwpsgXYJ7yc5+s3taLWbsi6L1wyRcnIuSzi6KrC19FraoCMStJn
3fR2bUR56Gn4dfanZrVipWpCafrJzNyRDyYctYgy54+Z4FWf3dlwZxpuTU68mFASk2SmpqaWvm91
RU0lC+V3x86m0WhbXHQBwep60bb/slUlN9GDuf1tKxBHg9EOTwXmuNEXBMc9zML06CxCAxF5AFO+
uLNEQr1kDtsEJuPAnUW7ZKI5dSfAueXcLfzTKcGOdqkBgc4yW/WlGrwHEEbiNDXgIzMeujGJpxDR
wtRXQRdLd2VzfOhHGGMRbtXtl+c6F3mkhwtEkrascr3mQUB6qWu7r0in0mr+RAknhEuPWPtB2drg
JIlMGSsdTn+1Z3A2guN2/ldoRYz69CQMOXyeZYTadowK9RkYEYN3HHLf0wolhFBkQVBfbBfuDimu
h/hetqQywRccT0BQPEppaF3KiwYIMw/F0U7fWzfGNE/rYH2wW1v1qUBYkUOsqQeW8hLJovnOgku7
1cA8tXVQV/JBRqPaXU9ZNOlQL+1gsj50WGcxcA90PFm+s9bIO1M4pRlEVeH4ER5MoH++6PG1iyEi
YRrCN+UYLfhBT4QH7u6Rkt/bTUpfSxONkDzLUiVhlgOoA+D1IEW5p9b9mYxYPFsEuhbPMaidBQgH
v1froaCxjqoF3K2X4MtRbC2xv8vLSQWD4Y8XGMKC/N2BTgBJvMRAvoC4YUpJomZpF0WcJanjVbiU
bMY4Tn84XNlpXBHY7zeCiBYh7as8YiOLWjBJqc7f/sY9aBCzUoEBuEZxWxJPrgRU7OsNFVwG0Ch9
pES4Ehfy+IBX4nvC1cWuvJedVzIkxiGpP8z9RJMaux+Y9ro8GIv2eB7E9MCD1RO7W5GsouuaqHYQ
GuUMPm4Lw5YqMx9kC3YlixN6Jzah91emsHsojTIVbqDcXv+SwHJy2EfX09BswcPAkeONwHUqT09W
1qeyjCUnCmK+n7CdsTSJFudFgGH3jcOmLx6c67QQu5Aowts6xCVB1xPKCRmzXlA7eh1L3ykVZNBA
QZNTmksE5PfiwJ/huYKuxrj3edUgS7ZVvKSRWe50oV+lpoKxbcpBuf1QvFIfPfspu8QoBLX6162W
d+z2z4fFwVwXvIqh6YSx3xvy4FE74rTzn91Om6nAVv5IyDwPuGk2QrLrVAyxp01cJVP3IbvqOXzd
76ZSvmizNxIU+hAS5ACM8JZtvl+XJmdoD+wSgxGR4qAHjQwyZFaBG+L0dMhvjtjjbm5dxdYmFSbi
0u8d/NxsrRTfrkUM6bscwtBnsTGGYvuDVjFCbcINg/KHeCaZkqlCedxWoBt9lV3TFXNhpstZbDoW
jmxnFOeEsYj0xeLosuN7wkhOMg4hT7sPHjd0jJmn2HAJ45Iwg97GDZCw6OuGOl0p6j15vc0sr/+Z
ZcrCiiRtuvsF2GX0YneWmb02AjWkL/jIx95kQK9ySus8jN3V1obu9umef2GCcjVL2nRwNkPvaDoD
xQqbys6f2GNT7zzszQXHnq8BMcMQxM/o0T2kZhE0LUSnkgpCEXgxLHSiZuQYQtv4/X79STP3rfeV
GacvMkpI93Mq310jiEzUPomBQNdr9fpqi3Hf8LSYin/Unj4ZPu4Z0rHsA2P/mXvnXpTccdXmK0aY
tmE61jprFynTeozn+g9oiI+NK4r+TYPObaIBdTmRT7QqYAD3num/8A2Pj01//GX9MS3Qg0QsPLDW
LhiwOScjzWdl14WgK/iDxL0K7GFVm0QBsCzpr4ookBUQx1Wpam4VgLJ685MbQwGjs1xzN0nbvD66
+v1scr8i3Xw85AYywp5hkQaX7j6fC7VfiVBLbvZ4gzh+Zg1+jnUIzOtE7huF5obts1dRGCPydnue
Pvg0nK+cDwEboRW2A9s76JM7PloNp7VPjZNJY96Ps0HT7btKmqZUwZN7no/watD9uI9b6q9NmN1h
8ycc61PV/4jX2wphRD9OvcACB2ZyNtiEA9IRPZMXQu34mzig1tVw4oNl+d2rMinOpChGjTkKN4Bs
vr4tiSFYXSMjSxZVWg8Z5TGdD9rKLMA9YBdQmzLBFWu3n8MgK+iIqVdQiq7cRd/dAE3t+H1Mvbiy
W0CKx1avrLw3NovdtSoqtigwCOZIgRgGheJbc7U3O+hldI26SEtsoRPsxy3rqwk7FMPpOwRd+ejt
x6b/axXKUuNAbX2L+pLuCyCVlSnMSL47+pQJs+GabxV20MWAHdY1wWfBEt32Ax33IPTA1jpZv2IS
Vcaz/CtyYdxeMMhjwV2uyOBkezjghp6Ek/0MpPBG/R29gGjwXdrZ7mm7xvbXy5SCE1F/E0dnLY0P
YIjDaLJnztg/PiuMp9WJuv0CAzUwbjcF9F08O9lMsnQ7asFSUQqU94GtgCBAV6LTy1klnFAAy6Eo
+c14BODi4RUdaKniVQluv8A+Lzs6Yxy590XfoUG1EVHV3coV//4WwzXjUIePc0YIc3BIEXyJ4aeA
rt47KpF4joyFBgvlnt4A3Zobv3vBzfTDdMNOZlXT/0EXHJBTZnOawlxA1kgb3S9rJEpTV5Ss3rTK
FYAlNfEjl+BGXoq7eNjQvpnoH4Vxqqpl6jOYWVAr9PagGkUmOOGTJSahX7PeuwrKMYVkuUV8rIjf
nnnsakdT1MBv/0+SXHUBaDQAw59hxLtL28OEjmUbbePvHTFV5PYcOWPZkce5TEbWGeCn9w30iyUl
oI4ztKpTA30BQ/dC9v75AtNdcE/RNlCUv1C6olr/lJQQHOpD64ZzLRvtQmmqHub0YKlP/Cg3VRgR
MQHLszfRtu43b+nuRx8T1Wppyji7MxpWLCU4un958SQt24l7y382f+QHOjmRbjHrtxpbnLhOjXVV
yhgsMJ4u3e+78/fQEEiKEEinnlU4bv6OfrxdSKSOH0WJS3ilFNikBiy4AIiWprmKiRcU0kS3EGU/
nAdaoO428//xgLZ+GR3FQXLDKNXPaAm0mRPsFGFumKk0a5EybAv8rdQ/ZHFOXCfWtHyUsJuHHpQS
Bq42MBJWsI9xr26nWWLcFyZZH78rqZ0jP6eSo7bz3llAoWQSm3idSmeT9C7oVvcGYa+H8PKfa5qb
y2ie+NWg40LK9XVqoFhGA1gTxH22P+5ZbDSakf9Awk83RlpuwJhxeuZdNL+WVTdTnoVGH1sK8Hft
o8qwe2XyB5RLEZkxE+blaW58aH5MtpoonYtTj1Itz6hZu9SHS1ptGunisFNgEsACVKxoSwPCQVPZ
cX47DZPhpuuBNgHoKf9m5aJ0ilskx9vbZPyS0e8EFl3ZITxrNQZE2Sxx6sGCPoLYb/ovFfzBUP/m
VbUTsxLcjrnKpxAoJNWF2yBSyuVPqsZh5bSZx78ET0sGn4ADw1kK8si2VGdFJjzKGz377P3jn2t7
JgAmm87kO9cCFJUSQ8lMer30X5GhmEoU+Bbcx9xU6v5zST5qvGEC3ilJDuO/HJ9U9PDj4VSJRZmn
1XCR8nUdr//khSVhEsLp50wmmbaWUigcAmFYEbhGTR4c6o+wdmVaGHyFO+Et12U1hEcV5GZC19Cb
RgiCzBs8GEXXQD2qZEus7ESWcuwDjAH4eis1CWpDvv26kePw4jTCjuXfhRBMNvmK5NnyI0hD4TRt
t9ZDAB0N1DnYlCt7uJ1pDoHTDtb8MN4A1wlIw+Zv8V1XT/VpuX/AxUb8tDzPAMU+KngkG37B5oNT
UTeWSY/VOt2gMcwoSbPTlSfA8nX9J/L4qxS81AfA0DPcahhlSjdst03exeu9Jo+NJWmUTC/K2+6e
RZcMNWz9cQ0lLy6BYSsy6w8FmA44Ucm6nUOMqCibXc/zf/c0bA8lFsjDeELZbrblH2DAx03M8J9t
wi4MUzI9mNz2st/HBf3sLm4ZWOZLMtrtEhMEctckMqOz6vVTRha3vpJWO6WbwsyLX0eAkZ28TyBD
vU72Etfj9UL3Ne5mfRPWH4gPvZCfDO6myHuMbMeKjFP0zK6y73oDm+oKvx63NZ48CgUq3004tsI6
QnB5CnaBYS2fY4XudSZ4VtNOdTZdLcrRYxgfpoGanKxk9B+cNa+6yiRgvrM7ipVeSb6Zf7GSqbjM
R2wtI9U9e4DQkx+kULoBE01Kt2/FkgbCxox4OWrKpka4rNcmeMVW+owU36KJuGCH5RkA+9C6ax2d
ZSn2OKFhd9BwmgxNl5E3ruaI2hTsBy0i8pSHwhR4qp25FeEB4AIg45Cdf8HL/H5vUfcQcVXII5ci
w1KzzhKYIJiNhJaZ733K6/FmW+ADz9d8c0n8NuhN/xrTgdBgnlh6NPpsxq0S7eONPv/Uc1cvetr6
Nb3N6X8Qypta52Rg1DbKcebRv8d42SbeZoedaxKHtafa7clDD9L24lRpdtxhbSKcLiO+fA+eEtaI
Bwc6y+ee03tPa7kGAXhnDSrZWyyWKwUSOGDYH0G0K8c0p29zH+oHJ/jTgSa4Cm47O9AjZyOSkbWk
YStwSM5/ywzglFatD8HRVw31PEIkHkq5C+LroPWyj5hco1/6cpcK7Qz4hqvMlAQIVVgj+lEbG3Uq
v0QbSwyYGlmYtyyAzlwXlxRLOrnNlW4fMlz1+gnVHuD3z5y7U2eCsM2TiooiWyApx4ej6OMz/sjS
0NgrZ678OSnOyF9FDOINYnyYY15tP37/UL3Wm/43Rx7ke/7iIPOgRfVpvfU8bFsklj1IifJBz0x7
HnsuKogyf85CoFUaPoOna/pJpvJ+WAKN8iwniJ5ypGnowJx3GELZYyIm7XPvuHG7AkJzMVxGUgnW
7VonOcMGVMJpQckUQhdoMUS1FRh11jRyTVnXvshzXsAagUoPlugwzYAsM7c8h3zM5VBuFjLPs/+e
St3nZylfeVsLKkpBwwY/LGk93++UmLnjY9bVkVGDy4KFSYnb6VruSVodXuA5vEMNae4pL2X6tF7P
AQ3hUQQGsmus5QybUTAZEd/sm67HrRg3JVXqO7Ru6Nk679bDTPeCpv5WRUgj1RDJ6D/iSaani6Cj
wyq6sp4aFkFsB4PSMTRGOE+1wpJ2/nQi2pIYre9Z1vnlqK2JEZ2vLkpNX3ihtABdYy+8koXt6PZe
oTjsfKRaZhU41A4rkzm8eXrInHMG7idNwk5QJbFExrXXaLvWnWjcz4WsDnRJQgGdWOyXG+dLFKfK
G9rO4ECIrehVw/f7QUbn78IoAz0GcKiTYJi64521viwZAje9p4NUjdfEq5xqLqy3C4jJR5fmxDi1
jIyqHQn00ywobxl+KK2+m7+D+DuNn/2HLQ+lhFrnWMcb7IM1Im/42XWyrN0mOhzTXHprvzVP6XQf
bQu9AlqHgX7AG3UfgHx+TAFBO7TUMS6pHm79MzqDUcEG2f1QcBcwBxiohBAbQl4QCyvZUdZbtgM7
bqC6MgCcJhVgzbooRstN99lMjJCL+NAoaZxVhg7HDKpd5mICM+BR1Fw/id+wfA2wflCyZ9imdZH1
FUBzkxT0qFIR2KYC9XkE+rPRVg9s2GC8Fhd0v72fPDJXdqVmntxrHXeCcQKnUky4BxaKFAqfwNmM
tT2SB1x882CcGsqDwRsBQDIWkh1lpjoEQ2WaYIbfhlnrek1lI2pePiKc1qh/A9XVRhzo7tyUCwy/
fuPim7ur/x5Ge3CETvDPi2i+xve7jBNhDZSxrKu7Me4ccxzuPzIEkIP3yUF3YmJTq7m5/AOI8hEr
rRIUnFTQSX7lA4S1zP+WPCRk7Btt8wWn1nzjDDtDBdhrAeA5IamsQ6fGSbdC3szHmnl9/Pb+9t2l
6Zwf7m5ytDD8nppk5VvlNf31uebMuA20IvHVikavbEzi6hNZbyMSE9t0kMQm7jAqDExAQL38dctK
WQ3PVTk7rn+Z9IpxaFuXHcLtrAsZUkCQvDLwfbQHmRMC3D+fMsli+oX2M9ao25DdNhK5boxS0z+K
+SOavoD4PUCoypxADwqBB9NWQ9kbjgOblVmiYr6kN8+2z71PGOQRDaO55QTziYZKPKvq2jQTvF4p
Rwx3MgJo4vBjK1aWLG0WSASoIMjAFBfkZoWwsYNEjIh5jHd2gv98vyxlxM/dEfnSiltP05L72s7X
lYQaCHsEAj8F7aj5PTPVPb01mk3nV4cRhTh+hqr7S39ABAvLdoZOkvvF9gKDnvY5kL8zrQSYswzi
AFa73S1peWlt54luicWP4uVztMVKF1kgtO5fpQq/weEHlHcBwKToQZEWORpl/j2xK6mscyjrJOFU
hMYpACJrs7tFk9vet/dlQItHMVPqbTZ3GBicyLeF/j2Ldq+eHGpnNipUM7NgY1SXW5/wNRi1L9Bk
RLEjTVfw6BCw6VuhJwnqjiNnNxsjJDi75VyHgY/lPu/U0I5W/LWlgZUje24//HwCSZ9J2nk/hZkE
PbztDJwJ2X0xIBEylNOt502LELR9rIIcTbcte1NprKyV+ugGDUTixxtF8TjkRiU3UZnuShlr+/n6
CB+Hpmf7Iy7JwO18et45wgdIDgnGZ7d0ffjjq/VdV5saZR6HxEs+Fu9tzlL1sa9QbPxmqkZvkfDN
7+l1X6WCQPnW9rEpWHbf5NWqbvQtQM5K8/JjdnyigMpJbwU0qVqIusNj8r5i5lWNF+dW4TJBZ/OK
1hAFAZNy9lPNtfvEnrxgPPx6HDHvIt1gKHaKxQK/bKY/eChg5+ZKmouV2QZ159Om4LN3aBu0ZJHY
hc+JlPyueE88vukdWWqVpiSNHUkWuHpCWu3I+fDK++//9/a/vwaPceeFqAXgLPbyKwpPF2PFiIvH
QAriH6qWTaSiS3Xjb+B8Vz6lee2+EYQ846ff4/r0hUYypm7zWqb2bAH36tnqCUJKbnCzq2gkx47P
ABWSKXbakQLE7DjSc+KV2xyYdcS+1a2J8nPkfMiQt6CExe8nvvrXAfr5AVp3yrSZL+eDXPEqE5j/
OjNuToCw2msyulaU2y8hsHafEYhj1mJsPeO2DtZ6/7O47OAmlGHOholc4GrHrL09ItfEV2l3iE3k
i13n6VLmRNwsG/HShlnAf1aaGpapiYUAOxGBkPoLcIG3fbBWRSlLVvhPPGL55ne/OxmJVKuSh4pi
e828VnFEgfSZOJO5oUTKZy0O4nJKkrubuamQRHCge07O4pkJOfw+XUVQZGhLkuyxUW94228qPS+M
VF99pHz8d17wK0IfXW9tIDQyA3mS/V4kndPkGvkDLNKP9uKfKHlgu02CrNXQNk9fbjbWPx735Dzi
OX1IZ5JwGpjGcZTCXN3UjQafQf4w1O6p+N9BbOhHaa+Wuxl41Kno/76iVlch4mDO56uUFmdpxy9H
BnwPrPt9n8qAcioXRiDCfTXP28cL73200wExg37vLbXJcAYZ1kycNZwJn8wshd4AttY4y+pTMYsT
eOIcDJiiz7q5h3fXUcUXWEkQH2gxz0QpI/Ob7EFWwcbRY//VSIGHl1MMjq50NEvVtG4shergeaNn
8wtnBEZLwWAQ9oxM02lZ93bfiyHcSi+7dtWJgcqsnvqaPh+bMIEL0PVSlViH/6xdNL/IZOx3XURb
5OKKoS5s3IRUTVOeh1i8zW/I7348g/w1NCn9YNYTuIYzTSwvMtvwEONJOmT9RxeBAJjRM1rEI9KW
zQzjuwhtPN4dAqRzEs6RV1aYJD7RZVfTlEadO2vDj1Srq9Ehij59ChJUl4Pnyk0bZPZBaPt2SMYn
n+tNVTSq+51q+jzRsZae949ylxhQ8xJNBQ1/5GnRgFfi5q+g/MASqnQPKak1CWQdSB3MW/HZRGa8
YhQanh1WJcTUTFqZtktiifdDfxO+PrPq6lyS044gonHdkhU4nj3hnNaFb3M78ig0M3v68Ma7CiZ2
X3ooYle0QDTebShEa2SwUtpWZK5hN1clanKgBVumqfuEr5o4ZVWPmCyrTBhEDl6lWYeLvoQ46LV/
3zJD1mHRtFg2Fia7hjKRic6HkJecRCTQuNk7JILfMtlAr0ymOoJ0JAFQ9Xox/oa2woEk85WS32Yk
WVvx7OuOepS7MyTMMkKwXegXGWAEF7QBafWIO9vaQVfmGuZspqr1fIR1i58t0NiFVw9LCk2vw0WO
/v2nEXejhoTKqMeFufsn2mLS3D8gSRMsLGhcmMBsE/gBw/hNCWDgFrGKtEQ2TdpNRiUY5IBkbllE
LAWGANxxSLjK5XY/zNQPFPuWfvxHR0hwemLLNx+BCqAWYDVbXyusqZHZN0M0EKHvY9jEK8UU5dk3
nq+ia5blKORSv3oOJuB0t4pZTMoJhVprQ1tEOVgtVLk++HUk4iyAcJ1fwRcaFQ4qJu87on2ixIb+
NJDjxbz8f0sJVWFiGszgBIYJqRLXHV0SwZKRi+4lT9nPhl+JXI2UGu6SxVNevA5sE2M/F6ESWeCj
i8xrxGTfP6Z2p/OTDx4cEKzEYk4izqHRJ6COVzhAwk1l3IOvQtlW/dTHHJl9apFwW2jjCeWDmf/y
s01bChAoftc67cqvLEsMnsKT44GeaRz2GVeKTj4uVbVo/OeffUJ/ieDbB8NRkIjijJ9FsmgwarI8
tSQxfr7WcrrIoPdd7esFxX8UBWhJdmc8eUJrEXaau4eTLQce36A4rtFUysj8zxtkgpmsPzJTCy/U
hTrV+GdIwqJ5KH8/9AyG4mWa0yEnSXMUr4iWJ9Kxgd78kK7pDB1lfoKnoduiSQc2D13y0Q/eD+dw
tK6+W536zejk5vD+01VLHZVqf3bxO2FljDzcnwDKQci+VOMPiqMY7p26qiFG4Moouq/h+kX7WHbd
6j0QAhkD8+xcLsK7+I6PGc1Z56Oq/rEiPNKMnb0HaUCnzEXkYiELl4v3nKLkxH2B3VGydM5kXzjy
I5DSYH4MIzew8Zg+QfhMI9hEVMuDzdMZ78rogHKdVE3WjGeynym9wV78LLJFEoli4eYZyL5YLjGr
fnLDnuZawV0+OOtaHtU92EPjPCvE6j+Pedwj6ByoLtv6PguBY/ZkvSBvciufQFxemjBv7EOmabVI
lUdMDTBWOxYyqG6bEx/PkPFcuR/eT26ikqu8BDqE3w1Yn2n7R1g0ri6zJIVAm1HiDrW+fawxs94Y
1M3ayvVYGnlLO5uQqIYTT4SbtWbYBBnrDc6UrKJD6y7bqzjBV3zAD4SlsmHgRMOJ9m7BLg35i4J6
VPDgJ9F/eHuSV6jcBwRzW0O6wl1zRMqYtvOcmC70MksgNcuku8PFzQRigVujiNclCYJo7wtbYDY/
GKKTzu5B0gRobeUjWsVcA8gcA2pVGVCCrIUqBM/bfyg4Q9Mwp+dTVXe7oXanvkGPjkrRdw0DGnS3
WQW71OL61oq7Y50jS0KEnKF/HYUEyny0Dn75rmXGnCQDuzElEucYkQ/Co2rYL6QZBGUBMN2Wv60S
ZLjEpSpoHN0E6kW1LL32bE7hq2tn4cOdHXmwxuWO/yVS+DriqBeM/bQhwpTNWKn/m2NS1Kfg7rVH
0BeCCbihcoFrAIh2BRS+H9Z0Z3pZ9x4lHTEo1lUi+4ajwgx9lghXeKJYTx1GK6eEHo+/UD16NLPl
Gu9xebNUbbcv1Ec6iclp7GEPpaLc4QsJywBCfQ4t7O8SZAtyS1iIX/UGOcWdG8YL07yK9biD+YMF
3iJ6mOe60astyNB5x88hwadN3JmleA+bFW2h82J1+DRBhjtJjYIiWwrWU1rilM/cioyFo2/Zsauq
4DThykJla7miZCKZ73egxiqOX3WDA5x0e/JcbvuitPImeIF40thaESGTWco80rSeahbgOB8lOLDu
lvQOU6Zlq4w76zTQYS1jqY+AMYzRPvfg7E2oaDYYx2P6PbbacfbRA68Cm73q+V4N+geRjtnQSM+V
X2yJzFm7O8aFGpiA7r7PLqk/Wtni+HNkfcFhFcaM75J89dNNUDDSOKclPLarum1mpqOOIdt0WTTn
G9VPaumBTC4eaAVt1WOEgSChLx1h9UkSNHRZGc23z022uPIxYQZTQqDWzD/eSLVG1TSlzhuOp/Nh
/tzoPlgdDP5WqghbASGbTqd1l6Gts1XCtUW/FCFON92muP0mdJNLqjoi4OnFwbK1j2iKoT3mH3VU
sbg4HoShCBXsDp6r4yQjX+HAAuLtS8/eYEIx8vGPZizL0IbbAzCrtE8663ZrddJyyjaR0SjHN2w1
eKtzBAuh82FlZMd21VPjwHTgPF0d5WS9/3PGNEE/sF+TmaFUUNlh66RCidToP/hCeTwAWaPJ1tLf
b0eKGdZknS6IM+bYSwWfFA1+ZgXwct3+7tJCSlaiBqKssqWOIrvmF+UzR5fReU3w/gRn13ePabgF
bgLmmZeNS+/R7go+m62UVgvM6//JZ019kzlOjhyS1M+f/9lO5A9uwfkC8q6yDy/j/KZooLUx1exX
7NFdWKQcQFImppBqlJ3+wyhjHXYGIYkgc9/Fzac7DjOPfwxkVJc9xLPSedjFKpGmWisdFFxdNO1Y
9LpXNug5x/Uq3dSC+hWsSahOMVoal6jZFYand9GFxZNl21lhKbJbp1KbgutQ+63crt32JXkEhuWb
X+8X8ilta27bjtoAq/NPZJzZD4PtmVatVohhLS3DNCXakzLsbLiOe6qM4nxe0Sinxgw1jaQJL6u5
oF7d8lNdkLKsbtIP2FWf/UydKC4WVZHzq1F0DxG1KM9lZmMxtil0mUhT3rzuToIHDYdUIU8/DnNt
NVmE7bMX6Ul/I2d01mVKulSzfifk0idgEz1aVyBSZgo5v757muxO36J/uLGWij+/Fgc9xxEphvH5
LB7OLaB6ATncp7uPvr0CwwYflFf8/iaEfwnfxWS5Wdkf/xYKuoJYv6Lt5V5MUCjKCiszi4nYS+aw
mDJj4PjjqfwEwnw2u04XQiJpBMZFJEzJxqdwQS9g5VecszEhA6sXlSRaj4+Ty3eun5hyF6QpycI7
8OawuBPaAoRTGwScmWJjXiLB5mCpntpnMBVAs6qVHwlBnFG9Jp0lNHr2i8N2bNoXS45FAtf2pdO+
YstiSTMaJZzUEc7op3BO2KCVWJE9X9BTJZxEu2k7zJEi2Jzf0sBqr6yJHRjt/kzB9xBDKPEOomqr
nWxTSA+RBE8TsO50pQfnSqzqxUzIIjLqUjoCB4yCsHAi0gShE2ScKQvVTAj8ziTHIJYTcpGB8+3q
9tN3uLsGNGFMuHJrorg0mNgddjJ06Xecup+BhPSMoPRF05/u/zSgEWOuWqgQAlL1WfZRHrNY4qf4
CvbF2Lt4a6DZQO/WcPjH8nfSgdFYvSr3T0AFyZlEAs2Yc9m7Q5fjVe/1d5k7NMTe5KukL9P635H+
RcmroDHYIbE7PvZeALYoqF0m6V7OkzMYVm3A5XTrEA8Eh2oqZehmTkK3owyaSamkaklM+egMdu94
ph6ijLczS2AcHtvTQN90Kh5tb/8oxOVyC5Fn0FNxMFfwcszzIzNiIylPiNEIG/b3G5jiW5gdzO1G
5wMCXmVt96KTEQ0bd5Swu7fumZE5NRkysde/PWQpKNQl6NfyG6vkHbJi2BF3geTncpfLte10DROI
yNv4mls8gEolNxirQB3Awbpda/RupZAIOdJXWReOWzSY8WTCUCzU8yn3jP4wjWR6byJHxtulYpzN
uPAueLAVxOGKSRfzkZXj8b8tlYm6bzoxy7xal+qWOp+v1v8BIzep9oCwSmh1MREiILZ2/HNg/ZrN
/NiDLLzRlTRetkl8sa3l0vW/YuEGUzxuAL2U5JIcbjFxm44BEkw5UgoRpwXo0uQCr/lH5TzF423a
bORd2AkwbPjoIsyrytnrAfkLWA3u/e93PZrary+qfjevtYqjord112r0p9+9B9MrDGhpdgYYuJQN
+WHI67hPqIGMt/6ps5Kr+bURzKuE51UEML6hE9mttxBo3FCqvNil9TZWX+8LAIM4YPd5UlkwZY5/
G86l3HmU/HnhTxcQJjqKmSZ98WP6Yf902YAjuMrxIeCIIl0Hs5CFhurT9i/raZLjbbQzSLtTSJOt
paixiGjGX3S75awnngeQhlx3pFfLGL6FpOgVSTvS48x6q3oL/YLu5c7WiEvx2V5Ati0NP7/jBJLM
7VSV8gkzsO9sgEpXnUTDQc4kHLyr3tSNNM0/0mwF5un5VQ1g92v2gQJf4MdmLQVj6sElt2hyE9b1
+wvV0pqx0dNk3kTdbcGA7TZiioN6oVX9vGhtrSo+KhLdSmF5Q5T8jqKsP2ZYmb8yVa/OpFdEgjKt
7wMDQjKAlia700zSYBLf1D/YdcIhqcMA3YudNstOaBquPaL7wiGICNQtEpKwyJMt9adDHa0+TPdc
TgxbkLjD3DZ0teLxiSvgi8Mf8WOsiv7HV8H8cHvmJQHI3IFNP/Q/fyJ8QL0AT2yS7LBFoyyPBmQY
kq1VCdQP5CiYCb8q0H1q3s+foD6plyA+32L/4hU6+T8WmAhdKULHNVE3/JmK7s/NjYzPYFyN5oSP
G4G5aHbdtkd6yzJq/FN1s1jg1aKoaEkAES6tUAzqhSzlEk6lGpMlwrVwR0mepl66jOvFKK1FV56V
SyvjLgv0ZlzGjvtCguuRfY9rqnVRDPYq5imjMqq02MEOjhjgzOBafhQs18daDMX3KZpQoYTkffvq
PdvN8cegd8xcrxnZIsnx3Mf6euvAGVJ9ZGt2J0er6O3VN/bjX9mQs32AUozCLcxRgnEv8yQWOnn0
Yq7Anl7LgfdeJXRNYU5p1XHeCF5n6LN8debsSnO7A28hqp9k9NG3/BgwFiZTTj1JC/+qc4g4cftN
Ei4o4ZJiYVHHPuJMNw3HA3U4mZjxX9rSUrIFuPDBli9MjYp/gR+qHw+ufu5sTDWB/fyEh5eshfF+
+ZevtSCrmFkBtfrnp9sOmqKF3TGMwJnpOPH350vnNFAvMMrTWQoZHcQ5odYAMd0YWC9RZHSbYewp
8lYgt+BN0dAxVXr3dfr0uueOqdK/D0DidubtpwShpQ2klohDDc8LDiUUIA2nd20P37DRofAJd/sc
jtUIuJOpadkdhEa8ogf5IK6pyqGIQAOy0BjbXUhSln33vam6czhduQKB5oILACFRO1dQaIKNJFxd
C7R2NzKteQaUsZ7p0t2ox4r6cNfWXIjGobXmYbFdz3QL25Uh9TTYbTkKlhKdvMXupL8ClEmuE+eF
zaSKtwxbGLxg4e+/UCpBMVKahmLSIm6T8F2o/q/oY9HHvHk1cTLQsDOa5hAJqGhjg4SJ7MrAyfZw
VqeUQ1l59fILWAj3aCwUTARhPbFCxfFcArH7MA+tty/ovTF+pOK7UfuHb1w7XUdTSyX64qOhrIGt
sB69ch/f6/J0sg8RsxUKxv+/UNrl0nwOe7wu8bFbv/FYJybvc4CikJ+eOgLkaKV1pK64nAsNRztC
0ZodjjZWoggYDUQ+JZ2bOPF5iWtitptbSv/MP2ON/5G6OlbmgzncKLLIYwYX0pmuH79VR4gVH8vN
rRC2P5HHa94eA427D8yPef/+OGTY4dpKwaF/uIkBwp4/CCvAgsz0m2zzgmzywkrao2A9YSi/z3Wg
CeimOvQkyyOUvQT3AWEVzxtd+Ku7fdBFqT4iQW55aYhB2m9dEDZgkv0oRiYqB58zcU2ZvsZt8Sjl
sA3nXW/9QcMDkMotruqfSvhPh4fBtFfOeKcbOEDgqRsH8TPrMaiRYYGNe9u2SMnZd1cWORH8vMWa
WTFNK8dWY1fKJgBu5KsNbCyquWF6A3TabyOv9IdGTUHJ2T+ub1SUv7QdABvKkvjCQQ2i9VprHOoS
NDvQdYH8ksw1cnd+CqgfGULWPQZOWQND5xi+J0AordagTLESFi7PTaSl+vCcFvp8u9zs/1AjEUbI
awdAA3tvG5WZ1QAHU96OQKSd18jwaAcvGOR3edtf6gpOD8fW9WKPTTlDq9r+Ews/C3jmAF/y9KTi
YhWrlUw7ynQIGA+a48A7/IyjmuK1Sj0Y3ug8JlnxqozgkaW1Tg3ocBMQupwem1/yAvZUPK274u9C
iJXUEzeMggwLqvsvvo1oB1ikZLKNc1OeoHq4m8kuM9xbxoonyMZjyoB7dfgNiwvLKAftIcDoWw8F
KH9VeeWDNmUby7Xrs4Bm+TM4zESIlDsGo2vOhT3zRs5hiv7jNPInB3L41B0DqqcByA5yImXCxAmP
rd6EBGssCtR5BymUxtCIYugafoo2jLiDSL8lp4wKWq4vpEASi5RqrryPQ8Ll37fMr1m+ZzAuAUbM
pZdqstXIFnUm9ej6LPG6+yrTVLO6LmsIKyZcEE6DToW4D8zJ8WsDfvFSHd3IRW9SwguSgq13xKLH
3FZUbLUt6ynCNLnBOCkqzTASENc0I+qZii7YxAXaUor9qP9d9ezfVMJacYtapgxiamkOsK97NVei
k1dZMvt/x0ZqD7mHzH4P5T5mf5TiRGw6IHnHMECAjx8d4pJsAg3gBqZ30rzsOD+R2cuOu3rwuVd3
alXyZMSEyJD/1EghZeEIxpYx10t+w+l2Vm6vmvWyUiBhKj7zpscdeCGo9fk8PbxwEJEdH9eSC4kc
FuMX/qBm5Y3ICRF/nKahR0nAVZcHo0k7kzwp9HYmXFbpi2P0xQ6w3wRvoLKaGJ/7Kw8ui88zKxQO
dRS2yFNRewluxzKBPltWrl5GuFpUhssJSz5wapKxjpgdlPHC7ugynjKSeBx98z71hVTwbUdlID9H
HEiiCjdWkMhYRsyx4mxgyeOacjVlGDrxOHF5wXK3Oyk+zHQr+k8B7SL4O7WaXMPEtJfQvgFubNRM
5KH8i8vJlg+WIAVfisz7XSoF1mz2qpVjVaPqR5bFkJFD9wVROh/xsAjL/JOFpJ/M/AaE5HZ3ITCJ
2ZySN9rAa321XyT+7ZobKjZlrv9PI0YKEbm/+PPv3cU61FBLp2QV8zcKdjumP6JN84i1QvS+JNsn
jkPdLBSxfyvkt4MNJDSvwhk9rjEqtV2VPhZUwrrcF+QmJ0goYbU7GI7dWShfv6XCYaB1SVNlhK+E
c+tR4NlyTrsSH9xcjAE0+GPqyUqFOakXA5Wv6EYEKebYiIGlYM8POSOHng032w3z2wil/apJ5obg
KOjBhkELKbRDOG7VHC9/3LasE/g06sLic4w2M//rKAvfsl/ndhNYyiS7XJ4wHZ7HVV1krnFsGNVv
iBcxTdeEUbWLVQwhIuMujphpJnJF7ZaMlGiiGjxirkS5gy5VTXGyz6L0FrlQJfTgfh1JY8XN/QZM
WiWl5dxSyYV69bD4DPdrJFno9Xvs2iAQ3cmGgLcT9ajnycYqbHnLxv64RlXgxK6ReMTeP3hePjWv
A9msg1hABK1U+BRX7zzcB7U5GG+pD4p0MLTnSBR7ZO9s9sr/H0DAtPbI77gmg4nW4coD1X5snJiA
r783Vi4iamaHqDZ+FkzNDFB/m42cfkmudOvm/sGTOSgzj+BA3WBLlnbDJJDq3w32LM/HjWSAHgLR
+VB80NHu08wKP/HFFk5jJqeB4I/qIuCjJSX1kJnHIH6qCpSHIxUzNKgfp39k+85Cju1/bCkzGkvE
U28DMibVlnr6qs+GqhllFnncHSodNvpFtUkrZzMELsoZnlhBw0pJAM3CSqnjkPyIB6xvJfHcqHAE
kSWx6HdWZ5PmO9ufaJDZC6hvWo2za6Pcq5hBscPCoY2UXTBsWHk3WXqjSS0luOJL3t91P6SJmdp7
wmpmPF6ZQkQXNih/O0R/A27nrfb2eJ+Q5WOLehwe5fvKV9UE198VjtSKWzIS0KZA7N5HM+4kz0vK
zDKe9l8LTK7/8IeDQi6XDSA1OepOWcQAgMdsjqsA32fkK+FAyc9Sh/rLg5Ij507bwCyNY6xVvzN1
Hs2Q4vM7DAlekwRxHHFWMuJgMDTccjeoPE7MmYeFWP85XAgaE7WPZICn6dhZDKhJ2fiFVRMBBIJo
ZpGq54o5B3ttqru4lOl7F1HUhAxr6I6m3wpsEmz3aHep6YzZt7zVZkfZoF69tQPeP7qSkW8gplbN
GuUlC41riKple6RBxRPR1/Otshhs8hHXxqL4pYuscZukj+46Jtx6Lcu+szbhXsATTFGLnwk1DYcw
9qRq4M/pjzqaN3YNobdlzVbBUmYc/Rhf6HMBWVdi6fa21jiThP7bC3lrVINdurHFKBSw5ck0kmA6
JQ9Hpdv9vA6JSd65/Ayb7l/4YQ3btpNqYk4b5WIjVYZk3Zmwih0Ze/iCshoVZtfs+fd/mKS4/j6y
OjZaw6mvJrWIPgJ9KrrXlrr21m+zuW8m63/nG7P0NKXf3GcAT2172NlmapPDGNEQSQ3NJ77+X9Ls
TU+oJypBHaaYIl231pffHW2+1zbzG/NZNjh4qVdJLcWqymRMBUuq2vaK41TRqpKAsRXFwrr8C9WD
VyNaUnkfe8/2e8FdBbjDe5/ForoSxb/w2fkCLnKE/eM23bPbsikSp+awSPfIKDX7hmec9QxspbBv
uqHKN2cEk0zMdC+5uM7D0LVAflNB5j2leWvg/tBzNuReuq4XECzmn/jXMMUXSq4uBHFhFwNQx6Y8
f6/XM6+B6vji7a0wB3K0sS2BaAISS20XWR2Z8nNlhDIrcPyG7ixRzeG5t8DqbHGRePAzO0uybs2f
mfyQf0gXQG7NS/ocXBifRMPO3WwzgOs/7rOgF/D4ZKUqUIyNjmwxVd1Rxl2EsxN8mecuawKO1koW
rFJSfkosQyM+EqEDDIKtc3SHVf7XOfApXk5dl+cV+SGEOznai+Z1gUpY2rdRZlGUniqdqx4ImOPX
EVH84SYPBXt+6v2gmJJZnHQoYOHty74SD/L6eluSih/lwoxtkJGoD7BTIa/whZos8+JKx4UsWMhU
ECoIJIVXLMJFRfNxXbvjD6OdKF4mMb+YppLx9rDtjPjnvhpJGCewNrGRIhMdsEsTzu3OE857+do1
I/9VFa1eviyLozyCrJTawH9CKigr9d5jzuuhARTZqBTD9NUW9pnm7bUikceZ/bXS49YjiRudSV1M
tD8J5PB4y3/Ufy41V2rleRCfYG34fY53AbWKBA368kwXU6i0Jazf3WDx4K6zm9+HVBztrV6+oONT
/1A+wuhwpfmuSIRIaTrmautc0LZvSl1iWTxzXjhEy0Oq5g4hO9kaQBoCkP+QIkMVNtZ+k8dlNQDO
EB3AtUTUf8gy72XWAxXjcLtrJpUxtUoWXleQwk1Zf0IXJgq0zxt7XiQo8cSUSomzesLfBG62PYp7
Z5cEyjMjg93Bkif8Ix8RJzhdQZe2OA3PRd1Cx5QTlNlYJprJUoWfAGFZr0z0LYWBkCPdUNFmKa75
L7bbmtR0RuD+V0SW0inAe4na+8l5DPWIqYI9Kuko6nNrn3SjpewsLTmT57p8WdASNxGx+ZTNbxkN
O2qlE62BKZm589w9TmQ5+seomnXlugzULe0Qpyt93h4PAG20tknlleAqNtsgOkyykBPsOt0Njzjr
0xT4781nEmwhhUKUgzd4iXI2+GsbgqpoZ8NxAGo16SFzqRLaVVyWT+M6sISXsQZoG+NNWx/CAoWD
qCSHCDtYcx6fNqCKcLWU1KTf1WV8DW19me3E1AbPGR24s6RdRP3V9zG7lcrGHOW1SrBRHa1myMLK
RrTiUT6r4TGGRCPlQpZY/Z59j0bfBVDwFCQjxdAyvbcUST/sQBcpoEWUAeTlEkDDly93GvMOS/OT
ZFAm7vWhBFQOFw7vwURvsgFGYsbcqa79jQSz6BYGTfCRKydNkRt//td9/M8M/nt7tiDSu3+8TurV
rIt8nIg9Pl3JYUqyFWgkTOEkUsvx4RRo+4gwbJQ6p+S1J1JYs0eBzZn9xxgem8caWE6Ikg30H8X2
LDvBfpagyMsNwWzOLCOdz0g9qrurMKA6E2FxfRkgJM676ApOGdYUnUGszDYE3WE3L1vH4B1bzpos
alb8tj3Y7o8n8TTEmf7CiQSIu7/gZJ7JppPEx6zFax8KnUNI1L98vLe7vnaHfv2eoPL5M7Ol4YBw
on5NfYSr2GB+EbG9VG0ywyP0lvdfaG7EekOi0f1fP9MrWul31BnffWZIg4hX9iaPNEABIXsdU4i1
hgrEf6sxnsIjxRta+bwNFXOcUparLENhXHqrdL7tcb9+Yu5kgM4gjkDX+7IEuvR62mg4ahCBdKum
QlIiLZjCo8q7SqD4kEQcczfz3BNaxdE2Kfmg78wiMSjZuyQ8y5XRLwsYUi+agjv/+RpYt1ym55lS
r2zuJTgNF9cVuSnkezxFY6Ze9L9CqyntS2GL9KKzzj+tokgNB2vi0XawschGX+kD2Cl6VlNQV5lh
GyAqZja9xGzIQ4oq7kb5PiIWrZZp3CMJazeWZApKOHzItS5eD0q2iJP7Bn8MYY9F8ZQzQfdrl+Sb
RxvGQ+fly18nAKBf1xyoWHp1ed0pxPbnUjKihut4gz5eRMUuBtofv/hLMCr75sDltJvZ0vjtUs95
vp+Obyt7RZbHVnu073rlODG8oByCECNFt07rhTxBxjI4SxH9qO3qTgCKaVSqX/HGoAIV2iPmjHHP
4n/lUJu3BS2GxpvlkOaKF48HjQWUCpYqNERUCmu3H2MSKqNzHDC1kieIqVRtMgWt7gj9I7Scr3tu
dGfWz/nOHssFDDyG75zPc2rqLXGjqF8M8C9BkGwfTCL22JZA51OImdYo3t9E+d0GVzf4bZfNckN1
ev7zUhXjVwDtSqizvecRUp/ncnqG1Iv/jFh3t5D2du0QgXOnPVvvGVnQz04K+AAJKFkkQHRsAygK
LlFKAV1XF9UcVfet1qZdKewW9esQg9YPwct9Y4oP6MHCSXoZB8LfdqrOI0b6wd8Ql/gTOZvBNJdr
f5NwKOW2R4e3eSCpSbbMgOTV82mHE6fsOvfqPJX7w2Pzy9RjkXvyzCxr3MqYJXeMg9Dvt88YmbE9
hxn5Ln7dGObkgNEswyJTIlVsmW9WFGsW780gceq54XbSl43hKksRgUqGzgvWU3/7ZxiJ+eEjomLW
VsWJCGr30sGdtSZkn+LT7CLKtzPUll1vAOw4Jv8TvcYHrhFGf8dEoIq5n4+roAV6f3kYiT3hVvpV
eMy97CpEnSokGFZ8uwxdDwhHJQi72hvyGQRASt7WfknAHrcGBOuJkwNhNza6GnCpN6zr+aoe2UUj
4LyLpj2SJn8HEI3+7TxjDvLiPQrbiGRDMc4jTWBdZRsp4+gysxC/2VgVmKmIVCAlIXKWI5BI4ZtC
lq2PWoolqKwyVyuKc0n50sYOoqQJIYG2Ey86fsye0M1FaACha2+572P+ah5b7QhmF3iqcndG5UHV
LG+7EVyeLZEhXTJdv6ibmrzszGmpMXgt/NQRa20wbNlMDfscIVmftfDzMba6tS0AC1ITwaHRYj9U
kTk1YSxRlVhlq5EsbC7v9hKKnhDaqcdXdZ/La4Ai3mO4ZeBLMYgtywLtPQMk+NCL+55m+atdzW1w
57YYkZ0/78S+yaojSntJojy67lFI3JbU4qoGqW+SpQeIp/xvvXaFJu1BBZngJIUk7JAfwTgT9sWD
hUDYPOv5y2us44hNPhq7cVkPvzxOWp/PJyOTGK3HCN8SVGg83HrrF40mxrxstM/O8F8p5fOPm0g4
LzRGekYvoe91ZMhuPqpx3BJQvIa7mZ/KajpWywDMNGQn8qrcxgYfZHPvAfA7+v09jPqcxaBkZbST
FvQnyjcOa9YCkDcxR1PpzB79GpResMjhiU87cGbann/Rr/f6T4DRnKTvYmYPPURpbklS+n4lvm7L
dj/n3yqkj1Pbsz0IjX6NGJyxRt5wVGazZu1vXYlz+n3yn9yzC/96bfuSzf0psaDu/lzW0fWgOiTM
vnl2n1X+MCVPdy5u77aVOKdRUPVmn/olmy/s9p5RKrJs6af9xENMmiqqEZLB+ZguKzqf2EhVkdSr
jO/AkdwPmKDyG2ZWCP1yioK6BXG8mxWgVUaQzEG/3hCFj84YiHS2O1lpbnUY97yc9/yLgFk5dxx5
xJU4r2lzCWTB5xA+xV24v0Lh2A6qnfZq0vdoHeuVC2A/xzhSbI5Mi40u1P3zYXch3C+ZD2MZZKrF
KCYYGgNp522dTu/rpzklmvbGcRYO8FdIY2GDpDr7DecMuUqW1neKYtB7Q9zFopRAl1NkKOs9L5EA
tJMlhOzj7BKi2u+WXlrzbg1zLwD9Zgt9JOgUMKbw/lrLLjwPzsSjbb+afi+kOBIsvkv6VBKTg2oO
7Jn+SBSFnwuzKLS5oyCtsDHr7g9hKVQDOdzI8BdpL0onpJ0/+ajGoyxPMXqK5CF5oTFAiK2CvIik
e3+FwogXctUwYk1+LXAnCi3gQc/5ELhFMP++OlU5OTW20QQRCp80EafMWaRHxumAkOk01JaUNSHn
YgaTYQpr5WGkEumvdrKr88FZxVbedMMUEsMazWPf3O50dxVbwq0BBW33rVGaCw7gBF00EhUnmlmF
k5Dcn74RLpNGV81O4+brm5/QMj0CmMzFUu4Ssj1wsUZk4hffatBE7C4dFjQV+i/ZHCFXadKRQhva
C0AfET8BBgHlIBmGe2QjRFgiPKDF1/IbP2cdvbiVr4/Ub26MlFC/F5RUuJsM/jFbc3KWIAAoJdrI
r62mDsQQkqpK4pzCEGfby3VJ35VnK/L2l32g7NPu0/YNTHuEcPFpj9FDawcQVE9I9QYNWt10cHFi
VLrxLJMSsTwCzU09COFlCHbAXRzKDCV3kFsJqT0KOrCVCHe5u3DONKymWUzjGY7goTA0HunPMkIm
KN+osx/+TnnlN3guYU3Oc/0zu/nPsjXayWhSpsvnDZYDQXgWHRaEWlmbTvPvUtgeNEcsdUzb6g+A
zI1cJWJRJ3WQ+6eWP47a8QCHksIw9C6hlkR+QnwBHNcR3YCPZ+Pu1LbLNOJ1FqOkGqdXLsh25eDv
K6BfE7imm7Y+w9wYARo3hjPd7HGmgA29R+L2DwBAkuEtW+tYZrfHGwXQBitpgYQDHMOoamBGOprY
NJg+IN9MWQmdPxrRX0URwbfFpEw/9nT40L1M48juYz+nKBjIEXViqo79JqPmjCAGGa+B3kpWWS8B
DKG4HSEZM4LqxtdXFAjCQbn6y1loWT6+dhkYVSO7QU9D3uMofJL0ENkWxPzzNFzRELYFY/hU4PDo
q5DGUerk3EM8x2fJmXDt/lbABMX5HloLBbaiEUaCwl7pcfFmq0ak+2lUuSelt+qgyLb2GdBnyU5X
jDud8lgG51fqUagnK4UNNTgUSPtuQRqoqqzK2w+MK4ClWIYCNFl5Ox/D5ZhWgYJuoL6hV1uU+MU0
VFApZBcJkl4v3ELZviI7KjraTUC0JVjAZh7+dWktrtYBHd/M7d5KAZnzq/RArgmiycVLGFQbYwce
eU36aaIBL3sdDnxS0YcnsGDuEsnQ0JUPGvAhfzPYIhMcyjwFy1/fsyhRTpv9bh1MqMYtSXuq71b2
qMjP8YeORwNEquUMm7s4a5h1S2c4Yxe24Li6tzqxInSSHaOvgE+BtXlLeDZslCupERx8KBPw0kmH
OdySrtDE8gAovED3GO1sm7Rrn/YIZYtNlGgETC9tVlqNHW3b0u24PshysR/4OSetD4jCJ/CN8Rqj
ktf/dW/rBGLsWrppDmTvcYs2SyoXVxdOD8Pxk893X90mK8dUVWSoNai97ZV72JHzP3nxGLBMuBmq
TIDlPA2vfxl2NoxEgZ2jd3NSagQwPRe1mAfIdp+iNJYrJtDLB61XB98V9bqcDIzGBc7MP0Ej+rAu
NfxUsM4oDZzVHoeLZ91TZt1M0lUTXcnIuQQ8fvslr+qYKdR4ui/KUD9xbsJ0NDYcnd4XiY/5b9au
ZIb8G9F0vvNyPm5+YRcdwlfE+CiUAiopNoVAgRmPcw7IpQSLzHqWGO8wpwQva3tataBX3x9J6IrM
jFY54rX8VW3fWOIsXl/Z3z2XE5KEr7lvISZAdlkNXPw/26g6xtKAETee0vsmHG6scAGJH/cWa4uH
jisalFKvjeQH+nOrEOjIsLu1kgGnMK67knt57yobNxOrZqeQpemV44ufQRSUCKz2TrOhlUePAOra
zWMPimm+tEVf1P+hIBDiYpEZcKekHaoPfGp/DvuLY2P4SaKHCziOYISruIgGa0Eosmw4UevYNJUA
k60bEk1++n6BUrH8Z2+h/CGbyZr9q7e6JUE6LAZrtyg34vHvEnOIJRIDhCK8s+6OVw3+TDSOsL5W
SSPDn73GnPh/YUdG04l+OlrloD5LJw4X+9Zfi4N/hI3wFosxpKJyDybJZyEPKPdeA54rarAbEvlk
VS/8k0LNzCN4cDpcb4embz/Lu1o5Ckdor6pJgrid8HY9bWZy33edRTcgdLotFxeUd88wUz2Fo/zu
pDrm5XSa+Rm8WiiIC9yOEvuFtapiAhL4xugVP04ea2zqhqtYJWDtYHuG2ewYTBPqUORCR8ohEnVD
cMtKl4hq7A3/52IajYfQ0PbD15E2KxUbj2UBTFwi3/G+f5xjmA6WGPTp8b+TJiVCAg/pAxNhevsY
+r4zTOX0inwOSBYF03sChqkZvL/Ip7EjGshE9SNBSZTHUyuRhWwbpR+Kna/b5Eme39SIYuf+PNeh
VnG1kPefTm1e98WwCKJ/6QBvq7nWpZukYq2AuimnwOIkY/m8Tv3GaGLeqs9+hLWeHvY0dh75/4G5
tKvH0CWl6nl4dkxHeQTiRDoeeOR/0TzizEwm5L83To7EqTZCuGC1E4+7qni/kCGQ8z0KZ86wankU
h3ojXydx3UQ7WjGhrO+QX7Vr+mmUzbxY5maJeWTpf+v3s9dBbNo8ZteVHR9vWhAkOd4+4qV4ltZj
DX56mDXWP956wgewo1Mb4iG+XwP65uNy9Om6pEWiPXvui+sF0fL87P2GTLWZtZjsBTqD2/lhOyNw
XeQI/nlKAS/bPJ0V47PWoO/NZaIlzpZe0przExDvVQVR1BFR3wrwssOpRptDL65IRhEmVr534j0I
kT5T+amCFxmrPHpHuzSyqcl8ntQZfMXyDp8V1PEpmziAPrFOYpSryqOTArXxVVq7c/OFhm5nnyKt
u1P96F3W2CQl1CdhHLkiTHdLRV1/XNUPY+z+GwqOARLbIWqhy+gXu6gzs2i7IywOr1IeTJ4bNC+Y
0cSvQJPr8ifb1vUYU4Y68G4ytex9TrEBbwUOQI9WEmkqKMCW38FjbbH7pS+gaycdGqgWOf3z/MRN
DHonr8iNmF+8hRU92SQ1kTSfARZXwaVDaorV3OBrFaMPSMDOF33O0h70/I5mNtBEDalHiatAlKCR
uAYSZSEf+KM1HFC6xOHxXnDqruKbrLxIYwMPHru5aKczH9lBQcthIYMo4IorYdCL2ClnCDl51zE3
cpY5zZEvLuC9BhjNTkr5ycx6qhQXl8R5oYySvm5s2PB8/ffcJ+YmyCA/vwXoTHDchwq+lCYNRZ51
hmH7o3HfUFlv6QG9UPcqjvr7SMz/TWAdU2TmjfD044E0hOsjcAIKqonRt22//IzpSr2CwTdvvxZq
/lzMiUlG0nDmDNIhApe7T3QMtxXIJzQ46MkWZDwHgfmH320TW81/QcN60XxazM0BRdA1RMBC4Ceg
ZPK9YQkejohCWNyWFbrAteEusFEZiH6bZKNkhmqeO/El3iICigoK58h7jInEvpGHbfRsqnVZXEFJ
MOVjjHbx/7SrBv1yHzQMFYayLfi7/q+vdc/WSh+EC3269jSW/90BCoX3AKsBM7uShRQE8wXKo6Gc
fgw+5zF0ylhfi+fkF/dgtVnoNDKSZBorCjLtfTTj88jjaxRhckefFWzEAaIS7aSJCehSL7neeHBa
8SY7TcuHuWgAuT0WWktfIrD7/61PBiIj+SVQP8fy9/hNilrIVptuY2NEe/Y91uu+CDWdsAk5cPRF
yf4GJTv/vPaq8cC91UlfpQn+OqVluTPrHrGW+lrkdBol4QyipdR9YYRulj7iGHQfx6BAAFUT9trG
Ud2vT0T8UOcyUEUSaoz0W/Sphi3jKleca7FgYS+ISLuErbI25Iao5moklw5WC7b38AQtGjcDdAnN
Pbdx4VOIyg2GXRb6FL/MBDdSo8VzWdU2N4rCVg4Llbb+8R9IhOptumeTHBMrDkhOAvfXHPsIuPxF
pUekc+3dmzg06wwCLP4aV6LGSuHR4wqHnjJi//QiLy5Jr7Elk+hUAulo881ldZ18BbF6TW0BdA0L
0qxsvRNe3Qkux/OlwYuZSgNyZRw7NaTdb4sjN9wUyGUj7tl7Dc4kZOO2x4L1tuOSshNPlRFkqmx/
Ew5sV9wOXXCWctNOorwAKM7jfvzWjnWPJpwNH9yOziuTwrJpYLSjcl2yjhcHRJn9QDz3+ret/0ey
W1sMKx/0fcR22dokoh3VTwALSouLV4khvk198w+ub19gAD/Cf5XFr9EsLKY6LqdB/LIvV/Mm7clc
r+6IrtjKfHAhfvpQvigWmBsQh0J6m2BKissAxA2990IM4oNr2367gT2NvW2KeZ4LmbYFP6sCbts2
GugpYrHD5t+OWEi2GiGa25dZfCDkR1/BuaD5vJ+Nd76Ec8CT9+kZbP9r7cOjo7f2PoMuhpdmp0I4
2d6ACqJNniz/DtPb8XUtrCGVX9mH+uQVzzwmhdXgCuIx7Riay+dweMaElnx4vf0glkCig/xcVSgC
vQff2NcoCYhQlakYqTz86NI2F7Ou4Pim0OHdNCxFTctVEqCbWFyu9eM8UktGM8h0cGNvJHa7xZVg
0BrmlvzVU78V46DEsjY4SP2lwVuiIMXkUJEMDdSNdjNHdOV8W3Ftvz3esuH7cCJsgJUJieaHIaEF
KwXg2cv6HpuzRliaL3TRY2XBOKk8o8fVXOW7c7Szdsb1dRNjrYiJ+KnIvKRmoU1lf+AYrWpMjUrH
ZmJOyGjb414aHaU3w4Cw7EGKeXpjnIaMNNQmsL+HR8WDz1QMa5hVkmJ0ZZZjxZKxq76Y1+YvsRr4
/stz4XUcIvmCWsacgbRX1xbylTTEsWLrC1rzYzMNokTfYeW639iVQIuFTvXGW/RWmFk+/R0OwT1m
E1uC8EDI/6f5VIvFDOYhq5daKdyC6KG4ngmI1Rk62WEXoMLAxzCpAX03WW4zq+aC82xxmz7LSvPn
KssMG6hPwRZ2MYpP4xKQyk/0+jTH6OUUE2+faFH3LrW2ayEPeA7FvvAAWnWEbMdKvTlNVucHiYvq
Fm5fixdYQezsWzIKfDtmAXOSnyxF1FOU6+j1t7kKcXwAlq2AM18wU/GVrpMy7823Yzy4qZ0C5ziW
znD3KR9WDzI79SAI2VERS8KiKoKx5rNXEvz9NXUSsgYh9phuDKDPyuAcG1tAnBE/t8MQz1b6a0zS
n49ZoW+slRyrdB0VZrdhLCvP+DwKL6P1BMN1c7f36MMWnJL/LLr3BzUYbdVvV16PMNLxd9BdJoFY
RHxzunF3MeztU5a7G26arAPuJ+SJmBnIaUiCu3DyKjf04qnvoN3Ri+vJt1fWLtizCnJCuHOcma7j
O8HIuh82Wp4so2ELXNx8yzLGMqxXDLGFdKJLc/ApjHJRmI9C7YnvOlbON7CbGv2UHLrvN5kuHV4W
q2tCJAf8BMfX/msFBSMUkQkVQl5dHd0V6T6iTUAa/z2PJ5r7pCwax1LaVDvXs5BPODaEH2Zvd4Jp
u0n50OHxfs8d63tGURK/1oJqfLTRVmzL5flOjMs5WykGqW5ZXUnd5y7GPWfag4quda+vi6e4IeHM
2XDgYQcrkEzU2ttodFfAGdH7tK/6FGBomTEHIAs7XAMUAAeN/JLUFMS7iKy3mdHclWGDWX37HR3X
jrklW8SRNz3EILOcox0rsfAWx+sWHgoOoj+lvCdBP3KAkCq1nN055c824SSVlSJ51qnERpuXt9XM
ALwCjNAQMq/Om075TLWErGqDNmrftGLaMT67ngfeXuvQg2IjmgXzIhXEFyB9KkvbKSj8IPpbfyTr
8aPZrkafuPbrLGD4sZEwhlR1h7weUjUp97hok8gAitnjy161gyQLVtZQ4FSbAZOxeiowHSkxJch8
iIVCEbBFnVIsW069KtH6PDPvOaKh2XFL5Us7ykc0nMTDAkgNOsgTjtOTKfeYbeWwb7eklwC7MikJ
Ao43/urKbD0hAvj/Q77aOn+zMS1ox1m1BAk3pEB0GkNgcEYSjLAy6WZDH3vYRy9I44whxJ6c6pts
4FVnQ5sHVP203WLxRicShGklAtw8+nzyCoZ4yPAxM2RmgVIloBj4Yq1iGETkJk4xa9zChkx5L1h9
xirBvvgl5Ef80WB8gpFN3zoFY8KF+zPJKKNM1J51h+ZBtNsYp1I1NIdI9S17l+ffF9XEuWhgAZpX
N4DOw5EYIri7kIMvfYM5HWXfTcV1OncqGq4KE60odeNtPAU3kcm0PueHFYhNOK6eYfeqAek1KxS8
KCAZ1eC5hyBuZQGV2tjhGf4GkjYagQAzyIsFGf+4h7Z02dd+ec/OXIjsn/gs17f+nEaEI8QkuuF7
dEytBlfwGYdRltB+kWN78oaO/EMn/WkARnXSCW4jkBKswXC7bY5ERWlZP7BEBipmngSOTMv/wbCN
PadcKC7/s8ZJ1/h+RyBGGVVt2ms5lCvPQKTLb8DTEhOdbABZLEPdoeX3/B6Aq3ML+0/bmuhVzR2C
R39cwLxu3fAG874tu89pp/eYynK2a32Ck25z+wElM1FUjuGcwUKAPf1iW4Ed7tJi+O1ZdahPhar3
dxB73GUKu4jYWWEBHL67klpMgK0HVqmhc0jLcZLRwLqmTv5KANHPuakaFtgO2cDYq5dOx3ho0FvQ
4Ds0W46H9lUG+QAbVS9h9W6eRDZZk5eHnaoUMvee7c5QlPddony00ZdHnqkM+9DebJanleJdsa/p
WzPTmsyupO+alemR+6eNInpcU+ObxBegYQ6aYRK5dQe2OuQiXtbuD9zVHLeFksP/ikEDmQrnmNvY
MGRPUn4u2w9qN0tNlo4oDv1NfURPCJqB7IS7Gf34SuksSD6KlonpHPde6Eb9vHTUC4vTUPaOebEk
9gtwzhIDHj/8LUpP2SPOTNh/GLQwe4lxjCVBOyl2ITjqDYQsFWfJTHk6xd1bxqTDuPC/f3/rVY6w
B9hoSNRaYDEfeOaP98yOfNNRSKkYpGT922CfZDKBUsEUZnm1RjW1O3UQ1G7/cRACXsCs2lbGDkOH
OSGq4RL28It9EjYFRKha+edMYq5XafPavf6S4INm2G0eqmvtVT2/AIGQsCtfYmkrWfsIE9XHT9Im
yX81uFNLGZ51h6EcxxNdFbCbWWay/6OfKF6HwJzDKpkPvP4Du5p6I7ys4V4CbICFtpRvWmmBNeei
RRntDp6NLkkIIWgfBld5/7LyJdBKWWD/D4pnNQW3/RrYt7+R1EZjhVyH2aHXGKOA5s3dYMUORs2z
Y5UjfdTKngFrUjVdAQkFeadj0yxSyABWesbCoHQBEkuiy1uo47QQLpu5g9XMCxGRkKFz2poL2OZ9
Hk2nukfntV/5K3SELDRY2aDwz2V/FeRub6U3nI7Q2DnAqJMB4SZRoE6jwlgDLbTnaQNjxR9VjNA5
5+OL4Xy4BNO5GuGjnTFmTveVm5AwblmTQxpxpQdIN6m+ZSiFR5v93jldB6tPaD57ydDCzJ03nsn4
kylvoqb9TLZKlXeQXcvIA2CNM/4YbVQy3m67JO4vaMB22KxhEOHzQpAORQ9GrGuKpSru6n0prSOF
cMJwmoXu48//84vcd0uUeEYVP3kem/xRfVONqD/gw9Xa64J/Y7ltyWZYn7O8qY/7y8pSM5wWVQsb
LesILRcOxfM4maOH53VNcjuUwbwtGhxkCNY6BZb0kw/NV07BWPpidc3pGyoqvf7f/lBPPeI8WgTC
T3T4dNDtcAO322OJ+ztl4uiaKJ2x2Ok+jZs1ACrT43FMkM3dhVzhzi6O0gHimiROMuGHNWo/83hy
OmnsnZ8sNFmEysyLzKgKuMm6GyBgsNosr3zKGl5ZIEUFhXNzNtxnZ4aw0rBozxFnub9MyV/3XkfG
WODv2BxvOyaoBUmBAbfoG/spb0lfi4GYXq7lib8t8khIrh4ZI2nsS5yWyOH1rL5jCg9dWFKpNsMo
sLq7WOWiU7IwA2vDzWs6Vwga9yr8ScPByc5wIJJ0HTxmzFrX5ctD/umd8YUHmLlfUucVYjI9iRp/
UE7MaY8KiheKAwzAI6wmUwByjSjN4ZNgQvKWfrF9ZXlX3GY6RIGOkoGkBcY0V56NyhPwXqdckcUl
1p4XjlPyCuKBQcws9Zm1wFtsooaobDUwwAs77v40et9o62v+iGj+Erukf7fqjA2onBbE65fg3y9d
MPxjbIoZrMignsn1MxsxGrjKwYe2zWs5oet6bDpVH8un7/1jVcQdUhTR7+p9m6cZTvc5Zwuf/MAh
nb7QQbaZEKFEcV4xTc3oD1jbanj+4U4RQV+dAo2bNfxUe+qj/Rup0M5+qQ7Kve5GA8gdd7GTzenL
9UMzswGBwyFgFyNfQZsdxEW73LQKK0IlycXFfbUMAsifXONsvf0Mh+t1Kp9sCR7TkA/T1v9BuBq2
MjHfl2jwZdj69jKsg259I4hzojnjU35Gj0GqChVBvcv2MfygfRY0IWIy4FRg2NuCc+B2jdRsVc8D
6DDsUpo/RMI3Zf4lc/E77+pytG8sV9qY2XfwyQofSy6xVNBqv1wWhMqrxYRmr55e3+eBVDOV/tF4
89GrM8l6SM/mU0uEeyPFm+cXhrmKEjDsH1jrf2C2ZafFZO1XOIZyqMzhuvVi+n4FCSRqaq0oSgW/
qIeKjUYoLHTJdPjHexAjXKpTnMCaWX9hwyWs0HnyLgZ8NNMomMdweBtHBoaIG6QTczgNFDm6P9ip
AjNJuaRs9Ka964wfzEOfe1UA+tE2cUBW93jyf7tvZGZNSFNDzl/6EPYMLFL9cmAefH53KRigXaAH
vY1lnEYLTnWQ1hgvGnZZXWfnidAuPBVtK09LWXaXpWFAkyZom0YCUK2VLmWpeF/FHJbiFB6FDi0+
9KEzZkzXZbaIaWy56XeNqhQvz3ab3bbdM7hDtyUv98BN0oDdOxmA6NfrI7AQl29uLqi1vPtdDnUU
rTV3ITbXjpya/uhvKpcB34NEGGCwa2v58edgeOoT45t4xJ4YEhBElohFs2qGrDG5gBpSguyQ47tg
/F8esfP5wFDwMYMt2xgv11Hd4iubNzjS1RHBtxgp0FK4b6vlTpDZ8KZrLrt9jfWclghhHzA2Wqji
If8LNU1nx0vtsDpQMu66uthftMje8ZluCIgyiLksYTKKv+hPYvw7vs4EJ1NJjCl7VVvOjjwts/e6
madUv4TYvqcGUFOb8AoKpAS+BRi/P5gcZYzmI3qFcevTjOHs4ux4v5hwyHtTiLeRBQU93Jzv3Dan
RHVCSFB9+VOo3UUGVaepYdv/RBkQcDN7NlGGM+Bhi9vKx+HAIj3YYHdjzIp/ELyoS+Bb9Mz78Wzk
7XvRRSCRJ9TdNDYhz7UzpZ4gIwl4YTfYgGB4DC6YQVbaosc5SK7h1D7gF1OO5W6GmXRqzX59vkKa
8sqCepzibuKySQ5qwWBqpg8ePOxBwSxj+h+0nhdmLCdPXk/VqlrhC3KrlZZPSXlg/dQwkOlIqByR
pXUCWbvDx3GyyyFpcpYCpQq1eKejmm+rR38TMv3pNtu75l+1+qdTutmw0jWwpwGq5vuBTKl5gSoG
rHHNNizNRJlkWE6/dVWS9kRfq5Ig+E/4cksDKTi0ncpHCQtckhbwsYeJdckG1D5reK4at9WkJa4+
AKTXPW9xtw8h5+JxBbY+D6lPs10XDgjybFNJ8Q/eYN774OwjLijy7ycLIhLT+57cbPIFVnJb4Djo
1OLp3NHZNjPlXoV2qC6qsNxk0aWgtXHJCglpFDkgzQL96eF+0dCIia1YBhvjVZCsK2NNTiIiF37g
4B0Rq4969mwGWqQg/Dpw95tVkJXZNAhCEskCctTX4KgyInK8Fqcqhl9QbaMz06nALswIVfmvRin2
5pI4dNjSbk5eaUOehxAfERTb5rHIjsqjau0Qzsw7/3BfR5wvC41OotS+FuozVMqXnLh4hHXowZTX
gDPQ/K9JYK7VsXNfXlDbdaDU5xKZdVdk8RIjL7mnqrQiGabpJN4E1dLS5MXIDbXlTfxn9h371acQ
Pepy3Q2Pv7u5y00MFP5XNh1FNh4oviKf0yMikNEQe0gOVb3FTAolOzFuzsh0Us1MP6DLuBwvajpB
CiMcFaKGzlfQ0s2txdvF5MgfSajsg87H+360tQR6YAfOyK2HoZ7zWb3Aw2cIS8/Up6rT+92c1cN9
LMX7gEWX+ljbvNhTdkzVWb2UjCOSWuBkKz5/xDgQ6xi7TEIHR+Sc9p8Dllf1nmDiWodx3aALWmBT
i3x+8QgEI6X/IN/IE3Pa45hkwJcEZcZmk4+ZFbCmhfKGVrPGmHsnIRMBuXzC2l9ubpiKHNEULAHe
dVwyXjE3NrtjIjW2f/6HVQSJ7Cm3m5bhPYqNhJlL4zagCtlp0MDI7MFcTNBJgaXrGAeP5aXsuZm0
Z0d6LhdPwQZ3FoD2xydjLYbgVHwgWlYS5BnNHzNpkVcxnDnhiaiQXcRMQK+BC1uQJkg/7koRW5l/
lKsu
`protect end_protected

