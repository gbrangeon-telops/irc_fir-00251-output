

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iisr0ydwFOm3eepmhOYSaxO3flYpViRsLN97vKyw+ai+x1TubmaH8qRRwK/QFeVsjlGTFdxookcr
olQwv0bmdw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dJvTzz+PoD3n2Ot9SgKfpEhIshJxklhDhS1tYcrcmprfs5wN+lN+5Y+o9jEEql61IqDkJEIGu0xp
zaDWEeMqwkFuovmZnp/AnbrHb7R/19zPRtwSyZ8+VQRLsRMgscwutXu29fTUST6Ribitutae85tQ
1okc5mYK0mcSMIggcMg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZijKIWnBSOuwn6R4ZrzJp1qaSPGZMrP8GTp+SV+Sn9xEivGxLJtGM40xMLXxiYuxIopDD/A1usG6
HkSoNT6OzxHJWKkUEyyVzrZuJdNHJ5q3s3y5LSNY7eMxN9lY4/gygh7aVIBAO9YWzsWu3HLtrHA5
2vsUFQxQdkG5OTLVP1rH68P4j/dhqr/LVHw+9H76c/knGyalpHLRC7tnHQcfuezFJWlkzaNGHfUo
b5cE1YTvtdlZVmw2sVG/GbXIRi5fq3+Okdy+JgckZ4dVWbI20rfa9LkI09/kwD3anyrnovVQVx9h
F0AxolVKVVyWNAaSu1fvXllqzrdJiRLbdnsq0Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LUajPw/jRTLlmEKb+9YylQ2jxw4jlSx/1GGaY1wFfWFdMwK2p0xvQMjui8K3EqJF0fnb3QNWuQDl
1vTtf04vcOAHkfRCeW7Mbp8qeUTtAsflGIPJDxHfVU8ZKprwANsENc8LVrpJ0WnjDFQIzJw7LDqc
Jj2TofWjKprdxXsMnu4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KG6kiSPrd66zvVpG96eKD+783ebVLVFNF7pXgq+rCyBBRoa0N9Hp3DIWK5125mkICodI82zuSq6k
C8aCiPbDiv4tiuIn19WDNNPL4ncknL0KLZTLAkq0BIQIsnFNRaZegM9aXOdMYGKYLpnjSD9KRWRt
WPXPZfwprSu2D7PeDZMiij3MY+cixttgVmNfcx9Kkmvg+1B5sTSDTVs3fqpJBBO1YslTmxyJAIC6
uDuGqvQ1138z6f4f+f8vMXratK1Ypo3jPPb4FTNLYJio5Vd1Nbpl9kRRtj801Ie0GGhbggK6IXJx
785o6wX6g3tRyoHXGJ4DGUmWlIHATg0KIAflYw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13424)
`protect data_block
H6Z6HaXMrKtvZSWZaPrlEBdt9kbeBX4CxVTJYg96CMfEPufj9bJu2tElY9M2iRe4dE3AG0YS8vza
PtrBWKKF09yn1RcE27enXMOJDQXd/57WMVvCzyI2vK6BL+nUlIU3rzT9blT1eO4adecNDEWmOqdk
/2zyarNlfcGixfMRBYB5bNt6doDLrR8wZgEv3mraTCd/WO7OdgkPvjGtx38TXE4BlhQTQ5KLAnBP
j0Ll8Qb7C4vw0WLjPup0k+xYcPdu1dMOZvhuQzyiJriQG0YnH/00fammnxkO9izzkDL+/jY+GceA
N0RzgN45Fal8F/uN1AVUPvGfpxnewmcz+LjBPdWJdTkAlETVfC+71/ZS8Pj3NirTTpQ5ST3kKacO
w2B1ksCJ5aEM5OsvS1qsr8+Tt6FD052FJ75RpOxG5NOovfXiybI5QvfCbGnynUbBzbzA1FW09xWI
IrfjuOOPUU+D7b53z4RYUwNf3zMDVdDX/xpCQoqgPnaYfgPs3N7w6dDxYuEq4kbcOLsm2o/sQP//
WKodfK4l7hickjq3zsSF8wDNsqNfITKcbHLO6171VUgLt0Dw23PCJ01GnqROjz+GZeFLvB6m4KEt
h++veeCMYZ8qprmY0UOJWVgu73L3CBH0nqjNtwxLHc57ERSkphJCKCMqj8RyPLleRTE+yg6Gbo9n
S68835iyN2mVcj1xjrr3hcYVDR2CqczBqUXU3lLecvN4peDD/OjFXv7/ea3bwVlFHMqx+bSRCFri
mOl6HnPxf+0eWGvPXirJcVlaOLjt95VCs7i3GICoNzFM/8La/8TPj+a4NJiSs66clBzP81FNoWrd
P2WhFIqcxuTlJ1mTq7nsh4Js72hjqHKfp986a1mR2DqGpCuIWXibi4h0jfvwF5XvA3T7ARE5xj45
ST7VnIWfaCQ2bLqCpDDFJ5d4LDsKscEqsGfT6772dCyXC3mpmE1fvK78W4Cxwoblmwc/oQ87XiCu
LaMD28QRDp6AJxlwzHGaYbnWeJxgZF2W4fHeKYyqJKkODixc1X86VzozknbTHppDE76yvZqozKgU
bFEheJMTXZAj0Gq/i2kVinBmY8FH+aGOq0OIBsJ804QiqRt6EGiIMZs60SMRdw2y3Fy3mgdc5Yhg
QD2qnPGhBdpODKOO4NBLEuKyUnaZtysAL/led3D6MvKHCbrfGfSMNjH5Waud9CbAuBGN19ue8q9l
Jw2JcsDhuTzKZpoYvswYRg7GB6hXeSACy+53P9PFLGtbr21P5ST5bXQwC57TY8/T8I63R/9NPIWO
R4wWEr21QVjLjhYj/2kRehn+iKOiQ/tkZH524Fz2OaqVNHQvDvF63iavA+iPXY7+GIDdl7AzA+Pu
k7XOqlk2G/DbJzgjffuHujI3cMsxR14jzDSFwpXHRBYafP7WBCZtqpB57X4l1j1wmwZ1g+iG/XIc
IYVNJwitA005cZOaXcge9TiWggOIskGf8ukdPG2RmVeq3WqV0YwQ8tK/RMusD+ng5U5wXATO32e2
Zz9LZmV50XeHVDz67QGEFIrvDUsKQzcwheI+DTw0K/f6kSiHHPeYAcMEZ8Pkr57wUQTgApekCORr
jq2G5/5yZbgD9w0uv2gj75LCakSos+nGiTOZiy8Fsmmq0Crstf+YJE/LyXocU+qD85CYcTXBGlGi
Bi5G6+RVpp7UqCLVDdSkcbIRAZRBVLCCPZsCBDJ7Z7N4UqWKZX4Zh51fNj5eYjF1NtMECIrby6a9
5rHpB5LYe1bkO5haIrEY23XYaDz3/5bcenVWTt9P6H64IL4ogLOQSADLyKmt1PiJI3pPk+fcah+S
2zjLRxPkjiuuS6GZjRQBG2k+sgGf6Evn3NzU+rjS6JCpCPubnPxqFVoNu3aYH2wBzhFi94GvlRFk
F7BPHp7L4rrzF/IGCewRWKmZWTiaYmMhzIGf+A4hWKJmzU+b58Q73c+jbj9iDBIkKYRBEUOUb/oX
9nmuKntHO+ub5Uctti7iT7jNptPmygkMBdupQf2OXWBuXrLy/CqV9kDUUrm4BDZRHFChUx1HYKmJ
yXQ1oZYzINGJVA+j8a+SUs4Uj54xgPtnxLlgEbJxrrCfTVCO4xyLeA+uPV5IHuPhFLyicvPOLAUW
yRmcPPlPjHlY+7Qv+Dvwu5VxqIoF09bXo0p/eb9MUvH/w2ymZDSFVCh1+HRwHIJZT1+aNUP2m+IK
rbP1AF+TgNAvtgkBpXoadLe1WIjjFKv3u3GA45TY7ZWeXnXcbGzNN/IUhTH1SqozKgz4y0qYlc46
CEnOT1OVHoAoP+Ih0udkRitRj2RBBb4DhJqHwGQIB+P1+B43FW/Y8IzlSssoSRMunGBXovxp7hbe
5kGWfzlcAyogCFVcYOwi50WxlgrmGVeK/5ejHf67D6Nt0MQEOhG7GgiKjuo0kfNmEUibsAyDPFXz
QAaFovbIEZfADMfBnGCIQE2Zv4Oh84LkLvRJSY7241+8RzstJUjtmJlkUEMQ1DPb2kJ8VKl8PBgZ
EBYvnE/4Jtz+E5AURY+6JMS3f1dx5aeTBnG6NOOOnGGKoDHhy4T+fCajOniMgTsJeBc/4Q1ld4UV
ZyMY5tiLIASEAFVWACog6HDWgOgP9VdkWDdqCETnb0Sm1chQl3kSQXcH89TC5ZYraRhQTW4MJGaV
0jz64ynXMu3J9rQ02ZCHOu4rqBUNqjfGuvFqX7oSYu4JXBvzEY4PV58hzxWqvD0p/+suAT9MWHNG
RVeyXrzA7emQukF8S5bmcGVGwBuISKR21sV9yxT9T0JHhDHTYpJTsyOW/dpsVkt2ffbSSTU4xB0J
VonH6ya57qczE17rZaZ+TVY0InQDE6/U2Tv8nMdPhdJ2J6+vEdlTjHJt8FLpFDB5oKCFvHHo0uae
w5UPFP9hz6tXk3cd7pesCWMUj0uwrRikvguSM8IWMj/nvsoNxTyJA17PgcO26txgE1/AXR0/gzwk
0c+1zkov3nNeJVq2JdBf2rHNfLGYmii/cQmaHlbv58Z9+l01mx9U74DrGajdDqG/ajXYFBrUbud7
cAMRrCFabyuJQV/EVj+UBlLpKAI0jF/YnhAWxABXBsSGKcAilp+AYEovAn/7Vr7BnObMOlU/GnnP
g6KfFG2AB8qtD2Xn8p0sUrtr02oifJvbmSwpV7lDXtttCwDJ0wfQ1g5nX4JzYJE3TLeJaCVyimDf
MgE3stZq1/QcKjeBUUwVwt+IQ6B6qIjSGEmR6eYGEpXysvAIGQgJ+//xOIPkdYjlQ3ODB8afjpqF
u8R1/LoIdoAQBSJ9XhkDCDjYncT1BHmzMyApYG5l30m9mPVpFsyvq9kj0PZ1pAcKHCXhnna3NY/5
4L85pEa+tbbRoMTUsTw9RlrI/VzGhveCV8VznekLsW6RuoAlRXt9bKSfUgH5bskTFOigbza8x6sl
fCVtGdQtzHc+a7CRPpr7sR4Dwaz6ZmYuiPYsl0SSvsd8jDLeXEzf7q9bKTyvy05oqNVfYBbQ8fwX
NLj9MgFjUrSKwW4Z7a3EMKsreuNSg+BgFb0Z9bYadf6g/DrwpbLquQ1Ijgzy/GQtAw0AVybDj/CI
LVeRnzMeaZDsO4WFmNH1Uq5/hr27rZc4gtW89psg8kj/6YZZUYq1hOGvoYjyRcbf4URkwyIJVxkb
j/v0Q4nqU4LmQxX69N241ZfchR1UQXzAwsG13cSSQtcJE3uoy6ZF4ee0TNxfH1zJqU4e6v8leo4e
GAtTOSdQeaDA1QDO4XtAHNyyIwMOX4MX1I3mk9IPI4IOKgFdWaRlzMoCU8ONrMWTMmtDSbiMDyPV
7uEiatcROVeMVyhZgBpNlcK7PpD7+rXIz4pN2z3yr1PPzVzM/T1zisZKRHKAQe+ONa7r+ErcPHPO
b3SrdCfT9T+fHGQfGUr8XMyfB1492Di18AOc9J9Dhs9MH1cmJ3Zd7+ZX3VDNjeHwzv52rd9Rj3rQ
JbYvYCKS5gwxVadVtUQZysX1G53PNNeahYwWIAnHlCXc/ZhOnHwdLbeHi8XJvcjpYB5byv9/mQ+m
l+i9egpddpsd5ZBwhdA7EXp11FrQ9JLmexA5EjfmXFkJg02t13aacHkzQNna4ma1wZX4pdW4JLaP
N75doBhwqsDBP1mrOF/IVuG+dzRk8kLNMw+W+zXFgoYeDFexVJH1fpQNUhaUjK7yk9J76fHoZyyx
nYTD2Gu2BCDGg/9l17cWEcn8kVyLyqC6rI51NyQfL3WAatiTnF5pNTHJ91shBVNMTHFwc+Rt6w0T
C2mlAwI3PVaDnZpDzODMV+Ai434JTs++E384Cf777BjFoPrnh4XOwpcUQaS7h/jLB9GWhqJG+iNj
pxkVZuAgtu4dOlcB1BF/q84F6segxFVXfuQ8jTMHl05MTsZz0fV+SRyNLJs2j206+gmHyIYQUUYh
PP10WbSPInG4VbGS77Yki70VYYnblqL4RbdTNq3DDVMNsKFhpRk0M3PmfL3CUnHiCwAPUp+7iiJF
y3Qwlz8rvcEE1843Y4fAESet2NLBXb5rkXpcMDwcTcw0Vww4PpaqTTIv/BtAqYD9pcQPr1ApptQp
ZAmb4qWEBo62fPQv0rPjf7f0KMj302WoDz3vY8q09cNd4t50e/5YjmYR8nyC7XH/yTrstlehLOSN
QVQx0nHFwtWw/7hN0nMieYAsNBH/FuRdtxX1oQWmvYipBTD6TZpb2cc0W3PNAg4FtAn9eSaJ4h7P
Cjzi/VJVzX+rqnB5IGC6qe5b+U0GN7/qWpQrCqHlpnfztSES+Oaa8doN5YPRSC8em+Y6znNMOZdj
1B+B5rF1mn9JwfFfwO5iWI9FXA7wFBkgTUR/vWbo3hc6WF+kx/JCB7MBzR5dpu+4yGqMVJN9liIh
5zxd1MKPmFqHrSDbdB6IXcAUCoyPRDTTFxp8CZhr59QwCEoZwV5gc97B+M9tcGJGPvCEUXSQZMY6
KLcZyQiiEdQptjKFXqfYvTrzlSKxi02EvvrlP82HPyi1plnyaEvzuzDGhc3h7LYS7I8+huKULvob
mHfR8821c0qE7HK5LEynA9tL7LfpdPZu6cQVCUBSdNKvh1CgqPBig2CX+5wZh0guwPAyXBhBqGoP
PMGufqPy0SJ2cdkzc6VqU+Ao9QafetEMF/f2/eB72T/lOR36qjFHUMdzqjMFxH7ugbDat+8AZSFL
Mv/3GTgBjDr+vUJ3Z4BX0lBizbt4U/eNvjT+TXRfcH91UJWKZKDu2DXMeTNFW+fZAs/IOvwVShGl
yX+OV/7kQklsVKcqpml2n5vc/S4N/Cl89rj+0N5M2EwreEFHrGBo8FmloJB4+aGwNjR+UqmNwuWo
xn4kzpiTSy202E/nTA8W1qGdZ0WJxCIEdBgjNCii/8Naasqkz6eVNZjBBplp2NHiwT3/SSWYDRK7
7eM25zf7q9LDzu+/MUexfJgzpYoHV6sQauRpeMZ8X1vwsnBbRr6FEhLpIFufa4kQOnCAkk86505s
hZ9VxLJf0O7j8ZJyC1wDJh3bQHCsYVF4wmf2gd+O2DLJFdd/4KKtGUx9FopH3yiRuWqPMzRUxo0D
XXXJiffuZb//cKBf2m1BfOYFm0Tss+/uCi50GRejiWwAwSWzDRel8lTBsFYB94cMCAVV8vrNkBf7
BfuGMODNVuaTJ7rKsrcAozYj8s5TRwyk4qGkbM38hXLZwJyHrrF8EMwVAOjHHYhlC9lfLDrD9DIl
Mb+ryNXGZomKYIrZAZS54Kq6p8HjXM8ApBGok6Y02gJirgpGCn/8idezNTSy6/QbsNcUqxz5Nd4H
wjpiMcbDTg8K+kjI2MMrm8L42F6lt/oH/7xexcyYOPxNe+5vSoay6/jWnvLVv1ozwaeNtWouxxZQ
ee1o/2KM/Bh0ldn4yAoKYw9KBt17wUsyui67py2kAuRX3aBxXswDN/TUa5BgOsvp0C7QTJKh3V+8
sJ57cnNgAEA9xNMgQfoJYIKhT6jgjU1CB5r8Q8jIo28oO8o5JIJsxAWoN/tVlsqwiYkw/p9erRYQ
9fQv8H6JabotJ0C0IwpbcwQNVGX1uqcjqyID2dLCNxsXQRZpzvLTO3QSuiIORXdF/RMe7XlkI4Jr
n8n6bO/Bj1EU86HLOC13adxZmLd9CBKcCunO50IOKB725I7sLkNAW7j+NtXp7egY3sj0G5wWtCbz
dUkh45lrDMoA23UM5CfRiifKkTtmeBIegrIIDEOuu/Z4sqOu3Ns40JIqHjxd9XyKHCDfUg31uilk
kRUU0iHZUos49wJsj33KPh1vBJu+PpFhQwux13tncYGnY2sFCZQ7QX5AG95qqOIg2UE0bCBFtVyP
sM6BXEJTRWXvaRh+hWczLibt/Mn73clSoKBmhSuqWDYw2SdtRAbbNPd5FhDuWsQAYl66g6LJg+YL
UXIRfeRI7BxHjEcjzsnH5/5GY/b5/X1wae/tPIUDc0Nayn2TUWZC9PwOwyzxKL2aebR1wgTLr19s
gM03ZJJ118/dNSLPcn9E65M48wmnlkv7vpj7qihdAXB3dqefkZ4RIPRJYyWqhwjRp665TF7v5tqv
ZLxgyDFcSApoAdOG2USfzZn3IL8ngVtyfZyxtEX5IXnwDIc5zRkMzyS+Szgx9LvUJc6bgTMPsP2/
rO+c5p2pOA9O/dBZis+AEc7U0vDwX0bxTme2AAmN/b2lniTfbPStqnVur3ieWeLN0amxif7BTR3G
gdcjnEGg5kwowRtf996SKXQNBhp6E/RiwftHZvsnXhnt5ERe0GRfRKHLjBOOCIBLaBvmiuy3TRi1
mnOovqmkkI526M1LVETi95r8XpZIAKxc0Vs/dfySiKzMSupcGHm7eX/h/pjTeV4jG/rrLV+LVVC/
GuOvNUtZR1hnARjNQ5/BG0V8jLUz9jqRtecCHY/pKCyBmmH7ppS4EW4m5REYVlhJF+NCM0jJhlFU
BI/IHFH5b8G7dhIJxknWX4d+x1UDP5QwMr5Osz/YrBzHbUDa5n9jhNzvsdM0sKXfkf9piD+QvchH
3uDD1ZUXxd75RaFyWvO7+/iMAp5PKi8nSwKYscvbrxNzUdIVtMSYw7tmGx6B9DGpaSQvD+ec9rX2
ZgxEyT4KOJxTJthht2BfGMYVwp9b8t8ZdV3nsWQ+8ROf4lMCeKoSrwMp2rRhgbeFR/wowAJFHnMV
j7M1i8Ld7c3/8Ws0n7zY4JC+SRSmY1p6EBQv1azGZ6Sje2D098lfKGE5vlCrL1tU4Smt+9xG+gf6
eQc0eoAUWN6OyuG3xku7imwNMk/GIPYBJWWNQiL5jCT4ZkFsPQwIvbxVFS1QDhjlWWcCpbx2FKcK
ULaFStJ8zYmE1J1OiI77BuTFOj2CRI4oX9qLZCkkoSbn9ixSDkckvOSxt7Gdihrxxofj9z5FuZFP
Iap+ilppCmmbkGTEVvVxDqpcSdaXm0ZPL7pXo3MAgZ+oOvVyenmmG2mL7UmmCx3S7pp/nm+aVlYx
cWpg90/9du8QDlsP+E/r+pbCtCpBWqZYsgSSUU7SLQEcZqsQ6MUO2HsfKOkEj5X2E8+n30uZV+O4
4lrjEmLmiOD3+qoN+SASY/RR+osfXalgEr7GeMK5QN5Hf1rysG/iDfk54its3P6CXbfBlniQa3rZ
p7qGxqvB+ezZenYDirLd9AnzYxkcr8qCC9b/h+pb9/pOXgV+rZwgpbTP55rmuCPP8z7KTWbHnZP5
nlj7H7rG2XYyG8B6cX39NNdixjvHqd966BkOQEW1ZfytSg6O5bpTJRuJTt/fWqZHsxZxlKTy7M81
bUn/eEYNmRQ6cW+WXH2qeEfIv2rJpjgW4TasAh3dsvcwb7hDtBtN+HuWWaAJXxXpJTSfw8npB6wY
CtmOaPhs3G+j7C91IzkLCq56GOyECkVf8si7KAchCE0f54aWE06ZHgRbL+sxMHBKgfPSR+C7CadW
5hfxjaUOICfaWtiIhiL6wLvO8HOiAfBq3GqDzTTqrSckKmR30b8IN+MN8vKT8PYv1QvzHrjQyAzk
jddfEBYRjX3cmt6c1lzW0/EJkcr7nOvY5OgyL+UeA3GcVbEcVmrs5AAcHo5J4mQFkIgDGJTUV75c
/n8CqZm29mmYK2N+BlOOrjVrBk3HWBl1KKLyAkxwQ/ecYpl81qIhD98IPG7I8X9NvMDwhPdhr3T6
lSaa6eRjTIgw+3tGdfOnK7S2j723O3O6PyeSl+hMzJREuy7G+yvQXBzhti2vpTTkXyqj33Z72A5b
3Abomnv8UoBUOMWHUq93GGvG0vvUo4EI5zsx7b7xlDDvrHINo67V6vU+CXIr3rjVpOyTji5xHxo8
Sxqr9cCiWcVI0MZqp/PUWG/9oewIDibanUpizl5Xg7JR1zGm28FMfLBaHRwwMTG7FAwAG4SXI7WQ
5S2qt6+Khs7UIl0Idu3/zB9LXT+xDE2rdJ9IX+daGNDeWWWFepFtPIDPQo9iNaiQfaYGAnUr4xpt
Fp9VipljCAdCjAlL8AlYqe6dPWf7mEjD/lpAzVXhWOE5YveXoxkgsrge1ol0XLChptKfhq/xWSlr
Xk1/AjMw/OsxvpAufX1E7QX847+Hb0Dk4zEv/9jTXWSE9WgvM+4h9NRA0AHqB29JqmeXifldvKtC
BpvDmBVq6wJCTvvXxxUTFFKq8PsvodD0U+qfmbOir9piviq515/wOWnwzqniTX3NGmKIQokFKAN+
eh9a98XEVLDhyhB6hfNQTwbT3R5zebbjCl3FtPB29wtJ4A1X3c3JQqCWsQ9XdwFMaMa/53pRV/ju
NsxtbkFan44G49JUwGtuQsv5DC7IZfbE5t5YF8/8pB2SmJ2cxgqgtt7hoHNpity7HdavrJKrjNNd
oOAxMMc0det/tKEKSkKFJ7T/5MHdxANO0i5vowJ0wy0ncQSceOEuYO4NDBCdhePdJpSyPyP7OnIj
jM+YcS11tlB9WQdRiQF9mFkOtgJPAXh3M4MQgKiZ5K7OVrk+3npBMiqV8IlgMXWmidpi/ww78e49
aguv9hC50ioJckzsKgj5BTo9jd6rSN6+S2cV1n+RtSZ/SQX/yxKxGcbHU0ndfl6/7EjBEvU4rHXF
v8Rtjp2EQ7Dk+dQKS/oslm7nPeKEpwm9dfj4x5TwA+ZXWwuuNd9rkcxTsE0VrR8/XRJN8eTo/lXP
2PPPvzVnCAfGQj/d+/xitQHCW0DLj20stFihqUxbD5hGzdmLvwVZ/TnC64C4/UOiah+kWawVBuU6
WwnoqzWdWbLLwo/wL1PZ+XpJ3c3FWnTZ2jjZeSJedZhJ0rYx1ZzbyThlM008qINGyBn5JqRqAIFr
WYpP2ZoN/BTtUn0WUStEISamHdOvClYamV1s0wcd13TBUKQkmNqsqTdfXojgTzHEDbRd36wPJhRv
ndwwLDWF3AvRXJ4wkEpNTTA0V8CrmDpjp+bmdirdjFEOkbvq8FomnnGtVuSYO2+Ti4m2YzvNdl9R
JOn7w8FJRHLQSln9MgHvWn6f/woKgFoe1fxowHV4LPiXnKhE+JHP3+CDe0gR8TwJUTWF1xRwMXAF
SJHcmTWPw7DZhHfNcm09cZssG5D6wmPcnOZqL4WiIq8LJA+v7tI5VHu9iupuQ5HcXvf0O/5vnFTH
GD97ISX8FaoHfhYuYsS/DorSoLlLLVcxv4jYfn6NlC46m1YY2p95L9XdN8G/KEFLoEFCd3A+46Ky
NapJXx683vmHpfLUtM8HDq3v0LwM81bpG7SfeqCd3BmRJ4wAAkU9KLRYVesumeVv0s1uwqIu6faJ
eace626CpCrsBUsF8M8xS5c7oZxCE/aQwoVhKcIEGKI7ZAQUv8nxDzlMkPJZe6BBZkdZeaPJFVpt
y/EGc13dM10/o928Y+TmJKNvHDMP4wlIbhDwaLIdINn05iDEkkRgMcunHlsUwQOaMcDOJqU7yOes
EIXmRNy/p8eCQ1UvTiQPjff+Bbn/+bN5oVlwGWIxASNb4nVYxlX7hO4mpEUPrP0TB6g4CGm7Gf33
dsxBgcDc5jTKloeh7f49XF0BGU5UIckb9Eii2EQwt1gZfyf88ydEPMrAQG4a1xAB+1tbKYwV+e3S
gZK+nLgsnl8qK6jrl9T4INhqWI4a3HFe0zfZX2hiIHCg5/Q5vhvd/4uB26ewi4LQEQIaxCaiX/81
PYt8pTc+mND4fq3D263MQst/xRC12fO0DaBGNSwo9qlTXmT5YdNy5DYaQFd7L54kK8egeQG+BJXU
B8bqOx5MYPSiBoAuFXeYFrvewTHi99yygwbwRSpPIIqLtbHsASbbFCxDfvuJPdbQZ8GtU8RpmhVU
zRTUhIIuPVAkVHBoGZWnGE7PrJC2MW0v7N4GE87/Vl3iDNvy5OlAmtYq/uihvT62yUpQl8yNw/z6
FN31ZYmLH8U9RX+RLJP7hP3MuMRKQegju/4K2WCFPxK65pb7hl5Ihnh9lfg4YDwsno5g5B8LO2pm
oRBKkOHMYpnU0SbbJUHAYsfEmNrVJUSc1ukboZXSzC8KL/gjvGXP2BOCySUKHEojzNCa18kqLFyt
8guYVl9dKEi7daNyRdBuA+7ng2mC8xoL85xbJV+J1Xo5psMuk1dJzxxLtzqfCV/n5QJEfyWgdVeO
XFY6WSP2Qzulild7tMVUhc8+ZmAWwagMBDESMnSiSJ6QKDMgcGjhGBP1E4xiHmj7K3quooXSR6Me
/3xBXrDOjzYb1Cdaux6Uy+aqYTuUX78n2dGOJBM22yWtLvaH6o1c425E3e3UX+p4E+d9S7ccDqPV
dYwsxc8+eJo0NRocKXhHFKv6Fvb8ss43/f9UnZ3k8mfLtm3YDIS/TTc2zyadM5vbJB+da/5breIH
Zf1VOB5CGVxHxOd7KnTbmtfEpVAApnTeUxR9LdaeaA5zVTfonDT9B4XDhkbnFk2p1eoIcvweHpCp
dkfufBpY/DYDyTIcmIpkzRxbQ2jlGOLl9cO7shBuC8lVYB4QhLBNxThCdfuBGcco6rQbU2Dc08MP
pb8auYJC1USfv34Pyx+Yj2Wrt9pn5bCbulzLhIKW0dxj+Un9OcTjgcfE4Grqs87XMhq/mA2fvM2/
ReJ4ukdSmfA+0BqZASNQT6LVC8DGUrhGIyzrTn3PcCXDmnggwkCFpApxLKDeSs395QFlXIWo5AnT
MCnL+GtrGgwK2JgPCfjv3fwWn0y3mmGB9a8aQuiP9VG3YDiM5YGRBZnObFMTwqlE/96VT8YeoxYn
jq9nfFZahKbb2sLf4O8Ibbb2Gw/aNH3+fbn1ZIFYwWondgOR5Xecw0kJ3ht+6/54i16dB+cmMekZ
P4KQopsjfQwMmydygRGSswBpo/wBePJNHkgBzBY6V/q1V3Mq82NPA0HCwDh/5dPWdaPuWf6bl0kY
3MywjNf8uXKQZbTVPZH5RCpCSEj+1aRZzrqZpB9VTa00Rxm/ORmZga5RGLhWO9x0xESte8SwqwaB
9bwBmiKE2J3lZw0H/jJGHeePHhCVhZV62550Vo/9HVwxPBW4+yewltpOu4Q43Bm1Co1/mvpTxC3V
DSTsN/EN7ZhMYffTHqoPWZ5x3MYOHvE3YMjUN+uj1AymHPQs/r5cQc2+vMNm55kSD8UIvLgbMAT1
0jRJzQfVAp5T387Ykj8gtQ6whc0fYirHZpppNqCsYGWgy/FjrVN5ayDb7y/wM71yPJA8T65v7SBw
nhdzBqTj1+RfNA97ieGd1/3B+oZWiHwFaTEnKaZikeqFG0qePYMjESlVS+LBA9aulYBfVXflM5yX
RKlGzG0LLqleTmlH/uqW4Dh2DwA9n8LkAzbC7PQnxMFAqLW62I0ACWDBobUaOgpQ9bFhrjE22mSK
69ZHua41tEQZPCvZIsK+U5gR2fkiwtFdFwiji9160TVcHjkzZWsCuFNufLdINit5/YcA+lZyByAk
o/kPns8E1706fVxFB56h1c4l+SI7+/xT7Dw7XYBRs703OnJKIty1BsG9c9bTD38q0zzZ3bJXue5B
+vkSBCyvOTpGgfR3PGdUFpqWfPEC2L6e1STHeVf8UpYewK+f4cM5kYV1ld1ZkysuC9tbGwFNIQpI
Y0+qL48Stero9mxIO3Zk6+Xz88pYMzH8dt3D9u1u6PkYa4ioBFYJen/8uIq2rURRRNdhcrfTuerw
zfxEyei6jETZZoUDcKW2jyuR5E2SWf4HQ1flglR7qPB3w02yTN7tz8FyEHqC/0O6PqsZDqzYKNZK
LpQyu5j955CnrjXWk9d0oLwIw11ArJrTmZpTNeDwhnysJgE0GkzUAHAuKACUg2wwvQPLvd/m3F0V
/DRz3lM6r79J96RpfF0Wi/V+u+wK8o14AQZz7MssU2hF3sxEgM2/yyeZaXGd21mnggIql/8FbmNo
ViFrDddfImxhphjxnUNIRyx/DTycMTIGuUjV1PKgEJJVzXp5y6JXI+HbpyPfzjGjC24DM2Esu+Xv
2LU+KYsPVbSOcd4S8tDu4lpCgaUtPvUd9CCUuZv/hD1EWAafBp/KrQPoQ1o7A9K2Vv1WdpKP8fP/
Z1B8MbQsbbpawv9zbGpZPrwKcz5VBr2644fRW0BxIw0FERRa0HO5MDfGTzGr19fjnYBXMSGi2/Bk
PhnDOE6+MqgFuxRfCEqS9eCYkiy3W8w9UwhFWa58NYMxHWH14pdusz70dbO1pdhTeu0KKiVEL80D
gThCEBE95PsMKejpITmaLgapmFahWBVDolzaY0lVypnCZMU5qcANqnkY7uq4+GnvyLCScc2Wz2wO
DTFxpw7hVjpTATSVD+eZypzqI2uV/vbqVIh90sZiDhCIC+vAF1e3of+PUjvtI5Q8mp1bLzNSNDgH
45zwMiMUX+nqE5uK32yrG/vTJK/Lb2NzwWFfW+IPihLGpqdsmbHSDWrYfT/QEkEHaugP9K7SZt+9
inbZi/88v9Yt+FAstbQM0e5ZYv6fmpU4oZrzHK6kdqcnRJve5qZL/Upr2AZEKte8RJt5gZs5im+s
u5QdNlOXsi5P/J5HsXp4diRg1grLGMtp+7X744Ksg2n+zkE0ckEr7VAvOMWp1ETMI6gW7uBZbdmX
NqNX1kJyMDBMlGfTDyfMWt11gosmKSdeYgkYcp/UUV/QmJUIHxr2r856McwNRjGmQcozIRxqBcud
tu0rlxKX0bvbunSXdlkHcsuHUpwu8S8PhgZRcBVzW5zVHNILZTEs2eJTBHid+zwlDNkE6qNiz6iX
2jgL9+F63dkWMWj1op3nX+tVz638zTIucgXrHtRoOFw95mXSTy/y1jvB4JFpjX+UYhOoUT5ca8LN
LEp1pUBaUA/QseuS9mcfdYdS1qbeeSPWSDmv/NRk/RuJ4OIYQW8zKrpMzC7e8wUyObajsHZiJX57
E7RtyiSjLY++rzeSb1hzuPegHZih0T9K2RWP2WcU/oQn0+CSxHBZ4HNX3WtfNQRxZ9B62I8lqMOP
dStOPONiFkO7Np/WRVBeP98B4NnDSc5x2ewH1hKp04xqFywCFgW8uxHGVhZ264uAMNktE3n+sffB
c0Ezo9WKsx9DV4ZFX3cJCFf+RduDhiZ/FFsV+3x3dZwBxQcpyurnZgavY746AwJvbpl+dK/ktGTL
L32LGO0Nxm1xJlM3wbdQv7iPWUL077v9jRFF0ys9TdGuVGNTGb652xlZxNYzhXBLyqmuNf6NFMCC
Cwiep0YRxxR2x25Bq8s3P+N60yx7oKTRnddxdzgWZ+Trkmo1AfVrNfs082+T4IYVItEdolRM1o0C
C94FYMFUKYwXe8X3PdpOumahEN96ZMLEZVlBqSYPds6j+8yqvfF+FyjBnaq0xcXMxitm5b02kfXr
j2yGNIMdydDaGAkz9kTuIpiDYGcGoUeNnbTJ4tU2K49BMjKpNwChUIGws3c6GNkl5o7HY5IXEaqK
ybihb3CbtEuI+/ounPiGMbQ7p3sf8aT8v43dgiTehvp5YdhDAVZLuSYEsir/efu0UhYz8+Q2HJzB
bfwV6Eo8O0H8LSBXFihgZaA/ovp6rQVSyy9DFg202gcXqn0+zHZne9XrdEzVVuhZ17avQc/UFk85
kTyNZq3MWXTo8GJP9Cr7Mrrc15zQWINfMyNaz6nJjZSTga6a69K+4dZHKok2BMsxfAC7xWf7ffJi
O1RG4gdHHMqT9xGF+4YSAyNeDPJewtMGfLEPGecu3zqR+SftOzwgWz7fL8iSoejDvU8Vrk6PAAyP
MNOAJ+nHFGZ8WL/g9OUYBxWU+v6qnaSlF09msk+oZh6eki2fAMqOQyvwZmsquSk+m/F/LO0sYMor
FL5oNVpUbXIKWPOdxzaIb99et/oGZStBDmuclmOsIstwFODPTprhFbMMU/dq7Cg1G32+ulCMTnx9
7zrCMr4TLRDFNV/ZYquSf17lnYk0xH/M9SUmb8GVxky3MzBoRJnHgWe3ybkW32MovSwAsEq8bSKc
2RYp4mFSWfvqNnRQywRYGlN0w6zrdiXbCa/taTq1hXbLz7+Oes6fqBIt4++VSDJ0aHMs0+u3er1c
IFcFQcYZ4pX9MGc6+XsGbtJa6ma62LE8z3zmh8dLgWJNxjba4oMRhiKGUvS3y0eERBdt0KK7HTIi
77PlOGH7myWoC7wI9evEkLlFdQswFMav+9n2EcSpwo4LgMMXUai0lbwbEsVtYzmzdNIpNZzir5NS
RNdYZAIBD70d3ke0UCBiDU6osgSXo5STsbqcR48egWB5jKbqXEl+9QLWiN0IhMYi6A8Itltr5hf1
En7evNK2Ctb1N73rik48mFX43aze2s4kCQa8Q2u6sOdlXW5OjRVNdyrozy45cOUBaCw1MjJC/OIL
E+WzYMhItP4m5m72h25zsUzel4WDr5O9bRBMZ9LYEnGLwp9NuFba9pDEGe6dhq1h8+Guwd7Qg70s
DCudVTvJXi3fHIsZFtLk+K/RiIZqzdEEBewQRLr0MQq/39YHt9XHbYaaZ/IhEugfdIIfT0jbqRYo
d4/f0JVlIXH2TSG/bcT8LnvvGPju/lXNosIxeKtB2phFbhaIRA1Vdu+pmzcQMmm1fkwq/+XEa271
gf2/SBZoAQmouMmz3ZlHN5Fd9jJ9xxPWmOGQ0aFLuHWyRZaObrMayEanBfNH9ajSVoCYFiAzeiaF
6IYLqCV/Rgm9csTf1gLqUhi3klp7BN8D8BPtHLVvfFAs5Jd9izcafU2COwo6sMJJbxrVf4yiopKP
DcY3uGsAoaezVqmjUM5HyHgYLT+kHn8lUU2VAg4SKewFGc9yQqLLuqCyy64Z2ReHQfNThbmgshj8
4hxWgDkOArdsSiG6CGDSBvkD3YAvBsB4pbhwNFm+lNMp0/HWDG602mTFRgujWGQPC8g4sq27ZRyC
PwF195Wun26XS7T4bSXfEi4G6Lc3T0ri86WJeJJeeNuGV3TlC4w0xJ4js5h+LAD1Bb4hPcHy52rZ
3/P01xUlT6GWCYjyOgWYoqhYmobCwrGeMGjCaKcP+0+z5c6VxLI/O+zfeNKakjr7zpRwxUgeffy3
uzog/7m5WY4P5Kkae9bFkmv+bRCLJirqlnkDST2q+ObUiaGlU9yGG4nOz9LCc1E5t+Q/1/9bbtRM
8Jv1LXbIt6AUP49D69W+eYkaMl7NxJzwYPDJctgNz0w8jKzobFyWsV3n0zC9PKzuCTmOqJ7VIFgZ
WL67TRvUv1JOjbpnrharOZinCzuJ2DXA5Vrzf9dQw6dm1m9blEh3pXfQIIr8rkRVNSJhShB+fhUs
yNRk/EIv6cHtg59FpfvItYPeWERNkZ/IxRCd3RdYMfctL//EVgP7aA2wTQV2Kor92Ct2P+HJbTUN
NWQxZUrohWXvIm2vvmXB0CVAbkxT8GR5tONC6rYWvmHjbr/S9T/DejwzgFNFuzm9oqzFNRpneGDs
rYT2wpNUOrcWaXOgfVAkcATeAEbzeWOMXKDgmsWcfMTvLh2TG0d5WzTE7aRpvrbIEwiHLCvCyi3a
lv0I+Qt0wDlhvQhLwQQenKCHxqHrf/fF//GSLwffdWqqFJeF/a6XSkvi6cwbw8TzWanuG862Lap3
0RvACjklGDLLSBAw9lOXxldkENlNdVKKOtdpAG/zehXM6cbW2+UEdE7IunwIKA7XzngMV+I0WfUE
PwkzPMHPpn3yU1S09a5a7Nyn6YWKJdl9ov9NuyzWk115DUsYj+LPm+pj8T6Mim/zzPaLpJSj9mWg
5JbCj+oricV6vDiSQE6N9fzHv2hxn0UhEjefM+SWfH76v8FOgUOqKb/J1kpJzdKNGwpedTYKNyJD
vE2+Pdiwfl4L2aWa5SVoq/9Jvem3N10y1x6Kt1KFJzHjWuuCz0oOACBx/VDcCcpwC94lXp0S5Tlz
eNStU1gtucDC1wqT1bYaJW+pH6/2afm3p2Lr6vJ9ySow+wftGJF+N0MM+anKip5T3ELYCA4fIxTL
BQ2+kEDQ20CT/VFAL6rwALQn7yBG2cCxIM7crbTKp4ZAQ9Vnfz7qqLsM1HhByeIxAxvY9HXfIEut
OkzX21cDAls98P827uD7TxwmdEI51UCIZElkZ76fZWaJDcs4qlmbe6ydbgJC/xiHilgwwDdUwJQp
+ywwaO5Qh/W36wDRNDWK6eQLY7G9TrB6M+xPj/qAzFXxkH6ntGCha8jOasNY+RzsqsjF50PPYm9q
WR9BinBHngxVDks7xhn7xLsqZnPTjlaMgl6SzZSdPZvOt8UbZThwrwzsi8TgTglszAFk3x44g9Vx
YEA6pmqk5fKqIxlkOcIybInvONajWaAIeTW6WgYjsLAX6QD596hIfyRim89lWkbAEex0jGapqDpC
la3VxptfoZBpPhkZsBor4LRXUADMGmmGih1gQlnNYrQyZjeJ4MOVm2+YRsI/S6R5AW2hdi1hdnSM
SVsi/oZ3hhvZGa2iYmjOF9o7ycBcZhEfIdsIuRMOXe+4D9+M9euqfxFOHza9P6CAGkMKQ586STpx
ZeQmr6t2onN1nNtftwV1gFSJSTcBKoWKPHBjEk4gqHKA6CFpIr/xg2cdNM2zn+IMcuZ9sOnszNV+
q7wSRHaWLmqNv3rAZKMiuQNZnqkn8V1LGqE/pZil48pCpS2g7RGwBJsB03u/Wv5hks6SbaS+wFAw
dqqiXbkUNPq9VWZDRCs64PWZgNqEE2Km53b3FATlHl1Nf2uMroxiUgJpmRjzCmNJKXTrmXjghrAL
oc8qJcvkM5m3bTKPkqk0q3YFNJjUTKDcWpMa01vheCcpalPwpW3/KdqrUfCdE/PDfL5uasjQFIaf
mGC3MwAuBv8UkVXWOVI8he4a3EfUydN/Qrc8GVKfZ6Al0g4a2d6yLl0uIUiMvNbusV86YrevWxRB
N59Ubl7geEfq0hnzP//emjwQ/x6q5k0TQzB+54UVp1WYyxzmClv4j3cnd2sEPNnigEUVJaGyQ1z6
SbhRVrGmiKrqB1f6E574TYXW4pNoDRZG2Ea5iGIjwxqLExE4KnqocG3ta7DuqzDCeUxJk3/uWuuM
EAuMCnfxkGSFF5PyKWChzOPwDkrVjkFffkM2vDlIt+eRKY6aqnbaeHw5GBL3iJaP/v57EPflXGqI
FdcSFNEDwZJilFo/QsMrZzm4If3MO2FIZthRPh+RThPY/2sbjmkinvHA4X+o/DP8cZtm2xtFnCP2
uDSqVUi+eDGXmezeXgRUy95jO3Yg1Nj5MrDbrCGPxEp7XOsO6s6UhG8dtn8w46npzNfkM11J7fCY
7SsPufkvv4+Sr1YbtkBfR156CaXRJ0JVQirw2mKaAAXwC7yGWKsogSTQoiLZtjakIf8yk3W/xHM/
sf9GkAmy+zSHKOoo1plHhzFZqON6FEB+riIfAg01Sg3zHRaYHFutBDiIYEkAp4zS//0ipOAt1bkJ
zcxlpWsy0BAZJ51ikMGK2RbYUzfua1fUSV4ZI4n21/ZlUGxGMvXV7md5WZ4Jm4PSpS2VXAqgByyT
EfzXAMfzIgrpZRqVjPXIZzAUuVQIN4zB1BafEAk=
`protect end_protected

