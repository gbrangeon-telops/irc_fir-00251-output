

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SYUpj6do5sFTflpbsRmqzQKFPQDYrJyRQArefGItBrRpeTStPf4iOexrlL2KuY5Tjxr42gzfz2no
s00d/SuK7w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NR3ykkYMNFMRKu0xHAyt5DYiOktc2YTf1JOlIURJ/ThqHJccRXVvH+Sc3vg9x993epLj5za38fd9
R5dBjv9keX+G5g1u3CtBsdqXK+hNOz/uDIy23yxr7rHw0ImE57TmiDkVMvMwv3eYKhw+6jZKYes/
orVUKkqCIC9qrUn5RTg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HlVxjhtCNCKKX+WIZOv4bglrDneJvrVwpTadJxqH8bLj9DfFux8A76EOB2zOay/g3B51jEHFXs1k
cSPeVifBOPOW+4hnoJ3TimbzQC2WXDZLrgI3HV0zvi2+v+260AsNylQU2ks3dLwbxExBHvawkhdm
qLdLQIFdyzjRMD/G+fo3ZOpvx7tOdM4iBWXd2qur6t8wJth9ryhPu98XGfaQXlmJP7Tzn+0ub08s
DCWHug4G341eF+dWmcugGtWe2Ca08XjibeU1gRioez7LDJacBlMb+me+eJNl34Hg9trbjeo+4u2p
UhjBKGy0TbAWhSuuGKcCtfIFOUbYcwT6t2Yt0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DoI+R7m0zbJxCq9A8c+QbVnIsy2kNMG29/strbjpu4rQhHX3C2LKQKMwC4UXbs35yFBTN82oCtQE
LCzB557xK8srP2DUb2FdCBqlo4nmLOUDlZKHLRnMjMktj2MJoV0ExtbMFAErwe3zZqIBchZgf5Be
0C+OuuK2xw443onEGyA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jkJi3dDxF04M0w5noeJKvbYmN6cGn5suzWOH55jYT8k6r3UxrWZdHPmAWJgyGzXTFa2rcCzw1zFN
8CUT3mqhUaMicnmv3k1IZXtmQp8LLIMHIhFQWUBUexg49lQQHlMizPzJBAEcyMQJQl2JrQBPC4y3
FtPjOGWfsQSXXVoSz8O8MOKUSTmbuzqKeAR7KYOBiW1PqJBZo+vP/teWIw2p1h9/ADBVH7fQiL3s
cyUleDPcPx934u+grxqX5IGh+uK/gO42i4Ms1tDDhMblp6piYQ998xcC3XiMWw8hwmR+KGnfqU8Q
VD22eRbZMxNB+D8sxEO3PnV48eApa0h9wT+rpw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30848)
`protect data_block
91PCBW2ezbrvmHLW2I2tMwdUpGG+ar4SRFCxEgTw+CCAb+IvlIe5WaVM1R3DTqRDprDo/Ww2/0gU
StIsR3/lHnmgEMe+QSN1wtWPJcX8ZGNYuzRRG1ip8cq3EC8lTCYgnDvk1A46qnaAFfC1pSqbrRZj
TgFI/s9IKxztleAZEy9a6Kix/CArqgK4tufgNAhStGZihMgSbIKS1nILJk1emR8PyPiMogyvxzMl
dy+4l+HQ6ehzcLTtdkKCTrBJ/ZOxwazpQ+YefqrYJvleseVXwd/8grEJIivbKYAq9C/WKyPBqHbp
jbUfPUfIss5v/5ucXmPJxv8/Jy2Zj2PyeuQkeP7hmhZiPV6YlOdRGVtsz3dCGBC4VaeldEuUlPc7
chLEegK3WKfJIqXrzseFr0A6iEf3IcCMeZCSTrhwxTaJME7uc4BAkdRAukLD/bWJ6muGwupc8jj4
sa58OSF5/E4JmdoFs/DhLsYtHMjloS2bzcFuvzCakZ+mwp9jKoLeVIDdQedFPlhmryc2A2+7kx1s
cQL2LaUX5uHiH7SwdotiOdhPmOdCT51BI66qkClt4AWXHenuE8wzKUOzJg+WGgdAlehFhUuHEG16
H1tJvmvv8EATgH80zD1v1mZZFo6abkM8pMUHWaBNHsrnFUhXFmNBWB3pGXn9lnwNzECSHOc9heYy
SnjjoxUNcz0pHYLjZ2cWL6TZEqS4JTphdDG6mzAgr/yHLCSVnGB2yL8pXjXQwSZ/BB8+hz8PHquW
7ZAjrqWMiYANk3nUeMCpZfcBYGNkV3rUdgNTjUgMeS8wFGc6owI4uVPNo+iU0wkm/t0iISpg6j+D
/laSCAAqHeWwkKwLF1Ok4Sftx5w4dg+zPftnBovZFbD11uODFjFz9psnuwjJzpLgtfgFmc2a7Fei
Z80hiVUDU2/fFBXzsykKe5n1FiX7byNkTQPd1pQqkxtn6JJjZKyZj5D/NoBi7vaOiSZwnrrlcTh8
DC54W5LUb+QPk/jHnRLeRGxBn9pOmtXdmHi/C+4n9NGxgtutGcbVXojoIdtDVjQebO7I1GkME2Vb
I4gdBsueNnRX0emeG0i2mSyUNgpYmLCLDzab+2VjBs/s9ccMKz8qqPGg4NJ1k1kmSZWBgwJmMPlS
FCWqtwgpXCkUy1VftFco9rE6oFCN2FpT0Wqzzc46lsfX8g5cTSZwwUi95aTDOphX4unI1a5Ry9ZW
9kqbz5P9Ph49vVlhhqXmnOHUOrKpN2Xfg7Nv3qP3yNcRfC/2sR5H+xijlm7kB4gLzss7w2WqWXd1
LEQ22JuQb6rXjAgzsmmN9mo9c6Z9ff4sM7a+hbXnl7Yn896K7fQnWQK4T0pv7v/wEWgEx6XNcTOV
dMw2bCqkRYwO9uwurgTq76qcd8C6xVetPwOow89qeQSYXwLAhIYinqs3sGgIHJ0wOuc2EDmhBKrd
DRw/2+1KukKVQEomE5FGeBWKb3dBfibaptDLaJBMfnDd19JgFskMG/ixW27RUzyhHHbAxvOZUkJm
HsczIv6GMmAHlqZK8QP0GwGNbhmQ26DvjcABXA9COMiCHIeA8jiZSBKSJdOvlmh4SDt8icBRonmC
egjiG4XtNEayNI15o5m/PmeqslFQ6CILigyM+wZb9opeWx/lX9iYEpKlTsZjR0CDcE4nPkhqV0Rt
O8V0VwtFCh/QuQvjSpufSFo3K1n5nYDnw2KOksX6xssV7UmxoNk4XNH7MBEoRMitY3Hn2P8ccPLv
McO8eF0mBHJhlMAEbketVEOwREAooYJz/ZeOG1l0krBxGqMesp8k5LlV6yA/CTcsJStn6EOHl5ka
8K2nWeFcRW6LIadbh3dkRufwVl5ha3qcFw0qOv9h0vsIEB1Kvfwf8nB7v1c+Zv9G6lnNUvhVq2jA
gzD3Y14coEpUbJeAq+KSxkAts5hy+N+KgJ8N+Q6XQIHJU7LNOdI5F9LDHjZonqxis0hIbj4wZ5RQ
P7Yv+6xr/O9rxa5VyJ1BEdbjr2nPbZuEwrucpPtRPcOQN2+S8t9BunBdq2kfHoNUMBIhuHEcsVUl
atFPOnbfXXSXSfS8EFkDzc+wuGfFTBm3DI9wRRm2lH6ZEimhKWMQEwn/SDldE9Z0+Kz2YUTWa+Bk
RH/I5TT0tv4De+3103YKqgl11+D+Ya+Lyy2TzHLCCAPYobs27EJA1cJjv69Xb95yLQVCxuX0lL2Y
v0kqqUqVASXXXcbtcoCwE0+O7h+RZderZzuVxWOioAF5oGS+BE16E2n6hhy9ZyvO3Ki5uRyJMoxy
XA+PoFjv1rm27tZmZNpFpfcgGFY6ZtiTmeT8M6Ob3HT6R8oDrA4EpGJMDqqcJf7MTfrAODFC781X
mhhzjL6zRR7t5646JDCPXOYdIxEUAinYRBZH90Fs5/ArYPiAWwNy9WfE4p1GSZ3oo/hIatjiyavr
LK2X8SWcbzCW70j5yj15G4iYlm8+b8mcE0Yh23UY7+jfXPRy475PRlgdiKlI20ePOfrTBEcXhHyw
rZgRrgzax2fe83pC8muAMXIgUObsFwETrTuwY95w6qW64XcnXqA481asKZRy/t/wEcq+C8ROh9g2
+RjbKf6JrlPJSj6FjVdygg1gRAeYjDUkKVjfX1Hc9aIVXI04Q395UJ52sHJAC/wPRFTdOcKl22lS
5jxKx92UuI84bkV+VMdz4NZ3RqSD1HWAJ32ZPOlqFTrsTpJXY8k4BJkLKxOKfUfxKObbV30WjQkI
BE29oJSsMQbGwopk+fb/5HqA8sy28B8ocGnjCSIE/XyLzQFY+sB8yoD7evBPDNCHr1RpFsGGS2ph
s6PWFemW69gsjPNR/fV8f+CHrGrQeJayD4iM5U7xI71elOFIjUBPYOK04aHtcdZi+Uz6ldP83urC
pGY9PFkScD6To/FoPowxQAHQM/KryRvjc8lrztPfm3Q5dTR0xeY1CuFRp43lDa82ONOA3wlHBmXU
nFjBxWHxZN+XstAbHofuf6NRcE7SPgM8sOuvA2meLdRhBTfbpKwf/sdT6G0IbPPwy57iI3fTNdvf
UyCe5k47LNFt3j9reyp5AKPtzbTH0ilvB2zuq+GlcRQFawh2st/jq4XAedbPJhRX5OZFQO7ybDOJ
lO+BMH5FF36dIeXQ/Ko5abyHjl+jEI9Ty9sOJrNAQE9mrLaI2fsFaoK4yg2c79rny4Fr0zwepG87
+xSQ5rEH+PpHvEYa+e/6gV6DEDumqjDKDsWF/Q60nH/tbybMXqJ4m/056rsLUuRIpTrpzt+hu3kQ
iepsJ1lanK49PGrCMhkMaA7r+eXMEFWuQ/gbf4k8pAVuNp/uZXWnRyvXQ5eBFoZYG0m9/8Ku6lO1
3mItbkVR1JUtD14v6g3omElF9Yunx7egvhDnIxXhK9AAD288aahCqB2qAyRf9BnJDQHWv4bVdO4k
gXJrdnS6rXwXOBOaHwiftjo6ly8UfUpFPFNm3jQRkOHHzC7vs9RzD1CiHltAdULpgThxjsIf7lCb
+7aAzp2rBhRov08Od+HCWAZCUdvgKtoOuEn72ZPXMfgjzlD0ntEjAqjt5MaMY27RHH2ocf5803uE
R48MkYnFgGEf6+Va2r/poL3/pjScvnMXVum5aclQ3KslWfzc21jpTftQohSrrgoJ2/QMe8zX5OOX
rciLDW2u1IzJtqJjQLWg/8u/ae8LfJBXjwv+co/p6SaEhx2DsFZcuUkr65U3GXc8rRkLmtDtdPwd
PLBNxNKqaKh5CK+zKX/xhgyaMBihc2tCCrWLdxBlXKUPRvIpkogw7VRSGUX/43IXPhscS2o9nkCU
70VddW94e3L7CjmY4ZETP1ZsQnIpF0cHMlC5g2bvuPaDH8BRpOBF+PmOemraLiZ1t57+FOyLenXW
pNYF8YxFfSWtV92CxO4RmYj40KoaMGgLpn7SYY2O/Xnm0nzfDLpxIGid/OI/+713hTculYfGkAWk
GMhksevUMcfe7438H9NO76xqUabTEiXOZdwcoPnRBTsA4BTk1oPXBjULkTkKp7Z4pscVjzdkQEC7
lQ+gs6iwZwAl4Q4AKgVhBhTZLpYxm/B5zLysvzmDC/I//9w9s5AEfepRXJlIzEUE9F9JPcWF9F/W
uFfb7W/7hEI5g054PL2YPJ3waR0GTx3tJ2e01RkFPx9lOpCybp60ldZp4Zp56Uqh3GQmlU2+qMAx
L5s8qVs858MPxxCNBaC3F5HezbTcUEVmgB9PNwEj/6MxMtA5xzSMBtb+wQXA64W5yfJ3WzZuw9WY
oPqOMZHrdZehLYcQdd61vcPA25CkCb/V8AdvfGuG5JXlId6QPcFzv9L99If8akKl7B8Eym58ee31
3s3R0qKNc6uAGl/XsOFBBzsppjZ/8dTLFtdDCax5ixGug/UUmWzrSu97Wt7IpxOGJvu2RzzdPAn0
YNRNZsncDXRPmkPFTvMN9Y0DCGk8WfhSYJBf9vlmEdckaI96UqK/DbnGZp+zLyxLAJhtR7GBYLzI
oMcbaTSqVem4mAR6Zj/Xx0u/FxKy2C0mXTYTZll2paDI98TLSe487lhaCX59NL7vwq0zhCCLHcHh
jTXBLzMyFDLrHR1WgwsLzsMq9/UXo00j6+vM2M8eKoER9wwLA1YI1gg824JV6oh6uEAUt3pMLoER
jVf1zo32AD2qpQlGUW+CX3sDY4OwDSukr2Vphq0cjMcMxZagAzphf8HKILd0xX48otA1Frdd2XSy
48PdHR4mxGLRfrwQcJB49D0EPO2+btmEgrRy8WgftFOF40yPHZCKBsPlJTeQi08HUJK/KLdKbB7J
L3SQimvuipSyphb6rSleX2Omg56b3uTp0fVp7HvZaKf1OiwuYHrwz7EMVrPgUsRkJuK7vjHs7spW
FXErleaRjwQ/KInRowZpntEsD5fORUDNOAZsJT+gxCs++OJyAZJyoRFUTAXxEgLmVtF0tFZNt3J3
TDmVby1SWXpQrEXemDvf2ZSAsPOt56V8OMRMEx287WfLGhT5uT9gQq+3chrrDqcq5RDyjvlSXRZM
/BOeCgPu7oyRagHg54pqz7Tt+JYrTg/R5OpjNDENF+tELT5q7Glw9e9in9xhbjpotpNL9VqWE7ID
2708Q90zOIIt1k+2g7kM7cAh5woHBQ7VgrQjQ1SAB0QTBYShizTuYamBFl625IqBfRJQJr90Rhd9
0nJ7XPrAIIizoVGVqbqE7QMi+bTEwo2vtuYc6jY9O/jWrl5RHd5tpttIxqUS7I2XysauLEpLo/bv
uqQIGjdzsmJHi0LFO1Yc6qgL8810hF1exJDvOgBzCC7I0WFqnkXsjUFg1Yih9R/W5G6nTXvSvzE5
dFOk+ZRyK50ZpNwzWaEFRvEaCPglMuiyrw9RPaoh6uGvROE70u+QJ03KggygXMh87job90NJ0xFA
+jn7HLzTj+DGTKppqehtgCb2Di6qPQtTjCZiYlzKv1jbBEokvJgOB+LDvT7U9jQYPQ6gGBMwdPMS
Sx53gO2L7BJUiTP1TLnC9ZDMEZNgdCxcwnajZMPP7yT6ItyRZsLTp1frrm183R3BNIPuhgNXV7F8
D5rhciMNF75iz+hsPFSR/oOV7Ybt3AeHIfy5Ai/2GNxhGI0rz3dtKdeyp7mrAuXcfSossqMqz5Yg
4w7g5iSTA/TzwsNlnnLW+7kOelNPuCxY2RJ+su1WDhBvAB0jCjJ/jT6MHMfou2RYsSn7c1/vFKB5
Kjn/FZ+CSiTRuni/lxnwVoo0To14aNBelhEaeJW4Z0i5rs4fdTqycr47TbJK59qKf9II5us/aMmi
4ahFuESXi0p2KTEKDSzLBdzt0CbG8mqiTNfgfwEhSN5KZ+ZwL4oJ/OL9BvfB9SGwCxyXmjW4Q3Gs
m3LNt1qRINRiZ8k4T4zL2kFU1H5N/yvb23kE+QlNpPkIYm7Ldt94IkidZ1dwWIS6PZvW8V4Y8/9+
ig700bxpGzXUcIz/ko5K3oOL4V3RirzNvCWxGsHOzrOwIHWllBtMfEeQeyXaCsvtXpocQbPcyOch
YcMArZUzWQVnyoYveMpgj2HCGAmtL13jGFTdNtt/ALCzrby81rtR7DQLPggvCc9ia819NQmcCU+V
qT8qEuvjNXxY8tbBkfLME68snJZ6ljgUgqORSOSd7umFqZASDqkqr6Ylm0J0IYTVyD5EPss+9rLk
Ni2Vp+jAQro1BZ9/r7uFF2i6oOOwHX4nEX7HWNe/eTh6a6T/LiyOo3sB7A+ICynSWJHgd4pyO8CL
n4BF5LMPao5Kephph38fE2mxUIiWMcPOuiABmoCtXu0Il2yTsXXuAhZ9pxaEw95MOGA2QwtYtZpA
JvhLN89ggv40Y7WVpOQlzsPf18/nJGUOmeMWziQRKPp8V7yUg+CbUkxPqnTwVdGkrANIuW3I6su0
XtbAtT1Q9FEvnAteY2RkGOUbNIJKwuu0TW4LAxLJhmjvGHcUBhRCeeQW3YYLgFd2h9fmIpB3Obrd
z/Vnu6A5Sty6NEFE+aw2FU/9snwe2lq7YMHOdPhxXekHTdOqhmlDmGOZcfVj0eqpXgPM82Ui7On8
mCPMA8A0w10ZRyyweUW248TYKBFmJFIgYP2X9e8wMVTF3F6syF8iwvQuJ01jGes2M4uF+FJxxsKB
aP4/ZW4eZt6UI2H0pRaLVe9YfzPoB8S/I90rpQ4y5DKeZYY8R7FeVNd7aHXoESQyF8Em9YNG29gz
RJO6v1Am6p4MTdidRAxX133lUBAcZTAA6zIVRrYrRragVGJewJ24rYIuOVhPJch4UZy0ypCF72+g
YKdbGPcDv0r6JjAqqDt4otbSTfJJo/dWlkppftM4NDR/Q//TvmtLahNPRSopKId6FXK8p0R1Fb/O
oX0ai5B96eWxmw0y81HTI3Itet19/3naz787BXNH123+vf00ls7HTLhJD4x0YgfN2sKx3Htkavot
CMqrhJTpyMhO9pwZkMttOY2SF+dfE/bnAmqgTlTV1nuPlsHdVf/xrr9StgFI63259jHzBkyA53kH
oC5Gq3xOV3bJbUy9MD0P6z+zBbi44Oltfux9OxG8a4IRjACH6zbMaTt6S+hoD+h7WX0JFhwp74oI
DEKw3bpM5oslgWhmeQOvQ9CwAQXpT++1geZKYHbqxvctuwucmZTgCViKVjbcTJrV45nKRfrfznTj
uGEQBAh/FYB9aYxuNu2WIVY5lW3vHFv3XF0OwHhCdKSq5n3uW+/j2ALyg+uuinIbdcUOfoNBEnXW
b1iNojYJbXZFsVCgEh4A2WDhiTKQQhwSRyG/KZCAerYBkBCqR/wiBVX+ktaBgvKFV2u7tpzlVdNk
ge1QgRVtOENMDIFIXsRM/8aJl9mQgo19KWiJlTnlcKRJX9YOpAbrOGS+R8tyHb4IQmdXGGRxn5iR
PaDAIO5tM0z7VAEy7HbehJFnbALgsRiK0yzxWgKGDRYr/XugcEHgudTooTJJ4pIRTUhcNqM5L8ru
/TpT9eyIVht9kXQ1I8bj0jED3HWGMYEhe1eoqKnIFEmkf0Cof2ZIgZ8HipS6PJ8f5u1u5nEbeYX8
ORoDup9wdkjmveEtnfcPQ0/ljuLDeC7d8fdYK2JMi1JggpPph9Mrla2U/bzsJSK/aMV+q6ATFmOv
elw/hL8GVCupB3DHrG2vLvi9ezIOLSodFn1Cbcna7CBeIpmxe/BKcIHqVCY9BwqVWpGOzYwstVw8
OBi/GJ3arDfIcWWQHtDUNvPz5Q9UGqOs2vzEs+l4eIhbZ93Wt3cO7nfu1lEFOdGZcBRRwa7v5Unt
OlKftcdW/koNFFUmuUn0ZYVivRo2uZF6xgLq8nWeKiS8Nz3PBhOOS+osrOtAfAPKcigpXF/rTz5b
JYqw87oErHoPe/p3cG/pQRpe/eix2pNx2HGR55apTOKAcx1WGvYP3PViGt3gAwGMJDk96761HB6B
PedkCLyGgmdR41xY3db688D1ITKi7Aa1ejgZ2+7Dsa/0nzzvNtVY7QJTaQjomtDPYsCzpYwFjW5A
AjWDc1HkcstE0cmBHLc9z5S9znLspl4rOpQrx3yMtRhyjp5KsYigL3Rq4ZrqsWdXr8H9taOoBv27
C0jcyk6Z/IpojvaLzPX7Cfo501kNuw3pUg+1aZeOimKSEeCIDv/i2SIjTMIaDi0fOY9AAeGvIBv6
fdhLy1sg2IAMcNmj5lJD5bTu2+LRgPTrfFSfLnEu8aEy+kYC50HGX4ArY1rxs/ENC/ZHbbax0ms0
zwuUyL4vNcdN/hQ8z/xg1Xxn6ERa6nCWdWZc0LpGBkMc3oaNCziGuHnCbql6w12CwTGC2KR+9iau
A53Oc2m3G7V1FbTKC/IP16Cy0GIze/ObcpHTu0oe8FSXFc02R7awgrfJr4si11DYtU3wyRLGriov
pbYZULMJVWgxRC3h6/25jB19LCHVeVE3DtLuzcaaurK/HaBK4y8pyqs+Zb5SXWLhW3Tz1ZO2J3xs
yfpxy7zUWVrwuOMUC/LcpdKy0a7koxXbdcEDbM0LRi4akqA7+WyCMLIzX3xEl5RsaMfINHaGPVSL
9oatIqiZvCOuWZfrjaxvUeVzzxbsBOAp4whBWo2/9vOGCuSg9oh6/2fAKL7v+/xkNyeJHs2Im0vA
ZdugYTTxdxo8yivEvaFtApUyM0xDkJ9Y3gnmtEWK9GFp5tge5ZzYnLGu+YA5llpF5f235S2PkXxw
+Cpqnw2xpUpYyqJzEqvUwTrhcENX/4yMAcPzYvpDXFQLfCj4Rjz+HSqzBn7/2cXZ7RX+ZKKoRTjp
E5D1bH3A8NGbF80YzbMFOE3RZBbEH44/IYbmon45HF20B7n7LJQGc7MGHoILDpQF/8uXj26B/j/T
peC1Bq3x9tvh12re2tJPRt3zx1znUfV5XPcNp9G75FncBfZEZWTLRPnqarbZO4+CbEVdIszcOZYC
q5FS3BNTxOlBYsd2JDFRBgr2gLSSzlmoMX8ZNd1/5iwq8ysXXyB5ygNQ1S6xzgfnxAxHa63QC6BA
focmpq1MHDtulk3Ro0rxKCo9XpM5F9/+LjWPDQz/Z1FaG7yROwbXFCbgI3xsnOfAa13jc5DfSiiD
G3TNZ6zHms307l2FRTxRZ7hMSVUMQomB08ZL91apM/mg3EDKNDUOoa4Wtc49fyZ1rPLEHOtn+XOb
aaILVZqyjehKCgRoDtzwAtSXsZjlhIana47qzsfF5jv49nXbcAP//ozwQfCIZued7k4MpIxP31E/
27qTgWTPgApBDfGkvzQWFh2JfLYbYAAwoQ/wszKvvDF5VpnbTBq+Vawec4uxhYnd3da/ikGqF5IV
qXONmvdHK9modVnYBfIZHimbhHA/ku8tL9mbIOPAF7mU/wfuyyLDhYpn7lp0Eu14FbFgDBwsjBOe
gsWJWmzUwse/AkHQpwokrkZvBVn/zfgk+4aOS3/MtkwVLkeebeaRt8/7XawE6DmlpBKXmepVdort
amwViDfBLCs8xVV/DDf6KojjRqiwvFZ0KcUGvw2VR1MeDL98HnnaQhQug08YptkcufR2/GUeu3Ju
+Q8Ztyy8cckoAdY+V2DU0U/ah7UH5zzKmlkd/gP0Rha8MXYk0y/ZCNyFunKxixGcfEl89vKHwYwq
oGNVDZ3+oYr2Tjep9nS4cVXIVOfDghs84ziLycAg3M65l6nUwAsVT76YPsH8cVA19XcqHv8AAKtY
THXcO7VYy95O5Wt0Wa+fGC9gQ4Iz4+R1LHSAUvI5nCaE/30CHJJBEUCHIGVGD6WbWzpAqyhcpFi8
IR4OT/hE4lGg5DKj9YtoGkxM24cVXpLI53/XTiAYtId+Ich/YhpNbIcHFwo2GwoQwhPy4VIKDlxT
sffcguWwrJ47sMyOxsVPnooErEhzCc4pSm/r43IzYdzEpV0+9gP9CCdoleHbTZVSuRWhf6JbJvaj
yA6Ruae77oAxrjFBU7vcPCNKuSbQScy1Ho8z9z5hYNyCFlKecixCHin0rxvNZvOfBeqlT4q9uE6F
DCrc2VfDXuy/1bEHFA+i4WPwJQ0khW+wuMEBf4FkKB6HD5qyS7oH/yjPSPfMmbwkMCL9CMA8pJlu
4Er9Qk4LSgaYmwea2NvX4EZg4WWD7y4KpGBVnmMzR3TXvu/sIpobWF8kP/dAB6Z5oPXbI3DkyjNN
apxn7RU2efT//tW7p83pBhgy90kJzRbuGnOvSvf6cZetbYD9IQa6ZkzKVj7zGR9GgbLg9UF7kt3h
7zWO3zSxEIoD4Y+vEYGjVkyqcigD1LP/bsgME66ICCw2f4G3TIofr6hYfGcTdbme+BLIPGh5RCSS
O4grEThH2rqSvTIn4W6aQ2GgwFp52FOBcdgvWEV5sFGMSaFLlGa54Hnte4zeCfPU1cwQSNSJMQ/j
vn75vFF28KfVKv4OkctMIXD/At97tzqOjWHRI9GKyHVBkP0ck7t/tU5WeajzCZNmWMJaAW/8My2k
M4f1N9ab2BlQC88skQuIsBHmuee5acti6uyOT+WWFmxSKvgvQoPJeebh8Kux7G/0cCY+I0qZWFgR
WUUkumd0UUKr++oBouxVwcIBAkD+WqK4M7AUZhRywEnZzNmeCVQo/hb990tT4funvIFyFWvCJjG0
oPg/Jywv/jDjiRMuonY9cggYSc449caxU8A8z3Vrhmk2m9lxHfeqLs3eUPXYQg9lpkYJ0iKzdrTH
Gz5lCKosKU8IPBL6h2CDDFoGUXkYXN2YmFKK+D5BakdIqWVu5Od7ofdIUyN8psywIDOk90UZGp7f
Az/OrsNuwo6iMdEBQB82yQ99XywSxe2JBGkueaomTRmdWfsMXuDGpTuLzxmrnUcbZn+hPYg+mw1f
l+19Fk04OKaE/J+HTMtOtVbRSiS5QB8jTT71tnQ7VE3jVqdsM8B+JnOSIPdFW2cFHGZ+4/ztorHR
UORwIAPxjyOgR6Ef+eFybrHbw/0znsp7yOv15R0LjKThaoRwRu6PcgEEsNsa78tWKmYgqpJTP0y4
3pPajqam717110//Q9Soj1/yGur4IrSTPwA+ibuuNoDRl3stJ6PZMgrfX1i0hBQPtcuc1Mpll2c8
LxXnQNRtfQMWBt9QjaEL5E4vNIxTQ3Pfu71EcknU0rdvDxuycRX/xVBGHkGkGioUWmv3AOAaMSQ3
i/MJ1lxDz5wo+lCeKvV0rjN2OK5CCXjrvjZjjq7dyr0LngLWeOggBUx68X09gi7lsCQjN9Vo+22X
fRya9Jg22BiizG3llJqTwhx66zzZzlzkAffLCBkzp7N73S/zeDNkCpyLyCLLwT5535Lw1kxwFi6s
3uuQZSTh9EmVM+BA5v+OIwnKvagm4YUSw4oeE6XKAz1gW2JEosDnaiFS02JJ15mMmjSdOUQ2iNBg
0gBlfF5NcWjkHQe+NKk8MmsM02MFqzVc+n+g9NwiZ6wNjH18BPVPGIJJXJUupYQnO+sc/Y51F1nS
noi4mIjUq5RDj3A64JQyODmAP5/LQyOY4iOh8rzS4PDTto16hvnO+WlhpL7Wd2ujdlP0COO0EB4F
cby44qnjKETx/o/MMDYSxPq+h+H7MIEM2NhemySR+w8EN4mX2UVz0sCcV66JYP3eYmLHg+2bGN1O
vs+sw0bni/65FfP8HrLwAqUHUOUkN8KBsJXVb4aBi+RRvedmGRjgVEBTULxa2Agc+2CpI5qFle2W
qQBNk1E9rAPeun3ma7a7h8ohPDxIJVvILPLfG8hEtPGGayrE84yZPpZXr6vsHuEQ8IqoY+opZVTW
/F5JQ/3j1pKh0N15zoMuZd/UFuBCWxjwtxkkarhzPxPgADzfp2ukg55U4Q/2y9vgolWzRh7Bf+JB
fZw9osYSCvhrc5NW0vqzmoSSNLOrg3Gc33WLY3KSJPbt7m5bsiqGaUlcvQ/Dg4KptL7x0OrkdsBQ
9ptVgHtihIRrQ98Rc6SgebU2L7tVBz6DIB2wNQvfMlMcS81Q5JZVz9fu8G/xI+7yKdGxdz0lur5v
NCByUtlp1iyLszBQexHGbrDyt4d6m79QErQZFRtoqTWQeWiuL4LuE9cwsMtLBCJTHBZrIphXSnJA
ZtgOpvGiAwochWoA1e+Zm9Jxr8iYL4pQCjuqHakxZoZlNuc7xavPa7P5R1c9V+4YHuNysCrRy2du
32Z88a/YRE5xgw+B5RS2YtmoqjxSr/XRWOML0qTE/HSP+165vtcZymD0eGRZjMkxkNQqzBE2iHOu
LNS8SZL4j9zf+jSp/CtWYZJ7iIzlR16kv1TAJaU60aws/l/UqpiviSAqUKGh4IStlO021nWuaA5U
g6qzfHDQrsompSqQfFHjcikrRmOl5YRg4fBPlUgKJZJL16XrkVidcjASyRTYO5x3QocTXKfv3Stb
NTL/ZQblfNKWjIbVkYPNJslMjWvTgkcWtE5ktdnbfA1bdLVfXiJmR9t8ddRey7tnqkX+/NiG85VQ
7eJ52ewJvabW1kcGlFBpuvqift31s5Prj++EwTvTTXRStT+yWllUeMDoTIsMOC04Dc6AmsL7VQAr
9kp2KHGQjfZ30hN/pJ962KfNXfNz0Fi+no577p3lvBiYDQdJCxVNjx6P3CLinOS5xaI3Hi4T8CDE
eteLczpw0LpOwzVCWlwzjkbvcXB0ICQAW4qQufqqJIuqPrv8t7ZNOfqHgmBuqJH7nq4YUVv+gQxl
RTQT/+o0P9WdvpK/DCb7jUzGbkZjm8yHfvIqsCOS+w8tugoexe0Seq4ouJYTIUH+MLEo2j5sHTmE
5dsIHNGDcTFOQQsknxVaEHpm68XQyRPZq+ePlxkIwAYxUDFfOE8qij09cuj8xiPzj/o36kVWyo8+
2tauoVSnRAQKnMa+HEH3URRBCPXMuJKa91326B7g/mwJ5W8yfgKiddZx0WFESEOSNaxACyIVeyYW
UByAJLfcp20cLE3d4JTuL2iYAfOLJtjDEQ5zG7djCBSga44nOrcPrvlHWG6KlJcmvuqu6RM/ym9T
DUBxb5+0fPCUuIUk5I9Sqh7bZM+N3PLAdi+gDf60ez1g62kJ6z2iVTlvxRrRLP+FXOP93YQqjgVQ
Yg2Ti9Wvb0PyrP44mLN/tC91SIz/wh8BLupQNUH01MNVKpFhsvAA8A2kGtTwLSR4+cXkhPzsjiOb
iWxoQ1DPQPFGrW5oS4PyKUyA1FeolxQisOVzDVZlGok6m8jqgqId/P2mSMj0leyWEygUuA8CEQeQ
NdkPndrvPXmrtF8P0+vkLdv8C4KxQz5+0h84/ImqphsqKz2ryGtlcByN0QzUDfjD+1m+Sle/QoPm
tkdj0P1PqaxrBC+jMTF7IlWkQMykRq44ZDVzd5UfV5G7hSnLTsctBMujRHGVfzh9JMUUW+ooDQ62
v72qPKTJg5g6Cj5EGuy4FZELMO6ngvnCkK/Z1UcCQh0BFxcfr+Y5gqbJONBwbMHS0XQv0E+vRWXy
yAh6CxjxnUh8fAqU8O/Q+lfbYWVdzjU/NpU86rkNkAqw9cAL0s88BvqaOKs/Atp9yJjyZ9Q4+aEa
oQyxIRlCnSptQbppGugYBUJeFzV3t/FoM3Q42PN1V12+SRtVliHLdHtEyRBG4gWdjTYGm3uTbSQx
hapqdtzS0MRI+EpoCe8muM300c2eyCGIBuhdY3Vah1BVhId+xMcZ/mxyKN9HT5eLNujhlrGlevdq
G+hhGvTe/s5YLI7dQG70/V6WXg7s3Rj2EGPzPfzf5Ud6z4YUe4C4Q2GYEHzRY20e9+gjrLxau7Nb
pAQ5DNPTy72NRMv8xOy/5F3XK0bKqe3RxjFep1OIZkGhZyM0+Yse6Co1sVFflpyztg+8DiwpWe2U
Ys+8V2EJuDBVN4trBIpzWOX0DsNe9KqpYsnxgZmHi8064iVmgZHhd3w6f198MfdTneEymZ6ylpVg
XLMRja/Y8RQZnQ6YgiOk/ccdmHdFWbYGKwGo6yF6dVWWjCrhIthH4MknrkUd8pOw3zbbaIP5sm3E
zTHaVzFzdCuc7tFAhnvCxOgD0cNjXzuyey01godorRKEK5ptmaMuGhKHO+RylMrolF9rhzlYx25D
1ZELdzjJBhUYoa7DWeRPdclcCMT5RVfspJt++w4uQ+SNy92mIYVgJIBUFdyy2F9XGv/M7HJMWNuG
8Kq/6hA+xHsh9sJFleb9D5LSL5CuUaJTz+jjTyezcVIm7t4rmm4LxcnC76mwoSc4Zw0tFqQKRi02
AEFgEUMNzGJP5BYEtJ/EIUi2AWxdws5caVOeWw2qKFPMu4V7qLkuleJfbKnQzvUxhZ03BgYKzrAN
RruQXQMJDk992SYv7Z1fRoKFgBcnCGU3BSkfKdy9KDlkvsQTtDUy17Po3huVhTimrlsMRBPFyHa/
moYZ1BWoY5RKFcGfT7MzqiyzmWEGwhDY88sOyE48kYh0Ip/Gws2IYzkk5Upt8RS4gbfBQWvRoTmU
PRn1oVVPmzQShwcaRxy9Y0bBqh6oq78dqyHpAFwcJiLOi7pFs0rk89+IbXFqgI+Tvq79WTk+8JC3
UKSsoQtIdeLhdtPXJU5195bs0lRWzKIe0Po7mbQBqHjAsVWDT8Fl/V/TR3axVeBtHxgNy+Uk6fxA
gAnQ/DSutd9i/WlRDnXbieYZW7q6Aqam9m5nVNnNvwpKctMnZT54lB68vLPm+RGomoip+u54uL8b
rScAQK5RcDszoZTuT3dTSyLG0OvnnT5tp3a3fk0nVh723nzk87Nv2vn3RWXK7bcQsaWpFUAxij6S
hXg9F7ifUx2Epzr8OgiIx7f+PDRbIGcSS9hjZijtPE7poewDgcdQOtCvvM3SCIA3guJV0rL36cIw
coedDviT8ZQcVQ/6M1yJWFr40ZETq7KK7yypRNaJxtLG4RI80R2MKnFlxdeCjqeJu6M5B50ybAp0
yGiVM5b2uNqr0+ttipTSnNkDDxxav8u7BKT734+1/uyvAoqNfiUA4dzuvqi43e17wRJ0v8kKe2ha
1ow30ISS78nh1P0ertEFzxRw+tgtOIYuoEpD4wf/6gzYqFwC3+6cC+DGUUEg/wTfGJHYJz4E8z65
Sn/G6jGcpuO8TRuD9B8O5wfYGvL+/3m06M5FkreADF1qzZURwcfGQq89MyXDOr8WtwcImyWxkqC1
ENKM1JqKUd3psjjHrWMrfWqy+SUxBSWyWB8UP+pGAxGNMhRnk4zFMijc5l6akjEZmXYslCRqw1Z4
sUsUZqqkq+uiMECR9tCJffLqERjrXlrcAs/Wx7WpDwwhdPZF5tqMYKKRo5AV9MAiTlhZFwKOBOCa
oWP5gSK3Rfh94reEPU0Y70Q9kzC6gHbg+C26MbAQXqEdj6symZuiAWBvIsQiaJoWgnAQPKmOWemp
+SsFVMV/HUDo0NNW5o9OhMhMpdO5SkpnSVzdvBcvM95gGXHc7vjPdxLfgQNVQ5cN7FwDk8oiiCNZ
YwilD9qgnvv1dTkeQMBH+Qzv7ghp5TRV00wA16daElw3OgeNcEfZlOvcvHYkotUqEkHA9wjdnv8Y
UXYEcKQXUPd4e108uJV9bC3aY0ps7n/bpeq6tfQZy79Zb4A1CdsS15QmW6YxfSrIdTL8+wDjzjbE
D5yJoNYQcvPYD0oH1VhEnHBJ8ZE/dx7bxUV0Gd+S5sSAxiUmq9JsN4p739rlq2CMBjrQEh7VQZKJ
E5PA4kF+sDQZRlMJpy/a3CQuLQUWYQsBIg5JsunvMOxEnEsXq9NfU0hldlDmwpsVa8DpUaieAbF0
H/3lXR6P2uNgk3mtrRU5PqJGTSHgROhG9ZXgYLqRl7QZIA/zevDyzxBcll2jPxNlZL5S1e8pwNMj
diFdYRfoAK7H9nEBX68+8G/yXAq2oovK96fx+tvua/6tZROCAYAi8sEuqYgw9vsmH+5lECgq6Sud
E37GkkPCZnf8FmevS5G7RV5lhZVEyxUfxCeaqMUDBJZjyAxXNQ9Xuq3ZrwGEt0639ur9WqbfR4Jk
q463Yyp3pOc47Mkd3L7WBfXvT2B9H3AEDMoR5mbCGtBPuG4XVQe7aQPmPVc0/eHFqm2VkNOo0eET
zBezQ5t3nvg10dtkFWZs0FcF5F6LX9NwG51tldXEKE6TmXMoY1VVAwzcSOrogNDwNbKSy/SidA4Z
hVZ0gB3GLJwJZI/kUMw4q5eEs2GoWtXjPmeGaFjdqW0gh4wtRG3KQbgqJALfd1kOvj6clz2yXTI0
OPno0iIHzPxZekQlzf2t+PCshVGLH4e96Fe//8qdUPn0p7uMO7DipJeDVI7D6TAwS/Hl0ciXB/CE
57OMl3nHjYKxIvw123bayZWfBL0MepmW4exsTijpCbdoO76va57zj1ko45ntZCwQlzyKdzhxbkZ1
es8YeMhkUbOyj/F8R0+7NzqXjVaQGHtvmNWn9UYX1uhE/KZcb/DzDNhRY2DCTThJkiZ/EYp6svU5
RANlyB4sGDFMPC7UpI2+qhnaLZ6PUovT1k3X7tku2oxzaTDnQDd9fZkr5kmQi2uFizPzF1XXrctw
fuX6NJe2D3AhT44I2/FdaFeJ+180IR4dSOZbDEwHIGZHIzzIuqkXEK0C+79vMvhsf/ztkoarmj1v
9ueaoL0Zy+7TzFwSyVG+h2/rx0SvpgVIhIfAmClYuHBEGwNQ1EGu8FdYKOoyVKKPpfmHBoGLP3VQ
D4Z4dqGvUJtyZdqL1iUa5tMvHJ+q+ikrVnJ4aq78rBNPz74fxiHOIaNnNNsVTQd9uuzSgkkhOvEb
7mJYlBD1JJ+VUcQRbZVWUpp0nVVKvn1sU+y5rBMNTVK9R+kyzPBOOMid3srIqBjqiJ169Ajrk/YV
aTzXFBl5E9l0YHKOZmyVJFtPcW6punF/T46/WbzebC8hvHRVMDAs/jyPs4ThFOxWa4i6+p67vwlL
fvG19CKW3R4nb7T2DHX8PvMTp8qkTvB6pYXYOwBnqiAzOdWV+L+Ua9ktjd8MD9dRtx8/iApH3li/
POaXV63qscgj7rH7UMmXSscaf38Vr8reNqawW57rsmT3f+073232MV5nONVLUQ764aeDyVkm+MTw
xnDqBufF/Iv31nhtMxKnva5on548nNBOGhYLQ9/zxSS2+C1PT9zcm1raSudefDGu3B38vW04cDov
6lfT0lbP5nEdfJNj7rw4FMoR+gIFTgB/pVHn99O1DN/s1f86DbgTS1aoyff/3tGDdRQGNtmp6ugx
8rbf/iGRZJJHcsEsFPdRb1OkJvixjqZH/1OZluJs5tvOauvj+cpnwH3HXaTVAYWZH8SDi0xiAHZ1
Di8QuVph+LJHk6dwG2iPiHj/T6VUQ8Cbd71t8GGHBJ/j/WO97FMUHD64d6Za7gm+fCanyWa/ryiF
R2G21026YjvcrRB6e8FR9BvgR5qtWa5nXqh3BuCHUg9VjaMaBHGjw8hkiDCieslsAZ/QZ1VPpaKq
2CvLJoZXzWuOf80frVBgLlBliNBR3/JBqszoF4ilduOSCGEYZnrap2Db8drZLfqULubYfeeHcgEK
vzb1f9MMp5sjdVhVYJFZUiv4FPpZX5BIBU8OCAeI7A+xw//8PZQTk+nRIOl89nyJrrF5WxqWFlit
i3ELuB1G5Z4GUWEdyfFmRTpvOErzQpEY66t/lknVhwalSbK35b9ikTGMdrR4WmpW2BZ6TeORvR4N
+1G3CJSAqtCp8iFUNycQSCUfpM+b8alzXTxouK3/+8AKzxJ4feQxPVyyS0RRwX4oZnIqIuv7bvW8
UfJCZKg3e8KGP12DfDzCzYsFJjQFylQr5gO9LGj5YPtr9ysTorM/5PtE+ahTYNJH3/20CrV10f1F
YKJ9MCbAgdWkiIvhjmoJTIrp2hIiMoCI77FvpNxuUFEPtM8KORd2MjRQepGOX23skcnq7nJ28JvF
6PLq7G+V5edfOi+nB6rag7+xLGYxOWuKZkihLCSOS1A4p8Mi5J/vTyVA9dNx5BKmHej39Vd7o5mv
w711YgDx1WKl5hoYF9oWCQa9enEDnhRTmN6HcJAEmwCgH1AkjNZEpzrV/OmB3Dpiad38xFeHzaNB
y4ppbmcbKE/UFbxte87PIr911d6MDLOA0CqXArHcA2Brp7xwheqmcxI89h+yKeuwi9gr5mYBbhui
Jo3HtlnWcoxD94ll+vNfA0sqq8nhy0WpKGU0IcKxXPz3KVrnfZ/WaVlmeo7G9gnMIQmodLVyFA0q
ljiRzC9pSui75vF2HZeZ3salxzTomobSjyRyO4ZTS0qS5exL19hlpQ6TKLefbX0SQqVVpO7Oj+tA
uL4jI6euJz3BwIBMj9dttXdQH/Okt2ZeZKijRG/JC1OEwV989EQruG9bo23t9AhEzOARn55oLM5w
UOeSzyKWi0hj0K8GlXbYGL8hG0ZpE7K3QtiarLlM8SjCYQ3kKzVJ24hXeqce7p1bJp1dEV7gQrEu
hC5ORtJd+wp58mWV0NZQ39vuzIcp5FhZXfx9R+rL6dOXgC03MPpKlRZ4K4MSaAfYmIL1jfFFFGLK
Zvf7SV+Vwh1UdIRENIcmT6uEF59ihF5uLkT3mIiVl1ejFlFQJ25rmOGcadla9iW6vdWsUiDmbdav
eIknKmd9AKtvtQZgINodQdjMiTAvGaBdWwfvAO0lGSVbUI+80EbehmegKigW5TQSqspvpdUnisI+
W5Nx/AGuEdOpTXqAPt1uugT9Km6HiIx9neWKe4hicEj3uw953jmBeGmEmoyLFzZ8myAHuzzk2G7U
YSwKlGEPSqWQoZ303T6WygYzEvgt3frqQFHLBDjnSHWB4B48FLezCI37nxdbC1oZTvmtshSGbBgb
4K/XCE6se0dO+IhLl9iBrBQgfZR0YLihtbJJka361L7lYHYp71wwzZ407S5p16Ebft/nn9yJq7Na
D3j2casFIMH8/L/jktafZ2u93FbFHkqUTRz6MNCCX1J6J67zG+CYmsFmp1YWgTl6gOrDaVVaX5SN
2oVU1dVhuKavycVLqcO59/73x2vXnsmBQpgqDlymqUxrorsA5BETPQeJ45mI02/I2RsA+m0pnYVl
JJU3rAVT0BfdkxWmU2g5chMxo1NN5esZcovWQ1c71KUPuFNNtjJWMcE0kkO8x1/5MA6A93AuxotG
8pMK6HJxgqWd2AtV7jc4u1/N6Tgh7cXhyQKO2SyQDGT01n92IQybgml2MJ5GQ3lHYVhBg3BVhFZi
Ytl+qlEIswY3aYGAp9EeEbXRhrhIvvtK8i48ZyGAuBMrtZoClj/EFTnb13v+nj3tc5gtmj9d1Frn
xh1tyKW3IlMpr3diaIbC1Pr1HIz0UTy9/Hyk2HSPp1fjRVO67Z2z6HV1C3gfgjxjF+T0e0MsJNJ3
GVVIkngdml+CxAAY6bB+Zt8wwj0wTSLGeuXaBaBKGDEqMJV4IeuzKG28VOg1CJeZ6SJh1r2pNO+j
7eYkqT4YM2awyedOnyK/n4pxWSiJm7u6QFUwH4krYG8zNCxBYEYkG0AoCqjAoTH3WNohzC5ZP6lz
sPtqeAE/pvJXLuQxNG7knB1ildCRV/5FvL51mewUOg0p5xMkCAxKEn5UEHAF0bovvlX6qdT4KY+f
7FajGVyMuQnS6A4RNy/aRUJF5londRVeihIurG4B6Bh4V8bvUmoi+DbSULglMUowwzn6vi+FeoA4
UQIAModythWitePsH72vx8lb2jab9y1vnuQZf12muvXxhWBQPA7LJachCKhTrdtJQC5EOz3C3h9F
L/aZXXf5Ir7XLYuw7yJKANFFW3LMbD9IHBbkGs12hMSfvgPYVvw1fabfyfGfbY/uC6CHQDyoxpF2
D4h7h+qNM479Oq52sFQsQ4hI+f/uFM2XSiQ/fPEMD1VLvb+S4gQwJBvh3ErxhRRZFP1FcsWR29jO
miiFQIdpyJnAxumt0gei2MR+V1eLlEeBo/uejv9heeVblo12mmrnk/CAifbQ06upZMwn944Dy3sV
AmBz0IjLpQ6W794t2ENEASZrTH+GfGpHbvg0C9CEfoE1m9NOLDwja1gnIuy8NmWeRjKFZzAah2TX
u0oMt2ROuEs9JM0pojLv22xiWuo7DTS4aK6EUfKruxbVP5uKGYZBj8SpB+LvDXlsSxMWDGriBXbF
SznbIk7AUCGQnMNsdjH9RHUikJvni8Vc8gZ3DcKIGYElNgx6DK+3AxBReqAnwfts/aeVaOs32Aj0
PgVBz99t9d14FJe+6RR/ktit3Ny1Ieh5V2kTMlvQwQeTycGCSAyfc3Ye3s8yqRAyGYiKmVNIh4Rl
SxUA02K5EtSrYso0Vr+hEgg/q/0UTwvA6GN5x9eUy6WsKHmMSksWOpQRV76q9ogCjsthtOYTXa8M
ZcNzfZFurZcFANvTMrl518OlAJKQQpqJRauyZx8GS+D1Z0PzDiLZDzEiqKv6nMA292BjYe4Jv0w1
+ivaXd+H9ngQyR1veg3z+ll3aSnefx2W9Gqz6XZHSSDim2Bxvw/bs4c3bKeUyZ0xN97GivXqs6UF
qKZd9y3RYEUjThuaV2lXOo9k/WslsdboXusbHGpGfmj/7XVXYFG4jEr8/ExzhBnj6uubRkFWQrix
PptADkA6h6DRRpPRweReQDT/x7dyoVhbQ9d52/0KV+KNv2btzSG9wyfjPm9TVclPJsZiLHJvceD2
2eetW7eChptkhOQltYpyHc11Rk3nt+dhQvc6E8SFxv5sTm2hCgQLXWM3s+mM/ziugXBwwPEpBeM5
wCAZV/ys7+RZqMMK81TbAonFquM7Hx99HCi6KZVuSSje/cbaFBcAbNs+yhhClrO5jX6M26adRf1x
5H3E26a9rpRj4i63/u1dB6/FnzusrMmTgyIPeOryHW7Ep/gi2+HxU1mMVh8IL0HiDCti9iHqj23j
a81O3IMMxeIzyOSEnlFnu14Vq5TQjlmXpQ3o4vQ9h63mREuP6qE54ModOa92Xlv47A8RWGs4ry9G
lX7OAfGB1jBbo0oz3xADvuzo1743WPquRCX3pi09/vLKxO+BrNO0sBaGHaY/1+LnHGuZJWoK62I/
0nT1bYsDZqE4mJwCCVjAV6syqRjwV9bpTzMRG1m18pUQvoqy4cfA+nDOBUNBLNKONsIrme8l5t2t
QU54XxxE3FaJU19Onr+hpmij9gdBIED1snawyy5XMvpKR9rJXk7jXhixJNqVoKe8AcB89KGd2l6z
QT78UOcmT3cn2FMR35qYyfF6HqnFVIl+gnUkBsJFc+Aj8cZSIU3hCxC301xkXcId1CcmliV29H0I
iH8Gk/F+YGLh/3X7LrQUYTiIu3/2EtVMqzR3w1ZDrgYmNeH2nkGfRC+7daXyh8nWkD6S75nX+4CU
m416501SKVYcoXCaYwQ6YXpnHxGxGxjdHBOsuXemdIsAOYKRjj4V2H+wtg/dEr2p6kv+lpadUGJo
/94a6Ht5a5IfqYO605NMLQqOgZND2PApnu6SsCSCFthUT1+c6r4FoWsCsRwo6JX0UJVrd9VUUJ7p
g271ux8rPh4PyazGFlEBfMuL/3nHMEPyUPHzYtOUjHQh/kB+sUhiu7czACaJS87RJreedhroufsQ
JAdxNNUP/6blBaWiB2WNhYvrBwkYD0by1E0FdOjEqBkxSOJ+KhOX7eWW52tGE6A6yYvI8Knj43R7
toLg1WfApqQxGoctR3e7820Y8+nNSrb7OzvAAVnufbPpe0KSXiOfPsgALQ6idXoHjFvkZJ7Ik+/E
0FTRq9JxHizGCi/EZWcuQhTVqrPm2NqHhet+ZuGx8lBejE/vlvnAmlMWdt+TqKR1S3x4DGjwivt8
GUR3JCTA4Yc8pLcoCv434X2GWnxVdNqdrPFHqdpGlRM8OJWgDt/5Ine9s0P3PEYuBx7c2s1LKBgy
i2Xwlr1TnT1uRQa1WOxRpUN5IUMDCCR2wDKeO/2gaUN+yoKGAbKoJ693YcYOrEsXpgoe34v9pjSO
dl83+MxxyJb2dwar27eLKzuMW9VcoGbUnUJm4WEwV25kii3hdveh7i87UQTcrljswP6aXC9LsjSD
toUMQRpAGORmmWTXGpwPhax6HEm9OKEgx42OZ+7383J0c6Y2+v9Z+j6Q/5FfiUHGBLf3jqC1Ez4N
iMMGE0/UUm5qpBLEQMynhZWW0mO8DQaxGFX3kQlKht8hvOw4Ys+wfY60Acx4SKMObVcSFzfCXN4j
idZu6gfV+atYguObMjXG3MoEpvXkHM/3n31sZUJzmv6UwuoTYy0DbyJx5/l66veEYg/Fr3dTz1E+
2sTyb4zRXCkAQQ11dbiJ9vScc2YCugQ6vIXDg8ngsSTc7qQ6e8cEWTg7XB+IAIvH9IHxcQXo2R/x
kj+wR9+Qgd5s9zfmOvzeoaddHEJ0TE1GQkUjByinCC1o3nal2R/RIEuQK1sTzgBT9Uox6DOpcLn+
RLvOlvLMf5iV9MkTrIPNCTk/mPxwKN+VioriGOE2QSkRQhT3U700Moyu4X7pVJCE3HXRrDhPCu/L
yS9bmyV2qgN8haikJF32x/D3NUM075JZMU5BPs9W9gmOENbXP2bO9/TuM4EQzgYpm696PK5M7uJz
ou6oGryYy6cGtg/rqvyvqPiwXB0svT+lg5GESxwPuTw/msoNlByPZd15jDeh8GqvkGwOFb/ODgWP
xfkgPL5ER1FR/NgapwMk6lb+QlM+SI2W2lU1sYWJKwoU+WYYnaws0UXsGAp7vepUegAGjFqbMakV
9I8jNrFlphD6iJU3lsv/FU/I5TTvLvilq7E27CjGVgZ3XuxB6QNA2jGl0x2DJ0z9nUsr4F9Jg85B
k3SFMlJTWBY6YEjpnXDfdDfIsTe6vh7tLbd/VWs5EL+3ZoX15Wk5w3+Ptj4pNl4z+dQiqNOdUV8M
nzwb8XxgyXuZ0nk5mjiykT+TcH/xUMuSUTg03wkhYHGpOKNuG/+JbpMMHIG3kTrShrANHpi93aM1
r2O86YW0l5quKZq7IDFsZq/+SqMsLBzjb11rc+WjdSVA/mmuvvap/11VSKvCSCb/Sw/nJWbPmXOV
bE0COVaMzhvWuqbNQW9+6Zc6CFtex+9PssNOoepzhBU1nD0oRwvDBVhgPw/NqJnqplxYaCp9fWyG
FMKga0UJkR/cTUVgpkYOQ6LeyzSVjd1HJ73VIIVKmJ/Eh7VyrVpBlQSdQHEn4kpTxkBu1d7duLkj
lfTISO91LLLcBrE8h44CDpmpEKLJjn4Nd6uMnvFSlP4IRMwIiYMV027xyqmclKLDWLEKMHUm0Ub0
RahAUdWUr2Q3O6J1zRvQcmmiO3//bggQvdCUNZZt0upPP1qrWQuMRk/KXB2TXInEvGPWwP7jNPfa
dqBS5LN4aUCEXzOXMMgYWgY4xoPX8Wyp7mNSLLc8qSsiaazOBPK/AAUnd3dmOhpLs9JjyT1pKMJx
uXK4ulaHQuGFiVOxSENwyChXfbvQoE645J75Aq5IfExwW29iG9oFbfQbUOmmxXxXKOfvQB3ZuwpY
qvydCwxj5rPsppmmY/xIHM736hqe6v+JE2PA1DD+SwQHtYIqCYp8kq5iXBS7+S0VePfV6gCD1TCb
zzdbj/LU/lCpL5u5/vf/rxlfTP9M0bJoIMlwxEXlFgkO6AFa/xY75zq0MIEe8oK6ZSZ99LOt+z9y
yTqrf0ZJBuKrRkubT6CEtFQ1h7JjOhTPm6kNqGGpeS6Zsffx+6uIEMF2K8PzZE9tY0iQQFqU6/jq
Fsby9hjzGwX3OeJKMeBGHHFpjcK/tvhQzY/NZR6CFI35C0Qhd1sN27GI9y2JjQKtD8/xPl0LQqWs
RsKaaaTZDxhm6N6jNE/RjmEhjvMwRCHVilGPFzo2aa7iytfFqbhBcK1tKTmdHkxFSUy56LjwYP3X
NcaWhP/TZlJaglYPLA7YHifCjgnfIVgC7lKNMh+5DeG8uPVVy1RtH43iRGj/+J4mdtoeRR0a8j45
tTFKaRGzTd81a1VXi6rZAMimre6jJZ1cRulyN4RIyZMFckkEqOfikxHsy2qGVdaZ6fU+VrPioTlZ
KCsQIMY9I8V+CHYWQe9u5Z222SEo98PVRgzxJHiLrteW4cPrJjE3P8CJCRvcAt0qDoWeFsxUE6ps
xg3QQB/C7Wcut4alhWzknHfkxPTtuK+UHqrpj7ZJtm50oQeSqixhAVN2kglFOrtOaMN7W01S8gRh
OfHHqwBHCAh+5QsplymZ5R3AuCcI5y/AIR1IV21YIgM+1ticXzMkJObyQMoQ+h4HrnR0MWlic5WY
kHDrkLrCzGWkv4cGFnZsK2IOAJPMSUX32N/tLJZSqpYhYW1KnZ4+HpPv/ixgiRZwBnhn/NMzkWO3
MBK4iJA9v+dg1IqH93OeqDaVV/US/6szv76fDsIJHUZYKmVvqGEgANiBxmVlcPK3drTsAqj3ERP0
/TJGw5uuPoFOISqvdgldSj0p21eYWJ198P78SvcnI8+nshRUeenDh47RIVLJiqs5H1SytTPbx/F1
c9NoJJRAbqhlPkdP/VGIh7oU78FAqW6cZhs8Tlk99cxGpHCFoGcFY5Ws2eBTxHgphHtqSS/1NAoo
esvWhtJyH0EPbsDDqqmzna+7A7wwkVrb81i86zFEk3IIdRG4hbtE0a9T4rUM7DNNXVB3Y9kFNsnu
J0keZ6IT08VPGmGWNGztKDkSOF2hgl+6qZgtHtGRK39Pgsda69SYTxaowAnjUB9BH+JuZ/Kj6wx4
85XFOP7ha/ZxxUx09JS+QOXwpynbumnJhxzJs5QZsCy3RP1LyvFHNHhu5U90ILFl+t3TE9Rt67eE
OpAZjn8JxuiJvgG4GD6uElk6d9lQJL/aEvdI591N4Y/r0JRbrfrIc7m+uKD/y5UhieOa7TsWzyeY
gCZ4Y2DERab58MGs4tmdA98Dk+kzrQIUQ4FuxrGtNQd+H7esFhMe/rpUo8s918phB5JA2s30JITB
m48yphgMUx4558Vh0G2WbWXKxHUHpa/+EvicLUzs331VvR8toGiq0T7mj8nTjJ0FsWAjOSv5ZSex
kfv6BKzPbj6N106VB6WQySsMrYLKpNCUtQtqUlNk73D2z2WC1HCtw0Cyn2Wm7mpNiudGwjNAblWe
todD86SZ4Rv8w5ePh1iX7IlIjNPMnI+dFMVbv6Q45Tn7+vW6Wi8ekJ1XzTaASLPTYGpV8Gy8w+9Z
ppqmIWJ4RZxmB0d+Koa1tvHjtutrK7rAkApUahu8zBqfJAnjWWuZ4cLjJlfll73UTo7GD6yOZgOT
V9jfZ7m+pfyuJIQlgfYHZ70cukyvqjjdNY0RXh9OA4kTwoQEbC+r0FMoTVs6BAdff13/vBbAxrDx
myoBF6wZ3xJsZPS4e7pHsOdqU7hH8b3DnF0xphR/q0m3GFteIQQJq4oH6g/18mhAcHzinRbcZuwx
/A27VLhA0gs+Nfx9DFeRbhXOUUnCjhUQ2+Mqv5eiQ3pTLQkfvDT0aa13PRCNHvIm5i97uQIJcyRf
rAsXHMu0IQtIMbwcxsp/00DxxN/PDaSDoDOHMtfGuV0/0+tiWAKwYDK303u4ic229aEAHhki7MW6
JzDif5AF9y8GH3IK1OZ2AN+ECdMuLrzl1k3lXJp0NHKV0NSbpOWgtG6tjJ+BLkhZuztCbCGyHl7n
C3YzXGhMTn902aJ2OgCr1A3pYfXjD1/j8NITH4q9F71ZIWHWhmxEonw10JrZG9y97YcgQeWulgkH
FyDYNCDU+xOHHz+4+vzo94MGb5clMLDKHS+niRH/5yYjV7Ok1FwNsEBt7pE1NgE9JowdKQ1JZj9k
tQb5gJfzL1duMxoMQcTlTD5mHtceq7mM7bqe3LtdWVvysIJjK83Camt2UJokWJLMCos0KI+4ELYN
6h7XwaCuzjFZ+VXe7tfV/SDE07syVjVIT7BQUQvKUnR9AdgLHF3FKYcJX3BjJkZeKym8dWAGCyRZ
srzu2f8+TjoBbr7QjIbFgJ446brDB2ylf6Wut7e/rE0CS8MX06P35v8sKZoca2IeheAX/kCTRsDG
B0u9tawFMpmdIHW5JJNJOG5Ghfz0NHAkGOHfUgAppEQmbsCB5nBYBwGhp4OQjtYxRXrPRsR7JLvA
lRqpgFwPYWnidGfVSLVvpSdydTdYq6UUFEEWLExk/HOAFiEQhnByuVzDlJkQToZvTCPEAnG/IKLW
jh92FGpGQtU6Q/h0gjCOzOXNARbVZnqy5jPY5lMEBnpPUMS56AbrHz5V9pnxqbIW1P32Ex68G2XL
HgqAncfGS8qh7KqAZjorU5rwlGe5V1vg3//KYDx5Hc/gxqFZoSKVIdyoGDy558xPSBSVC7yPANCa
pVyeR5LumCEASdMDyPl3x6V7O1Papu7TjhfcBlQFOdoN475htH9XL8z1jvMImHAZL+rLBmrd2jC1
OWiaLNcR2qSuAhj3rIVaOAOZyX5r8eCy4pvmSdBOComD+1eZrtFi8+yuVZjWPZWlVK//L2/wBgQv
7+TZrzoSiMREsBnynQ6FWozBUwFznRtHMFAoVnfAk68G12D9iCe6gZuou95pp+7qVOhY1db4TDVK
NyK7u2Mnp2zrUyDIrICJwUw+9L/qO/8WrAT+aRtW/1rkeC/rVlfUCtBDDc5klbLExP3SgfkKB+zl
To2asnZGWZfvw+QW/nO5IDoXwick+uP88JB1JsNj2S3DboJ7racVtO5eW9Yt0uhvQ78C5nBGk8qW
GqzpDd9jYQzc3UjrnXYZjYjrmquuuaTM067JBKY2KQQYA2VHmovGYw65i00ywfMIFbeOJNp9EM0i
ZYQcMliwqExuf5pzWpJUw8ZFifl9SpDIDJ5GGXqYNE4OXvj6iAZVKaw8IAzlS08VcTQFricZzS3t
UbJrIm8bq7l+XNPH21H3g5x8GbCwgOaVMHa/ZMjzG8vMPX8+TdUeZ/SpWmy0+IBPnCmRb1ccprE4
zBGPVGRZ86MyNpEr/VuIyFtgEnM/k5OVI9679TD2lqciMxRO53/sekSIpsCUG5LKZFPb+gnW/7Ja
tqSn/PdTVd5K3Ch6uvqgzROxkN+1luFfnKbsqJwrA3/Rg3LpRDDXFK1W38WX3OJ/Zq+BStco6bZq
TzRvR0sLio8XR3qOBn84EuH1xDfDRnHl/CgRGpXOEpBUrrLWVabJoWnzNZJWNow6LX5l5BQbQKbh
lxECFMRWOCcq7PWMO2Ea/LKewvBuxFTMdvbGqQI1umfflN8/3G2MViu8esQsI3DTI9S2cIRElzfy
uAF39g/SC9jSV1BCMl76Kv6ouHB5Er9bdeXJpX0wtdjcpWw5Ho+VG3x92nQyNQTHW1fphpw9ziC4
fK/oG9GI0JOgmugfeNlaNRMrAm4rJlPQgXfJCVV2E3wVW0azlotkqmvkKERH9QMSSgdJtVPcW4j4
iNSNV9MYpbfhXxYeEOKjdwGsdJjLtbvP9wRhXXrYJUccfSTiaS6SfFPthq+frXMbqEzzNgHWwOUl
WuQUdQ3zpLGY1meBDd8G+oLpf/heykFUjzXXZTIGjtQT2VSROfCXDRgCjo8c524HVl13r2ThAbRO
IdTSf6ohmHAMrzDxLCY8wckWePw64kFBIbVW2jvEdQYGalEXrfB0jkU+WzICTBwaRQDfQEiM4ttc
byGxN3jJr/43Eoj1/4ndwApSEDR0rfZ/U3XoDpyQARXKz8Pvzjt0Mc/yl1neQNVFSAXuzdzucDVx
nU5+lt5BrytSh7KbZv0PpSa+GEYoPyUXYqOVz3O1XavWU9MjWGE3fgA6YKOjMFOKgRgbPP/JcmbH
W91Ug/cTDtsHOp/6kQ/wGgi5uTLPHFVFBiWAIGgJs1TIurO6hScayFLfXCJjfLV5/jQjAt7UGwCo
5QlepdIfyQW9EwmBaE+vxtBeVaW6omIc6zO09IqBrniJaA3FWeLdZPGG9pRMkV16j6VROOFs6+JS
Ddq8YT+1vUNFxYLn6mEZKJ5ta+Fp6EM0iYxN/a1w7fw5cXHaxJr8RJG70lVLBsBurejcJCEHD/D1
4aBT/JEoKLZnrkN/hlfsiBURSF+NP4NRn5X0yK6HeQvJ1CY04BIwQxMvE10J95yLGWlN7diSugwY
g43dNHjz89rgL6TvrqKaZhIQT2NwJarjvVesDbxsJYTmNFeSZj8tih8SO1VFDU3EKO1fWs53eP/z
E9z8y923qL+hpXmw0ADoE44sG76Y0iwDPiqY06Nfh0Yzp6tvfq3AKy0EiSg7Ks9v96go0KhAAXH0
GkpZTTZRK8qB09KjlmXS1alrs00CAWyNbIo89r8ZmkHmLcEnTvqhvHpKrPaJj2x8DeE0lQbaXeyH
ZFM98yGbYKCWAElYTeGzycs4bIPqA/Cvy2nREcGn8oKN85bzfBsw5xcWp2Jnm+bn3XtpgXKIiQgw
n7LB4UyZrVhx2WtlPO6cHZc4ueHH47QrwxUKBmReH1cq1SvJkxgHWmfcshshatGEpZrEAp+wB/Mk
YJ2OxoIddylqH0qcCBkqrbYJ8n3LlGB2iXfDSZZZVRv5cNJU+rsT/pL78ZLCtPgtpBDxtG8bujcr
ylriZsB9WtLR/6tCxEF/OX/wK9+A9Afby7gs99Oa2oAHe+eN5dSmaHkvJxtF9rwFLfeRyICANfTS
kz6zKPLtaikjQUjGx07r1+rnqI7WJ1wSmmDz7lg6Pi0ywf8sYTGD1kbhNzvCtGqyGj7v9SVSmNjW
2DatwX4EzB+a8EZJu7KsXAXHdhGU0/iO+vhqXP3scHKI1dOZllyj9uzs05xNU9JebI7FI3T54C5Y
PAgdip8xbt9LMiwuMp22HezE7IEf73ADskgCFtysI+5oJtN0fM9Sp8RyHyh6gO+vjalY0XdEUPyL
CsTWaWgQ5SHG6wactcpGoiD2UR9MUem3YN0PdLTGZ51fd09J3oWd1pxDPLrQU0ltHnsgoEFE74tg
CNjtBaEkJNVDkyn7TCxFND8rNhyE+tsPni5uORyNjXD70JJDhJk1Ccquamnt79/mXdFmhs2+T7S2
iJAinxGUF2hjehrdXKoOyYbCmXeh5a+gs+LFRZn3SYRVNSv6rBGSSEbNLhVboiNUqxrnm/6Vlke/
jiNJA4L7E2dVE+VD3vvaCiue2FKWOZb1QYHv//3Ti7A8SbDIFKs+BdilL3+gfayVdYQA8PW4SCz/
hRMhURHtRQUXlv5seG7V/uC1Q9HA294zQKHmYPRNYOv7zyLj4xpH9loXizQzfKcZYCzngug8S9Uc
uJjqGS1z0P/lPQ9wwBFh1W6W1KmvONYAG6KPlg4J3kNBwZPM9yU+A7+Xt4IHM5ezd5HYxdUTgLz9
ebGc1plKMYy8qibJhK1Jpt7imicpR+bZ6stal27r9XGdqc3zGH1AfCHHthyXNXyqp9fUnagObXpg
XoMrZ286OSLeHhotDUIA0op5zUAzUts75iTOTZkIW7wku3FMCLJH19Q1kRigPrL/k7D4aI45hb3R
J3WDBdZN6vPVL0yjoYScf5nuf45SOPiofAWnliML3A4BzDUucFJO3TAl61OabWsdAQOw43DlU5fW
tL4K0Le4LWTQ8Oz8uGua6tLz+zaCHBxhuP+tcxuGehhLBz4gAdhO/NUrRRpSGz8vRNS8w1RA47c6
k6YqmNB1UqGg3z/YIN7GrJ5SJ9oe3dNK+c3xGWAfCOT2ZtmYDb8CcydYq+BjjzxI/Fpukr2TAZCR
tfh3S6QQyqNUct3+vrfuXVaqlHnhSHc0AV4Q03KNWqDc3RsYlomxTiafjxKt7esD7yMfkJDv4kdl
NygSdXb396UxRzJW9f+zyA5kxZVxg5ZfXnxtAXo3+7bFX7U8zMY1KXMy1fmnhsY/Q5ebphezGAnV
yJJc/Ybu+39AeYtBVeGRjjEwjpvWE3D7XughTezO5rUVMR4YYlG/ymdp642E9QiafDJ68DDC2k1R
SAW5bqyR1XWyU9t0ga82HAjemfJPn6CPX6e4RbsLHZE8ITIfS/c080030sVbNTaTaFm5pYqVaG4s
yD9TFj1xZglG38gAlSDRR2Vw5kgCHEEcXNTMaTf3Nglc2Tc0sm1z5JpVu7jBAucqAqpgm6FReKcK
WsNlt6/Vvp5/TghLUlNCQPV0I0wHUAbBbjZig/hNipQ+wmaZR3cl3bE/BYA4M3rYZpOKGqh43Snt
qDUi7Boz3yLI4nXynkO9DY89GidgKWX6FhULuB9hcAEn0zGvbjayddA/qrKBJ2qo8VrGQKtKgNak
m1yiOzN5VIk4gNkbuILwQt1IlSlMffUidKb/R5xX5Xi5CXK88ab/2q6xsdVFaOPT9Ui5NMKHX/rg
5hdC6kBSyIA+p0owek7/BvqMFfA/3LaviEhlNW+HXWPX9dyZfqJq44w9GrHE/6sB//68arZHd0kZ
uB8gWOslAJju0z2N834jR6/Sup/A/dSYhK9fpAPwLspxRt/shzAeEjYq1QEBJr9et+N0ATBDtW4n
Lc020OMb6U9eekXhmJiJMNJ/X+UMI48I43U3TomweHBLnC4PY1JyZNswRfp1i1YbJG4cnmXnWLQt
/2pHnbh7cLCPhAen9Uf6mSolH8COcp6ESncZQa5PgxkztJU+QNN3n5OI8Bg2MnEiuuLYqpAwyUIC
kOlaPFm8qXkTYD9mR0oIyFQwj/KbohudLG8Jd2skasVO3qSznNF3Sk+XM8BAIjWX6oLbsqjbppba
z11IINTia0R1A6BnQ8UbM+WXYhPaTHJSBuEvI/sgVVWKvq7+gEK3trwLAnd2rzK7ktjOoqcKPWkd
tvBo++ipPs/1iGU0LEIUNbt6JAWf+EgzAjyZ6yP/S0n39urByKs2TF1MoKO63bSNVqx8qm+J/5Va
OOGhTwoNnT5lta0dQNrpOVahvyKXwcNNOl60NC1oPtr1M01cZtvbo3dbqRwvunb7WpGZ1sq7THi3
aTOc8CRBG0hr5BwqiSsU4BTAU/sbvFUWxhf5A3Pp+703QX2uUBPM3xoRSzkAIOQFa6jnGN/JlrSd
makqrCC2YHlyH1GyJesSwfMRL/sPBT/Hp/l7mON599aBV+gEBhn2q9ve5rZ9FaXQZUVonBcqDsm7
6sWpKy9wXWgw7CrJgvIQb7TSGebCuM0DIWWOICgxPVoVF7YT/M7w3LbR2pW5etnNE8+6uQTMyPlt
qsB4XmI4FT/4cuOlTf5CYJgBkyOJlJ1WlfhUOgP/QHLIeFXqkEJE5ZhE4X0chPDQED6sok9v1tW9
Kac+P5QVq+1UttbyqxkDSFoPR6TOwdAwV/HjyjDYlwJSw5TARTbJ2V5Gs1OS6e41kjWRCLeSu6BI
55ZZvL1hWYJSnITp8PCTAi2i/xJQbvsoLgoR1KSZ9T4IBFAFi+hTtJ/yf904tNDcppyN5uQf6Qif
qZL9fFBnMkynAACebwo/IDIvOQw5WEBo2i19VKMW7rqRJcnTgygZubDwhR4HGSXelO9g43QzjXts
7srHJAD1Ps43z+JQCcwwdvtwpEwICpzHeWRp2AegkQWMlkPc0uvB3yHypJs6qf2sBYcC+cZjF446
P1dQBvwR3Jtbugx2Hf+S/Y8RTHUkEZoAYxmtBlyJkjYYjw1U+v488yOT1Q/KIIGgTBrSaJgzY35t
S4nzXyv2LG5svtriyepgR5cma9G1NdprhwbEKO33fytSo9uB+QWhjndXKlpyooixSVf6aRYVXRSU
WZwelSTqW46mtVgeelSxmD4xUc9fUwIss1b7eC4Gk/xUVrqFGP8TVh4tmYcT+7lvu8CqFDFYyN1k
0aMKfxm38wgJvL6Ek/ujzWiqHqpBNFD0KFHOqaoh7q+ezaE2PCdpjzMExXrpihow33DzCeyQgfcS
LEF07+hngGOK/MGblhmRO6AfrcHhNS7Gypiv32uG0mDP081PQagCNdy23Ju2jHxKhMhs+CP9zJyp
ZyNyPak6fvyJVFeYrDXB3wRe8IkSlQs2P7cnxXo/0DoPVaNgp9u6iUGX2BF+e0CFxZmgyMqU1T1d
hFfYxNp2li8Nhbq7+gwAXDVrA1iOaIN7neW7rXRu/o1KQ7hgU9rHJhdHDzQ5K/PdOWr9x1YbIp7X
rm/HmLCxHpdotPoa6U62kmrtdCwbdlpXeAKzQNAQeQRkfrdS/f/s3L2gGH7UUPo6F5hjPzYe/K7B
MPSqiy7sq1L2Pfg0KJ80h1YFNjyirddmOV0LSApqAIUdJbM6DFmaUjf/CWFWCdR7xm2jX188Ar8U
oBDr/Az6XqoiPmb61Pf6ClqRLwsHh83alVJEs9cz1/GEdVmNA/71Aph+VvvM5zU/GU/KliY/c9A9
jjcu3o3RHaAa5w9m9fZLCepucCinaEqPdi6oKa+F8aCXb8VXil/aRkDGEj8tLtsBxYZRw/00u9Nc
waYwBpSL6LxssIYQoqDlg54Cy39HaaOLzryHAQfjoyNexlX5pkE3hNsJ9vpHcPjhrXmbKXx5FUaU
1cagCkpV6vm0X/HaxpY5XiZZhWFrEASaDR+nxgaCovwyP1Wf/Weee9663w91J0bU9QpCAOlxUnoC
ULUK8HyE7geq6UaDRrQnqPrC4cEzo74S/4NiMOpNE+jMEcNth9viYKvy1JBmBHolLGDd9gCYt/FA
h7XPYKqs/boarHzVT0oaaHNSjeLtzscLTq9Gb1a+dIU8NaUEZD8uT+rKw8LAbZVN6Qo6/5Tp3mAH
PwgohPfsRfbJ9q2rP/UmhXxeEMn0VULN2nWdjZ936hCR/ZZx9cFlr5SmCabPJfqrLrf2FlB+Eh0A
2tT3l5J1q8UiRtVeZ/NCDhrL2d2J4+8xjivqNFTs1TtTTKtNadQmXFoAqSrUBl38DtvUDFkA397P
SkJd7LUV5zzYYYF4zzirI3vxReLPlZ++/wQPvLshAYdKEF15G4wLYdmRe+VGZiWHYEohu8dKGGOY
qcsIUhRXivKFP+iJ+bxA7ne4qFUk8+r8l4XtvmGlbqKJNubpijByK7+Xp4u1cGUf6/xIMUuBWW2e
//TPvaGEGRj3uhPpOzrkEaoIIXetojjFDvFNc0Vn53ASTGb3Huj07GlbCxCyemFE9bUtuyBWSf3v
9cd8kKPyF83V7i3YYA8ioe6Ga/5hxAMwnUbO9bRqPYH6/V3vtCllCGGPzUbDjK/UotbcwUZ0Tr7G
QVj/2vg+vcZsCbWyhjSDo1LWcNVpEezNT1tPHloqKu+ZkaYfJjAq9OP5zO3ehteccQhYbZikvRrY
RIPDujTnKphfuknSD2QojUVugGR1UOHDP243LmyHCdxMGiDuyTYhJLKmpXlGOAWDZ0U5vlQ3cyXk
CNqeausaJfZXU3eYlL17yYtth8BQv1xRSOwWaOg4mqDxE3ZnAJ7JoWP0d7OAySpdbzmsmzvs3TU0
g+1EEmSamuyO3QamSHGc+LSOO9lJEcJIswt21LDmliAb7ht8wK/wNz9TfEJTrIZJKrkiM383yh0v
+2DJiwPoNq90+/dGy2kwPm/3NEuTAQfC30sFUIq5+eson97KWQers9mFcRnYn9pFan5AWGl4vnwN
sktL0FuPQQhLNYcLFCpTBMRrow2dYYZJzPU3dYzq1am+zdmwqoU3jdfBG2uIuHNGCzhtA+TGurr1
PEZB+DmUnsIO1NMvNsmXbVfk/FffEi8lDEF0aYk6XStN70gaAQkqks69pIyzmW1eOzsCOHwKSYGO
ee/Q8qHHEjlIH584SLjxLcY3q5NdhOpWl0Fnq1Kgg1UdHiv6KRdrdHwKFav2qtSH9HYFynb8VcFh
kXr32aIv7599DhroiLqtuomfa2m7qFyy3Pc5U6fuedF0RTTGmdEHOQ6/fgljjX5C7epV5EVBcgnM
M8m0WiLboV6S15cTqiqR0EEliiQvctTHYZmxySfu4QT2WCQGsVWm7eVt0IBbpYGmmZKt7bBeM0EC
NRHbO8qWMGnOyFVYqiTLcpnwrRoe3obtXS6Nv218ix8+rdB/9BJ/Zyn0vsg+IiDogzOYb56wz02n
rQGydzqxim+x68IPIU1IyPusrCsu+ZF7YIRjGJd30ShNbeWhseYyTSA69tVWHajwc9UZhTIQxrnW
FUwuEjiLTk4MJvPlcz4NrmEv5/yk5JQNXXC32p9+YLL5yvz3GLF3nY1pdVkrxDKth8KVFow/8zaT
YItegUbwMunpTde6klXGA+UWGk6Zix+BBPK2kHXSy2XzNTTd2+bY5h+4UJeHK6uvzsWWYHAqccjM
D+nxh3fsV3wHvy6PT87OSKNQfjX49l98xPFCeTpkPXaS02tM8LWEwpYtT4kyRUGWzCnSqfpJI581
IGYAW5mYDrLNeSTiCdifbW/26ZYTi3tDOssrMUhceONbRZTIleK1LxfJFbPoOCUcId7IcL9+4y6q
Vn63yHwG09NePg6R/omnflmnRwuL6d9gokYHh0Mfr4IU6L2RBOs77Zhu78Kck3PkonsyP4OImt6f
heDekujcK1pN94SD9w9EnJm1zoTr8umz/j2ZfrjHpY3eSlsXX+F3yI6qgKZVIgjtN3t4DYVJnfev
JzrCCygmwi6VKpWhEgXc+KaArOWy37gFKLORDdLweTOEUNLo59FYeeOix+qc0+fUVOCExWFU7e7R
leSkM34j2UsVi9iN1yzwSBsVpkydWuDWSjeR8Ge9wIObNhCuiMpSFEEqAFC1osOKBrwtftvvBMPw
w2yvMr5bYgxoa1uek77FnKMUk1+P0wUC3yWKgh25RrxMscJv/B4rrika9aU82GpelMhiNJvE3L4c
zkN9m+M2wGZO4QYcfg2s8xGxNHXsZnUqyTs6s3wBNUjNXy+71NXjLCVBA/ql2BA2lMHLk5tRhxda
tdzk2zEBmw9mZMHb6U+GGHPSC/IYZOeSiPokni8+iTk5JdDq7dWaB3IiEn62BSGqZ83fJxQji7Rv
F5akdzigRff/4+3OSbSMN3jVcR1sPsGIYYUSd5vKWJ7WLYFyhPpJC3wh8Aj/hXe5U41OIBmK/3Rc
RGiXs7ZTrcXF0IVBqaAuFTeKBJtV5du42pYMoccSzABWw6acImtFI7ZZwZpPwOd+X3bBvEalfs0v
PIHG+ouluj8C1yrmlmaWldUrhsAQCUU2ZN/HLtRw25gNG9M9CpOruU+TenovfzBP2JyJae6Sj6Ni
FpeSzxR8dP/tE2TBVCOecU0egWfPL107xw4X1rx6N1DUFztKTpmElM3jDl2Iwp2Qs1nYtTFEU117
tgdYgPzYOfsWkCTsKWGdxaGuOKkIs6RvyiHGmREsa44Lq1iSCBQGMIf+kYm33uR+4lH6i49e0w1x
j/Zg2+fu+YFRw6bYfVY03G0s7WtKBwL9hWW5vUTB60Lsc3OkqYiVD7hei6Br2Tutbot5r99cfhX6
gjMGxRMpZRiAKY5sjjU5nrFlx81/Mwsah1NN8HPybZ+hnFiXkkQ4mhwga2GcFm5cme5OT/v7IBb8
QeuTvhbKBt7eEuVo24eYZI5RZkA7Qsnrxi8ZRFZcSesyMeubthUAGgpvAxKqSfEVmRQVpUJZhzUO
aaMRykRPMbvWKJ6siJIS8hlTYppn6P2b0Ot/q5y8lZT0fGpjOh9aCmQgQrMn/yRop0LaO291Zjjg
7TmH0fEFBB1Xiq07puX1APnZX38kNvtjTM2qhbal52VzfS5waKuRGOJ7O2XawDB0rXZf96BSUv3v
QguYJcjeXBktQLsC1ln/1P5e/FMNR1hSczeuoumm9bv7Q18eldCzknunpo5dgtxnUBXAg54fyszG
jTR2l2Zmibff41n74cT/EhZeNwwv6fHgmDLBVwEZUfY3JQCN3xnPcYLhuyNrIwUkUqaxbvYOLdRP
MkBvtBoUB06zXW039nORcDrNqSZ5wyQ8G5HnP9jOboMcq7Pk0hW9GlJXaKunl8kYCoDW5MuO2GB9
0ruxLWRXe5/BRVpLMBXt2OilJ6QEFr39LnFOdLbWdw9rFfrSkZYcyZ/bKQtYfPHpU0JBI1Xoq3l+
I273ZkMY9rrOX2zhqOZXPOHKw7Hm35UCcFDp6ZfNHxrZUz/qMgfNs1V7Ihw5ke8eE0yhIDXFT1wx
TMfBhkQQKf9NX36AowyNhSMu53iYgQuqhEMWfI5B2oSJZYRR9KK+YqX2NjqG8rw2F/ieBlU23+qN
vVwbNUx7D7fxIqG/P8xt+lQmAa6c/JZGfQhsxICtzrO3Adgbpk6dhABW9Tg1e4zuNcd5LI7XEq3P
24YDDsd1yHDojVRU17G4lmQJzKehuXYfPTn0BvuaBMPsP5w4tjL3LWBJzbyilCi5qygVhLuboS+N
yT1zk/Ol88RMhFNOGxKmBljnOrfBHz2t0ZOsjvh5SgEZkYUqOUZ0JVTR7AkXSy4Tfy1IGu6prxpj
m5N1TY8fmRUD7EhN35ubd6Ls5WcTZZq0iRNr2GDp1C671OiEM5qb2dLROFXwtaW9ycySt81uSc/K
i/n03faIgNq6v1OQ1W+3k5FwxgVgz472NqV/2+CfarIMo6ERhSyBZoAx8AMf6t1DtYYsqqlSE19G
ql1LWpE6fZHUiZ8PlH24aNMzCKPI4pTjNwWCJ+w0QRlgNsfz92bdzVjoOI5Vr4+SciZbo1ZT0ZXi
DWhEnVl2Pk9/MaCCmRNc3qxZL1gm8pYQIT49D5kncyq5y3RHi8EXwU8wpsjxPi9ctWYVcfgS0jxV
7iUcW7jIr104JUGAq3WsHvKQ05DskPlhAZjRdt2+aa2CMw/3/DJaMXaGWbNF3qqrIarQaw8efCDp
u8X27/EAcEqAK4zaKmpIol1nyaLxIFFapQMmm0eijKXQwwqo688QxBo2aAPjdEIzjxx/U8T4Nk/+
Nd3VIAdx5HzUfg/2QzDx/SDotAo6SxTsgGcN1+HDf5dF7eVsIIjCPmLv84DoAdPRUGSKU+lwc+Fw
XkfjEH/nzSeG0W453ST1+ND8ftwRqG6NJI9Blr0zAzgn6iBaxCMr9aYH8uaykSPHAb+BfnTKnxQH
ZxntpTPvVNEE/8KhbnjkP0XwPiez7Bz2wDIceJp5EYi0DLOJM5wKxty9NLuCIQKHECEb5Lf15xQW
5fQ6BWDUMKngC00umeszt9EkAYfHVmcewKuvQZy4QUBKaJKhryuQJYAbZNizM3ORMelFdVMWSGf2
RkVYtzyjad3/po/ndwr5IblP9eafaPGlc5soOwoOiZA3pxpAPCuzYstTK/0aB51ks9n3yYV8RWBN
P6vDouX061yAsLc9qKVYUNtgtSymHxYzfy7iew5UiUCTStAWJZ/G1DdgiOCuCz3EzJert1A5vKJJ
pI7nS7ZriyVC43kKAXDTZSC0obo5OqvPr19Dam5h4CS06tNzawfec/Ktjq4LpCEqWXBoDEgCK4TM
1g6oSdGuDJ2tTU7eudOAohsEFxvV8dGBJj89JLgALTNJYEOJSGJ+07JBTymsWVxXtJan9vRvBkUi
bV8eCb85HUUQLYRFsfwrGOZ8UiNFNMXH4RXVFNLmGFHaJP2dFR3UoYhG2DPb7VarEeOFwfhGd6Y7
Jg7chUlQZp2XkJDGylDzNqb0xwJcWcrL5T5Bg860GWHMCUL2TIXRjDsFYSrct30/Kjy3q8OgpBas
SdU5dewnL+o+INRW83sbKNmJurtxyGo3RRJrpoA157Dh9cOUda2zS3HURziYgsUyYNQi8DgoY3kT
TdOlgagAfS4KJ+LumTL/YBkoU7XqwHvINjWd2i3vymdJGJN6lTK99u5E7WQH89uYG+bMgTNqn1Vb
qcanOPIYv18zK+ghPd+9fnQbFnuz2VVdVs7UmNJE02DFgjBaKuyyBwXL4IGYSWUXHBoEghXorIri
DO30gJPQ7CXHw+PpCUAkKaBsCVuJRgADz4WG872rrTpaN3ACh9o2KDIG4H/Z3hOYXmO3oq8yXbB8
A+EnXnADLpxnxETc95QdagQBlX2d+hKrM3VVBMkzeK27slRraTP3hZIXyDNK/fgGwMX5q52LVzYL
zuRtlkTxRvjBS2n7EgeUCT0mmZL4mRyI8x4OB8WSQrmzgeqM4FEBYZSv+QXC96luX8rYllU09tGe
4+AqblJKTIJlWejDWgcexdAYyYHDuN4p7ekWZQtN14PNksSCvLEouhLIoWp/rXFptJkflvwL8AjS
9753weVa23uEDU2SGQiphHVYAIloLwMEb6oDrZn36PTRIBUf5OnNF8onpD3mrOiA2DvPQAowcnvQ
9OcB+JxVnG3Br0HnrBdPn2OAf6vBR0khqAlz8dDufyy60Fr2jHWgEwQ0enugwFhFRBvG3Pks1Ra/
yxjataAnBWR7USgLEQ8/PTfLM9ZIPkUQDpuLJSYVhlAwP6RH3Z+LaCX846Ud0H34ImDJgQwT5y76
svXL7bXp/3ftu7+Sy87DdYa8bghGEIuv7P9E7QOz5YgFGza4gIEUtpxIXa5hSX6u3dB0w5l72O4K
roz8itD3YzCrbGZCUmPZrv6vZFW22YkRvH2a/18f3+jX68o/qRJgGUCMEaXuoe2ZKIAJfgQ/+eCf
qTJ8+RybZvk/lZUE6PEs36DjCHNSLEqHRCBsHw1STEVkOMv2j75pkU99S9hwZaSmJzIrU74ohe23
f84W59rmIE0THdfETKZjXTJzQFz6XG4rY4+X6NrYl2w5z8aC+defCYsmgV6AYouU1rkCub4go2zv
9nl1sWNGkLu/SZXPdDg33J3gsBbNsIw5kBQdjwmva8pv19MrdLgC2ZQyN34JJ8bmzWtp0YkmTfoz
UtJbRXqFKS6SnpBKsoP4tpnl1G3Dsz94vQHp6gQedprAXSTT3ACZVnTEPv4fKcyCM3LWkhADpXp0
Or+e7OMFDOP9kIA7siUXzZUAc9oqe+hPBlo6awNeOm1VtY1lTx7DqNbj6i09fLlNkxYKLUU7VCOX
a2hePo41990XLrpendudR2+vSZ/aF6B1s6ViWxu7cMfxW5rE3IVD1eaeA7cJ6fVGfzvzIn2wfThO
pke8PtpGoVCAkoNTqIirNC/3WmzGAOozjpxqGkJk5ugpyAz1mI/ZG+yGlneELRBwttGtFcyrAK3G
uRLBV7GU4Jz+Dcjz5K2bw0sQN3xpdsD5iavRusOx79ewI7dO6W/C903yP2CO8nLTqPseqzHrP2Hp
3Iy4AqrKvLHEI7D2gug/vpaeb4E4vXr/aPPVqMecdQnTM7gAt7+QEB1RrbaoEPqYOIhBsai2GXRi
tWh8JvImnyaVO+dWRNDOx2UAmTyy7pdRz0BB3szAw/9P68kvQUQtHdnmuJx1UebnMtQFu4kHSmDO
1oIhIMBXF9HNk/otGjsY5KmjJBuURV9BVNtasFQT/KrRb/B7HHufroPdHkv5itfClQInCfQJ0cyb
jo5i9jKXkwX5tx1I+PclDLQtkag11VfwoK573FCcsI59mnIyUIuvpFa0c2SC8togFHSQCmP73GyT
EnpLFYDIxlqn5U6aIOx9juCcvCZkwL7PIn8uurdy7JVit8AJvKCSBaKCsrbR/hsrhWfOkF4BWfyF
jQ7tABOsaI+iMe9TqM1s10VODwB/RH2DEVXaQi5G393/BiJjgYMwGQAuXxY99WJCFtzY4+/rNs9V
4ASzgfzq0VOW4mHD9INIyqh6HO3LBVdCGtcuu9ENwbG46HWFCykHxgVILWg6yBwYs643fjV8+LNn
BOtlchWjbiwRiKVqQsfvw8Gu91A60p5kUf3118jrf3XHdb6H6miPAaGWyGp362CW4S2PgyG/FVJf
15dIWO6IM4PgJWtQo8jwbVBPbSkZKvqbYqipC0Zsjp08wODtDpgJjoWooI02JhNpMAzgN5nRWzBo
fSSqNe9i/JwAM3RIA899U+cLjvMRsQiPmW6ghHvLx3gskqD8/VoiwFW9lhT+iDh8sOKx9UWqBn4n
hrk1mKyo6WJzXab/7zuHnjb08F9BRGkdt1KXunuF9QYBJ+cl6OJ9OrARoV4iqsE8gePbh3SzkAoc
QTgAoyfc5Mzc2gSB9OSQFFeCZrHFzv7C0XwPZktq17XqL02D7L0E8kMY2WIbqAV1sXYYmneEc2LU
0O9KckuBjBx9E5mvzeD0ogi8akmBQPZQ6pn0vjPPamXIPMcByp5NVCcnWpB5B+KoPE9IcqEbWozZ
qxycDzqCNpA4Lks7nGFKYoiwAs7VK83iSYUVXb5qmcx/TbFhRTh5voLRHGdsmC1Mbhoh1S5Ml+8I
ZTPA4824+iNue5Ys0uFFi5j5zVzn/js3shggtzoPK0vJyXaQiVY/c+4um/m7t8AyiDCktqKndall
xuNQ2oHzb7aP4sET4vb1qQu6IHzL96OSwswXj/8misI+21gCA6ryQCMi2okZTjZD19LPhncs57Jn
cmvipiws6FD6u6unCmIz2bMdc9EPmVvlqM8nODSzV0yuxhEEHslIaerLYwPPeos9N+Fm9gCQ4VDm
pWvbvBM8uagKmYv2e7sw58tVAdqCSznylji/AgG7wfOCD7kOg9KHubtrCVutuRM8oCczkY95ulE1
Xf/zp8xESPNihZwY8NgyUZhZZU/ourldGb4Vt8Dg+2P6S0KZwCKDPXpqLULnatoZIsdLuEHX6iYL
heGyY66BFiE2ZPVrO6czKvO4TY6rlS8Be+4DumMTJ8avjnwOxBoVaw2FVsWfK3VdDFPWZIq3ZrRO
6iFs6BeIlVWQdfXtM1ZvISWc+Cb+quP+tJgHOsXqRkoFWZRRxa3Aui1hZQGIhC4JVnsEyNKkqkHC
NNcsjYv69GZ/vbGbB3QUYQX1ieM7k4OrMmQrp/pkX2qWhN6qrEdWUloBR+/uct7zQPaJkRvUSZzL
6R7o2+jBtL0ojM7yRpLZw8S65KF1m1+hfqr7H6UpEe5NSzJodNGBpBnX8jYOf9UyeFQ3SuC2Vt9J
POdfG5PDvV83TCAJV2kdQ+Vu532QigJdKcqHyVh+AFKbbBGLDCkuZhvoPkWcfZdPFMZviFG4f+OT
cd/3kg2cRGrTXpLozF+CThTcvoifA+WnMkT3v8yMX+Gb7b5E0UEEBUFJuZjzKuxOlAFQFgdUT5hu
Kkh88Q1jgWTmD3PtRWj3bCvAUMwFtkq8ULDND0WcnEw6tBwjqiLiCc0x7WoLSbz3UuFmUG0ZfAGy
tF1q5q9rCqiEUyE+R/zmvG9Iva6DeVWEEmqDuglBVmpYvpg+wUqAfr//z41oDhfD5GjloacvSXJy
tUc7Cyu/c1cKYcnpVu3rIdh0q9VCRCAwdbTh9ToT7J9g5jSgMEDWJlFV/dtCKuP1VIgyD6HC26Cu
lo+7dwoIr/S7kdrJD+doTp3LtpAx8mPQ/9nLt9IG0Er1jflQigP2p3I6UnB7yK/1EBfUkNY08AcG
HRHPZTaNAXlkGGufYYuXtEGpMkHPgSGSE5xyJAiH1wSC3L/1suSriar57r1+fO7uTX+2ZEA2H4OD
DgMcUqvV3g+t5wk=
`protect end_protected

