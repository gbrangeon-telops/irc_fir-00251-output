

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MxpeY9fwU4EddFSpExWohS5o9i8UPinR6kQv/f7rVpVjW9v1XPHFNv5NQBBqnxbGk/3GroOhKYHi
zeZXd9sb8Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
genV68U/jEyVif/FXdfTRcDdNLXMaB4JkzDnEPHISJLebDAxHBqab4xQb3vzSMzS4EZxJxM3czS7
l6/Pa+/lUNH4iHFgH3/d34ImoXy9UrVsNWI4O1k56f8CO5JZkX0ENM2JUr2+jZNnrmepHCpz3pyr
N2xknPLUPWomWT5p45Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
4dyOi6X0ND7jxJKLfQYpMzBQUnXRUvqhIlWd2qdz2OgGY9VUivCAp2239OkMu2rIWSpkdV3gd8Tn
4E+XnpveIi4nHAn1AdqR2yW6qJRqYI/CpvcG8E7ZhuUiWSAPiQ/jcxRmeyzLFdVhgEV4hed5vk+9
Qi0C1DUHqDNPvc06f+xZUSTzBSqXkxyUqGIa+j3ZmCrjq04hmRDILUEkjqmR0K0TOLNdsLd81gAl
LqIfeuzK3hLcVWnnJG54RzS/q6bahPN8UaYhtJREcAC9BD1S+QEdDXRxFczj2T1LQBL5rSryR8bI
LV6YqNl+85SCCMZmZV8Io9S7fDVIrhzNm4Kcmw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PIdLn+S6alHzFt/ir7zZvMPdMeYQTL6BrWSuIGxsOazGugSdn7m2jtyII74LXXAGUQ0h11spxnUf
W/HpoHHxg6pfmAZclwmfvLsFiVi0w0hNMmIWoR8TGPdAC93Y5+aRfoAJNuDfUDfLzdBM4O7G2ZFx
YGYpvBcNhzcFFuSCCK4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KkGw0OOEdMUjhZKEmICwPPGTbEeQxk+K4HH0ah7Z5cm5dbbyDDJyn1CdBy6WY7ZD/SXDbXp0Ibi6
BH7Y9BzUsE3rhTUVWQo0OMHXc+hE0CnmrdIq6Yy3Wkf73IKl+pu+66Qo9W7SdJGNPpreGME4X4AM
zBwAv9xByRwGoY45EIIGTaE7VL15piKgLihjK8Y2Ee8q921qHsI62b9osdj+stH9M0nIgGIwpsIA
DiUOa8Naw0kRMS8QCXDqKr1fJ0jPj3cnclvP9Taz8J5tp8Sf8I6bs8irg+MGD1MgQIfeKkimA5VH
MerNz8gbn3+/Vz2X2+nKanM3LebAMLyCO8EBfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35024)
`protect data_block
Og52LcMVV58lnq14SL6GhT4gh60vfTKtgSJSdL75KymI+Wm/5/SWRemgQ4KzVzS9LASre+m1qydm
IAy/Fgww/wr4l/8gATBuZFyf8wS32cFmpa29FnK7DNhtQZ6pCDITwhvu3x12LPmBida1JF8Z3XV9
OP3sdbZj1/xdC9ORNhpzoQCI83whklB6pcC0/e1Xk9uDfPxbuFIW5FAcMSK63He10GUsZLPobsEI
pW2frLBo7Af/r5qTkclPY5JPxKiYWifWmiiunbzU+RIxOGrzXLoIIH8q+DanuV/jZ6Wm/UXbZqkh
BAep+0ROBJeYYrzYVFz5cc4sQKVa7XKZ9C01E9vngfpxQvIJZk1uaAplo3m7hyu0A3+XSrod8pUP
oj4/7xbptchGG9wMAvkB9EGjuCLaaSSmXuQ/A9Kxg/mdIgb2y7Sp8GT0yehextk+rXnowniJDkxw
rT6LwBSCDTgR3vjeGwn9Rz1iO/7nWaJb73FaQ8Dj0Qp9bJS9owh1VFR0wylSuUV1ocO9oQxqGHUc
yI8ov2s+0oKmluJCJcl9OnMJ0rCyygBP0ilUmkYrjBaZ/xet0wCsJIOUDcBLeyUNswHPauex50kD
wZg25/rhXIiB0dAd/3vlyF451ayGrQX1jqMT+MauO0uZQ/bM3GA45ld+81B7LPqlxcBjt76Aq+zX
v45hfgNxlmePBT5k3rA9orPZtjm8zIDfXu0R2iGjUC3aO7BC03RB/mlYXjdYVkOvC+G60jNEsnXF
9XeYs3NgsLGMrW6lLVy6b1YiA8YxmxHxx+QNa5BBRsbDdyE4sclMvC+EzbeuMeg0B+Xsdx1eNa0l
fX1+SeVhEBJRUnUJm2Cg6HoyutzsRWGMTPDQbreA5I2PM271rTRzDvyLAGlKX/RkwxXz4uitsyQL
vzk++JV462Qh5FA9zMyGpQflawwgz9t8vh6Uhy6YoGLyPJS+FzGGOTf6q8dqFafDLJ077funqbf+
WTNfI1rRRyK1/yL2CvaThK4TyMgohIJbkoSXgwRkx1WlUK9YSZFqOZZdv95ZRWqebNiQasZMjI0G
blWiuZ1SndGP46Jy6+g17R2BeXS8GDsRFeA6aRbENgGEsdNe9E9XdT1gNbKUgM3yDYDyVw1d9cLt
ViSUbpUKE48kyeUz7qX3GiY4VzbI7pxF2902CjSBVQshk1IukUJ2OHVh/yD5CHx0/lWmkd5PUJ3l
KF/hEGF9bsJftOAAjwHIDjmO09XRYgcG719kbVmf4CCyrwFRotWPLMLdt/U3cw66/bTUQ5EQ04yn
S96gEdXGXsOGwFoRDLgd8KvoPAevaFE5hiNWrgk5pWFq5y3NTeGvTDdyZSe50cf9cyJv0vS62hMP
KptJW4g0oEtm2kvbQYIPLWgbtDG7xTvoH7j3qo+fxVIwGV+rSbIgWybZHYHAX5Jkv/BPIoef9yvJ
noQgXk8WMs34n+Frsiy8j0lIIgKWXqoi/DTdKeJBp5qJx6TAueRei5o4CcoJSksXT0PnuVjsEW0G
IwXX8ArCU8L13P6CJHXSC2j0LHF7MSy36Suf73GNWkcdrOXoLOy9R/R41jr7B3HlkFhDMB+lYmTZ
qQFyP0JdPqbOAF2InR2KRgYASZjUzpfvVV7ORBjw/nhkwES3GDurMty2EGcLd3RG5SGQWzje3oCk
um11NUx9+6LnHCNDdp5UYYYPAJw6ZLJzByuWyHAZJiRJ/LHOisjwyTXC2phbo/rr6GG/7ttx7Rsd
ZLDHRCy7Qkn3k6U2zBmU7sPwEKnwn+9VlOblCCcxKSfL1iAA7OzpCyCB8HV77r3ZOYXsI5MYCoq3
wAHsmYXepRhZBblTWDSHUUsP2bHxR+++Xe2Q3hcU+sX87+mL3cKxoUHav5OmeIo226u/xMiUgM3f
Lj31TkUQ03y/HorMECAgCvYt+JvSei39wEbqV0+Wk+JIJqdioytU4Zw+wY1lDUcz5R8hoB0/zQ4v
ceFHOUoQNQOr/krVZjYjv69LXEJLZI6LjPlClVZcoRFx42AAb6rYg+QhetHb4hcDMHaMey5k75tl
fdl5X5W3cirDyqzw3/yQP4ZEpZbId4XYavdVxcPm1vsxlHb6nYTSUf7U2sQh534F24mkz4OZdpFz
Ld7v8GseWZzU/dM6lXmn2Xz1bc01SPU4Bg7Nyre7NVAsHG7De+g9sKpzAGZMbPGx6Zb1F9MmyQFy
/wZe0isz80Pqc5fGd9uyuvhTOr3zR874suk0ZWSquV5sOeCWEioS2eDWegkD9BDMhKtOo2FazdLz
/EG9pqXXCfsXX5uUHbROx7NzKwf1qbzqra3TYPwkXRGdnLwZ9liRSn6/iB7mIqpleJdpZCmHTsLJ
M7jNtmPpsvJuDFnEF5aO2xeAtj14WJQLO52bAtYfIEEYwdfX9A5xIwnUBcpqd9VktGhNmn665omZ
4Qw07sI1Ct7T5Sgjs1pHgnvbE2wauXbzuS7jPcccawldejgdzgQnrhszs7v1ZgCbHQEzj2h8khlb
3KwrrvpsV/d2txacTrYozQ7jfRTJbNOmo6jlSl02aVcyWYww4PTP5Rm6ySqKGI9jCJDYWPbmYoLl
zLJG6+jeXJW+js52/2LEdLfVtqagUiWYfCMPvhriPywSuBTw37yK2EJvf8M7JPajsjY6SHv/T9+a
KTZ+RaA0xFN9Yi1LQluvWa3De+lvs41o0WulX4DrdYSK/Kl7WL/+Gm4BckPE2U1XnewvB4sUbQCQ
b62F/mROqKOuUm8vIkxIyKmqmfS+8aFMkC280ptCZH11RpEYrh8EMMiv02cCpyYnkQgTbZAyw5dg
lp6BHlLmGe3xAFag1jKpTU+eWw5xw3loSdRZSuBq8BL7DfYxghbXL7Spy5tmbxO6aXeQqSVTY69O
xfFy5oZRUFQWDBpDKGUhGCx7oz95XgmTsDgK+jAPmYyloqACHXaavmemUt7be5fa9VUhAqDy46Fy
o/r1IbGeeVOdqf+jDupSDfnaR/Ae/e/9IZbJbkeOuiPU0ktnYg2WQ3qVLQYh1hQfPzlH/RWtxKSx
eVt16tPVGRKv7lOgvLVMykc/j0pzh9k7Z8om56t49n928XoNJ7ThSSvLGaopwBLafy7rskAVH9/f
Y1pooRp9pHvugTMC4r8fxSet+zLdzQTjNch+PgjjN775lFKq7EJvpZPppZKNSpQ2BZ8O8UWxffbV
NHDwv6B7FMAxWzD/pzLVGAA9ZpAOH73WJd2hmn/nmzwHz5xKcHJwY6xmGlgwvHBCT4AbuUgTupPB
g5R7Dw7GJdJ1hTQcQm4CSGbUIJzLy9EEcN3RlOyZojKoYXhigfb/6/AiHEVeLDjBfhzfbild5Ne7
AbY+itbSH3o76k7QOw29HiENknLoCn58qXWWoIvEoo+4PltqxJLvdI3VjUQGYRHFRonSy9MjpzTn
SD16Ly6sz8P2iA8GsmhogpTaUVHuP7aZCXn9Rv7+1yUQXbEAN/wXBWfKQXyULhWbIBHtdoaTRIDM
QoWTpQNN2sBWvRP2206toRDUjBXOiUXDEA34rlQk1jckb3ZOPP2+WZu3cD17R3Xxaj6KyAyjxld0
gZAZUD+fna01uj/iUL4kzep5DLnEAjQ/bkYc1/ObZjtsThW4DiHZJXwCXtM9v5tNXAv7eHmqp6SK
audaUAO8JIemKODkH92X3J2OeSE+L+PtX5NBmGoSB5njqu8vySBg9eebupvvfrzrTixW94M6Ot1W
+o4PwVldNaMWnzbeV5sfzh+qCRnk2VcpSwhyCLs6MARltiXRV1W8rYMOWD7r3bAHQgcje7LvnnKM
DEaG7c4RKUfQkE3vztrzauOKQCQ4Xl1afDEwWY99ZZx0lxxhOvwxcKw9jslifcVNvUkKFbzjPw8g
Bs4/t9pk4wNg4Vdb/kdow5PSaxZCjA0DR3T0sNKAUR/qHfj+TZCQ3STvZsuDtjbifPY1Xe4QYfhL
9vHrdBz/k9nGHqeU2WWLivBZY6yRM84AAQldXlexXXXu+peq5sXmGzdk8+d+5WTuhztCG5hlqEwz
zD5ZfenLjmEkq27JLyXvmn5AhzYvPbfduHotXRnLrxBtSc+m8szHY443KXYlStr5eUP+kQIBuSoJ
qP7BHHVQk7h0L7oNhq3PCqljgH2bt3ZeXUJq3kftgDWKr7nnrBV+D+HN628mvaZb6vDud5K79jmj
HkRlzQhsea9z+93Y+tW8BjdVlzgb1wWOMGLfmP6mcTtrfC0t069Vx0nSt50q0mvpeq2C0AeIB9fR
8Sjg0JW+hX3CQPdpygMbiIF1kPdXTD3RY7hSD6lXoldkJcdJ4rg7dOXZda2Q1m2lRTsiqZGoao7n
6FiFZVaK5+4CVEFU4XNXUZvnELmc+YMrOe5UKiIDbo7pnS+uj9zIsYmeMsG2adHFt9/MoJ1UUKsO
DHI/xqeZvWB8QxPwJmpx4iT+rYDYQlsg/uRM9Uk/ZPBRtKcSge4TrAz6WnGw4QVrZV8t4jTWC9hS
TzbdP4JgBBj5paXKu2GDL2i7iEaFtdsOnTgbqX2REaZlRYhkMghm7ojsn8dn3O4xHNd4a6UC3/KP
nocp8RPvr5H93vToyBi24PsgCXmx+zUfk1nujYb86O7xe4TQiG0ircjJmgznAQEiMo0hv3EukRDU
2DskeMbIvts0+hT0JwoHrNzcIQDxtOUahXyYdHLA5hUrqbGFZHyq6ODuxPg80rdGcM3cm6uVXoXW
RYIrqJyAYtzxrAs5p1ZzUc6tgepRcQcl/QrpVRYwf0axevpJZU1wiqV216bWJSXSGtXyu0vBY7Pc
s5OWvKa1zGKr1WsqzZRz1gEdwm1EyNBadCR3ZFf6aX2NzMmpwPKbIqsCiNuGvQMm2kRX7u+J5+32
vpIf+i/Rd+s60a2kzdB+n0oGj9+u/H5F3611bdI8R/kDDRAw5fIx4kbRNEk5JDGOiJeqE18qBxWZ
n9Iw+vGxUX4FoPTe3wIbcDumOZ7j36rxnX8zsiUtTWBH30D5ljJIuQJpBhHXD+T4e3ZQoNnORkKy
192iDdI7IvsAhFX7gbJdc/ubxr42PB8G5mPhKMK2Uvw9D1cb1GxjxS15fHFYiAQn6mxOGcaje96i
KCrmmI1f+TV4xaIF7tZVLQ2SWoxae7WP9jBwCQZrWufX2JTEnOzflpZvdNmLuFGhAacmeNtR8GSI
/ZXM1v6cQh6zQ7O4LoTAywT2FzmoWqqGw3j8yduiNi3FH2p5O/QBI9sJvIAulx4g1NM+L53pAEvr
W1sIwGW0ZF7SbXh2ucGlEu3n/p9CEOyM5CnJ7DtI9kXPxyjsUD4kitchXHfrFzCNc/C8n6eO9RcQ
2beWK+JYCT9pXkspiz4WoUASYiHqQNLjIPYhqW32g0jjGR9ItQ/T3zeoqaMfMwosd84llTYplSL5
pW0MuS9zzd8XffQNPQrth5O0zxz/EPrD04/NjbBe4SLf24yIrhoDRa+95vz/+UkDnDCFgUAoTnvd
CF0rInPo379hLBsIgIqk5J4fSfJvC9x1uckW4xq8JBNb3c0kQPASuiBH9jAlAEL+kRq6sdtBUbeC
mOV4m0g27GJpJEuBuiUNXNppnTPlDp+OIvsipzb0oOjEDf1JnwkY9nZvRhMsRoJRrX3IWePXdZOx
urbv7U3Jct03IcuqG+oSvOmxfR4Rn+ZNcmscMllS00VMb6ZQL5OXhY1erY+KdH8IvPBKFay4v7ZT
Lj6ag9EIPpsh2B27bdzqhtNl1HOt8L6B2vLaEPhLKN1NA7AK6C7XbhR/+GPdh0yVDajWxkXUHAPS
a+hEvcza5j+MMtxGo1vapSg3996qNrkaNElJUsvZqhf+DaZ8aKRUyua1pPz4CxSHJtQmAB4QoyP8
xOY9RQxBfqJgMTo1Cu+F4xpBnqztfgD4eU2DDgaRaM9+67p+WQrWYKqEYsHTicjAwm+OBAWp8krS
3+bpq84DIymTNeSwceTnR+uqMU/LGMfKp7pLiHe960nGC95y0zQf2VJ2g8VX19ceI9ucVhYphUAw
2m7W7UU1xrKFNc65oM7PZ0FCYc6MeXQgjeuakVIGmOnD+LwZLhYpu9QEVqepFaBKquo2R3IsAugU
aOCgpaAjdKXXmSGtt9Shi5PDcPi2AJm24gQ0iYs4lOWkOQHgRbsBFrPSr0V0lVl1hAjUAWIFrr4W
V6eGHlD4zXndnEdGUZJDqTIUWOsB3O94kGecDFKdWevQfsUEY32lFJYXdr2KMCHJSECvvKfKUNKT
c2ZasvJmNrVmtaQ9x+BaTQbG/vncBQC+wAlo8EeseDgy3Ul+62ML9WGPd5k09Et6pesLakkgTTJT
9rvAfq+4EP0GN8O5Da158fLgme0xbiAXwxz5CPtwE6jy0YgaA+Vl80/YB9g4TM4IgOv9L7O9DVq2
XPQm0WYU3RvphGZXfFYybNqSac3sKEF3pvRKba+gzqIgULjT9FM4xJfaUlIbnBJrCNOCpGxpf5vH
SYw3lH64YAYI1chKNgInuEpfUSlExQufyHuG8jJwBc8ys6E/N8qJV3cA5hlwdH6BXxDVui4+IzBP
ckph0PYru5+3dGUWoO1Vf/wqXjeL9Tysoyj85Z9Rp/ce5/okIkO8XU5biqg5PYCoTU+HiuWbN+It
VkxUpnbN0eupMJMPygCn44eG4/yd3GLLLzHX9M5nuXS+wvNLeTTYOjpnm4mgUreNwFM/4jqaLApR
LhL03WDVk6FRt56yBggFnUddoEhaofBodnKE8jNetQ7GR2B90RuKG/NeyDv7Ml7wZtDK73RE4Aoe
EhovjW/4KRbx0gr9JE2/sf95zhw0IogmKChyklgaww7bIw9hs7q6aQY7/1lEqMtKfd4vIAl9/H29
NHGwjgImq5JtKMwJcPyi+ZrEw46DTGGUOlIuSgzqDK5pPibSi8Noz1VzjsQBcGn4xeG3H0Nx/1hl
UA/apSOEourhIh9EiULSaSDhDitxMp1k4/Z5rWitP+9H88HruZthhcW0dbS9us7wznwhNftiaJPQ
xUMQuopjc/2Yjpv0AxC92uthA3rUEEyENcKKuXOq5LMRO2UlmzRwXB3zfsxFnDsbOzzNuYlPT0g9
nSVXJEpJ5jjZp7tVYhste9uoXieZvMjEqUDltjv3s937haz/hzY6B4RwC7dJNdasCnROMOenYxvM
qTBv5qlVk4E3txFh/Eclsh5MW77Nv2fqLE4cd2IIuBaE8ivt5sZ5QCnbw98wL0ohGcr7w8jVIJFt
9v88pmZRT2CCbBPxvdGAYzwMTYLAJnWguH/IDslEp7h+7JFR+IV3PylDu7WyLZQCEWdCpwBdc3FP
xkcTvHEmITM9JEB5fe3cLvmKY1rmD2EQJpaVHwuTjlZjvZlioADxXOl71zgoRJ+j4E+sMdEMSjYo
nevo4T9DNEBz2D9ZnrBHG0RvHF/bGL5GiMpZYDeIyeA0t4bLBZeg4H6avzd79dA+rmzfRBQGax4J
ZoKH63we+VjTGgJiwzuDIb3V2PSgI9jgt0TCoiK1Uzx7Kty8CpRpI58lqmCWUWG/DqbGZiq6+72w
Mba+Deb1eJRZBXmRenNTNWKAHfXzDmnXVc9LUjATiPRu3qaRewaBSGeIroB4966A5snl6P1jFnRZ
AIfg4YaTtL380eQxvPB1UcN/+mCeI6MeJ31RPnGeJKBh7BTsTJJ61Fmm51S54Ltn0MhwpX4eQRmL
6DDr4MygwnMWHf/z65pCuLen/yKM9Zfu9mx26Eo70sVnx88795Y0ZhlQLqNPamVXXM0cVQc8dtzZ
SrxVDnETLsgwm/InxmoDPhg/ANmjmxbIVA46VfH3L6zzcunWYCEziH1J/GkPxvdns/ALi52pM6ZY
OaeOJuxdZNO07jDWyOBPdo6F4t2gjtvm70ir1QrSEOU24te6X6DX+qBk5lv+7UWr7DdxBdi+J2++
kCGp7CFVfFfV8X+0QfKxNA9B05WHtMmpDlyKwJXeKacS8ZV1kt4UBCJxH//CNmRNpSsABeV0BIsl
vvuBRwgRTT1FVBZCe9NnmATDSB0uIgvT2cuxMoWLiEPnf8NbZCsdA5YTJXRnJSj1hPw/Y80uzfn3
h36YgOYQXre585EhffameJhSnA4G2mzlLn3+VAhKPE1mtThWig9bN7Ive62hyFD8m5SmhbH60oO4
ku0ab3vHzDi8vmBmuCzBX6Lc9u0rnPdF5dtlpofBdeEdCF5hxJX274G4jCAxt6r9KJN/zvd4Qf5w
R0WhC9pn7nO4+X+rjOPDnVg/Ul7NHm+G8fgLpRLXe7l6dvYqtIHAW6MLJao8Pyh2aJzFrVpP3JKo
uCTYwJUevGuxIklzRleQj6uzlrkrguP+nXAaL6oxO5KlVja9zoXAs9LcjpnwVVQfZp4iT41Ic4uT
VfeSXMBAH+eaeP327CxsNLGYZMVBCcZaQLdy1D2W4AlOcfqVtuPZh9lrI71AK12pJqkF5o5vsvXi
lFzpPS0uq/ze8Sh4Yr72VFg8MVmmei9EFSCnorxcTTVj+/CUjFKs5UgdUGNleK0nNK5UGLnCn7/p
aPSgKO8lSWIFTJxuBAA/QVJf/9x5+5aEspHuYSJSKtKkapJfDD4pNIcNEVHlVr2bs/U7ZIdQ8vNC
wXL+zlgr5XKx8bZMrhzuc/5Ooys6QLYQEJzSLvkdcVzlji3ye6BDe6TKadpQBb18hmJtg8B0m84J
T1QTXhw1Yo/YygLpmQuU2o38x2HekhnTvjKtbISEJm/Jd87kIROMBU+sWB9V4rRqDNmDAzco78AD
LI+WMm+bLp477MjjGEeXmLeorLIMmtAAaDoQc/Vv07pa2Md+FwnLkybW2bQApfARE4AJo8Bc0GRw
Q+No24xYatvjcRoJRn38lboaSOHKaHUyu6k6R+itFGNtmCbq48aL99RNA0bSx+KNG5RLIS1TrCzL
vRI9X/4lvbnSOILpxJaw+TyKFqyDrI12jvTas9DYpWWryXXG3pocTpS9oVwiVFqz0q5bmKNTXYfF
9OCsXA58/iCzry4Vf9c57PfSBAos77CKp7JYK4HxJQ9w/pO5maYvb1p9iS+3IQtu8oGqcIkL3APC
8YkhjWCTRWMqkJzFe0DI3bbZ3YU5LeFMr2j/oVmLssl11L/uYdspmfwy4wfTYgyNZ0EuYKw4GeW5
Sh6GhBUo4/oI1zgUYIDS4Hn6ZZSFBx83kn0VZ7YpKaxDpE+MbNWIvN4snVLMjYr/ARZViU2QSg+1
fyl7BnhboTpswOnuECpzZrnPx9XnNbTlSkHa6Hvg55bUBA56AZEKhu0oyr/T+qpZzgRRiRgOcSne
MPdUZKb/UBs3hef3PDPpVDuau+jetg2fuEGn4NkoRz8fMawfs4+Omeucp0CmOv6dqx6EYwrBgMmP
MkXWD7Lg+95hIY5ZymlUr0qCP3IeNZXVeBDz+0DUaNdVGJMggJXS49M9LFx7/VCHbZfvhNVVeIuK
IdZvzDhgVqKOovjRM0g7MTsC1f+H8VIt6RTqHuYtuMh1mKC2Qbhmrl3C/RciFgbtQu1+tBIN4lpv
jT9wH/7s6l3g7ZdyG1JTiobizaVQYQpuqcHkKq8Z0rYh6ZFtPVFwAKo6PT1+f4p8vLnVJvawjYIG
8Q9DDe9lngmIfHgCRCXUgnMyQwZXcDqxNOOTl9NIfn0gfEoujzRxqdJdXEpJTGYBtm2kAwLOPL6I
0O40OhsT35jA4dEG20ssGb6XRN8sDtDqrKnD2fhnnhfUazUMWbKH9zYFUy6QIrisEOBUfTV2nHQr
2TwAwOb2C8BlTiZcRCqMU10V4JddSrLOZqqkppFGXghQJG7kWGW9pZbhSGE0Fll2b5JcFxeEpAPa
jy4h9L63AS7ktGWCOHFPTLqDWF+t8yAms+kUufdemviBXbgTFSU1tjVW6t7Ni/yuemg2AJn45R7h
bHvlz/I7XVln/UWhGk3wYZg5MBnWRLWom7tj/vB4HoeiLHRDDAygMjJQ5FbszFn1c3QpWgIcdSIf
KD5AECqsqEzyOL+Q59t6etr+Vpyejgv5aH6qIYn8eY0CnDGN5kOLTJRz3uoLSjVf2Nem4+vSZPed
w4/NZlhuHEFlnpPGWs5dNOh7k/YUByix992HPQoe/zVIBsjTPt7UsyWjPiktyvspt06mz5wNUYmn
RsLoLwXPrJD77FpMCzFMv1U2hZ8vCcev3B1m/3o5XWqhMI+ytvxW7kp7rrxZa1lglvOu43Zk46+Z
qi16cWLhbONMPOxqIfJK6le04bla63K0TmTRtVExLBeZ9xvYIw8Ng/R068fBwcN4X4e91jupKS9d
4sHU0NhDFJVHsJgFS5IfAvyaSeVXHeOULA59itgD365hQNfj7CE8AnBhyy53Caelmo09mQ98T81C
Akr1d1eQoMlpP2tsv7jsT2577OIQjonBwNCAge/cgqfewPR7edsWVLV8p6LyM/yT4hiGVxNK+jfA
NCBS8R5oihpkG8wFxnoxnnM12kLXfXZS11V2PwOQ/qvR93h1X/Jeug/svrKeJT+0r//d5vlNi+Om
dNga7+aABP8SqQZyjgXVGxSGoOyuEa/pZT9EZqJeSV23hJO801vk1g1pbDviXFk9y/41hQ+Y84za
dlWIt7xWR6kKFSpfnKJZ3C4XlWcu7njfC55IQRfiWlnbFCTpiw6lNhW5u10nouNUhoR94m7WuykB
SEMxKWmOp4cyuxGovd6zL5i9TYQpqYOKVz8fWKlIIrUG2ZWaOSnG3XWmQpMANR2owJtFChPCW/18
mCo9cIzpjmGIo6Irn8iCThJ1+bh5gzTe1MOnyFcAurVvsm7uNDGxBMPbO+Fk59SIY1kwIHQtTTKN
8nZ2utCf/zsNJbG7DTv8b3yndKPrXZ9KD1dzmhPq3+1gu+h+H3SybdjJo2oUrOpb7FUz93hCpmpG
7IRXGrTzFUpHViZkE0bJSlepW+s+gY5Um8s+qNte9l7rG8ayOMim4V+YJPh5Bij8HgxEfxX2leck
yqSVofMCdXnFyOUUTsJCHn9BkVVcmCS/o8bVWDm6/QubBgk1up/aYKdJaC7EtX1r9Lz1jM8LZVw9
B9LOp4HkNyzmhS7uwe3AYrrf3p5v2MyRGBHIxFhDoSEAOVdsshQnkH4QdK5fSOPvVNtvAg/OK/Rf
iU/v2QzI/CMmFplERsD67PB8WHVSVWhCveW4r4BePJDib29vSP87KHBwnMcnhsbBBDo5IPteKTK9
+Bae5/YFxIBu08bFD/m21Rt+tvUn7/1kHs4tReAvABLC6IHN9dcfRt4cbdMLaO9L4LWbfK5YfOSp
I//j13py8K93695SB146VS7/hyEylUzomWbuwY0luaWGWH3L6+MhKUTQ4UPqfnVfavmYM4cv1V/S
YVwaFm6WvJoRv+3nj1OrOdbEvU0YTwnfZHW8+SDRlC6KnOuCFfs9BIP0asti803iLQaKT28lk+x7
InURVKw1inM+isP5cDjSZep6ecrZ9LqZJnR7yXnSEnV6w1YENHJj2UxHg4P2El7b91w/Y8PHF+fc
UIjVrJ4U06Q+3fpeDtSzd3XzVG8dviuXMlqfM0O5YkMZh4GrXuFlPGYmyYVNxHN9pvShHu+2OJcC
Xi0SW+ucZwfvRGGvHdGHGw+XcGByFlu603rLzKA/EB6fQVdP47bbJY/ATEeq36BX+g4bBlTI54Di
fONdfKlbXl8GEigsLJPGv9VHeYa6hpdhwbVkw9V1u6WkZemGcK9cDmIRJuxut7jg454Hrwpg6mdg
1R7Hej3TkPKWvGUFsMGl5wtmjU6yZvL8xctNxJgtcpPSP+2ArEbwkrSXLWq5F3x2wqLeoYzaawQP
rcmd97btiWi9afS2qe0kfnOwFcm210wlno/TCx8SPUpZzqMk+QU1albMlmgY4D6VrU/6P5c3S0hZ
LX47t2Bwc8bDtQapcuItJTm8v8aMoGfERIdqmF7SHcRhlYHuQgnq9N2tmGammsM362Qyony8arVE
EPJmMuNUbLx66Bb/W6byzZSHhutwTs0v/jO8xVbZ8gP91GKcN23CPdvpDADpC/VpYEtQ2ZpVIbmW
Ej9SHJGoUwDU5PQPVe6a+1B2PXO8NAWI/cV0JddoWpArArwVvS4CfwHWIVzIHeZdKSn0f8x3DNgn
fVA7BTwThCgUF1YHt5OF2osxo+P/zyDEbzDEbboUBsNEG3Vn8f/XqtbgVaU3SHwyQjQoQuGjd0Oj
lszvOhk6Y4yg63Bx4b36R7/d1yATc9469yH7QLM/TISmIg02RD+GhrHG6YNYzdanF9skh0e4h4jW
4xhd4Job3JLqeRLrTDCu+ULddQARTpeBJ32ZtRj6DhN1mFKLXAVtFnlZM91mgtuPyK+KeabcthU0
p/JpfO4qRrQWf6uxDG7OxlOK0ahPo+fGSaDoHZYwEQsyadCa0mIdlt14dAgWpWl497M3cG9O8Z8K
dn4lxOLegMl3d5zFoiNdlDa/Gk+ucm6KiHLdsGJwETIU4i+ZmyY2XL8d9HrwzRaW/FQqoZuiRIk6
mhWuz1rL7wiupto9hi1Lttk8qhTFkX87xZTvISLrGVD7hQGtauE1lSAP8b1Iabs46SKPWSEm8uSD
Bf9FLe6jCIQwMxWa00XoesJJFd0cKFKJQEDlGb4rAv1hEiopwkT24/W8NmMmw90RGUsowWUHNpCc
0XY4UdnGyjvBbg6GUX2L1+XIJeg+vsSKqjcImSeNqxrXW131ZFLBe23QaiSmopYnorNHRWMebYbm
wHl59A95EGOfmyVlZFhNz9jDyxep8osAQHWVl8cGGS0wa1FTewDzaJE27QOvGFJcKc08aF94NWGW
Bm4CiqsiSv6+lqXlKaPC59lRKLcPQ/O3iVKHu24lLpmt6LPwPHcc70o/VVppr7458TTevs/qu8sh
na2vonjtGMeATFOo6yvYtKIyrlXeirGFcXdRcym81jDMxnwuR270e36rir29hLt0Ok3y+oEQGcxc
d/UCsDua2zWDW0CHhDqScfPa90tlmzOMhyFwTR5pVXjOviDMACwndh23apVdjiWqUIcYeCg1HYty
x450VZ+s9JtRwyxO3fZ3xk7BANKFVP+/YEZx/EdY6+OyWJz7Z5I1+g7IU2dg+1Wg5xrd6/Gjw/AQ
33OCEdS1tdZ0eQImT3lUU+uFmSLV87OBziw7JqVwWMao8ctewnyE+QKxFwihiiZIqrm6r017MpFz
283VHgrmPdbdnrest9DtV/3noJXkad91gDmDdSqMqgFPFpqQF1hjLDiM+jPkZDziENbj1VNRkRaW
gkq8+NnzM+YzPfMnnRAf+E7US9YA1PcaajK+ZaKjsHrTYgBvT0/RJXlfYDdF6+7eH8PzneVdzl7L
rExxVzQy5rxEPJkShlDtXOux8xHxPz8X2NNSAJB4OqFodDryWMFnhro9p3+yEefsHA1Guvq7UhEo
ZnskZcBBb/ZV1xXGP8co6S8EKTUY82i/GeCGmhrJaIMgzMRxqQEI2w15xSgxPrZ/QMbHow8XB0/O
STDG9UxfrCdiUXED9FT7r5vN+uthJRwRcvp+w0xJ+fjhCiYO/1dQmDBsG85T1qbZ9IlIhChl0G9M
iFOr9QSd/hUvzXQ9JEHwRXity8nRITpbVga50Tkj9ZGmk+tyFcyKC0qfF+NvzSzgfTfJcAZQpKy6
HhfutENnsZs3fE/ZCeCgZZWZUPUXffFLbWksk6WUQ+dDjXt3TmIz7/rad6gYZC7UPWXXx5puIm2C
yrjvHQvESjidqtBk6lhGfQPFf/OxFdLfxihKWsTsd54PCEnoLFS92T1jHeTJ3ebl/TQao97BG/KX
qSqsPR2X20EreKuAow3S2frSN+WGQG0zDN4HTj4oey4piWqVMjEJvGdTAEJhpwEMchFS7VVychKj
3AsEWIS3OXkZ4IRo+1dvuLUzofME4UzRnXECz0nqiVafXASg1i/ofRYh2r0qGynEmb4UguPxSyXo
2B3lIQ0v8LS1TwHz6PyI2zKHEPrRFXwLXRRSNr5rZkiK48wXYXXhal8HeWBN7VbOdFwycTPnHEtx
4DqeEdcUTDYyQ7yGLul+d5U39hsYKMmKAI16e0U9wp2dPucekpoSGShBcw7rxfcaTUsnjDiLFM1I
nOMYBezi+BJKoXmS5xbWRNImuYcfOS5qrKcFm+hsC2aM3/obROp8qNr25nQC/aFi6kvn+5jnldus
9QZ6AVCoI7kikVy9et14yd2/wtfVJqe8b20Xuu51sahXKHWu3VzSkm+yeS33A7jvQKkHTHf3Q0iu
KmnWrqbS2ZIXcwODhVu8LBDjFdcD+aiGjCC/mK1i7UMppwH0aJkVu4h1QYe0PjA9sLFM4aG/eUsA
8irtsdCvzPCNN4SZzNW+K/6kO7jbI9FcTYsc4mRqZJHsjik0Iu0tiaOXLawyJ/PpvJ0lRU5bgZyd
2N71lv7xvtNulnNKUkSbBK1+X4Em/kfp1N2mMU+XJ5x1eGTzPto9JfjdO51W3WJKrvNLTUPKKPFJ
Vh5SxGGx5LrR4qWR1/YDcCFzqDoR6ELG9di/rK4JwS0zZ/UlNahxYdhQaN1BzA3iIyIjG5SBo/l1
82priv/fr/5cgv32LSzHVajY6iEBy8WYFmYqB8NEiw3BgWe72fzBO5S9G2vDJHnBoQEUPWz1w3xh
GmvxitHRru8jjx8hEpgb4W9XoIGIE5vyhzB2WoOMVXFFcNX/Q5dhtO7qAmNpU4M8O7ydl0bfdmVY
SA3wKL5W8yF4CYcTpplG/y87O2WYmPpkwugnvWAsQKx9dYIesaYaUN0kMyJGDPQe/skXmUCVF+hs
ajZ2Ee/anO+xF/b4PicBgHgsoW5iHAq0YRuc5E9qSW2IeB/1iBibNllOQG+2KtQs1E5LWFIunJXE
+c2g37elmQbXSuHCcctEe3jCYaPEnVycI4zJaRbCwZxBVQZePqxeUqR8z7O9K61bxXNOyo/7/PYa
2QFj9kEdrInoFNaKSyasDxPf2bPh2Q4TEJNchkWzJ7yduuk7YQzZbHgyN94xBxKKIN7DH0EJhFSt
5xrmYG8ZLTH3G00NgN8dcrN4ER9Bqi9tspAULbePoZMM++IKrhNGb2uo3vqCD0satFxMzz4h4S1S
7krTr+52kXwzUKum2/ga5haVEJbNP/fWfMu9xP0xx94QQJerNUaYDggI1CvJO/XiFPRk8Ibt7yok
AM4mubGM2uCYe9KhbJ/nTyQgXcCW9LAIJ1428QXTkZevNTQSyE5NynCn9ldkh1ah/u4o7FmSCOgs
GbOKOaKkMFK5ozpA10GVyJJnLpen9koehHmhlbKSN1+nOP2aBCp8VCdiGWkrZYT/0izrlblMfZAD
5v5ZTDI9j5NwAQsyRyOr3HG2NFCBgzPF7urwovGZKaMwbSyyJ2hffYVYHv5keVY+Z8EKtfJ8tJfx
f5G0x97yHyn2nIYnwhG9+7TuU/Wu9lD/QAGUbSw8Y4G/MWdYjYCngIYHgK5gB38S9tMR0SNUNAq+
gxy6CF1msQyx9ZjbS2baoFvVGkcPW3goKtcNkVXIhnXvlcekbNhxSxF69lYzr3b+KPIfIe2RwowE
vgT+w/dcHwl+9wZZeR8BeVZ/EiiiqT7Li818zkqDZGplkE+1JX1rtN0GyOqTLVaIuh1lB4rM0FV7
dW0l8kGSl8ZYitWtRj1l+XdQ9870vbyR3dctKnwSooBg09oqI9xluUQiSgYAZerdYxRPbXOd1bmw
vNmss4DALheJXrlxE+rryLvAnZb1L0PiRvtYWfK7LFzre3sHRnKVS7EqPY67jDoBNUITtPLsTbz2
ExhvmMdAsU5qCYbbTC06DuAdcZa1HEYF9tzFj1h/mRq2q1IHPnI4lffD7k4lwPSUjvfX8QB7PSn+
6CAQ9aS8Nfclc30EbIwsMhJu51vWQFVoeNTLaN/aUQaAZukIkuiyE5vVC3aYhSOHSUH/QcTGjJs7
GU8TO4eaEtK1JjgU67YGnO7wWFWc33xSysZFbwi7DmHp/GqsP7KOZlACPj+7dS+Urfx5SmHlwNXL
cQeFsw8ykq30FhJloqMTN+7PHWcK4bvJnm9jHBHW1SO1msLnZvwHDCladOKr1yJxHOdtSZJdjxnC
+D8J4a1CgbXcTpLrii17hWHeEdrOMCaOhpwsF8DNuiaIH/HRA8+mMHkWeLN62QbV2fi3ZmYkvRe7
kMuc/45V80mXSN+qAU0GB8KfQxWIJgp5puQQ+/Td0jbMNSJKAaEvOfYN4bjJBE998S2yjLGfIPQ7
bcXdyIZ+NuNKYUoDzYBG23BcN1N8X+3FK6UBYdFrptMogv2Dd4y5nO8gA16u21ZYfoJRXfh6pT75
zJxN2S2irqmcOqcoVc6T5WvvorVXr7Pwrx4eG0dWVOm31O0WmVIo5+e26XPnN9716+UYVdorEPN2
p7iWmoM/ConYcRHpkXjPe/35wF7f37mcUdZU6fSrAm4tLFMbLxcX+KLIpQZCRmXYfK+z0wP5qyMn
aYUZdvSX0jyNmtHWNxrP12ievzbegeyO3iETRglQPSS5pE7jDdVaAVUfM4UByWj/Bq6GM827wv5l
8totWFmApxi7wmJ2Dav6d34fqcoR2h2RnQ9F6jVqYzXbgaaD/qWzSYhAasd9xjjRvANUoI75sApH
Ael1Xwbxxd54eZdZ87xL0blxtMFjzqfgyVoiZosYss0cLu9X0ZkXG4nIDfL1tdLrPwm3MC/J6orc
qCCtDcBS21n1fK8I+oIR15I04MEvzuz97OVCHrH4tOtS4qsYOIwx1QmGxmFjaUXYuHHUvcqEI9TR
R+C+h31OllISV/WpnXsXSUzdk6Q8mNVP10B+N5T+BJfniA+LoTORVXFXL8ZBY+J/+iY5Q361dO2I
akR/XscaYHxm5c00zdaC0mSt4wOK3kX2/EjivxrKnR206b/OIjK9G7t442U0gJ+LEJSCi4nLyhUb
qoppsYBbjNSi+CFtC0WaEg6A0Q37V5mTCb9JWjhBnhyNnJd9m5qlMiKk58n26nd3Ucc1qzTnrK6T
W7BOOLRyQHa6gi0+w+z8BF7njyfcQUauOZ/OGSQOSz1RKzNOG9iiNmbqoL0/otXwQg8J5TWyM30g
2MVHb5EU9bFpSMAuz3gb8QPS6xo2hSEGA06lT6JdpueiZCliH7041LfXu//KFc41zAxXkv3k+dHI
t+4KIKGUHoe3/1uk9tUX3ACxgsGoIaly9dIiU8DZig8ygfB6Hgn3ZSyjSLIjJQujzLfQCh7N9N36
BjW8fiTRz1tcfeBlISqVEdnAeQVmoy+76JH5nyNhfgUJSsatYQX+lZWChoK8HN4rQNwLJBuCgG/f
NuT4TDrPo5GbsgYGwgWpVurEMGdsMeW/g5IBV/mbbqPwBdmpdpCEdM4BHmeUQiOXmSIPbiz9mHK0
qA1s87sxanlBgSf6SgfcIxO7SYV2PX6gNmPZb/E7cwT84g2lsjK91YsXwG6uT4jJ0zj9Q6z03gAS
nYavAhIPI0HfQg/msbxOftYgZrO+lwE/RnG6J/vZJ6w6kAY5BaWMUMDbXluwEn+n3KO0FcWH3PZl
YY4HgJdxlCd1b1ZFaX0XLGGaxBRI6erm54Ngu4ib+og6oo7udCyswztyCBsMdxxWV4oHY/vo7HgA
YyGcXnpREJycdBmvrq0gVHXcxtroha/V2L0ldWSLgLhRj4HlO4CNvQ1RYbucpR+V2TivMmKF6GRL
8C89/Xr44Y4VCbhhipbFRIcwou4fNBbiu0BhG7RriVu0qNXxdupRFvSc23z+M/T/ds83hJfOg7Zb
F2DY07K2teOHPDpuAIj7HILYzzexWi+S67zKx70Y5zsZbaBEOILxkWrJXWz6zWN9NnMt902FCHrP
dgFFLR/zSxRJuLvOWwLE2UuxLKGSN5Rt8JPurfGz1bLcprZsCy4XLZPrKbUKija82Vj9NZVSVHG+
gyUUSnNUXa4xxz6rrtW8pHJYjqauBtoVUFCKEDbFq/ugScpEwG+gT+VvIUSknXZ4HeHVLRQVPOff
s50JvXQee2vhelft/QQD8puvt8TmZN/UpMiBNEiJr7TafzY9xOQEhLMaOC03+bfdduiwLPwN6lAq
WHup79HhERttaQuKcKctwgBsJ5CzpZuk0pLTT/C+n4a6YqukAB5j8uDAlXMvk7piJToDEBacjPAC
vJwhCRI+GCp4ZFCiV/OqC09fRW2H58aZi7lTJ9fP6eiXtf484+8VIB971bK3eISvtbSLHt8GbaKx
M2/ZhLceewIgdhvm4+l1EoGoVvPdJ54bYtrdYMbViC5/bLf2679aCRNA3PtaNHoNe0wV6zQGQBnI
j/Qrd/rWgznLaMfrvVNwTrSr+KcHfqYGyZI/cS6+JgFHALXQC7SusEJed0QtmvzOWfQKuKHRXEN1
3XjQc4bQ/VZlkOs+wkKxzfE5A3lUX3NVaZaOkx1yjMLZg/eqNj0DpDgFimyhX0VLinI+UuxE1Lqs
SK0WYWQeEW9L7nedbWrhupZQ8Iogdqxy4xXtRMAeP+3Hgh/X/deZbd+0uk/qpBU+UYOaeob3TV3x
k4T9gDl72NgU9XnGQfOOMdYjDNBJ75Q8jMy/lDWG9OusA/S3UgRhUaXyxsRDLR/HwQJsOJrC6FH0
MCCSh2VCoNQRrPDCRAFVDWyLFE2RofhnaByu8t0hws6NJQoUER8BZfqUDIZO927B+r5Q8JM75jUA
cBr3d67CPAvo+sXKPyNSI402AqbYZCWNoJNhVx/wKV3pJk3fwLJSgpgeagoaZ1KiYvxG5ye+jUrg
YfJY3YBxLQK/BI/ueE6Ojzk7gLQVpgH2GOp3dCvbtSyzlFzGhkBlcWELJGl2yJlXXAWCsr4xEFW6
zvf2YlEmIHxoN0bpwl2WnnnZYPaRhSAJBlYiCkq+emi7I94LrtrWyXgeyaoVS+Gy2MSEMSS/b+xO
G17EoNo14xBvpV1PjaBXnt49IZwpe1WffYjIYRsdrUrhiDhucFnylXDe8TFN6USbBE/igQYNXs34
7YeuWASfZBe43SfM1zV8qSITR+xYrM72u45/IB3Jtc6c2QY1nWDflwBrvQpqZzJgU2iZdOwWTkM9
D7EWWHIwK5ORIS63cUMn80GxYGQeD72wDYrsn/DFJLVOjjpN3vTZNV/pNq9vIATdiLiB+mQMHqSC
4elapoyR+J6wozMFSNujTWtl/GWGIF5laeqSpPUpMRLoJqRFdlOT+2ZmR6UuGKhLtwbTaMrvKU0V
ttdCUWE7/ceaiWdPcnl+8dG+6Ts1ZOtLck4gSLWg24WmFNHfWX1T+dhpdXx1yLRko69RkX3U8y5r
iqoTwtm4X/LJvfa3fKwmdXPErk9uaxLLFMvr5ecwldUZ/uZ3xYEAiCrqnW20YckshVZl/10H7zVQ
VgQMafqbj7pE/zCoTyHThP8b7nQWP12Byl/VLbUIdEeLUxQPS0L8ewcybKkTdf9izZDRxhn5k0gg
yUzathvXhIOoJpKFALes/vSMe6Cq9zmQrkQBrZYMwLbjtq7HzF79gAhAO9fS+/XTg+9blWRTzmKN
3IdecMSbAJ3+1p+FE1o3D1WdeehcUhIotxcmWKCqT03XBDzzfBwvc6iA2brsXZjHuJ5XznfV2cC6
PzNApz7QfCrOfhwkw73vIdPvbFJ/XGi9NMrevbZ985K64S1kFNiUk29TA8zmKPM7L5Qo71H2eqUf
8y7aSZAC2rsU7TyvjOzvw9JM7H0v0e48BtK/4wbkl0ay/vvOXLgB7V/XzT+cRIh6NWmDZeh4BcXD
peQG+QN2AzIrhgehpXuoHgT7f3GevYCKYspid7MiyuZfRm6aLutifKysAJpDW+V5tNyLkQDh5wpr
sYUjRWC021Ty6tKZzHd1EXCWMuF1U1XwNIOfCIV3ZsxDcukMYmKJihavXOA+FHoQKCegBqvQwHXN
/Do9kd9f7wZY0cYU5c3dhFE/0Lj1FK4ak93U0y8EEnAJaj1Nnt65nP6gPssU6azlXfhMeeU9zDdx
am7vIxtryCpJGivBw8TbexkB1LoaEDkghPZgCkt2z//fIwSBPrsMmF8sfpbV/UzyF/4gTF6WrQS2
zjMrrLqCShKNHHsHZdD832f4isgd/wb7Ozgy7uJnRYyk5FnaU+d+RHn31/Y7po+CjBA3p61GzcAq
MTVf1QR3tRFok5hZPg4Z1A+LiMvZqY3iQQ7cCDP4bbZgNIvKee/jz3qVZFgytQBCgoV64CrvQs+b
HI52H4l1sgeDV2GkOmWVgG7jDhbt5MPkmf8982gzOIhmxH/kIx7I6ZVAZGOcWoSJoadJMbqzY3/S
/UAqyABgeikcwgU4fd9JVDC9O7E1bQ2WfIMEc15Ht3IohYUrAQtE12T/j/svOjeVBliiZSeayo2M
aD0DSMh67Nm4axqhtoAyHaZirWk/ChpYivJtm8cpyecKrM8So/zdtc3PW10XQ8uV1jWfMdRQZrFL
eADEGzbcutASd/TIxx+JFK5pUhR33NdbAVabn5IV+HVuvBN6bZF8slDmpAlLdCYSJyJjmn2UuThC
I4YHHdazxO8C3XXcN9/Ntxve95ExvWk3Z/Nltocs5Kx5ZrfmBmAjtlWw9hSGfj8JSpS7kGjQV77c
MCswB3cALCZQV0nNeS3eW9Gio6LAn/dVs9FIiF4TqI0uljkidr4pjI1Bl6ecTCJcRYmsRumrQc/0
dkG4+nxq96yhC3yvl0WnHPNWZI2odrx+78rUnNSRnTeCEMwT/sDxDrJnKXIC0lqVIFojIPfj6CwN
81zHqmapHLxeRv68LHHGRe18SipTdhq0qxL90rX3oNNEbnEaOJIQ7rQrzftIf6AFrpmJRMbXpR9v
ivLbZ27qcxvLZ3N33NrCsAODk5mbtQ2yYhd43hCF+9SQmHkzzqzXOW0kzPRSZrX3OAlILO/GO5vW
139crNVil8trvSVlYayPtOS8J5+OEWQM8NhFR925/36VO72mOFPHEAAWw9FxWEzwV16P/ihLybmF
Od4VJFbiEOKENzb28h7VLunRy6ZDbPReDaftzMCQO6t/iP5PQ5lOiFvmZS1Vyhpm9ySf8gfgEQHt
jukN+/d6FKcuUsKKulpvt9aRvPVdF/8mH3ay5S0fuYCIAR/nIpEHxXe11FDArhxSnLV5Z2edQJ9T
Q26rcnVbRIibNpKrknASedVdMMikw81DWaweQQMfVVObGVV9rHTLeBo3D5FzWyKmODYmYILC8eoI
DlJhphM9xLQGI6w2AYXf/d+Clq2cNyBX6R/nTXmQt69xusfFpXUpmBPvsZcwVSFSS60/FNnvT/5w
OQ9XzKdUZcLUOCJ1eXH+/ZbGr6b4popljRRLf77Xcwi2kMXmcqfnYtucazCB1GRJMVsKCsVoebkv
yATgxZ5dUlJmxmqPTrPnCkwbO8UlkEQImjWDzErud+abN7R6+JCuutJykaMM2hB0EMZL6TZHEtvC
Vdz5y/CNA9Nsjp7QF9BwjaxCKMd87wuQbYlqi6bXVOPQfeuPxpN2NY6egLX4mvbXqwKWJpYWTeZF
U+PSDtBW8um1ulTw1iv1pWmGCoV3oqKc94szhY4EkvTXqi8El6m6gQ/FDQHKq9TtZcpKQP0pVZbW
gRr1xkCBZGBaMamQ8EkOFZp0M6HLcXSY7Oav+VAkNVoShPTXdaPKl8vZL5FZgLLS4H6GLr3MZvxe
k1yE390vM8a5O8HWe9S79TWx81im76xWLZN69yCS5maXiFxdO17xtWb/nXEITTUF5K8nLahvP9Kw
pBWbmZy1jMCcOATQ8MKUO0ecqPU3e+FDsiGUIwKZtsdsvobjRDLVfZPq0WgaZlQ6IyWcn41+mUvZ
PTGj538hKhNX7TtiJkZOjsu2NE7n/0d3iwS6c+wlwa/acE5A8wopavNp8e6To2zUYlB1UGiAgU+Z
xPqZpVEItcvcQJ/40u+z5azqNbp44GcudMoLHTiHVCx5lBmwi4Hw0JUP6xlwdxlHWhp+eMapXtP1
ahA+4R/CGtaG0UtbiDeXlU20XChgSUcrC22DWDlKAdOZzXxj5P2evJLWaAvIbcaj4JRSgD6jOe0V
wCgqp/XkJBqoWJ95Rzz1x9USKDfKZ8pATAwbvfFMYFGhIt3exbgx5ftu9pWwj3zanrwbHSvArtdF
d9Zh4vNk2xKfkJPROBCpy5mOsvPwOc/LWOtQwxdrUJPOFWQunuZBl7zCdPb6H7BvWEM5c7TJKtFe
n/pMnef50ZQdyFlyNmZorVxcCEZSnbT9EHP9v4QuBiw3TowKB+FPZfJHA7J+5fSUVPFEhclUCS8l
bL/Vx04Foixe2G4KbRgLe8i0C8pSnn+o9256fOmv+Ivn/iISF5GlkM48WgflUVuRavct0/df/NA2
xmrYQbkRgsX2gEf/7cppFxekNDPckiQRiHtWg18Ju34m74N3mFRRHFD69f6E3IOlu5SdN7lJM2NY
VXTLYOSkXB1mz73ZJw4qlyYnTAk0DZKfDXPBJ8Zxd18klm0KsrQqOWHm2AX23rPLMBjKOdn2umBM
Q/gp9q3Pnefz+ghRdbN8vsyGuVcP0aHVY/1Adm9Wsp/lzp6v35UEQ3kvABzL9+hxIzwwwGcXYjYI
E7p+XOFyKGcNodEH8CvfklJluJYAAQoDzGEjp2QN/5vytuitNAgMgWJxaVAkW8M0vl+htqNmsJyY
ZIKqiZwzQgWCUPJh09Nyk+IN2oEbaEzGu6k60q1hgnrGOikXObk+CLjBLpNfvJCzvtZrEcZPyGHE
HT0hDyEqWxdCNxK4S6FSIjE3vrxv9n24+rEGPXq9PnlPEurNQjz3Qvn3xwXNS7K5IM8edNhTF6Vk
DhzV5xeXd4vgRJVZZl/7hKty0MTmZrw80Z13vwmgwDHYSNjjQC7oG2vkNjNNevz77QyGEfTVFSFM
YQCMb5ngBngdgykLJ647l2tLwejPPRKjqv/2+ptaBR8ASz3iM3fjIxV0cuqp99KNAXVBtBoLoBoV
zSNKQqCTNxXShbbc8L23hF2U3lg62O0kfPF48pb9VRFO+wIxCKbbcjloigFvGzMGbasrrIU3eqrr
2ieGY/xh6ZndtLTmS3ZV7HDyZidndYr1X1YmvlI4l/KsMB0A4b6rl1pkUBgT2fuswTBRmUKEoNz0
cGefyNOb64fgjuj/Sidj/bv16qL/LaY89r+t09PYer9HVZdxuL11xeQFxOnuSvVg7RVmKwcyxvLM
TY8t4/ETM3k5qgEMidGxi/CR3lLxOBf2J4lL+97OzupwimR1DF3aonJYpfrNdKBx4/k79Mwo9W9Q
+yIO/mPWui0w5rDFF/lFM/iLTyv0JHXKFAJzt1iCNlpndRNbH1EWHj15gN8JB3vOZ9k1a8+uEV4Z
mi0maL9qpvY282CL4oI6+j0EIlDUhLxScR2nDG9QiD2rMHBkW0oz1yLAcif7c6HlWTuotaCDxG+c
FAIMNvVDgHX0EOkqci7UV/qJjzsEx9Jq3PdG9fs2RUHYJ2i5pLF6Q0GzWmJDtKIyGjvKzLqvVJRo
myCYdBZkqig1ZVpwxfYYWwGuWqGKxyIu6TK0eumurepflQvgl6a5A7XAtv5gT4ESYMVNFp5U65oy
yvrgXWcudquyP8dmgnc4U/p3wlPwKZiWNcmYsGrGihaXjA5CUpGhL+tK8y9o7dboa5RffPR2dOdg
gReGTklMpI5UPm1vskd8dMwyPXsFj4keR8cxYcY6AV7qODhX8dATtiPoLIrBdWQo66MkYGOKnywI
3yg5liSAyY6ba/0i+OkHn4tkYzgumsPCzpAlTuX9U4jCaUE2+sCTLsYzji36BDoOh+0qu7PbbL9Z
tGMUD29i/iSLE2s6s+iEnyHOahg0UUAqg2LvtlS2SoOdafTUGWmD/hEwU61BIoSAEmCeI7ZBaKvf
25mq7ulDrGR8dA97ipTAyS1dZyJjjWLXAOAoXGF25VhvfAE0qzl2e1mpg5z8z8UdL+aQHOPxnESl
+kWh6tTbj/CcN99HqINuA2iopMAgylCGIUaxhHszP9HUcYTdbBvWrT51FiBrI/lv1WgsPR9oyJhq
EYjWmrm2o9K9LUlsILREZLuvovEmNzm4z3/LHUePATNr9/FfV+GSOb2laEqe2S25SrVjUOVh3WbF
0BSjJFCDz0rgi395P5Zmj/eQ9HvdSiYJ9w5fBEM6ztXJrPZSmcLg0NIvx2+Pq3mdUHRYjaKGmYn2
/+lriyhJpSMgdKD09scIVVzQiJvGi7a2WURPdynQbZTUzN5hIGDoZBwhEyOyb1eGD1BLuDpu8GIL
LoBBBD26PuohR+dHRRmdd/Xm8EpkTuh6wh6DBKcVMHBinSFOLOTC93Ak9MHzSOaxbEfpQpaspedD
xJYjTHZz7lZXM4ZQJUd8Jv+LxB5h9B8CIH+rrezo7OIkknbVdKhMXwqIuA/Flu/c0tND6TA899sv
xzNpln85ZFaHCpFJcWPXYdhTCcqz2ldy4ImUmBxIlqXuHgJKk5zAHo9fdAEsOhfWxcKbBFVrjVQO
CyFWsKhC5vs+iDN4Q90fAKgWlI8SbeFsVk3F7My0vu3+Kuvj3zMKLwOtIW7eLzUpcV7wZp7C0zcb
5Tj2CpR77Ff5Cq7U/oPh1mKNDHtm+xiyfB1fv5+Ul3OUNsbpZeJtDtfPKonvt7AGqPk5z8OqYP6w
/lQawgZ/p9Ynz7oUbqOwDhoOe6dfDAZGqRnTP4tZa9d3/EOhowNZaGuIswp3GlK6UovCf03y/FVn
y4pC/uUm66533iJfu/2X0gOEWTl2P/PqhdUcrcgJ1TnJH3nr7ooKAUY5j3VjJVY9SynvvOwljbC1
BABMOBpnsGegB/llNNb2Hs+VJr3YB3ijI7p3oCyzwsgpGaaxXVeCruwohanQXC2Od9BZpdG+ECdI
d+c0r8LG5SpZTg1Li0koIq0ncHJ7XMEemeUfkaqZhzOpOICIeNB0AxGdhBi01a4SIEXDuSsl5jjm
bonfcBlA425u8U1wAJptjEbkRxaemBxEkoHtYquzWkTF9IB09msmEm985/fPJVHqEs5wYthLB9p9
YGfR5QayZzoDGewWdnlVuVjM6s7d2ZQtsBd3pmK8qe+Q/1RzFqTamfQ65d23/bIrL5wGFWD/Tske
eQjSqy02Y6wVm8zXnSfGfw8xdEyaRiNmVkvxCdbECnL2K3vqpFLIbI4/zpoYCBrGFVnEFF7CB9fS
vgXl5uKViju4hrs8ttH2lnCxX/RY30vpDMbM7I810Od04rgQoaaXwbMDD2fCrEib3bt3g+1+mxCB
FzoHeSX6fDhNXf3SyPjiHoNWU6lTVUFkgn8BkwURxs+CXEeUGCA/lQ24f1ZRuaxApZjbqoIaQDBl
Yj6amSV/mzzyOMidV1zbPCotpBhnZKgFRidxHlojxTYQXEogPHhXhIcen/oBQk9o9sdxXrM7jloj
f7GcqBNd2QluLDOSeUR7PSvoB6qLkwwtKVVX6dzoc2nnImVq63r/frboo1Nzg0ch57Gxd66dOls2
ZHW5jD7evZ0VahZfok4MhoZ470VrpOT5wmYL+vak58pAAq6bzDMOVrutRmDitQFebiEKmujet9pB
vlysPFQ7BeGclg2aC8mSAOAx9C7ZoniF8BgshULI1JJ7yR7JrxyHYclI9sg1ZQKX0iS4Wzs1MDHb
ZrubyJ1HhLOMiC21dDv8iL1cYgK9gnX8hK5j6vFTAwKi/NQt2E9MvsoLS29/GdlV6KeIo9khIBWR
c6oWNSh6ae20X0R9BVc853a2Y1pXWzVXfkbouJbqOrLHQIZH//3TpR4Bs0YUnBq6Qh0RRidQIUwR
YTSratmrYIk5/jUq01EHg8X42rhntNRQ7De9vgw7pwCHv6p+ZA1o3OAiYI1/UdUpteUtrOeahQ5e
PpfZ548bkrcjrpeFTpK0r4Z8KNecuOcdNIgh85VyW0ptIr5h2Jh23M3VDMOaBdGr6+7V8vByF7Md
cZWFbY4Yd3JUockbo5hP0E1idECyvv5cSkHYEAse/ozMgxpuvZ6GbHx8FqLsnFYcBK/H+IMVWHyK
X2+T71S1SWiAqaYAhFduY6zDclaeEzHjHkwzHl6djgp9MpYRuMoeOwLanV0te5D7/hkjy36Hs/Oa
pP7wwBphZTV4n3MA8UiPtyvOFjdPFin2gf+Q+tKBrHTRwo+nZwCbA5iC5R2WhTcw9szzcNK8SWF2
fZbnda0eGJDcddsp8sgeIbA3jeOe3GEkSYsoqM20j+NDQtQC17aCWd3LQRGlHAeb+ab/P2GmjMHV
W5ZXwd1bamUTOARVEe9DmnFUFbiBb59GoaFD8VMDSSFB6I3yPTV4uWoRlZgEXI0a2QaunGTVKEZy
5uiVtE3fDTQTmiptwJyEjzasTP4sNn5w2p91TQLkSmbSljCA1jkqKrAZPVcTvEYRvO/5x4lTN7CT
E9k35b7LuSbm6bLqyjRAIiLTdEV4Y91FJkbchCC24VpDfZEkTthlXYjCH2dpPP4K38bZlHpzgQos
4fBmEMaWNPGlphOIIXBWqfZqDnhxZFNnGcukJCSZihas8f4BCby4BUCzsmlQivUSaz0f6PImFOxM
v5CDZLjKjQzsnprAO3gerEmNSrUBjN6dGUhf9Fi2lruvONrx/2UJnsIq3oOP74noftMz1VHU5U9D
SE6wCSLis5+VqvlnwShOi0UlGywW1Onax5ZJ3acbmHdj7RaZt0WfG95pjKGki9USafcCMc744s+h
Y6DAbogsiWC0LBh+wHQ3J6n/M3sQp8JhXnWWXiWe0J3/7H+qm1G4sMDPotYHIoqHReBP9ipfhoPf
C8Qb9x7qC5pYFWqrvOts06QKV5vpfhIsCeAvqicUmr2PyLHfooI0zi9Wk5P5GKK97hJPhb/xVZEY
WgaGi2TCs3rq+RWBaAdF8FJBRvksGa/apFhuBpUDYWfwRjJfwTfw2X8ufFfOuklNY0NLFh2QJ2KR
SdLKD/odVMVikcz6hovJyzQZvekxJAc4D4ZhhV9twY9yhVNIiOux6DkXK9M+15hNRrBv6FoKPyj+
lWGNGS2lhS3iAwZmGMX/e+PVvmBSB5UgnrxonUI7LyRmtPupEizrGj7WRf+TKuRw5D+mvzEjZlF3
16XbLljFxMzNsdnxqgLs6ETaqSORwOeMswRxb5NLWufVjIdDKm8ze3gfBtRRCgG07r9aD1PC9Dl3
iS5tCeRVZmJosdFJxghF/GDLYmfbvNF2pgsUCIAZIL5ij27agYNwOWygKuW0FDAVREqu1x+ikBS9
5NjArd2GEQrCadesGea9M1rdsg93rTj+7J6781oCZxWqyYchRRcN2f+l/JAfvBQkS0s0GYeN7rog
+ctoY7jD5SXvj8Chd5MNmD31tjIcSygFoiexYKiqCRZd1JvNaBskalwqOVO0tnT4mSsxNM514YPD
nAo3rDuiSPSe1clk0bWokoOCCQpK/CNR7dAWRV2r6AGbWhGWw6VvRYTPVLmcZaEL7bBa7CiHnyvj
il22Y/plwTXc8Dl0mCXF2Y1nY7Gzi82i1PvtwqKaB+Pk0RuY4iDO3U5ERk5biW8ucSx1NRUOLRyj
niyK67SHYWhWqNtUS/YrgJcWY1u1we0l0De8mWw6EgL2I4h7nmFI6fzcBcnT07qnvg9VyqY4353s
WLcMZ8SR+xqME5g7VUexmhtSqNdU1TBV+ztxRtLq+XVMEoEhSbXekNXywwq6Z5TXA9UoHZ4/7lNu
kR0pgQegDspEMyUrBZXM+SPZs9thRR8FscZ1njjx0p1TD2YT9ftbqZgGpemodbIu8VAj6FLC/SCd
DLBZa9xKSycRkwqTXEwuUPqVi30UfeH7XYpQCgADfMGBpxjTSmruyHona9OsxgIAA16ofMdIVBPp
ujjDj2F/qWXQUWzokqo+ZChQcpNf12+iXUQQgi1wlDhOIY2uPfsFClGwUU0LtjwiG1uKx1vQ46pC
IRpRKI4cvg+ojaHsUUVDBidqhWEmqOa6xtVSZ1YQBz+qikNcpbzeulgjTlsDwdKJ9F7pfffSX83w
b58YydR2ndS6aLsaQ+9zdjg1WpTcVzEkN7Gr1CL6ndQAgwIS5TfyD/DDgxtzy/YZvJXMG+jZ/CbL
1xSOWpRw0AXzPU1dIz2xcGk86zPCVLsSZoGAROBGqLX3jKn/yNGAfGFiiY8XSivct9WGwvO9cws1
MYjcwK8ANTOgj/l9qeh57sMXDafAnT0abG5//XkWoeqwC/fZd/cZSed3NNsGxIHT0Sh3AIRAnmEx
np0AJMfn8nZHq1YTTRUooD0hq4gF+DGFNgeUyyfft1c3rip2AnmZvJys4vRtCOHww6bVJ8CYC4pQ
i4hXKGAr6WDJtgZWRWLOzdJ7ejFb+RbigKUBGku7ZuJo1Rer8t/p2d2kW+Jx8+BtIfHFDYgixRB3
zC6Ofr+AWJYBYvzFWdj884/a4nDE4Vil2DUdUsLPfW+v/Vh92Na2e1ub2i1Vh9VLByrtcbWLy1dw
MpvNNQo26qW2ME5b6QVcQ/ENLlL1Djsf+59PHLokqPMnx34wKf9jQdh3kvd5S0MUtjR7q4KT8rTJ
iXTTAFxkXTjcO3SJNagdXOQjgIpbCmBFEO8se6QGZoER4+L26g5yscc8UaUo3aKz/gsc5wRsSIIF
dKklivQ5aTxOH4Q/OI3K5PIFtUwZqhib5o2/9RqR9an1sd4MKPHCzk4/86fbELblE8ugImk69A4s
cR2T1KTGHtx6f8PN48Q1pKKIdQhOo/4PuG2RZu2z/fGmh1nm8jC/O0qA1uPnWN9T8bpTlQ2Dw8vc
tFQmFNabUtGdghhCO/aoADi2Eff0aZobh0pPZSf2ZjV6dNXjvs9PzL8qtMpoScAiC35M3dPJH96e
doI4Sl8Vd2qQ34GJK9UYCRj2/0HhJi8wbZ9ekYKlCJ7E5qE1zxuO8dQ9QnJPB64TKeCscL+/Fyr1
MMtJuoDrLnswhMA+VaU9pJspgCa17UOwHq4MbqJwNS0vhDPd12FGDdXzD5PlzOSmgErb4VYNireK
5AywcOiQSh+Vv4CNYR04VpDQXOOMHzv4dLKeQJtdytzSOX1+nuoS5OsTVbaFLdqMW6uLVxq3aUZY
mDuHOHVHNV5pTLR7q9FRS4crBB/WkfIfdEJdygfDdeeQLbwsqFOqLQsEJT77Ml6rI23s8DMLmMp9
b0Hkii8iLh7EqBUSI/GC5c0g+Axim8lVya83X/To4HA/6oFwf/PDTC10qMDdJpL+m+/V4KBcAng4
K9UB1ReLynb35Fmgp0uwkMUFau8hsy0H/wiSXLhiztdQWBb4bdHg5UzJ4cZzFJ7NzzBSg0OCp3zc
lvMLwBSO7crs/pHZryt2nfCLBvwBN8wIieMmaPBbQmJi0pykM3W6v6N6f2beTEBr1Ij6E+D82K0W
M7dbzeG0X8TS3G5VJ0VWkwV2SKmX83GrbteuqAP7SxqxkmGXvzJQcA7lEN6OJMp9tKroIAdodjm9
A2h99pG9k7EknLt21R8O2FtGrZA7802I8T/GAdkB9hGGThigFKNO03yrhgy628PvWHHuLmXv0pTU
+YH7bOUHRhoda0lYtRyWHjbj4hK0BgmAlkTVmEx72Cx24Bo2hTwv5vkQ2tCrgmNrpZM1kC2pCkgA
5UDuPph3HpzurXOA5LkZXZO99WlsepLuKhMZ7xw1cVYZwOdPzL8Qs6Yn/fzO02B9PAY3gKEnclZZ
NxkylOGI2um9bBgBW0bqcl6be+FDFZmnEdpLSD/iHAqnqNcYxHm6RYEFEhIQiT98E8zi+C4smNr0
OIro0i4dQmp0Mio+gn6SApiCI6W34r4HC9PIK3GYiXN8uUM/bNhW7KR6NkQPtroa9D2jWV8vV5P9
09uC4bDa/Kn4Oi9IGCSZ07jdR+KpUTlhhJvcSDxkeCBafJb4GA+za7admSPWVJ2e7hB3ion7UoN5
3JHPyKdXHlrqGRUd4qNTeKBMueCDuhnGWe8XEvWn6kUYxmO2dfZHyRCALf/N7NXT9GUM5+yZ88Q6
jB0Z1BmyseXpkD1d3jR9oyNdKuQFYT5+bRUym5lZs1C4PLjdVo13Rn02fEiVgZzf+fOhbMZTN1SK
hYHzBny1woxtoI7pf8ln/5JzsZuDV0I/KE9o/p36rgKxmKiegHNPePCxv9Hsin2HL/4hysmS2kYL
2PXLBFiiDg8za9y4IU/slQ4kv3q2sCtVszHuEAAjpL+6NUctmRhZ7SNFYaV1h0NeEP6OACyX6FuF
0BPkN1ytzoJpEZjKxA17+iJ8cJ24AV4vwu4QV9kl9Xqo8Ez8JlDG1F/sZBwJsn7/mGQMirryh74a
3fh/Uo1v/c5GQ8N8GnU32h7Y2f3yaChGmpfgqKR9riT3hs2r6ykIsPDd7EEnFwOr5XMTTKSZnk9R
cZzPCbGs6Hf87pTmPs3cjFTP1C0YxBCvFEc3coYVKfVW34jfdu40RwXXQEzYKaiSJ+m8SYLciZLd
yYhHcXbZpUiQ3fCDjBpnu8mXNbS6rVD1KMoWGaCxYjfqFdvJbBPPxKVw8fLMz1DguUe062ZXkuIV
MycDEwRE0/7mWHfbIwQKfjWZQE9l2BIlC4P+ViV3wLoYgyNbOF6az0/M16/HBYT6hbkj0bs87Sou
/C4eL4/UQ+FIOdBf9AugGSAX2ECHh6/sNUyG+kKyhhtKxZnL3f/RoUnhe57TzgsX40ev0eSHAKaZ
VOtJM0xsM2iZvIXOn5YgIBVfqrQWDZN9eDxKau+rFYzxJi8dJkj7ZSPZh4HcCArVYNOQGPDzDsZE
4VRXL6T8CSeZhExVJAi8ndemsYLRCRZA8/c1XaogSB83FyykmaM9LsbFvhUP2Fp5yL6/VN3mhtfS
eWMb/jXYWhAZcSj0OEzFYDURPtReFeNZe4hTuE5iZ4eRq6o8x5r+FEvgEf38FrrvqnW+qtco2n0O
U0eZdflVf0tFaLnmadYqlq6TKDQGc5VPK8Zm5tGrHZZWZnSisdsEcGs+J2o/CDNszmXlj65qnQBn
wEmWkQ4ho2AoRVW42AxvcGlzz9SCD9I/4aZJqf5L2ybomYfRlp06HZUmYPsIF/6EW+M/XsS1Rhyc
sBPN2+XcOB40M57hkkkcdB+/q9hrbLXUJGXi/TzB2DKzPhJHV6IzMYd9BhIkxkYOxupwjBdJIesT
zQhHPWT8Q86vT2Ejd9vj4MaQUTyJQhe6GfgMRjLeNplpE0lUN14yOumZOyktzExn2C6FD5Tho7Uv
mHX5uSMAetZGDB5sZVCJgOSJx10ZvJd6lwUSyWbKuyG7nGaI+G4/Lqkcyc3F8PnBGbFsZi177jb+
uNbpAQjosDTd7A1kGmpSL8z4Ds9MXjFNuEh5wVoyf6U59Z8fjSAspgY3wMa/HNC6nUprYvn0WsJJ
I1Da0IuVZgJrmGV1fjE0tbR3bYE4RR1FnkGbuW5j8tQ18iijlS/O1ZAvASHqYUoxjudSEJfmLEv+
woVxQDjxdsiQYWwO3eVyyfs/FsVfiJvMgXzOVOk8d8qKq+Zj1lA+Mi+BU41fq4BBaBJYLGYeK8kn
BXjQXeC+E30IAY6c52zu+MbXDr9Yi6dUwR77VQIm1u+702flO/pYoVmZZd2bfx6UF0S1sJYexGhl
i4Inp2bylLfFkRQBeVcIoNgubpv3Bc6OfF/Qr3eHiF0dyK/nXOpTBroQIqCqEdMCgoa+/bqdOZ4D
uflnd+AVXfdhN67AWjce5I6wcnSJN7ZVuFXATc8X4qJ3uOiwsDBPBswyb+IM1k6tGCMR6PNzATMA
Wwt9xZwWLyyyZbIhRPgU1dtF9qwXwHjEd4fULfbyDfz9y8B5bDQ/0gd+WYxZtSEGTRmVFMT5eIjt
zNIg5wRvwwNFsl7ylrjwu/GcrseCWvbsmetwKqbRjyC4IGvNJ0jlQ+DX/O37RY/HsP/QwLFx0n+Y
Yz+wPHKKQdRMz5iEmUCglKfWCuKohGEc8i3bSmxB7L3lRVlDbzYBrPK99Rh9nb3zDq+Y5hH+XDjj
i8s7yYFHjd6wulvnPkCl56Mk924Ry6uXh5c3O5wtQshHAwr3q/7M8bLl2Liqor7QfGX1HcOIT+Gf
RjHbuPPiSUUd0f7LR9rsi2PjVC7uzgPeNUhC+86Mo2nzauW+qA3SOa4rTdX9yHFX4NSjgEBX4rXw
t2VktKmKzVzyKfx4m7XsMwHd4yPKQ1jZL3diqY/+LRQkHftAMSO9IxAmymdDpl+vlf7AVJUt71En
DCSrvlfFqcFcQm9OGy6aBSF2HSe06mTx3bawjZERKk3VSQCyur2RoJdxkTbieVnGgK1BCYnUsrEA
ESLTm4BPCMh48f1aqFoExzHVXnP+EnPmjMJM6ygonOPzjUHemn9fSeGsqqNwoxPmKzgbhkWUA0ta
p1tapQry+5+Wvzyqu742423ulYxu+Qd9FaTQMc6PfqxWBZ8f0Wt6TxGKcFd4376fZLXqnWA0jSrX
ilSYFdSjMRjjQv0ZjuYmhZ988Uf5/Qj6Ac9iK/7cZl4Cg1JdxVM6a6qq1T0AFzpAPOgjpW32VOYq
41uYWW/47qvJ+c9qXeecK6wSq1ZJWwx9D3vrb8AZNzqyI/jez04rZ8TAsVB/UeQUY/Zv51Dv1QdA
8cRKHDecqyyAQSL0W7DcbIJrRH9mqMqKNEgOSCR81nMfOSuzgiYl3tdIVTn+7LwzZPH3tdnawK7H
GzLucTccsx70+8CgyOtUPTA31zgR/b7cF1bDgwk77P9kXweqBCTCN2KGGLP5IlN7bPT8jnmVC2L5
G4NiHHz1rDxOIZpSgV7flsoDZ3aQpB8ZzbUPDiL+f8uOq0MJCqUX7HW+4+BXLuBfxIumOuC+A76f
hNIlHS4bB+vFmvHhnTpIqfVgeJ/S5sriJb05km77oWE4eqxpStP/WLualPqq1WpdoPPX5Z9N0v3+
tzjSCQv1CynIDOZxWCsEjoZ8S9IDhb/i+g6DYVaBzUULMhRSbSG5NENacGIPN7HQ1rlB9JWYGsDx
sk6MMjzNYkTUV6DUhqGECnOOW5aUfA/OcXNLH5QcFydOrWXnzgQg+bR6H78PdWrxQqoCQbfZdbkY
KfagqgqVDlSu3v4qODjT99Ob2Su3YwKxnXO9yIQlWys5oSFnRahHgDWbRff4m63FuI30m+Jy2Fy3
+pCkjbZ4BB2NBG3VLZnTWX6J0ZxWskQEyrMPFSNAzBmAH1OHm0UFDLofJW3jesB00XvNCTL2284+
qJLJ2yJcm53csYgCGbI5XxGCQyVwDMhEppepu+RCNAsH+CxWmkR3LPa6U/CKft0uSUBeoZ90Li67
XOrDOYfUwhMoiCEL1NI/Sv7t/ebZ+rfnBdXGioXeiGHiNebq3/dzly6Ym0ivQTWmnZ1PVMtT+KsX
VNfnxKNgMSQoSvqoNeuTzHims5DIxlVgMrK/w1uRpAPmRl44ISS2WrEOSyHGFIx+zBm0b+qCp0L/
TzmpmICnllfdJGdD7VaEN82BWAQbcveXUDsEKclzVtg7l+KPg3vKD8dpbc/eETwdyTqPHZxb+9BR
ZJS5haEKV9pwmFOIQFtMn0aHM6pHNkbrk0CN6nNDZ3J8EHWOdGTbNIWlm0NOlsOvReHYnhTqnLFK
GipUwfozszGS3dCLIzn+D1Rs4pWU2ivDhhqsPtRD5/FYdd4zsCZZdLB6173uFc1tRVjXzZNAHCzh
J/M3+XH3MThmpyziHLS/kvX/Kv0WLwdFHNvCy7mhQuaXK8wDcYMp/VtbynQEGk2LorGi8DxcnSH6
lxmhYcsDSupQ27t9J7QOUZ4koT/nz8685xkzbJ+SKExBCFe+gVI2ThpeGxcVBHK3/LLXsKzIx7ZQ
B/AieKG43HQBouLP/ZjKbV4YRegryVhUwoID7VLGVu47S3ScB9wbA0wl89PYDwqDEgTV9nubYM3c
2Hje+wY+IDI+iDQvAlRhUSgJghRhayaGscXL0M7je5mCjOWqPhogFVGKVKdBPa+wNCSJinLnJaRo
+scmghNpCMEQ1AZ8gXB6JjDOijbQNnXwgarPfoQszNYeUWDtWwi70THykqeBW6xL7fhGK09pau+9
3Y3tPrnXK4CUHwK0B/AkHCE84mFwF+4zEyGxU41dU7NvS8v6oD7AYWY0hCBt/WV+SrjEXl3whZuT
SvRjUOvoZGHZXISgpRbR65B4vGdGUqH2aqyWoYJiREBCE/8KGyct7oy+QycbzFDcUBvDny3EvCuU
4h+90bkrWm2bllbme13bXuKAmsHimQk7u80vdT/i3JSj6Q/Wdg5a+WkIs8c5Nl77r0wTb1FxCw6E
cEUXCulIG57HvxvGrrlga2fvkVdyc/bjsQajpLTdLv7M7q9TXP3xicRv7W8ZKB+MA97QykNuM80G
3FkICBvEfd0imX3hmLMXshX7IfLzuzBwJBJgfCfHoX7phGc+qRLGqoTlAQac7vbfliIeEP72u7+L
JeZsJym1Vu+KbCJcdxFC24IP9/Mh6H0CIhprKqpVSIrVmKYMX/noHUQj6oDp9tFxHYuFMY7Lmc6o
FfArqZKdvBl39QOZa7gHGFCjzfJSvnhWnDiOnzQ/CA2NtBvo8KzDLKOMK6tA+O1IrV8aR/Izd6A/
VCbR4EdERsugzO0xVnGIcFk/eOdJFDHOcKov/x3CsOwkZI7UrnAZCbIWRjyf9ftniOh7AWepYMR7
1nFLwHhbfesnzgfdp8A860dKduefLOEWNMe8Y8gPQman3swoKzi3385fiCcGlzVt3WV33PP5hE4r
CK4lqmbdpAMgtOEbA9f031td726E6nRMkgHKSjlB9HNJAl4n1VPRpADYQ4ARbg/bwopGsOjcSU/2
mDqoTqbAVC8YYrzEPhQuXhlQhfYm+fYADsTKd8wsXnwTuQ2seySzDfi+OAnmpeHS8iA19cXYJ+TR
o1W0m+aquim13uHUGlabSfRI9sp1LmDFu2d7thj241j9l1bYgnSu2pjd49XHSjTAJPaBJBiRGvL7
3dXg63GxOF97Vs4HroNx/sWsJ1HZFxCISqezDz1QIetiLmVSjOgm9x2hZHhcFg/q4DkdkoH8SnO4
huYoXeDNEmqArhTnqk11SmXYUkD1WUv05oD/F90RWkYwMsIQDwC/6NL/3At2uwLmXbczacun+oK1
GX2+Z+j4p7/UCVpMFsxb+jnqCUADYlhwnDuEfSLHucAseDeXy7YcHlrudZ1gi5LIszGdk6dM6SAr
vjJHoFjvu22rVXK5jYzzeOlVa9vEGEQUS7eNnGKPu5oMLv9FnRDeuTY5YQRX+6vSkbHxkJntOwx5
9vfs+1DbZhBDPUhtZ9V/cqfBOtQi1TnMVf/D6z0a+qbxTkglraplV1cuI2/bFrGOwdSUFTCec0Rs
/W02xiwdav05p4daYoAIFiyioFR/gEDdHruzOLzwgAYnzbSGJZ3Nj0oa2WJglOP4nVx1HQL2yB6s
E79ERNS3ftbV2zstL1PyRUKvE5yc9LApEnr4/xVQM5s/GStAaoMSJd9Eti+vJGXce7uQ+XPCBN7l
m+gU70pDsoPtASS0pfE6in4mmZUanonNdmwYmlduEPPatAjjJa3MACwXyH9QFpZTbKe4L8EhyDR8
EzfmrNB8MlzkM45eszl5c/kvoll6GQKGBr5asTkfOu3fOdjor82RbcdWb5F5FUPgPOK52TuzRmZF
913zdaELt67uS6vFqyrXG701ZZAwTbymZaAJwKHITPeJ3bCw8Emsu8kbLO2mKhOV/M3ruriigX2x
n7qUfnkWVLQfpFUmjh0rj0n7GzCEcaHAZZf8lBnGLgPLbjJUflFy2s2Sv3DqhCtztsUGSoEwZDqd
g74Ts+VmXIV2D5OoNH/oGk4AeKspoNZIdBxLN3UmcTcGoJrhE6g/qT9WIZor6PuHDzR+ZTwVF7IL
yjVkd261CoJ0WCTqmp71swIc97/xIh8YrHqHATPYntwXtDatI0GevYAmiB3PYJa5h0U9FktYlGgt
9UsIAnNS93aBq5qcnBplQQqUO4Mcwx1h0BvUQmqk3CykkWpsQ+qR62eloNk7H4NhFcfKeYBUV90h
++lWLjz2DQ7RDjRUxv3IfqxbYfSwHabYzZtFevTd7J89ejADh1ZR73CVdbey3fCmPu3wpKQ2RO1g
6zKtKYKBAZwZzaPYYx3PE3W21WGkW9KnZI98cdKgzeAROpQGbdPLSv0ongRQw1Vy3DjignK02kp3
KlapIV47ev3eaXk/l3PW/uG4OGwr/x2e2v1uO/GyBf8Up5nhXMxu8sZT2AuMFWm5f9PZtYCQs5l1
s4rk9pmuj/GuoQlAJUPejsVNY/3L14uCtI41fG3IZ1YCMy2MV8n3q0VBN7ZiiKo5j4XFx8kg5yJY
AvTuNYiYQUFbcgO7N2Tq7sHkCspmxAWy0HNZTqefC3Ipd0KotlWCYBNtioE1HOOBczmrlOZbznta
Usud0a5sPRhcS01QEg9HGaNmodLVC1AscqXK+EJH7ogJrZ37h1jcR9ip2fytDmczFpub7oQS5fu5
Tz+BVnVWiG+GtsMF3DDXIM4ThnoBWVVJkqwPoQuniD7j3oG4awpHRc1am3H8EjYP3cDD3Xoj9aPv
n9FUo+rpHpoj8nYDfUnpynWp2UGmk+ZyuFGDW21JLUV9IwtMpUltbHkhdzU1BvT9rE/j2GkRF1Dm
dNktcLtKzbB7sInNuQA6qvok0qzyS8y5Ea0Ldov4HI7INSN1HuBQb/3fMfFXkx5/E2MARuOYovr1
U5btPEhSTcNLhw6/JCcE+V/YxplthZig712tc24Mb7jFfwsNlerAGVwjSDUxMOL/xayn7gfHMpJg
EpJODWodKviuxHkq0BkFspRsoiI5Td7gVZbC4EO7iVfxAuULNWV0lRXsQp3LTeCrTjLT8KnMJ3Nr
UzCi27xVbcTSn5hqgcYK9JN6CcP2xtYlQOOkG9AJdfDNgQjMlHbcyZU4bM447dJIQTYzoUS0bkx9
GFZL5O5ntK+bfTwnMTaTXVKxxSl+klClUf/WaDaxJG5FEpDbfAAxLQjjW+Xo0HNYl8SidP6s3x8O
bkepxXZgUo/C73mfBY4N4bS6guUwUom0Xzvei1hs6X+Q7seOjDENqBIZky7qgq9Rye7xOnY1cQjj
k0W7p5/AWXF+kdscYVSBLpDYPN5VLkv0D/QWbKjEHlH+oNHD8mEgRQgmLsMs+pmjc5NgUg0YVFzN
gUggGkYKkSX0QP7hD43d2dScK3yDTt6+FRZI/ahO4i0e7x+Vj+hqYXgXYwYG3AXg2vEhj+nF55Uz
rLH1xaw77iHivksvnDyYSAyiCqrbGszm39vj78/SEZeW4mcv61CKFhakzAo0JqAElyMqlrlMJ+wH
2v16CZpqVylo0PG0n63L+iTkzc0HRBesu2x4JElQVm54XHO/RGXz8IrPnAR5OPtj8ynb1k050M0I
tGkAzL8W75IASqzDxXPQGSXNHAEIdjl47JLI8gli3YblZioUNvFv4KxXLiXgk6xLmWX6FjZsURP/
x1+6tJmUlv1mIRdqt4PUxWttcGnp5e/tuBs4wECFtbu3fx8HliKwipjK83acRWhYBZKLHXCeFuCp
DVhQ1UjxPazuj6StDD5+fk4KjYYbYYs/2F1TKX9ra8tC9ueH6NEBAI7HwMO/F/z9FMsSqOuGerH5
pJjphpmMavgj1/YuH/grzxGpU/TL6kbaIGdkJIqRJe8hHPf1JlAdCIq41pwvy5lkTAR71lQV1664
bTcharrUwO+FSSBsZiKdZ5lVIssWfE+BaUI+f4OYuiX+RUOVUuB8SAiW4Az8+ynjxL/53YPz1wex
NUjuanCmXZoj8z4R2SVfkgctrFNXPGyx6fx32GurysBlGQTORkGl7foWErXB4nbp9KixYWQ+niLt
XPEc8dTDy3TjDVmwxPd+zUi3eB2CXvg8BnK11qM/t7bYbNaCEGHRm+7neEcU1/nP4qTmYsfgo/eb
y+6gw3xq0Rg+b94pcolfvzTWTluivwajHKqM7GYBn/sh8hMxeMwLY35Fl5dGilnTfDsDqt8T4TEX
jL9ULoYtjYOmH3HdHBaLNFTBZeKrITAqmpt6QjHHAF5vQzr9t4PrnK1qdwYW7OIM2U3XXYdJ4MZy
qQtIhUNRLxc8OyDlxekJFc86W2y5IXvhFm4bdRpPaVPc4h+DRQCruGTFlbIcc3QIKEF8OZfpi8cC
pYFRKSbeHbHJUPC4uSbkDpIh2i6w4jXMit85lwMUT65BEeBu03iTTIBpKueUv8DZ54JdvbHCVtDM
+Z7BgthXufPmpXJUTnOS5nGVtcg3okccsD5X3l3BVCWjRpdD4OiBrWoIFDBZV411XZ+NwgDicsVh
kZVPx+MQrRZNmbiIy8sSzMGnUOuCL5v48201URA6ufTyxShJTWkjOJgHTqz89fsgraMI8sX36lhO
rgjXMvP4DLfshr0bafs56GGlSMn7p6QZO7OFx7VeDKieVaTP/plLwwI05C99WLAJaTQkbetkqrU0
XaaIpAiLcV/IlnMxHvHxdPIV1zDUKTheqm/nMipvaR44+YUSuuX+T3deoPRzOnmuxFu2iE8j1+bx
fJuO3WYcOsvRmmGRGHMmABRlJVXS42RBFuyOox7/gRI5eWaS0nNzV5TWZraSoRjcEV5Z2e27CXfR
k7utwtzsITyeXnVmEzh+ZU4QAjc4AbJHpfrNIAk/SyrekRPj6hDmZeNVnuIpo71qkhUK3hAc1EL7
qfXfCk2t6laK783o9WAzO9uGdNcFI1cRs6CMR5UBrX2q9t5xtLEEPCP7Av2mBKSNZsMxB33P0be3
MlVJXYdaifilIVIVlAQk18/4Dz4Uk4K6uOf6I/jiUQZsoUzYBgD7YnzZ17Jayd8JlY1NUfl/nKab
ML6r3l92b4mOKo3xJ5YP6ircJ7pMwGFhproupugDk52eARu220fVXhA715NvrLrswLqoJ044LZ13
ivy+oKdAUpQ/ZOkQ37ndxn6QSUuvcluTA2aAJwCzJogVdHopU8Pl28mxtORhiyGHCTGo/9kNT8wD
mE+bJO2RtStiwg+yVkYF28aOIjmhMQcC2B3HYacZP8vZq0Yifwhqen8J2UrQ+dqGg3iN5NyMmBLD
jt/aEYwvviBd25zqIGkd20QfuGcA45tNfpuMl81bcMGwbgwD3PkFbtpI4dMQ+70E9UfCyTaRfRe/
CRxRjefoasvm2FtqHmwmt1/tpLDHiFi/bRk0beXR6FgQiXdOcDkSFQWCf0czUbjUhe+mphL5hM93
nlEtHq/a8rp7gSv/ss8wTshcxrS9Aj4lYoFKq33Uz4hS1bCFNj4J9DLxhhPfINt0SAZZ3unrUR5/
PT9Cw58wLIsgW1eOh1hp6S/wpm6iWoAF9e0/DZcS9wvy50PVVKMMCu1LsfcEwY9TTHZeqF7v9FWl
Uw1vtfbMFjxuvAC5AXs2ExKn2fgieVMMvgNY+d/ztAC6rGaiRFk/HOYvA4QD2VZy3JQrLI+/j4R2
LFsS0Ig/D3xvITTg5QMKfjYBXJgy8ymZaYqILmZ8nArV8GLcOQV5kKgRXPnpnlHViIpa2TUMT74I
7rzkhg/UiYM9ZurXj1YRz6fbMatsLNTnd5zzwfvIHWEviqw+dk+7OldjJymVG/On1JcbU2emWwd6
w+I4UvFuGR5VU9ljZ7v9LsFpCY7ltT0QI0Q2B4zbWdS57DALYGd1DO7VK2BA4uUjo4LPRhf+bG8q
KJlSTTjdlGMjIGI2F0tzak3WijmueIECFag2/eDjWp9NmKkJHnYaBS9MVLsHR3aN0fUo7mwGEzpG
V6Mcc5RhMN7RR5ZT6VMPLtNdI0favhZi8mFCHhq5CmwNTcI6qfts5RqWmC4MCeHeivn5Nrg4rFFk
hic3bsHXcs56klC3cbb0iomuekbwQ6u53vkZKkfVwmJ4q8+jm2NicNvsBcsT4346rNOoYangMu1u
jYzp+0fgE6dzgbFNOctgFFSnaLtfijt/YOMWgxMfZ+2yBCwzz2Hf9uz+gZcu4aSCmo0r1ATR3h0f
w4PoDhaciX2S2PjAHFgeDpEvktPufZZIV0nGA5RkaBXBGdgY/sgLRBpA/5ewqYbXc7n7GjLNAI4X
WJECS3t2Qg5rNTEpyLCkLBQeDKg8T42FuW570sIgKSQmYnq5uCqtoDfVAwxYNjod6Yz7yRlIMOCD
+nlY1rxExCZym6S/d32TK0weyLS1D03pnpIqjcRKrbHpXOTcPA7dXD2Jvx4Nx/uNwzxH8ETgY1OM
0yZgUa5xYc8KQcYcJ2TfTlIUt0Z9yJId8WqWc+F01dG5EW7snv3mZx+CCGpMN+f+PPivMp/fb4nF
qVFLoxlQKhFXhIM9ZcrwoHHZJN6vGQR01fc5+HNK0TiKpJODy0zJW/8/sUz36+8JDkDCC85/RD2v
ZYZLYrA49S7VAkp4PQyRR6/nVoSiW2JKQxKs/rDBCzKFfuerS63nJ6cepaqz4Web77/TA5IzLf8r
yfhAiBuJJTGRyukR37vdD+4+xFR+JXPRUvR3911KUAy+x4f9nWQzzasvjF/Sd7+cWDkILvUY8PXA
O+tc5gtQ2vvVRykhh9E5NlQFGnCQWlZxBtomJ5P9RD6RV/q3F5fD1zEK5w482YnKc40gQXBqcbeg
0twSqZymw3Ye64EQkk/DwDfWe7nPCgWhDiYYstnxaNFxgp/9z5WJyM60jyq7EhpxIFsS+Y7Bj1Bs
iIjEmHU835zAZu3P7JIfSx0fcZAZGr8TDsTq1rJLSfupUNd5xDYciR9JCk4tQiZp4xt0E6rw9U+6
Q0ftaicGtyFFwLbsMIKycRVJEQi9yoNRachXiE6jwK6NYSb1TGNoQeNZ5yXDN6FxsGnsSqkxm7CS
9V3bsr44kKeAyHoPbPn0iBkdUJhc31+sKAYcaakForOqMdGjxXLTPaeI/UAn3GbHtZBX1DhM4Lh9
4Nl+ugJOpupnc5M7CYayZ52+5DFYjTt/Ag8Wgt98FB3bgofj1uuzadkG/NlU2IBPRqrNHDaPKaKp
oUXVOOxNRUAldWqf+VMr3pQcREkdjdt8tVRUoFRPzyoa6WTLbdvYO2KMoO0rIpdp8DDrgqFAZsvZ
JFOdiow59SjlazJEaLwH3c3aag/Rc+cVe/0nn3XCLWcSRdPVweW9scPkN6yB6cBA5UhjoW5pyOg0
QiC5zCIl/EqMppte/QR1CyzGpIeHC3jVy95jul+CslwWpjhJu/R+TN4qTK0BOWeBAcPh022pPXs4
qGYcfc0GLjxB+4pRPFuyojTaB3eV6rC5piqGkU0oQT0KrKVZWx0mI301AK/qXrWmGz2QY401uTNx
HI4fZH1Eg7R94K2nEfkzUZyFRi39cKslDGMEJMSOfDbAUm8kLQDAmjhH/dBMi4lABQ5rCr6hNZrN
cTSSwJ9y7N9C27LsV/Vd2hB2b04VVLrepE/kC+GJGoI37Ncx9gzMxIMKrqKJJLmFvhckE+szHSgg
T3wjy3AvutuGvZwXW/iMaHy/ZgVdlLI7rbHuhD6P4cUW7ZggaTj6apJMSih0wO50dlEq/o0mlcIR
pN6SZzyitqXLkE9ufkLGcLzova3uVw2RDWumjPfr0t4OwRHidNKAg37RC6WmpluKixF4NyJE97Qc
vhmufmTgvSigQjxJP2RxZRNW323ueSH3b6MlUotw/s9GB1hhyrXksD/tl+aDIU35F/WnBOmW/giE
zFvhxhKbx8Or/Ni4YBGvxPtKLs4LodU8sg+/aAsoR6e5wfocdZlDJ7C4v2X4xx91L/XdeIIVFhE2
MkawjIgy2cp9i+sVYCKpkPP0lpgjpLCCGzY/1CeEpWlijxYhfgsp20AHP/8IKvr8YD15+vlDULYO
+lrnPWWin4muS/a9CHppdSqH1sOmSWQet8+dADP+6Xqf6kyQS5Wh0ar3IdeQBvrbOvUhPQJ7cyGn
DIJh4FByY7jf4EwrIS4939IrA34uQcbHuuLOUuIvkKFMU6LdsRh5AEBNeR1dBCSK/zPvpC823xTf
xt+2DTh8HpdMII6fQKA4qqRGBPYp8tMKc73V6w3sYO8A3UxEbF2g5X0pSOA+2uiODoSG4zc5qnEq
n9j3ku7jMDr5yCGosncKFuqSIzxUk47b9qUcArZoX8JMPoUrOAs+DTxn6qq/hj7CGfD0lMtnKX4G
DgR68doh/GmNi5LIWYIpaUX0xhpng1Y4iVYuE/uCXO5myPaD4ygHJkLaGiKiMvriJsMVppQKOSod
Be2VONwzf7QqxmA3MSFkeTXEmlndsoEktERVpEo7ERz368vnKPT+AvXiwfosBhkCpLNpKqOLtJ2t
C9jQelNmB4tZW90NLVU3q3q6IZCYtG/ChpNtyhPk08OSLj0Z9CX2sNpN49YWerZvHNvgTBG0GzqN
a+ioHjT6bEGW9r98qltm6DP3VtVuEYRXwT1S2kCgYh17ijYkskyLMQb2rWSVpRjVVeVZRf+3aXgF
5TvplTsJU61e0ZzbUy4Ak7Rb3duU7ReMSrLk8Emd1v2qzOxzzb+lA4b09BU3hf9DQnAWJ8RebKWU
tl5lRUzSDOxppOXEh//YcGWiAgLjFt9lIdCQj7a8L1gt8JvkwekXsG9xwxvPYzQwZFnnyjPnawlD
6dRU1UUVPm5mKar0NqHO2KsSQFtds+pY+s+3br17rHQCArhMIEFg49YJnNLre/PFeKN3d9IltIO3
ERjSUixBOBU5vY/bFjKT3JTCnt6mqY2IqLu5UBzPSlqAI/zyCiuXjbl1y9JfHbN9Os/IsP4iwi/W
SAORKrqxQ7lFsntipZQe1OvrfX+I71WZI6UY8RNPiLHRL2iC4bo6XmNn0jMc6sM0qBHGLoyesKfU
Jsf/Y/C/uE/UKD1fplbYlczb3hAuFYeDoLg9h2YzVCrg6CpmOvS7neEwjF7b3bjKEzTLzFBVpV9j
1XsikVyhw6PZ0fvjhPgX9lBbPe8Gi+wezAkeWIVqmy5AmHIEjPVgMjZV8hwfK5QYZyqY03JkoAeN
BAz1wPD2jxXE8UhPrHjq8ma0V2pStkWt5o+/0rIYHvu/7pq3G9jRnNZ3cEz3nVHt9FB7V3UY0B99
xiNaDs26cP7mf6cMES+Pbfi0a6zqe8LqUGS7cq4l3nB+lhsGYHkSwUIGZS3PlSbr2KtnMPXIcGrD
OwkUfUzjAWeKTlo/2+WQJ1yhorPerrHyTKUHvfOGHebBstN0EGArzIx+9Nu4Wxgs2hXXGldrLygF
2OcEuxlZD19MvYkhGR0gCKVMNPmpW/D83sU2S4PpH0t1ZTr6iCQbHUeo4PjQggRvYnm1pXlqTIYH
ehVgJ2N6A+PXqAQQ9yxYKcy8AFyXLFPmUxHcpjpcevjVOR8yN+lpbl1yDsEecv9WN4zbxZ9VqG2V
zjwpE77CwmYbZ8Mr6DzO9H2hLhHLJokP4yr3CP/9ozmbAKEyc1qTh+rptORGutEWzhzuTpP5ep1l
6TkmIIdqMHVqAqI8eny3aUQrqU6PX2o96NrdsQq6JCtezOGwKjzEepe2Jtba9ixiCzRRQ+drT8f5
Mw6evzMI8aW+KYXVUoKqpVPRp5aYECwethzPUqF0nglvbMuIyjK7XiWw/WUbHNfFF1PUSW4+CNcO
uCQBHx9VRn6WANCMkIb+jv/mYQ2MPmC6hevAXVVaCL24EHWZNDvzMQgs8j4WIhED/vH/PLe5gHes
8NbWuUAmbhTIaoaOOJhh8UEH9+SwJX9gUXcFkTx75COH243CbBLaNd6ss77oCrjpIJ1DA8wXD+zW
rGvOSO43RcTVSVoYaM54S7Ybc7DEsN8PMvHtocPLVzfH/7F2S6fu/MD0/PXJ6BVmuCyW57hroejp
mK4770bzmxDzAuFRB0EtQ9kb5WbAl6bUHE8JFKaRXFPcAaDPj4oxFngQzZIi31nxj6J8gY+WqStK
GTt4N9j2yCsmU736k7muWTQioFwYNY0jCox7ACAYQuz4fVosKkSPV4mufdjQaaA0wlQfzP4mVk1q
EWJR2wPcftcsM1XlcocWWzW6RN88+plC6/09CC2r7GaJjCeOzzuLYQ17E+i64zegBx2QcM3rmF0K
CaotJ0l3TfI8S9bWPRr7u+9gXSNy7qJ5HQ+1s/DB4PG85K3XdztjIvTKrW4oJ5vq8AM9fZFuoiJv
lolZafbkCuDuQ3ivTtBv7VO27VeY408o/BaszksXW2gRe9bQHJ+5HdpblF92UUv1nwzfTmltVY3y
fnQxgKC8PPgVtEjjkciGifZwYeQAd9DGmxSUlWgOd+MxZOMPj8itgDq8quob9IbY4a8W1XMPBnDN
X2pUWXQvipibpMp2BfAucTgpqXT2d9kKcaYWsQLuuC+694otR+nHOlSpwN4xksg3zf7Jd1WLY5tz
59ezezjcfob9xeXw/VRnvHNhg46hA28q76Sx9YQNgL2g/Nqbae8orFCE5qKHcz4goBZcNRXKWQbQ
HNU7VHxqGsUjNp+RL7k19WKlwRzMw6dgvA/KYMES1g86Cx5baae2SPQ9Q6KI2LvzOXm+qioCpwca
2Q48V414sxKPlwytl2n9RRVseFQ5pLhrdQQ3DJQHJvgJ6Bpdtwsi04J5DZo1fZ0UgLOJ8ru6CfQW
qbTZBC7vRp8YMiIxKNMM034JYpv2IpDEuKmTWBsdpTeTCjhF+Aq3se7Whhj2TinJLCs6DRsbTjv+
wpQzbjkPSgPnw+5jS6BjZ4wown/QJSCQ3rzLlj/9LuQt9g/J6ceSSw3cBIBJDpyUsjfFzo0O0zkt
liITlRLckhQrRV5PN50F3+/zFe1ltT82xx/wcGROm9IkHTgmt+sjkQOBk+Jsnzxmqb792oVpyXpF
Luk5F9NliUcghmL2OAT8/YllN9Nk7qKFwxFOYLL9yzRtVShLBnjnJQ6lU9LUfXZ8RYaEMnTsQPff
T/4Xdvp9wVq266kaL/nXr8RBjZ+mF/jOFiUK+RfI8AcrG2BPIsH4lro744uBSzvcb8ofzGIA2/Fb
gJ719XcGGm7DoBSt3Bo9HzUPWjLkaLyro2L/+PiHeZ0b/L7TA+TwzOLxEh4zjUEEViwkXnVfamDE
D4oB5PEZhKpND7c2T0/f+h1O3+8DNLjf2+5WkW6p/2UN7kwfh0jorbGwJ9+QeccDrZhEFMB3U1Dr
gPiSM3QTMohIP4/aJ/NZDxhjrElyktOIL1ejRIAclFp6HFPU89HOAq8jcvu7M73TT9leAhFS15ba
Vh0HaWTYInyBDUgh7iseJA3LeL14/wDkbgHstUcRqC/msFQNEQ4WY8pe5KWtHRItFt4TNOrx8wLD
ZqWumjbtUy3aettNz11VGj3YKHNHcJEYZvxGvfEmZ8dFPvQhqp/Ai2cN8s7A58Qry1Of4NrSCnUL
NNVio7KUCKok/H1+XxGVAEHf1kbVLpaaGKzGPSrCXh/3gbY9sqbxfC8qUTF8qVOifA/4ncpKK35v
r/L2eRz2WtYw3gfrwyQvcRoz6JF6goyPRAF+gBbe7Oxni9LJxs8ilFGnAJeqxnhQ2DbSvMeACvlJ
K9kawmgTHGufbev+sEGYYmlNa+40kKE8OzhwC0y/t7Z0CqSAJf3he6Rv0hiYoxCETtuuCkB20/Bn
2xNEsXU3skYIbonATQWRnrfXbDhv8m/SjEyq0Wa8D/oOaJT+oK6bTXqd6Q/RlRNfoA0uohwiBb2X
DvghRtKlq0ETg3UuF0sJIQXizJjqX+8QTBMLjlTUbhCmW2WutJcy/6txchk4Zt/XtR6EGQHH8O1D
xEzIkW05jTDzIEcs3S/zbL9X6Vup4uWORxa1mt6xj1Dl3JyLslwhBnuk/E3Nw3p3YWtO3o3Hxjsw
V81k44E7HjEHBHdhxLc1MqBQnplG3RsyUZbKok/KOlothmsyNmF56BFRfmh2dQRaH+mguUkViF/q
aYAMtcUDmrsNWBH3gaeoChzmhNC/eLaAGSuZUWR+VWX5JUBwS4d4P2JGLhPlexf43rGawpEJ2hy3
rQg9n/SS1Rc5dph8kd6kuP0WFtrLnqR8byeYlmcOUnZ0hDn9aJqeQb1JkIkXrdauJQiTzHPbEHju
tDWINKIYwUpnYTGVAnPRo6KMuU/V3beV0J6EFi2SLjYs/S5+IHPZzazctVt+T56ysYp9ym5nP6hj
xox523xwIFwYgFVox8yczb+DZgmlxpT286JN5QFfe1uJSzY+qhsZpLFEgXQTfIpeDidgb71dvLYh
9C38RXkFSiE0mSL3XkrH1yEoiUA3C9oRAayMnRauzyRXukR1l/swIl+G2oW4S5hQ9QxhX/ug1Syw
Z23q+OnJ05r5dEebIoiW+mq1ZGKPo6gfa2lMIuPT9VHsma/nnxKtrutf7iuardx0E9jglhKULEhz
mleRgRihJazs14zWCwQUk85nCQml4FRcIOemqGiNZoYf4gK70mfdIRkE6kdNbPMC3Z/G2474Z1uC
RTI7WUZDBQqdiUkktQ98000X66HkSg7naggifSRP0+9xY0RjPul8vi7Id+hWiXGaQ0fDLOHl8txf
yP6Sayr5pJhOaoOLH6P7UO8XhlbY6GpK+RXSGrWyJeGYWAD6GlBdShnbplru7G6YwBcxyYvl84s7
LOkOMu1epYHK4OzbSgMisBFUc+wPhp/wEEWc8+FbXUtpZztSku1aA+6W8Gu8o258HU+15FtRFHDr
cfIcVA648Z3W3KAjhAy5EdUecJKSGfPPmj0GzYyKYs/Q2SplAKcL6RL5a+xbM+ugO/ZmcBm2sTOh
xNp8RLSUQtLGkIL3I0UY+8K9CPTES2O9KURC1zVHIF7NSx8MLDMIFBcQmL8rndiBpL65nB6SkivN
2l85cU92e4i4AEwatSmY0L3SSR13D0ocYsZ4WtzxvgrMQ8eOVfZ4YieIb5hs4FbDVpj7Lr7Rtzmj
lvw5+frn6RopbiclotnujPzEu+8AjsiCLzw=
`protect end_protected

