

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JEmZWuLCZazscYOT+xp8tQcgcJoo9xw+tt17VTk0Ee/cpOS713F8lYXKKz7qKA5t3FpvNSj+LwOT
FOkmwv2alA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IW+w81BdrtEdSrXT08IyeN9itdwHkCyvXK5q8xF0K0oVKDwJZ55f8rUD3UDvvDXIcAjvU+645JL4
ch4hQtC7Y2FokqIuMtHZi7cNrCDQXzP1bGPJjMCZbuYkodHhhDFZq0vnJHG5npJwjfiUcFOs/BD6
321VxRY2LE90m/fkP5w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mn15icVDdA3CjzJnkJvEX3d4TytP/AnBNj79QG+E3lCes2UF2pZhqISOBY2uufaQ44Iz0NeMSC9n
+tRGbjECz4+Qnwa3jPWzed02j/IF9RX7XCNKwHKcmJw/yHIa2jnhfXGycV+rW2BTSaOcvd71AX8c
xlCKhnyKdiYayGwfRy3hMXLuu2cdwaKnu/UJ1yLUb2SMopRlt3x1/DS/ujprioIUaznXnUPKvPI+
tY5o7OvS4nta5AxgAsVoz+HHq/K+cZ5D10lOXIDOatM1ESgBnEMFZa0ND/EVV3+YXn7orwuIkC9e
CVEV4WCQjR+/QOWg525B6zV97OAe2sVt80NsNA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3K+sUBRgBhLO7z4XKbbFj5Dm9dnCnLXJtz9DyutJQ/EYt7E+7VQGJ2l3bkkVJ8bn/YxKZD+Rqqzl
gzUxIUqSuvPPGmd3z16szdtLqj5YRAEZVXdNbeQ6P/rYfI4kn/0Qw+0hS8K2lRo5EQLrCely7fSf
ojGqs698Kv3dVxOM2uU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EHFOd5L9tY2zUSTwaEQFpNSik2aT5WpldK4px9GxR5cWZzjNzosBm4ckg29GsE3hW7YJVXJwn2ft
qvaRBZQhqD+DF8s0vynZ8IngOkOgp968BazD+XmnNms7D3n8pwwWq1DBwFf103zHNgk183z41Fww
ghnhfPrVLnkJtKMArkX+0VsxpoDgdODsv3fsT7CkMz19ja8WwHPQXCAKUD3p2rptjKIU1LKJfHEW
xgEccgVmdaHJ8o7kwvdgJQxZnf2Fl62jKVF8AJCrqXWKtvakZCxpEqbYNpoJ6R3Ns/YvtWdsZkRH
TW3+uPSDGYDVS3Az7zcuFIC462DOhpyBpwOGGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31872)
`protect data_block
5+hGd1aP30cb3O7GzG2eGqHxpMPyCIzrW0+NvWGIFZCItopWvEx7YkxjNF9jHA3CyjkHTkvONu3h
oztuclnEpB6znKh99TCwhZfNZazLkJmS2eqzR9RXkZMl+mgOhzX1Vhr4O0iZej/NQL5Ez3EoITa3
COdEBc0PCchfZo9nhCQN4XCMao925QlqpnblunfLJ/6Ta1dKMPBd5s6xAPryIxJeuoCssLu2AJYK
/KdHPYgnwViWw0904i/IP8Ak8KsRqAoxKqoQ3q3rzjhQzix07k4KgJBYSeDlO3LkbMxWJI/gw0xs
0VmxiMwnPdvkCBOMQxeS1F9RJt2iyN3lHKsfRVW04cvNqRZwnLoqxV4lctDUZKfZGeb0sQX67YQq
5fLBUg+EzZe9U/kIkNLwv+fH42DY1BYEV88b7b3+y7sex3C4B+vg6N/hPoRUVROMvwxldz+FBVWJ
gEP2BtkUFjsqhAzRgBuqvugKWpSDYYhSoeJg2A/CKzbrDpEo3fH9nxelM17sI6nerFENaaDCElEu
i6rVykcTKJ23fZOQqx3FqAGn7ZxTLufqwHubeGqRUZauQtXLn7SQnhurv82xccYibF0StFWil5Zy
8UDnP/aFigiRtIt0uRaKRTLUc1WHS/ot8bSIoQLRw2zrwPFc5+mV1TP84mccnTbQoXyokD89biU8
O3jEVCFsM76pHVQoqzb0ptyKACKAdMgLuZIQMYr6jysle3A0zd8yTvfXcEZFxnhR2WcK/5xW8p00
EnN/yHhRV6PInuXCD8Y+JYp4SiYa0rt+6VRQtg1WJswmUFpoMfo2NA/VN53iu0iYPa5f2adCsBt/
qwltUWWksIyRjVtIvIqnpB7dNqG83TwD1y+hn1BQFYXVSxtGB8rVGAZ6w8aiHT1c8rffnlclh7RA
POo6qI3CxWFU5JumedOr5gyF8HlnrQXvL8hjfTR309vK8Hmwy7XAsqw8EA+kyt5qWO5qeksmKlEG
tus1X4tbFQUDOAgxgnDsbn5k35qsHR8iiWJ/mx6Le8z7qbtngwp7xLEK5MM/ceLOytifzXrUXHV/
5mvKZjxpe4psvwMzZhf+RLNt5FW3UtWpyU5tFDXQ6qtXTENtOD99CwUCYYFwrzuF/8QFuwLW12C/
X+Igo8Fg6g3T1Zv/CQK5AVFFBPxxw+F8uMKAZ1Jhu+AnOZuNpOKDTYGyOJqt4Wv6mxOouWhuAANg
OLT00rekZT4rzbEyKO+dD8uaI64wFcfpkgQ86lKE7fPsfVWPBJJonTrMiiVsGnPgkreo9g9UdYiC
3Qfu7qtDiQHko4Q1cj+PuF533RhSC4LxRUsOvKhT5p0G3a5QJm+nheSG/f4mTd/Bx+F81f2A+lv7
mUzkvTl1t6gwld/rhFJjL3d0ATCOd0Qof+eZZvHM2pZUrEgLVmCaxU8XNer4YrxVXYw+CpPPoTu/
p4YaA9/KgU39mXiVe65vx5OgWT5Fgv6L1B4yLZJyBIwUC26DJFokGjQmMIwCt4LTSH9q/Uq0NaH8
KJDM6CV5Dp13rR16EQcKGxtVuTpvTpPq0QRqpXYmkAmwf8KlcK1qjAZ2jSWBwFs9rVHnQYCsIoPF
8RGcyQ/8DwXvd5nzhxQcNaMYhpc85blEtXSMEUNa1bxw/re8q+1mPL23TjqMoSq7oipbN9tEEUZ0
wObisyJTcRXpFMD5i9JIQ1wjmMtHswSv337myzZKrpAQfrGzgohMNLG8XEZo+nsBKdU+KZCWZ06A
PyYRHIBzQ5v2ubFyYGOXOZc0gZWNRl0jZiOJ14pTvHZoOXvNabFgXjsboR6kcHIUHqsAE65MWJa7
fFI1keiHG6LDxGnCOjxgMbgy/AMHJdurHbFql43dm52Aa8BUOcqO9N6LndOLaqTzQlu9PXdB8/Y0
eA6NzVX5q5ElJ/V4lM0qu4Q86WS4E59TfXEZDKmLLAM/yzkL9Xn3lQpX/tIz+YjAN2H30Y1WEU+Q
TN3KxV0VAm9xTN/JnjnSllv5RPRlEuh7GkwvXuQa+PfscG0x5IEuOeWc+eN5edlMeL9n6p6tHkto
lKQcR/kp0Q0FXwVphYdzU/jkzWzT1s4KcoFlP60tEbofQka3C3+PJ7PNNslhnrptNLe5kc23bF1f
m3UCs6bBgbH1tXofa87WcgdmR/C331QhwpodgskhAbvafEK42A5Grx2X6/sQJ9OvF5Ox5gWQfJ6J
f58qAuLs8gT58ftLOKvPneYyLYyi40CA3A4vOA+IocWeHlb0q0ohI89o2jqx2n5gZtAWly1+czEr
gkmGYYTVWIR6ah/qzRJkpxCMxXg1F4QiTpxMUNoO9lihSiCsceLR+nhHfdWaCPtBAZTtJ6e8lGpj
QfT94GVAoHBvdOfCQ9RDTPv9WCaNI18UmZ4Uc3a89RHoOEP6cDRCS++X4boXhURYT0myIdfgvmXT
sEFcfG++KovHZYqMC47l3aAs1JuUfA9fNf7mfJuSA2xEMLfuE4NPDUWpIDJuRZBmOD2KhvbDBwdc
4OL0K0XtnoOk4Nqtct+ysW/w0AcX5CreUph6/NTt7cS3AoklEAovZFqVNuZRLvk0FlS7thxbj/r1
4/a7ox13d/zQer4ose1gy7o3hDgLM+RtqYyMUjVbkVigHHOZKDKqxMyL70FJBdwsVP1WZugVxavf
5OraRohWq4x6mI9lRMmFSVHk8q6AINuqwrPJ9t0UoNN7r2CnM4IOCI0IX1tPOO4V6aSBmFXXhBFd
oAnbsu1QX3APRuUGHh09J08ILFikhu9O5pIa2Lpif/XX3+MNBYqXXmh4kvfPp+qfXRZuJ4UR9Wpl
phbZ00YvsnQyiejLfFfUyZJksqO66cWAOOx5tbtdv5hInh/AEYO+lnr31NBz10lToYufGGX7KmOv
JfgP2qA2UNRTsVES3dOAWVsOJf7Xw7FMixfJberc1UnY4mtp9K2lAe4HX8byc8Ij+pANPqH6MZms
ZvxU0J9Olq+MFyTwzb139WjW3V+0RS/LNGLZ5VD06CqmJsK3raOlQX6P6z6JtaGfiPBgBHApl0DL
6d3FSM5GnZldN9ipLFGuU46T0rhlEY9ZBMRSRQH6iiOk/bvCLXw56oh2wNBT+Amgc3ZBtLYOaOCm
a2nRyGFgVv1se+63buL+mp+yOUKvXSWoLJAO/4ms50tEgoOuSrOAPDFRynaAfZcb8ibTMM0xOZt/
upLBfm+zFxoNKYc2v3TVb+xDLxbCraFOKBa8wZn2ThUxGMHWngVZeiaQzJp83lYBSBQ7JbsBjvg2
yYuThc7TpfHfF9sPODmbIYT3NpHWoUCOkfT9GyPccGZLLm0OevyfnpSziJ1Yx6raDL/N3p6/RQZ7
D1l2viuJSxCHvXedSzav/r3nOxsUUg5VqPDP3SGotZrLB99I56ZdSZLnCjOFWwXsKO2PXINUfJWa
YjMRowboUaZFw3yttCv8b6MZqOGhu34TMyNEDimgFvd1CUzSm5O6rUYHd0RQM2EVPotx2OhOLPJn
LcuRU4T5X4HGK9iK4FViR9s2uloGno4cL+qhedulDv1zuKQPrElkbyentxWCoEAl+49YaqnKx6DT
iCxQ/0TyhFC84HJfsRiH+Tn5vKH5A5VJCI4ZhAXhvK/7jglE2lomLKrpYW4OccJ6xxOCvYS8v75x
L2KZt8sMF4XbY8wWIQ0r1wKK2BongWod0n3PND12hLeNeXJrVMwcS0ZxQzsrNlZH5rtEljDoqBhp
E6p/m3RfWa1UfbFt+JLmjpzl5QWMkEgfw1aYPoTy0j/eDRkDjcvAS2+OEwK8D+Szkvlcktx0paps
9Z4f0zeNazJAuvtBAUtS/NtBDd+TdHgzh3nGdmotkh4e+7QCvxGh/GfVHFChb8PYJmEmkZEjH84V
R8nIry2uB7VXEtw26zGhkg1o5NNfnuFcg75Wf8PH+kgQUPidGGGisjGHoEzWSN6CDHs8rjYYQnI6
9bnjjt+YSPkVMNPtwZ+5jM5hcckG/aUPjo/wp9RfbKMj06b/wmPC5w02nJOGPT2iKqTdY5dYBJ0J
KM/FSw4FD3+XW0C8sfBxd5/uhX9moM4VzqgDc/6fP0aUC4A/KXUnXU/CqiPM5XoUV73glSI5EHIp
6fieIaCdJLbUruMnHSuHLfO+10qZx0HPDGiyBwqoACBEeVPx6Ktdw6rJGJCW4mvxq+ocjGRW9xst
C1BwRQa6/al1vywfyvhyUE5osm9B/p/v6yhjYBneJNYM9k6M74I++4DSBkphbMQvW7jifjNUkmhE
KJJu2KmVV94/DC9HtOHRdZwkt0lu/yNCATYQovxGEk5gwH2DfIxImU/sVXHs5hf09ouqsz1czV4A
+MWZsmUS/pRsuAF1M7qOwYCU1lIOxJKg6zi4ipx7qh8qz8ghXBijIGC0jOSSpESxtS9PyH80HFtD
bcSNF9QE/WQQtqWhccYGpcPxq8OTeoMPBcj7/YpD4CSTxnbsCbHSViglwE+hCYT83P7rTj9xl5IV
lphXQttxA3wJL7evM56pxkNcZKgPS3PMxEBoREsK4jZIQcbhiPw2UipKzMonB3p7IsQv8zOisZkn
oRDtAX9jjym9cReoSRKGVpjYexHQrix4mwN7IFabTcO3QK/nFdMdjpACpjybdEcEknr3MRtzdTkv
nE3dJb32k17nBtseAiZT5m9PKU3sZldXgXjU43et4xxJJi9rY6W/RXD/k9AMJEKk/opdtua6FULM
A9JSupWGk/h0PM1nylNOZcizlenF5FJddnj3kUp4q2csA4V4m+z/klyMqSMxUp5nDj51Nyd81kAF
3l/05HQ2X3HiXAK3YYTekkFrP1RNLbTQ4u9U6QDEeJ1Yz1Cvnik+R94ga98FHCfuRkW9J2JMlxRb
60XWN/Vv2tfPeLlIB4Konvvy5tpRQn5gN8K6ixdnDxHrwalXEGeo+K36w0HL7r33OWjL+/YFoQ+r
HsfMzCp/CH8MHwRlWpUWkr6shXij/Wj/5Vyzs6EkkIHd5w3xmGkBWCpJrxSZCScIvTZ+3OaVLx9z
YwFcW3BAyD9AnmFxaSbeJNOZPRb8tZjAX2dDKvfxKAxFeaIldOQTPm+/AtGbTkw/q6X1gcNlDWND
uJQ9NKB1dwA6uDiBzXKaYtQH68qmZ2EGHrAQ0vq85+czYaEUAzT63M0hXnpjZ9OcWLP8OXCuYday
uFwk+/3sKs0hz1REYn0xHJsbq9lmQGIcb5uhgXU5ptFsDpfk8TKgWr4/ws5YRgmdbxcMHCi6VaIN
sn+POSK4SRLLJugpYUkT1JTBR9QuF4I4CT008K7QjpLN9VvK8isC28lfXG79oJGw9eIiacMzQApi
Rq1np13xjAkBkicLVNGduJDrpqhE021i2s1xPnnVcTHfrq/FiA6Ke5caTxzy7tQFrq3Lwl+/NZbA
TdoVdR7AVLoL+VSCAA6X0wr87xXwGXqVzHMt1V1/kwA4evF/ZY3S4vjNozfLYP1UDqSXEt9BOYde
bvtH3IiSDNWQH4wK1CqOWY5A8o7cMwqVUBnWxvg1hZd/cTi9gTakjHB/tufDzIxMmqjzd/W3kINF
Xe1YGl7zLcweIWtRc8TGzmXJj+fa2E5NMZBKrBMzx+PvUnJ9N/P4AOeISCVEtd7I7RqysQK3h4DC
1pxPlxHbP59NW1ByrhUbwkclh31ZnZoQa4+vnp+A5d4wssQ7Guiwu0Iz85qoAw6bOQvvAGWrbD5v
WAch4ykCu2axt0TK3H+LrEEF6MEsTostlRb1Bv04KyQ353nP7NDOuBVoC5ZyqOwUSPBL67ERjrv9
zoyg2wrZvxAVrGhVzhb6HO+WDeWHwbPg/H1z7dYd3I7ubqFjtErZcYKX6oJEM1/XU0idvRsiYNKF
rK/Pv3+3YOo+QRjTgV+3ZQxA57UUhvJbO9S7efQk7yBLa50peHSxs3UomGeMgNW/zdve0h+xfyow
mwHqUi0ObtjCSGt/PdnAJ+DVuJzrhxZnnyUCTnuJetGAdv8cldJXwItOqK324aTLsg2DBmKBkzJu
wRJAVEJtPlZh4wJ8vLUZCVXelqJYxRR2ea6HkWhcERem0a41IleBOwUP6dyNUmRX6odqzDn8wwO6
zf09t0Kt/9Fm5IsAARNSpt3Tl6lwz3/ojF9cD1pJRPRyfNoppwTShYDDtlYeig6D9cqOC+XhMRXf
YpRB10krYEIymxM7fDe3oukiH6BwRt/0Wx/vKROmxYah7DF2pN0YAMVxkCjwWnLj3scZv+y07feD
dkRuXt30M0u3pNg3w2Zo7REuPXp/KMbbGWisdsuhm72IBxVmMQtBQrMDyyof+B6l0TnVPuvZZS3e
Et+5b3rLubcr2g7njf+CdTuUgFcGiPvvLCBXYid8tIiDfgEhOWemUqUBRbYsKPMLk2KgGLW3QmT+
12Z9Fufi+nhP6d9tiTrBzzSSxL5bleL4pjwddRRStLfWZUkFcsY+h/qa7QMoD9wGeYMlv7ynzT/2
qo8KNCcoonlZT50gPjmrpVyQ1Kx2VWLa3UeMpmj6IbzM3O9ROlc/UOWP2VGiOEMXzMLTYFZ33e+W
BNUgumWvdjlwyUAKnFFRY5+7dSp7blPRcOVynjNTYRxjEd7a78J7XRGdY0llPSN+X6BGn3RnXoBp
pRoZ+xFhax7vPqZtjTmsDVip9Vl6WqPKmYo+h2nHHAJK+nuCr0x2h5Aex5kM1PdxiKChNNJrPyiX
iCUgpdDONzVfj1o8UwLcc0S2IYGqnT250DH4wDofQTRFjcadowTH36L2JG3E48Xf3IQJfCQu08Kt
VHaHDJyxeS2KV/fryRWb3H6068KErpd2+EWB+d9RyCdgx9+D5ebVdY8yiUnmZ7oemtMtE13ZE/gx
yDBx3myLDDgbxRCCoYyQyUmY/DZc/FSaFWMOMZVMJqzxEKlVvLyDUoxhN6YhtGhZu8RKhEVAiwYy
riv/AfBVIAEq/13I6vaWqDJv46XT5gNRxPV2jd2A4NlpCjZ6YnwjA2vvSeVsaQX4aVRcV9D+vhEj
KkAhtC1hdI+PW7umxLkydCpI22YA7EWH4LER1OkJHqoKIfh276YTh6HoYMrUis9iMktDY1JOm/ou
dSh8vJYlAuKdqRdRFSahaK8oUNScSA/bELc3/A5MusTwhNHDOK24TmSZJ8JcZeZFa/Rkz9TdUjO+
LG1XlXXRXXGoI7DjA2kmgkD9ftYaIXuccCYgkBbfyCDCBuHbYrJVcwqfbn3sKUyBo1hQJumoPwUM
LtxJdDotxE8L24pVzlx5A4czYTXGPxfO+/dGc/U8z4eGWln0czOHGGYb/CLDLNbmWR6fiDKaIRoh
1uUrGMQlr4EjAfahT8udyUnCsWyxEnahHd/FqjVh1Phn7zbnwdpjtm9/cnN60fQq3hJ5aWxwL+oY
qgVjteRNvhSuOD/ARUMLYxeXeM+dW973qkvmOg+wP1PcKMiRFYuDlkzDnODILS0aOrt+HqQoIsxy
6RnzY9+QxbpcL2YXPw0Ba4Cykm5yPcB2FUIx90Cf7Fm3oP22KkBKHRKq4+7GD/+iNZi77VsxaHW/
dXpZN2t2AI1m3I2tr/V69898rz5yw4gu+g5S7WW9SQGqE9rQEiH7u4lTL71u+LUFlrWOilt2pZ/8
AS79OmnE9003jEurPl0QueE0hPB8Crc8NIaR2THYt/+vejpRorv7qpOAeznL8i3Z07Nzy5aed70A
gry31WYk+9CvUOIoz+da3dGq9LMgep3gLaTyzLDU+Xu3t1QOOtt6Lf6u4mEACmpQiP/h+LHeHQS1
nYSkNxzVhZzya4X0I3NpJGYGVBcOJ98JwU6+BHnSI0q91YX79BKDlWP7XYW/rI2HgZUkMNvxrrRh
R74jC13tkWgBq8siT0XrEa0DxMScss+A1NJguRk31R7J2rsChorrnF5ukiFAmqfVIRxzoZnwLIQq
azyqsEKcQ9xxCjdceoAz1qmDaI1eeC30yPr8aeDKlxh4wzLa0iNuCd3vkD97LC23tnSzP4cd2tY8
8U5UuWeQjeiL7HZRpIB8GJ0oIRHytB9rSSfDuZ10WjDy2InzCoFuE+C6snPu/pPcecRx7dlTObPW
L4tcV0T4k5h40UtJZoyuGGa4iJ4ezj/VEVbXIAyVnOsFWphmGbr4V37nqBe9Bf9xHhT5pc9xmXj2
l8lbDCB/jIs20gVRgdT/QexnkgmgeVZ6ajELcQ/N9sgxzIhNvG2MlXVt4n/o6fSd60g0nieSptAB
Zf6MZ7eV8IpYdLk5N6h2E2HGBmjzGUUPvRlIyo3E/cofPNKPTsGA5DeLcU/+PJ2i+R5LpcQfh+H1
TjkhTEn+wbv89xVF6bS9ScvzjoI2g94tXc8JAOOf8ws+TG87ssiyERxPwl4uEAfEEL18wcFgVdUF
zDIKKXvOJjGXEDRE1bSDj+el/UZQkxInJLeX3v4y0UWuuC9Vojwz6aGRHA/PFF5ef0LRKy8lL9u8
KJKHc+1lb3CU/tk7YpesxBVxxyUPS+lUOi803Gvl3fKJPlJHLasmV6RDg/FZqWvVhXvvEijwoIbl
/CcL9fijqixR+yC8J48AfAtpqsscBazqOVqVBK9WTVdjb/+eLIFB9so5g9F9klwSirBjnWT21YLG
WvFLWSdfgMYnuTh/Vkri0ndCIyQ8SeRoFp/B6E/pjgao1C6bTQO4alXyEjY3kB2oQv+pxOSrVlKR
2/UobAwHvc9luQfSz9Fye4MYIUGtoOlSgyz15kB8J8bunyPRqhZU0wslEU7otJ3MlRnMDtpckE2D
p6fbLUGhHo4S4NPyewNz4gBGdTN3M365uVBWaBuTB5aItH40UKBnIkW/+x1qT/Aw+ZGqXzvOxvPR
aDaOVdapKbIwbuf53/+dqq9UiG8wR4xMDJqVZynmVzJk3s8XAFyj+PSwfPun0fryD1Lc/fFc8vjj
XYfVYK9eO8f6Ranfq+hUnPFhKeGyxhByCwKcjV4yhikC5piL2LrNW/FA0/hEhYbiVk07nsAqfpMk
yGhPvhoYBD1T5kdl3JHYkyepAek+WwlUEg/PR29zEKkqRmUtq1AQjxBusv4jYuawVXvGePm2cokM
oJQOOnfaeWq4TIWWfzr9oXURtHRpeuVvl5U+f22z08dThDDdXWNWJR0RkjYOmV+G8t1eCTh2Kbwe
2+o0vYq+82i66+AQkbIm86ougyjoHxN/1N/3qMdU/6VKgM3canMLY3MB8P3m3x1neLRrOI53qJrX
woiTypJ/hGZlyv4c162+kcl0jzQ3btO08NQWvhs1PSiMeQAKx1h0giGo/9SxzNN0S/S4GLDkag36
6xjnmYK2kE0e6pOy/gwM7KLq09IOOdpojl1SiDY8jnxBktIqzF/84D5KFaszcVU56sgRacFyKfZU
CxdeGCQ7rwENmv8qLUCVYuATmCgMr3I1ngsVdnW33QYLrgwxjoEnEdN79euzgrpX2pIwl62k2ctK
Q53Stea/z7FLk6wWZaHXGKwJYrc/adH8Y4L+hNuUent66brwcLdCC+tbmp1Nv9AHw6zi0dAl25x4
XQqx6Udqic1muzLtyLAONvjs/eZPr6YXtfdR02Up/cYCZVGTo+iSdWwqGyR41yJhCiF2F7MzfpZj
4fmT0cLCL0ugHl1Su/8YVirdkxYW9FpBWwDbZy/mdjRnw3x7/f8F9o1ikoptE0W4gnADEXAWzTnP
EkhU7MdMhmFeRs8j976i5E9RmX4tAMPgX3ssRPW7DHDa9cx+s6IYiuyvjSNXpdCDYznlHe3H1J63
fw9KyGPcxQImPK+WcVBJqhYpzCPb3pQfxbw/9A0zp/RZy0AlPT2S//667eSQqEjIRa8B55/YNk8x
HU/EKOoYnwwbWLnVNGq30GmgNbGiwKM6yXXgooO7/APbbOdDi/pjU/yEBkk7M2pDbRfHmqlSYOpn
KZyQVBIiY3cm1AZdEena2mwSZf41cBMiD5AtjkIMBQaHYdkBszr1/aqu0bz+SAxvsuvFjPDJN/3E
Ayhr50FfDPGIiaQKwtN2bnSBr69zOPsdjeyNnAfr+oaOlWcqiD3iw5hcFwGgh9U4jnGIZ/g1AO4/
2SN3w0Guh+lg39DsU10kz36apVvfDd0bXWV4447mrlxz8leb9HtdRBKQgnU2PkmNUcUemdtm/PIW
DzjQixXNwzTI5PSrvsGNVvk59MG7KFXUrVneCFKSBrkg8i2VnKovOBgk1J3eQjMJu11SJ0HqV0ow
M/ec2UnBQI+gNk+QRxLu0dqlE0xlO23TjVxSiopWotgNZH1FA7eipG/SRfjzFCDTrTZQl23QUhsh
mvsVHl2BqZKVzJ7m8SgW6fJv/Wlv3J/dpT4k+0j+tL4Bblh33yRjDYZwN9fkL3WJ5sePCUQahJlT
KeupAXpYABDK9k+wtPTB7BqxtTHArQgro1IbrI8HOzgaxUSMBhjr3SFu/eTN/fujgJS24T+BLagZ
T2tFV4wOTovOjFXJnyE9xPL3HrHRZpYgatcE/4C9mgqtn0SSj5S4vb5DExhgvuuSk8S/SrSpyiyN
WZ2ou9UaVkDOF9CNmPYM5z8Dj3zPhnwaUeNM7lreyg2s1fdXi4tMGhdQbl5IlM6YoO61OLV2ezEK
/PjCkCW8CvTFfo0qghMWuNoDRt6GaBIWwMa9uOHn3GZ2PhWHXGz2Nq8qrD/rXt87i5FoKjYJ/bOU
xYmwxLVU2oy6ZWPnBSq1wvw1YgQxlczkdd3usOYjytF8ARh9XQ6gHxyDQqPBrGw7/LiNqvG3tm4n
zwM0JLOV21SR6m6seUYL+fMyeR7/DavgyRdskg6YGNeWkcVw4PuKUpPu0YvS4PvsVpMwlQnts/zr
Zu24uiHSVWrnUGMmSScuds1sDF3+Ds+3a7COyQsoCmTEk60FziQJNB9wX1bM9u1AdZo73anchrR3
SBHTQsP6fY2d9xQVxZ4tUOWkMC3XjERMY0OWuTchLgT3vdKOzwS6m35inPV/FwWckZV9tdubF8B+
8lYgT0UfBmgEpCx19s4X4ikS0++FnMgtWMO1x9BeLWEkxM3x0tT+0O4gfqgQvPrYgm4v5vJxztYq
UspmEs8VfJ2OL9+DDA2CY4w2JhztA+JQjL+eprgudtn82Y6soUytBYRbp6c2f/Tyr1lg/72YnBwB
DPkrEJJVNQ0OQ4v2TlSWEP1KG1gQul0uHkhiwMb9ScM2D2heJKtLlndpWqojbVG30tV0iUi+TgC9
N1mB2lIaL0PtFb7wORiXah7TOuFwKtKeONlMzT0mJZmoga4qmfysWR+Ys+xuYEFqVIowbCA403zX
/xY9DWDjid/cvVO1aovh34VCulooQXwQwrfqi7x0AQ3X02IQfZ+Yf0gdjzSGGw3Qy5BL7kAil/G5
wnnobvrDGktSPO7BrBSab7tVoNAW8HDRVDRtHCPr/Qjd//8cn/9INfXpyonQHhUoOcKQH7E7tZ7q
HE/b1qMF38lu6frBds+X1X9CmMWLkt4n048dd6sMWsHtri7o4+n9sjKAwwH1lXqMwDfR4ol+vNug
Cr9Rp3Mb1il/+X3XFmIIkR8hYWso3e6zbxHTy8YMTLtRJ2adTRNA8vSTPYwWq8pE3uXPEVTanG5i
OCXGF+1n7vlZk74gAnsXb/vqgch8hsG6WNAUAt22I52Fjil6O1BwgAgFYUbAVVGBwgFIVnihN1Mk
mL1s8Q+mtTFWauufUWKUTnEfgiAF6MRTf5z5j7u4rwcK2uEFhGljmdqZzh6IWAtbKsKv/RYFOkHJ
1HWjbGV5fJQuctrTt54ghp05xVN3mWXkJ9MNfm/GVyYn7wQEN3Q/c01I0MbMXRwefaAvMzu4N5gz
qQG4+VIOpBkjsUZ59+pD2Q0JQ1ehWAyjGDxL3w/Sn5gafSm0tR5PeJHTYxCkBX4Cunp0XnrQlrPa
fiebgPXslWfXgK4HfGBCJG0u6DhGDQ3+brDUaN3rHv2gOxPDwK9BJU6FbSMXeXfG3NlHTePJxs7K
10BG9fMYDW0Tuby86QZ+EcxZw3736H2D24rgclw5qmqZV6WIJJRieVXVAw1MFB8BkWj6fCnuAQJT
LlzxxEgZEShJxHIuyjNShgPhlCX7y9/CsNCMmZfgXMZebVdxtboQGQNsY9IwW0wg8vVkUrxVZCki
IsWA0XtmnVRcsT53Upeqry13HfU92H9qgZHGlZEqV3rZHoUGn7gZi2t2BQNBg2jQ06BFX3Sq6GXM
JOdRAF9/UVxeHdC8v4Wj3ZtEj+iKDyf7pgkGMGrsE/YLFjAxTnSw3WU85uPGLb1eOA3fFNAkBMrK
b9oIErGVS9d8BKjnz3c4BNH7mUmppS91SbQymug+bdaLz+MneSityD6tXr3xV04q7iFHMuNGmGEK
KzZLD4sscrFspXt06HJnOnf1Tb5pzGSZHtGJQKi6jGZZNCiMHzxkZ2wKQq/CNIO2PqnYeS544tZy
nbOcA5PlaNElCQvbEzoGpcGrxbb2LKP3S6+9+iDOIzFNMlN401ALlutUleD7WsGHKEqFVeK8iJDy
jEAfsLB3VHkrppMOOlP0CEfSd9nSzWK3nLEgJMXfhKVnlPdNmLFR/utCsJKDZQi4TxlOHWn65Ae/
zyC4vUostgEEQVcTAqcZzv2LuAt2YXBmKXY1cEw3YaiY3P15aEEbp+qPcKQNvJKSX1EySzhfAk2+
wzPSJU7Csu05kFJaTJXsYHExPRTlk0q4Co4naAiu2aTdjcZLeISEKq5MU8S3oi9dB8ELlklKi6xJ
UwGCD2Ar0/ALpC2BuuncAYMW96S8zn5INfqUkwWGd1PfqvtsZn2Nf1k9kzyOWxIbWR7qtrJfe9Xh
I6fG6ImlbiOALdnNb+LruxJa0LrPzLDRgU9/dZ2ogOYTAn/nh7ph70XJ1tzZzSlmJDFVlZrnlx85
+XpyeBxv2pjrLFgb3RK5hRwYNH0nMg8QGruBflbDxjlxAGrqSoDZkbf/AdQpZ4d36xi6bldra4PO
B+LQqLojIX3Ycy3anZXrKQd2P+UvqIcdzYzsxG9X4+JTvbv+s6kqYlBifidTqRrkkE6I7lKr5r9H
Pd8g8YKPJ9A4bmn8AEJuHW2SrIEgB6oZuGGPW4WxyCNxM8sRuLFncqtSWBSJDxox/kUgypVLhDQy
LNetfSrOH7b+uIFyj7aJwWRBuWhxjv3VVAe/5SEavmw+bFhaGxiHxGcadjiANd/q0RZbb2vQ/njE
pKvKuTaLSLFQA2jxIixAepZ6BLcYy1DVKE1lpKp9AjdNfkLvj99CUvCFeJcyy/eMDfV91FaxeuMe
Z5pkc6Y8MlKpJ2eevZRZRjpbu4KLgTbbQaJ87zGqQzhsxUDtbIPzNIV3AS7vFfxYSGwS9yQ7F7Lh
Q3+7SpYkxb2BM8me+y/IxhCHXmEW+j+uYmi/LFZlKvCdhcuWU0pLjPK+DmCICXd9vSzLBKKReJeK
+5hvAkJBMpX/nHzaqj5FEJRqN8QcNFxN0leRTAf+eD7KUQn9G1hNsVYkr0HicfgcBjG+KIu+SVh5
mIjeNAnHjXVYdtZGBVKLdTrrs8DnwrrE7Hj8cDJ5QPwTzx+KE4s8imoyQjb94iK/hY0VPgNQbqzg
w3k6hieA+HGJYa5ai6Bijg7N97x8g0sljJBo24q3Vg9/XIsEJnVbWBGhohuBmv1HgM9yr7TMS12m
f8OMRXCE4+RY8gPqDnIyvIiau/vchkI149OUnePzLSpZScUBWDxnGpfDeYRpnxaBsc7eeM/2WLoD
vwTEI9NfEY++HYe6v3k9m0uIgOJ4ZieVOvPPnrCxiRYiJnEZAb+zjNzfXjXBsOURygzQJ9yT0OtN
vzb75Qx8HVXAh8zw4AzWRZMNkoAt/xnlKbCbyeCcSGEGMTljpjpXbbpVjgFi2tuazfBbta/1mO6h
rT6ufyvkI69mzkJykCirDivEwImeWtwKmnr4H7nLmz5awouViVwWLOzJRIV0dSEAmELGLG6Or9I+
vc2IX06BWVebPARm2E02VedsvB+zjqZwQAFFyXrMsArOwGuMuf9Z7gcwjEMu70YQiq6uSBHybauA
06SePBIkYCZeqCcPN0axwQDutyf6+wI8aQNprULtqadTU42HkYSz6/jvkcaIr9Hf8WH0zp+MeQBy
SHrWeegELoG/5WWq8TvWlXokQ3gsFtFUO861YALsFVENMQRXhMwdUGfALDHhdpx2+UNpbEFUOXcN
U6Zl4v5zyRHOBPrtI7Wm4hDV5JR+9FUr9p38FR0AUFvmZBf0qa/2tg0jhUsTtHM32ihleh7WrfXi
S/cufdsI2kbAr3sE6eCTm3k7MsDUs3FAnfhVTGbAmmj7fIgmpA7i5aQUGwqXF5o4z4Pk3/iNbb/V
d4KSuG/bsekuoA8xpXGQxSzoeNnGjr4BAeFYb7WVlo1YEssCchmbuFUe8fDKdZYLWbqslL5OsKhC
WB6Vxm3W5y2m2oFvEGeb9+D8Ocn3xkmoL4+HiLLBxAa1VKDZbzw9Akv0VaqWHO3TrqVmGcgscZCk
CBpcAha70ig5zbB2v6d0wcuHHmKw/+Loy0xZamfrs3CfqbcOjvrdERGJIJvdHnByn2yRKAse1qQq
gtY/nD+9YIaEDXs/W+WmWJMHZsdovXkGbITNDzN+XGZHfXO5UYY7fusu30SAr/96aEGPLQz2y0p0
p4N6SmxBNYg5fDGYwmvUO/dLZoqTvA5g5NWI2CusouXALvWjy7Yw88shPA+JonioLIQrjfv6mWzM
gL9ocHZcrY4kvsAWPwV9rZxJ4XJWPzaRW9jE2AVD6UbA1v9qDcQXosAuMZ13dH3U1VTVlkZdvBvR
+aMTpr6vOoxO4xtdbmqkIkyRxi1dXg6fN9b5ko8fLBZcuAQV832ecwHsDoGF7YZpjpRlA4opaRMO
KuGCFiH6rdSoAiTG8YchattOjtMusFayB+WORhnCFYyZ1mbEWjIPGHiKLrqnqnR8xJmwa8uEN4SC
rR1gJnzRJ24Hcj9NajJ06/XHap8T+jayJQeiPtD+akX5ENrPLLkkb26Tjla9QD5uT9ot4mmlZcEV
PyF5NzddcwThK7DmNZWkJeScgrfPmjpSieUm+2fbiUO1lbS0qlG1U74wRz4b4NICN5+LBW/uQkKp
O49+YAcSLRSFC7eIdjoaWnwb0/LzwWn7VhRcwoTaL+azQLwyjEcBxoPQuRTWSBPVz4zTnIvT5iq2
3mkZ4Ayf/mbUTb05ZV6bwHRwTKha0/hh7vCMZfJmS669yTgy1HyVczP7Ug0UXzw1s1t7ZOa84que
IscF7UJHvtA/6jsAD3G0DsUnNfbLGpl5akDsxRBSxZE5nqNN07NFfgd35Gqqu1BrygGmAIx58p+O
mecl/gR8njZgj14HrdGiDD2Bon9zUhKsTKFMDeZcPgeKOtkz/g7V3vwxkfe6qQKBMIgao7L+pSbg
/uPWRYx4E/WM7UhDZlDSi0VI+7SkSrCdSmZ71A+GLTevmAZpoZxq053E2ar5WmOx6wcwdufOx5SW
ggTK6OhYcsNO3AhOW8kZ+P2rdCg25ZocUYtwmWrtz1YEtESgH30U/DtA+Q2QVwk7RQq2ed2fR9be
Br0uUdWd6kOqNNgkT0ELPuoKUJ5DgBCdRquE2DJEbWOtm2dCPOW8deHXtye7YrdlwKV1BlJE9EAa
ESv2m5+GvJ51qiKY8homZtkrYUMYVo4BYPOffbVizIdAlrkblv4LtRA4Ram2zWSgdPqpN3J2MXRL
Czm9SK5CtNcdfu72zOukceXcnZAFTTT+T7iX6MXb1GwT2Dn9dZE7/RkdqVsOGoUfpvO0sZyrMCm2
HpCkB4X/aeODk51Twpx3XP8qsf+G+7JQcuZfdlxSOaGwD+3E+csaHYFomFto/xq1W6icvlIYl5Jm
Q+mWCASkq5Xpbfk1/JLfTN7cytCXEtnRER8OWU5qvpF6ancw1gzCbNB7iwDwkV4JHbcfoZJK+kEu
siBqdEQlCiT7ejpx7w0D5FhvBqz5bGNY/77lTZKWAQMBbbDuKysAMPkmXVGhfkpcLCI/d0ohQEGw
+dW7D5uPaErwHh92WJN/+2b2ieJW+QZOYwkHUZV9UWJjcSJDkqpXSa7mCrmgurEE1uoC1YTAJ2+6
c3qcbftBkkXiiUzF0hxgeBevvXfZJYY9bCUswoiTXQ9VixdRopRxHlIUtTkrBS5iNJPiDEx4aRpK
FQitO0OrJiabX0BjbM6hHwGrs+vMrtGxyrkFegZk5aXAH9wVZPV3sVOc2HOqsFhxK4J7uXBXH8oG
0ewOv5fAZclGVNjIB5QKz9+azy454hLLU8/knI4XbArdub5ESurjfO24nzK0hYsyms5TDwvimHsR
BVcTZF+T10FvMH6slyGMPY1EUJwvCDAYRWwDzIlQMtN4HxVk30D0yU5avZ7JSaITVRsbuLCDnsfj
WieJ2ALBuyXT5A+jrHbnGarW/OM5n/0fDVlyBBetLUWpyWqRvR+cx9LuzEbmDWLQIdOch3NA3B2m
a5nsxLACBNrWcbMx0qOR3zt9p80Efu4vCKNbAmYSWD1ez/YUTwg5/2fNG6P5EnlfDXZCjk3hGh6W
Z90KpTFS0QI5Yc6pR0AlV90Frhjmuoc79BTl8yfpYZ5T+aWS46fYFWNX/S/lG1Kk5EVU19F6w21F
3CWo21cbpY65ATNefghOoLvjjdRWBbDEBcWg2MbmQbFZuv63FdAJoKMvpFeiNM/FarCq4lBfMNy/
oONMZDin/B4v8Y+MbEL3Gsgl3cNu+7qhYdHZIz3tpZzcp5iWJkrdFFaEfEMUSSqwQ7yEOJgnhLPj
cRNI0rCUS70vnMrvHl7w10xG4OHtQ6Lz1/aWRGbagk5VsS96eTFvkupbzCNdutlotGQFqZf3skiV
sDCGEZLVZTYk0KYcvbrx08iRreagR5YddoU4qaywxcbMBS3Tcpnavp6d3guCYGtndnJggjm5ZfrT
LdGW+BIakHNlqZ6+mr5XiOTSqvGM38oUm/vocx6XwCdxHULsXcO7R8egxNcqA+QTW6keZ3+4ei9d
k60jzAwZp97dyTN2eETlcJAuUZ4rAj+ABlDLexyIXZd3LQZR/qguFHWoGyUrasJ8Toti1DVwYuLF
zs93w9dxtMgK26xtnNzVOO1rR0uhfumVbFY+gOOtQOGZcXCFs6BO91RGvpSl94x0EKF3keIKYPzW
xXqhquPLCvMyGKPpB2VPflwlqwEAXlRBZ9izA/mXwDMGLbAOTc0WmVipEU6kv7lYW+CuFWh5LZvU
fQmOZjTYDelB4zFPwxxD5/yHLpNd167loEAO+5C82DDUnZp9vzEzQcvL/MOhuYW8Lu00oQzqqcD7
xggWUU+sTMq1ih6cQHL9mkEO9a1cdDcNcK7ZkdTQ8o6QSIu0iIp7Pwk0Im5CSXqmQlTGk8On4AuJ
nXl6F1EXtUTLTnGJcoGRE5X6vFz5jkz5x8P6GOjyV1CEvK9CKQbL83Yho9rcQyrNJuB2H8JD5Edf
u6JDsABy8+M5CvdAcmevSb9hjTsMkB8ArURrC1zkCg9a//AatoJsjAVICEmAX5AWniuxfP06xi8L
Vh/mOEBVg+joD3lE49Es5dLgZ2VFvwggON2Mm/DBlro20fUk7fT8DN/93O7mawKnYE+pAnQHa5Ue
PbI10VBezG22E2cCmeMcMShBO11kfYEQtJiScfNy8xvAjKCObjaQEhn+wwwnLN0+ph4oRlOPDu7l
Hni1K1yg89WtECqZ8XqBEYAKYyx7wN6g9FKDrgF38TW1/0Dvh3OCeVlacas0oQDDcQiA+9Gkqp1C
41syzFRsaurgTu1AtU4bvAoQSg/o6CcJd/3qB84VcjmYdeglaXzYaqesS/toeIlN79Xjbnd9ecGI
54+8gAxz9RZABSq/nlg6++P8BFuSqZ7AzoFFhmbpSZ9S9mWm16ThfxugcLB2PiOtFNdv6iGKnjwn
yJB1c/IUVzV9YmFK4idEcfgYGPxvrdbf/EvmWh5mO7ncCvNmxuYRHCqnT+UFTtC/LuJ83hN2JuxF
nMJxtNCgjEHBclyMvt5bMc8m1+tsDNM+Is3NB985SMv3gM+UlsAg05MWVlf73sm9/kbaUd4eS2ef
59vmg52dAQx6Qh1KGTSI6AFz4rIl2kXc0nLuakPoTZ/QzWxeNFcG7xY+hBqQ5Kw5URdLCmNdb4HG
dC2H/m/myDUOUDvmbo+qE7NmgfEMrCxh0HLm7op53B23x3LbqrLsGPUhmLONvp4FiYey2K3orLaA
lw2ihbDstlKMvQ5iEdm4CfPp+rs4IcRUOhdaVqZCIE8gM5ig84COpbRQYS8rTLX4oN8die1WxEaz
oyJH8yQoWQo1UHPIrSwUSs3a3vOqbbVAdeK+pjbkEHn4EIHtDCUQCeEA+GGySllG0eptDKlKLqED
XiGxSCOnEqsDI/YIvVEX18S9AQzLB6uTGIwaQ/a6laP+pGmaTpgEHVUT5FT1FgQL+9zIEGZSvkBL
N7yD/CU7DjQ7okh+IjvDGpdCaThtL4Rh8u40O303RdckJfOYOsocbNpiWaorpYwclxCd/BFAhpsu
VePmUjvoe/bHUi61irJhWnb2QmvFl6rMugHZmllZCFs0e4L6M0lfWxeJKw1P4K5RC/QHIhDyPDio
99yzd0NDCelqcaNQSsBh/P12YwLqnjxuhpO/8M4dNgg0Hh2TWpDbKvy9FZM/bBa/+y+XnDao8R2s
19HXp67NIwZzEA/Iojxq7QjO9f4vBOZ0GIzYqw13R+wlB0KhaPa6TANsHkXCDfXDKXDwAFP7aPRI
aMIZxTpBv263V5tEW4zpsVAHlIq2oCZPRkF3jabrVsF/jobdmXhjWbzhdCgNiWjevwl6whechH3x
mlT9SR+54KWp2hP5F/WvKXsCsvsQAsiCCpvi0D1iFNjv+Y7rhEmDstHedYuIqTVpS3sP8If+F/uA
6GK58r3YhB7kHn3Cwe71Lgallhi5smfmeZe/Iwv4GhS6cp3B9D5gAFO9dJQCgAKyUxtUsnHNbiEJ
d/hI4j7iUmYZuHM4r/7V3jEVEM4DVOOwYrA7OOcLQCFz6PXLLrFoYPlIAjsPk6dGiEbwEe3PXimz
+Y/qGO8AFPCNT/kKpX4c5y5rR2zmXdATjjuoTxT0sUWzlUiudfBwEb/+9nxsep+rDDR0gUPeowPx
wb+d2xOxzFg8YbTsry6y9BcX4RQlZfGUPAlB0capCePTsLYKfASo2qGeafV5ROOU6H2VFifYQ1lN
tf7TmnYWuImw+WV8V2YOGTScDLGnOq8X7Wli3Tbk/DDywtyxejHGFJT9Oxm8sELOzPeeH3lKbiCG
2PR2lX8SEMKsazYmvhffLBYMdFQz72cTUl+mEcl8/qqtD9EWzPZ/Uc96/YVo+jHplhzodS6XBsjD
rZ3v35MpRL1yMaioRoCNk6UGK6SwecO8ItW1w81vij0+ybU42SvaFuGIaBsRYTtUD81Pu4tCzo1H
WV+poKepgYj51Xnj9kXMhXaeHUB5coKr5svD8xczFnnzv9xMQ1PN1PCN4FUuxZP7/X4ob/1NC58n
bI2LAdSXFRTIQOngqsfd/nQ7nHxGx++WDUL8pdDn9/1wpdWhXmTEj09WLjRnwwZG8ld1ks9VUJN3
z9Yj/W7IcN1oGFzOg2vkr/XEgxVba4Uk3XQJrSugiNrqmf81Licr3PuTvjFyx1i8UYWRiuJ9b7xd
ib1YFv2Ar2QHjHN0ndo5rsM47/9K4/9z27GQrgThX/HGdo3z5kiiMEj86ZglxSmNjal98x/IVGkL
Ee5mzuUT3Qk6XRMJ1Ozz8cL+8v4muMLVP++XrvosDNM1IcGrMJtf+KUAgUliMUK8bopRPkFpJxmF
Vt+w6ZFXpiTBy9vKktSmntO2Rqp2tQuDOEJVeuYpJCJh9fPTDpxwo5Uimay6NTnAGLLj9UoYYCaw
+joGzMSvS/gFkwxFx5CARNyqEhDky1qswut+u5uvMhx/62Y8cmNmEw5JOxLobqs7vBIinQQETrLc
rIBDfqp3Ht3euRE5zxoH/bl/x5zNUd7YFexjRr3oYkkM7DVVDuHcgFtIswn2kZv0r230V8EBpBE3
P9KOccim0gEfTXTYBea9R/c+Px2qP3jTFPZgG3zikDrSWkazXyTRnkJzqYVMJRCsh2DchCeoh+L1
UoNy0o9dZfxADsq1YNWi0gHI3hLba5W6i9W8npkSR4CjnAsQTV+KPIZ82jmGn7FcmtWdNceurSlx
kr2k7DWLDiWWuPjWoTs0SoaN0kuPus8Zg3vC9fsLLIqWIrhXXMm7ueR3jS6oPKic+kuOi7SYe+sr
guxnQdLI+6b4ZGRz+dtwpzkMqTrdY0GYpqHQSMtekXIqKUDuMFLbUeafyurQvAwVohNfyjvZ+lKl
lK5QtwvRm0q0KNKmaCNOPUsuhxVPUKIq9L58ELwmdrztBeWUOfxj/o3uVTU5SEPwmQHpXu5uRxA7
7IGE31B8AMKC94N5J5qQFeq7or35tXuIFtbPNiKTSiOd0oGIp60arXD0+/SjnbRQorS86XWUQDvn
B7CzrdHuXSib+xXAYw2P0AZozPYjlgXTN6+BSEIP5jB21utmriQliEJ5F/deCTyQufXLYQYkJXXq
ITUMVCEdrFuiVcZ9IGE6bQHJAVbdYvr3Fpd8B9AchKVhrrNJOo8yH2yBg3TlH4Ed7Ofz5TRNlTQF
qKzATr8IUzkQeV+wgVpIOrkx7rp1jWgOQAP56rV9jJTFhnyXyv/eqp5q8xCNJW8M9iVKioxTKsFg
4JOnYwLrz+bqKe/lX2ZxwMdtcJqrnkyp45PessWLKGMIMmXgJS0bojMAk59jc+3SIpatODdcktHd
8+AN4KNGrxTNL+Njz6SnV4QEA1G1iLFZksB+jRswuTPYBKLlqoyvvjLs/E3We86yT6p2H/ZGSkHE
t+7eZO70SI+dIGyJWlV+bFoJFxbBBA07n2mw60LH3Dj9EXxBjZWwl/Ld453b1ogdhhZoBI+T6+it
ZFpL4fpyPv/9qVoukFf40v2RRVtmLyonlnVu1IOBC5LdeGjebtrGlYUPP/Be34yXAz6fJm9txs4r
TqxPGjMJi17hNi3CMin3zEZ/t+rs3QYP725tuuKrpKWqoeys4lsVgMdiDEdd3HOtfsmjlx3qswCy
ZOqxzsyiVbFhX3FNH/9qIH6vYQlMiCVcBxrlu3950LyZrN9ct1eEx3QltsVaDi96DHiPe91WqJTE
SoTnGk3DBkEpgwmmGlEJi3Im8Lg9ZCpB5OED7RD57ueGKzjztXWUU8+ZL54Nu6MMSqE9bwo8nC9t
CSsYmqUTs+BFx7B8M1t3LaJ5TH3QgOELhK3IjccWrm98MpckxCiigNcDIk6KtPnYz7Dlg+bv1Bv8
aNAydzfUaC/BvRVrfm14h27ZBr9PauJMBEZxQYELJzFSqFJac0NSd/zpllW63NJ0vFWmQqtoib/j
k1QXppVy7eA+t5IsB3QZaSUsOVnHPFF9Jmnkv8db8IzYgmwTNa3GqFsunU52Ub/8LWyK5c5JI7T6
EyB9lq7Fjg18GtM+hmlEhNKPuvIVcGq2/BmJJNxoPC5L25jxzIDJtN9tNVQeh/90dZTFfRUUbQD3
Tz+d4Jk82ZkVDW/BgpA4qSwhgC+zg3WsTe6bW7tWDZaTEtLVblFR/5xq9RMK0+rJYhjtZM0BBHjI
YPauFqi2B2Lhjk9YoYssjK0UyFEym923n7sDu1jb85piIFEaAVioHAWVI9+HChGIrRVSMd06/Q0S
VRPLL4pzqrGpZPcXSb2cvbTpVQL7d7CrAzQGF9fakInzxUAK+32ks4tMj39bDD7SVrHS7xfL/y+t
ozAvEhE+MiaT484txxGzaZ4jUtMdM9b7bSSMSqoUGHTvH+ewV/CJmvvERLHMal+aFNXo/uh5sGHY
GFNMNrq2cGFo05YcLQDa+StnpfD3n6eBK2h3YXCEo6IiQWOk0agg7qcJOA7d6BLNWv6ZEOKXmEM2
wbhpRSIuk+jCco7ezbahjXyK9Sw2J3CcCUQKGNwWsNPagk83z72cw9Ob3hLUE7hX9qwPYK8dZRsW
4B0kGD8iY+9eDb7S0ZD9PJH4rJSw9JVT8z3a+U4XqznwPebO9B/+MA83Bwng0sF6gACyPLd4s+jP
fBCHBLczxluiDiz6fPaVHkBJwR4ldL7y9ktC6Cs5bT6rPKITi/wUBIOJ28vDz7s/72w8MSe/MBVE
47GL9edbpc6fUf7GAnV/cVo4kFYjUOIFEUOaArGdWVNZbkmhST0+K7ZI7p7NS1+5C5xZTBLsty3i
L5qHD1Cr5ijjTCkHzyRLSWzyV04tthK0Pwa9i0IlsTrsQs0nHLlK6Fsj8fPkeeNUiI+laPOtTQBG
9N/mC+F7rp9DJWQwF1Zg+qtLmSuWe3sjxKTbCvu9oPvLyWHxN/2cvBZ6qCNnbS3BV60XxZd4zc6e
aceGRqvgVBoHRZQhE649CXjOhKX6Cw8Ea4awWQR7ZvI3nWaPU9y4xH398Sge0Hki7w1VANqN40er
jOZlge2ICf1+KubTV+cgFwfi+icQ+04kWKC2ws+LkJmdeZ3tgWo1PC5A/XEn+jfGI7J8djIKE20p
YZjbr9kNe/R52OKFawTfwjYa+QiLj2ch7+nbCIqEfee8Skq+JiAJB+pcngXGGl5IXniw1XqFOsh9
kHwqN7XqaVvTGIo9M/+t2N8103Hx8wdFaYryIh/lS9dDfxk2NQI0rv8FYL8UdLitQDOQJEDfR92H
4NfMcM8kCSGmN0jxzHTuuwy5fzCk3nmbmXP+/SaPHX0Q5zIL7cGlsuKM0WJVH/Qk7VPH9dHQe9FV
gVwznUAqx4otGQkLUbSP0g5zxGtFadxxbeSDTykUhtuWLHbgTjXiAgGlci2ONLPwGKvgx6XztZXd
CwKN+gaXFqHkGYQyyBzS5bE1P4lcSlyhLFm1n+HmDOYDUQvL8hggv7jobuudnCdGsUeFXJZhIWV8
VEJGZ7aKbHXlH+BjEy1zGALqphI3BizmZBgDNPHsBpytrKJp1AsYHCL3xtBnf2vLatft2DzhoC3k
MkPt0hSmDbmID4Q+w8ijwzNLFBKbWxJRbxRTAom96BeqNZ0b8JJJ2OgllWoobBPz+K3NLUbmAoa9
785G242f78/E0XjRK5V1Vku/Ue2D4umB3MllYLa3JgYEZkvZQsn0QfmvCM9raqI+GXafEkUqCvCY
l6OZrq+6bZjSyqTZgVoPWwm6MbaOj1d8pfX2RefCkyaVq4TNpKM9bk2GTzJi6HnXzn1Veled2TSs
3N/i/pOsQ7849IhQE6LtHb3gdcqLG1E4W6gWwwxH21oA+1fwct2Xu/8cfg3XwLkfiLlBQAcxO7e3
SufzG16Mgfhh4C4yn9SzEqZVRyaR63zog7ZoOq6Y7RAGLbaW2oIreZGv3/fhBIowCmk0IR/sINnJ
RgXA1UluHl/fwTVz939I9SWAb7Qm+5UxZPJJE9/8+k6ZiBcYUyRqauXG6i/tyT60erhOtRuLwG2y
pdXo/+EFCJNtOdrzhMFcLeHBU5xEOuBFOtkvC7D+pBz77e5pulkxB/Xx61ukkgUn+wpP10jV93Xi
irvyCzLAJBTNyprr1tCgFoKAFXmloIqSzVA9nPBM4o23Fs2tlGhE4XdvnbGV2vCe/mDwT5bDhXnv
TO99aG7zT2pG9DJilPvbdO8bexPuOpEkbpdGtyHixMtVz8NtKrKgwehV747VDge8FCBmA+5wtkyl
UZ/wqKbk3xHFuxZRJ3NswNmBTi2mZufeI2VGUaBnsC3jnMcANi68E4NmBJGZJ5SnG8DuJMtqwJ2S
3OFVZbab+yeDSUJTy/WaK40xt3oHWIjStpFgS2LfGjO06guJAeLq95/dAODPBC5oiRAVspKe8QT8
lqapAIVqJRnWXBC4/3PTf+Efoq8xznPWtFibdpRx9mWJ3OHHQPCI8ydOnpRBVC2w5Cz2w5SPgvNb
ndQotCLk+cTJKiCRGDLyAwtszxF/t13kM1cVBELK79vNtpFTaebhfs/0m/OfMpy78bT8TPlZR4dv
i05ET/d+EFK+/THtoe5jlPH6Asbt3IrkMxvVtAHJyMl/abiX7qUXLc1rGac9656gx21z0S8TCGNn
0l/2DUHxpREKXdyD1tT3jyr/06sKAIdbORoR8rg2tIagG2b+QbOrH+omvsuS7oV+3js3/W+LSL2l
R1WAAw6muoPkXvx2jt6sygvKnVzMWUGgO2BG2VWCxVclhNv6BGF3cIofsWS8PNPcgaia7KQ6s64M
VHohpESLEBQvPvXasomkFzRVaKl/lz1nCyZsR1F5fGlKg/Ywh7GacFv85XIuxQS/pLJj/SaMOJmx
cXWueJZcHwu1dTZinnSp9uWFxE2a+2/fhUR+lXbfuFd4nD1sq1lWbf8t21E7RWI8k9LKf4kif9G/
0c6gWjzNV8HS16z/GKz2FU8+d6hON+1Ac2R/AIL3fah5cE0bH+4vVb0t2JJockRArS0n3jy7pXnx
v20dfB+qWMRia/NVpwAOxrVHyny5eURyoP/DqPjpVYluGAWFQq9JKZismfPEVvFES0YzgZq7stUO
717MNly8m+2QomFeBmmj6BCgE74MWjWNBqe6cdEFTzQVvfHSLFxXtMdprwj3rBAIpMngLWKqG3QS
FTYh8iWAAAiLyYcrKNkbIyKPYW2ltKBXpxhd6jMqmquDgePnK6+993IH33xaJO3adzNHcUmdOEmw
Go0UvnfVPDa1gH2kunOQ1AmiplKYkBrsrrZraN66Lrvggn2zHEypvJmw67/IwcNOvfUeNrTeL2nf
pLtEJyLn/iDxFZ6Cb3A+2X1MsBPRvt6NEyROJvVaJsyzXbXRv09VJ2KWRTeNTE9s1h7JGIm5vplz
B3hfgSFrvHnatuk50bvWcMsvrkh/C+b9EIdJjrUruMFBQpTSdjDrqCsRI7yFfiRihDXNC3m3mdEA
XaRoTBDmJXhzCbZoEv4J9GrvIcW0rxKPQ1+E3Mu6By9KZ4M/o9QZyj5ENNyRp4ZyzR7q7dOrIwfk
YbowZdSsXJxQxGGKflyHhGgHarn9K+O2uDCHFb8cQOgsy+FxC/qrrOAb09hkCX5C+72aCeLxZ2vm
hmq2J6mauJyyxlZwzwLOU9L7n85SXzFPzGJ0d5clTs3n6X4pQhHWIJnx0/Fg3zHRF640MMfEUtWR
lmOQfpZcWH2rwklwyiMaQxOfF7bFSUGN1CIudwjy3bJLM91uZczCplxKJaz3G1XKnQnU7tsg1fH0
RXRCBwqX73wkpo8B6IehaRS6NWULMLg5H9QSPURaJWTMOge7AZXdBoRGJhjgJwLeyUIk2y4T2Q7J
5JCVdBk/02cePDNE+Klu9S0SQs2x//wXBuvrdWtLl4OktdQEyl8nKJuO4ZSDU9J5+2f6llYPsYpx
lQqhSKyJBUP5lY2De8jqkodsRPizMMvRznWxSnNsIwRHwbxS3I7vzfKzSnf4hf+/O8sjmnh8mSYQ
gwADYKxcnGngVrMuNy1LDJZyCY4Pre6JfWec2uY02OZEVmcdMtikEniJt5flQLsrmxSgXevaTkqA
7cJwno785Qwssd0yxjDDxtaOQLE7mm3nrCu7OEuu2KJlwSDIz0YSfCsMWhHuExiU6ethRxZ+1Qsa
BiWIlnlcrNtVjIK7WyCNU8RO9otJQMAwnTqjkgA2YzeP3+c40Ifh8cw+tapZsy8V55hEJSTiI0+5
NDavytGs9AQZF0ufpwBLW4pfbDb5rfgshtUyGopIpUnr9SV0sVU8sWQYvPXJpGQcWLGrvxx00mI4
qrVz+AbIvgRo/Jt7t2mrMWozE9hmEQxLjmLl9JHMsLqN89Y3PXnyq4kcmCtB6o/wxQglqDKq4ScP
jRLBgNuz/gqXiiMUnyJtl/HQJxjx8XaqKxSBBkdetecBcsUVGvjzmxlC2mbpQ91+w6nlh2owLcSG
YrgW3qEmVS3dBZ16P5ob2QjsUm5W05ah2do4PV8VseigGpekvl7pigLGiZ3CH2ElPO+V67QPj4M1
/aotn7fVcXjCQ5QMRsfUVgLxG7Q2HryIUbuTOl/+DzixDpKgAg+80HpuOSReXLUtRD9sPOeYykUf
QDDFsiCFtvrEUCIeC55lS/ZmCJjzSidTkd5Zb/YWWHItbGethIOl8Wq5gQb5yEUzgKSv+VDKyUQt
8aYMJ2ZOiJj0BJggsPMHMy5At8bOaQPo5XnUssZ08uQXD5VSeb4XIMGwdnLnWevxQQWN8EKkh+nU
O72UzD3EVYWK78d418II8ttoJsQfKMestraDn0nv4L/26MeNnlEjZuwl3QmtiV+9/Dn3kKmaPLek
YiNPUMMIcXrb+TdD1d8D6kk+UXqZAex5J0dX1J0HWet1YHhSLjls/bcXKXjoTH4eESLwwCSqppiU
t3pF32VegxbMEFJLkvoqTSTTPtagjbryFWKf9PrO/QBy+qYFXD62XgRxobkU6Q+N3eSVDDyX9O4R
7WkzFDSj47329Eb15aT+UG8u8HPDjSwMjd+TVY9gs7mV0iLvDmUXNBC2Q0tsDJ+3YgJHwsILEL3U
nWw7Iso4C1OKsqyNLUq8YrnRk3OWyAncI8tNBYbzWN9z1IS5efvU+vla6GKL3FC9Dh98ogG6J4gA
AFWEKGsEl6AeVzi1YKyQG5QH86fxepdNXaQV2TTtKMS7pnZydj4XxWOahX2kvzblL0NV4IOLl63h
wT018uW61H6CDBXjGL7LOAHA5kNzs+Xf59lJG7qG8UjBrNyaTcfnhyPWFLg8FmLMhDPgBgSXjita
RF8eO3lnkWTR3P4agCcYSF1SmK239maiIVZUQTKWK/X2gjmw2uw2JK4cImhbyrr9+fRWwCF4Qw76
trQ25UUaDQu3r+I4wP5vrgOdsTpGZ+liFO5Uojr9F3ZGOQg89Q0nedoNHCT8txOOoG9WBrZ+LfVx
7iSvI/N/0OaAiZEuRrIbS1SWNI/sE/k/W0lYQY+WCfgc3qDy5aiprFyE19ZcXqqATRfhqujr1dZq
zJKl7ZOCY4QkuWK0g/g2hWDqzE9IYTdF4tC8bi60BPfyBrv4SDGh2W4s5yP1TZg0JePybdEFFEXv
ytH+U76g9y5BkuI7rVFNLFauhU3Xe5RZP5nUDCdoE7qSp11+ZCBL3BIPcKx+IbI1IgDtBPF5r57E
ldf5By8eb9LcqHz1XPR3Yqg5/3fQPMjvth4okAHztw1mcPLAqutPxrz/1NtqVxv2v2C1SHqDoGws
QIX8onQGCUGdbJV9x2PMMnev2vmKAZsuW4/6hCnu0Ip7C8E4S4YDtPBJ3ZEwez/6vzd1oWdifWqV
Tj+tRRiNh+aECsGfOQyn+0JJObl/YRN6AecvVhHJ2HuZnBtc2RzsUwJS27hzYSvoDwO6dvDEecl+
G5KYUtQSWxYG+Wn/Q/NLrZrhb3W/Ffd63U69OjKfJolutfJyDVNtcS9Cg0JdG5yhZI5yMP+xo1Q/
qJBaOj9KVG5qSdWkAAwxAbfv5A2b/ponTEgzQW+BPCYeettpgX8j8wk0IrHCeIkkD7kt3BxuabLK
TFeVruHOMp+MQIwpwc469JafZ+x1FtKILGqTzAN6iTKy0CqQMQ7LTdDLuN50PqEmcHdB9RYTKfN9
KWkHOORY6Vb6yAQ6vZmrpff82AkbUCqFGDD0DHsuIvU76SaMi8e7JcRvBFzHHw5ZVsKq6y4yn90b
iYcmaMQQQ2L1WQ6yRMeitzdqcCURY8mP7FVpXwY+hNO4kH6+UPxwodcQMjHa+zoUSL/2YKO9Ge7L
ANiH+OJc6q81vKo6sIywz9fb7q9h2XH0VuaziTGaQIEH7jxPXXtOPl6RqRKSWzzDIRjws9EB2Rzt
sCIlp4+HHfB60/KSA+f/fa24Q7sCCSwoVinJ74+5x4kernClgBO8UkNGchvorK1pzKhq55ybN67D
aErTM/jXXo3Ef2VktmP3QVF1nsQPnJk32FblW5GCbGpHFAUl6tuUKLodAqznQchC+CxaorOosV5X
lk7di4ScRiXIR6CHBTp+iTe0DFJrm+a7+KUluXRM2/uYhaTxRQPfA6OYy/GoJce2l1G+xye/QVuL
eOwPzX7DdUiyf8+DkjAJA+bsKQk3rw16K5+pOUa443he9NTs1C5QIUyC/AFonvScYmYjpz+HE/eM
ai9c6hSqxX5avTf+/gsuDmz475QIvOay4mFehbRQxrWD6U4B0S4asJ28V8My65qhxm6LU+wMryOl
772a2tejBmfyAjOSA4aTNkD51r704Yp8IhxEN2HpqPgAutZLUWp+SytWkDtOd37kyfRU7NTb3x/0
9nWyS2RjOmZo6DNpnyde/U/DmlJKw2IQK1ah3kP+kwS7bUo/wej8YlQICxuwhDwZl7OV6DGEsqL8
WV6cBSup2dyTx+oCEhwHUNQe8Uv0pq1a+xQvcLqEWnS78H1/A3itU42F+KRATblOlfdRtwV+GDfi
CyWL62NmV2nDD6RqWrNo5d18Q+g7fJ4cg+iWHldIyTuQXfgwz5D5RU3ECIL//9XFT80hrLSCc+br
pvxuYFksrOkbh1ECwLErqBZ16iGCab99Z/zUs/GosLxFwL29PPIbtQZXeOxADIH5YQGiBvcb9/b8
CF+igEON85IDzscc1Hu42m89DuQSZEbbq+UhgCgeJuN9XXzXbh22lMoQe92jaXQOVPHUT2FFH/BP
28FzAKXC+S+rgq6pNeuE7IamLVHIlJOEwBIgWVL42BME2fDmlBqYy4gWCOpObffdik9jN1/OA710
SXXmsHgpCRcaqqR5W/xQlQmszGltH3XOIh6N4yhZ42COCNqB8k2QUufrRBx+40BQAGZEfvxxTYnH
nZZld64sy2f7YuNFe9fPp9ilOp7oD39b3EsH5nE3+Ir6tJzIMUtXpzv9Xd2NS+cTIYZrY3bu8bmg
2wJyssiP55tCOkhqJCsmwfBopKOU6gafjTxB/ALEmSa9J/QCaSFveq+ovGYpA6ktWvIcytuhZxQ1
t45W3ugYNQjAgDgyLTZwxNwqQNSNdLgi3k3OboLOzUqh0MC+4uA2633iTu7fIj+/FoAMkXZ6QekM
LyqQleSER7CvmkT/tW/W0gAJBMqFCerU6uvnm7o7reV6vxkivBcKVUgmnVCKPloL6MAGgD/JzvaE
kba3fahlE0b0mYw4B6Zi22rTV//vaF6xvBXg/s4cvyMwrqOi+/DsSgvikQa/NZ3Mhd5dpXyQbzkG
GvG3/FCO5z9Dfdxg1kapBOEAwpi3K8K9O34DetKjyx31c1aZA0yJmC5VSr/vj+8yJeNXx0+OISVU
rPbVgRvxGmfANB3hGGcHCuc4eIjk0hq17uqYiTOeVy/7XXktWD8xJByfNJ7tbTwdULZ/p6xjnst6
20rivJWPIl+etD9OeUcCGqEvwXeKbOfZhtjLX6Zey79wwzSvLXP/VbZreq+ZCtfQkPpqAwBjjs7h
5Ewzfuk/DdWzllN9TwK8BhQL+r74FWXS3v00nbbL9GGaDp6pTlavkgeVAat2YMRh8yWFJndwrqs5
dsTLMElGzqEH+AnRMPkTmO9RwKcfPaG7TBdsXMUnYXxkwvP8U9Lm/MB8MJn7iIsFpQJnZo8zdmt9
1U+kYb4oLowjsB7UZdiSeS8WaYAWQjTRpAoaD8wWSgKnmzhUogTGH8a+w7eN/ovHxgugldbBc62H
aofz1+X3862i6A2tP0VBcJd0U8FrbRgIhwpYKTTeJjN9jmEAcMqePx0xd6nAsgiUHNrBwOPxxK1h
gBBSOq0OmsjGwQCV0jRSFnHDnn7aLi5bOgl9ZQ2TrrybGq3F6hOu0FeKK2XiTQANuhPj3iibPXXC
zIESXXqyMjbEIx5k730F9Y2RDEnH0G7Ut4cdIAyj2JGn35I6g9jleW7KPhOJmGJdrt8LSIfOYmOu
K+bpIpvboLjQtZrT5tdRao2iPxRnVrkI+W+wc8hq/1EuApmKE9FXz6TVbtmA3F4Us9FA1QAG2BB0
H+EFWOB/IU9LpfOMPwC/G3cH24PHT1R2GoWJnGuY6bnf89YSbonF7Te/xAwbd7xuXmDTbvu/LIhs
FeOAQLhuZJeNMicOAXhwb7DW3TFCMuLGVN7w5bslEMaqUSA4rifyKP4HoFv5HU1905woJlTnkHFL
wd/EfKhb4p03l4/h3NjXFwhd3kp1pv0P7gGEj5PYvUFFaCWxJ52SUiBi2ZL/X6+DowflzcnX3bMj
6vKZVSQRl7Fvpu5USdcFiBfzvJ9u1GjEFvgcP0nOkzIqq+tzfqHo4nXMlmJzVjy/Q0o6V5jWOMC8
9xmOR8q/HZ75C2E90jU4flSmSMw26OVW1YEe1NW213AgntUsLxG2sgrvK/f8UCKnq7fBV2VpIEx/
ZUJfWPkGjOAGGkTnt9bRSDT3F0TyNJCmWA2nh6wiQdQ+ey14/otp7ll6vLhBUPGxbSUwkGe78DcQ
57Ivp19QKyjeVRhSrnDtAk07WaSRKf1eW8831pyrHtEONcIqEM03xhPe7Bv8Nl0tUgR+13voK8dc
CEM4WTPzYfRCFsHzAJ/ujjOOjCz97pxWNMVTrE/9l/L2UPc6YeEQqrYUbWdcZBqPw6cdBmXaRNqK
zn8VKgS8hukMX/j3kTEK+3zFcpdDKePR4V/BFt7xBRre26JK+41WXgkDlrN9PJSVF21ra18g8RSz
9ddTUeZiom5A3T+BHOX6JQAI0sJGd2tW8joknRZ1MM/k7igAkAB6XZfhgQq2lKWWd9hUom23AbmX
2ADqd9MGpREvM6LfEyL03o/YdG6vvaYLKniti9GfOiUgNPVcER5vElnajiOMcUevJwQXk+knq3gT
PlMl7NhIGOUrpnMFJZRJoWu9J7yABEqunCKKJa/wvij6QI9vMkYAU35lbcLDp7CxvZ0C8owA+Y1E
kYBCgEgpAyI9bNNohuMfkC6RfD9Qp+3+tMhqW9CHTvfC7ok0kOGD0j19xtuPoNcIgcJ+C8q+G2wm
+ui3bH8jySclriyX8BAP9osxVuytfMO/RFfmFVUbPJFWqKN1IjQTUGhkf5dA1uC0WwIDsiKdX1qm
cpvj8DKTTwS9zR9YdFgD8AbGBRLA/IPXqTK1PSHqZ8sJJ9dLPu1n4QdrpWWPPcOu9Ix7i4XyRGnb
HgvIctaUiAv+umS+St+P5p3DreOkY2DGAIgDtJ4zUcKKwt3Q/mzdLQ+TPzidpUBjFyFYLa0tnWKb
2LRM5SygM/xVCUqBcXGn2uM4x8NiqgxXOgHO6knhIGvcRBs5NSm0NqsrwdfEmZiDKU1t5ncT3Nve
k55iBeyw9zUBzaqgP2mDQy0mjDTXK0vIFC1q27AnL9VGt1NirDQlgCmuytyxE13M5Nx6msh/E0Cl
Gq0lCUug7BYkpmaiNSwb9bRnw5mKx/ZxJ/6ikTmp+RqHAmkvYnnwW1ws2i/hGC4l+VZeW906Wz3a
VSVZTZyyJGufSoGPRdnsRSlHnejDoKjbPryJU3RHz2oOFXuOXAxYD+FKEsiKcNkJZh9q6A0p4/TB
RlhYVSPTBLTIALxW+7FqjnDbDtwKxxJs+Ebh1US1m6Ty0aBFQjuXUvfxINHXrUDOpTVkpZcDdlny
SxjIdF3fqojQb+dM9YH/HWS6hc37m3uf0esgW5TLMfaEYwH3LgelR1gHBsgLQe8bp7m+iF0Ll/6D
iAzu0bJsbLm0RK8BpwOCmk1LxCI8PSPGy2nlbkFh2EBwHEf0X/DbWFqkbfT3vin8gxJpNdFtNVBr
SIsMyFCfJ5T1LRvL/bPoITPc6ddeqj/EjcjOgVRQeWfXP5WTX1Azh/LoNFNQZDJfZjlFoDjY2BHG
wCWzQHah3Zfn6QXUF9uwD/eQKU3u5ggyrWRrWySFZpj2e+t5S0unLKsIa262qk+4RB+1Be1TLmxD
Zn+RFuB+X26OsHOfxJ1teYTMo6fx+rrgmWEI5TP8gSBd60RflNDqpt2cIpNSmmnu7y9wLKQe0QYU
P2XtgVXW91nkJfX8Gq6X60QbfWTDrQn8zikUDVVbRvMqmKLlrONvqEKnjJpI4Qz267iUpnpduSL4
EwSyuKLjM6EpAJJ0Dn7TTfxBD13yiQclmDeeFM/VpjiOKpa08vwhBG6PkmoP6NPvykIoOJX8muDZ
obEEuxV5vTyEO80sTE60ZnLuvuQuxXRT5dezZmPXpqmZxMNCXA9Lh2o3Flier3JOdlxwTelq7zIo
94YuKgRpzYZzEqO929WWlHN+k5RiiH753hL2TF6sZn7FUgc3lvLaZKbE/xiJ6XytIX3paMQhsQT3
CJJ85uqR1gWGZZriuzk+QJQ6RspGVp4u4khIPPGhJvoEFvPifK2VlAx44ghA/W8w2TArRb6IrNdS
tKzQVDG9iHFG+k+U2FlUWL2DYDTOo+vLJS/Bsne12rcicoJmlIRdg2jLuTUwQ4ph52IHIR0PJsMu
swNQFJQRLUoN9wD0xDGwivk2mcWh9HolOeJ9VwqR2HyHwpbdIERpJpEIQWedevguIBv1aOWO69lU
ccEV87VrkhAw9mz1ZuKLC0S1ksBkXeMZvbm6Gpok2tGB9PiWjVmXogkohHmBkTmflwfM5iLRdcb6
Jneaj7IjalFpHzvCdD6WWQfyYmKlMPQbqyDH0fayvYz/xaCtYQ1VmeypkaJFeMBopbwW9PL8g+Jj
mh6u1s5FbM/gnZV7zBTuGRem47V3IwVU6lztiskdx+x/xkn6ettjtq+SpqupybRRbFlWfmoP4an+
FJJJpDtcNovIVmPKlFKItEl34X68MxkkxzV3DyuMUpXre40s5bfraOphBjsONxtdih0QzI5CWhp8
xLYxn1hE23Lp50LH1e3RGVxJzXE7jl7PxbUkAgLkdCAG+pfYerrZ1s5aMRzBl4FH4BNJD8vpozLP
XENJWvRDL+z4yutMqblRL4grUlf6xFm3lWIoKO+lM0b6hyCVyQ88EpEt49NrVx9Vvw3W+XEsx1Fq
iJF7a2DWshiws7H9d32MKYAwdrBDDr5C2BOy7lvnS5YszbMf5EPTcncZn9m8cY6QcH8wV6vK7zMh
Kz6fiWVKea98flr7NNF/0vW9KaK9Dh3ZjUJ/Pc7ua/+kdsxEpIzbyONj622wieorSR/ARTo3IL53
nm9NBmvh1pACnrTxckCGpIQzX54BLdUOgFiOYKvd/ElpOAHv2kVUyRHZN9MhtY96nGQUk+nx2D+M
n7FLb/xf3n9AKnAeaXcTy7OE7i9eCN3XExegWIJ/bp6rSXcl+FbxQkVPqWEf5QHEnMqIQRjDZI0B
NrPRapz1mjDacjRe6T3VM5W8D+AgTAeN888upXliPpXLUHp4pFDQgfM6nBip9xmWpXbsPxBKcVHf
5C/Udfk5+3oK2ouUw3GnxUvhKBILnSP7tXGCnSDOffx7mj88rPossdvJXlOkjNNQom3XAh44aCH0
e0nmSvxDnWWlLMcTs4tGGP8JXnH0hVX7m+p34R+kARUjEbW97UY0vnC1K0rUYvjT8S4RnurCsSUY
yaVJZx3xAAsYzaD5ZTMSSiDMsjNhasMEoi6m8wfTMxOmav0yUuw3eF6oLJ+TNPsGWTGXEJCN/7ZL
9kjcIgxE5BywuRW3oHDpxLX4qXe4DNnI9ykiQmWRp8hGJoUGlnL0Vg7YTa9fI9DAVD9XwqfSZghV
ey/egIEzA2FnyIdDTot986BmQEGa1XpPdpDqJSBHNetGJuD3dM8mQ/3uRhzEnkviSxFPZUEtrBny
AmeSgcRNTenVCamDodK7RXqOA0Hi0ixQbfhS8ca8QdqwD0SYt3vWAm/6h+IptQRP3XduuO1EBn/8
ifn/5FjRHjDIwlSPOfAqqzF+qYoRVYVBowkRNHpr7cYtsDTOxv0MZtpUImoZq0CXL12wMH8nmli3
x1eBJUGE4vkT8FiDFOzIwppwiiK134yhulYuna7x/YOOQm7E8VBCEVm2HmStL+nxTppBO0oN0IW/
RavbMYQwcehzXCL0dyozC2klQhhCmmqTa1ZCnCu0zP+mqTKRmV0them09mgQ74qAKWdy1c2adG4Y
knHlqnuRezuyBILleYAikficXGeGWpvDzObqhB3HO4IiXFREU3wCKroPHtapH+ggzZjtmn+8DQ1D
33kLv0hmPmd+d2VYEu5tUrOrmJfdt/PTA7PzCrrEcQ3p0nQ5pSizN2QEP7Y5AxFVsTtw0aQ/J/kb
wphqaodTweAgSngErYI5QfqUeQUK4Q0z4Ta74/giDcGhWrIN1MGgcYAiqUw1fhwRf/V8ofs2Bt72
pa+gGLw5FEUC5D0RVjj7f94qz/gPbOBfHUHoNZbpFoQJGS+cbJfhqG7wY2XLMcfT/FaMMAWOG9fh
Hic5Bn9ZtKx99gQPjWxFoTAynyS48PJsJKdibbIU68sIfpKysnmTbql6j/grI2oBzftrIa0ExvjA
4zOANk15xuxZ/ZtTH/mRPgkE2Hj1tds15CzxBZ2yFkFoWG454LCxg4OgfVZ+EQiLBu5lAT82+mY7
zmvbHu0rsbvdi8xABLzX/j7q1+lc94yADLc8M81fik4WVx/twl36MZedtPRNExNhsfZwHAHZ5iej
kr7bMk41U9YPr+cDeClE7VTE3M4r8/UXjGqHZcfZTtTEJQitM7U7htrExzV0jA9AYA+/zYK/1yoI
Q1VmPj5yGyM90Bd7WTBscX2Ee1zdSIq8EzGv6nmgkoMD9mH5EdXCiFBAsudTkXDfzsXZu5sJNrYd
eCnHI60TUMGdpPAqh4apRGL03BeiH+h7i7gULKCnUx2VrTHaZFABCUAR3bx94uJzdvJxvQOGS3bH
NU3dkwoCcEMS76JgrDaSIRRa5DJmdNRNQO6gjApVIc1dEjVP9IEjkyBMJQJv4KnKToHbHF8mCRbl
mWSAL/m5pzjCOC9QbNYa7Qw6QvqS3E/P/7KCJdUM4c6lyKjMsdLD6/wK12H+SZ6rnokc5BxBHLlc
eraTw+HloJjzMUknDIzA85/2Bg+jshnPO23Un6L44Lb6j7qcw+NH0Zw6knizLDhCsLZicFl0tDdp
CecyKtzsNgcKwFubJ97QWgpSOomSHoZejHjkEYRDq1C44gU9P//xaoU+khRm1j783gn06CrbsyD1
YiFnw8r7pQuAQiADBIm17N2OKPzRBQIfh4i0nUJcmdIAZMlBj3UNMHfxESbb6u6XNLfN/hTuwSYn
Sm7QSpT/WjCPCmk/xKNK+fZ/Al0ikpZMSfd8ioXcuECqTfmvYRy393bolc+8fHapf6daZA3GeOEW
u2FIIkQlBDet29Pw2cDguZzVBmOzdvCP6rVyaMr5iWAT2QrjMc7iWTYn/ZaYcUKRFyb/76novvEX
pZjYd7EJkxaES9hm0cKjpH8RGf+dodw5e23iMUx/1rDJ2gk83bXKwdHdJmeZ7v+gnMoXlHeZ8+o4
SRAj2dOjO1bAQq6Yuizk/8SIkRfjm/wTr39sjFTC3YqjIe2C6YCN4ueGAw9gMF2NIfzXRX5At98I
7EOabbbA2B1oU3Rw7itavxt9YqdGbg2daGhPgAyKUPKolYWpjPtJGg+RpSeGZHp5eHCdwHseaH82
7z25/EfuhVkLvD3cVJF1t6+lU0boozh//yvO59NA50T1jQ31EUZpVURhBTk0ZEKU8D3AAyxIZPzJ
+sLyt1OplNpxdUsMRNpmHPgaCwPFktR2qBcW7IiV6ueMwWTbCuT52Geb6N9fjYK1TD6i+b02Uwsl
GS9dorZAFvb6a5FtqYUS3QuMPSyVc1M25vQA4TZJkNEsTUMrn57iQC35ZkPnKwwQF9rxYSOoeRuu
DEyzHv7cH573pXwBYlA40IURI0aCVxwNiuS8hzw3RJL8WCkSnqxuPTlcwVebVRx9GxBrtkhjqlyf
JwmdgWwJEcYQZnTNzaf2hWi4HEYLxgM8sBc1VDl49cpFtb2bo4T+AnrxMQKq+jobUrS9v+JVTfqo
P7bd7ZEr7v/7oO/moXk89XnTJUqqpibBHN5aRvEQnICu3T5iiFugVZLqsoOn2e4yQhb3T6SiLxV4
Zsl+mFXgthU/cH9uBS8ffjZwlHBVyOdrauWNzWrcGQ2VhAzmmEX4ASxaUKFs9DyTjDOVnVWmQK73
acBgVW4LR1VHGH9sksEZ5Ocu/rQ4ZYzPUpJIUs5YiB2PMsUhBGbGzmpbVz5mEUSle6a6eFnnA21l
Lg80dmEGq0OMC3i4E7fwzz6SorVIGnDEeJWV2LhFCBwwDuSX5opn+Ps5wjIC+rQiDFukl5H6ny+P
mc2SNe8vSoes4eQGgBDiSlLo0EoJnIOEzi4ydqeFGjf1+qM0EmhAQQY3p7FoDdynRfNfRAcd82Dx
LjJWPoTBts7HrwgkOkgumFyjBtq8bygGiC1yOvJO8rhKMHKskCRPSELGesW9pObIVuvbOMJLVdnV
pP+m9wNIR7QSa0QHiT5ZOhYZapcaLyI5rgJcoPob7n/9hFm4UAp1hK9MgMuORcgTTGdl3SkilCZF
/I4U1rLNPzss18JalMj7Shsm5JGh9Y4jlEf6+wVHb7bGEmoZ13q3GkW1QMtjTVCiBRxgB9zEeLTH
Sjy9ml/VhgQzO0BzQTnkucuRjclrk/sLcNMJ1fLiu62yg83CCsDoiA65PMgBEel5iKFeCK/7QtnH
KWuM44kuqtZEvsGlRTZsUk3g9060XLZQE7x7vsGL+ukBiwsQdnGwYy07z+SX1+Nt4cloCkzgxOWo
eJfCObrgE0vazIYq6xGDoxEkIQrFRx5IWZOgohh9lZHv8mVGRQzHl6HT38ZXsjxid/y65ACgex/W
TVMjx5kugmby2eRvSMAjogCCYaP7eeluptPQ6PCLHUV9zMleief5i+l30Ch1IexZcplF/zhO8i0O
WK/97E9SSwU2F0YlFzgGmlR1MfSBGRZTfeh9C2r0ufLEGkTICJUtXk6tOu+UxhYKKwsOe58roXum
ov844AGi8zVVCJdwVpYSrdnYF1ncJ4IP1oON7kuH+ZlOnolbrWS4tg1n+v6csu38OiytkB/RHJnj
MDJKRQ7hABT93wcmF4Taj6gRFO8m0wWANuRhMjXvSkEsMk9BgyQY2eJr+yc5pCFtd858sC5crQZC
/zArSQbMJpDMmwU8afVoxRA4Je3sSS8PQjkT0y3kn/fDx3VAkP0d+QZrkyPGXBTUedZF3SiXT1l9
4XxWbJQKpFjUAhOXBtpGYtLqrda9DlhMX3DQ3UL+466wK+UqFzXLGeKbHROm+3PfhgiZzwtdrubW
TXK4iUyH3G63+XGvLOr6oYP5kmdV+yuv+ScxtXjl3SpU/48sQzVPbFvhonaXeaYRd7NpdvSQhXOs
PUP+OoPL2Ihsry/7wlNPilpw9EwqfPLpWrECdo6lHFoYVxNkTsVgFkbrjDMrRd7Db9fpCaojauQe
CvAwtCNJ2WVPjIVl2Efmv7C89mhxDNkrnRHqz6giC2OvmUNx9cBknjlftoEQC2TM9Mc6s17H/Idv
MfRxXJ1mZEy/hO+PwOxCiVtLR7AHDg/mMGk0fchz+S0dZSww2YdHY9k2ID8V9ilZj7qwTJEDQdDG
W3j4Dej/PwcaB1j8E2padIGoZd2O/FVBRCr2G3zWitXS/SAiGxg/1tMMA25i6usQbfNxaerbKhff
tkXJeDy8yNnEH/LUcnT68htrWK0E88Z9vbPzPQ41UlzlMITyXHb95xwOR+18PgTDVLJcUiRyt2fG
sW+aD0loXALVGrwDdu1pu8jgH9uLU8TTnQc+6hcQY4zuW6A62UbY2+2qY3bkqkzhC3h+FLD/Rgwz
f1O/+Q/6QZMg9G3H6KI1UGp7LeIApy0j45Oj7x/xQRAuPzodIv1MmgyoMNblyU0fCyCI2I1+Q2w5
joOa459vyXhkdLzaF+/18tI71bYN9SZDCftCWwROCtIFmuI156ndQ2IdaswBrgdxYcYbYZOjBarP
uk8wX5tDYGTrtdVsf2042xxozky5RtKRjYD7E3WLCqdUgGJt6TgkYRq+RLeRNE+fWg/CgljDfBk4
o6r+o7fmS8GORMhzBGUqXTE8YqdB1hv1ZFiIRkPeo8+m3S8TWFuIwuhv/Zko/Soh33xacnmDwNwB
furT9tmM4lxJ1yDW4x3fDcH0gRLs/0lHL0D08s5hYZzBzcwVhcm+Htv88pI4Kh+A3mxFji/1ONLj
OaewvDGhughF0l1d305tj9CBOOtejgDC4LbIHtWSOgFLFvLoH6TDrkSGGgNcD79NSaV6rEwuy0T8
6076va+lQO8pqJD14q8OTbk7WjtUYJK3SD1w3YErI+sygSTVWoEILqBcPjOjYKdL0lTGFZ0oiudy
rKR0OrQPPN3j8/VGQtm6p2xuVDv49XHWdSVqquQ6uiMGsUl1GohMYjYmnngSi5TcEIP4jOsejlHB
XoDYgNQnXZG4LsxHrA0Ty2l62E4JXRcI7FfYOHdk5a/7YxFyquM/4HB9tIJCCTXd/R/exrLvCsWM
kBaAaYjBZ/Vrw/eBY7ghgp6/BUDc+EfEfDyo4eKDaKsNhRguyQlM+oYxQkgWr5G8Fkyh36uRFSrJ
+iSJEKJkv1tt392hYaOWsX5ShTO6cmRucfbofCe+/EkDyUMiucm8Jqtu25NgUiHLBh/bnIENENCy
WxMFA8V++fJMBkt/iEMzm8EJ8LT7aO0pS6kx6TOSfV/Ewh6NoCeQUWnkbZFdJKNz1x2/JHIfdc9q
felE3ntpjWujNe/CBBIIi0kPqThSow1pJqxrFKx6KgOSkfl+wJ65dYtu3wpygr1MUP3D3NfHZoBT
5MNo4/p0R2wRXrsvOjHZK+MrLfk/GRj3Rx8XQsw2z8wchzMOoDVps6kOyykkXv/6N6ZlcxUurrJn
cra0LjMgPTENllsk2h+QVSb0SvrAAxGEPAAhHVlK+8wZpEgjxW0qIDamwOlzZkaLMn6nxOowXZOU
622u4DjzNcF7TxYzMFMqbUxJoY9lnK6PsPTmFG4tKMjVxX9br1BNfcMRhdUvChj6N9im3UaxFoJg
o91AGKmKp/xKNszft0FQyTgJ7A5Ysc3V/UNvK+lXgJiP2XTH4wzkoQTIKoqEtMyKKwNh2NMbV8M+
FNfXbfjFcKUJut1Y0CDMFq0PSQnWi/0f6m18ycpO0tDuCFAfdup5+j4sHCFNpXWBMRPWaA8055fC
nQUKlbvfCXNf+vztnc3z0EuP5R9MeTeYLjBuq2NbHe6J26KQ5U9ckImoU1ATEd8Mb8gXBBl8J3r/
QaisL/wsHCfisxY9DK5MVTmATHwF51I9h/KbZM6Oyq3/ALj3p4tRFH3uo+KHe3TxtcDJNVl5PmyF
F6fA0/G27ZUQk/w/BARi1q9mGC1O3+g9T7RRHZ4Nh5zJBzKW/Ipq3MXe9DgohDXWuI7urPxoplNe
NMVe8vEILBBEQaBbT2dXTZ6BA4e9XIw3blvliZ1unQAktlspGatUTiuqeMMT6XQB+XoSmYGo7o4k
Q3wTRqORl7J4+5xJ8pRR8nTZ6GCCHo0NYuy4jXtVlFvKls10ItIUOQY2KRH28bjYVCg69LZxe/HI
xii3ZvmSMbH7pP8yr6T0UkB57eakpA9BafuT8ArBedeiBYAy+wMSda/k+g1gI7Y9Wmh88ZrKyi0X
m4xu3PK6RY2kN+nmGohw8Ed74aX3XiAtrgtmqUjkollneM9D/741VlW/D3JTqQ5J1p2r2ln0PQ1B
tq0CZ/3mVWCXkd/kr+Pv5ad43luJugSL4AWgNQLw0BAWCtL2bAEeCvUhzz5FYtPvFcYgwXxWMMR7
aUZm/07dU8VFqTsPOJ7SuYA/msBhzJtTuMLlVXWycH4ThMijM4y/C+RBjiG391JSEJPSvYkVFNTN
PecwdPt3cBVuL2K3n++jxSkqNODlgaiKpR5iJYXQ08SgKsYZfPxc7oIZkpzFA/kxjSys7m02yxVL
DC39nboy4GLOSh7+YeIwY6avA6DD2BXmm4UvLU3LIMs+3OtqomeJWmGZLhqh+RCKOgGkY6JXjvxj
wS7v+8vpFFnybvj9anDrBJNKHsLCXfNt6+6ZAEAumiN/3sitqd3z+I8qM1DS9v86jL3aj+APR+3l
rsMGHwZQ5KZiWd+mv5AOASnVn5kPozbz9mSnxKdw8nt3tuUoGKK4DAdOX2V9yvt/VfZBUtSoZDrz
n3u3UqQvjNmCUpkPOj5iuorPWHIUhlrJOFYUa+W9AKOZ2FCiIV6Pj3XWsmTy4VllLv9vUxNEQ5o2
Z4mELilrau8DcrpnDzqOIM1MdzNRdIa4AH3qCk0Hqv6ZCKtv0oaY7OyI/mv7BBJ1eOS7U1RP6zpb
9pczj3mrAWzx5Mn5aVjk59bFbf0wAtKgjz0E3ixqYziv5eecrMCSwV8gtqXhYTm5K0HNIvDURXE+
sG5ujGzsgdxsfBsYPHKCfmFMA7dvGIcUbeuIOGyOgl2wannG5ifsOUuJ7rUSJHoKdPv9k7t9qWTM
O+InM8XrmKFDcY1fpNUeKO6EVtBXm1kRdvikog8W782t3vV0hdOYQ/lpOs7VfvBkk5HjqBpmD1+x
WjsDDb+mNnWhUupVbyf3BoY5fbyCdJtOGpV0jENuoyrUv4ql1Qy52I4jJg7E+EDIU+cI00wfw0Wq
fTUsXmQeJTdA8OIVdfS/Ak24QfsOMPZ1vTLbQJyGzVQeiDD4h4ndBrWWGBooErztuQ0Zf9sPMrjK
PsoQWLuzKkaawE8ikUi859pBWINvwmnN74zi9JnhlU19OPI+slBb/vtkEekd/d2fy8tY+6VJEd9L
y3rJHfXP/0UKXr6Lh4Wr/I0UfjyULY50nUp4WsKOaIJDTlZcu5ly4WkWM7ky26GaLJfKxYapOkzG
Xi95pW6AXQ64zpfYV40r8BhAGn7SAH5mMaOEw8SUU6B143rdEJsq9ddu2+zFd6TwbwBargyWg8BN
m2FRGz5qzJpPHX6P2bytNWMihsl2pYGu6kT3UN2w5fjfvXuX000bfup72c5GDca+eNm2H/xaozFN
LvZPtt+wipam/MTSw0EGCOCTeJc1AMjTl27b6bHKi1MKMT6xd7wBPrTlDnnYtKXE15AaPeIdP0JV
b1bB2uonQVBThqJxB2EWnXDiA2FpQAN/sj+M1yTtElZM0dlcxCUeGeEHWeAalnntEnrZRJdyC28e
s2vXXjn8niRIhqiWmHZXBszXFgIGE0ufB1mlyrqhglIx8g5ffWw5lAAzOlOljW1WwLK5/nrEgSe8
JvlH2yzCUG9FDqLDWE1V3HP60SFo/Cp2cLCnmFu8o/DbtOcp+WPvsLROO1tTpa1vW52b5gAIRrz8
Ejm4TF+aDMLTUF94kZElGzusfcIMgSs7YArdKH/5ENywHD4amvGM4x74fvoRCDzUMKiotC1ZlsXa
lImn1x9bqOlmWps0uzJOYAHW5n9if3Fial24pCmlq4GvnSwXH+CmYYJbyVA5HrFw7Q+v1BlbimFv
z2nM4PV9j99rbXEthtk8gABXQE/Y7AS3TRN5LWQ6/1dblDohBC79PW/jGuc7d34T4B6jeFVEzxu3
1uzHnmjejtcqHaDxOHJ5295FMv4Xqi0/xlvJ92YbQS56h/4uoDTEC0wC9IytZeyS+Sl3ONR+rxCa
QxrKpl7xcQO6lywDuVI9hlazkx3gD23hxvKJBe9U2xJOPFtzTT678Onp+7fAR3Y7km1r8h+bvQAC
N6pzXToif/eVAyzde60Hq/eyhQ5r4J/c0exUCV2gKgi8fvbpPn4Ej7WdWgN9w3NkemU947ZcnmIe
eJn6DnMO+TEeNwSpxL8T63qW4cvhJ6JU5PkGEPeX64olkkvKdUgeq1Il/dWI3FIKzqKIrpEFIQAc
JQXDsCx50znw7sIxddMabfrJBs6Ym2ZVO8m+qVhS/otBW80wblpY9QnHXXP56K3ao4D6ucMnGTd7
iGzjYdLD+3QkcZeCOcBEodbgRAq+ebim9EahCdl2vUJhNJ/5L+DToPMSBeevWg7s7Oi/spceHwFa
MVGfLPaHUQfCiupKEFa/ECwu2pZJmZBj+Zot99YQ8wDId5W3MaL7+JWG5rbE3FtBp6rzW08g5CEZ
fgkuSRbP+cPA+KfFxxIab6YKGGFomSnPDg/n+tlIU5JC9vVNw7BL50YtWiXv7mGlxwbFL2tq8zJx
McStFVqwXwIplqH4xHuFnJwY4724KZzMEpnfhnII8d2K2RuFOtbGxaxGaSlLMgPJpMaJoGtwMblf
srLN+ujWjn4lJKYunrxLkGCIKgDAJrjj8TfQU2LXkuj4GJ2A5yI6Xr30I4KV9RTqHudD0S9Z0z8C
hQv24mxVc9aFyIqUxjdyVJisNxLQEI/4+o7TZdZ/AT7XW3Nv93h+KjC3nbg47woXXViDHzrtxqgN
eLJx7pY0bIaQh5zQ2guV/X5NiQNrqbXF5Dm7yqwCaC2LqCNhrGgr4bp5aO8gOZCyZe4qUf0lwUHW
X5gOpxetOybXZSZBPBJqf3FM5p4sxeK/OrVrKZWYV9gppo3RmQMEkCZoZiqFiQ6FKTqmZGP3kj5M
L5Q/IpIl2PJ/miCIZPZtxCKQ8fUE4Q3b5b4UJRi69ZhXfe1pRWcHy8mARIzrmR5J5RDwoC+iRKZt
7TainxDr6ZRv6w/tBCO3w29KP7iWz6rcHAueZMX9g/3bddnZRYfFF5Gjv7knhMK12g9dz5jROrxE
AsEOkoQjDflX
`protect end_protected

