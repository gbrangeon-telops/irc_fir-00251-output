

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bvOwtDo+u1XQuHmmirIW0G1Eep8h4q1lu6sagQVNOpqoo1dUL25zlZCKWpryXBrbavlsSVZj+/Kj
u5U6Rqq3pA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R8VeuF45EN20zhkGmJksRGl35KTSV0YbXBmOJfN53AFOKNxf64co0R3kMl1KH48vuem/BXWPzNwW
17k9On+EP4ryAUZ6V1YvtlO9Er2xv4nZefuEO+pELxS67R6s3b0HhdPIKa2fxDF3e7AwjfjDxMiG
HOQbqK01rVOmqe+2yps=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qqYTedtVydnDu0uy4wgVS9xnI5W4e3CBu2tom9I4ji9x6Du0u8YzLw4sHBXlBjTr0CIBWi+453uv
6i+HBaHUw6WLmgP+uD0PvRoMp9iMm4rcTjCZCtUo+5bxaKDQQyKy3VozWJN9cYsOEXUyn41sbHk0
MfnFQ231FTzHKrD8+sW8iXzJhrvAxVZSOCQNc8FKSuvFHDKgrQOZi/Dde7fskgmy7Y+pQzZQUv6h
7xsxzMyVpdCwJjhjdow/xj17Fc+yTtNKSxkHMIxVK6RXkbOidb7jBkIw+8aEzlqsG5f5vpboGqLH
6uQ8IqqBeKv3BDowwIwUDotWgCgTdyFmv35LwA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xgoCG0tChkhv+ljdCxpV0I73D5nOgliZqF/G39R6pkQNEQixpt7jSEz4sP4s78dR6d8BiB9A3KNg
s8gNghB9SqKmhRG0Jvm/hSIBQCWAqWOwg26IvTnT3j3MalMVsj1r5WE9uyiqdJ+QCTo/Y58NBx8l
pM5ABblrTJM59LnIcqI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VTcA7V7opij8+vJ+tjjgJGiOJ+o6V1u444VHa/k01STvZB7T6/Ztq4KXHSVmD+driESiC+2EQRes
dfVcUifCMaPU4kNZrlpS+Cz6GGzKHuujVBDhNOZum+ncGM2VGmayYd6F9EbhwKFTOVOkQmEz/eFL
4IAryyIE59LghhLnEgKJ/yOFNS6XwipLZ1ztAAj7QDruS/h8wJcmBcjwC4vXftAO79YXKmVgRKly
SlrrXAPgfawAm5V0hj7SI23oHUFrT671NQiN+jfhZylivDC/aANQXHsoSuY7NkiKvHESuXKmJ3iX
cfk8aGjoqSspgWZUBuwV9vfaTHDt+AtBbt97TQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 174368)
`protect data_block
y9m5qsCNo6RjwGRgSSJoOLC6LYLBkTGvt1DQXQE71KvhRgX0cXzZ4ZnknJ2f/HQG6IAmRJjFPIOd
3kiBoeecyxkTfH2c8LN/7pAWC9nUPPfNCXLL02yc/GIbxkLE1+UfsqOeAFSYWNcbq3cAeJIgzPPC
w6nF1685sO0erRGp3NLHkuU1hn0swZvtSggHI84tcQFBB1yQgZwMW3CoMpVRmlk1NLHZVrbYp2Rq
cxZbxO/T8G1KV2dHo8zgSKlQ/Qk1MI6YnE73xuceuqGJ4rUzo6ITY7Ncm0fop1RrOEDvN9Vcxns+
W9tSUXEgywR2M+1QkpeOVTsvXEREmcA0s9sB45IA0xUGr38TNZoDKUTOGLh/8JCnmTDEeIWaa3Aa
t3ZH3dbkRj+9UMGtT33UrDeE+8O2QD0i54z9Xcq0JeVxLH5B2EYNgRJ0x97olE8kfvZI8Jm16UEQ
Kc9+lsbxgYb8TFl5i1W1yWhuA9De357na4MaQtb7bq13H/UOqScl2gc1h/3A3fXB15C63iyyuDm3
HNEsRbmMNkdK/2IDhFk1ctUf9PskgPpftuaIRy2QLtJ76vPxNAYO4jHLnSdS8m2pPNQYldxZ427U
8Ya2nqHfGwqJMlAALaQelYoiuhW37eiAD2RuiHopmtEpNqs4yXT+s2CEf//YjeomSrkF1B+zAjtD
C/u5qBKIc0FjO+d32HhXq0JbM8VOXFnETb0750qH8otB3ENaPWOjw8ijmk2jXPN6FYIWwR6zyWrt
yVnQ3CRlr2wihttegCe9WCUi1Fr+HEGz79S//A5j1UMrT5xfce9cdRUnlZBPL/WC1b0g2Sk7Y3JL
ol2Ux0NhofmRIuL1eV5o6i/+KrwZxdRkJHL/cil55DlCfN99rS0P+2ijitC4LpvPrYLBQ4Sv8y2P
aBWXxaQxAXmY31CqPsm/E4jH8AXJgwX4fclSd+qqCnycByQ3tuoONMmeShv/6eNPVcYZ2ckX7Vcx
CrG4EtofcVbyfhm19r9HpfQIeRu/48/Lal95CXdQXOPmHR1JxPLFOssn3QgtnY+PchOSIXX+Vsoj
MR352pioiMbG8r1S5KZYfmZPKwjtUBUNF9HfN11aBGoDEnYN0sZn55lIdyjeF9KdONQKe9gACJTm
aaBUf4jRez5U6hGQXL6qnKVNkcl84mD+lLoQw1lEJJjZG+2ieaimlwQPyNAPHoZsSmq5JglRVyZY
tFKsO98cD780Xaw1dd967QeaRRp56ACPxeVrTM3YCkx9Wc5VBF1w1Mm1wpyNrEOeDIc5LbFu08yv
/sAWqNsHmZu7UzfzSmKMnvDaiQVYcuwDX25F09AcL6S+/16cdBSRqVbOcpZ8EJm87BElSwPS/zBv
WfNK0oziiC60UN+4rkHw+1yIOx7qJclmvzmWIrjetGXUYqkxiY9TrJfHPdrQ9WUakmC/IZPEyy6W
z5srHNc8a91zQaZmXKflowiNIoZeS62AACmqAlMmPY9m+ZNRXHqU0VBvLwB6qIGl8xAH7PahXjgQ
CVQkWlGF/rp+TCUiVL+fduspk6eP/Jb3p6VMRL7KX6fca7jt0+Dle1nJ4JL/9FwRyPsqjh7/+9OY
d4ByKrGjqBixQjDmkNhGf56Bu4WEm2+3RjXwXsR1ANDdl5El1Awh/sOP2umGmxiS9FinkUIK/AS7
7R5P5MPfc/UNp+/1OJzyHN8mPf8Fjq4BVTbDbxa/646C86Br4ZI40C53tXUVNHmVmkJpvIiTQKOU
focNevm5uOAfP6EE3YfMRfeSobX2JT0FtN2DaLLryV94jKatLwXx8wMMH+wHD9zBRfN/oQ7zCyXU
pKRrcx7o0YoD7+KhTyI8sq/eEk2U9XJejf1SG2Ggh34g9V889ARdhSbZ7AL+H87zwMbdTYYOpRDj
Bd2f1caFQY9GWpFTXljt9AY1pVyCi6zannu/cwysmTjxhte1c0GBxcQuwSISFWiHn7DV+Q6i/WId
SA6yHhHpFwxU7MAcWeepGFPFGJgCeNMKDsXpfv3jfprtRuK30vdBVrdzCVInK+XyoBB7gAhrMSQb
+cEl9GumXqJ8MqYj8z+vPnDwxGn0PTT2oBjcvI1bREDCqf6hOS2iqgD+W5QMq1DO/bvNyLl7sXSX
4bUhGdeLelPWwuJVXYc9WySYUV941hwI0OYPltBFmN1KotaqTtmvV/hXufwcVEo9b3WsXU6W3C1e
a9bpPqnSbmycntaemCVE1yijGbKq08pmYRvPBR6f/nGEaX6qu1CrsV7+iByVvCxXkO8qoOV2GER7
yhqJiFGGjFZQ0AhGcelJL3lf3tUkmwf2FOldnH+GBpuCAblnxo4ueMXWnmXrd9GhzfA/xNgNBsUH
+8aY0Arh4DfuqSW5M100rzE0hW8DpvXkjIEYbX+zbTZ1fuwUyvifC/nWMU1pzRiypwtDpzPNRLg9
7ZN6eg54Dax5jxk5+wUc8dVr7N0sc9g5wGKFYTYF787a0dH6wFStz+h+O0Vj30hdtbh3jk3GOgPC
G42yRW0fjJ11fL4t8gWGELUCvxg8vOO+WHmce+8TbdJhnIHJoiZOhaS4R3iX+wMQvz1EYOti/mKi
rwV361C6Tgxsq1UEKVcUAugBLSHjQbxKmACaBa8HMMYfYPJTas8rZuvRdRLVF0M8loGSaimHmcI+
dbkC5L462KuD0DMN7QZLeXv5YM+agdYXSxotKx1icMx4XLdZ4C4RkIrRSw3rcJl3mdIkEajeGkLK
29/L6LHG5BLWMY2eMOVb+Qf99yIjt1srPhB15Ldyig21l2bIuUTxcvFEKS4RQkG8xsh2E2Gc/pbl
C79f/ovqfVKzj9aGwDhLC2mnSzkJ+Bbd25NEQReWdcyylS3COps5FI0ToVGGac7v5K6mieLSg8ss
7oEocI43gcFqnLuamZGf0JOxfxWWovtifeEI9gV/3kKqJywPbN7bfA+/lGtmp4w9loVVZSobjp/H
pYh2THFftkP+Sw5eTDOHR7RdFBC7poYyyNjEAdJY3CLf17rVqd3UtUaPJ+bZQ3E/XRywVhjxm+Vn
zlEC1vAOcZSqeIbSRdlKp6X9mqa92KJwx3yHAMZ6+eGSPD+M2oEkcLZIQfI6hFToZcRJa2r9cUuA
bzOVBvIHkP2i3Juro6tTVXlaz64/bAvOeIcrp5EOCpU/cSfVDbOGaownM6X5iJ1tU17VMZ17e7ov
dkb5HxwtwUCoT1Pe00rrbz6z+D6MF5VceqSLcJl2sMp8wzhYgzW5hl/rc3yfJEzxHwdQRUiiYQfO
R0gHrfx+cr5TUfR219PV/N4bXqAjMX8cpVpEFGkADACG0s2w0O1OQiJzAIbrw+OAi0isA3yYVRdv
Mv4Cj3hmE08SK1WaNfNKZ/pTwOWoxmF3L1juRo9UufG+jfGeRGqIqItgeQZePDPh3Ct+L705oBG4
TW80wAthwbw+OOWEj1s8/qQcw98QXmeqOGpWEHWoKAQ3oIjKeORNH4KjYXZLlVZFhTTZMVNlPhOB
JKuuYrvnhGM7u1zJf7Lq6GuypstIpyik/nu0iArTybamQhQgF+ELhz4pmwFizfOYpIWI/uSzq74y
CnYMfW/wtwid8StById0gWX+OToAe8ZKk5we0QldYzF3V8Rbu8Pok/zuV73gSz/ZsV49LvyN3DAX
P8OCaIMKTT6IE65YZXHqdV04ibNf4CI6UowK4xIVqVuseu3dPDVr71LEegZXR7PLm+Q953s82W3d
unKBOmAJBuT+0R4GJG5B4yw2otTTVZb7yQu4w22dNkt0BqiKkyC54gtCSoAMe35zCYEcLeRy3++6
7KLlCZ9WVDSNy5l+0fQlS7sTx0oPdE3vS8b1nkjP/lY6Yv8z89yq276ES6ZdceQDduaXJVre980b
IJS1/RE4l+/CqF/8oEg3zXsRDXjwg/LXIq2UOFZiYZ/FPL9V3+vcbnVnhLoKsNem2YQS2hNs+1h/
tcWHx1y5xkKTpPOf4dHAM2/aalgzT7mF/aOkkYzo44qOm2cwvIKXLuN5XcFatqM/ETEOjv5nczuO
bVHbHKuET86C14KhJEqqt4452BLfobRd5mfiP/2SZecgyEIkLvdUNVxphyws08QZgJwa+E1an0k+
bHn7hdlBN7LnEB/kgmoMBWEPK80eSz/DNoC0HLjCzcWTQIvEImStviJzCuB354tF2qrvao4ZOQXs
ZZ1cBljw+6QwfVdcW2h6tiai7p/A/Jbwp4cfsYtv2A7JBtesRrMXckwG2rmJOEpDlR2t50jqVUD1
MljM9S2XF7bgx9F3WTcey8eOS8Usow7OmOPtiIMH08Q4RHLO1VCzUR+OV8i4+U5P2xeWYsaUMYTJ
7nhPvY5V54yx8A28lSgBwJFe0vQG69JMDzqOy7PElNVhMbXpRCwwHgNv4PSPsWLxv0/irfz5hLNj
LWKzIQ+e3yudamS40RSnO4i/KF66pPi4SqXxLfyXplToaOV9Nb1MQ3BqI3zCanMzM4rlhegAePSV
w7uWgCgAOpLziD9oaulPxf3dkhWni8OW0BXRkLamPmyXLXSbUoW2ihNI0utgQzEZpiKN9WXqlDTK
Sai3L6l+1pvQQa5s1sC8LJR3WOsvCpPRrhPygJ9E6P+sU5zU009zeTQr0ZmaPxflmzISHRyW2+7e
aF+pmDe5jtpcL+5VHNEv5LWdqxVUBxLrIViZz0gTnBO/o+haE9OdHQ1ug+k+hPICxsXrdaB3EdGa
kTGNV6ns6SR9DtoTEBQwRfeu2Hp4YB5D5nQRSDdFwnLlWTtfwBo4zlFWKwQtZhw1ih4tZLD05Q4q
Jf8fesdYVX8HiGC3AhiKou9cQgtOV72nE0JZ00UnHJdRVX6WmfEhErCD8ZAu5jqzdsNNZECFIQbp
niTu20EBSBkoCJ0gK1qyu6MtEkSOQgvXhH+2RvAiewq3EcEmzkdMFTwxiEtBsWA4BBv5ohIR1NvI
QQ5KCVRMWSxPZmUkEuuvFwNNreoMBuX4F0WF5rrzLQCdB41ol/r4tpu4HHgtfX2dxKXMv1e7XPFF
KtCX8Gy8/2DpbU1pRsQPvhaJAniCJXMqKIrJRY267MOLRPKZVp0TjauHDt0ItOWXjMgQo6QFTPu4
vJ1+5EL47zndut+s8w8gr/3Y3peJxU/svPpxCbUvyi9cwZPRZlZbUa1KbyG0xb+ugf2n7Hud7ErL
tHDvpV6CdupZsLW0tolMogh60U3xUupj4h828GHu3XR+h6hTBVoOG5ZiEMNctMT/O0wcpbWvRkWW
IAbfV339teOifzTDDlcQJtceZ4wGTkZE+S0h3z4elSa0ishCaj5cL3XLM5jYZ7FyYxD7fEFmCDTj
3hGJ5ihl0/IkyvDZkvGpysw1H+8m50k5ZWj242f7WdrBjbA/MEPev8oGob91MVJ8eB5smubWhGjN
PlCPBLwMta4wnPia+WIlRRMujk/yVQgNBEJzcwpeUU0+AZzr56jPAvCTJa1QWQEsX3ehPCaSHRDB
bq5K73oQITnS6EmkwAQ1jFwTayADwXtZoBZK7TmaeFIcPPOZ6sL1klcAdH3ih33cxetuesJLLEgY
0wNUUcVPfc/OyvHQ9jTE+S7UVYMdeadcpZuugubZCy39eomiGq1S/zstpGf2MBGQ4AXSGoe4AE1X
LNNc2BhUib/UNty2XwNikyCd6EjEGquzWHXE3dF3NfmLFqusBleUvVWXQXWwVDBRISQqdC9chDKy
CkyT6cJzoWahNdHdZLuxAjdfvvD3xp3P5esq9dU8WZv2iF2160x5Zulz1ETC12Kjlmq6ZU4SIHUq
Jf54tv/ZDu91bUEvsHHlyT6Sx0Mvbej8WGrAE1Z6gndxeGTGoXOiDCqZMEGXTu5ysNF0ZbcRaLCy
lWRbx7R3TeVq7xvmLR8RRMJdYtzwu5LqyYmDL61yQwxdu0sC3ovI/qfmQSLj+rKqeku1mQ5PmQv9
3RyIDQF2MwoghQVBcn+7cDs7c11qODTG3L3dj9sqLZmcg52C9uxSCSAtDT2/75jzOqcM2ro5n53l
dFOaU+t75woqMlawCWvpv6bEY9XWy/yTlN//gT1jiAO8qL2ll/6rAiN3pcZMMCMfKUAQ5muPwtPi
AWBgXH3e3ZjIVRd/5MU+I9keHheNaSB+SckuefJh/4MADY70NlEkj6P1ZQUabRTJdWbdQwJ/koHa
GvXakFqJkHq4x81ABAOe2o7m6oyoIkeG2VpfFgsfBnOn1PNM+7bV/1/8pIaxWJ6f+iGTCZoLxxf0
PgLZMGs5PcX3A8Lu8BtPpo6tJUq3K+yNYvEuAJtXvojD5avf6vP9E8Nc3rhQVGYWIaosmf11s7Hf
NzcXKREuvxtHHMoGZke5DGGma/AbfOT+RZlsuAMFjV+depa6yf9qC0/sVDno9rIJTZ5k9XBnAbpv
BeFiLFDV+NCklCGQ/ot3nl35T5fLOezCPceu1Hv72+EyeJD6CEfyaTJKreljJVpkP/UQw6BtrRkd
Yhr5V1KKzQW17yhBuXheUYzrwBkUvKJfgoCyXqz2Wyfms/0Pld3MBL6HKTWbMpQEJBbgIA4zuFSi
xVswgxO79bsX4st74lITTj8cmHSk7elUKNzYsigERbyqL3rs2tPtuErM/9Dme+T6IJX66Nj28xG2
+gqyZdzR3r1EJJ1KApgncN0yrkvwEawwuQThZQVSf4nfS8JH9Abjw0Q78G+mP6vAh1CARPSNPp1O
t+qUcdrX5Hq2ud2oMhf+OH+UB9nWPm9a1+KEZbUdnLCDAve5Xz9qN8pqnflq2o5FVoMeQbjk5zEA
K9BcZcUq76MXr++oCzZZCIjJKJPJ9kv5yMUDEbW30qjnWysp+ctHzkYHsI46VrIGEaZHepMlA9iZ
Y0+81zA6JBJ/IZ4hHPwp6s/uxkWoEk7/wzRkU0lWlca554XvY8oM1A6nwXZcokc/VCp5Wo3W5bDV
hG7zicWw6TPp7mz44q6KFN00qZL1fXjItT5MqqyQMw/kQDfneVtvbyZ24qyi6w9Nknaq8QW3vclp
9gGj0PVZxMIX67x+kfhNwNMvPnz2GRYdPwniYO5PMRX3eXNxxiTjSl5Rl8+IFVkKJqoQQ/eSxnz7
BzDiaPUg2IZQ/OJXkTHIgjM6GgYTmOQEEplOucHxNjtMcG+6Bk9boyB4mgnqnOdGx4hXwCJqgcyt
4AZ4V6ccXqQpIi2QHmycReKmrNRPGSz+9DYYvROJ9Os17ejov0oCORgzNb5qQvH5ruMF3ALtKr3f
Ey/y9ZD1EdY1/mlH9I51byzdBICGuPqMOk4r4FyLGDYTprXi6HUcGrQT1sdEFS7gXW24F27LXkIZ
IQIM6+QBSxa8SmPcWPxk2Sp0HnX36NKnEgc1SOUm2iv7UxKiK6zNEPcdOmvH0JVUxmVnPuJ9lE3n
+OJGh3c3g+HXGM2j/5VlIbCJZYXT+bqxae6JIklrA4xM4yp3NeyGY8l39i2S0uPY78u5LMP8N594
w/FAD6g7JIfxdDBeZc5er4UhqZ+zxe7YC+eaLQmPBZLgp353ZRAgmqFdrcW1aVRvcyi6yp24wkfI
g1maVJdLaVxlyBi6/r0+iCrj+rFd5kKEKTHfGEsq4MDdD5x/pdJVrElksyvvj4h9LLhJy/cnF94F
7c/Y9bX8sFCy6v85f//kQMBYuDXCmVnPM29IMESJbofU0ULoH44d179KETT2qB3Mto/6b/zB8CVA
NyobN9HK6n44EKJ4THLmlR44nnVtz2BTqWQmtg4k8npEoQ9x+SKs1O9MS4bFkhi+25eW7Di0l9Y9
2KHvfxxY93x8XDj5pieL83CPatOrJC5OBdRn3ksdv9QqM3rIkc/gCq76MxxHkV+1zKc8T6Z2HIur
+c4pgfZpfeNUYE/JrqY7zPLUlulY5o6KO5s2bBhTFIIvpcNu1i8wTIuiFCAHfzuIvwE0CfLkTp35
GD5x5neLx5pVlfK+Vo5djybvlM+GUkzYYNAdqYEIWUar8Ga94a9Eh5/7xHLbMDx9YRC3qH8UC6aI
2SAZw1RdsBOb6IILQfhTtdr+cYLIu1tH32KnixgFPxeWlfFOFQdzdpXKIGduut7vkGi7Xmbm5ko8
zrrAzm+7HrTSUXDTDQhCYyA5dtW0Xfvj/wOAhgCtDqgIfdUbt2arj2TkOwbaq+isTkwmFNjRRW4t
/yJ1npQRD+jilRE8eo4QHtgvIaYF9scj//lT8IpfwI3x+/Xc1q2YS8p1kbc7KLzb0VBlyLHQL7Ur
7xoM1hTRtVXi8ukHeEhjKUonj2k4bdhVzox7yQCXwAlnB/9YNT79oFT4nEwdr3bqVEdIZGpt9CJ6
QQRpRQWPr6t8NffOz2CkXk5fi0pK0Oc1UfoOkrgl7EQkbojWum9CzB41u8OPDuziMK1XWr23XBzn
fpkfFf88Gn/Awesa6ASaFL/lUx8fktJ2+fo/rtax/j65B93136nq2lwzsTuHDRERoiFhIloIUOiK
9Qyeqekvi2R1pImulyzuxa9qqvLo8gRYrn46IjrwtIpMze+iTW329o9KnKaukE84vUXptxigv6gU
h584V45weDjkn5PdMxPlWjiQQNJZ3h1KkkQnREHFC+mZKMrrlsNRCCHC0Fslv2TuR+iKHQPettJk
D9UgdN37tFCgB68MK+4C1na5MYfYqUKKEQea/PY2SS6hvsIppDwK+u4eFoa3Irxttv09wh7iwJbT
tTZT+YT6RKSeB/Ki4R/tDwsqTt4+zetUd+Sf8rGZKS5VW2MaCuhiO6q+n/Ra5zLG2bUeFUbnL+D9
Mjj9MK63b+hKA7JS1QSUcsMb32NM6K9dlLeTxxvLkAafrw6C+/NtLagFcvjYO0X3NpFNJazZonVL
naYuF8+DZmk+cq2KEM6p9VsrAqyYnpb0qDBj75dGAXLbLSZfAqBwW6rTz6LDSUBFnsysdgvcyXcE
sjLhehBhDTCkG4lvXQ7wX0YxTKlK/5Mmsna5ErrYNSZZCaQACL/GjxZzbwHgpjFB11SxlG19JnNL
vNEXbxNvoO8g8mDajVpas2NXI38wI7ZERFrXPO4Xi4NIrgtzaUIP7VOYw/plfcOktK8smW1bQssP
M3Pv5fYcZKvJu5ymTalWdKHhmw5Y7T+HEbnxNc8ew/H7HcTfgr7xKBMBKYVYK8v5my6FiNRLu/YS
nkj562JaCyxsK5wHKQAdN0WUYH5X+IGG16qJzH201D+JeShuoJElMHQjQVUWUS0l6Kv/PskL2o7O
9+gkChUbGcXkE11kH+ZTNyvGVG4mTVChPd90ycRjn+R06vzDWNBlD8ADsod5AFaWCrHpeNw/ecFV
X7qAGcAyNYUqNjRUVIzC8CS6sXj/dJrbL6+kBn6g2Sys0E4CiY5+5/iBN1XcReh9WaYQkSQMiqLx
cj8EN7pVjyrKy80yNDmWeKRIC70DAeWSI1pQLIgoj5GnQNOFpgJDGrJzRLvmnoGSVLUu/3sJxgi5
WsLyvx1HJBgVwStDIaG1WR0s3GkdfIX42+qR2JWWlsiIbyRb3VzkcFW2KRR2njmsNBPgtD9VoqIA
w518hxfWF7irUvN5j0fVpCcvf8m4lg4clxeCbwD7aC0fVjKSpvuLU26MSXHGoZrycMtATfVea+/i
cnmsn0UHZHzk+CURp5v/0V9eLd+wHGRPT/nEXNSfeFHkTvVFFqAcu0pOm+aPmq01KrLQHUmSv8LQ
CHk9TsYsaGQffWNZi2IcwhJvl8+zF/dsFw/ODCvv5rLeePSSRh6OrdapfEsJhRFMWXAXfqjvrGBa
1DgAFgp1nAOS/60q5TbS6DESX3mgavWLgWu0mwWvPBwkpZHpDIwpJPY8MddUwoyTGlDQSJH+4GoQ
bczcjTZMzwYZNyqhi80KkbpgOX7Vy01mS59R/5JVIPeVAEHVBNM0Gdu0cj333sy+a5p0tmTOUCET
8bPGSj/AfuLKB2D/RWIv96oq0OGzk4f9s+NaocV+mvx1eSSL8OU8aU+h+47gT3MfFzVGsEBdXWo3
QgQCb+fkT7Oz4ab/i0A2MrmfOEBP40Xqn1oApen2ZsSeSOFFuWqKCJ5ZhCGMlwgYwAj7nUEA4JRL
YaSf6iAQzJcDUwvvKSh6cYINAueuROwxjODrGZp6ufW1UkMoUyb7qiBVGOaX9m0T92fyK40SVM67
xvJp0eX+dJ8L9AWNjIvopGpfwWxeG4qnnQKy52Qje+tB+1eiTpW4qnpHm1fYBshb8MoP0no4fH7G
bHfGMKjq7rSN1sKQ7QwaxDUdeqUOBVjgNUoFjJGQ/lgGWEGEqOePez7uYmli/W043AaVeEnlczeT
kYFmVKg2cgWNK9ag+Ti4VsaAqIQcMWPyYO6rtKNeROARJheYf9OfeCXFhgNC+HhmEeFycM2Ys3jQ
kXvj2bqRD63WIgVuXKdIwvg4ho1JD0YTuBzyrLIDTNRIfGmiAS868O5MGw8lc6Fjuthrx3KcJdTd
D0aqSVwkZKEChRoZeIorigOfC65fW780MXjiJWDHDdT24ywlxwNYDeVAEFypfTnNFzOVrJbDVS1/
H+76Rbv8rPjm7DvodVvTG88pCeKnqzWPCjBzTn/k9q+2gWjBtH0RCBblZ2PeG0v0LvJp62aZhG3F
ZUwP0B+L1KllzGunv629WR/KyeqZV58tladmuMbPcy0BvH9ro1Z7fT0cDCYpLdx9wMuKsaAUbQLt
NgTnCkQA8hp9m05nNYGASbgif58ylUEe6ud4ya1+6qcN1mS/QTsptZqwN6Ge5YSJ+N8QCHYoOdRm
G0XH7X1JiI8mdnWdF/1dluuzylUca4y2m3pEz+H5xXDYLoreHVOwb6Wd1gpQ70AiLNuz5+O9s8ui
vWbKOGHN99f8bWBAvB8i3tzDPavjiLy1FIEBOPYfnW9PdxhAUt3Uh4MCvCbDWLNVHftjEb/5572E
iTysw2qMt3AR/tGjTMeC/X7GWWbSCevV7f9p6bpreCSOegUjWFPBdXL3R9MmiwQQaByQfXPeoLOt
hhnpnOx8pmVpiz+J6wleNAEyvR13M4IVFUAxGw+4GFJKtDXDP8kPU+DSAG1yvBAE8SaiFzY7msDB
cUD/ftZcgEZcLdZi+YKxuLuxrcDII7jFSwbsXoTTyL78k+UXhsm+HD55VhMqcXIqXheVV4nMXehK
nBE1+448WSrN665TPgxtrtAVEHiqUOnKN3kaYr/tHPtzSi7a+M/2QQXrPze6zkrcTkoojyD8Kehl
XB43i5rF2nEpooT4i9qI5LlKBwzoc+0yhMlofjJnm+Bro87Egm6j8vN1tX/+8F0e30l46wSenhC+
zd1zWRK3Ho4+a3Ou6GBNsFq+OwlsEEDk3HesAyOlEyZBbum32XEP/UUf6Jqg3BBwpvCLzKUfKx3k
bw3oXKGbezvfuUv+MiDOjph5g8+EhMIQpfcbKl47BvVzJs0PZh2BxBLXGZwg0okenlAmkfh8QDKN
+oF16VlqNyNiCDuhG3ufxtuhHB4N/02AYQ6oeGFjtBWQrRuwIY5/AlclbMAwTOXSs97NAaWu8p25
doyUGOY2lkvcY1eN3s+JeKFey5gAn5iIwqWl18XswgE9BRU+GpKHtIfZG7B/5ovs8a1OOvkGwJed
AwYYtH33L6AsNL0qJg0tizC0Tvzp6n+pQoSmVuSfIVa6j+IP0yJI0YGpsey1lXRd95cfwd3pellY
I9WTpcffhSEqC/OZ0t7+Hdq4ZGkd4vzYgbrTzElEKtxS901zn+VEici8NhxZ07uWa5WqX+zbR9ay
1QtElCRM3apMD5U6pjMuegL1Be+anuZKWZoY9+JXmZV8k4DK744jTChtoDoYACB0u2+IPsyN4RJB
iaeTTd6ABBSYjMSrZEZnjh34aIt2474ThyWEAR5qvM34K9A8yRIZYCBntt+ucv4s/EFn/ViLeHHc
j35RdpoFq66f87KBcykO7OpO9LXI/XxdBzAddqYD8NjiDdbDjnOW7Xm3l/4K9O8DXsf9Ls6IB+LU
5hEgzpBm7MLAjMOb/BcqILwSbFuEZ+Cy2xyANNbRDFXI0YE2nw8SFk82VCRDC3n/6NIiunWZ5ik6
Dm555j8RAxEPX0il9Pqd8zyU/LWvoXMhZjEpSUt2ggo4cpVOzNjDuGD+Em96MUMKzXr0IekCZr9w
MB9MAI+oVpBNn5Q0cGiyltX+SsQdlZNKMkLwUEF4kL0dm+U5Xk5zT34+TQuZjWlOqGvF9aDX2wRX
9G5/5GFEiPObqg1JzbGfJnfgnLuF0Rua6j9S4Wsu/zhWp2XBQNm/jmbqOI+kkUHlaH2lLmot0GJs
qsus48DMsi6N4cxQ/hdskX0fmmKI2RMsTa0hWjm7bUaLaHREwk/itlOGJ2rTyUc9R4FHU/ykusit
mfPqCAPclHaA9lGvHuA9GIiNhfs9c3Mr/QHFTU9enzhxYtXp/bqu6R2PuVW3UaIz4lvYONh7PWpH
zGAS/FFHLarmu3UNdiyWsv7GpYQWGm9AWL5+nOT3EtDnwE1Y4ixvHZdmf4/a+B0R6i8xMpKEk8j2
HUOJj0v2VHhjvI/gABrz1MHOKQtQG+Wkcswv6po0388jYVAE4kTvhiauEhkD8oLUf3aS8nCymukj
3/ptFDkja2M9y+jtZhYWpnidkPGlghYpJKKOH0LrZ+qQl1SXOH42i01nDCrVjJWpcC/IOskohibL
okl1LyznWYSZdeB2y2M8EzccQwtBLdCMrRaQpVO1G3uMAOwM82/TwmccZ3ZCCQBXL1DDIR9WLtZU
XIO/eW18HchzW42A9IHF/Aap6/SmJNdjxVl2F1FA+HYI+zZ3S2ExvPHu/nLV8zQeyjV1e9O1L5dc
Uix+Xu3vWQmv3ptvfUCNT8GKQz52eXQVxncYgjbMt56ihRYwrOsfQq5VsLwORs7e4Eoh9YCbuGJK
aTYUtPBZmtQu4VWlD77swr7wQtxEJEmkr+lwr+vnzJVRsoPhVhq726ACs71j1nBPBorUaUy4AFDW
6QQdcjmy27yKEfCLb1OxqDEgaSADHh3idNoe39ezgEJTEIZW/W2WjTZQ9lV7khPWker8DZf7xo5Y
YXy6v8uW7cerHi18OU34cjn5/9m3g/6uspCkP7bl7UTDYqIOy9sdNMstpNnhN2YG3rfPnKiGnAVM
5recZERc2IIL73XYPt8/DL3/w+GeHezYpkSp23M60JIjAh6TBirPEdWzkjmsJDJ4EjEs+IKQYNUA
KGd0mePMImHOvTI2EUX6zZDA1tLT2a0RDhzfQc/rztuO55excd9FKRqh4WGeBSUp0DplYHBuBDOO
pPeWHH7JseUwccH1HgA4aUOQ1eCufFuzk9hoE0/b3Ttyh1jDQNnp6LKcaj+iRyiiCpb+KxHfoe2H
Po23tmz1Rediv3Mm/GeSz8moeKD7GOkqrOkX9wgQKcSHC39IeM1o2i1vrYGtIQsve0Wx2NcDIs3h
Jhx7UXw+nGVycr27ujXmXpwFSrbdRdKLffFsiZbTXbyC/E4rd1x8hENBBfe0dqGxubCpxO8Rbfd8
UvUIRmolM6t9sk8hb3NrusykaGTsd/iJ7js5UsU/+oMLgpbtAwQnDU++1J0Tee1ByHAcpZqt6J5t
e3nIwvGu2aS9YcQ76G8La0Ft8m+6fgFMRCQpbKr4jNIPIOiN20iYN5vP1/O0qPa8sRzhbLSawE9R
nhCD2wVOLcGHH9e3F768PdYVZu6i2l5zlCLjn1gGG2qOaCz038Ch1zqvVSbmyw/MTknUgp8pMoDR
m1ZtAsHzuDFUjXU7KpNcNmMHypvAqdRKFbD8Ir1TtVYUx8uF7PbYGWqmy5zF55ttzyo2NwZKt0hC
DejnQyz6EO+h/XEDKbj//4M0e1NCzR2m6lJinFYmWl+ai/O1OcIaA974IS7wfqL0bDBxQX1WwO0f
hkwT7KWqmnFZkjO0DShJfFFzaM64XbWw3DfUgOb4BlnVWzGJZDo49pckJlK50+Fy/u6rajf4TP6W
IzeHf4YtizW80ZsBM6u/qbdMK87Ebf7vWW46ktCTuCNtZ/bHy8vFxePu14/BDa7LTXU6ioN656fV
95gV2tessVagb9wC4MicBqF/BhyuNapP8bN01QZcjwdwKfM1kUz+nGz9URPAVvm8lvVureszXMt/
KxhUgTrYcG+fgl3QHwL73qjrq/0lU2EdAOpDK8bb1DcKoOkZ5gOVDFxF1CYPwaf/kNO/0RFcUdLb
fpsJNrDpoJq4sSvKcWlI8DffoRxJ+lBIvQwa5OfaqyIqKmjDTxELkqPYE3omRbkaxtG1CB0XR22M
Zwwrm9s6JIrUQFa9Ffwt5Q0MsM7R7wtWYNUP7mbtFuI8ujq7K27UvOnojRw/ca4bQCm7ncdlnP/B
LyUSiHb5uC3/yuYHkWbNdXUqRHfHInWJmFXt1szf3WkV0NM2IGI1KKVf34uw2NNNbqawh0DXCbdQ
TnYXU8Br8TJ0KYVcmbw8uKFdpHD2z2P6uQXLGwK2e1JgPgjvAJD9lk65jELuSwi7ETxqzKwW0QRK
1mtz7zelOnAEqQE6nhxfrHYMXzkOnbMlwAKIvzbbjHKZuQUO46fhWAEZE0YkqsAYGu16C4rDNTI9
Vplat/fa91cpSnCRux6moAqyH0CaguxDqjWyxrJJWKzedMmUxRut0XOMPncL/kJfDqT6dXLg8UDG
TU2b8hNKlI8FfOlVi0f8VngUBO957lDqkJFpyNpLx6qQRxW0jxj4KpOEjUAYGTKAbmiM0hkFPhYH
YiIpUdiBRsN2g6LUWtiR/vRNqYhGE3E2Z4Gfztz2GCjJKkf8p5fTadN6KY64Eo4Q4di0jZr8du95
e1Pw4PlnvSnQG1ozzCreYkhlym5cnEK5kZllIxiUjqv7vDjxektBf4ikAIO0pABgxMa3fpQdwPJt
cw5msvypHF9EQUvdz3ptSCRrGpbdfk9fffrcFP0xipKIMaOTSVu38yQCGY2CuWExOg8JCly6cA2I
8jmkZ3CXJ4PHhKNSph3ocmpXkl2JGTFpfHqpx0Ozn+YHlI5LHUgc0VitbIzCTDAZfbd07VRDEhcu
uGjYwJTJZkAIR3zzl+EvZsKgjpeO5LsLOnve2mMB0G0KZEVMRxcOjK19+FXo3blsszu/FG7NyKZA
kYjR5X9ZZVjfVQKkdTPO5EkG9BPVV9FEaN7/myxBiVlvyQ1DPgsMrf1kyVaFyFaKEG4pj1X49uk4
DD+c4JOFOA7dfB7bgctTpWE0tCOw8AiHbkX6kRP7S1UU7lCiy0D3SA+rr67MZsvddfMFlz28V2Ji
46JANAQxpg1XVl2E4Eqj7V9xb5l7NVU+w1yPB0Qu93/PHiBHenFGLpi717f+VVsuM/7gq9lM+xxu
63bNyIWAIuNlH6nnw9308sH4Kcy74BmaEUIn3jZ2Sm2l23v4FU2JFgl0qRHep04wDBy0HD8LF/Rv
xQyNCaQAou5f8pkqLFIvT/IsyXTCp1sZOov+GKVGAVlW3hf37+TiEsMJEKjx0f3tfUMDIN2XWKpW
OZSli5Z/a03ISPpcgVBZ+wrDydyP2sF/5qG+cCoPCpCDKLSjPlrjmW2A6dqRz6U8A8xFlBG4pmlt
l3AxmdSI/RvIyWt5cCi+CqIBsXMxYkzzuDjeNHcBQO70G3v6c/F2tK8nbSvH4yu/za/YQ5Vw/mfx
qZezFVGmSAuIwSPbI8VtFdR0xwVwFR7Pn8zqfANBqPFYhgrpo2OTpQkHsOyM3cPOJ7AV1n6o355z
UYRtTdwoSNcx/98ouqu9qcUQAkggfgdm8pfK2S1/8/RDFr/z2SVwKjmJERE4eaTOK9FbiZTiz7hr
hwG97FJt8uga+B6gY87sOCLEcdzGFjrxlq2jTAckactg/P8RQ19QuWZq77wpJ+AduyHjy4jKvSEd
AN/4897xUxjfLJH0znfWDlwzpUSSy43zDiJlJvlJwubshsdADsPqWLVLX2/lV0zhQCqUMvUuxP5z
eU5HOf4CYlw2HYVj0lmPZFvp3lTbBQ1ZkDaXYhmJi7AfzJPDs32AgonQttFcJgDlBF5vMn9q0JSv
ZJO8UFvVHhmDqRwA28M7zaIgOuy+Y48qRfT1ryDNkGy0IkpPRNT6RzslRHUXP7n/IKhfwRigUL5P
Y0t8g6VELj1OcJ8A7NkrFG2/lPWbKCiALcNU5+O1L8y5/osmn0m2q3wsr9LqQyD1DOSTT0ugWltK
lULPrJu3bDErTawYdzJxK7fbuVLnBHJpyiCteeMC/HiRDe8QctXfiYLpQHZfB/KUc2xUrIdc6BOo
tNJD4VtF/SXf3swMYt/jY/he1i9JmMclZnxXUb5zKyOtAb0m0nRvIvUpH561jM7wJwThoSsPt6Wm
mLiXJOR9q9GPAuM0K7kkxqHxbRPDucBeO70qrnCkljGAgZuk9K1vW3ap6veQsLeXqJ47Zqt4s+Ue
oyMZLqY7YybtrsgPKRAontrIU9rPWAUmfVstDLp/K3VhH4/1kpmEHfVcNIfYnnuupkMCcSt8b+WU
6pxFkY4IffLmj41NpPqxyjTqP2t2LEeHYVMdzUAhr7rBjFkjfqArVQMQwxi9ZV+aL3WyuoXFvEzR
dzitVwHsrtRz7BdKRrT/zmuIvfUtiaFnhw7PAjmRc9ACY2BhvGq0T7Xx5f9nVPgZkIDHsBdS6Wl/
miFSWuD4mvya4jP4am7stH5juhfTbOvPVPBrgW8S4OEtcgYbfeDQ5DWKtxgA/V7a3nfd1osj+sgX
nFbmLT4m/4IlEleSYvZyKUfzADWB7sOhCLGi1ehRQBDv+V8JusdLsb32SxDDsLDVrlEQYUqW5+dM
2dvXpxLngfoE5gr8eCRVLb308b7+X6MUiIOHbLDlywDf5RIwp0+eWvzh6yEu9U5uzk1Gz+17SCYR
L89GHuJhn3LcbM77vg7eluU7c7stU+TFNwPX/qAx0S7y4DWqjUQSfeCQ5qSBErA9+mLpFIpOpF/L
FtCh2qgTzOwMpqOHEwkG8s9gavg3OSKif3kAWhmpK2h0N+hjy48V+yK5GtZ9A1IuWYjdT1V6shl7
yIJNXzSLgehtdRdzDO9hL/rnSrPMtthKFwn0YWeauSH7HOR/4vPdalamBgdSJ9zhj63gvaseZHBM
fqVsprBGGP4GzmWOhivLvOoaoijhWk7u9TiMTIxQs78aX62mfMbagAN5MihjzSHIubPmZtcp6K4H
UiyVWMlnXmjzwEUqDG98N8gvo46lbmRvxmy3HMcyj7XqlF8+PfCzJtJaV/7C7hruKfGqF6zM72cn
nJo7TH56IwQOiYCOImHjPZB1Tuqz7BGA/unJE+fVj6a+8xvuYHwvgmo0ne/EtbcdGumYEWffYEWF
1/uPAO1J5MGKLBr/mdSIA9Ts5nV63AATfpTij4VExqkayRRFZAgVOhqWTbn3wc7aPSzM4EYfpRMZ
N9AxGN8vPZ3q1x7pYxtFjzDmG8HznYxxtTsceMco0tVsrecz51hocIQ27zofhlRsuW1PWleLsd1I
MMTM9T0Df8Eq34APC4qms2bJIkvpBIh97ABw3aN4ElX1q9rkwUCFkPA8XqUGIX+3VIMdZQv0KBjE
TCh0nzGQ/LRMXVbvSUWlZPHJFXa96vr+2MFGchhry3NaED3sFScYOjPyHoFmx3gfoVw9QRXOD9Cj
+BUQtfEbPEH62YF5a/uROLCCN3lHMYlyBRWRDgBMHK9b7j8wGJ8fC4DCGd4eqBPp8VI4muxpIWvO
8KUG9r2gk1l2vLIml8FHJ7f58C0HocZ0Jw7uCweAcLWhNkelyLZUn1U2kDGPyFu+41VX860nzkjM
cxx9OL8qJ7ns2/Po4Rba38IHgFxPNaCp7uneaRF9vE8Vy4tJhqg9iUaH1LvBxxtGzD/TlQ4XUbH4
GEVaXqmk3wfntUAkOLT9/AryrAgsGvpsbfHhdQJ7b+PspEmzpU6VAPyzOa3mD/Uo51e39Ooeyfmo
PzvQHGWEW0o2w0ruvo8pLoakLN88eOgi5zPRlWpv+l0Bm0qN9teflMLL4HeKQHq2V21iyoLw5sjf
xLOtl79oQ75K86+ih6LayjCFrS/r84mgN9erc6s8wwny6vTr8idvSZgOnIRAm5+ixUtKRV0DCnLG
owjOVnhTj4PyaDPOFNOxFELs8QkRfHmLAZGLLl9GiqB151nl1Jv6wfMaLOaUW55iZK8OVDzo1Xz/
IErtxIf1qtFYArC8UHhGM9wYH1sxYldk8ef7xobP/Q10Zee/HnZJpeSemW3HZVIZD9pUnZxL/1K4
9FXJcpAxOCQEmSHd4u3Ud1StaCMhACW7rhEB6bsCGNPDG9b/VJGyxLo58JmJVI0t4qD3osFprHa7
+7S1zkyuQUPBx0p4yZSyBItZMqxWCWLU1BW2bD4GW7c0/0llF9SHdHhFpS/fSCcPcwBVRDIssSVz
mpMsv/DjiG6g56DdufLMhREbPRhIP0aQtfrfKInsm5KioNfUDM7AdY3dwWWayc9d7gGxfJ9pOwjA
USF8s/BsB8A9tvTezxUvBiGm4D22bXhfuFvHGEV9vq16TG9BQHvRbTR5g5dMDFOdm8QpQrdI5hFx
qPbLxVCnCS3JHgEObSAyMOSp+azJSPXqI7QFWYeEkY+8aF1bSGV1GXnxJ7Ir+vMK2noSeICqCu/S
8DUu8KLL7UDOuvMP0Jttj0FN3erV8iuaYPNEs18GxFB5UEqiqyuKoafVyMzxkZjCPkHbjHUTF6nm
Qc37n/FoPFHD7gSthPkqJjZ/sdxwZ6KIkfuSlms/nAPRdVdWKMGb0Ij+eiHACgpiiztav8esYmoF
WiEsa9hzt7A/uKOXCTyR1Svv4PWS2+YnvKVjx9eZkBfUg4wer7oVXKwW7oH/KV438vyYlk+gDrwN
fFPMY1yn+HNGxdOz3BjuD/Ewz5ZXCfOuDqkGQEr9xaprxBmA9NJxeQDZMpcwa//wetUy9qggLFA1
RKBpDq0apDNL6JSmNkQZha2+0tvPojGDVY10t6xkI23rABrB4jRJTvrqbp7Xn7HcqhaKr005v6Xs
g4mEUnpEYPKucHcmcZHA4PYwjaZh90GR3CJNTa8hr0UOlOanC6sNc4nMBErs22u/dMZ9Bfb4Fz6l
h/E7BaRTqAg3iP50Zwa3gG1TNCmXsqKk2uCd+ZbCYynexmFQgLOWa2LBQWRfsbDzbbxKuT0WtSL4
h6UnmWmD5PRDtS3ME19iQGcuj9fbsPaUnkhLjuVk/MuR3zy/WhnK75zl7rlVue1bLWN4LPcA5d3y
LijphtPcbbhR2b/dhTuZb4MX5oY3QKqPLGWgV+xCK8w0fZEVyFyRGU9rhl7CxIa6Mn4x7/Djku6Y
AmR5OHoFzcJsG5iJrKWJEf+NPRsDK0wrg5Eivm+dtmNQ4mfDQ8rRbDirxrPIlwOtGnMQ2ZtRRRYX
uE212SmN8YwBnuSU6k2w4f1ip3vPDpkRH5UgoXpIr2wuMr1AospczNgj/m2NSzGhK8qwQ9Mswb6v
RyfJG2mVTNrpfpvAozwbX+0WsX3ESVcUCfi/gBw4uD9vCieUITsCgaaNmwyzhKibINLC8n6h7Jso
TkonLX5AzE+Du0cVcr+lNSHr0oAOjZ2236LmBCKBBhvVfOV5FwGrjtworp6X0ayeFZsBhENIaaCX
1RkENLLCv7oRXcLIU9fljhkP5tDFsBS4hUaLBeXaFBQ0+MoDIuPlnsGz88lgPOgBp/JQ1cKDF5zo
P8oV9q2RHPmzcaeMSwtt1/IcceQkwpPxRugVcHBh6gBjoR6G25XKutHAR+pZjVgKJCKpR+oOzNKE
4Z+c/u1invqdcLHjpFgGLGbShrWT7FM33fSIaoixEGMRICWHGAB57Vl1teklaIDRwH8h+AJiHPLN
t5dLlF+O2nNkYF2QiFD2VUKRVU6FP+cx1CLQ4hl6zPqWwUkft5we/6Cj/g/G7grwt3fS8tPB8E/7
88rzBsapcN6NaYgIXp7GQ284d3JtCQOdLFT7tpUJi+UMnkGy6DNzprIAcZz+Pf8VqETWZ6bhAJFw
/5YGVwWoDQDajq1K7UZACERWiJtGWr65Ju04eIeVxOqOh2i0+sQ06MmjhJCO+ims1iKVeYYvn63t
DQq5miYr04yxbLRHFj0ERTDeZpUPSdlJnuwnuPyXmq2db0WTX/ptqt83Z/dfeCJv8xdX79T83Xvc
7kPVS4oPxPxg4aZvizVUta74LXAd6+F+d67IYFgeCh0ib764ijRgTLIsUddchVQo9e+mWYZa8/54
tC10V5VtKoZY1xutDYbxOgzYP3VoeUqCHkwiVcFFctKGEQ3p34C1QVLllH7cKkhopSinXC7ldeSW
Nth1UAfIk3I8iopKYG9wBjI9PhZ40fZBFloD5ae4SMN9TGOxFHL7tW6+kNujFaVj4ffDRxhxGno3
2zBWGxxfLExMfvRNSACgI2S96HrlXF7pJaYeVm+cD1sxyMwR8nuUo+SKjCfqUGc5gq6jYwRim8mV
em2M6dcsMMUYiRwbMBuvDfcWsCvBuaRoIiQFaHf5Nz57fu6lozFKgNUb+kioE7awTZO2Inu9+IkK
ivis733rAjxNgj7cc9ftyJKgrA6SSwvjTtpHzw+9rnWBe81IsRY3hz07oxot13ueRlbBm9/xTQLA
hiLUi++SdLuObUrzPJ3vGA6qrCRnAXophexTzlSh0X8k9XMu+HStDchW0v6JpA1qzPBb9nbtnoUO
PpOa9UG50c+KB3ZkoQTvEnBVRHMl/YxjG4iYrXpPxpo0A41+eQTmDn/LA8cmg5HkMxFUBoakLxpa
NcGs2C+NVanBZdpBJHJR3GAe32yG9zxAsYtmgVm3TyS10xS4yka1CTHe7u6y/5brxBD4fdWT76Ih
C/+AfrnDNq5mp1o7K1vWiZL0gjGInK90Z0K3CxVUTnFdTtHkigbIsPOK9seqeCfgE9gsab3u0WIe
u6FAYuh72QfQi4VXqeF9+rFrF7jrzUB6lXLxlfXQpF9YEvUgfjrb6tsfhNfT2Pu58ouyTSiOZvPu
/ARwIT2KrtOpOmPbqr2aHr6DH2fx0XOkp1m1GVhkNvBKuULpptVTO+YgfuV8IePScQngwHLbkavC
mwYUEqIeag1yhsCYwHf4Y7wO9gltkcdPPQ7bzHDz5SIEjpWPxfVez+RmJuUA/WV2BcQ5uDG9/nqW
BLdoO/HT1jH89j3l2ld6Vz23nizEw4GL4LJyVczDXEr78vtKT1PJMDH6Lcd+WL+DOBgrUuOPLdHx
OvV/ylA4SpQf4/LXvXOFj9swXaCqlysjh0n+vl9lJ3e+iw6y6aImDdCQBj8wkG4v6c81U9tLxAJX
0+qYE+FTfSHmJdfg/plhdcWKYkb4Qc1NhEPx5E2yNBw4y0ZYpDSOO6/Dz4Ew4HPX0raeoD20O10l
JoPDIzWqePAC6+gTZ2efWp2bpPPZe/IrKCFyT27fmK+E85gsnWfSHxoFxP2WQG/XiQKb/zBNMX6K
N8Xp4L3NSAczWegWeh3W9cjRobY0JrGw/gmPRBUwb5BJxzbOxSN66svUI980zIupXp768McNWodF
2hMbcvkQmv1kZygzLczV/ahy8nSkpj6t8DVRQgHkry296cV7A5sVPBRgXJw6skghDQ2S1aARMSAf
fbJgIHrhyOmgRJSMlRB3ncx3OMX8XiV9bUtmAX6a6PmU5OPbKp/QxFC7UTsy+fobsZK1KDnLxCGe
P08k1HVy8ON+EZdUHc63ubePy0UvXtSeRaggTH2wqYeT+PUl/lHt75nMIhniw8wvwSsFIRqjc1Fq
U96nC2c6UklUYsFoh2IoqpFB2LI05auuj0mTMwNzXupAUMpX1t0OVLNsJ1+SSRGU31H9xce5kWzN
hV6VLcGLFwLXt7emM9WPHjCoW4Z4et4jXSe/kGI2yxjGsfxHKZ5+ZQFHuwkMDS8Sx1eYRCH5HAPj
zH9/2ifgs4SAti8wz6peNXTvaKtctFVMkH12zv8jzpHePKs8WLvxbIbfKRLpRtogUo0gErlhRN8Y
3I5aDT2qqo6sEzBwjdNKKiwQehpD11QDhm2GKYSyy5uoox//QOgIl6TzaT+vt67Jm0c0hFgMBKLE
ZYP8sKT8wgbFWYYm3k/b47Kfi2LSNEzI/67IH+p5Xh8fUTyKpHSsPnKFPztSJ9P4rQnyLiSTDK/3
nsdT793mLySVplnH3/C7e4e0ZtwG1qlaKwUZPfhW4u88vtsGxYNJZwgUZ/LS/eZEsiwgmbgnbp7A
EpB4E3VGsxqdMz1YxP5gzov8VBd+mpZIno4BpWO8GRqUgvWA5SwM+mTW5ALVP94mFwKf7GKBqia9
VTg5Zk1ZUDJZpr0XXIpGtpCFakMRkIBaooubZr9R+gU7BDRfdfWwNWmD0tdWOONnI1RpR7V6mhwo
ArrFgE16KtkaFWqsZ0h/80bzgYeWXKLbKZPDEyOvjnmDF1nNZR56b3E4QVrw1xfLfQRQFomHIWQU
9CtpnhnOFW7kHWtWTLElQF87WPtUQvZcP8ZWW7UbSQ64WcBsPKDxp6uJjLufDq29If7Ghv3pPp5Y
vIJ2JIyM6TpGJYTXdkRHgzl4uPrz9LtP0g6XilfkoOniSSxXsQMvXx2xnRBqQkDzonG6CexRYgsu
VLCm7hGv3745Z2P87ClKxHHZpH+OYNfpjopFPQNQMBurj6h462dBS1uzmUjne/D7m8q/LcF2WGuy
GwLDQzjeQS+1wQErpuNXQ9TrQdYzPwBPciIefQsWGj1wwDIIvDnX9yLqqG78ssHP7PTrWVDT3uyJ
vQ1tDfs63XkNYFRzeAEKOAQiNKAL1Y5V6p4cgOR/F9jHskHSWxRWfIePKXG9ncZTicx0SgmZbLHH
tMLE5OG9usoLzFlxMSFxpfnMI0Dl/TGXmkU/+ojyqIZROE38ky0tlMWWZ3V+IUPpz6ttPiLeIZXB
cbagzVGtlEdp1bBSn6qbAYiDYwxcq69H598ztZlFgCmXJpTXBZAsCUXZfmX1dyACmMiCyNV3VWQN
z1vY9uw3b3F2++G8E1p+GYhFtuuegKZXheAgeCOckMT7PEdlA0E4h5fqrIhiu9sm+jUJx8MdKo00
zfeCcGZZMUg3zOXfLqcCpB3qbT/P523jZmWrW1O38//LrfWd3JFcOp2px9YFCfb+R7yulNQLx1tC
eGVBuAR0j6b1lDgdk+8BwnaTzPXGwku+6tsUEO1PZEpWExFkR9yTljuLUNaofclE/y66x9L+8V9e
b/ciIbk3wBfPzmmujzo5v7SyVxqqfy+uGryiWvq2KFWMq64TIUvX3A6GTPA3uFFC3UL8LvMrJbcb
aDT19bmCzuwmDR5Y7NABjosGp+HSRn+qa4rG/ifLnfwQNLdICxUjaOZLeyYLBVtZJl3mxIUiDqAS
u3xrMwrP0w2jGNnzQ+caoPyTZNTLXsTZLtOMbynCDXQZ/rSROMJSbmAKM2SFhXHvwrwMK13nWbfB
VBCve+RlXcHBw1Mj4MkEisypOA/cHcdqVQk5LnY+5A7VuRIwHtx/V3VsveFE9CgwAEQIHxVW7UmW
TN9ZHfKxl9AxcO1eDDX5/mOqCD+rPv/L7V59YOwcAhrx/3YtBauYuC8TF5mTHgfQIrPJq22J4SBE
J9YPkU/3ME2OAM7zhWFMAr2tR4JpzEws9h7TgHO8Ze40FXeWQd46UvWnkKCflB9qZ6s77RLYFDef
nNxXx4NpA8sPGnGrCKLfxSR0j0F7aljPA69DlKyPgZIfXpsxUc5e7EYGdkHdbwafT2fy8JG9p96I
rmhLJlv4mMBwDv787N0U9N62Ln/mH4jxzL9HDD2JgjwW2257CHkOBr17zNKBn0NR0v2CQXDxE3Kh
AQgugAmdRGSn6BNsn+yw3j/h/wLkmSOTc4lXG/DuDeYpM+2bilim4IAA+e4uk4YrQ1l/E3pidtV4
UxhWwkVJvA1iqMRXpoSJuz4RzAwUEINKBf5fEUMPxN/NImYf+GQ2pLHlUe3Qgl9XCDSRq6+SB4qE
pXfAjEvN9Ixk96Gxh2nw11UIeZTW9NneS78nLFLE99MWtYYm0S1XAJa28Cfxzz6QF7faRO+Jewmg
vZlacguI1PpInC5uwpgTptGTQNEWD1qceGfditAZYQEoI3iT1GcWMZSuGz1MjKT9IKqPoURUxnFA
cUr28BvrTex5ik9UCYWShOmeTPynnXLDXW3sDMPvu5WVvvnHeRGQrR/PlsA4Kniz3uGOtFMpz2IG
09Ip4knriQ+WCqKNTwqa5tcoza6uyIGFPfh6d/2TcWSF0ePJRxhvuoJITxGi/8B+xRK6g8ZqfHtt
mMN2wgR0fkeP+P/tH15at2I9C4Eo4C2d4DjqnWo+v7Qo9dSPLOoo+5r1H34ZegCsBK8wXO4swn4C
ZKQA+6Odj+Dy+o0W/y0tlOy6nNiOthvdCLmSAB88dXMx1QkwtbYvzhlXU+l+ZdJ5XjetkdRrIgo9
ekDcTo9cuylMfZAPeZk+PV0UlUhppCn75z5hUDDfvdgLIPcItpyTuw7pzhOOVASMgaDNQCxKs41B
bz+c1zaM8nrYfaM+f9LzT9R82g0ATnaRm0wPbpgkGDl8vI0gWxF61O0LAOu+Jh4Sa6mmaUNiEi+e
3yiOnscM2D1OtMQbqdE4iPOKQwskDKiQinsP/nH5q0VuqanNLbeG/An2/1oiHVh0RFo9f0cTgFT/
57JLogfM0DhEiN7vT4Ss0/8RpEAjNtUHXhIyy9TVkOA1cYmR/S1aPDyQ/mzSXwLy6M0gi4aFRv6W
izSyo2zPxSg9MHtKZAvIGsEbbQk6UfZyd3x/+as4i9/qq3JgbAgo0Ph/NHFaZFvzucR6DskcEG6u
61gHWZSWHVs2kDxxzVu62My1Es25cXVpJOXwtjNeyrps0Gorfbr0DUp9lLWR/St27C2PmeZl0J2R
Uj/hbtNsIiTs58hZ9fNH7yb13JdSLv1C9rVXcIMPmHjYhIrOwZs1TBM5EZEjh++nYgcGlFbGajBi
T+ZUud/0j8CPhQWBjpUHqsouBJtWQmUQ+kI/dk+Uat8g0bsgLLSzjA7NtyNUHLBxQOP0w1xYFW2J
L2fMxAC+9ib7UTJdX4DlJR6/cNgyN75NB8HsQIZ9u5uf0op3QSERgGoYEBNjmmqJgAih1hRR1F5/
f249ixzKIePOUGtKNm31t2CHLVURLJU/jUnaE5h6LOedSQldayS5CPz+J0GlRH7Ogpx7BXrVgBX3
tl9ZOzThxlhlolE7X8tLgcxMdUjR2d0lbaY+Jcth1e7xG64lyAx8/NSh2Lrkn29dyfaRXUmteoeY
Bc2tcxdk+WRSQxwMuuZTjDBChDRa1r2kXZSPzxgtV3D8+XGi1ljGBPuhtUZqOWOZsW7Esd9KJtU/
dy8XKKCc7vdgY4mdgC674kwLhBGbRDT+2RU58gIWtPMwaZ6xb6vrsUKBcvk1FrJvF0Z7Ix7ahLaL
LvKFjSnz35b14nPduLjyLCggtjvphSHib0PHQFdw+aQC5y6cs5Tqe3ZZ7FV6XSFFT6GHDMifEEOl
ZxeyQVNKYK3Ahai6ZShU6YUoTmHjYC19m1eqwNVFbpCH7ImGIa1jO41ClVtHLB4vP2cVWCOpUULC
uIAHcU8XfEkdAniMn29v3DTlEjlv6pVfUcBx1g6u8KMk7Gb5PHJbC3HsYFxz+JHOrupTIbjKzHvY
ayEYvI8W3yy23hJ9eEbKQrbiH1vEroW4buDzNVA54FC2/9TK2Fwc/3JoQjTPsL5VcUKKJ/zgJ3hz
qNXmI36myynN4YGT10O9BauNFj6yCLgXFwZ/Lou5gxbhW02pMM6mH1PwwUNgTDr6ZhCmq66ZH/Yy
Kf+rlmeIkQrg+0CU5HQ2SOjpUWzjQGhc7bHSCTvcfcs7qCRvjdBGmKYhvNh1hpoaiai6f41/SPTt
+RZWNhMHk2RHhhKjLOQGzn7RhMjHydFgqr0LqWkoLFYfgMtj+7qXTd69QUSwcn7UPKo6p17Q4i3p
buhs/SzUdvzYCMf9QRDt3Oa27VQQesjAiMWmAgLN9Y9NKzADANzQWmrdcOsl8JmUJG/XIkGApGXM
wl7ZxltrfaiEjhi//arpAYF0tVA7i3wC/nduM4/QS1IshntELpUGz8iabT2Zot4pQ7ihq9g6vtBE
TOGBxcI812vGroOzNMMKoww8PVNIwt6SRSyFzm9Qli3hBdafGvx1LYmnzEMTqJjo0eokEQxUO6ER
zvv1Aak+gzO0kLV/VOrLY/nth7UBSIQIbHoW4c/grbfvrN/l9fsFcb0SCu3cx7/86c3zAqGM8znG
LyXRHjkb1lZL2yPlPY2V+SxkTbgMjBN6fdtPX/ADQ/Y3PkPszXiFVUn44EMa6gdAaj8VS9lm3GNG
sksk+tR91LrDgimA9pB8nEE2eRs0hU//WrqzsiIIKTkAe4pTEHiBLY4XRhvYt/8nGEWUtm1ze52R
Mi6IwIsJPjIz9sKJksmDcss8kn+LhUnc0f4UpD9PC8wMa015jFEW3cL6s1WMzJI0XdargfgAI9Ec
EsumjXe3U4f5w3G/hr8UH0/CxVUkbQIDkLf7/QReSNE4tJQkgfKoX2tnht1p6EvTJXVdQg/msqQj
4XJovlx4DLKSpLaBLyMYg1TTt+SjG7TMp0+HMMAH6NcwSoheGYhtuSDGPpSJAIGD/vkcDVfSntdx
jFFVIZeBbkolhu14WACs0FWCOtT+UBGP+74uD8l7Xt2u2onnYQsJkQ+Q5J6Qs34wBklkljlec8fX
cnF9d/lf1CvfCOXwebLWnn1xhscOb1zY8hYfyQr2eIVrrtefoORtpjrPT45R068WiMGZJJKejhJl
dBVPGsoNUb2uExZzPYn3+eBYpxPhDOTXL7PcJJVni67mEQBKA2QMOXkuH5lke3HKJXYgSXfdv0Zv
k014lxPNq0ia1FkA1he25O1oQfX/iqCkrALnhqM7JrEs9kg4OtVOo3ZCNlfJEnNelETOkWTKclzo
lrbW+5gRAxPeX6JDn7IZeFGAWZ+NO0XOsSD3dFxEzcs7CSXFikwk+o11nYb87bOQ0pmQNh4cSz2q
y7Hv5I8SuD+DY82FHagRM9+HjsOasC52MSZg4SBkguOL4azfCosEm0omAGclw3KQs71TNqXPq54z
g9cBL71XIRTXyQXCstZFcTMfLTg4eJpCau9UDVpP9et0RUKibuzjjqh1L8bxOBR3rCAKpQUH6iHE
Skho7CJMcOL55jg6tqeohgaG6OqItTUs10g/4dIxVhzHqExFHxe9WcJ30Uz59U91G/KoR/JGnGBl
/qb5Oq/hut8OL/2ogJ8DF4Ql7rnU/MZcD/z5O+uzeml0e3R9iwh2NvMF5Y4zM1q/vgzGSahzBbk1
dOAiZnt28IOQM80WBn73oaiSsvUVAkdHV505db4bi2D10wjoHwyFKdhZf/HCxi1EkOZ/UMWh7DKj
VmKVser5XC8Cc/ofr7c97xY2vk/1t1HlT3MxLcgT9hhdR2B/FFITZTrAQxzga+INV2sGupIWaa+Q
bEm413erDfEjjXg3snTfUIBLRW/IEaKiGJTu/zgBn7MBD50LWgO3Qd7EOWATE/xOvY67TO6aiATn
BJUf2IMS6YjSPLj8DOorr/c4jPfAOjXvhwFlymL1xQjups36ZYH/pe6w23Pi4bIwvoD5zp0fOs85
n4iSVoexzScFP5GgC41ws6+T+QAZ/eRRqW04tv1HLXauzKWH1+bwhraGqrWmHNqaDrajcDL2wjYR
D5Qm0/FPMD2h6etlolV5ltNIf6uzmEAd+vGbQIBfnUIheji0W7snFkiGVm0+poH7x/I1DZNfJGLd
voNKf+2q+ljCdTyHiytUcS6a/iMt7CbqP57PEQ0KWG2eLREjlyQHg7skJ+wipCtzYx7WHP1MaRz8
lD4Ll4DPqieUEVK4/m0UCtDwCNGak+jVzjKCRBv8f2Y1ab6AcYpYp+cC+vaMZbncnLGFdRYOZHsA
KMN41NjBxrwA820Myg29f4wjHPrlOFo1HgVDAEg0Xf85yJwY77Qot6aVhDvvrpI2MKfgU86g7dOX
g16QBtYu28eE81H369MKy09eL7SqA4ZesAnp41I/+nfLGvf1ciB1EgqNm6kdtgeEY4JXLoUUtLzF
EdbBDlqBc5mSnDwuTW5tqFgg0ximCiYHai4K+M4u8HCWIW9125qmVlv4tav5NZIO2JxnVTr4q0e9
wMuOfZiJaHbQxaHzcaaYKec7meFr6Iqi4IhGBu0phjntM3b7JLCuOFL3mGCujY/1ih9WaIIMmPWL
fT8PRzW06E3puLQXrBgyq8Ia770j6PyHWikP2FuskiuIM1y3gYHRqg+Z5Lg9tTZ706vNfhsRj146
49kYv9Q6PlXpqsOdU7z1j9K7pXzB3OgWe2SQQ4UtsP+T0HDYukBTnJTBZVRZLGv1crHSfIKhWz5o
TluDDI3zbdSOZh7PkuFQcTsxVlcZ/StfpmGWzxDvh7bBcxfEyNm7u/AiKn+61kemM3gG0yo3jqO+
AUKKMIxNojNLqTuoQL1bfPnCZaPRRK8C/Nk1EKP26FjKllrXud2CAHu90fVjcqTH4lvhUeAlEEwp
edibwP6hIoFXgZ77lCxSYA4hHlD0ThACqvukb4cSj4qUZnItzx8qe5/Q8fiEMfmIOBkM2MywLGhR
gQx1R5CcOVlqNn1QlrH2VEtNCnlB13agD0YHv96/Omq8vT3NLOQixEyw9AM+8BYzngMWXVq+bcTd
Q2jvAB+vjrSENTGOpUN+UcEPk0Ne5jLCex8g+vz2LmNg99lSE7svlYEFeVGPDeYqrBJe1UXDqAwW
XwZMTLDOtzrqusB1EhoiSXcQ+U6xWef7giKcU3WAdzHia1cmPSxR9uFURp5ssHqiLtJgmo1+KEDQ
Dqc6S424828DGkl0BoV3zZ09uIMP6li5QqB0ZkYQipTe0dZf0yWC1nvB9mrD7PceXYnIbeKUEHhg
PCr2cswj1Lm8XBYyfoGZHJAU2NSdyYTeT5AJerG/55y6MK9Yjw0JBw4hzB5ifthCjYFHq7WPOv1y
TnYSlPVTFWK7/83EWh5ct3yZU9NfESZE+TKzG6IzpGdpnhoD8oxsjZlU17Fev8XVNRGYMF9PgMlK
xZYJuiicZm+fmC8P8RevP45340j4jzKVCGWIBhVUHr7EYCl3H6sDSRZonm8+o2TqKW7k0J7c+YnS
RR0nquaOk2+1OtrslhrEE6XeCbY99oRxi4uMOj1u94M14GD9n04t9LtLGYD3ZEow+Qb3GbhEd1Mi
8Nm2H0jfYT46bkNuxKYdGForlmRa/2uDDVyisDFXsLzN/7B/2guWKU0DL5JaIwcVpCHj2GmhnB6L
WP1/RDwDSZDW364n4M11S/aIOxhqP1mssppwHnNFoBhIOtbdksiNjWc5vfRjTLcI9gkAjB7SCH0i
mADPY086x04zQZ1XjkY0drlEUvrq1dLRT0yhRtoBZtnaRgd0Ce2Ym4/naMGthC7dikkvCscRPdmH
GeIuzXB3GZjuHBZWyMO6IK573FNWzqKJPjofCuYYwwQcW3jsVDZO6wQHASC9WfF82N4g8M+kVRmZ
OUyk6QWcTo4UAyu+mGkPtUD25xxlBJpho+/MpjsKmHSzOJxalBFsX8AoAGY9Rktw/3CO5hkWXZHw
qgzzUGwifGTLcJYS/cl4ZaZpIsPler4dzf/KMOoW7fUrfKzt5MxQLwQMIgdA28DMqb9CmPKp6HpC
ALVcYcJJNgKEiOJ4utz9R3d8UzjyL130z7hE/Ijdnsk9oOa3ZvH0608WCQ9N5Cg2i0YrPMDeTQVg
xJMwvH5nCXUyRZUKRMd93smoY2BDtlA7/MI0Mdbjlzfc3aaMzZw4b+0uGX1zp1+sUHiInrmDoZv1
hqzuFV5TfaGa0rZF9+81N9d8RrGMo9f899kZ5gYRUwgsn8mHdINKWNmflsZ/BvSSNFmjCXyFovo7
8pi6jJTN2Ggs9brpsVLuS3IOp6l45zjotCeczh+vckRHdvlrURlsNmQogStM2ntXX3qDQvofWYxa
ejQhhVSwOoubEwZhj7tC/zLGsiG69fUIhIEgRlS6vYrNBjxqYf6olSPuMLiIroPdusOjNVTdgNQu
L3kqE4ceuJQoDgmewb/R6DIC8CGDIUzXvW9VzWZPCzuOJxpHR+QEu32T+OzaxOLRUJSOaJP2T8Ca
EMRKOyfBZaznwzhLzIzJLD0c2GeecY/Gpt9VLSqTKcGqDKDlsWQ3IHH7x23ct1xi3chGg84HQN24
OFXu5atUA59up/G84Hzwlod5SlCwDTg6lSJlxwImMmbo9vHpGRg8rqj5xJ6WwB+WVpBFf9xR3o4s
ZtFE3NO/dqb6Sny1qGQYlrFhbOj08t1epm4mSHlU11SIq8QPFRefFCj5+tUbamwYnzH6htutvc0c
ugz6p0iZATufTtaS7dWhJFBKiEUOACqOK/+zVGaYp8H0X+MfPV8ciEDPpYDol/j+9RRin0wDnR/r
aG3FSZtaf3zi32HUEmfSJSXZyzpjbPlRc5WVVUpOSKxuuyTOYEDbgsVGgrdlR+/C3eqEN2P0LuNc
Un9p3JYJuCp2gPzPPC/Jihc1hJWvqd2AolRWvX4Gwg6UvnLWvbMlisJqeLjPdia+jsjTrUqYgIHC
xxjXBsbQ+hovjx+myoLxIcyuHkLSftA/CbehkpbKifQ5r0PlZr4UmUSrB96nSyIVtSFTrOfzCVJ0
alisHzMbbrKnMxko4CriAIghvGG5+mbAYCBGL/BZT9J5P4b3Kxkasd89swyiBpQye6XZWp4xyjtU
+8nZVLg+eSBJdT15JXTDHp5YaqxqH3A49sIj0Ip/UTNzpgh134iwZQIKjZa0gM5+H6FFbEGjV1Bb
ogfLwZyF2drjMDY4HTyd1iqiWjTSzMp4zpep0x32FXFDaC/c7nnO+/z3zGW4aiM325T3hDsNx2+0
8JpTN5lNDcxUZ7NApExMjs75Saxh/NqVeweJXiogG8x2udbve9LTn9VuwwHAeVEk3L6jqZVOt8On
/yNQSMwOTBVP9X8cm58blXc2ETvVmolPeMe1USH88Hv6+kC5W+4HhBHOYiB/2Vq1KZCurmc/h6WH
isg0d8LfCiSog4kE5KnUuy5ePP5YQlN7wxWQRf5wy8i+5TjvGxRa5viFxir1O/FFXJDrBV61LUNv
L8iAmdHvi7GqBratUWrwrAWbwDaXDNsaItfpyDKLqWQU8uULHhyOU0aKC976NsC1Hg94km9FbjOH
KtzzyAkb7wUxXV4XPd5pBCHd42h4GBEC5Gr1lPS4Ea5/Nf9DF11MLeS136F42Tcyr+nIm7bLVdNZ
mBHtzBUNtZUAcxigjhTRuHIsKC5mggKcbYzp5bec+BuIH5gYP8yTOIxZ/mbk/wPFWnHAKKxKh6Nj
zhrXW+YouXVk8ImEAVMsJ9Kyvpn7blMCXUUdXGDBx0JQnC98ekERR0WY0ejWbmG74JTYymUgdt0I
0nIe4TxNl+FuSN5qDiFNdVpEckOkyC4QHaQOi+YwpcGbBvquebvvyz9BThM1tXbRtj+FpCM03ALy
DQ+HaCaEHXfcoOif9Cf2G+/euli5dXt3jk+inA8R4/brHGp4dMMMN2yw9h6rma23JIPDm7q390M3
MJDTdY3DGbQIZBUxCIx9bqneeW/z/P1GjaABR7WLk3p/yRxUgksTee2pfgwc5t4v30kVhlU8baf1
XMUIS/cZZJOxBNyZvIgUFwDt5FIruzWoBSEBZOXw33vLnGgn1mBR/7z7xRQCem8sKl/2kN+QfdJa
IllypZQfRuJnCS2ldHc22MFUDZX7x+H8badfTXBwXcXwL8fo/l7PGApohd6hp/Gb9CgUCSBT+lWK
1JvQmbz2HU5PiFnTjs3DwSk7DGT60h/6slUpOH7a5vjxdmji9CqLbRa/8GHWKGJ1Nr3Ws2WXZObb
pxnMXhzgXQUffjopW7j1w48gZJzS9rKA4zQqjDMIDnBl2v9YuBytWnjCxSNSdlgLO1vQJ2JNez3W
OI9WvdEFkqVhMKLsZz0GvpFWx2n8C6r9zbGUpxF2sKHcZcza6hGW3enQ96BTPvOmWmEQmzz6QcVA
RHq/TjuMA/cTFyjg40AwE0vqsNWwpsFpAENP5RtwOPukSfOQhc66nnmMQatdTFG5/ITdcZas5B/z
7bsYk42wOisOksNJ1jIFg80LqAq7GgbgibxjIFOTvpmmE6EfcHJt7dUitCjJDa/KjK7H9O97fx1E
a7OrHQDRgjSSAR7ouW+ELh8AsDoD5HRmFt2HaSM0AaLpSTFRY0TPSpe0wzQxeXvYJ1cOgYARJMXY
O3xB1UTQ4SkyFBq5+cKRsDcpXKNVbYk2S5XpO6lVMNbiUHqd/rvMqRwmalNHkd9O/2JIeoCrIbVg
UszNSJC77vaBrUzwBIemY5wB87s+RsYGI0e5YpK67DtHydE+hN85909NmELGADVqqKsTywBOoV7J
h7sfLP8hphBGX1n563o4m47ZE8bHiEuu2vZcqNHdojEDWYkcVC5x8cBIpelvc6IJW64QXJBJw98u
Lqv6HTNeOVh/kiSYbRCpfvK4cqwsbqknk+/dZPdk+54fMJTl5ACnIneDYZ6wIf/qXSd5ZpHTWRY+
HyLtJpuqCfzdQ7rRvU0kr/1bUHAJ35XpS9yWvNyV1Z5JkacJ5HEymJaPVbLpHD+VGIWesxjQdEnL
ap+8jnykdEp4cVUp7+NYDpUluR+lj41hj6ziPCtklQm7agdI0i5R3feKpXu7E1uIBL2eKUBX0Z6S
inBJopCE5oTbOm2gdUcJDvICNIVaDgAGoU+LHYplNKWmuqgSPs7zixVASTGfe2APYM15/BQ4ocaM
IQQacpQ83MiXX0pvXZe5m1WV77vqF4BQdUdqJLLXSpiWt0hdiPZG/i39eZSdxdaJ5n4tAw01hQWR
VkmFm8nKGDVn6q0VENZDEO01S5J5l7/0XcNdAYwslYV3fOW9bXrBfLr1QN1I58wlCar8OyoEyfmc
wkQU1hVt4zyLV2XhJ5fdyFE2Qf3srbQU2kUITQV2e2PP0Zoru29i6gq4+LShBcyYaYAQwfHuE0gw
NxYSAPabwtgsqOEKrJfzthLeRcU+DIUgfS7UuWCBjvGPBE66o69Y8woTdCDEfJQNFeEM1+3cq1jH
WkFcqKLrcskhMGouHYMI03PvySaMr3LJfO9pQD0eMPlUjQPt/qWd2BKrVmPG47UTho5fFUj+/TdH
mkI59gpOkNVBMc6B7TpBKygN48LOy4W0S9V6Eh3qJLsQed0DPnsgkZsfzsHj2kajmjSPkU+QoLS5
nQhErnagcNjUBUVVcFj7574+lZ10UeVVZxHh8mv/VyUKD7gvSEn5y6+ZYBDLqBucv7OBiHIkgOr3
Rdsx+6b7M9H2a4UBL9G9BijFT1eyvj4ShHUqT0XcrKKwYlwgZhvU2P6AoJEtYciGtbds/jeytkPG
qZhFpfWtduWZDel16PZkA5zOc49zRkAG+MdhB1DwYGtRl1Ac7npSrGgPj8PCdG4YkcyCWNW5cwum
ilt5RKKcVXnL3rqLJA5W/dBv3S18QeuHxj/P0pWwbJ/uGCd8TyQZwPR5VU3sY4s0GYaVT8ljqXOt
+tNYpuAfvUWVzh8aJi+iFNVZTf7qaWNOZvTvTie6ygWA/2+cbbzr6xPDBDXnFVKnpekLUUfpdhYI
VUJJ/a5xNxJgeHIjdDV/DyGAHUUwlEAt5zvRibWZhp8WxtiwLa7dm4O/8x0Nqk2jXmJeMBm1nTj0
kuCXmvTKgzeJ/lcD/kKUHUco/DI1ucNUwBC9itWK6QrryHFh0mX9O8OklQQRkQIpTD/fHO9E3hfn
/0tOJOBim05rwS7+UgW37gk8q+xkR90zpliIJ6JIbdWZZSMkU+zXWPupLEBKxGuxyfGeyTAnGcdM
gwFzJhQXKmr0BI/b7BEUhGUiKCS9Yw+Uzg7WEz3DSy22hfwgfS7qn5kSh2lPdrEsTz2UdXYW29Hu
0JmHrs+TyYD8cCGjZjKNhJg26pIAmiikD/5vhi7dCcTxZlP/9f0m/FEf/JgQnQTgtT9GqrasMDnf
wObOwrwg0gqvw6N83z25wCE6x7GJK8Agd00j93cp7J7KQkQQGkfRHLipOZOm58zA+AbzJJYpSZB0
HC0mtIu87ecpW0aaIrl+9nYdhYHACROi/hWc/PiAtztQ+CKflGRrKNV+c3sJn104Yq9saHp/H4aT
2Hv3aTo4yjOR6e/6tTFXXnoXrD4/RFMsW3jDRxqQsZ0ixaCTO/EZeKh5R5KA62r8h9gs84DffjQm
VdLirZTCXynSUx5ranexk+kQNOb1jiTRCD3I8FvmWcS+qFtFyovAc0unspLuO/BTo7dZ+7rS2Gjs
UnM2YuwR3zGEJERjR4OPWaWw063meoNBSyClfx7qQNwEYKSVuBjktu+HqsE72pnx+f0Y7yErzBid
WDlQb/HzwggSaZ8e3IwkZQnYTf+K+quq0qeiJj/ipG6TzT765L/7aoHyLlCh6mhqHuvWgMYrWK72
5LYKmHep96DCqbEl12xEN9ejxrgAYOSyrAuY9f8qXg+mstFqfc2DREJSPeTVJogS1KX4WneNQoC/
oV9dyEXox6NqWlhSE/+yavqQQ7Mh+Orb1SRMM5KIUnPKHcOoKPGL+RraeE1fE9z8ZAKYINcv2i5j
EgrPM0Yz3q9U9EC3ThD7Zt1voEUI902bMaOhkoUcS2SIVcjsjn43apHiYAiFpekBw7DAkfbeO1+O
tY2YAiEettpR40svkwoCUy61WS2vtRy9l3zZJ8nPZkJazRKT/6Vg86mZrzdLQUxXmjACIPIsOHg/
heAGluiZnNxwgn7ZRF3yNiWRwiQ1EWwwrNUytFwpktvJuOovedGiHdv/Hjt0HFFlWuLdRgwQei3n
czyzBzBOQ3m3E7s8Alfx47hVfSEWt2hHOEgjIt4DZnIlDSwoZcPX4m6Q9oZhTojZSHCAbuec/67c
HXB3Jtc12WAdPUFUqwIXwMpYITdsTQm4f8HXpqa0rw4uvxfLsaoi4lnlsqW0Tf8nvnAtS/Lcn58j
kh1e/BJq6nB8CCaY23ocQ7/kftxJjP9yc1Gzgs8DhzGtpJk7KiT3V63PsdbdWGjd4siXN1VCXGWg
sjCEzkUXC81aBj582qmzPWrmWiVmW1pEza0jJv2b+FDX7trFMmZcwugzivDvCX9106sDlldpnXdc
sEDw2cFFmeLUmjuemfaP/d+XHNp+oyUDtxJz9vplL86gVwMQAE6xgaSnLmhKWb+RNu1hg4p7YT/C
4jGHIafi8vfprBlsy6EFfR7tJb2lWDG9cCs6JvDGG8SkafJFWxEvJcu6o/cSQVSpcBcv2AbtuauR
0Agway/AlqTaf90MmP6jbwN8bEzH+DByQpLHIVwlQO4MH+gJmM73JH66gbrdiEs1U6iDbYXpTmFy
5O+RPKKmhuL/FdykyOg1rGb/eR/PY67JxSFA0mLGpZNsMx2VVxNu+mR7l54Somh4D42W8Tq0Tzpq
CDJVTkk0NY8OvqQoOZRDEAPgvq24ir5AchO8cykTN0B4FNuVE65DyI9ujqNHgCdHOLJGTjqmPtwz
VFdTfIGAgq6N/b8jord5VylqNQ8G0Px5IoEftuopSx4AIxv+p3uT7sJH0PyN2YdauKMl4lhWO9TO
eGHWhwhqTYQCphvQ13cRcFacsf0XpmXQpSdWOmbe91Ixbxpb13boAKt0Pg/Gryjm+l8Orx3MwaLA
+N6oBfwVgnD7kM3nbYbw0fMTYimdmuREbawBL1v0wvPgdmjZ+Dwlzx4erFkADl3er2taRBW//aah
rNFfmh4Y335QE30aL66L5C729jfqONbo5NBEV7osC3iczubG3CdWTvtG7Wjoiqw2ZX+qBT/565uW
7aGGAObIbdbwYn/tvdvoCEueuWlgx6wbwnbnwz0RvfQEn2hv2PAwYjm06EXP2qt4g0LHnnHvdf0t
M4CIu+y9rKHJ35y5fmyp96qR8cF4zihO69b/2W+rgIWlonOpPfvXnSqtYVpfCxdfDq6WEEktA/ly
XekZmEuvGlN9pnNQE7TlEk8rr22Z3tte+V2CXXKpxBztHEIe3AgB7WOk1xWeiLNNgjJaNeRtJpoS
nx0RU0lhhkPhV29e6ufeIm38mu/hcRmicITwcWRdZTAVQyoAZP/rqjDlD1G+t51lXcM1Ru0OPCM1
3n8kaiGY/MESvIgWHqdcQMRQCel+r+oidxdy+DuEsUP16x94e0vjO6/g9tHCzesv4nltW+Rssre5
PY5dVV8ZgslHAXtMiDvXF2F67Il9Tonqep1zp31E0ICYFCFbo56b2lb0wx4PkMFEilXQzJWODD+k
OYYgjN2O1SH6xLvpFQeOOBetzeqHCzl/0cdD5efHgb/SpQXSBLtLjN8y5p+7mIjyrHbu8KwT0cS4
pUwMJU+FuVsrKX6+8mq+tGlonUm1R8UEFGpgHwqg6Pt7grcn9xg8ozdYyV2Gx6KtSrEe/D/MrIaw
6M6rKVVw3Ywt/VNtjY9CakdZ+nUnlkAcDCIDj/4rf8WjwIh7lgCdEB27bKplYlMEqzIwElAn1tmE
3fjxOH+PYY/vQpM5Y4vBbuGzSnQ7WdfPQGQUIYG/VdPl/plF6V2c9U6DONmcLDXEqcT06w55CtZf
JC9WD42o83K8mkXElB5Mc0ogvjnH7yeoFf3dBKekO28HHPEvvx5LYfqkimpYAT/ITMdA8r1KQyqv
7Hbi++n0fnb2NvjhsbXFLtE5KpRIDx3n/bYgEhdEuxnFc9yvE2Z6VLtXhJR/KXd/JLv2JxAvikHg
RIcXa2NrsDduyM4cdXmbtffuBsO7IOLXY9H5X86NB9HnUQYqU18N38W3Kj3bi8LjWm9Q+sr+HdGz
gyCyLC+QO5cpNJielWS5MfRj2i/M1S5EXlsxLI65QqryxMp9zfyMNVKkz3QxyBU33Wv7gMuxHSJ1
HZKraidOULVLeDnNNzzdkDHp46hwEdp723M+MWPL89/pQ3q4DrovxEJ4MrJdy0/NXQmNRZRRDiPH
0Ifniqu1HC2xEAE8/xlife6XYoGZ8LwAceVYJBGcudN07b5XsZuAcxn8D8KtkOQjYYLxr3k6XVbD
F1IpzYG04OdBqTois9tRri44rBqiX8Eu0xs8KmBsAmSNc7TyP9Dp05kzKkznowzea7La0fL7Vmmm
RHr5HRn498WaVNvypul/sUxMj1P5OZPNSjvROMSKQ+VNG7xSNZbxM71KX1hn4ifO0nuP1/KpllsH
H0bFk0cTW0s1BzGpzEO586fEFXZs9V9CeJv3sEmxQjlm96eYNbobNwFiad6cIPQrve/QirlfKBFk
BWNtRSkeLNMNvT50x9UmDXg9hvQQdkXfQo3yTVvM9LhsuK9A2qG22SXGWdapNjhENaX9+tcGXGn8
dpaeVmrXp2dKJebstVm9LaQKXJpZlpRkZgdiVACAj5A/pPkdGBV+RHlYZU+pkXCAVnlaYuZIKdn5
M9agaVZZi6gE0fTBg3NcVuSlZwfpXbBjKYT1OUSVOhLYrLPawJUsx8BVphT/DaSS2H/3MKbOCwg5
oFOUR58ovxolrSRX2HSOi+O44tHnz3DpenOqh2LWOg9SOip/MzEFeljlhiM5tsv1H24CPYBs7ToP
IMunAralwGHnLjm2+isppFCiis4UB3MKGv1wl9iIMSHp57R09vNeShTxJLH3PIpd9xi7FfYcZqtb
b8qZCr+9PAPNjesQzAOpCVdHR33xsjXsfe5yDT8xAXyU1VKgihwt+7Ye0iQbjcVFm/73tkT9cuBW
juzCxFjCQCijx1NgVSh4inQK/hySg+lYw5MFWqJpjAeaQx7MX52ksxtIzC6PHkmEs0yO3wsqt+WG
zsK0pCLyYBTmryF6GqfLSpAnnLE7VHhD1s6F9TbTR/PFk+gwPblXDIE1QNNu+rTMn8wyM5HS15ax
M6LsAqeK3wBjxD5iw9zNyG03Q5j1ovpEpT0N2lp8yMqZHFrpODagafqox7Oz5/McuvroR5J6jwyp
NOJSkAoM88Imc9/VT9hvpZkvm2h8+2pfG8P2cjbn+n5R1A2fGU8pTrFP3ROF3ehCBT2yP3jzd80G
fiKcLjWmCSiXEuMHVxRmY6wxRW8DppmkhbWYAQGVxQLiKsxjN6a5r0UGxkyawfzI5IpAHfg0aZrW
FsNYTKBS9jRsjcVmIscwUaKlgVfIK81Ujcj+rT46I7wdofeA+0GUpjV9ymNb2IAw32vtsZZKSh8O
wwAO0faN8VMDpaJSCJo71lOi3MEwmYX5OlGaorcxSqjbs5qO9m/ma+ZdSFVVek+iY3pQQPPEr+OD
ztDU9rFEX8FoBh4cetQUkLkQCDMyGMOZEZTF47JibffrSuKJibZmGPZZgKmXGOK9uaekPDx/c7/M
5/S7RGQKadRtc9EaN8xsPEX3Hz6tuhReOn6dli/dBppmFFEaJjKndBVpOYfYr9vu5irotYTi6BIG
KSu6Aa3xftITEFL/Y9Y47ysKE+anwZPUd9hA9PzUi+a7HATstUa7eFzeLrFthLb/SB7LNGB1XOxI
xtRuf/J2ixHYsH6WNPErR3pBFJcldvPyIu2cKSxT9goqWNlj6nnMAIY6EmOwCj6j6WHitbdSdOdN
4A+Iqg8jrRABjf1iPnNPPekVLSnt9uXHTmsIH55yvwaj9kEIoQEAGt/MzC7UeCX6gn+AwTddsOdF
UvsD+FGzrvQ9v+xJ1Xn0Vv1jIFAQgLaSPDs1aU8VdTaQ0Ca3N+u5QvUST4BU4PdahtgBDS3PBOKq
bemSwazDRanIllnJj5ul65Bczk3jm+AuBTLK409K/pTqjojKjeYNbLw65sh605sJcdzMbwdYHp97
MBoq+1TVZi/YUnvd6maHz5grKIr3zc30ZFXxbOGEkufgOBQouXj/gP8UFsjk68NuEWxEzpMq0r09
AzC8C/UDOn5YTdFRBXDFRJDz+3G+Gs4Jm/fPg81k6eCLVCo5f/vGLCTYX5b7dRvcu44F/syIDcNt
oeGNUzENOBjmxjC2eJz0IZ+Icr+JDEUApKC9WzJby8C3TekirhIK9UeRuBVWAofc+PdjWBwkekwL
LlBNx62S8iSTX2n2epMXVCGPiJN3aoI0fYRF6rnxKaLNSc6vkTJcrZvXvLG5Ur5tIp0jLxxSFchv
puYY/oVE2/IDUp6qNgkaT63Rf48LvFVhEeg1VnUiFkLahpIWAwF3FtaUu0nS6HwAgu6HTFJ1zgWl
6KmsrYhiEvHBR9DM2jrma7Zc94CrX4CHZ2m6xhGaioyzBAMFvmyjCW6RAkAhnrkPeWO91BGMuJnc
63fm735Xixvt8wRZUiC53l6ilCxeT1cpGPs4G56n4fJxfPe1/KPNOndsEcneURDym8S7f+du/y3s
4i7PbEYKtWgEWIi4E85LAu5GzkFja6IiBLyh2QU3EwloxqycQbjYvQ1j8DmGmN71enUsQjXBeJ9p
hZzDXQWYWrGpnUgTAH9aDBqqlRvxKSU5jMeYF5fxCRmqO1TelSghEZc2MjrS19eud7TJkU0aSoiX
jXabizwOd8gBNVJKFLFyJ9SsfUiyZv+L/yw4+3JIqTNXE3TKVWKKC2m2Jp649A1uXnrE7Q54xrx0
SY1Plu+jJq1gAHv7tF0Mz0orjhJ+hG8a7zmz5JSvKQ0XJfVIC//cKSOHmQ+0JvGov46BzUhbGAbD
z2nx/ZN/JLOfk4RHlB5oQC2XN5NLsF/f373gvHErOnez2c0nI4kIM5QXADbV7M7VZg5hLjUVrNz0
F1n+TLcpgOm+gWbZhPAJlS13CztLw75II0RHvmBjqUaV0pfkrrw+qkP76ktVtfqQ5N5bcBQRP4sI
kuzwnQ3PTtfy6i00Q3j6zeNdyByIwZ1sWVzAxMuXc9Ecm0gMzzSupno8WUB5n1Gy4yn+2cHXQx3z
ntijR9pGpEA0oe9sT5WXr9kAQBkLcAv+x4yLqEVCzBfeC+wR+pmsL0yx89uSI5urI+KUzgXRUF5H
serWQmgBAm8Psi6foJsjc0DIc2fHfyU/R4Gdyu1AEretRZAGjpz4SCviNJLNUP3qFvw/171N5AZ+
RuZQiHb475XjxdlQzt93PYK9g6VnbB/wmP8/f1yBKVCZXbQufLFBS5fL9cpwrOQDAmIjB15c8qDC
tWG5Bbi9U0ne9w/zq6F5ZbF91xLD9Wn7MFEaAHdu0f7ueq20Qp2ATK/7sSsF2n+JuIsHy6Nz4VuU
HyEihXfx16hCwBOjuS4STqtN1sh4R75ygMLyeNRfEDN07b5+Gsrd/c6pC/rhYi1+mcSFecdOaAwc
r71z/gbajxVjpFMoO6YpRZ61ork60r+1bhXNNtguz9HQt8VwV11QtX4xIttHYlqrr3G91A1K1gab
9OqDHZVnzPe0FB7E0NFr3ULIJQRQlh+pxKcaNlfEAy6SqhbNNGsBkLyUzxMl8nNZF/om3HdDEw17
UWl+a771GrImW/EXdAj0AjUvfIqnN6KMKzi5FBB+La4rRPcIKW0fEIqvn9IU5P9seHH/xC3j3LgE
7SKcU4+bvbqcLydH8WQ29rZc90UfpEXwVzPbPjfz0z0jhMGifQ4taciwuIsjfvEsbtDUZTG9CjIZ
1nRezSi4LOAw/jEuSte6Q6+tf51/OxIYUv2ae/P4wqNM12fjcIWTxx+4HUGAailIor1/7mgssKwl
HrlA5Kf9zMXXA4UKWu5NC5bs8c4ZR3GNe9YbDzd48DTi/WLAQ+nZHoeKc+aPwKPJ3EOWdFiOhOtB
wr+8FRAYWtaMvcDR9NUTI3atMbZwHeX2LeI9Uulup02nODWq0rnBgvWhjUcJbRD47gqdgPyfga7T
0+hUM1wCNjAqfw8VtYAILVYeQflkWYjmzwNgjLinna37pAkDM3butlndIV/N+kYIXq3AGrlKwsaR
1IXqwtxLV+X3IhsXNHNZQpndkYpPbA+rFW4SycydmfwJTud+P3Tq8a9easfnXQuX1lXHCs2MyfES
vG8qX8VeYcb/8IPd7fb+Kogq50twz1ViPdZnvt99BOELILDwRWhY5UnKRHDsNzJc9huA3TThv01v
oMWKExcHqgMHqciO5T/WYdcMQs9niTZ69tnfL8tL1AC0eOsWro6rOfdVbjoZcMhb9HWWm1+cyBnN
5c1ptjN7hsQvXumCNb1qcjSgvl4i9tUv/9vUyDW390wm4+cGEAfZcc5NlBDYcvaSenSJxIHYMPVr
qH33SatM6YkQsXkZ1rLKJVT9YKFIrY89n6XtYt7K7l/iN040PQ6vze7y04jCYsI+RIFca6Ulx2yL
ECLb9f6phdmRFe8rXg9UBCtXkQBeU3HIUqYX5isHL9efnsbXlczt6pYD1PaCtK3SUPxUL8L3Yec1
chtERMDX/6GceWSP2hJr7pzk2umYekDDYzAgZKjkvsCNCqQjoEaAadxbAkyYR1+3TDbr6/j3zZoa
gt39pL4BczAXtnLFzfKGdE7kx6uB4hT2mM1cuDSsAj71m1FdNVY0vdOO55oFJk5smvk3AMkM6v+J
phHruxLD7X2syomEr22SMpCrTpCkqVX48PMFGSKi3IqvFUzMR2AMYLKmBJ+uu2DdlR+blikkXMBc
mdoZhIqpUtxiXlAoUAG0iDFIm8Djf/jznG7pXPtKFmZ7Iz5X8XYeoz+MJA+VjdiK25svFtXHtlGz
aCiqCAkXy+Uv5GH4IMFTlpQK55eREOeNkiCoYYmKI3EIjEZWTXWPsKqEt5jM3hVljXv9eAf+zadf
3CdvDcQnrueLwfjBNHX1WVdpcVx69o1R4TLnvJqmYgQyRCBXtYP2UT6PbgvryYcOy6cX8Uy54ggO
luj4keul+GXKywtZxH/u2Cv+9bBCiPv2ouEq0RBHs2at8kRWpdQaTaXs1BCpV73EZQyhoPoGdszu
qoQ8lLdHe6ZEPcOiB32UicXtvvOJ4ZfKki0Zqu7u3+S5SnQjLYfmUJGr3VyaKKxbjAczMCXt/ET1
VMpS8ZVUfFxfloH+tB7mALrNkzJd4iFqYBN/O30PFaByw0DlCYLyM0iKJWRc0drZuDsi9XKGRhvv
+SWK2mGwsKB+oGn3ouz4Z2RVvZBZDPTk6LNbMuOFtGFWq6EsAiluLbbgMudTN3rHNPclRUtjJyEp
UDW40nqDD4BIcvgs10wjJRVPKZdKDSkSs6RrD5ctRF5L0hJCaMAoGiA/gIMXBuJ3UFHSUdCgEUHm
BdCBMgKmFHtohlDsfrSgkmVg6LwR/ikF+PCVR4V5CcMKgHXpLIlPLEkdK+Lo4PLpGx75bS0h4YPV
vJGajfegNPS/d4Gi5i16YhmkjnPX0MipCR8XpFj2efea1beKxP+9/CD8NLdEs7YD6h67DIxke8vW
U074+JWbQZvLR210j2x/qY9Z9MAeWy5RRZ4l306r69zBfzOBm4jlRpGUH/fbGQ3kStS0lPxWXM52
4zrlxQwfp0Fy5ci29L/8rX6AszUcKwvSCe62FqG1b4EdMHk67trgYVwWEErLjNi051xO4tMnP6a0
niNdUVOn/hKe4iwnYX40ejA2jQxkYBTOtw/OoWfpldWEay/YkylTD6VqxJlQKwIDNCrzAE7p+EVg
Z4W43HeSUvnLplpfg6z5BL7224h23vNt/3hh2y10cHDqKDoZBBnpMcb9Vgku95fjsno2FxSG7vZK
fG7F2muVfATDowdtjBzzmh9DVyei886eokGoJMZ6xK5YvBBNOhTupNmR4CNJA7cDFJ9CRcC2zG4L
epMWmAbxvwARlvX6WwPMATb+OAl8PnUXfNY+UJdtUIwIwEPPBX4EdXaMx8Df8sFPCtDpaV+5NmsQ
8bbhqfFbwJW1ztwFQ0p7xN6nVuuPgAzdKBPa8vdfaV8Idj1E0jc2sg1GsJwUP3ucqe57LYJJ7xof
A/nV/+RzTaNDBXMTH4U6AqgKKB/ziVlo5JkFCzHlXD0YqkdFzIpBJO1pYg93RhRx+6H2qeF4UoUT
S4JORGMn4VBHSvDH9VmO3XmfTGbmk7WNQJa4tH4F0fz+y5tb0JuqWfllx5SJb1Cjm+VOfb2IdrE1
tU7G38qlSyPAQMgry//EIsfSD8kcI8AGzp62oW8BCyxd3tIy0I8AbRjWcurhBjf/DUVy01PAOan+
zd4d3w6j1/rw0/mDoBCiYAZMbVihzh4ZoXifj2j6vWJiRjyBa7pUyXiyTuCZnVSX9W0ro5FedWqM
3EUy2vAw09NRJIyKV6dfglDQ80urt0WfoLL310Ko9NYkCL3Euj3AxTvx5TlJt/OuYbbeAsNA/akW
VxKp1gam8ssn1bdF6PYNBzT6t0JqvyOnoOatcO7PGHULDmHNbN880QkInaaUvqfuqH60jIUVa4mb
UQRepJGuUghE+qG6RcuN/7dC/4EbNfoKmqwqk3N9Hfnal17b45Iad5+jZHpRMu3dDdc+2sI68meU
vyAj4EIvysfJil6QKvQ5uGUVMg6fWB2JLZAxasXv5hrzg3w+nOMlxGnm+r42bAzbUQM3qzUNUTn+
GFQbKOsa68Nl1ytf0suUeeEr8TPED6bn1D0hXqlNApe7RYBeXp2cUN1IKk9TfXklXMWqYISxFefL
SojmHqVzkvSonEJQOIFoyV1ATCOGVGXejliqw5NeruuLho5tON5tEHLHlhokFm9ZR6o7JM6lN052
p65PcEQqLnUK0CwzSHaMhnkIjP0t2ad0MLOuoNBISryWQp+FUa+CT/9Cjb+TRWpZeL7juyUTG9Sx
tL0dN+xwKc/ZJAKV2E+Fze+GAOy7gi1cH9o0w8+zWn/7a88ef9nbhSM3L8gyxHV1XelssAjjA4lr
A049rlFaYRohV9zsHm2ElDXucBl/FD1IJaLEfm1DqNBH8wrA+QOsyPq9jwiLW9rBtEjNSMaiZcgM
Y62jFwrGpHK8/+PgrdLzD3KoAmV343T7BBbDyHjxjr3Q4qrJqQkA7QaqlMYqmEEYQ7MQStB0dyfs
YUKmVY+QSQF9K9o2VwIPBk5WVOZUC3jk95nOKiaTm5b26gQ6U5eUSl37izgWBjtgr348kcUbcamv
Kmey/iazn1pfzvfCpuqBle0No9ZJf/5vdktXkHgaOwabMLBZPVvSnX1XJms5jVp93WQ/uHNsfjnh
vM9I7+pXeU1pTb2VyFT63CKul/5h12fqK9hAR+/uCet3IfVszMn1ULCwvjxqzVS3qPh5d1V2Y1gn
WRDFWmH7h/it/3ijiDWKRBQrlFTvKdn9rdG4RmeTb85tyOWh+7NUNgJe4rn9x/ZY5sToTcvq6Mhi
UuP5m/8NOFT+QDSfWQg3fjai7/DxP5JIWjnFw0VUAjNokODf9YKPSv6YhZZ/VHhsvU/7uxLJgOPs
zEssA8krDNwQMGGr3BBoDwr3aeqpe1/eh1btFX0PpNz4eid/NNGhojazt5wL0fFKcCNwDh+KXfAv
xQsV0NeUiG5Va8IS+i2sG48Dz9L3VJHKaaUPSctqtQru8tv9QGyX6koFj/5nUiNLMgwjKMgZVZMN
ZKPyUM6jJOBOoILDmJEs0E0F4QgXWIdZPh1rERwoQdo22Nj6Luz3ysGzxQFCSNCz4QFtUHTkl3FP
me0fUwWa2zAycm9EgD6ZHEvPS96YhgqwZPyMoTfaa+80iCXWg4dWN4mWf4RDWKKmCZWRj6AlM+Ek
G8hB0v6mfAnap8xk0OjaeBaHo+KqBSpYZj6a5Trn0mLNNF9YeqcLK5w3qJ/YoFbeo+XQhCSd+05S
RFm+//E2Emy+B7YXbtKvgCIqx/4ibbu2FgC6Z9WEfxtVS1RmeiAJff8K4qhENo+egHVWEgUMfCwl
wt538fub3TmVK6xI45q6nd+PD5K43As5ySPt2iEir5uX/RVMTmDAKjZnp9VNw+/cBjn3c2FjX2ry
Zjx+obI1L0jsNh+DrG+jLdVLstERElsjpGSvRTYss/cNPDMFCv6YPx1SeecI+ptQy+ZDly+OMB/1
EYcjppSpYpttePjpSVCnY/Yw3rEwMZScdn2tMo/tJkadkdiwx/aw0ZUtjrfeJ+hx6Z53XW4ft6rB
lsED3hZ2yP/S0LKxH8dM3k/cgltBleUjTAjNjCgIVRW9Bq3zqv6dF8HHP9QWKb2FcVHHVFd3oda6
nv49hAdPa/LR8JBuuI9P/lDuYgIOULz5R9NHz8UJDEqOvN9k6RawG3Dpz0KsjAhrc2eJW2yTae8a
334d22R2+XrVFNKpb5T0XrmJ8aB7aXe/+NhtrWq6eccFI62vBd/ixLRWy5hK39eI998pntbJbMY4
FMZdSewoF+H5peQtuZH2UaC8JHIWYFg+f+4aDXpVBa6IkBzgwzYvrq3u79NZhv1XDOWKrUOU37ki
IIV+bGBpDKWQb6cF6lEMEQP4OdHzy0ltFWG60zGtmo88sFr6b4QoGCFjZ8C/LgavAI2MhZUkXDdJ
f1GzatiuKnKcf+6sAYgJNMyRoV7914I2SQJpyqN72wB/2CPiSvQyEzK3IqD2WYlpLG68/SykmjYZ
Ar39Gegd4nlPPE0GdzT8jza9qzAvKN1psLLq0haiHSVU09gMHmB1jVcthf8EyVG32wm18r18NU+t
2IgZSLhOEls3XPxWHwCMkS8lxUCB5dUSxljNHyc6e8GOg0n8d9iVTUj4YfeVn01vLjhC5sBRzoWE
2mpFTx7NL9IIkGak9It4nOMtkKCQ+up4j45eN0AtVWUCYkD5XkvlBGUkiUv52Hs9A87mKremft/f
bQvpfEAAXx+GwoUkb8VGqxcXxUzWkQwS//TRD+zhYjmh8agxkkd4dVtqO8dGOy6erBWO2fPbD7Bq
IJNdUxM6/uYCFbfIqpwjTZBswrtYkr4ViY3m6HFnOiuUS8jzP2EXAeIsBv0dK0z6muft4rOladEP
0gvNQSZlse6pT/ZFMKT2WeRmLz6WD6RpOIrNJByFxjRxte5mpDd0BIw49yrBOKrTBs1lXc9yG0Gm
lXuFMBlmRHpVAmbp+nLNaN9D0GcOpv37uj3YZOpDwx3UfGVxouw/+nb7P13vewEks1f3vINSFrr9
y3bcES4vrygT8fVvvLP+2godjx567S3FlNIUWrQaQ2GvdWKPiUjKIYALqtHLYGb+z1g7e+OB9/lB
9qq4+vKkSw/j0MfL8N2mAtGxynPtK0eatJov9za+GNG/uSXvsRORstyRzHhPUgGQc87rne6GUhaS
1M6eh1CFXE/pcspSEWoRNNqclYh9XfzIodXfmKRXfEL+vBMtg/3MxqT+bbgbGPQR0dm+jH75PQ9E
JaDtTMd/W6UB/74VODl6UTdUx8XIL0TA9+5PdjW20lAuyRIKROS9mdQpHLCbm6sTEeWOagncok2n
Xh4LDh0s4x2/WjJDgWhpcaEjtpeSPi8Op1sQmkIyzpMd5J9Qx+roXSShPmn5pYdkv59FB3ivHyt5
Us/fd2vSv+JupOZ94U4xYmJoGhhtcqVCdzb7YCdNCJ4itmCrsxXko7oAWSzK38a3n3muau9OuByy
+OKyUGFJTXtPr/csbDPsMnd369hJcMoxIowwFgLm+11NCmVse+vUz5nlDbbZfnbYT39iqwUqeBCm
TR2Bcahott7yZ87F0nKp1hWaS0Qc6VLZpwvVuziFwDIr37UI0Sw4/BNY06NiJYBkR7SL/GEsU62n
2cyxlzJNgVBXxYhbdqtnvepvW4GAPD9aznZG7X5VHK3QW5+EnRS6p924BwbWEE4EaFL63j6sLkzM
bmFGTRZWtKV6HumcZ0MtRJBNQh1pXCU2tPW7v5n92zmpVw+LFPLRwLVYljGXTnqMAMl7LIj/2xGB
gNCRK7kOGWmPzFCcXIYDCDDnBwJakxLrcVOHKOwBQ/03aUIum9wjQHeL4msOVYt0do5LvE/+vCJE
mYlcM87C+UgANwGitNpdbit67fSfUfYTIm/4qKSRbHuFB1lCp4JRJvj6kaHm3uPtSUyUd+KqR3MM
cipiNT9ZtZALNt57H8xEkfU9blODn9wY+KGdm877rXQTmSFBG+KwIt2VmNibJx1Evhw9rrkhEXMQ
6eFmZRpfahzb+KSLD5Ac6BOhSG8TQYN80rsTaSU14/ofSyeYs9uAJ0QJH78lLV1/QS93BA4JEgLN
pGtUKPL2MzZNkznXZVDU6UhMJczydOq/v5rwA2lbrv9E2Fta1akA82Lh8ahgAcNhaiQd3U5gK/39
I7KVjtXtkgCyOld/tOmSCQU5hbQAxyKplfSlp4k9uwIuipeXFysPJOigX3KbTYHoKPXZb+wfV+ZN
V1xFfJXTsbASTcvsN7ZB5JBl9PPlFIUMiFHZ9mBbh2sIouVfBIH3YMGyd1j4kYDu3MX3mFSgYEIO
DESFvkxH0ymVvUOIfotxZ7VIDl4bkl5nkhbCEUZ6lmNtI7hA7TKPeKrXC2xef1xqCse43DZGLhSg
irkua7aJaj28JWdUc399fbmVg5lN8GqgjHLuo/aeI4/ks5KZHghlArclhRaZ7hTDAMCJaqTiTp44
cAhPMoZ8HpFMte8835ClS0HdluiqgoFqSadXYZtG5kcvZ/CVEQR5cKZ0jTxd6KGkDyXC/7Kz/0JF
rIaFUDC6yZXYzWnEeS30ypr98ihmdt8kdStvBnB+rfcqOP857MPYHoaxn/GTw4wbwN/VCvGE8HIl
RCDPJUWPsmJfKUovhjLNjOeh99jJZ1y5DE3/CnW5Q5REWQLQ23xCVgrntc4bvCSKWnv/DyFrtmHl
XTdiiNh+0N2LTooT2H0HCx93PDima+1JdSxJGdT4BvD/Fw38G61+YriRt6kOeHFGhortdjuSG4eu
nFCM34/SqokGvEToEWguEAXuWTjdz5MuFqXLYu5fgRCAi0kM7b9rxWWIGaclXnVlxMy4cuOENb7o
a4ZPqOSDtCD/dtHuXZvBSyNXizmpWWtgITN/EIu5t0/QeKG5zDjRtPaePmIYbKLiCWN7rn6+T73N
Wv1Thkgufl0/TN3l4/4keLj4RwLv7WbtizNzTBuFNUOKFDbHIKq86WMYbtV4N0/Vh8THON1J0mjp
IUVTJbq+oz/ahlc7JyFghTf7H9sZ8vJ5bUmLLhjhIQ8Sil4XNM4cwgwcZig6bF4Y4/w85dUBupkD
TUqhfDxIEzUbBKNtBJXrcJxvfOjxQ5mcvz14tQILrsvHGM2FLowoLhyFxe2kBwqpwyhgsGe3DDLI
opRGeMJc301HAln8vxynMMlEqtqaewLRxyLjigHpM9rBuHPbwpsxz5LhBjZ3wi3RkjdBj5caQTZL
iEgLw+/zddwhk95Jb1ZzFSTvG/igcpQQu8sOaH2/bfAPW/yxlAD2tPPfrAaZ2BypEOuOHtJ7EXpT
r40pJnb1QsDexfYdmRShjXQ/xsWX02MbDqcAh40/1opNrNIPWumEzJkoB1gIiDvwW2KjzsKyr2z8
xbHv2EqPXhr/ow20gVUUTJFxYVAVEpCUszr6H2ISbcKMFlcqzaJU9jeQLnL3YK4nBny9FUowhOff
9CRMwnJ/pixXpaDisiEOyFmry8JeQzdjCyRZXnhFKTKTfyQgnOyDkPOTV6n2F4J9lJBxXDmf2P+/
TCs4B3McQIPujne2GNbxFPav9hnYfROcTFiHNCBKZ40jDVbJR3V7ZFzYdSByqU4FpDiQ9AOlJ6T2
xXZxe9m4Q0MPqDl8s9D36kHi2jhYVFiIHyOYKfkPARQcPPX1fOnCLXhxG5GSK3w4D8mjOUE/Akr9
7hQskz1YaBttkDJnBURkFiQp9kfGcJ2dtDxrymj/87s/oZmyNqkQK23byPDaiHSM5YOBxYfYDm7O
HcZSf6nPY67y41MqqVM5HgJEG0LInYZLdQgdIRAoiDK22jtIZvqUddjZWkR9qlPSqA8+opo7qI90
hyhs+tWntlDpggd+KrJzw6U6xqpTyTjPjnZW/6PHttUYWFf+Ch/Zaa/htZ0nt0iWDL0EcNf1LMon
pw/6WB5S3lx5H9EdtTLWvPdyXlsMv3oah45/Ds3fwygH65A5m2WZdqMdppIfo1U9dcAc0nteOGck
NVK4gbBVUl8xPD+828vAKU3ikm3DRf836fTajyDjCPSgVh8YlZPmN8vsqhBNpYxhyOlWq3vewRyE
iTrOQ3mg2ACIOpnUALuZ4six6tBP3kCl3o7L2biCM1QOxOa3K5IXceGEu5stP1LDMrLmK+sC6ZiR
shqpKsH80vtSIEPwLdZv2bSKmOnowHn4e715D9tOQc0c4Dk2byOoQHojU2i9TS2owdLY6NtgNmME
sYKjD5yglyGnGPSAoR/VRQ+Vwlu/GThzMJ4In34/9xJrUO8XEGbkH9axIf1eOujSIsUXi+k+b2rT
yLlzLe+TsEPUcN75gwPXl1g4LjrIBafZJPxmeVM078WANMzm0fWh2TKzUFx470JEVB3B4eHeWcRP
t79dkCpjEUqxDHwsm/X/qRPC5DLtnqUEPp+5NB1J4+FgZNBxGa4MOtNic0D6dcEE4KaHmmDxb3OM
JH9FlpWQOu1ajkkMDjPR/z65Ffu8kNciAo/ifUqxJgVE4AZCPg5lQqQc2IhmZFxdxccT4QVafKx3
kM/kh+OAaXsDdvxXxgtyZyMcpxzzgIVIarLwi+fDYFdZvS3CcLETxmsLBz6+Gi9vxsexzJWMIsU1
i7Q6HUXLBXobHWfLG6TeEVsTUnO5Min31oDKnshynnciHlki2xkmbVEb0EZxu/ZSreVhPviMXo5p
ewC3bn0oiq/TXC/1u18bBfyQ1aLsztFxemhfEm06ZiBJkJ/zVzzNDmNyQnvwPnxLOVlSAnsRI1x+
KSVmpZcvMq0Hc7Lmz5iYCDGGMWdb1eQY+0eFtc4DM6t+TRzJjZOC4AjgGiGpUTVZzUV3JajM+fy2
HGR5iidSgkt/gaWtyumNML3+L96HDlasIoIBqAf2J6WaPFnHkP6BIu2VRPXIGmWhxjDQHnhRH24b
H1YVcveTrvB7lmE9Q/GBxxN69LimgeRJDrcyJpmP/IjFQ4yvkgqyWiTD30Csr24OjTPBHKqWzfNH
MOb6sZauxrrvgnxNWV8U5hHiSt0bF9TEm7vhhkomX7p0OEQCmHogDLe3Q90/DQeMWNdKhrGXurlR
XLSlnVYk3YBMzV8jWqz5otzZS6iQV0sTV2J+xDwfdouzPdWqwi6YKTlAXmr8ONZX+ms9t/Ukbuo8
lhv1/O9Eo4njLMl4M+ZQSTNroT5ovUVhjPY51jpfhsxQiJbNvqb3nsjHtVt0F57kltiDijD6ctPE
MbSh17jZfzlYfqOrqz2RrXgAUsCyEZE7RHIZWJznhRGyr/dFd2GNhCD48MSIwGLNubGIniTZHk95
Re/hM/nOQwmsGJH/OLzY+68Gu6yit4yEG5u8IivoRNRsjeFm2gzUXQPORjUw8xJP4nAm7xL/VFEv
/nVpwAQdOlXqR3dstojcUpA7FX84Y08um7XQ98tskE1uhr72qE1CtxBHLxLck6u0yObFZbEz68eo
bqC9hmjc7zrnPX4b3pgYUyMGJHyFD43ukMN4/LRVa2OQtXTPMgKcgiXkIxTS7fp5Q9ICqeT3DxUZ
VXOo76xXdk4jxE0au5Pcp1y9g7zk6BP9rlpqOdjTE1G/ny4r28pLNaNihlfHV8OwmH6ESs66Xv2L
fK4bJNu+ea0v3KM+7peaHvkltBXnHhUsmvwnuaQjcsUPeKOLc17cz6Al2bHEwvv1YZUSqS73qZQQ
/PmxUdenmPCvuaPSgzKJZHL9sn8wRMb4ifF3tQLBIqYfkOqJeznymb+4A15fzj5U86v7nZvIg9HK
RUCZpiO5Q2UkzB46bSVNiYvI/gCmlwpcebR7Ck2RApsOveHq0NcxAIfzhN5TbeCqn/AYEi+Wvq/M
04GZVsXWZnZuUNW1igDwP/2a7TGN3Rq2gGrv9OUJVP2qA4anDFaWmWrz0y+cP++ch6wfH22Us9fq
HD6iDFpM/QZo04VoutZZnvPzYFPVQz9/wpC0io4viXmVQuUcfs2eaVzB8ZQwKJNQqwFY93C0a93Z
s1JFW/i74myqI1JbV2dARYKsCBwpovVY2Qs0PL3WYwWGfveO+ROlbtdxEipA8qrNr7anjI70J21Q
OTlWEyu7hKft5nViWtgjiWb1wHK71ZxSNUzuL4Rqfblq5bTQceF3I/g28DzGICMihqkhsmySuMSP
9jC4o6zlo6vOXHcQZ6A4TnDXW6xQ7OJvffA0Nxu0hpmqH5tz8XnVDwTr2694ltEY6nKkl05vNQJP
ysaNdHXeMJsirHWNRa6wXtr/BK9TjxqOp9w1dlSUGQJ6WHCvTEy3QoQ+URQb3Ofx6QImzlTGklVy
yMdXXu6NuGi4puK2lMq5vbAxF430GuvHeb1gLHh9Yg0BZhUPLuLw0pF4D5ZCuXzi/dFbqW0wU1yI
zGJDlGTFfgwg7wzl9RYh7D4W6w1ICJzaceD1ETiNqE0HN6lpFJ6PrIJa7LPPgUDwyHYRV83ftuE/
qM2EZmw7c4qDLngMjmSIHXjWzuAtFlnQvTUMObTHc9K1L/JpjFylRvdOLOuvAT1wtIA/o/W6qz3N
nLl+P6/TkbVurDV09/ZPoKYHm+F8wTp5+32mEcv4a3mriIM8HgN9zaiMc3VOZlakkNkQy/8MoV65
U5/eafHZ6oVBh09aeZz85e2Hh/tl27sdfNVfNSaastzqvYD+0uk8pJd1B8+X54Cl//23nhnCCkih
WezDarx76Vm+uvLBHSqFFYZ+R2KvOITAPKlQRNBA2yF4eqkASdSAoOD9yMNyXv/rzao4j5x7XFTD
YoTK9H0Q0EJzwLpGMNr+EoZ8YG0OThaLf85Ex760EVLNQSU69G2kcotjvScLd8oOq69tkQ76EZtM
t3LbKRtsY7qOSPnP/br5aBIVj9fFRgkwHku0N8g3gjDoT/lxh7uFwsgIuUqCvaV/xbpSy2gcqDVk
38TqyIlghKJf2ODt/3twl3Fxg1X1uXmOi1CLEQxo663rVOrr83PJvm7djZWLTHolWeqHsCOVa9wf
cj+DG5VLBAhYVeuJI7KyDeOww+MqXRfDcsSUDCbc0JG6nkDJWrVA8hhkFnd5UrbFEnNh1ll6McHt
FH2HuaxkZnrq1QKis1dhl0tb9u5d7ghbwmspIwLUpstJjmU5zAMKOQfIBI82hPs01nwWpdoaZ1jT
4zFCU6MQAFGS5d2RU/SLpO361mEKKycnDWTDOwWERS9hQTNu0zFBS9GpJ0R/h7DgmpbC+kGuz1VH
0NnGa/yCqoSurIQkHiUZZOIv0cK6axXC2G198PGtka+8G+5s29Q5y2lpDJ+abpPVHSBWXwmzVCf7
6Ev4lwyoOGP9xYyAPgNivfxXMhzAj3gLVudpBEA5IsVIcIWGkYvKHQ81CobAb2VUMG13UV3p8rrZ
zfU6kdv4QG1Pn4lCyKxbIyu3UtZISMFrxUO1cOjYcbaEfyZfqH1TUuDxHHxqo43FT4Z9hIMQa67M
581gFNCMjjHhcoJkpFEmJMaawE1PTe63+pxt4P4DroML6No2WNZJJIoHTM8+y3nt/bEq2pwGrOZE
7oBaq9fud0AIR0L6UhG7QH2L7W8a+1jl2o7+pkhtcFu4DiY7dGo9DUsCskjZdqQgHFRNvI8sTuFA
muj33LYfgRXhrUFO0yrMKz1u66bOtKMlmVumukLZIaqUqQp+vwooGLAc1xmgrZMuHXVeeLXSm879
IbsM5eNQkb4dm7kdsvCyzQxnT0dabA81P1IXQr4lGEIcp4yA5NH0O7u45pTzlig8hl9tM6uOSMQh
6gbsC/LbSrhQGjfOwf+NkdEVhMIAJOBWWtsBteMeRZXqRNa2oNJtx1PMLMw/quWyJXcdKV5XqU3e
/2vCd3p2cZdtsnUOPIt+n70Shc8tFPeU1mpuML1aWHVsy334gIkBGnlTgfxfZ88K8tWKtX5FY2KA
X9HVl2yt7HI1qNbCQNnt6dtoheVNT4XbpGLgdi/kNMWbwvBNJfpnx9zvx9QJIwDuHXgC0B7XgLMn
MSDHhmMJjRZtJL5MhKVeBhqjJ3BpSIKXcPBmHInnYmQ5ow/h+3akG06JwaIg3PoCg755yHfMvvKd
WlQoFJ7sG1mLTvKClcj4kx7VOXTC/CoDPNjiIgit8zN8grHq6Xp1pzYyTBsMPWsPXHP5CVntkQ2L
/LxcedlpAwFqdJXzMmVwiw/9j5owhEKoTFUEhOTbxhKx1o5AKF9LksudPWHpkRYjlCdCb3l/i/vl
1Sdzz8AE0ayxJLXJ5JYP5SAoHECmdmkmU/CdS2+/hnSzW+5Q/xvgNaKI9Zx4fjP8RULY24LPjrp7
y4Eaj1kMv3xcMbDgCdN95OfTlBEFMTrbs7caQ1FWTYw6aMr81fmSnR95rf6LFSsAEQdygdA05gap
9BpGB+IZboFm4gaUXM6iPp6EtXsitYIDo0sX1XbuhrKhUGESqL1PncPvdVSjJMjF39Estz+nIklx
93N3xGsURiL8LL/02tLsSLgiO7Lh9L/Aw3o38FqNj7urFuvs1HwkIUSyrOK2iH/htDTUqLPTuAEP
uDXFj6AtIZsXG+nIKckKfT0DIUF9ZImv1MUv/fjLYyud8nE0ebetTiEGtQY0g9cgk57wls90q33d
0qsLsKoL0iVlSdFDTNrjmc6GDDe7qI60bGgyaaB8kj4uwlnI9N+0SMvwX7Rdbj+mCPzhMjiZ8shV
GIYKT71BZnqjj7+R4yRGIcix/xG0w9p/nleQ9tkEsOg4cGQcIkoG4Qsii4eIZVIze5iMLHQQa5lk
UhFGCRuS6XRmn9VtMP7d+Y+HhAvqXc4kiWW1BF+86iovK2VKD4TmuyZ4+ghAqDpfyJAxRirP/FtJ
vkpSZHV76omCNIBlb5+MQeHrV1jR+VRGK06p8nhBQokqmn7uv6q1rIjZKaeLMqJz+CTDEzCvqrVB
R6ZjCucCIQUxZy7rRX9/xqFCZEsn9iFAJrFykIZFczXJ//abN/rAyStt2WSEFlHctD2fPNRofQYI
SIHscOII+e7207w/rn0auLf9PzFznJixeU5WAdn5w3VTVWPA+XyKovXzGc/usA2UUVcg+vEyedEQ
II44DwIthE91biwkps4bIIuj4SMeHPtJIk/X6lNf0reKI73zFCDQfktEPq/38fFXG4ueL2wx5bEP
Ah6KfgI/PtZkTHTx5XpAeDeO3KQsXRTr89zFTJhopg4a+f8dZzNgGrVHeuFNmkFzcoiUSP/Q7+pZ
YJRBndlMZR0C4yP8vbgupONqK5mpes2aY0V0bUMWYj3j7k1OGhUr4dthJTYXV3+6oBVEDFOG2ak/
dv8jcMu8jS1tjgzj8mZJCYLmviMJujqHP4QrYHP2SaEevC0Ug8QWe+lmT73ADUT72ZKoiiDdDmL5
dMBFSkFEqsPWrFkwIj0qiclyjn+P/Gkk3+gK1EugdV8NRw8bwXrk0Wu1LWf5f1Wt6rGG9QvKxz27
L1XnL4j8UJOh6TKXdimI72xUF120dmlu0m1hNtEd2LHOy9EWkdR5twfEY09bqkZrkojuKKduHt6i
iQy26aGNKex95+LSgcFeCoF3mNydi9XiIewAx+QlXUbdhrpVWYA0nncEOA3YJOs0aDwPEFzKkW0X
2MCyDH5A5y/FdXvSDfILkZtakh1Lk2CG/M55uGYO9KWtos7JXlRtYJGs/pC4jxozuLYG+MivjUCd
GM3aU7JHH8augtNrYVJvJhDjakochByP7mTQ7297NO4nsOgWIxCRQ455kBQNugJf2WKge/FFzvyR
CtZ3Wggev4F2tY+TZGb8cCYLhrW/3XbTz+xV7cIlqwWmDtvo2wp0mHC9d4xo4bHSTgknD3ef0JJ6
/oRHU1yRVVabjfaNPJYuJUNIrOzT07nCCzpz6goOZwKmgEpR1/0uTvA28hKS2w+oq8oWCOY/faFn
DWVh3mshrM4FAdtPCFkW0wQ9I0y1xg1GLGhjZ91AY9rNFIl3E7RkGBK1S8dcEa9zs+Xih7m0Q7qS
8WlZDkuPlxZ8yoISEWwDP1MgyJwcBZa7V49zEh1pE42WfpMay9ykbyFL7ZCRzGVOn+pyMboN7wqK
oZWuILQU/kdo7IXfTej3q1TXpNV9AB2K17CcRlyveJyFijhyst42+n8WvZoK3roge2YkSgrn0rkk
eejcOxTu5e+QL9u0F/+vl8hd4TOOF1OotJAc0PmV3Z6OfmpIysUzketUPslSafcuW5LE+rH/7EA+
dPpM1EB70exA42/Iew6c7f1ymrixXffegXo6HB9gpOWd6K0DO6Acw0lQUpAXmwi4tB7IMLpnvMv7
3x8iSmh5ztZWh+iThpkvPgkExkrIV3czJ8EQkYQ1xyf8kTrk2jYMhpzZLZFXS4WH0zZmAMcsBrgz
vm2yQ0rTZhpjq4D2ajD8LWNx3mdZbydCBtfVmt0OthPJPe6JhvFQoTdaiiEKRZW3+6jkTRt35j4I
nvl5tYXqxCW6wAHmjIU0OVbjzUf9L0MDb/W7/1UFRACtuXqG0CucR3+xRvD3klVVvh8f5FN55OHl
bTmaIpUNfeWPBLwWhAhXX8K+zxxRUUJz0k2g4R5OcWPltZ972PYyNw3EUC+eeFG6See69EXplxB9
eePSLUyoqkkwwdg/07+ol9Yhs3LOe48iPTWD215vnIe3hmiPlIa0Gpd6UqWUuaenAa8DraCEVUER
F7+VuhDOGw/MVcgOiSujr2JuQ4GByguSWQmP/21wfx6fel4dY7bJlq7rellTeKSJrrcFY/USF3g7
umFIIuPq36H+i0CGWi5L+bZRd1NCavpPIOTvuQmCvrYi/i+5E4+r5oPFwIZFD1R+aZ01LSxv9BJ+
i7GffjCPrgB8dnfdhvHaALczhRMtoq8/+MzuDFMXBF4Zf6kxKMOyQRLB0rSyWwQMtD40jJtATBWt
PdU5F9fQqpdeZu/v3ZNAMr5XzwNPNeJSSY7srfvJyDvk3xoRFoR+qWi5TD3umoWJfl7MGUWnZTCQ
Q+4AK257pmdMQgmfV/GxwVTZVISjNBtSAbu9IK6uZh/V/MVImr/4k8wLz1rWsvQJQVAkfpAGZ8bh
Lji2JLyuRyymxaKLLbe+zdcQm8dpJbt6FTOY9NKE9a3T91h0iRHraozdA6AA3H0f4uVcBGYL3fPW
ctvpvFgTRrTatc6RnaxT+OqCTO2NQqzFOAgWcmyhdRKjjTBlucyHvxfRUUBJ4mYcX9BGGwLlLH+g
Wvvq//+VdmZN5k40vxVTes9vTOJWCjkawQDDkzoSN7LYFZ22UAhsoSrGhsvctHcL5bgAWFrv1OOl
beYaQBtKOv33dkzezYbIee1iF8gAhPMkbiilyWWj+/rKUsG9iCnVnUCnLCZB52acmas3/N6xDbuJ
M4wbREsnvQR7aNHQNmwTaCeb0IugR+CHYGzv6wCq8iRTItcHb8RVvCNv5NWOGypaGX5TUH6xr6Uz
GSXzJPzP189bbHny6wW9yz5aMi4DpOJG1z7/7ITXchFFR57nlLxf7EUQ87eMpB/FcL2EdwbXRowO
KbgnFtJHNfMT1nmBJFdsehLuu266LyyLas5UIaGz97BylCllDvKC53gEVZGmAncmhz6TeEnvXDYG
6BGQJ7+1JhF54Fhlg4mbfXW3Xaf3UlEcZ9xlaud7guoZn630JgIEIFzQAYvkTvLCpKD7e6uOmbiq
GjhuhbzpRATJYk6EwKUl/1+MBlXKpiX3jUEg+pbHHYKVBzen0ihqNudsxyQltUjFb5BYKh2+Low4
Pnbkn97QSV+CK+V2ZZkFGWypGE2OonMXiQs+EId1OwgS35/JqPkmCA8lgjM50vwMlH/721am1PwQ
1JQnDEP2ExbQdN7XbatoFV2SBbEUb2DlCVV90Yn/AsxKJrYqqN6V4LPAYw/VC3e2Yxm1s4Zhn7zl
CYSbcHlHbjRsVn9zefAEMEZWy9ZBD+LBArpFNVf28eelc0J5KLjFZq7/4WB8Aur6xq40zeBrrDoR
BjhNhUEMLhCgMTtmVhh+rBL63BCoNsii3ogaYu0CIXhYRdbP6/Fk7gL5xJi/qma/DfTHc1HbULaG
ggr1sDaomVZsJNbHuprgHWV44qmhHROGIk5xDmuEu8dBOi4IEkdBY1Hk6jAhxbiOBcIZE2jFyTzT
B5jxvOF1r+xFukiCun+yu3qmwt5LJMMYpiwa+Y0nLj59zTV3oueAfOvBopeQJjUcHr7Nt5HPCZpp
RgKEpFjyzI3e+QqXjhWg/i83buc5Tt/FqdPrIXIWrUMFU/jXuk4SZNv65d1zWrRa51OqIRwZE/cc
CZMkDQhAHkde7+gDkC2ho1OJR9YWcHR9+AxzUqCC7teZokurjmug4pSiUZfXXypPcrfQTM5o1TmN
xFqUbDPiF6kckwvQseayuSAi/kqvZ6DQpKDA4W11hwDSEg+WtmBDsk9tBLZePovFKHZjnFqyOVj5
1vTR4lQB67vYqAvGQy1H0JKSv8wI0onRv7xdtnuckWAAelo9+FP9WWy7zr5nThMh9i+Na0D8xpNp
tTb4U/Bt9JyiDv+rwXAOWBLJ4uPPTubdQX0Miy9I3HPFwo7RRr6t+/Mk+oYat8bXxfwmzDbL+INh
oJwwCoSVykKS71QNNjtNZJHYnDSV3Ja+Bi9XrwjFeVDoEGTamnXBiyBrKpjiNZePMxD9HC7y1JUe
ByuonGcUoDcrGQ7EWUjlspkmvnnKRF4wjqQ26UHPD4vihiuX0ZpkL8hWsiLuXlMNqSQiZbFzSiI5
Q1RO9o/47/r+1rQhY0kPA3kbPVNbxfjLaDfTH0cbJntDKQWLxVUdAzHnjCR7pTseDf2wE6MarrdV
qDon59NX9xk+XH5Mu1ffrYHCSMb5LxM73Qw13uNZ8ras/h+/RXpel3k4m3cVuTI/LP4Y4L6dOG7s
xHadkv3vadTNXhwsUjgeX5UPFj6YXj6WO6xFayChSn7Yhm8t1VRe757kIkWqbJyazTSbZBNZ9rXw
j0Ot+OC1KftxepPgNf8QiJVJNEViA2l5zCWqbsmPI9N16TDTl01+ThvpbAJ9Bce5Wi3g4NXO5oxW
G/U5OYePZtxE8+stlvUW73UrjwERhh8chhXxICcUZZTZnBdRynlWlBpQHhzwcuLmnDixvcJ4y91Z
GAx+FdKy1HJXgqwuPiJinr1k1tVGgaX3TBB5CW82lHqWS3pt5o3TYkzXLASHsessHk1jfryWv2Sg
3QRM4gUYWGKY2S2ikDY0KY2xf4uOovu03rxanW995NyBZzL8XbMyIefzrQ1oXkJVGrhiLPnJrPG7
YmvKC3YeLdcUa6DFEEWrR8/NDDQ0MykQfxA+wf6UoTOF6dVeC43v1kNob2JBySFv/ftX+pGQc+WW
Hcp0aQs765t6tfFEJAsmt7G4AFy0jj7AbnvtmEhLmqCM74eH0wB0UuYi2G8ktYBasXPq9CbYLPkw
G4Q57csdx9+cUde8FM6O95Cm3VPFbWliknxrhG/3/aImawak3nhWRj6zbWg5/kNTjknVwVfndBlT
MaZxDjYBfGeGg2UiXptU3m/q3+KcBZzT0rWEdy/C2YqKTJlwezZFHWu5lXie01Os5ZZrOE/zrFnS
ACxsWgpPNHHJ04pPIuAFIkUysmYuq3QLdkmmJeW+rRnTWjAjMgcIIx9BPj+CNjSrkVgi0nCry6bb
rWCFq1NOUjkHlMCrdtoxcBWBcJ5PqtZgr/AOHLmWkqzGDhv8m0DGGZyQQwhuyQFCW0q8ETSaA4PJ
3ajrDxonG8h3n6eoDZD1LYfwRRk73yJ+t0Vr0m7LEumB74tY6u5Aplgb5yKM3XZu4JHxEFKuz2ja
A3Mt3Nx6DPZYpsNb45lLpmt66wDxR5yzJ+YmKjB8GrIXZvgtxJtZMUju2UeULk8i8QkoQS2bcvPO
NZ16RIwHwmng3onDmifKg9pw9EBmUjGakm5/Is/vlYJQfk/ax/GzYvbj9/y4COLflxQjlCq/mK6g
KRJUT4dMa0W93MvpHotSeT47yJbFBDP3lZdaytktidthfKCbbyvVB0v5IZ1KJIoXzpUWsjOSRqa9
vcuUR2HRsl5NVN1CmPMV6ESSsZR2dxjlF8DKP14iVDdyewF2aDZekfsx+6Qp59cDED06sD2Wjs+0
PMWdO8dVlIt5UUjejsQyE7gkArmf2AKy1RBEHGTMxIrEqrtZ/4OcIiHo44iTIP4Rxv9zrxwq2kf7
RweHVm7HYxWJiBMBfimstL3D722lPxxjsE1HRtrma1m2DJGenZO9Q3/dalLuCURCmHzhB3dQvWJX
qB0uYlhbLe3hiEnlQtNPMMov0X8lHLHZ1L2DtEpx7EpcumQAO1g+iwQEyU73TgDrt4aA3H0yy5wC
FDswCmhk7xdntydPIdFvPrLC8VF3Pvfd+2wbtRd0/qBluumnRxj5UwUbnO3TIZxEUP2AZcUMln9m
JOdQgQGQHWoS+aI4Nysdmxy7B1Nkn/764OCb2lEsGOOodwd+j9P9AVmye3QM52GPCMAswZNHjuJJ
IxPmdoGuKaAt0wuO2BmIC3n/KQUOvWQ8ieBF31lyyP0ywNY+Z6UeHNd74D55PR9igKxmLHESMJtj
dnu4P7Msw1hSMRtDObgv5R5dFrAXfTPle06TFyBqvnfUaK+cM5oik03gKFuYR0rwtSy9JIgTjhES
xjTqryoptjgKq8QnjjbzsVrvnSHAFPg46IFbn3bF9NPp79w1fIxrT5Jrc7z2SyDTSFgvoFeuf8mb
GHbUMwa0Cb46CpJw5qZyC3FDTXTW13utAyLOv1VSicPU7vQ4esmUXEmlM/IWQF6rIrijkOBOdAct
c7V5YzcxHACaRxp4xefQ8MyDxXQ51q7jW/8MCLTctkrbLgT6CBv5ZFTMZ80Q1UTLUQobL1nlDTnD
h2VrphCQWlql9clYoJqEeF3cvRkEUSFN/BJAfrpmRoRx6rJNAii/CegZrhzyHf+j1GYA958bACx+
iroHnt3eU6ZpMULkzNxecv2yo0B/ctJLijzdUQxs1PWfmaq0G0CUJhdfyekI9DQvVcSTAbIw/1OJ
ExqIySAbpVE+bF37Jh6B8T/7JYfo8fDl5w3ogu52IXbdySG2yrnRXjqIKUmmOo5wTE/cinkQ0yrm
RMwo3msT1Fbmhu551iHnmBgstLHXBe8QhAOOmZQ9caRRUYEAGkBZejwr3n5em/MyuaPf/TEqbOMd
DvOmmMCNhJeX2P+QG+cMel3zYRWwWEp7ID5OvvFStbiCOvqBQ75Rh7tufEvlCcM83PSzf4T7u/6W
kMdL2l0oQr3sW947WuWHNTAjE7Gfp9npGJNdtpFK0hcvURv6ZyTKgsquteLZjmsJl5ELVFrdK2kC
18s9/IF60Br53sNYfLIFgO9mWJUY0FgCSx3xIdd70y9x0ObzUOob/Ys2zI2Z0vFEpkzaiVgoDFLn
vrBOUcm+vWMRNgJe6aBW27umRuKpjOGmLtktCbf5x9JCOUhpUSizk7nW9QpSaJ84fY8bJZ5iMhkE
LSCho1lhK8vbtfa6umFx3BZKM1sOhYYiWcKtv6PR4jmlHCo5o1Uio8sn1eE0kD9LzXKjo+4XtsNQ
8g+mFTfBGdlaVrHkIkj06hMgAm/JRBrL7fdb/qPnJSYGGSUvkuBPemWF5t8rNIsbHz2V/oXXWsLn
+Cn9JqKYlzv8cL/DV6h0do3LCk7OVEPsY0h6GGCyOsLZkzCNH2D+r61CX18y9FkGUvstj5aHMirs
vmwGHSXx0GSSGjZEN4m9yiw5TBBlMJ7ARTkd9Xt09c9lfwC6qVkM8Go4h2/ooSs4Y+TUmc42aiH/
J8Eo12znTQen9peOz6cdl22/CY95lZGj0am07xKgkV10Uuq832enK7cgzJuaWKPeXg61OYqZ4AX5
yoeXqKn6SBldsHLRk/D3G7ibv4LFZP9BBOErOe1w12+cgqiqO7Z8DG9NWyA25dyR8YiEYNeebfcP
zkSZqMrEUFFLhE85dQ968yAthyj3Y2+42mMQihIk+2aqmBubaxQpP5xyi32K2E3b9MGWszX1rGcz
+iCxUF+O71x3jYXey99Q69o7uq6Ey6xzm4GqOonSST0bDoG1yx8wsY1t6tHR6VgOazWsNGJw18m+
KarY5ljb6s4roHUhfOpFgAiVOa5skxGWc723xPUzC9kErzGBHKE7ECQRAYcYFu6eTpJVQydLF0ie
RmXCbOrtaXXFSWRdNDdmWRQXlxo4teyfAk+y5Yh8iT0aQwk7t00fHOVVy3F+FoHGyz1eGH9G+BAo
/GY6ycNsPWDPUphl1j/uoYOM++0QyY/zIbWXiUq2cYaM35no/0jEyoT7P0+QsUiYt/sFoUb0Vb34
HLKdLvu3qoqNvrCBM7vSoCTMWsSYOYaG4aibZMxEqUsY2qRzsVPwlelM/BtgS6ZVkoXppy6J8lYa
8/aFmIgILDraPPX6gpajQ3mb/Hicaxa+wXIEgno3ZP9dnCAX/BcSfX1WQRbzN5EcbY6NxGepQWY2
jHeKz4QR2VBqRD29vjJPd5ajlTk9CW8E1RWfC12TOlkIc1THkHzNxkDjNkQap//L/T/6v+i2nG5Y
Fco7vgf4Ik4UIVlig4l3yuvUz2/HyXkAele1Uc/ah+Ax2hVrkBMsgRiKLez+drhRtDBN4GNJOJ1q
WB6S55Jm3zJ/4c05IjmH9h+ZSa9UATe0aUpE1u1u8aw5lldW655bAXyqWOmgxDQJuVO73MF0Gpmc
vtbb19io8+JbPyhYCgyway3acKvnbmn1PVUbeul8Xo/lMHVn1zJk3cP4ugN1G37T/CdMj1Jn4//w
6UCcSsyb/OKF/UioSGMhQUWiSzzH3cTJLFJR6CRJDEQC6nmVgIPttkrOw6DAf7kmhLvE7G+34jrf
ujdIgjmyVZTuQX9gltIRsFGrhy3PB61cPDunbfpM4cmuJEiomwv//pxqhPCDPaJptwP7UqEc6XeM
UaGIkhxBrSqyMt2kKmO2uzvK5BYvfRUDoqCpyFjka+NpjtO1Ya0nQqa9w66f7EwuFC12jLaBwVl9
B8BGEcevt2tDw4tVvUUyHnnB4POIl9aXvNmqfuwlZOtdajlEjyTZA/iYH/KSj+cvB0VxO/1DnyXA
PlVnB2xDf/6wmoU/RGKV/AwXGnM2fWNEVWvrZEcj5WCT8DUfSF8H4Yh7LDairv9xRRZAYGQSEo1w
0I2+U7KCqgU2a4NScXwxKp4dcxtOcXpGKD9cTP1YjRL6qaIl/ueYRO1nWqQ/eyg17CB9K1E3H3RJ
aACHWcoImiPkvqVs/2GzfR7wzzl10YKX2I5HbHfoxD7EFvdqsRNRPTUoWiPK+lC/AKwQT6H8LYjn
PjVmnLMJJ77ukwew3+4goNjQLMbRn6JnOfLRPxD7IBfnejVGc4VjhYMWXFExgS+xzgxnaXMNv6ct
6TtQrJysWHqRE8Pj9jKXbzEXUfLn/rmAnnUt54hnVdop9ZStzt7tYG+WDpN2RoVz1YsA+pUQdNaz
LeYJCDkbvvGnNwpNynnYYkVzZ8/2DYm7M1cA4WaVcMW5yyzAolvqZtG97voizZpW5MZC7uLhGeAH
D5CV3JCdEIOoZ3hUyD/UuHFQSxwv2liB+mZZZrCnR38oZ6j7h4kacEIPAPVRmNTcfAascq1eSHR4
AtY1YkVmL+HYRRUZyey+99qNXosMxTY1ik9rnt4j4opLT4CxdsGS9GY30yyYgZL0wudfSdy/iw+j
ii2ulopr/UeARRYhQ/5FN9JfT1j8nrrcAUjPie5h0UaWGJZtylePBbPUA6FLG07whV9rNZk6uA4j
b2wg0Z/QSL2NZFaPvt2QziwYc+UOp6fVC0bDuBL1BShQpWzoznq+VAUkQRjOfs26dQ5NQSg4j59y
vmaUOruIDjiVwLNdw0F43OSIk5txOxh3Vdo6QDvCxt2+rTVPHkZ3zbqdzvSVImM0TLXZzRtsKzHi
KD57Vgg4ipd6W/ClJAyA3/OsSEb2O5ZYi6EolIezHvJY8i+D76dyMZ2kaP+78voZ21Iep+LPlzTN
SpKuSZM/Ykv8eq2a/gvr+HojFqAo5bHaU6PpGIe2Spf9eFFlKijCI8KdyhUUijmpW+bJ1ffdt5jt
Pjq1m1cIOXDeRV8OT3PfDMHKSMd3ZNOCp60ObBTR5EG4QzfWG69NfPv9QHcFMqcK9NRqhobae0AX
x+EubyPLirjAiu+nnf6gkiQQmDgjaE4gQt+1YSYKqGStplFowX83I2DMt9V/Ki6R45kPwoRzFevI
fXP8gcDBJc2qPjkm3qVvGgp55m/w9Uc7BRiDoSFz/3zF8gbK6orKIJpXGU1jHCiVjR3q+rbLorMl
Q3l3htx1SAZRMXxv5oLwbA6L6MN09fOpRNTOvcfXU9lZVZsOOndPNPL4WHXoh1Z1qaGjIKQp898e
IppxAXE0N/0Bu+DmuBao9lVqDVXwbrYKm3xAH3n6jWnmlQWfm9JaC6ynl8cQjk0kQqr6dg+BMe+V
LMoIOjRGAAjFJy2sEnnFleljw3ZKFqlNk/A90DzIgtJgXJF6ePjUyQpEaM3nPMzLbjcrdHYI/kyC
RGnVvJhdfyBvWibnDMcSo/49Q7ODWba+aUIl7qFNYNqFJiG0WFLmvPG5fPK/x2KZYuS2lDExH6ZN
1/KnJWf+GCDYGlk7VCl7ZEQ5fHhhQjkRSkwDqod+NhL+FMN9OhguNf/gwHC46MTZMIUETATPaE3v
9loh51RmHmzdjJkB6FmoDMvYBkAA3KQDwygdf91Q08PbYC+4U0LzuRxObpUPc1IjiaZGr+wjBxAr
8wwiKydNagrIxg9Q71x8PHkDz2hj+KecCZinOi+t0OukxaIfyT08d+8vW8Zi9BZg+APwJyAuVRDv
3v0T8ehB7MPKzZtdRxt62FGWXYjMdeRox79vvX/969ZtmUZdlaW1fZNbKygwQegZVknuAvs8yaHL
QIvlszEW/5J/ZOZUWqiCA/0x9Lzddn/Bo2K3I2EF3ni3v6V0g/ooMNy9QXXglrgkOciZ8j7HYK7c
HiFkDh3A2WSzbl8GZoln8f6AtZFh+07eW+4VdnbRICBa0N4wiQRv1Q8hWox8q/C9OpDnH78gySq1
TTOhDQGSTcIdZ/5YD95zK1uxLWI+czCeZb1S973qu4P9GiQ+8j8Xs9rESej+PZrMYQD9f/9bKcnz
X7FYln+XuPiwmcfhLeeUuxDxz8W3rg1oMuzFUkh2S4uuF2w5yqHnhM1qt4xZ9N7bwYFbsbX/B96M
D8VYj17xJl3D/qjD/A3Jq7PsPhj5nzq2Ph8T+XvUx5IUquN63eztEEfu4zgWBQsT7EYLFbqOnCtj
fK5FnSfQv6nBqBEfgSyUpPd3i0mDj0BTkRACaKOfVTjyv/tHcng01je3ea1IYeJPBxKyVGLaEDIO
58qUWop5s3bx8RZlrF7x4xd8ElMfy3I2UUP++Yv7Qax9da3T7ZPpJ5ClPEaAVREVyS1+aO/cbiCR
vaIffPci+JC05fWPTGjRCJoSKFKnGb3GTBbV1wts22NTvwbP0dLFcq5pFQTLNnivhKMUCktxWmkX
ZP9PYf9+HxIqXBZ+aAQ7gqkX54JCGAO2eBTp/+ZPpdDsBFWTI1RmCUVbwg8sATfdiCcoisrJxO+0
Nh03ANA8+JF+cXPzJ2/qXtDPhTn1bH7SPEBeDbtDeQDI/Y8pup5G8IDAEcfIgcm5OX2i7e9kMSWS
/YOJVy+JMCQVILFXi1kzmTmaof2qO21WP1WJJ01nKfgXV7chYMGc4M3fRdgF9vgn3sbJ/ZsOZAPX
/ePZfFHLWgwK6dOgy1zbSC4p62Qo8oHm3E16fv0zEwFVsJ6YZCdrM4GMRBpxEk11izPA2xgyUQWe
tQiC5w22jUKK3bK07Bz7sR5IMi3TwtUPzYYS1tdznuArhfu3DVPkatRJ42wo3ejaGfg0WCZHtI20
keOme3HNsLrOsWvIrlJJ1E6zUNFyOb/Qk3F9a7tEVPqmdQZRjlPBGSTgUE2FxTazPFhAiujG6eVO
d2Zy087TyudUeYUzKmmcDBUCUgxT6PM+UfquTpt6Zeobwlgt0WDcxH2JLlhq31rp1sdsyOzh4Iqs
8JGHuCmqzv+t/e+yk8O5RtcARh4pmAUNFeosWMpwjNx3Acc2Vqn36gTm23YOorTy8jU1KD2iQBsC
vxaSuzC0T0wTQIE9uGA74qenoJmOqK2w3rqGPWB8It4JrPlvrQgTGTRyHYtuFWFCfxUw1ch5iich
As34byNLRD5pJxf5XjLRcjPpiFBPyNL3wW1oGM8zok8DP6WrjIIgZKCJbPaf3Ps0LhP57o5mvbVJ
Yq+MCep2Xi/3BYbrY+R/yvnqxYuWg0IHJqIFXyW/LHUKc8rmmqNhVP5TghcyxrjLcIFSZxWiT2Vq
nBY3qO7H3+w/nLpieKU39yJsQgn/2aLXuezV/WbLdS3+9rJI0z/eyTCe8N0JRus7bEXR2FbBr1bz
XQc0Oe6WgOook3mJFEVtdy18F/iHiF9cY4f4vFFUoIuYcr07VbOyuRX3SiwerBKxd7F0tGqLxnrU
pJ/VqRC1g2BIT+eSQkt+fv0tMyhr76vbyUVaNlOIL+xDIjyqVNJkkXy0QwotQ9lKzOFIS1VWhtZz
JBK403wtI2iZj96TSUK9GZYtRrsoP2s8Fgiv8smSiUuMhIuu5iZ4p5Dx5sKoKeSxAMoqVCY1qb8/
QWsAbjRaAUoF51pTAna1dJgXaxYz56DZ0btCGIbWq6tsv9OiuirAke4RiWNEAYeV9Sh34/XGH2Eu
zLmkXtmiDvn4ld3V3jNlQak0c5dxXzZOEO29ZP8Yp4YFzFUIq4ix/KVtDJ3eCvbMJYWPa9JWvJ/h
s8Z7o8wFv+utoAMpt9qw/Bi1worgCEHYihqcOQGtfDjmsDwiPzrjQNciludQMoJPZH7D0YkJ/akb
jGJkFHH6Xd9spGZ590NcgCZ3jeEP8Cr9zKXC8802Oc8KgOhd7r9rgrgNs/9LoqdvLl64icOg5Cmd
LIHkGlAYVC9SAaqzw7W9vX2gUODtO74p6TL+GIcPijqCzE/lrtNfzKOT1gASB9LyX5VLpNzAJLB6
vewc7txuCU9MkQS56fTquLenfsiN9GUpCK2UciDdGszrQANmmJDdDLF92cxTW93x/xh6P8OOa4f/
BD919b5rGJq1VH6HVLuq99MZMWo3GNjbioYmBWsBbSE+qU4+HwAvWmG4/yEdMfbKf5Sw7LE72Ja8
2NS5SduifFVB+fuS9HXvkrVkH/2mmNe7Ji3DerN7gVycbbCwSgWl6xLPkSuwqZOHZY0pu+eEhJ+b
1Hk3tW6o4m4E0ZoiqnM1BalstW2trNlZpR1N2AozTM+3YtPciImTBMw+EQ7HANSqF7a+Jug2QQrt
4kd3JCV0kWa/lNfvFMHmukN6nnYoFb8ucV3uQ2++bpOvyLakF5qwuVWFfSJTXTJDobcL/HqfBBWA
jsZtekLG3rPPGDeAXSPnLIs4hlOeJC5YFOz7lu3jGcSI1UvVGejIAegPE8OjzOYXRG1U9e2lmxIh
bEasBXgL3LoQ3W7HJNkjV4R9QS5L6/v7eYmjHxjYb1zYmlAmx62IIyjYp+nMcFbgbxPsxX1HfneU
6lpwRM/3eKOpX941aOboy6z2zn9v+Xgwgsi8x5/T9JNxqMRUo3XfzL+i/ll6Uv9u2zC5AVlynaLP
BhOl6I7JOITFj3BWrwohGuoGJyfClu7FdFdbXg5JypM2P/uY+XyeyEC9MkH5GsJ6RJ/wofoifmly
WqXwo6Sd+NKEUa+e9squ9+Xg4o2slYVzQR3pm6lphFrg4vVt7mWI+ytUQm72tHgeLLBt1hG7qbJG
LvQ4b1vZJhjFCO1wjg3QCwIF4DN5gANyxoZkx4ZQ0OlasyJFcEQp00v8Fk+VfUtWTLwoJgNEeEze
uvcenzJwU/n2Fh2QH3/2ijj2i1ntW5wt/RqdwMlx3KnyBVsGgjAf/XMhxyMEKwmXLTmNC+fxMKCl
a6CCF6ab1md+uMJEa/roM1XeZcPFTm0oGo/NQAuAo1h8Z2J6ht81ITk9hkphwwbdzogAxVo88SQI
/M4kquNPAX0sm/nEjMuU8gq1fYfMaEKmAlWc8BKz5zJ2MrMVnQ+g8Ixg2nWVuvcSH2P3blrZkxVs
VL1uHAjJJ6GW6MqEfrQI0QhqCoyWB4qoxiKxVU1BHk4Fm7coeQRY/x6aEr0OJrJYglZoeEs9lWeJ
R1t9KColYK+60J7zwJyGuLJw28lKqHf7/BomgLf2uTOoCRecg5AICaU70Wv99cMEMwRN8N+AFzJS
n5nEMro9fLNTeTr0GRlEvGOkfL8/PMKvJRlCjnzSzr/ZinuY0JNq/e8IRS3bsHkWubpz1Kx5VT90
Zt+quq0nFQOzBCcplk7CIFNg7zZnWEtS1AuIz+SxFi4dn0Ibq0B/aTZ8P7KBAAMOC86amU8eOtnr
vphwiMhCfn+i8b15S4hz7UzDuAXnHUJERqgRIzI43T/nIc2WsWBTTNCXRkL+az7EgQBi09TCLRkK
4eB+J59Rmh2FulrAbbCvf3tsiPaq3YjBftLLytFytoSxDRwmOCRigkZ4yqSpbee3iYYA15wm2T7t
878i9GMBRWoLVP0l/JPKmK16tppvrCj5B/RlzokBBKhrGY3B1UVUDftSIV1/RCUD11j4ve5svZ/z
LshcdtGm2u1DUVoZhE8mGuD4qiliKIvoCSzGnuG6D84XpZtvChjZ5Tn9t6lePJtdWsKN3YbH9e3t
zzMM0Ch+HG19mbw86BT7yIaYgfmEDZw6h8oXbLzSpq0lNJhBOIPgL/syQL+DqF4hcJ6/STTBdRFj
rrPhTMMTDEe34GyshLWEl3eTVO3f9rHlzfyc+Lmvlb2cw4H2upkmWz/ditGDVnYZ0ShvfjKz2zAo
OwCjF9dpJpyXUcUKvou3WW1Z/REiXH60xDRIjns3rUF4el8cHbeCRVk2KULfONHYRsU/mXbqzUyt
mS7am/7Fjw9yNKWhio8Py/B1bgeTMxHTteUxfsgxs8IS3SqzKO7OcBELr+GPrU10ZzzSL62nqd+d
OfPEui0DkUud/vRVwkpw74EuvnpZaFzW5nt1Fl8tRqS3BNdYW5wYT9CCX49+AkVsT0p4AD65WTlI
wYSEZ9zsR2NY3HBDnJIP6bIlrq876e3hvLhOxzJuv4aZXUMWFcl7QILtT3v9J6pvlx60WSIbvVn5
gMTtrjzbGA0+ALuYOjXAMptoBz+v8df2fkbEnyKzgj4SJXVxZEHYl8pFWfgS5DRwMVzG9hd4LUmW
GbUkfqji2uceC/8OBgChzusUHeemL6AIJfYkYq5XLtYgx9sjkKXZyJcJTmR0AaEdEI4XdgY5WKe4
0vL7hQj2+q1YJ04uHvZtCN123Vt0Ixd0v/yXDX8PhIVe3kSkV/B5BgLsCMoU2sKK09gd9jiBjcyO
pKAEOuaTr/0niaQxnY8LvCcLfPVtAd0hNwWFHvmpDQtSd2gfyv0R+qZ2ti6B7Sksm98ncv8FBhMr
PSxYzN5/rBmqPBaXZ/LU9onoJUXR/58S/eSyZBB6s1+9NxUYKmDVKhVbB9XulUYXJCN6GBFRP612
6LoKIcMnX9G6mFQyenFRg28E21TLkBvtKm+mNNig/Nm3qIOrTFta2/pWfERy9RqzEIjoDAUGrQYl
PTuUAYYZ6KPIZDpDFOqjnjhaTcybEV2ZkBbL9jjZa6pM015K2or9dN2JZBdA9LTkYgfYajDRWD5+
lv6sx2HqTIm1ywAXk51C0CtmZYT3Sarwl4QcLCqx2RbKjVU3PXa+c2NSL3hkgXc1/EhFZVzTcS9H
TfSla745ZZ7zDjZoe3xNuVeb1dg8plKlI5hqCKgysIbW7q+hY1LtRH5sP85zVbBTlDjoyOpAF6fo
VcXxNb5tHDzqrKgz5XLq3Xs1ILV+nKF2GDYNtQaU+ZLHZTNgsKxOKqAocmPP44IaTtGWoMj1yUM0
serl8hrlKL7LAVcqa6ReL4MCDh2kDnU578r6Rth42z1x9IgqEA14cZFU91vxNxtd5rcYdklc94c4
TaP+5aJ/qwmHPeiC/CO1OlQpkzEw62Sr3XUQFGXMd7nXkMVCnuy1tjbX2EebfwYrpzLgG/NbNs/5
1wa664ielemAgfCAQFmq1UsATJquYY4W4bzdNDYuce1Nc3ICrQytjHLW8WJlEBIMvjfi2Q9aE28C
57tGnQzPEjpJozslOeOtN5boYr2HDfrdG25mxm27Djh5QgOJY8+ftFEIB/8cFvc504W00r105xBY
vrS4laGiTb6CMqg3Ne5wUCpTB/aOb5FQdgSKQ1S5sjpc2y7eeS6smn1xQRHuJVZ/1Rr38+pQw9H4
VJK1F9IRVNZ3UqcLNFO/OOQSLleXFyRcPr/Pn32dEaxsVMziuRnDv1d43doyB6W8mEAz5H82wndT
mBJNPF4IzSB764VWb3ENL7OTj6dItDqaCUixRw/UnjkBNz/2llqxb6odqDR7LcrbHyj7uwgxSBh4
niJYchh2eB1HaMajnVf99TqTlBJBOOtHU/LxXZd4Y0DvB8ghWTg1YFNWco60QaD2zAjOo/9Q9dZ7
rNd6puf4NnL3ZD7886YwrLA3d5UIHhhh6c+dB8pROKICnjU3rOZ8TL5D4wjyFVE74TbpH/UAvIsE
Lts6t1nVr7+2Gp+1hzaSX7/CnnJ77hNfYflE4kYrBaa54ESu4IwjZUATAfD2aYipz7+EuUIqkZd7
JrV3i2Ud+gbgWZF+k1oJnApU0nFGKZQGGSNLSP6UwzVh0FQPtlYn4MJgLN8sIJZSCpQbo6jRtJZw
UEVJ6dYMPC1CUeMJrvVWk9bOb18LoMOSkKbZpNI0sRNFXD6AmwWpaRvB8rQU1XnQP9gs/HivIOx0
yW7gkgYbzcm8AhexWinwxEzymz45wwWUdh+DFohYBh39BVPgSVGW6Qj2gRTX1Hw9oyltpO5vhI+r
RmpTgSAGyGuo6cEPEUYNr4wgJtH8tENxiLC+6WlYwocCqjaD/Mh1Q8rq1MgravY+Pdf3T4AuINWD
T1eqipfJgsrgXduhIELFMMDhB9a55pTO2pXuKDXy+pE7Cytp0MZgiIRwGC2DrHxcLbEWdUWytfHx
pIA5jpiqqsB9L9HBtALGukeA1PLwzI1jbCyiGQmMywIQtMAk2IHOpMsBGkamlcGBx8D2/sO3A9/j
XopYgFI3+PjU/0UIr592/n7ANZkwpG1EdfrTE51SZ601+dmIpLCtiFpF4lZ/dwYRpHBoGeoy1ctz
0ctuRxPzYBdXTjLK7BPJr78DPUYBykC1keVdJBDvovlzvhAXDy9cD1zqBAF8D+uj23jzg00oiOPi
0OyDRlbyFDTZjw5RJlb8I9rDSD35KkRKWYUvoHd5ec9d3vxnoZaGFIvEAf/ENcRlKS7A/1yw1f6M
wq89JYogjzyl0X/NnCi9UDrY6aIGv7SR0Um9RCNjVXYQinQwPp1kpUD99TaALlelAgL3wZ4doWd4
+uRdHS4CdYWttJtbfb0lK/P8WfmTIMxf6v02eJK3uOiqUBGo3WzKJg5Ld1R5luPy+264Up52t3EB
YLPhif4uLV81U8DBIVF8chxhSFOWrpS9FD708a3ghdxvSKr2dEk3wasJmGfjv8AVV++QHz5j7wgI
umbh6sXZ5iN0n3VEto9qL9qPFOUe9yXYdwwa1pWg4nm8YN0k4ORyC2E+GXyTqN+BfEF5FXiwWmNo
zyzDtlNGAJz1+vOsM1hoHc6g6Q93IcBkU7LNzc+o8sEDCzK/IxliJmC92QSbsOqmdpNtZGvxoACX
xnzowsrbCWLoFoIfcafbEaWPmbOCMiSl8+dUeh7mkM9OROkURdpYhzs1F9Xxs9gV4q78YHxOJnWS
6fvayzvW+b+MBXloKaolzQbQgKrleHGMmTK9YPD5nsXoD2294G7ALmd8d7clIjmuXD5RRCnICmlr
fkE6fsz0jP+uQAJ67hLviAqKeb/aSXh4cRhedQ95LFRvc8xHTjscM4NvOXLx+tRbN7QmNVMkton3
QHu4/6Bmy9/YXFke6WDaEDPMZgUthpnKBY40XWNM5H39OoYo7qUH+fznGl194I7ENG3MEudn3u94
afLOvH/51v5UguLfoKp7M3Wi8f4DjX28VCsl923xM2Kkz9N1GxP9XHyhIjY7fjsUr5rP//BQT9+R
/gKqDps/aeH7jHjl+sYZKhJZ4XQ9vagimu/+mwVQNGhMussScu9dTcwcmmVM0FEs2+Lg+3lY461K
8M5P/BfYNNlP433SdVnT0QEdNIFcl8+LgtfaUTRRZ+2byFN30rx+MouFXrEbJFiCYOF687/5X0I+
PYDQwy0lgs4Z2M3OHaSfumXf8S5j2v+oFh0EnXjMjUEmXRNngBY6l1IFXpp1w2oTpsaHG6rrYo6u
FSqCbzYfDZOPy9EEP4l1dNMgIQkw/eH/Pw61Sc0bUe4nZQLKyZQiPbGTX96XIN1D0JSAystH6+rJ
ZftaYvHVkmU8COa074CNNzQLhxxd8leWOI3v0QpgWIPQcsRaRFTwbevP2ReOK9B6h+9kEMRYmOMZ
iDt3tes7PtmpE9/+QqYnl+oSkxpu273dvEnnH4RKCbehoVcwGauybc8V0KpkW+VuAgu97KGG5NgV
e94D+UA4bGnoLBA2dSGoWL1fZA+2SrUkNT0/ayvQpTXbx/dtpghTfi7wvMBM58lRGPiHZceu1/le
imru7TVK85qMiiQe1apbZy2O6rCZSGJQUVRbkMKsIiB4t2B9LxnBYWEn9TxACSjNxbZT4VdQHgFQ
3RkfsKnbEH7b558QZxdmo866osDiv3yxrvELx3He6dNMxKKEyJN3XyhaaJBwLmGUectfWbK6GTwd
4tkbhOlXNS/6XIdKVtL0b2hpkVMjD9Cnr82U57l4PcPtUnhQCMawFGhFT8zudxRfEpb4pnEeRjto
Jdu9qGwanyw2FZ9zIq96/+0KwkJnQkFPum0F8uq2Bd3DsUyenu5UAWAKZGkaXAiVgJkyL/+vqTdd
Ctkn00GAQD0KSNwlZAB0qjAgrD4ijukrLPJq/Pp5TafmPEYgU6h7Q/850hRiffBIRCuLfUBFi7RU
WISVssH+qfXTW2knmGCDHVwDhvMDQFW5b1ax23El63A2yw58tMeFwPRskJ80Iy2KHYdA2WblrLbM
qpv1MM+tgyF4pwRCInbZQJnsR/FjQ1uj6nXpcY2yMSESZw9ycLn+xr5Re1yUarTK4vDr6mFvOpnw
2Uk8PCFIQ4RAiUT5/CE4Li6f9n7bRROV6HhoPC61/ExATikGwXmmGsrANQmNe6oCU5W4/jSNCq8t
vDudiXbmNs0auszvMjCqOl2IaB15LN2j0NesvWYQ1eAyayGo8hqf8mUKQfmW0sLu1Ky7kb0J9WOb
2eNo4r2eJYE7fk6NLQGOwavaWwSwiiozot8oEGUKlk82RB8hUKgisrB5rREK33A3oKtLYx/0l8Tf
yiKXDGvo/cOipV23gxYOBp/fYWNYlO+POnVeo/sXPI2dse+b34m/Zh4e10VYlgyv+nclyjT8pBP/
MphWRp0xgnUI+MZ3XA6rBJJD8nOsBQJ/orOKIF3ZS/T69kFRs/jJj9WZimfrmKzlSvWMBPO0fLA9
BnlqyUIhU3UsUBWJdwPDdIJj5cqdLGuPa2gArR/BC7ySEl2wfmYSfM9OaN6OvYHVp7rqjeyOCr3o
iPsFjc+8vvko10s+pecunGvKSDCxX796csDCP4AV8d5iZ5CiTRSllUpi5Jopa7iA1WLhl2H6zVJ1
zCs5Nz8pqK5kwTiFV52kNXg9dZrHcNRa84nUyzvZnEPcL+LgaMotML86Vr6NeCbiZ+/EMMugTtjt
i7Zqvrye3G7ZOwVbBGEcNVPvy2o2VBE3VQ0TwzQarvOYOH2gw+2OfoRVukCKoGChhudr1ptrBzEN
j3hJZiZAyJoYkbBM0RccyffdUtH/VYVHSvmKooOSUk2Qz6uKzaTbZ7CUHbFdNloakeSC1Bca8D4C
bmIOMuuu98mldxLcKxavqSg2k9jCHXVxFzbHl6Ct1wPE3yk2TkNIDzJ/kYlYAlQ48xa0lCpXOsdc
Rq41nJOVwimVvWKEddAG3hoSsHNb/Hr/AwDNcIh2/9/d1eBJNWGs/Vr/fbHMH+r6BU6oORhC9Lf7
6Ri7FzCncxYRL2a5FEXCTjIaxX3FrEDWV37l8+3+9xdwBmmVxT50jz5Rh2D6sk/WjLvUJKyp5VCm
/Bv4Mrk9OlFnPJzLji7kDk9093mMFHd8BJOxuC4OFFtrqpTCSBJZDpJ6/573ZAPjn9/qYapN1/94
Rq+HcQuYeXVO60S7h4s7YaG9rFFNAgwjHiCr3enNxuMxlxiw5s921zg53NOSrxCDkzqP+xgO9IDs
A6N89U7JgDOfEuwUn4166dmiT1hJad09fIFll7V4G03usrKsmmUPEEWmeRly1HORqGyR7GtezAu3
41OzH68iPTuBtnAq5xZnj7VF9NyS6cGLi9Lv8Kyaej3TRKZztgugsDWax7P3pLLVx15AdOX0fdis
bUqfd2pQxtusVwWa+SdaUa+MDAM4JwCv4KphNOhbUgYVB/CoUMOcYWE5ox63eBS8Jxi9/hvF3AnS
D+ypcWI6YdWTv9oCX9O/r+pPqAanCrcvlzm0LxGfnFgzJQK1lL4t4YJxIH5sngNk4TYv5g9Q0o2Z
GPteyn1ijKBrU1H1j3/e0mZLK2ZGrrTTz46U41AZYSn5DravCk7GBZar1AWrcpWV3lREEcGRkft3
EbmYuUDKldtlz+9RQQ3fr+tj1CzKM1tkjVyzYRzmfNJha9dA8KIhb0MFU1G5uKGae6evncjdQLR/
meBPtTl9TSmHW7Q+KV8vTXxIwF+p4FkRxqBqUGOJREqxRKEbgVFGCvIjkQsqk46x/5z55zOMD+ra
nFL7nQB84Z/AgL9DRcN8/QdaY2RJe0PsgTiKMEPoe1EpR6XAo8jGO5J8dc592Qla/dquAa85cKWr
zLmDgJ41tuByhszpWMD2+K1Lp0Svb6N8jB7gAZrF1a42sgxjBiXZAs/+p2jJhryuYc3hH/JOFFg4
5C/H7XHYiyUWIIlZpSQJIz1dGD0Gd1gYHi2M4gbqgDpt5v2LPpi+lbmhy7adGuNk4sm7v1yOAQBf
tuJfGIi8DmkmNGNgF6Ze/D2ZzLMdq4cpmc6KeJOFbwH4k4e7rT7e7NjjpK8KuBXjZ7db5Li9gq04
7FMS4ABbJu21Xg2A1pGt2JXXItkNc/ijitdfZgS6UhSN5y31fvjNwtKeyGC60qQnddi6clAqGxXn
aXNhOQJxKMUZUPhkst8x5OEiHcT2qPyUEp/lP46iqKzn/ZB4MJib2dDcMD2ad59uIB8VyTA798qY
VCPJKG34UgUV80ZzECqEaKjywARqzN7HZGXcw47uSU3+1hWMl5TsIBvojIWg1iGdbUYyasJkDa80
i4X+xJFPkwErp//1NGRaiK3sCqDkkrgeYP/8wfhgYUXxKdYgmt+1AdHl92AQz29S+7L5OeSsChoW
/qhfqW4SFbzGkoUEweLaW/Twx0c6ZZREoFn21/yLdyYcmdlWdOn0HBWKPeHnvZlxWJeH1x9jFfTw
JGtOmYv+dSsxjk3wa3qK+Gwntz6m5Cq08kcWIG6dygXS07w9cnqKVgvPv0hgznHyLMlBf22/RGNy
UL3++DCrT0nTv6D5s9vrZR+lOfU3oJikpW9IrJuSxv57QH+L5/JJVOdhgU/AdonKi/hxz8VDaMPP
oZpHwFlXq2W6KzM2Vu5wmvC77uWi/AfsJ8czMntY1f4wKN/pGidRPzjVtIXwTMNdpmhFbUnD8hD8
XYzE1ggnV9BpF6TaLpO7S13bXutjB/HuXqCWr6qzw5X2kaQR7CXmzK2y4XBOZdfdwlmdMXWjeJEW
iOOsYwSyiZvGY7Zpztuno2SkzKIudVhnv+88f2oiBy4ZxWjF3LHdXNowKgIc/r89i/M3PdIsg14G
Sk4X7lEDNz8F0Hg1+uzpOsOHFwoJVZbBjV1ywPaM0sVjQWpVlISGUoG52wEYwmTvt6J9cPBiyqEW
c2jL+WnwSIUMQTbnPmIC5Rrs3xjKz8rFcyB+QqWzSKbYPKvH4anVyUU2D/lPzTbU9f0f2zVzfgpR
dt/NdWnNHL7pdjW3IPdEZMvsg067xiL86FBZDAv2npEQJ+hQJWQ2Me+QEziWqCzM1YJ+o4z+aPI7
89cepQONhYIledvYUrZkmVzPNTC/XKa0s5IEIyNw0tMsJdlnRCcmsxIavU0Cxq50W7e9Xk0w0eXJ
ni0UG0vRhPDrdkuxruz6t+EMFFQU2CkEi/VYXFQnBtp4+QQicJcH9VDXmPG/x9DD5MFsZtPJDtVG
o1klvYra6gjn6iBrNgvQ9ImKqsmToIFjoZU2nfbSiGu4GMwYl2u3z8GvG0+7VqTeJIo/JREFBBEG
alVQhG24qk0o1QYRH2BC0e1etCeTkkqmwLl0+08pUav4iNhv8q/ZT4vpjGZEft4FYHDAYVA15XAe
xJMr5NnZuNjkHI8qx8EJfVAPCX5pyaS01zikLUeKfAuynFnAVL7bz2coyyzAKYAX8W8hzJZWaRzN
3AZjwrb5+cIo1U0fMFp8eOyOg+xRCMh2ur4RAareVUgkD7iQQzlB6bohuUbrc+2Uc5oeoOUQqzAw
DwZplG3d1Glc71uQtB5kh2QcHG+l6Tnf1CGmpgJIqNAHgkhC8aByFfYDq/WBvHmLB6QkV9DS00GT
dKLQDgESH02dytLwvyMJpmSy77waJn0rqdx1eUH6x2+BWQwdpnK56DxJD/DBDkoFdywxmY34X8Z8
FivPbglYhmqQ7WvuvPndJ67icMEOl4Av7/OXUD2B1tOB2joP0mbe7GzFaKOXPZ8hfJSB1jgQb6vX
POFlYuwJcLlw641WZKYK94S+j3eL5Dc1H1rah/W4GPoJeM/gMKk6TrGq7VDsLFKPI1c5HH6MB9Bk
+Gy6N5VbrrL7ENre5iOjVJ1qQS8xyScsAQR6+4SExPORVorHpJawX5XyakLTDSgZ78/3IRa5Izwq
Mp/Gp4BQ8G4uVNgx5wE4jM6hcvqVMSUJrAUoBaFNByNeIYrQ6S84/s2iF/eRpfrTYVVKT6jdqTB8
sKT+fsjHaDpPRm/5gwNXsktPf5pQu75Y+Tuu4EJz+IHvr/iN+UsG135MTxV2JlmpzUtfpdy41px5
VYJDD/BDCF2UzyR56laqSQ/MTU8XSLJVq9c4V4lhLqhVyj6ugYB41JflX6ZtM3/qC2FFhdkzsPGf
1R0hhBndf+2xjfKQwMPcPvyJUbFKUSq3ylSWXQH6kzomLKfNEdRhUyHluI9SBqSAyK1ErgiKZKli
TQi6g/oR6moPFTUA0gNRGP81lin3RsEvey44ijRrD+8UHAAg8IOL7lrezKBCyVoXb3goWv8W8I4F
68X1uLTeUr1yNC/KNQ1D8Yea/dtrHn0W0WB7L7JrL3595pxKUhUIohHo6IDZjWJEjUlLKPGUkRc7
1fziyyUDYeZ9JqWD1ru80iUuqfAulLyi+cxCz40iUsuSJymQEgYI/0njB5fo3xETePbNdFz6apxi
uh81x7wxliFxgk6lw4u3R6Xz0kmzBGNqAOw7NpIXHDtlDVR5rKr4wSupCTbgCtCXVG0bFEEOTGFX
aNptBUx8B3GyGUO/WaWV1txOWCWQjag7xsONMJPtv7JONjzxWowGXmW62wxWp2LQxL5cGSKMTrHx
aRUJY9x5sBpUZt7ElMGhIXR8vHAfPM+F/BGMFmL5BdE3AGf/ZQMqRs4hd2s4Cs78NRjH1srUNqB9
OCBJZjOLk30iXZWR1nBHXQjkHoMAz7SkG6JjnnImzFPeS/xBhNKd9VPABbXvz/uwoi6Bz4TB+ITd
hD1KQdy6OQy7oHy49ZIsaXyECF0vxsy44VX4m6MSF+WKUknnMIrQhltPj6AWHO29daAoC470sF17
QuupyNkg8D4DS1oHs8TtGBqhFufWP1Jp4kyd3bEBMQBuvHzlKqY9i1UWrFGXgoRh1VBXm2njskoO
cclGwijVEmiYW3xHCrue3Dd/01SZaos2lbP9NEWsc+KeeQEuIz0wSn1qJ4YGOJXHAJWJFtoUyffO
5nc+PPbnyvysN+MWJVPgxg6niCs3okUfoVsQMtkrfSdXBkh74T/hMJH0qjUgcWqf/XKV3Je69kBe
qyhRj1CM0F7ynYI/4sKEpGsyI1KIf0kErOIznq1Q+y4j7WAeJAR4iRZBuOojgURpZGhz35jyF260
vxZ18A0wLE8dz2vABJQGs3Xehqkb2P4jTGOXT1QrsPbHV7ZofxZwpLozC8mxEmEucjAmKx7wtO0p
q9i4INOAMGT4JXAfucij/fRIwZmaqy3uP3ABnqPqw6BxHiFCmMe4OA98do1vhHYudWO/NiuIblcv
GAUhcyZJrowTE3DV9kYe0rFkPXv4AszLWbJPFNIZFu31ryUpn6zN4bi4CMqYUW4b+qJG9BG7bD9j
s9eELUdFqeW1Qa5cU1xPJ25AE2VHco8Ya1CUziu5uR+ORYJs+LVszHfL/NM8DK0P/dP+tofJHAH4
XTezpqmsjhoRnXjRvhojXUsA0JbNfq5nTQQfn4UYvhRFqAwu+cmNf+ZAS9pGB8zLhI/0j0aDzlRI
8XAjmTtkzjWAWY2B/F////X4MUTeGQvH5oT83Q1igdwNvDEgywEmOyTclgZmhRksp7a8Tdca2xcp
7HWEFoDhVRTrwcZ7TACurAmg1YEkwmBw+C01PElDJ2/LsFLiwVm5kbNlEIDBvCipmZrr/yFhDje+
YS/U+j5QzHPbzLWurSmOtCndQTGLZ5lLccPg+1GFhWzdIpBuikKR5AvxhH9mcd8CtFo2mA/PlqzZ
A7jPVBu5vNjR0qR0Me8d4QMYiu2k9F/AuHhyKWFDv3e7X+6HS/9bTQmj8ceNBYB2aUi0Iv0xaypa
U2A6d9cuUDBRxK8odKgEc4XKZZamDh8Zec6WCgz2pO65d8cCcqOHDadY/p5GX8vNhT7bXygbXR6C
MbH/0UKyGR3Ue4WVyn07IWQ2W+B8FIS1SNPhM2URu80ZjpPMzwPNBhSkJEhFY4gby/qmjTfqTNPw
BvQYKPqIrYDmASuAFWi26UvCUJCvw6eBiTQ8s0P1qWL7UeTj1Yr1ub1UzqDLcmWB8QkJUdyAQM/O
xy0hELj2ja0+/7WT0BDGWmgjZYHxhycBUZP7qTT+123Xw1u/G+NEeYY49wUyUvSrOiPqyc8a85sI
vdkk8D4WHnuiWsI8ImJibnOI35w6yw34jVnZiaMAlUn7IkSKy6/UOdT3KuUSXuV+lNUL0NnTMD86
4zRaca40a5XF1F7YTO1CsZXP8+0HZw9JFdRlroIIuxndEXAAwOO1MrVxRWq/xHCM6XmfSeMMi/s8
7k/MkIwiTXoBjTynPzS4DY5tiS3zg6JHQW6V+RvJkn7I29zrZj/Svl4FB1ts2xZn7hbTJ6p1eIBX
ctk4lzNNkw1zL2oogWzVy8xuwKtXriZbL66PuZ0Gho0DyiHDxgENOmPgrADXvlRBVsWaGyVyjPje
+fey1A+jw88H4kPp79AZUtxdSKZwY0qbdmFIZdJQCJsqhoZG01o20/wJ2xRYjDJveMLrUEs7htud
my1g1N8tDqIS8wnC4YunKuz0F1TfcNiG1kBRaxwXKSZKyCyvEzkTR2YalImakn9DKlI1iaLFRnay
1kZKQn+WE4OOAp+KNtOWtvD24L2qL/hkZH3mLu+A8AVoFF7KK2bvkuNp43WvLXUz8LZigaEtqR67
jvne8Qbf84/42pGRdOiR8XyqPZWaBzJlnjr98QZsbmoeqmofq3YuRy8/F77ICQ8DZCrsOxPBREob
4syhjqtyrDeK72QFNyfHFLB0Jk4DhuX0RU5/0pLztWvu0li9Xfh0GEjP2jY7S4LCH+E2j89fjZY1
WbzMCVwY+xsPOwLgAS1ZzbRVS5Ivujwpva6KG0urKXwmWWujyLOUruQiehKeKzQ8yMZSTfoP2ew5
d+9tGRi4nmuR/uDoY6sl8lev/RH66jlG4xCYHFnwv4Lm7s3cjRyJ2RhIhhpDt5VtUtri8GHT4TBZ
ztTFWf8vgcgg7Yk4DST4ip9S7rcFKj5nlUKKAo/ge+CraKt7tRniQ4FiUgnrGq7qqQTJy1ngkHp0
ZQyN7q0i7s6K2t2Ez97vtUexK76R67Es4znaoxSgDcThJh9AA9xEDiuOIG0nwptwMguLQDy6ocRO
tzalVSDiW+8WO8wwWEKbE9nFr6AAJv7uvT8Ac67759TRCueTnXiI1KgsRZQUFJ2jlJxJ+cpBIfd6
MeYrcFi2fCDGuzDy2gIMRs7Ducawy6rEsYlMFLW+SsLVZn+9kYlru01TrEPB7z+fsxA5X65MzsZl
/NiAI+zXod7aRjvuH6e34QKkAqtsZ6l6W62FQVETWiduzHyldx7UcuMlxtypKAKCj9o40LpBneai
5fMR0rzBg7nVbug/yh9GTFD5FizVN+AhtQlkarPlqabyFBWE4l3MOjeVLmaAB+mpmuREJ0F/0rZV
eiTG2iMiHesdYfRaQFvISaQcJ7yxJccPHuWj+6sK7Poc6IcXvcfFSZ2x7WmBmcSJ+EIEeyeInEGu
8GddaL4/tW6DaMEii0FIKeGmCXeJivYWSbQ324GuXrz0559V20FXCYHvaY4eMp48DhJG8HEOkGiM
xERMaQ9Kn6JSoWDB+6QfC4sDq5wjv0f/yzDtXBT4Jsu7Le0mrPFrYfogES09vnM/gZFCiGCd8YjG
NZhS2WsUWNd1ESQYWNQnJ2HFEAfn434P91XSrFxp4CvYnyItblBgrlIU0IcfvVOU7nz8Kh8PyBpe
fJ/sTUVpo7Rc9xDlsFE/GDahYCVcvKduF/mkuVhMm33dF1myiGRRVKutPw2a+nuo6e8LG7Lo9FkO
3/THDUcR+nO96ZXrpJBw8luBzsD8ldCHHJgCHs8AmCJDITYaNyxMJ39R/c4/DGW9vMsHVJHWuNpn
UB8w99PcaIkxe0HMGg/43SNflUCbYs3+JNuavWBHEnFFfPvgj6olrTpKo2j+GlAAUavpNCv/If6d
b7X3PFk4BJ0bGzg911f9WUXD1QihAH+qFTxhiXoJrNKDVOJuMtc05sEJb4QcL7kInZqtlOdDbsQ/
p5QcN0y73HUdkzSzrSKpVEr0GN7yT1zGv/YZ2xpbicy9ntLpQ4pbfOXvmgtctPrgTjZ6XoII0Gri
gTX1Eog8rhrm+Navh8IWVsEyZYdVCeL3QwE9LEx+T6GwNiqP17BjIBI1kYP0Z82DAMXiinVyQFCV
eACGV/9tyv188jf/zgmiZE32sQfzqdMCdNSpKtRq7weIMvSt7MqDrIv2YvWl5SGWOGsI/n4VgmLX
pgp2iq5zAP0ZGty8wAUjYKblN0Py/EVMu+Yu5RnjNzV0C3+b1kXc1ORr7jBT5bW//iGKJ0clqIFv
bbpbUfepVTfsSjMr5Oqy8tWaDxfv3JO344meOkxYeCZH2deTyKbHAm+qfcXF6Akh54NEyaandvwf
WxZpph3Wc8TWlqpXYWdeCNHI3I72Tm6cMr2Pg5a3LPu8qKLS/Ci4GBulPscB7ziJT8gmVLVrgZ/q
ltOO16yVYQ9PbIlL3gNmVj+jCyL++TF/4KqPel9DU9g941gXqGgMbJr35y8ykAa0r7dqXDwFCvCp
g1TPDUgsGJGLHteeCZd25ayx2zZPEQpciCnp/BbTUolYZqVL43CPGOgwPPbwaF+ogsd3NuldCz7T
d29uENp6D8eadskDuxry/oeJlNtzCA6y1HzW6oYFUmmHyb6WQ1i7THt/5Iaupp0dJCJT4Tn9vG7F
uU1h+IHsSDo7+ZreBqqeMoSCJzxktNv0Vc0MZG1EzVJd28hs+IZrsuirBKCKG5AIBcybdmmKp5Td
eYkrkeFW/kly+vNPXaMgkEG0qabk9gnZeniAKHAnNgZ+3yNMtSyjQrdmO32EGJy7ZcMaNg8f6Snj
q/fP+gYB9sCer/mWP8AVv66K0b70UCo0JN4FNYqPLopesqhWjWZHWZYkOXq/AbTbb5pv7s3AkvUY
AKDVwOesRCfNi5YBxHO76AaLKVkk+QY+Y5P8HwQfvMIpXEk3Mx++KH9PTFsmepKOMOuHKOFQJCTY
7zFoXiV25lYfm5jCF206WhY2UtiUDrQ7E7wXGoV5XNIbXra9Cyt2+uWV7b2ryrBM9IEkUS6ZK4WE
si+ctkjGZyWkruTnaLh7ball+yn781/FRLp5bjI93JcYBXMU9h3T1lzKXDq8gJxuP8o14hh9cxOj
jd8PYgfClUXQn25wX3Use1iR4qYsbdrUyLG30vr+IkO+FyIeiF0TkQPWSN3pKdKRuJsPgSmOlB0O
D8qsGcwnS5GJzl/cceLlyw1f9DQBf+Xna+vhlEUbPEkrRt95iVKFhJ/303qZ/ffiOOf8kcCp3tW1
m0ORLRRXX86eciknwrlmMTtDWddjkyUQ16NX8z5AzwwOfmd0brb/eTMqrN2AXTGLWhi7DO1jDtlT
9A4UxVb9OSnI2Z0YfD62I8Z9LwebLs6qFobxCivBvtSTJnPMkZD2ewPDxGGk4zRcuADywwiyAmt9
/pkPtfi/tgOHUVchxumviwv1vko9K0QqL/nRJP/GSmM34bjUtTWBNXPQHyDkdhnJ9xYwsK99kpDl
lDNH8hb0u+xyX9a3210nqTsRjagdUsg3aNIwvv9C6aqOLbEMc5bhnATt5aeym1/vMMdmy8fc/iE9
1z+NtScB3KorInlNKCTbJiY0EztlH6tNrnci6RTUNaCUgfBh8GrQiHm4PK6yirFzcouwHa/fdnaW
k4UABqNKuOS/P0dgORkMelLzHm+nNg96Ou/nGmEVAMhXLtsOVn18QkTysqRDvf5/i/+b5TWxlakN
yk4c8IueVpOWkw4iYWXMJyEzAgSczOOcYp6h+j4cqEzcNLwM8dj923RNRL2WW7rQuifFyo8zqTb+
6EC5ZyFseG1QUtgEmWwPcX84rsND4tn8pOxUJu4zPhGaqsYXexfDGRosXUIpsI9jwUfcRvHxak3q
M7ztkKDz6auGMGbm0DHH8p2RV3cqBL/BcfXb80tfcLyShzNkPldRKkaLXEH27uO8Cn/cCJUBxAlP
VF+xZwUbNDm0GB47ZUTZ0+zk7PdaaUsrMgk3Ovzc6YY7thuyRyqmTQFU34ZmAE2SfH1Wn3zQ+Hw6
nm16v3+NiqrOdukJeVEyAUBTdHORh4W74GSNopf9c+uXN6A6947bPKnv0lciGB53ei2aoPaOCb8z
HcNhGx5Y2e25wKJG6nwjn9KvAC8AIROfCJqLbZ3KJfdWLqKu5BTfRpTUsfPCZAXA9dHT9quzgg8b
PcOMkezAcsWWka8YmOCrqnUHyJij/eKnvsrRhOM3CuBIDTdLfZWRZHGq7RI/SbmGpDIMOcgv39dq
4N9Z9APxKdDVzHmuZL8Y5JRbqVw8/7kwz5clxanmlcpJmtfNEqrZIHXkpPE2PKoRff4wQuDjli+J
GDykeYKPeSGY54jRcc+J3JOSnKrJSVx8s4k6FiL0P2rmmfC36oZK6ya93bDXVI8xeohTNqpDCE6Y
8oBKx3gX5SuBxPuHFoK2xnK1O+INGoW2H/yDKrwuTBwHAhg0yZRrr5qNR+R6nJYXtiZAaI95snQF
+v+Ce0GaTAY2QXySiS77ZY/etwHHR53TwF+36jaYXd4Zp35zXD5jJBw6oU1SWV7pIlXhSwRP0WJy
eGk+tKQReH0AlJLsJjT65pGhjxJY81O4AH6CBrBbjWBM8euNEP8CE8cPcAvCZUdCras4OxjS7sFK
OPXTkg9AmfsCEiANzgD3sh+t7I1KYo4pB5mCNOrwIRZ0KOfnRy8AbTG+rp/PrOLqP3J/giMWnjwf
euVroBaj/vB8/aYCdC6Q/ka6lbgtOeDUQ5rmmTFKw0HUhswe2FQaV0eufWU1dfo6IxRp5FQ/pO8F
IQ19GVQcV4OsOlhbBVq1IKHmfD+/INnGO0M+sLd7dGxGN0qjX7Qmp9b81mmV7Y3geXQtdQ81/uOr
0joV15uBACgiUOnZyFlOY7Z3Ws1lwbOQgkoD6XZn7XaeDsThlzbYcbNwwE/5aqY45S260XbPEYOm
62KBK7cRDQin7YEQhyg9a7rQbROKbRbI3fFUfPsFJgo24qtavTucgauUvYzi0upfW73pVGcYp1UW
mTkTYhOPFIacYRurB8ji6RBr4JGtMWdAWhrivR1DVrSKCIQ8czBr06hcymf2Nc88Fjnzdr4rDEav
vqXob3YkBHx9dUIoWMNYh6g+CeyHJroctPqd0Sex9GCD90AfsC6VGzHM4PjMy6uCZZDfzkuoaCw5
VooukwjvUY2zxmc+8fsGgC/UHvCZCvtUTKKisRGJejmCW4PS30c7LSwXEUXHqKXU9QdaAPt3A97T
wY+U/AFeATRBAj9ZG7ouI93g1zZ8f/X5O60ARzSEZHeYW+ZyVJgXNl0KdTCEU9ZxC+b+sKW0Dk0c
spwYS1ffeGGLkAXnddPGKyanATE/QtlGhCwyDUFroIDgwUglrv6VF1mGjZnD0Ltq56tbZc5OS8SE
XeXZSHm2htARFYqxrIrbOWiG4ldH+boMTilpbQvcf6gfoIQcyFFF2BXANlgjx6/iJUuyASK03bBA
Qi816ldmsdzn9fC/XpViFiedNUQ4fZmfXUbiA6Epz0GoD3/yh/SbIzGtcDzL6BUjahC94ezQyFUB
uh1qtrAuT4i0pAPrkYE7HoGmj2Cuz+cOZlm8GOvuieieC/UQcRqaMmxPlaOEtLimoGSVq/fWNmWS
erRu4QB0yOZgdAuJnHZ99GTmmgaeJk7tcO/y4kk6JkYfJAJBhxz7E1UGe/ILjvPPYzCCPJntjL2G
9Y3rn6Em3NzUJkFdFHe7xHEWWDOTpTJMK+LhhdCWQoxGy+AhcLIuo5ZaC9enNlS8S+l0oqzoNM3K
awQc4p/3dGQ27U5t5rGrat8U8W/jIZgUURr3dZS+u5sJraORX6rO63Uxdxej5j6vUwKS+556G1Hf
rNxo8vwJdZxEJmqEBEl6+SJVDQeNrA4528e2q5mBCzsjKzEmzzvsMiWS1MsqYamkemdMovscFY/R
keMnSxfDq0il2N/3kT79o2FugJWz1XraGvjne8wdVsF/gi4403NtBdU1ZJzCWKIpVqZ5YUZyTpNm
epOIb09FXmizi4snQS2rY2v4S7yv28yZIw60IqN61blByAHl+UxwitO967a+Cy621OKaqkykxPwR
aCIeE6MU8v3zBhn/P3U1HdbtE4WNHdPPcBF0RHOed8RLCutaViscDAPRhRD3j/lFb6EdGu0Zwbq3
YqyY/s1B4DyZzfwUPTfyUeo0mTXNLpCLansYfsnkX8VRy8p0NgmaU022mLbOuzL6YiZh2xd1G0PF
orrUzq1uch2u3fjzmjUbhhygMPVllIGPi3TPvSWAekkAnz0+9hw2YJBRzUvo29w6rLxDSpKZfgE8
xYawJQjWN62qeUTaau4FPaiMu5d31SfqICEs/zIOLELQA9kPRfiFhI3zx3xdK0Z+tbh+WhW4IDQE
XoVJpQkEL3Bqv7NxkIR97Rq6NllfsVvBEs7o5jkYku7J70nIqzTNu5fJ2zX7/JoZJGVuqsNdQM2N
J4EhpXnGciTrddWB//jmxQ0npNITiLM5aNo4CksWGJIr8t0CqcBhJRNC8YJYIu1K3C2/KNIzuvfp
+SSVWXjQdFUaotJkKnedzkDcKxUDQbag8mA26ccJhoykBo0CJv+0hWzejPuW3jRTVUMH+nRIASEn
gZtozOX7iY77ciI+rTXHWKWX9ASpVt7xS0e4TuToq/e9mMf5W9iB82983nAnuoAhqJWjcKszEWO0
g9XDbVrEb8EsiQxtbccX7yNhOqTiZCmavW+Dujwmgw4RRdzJ4J6LqfdqD6Uus0LzvgvE/lpKQP+7
jNMfi8hWy977t/8gKCSiXBcxNAdAmPZBo5eCffh2mJ8dd87Hwt+J0VgpF8R74Uq7dfXFafjH7neI
P+HDTvNcfWB9gWGq/7MgcRSNfd3VTxOLnHUtVP+qfwxROJ+oPbsA0cWS6pSBLBLLVitSg6IeNikC
gSt1TInF9Av3jR9Q+pDq2v4QdoEQYFAYXlN6P2fpAa+qPoLjnNb6n07Ud4QyoNFMcFbsNsGrVJE0
YroVoEirJlofbmLUeNkz5l+aDXZ/k/k7PMCJFZPLzA8y8b/fSnKA4ids0NGmVOiCLmO51dZvndf9
8uTOmj7cxvQ3SOvwaXresAnq1FBInF8d5X/EVZex4DHfsKomhICjRL20GK1Dd7+lDCfz3kI0WFn3
J+eU+h/X74X/Dl1qKXAa3YsaUg73362xrugFhntq+0Po5xT1pTO5AwAAbem6dKvFk+2jmzIZ3S25
FyrSicVyXNWLoLqDZ5PG7sY3Z0gOIUiy/SNsZY488JgD6C+uuLWmYRRvTESks/L/loM3HtBJrjdg
FNuizpwPrTiIWL9N5JWpqEjSvHyQLAu4N3M4qVYeO6I+h/d6V5X4tfjbUnYaOC3CWLAip9PSzUMi
t6uZjenftTA7mufoGsTIKfCwnI3hccvFBsP3A+9MDwE6VjzxBasvXUjAjgdWMje4DWhwdYTx9nix
lrKmGcwmvEjIPQMORSG8ROpci2A+KXJs8CXm9EPWJ5cr0OIj+F2zC0SAl08UL1zIhJyRf2kEl4B+
qqTJUvsWVbKVkr4IXuh15dqS8h/ocmujxLl5n+y+AYhcDHnLGU3diVYUNxfyjHE4ZHgE4G5TxBE1
is1BAqL1kqPwCPSqA30C/K51pBkbwXW/u42ZTGUAV3ExjvSgwBic5RNhsXTHmTKURF+lB5awwaDV
ugKHeAvrDli6B3W27htS0FK6Y+WhhNpGNBpkphqtTZJOM983//P5b6uQHjCbyBNa+z7W2MlrR77x
mNjCrPHK1KDTlVtxoMU4+cpbr+fxuF9UF8G8ku1KNNZb4GAUC0iUXl9S5LVS5bQ3wiG21vKeuXst
tb3ldpXFG6K6PL7Rz+pe3a+vPqQbjGtdz6GCPZf763Nd1dZ8nz8RULQeTRxKAiC2RbSxGy0JxIXy
h1jRy1tWEC5KQt4BllyDlmEEHDV+yePbfVaajF2maihInwcPxeSxpz7fiXVqwuGKIBYkLbnHQoQd
fbDGdZqQsTeYGvTVKPzjvL2NSYzXvF8oxh8pkmqtIiZA9T7ASzJrG5BNhSzLI5/6LCm3et2qjK22
MmYIHkJypypzY7n6ykha2vibOpmYRDUiX9e+rp7Z8WUxCqCIRpZhGkBq9SUc3/Z+8IMmKU3HdwTh
G2h5CpFM2mkfGHnp3ETYPXVtesusN5NpCJIBn362ny1O/GZtjNdE9uXFmrtW2B7zyqrAjbGCGQQa
Fl93ntF1fa+6QDFBPerLw75kmNpI2AQveknIGy9Bs23NYYX1IG60OKDfIykJpAncfCHhQ4AbQ+yR
D1Dmu6M22S8X5xPLaOlmFSBR7SrDm8SF/pD8AOosxeV7zm6mxQdupLw53gml3vaRUMsFSEWuWJZ8
G3syoodEYV03taR5D89fC4/5aQyn8Ci8P0Tx1Dlzm4sYmycGClMu3zB7VNZT+Sf8SGjJDLwreKT/
M9aRq8bwZiyz2G4fXT7qDfkt2ilhOze6LzLGDQEsJw5NlC1DXsX4wE4PxClNnB/QhnuP1S3wXcs8
3rHoXjqvGoKoTTl6SH+RhnnGP2VVPnRK3L3YLxIUmc2/zYUxf43bO+4pWvt1r/gxt1M4rqdecHTD
5pGIWiOwZjt4FAR+/Dg7ae7eTKuJRkt78oCxUGe7qBHM43DY0hKbCWtu7vmQfpFrHn6Jc7OyndoY
E1emmVlWfIUr9KXvFxOPqoxOHxIK4Mq9CK/FE+3m/08S1WGtCBXM6LE//OjoNyNe5xhv1QWRoX3c
tHoPnHcWaoK20o7VNLh7Sg03s5ZTrH/+OWdyDkKf5VWEWbLp4Khg7ga+/pWMiQjuZZFM303cXoCT
YkDwhBFb9UIYDQWRPGdaIYwqnLeRz7QNR5yOo73FqGZ7QAriTACgJgxgdYyJvyMteqV6NiBgwdep
ywzqQpsX2pJ9cVtP/VnWm2ONpilm3IG5CRrkNgouwHcXfxah9cWEy8h/whMr9CGHpnKeejV13cD5
J8ajjkApxX2ON0qJKxTk4dZxj8dOfEgPEKWfoOi5UVGO8jR5WeDl3jFyqbAB0n4ib9ibRy+j8SqU
DqJPisKK71D+3KAOcEtQ/15rXMw5SsTUGBQhOif7zuxG8OpFXMKJmc7yn25Cb4Zl0awSNHuMN469
C8RNm4UZ3tPp2kAPDgV1hOIyOLtREV5niLk0ZR+fLK4TJiJa/9VxMbQzGLBoBQe6+VDZjYqfh6wQ
LS/wgpAjolu2S9zliP+5rSdUFWRHaic9fw1QG7WVYcMoZXUl4kYTx8mlAnwth74BTMK2mfiIEfAZ
NV2hF9auqHSYWkaiSXvGS+dsO5fU6jn5oDOjeIiCAYSfJc6eeXrhthyM8Vju24miHVZtI/ngnKOf
FO0SKMB/wlVLjz0CDL3RtmNbwTVK4QFekbb6w2bIh9xiN0i4GLNykRCXHF9ysCZ1DJjX3n9S/IsA
LZjsEr0al2WQGYAqIaX+SIuMejaKsVrqGihkC8Y51x32F4IzaRWwdBXCKnhJ4lwsZx4pJ/L6cyfc
RoznOjUnaEQ+xOab3jTbBji/+omppre0SPmGLc/e4X8DekEQiYP+n64rMej5DIShAc+UT/vpKmAC
/CWYkpsOwwuXnYg3iDv6t0ZYkObbJgoO6v1ri/pRHa8Q3RI71wKu5+8SG+HUg9ZuQoeQjcdeSE1R
qx3vJmW0wCzXK0IQgLqHKo6ed0ATwNK+9wabxdCGyRwxqb3/45Mk82KR3vTMCO1Z1ka9O+VVaH4k
whdZWlP28EP9kbzLRJrSSTEpIPnRRfOt974kOaAHJuQZaZ5EaiphmQpmVwD/kwhETiu8s7PD+tjV
8DmvLgNOH+19TEvHO9QXQlaGz+RlsFGQWGAtOtuU3ijmE0BeQo6peRiEVE+uka4DNupgwFpGhuX1
WzsvaJsY5k3JWLqe7B8CZA07cAiCu9L68yw3OtpKa/OTdDftz7W2IGE4sg+bUULQmJ8pTT2hMzoR
E3wRIWybvkDQI/9ykjm+ozCG/JwMqPJO+keTGCPaveoh48/es4Xhc3m2A8p072ksid/PKnh8dtPv
FE4X3QiYUHgpTYrCqvNRIAB3kGspXtvq/4hof030lQ51rnK0XWd6tW+oY/DpgCZHzbfGEbFsEUBx
h+FD/ClKnnnKd6kBrRkcHUfVK/qTRtohq8fbZcCZyckU5EPt+gbzzwQwSmCjgAZ87keynForSEg8
Uba88PsPblq2p/vRt7SkMwsvsPKy3NtRXGyUMGdDHGt9/nnxtj507XRd6JybmiSU2rN0Mdq5FYeV
qyXWGMYWLx5mAczXH96Zyb7nTzrM4Oe55SF3+K1rW3FCropwekmkCUBCw7KdI7IRaZ6NCNbwTGgJ
Dj7MpLgyo32EuFpaVAbSdI6c5Zb2SqJ9Z/fhAvFPubbQ2gvkonEcolTOxwpiSFcYDJsI8gbJWLHC
/tY2zrn0/3lGHqdbGg3tuAjdWScnjUN6bfdl3VItoZJUpGHY+MXg1uqKJf6XCJZg7SbtlgEdoLpf
zocZOaZw2ZFoScJuzO3OKIbq9PxSjFIIDF6Sfc0qf/M0/Ws8uKHOamMHXmXknC6iBZMeNxpt8aaR
5wQqb8vxa72yx0l0waFb1wJ4F/eCP5qMSHzr1cYRTE4vuz97ffzPKbXEMk6VlWA3ZFTAnEyB2Lvj
58vMPjIlIt5MpXvQYUBVc7yZI09ZApLQD53Bde6a9vcsX63PUf+bDDFt3NAZmRtOwddtYHkgpKzF
Le7RGrvlppCLDRbmVreJE4C4jOVCN7imz6Qdwf4B32gSmHJUFzsJ/xu4VPPqAFI3/nhYlxW1b27D
cEvc6TckB9KaP72Q8QPRM80lLt5cn2A2xK1RVAUE95BmCF3BNBldaPcjJg8CKR7kKEAj//RGgQB2
m4XDoh7fc2H6oFsbAMT00G/8GNEKtLbT0wvcqoNH44O2TGSaWkl7SNZ+r5dk0p4wrI2m9nPkM7DI
/0z6jPPFuo1rZD8heCLQvqOG16MwlXTjU6qLDdkCpbkzemQMlRNV6q4Pdyu8GhAQg0ouUIRhGbVu
Ny8ZvGAX9PtpDp/kHejkMn64DwoNMFS9hfWKBAT0VLuxDghVofDVo/nVO9Tdnt1kUFTAV0ijXgh8
6gewF6KCm1WidC89Au1kw0oIz71iAEcAQ/1j/ocGOl8ToWLgpr/Nfzup6Xn7l6qmznyAAUgfLYp1
c+qOl5CnFFdDM5SvELz3NkfuTbQHZL3l5HMr9wU3+2xnKRtE37cjHueGIzmjbeR59pUzN9/680N1
+BLWe2IqrYA70RUzd/MVSWUcn5RTuiJhF8mGz/N4CZjpagaDBQbOk4y26QuQCbbHZckoLgpYXztC
djRD8vvt1cVMubUlyD8ucbc4KoLlMhYfT90vKWyplCt4t8kdKmUGuJ1Chcw6J5bsH+tpDcem+h6b
beYoS2wZFw1mTCwqqikwMb/ozjyCUX3vBsX/4mBl+9sO9EQ1XJjgg+wn4aZqkY/4KQldXkYTqJ7Q
tAQe9pghBeznjTuzyynyFJXEHSPRsJvOok4uxS+/WKDv0mtb1TdzmXvzhcCnGp80W7iYW+wROR2c
5yPei6/8QmlocNz2curYgLNanWKVWkVjujb9YG4J7lclvhqJYFxbTpS0wTx+KSsrN9eUYAavJCeq
DujcbKYYB88y275SPjN7HYmVC9LTrAEPOTRYAm5eoj3sAyY1r9ri9oLFzBarRgY4kEwdDXBaAgr1
g0FeJbLEYjf8xgQqyaad/7c7P6M3MD03f9fr1Tk4O+3cS76+A1qrd2QpN6+Fg2tgY5X0wY7UKfLw
JQBh3AJ20PxWDe5+vzSU41GYTvOnzUd5egjNuqWCAQXeIRCCnVEolHge/kOs/osVnXpJ0ZVDvgyX
Z5rH7OUVI2qhan4ZfIxFEnaGfUNefCOPR4xXyDu7aE01p1HwEYOJpN9I4vnCKQEM/CKUeVEhRa24
TY2voAXsFBYlK2yyKt6v2EOLvNHgd5M2sMQSCB6cnlEyuLiTyoSQMQrhNAHL63XMw6Cpeyh+LcWB
K+ydKkUS9yjO5EEBbYmnIsGPZhLjtbLrgLqsdcotvYpbpMff8Q+FsdXVQVYut5QWH/ZGEsBDWUeM
ZeAQOG+M3BsadKjZCx6bE6XUiI5tfTbeI9wDl+z4qvlexbFnU9DUAbyRHCBk/w+87FLR84V9utw3
FNdJlERzi2W8k4hI7ntQz0OGW6IndIAfk6PhhQ5bwdzCfQour06u99pMu9sQC2WwPU2k21pSCat0
XSU8f9/LhgPJxdWUXdLGlJg2KJDg5Q3u6CA41SfIjZXZJnOg4i+2dkPrqb52mJdNLCG4zy00teOB
PVva9+3UrBe9W5+TIFFOH4mE109e+UKq7hszAblXacrzCCUkF1L7SxYP8IhEHAc/R9VSnoWKsYL3
TwfXZ7hq+VUqFf+C+pQrIuARgpqOj7t0rim1MbngSyDsfVf0xcwF/uUmONBzNUnYx/XSeWXPapVt
tpmFH/DGv9gVKq++/2QeuoChc6mo5aogIcoJRuCzIxxv0JV3cqsjDtHKxxJSvWlmizOrJrIjwOWd
NZ9dJJu98olLiy7/JN8M+pHeJsEnFJ5FIzmSH8ln4cYrNExp6MB5QLPRLM4PqJCtpEQ2NASkjmSl
glDc0K/ZbM2pcV+p6kmur1RrLQ3FH8Yrsd7bYo6mz1Fbdo/YvjlCxEBrR9SwniWUFunBH2MzYaMW
tZA+xSmssZUChqpKPRVJOMYlN0Wnvt2TQ474bzvrA26siX2PcLq4fzLi4EYPO9vtQtK5QKspw/Z+
kjI8qbhHk8DrWdVZFS4seOcQDEAd+d06IX3zb7qZFzxTtsifWLT2tzdeujK98yeNBKDzyTyFHLjW
iXO7L+yCCRCxf/PYPk9eyN/kcesLSawlJ/Rj8tZZhaxzLGKrn9u5zJ3V3RDrfkun5kMhX6oAgksT
MC7T92/+bUpO62fLhQ/euIEzm1oq56bu8jr7YU8AXSg3+PBDMT4oy0WIuA0+Y104zuPSsWduCK1w
C/f9go1a9Vk6c9rfsBTECbw+YrOxdgBE3lz3uZcToLdcGYeFkWK0uwDj/YKt38PFJXuqHsTyys5a
WP3Psc/d3sC701oCWDbNbVuku0LVbkBvwc0gbNwJdedsD82mG4gJKvL55QGGn50dhu/zUDlUAfzl
mzNK8hKXe2/ifG0w6GFf0waQmtaDYAzJmGWkMYIUFSTLVrifeLjPEz6U8vGXIdw1lBkIKQvPZB1j
7+EN4zAXbdGIM3QcH6amAB+OGl0mMktCWOJNpAi93pF2cjeKeipjlTqp/pRHMIkGdLtPlEs9UcuT
KqFb81tYIePsCeuLsdR+a7a5L418mFx2KnEgSULSh5RQJL/wZfXeIfvMd7A7TqMD4hW21ELhrfIC
gfHE+yL6ZOfyp6hqc0yzrAk0ZwP/K0uJpyONmPjG8GTAdaCXjYCXmubV/l0iX3XoeBrnh5EaNMJu
cVTXqZmPaJVm9d1npl1aKIj9zr1GGQ32PnZDLXA9mxz5axDN3+0IZFJzbPaBYypd50iQZnYovwAC
QeRmXNy0QYE+jfvkQ7Zv1Hv/oJDkvOsuck7vXBUdTFEToe7BUlNUi4vm5pXbdcqLvcLXTr+D7TEl
2ie5jUZCYDHN6nQfn7yz1mV3VeC118b6nv84/C2+jdHfSYDjVklvvYXnI361k3sygQsgHQeI9OU9
m+r/j8PXNx49g9mHMw8+Vi1H9iDXDUsjhwOT57DMvUJMXQ0q4qToxIfzrRgTbmxYlZOAStBghSvC
Z//WAQcaQkqZhtZBNE7jCs7FjhZ7uUZvM3L6Fug21g0mU031NvGMxIoG9eWu8rVWVQRGNq6eflMQ
pITyXit7GS6nHRF1xFZ4igM4W5xrEUvWtu0TzbelzSX91yk+VB1EvQnaMK/gz4uMu0xrQ3AZJcQF
btBo2J7XwHwF5VhaVII7oWWxhlQ7a8BPb/cclFRa2VBZnr1j1OTpxSdgHok0ZBNNnuQnrNFrtLKg
D6uxJFIdNZi42gBivOLZpnzqzprcWfI9WPp7elyjyeRPSSEe7WpoIBmoy7hYKyPT8HMNUhpQr4Pr
EIj4f6tPMK4mWn7/ZANnwollBkCETjAJcATIF5dOiiCloBlMkG8KX5mg7lnoJta6wDptE0MSWbAo
JgM3Ga/uUBmKwkZWSkR+n7ezqVVJhFtM/AmGlIYmEMTv2v/0nGcmQXU8UzOnTi5J8lG0JWQXLaM0
yqz0jpuuwkVBgO2au10DH4Ylsu1JhExkYaMkiBCrB9vi0wDUKNhnO72ZqAkncjrZs62klOoMlpBh
sTWLFTd3GA9HNRmHrv/+Tge1pH3FeE/DalVrY61Bcve5gdWT9JBB9DDab7GkzzxDYI+oY+g7O8Yr
Ol7Dd8JoZIT9jslz7FihvVOXH4/tawhXQzH728cVZQPHRl3IwX4pNyZXvIduymzLUJYD2vGZZRrF
NYKQemZzoAhNdgO/pTG2IufF77wioJgH3CiqZ76sU+OVWG2vtYeypVXIU7944oCXk2VKQvMrz/CY
tXIDD0hxvuCaic1251iNrhU6MeQiq7AD5bItAcW3nLyoIEIU44wlEe0SoVjgsp47IbpTLOEiMwhS
MIqd6DNv5sc9RIohRvVmnST7vT+ShaPuodKFrijRu8D3f+KXgQ962k2NXmiTQXFD1qhFVfzvc1xe
KQzBbqb4vIAGn3x5rZ4+Z/sHUOpLNj+T8Eftp63SM3fGuxN3/h/AIzcZVjsx3ZG2GWXMMGpUdC8D
8XSNIVn1eygrsXOdRxJJcbMYaktW8PjbU8SGEEMRAXXNdGlDaaWj26OGpwB/PqC91mbIoKiKF7IO
NiV9kBPF7GU+DKC1Gma2NsKHyj1I+ORNBn8Z6s4m28yEfjUVOMvZJuCptxyi3ZEtt8aYEu/0nCeX
PZdgjamlKiJ4xJ6rIvBziYToAWPwyle/mMFWTdUP331SN79k2eKlmiGi2aqyDTcQyQ3Yu80OmTff
OUaECXGwch/QuhoRjiGy5Bnfljm5JNqbUrwxgZB+J689KCWEG9VsRGkaoMaL70z68kwfTw29BGL/
bvipeq2AANhxAAk6ABrM0CumLdAVYgpHSkpzykiYEcX0F4OEP+qybLXXuRKIivIT4A3B1vRMowFq
tD4me9Jgc13u06PUGKQC0U4Tcqx3fDJBfrVqfKPjT1sKRq09aGyFXV3my+aEuCjtR31FuNMZ/G01
Ur7d9nhMN3JkWPRxYJotKUx3pyOyVeTFgGNHtf/LOZU+rB2QWwdjfK81Hl1i3884XX/3gkNOkbFV
ZwNNdmyYJJCTIIMJLJmQJbauAerzKiUQ4OBmDBoGCOH2olXmotTq/cWzpIHrxPxbWh6G3XFuZwDm
JqHIowncTmPDuST11kJIWLGwlYXALwC+IQ19cZfrh4dZBw3WOzmILiMfZR2pB8IM0g0mdQX1e7w0
8MqgLThIzcXO3c/i7DTVKt0m/5Myq2lymF0rDOOUDmMFHgQfzoyRpJgYbId7qPq5HB2A4K/sKpjk
Lu47J6XfNUBL+Bi8X9+mG4tqGrrpDrPht9HMbrOr/+3snN4vDVeZ9/QipT0+TI8qgXEuQN7IrHuq
DJwhuWEAWCfQ+ThDWl5GrqYQ1pQ5Y3uWiU+wCLAo0VlnLNQ+OaebnwVkXqZnlJHo4OQvGcOcfva8
8nwZgWaAIwlZbJg70TVFM8elkAMz+XU0SIobqmZaCYf7WiMBBvfm0eS7trne9OVLbYR9Ky6gVOhR
38wSWWDxABj6AyaniZSsckvsPe+aLioApbYS6mo9tJyhXbwarU41evT5LGsjLrv/YvOuv9M1tjd2
95lODC1DFegS4BoGGMN99L9L4m/rTIH+Zu0KcZhBcUoe556bl9L0YQDJRc5YzE7OfIplyWa7lr6c
q3SfUnZuVhwly0iBOObE0WaIpXpgAznkFnNqhgcjG3tsBwdBnsDnraqWig4/HUKuX1wVWysKVo4f
7pvJDTPTclUrURn5SnFBg7hb2/O1LcsRylSF5+KggermXC16+0b2dBpBKmUdaQNUMt5sCqFAQ6zk
25oS+QW4c6GP3GR6yKtraH5Kfa/58jrT9M1k1BATkWmsw5FGJ9AUFFon/PTFHZngMBhSHnAFfzpY
fhoL9bZdO0wgI4oqlw/Pc5MzL/yNgf+9rEwM3I3IgDAyhbSqkGOpZvr80/sgaixQj5db5LvQg8B7
83IJxLiI2UJ54DKagWD4TjIlfdLu1c4PdGk7FDwKuWtPn8VUq79cwlXAQcTcYJSf/H6OOOHYUWzY
zws8vQfjU9PaYN1igjQjooVBzKBbUCdA8J0+A2K8bBH3DUsKgv5vZaPV7bIPVvY+3ofkP2QytTsL
Ie2ibs9LZ12WA+KKr0YFhIt42IglzyO+jK8W8F5Ujb/wrm5w/gu9gtdLN0bBIXnRCI4Q52lGZVl6
B9lSq3kn2qzSn9Rqc9ZVCPSo4vgmC71Pxi5FwvPUCKx92Hq7qgzBKN2qPclAS4xSMrdz11hnx50e
cpKCXivr2CCjlXgtWrp4hPtMSFL2L5juBpesJ4ON+XT9XORfodAMEszB0vOT1TI3fQ73uu/4IPtp
bB6d8izC/GRer4jWbv5zuxxhMvNWN8tw2Wf3MFak+01ed38rT3ZmolZsmVQhbTbK+BH7LBumAPF/
2aw2HmebM9swMiiVgaCF1AmjN6mYLCZTADdD681QYSDC2CkY47emaMW3VbJCqnXC9x5oR2jpBsjE
pwQ4MtQ9MRuA7trSC66mn3MUBeEVmg0FfT8Obq/PgroXCRG+Eg7o5ZQPDFCC3TQiCCap07SovQW/
I0QaOFN4kCDwYUgOl6XJCifscYxGhEmsktQxXpOKlWNpdM8PoXqVDz8qEL7aGp/6wb0yjoIb51oa
FlMLNd+OOJ9brycJEQa5XjQk1iZ0o1VYTCblkgHfjJ/dx1UefmvyHdXrSfZ/OcDfdgq+ZN0HKWEH
PtwhGQMbdX/1HnGdlGA/+4ZgGe+vh6sTQi4pjla5IFcWb09tEpSlqYgcT3YQAAfaZHyolCH1jtui
O+72sw8GqiVFqpBtrvny4i7TdtUha3h83Q/wE3oQWCienrMdVVMtVB7y4SsSNas172fyWY3tnfYV
rlpaBI1u27iLK8tV1NjmvQtGZUXBK96gv7cxk+ktkAZLw7My20McxXLVnRj7lAOaAahSshpgYl10
Pj40697H6RNBlZQuwT9HTwHobnqU/kks4wD7n0O8IecGasv7N8epYf53DLZBD27JsuQN2ojcbkwT
d8jM/rdEHH7MwDz2h/QdCun/WcnrmPZCJM2zRLUrQ4JWBqIxDsEdICUYxBajKryY7AW4gjG8wgH4
kdmQi+yDp7qCnVknC4IFNuljwJSzK8EhcXFeCiriZBYVb3t9spt2pG3YXoEospA+hLxPym8/ugAy
uhi6fHcbYe8GkXY2PuzMwt3FmJEcB13HSl/tP2rkpL+sAOFst3hl41pw0CgBy+BoOmirjtg8Kjcx
0ToeGf15Srtc0/YZ0oAoEWaj6r6sxEK0gXu0bNEpKs35Syj3rq1nWti+8x3t6EQQ3ZjZm5u50p0+
7+bHFtrpjwRUPjCzYDqpDkBoeEQ1T+4BykEuP16MHD2IhroqOh//bxDXC5WgqkC+M4cBR+3oB2IV
QpCu1NitVoQcjhgiGSmisHCrN7cYq4Wei6Sf5kcHTxLJS+SXJwyqWobavdYWwzz4fnL1MzH995uP
TGS9VQDi4UhaXQhHqRaPh6MKjOsnMO9ifMe/pQtendIzWC+1uSkh7NIyB9rUIgPw6lgzQWEVfcN/
cLPCubhDdRwYf4NpBk9mcCRhsoLLGXqOKrSBg2x3/H5PvJEaPSjSozuqLBqASRom+g/iGM1UsLuZ
aaR/3+Xi3V18N21633XEgFBqtkc8wwYsvhUnT75nxvDwUZ4yNWyQ4WisMnBfAxFOhQlpTGuewDVn
+sK4CO1IQAIgMq4nUEb00uD//zdZqbD4AZL2D12xhcSeprQ8+R0A8grLidgCms0+R6zezx87F6Ox
GXkaeEtvdKwPk9iE3WSZIxpCiKQp9p7+1B4EZk9/edIoVfFwdv0UnuIx9KfhtOVu24NlYAh9zqj1
izyYhMxTL7bKnK6Ke2s/N6VGmj8np1Bdyzl8Biphc3S20aAlk+x4InKSOJDTU2Zl3riVuQyWdiJT
kY22MT4kaTZxZR2VYZD50UxKPMlQn5j76s4z5X9Cqxewd+GX/TY8WqdVT1rt0r9dRT4IVrpE3Vyl
DQCagRfOjDddut0DOOoZlVuKXNHOHajDC4icd0k2QEB0LyToLmlB83A9WWwC2ELqZpvkantbmKq8
rpCmIDwOdUfUCveHTh/Da0Hr9l/35PhpvdEtirhGXyYP5aOvrDe9jDrCbssgEnGn+yDcdG/GO1Sa
FJVWcwxA7uoVGbvfQI0L/05aeQcB0VDsdI984laclqyP/sejm5+9ohpIxAFS40Gmbg8+rFGxcC1B
AdC4GYjNWDFu2XtZiCQlGurqz2bK+ZeBgs38hYutv/+354lqHlmwVRmRqMygzjzMkUfO3WAA1gsK
ox/O3movLsOa78hK9QbbF+ldmzhe6r3Qz1SLIAA1R6JDV9KqA4Ieab3YOSH2UO3SjwWQG8/gfiC7
Y2rQDDoHiglafVsel8wFtmNFTUEGOma1j+QTHWg6Ax194Ga3dXLCQtNyamWwgmmDPsxQKayYiJXc
U0+6ToPYgzA4In/t+A9VIfofaj822QVCl6DbFs/cInPVff62CuL8c5C+FOHUOJ/wGtmNXlTOlfEB
wqZPeVmiYIaxp/DGy3sS9ISILJZXsTJG8IXt6187dA7FR0zCGnqbMCmVhazpQOEfercS+f7zhf1b
fnP/UvXTvGyz8QfpRTXTvIqc3h6vcSvmT8WS8OrWYpoddx+twnZk/1liDNUabdcRxAeJKFWI8umB
dW7GyiC7IVvLAc8kE6fJGZblhMwe6OqPifZ/H0OXTrRT9sc1vkKJowlL83k+2eyH3qwi01Z7EpHy
izVIPRbJKg9oDrW/sjXdln0LSeWrPVuOavISA3/hTaCDv09yL40y/SEld8KrrjjaxBameI9Ywxdc
TMerh9dRaq4deRFNhNifMGZcnP1baTQtYn/ijufomHdn0paV47ceYGGvzVt5Q95XwePwT9hg7jtx
bqEfbynXApO4Q10cM93uF33zoFvWgLEHULqXGCa2RxX0iSQDPNL+UzHSUYqXy4/hT1+zj5NYvzok
UCY/anBlqiQFdF3M34df2GZwcf5htjOlp0vttEOC6cyynUPWJPf7gk5asAKpI8LoRjfSS9kzg+3u
5oRQ6TgkzYN+eP3RLGRd2zgz8Ry7Qi5n4X57XvYl5JixBF5kMZROz4epNf4xAvNeMJG20DBIbP2P
3a3s3NxMB4rzfY8+cIqK+FrabttIoUsSJjMTgU6cRzJhfoPAKIcAJtvBVqbODcKvsCxdc1eL/fis
YLj0Mg2vWBsbaFWV8v3PGu6Fo7aS7BLa1++0MHBJyHyH1SZ9RH6KE4gd8n1YE7+bSDC0FIKz2QN3
8UTCXMY7OJbsEJumg0GDZ5qQPZ0JdhFs3ZUy1ApHgxXOBQyDNjDyDZFZtKU9UE5bzZsKXTN61AhA
RkAAHsaTXl+9+jMSUUr2SatdnJzUyDHdZy0e0vgR+upKy4DMYxNRfUbBlzTew62C49NhBL9d4sFA
otsANbTh4EPnfuWM79WmvBrPboMnIFmHk8yEYQusdEXvNhu7GYCkVm9G07H8hRl2jMRrsgBYi5vo
ck/G1qZN8xW+8hfYFyHhIruZa/xyzoSoygqgABSlJvXG+/bkUwXa8vkPdL/LPxjP0swmwUT9yeYw
MbhEk9lnkD2Lg66VcdTbLi/UdQTdcsTKUBe/HvXuQ/ghvEYC26I2unCF4mLZyiRIKMEhOcXnXoIR
81zg5Y+EURtGPtnI7mY7EBNTJyQ5UvYsri+uBlGNyDUGM3uihYHjjI0zdhGVZomgbbIXXjkBVZWJ
FyWZzX7orOTOO/oCn90ZE+9opaptrBr9GY1BSdBu4OGmUGbSanR0sJL56sm0dC8FY5wR/+8kP30t
2nt5y+FZVUy/6YLd+VhqLoAkopMtRY71RFPGNtPy6nATjIvjSeima0WtHwtPjfTg9AhW40ICLKCT
kgV5JaRw9gScDcrKJBlXznmaLw6EJI+ALOdMwXA3622zi69IcSFtgkCW/VUxX1YUsRnrWOgR6NAe
iM0/yjlMJLWhNKuHLm3lmjP13PaAw7e9HBPdoj6nbBzSr67eDKQAFxkt8mAM3OWOBuP12XMFpsRd
SjUcbqxgYMFk2Wl/Pecmc32GnhWubtWY+C6nVUKyNKaM+RLUtQS5CCSbdkgU4YuFZV90DsjdAdPU
JK+BoYT3I6oUR866OTd7KiPDP6vSlGvVIrHiU9qJFNOu0hs97MJOkxYxfr83bquAwmoQA/YImBTC
VqzpWCRhZ7OiB0A6l3+Ggg0mAWAdjGau5YhDVCnh9aXxJb+RnbW3W0fPZNEajWyfnYNiCcCDUkqL
hCUow4uc3VLaoycEUFeAKs42hAinbgc58S9kQWCW9EQOJHJtLN8UMI4MuW3tgUjxu9TrLuWhoH9D
EymW9maaBlyLNZNc8PyhDA1S1QQSJKCBxJb/9qsMX4eWJAtbreGFeIFtNdvxCq/3IW4sZm0BP8Q7
Itaw90ipk8Srq9ObSN3MRyV/hgWEwOoDHeNV8e6eYN1v6XU6r9DH3RjkjmUetcmcoYAQkoDUsFtw
DS6MAad54cGqlEcpphMOAwlCPUZ7lgGOoY0QaGc/5ANJHKYcllNs6PPXIT2pnrUK956lc1iZmPqx
CQ5hxj29oX0fuRrbozPhE42CKZBV3CnXSJCotBY3ladTSDFcPMkGOiCPDHkGljnas1nb0CA9j84m
HXsktxU/TiC+6G4X42RDoMcG/W8s44QLSdFYfXjjwt7ifnXfssiGPb81ofiqJCjW36vpi4ajce30
dpyNSRh5in+sKMxaLpL2dZtcYSQunlX8BlkA7tiEzZPt7+RrqZzlNQ3ZiIvUaK8yrechHauqVxtG
GCP6rlqlXUPjk4uyh5BCIN8xeCFzRaX6wQSyqtZIwZWyE2hIEtZg+BbTwapOk8+LQZpwFyoqRVH6
kyhth5pVRg/nBqCsmoQ3IT2q62InNEzgsF/qD4LBqLMCHbdZQjE6BrDUMkEsRM7yB5ma+xsNbds1
lvLwTwx4wD927JaCTRWkB69hOatdHvAS44ihtMNRn843dc1JXT7+1htjXrX3I1ZjeUJGf9AtiuCa
IuvNJQj94bHsZxWDABYMeTcfClZEZqKkYAzmsCfoeiEHmK3JYbkUlVZECBPNexu+q74lmLsCP/8t
Vcnt+6n4M4gk7nRJtyNFns1PrhSsnekSYPkjylHdRGSxikWvTcVixcM/51rodIB2bY8Lbt/I9VRt
kVhf0p5O1KvsvKlZCcPZgnhhREY0dJTMkOhUBAl1PSJzjZ7rixTXNKVLAnGEG9GoXfc8T8AmkSfv
2fQOVyJMQKIyqxJdY+wA/H5XfhgkpTh/WOZYbThhOY281aoIAse8kyaIAQkfYsdcQhTQwKdhWkJ6
ggoGH6Clbhi+z03ZP0RFZM6e0gU4owfeZ4JiyN4/53eM4eJTmRstf5nh5/cUdvlJS7HHRo89P1+m
3oMLT4FbKBENXbqp5Y8GvWblDbsimKG6UpeFQHexGcZ2bF93U5CsM/5v5HPEHLbspRD5fV0VQzDf
x7OulEIVf6i+7Ch9Exqn3u72+zeikWDapPLLVabK6C2AXhcwjqLXs2bUoWG1jJ0Vh1+P1nMFWJIC
rzQexr0KSF60GveOcpcunORxAbz8CA84ksemR2ipM5m97Gv2YIzg2+Xj9hw5OcU6Bn9sj+z9KYDO
F9yJHYrGiBFlSVbcDgKwJhNNZbaRoS42OteHN1PLjc1TpjoHXjNwXEMMkaBJz3QffhCVuZqNBH2j
gHkZ7JD2HlBPuvWSDsjEjEr2JCelvOUQ3rxaqZKhgyg6jCvao6shkR3GAPN4Kq9kOGmZ76oD206r
uY3kmbR3IMlWsq+l7RO8HSn60DKicGeYJue29paICpXk4s6011BT4H3JQlMlRUkQ8D1x3CBvZjbd
Ccs4057+/GBrd14vp+CDvVuA6I4SxFDomKvnCSR/ChfjFa9YLg8AMOkizYVq2+8qss+OYJ/RfTTn
tCItLYZgKJHGO9vKwm5F4xVvalT29OGKYYbvQ9JTljggapL2AxWXfp8jCsoIZ8/bJEffxfSe96Ag
uGD8hdnaqSRhZfENhU+8oRLTUFEai5t4gNre79vbNBMir8NdfadTqadSBd92f8N0G1lpzLJVecih
wUkTae1y+6Gq/PZ6UTnbjQd6OLGHj6drAxeifrSfwEoQUEloEABhN+l3sA4iMRHrDfD05ghXQTHF
AQzTTjfBJYIKJ2NhZhJq7a5oaE74F1NfZZrzP6syt7DMeEit0JT3k32tpAwvhhDifQxjbC2v47Yv
TRbYpfch3i73AFgmUWOU+IduHFaFITXD4wd5K/BzZVWy+AkQXA43KcUQl1vyToVlygdL3HIxaTcz
1q1DXj4Urtv/2zU/LYV9mKRL78tEZC6M8COAT5oA7pJ+wqRJQv1E48SqHls51HDUP40+DHclk8Ad
U9UsZNfLYfwruWOf7rSMzLp7S0a/mNjm6WkDCeCkK8FYbfArnExX63ciLgFqTIISGvxYal0Klli7
m0v9K00LMIlNb6WQmPPuoS5iFkkg+68yn02x5DY2w5wCOgkOrC1vDwjqRfAPkdgn+grU2AIAUtK4
V+XF4ZKJ86yKaFtwL4ldY5J4JhcAFBx6hTVBr+Z2iBav6Q0ZR25fiwXwK1zIQECWB/Y+iY4dCw5Q
LfGq+4YGjKmf4xwwLhh3WOPoXRMXDiXVCx3cDzOJSjcHW6O9nIwVuGK8a1eHYDxoTaJ+wLb8dXqM
1luzv7e2RRVo+u5zT7JP+3cFg+tFEdh0UHbOcMnLkEyN9ie86sQEK/kjaTL0MnQjPgsaz/ReMZ6l
BUkk6SR7foE/zRbPSY3w+NCnRnyXw6yFXjIPYwEvrJK6U85zbySo1T067E0DnGnKMmOcwlCyIvC/
IPS48bxTtJ9DBIynrP9JA4biTWcN8kSvv2VQo7giBiUpwpmNaD+otG1gHcmh5aMkj0GKk13U+108
LJ/BnS2+GJl5AdgvL6s/oVw6cfyToqj/N6SDLnXbU8HvjLIc1tswL9mDXPfFuolJYZXNIQWuAdDW
94yCvaCMsR3XkcWjlose5VGh9NdC3lrePg0AhA7AAiE7OtZ1jtymeA2iHzOd3rKGqSHukvngGEMR
hXANbCLrgoeHGD3o82Fta6hV35MMh1kab89Igqjdj4Urb7VlZ2CXpU3Haef23uWrR/vATB8SgqyX
QsqtvMPhK8TtnuAEK7YRwxRiNjFB0nLAyi+r+7k3S08HVXrm4SvwxI2IDwgZBOWPKx5sMFnnHKmY
632BcLPgrH6o+DoRUMhb4GFGPA7F3v1x6BKGBzDqhgxG9uA8ZabhOh/90p2pCwFUQht1DzqIrd+Q
0Ib50vQfmX86f3vOIWWAfHEsE3u/gfPGSAJm9CsWRHCDciJlUXwZW0jZMCm95aGwxVo1fMg5wB6C
nbj8wgZAaqZE/zutpV2r381wLX4CIH194IMMnKqoOKvNX++Uyjh7JoxD3p3RklpBc2fv//tbNz4I
FIfaEl4ESaEBp8xmP4unpL5Cqu83QNiHXHtLKTfTUXLAnrNdjrM6TzMfnxo1Di4AGxSNts0JgWnx
QjeGnZBHPI1HgnvTxS6qER+V/WDw2VgWm/aJuSFrqKXkYs/E0IEx0EIcJpoppyMj9fppc28g+Nom
JDQPs70YzwjZdhAzRC36pIlgTm+5Wi5RzkZa7M3OSQT1H/31gqs5ndl4wqN9ea+G3AYmzV0H9OT9
6WS8S9Mu68lpeSYwlq0Dr0czgpUv0dzgpuQC0NS63OKMQ97LDyzMt88ljmgQIIlIsY9EozmD2DB/
kOx93Fal7DW/V/AXP5qycO5BdlWgUOoivfP1CjuLW/WFOH68UcesrlvrKvEiuasSpscJAezeRrzI
1IDGEaLJHnGgYzqBMibJEVudTXvwVdyr6IUltWV/wt65l+HQ9akOKhreEnuQcZ2JCVEpf6l02+K6
crG+X4L9BvM+VEm1p3eFVzG3qEi6VyUqMgYUauAGe96M2QMfUnznkUfs4/CvnJs1ygAxlLQG9CCW
3c+UTSonXyO6YrceDWbjrpS1mxXl+QTRXZRul8nuqlFVW0+WPuaAD5EtAzPcIBzjiuLa2lt6BkQj
avtf2ZlIbmBF17cbmOoaJGIAZfLcgtQcxXWr9y7vqN51iwn6687pLkhHR4jmSihK6vHGFFlml3ev
+VxxeOkDZLGAv2DVzikMTQft/wCHq5QF37e92dzjnkkn4Y/HxwYiDw4Vt+EDEr5RnTimaEkaC30K
CP4K0CkK1jtQ3C7svXPqt4QoWiYJd2XU5kFAirTK7OwgQJMqogGXa0Zu1wz4u8gUXaY7rbvuNOLz
Pd6T6glRHQ8X+5EFbelUW5j7z0H/asvJ5dZVarFKl8Ho5s5M8ToPHrOf6tF+MxSIRQtDjI2rmQkr
IatBBbMoxlj53pj8+0BH3DWowY5mS831ZZvFTLU3BaViN9Dr6Xj4G9oeNZRTueMWX7qtwIjgvcwl
45VoiSVlad4ewYVZZT+X+YGgr9+NOkLKKk4LY0FzoiKCJnbitLpd6zeL5amdjNtBKRsYm373nu/Y
Z6/Rp4ulB1cHwYwJii4fVS0JVW5solYh46g45czbMVeZnHLKCuwO88I/bbpWVoJLGTr9x888Yzo8
IlqgZ48yJlbJUOqIuscYPCnZdkkX9QBcXNo05/Xrf/Jk/cvrlOWeJdFbw1PX0AkFf6zTdgoDZgtq
a0TIN1E3zucxtxioKZ6xA7tj2dYPd2DY8rQxH4AYMKh+PWKiLsI0U4G1avybjkvLqt4YkKkcu0IB
Nk+EpGOfuh9PZSF8QGNrjhzK6gqKJ0N+D53WBHwYSlCVPk3/oNg+x7Kkfmyz30f6B6jzfCs+45YU
JrW7CVtqZVEuYsstBhWZF3QbOklfbOb0VsPVW8LV5O59WVsQWdZlGA7llbwN9qvzFhvbCKf+paFs
iB0WJ1UaYF6fa7I5YqfuCJTpSfqFoDj0WbQEh+68ekUB+Qt96RWbghG4ljgQ2LZE8C7iQPGEo/yw
m7BTnBuTV8xHCo+mTRoM2IX4Fpln6YtPJJ+x5t/XJIwWtpYlYQnLbj5cZxBUD6oXzf+g5WKaH+u5
7nm/+ytJPnibGs+J+ulN5Pu0em4pymIPaarnjxQk6DkCkuXI6Vj/YgI0lM6UpNnfbwRpxwOfaegU
lgVGrrZs4k9jbr2nEORfrISXZa0Bq3DxxqisONxBKKRcKnqsEgM6razC5c4B+9s8HWwQdIZhHDCi
7of64/+YFl2V7eZZMiZnrDiAnk7AMWieTehzx81D7Uc0z5qlgfKu7j0YCjii5I481DqjE6jcSw/l
SuOW7JcTLsN+4efCksA5072Lqe7xssBG9EfPJHexCHCzmv25CAkBFYmTyarQeHbgF2xFokLqFtkx
JOo5pXON1C07z6w40Bn0T2rgU+saMG4z+AzzRiMBa9g2Fd7d/XkcGyFgDMm2EsAi2kNdpofmCl4O
aB4l6mGzeWNuvispiCtOLlV5lr8gXYW4EizXdbcIJU2cTJ+H39DlROP8JvtZz8IKsnUSl9B5OvKC
/cwfvAOMtGeEWJE6Qcl9M1OAc5F7FnKWE+pLSKNMMLAUB5UifX31II+KYAKejZyC9UXdF/ZCuJeh
iGlmk9mioUYwRPxFOQGAt2nN+/08vpXOtFeabakSwqYkmOzMMYXgj/cGahSbPj2ypp0Aye1hECoA
eZc75rh+I1osu/KkQspFcUW82cnATfYOORAL+kJDHmEDBTbvEe6KKVPHC4Vq5NG/J+Gz0yLMo//W
5rSnnaaI14MW582Y77kspgMlFIka6V3V+q587EX0rm6pJyzq45hrLXzX/8lWWuVyOeBy9aOjYzd4
IZkqhheyikeQNIJREi5FMNr46yG6DFHE70X2rRGQOBXnXjjx11eDSir5D72E2noJTv61Z4N+n97O
wsxx4iimMLrlloojAkSs3YHo5CG2Ih22DJ2AgAEzBt8uVrP5T0h5vYpPVy5cbjUbcVlmH+7k+yBu
0FIeVAgbRgyGdTZLZ53xvfK5UuCtet9UgZafPMmwaq4u36w0hn83yMmbkZAMGsq0woOHQNr8Wv44
4QG/7z1aPMpkg9/SbS/iXFzqXyTESYQoLwur/NdKn4TXJNQ+zViJ5BQE9mAuN4BeOYRooYBoE41a
gUe1PTueCUSsLFKCh5IVnCSK7TAHiZQo9ZN2AZpOZIk4nt+N5DuYTD22PMkkSEze525xVQ+AnEi1
1tDPOBGAC2e4n6OhnBdNkp4B6GOXzdoZM0TDaAxTM6V1Bknr2KZpBYcvP2ZPzGtMUvxrxKCeSEk/
4twFXqjV6HZJ0Hb0LAyF8JWxxdAJwRPFRre/fUfVLr+cFOu84t2y4bgl95/lHks+NU0jtc2TkUmV
ngs+R5/xjwi94T6Z55Go4ZmP3I0vuta+FGw/kcBuBDfxDW1RkE0eGFwsnHxStuTogww+Q7FN3md/
2zTeadtJRRriBCUpEQ4HmzLphkkXMLWfnthOqbmkAPTUTqwSkxsXpBBs8VRYL2YI5Bx020+Trwyt
0jkdFGI0IF7vjzmHuu3MDJwL8btXD8xluJVs/KDb1llXFPdcZG/vAh13bqhp7spIS5oXSaHXx6nb
e9vlAnEVUE5+devAXCalgxwjaXlWiMPTZzvVWM7DtzkeR50VRHnEw03SikSRYH4ak+PdiBk/+bJn
N5KdmIeL5Cg3NXw15hvIa4KbjaYqkIkg0yqnAGIVoEXBQOJzJh4ORIGfe72dWtmxW5G6LO4IUec5
V6MU5ifbCah2y4adMx4+mEYKDDkq3GR2WlOVkpAkVw2bNHGWLNqPMioeh+WeDc1FPD7l4hK+BqCP
SLDpbl1Y28AsFZTMgUcNfIjkJuTSgtXFeF0G0PZpmQ0Vqp1b2rZoLMzWY8S5LGmYAhEsDPvgk9Ko
TKA3vYhAp1SNJNoihJRgKxQVxWSxXOVMzfTOYvvW1kQxvyu3OmWXgWw4PuimibpJVrLBaz5wzXvs
xvEqdnnf0+wZR4wnZNJZWIwSZ9wcW2xUFAjBxSjfHbCh5v9/HdmMdkyRMf/NMRy52ld29RZYj2HJ
MbGsKJJ9fqHTAKemtqNj6jCCQlQX6K83jYtvFKaho8Fe/o73ItuBu1ow6ywojMoF7K7RL0q5vnGR
5mhurSEY+01K7rk31HRRCn6ZMr8Irks4mnrkNRmPglQNwVgKvuqLHjIOXzNIG4u4B82ElB34IDse
eIrM2pxv3sgAr3BReFPHGApVPxLNGjcBAI/NaEk24DY1FXx6xV6wEBlco5x+GkLAZBUKLiZ6XSKZ
EJyjuFAKAc6LGgWaK4BSpH+6be+FOnj5yDmzWttA2/+kmuiB/FJiU9uqRdPvqSxszeTX6+7QuWsN
ddnZ9Rknb28Vy5Sgu3Osc3YGJh9lEDRnw814Tenee1Eanx5KvhMfXen8ZDjh8NenOV61rw2z2tjk
Wq95A2nBj8QGDE4z5eJlTVTD0BtIAq+bAT/H46+zkAp0HJbzBI/isTzsOD6+PRUattRjyaH6jOjv
FPhLy7Rls4ge83KFdIFfRAIuIur7a/zIXtQwLCS/mIYNoOfwboQ+uddccw26oTTi8GiPvZCshKfA
Cqg5OGpUX91KSk4vunQy0XEmzJroasiKzcp8Mv/Df6q3t+TxWA1AeEE/8cqiKG5zlE0WZpR7lZKc
33A4X31/vzUSgTkl1n0RLIys6Tk5KGxHqHUpO0/Cjg5QU24fSSYhcht53I6QldJOt0LhR9LTtuQX
h5o/AaTYk7I47rflBobBMhQhVudYaUoNf2eqwDWjZ7VrRr+VlUJ/t1HVsrwFiZR9qn877rqM2hVM
U1GNux51be7bIfVwjWYMaDzMUkthSy880JM4PNfUKkz+LhnsqIX6MKRsMpUaiP6chrtuNAkVreaU
SeCcev3tJhZljb8I3jPs3kPwgnhL6L6U+WkKqdzvWjjbAuMhx4k55hi8ddICteXjQ10htPm1CkLC
4xrbBDEvn4Tip5iDz45H+Xv0qtDnEpVmdUPobcJMMdihIrDp+MRejp6frSirQXygYmA5bHsI7PDr
GkKJoJZT9N/elmwHXLVnFgCYuvRGlSUet+Hrul8tPWCrSDwc5wQtpwHH8gDOIK+mRyL2bjKp3S0g
xUURp3AIUIlNLGo6UTCVtfavKdLZbfpq4Xa+IK1x74AW9yYu/L65uRdOvUIcj1y9JnkvsiEbarM3
5eT6yK8JQLCnefcvtVSbNXQcpmgWv9saICADkkndBXkrx6nymESuXTyt8cT0y4g03+a4cXi56tZT
TA/qlzVig4rWXqg3A+r885/azWeqGL04AleePKvKUNseHMaL1+rkf9uLq7aEIr3va3PegkSsJeCb
l2cj9OQbWxnl0KcFpyaBSeWvdumlVDRi5fqvQHULuUOBUsSkOTceQZx4FKQYjXB/bd2AEdUTRXb2
18uG6rsIIOEIYA4g+Hnqruf0296taf8Fvq4pIhv3KrV80MuTkzPJ2GTJb2YH5eJI4zdf9eGYAaLH
ub3vSHydgsvrl8Zp0M0EiBv4mfANPxHKlBV29uC5ytkz9qVxl08txAAwj98g8ixIopnNuCqERae+
6QaX6xnZwbo+im9iun9K6UnTwCbyhUjlRXZ8ARH4vuXwerVFSFoP4SAn0qxQhTgdBcuQvHoCdz+H
QSEkfo8wCVgg/oa3sRq9F61FmNr1BE/Dqn0KGplzfYcOTlnkhBz0YQ1r5QFDjYfee32vhOMtyWnV
7rrDmlMrkFXrOvG8kVuMLscbUWMNjfrcsGRptBySNYLLUwrC7ei/1BWwv0uqATgwWX+I7BEBD6ZT
gnN5EBzJD2RHQsaqdqgMjh9JPR478Ly2cX3kZJQDLQ9I1jeqO14uGRRu3OOZcNCMRQO+YoCpjc0r
K/+Z9aH83dZDxSbiVKrqtqpMn43hDkWh0pYT1h8zxnRUIq7EYTf65IvPRsbnhVgI7pQaTHfNoz4d
0JQxmAYW/DO8W44yydp96SBgsT9GjR5Gb75ia5LZL34HEI6SynyL9JOZkJlzNiQ9Z+Imv7JDVOXH
Egc4ZXOm+9XXIskjp3GOfhb+hIg0OzzwvMSQGhL5pSobdPt+X/KLX2F+IWHp3KGpWpzaQQ1Pen2Q
5lmd3ks0W6T+lYDdJmsG9uSOWms8wN7vK1E8gP7B/29uU3cXj3Jx5mWZOr82a6l0BvVJWfuGOrLP
2RvchjxIfruUydNuS4sHInbiAzuY259QQGLpGAou2YidO3sRf54XOexknDwU4qxBR0ish+F3WNFm
EmPUccXnyy5oUMuwAVJABJAPnEJD0gpXo5UVfQN9SPLeHR4KSbklf2oCLXAUXoi9uzoDiHtsuz3v
AwrRW2fGNIYoK+kmSCmKxSa+WDiwxBRYuCe0qua4u3Lshm3+8iq/nrVvvuqjj6qnUqAtNQyFMEZB
zaBKD9JtYrA8C2kk7cOKp7h93sAqKVTyRAPHtRKwXvXfNKx0Hz2S8wcMkvlpYTHz3k5shtjmyElf
50mOx5hlfEFFc2iz390Xkv6famJ0bMFDnLfqLf8vAfDGwCYPY5M8I/7Gwt95+QRe3Ujk871fdc2L
QBO6Jc1FEPh2Ts29fyR8nHOp/B7iBXk23xyPUodt1KR/hudH6WOXPMedfxXxHw7Yhoo9xVuw82Nn
tIswgPojQZDH0PICxzl+iI1hgQiC3c7u9pnZEkmovJ2pUN6U+q5QAfvVUJxqyQ42cdXjsbYem/EL
QXLMqXAVPYorsuyT5rvlwm38TE6t6CXnW7eDfw7L7/AkqZVdzEym9FAtJcqtsEvEcKuEc0vApKLU
Uq6LzPn3lL5kMAJUx9chmO+IJYOJQqx3BhJOdUs+UOjhrU5K7+HD4Mo2xGbjsF9biTO1LjvflEfA
JLZGbiThhh3SW6mXtZhHtNis2R0RqSB60S22zmw4SwkKfds8b2j4pgYGa240LrrLj1/CzLQaBsO7
+Ry8lO0CQVeaHrDJmX7CRgRya+g5Is7a05LQ6IsTYxGSnirmhKC2Vwiy7N7pnJqJNBsZJWEht4Au
NcV3iQD0XM/YLDKlovned3vsf7lnlLUhql1sgAUZkEMo8Gp8smyJ/DcrLqKZTsGnz0zkTeHm49UR
6zmaS2FKIa2c27ibA9DFwrLtnrHVNbt91HrIh3IgXzzALRbtCihcXYodVTgAuqFql+v7XMYhexRj
U4jVuFsvsZ/2X6ohOwGVr5SJFUOuBKm4byWxMTd0B/jh6TdDNwa3nRzxOl1h2iQv/wX+HDdT0kqO
XCqLCLmvXOFNpwQVewxF8MOCuZj3NsvGsitV4ItElbTOr2g34DUk0SBNLaFWM9oFQCaShPlb5uMQ
JwDhPlfLSJ1JpYnWMgSATpU/wVDfdh3L0cDtoxSzzlVKyrzJxZ0KEsB1jkL1L/CaQz/EYeinzq3y
8IBAlaEplQeIEjWwxftb7gWdX781TyhYPMfCUZbVYMmhXiIONA31a+Sd66SUHjVQ/Iic0wMolZDO
0A+UL274Rcp7I3sG/4JYNF/8SafMYHNKd3UyNadbz1ZL/3s11RnwQ04slMdeQxORXIAHKhRAUgoA
d1kdf+rc1KsT9+7NtBHKKkDA0SB3rbJwAFFzl23ITxjzRrwBHYIQ0F3mPAhIqz4JR5vlOwIKlJEU
szhALLawM+Cdsau7JHu6N+b4plhsddTLLuTWpSU6mbgy74MgP9QvEuMavmy1pV5bYMz2rNBnGUAv
JBaqjbA3amjL2N8Bk3hoI0UmOWISNWst40RACVYnQ4dV1PiX0r7kwvcPwS9vuEAtNLd7wk895mxP
Fz3teml0GKL2ojXdlvfuTesUTPYlnbTRbKEpXQkBdHzEg4xWPhHwoF/fqlDyUGxAFmJGKzlrd2s2
Yj0kG5OvBXYpz9jt1eSOP+pLvuDeiYFv9ItAx2k7cxwZBR+I98TXYPc8LJVEC/ZeYdYmzWQmLVDZ
BaDnP93NODLWPgB0MwifcvDTTRGU8KFAgx3H25Ysc1UnQgNWGg3xG/mIOUsRnNaRkLwqsumCqWUX
i9ZPc+xYHnT7uMk2DSAZ8rPvRzI+rOES4+hzP5lhYFsrsNmUvOYVhygDbuonLEUBI/bWtZrAWg2S
knBR9Gx1ffjLg2LUyviW0L3grHshVMqhZhbZTraBSZaJEB7VV+t9g/wr9rQYEqbvl1j2rzS0tRGd
mx6QSvg2h1nzUqroiT/1GB16f0O/fpwOTp+daGXUO55VlqMFYrGZCvc/x9Cn1852M4jNBcl1jutd
NnavD1JBf2pdooU+imG797cdaVMI3+7Dly90weC4/cRnqdtJ4bfGkYxApD8tj4ISuqKKyD6LV98c
njzrAzTe5nKuEd3aO9ePdoF8KRWpyhdz3Gy2f/o8Xfxh2FcEvceIInGD7K5n+MQ2NUybXUfk2LLw
c1CMxhgfHNsslv3Wgro++kag+8dFS8KmQ5cFb9oIkbdXCPd97FwYqGA+fzf30ca+giwYAvQAsyfv
vhodvbBpkFTrbd9Skj3sRLnbStc2QGMy7NE6Wb1mV/pycIKEhqHDRLy0rfFLhlIXptzt7IqS09TL
NDepTzl37yf+Pei4sP8qaNbz1YZQvnESsnFdxYnYjdAaJ5TeWIwpm/Ex71XZCoDAradLVOIQwl3I
V+BtQZliW+Ucicaw1awxEy7bDpeItciv9JWuNntyvB0R2WY594yoEueKZEDfQJiAnWZQmerEw66I
97RjlYpsDBlc3JNsHPVfAzTsTdZxxbXv5DEu0zg/IjUhaGBPP79pXXRN6nDErsi+FQ5mJHDQPyGD
cMax+DJSJk5BU7I/IQG8VN2Z+suTpnVAl+HKE6DW7T1RWLyo4cc/DDjlPbuFj15zFupKCaRrS/8m
32KlGZeXmqTBVZwxdfgq7sXXEU8Fzbv/9+OfD6wvFEmtEoBlt2IfraxH9r3iba5H4ZAItaEHL1B4
q20kmrv4/vxAT90WJwCmCRWuSsy9X0lAra+AarhP0cmuTGUF55n3WcLi/0/CQo6ANDQwuq3ROVAd
TEtV3n1MPOix9kxHZSrFMrlYUb5YT7KNFwe0BanFU+oH81/RZ/t6r4vTLcdvRXJRZnvYvxNhFft/
MV+u5trxdZnCWCdntYV9maIbY1AwShMRptssmRgiHAJ6xlGBGBpbG3fzi28+W9fvJiP0gqhzWSlD
OvFMcrYfHReqEoAxvhu5fi56t1BRSDSjqyu5D6ujjtGw9YaLbqzwXvkD9Wgaj6cj4rnPe7x1ywV9
vBdI7arMOzf5Slyaq2hR+eid/a7lSJXEvhWOPN1gl6M/T4JUaNVs7peyZCDNgtBXmH83M9Wqg2Df
g6iHNmUNyeAweuaRRO0ZiXucKhro8/D+C+ti16NBjzPP12jZQRncoMra+ghGP4MBtOpyAultfofr
oNgpB5jeo1ZSoeIg104/kQ2pQWq+OhXywgrdlJgxP0nA9kChWA1CvE+42Pl18W9xNcy7qx6KNd9i
ga3bTDw84Pj5XmQPsT4z3RwopdY9UcRISpnoBR0riQh7Ce2x4+tffPWukJ5VJE33KgEz2/MdkyNT
LTEFlgNmYFukYb2Xm8GcuO5/tzvsEjRJzKznpFxe3AyydK51zsuwWJQeomINCdYICc3VPqRD15W7
5Zt3WVMBIIKflncZQrWkeZSxDl/B5GN4vPpfTDpUDn4NqMympV7EpdoPUnFqGc1whzp/XnoBwVTO
OCmXIayrvIbAqFyhX8vFPF4TP4X3pp2Yr0B8UYq1Dxp28lqo/YYQYEAY+h8G0ZZuYYT32Ng4Afd4
eVx4hTJy5pKuB9pvXc4ol+uaERVcpra9mTZmJKE/TT9WANgI2WEOr+Vg3CZYRnCCuWjr9OxUqHj5
7psuQIzw1meOIQpVNYXrTalKrJi6nHlOzYsltd3iy3m5fpuLKahZ80cJutr31iX3uoyUxXi8gFs/
f7PIyHWlstT6B4H/sqRYNEyIPOgt6jamF7d15Uf/jU2F9LNvWYcfCBUHWdgya/f/PbVcO1H9TwC6
aW6JJTL24B2SRsq1r5G0KCoSLsVhPpSjaCTk1qs6dUJIYlI9qk1QLjMZ4Lh+ZuvJ0flaHGssxFG2
Lct6J8CwXvdyNgEm1fSuTm/jmwUOOiSPmUyiwgiDomZM6g/B0+A2C8lIqHk2uLM0KnUrFiuDigR+
5ITQvd4WrsuVjOe9AIJn44x4ByGoimTFMUG2zxFcQZigbiR7ed5BfyqXPfTTBCE/SsV3jfTEf7ki
cMn6NnvIWEuXYpn+HhtuZf0DfR/8Qo+kq664d7F2WYg0AAaAIwMJN2a04XNys4rP5FRjYljvAtJi
vE6yN9Fs6rxpd4nSudvGhJ6WLLY/jfpGm2ah5cEPVVF2GbgO/ew6sxPq4g4DnUiErm01NZbXJGuO
vq0j9xydoZ9CL01WstFaD2EslF9f29go+krbvvACxjYsdSA9HpqYTFJSAbngNGB1HlsjRlyXIj4A
UNbTAq5idvLxx7VB2V6ED43fG4BAp5Zm28vDPJuQWrDF5BseT+lmw8xsXV16pNBoDbH8cAZ2b+8o
O0fb5+MTScUUcIVxuRRPKZjsquEI1WbEkSfltkwnVeXHTqcVR/0udrdq4QtRReVsbcSqeqMClm58
q1kLS2BpV0qJCGa6AarrC7V+3xbXGTXvaoMG3dM37dDvWDXJ47DsN684tmaB4Beo98b3tfR5lfWg
IF/nVrORpD33hHbcEsnkqpDutff33ZlDnSdQJuus/4O/yRABO6R03qjJ+N6TV6UKmb8XBls9tg9o
nvXqsy4ZSgF2N80Pe5d7er+RybfGFKtDna3zdPMLq60GmgxBhxmDHGlJgZPBbTCgUNgqzyDMGkM6
uBZwX1bocJDTzgfeZtuJ/1GbfEyymAU/gDk2pFQfjoGKwWVGiZwe8Mb7SAXy0bQEMkFadykHNP7O
fTYSgySCnPSyNTalOB3ct5ZSZyYutn/vwnDYZqv5CFkrh6kezsSBZjwzpfJ4bM6u4r/kzBxHNKHb
zosch5323oGS7sL5SQexfi28Qej2RW8T5HKJwLGumsLHsU1fKQNWBLyGjdFrAU7OPwuDU7coUID2
UwCv9YmRtnVYoczezzdxxryCvtzKDIW2fDsphyrhLN87ZXIPIVMwHjhDXqt84OmjHpREzL5KvkF9
yXrxXF00xvHgIHdh+nScik0HODKVewOgO6/SNNBkYtd8ZRg8VhG1ww0BLWcHQWKa4lTeE+Ru+lY9
nQNgN4zhQSD/1uEQk8KZxETJ/NP5ub/aORVDKFd3HbNGaHGhIn3YoYogn/Y7brge5nuQGDSzjltF
mTpqyDIxZrAYjQ0WbJngpVagz07/TxtN6u5hJB2nHuhMntsHXJccY2nrXjlPGgtyf8o+QsGI+Qc1
zNhdLtw3qhanpJrixiezwxzGUDw4uZbTXXcldnXUCCAZrc9+fu2oADjglOmFwycpLNlD3jDLnr4I
2HiStfK6gHgRmb34y7GtZd7VIpPRVhvzwLraIJhb6tDqNoyac6jJal0u+pqtOngiyT5qH/A7F4DJ
vVJieP3SOvcVJGe2M4UqI/rW43MZ+5z0oT1bUh/8DFsKUnPQBiyI0XglqKbpcBE4Xguu+5PwW8NX
FVsNBO8zvPfivENKZEXjOwTOjOaaV+Fh4TFmANT2H+EXvpYisl53gNcw2GhToryHx8tCiYHAUkPG
TKmKc3M1MX85IaKBMkhQJ3UfSaZxwC/q3iemzDl/uYFrLj9JVOgrKP8+6fXCssjbEMDnnB02947i
k/6lU4Ss7nZzsz82y7MOu/PYJ4jasAzwivJkdcdOdmLjIN4UvtEoQ5xG1+Uv9nZtVTXyA7V5wKVh
ssH5cRAEfdrj64iF3N/tUysXSryZ8uDiBV7m4N0sbXY6sQnlV3qcWFcqw4Mv6f/RB3nh4qPsoIER
w27rop5h0ppJspC8RsGNhCWDHaYoJx7V3liPBo1rk+KWrdfZY7qOpVSMIFRZ2a25MfBM5Q99PCmz
dvd89E1tMAGmPO5EbNsf5sU7BnKfoe2juEha3pld7hyXYgAuBxP7Wwv7iAZVLTYXSKHbdfRdsaxG
v3vObdCct6YVKn7PPuUgSRAif+C297ehfcj4XUOMSotEcrDUCxdSyvi7NjX3cg++eWlMl06Abgh4
tDIjfVmvXRbnjuQaebXg9kEWefBGN/jBqDKHMBnyZM2DgbLzMM+/dN+RIp86qud7HrwNyROidSk4
JLtYj497psC1LneKlmCYXuEmJurNkSiXSN6eSi5ow5TNODdB191pSkUk7S6+aknzLVycA/bAeygO
JwyRguoRbQ7zdpZ23vLQZ8LDjdCb2TOmcgkkujbZxG0H83da8/lc9XOrWmd2TBPU3PRZOLAWQwP6
h1svqDHsFknfunjHDuI/9VjoBamINWIrMc6shPwqI+5hazqwuwUb1GRhiLtXuW32HhC7q/jVkquW
0GqloJ17TSE8wj4EG1l0jRVe+RjndJ5Tg1XQaYQNPG4Q3Rm5lTDLrlVPVp//wH4h6WatlJRByxV5
yX3L5kmAWyJbVZeyE86CeBic3Ypzko8/8j5Y/TXFKFggR5JvpWK42Cjrz7MqYieyqyW/BdOcSoG3
he6aJ0G2cB6QCJeeavD7IFgQcPp7oiBsBQBm3OblTjCoOrHxw31cv8XIWwp2Etadq/h6bij5i+Qq
KrB1sPWhp0TxW/R8Oz3rLyOyiqi2q5/SZW3DXw1JBMgcdkF+f/TxBY36p/8CHAS7Xzdhq1dAalqe
rz3n3nqHeoJVorP39B9sKvzB88pBcvkxUndpkYA2M3VCPwfAbDKwz2MzaPDIV96OPu71nvDd0kq8
ckDXTUyErOeiY+/Yfcxb7y6wp1f4FIlyRtNqHCf6m3tAXjtj492DqjeI90QL9W5aPesCplUhlvS8
ssvVM45MlGSk+ZuZMNLwcSEkEd9jcrfFAwwAr3gqkbpWlNX2QGVtiEorn+ruNQDEShWln8rYOcj7
iAKb5FtNJFtrJud/4IISTm1BdZef7bBUOMRV3GOd8KGcGh0vDBync+4OPwURDA1J1ijKLpHBNsDo
qKA+6wVmXRmv4J8LWgCTxPPT3DQlpkUJquESsF7SLEev4M46/RTEMdkjk83o5zhNUv82Q1Wr+Tlt
BaDebU4NU08EPfSCWRI7BebDz3EE59346g7BS570wkvKQ4LrE5XX/Vm3KtkJZTdWhwTno90/1p4l
vItbHDb/Fi/itSX5gdAsPGOxkW/nqy5XZs2Br8pZ91JcugFyLjuCzsQ0Gv4tMVwOvlxJkhwityAO
LXyCsYzrOm1pPAgeK2bOgBFuYxN7BBrutfG+1vjOBV5A+ausQnVLOUR24I2BrhJJ/gCKvt4d+LvZ
9Mwl2wdoadEHMmTUMNMEqYQAksxSAxwqGJwapUDiCcQGWZj3Cx2f5lkGJQw4Xceh83jPN3A8Ic/U
cm80fEio2gOicGbMlLEe/S5IHSU7GEF66pz13HHefkmkfho59Ya23VwFrGMYvipN5nnual+NPYcN
th+V3IvbH9jO4fwE6P8h5fZSuP9copwbh6w2IS/CZmJ3z33R6RtL0bIAQC3N9xXduBiLzvcloJb6
zdn60wF4YJPNAw5M9XoFtiLGpeKqfofAxQGTqnNuFHxk8m4xerGxZzQ6kGqTj6O7hbgcU+t860dA
nKEm3OKxIo71gu94TFz64023qN0HZRNYYOmmrQmkgca8NA6Nijw8lgDU/ajdnvl/swzL0teWa0nz
HUIr6akxPqjQurfJuFq1U+Skfk7G1JhgNq8leKKYAoNUa8rQVdrk1y7KT3UzaXyIfd57xx/Z09lN
XKLhmt3xc8SJYcYvu+Fmrd3GvSL4EKWUWTESvwI98RkQNDGB0/DZtsDblfgN62NcPOLbbp3cncb2
666avky+j5oKgm0il2WTVspGVON44xlxKZo12oZfBq9069OFHoBNWe1dSvZvxHsKUhdBlaujo+H/
g/1btsiKA2G4csxLSbX0nndWI9rCaA9L2sT7oC998Q1jf6Jly15InKyLSRg/C94LLCI4oizyBKiw
57qqpmOZtD743bEO1Yd9MJ2wWwUs45MS6J9M0enZpdCShYkJ/Py1pyZ6T2vOnltJXd1fNRPbsSKy
NQIsDGMOIMgeDHM1mIExbOp32foFwqcLip8QaFHHxeIuGCC1KGLs0bxMW+b30zT5jVsDdCVLqJN/
MBPDpJAHnk8j0g7qJbE5eyr+Q84F2RWkv+iIGuj+GoCzEn+wGzvvflxz3ABBaJIBeTGze9JA2Ets
5ynk/48AYm53Y9Qz4TqD6ubF8Gc7PGfso0cXgoCplcYZgKYEnSRTeuQsvPCEScj4tyjq2g0xQnFt
cMRFEy3P7rS0QccV7ojtzitEPlLcUJnQgV34lWQGIbTm28gXvkOlp2AnpEg5raOzrqi3fZvcPCPn
um4XtEMi4B+en/irZRnW3zDJ3uUUVqrVy0MQ+wWTyKYxplS3T1ubYRrDoFseDGUvfgIjKJtNDZwC
mxnfEAjvFrhI4GLIy1NS4em5jLerkIlm2+YahomCHmYue6Lywmh7x1A0/L0frcSeA33qBHxiWFUc
kuAm5KL5N4FaeIdnkZBR4RhtPBg3XSYRFquRjo2ASfUTUgloK3ZUEMyXIrj06aaPpv11lhAyXp3T
Lz21ddYpfma1b9LF0u0IbFOrstOibuljGD6deyw6g9n17nGNUP9xtjaxJZXuDUGBXxBi1fE36K6f
xXMCrXGpxuudQz/Z34b7ga++G7WchGxa54rBs4rCTGVpR8qb5R95ivYunkFtw13BOXOXZg9tA7WR
yIHnmFZrN/pYdz+TX8WQqfEC0Nihkefp1cAwuOwqzPnh+b3WZct2lmneq3csacuo+lSw2qj5xYVK
zW+iNKRbaOOUIhRFk8WT2sh520Qn7i7dx5qOS3BOwe0pRJ2qdSB9VwZDtKnH2kiJnyam30GH05P+
6o1GBMch/73avOuaDzduIUsupBKr5oQYQ/CsjDm4mujPtPWveQxVmDtfbiwQ+NrnvpKVpEMWmUU+
fPShOGLg4HypandROoSo7w8Gg0DCOV7NhlA5xjoL/BF4oCdlpBCnCxR5P5nb+I/UzAhGSbKKtbRU
ri0G5/QoZRhXtedsPDenbrQZ0D5sXJdRl4n2OZpfXHKFtzh+3XLCjEnblNPfoDnswF2InUAbvzO+
VCaAKu6axtrgAp9D1FJuhmLm17+hsnXqzgsXWNuVQsKexbkOMaDQxvEv6Z9M7Y5aRN782yEx9GL9
HUJiIx2Mgi5K7Irt6a84zxzD6rd848LVWpojHv9dJaIXHBvIaQGs1gUqeIwJfSY/pMzDZXbdfkaG
AToDKSjYZbMGQiqvChLnPcOWZAwH1PMNraK1wkzl7ksokVVbu9dnd6y6sAnnSL3Yzsk90DZcRjnU
mASy6TGHNu+xUaagE2hPoh5z6PF9I5iURAVG6HVVkC2iRUX9TdUPPGRtl00ZlNUUf8K1RFDFNIXk
Kvn+hHZFlqYgIAueTt2ornY67maYY13eIyzzGfWBPwUr88vq0mqJoYVfhbgYyzZSY8Kzgdbp4MwC
kPggD7NUxcWmpYDec+nRXEQ1NWQse7rsIzW+T8xg6tvlnfJGSWILjFArUjlgyDL1DlUwDFCXsCBV
tOrMWyNqa55WmD+GToBkUV2MU07dha+SO5qiAeypJ3jVaGH1Aza6nYWsGecRH2k95t0Qi+cFPLaR
JADsLYFrN3dYxw9fxFUVLp6qQHXJQY1IUyVdvljXiQqo5Kliela6Gj1HSNWR01ln2t6js1Ql47MD
WL9EgafFe7xrRSu6P/hQ9qMHegv6UjvT7t6Ggz8kgkHIllCBXb49bWEZoi1oZyxduv6CFb1zYnv1
aQAPncqk39+tzqnbroj83dQ4HvMSc64VwzxqHTfi9DrgJUNczl2tEPY3r5qFMaPSlN4dVE1XXbSA
pTPJ64DdoMjLpvMptpwZrQPMfrs8FN5nZ+hMZwTBsZ+iSLRZyegnFe9FM6c7EllDIr0Hq8TM9ije
qzoHSFi22FzyUNWTSykbCXq2B2bGPct4QnOlFKeTemppJB6PPcmfAbSlcuEL+LbqM0CoX6U9ovYK
Mx2AZww96MxpZHIQuUla0tKRGgGBn5rAJp3jtqLT5vJTlz/ib6p6PtatQzUcIIht9PdWeRamRBoy
91OwtSLww5QjaoDMCe00nbErXT8PS3lxuBzbfskQtEVaJRlEVmY8ukS0Papq7XQT8+pxDziiZsOE
sF+jnGdAUvM/oDssU/8AyXQHmROTeWVLqRHJsGWZ5DINn03Ti7S+PAgvIM8XsXSJRnZ4GvimqSlg
aJIgKflNz997IaJzN4dHta8AuHK7iRhXr1AanCb2MEa9VAbopil2yqq6F1PnMtTxTe/Jb8WbDG3x
P5cAuODlCzFTFh1DM0Iun+6sNM+GcXmQYeo2EL02DfCiVnkWhVgHJmhk0NaKdpXxtOb+c1gEgGFb
qeozBHGLKTGZHsXt3gY3QcGm5sFLoaqhT3oNZN7i9sYSe2lX7k8QwXgun+taU7Pe8q8NRuS/VBOx
X+5Uyjx2eAq8avhsSoscrd9AGkOSjHr2pBNyJGWJ+tpAWKC69TDuAEYFY0A5vIOlK+aLsSpW45HR
F6Lg8Hq0b1M7ShtYT2U7GkppZdunYCcmja07ya7nhhDmEomXSgZHqXj/LgCpbSKLAsY4NB/4B19f
Sj6VKfoOPdmE2QEko8+tAEVKitlbu79C3ZMOMSV+ut3Bj3gajUuVAU4cV7FKoJXHwLrpcGLgn5wk
RuPzQitRw0nXk4Sfc3hwfLO6GQcrN3YGT1REm6KppZ359Jxqn6jiuT0IDjMAikUb4md9I9Tc12ay
ttdS8j4x88r6YZfk3YWRBVwb/cvZc+fofqApR3JTNq8SjqMAVIv/yOuYKDQZahPczzoUqNrjODbv
SR2VUpEcNLExlekILuv4ib2JT0QTAnonRwew6zxxTqUovVoq8AbKMC8fkMBnSn5VaalZ+rg7eeXh
3jvtjlfbA7TVRAQaaUvRqfx3FQHvp35gbo3HoQXuzFpb97F3vQzXukeXPlEnVVTHQh+O3ICKihE9
lRvJuh+rNat0xixvX9bV2rJx26kA7/XTRN4DMQuyvD+3WgfZNRoFe1ZBbQxspRIKoSYbQZc8qai8
YmDM7S9tkAD7AEd8DzmZM5X2Ih+En8qRHjNEHhTHF/ewejsY18HKkuQI0M3dHCf56noTbfLcEb0G
YpsIrP6gOOACSwVhO1pLw6jwL/2e/xX3vv3oy/BiwAW8f+u+biVUSYaAHWuxlIo0yJ1VzAKrcWY3
dKgJbSZLG6tFkcQprN3aa9aEOsa716A1ZHlzOm1OgRvQOnAgdbCFyAQv5VCg2GxexQQwZlU7eunT
fhAVH7nscjNLq+0hnpsum43D/XK3M5EdixVDr8/jiATsjc/bVyuDYG1689PCi1mTjrDOa5YnW4vN
oR5edR5f5K/TpGlapF+uyF6xaUB5SlZQkVtWd6eQAOvMnSEPZY02PRtKkEEqpNsyMs5X6tuHUp0X
cxLzZYR7ogm0ktV+GJilYvviogr2O0cAQl6xKhZnXqJfrhQUNnkbqz7tu7PGcKNB5bitCqn+aTxU
o/rJQbTQTIOLMMdioC9HaMn0y1wosTp1CWyCqujK48kpWMV96y9vrxsVkIuiLPud6J5XpSf+/kdc
oISnGKxB3AHJpls4TJ7tNHGDhun5P1409yBja43Z5QBWb/2q3h0ei8eR7IGeheRfs+ZTafXFnf9u
zeiSy1kjZjWIO/JDMr8IjqMUVBFF/MT9yJIkfPPWaKhx+Fgmxt76Q7F+W8e2xzE1Jc/mmcBtbwnp
GMlm7y47l9b/HykLUlRuJDNLKrwD1pC8B4v1EvboFHL+Qzut5QMZAxiM+61UOefs3cIkijCFFqWG
sTu7O3QVFOVy8/24kR7Hv8epGdtxmtOUCbn8rVfJ1SDoZSKRibOdSYWOz2sDTa2pN5xJBDZBtXdD
l6pnI7Dfc8yEjU0/4A0w6OQxvvp5sA0B8zi8rRdJc5YPBkkyOpMi/C4HK9WsmK40ropsS46rr/wG
qh+EscsJHPOmQHL8sayAiK4vKxjMb81sBoMXA6FZz9B3J7dKbbEiVEw3b+4izFsRxEN8MfotHFAI
o+6weH79UCrar5g0AhQZewNBKU1VgjxaeVW5V+fNW6gtc8Ti/bE1QXei5bgCTsZUXQqDUgnfVcs2
NnNR3B/UBBTthtL0MAxYdYJP9fibUHGYv7imz//i2KCxXUIlcTSmoPUdihHXsoJLbZRTBh0O7eQu
7SAr/k4kniLvTKY4BQBBL7aF44IZFRLKrqpPjL7W8TlPCHcuFwXGCwKSjudQH6ZNvkVgCkc7AlHA
RSPNSG9ql7mqn+20Tdnt0rrgP+wwL9ma+iagmuFPe4/4NYV7GQfeNp66xmJwyWdm+A1PcsKpjMPC
d9OopRCSULjvxeTNzXAUvDPwMxAv+iLYuLD+68MBdsrUvDBRc3pZNP/OSgX1qXbirNcmvk91JZbH
VY27mXp4CvcOJPwewK4ZsOlFIGXW2GpSQEMTooHIhXBcYDit3H8w8iDi+2KC/NYunvSS1oLcxk4V
ieSeNcnd+ayyPRq7u+/6m+KjJlUYXMi6nWCU9+OWTNh0lotdzXfqP/Ckj9cu8+u41ooyoPeJUAUA
FqkFcPeRrJOADMqwmi83hFYMxXwwYfDBaKpSAdP5ngJYD7b0fJ+hdkYuGl9Pu+ecCMsvOoPjISS1
WkrZJxWFnoK1rADnqmuTUc4IwDVhqsy1I7JnLzvMdB9JGT+Vk+pCE8RoFZs2ZPC6wnuEVscuvrcG
oCOcIsI9e0DvQ7O4qSMqoGL4wPw/zc5Ot4pkjwtSbdPQOaeJ7wKcZLD+qFSHVQ1fdPuUWk6pw/CA
ESsmhrOehePGesR+5aSXFDyonpmHK67ZpsjrXJ7FQJp3rqB7jTFdygYiYMihpCRMx5TYneloB0OX
FBosimpFPQVy8HXTkRVzMXvZHMFKFQWLzugMyMN4BQCwnOlycL9E7qV/enym8Yx2XBdAbD/Oed4j
EpJxhVU0DTkbfj4gJHmtlZ9g9ANsx9ROLli+rgICb465fYNHLrVbm2/T+IZ77ENRQWdSs4iNiF8V
x5nIyKcPAp1nJjVB9h6NMbk3tr5vNJLgfAYXUgK5GClYtLqyZ7uIWRiUc/Uf3WvhaJPrceSkp3sX
lDExEy6dvy/61Ke+aghgTbJJbHRqNl5XFQYHd6B6WEnZj+r48OLHahOUxTHAQ5DVEUqtYuOc3hdb
Oqy1WdzCs7TkkEpFtXStBlFD/GVyE4J27NghsEayAxNO26t3HRi722nIoR/unQ7rBLh6atVijGxv
cxSwL/DcpnNBYEVquNWB/TXHKy/44QTY1CgBhPbivwQoCZs/Ba7cQwEyldIl4M/LI98CFx2itBDI
jkD4BqPkII7CxBIQ7OT86LygQ+LkLCS4Q5b1q6Xb/sgYBX456IBPAvS2UpG+IC7Jv2nAmgIlRaXM
VAkxT718Edc6+bkOIBFxAuefgE4as9kigedHg8Z3ugnTzD5zFX+27x1vcQaXdxXpD5aNy6GnG8BE
alslLmGtf9rL3MXhbOCeGbPVxnQa0g6EWUv+fYz55308vbHdQX4KerqmPp1OQzYgTYWDZ9yw2o/5
evXVOuJGlyrjxcgq/F39OOPzrPwA7cucJz8mINurk8uaKSCXKPudrtNZXPEotK2O6b8cDQg53Etx
RUbFywA+ZwjP+S6IdD9sTW3iLnhkFPqSzmTvs5JPdFE5+ztOoqVG1QBlrBRmVDU/bKRdTfI0I/i9
J6rqq+5o16+hz3zX5MGfb3alU58pOlRD2CPa+Qcb1f5p0KLdUJEETJRbykIjwHZFmVnFcm6ZJ9bc
fPWYDiZLFyT2EY9pk5PnZplxk9Ntvf+0PdTuqCxi35Lz8LdBPVEU0cFZ4+7+7x25gZl2+f7OR6+J
+lXgHJ7GC8BhN9AwCBcS63xUCxOJVPYk63LanibixkwZwwsy6r7tRmsROJAoMKtaQp6MQ9yYIwzn
y+HT12+WoErE4sisosD19bnf3UjF/lDTKQJLMjphpTlSJ9R8W5CFZ9KxcwyRd5gMO6N4k/Wo84Be
z0Z4ZMilZA5tx9C3pANfRx8vBt94fDYNhFk37ifwmVxnMNWcvMYMeB197awzv95pMspUbFRCrhz+
/iZqWjdf5Q0rhtPLYyhUetwxmhPQw7Jm0Gtfed+5Khv1oQ4Ww6EFp7uMpL2Bdq0waPWW514gP12T
1Ew6pFXJEnIzUrlbYNuLHVFvz3pdR5GdABPt/87TAV9P++IrcMldm1qsqWYZDbNoVUU92vJBR2Ac
Ni7FZiVDCYOYd9PhX263Y5j3HEYKxOtH7mMcqU4O8WbvZQzfgyW5DbJ3qwyTccI9Qja2HaHwfylB
BHrzae8rEjfDLbieI2m/18Go4p/qFLnzqAgI6IvASsKpJlPpfXKidXmcP2Fd6ZVq+x5WO8SqmQLQ
k2uhOB5EtmmEq3L2tLs9b4U0OCMDitjq+ytEbJPtmdSwLjbjhOoZ2L+CwsQ5fkoFJI2Tjb5yVsC7
Hy5bjx7xUCm+KyUx0nTiVV5QVIVeuCRqlVfP2zHAsRV4rmdTTK9mk1tMJqpvnxJDXENsVr05+aKY
Z74DzGtnJ63OjR/0Iuq3lSt48FKHb3vbCBsGsxpdQmQdbzm1bSseOttpcXdgexp42MBg+Yj/xdxx
Kdc2Bg6r6VEEJd+ZZMYghXmQJzpveHyLRQBvsYHJjYFsSlJZHKCV5IX1RATAN8x+NtFLEYhEb4xt
0vFptypmg59hOkIB2dg3x7eoqJUm7OS7wUFMcOqn3NNnY1dIGgNjoDUswokBjez50mlkIutwI+OT
YdDFLS2fOk7gAPZz4IAEKoFkQQuSmgkB/wYPXiBURWfLIxeYI69SmgbKF0mgmn5vu6sgRRCDOqUG
ZaVJN5zw5IWGx4N5Rp7p7m9WHDBcsKeWG9d5k1EuU5lXvF6y6TI9pfnHT8DubkGiYs1OiCzp+kk2
3jQrXoZS8FU2tw24JqwFRgtLIX13Dqtswx72/PV8z9ndYVFMs0SKsrnDUPEMwxtgel3ePyk8OuzG
Rn4jTuyhyqdh6hkjc3WJ+ddvrzr8knd6Rf3k9BeQaxNDcfUzvVIBhGfb+ASAG87POr/N/rK7AbAv
H2cPxNaoHTsD/ECDbQAYdToHj25ClrHKVoT0n6x1YmM/19SXDdxYvwhLeht1PjvxhQUMy1hFePsX
IllSqpj0jFN97LqLpnruvBJv3WVSWWB1dK6xSy5ePwK+E4Jr1gORln6whRNoE8YJdkxilDqJKlED
NJB0SzTUBlU7T575giAku8ZteewwD9fAU+tpfL+rycPFiwkj7/ZMx++kwJJ5Hj/5cn50jcVn6O+z
kMR6Ug+zkH98JgqGnHSuvITnRE8VPnUbB983oQmQ5m6JM6L3WUnmekGHs/QksEEjyVw5VLnQgact
O/aHm2QIKLO1j24PVxpMv6V0VSDbb21gR8lmVicMSeUkMOkI7YY9l+syzw4AHxUXUdpNx+6/zXeC
AndW++Ouurtoldw3PRbmwQifWAyUApynE6xpuAJy8FExRHD5joOhhqidybv48ENNxzZ4jdcFaI8F
BPUYYT2+UX3/icvyJf+SXHyiZ4yEKIwR/LuCMWcL14Z7AsCTR1o3IvZ8YXu3M9PJ9WNPgkVDVfAZ
w5NFucmx4N6d4f3rSKMx5R+WqlP7zI+DBiny8rnJ8GoTVdES3d+zl7NoDVqn9Yu3EHh71lzF+ed5
EHmGhuhJ76jm/aWFtizKwJL2VzLL7WnTsFq5qArxdCd9eIA40Zv6ZZLIqjDyV0UyeKDrSU89j9tm
maUQzP9QcJ2kDWt4V0zGzARecEcoRhnMRy/XXLlhKRjqq4mBdb5ckmo8moksD/+SffYvX6iLHdkv
O7VpBTRx+PIRRZE1b7HRtDtdbHjJAzd1CRaqK57pWIW2XWOg6FXWxERrF0159T2bXrqeRfzm3R+I
aYaOat6QSve44EyUOt09b9Ak3Ph/ey9jvwUzn36UqvcSI9gEm47OfTgbVBed4psCU8P0iyGVKZNF
HP5UdFMdDNkiY+DS3lD4iowDRIVAFhqixkNjJJO4nOTb6GM9oGoOqf7qwboLWoMXxn2E6i0GKFbs
0Vi5qOvQOHad3tqmNkD5dsOxTnCNl+rIx47MDh8IHSUgXj8WX96zPgH9HnmHTNRLl13iB/C5E8/F
OM7iM2s433znpQObBZ2zYWg7TS0Uosc5i/sU/tyK8W9YpFBuOzsNI+f0/2rVSqNX7mkTYbmFOwgo
maM9SmqxEUYIVrkH3NZBB++1dSRQIob5VdVEcL0YF5rkceiqbUFncHON6GSR1ygpMvvqOaxGSLlC
GDGQq83JUAx5FQqY0H1ZH89gkovFPcCWSzEe66oUPBGlVD7V9C62lq154P8+DID2TjIo7rR15kEE
p6S8+knbXAc6YOEB7/rFXMak9emiGEBcSXV3tRZD1lXauO07qpU9ctOWrR218fUPXGyMChP4h19B
VesKglxfOONbP/XYgxxOyS2usSWhZq5+WChvsajE8ascli0z+CLnM4RS5MCdex58iNFPUqP8UZPs
RlKgU22BMkJwy90mpF9Tn9NbYu0YnXtTJa+X5cFWJ6rVgqm8OnJer1sp05UTJqSkb/Yu2ED4N1RH
9yA9NsT7Wp5rStuF3YAbJ+SK31TmQeTYs8ukclNp0t9jXWFq2j/VZ9mycHPCTbiIKMskm41yXAso
HeuSgXLy2H8W7kZ15uvpQLWhV2X/Y0ErpEGa/zkrDbZA3ZSsktdJ5Muf5I1E+8krXM+938BIMTyk
DpLRLdDmJJ5LTeLAQ+JGTjLQUgLDCjmfkwvP80JZXHYULNgcLM9mi/UKc4rKG3tP5NapOi711Ftj
uDjP0X0mu07NX97f6kcsDBlE5ZM6C3wrQKI73Ru5T2JGS3jcRi69DC3mZxi3n0goLjjm4+RUYkWV
YsIHD0kI1CqFuWnTYoKTAyyMcnMLwdkcSW+KJbn9xJ4FakbB/tatJ/+FwkOX8j8LbfIhVen7yxKn
HbjSq+Xe+AuYtMNhSaU0ZawHOB2eKXHxThUCMTlZbNpAD54uAgLUeIpO6XheLLAhzCodpMxLvzIO
5GEYsLRkPMUy9J/ra6R0dOX2/nmdq2yVs1wj7RwYsult5H6DHqrj1OZIn2HRqAaA/zgAyNH/PZwX
+VSSMB5OVLK8gKKjktj+JXYCBYCTK76CbKhx73QpI0rLFYWMuzzk6B2kY2VoNrfRlGmOFjkaa23i
ygM9+UIRUegpNAN62BGnRYUn+w/4wNCPgPhRBnftDy0PKyReiaFFOcZAvPvxF/BHHqgV3R4VXx84
jc+MCFa6g2mEUjFkIEBDzRETQpVZCT8rxY133b4j6tUB5FRUpLveQzX2NT9uf1K50BuIE1yzvl8x
i0Vqa/94a4O3Nh1dcPFjxsP+WABEUKrqS95Z7WkAfhTqux5jtaV0lyughsi/NkVu2k1kayuNbf3E
uWWLhltrxWUV1aqqnTMfdNBQBLq6FzjhG719AdU8wTQ3b3HaWzwOJeRQhQXI8T1fAitS3geOV6s/
je/hmf4QM5XUsCP/TU0OkXCpv7THE6Yge4oAEZhg7gqPF1qlypseYUYToZpE6a/eAa6kat1wLNn7
UIXI2Usaquvu7whwlaCUqehhKf3H8h7IDSJvy64i5OC/chIzq1Rtxe965/0O9rMY+9WLBJDrkGkl
IyV5adqXFSOTYRbZoTfOAIqt+ed3cvSxAK7dh7azdQ2Lsa5S3PO2Lv201JR5/9SBj2VBRJDTNikf
kZG9hLZjSH/KkeJN6jJX9M5vJxVFGsRiGzS35OreU0+WwohSgStByM1TjOSE6WNVOzhvRGL4RsKE
vw+708vmZTzYf6o1nceURV5PixO1GYKBDfbrWc40zevTonLXBwR5mqO/Siz+QXjHiSGizKFncVFJ
PfDjiHjWv7CA3MWPwQzpMqzdPp2200enm0lMhvDyrRwnFoIBm7nvloswW91mCREmQ2KAfqG/mkKF
YKVm7YcvSR0orvLkm0z3qa/yUnLeq2xkPFRbh94hNU8axLijY+KnzEGhVdYPHwN9WDnyMF5Sm6YY
y23v8MQpLAsfeGxzV64rBcRAXxbBrQiQuGLz3kTlg1dO6z9aRGOA4rBj9EbVAiRsJcEyaKk9BefS
k3iocfktwOzM9JTPfeXyZmSaTFzS3jR4ToC2d6NPsMzUqmDP63K48BlMNd6m8JhOinGdcCoq8xYy
6JOnOzhoQfRKhtHMUqkm32ATaGdXJGdmZSIPJygvqQDsSUk5Ubngln5glmAIpDA7DDDFDQojH//Q
4bgiTUPf+OIAKM/YevivMzrthCuY2n7Syumo2g1lkjnDwJxUfE2HgN9Y4uZjtQSXazV5OZ1t6YIR
nVLd+MdhLSM3m6ZgAayBCoh7GkDTflCYk6lum4NG54DyU0IBXwwheov9fUTjufykGaA1Aj+qIw1Q
TcYTv/nnK37KIlzf+/NabdyS3oY1S81HNpeMPzc6lso36C+KswWrT0tVOfjyKCuu026J1uZa6Nbq
qEbS2QQZMA15lime0V4z3YNE/lhDz8M7m9GSBMDPweA+uXRGhqMACqWSWlQG11oMImF0EwT6geKx
qqCHsXEe1jwuvqy1iIC6AB778u4ubJ7AP2Zs5cYNC5q3eCUcAmS5omO0f3h557NXVKqhNjcFcucL
VC2Vl8VB7xfmR04koHWCl6+v/yFu9nvGpEJmOH7//EWS88U/rCnV7oEzhxA2Li3gs72K1Zl+RdHg
xuTtYZPDu6jg12zFp2q3T+Cqs1t79QiWCWPeoNdZinEIKtsKGnQFoVubKJ6CZL6ng+VqOWveARnZ
Y08draxMMK9M0cbvRRCV3sY+DlI4HCCrDNGBE+Wxq2a6V1AQDofjOHctrLS0QpRruKNmQ2cDZE8S
hOXYFvUEsKyBIbwb1k1m0ox8OCxK2YpVeJkFTjOBMgJ2EawpOFloClthylp+W4KOdvSECvzD6M6c
A7GFih6SmRX3QJ3feMx7jFGHaOTiTq7KbLGH7BuQ1l+oUbrbeDq72SLTO0eII0xfa4Af+hrt0m8/
M5LC+q+uWBCi+o6o0ovyfwAz7CI2e0O1vp2mIWwgSDK6IS5AU+7m+eVkpq3+XKsvtz79bAmbZqOd
RLvOiNWvnM3fOE3PmWV3xTHnVCwWlUrITR5YNUpt2xW1K3FP5BxrbFANxNszD72pryfR+PJeLeQL
IWXAMmTV0M3NxIUy70bJP6Z6JsTi2VBP5ZbyKvYl2yPG3oH0ykXCqfCfK3FyhX0Q458rUkwQdakb
DDRv5w1jxFqNEyHwFoQ2Usm70kcTFa3EuQ6QyAiSblpV3yj/kRuVsDek6gvJqoZuH6HMoy5UjHaG
5L6GLE6GLjyf2KezypjE5VxOizQsoMyRSniZ6l0W6Z0nbvCkLN09MjkUMRiLsF7F7qsAqToq7RI1
ViDETUUhnics/F6KYw2gKUo5XcJw/MfbzZP1xIl4KakGEc9FPHue4CNAiwFKgqgdXr4PBh62c/3n
UDEnxv4qJ+H+l9llUfzMyglvw5PV8eFF/0dAsl2Hx8ojHQGzPGPs7rZ0O8I3ZCOL9yfaB/BkZrjN
/NF7f4Kc3s8Xlj+W++1zRXm/hFEyNCAFR3odyToINudCgZLwXpM53bv9h6sc7/KEG9R5smXl9CUt
AzWTwzhmf07DxqXEie0XUJ2QuP+k755b/KD2rWSSOeWUHYs+Vmc1rm5ySpbOFkL6Cx7bIyClABx3
gPsQNnj7hbbyopqNcWAT1Mi6GeKpvJXvlpQ7VQXSuYzPz9SFjdkWF3zXVxB1AXFxp3iFRCJc9CkE
bBJ8xZXA3j2+OZGw86ZhJs+Me5gOGVwHzsADE83SeMf+CYCbV193mBgq5KoIFSWynf5lDDYbNnc1
dbhHylKX3uChN4fFQjUIQ1QGUc9GMc9ylxhbdm0KUqDFBQ5hNum6XpVbz/VTzYNFmL0fdO/QgXzI
bgVWjT95LD2JYXmyDaip6N93i7lbl6o0pK0l5d2f2qSXksabGcAhaJcGeDXG/Z7+ZQhpkyVXgI8x
Nt3QQq4b57QRj7VWbxGqjMos8E0EBEvuz9N1m6u+tDwtVr+JlbljDmRYH1uK+FyWkRMCBuEo6VST
Nu6+kWHOXd2Lbv3tSX+WM5odG7qrmXRpfDEIaFiYCEG/LQS8ayPnQU5FhiZFY3qd/ddWjo7wE5uD
+oAXNpV4s3RszkhZ3IdJBVOHPkk6/OkG9fhfk2HChFDjqhHUEmkKnsqi9AgySBUAAZ4T7cqPm/tc
I1qyuouSNOjgoHEHgJCo/HvyG0HlmI/hH8sq4jsaM1TxJzZfca9kIvem9PR7mjuwikaqvljEcMRO
Xd2mx0U8Qn8Vbc4+MD8oSe9HzJ/IcZ0HmmlLDmtVj4KO34rBOJPSrUHnZIAzPpyCa+pjH4yCUcze
4/fuFLzEtJLsb7BIyXNeUWPlvzgIC+3Et3G/Htt/22jESWFbcOIIvfiV3IQ9MwQ4mePSV1eIKmkr
davHq4cBEMlqcXBsKesZhepDOmoGGF+ksmtQQRB3nBbylrHJo1J2gI2HHgCXV7tifxEhl4DDeihQ
mzv3x81zuQcDuZc2rr56P8MmgYqMY1kFx28uFtRC+cqDxobdkCXLqiSqUxxSt/SPrpuNbYM0aNp9
PfiDCOePvwIjny03uoZhJxzOydjjihS25jfBXHJEAET5e3HFJMce2+SkwDUaLlNQoZAruoA10121
rf/4dwBno/wyiceKmtwefjcKoGYkWD3dUtVLPu8K1thgK4XfDZhRe01bPo04nJ3z2Y6M/lW0c3We
W8QiAYZkt6/2jXUj3pBPk5bRGM6HMQxsqDSLVEbAxDzB7nfV9vrnTo4S6WVyJIkkAJbkLINjXEI/
qNMkrkH5ttobUrZnx/hhAjvE+C8KHPbKVXJtV6EpKOmz1nZhAK6OzsDpzE3V6AS1bpbAfyXB8Ag0
r1xX3t1SrHTyFUxibvyUipK0TRlx0yx2H1UqJq28He1glltNcOVpsnAVGPHSCY6II9Ex0zGg/lF0
YZ2299eetskRnAcCAmeR0QIBnZD+6gtUprvEif8U0qvYxzmIDIt7+m5URVD1kRtH4Jfy6htLtIda
QUEnf0Pbo4+Fr/ccToIhcYkzNauH45Xr9JH2cxqJF0Nt1QeiJNstQgvpwo+KRsFK5U3RiuCJvx51
Uttxs9m8csS5EaohI7kmhBWfjYRr9VMk3a+7x3QOmur5qcpIe3AuQvjOmt40tDf+tVA5QH2fqlQm
6iy8PgVCXI9GQS2L/arbUvpNgF3MV9xamfH+cZB2smOXwH/SmmFo3vEM9cb5CBXQFY9ktxqhMyD2
ENRx2JY4ETM36amlJRmDMdN2PlMVuakwdyHdzyzGFBHuCqGfZDcLI5CNQX1GrLlynuqqceMjLn2Q
9Aqm6GKxOvvXR8mcRiObTeglkjckPA5HDK8zfJ9xDfTj3GKl4t7z0K56owkJsjfFX5YA07qlwvQx
MpFriWvCv0PxYY7/0OAhLEcuU3siIf4L+eOeAXqiHaybGzXuhOG9aVivn6G5rtQJkwJ2l5LuSEow
6/ScakC4/6gkYEGWPGc87024HqyhSFLLRY6ZUyENUWPelCWEG8dMpS1If9PALlfYM+R0eyE677IQ
fYnqlqEA7yP1sv9ToyRTc/iUyhSSjIixentKtzdVQ//wkhncmyQvdulsnuN+zCxCvXlqaiAOXeMM
iYkL4E6olgjY711CrsCyLP26z2cOqw+awwdWtnP68qTRV8p5igtw5UZF7DFvwu/XcafA1A7EBtVY
sJqF/mwSaZHqCUJ5pzqMEqlESyzuK8YUtC0vCKNzet0t/Af0MOoLzBg9gaWk6gL853ssfkiXjg6u
6sctEt4pLpKJU7kl/0ZcYd89b214EewPsRm71bs/+Ur+sYGT/58XSwCmbU+jtQte2OW3GeffsnBK
j/8TQnIvIIDPj0r7jSFgC5mhZakvZGUhy4u3jLoW03yZjMQyDypq+0QecQMgJl5cLOmMbR4M+t3t
4dKXFxrbDWXo0Q7JYrZOnHYGIQL4tYitnRIQn39au7sfmqanF4KYwu5rqy/GILlVLNYyRdqpWeQa
UE4s7QldLlmkQ4nZSfO0OziaA6qzpy9A8v/z4YFB2+E4l4mqvb9qSrMPcv6Asc9YdKRANyIEogpB
uJBl+s/B3OmAMwVOLmMc2REpANGs2QHTr5LId/yD/hm71FvjAN+SHczyux0L3UsHvyd0UiFloDbO
XeaPNQygab+4op/bkBCTQuW0NeL3Nxjvg+w3b6Mu6fUv3U/R/QyeOpJpOgwIKkiJWvJSuaV7kHQ+
o2g5/O2+PUdkeOBy1cHZ+ik/XHktkR5qnwx23VMDxdpiqhm+qfr2XQW2cKH9OWE34ZwfB2GL1ezK
XnkMwBHLZOChTKFeGyI8INrT7hnOgArxxkuhxjJC8FGVSxxDYpyUzHh28XYeYeSJOv7aBEdV4mzd
xOw1Vjz0xZycEimlLUxLAHaoiD3eo38+XVAtPFVnMEAYvuXu4NL4bWTrFhczp+2guVUHeSeXVlSt
GZesugdQh9D5dwfdhWeELxqdaxSLoSNXgPuEuAtZ4VvFmmelRU76oXuLVOKBK0dCgcVEDWh2nd59
CEtiE1exDWOtI45g0g4entllKTnBFYPH9hPPT7ZYkcd08/4IOySyEpWT/P+yjdvMWgGaWPMhRDal
2xrRh8x4b+Ck0TgQjTdIqdVFguo4dDbfQo3+QiFIqTuh1xHk1Qkva2pMUfGmVYxmJ5h02peMaYqy
J4Fq8N74vAiA4Ti9YSLOemvh8RRyxO4qmOCwYd1Z402ArvT3D979ao14iEMj+4Qz66pK0+68XG6n
eUl3ByPDe9rM3PIydoo6ZZCAxB7kS5P2IcALlEeRtKXUPYzdk1i6hZ1+EXsyirOaV+CvftVNiEU4
56FXhzszN+z/Tp4AhyDDzOYdgx0X7Mv1hZqLnqXs2twQ72jv+KHBPQVKAaOTnc9grxIYTR5V8l/I
pSsJdCkQoeQ8MgwYpiGQeQjz20DqTZ4gaZqN4rJhHbgmnb6CRYo5XM2o1zfJwTcGlAewxQHTkZTx
Lh53J7A2g7dVAkTPdh62LVjXvtCHtRV7SpHr2S05Sjly8MyCq41FZdEnyg6oiMNX4m9kmocDIrrD
UsVl/XimX/blRyP7ZOazPRsHKwtX3+vYdt1jMSxwUlfVbtDgFTj6JslGOjXcHHxFAQom+MNezbWX
EwlP5GTufv7WfCSHj+W1gjNskxbHa5XN62QDuYB/JjTpoWkjlsRUjzRwWL76B4iZHXbMzKD2znTb
tInOpVZzG9fPDuYAM+9Rsx1RKH+3br+Ca1LqASo1FouKLP1wsv7QptCmBd7Zb9E/3uhSLGUWtUJQ
0XHXJI/q2fwwXQvG3/HGVSNzzAJTnrDMVoW27Fc4VpfFWAbq1M0ncwo9lzK7xrYR0lvZdSr+gpvz
lQxFC7HldlBw1eBfvupGA6Cc631dqCDiPTRXQw78hkEUHtzZi9EEusjthfn1YBTbdO3sbj7uV4c0
+E4u/hz4PoPdAkErbGpBeZOaoW+lc+FVWGtzm1EchOeXyvh6k7qropdMZkx2cS5NjinuSAlxioVH
IDRdsyeHQojuHVKVLtaWGVSfVkaDjNQzumjEdIDYgkuw+eIIthcDoWNUnDyK3AiyseVPoQdw4J/i
6JEJvfHPsjXUcZS0N7lOdkCduVkfsK4/XHx4jr9fmBwr0tAA1YiBvPxmOpeSbVsVfsCfAvtiO/TG
AsJLqMr2L/H1zU+Op6mLnx/gGvH2kJtL5EEsZRy2y1deRwjFljnStViAOIZ/7HUE/3yRSEnBRUDq
p8D8ZiOuV18qvnA0e+u+VTdTCOx8pWACkhrGqEzH6WipBdEhDqirME983X5/dvX11LjnPhS/iaRt
nsT+PqDkJEdT6zSJY9hcGQ8zlJCG40dTimMYtl5INNwfIKEYr0YTePMM4BcAkkpBjQL79XyvQt5D
fOYB+uXIgCM1/fVY/EZhnQuXYBgkDl8vUCzzb/hx++0ZKlw7NVA27D3iT/8PBuhWO3FDNi9BkT2S
z4HcCSoklRlscCxlH1k7aMOTGVRVxP68/svrKo/Do6JtPK8KmVQd32gaK71EABb2krROHCY0l2b9
IbuetqeqMB0rK7pUPSlew1yZY3uWuFrsaUU9hUhL/hJIi7ffH0hIaH2SM7svCQpDEFPYQ9wZuioH
efony7X5ZMppEfqMqh/h6iANq2ylG7PWXpZOlCco65In0WGQn769YHh8uDzBNI9f2LI0zqjKLmGZ
8Jxm5+ArQ/gvp0LSIvFJ9TZUIS2Q+4a3sCXLBNjd3w/lPS1HLBX4dHeH9fXxELVH7dlsuQA/wzln
tWcsO1MHlwVPqmYM3QZ+RrKOf6T8AB9BOiMM5h1tZtrk3R8AXzqQa8V0VwIzsR/AN2Bx7xABbyBu
m4xxsJNQjpzwcU1zk0hgMTyJ1nyy723H8AZtenZS6UNSi6YHrQkwSl5ELEizfTdWy4Ry6BsQf01Q
ho42hoZztsIUBFqYG/BD/lZ0cwkNZJt/kgbyOaWNIi1AtHWERHhk0AxxY1jYv1KEl9ngV+5w1BVe
hruUzpaCDdTGdPwOsoVq+dVCY9cPdcUTOmhQYV1BFoHACC6ajDvEXYp6N4ikqBVbcKfcPeUtDNd7
BxRJ+voTkXC5vlmSSFp285r2b6I7DPqJpGaR2Wx994XR/x7WzxsZaO8nJMKTEdiCLPy/OJreVz0g
tItxJpK+vrlACnkAeiYOuMkeh/MM6Y9lH/m7XsYwItDynWkZEdxVjcUptNlS+EgGPBE4vrn9OTZ7
W7B7c9tmENeXVzbE1XzNqdgwvZo5cI9wtwrmnMIL68tUtjupqdCAsZU33ayKMPbeEviEk0p3V2wv
nn4N2/i6Hky9gC54li8nS7TqYxBww//iBMMsoxQSDUBXUuJ/EXH4IMTFZGh0hyCu1iDWFZAPwDw5
sLKJzXzJousf7a1qPY/QAoHYo9kSZxKWFCq2StEIK5sAg9QD8QLqCCWnlTd3lFZ40+dC1T3pUIK7
e+5M2DxCWxQRjYiUvrEALgfnAej7P9HXmYWWB/4S9mnZi0kmTpdgQfRf4rhtvr4FNSvpI452+ryM
fCwygFVOfwunqG1BIw5XRmrcshAPeYENjes/lX1qJIrQc7rWAIW4RVsOOOC7y+0q5PxVgNfTdqRY
PLmKFebSXqqeZz7TZLIzjmI5dQpYDpkSKHGdgrZ9ZLf5GFLgZOLXDMvWOzOrap4raIB8LxCUu9M9
M/uBq5eaz38jhwV42FoGFgnjpcGfhHEeeL9zszUmloq0WPaYwV0a9jTnsM1sS7k/JpnnHQ9Nkd3G
nwoWI/RNfQhIJQ7ceLJAPFz/mG8MCcZ5jRwQqAQ7PpROoyrTQYC2E7CReU9Pelhm/I9yCKOoV+sc
FYWZ6IJZnZaQ0aiosY/1Hscp/bMhBGoJf2ggUw0xlvMUVONlOT+nACvi8SoF/4X8cXH8yfScy0ba
2XJRz9Kpe/lO8ZMBVb/ZRDbbDv3szNVMQgERt9qGi7A2OEM/mMDEJODe9CqnAt+sdbZAgYGlKnOj
MXhg4hi3HoF1pQioLqFu0EHhBn2A7MEpsCMz51NJmF54+ISzeb+fCD92GH399Qn7/6muPbsF8n8n
0hm7H0YM+wrv63d9goxQeMVdLqN9PNgqASC/ZS3n6yCMqnNT4vYhRusdu1W5iIDZTnSc/8N3LgOY
0GrSRDORcYxTYvQAmfPNi/Fk7bkhSPfPT/zr6oNAMSfm8fcgaxbu4EovqxYNN6SDQPsgVn019ntH
q8sfL4ZkltmNivJFB8+Ygxf4Hct4WsfNPtXClGAkCeIIQ9SAet+SVO/i0GGMxpVuVIjmqiuPO0Ou
7RZdhLgmsnk4uKDFirT+CpMP9Fqtcgxfn/SXnLuFrHuo1Le3cigsCBmbkZBh6g4tiOKGvUTAQwU2
L2n7gFzW8Mf872NFAVW2igLGzMP0O8Vrat54xaWSXv1botpobDFSQ6ETpDCd+o6bKI4nbUGu4w3G
fbhep6kfzehkjSPgEfNT/KvZDM+eFYwpeq57hWeSFZ9iYUw87iV8Ym9AnopKqovRZZHoQxsMEGvv
3AbBxmCaHbgTkRv+mwU3MubCdVlK0lTzkt+zkCyTZUdCsJ6Zq5iw/GcwWjVVY/5qx6G8k1IdpGcM
IaM1wtfkqHZQl44Mktbb77ur1B17foDqjLuQg52Pr0mNZCM0jMsA23/YYKzMlRXQOpyueLqoxjPq
pbtRFQPYU4c14/2oTj4/VyhhGRWYZl0nvYs851WRmbZXUnulhVuQMtB1TzjSn5L7MAuK+OgrzFlp
FL/HSpvVP6sNfwRhzgesYuyDqWJ7RMv/J0qL4cTBCvGDlSvhsYOqWz0xti8uHzP9dwIxQMhMvnok
ZcpZauz0OvpMc17AjqNu6K8Mm/bDL4ejY3r4BbWf7UbwVE7vRucfrE+X6mg71wWLk7TA7rJWItB2
tXYRDt5FLDaLCvlxGB8HoePyM8spY+BF8Mbqnu80lCsugPBxXDOM6TGsLuyUASbbD8bu1UN+TwB8
zHEnqKEQVbo/DoDYmmWby0aP1r4HREq9rs9RzfrgYHwm8Gy/i0FBPi3XhD5l4n/nkHw/KC82smfn
lY9PefO39SCnd4iMBlUZstGXMOCISPo5kFEX8hEBefJnNCGl34eHfvJBADnr4T+VnxA4kAYWRFkF
tp4eMW+OnQsx0WRyY89FF/hLHEYGJYZzs9nouBgvPOA1pjvYGBPSbPekiu9f/cvRor2i5HlFV8mq
atjAHz2NwyqUprKoG7AClLIIL+WsHWOZQirK7QnaTMO9WCcCGhTtakiqubYrfC/nUHKx+9TU9dDX
59sl485ast/w4MrcIAm2UMYNP8kIifyqWOeeBYeQZWw35mRJGdilk3vnnVaucoedphwr0sEi2Bpp
+ZzsHDiRshXjrB5HEGMYHx27VzB223LsKmRSqEVQicl72OKyUyT0H02eY4GBYOTR6BfPrrSTIqMK
4e+6fx8IGayR0Fswl1rrhqAkVdUaUtfwUx4cTQr66awti2ER6MmlMuBLfz+Fu635Kc3o5dR7+gfx
wJhR8l8RRU0wbRQORXbPUo12m48vc/CCSZsoez3/HxXWhz8CGOuhm9i6yenz45nReUs5KiJZ9Oao
qQdI6jgu8ysPkms+tw5l1Rrqj4v4imARKMWFOO0OzzUi0fZRfSvoyQ6FZVLOpi92y6MPcP0asWdD
Lcm+OUwR2Z7+DbOyMsylKh96i0ZAY2P/VrShxLn0VOs1zDiesouh7QU0KFmaZ91trhL+FQV3H2Y3
sT26d/rWSniWdV1/Nyr8KpW8byaADPHFs7TdS7Rs/qE844iGqw83/gEIozUDU1kJ8z120Ue63uPz
Nlcx7ty/EHcP16fgy6J8k0slQedEqvQAtJMw91rzx1Rwv7QI+QfTBgUgphVgtbir9i+9C3g6x3Vn
W1aaqaQsH3+vbgUCYOBse8FF3etWl2jNDm+igcy18wjtzOG3f+1DlSkvrG7K0fBHCupqwzXUgXGz
815MxiLf7DXNnQC6q3lVy0YYex/EcbceFwmG7vQm6hUQSOfFnvaHsEwGVpuR9z0w3BOYfSmS7qrF
pZBdDxAc7QSz5RKtqqiywGPpyjqFOuHYNdDYoxZLAa2gGuLI93cwxQjtco1q70tKAEsLKAVQaXYn
N/BCDNjZkYD/htNyMQPowGGQ/ER/YQStiI8cC1p0/k5CWTx2N5qVDOc+elVx88Pyi9sZTF9GcImW
HfPrTVMEZO8QyrIMJLTGGizka9JqDCcc6tLoHkGtWdIkAoeTKnKagwwKjxS8yjMUZHOhCVS4E2UA
iYeyiCbn5sjoWibT03syQxHSgSGStvRgZhJNRaGdCWnJT45nnz0rCWUyy9lAdTfD3x/rnv8xVnjM
SXO4WR+uKMaeqfEJaSGxEiQ5gXA68+bj7GLpdlo0fYsXbc9Heg8Kou3zh9gyINh8Ywuk8YBwLCFi
Nn/CP6ZIUqzEE820mZInlCE8bAT9bF5ZhrlpMR6xt6iIvldXmX6b2aGG4YirXeV7amcoWjTWf3Ob
xyN5vWDLx4Hiv5ohRgKu10Y/OQNbc78CvTCqMkhwGArlu2tq8pUJHKPY3zeud8Z/85CtH8WVHGKr
Q0GwOB/WG6EYe9Ar3gcCSjOVgW/eHc1XP6hWzyBUcNtfkxIWJ6VlxCzMDbWQrhDAEJ3492lhaxD1
eTKre6wenET8ndBsHfOgoJlUa27WrmTk5cza9Md8UQNGfw0bIe8BgU1iS9Cv7ht7OqNUwMo3VmIq
V7x4f9ua8aZUpbGjpgfA2zqBeO4SB3Zb7zV7nRe1Ys9hTWKHpYqry6iyW9Su2hsYSjq5i2xDBPfS
E63NF41Odd9qIPQ+3GU7sYV9neC+GI7xMPvLWavxXog30OD0aVfXuSQRtduLbflaBkvLeOXdPpOR
ZzlyhYKA2fL/69TTW3p1l4HNHKbEGZoJDX90MVeqZ95JnG6P0JEbGBjV//Pv6ffw6MYlZDa5hIQl
3KJlHTgMjMNA7C5flrgA+scBjIWbxWKCaQ4RWjoCW8YbjGwMVyfYmQqQwWK6DZsjVk5+BWVuqAfb
bpDATWELOV1CmF2VZs8TB7QmJEiLcSvw7ZImrGCGuQhHvaalku3hEtlhJpO15RKkPSJEzpivYT2C
KkWjCoGsXorVapVIWPk3GqGwhfqyHsvebSZIHjrFbErdEjF+KheQpOB/3koOAL/D+QMPzcqOCLQn
af+sS9c6tKbGo9Zevv0+SR9bMCnkeMXu/UQQPpJ3a6LQsvet/92wGbCCHPc/P2kFMWvN+g2t1ZGj
FYc1F97aBnKJghiXWjXORsX2nNx4U2ZQAAfjktglI9ZTf+dVjW6DBHTZvDul9brqhlZcD/xPaDwu
gHGujQ5BoQZB2Mxk/F3qxTNvJ+eyxC3EK7xEKBT+AztLi8t0LSCEEIrODwuQ8BwxF5Xe2aW+ZNeR
Fk3nVxYI1Iufl92MPUz0SJVpmjJBpiuEbgQ98ih4K5NtPQzk44MddJTnA3ve2TRczW+jVUFDm0gO
ZHVqinTlWp4x97L9/VlEmULjgVPpHpDvfqJIMFkbnnDFVwg0Fcy/2ibPdGIpGZEYf/UUViHfCKeX
UULgHgofxQy5y+/f0ARhaUK77KE8OrG4q2Iw4EUMZqcT/oREecSttKP60QsJVK52A+jOQAAhESw+
N4QFdg2u4DmkskfGY5IurzoLKWp+Rxpg/zJL4HRgShZ2Slc0O9AeqS5mk71XnPppDcXY9LPsxVUo
Gspvi5rnGhW4zQgPTkRzJ9jLkYVWxJJRmqa2pVRcQjF/ZXuqAEgRYxsafd6u1sZZMR5VAtEkoMIp
mVLTCZ0vci31EhHphD9WcFTVDha+dqX6359b9BqQQBwDUB8kaVSQGJhmDPNnjSODG3IPsZg/r9Dl
4h4IVQ4qYkjEXZ7cpPb5ktYBbTGG5/EAVAfhah0ko+ETjpRzJkQNwZa3a7n4DxjCRvTKZGDvxAzP
DnFmon0bo+g2kvShFmZJYQJeF5G+cnpe9ahEslApJftJBoxBvlUSf8XkkNlIW+t9uut+7QHUBBda
+zqoW8nA8BVfDEM/PTRdz01ucUMB/vBru0ofIYVCMBlTRPdbdaGJ1jr/WTSydcD2g7cwQhb6i0gh
QCJOnUtr+UxFVQjnDjIF65pYDbvFQ4AFnfnCkPSvxiCsQ53JFOIzFQY8lYLT2ag9GdO1bz2lW2Ek
d9LHDu2jl3nH1KvpLx7R9qK3EZys7XSG84GHupO2V6yDXTsNSctzPEBNjUj6jHm6cGgF/Bgj/T4a
ReXGsGCX3VO2bpi2GtvbQcNT8fvDm8/h7ouhMhCL7ZXaXO/znKz4frGI5OQUpNSPbSNN/Kz9geW8
X2amRPXo5e+u0h12pS9vPYcTjNC0YwtwYuibiineZgqIhquT1BpupW125TRhQg8VFDspUauJJpVo
BtWudOY9qHzruV50RQPs96DUtUpsgbSW+P+Ck7enOKAs6P7UV8Og4pOuBNRluxwyE3G4kwltijf5
WXZZnItW4bntZ3hiQagtHl2axHVaWk43+SAklV/wRL2ALdWedyg/mhyxeqfLcgHneFnxSRKr+1bB
A1g6ohwwNm1oEvc6Y0gbD+a3d8f7qsV4hay6bctIChg1iIrLQJPNuIKr+mLuA88mvCMtXE0AHmlu
jdQ7CX/zDo63GNbZeRS9ux8wgFcQY7X78SXD3Q7/eJNlixdIjG8wJjdyCDD2tqSN7/+105A5WcY8
drxUITqv9Mtij7qUhO5g797/9IQeRAXaVSPtXqQl00Mv8+5dC3VJj3N3QdiBLHt2k5jTJMYEMvMD
uxoGcKjni+7BmZimZ47X0akH/H2mKzU5eu3+lGrOAD6dXTC6is1TZXOWz2H42jbPw33natVAiDzH
ArXIyz+CnmVxXkXgbzDcebbauL7G4Dl/KttLsvbNPE5QNn9sEGcoRXS588JaDTVm5+OZNiuw7Spe
gNhFBTXh0u1DOlkA5YV0zxuLV5u66mYEVbfr60XnD9NVqYLWmRmmNUsJ8cXq0OPlwSA40r/574a0
5Lipj1tchXHt4sUG8rSR+HlebEqoG2LLDFRtf4hqrFjcqFSNr4l3TgPEEpcg5zNtQXmvdYMVXTxd
i0Iaysn6R/r94uQXlzUDJGX3Q7dGpNJ4BiQqfBxbi1TvKUcAvE0izgK4AyY/OK5MvYG1cA/ebXtD
UWyoxOIYn8I7UuC/MlOyo7eeS3cNaRb/n6sGi3rR3kDYXlks1CS1qVqraPRQUtgqs6SDB4Fmm59l
hy9pzv+SRVTHc0/D3yI17LCkyS3u3KoOByGt+TsvCYgPL8KhklDZOLZV9hwOJroSdT7Uv40+3TCZ
nft5dvFf5Firs1l8R0hjhrDDhxpSTqHM3o+aiw86fXnJ3fygnxT/at8WMX70qIBtzs9zTZAvi9cF
vJhc170m7LNgnIKgvH0AYAiUEM7sWum3YJbRJ1MnVdD3/sVTQzBaWDbhXTINadqH342yXxV1huyu
pTnfdSJiW63V6UXpdwq3vatLMVmfqobp6eGXzRLQEipylgIDJ33WYRMGmyNsDx/Nm4c8pOLhVmSY
d88JrmUtVGda7maCrWm8eVHu+IMXe6srpF2whGBZy9IJNbCHxgWLqUcJaWrDctNV+09wCbO/LdMS
fIsQsmfvwKcu+PnVon/C2tlP2mdKSpo5tiRlLQ1oYC0TT2QAyPjfUdvM+wZZOABbSPn/HKLlDM4/
AmsUzIwFCI0e/na0/m6ysKoxyGXu1bctE9sNDVuFtO0ebZfTxIJ31enBk/YTnkTlluqrw2i490ai
8eBYy7pqmclLeWNCVykCCty2ktQbauBb7fKav8ed0vWv59rYsbZkSiP64xWOXxPBO6IalBBWfCxx
o6in6E4WaeXTolMl1iMO/84t6WRxNnJ1HVwzlbGi/w/iCOQWUdW0dYr/zUkd6BO4TdtuZAkg//cz
Z67d9S6lY+gmw3LTVeAFHRFzF6rZAvxzeYn/KQp2yPmuQE4RzOJk6Yqgf1pSXR1wqWAqWgfYjjHs
SCQx+O4WFANzYhgbz3B1OwX49iUsJyq3ojwmF/UUP/5jhi93YzDbF9UhTJoyrpg0X/Zkt/2iLLem
FOYpEm3J4VdNWLmUZeChQ4SxRCRF5jYT2hgaOoH2Q0l3Yz012LZaa5Lv4u8NjhTNU47APSD2liXY
lxfKS58PkoViweAkJn/jYYv6rgQ1L7Gu4SGaDw2spmj0YjrNPY0x80AVEH6lixIgBTnFR72+bmR/
23GsgqhxfkFa8Ftm5ysnjl+94I2UBScZVCgDmcRTYUpyri8ghXTpq2OOxJZdR3RL9V3ma/5VGqrm
ro59iAAraZvnTAAzJbdffgetcQsjG8Dckl4p6U74Wrr6/8VTc2IqCoa9z0dxT0lRxGQwAAwvnQTB
+/9pGpvxLeBaQHyHhfCRfbK823K9ENyQUjS0bheWNUBXGh9hNMuADlvDXCNbegV5dsSAKqhEPyEo
zuRVAT7CDtXdLZGlWgAiMxDmRz9bXYcNu4lQ2a4hxPN4/P9SEnMpfn2PtvJcH9QGXOitbdrAItZv
BLP/jeQ2kWiiO9yuGPCsScQssi3T9MPVVo1jvXi4olvd39C02JM+z0+6Dopjuz7RO49uZwt3qXUd
reJJYa/IN1aJJgbeYBTdSZigbMu8sFuj4zEdXY/vHOqLFUZI3c1ZqMERolD6b4Slcj/RwurII2St
xMhpDso/hZ3FST9pxzYxc57Dtmf9jzLs6aJwxMf1vUQbKugGQE+FaftNSGQM02xGwfDHi5C7rpat
JLwxIV1ZliE52UtCwb4gpX9LBtpolriASIu/r4o9xPglS/Lng0fTy6RWVkgJKcHShqUISPufgPo5
PJhIOr9xbKFGuh0kX4cb/vRoeO71fAnU1A2j64irYvpC8BW4Dtdy3N3CW5bu16Ca416n8GfpaEl/
TIwr5N+QxjORkFWoYkIGoeHNKRuSjIkP+2ZPw6kmsZVQicTLo80gFvEeKuughl+4of31XTIfpsUs
DiA5apaVsYpv4N2CrcMyFNl/wb5g6FoKuJNlgtMRozIbtWZlHVbh1KdoRSHrFZEU05jzd5zmJtvW
9pLLM09eacG0YOMQMdIAdFRGDBXSnOk5Yjvr3U4InvnOthsQmkmXX8E6NLdtm/uZNH5dli43ZnSp
vzZ8gs9sfrFQ8qXFFUJ7ynFj8xOsjUPpuYZy5yfZ2CMtsih+Vl2YWhXO4THbBFz4H4elc9GoXXIB
HVNsMZ58OayfvhGJmtsqAUfOeJdg+XUwDs9BKVW454zy6e047MU+/9lU+Rt9ic7n3fLO7tvN8F88
ieyuYlhGrjL0ZHfX1EOlYgwXKJybx9p9CKpm7O6NaXsZX5AoQnb5nrbtbRqi8M1Jlh+BwmZHJRmB
st76n+oB+vk9r5aTxibqfvIREZ7lVdZhtqSUzgGsvzKOePXTpDTjWhHQjdBO7vA0nQt2OvPmIlvb
rE7qgq8RP19b1is9L+uwc48/PhN+MqtJVwDFhfK56gR8shoSU9wPXZkagBfZWfnNOJ5Wa8vgbV5T
ju1JAwSKYMTr5AUmBXg5TXubFbFpAh1Mg4X8w1HiYk5qnJohjrKOM81dJfSZ0smnvlzpJmIzQzFa
sVnAZ+6d0toYiwUATnH75aqMSzgGdXMjn+mSinSbPUGO2QdX04HUeHuBJLDTqcSucSMnC0ViG3IP
gglG47XH3YE2sYHeEzoYhAcSPIPBf+7D/AFWrCPZYFAA3oW70hWxaBcnKsEhrgUVIK3c+HGJomHz
CJVfxejLWXzxvS5FCQU5M5RV+yHlbs/WNU58fjO2o8uvMbwHS71AXlWCXZb1/vvMsrH2wdYqrMIa
h3tcBGRxI7puLUhI4yGK+8EO7GRET39wjJbezSHKwkQl1n4Xo8nYalmN6IxIGn9qWM4A23+Fodfk
4TV4bfK73AG3FV08r6NxQTHVIsAMkevakSc6zLZEXTpLmJNbEadeocPOsBdwbk4V1dOfPsIKZ9Yp
tzE/0+48CBcP6tYvazl+2No2higtdRdQ/msdUa1TCwqmq+aM6CKoR9paKQDGL/vlkgg1l41xIFxR
jU/fBMdSMUfMWPZdtaj+P0lIbIxu0KzCC/xyAUnVliFjej3cXXgQV1MIVrS9ZFcIwHAGEcwUafFt
b1w69thdjsOHNVPsAnj3vtHMWJOc91+vmj0b2t8CByd+Axn501gz9LCESA+MG/bqI4x3l6rrXfHf
zOy+o5Zl47KaFRSUFmx0npVRc/BKKK7VemJgQupDx0k0ZEabQSLBwFORT0f0DT8g+qAuJn5z9H34
CPMGLGbFUCN7uW9kcn1fA+8uiNtOCtfuqJEHbSQZws7UDnoXTKUm9v/Sp0KkcF6W9AiKWvcJa5Wh
EMRIx4p92AGHkmwp5wthD7ivHjTwZd3GVk4tM3jwHuLVhy2n0d6ezqVk5bNMOHoXBhx4FVd5TCzx
zQ9xN8OJfkz9i0Z9ztvnhAbXGf6cVSxZtpikd8xRDnbp5P2mjkR7hNJqWXaTjFJY5mKVDx+F/o32
MXoKF55zwkA97sl3wwUOZTGNwj4nUS2XbsRwAzwIma+znHcJ+femzz1+UQbaUvfY0QegbpmMPXVc
Ya0PKJeIagqg27xsA6gAw5Ih9HCebVQRq6eTcrCJd1V7Sz3RLVQ7q64jvSiseRouwlFSpkYRLLpw
3bCba/Lp3MxYiqq9ud+ttoBS0EzR08jLoJCPQBhLhJm2gsj32t4ULeESB19WkffJZKqlEB323gVF
ujsR7p0Ak5E7/CNBdKt945syUG+C51/susGG8M6/L4T2z3apleeXi3pU6fprJ7ZjuN8F3bzzwIfD
9DgAOxeiCDWffiEQwcAK3jVypY6hFTiP8OPFiaPcH37iNtJoK5x26oC4c5gbMvS9ZhN+HEbqBlp/
/xtmPY4qeTgZtT+mNEi4j+0RR4yhBpZN8URfC7L8uKXBB2ssF9q7ntQ+vWaCqfCi2o0IoJgZaBFn
0Lgg++PhmiFk5BlXPgGMPcaI7Ngb5z/4fOiTMSNw968qZrs2qOPOZQlAfZ/IERisUrqKye7kweYz
QlVQQmGG3Nqcbf2TOslZHlW6qLnnX5FrDATZjqEJd7G992JvORYYmHIEQ8gq8gGZfflhSW/crOgU
0IbjxbIYHDbsedNstevCpRVMdxJJkqmyRrzXTwISle5+RWqxs4vE0w8yA+iUPHwHRZR3W2iTHfjS
ipLn0ESw6EtAG48dHQPVkEGwaEuPOS3xc4N/blNtEikN91fgGhewfJqdv8DYB78LQcMKDs+c+p34
LEEawQtgw91pvyRkHigCWl01BLzm82/FF+dSpI8WoipFcbjzu7j86y0Rz83D7Dm3G1Szej34xFSh
Vu7tBqvPE6y6nwbJX8ObU3+R6B8oG/K/M9S5BKsehFEGtB3Y9+FdznDfvoh+3RMPtxlKwoIkVu7Z
ZwhfFQvagp3XpXRnJzoHyr2Q2QnaWFN5tdALx+jS1eBQuZQckY3VYP14aivTn3/iOpCqXmSR7L5C
aLS0ePXUTgGgV0z5wEXsG3fqVN3wSUGR9japgY6Vn2fjorPwLetF66r7vzVce4cbBbFoA9JDOXmy
d7BpUC7HAEWKWf8I3YcY3Z/2qy1/FxUBj4itIsuKJJGDUdcJtEisss6Drw7gAIjrhCkD6Qo/EZcb
6OtFr89RTrhWAQuj38/PrPm1zU1eYcChllEZo51seFzThIbihfBueoFf4VaEj+FoBrlmF3y5Vigh
6mgkgDagLtq0YURKJHOkc0uYzQ6RTyrgCdnv92DLzuVuM9mmZvS5eAX9xb6c6C0JCEPklKk68nxb
rU6ybOvIdqXvPmfHrm2SVhi+Hr3oCVAcsFqflcrSs2fNdc6pf3E8rO7HXcyFXl5rqS5ms57js2NS
ic2CZaze8Awc0YS8kToTixFWNKe1Yv6JD4jJJwZsJ6VMWSUW5NLoWehV3zXZxWEzdBJ0CZNMHuG+
zFy6w3lb0B82ljquDwAv7WlbEz8QY9Z0fq2T+10qC2S3/y37A+W7ZRw3Yh9bcqzUpN4h9cW5TnqM
F9aGhGa2Lfp36kn5mxkvnsAM6qU4Ii5a2MqfKG+AMXa/kmw/lAx7IePdZWFrZLTIKYnRtVXnrLVZ
vwtjU3r48goQNXtMSIz7J8thiHS3hovudDz4gcmp3HzibAAVZ8NazP5LG+RKPSIDLEifUGZB2THO
nlXwA5WiUv7/ib/EbCIdpCF4hATxhsLlx8rSJ8SAS9NAsvZS5N/4qy+UHLORCB4V5aFnb5Uvv6xL
Oq/rgElX0KIY5Jr6jEQ0mIgXC89fEh9cWGp4VA3HYyH20ptgETLrOxrMh3gSZIBJDfgbh4L2FOyP
DIc+9mfZP6dnfTnwAUWCXno3qQaKfpX4nYB1Ngpb6SaVAkH3a3ExuwkOm0A5Dzjm5Hmd9vfZIHi4
Edu/SW7QJqgW1MZmaP0vdd0KT40uIx0Iwix2zBfaRQf6T6B3ep887vRkyHBtzdFTv9/g+cjo98f/
TrgSgvmdByWx+ZrXwCQdQmhYQLpfElFQCM9i8yJCyHKTDQMR1JWj9WZ2dTtm1ORFdCjU8nz08PdF
eYLpsFpUVjHKXucuuiBGgsWsC34xKB/+W8t3nZmqgqPgIIXYusVM82zZmEr9f8uXgF/PeKRS9OE4
l1dvLDTOFLqPEJiuSVAFiv+4U2KSDxswvRKZk4NgbqE9aQmghr5/DVvHVDMBPCIs4VGXsfwyJfLx
j0Zw3LJbkhVKwt9JJ45xJYxtDp1t3ZQeesDwzkx92VDsqio22sTcTUL1IwJEjJR1Oi0SiiLs8821
vFiPtgQIDjQxrZJJ7SrIh125KJcLdfEURIAopJxlD+b5xi/7UXSxF7YNN/phvgXlZxNqvgw/5BHx
RfC+yrCRXPsOGauxo7b6o5C2CyPMbCnQVS4KSLEzLiBmoxjviyl3EZ+d1vk6WJBp49TmSEUnQyTB
QuEaTvVCIL8zRaE0Pw38EPSYakNyEr73E4NWM2R8IH2vuHPDCrQG2GxRGjZqds6W6kjU4oNskpO1
YHFjmEap+Novhai+QsmNwevUJlwoSvBW3A0qZzCGl+2wmG6wBZFOQ+Yaj5ijnJGxSXnzPNhR+uAo
9mDxB3AGvttXJaIPLwVck6LiSYx2SBCMyFCSbRH4zA855UsXTu9SYIs+Z7eoksFYMzQgdxJkRmBl
wGwlwJ4bh5PV9JzpJnEnhEssUU4WdLgSiNvoe8jT6jOvXakKr1WM/YO3rtKrlHEFCE4owJ76hrMy
ndmETGjDY8wJlijs0fSmOx1Tty6+6zmKhSaebFyGwfY8dTfkZAjY4RXdDVHrwV2c1a6U2MErE7V9
KRoLcS+Yi8aNfyVuT9/kRMgGP8exJgZy668XxraH1IAkVnZjQyH9pYIHnUiknEx3EGPTbXFd24+H
aOswDBSaTxYB9Jj0fpw3RAMpE3IfE5wQYwMZZ9JdbadQId73z13aJgmgf183aVk8SYDnGmcEOU1B
6LMUGk43DWPEuvWiICt2oEqcY4oLna53OsZ1vBGHShnl8yjyVQW1KbSGmFkVdomB7VKuaERDFwxN
XPrXDUnXDHvviWe+UYp9pLwZ1lM1IANjDnjW/gWqVcLwQyAbmBd5YIzFy/6xopxK0DXw2BIFWDQq
joo1smg9MaLaGc/CIiI46jxIuCn/Ye/gW0v3AWXYApv2i3Y+Cd68IIw6Fv8GXSeUQQFbpn0eEMnj
lQogdRTOPEIQAjWqxd4lUE+XG5KiF+n3XP+2J7I3UJ7lS2OGrXUo+lICT6ZJ/JJTXPhxm8eL1N4W
+GSGAO5YVDYB7WrOsnOWSQ3WuRILjelIiwVuFlkVAXZjG4YDsC+b5Wtu5h9SNcYoGT/ZizYmgD6p
NVmOG09xUQuNrq5G1Wp5kAB/vC6jYv2sayuNWx1BZdA4wTXtDQiCJFTAyzSazzIcra8dI1myoIU3
c/tLr+l9Squv0aMKQ434HauTNTDiEHdZySIIS+y3I7e47JnYoj9qHZErPixeOpAQwYtAIlJBUS7i
YyQZNhgasXQfqlyNsgskQYFt7E8+lUKDZPqq/uJGyZR/KOV7auZENf7rzwSYooN8/2asRQhhznLW
b1i4HdN8naWLNNcz0HN62XJa2iUeLe+v3VakbNdXVh2x3fqqnOgfYbvEwJOLqCWLH+hOtf+XdcHL
+kUH4vqyb1lpPJwyxdiJnpGJp1X/HMjv38FtDmf2rnvzHmXhLy5qj9SLnIkQzPX0FEoAjPCJ/6Ki
GZa1Eo4EtTdmMrrP8iPhoDXqtOzkZUX691xdaYcQX0tDEiQ49JUxzPJN0rsAWd6e8TUN3BljARFB
EqTPdR7vxX/FqtgiQ99rXZaRnoa69DbYQ2+p/6Br8NASqRcREMxq2Ap2bhYVbrpSm+5AiEsv0YSN
2WGgmtEvvs4z3XdMXOXf8FZcOuP0UWWy/P4jRkOVCeZzyIGpkZaNq9Pjh+Wv0U38zxtPCjHcUZ59
NnguNZKchLffzK/7Zf2WEhGumGp5T6pjxyERDTfWNzQK0y56NRR89DH2NiqyQryqJLt5QPvkPCfm
BHtSLaRZymmUbd+fGr20QF1xThp3N73GuVs+SufmYTAFjgq9HnBIjmprXpgojtmOdbQ0WrdULU2v
eIUEPftxBXaurg9kbRPecfCwkTghI2WC+YTlkuTF4Wx2faaAlFmgFOisrAXEbORyJhzYERnV13lS
jGzLjWqjd5Fv5PatWmhUi1l5fxhRETQ1iEEE7MzFdt4UyANZP6/16eOf/mVJdzSRxow5wHtMz+tg
HEBet1Eu0PBym8fkVHz1IwJOiUbpmByw5HvNHAKpqq+srA9H5QyMu929qcTBEimwPRvc7PQ0FFT8
d226r+nCCGQS/6LkOeld9/Rbuf01OGVbj5hkjtw7o9p3NWdByg26+luUpR3HfrFo3vNjhp+tFSr3
DwGwkm/a9P3c6SrbBPDI8LEZJWvyDggzTts9GfO+y2yGeFZVB/v4PuVgMhDwZBoYE3KlV3SCOIS9
ertb9xVWGQdVJLwcor5I5jK2fzXq3xKlbXaL6jypc3AIWM6eKvUsZJX2ItEPqGG0rLeiIQIqcpFk
zTHEmVRKZAKlGdhASIMCLu9BFB+Gx7+JWDgM8q7oG7kaGioSufMAHsA6G7hnpY6/bysetx+VPme1
pjygORVYIF883E0TbCdic47EC3wmzy2/zgGBQR+PG/fveYTj1zaTNFKIoGq2s/g+eFfaZ4bBV99e
oA/akg52o+APq9kg/+BpXeUx25G6XZbvudgFr3qgU1/Uu7zMOV0BA3nts9uQOmcUDAzMq8wfaSq2
RvsJi6fyoMwAPyNKWcC0b/aP+TKwqgXH5atrjQy1mYBvEAexYUNO+wbLKqy3qRbTAz3wdP8OFTyc
OTgqvnhc2hOnq8tBWLp6HwgzArpcdp3O8O3tPUPTYDHfIBcMriqGFNt7Rwzg6MXewg6/6mKMDTgA
F2c9mSuC9B3rsiyxzbsLEmpE+AVBuF0voW05YDDLQSoHKGyzDxWyEgPf5ix0yrOIJRqge8PlRk9q
CSyf4sBVr/lU+piydNPELhU14WfhB3zDsSwmVzeRWM0/3JShGPbhTTr0RrA6KCVNwU22sIjOx6qQ
N/SLImgibxzt7EM7gQG2lkkd7+GP/i72RATK28CiyFyjgfL5S05XTu/+giW8XBSNZY+JXf1RiT3J
Y0bZIOsuKsYsbLVL64ak1K4kv48ZLGcAR54uG7Y9oPIqP0rWWQ4bK2bwEpT3suMOjHBxkzmPJOWh
yXF2QzZq1etOfqi8MORWe9kC3j4IJkJfuRP/DgJutK3l69yMDMb+9v9q0azMF4ebdk2q/SP8rKlB
g2gllUUwC7LgxyE1Byp0QJ7Iq3aSJB+31PuETQjS357BhlLiI5FEUWuk+fLUozMzFrfJH0rl/Ohu
yXGQaeEUy3O/s86T9cTGNUAnFTWwzp303kYfAvzzXxsDPHNGmEn0lLyQAbfK/FoCI/QKlSGwA7Wu
+YaYXlkyrxwmSjoHNBEJyZTunWHNJOE7yHv5yeQOBxnCd47FBhgwNXw+AHtD0R9eQATGj01HZvwp
EE4z/Jd88pVd2guFT6HImYd9iSwWabmk/MIqg6c1Vq3DzO7zlTIosxglfvqknh54ziJiiuqq8v0A
TRC22ebrnKQoeSTB/OiPvk4whp3TjURg7z4XOZv3AwVyyeaAw/OqsX3XzCTIuLuqqP6e4a7jWd35
q7yJmbe20YFo0DdfkH5st5+PAj3xh7BwSxdEBx4mDWfKLGZDR1ele8OQg0+eldR7RLP2lOhjbLeV
aK77FbVEYh3VJFqI6+ulJceZRA8ZM8U7MZQTetRGCUWhoXJ+PVj1myOPEIV/aU/CvFSKI9/EmqXa
Uc3UZGVefdqbGcUG9xkpdvSizplAldM60vofGRISAOWB7/4NYT+E1FTukehF/0UvhQ9tW60cCPXw
D/oww76KQXwUda22WD8DXBJxSyrYKh0eFEZ0E/dfxs/6Jf5mZzEWj6nfxTu4rerANN3d44fXJ1h3
RxRyw7b1XKQsFBZlCh+loxSSqIXG6OmkY0ZD4ZaQr5/M0NHMGvhimAtcf1KpBjH0ZIQIhHJjFZC6
JzRkwtSj9xNTTA97BJk6p3iQlwmNpXjGN5/FNQ4XnSdmiebGXtDMPOeatdXEmv9YLmNlrLwXeDEU
1pVamHYxBgPupSPpPwb4N/6BB26JwaUxlN68WjuCuh152VmZEV+ryWgwOTchFYcUHKBVcqDFBgE6
PPWaIG7dbJTO44i+gaBOpEFkk8r/AL7DXTeKGo2XrmliBLgzQ+Gmu4X3GOryLaYl+IiVzlZ3ZD3k
sHdtE6VRb0D+p/deokWo/REK/BDWUaH7UkTrfjSj3McZ+eBkBxqqBHPrDtAMMec3++NIEQW/NK7Z
JhJu1+b9DdCyYvD12WkBypBzm1vDTsujOsVrQ2x4/GB5Am0tLhZxQxlDlKH6PXCZBJklzujaJwP/
GPeqOGn20I6Try8SMQFfEIHk4OxGqiMS7VQblBFjKfco8FcxmegpTpRbxma9o6bIjcTy6NkJEYtk
RP3CNFDn1XmG4JsmESdld92aWCWFSZVUDVmtQkvUH0xnsrUvRrVuVTHa34Tf/2IoSjYCZsaaUntQ
MEqbFOgkFw1WkkxjtDvJINVyZkCJGFKH2moD36GrOvERYokn1SBLWYDbRq2/MS+u5GWrBghPPVaX
wW+Ocf7xSgv/Akj+qc9h8uD0XpF7v0alwofg/qtqYOa5BDAseb1+zeiymULIlYjr0jW/o0+f3f2F
5kj9uZzbK5XAoSwwgeH2yNH28E6tTHMU43H4VjB9h7Lk5/N8oMpoCNYfrBs5V5aM/hjIf5e2ekKa
w9SJSnoLvedtg58z2/VswQYgnZw5L7/UhERR99OlYAqdfJaJZXBsTbfwg62SXm+JZ6xN1RhWKlfu
MD655el+sPFjkj6XcIFM6FIsZ2B121ZHSEuyfMAn8+LnQW0P3PyTklOxZBs3FSu0wnze5wy0um+8
xBRDNwUFOGOWTCqR87jemgqDsUr4t2dQesI0Uea+NPjJx3eIOYHIxtyApP9oi0wVXQugTl8kyvuD
vTOoC9DX66nxtP10ACu1nNCF9qM2LefrgjTU91L4qyWpaK7eN/hJl30dCFx0pq+rA/tyWx7sW1Dx
HOG4g0lpBBAEgd30X3925hooXR994l08h8oDDo/R1cnKNdeQEgudpbkMZYZO7fjP0ZzXmvoR8sPj
YurTNzC/7WS4rI57TzFNkG0HeFu3Kct2pys81D88JhYFs+vm3o19Z9y9/v3qdgz5ShwKQzmkx0a/
1pqv5O1zsQNOcceReXupGzja16TIaDTb8iX5dNittXkIdKrTqQZQdYJ3u0revR8uiqlaiA/LE9Ly
3HPCGiILvm8ICpdN22rJaDw5gbHHNHuHyRmUA0mVmVUfBsYA4ZuHfsD2B+J/JpTcZfHoCgTQkWzw
xnrK9HSmTeCvkrv7LA6xSkvnkvhFE2lrPDKMjxBCU972In/rbpCDyJziTbjjmNf98ekmxOG/YHjP
KA3M6VvBat6s9cdyi2yZXbJmeY0LgFkbp+30Nq7ZY9ke7racA4LND/XqTYjia9BltzN+T+aZdsM9
nM5y5vwtEbYsBSGxQHqYejfaSyNuiRBzKFtIIezqOi7gubsZvNfICAYY19PYMZs89/OdBLKIr0pd
mcvgIldLozJUQpLhLecZ1Akx6JigRZdEXJAQj9qEnIK9h6v5Jt3JLyX27nvXqkbd3xbmofEEQtfy
ir3DoZColQkmnHvHeWFvw82oqxwtXMWOQ7UlUL8iAbtKYZd3fVkJa2IbigfpdJUshT/BnP7eulH5
cBdYKivN6ytUAtOqrPtwnCE+rZa0PbnV+9XD+/0T6fNbePeATp+Am5G+turLpLXT6OrKIIGWEnmB
qLj6hHj9yjcgoU9nOH7+vHG3NcOB6OOlB7wrXbc3S4rTyJeNSZAPXj19CNXjAopx4sGKuG6NEovG
Udh08cL9kTxF7aFJkrz+O7w0IqbBbz+xfsQpWRSnPvwiy2/HFuERfJyoPs1PB/xELv34bu5z+K7v
IOIs1rqFqGkq0hKkQbvAKSWplUwfrl+7wws9rGFERowXDULHk9XEig/jBZxTcu6sxF2jh3d/YG85
DrZKb1QyYqMc+DSUMwBaKBLPc3wEaPVVRtfacgodItwMOxbXADcEGSFBo/ZmQOBpTVYiv/8jbRlD
t62EWi5hLMdqyyL/uxz2IbTtxtgK2R4kwD+jueZ+fs0dyZDouH/3BEIM85db0uAOLi3ridTlKrHN
ikhSQQzoHPLyUwGPuX59YkTIv8YKmBE1QFyiV+Tg89lFExluO2nwxeXDUJ1uS3Z57RD1VeKoXWOT
5C5xwpKyM9lDJbJ0A7OvV9wGoYT22uw0cGXnIXY1vjnduOZyJFaN3LJMkO1WB9GbTFIEioaHqCIm
jIreDvr7rD7WgoMhojwBp0Z13Io6kTdYRJmedeAN0lB+yvV27AHGT4zHfqmtEc9+LscI+zmy/13v
7mbu3/i+0HTrICdukULbfn23RHrg/Jp9or9e7KtDC/Mcvlthxmu68qPEXbscZhinUw9RDlbYK3oM
Zt0RdDI2Nv4BLAT/nu8jJg9OdCR40kXl0knZ+nBVB3bPNp2+2mTf4iBa0KZ75wmXmaQHwy+mZZWy
PBOTOnKACVWQXMwjD4tEMm01QNaQsqtjMa/t+xk5m31VAVzOcb7aOs+rDWyJEWZRHkF7C5jaObls
Cp5R4ZmOUZY/Az5VX47ObDNQ07cKHGtH9tlsJ4Fa0vbTHwuVAhBdAET9AnRsVCkSdARYwl7aCp1V
m2nNwH8VyGR1Y9/Wp0+iUUzIzDbe7YwdVmtm+t4ZpEGeNg2dwc3gPxZxdirfYK4qydIg65ZqL0BM
uxGQ9zonEtJ3pvss9tZW9huv7JlkqwUsNjnhNZ71JRHGqIf2iBPspdRQQ10e8tfih5OhasF05nKo
wHv760sHeI8GJHaxN1F8/WcLw/kBDcz6vzYglEbRW2374x/E/RdKFQQTMdQSt3jstjxQlK39z67z
W1lq9QIor5NB83TG0IXzR+e1CJnG+Bj9SPsa0UCa8UqgWG21gMB3+UlIbXCmqDMeVBRGjIlykOU/
JOTVjfdTIO+aaKUoDW67CGKb8HcT9x5/p0geH+RgeiBWMUnD4i4DVDQtpUkWjY8XsUK7vthtIuB5
6xhExKKq1X1Bv6sKPO0dV581VkX1Iusr5mAsvuN55GE583nEqqSXj3nQQnaQ0iBuZRc1mZF75rsZ
giarPJMZ7uLLrGc+noIfz9WymycblNe/AbKiqAJSIjU60fViiIgNOH8WeMYl8BJsPedM7gjc87Vt
J9sAUxgQynvr3zt3VN5BLH0XwxQBYoIsmAxIBDPg5q/eXaiegEtawcIQIXfRUPXHqVt9TkVNCFMY
TZRnasRfb0eOj7SHF1DZRCDFGWs/XuO1zkRH4MKlI8u5Xub25YOGC0SKJEBycudUP0G3bEjYwpZi
gYgW2xIlmWGOn/oc8SyzCQyFzqs7jgKq0HP28qgmMNHkAKotbe8Xg0GrNs63e1Cas+9FjOVJFCeh
IDoxZ5Kpmqu9s+6roC3gku/+nBredfWlWaClDnw6qUX9wp3OfwOMZPLFzwRI9Nc5ia/4Aua8bEgs
DzM8RP8pf4gQndSEXF7pGhAM+c0rYLnrdtQk7nkWXFBqNFnze1AajzjVBUCtVI662CPuyCEOIvhK
kGWCbYG0+NQ3T9NaBFRZA637g0QRo5s0CCSqeY2Ln0cMrn6cl61ZWLTIBkljyMCd5KE0dpgZIc97
ZpdL2BCGuvkYsPnnL3qlts6Sa4q2wb7MmfLzP2YOv+QG29zJTY1Zd4dlVm6j7BmrDCWmqoiEJi3R
3W+B1ACtj1muAC2yeqORj8h739jGnNCwhXIs5HvUrtDKMlkmtdsJ2gcXIveFBs3Y6Zg/F1+j3+jM
bhGci+MWljBjmecuxgUqxdkI2uABXqnC49VPrqvpMB+oIQxyt9wuvgApw54Mi9BOk4ilcFIhGjZc
LG9Gc3wSqJX8P1xcOEUfsUMkgah9P7NbabN+aBLmUhpjrI2wB+VaqQS+yiw7Ejn3kONcR95kkM6F
2Cx0yjAY86uf2xglqULVtKXz6xylSOHGlU3x3XXF4SEeEuvbApt41RBx5ET6W04zgsadDGRTMm79
TnXB9qFcJtNMrqZaGdUoiessbBHnPLemw3o1oL+5xqxKeFuxC1Sa+vrVINM9Pd3JDc0UqsQv+foP
G7nkPxGEKb5UkBXMFrlrUxBDxhyBxae++PHkFi2N5X9K8nLGaXQGiZLoWUIUh74LXiEnxSfYvbLm
4VRb6nhfBND8D+dyn5Kdxhx3oNuXa+QAHbsPEOvbsaIZ3cUkErHxH+QJzp2Km34hChz/Iv8twriD
wq+glb9qBfemg2dSenntmgzLXkq+lmknlQaS/N+omvXY8Cu1Q39OJvRInAFXjkekKd1Zcx9zf1E0
UC+phT3ldRLH6PLW1v7g2fNSV38LMmIxvM5mg2aXhwyFwvXnzfHVRmbpddgVKurBK2LN8LLaLKka
Q4iiIoMjZRPzo+btTC4ROCfcu8KE3l5BYXDsFzGotTgrLUU+IzysHxrV1pzlN9HxSn2JrEFwk3cO
aCNQY+Kvy3bgksXFRvfJlcxFdRj3vdHvPD0YSmi5zhoHRqikD00WxMJC0tR9XR+Q0SI80PaFT6XB
jfbbk3+kabJ9bBS2/Z6nBLRkSlRESZJO7juoPJCM2U6m07jWT0uxVXYx1QeEVBdJLBx1HfMOWqS9
TT/vfy9SzMGTqxCy5MrURh0jCgaSDuVQG4G3js5D7yRpV3CTN3bfPu6CRbuYvxEpBGHwjIPmoCzk
DVivK7T4ZGJnOZMKfLwO64cYNCn6IK+VeBIGNBa3auN6Vq1+5PqQKLF8TAwVXwwhU0hQmw3Q4S7B
6OTMwm0MHKdEf7Y0ON5uZa8CQTbiwnXOPvUqhJVmvkbIxjkE5vT3KbayvwNpY9rBOMeorq7RJ7e9
VXue822iuRWFaZibDuEUOS7Rt+ZnzU2it8ZRs5zZfipAsiToPmEVjhIxHrVfsZbPLz+bToVur4LP
RNCQawiI/SI1teGyGcyEF49TfDBpAbkaeQcUF4mjx3KLKCnp2HLMMeZvtxDTmp281B2z87CYip0c
LDcRfZxU+oRszde1QB+0v3pSe0hXDtOEkxJ98nTm4sO8Hf01hypW/HNe6mPWGSk5hsGXwRbZnNEc
DxPT7rlWNlO8Fvo28aU+/5aDXufGhL9s+7HlBhcmzPuX7MIQU1izMRJXVlEymMAy93DfenLcTN5/
FYn1vaFX4ePMS0RnA1SEAZsUKkoIkO84IkYL6rjHycE7xSRl2PaiBqvqNqsj6ofv8GEKTMdQM/rd
I4ZP6jED4Qdnq98nqrVZY0DUYO9JxALHjcq/I6gte36mxx//y4j1Jn5rUi8eqgppNLr2e0GmvsUC
F51w5PZEGY2moTNwFkieKWXEZyWLh/Do7a1CoCJq+C7HwcueNS12JezrtgBMlJ6vQVsLa/GogaLO
ZlbwyR0zAnPwW3t/4/rfFF7QKuGwTAiohErIWGvhBuaV7pH4RQ8mcdOOXuZEWUGpRLxw5YRiJleU
S1lqqhLZtJvSnNJ+BLMkKv0r9HkpEPQ7HbVQ2wQXVJ6yUXHXW/G3fGKnL0WJvyGLkawxD10T+e1K
Shjgtv05SGFS1B7to2tmNsB58DDzhtwMmcYu9C+7DBfO6VmTCZdsse+vJLZCfFMCgGmJ/38CqYkd
iflQKTSHdg1WsA4XGDVhQySPkMTc/wvw3y6WuGBdyMcEp6sTVGh38mRpIpQm5EWvuUMMXn5zXxOr
9YFG3lvAV+Lf3qU2lWnuvNwuNw9dEqea+1+wqlypWfBW1DaSqLf14VzK0pgiqJ1+tOX4krPINfFT
NPwh1xJfcrzIFmByN22dBh0ZAXfZvLVtWMjvGrvVyL5W74C1iNfwUCSGA3GJD1PuB+C6bYkJj8+g
Z1rYcs2UinlzVZpp+RHNFWAOT9/X4CE/SQuTLztiDoUneh67SIfjYBc+qBwkd1wzBnUmM3MdFohj
9l9uwnuZxy1ElxeTNquqZqmbTbWuiz2wusBr6dqbrC9+b9jgK7YjIvda7dTAonD3hm2TrCeuTYXI
uABW7zjXXQYKoYiSG8utUpoFCxHHE2p59lNC7A1/271h3gFWxBaCYZQS9IXkrYBLEWb6rjJQh/UR
PqIdy/KzD8SOYqtW3Hh7HSryDKlreUbzgarjOK41yaC312WWWl6U204HSZcPLokk2R+Cqf6GNsZU
VyFEs7APg12OL887EP5T1P8pZbNeb3X1Dn8f9kvm/gtdt/bcPpCPR6Y/4bX186QnBiAWnaDyw+j+
3F1uBRneJiwyXPYL9wwuv4kkXC/MbC3s7y25UHa0Jkpw9t/qzGd5TV6kopu99bEifCG0eFUtWybY
LOmUdqjYIQBIblD86wfaLmPghXhjH3FQjFnWqeDagZVt0kmKevGUotXvHNSiQtfjteoCIbDedhQH
uBsakOHdRQwNs6Px/0F7otqbtutdstpgXNQ5/khfFAcsHMWpFuwMh8FdjEWwELb0GwY/fey6nynN
ByUBdLS63wXMjb/fUpkCwl9q8Gy279UFp/qlloERFuNlUXVP++dfQ0adguOoboQnGo50zzynmc7G
QvXBRh2GKcJrlvY4/u6RjdmTLYlqxyIGhKvLoSlxeOv7cfQ2RjHLViQ86uzwIjBzkCQ1sKbjoJQb
Ug4l2A5ijpRYal+/osWO1olt/VWP8SeU+wSO050YMdomcS4iBa44DFIfphWzuUyCpkPtzknw7HZM
qi2Si7iDB3GIYHKk7onvuYpZJDbeeCKOkvvxPwI7sYqPK9UxfBHYMkQCy2EjXKFzDXw8mn1iwHAV
MHP25N85ECMVWq6Zd+ikMyYqB9R2AnwL6Ry8rl/kgUYAMe9lQy0RCn+c3debz2zDpKG/ldt15w4r
P4hpvu06KZNHWItQ/y+6Z5nnFoKk1pf+5Gz4KJrPmCIBwP0uAXbekzIOXUw+g8LBdaDunHO3vG4j
8tbI5X5yp/3LKG3Gi63X7+2yvMWnTKtnq7RtqjVv0Io1eYftbPUMLoVDhpPgkJvCGGulwkW3VCaS
wCY4Bg9lQ6eRIv1oLy6cOjup33bw90lMMCns+uTZYZXyFHQKlmv8Zy6ANccYS45xAw7BPiLnqeq7
jcKIAgp7CSgyO+g/Te38opnFVHqIvS3aZ4erlrAYIPhVbM5xSWyoJ4qNN0DpB25mCGkFOkxZYf4D
sWgqODLyMlQPHAaGi98W52Qryh4lav1EgsFpedIBuB8daOYKZa2VfvMGxqzrBo3TE9vO0SQTug8g
uGGq05Kiw4NQ4VceK04PD9avNRzoPQxapvxXzjPtYjXjUIgvZew0OOU0yJIIllNvWbOP4NoKUJWY
kzBhYFpJ/nMg6GCtzZK+4bH/Cwi2/Yl5h0VB8GV85KOvIWorBlDUgaEhOllo7W8E/9Z5ORb1gDAI
6BTqOGnUxVHV/C9hddDmexEseFigLGgsA8AZ7PF6mJzI5nZcncUvZpqFAe4TBGHH2Kk3wkV7jEA6
sAuP6vYTWWrmdAgZhvG4TxwYu3LdeuJXCAkxck9oQFtN3ACGF94u+C9ETRjBqVOFTP17op6U7zdb
mOKtM2Y194NNUpPD1tT/t/p7wnodZ87ygmTl7viz3bz42U35a/BXCBz1NCb7BZqZSIg6MFJO5Mgr
kCQQ7H2vreTvkiFsxMkhCAQPjpcTeQQavlnqLg4IYrPdWdiBdj5kNePC9NDAy8fLVOlS+L0qxlds
a1vqhuUuS/PYhQgYPvW2vdUWen3vhMNbeCL0z01wdSBCh2Pkp/EQQUaZreV/Q2LOMxgAmBE8fOIK
N9tvWM26wL9KIkbQ5KJ2c4XPfS9F0fUcquoBWxiM6TMFgiIY4lS8QNrb7LVknqjQmFFCztdtu3b8
FTLxgBgv9XzGQcr/MwV9JRbGeW5PcdS25YOdUz1Fub6l5n1EVAqHcVjRkDkUzv4FTykXpzTdx1So
43gc4QNVq4XBNZeLX46+tS7pgX5AhJzY605Jo3U1o3RZ4WbnIsP9937nPbXSFhITRZB1D6Gey0Jj
q7zVJsbEzwuOWRa+ufk70vpNQ5II1xAEhWeJseCfDOmxjp50EtUarHnmJvw2nwZmDqZCH0LtosNM
zay3PbG1ThFNOueAEVa/AUvZWkrAkN2oHA+enl8qv6bnostXUvmFr9dE7oAT8MYS+p5HVFaNVS/U
450U7NI5Xg4jqj4MUPUjjsiFolSX6MxafYbef42sYe/1e6eNLTHTRZ+0Gfc72aWQOnrvk8+yd2Da
2xr0QC3LNUljoyT8Cv9XbFC2DU+obdhSW9WEbaZRCcCyX8jGYvSRn24DxmiH1dCdIscAfz0+1ltD
tBuoNpycKkCKg92iKrUwYfuBSdefV4Y58mK4DqWMhcJn712MKLnFz6g1q5DuN8m/c02QZy7AVasQ
yvIWre47wXURXuIgy25JzHhv9i3gNtl36oIXnIlEzQFGEJEhSiQ+stjrBbtEbcp+IOwpMJ1tqAQb
Em515WJKhQ3sG+tucwbdfQGAp/Kps9FKoNb1rtnisQ8rnHJU05KPxavgD93QZnyNy+PqpPmSljgM
fc28XW2cfsku+TA4mQlW9YTGjQPpHAZg+R9ul2QuWPLk1RIn9vLH31s4zNGcx992qaaz7vpQB2tG
8dfKAPfOlQA98B51QLTr4AEg9KsN6+xVmGTLnr9p2c/G/9EdNY8AIToTsPnkcXYxPpBYwN3nel5d
paEZ0i8vu5/zzPe4WJplLyDgCcM8C4QC9lC3OY1K6PE0VafdKChzVnxjZwDSYxdQSnJel/+ZDOF3
LYC6r7tMOQVZ4im9bMsxBdh5R3jFvyCOHcli8RfIK65p34cpfRWyjZ69Orla94QYHBlctyNJ0xM1
fiLcRVGODAlNG/k6pnvY+9wGMQ9xvZnCymceg1DPkikajNvV8/bBDzuhHO8L46RtmrwQmOE79P2P
KOg1J8X2oDRYdkEqe1qViTqBO/JAKfwiAkxbq6aBNx196ITjlys+jGc/VnJPKLuvOQjxgT15OkxX
Fk9pXmO4oI8vHgFmxUP+gItDoCRrqDj4i84IaXmEK0c30onwO9vE5xGCw7vAQrHTCixu97kU1bQW
N5k+/Q1BdkpEf6BP/d8DICOrbTy9HeBayoRifGv0vZYcySW8whnqp72zIMnAe9Qcuy/hqlePDPvA
qPNALSy+Oc+0xA7YMn5Xteu7vDb9UbB/BhqTillNIf7MQB5Bu4Sgf2GBSG29b6G1yqjE8wvyzXnC
cunqTAbWHdgIQiJxoS23QdsnG5OHii0WZelNSZbiV+6lAu/dxhji+vP/qXOr4/OM8xwuc87Y3PTI
vvEmdVYzBbS59b27QCOcIpSb4LNxNzqcn9pUotTQH61cX8/yTcvR+o48Q2xRFC5K3+WNpNKrf2e+
3K4XaA9EeOg3PdUr6VH1EDLM9JJgeDQgreoSJQiM9Fnj5CcpC2paqbL/r/h+xMylx43Aqt+W46Xg
0wixa6X1d4vNCrtYjHu8zSGJJp23rT8T5ofM8sBROLRDxFFyqWFfS4IueIbvfd0AeBmR0hC0mC52
yO5wM93F7A08v02qp9eFMGlKT2roEwaNhy3Gh5+8MPulbYIeb/6YmaN8JIln6XIL0hABU9H7ldvA
g5ADIpC1XzwSv65TwoxEbsOyHYh0p0F2OwB0gY+hz2OikkncIEDBrIZIO0qFpdViDgItQ2w+9F0r
/CW0tPt8jyJCrZP/o9T/k4RE9EALJIucEwdVaWrc3EfA3ijaikosy9cYYuqnTC1gcaJOjFUYCqQi
Gt+stE2MA9WeBRmELJEwoQOipCYXqfDrXM3eebFt+RJDf6sjlg4SGkMDHZtz2IRQnP4dSiZoQPKW
mvDLxjoQKfpbuOGZHGXoK9wz9j/DY4XyFEgudnvrimOhz+76kpazhY0MT4UauzNDsaX4A6bhCMS3
pDKHc9P0gWZ2L4jpTFLXPGaFSxgRQqywRcFKQ9mq6aeR7Hw4flnL2ROvEsU6XQ88Y1ZQTuks0lKz
DGLUO2vf/fcu594+ADz4M9y/Gkb89LezoH68Jf9YR6r8Zh5AjpdvBwgJrR1INWodwdCOz09o8DOB
JdGtrBLLvEXwZy1dEn0kFtVzBXq5twQ7vHrkeXhBr58jcb2ppdLLc8pyNSGdsFOOFF9pUVASP14J
fB1MYBnXnOQuc2RGvkhEx78TtSQqIpgilG3JV/bVBTCRMrL+33g52wgvobNtNr/KE6EFtcw4exoS
HUoKdZBaGVpRs6dbDacK8tE08H5ADa0S3XPlK9ojHdGEEaE4c5HImCIpXDwH9HE1z89fZUIETAvp
whOAdXEGarlxyGanpH+eJxp+5O+YedOlq06FH3FTJMoCqPgqi2ZS9lK5B3xiDp7fQiZ+vdFlEKzD
i8wwXJYWgmKqrGSiDf3eXQuQmmSvi8to2OeftdMNc1SdRIjlIrNKLxhncs/tdNSeNu5Buuwh8CVi
TSaF7VW/snI/HkPL9btNbpiZtMkdUINA1SIyH7jrteq/CUvWzD1YjzcfUcJSjSTyd+kMEW0zbhyd
rjkA7r3moWo0KDk9QKcxWq0GIVbveX4CKTHrzmAnRbPWg1p5vUnWOHr4h1uSPtVKqutnujTeu4Z4
Ihs1unbehVME2NWJJG1ZY0gDH67lGrR8Ee1VZXtibKL1BWIopxWa0ccwcZur4r2iyagvkv/bcBuS
LAW32PSB6rb/cMSrw/Z4A6pnC9pnH9Vq+Gyln2p3WhVNhslIiZ71CCcMjMNyfgUwfYdYf+5W96Tg
JV991fOk+rorRf5hIzs5SkyH7j45KkSwDii7/N2flDu6MVEopTOy2yVQMdSODhruk1aQeqf/9pEq
dj8Ujk93+9Qz6Z5ZpZ17wsZz7WgSmn06XouXivHOXyIDW/Q2lMUY19EhT8U6RH0VBq/DAJMt872L
ZES7oheCO/Fm9pAny7RfRCZNQcGEFpMLQOusOgqKRMoOuKWgS0JXAH0WYh7DdMtllQW12ZH2HJjn
H+ahAkshos48bX121dfPzWdpUS1AUX6QitbbD4WrH1CL5FQlTM9qp3OkScyAXZARnZJCUZxL4S7l
bfEPV6IOf0sa9fS+FBHEz++qQFSgLnuhwafPgSVZv3k/drmFnI2AVgBWvYpKdxErel2xxXwIPVQD
jQuFvSu/ApXHXQC03MSMiVi4EbtnPDmuGJ/8Qv4P/UbDJ2tEgK+VpTz7p6xuuJs5mY7jsjiOo3RN
CgrsQhQ7kapcDsI+Cqzdvg5VA57aw6oQCxwBDur4LU7ofBu7R2qUGu9+3F6tE8LM0jscrSYsqBre
Z/I8iU5cWbxBIb27nQvSvvBwXUk3o3P/2FaNYS9YaFyKs2wRs0ywBJ0iDJzvRfBIQohC/76A64Wu
+nDd5YhPUBkep1MZJosHl/zt7BRL3GymQmvmuEPC5XyqGdaiSffkEVgC7Yxz0S7wgkGp4FwrYFB2
O5cbSBSJXBDImqEjxntJdLYt3If2kGOsfhaOnwM9F758gZoXxEalEtvxmTmlbu3VFMTxjbazv9Jp
MLh0v4rI8vJh4rQaWeuEsQT9gc0NULbVYGLUeWLh6Um1bDo/gkNgE/CxLHIjhmTFebF3LYb5k4aT
uwzdtjx/2jWRxlaE/DKFwOg3yzwRkKoRd2qgwfVRwgAOybgpWumjA0Pd58wJYfd066cfrUgXT2po
dIWyP9kq7qGXIiHQ4Q2Dhfk52p69MSHr57ce6X63G7B3qwJZ4zGL14jNsX7ajRlXWTALeyPWzkP1
WpQn+c0SO+eNsDoVOG5JryAcK4pVIhfPtXOW4NxS9ezj+Dl353E+gHNXjsDsHmYJcXKVtoP0vZpx
S9IuwyA29i4EvfR2xRY/4MeEq8dpKxAawJNjFWvH2cE39EkAaNF/Ppu3pjojFGtSMdOIK4G5W/2q
gWxOtsmfJCWSW59n/q51N6IMyMOgGzYLqXfvFxZYC3LGQuJA67Pi/wNfWSldRglDqihlTedpXQpi
fKEOkXhfZ4emnkoCdGJkNd3idZ3I9GBpozx/UN6I2L1N3OTVGyZwDbjXI3WSFQlyG56j02vB1fHD
3lzojqUjynvhVzQmqjWmZHvhzTObVjaba0bStBZX4MWnSf87IHSx0gmwU7cehOMw3kyXt7ll3Fri
jSO1besgiLwIT58J53o3W/0/L/FiRv2QOLp+t9bm3nbxgJ9feosG0kdT3M0yyjBnqS4LgO+uZuQs
u9+AOYcn5slpv6t1PCIxgd9ciBIlBr5JkChbuU2xsVcEU2IcTMveUKBo/1FhWmlNsBmknaIN7OpP
G+uqOr6xT/B8uxl7jlvJ4sT4MK40eR8IbIDWVzkfd0gCsyDAAba4mYVTcdxS1UoslcOgyeA4uS8a
OxzVzGxdHqlw0DbvK7xMrhft14xOpozALhh5ihdVihZ3fbNvXYZkHGLXmdoExiFzo8AWZUdFktgk
5lvMzjQPpGxBobENwk9saAjq2/wXKSG14+SWtUNctd5OMdphCY3Ty7Mc9no1sV3rF6UhKWGiBAAW
S61wSnbo1IrVyPfPQFkgPDZm4qDrvqAtTkPNDlmepHGdm+gFgw4orHZhYeS5sfvTGqDdkoSrxoDH
2RsxuRi6AsV5h9Ut3ATzhveKZCUBfUUcSr2fRIvlJyPgo9cLRKjunLbXRzuR9aLVAoRRkVcyZM0r
KmIqPD1wXcVG8KFXq5f1nR5RpD6AJSbOLRo/aYoBBV0V9hVIp/JSiebvcRXYhnnW/VYy6PdqfuFr
09JW7lUWmlWHSRfLwzed/gTHFDgEhwaURUkJbTje35fgcKqO8O/3ZAyadXXIzCp+pLcpQcFdAXji
zKVjnEVBFuithZ5KlHV/FiYm42Be56i+YDetQANkvLUHWB/MqXdbsDEJjHR+dPw4/feZrreEf2H9
ZhvPQFlzT6A/6PsliohOwVBVCKorcuarOhVpnym0mw2Y8Kf8sXIu+Bhq6EyAtirmx6KnafE9/PTh
dV5YZGvawGrPWvYTV/IykYozSffyLp+AbT7DJkszXrwTu9Zp/z0UihCxw+mLvcuv3GWsaqeKevV7
/wX8ZHHrz/y1RLjNqJRz/8/TfqrA6yHf6vcMfAr4ztIl/33uSGERA5Nabzf1AHQoIbSHwMeVVkZ6
e8JftEedNDIKXMSebf+C1lLOrhPP+kunZ43OSQBam0mVvr/GIb9ROgnM1MKohNOHrvB0QXIITpKj
FDqVSLPLlB6aERjqQ0EaaTC56sYHUiC0LJSgvwAPjYhsstpzvREF8SZp1Wx6XEu+n3LVHYvsLchZ
Agi6rSjGbyFB01XKzkSWR6+BjSQhdI6eNF4z4CPGRl5Dp9mNU/GlgKzfceiyTEWJ8mDt4iYdc/9e
6HFKZqY5mlj8KdQrQaEyeb4FEl2Hwul6YxKMgDxzL0zEN3a5NM37i3WlDYUjAUbwUiFPfhWPqIKa
GI3VF21GNKcx9l1n/zkGhFyF6x/5gyvquH2DeisHYGXGe4FkkVJWjkAU/71w3pbeST+xvrmrdGjc
N2YLWyms6xTnlN64tMvY0zcHnaGd+l7Wu+HRLQtuWro2pgKUU/fUAcU9TiZ+Emr8nHQuGNaPirM9
AqSdDeXeJyfE+L7004CacbmWibHX/aGbjdVAp3OA1wTkOYPb6YkoX7mSse1afwpktOELaWHmWX5z
R6CFnemPz06sWHvsFucd6W7TpHWYg5GXnEq6bcS2MIuqFfUnWOnnEhlig7VO01gWiruOe4Ja34wM
yJEiuDuz8vgObVcQbH0J1zN2R0YBW07P0mCpaqe9aQFAxELRKf9L7QkzEpjm24gzFiXk/ePxZyup
CMrGJKuOGnPX9LDRkRb01edwdkbczHxxp5Zj+Axp9nR/u5SMj92L1QokvBCCrThPQEgZWBM8rxcS
Q29ecdQBYzuwUcHTRDwbuvDNu/M6+p9bNmcaTgqtcnTBmlqxzSfYsPLtPUiUV0O8jgIggV06yFjZ
otY3hFX+eLDZ0JhhraNzzODvGAUjc34vuw8d1/xtt29NXWBESeWi++v7KOd/hbEpuaIERbfwG6M6
LFnESIZbbZunIy3xHp4okvHNHOq+OVS79wuAGenaVGkwqp+qUxbBLfFB3Ng+dKahO3rPV6Kz5o7l
jamGMFLGiPgD5VLdGBUv81+5Row0huTbqgsi0gagYZ9NwPCPbz5worQ/cQa8EwBN6CG7kHDYvqZQ
esHGczxMXEYEHQbhExbVhS4eBVQB4bGcwYIf0PEokJLXI1+BD+dkR1TR8PN14rqazPEP3bdHvnoB
B7ReSV6N2A3xC0v3FwZGmxRI+ub36Gy8q7OJF8U7bR2DMOHEZ5WLQV22vXbcDtzdZejrUs+XXcW0
1oTOzNWo/gdNXiQfmEYQYMmZWVhGPv13tpiS3TyqV5HiNTRzaC/1mZ/x4yDoV7I+h2cOaEt0I30l
RfmU+KavdndpVgOJ50Ufg0YsVC0r1DSHbvw0Y2LPRb4d9SCQ3YO+5vyjyvAbpdNe324D+5oxk+ub
yGgfZQsFAZA/Qnhfcz7/nbk9T2s61znbhIVuRzTjlyNJRS8rUrrKtRtHPD9oTsws37YOXRqvaaMo
i03QVB6rx7RSwhSwmbJ6DIwJ/u3tQ4xP/lHDk6qrzeAekTpVMuZrSt2oeoAd9DrlGG4Uh11PHRMK
WMNp5I1T91IMGhr64MdcA2CLzXy4894UbV5GHK9aV7AbodEYkxeXbk5U2lJIWmI83FjBAd85A3Fj
b0k2s5Vl7akqf/AjX3cGOnCsNYM4W4S3IXmLRPxN3f63YSBo+1WWJya7iWvksw3mZVmgj5A7TV0z
VVtsw/dgNv1EgzDtT54DjmJG4NYmFre3xedJucHGb6s3r2aQ6y/byx41TNYd0Li2LzaKZ3eTKtVa
QrWgl0Hac94LcG/N1u6PBjeM3iuYZPvskPUlToG/LHZA+tKoUNXetg+lW8slREIWXli2fEj/gpPO
QCbPq6FExY0Q5egxCtAGf/NEcnUkgvz5F1s+U6bnZEH5QsKm+Xis6C2/uu/Em1rKqnn+OrP+aecI
x9uCQ4wM/uzogR1iz1kPl/LJtF3vj+DHAlLkGKqjRKZIwBzQ3wD5ee8B1/g/17wbm5oaeU1iB7kQ
joB6+7Av5MITE7WB68JebIVqOjH9rbsflkAjftdQSGHwAxGNthgUW3aYiTpDUdOOqr/H13crV6db
5293Oy8VjO+EuBAQR2g19y6/kztHlF8R4FYGUPqaD8gejM+uCOu/Brn6cev/W7cd1B02pURfOeR4
7cTgwAcJUgEUHT4V00mZNtxbs91S4FOHGxLKfeno5vAgtM0RX+5FB2yELKO2qvxayC54Bv4hR+EG
L1WbwI7HYtxQ6uAwqgI2wAC4At1Ytq4o7ifU5cMU8pnVjmwv3x+enQZEdel3WlizlXxlcQ5klACr
M98ZdeRzNTy5NKZwW6qDpfLz7R4T6Ge+bYAvRAI4s75JUZJ2sbKk7yU3rCLV7LSMbrkC7GuBv3Ah
Sb1gE7XMFT43rfFNiUIIB/slEKbMPuPX7uZipztJKQQAgqKZRE8dZSiPwlwcu3nmu7lmDoyEaIKB
W6fikjgjQ6aPCE1Oua0H0rMD7mi6f3r/bP+l1TOvjhm1NrdgojBYzbATBbm0GW9uDxyE90xnRiUB
AEORtyLOb13qf1/ELqLOud9eqF2HpJgo5RWYyGPWOW0F2HVk5b7uzY5LzHoN7buAsSUVw8d5PEeP
uSMPZk7aIR33B0fQWhMP1jPeyZhhV2kcXpnG8HhxLj8/gCGfO801RdzD/feiK5TCrJom6NehSkCJ
h3JI6AXJ5TkqTJEMD0iHAWZ/yeLTWIIheKbvtW6UlKYC2xtLp/C5NU5UM818ltmzIUzLNzEpZfOM
B3/9h2CnG2NPTQisVefjdZUIO0kkqrVGvMOMp1fmVx8SEmONgVXYoWAUNG/yfQtUSQhq69XxoIqe
5MA2/HaWyeOlV/0jezE5M132fbafR0RwKDJAIm22/d/Va0tzinrmqqKOGEQdGGZgdZ/ANwmxnmoU
6oUxASZ5DzxLELHoqY4guXG4cD7OvbV6KLQTiYB1YgVH/jDZNuBQJBLJnIajOiO3H9mF+f85LuDe
YGibUFKoKt5Cf4VOvUrbWKi+Z414SVFEhVDcpUX7kvrZ4qV4+gyKA6lrO0vzYrULVC3WNdvCnkHW
7rt1+kYDCX3T8WG3rTvQYvLGFIP+CmlaDPsi2XgeS+mJ+Sb34PdLLn7P5EYM1WiyT4I74fxHHT2N
xUbWaHJi+85kx8dzTNL+YeISq759NPO9uBB+OGNTdmP7F6t1Q9wGtnluBWzjGivUOUQS8f+7os9d
uUko8Ex5cPoe92jW6yvTQxNr1bZv6p0CNaTcpou7Ri0KxYcuBwcPrRa3iwiFnugRgEuuDy0Ovylc
ZFG3Nn2EdRwFd0JerLpibIdOO3qC9APKxDCHs4s94IZY8FymKabNSpPycIkAgEnChCOUQ2zdCr3D
hd4mIclrwZoIJuTLBWsrv8LWHqzfkghkuo4WNNxHlanIygKFgREoLpANobXRhx3xupcqWyCB4p5K
m4+aCyhaaFF+716j32tzackx9XMFEz3mcHvATMH9lHJxFViH1Nl7ucb+AsaglShbgLOhcZD2O0FO
NLrO8ulCmkx+A1uX2tjSxuU9X9UoPekqDr+/c0yUofKiIU9Tvo+jpMkbkotU3O0lePagLp66L79e
ImFlsGxyD1VUtW23UaaJC6B+N5NZ97K3npuyMiWi0gFOKptY8IFgb5Z+A5fykaX1BiKKJVbcbXeN
2QjYyMEL8aXNgz6vLb5aLikp4xVZAG4FFtLpRR/HoDHDaLUt6LSrlfYHCrvG6d4ohYem1AFVaQWR
kenNmy1HMqrUvT0IaIWc20MSE4+MWRF7a4EqeCbiuss6eVegomm4oGhALKq1M8kY6NI/ZlqMPSuy
83RZz+KAUMnahozEG3OTXJGmZs2ZPTldRvyEtgxNV66QbJUb26x/wcMFyHT1O8mnV9GdX4QBGLQM
8NEujGZ4lZUyOXXtiRncFq7cezZbbTkY29zTzGEFmdE6N7VblP4BaFoPnOTjoOdKkUT4EAAcXIWj
l+A9f0cE9+saZ+AqYk+lf7XK3SAkrArm1ikwWiWrFjBcUGTsSt6ABJ8O9OgyQMsWrE+ilGDpjbOW
lMcPcRjxJXxcNK7CYNjsWme0Y2fFxJKL7mg/48hngbqm8YekP0dO5AGZTdXWUaFNPZPI049SNMsh
zPfBH3J/xkbW2hdvX2RmQl3pzVcV3XmYubBrkgwQGGXk5T+eEh+FRugT5DtGuM5xAdR42XXIqyZs
hcsEr6QD9Iy6i5nLlveLE20tvl7+qP0+jacaFVLBZ2wbSZsYJhAohU5E2FAUgAA1gWtpmh4k+wVQ
1+I7Kdd1qnsTQVE8NdbEBk1b98isJAqc9msVR4hCFXVgduhDiQxgVlzYoKKU7GaG5PNdZ6+pm2zA
7ISZC5mlz05hVU2TpEv+V0rjYtmjTqOb/BHzbmTFuCdxtDHZCpsTrYS0XPOV+7pWBgrm0rn/zWOr
7mAyjUaMSGx5D1nWwJReK97525+NTpz1OBXfxDmXdw86vZ3gkAl5QP0+6uajrIE6NmZr91W4A7Hw
L5CMaeFANyF58+YIpHBKJJ4snRDDEoWfWhRtgD1+NZ9t7caB4oq9mUKvNMOQiOsFQjbZD8jVoIK1
nTkv6+aEu8EdctDcv1aoiPbQWNBapKbNUwvfRa8SxD4VJ6fzz2QHM3IL8ckeNTzidDXB8Mm+p2nz
RrbSjzfi1n9uBjb7qLFKgAtIeycGHBIw3E0d/EAwcTQMpnfg6aFAlZ6PrJcmFExnyaJEvyMjvE2E
didMPrKJsUBoIE6YRJgITZ3j6DjK4fBnuiU5Q1vqoA72X5ZNu0px6QSgn75Xe03gmX5dsfi8AQyQ
1Q+BE6fQ6fZgnLUok3rLJhftLAoME9LtQ/sADy114Funy5tP+w4sUzBhGVfSO0tfJVKRkZtUGIXm
f07OKKmx7QZUtbgEic0BdrfK5FEp6HNPZILp5/ukLgzACQ6htl9CMfP20UaRrInKYRky/M+hc4AD
Llapn+OH8dDTLH5Frjsx/4BRDeWUWFNQPjwNtyZzSssHZtmLUHy2PmcxDVIkNzHSNfERGADdMdyF
z/Ajce/14HJ6Z8cF07uUsQX5vbhaYC9xqyTXGgiUrxQMoRRtJ2p4PAzbw9gJGscmun/Hy1VfJZlA
S/7YqEWzAkjMN+8DQW5FLdHQ79POJrEsaBKxdUHN9jSo3eIdwR1rpEyQr8ZoF431My5L4N+ko+jA
jWoCO17fqDW94KFHl5q0w4+8p7W+QayzRy5DLI+fVZYPfAGqMAmvOpkpW3CpLIVXbHP347Su1+kt
dAI+JbjlH1aB265h+nSF+Sdj/vHbKel6Df5EwKCJj47oBH86vlo3IPOXQpo0pFP6UvkzdqZ96Ypo
4XqI+eDVQSDg9Pf7eo6SihzYaQgm8aO/Ef5BQdgyynA8hkSF4N1lJxjwqbvJq5h6XqEfRj6R0ya7
AhB9wbYQxJIubmYNxHKpOc4sAe/XSb2/Ery8C1mpX1JG1XTzU3C95WRtehG/2JP3uSAFVqLOxMKl
AkXf651QAyX1nOKUGdUx7butQD4bLOJjz5EnRQJxfaGiOamqgYyMKrLrfOl4zf8fuoM8a9YPXwR6
COCcLm6ipNFnh1ORpI7CIkp5+WtJYpUYAj9EiNWbZHGVI+CELKKtyd0dLMtxUM+e2PbMH9gEKQrr
FRWJJjWDfZ9HIKEzCgdVB7zeJzMgnthimHooXwhEHnaGv3h3Cb1RNHM3Bo1tJykFzx1PCl5KUUQq
3xIfA3qds3CoOQsKpM+UuHzAqGvWdwld23VQ68FSY2/+ZSquZe4Lt1R262S/lnRX+/+keBbbV8TW
whQkneapeb4HxQfvcvaiTedGqo8NVwNt5Rvj5SgPI1CiZYWysECQGZzHPqMioeK3UteuMSx2r/eW
LjfGoBN5eyoSqqATpu8Hqb6VNRIT6x3gjsAVycWfcgooaN0J4d9qNPDEdO88zIrEaykbfjs3z/dc
ZtMmS9GRNdqSbxB0UwYDN2U/RzZTjPLtya0v6qiXBtiHJ//FsSNEMoBHNqQFyLCXeDPtcpsSYKK+
I1GIbhbQ3GXUDIi7Bi8XTlBIKK4jTLg1tCsQHsULGZlIdAxdbF6mAm5ANW8AHdh5tKSDtQDYfYka
fYj98G1acP8xQizhcaiicEj3qNcg1A0gr7+CYDLaDR1jGxSLrw9kefd2sAJHvPP3LWzFczLMxRrL
RoS3QzkOxm6jLV5De/+d0uap4kP94IyNNAegd+Hjt3hOyxIiCZNGroevhvPSuQ45hkxWPn6/11TQ
le4n7ajvQXUanS0CFfg9IaA7oHAryFujYbKMSAAgJNTKt2f97sdAEggwnPDNgfnrjnchnnuLUKN7
gRgQSOnxsSEmbw7DOpBW0vkbuxJCeWDDGv+yJIQZJMIxzgGNucAjIe1nNnRCobSuT8lnjoLymLZ1
ViX4kICT6Ec84w4+X6WASHXuErv16q4cKNktuxn11W8KV1IY9j4zChCZJs+wLjKEq00VWcvH0KSi
dr/KhRI49eRvn6XAV+qnJM94afRNpPwbKwOZTDwpDSWL7hx21G2tIjDTftgLhz6+6W1kW+1BGJhA
ToGYY2jtgbCllmo25Un28rzks0bGPbNuGvqxeZKuQdnozvzTj6gVnQyCy0j0yop11Nb3b6xcRS0g
0EKrCODawnIcYcmqtJqqLMrplJ3bjrhsDbM1bXJUDGTnJuoy2Qie3qzCjAsQBiYRWsrUBhAeXzCa
x0XyCRBUtB2bRaQSmg6fK1x/suopnIe8i4p3p59gbMzD4D5+UUzN2a4XEWrONeWvakGFnF7uI6I8
QoawqNorktmbPp6L7N+3fVKJxufrwYxPdNPXJpn1CZMZyJ1K4vGijLHWx5ySXgOHMh19nu2t/hOT
LofUVI2+H/kiBAABG2UFFQV3E+Pvdfm88qnjn0LAEX/l+mKf5gMnn9afdM/F1Usm8x/UVRNdPbhK
z3XvWVq5s+w5Mxeq5JEwp/rCIwoKUnCfDTlYWqYMeJ2ofS+SK8c0bf5MBTkE4Yr6d5HBo9/qmWoL
cn7j9DySajdGzgPrdXAEYkMMEE3bvipkbQdsTTThpVW+akTYl5mzM5phXLoRe6YsjNq7oY/CjuN1
epDf26BlpgWm6vULA47w3EBtS4b2hkjGMeobid90u5JC9TNoz9QTAmp0ICbJJ049wedgwc393PKh
scBOQvPtES9PW6Pm5j7rBt5yNC2rYguYb+oYRklaFyYpjd5Vk6YpyIXFH9the4wB/PGlIpq3PB9b
fSdOj2XsdY/bQEF7f/qM87yqbflT8t2o38gntWZr70Tgot2U8+Ugwd1dh7Fwj5O/VIHFn8JZ/CZ7
SxYMJ7HJl6OjMXo6FLyPgBYMPBmHnug/+n2N0i4N/LXUQVafwKc34ubYnWu1H7uJ05NzqyF5xLt0
+oAEXgLM4rjTzuhhjR2GYKee4B0kUex29PCFZ105VliPl2T9OLIYrInZxhkJDsBCmgqhCOlIrhZR
zmUQass6o/EeLSnmuCFLY4a3BNd3wcXJaFOO/w2C4j4XdSEALjjipaP2chdZExUCT93NY+7xiyzT
UFelKB1rPRGM/KlaFFEsZIpX1kpxydl0LQBJTTP7HQHZZJ0kv4jrNIafs+ptRQitVNwW69ytN02C
EXP+RtsCOMcFCac+kwVvAt5P2AHQilq9gY1Md6NstmLitXK6coGfJSIF7OK9jmuKq2pxvaMgt+yN
lMGie5Qp8P6Z924VCgiuxAw2rUhHerwxm5xD3EUJg0qSVWC9Uwjjk3DuOIXRKdB7k5DlxKAeLBP2
SO80Y/pAIX7d3vXyj6UkEGWV5rT9+i++d08Y3U0PKqik6U8N6sGmiLhkNObjyBfhGock69AahBhh
gDO3NFWY7NcVpXblbZG+GJl1dZLiEhOrep06vLZwvyDhxTGyYbJ9twsu6uEFTS0lDoMJT5dcW+mL
Dbe9j1hMPcp4KL03uaOHSbUudieY5soDG6BBCgVGcXmFDS6fRvrTX5Y8n/Kyn9C1W72JJ4H+Q9nr
7KnnbHG0OOUBpnkJyUqzVdFiM0UzAPky3cgX/y3B0//OlwfErXk/v7jQptuq0wbdZiPxqvq1avxd
EEF8JEw8QxitvwEftN9+1k+Vwigh2+YjG2ahHQJgJqiHGS+aGXgjeI+8RJkqDBNrfJvNAAYYFPcR
pW/QOcv1d7twtAKksUx6eXi+iuyttg/ANV1fcY2qKHouYtJNZjBcmOmauZ2s0L4mF309YevK97Uv
iw/qKoH6y+2EY3OIrhZOzPgQLFFN7k8nVm9RviBEuP291LCGJ2ex1MHgjN3b+/rXFwX7wwRQoCNE
KHX8jQ9VDyWAkU3So96WaueQMWmVA/dl2TaceQLk+GJWIZav+M6rbBLMTjAxp/N0pXTcbh1jX/Ws
HeKOSgAxcnwMieW/N6E1p566boGpvt9289TOpFyYCau4Dnu4xvAJxx+Pibix0XZxXZygIuHZbMD/
X/bNm4eErDfRnaRGqVdZtqJfpz5y7tKS1oCFmmTjdy6Rvlnt9ZEcEpsnpbn56tWWtKjnJETaTYYd
2BT4CMF8H+MflkS17fkThCW90L4XBaoF7e+HKv/M2mKGxuusM8GeuS9yPqeRWH6VNYcHxG4Qoup7
R7xu1QQ+hkYDOnR+B47fK40WhMtqcCp/2jo7VvUCrN2RYACl5umXZwwq7NNDU6hi2Q8vNsfA43S3
VOrvLBldLBCMfzqk4fzoTcMn5tWlNMVnL2NiFqWsrO0BA4aXVNDVndl4J3Fh6TiNW8kO08RwH7dI
z+JqrcLCCzVo3dCEDrI5ycRUZcxRdHIt8kwnuTOZxIjNfJ7R3/2JPFd/ToLpdnsYNCf8zkl/NUHp
W4LAEXMayWmiTFZVRnBjJAiKqyo+OtMLG546r9dcPeo2j12pwGx5caUdx/ERTb5UNARsoYa/yGwR
oDcRcJO5NWKzctmtVbld5m7vvk2ZXOQcaYvgJC74FWxdMLinyxTjDvN3m2tCmHUAKE9ev/wJCaPq
rrCN5Wlgh0rkDWtSaFHkBhbsrTaAXroZGWcVi6S+DAZp1fYBtCs+tJ8uUKoWEo8eAjXsT1rQmzGy
3kzFgDzrrxfmi6Wyu/gFJ8kdgNHrfCthyj4hzz1fThyEnExrfXWM0/ZCuvR0MDH8SeWssRVM8aoo
fknwczd4PmDB6rp/KY1bvQQ9Tfddya2X6giG0uOADYkB8DYNPJ4tLCqRWZT/Q0fVuhm5jRwc5UtL
yDwXiJtiJR4/09UQCneYETrXljAHD618T6EkYKCj/+FOq5nDO79qbBXNujdng9cPiCuRvfTftZKX
33jFHw8L12EzalSQhp2FjCG1Y5mHUWHatG8IovFAQ6nNJOtgSWib2QKsvi3DIFUq6kQa5Tq6g22x
gY7fClMOsjDW2O6/uTQuCAiCTxpB4wS4QpvBEhmqCRH3pLO72pM1aOTEJB4P8p1lRRsCOPQ/tT3h
LOElZ2goHRtJU46elKGzJgKwyoE9ttIP5zCn2v1vzAp/yyzyfUL67X3VAyJOx1kcMgkqiG2Zk9WQ
YamR464gMJ8pmXYNzxyyl9Zhcby0P8XJGU0JNpXDVQeEIrA6lciQaV+W0jhJdJp8OCwEHDz4jToF
SZALDK/rigLTscPfnwt/dwR8U4Mxvym/0MxJN+yAXcJkcoEE7SHC8kbye7PKdgtL1zPWWz+1uHIY
XTCSi+KFr3pVePMGviItiIf2HLbYdl6TNHFYwMiVqoykujwbs/3YcdO4gBLI3n0BRoFnpgP3MnQr
vfF8/dutbR4ySRO7/lQzM965+Ofzb5Uk9C5eWTnafMkD15xpcbKMuCAD1C3qw/jfiyAErRq77YtT
orYI/ngv9fT1CxKSqXEaGXDlSO+gPlHE9tocxg0SVEmpRIHA9l/5dUf+2b+c3BnwpnE0jASI8n+R
cX79KloxwV+o/WV+MhWBgzqTXcGAOcUSpvUU7QDas79jH/TcWG9DeT7JFRqTsfoRvcb5BOBm1pyq
XDy7DsdowmpKEbsGc6HiaSV2gwFl5AJlOf4H+4wYP4yExYZtVkGo/Bv5D0PYxoBdakXJUPpcFQXV
Cfrfwn+4uHAQPF4xqd+42NKBZv+iHUQYF76DA0BaDehZfQJdJnwhq3Unf1okpC6LlyBFl/XUMo3P
0YFhD0kg9KkGAYcJKe9s+08blYTky3iH+550vvrHxK0GAxIG7daKnMSGFV/mC6fGEl7d/TdUyshX
e1x/HDdqauUVco75MAzAYauvfygaye9fG7UmFi1iGf/k3/xyYOIIrKHR8DsHMOROD+IFH0HFNZLN
ieUOHoAi1LBWOr0eXKHEkqRq0+IYxFicfu6bBMYCSoU89KqRG+NB/Z89HyfqUeYRFY8LPTXU0lBM
iMbo2oXykSnJ+mg+BJP8laxockyTTmB6GwG3bIY+0vIWUZwZNOEMsTr0hsLd0Xbfo/RH9VAt6o5X
3PmTNgmijRcCf8pNAS2m3lKAaPNDCguSnCURhB+z2x3niy7onQYsEimIIeQVENf4P6YoH0nt3f1Q
CBgBFXL6EckEYgsNP1Ry4TMBWGz7y9D2QIKDJKE9Nl5eQp2tA2lMJ+VCnRdY7hiD32WilzOQwVFj
y0CX6HlW7Z/SF8aktpgr7PStHzUR22USrkBfaLAU3ilGdAVdoBxMEzFM8m6MK+Uhvv+foEAf9q3t
FxNujc6CaTLHOn7C5i1/WkUo6kOUgMdgCPrsN/3UjRAy/KxcmPjz0qmspFIWeXJ5btpmCxdts+xB
G7ptALGhmnelvDzHJ7VvnktB4Fx1pMiyxg/vsfVoCLX4US/6JEfML4IbwYh//ytfqB1/2/jB2lWe
UQYpaA4AJvlce94x9bRuXqZZLEsuAJ7rcwdFHjhy2gr3CnzMwlNqjff5tViSqOJUoQr6NoAIbObQ
pGgvnxSZr3RgD9w916V1K3JzXIn92h2FdGnuzfIADkKyX/lu0SXCa8tPveZcRJsgToLtuOhfjSw7
gqfWJr4zd6Ays/RjurpTzgeeleTfU0YyP0c9x2Ql+55aJPHIvsxMUbXglbRwO5+EFQs/J0NJUNNg
MlIc744BVSBbgNBhRDHl2nCoF8WvHpkuXHF+ilTnALBuafyHXWeBn+2y5kXCTH8ZORRnUZLGfl0c
EYAhU6Th8eBfy2cBcxVjSeFN1ZkuFo3glbF2i5dg42vuDk6s6yV/ybAShQLwn1GISQkEhyvBbDJK
DR+vaqm/zKiow7NHOr9TtNOvDDB6bdh/vaLG+pVhAVW4TalcNe6WOIR4TS4vx6DkqBaZ1V+dz/5j
5utYPRYUm/JliRaSUYjr/xzj5HGyjw76ynjOeHxnam9s0dgbm5LMq8ZDJzMN6DzWjC6AMQiFmxqK
/uUIPQDaa/kpdgK6GsoBhF09Vd0j06mrI0c6iypaQePxsL3a9Uv8IkEdRXaTOFbskz4gAxz6wlP4
ROJuFT88YICIuTUSLAEZ/hSG/f3bSIbKyumV9pYmJEjuU5DZcIG2jiq4NToAWnwljt8+Fy1iW0ZJ
D5VRHEiY4cR1UuhkZKZHokV0MFLusQBAtcqkcvl/MSfm7/0bG+2cHoy54HrCUFPMh5Cdx7ubGcMn
1bUTEuxFd/BdHQnrsMi0xaWHMUsq3aGUroGoOzX9HZ0TLye8DyZrz7WrOmWgRsqhBzF5vE038dlK
4tX/TH38Tpx0GBpzdWc06pdrqjbo57GDXGn5/YM8r5lUPL0EWgWIEZ32HQR80N/MyQ4tWdgL8wd1
VpaurNSM6FiLjoQ2vmeGbvHTbx1W0xSFUE6opp4qdfaG+BRgwrxs+BLFeftZyZDnnjX72HN+JGUe
XdaOKrqw6GvcnEm26kDOGvCI/H7qjC/5Y0wclZ6KlaRWoBR05HwFRDGHvl3YZHzptvlRYrvZcRFa
ETuOuWrll+UYvVJuM0Zm4PzzfciwBfW8TvJvHFeyOxOccClQmFJM6NlLE9PRJGq8P0FkLKHgtJOe
TRj/5syBhSvjw3zbk7Q6QniJybbcZ1zeM6EUNek3MoAgJsZ3ZjJq/w4v3yQLya6UTxagnBjicpW/
6dB5jhLXP0yGOTt1qbjLH7xbbh8PbKXu8wrtL1KETUhc13OmjGBpDcuClu1wsFE1aiduvyg+RaKa
m5AhFRqnNi3o5pl+tiZbR8xtVJjRg/D4xAj8alP5A7HInt2cIfvUWpYMSs8U7mNYIHgh2szvYucz
aT/AxJei9UzCTV1VKnt8p3GpYZl8Jq8v2d49leV7JK7F2okQvZwHnwlEfy6fGt6QFMNNUx+KlQw9
JRp408rJiPIk1m/1x6wfON4oyFuWUFKz/fjGXCebUvIaXwZsPCl7xEZkpCpsTaFF+Mstq7bt+1+A
FgWUdINYLJHLkC0VHesorvAefNGXxVW93lysV1mzQDPebV6Y/56Xh1DT1EkVWEEe9bfYKR8bYKST
5aThcs07/gTTX0yW8SbI6ttiCX9NRjtkPO+3lZfl8hA+qIGrA04jPmMJYasUwBxWlOuwSsDCkIfw
veY47wlBXL+dbrdAFBConL/gYwtUPk4uveITfo85eVOdTk3YDC+eVIWQziSncSKhTBjFtPuDzLH/
hUXcjlk3AsljihgZcwgQstuKsmSk0ixbUy17cAsiCj2cxHWSsJxgDJ23ZusOvd70UKkw/WZrBjrX
3Qh5jn5ueQvdzf9l/bZhMqdpMtZ0WSXzmHUV8eSrVZd+oirlYy0Oiaa4EN7SDJi7UL5kYajMlUCq
IuxPPKElvh2S/W4nxIWI2qqzkXrPJ5sPZlSf+V42+ww2E8vFU8l+mgc6bMjyVnmVIC/bsLWuU4SN
Lh/4PoSs08+VLrRMIPrtwUL23EgBhVdFoWnNvWk2Y4SwI4VPV9hJn3eBVDHI1MLSJ/mqMBP+aJ+t
90XeM69XR/WRcsF4NtbTNXJQAdW3PsF1FOfObqPhKBodPrm1Fc80tiMa42PWd7OLQwCxmmb+a5ib
8DYkxGYI+VcjvgY8M1Z/p5x5f15qU4k4jtGj9jDDNDXhLJ8mkXyclER7X/drzuM7NS2ehAyt8WvF
0xFSS5OeLOLqhlz3MztUXNXpuCSjWnjldmpy9e3yOAO/CKHXdMaQi5PDv7vPXXEP56K3C4gIL2wp
jyid6iLTRxihfxh52G/juF4SBbiBfZA21i5s+1KoqxrPp/cRnqcj2El2Gl5rtyNpsVU1KnOk0Lth
VnQ4+jCrb2yN34Hnhhr+69IBOwuPWgTjMsXG2N5FMgPikfqwf7ERoJ3Z2SnalphSRQFN2pzFDIvs
zYqBYqWZvEyZQtx6fmuVUg0EyHVqs+9mlXqUdhjCkiqWLe52u95lDUhk203/p+21GJw7AR/1UYOS
/Oe/af9vsEavReNjs7oteB3xENDL8BWkrfMNn1i4JKhSz0B9dbloWt/wJNWER/DnJwY7wwQObBVf
wvFuGMN8AzkY6S33GXJP+GNwHeltb8AKQi09gKIHD/j7KsQf9p92L/sdsnLw2Xmk/Wvx2Nu+TtTI
IhFG+c/O/2mHe/HBcwSPWt9I9oFQIcrQMpATH7amNWIdyeXo6AnGojR0TDG4bweZYwmMFyBvPSYM
sGSt67NELwVaMPz2TaRH7VDAOLSP5UAYK14C+3UDJzBN/Ksnksx+ir+Nio/yfFtciC+UpVTi8cvH
bdJ0+rIlmXiSSZUt20y+w20BMs8K4YKoSW3Mm9nikhetqpQoxhxurj0iXnXCg6n6Jljlb+zFyNen
j6NnLmv12hbNukEK57qFO8Il4u1aJDmgy5WRe9DH6/wp1axt4XMUtlp7f180PgCB74rkGWmhISZ8
0OQs48zSurT/JnPD8uaH6gLIMhUi9UrlxvMjJxpAq+1iO+sjpZK2/5zW+rdUx7VOJGpTntxcYUzL
NF/A2VAgoGl0cQAWQOVRc3a+oBgC5QFGNYiXVwgL8yZyxSmtv3c+h5lsS+GvQgVReOSAPBS4sR4z
n6MID4c2aOzWSDDDvPsoy3pnnYKDuzVw8jak+Cq9M5NUECXE1u+kzG+pw5hBCErFkEoFmgxBgUCw
NmJ6CE+e0s5lajdN8AW4HmCD1QNVKSW4W14u1NM8iYZJDVz9yVCva4jbeLG5LMVsI13Zp27DzsXg
zeTl8EzAzT10hO6WFQYJkZX0ISgaFj9a25wHcT58TCBGcf5afcNVZJ5KA9iDSaeoElI94HeDXlby
0pJ2b1cMYx02vDPCbtxU2yw9S2gM6uVkE+hJJiQJVpSC5uAjlIY9P3cVEg+nZuRlxA0AY3vjqqja
q5eLiwhKw0wgrt+YUKPLrnBj8/8svxRDoLBtsZiTx1NN9G7+buA/nc32QcG7bXBY98wwq3ieqFWE
HD2aK6oANy2WQvPcv9a5PwTa9HIJ2BCdbjZ06AMO1FkLX0Nbk7aKS8WT11fabUZ5a6QhL/RHyL5l
bslLcoGjiaA5ktk2WBGzK9Cu7OFMhy2t1lPqCvyK9BATfs/MgOhH8oxlu4JKge5+xNk+kEofOqSm
WIgxuL6X3lY75xvM4goPB5941Wif0RGPJDZRUyoV53xOjZ7pbwSCPPEOKCKb2Mbm75XJgDDC5m7J
sfSWbvrPQC/FWl7svpTsow6ST/KRScsX1+nSysDUWFQQMdyy0c1dNm7bZrHWebumIE5Id3XpoL80
8UuazXrWEWmuYGBPdBmt68hOetVdDKbk2a2nHl6PhDTVTAcOM4MWkEt13TwalOa/BdW5nEku52nH
LgAOwRArK6KXIqaZg6G4mKlDUf2u4dTp8vC3mLBQu/oELhuXU6rbTYRv1iWjW+r2vNu0ZY3pfr95
I1jOCYJY5aj4jr3Xqg40GMR9DzrqAi96WXu4cOGNumVmXmXL2BHNjJfRX2pfxtffnHZ3ddru3jiI
3YA6UJtt/mKuAzkCFJNrpkbIKvXshsgxaChoHW7d7MLBUWXOxuJFGOEcx9xMYcA8KScdAffiBAir
g03MRsb51mHMjagwaO36TB1wJ+DhLt8pUgEh8wcG2L0aedxZZACiW8zDyk3LBS3mgoXxfKxSvTKR
GTRP8kCWzo8/dp4uop1kaA12CNM/aBmgPxmfEBYOFCnm2DDU5tIY1HoRXM9vEYTo3BTkvH8M9ni0
BqkNSpAIMZhiLhhosEdeDDTj6xseNGLWKThpqhppR5MJJyOpntmEW4WV5mroH8YHMzvCQzY+vfzS
qOzVDx26+XwHv7EV5WojTdgVdPFh65Ptjvj76farzQvQRewWr12znca8AwGigP+Gtgoxsb65/tJr
tPzDOHmoyYPHVqLKFJ+0iWou8FLljzQpbPXdb0Cka1VZrvtl2eRmiYp2JDc1ZwXw/xRw8KhzyoBl
YQFQ8mrcl4/EEs6KOR6Wo81fFc4tqZ6xYKBGEHXh4ciDiEysfzRO/BAMN25c0X4ldE9iGZk17d4S
COtCI+ZsTffN4iOyaRwZ3JXDjOucu9thsGjcvxE/h77cfpKmk8lUJAqoN2GCAr5LuPvocBN028vx
a8l4VUbGfJcqqPShyrCkAZoq915vwRYWVE7xE4vCWHi3026fb4m7d1U/XeOHfMw0Hkt+hxXSA/PZ
PXTsKrMVvFC2cCzOu80aNNexxxhVhkj+hXzUPsURczDineC82q9tn9YG/JQBt/TZ41t8JK88XXKW
WB6I+KvdT0ZgIlYAJ9GtIDNUPOtVdKovFlhAEzi3NG+h95GOySTf6QD1FAG4lMkvC7Ag8LBp+Ojl
HY2hz9xRXJ8u/NDSsvijkKf3Xn3lJj72g10qkfJToXc/EFiZaC+Edy3Kva0DjnOcGuW7m8na4V5a
8LT1dMRAkFh5lVSs63HIVErTM2GZ6vWBoXjkyNLWapfOlcMcxNCRcfh2ZM0ZEeGzhZi0Rdc4qlvt
sdo+83U+Y8WHISA1XyYuH1fmC/vyWrEXJNb5BaQwUqvdJPznWovwvaBDYjRhDN1gSkUnhLeTdf0X
LWmKNoZaJbT4Jxaw4xtoofl4VOpOxTy3Ud0czOTK0jjWDBthE5j24qZcTYyKMX5ZzBXGAMg62P1O
TpJI6OXPHnMqYQY/cv/a6OPkeslU743yrwS7DDgi9gLHKo7/LMUecQZ5VkvefiY5KfsUFCvvF5py
ZzJxWBbbin0GymHLzzoLZooaYPe/eYkn9I7spgJabftjjmWIm9dM0Fn0td7g09iCDhAaJ0EMecJz
PG3euJjqwGAVvQG1CxHNt0zmOgPNSEB7aqoSSYdiyuINX8i+0rKJwbfCt6H+2kiZwl5iWjTl5xhK
CSjjzkMCVfOO4TrEwwUTiEzvH5kTUg6prpzYbQOKl+6PqCZdY8FgZKatS3BxuN24yni1/vo1bFf9
mhANjJkviPuXQ2MQT1LKkhL9QjmcQmbAL4n6MMm2QADCkwNGt7x0SUDkUZ2NlWhjCpePBw2HL16R
rfW1WPg7gdPxRNhrKYF+2KfbTffLoQgaNFLZD2siCn+/+xwk/rMPgIJkRvgMKXAC5eEXF+p8ZVrB
YgoClQ+ZUTTMEBXvbnWAF6nuL6aXtJdrCW1Qmho4mBK28mrf+W33DrB7qgUiPeeq8KDwF4FDoGBT
vg8ldLZPntDUKVhVeRhb3EqdbR64iPgKH0C+/dJ467K9rK7Nqo2qsG50ez3Z5QSy5dWMu3spzXNW
GF4CJODc63oC9G/3Dnhwl15xmUI0OC1/pSSDbdVGVQQLG3oPmkFZYJNGasyr7Bf7oLmYr/v+kSJ3
nL1iBCKslBO96Xf8+7P8t55TOZ7WeaTTzdrijnkA+96RlOK3vUfnI+ZUiyDVoJBxwY5i6UjAAPh2
tLJpya9HluAv2vUY6LqLz5thAqyeEC3PVSa+YijTN6kc+J9kV6yTSukLaAiEUk3q2vJhjsB+gqeR
DE5UBPGh0IHz9q090wIl+F1ZpSYvCxo4xvTdIShNW4T+NNfobeFkNxn9uFCmOgBn/R8KTIhkL25L
/izJvWqQeebgKQRB4MzEVV5kU071JxrmmX29Ba8uZn137tRV2XzfBWuDYhJLHpd9zI91cKggdSaU
G1+JEut+dpO4ySbX7hpr3o0QOPfP1reY5YMRg6+9/fCL0KMnMJ9ol7fVG429YsEQLmwFOodLbJOk
lCWO/7lk9bGqQBZut+QZapAVQ0J57dOQTY0IcqqkOwB0vvTMiSivtJbRi7amMNdcUGqPTdBUMu8l
PrF9E6CKlsJbf+4iym0CrexU6ht3SnJ1+JaTWrju2J0ZeodCVo76LXDXmb2OU4xuJBlj1QPeR71w
SPAjI5+fbF8+6DWmn1kJD7bFQbtwL/yRPUHjmmS+RqyrjeZtVcLIAn2+77j3KPsp4ic694AuWCjT
/T2aCmByCxrpe+8s//Dv2y139+tTNWgCRy5vpRBTP/2N7TDNn3bTY8jUjhj12OgXDki0Dspn68IL
D6oUWGX1OnWUyaKZNfXn+/Tf+PHgAIMZtouwwbgmHRgRzVD9943JVeTur7j0fLkC967CyMS4vk1/
AQ6+jP54pIbKWLaRZLhARmaTUG95R1EvaJ1wOQAVdIZw9I8XBrGfdjqj6sqN4BE/FYrhjAupmTui
nPU56YQD8Mga4xM010q5KJazRD7e23q1diiHUnhGEqlKy5/hZryHJshnv1Q7w6DbOFcEoXftcxC0
neAKZQ3DafIaG6rubwW1b4YlVQy51QUdEH+xsWYV9fy6XIF+/3uB2akQxgUs5ISiRsUQtBA9983L
TgHph4r2EG1kBK5CynG4CmE9sURl1sj/y7lbmRIbuossMsxWuw8CGH9+ntGCaDxrOohlakufvOyF
TtUdEZJpRTzKlNRz0MLEsidn29SKUreisRvMeatrqMdOfmtERp5082fyeuvMKxk+YpVvfn8gg2xU
ZA/nNFuk7Cw6M6MN31N1FJvgcRqs/LKE9e+vr56Vk/p1jd1Cpq6+LtTlSCxIeeDjHXyWzYM96KBQ
wwnqHYrVQXGAs19BUpeob51u8h+IYodoZ14zp3k4g+LtfK5y3MlfJeJXwe7wek8HyaVPXfUYL/Kh
dBDl1WTw9sL202hpyfzkyaMLF4UKai2B9LruZIMb4c3L64EEHIR3ojN94r7AOC/2wnueYv8vDVyL
ubqTEXvyPBs2Xk6NwL+DmiNHcP+K/FhE3zvCaF+yVocUucdef4y1QPqU6zJ0Ts8Gylm4kNcgdqti
rOVZlrUfMkdgXDgBiohUeEthzyZacCza5/zXxxO0Dxf4L/ZVjSwlcTc1rpeheMy/eULE4xSR82lm
29v4VODu7bJ4SzkdiI9B9mR1XIdcJjRg+JaR/OUFG8BxWWHLqL/8dIEhdpiOtkVLl3RwMUh3pM3R
BL5YMSyPPglPtBPgtdjDzsVRD97Nk0OTm1WpwT1RARWkINcPq3urSC/Y0PjyTJXwjWWOH/+dBbv6
8GUTsKaFPSY0Qq9RJaiNCS5XGoC+bZwRC+tbfkD0+SJEBl1sb9f6kHhpUfLI9oQIRmWheFqY6ZSM
fd8uJ2giklo1WFLz/KSCDu7JLe1OtGRo7PJP2jNR0YIJNVyPgD3HrYNivUNkLv3dXAtAjiL60bzz
g3zezqV6Z1+AP5nuik3ux4YTT8A+4tl+unSFuWAg7NmGEUZ8PCkwud7lPpTvOgbLYKKbm8unsJV5
XWka485GlsTLWqVzvco+T32hyu5AFqleD254Kidc4RiTUWlRxchLQ6j8G2K+jSSEMhTgwT7GxoTk
ErENTmMI+I8Mds43vWXHwqiC4lozs9R4XiHl+DXRZ1XbH8Kd8h7e89QeUkqdOZpNKAY4ydtCxXk8
LnS7Gpw3J+GIKjQdUzUTIt6Z9zRrZS0npK7Y2aUNSg78h8pv7vJgGd18742xRuDtzJGWUoNDV+JG
M7gyCYWco4WSl552eeC6Zqb7UBATq2qDO3OCRJADhBgr1WcmGVcCGUMIqSQqWAcdNywbq4cX6HUW
2aW3KFDNcqtLkvRWHmtQ2lDwl5lDY4jsJ0NCEW8/nR3N7QSiAVQ1WTXKgrrlI7xO0nACr2J0K2xn
sG3wVg6RNXSpaY+qX/LlFHzHvyRCaYcC50+v69V5jz+ExJg2qp25Nk8jayHqmN8KaAUGfMfnUrW+
vbWimCiGeWqoXtlIYOOZ13otthis23LKqIhNCu/aG17DtDnVYeji6Ps/Io32jVdIyIrkxOywWomP
uHJHkeXym1Qka6YQyca5ORjvqMF+N2UuOTVSsYsFJUknCKUZzyHLi7YFh7+dmjEbnYRfhr9PZsaS
sEmaU5GM59XB8jmMPyY8gsqUIKTQKWCtk66+y0mIWUgiXRltxlXjGcYsSqxSnDFhCptGDOCMYk0I
2G8kONHAtqDT0+oWF0DNzhQVXG4Xt4gYUNYuFBJdrDPcf3xJB17CK0XWCpkUeH89xk9RFzy7Mo6G
AFd9xiNH1xRqAO3UIDEcAHHjwPP1tcSuwAb6CR5r1yAp0MKWhJiIT/xLy1oXAHE7pVnL8SlxIftH
mH1R3uiQqdseeR64IXOf5y3radFaQFzVki04wsk/iecpavItQ/GKaYAbCxUh5RHkkhpn0jCVHuuJ
PaB7ZRwn5U6sk3ohX39XY4usvKvy2b91w/1IpteyzuUZIs2Qq9EtJ0HhAfm8nkRWSncAsQqrYuqX
ruD8ottp9PFZ25/Y3aFj4RNBKNqNX9qsh5ulxFnJtXEgcQEM9QEKga62K0cL4+PmR7XxhP8+YXQo
qKiyw7OLUIde2xTp4YPnZVjxQWY0B4lwrMar6l/s7mouMQrUJXwgk1xVut8lQ+T8VMF2lSltiOsz
GQgs1jA4E/H/znKINyOQiRUMQCl66S5bZNT8hyGQztQzX8ZT0gkkuzSWPlhj1/Gha7wlnVShNioL
MrgdjFZA1ZJ7O4NzScC3UQrKTEgEl4nWwd1MYGVdPLxHJ6iOh61Ug7xVVjWl0dlkLWHEyYgaYaiV
Id2DJwnhm+OaqJrhnJxNZxE1gkc9t/SAlme/5doW/D2z2iGa/16YA7gTH8WW5cAPtSVkXQNImJuj
J6B1xb0tBCicSbU5Ih2csYK7y0XDDKErW0kKIDSYNMCG+ttqkhuTG2ynw0Wc+Jv40MUG7zZWOdhX
zhZHrCFIv1GvpDJZce57USCKHUAOBkBM8q2Z6XUN3BZTM3DcTL3RsO4ELqYcYSbs9VOCcpEZnAGi
1rQZusI6twkfCLEVyZ5zBPPLUGNzqxuvi6gmXe9WgZQh76Lktl/QSyU+BEDG8qk2D0jARfjrWhfG
xCI+MmdZlgNzIwUtixrWZtOuzHcC6tXDGCJMNxd/OBXdtHAaklUmC88gvJp53jEoX5mKl5smy7W/
7o5hbQDpcdZSx/TFg+Mw/7++zAnEm6PIPBlEhw3Ei2WXxQDbZhoZ95Karv9kbXKvW/X5TC717Nu7
bWwA72YYc65LEbEoHnJkg/x6gCrukDBn0VZVIazKXswosYqWSvWFLk1Q6jE+SUXEnqW2Sm+Wcfa2
53L4Oj8f4sWRZ/7c8vm0w9dDP9VzhtzCjyhQHufSJr5OF3mMbCI1/0q2DxKEuiI13seOZ5x8uMkY
ZtaKks/dYZGwKIOyB5eoPTX04FNpPa252MucrUePssK2Mrkp93NsKkh3YHe+YyPB0MOD3+gVkwCE
JQMRKqdlq+43GPuN4ujHS66dNxulLL27qKiFvAaUyIgpeDyjE2SIOB8ZpfdQX6YtTY0JqruT69ZT
yM95IwQVeXt5D2+jJU1Ii4PX7txozyhqeC4y13Beq5Fi1AnYIduvH42HOoiA/+2GBnaai/Ynqbak
qed2lN+CuJLC9PV+vAAaSCFI2nMsBUyjzMQGKpPFLY97pt8LuiaLWGzIFAQSDQa6PhmRR1LcIpr4
47rVITcaulJjgvAG79E26JvytNhFkvQ4l7ZPwHilHl9JPvxUeWrukEFDgmx/uf6aFSUT4WQCB4r7
O4hHk6Na64e1ZHfSOlkwHcL0lpw0SAaJxlFbdSDstJnaUIj5hGTlL1lhZRY1rc92+pTGsfUpW1qr
hZQDBEurCtfxf2admrcvik/2EATl7EjAW4T1SKOKM4vP8bP+OJoHvia8BimFvhV/JcvJ04txkT7s
2cOY+BsgifOnDaAajlDvNaIgx0QU8wrwl1nr/yOR4TKRpaS3S3g6booWL+FAdnyTAzAf7+LNnZmO
1T+AiNRIQrXIXxfuGAQB7FXKVoDuecUlzri4RiYoRBzePOresQUrIZhYMRlk2FrxUjLWeflcXTJi
rfQuup/Lf4EmQQl0GGm3t45VLhyMMWFuRZEBtAEmSRsVMDXScpLRKSVX+gwI/r8GJHxfhBNsuBvI
kGbygU9QINAtSi7kaWfUWMS/AeLn3F3AXLRtb0QnLZBCteLXBhiqV7yeQAxNc/5Mi+g5IM8CFV0c
EtoB6eOk8vFfktZIxJFRWe8ZonAcYvjTblX9nuu9T/cspCH6C10qjefyw0Z86hAATmsQN20lGDJw
B2vKF6WpW/SLGuFJnBrvcf4VxpfXfVLrlwKkptm/cph2UlGbJHaJaGJrk5pJT3o1pZFLwqKGi3xL
0dJVpmBILM3w63csulmRwCJMp6qgvz668CYtUVWcNZm06MdTZpwDKkLd9n5lyMKH4aBu+pDalpmy
l0S6KuDcIjSDRJsZsa0cfABBcTMtHxaoLOzGqij+rCZLu3yue1+l37IyeuPyA/sR6SO/DxgJxUlW
7dJsR20dYiyPCW7F3P3E2QnPTwOxeI7QEjqEvHYu8ttTv1xcEAgxfkZV4KIILMEzhy6xP4PVk28g
HE9aPSnP/eHyrlwFxhGSVb11Uw8+zBPx3QAn5pkDwcfvuGNyPI7p2uwoVg6LM2ROKeF5mG1bnlu0
qGUOI7vrbgU6MhQj2/VKlS0Mduyd9nwJAUMgd6wL3lMgfL9QE+bD2wz5I4bYWWd+x+Q5L/okPMbq
gQ5h4X5nP5SuXdkVjBcwH//UrjlMjOMzpKCpbs+SU40o4CMw2MXmFAM8x8RC9mpYVjsjzD7+n2U2
HT+6BqZ1OEvKL2Qx1i8G5HoNqstipqxB5FtBJdGa6SrGL4T+TvoYvwQCkSLO36EdN09j4Px/rbR2
1SUhnfb76K5CEUwQVVzqSXT5krR1f819DTiMDL4zzx2CqFeaCW/SJJzYRhtcVynoQZ7Q8iO8SvjW
Yg7FwscYpU6f9hGNoOo8tVtHjcwk8X3XgLx6bZxXlFK67YXOHjb/shxH+DEOCh1irUM1Qr9cYAmx
Hgp2fhISPH2UPwIuAKc53fYPw14FFzo43Ba2T/HmhaUOJ4Gal8G1O6XwnTA2q8Ae+tylkwBXp+x2
rCRupbNHhZ7QkbqU9FYYwqyiFzZGBsjq43kPKnORhF9kva1rMZLEjK5v8ZDL/ixQk8dwmusjo32j
v8wMLZIEzIDq7/muAmazwIErDjdgTjE7zkwrogbaaC8tBJla0w5GGrID2DsTPUVrbPmZDCZS/Uba
CrBeevqrpwUDqpmaAH1Of/uH1nDAAhMvmxG/vPZ2ovUDmyo0feK3Af68/t2P7m1FpW1qs15bELIQ
yjXGur+BHINlshmZMw8WFaF1TP00pw1Bh350agCS5p/AZXhEDEZeSb3u8y+MpHmVHsHf5Lql7aMX
PUp3kjnMp1PPthjXD3FLMKsWOOuJP2oIYQvgLla9P5RALQ2zjnsHcHhWLBMQU99VIJ2cVImITCQr
TWeKsXyhPW+KZ/midlMnKG4zv1yUHz6f82hm0ypM9EIIA848OXwkg9hFaYzI7fENBIq4yXEzR5DH
Nb3BuX1qnkdwXoMR2IX7qUGdnfH9EKmT4di9bFRY6wcIky/zWVpxL5Z9bVkCXnTAUGTlao/stNQr
6iCiT9p5uVe0PHv4X2Eic4LMWOQsMgSOcO4YksHBbw8CP3wUlJ4RIk9EqAJg7BLKdVLpLZmiuW7/
Mv7dlamo2ep3tEbWy7yvT8SLVa11itrqHEn6mSaHclKxipdyzvXXDbXWbeog2RQ4M/AFkueG6Fmg
NmdllXze4HeQzgEzd/0aGIidWz3SarEDnycWCteWzRD5ZlVN3EYMjDspGh/TSZN7iK5UbQzprQsC
ERKJkcGYY4uxjlCeiOl90mTS4uG5LkApLmQFyORj+qLqrV+JjsUXxHeE1vdjoe9GrpZexxmNWxol
rjg6LsUS5rZU66UhmCnlsshQwqKsQm3W7cFCY4q7BQq84vCwAD1r8Qz9Dtjqb0dBMvasahZ7ORWB
Z1P6DKdMIU1kV20kgqLgmTukBOB0Sc2g9fwIJDvtpz2Dg6gB8geu2o8YW9u5H1R2vT/dm1NGii61
BbuonbpU1scDvsO+9oB/2XX8K1V1qapLuoD78VCMUKnX0Bu2zcwQElLVr56xEOhPJxe/fQzfKc8k
W1+bAaDkS0RjcgqR4IwCWaj6KQ8TynyRxCgh7TJ+r2VHAJIX4X4HduaHj+fwRAPyIDmlneT+A45R
wEbSr6ajo1ZrV43eI6ltCpnZ4KkdkEmd9GPeM2coHi52h03jfJChvEfAZ7mThRppEUEL6ocTh833
itWVwRy1WArlRlBvvknoccUYGzN8VogO8s+OQLueCIsJ0Iv6+MOiKBh6cuXCpw05BS4MOmjKP86f
8idgndRJnnYDJOseQY+ekYeiyiyESq0wpOcid/h1s5ucfTQ3Px7SiFT72YSyJv6QzhyfRo6dq/y9
4FhAva9K4MiePSiWkN1SxCqBIdxlwZCM7Or78SqxZ/9ZnU45fyLDUVperJDf5chGLkpnO+DcWqYM
Ypl4MIuS+1AcoWacI0FYTW2ART/wDpM0lsLwjMg05JtDlku4+8dhMBO0rOY5+mAKvJiAh2k0IK5p
OfINt32KsxXq+JBJVCFg885P+OY96wf26xOSc1qDSNpN/xMbV5pi1VjLNz6qm0sGwOHJPEyxaIyv
EE9K+HeKGDjSLE4mwFAR+KdIsgZ3Rf/8StzYwmr3pDmHyrkkS1x89ExCUZLGg5i0fsOW4c5YUM0+
lGOZrOHv7PpWQ7owkRGTTeFX0mRV8uQWqDGuTVLyZ2ySwwTIzyVyzvQwVNfH42B/9mb9TmTVYs9u
ksbeVASnsAssd2jMyZEOjhiYk1JrK6zIGX+PpJSbaFXDJ7sg81HRCYddqQMqfagBxvbQ+cHYJNWY
6OkJEBdrngnwoP3OEgDwZz20e9NFytnqOtyD6Tke1kB1xvPQJ915Q2f38zRdlpl8Q7yZxqvezDgm
6lccGR7Hb9yoOxIYX7Thzt0JmVaortHXzuA92RbCOk+pwwx81U5U3rCrRb78j+BIcZCuymhw8NyN
wZw29XE+HBIbe0M06fOmgtdYK06f25FuUJiLzM8aoG3KJRRfr/nIPRfmdUYuFnhsr9hn4bhbSnsd
QvDwIPwePjS9w58O+VX341Z/nPRj5rAxQrXdZ0n3ZjNYUp3kl0FZCNuWTg3k/phtWUZAJ3XrRVzV
HjAaBrpBaMi9RtQA29Xfnd1NKlaff87bdjGvrdFUs15CAQWGw71ByycKvEBe3pFFngytgQs0Mzi5
K2rwzp7T5BwgW9zB/uE1mJs9bznTGIGkgP9lgXwfEgsm3lIWzPzBJTfjMufMWuweL9dOlmzjIlIA
ARHTCP6DRHi2P8HVSvEprB7Cw6Gmzgqk+H/aNqOF5G52hFU54/5DcN9gTRXZFb9bcwZrVSTHgY4W
7HFZPzyXXaI1iSUmm2p1+Fq7QcmX/7k5HKGGXUDlikpnTufLTTIPlpL0Qmrbnin7bRGSRDx7V+P/
QKFjNn9r+MNVXEGaTtOABnEK9nQGCCGWfg2N3FbGowyhAScZ4KOx+KlPsmpBu0+W9WKuLYGgtciD
voZuPV+9zhqOfQ73qzZog7d6B1SmhI6EE5vNCFLWj7LfA8LpPwPmubzNdnQth6K4RnMbr8QNgNMi
r8F9WdPM47zZHTo8h/e3jBkUnH5ozubpd896puEBRBM7CHaVEJbdQKqBG4TG101fT0ztSW5f4MC3
WeXYdJFKSZCAlJ5kpgKC3MgZbmV/2nJgepGEWcbVqdo9MJHVbc+Qkbgyg6HGm9Z4xfRdfPU1evoF
TGMFUGkH60XtftD0pWC3LtVDI0AmkCSY+9cLEq3+Dbt8wZ2b4Y4QfIQn5FKu3hy0miSqRqdim654
LX81JMOU+9cKMgDQQ5iBOdXpCvNBfRezkL8Dof8gYFBZhcDHCX+vwcFjJMIilQnoyIdA51ljSsR3
0lHvIhHQIdskjSQlJlrC790S9BpHTbNd/QU/NfVuEvA7Ck9S2ve4zmXgv9hVfhEg6ERaIsUB3YzK
cPglfIrQf1DWwMi+h/cXOf4kGL1Ot2bHrsw4E7rTaTVJUlIdIjrB/8T4jx/afzdW+W5IciLhMFxG
cS3Ty3sXANFtQdZwu3XFhY/rfKCx0JPDGdd3z+THcgqWSwEUdUDJIvQ8KcNmooicfxxMpyIOEhNY
UYecgksOGsb+VXMgTtSOlAe7Y0AHig1QghpljFstBZYK+T6H1bygnRKKD7UGtLIg0kdQd6+8ocwQ
DzifU08sc0Cyf9wqG5448eX67m/zvfVhMHIsgAwA5RjuEA6cLwTAs9KGFELXoUVTjG/OT/1nDE1M
uoebzxTL91yoh4s7rIZRtzwRtAcrP4h8POyHTzGmM7qCdHiD0SLwP2f1kyBAEijmlXqwCN/1HAqe
WXVIXgzswqKuaGx9LveEGrY5KSUJMRrx4/QqUGT1eRXUm5KNDL41T3aNcfRdhYIJkihe2r2CDQDn
k8M3wkwI6DIGiK5jYa5qp0IEMaEulY9HBJ7/3XhxDX7h6vVVKVG4d9MvYC5+LChg3/coisCDarzr
05rMssV4jqXW44WQONh+1qtDAxymS+5ejcdg6sUBqZ4YjSzhax6OROBIDiiCNK0PvRzFCrnsaBf1
LiSO1vZKrGH3IULAQVxVINolunwT09W6+QIKJAH4ph/arqhyeJdnsj6D5ZA/aq9WikDUVRaCJwX0
b3QONt7oWNk0B8hnLep3WobkpvobO6RDta+QYnM6TlyY92I7iE5uDeXpnzQ6asfqE5YUMYciea+Y
q+fM4I1CuP95ZtpmFwUNEXqOPRxAaoYzp9uIM7MikDTp0LPAgoOIUocMqGZ86MSs0fB1G7YHH+z6
GYDWYaKD7yIkSBKzJlTh/olpHWwmKV1KEfItI9R3TxRL0M9IE5lZ9efs7I59dZefOFSWWb2YWhJi
szyMQUOAukhd+MDYk18mtuQ50cVUM2Xh4Jz89FzmcH2Eio1tObZCn4MQxY+oZ4eoH/x5XSXlZUYd
4ZsL7Ou79cJs45YjtGRjVhUcL5PksX1mCPe4mWaN9Ozj1hp/b0eSk2/lJePAeOzjkZgh0uGK0J6g
Uv9b6cXkGD/ksOB2nIuGvl3CdrS/VJSAN+GmKaUHcrbDzrG2NKuCuFeRHuku9WDQgVglyLBfYqua
g5LKy9fIjX3WN8ZQXgSW9OfWEJd/y+LSkviesG7IWc548N0lhcflx3ATEbKCgzmB5Tog3ogGvet8
yCmIBjcpNjihtCdIEuDXbxLLwJ25mz44VFf1OZdR6zNuAMeSYSEguMpcp3BlFpEdFP3p6mvD2T8O
F+kK68kIfXX+IbZpwwHmiODCz/5OMWX1ihX6aQyED17iFs3flEUU/EGu9Qc7VQC6Va8e3AqrOVp/
pTlvOb4aCRRK2vz2j0oJtqTr5vwWaLfWiwr15rO3x5BuhnjI/62pn82KMcBQhUBNWbDPCZRnVidp
O5yohV20oXKL3uIbZOSepGiIv9z33eRqIJYGsTaTijv0DtdEikarvmUtDxJ4WX54CInsiIqNRyJw
iJwgmNH9MrsMIoyr6qsKlnp9/zlyEBFB4hLpAcGPV59uOhmsNIQo/Ah+kzkrY+poZ4fkHwdLLcWy
rR+YH8dVzvP1vNlxzk1P6OZo1jQwhhL5qZa5ZuLfOaNiA8Twp4zWbWFjIGgY6fQw1yrE1DZGPen8
BY8NKUMX0MkpCB5sGuYniHkWEagjBb4IupbRaSq1ObMVaCFe7DAswNjGQPjfjjzupsli2/kcpPxd
ECNT0wzjx1sMzW9gDrO96RHAMZze7oi4aR9ZJl7iEdjv6kJCunufUih4gdwJ7RKlWz4HuzbYC3Dn
ZtAFaRCRZ+HCmw/qoHEgN25x+kIOxfy5yWfs4o8tAjrywFxQ8LZHxhtJuKtJ5GSgYlHdqAB95uHk
KVb4PullVqqRqvT5wePgVlK8pOy8Awb39GGCfKfip/l1AS4Uh8lDfPywlfkUAlQl0o4T1dvam2v1
QweR2hm9a7Yh9OUQ2W+aPUpwPnwQWFsKEyYvh/BI7OGjkdsnJUpPPyP0Ds6a29bBLvZciYA72skd
TuqwSpkdKqA0ZMUZgfuNEyc73zUgO5EL2jIhEwmrST9khQJNr8YkE0O/QIlLKdQrvtqMZvvI0Omd
LXRAxSiWNMA3I5WAGyyNoS/EAtK87LzFhqhCQu1+bqXBx9wvnr3shj+gxjxok6ekOItV5WKdGMpt
+SfbDiBXBz8VRg2ywiBKoj4U8l/w2ErOpLQD1DN2mBjv0Spuf292XMDlyuJ5/wcbxUTg7ZO6a1sE
JDX/Gg/++tx7eC7bSfH/4sFEBdL2VUQad0xkv7tn9K29a5l8oNQ8ZvRL1+/JxiwmCJSB4OCBmjax
N7XEtTOi+QI+6B/DZa/Y95IaFMlgT3qnmgAGHaKoYksm9KfBviXnPcE4dEuuXjchVVUChuyAGf8t
x9JK3yVuKXvl5E6MvNHpSBTjli2D2rotWQ/1XsB72QzlGsl5rQNURMHCeZ5w6oz6jitJ8xMV4Jwp
PZeBHQQNso9AVTUdhoC8RFwVpsoTW8KelrfXerNi0xJmgoz2I8Ud01hiQYmcvzmCOiYHjQN5+Esk
b5dtpyS9MEx1bPjN1ERIXyIXeLgEehrv8fFMH3nS3oR4kOHrecwgblYuQlMCJfwVJ5Z9AZ7BbpZt
nPo1gVhrKyWy9Oi1kpInYX3KkaXCv2MOReWX5AyRobR2rSo4S4mtvnfR8Hzgu0SdflMpl5VBdwqC
8RybgzOqxqbbHEM41ying+Wch4TT4XyfEqCfIumK/+gcSmQMgtUE7i6NXzoDK/YcdaAUBIaS2XJQ
4KNLKXbkwCZwZraNaGCwXLIPxRmYeDJaIpzK1sOdZJULEjpnpJT5RXrT4mIJRHxctmmBZ5pKQS3Z
2xBtN0NBG2AG0lInOTTG41EjsZEtvBiq7nO9QV0q5ChZjclPhOQwCmQHv5BZjwcrp4bDrQdD+1hk
IL4Qyk+zRLB7v+P1dp6YaPhCNvBkByymoLovSBQldiu6mrfzfquqHCueDO8Kr9uEEM+aCYZ0Aw3/
JMuUaLwY/a88c0fLiEXbMZ9aA0mRdfCRqbP3gagDUj30HMCZBTMeuv5CaSZGJ67/H/D9L3iwf/9I
5wJB1vCeYtVxyOzKLK/MFccN+CNdOL+KsueAgsyEbC0jFQr/Rh6ez+Xkq29u+WIn5XK+yiy8lkHo
SKmniGc1de7MiOB5JhHjUgOHoiy8THnCqYG79B+U7aYMve7PvpyIGlWK4kkBePjxUGV1MxANlTHT
XvhwiJ5EQPndS9l6i081lT8jibelusHG+Ots3e7cJLWF1DRYuaC/gfWmtvlse4N4MKrcPfn00Hmt
vMTuRTC8HyBR/NhAGWKoHe76DSDua5xemtvcAj86UfWKJCScVfzS+hahMeEy/25VJjn7jWFVOWsZ
fJXpx21EsYPkbi9JN/HhOYENPHCf3hS1Iv9dF2NcBA648vUkLGSNl8Bwp8va0Vdbs0LARUtmYNRl
kZYQuI5/gP+F4vrh5WvG4MfTrJxjgRh7nEv8wgP+u8OD/zIl+w2zw3bof/AfApIWvdXVaq/Jf6m3
rd9VR7klmwwTwvaZeeI9d2zWccE5mZz9bdrVM/m4T2ryMntDDDP9a1wCIlYEAHx3xMjCJbFwlX9B
8sOmqfL/wUKDZZKEhi8fP1W59Qu9CAKUgH7iT5QVgqUwG5KxaIGMlzj7f2F38AjN0uYk4An0jour
/LXuCvmqoRHi7KmioUkBlc5eOrr63L8fA5qCZoTeggiVo8zXu8d+kBMaaolWuZq3SGJi8tC+AVXy
UWS2p17K+4aJE55gvxOv8C+BA7issz2eEG5lRGQ6rrXYG6nXG3HvjfBqfKKjtTVSB5K+JdVwg3rV
mJBEnE1e9gOpYiiYbEWvd8w9cl7Lyx8hhGhat/RYjZrCUrseO1FfFpOJh5rIEeflapWunm//Fjbh
LFl3cKKpb2XzrjimRquFkCi/PYUxwahwjYydnaTMxq2pmhzZZYWlge9PSsetwdk4gcvkJray+F8u
eGT4aLkzarD2nP0GHGzERdOT/apnlwBu9cFO+6AY515DVaMYAHq7eRe7fYa9D/RXr2vYSdRL7el2
yZUSAkNjz0JgNEoafRsjDpQJwQ0Darsx3DqIBOy3jNg4MnNCQHIjSsxnOXVismBkVpR2BKqqst8S
JApQ2zFIYU+pVZl2P1Xg8NaFCO8Rw12PJkMEgPoBb5qpkpzWiQAdaGoqIJBZ1YY899hOqiBJqxCQ
IaBL6ONEpla7299wEpxkviX8BGdk3H/L7R5jl6dQqB8kOpKl1D4lgsl8KiQwzhDmmfntNAoeaR4D
2IDar6Q8PUFUMUWfHEmxHSCLR3x15XWqXPs+7JdzqpGZ6oTU6j1R9ZGwq+0VhiuRWjWJt///Audx
Y9+/79mB43D9H5HX+oGnkgzVx4GRvfalYoL+2TyCDyK8tpas4mXykzaUq4beAhzd1PtCodpkACcg
tQn0aJiyfDHCYn8ThzNPZV+S5dFESFDNEMvUHMt3WABusARW81QSGvslRDInNwJB1IhudkZNSDOb
s8Q1sl4VV17/u2gZ+uDLPQ94aUBolQVfFP11nNHvmyS8MFm5wDV9dcFPb6W8KLXSbWkdlekvmoAE
GoEznWwzTsN6XCLkGw8U9oBUJUHikwdbBDg6RtXy88PKDxOqJD3b9g9ZbHzAl56A7CbPK9fAQDVx
6KaolIkVLU8qcOOR7AIg/diHSI0/1IqaqrmIF3yIuRdZcIyS73zThQszuruGbgBlqIARUju5bFqd
CJp0nKiRIWV2kVdAbEOcL8Puei6iDRskcDHucE+l8EjlVWKrlU82ljxUVraugMCNWGyEMTRf4lXs
c8zpDoq9KS2Q2HzZWBM3XeOWn/E6DzN6rtekcDzZLpHDtyozn/RdI11ndpMHlztwKv9m5jlhU6NG
ljo3PGCWSGIkN1MM4qctOhemEqif4wOBkGg7jFh/c0mvRZ+DgofGkcvAC6km1HSQ5Nra/7xETINW
DIZJTLvdnObe8ZFDOkiAf/gDvexnaozdlVas22B0wypfkVfJmR93zf2XQNwUHRm6C1xrRsc93XgG
wDIMb3CjJpD7xlnbcVC2pUGVltEAwj35Cf/FMbkl2Y8pH6OBJaEGjmqZ6ZCa+PbuPQs805mPhlgw
MHixEpS8zPlPxJyGr7Xey1zk6rRk9RHhEe6ayt2+AGI1YqazTqonB25xHw2qEW1f6c0Oh/0BBcqs
iFdM+Tnm8b62cczW63sYi4fQsWI1ocGLtr8QbhaDAMFszDFty9ObMiTJHKdSBM55xbd96Wr3Z9A5
t39N2H2rWQC0SGVWYcJC7j3w8MG2qGNMJplnxRtqPgp3uaPeKYfxsJGBUIhQ+28zbEWyO5xsx1ff
QRRcFB93pGBgURPhb1yEYYK6Rsi24TE75CbR3+Yj+pD9JB2DZVPDrISjjrEnjTfh9zIXB/anCE2i
0SdW9xps0mLBjXW6s7Gqlic9PXGjkNBfD8OxAm0BaVv+mYRrAhP66tV3pATcbsxhKYsTmmgrQYw0
TzjeIBgC9PjGwziVTUse+ePPDpzPLsuem3sQwmlv6rLnxvQ0e8DP3sX09bcfd6pdyEoGg3QE1hkj
B2Aw5vo/gf1p6ACcu7G7Q4lNbN/NMDsEL/sQdpVwnXWdFzPL1zvm31VmucAK5hn4rO2+KzyHJN7p
x8PJL1Fm8M5VXP4Z7kmGX1JkcyTgAjgo7REp7uHp1qapaczdZVdh7RODU5QUYadbpIwHAKtu3Smq
EJVxLLonPR3n0RS66S7Rh0XmOI7hN2CNhPqt8pBE+J5SJgIF8BXN04RsCio3oQ2+21rKjw5hPp6D
rBvo9xqREc7Kg4vbAzy9wAnrodUCIvr6w2uQMaZOsjppG4f+qaGBTlt76B1AMMuxvHx73NvFqA0Q
70nWX+wFoE75qOTr4MLF4/mhNv8GkqYKycxHydqAQUtJGih2UssLQeCp6tj9bKmXWlj7uPi5d/R5
IScUq8Out0BQlX2iCs4OmsQLJHbGILIIW2i9p62787nBHXO/7O00b0lvRUGCANbB/bIg4+8vko2A
qOpuUuGDgGdgLq9w9gffHel5wbtl7DHDVuzd8fATPhqM5I5oqKzpRP/iQ8R1pNt/iVr73p8t7k7y
XHLcYuBWD3d8GbHl+jXXCgFS9RpQsphflGYGVXq0pljoFmyLtQmQexYpwKKdzKoKNwG73DpsuC/f
WudrkRk1XkKB/TsHcKyjsVLAqfyJ02QO25g7E5Rp38QYLbEc3jKxpcL5JxmASYHHmPkz1yqusSp/
LvqB9f+UeraODTMFzXwRuF/W/W3Fdpwyg3GbYHRK61K3CUs4UwH+tzgVNzww6pe+kyBfeTYpcwLt
QPkMy/akJjY+2xOIBmwlRpIhbsBK39myMLilDvHgTuMK1afMSkC/O8Fu+zWjIW+KDSQouCyAuCOB
XpMhSXW7qSxU7gonXBAqjuTz7vVhKyM5FxlUCW61tvL1UF9JRW+/75Gxi2+dKolJ7NR6TbYScwFO
TQ+VsNZeNuCBPZLd5JwxaN2DG48VEPAqEmuLO5qDtSaNKZAhLmHpPBF2yVxXPSCRch3Cu3/dOT8K
YEv6SnxEk1MW8x/O5upv/pHyUkAOpwOyEXNIGuDue2cRDR/6SL8UKlhAAqlsTP0JuLgdBmuTSy0Z
vBLktrPKStK+T6AV70JBrLCPbzDY93DlUGrbtqcB3Ds5LOptRLdwvrxiNM/z/BUHn23kYJR4suAM
+4Vp7mgrMG/ud0gKhfAVsGyRzmikPOBsW91WsRX50hz8Y/lF+JeuiWqio1zSwUYxlDZRhqrWOpXE
xWDd7ztCqTnKvZmt6a30yKfUStoCv+A3S4slrNqcSClAwccQ6Bq84N9XagAFKpWaAmigA25tPHw5
TQqOBUTHnVd5Nqdk+DseeMfnllYsLVyMAusmIB2HWJVZ0m6oE8IAxux1lM+47bMWWUr9WFMVd5IO
1gRSqxZf63iJqDosYMCN2ofMjsRYa1z6KuQ7k6E5hyxc4HpwVEaqqy4ZWGwFPlrz5MAQS8Y1Ctk0
jAf92Hl9VbB0wRo14qRmmAxZakQ80yCOZ/77A/GCcTOtD1Ntqz9E8DYeYUJdzyfPHG+W64HU+o+J
0SfhV5/wKhRZNaGY45il+ppanixU1Zl+cg1UeN2jx5DpBSAJYLP1gcw1PeZ0i/AqpO+6UwMQO35S
6daitxfkTi0he3u2xSniec4eSom1zHvX8n8/oDJiwytvonwSzI+/yOFwFN/zXB2oOCqgPOzmu5e/
S8Or4qtenb5f8HVulrkyiwBKAg9BdJIqSVg2kAX2/uGlHRajEBjBbfzrV9tVLGl9o9/1lqjo4p1E
vTRvxI15aCf3JOOr1Q3vDHKQJEETyh5jeFtuVjUt6+3ADEU5Z0NQ4QLH/XcwwpSMH8kAu0/artW+
nyZL+MTjmMjNioqoLLBXfp+gOuZ+mp0YCfrIb9G88ffLvy7UlAP9p5BWksKa+twEgpDMqe58wVmj
C2IL5BFJ5+ScYK6FhxxfwsOK5zeTRn7Ljgua3q4k9WZbXyzN5ceiiKYxYKzj8PcA43kiVyHkK6qV
vAnRZV5u1TQKifsRUoEYbzqtWfEPVvYnOyfS36TtO9SB+krD1dkCKTbIB8+9HhQE+VaocCyvgBDN
FKtsRxkqED/xKNJYRz8JmjvDhpILQsoTD91Fb3bgzhdLi1SJVOwmmIkGqTtYRllv4N3rr5qyR1CH
PJ4ZebWwB7pzaCvXN7gQU/vozqWaETq74XcSWTbQEb+PVQYM+DF/r1WsY2M33e9uegviJNjrFl3+
qu6mm+vRbw8WWm7A+7auatf4M60leaWF3AVaoeXhDuDXa7i46VF/AFMWSWNEOPxA20LhWK7cCGC/
ZkmK4uDRqlLVh/aB8tWobdTXPlOiSTn6Jy265KAJc4tLJmn7+0YPOvFyFkwBjMpxenRlvxrHI+2r
dIWJaNzdQeHPHLIeHPwV+odWJRBp6OCBaQbLGBfdvTexK5t7HDyTRobzpprFQ23DOMv7ASzmFv/K
LMRiGiNl/gsU+p47LHdhGaFU8lIajiujlvVnZ5rmahVPEd7VE3L+NN8+/w3hX/IDaC5Ro8t/q+xz
GCK/GVx7JnKJR3fEt4dtTx4HbVFhUEcbtmYLWCXE434/xP4WM6C93kc6A3HGZb6vtVimP508R17E
UFzqG6vi3zM1PNCHd3dxO/W/w183cT5B9eg6S8RT1FqMBbfWoyAePGrDg99YaUWdf9NH753q7WD/
GQoEjc6wExkf81h/tkUnEUP36hVS226cQo7TclTZzEclbkjwTq5Bb6gfGHUvx9Xd/ugeBgMkR7jI
ZYtaHY/MSfHkyLlbroT5OcT0J8N7ripO50oEUL2TbYPHDaCP40r4J/gOq2GFIJJsVsAVplV2Bq3c
/g4MVqeBrcTMpfQr+awXzw0FLd3ioiF5m/ETOuMtkKWx7gJZL0rZ+AINuK649cto7ihVwo41IYYi
GgPjKrx4XJtfEyzY8mc6JvCA8JA/+XaJPe5kNkPA9zRCeqf9DEtvVCMXCIWqwrQt3c792xe1NYte
A3+xweD9aJUUIiYdK4+Ymqd9QtxWOxz0r6jpjNgrP4PEuliddVKht1oZCkAoxMkSclu5JHmD1el8
IzogeATHQN3502DK/3IlWEHzK+Xtr6Q1DvuEcLFixQDD0kaJMpJt4SBrhXF4cTPMIly+rs7F1Bp2
2qUDbWGHJbyg690/0MA9N1FSKf0+DdengOWjO0majc9ajcSqeTqIaD4kQ5ZcTVi/ywoVz2CaZtX/
pejCcHM3Z1PcgiWXhmLdt96Y5++0/XjocYbd40cQjnm2PIpJjIU84e8NOSNU6MB3tTj9tpLrJ0am
wB3VP5jCTpcMY1uf7LmhP9eeh389ufVDpdUW9GIFqea5pUE8XgL8OCB3PDcBeOjG/2Chbria3PXM
5Xs9poOCgqUcCjf9fNrYNKldCiGGcPczh81dD7Tw9szziE8PvWrFacHWCQNEl8Pmo97OAG30FNEC
gg5aScn1HLGj+KKDlBezD8jUA3VKyYNGD0M/quGfIFt4DeOo5HKzPXvDeRVF1SEvWcy+imdF8vwp
bWs9NXPBvicCiOIJCS0vYAgx3kVrJfNeKdqBWrEBQAkzcYmUENKiQgii3uUnpkk0DBjM9ipfSOsm
JiNOUYB0QdsTmaxo8ceedsCSJQ0QcoIvsqXWU/H6JNNEf0h2juTSqlkzWK4aJ3NnLhnN0DXCBMly
IS5I8kU/doqSiagSEcxLQ6T+qmJZg4TzUtn9NAkrSkg+ZKFCw5AQ8f+FmF7/mmgCHg548Gg1ilga
iehtX7VRbccwC1kssFLJGCjB0HLiPzvlpRn1TlSzuKxySG0d11s+M5N/5jPv0+5qLL1DPKJ7fw7C
RTazKzDYqwY1T2rFTN9NPLTq4mdVrMEUiK65/FhJVSbhVTGlsrhcIWN8n5kHPgKADz92bXMMuBgm
Kqkje7AKTGmJ65y3LMyKLfuRbFfP1fIyEELrug1WVHYut3RzRCGxLt+hgov3QupWQX8w8u7N1Okn
IKFr7ZxzCiQM5eKGvXLCg0CMhmFS0vu6i7ihfxPILwbB9i+iJ6L8AsFNFz/z+IUdwnStfcv/Bc5j
UguIKDMnBHYk7IRMe2PS/cRQpcIJgnOY4FHybF8l9PkSka/PKxiM4azGbQcIFGOOubKm9b5bgxSC
hElZkPnpIIaqopsuvh9pvh7AfdToYDUV0Dv8rD1jtf03gMu/E13gQ56H58K2Nvfzu/4GE50suWyI
2Y5VdZ+x89ohwO0FfKMmQyQb5Uu9qTEsB5UFuMRGH9zIgurkI3Iiqdy3/QyLZYRwb3G54gNyHeI9
MO1jGRqdGHdfoNJjDPACIhR8R73xrFaym4IcR0Feskt+bmElFbKHfu+pdRxnZlNaApodBJ1X9Uwl
6kBlvHU/ZtaUFWEj0n9DEyZEPreknewzaUGYG+ZjndmIX5xUd2QmkYibLM85MxAE6s/5I5vWhU/9
1ErPV7z1ho2XaoDeyqXmM6AV+KPf1ZW+WZaXLx4+RPQLpS0WQtZTTe/IJ333th7GU87NA6Xscjoq
Iz4ilorCXDi5Efm8P37/FOgo4X1roAJwBds6WxP9/bBtMowYyMT5YhNMFb/7xpK9hyepdA3+ftrj
lUwPyjBL1nS53mzJYOTZU52P81TH8ht7l01sZtmZbYZzzi8Y8/D+o7nTkS/NfycT5UXkPLlS8uES
UwsSeiI6ThAwXMZNJcDa1rdIeRHal+e1s6ci+dvmDDSU8ufOagSgRogqnNWcufwGyeVBYYgcfPUF
xZPyiQDFuUOBZMaO6A0TFRGSQnFf8yF3XTBvXYTQva8TjMoaES54DgRnJXQfaTrnJGw1aOfxpJC+
/8WV2pXSepKBD6w+vLFXa7/POkwd5jvhzxyvmuzOTG2T02PL4FPtBqw6J7ITFIUeFIEpce1x5vvG
vZbkwh1xcvjgAciymNerCAzUmkCt4qlPRvwJB5m5RxeFMEezTriKDZ++bVeGB1Say1XXbpSzmB8e
Rd2Y+h4ZwXw4B0xiGhV4Qr+5NroCLWZ8pt6W3ehkbhEYwUdT8+TN9FgaeAOVV8b+btBSJ2w/XFF7
+G61OzTo6KX+NV9/UogE0t/co/AMCz8LxzZsFnn+mOOxRez+0ehTukCqeSlBpvQmjh1vOfc9OGl8
fSofZfHoFfYVeeI9Ryp8qIKgKy+P4GmvHhBAfBdOgNgHh6oisp9oNIjNzzzeCHLq/eg9OKNceeHy
sww4dsvdFo5M5pxwnZfZa3wCTLh20ZZluKmsICtHbpE9IVrX5zsYXfKJ9wIBRvc0U6iKu0Qfp1hi
O6EMjf58bb5nNxuPLy7h1VSN+UkkTUxfzB5eLhB1679Kwexew7eTtI52EXYPNpIghWIomQ2gQL6D
GHDcr/juiDiPfO9M1Zd/3bF7gFFjFtQ3HG52znBdTOhzeRFl8ETmAyNOkmEbFFIeKqG164poeOp+
VQzleAtjdZdd9UQoKGADKo2shucxIPyXJlKvv2Zm3ovrYR5SpxFoIrFXb83ZLzQ/+69myTsAqNUT
giK69nIpNLVX7suK1VpwjgmQdzgBXw9wJ+pLcGTbd/suHIsYMUOSLDF0Gf/arxVnSvy/voXvnjVB
0Z4Yb1QLHh5jWHo+Qd3EZRI2kV0gUkTVSyx1wJ6G43UBonvkV860LsDYDmfn0RArhX5RsA7tZ0Nw
nSObK98FWggLfyrTjSk6kWJ8zA00I9t5v48lJIpTh2tkEIRYdKFO0C8oTH+TxN3IcfQPbxHY9jwK
6NSxY9J+pWwEK6NNgpcJHYxfQthu2UMH7sS1B+xwnI9RRyo2MgpEySVPXeDT+yDz437dALW2H6Ac
OFluDLuLbHAQX46g0U34dBBgszg+kZ6qFvN0PlnZazqhVpRnnkUijXJLgJb5MG3t/hcTtNXPGqkV
kaYiZyaEYsCXdYFBxbT/VZkak93tXEDOcqRwkoY1WJzbM9NUa+BGztpXnk/ulPDjoTwfKH9HCDxu
wFpBHPDpFktorootv9CAoxEHJPM/XWmGbYkhgJ4bsojYwBG700I+QjH7WKU5lsidEs69XKrZTZpi
RIed0suMl8sbYZreajlJU0NtXZ7Vwl7e0qKzG5Y/jS2Fqkqr2x6tbPiQpmI49YMkx4qkc3AT1yYT
XzlFkaXeNXclO6l9ud8dsIfsWUoeJ8fyRsY3v+N3A+OZ0cMRPQTq+oK52ROiVE9oqLEbnMULIZlG
BQGLM9r8XcS4FxEu+xAhkqHf3UWGHD2Z9cjN+pQlRaEu50Z6W8wwpwHA6NXkMuq9cR/i0DpwSwKF
1Vn//rgfmKAWqQXH9nCGxUiVTtBcRA80tc4JwBT38ELIZJwNrCoLyDqGQkD3TgpT4zqIMxQTuO2L
+rgSCJ1uGY3xGXvuMHpfORySd8PcDAVDun5a1QpHwdLuPGEdxA4VjI0wTNW5DwXTUjxoUZdpYynL
SJ8JgD22SQFBv1iGtU5SilvWAthN04MGOmjrjfTLPyba+7UoIWm2V/PbQcmpK+qFNF6GUo/0Tvye
Qh8sFnjfajMRZ/pv7VHucdIErlcvsHnt9QrPwHeVms6fNZNYqFaAg/nWQXCMUlzAr8d9A1jz/tAI
OcaFo9V7Fh6piEYJoktIjPQV4eQcDtYTKrQJ0uGFZuX6Eg9M6yBzaeqk0t3YCRwMVvuTFjS/ud9N
GhuKj+1GEetPtRh58Zd+KHrQnaL87fd5y7jLq2/bqiaX5gCbNShxjcXljjElpTC/xpAmKT5ZgwSd
EvxXC3u5yuWPgs/E08ILypQEEtQfYbVCKFaVR7/Nb3zjT8BU4WfhaeE5A89JdDlKvmDOLlBuXPZ2
bUPtIlLnuKW3E4oU77//Tzt5D279T5R09+aZ5aduDz8HbpqOXmc7FhjIjbDAtQd408qqljWey1ya
fiAKZK59DL/p6Qq0u/FlqW1RTY/i9vWBP1ybEfoLG21bLI4XAnJ2jU4RWrjud1SkWxDV8x9/eXDO
0wq/aXBgSfJcdlq0jGJpKrOMWAcEBSOJ3d3CcGevAqiy/bn+2UaF32kGPxS4H8yodNS1mZcHoCR1
vI587ixITHJrqHLTDsopHegzu6Yx6jGtc44W34iyhw9s4jB5H8HgklXD+EjKG77pBaUg5Tm7aZZD
G8iLt631dROC3/GuLAxxf7ZcqhfYqXK2lQBDjTn0N9pwIpg1Ftg+AX3W+X+HajXBljm8f+XIm9JI
cp6bGI/Fp1+b0yo2KBh7cdL5Fh9pxFDjUV6bjYAi8Vq5hLTm6AxesVTapIky2YVsWIo2dLiuuTb9
pObOKnLsUG3vruCRwb1qJWuyJ/o9Sl0l2bbat3H88Hi5bAKTpfXK+74MYokohL+LtMZYp5gPIxUJ
i6/6bJ6lKxFn+6PLDxQxhGtjmAwKpl4AmhWYV5xbBaU4mkW31gTvjMOhrSyZYSvoa4fU1itOu6bX
/oXu7y40fcFjN8mnjTdLqsMVrc9xy3Iy1dnsczNPJL5Ya+5ktM9xQbp077tQkrRTohxxgiUKTOXF
S2dNSw61gtX1mYduh1495JqTkrE9PIGo4A+rYvrxC0kk55odxT3g44a7dPrD++2vfgq18yMb2sBS
895Up9qXqLtPhWe4ixQD/NOyLuMGRsxgI/WL0a/dMICjxmHODDrFTrrvBl3ghZt+g4WJbPgz8F/q
oNk1TmCfY6wy3R3JUye53g+2J5ma+jErWSLTCFVFhO0xLIc0y270AY6jj3zplAhrzSUUR+/BrrdB
T11JvHaxis7qMGm5GhKZhOsLKMHUfEmoYFz5zpTcG60vW0xq3AzTurTZMjIZdgSxebvvVkZwbGXF
N6E6KM/A0rShfp1u18C1hjgP1GXfvjIJMEiZ71ke/1iwTAarPKHD+qvsabJk4zEEIOKFeP7YR8jG
bhvkG+Glv1QjUsnE5xJGQRGZN9OmMmA+3fQN4MscqO3dAVMxzCwuvPwC0VATGbVSt14MNtahaUJ8
SGFwb5rIVcUfKIwkeROw1yVOiGFx4uYGz2nyQKvEMb08cMD/FShjN7osTnNjiVX4pGViQbgfSOBg
WR6LSgHIIwaCgXR1dmYvz8dbdxrYTXxpmfsCzJXkx8lFd6Ji3EIGHzFUNtvCzdJS7yABpc+g6748
25Gr2NTkFUIvPssM832yyffx3e4+gUHvAiF0Bf97AuAX8sSs4dCZvD6pe7TAatcA+yWdZxKcqTpr
eH2MZ/uaDergJu6vMF7+hFFZaGJhGu4OLwuzLjhpCtwXuR442+jPiFwvPw4VLU2frN7SVdK3m1ml
EdfHS3NcrbVfLIqdPOOtWy9V2JTnDh6KKCZqMUEuqL8rIR0UrXGryLSSyVni9fTcPRFHjwUzt2Mv
T/9YHKvDOaNF31iPtF3z3nHqq9SGfNBrvf16psSCtWs1BXLSs1xkiuKxwMEV86U21XsnnPN57c6h
UTNNjvI2xJbrsiPicVnlghXFMH8OGR81NNQMD6gNFdSDvxmeBg5tkSAH3aeUmEIDE/BGOScMlj2U
ydlzT8hnfrlTvG+E4nDn+0oQjjWdHvuKoB9e4FH5Dc01Xtu54/CIRbY2u408IfN+MLG2/c/SyqIs
ujJH9GjFyee7ZLWR3CniNGbS38i5aNDh0CPAqssiR6qi9REWcmz5ob/2Hs2003Yb0snbrodmOsqg
1MZtp1yN4Kb5WM8DLEYPY4BR1US602tb/8KzIhCe8ZEpCzZl1Nm2f82pqzpyx8xhno8cOXSftkHA
pUWONTbvv7UUI2Vgfggn809fHjLlRg9KHH32RZgec2UMXOBJt8+ZZik7WaSJZrQQN+/bUzIY0BhR
mtT6EB0Wtf31tuS1HQ8cTTy7QzaCRH6TJDREClUdtBy/Lia3jKUxjgx1nRONo478mOtiA/2JD2nk
c8gwSWWPatN6/cLORqxbWM6VsK8Vr9+nkOUJ9lMNkxTeiiEJ3gYvlgEfa26fLB+aGuaAxRUoULqK
9OVWCF/p3dl2hlEzdfaGiygCDh9DHG2N6QSXZ0jbPgM58T5hiCpmlGHd/ndncMMq/ecf9UIJAqP+
UPJXPyZws5OKmIQVmPpGda825pTMPYJDZUcUpuA34bAX1oVhIpUGISj+y43h4Hcoh4hoGN8vWpTz
sRgYzCQrxfFTv3PlaoVGCbl+lgpd/MQy40Pk+FWtnjKUBVYreTXzd7fVvyqT/kgFdUNFpbMD7k4U
nNeNMm36dJ13CRUwSWLyAJhBKaIMJw8M0Zn8xicLYJY/5+UR007k1wenKL47MTXadFuEVl5v0FOd
TiiTiSxFGxBjkNztuZJdKSwvqASdQPBYKcskDpR1AtW7MXmukfLrsVZaL7qitS0mpbD286HPSATo
UFhXc+YoNG0tDMArlvWKCS3naC78zuzm1C0TF+H7p4tGPwJM+3rokGbG1EtsI6W+6lGnDVMTtZAv
bTAZOvc6oe+9soy+KrCB+ea6OM+iVUMANzPkud+OB46cXv7kcDQTnzBh44s2gTTrOhX2D+u04MLP
VvkbucBGI0R4MtTvy7buzEiq5a1LTpXjBkcuK0lEEJTuqhtCogp2Pz2SZYD1O+y078WcH1G0137u
xZyipfmo3SIJ2R/elcn6OJIye8KtkLmg/0cDbvZ9wQ3U752zNXW2fkKJfXAAhB6zLzahcG6Dgt1v
lScXRmPtgbHkcOnn7EVU42JTf9umu8dGfEK2lb7pRh4zT85yDxkFsmlYwsxeCDy84Sq4hTRWh0KM
XL6Rc8t8z/7TrfUq+UTemoC/nPBj1vwGRPZOgaim2SW+u8943yTXbYLQUI09fgEJIXdBkFUq2kku
trcvQSX42TdkV7vqbEw8hhrOGhCzUJ3ArvRhBGjhE5Kpk+H80ohy0kGLCWCfw4y806gt4Tj0/f2k
B7vlqa/j6O4PrDxb++TWqoCGrObkB1WntvxaSc/WYQi2jBIIOahoJo6k51iSCB5kiaHHnom2rmWm
u2GSSGNm7n/5fZRJJS5OW5HEUgpMm3ncERecNL9ired+Vz5/w9MbpqNWi82r6VhMIya3X/1/uQ2p
8BkUFPpJxNVHZHAK4f8dg5vyHP1xmYGNIQcm9BfLObhKMxHZgrQWigcxwQJjNTwe4+OtBDfi6u4Y
1WSdOzET/k2ZzBqodp8EgOLMQtx6VgtsSNcnW6YYyxieYt8vqly8Xl742ixU5TTYjP5Pbfxw5Kt3
6SFMmoYi/KU+j2KwBQAh6Ax+ajFiwhjunI3Ps5drTEswVlgVsvq3IwYoUw/7dfSJFlvDEnJGjY25
GNs1DZsRdUDr3mdbEu3VwJg/oF8rZVJPOEiqTbVirhyA+Mts4TuGn2Tx2oX+OxDYCh3eosHUApkC
/DzhelWdgAXpzhHzhZRM/XYbmWXDdBYLxD53q01bnHOAaIhmjogyTc4sOtEFHjXaPPQcNaLkP+zD
1g4e2D61mChSHZgrT8oeWuCXlBb1iZEc/8geHvlVk2X5AtvktCCa5Y+/LBmcoSGe5YD88tnRUL4L
HHGTDsYyfWixjBmvo3EJzbSN35wbOFO5U0pVvjv0E5JAwjoL/o3q7dhnbjmTBKkJB7jpn31Tpb7+
eOnCS7H0wY3RwV6ZE8dW3CsaSQ2brYuzqouRVkATJ4HJIJnrjyDKUenv6umB0W7UvW+/9wSxXYUx
5ExLPfTQ8YncHwMtXPflLaCworgaFrNFVLdkTa1P7FlTXI1Z67O8BoGEWi224gdw/kucJe0OEocL
5ItF4jgvkFhlRSuVDPOgxw7WCdej0M46XtYhEch+C4KPOYbSCmYOFlOHsT8Bc2fQLVAAG8u1buIm
f4lDsrEnQGLYxKN5Ae4+QUEZNwtCAjxQ1ZFBsruvx4JHPuXiKm6+OuhPizmUeWagmKPM9oQ2r4B1
pPq8G4CosAa8hUbt90V1scd2LRvsx5LZlSQqCUul1df4l9+31m3qoRWaX9ykEWHt+tCFw+oly72L
r3PuwZApf/+K2zYJo1wJGtd6qKmEbYcqYJkmtKnB3Pc54OKUm19EPj0bsx6L0BV82ZWkhFPO4ATD
4jx9bA6J5Y+q8RMcGSeE0YOvzOOvrZJ7qRElwlJa3oVJAfOROgY4ddQtQEh4W2xZIiXFc5SdBTOD
/OXQ/HobYxKcaoLtE39yrHh+P9LvTTtaS1Ta0yPo9u8KccpO1hfw5KJoq7Bmzt7NvZBs6vMJpUp5
M3SXlj6H7IfIolnzxsHFTxz85lhPkhNuV8MrVuFEatCL24G9DMBRJGRtw5cgycHzfXQ35FzrPwh5
0dUIpAWFelEK1JqwI3Rqbl/rJxCaB5+YzhujlwEyIdUiO71kOLfqlK5AJw/FmsF2e3YdPFXvs87k
4gcGIH10bQP9ZMI/En8MUzHD1OfL2C0otppH8XtBelcJ1THuzPxq2prmLIoW8pPmyt+uvymSdq80
8/caV0faxiibSR8FQ7gcSN306hOIDsPBJ5yyOb6cii1Na2tsZFnWbk8SMNiqSOfgKD5XrUC+n95k
jVAGmnjbRFRjvTHbQrRy7wbOVvick41cJxDUHxZY+uiaRUpGpT1L0Be162vArd+2NUpa50SaEjn5
0X5C03QfLA3WIB8QwO0AFc0dZ8IyTs0xWULRnk7rcxoKbgO1FOm8lIGPLU4Qsf1uPV7jMGYXivUW
es6qhT1esFuQB/HeZWdkcyIcfJCRHcP/O0pRhDavKVWqwEfMZ8E4sZFN9it1MfYao+OQ3j+BayEP
GrXZhaLTHozv187ZQU3jfLFjCiv6hXXbjOnBHcTE0l36c1MeNxV3RqJEumvy382znBYIgFB0zH1e
CcG1aYYDCaW1umqy9cNbAJBUgYFadNoaUezyn6W3TVkDj6FY7VGdaFC5v94j6TDi3EJ7FgAcGzW0
AMzz5fOv0gnDy6+lbUX0SC0eE7kAtRK55pHaklgsqVEYWkFKYRlEnn3FOcNUWuMhXWjqZLTJNTKU
D073EO7fyqYIvp2Pdt79fg/PLWUGWwLv6H7jJ1opFHLk8lgDB0Tz+E3hbnAhQRE21O+Onz9rsfht
Qh4w4N+E6xC+5p5wFGUbFKkeK8byRtT9Rf++UGSzSf4iSwZpkz505Q12yLo1ZI44GTysRo2bH2Z5
RMZGopGgxLDGov4vUfJFcXTjC1Mcbu6YniaOI6nInA223z5t3Zjyu0j+hbv4uoU2O16Bl30LhQDo
gyDCqU9uQYSzP3GnWCAhLVCL/yB/peChnYXexX/teO32oEvZHqDVYrMp7jkWZ565Fk3wGDXj/FJ+
LkHvvsl82alrtyyM4rNcYww93ZxzIi5sJAKGhBA34ePS5B5jdSGEFmfZkHBqD5w1yyNDnTIlYDDl
eBoUVQN+PWyQ74Vk51a+HrW6Hq3Ha0q0octtaYJeQKTcDlWGmurP6uDef7FfBZBGDM8T9utGMRGX
vg657HSY+oaHXvnNOLc5qa6/FgXv82hdqdN24nrCsnMeA7FHHhPEI15VVUH+SlaqgA+YgPTxl5Re
nf9RnMXImGlwR2GkTmbbVODf77NTz6eu8I53oDyxJQKLprtveVSqg6DVoyvqW4bmG+bm76vV+XUA
HOdMe9drQoqMH4nVTTv3T67NErGZZ7KoQmMAXAvTVeOxYEgkrAHiMEJyMVJ0Qj72o9nJsiuUjW75
be6GFifkg2isxm9QybJRd644BMK7I17zbVcClhvhpQQ/svpIAlZugB1Lx5LWf43vRyY+WLS+9dMG
/tfSAjmPEJAnilKhXual6HalhDcp1+H/G1m6ztFJwn9HQqjm+ScgSG3zBM3AAgFpZ2+h1SeZ1RsI
euhswXFdP9zE8TPDcBuMBVkPMzaSS307Ad0cdjq80v9Cy59eSGVDosii20q7URsr1Aq5VeKjXywK
mJ2ILhNwhlvcOlBmJlKMFqwfyTkuiWnd6lcRHwSb9TXVFCuBQqm0cBHLYo8PpJjqSphaJwqcjvs9
gvRTzzeYrDFWD4jiKtmonchetHlIcNblrfV0s4QkK282TeC85/zpAKmL2cx2P1Gq5bV3xqHjfrjM
J2qbIlaFbRYdfNbZIiJVV9A5vMOCGW3nKlc+hN0r2uYEnghjkhjNXN/qmvcUNLsVkxRAGW8ux7EO
vPzupKS+OypF0Yp8KflbeY/Q4VTljUvMVLMb4dE4VRiJwaz9Om316ZRTviVedZVijpMCDsVyfiBt
aW+zD3jT1TKBybHwkNOBb8BoxUec1nAiTH5NY/Ay02SvDAGP9+irO341qNhjGC6asTQD8Dh3khs6
re5pQrPLv58+Jg6mSdsoELnnLVJD2uOQFzSQy/dLswUaLaeTR8Q26lU3yo4osjOvTmY/gGUChOvZ
+5sOaYzQkbDQhM3odxrw7ernPSJS56fZ5zeS0/7qpmsATFnDPDHCjhvNHbjOGfijhSCqnuwFpu2k
dIzEfFaHkoqW0m+q1ByKtN9Af/tI0OT+YulvRm82vbDXztOyijwdZUH+NIzN0GHu/nZ0Q1zRYiQY
jVccfWNAKlur7W9/TaiQuTTnGQ7Bt0ojZ5ncSGSS+Rou1hPT7jM1F76KqGSEmMd1vkWr3rUQOb9D
WMs5lec9CFTqaV49U9Ovg43Daa+4O9jVYfCRR9LGvUcIwlHdsCMjBKTWQa+IOaFnVPVOKrkXDo4R
5LAOgqtPMz5XjhR3vrN7qDnSzFysmzfObdtPqvJqCOyscMquMlJn9xdONeHDLpbGmrrF93EPspCe
z/hadLptakLC8PBibdiZ9v8qahYtnUBjmMrRVGUtR4h7qxXQ63T/Sc0MlYNnfBpBsABjPPjNrLKT
oHz7N5BjaAp9+7Yg2nmiHCDIpDsyA5v4prY1G1uw7Ffwl+q0JZpGXd/HiAWUi254ArO0ZdThxL42
05BhFnZq9WC8mZF4k6FPTDYN/NEpNF67WfMLN3v3psviBcbJZh008zlDO9ti8Qk9UUoyDUKsX0Zf
UXZm6H4e1zOZsx9nVtoprgtr7zm9/6Nhg8eQLd4guprMnforLVTiLESf0+tf52HAn+y7nZRVaPxB
rkmpcQoWYjChQAjbVeTdUVbac6lmY1rGykJqg5vy4R8tBG9g66vAI6oFPrufwb2IAEY/fWFc7syH
awQQmnT1H4dh/ebQd/p1/TZtDSM/7kAxWySWCyhtpewTJEEsjRR4itVMUNpMNCmtysW45PkeOOOo
2dHU++tbsS8t8jA1pAaQneOAdZGHUqB2i8A60zHfPWkbk8MzgaW4Fbljwa2VJ5Y4BbQ5b88JFEO8
WyHq8EUrWc5CtsGhbpJiJq49pNf+MpywncymoKNuMEM5tIJ8z0Q/lm5JgfcwhZnO5btT9/4fTLRJ
X5jJGDmime35pXeKrR1q317/cuTkxYMhCziWDI5u7KXuzL8Dcmn5hsQZwxMPQAi0GbbcoDeHXy4y
RijY4l+O9xeWIAs53DgIjQ7+p/vh3D0GcytdEDZH+C1MECdOdCDrSC4Y4Iy0xzierBkR29SO04jn
axzXFS291ufMxsn0UzXtLNjp3vpOjAqlY8sdd9fFisrtA8R7fyXAKdV2R42cog/Fxm9+rDgTrLak
vJhtbYTAu9PXREBo/PntFyxEMDxBUXHtboVvc9D5pq9NsgW+ZzjX8N+8s/r/A3fI9uw3yYsbuQ7M
QKmJqFDY1lSwJhRDBgsMdJcRQvi/VbDUmFGY+zjzr1MLw+rjkTLNPtneTkqSqrtjxdbsSO+jhEFb
GwWCjB0sfVOVESWsg8XPYfhfQQM526/+Qm1IOveBNbZRg227R2SodybXOmmRZRqptIUH+xwrHhxW
8dG//B5zjZq5L8E/eME7RacU39IR6BUHM24WBEfSnsJqe+JU19qCbGtAFveD6Z5gyTdEjl+ED5d+
OEkv1/LCdtzz1ItC00XCUgBErO73lTSr5kRjnzrL8panaXhh1yL7V0z15SuMqjEjwiJFhGscSIYi
8XkL7TrRmoNBB63WnhllUBOOKnB4sZjImbE4FEEKAoJfAcM7BHH1Ge4AD1wAihdZweBJzAvBH1cH
RHHxrDMdJCdQlhlOuAEfb6iE2PYo7lBGVePjThHX7Uj4Yv3v1tQABEpTijCuBajUcf49EQZ9Arz7
2XsBN7yHsKiq0fIOWlfXBjAArkYaa3VKKNa0mV2NM/y3yskwRQRp5sQgNPQWVNdla1QuFPGnZcIy
KeP1Zr/vbgn0OV+l8in0MB3fbxc6W/77iQ5nS6B458JnrGq3A+RK5Y9zQC2v2/86vwBuCcmq+AQT
SJqyyaAuXOEmwvXDYuD2Tl6IxQQqcaPAvFfkUneUgmlBbiya57MtKMP5v0iREgEGrTFqiBI3zf2s
qmfDcmsnvsH/cZGmik9dGS//qPUC5nNX/4LfklvEqZDO+XG9nwunq1jh+F4iBXZfdPVebj+1lRD1
gv6ZzssxkPT1Cq+rsUVLzPnngGN4ciQWyQPBgQ7ElDaV1jc2aHgofmhORaqFDCKdMHgX+QcafPKU
lwCUWL8bgVQs+wNOJBtagNTH1GEM+PMXuKzQ7L2DgEdwWfzL5faAbYnamhvAzAltpFR1JEaxVXXO
Llhl/H5XDJNkA3mWea0Pu9j98ysLdVlwdSXiXv9Uivf+2P878e0afva9zOWDXdnVZ/uXEm0uPvYz
q2ulHT0lSipkn6TkrjXbAnadt3F0+ynlTkmRI1XrlvmqLqNE8AEDle4HKWebbETVRsEuy8m+6Sr/
yG/WeMQ5QAKirHXhsKDr46m9IQV01GbkzEUgBAiQCpXnD3AmZ6H1LZgdo8U7wETqNruMQqWDwDfg
BHCl1bwM9PQ5o14TDsqZdLmLNadNa7jy+2cMbxg3qdhG0qRumM20jYTS5c5nvVTN9sLctnbW8S2T
vI8IGjuS74LJjRpyD06jST2H8hnASvgmYw3E+9aBnvKymtUyLYvV1+7C4UJPv+MjcIz9u9LeWUX9
yPimBcGNosMVgVerSsLU/PCkPfTU1w21Sedf/RLBjIjVuBR9Hij0A2b6LWjHi6bqbKB19Rymt6h+
bbuPDJR9b9IITSEw2JkCcgLr86F/ZZzS32L1tx0RXmNwsqY/5qrq+X7L9tg0sdEiIAy3pDcUH8IB
sJViiUeli/BMF0jd8rOITfI7hRDcv4tpErBSdqKBOOv94C09MOy8qIpwv80RS8xFAz3a+ezCsG55
ej5zz1dfHFDfxzqdWOHV8dpvfm0VrMl0LYZtXdoy57sI32dvwhRq90MJTP5peGkO6LhW0wjhRo2a
oyFa6l98m4SHGWHZ8msi/ICgZ9w17dGSPBTNw7kRq0KOtVMC1/vfs9kp3rGFYr3McOX2+dZ8U/KK
TntgQhf+nhUbwAGAJsB/4yUddi795eZBV+GDqiTjgluEURG0/CcitvDwk3TiveDPsVkJHgfLzuKD
8t/OLLyz6Pw+yqr+4Imd9Ih0qHLTunJvnpURnOYO+H3WN88cmZg7XoDkA4S5sqWbDjhl8/7c66PE
iHKPHUEEHPyEG16sc9XOVvFUagJ+usm5OHe5Vvd9NqnrY1zECIJahhBiEK22yMeGFWyQYZt7qvRY
MpgZ6SrqN1oCx/jCXmJt0t3XO+qpKAXG0MhnV12KyuBC0bgbt2YC/qjZkzutynlM4ZU0qFYKb/XJ
PhiE/NDZt+EUhZ23rP0PCAt3FsqEZ+ZNmYzV5yw5XPtH176v66aGJN2hB6aLEm1sBa/X/rbdOaQE
ICCXB8/7H0n15pxx8k8wU1KaNQ+pEWtlOyx+dRhYs5pPkZTM7wvvzZNlqExgXDB8fpCI9pzKzMFc
dhyVsMKPipb8d4hegowndtzd6oigDZr75dzMJ7bmT/OUAyHP4+4WE4EKNYHkOgU+FEH3ES30X70S
+t9m6GXJ8Nwl8BkiR3YmqdY39sSV0YtvVyUvUmN3S5ZRyNILvb84fcgjv521St0XVtdKOJe2hH5W
E96t0tQag5befZzepGvfA5muH6u8geSblEg8rmymaBedP5p3mxRtUt1vDgBmSXFM/Ulw4KwsImp/
inwmD28Zh1u0QFH9BdJGJTwKt3x3Xivfg4UKnJMz7UAsu9pe7fJh5gQR81a2RkGQNcqFTJP9yvjW
8QnkL+DExqOZQvW6Q5oHwqICrOqQgcYr5xL+VVR+MOKAgvstp4LddQIW2ose2ap5LsrUImCOk1Oq
Vh7VZmosIiYlSDen6lwNzLJa+ZuZZsU1eIbDkVPCqeu5W5xXvZAGehzUSC9Kio5pfzLTe+AJfpUp
tObEc//f6JQe2KzmwBo+uUjKTDu1lUq+vdSQaPvYiY8z7zfDx0WHElJl3el08VNnlj6UaX1SuLZ6
N6JeJMmKN0Y13UOgDKN8AkXPpfmiTpc7VUzdD2EzU5Rf2l19h35d9tqk15XlsPwQK3wzHGn3lw7e
kMxmxenLy55RQlkH4ki5YQtgmt/NNHlmnhImoC9Qy6gvtMnWPDf22cVIOR2KNeoWq6zktW4MiKhY
czYyaAKf5JxTaDqLz0PiiKOUaMw9+Ds013JltmCoWaVEY3IKyftZvT8VxhIIYRRED/IqAwY85m5o
Ud6p8Wssjg8Aqn6QN/onSbZQStiuISBqAwMbzsPx5f07EayGpTu2L/TUDDWp5ypU82is1CM5IUzr
GAhTn+8uuCgMALkt+SxRO4kFvP3uP8rEFaETpJI+fWqewPwUfyQKxtRFu2tRIsPQNoy7Z82VAOOn
FpmAoQwx6FHNzcxb3kIIHfZokGAY57Pd+Whe30VZxrP2l/kHDG9TuG4ez2WaNfRpZUE45t7P0vq6
20feiqqkrhROAoraKJrWY2XPgkQLxoSxVK/fIClwXh5tdPIXtO6kTB7OmRIFcRDQSi6TzRs2u+q+
BxDFB9TWvJaXPcmDsGRZw1JydDSiE0zEsqTW5B6ZyOAy5ujb76nkmyyi58yDfGPpS3Y0Mwtsz6ib
0f+0ENgaOlY9WPk5kQ6SJ8UksNXgJQ82TqBCwY975HjfHvtg6vLh6n9v2u/h568oITl/ex5Okkf0
3qgyQeOXeMZJYABUEZEcM4MvinHzE4V3CukL8PY4QYlVvwxvM1//pzzU8t1C3gRZf7sEZoKp91Vl
FhQivAs9TsQaeqMvkCenHU+SCkVMkWXUdXrLx6cjw+fiUlDbxrQJZFD8/xqT49D5ZWR8AWljMhKB
pW519ndd51sRYMOJqHKYyclaJgWG6PexUbj+5Gfdua8ZakHapGF8Ujei7coqSHYlN3oZTYkdeaT5
ggop7OrO8vjo+DY0pn3Ti5f/mGTtt3wu4CI4OA3gdLqB1p3W634L+BTW7EFWg25q8JDtVCiJb0TR
uNp8uunY3w+mmnxF/BHcmCN0rG7pd5/mGQoxCtkK1CExdpxAHcC+mrkHdfj3FvkJH5LqRGnB632g
UM55vzM6xQrB2Hdlc/StPUUu5Xur8TaKnj6YDqJ/rx53FDX+VBBjGrIyjORmcub1H9enNWebFv+7
pLk3qXTQYxkxRx/tSs894Vb1SP219Bo9SxNxxwi4y3l7riAasEleybH/ft92myS5xiWnvzuVLqkm
gucHbWCWDP+tCWvd/DCCDl7K0E4WWD485bB2L98HjyKePzPE0sV+N6ENNgV7Qu2mbjJDHGxiRsdw
evGfB6RfNtB/XUtT0F1RfIBvN5A7WS/R1uRJIfDu4pF932XwvI/bQljnuFnTOFF1qRNzVuOIDzUB
37cxDSk2JwTrHyyu5VY4cy6aF28Ey/CCcekZmFqASBGZYsg8WjNDYHcee/Yp2BiWXyu9hW1pJXEj
Af9hwM+dtTBuuxpn+zKVRDZ30WyyqeEWG+ZZzcWVNQ59HsuU8o/boHFmm6iq/SujrgXFDCynL2pM
Gm9m52WYqiD4Ugjke8B1UQ7kJOy6TwFiWnsxZK8CGSgt3GS8C5k8QvYY5r9FPNmKf5Vb+XwSlihq
Gcn2osxe/t8FIiAxn9eMzp7q+8c5hmr40wJe50eBms45SpIKKGqiogkG98iHzgEZHZR9rP5fdeKn
Qdkj/KCcIzetv0CWmabV9ZjQmaKjGsUvJgonXhiPocDeHGOr/dZfbJvY5LD90t0U3gpl1juHLkp2
7QVOscyMMIxJ9GB6PghplS9n61RkgC/kJtKOH/lWEjf33IezJKnJN/qNF5BTOlHsEqefiBugqgAP
NUEjpy+2AFSjn2Rvh7uHeGnIyCTxspfDSjkjzjjmdVlv10U5EuvFJ2Lio4+d4xcuko6FBDA6+qO5
cZWnm0joNtLeK+5DS7kXc36HB3lbaOaujsR4n8d9mb/PaA12eJ9yXUThwfjDBaGkKoOBzEA5+g2Q
nw0Mq7j3EvNpuq+M0XSkwOqOGZWwkK92jElg1FTyfqhSu5nFF7l50d1awonjMIJgDoXsa1W1OCiR
QuGVN55UZ+5OvRpH34hFUUdY2V6GfO6csf0KyuB6k99RPDCONYlNjPatt8kkhwDURXV+ub4ghrFL
+Tfjaxj4kS4W7Ad6sbj7pa3DgRQALUByzVqhCMBYgiUbv+BnD20aRTB6O31ad8rfAgFr/6B8eVAO
ZWB8vNDPjqXzx6M+r65svJbO+1XMZJTIXmbllOoPMR3Hb/cjw2y1MpTbyYx8XAgpDfB+v96xilH/
AVD0JPwhkgGKk1Xqg6IdbPAmST9TVfyW2aeL1+kEhEl4bcrh3of9718BUQQPNvxVixJUGpWYD8h1
NhzWyNux2VYA2+wkdkPcu+hVX/Vo0c7FMNKLqVfY9msaltDE/sBOfdDDzwHTks9YvPxCcRiYEp/y
uYkYZQ+0ZdekZHsmYT04sc07w8unVt+n5EqznOd0qPdR+U7J7DSQ1teqSuQeR4J1cFkAPJQiek2K
00EzYqs6VU22T8ZstWyNDajpp1COJKV5jZHl0Pmb4RTdRRrPggtH0zMgBhZdC+DX/E26uUA/SEcm
A3YY558GJ0SK3MIFDrCD+ym7Tw700RimxlYZzw8cQiT7f2hYIfTOfRoRfaRzUXFSdrVSfWz+lrE7
4rk3mAlEtVZuB08EGLWz3roZPwipBZ5qyUqWqs5jz7v2JWNCFA3Ur3ONBfpOuDfJgzQpHoRvHdkH
8wRJ/tNpxlCnd6MfQN0peDI9APFPlnGT1V6ZGQ5LEiG6H6Mw4+aWcaYJaqLnZTopU49GG5i59G40
3S2PZaznvkvsgpo1XhluyTD6rWTJ9QVS7vPftVWTjetQW35KEEI7+REkoAXikcCjLh6u7UwkSbxl
uKMZMUr23R3R+Vz8DS7faIFhNcRVis5LmPxfyIyY88uq88Uc/y1QXSbWEkqpcCF+V72skDdY9JIz
Yd/VkK3Rs1njJw4IPYp5OiD72UsmpKQNX+0BW6tOSF2xCph/K3qg7X5X8g5vfhvPHGDm8O9+o7As
Rh8xq5ipgNDSa7QiF5Y+Bgu/g5gcLRnZzO0pGLy1J1K+d5fKc5im2mukUHM0LD+6N9Wv5qaYq6QV
FMHjYTKwpWmm+j8zq3ecTHihvk2kU0cqDeknFutzCRgcdV7vRxVU7tFNd7pARCtzonNrruEoZZxZ
650AeNGiEDGVt8ylmEh/OZKJfDoulYhUP72TUYq47KjmN2Vhbpsf9TOsUhalw623nnvmo+a3SpM8
dyVaVOp2eeYmMXzjuWZ/g+h0mfvDkUFg3mUwVYejeE/ignmzk1xyTrHe38ij2NOIU/rmDfQZPBaB
ZWpSLRMCruQpf4azpl1z6MArkWKEUGeeAmgy7f5l78/HujhJ7cJap0IuE6xzRme0vlH7PaG3yK0S
vcXFXHaRgIjcHVacjHNJjUjTsSQMo6G9uwIVTMiLWdsGSsca5enS6pFRBb+5Ox4oIqvrc/JaK9th
A/ulIHvRJ9sruNGxhxmUUzu+LdEzI5PMrqe6PQhYd3/hMlldUpICMbYECgnPTjX9VLb3YLKNIKnO
6tdn/g20HygK20F/3xhbmV3U6X75/F1P1u/m81vc38yonBI/3GKpA1OQIk5V3pHdHI97flbc1JQj
UESMXOFgDiyfuXi3C4CFNiXQdhq77P8UA5mkJN0HvrGiFM8Zzuxo82EyT6JEFKkG6uUKDY+UzxUP
PIJYf1Ko2MpY1DdXhzo90t4Q0xRwjR+z0p4PvrnHAaVn2ifHmFAzE4KIRbSwPlxcNnKR0tSeTFYr
TqdWaRNBIQAmqy7mvN8qE435rsXEJiulNPd36fdSJCkLfJB9mNb7/c87fDNZX+f3EexQRoYT2lWQ
SSzFzxV6vjCnAq3irQ5dZX2eFxV82psjQx8Iowjo+EDBD6fu1Ud8NT2xs8fXpruegChzsXJzJJRT
C32Dub0H4bcHdVyGcKr1Pcos5FoHUx7ZNpq7dxuevsqky5UkNciG7OtQ7TF9gl1p75xCCzij0ZpV
gES7XpafAJB89Cx2Z12YIzxEps+DeqqPUUUphHxnqquvGJE5q4S7pCyIPVhSBvoaSILDe3lp4EYM
4OOtG8WdnYk42Y8ufFOvNGi3RewHAl1rvj7IAmEryUtyno/yr1OztdxXg2fn2ThAUhvBPKcPbxA+
UlwAMpwyzC0EPo8sosW96kCAp/LcUZu9W7dhg1Ixjy2uBZlZXosbM2JftAU8xfm2876OotVJBBoZ
1ODgKg2HEVBusbDqnpkb0yhyjlDaD8sgj15yQLJYg5dqnVptXfF4cqQRCxgGAtvShbbNj1DhtHyB
KG7M+2m2FAZpuLi47vBFVLx9pp8I4Ae8SZX/J+14WRW2YpkqycyK9WhOV00P0cj/SIgUIxwyvLYt
gIg6D+iWGK88SSpQfSjSe08LI0/65YUsrE5q0OtVQDOIgdUmLhruz9uuHw4hG8xV4m9UBKbSHmSn
gMsMElOId8qvWpTnwrAX9vjUXUFph9nYQ+nj8VIT2bDmibiOfciuiwXTHhMH9r9PDk1ilmijwmkk
zciYFbNfibLpio3FrD8BOSGhIHveNz6tjEo5e4vAnpaQjwXH8DSy3sDRi9HKclIXwbsPIHVP0DXV
P4MccGyf8kj/SfUqQv6J3JzJ3E5jprvIKHmQG0VnjH54OwitjVLIqgTYEzCyT2U6nEdF/tZXC98v
D+1DuoSyFSjzLQspBamMA99J9/4JDSBcGW5u+unr6dOryzhHcjAVXCHjMo9h258AD6El+l5Y7YJk
/XWqp79tCH8aCYXkCdiEXJATFj3n3hVia3frzK34jORrom66T4bWkjPCyCoacctP3w1V06H1cEgh
fnl1v41DSdeBDhqccsSlwyzKhm2ypNNIKJaObqRMp/O6suopVRoggHV5lki0NSO4/h+dwMGjUKg9
rGVUcv208NY3hNNaB/9NYWp+GYfQ4UP7LNigVzGFyH3Dsn0/X45ly57ZETqg6sz2gF1w4Aa8/DXN
nDOmqqs3wRBRKTYsrCEPgpuLhlkrSZ9y9+ec28ef8FAzH7sPKG++q5H5vEzsmPrSXECgKxyimgm7
JYT0xXtTnrwvKFzO+kagx8yzG1iIGw1YX3RfADuAgNCJ6jhW/mgUNTDHbzpf6EC2EGshHzV9Fe/1
ePUG/AAgpBewGiTTEuBLD6pN4B6xk3x8OXUhohE9i1Qx9CJJn69uOPGeHSKDMgmfs+YiwEj8Dhg2
cyqfJlNiN21pQqX24OmytHky6QI4gM4VSso72k9FA0mBT5ym+0sHlFjcot2KMroDHhWw/vzrj9oF
M6N/nBXsfCRwDafI//QcpnzUbUyhl/6qfpIEuHgRVVKj17HkZOBBeXPVSpYL4xF/+778OD0FKTvQ
d876B0W3zNTzjUm841zbD64AjuD2Dlk2dFu6i4fX/IlMXlNqFn+M6h/pp3DGXiEiv4sv+qX/S2+x
6M7spM47EslIy6kvMj9A+KVd8omVOjZ2WFK/GQ6FU7YdGqbW5tmsKEDkoBFnF3z2z/JBjD5iieos
LyFDF/zTyMEdnly7LrKrKFqEDtWVZnEbdNYbxqnQO+7KOf385A4x1mLIGkT3hIJ9upWIp3qDoj2i
xCGv8+nbJJYJd4waSlVebRZydXt2SMGilpvmt3nZBjDS0sVcmOCoTCtLuYexDeWoXXjXwYajN6k1
AVCwZci2en3zwzc/vLlhpCGoL2oqylDWjAPmWGdKD7gIBh7GXZE+k0ULZejQqRYnzWwcIznKGqNf
a8IPFzD8kQcl6iqEU1rW3VfxLSFu3RBTln2XNDg9OEMuFfoouZgfW22BPK/5K72JasR1tjua21ZT
Y/oA6vx7ZowqxGlwxaV73eBIBuifirIO3s1KS7ojFtdM1ALqNnmdzTm9FoRmQL+U6B1P4lUeIIh7
PH66bfnNZ+4ZoVJG2w4BhxRSg8dghgNAqxKFzf/xXLO2gljgsfWB/YCGRHVaWbNGxNR7dK5yQt/3
7sA72E/fkl3jxTnD6otj4nWWs3XQCDmh6IASq9uT7/tbkHhMAeu5JVqYZvCAOknp5Aq8lTl+D371
DgPc1KhqIb10aIwvZ91cf9+fRlwJf5dWHBkcVCq4Xx9BLZyP/ZjcAOfDWOnA6z63Rhk79zI/4+I4
zQuKkTxA6NiYWkjTLQlF9Tu4VG94VOzEpfk34OXngn8p/7ahVw/gIY/xTXcsbtjou/r5RcQ9uX3g
7TCyRMVWv28ID9SHeDou+vj+F499T+09lz97OQK0W6yeVR052yPKv9Q3B3/91xxz7p9QAzr/hjQN
7FnEWbhPeIteCX/Ea/zoWXhT5sC78/ffqffxayozNfBlg0xpVvFL5i1LzQaQnyWh1c00EHiC8/ot
4wKP0RtgmosZLIFVvJUkIAT1oV3IwsBFDNuxxZUqzmzBpaaXQVV+ckTM7S75I7bnZxWJ8sarxl73
JaET2vXUmZk730Ge5izxnbcN8H8UTr69djQS18z0XecRubPOeSpCjn1CwWl8nAlr3ztmrJ+BBqk6
+d4IZzNfup7wyM7INZyttCx1ASMWT+pw3LMI/izH+49r1sQtcWc+P6HVn36bcXbCnhyJF93CQWAB
VFrsRsQxmqcLK0+4FsgCploByVoFx5baSd0OPMwd3EkxbXAZYI3QY1RWfIq+/3nig/qxITp4FePj
vqpmzVrAleH7EGrSV5EyTDw7VThnJY6kmZaEdDtPWg8u7FQcDUmBNxq2WDDIiRcnrz+tsFB37sQ5
MAclGuDIIj5acvyST6mpQ2t0VFcemi4la1bkB1hbhrWBR4xfg6Sh2iMnbtaRHC6dwtDztSKTqo5m
KhjyW9vmQDkrocdE080hOUZFArCO0RKw9LIJv3z+KLuU7ISTY0tqA7RjrLGMZOfY2qT1aC9qGSrB
koqJxLP3trmfaakEm5D/vtJOzyTNc/96W5WbWcx1V3N7fCHM/BnvaWKmC1odZ2KAVP8WvO91Uczy
sthhr1r9t+zklv+MPsESy/v3/4ipbkPUa45NYnEpx0lnt+y+cu6+KaTde6xzaGSGaY4g7jHJhd1T
IzjhCjWDx6BqQ0AGyra7ub8qkeORKF1OMOCFAfOzUKrqHBX53cPg1uGnpbKSut5+ZnZ6mLwNWDV3
R1YAkJo0YcuAOZHN6WY1Ub6X5V08oQ0FhmyIFjVBuLZqCuqJYML/0NmdTR10f3gQ+nZC/ULsgWmv
6Jp2RriSLdPKguDUYBQRi7Kcc8o4ZsYcS91P6TuiUNUf3E+dxPs7Qit8rOvjjETxC6pelRG06Nz9
sEoko1kG42XyUqK8JckB+MmVuH/jqEvN4gw/2Q34bBtkKXdHbybDRIQwHX+yGr8YdhEfnXiQACkR
+mDdmyXtJcO77QY7wsCWfkbGiE58JQTNP8SwfCk2myxAnyfT7nw6zXtDVVbp4yXElTJsPUmiMycX
2Cv9RxVfFI/wDDYnaUi6G4WxlvdX3i6McsvYXDFjTz9/fP2FKEYfS25SDAWGawYo/JLJbPLJv1k3
ZUgfBRxyXkB5GojSEr0paugJyQy9rNWy2vEe2zETff2YlFVGxk9uHUFZsgFFBoJTp8n/rZ5AWjGL
6BPZjuj99jzTjDqRIXPbmPVgeOZrEfXpPnUJfMYunR/uaCeFmIy+XjtkeqNUollRSZ1McJKovrTF
GgiKzSh6sJG+AHMyEXIlMHTtrpDr+Jl7y0yr6J8+UA09a7b7WEQSNTEUr5aYEkBYgqRm2SGJ9oI/
nAZVV4vp2ewo2fH3wRQ7NaSE3SVdpLb8vZM1Ul7l3VRKA31aWcwCFL/T4Oydcihcil1EwugsPIhx
GDx17x0ZEzL6q30avB8nORjFUwCHEuy2sMuEsFcjTvAl72z+z/f6o5BCGZvQe4hQfKfMHzEICElI
4x2nOFS9WcORNkC2QGhho4EM/cyF8790wIeMwj0lu8mC+PrkIB9xSGyf8DjemfwEM9knNhNN4982
V9B3hD7BufaZnb49HRXUzpVbLtKe5mSUN5T8OwOvU3oMUama9WrUWpvZaeSvbgPDuW0Lg1zpc+pi
G1/F7LR/Wlcza72s7LB/JKpqvAkLlmMjk8D+/wPpCDmffimshT+ElOPa9N6xAnBUBOLuVF9rTvAJ
fijqa/g2pGG6Cs2q2yfT0byrN9E4RyT8WSxqgISLOhaMDUZrCGMn0+YWuFV8vaSvzceJQUbaWNV5
q9V67bgAlPQOBnGthI6YGsnTvp6MMtjgiBCGsRkEHsscVXKWBZLm7pCl5fYqle7Zd9dj83GR4THL
XJz14rOVVhaS+CuzH20tpKUBveCqAdt1HEt+GwIm0I/brG3cBxHjSGKUPHqPxlAjI8AH4y591RD6
6iuGnJvcxd6M0ZDT7D59t+wChJdzLb0RjIPWwYqmPTBLmSsKVxOHYg+L0ixHmOrNlZ6NkaYCIs33
tWj4v6iAshPz78Rz0Ombg1/jtDIUZfco/1e0PgWAv0B6bbHuaoEuBK7h6PRvoZogzOyaQ7Bg7i9s
EeORf4rpowFDWagdOpf7hUgs+pZ4zHfTvC8eho1stsJ10THsHO/IcOiXLio74RYkuZ8mQF3+qNft
78ANluATdfY86HAIBveXWX4NJypwWqn30rJzBHctG25SrUdJN7852+rVtxXCM421PmFiAq6Gc7Fc
lSzvidzAIqd/ucTb627DMXvQfnYLYUhoL46+0v+oGAs1Fv3ZzkLRD06tj4CyMwNjFM5gTAnkr0rN
bU9MtUHHNqV/9ObNxSw59vP0pgn3aVzndvKQiqGYr2RaJDzloL+6rQDh/ZLI0DqpK7MQypZ6AOhy
Iol3oHBQVC0Bq0qvFegmuAVYPo0HZNqK0M7Usg8y2arSXGPsKQXRFwQG8cbTxBLyD0m/7IOW3KdF
20adc/U/8/Vy84VIQxKylp5MuTw0rS212C8gNYW4KO5CBlCMQsxcuWR4KJIt7ZftckE8SEuqkCyf
Ih18MrdyyRCtYzVS/pHhDqnKb2o+CbnZO5ZOnBJbD8UYTZ7LoXHh8jLATk+xnZpXt1EPo80rb5BQ
dCJ/XtWwHs487DSwmXe+jzZ353wqnDCDKRnv74ICV5OEDFzy7J+rEsdGpqTNETDiYUov/vIKmQDy
Ymy7/O8NTPreYiH0mf4MYKFdBA9t0DgHhYJLhZoPrKsBgzTc3xfhP0aWiqtKg7X7AtPaiEwiO+4S
gs+4HH28A1OFpkZeBG/cypDmHJtx5cCec42Qq+ILb0UQaiGzySICgRiiuTBamLwjtv0gtWRJZ6nP
MCSqTTOVE+af03kXc4tL1m1OKGJDHbi8iywwzBPSv5NjY9QS/ohbmc9AHHFu9SzajCm1M8TZ7QzE
ba5Uq33U/uO1XhliTzCK6aBxwkS2pAdQZrFyuZRUS+/cT6uHVyvt5wQ7O1f2sgoTpMyJapxh5GBu
3g25Pdm+voq+NehrXrGDjGPU8eGHVd73iePMDPkV8i9xuPHA8dWxAPdxnd/DIkMyTeFGoPBLNNjL
qlwXbIxQOHniHYYNXidKsPN5uVMPA0cAkfIUDkws+4aNzuHQwTHcN1BQvWhPhCEikwB6q4/Il2RJ
U/L/wSmrkSpVb0XmhiE5HEH0EX0e3nPNGPxjCorUZOG5nupZ2Sa3bCJ7MaP2FY+yf42jF5I6k469
hoOZmDT4J7EvR2MmafE2M5e/fXUyhJSELszdwPHhKwEOsO7ZaQO7xzBI1xjirsA84MrvvC6yRHLX
1Gl6f0LlRpybbsIJPBzTsveHqpSMAqj4WKRwIYYi9/5f87pjMj/kqYegNoa2CDqkqpHFXMy4mEQa
JJQ68RFF8M1HxYxJUbBNdIr8rOLrzeZpSO50LupOmWh9NvlcWAu9+nNvnxXui2PAaoyqrC7mWj9i
nZPE4YVrA2Tkbv3j7hDOsryMGED5b4NVWNSOBd4RUAWXmJrPIaW0sDVzD1cZ+kLFU9lHuCZXPVZT
w0RzbdYodB+hJOsg21ExKv9G5wZC3oWHP1bxpMN/j4mcs2OTcWHmRMrVmSLpUQ1Y+n+wBVzcoN49
5X1VgRQ9U8MgcqiFgzNb/duULqDn0QlfMDRTTGiPEgLpKTXvws50SYmYhqSz1Gwp9VP9JQnaNQaz
EL5TNvhOyRHY/Vv/Qmn0Aj5/ueMacXSmLF23CO7tZX4EPqYHoQgkkUtfM3EqRuVo4UEnxztRXpK2
MzO6HEbCtOTtSAiTiI3mFHLcbJeHeDMMmM5pcokQedpdTKQJH8GurTiluuSXiOifrOeLdMXVrhQT
jzstH/VzeWM2oWbauxHFzq+9Xx3AevkUl9C1VLQqZrDRKW2Br4rmk5OyKGwcyP4cKOr0EENKiu3/
btb76+Q8BbZRhosJeU4B+ThQh0ZGV2hhQHStk0ak0MriBEfMmRhDRWXab5yfm9vlv8Vnz5bLO/aF
vLetoepo6XDRlasXsQadjW1QDbrEr6GxImbvDG/RhJK2eoymmUqgvc5uST/uzSrvUY8Mio2BajWe
Ph47Mo+j5KCRCoTWRXP+DJzrn5yAOm2FKk7EBxRuJi13dX5QWYXj5BwoJYfFUGipSCXWemOfrj8i
yVqXs7hPL5tIiG3zHgO3xabF1j9sJVjmkCPn9jrhjai/qp/wBDCAnMdw0NMxu6RhngTFBf9ST5Qf
AT9ybuCnLvGX2E9OCKnAZdW0sfNZihpeL8HowROstOZ1F6Q0NKN1S7PQ1EIcaVHwDD2XWdGGD2ok
0sT11NjahVfGgFttHDGUkmf7w2Cs2LloOHZ0TvQg+KdqQfcRGVji+XMM2pxUgNb2jBA12fi7Mxok
5VGi/v6eT6txt5jTDBRLrJi5JjoSlR7JRTId55JWM6aDA1mtP90zCLKH2w2Sh0MifmPL3yImH3tz
pjhutJs3qawpmVzB6gsLbIFFuwfX1S1CQ6OAmOdWoDstXYArjqwunh7L6DeY9Bgb3ZW+FjqMQ1D0
8m6UnsA+hY28pS+PZCTeGcWXTIIWIhek1w9leQIaungsXU97/uQM5Xt2wsFU423w+6kMh6upH+Iu
qZX7RMtABV0O4fD4fDeYuh4vBTqkCcVipPU3kYaI7+tz6y8Yrv88DiuVcLpP01Q2jLUy2sP8kjk/
U2R/LWmDh7cQYF+LXdVXW6RQyaplCXNnLF/srSwhWziT019FXLlw4oIdUKm7tnDoP5jw3Q3Wq9jR
PeikFC8oc2317MVF7+qbZsytSqo8WzUUgSCqgu4k1xkeubbxz8IoDr1oXls+BIZZB4QjhHFqiwdH
kR3ciTcGSM8h7JDYX6C7wC9ja8QhY+4MKUYylUQCIiABVsVGaj69p+pc6gS/MbFLzefLHFEWpwqq
fGXE9A01ch5m9c/y05Fz4J21EfJ4pXkG7rhlf9/Xq1wb4Zfr8XaopjoUMKG6UC4b0CUMFaYD0hTI
U8tJf1lhc4SUpqyL1wZsQXB4YCSTTQ6TaPdTUMsrHttBpiYBWHOIcHws1q6U5GNnDrZ58OKLR4kv
6i+CjbqpfPRW8uNzNzFcKRUjTwNMhRZkGhpegpkVr5kFtm+5d6Nj7eZk8PLCpcNi/aoWPNZmcif/
k+ghTUWnQN7u420K+7qQOLjugBnSs4xv36HdWaRIfhtAaoVAEozCwD99Jhf1VUfImMYz0eumVk0R
Q3QntZnHsDkXJdYQ1ol3ybdG9jXpZxwsg6RjRtjT5j1yo2+VAvfrKYutF6k5VKG/wzYprCMo7gwA
M5+c+/X4uecopYPyC1hTgXGE3+vnMGOHCMNGBlmk/5TjufDVT/4qvTDKK2Qs7C0Hs91RgVC797qr
wkC9HXFznhG1H0xZKT7zontjOJvtlVcAqLnGG+m8jhZYLLjUXTjXeWYNLOOvIv0UnKe8O4lVLV6U
nakwL00eKPG3ezpMf7cK3xrdJPhjZ7fvLPscHQj7i16y5p9qoV/t2+8iZ+nCGWkTuebGZK+STJ3/
ONEHNiq2g4YThCN+8pS2cpVzSUvUrKjMij/vhELzXtL1d/MIhdm/quIQfGS0jL4IKChVHpAm3Dub
orczjvblyvE+giNoa5n0oVj8XIh132scQ4diokO6Zxn/xFOKi0r4hTpInjaOeiMYR5ztOO2u6BZH
K58kdB4/JkBTEoSh9mgJ/1TGy3YDQd1Z/RgSXpOx2z1wucwpcqTXY9Uyqw3Xq0xauD0Sa7OFnhqc
GpXTXEpHc4blZHFNGxDexpDIq6vIG1broLUIGyqkfiuHdf/BA2fwYqe3HFLGJuAkP5NCk5JQMytG
q7w7rl70t5KDQHVD2yDg8QDcTlSg5jXSY1lp31cyqJUBIvaddPIuW8WY6kYph8IFTknSxYMs4emU
ny2joRLVE+bnV+xk25PXDntx7lQUV8Qpwk6fU/ISFtSdglBBpc0/OSTWPJtWISKKGYmuBtWsDdZo
YpANOMFeE3fXQd/+J4U2AUZo5eg50Ap5eWy9a4iZHcMcOp6e0F7ABhLph/iG5+MttzB2tfyYRKmI
FBNR0H8xSi211essaq9MQYQPnwgvmbGQMOBG2x0pYF16hd5+T49zM1Mq5h3rP4w++kkQFJeFnVG+
52/ox37HVFbKnrpOTGzjrfemD13oTWWij/wSfWq9Mf4X+c84/SRVF6tP0gv+SfMHXkrN8njkhXBn
IOjn3qPtBXeQJ9cHpXoaNMv7C2rJWxYZtU5K1CqG3IXr/ZOWSrww9GuGfb71JCfxXHItkDMAp1q2
8kQIF7NIIejndWyLR56RWj/skLQ23X8ARkYJnLjEwkWMXyF4pjpyqDDfMbIY2NyCPgEVNq+nWrKp
O7tN75SwuVkjkNHyphHENyUKJcNVpY+DgXNpeaPbyrL+ALKZvtbFWAkqrmO7ntH2YSu9JZUxx5zK
dxqLXvaKEmTMmwGWw8mNJSe+Hv1XkTlwsCMj1tfE9Do2ggNxL8cKnJAeuLoV9FC6HpHHNIhJ8tEr
9y+DEhqYffOWjDyX0rleXOsLF8VzgVVoSOIuOwpIuIvgyYbQsZjdpGfhiWBcjoT34vZO6npNEwfq
Ze0peIKRGhKRrkPf8TyKzNCjLOOwmsPj8RWNYa2qsfRAnMlN6tDgbKOgQoHb6YGODKtSpyf7DpdM
mcrFRzbuO7ShN4O3zJUYx8+2HLdkeOH15XdgI0n6DD8lrxKYcomolVnqAVp9sV9Xk4v+1nmOaj8j
rtLv6nqyDIxovcv0Q4C1cVURFcdYg4R1n6k/0aaUvH52gVZDse7DutwpzK8BJInn3exULXL+ERlI
5+5YsasQqfCEN5VFfLCbgsui/sogpsd8Rnp0svKzwKFTFI+h31kCKYo6Fah3e0DulnyijhzzRToI
mBN8wXZYF4aDmimprp4VYLEqdHaPcAPMFe0F2Rlv1+hz8iauCh8FwOAg5EW0yjgvX9C14Qzu4OLp
Kdy0GfYBYixiszjhSuOWLN61MbCZA+gyaeAf+QrqG9lv9Rk4wQJyTVh8l79iS9LREDu1DogPX7Un
qKUzw7vuOXAlQ2ASAf1NeFq4uFoJwpE713AHlUoIaJeEBg/wK45px/qpz9wqGnb+gYG52U5enIwl
3xziKHWWs7upcNUKggzddBB6KcwizhG2LBYsp8VLEhrY69uAzvIJB/sBYbnLg2e/Txo2vbJKri52
vUk/oXIs9nty0HfyYvia2mfsxid0kVgzuMoDSa3Pq4idaOuvCkHA3EuIg6IppnYW2zJbETbuQkhk
yEPma9MORtyFOW/vmR0w7aJH7nqNQlQ2B3pFoD44krRYQuDhGLTrmNcSQy4YcWxfOyj1uQK9ijQV
foMvqbEbq19kCnKkNB84TUpJMYbj/9hGQpDoVz4Rr1QjPAWYAkF5JhRa8Q0/MFZYgzufJyDH9Jxx
563m+f14JVJki5lIJIHID54K7qbOxEVwP/Miy7LZrfjlCMk0RAfKchgKpB24BZ4Y6eGC/Rb5beoF
Sjs/1pyFwrvPzP34HgAxNY9E7VdDhvF5Ml2yYsmTCq0wYqafE1CWXK507IpYCDbTiZsfHqypr7qQ
qwHHok3EnLELUuqj+HuJ/jXr7HdKEIPb/pxR2JO0+PBa8Bd222VTqccgfMVCyCbGgfHpXqGXR91J
j4T8Z7UKE8xErRh/OE5uY2Za3ld4YWuSMmg/k0CDVpBrc9zXVzEtiQOjSTXzF1MG5OxDS2gQN8fB
0MZth9TdtySR0tIwvMPIRnQ5nKJB+4LpDy3pcAumTp2Ze7tpDqilSG6Q30n2UsVrzbngzScHCH7j
ENltU2Lb1JFu1Vh5iGUT9iDEpYgy39p429dJWN4VtS5pz8HhdjOg5L3nf21oZL4EzO9LKKNDLeVf
ec7Wj/hNQQBGvJ/UgQk9gMYUONl+N3bFr47cL7W7TeXwL/ORqfuZaQnCEY0dvW8zi/8n1yXC4eht
aW7zQy+Nx8Up/HktAvhAMBlg8gJV9Ld8pn+cj8Vfr7qucJp/2OslNKdUZd7OjSyZYX9l74RPac9w
9XP2nU7KFspn48v/UqblM6lrCz2DdNdcxogt8Ct5y8oIcxXcwsYsThxekDxVZfh6gaatzBus55OX
ojbTwRRrkvH5nCvVksbMWWW6iVY2aMkytjc0I5yztDHHxp+kvjMV8eO6snFG3SR+Reshw2p8kyYO
P1ef92hgRUkeMtXuCKe7d5x2Ry90S8ZqlSA8Y1/JG086dWsZwg03ghavYIg2689B1lJA8sVA5LCx
3Qx9gmSQ96MHecUL5V/YY9Jlhe2cVfZUwb9+zi+JsSqkTWRpkCq3DKNxDSHS9EAqedaHJNIR4gtP
Mrm7y+WtYCSWWZbEf79KcLK/fwRf83BhgfUKIpzCHal71rh/bYNn6Gzm6LCSmYNsHSKdJKqVO1qF
G7V2n+f+5WEgw5uaiFiaWy27elbuRuYedYKOQ56usR8ruz3PaftepU+2T/lTRF3Ffgo2PIUmGHPd
7e1DZX/yJBFXig0kCGAOox6U/OZ2Akgot2RfxLF4DyVyPJm8HeKCmLpxSfw8euWrMlkK0kQogu0s
KwgYU4fBcAbrgNmQXx4m8ikRw+n8Sp/XSclpBe72Ew5Sh6rtziYS5rvo1buCp9u5arrubS5ha8JL
FDOnr6XF9vET4zWU0lH2+ZzuAjMusvGqvsuRJ+YLJ0Bov0mOGR2FNYCL+BAOfdso+VtJOrPfSFMH
IZXkChD4R1f8pC1IwLAQ7toWGap667DXGU1TFuOW3yo8V5ka5lVEM62IRP95tsKrJtaOk7hZoBUI
W7ruLFGpLb8A9Ng+D0xQxnG1VJjFlDpron6wR2VUlPaeUvPbgiuL+5hp1xPQjOtgh/I2QNgIGch8
MzxJZDiq6IZumgWs7uSS5XjRcmXraDxtOHMY3kK2ilT8y72tC1dAPxHaacKii0AdTDoML4KOkTE5
68h1o9aJ3uV2G0C3ZiY1XZYGz0QdhQ3/7gzGzlOT8WQuvZhZFzsWehOYDOmTWyx7U9481cnT2wSC
+uk99kO5E9pvIhPsGqeiiqw54RsFA8ovUpK6febaaxkkwe5E0oBqHQJy9pPPuAXMlcZM/5AMmdL9
e/NFxlP0T8QbKnUWfmCLKMQGVCMXjavL/Ne/3vS6InesCA0DS3Q89QdIIvPSCIqNN4wyremSLI4r
yhsrNWioNUhRNqM0nRnq84YMp8E6obcNXCct2/jUwv/JZg44oNq/PPrRTV9W0o09d4Ub49D7xgz4
uswUtQpL0JqHVOxGVhy7QmOGEcS9Mo2n1ik3ehUy8LuTgO4NQr0/huN0N1toRyEnA5cjJzTmuFT1
xrwmskMOPxZC7jnO+gP/8uoY9l55KUtC2FN0CYtaBiVcjuqgcrB3CSLoUN9/b6kcABdPIBeBER5W
YYKZiVMh0CpGsVdArW4rPSMM11zdI1SBGMtUjjpC1xm5yTuTuaEQOGTL8RbvfDVQIyZ2e/tAfj7H
NHs1Hnh8KMz5FlgWZU6TrmQsXt3GfcS7T67j67dEqJdRiLyWlq9+tYk8Gcm1r4+tcr9H/eSsfA0u
ddGGA64V79KRoxZslePudRJMyxvmdadPPsA29PTlODmn9pphdbCswlo7+qVERmM4OwXrDiXh1J2m
2/ojVH5KEIAM9OXRJ+pdLfdNeIhEjlVpvmz2cLRmNFfwM5OYOMVDzVh7yz+TCvfra55wFFwbwFw9
21OzniHyhHw6SRJjmk37YMfNR4gqENSQubBrk9XBEMk7Gl3KApgAqQwthsZb8hBd+IwKVkge4+bj
9e7Tp8vz7YNVXJCiaI+nj+DFOHVL5Vi+FdF8m3d6n64sllfsmfMYdhFZFpv8iI4ByoHOcbU/0Af1
zgIg+MbP58wMPvP4r4vTone/NrjYZkYwW7yuPtXCXG4d1958f9wpEZqvkn2DXY9ixfe2YuiyA8Wh
eS9di/BWmrEYq/ZK2DfIsg2EAC0G/Q6PGWEYoO3kSKoys+vq9Tv4bh2TwN65cZW3QUkd0onlpQnm
mUn3qaJB0XapRUf9dsXlrhpdIabMFCA/8rXTVJhJKKjV31KUMjpS4bdYUffPlkoveW2Po+r6f9h+
hK78R6dqw/mROQTXUFXbGlhYzpyVNWYF5wAw710po9oOqmsQm9ku/tNvkKzG9+MES2oK4tN/ivOK
ELXhMbpi5lSsm/6k+sWQajdDtBg+UARenuHQOGCBUTpIZx6ORPo3hrtYctz9I2u/up5i4wqiLg2+
ErmBWdNt1XeA8mtBI3Gq8pTUokCVXp+3YWHjc8vLaNtjC6gWvZH0rWFnHDPjKmfrpIwPbfUcO6LR
gGAJtkFJWvErSlcieDY4Ue96CKQQpgwnRpCcgoK35Livt0jXSQ/IsjtYh6rzbqbBN+/QPqtb5yec
PlxMWCOxtEdujjZ7d8hQARttoLY8Eq7PsGXEMHgLPer6eUQngCJ64Ynrl3LvcaijE8LAaSLPqJzI
YRAQm3zOXgPnh8VKQlPx5/A8gG11KfZxisST4nTa0ttbdzqgKooOf05b5ywbKRxM30jcymTLwy8K
RFh/gAOQIaC5NvJs/jXviqSVGSIx/1CfBJfRuNyoUD3DMwUyuRC+dLUIL7SFBE7Sf81piPHroLZW
yM3X7ekXe1bWWY1G9z08rCu8MUhMijr4on0hMrYSKlZnFFn2jZNpnrObT3MQo4zwRgqrzix40a0c
kYdYbkUrSDdxfC24ek3vUtqwx9WuOtIZjwcEsgXk8QPdrgcEcBQ8eVFg63dzAao7oLxYYDJuIbOV
N3a93Evl+yH2bLFoFOaQvkPtVbE9Jt98WG27t9jUyl+2XhjxLAY/TkCkIZAw79kVsyg/M8id3Slf
9iFSHow9pmZcfiHNKgVDH1UT6WjjZgbRFX6P8mtlJl/9oZwncXK8TRgMtabyXLNy4hV9RbPbZbCd
G4tpqjKdN2BHibVM7B3ywdknXRKmMckYrxCFfBuznKjgxlkRLA2f+40LcQyEe+CGkcToaf2N9StE
csn7ko0YB940THKLRIO/0CW7jVl46VTzYHQqNke5UGNJG84s4ic7Ck8prb/LvHrwNpfX98cUdBc8
9EW7GV4FCcVzbbm+D87tGw1Bl0CLGPzz+7jodWuegPnxMy8Q5k3rj6FKCQTU3r2CJ6Lv2aRwXW5y
3nYodZSiU6fsEfWMAvKKiptIPf/j9PAmHyH0co/omisSYq1UdfIjO5TIsygdzzc401jEIRLquh/D
x211iHZFaA9VS2jT//GvEDojnnnLHzYjR5DwoHokEqRc3E2zPiOSbG8gntIfZMmgogl8GjNGBzdz
+xhQIgIHa3RhP/R9xDBOPn01wlo/1TigsxTsBFGS7wPlSLjwOXZDkfcU4ww9XG6aGw695Y5GA6tm
nqNlDF+Clghi3rux1a3DlxGZg4RhxiPBwCBxQ+Hn4hZ1QnY9h2aRzFJMSQ7jVLVb5f5BH4vOkWcJ
5iXmCGWUHXaDPVvD6DtfaTnl6YA4YMkscIEAJJy+3QrA/mitychpDaovIB9KDpwzYzNavcD0CFAp
dfYF65HaQoqyhShzQ7ZosLP3PbQGAmSE+Yw73r80KBOUGjErcKsm5A+J65GkkrZV9xYx1GIYrOJr
3CFZs/50MFPgygzVQik0vTFB2DFlRhDW07sSHqp7IIvK3ge7sM5MWJxUn4liVAmx07ex58E+l44d
6RYB5HmVK4igYDUSvPNEUM/qaNcNnmkd6pldY9LYcwRlR5GJjF7Bj47agvtf9yRI3sysW1w0Hj4T
pxCSH+gWwKm3V4QT0zBMQyEVVS1HymN5+Cn/di9v0Vdo7hQtirsbEG68nROcCHP0ilXVDANy/9EH
4KdPuJSZVsQW2ITCVIgDXSx1DrvJ826AI4lNFSXIXm8PYTpeU71UaPTZ83YvmDOxVnbzln0lCTU4
P1Kk11kfAxNDGteqIDAIrYrimG8rrGUck/a2mkUOk/lGhhAlkcRQwN/uqFTzFlKcL5fWlhfPVfS4
D+72BIMiJTVdI4t9mG2Zug+0mCXvVNohl7on+e4j+eYXdxx/VkxDnL34XBX3QK2OY4ilD9D10+ue
qzAQeTXStbRJX5GC7PHEftwR9yydRvxc096tLPswtObnDQQKpt9jOg5JwdFgqF+XFOBpct4fuzyk
Ex2s//yAQXxDk+SL/0T41E7Qu0bjZWsty0r22ZHGIMpve6z2tgapwXtnOpZK2+SM0kw9lTZ9u3E5
ddhs6AchWS0wJMkOo4iDH/abHTv6utHu9PwhCtNrFEB0bYmLEQsckDfV3Z0IDLaJ8umFQFRRFr0z
eNFxbxEAt6O7iO9/cuSIvG9Gqkp2ja7vKMGrq5SKvHG0R1wbydTQh/iK+ctXo9MfpIwljksyJVKf
6MapniiNAsvLke2vthBbU27mRsU1oZzZ8fyBHPdUsWdBQk32/qt/D/aOViu5Uxq9vULOc1S6CzD/
FgyWsAD0zqdl/XgZ4IFHjhaYtAZhNbvnxYfYrDJMAkldqNZWypAW+lCgRh2g8sQMQoYeDTH/DxMu
eVeHNjNlz2MgjvodXSML9C5w8DQpwrBUkV8ibB/nPkldmFrdBzNUcfptt/UTNSKh8skgTR4XebXE
t8EWBX3veEb4TClUKthbjW8ExsLrgqyYCJS2q+tiYst/MIfJyAwXsoXKgFGwwpA++4Zah7xAR5CR
nrU60TC/nqd0IimKmokPS/toMEsqmh6K2uiizsGFekRntgQZeYMheCmrq6nwySxUhCcpRDe2jz/M
W8DIxZRtgvmhunlvl3nvOFUPGUu8NxDdrObsX49b8r6gqhhMcL06Izu65XDxVs9CR7xBg+ebCRdf
sty4AJOz0K3VqoVVPC4bXJ9gwmOP7BlZU3PGMsHc0pfKUHF187/AhY2EIFCm7RJOzDw9kvBrcK8k
CtbQNxJimD3D7q+uODMwqiBH9cG9oQt/3nWRqGiJe8NnX2vH6l5ZrYGlvUMIQp/DuS4BqZi7LSe/
hJqSGDcSj5culB3agRJqxMlsBWv4DDT4i5+fAQTTxHfNNzcirBU3lgdu4TeBfEDqguwvTctPc2Q1
Aka528pZkStLBNtwtG68gRbEVIWZcHkQkLTc6nYt8KublJ0toLAuaKBD09CoVXXG4dqQoGtkBohl
AKIiecvBnRJPXkwL1V8bWAmPRf2lwmFXl6jCgjkuzfBclXrOkZGfVMMAZNNTbQyHjbws3CKiSxLL
JXatFblfvLgE/OiZhmI0Ip7ZHBWzwd7pybsCZXvfQFdSufSVFYa51/6BYBKgOaBPmUPgmXwKst3M
buHOAzNhwTw7dDLKQoSRQuFEKm1h0MuyAWTt+5oVwA2SOSASGaDidlZVZfIwF3dCmnyZnCEj6mEG
w4Enm++ccFYwjOuMWduSUINYuDCgv74sMHflV10RgjXA0n41OS5KS/WcfZo+7IyvJjmKy+wPGCx2
e+iwvwQOeTX8bMyoZCK5ycwLiF+9w1bkNkSw5CECRvenZoQN2ZB6dozQqWVfRp4MLpq1l4PKbAqA
u4EXd8Ul/yp9sktsPvn+dSA2/ZRHbkZM/APtEOxt6kWkYqH9VbmXrkO0nqDoMQV0a0jZ91KCRo1+
6TRoyEF9kwnbiJoKaNmxW0fkSnOzcj7uIv940HghQhlZ09IB3GRF4zFJiMnYChkYBxaMILqKdK2w
xZP/7MPibgaXZRQWNqYAvqS/Ug//qwSgsOuZbBHoVkXLob52H2Suv+DBXnCYUnKXNmdN+MYUvzeo
o1ID7qe4n2gVhW0T4jSJNltK+lvWhIyVWZtNpF4R7OKbh6mD6iDG49Ym/25vQWrpBJyntU5P6EAe
WeKG7Y4upHFlRFwM33NUZmj5Jm3tpazP6NreP1gchyrtHR1jCdCDyAenNvJ2ucFEC+Hq991gVEHk
THcmle/Dtf1dxnOBfO2CW8wfjPnEbXPDW/uGcgCJUeKA8/Gedh4+Bmc7DLpIHtaFaQP43/WxZOp6
C85449uhJO7umYYwi87ps//VLi0UNHsC9t1QREurDNoCcWJHXmRAu3V62rHQYHX8ByN31SG9u/OS
Eaylbt25PU4SNMR3Txd6cZhGj9IdLfvoCAqtWDV6tiyin7OM5gFT5sHmO5yzRWcquSVkuEJ/1t53
dby7jH/iDLq3Y7JTy3A3+ZFpFUXo15vhqYmWqNhAGg02eCCbjIfERcxURNNZXAOqW6hzHYxOL6oo
z5HNpDbPnJZsdbDEOT139gLdei+h6D+aSIuBxq5hSqDYxosio9pgY843q+ke+TQ/+QveOEjB/GQl
1CAkBpYuLVj0pD6tAxbKvl4Rr88sPHZ8NKm+HlZydW5sxPZ7l9GpComdqr2zG9RVVRSyVu/bLACu
DJhygRzNW239heq8RckzoQIq+Pol28bzF6QB+i+jiaB6acYyqqjHJOs+IGcbPtsNCpYlMGFm+ULz
imG2clENK4H6LEoRL5qoZw77AzHM+NcKtUUiSwzDfFaAv5YwJyED/HJf+kb6EvCG5bA2hw5VgbB3
3Beb2+f6WCtl1nG2vKjdnhgXs9ccpYAU3+bYfWgrbGCffe+eDBgO4SXdH25v4BwiWoJ0SVsHmBvf
iVQXZ3sKhZMDB+NMpWgLix/EACZPdowyKyYDqs3JMG4BEaoy4hms5K6q+hzK3OnwCnhrcM3R6r0r
RRNsdQE4sjgc5b6atRw49hx0J1iE8mGyRr9DxCjjl8MOmDlq3DANE5dwx6x9UJEU3oZKaVRmBwdm
pPGAIwwvmcaBNMYLoA+ipF48PPbnWeOG8lkj2eFE4rqdd/XgIo8Kzj1SBLt4wQ00h/zmFdgKFmQh
UG6cB0ja8wA2KXf28RdR38p0TWkQbRAhYEJswfnhrYLG5xo97BGOvxEYSdbifkTfl4nF3BMwEZBY
/UL6NMY1cXmHrh2e9YmCOQpIz9m+QWW5cawWj/CobRhOI98w4KVuaDxPfNoyGPrXMk7P4FfpPZJN
45VLp6NtmVFH0Pcfj88CgzhuHec7kpWQt3Ve5SCMYnW5ghIXnUlzy217pXhJYyM79RAUm4DPTIW2
Y4jlp3re3PQDs/SS38dvJ4pc1FzJ2Y7ld698QQggsiy0K7TlPafjPxyVIsGEjNXdun5sMaI74iLZ
fLbZvivl8yIoU0igqG8E6FV7qgDoF6ejaqjE3nlfSv8g2A48lvBgleC8tybPBFSzZsYrXwlflM69
ncKvSdV2yQ/6/ttRXZemtSCPMiCskfSPsksIO5yMeCzo+HuLA+VpF5WqlMv1V3tv63I2W9sn8c2k
1QcZ2sVUdLURKsZyFi+diUacnZQz+aC2uMjvMxQFHRERCYKqGQ6+KOimBfNd6eammiRGl75neSFU
rcI7sC/7XZGxrruWQcHoarxpw3zjKNWfM2NpVfkiIZPFxqxFosebg9nn5J11ncvSAv3GIi5b5UAS
Xbmz8kwT9gz3cyKYhueFxRb3C0tjuc2S/JbaDVYMgdtnjGs8UkQ9SsgzVHWCD0LM5NyeywqKYCMF
EPuuDqxNH3l1Ok1685u24PF3aWWNF2tEiStmRsMoxy3WFmyICmkS3wtwbKkFmmIirsga9I7ky0y+
X1vV+b82lj4rt6UrYv7JMp/5FAw1NzmBFQv7ZZdyqgg7WQ6XRIg7YyvU0QwbmvKuR3COuJnQvlHY
Omc0cQRKZG8fmxwVWl6DZDlrB6T8tE5AqMQ8+lji6WYXHiNwWrRnjBhsDVjQ3Sx0hFVlnT7ZQDD9
XmeEZksIwWpne1tr0HYMKviA3LF3IgbUeiZewQGjM1/QSqSFLXwzR90OIwIfLOfS8DpLFprSvhX5
G21lzHpRk+JBIHudOrs5HuhNQAxsqfHPfAD2vKwlnGyLyPt7T17/eAOENhehIUpbgCWpEbEQg8ha
DVAL2MF7Nzcvazko8wfOdeicra+JcQYEMO1kkojJMOI9wu7u/Hd1dtm9sOv23MsbhCNsvUQH4/Y+
evWCf8SS5EKAlYuYg8Il14GazQJ1LQ9LqGeBFIU8UvZ9Ao0YRajOlmDJO+V0mPpEY1Tq3kTC+SA4
0nXpAexsPeSV98TMuYTStsc8OuwyM4iz6ZDbuO/3c9P7F1P3LcGcm9qqXqaZXlPnJ1pTacqqWgbM
U1G2OjH5mJvUT6D0yU3XR5Uv/kulvKCnTlD1+irJIIzdbXZykwNvjJRgtcH51++PcHPKm0Bx8hyd
IvH6Mc8CECbIWizh9A06LDOmNpXxoZGxTNWFx3NA0Ahu0nyAYTHFhWu6ihstWwVMY5BKGq66JQCl
0G6DKXVSt6jI1i7xNelVk45WmgPqN3GTFWM0/DadDVA/26qfJzAu7Z2Qza3TEc6Xd7uME/NS9o2/
JS1ob+iuivkHp8vdEwchM5xkayJIVrWOT2yH2TY+RYLbjmjfivtp2D9p60dfonzXO1LlobEKesZk
9FSr6ubjWNO+FDA8TbaMeeLV6ouFCGgOlpf1KaFKz1rA+cVL7YSwAV88GmiZhsLx8cbWcZSweRpS
Pd1Kj08UcqizBQJUpJ+5nb7UzD8wDrU8OYf/Sz/tgaKWIkn4Kpm461Jnw68s3Ih45k79NpnO5lnk
kDKJgAKq20KIXnqnIlwFRHnCUd56WMxspEAZbj0st610POSasS/GN4w3ynSynJ0XBQslAHYUY3w4
qdDInWTkrzP7ogVU61OXEnaEIHkb9/8P3m2zdoUWPUUQOIttJIrpv8W28jLC5X6Eydy/6NebYR7O
c8prOyjjGo7m0L3PSfoniqirT/ObgGppv37LkFw7Dcuyw7JM6KedIzvyE630ZsFZlLALQw0pT9jl
Vl2gClbDYbsR7JUqygdY4pE2o7wwaJq3iceLvg4A6j0oLi2qMOVlgoomHr4idGHAfUGvP94dE21c
7ptcx0r712nETHnOGUwIo4jPlE4n10Z2yW2tIdQImqZ76QL4fRuSGHxbNmNMp9ySDfrMm91R5d2h
6YEMwVWfyP0hI1Vo3T3JpNMPoSyViCcc3dsizeJ27D0oeyUVGL2fWBRlmGQwpTfhaolMJ6GFQ38a
5kcnnwkk1gzjJ0743m9/Dn35Jv3lKIO05+Zj/0ECzYl4H8LoEZRWoHc8N4d7i3pK6J11WYzCXfKO
AhSHr1ldzp58p4VJI8Ga1dxDYMLTDUXLOcssjyWW9XmJ+3ldjuUpQxOCUjFVSAvd3jfD/q0BqV1h
xSCqF+Aeky+mVOX1D56It4B6eguxmo7Tr7Vidrw59349e18zf8+iAEYGp6Saww3WilsOH9rrLkg5
gDeK0qNghFYU7F/KdhgM1WuUSg1shoyqtrEZxlkApiYp6+NLUHotj4IB67TKSdFucYMECtabkLOT
h7ErsmKH87yHbc2Itt2rmF0jtxuFnbjiYmiqFZnWl7j7opBqbW816+iP9gpboXVZLWjoKDB5xUbZ
7g9rqGzIrY0TW6liINwNQyv6FZKkdlFnaddpumRm2LyiwgRCMYY801WP4phoQH3k2o+dcB2TpW4D
YbLn8MK2fRZ/lYHVu05rG0Zh4t8IC9mE9qRHiRibDrkL40iubs4Ul2JaSVvSaxHjVDYK+DAJJtnV
v0B0z8zYtNnTuSfUCpjIkOhUJTUFj/QiDvR0FLjstZ+wziJvJ6/pQP1DWB5qg1hWs8YrCowAUjyo
k4F+TXVQP1lJWyoWe12ye6n/m2LzaYuYZPZi3xt5w++Ff29lgCDU+PKP+up23wWttJGo1Zk2yeJc
FcmvaGw=
`protect end_protected

