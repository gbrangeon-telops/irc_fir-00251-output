

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pabZO1I/O5UlEfYaQEPwd4l9eUai0bqYoMxFZDUmBPXyS95K3GW98Ld97MzJKAXXnSlf1PewGW2v
0RIeWd32HQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MnYS98CLv6GUlLtXXj0MDq/aXJWBamrEeFXZFkhzX7OjMU68I3JzEc2/1UN3CHInfTII6cQBis+f
MSPPkhHYfjWA/UnlZNCfIbUjCA7v4zzzEDOXLdUwHhey61M2PDbtjo4F0M+PSYsHQUE61FCJYZr6
+aBOwyo0CpKkCUVEbxg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qncW/Cwz6DQ02ZtEcvyp5WdAA4sItotGPpP0REUtLyqefQhCtJmFILcg4T0iyRUg7VuYEwIANO5+
QvHNNc39qIJv9lOesalgHBZQgvNRJnIdYWaRfS0GyacwI/2JQRwAkuAQstvDCp4RTc3l8lwP6/ls
9Kgq/wnF0FIDD2zIsqBFYPVau5gOg+E2Yv8daLhsLbgUNkGI+w4/OZjRbQGSUjwZLuzAjcC7dEzW
IiD8iCe2E3P5aTpTA2tXeuvseQy8KOwVCxJQuur+f/bmnE2QrPi5PPQMRcOyc4ok7k5U/64SCKlJ
oITfL/xIL/xwZa26tMPcLgkkx7p0G3RLvL/tVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Dnf6vaqe/V3pNaiPDsCpL4mEkUhuRTF8jsptuAsYR5QlsF0hNdnCfK2+aKM5H69faCvd5mpbM0GP
Pqz+qhNmOYPHdckgaTUGR5o/7QyV8YKLvzwfyDMqTu2isTv6FP6Q6welH2CNBnmC1/h5T7i+fy/Q
rlaoXYJxfrB3B6n9clU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IMf8iBP4Q72XIQn7cHjsTbT2wNsnwrpqWy35OTpGthg9IgmIl2PQf4/c9imtaZPdkPVpIBywT+vW
p0seCgJeCim8uHSlCA4Yuvzi7NiJqnEZtjEX9xSzaDj4EflUudOJTsvuYMqv/3kxvUgkIK0AS+U7
CWRV3RwJIjyzXaV3SkeD5i2xf0d/bezTocOrvt7wO8hz1n7ziicW5bgdFMZpO18+84bLDi0MzKYQ
Ad5OLz8QJgoCqRTe+B2lLXuByvKd2+XBYArz50J0pDfy4RubYe7FYpZdW50ze6dgBWVP0HOw0tLX
Pt7eQrmsKxnIhjnIQBRBht+Bb5QLkHSbaJnGbg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8352)
`protect data_block
nv3gr3ubjO+GNW30EEY1gPvuX5MVbQLJvsURg9qK18DTCew00TVKIM+7UbNDTwpjDjjFWiBdZ/ZQ
jFXfTCvLhBVKh0S4tqfCA701I6BA9DiJUilnYpkogOqcjqSxHHz77enE4+GAwo0kQwIL32UAq1wv
I/mRHRbtg1YOVhwDAd0RgGR23a2K3kjclLZiFxYR6YACDx80g95wDOJUexsJ32g51wuRaEsicLZT
OcdBFq2cLUtXAEu4aNZgo/mL80zfKwFlKkzGFjK3NTimg1ShTx0mxg0Y2h3ir8zu+z6OyipGGSV4
sw2mh5zFcOV1BsBRGC4OEz5CIaq0Kj8yeBl5bEqr6hH1OlhYaDukz0/0GA4Y1nyJGqDZ2EguAHrF
hsq9w4vyL/Gn02XULtkNdVn2yGnUgDDkg7/LgHLgqw15eEPMbbXnbfUsv+L7Iolsl8cqrWUGCs4D
0l4QJqF2VqXqBB2nt0lnREvpjzUbkgRC+TzlVjq83bPs6KGeImQiHB6KMppvvRDYzjdEAZfqfTge
IFRE+d5wVAVZnwjhbX504lHlfTvHu8an/LhAMIry3rwqGiJnHFkzFWpn4sAfgI9VwuPT/DhOBU9R
5Oq0giborElOXlOHZLGPJ1WuMYMCoGn22V8OcimKhQcU27fcAHHeZEG4nZueY6Lt4jfRcUItNKik
OQUzm8++29FBVFIU1OD0vnMTRagY8ozUr3oAs3w2jjVCfDJMjRsJ8YbyeuNK1AoLXZdB73OvqCt3
tE2otRM666NfMvt8lIKvAVHWbmVJWR3UC3ktnfHKQFVarShbXGAVqY7Ib8sD8tU1oUC2mMt1PYDC
+gSW1I3Q+MZJ74LdezS9nmywBTyKASoqfpMufBsJyPsJ124z5+//HVSaLmWzx8U8x01uAuL9dw1y
xUPGXtEEfx8GUPTnddDZolPsiypsh7xIjlosk2Xty3cjGAaipOkrLlkC1W6PCAIiEmn9I3mhshpU
7acJvRXtzTM1rKMNwraK27+l90FJY7e9ppTbiiuRlB1aH4f++JSfG+InGDGTdAOYkD7eb4pBlK4m
ssIlcanISJR5BKfSK0h10h/Ij2w5l4GvkMngKTSEWnhFbd6nz5x5wWtHn5SXx4Cli43cCuxY/oz+
hA+IFaAGDxVoi7dEfqjrIkAz/b34EC8FWVQdWyeyx9OJDPdOGQQClHm6tgu4CYjK77QLNVcus36w
exLmBhQtOi9zYoQRvhx0JJMXm7s2we1+MqINSAGzv7nRTbDMcrdtnpAvs+cq6Uj8yFOolCyuwgyN
6FQTSEBlxuKSJyDTS+M9p4OhJ3Vq2l4Whx/E7ZsNuL11Upbg/kKz0b2ZbH4VgS1LVICzx6DxT6Jg
wP+7U7cllCEmnOAiXUrvxRscyAkMwQrqa3uItqlxZ3Ze4zAvMrA3+GKiWeZVuWmnl+hDrmJMiFqj
VmDb/vOx1UiRiOVfjTLvTTFLoeUE1EZ1e4wpPpHzUl9zOBSnGYazBqZu1jhnSDM96f6qKEHSfCMB
jgNLQtxbBALs9j5btUyJDJmuq2f5FsBRUtwA8gca3MYkzC3aX/sq4rewKkDavK96E1/Vgb7cg2FA
4mQHQmKsI6GjUH2p5Xintuw06TKVF3xaVv5b3D8CEs0uhFDSU0AAay83/feddXRXu4zZks0wntj5
Z1s1x427GhuSZdH0QfeN4lMNpPzMZ7GzjzH+catHR93pMNCBEStTRPx06CPZQ0a2Jvh9T5ybwQh9
gkNmgoz8OhuGoyFdDGWBlNXFWdE3CPSfw7VxGoz3GyYb6nFo7E0+YYsk/hvlF45zjZ79M9pHrp3T
6KZXFT892MdKUZhM9h42HRtlxBQnKcGPJRRCiyd73YH/4c5XJumLn0AaNqaWC43hYpoOy7rgsVHk
WMg4OHkZXth7cy7Y+IzyOlHlMZ5ku8F04qTB1LfMy1Q3mOnYhL02wOAHzrg3gy+Ct/SpCS3B0TmN
fD038/TQsFV8DZb6cX0vDmbUpynUtThMagzU77jcdWBS74ZpA6EiAAJsssZYzHlIK6ub6e2hlaac
QQgH82xWwTMi2/ng3HQdVPrYFMumSi1UnD/z54x2i36PRqQRt6VbBnfn0ZU1RubOFAsWFbgh9VPw
j2BzHmfwKe8T89g3BCwmdjx/rF9CBBdn076qrHlJdemR5wrCVJjN/ZHi3zD+HsunJ5nlq6IGNc/I
RHEpy0J7rJdAxz2KiBUADk0LN3ChMS6TRc2Y9+1EF/a8hd3NQdia7pwlHnn+5wFNfGMTsf2SnEiQ
gOH/IWg5k+eQPTHW/zp0k/kBMNDYPTwf/2hDlSY3wsPfStRYPhsfyj/GZqhAv55URQTNgklYvkFN
b2ofaQ/OXCujOdcMc89eDKqbnNk1IUtesbnXV+PqwaEJ8HLhGmCrHLuyNXz3uFS2oMV+Lhmf2vRz
NrDTw9WkdHG8p1sVFaWdvNW5BlMBAha0dCLi/SwTSaSF9OFH4CxEvNrPnSF/RgfHbD/sKspqjYHw
lIYMN6oA71SMUXk3CDcouTcN9FYQNT+ECMnIT43phhiQne95IDyM4bIK8qQCZVYoKg8y9G8M2Tj4
TA8NgnMECJepvkU9PrZqPw0IRYgNA1uoHhtuCqVS0kj0o6xo2Fg2uJBTJ8VestEJVh7widOKluiW
YQ0RdG3LHiXTYYwyN234WALuoAeSOc1/15+BlZkVacMx+mqoXgiSP+2FoqKvd29QJZsATEche5Bm
1Ka8JPu1YrBnikkkrDYJVWMCgqJLowVIy8DOYkgnEmDgFH7TB9hMHpZJ6s8W/Zi1DABPpmchN4C/
XpYkz8r4QCqzIpVI1bCbTPe0P9nJi4hmOTdwa08Z1pBoYNQZyazj3LoaYnMirIDPuRdiA7w6araH
PBF90rDY7Z5fd/B0SjwHjmSOiuda3ybI2oyTtv9gNuyTI6riVvlMEXzhgh64E7Bp8LQwD+FCV2WW
QV0CF0pzinT9F72fnVudxnytf0KqaDrfKrSuWV1WVyyYjz7lyM3bJgAg8QWlIA0fvt/4jKuPEaIX
iE0SjpvEFxZt7Ij0x4Bko/AiROLIq41dqgMsksT4DV8dFC/4RP4bL+Y/KJdpNXmEc18GTvcROaaw
Bjz2Ze5yga4HWYYT8coco14Wb7OR0felDvbc4hmn8PJZAvA6XynB4Kzc9BnCL8UyPSzPweUkxyPH
hD38kU8wwxkLHM7ZGMr3OgYZYJ9+9wqW5HARK8YsR09D63SXoPAtVL8pXPyxFZPoS5VtW2UQGnUT
GZwKm+PgEDIbKMqAhLxBFuI9hRqOgwUE7Tyg1asUjsA5WjWgntipJWtpIfmsv4BX6hVrmNqsVDf1
xaA+DuGWVNZdWU2zQE0jDFgW4gpb1xzZtOxn2xQxAV3yAwF1zaKjiYaYyf+Y8UiqxAWzGgZhWGnk
KT2R73T7v9AKEyHpCGtIuBr8NPYrkkaPsElS4tjHK/3KehUCnSzU8cFryX4wAU03dQD7ehqurNAO
zFCME9Kg/fmufNwFv+OuCC1NOe7tgFF2bjC2oagt9Uo5d31RpknYKfGP2lev3g6LStKA5Y7L8Fcd
h8Z4OrYN2i1B9A8JnOW5IV+7rkmQGox/kqdsi7OFajHt5LiLBZBK5sB71RnV5G+M+0y8WwLX8zWE
4KCLlkeOhqR46v4ThK0uiFP2J9hEvZyZK3eG3ajpVaokazfX7GQ314nPZQl2Z4/fitQr2VRXsQby
efpokc/HKRb3n0yG0DLeie2uCEkMlyasGlqold9CaXbrqFi7bg3HLQSHDElxgBxRRd6Uk4CFfEed
3Yqv/fonN6kABbaKxFlwNQDF7Ye3QrMlBPDNqCxwRhz5PhIWefYYIRTERgdMVm8V+JgL3wAsZ6ho
xEFrk2UKJzxclxK8Gm4yXqPZWMkLmtKNij2IH94JUmO7NB9rPbFLj6X6leIxU+h/L4ckedPS9veJ
K0L9eo6ZuuntcylirY21I3McjBRxq+6K4pElDBdCdZCVv21U2k0b/Mrn2cYJIAQ0HCTwnDJPNLXp
8Dn8OFamUPmvjIArpQ8GivnryqeSfPXtSOK594zmo5gLTELz2oupt7bFwkZUtxx2ducu4/VyQAiC
SWBpJBh6tMyTQVAtGE84bDmzygAmchfhWfgX+bKnc9c510nBQl/TvmRuJtCuY06PpFiu+FutjtrB
X61Kv1vPid7MOmeTllzMjjkQj+thIYXZsfEG6RnrHSymqtp+dj792aVfU9xCO1cyQaDgvWP4Blk3
FUrt1drqgx+GsbXm9IR0Zrxg/Q0PZBKcYiRkCzg3UJ2ib+XDmQXJe6DaIOujh3ryO9rXyW8vdbTq
aSlQ1bEMtH3SivN6kbaNcNUH0YtJfXAN6HbRw3T+Y5/OGRN5qHw6qoCATtcfvoLSqYvNSnqMR8/B
9FBvJLiKGFqArVnPRG6kUw1Nfc1d8+seOvBXPUDrq/M8vjXPz2bQtL4VdJqRM1hjUvAr+/+/UiHi
uI6zK6TItGygUc3OTI0NHRsq5nJ8q96c1Gdb2I1ANVI+DRonos/2J9Z4Za5Hijh2ChNrFmwAHH1V
4a5l/HM/B4hPmyGGcH5Z38XR3PqGoyc0w+KlUk0Dql6NLlFtJLAuR1MZ5s2v2LcUC+0/6yMJGqE5
DLpAouFyCNKFuZN3Pnrcqc9FkmT3WUykECYnfTgSXGEQGu5rW/o87dB8RkkJSDRfHN9+i04kw3pw
dtAtwMN1rQZRPzsM/jy9vOP8ScWrTLrm3c2m1vuGNl2XR9f6Leo1FUN2XZRMFzZ1eXYHhOqtpiZW
C22i39lx2491bUBVOMOH8Lrp6iybx1JOTa+WQQZY0aRfREBjzaHYDYP/epb2QDg6FOZJ2sllgi0+
yrQi94A5v5FBzu3rVa24VX2iFvcBMFS39SlgnwqJiLH7lo7GLWcxy3maYLhKtTv/KePAuMdPsXjS
q+FNWRoumoLafzykDzSKnXP5ZUcverTcoBqwoxXNCHavp0Lw0BzAkHxtXuBBJKjeysEs2IYf4iLx
lvuXImbVXq4WA5/WmcABvvk11rDle/rg2c6uTkXdW1oitKyTZNBuYFgyo6hMtIBagiEZEiYiUptd
y8dFwrfOqa/Sk4+mmtvgYONpoQdhHafZTMPDUOEcu9y69tN748SjAbmGIWsTLEL95ZT5Uw7Ml4IX
FEO/M1GySwKz2fYPSJp1vx8kZG6E1WZSdiB87eVGgY/5KEgQ0BJPsMO9OpDbYeyVrJf1+Wc5z6mP
Q7VZ15Pg9SE+nFTlDh311QB7RnORRN0Hj8nUJx8BvmK/1o9KEGcQXMIrZypzOKTrfp+Dmt8NA/Tm
PWvA66goeD8WXAaBVypdAs5DaelfjVsPgFtaz6OOeZZVlP50w8c7DYbrdE5M750+BX3x6pTQvgm5
QXTnnVDKSWbv16iXXhFJidFInav/PdTzt9AaW//SBFsdT0fBzpkXsZ9NtLuqfMloYBawEMvtVKg1
vJ1sRwA7KbCtM+PBkxZ7B3cbPrQ20FlVoavMp3KcRHuxQjyvi1imIRyA1zPOVBVFB4r8Q7HrMwgR
zJ+Dl6B/a8hWbA8WuyAX0BYH5f42peCoZRJUZuPENN5ZwgU6ywq5125jiXrQcApxtvj98nKQ+4y3
AmYu/CIBMXy7LtlYc2zRQc/4CD48kANS10aSheT1weiB9Nt1Oi2huyvV/eJ3DXCEdycUiYZCMBTK
fU6y1kY938JCzG7mqu5+GGzADWdgXyspRNv+MG+3VILaU/zBDEuzBSZO483al4RywDC4Av3wAphh
kMO578eIQiy2WW2MfM3WOgIk17USqqegPp1rZfnwKIZKPtqtHdUfRM96b3enKxIXk7i9sT2xlcSM
vw8FVXgfGXpwjxQauPHPB2AV+wvx/S07RNFeGWUqCY7s8JK9RuPgGtNCm0oasChFf5gEZp/jHn85
+SINs/PtiGRNZlbUTYzt4fwXlP3Z0JDWJeMGQ3feZSjj18XIlbQMsM0iFiAoHmOzy2hVz4f9oAGh
XwlaOe5skqMwmqR4MOyO4EIGarRheZsB+fKaTYRnmu44CAM4xTspriCVpUtTXg99hqS1nhjpxYXi
vehbRmgD6uMbOT/W+kQVKGvOeBftHowRqJD/WgYLEWS8/pXdG5sZBS9gASvL9igwzAPdhA1XQ8LJ
ACOLCMiLMPPUh/6BowzTCr6LSV5b/usaM50Iaez1iBZgV+KEJ3L67eTMCcEre+qyyVZphjqqXMnI
7y8MfA9q1yHUtb6E4cpG2qZhfZOlwINnhaIy3hyGv3Z3zyIs5EJzeg7Vu15wBPT/nQzskFI2MJS1
bZ1RhXqwU6XSKwAqN5A5ZMrYSHES7yax//Op8bQwwtJXfR1efsCennYPl1oMS2uRg1nzDu5soJyv
wnz0d7JvLJjmiu2TE8LE6RMvuzO1IiiFhfFiuD2D/8XnBETV6RPsuLijFLyA4rWdoKo8rdPu6VpA
Dk0UDc4UDD5eBPnob4/nlhbVO4FB+KHDryteEHhOZLBp0DnTzSgfRPI62c39L/pcLTk3vvBB4f7P
2kE26CPJot2SI/L5XR5E2Of6Cj9lQuUY8sEl8z3Yo83OQxy5GaEqhwggSIh6/1LPDoKfb0vEWZhi
QkaFxkVAWcLxxtTHDAt9FZoSMi1+WJdHqmIcR60dyBhDeEBxUb6ipnW8hUfqNE5WlQxgexM5Phbb
CcLtOmipGL5L07vB2P5raVPbwRtmqkfl8Av7e8KQboZd83LKQ7pg1xorAPDGKJ5NCswh4B0Fhiwi
QykkMo2b0xc1oXUZPP2KSEb5uhhfHiaUEp7UH4hknONztWImhSlkTmzzeENjo3eJfaljqG+qatZE
NWKg/WRKOCB078Y/lIjQA2D74vQLHqYDD+hmEwI9GRKS0/jHJKusWYs2qIpdmk54nNLDiqNfY3h4
SwwkhSK0lcr9WSoBUflYKNjAc9LxZkbRs1G6i+q9JStWWXQxl+oBG9Qo4Kc7m0joZpX5/+nk03UP
FiPTg/1QZBHQU8YtNqGS8xzI7lfm4ALPpToRkGnaXq9TTOwS/qEyoFWTmx8BZTm67mfam1u4OayB
rAKA+lFBUiKPCfVB7htcdrG6fi8aW/HlRk0fya2PLHBWKeou8KVMIEYQ6OuxlTkrFiIV45gvhaUA
Awppn1kGcXJd9zFrvdEsijAQQNaM+cUt3GM2+O+IDEkEjGImvA6o41ysMUZx8ukaH6Ha90rcJWYd
1S1N+IdEhsHOazsB+gMNLr6meP0u1w66iXL+qg5sPyTv+lFLISLkZUtknMwWnKfRa0yHn49/QM18
Hd4/Rw3bGGAzXf9arS6u49JrLF/pPDHRZwcSEvQdywy3Tg5bCJF+ohI2rfE4wM2HCxcjMgagiaEn
WM1ItW57I83j8piPdluuFWUWQnS+wuKL66nTsRekVhA01lSJzPjIYnqWw1+jf909P+E/4Nv+Eh9U
ahmbTN1f6+P2mLaFwstOUlidm6K9W2AFJCtSEKSSoEuIvzHqoAUJpzeNf5pFReSYC7GiyE+25Dvo
/xJ5hZbpXyG1H/NB7C8V3797HkfGd6oV/FKIGsDi0LbeT9DlZcyU1/3iswXJGP0W+EC5FmSpR1Cw
Udni+D6eUKR+fxF7TN4arzsJM5aPDhC7o6w9aGB34+Pb1VR7xsa/u0xTzAd2BQuLJ6uTZXD4fDck
xEJVOxa/fWlAcwB6ZryFb/nSkQ+e3C40P32J8ci8p6/CWu/2QzBnMXWtOdFmuav5qVXP5BhdkZrW
ORGFYAi+0+x4oWgkyuKfyvmr6BhiJfiSJVMIwCUa4b4kSXXidPNkhiGY+v03LdMeDlk+tiBJck9g
lMKid0dsJpH34wVR+hcbAp8UMEohDiTejwX9kwQNLQBavVjHZKrjtHl2N8JcbF1iUdS0ZTDtuJXK
UYKNKqT2YDZcH2fxmcC29/3oyH1+1xd/msMtnf0dlNch4zpzP6SBsS9cqvVNcZA3Zb5A7k3RfAwU
6YMfKlqAL5jvd81PFLC3YdeYpqIbi5hLraBPn7vzDtfj9WufLyqRTr7mALjpaN31laukeUUJ0FCE
hQRWMda8IlihLMb6rasNDs+pD4R+/5DPIxH0lZaSzUhdJQDw5Th/1UmxjpQYB8wMlvEKsnjvAjpS
45OjOwOS01MXNYVsw7bzgiNO7KNQ7g1xA2OovJBM7oeo4gmn38LRWkULQmFsr4JfTG7YL8wmduB3
jxB8IBA9i6ZDbQ3uEdIwCRa3KTqeYzrbX7fHghqdHEx1p9qyUsj7LCdVlIPzKz9MzXF9eaILFo6e
8c93HjwGQYDyrhiE4olYLgyfxd1SVCeC07GKpOrtsOt3e1XBx0Zl+JT5MlRmvXeynjfkpxJFE6ia
jUTHUXWWFcL1N/XSQM/iR7RRYmJliuN4Fc7T3IrqKgIkufsxtnQfHUaqNYqMZFMwLiiW54FvwqNK
DgP3rsghGU6oUbH4bl5U/cFyYKxhV2jJQHS6z+3jjPNelbtEQeu5KDx+PU/p/N1dpjaZCMDr7xqZ
amPuUe7u9TvL+BWH+1q9/XGYpucc/rrOx5mIuhywDKy8GyKIq7rQFpl54DmZww4TuOOKV7U9I+9z
7Z5eevOkkvJfkDBMNZC2eRgnZ+ZrDvyZ1pEvXTC/TUCMfjHulEtW44MI175m5qsGcgXKJHXCCY6r
Mftgfn8uryo7M3mBdplMwlUt7Ol5lB7PyrWMIFsZGLxjA/zsqBiZfwED8x5gFbboAsAwDESGP4LE
3GW4a5GwE/ObJZumZxFTiWknUp5zWzDoGFP79dYPvnIRGPqZn/qoCMKbx1kZYcPW/OG0xafHuE6v
Z6PyIaEpvNwSGjRCm8JC5xkoSYcx3Z5chgLz6jv6w9Pfxrgpi/4Jd3rclXiDZOuRNS9OmFNYv5Xa
PfFj9AI6hZ9aqGQ/P+meGIFk42nK6YdeMbDUTjqOCWGfs87ve7O5qjsWsf6MvS0Xxx9S7178bgbu
5yiw9zoamXbnoYdobFWczcuMejS2vhi6S+a/PODfctyFAU7TFb6RKtU9WUwuQsNrcXMsoW+3wwgy
D1AJ52QX/qI0TkSIv+gc+Oup8/AYJU4o190MQQL2cnRE2MWjwnpFa61AyVERs6UI/Jhs/rm4zKs7
4A/5J3XerAepqeriZ48Wn4cwNsgp9rNEekx7RwYChb3l8iDp1FWtO4+IGiwbQ+s6XTx1PrJvFEEB
QuxAhG6BZHN1iTUNqSBjJunpYpn+v3cdxJjHsI3nBseJrxiJ8oSl1hTu3PJBES1en8Cxa90oO7bY
EXnnHgXfmIPFIhmBOWLvdBNJgfio5ljJG6uz/6gifNf+H+AoiUfHhVQMWlentRUXOT3GwPQO36XX
Z5P/9XBepBPoZYSa4CsLM2BeNftxDugSohtFAzmDjCn9sfCLiqTIUt0BXJGwKjx/zj6dEju0IuV0
ov6CnKib6xO0CfWFntYr4C52tl5IBEVd2GJJG+uLPHL9g7a6OXBpFYo5F2d7Dy2lfzkBranuXxNI
MpmABVr5oAZdwuB7ofGSBD9Mv9mRjHAaZwag/5cBuwZEmoItxZKl2CnFPESRFoFY6s8nz3zovS3/
04Qqn6fYnmMc3w8Je2jRt7IFZU5rSwgUBHeI9KTzp0tbaA4pxzkSVLaLav6ueDV1dkvSvfunYsFc
bN4pW03B9CYOiUCtPbkcwkuVumzcli70q1+mb714/4Fq2T1igURN1fuvlM5nXpX5CzBctSmnkqH+
i7P1Y4bbCVk9iYOlURSMmMe9Ac6SrRXEPFaxoJDfBodolBKklPr/uytyfwZ7bWNrR0CPduy148s4
POE2qp3VcEb8GmKwCpUPz+F2B+cSt0iuUJywwPKsgpNle0nqR/e6D+AN0M6G0b2vu0C4VUJzdf9A
EqXSM/RlqD3dZrtJDMWSqkSJ6h1UlTb1rtVlBs6pMwEVLfwcdeWpV4aeBUpgpIN3S7N/CGKWqz+E
RwHGmbroNvxHVlGqfA56IsXGMMf5pRmXndBxsw7GR7WbRNA8CLjW355On1+qf1Nxc/H+6iRLhvvm
H0sXnnBVksVQTVSZAQH18uNIn3P/nMgNaHn86QC5n1FlIMeuG+nsklDZdDTv3E+LCwl4cpI87ob7
kexcoAC2z6i3QHKVegpNuHVg4sEHPoGXZ4boUmpBAeqeP4zWH9TbTivwxiAhahb+BrnnPYkfhCQU
sdgGh7+EV0mX7V2V/HmwckXqafCyzgK64uGwLQKaPHg/mjpZiPYICC0VdkbLVWjIc3WiIkgZznQY
xSag9BPtcQRCTtzbMLqb9tynYNqtrUA6ehXKd7V/76/v6Z5ZpCaBcSN0aUcoXKC2/x47DMwOk9Ol
EPL+kxndLopZvYwftkD41VppnuEgqFXAiVSuAiiwzJgDeBxAUBW9yiWb1leVRXeq5Pa4Art+1hFB
DEHgNCLBewUnbTymDnfb7+moKnSZ1sqY+Qo/gC5F4ZoZ3N+lmvYQncNHPQIRwTwgN5fQyhOL6TsJ
ng4pRBh6+2QRPxaVcFB4xpHgTUakAGJBhHq1jV3B6dneeJ3gs5etULxFGJIgw3WsWFvmFW/QMIhw
OlUMRtx9tRLrKWU1Y9EW8ouKD+pHC3mTLWSwcy3SOqoNpCTMFqLINT78wtfQS9zkRjYN4GYNRPWJ
5v7w694K5/d1lmBlOGAu2WbY+a64T47+0CpxQA0WINQxmE14pIt/ATNdbIrwydOkwIs3jvcoGYCI
nKmv+OwqTB0YgtE5x6K7cfDaYYmVdGb4zL4SJVdeYMgVPoS3dUWIXFwDt6/DPBU9THLZdh21iFPo
LwRmmBbWYimC36xajoGcE4jK/M6Ik7ROru1p6D/NBdYUwQjOg2JD3Eu/EahwuUqy/sTNwdQR7NxP
6u0KWocZRvd+pAaanPyjSTwmVxQUxHaxPHu/mzk9JqUchWODqYOP34JboO9GrzEYt3NLjoWQkEGu
gZuSSpGKvSwDOfzd/CwznfEnSmYfQ+BFm+NleH4AZRgdb1fhDEw2LGKuRYdT3FuMyJLYpleAcKbH
jxqtjfJ2OLznYG9w9ET0riMcqHkc6PA1a2wSwXydBo/+SUi0y15xW0mewJQnG9E9luIrmPWs8r8Q
W7YMfN2z6NwS1+jCxdPAdvJkLyCt8sRLbnLgSCb7
`protect end_protected

