

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CmScm1EG7+yOvSHJHM5cOhdqnLzZOcepWxY9DkMOyN4kLbgbdLuAH/l5P4gSPyg81gBN3kT+DB4u
PBXNo4263w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fwqNpFcMm3h5oYp0iLLBA7jw3Gfbtf9OYXqaNYQK5M/u6ozJ7zqm8z/7Gi9eaTLXS/9fpHpwK0LS
QxC2diEfybnFW6aKTP/iU4AM0T8Jfwg1fYYXa19VRgeHNuXnOnQbGrbwOzyL+M1AE6VgNshYAcke
HFUgdv42HBSaLBuVCGQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D3xIUFHSYN/tuU6xykyZi+w6uytCi8PG1RRIohuMCP7mdmezS82HpITZGe26wOIBAYGliyfJF+bm
//Xu42+HAg7awD4lB8/Gfse7Vws0SwmUepHhRYxtuQx+Hau6aq1uL1eE+GMEUXgxZ2vOXH0ipYrS
hLEg3TtjTbccTVimoRhbMQB8xVTXKgd1xaluMo7+0fNF3EBfFdhrX7VNbbmxpV636ALP/wC6VRmP
XNe5xXQjiv3FP3uE/Bt2VYm+z78C9QX2joRNZHnjI1wlv+JUs+OBnQx0uieg97dZpGTJDWS/ROJD
yUMDQnx8oeo5Aftp86QvBAbfaqE5X6J2q/lamw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WD1VRz/pLvBXDYk7fWsqqk9E+EKCxbcP63KaJV1ph2old7nkwo7SBQkXHtT+4KqXUeTJT6DxPa8j
tS5RCAcDnWldx37xHa9SUujjT7DruuKAJejsjhxtSfv6A/nEW4C6nOkCH10rAuqtBTv7SUZEElTR
EXiyr/yJfBZig+juuEc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TO3nxTWXykAydBE8oLE1lWHpTk01Db/e9HeGVQPfEOiTpRxWensjccZLTO1P6wLTocrobkWdnzeG
BxBt7prIiPwnDDfhHMe/xea/ckp4CqeBr0GVOckjbocHEF60X3dEzewbdNfFWYT0uATcWRkKB+5o
X3VNEsL1+rzFW3yXd3oxwxLZl2hrAEzHGv2AAZZgDP43u0eLOoQsuloFBUh5XzvTCc38IZkfTB7l
fBrAnLiMxoJyYNeps3ny9evx3MIX3RbK+6dmn9Aviq++SNxcoN8Y4/1btHsL6F9ez079jTeANSEU
ZvBBfKlGq2n/FXU3NGHAnGxirPn//Y4kyfC2Kg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10960)
`protect data_block
zA8mi6PWRxog6/ljI/G5/EJYHK7Wgy1um0hQTjlwtzWjOo1Lz6ghSt+4TNIdixdCGHFjMTmbi9TK
UcNPbRtnKIlLyzPowH0UTf3hDXf+PxHfd1rvS5SHjPyL2OnU5br9XTgvpSPcfwjZ8/Ml6dnDvh12
ENoNmajMIVu2dk2tCOTp75LdcgxLOa2pABRUkfB8vJdMvNQRzkRmXgwb0ccgaMebOvhELzB/VXrG
jr4ghY3gvGlSYblfoveuLUO9NWrXPxMJtUM9lQgXwDMfKi0eh5QGW2COFilyILJglkEEl9wwhTpA
MPWpb7Kfuzl+eSEk8rNgePRZH9Ji+Rk0aFT1mJ50xG5Xw8KXyr6Vq4z9urF4t69ly2cSbdgq4UuI
6Wubau/TvewvpxaAM8+Y09rJ9KY9CuP7C2FYEVDmIKUobI3JBr/j0MyJYfuQ4rMXff1TlzPgbfFc
jFfcm1XEvUuWR3hsjcGPdo/SYmLV96Pz1TlzggZ5RvaMsThhTUtHOsB4jL8g4a9tMN6wojqqULhB
Gc8dPiSia/6JXXEX0N0iUTEHCf4pJKRQE6L7dAOBmggAy6aD7gFttL9BwkpWt2TkCmXTltL1UJNe
PiG6umpfadfVUKtD3mtNFplqPtDkGA6yc0YdGOvAV5XTgzS1ZBKZq9XqCI7Xu4wcdAyWmk4Pj61u
2WXU9Hw9C50oaxR15OT++61lKTrjn91b9+ge/MUhJwAa0f4mpmkCm4V55SI6DFE0utl/eWNX1L89
ka4k05kb1pwPSaFtCe2zdNbFHPgMC4V6H1kNGrFqfX3R923zzGVRAYaQ2XU77SNOI4sg2xQiHtfe
sAx6jN6wL8lXBh2aw+EzNO2io7Q53qu0kybJKJNZFrMiriVMVQ6W400JkrCg5HvjdBNttP7yxGQw
1AkiCiNSlakHAqt53GxwlPScL+xunjjyXjhNEnIrQbcnFNj1QO9kYNNxgoOiMKdv9/hbhKm4P5T+
2i+xH0GPOipcWu2NpOjGKpl5J7FWqLsH+t9tFOdgAVZAYPg8zQXqQJqaA4+4c93cMHGZ31vbwJ37
stgwrKpRN+xjr8IYeDOn83aC6R6VOXJ3xmNdEPB4rOFYudDe/s7+ybnutrRq0vnZ08Bk8ep9Pciy
2OWo6c8GIl/o9MUJtHMQFhHxLMzsjPpzfjgSvjH9LOY91KrqlS6OB0cZCd5qVf09i0vVVfLbtmYC
EKLzncw8N2bVhIPTlJI1cQbK//w6H3m0EdCK5iIFIBwfN9uFA0+0E8KtEvmJGR1r42TPYDXduGuv
KjuPgrqQc3RbPb09+W0r1RhehJ8aA1guMDRFk729RknDZyiThe9zMqkofDXHhKTxamcazxBIjkYM
RDfQ5iVFLA6dM2tUMK93mAdBp0qJySoONeNsYRBLigzeuAVQDuXiThU1R82KQcGx+0z+it/dQlA6
vMDIkrwcVxgXd7j8WfsPG/1cXvnIoms82NRJVQP7oV+cj5Vk9+s8XGNsd3IGomaH+7V7D+OujXv6
iaASX89PsRwgS5hnK6mnz/sNqkv5bKyAgoCRCYP+96+FmJwU0rRJsrxnO1kCgJHJxygHDBCf55iY
VEhOATg7HHhKYBM/ALTWKYMaWcBctBBzXUDDoDUlGlPgtF9YZ7czGtI+aBiwhAd9ZfA1hn00h1fU
+rmQ6a7oYLEdXb90VUxf8jPZPjBFR1JrwPo3DzoOIlAtzll92SnE0UF0cIZzqIwKECs42sF2+mNK
5fKdBElmRlnBH1JuppwwKrk5IL8EjN4Fq6+bzZUoU0ZfE+EYL0HweDxKu8abgYwBAkGaiOGmd5NH
B/6RRZ3jcbhCcxFCX0IefdcqoqcN7S41gVoeyADBt13cFXTZiUr6AKmLhX0GQJeOOi1nNQLR4uxg
ZKH4vdSYTCQWhI5m/ZKdu54fxgUPArZ5cUA44uw5r0djRxqM76OpjJPtamxmtKh47nu8OVDVP7Rz
jzK1WOC9dFeidr10O3h3PTUETMr/T6ePavCNiQyW34+EUtM9yXMxQZ5qgDFN+GhTgM6+YzXfS4Xi
L+g/Y0pvGFlb+k1NdJjLHh67yprtAnWL+McdcsYUmONiBuZCPyeeRdW0Rj01SFHoJPrcKO6FG3zl
Z7qkO7IriFx1puCqf6vwXi0De/7YE/SrTrsXNtkWq9tAt/s1XafBh3qAuhQDadgsspyqBM12er1W
nvswogH6IyKkCzYOcdWAm7A/a1FD/8Zgbf9Y50Yp8xK1Ki8hYMNMQ/cZwfYscYis4g2GZ/83ewIM
g3zGhRL1jdnOfjCKEvR9LfGtWUD6sT7C19dVLnHA3TvctmBQKtDFfsvnpeLWweJrpG7Zsh2CKq93
ikfU7R/Zrj1deyYeRRMKmDpOZe32NuycEzUT/jEzSk6GfNqfHfxLbjDK9AdsZQaAsB/Ae/s90gkD
w7Sg11LlA/Cvw38tXvvwdx4ppg7/ujIsP3ybX8waKoNFYAxE363PTX560t4zPPY/UUVwtQIY0y0T
ySZNUtLM8M5X8vW22265pHy/hrOvHoShNa/35V7LrglWHbE7ey2ETSnmETOLCXg7tBnckVYr9nTY
0rpzwklaRNdgSpsC+UqAeozaSFPEPbwGAVS98QxMTc4eE6SsVsUB+zKVkO4iB0rBu/3PsLgyQBAO
TJk9UW2MivRutbNsMymPzJ+1u3ypGSMCzqvdLFd33arDggwQdnQoABRziHpZFyGKND4lxIssgcBT
CXpcPKOG5rtjSwEzgbuWncxbrSpaab/hBisMrEfu9yRR6xybkKblrarA+csyJCuxQdwg5xLyWA2m
4MEAD2WkCJECCW0ChVHG2Xn9N6SMGGh+ZAOw+MLbjxvcY4OslbuaqDptQlEF0rnKhL/qCTXT8dt1
K4r4TZP0FNU1akQ1uVJP+C3TVat9RUuTK/eC8AUL2kaLX4iXC/wJyVFFSB/ZkM8WCBFaK9RpqtC7
fu/3Qo3kE43bs5MUV3Br7k+8qmxAzxLZbBV6bVYfbkUsTSaWMTOxsIe9AQJfRA3sf7CTpX7p9L/u
C8IJrPvwY+1nhbc+rHTLYpw93SnjiARxJHQSQ/kQG8SCWfY9tW/RjeOPr8XbnqXj1NlXX2n8bdFW
29cwry9SuruqxLSPMf4ikf/jv2GL7etDvJUnsLnFeRvpo8GdC80U/nowdoaFkL7PFQ7l5/Iq73lR
hR8SIRACEyX0Wf9yL0ddeAV6eOBf7fMXrVB2yyl0Q4z+vABD1m4SffP5QoYcKHm8WPRlhr+SmMas
7brJRXDnNp4ojLM+RYDsCVeOJ3rJ6H5Ihbriy5vxBrOsUb6aERZA8FUTQULOVvEIu06ET9tOcQUn
S6PmBHTl1ZNAFKKBAnFQj7sS0dL1BW2A/eL46CtD5smqBaorf467/pfb9wtwuYH0YDc7RlGrounf
Ua11hNFfPwfgZYdUykRKGTYZ6tKfsW9zyGBAEJy4qQIDtoPPVljFPEVqGgKPvOQRqfjbha5JPrh9
jnvBh6QaIoEc6sKrqqUKSrwdRfK6vIAfXwgmZCMAsp0d2HQcACUFdIUm4KcR5MyT7YYrgoBjsCOU
RybhdA8w5JZBq29IGWR+BOVZnTyoVPWZVxq10if8FkXkAxnNBdXvfuCYDblTgQr3aK22217pSNi+
z3I8fffW6Ec50ugtbS7rN9MvDKfvkO0EgvpEYsUhbWm61xFBgKJbWwzFkjpvEinxPjsHVj0YxnyV
DrZkts95cmKQfcQekpbnmAvBlKvQJjkB/Tqypb39u3CImFj+JfWGIddknBC01lZBnsHiLuSc+cjH
V1NCSeCN1sLkfbnVmamALcRHKWVQQVkPlagknBFza/yvHK7xTkp0hGnaxScXWDqpMc72Eba/guaT
7Msl965I615gvistyiuN3mnaIHS5VxBIykuAU4NqsXVCvGECD+T/8Ycw2Vse3n3Jtpj4/SqYLE+t
k7xQw2KSnTP5dxXM6wXibLC5DGqheFb4NtLUGazHiT+HlvW3H0DKw3kqQwGwCLNP/Q1K65AymctY
eomdq9mCcawXNH8Je75OleXlN+IwIYxdRGfw/98oVAHrKSOn9HAR/bk/TXnSv0Ou/aWJ2BUjJbg9
FciG8zFiZfw/4tVaYDxzWxk3aM7uuRCNFNGVAHDVBl9Kn4VorxFLtPfkXmLBOaUS1bfO5PJr/Z8F
kOeTVW0ic3fIOD/LT/nnMpX1brrNCG1rR8bt6fGSDC1R5t+dwmoLrhgDmLXa8xF238058lbuqIjd
l7PaDgLvzJwd154KdwStIBUlt5x0qafZPHt9QJoxr8B+WxI/J9+fT4qr9CfqVoPRuA7av+wWdVLv
3QEoPV/E2Gsbii6OBJR90qE9uH3ZaBePcrCQ2J+D4ir4bKjAgDyFbQF4x9RLYrRDflwn4ud+x2zT
OoknAMO1MTmaYsRDP9j8yn6e1DaWDNQyAQvpwyEDGK5cnyYwvz3cAUKmy7y6RDKqVljL7Pp5NnQ3
mTpUjQ7arsr0YyAbPiHEyr4y4J9YQlK0hVz8ZOyJ6ykQCUEHI0tXe18kUeM1sjGar8G6CXkddSpL
5NJEb9gr9UD49K8g2TStG9Bp6/NByuso5uicL6Zguakq9Nmh5QJutUzE/RgYqmoPHhuru8L3uait
sqBvnoo3L3Km8BujU2UsFms7rLTJD8JWVz1++d8G+d/ANbL/56lk+oCZ7CUNjA56BPG0d8lLs8Ex
WRexjoggbnLmfkkiNxZ5APPC1IWK5uAWt70S5zGnt4i8eMcp8Q+hW5hnA6LbvwztBd9YR0yGhqhk
0tTM+lQuNFQcOg8ozgHJ74+hM8hNY340HoBdmHwI/Jzq2MVxVdchgkMVVK7Qj6bcsIcOPndQxDhr
iAYC/Iq/+CydCS4FCcE9G6+pjyJ4nc6pqbePFPU4oFLinUePyPgwhJsM1gv3US1IhW10bTvbUJyk
pvnBUP0goq/TfN+lnDGx8C6QExC1xfl5OpiicxLqdY33ljW5VaLQT2F4naeRd1cA7cDwnqg7u3iA
00fiGBxGWDQWXPQwhIUPR8bPtoKR8ZQO6AKo1uv/Nnq2hwOfi25vAflxWKMqPistLn65Vf9e7Rzw
klfWctB0S3Yc+gy4Lgd3COTofj/DXIrGQlwCSYADeDpiHKh24ZRqmIiEG4te6GXiAVLjRSBOb1fj
B17F5IMbCL/QY1odvIeDuPWuy1EsVSUdDKJ728nXw4SBcxUmSlb1oJIzuHF7w5UGfnhwPf1eOjM/
x+qlWEWv3oXA5cH+vO7F6rYP1BwEbLu1mRj92DimzBUwPE5rz5BZd6c9egBg275f+2ZFzZtI3MU4
qA1MOjeJAmaq8nGuMtFa1AB0G2kUi9MY9ZNlCy2D2UPi4dCIgH0mYPJHZcDc36orkowx1BaugCfI
y3skuOaqX+5pq3ZxX4NQ89zwIkY2XHgHBBeETDYttw54stJ3Dl8Q7Wb2tqBUTZZ8szCYfFpm9IJI
6E5pFcZcmEMzBwOmG+/SQGEAvs3S6pX379D+uFSEYnWB6cEuwgkE3bTejcGTFiT3r2btGOwNTiWW
wQ25utryRlyjMHw4rJvL056Xc1pNMxC2GXUYLCygXW+sm7JPqOgl5zRBGuW8irSMO7uaeMkrCSak
5UdVQX4QMsI5Vn8DdGX+IrRZLwBDCATjCaT+OKPpYGV/yi/qjmP9vBsz6F9Ao8Ku4RvaP0iRYMUp
Wb6782A6xyfUSjY4ZoHz5dDJMeo7uu6TO1TURKTuLrg53QBNojzW72aaJ4N5l7XFV4tT0y3mZQ1U
T7b3IIf85HAV6WOO5JtWwfdAfjhXp7vF3ahTp5b6K1HqhirONgpYhTS2L2z6LFNZy/853FWBOta7
0HFRVHOg7QM8abXYbeud/k+ZbmRQ+maj5edIIFaWq9g23Y84t3/sCxDXVk/N7y+fdN5VM4yCYP0G
r3jHWpFOqjhnO3vL61wpy1J9q1L+AJYUQUkJmtlNJVSvl1Gjtz9irI2b3YLh/clRq4cgu5uQdjap
tgUcT7YrvXFVbq6Z1r5pdf52rZBa+/XPLr5lsLRk2D9C+kFGqAA+jioJd2Lj4OqPmxQ+jOYTiv8y
54gKgV5miOga8sjPTv2rFKtFRz71EARaPvj58ixsdNFD54J/nW1S5jTe6q/vvdMfmYeG+M6LAirK
fP3aMOsCKJfg3oi0BPIzIodhk2k/MfQgGSmxtpY6n3t9nRWvT62Bzp1NQVqEmtKbVtb1M7rQlvbx
pGjo/cFiEVUVMqUSsb4wNXKR2g33zor4Ulax6RC5cEOQQsGDoDZy1yRP72Uqm61wUeDpKl60t5Fn
NqwotmgGRxYCszTEPpQEXKO8gVPr9QFT7yNE9IksePBBuFZ91vOxnjbTfzqeAL0G2XTjZSdU8DDt
zjX0VsKGoye2zK6GrzoyiemUC7xDuPlYpJPraFTv81Cqm8oy6lxVXbRqD4VYaFx38g6v0qDHLD/w
q9NwWFj62OHGojxaOqhvepa879JiRJhtYQTnVfJ+fkrUNI83LEPBB6t+APWizfIl2xeUOqwDempe
o+sgmlZhvOcReq/KRwJA9M6sIXgI4jKKLaqXr5j9m7taK4OqydBZwaZSdpIBzRNvL8NnRbnMuFH2
Cg1qxL20RMUGqqDuwXGLf4GccMYSEhSg5UJk/quNcq+DF8xaxjiiQzxwoVlfuxWu/TG4Pq7wLdTP
OMV61zj3Py7q10hFevVVtqAWj4NcJgCwZ35v/szTFix3fP7eOeM0qmM9PR4SiHQvr1I69NxFi24c
Y9GuooqYE2OXcJoq//rE3YELlRAtnVJGSa/YZc6cTFL38O0UmT78PzrbabM53RRHcFgyuqNlZh9k
Fy+1pT67N/XapgLF81uYvQJktJ9iB1XfhvaDHLiddgFYS7Mj9KAe4w552phi97sojNGqJTmLmN/S
5oy3NkcwUeQRoYBgJmNzKC4PopcrFiBTv//7kxWRxpMB/4c+8CCzHqT10iJnSzzAWqVwRLznfMDT
v+VVv8jtnmwadQR3cOFIR+P8wuCq3Dv/Y3mIu9XXAnowEjygb7tqclv8eRzjdBQu5+YVZgqrF3v8
t6qpfNiKCslbsR+cJAoZG9HGfxPfreRZGCj9Va0Ys1KWkLhO+h30QIZNr26Z5hKx6nOlxpUnJfNH
VcYicvfWGkoDsw+9TFjuopeTAkWIIS9m30ZmSdi+YP6yboptSEo1nzPj3Y/HBRnRFKoQ4jpHeG5A
lKx1VG0hmuVT++UKCd8M5EqxJvh4KcpUBhYF9V9PeWalcAdzoIN5OyGozlu+WyKFS9RZsah+fYyq
ihzToVQwjnfCaChUS5FMOV5dT7NeT8jen4Uadkhw31wKn5GjWvRLaz06Yg0PbWmh0y1ynoMVlg7y
Z+BGrblFmn0hdRTzVTS+LkDLhEc8R0s7qRJKw8Xf1ik+OhE5Z+9hj62UbXFEMfJV8JN7t7zIdy+M
wEe07sdDJWP7t6GtO1fNPO/mQGw+DRRqKazKV2lAV2IqN6tUTcedD1bgR6HCGaDHDkPFjk4VqlA9
/CNlsBkpWRhTHhYAHgQoG14XRHHCxIDi5JymoDdC1fdWsN6rXjI2VAVjrhImwEHM/2a1MHb4naYG
jV6HrkrSJBTWWPMbo5MLSvlbn00R9LhKmcMMt4mLVClg4UPViciapghBRyjL9U5UAm7nKzeiAbwq
GyHFy6+BDJd7SH0L4FlECf9uFgACs+ykHVUlBp0b85wFewhaookrq9CVvI+ifd87h0YF9HTFrb07
Tc2GD7RzoT+HvEsVRk1wokZqm58pvbF/A3CMqfX9gfmpyVzC/PbcLc5GhVKXyAQskrCXgRYQxXXn
e+IfaFWFcQEY0h+i5pYmCCHblTfv2sH82mT8MS9ccTnCQCRPZkb8bC9AVFoeffOm79HyoAw2g/yw
Db8SJzNTIRwOTksEyHEMb3m6oFC9hMMjYZPySUEeW3tgL8Og/XllGJ7QkA2S8MTzTTrc1I+UfNgq
f6ZWzb4N/rYVG+BEaZAfqGuZDEVz3IEGzfJdhvgxOR2PJt1U9/26ngp/crejkeCHYIXL3Q2DPbGp
Wgw4TUlIdlsDch/z85noZJ1qhqJhoB0Stm3tq5DdMyk7kWBuH4IYLYiVAn+qlO4usqpfzbLOvHk+
ENczHV64TpBRwXhhaLWOX6n5YGczje/Re4VEiS/3Cu5uPoQdEipVsfEiWl+AV2/Be5G9zWLTBVlm
hxxPtcZjekyuAJMDx7Y1sU0BXqKFr9EN51zvmurqg5oz12evD7zHHFpY9nSyhMpEfHVROB17ag49
WtdwOVzbnyWJw59WoVSl010t6g4uL3oAS3N5yAYdTngWO4TsDjJuLopnnFrbjUwOLE7GND2u8hDy
awKsA7jqfds/SJEFtybBBVvV/yydhClrOdzC2x1KM5nOdyi+6uGdSSYQvP+etyCTLIsTDnu5wmBJ
OGvvGL+tgkucE60QuhrnKgLv24fF0qs8t2vs6ZsT9g8LG8UeBuzfwLKJomeMyLZMhs+hU12ORkbb
X8Ddb+/VwouI8PUOjU1Fy0JEVzjpJBVA0L/wYqX8o7NGWX1fkSv+xNVfQYsQCwRGIKBf/qqvoOev
VEL+Yf+fpUdUBXZXxn98QLXvncKBmFeZbFGyfvTC3JlyJzkiEAlsIjsoH5KKVn4XkG/yxM6WwpSp
OUBNoVYfgBJ3kvSS3oPQ+QJ1dQcDREYco41USSNZxcp8ZVvo1hF6fhD8axFgrxBLm4UfeEHPC27a
Ap57lHGEUwJHCJDvX4fXp5I3TvnGIpp/PCQdEo94FYZHoTlEvFE7LDw2NXf24pdGl8BYua0cEng6
YHwvEdDWjYCzD6JViAAof10LJeYJe/zQiIpisulJ6kHCsD+4pV5gi7fDGMQM41xZAXRSqgSjAqHa
9tz6zUSbV/IE+0P0a3XHiY6GUKtMhAqsoZbimf3i9Rsz5+6AW/T3P2OA7f4WgQy+7HhQfOrEojR4
CflVrvaLbOdQqjFveQ6YhvtZztToUkxEklOLN4bHs0N2nBOpLWjKTTBLui3nL3P+KEmGbZXKCCif
CQ95zl4rfxG2CU9KBt1nqSGOw9s+Mnw/UCcbqful3vgtOq9QVc5rZ1qF21mwkXTpQC+KbxSeh/VC
H/lgrIg23jiMtgpGpt1qd31CpIzuvdyT4YpF2m4pyOUniihaCxEVDedfjlDPRhu/17ze9pJm/CAe
S47rb96le0CZXD/HqCMfdqaUGhnrBZXmQ0DHd8LEMwrn2pqrR7nXfmOQUR79e3FmTlNbAReMcUfY
JGYXRarDPa/M3ccLe9AAT4+yM+waIbN3kJsq3tzoZNUfNuwN5EF/7+dJG72LKxPmI3FNV2DC7L+F
z4g5qE8pSkfU80WXvEhNlKvs23/jbx2XtZeJ34hp2BpO+x8hjKnznmhlq5hS6kLKKKvFxTUUCuhk
KtcvqcOmIt5OjXk1UleqsWsKHEyAUHg7aKLUSvCOptp4t+U1VA+A2bI6o7D+jb59hJ6gELXTTazW
GZxvmoJicP1BcHLlx9AVKetqnOvh7ILG7e9hpLENQmYpYtZ7dGJnzeNJ3Cg44txVZnaejLkX8p9s
DF5/NA68Lglkk4cLRZzKxSB1sCddgexbmKWEPwVoESg6VsjoDesw/kW6Vns/xXB35wGEP4ciDolC
Eq4DWMUBgi+lc6IiCwAQZ2Jrhlg05qDtLVoIYUgWc5AJpt93N1M86Mb5wrR/zQCNS8Ir+R6JIA7k
/LFTbfN7hZecfNa0qq/6sXq5NS6HmJyJJQDqV0vOTIG2bLvkDqB7r9G/dJH6LOhpXOyLEDiLWwIh
wbyHqr05bc1a3LUfEwHm5lrPMT94FkFhuoI8LJ+emPI1EiAUjvumGxnsJL71mE7X1i4ropal8iS1
9yXr8y0oDKbdJMQ4a1trmyXQVQkEpbZ6RQjodGe0u4X6nwaALU4IbDaRpnY6viDYnuqwfORYo+Dk
hn6Ei7WiwpJGXUgUwyPHXZSZgs0o9xeWz+LXeM8E4GnkMpioFzgXlpE+q6ydfX9wsmPHrr0EVaSp
Kj4IodQgPX111m0rRUrfe2wJoI/WBCwWhe0FIROD4I/sFczR40g4+LmPo1LEZsRfvknBMQKlWOy9
n0a2Y9knxyWXNjA0BP5BBnn5B88vfRf5xZrDcwOVFa6aDT+x9kGhUFbyN6h7GyE1I4Y02jP0vujR
76VHZKG9QrGTAaSHdKmdl7HruwYah6wHWMARRAG5s7RL5Yv1qYmDifL2ROOEW1NHf5OcPy5Zws8r
quAvcEm44aVyNBvHznPobbHDKWfI1CvMHSkugVVjzraZAdy91X9yRgzcmDzi5KHW3TainvAG+EJj
p9Mt4EuZE/I/jRuuUCZ517RWnvlDCIITaUxqOYOG2TpheJJaNp4Gr5uA7b4zlS1qX3odqi5aNJKM
1wBZCCpz7W6AuuEwLEbVlvRy8QGxQalfMmopb0Zs3lFFwgy7TVjdWZ7Hnd9RYg21HSKphJOhx3Ia
+mVwh+oF2DbGtqndEue0hGJ8M8ZoT9OZsTiB5juv+Y8nf7Ol9LZLvx2f4jgL3PV34wykvEa/GlW9
4EBAGfVmjB+BNH9FxI22IDwJgICmgc2lNnr2Dkt7m0kXYTYuEA+YrNzAiH3oUxlNp12VPRPsxq3F
IkwugNl84abEqnyAemGw/bGANkPiyol0uJQ4rW+QpivJKXw/3jsFX3DaT9UW2fzUgFUaRScKNJji
RdjBFLRFa6XqZLJ0NBF7dOG0AscSaRNDA3nHcleh6HyH7aejoZCvamDYc+Y08ovPabQQqZUX+DaS
nREFD7z6GgKQDwzH1kLxriREz5Jvvx14HPCAf4Mb8n1F3yxc5CjSv5XtbLhQduKXnVxfWjbo+I3V
/J8X+44EvcUxi0NasIguJepJV0WQp8cVmT2kHv7+5qprTWpcNJZ0HD7eENV7TtaN/StagpmLjg/G
Hrkw4/od5fTayNSO6bGk5yFelY7mSCjIJzaa2RtH5Q7TbjhFKDle2Ofb6vn+MlGDisiz9Wgudkx+
+vMsnhDkIN0zc2mAxpuX6mSH/qJWS2FJOyyI8L6fZbAxRSK9VxQifSdqzaOze3IVdjPguUzMnsSW
GLofXd0nu7YtLEQCRmlojdsNzTo0+WH3uYc9JVEx8NuY/sZyFwOfejRpG2B8mM/WINl8JZrwORG9
nfaRvP+frkt0JdIpgiVKxUNRRPOGvaVf3Ajl21zGgoPLCyVyL7ZHUsRYzmZGzQRHU4DcX4o1bQFg
gEt0oEUat3mkw8o1jeNVzL5KMHBjHJeCM4o4L3OW+a6V5o/scqTowrASI7uXhEWj2nuAFHgI8LBs
htVvWUna81QkDUjKG7pOWTI3kqa6ujnpnwxzc2bZh3d9Ws+3Df8A0IMaUe5aex+51S4lEIMPoHMq
nTfRyDWpp3q23BCgnXsEAd9kzIA3NTH3W8y2FtToE6x1pRNr8OBoJv/ETKDzqqfdT3H7iBDJo0Xg
bXELKZtZkV6n6XHXxxXoXj+++xRAtEjaszeaShCebz2iZkWHu25jdH68gfP1wrn8dT+QAd1ZffcJ
S/cMfmtSYTyUCSSykOL0/UWjaAuN8oRrC9WZH2Wu6vY11Urks7H8/3iyWeDVXNiIIjoaEXc8Ns5W
ANdyOIGNXysT/GI4N2EcZDhYgNWnJen073lH2XOa7huy/4NP+nliUdXiZtgLZkyHzln7yloOf6oL
VG0KWKDXbATaRIlYbAebaflIObvELQmDy+oXTgEqvNZn34w6NeHtw82wRWz2jHUmJzsPp46oBfdl
MEWeHc1w4cwER5GcBIQhkFUzAI3om35S4r/S5fa9oN6EiJdE0TRBsFTuuyyIuQZ3/KpRsmf5R1Jr
Q/1VBLG6pYCMS+QSFTB50alMk17mnNkX8FC8g44SnFWbNmtKQNIT7CKon8P6Dgmggte1xJFpRC7/
+MAA2xtwJjuW5J7thHulyuJIrvXvGBM7y2aFhQhR4GCICAWgD3PFXnlavcIvJ4dXNwyvHk6Gb/4a
1S+tgROu0OHiDFy0EEWEPDFXgkZZYYqf33eSafq60cffTyVv6hCpNIQOnvIaBKQ3CCxGohGEiupo
ZlO8ksmnIkU9HqRu4TBnSBpFUk1ZUYZoUz2LN1OP7C2PoaZP2n3sR96XHVTX3Kk720M4yUQuwaPW
jil4NYkpjsCbH1JmS3uAeiX4hDjdyUYqi0kht9n7LWDPstVkaNXVR/T0bwENsA9cfMoZdPhfoOFM
1YUjMwrqBDv1AnJJvf4G1xgs4Pc+b7msiaN4AV541jBN2JqDJkhvH03QlyRdzujWgYiuvMhbQ5rJ
zIVRvXrl+SOl2cxk4/XToLFiYgYDqmRzGQ5jnHMbSjEZX915Ai2d3CMm7i5r936u4S4nzpGnyQVe
+CDLVH0+LZb4ve6J8AQOi/Br0a7asUhatSZTMBEd9V2aLTpNA1u2nJQywwKd6ipSKjS0Do4p6kRB
YKHPaG4UTW53kRFHuqyXRSOqeEQhN36YtX5xCtWwzmNi9P4IHhy8cbmCxzzlPul1K+Wo2vustmJV
fn3vUibr2JfOpYgZWXQaRBp/+fG5fH/QjK63SqqlFgG3+x5HCkBtbH9jeVUL8M/5WsMugBhlELKY
BlvLJsAPe1DjsY39GEQkd/IdlUgMAOuVCwo6v2aRehyfYid5HmMf6Rtehy+FIIukEgXW2A5B7Byp
T+uauh/AyNGgHtpoS8WTMEKUAQD0nlQWZnjArqdSOp1bFhwqeqNRKGwYSFHVwnqmo4jTSPDyegax
e29jHxi7LG2obRwLhe/i2HIqSZ0YqZPFLFaiexwBaCGN2fkamRAm+cdZ3QtyyXuP8ltX+qxLMezp
Rc3uprNxdxxQuw9ve8x1Yki39nDpJjG+9b6F+cYc5xbXjjFGc4sPd8YQP1rJfQ52kdIPPxUQIXTd
gE6aJy5Azst5U+xZP1PZx3iNHt+LNhbx6HztAlEPRvISaF4pm9YrHrbPjTqyNmZMPls4N3yZSS4k
RloOn6nLIHTIvJzCEU1O0wsN6ukrLqOAg4brHOxEvtVA/k7U7FWx2hzjDi7OkQ9Hu7BCDmTplWMY
BJ65/UYBDQXypVidGsyaMz4Igxtn7f3k6SjalfprBpOOb6qHluiidwPFJCK87BaCljQs0EgNkav0
5z4i0rfAyVc3OPlSKK9URmTpy+X4YA8ujV3cRxrYIslItB5RyAFRe39DEf8NpEkns2ysyvxwsjgn
NPjEU23gIjjIDI5RY//9UJEJ7kDTTGnpbO54QxMHOjedK/FGMY0J51hwX1XflbZUWlt4lUtufPfE
vkQEyKbZBA6PYYBNljRIRKJJ5uaz2KGIjUH6TE5lc2jIDULeynteVBzXMlY4Kj+UE1G50bG1blol
pU8kibbZ374NigqMl4ssoICnr2a0LZaOx20VYnyrgr1N9KdE3pJaA/ynWCgJ7tIM32I5jhoTf3Sk
b2V3cbVyzZuttTyxOHoar9CB8wduAVLlUszaeHqYSimPnivm/zMJZ+tbeoxIfx58MamQUgSG43Zx
whMLXigv2BFijoCI6JoFD+uXrJ76Vt4PNilLDF2OcDtNxP4kujWL3xLNujEcRlmxr0Tt+NcKpQo4
N4+WjfoHz13AJZjq7uRODGZnkgGN79yYglna/ZmMbRX+5w00I28+46hCxOmTGFK91OQtiw1Cy30Y
7MWn33w/0mneqBeqHd+MRco5ZkPRT3ts6CWoOIN8+NTrBRPSRpI7OcL2Dts9GEZqiPlgrEqn1Nj+
8Qmu2zEbzx05Icrn5QKEsPb6lyqCinBd5865Z/Wk2oRENPwy9+/3G4KT7lM3EmEvD4Yr2tqg732H
2DMb3iULBi+a+yOh7XQN/EyVfS63aEUBtkGm27qgrNHyvcauUAcgsUx287o4GnVeI7VPHmcnCAvL
8gWaXt3rJnLNi3/qkPurg0sdvTo9If5Iz0HuhJYcmAz2mXxx2PcY/vrLtH1KUsWvELvn685udJbj
04SXK3A7OGtx9c3fSn3ekCHqMUHccCakOmaS79nBIJp2hhvdPy5MyBbnRLQDoVhNCyy7JDOu1ST4
6Ky845w0CfheKARB7YplgLOpUEGKZrsqI5A+koE7iVaA6pG2H0P21gbxSaer1z6OGpLIFKMBaJTw
TgHa4HdXgLcS9rhPyk0SGxkzCqkJRTYSY2i/Kjlp8/I+Mb4F6UIIqpuYfrrNCLI7nX37z0S0PJyq
UyAZ070Ck/R5Fj3nSVqNLimihYYtJp7RuJADBi4k0SS0sd5KDA4+5FHQvx3w1rBn5InOirgHnDyt
fSJgIvTcousU9IYchz1zmImAxm3K6Q9ZWmqJ/NFKQS1fMuGdfntoO9CNm+FJAL5gap6G8U/x/iDH
oovmGHRCimp3FOisFpJVnNYEAu7ssagJlaAZgRpHFy3atU1+6s6Ach4mdC9QggTPciZcSwSCG2Xm
5BpV5orG2j6FXsHoxsPPrWPz9N5wHicvlnyEz8CICU1eO9+m8BMG5MJxOSSgDG2vFgWzDSEHDFaU
+Nl954RA0EFh6ur5GVql/V4tKO1dMfDOFS8kGAhOdFiWv9LVinSryibF0MC4znmUwPqSArrG8A94
9DtbunmzsZ9fw4pRzhwrog==
`protect end_protected

