

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cIiYfk3Xy6N5OP4pq3GmqGiiVNUZ6H5+UojetFJBvbKolIu21jc4BnJQVK6clVlXeOqxCwUuMeWy
2HOHrYFv+g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lIziGPDmnLk8lYYpZIaDaMbL8fBzq4Pr1Jhh0ulXet+pjCJLyV5jakxS1oSptZ+tHYCT5i9DwoXk
484l0YBwGxIV/F50kQ4mY5SmovR5v/32XWyGw8Sob1+z/rA/iYbfy53jpQjBFTMhONxMl2jPMKOr
8b4lWHN3CKPgzR7gpH0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
htRzDc7r6AHMWLJSZlCSE/9tAboPhTxPArTqmJzMnfBntgIxMOX2YAPT8iZ7gZlglNlT/Bmc3ZIa
nj4bYkmP/Ed/Ze8J5Af7OuS/hLPfbdPEIMVOJrAzPKtgRUGYzZFakpIpDVbTLnXVCXGbnWwhbHOl
N+MoLyC3ep/1xGkMFlPyLgKVegokAfOd/5ePZ6yal5L+KR1ET32v4t5eGaONowzpG0O9uY8LtLQU
iVJDGAf4BzpePmtzOyeo5v68FfUFTjm1d6csF3e9pbQ9fEwJazksjJfyX2XYuUZH1eu5bhyJMU/O
c9/o5sfORhKXoxNo0FDKepouEYzneEXI8uuD0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FHtFxX6m7YezwdeWAQ6jmWMHTTCQ3ATyb5990cCrfHVNkzUwGdq1shf9GRL+uR3C20sVQ7v4/+tb
aJQn0JjlSYvQTO2Q6FVyjXNHAr7wpM4t4p6I4KuMXkNXuNp6PVpERQgKViWQe974sEr/n8wacl6w
0ZeeyAlvAxPvOHeW8Sc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WrHRD4nLu8DRRwrUtiyMH2ZN6Vs3L2kgyFgp5P9DMlNKTdIDDQa1yTQPpciIt64OlniyoYCatBqg
Wt8N5KlawExwntwLmfujXap7EAFuw40uyJX+yki/gczIgekz/25Q1+NPVfIAzqSReCro4UUW45VQ
4oIxLBIF53PvEJm3CGD200yoSxIl9Szkkq1FCyNtIufy0im7xj9CnEg/iFEwxzn8s8Ge79lV+lhg
fO4H7eA/Qsx28fzoVv2RYnMwC/Ln7iTt2527VU0KjrPDX1WGbNCJ5ny6IM/daMbuTMvJb5fz48+S
KUNyOcNxuhu15WGxxGlN6mcj5zB0r8XxgsnOfQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25744)
`protect data_block
+PBj36KvH2O46PIxL9MBqeaMNwiG/xO+qczVaeMvfyI/ppzrf2kAFhAOUut2+mJu/Fp0a98JHcK6
yQI8Jbmsp5jyX5M/JoOu+4glArNVoPbs+NG43CydXj9wS3rLOf6/YGHfVB/Sn6xLGncBkHKynOUO
OaEIMqGEpfrfa4ZclNwyFxoX+3dFTWYyd/CjY8ypeM2OL4vxoiuVcKVDCpaWIiCyc8PFSKx8cN8Z
yE6yg5j7YnXNCmcekf8cpiZd6BYqX+cx5rxKWN0ssFAqoo+e8q8xzjDS1k3GszZfO81XuUczG/uw
fr1C0sEdoNQ+m24mN0URyQgruy8nWII3yHyIV2qPbukepGHs41C6Mqr1JMno0jmbmeOiJ6iAuHMh
hd0itbMplLoJRamVn5wBdr4jal7EExTRWzuvylpjSLNNuuy+RZ80KNO0Rd0lzlUC1lQ4xi0wvt3P
AmjsK3Wj5fNAZneP2HLyfqZr3DcJ1sWrDbXN7jsdH4lotrVJS27JLx6uIZ+4lV1/BcOqVuEghr/m
aOeQ0hzsBvBRnoETwMhqZoKN7WeZlnZWVXE7diRDDDczDCEQYam9mi1c78WohkL8QvIbWk2nEkFg
iIJykwgl0PABk5TIeJpfLnXIiz+6DiMl3fc7rQsTwZhD8rOg1afvSObsxIsCAYXMClg6/HIuE7JQ
wlVsz5fOU740UK9RIstxgW7MZUvQ9nnu4NA+/6H394gb++CGnZfK5EgPzTzpxvQcEqWzKxjXN5vL
nxRFvMe7u3KWAw38dBN84oEmeAUfJcezXncsD+SFIg8I/rNJ8PdtJ1f9ghmJMCwmqVEQcgV/WDHG
E3dAR0k6UqfhJ/kGYfTlQUGHzPhNyHTNe06wA54VHzVAMj/y3b59+DSi7iMQAyiaOqRZ6OMFm+9B
BZpHkvBWNuZlkr+RHmeLLvefWxgC53PovSJFjyWOow4x1q0MuftJIYagRnZKh4XWrhJkRDGAWqlf
YxiHk1NtfwHFsL5iixp98YeZh1YASn++NwhCQF6wlF1bSB0pN1nLaXTNONXVinpbN0FgP5W4mp/K
rjXzvlfHjR5zZZy4KzUQlsKP8Rx8InR8jXMNjbV7971Wu3hRTL9VqmlgTySWStX0GcgAzA/CHqKI
uuGMSkbnnWJ1zN6ntf3pa4YLRIM3RQaKGcKPLafPgIXHXyrUAev0mmmT86NsFIZ2l72kpZ+a/mbl
tsCigseRWfHXxmeOE0+Uly4pxVIt+vZnWAn1FjMUVX0Z7G6uvrj5T7zu+mBEsvgXxeeHStmzmETv
1tE6BhAOJdvBAkilJbQK2BsXT2nd7zcHx9UCIRb25vninQtVTGXCyelORMvepYGBBwtgmhnxTHwg
a9oaamvEm4uNGz9Yb1Qih+c1czejXHM7hxQB90wOo6GnidVCH2cw2ssopQRsy3AIiiUEdX5Jq56s
pAI8vWYsk9qZa3qNUy96hAHFtNzsiyWWMN5fjBet1hh3KBDn8vZPvKy9KmCB06KQJTt1A4UxHE+3
GSzGgEI9w1ihpdUUwTfsTKqDlSsyMHxSV+DfeHqOqUXrXDuggjkzh+HcpQKR/RgUhuA3ekVFfDdy
BPpNv4bp/+nlZRDXObDaVagxD8qZFS6kTAGRvSqUEss9AqHogPxfUZbA9HqzWj6GSlMG+D5YXiyC
C/xVjtWgFQmbas/k9eB3Ql2SoSPVqWbafvBSgHZDKWkYvU+YBY1UwrH9N6JCC9x+kZ9/9cUgklnE
bvYKlWjiLswZO/zNZ30Xanzp6ZW+KhchkB9licITBQ+55G26wsAk6BDigJXlq9n3aa+qRtZn45S5
6VqQDVHgsFQFEXejIl16+X35/qyg9tBG7T7K7Qg546rbKOcQAa8/zIOMt/1TUt8/CX+HJ2yUGDfW
Y5Ch2D1u1At6BBE8thtX1tQeAaMG4vROfnFQlT0/616V7y01WTakH9Tt45Ol2CzQynDdoYuGH0zU
Lok6eMUoWMw3tfcNNrh8E0tb2mVJSA0AqrTR9ZXyxj4qNtuzt7zoHvf2Gwzrtv1UHY4PhPJ6gXk4
OyNombFTEaN7o/pyC8ebh+G6XRx+N1OoXjFdJ+kvtfrscZzZt9TlZsVwIwmLiehgn0aYhS5GaktU
nxUUmT0Ic1GikL8Ogyb9G9nbSONr/9JzR6QowTlg+eX56V/9e1uzOc47UJXCr20jnj8jxwvJBThU
YxS+zcJNT2xksCIdumaSWpVNhrHgw1/eIDgorxgI73gvsJ526vja8WXACzpSzp4N0hpe7DuqrWk1
whmJPoyChFhHXSdNqiv7Dke2DGQmSTc8FhcbHYovH+9U8ejiFXuKMM0EbtaeisgJx6ABKfAhEFQ1
vAVCJWVMOtRMao7xvpQ3QXY7vkBOr7fF0TGi1Q3tlKseg9IdhVJ0Zx1r8XtN3/ao0pnWe/HdZjei
T4+dn8zMXi7OZ7oeM444qp2/nSUb+Tz4M+XNdxrnDdarZ356T0LUwXyNJAiEJjVZrNirypOt5dGG
Yh8auKiuD5jL5D0wL/S1eEOOQVaVMfJuYZe0gHoQrz81nvWhzvcPU2LSmgn7qJsdG4nZRFOLw3KW
/eXlZL/l6Pnl6EGHJ0uAE8jG5yzEe52U0/TXIiPKMFrx7scZdfvQxjISxaXfJ0v6p9eebol8Wq7y
LlLzxG1qPz+lM1R5AIUSsb6h1LnoE+D5URYmDz9aLtXoDAYi26cE4eciAxdXqoZNENQBlW1m3d0C
x9TFEAXdLMjHgEcMBefFaVIpeGzwQRJt4qrskZnQEz9Zq/rfA+M2vVPSYZHLFr9HpQUHmXAoVuzv
4vkthBKfLqxN0b4K8xvAplCFDqyV/kNAo10DZz+poAWCNslJBKXAOtzwnfF6zCn19LDC3AM31wng
VQd37r67ZziA+ZPpGd3c6sPR655l2T3eKS4ggZfYHIF6dmE9OL6D3c/S88eXI60DQPF5EVjgGq0H
emyFoRUaXsjruD2fxqqfsdteGW3B+0XZd4qefEOR6J9Dki7riKOdqX0cHKIytbTeN3cuEtSXdZK8
UKvKocv+T/EdfjxtEdNQin9RG+2PDdmMyNKBaGKxi5R4yYnhZQnURLHB2hUxBzfo5hesAUbHclKu
NSthQ1e+/11YYJIa4XXL9tKHsS3loQaNK9aHoavnWu/UaLIN2S8AlLPa76UyG62nD+wmF2Bef6KW
Wi6lGUNt5gPL96QLv0khDxG7GZSlb65IwbDvzwQcbgWCFghbM2Mxs2JzEg+fc6qyPUDSDfXMs1tQ
sg+u3svvROMWOpArjtu+hnrdOiGR7hwBitTh5CygOLZkdEc4vOeRV2hQ/JUiREDHirMAEhUFHSXJ
rjiw8tgObO3o/RRs/bbAAN99kiRrBi/EcJDw+BxhN4blOryqTl5Qvt4I5STeJ03MADX09ihMaEHE
aPTVKJoVsNnJ6jGy+F9MmTqh4FPafLK1Wmt469a+YZ5HfjdgjVFx+ligK7tMzApDw7NGXtY8kjWD
4gR7jbb6EikNsejPp5ZUDMFRfrWs14WUPY34uFi6d2e8MeElEAho9Zlfxkmxv70dCDhYSLppf6YB
Sqw0SFDDB4gU4C0sjFQSpMVZ/JhCWO8HKpxzpc/Afk6Q69cGz/mrnOyCiPhVaaLpwDsifxV77RLi
nEwmB3anY3SRQxhdpmWoOzN0ZM8bD93Ghn2EOYCiCqiqku1lXHNF2Ee2LvWI+s7WHLJgo/rlBWDD
i12kpYMMmiPxtk01iSOTCQ6fpj8B7DOB4ZXI/9uunfa5tSd84RmlbN+xpEsRSzpaKg/2tjM4WQXF
vQaO9eYh5S91u3x0z/mgFUrzVgN9Ds7fQ4Eyn7Hs9t/sPp5arZ71zcU3QwXkeUV6tqlwWNt1mhRt
XzDlU6zrxi07Ya708MMHUBS/50Sgf4awO+uyg1ZjvoPnBMSD0f5u/U8/uXm/BjJQWEuij3IamsFi
dgLOry32ZUtm7YIhdHT8nqeyRh5g5pUKn6DCtws6/hpGR2x1DK+bR3kATFo2io54zcTfJCnT733O
kDJGbIACDnuKl0rhl7ikeTXlhUX2Xv/XeE6hvhiI7fTPoy4UUeLLYa9rUEauUAJhqGdiF2sTpP94
F5+BmlyuxKJ9vE5V06Y8dnFXjMlqfqhY7qirnPkswMgAVuEszwzoiGhNmOOzaazpXbU6aHEYpVO1
Uvv5uo49e61F+B3rmVMhNTBpAYs96zeui2uhXY0x1wahg9Md7nmb9nENJbDjNOcDy+NmfUU3y1Ms
XS8HhLu7EuiVWkdPGTZJvGDq4aZTNialzJLzNIjqE99JM6WL/ybLDYTNrK7Oa/vs7iecwwkaYOez
qpabNg/pwy3tLyyL6tXLex5Umw6lQlgc6bhfQJMdhkQIRIpKCrbHSGSyr348s82TIMto0P31Um08
ze7eUhcYfsjjSXrWTY+VtRdY1wQdgorvLKY0IL5Y/IfoXSfg5475XgyzZfkWNr2F/OPCj8MgABgM
yCFjeTgmTTELhZjM4UUW76zmvCytRfVWchqIe1MO5gUSpuQpUcWLYUNmbRaLghQOTOvS9bSI9XuA
02+KziFDm8FwJ18qZvdm731TW/Yi070EvS9z2C2qKck/QAqF80XQVNIdBm/njaf33JTxt2YGmGGN
Wp7r9PWzvwwm53G84CHYHBBpUTgcT7U8ctf6OIGSG9GD+JhS/bZsSQinzysjwP9lLGK6ipltl7bm
+Y5+XKonhImy41LGbILnpUl/o6uose+P7fsz/o6LbsNvjrYfl9LiDUSOjTlyddtcd2G8TNndajLo
a/N/fgupUNIewRpXEOE5usUmw8TCPGNTKhhnPF1RLL9hej8ez8i5LjQfP/ni5gYmX7BFWnqkmfh8
DPKpjmQJoOC0wVseB+vYBUrgjNwJbk4nAvwOItKBFRDD/6nhvZh7zmJu7lUvXWI0p+yNoASkYPqt
P2dTnGMjMQkrTMDP9esk0fEp8LTzSW7wP9DEM1TP1owIIWBJJLad99SjMtT9qiZ931KjjEyfLa7x
ho5z+UBYH7/jkHpo37mOM0oPJlQv8xmKeCu1ZFYNusHTarYI1dqOtpkdQAouTPUaPknsOnnbfv9h
kDPR2vCdxAWUn1Uoz52MfPX9C8mGNnAWPQ5YfBjDThon5Ym8MhQV/lY1ilJOb0QNBweDLJ0q3Cw0
lvmMwx1WINbjURNiMllOvNxvpIeS3HBK2+5DRkOBM991+x3tx4TqMAqS7Nax1kPHCKkSpmRnwJQn
Hzbfje4X+PZcQvsEUZ9gR696njuxaz146bgJOeMRz8fNpMipC7U11nfbkxvvin4DiANsXur6Ma61
Lt4bC8fSUxq/aED0i5/FwzpSD8Zn/mGhRKlHsKM+yZYMN1kftWyqbgF1VxuSC/UlY6/Q44Xowmyo
zIT6nZH5OQfReVfXCsD3/bj2JIADc2R2Tb81mdJfYUs2Yp/LghNn7083G4KAV1b+1KXr/KEkS1xB
WrBqX8uHCW8L5lFWHGMLY40kxTCuPXyDaMOo/DEyvhmYy5hEd6Y8LCT3gdSly7OAvDbozfGw8M5H
Qel2Bn9dcJ/h8RyH2guB2DZJGhTnSSH4yrRdriP+FIcypQMMW7658mb6HgwPQ5WaVawINTBSKjbu
ln/mHsZNW8sBDgkdvoqmVe6yfjAo+I9uRvIc5tBdmkQEXIAoCdflgSj9mRtKw7gC9tOE/whK8Q7I
5tavL/0MjNyf5hoUMp2cigBQEi7VLOtbONvZGhJchEjxlvB+3lluWHsHsAZEkcXZOIWa492gInpD
d/y5ZPHIcpfPSqsjtD/fxsSJNMvOC/OFNrhZn4KL7uS7vC+qpPuaj6w8AZYGoA1+Il7CYhDJxi8u
Kn5qWXw49WYQahNpRZWnC78RgoSDbFU+xQGf1DUzhAoE1OvsEa5UG8+JhfC9YC1gHKqiY3A9QHC1
G65g+jgaJGAoPajFMMpvDk4Tj/92RPAo7ugB+14EFgBtDj+2KmulDALB4XuK7hlHYURxx/oKmHue
tspmUsxQ+WO0LcaoFDeXybaYEtwLJXScNh9JCqxXN2vpOtCOdZbiDWFTSM3mWZyKuDvBnMKhB2bM
CcBNCGPecGBD72O+6OCZQOu1czbEGkDwuozxdAQWiudqLnKWH8Bib68ScKJIacMA5mp08r/eq4th
Xhw1FepKALQVRU4Eh4USmriGATie5LV77j3aWYPCEwZiXs/0PnG27sAqS8/DHk597ef6ksMIsOu8
DhG7zifILwYF50UcGyIMInFPwrBt65Drplgmt5kK/lj7DpMJUb+QRWNyJ0oJyFGB+11qmVqsP2uh
9aWq0m1H1nj2aihoEYxmJHDsyS9Oxi5v8r4lJGlR+qFTS7qsuFgU2tFL/MCnny1u3ncWIiEQpmi6
dOajmCytPEb7yty1LOVmUb5gc1+DEk4hZX6ogXZ28i1SmFFyzhU2H4t6Hb93k3a0K9PiVCF68Phm
vquco1KbVNnWO/Io2V5nMrtIpvdwaPACV35ATaw4ez+FSYTFDWkt4/BjDEitqy+aeBTb25/5w9O9
jtoP3iQHEJIScWWgmKKueTdEHTb8Tf/U9C7RzTi9bgZeFT/BClcODj4VNjNjbSji5MjT7tfW0aZa
UhC07fj7j/miCaYDZGNEgnUZZSrk1OQeQVIpd8zYaqTvGiPb3LSNdcYyUhCBVS1+k0jHmNNuTOmq
jm89lCUl8aorpf4MdoWAQ4O2w8mlV1+ZnMLytC2sRl03mkxkTXpXBU/5GG3cxa2RYFQZjbKvo2JS
Na92JJs4+mha9BkyIC89G1T5vdsEDqrkcZWi3Y4JIU8R8Kkaouw5fG87pBrX82jp0l8YaHGCqXpP
QhQnvMIyv979psaPKT5x3uMjt4D+b5XBlgPDTutFYJQeexuJ8/OhxV4kaMW3DRey54lW4Hc9fPBK
SDYiDHxNNw1/kpc9s35/uLAMkBWvLDKWuy1yGUGDvu2Itr/XX75Q/5PLIX7S9XJp4hM7WVmSWUn4
gK8iye4R8aVDHe9sLneier42jKVIlktEedLj0pyZh/+G7L7++E1D55r2KyWM/f59qZEelYYOy3Ub
k/xmn4EkepphfqZ6D2CWX7F1PE/a18EMs9zQ0DHExJ6vUY28V+p5+VqaKHzd51/FfxHheNgsFMvS
wtZ17msQtlE1CEDBr/drSIm2PYSQO6gdZtOh3paRLo8mERO9VuZRqdyz8YvuKqQYuxANmNiy64HW
fl9HlJNvNGISWHjoAp/hSeHqCf06l9fWOoYg/KCS8tJOREmzNSOW9o/IOt2FhVRogeQv0GPKczPd
nYqga/BfCCFkx2GofQQlV0vLopL5Yc08fCOzPgcrXUCabKv9diXnOOwjucmZkq7Yku+575fNtttt
utTfoYlH9KFmRf43JgZtJtpE8rStdQtjzE/Y8GWtGQwu5lyoYKIQY0Hg9blLUo2BShZCRCNMaSmW
wJaMws3Vi0ZO29ec4u3jZg/lszzoxjtjXHjfdY/FNgxijGa5M3CgTXEg5bU0mMrA/A3qfTGgknFH
5oKd3PJVOn7gs1/ZB0pLzU2c+CyY88NHFnPXp8S1qnVrYBpZGRZZfkCGIlU+am8vKqX+McTwARSW
It5BjxDVdZr8KbfBYoXcs0auF3E2jfl50jLFmIzmC7a2FRK24ruSXdEdWl8PY9+Jf1OQImAe6tAj
k7QUCz7O/H9jCucK2x92HnehMw+jR5GoVeZMPqguT1pvgCMWZYLAqytug226vQZgZ1d9CbAumO77
vQS1RijrytHESxQCwTbCGccq6gyO/tPPkZezIXbAzEvw1QddZYMz0SaF6zdLb5btFYBPoiXlmlNx
WjDeNEWqSLZELxtyO8ySHAWJXtZ4cN9hRo4Zb8iiRlNTvFiNmB8St8r9CLnQU4ZTGLu5/fjsQFTT
wXZvlhmwHkB9yPf3Fjr9s2k5zLkSFbV1Bq2MrUqTHGBhwrVdN15ZCruoxQyTkaLuX4khfxevJ5un
gNPCnk1vvpqN+6z9ExFWot221AYTQplcnyhLv0P5gkbp9Enh4aEd0cN188CdrwyRR6vN2F0WVzYS
FjFsosmeDuWZbz8J0OcTL7I/mCjhNL1wHP4ptV1QzlvI7o0D3mxjhvCSq4jK3qxbYQ5WtoNfFuQq
1TYNhtJcyKXwIzAaCztZX5hIgvw1WD4GdMOt+AWbWuuMyKci68LLEfwJKVD/ZLkP0kQKa0/TE0zc
FUDUmAIOFHnn9uwn9T4GEKv/yBodu/mY7q+NgFutqX0C6E6bTfQ0Swz9TBcXLeFPTeDJblCKqaNx
fgHU6QjorIZglGzsely8Hj4nqva/tUCD/yLgxeij30m5C+Vw6oeWTQBM/QAe/e2gNgrTKflQ3Sxj
CP+/KlgJVWvKQfYoE77/Ho4lCmJPN0xrn5jnSCs4O9WFcVz9J63SLjwPsqmiaNF13500V55CJOtU
KUYXsrBQRLdIIYNYbxpLX2ru6bxTXg3iwA1DQmGp35zeSuE3EiRJQjq1uVb5DQLJ8Nz0Oo86uT6e
YE9+xcqC7LTTeHETn6wrFTykDHuq3ckp4ptHe7Kocbbl+/fzg0xLwkIYznSD/W6mOn6yL4p20DLm
/PLeyG2ewbSkFy/jVGM00sqbyMHHeEpUplIWfcvRzCiitl0B9THUyNgw/MNR1L6y3mEjgpqdiYPW
QKc+5S5F32o81DQyCWeKhuYTM8ExeSMyCeHRhT9LAK4V8rVBGTwJ0slTWthCSZWHXJuIXL+blq0r
ltA/zzlJKH4C1/oCyeqJXMTeN7UCamZxcZJCtfTkcJyVWLFJMi9nng8kmf7sVD24DInV48/PpHnL
zK0TdUqKr+Qhb9W6Q/LjkGFBdXc6CleRqoAV0NWiQGlAcdLpXU56DgNP4F0zUGmGBU/AL/5Ou8od
EDN+wapH/VyZT3fSlMcgAPKrEq/OXSN+WJkz+AshFJvi5j4L90Ui6uM3bDD6gqZO4WvPSeKmLbpg
Lr5jt+bAIV7xZiGv1Fo5QNpZkOVG5GSKBrrFgTVKKk053ihoc6Ylh4AmeKeEn3q+XvM7urGemDYB
lx1ABb4dR2v5t0V9hJISPGJoLdlFP8yyxK8gXtWmjAS3U7cbNzUKX+3vJIrtpySY2ErUFaenBYy+
xZhE0ufyFJ2YR3oq+my5Z5ucDsQmI4VfXz7U9+2JRu11AXf3Ie6qyf7qTCLzDRdwL1EjqgjBTIbb
D+hP5oN5niqZp1YJqbO2rgGHYPfItionptQZ0uYochTiH/6zgpgwS/hIfpHlg+4/vwEKW9lLHEEm
mjh67nZTlBdBn5KMG63uRCpWvz/jHGiem1jwzx/n2d6AyZsXPOYysteGHUPJOtFQQJBSlYeFGHQe
WkklaaLwc+p6tjIpzSC1L6FsezGd5ML0SFKA0d8dh+FNggx2qmTrTYrjC8q3lolUI9XcUMaNH5kO
V5qwoSI7DSfHBJSX+85+X1Hzi3q47IyQBw8pYB49SPu3on4jiD3IWs5ulWcSJhO4aLrzeFowti6E
FuBdhLxhpJWzFEYpl2cXmqqufbmv9E00Q0k1+JeuJz/7rHjnif4kB101hdBRUnOX4AJy15KvzN0c
FA9cf8XAcMAc0jmC+s7ChaPS4u8Yo5TzptcTDUg7sfVit7uNNHlasiiR4FjLwjVJUX84rXAekOK1
7h9H+VltNlubhniGxrLV2JITukqaTrSS7jMGOAb4DbPFlH2jcBABOgtOT30bmNZF+VUvrKAxAKMR
hiv9pvBuEEiadwFvHycVBdOPxcrWGWljaAsDH+gvBBRzz+UQgYT56t9UjI4PO6d0PIS733zG4d5Q
rjeV2TU1JJpaeRizlhKhVUUzf9cF9GBBdHyB22eOFmnkF9E4cbILVjpAL4ZY2ZSPU7muvkkI5ZLN
Rlmi8/rSqUATH+hwgU1S9lx1z0v6wtiSKSu5E8Vblei75KAPVXTm/lp4Fgv0+3qIPCag1D5GddIo
fhljw2A8TlvdPXuhxK+DS46a1rE7Yo0OlPnshVrh/qfXLt0WV28QTEAKxF7ZNww5qRXEUpkaqDso
cPR6FwjeGxze2a8vNJaxvmjQOE/jec3GOr6DSwsHXbGI7eWRuoXbktRKn8B6MkRgl19rAJH4FpWy
D9dPPrXNVkjnwsODBTfm6CR81uD1Gdf2KXV3Zw66Bpdf0q8xUwoPbTJIAuK/pP9pK9eaHM3iTSCP
Z2AfFoKYejFUMeDJOye8+IdB3d+AGT72cMUbVBq++MCg2cGnKaGlA3S1U/9jlVPwSF3hPr5Ru382
sJmcfepiB+pVdzrDjzy1903BnBojG502xRqajJEVU3BzwBapQc/v88AfSxn+FsnoeTXq2P5NAZnd
rSI/5OfSiKEqF7qEnV0iE8QslbWW3bWeXMq1lbuazYhjKcGt9HR+mKJfXdFRtgsvz01NYrVzCRZg
r4h/1r4d3ppQmPV+xrMmAn04NJa2Gf5J9h5SVH0YEJfFWbxY2spwxaU0B5o1nPBoINuNKrluRLPE
Y+TFjij6uqdI0xxBIHaAQRLEy7791XS+NXrfczjWMTnFy5pU8hrSapziEw1NWFSPtn6KtxQnbe6T
sFndyyRybOSN21aIxxS5VHmacq8+p+6GYO96qgO5z+wWvQTutxnlIwoA6qotCr2qMLGHYjBAyWVo
44JLR1I/01c/34WN3xP3/KRT2bYAK6ZuFiTbE1QWIiz5DMSgLEpYfGbqPPwm1LlT19AbcY7Wk6XR
g/vzqJMLmXZ8KF2mLFIBVv0aIjI0JATEFQ1oNeYKj0ivDSRjmBDPypTHb4oQFohb9kE9UtFgCCw4
dCMrksjKvkoOycDoLGvTqLcVy7JF5aj41L6Np0x3UUyX7gQNp8L3yCuJFA3oKWxKgOJDNJSo+u2U
fOOftKTvC8+jE0oMrMXYqu6nDHbhj3DRhVWJW5Nrjmp+ol9aYJnPGK/OTAO5ERMeS1i4yBNo0RKG
I0Kwk4lkJTi3Ba5pfSzXV5gXv+KI/V2bmhotwHoh1ItTYDQ63uS+l4//F1ZmChBXLi7X4G3j1O3G
kcR6F3JgIsfn3Od5YSefjnDDT5ORo473vXfqDcZPZuoUVJAiIDfCmpuWPVoKBiRq0VZgDoA1gkUm
P4cFNeIdfHdDqK+TTOeTTCRB2LnuPd5BqBd/lezemVFfWi0/EYDI6kTcuHg91SovZtUP+ABhHOvd
Ryu7/ktqbswvyauN/hSQdkvXXF8lO1pYS5sIgHhRg8wpX1W7lHiH9/il8AmRHCrp8OcpPiRsbHqO
C7bTN3nKnwSUQu49vttMpIoKqoJxjJHOdZQk9LPbW79z5Z/AHXTQMEbjVIGj73kZ/s8407Fd+ahv
QteQn2cAedYnBYxYCChARE7F2y9W3Gz5X28IDFSX1oydhQjN3lPxB/OND5comRrjzF3mdq+INm2Z
9rhpgy8Rp9ADyF4bEOXO5nQysjw5RgVDWj4X8vd5nRbLwsiV7sXOixlmDQhdPXE7Oo8whcNTtLHs
QC3ROWnamkkSX2QSveDErSBVevV1+QrI4sfDozAvcTFPfbW44E1dfqNo6nxkQAOe8SGy7MnH6poT
WGUPHEDhqUlzuo1/vkX2WB9VDEPooPVfP6ovtTrkv3/OdiQePogH+xLtJ891jTjk6xcv0OqH3cfd
L3cDmBQIL4/Dl2IxjMpLJ4v6glrsP7U5k/6AkUTgLOZJvuEwPeMGW9L0bdFR2XM96hpe3epD2deP
1ulQKzWU2T94BuanvL6kiT3XAv8x34v4haw3aCDNB15DCSfiSXZeMK7q3ICvK4x+aLdHjSevgSBi
k3vjvKX2vNrUjtzUTFWN4FJWDoAuorDpjVFKGFRyxyg9K2c688jvmdXBmi5hF2D6gq5dWTiCuUco
pJ5RC5ATV0ju6xx1tN7HHEropW7wRkgxtLPVRvWaatYagYaYDOdrRQI2zwcB8xWylxSU8t+gb4p0
7X/WHA7f2bq/fQbDa0Z+PWRXn9pl+6eDvNTfuctmEhDdtns0bx8FaR+eU7J2jKueHf5PKlsRXJCp
kRx4taxIl0VgUoFCxHTWCko0f6wIqoad0YOxdKClgMAztUcugjmKoOEyeg6nW5ztkR13GW85WGmw
Lh8Ptr0MoteFL37ZTYwVIYb4sxmtsZwTcJ/RE2RBTi0pmh0hFguVFVDbxHNmzyt22gWgE8nwKa9p
+Z23NT06wPvnhBuW97tTSFnsHDnEkP8S+tI8gsaY+noiZlwaW6lnj3deFExfGwzw0WInuthi/Y6w
dkfPNK6rvxEyCHts92y2IPnDDMGfMeH7IZsAJ9qs4ZI6shPtAUtFVEpAF4t4BBqJUuFN3QB3HzT2
+QgnVQK18CjpyPpA4SMkIsiZwrqrU7z0XA7TQicCauCXMI2MjhLJtI5VOMQ+y4t4/DtLg7F2kr8j
72dCPjsKgy8CfDYqzK2tRS8WKtTaUAZi4y0TWjl4t9JmE5UvRfqZZLWEjtug3AKVxUYCbXu+zda+
B0JaZY4ZWymixIalUPU27bK8Ge+YvQFPEp8B6a5VaXR6dSfUGGprPXdwudHHuE2UCf2OKU9AiAsH
NVczAStK5oAmJqqXGiXhAmoTkER1T17KNrauOON+ErGb8SpYlhOYUJ9kuKDHd7LvU1TuJzSBc7WD
tWrTKm87vlZAJqEjpeIqri9Q5qIJjDplBLEP06UnlAvJlQIBVnlhwhzhR0w/m+BiWG7Dc43v76Jf
swanak4ZnxnzU1RbiWtjA6t70UympZo6OzVLLDJzEqfN3Ccol7KnXEkjcoDFiAGNr0dkWtk1Q/sN
P1+tH9WioA1rimd2NonNq8PSPU61I1hWHdXEdSXe1bimBa/5Z+dtW3UkYvoHS78tV/DEc9bvoldo
67IGYdCQq8zk8ojp8rZtYiAF4P4oONT8wDdCsPJQ9C31wMKaEMMdb9NzF7ZNe3FVLt17WupEzOpR
6yia0mdGVdP76YuYLxEETi3W9bnVRn/tYJ/gbh8Dv1b6W3tEyYycCCSIdl6hU4U3pFM5i+AnK3TS
SkXXLVNkiShiys7+Cj9jY1h5G1h87BT/90nS1vr1Q8zWdos02j8twfCDjpf/6As2bu/qwecKlRff
BDnVYNrQz0nMi2VtdyGB+s9BaBPAc8j4pZORxDwzxa26M7ei7XmLY7ZnLQJFf3FK5d42jIq+icnV
zxGJJqS9m85SOqy/zlKrESYiXG8OqfVkr1RQuen/FaFGnMQ4fNrgfOvSuQCPsJqe60SbeWbdQTCL
1lhH9rceLYCFeVdQfzY9MqT6RFIi6uvikcnYrvB2FBgvvIoEXAaArzpNPuENGdnO48xl1qYCOO/p
yMpSesYkj3XE0hyjF8v+mrT3fVMbt1qkCNZfup8UfzXAMUzQApVTYZI+wV/hEXaP2ddxfXxHuECj
6qWNHTOIoLpwX1wsKRKOYo0/0kvzQkd6lutSaSWL3GAJZj/aym3GoFYdHdqQJ1IizIEUtX1CkI22
8FaajfIqY69S5r6OwYPPyGgMmCoCtTlMS0o/gb2cJ++FdtEFL73Ga3NuxodZnilHGYu0Urw736Xw
NjP+qwH9ozGzO04kB8ZR2Krga51b4efKozNDeVJcwTS/elZ5LK17cZR9AS3kBTSNaE93e3ea2VHM
VsUbUEJhu6e0U60YN6igJghKTIZQWMGu/3w0Q+NAr5FgUDVcrillwJZvRdgNvOlqnAX7K96E/wof
m8BE38sikcYwu4ljJ5mEahxBfAL5ZnfIDw80NqMkD2gUoqo0ZQOhFLccK6ZWIwpSGhdtqGBHumo4
Ce+Y+fxNdUuq7lMNVJ9ounnnQwAk0EXqb6SmxGLtgPv3XbNBtTaDucx1vzbjqZsF1K+BWSHppqxU
Bq+yVen8VnfRe7EhdSX1OKcykpxafES8m3Em4917IknUphho7XJddFOq4maziSLTrDAA9ACGySRl
VP269wD+mYKNwKxxGZsXUa0CRZJQsK8fxI7l9SnLQ5RkQVWOsUIBEBbXvHlgXL3P3e5kM0vBoBmt
dnCybqiLyT3yxMc30v5I1LLo7gig+HCy9ruxjhFmvHV5G4r5+TBPFuk+ECEYEfX1QB5g5foioz3o
FiTmJgetYDNbZ1lpHNtA3PQnN/D+xocDMpWyqIFyV7uuEtDC84YxhTUxjvTf/I6/drVHSkbhlCKJ
M8nleS4BrfOKG2vVAnHa0vhyzYuWCyQ52Gg7wD++f8banJFX3oVil1mwyca9puS/NQ31SLV7e7ap
qB2+C+KfdE0SIOQMuHsAV+ix5egiU64op4rhLclHnBxkf0j8PdQow+dwxiPRZa+ic2Ylc8LLKDgO
GugxNlvhlSAx+9ckEE8EkcO2h2iDlb2K68GyHiPk6ozTE3d0oH7yzS2ShoPJDs54q5JXD9MAiogH
87l1Xi2C2ANu7t+HA316s0fsTrshuKqjSWvnvZdjRHGNXMla3Ec37umYE/o4NyhaeLgi8kR5Ptxz
Vhjqq/5MM4EeJovcQ1YcgrWzebG75U1vv0pbWFWtsqSGdNdGI2ENR85+VaKlyfiWwr9YrYUdKqER
WkA2qnf9w+tF8h30KBt8gaF37uF/48JiQco+LgoPYWxlatkV/ZkEu2qlKqMqzPFKs4WZD/Mp/B29
6aoi47WXxShyB+Cg1PsJDAr6i4XA5HHsRI7KBoJXCUCfck2CNQnnfRpYux6ni8e/oFqIa50EVikl
X9zPIjRN/22SDoIAjiOGMf2aNOhtvsr+tQBmSTOw2n2hgNRvmTHcpEOn+cIL3qTBLJoBvpYCk5w6
ue0lLahfyZ1EGkMSjs7xHa86Sej+hrNEhM1CUZlkMLcDVAQ/03Xbk5BnCfOywR94Le5S2hK0TxbU
TBzopQJX53kbJWiHHhv52vrBWK/K4cbQRVz31pbUZSIH+nk2Ldxl3oMto6yLlcACjDgXfPU1Tow2
l5pSbSC4wBz52EaKJjg1gduZ5bCOZiMRmmyQxELB2ztXe5g6SLxVDcR7bqkqjRkMgIOkoCvCoOuO
rmuv8rYGIum5kDTIy4E5kY0mf3TUwFezzxD0/BSSTwj2gUxdIEI2B4zEvV9B2Uepmj86DQ6hWH3N
WRnA0N0swdOZSKCpF6t5cXC2UglSWihLrAkezhUuErBawVWPkvClFemJmPEEkSUWHFxYs/NOMeqm
Jbuo+a26NXDhQJgaaSJDmyBfeJReV76aW6tPM6HOiWrLnlIBQVBq+RDk7Or3wOOtcON5gL51IJnv
EaJbfHDsiGCNP7KsgFqNdQHW3ur2euo0L8tBCaRLgQtIJnGifGmKYgFaZgpCZoN4t2gWfJ+fYp5l
8Su2typMuJYz+jjybhohPlj4WmM3u/sPxIu36g5npkQTscjFLGI+w775/3F8VJVdFSYdOFVMtHem
FXyuDq9ci1j9h7zyuKMveu9STsXarXq85S8VTpc2Cxe9xLgyJ5LhLFkZjHAEl4iLIr/h4TFCrXct
0RQGp5hLiYORSyy61EKsc67schLg92EP6opdTOq5e6C2czG2LPShLULCQr5XN49BMfHOxW5aTz9q
IIbk0C97RilkSko3FO7km8GJoOqXNkX9k2z36ad5WESRMkZqg8OyJSKVilRFJeRD4/pYnzMRkIRj
YY9gBT+Tm8d/kewrUrlWM1BslLUcL38Jr91MmOa2CuWPDgJasJqDYhosBVyo0exerWSo9UYVEEcP
vQaxF8XXaW8eQfiB4z7S9PFWNxqBM+xR2VTaDEV5X10BeJBOBJnYa5Z0Sga4LFWHvzpaKtLkLUnB
Tng5oYagFUllHGSo5ldpn8zbShyWl8SphLem2X6+4QC4HItATmZ65vu6UOjSbN6Wixk/9i4nrMn7
eumhvBaTDLZcXHU3XBAVZ1HfwbdeQGgq939SvCoaxsPGGB3moRAi8iOS8/rNeypXkZfixqci3EAk
OyXljJNrZ975Vkq0+R/UZe152c9dqpnO1zpLVnWXqaJZqdEGvmwHRDq4njbULlME7Y7TtLHPXmr9
sjIVwVj49rD5GXv3jJnuUdGrwHee4G6kxM4c78JZj46QaqUlJgxxZWGVyA221WQmoISo9ZJP9Zyd
7c49DtqDuoOoJ0B5EnnL3W3X94sAboMZojFAEp8BaFJ2C3KJwR9GC1udxmLyJclTQH1+t/C3NfI+
6R5072++SebBFMqJxygXKDRf0ngoekYN46H+5TRKgK/nH3pI6x59dpgS9YL7BJnwKo2RbSznrUdX
9H7xNaWXv5M/jLTNEoAKKZlcQZ3iL2vUwtAlGZRiOJ1FMkZQ94XoQDo4BRFEWKHim45curyj2+UL
gZjzwOTLxHGIL7gho/Bpwjz74BCbCNHOuDMuG6LMSBKnizr6ykHrJNFlD0bRU8EG27cIv1ATrU2A
vDMKSzmZN8EVWicVR9KZzBYNPQZr6OW9kzyP4R1X9MMz8hyBrcxwxr9hucFgLuGhnl4QR6kRzqll
y0hQXTult8e7GIH8VTKoEOYAvYr5iL/PH94QbbgnBZqtf5GmD21qmL5NLYN04yOZwSLTKBZZyHij
TJXj04P7QogpWj2shLFOajr3va3LA3Ep8KbwCc8YMShmnfxpOL7sS39jw81OyKlEz8YE9ZsZGsBD
zpLExMuWHCuXmZJy9e64JpxrXwVYaVYO7oaMNh2Vj+0tgv4i1gNM8IXlCThr1F59FEaCsL41W/dB
PEfCyyeGyMVEs8WUZPjM2oF1lne7hHIlEUaeGFe1gOoDVFzFLBqcDy4VHyXkLCe3Sukws9exz01H
Bf2tPSJY+ghb6Xszh3un/djHPplEAiivT0grrx4KyDx1mkm+aGczAVlpRqLajaHfk2qJOk5gX3Fu
qjjo8eN6rFFD/XKFd0cNDljtVZxcJeCnJnMIOLk8Z6quzOaWXc7Mu0flds/rFLI2yy21PUdkQmu4
aFOnKiJZSH6mOEJZ7xIelPORJY/+FHfXnSiPIYv4wHcRR5tlHCQThzRHw9wLAjZ5O7xTVn32JhnV
nuwzs1tbcObyatYFAcYvOluvQ/rlhAZHezyCSOTDdhRdNrbpTr5oXx57CB2/qcRePSPmP9423fRs
kKk1qDn/qQCNe3EQv9B80w6GWYhxsZkI8hIujtkgOHupPUhqLFEt0pm4CZR33z+O0GSLUZWnqEt+
HiZaDQ8/6jhcPOn+6mMbaCU+aGNjJFjGCLPQ17dUFYJFYAEaAsUxAiszEmO/GY3NLOjbHwPlN0gI
tTpIMAHbwCd5CRTKXGOEuAuVPunN77WD92LHHHyJ/fLw9R2hbpiMFAV8ifulA1B6Kas4gsTozYy+
iq4E3FbkP81cBzeS3n+l1f1rTt9GD6ZEPLZGsjW6rhbxj+3s08e5EW2bOLmT05Y8AxHWenL2ImXa
gRb2/FVd7eeH+WpcgJ8r7oWqKu/l/UzD2SGDOvaJmnzJCDAGcbkxQ3f3BgZ9k/f1lNnLV2GFF3ml
NP3XdZ0Uvk/AjYK68UJg4rcUMprbpwYUCd+IY0hOjDZT5/XC+ybOc2dDSgODlphARJUTpM/1xVHl
B+smWL6zlehOHZ8IXuH8cIUjfchwGVG9hhOA3TpRo1qlUmYDHyc0ra3PQoh577bHORGfdCUknVnP
YNJYpUiG9FamFGiraavcC+dMicztBfItk9F8kF3PpjSmwFOLaI7ZistI+5NhwDCw8WWht5muyx7f
MT8Bfa6ViUs/02IvDn00r9Pe4uxcg43spaSfMPoPhxO5cvEsjmo7n6fFmJxpqQuETUEYGpveJpKH
mXOfz1iDeNyUw06KsAN3T2Z4ens0HzmTJdEweL4KFEj1bPaIa0xMb7n3FKa9dDVmhrDkLMo6Ez+B
2q3+DKFF3So9PXqXfUlX0cyXToyKlpwP1v8ESOr/vwNCuziGyM3CDbtYxMPA9I7vJZCdsaT1fbrS
sGFpZXp82xurcSDhQ5pXBOz+3o9PwB2XT2PbzJW88ItkmiwXGdYcmwkVLNSpXbOUGgtubtw+TT/J
xC9EExX8bEALVGqb94JvGaLU9kw85xshgcQe0y+zQy+01zCwEJTKJaV0LVxHRD9LEyCH4mshs/eC
QkGrrBImN8vLud/3qt+ccYss8kOWHz4SY+jJMxIoCo0vWy28cKW10zbOHZY/5pLjsOdh8bRDkwK4
ooF8kHf1ZdTH8VsXYiZvD+zxDegD4cV4vVynHB5AUqav4LeF216wdfyfTPlIq4pbvg6/sKM2UUPX
aYnbgiOr3GobRghUpkDnR0Edb0Tbe9mjFfkiHJbOVdGZUv+UoEoR1D6a4t7wEQzTBaK206V7BPJg
msvKOHSzj5XjeaVaZpLo6hg9pG2CClbyNOGSaUvSarSnYjUSRMkcz58MXA/eOs33mKeM+qwKknLF
RU7ruqkTHwD6iiypdR0NUEUl1pDFWJcFN3sU/SPqsS+QG7gZ94Ki3WbSW5EHFYhsUieU86zJHzJK
b/EoOGr1Xqg1bkRaqgIsOoiBqZDNSddpP+L9bWZXvywT0Jgtk8e6E8sIZpQzj0FXlicCHGlD/5Fp
I6QWxdAoLsh4EgoiqcQZX8/4YM5TmsQLGWi+12VKRaeXBa8+TksMY6jByGUmhcBGrBGSl39Zcp5x
ZDKnDx5I+Xh+N/4M2aDl1kAqZRNVbU/LHpU7YoWpJkoG9t5sonVzwrfdFUakCr5qSOt988/s0lZL
E6YLhI1fDcHlGrhU8C14FRFKaWyyWsZ9lIEQlfZDoiAAe5M2vdbz9rD4NikFymIN6YU1ydd+cZ3t
LtghlNTm1PtCU4zZMH3qCdrl+9iGtQK4WDM2oOi/cj00rr03aqWp6Ak3x1dVBuSOQkYZyRZX3HiD
1DilTidv/+5CrsGj3tFCzImLRXcn+ikQh6VuD73mcnB1e/lhMSEWsF5SpNpC3qTh8oTeonoZp4gy
XRlzFWqP6o9SVuqr+atbrlSk0hJ/3SjAlN+VWOGGAOH9+EUcSqSEo+grjAYBCrQbIvvYSKXdjcG2
bagQqXk/8ERFwR3qu3pHJoI0s5WexEX/F9/BbxoiDtJN2M87eIDs3A/feMtpXHU+0wTmwuCYFqC5
kZYkl8v5/shjf9FWnNLcrgBZvAEgV6ZyA0ziJq8tkTR/gFQKGZanH1CFL6ycU5K3GtIm+yz8aW+J
ezk386DvsppOZl4gsea5IC5yIOEuf7T9jDKWC3AzqIoEdUtv+Q/sTgNiyM30ZjZKP6y6sqIPnpoF
ohPmHQyzbg3AipVjgEQjZqI3BUtMveV6jpUopvcs44hcKifrqDj4tsepJjsQfguhlo01wRvxidtw
n+56L+21mOcSXrwBfQcgKt5EIbvmtKli4SJWip6WZFTqE8taEosviNOmDf28xIRg7BWLwT+06H7H
e5fD+RGydc+Ubbdz0SLF0t12tfHk+ewKA2h/DRivjp2TC3hg5fm1maiiPjeskEvHk488NEzWypIn
eUkuQ9ryftPms+zfqfokUdsCZsmKlhN6MbHmd38yI0zkK7xSVlqTneistQsiiWxy/5rXgPuDM/rT
Z7xyFR9ESkhsSGmkEw8JsU0btDZfGSyhwcizsF2Y+Zit/PpLGKrUaZ8XoJNn3b944Jtw+9afwsfT
N4NzJX0gZKjRfst6Xbv139FCd1mtttNrarLGaeY5C1yiSAZvs+oTVeLA2v8V+UZ6a8tfw5KNAkRD
fEh9+TqOcxMI5//Hn2efwvXgdyQCnAlL9yJDX5dMJAOy1Iiqb7aRuCUojRkticIbdxwUAv03Yb5S
Nt7qTTSXzBFqrT49IWIw09PdevyAehvjXScXr2WReI8ms9Ep7nLOAgVvygkhp8nLNg4P1JjRnhGn
OzGOWpyu/1WDDw/lC2Xfljf+dxe3UTatsI+enmsAosWpTeLGJtJxqFRyDD25HnBGC2BFdEVQXvwS
mIgDJ9vYauYJTREp19O+ja6M9rzau1C9+pfKE5m0uDn9uCbih9RxH1GV/kFCXOWm0yvqSWkWwk50
b9Okdw9Xb4JT3GAER2eMA+fUKLui02ehqFgyQ3REsPBVbQ5y6TTHSx4rIgGcudo/VhIpaIkQjtrk
J70b/wI2it6sMHevwxGkInq5wCeeqZmlNBxfraG6NK9FiBFHTa92WrDNW5Vd9ZiNs933Z10GbYBn
H3hxEUM/HHygIH8MicrSFt0ffl8LqlTz2aAYf1A3ieA8YuYSTJDQSffzGwzMVFGBDBodYIhGfosr
6D21gJbYOHNEE7dm7PNgwVXrqJkSuJAhtz6mykWWaXb1TYVYvfgcqWIyxt6bFpebx8mkQtrUpUzh
6ZwX/xv5e+n9WRk+xnpX6iQLspdvVaDpPhJ/JhUIGXQ/wuKfLPdLsWxYuhmc7bg90I/KKFB/3W9J
cMSGhEnNMA71RreN8oRbQUnUxDpIs4xeKQEw6/ko+fRTnuZNdV5OCvF3njSDP6NK9Z6KjT/lgx+p
DVBeitNfLTSbHdEOz36ShHmemKyLTg7Y3pN4kuvfW155tnGEbILE3R6glc+g1F+CF/qJGilcWxKe
Ua35DRS/x93gM+EPDQPdsMl7YYSvbx0+z/Nb+x2J2vKiIr+P3TARdjO6rCn+FG1J+mtxNP6EvRP1
Zwsh0DNgkxyNPLwZGIncOp51fjkqstcNmnqveDEN2hB4iSEyWhJpwOL1EkcHjkdbhe2HvmNaqJ5f
L4hz6AiWKGRgqBniuztyKzwKFwDJhG1yrSmhJqfIgizB6W8bWjLFhyo9oqawVhp+YnYX0zCzakaL
IudtMHhT8JyDCKFxSRpsne7LSC9SbwRFcCsjub7lAHpG1lN9ceDd10LBzIsrELQmE25BWtx/eX/R
aFkW1HNo76szqZWmAWPfiNY3I3HWBmmq1epcVR9adt+8mUJRbB+CMddJasLkOIisZCLDbgch783b
jxyj153vRpPQBRanw3hpzKk2Gg6TGQ4SpjrrBnRSQJAOWuABoI7dRDxVafDImlCgnveKY3tdIXF9
J1gA2lsripVgGBRg85015QQUX+2eEdYqzxtbM/CuoL01nnY4Ey5Blb8jUvSDN+mfSt6AWe3y2U0F
P8J64ixnE9+0OayzXhSkaVWVv5UeDUWj8MCdycGfwgq/RYktT6AVt2hzzLyREsr3/IAJi0KzAzMR
rMl8mBJmQfdK3/8gWDnUHHPHr9oWFMW2qI3lFIFYBH6uO1GpUXFshdKd8kCVgfQFPLiHw2TqKk+s
3vN8LBe+2LonvswD2iW8/5sBHniN45QewQj7PXZROkLElR8JWc1wPBWH9EMNziOodVLssDe3rHZi
pQ7+t4rloOYwHRedGWyYqUN3FGVJWdm+1nhi1XSLYZKYIilaSZQin8W1DZc/abY7SNynjb2w6rXR
kijLIIGo7K0WWvYICJ3JC8APei07IIePqSSuZ1VgjeGOK9wNyUXtbTqM2u7uiksGiJUF4QmFaBvb
RH+LkBxYmpcfWAsXpwN5ZMeB9TiE34JqS2/Z4dN1ZXho0qAGVuTyLy2s8/pHdVGmcN1XnmNMm2ES
ApN2SSDr6mFRmepgR2PLHjJByihoitx7Zr5EhNlONbgZiIAQeQMSCT7deX3vO8+eBiH8SRpUx1E3
0I0J8rPBgHiLyImisQlRUK5msLPrZiENYsCPDwCxlTQkBkA/D8bLc+XMiZtpFi/mDZhmNq+r/6cS
5pLQJpXmXcJCQEwxe1uNOV5234v07LzAt/nM9Oo8nCky3OlKOXpUJMi2Hsdheq1j+9KXMiSs90Zi
LfK77c3LJhuiWoQXuqxWSLnKG4zz6q7bo+/9igL9pp34xzYkYZgWnGDyR6j/TomnLIsNc9iioICi
jFJjmxirOsUJyQq4Eo4ubeHeO/U1ijUPInjvFQ+QuOJ9UUews+zORg/cem3iSfGS37uWWSViqLyA
fR22o+WaEFqbCQK7xpcKXc8T7Vakllp/OnqPHuP5UbVd1ZLCdBNXxrbo1m+tXBUpQlcuolOowSTk
90w84VNWVeRVpWcKFaV/y+pbim4cMez2i0fauJ/S0y5Ibv0e2ohxlakFtj9c0OwFOGX2ZPHenLDl
eGAWV58GCnkDhmD4SdnsrgaBYkIbeVrc7qc+x1NQpV9AURJcPqb64NYeCdE4mVe8+qDIqwPl/sZK
8+4GpMdVH7g9ZcjvT14OsulcvgH24vTETD9aDYG8SB6E4xz2OkiCOuxMPwuBOUo6HXkdazI8BxKu
/uIuMp9CxEOQaUX6NIs4Wntx53YUKJl8P7diO8l7Y8ghjc2NXK3NC1p1Z4jcL4+Je+B62HiI797l
TThKbh2hn9tbp2DFGPFe5rxMxGvZ1BdY6NVSvD7MCoAc2kqrqwGxFt6NIx3cq1+nRY6O2f6srXaT
vcuafkhe62YWFn8pUfk/6nyP8tW9U5rSkY2swguNIhGoaqsZuNiU2WDae0u1XDhhYp2eSA4ysLBH
dz+D+6c5wjNDLQeCtTVEgNLqRdNN5I/rRkqSQPi65n4uwHNV6KUoiXKMFIx4T1dHDzVNO4IQnNR6
0ieqBGXOjEFpZiTPheyzMjz8hDuiKIWCly8a3GN9B8k4FfnC5mcsrjKeGmduV8ADAGKenXQX+hz/
WgfJWVvSPgAeBpU7yqhd8WcDIYThMs6MXI3i22VVz/CiclA4N+D4T8Ro2vyny5K/g7Bz+KJmGavs
ChrgKAsssIR4cx+NeGwwcrrLPkK4gPRZGiLCM1w4RXtYFH1vNGIQAAWsQmW08jG4aibXKsC219Pg
nVnUB/zye6g2WXNrot7AttEYOXmL/2TiLOoaVIlFpEHunKy4ffsvj4hJqjKttWqHTW/XGVGJKUo8
ldBpAZQsHmpPXnt7RmV3beJyVZ6FW8Fmw3yvZNhoUMWmqjh8MfzTrZ4sjXgN4Du0waYBGlAfKW1D
d3quslxAWcK3DAXek0QliMo6FblY6+f3h0FLCOA5rlzigyXyZyQCN9IPoJrSJLohA6OGlXU1OWzI
cdDX7nk0GslOcz/y17k7cmTFQcZfXFL5sgv8C1gTkkEqiGMKhX2ny8GJnkWm547jGT80EiwvnmNE
Q3eWXqtkr/bIiy5Yumau2YiZ3sezcSv5rclFBfI7rgXV1zVyiD0qpB88cfBIKoM2wX9soUrkik7m
iLNzzZi1wEpvPX8TLB3icCe95swU2LzSRRfXf2Fli9wHbojEwzxN/OHd1hLEH95uAqRt2r+nEL+2
l+xUfvAbivcgzbSkU4q/bITdgzUw4TJcocO3Bi2AIJaRM26+A7nRUPYtF1OZnIV/9ruBQ9J3MZkx
f0zNqUAs960vIKu0dFNrELovikiMowtQsSBjqoehNtUvHiEPHxvdKfvFeAe2RFTWsuIP9jC4ZXiB
CsPbO8JRLGm1BTaChUOZCmbHg656u1EQE8Cg3dPnWkjS2TVFwHAMZ6BS1Eash88ajV0/qLKqgAmb
nlYjVZVeNhcxuZ1eVJK4uIplyUfp0bt48JLKMfr+uGih1vGV8iCjl6ZCJVMxRPLtLYkGnT2IV2o7
8sgPiQD5iWPyrLCLOSen0grO7hAPsz8WalKsinqIrjvKWm8MrW7G0EYFdY4B1Ix84uMlj6kJtCif
OsMRkVB5soM3j59D04KsfWtzJBspxWnukmJm57ChjRoRjlWMLgF//khkLMB6iYrLBA3MffAiSXf/
0CBEzgnZeX16nethhQKr7AFMhuhpOJFLRVlDq2x9DA8veKPabIuSbUd2D3135yfdaACgF4h+tp1b
ot3vaRtdSW8JR5QAFqb1Mpo+sVRCDDyj3nBmR0w7RBYrWsMve8U+dUcTP25wK+bbUw8Oq6xJwJh5
9aiOBuvnoL29mGj5xiDfmv82SZyv588qx3tzy1DubtAV/WXEeY+XqWuUfv2zH/Ihj6W05nAL9NwH
QS/26/h9XtIWN8sXpyIeR0DHsoc3eomc3j0ivcYyCXiUSLXKwEMYcBW1Bmm9rYXQ6Nk+NS+R3oD1
LcfLPYUInmwwmmqV2jw1H4ea6VyOfvy7sD2lQRNJpH7wyI9vbP6kn3PDiqfFQtONSEReiNuXuGNC
fI36L/SAAGEG6dfBFeIcNqykwObpNsD+Hp6ibstNygGyZnDspOu31TnHjaY7p4BeMYlP4R9IlApn
g1XOrnytm1+OnxoNwuPaJ/QipV4ILmA/61S4Bwk88DuTbQAAwIPPSkGIFhNkQQG7CS4FdBOon/D5
VRlxVDObtNKAs5xs8KY/SS/TJfhcO4z/G5vueN1D5zhStX9+X2F6tkXsSn5Iv1dfSUPGm4MwY/1J
AwR/NoCrMJhbvGMRMaPxI6VzoG2m7G9yfTRFwIYsADB6BjE0cFbMdLeZ/g4KnaSWFjbFV2n9AE4y
sMvJZK9pJNVRcVZji8+Z84Bdme+NQzu8QK1d0CYcTaWDiboJ+d1A/7WrgtACN/bG34fTIz+eHYuh
X1X8TLKx9SmuU2p7BVGHhNF263Z/x69KIvGpfZAtRfsS8dYjjk/ITuTF+NMdlQBLVclYBa6bXD2r
l9cLbbashJeok6z/2mB3y4oEae7pqqimSyZ0cGJbLqIAe11iQptUKjgbxchYdd3855xzjvNymZ0O
YQLeOWUuUH1gs8hGjw6nd3sXf4B8fgrUuzxcvaP3ZaBOA1veWpDge+ea7nkBO8CJNtIJM1FYje95
3BO6mtka2/obgaVTH7jDn3BlE7gyqknsZVblzI7m66wgV/50pKi2byN2DiB7u5moZvq+6Lq0iKjS
Co7AVw9OQZz9crLhIo8ZPFoT5yNwF/Ihtj2KjKPsHsUVoYZtHDfNk11kZuImK6gZl7KCT6IIn58p
eNs1q+Qz49yTLAWvzq4qLj6Wl+zvzkv+FDPMi/u1EwRyi3EP0BUqosPDz6FfrMJ4brY7Vg/sPmny
qfYnpRJMXH84fG/RXVq/A9QGK2fQqaHsMp9p5I1by0PXSIIVPwyfc+ZWxZmCSOqDPV9T7IUMVcNM
XCCyCi05jvM0S0AauvbVrNZKW+E02HG7ENRt+PEzIO2PxB0jkx5fsLvWop+ozfl44DsmMMS+ZVS+
s9gqxVYhGpKHRIU3pzx5xTLK7JgvUqAcVdcsY2/PzH3wnkkDIvajFFoaVrtr0hXSnmHxwk6s0Qn0
JzZdAWpZue4492iTRrWWZq4KrxzNNBecPWRaRmpVaVYq4/M+TTPJY57Nep78XGVo5wOmiykBlBwV
PLdA3c3nfRiWlb27mz5OIP/fTRe5E0CcO7rkppztibO9YLt8HkIVS8e8W0K/iCRadGX1DIaYlao0
m9M7MsQS5sl87ku3fWSJH2X1UWXbtUguB4+5zp39jXlI2sEpaTTODlnzh9GbaGOT7cOryvWZQUgI
rK58B/+o/mg63LzVFZD6zb+CutBmn/4lr0E/1XNOUIlaNgLJrywlVQTLcvW9bSG8T17ynbH0f+iG
FLUP30oeG2cjG4u/3lmPlh5JO2ytMEecaBfmQhFLozxpPoWE4ZD7TL3Co8cm24C3Tx1HSQEqBNtI
1bD6FFa60fubccjL6M2VCu18aVPRaziWHipLTiN0dFPN2xURwyff9ZAwAKI9obCI/dDo86B0I56U
yPMWnBNegCigHVY4rODE0Fn2P/rwguR8t1FSJWw4jh/G5uw4tcYdZQbYJtrAdKBkBAqg0SLQOqwy
6QcdyMHIDj+DxK4h1JNPU4AnYwYMjGi32bFyfDqsoAl4CGg3h2J5XJ3nJbHxx6CIkHFczd32P7f8
8P4mUAYtJthk/AkPA90/wnGxH+vJqEEIQeS3WQS/rMdN/EbKznW42ZgSgMjuPVNWkDLqeTi6FK80
1g/ZO3kud8gZCwD/6ohfILbMXKmleHZJTsOmsM3dC9h/XWLtEPXefc48ER+OpXiwiDW00Jop2qX6
0WlWqnnBEdrp6+miKyEnevbEhOE0YGVa6j7D6Th9jK2Wf5WU94nMt+DLOa74zPL9qkpjybmXdEm/
wfhlVg1HbjOJsrz1aqMQo/Vqq8cc4FJbXKb3JhF7E7PlU2XHTdcUbBqjLZtu/huiYGayTTY2B4zi
qELD1vhvugkFUVpWIXFCZ+0mRvtUpOR+urxoWz6hwIuo5eHY7mipGXzpMjdR8ISMj1FVfRfxvycH
2TpRWlANc9JuK/AwQ5ydQviTB5o+kzpKPnAwznmzpUkPVCKwA8Auq2Qw/8W9K6myE9762Pju0Lly
EL1bLMBu6/VJLsZtNDdr6DgxunSGI4lhnf+AMkmU6sWtI4eKMfzm8sH5jblW2LriQv4rgrPaWobS
K0BS10C4iNKhGOhHl4hsCOtdCe9Gr0Ohgdsq6hJor6oW3QLBHpIxYGfu2F0JwBn3mw1E31gqFP95
Vmrg0SmRwLPvtblfa3yxbFIc2BOiKvEBPJ2BU+aAfdEAVqOTmVslOAoW0qRYD4gs2E1YxPanbvZ0
d2CJ/qvoQT95HoVRMxyiPAkE6U72kCB0R5UAkKkuu6QdBb02fBSitb25aYb216kq3d4T2UF9VV8d
F14oqvwlUCXbmPuyHgfE9aQP70LrbVDE3GxZBoztcAJacXEfl+sY/U7T29OA6yyzzm6UGgaa5WJJ
P7dbtPAsLR5iot4+yInq0eQdNZskp0xg/nQa4+PWR0Z7q90O1k9JtOAUplC9786sCIHF8+PXk2m/
88bM2rj51h9lSmQwIfDJF5o4wJUT4OfCXta6e1rKT90krB7QQFn4rvsHOZbxQbPnQe/Xsfi8TP9E
v3/P7lrvN4pDNhtoOogLwc2CKKgvBzrMee3N/KMOKXx7wP+NY0EQQDcp/XM8DuSH/Koyur7EIhhv
lAalNbp6YezSX+apPPK0W9bxlrhv8BfXDmW5+GVGTrk3hGGT5GnV7JfBBUN8cUxkUQ/Hz6ixldDB
91xoQJltSE8tB7guNwMnpgWUi0ZRnX4ixs6AbelobjV55PTNq/cRhS6VijRbgJEiTpWKdB54K8QL
v+aMsRVFYbYVytzDi99VZFJvc8hWlSztHRqPTc20zkAPmPBW7arSKPaXoDMM2gx4J6AnA9dwXuJi
LszVMcqQLXlwxgV66AUfBpz9Lo+pgKk5TrLi3u0bAodBr43YFVCxlteA9cLP1bliGZTl2bnyQzgf
3GRey882TCl4a9SjOolzpQPWoMPFWCKWJPg8mzf6eZXgfL7Mdqv6LJjyOZ3v57B2xIS9XR3VWUte
WJJOmEEMh+2mAC1gub2XKDZHJv6gn+u9PPCyu40AmRXDQ/nCvifSajdWI868UDTxDLlliEmOgx6k
LHKlgJMyksDPM+CVSInlxZo7CZAyCQhVacFurL1+FUslVjmbBwf6D8Juu40siBqK4FSTzWjVVi0P
FBHdpFf5E4ZXbieQkCZ6y/wR1iKVXvf9hutakS5tIGctf3xk6s3RX9ua3m6VqH9GMQjWzOwS70f6
ZDW/af9Fyx+2SeeQaQza7A2Fq3trLkdKT1PPNSfGzEos8cQMTWTaLaRQikS3kSmtxLNoO+kvvcqU
gtNfC+FJogcwWxwAZ8gNrmzo1+phggQAmY4P7eCKiSGye6eH3suNkyq8p/YICD/C0+h6WkG7WNY8
ELytCkjpihXuHswlzwsab2fmDs1LTw2TMVQIMIbmaBdX2n8KaA3MoFmgQc8VDSbJ6Tp45ndEDUKT
Usf7nqTLIyjdATG34QAhmlgzleVJKdQ4yC5OR9ETCsNiPOecf53PlKfWGl5yh9meQ2E8yKlnJ+lb
HkVTFbjQjHpfmw2hB5HI6rdNrd6wx4+b7r+MOFDjLYaOy0kvb3MSUB21PDK7vAHH40hUTEc5MW1L
HPdpX9SlcTmn19NjUy2qMgWYN7XoHpj4ABHoAXsiCJXfMs8XMKxpK5BmNA+A93hKulZq47eywqoy
ASmC9+E7M7FymNyiCveDznNIQCKTxTfsWXajcRlyWHlycFVUFDBDTBLzMRUKpU7LwVu/IobjNcuu
g/aACNcMIdTGPoTr8fT035r9mCpwm4FjzzmtaBZT21kgNA1LK3EXoCyFa6btG2kzjDzuGsd+1seo
2GWVZLdY8xw0QTRWOHTjM0oqoio01bfIG4RycUPA5tK8O4rYBjUrlI8FYf4N+YToZwxMQfhjD+jk
HBgb0mwTPWwVw+TZdc0Md8esNB9LyzjO1OqeFFh0CS8byxEvzacnUPnKIeeo/x2g97EIvQWhlKzj
ZD1gZJmIeVhZSwaPcUeMOFl5qpxe02wTZeNk5Yp+fURDDaKR8uaT99uWqow1iiFsh3Jr/5UuCHAK
kRLnn1G4JmKR5uWrx88yq1AcRP406LxZ5AGSx4/6lFKFNPBe0E6Uwdkt4NReWpnZQDCh8Xnd9LM0
E1qF7poFiGlr1ioDNFbqgYo5Nulnxo0u7qSbnDzyaVtjM9MO+1r9ASEFksTC1vpW7XuKfuTsgKKk
XgPyapqMZqLaQzXAgV6j09agg86rusiTqUtHiYmvPISBp/F8OReg/OzEKy+6+SAVuKQ0E4NxGd+a
ZBqEBHd+m5BtYG+egUuOEbDrpZo+b0EivuWyU4USaNvjbSBiWKDccG2GXO2i5fA+HvPg5aS9Jrsn
PcJUQbUpZw3m53rjgCPqhG+RFEbby6sH4oLYtJxpRN69/YODuU/6wAw6FN+mB/+1hPYgcjNpb1Lp
Ake+x4fuZt7pK+yGKiPblhaGd2q87RHZiLvxdpDYEe1WhdK6u6bxHH3NQl+QBefAoilhl+aQGsVc
ObjzSgEms7h8UFDb26TeeOMC021ptzwdq2v31q/tjoqmRfCr/oXp0geIYX4dZd3bxZxyp9+rz0l0
6//wKx8Tc1jUy6F4u3hSlSspte8a5vBVUillvXmp1EtVEW0X71rC/9Mp8h4ss0mi7o6a3epJbDMX
VlFQznAS3ueJEnhaqd4WnZltfjfSeRDz/eqMwgS89MEqJPAMGQwhqRwTS58hPH190ThRAi2recKP
Ct9OifxwKNataKSP6kyWz+rWfeDWszmaW2dk2gM4x00A3/8lRLOmgQNqE5TK0DyJ7uEzyyAmuYO7
DHx7j22QHdH4eSLzHxMrwCOIQQvV1I2XlqBiF0ekGAS9VFPenK8w7z+Euykfc0ize2W0vOwz+R64
8yepCGdBcj5yjP037cz2d8UiLlkSWMxmhYb+yGnNBsWW4olpqMaINIcg9CQEaPWxiRvRUwM4kbkI
SD3TwGn0Y/lN4gZWMmcoPkmI0TjVKURO7EuOcJl/Ek5l3kvDe6CApcT32UOeelQ5mwF9oDDTxwvS
Rc0DboAcPtVTI/ses9vCNWHrk50+YNvk8nRSuMy1cFBS7byZVCkfe4VoufGflLwu9jdAa3Ox9gP9
q+ovKzlr0ZRl5bYTzZLoOD4CmzAYx3t9DEhBOuF83u6O+Jo/7HPJ6ELu92w88B0gKg0GQ2tNlChy
b539YdVfyS4u0CmpZ7jOVCa9WNvXlnSRsSZZDSilVhpRZx6MS6JiyEXPX6KyA61utz+/c6kb+i9x
lG7bEYkSMAhJS5ACmG5mMD8dQtTywIDCJzjAIabGQ0GKK2QCgmYmLXKqZ0EUI31/7HdrDP1arMMe
+fL5+YmjUcXFzc4D3nZIwG+mqYp1SUVdOGHOA2hRz2Xrax1+LjMvl8zk1Noe7kJETsQBIY4SLAfb
lJi9khWzxcQsMHDAL9e3zQixWCBX8/B5YBLp/aqP2pXYGMHk9nF2tCJ0ES5a9BTUEvoQocMITw1E
QNjnOBEDflw5o2l55k4LbLGxq2XYlLapf+5+UKOsZE2dedoFxJQ6X9YpPGEHlyjBKXiq1BdYMqrU
tKMBiJQHhNgkNwucUe//ZnIbOqM9j6F43LWQKDGTd2kisc/jbvVr0Z50l8oI7OOqLWAjcPVEuU+a
6n7OlrHSC43T0gabzxMK3sd0w5hy9LpeOJx7ay84gDfijz7Do2TtZ9lvvX+YiwoX9qdYl14MCN3B
YvV6+Ja07uXi44SyfWP1DNE4o89b9VDcjEw5jC0Qwx4b+6G1EunxGbOe7JXrW7EH5APM4cBw1lwZ
+gV/0hLor7KwMeuW/DWgE1KlBTx2ug2FEKsvA6LR8AHjQvccQI43VqR43bOwfLqhkUAm3X12zNOW
5sooa9SHawPdOJq79qX6A8hm5gcqLSXDhwsCjrWmEwgezzBBlFjDNOs9Ao3VAfrdO2i3LYZq/vZI
ihspfChSHZ6eWEuafaNQHy0LOOMnmyCS6bM5L2xGJazAzljqma/k4kIYux6h+zEwzpnH+/ykpRcG
Rf0AmAHXXbBWKW1DgUVUhdvSCyPWksRNpT1fwnHg0v0sip3p7qkVrCRx2C21f5JcGVpvjR5gAB9w
cLyHxdtJP8aOm8k1Y3gwCJapMS2pUIGB0P0DAclJLBjTu00+0eRS7LPse6kzvXF9dXDQ/aZruJl5
eTHdMPCajlteJMKGD6GwagPj5w4T7epJt8leSUYQAHrtlc7Z+r1/PFbJwqtcc35BhP2qxz44ywr2
HI9QZ4uJGmw3hlxV7zdF+UajzA3zRvRDOqBOuz0nD614oQS1uPsNrdzhi6heGSt1Gxbr0FVICzO8
6tfZcNXZi/PaIW513tcBKqS5F/AVaTmKmM+ScdJbKv/2fmPGtzKqR+J3pUwuuC7ihxdNHQEYfO2h
U8lRtnPyCaqEZ1uPhCHP3iQkWeU7KyvJU4r+k9NKDIEx+zew/kHn6AsMmz+TfaE4TZOHVq7N5SX6
9xR0J4e7FHWSyynU7gyzs8UV+/5OCvGMWT50y8miGPZVTWfEqrU78ulbmbC6yuaNMfk7OLJB1Tuq
mAgrDeKORq3j8xk7bYcP1YcVAvZLTcT1WajSlJ/+52r+WIsY13AeRclmqux5lGIHe9s+y72W2pOD
YadIiIgyqWk1ECHSbHuFTDZhLtqvjENTf492OXNOUldg1jrnR6Vw0TrzC3HyyYtlb4HzvxJjQEb/
Ik7GjwtHBMLpEvOgrGWyldt01U1WC5HHu9MY0KqDCACWoy4ifEi604KB8n9YNX59REU3+4y6iJ+J
I6fvGBaxsBhJHHNNOLcqiHMqVSuccmIrTcJSh3vbodb2cy4hWhoLZIv1vuDFZoqqXAV/SrlXi/7K
FLzbU2gDjjO8yVIw4YkGsMql1HS/k4OsgIIwHraqjvOlEXlCxrwZroN9Rv3ZioOW3FKdPRyHh0XI
9dkdPPq1eGoi5POyGCk3NH5FtqWoYaV8Pb/fPYNCPGv8Kf/vl8B+u+VL/S1VNrfwEZE4ye1g33Ua
jYutEa7rjbEJavOXyjqNNE2qjgNtuZgahBm8E5LKJIfzCtIayB4RxL7ZcG1qHZT3l24mhayRM/Ib
Qy73o9wUHOHC7plUlqcHjS7D955XFc6siWe6kMAjw3EGn+7f+bBfqEweIecYOpeACxOp7eoOU6mE
n5Owy6VLNp3yXvosK4QwnctzZ99l+W4EpQBu8TY1qKzCRcv3CPxH5Le31DL1c0qSMBz0d8B91iGu
48VFHAUD5htv0Gd2/UppEslBaJxWx/W4q6i8vAhNgF/6rnNyq17zZyIu0zdnUE+UBN/7MYBk5tbn
cYwTRL0e+S/Y7uy5wz7ORdpQ8Ip7wc1wAEWlg+kZ2AW0xdoS47YjTS/mZPHeCnduKIVyUy6/cLqB
Sq9yuNlY62a3hMezEr8XMhd2aDD6lVN2OSPu5W4Jy6HfKrit3GVxnJSRi9CZTqa7T/U6KVL7buF4
hMME/H2fjKTZo2t8gMYgt07CYm64wTzvtkWTw9lW6pR7Qj0k6vrPbhHosJ+TaGO5P0cfC2ZpOt7U
XjG3tfIIjapD9tpDg8u9tjsZlqfqnvKHn3GIUFtFXnvGdAZm09YIVztHtTZnMsz5Wtt7NOVAijDu
IlBxe0eWwKL36iQVkVgi2xXAVrrZKpK53w8KhJqTZHB+C50Dl7CDjR7R3X4QvLH/9ywEVNbNNyBt
mCpgrV3T582FHziAP6sNp/LkWvZGtH5yG+m0JZVL8aU/yaCr9NTXhwO+2vsij3gGSwITto7WRSto
ZDxSVjgIwdLBrGjw4kO8ASZYz2NF5wteYg/9BLI0WBHZaczAE6KnjgOqeYCx6Lii36GI6BII4CVh
WWo8Z5ZqUN98djBNnjusFaT902nxfh7d+Yes1VG2jSm3r+/39arMqQvfpPEkwlaXkV1UrVUoawv6
NKOpxFC7WhvbmF/5olcLAfnXexFNjp7TFfOabapr9kVu39aQroCuPrRAyWS03x4YZKr4Jy8rNjUb
EpzoUXRtLnDHwcDRcsF4oMHSafBSXyZj9jraYoMjHE0cffI44Fod3tbIoDCU5h/wffKQjxUH3xf1
VNho1CdNuQrquKkb0HqFoh5ewIPhWm2hsGcN29JDsc2znEheiOYHCgO8Ndx3/T49iJrynikTYGJ9
ZQgnB8vIaWF5iM230BBmDCweskvUhCsI5F58HsH/lO8vBSfLZrwieTwFFWqC+O31eKWSacMaKlFq
VUiw7Lmks4ehElSXxBED5WPg6UQXKp4X+AP/jV8S0tNxxb1WE7v/Sy8FrZxVitZ8qokBR9Lea7hI
adSDMBa6rBhYElYnvmF8aQbFDSFStqL91GZzu2X1BurSTDzeanwSTgAJVTN32nv0or4UGy+sTmW6
kOh6SRAjrKaXPJCEPTWiYx2K8SKrrc3j/3a8SSxKENE1hkCPVO5zBx4J8qO/dl8wrDhb5kKQfYaE
+axjejYrd7z4K91FmFbl4jehJK6kDcX2BzNi+wF8HW5WNQQJ65qUIfB+fmqOglYP8BwLW7DbNmgs
4H90sRh5vHs1seF9lXR1ImsTY0O7H0pDpdm6g60E3iCuQX4CxFKLolL6TSgORSX9qecbXWAejEcv
kMn4evmRJj9nAVHW757MdYx3fzVObEnj9H1usDC/w51qdd9FY4T5zxkcSzOBSmq2PpMXaRNpBlsU
QX24OfUoc0Ppz3O6FEO72N1FBGe6nJGe3r1hJGe1PQWB1Zh6V17uix0d7f7rSa3mmZsffNvbg//D
46APritC1X4GAB6Q86ELkH9A4IL0n0liqyC9R4lkjc1sNJ8KiKwrNECMG5v/mMTR+wgoCLU7zsNC
lCyjkuqajTvXaAN+jEa1L1Fko0skJaxWS6FC/u3odVbId+I3DiOdONBx7HlM2NvNIoKyZDE0rydD
ANu2w0VeUumuoNkW1cUOAmPiUzCreo5giNYaugA1Shk1/xqE7QEVwLJuzNvLh7ID2rfjQVEXEGAH
CX1f9fS8bT1JBZ4Vx/u5/Uvk79MQE1Y5aZV83STw1ZPQIfUy3GdAc+B/WB+9LNslRjMe7b9YR7cj
DUyHfUIMg0CQrnuAt9pyyGadd7v0zg3Xf8/R7NGGQmBMM4w3IogUORBms5p8YxdUn/1yDRS3tv5I
rZy0ZWyyWMN/vGHJfSZSMBuokPpGVDTDO9D5dR0p/+ksWpS3ipAE7xiycURd6waIZCBBDw426eAT
cCqNgigfYP+EAmVT4LgK4B4ww6v2Pd0J6dUL6Do5zPNxEZLTjvcxWXbJFpqONZP+yZGpzLZaoV26
7myxpZCtZKec1upn0eMw94YGJrEpEkX2rNwWhnv18O0FaNQzDIJgV3cVz7h8FJAXJX49nGaL1hrr
z+KBENP2R312CJGU0G5A8pc0E0h0es8Lmcy0jnDw2IuqtkZm23gPBX/mN2VsaGsqIpi+/SuVZ0nB
0rKh3GIAm/C2PsPH9rw2Xnh59bsO3xk2x0oGctoxiiHrw4uQq1bb7W60R00JXG5bmi4NBae6pn1s
CwXxxVhQsk66oG4PU1Myd/210/ZFUiZNyXoDTsmkZqCpb14CQz2U7pnBXMwKCSaOsvJSqc4oPiWO
UAQwqTX+yYshcVhvf7sGr11+Y7Yn372n0SiCsIKmidD+1GJSq3yzYouMly+pbJDQZMwZQQzWmgxE
2QfF8L7PQYglYafYkfdTKDUEzGUNrGP5Kkj+N1B0rQgfjFrQb5CXrXFGR25Dp0Rnd7o7vGvQ4Il7
fVp1eBqokbsaVaU/vX4Y+XIXPA3PiozpNGAvR8N2cWM//WJ0MH7TUKjzrP9i5nqPrURExg/D7iBx
h6UASaQZpX80ILqyvBfMu9/v3oUyPBTuV9kYInrZHp5CNfKSIh0oxtzCWWOPmEYbpxnccPTpoSbd
+80CAVbRXZtMbeFKCzm9J9cCE9G1cDCibWWQNtn38htpzZTnqJauurCkto1RrjHJDc5SpMSQ3vwO
oGxTrBSJJ95eO5zyVqwR5HcwvFxPbbV0spNI6oYHq5ucyDBx/X+NroMjdNerPmw3rS2aMoqZYP8h
ahJr7DS60V926p0lHSNGovJZeGm7BavgLhNqsOJ21fiD9WvZZvVEckSXdEVb+wl6wtyfY+7RywMn
R+6nppiHEtngcTSVNJ52izkDNTXCYZf4ln8VJ1jms6AeXfMSzIhFnr+vTnBSog+oZmZb4Doj9Nh4
TOpVGOal3D6rUraKh+sIOPSalg1/T2lXOyf9DPFm79hd7BxnyA==
`protect end_protected

