

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IVTcVKz+qqR6KelbIxn6hKss0fyLwIejVgwej+TN1ST/vU6syUW6hxZyGugx/VRu65UT+0QU+88C
5SDN434/fA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W0uuDuJZlgdtFvYMz+doOP0vwnGc2SXfLiGH2a5FulZQF1GjNx3fjKnarWbbCm92Rksm2FFSGof4
SgtGKAeCq4Yz/Vqm5xuP6QHmdBwou49vkKDs52HUud9c3EaEYtdNlkb4+DCcueqZu76yWN8rf2DJ
ekmu+LGiL1dmyzv30tE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Da9hmR0COgf/nsNRjZU5mrjIzRjN0/ufJQ7crbPh82WrNgInUm192216ks1D/Quh1gQ5TieAOChY
26CHNdLfPPmjLAo5/cOIRsIuy2JD7JAEIDFhFO2BcC4GrUAhSArSC4/9FyqXrVJUKuDybwv0tWSf
qpHjmJw18CiVw84ne90mESBOJ0fW1ujayfbI70yaGaFjJM/DPm4Lq+TC+TFlaimxpTFNrAUzQNVF
VSkf44Zb11D7if2jaL6ua4hPGgYpPcisaJtcEYpURXS8Lw+NjmMExnMpUW39NqnMiTEPom3YBwag
JMKm6/EZOnBvVc8SljH7y69fXiGUXgw6Z6POkg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1/llP5a+sEX6Ky1I5ak8Fr3e35uMro1bXNqkrntPBRVTqUhQPFl7wfr/6Abnu74l73YggylsZJi1
1Erm6sC9oDhL9IE4pENErrDQRZHuFnl4+DlguLd11swTlNfBwauGoCBXbTtZ8+O70UI/sRzXqbZc
NDH1RywyQLhMRmSOjCU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OI4vyCtRzSCtjYNsCqL7rYkcvPw30aumOHoxNPQx0NU0Kc5/zvGo5pjE7sDqPsv0b00mAjKXUE8e
pVllo+uquegdt9Smrq3DaiQC/9hKGiZzOG1rJH9JbLcfPMXDGpwm1inP51BNgkQwocfUEAVndeWo
GE1Y28I9gt/5q5Fs/OUAX9cAh1VoS1OcnYX2wbgJSlzuLqnGWRIxOHl4+NkNkBq5Q3Xm589bPnnz
m+d2tBEPyqaCTvb13xXW7hqIf0ahuv0AQTuiClY+KmF0GjLdJTWJjDWPuRd9WYhybCp/lrgDnhAK
cnRXJnAOwP1Vgr7EPuoyVc3UkNsZTxEr3wrouw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11680)
`protect data_block
c07Y4+ePS6PnBZjEvCwNW4N1r1Ba8mnSC5OSqAYtUJ/72yn4UyZvgtt5dg/pGugjuIiCw7VvqgMp
Nxs9G47MdpsGwOHjUFc9q0D87wEw7j/Vo/yvTOgxhv3ej7g0Dottqh/vTMRLX7zB45vC0KviqIan
9DVq3AQgnBsV4mfIeU0xfkouuGd8P2OsA9tUZgLyKZjdC7GE/kcY9cBIFfBo4HdTwkNtKvXgrKpi
fxnzVAOdB2s4nytuMQIiw+gDk4pPnqzHZPghzHHSJIZDLOlK7cjuN/FgYeZExPdACHgt+Za2ldVR
NXiKpzeZgEE2aa0bd1Mdex4UzQMN4rQCUmPO+UfTrphCvMB0Ty1h3x0IU6AzWCKbq+IlwmjahQck
4ghmo4G5iOCKsq6e5mvOErtga2wT3hmb6GqPkqJLzJkgtE4qbGjbCnA+V/gQfj02LwxHt6HmYPc9
RZjmv9Klrnuv30hb7fTL8T5WACcp3ID9Yocg714Cy3eSWUjw0kaODhDtLb4xVIhXm5FNz8m46p9x
xo49bwvFzrZ9g/ALcWrlO3Piq/8/nKaU/1NwPuGwg0B05VMmtFr0pFogZHGZtXkxFJjTs2mXU8vT
QmzX9jzLP7RqrBlH72uXZf3XHosjBhBNksqWDhiv6VEnCjKP8kDHTo78VeMlAVOVyGr/zWmNTrQE
hbhMRkfcohJHGtMY5skx/CwArj0yjJHuRwtBY/fYlNGN4W3Q/i+re1YUgtMv1xaVxpIHQ2dW5gbE
FU8CxOKUwwKMybPEBoFJ2lqQMKLgoWBS71HsXKJKa48kXYd3BX7KksBVD5Wkb6CmarK8Bk/WBYe3
sUAmfRJywaBkq0B3regZB7Do+ipMlG4zDlWhUZi/IFXIXJ8uW01rO6MeuYOpCO/k/TCKGpwy2FbE
GFw8SaUW/EqTcB5n6AFXJ1u/sBR3UuPwq9TzT1lMKsUD3jW+4pFyaEYrnl+zLZJ5h2P+9OxPsliU
/bikcIAYm39B8uC1tISHp1cf4JEhDcK3BOVWSwU63Pa4sany8hIhtz9reoMNOksw3FIt4OlITso7
Ras6TPEkwVGB1oPnCDAFYyj3gbd5UK4EEOJDGvH8FmSn7goPvk09QmBtgF7puleKlWyEwOA+0qgP
HDoQP6e1wF/ELSmz/1kZP9aREqIIlIG/0+w80t6Hvj670UIh9D/uYYbXik5qUhCK4zuOsWS8D90j
MEoSB2mZsOJDJW7OIBwDYCKwzV2x7QfGZWUZSgV0wCQPko5S4HTunYH8/HSJYYPJuGI2bq6gRszR
DRhf4QiaGLi3wnrysYzYLdsI1N5LxcmWlPgcrJtnvShvOUcRF5J7ZIxuwVArt+wePEn1uZu8RzWp
7cB+FQSnyeZ7ePorierIqbhjkmRHeC0B7xk0jkvQKZKFiB5LuK0glwElc+Gaxe7IlAd8JCsjRdyg
XokJHhkOoWMzElr+9gEJpCIgKJljpbuCi9t68s4wHYLtdGLSMm9toN+ep0OkXgKHVmMNQsCR86N3
UbaxS3p12LMrSbNcYPUoGpyqKGkMlfPAhXEsPiUgHC5XIZGzp6V7pkhrn/hrzu8jIuTAKeo4pW4V
BUM7LfAQIhPc7KzunULn0991WrolK0J80Pojj2XM7V6NWDp/GFVoUOZuCwGAIcAoQ/F7g69d/pCa
8CIXO++/ZHboaz6bJgLju8bIbykDsmdF3yNubMMVGPSFW5b5XmBzPtrxfDWwtHzduebNzckA5mtj
O+ONwQXIUkCZtuRqfoSdxhLDMd/5e20QKLd5U/IJPG4WTiRVBuT4glC+h7Mcj0N2X2GhJeL+PwI/
ouIUP53CIB3Z7KiAjmOVvtU6KDVt5qX6VUUjChtFI0gYP4Xr5l4fZabcD0XmUCr/d7q76uZLO4JS
jxOXCVI675f4KQJgBnW27i5dybuLk/bTIs93xIYnQvQ4Ywoqg1oVJF9WAJZH+6o5w/ErS544yU4C
0XBNR6NohUQ9orfMSDs1MlGmPn2eGRJPGMIqjuRE7UAHX9AcUkRL3K8F9YwI/PccsJxzZo1rd+I9
4FcLOHHmjiruGu/93bsvp/xClB0IR6iI40A+ickGaiz5Ri6RT36RuDjq2gIVZkSFd0juCZRVX+7N
WoVBC9k8vTl/Vc6jE9U0iGg3puLiAcT1gbKJrXmBdgpLw0qVhMIH8Ccap5GhViH+1+jxpCEy8oQf
wnI2UJgnSI9TUQtfaBpDGUC/o8PX23sClwI5ckEVYOFE/1Kn+XUxgNGw5g45dfP9+CmLVNWAT84g
hjsHpwQAucN0ckoz56er1UbKQblORVgxzSZIWMvYD86apf6SzcwIOkYwBRKi7D8acLArB24/hLeh
jldabGb6z+OoRVmU7W7BtGwvS4TXn6oaj/4rGnKA1/LAU1+AkytvLpcdZLNEa46j5Q3RS7c6O8Xm
3MFPZjAgly1bt5lwCfHcJDm7XDu3FEql5uO2FvtNFMfAciv6oWjchTSUSeelIfrGhh2BuudFbL/g
c8DdeLx6zwVO/Y79uVSZ8LSmE9VG2ha9gmbGqdz6xZaxdPaLSrHfwlQRj2h6366cbx8T3N13UBnY
3YAvNZbSPolHg468FyFfh3DEtnVCpHUnknoE1/Jag5ifS7vklg8TqeBQQlTCisPVOBJOJGW5qRhx
5DHwchnzCYj+hHTWOfo62JJyapkgcPBFhQIiVqp7pJ3jU3zoOLthHt27y49L3r3ZY4IAh5ywXqyT
nfSpVT7rMzX1P428oRc7XTiWDiWshiqvrqlOmLhOqd9OfF9tSUzHVoWvsyNq7Ov2zom8oT5pL67A
8g6TEkGaOIDfMFfhmPBsv87LUFyQJ9dI9fJ7vWcofm6k7orVKUiiEPlVbtIoYMjnwlPSnnUbbr0X
LriGaMuMZcnrpYQpYKtOjWEz4HKANewODxQwC1E7zlR4YvnVDe3WjBbFv9/VOs+TGVMhO4b2++Ls
WFAH3eNHaTHQ+1oyq9sYQZQprlMtbrGnwOWkqRNqO92/SNPQ5UBwhKOUIgeoX5kiUWoqPFIMdt0s
XiK0XqYyU/BBBcw225bwrfQGtTax30fZrqcV/Xk9mWxhwBtvV7CTiLJtLovyAir2ZITH5RU+pp2D
8xfcIngWsFGuopcpKN4NN7uvCA2JBUkkIB0VB0P/hsNrhN8lbwSoToYGpW/YsO/AloeVrYTtJSK9
5fbsO9IjykFvrRluugFf2Tn3Cg9apO0sTKLZjOmK0AJqytCam5kuPNXEJz/Blw0kEON7m0Hv10NC
BtGmaWYXL7D9dGuCwwuoBGNCCxWQTmVrK/jbLCqR6WK57blnxs5sL2ry84n/rIe6i9t+7BWr8dkh
E1H0yuN+AjpvsA/+O5D5quM8oB5SCdQdpK0HrFICYHJeCH9rDfRBNCqE0/gdiBec8CrLNWuxVi+E
FCJ4P3lk8v8/0A5eEeDp5PbrkELZb7sUF9bRvJ6oR69dts7C3HbSRX4vC43PqXGc4W/EENTbiExu
gQLK1dxSTfSlXw23HnQTHqryRt2mL+YxAIdIo3HVo/eoiPhiS5gnC8g4TICn2OlgAdoL/UiwVPPQ
eAdWlxRHoDn9BfsyQ6xqhC1ZSV5/y00G0l6FiaT8DZv+W/h5Z1gdf1CQ9pCUJEiO1SqSTzSWsLq/
7nZ0vtU0WkXibc5XeA7s46olLVS08oYyYoT/WWQ6vFsGjzX8g3olXW7928qdS9iT+Hgm7+zql0WA
MOme0j5xlrLg7VchQZfVnfDw2Zx1ulTKZNmbknXKUzSZQlyjyK0puX6xVQwKGBoqE1vygAOW8d2E
4aO580IvEOA2No/VOu86bAON3Wh3Sca1iksPLFLk8VR8sjK7SBGBoFNyn921kyTEKAuiJliGRVVO
g+Nz9kpgfR1zPFmTwAD7+7olDBcRbr5L252VYBdfG6o1TVRf1CVk6tWKw5Ah8/WIutW2nZW2T9ZF
VB+jr19Hu7urhPIPeygYdi9bxr0w9pWGL8b4/knTzxi7N7wHOq6wWozbD7aTEvN15Fh48bpHEvKP
ORF5Ri6c9R6eWECsvekMB41KYV3WXVMpxaesLfIbHBDTHg54exPkjPJ4fOltpYADHaHOR+LXjJK7
Eb0bSM4zpk0pLEEvdik/rj5PQOnTUWffuxjGnSUQqyOFEIZDeHovEof1XzSDrWi0hXGAiWIeOTVb
I8EMHku47cX/gcTIh2Fs1bgTPc7vqBE7vkC2uuQU6AoKYMukWpTmAVfmtgEZ7lxPNd8s80BX7Q/Y
PCK5wdz5mGJdECI8zNBJIImWF0E2wZEn6WfliL/6rTBY5ijXXaCFzqafKKDfWxGdwrgwPGNmY9u2
hEqN3Tpnnh2197Z/1H1t5tI2CSHA78FPLUzH8mC2IAwHsP7p6PRJsLigvEaQnI4R2t+B+SiFtj/R
489oNCU4eK3ExK4Xd4xIJ8Ga2t2CPT2BFmfB+V3Jijlwo5m1lt+1QxXsm4TtrPuv8xz+llGVUBli
2gnKAyYF4Wtp62J2zz8NOkLWbQ6/iTogpXz4a5Y9rwObBYkFAz+hIoG8RlwAxv+T25/Js7r7Omq2
yR+R4egkwCIru/S6pJhkBO2mGMSSXIKTr5+9X2cJUfe+YTHTAuRt/ziSLCWaNYrE/FDpKGyfrSaz
FC4a2bmBnA7JA+Ce8WxM3UyYqU4kEEdRPOmNLfPHBcmr6WBfwLIxbvj01+z9K1HkbyZI2YK5rOh+
eCzVJbcA/RCD3L4ofEn0ZHnwsICbd3sK3d3/3tx9JLdluLLrp1Q9tM9jcLMZkeJM2p0vxjyWe523
oXRvZqD9IRewlRZWD8QH5BrJJATVqq2LJCgQZ72ua5xy0s3QbDUsj0LButUq7nuFmreDtBHXq2eO
G64RgOWRlQ5xDPlvBsx/ieQlZB0ne42f6mo8GRBC96pEuTXyJaqfVAqrcWWF/QC5/LYvQNoYPee6
RRahnrf1L404NPwHa9EW8VRHeBXr//t1s3BdVVNXWXsOkDwmfLJmZ3vCxch2eHfJTTHplhxmeUZI
5/OHV1Sm4468B2wmEGI9AVITEPbEq0ZcTLpED0YgLpSog6XPb5djp3towRn3FHQJyJ+n0TAJrgR6
3uYsMjhkpht30+GbBE6Uf0jaX8AVSC/RtWPZ8i1crjmTbSDAJ/fsnakBfuLDxxgtZxfxOmATE83c
2MQyKEvPuckcmDoAsFxfAGblnHwh3Y8f0wpXfzETjiuKCg5xc+5uTZr2Eo0I9ZxtjDguPnaJmmLf
XwfcxqN4a2h3iqf3VV7oQ6OmzdXwHJBm6C76Dp13W9Hire6kdXDGD0NUoUtRRKAMfDsdCtf7YKCn
MxkmxR19pFGqNTlMRNRjF9cgYQ9ueZ/49x7PYlP5+nZ9LChaEe4bwRW+KS2cOgjszXsixQjHlzz/
epTRWUiPytiKS3LNNe3ObWEj1cwnQjjRg8x4nuSIF7JfJBNU2uwrWeiLa9Lsczn+rCcsQAxo1Ttz
3jkxsMGbqJIADZJYWoPvrKkNCWk1hXshSnL7KYJmb8SIFsW4OOEz88njzOtNmC4dDPVVCpPaPJe8
Lm0UtjIYS031Tzat7uqaeHJzeaU7wvirkqatm146fwbtugAqcpJlf3Eec+gIsQHaOrY5M7tTNTa4
iYX38aDTFBzP5t5d8t5eshqijR4dN9lMYqq+qurkF8O/b749V6MswZjdbkTmw4Xur2uliDub+XLA
Q7ue6FqSUnt1Q0deSmSjIM5TbibcL1XBRespr9SM8HqHdSz37vgHn07aQ8Nx8nSmPfsDv40Z3ZUh
qGhT4YQSFuS7VAfq1TyYb256qLr8a2Idoob96g4qnWo1yPuKqui3iIlK9fUiRzS6lzpOT5HNmDVV
1rMq1L+TqhhMdot61R2brq+VNR5oxThhr2dciKFuliBwFy/Wv9/ex0ZpwGVHtGn9Sv+cwn/SRu6k
6VBfO4Yv4iQxuBCOxHF8wsC5dN2trWhhb1MnmJNutXprYNQuLubJQbG+eODcKUz+sk5huvA8dTYz
e0tC+z6sD7LEumx8gfmNR98iSAtWKWLJLlI1f1pXCvShgHwoIMwCKVw3aOGKti/+NZw7fCQMpuzB
IFx4h/ROJoXF/DmQ3NYeydtnFPcl2fOVnH/GjZdHAywmuYJx9Oda200YSlNmS4K2gXw8Vo6fdm9i
tvEaaPbCfLgztOK1A7HvZWb6KWr2xqaW1I4Cqd80w8qhuGDFjsj7aWnCJIJVa8IBJVjFdWonfSgY
nVBze1uG4MGjp6D3u5czVha1J60dIOo5MlNQMG69W45Yuv51ah3wm4CoFQiuy8H+Sjd0TqgzGN9s
UszyA7pqjIMWEPoN7TqUgu6YDVnv9/ZfWUgUu0WG2XnNZPKqs3jNeke+ePXNHOmfo4TEw9YNCa3t
kHmbNB/UdzurAoBetWzJWWkBktILAdM2pcY/Gj3QZxBnUwA/XpKUOZhytWA+brEBLUA5G/KrtkVf
uH75LyXdtR6+EPlBHfJ2tRZDpjXEZm1G37DQbTCLoyoezNoeWTgQcA5g5s9VREnYGusgYoknQEDq
t69RHsMrF0VwToi73POak1QoWyoCfHrG2JjYJyuKUnKyw4/7cKHTBnpbSyMS/cIFx0j/0GKi8Zz2
vVi1k3htpwZHQ0ZGbu0D2IIpNnvag4w2O1N0beNJt+MX9xHND52plv7FMIs49idtfiSFpGeXQi/z
mjpzpMEV+jRQyWG5dgMvLceQv0wtKzbnrPes4yexDK558vULD44rJkkmeeqTdGSSwcM+g6Ev9W0Y
YE9jcY3lKng814ba0h1Hxd6C86NdyYAVJnqlNlBcqxFxMwdySSEfu6paTYHoWcMcxcV/BSR47bSl
CmKFUxeUQ9aZkSNDDbv2lYW/INlsOOGEAODvZoatOFgjxPGHo/jJDnMPtNvCuCKv5jFt/BfGMOO8
oN34inamAiZaEmZGtKvHtOzK8beGYPXFYkhvtz/c0RYUFR557fwhH2sn/8HSlFnFCCM6EscWbgS9
YOBSiUIHNW11shNPmy9X8G1rNeY4msu+PZrHP8X9BhdSVoN2HCjN4t1oj3uHUA8/znpFL3fDpGZr
YMEbp/UirJyMfE7vwKOWKDGXWJmh4QAiHunvgSM0xY3JzsRRl/3aj79Cmf/seUHqwRcJtFbUG6fl
CUEVH0cdfuwuFa3E2Cq70QnLknSVYYXP6N6LSHKTVeN2Ux97V0JK8P3jXG7qRXbY/lRbkh/fOr+y
paZ9tXFmZmxW6LMH7pLf97WK5A7UYuCmT6JUoAAhZ8n+8cFCl/RuxRtWquMJbw0M0PJEJcD+31At
y/cJRApOKLI8Ip6xMbnaiJ42YO4k5RFIdP/HNk/3fmNC+n69QDRVDvDV56aIfIBAOo3lDVCylRQs
IpUJUaCa6XlWVUklFRZann/W17vKNyJx6NhXymLnIl76qOWWDqTx6pISNfcbPvZBCEY7VW2kzHxw
FPyVaLqql7uhTGdGnMz98JrFBiRfQvAm4NZ22JVmaC0Ff3MC3Ya1+XpbR/fyiqU05WdQifTDeEXQ
8rajKbN4a7LtTHuC27dqu4y2pmFUEBa5uNqZNhF2s3Z7Lc+1Hja1rV4NugqXJHUDg+8XmAnkXpa6
LedxOOKm3TusfTjjblzsDW070VwGxc3FpS7NI4Z49fMv7SJt0MGOaoOWFN7+ER4XqugATEkydkmO
g7Min1OFV0tjj5udkMSpiGuRG00wPd2vF1thLkH1pRw7LstZ7vJnyzO2dQf/2ORTZZkLW3M6OiEU
5XyodQttuOEr+De1KFzQM6NZJQOOpa+nuPOdG8c7qbdM2/DixBGB5vYS5JoCXfHj91+NNOCSIl1U
ALq8Y29kJGCQM/4T6miR6+uqbnPT63qOgV3JZNukAV2JEdXOfm3oztn0bwmyo6qNTM05dnU0fNqq
1l/B3D1Av/AIVU3cD4aOLPhiwYG3xUKDrbj+CBdN09JNDrShZTzKIQPsgGWc1rsiQoyNaTi56jZE
XnH9GXb/sRLFukk04ABTTZafV8wHhxW+T5fRgvGP1BFPXZrPoklqPeErkkz3qYJZN22D4lDWzJqV
k99Z5Bi7kEBBvihAkMM1kefUvW/Zbws4nWQsd0YkHpE8+FnuEH3g6WQRA1WRfN8Q8DmFzDWrgbfn
g48tGJN1nPt//NJNUyP/TrNMbtLYc2iB8nLfxvtWG0RJGuNzOleoFpeF0VGszlFoFZB51VxbPf2l
/E+/Up1YNlUJq9YseRFQFLD4OmNDAvGPqyNKdI0tCLXOofI9l0Z5PDgO+uiwAvXzywUk9JP+J645
mMMbrxsOqOlITNblgjL9hhK7driqKoWg0ZNduhn3pCdqpkh0OM4Npb08ZDUznv3QYDL/IMwzmBrs
ifO4ERDsWdEpofEoFHTLe1FlfEs6HM1+qOxcj8tlUhNIRY3i0Za6XKydY5PMX6ZEoIceZPP4Xlhn
8yZRE7QZVqItgxfZhgOYP6himA44zNCsewiWb+ixDnWTIMTg1VdkNoSOhaIIkxiYpNKkqAj/+sKS
nZPV8wzRs+c2QgBBmHOcR4Yf0RCoZlxVVNUsNM5S07+FspexKxlcCq+onploctOTNNh7NGdF2aH2
U6NtFwpn7pYROJe3rgork6Nr+pYuR4qJ/SLCZbKqnOznQ4G1hEQV3kqnRBqJxRr/9keOqck+QkCT
JZn1nc6XfB7NML8va6cvUo0Z3Kmj617f7rUkHhV025Pd2a3+pSM/vpRJYd3oSGt4/B8PAkb3RReH
psUVbuqCtirP4uJTOjRtOmQc2QLDXxa3Mbz+UfetpTNBMcy/JqgOQRnVBRpE/bsaJ0ge9nuVNW4C
ezcI8lK5FDfwQHWPncrI2B9D460z4d5zGPSABNNS/c5Ly0Nkz813eG7LXVJ9t+i9vK3ZVrU2mG9u
WEAsP+3QyaRpYJ9rcNlhMZFljjmSX9+AnZE4TZpBIbbhKYUyRvI6OxLnWBMp0iD/m/SaBio2WU3S
OLOx6vaSPyAj514InMPtJpwb1cLSNQWjEuPeNaK7oe1xCYUi+UnsIvNK+EtQytjfAUC9sVzyxOQQ
v2Qbh5PeVDP3tQVUWRDcnAUgQ7mBNcdpthOA2lyZVD8OJWVujOuirkTRNTiLx0icFn579NCNdt4b
0h7lQy4mrfmO8YPxlEgLdETJd50OJ49O5KF63DFzXB8A3gE8rC8104Xuf7JGNXjYM28LPYO8y615
BCWV0ETt1Kf4qtSuKSTjHE+hWNoPtKbcIPp1jY+kBr/7gJB/ugoEZbHvwByXQj2E1p38PRo+nruH
LUrU/gFSAcP2rKh1XvbnA5cKP99cGh3CzkqlboF8S30DlRMJUENn66V5P+BD+VDcIOAam/rwTQCB
ubysVCYZxmT66XLSrr87ir2dNlipcKhkuTO0irNZcgqZLKeKfKbdiycbXzwG7213h6DdOi7Ss9Ag
vS+5qQ75Ieqh/QIx1kGl4HddBVo9ZPEVvlppJpzHSWk2HaL9tvMO0BQ2VZvjM+pV6cOJ3moJV17O
esuO6jBvRSQsLOmkDykrSWAGUxxnIr5EGNUrBrS/KRUi0722V+8M7Zm7YsAM30MHiyTpAYDilcbL
P+Kyb+O+vvy2IebIlgusxPREI3zHMpCom2tXtuLD3JsLGES0+L4qCKC6Gmb/d/MWrWDLLSBwe4RB
k9OBA/I6Shy+1NY3mAgG8BpobDpTcoavEFwLf0YNohOKpVgeKETEm+7Gkrn4vTNBJG8M9Mo6NU6x
fuQJeej2wPBuE9xh0JOWyz0HgWSEXOlMDSEjigS2TLdEGivV8xrxoghmIlmmzwjAT/NhR5CD39t7
y9edYfDRrYT0VQWvWLTfdLu+JTaQArKXpM4A6E0G0qm4BEeilXHyEjBS94Mb0G2C9cHhF08Sz3Jq
KCGoBNLatchc4VE+b9X7ROpQ2JhIaQ6yeaIwx6H5ec48Kk0UrSacwVez/fe8jodmHO66DHVk1Ok8
NTBkH5FBliDVQ2ukVOLEYSxWD4Fx7D74hxazmlQVU3dVl8AF4VS1s3zH3Uz/jaCwOWLWeXk+fE+G
y3u19PhTPkCcdu01dsZmbLVO6kOby6+h+aHVTuFgb4caezLbfNdEok0hRjrMmAja+EfHUlSOXdtr
rG7P+4z5KODyhDYhr4Re2jk9wCdOOnsrUW1h1pLVWwY+o/xKqr3rFzU5xyZ/2/us6avgFnR5ugQU
B57FP0uNgIsH5d9PrGGZqUt8ZnQoiwjbmvFGkCqPTh7ei576sreaWsAN9hzr/sPC4qMdWyOoXLxN
m16bVrZPv9orXV7MFldTZ41RonPu/7NpTbBlIpDjnPhEraR8xB68hXFb0u32x1Pql+HYucq2KVby
NNo4kRMHe3UPzEpRG/Ugocldsn65DfxQvSDgDla58D3Z/hfzMlOc2b/hGix9hElJS/1Xt1g8ez6v
Pj9PuZ7f6F0KvmIh5Sg/omHbD7aEH8a7RN4vS6ZN8ZuAH7fKT6dydR3krWFypAK+AEb9WTpicDG0
ayBTOV0RylGTU9lHBAXvKILcRCpiXBfroWq2feCgzfi+DEpkcVBDTKsIH7/SAsrCSAsMN8P2hp/K
V162RrXQRNfYwStuDptHudi4TLuc1ahiHPYqdkwa5PxvWuJsFh0P/JSqB1320uhtGAyLLrCmnDqL
uHYMfHKTWb+kBSljAe2WfdkL9UNkuVUAlUIIgFPrzDQcelztkbmYHRLT3vys5aeUPWhlDrHzqNCO
Y5/ekfaijs/7XD+DwGK+woWwSUlpfN23vDhW/5zhAHsde8zncKviM/djC5q3APU9FI3qNlbkpzy+
dCoGNZ9Ty9XnrQXJ5mbtZP6YE0ThUSr/7RtRoZEShQOh75YIlhVQp99GBQuCHjVLieh2EeN5O0xG
sWZ4C75UX7ieQSLllkItkmgWD/YuiAwb54HfWDF1xi3YSkg2M68sFuIOJpebIzv0F0Lq2mWPU5h4
hhqvjzlhUX0TypUi8lx1zRR1tTvucs8ILKxZ6hTcVl16gwtEmeHZdQ2rfJSO/LS55VYLWWOD8APo
MAE1GSss5egm8ZYnfQXNaW6F5apm64LGDaTVsOivOtk//JIc78XZQywFT319cQGciBWtyo1uwg7K
z36dh8UNBOLSWY74QZnKgNqdqltplV32fK8dSv0W25Om+CUPA1zOEKyQBx+L58QoLgfSh+AhICYD
AFP/IQ92XEKpyc4Y0nPUgB0UTTaYpmuI9ozGDfQSUGOWX1rtGg9FWRwHlLMMmppFlI/cDaRs4/Fh
GGngJYgTjzJurragjyzBn18TaaKfdoM02stJbFxxkUVjKC9G3UxmJZAJ8s3NSScUQsA4eW4SlQKH
F1Anbeqy1zlFwlwGEiTXDqK2lJohzZ9IZMRMf7kagkQCt1n728rOwmMNa9InUmZyQ3ts9uHNtqSh
8ZlUenxgFBsCbfeIy8N1UGxWgQDuQ/IiObIYVrNKub6EYbvw7m5YLX+UyWZA1tU6JRZV2W8I/Ciy
caJDe0PUrqcuV7M9Gp7dZ+Gp2b3dNEiGUoQsasHBGWhusZg0r01KXcyIUvUPTlid+ER7iMkZ8pCf
JZraTf4dVGjKkBI7IES5UISzo1IVVxN+3STOl16zpx7bhz5srpLDqoQqA3UsE22LytaqU6x0tnr7
kEQeRcn/1OQxZarzRNZdcfBSSmNU8a57g3UDKRfCuVRymXurfDHQtt+eALljk+DiB4JDyXT2BJyW
ID6TOOjWsSFF2OBS5IdjkvRY9bY87oee7h/VSVWztzsKbhAGwqV5yQP2yP0xLcN0R+V1S62F2TZX
P8wucy6hJQ3ikFtakc+Hxj+LpIkgZrFBI4v655AFn3Gb1UeXOOia5k51THN2EUmaMT6C/QYmd8Mj
qc78tXL9AjKfU5CKFdcO3wk71knq4GmxMc+W29OWsOJRba9cNJIGFrNy2wLDdKOGwaxzXrs+rT3d
kR++f4vF/CqI78j1DVxLSBEyj0pivP4i7Nho6Md1BBgX34md39zRju1VzIoWirMqMhhgPZV0V7cS
GnvBOvAfeSrKBr18tLrLcLIDR18jx+ExnvNum459HF3kpNaS3Ws3daKDWo6tdTxAqoKG12JpqLLq
2Rw2rfVZLbIXeZ92YCojFg7T4H3bDWRQcqLe/jC3vNESksjcS5r81qe4EIyzhXPtzTo2MJCkVBhH
gqbpE/dyDe4Fjagse00gb0hQ1+kWZDHdPJ22N++b6s+T1C58xdxTRTavF1zoJPsH1szfCw450Vft
0rwT4YSc0H5mIZBRwBF1dBKiCS0hjgFb4nDgcMlWVcga0/wmZIdq11H2BYmCARamwrRW18e/GN4h
VIdHOSACOFbhPvHAqh/O7IghhrD/PNvB56qz8P0hKIKZroolRLFoPALwiB9jumwWcNL6SAaFduWe
bE+ISXQXS7vsXeBbYnTdeD55iaRHMV3UvqWZia0x6xxzFY9mQcmTRGycH4Vw+Y9eGohUrjicELVn
cebFGruRL2+bjVsXm5YYaZ5flK95Ph9dmhPdyX8HDc+0+xY/DAUDdHYNZ9cynphVtdLzwcBbBvMh
kj78lkUtkHRK0ZRygU4/0ZChjcF4F6JGjSxzqWJqGu065I4UwPwlQRJrOBdyvyIqRn7hkeGZFkfx
H4pzIW5izVNANneE39Lhe2XPSr6cCbKe7EDwHmXiHdkMf/ypGK2wGCI6lfqIZONEjBFh72ypAtFh
xqoY6scbHQs9RmbL7cRqzXjX+UmROYNRZP1Rl4CA9p0brM2ZofhPOvdjgAU5kHLPpbrg7yl/y57K
/6OLy0oyt6rRwgr1hynAnMkfq9diuJI3nLFaY+2PCxCnGiBM3WWdcKuqToUyExvO+rkq+S5/Hp3G
URSbQqzmVbdWmYchwMFfc3wphxhLAFch7gWU41BCckRCt/5mQG2L8hRtSgCvfDnfomStZqEKFApZ
V/bMC0j4AUKvFxEQDnO5KPsRAHbQKrD+GMSqqYt+28dr1xk70K5T9032gjjCSrI0cMe0Vubm2IS3
cF02dC5l6QaiglatKI7NRkv/b0mgp7ry8tyxMty5Ga9lRu8NHFw6TPQSAv1h/6xfNBJ2prsJXzDp
x9qmJ47OvuB+REPpPhMgGR6aqsIwYjogpJpbIoHctCeKOhQbeXX0KzqV6ErOt/n14HH6K/5bNxb5
vI0OmxlbLu6RBUhW2JznSr2tV/tn7N5DB4f23/SDERErMWB/jcrDFCteUq52e/TuGxsmTwz4cjAf
hNdZzFyIqafzw4KlIPuxly/QPVioK+dZ9XK2hftmz4CVscf7e3BREhRtDIT3T0wliooIuuHJSRUO
QW71y3idl+8TPkf0qI3an6LYlMGM8uhBSxIPUl1AxP/2G2PbzYyQWrCuaxjtn04nRy95Ul2IazoE
ikqR8lWTQCYJ/PDvVECc7vkqaAWQ3vrGH5AZoxKfU8Wy/8mmdAm/2iC9sEza/Wgi7hG1ylOPMR4v
uELi8Aq9wtipjRWcdUTrlT05LSEcp+8JoivfdFGthh6OGi3ESJTk9Mq+U0KLEFcKke1PbsDlLhc5
yJ+ptab3nkVd9bRURDUBlG4AYXOkQZ5aGWEajrgpb7miU4IDxwySYfN9ssi7NsvhvtO3Pv6lpMXI
KUqAYE/aSmdzRf4RumsHM6MXZEk/TxKt9H5+3xLLJYIz1XzoqYa0mrixxPQYei9+Uksxa8w1Zq81
6SrxFtimgW2WdB20uoh7h7Gvpl7ZUJDQFyagTJRVy5ZdFfZljuPm2s2MEZjds8M+lLyUmTxm/uT4
KkSl4OElNKRS0m0Mc2Y1u8Nt/uzbaDT7ozyPdNoyuNE+C/iEKEAiD6vBgr8XAKkqHg5GZ2gp8bo/
3hKxvlFQu4zrMO9EWBj1tdytIcqEm6aYOb1zTYbZfv5UKi+pTHGYtacFgoj3gkZQHV6Do0K9Hlgu
hInTpzhw5A5SY3xDWIqkhdMS/mncovYJqWKf60BX7pJldhO4ciBzFzEtwAFFqaW3zY/uIJxdCVbj
HPH/wIcDotgznd7iBkJY/N8vMpDF4CG2mf2ctux2S/TGzYBh3oeq1toa87I+ifMowlY657pJmvbB
wKzr8cMFwaWw+4k+sSsxgAnbx8g3MXZEomJ3+RxCPni+HYQ4mOWx6DYsKMz3kSFK0581x/gxl6va
JmKMAj4HCPl4a6uUQ7D/POHuLA4i4RFO6n7KQtk2c3UtLvif7KcNCOBz0bxFIo6oJTSvV3oWQ2gS
Rvqb2rw/xUdhEkLi0Q3R9qKW+VXKZy4iGvk9JsYUT45CuS5d4IDZ6PdixKe6KRSp0uIQgg6JbCE5
jEalF5YEajLONfwf04Yhdub7eDQaoxu4Wllsee/auM2W+Wxe0w0hokDD+keuN56BDR7sRLgwfcWE
w+cFIlX9FjTzl4UNNPjoaTa9aVSrau+s3YGTXbtczfvu31oaM3g7CcZaw565ZwFLawD+JX6xPIjU
BFunYtH6Oa3/kDwfQmqumslkM3W3ggMmLsrbLkofjCNYyFlPqmZPfIb/UrTtWJfRI2/xynytcD/D
/GoQJv3AVfcMx0RrkYOermRiyy+E0Pgo/hlji3LAIKDPdij6s4TrPWECXAEM1YFjMJUJnwqmCETe
+jOPB7CXMBe98sg5bBH2xuKGAAW6MqQjAekk9T3dWRWTKVxjOMvxShLC0SebppD0IL4E1u60IeAX
SbiHilX7NscXzN0zncFYonOwx9J8Cu1XR0UOD55cA6GRB7H3DvCy9sOBHD1CxTg6degeGceLJ72s
BPi+64EQP1nAPx+jVEX6APlm2sy/oSrxJfF21TgbuV9hv3+ea4UIzTIJw1OLJgLhc7dBwKtCZsoG
/ojR446x22F5NnI7+i3kcSGsqe/2Nm+rRzyPF3vvH40YhbUloY1qe+PKojcMifI5kADwVXBNs8Ei
S+pBINl+nKN869bwkZomp8Tkp8WE5E/ntjta5ZaGntGryFzxE/K84Tm2coPl+xWqVaNrHoRHdbW0
bGecC+vBL9LOTpjDonDNfOycf7l26jChAkFWXeYoduqGnA89O2NAobuxDKkNU6KAk21CW2xIRrhH
eQ3qv+4ZPljKQ3WYIBTK9kj6gtAV0Suk3QKQRMGy0XXfA6UVx+qJfDAJ69treB/Hip8w+GmjO5rQ
4LydQJhMFFg8kvaEgsdQHMjM7A0X3Y226ZhraPjb9r/kPc/x2bNhEmgkPw/JdSDDOInd0OvZ+za5
BU7c7Dyht3fC2Cml5JBR+6CuTfwSaVsoBY9VC2GdpDtb641J1ucvFAtlmtTgUUszbRkhuifvZrXR
n1f20Q3dFS0kVb0QiwKvenIdG0sc4I6blkOLfm02tvB42GpUaSq0aQrrq3LpYqyqQfp/wKsiG9Ak
zw+Ht6wVkKnpf1yvK234ELPtXLS2sXQFPI5qfYG0wD32xJ1wFV9AoBkwTwePGnm4EzXxF7UGY3Yk
3KnTctgfe8J/5NZVuVZWW66F1mmGbxI27uRFnzDIQw0bweFzXyFKhmcdQK1NoCJJDmoYcJE/0mL3
Q7KHoIGqtKa8QJGb29KyE8JTEQrh5YspI68tR37K+sJGPn1+JbQs1kXY8AsaAcVH+vJx/Q==
`protect end_protected

