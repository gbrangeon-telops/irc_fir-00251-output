

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bdlZLEAewQqpv1o7OoBr4R377V8Hk5Fd8+q/Az6G9nxroFaOnD3V9+lWQZaiTQ+UR8tYlBixiDT3
2rrbvlUYqg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PNj5XhRRPylbuLUnq16m36512+Iu+tuxUNOB5vui/U9Vyxliy5LDYUjGyTrkosJ5RLmSfgYfmdaq
x3GXyG6MVOiZo15XiDmGz5Xa3WMM3TuUhfpzNItvR+cjVJcfSX1Vpo9/m4Gf2HbgWDY8/uge9Yz+
pdDWTg9IqOS1f9m0bhc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tfy6e9ewB1av8IAVBQg5F0wJVpezM47U5T38niEmKqoHE2EAQIsVtLXdGuC0EVCv8iR27vcg17Oa
mBfBXWB60tzPu8Q6DSJi1RmV8OgW+NgUvCiTMpLKqqsw6FnhMEK3lQVXfOtnfyh9msybPw9byzXC
dambJMmCpKtH2TBazWP4yb5ww1Nsz/1jL5i1zPiiJqwiUek+yJBHinlLsKOdmxiEOjEIxiuXMNyg
LMJzb839xkVhlMYTWXZYlSQVwwm/sLGnZ2Znntlf9sYBoE6D2vYri/PUGcfI5TqvvhrwG3MMHoTN
rPYZvU5TTqkZ0UHzprP9ZbAAvBMMlhHGjyKLgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
enscaK3Um9KpWwQm1hA2XwO16XJLOAeYZ3URNnasJSAORmdXiuv1QgNvxstTqRmJdf6aiVcX+SBW
QAS4XOQmaHblVVCTrTFxq+i8/M/uWIiPlKdwfgcbq6W9GDVZEH2g71B4sNE7sbY88daOW+dsFMn8
evKdCCrOhrfApxD2w7E=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qn8TdDpu0TmAhfXr6OjdWoz6rfyBW7fFZKyqPOjjqWteCvm3OM0JlharuS1oWtO6vCpto2FAzG/S
BlRFnD+qM3W558gotDG5xKLXH54U8vJ9P7HSKDrDRZfcvgzYnDlLOZYqIhF3QcOp7QlIfdgIFJFF
P1RDJ8d43uSYKR66QV0gPXuT19+tneyhi0YpcaupqD9/Z/vQdGHiorXfqzI+zmAX5/7dF89mvr3v
Pvp32AibqOZJekU7QCnp4VkIAFQi2sNR2R1SirejbeSwa+gfCdYZC/MT0OFTfQjM0uxBSK/I4IyT
gWZgfuPijqASxDrsrURmKezc4hgCDujIExBWaQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21952)
`protect data_block
6JDzhlGpfSblxEbiwKj2vilo1AWoaI2h7nCZAf6BC2iQnLdeJiFCj3FnAgB79+jhgFYzwsKUah1t
tZbzmx1Woi+iBY9Kth8pD0X2clOY5RCYLmzSSDGVUlHd+pmxEfzho5iilofPNxEimUOP/67aZvN4
SiOuayKQ8nhmu+TyFoMIJzHWlnJqx20fHR+T8NYtgLgEQkDRuA17E99xXIn2EPbJD/XpzefTXxp4
cfCGOLMexDLKYwDQJQJ+JECtQS9VArdOP2HIOwguVKgJ9TM48q+VvhCxfK+382erOsTV2uNSbZT+
lXJ4oWcB34WkNK1BAnZqbyk+mwnYPU4o+U4iF/72uQmRpKmfimgCnV/ZusS2z5NxxGRUqydEH7Av
vxc68VYkgONLtC4hn2AaZ+xc9qzSJyJ0bVJNQucL4ca2xRUYl/D0nx+kA/MmDbomGkhZE+in7GST
YowjFl+3HHXO5ZwemAUbgKWUtizeMFm0vsxYZexo8hATrXv72VkNbiCTkxXF3HHSm7laldIs+hTL
U0satAW6bJzA6xI6o7XFkPlbfAVxs69eZnPC1/42YwjLeIQhamsN1/Qj4UD/GEcUqLoQrtR/SbzL
cE8fpHjcIElxMadSMnodstEmP3W7sCL11/lTO7QbxqNRw12QU3C2dkCbbpDUfrmlHPy/F1vtxmoH
oUBHQvsImDCXoWTj32JX9VlGpKDLFI9cvFdvrOeAbPW0XFQ2PHTF0tHvV1wIRtysGB5GoYEOADf5
GJXVvVV+hU7DV2yQQYmOEvHtbwgkjBO0LqWQXqoOFm75VxuCU9faM3Mke0+5tH99/Zj5vABOfs1a
kW7FaFplqHIiLVhquvAi8Zud31LtwyZKgAGwH2sxO2VmEc0H5ALjPPT+r/hT5Nc7JEqqKAmOdCgs
7LFo7/n7fEEdN6hhqiA+YVnNoz4aOE+OOqMau3kuyNtvsXpwv/wm8flmHY/vB/U8hmAPrjBoQmHl
iw1GsWqVe0BKmnNI/s16qNdVRlTMX05cr47zWc+MwRiXXbHfHjViQ7nMZuAzwFYPp7dlOpSgYQSI
eLRUbau1LaQT8E2L0Nxqfkr28DH8Au4d99eqVBmIRRHHKn+KwM3nyWEMzpuYX78TtC3ZEEBBjaV4
q2jS6aK+wv44RlkPmar2UD1tiVt4qc9/hjEGaFyJ1ici12BBmns6TESHhqMuuHxkWXTaAz4tbFA3
SUdtRUdkFIZcFbqbVD0HYKH9CLu0LYDZA1J/BF1IpwY3ZTPg1AmdwczqUacb3X3gc436nrIHZRht
/ntMY1nz2GhCK6CUHyWhSHP/P0McOxyXb7K4ycitiFnB9/xhPKYEWH192SKKXRmSJNv9h6x0ADLl
K6aKRArfkk695BlN6QLNwbBSziyec6kZxvwJUvNEmJ/2Ur+XTTxl4SopOpdBA9zebz83o+J5/pEo
jeliXjJetfVUlDHYhsN0lfS8bMeHneFjYrsbT3pUsQSoP4wGzBKi14kbb+4SqF1moO3ZkO0QpSaL
crtm73Cx2R1jjcvkW7XtqRRW4EMMQY+PIDTF5vAtE/aU9wmSm/m9IbVa4xY66L/4+xwP7XUY8803
bFVYduaHifyycOpxp2VaY640HjcKlYj6datd+MHlI8KY0H0bgwOBhKv0+v3x/y0WwhPPmMKuTYdO
Dtq71r8EGGBeh6suEM/CPFhhBoqs0lATwmJNAjPKZwusRutjqLgnqZzVgnCR1wVFy2HKXfVIVhyg
HLY4NIZZte5QggdBbcuuNLNxBzxLyLkvfEZ7VuaB+UHSp0PEU3Jfw1asH05m2K4sw4BCNYg5GZb6
9XuvZOrjBinSvY7neJCawYdgQOEq2bDi+lYFUJjkd/ON/Cffc0T6L1UoZMUlXx40b5reIAUOeogL
iyEgTAW97vOKX5i/u7IZQcG7OdOIeN0DNJDctC3cZf/08K7+6yMJR3IrxawuzoFZOFwFBcXICol+
b6zFeyll9NnBgB++BEkIyrloTyS4FbyBPnl0WQ57HTo7qi2gT2rRM196U12i50Lkp+fTTFvWa4xT
PbpdGS0nQVjAZjLcZ+S/0JqMoea3q6oEVlDu3cQlFUgjsGoh6gL+iwJrUy0A97Aj4fFSZDKfyN/G
Gf5NK3oLZpBQ5PvqdOIGMHiPO7OZnc+P17z8zG315YY85N6/3c7WKNm+4+edoDuXQov4nXwhPphY
ZNHQhOt71E9xT+tmrqcEFq1Y4APgBinfBHdrPr+BfoiV8OW0Vph5InWx3wyTnRS9nI5xj/DNHE54
DtZvFWGULmTJ2wcxCjTISclvyqZ8Nz/cn3/+8Unpsn1Nr3OoQ1Ku49p4ZxiaE7lbyu89NtOleP01
4WgNmtYB/rUsy7RLRodOGoHQbATmZpBmE5KjMFQ3jCkqC6rlGshI0A12/6ukIcnM6qEJu6UC/unA
jZ4M63H/m/5fcJCecJGkaTFHZGtahOxoA5PN74oYu65ySETkXW1yHgmj0dRDQpcIIs6FILhFdnQX
8uD+ASjmux24oj+rnWbSMKnuHqfdnrxpLM8fZEK+0rwsDHcjOZ73NwJC1zvEaltEbEiiiEV4guvf
uT1EiuEghgWxQ/Xgw/JZ5Dp4d+a+bMOocpmqTHwsrh6bWzXGF8CostLd8/wgeq9eY6qvgtwgLI51
VqmipXEv9lcj1i9r7PBeBPu321vbm19Ys8tV0eKHHuybEsjs9uB9SapI8C2CbxyeBFWVkUisOFeP
HvKsDRQHKEiXHKblO+944JEcPFjixlhnW4nEHCrkOqhslM2YcQSUjMYs6dclxeLlfpIb20bMhUrX
ek6NhmnRIkBcIzUeefjVKKgZJLPj+FulG1+o/do9GDMyM/DwkwsUzIGDAmAU/ci0Ulby7hhY4yQs
1VyWtzOJfEQExOTfWg+kaC83L4OtnBeKic1JxhJJXi5wdmmKYymy0SQ2LbVaX7pXQ0O9GKfP/9VP
7PjhxFbr4BL8/v6Z/BHy/AdvzDerecpbKwnbTfBNHJ6piw474BtBGMNOlfD8fty+1EnZLl8hel6Z
S3j2fQG8wWvgpSk+f4NZIBd3tiVbr4NG7fhHm34i/rv0+i3KiTgYRLHkv2UBqJRHvKHKat40TAPi
zzBdbNXeaKvAnvWdVwO7S230BXqDVfkbMdJSwZw6HTjc/urBZXAJL3fin8YKikPec48lvpdoKJ6b
6/eVoTGF5crxgvjEaX/48l5RTzA3W4aSflJ9AYPb9sGvsE931vdltBq4FYxCPGvDXXLsPO5+vlEX
eAvpDLCuEmr+5zpzqscHF56SBRudLNIttsQJZGKzmsXHUlZ5hHg+N4iLDITF9/o0wis8r89FgnC0
j68rEpsmAlBkFEUTPp1WWykqKajit3/SCCYP4108cm5nqlpBmDWd2ojQYWI3VOqwxRzdzG/l1I0b
aih5/ouzTWwh6Z0pGROWzGfAvYh1WDzIqZO+EwhbBDtf8EVfKqXKJIRmnY2qD1qrj4TPYGzEf5Br
hse+RZbaJF3zU8fXJkQ1gABBAp5S05Rqq2YoNx7NiNin1D+/sOe8d8WzZAtJij2aNuUMeqtAFW69
OXEW4GvGFo8vikOWZq5xWUxDyDjKhi7zWwtGPAYiwREGtGFrieWRwsZbEId69u2+kKlJQA3jxwj5
e/LPxg6ESBiusAwVF00HIKwjuz/zsCnME3xSe51cQmELIs4hke8shZbdSNWhJB5Lje4k4UOcyCRo
NepFAArhDDPjk/SSfIyUqpNyOR4sturQ0jpOganViUUhWsOaYCPC9zpkRdjwMZbuNZXpQdqiFD8/
DWViPf+LHE2RhNk3epSpQmThXhXAfdOXH5n1ElVNqS52R0x8+Jlpv4IyxbL3Kp3gMKb7oH+T7uPh
ZEBxXZOjjs2Msh3nMsK1CxbJdimHAbwxyYHq0Q94+PkZng08Qo9MJOSXGlqfTumZYE1D/5bXYl+O
4vjfS4Q1z3vjqHFmbZwSJBzXIXINc7Fr9aCz/UooNLEfNNhg9Qi0LbEuGZ91TUajQMAbhh8tEVi4
ssUGad2LrxjxEqeoPRXb8PZPh9rKOkf4dAPMhk2h6kYwxhuWZskBbi+qQxw71Wzufmd/SNVTZ1G1
jx4ZwdN2l6lBAKKO+98zCkFU844MAf/PGD6CIGPEfCgABPYPheqYiAulPpI5EcDij58amHoFBzZ0
h2p4uUofNVbcfkB/Rwbk6gnMltiurIESdwiW1R7WwJGO9uin+rNMR3jZHn9/lUFDhp/s7/+0kILY
AlXfAos+lNuCe6SQbkCDrkPb6qGvMr3kRQldAmxQrnoQJhqvDlz80xm/ZFOIkyZYmMeTbj1/MTlo
dhbTfrryx4D70V7x3l1PtlvaxUDFF/rkdSd4Y1TCO79CyRHNPCry89+Tqxce3nlCAi3kWVNBErUl
c18EA3pumw6x213mldomRMmI0OQJ253IK/xUOEI3Yv2ShedLl1gr30PWhKlHPicYwpMmKdxth/Pb
uaPrqGvsuQwBsdpFoWox2bdpb0HK3zl+Mg3WDhURprOSK81qWUKhYHjF5mw4tindFMpmPh4G+4Xi
G96EFtuL8YiF+yj/d5wxQqVAjRN36C+xFkd9Bk2CvBrmBvLzxY6cR472tuoHcR2+9AdGJJoccUPh
S7isCizvkxa1fWZI/qFJAhoHTbaZ9aDbxRmj7yukKG23Cn9yMxSO5pLa0bU/MNKRHrvk9zpEwcyV
OKUzp1gtRI+JHqpsupGgZ9+YUEx5RX8Z2vHX0NZ0Abuu5ACwAdcIfxFfm6uqJj20/yq1ui9KeXOG
TrgkP3ubTsXRdTqKd6RykBK0AfHybDjg42Po4fS9gsx2p6sA40nroVxacCpiZMXefQzZjqqzpIdc
+FpyGuIHFqXjcUjqYhf2t9tsPfQyTEqen02Iyo9YFhucCpfeejU5IxpsEsbdoV4FQb64mLu5cXh3
8Ro3/9qlZYueBjN7wcI2kq6P/qSi/jftjeyOeFmO9NRR7JSYJE73PRs1C609snakTF3e5223fmyx
FLFMOfEHrls0Km1dZmZzKkJZGYw/DVG8PMO1CB+QMJQt6WArhhiN8muGwwBrnCiQrYGqf4oEBo1C
qwCSkO3gxb3IvaWCczFYw01DygXmWFXM6iYp6mONLUK6kjblLReM+0UMxjyBJOXsckWH8CkZ/BZ4
8pdaZ5l9Y0IIcMh/ncninDK9Pifai4t0cq8EHIyJeQ55K7eB+JxP2QJGCyHeIn6tYeAoeTkIpXPo
FCNoiLUOvtJsaagnEIo2X1/ZQ1dofjjvBOEJUQECKgVDMwl/r209pUfoamYJDqtesAXw2jfuTlv9
XA3bKfsg5jO/UUo6lEyyrEwlsFhvZyo2JKTt9synfxgyLP67/0ieaYggRvAKfrRNmPYPw4rUVD8W
YwG9kDc7c8OKKVHGgaHOp0y1hYcvBoeKI9cZ6+Or9KYEZZaRJCFtlqvgRHNJH/omNmM8FUCBSBbx
YY2rNCEvTNj/TK5uNBAU1Av/miaryn5qhiQNM6Jv7CRDx0SXzdYWqCtUz/Z6H5pok9jxPSZasc5S
QFrsvDIORsAW61nsdmqLVG8SKzOfEDb/jLMrpjaa1XqJBw2NsSf6TsjxLSVfuKOFpDxanbPSbS02
mRHiHt+8tAYb/cPNBs7aVUm1Re0Ac5eeoV5iClRJLW9nYZmzyygleZ59Qi1bQAeopvuQsw6L55/n
IjPPNVBqwNJbjEqWQGmjX7C+nUTHT7J3KTkOrAHLtwVaHLOuoffcl1MQzeTGYJD5CQZ6asZ3tYYZ
IXhRjxqjmp1HLppjEYf0/XVZuzQQtULKd2+6ScYM+aTRI081diqtSH9aUGpHh5jBveDiaCaWOnPj
sdkxwzl/laLM8+hrr5e6VuIhNyHNblqihvK4ycpDJD76uO8EXoBp6wwgvWwtwrxAmSi7KZc2K3bx
OnsQxeMLKZuE1R9Ta+bxRTWHs7XRpN+DD4DzM1DcVUSvfjQ42jZSrSizTMOSQmGJE2mDusgg38AG
ixSq8Q9caFhBbvxwskTjJ4RZAJ3vRcVPZoDTf+seJhkb5ChLXNVQAo4ZXaRRi1YofvyF+1h6lHPe
BZabZ2vk0D8JEJNB7fAPkk9YKSc11BDApPQLIFgv5mWmZXbQVd1tDRJPiM8X+ZlB7xDQ1h00or+r
b6PhtLEAzFNMFVR+mEgFgmK8u+j6JglsFuGPfsPgpBD1fDxiZfvJpjUFP4fG13dNguqkYu/fjXMN
7/VIdYSUiGVm8CT10Ph/QwaAXaf5yEdZ6yOkHDMJ0hIpQwQBxIz5jEHqMCUwkCPlSZhsAjDKiHgR
hxD4tnO9eJHN0jKnowrYzajDK0ElNEVCnFVGhzfwG1JokiZqD+wqUDpstRquHB8zMyPsOsfblcY9
Gj/VetQT2c20XM/DLpByI2UhymBQRgDTpca0hEtUaqK+a4wXVM5oG1h2nEln3yiEFiXCRYmtDExB
4+bcQNWpsQMsSYLBrGCLds/5t4tXOyuNIHXWEXBT2rBzTdUBIfMA3WYY7KE2QffoD0X9S6JeOf7u
BfFoZO2biGnpcutr2gnRWZwNawdaDB73vWcUhnQnmiDwcQn0lfoh238WQcfBpOVAc23Z4yOhe+fs
njc2GZhGdJeD2cDRl7k3EGJCfjbXta3T8HQIi12X0gvxis5k86TPwIYKKIAmeKJNIPxwDbsejwv8
qUfcQv8uxZ+woZX+zrG8qZr/PqmGZmPi69y5L3LovJx548Vl5n87B6Ts6k0+QSUUZqKsM3nD1zES
SCcUSyKQAQM9oJtCIN9TXhw0sVnKBnAloCxpPrOnQgYG/kLiUMRRmb3ubnKImGHtirtBXAeYyB1V
DmNBAoUYMiifJFX+F6qN/Tqd0l0XrkYHzickUNwYZanKRbroGSPXiqMYxiqxiS4eUCmiGgRY1koj
pVCLt63CEYXeXKkYyeapwni0YPHZJA12ie4B4P1L1L2S0DflZC5M61pHsfUumdzXYrhMymPDtw4Z
Sh0fTNy4hY7x+Ih4i8RzPaiVG/sAJuJkIkyxzCoZFC+Z0EvA2lofKM5a2uk97ModdfH5HH+EMTDc
waGbczZaeQNyMNUxDUIBBpOf/9XhoasOR3WqH0NLNjl7cz8ySrXyr3Em3qsXs/JXY6/C21F1qEkz
MUbBHnQv23x0DNon2NWrWiM+a3gvUf/+g9khWhFhX9Y0MFS0dl/oD1V+xCNlRTNPx2E5MGNSh8sp
cYPknMQNQ4w1NTC5bHlRoAljdhE45dbCW2C84uaaaV9583c6xfX2eFLWTkR9rK9TFORXolY+A/TV
4OZT7qKeFqFXDt9Fjq+mMnY8rKE5lY1CgUfkgPV2WnjsLd4sNBxr+Eg6fa/+PN7Jq5toykpiu0WD
9x8xM87WqBVlnvOWCaG866aetFbN9Dj/FvUAlgXU4dExsYbkAFlrcamMeOjRUQQbQDZhdRAS7DSr
ieP05NGP+v71iToqimRiGVI7IbIcwYN4ZfnTUrdcEFUGxyIdf/RW51j8/PJyK3fdHdIOC007Ruv5
TpygCXVx0TB+Gmxv2Yy+CGCoe1HsEyizREF+ub/CmDcJyLbfvJjkE/QZar1b1rfHvliyA0BxYQxK
tM9DHDjKIj6eO2NJXjd2R4xm93jYB+SNbQg/kJ9649b1ORWFrqPUKLQ/eqeQbFp9o1alR3B7Tjc2
WR4gs6Oe2pUT402MbfWY99Vq1/XA1IRIp6S8gi5TKE1zb0mNeLP+Kw0aQJflcxy9P6O5whpLpu7c
ZApP6lBZQa70IOTJtkUY67jrSAsHK1a2L8wtEoWE93s3iH8nZ/Dt6S0HyLKF86APTt1HhY3U5zJI
RzmSpiDz7MaHX7xSk5V0mtk8EPlfQm0adERVY7pU9kbMD9LA9f31zNOsxKEk4FcthACFQ/e5cxKy
fvtc9wpDDWRI+rSKBLGqaEQ4sl17bpSq9Z6kSptAn8GBUBFxaQk7DiykmkO5QWOy/h3wYKmJNJ9n
WD+IvyGQpuLMgv5j4nWPBwfSCaqPMubkJ4W3ans+exPjqaw6sm7mSCQAmz9OpsM6eiFXlj66IOX8
IVLWTDPoW//I/5sMyTrPXfqJh1Ax+82hl/1LASvgfHiUIOXvwxvISnMSQr3NpUFUYjv3JDVDu+At
BpZYK6W+xmx0AS1V/sXLC0LQbknihXnaVSUgJ9CLf6s6zC5MKQFh7/KZkgYZGM3q22IA8KZqOX9r
rCoYwqR9FKdPlcH0l+hRKaGkFlIY+stC6pz/WoHwnxkiHfM8ECYfC+N7s1MueSUDpCjqR6eYIGla
LqDaPbCf5IGUzLn2GVBuGBOdkWu5Hs62y4w5icCv8nEwxub5uUbGpYGjGgc66IhaGhS/t7Aqlj3/
E0/rQGBxKX2Hptw7RtOHh91p8V1DuAs+GbY/EBw4fVO5S76vPh6uD+Dfw2JkD0UlbdsUA7j8ImJM
c/gEHr3acLt8/4Q0Z1SXtQdjcvElkDxBxmeJd9GV5YkFluHweKz+HUgI/Oq8lmpxFVkov1suxAjr
iNARd0dfDIzGoR8etvtR3eUneffhVeNs1/3g+OPkJdJ2PbFeqD3ejMcGoNY5IhqsiCz1kTU+D9jE
8Z80eVgVBA0q37fLS7S6TlsYzC99QNzrc1p1uMmSBqZE8aZOTqwhAgBrvujrPwm4xc2cdHoEePNh
XpYn9c/w/AHxe/kXdXrK1Bjyy/V3n7Zr9M8oyy1ku2YMsDKp/6o8IgEo6LmWe+WXgTk+e3QI7lzs
t3Ogfx/9jqgQ2Q6JYhBWE2Ry1vlML+2nFbSB27Fj3eLWwiNms+lAiPvE2ukZHwoUKzt536OA5H57
+NJ6qB4lu9+RjW9bMdB1y6fFqmZfvWInzE08v7uqvr8sYlZe+Cby9ghRvNbw+bP4Cc4NXjb4zocs
Iza4jHsZmknuWRkVkKygJYK9SqsAcp+zvV+GCp2Lw5XSXc7AeSSDatrXtQy/qoZ6JOg/4ZA6q1U9
BmaAOzn9fzqzz679x95AxUzIRFfyKkT641v9+3pGIT0JRuHND9U3VnD/M1o2FvvSA1lUZXjewI9v
/SZ9NHXLq/WiBGjyFNxTb2Xme8rqLQ02uKx8mblD9NHDZEKZhUY4QB0E/SZVGx+PVIhmwdMkM6jc
20hAgVUa4ATADyb3gwpfotEW4AIllce14bS50pplJAC7C1SZdzrcqCkxpbsvnP0VlH5yVJ5YBDM6
PsKw+zcdQstO6HnSxym5HrbQ2xLSeEPezVyrWjh8WhsvfXqITF1Xbm9MQ9qg8RSRiCdaKY/j7NTN
CMqildnEHahjwcnpUSwZAxALnAhvj3P5953wcGmJ/OX4m0+UQNqWT042Q96IIf9QI3eO24YbWLnP
7eJ6P5KnGedRSvZwV1TFWRyljmSvKDJLFBoYEyWFFhex4zRIYrBU89/WK5dRW5YdV9AYWmplxtyp
Y1JxKVCJbqbFanuI4HtHFTNiOqbIWgVittjJRPyN8x0zeVfkiKcniMv6y/F81KEhUFQKqAuBy6SM
kCSTaO1xN20IBtnec31S+1avsW3TBHT+0qlYqFWs2Sc+BvOFJwY8dRqvGINUG/V7yiJ3Fncb5m+H
lmbsTizTN7VkwkSCpK5aA90fLaDlzsm2IOYcRLu6vblCfd05OtrnsBScMG5nVqBtCaHgDbLZDxZC
SKAUykj9GXTjZhvLgfvP8nv19hA3t0GUwmyGiv4CPcYekbELuYcadCXYEzlJ8x0uGkHtid7Nw+j4
jfDSMGwav/xapq9dxg2eVwnZv0GsQU5PgIdtu5Ehsx+p+Bk5HEW8qhVyjcZwYJIp0pmgqXRv+JLq
tl7ouHLfAz2CgAdJ8l6b/CsDxqEjZB18PAvyeWIGZoiEemBORWEB/gOOpv/wn0xlBdr7dUo7WfJC
xlWZVxFoOV95CVugP5HkwJVoB9HZaQcxhiB4eFtQ/ER1jCqVkJCj3quqFDFX9aCito7SRc6FW3zG
VNb3xD/wRW6TuUVMtNo926GVRED8V0brU5Ta8XbqYtwVCxDsuae8qcTZEtDm2l5x8KTJ4SsNUD0p
Wz71Lj1WJkIeJXXWN5rCXdnap5s1QG0xIGwXMjBK99KbqJ9boKXXl3WwSTFK0e9w/U3g0KmAQyPS
QYkMgr1cDrIFiYQ7F6l1fGqfzPDuv2DOKWeauJ8BXoRuKWGmxZnnyZx7edusBNe0xDaseYYeXEXw
hVsoWiHDH94laxDL9BeaNjaXkCZ3UmSKPPrmiIxOD2o1asSWIATcCuSBX7P4ej5EEaU3GLGs19h8
b2LHWNPfafhkWvsDWDGyp2Fp/U61fLzaNC5eIS6Jnb3sMDuOXgIA9Lxaxr2Z1oyItqQEYo34kUhI
g2pmQhFIPuoDdibL3kKsG/QprmEALApXM6FPKa4Q00SwEAoxvGsfV9TpFkDDVa6hYGicmF9Y5+HC
Zxwx06mxnKzgLkUanAD4c4PnF6wbA1bTDhW42hJFHWip9S1OmgyT7sxgiDXn102yzHyZ83HAwjeo
G9mce8qMw46p4pgdk775P/0xXG00St7I57Ewe3dHauddcubYTRGkeM7WHE5PYxqUBh3Jp4/ryQ6/
KE0y+LQOgzbQg2qAOapTyJ2zVhuaux2UXxwkywrptF6zj2c/KoFNuZx9EE1kolKKA+2R0x1Ir1NG
lQ/egaCILRKPjGa5S9EXv7XY7w85kdvHHNeAW6wMd/pLXOXOXvGuqvRgLA7OtgWyt96xqPwNBcj0
fz2SViNU1nU0hW+/G0yudI1wwIaDrkNAc/A6LjxIYdOxWgwAhjaLDK49i4xsIVVSAHjAPGOVdA56
5kCkAg22BYwJF9hi0PdJMEpInI7hUoPQkS4qN8xsgA6EzFyayQeQ9oSgKeQCWbyW0+48S1Q4yyzA
VSsR9HhmpPTU0V96UxliRzbTrRt5mlTIMqDPutmGXCM59fBVVCxUgFJWRCJRst3AVLuxLWe6kG7q
No897NWJlh61lDqLDYwIXlzG1LPS6320+S3okSjh5klD7ic8WQ5Sr03pxmG7O6kFM7uG8ZvBF+Wn
OZJIG5ymTPHCRa9vi5dwB9xxtQyPasD0YM8ZZaGBtsmna8NeY9xxgVEOJuaXL4T0sxcveLalJpBP
DKeD9Z2Rc8LkkMJi0U+6Phinq50L4AIYFre7UImsRNFxhNA/rGPV/3lk75uYfG9qwKJuEzZiIgpN
RoZ2BJDwlWWtddZ0WfsGiVwRr1zHXk5PWPfF8YYUFgFJrtiYTK7rUpwj49E4poqdUmLiRY3oqXJz
r6cHtEjJUX8lpVaX98Tgebgb63P1CXyC2gLhPzXINMz/f1C3uRviqdi4UHDeJY62MBZq2FZrgLDR
T9+Daqq1Yu6EE16Uh8Ql6aySnxoFqEGb0yiVZ09qWLEUOYGTAjXV4OOPWxkcqSu20vXxLDJ8egnq
R2JRmCCLXr8vnU9MmfuSz9JLYpKiIVM9oGYchRQgj0S2jXGnnCI98a1IETVmRBwVds4g4Pv0msFX
x+LHCGf07kk4xNFWydv84iLoEbPd7DoFrIc1C2GltgmtldlRb/30zvHR6n/xhVO1bVfaUsHnQ++4
8lR+k7ZnYSTRSeyVX/CvqHyQgl+IKtn5NJQSfWv3axJABNR4qT8de2tChAza67w+9kdUXHaRONSy
grOKXZ2BLGGyqVK5ZupjWp5Zbh/HegfYahW9C99O8VHJCKn9orkF2okiaA7Wk7mTVJemdJXK16jg
m1kMqcZejRJ1kIJuT3tYMPpXv1d15OnltO38n+WO8Z+GKtClrO/sb3ITHdCMRnESEQm1mO4tUQkD
I4qp5UTQdTZCr+PhCfYhI6xg8QAlq20RkclPiqIFegjhaIEJIajJpFOl6vaXaQlk300pJ2WdUOAh
/JAE4Ejf1589AUh9+7jCYtP7KxXgOhiBHJD0P4r8fOflGac95wF9AFTasdGh2S1lQZZIAsDlpEfb
0+Fw8RmYpUcdrzalI+l/6lkvcYZ9Jc0HC+hJd9PqaZiSZVADihrTCH4kr7jvwPgp/yBwbhgnM9rI
UvNdmsNR0trVaZSC63N2I6ICOA036aD6+kQui26aw5XLmdICRG1sh26OTmzARHPJXlSo3MwOsPr3
DCfMZ+PKPCFN7LKtegAZpX3qoNjMWsxfcGWM3hrlPYY38mn74IVnQ5MGKc5VWuO0CkDKQG6Oe/nt
AWgZ8pIa/K82UN+CUEIgAUbNJC5hYet86yd2Qlq6AQVxgvf7VW0KquYnTD28WNvEiwvgLLfIMfnU
llHZye0cyWnR/hMb9f4F4f/UdqObBCVVo8ytmalffet53u5jh5NygUpeEqu04hPRLDjLEcrveyzU
PGz4qH31NJYnI+8iXyk9XZnN9dIyYy2X6e3ACyHZ34WsN3WHNwIHNUcfPO3RAGkXmJMQg8094QKV
SM2SE26mX+2g31Rbph/e68xvnI+9V+Jtjm53+ZVaH+Y+Wsf7C+DQYZnzwCcSF9yEySZpv4i2JKsE
sST0TjP1/KpbARhKfbU1T/oerWmyDy7w/eo056ftJLN1Ai+3nRYKp0QOImj5XWTYUXxqGuFL0jSi
dDGFqieoUV3sN+TGGEbXKYSjjXlUHMvurj4F1ItSzFQlpaqQ1XNsbq6tihdtqdQr3gfqv889k2Kp
f1iMb/4s8mLdWUHvaYNjjQIxQgpKBKMJhRt3wHZXb6C53RmkrZ1fIChi5YSuMDWYA/lnHIvsediy
SUJnPtCbENKLVHzugyH3UIru+qdMHgESwspm/PcviZ8nKHE/FP4PzYLmCykw2OPQJg/2JmYLESyr
TmbvO+mbtr7ugvXu1t1jqj2jNwp2GZau3wVJyn+EpGLHfOWPuy6oe7Fy7zHxyI7hizYc9OHkKYH1
oLXw08U/RqXCYtz535LJPfFyPMpgc16ZbORsOTC3PbNkihgzKQfeCeWFEThveurLaadqK9Ijfnxv
ToAp6ZRlAcWCPHyvQeSKWFa9T/9yAoKLSaGytQUmgrZ28sY+OdUyo+EPp5zp7NcWrrKgiglWkQuy
m4ZjA81w9P1fTTYeZZOYo3gO6L/bwTQp0l/o5bXHdLBwFdA8Ew58FwY8g8mb6QA1TfqKZA4VAZLo
hMRP6GHtSNPpOEnDlSbmOFFiAzK8q5nIPIjGBg+Pl/o5RQHfinWbymgDhX8bOiHasJ5kAx9K6vyi
97LPofI82VPcMXPyJBRqUuFzY+As3Ck/wuMKmDXtElaGylworpjoerQuL4YapnjJjMFyvRyg0XAc
sT0XfQGktA5iX+ZHKF4AilFdAP6yn1/ogFbhkWU8d+R1r8613c8qlu7r3Jgn37mX9XXCURfraZkY
PJcRfva0dh1ikudUkH6hS6aibJfNhryh2qREXFJLA4QPpzmZcazrS1NKpjY/Jib6dT73ZYwDMoi9
dqgv8gLhgGZx6l2iz7hyuGlScRqovle5zTl+xjoJtl5Q7ApmHFH+Ng5vHFzvRZerrara7Z4/q/Q9
MJiqkbJ+e73MNnHZi5S8I7Y/BWoNkfV90kq4q7FfWdOQbgHX6Mr4roswyNfWYk0zojglg6AOep3T
0u2GMRC9py0kSI+tlu7G7vz3G5DucutapjhNAraFb8tGXD54vE6V1Rdn5V2X+PZi824SJ93L9Iux
j3TmAlbOvuADBz+FiHH+q+mfZZzlztoEUh8txPmYpm5C9XWKyHZHQvVrFPT7iOUcYwWVKfk0PjAB
4YL6Dhz7X4MayXNsMqZWpesYVi5QW+ddpkL5fx/4JhBEtLGKwnfJhcjLdFuU0twC1OJPC92wD9GT
aUEe2iNd/n0WBquHSqHGzsFyxIeNtrJMkntnbfwT3fyKKQrQnfuBIeqWvR1hmwYDsS66BMdeHIxl
w/no7yrcUGVzZoDv4aRUJvxPkpm/G3rgT3ue8LRV2ElgAU2wAU/OfZ2v4pGpuTc/kTvoe24bip3h
T0aBNYM6IiebdQrCncD1RuWHoxjAfghUGqpOrnAr3NTFntV+xV5XdjgV9cSjLDZ4+OKCD8mKb/u+
9PlyZ7l+XDA+l9un8Buno3rzecROEZhhz8BxAQSNmUTFoklYQEQvg1tcGFWlhM0R4ZjdTdIcXEqM
BqTa5LZGigmgIcbJ/WvhwOcFkEDtbPTQj5FbMxRUWikatytZHWumaeh6BOIgU1cpDPZ5i3W3BRIE
j44Ds70H2T2E99T8vuN4eEWZDMclblNf77OOB1JzKTKKFvnD7eROqN3VeR3PeiVeUlAEb72u+qHd
+y5ern6skVIF1RdDaj2cdNnpAPret9rnVVo8flKkjU4z4m1YR2KPjVPwjKg+XnlFq55/y0gHGyF3
b5CtF05SAwY8tXxVB3yH5tw9vNqNde3T+zEgNcxXqy4DO5/RUQaPKL4jdlD2BI/82KD+4coknvN7
VcAjYxgrHy5gio5b2GZU8nLeO8JZr7nQyNn454T+V+YAaohlwYAUsMh6KKcxKZAKqDTRahHCB4Ct
+ipr+EBXr7l3X6cyDzeNALz0qqkk/ewKcuPBNvWL4Wc9ImrdLJRNuwjzROJ+79g8GvfiZIuqc+w+
qj/qP/1Ehs45sGWUp1563F4/LW3oIwkepoRMtHB7urTsHD8NbCpA4H/9qp+w0DJvO+SiTxH1HCfG
d7tJX4nCRynoBRNKlQv6tPKJGLJoq5IVTh2vCkNlPIN5PpIrjaMOYbeLWE8CMVxU1htmefiF0lJH
mcSOt3hl5py+QPrCy/6IU/TauVIX/+d+KhAxKyri8tUpMuM8uOMFAde6Y3PShpnfCNTMT+KgP6Ks
lRKab9wPP6LCcAHddOSWKSQtJ7J2xWs7a2M+Rys/ovuBC9qsg4eAl5l5+nVoH4wXON97QZ4RenCE
KYvVpPiMER1sjv0jTOBig1SDrA0EGDHJYGowBd9TMCVhdbED7YLvdCgUbE/mPkD/4Zw6MEsqE6+b
jqdPiD1GislLz+M2T96a/lY0GtCLOwpxliGttMCaHhGqcggIm6x8GqZnGgTTjoo5ItKSjPVMPZlO
B8+nN4Nf4pPkfs4OqAs877k/ywF7LYwF+TrY/8v3wniUwM4cU13ViPt+9IPivSsN5W6RYy+Ef5Of
Vsgv92yd2eLkX3sTv/a2XkRv2ww78Fh4O7rWC/Pn3QVoXP65vrhaWZCQG3TRHEltLhd+dPuQhK2b
L8Iwb/pzU7hGNjA53X1N/7R4KLR9woibEfo/5+V7qshvcAcZT0Ftn909v3+Zmlh60/PDe9Dt08yu
Djqdgq1WVBCW6BtyWaJYGUfT9kdvMIfjaEQR8deXI7pezts3rsEP/fQbyYwC2fpf1FNMnM90xp6R
mvTTxZv8FlSgMStHQpv7GzFA5uxLXtHw8aPcLA2b0Q4K40FQmlm9KicJxzEpFCdtzTf66IwVtVb3
8raDwgM6mS/oNe2ktf/+7KRIOt1wBYerhnhUJkIjUBjDWnG6krxLL8UgqFRsl9QsOmURb1mqvTqp
bomK1k0il5jjHXDK0Xsa+lnEaaNQocgoq3ozo9ESvF0CaNUd+L+yFZa+8FOMLoEpAwIBXnUg99GW
38AlKxYG5uOZFkQtIWbN1We722RH2fez7qNdTL1TUqSBq+g6ZIF/MgWRNaqOkDfGV2CdZ/cLdeVd
eXG+EH9ar8G3khiyHeFnvxn5xeMG4iAWUX3LuPl9lqxsaKHyVEcu7O0/7bH6ZNbyPPc4M4qAqUoP
wm9D9PXgjqIfDazyfTFvL9Djn0Um9tsPh2N+0vdjc4oYWx+wczrMFtExIJPhqOZavqAziJ4fuLxg
76LUDsspjYPLpcmJGUa5lbIw47auNPgQ+XPyZhbs7DxcfweYP+g6r49z5ogPSzXop8ohYBc1isvx
93YyuAa4JPEBC84ynSAqdGoTvCHGVvruTo9hdmHEC+HODhv6Ma8Nn7Gk4buOwdYCj+gwtc/u/Fi3
99nsXm85ym3s0hO2wge+aIXZbcduhbyOZ4OXtXvqC11olShJlFfqD7P49bVSWB5TunRtMQhbk19u
FLC/hEpUsJsaOLLTRTeEivO/Q4yzh73Jnl5FmwwlmhrSN2HP85YjYrdXecFCqsgPFO6rtUZ+tsrz
3gl8NclNpXAAyscTYVvbLmzRgrvkA9/3I88Wrlc5sayg9fVwOiJ5NdTauZaCC7SVIxujmED1k9qo
n7S0P82Ssuch21V9uyjzCVxvhaA5LhXIqQJrYK0BE60IJeWDtmGfczFx6f/9N+3cppsm6p9hu9Xj
grNXqGCQcOeAlHf7MvjPTzHGysdU9iOxdGoQ/fphFgVGLSoXKY0o+oEWelgEw7mZyjGq6rlHISjW
IwgIEiF77f80LG9BrMYYdVdcDDrG/RxCQ1m/4i+9wb30h6QEDPY9Y1yaOsmzIFV3TDoBEPaP+pm/
Mwm24Y+jjYOiSHp0BrpDJaVj1Zo7kfetu8Gp/G66zff5W6CvUfoB/b+MB0NRT9xwYF3kyqb7Mmdg
7PtOE0fHjnboCX348MeDLQflFmpsuyTKIFdSz3xBNHKUiN77x6G782066u+J07GV1J2iCHv+o9HB
ZoC+Cr9pkubtasUb9cAecxMjAp+IIx/Fl6iQm053uDeLFea/TAtKDVsyxp3LrRBSZo0JHw6upKYC
OBnCKBjJ/S2xTqGqAoRgKzfglt+SKpBYMLnvWq3Cnwi9xDSEYyIrbkwZv3lmyYYxVw/SqxKYYr+/
WywmKnnkTUqeo/tjPwaeSX3EoGmNnOOHO/5fT17ylU1YqKtCHpWw6dfBHzmGKqSHbUuhjXdF92Q2
9M2frhdz+S49fBcXMIAYX9erpLmOSO6y+5zOGh51l5iqFEtUlrB/YczVIVoVK6CJ3VSTUBWb+SoB
bjhJ5rA99tIdGZSc7AZeCcHRPEhhO1K+fLAiRRMVkpuywyPl92TRYz+kQUg343rGX9tXkbf7L+wj
zbVV0SUueQ32DhWDGVcfX6/Mkh0JTopDN33rtcnUX+p7XoV7/tE3tfzcK1Tkyu3EOLB8NzIQls8M
knZV4x9OfAy9bmUzBYoj7NZUte1DicEQjAQO46kIwTtwKcEdo9R1qiQV63Widf/pMfe6KfCbdaw7
LhjG3w8jTEw8EnIX5AwDSukXHnQ+QtT6NR/bsAKggxpXBaLDvFFB3W0cYnSycuuiY8YJDLcuumgG
gyMIXM5ZNWg6b+vT3yhU5Slhb1WatPFel+iJ5E8myNZ5MgRIVoYrKAtD2qiUMZAzJLXUN1ukCp/r
U6XF5wM091c02dj8AHMAMv8Ko5Wz9Q5jbUuMDgTOHyBaRcqnRiSR5Hj7t4S4++lLbOW7dCymqMAn
q/n4ycaAEpsWBDsxirRlSPjkh5kNUMd9fgt5u84QzGd3sWCEDdRa4CCtjRiy4eNwu/9MXhJYtJGa
twCW7iko5kAuty0j0TpB5Jbt0Uch67RTw1Hd5t/WZrT/XOwHv6jnKkZ2nhyrRhQe897wEc6yshUs
CaZC1U+JMBHtyibZasUjNrRQLDlIAmYh2AeVvZOMPeR567kqs5qAOnT8kLqK1lZRkbFZjMCTpOmK
fZEJV0nO1OWcMGv4PwcDWPKWO1dhy4csxkRUQlZYBTslRWCtVJGfoRLa+CrGTlp16eqDg60ShPmV
WzRZF8S0nHHYAT2vqx2DAy6JHYVuPX8bbqARK3H21TQCcl992zDkh35HkgHIEFB9rELy6kASk1pO
6tuW5FMI0PZ0XBIJoLLIbETBBZQ+Nc9BtuWyo8j4/IWiB7N5BLLfZfkAofenkcELgdZEb1m3qwnP
giRuVJod2znpJ4WZbfTtVWzGjhOPUWq95mCXZXc74/33Ir+nu7wEDAutoMBqWvp9zIPcpokMgacJ
30F8HZ5QVNAX6ny1PliWqiimUNtiLtBW5Nf6ToImPExH6yp0kwXpEPhhnBysd9o2E1Qw9EWMlVmc
J+gaFFPoSmVjo20rdsoAYfa6bYctmF2l+BCbLK//pYLKhFJLgVTR9tX3Ag/P9mD5tIbl3DX5+Fdn
/2nRKJWcNIe3QfZ++zvmLUnUnrMU9TIFODGVhb6+U8KLyjqW2Ap/uUUoOX1jWaB4mdfBqhFc5pMJ
WD+8onsI8PAFI7bmiVlctIdcybKawRFI60gHuY8k0UanM2lfwwzzsst/svWQePC9UeQWESlO33xs
Y9v55/UMuFJ4CXhXR8nnAvZOxwtMyNligUK2Y5lDN3Yr3IhGXCvl27xyNuNuASuo3hVU3vu4SCfR
NYi0jFq00Cy2YuBQQg+CCODfdlsihczmcFSPjGephO00FEhF25AwxPegJM6XdpWa5SPExqFH6LLC
ugx/HetsM9oko4Y2NUDRfSDinhDHKJoEl7uNp5RGWpMt+EkjOniB/PV6oQgDAKzeNgZS5+NJIiap
ZlQcb4sao2Ro/ZnnqPAb2QCMNYW27FZZ9/jcOsruaazZBCVMSPmZv6peiqNBKZOJ6hDIv0oO7gcv
MjTqBOJmUsxyz3XyJgFwbpoSPaJamNhg28oMJ8ZPqrPNEM4ZBuQdw49HA+TXump/GfoAxJEaFNRD
6MsEAR9LQ2tYj4F/rQUytN2AdQVYGK0bTTtoU9h3pFXsTmygZWrytOYrwQ2k5d6ePjguXj48Zs4Q
3ViGmt5Yw5USalOUI/9xMBhZQiaB+O9I6MqadsSO7Wli3sX0lrgaRzX72GDnVhMI0DiZNK2NhsBh
Z49ib418vYgTOmG35KmQBvlJQ60zb6wmDMm7eVDS7cUwTUBhLqICv/rO2Rygy9Cl/HpX7v6VjcQ0
CuEO1xbgl00Qzd5NeXLNWZFqKF9mIHbBMjUiTbADh4uw6w/l2QtgdtzoqTHT5LICTboPLwq9/mmQ
VJH381MbFo2si/WWUnNwrAmeXxdat6eR+VNQKB0NE8eZYICpvuY4cr7LKEi786jy5GCaikxEhoFA
ZNkQvLmGuYk97cGKuII7vSxMYPbB7pcagTcpIybjP/qKzcqB+xVwjqQlgDp1udWMRKPYLox8WDSd
xEtrU8bwnRzyZE1QGaR3EvLzvOaDooZCAX86hmNDzy+yBx38ABGIh39ua8Bu2yP1Xmji8DqWuWlO
SIwOfPQ5Unuw0gzo43cZ/WbyHBjmjmmPFmAhV12KwIXoN/0ThYu3Bkw3piXVSlhjoKi8CW0yBJx2
IsaXNZ6L84sALdjp3Lupf92sbi0y1BHMLRTgnBz5N41ODkbtYK2XqXvtT4of0oDInkLqGuoQsqvl
PCBxZDcgR+ne/VIYNglUzwZguQhhL4EU0OoIBY1zC7MCOENP+19EjYRPxSu1BsGqkTx81gOQGpkg
bGWIxy/5YOQdEA5KZ+tsWjKVqKNikmPeU5/tjooUZQjujpnKItsBGEwL8+voKehYykTzGb/xNoly
jahl1UqCUQZzUI/zfh7I0gs7Wnv+k/sd0kSoVL3z8Kc1F7ABy1jQjcvXcciU68A81NfN4CeibOmK
qEyaxWUDe9PpBjvvUMR1MO0jLz2s5OAA4yRzZ4HgNBsDRA2xuCNFp67YF8NwHl28IEhIfPh0MWyz
3YqRYt+XqBAW03qnGWVGvnqz1qbvNsi41+x31CmFd2deYhWcqBk35Z42AL5gee3XrgsrK+kE+ASh
B5v3Z3V229X6oi4jIEg6mMl/654OaWvzyfhpRxZs6AfPhyGBYSk2XI+f7q5bSb4/kPHqqsjqPMPM
Z4fGS7E+GMdIKlnSJCFwdyJZqI6eLskqlPT1kKODDlCOoeJbR6FOhfQs2Gk/hLpUDoVERZiW/RUe
XFmMxd0znEMNpAoDgh7cZ7cYU/gC2TvFstVPvIWg0fo4YFExvts+8ftvZSq3yxs80X8el1+9o/y3
QhmPzyq2BjJhs2jGdAAjJE9Ys8y7bKQ20B5McFG/8gPWhHFC72+YsJdS6A9FTMoNLa1pwP0jm5ig
lUDhOBOyTuG0FfFhUqO4TSC3gJYzJG/DBKSzRrbHAiZzVSlNVE9xoQs2YrMoDdb2DVCi7SrdnzQW
9bmnSQkvGkxovIrJ34tlq8y9eL7wdWySQAxMoXyTGRZi58JYi5nbiHhnDKwQ4bYTbKZ469RWXXlb
9ZBA4wL91C7gxypDbA6ZpJKL9NiK5mhnJ86QmLCQbc/AtrEWz0SIhYYsrVbF8isvXciniKLL8l41
2fjNcuj3tpVFqoGvsOMe/CAIX3IDz0eFAO4MxGZu//v6U84Pf9uodFbzKH7HqEgvYFPcPCVe307E
jW4J+p+WGEKMcVm1gJgSUhSURVeM4TCbLUbGW1tKWVBzi6ojVR8GlijjEM1W17poZkeATvqRWKGr
BH80B+3dB/q5Ddb0Tu81aO2A6Cx72dTm1EluDtzFRcIWDiMTMihz6sUDJWy+Ca0FGDn67NhEpqPS
mQHKVrA1Q1piU4GRSJ9EYWX58uJM8kCsKYqncpmrTArXy0Ge5TjyFzBY+6sHfxOarecMz25BJgqm
M5YxH6az2uWqYmZmvDh6iqO+XwmxQvVH1qZHH93lOytdVPvUuxqtcdtnKUQl9Lsy8hmq45RpxY/O
Kv2cxWV8xRaH25O0gpDAorM/VGfbXN08gaIDEQl/P4k6SgehHWFRRaWT5kBbdm+kdPbtTLTiZFcx
aIL+uOUftIv0QW7bRDy5iFKxInrFANZFlWw+3YR0hIuawM00UKIiTUegBuDl+Pu40JSxHVgol7/F
iBvLJpTnOuo9kfOM87U6gLQQMPC5uQ3pXh5Am5Ooj4PkxCcsyAVIofGb+5kFKyEkb4cNPM3I87gu
Ldrj/5LPWyUutnmJ8VdjTUO/i9vO5DZVOcCcgd9r134U1FA8W6Vf9/1+JPgV21DnBZCEex/kNfit
1gIUvK8wtgqUAKTo1sUgVYbtEavNY0TyivfVCNKq9k1EuZ5W6jlvcygtKIUByVhaip4KIg0X50JK
3BcISOTo96vDoLJmzzG1Fc7JgqURRNF6XDALbCV0rXIYa8OCwnLgQ6DY76XLc9sUNZ82Qumj2pns
1rAD/MWuooqeI71/UYSj47cqdG6Ho++/3m0sOKtEcmr/IrVUlYhWUWIFZ7GrBcw6axQ650/MLT+N
z9GrhleYukF1pTJxj5HkdBtgoOldsgMLqFWz8Yg1DOujaQT+hy7iWw6OSqIStf/We91FGZkAE9us
lcHddafUnPCEHO0A0t74hfqwy8lXcsPoCAGzxDBz/XEGQha0dI08NbMrAzELp0uP0f4ZrQ/DTYGW
Euzh5Ywlm0i2cPL+jd4nmeKtyKpY4nQdbjEFL86tDet6SVYZz7JnjQQ+I7QZGg3YaFSbS6YlwlZU
0iKEIjhIHsKyiNbYxruwalWdqYa11KlxYyvQ4yXJyrJmwKC05t+8xmxoyDJ2+l3THlvogzAURzje
oEJSGaFYzRzQ3Tu1EGzQaTlbZuOAHZu5nkYpeQLn3kXxcx6Q+It7uDBKnFEOrvOGa+UOVe9H1cCU
a760HJTHnRRYkf9zgBD6+IGK1d90cmCHnTZb4hcPOGNkgklJ1ggXjPDijMIsUz0CMw2KkJnL3G3q
oiesy9uyJ9YwMNb8Nf/pnWWCbshEdGl/SloQdt+12OxDDzdaPaKFwUmFqoRGSe075V4fwXABSrNc
h2mC62k3cFAfUdHh60cvFJRBIGqOuHqQvpybViO3bnt16NSqqHloAhL9AT9sbJqdSRILnkRA/N9+
EM7qXUn3f07YQLoJLqdYgX5DONhHmbE1SnanmmhO0j4Q2ArBJyHzN4tgjs8jn/Ri8Y4mwvYUZ8Wi
hqB2f1mhaZWdy90rj13ToGUd7JDVNDgWJT5wOVyNknF688zUBps2mg9+ZY45jrpOFMV2CFmx27AL
CFoUaoYDxas/cgpA5BZ2Ceo9jPFJ1F0uluS+0U+NTbOCaaXEv6aDQhoXBhFyOANzHvOkdrr9CTKy
u4DpI0ydsyge0Fvld/dhlJeBcEcbP+IYpvbl32vRsthT6JQrw50z5rthzGzl73aLESXLKIdXu7YE
CglsWei+czIthpR9Hp/yDyp56BLBwHAcKg7N0dFvVq3LG0afXNOQJMhxv7wHsWG88eFsnJ2CtT1k
+I5cJVyOyipUSgEZsRAxSoTuEERM7g15gwSZJ7mJ851ei2Q2p1TbS3ZpPl85zvJKO2tApn+wv9VO
tBLnrltHrahmIkHyDWrdvKdj351ZkeTZpgpdXm9fRUTA+cjKQAKjLHKQ+269T8aYNcyM5dwdFuxc
OzkkCwX3e7La5/7WvUZDi1iVwB+wFGdQboOIfAbOhvkj4ugdM3d2ybuRsLuYwzlJSB9elLHZUSge
G8OL3/ZvBzKkYF/E1LfrzOaKuw5tONFX+f0szJoU2J3TuEpYowz8X0HSkIFR4VfJvLdj8NdxiUKV
Zp5Qy3EEWI+SXO6S0p5vtEhxhVXLgdx1JKfw475kLprlASm+q+B2Vf7Sc1BKTZAmTokvAxyposZX
Rlyf2Qv6DZ7skWixTr1dsH5oSoOv5+Ej4knfj8t88g85K4OIkB2DuYiJ3B1f6LjHgoidVOIl2K8M
kVMLg8yUdKfyK705y6AVni6AoO7b0f+C0ItoJmXsVOG9lckhYxs3/PEPEem9BUVWQK6Qvjnws7ul
cWd48uGbJujjrPDcmYxVRFdnZd2F6M9Kv1ZRNwm8XJo8P/foBibjFSOiqq+8Tf7oTuXr9p9xhy+w
tRP7QAIqC2ybeEB0ReKyPdvlY841AhijK/yRw6Etv52Kk9zEkVocjCGI3XCmGrSOgr8bxhOuXqqr
i8v7786aZwVgGnyRhLyDQTQNEvFP4AwM90hjh3ixFskGAy3YAGQkYrLV3eoOLlIC/+meVAFpYO5Q
kTFbx41VhHO4ddEpO8h332XxdHdwUvpZpJe3OD0GvADEa1b5BLPFltpRy/DzV3fdt7drLWSPwJiO
KuNyTIW2oh1hdvsQ0bgLywqbdzleRILh/BpnpMfcebcO3EitzIP9Kxm5uxVdeBGSyUdIuKU8+30E
tcL5Dl41ls9XUWBdaP2SvGSF0KRxEHEBZVM/XimSlVWOcUdDXBWb3bz/GbQGkIGK8F/2rmrE1gto
LFStkv8ch8pzE0lRJbukj1ER9LqFEGLNpmVZjehoON6cUnpjXOAZ4Q+VcZslFdA9yQFYELT2tb7H
L1xu29h0blPjUyg5Q176eiBFnWDRx2h0FEsJZ8DcXUs4GilqNYdjrMIf1iUi/NjO6YO3GPVvzhac
IMkG0UYHall8ErtCUZWGrn2xNn9EZr6/WY9SsUbG/bqlDo2C55B1nLtOqQhQ3wn9LjhDiXwQBWxZ
KmTjV3iw1LEQIxpsbk/7gZIJRA7WIJeF9kmzpvFJNbWnPNwH2JnJMszEHJYCSM21K7IdxQoSEskx
UfreRejdvxrllwucHLsy77hPjyEUASmyXLj7QKVh0cWHggDoJ026io4Lf0ug+5VYCf+1SwzYGvuq
fYayxA3VcJ5ub3b6bEUhbUpPCi86aE19Tcg+2Z7iWsAPZGfUg4ue1nRwkCuTKu5AC2x4YKymWri8
cSx9qZT5urFfmZqyFCmyxYZkk7gfGdCZq692o0aXKrELJ5CEpv4du9POjFbDER//ypmI6h+ibARe
07Fc1e4ml//3Mvg9VBkfw93VskyeVuVCtNnD/GhBCzvPWxCDZlIzmem5YniFn3p3h7fNGb+WGMLq
6iqszc6IEMGV4MZEsxd9lMc9FRyQy5hANgo7Kj1wpQGGEpQKxcEAJWqYBwH9eRXMlA0DXMu/dW3f
pT6kxppeAVDzEd0hAHj8M+fsmFgQWmV8lh5O43Rl27goBmaOV6luI9w0kOOCW9r7j4xN9PF6i8JA
4zOihNuVrXjfg3n04u9d5QpAIQAy11WKh5eu3dG4uIB2T8n6zD6q4XN9vRzSg+PdqH3F/WKhZ2/2
M1ZdKzioYTHj2ZSevikFdL8xz0EUHVQGZpdANG0tcpw7F34D3KenzgvQcRfMdGKqNRfchQwbBKYv
LOhk6Ek0qDEjeqmezgZ6Y7dNqcYn/LQcUZrbR2/aQ2lRAw6kmVKJfi4kESTF/JqTrFr+KEbeBy9R
mDlOIajMB5+5mc0RFxrN6pMC3FIO0dWoG/K8reVd0t/6L4PU5rjioJO0/8ekpAq+4x0CIt0Hcw5B
eQ247oWDs/HLuHlmmtgVTefZnBpZR5FshC6BVUkAGrdstBadrb9FDYNNUwcGcvqRy0Wk2cPrG10n
sORQCn5lh0R7mvTj3ej1n4hod3R6mFa0T451LkIP9z9FpQ2sK5Jwt7SxTIlQD6ZGA4Y12AhexUX/
hJNooJYRJOxx2NYpaduiKev3xx+HEvWExpEFYxkUw6jCE7klBlTz7IA1nnswBMdt7cyj4riFrnOU
KpjrVQ1HxtJYbLxvWlkhfmFVJZSEV80f6qImQa0Ls4cZdK+hwxAs80r7PUm4q25kKERnGpFNNeXZ
0HbO3y/9oe1KdHWU4GNf9Hm3rqGkkHfPoeNcfGHGcEK14HPrRQbwka+T1tWwtYwcvGrDDiascMqm
4gJVMoy4extJWZ6axR5He6rxkL3Ic5O+zJcUf3ovR4f8kE7GkOM5a86cFI5pJJPjyV+aEL+ofrZG
eEH3voHRUmUBEljjwtaQT8bUoWKBSVT1tYCvxEWS/EUX9oUuoAs7p0M8ilRDMXH/z3PNEKit/yLj
/J82qrERfX4kOSmG/163PFPneB+SMVearXpY6XcnDm1WQMZY/rQIDseMLZy++59agljw1Cw62rX9
nq7BGoYqGmoD6GTuXljNMlQpdohRT/3PVgsNdMlmrWjdpgug8lLEgn2YdYThdcyz9WYMKILO6DuG
PBM8xsSBooRYtZG42i8Wy7312IpAoaCQ0kY+xxphCw+ukQLeG8kqxLx2gfqcjECWWujTRg9gok82
iA9TWze1FdvXhYgwbu5KkbaVcxxvq1IMxVJfcpG4YRXeQRnoLAnkkB7S5BSdZxhrtRLNpZahb4wp
PgcxB4tMKcIlH2rrOcZGIjZp3TYoNCPUMKmUZzqscBk0rbNlho+AeGibSaut7EwuggsDJE7Pf097
bISY3H1m0zOgHqTmdPE9rzc+UVsF941JZ9+RiUMxRvv0n1NCmZ1rz1dMxqVBQs7IKgoGjk3AjFVw
R25h5cp6ip711Zkknd0yOSpWbMvN6ttD+O+iuPqV2tPH26nHdP+FnghQZB+D8GkzPbOHXfNCDC+e
Mg0ZU2xGm8JagdNep6Msnc9SyLuL1Gx8UKbOg/unvGD+v6R6dxQtZFM8NKirEdlejAKgfDcJev42
1i4RPkK9v2+fQJeMpza+x7ToBz2oSiQg45qjGMogxQq1vd1O0zQuy/WW8cWFxwbZId2VmqZBvwLw
WYxNAQk5yMQeeO2MhzHCaHl2Imkp2qfHXShRs32ALeXNINmwsrTz81nzl1W7oQDqwTSXfdHLk5pU
v2LGENR92FGVgoEkdcLkwuEAF+pC1sM0RNfHt4WSQn5qvSB82xFNsBWMqC8L6K5/NxnHu/McsBeC
Mox55nvE+Fff08BH3Ql1ccdQ5e7TVFGgWakoN8xtKNYL7DMUh5etwCCPzmLdXBUYGx+4w86HttVF
scjsTsAXJbwhK2chRmBAHkw6hPZqczAf3S4lZtw1+DVF7z8WczKFb6iifCt/VE6szzkCfkRZQrJz
UZo0h/Poxv7tbJ8z2d2rj3XoOWjVQmbd8/0i111Zx0wxJDOhK2exlBi0nblQE6ERo6EH5vmBsNwm
/589hXPmKC54hUwQawFP8AI8RoaEiaHH780lYFaCbs2l6WD76SICZsj24PX+dNNa4ZZVIE/4bWYG
Mq8sDYwwoitH6guFerO4elpu5JitE4ciRngqTbW6rqvYoyhFnMxbNSrch3fDj6md8g+A+LNhwdEu
rJkyz9V22CxXwTAGsByud5j5GKxNmikSLSHKo+n6N9Svj7bnnB7VGA8zQ8riAzsMjtw+1KF/24vO
ZXiosTlECQsX56CY1xcwgmfgqyr1EH/Bj3PFwUEi7+8K/iQB6AE+0eL47lcnmOa9IijPMaWpSJG1
qTG7oKSXxzdfWkGvvHURLu5xTVYbyj+pc6UZlQ1JAGFh+eMgNPOwQLAsE5Rv7V46/GIPkIyZjy7O
J40fBQKaCM6SJhIN08gk7bBpSWLqF594Sh/5bmH1s5Xh0PkkzhaNMUe24zSjumoPHqOmChD0JSuT
wpcqbfqDmdcyp3iBjjn0j/399ZUaKkKdl/7lWZzrhV+zsdKJOy/gvfqtdaHpmQ9UANtE9b3zeyYw
U5IE5QcYRz5DEsxW16D5d2ZYjn9pUcFyJcJOFH0WtehFJ1riGHpg8jbbF8yU8vqYhzS0rR1zmGtF
UMfF/omaZB8sndfVpk2uqtw5RdGY6m7ktppOvaSDHtttAeQrL+hmV9240WsA4e+XQlgQTPQtii47
1jxCCwy9KZvFvRrjofMnqecGQQtBJ/Pgb7WPZS3LCM5okcJH0ooT/QTyV+pkvoRVqVN24u8OBImP
jJMN2wDj/+r6RRChxaE/fNuyDvfdC/PfT3JtGhxoz3jadzTLWjqk/7LSHKgjCy+H/sRNyu4cHvQ3
B4q8R2MSfGwXdAkJRkNhqHpo4mi7iEBdC8CuGNihAxCplZGlMVmKLwT6trya9N02+kxeMIbHvBZA
qnnt8eOxCOhCYSYQJsG06GJGXJdwt4DMPc2chhjhPzzr0JefB4sth3Q+gQnXj14KCNS7PXi0zdmf
NebBqGOa/MSft+TL3mywu6qynI+m03ZN/8UWhEbrdQ4+mWuv3TOAvWWsulZjzs5c5Kgxuf2UvQjZ
8JPlIddkjRV0yTDCot3BRxNUiyWF43DMUC/cgCM1l9iMzb3Kj1K/V7JX9F8n3ay9arE1p+Wh+VBh
rv04zHC927Y579nOfV6Nc3WHwvGIHb3ZWhD778/0lU7ipVjVnqpU7GmpUggBnamKSKOx+YxZ+nJ4
MAi07CmRHSF8HOKBxM4u0Wstiy+PTOkFaetuvJwhnc321QKSGcVcsfW9n50LhfvbjiS9arpTdT7p
ckQ41k81oG72fEQuvBsuSQM5qjluNRlNfKQ+sPeTow4OxoLD6ansrk5HAX/deHZv8AYj0na7nZgQ
DM2kZ5PPQU5E8Bore46uyjnxW2iv2elrYbULS2XgcjvkGWymHwMXNyE05YVneN9/YcGwjRF5Wk0f
gqhFGJIRpNKd+HC+gbqe83GMahjty2l1UyIoLQL+M41cYM8tn/R/8kMHcF/0AX6x9CSvkq1oh2xB
YeBjEh8T6YYbq34kLP+PqUAa35shm4OAQyWjNhxwiqr/tlb+nGwv2uMzK3/YBRGaj/0pnXmhz6Dp
vCwCtP7bA75USyVhULtCXQq2LBpk1YY/Vn22rFdUkK8LkoFq48r/qJCQYP/EMyeI8J93GiVfzQRR
FzR+AvEmpbUfGI+4gIF+cQwMdzrPYB9IW6tWf5675ANSYNq5elWrA0pDMm16eG9lA1ELWQnavR65
Bn8sSEKkKPWUmirNiVIKrNjvNsByQAzUhTa6ig60geKrnU9qYkBBpH/QgjTj+TOD9E65kKCMjvba
kvOc8DHuhNEZw77fkhKdDu+WcICijnkwq2+xDfGjgmrya6xKxaq+SKhxRxwei4h17hTKCCTRtHlg
Na64OD83fpNKGNjhk1ZWeElsAHuHj6Oke8f1nBqbVDEloD3TkC4HR9EP9x5VnzGuArbzcfn9gneX
O59zzMqHLgaECDKQ6goHTeawd2iSm0t6DZ+EuMCiuY9gcy3o9/knCuv1nQocCp2I5IiGkJttJ+ot
4U9Lz/c2nRqYGSnXMbxY8k6BcfSri9Suj6Ez1ANhyMN34AWiaX98KuuXD2vTdKSMVFowci6vHgsm
c7Bqc2PsB5W7y+1kmqEhCoVjqYyLt3ds1ftll6optyAgKUyoOVg4LXdhI9gwu8BcS18hbDbaXFOD
d0dHDzHb0A6hBvKs9iLg0iISSEv7L49HK3rsYOsTXtbS/FlzbenwysaJmSlgtBpeDmL82bQc//17
5UX68UVHhK2BnNCPnWy7tkLieTu07bIlV1XmNjCF5n+hPHqDKYi5bkq10gTP4gt8aDqhdPVxgMeL
Yv0idr4oKe9GX1g2uapzC1BTY3gySZtOlreadpDJ1oFU5/x2tNi9bWyyV5XvLUXn8n66p/qSynK8
ATvNblgtLD9vcdOlpE2M51OE/BuXMAQcqDcYBgdOysR4jk23vcxG6aQfwovKOFHwFpn5exShpeB9
Pe3HjnabSymAHk3ngJLxlm27RUVfyBSyE7xRMoMTjXUiek4DYsb40qlcryBA03Yi/86nQaMuqlGx
n4258eMLZBlsXnybhAz4/VPn4yjWsy8aRJBW2J2NIylhXAC00Icutuf8VAEsxQzr6nO5iantlTjA
mMR3AjUgBRCqzsr2QhwwYaChsVKPU6u3Vf7O68hr/zGHJ/hJRO2K8gSdDC4BBQGoKp9cRc762bQe
vMo8Z+gvf4XgN2HullwUZnxeEpOnhFl382Po7622A5jLOdnI1Nn4Zs9ewKkx3c2+pXv8b3rMGXFC
mwhW6oKGp7PNEL3MZnqlsFm+DnKBXJQoBa53mbAG250h+3JuJlxbO6Vg5PBqkcTPXD/bFmi9vslu
7mgn/VMrV9SOBMxbHOBCN8JpURV/yDTzneOVzx1QHY9e3n9TdqMOo2ryi4t5637HDLBVMkCbbiYw
RBouPWcedPonpdhSzbHuk8CIZ0I6vG6wq/U/xH0KeoCDJKNrEXh8DuiE+zed6l+IGHPJMVpPzoTu
iAIC3CzMGjeU+gUzYOOXB4HpBHAhDzxeF2Z+SlnL4uLVZNQDT+2qysiJ44hgHnXg4TBeZ/5fM7ka
5+wSguzhBqucRawi7ASUEBbUxxX5HRI3ty2Rp8UufL7qTvq0JIJGoZ3ocThmFm+06FOiplwEi0QZ
FnVjITXnwyQEFfmbNI54M272oHqOtZZQxYm/TNro3VCPY8lsbCSQdMg4HKVMgbPTRVkpF0OO1dZU
VzFERKHqzAuVZNFOpgqSFp30M9sAcmX2R+10r1iFUj+Br3GO9mGoqlhjPOUnpAp2aez1Ug018sLk
zeog52kIe51Xo3PQGgdp4d2YF9844QRyiUk3YP09jcgk43IXJgi/1HhoeEVVAtLgIAv/bG/LIoPG
AY5urFOsL5N7lzZGgC6h2J6MY7P9ovHY4KgPxGCepQL7DwEjEFsHfz+wK3KpvXZHsxrs3HP21pwN
5CrBAbC069GB6Ez4rgSAaWr89j++V+9YZdVK840AmPgtFUVvq2pHOjEMPoa+0Muq3Acwr6jnThdk
ua1QJaMUClBdylT4trSlqE/DDt9yjxvB5/EN787SkH0sLtrRdoH9dNsK2Dr4aceRB7ScZb+VgaaS
CDDUUCCoTQ==
`protect end_protected

