

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VInMykl1cb/eyCcstyHEIOqfXLtsMYAK+iioa3bPNZdsHyKysw1sMYrwKEQhbdDvFZxexFV/BuR3
E2V10xNsGQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cUXIMbq/fNZtj1t37ez/ki7n1ShEuWgIH8yPxJTOO6Au2Dmq6/c17dbZtzNOPZ13Y79JsIBKn47t
AJMl7N429e8DmdtbuhhwCbJ38cBiFdxfH1AfVZI7GGjMAdNcJoTCbcfH0JfWJ/S9l4OVfdRveiIb
dXW5fh7twSl61WcUJpk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WHbKIifiSnVyh9VOrHbsAOJaiYfa+g3aWjT672CoQFGtZoHYX7lHrwPeDjn9R48BpRkqqMyy5V1E
kZ30rvMKCifKQNzf0TevcVrl3t6QqBIPZj7dsFAaWjY+3fu0RTcnya994wdnAwJ92k/2t3MWJiFL
8UCO8DDPNY0Xt40qfK/53oP7zxzhOh1lPvsgCruLCaYCAr7BplNWzKtgMfwt5ZUX5jp0hTpI0y3m
TFH3zhFRvsKAbe3q2U7sLVIx7P0al79lRmHpf3nBQ8JKs1WigNl/h+LWFmAr0nyU052Sl4nQmc1V
27CTe4+On+Y4xMsv2u/myTqMuXN6bcLrIAsu0Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xu9pS63o1o+cY63azBQM+vsKaznHACPUqoNT6W0vN2jhydQX/sdcqaY0W4LMPjU8g+1LDfLNYA4a
7f9gcYfJbb3zaKr5Y84jP97vWDuvkp0JSopB7FwosaQhgC9ZFFZSHrzYGBzwuhbZMni9A5RqvV2b
bQteOe3Z+NH5ROjD29Y=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rwUkytz4o3nSG3lKXYNGBGGd6NQin1yD4vxAFncd1x1HAH4uRN/6Csj8O1eFBSdgBZrbzYpSigyS
irdheULjGWq2hoVKG79mqHugwoJaQ+RWNnILZnDjYUeFGEu0ddu39e4LQ3yMfBCfQxRQcGTVly4Y
EDooxEh83Mu9Wm4Uvi2+2y26u2oEwtbjgdJCVoicm+J7JrH1l744lVTCHFaZPWdZupXmaLsbDTF1
IZL005EF99uQ8TMXRMkzqTgTLlajCuwvHoYLTNcLy8P1f7qEEvcak6Aw3luT9m7/agpHKsss3X26
y4VegtaqqF/A90Z7VEb2715YgMpxzFEM2FzMyA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15264)
`protect data_block
iRvatxsLqWy35MO6ja2ADE8GSZ9/09178OAzRVwa7N08ayGbjnftKvIPHxIa7ONn/d3dR6Z86Hx0
3IsIZLaLejkrIc8QeeDKs5dNTXBC+sFB8Sveejv4a77z6oqYywnDNRK7F4IugS78sG2GCw61w0Ix
cMxDkCTXhb+W7tNdkxZuRAq9sDeBlLfAyLYTbJwQ2OfMvw1+TgtQqDXX8gEkC+IAA+Ts5C9cvyVw
rO3ssYR3pq91onKWwj8Ap0oxRIwhUleG1zC+q/Y/yk0l7w9xMC9d3RW/Bt6rQF8Qy2OfdN1GdUq/
rDz1vO/tuq8bG4XQYIer+GTRwjvku24IERXpLbd72q/GA58xoXssO1eBKleb9stpK0E1zTz42Zo2
yn51aoWN78H2ztxvvqw1z9XXa74fg1Z48g0hDDdQKFsoRMoYTTSfnM39bhTR5p1H6dXob1TN6G9G
vlYSRrCRyflhilvJZYA1QJAkLFEuW4AAVHXxCMkxOK/PM+LeO0ubQV6IAUi3TR0gN9Ku7EG7QIu9
3n2P4POUlpMj2yuUIL8WLGklVtRpo8oz7kidAFq5s/tUcZy+/0bTy67w8nraabEKVQ4Mp30kKxQc
I8k+Gvcqoe0ANIKpWbGYX5ht7OPv6eFtkb4PRA8ajzdvSSEuDeCilBNFOXFBR9umzcauPik6UEwS
NSWHhgfxE5TGOpz8CYO2005P1mi/4nFWnjkwsK8FsskSL2u3rEFRLHJoT8ExtX45tz30aAZQURgI
wxX8OJHTuEWgtffW+GE5bK/ifKSR+RUuGg2AakoPXF8R7heKFUc758SYxdtxNQqYxrQRu87FGzBJ
hF6Se7Z8l6MDvohhk+SNBRtCXbvTF7GK+DgPJ9H0pfmg9mE7tfwoZAI/Kgot8d5R7cObw28clSEl
789cTh/7U3PNhmPyjU/h84DTIM+wsd3vAiUdNNxsV3UnP5tDqYwzRxJ9b+wfT1p0WXnMeKo7hEvF
H464o1fvB+13fAL0/i8E3n099hN4Q0noG+3L5ZDe4b5evqdeEM2ptsE0l06+EEBER9EFyf1Hjx1f
NtdR0t3Px6YAuRqWWbUJMQv9n7lWadXe1Kw9bwqGhMZM0CTcDUvX449zDpAqn3opUF8TttevJmiA
rkmnHmhwVt9qH+s/p6DX1jJt8rw5alvFUhinffn5E+SprRPeW8lUIx2k1yuqt02xUjvYYmVV1uEZ
yP/xsvNCu5N5ZOQDyRwPdw9hzyjTG1tdA6yelcgZAlpfV/SxUhw+KxpA1HtYuMIRIkXyyrbixMeo
mxK1b3z9jA4A1laphaKFv+giomWj3BdJXy3saRGhcYbzXg2fR2bL1qs0I2ueX+a6Sq7/KYURbW7I
gx2+kBcPfKp0vsZrO2OotdUJo0KnJXU6HaNDL8rSd4cN8LK7rozskmc9zV6rwpYBDwwmAbwTh6Wu
gx//hgGKs1wUw14xVn5CipGzeHkTEJmJNvPjv3vDTVBMnrb3Xf3HKOix3MP4RLVnLsluO7AcI4N0
L9+OHn61WrXel+GPpFAjqEAUoy9fPrO3s/5pDdPyJmH0L9AInEWtocfCngxoQ3UDhMRiB7IQn4v9
cIGynegnTv8jy2NimZ/qo5wd+zKtHlN6Ib5LgMOsYDXXT+1AcGRhmkdBImymOfIkdqbYYF6WW2gQ
a+KISabhrzPfHigGuKkijVJEIZo6gyEOSY3Kk4cQq8GACKepmh0c0HskSpbiupuGsDAMp/jT/4qS
k4MTET4ql0Hl++x1DhwG13bji99e9OKbPpYwkHX8IAdg0EgZJajETtbejcSDWUjQS5SCSuV4XIQx
x7VP0XIVUfdKKJvflclrll+eVPN12PK09CYL0QMhwp4g3+6V3Io0PQE0mHvWnvdsWsW4GlBpIx/t
4N1FaUeJe081iGMx6edtMCTBpag1QIK5pZOyLQD4TLodogRnvFsVHcEiJFzjUvWx8xrcSDGiwkup
/16sL3l/NVl0bVXVZZaZMUpZTROJzuHcjCm1h35pkZLju5eqz5Kp9s/8NEIvXF1XspZffeQteCjW
awV7ks8AGZLx6QR6COSArV6IMKaPyr+D7BRCxdy+ISmQmLUooJmgepjRGgnZOZS86hJLlPiTQYMU
72frPxmioHU0do0vL+CP3L6ok0NuCDXnvvaRhZHpsv3I4GXCsKlG+27cUQrYfb8/NTktElGo1bn0
BzgL+yjQbRUHpO4HfH0s1xsOYJErsDSYkKn1s5zoHa+oZnIJlmc7jZ3pZQ3giH3TZ+EhTZA7zaM3
shJxxEyaJsikKogyMmgoyRNy2QJXxNPRvFB3EpAATZ7P0iGJ5QJYHhEu6nsBD3rViQ5/JE2aB4nI
PLoBjcIuv+dUHtc96wYSaqdRi4ndAnPz6FmGO66d/Vqw1D88taz8Lsm8Ywe2hrN40h0TJB226SZH
5Iuhu+08d2Y6JjTmhe8HzKC8/Dc4O7rILSwu2dof1VcCl9KKhVHWoc4iu3faBj/2TXFIRABSYGpO
4YaGs9kX0NC8wEmCuu8hD6TQVhE3LQGllADkxqa8pBlHCInrbN7utKkdwklfi+njRUQbBDQGlGdj
iC1ls72VnAVvsd+DCUE/QqV77CI1S2gtGs+yDJRLo5h4VeJAFBdYXvliE5vXNIdevSZQEcbf3Ikb
oMFz/m75vOQ+nazlefS3qrMC//28OGp8opXVbQI47mPR2egFyw3JxKpNa6W4H3s7WtRyDfwzGBAl
L+1q8vid2KY5n9FSwnw8EZO7INlTAGIKGYg+OXVnFTHHEYB5H3i2IkafFnA0HK8IV8WVGjEREL1V
ZopyZGqaQ52u7Gv0yHfyHO6HXD4E3jy0IisLEowyWpZfnK7oTNTJaynINusEvaXAtdI5vpLxI6iV
qimuzhJVEGoQRbtIX/iYgQV2qxd8FlZUloNf7R4RrsxW+kOX711DRVYcsuVB1A+Z+ynCOYAl0/Os
/pNrBzVY+iIEVOHE+7i+K0I3LpEUDDreqWsygoP3taylObUIOPZbNBAmrCMgcDkDI8ik0xmQVBcr
+PwNj+22nnfSaGxZbLAH7GQ5+u1O6zHLyAZnLsQjD1fZu7Spo/oXtA6dcRrIf3N71LQUz4BB9k10
xhpLki+UmGRT9/aeZLEEy3RuEJUclNmVSGOhTTW9+DAzAzli/algUQHyVsSr3jp+rboMcWUlnw0E
UPho/GIMtVTy3TdlxElv0gDQZpa3BXRnP39iHnJJkNIjm1Q3Vbwl0Jkofy/lKoi7v5UbkRSeZDJX
e0k9wh74QaKQnmOKc5sWTE4S4V0hLPHbyoln4ug7RI1mBKb3aKgQTI89yrjl+gBlAvsesbpNah9L
EQWwIGfLpzSp5079fsPVHjx9LBAZYOPixH/KDBhi2eKxQfrfwON+PmM4+pZ+N+rg6+T6BxCLzf0M
ZlMktnrFiK4RlFUlgJs49JTtc/o5qbWVT20tOv6tMOqIl4E8O7bGj/0aGZzzxPvQo/5xB2wB8LiU
eWwJDZWH3Utg+yG7rE0m8u6unHHUSLHy4FaanJO6JCs2w6emCgLVOmv4fEymXEpbaEay9m3jk/M1
Mh19FDWsFM6EjSUFJL7q8WzgETQ7hKjSOxZ6swCa93CTjDKV2h/lm82z2yLqIWeFfJ6VamdEAD42
fiYERYj+9wTnjARnKxB4cfxu6aoi1sOrfM15QhrngQBSFGvyFw0Yi4Aa0lPWvDkZZ6ok7PYZxu/o
ESpDTigosKoEuTj6YXac/Be+xGlHYCAxhZWnzqrSaUxlmN+4XAostPp1ngY2xQKbe/WdmR+6TQeY
lIIEpXWRkeXHLfxQwHV7RK5SSl/8ZJ0dJ9pPuBIq5yYwD8w8QyOuFvneC+fkBFWsoqgTWkTUuk8I
I+G3x6aSMj+VdzfOg7Pix6yXc/4Ebo0s1gCp/0enD3CzvolBLYW+sQhqqrqJgaCCCR2rU4md/fOW
SCD/QJEGeipfxi5/qDgv9Kk8uX5c4A5caUKWmlenw/jieSPfBoHZ/D9+yz4ySkpyp0QldSDouNI8
R/622pekVw1YR2SSEK/ruRqBXJhRqnL5SMarwfSYE0W9Z9XyPtbl50gvOrHt1o8KxxOHhinSalFp
z9psqpkKULHn1m0DHEz3bFyktDhEDNMKDUU2uD5WBHMv2EAMbDw3HcMP9wvqdUh5WpcH3bHkarbL
GcHGGle3E02dy0ptBzb7SR//7LDucRQIa392cLleGd8NV8ZAXqr4gIe7meq32GdWxGClT3atvOUM
GrfdQsHkfZxG9vWU3wO5uE7NWSDYGZtaYYUl39u4eidOCJOOWCn+Ua/X+fOz2Qeap40xnPXddPMk
8TrCLFZCBQ9V/AK24YSfHDdciHDYoAbiRJmLRCikQcmCpdkI+pNIjxTk/mbnjNHl/TCCggsL1AJb
eRIvMawmjHf0e9sooxca89maAkM8N4nRYeMArPevkn93WEvBNE2QSHc+FY4NJlbxHZ72YmHS+YTE
mJbFTXUCH5lvndWjsomgpEFNZI88e37qWgnSZxU8uMf8L8DWTNxdvkNYTYEVE7Z/AXFFFWhV8ghy
QyH188Sm6k1FCN8oh3hLtAH5rTFhVK252bEVq7ZxLWAalrYhPxcJ51sPAMY5D4fHUnFI8mwD+FQd
Kp0V9IAtOc7AyJKncYGt/gEengdYpbnEkDoc5ckIYadrInuZ5gAacq9A8MfGPGaCsLK+EHok6t0n
sMs+3tY0y7b1RyV6ALVhr4vjnL00XiDITrJxVH/zVi/PcZcQz4P4sjM04oUtJPbDlIXgRblCc61j
ZJyXzVuk8J4Hzze/lSbxLyT8PJ72r90G44I/eVbzo/hCH6fOJefnb2QVN4qA373sQUpEd7IeDngN
KlvN60ZmbyL8ya5O1kvk/9bV1PQ9GvHAbarDOXLb7eA8iA6dw7dolInlPpMsEGM61lEclpOediSG
N7hklnn4Edr4tgpBKnW6AZX14yC5lm08MjqMR1LOHTuO1Ijf62mu5DwJiTOfjNe9DdB4bD2WxsF4
Tq/31Qbwa6V8kepr5timp/HlYqJc08qE01iwO89tSze+tPnxhofAJyWDJ176tTdN/O6LeV2Cfq/r
SGGzLiAYMqwNx/psSw2c60ur5VnxNg919mY1xpUcbq705R86qSAwRpQa0+eZ8Cdipw7NwrP7dScH
dTUhNv9nK0Aa1lei5dyJ+H5jjc0wQrQuOsqLE3lWCxVVuACD8+nNJuvUJ+AS78qj1in6tpzCUVLC
fr6ON3TRANM9wMJGI+pXWfKDZq62obrjD1A6kLhrdg0sX05Byurpy85AeorCsuUSBlD1hrswFxKV
LUJWOWwtU4WIJPbhxDSkXBGFIwTkRrIsP8NOWVjeJRns3+PWl/c7RCgBiTEj06DsxpqoX8r1frOX
ZC07pFI2WBbES/rgUhOXAr3wp+iMe07gfm22BQwM0Pg5kiED7qnRuXtsrXZapUEoWbd6H0k1jk+I
a25yIqWJouIsyB4RVMKxaJUdjL/MnfIKQG12yvH/y1Zh0EwTBq9ujlmdWfdoS+AEpSAwEfbmbQKn
IkWrR1RgR2yBxKePBaeSaRD1g/v3Kbyn+npMfNUSsEROXX9tlx1vs+cTL1ZllmJW6Q5Ia8P83T3m
QWHqZKEmzZ7PnmaRfLVH7zK2Xl8Mb1Ul4MwcMEEmWBS73cIG5L03eJqNtYkME0jjxWcOj1XZeaDx
A0qXC23yAw4ZtvCMY4uT+WuZ6voQ03OQwPP56FeQjiyd2b6j0yRh8JPEQcnzD7DUoa2u9KNhstkj
YW1OQhHmT3JsmfPlKmBhYIWhhf7DnZirpZY9qbWe9iCeQXz5Ma6Vr2BFybG2db9S4inp1s8+0ZGE
t/B0er68F7Mcp0aqwZuWhdXBrxfeDo7hvytKH/cnAKrCnFb6FHY4R4sEqHrK3bUlj/sHNmUzxw3w
mOHy9b/VZAlIEkvmrxfLSG0GDjU51YSvTerX8cDrd5313WcJX3YFV0rtVWpWIEiwIw6hz8/CqTT0
iRtYLHkA6wj8UQhFRf0jKVYW72VON5ui4o7bmGhYtV0i6MKWxtnS07fgyrvehiRcAgRhuUqfgzOu
k6xZSD6n2WJR0fuX/DVDP2PXfc4k67PhLBAsAhG1htxQUEWEeStAYWAHuRHnXCBA7wk5KrzS7wsb
NW3OsYCAa6DuRjYUaYGnwAq8rBDFf4Mv+6DsqWpMcytAQZese7P6R6Wd+lcRgX8xLT8BSQdWg/S7
KLG5yjlEHjUG+A7jGQXKggQYHwavVsRjKsa4bycBytjRAfeBfMWgEvpsI3sPc1G9tqV4BXxLR6nI
nO6BRwl5fFDs3fKeXQUmD4Y3siut3aYFbmUw+9SohNt6PfogVg9Pnyb6M8aQaswq3zOMQUAV7TFW
AAWHgGJnZHGz+GnEp6+XrI4nDhhvi37N5LWzA3pMLBKQzT7ltgEC7zRYnVbsrCj4ukxNppC2l2Sw
3e2JtJmmF5PyV2puSN+KyyBnWmfds2Cc+OSIc1Ib23vJWzKhYVaPF7MJGZSkxEuKcmoYte+gqUEV
rkW2KDN9/VCct7D9Aydz55g2HhdRRr6N6VCnVxP1G/dTVyctPIqztoNFmCuSjycnF0/7XpjA6V0m
A5MUcx9t8rT0yNb5+iI+rTrGIiqtm+sXL1ARI+D1kQnoauXTK/dtQQqEAJg3Rmey9R7LAK5jyQtd
m9yN8+MsyJdEg4CpW+NxbGQvF6kwj0nhnTculDF+DL5vS8hco/IO5pyNRNjWTcJP0gklcMsvYjlw
WoJZ8tYdozfzxK5n/4ZeH2XjCj5R+nTKWHRQUnjhzNyssYD21NVH+GXNvsr3BVRmjo8YRfRSqDFd
FLBWIVbI8XjHb6+OoNgIxBxa8ZHalv/FLhRLbt4d0fgv15oVnzvyh7pYafNv8Z6mKvqChiFjtjd0
A+OXHguMM38/zPqwtjTMt3vgjr/2w8qR/CfWOBhFzYZtGUNL5LnvHUxXQ3mhvp02YdrOkinwOl5t
YIg/b/6nsAAny/eBkYI3KamdVWn00Fm4FzvPGiPY9Q9QUTr+fZ3Got2wuJOR3OR4MheZQCb4YY83
9x0uiIDcIaVxWm+sqP3Ud5aGKHPmX3nhHd48VYxW9FLjUPikOZlvormPWY7Mx/AZvXX5IRTk30V8
SS6aj1fWcqgW8qdWKC1BOo/nmnqhdjeVl2D1BHekKRhdbmruda+rr3sko/rRfw2u238oxpXSp3n8
t5+9Svy2vVThx9sZexm311S5f/uKgfQXuSIr+JheaAfQRmA0Nnq6dHjaSiMNG6H5hdzyQ8YAQBEg
hsZ+5GApzPlw9RYr1TCsaEoB/zVW/o8fuOG2Uz1Uj7K2V6svT75QqRVV7RdXDVyQae4Iv+7gPnCH
hmGdrYi2t+X0yZ38VhoHRG8gXEWPfuoX1dgfnXYci0IdRhBLpxBwUNfC8hotTodDt0BYnofS2+9Y
ZmiwixTdz2i182yf5RlX0P9nxj472D7hOhfeEOhEgBV4Ca25nqbsn56Y1APGpaEyww7Ly9QkG1gi
8DE0FeTdnBz0EvTAwe8qju2VNniZi51gCkCC9iBhD3lBirEL5aSdjjCpCfakTZXGkkko+tTYtclb
52CIn8r7AU/VzP73mhE+CHFGWbL0Fpk8GzL2onJXKGe1bKHmpL5Yqm2eDTJ6YjMS6JK8cleepr3i
pPWZiyB8GYk6gMRLh4t1Eo7JWAbkxHhfsbRUPJlffR9Ku1QPNkDaJXSm22IaW5G+iSJq5wp05R66
E08nA3dWxInwvGKcthFf8l5gZ3DM5HbiriXuZWqBZdWD+50x/7aYysWjnhI8a8zbQvFiV4tNE0xY
1Ger/KvtvgY7z2XCQTjxChv45vde7VZ6K7VljD2utkEWSqyju29FN96kR53SuhQMQrMmQNME2+Pq
h5NxT6rHV12d2HhRAoinFFdPH3DfLi1Yir67YVYZKrJpt+B/UNltzWSNT4Z1yE8zhx6wZ13G81AU
s3CVbryU8muXb+bDJM5zeIIgyTHu/m9nfkh4kmhcwZFcHQFlkp0SblIvSzp3ebj2iT0c5j0jPmrz
5Py3K+FS2cfKY625Ibm9+Vpquhq8hbjTXMgF3eRXgQLZ/Ion8OeoH6xfzexxV/eLA8JeDpDHwzXb
wzhgaGDvDiwVOrW6NR3ialpGxLL1eQCm7mcn60LmuREivA5s53FoEzdjaFHUA9CH4QZAazbua1iF
AFf7duJnw3X2ZBNGb2C25hFdgh/fN1Z0cvD2dnG/HKcmd+z4G2iKTIGQ9xP0BcIBbhJHIXUfEmGv
CjwtYDHnrzuilkapw5Z2ea4X5BauZ/PoeuMDZqHR1/2znIbRLot0B7X/0NOfM1BCydtNXkLU0Ord
0SD5k8zZ1d1k926vqS6Mp/jju79NmvaTUuYR66l0A7iuRadlwq7d6DoVlIC5wnOd4SRNKnBOe9zz
GjoV+H07oMgph5bFV4dbafei+HG8gZnY3gtOmcGB8Em6VOxkVKoPFhzV0p72NY03VXPZCHVyRuFN
4IP97DkbLGaSTzmidt683ilicx52vF/SPfEA5b+fCXiH/0i2aRGraQCl8tazXKJPGVRbSwqftpHG
Vsch0g3sVQbD3dY9GLqa0Oq4Id8sPGO7izd6cDyb06jPafVxB3vKuHJoDeQQ93IYITWUj3or4Jau
V5EQ+x9HU5eHsoG0N9gclGT+I0FU3KhXCE41LPig8AYZUAKCpdlTEF/LoS7DghhUL++hIiRawdQq
iqOw3SZteTbteVVKHE+kZwmuE5yBNORC34XevhKCkPOSq5diYOM2gCbXG5A6xPD3Eb24hE0/UOiL
pIW15lPKdxyyHJe14eeh+dpT0UjSbPLhUk5F0g6qZoyg2Lc3PcLYECI423+mVBnojb5a81o00SJ/
JDC2anMMyrdLaJf40SxeekeHtmj0nSbI8+uoY+wRsk0+ZQlUNAWMNrtM7d1YjqHvD1EfOIivhdVc
czFceb52Q3H+cmSXa9FOt2xtWsKAzmryJ7b6YJMpZ7ZN44WWV4A1lqSx24CwbxjUd87vSo6Zmmrr
M/8/aHxkPa3ruI57ykLzhV7tUmaOQytDElaSgLid5uNNvGfbtifQuSKbonfxsifLsiQg4E0CKaiB
j+ukYB5dtbt9FpuKiurrn/TixffKxa6yrZDBywH6cvKLSXG68pGog6ZQKmAgK+aVGIFQZ+zWOUME
PZxn7VkGdaGrPhmxlPl8mrizKm+LCq27HnvBaxwv1PbxCmmFVROnljsMntWy9q5MAVN8ScM7XLZy
k2YnVoFw96EccMzD7bLXHnqoKpdEdk/0tv+tyJfr2/Pfp7I+C68CoipKo5Ut3VHGfY+WoyZHHWlw
8jylqkBXaA7kfFyv7u984TE7UzL47VGw+SRXY/st+Omik9sJ11PCnhryLdT67aFn6JsS6ZN0TLEt
EdqIGZnP58fpLBb3p6j38j9lw0CyWbyM5IUTlIn54mwknLp8BC/Q+nAIcE8lJSaTuLtBDs29jMKa
IXoLA7AwCxKMdCc9YBWqjSQIzlEpquff0qDyzyNtaEzfGhnpX7TnUi4g4bMKmtJD0/0HXv4V+45y
hUU06eumilSgtIJktqItdeTfD6vMcmG7UeAZq0GPROgvhWekc8gB6+MM6QWokYzo2iMVrJ3yrbom
7juvSf8oMydp4YsefiCA3OQE7P5Ec6l4W5tfVO99JV9bGhMD7SVGwVhyBbVV0o3IdHVmsZC00Pd4
zNKcREjXkXWkoWJi6FLFYnmQwKSSS+XXm4KsPITO8tV46q9Q5Ueqg10S1/xj+zJXXXi1BIqn2EFA
JnI22qZA9iXGQNfi5F7cWG8JT85+5YtiOsgyRCwlfV44/zViv2tDnWDLqQyEuk9SulPl+qjjvg4L
bL2ElIkynKGRHHc7OkwfSvPwgtAGS6O6ay1PHOJ0nzWebPIcWDMnXhtoJOa+iGT61yEPqCYag5Us
/K09pHZwxeuH/6+xvvrr4GQIPFqOmPtkW5kXuLI2hnHAdz2f+uaea3l/GPNAJ6IVapV/dx7DwLFv
Mo4IG0bJvTjyMKvBZlb7NOe4lwaFHHNkXHsxiadwvl5hCU50oVAjPQMaIyUT3I1oF5OZg/73yIfx
mmLcIPkZ/4Fu7O7N/ImlV+y5Z2G8ZdyQFARwMmPv2oJHyv+nAjds+/RVmOmtJ1o/s26YqgaPIeAJ
4+kJ2EfsLijlWXs8wJhqTn2SeFyEUdJl8cYZTDSMVZGf52ZA0ouI0U+79/3HmthAkyKhx6+Qldmi
nckOsGvK2NZjD7209cowl5om2J1tTZhw73Ukucx+4qNe2QfKuqWUd/X1kkKhrCKstAWNyFg7mx1S
HW1mWgbyLDRD9/pOBZrs4PlzsGZmWN9cReHhDE7/xzUXZSynEHkPu1S7qc0dfOcNoA00vY7D1BYk
34MrvpojoZqmnjQkEdfGZAemgyXKMUMYjyOkY80qSysZ9ooEMQSU54Qpr0sg2zyyA015oK/scy5a
hI66faz/NvZRIc3YXw6VZHCXUkoO17ppnixZ++nbDGU2cIY3lmtZFDGDUeKa1spvMBai2i11LDyG
j0BDmHaKu+108X/QOLfceL8R6rl5lXVu6omD3U7tHmYYmVspNPtxsYqnMWfELVl/B8d7dGWUb+Jr
8wm2dQm6CfO7wpe0uCOuO3IUnN21QKzjl7g2GnEDM5l1+VNNiiRQQqwchl/QYlVLC+lOQL7l/hSr
VL4BZchrtnxU5ZGqMo+GTe+tH7mItDsDSXQuWGsuJ2yhkCsx3Tsf7+Iu/kIQo8W5uWJQajyXhhAU
JHdLUScwWsjU7GUDZmrjRux5UoRZRUpfkrDqV1o8D99Eq5Np+WX/mqTqFwyTgmQIGQqx7n2CLTic
1EuoY5UierU3cbGMz8VmHs8Wb59gozomB+ovqUxJLu3JRdkkgq0Q1vCRbgr/eS7W7oeHmYT2Tr0w
Ucf3pXOT5TS+72U16EDhPay3BtO1S0pmLqfGhWgKNNDx3ZTT/cAKKAPLfStiBqTzfIC7K5Cj6Cfn
ihMmAP7jxeOGOWQkOp48E6jXzXu8aOpBzYgA22032+VtUzYZv7l7aGFik9W+hbBJLsjw5SNDOho6
7kWYbN6MbA36B+LcYAdZ99Nk1PomUYlaNCekZg2MGDgGbafSE+j86UmxMdm6Be8iBsqBX3+FovI5
mQLFhEDDG/vmpWxYX0bq/kkZJE4FzQ5FKm22MnjVR91GIVEYjkIhXEXYGh8JWwiv+/C+XYIxO4r+
oNC73JbeR8vg8EmV0pTlRKmhBhWL8jHKbS3Hq6+F60/afHtSARnKCGOPlHhy48A6CoILzybc0ZjA
iD38tg4U/8rTEeexkhTgEIGybo1dLBhnRoGN156ANfLawDtbkVFmCSYmRuYhVewfz58tcqobWgmP
IzSiMLk1YgtFQiwH7/syHWZ8Vqm06hjnf3PXuwneRFEjILpAWAGvlsBTwfP4ac9e657ubMSS6D+a
WjFpQSUDybKwlNs8VHPFQ3emzrU0Ak6xhGf9XUJSipEmnRQcsIc7hnh2zTakz3n0F2VZGUnWngyX
rzd3M03glokw8afLLxp+WIwgO2X8FGur8FzzOhX4r4eVfkdxYZ4zOQKjr0/5CnXpRo4SMMFxgOpA
KZnTh67bATINfqiv2QCvYAIwZyJzjXJQd/MU6kBY2ezP8zzXDU0TyLVaJqiu80otqeYUAaXBpSXm
DS+DPwKmEex21KGBMRAk2rMHnrioMdZj7sKhMrx2/ws/bwpOQy+pyw0Tdr8PxPngPJG3WAbi0Asz
lSY2cAfakgazCEhFp8y7Olc0cRffN72gDtUrLSCBz/hp6s4yJi79hRgIedgx/lkb3NllQ3xTPoKJ
ilxS3pepUzpjPf637mi4wyMcTkYX1KDdhuFUfm/SduUkBS3389wzliTAEnNZTlBxV6sSilqZKfpw
k7tl8XPVcbfm0JnigyObO/veV7h/E6mVMPNBZg/xAkHyBscalSSZO0tikZmB+YPSfghvG1LRZX1k
s3izN7fntcGBKujxjUpQNJnRRpp388t2sJrVvhx6K869UYyqgHnErMN3GyhvVeVPRj/Rwjk/zUSg
AaTL/EXeIjLkuGIUkbD3EA+A9qmrSA8VaEUbnCkhSVfbi6JrL157oOds5R5/kD27Uy7clkM/a08X
Lc95zcVym4w2/n/cFyyBw2tD86l5eOkv3kBArbL+09XaCNf/RvvKJ2j40t7jS92ih6PcP+9SC0a5
/1LHw7dUPdIuQ2tu7PircLckBKYbkXkTncQjnBZqHK/QaL1MU7pI9bp6bxCC2eNxEDb1nshB/WvQ
TJngvCtcX2yW7ZkBuv6R//7Q7i9f89Qc8CAvLaOrrTXk/vuST3YUQhz9IvzpJdFPKQKNjhB+ME5Y
cPa+bnHVbDW0KuN2exr0V78joLza/Xiu0NsSPIsPqEWw/SP5ulF7usLjCGGCy11VkRKWCvI4UavX
jNqiyX6BQ9uZjBugQ7YnBlqUQhxUFBSCxqJhbkJXzCA38+K0ZWksNnNKhuL/E/pAKQQ/X+sc5kc3
OmsLzL//2/x/L55oNhZdDpqg0CoFcGpzQTRA1TKbde9reJWV5UpjtvinymGcSOuG4WPOzRkPTP8Q
Ywa5c+a8WgLiEzltlve6LZ7hbXokhLvsitVakfDmliA/IZtni5F37E7dLjrLD7za7ZEq7SJ9Uvwn
rwXjN2uKTQq1WpkibIfvDZy8SjuDvoIrld604/jbO30RtL+vO+TuXkfSakCsGms9K73o72Tra8GN
F/fmoxBb0jTMCH9yVC9b3hDCIXkWeSHpI5w6nBLLTQ4mQSBL2BYY3ryILxTfLDoIpXvcUI1CAseO
G3x29yJLxGzuoman2ld5lyM0GwJjGtSw0sRLR789Gs2Kv4UE7Y+IUH9eCFJMGbjnxwPaQDqXN/rZ
E1P5Di6HgOymGpPJU89HdjNj08A1oR5SWy766TVNUco0ldgCt4uUY4a+mm6H1jxfLJM2mmVbHKUd
WDyY1je1ftK3wDFB/Rhrw2hywRRKkTllWW9jjQI8rptSNSCTG1Oj+aQLioLmEfC36rygMlsgnwfO
5b0cuWZNg0uqYdhcBpr/JfdHGRsKt2+yc/X3FL1FcQ3E3D6/5Df2OPLU1GyZmVgiG5MKpV8PsfFe
b4HAmI6HcLO68JskF6JcUFjylUcujNLPN+T4inRqGy9w1vSTTAotF/cOyTYfBC83htzmYHJC8p1A
jRLRwx7+uFM/BSlsXYYJf7dQBbflrHNXYvHZf8K3ub83cKHvtTBoNuhnCk47aqnwD39ranPBhXAD
Q3aXl3QhGXUF0c0lvAn78fxV9xo6C6BL1lQ5U5a4MoVphCNzF69m6nKie0abH0+PBaLIvMtK2fXD
DrtAOLFQd2T8CGKTinH7GTYiIeNV83Ca5JPVw7Rvrb013jcC+BcPlCErF4o4sAd3a/dnIXvD2JQt
oC/xBP+KnO4ZZT9pp90X7UlZXAECkyaymrSprT0KYbbi5oeWrgl/rraPk/LZJoiLEjOIbygx63Ts
lxndYKPqZP+IRifPSTNY3p5bP1UzyKXxXTSADNbDHhwyvBVfb51MLyOtAR2j5uBmCvun+hIY8N93
wgXlpv9EhwZ1xxmoQptOQHsCs9kSAktvXqKp2yNboZUGRbkKnUxQwagujlQXNSstCdZde5U3M2uq
LCsYz0trxAcGJsE8o4ZyrHR2pAWcpipNjDytRVFNlXsP/yp2j7wU13yzgytpm7SC+Z1wYhU6568h
w8CrmddpUE5n5W0B81gMUKkWcuU69U3mDyjdRlUU497ejk6z68ULgZhhehpd5ZydZzsDyey34KCA
t2ITOX5HrD+eMV+m2b67FRp7WpWJoFpXIF1tbh4bX2TkfasGwSKjy+yDJsSnJ01fPwy5n28C4Lfr
gFIwrhBmhLMnOOnhqbGg7+2701f2DzXjvZ9JMGUx4EAHTZCw3qWTjZ5x8iKDjlRlpgiWQsy3eJbc
E98itbsgJJguuKN6h38tp/ZsgSn+Nduna6NvgfbyufwDgHocWUfYuVa69QTO2jh4SU1FnEblEkJn
xpbs8PWmLWf+rjUdqX68Q5jSpukkm3eua3I8UOhwfGZG9MiG/bUhC+/xA8M6aQeB/JBTZ28FXEaq
j8SMbwN5nAmKDsCbtn48ud9MtRtfln85m/uck+PAvcncPe36dLRgjQXgY4e8wM5VncNWpnA45mKs
rJhL0d8rMSmOF9a/F5c2Wdm1i73BnnmtCF3mnmfu1uh4Bxc3FWut+PgwJfJnAysMXiJrHkzTDeTe
j3IF8YtiGEG7Zd1OphB4qP7ZVzMfFlxdvPhq05uMhMM1wuIoSKbODqyi+navxYUd/vFVX5icW9bA
8TjiG3w0MnzeuTrqcMiTBgO02hKWLm6jVbzabm8nbH7iBYM7ZFN7SpMAjy/ShrwApzIX9lgiaPmF
rBDUdNVYftgUWaV45JPSLA/1e4jFHiCd8s82opo9gW1RCGIRFTbVxfV4PeFrPh+oP/bfkyvsP2xl
xCE3JIbYH+oGotKQvWc7bOukWY0iA6g7V8eHQQc484KhTl21ROdP+mgZFgauN81cN82tLHf/xK65
ZGv9OMeszQiQZ6JOJJYSOUVos/Jz8IlfBEzSfUn9nqVOoZWbmX4QBwUuKuUrG3KgPrAN7HJsB3zT
QhBPScFdQXe+llFKJTSWoSAeAhojOLLNT3e8rE1G7SzUeMqGjRIgy624l3c2eyYDGdsdNP6FvNIR
uvl6RARdnGmT7fiQfIKfdhFk60isJKpgKv+0sUKcwYHnmdunNy6bTT6HzFfwZmlbSopLfB9wR3Xi
UXrs+5ojuifhiVanAm9dZS9l3g7bSqQr9EvrqfqQlcjWUFUaEEVSVWsH1UqKBYq9YAC9Plqw3Xe6
I0hSpyuY3erM5ynQ+9GJtikHngxYt2gtdfcX//fsyFBUWAZP9tvO3DqFeKOfWg8PjPdEE4TJLyAV
Yb/jHusy/vx3c5H9Xk66EvK1cR0mdzy0ALw1cvzulnV6hpwqcLUiQxtD3F3ysBO55r10qc0omGQg
FHQJTNAwPSkd9wRNjdlkpwS6lca036JEPkn5xnhDfdwQl/+2/uRvG9usvmZ35wX1fRQPdwIIwXB3
+9YsBkuokMkEnLJUj1mXxoVu86pD+KSnzxtxNmJl+3nGec+vuKsK2a9SoXaYtqyXenhe9DpOfR3P
pEuIJ9xuooErSDb4zSNI02fC2fPj9DF38zH8dYkMaCys0YjZngGByRxeWknIBbhsFiIQafe9Q2X+
QF1D0dIHy3f0MNb9MYTC/7z9VIhvFAsauKDQ1fDooAseWzjyl8yGlkq4/M1056LRrLRmJLXhQRdb
xc++Y0M1L+wE6Az2i79a67WjqkLNQDn9srJeI2RqNXTh2xYSK/Q2WLqRVEahxrJTwQWVUZFWJBx1
a/HFh6/QbEcW8uW2attJdc+au8HUfY2c9nn0X3ytGB+/fVFPyTw3ZbH3N3+ezkFZ2lNrLgHBckHl
s4AIRaknfuqLMxYrrHX/2c9BnKeE8CcMlfAs1V5LERRyEElQtqAatkaKEVjL4IM8wV5c7mVgMNQB
6J+SfinXmCAR3Z17CypP7TLMbjynB5XNl9OX0rhNB4ODJk2J+vAL0hPizM0BpEOWBTQzTJ3YK/WO
Takv+dGEExcwGKAhTAdB/qvM7zWfTrzMRC9IRFTQAS2br5rBm8o54z8IY/uv+mG0zgpmGKYW7zq9
TFLXvEOYQlZGqPZKRfrrtWxiEAUOJPn9y9drMbi7v577Fi9wXDvaINmhJDKMMWBrzLR9q/WRwgRx
mMgeZXh9YOODyUhoZFB6F2jUyE65Xz8reTLqaeyY4ezwyBvXipweE/YodG/F2aVXB56rzYOtGWlS
uOJXZxwRWqHVf1kAxz85H7uIIYiZy/1FXI8RLSQqSN0emrXLkTD2unXlvFODMA5oHMh/15tPVC1/
HEXw7+20HOLhWMjVwFidXF7YeURsF2zspAGZhFGKRzDRS8NHnyO8vQca2FIHAiyZiNXZRBPruRJ9
XuZMqud4g1zENn2nUplvfK9YmeWQvb0uX+GHxAnt/BIVuP69r/uWa64wuMmj5jzS/CleOi7skpbc
Xt9igCJO9rA/NjOclxbFgotYtlO8aRxKR9FA8uqmviwvaJiFidNAcHqXj3zzrQ+DqkHDXlQFmTgA
kMZTxLjjw9v+FdPbX8c6NsnI86ggHPpncMCVj+7Yz8aXrpfBJ0Ai4nN/lq/9ej6iEmF3BtqJfq00
mrAIBR5loKt+M7H4fu4s8iMHIXuiQ621EKh5fOavHQ3VzIlNsu3DFU5tWC7W4ixJyGmkTwzWJsPK
qHMMfknl8BnnI0uGOKgzMt778WX/onRmjy+ZMkF3rzn+jJGwKlPXXg+62IEBf9X7gnxwH+2qriXy
Wn2ow/6dtzZ8+YeWGSnas3E+TVmT0ocDCpqrIo25H3bPMtk2JmH+tx/7XaVdYY5FRxxgWYGWP5um
/0ChAmrNhvUZ4wwdNU6rvz5DNEfBWZK6mPjtyExneCqiF07DcUJJdb6e9b7nCdxSpfuobUkIMV2B
NdbbMm/jDnn0bqvVGdi7xsoF8orrad82uHMbl9oFpAgG+FuN3MXitstkE7DKYJkBSIWvU8uHYa9a
vyfpCVfZ6+OAmKxUyKVdrZjnOMNxqPDlVI9MAPpTOaWZxlCfeY0LsDNtCVhQW5biJk31us+JIvYv
+k/QE+TdHulluPGUVVbwt+u+xiVEpyosASXJV/+LoOxx4Mbl92/0Zt5T61l194HhJ1ot628lyuER
us2i67PqHTxS4V7E+9TjZtBUw6ZgXulons8je7YH3Bo9TeLvWf69KSpNG2ikLv0hWjelIqn8MV15
rS57eGlpEzr6V9/d7UulN0r3uCbdyEtb24YQAa5RwHG+baDf/O3N5uUSLrsc5X8FaPswhqoIZUDG
Ei9l6HeUgA9smcTNXPePUgAdaindl14hC7GvFnS4s4WAabeRmwkC5ATOCrsvNQxrWBwlSY+/MOMQ
q8j6+r3jALKeWOc9CGUaUwSI/6en5dYO7ZAGCDJ7xhN9Ex/nB5bHPPMjUHF7ZU8D3dnOCd4RBoFa
s7TzfAJgz5P3XmY3v9Shmh4+22XQpLqb6G3W+6IrzLywZVuiTKlEXyk5s5hPYH3Q1mIUPuerQHmz
/tEa8NoDJZ/U9Rc0ArUXsUtSpFXpdE7B+/INUMuSnRj6Yn2fb3S1NR4Lz5UeHdGg/KLjt0C/K4tY
9MqHXr5MHZY8NIQIMICBcA3JDftBWF2AdS6WO1wBFjRRABoSpuoepQ57hBNq+07KTBnzIefqboNj
Gz7/SdseVvlCo9KlvLVJuIItg7KkmvFSVAhh0nmiQsEzEISfApkpFEWTtNWxgO7a+w15ba9UhKLV
/38lZaicufVSXHEucqswptTg6My1NypZ3XCWgHcJOzBrMehRE/8dBu5wQ5qg6DOdfwE0hFj3hoRx
I4VOvfM3D8T+iRipLG29XnGhhTgLXWAKN/4inMKOcrpfhOWLorOvjh4ihL9PZITkjpoBhXeFw1/c
1z72dvRLV55waCaV07XaqAfgS7aM6MZdTnQvpMLLX0xCYQebhNmlN285G+jEYS8BK45YkNuUoL5p
aWM/ImroHIrtnjzjjW97CJ69xpPBcigqXacq4YAQTPf6YpiESxyHNCOBVWqyIbb4ys/XT1ZrfOrM
8/qSxfuSDeqowZmG6+LXV/+iUpYEhPyIO9mTWiUqTuX1gJ33cncjEwZ6t5VMg8MF443C/g3NivO9
JiWjIWs7REI36YgzcuyqJfVFuT5MzRlOTbt7dGrDgTRXSkDudNuFq5hT6Un0GA/HMohjYSVNJDbt
RB0onNfLsbEJOTdhbllFPeg/uyOMkZFEDbKbda9V1n32PDr+cNbqJ8wzmglw6IHjEawnaa3nL4C6
uu7x/kQOHBcmEAoGnLB0bUsYljPlcYu96S3hsGfa7OdKcO+YlcjFdNAEE1Inh74IQ+gxuRZMzQZ8
fc5Dc4jtLL0TTz5eW5r4tRRCWlIFqijhFxI/Or/UbpInVQfmdhoTKvDXn/9uH5n2yfLUoNuJ4EP3
SJTZZ0GfiLYGXMSRhuj6/JnL/bXz+NlQF56gTqQ1UQtPZHzxqaNGZvy0yF4INhLgYPVl1g64GkKl
VxMwrBKIcKMdIR97qbXqq3WcqUtb2+DL695vWBiBxhAffX5g6yP413/tiwI7rrqfF7+qalL3cAE0
u3oqBTyPgTR9pWFycc2Vpd9NPaxFe/2pMKJzhg2XnhhcdfCSGc2UBeitjD+jz4gpkop9IjOS2mGe
RtnGUJLb2ELgPstVPPzphM/Et09IAwfFBHauC//DYzbgNujZTEF6i+tg7fof3bA7jB4tPsD5yfuf
Ry6PjBtPl6Tcji3DcsHY4s98xzy+58vO/RodP/GZ+f3zgh9+NgfrCKqcdIAOhq0B4srBfvlT7RAT
WkbCIIgXsjh3Hb0M2Q6ifx2CAJsawJUh4oJ3QRFhzbZcBYbX1gWXELbWvfF31mdMmEnYuOaT6JKO
w3Pp3/hYWjc9y0P8cFRJlbL+O026fKHZQJBDgqGzWvQJhps1Ja9v89YH6LAtx6NjgLHj5Do+wjNx
Fg+eJnzmgFqlU4yK1kn3Cqc4Cjry/mLrnQbmE7cPkjEJEBokcMx9NGSWhLniC9CoNodnoMvcRWvc
TFAL9CLRrDNvolxxmLmaFPcZ4d1KC801j3t7qCXnNsWtWSLQzQ+jNqCTrP56xxeyeb7AH7jjmn4c
bGKINQHb/ccNM6VzGPpLG/9gZZODUkqvVYAQw/3gnzE8Jxb4AXEekLTlbfoSb50GhB6xjO36BYf5
BGpdDB0Tmx/RIWGYtGqe/+fZNV0ch+FKTQYYeZ/HXoCAEGqKcGFhfzgBYrgcWDOThks0bWExW8sR
vPA01d8DWuMc5rffzlKr5n5i1t9caSKTlixb9RSqLCH0psrbdJKFB8kqAfLY34ahVIvUlgEbgN01
DJX1xI5wr6km1+Z5OieXA42pdTzwu5fl5yc4i+RCoUKA7HkDpfBi4w1qMFAGORfYWI/yrDld2jcJ
h5YpvIpWLwnyFLz6rAVrYWIcDmfwP0iCKIzwkfW2Ox2vxi6WiqV6BRRHQbPGgjafgpf8VtlkjLjz
vl2O/LhGPR/o4ZZmaSEV1zWohaF6BoJSij/Pss6kz7yVI1v61EabpFkpkBhnI8SA5Jd6BFy4UXl2
0YNuJhrJHbVUIG4509eXC0uiwIDf+w/xmF0/t88CMTSKpu+mEgXsGv+DU+PZdd6KFeMCh3/c212j
fyD/RvEAH+BHcqf0PQmn6zejVrniP3mOcRMHecrP7cEYP9FMID8VbZjqPV8Y9krmUb8H1miLcMug
DNt/tEGgTp4/LqDa9u4SWL7jWyjRkYzYnvKNPukhE/7fpJSX7G4dSmhVhtH9dXGZ/7ge/CMRv0u1
n/9Zvg86X3TJWFG9ddRfNuOkZfUqvbB0xCO3CBJA5F2sDDh7wVjsIMK5F0V1eLhMitaL1DCGVAQV
RxDFSh9vfFBvfjNp9O8OUqLAoPnAdWO10kIgQhljMCxmmHHC+FU4IK6wnyYtu2dvPivwuiqyx3qQ
Qu9mHJ8WTMzgn0dbayEaLmjGscICYv4uSAGrJLthdSLsNqcoxhnJZpYgvZ9GtqQGaLlWw2USLIZi
uqSN7v4RQ2wjXev/IagVJxPPlJnMZKx8afDfiBdQy9AWCBcxk+6KhwjnDy2ZFrrHrkRI8tx6qCxv
OHJpDNJPp0PkSNm7af12kgvLj0m0oqmzubQFyS4tUmy7HWNws3TNtyYaq5btr1cC6P3R3+i7/+bd
Q80Fpg55+njehp79ozgqFvPrqpntF2hYGO/INib9mhQ1VjmJKif4yXmgakToJWI5VuxzFmxpRF+/
a4YxtKOT+KWnJJaUipAiqkclFlv77ZmJJXOgeYyOVa+hRmQorcbcvf39r4AZccny2jZvDQsn+vMC
WM3++RUGnijV0ClaCA3XBIuCB0QygI8y2v8jc3FfDRrswJ/wq1FLm7+l489sN9mTb5q9ORL/O/ch
zsaSo8Z82su1r00mhlHil16Td9TyvJWVW0VNGgnAzcmaLP1OTRzmaN4CXqeU/Oc9pYBlw1GAZy81
ckJ6YTikSHywiqxwzzqCPu3+kSTz3R3DH/c92xemxsXEse2wdWaJAo6eq1V3bmUoKQ447U65/v47
9LEtpQcBLdCSk6C7wdWsHQ/Rneer0zgWjYsGP5OKUybOcnZNxKQ53yF/NincSgkPgPGTJucPpNlY
tzYcVa9ziONfEyuNhVqplBdzNaBEDOUAcy6upPX6n8Gm3RyWTF0DUKj5Adt5
`protect end_protected

