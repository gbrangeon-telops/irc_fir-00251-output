

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CJc8rmbxQK7PiD9FE9h/V8z28Q2yjtwOLUGOHj92X0D4bGhAiTKxH6Gs6WbTk3x8dF6WKWHXW0Xd
imaqryWs/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KUGgnJN/sGLwh1pfD6BBRkJkdz3qYXsMmFAG0D8TIT3kvn1DM/WYFdJfNjuI3TZJ+GjJhgQt/TQj
vszszvccproNtKL+iK2kDAI+dODbmK/3dk8pZpjNIY8iqG+SZd4LOHkCbGnDn8J5L1SCb1FbgOpc
lYLzGKyKMfpMp2H5zrU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QPilQnlZ7SkqHJ+uQKxasOWlKPf9SmSQp0r8PPqOPGeQK2aUl+9gzicjiy17/DdQAM7rwf++nyUV
Yi5HrcGStcw9bK+k96zmiNT/NPvXPX5xeKvpNagObga/il62MarkWpibvt8B7D5IQi80Rp8/xMyy
QM6+TtOf7NVahw7dZAUwr3krfROulZTDfEY3oalO/PlnwAGr4Z3udXzac9NTOUWxkjpW4cmTbWcJ
unHhHJbyMO341XtwkTUgKReezgKFOpi+gREeBT80YOKcPQyjGyGuc28HYVmxKisVh5P7BYL5neLX
P5GVK+HA7MCB8DsbsorDqal6rxwDeaIF/kJcyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZE3LPHWjt8FXIcLXD6pONgldgtzqHVcVbUx4Qj9ztf/3D9DwoYFB/m8dT7Cv2OabvKVMu13QC5lB
rxR5Jhd+fouVouDNKYwIESeS4DEkgnwfSJpsmeVaPW2tqCd21tzGTVfcw3Igam9PcTjnI1q1568h
X1Tcmu9paLkGRwvQeII=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EV5YorhH0risCTPPpyQGO+wsA9egdTVjrRAwQuEDG89jVsb2NsTih5Y+XoLrashGMO3AtQzajDhF
KB2YGM3JfNSzKu3jU5R247s9Goe6ZA8J4KFFzdwq4blriCHlPX0eNqXwJaOF7SeF++njAnDs0TkW
tSOb3VJRRI43LgFv/CHX80X62oIhRm2LIRAjPrPj7KevSjFw7diU9sSURAffWyrhgq3XZsUY6ovy
nAWzeDeWY3xrRDkxjxQAN8xOlyfUxlNsf7am6Prp3DCG9ANkw/MCyfCVBJXBbghP4T6GS/pNjySW
+j4cMtiThQqIcJCHVcAXQA0FAf6PbH456gYJfg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
O0BrY+7M4teatHcv3e8b4gVawTcLjA/NrejmxNsSTzQFxiz8ecDGm5aaFkVaGJBP3UjCAe7ufACW
xMxK94MTWYmigoRWgdXvcbzio693tDZgmONPSa86ihBZWp75VvUCkRm/IKWtTOvXe4T2osoMJajC
oMKDmkzaw4QPM+QTdldWMbCtfIE1PRGKOtrUslxpUtaG+0pohifCSgDpnPyrweVKTDtp7LipjX2L
mmQrX4ByJfOhC1h1yv9iQWBDRvA1izNGy9XyY9UQy0kiGZvbsMWdjz72HVz1xaELKQc2t8qyp7cw
4kvH/tnUoT/yoIkdE1nJ1Zjh9tpmdvvMoalVIPFitGIRT14hFwm+oSUI5GNhUMZq0/k3/TQ++jI9
nsopQbLdzi0iLnBxpHYz38hlrcqmBS2gygmxYLS3fCLF8rm2uRNwwS6QUh/sa8MJqa/ROG3q9nS2
c5hU5haLc0n4anwsPoOz6MTeCnv6zZQR7CmcYqsPZcLfmlIBYZq7RvBfgxGSSG49VREP2PTlvM+e
0chz98Z2JComfIBd1brC2wzbulj7uaU7ZR0a63B1tvrE6h60wHBP7QmZtAJBal7zz7con2J+HVrJ
qvc71JRddikpSaAz5Nrs6K8RJIlhHBTs8mvN9f6ebElEeb/uxsYufl4CUhiQpOOea+sFC3h34Ptx
8QWOOr+g77fZwiSprBHCTncPDc39uvz2KXFBhKfq6ImDGphqTec3u7oEmbLQMERFJO8QMcxdVr0k
uhdiu1kRXzhyCLDPN4fmj7FTlyJ8gEMxFtk7lT4m0VBQl0JG5Nua/24edFzbtvqQ9OclRag1Iink
cG0EQxQFyQNkrt3z2NsXujWQIWUqDSqjcZqdfi3yXv1YlzlIrofXWGW3xhKBw6VgVeACyrl2rDQC
mDTYHRm7O8f4ibm/VMBXjyz0/lU2MMiky+eFR8SdK2uaWfCh7Uc09twcLDc2EWeJukMiy46KM1t5
QdLn7FFmwZjFapnQUn5gVDUUvWIOe76fiPY+vfH/3jXT+28NQaiTDZISlpqbau315QqYhAY+ze3O
+wK0pIT4F5fRne1phZ9exRx+S+Qe1GEOCnJy34s9aZm/P5jvGHXxQoz2/qEdocf8bcMEeFAv+2RP
HFTRM9K9CzRdev37w7PpyVbWe4hvnlVaRAlPUIcxMebOYHSthKn/vsPVDD035Im5Ot0PizIThKR0
AzR0sgC/XmDeYBUwF+N5YWuqW72XX+AVVMOHM/YMBeg6/Gs91qWtj0JfkOSYaMwQGZLRNt99S1ZE
8ddOG68kKn1Inao5yxPa0u50U9+o/W6fV6lRoXC7WaxbfP3/lQstJxGTCCXXHrh1WcJTDyM2nk9z
nS5TDsYRhfEA3tXjntfCdqPxTTMD1gjYVza362SZE7ZPbtmW6Mxo3ss+ctKKvxJt/68BctRbxGlt
AiuxoABgpvrPdj0Jp2Ns52gRU681K5by7pN27B5I8TFwZsB2GSjwG8Hj1XvOgoIhQDmTVX33Aa99
u51SjPvO8qNjlqhgZI1iZHSoNDsn7fA/ApBBxzzonYXYP+PoBkLtPBIOmwoTw5l4G+Q8yVb4rDBG
Yci3/VCoHDd/htj5uowvVBBqwRIrFveTp5iVa0oZiLARuEeMEqwHDUuOK53g8QfawErWG6VtGUN8
uqAGDk4nRcpuWa7faD7jzs84NeeVpz2/BS0Vlj5xKKfWF+t02+qTSD/3nnQoXVo24rfbPb5rljgB
JgfQiNTFJ7dkFTMF0WK9Vz3vLmnnNEABrDKIvYh65pIVowHK/Huu3cNAUBYWH4MWt5C59Uh44ecF
8IcgVbqGVXS5mLdChsfX0tunEtbMeXGc8v64wVgAUXsK0GcBxNyUZ/ZkZGpQPjX1kN8OI6KmwMdg
d0vNLVZfYgMZHI5QGUlrrOoIKLXYgoObgxqOkk6zZv0wSLNk9rAV9Jx/REENmfBcXob3pDJnGpUS
wFyCm75Apgj5+hGwpu1k0mdxR9KaMRIYDVqkjHRsjiK710kup0oLTRUa4rjHjxrERMQh18ucsAnn
kvXGfYfcg1Mq/3p2sCo3riBh7KTS48DjdSCFVCVFQpejH89caYDDFopsNDjx2XxE9cgH81CbCNvj
AAml+s6Sl3n6xYr5Y2XLcNK7zjJ5HXnuZrsF43uVqrsdhM1DdU6APkr6JIIL6LyASbRmYYB8fvfX
9tJduHkB8vXgagAaMoo/vCHC3ZmDVwknh4W6NP2kfT78jjQhU0CUOhALjkET4MR2roPtZ9ZFvSjj
rbmVsKXZJ3ELzR8uxrWZxj5bTI3fRGNOtw1FjtJ3uvVL+oFTLjTl8N/jgfaZSemSVWqQfTcEdGKx
m2VqxU5Lv0sRijtOVS7NDH3IhiCZwRp1QPLLxwrqN2MBEmVHs9+SX1fLC1SOk0sROgGCo8SkuZ3F
RvIfT+cbpVjsMFDZCQjmtES/eBYJBThtdx9+eHZXzcn+2pZ4bOsQ1xSZxzg4cSF90OmRvRqRa1lp
/UQrkYEXGYonS9b+H3QYeyee2ndih/B3xlPSJYtEcvdo3xHzDaJYzCHNklJA/vlfQLJqRJZwNsLX
iKyWgHOEpF8AagCeVhJmLZGj0aRO9U5sqEtSoXWsALsOFFRY8Fq3n3fHIZgSgtNTkOOh9HxRsty+
GHrKp2xYhADBmKuoYzNC8175ffwR/yPRISTd10eonvBlZ1x+fd7vRQlwOnSNEHjGKSugwL+QTdqE
yKNQSaq2X9qbt7AKrRFGm0jOJslzxfmgBLhDY9VMfmD/LdYMVfonapTE1IafJLHGeLpQENQPu9Nn
wkAWDUfXb0IuMuZY1xb5UUV0C9xg528vTAiBVgjKF6SCMNdGKrLSstieKGEofMHId2iDv4YAUt2S
VY3fx/AyMQJORaD4OnglKT/1BFxDhsCY7GTQVVCDKDBLm2n/TWYJFXH1kRNeD2Rf8HFBkq0NM//Q
Mwhk/viezkqa+v64ExwnXwiIN6XwDYWfKblejxWXjuXXSvesSjH20qSSQaec1eroOS+y8vwahwW3
B6cJAsML78kPxDNlWoOHWfg1jeITjD7iT979JkQhZpXLo06IuOYY2fjArjWOOjFc4vlV5V7cyIY3
D8mLpi6GHyPOxnY4sXRwsfbFOO9uX+9WK/IWVq1QpwWu9nkG3hXD0QQcqjCmPtbI10uM06vDyecw
zpkKcRMNVPt51rzKTQSZj7IN9DYCXY3NQPXg/AFHxPK0Ia/J+SqYPavvzSWkRvcTv/iOFK0UEZYl
xumdpRlur9sASTZRwDUe3JppDHguDOyn6P6NJIubMScW9o1zcaMWw5JOCbADhtcB/wHP2semnNPn
S9aGl/yhOFeepoX/zfbaMJqkwO9hYmwBJacaRWR4dL1z93k+u7/DQ8JzZgGqjhipHNPI6WC3yzfX
TZd/dVDoQ58YP6gviiX7HI77GVurQ5vzXCE+IBqf33pTuCbUGkaECxb/l4mr0K3LvxQ9KeAP0XJe
iGDziOTCDpO/xrtjQhrdDPjT0n+YLit1XYVpToF777IohQWUaWSY9wDhMAG+w8yUF9w3rapiSrs/
WL+csem7PqzyOwutfTMy6KmOnJHoUv9SqThMMqW5XaH+4yxmYnP9gkshBrfgVecCyXYDovkdnouC
pL4iXY+7e4HEqyFG+6IkMxzjC3c34u2LjBnLNsVJtp493iwB7Ff6jbIoHmMAWnC7VFehc9r/nAVI
sWE4vmvIm5kBrKX88F2DuJEnQ3Omw4nWiyEapbYAAIdK2gNEM/seDZCCk5lPlu3cKYqUEfj8mrIc
TZnpXARXnm0UaWgIa5+4blXfFT/8isaAjTtCbhEdoPfnkLt8Y4HAFyTiDJ8PM4YdLMQNfYk/J4Gq
dQVcGfV95b664wvBoWw5eL6Sa0Ec/TzoYlxkDpzxO5hNrsuNPgUCtOsmvyQaH18lz/frKURm3YFX
1YE4mqpUnL61Xa7LtOA+w/2cFfEsMAt76LVgwzEcKZNLGTbg5P39o6v43yaYuBOQSERBO+wcAvh3
iEhtlktOHBIzfMshKZK3/dfBuoEiTMJuL5FiUzJs3HaevDnmUAa+51iZEqTzc7elqoMsUR37k4ze
YCg8qDp8a9lg+NxvTnrzsJ0jwlORgl02haHoYRoKuSO9WcIYWIL8RceAIvBfqfN5Vk4zeh+JIlsP
gFx7uR7oMt6ql9/+10kv1BeqzSHUZHchPMIz1cq5IUXxkW0CfKdobx96YURy51vaVHCEjIqCZI8l
srhD4d0Z+reBgRq0FT7qfWIdy5EMdQgOzwkb2PN9bgmwBj/GJ0FXZnJ4Da9NhitQUwCMDU4w8wjp
xkZH74lDwCW/IFf/M2ERWsgJnyJkVv48OuTxedXsFBmHJ4PhePFmMA6HUgtqd4TxHtBT6qYyRSep
mhZ+JOzutQP8eD0BvjLiQzCzvVXjfa5yBOllEj/0/LBUV7HOnJ0EzAUuXsF/Aerw0VcNhpMmFS+e
aOPByHHnFUj5bhPeAp5bHc4U1Js5YQm5RKHPMKJOZ0ucZrCDE+xBSLAOsNgyDcyEMhGz8ZiqmvsR
S+X6xgqYmFxsqPMeaviNxvhIpdFsDphIwycfe1r7JOoH/FJhzoWKK+GNi7afYDxy1zw0LnvLz9uA
ZpHZIsNe7SSJ0YuMlXdypEBV0EZY4jXQXJcXTow7+puT20i87JXJc65og4IKF+2eIQljDBrUd7kU
wGezJeSHpmlFAZDaIpdiVzt28QO2VqojoH7SViPHWmLp+JWL43VC4n+hVMzXNFymLBhimxUYh01I
AiCzOmWGSDA7gWVu0WNy4cqqRDbu9A8qeYNgeQ/vvKtgYaMBlgobQ2fSmlRBchq8LcqKi+xX2Dxb
CW1bjrXx77ZLx+4/WDxCNlBYz5D4mHol9CbLL52cOdPN69hE7PA/6RNWeOo9C/nQe8AKz+K+Jmdd
93AX6DX88d+3WDNWN/pnA8F1a4HcnhBRufxGSXypJh62DGQehtcys3a/LPYgmz46681mZdwfaPb/
E0w/qGRMea7o6L1RlIVkszZqaQhDEPiEpPZ7WpgD7kEMKibGVq37CTewboSL+925EEXfSDELgNr3
7ewB139ediuiGl7qnZ9yV7nwKfumv41JAzAdujszbqsifltEeOZitg2XphLiBBVzu7XH9MBJ/FWN
qZvr5VMlHzoaGQ6OqcISGQvbMRGdrEhdlxkgI85TEFj/dC4qaV1NJpxuTct/V335AS/rD/oqFAIK
fiXln6MsxT0+UEhM5+1Gxhno5jwZWcaskvoR1IPi2telqne3Dfn7S4x5vRu5sQi4ReNR89HKEGF9
VIaCFMXAPrFZVGbBUEDjg1QyKaMTBdS5tkdujwolCrKb0rlctbXOWA7GB9N4b+sCtGD8yFNX7Ewh
9wxcAPEymABkz+Y/hMjFqGanq/3boi1YDK2AAjH7kRwkHbn/Naghz3V/zIzSYAesIzfHovQm+2jt
/iF6IW9AM4dKgCav9U1+QtQkCaW7DDgFm30aKKk0qNCBlPrgOXa+TLu1wGfxjmKGF3Ezpfcg9kaW
46FwxumspWTJ2lcv8qC6kSVnVvHIDjQEAlt15VJarxa+XENoWtYAmp6AEu8t35OPbY2wLQ1ogN77
Sfe/toSjG7CEOxXaHGnErTEtJKHXoNgxdjL8mA4PLz9G5GGEBFDGmlz5MhHenGoWjpYpkH2wL0s5
eFjVNPE4V9yu+beeMI4IkpPALvhADNpdi1eUVGgr25C9g7TgsvEOGs9H0D0XeMXxkr5VKPvypYDs
D8kO/mJ/+D31sF1DXGlu+UgpFuC78SS6z6pZnMhe1uviEPIL6ttnwmsH8sSU6CYk4u+K++uqwjxr
k7CnRLvK7bZq+CQoMijLZon2bG1Cbp8lJPTi3WzCgx52Tz2hy0oZqLv+d2NbpTYD5lVTVCqlJuP8
1uXlHKKYfVXpY5JReg43PgzKXMuVXZgwLs1jOpLdrWvuILq2ZzZa/XB7H4oLrhol3RbArcr+urLU
qoWqbUD573eOpyEb2cnzFgnglOzzw6+tJu/tg59uL+7KD+CD1mJXmoWu2PjGENesucuaC8bbTin5
Lvtydi/SMIPHiG5RpPp+JKe8d/2n2f5rJfyFwK+yVmyLo/AXlAT1x1sLxdeRMxjCklRUOgZLGV8C
Mtxv4dsIeA==
`protect end_protected

