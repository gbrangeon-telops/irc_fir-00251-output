

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AEDf93kkZknTAYDLPy4q67UmP9O18ta3jK/RtCkxR3ZqpY2KlRt7rza1H96MUf+qsK6643W9A0n0
TP4few4v7A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
erRjv8zI0elbdGyufePGLqKRctW7EMRy4ag4V3lsqysjcz2IbkoY32VNXZB9TkYq6LxuID3xgPR/
/dbN8HKNlVJr4fTV1LqzlQYnx177n3iaEwIdtrjwP76G8DtyrbDzV/JISwzd650MMmyKJtHnC2yw
alWuAIIBdbSW+HbA0I4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gdHY5LRWuJLwhBPcRYPMx1NPD/GuGCtHF8ywmbYLyoAM0rjTxb8zBoSHfJbS/2vKpgG8RCdZOknj
FMJ+fOkJbpOMFaFsosZ9XfIryZEhroI0pt0zugw4Ha2XsmQGqxGDd3IyGRBNvDMKRw2cnjSZz2Oy
H3SrajtWuLhpP/vuSzlhtnqryvgbp0USaL81fja6LLlPm2jXTcuqgEPsJwwUUhxjUSQyRtABTEvs
3Vjc63pIVZUYkpkoaKpA4243dOoRhazlhTF1c2Dp3uyCrdGZU4fWhJHW7m3Cq9Aw1murzYGrPLS4
eQrf4MTXbiMtIPpNK49OUBbEpUuLfnDwfATFaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fCQs5S/zt//IgxsFc+FuMl79LHVh3Px9B+S0yADLC6MfIDCRddIdSKbTMZ5DlFrngWDJwpd1JzqP
cRXcul8iGoVMrVmrEStKWXi/mhtK5UkWTAd7hoyj5zcI+N7wWWxU1eBAeKZQ7uML2SLN8mYzQYLY
98ufqGLyMQeFAWp64iY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rLzkYB2xv7C/3jKaA9rJ0Hz1NLTW5YORm+QksBhLo7WkyUXUd0Olk6yTtcSIC82lRfBo8f3njqY3
dhmWfikGbTNV7gixnGfPYVUvZg+xsJ7adfqwnApC/cK5eBJGeWXZ3Z5gEbLOhuRw/04o37fRIoCo
Rt8ZH/C+LE5As0rIpYw6uzjL55RYR91wP1R/rUwMQTNJ8XwXPkAbkuyw7FWG3uW7vEvZ/CGu+T1f
VDCUznG/Mry2818W/OOR+t5yQ5fYiXNh34gzkO30FRWgtIR7ZfOn/fgLqv2Iaq5XPzTdULGOHjv5
Pl+0fdEaYyo+sJ1yt8Il53T+ZdgLTjEgv9cjPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30320)
`protect data_block
YBPQ7Jw3lhLpDre5nQ0PZ+YiLtseFYN6VbGYKAGo/w4uPcFwMs0RfjTDrb07PhddnZ3vzEsrZhyp
E1gV5QBrqYXhAakqkpDODonXVHfR4W5p4oB2fmcHt96FfeXsNi9d6DzeigTKWp/NJB+7CYFRUq4Z
6PWlB3JC+qhpyKoR0DCH29L5KEq1oUb6C5uVeJBOu+SBzMhsaeyQ5RtuvS3ZVZvnMO0+7wra1fKy
h/cs6R2HR23ZnxBXd2GZJuY3z40lLAiFdKQ0OlsLTP3mPs4Cpe0gvm8CD/KNgBxfvR2zbb3ltEe1
c9CBjjVqui554bJNt1DsA2S5KINb8+HERNHgi+QPnhGnfzHgg1nyIN80PSDqp6HNEonHsBHGemmW
K+OJvaAAIsEPQZ/l6X7ljYRoNDtk3d00Erm6GGCZcdokVc48/qj2yO90ZveyvF+xbBeM96GLMQsv
nsornilsKdmUIM08EBjTbDNtgPcEspr4G75u/rRLqYc2FKKp3MC0KT3eW4tmG6ZfWbr+P3UCCRMV
ZthLzO6zX/ATviFE1ofrtWgig/r9iuSWmyhf1XwGqfPN7Jz10rrpIi1SEL4v9QSKwWDbhHdO421E
AdawC5QRuZJaOuaXREQjlOJByyye+UR9bzlKp0MSPThHEXiFtndp+RGgDgZHg/nYBbf6EIdopN2f
ULlFRJBMXJepucN09E2zL6IanLFACttkQm8jSCZG3nWbLNRW3EI9XPqHwGRIMmR/uD6BnoIMnP37
6raXC/apUOFqDsrpeJZ9vL1tfNZc1o0w39sGXKJRSUv8pCBMJiMmOAUAzrf5h80jPMgj6Xfoj7ez
FJdpRLyDPJAc3k06WDYIOirfWR2g09pW+K2hNY41D/kbU6PyyhomtYwKggHZMiB4rNYExG6Bl4Zr
LYnW2EahtWr6wnYRQZOi/8XGqhc/OTa2y7MK+4vpR5TIdMbmwuZWPVoxP/mT2/XlukMmFY6iEtZS
rs4/s2AKt0+D67VmVB2lQmg8/Ij/1u9pBqGC+m2+6778ZIerexC2VijnFj4lYMUftXzrEKmkMss5
i1NSQRoR9KnYpjj46nkNdMAHhVkx9vnBvGfnGB0Ywfa6hzTa6HpGiECxQG3nfU52dEQSLJsxBCxB
U4Yhnwab54Bmf9aJ7yxS7DuzSBc++GqhQ/2jW9AOi1XHzFH+1KRupLT9P/DYgLj2Vwbpqlto0GNd
4SbYo6lJQz/wG/JFLLeRQu+kld3u0VDCT1CnH3V7W6Llk11myCLXkpBJy9XgyGP0IkPkRqyu0F7f
mF3jUs8BetpvGxXxEgu+aT9+FBmw7jRqgGO1zGHNyZCtLQ9dNC7zEzPMwkySZdNy80Rynq1snkBA
LfTFb494iRU2OcmNesgGsEkiaA0s1LyAUkTqxSwvsMhsTkFaQ6G+68EnUXQog8QN2vSGhoAYLj+E
5nRfHn1SvqlJP8UdzXXKziYaWGYNqzvyk512KV2Z3xcr2tBaQmybLuMh7P+C7Cdc+7M8VZAc10QA
YXiJU/dmVXKoGkGmDm+jm51ahMRSTLA03v3TqbKRNFaD/1nKk/NJA4ovqYpqfM+YLex+Caw7PSPL
eQOHPTHFR68C9dkWuKQVUpbPjN2y3tmhEd0yPUd6TSRjmwpjb9UqBhhXewkJAyJNCTmGixV9P/2U
gbfbMGi3B9q3GKxrTxGKDcOY5uftAuteQx/5JFfMFhs55daIQHEfJ7agD1Gv9slDXR90ehM/KtIb
1glBB1aIsDH3XanYSlZdJUfJibauVitlq1a/JVG89zVOxiLkpSuWQ1whz++dqMfDGnZRkATKCcGN
ItdWRHkIN28tWfDXUSsJinuBT9f/uQkctO/XDvaHfVispoznPqmaC0W3LhU5nlCfMSGkm0iwbNIq
ihQss0QfK3Uh/BoM7KGCmd5gNsqlZ64eCxXJWfFr5X5/co52MT8vav7oxL1iZG4gt4tjIpztfvwE
1GJALxdS7Hp7GaQGBLyd1I0p9Y2QfLlMYGkK8dU2NPprOycwRwjPlzQZN2mGtbgXysWnrIje2fAs
TV6/RZG31hUkSrntNY05IctOs8qemSgAt9JhP4sE6pv+9gkXisjIiMYdYZMrIYbdANmwq23tUoVa
NKj877egi0Y/zamW8BouVqMcHw4U7jJQmcj6iODinebROMXfBF2Jg6AcQzIkRXUJ+MS2X1y7+h2a
Qa9Qt3Pahli/BEwmkM1rawMHk76x+0fpqIBiNWFbn5ENn3XbvO1jZj/nQlSlHwhunN3dte/kJ8wM
1fp0i9QXoQ2MjAASr58fcOoz94aEbVwUpxgxdzOZFWoXAmuh5dKsg9QMTgbzcHe8iwi6tdWCU7gQ
OiZr2fze7+Ijxxrhp969meaI0o5dYeYBGUlq0xGdAMveN2dJ91oABUkgSjdGsI24x9JJpWMmH8fJ
GkCAcb1fli2OmFNwQjSfJyiF0sWuoOnlW6lkgq5eABlaxMa+ZlY+MPatm6Jvd+XHfjGBY9af6Tn9
TctOgPyeZ+mXAZpkuXm4v2HZGtPRJ+h9PzDhI0OBWXFpWKU0X3XGsW2ep4sNb69CBqxLbbDFOj+a
1kpkVSnlz9j77tdQIvlQSf4CmZoZjn5Yd6gh+HKH1eN0Z/bDVsO2MMPdY+BNjzIEXsvlNE8LT+70
d8YYLtgkFkvOqoXdFLhN8x0b1jdsxYWOQZhla2ue80jXUBjPJ10b1E4DKhDf4KYzc/76Qw9QboCa
aQWQX6fqUGUJ7Cdab4vHxd0H/TOiIWNqJM/FCPPA3PQntV87bcVVDjj0Advc+M+WOrQq/8KidIGH
hNNJhPn3gqAzhFdooby5rRCPTj2KV4lcpHkfRooDYryLIfD4nO5U4c3HzO6HiulfLg5m8bJM2/le
18WRct0ZfHiOsDUDq/6TA5BvlefUabaZXUFlMyzikHpPymhWl7vL8vrRs4Uiq4hbX/Puf4fVRPN9
0Y3kJTGdyJ4DqGCBhhLfSZnPC3mjv5X8NH9HVHQvai6S7slXMza4J0Cyu0KEl8bYeJvacY99H4Af
6gvbDjsUVyZy+v/PiUxCaWWusGBDvvPsYrwfUclV/bPKXzZA+ceq54Aesaa5iDJVS6WTx8WU4meF
4p+Mb90z2yojQ9iMYYck17fJ5hfytLNyDcYThmiyyHJ/fM1X8xrKL4M8RpAKgJotrLa+Y5BR7jCF
v17dtU23INQqu7kE9BxM1hyhJ28ArWw8NTjn9UpoCFkOFQALPN2gWc2v/O6zQttf79Gk5p/rC7YW
jR8gkRUSVc/FVQcGCtrJ/0ExzOTolAz/MwPzDxK2YkLQZcqxwrRT1Wh/YF4ivve9HwS/Lito5JuC
C+HMRIQu/KGRRUHMWzCx5wkD1E4Wf2Om5uMeTmMpDg6YgY0uftjYQ7u+GyjlQ52nsiT3Bety+Arr
9RX52SGfaGUPfPx7VLVwZwK4bVGGgLLY2yEWTJHWcaQFBeswlwjcqn7iFWwWkKtQyqEkLPwpYo0r
4rDO5/+2zyQP+O7uHkJYh8CElAAKGm4sCCIti6d80nzeTrgRUb2QFLwpUdFBA3KG+slVLEYETcLx
pTsT3UJIws2scQTXeHqbANtSkK2CYo+5iKgW5muYsxvdw6f98rRhvR1hjg/0uWxg/A4GClpMa3YU
6AoQsQnJs2X/GxdJjAOauV+BABfkb59H0x2AOZDLVW2OycvhKldHBrl/nxlZanXkecRJhhongzle
ZHvg6NoYnQ6A2X5uxyrGNtZ9A11Z0XHrjCxR/3EBrqNo8XIT5BVfLYUxcnMX681J/oJXIs16S3My
5kIeodekdFU5bZoFNM1OSzCIPdul1X5ELc1+ar73u9AC9SzKGHBQPuyWtENruD7ypQqKOL8paF1N
SjG1S2CFdH9MiRPmi6WNiUga9InPqB5uLC9OfpONKpRzCOovfL7FC3h5efCn6i3WRxwnpx9i0Adk
HlcgXXa5CjObLjV8atNbVeyVKVDpHRbHdNDNtHpe31riCfNyG2iOR7QVdgXpS3tm5iMKr30C8IbR
wBSL/GbBhAYO7EQNUbP+t7gsm0dUXY/J8JMzdshCo4hJ/YAckfxfyBn3T0kSJY8eMWJU3c4U2jqY
hz+LgEXqYePF/8tj/2uzZRmUVblAzgQxpIORQBVV+Qmv1O0EnzB9nnzI7uWtiPbrkpeAjYHMWdu/
zVVcvm2ofCa9h5SsRJ7J0PRhFBPRtQ16VogTNz9wMceLwjTt5pUsezrShm9PiqLUmXukoOoL/1wa
hZIFNC9W0bkcPBhiCg8+XrFSHclfIrzi5gyrySygL/tqx+3tnz6JoJsAZeNynJu6z8gu62TZu7Of
Z5Rlo6hwnb0BlpBJXxqcFGhjEhzW7+WH7yXKfG90Nzf4WBTuSQincYbfKNjzsgvGdkkp0nYCGW2y
pxnkBAaIO0Ou6e62MC5Bf0fffYw8Zm/TEv+S2wPbsxIsp1ZzpD/Y5uFgDkA4oG2jrmp/PogWQPpH
YxKdlHx3F6A+vqrYCtOzHMDYlZ4KKpHjJLkeaOFAXC8+VF+8eD0Fq1RXl62IggCH2h0ltJ9EeiKc
Xn4UChIVhk+f352o7nboeGRBut4UF5dPP7g/ecmnsiGFRCtdHvHFjxSZM4o8jRhdfsnUqz7fG/vh
CPUeA9evRLG9RRlpDlu3JEJ8TjCp65s92+sCrEJ3h98jFLt80cHFU/HOdNdj50px2aCVMpFyfYM4
39UOVIEze2LlavZCao++Xfw2RPyUqPYYtSlogyhwzf4pSUnsMwrP8eiG4/Aynb0F9OYMqLQMUAZG
KPL5FS9qREXixX/bfEErbU0JSbhHEoKyRIA2FLKkexH/rjCzisnZscx0nmf8NpCK+3VaxlROXAYf
StfWov30MroYnj8gzoHhX5n60hJ5La9Ay4PFiScsMAclKvGivbSOk3PaKQsdbhmvrP5pwYy3M2kj
/7Qn3n245CaTRSzHRxlR4uIIHwjhFfmyxdcrvze6bDBwmlEYaa1JtvZMq00i0ObCiJKduJ3xFdW2
uBbaKxX64bYgi0CbF3CswZrBnTfFSTQIbiyQINEklHm48MFsXW/s8ir6hcVl9dJSy7ocuqguR5dc
LZyyq++9CvGNe5FIqvuqCJ0ADGNuHu9nG1sLwHusO7I2ixhudrdFnIDGIwdnsRoeCs5UeOuH2QJE
u5Q2EwRlqMkbBJ63xdnITdD5JPXXyoq7fdSh7zzAcheLmWNAPwdaL6NydhgkyHiHzUhasB0F8xWa
2zQyMpuXdPuGq6qiP3g7tKGIoahyO1PToMYOpYmjzBYiLrjCWS7Eb1JjbM49yzkDlIVYoF/W/QDX
UFnL0R3WY4nKX+48slMwfPWHupel3W5GACCbtriMYfkxoEsw5NbNT2edB6uv7lJ1OOX0qQ78xyoS
1ReW7lcwRmL8bOWrr0pT5p1KP2LZYLHRspXvs+6DjBVf9PZNJ3K2dpHi0BhsiAbfDY94P7PIpZyE
5yrkzV4JKFpOVDrmjVAnmFzmWmI+wXEPWEjTI+9iedQwVj65NOaYx3aNKZ3sQpG35W926ZQciSlQ
vwo5jnr+75z3qh03MzRHsKFILCioAVr3nHyBFX2x5zpXkZN7Lw44wr5vNNH6g/6Ir54winEX2lOU
uStFBl0vmWjooiNWCOAMzN/UeDIphneciKfL14Ps0ULcXsJqmJdmh6dT/n3444jdRD1jxgVb6GbU
uLxP3jFJdExw5q0GIpBsxb+tpLImZH3hCUHa7aqtg2gcNVqvDMvv5kTWskNsJ3UJOS2jKrp6Iup+
Yngwavyw24jDmmT4O377yOy7POqywTKE5xtquhHALwDhQ97PZS1eplpCV6o2pUoLpw1yLSi6sTtX
KaXY7ea+2SS0BGSofjswMefeQQr8DR72PD3buc6/XzcXFErmiyhs5JbgPsa39k2kEo2XLI1RsLE3
Imdcpv/7wizN7Vo3+lFDwpbOK5fqMhugxIALr+2Lij1yVwbwNZuIzk0sel47IdM9lhKH1u09igXR
JKhjwOPUwUvR3Z9+RK8LKVR1RhE+oFE55pn2M//EFILS3QmaRt2dm27+/wm1Py77pUtzy3kRAGrr
kTZwAEMfyhjjGPXr75VtkiRzQUSXswbZzrYAP0N3+FNRZlnSNeW2k4isCahVZIKx5zdIyXPrS7h6
jsiehkRQoOBjG+BeXzLL2nXF+ACbno5z0nh/enJNaXBoCkayl9fhonhC8nHirlQqfAZWP23TMV5+
VLydXWsoljk3Hh+o+X9o29ZIxXW/oJcgv0wBe94IdVjVhiNiaKoC0ARFtXYAJHsB4TpYkU/GqBb/
Mc8XM/B1HjdlJkQ6yvXVVqCwv6rnYoyUjnSV0kWSXnl3JquJJnMBiAvFSTb4urJ9eKIu7Wik5wbC
2e8l4/vOpPUa5VDq080CL3/qXqdBF5mdsCUMMAz+nka3nN9APLpN6fxiWS+JaRFQewhxdSEIgP4I
Zc2F12kbJnEahjpjd5hRkhPktPSju5AOBmRNABSCvLBsCRRvyye95yQyCV2yzT185Byn7uJsaiVo
iSH/7xWe1adwaf7ZHsKU8I+Tk5E57IIw4tZz7oaXkH7ZBEmIweZoOEqLBqXw+r0QBOEhMYS1u3lA
GARA1/axzXh7/YShA79ZeJ2oGGXrkOi9fKpvFuTMSlhezyMujsYljc0kGRQi6/rDsLhKJ+WkJmOA
/fonOx8pvbRj/TJMG+qEq/dHsRdDz7VGmLXawQN35qcvzzbUIws54JFmFBKpYtzAQWJGVIkOm0dm
D//Iaq7TlfpZyyN5uHCO1Ic5dN1eCFugKE3e2Scs6aweuk+InaS8SJmRSIqRyvtO3Erc9lE1iAYc
k5kTdbsJwrjcPBpWvV6JOV4CGpX7CktY/JLMwJ4PsOGOQ7obfSGNIJiJTSSdkSNMkYwpgNjLIW22
cUMEX8XN6v5eFfaHxGyC28i32fYMmfqY4h0B9a/IH5INN2pLUVdrw3eK9l3iFNbFvrIomEKs2Oma
kH6JDk5z+M21aL5MCXsrkpFr1GJRRvgsP1NYsJkvFL7uQhi9H87+Zhfs+W4EmEYS5F7HE/SqyzS3
rQwjB/G1PmTYyGW0rzxvu7fvwvH8ImHA5Va7hHUNZrg+g31lBbYryHm0XWKv3w6YLaNAF208EAfX
/sz2Bs8xQmhJOroTn4dOdJpJlXYvE9ofRwZWBwsIZKDRafXie5PywyOoSK0SrKIDacxlcILa6cLf
+t7dqKDtIYqr7TK95DpCFEoyKyzDy50s3CoLRy1pi8aukZg43oEXoOGs9fUpi/sD+LNM/QrriKb1
0Y5SpArq3KP3Crub9IiNDPBd2sCYAJkgHQOcXr4oXxrpcOkq2MuGhSQNlcnBSGDC6j42XyTJy4Bz
CcAFIBHUUgVFmZm1pnwjPwj/NC6Z32tJyWY1Ivb+6Nz84Oc1fRlzWlXI6n8gxQ4kB4U8nu7kG56K
W8vK6SXKiYhpl5epN9j25zObZhUSnMLK5z5b+C5pYZzpETkC3nhRANXFlO/EU0uWtGyh1o25Bdtq
ENOwJUM0B5hbeBUZR0q0klCDZ7Yz3Py2k0c304bV5ryZDKn9rSScQycznn29/FI1rzRFM+Fr8Do5
foTNHaTFfNfe37SKTDWSA38FhTIWUcwlNmt+UI5K439LynrKA5g88PiodQKUl9S44Q5hLxUTjKTD
779iEjj6yhIkL+5EBi6REhRCykGUoaJSPV9jQgeKKIBBTM4dE7hOBMe13HApdc1DXWU8uHnX//DM
YaJgJAKfYnYJI/mdFnJJANF8DsBk7W/vXi+n/PwdIvlMtSpsKGBwilwLAMOymkW5UUtH7ymlgF1A
G9ocEJ+BANJa81p0MJZYN5dKUEcK4Dycp+dqrNUsCPFck+v4tC0gFvfeUQjNVOhpgeMAFhQQCocI
NzJrqPazIzkSseEjsqBq3q9TmA1hTKGo8RLqYvj94elKTPw0wsaDQI/WSGlGWNC3t0rAaxiaFmBX
C/cBJq+OJtP/JqiO4WfeOCc2zD06YVQ+RXm9vx6r5wXrH76hjjkmqJOJsuzSey/kUMMfDbTnwASc
roMkrlbDpj/TihYlJ0yPRuf+d0HRArWuAlBe1LQk0lv9f4YxuyzBZCB1YIJx7Yl8R58CcPUVj+yJ
4IXhx6ViZluSkJQHnW0w5SDUm52q6AkoH+lXjCGdx0cgenLGkYWBKu7cOW+PfALFdNGbHndSuJXH
5JnoJlTgijLnmjpmhBN9PHUg18NYUBmYUH2nSc81KZXY9Cs0rcH4cyatHnJ13tObFM5xJ8fOiAHA
ersFUvAKzUN3/g2fuX+foLlnerhUnqxZCmrYzbN9RrcG0MEDbTck6fMcdTkyqT3FfeaVEXRmye06
/yBnaIZEa2SjSAGHNNEE6AA7XpuIRD8bfFxUS3n0Y5+IzYCtOOlI9DYWmZVT+hCDsDtF+5/sMGGK
N+GunAOdTsbaFiS12tuJ9Xo3aB/Wmnv7Lelo090z472t/MFiIvYJCGouT7ZOqODGZMsoRJB1qxOe
xrgHVaVvYY4t6Y42/jUtYcCrWu7Kn855fNf4/FVkshl82IqzBIlfIemmKzBu5aEqWGm2gGP/qAVg
G1YJ91FU92uMb6RG+ArzdnyCcXCsZ/QkjsIM4g4XGMaVtc0enE2vI2uwO1w7T1xEeze/+jHroGJ+
Vw20IY3N8d/tI16Ec11OpglI/b2a5CktrcQtLYLpV5MbmMJCeOXlft/tgBmN1Mv6CCywqZCxEkst
W09+OZhjl1DplMppcqM9+uku4YQG3syBc99CLz8U597Pb1l8kcE7ilEvoxTrRBEz/IxL2Q1RYQ9V
ZGG+eSM/0bNaZhc3t1gtCTgXjAPu47jJq2XAAZMN14UUldvd4CT6M8H6yPDs6AI4tiX9oWs+HWNh
qdxbv3WHsPQFLnC/QvKgqEBuCwe1Y1a1HOel4fIJ+NGJIWjFjZbpi1jPzGg+jyeJIQ+DShiKd80u
m+4s+/BYQTKfGboRQSLYQag3GCUyVAxk4tkCE7v7OpjGN/v4YOkAXInxKSGKMaGYAfmdRNcL+8Od
NF1fhaiJ+j1HH4Q3aDmQJISnUcNSWjgyWJZJRmGyO9h8a7wKbeOO+mS8xA0Jdoz8x1DVMcaRMwd+
16pHbWrQpbV9hmcZ5+HxQjeycabG0Ik9PvTNIpCfrxsWx0eMVlyRjVI/SycGwo0K4t7ibooWghJU
Tmwqd0P/4UFqvGTS9Xi3wqVPIkiktOdAn5wJxx5fZTGJSiIAvoz5gNr1b2vNuYgg7JZRfTvV/m/D
cGPJVzHSPtQgCFIX3OfbL9h15yTVsTE+zGWIEIbsDWpAvRu9Bq84pV/6B0yP7iV/GdW5tvBznmkD
YJN2mFNerAl308hj3yWjgnwNKKp+X20VfpTR8kUJmq9Fr4MWPUWlSScCh+FY02BQwoBCv9XO3pWz
AwtvAP0QrSfciM0Dq+G79I82/KaECli1S0fgyJSSH1h1FDYWJ1fhX2264PIqARyB6yE4w5Sw+Yp3
jT3uoX0wZcOxhYq4BzVgXAuIGx75jc1USu2n3pRw3QBC8R5qSPuTmbrJfvn2VYgGL4g/N1+M16MM
ELWzlnGCVVt17CsOInQWbUUReGnHZRrDJ0A26z5OzCOj5IXiacs2aIOzqimeynNyrSP/gubRi6Hx
PcAOvAhMNjHwlwP9zBFjBAFr85zqlYpKEUJqiZ5zkYhsUn0gh9ZQuF4dLkHZMjb2zcePKHjt3WOW
8WQaMy8Tb9pfjEeIeFH7CRcSDEuznJrsf0g1j8Du6iF0a1kGdnLiv+FhX+gdiKQjr6EJLt4HVbMa
tNkrboHzltH5Ph7PffFI58/25NaaBz1Fey+OnHqN2hVUGoTJLN+hPCZgX9dUpzHlUSkSmylcM0n3
+uq9OGxvo9SpGH7Sw3tdOw5U3f9GR5vwegdx0RwXO4XpZ7E5ApG+nihfsx9F56Mnc4iUNYKS7FlA
dpdyGz2E+C4aY2PperSvJ3qMozpRMtEGvw4+XreSzOUxfJB4QqjDd2qk7NjFe92hW7higZDiiSMx
L1FRE6If3/EfE0WQ/WTKbms3jDWviYDAYKRPXGJNleLDVNpSprPBIWOPgvHgkfDqmvDjdx6/K6gd
AWoQwSEQNyXWEIUUmf0188khE8E2ULTzkt0B+76Eykrry645wmlYpnK0W6JGt4WQaD1n26Iq7b9i
TlurgTfNuAys5x+v4uAhxVNLUvCunhFdhMGJ6l31ZwK9fBY2P/SMf57z/5xTFW2m5HKacUO88Yyz
/E71e1meWUcO01n7QcYh4ZdTsvNCALi3a3Q94kRaJARYpdEhDuAWLVWook/VnN33hDNJUtxGrw+J
0JPO9KZe7VYT3lpoAUGzpOHFMKXvAukuHdcnG7xtM7PKrpimhDBPmMRagiCFrWXE7fbvwx9tfRZg
aYwKb5la9ZPpMFwp2XYZWJUnZSWum7d4GdFKjMM28iy9yEf6r1GJ6H0svKggNzXsZmFUjM18v3h5
F3/jK57iXxVrCiCqVzZdkDDjSTeHNeeN9gxcCymauK3dxIWY4WN02yCriIC3ULnoM0LgACSOHxh1
ZapqIEFDVFO3hg6J+Kg61WzrYy/edIBDOyd3ZwDhFVpIXFxWdPR2LUXwWD851pLsIt2FSpZ5PXv4
5sFAfclbVs1Mjidt3nckfJaaajb5YAUC3Zk/KTo7QCWzFWKhfcQsQE5mz3SmhrmTwCK+8oOvC4Cj
X+CPrI0uy4MkmdOOh7f6jb/vpRDS27GlZIBnapk+f3XwFuGQnSmcYU/CUaya/CK47pOjS1KE9rUO
1TJfsP0XWirhKThBagHqZnE5fm4o1UPAPq455dmLBEbllWZ0bvTjLC4fuml6E6vQ+0Dx0RkamS05
FJWplU6FLoshpXgWh8DXaIKJpK6KmRQXUV90yBACRFVmvkzIKcNOBqfvvyirMkw2+Zs6JUg/Iyv7
SYwri6xEGbcCkLVn0K3UKZI7s1R0CFP0a5tDZXChS6rnHFZApHwJzs4u6uWqW1fBmMlC+hd79MEK
dVNZaMjDddc9J3R47p5YVMgKc5XNakxwFzSITdimV+CT2/+0Ua99pVTJHKLodZKWmSpFf2spXSwN
Gm+YOZdz9PA022DCIg2shx06XI/Xqhvt2ifygtdZSpr3gi1E49MmT4s7TdVjfyiSakThy0FYhSLS
vrgI1fZaNf7FSg5Fj5c7cAwJQf5dmRmQWsSD3WoAaYWbIaMo4wW6Xw5QmZI2l1tkYD+SgYBHMjrt
OHFBHXkphUGdT5pnB/SCl9F9zTlij+Yt3hcmAFZ77rgSgfBT7HctzlmyIhrYTYO4t8aPidWHeW5l
ES4FpMJGBNvls1R8JooUT3tEUV0WhCxoDcimZd/r32+eah2s5dLhoGwNIVrlZEOSVwSlXvvPP56f
B8urFZAa66uDyEvI/s4hg+oMj3lQeDHSHocDlfhhpsQkJFU+bfQhuAN/hrX62onwGZnfBnsqt6fr
NnjyZ+Nk8kJJ9crYyPnh+RQIKOwVZEugNmplFu5pls0yf/WZunW/L4EM8hORUb0tOmYWX+d/6f5+
CaAUM2/gOpMCmjxmJucXzqGXdtgmaFJEObnJTKQbI5Zxu5PmupmmwEUHYwQcqaglMvEgEAt4Un/7
PBH+NipRH5Gyz9vBSdblyRKmHNA/8sPVzY5t6lR/pKeiozvzeHzSUdcLq5WzgBbcLrOp/G7DwOPh
nJIaNG4JpsrAz/6dCB2vVlvgs1ISu8CJxfKgmAAomCDzANtbrzSc0lbZ3b8d61qfJ3BKGIXJarhp
LnLA4GCZpawT+TLTH8ixKcMuedEf9AaVkTC5XgUtWrbEmJ2Iqu8ENu+VSA671fqrsTdlvkhQj138
Wd+M1q4SG0S9SBklgpsZ+W3tQL1fhTcbc02sUlAk8gDTA1sDjOlNMJ8/kUH4IvfT3AxyPHgN1qJd
KEzetr/e5TQyxFdaGaG7zjBBK6x4MHg+3mmrTyGeK3wecCPE13/q02tJ63qxk9HvTafWaCnyXO9W
yQagw45eYRNtB/SCDf64nZL+2r1X6UGb/Oe0nUGq2gxL9jaHLSivGPcZrNOQcWaSyB6uSRchdIoZ
5agmRztJUp5/gcHd9jI+TSww8yRnecp4iLIZ8Ej7jo9fwAmjezowQMChnPWLzAojZnsmkgepjkGK
xmurGfith1uTiAR7OSmMZuCN90TN2AbnUxejCj/D0uzvyUl/WFm9o6ryhZKgftfarPm05Hfidjdf
m1izfsw4ZfoPxI8rbOrg/KtP43mv+hSF4PJByuuPxxUSxMIvSBLkb4SetVcD6NmHJTROrTnY0uii
m4SeQgoIUlZ6Q7GOK/z+LBuP9krP9n3gvEVxUr6Qtjt6EnspXR7iHVMcSGHLyJkrE/wwyoVxdUtI
EZzqMGKchde2b8qMozSo5A4plux51ugmYqAyKA5HZZ4Axs9zHbO5cZlJp1uNcqX1+0mi374keLBA
2LZkLBs8w38Q3vV8bfMi3drnJaunJsTOG4qklltM+jzfzEr5+PsELsEwZq25qX+metXzXnomNQbP
fSTSuA0nAIA5iiGILAlvc9PlqdCBHIL7oS/vnUObwPRolTLvJIfarrI8Es+3AKA3uSXlS1VHgrZQ
k7bZMTPdUnt8D0SoVRGUHHxKiZMkqMWFFyQRf5aTbG5VOoWT31pN9xp2xb2e23MDttgsgd3w95/Z
ls+d4R5Wh+jDCmMjADQpAmOfZ79Bt+RjoXjJ246X2NtBZYwtH1/ix5EkeC8glyBFJTA5dsMY06i0
/fPVuBHUdGcGQqF8/exRkkOer32eY/peLCoax0WLWvLkHnduY1lMuUiKE7CfRLl/bzrsbQgGPVVl
HS3U/vMdDoDWpZu1wuqr2ZzoR6CT0OCd1FwcCOiei1PTh+oG5PQQNSm8KS7RCTyx14UzflviAX65
Hsla3hEaJdEuXUt1T4ydiAZEBMKXTtpprpAEKWUYE7/MP5fr3IcyT8jBoRG9bGSPRaDDziDKm1GE
OW2PqiBGn7iHfuHWaHKmD8L92Ojc4wUXvRsLZTISJwUnpv9QKr23sRzoQLtD2lVEuIPXG/ztvc/8
hx2owLRGUkyIeAIhCrC/jdWDPetn4Gn0uO2jacZEZfzwrQD44VwmuPYxpSQ5L0jhAdkfQ8AuRXL2
LvkuGLXfZPPHsilV8y1BuvG0thwQZKBCckzzP0wWehpiU/Kz01MZp326+KwCOVXyd0ndshnIQTMr
rx1pbnkbhWBrDYI6ksnyPmUcwNfZsd1YjyBMpbT6NfXK/+9WM6SnB8eeHn50bDJ5FalHTwgN7YDj
2+KPDG1u60s8xAERiiLGtOu4sreBqn2Ifs2TZvmZ4drgcV5yoQMirK5C193T7GpliqAZK7EyuwYi
czLG86s056EbsAstr3oaWcJz+pLgKYmx1u3PHpE2WTUNxAirnA606RzOLhfv1hncAk/GIzVecjn+
hQZEq6vYCccfSVKvS6IzWASeGFlVwW72bQkUqb72uhUEy80qdYVnFu6p44/H9zvRJF8srsJPvN7d
CXH0wWGzkrmAvB6qRv1DhxFhNuja6H40XXZWpifY01Ht3b3Rqzhah0yzF1sD387xIGH2eyY4B4pn
7b1SmLEItE555fwp90NTV4fby6T2Nlk5xOEUI52DMJ8xcpb81JXhNO+ozLXn0IRxypCY67kSqNaW
QEixApwhA5BJ73FoxhOOxo3P3roAMC91Ap2Yw73MqyH1b8a3uAHM8Q91Xg5qTlpqZ2jYPX8xHQqf
1h41fM5hQf6+XLjKYzaggJSWts37sATHduWe8XgLW5nFL3fqUobGC6rltNISQ1UQP3iZW0pfubHd
waNvO4k6whWgOkjVqWcppuuzTWpKQyU4a8UWG4KZBTcAL6GNa0AKou/T2bpck45Xw3ipqS3EiDsy
48cO+Xcg3wNK5qYBNpW+whLNfUfZi2Tf9ZFQl5RiFVAiRxIQeCTgyxAWrbLDgSa+mnfjoD7kx1/B
B8/krt4ur3jvKUEf4O6JjP/TfgYOnI6bq5Xij8C7bo/fN4xXVQKv2ZRjg+qBPUW90G3AIHW92Hdr
HoEMADLutUf/QRuZWsrDDEm9schr1g/zORgJqSYIkHS65J9kJ7DVcERRcu6Q/W2aWDAfXiwjdNyK
DEMxWZYuVrvIsEHizCDVLezgeChHQpRvZugk30mZwB2rLJmtUFq1hgIiqNg0qcokCTd50R5YjZ+T
Aqf9IKaTuoS39lskqTD66UutJ7AfJs6JwtymJ4Lf8Dxqrg/KJfgvZc3OCkCje8PETn5/y0kh31ht
3f6nyLbbPIufBSM/pSGSB20/uMSMUKrjCxmCbUXtG1BOPFbhIYeGaGZ1CYyc/7AhAujkuYBmCVYc
EQQDgeYYbjNDJVvoTPxBGPVlXyV0uPGHj3PwapzzDU14isaJ2VjuQn2gIj7WxGtMeoZePXSy+Z1a
zldmXCexpKs82jPjYOoM8+YOa41FUbgIS/lqOwgal6ALID7SbD1daca9UQLTepJipCyU7lDu8FcZ
XW7OP4mbDb/Y5b8qPSgEd14NUVT1Y2eMh8Cth21jrFCOJJKFLGGyK/o7btUavOkLYsSC0ie4+ENX
Xo4TlCdqcADFMGw5whqm8YmnR+FbUtqEWUO23FA7GVseXThKjp45WiEcnapcK//W9h20mpUVOQNl
rrU6J28OmTOjjj8pdTRpNRBIbfPvclE7BfKcBndC2VGxLoUEzam0guGGjE1TtJVbN5hPOAife7+X
vw1tYbOL+opBOo+CvaZ/6tYcjHtzlGbt4VSQkeuGwtba9pHOUwM3orpuSbNlEYDYO8Fi6Zwb9kGw
2Cn9f+81760Ci1llsbOfilabO7BsRGCRNkS8sPrriN32xyCKGPDSeWTYDPFA0IX8H7URLgGOK/P7
xDcC4jSaKj7G7D5GxeDVEnbWL2ERbhfjPEWP8vQEaovypFiYJdbmy24OTcUkOVm5dhs/pKJTFe/x
pgXdR7Qi8zYfx7LEdG6KiY4k1Gegg33TvNxODlptqxRf8X3qDphKqemwzn/irOv9CJ9BS5L1MwtV
ovT0Zn1S9ZbqNeOpHpYrD7GwSLEBF3Ilo077+e8sdchwElfRJ30kyzhuv3i9azCXpSpVmmJgw8mv
PR8cBa4PoqYqvxk4HHSF8tgbsVVN10m3H+WH5kLNcU9P2S2iisKY7Sx8JTm9FNxAaVVLIFADduEl
x9yBhSUuFGx6xSVvsnF24oM/qzMoKs0ym6zHKdoT3kJosfJXbXe0o7fcrNRTBbSTkZv9ydB6VcBn
0n8ixViijp9++ZwJkCtF+7vrj27DKN5amM3SWLbNszV7k7HGX95bSHqEa8lJMJVlbPO7L6ZIOQzR
7ReqxiXvuMW3+IHlTDBhJn/G/10aCU9qVTiZGVcu/h0BFT5sb1T4pUoUysHlFd8vLAZIebFkRgqF
9ilqCnUtmgk6jSuw/TC9kFAoJ7PKt8i6YpSK5VpH6u5lxyXgFZUqdvsnSCa+Tpi7qFtAH+YMaNh6
cpMVGVmHo+vsHKLy74bVqgXJ7bcFQxCKWYsuy5hRhg0joiBJIBW1IoxLZiDkCr3yfEKZeddw3mFQ
runDjto+TjY2CfiX2IQlzw4krmFvo2MbAt7tmV5twHaKW4fwCCgqIgPq92vrKkfrUjxRQSWaQIOb
Fb/mcgzOGlOrTa+niPEfFgOdejZYXzXGpdl9ECiZgjidK0+KKKNXmHp3Kp285u8DfG314XRsOJby
yl6/8aOAWl6/8IVAyFLv0eFuuSPPPDKXeqvXbn0ab5d/PSNYGgKlwJ/41NvPVOW8gNUStiON6UC3
RkyWUgZjh2WvpQzNK62ti/R4AGohB9jY0tQ66gcYPrY1A4qUuhdR+UU6x8zeZ/acveo7YFupuG/x
2EGYpkSRQidJ3iafpo7iT//HZtHbY8Lnq6mAsnFZb08Tn+VIal223fej09U2F16x/pScawapIM0l
V6uK+O0b1yZK7Rm16v6R/qosx/jONUtZ84VdA4nSpRne2wdGCqiDV50gSXq4e55FjZVVm3+fBNV+
sKNn/EpysYym6OILpANvL3PwDEavNAOFyZJuOY/QXEy+kDzo0rNTvsYAwwRi+yXsIzyUjrGLAsdK
iw8CmUAJsPDWUSZ+CyBHPWi+TyVrbR37k6UUx+cxDAXunapww3vU6+sxPjpaMkrc0P1jf+ue/M+2
GZW3Wbmutd2J9916IFKi0xQuaJVLlk7GB1CUF1Q8UGJnPd2EzDoPcCa5fvz7m0Lfvf2otzok1pj8
3Q4Guf5JdJbTSBUyzlhQgyDYvMpPR+IzVBrj3uVoyAKRUqD7dVIwmf4LVNcSmA0e6dO6mfZ+nKhi
yE9+N5QN7jmAarwI4aLNXX2+rBogfYIeOmUq2ZIydWyUdH4lqDzMWQS0EjoJ3XTfF5/oyeoIIZmb
3smLXbO6jLr5WD6u6Vfd9skXGWZGtJ9uBdRixENtrDsRPmDa3GsYBf64rslj+P7Jhzj7gcKnZfzD
fs1wilUU1dosuAzmvMqYk0EKsQn1wjr0C5kcf8x7u/aQf77tNfCq5pJx2SeNCMUtPmZQeRsedw+x
3eRRanO4reWkr+/8ORtrAOZpK/3Bb3U+UNIWjTlnqMSZiQhphDI9PR4f0Td6DFnmaBTe1wKOqVno
6XjGHXhII18XpDzIKILdurn16US0gd+aO0RQTauXQ01sECjwWxB58yz/DnRfwOyzZEK8mOJrMyaU
670aW2MeAwuUKeAKHy3MlWk7RCY02mdj3GYGvTc3oEj/si0KNm8AWiXrgaYfxeY8wKaK8vz8xLYn
Y+BJL7Uca+mbGutKXrUXqNrXpxsfY+CC71RVo5m44MA0ym6X9iVqqvbJU6V2fEpLoYm+L1IlaBKH
r4NC6sofnY9Qh7xJjN0RKh4InLmr0oiPOX5NIekLqc9Ld1WP69SW8IaUfijDaPhRoeWiv716SM7I
T8FLnIF2FH17rm98VV1ozJWLW180fx0xChXzXI6fZX8/CBtB+9ZvEUGcLEKMonSiGff9nxeJn/OK
ykTAE3VG0OGDv8D4MdeVWouTVdf9s98VoOQetw9bGBSXRtkSvyFFioJKDuJgEbCUtC199irIum3w
gqZF11aNhKGh9nK2FaKTZMJ7fa+AJdos0jUxG9FFD4S4sVwriob8msGVDaxRTGKol/DuMVAxna16
9tfx+/cVUE4CBrJ9KscH+kZNBg7rvgsDB6Mk5DjYq7TYDrhB+U+CQVOXh9NnkZMwflIOlzXtojgq
eJywuo9yDe39sFOXMrBdQ6ruWAqls0aMr6XXKVFYvBH5VOtoFlb9ZkoWXcQOvjIPJBErXmyHhnwm
SW47esZ308brDnFBYsi3Oaq1gJEE57SgeAtWHu6Gvas2YBdiWi6/ctiF1YH+K0hbn81BTMr9ZGLW
V5cjTF6XBxaPnBX/RYnUo62fb9m/6N/h3584q2OH4SgTDpGUvwrkiYXK3ODClFWiBuJ/LnrkTJ/k
AtjqUjVQ74kXtYvnOkptIji5ZXGwa30ZDfUzx7IPEIq71R6jbbUMK6DHkhJ45+wXkgD1h8lxRx/w
hoP5DC5mzWul7vxlMxJFFmTqofDOR0887FKmqUfcB4vCVpR3vHLj6QCnFZPrEkI2NQVbd+NYQqVq
P75K5iBy2j5iVh7brwdi6XXBI9oIGMSRsCIp53Oe78pxxYaRY7P7sf0i+pgOdRDcJgxykrQwCFCF
BZU/BN+yNOQ47H8IF6TuyR4+3QeZyAtDOcaD6c+Qp/CJ+ji8F8yPJ4ffKPCvzu2QuCY37rLsk8aY
SBvkGu//0ojRNFjHwG0LXfPDDeU4PCDWyfiBdnSmSCOzIFkrYDOCUNcUOGj/0wOexDoq0qOHxW1f
HIjeXsRzOIU+GeNOkP+A8hDt+6KFz9cK/KBoKKx4A5PxZCcbp4dGPyZdvSdXPXNPaoyGM0wPpQEc
0gXkHwxzlbu5ZgEw3dGz/KfYmVRkfpMMU6rtpzK4XoBgPpIs70eZbVvzCwhWN6zfmn2u1wtH8oQ7
oZLBnO8E+2f5jSPy2PL4kNJSzmWsHtt1v6FKrSklExOUOWvw9n2kKwCjyvOPlfuIKbMgIeSMoLAM
Yo3SdQD/KsNzr9oM6zw4lQYkVlzzikV/bLntznn8DOIswwtr8eIquBTqgDJShFe1+4huShR3XK+D
fy9mi/BG24OnyBsIBulipy/01gcPoXcWlh87sV03MN1kyKGZ2aQtwRCk4mTMSA13Hu6uJ365SljT
CAhtGMp9YhD1Zw+g/o8No7wpWXfvm32bRyLwu4mKxtOAkhJoz4Crfe8ZQmSB/Fme8rgiYW8jEhLG
7+VfVebeTw+tHO+6J8WgaCgqlmNygaaj1Vx2LbRcDhIGZuZLwQGPMcULO8Lzufu+UUtOPhlhEIUt
VGvT/WncvtJl0J4kVeph2BqucWhuubFs8b9/VT2g259EBnepkd3zP92uZGbcwlsjZQQmKe1BipI/
I6qMeenbGcW6K6YDE6fcS68T/3hWpPQmLfQ+7QtPO0hJS/q6RbdbE9iW2df656qYADAiAhSvrD7K
qq5DEr//Fnj16Bilddp7uUQnI/DxSsdCIUKCZRnn8TG4eFJFpa9Jkb0KZn3rDuQLeS4MVhA34C7U
zgaUWbS7WIakdEJM70M+OkpoJGvsMrZlNJ0dlTsg+Lxv0M6QNEugHuyuJbcBFk3CWJzOcxWgjfbz
Bh6xGxPXinECGW3Erf3Ak4FzYN4rjbKs7RSmwMe/b2Pva/GR0ZL8p8mbidPrYHE9D0tZ+1pYn9cA
jgj669ktT1CvPykbuBivUNZdRejfPJYFhiqF/M2kOJ097Mbc7atfjQiloRQqKoNeMy3S+pzAzpr9
r/WIyN/moVDt8z7uVCLnbs0k0Q7qBHz3musUt3ade4AOH2WGFTjVKCNiAJ2iKy+rxCGeFL38oRen
JuIjBLy8rd2UkYy3GgFg1Z5FL9JDfXf7W4miTRxIHM57zoQsjai87EPlIYxEZZrkFmLZsfVZc4fe
C0kXea86etmcbXjbSkbzmPLMGixbtcRP18KiVnQmCfBF3xNYQYARzKSXeuLE/2KQQBs1YobXFjQ1
dqq1APzdm82taGxwAN3Ny7G+VI//iDVxlYS9bL48yJyOcK4bgrCZ76JcozRHboCpxhMpeG+O6ZbE
F/4CLp4N0tvD6reNeuO8GTXbORa0oAc4BKb/LLM1kr3ePqf/zvAH97VhZxREbcC6OTHV6ebHTEda
HSLusqpYytFtolRgrZuIs+BtZZz8kALU3DZQAQqwShKP1rwYzu6ODG0HwacKq3aWBRnRqb4r7veG
w6DfoGmkYY2ze0p3ISyayIgSSrUl4ZKUbrm0r6vgwpjQQMOMQia4VkCGvil9ijhnXFaZ3AbF8XUo
q1funDMuUSfCLQI86mg2iymfLEvBICST2PzN5gR521N+QIa7AeK1GZp3bWxmepSqhO6iKb6wiONx
r8teVSVjAJkUdNEfVGlKu7713P00JR7gF2Kb7ZRQFwAfav6MgwFQp8yoO7xSyU8wA0JpzyO72n4R
RzqJE9/d7zfOd+wOUotipkTGWlsW0QgESSoNj4kMCI/2jOdFuR2bvapOCis5u54oS/SOam7avyPK
9rrXGE+Nnpofcruf7MTBPCKRLzX6/BVm2noxrLOTyrFM8xqOVUUf4s1EzjILDbtHCFZxkoWwokso
lxBN0X/VCcNGVv0IRchngCk5HUDWSbU86VWoKYSrE4AxwE2brdBA/wvHaDgTlxjHyCPTd04fuYFR
lu5kraGY71ERNc8X4GMp5/xba47YUCv6J27rImBsE2838ys3EDx3GZUPATP3PQne9pZdSp4zS5OC
5JGoG9iC1/2zksoTelygwsOxIXdFLuxfUPsfjrvnA0OAOOGwoVR6nBYWTmD3Fqe/ggEwg6Vc1tV8
YSjzR4MJ18GfmmRttK7KHpmdt3N3fL0rlqsT5YvtMJCvpRf9PvS23uW2qEhj8jGJeD63ncmQhdbZ
G8D8tMD13T1b5bLRLk9E7JmMU4qmraIlUajHVUY5URlkok6H+QERyPYkTACe/sbgYqBXP6mIB63G
9rUWJwJ2fqqtG81iBDzuEFzlf7Irtg9Ja+qsohbSnPhVKQCBZUDPQELgTmtSJgK2m/o73J4Q4g+R
/tQh9W1620HAleggqkhjdZ98Bv4bSpwacFMtWx57vas2lEE5qwEleYxqULOR8fHpFHdeMZlrTaNU
TjgopQb8l3/vF+PKebqNd7oRWViPI+npXUuuJpCZ/qWMT7FOrLcDCMmCCiiaxnPBj8cKl3qJPK69
boZcjaNFHmmanO2ggHJtLiHEO4/9+4zzAbq75s3tGmhT1ecTZgCFmmAR81nmZExarrLZbfsW0WHw
Izydauo8SCDUaqyvWbnbWAt0Ur4OGGJ/5ufeNVWcwpISzdAkfudF/KG74XXdPyxuL6ALtOFHtKuu
xm8TUsER76y7yZAFKxBPBtm3mIu5y6hRCeBat9EozbBFGY8fYlWu2ealAOlbYOqE+zRTWQWVPmzo
aUBGbV4isqERiba5RXLEXxqpvDCeHQhwQXQmXNDvUrDOf6Doa3GZMvYXBs6C33pzI7J2nSCzsaiM
4HV5XBWGMJI4X03P4/9Fq8SqpELEgTReNJUzBt5l8r5T1EelaDu7qzFx6L2Fk3OZbyl7+VR/7HLK
JbgnuABW/EslbmbwKGvQoc3p+Nes04HAzM+ANJ+UN9tyQyGXP/ZfW9k853IvVpetZavsp7S3x+HS
AVQe81KG1GxFgOSm32gam/poittFas9yy3ISetS7busTeZy87q8+QeUBV9SI791ulH0j73mGrZJ2
WA7RYAB+WWhDbf0UD42K1ooiu2DqQ67anMmBDUBWEwYcSW+ZGWvJP2PUhZbzVNziLKKkz7QxUMIn
/0nCxoa5hC2nSRB4NGckwinXhIcY3f+7hm5PiFIIUylFV7rwGwX0TblzljIifoBGOtUxv6aIROKT
LbL6CZpEJL94u5QDHnYflUolGw9E19mdMI4tAxp93XvtEv8bqAAomWYvI4AxdNiBSAYy6T3T7GhB
x64vM4lLGyKI6YheRXTzL4BzU6/1VFldDWJB8v59doPg4Txl80gkmLzeA0dbVVmlIkzdB32oZ4Pe
zgezI2qLFg2Qlb3MgjXnr4v9XKLL821ZVszWdfcd9/XmkryB2Sk64cK8TmwNK/ijoaDACbG0WwDe
/p8L6fGaHLpJn58MkzPGDJ4+xzX8X3LaZNlC4NPpQCrgABHUC9dIwuTIhUJtdR3Z5TqgLzXhA5AC
VJ8R+oQiNtg4+vyx28JftNS1wKXcC/vQJigjVoM4a+Vf+E9SaRnMGG8u9enF27PwASvQWhmuN0lK
8x53oZoHnzqFxZTcqdRaWpVOLDu3/c5Av5WnG8nyPGq15ojjlwFdb3/Bo//jqi2mqEboXCYqKbqH
5cNreuaxJPMapYtLrEc0K1H8NVqk2yqlKHmwiDUGJvsGyHEYtYFHTYTK5IaGFe2pPCJvTPALOlVC
ETtgznVfnup+l3+ZrF5EBpEgYf64AvoQiqxwwFsSOsT4Q7VlFQMotHuh6O6HadW6UoCWSxom714K
gpC5IKoExqeJdoR9HiFWTTg1GyRrbkED/aWfWdvB4vr3MR/ImHmJboXdNU27Je0z1H0xXPcnuBQE
BfMAF9GfEa8WMB93MVttKaQOVs9n7ufIkKGwc81Xxtphza33utybyFwLoIizn8KNP5ZFr766aFNn
CWFmW0u5c2CuheWnL/Xjw0jOArGKvjfxCsf8qnAKb2mRTarBrWKw4s34FEX98v82FoV2s0bSeCRj
s0nFqzrx/VfIEN5wJ8pCU+/XfBlcj7jnZF2UublxJYl9mJQ4BDeB0G2Rt0lULZuAHIXqSbVs5UMj
CPLukAOdDNTDYAf5MKWjmdOJUe/APzBgM57XLvLCNNr4E0ebFHSg0MRq/u7FgWCmigyCVqGx4EfH
dIQIWZTOklNFt/4mVMoZQq+dMKhvy4MVYnUf1B6M7TKjzBBcLSZcQEXKlfPLK8lFQEoEI4sDQZmz
kqgXGfpqKSjEtfPRRIxeBc2HHiusK9rvPRPgmhW1N9SHOrFJH/btefPoZDX3yOxA4iMaPX2dQz0S
GprJ9C5DjJ+WZr2vRWo+8bgj1S7Aq4ys9qUOlxc0FVQd9Qs4kiCOLL1uxsZ1LJxW6b9yc2GBS+VF
H4GAE6wU1irWxVYnQs61yWyLSywk6VAAPbFKdTnPRhLcxnKLCp/XrHLXNHkyrwVTyVuSHELmd7Na
Ggwz05Ajyo8eyt3kEyWdh/fCI5L0v+p5X0Yi+iD2GR2FuVQuSnv+1pbxGffbjWFWgDsP2jvrXVEU
nAdVoCUPsKMSTcZigpThP6oUM2E4mR1Lv3HudaHTSCzMAp6URuhQdKTYfrkITIotmNPgt7ew5Dm5
fi80RsEB6mqIS41EpqU+XlmONWbg3iBgqagkMNxcvxnxELzBhybydx63A3gRR1/XrjzfTVqcIIz2
zttup2T9DSPO2RRdW12c58s1nfpQ/crTArT+tRQsqlWFHh42dmqHn7jsdNhYqRR1nucrPxGyjdGi
OsNdeUetNOs7yC09GL7zuG8WykDOXDBkaE6uS0VA/vHKNljtwq6WCsUUQc8g996CMwt/GeXknFg2
GCcPx4DT8gGqOiQ4dUPGugKK1HEldHWtxhR1m+R4oo1NJHCgf2ITLxvS3VqKmT9Q+Osue4MyiWHy
qJxXcK0uRMTcHnVAp0d6X9Qxwm71HPuBQ6bdhY3nMzbFfqzmc2qdn1tswRFg2Yy6g93JgY4e+QPc
2DAQ5Hrqo2ggIYeESbIQz7mdli4DtDSffyIrey+cQgahBzv7PyEllmMWx8Eg4CZ7nnYA49Yvltek
2wmA4rH6NCwpQmF6OuGzpOLVMyGcr0K9K05AXIyYQ8IOk8/93sE/r5NYMVYjZMcy9t/Anxq33Z+Q
XC/AjKE0R4HdjA78GY4rDpq5fZzcY7yTi/7q75DQ8N2CgUgCnZDw3VRiUKOx78BKuSzuYlWUj7fw
vGnnvFdzD1EZFWZ0/UbvvrpKogLnWetGct0w00cTO+rtpgVZbgyO0XulBV2RrFiGBL1PmTuTAGo5
HmOIjWU3ec2QsRCt8uIFhb8mRrm7Dg+Abo8/xJs20Z1xFe1c257rY0TJttSb/WFfWIg3ovkcms0R
FQDl5r9Dh0T4aMTH3hXJmTdGbcY2zh8UpX8sOK62usKGuPXflp+j8P8sTIbbw6p+2DE4r0bD4JNT
q8XQWmxNcXwO45UPoOmkRmdDqQuN8BGQ6mftfEu23qO2UoZdICosQAwOzwkUbf6AkQdYbY280JW/
Fk35kMTatt42w9dL8WyOxexkxS6/J8j0HVoBlO63AyrQsiFz9nrxTVpnUD0Cb5ahO5+WmWmpyvc0
ad9+eRmrD+o1BQAPhO3CNGHBlLHX+Wa3N6hR5LyU1MsxI+hSOTUTS2AmSJRZY4UY7JVs1GXoc19w
KLk2j9AO1wMG3K2YdMousV3/DPhewplDjsUt3ci310VNfKwS051zrgH3JMcISf2aaMktQwXGJGiJ
AsnSp4/mMQPShl9/RVfbJf6bRjJb5vplxdoUcjhaVsSEUoURkdnw/NHHNjRLWMVpj031QaYF+fmL
CyCdX2coMMTrIgsgttxD3DxvZKUc0F/WwhZzxb9LSrgBZRwMVDoHHli2K/fYNN34J4S8pCvLvkJ8
z5Ftb2Y5GBj5RUfQv6dZw6GgyJmEtQfaGWiENCSGHLMHxyz9EoBe6sTQE/BEGj4FfmyaZgVMXLx2
7c5j774HkFGourdEZjtFOf9CDg+ySpOU6qrOvn1iYPk/9SBfEAYMxEu+2Hr/NZDbliaMmxm00D+L
ultOp/dHHKmhEVohLVPZBQKJ39nrnlOMD0fox9x7C/cVzWpBhAnEwL2GkCesoi9pBdOd+fyIqvA7
5//wYXjcZaiDPkPqL2KNMIEJmnrjrVI1X+TGfy4pLrdNc/p+BJC1sW+MLNDaVMUWyWFqAH+5+cGi
HmM6j+i3JAYcEA1UBzE53KIjEf5W3tp6Amk4m5dhSIY6EaWzPhgG8T3Ux7rbccOUMd4seBDFE9xj
D0dvGdQkoGosyr/o+p5L7I1geWvleMzg7+PHjuZOb/VWLS5i4NZcgsMBgVQhLg0QX0sz74xEmMOt
KQJUsnCq/CelXDxTeSN54il2kZTrHBv9JckgdnFukOE2COwUaofkclnkfdMyeYux30Y33z+GYMvW
9dXWwzjVmXy+5ROkj1vHgoGknGUOq6I18/rzBxHTuoeeaJ/3mDlh+qcZYNyOw0lHswFnb9KpTj99
vfYU0NEdHLmzWbpewUwjC2uOcymw2bFbtb/vmfGb58o8MhcOwkdYj4R4vuWjEsgPRkr2VMvD2+cO
EOAUyUE/USyRM1/9gpB1Cmjcp82w34On0fepJBYzC2wYahXy1ilXCTLKSdCZPzTpfOhAj9zoIHz2
WiVVFqM1OqztOT/NEPn6XPcTEdq4Z6LZw+EIve7zdNSXGZYOgVU8L4SFk1dWc3unKStO/VQEKKRG
uKh64U1KPEz0N2nGP+Hzt0/sksjC5JkG9n2QZaJyZs/8w04P6+BkBdDyxE5G6ShODWul36uq/ZMs
YXTWk78G43usIR6c14pB4sv85qHyi0+ad1tekXuE22OToAea2SFM2s++0Pofbg1QvDnrW8Ax6Ggr
hUGnLaF9ggEwipoaOyb+nTyc+Nfn9Dl0M4fqloyUUmNDMv3uegRfga8e7T5FJszbyXhP0i0J24yH
IGDNCPn5lMIO6H7HkSwVOa4OH6pm7Zwb73zPR7nCp77FPqiQHM4fM9wB4e8NZT1qVfRr70D6lWTm
TAUuYHNy5kIZX0xoqoJUGb2oghHMEtu7+nWQHuSX1jdbkB7DbDvlIsgjSsIsCTNk2UlPtC6GoLUr
ZrKMsoSrICDH+R8B1aUpy1Q4CCyCyS4fAk5+aRVc9ZOXlsvF+HwuVU0++siODDTiKYjjBNIgu0A3
T3f4SIEbv0OuNGht7yMRvLXQXS07rykFqVR2JjeJXA+5SSZql/GNM0iJF8aNn04fh8mKB9X9XH6E
g59Lc/4TEhKBub9Fj38BBKqya0+Sgda5jEZS8yn1+V51QOlyHwkGKN0STR6GSHNxr78G+cUOyoEv
k7E/agVWIlzdSulqVVOQkcnKPdlJPnShH93J1NBH1GsuTrsL6yMOEUBse8kzIBRQhj9hlCSkC/AW
cYy7dkC+3CVJ8kCoiinDzOf5J+cBJCDmFaO4/VbqABwsQ9gYuv6fyXMwxdR9jsnHP89NoFImSIrB
M9ju1HNTdobGFZ/OxwsSDGyibdYunVaiuQ+ZaP4AT3cWr224YAHPhfqu5iXHkCgvSf3T9fReCvcv
tf1pefcvVmxlDQD819flBmSZEHMgodfj7Y0VSU6QKy7oz9PsQRHl01UR13mExnoJIUP4BVdKcuaT
fFvBsW5ZhscTQdYnCZSIPKNVdLU+mPdonRUemxgflGwdCIMWwgXZgjDeR8U/PJ62yCp1dwEHmhnO
kAtvHDFh9mFLEAZvJO9Rq5emaNJhwa3QzkxAlXG1JfTOjYJKs+knsHNfmryKhskp5LqaZqwpCfYI
7TOiC3FTOCZOrMP4RpIUJ7uIrY+w81hYf6XQ5ucMXv62tGpI1M/wu3vNXi0OyjZNO0v/HBUZoPHW
6mEFDhp0ccwh2xpSIPjVtCoJrQF6oxOC+dFuGagxI+DU8NVdwyEVBgkIF1licAjD3nMKaBQ4KCQf
yQy1v91gSAd7+3q0yN0HI3n3uRDYYAuo2n4e9cUj7tTG8M1ZQo0MxCSYNzHvIfCN09xt5SIZ1iV/
ZZhEMVmH+ff8JOSOWuB1nrGXqbowtc4ZJuwzxZ9IvgleFLvDrAjiUY/Rty1CdPXXAkHTCN4dI6Yq
jxHfL2MCDHPFQJXOyYW99kN/qH2dMdmt/s4XXGGTrsZdLV1a4ljDwe+Q3KsIud+RvAva9iiUDxeM
nQN0Y1V1BQrJ4VQ/1sQ81qYXQCnsdxsXNYCSh4Lx05uYvJhlMGMuCINwCLn6MQkO5bNt5ZMQw2RM
62QSc6U5odFytlkIQss4Rd2UlZmy3PV+VUnqnH0hFG1dbvxASlZvGirRPg3BAFpfchyFZNFV/WUo
AFzKKw3zAZ88ltHjPdsh7uLJpduWXvxfurobk4OMAkFYiaIUp6PFqW84HHY/LKid9AtPeMgYVvy5
FiPG6VIdrcl2p5ixIXXVPZVufc4aL/Q/3lKtJffPROqQ7dBzq2Ak1tFXiR7wI/GU0KwIRNgmBoAp
tpMFiMMa/QV2FAZuBrq2UWTaP+PRflcfijbFByMdkRSOJSNy/oLYZM6PuxgoZmz07CEqbFM5BU8g
UwBAC4kB96IRD4/oS3KHAGRvQiTs6fRyar7TPsnWxgCVmvbgkxqH92Hl+2p5Y/RF/uw23O3tX3h6
4dyjAVEYLIYLdTe1oHTiDlrQQXbup/isxEn7790I6hqIjiY75oIB8+WAdg2dlE2qHcR58ikTDvtK
NdCgbY9by2M+lSI3ibMGxIt6dt2nVq4rUsFHtci8/aczgVCUpBTgPONO+/rYgDI866Kk7jbTW3pV
3JIkCkiaGyQeB31c3Iu3Q8WchnZ6uTm1gxRXiKoeKz4nw0uA2eiKfDRoSpRgjjpPb9Bhq6xQh8cE
SNZaynCsgcUPnq9nejUFAivJ1EdsG5/akjTCElLbpA0rZOd6aAnpuzpzSRkpfZ6eOKz37Nz6IE/h
s0BwwiOo0Tk7iCpoX21IpkJYw/zNfljGpUwNvgRx+b/DiO50Fltd9Bkkq724UFO86mzEKgMhtlKT
AtGs4CnZ/cNUocZUCe1B03TAEyjUoMTwiEHMcm3zYHw2Kyq0+6RDscJW/vW+UULZpRkxMOx8n1fm
36ufkrDis1t7hyt838kV5/ER8tB20s1NCAadGNHSayFCz5MyLNyzinIeXvYKgkkz09pQvWo3AsKT
/+5uJeWcP7UsYq8feIEowJ9LCauH1xw8FzVfbe3e7oW4O/c86OvvoxeqxC3N2/BRHBdEto8AOfZI
X7nM0wvMPiso0NrndamUOCnGahyhmHB/3xi297MLN2fklP08JjK84CQV2CPMgahzPpQaSwDAwNQL
yi99kVxlOsMUhr1GnqemqpFYEL9Psk6xJKMZ3osEVcD+ImyeVANdI351MpI+8521ag68IA156X1h
JfQBEhEZiuPJ0cyZC/nH0MDPm6AoF6A3u6NRJDVw1hAE38KseDPAiMmkrIkhFa2VQgcWEN7fPQb/
kPUjE3irwha1LRNIHGUzu06RvDs/qj2DZ/Uj+ddzvwHkoN2QO0JjgM3kZlXaqLLO8MLZjcIMkf71
B03BBi3frJkfc6CdDo0bSVKLBWhEtrxgPLJbWLpiYkXa2SD5rM8Otngb4/syDOJ6QMii8Geu5jgC
eFlQfEvp0V3y3ptSjKaIEy8/qFdXFiooxuCA2egd0urHnwFH93KYB2rsbSeajGQv1msYDpo3x50U
Ler6jreUmUABDHfa5pG2zsxYKXOT6MJ2n8A2HDY1ZduhZDeu5gqSqSn4QYoGQBAHVg7RFwIuWozm
f1d1smT7WwqkZ7FPp/pf0ZlFoE0++rFgaiE0CrHZZg2gqBrJp/LlwZQ/lWxmvL1S69WkOJsMsYAa
kxOxsIFdimLsL2aZtX1jh7XlVAw8YFVgAJEWuDtVCaAX+ftWiFv5Ar3yj6+kryQh1d+NBOC3x2vH
4Y2e2SlFldBydJxXHMDXxkjQnWZiHtDS7pSYRkRwhzSctvg+rdDxhgxIdohO/aOAQF+BPziC3IdV
ikGUsOvNZM/y8BnF/liK7W3Ze5r9XmhKucYn9SsCCCIjv0lxvydcks44jjG+cw2k/5jJIt0awpkJ
pinHg6vDgbYwV4Y8gFu8WeGh8I0QphEmR8ZztjU0JzWQahn/J522ZTuKqHq7VfCHubx1DHPpFI+4
CBwKY43C+kXMUSyJoyc6bMTT8cOazj+ITDvOEatvY1dAN6/NpS0s+q/wNPTKPWlzMEKTvLn4GAh1
i6a7bjYv6Gp7xgwA/yxZSwQPNwi0jetrPPiSJgtEVz0rqrHT/eUeZ7SV1EisysjUBDKzxhsmz8ky
Xy7qKZmJbM218T0BCDUPJwUX90REc4P33mXpXxsCg3/K/SF00EOOaJ5RZsEDEy+Qwpq2bVglB8GT
2A7JsXUDoZk+u59IcV50IYsfmr41TWXqJVnrxWWTzSG6gLf2utH4t9UcYMBLV6eUBHMUcHSG8sXL
eMxhepVyEuRUXZBTW13GY/xrZR8WP1I9RxCkbCg4V3O+eClxB0blphiy4+qtJ5mOBxAJuM8LuCkD
Ov9AeuX2u3vuhJ7f0aEDNkFXn7MFxSURajjRjkfa0aiowx9kTKL3hOm0hcIceB80mezFTeggj6mZ
x6vnXYoT4R4W0ink24wbEuBwz95m6CM7XJnKRr69FNYPdaO20oqyPZOdHnG9ktXGmUu5otJunS/y
HdN3BulO9FiFhatOfNBYyKjmNSDuH9eqq1wR5rAmEzCLdsfgr84GG4wLNQlPN7qwUjwnhxefxatJ
DC8df71Njg2aoZm5eYUu+0c/2Vj5lxCm6vgRq6o+S/hPnvsSnFuFX2YCAP3YjV+7h66hvPK+154t
t1k8kWo+aMR2xhXrA8snhzcdTfgjadGFVN8wEAskv1DeWNQrETGl0TFLFjZuQpL6hPMUl70PU4vy
Dn2ofMi3Ex8v+Y7BD0aDbQHy/7tttNH/1Qp/CfkYuhH/ppykgv+fIXxV12hnbTRfpktzmB5ID4i5
tMvv4VWsSlIsP6KE7O71RCafxlSSkaq0JnXDjD+cZkftu7ELuDKUvED9mbaiJXuj6v7dlOzpeV87
+Iygf/p5dkVKIGDlzYKdnY4dTV+IPWaMoPJTaV2Tgo5lhOxmtCl685UF+F+HkGrfCiFt/VjBkyFu
fi8AUuJgpqv0dmNEqzY7+xVgVqqLfewqAdv0W9xNwG1MzQj9iL1qm27VqXN87bXl9X/tlKkwMqVV
zU4Ph6shtfSYVRemFhn97iw5dJ2eUabTjOHXqrPzzwyCl5JHV0WAG4Qy0zxdmzRfpb/IMTGxyqp4
9a81MDhv6EThGVEd4C1wJgR4E+vGLV1ti3+pkeb1LMU4fT9TdCGAv8o348urOb4FmJwpaFs4HBuO
cM/ASW9xSqZzShCEyiMcCvBlxcRv5zleGim6e/NogXV/vVnmRwLXFlzhztB4ZGfDAhxyUGPFeECW
kvJ2+wY4K0G1rqrJ+UwBS0z1etcGPiocIvxT17Ugq9IR4h+DeeWBKaGPef4vphKziJcf22flNqaK
perG/jUEt1IwTtWNCAWHiqk01delp4pjXOddbdPIn6OdSkUZR/mzyBd4hbncFu1JWIn8Pn0oSMVd
vpQz++30cmhVq2ZlEyP5OBPvEB767gE97FoEFZjUepqE9Xp/A4VOhA/GISk0/lY6xvUwPCxIupVk
qwC9bTmuDwbXoqz0u0Hfg6j1cn9EACk20JFipcGJjezn9aD3mCtOzzMjsDBg2MN3rp5TH2Ns2TGN
IWXUci+vapFyqWtrSQtnKGTEyjxaNS0/XBAdGazJrvEXelCvJQKheHHa/e+LPfN9Mhz5lEXTYuYn
rDbUH/r6Lla1rD5gRRsydhFnlk3mg1nGUF427awubHSnv3mABaXWc5kRVBL0m4Y2PszsPNk56NNO
pIoAb+ZlX4wUuAiVVhvO3OhGi9ukHMQrnoZgHG/KqB/MZekXi6jylxFeDvIwKj1XqLr36sAdJY/W
jchndJ2NM5mRC9l7YWpPKvcECQEHa3Q8De3LO6rFmUgsfKoHrNIcawGHbLirfYvJchqJsbDyu7Xa
RFK7Wi/w8mNia9thV6OeqegW7wAxmsNBW15TwWBCS9qBToq3y8AaniknBjh4ZhntDeP89lhvoGVy
4JF3QhtRLlQOu6rI+Fyd1bYr+KxK5+VKiLSdQI43UhbZzx8+AfTvxFjGXO/XEWfKHRWK6+EDQUcp
3H7mhqJqdJDPZqwLgKD/qrF/ppSw9kLw4qrjz6esjaADhdv8Fv6ACF/iwrRbkbxP20sqnEsHwEfs
Io88FfZbj1o7RyNpdZVDCic4JgmwCYl1UR27r+p7uj24GxIqu6wxfbIyb1lgKDr1lYfuVuKDf5Zy
IAuXBYBkJwMPZdoYuIsF3T2GsW8OkeTuOoDFwiWz5AW+AAFv80g+ExIBnavev9hbwDUldXJTpAde
QvYrrQfQo4iH4vdR/i42t3s5+5Axi1veTbA2Lo7QQ1PO8xK9WqmhlMhI7alVJuItOasEkOZj64KA
aqSQW1+FgPRRqQ7B5SNvunbX1Y40HY4DdDZe0r7ofpYUnzTgYrOhXOOxfTWc2yhGYnLZbyVQE1iH
XYKZYbY9sKxo4yd8N/Z1h8Q+oXstBtL/wKdcF9fxEgTgYwhRJW7NU9fspJQazQ38ur3r3n1dSstU
FinYMZWyErQOOyeK2wLVkzh2xGJm7pXw4bEKb3OisIvpm3RZO5hBJ+PvaSJPBypLjRY5GKIOuzYJ
DLWedtog1ZAImQOIuUifJo1cLkyq+hVTFX+1IxjXzhPSerMgbx9eutqNYPUJ2twK2M+xfdXpp1GL
JL2y63hSwpOhc5kHQET4+hpmdb6yzphmdWdkk8j+5S0Uv47RGUu3PP8UuW4Hd2+W3bq059RfZxN3
fS2z8+L4jpqo6meCWGWUL8Jwj+KwSvFSviNII6gNGk/wr+J83XdJzDP63P0fh7lu8hvIxg/NZ/uM
c0GuU6nuFOaLhSdKaAVBlmoRTExkKG+NEqeWK+sOGKGVQggxRuWODJC2SFUs7Qgt+HTHTFLARcob
4VQzZ1QcfYm02KsJGx3W5Gly2HspfezemgA4bW2+6Thxv9f1PAFU2XyDMT4U+vKCxBQaJOgYwBDD
RZmxAcjmJXXNUEdao0rcKnvjqnE8yHrTRYd9UnCL5EUrdysmyf7FKYRI5xHP2ggvhwvpJnaW6DAd
rNZWLYbk0N4ZeT+EtJY7WnuHXPvIUWCx8vGYb5JsPJscONry9m8tgq34cIoRJ1IhVyX5Xd/bR7tH
6jmNvk/T0Gek5+diEJ1Q4jyXsQoOL1mM44RwsK5UKxSFTz8nFAWPJ7QC3mygngrcd6qYvhKVDV59
U04DVSSyMxvIL6kPwsdMLSeMBfnPX1UVAGUREGmuuo7B3xfNPMPpEhA3h/JaSUfaD+3cU/M2zztN
YR6t3ozGD0SzViEuKBHKDzz4jLFbcv4YL37lmeGafmDSWbb49MPp2sKMaKhZTG7oFGi3uq/arKc2
Zt5f2y6bW+s3RLO+LzIV0sVYhIFLn5u3NLEOu8rFr5QY8oeyF7A29ubrZFUfnoM2zaqr5bSG2iGj
2mO1PQYIp7jnFCK3M7X5xgR9WVOaUU4hUt8oV8IQRzHIJ51zAjd/nhCfMlO/Q2GQlupPPYeafYz3
KYky6ehZjKx5oVUCSdIZlzE9KavkXeZxgNhlA9eSv8D7jTrc9SwLHBRnghPHVdajar2tAiv2h/Ky
cJguaDd10m7Ua2VZIGLuB54TM3nT1p0X0Ls8zWt6SoeSed+xpQm4K5u2ugeFCX7t2xmDVtiYKOAN
2f5QWapTkXrCeg27pb/yeLmzH0yiN5/CrWxrMEnrcvJKfsVEqHK7mwLwEOH4mYhJHDQ4AEX6/pdr
gYDfDsattjr1fHYDhabxZd/DdolcK9FAoc7Zf2jQ9rZtQ8Sm26Y81LBxmMCbBAFQ89qT6xGE6Ssx
nVDTLTEXUJUwuGLv+i7VGB7BtDh+L8j2LQVa/pnpYd1hP/KJRLnmEvYrJpGCYRGHNebpehL3BYBS
nYIZhdEdNTjzfA5bsao07lNLlvTqZuM3G+bK2wUFeRVqDNg6imsYH+VHVUaoiYuVf0swDpj3bXHL
ztZcQljln3DNkyA8f0uKWieAFiwFdmR8lDIRJKr4uyP9YCGLckB8NIsDlaKuuq6JlQK3vhReH+7h
Cu86jqrV1ypuEQiiNanmJplnqFi4k77RiEuYurlcoOV7un31LPpGDtxtzBLmNsUHLe6vZ4TqM2AA
Hlt2dU0T/ohaZsxiL3xMgV5oXHojrAogaxmNaWhiwbIAUBFzTOfi+izjlE/wSMyVSfiVqTkdMOP8
Zv3zBf3WusSvqgFz9BZqeOeMhQulfAy9hYfJTSmJda9TwxPR58Qjwg0wmOiq59azNCBJs/1Rc7mv
FvoRKtgmf+IQ33fUkkEhFauYQJc1DYsKVUsdA1/pRxznZrHk9TLFB3ikf3qQHGZ2x6kc2n1jzEom
KeqmDz3QFdBI4Wk0L5zl9LILKbI30+3EdgvJxeW+FkpADy0ZsVnwY2jcZ/yBT8+78/dm/9u4Nq8Q
Zsq8/DDoXiP/GSU6GBJe36nMqbRLYX0hqjHLe355ByLwzJUuvknOSjSs+TE6abVKq/9rAOij0VoB
HsfyFXC1gUMFlY9foSUWaBqI5Wfb5TEkZrMnkcMxmoapMjGEzDCI+Mz5GTyAstxpi58B7wkf8mQr
GLGpkkEjbOXNQk+SVTJFT2lalwwN0eWCUC1pb9rGiWjhkiF8kVPsB1nY8XCwTX95bN/5qwp8OTs8
/4KnBxGAfiEq1vMqZQJWu6h7CiW0wl4gHeMggqvFSRUS0OFQYnKjWln6tX2dwfGlMR/2M2v3f5l8
W4mn8mBIagRgEyRVI8wtZZiwvbaCg+dBCBLxlYH2L1tSKHhBTFmCPAcknjU1BJiRtxN8zIAN9rbT
hp2lMP1mLyZBZncGlTFeVmhYVyqdTWKWrjV3le4dMdywTsoNa4eu2NezPbrXOdgnlVzx0aBljDIq
Yyy9IIjmSYMLj8i63BmBNq1yOqVOwo4Znfj/SddIAJ+uQ17skrWOTkbch4xy1rl2FADd/6HeGvV2
no5iNvhaZOVj10CehBGwTn5USlvddagWNuiUyFCzOlg9SPnAU4eFkMX1iQt2hSvgt4wwkau3xy/r
zGkGC/Xq0gOsc74wXU3UFvsCme/iWYZDl7SXalPcMiRKuwwPKLCGiOaXhJdxOC8+YQ9cHybAAn7V
/HVzUof9CFmwGjg3yUdMGIitllgF78HmtFppXVP7wwjkWSypzjMp2rvb0wqlFqB2dPcSuIHGDm08
HwZX2dn2ZLQQsyt6P8yqil0/Qt++9sRdDX7MCQyvOnQEzlRW/QEGLpUrK9PLu1csZBboBfm61HBY
ALnQTcTNdKsWyc8m933AnHrglQol73NrcoYL1J9WgTAPVzAfjxZwzIndizTGDgLgihWhlwYhMhFv
W+12Mpme6QKSYNQ8VJwPAvoJu68OoQmPhTmsuPrzGiqL/VNTnHMaC01bU+VefKkXj8yfBxUFPq/b
tSr7Ut49w5ulM4Aub/xR9K3iY2Zla2ncme46BazaKQpwjsSizo21H118TgqTXZ3cljZfdC7dkkNx
J/8PIxCEwOR5GvAjtZ2dMU871Km8u9S3MkHVbGExyCmmnxr4G9iRFgqnvvoffH1m7ZBr7Dt6Rezn
OHUtSkZDJOc7uy7sB2pljXiwdBSf3jIU7ZOHUJP/0OjLO9xvPS74Xb/Ygz7UvRYgTgJpva+9f45p
sdgRNWefUyHo11XHE/KldLp92EGZyU6BuSCNhqzpZeZIhBCi8I7KsoLA6DVZWBn1fEKbxNW/qJ9U
tSzA+ZTn8VL8ZCpIuhxcmz6scqYLPo67i12uNvuBkesqye+tDblMQ2xpSNHOZbJVNRPRkt2YUMBO
tuycnNJpd1Nxqatae7G1WRWW4xXT4PVo0U5vtyLqcP84NQ3NB84cl1YH2kovSqVFT7KiLNVgWcHX
K9lUBtbBV7vdufkfAGlnKbMOuIBqvLRC6wRFXnOVNC0zyAex+rJ/EloJ2kv/XGRcOY1DybHWErph
Tf4uTB69VS0z93tLx8Lh53cWzqOQ5ymEjAz6UF5pbtzGjSVtqkHDClnHB3y5mDv/nNZVbqToC+Q+
6jHcL1K6CGLTtz/3CLh8uwdENTgseAgrLCU1g2klH2FpNmqRvyv9uJAHJ+FAGj8AdqJX5vSn8Z9a
sctJIBc+yycGfPzLPqFpOShl7xeodP7+L8HnCHibaDw6Oh6arG5YRUphERsQSyCvr/0+dysWGA5a
28OzI0HxfImAy6nIO1f09ufFCW+LPS7BXYitjlTrw/iIt1oEWXE/c1pwixEx2ag+EzO35l64Fr3u
jubIEQanjMizpoGtzibMrMh8qU450Y6mxbVx7uJq3AJEHSbhbNEDgUQpGtQE4jtpnjHRocMN7Gg+
IkISaUiufj8436nIGFjx1JW71i045muC5Z4nMm5eqgHw1M+m1lDyp0js/qzPZjX/SewO8DR0SVQv
6RrP1e5s+eNjg2g8HM2aVAc1WJnAk85esNfsz37l0wJN/bUjfUmpNTGazDucJGtKvncJa7V2fvaP
jJiTkLNMokW2xn62r2newtMGmLYgXE6jn6kv4pdHLKfizoZ01zDv1XeqPxhuYvdOK5ihWusQFxNE
CDdlFKrP5vhXMCmIiLI9sqvXyqY/i+ABvf9vXji0u/1PBPeXJJOv2yke/TNXcr4nCPo8t4Ta7M83
ioIXVXi1OAJETL9yBQ1err9saEaqujRrQV+skoKQf+MLwkycj5eFkec4mQjFgPvHo/g5RrtueWjn
E70WjUFxZMOBWNT4Hxs4HsXwL3T1q6om+MvDV5w+jUbh2fCWnaRATsBSwttgIUTJMp/HkOjYbNmZ
4fdo1LQ89Kg/FOcem+h+CH/9TJzcg3nOj3uxPSOFuoNhbIxxx9sSrmzDDSkJ6i4GTi26+3NDL2s1
uksvOptCaZU/HVwfe1M9/3yP2U1SI6JLPWGcxbXEA1oCJ5jOe/cXlFnTfOXN5FUA+GSoeS3tUrOW
uA8xr7GdErbkTgkWp9etoJdqwwpK09kxto2MZYdQn4vyjD9L+IPmHTo32KXXDWYcQYzrgu6Bmygj
gBkLgVi2a97XlpptYdiTRGNYoktQ/c9LyUk2kJpaXBTvxaPseAiwR3Ewr3dIAw/+YQqHlxfBDhsl
0q1KbKTgO7APOHMGi0qjzu9SU+EE0igtLDuHg499yYtz1HmsVflX+J6Ie1Eq0gRbRbGFGzL//bDm
fGPMZpsdnJiW7NcOEhD4p1v+vG+Z0j1UCsW4uCB/GA1eT3jgv7CR3hblCPQz1vKQwEeayOUpPMm9
SsWHkghZKo48aEsidhCPrVEpsHlK1qH3vlC+mtC/5Ra7+p77sosYIeYgmdtsJJup3kvZSI1BdobS
AGhiRCQxWrdYfcF5Pi5h0q6DurqZzAT/rcGe4pN2RXsQ+YZ0ic6GJv7SR09o/36+UYEasC25JXtr
Jy09oIkT8vB1zDOX+6LqpRDBz0rlLTewyzHjAcKnurI5HZpkmJU2xGvuqmo+PVU9qA70TexVazi6
Px1KvumoFT9yp93ClyKFiBtWGyLxJlMWkanDUJc7Ku2ezQjc5VVTa0Tg1oqCTYnJflBlGIlHt7Hh
GOuPc6deMPzsha+B/ggnj6ZifI4FrtMK9dHZmAU0oTufoAARcrOYHxmmn4NjXtMGbLnn1ScderOs
LFn4Os3z3jZjHWTd57oG/2xiCQWTJkQufJyB5WFAmdqPlh2Vuo9Z/CaX1ICzkeG/3ZRW1Wd6LKCG
cr/2Hi9JOmLqEMRPMXe+JYSAxLm2haz5J4QGmc5159AUBxZVwaQ/Y+vl46xicMWNy8QVX0YW/0Co
FiLThQoRiU3sF0qb6yRuwYmXtu69oe6PLeg9QmPPPdgsypcnfyJaGn7RtgLNIZJ9gXrFuPkCGn9m
/ARzURdkHvijvxNIO0Sp/uGZQNuoeAL3AgoMfTLZfQXsBAfvQ0JXuxxDGKAzSpvBdAIIa/9s5p2u
Gr4+kQg9d6h9VPwbEvDNBfS748QLcoCugsSqVRCewn/jdQXpDn1249Nl0YeYRVgTGInqO07p020v
V0ntBUtV/W/o+Xm5oTuc72u0zLpHqFv5F9uj8aspithch00EhS769bIJ9J2pk2P8N9T2nr7i4zrW
HNg8seK0BXHMlvjhGmNHSHbPFwaZGoZEiA5gIdCUlmEeYlmtLvli7R51Knvuz+qcJGUvqStZlJA/
7mrXf/7VA6WO613Ncm3UaOlK5ywPonAv+AEht2esURNU3Myr3o/CtCRSZ4zDW+hBONrGTGV+QJnV
VpSyRfTWo1HLmB+pshrAwdFkWRGBiWXsDv9Bq3D1hBzndWfbh6KAVCPP1jGTSjICniMfkfJWlgNl
O6e9l9Sng+uRcsiJb3sD0xdAUukf6qMrOc8t8bLTdwZezSj9/QiaYU6+h6jkDDIz85xcpcz0dJ2q
MCUfgoJLif04+S66sltbY8aWiWWEHfX1H/zYE0WyTESejrqgdRhRblQCze9OeEA5/xJKhq9KRmid
O87oI4wlTrncZOwksoK5FxoD9oK0Md0PnY7eoK9nSXqev8p9SJIQS+1AQOhGcdZDCld1iUAGpT2E
Bv/gPhbbOnQ7Hnh0uEx/ZRY3pH0u3lq3hiFza+g7kZNXOarefz4/Yx0nTimgcy/i8GuN440e6k9+
s90B5/KD9LXjhbVQ1o52bXQeO13xH8DVpPwsjKYDhfBLhm5w0sFpMYJByms8vqWmYB+YVGkDu+lR
xkqHzoDeZi0jwoBOZHqJGD8t7hTUG7aqLpGX+SkcWkcVvgy9ULfiU1cWDkl0ZCA/B80n6oSPTr8o
cfW640PyurA1wtauleXGupVKT+l7KSUVyLs4X0sPqhu0WX6oaY9JsnuPpMNqgIe5Jod85MaFhg2V
8+15KTZiMR57Ku51+Eubzc6ACTJb5kvX/FUYX0V/1W5AKN8ePHfL+dmWRs3AY+eJPIU7MxY3/2xk
5YYaF3V+vZe4tgVpsXWbXbN+j3Q4lcQvzSzO8XVFt5K0cCIeMNtBAlexiTIgtHsEmr6C/ubxfF84
YKNGz+MrpSNF2cWCi3PtUqBDuidrd79YslMb6V88sBuFSEn0u12o44qp1X2RH7gL4g3QELYWZzPk
l9Otv+OrMnnW1lEHN/Sizpsv9+omhkm8bkJzlQhaFKlN4/OKvrFGRF+kCcDLTGNks1iJjwJWcb0M
euNtwabEnaewcBGvQ66NVNmTw3BtZahT+FEgN7n4GzK6BNRNHytRnE3vwOaeebkQCZHs5fBEziPd
pifF+jUYPDKnNOUxrSydICcvpAoqUDGYqYuOXzevItxDAOBabKqpq1q9u7L0vTPE+0PGdHsnd/w9
nQNFQmjBgnrlx1RuQCEI5m4Yzm+DiK2zs5GNMEbfdKlQ1t6SWG6ZlMgrkpDMHIbSxThjLep4mYEJ
Ca077ehGcz7aOmg1H6W9KbV4Fgb5o3FGJ8LcV7v/6BSm4wwI1fgSQFCSxuYpEwJOD/Qbpt6HXeni
sS2VNyHyfVzBSkQ6FGNvEGlLaJBxA/qi0qrCXSL3JmfYdZbKgDeDXu37i0whpkTzOm7vaowLwbgO
VILKfTkRZ+4RWpvE7mx5/CMkzW1y1P07NWbTaUENU/0CetThaA6Q1KiXwzr11Hmfc0IxO5FDPeEm
ffy7SYezB1TRQFqCijEDk0dsiiQO4mfXiTFOPFmRB9WgrxU6MnvazwU6CD7SouIj/rYXFioYpKl8
q3YiK8R2BSpsjwqMdI+5u78ECan2Ut7b9qQxbzT/37UkRJ8tpVfCZ5fgEMOQNGrbkTn6R3BUo1RL
VrFwyX1YDMyQvyAu3gFUQO+EgG6y76JysUoKSVtZQDFrUh+AeA415j7aQ6vRGSmk719z/GefmDL7
Q8kKsTNikdrU2xaTM5eT2G1VRVL23LoQtrm+s7ygvdre6WOftB42dJ+DuwcwHhcUg2xBboLmfU1b
bW4GSXj1tjq3wf/DUMXFRnpwYgBzxIt85OcWYJwyZS7bapN17hclHBwmBVps6POkidJIQQPUl/N8
ErxUIuF8vaBq1FXzlGab1xkLywEg4feHmo+ee3crL0sqaIBF/x1I/J0yvIaLcHboICmEELSIF63h
nB05bQJZb8dqevRgdjC2Iw53WFBh2vpA0E49l2GxGfKAVxDpUSTckJMjyp3HUzOD9pOtqSVtqtk5
2Bo1/q0b4xAapgMCvOjzZBqCfYsVVaYetH/vDXH2EX/TDAlllH/kBSwRIhZbdjzsr5NZBAQhxUPP
LfmXF8JYI8MkYRo45ElX9FdL37PXjrVnPEw5qYADlkSbEQJKhkhQ+cJU3ZDmzX5LXPjdNSPY3rzP
2XxDT6+EOo/z2b37hXU/TxTQGlIm/1KpYh3k6o0KnyKlRmAUQBw0RnDaNovLZjT48s8ygvcQGv3Y
Vofoj/BvuuD32amsHAp88As/wOl57QMkxJYU+AxcUvMfvJI4TNzbHEGPJo3FCaHh7NF2hTXon2Dc
16TG5WRTh/hK0qmUCkMTskG2R83ck48TAW7b0myACtQQaAtLJLMVhQOMaJfXRaXPt7QjYWPRYPAO
6Z8oKBEx4h47aYGBgC0NrrNffK1gAHH/A4O6fwmacUXQyUam65rfd86AIJRY3Ln8WNWRCAfSie9D
P8gZdj63u6c9zZzjYCVqOcueSynqSgBrdLZDJW9FOqguRwwEdm4cN05+Uq9bDbpmTGOk5FlbkOax
wNlXRIqjMOR8pvawdmuxMBM7Dt1q0yMopyN7ScekkOQhLwHe89RM8aFbkaHZlIVPoLdZunzB8jQl
ObjH7lRyAoabYt8Bs/bmuifH5S0FMNLttBljlUr89aHLcNDAKzo0HvM9nUV1C3TJ0i9s/ukz/Glv
tCFgZviB0Ru6AQaMtWMxL7w8NY0wSTZ4y8PW7wbn6RtYrhAettIm71wPWsC9u28Vj4CQ7oh/7JWL
4/QKgwwlgEY39+N8szw+1Pn6CeqCrDhsx3NBotvM9cPQUefWCXXy62POVACkcKlLQSW49xz7lz8D
u/u/a2exhvZZIZ2lf0GAiNx1+DPkFKjOK6dvGZl2Zvd4pMDDjexsmS0vLXNCJZ/MnZYeijMUTOrg
lEZrMBw6N8+KrDsGaL4TuFZB9nqgqsBJ4Xxtk/b41jOw5Ba40Zm0VJZ2jUdCtfoa6tQyQbDXsxZZ
EcitYFt/AxrwzAGYP83fsQ1S2w1y8jkfKICRn9H5ydIkXaxhIWAzc91pD526h9gZdEOHqkx51ROd
FYyT4sIehA5hXHGvYFNX+7wYtZQHQ+fOgyPG+hDct4pw76fdPO1dqSSrQws4vojfYR19/H27GmnA
K7dfYDy0xeMVrssj/NriqhQESgb0f3DbhhgvdLd2/ngYIM7CtJU8G4or3hC50gkYTK9LxbitlB18
eSHDRtvePbh0qs/abeEnENU0Bd++cTmUv8FkmmQNzO1LYsfZ9ocn2Xno1h/Uc8vM5dtOYpdN7fGr
0odRb2vbY8TEwBsV9o2YP08ocYTlUnNspDN+IAxe6ifCk3N/QtX21iwRPp7YM/aJU8KCf0gIR6/g
mF1xWJEONSDICcKKT1NwIdolLEWLjs4iOaNG+eXU8XN2doKmal9Dlfhiwh7tTMvGx2aS3x4I1nWd
o0ceFsEbSbo3/OPe5jhYEvXDhIQT1N1KWiiaXZQ3GGiRUW1HH3AUwAtv98KLxyXFMw4X98vOsCYC
BJtL4lzJhTVaSIuKAqrsW6X5IeFEbbcjrO7aWB/vQMJms3nkfElG0NJJ2D1uBvUa3jErHuJQ7IPl
SO3Kj3QvoWYQL/RoIHsHA9GaXPAYlHo2BLzjf2bXAI87plE7AHYAjoO+h8hU/ha5pJbPYh+jxpwJ
Mn8Owkb6PLVj3BVJOzfazxZRTWy0y6om9TKTsMGHY3eZX2Tt/wRiJBE81thM7DSUjJ2v6xH7FODx
X0ghMzG+2V2ZI9fKx1y7aLgE2Tfl5iv3OsA1LPZD5VmBJH1fhzYgq4dEkvszX8avE6+jHDw8Kk0D
2cYUsia5VfZMGu8LiknuK5GCCxdqD002NsC23nV0dw7VRLCr9UP5YG/UiNOOg1XXPqhHTngF/J4A
fNbLNa/3ll9aDzrz5VbgF+jOjaENXrUZgXL3AP6bBKTCyke/IEeg0G8bzDyca9XP3GPk/9bKKzSu
1e98RvqBQy9w9meKXNCiM9dHYz7TRIutQ2kbO1Xs4i7YBIo8gTPS938qT6yXr6YZSrjis8aUaxUd
GvaZWpm1Zqj8I95KRHFfTrqZ9tmz5LRVprL4VoEu+P25qjE2Z9Fk+nzSZN5AwDg3rVBpryMmJtKA
OrvCwC/HSh5ywx0e9gi0zLMcqMfTH/IlhXh9eSzGlv9lbOWCn47ff2jw7n6803ZVGeEcam19rmLa
9jaX00hDZAHtkyJ6bzbYkSRAqQ3MtWsPVxCcTbKDJ9XMxarEvZVrabwIFt+3FzR9zEJ0aTnLNDAz
CSkm7Xnzvn9QyudmvJt/PXfgxMVlOTniVtbX8C3vZ4eSveIR2EYTsbsNOfOs+XE6q8x4GJo=
`protect end_protected

