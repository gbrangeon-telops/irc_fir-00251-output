

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YeJs3h9nPnCnr3aRxIBZUXmhDS7WeTgKjgxxU15evXAwgLO5UoYuCJb2fGld8H5MyDQGWc8UFp3Q
QS1bcwQeLw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QMDnsLueMbfhPqb347LcBnHgrgkl6fbZ0QORe+igLd+Fn4pMYglXhNwzAsr45PWnZnHEuCtMe3Am
9p5sJ/ms8icpsPjNhMihj0/+LhkVUeJEYGJR6AGOi4DauCIoKWFsirWy53ZScEPa2MEe+a32HUq7
sCpglfzmrbsWEab4EEg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F3FpAl1oCeVkGEm2PKCJ71S6Z3CGasBF9SuzLFWQnXwmvUuKd7HyekhOce1QfyX+pLQcgfmP3XmZ
qpZIDWOrbZbtPCk3pZcRYdM0rjk3gWPTq89GN09GyodyzYH5nERal74RXFzqDSlXYzgzDvsSzAku
WQ8fc8R6wi9d8ZzaPtv7Mn3RMOg32FvlzTpy40zwgHFS17RZjspNh23gqb62COtY3bIw5wgzOnnc
pwYSu+4rxmNM105eSJdh2TJiSEN9+pTEYMITQ2PUZ0OLL5Qstj3GHFD8/78u9ynXfzh4PnzFHX+c
DtImYoh20HOPJeCFpBeWPHfekXHEPhbC52n0dQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lq9ua7Pc8cPhzNKkRvioUx2DGTzaswIzLnIP4rJJ3cLZM5wsk5kiUTKl9rdBpb7G3yE/zCnmkGDT
ZEvIhQ4CGdpOb9ZjoYg0BIc1GhYnGIexWpvkFarqP15NwctZCibdBpj579M1D8fvQ9Xw1j6ILLQ5
gUYJd4OzxaJCHTNx0vw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qzr81pSyvLThhRepJmzjPLJdFa8x8hA7KFKfUSPL+CaCFf8sC6XyXYts+1DRzPvdthUp8ISKrFAv
jy1EBIdnZB3D8J/YmjzA1s/E0S3V/3tyfjjyCDrQgRkpjqKN1zwlXCzBMyGSBWpl8ENwa6XmbY6s
fYy2IxFIrKpit7mWPaxU1OjywKhHRwk63dw93KzE2hJmtDZhJmXSPJNkgusdN/mkZzbIYUj8bMZ1
mRTDgqzRIp9L2zyHSB7GfUn9cIiKtJb71ztIZtRMoFGfKpLMWPUiRhyoCIz55vgxKfE+F3ghCh2A
ig+nnH/YWVIR6bKztafV39mEL7utiMvwk79iag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8592)
`protect data_block
YwcMlqAQ4vUKmq0OJgR+VBWc8S2nRP1LQ1Sgi3K8wGQDu8NI5Xj2LXUbt/txLuifuMeCpL9rQRrQ
XKxR0woekhjTxXi/Vu3oJdMSQQlOf/fVht6y4cbwuG7izTdgN+bN9C0uxLV6Mdk2YxtXZ7A0+DxJ
f06IlaQ19ynPgmPdyf+9VC6wNyhr7N1aA3jCXOBkAATsNmH0BPsq5K1tmS7RvVkXU0HUJJi5NO9O
9CVQFzyP8dfz09qYLvlIlIsukvZQehPk8U7x25dt1pHRLihaW92VFGDE8B04g4v4tsXjBXBeFrAE
7qQYByda87As5XK29mJE5tIXges4Te1/p7pR38/ioM6+C28TUBNaWofi+pV/FMbwxogAMFFJr4R+
NivwDt6zN1Pvy5VypZTIUQcmMdaKAuvSG0aUAn/RurrYhPapp4qSXH6gS37j4OKGALjS9Hs0zT9Y
0QKXrVJeNc3AnC1PemQcVt+Yul8wYHGAMMs2PKZBvLJgjqaG7D2AEsFQctyMqH5Kzo1/qEWBxKcd
xUI8H55nTr7Qn3Q1HKrrHlaE9HPcfqtEqGD0wpghUye3mhhUSpKE03UlhnB3iG4Xth+G7hvEdSMF
bJL/zwN4KvUJinhuUttk2eEADVSsicc1uSrPiYM7rKx3J+oTdFnFYxyGn+uo6FjrOTMU70azZMYE
hLLP/N/x/+UDnKaKRGebUY3XbnLUQynGtDyCzQXy7K83Os78azi3Riq4jPyOQYgUJryOD9Nhdap/
5pbMrswwreVfucz++hL7KrAMiTHcWUllg+bgIm0SREGKn4Lw/dIgYvh4ftWmH2V0ol9IVsPS6wa+
AQb7IOiu1fuRzGb4O9+UZAwYMUbqx/6b9YYHLSg4CmkjLjksZuyV1SMWfrR6Z4OIui64ZnE63SRw
RI3kL52BGysEzMBYucLqo5E8zTmHucT3LmkVpybUZvlaEwnlwH35wCmglLTHq2jrzyxgeleij6EG
PuRnx6viZbdDGHlYE0756VkVyuYyEwNQX/SbuDvUdvDxOxF0HgwohgSdyTP9Clj1Cuo7WPIpck37
BBJVdZEpxi02KL+alJwIH/BInpkYxGKMaa3QQ4P+zFuXHEifvkz5aQAEhNDLW/Bhwrbd6q5iRl/h
bQH0HM1Hh5Gs1kPqFuazLGKYUHp5SLTyQ2OE+pc0zBUB8NPIJYkW4c+x49te+4mgSrMNoWj45125
6UqA5Xb134/pFPf0eehzG6LNqh98Hr5RUTBi+iUxBNiJc8MPW6ulvVAFwQjMvN+TrHpma+I4mUPh
eDilxbAeM6LV3LlKGLPft2ULm3PkcHMRZWVNglZ1SRhUFq3EAKE+ejjVdPeFlvTSk+GnrrM3Tmkn
TcEBE+l70UUs1BnJuQxdLrbXcCPA6iul0b7f3VVI8rHwAnIrUwXh8OorKvq4TqZKTXQmIqCDKKCL
DF5qhTJG/NL78g/mraINerkfmkCpjMG79B+M/Mx9wrj+PQXtLNQUbE8x47xdVHeRZNdE4SAXX2L8
JKfd0EmnofQfnkT2L+hgr9ROjl9tUe6fgCIOfpgFG7CjVnS5JtpptCRSObDSSeOjp+F2FsIX3jh4
phNVVE0kNmvg3JdFipLsoCOADppdDqxG+xfC2ER1greblZJBcVw2eYgsaniAIGIXJrIezK8Numiz
E8NMB9kIhCclTIev4CNRcPAT1ltZQXmphm3bBGXZ38mVWqm0kyvGve4vtUeOJAEFDBtvwOBmjBSz
3sJ7+MMYla0LmGPkzLIVUg7ngZv6j6qp0vhmnkyGlkx8UmwsQzDENzxcbF9i9SXAxphDh//1pctL
C9wWNuurl4xLJlpwh5G5hwM+krXjj61m8qX0g+VMcXqo0JGoo8MfUXp4LiydFX0LUJodL3AguoBg
5m3cNpTZueb6WtosNVAzZPYc+uNHNV2gzZvgzKLQNsLJkqyZQBToj4nfboonohGrlZBDbdfky6yQ
hIm67J9ynw8oO/LV7m6egmyeqyx/3ltDlD3esnAC9TO3R6RRuhE7RrhJE4FpPfdYY/1gNvzeIH1N
iXIV2VIgcYTeIwv4ncC4/xMdhP9mVEVFthvghBx6RXDggNH5XhWwhTDSbH68WqvZZbftxKErUIvQ
bXSiOoHq7uu1KafV7r+xw5kLsSSYbqqp1OhuvLG3dXXmT0vWMEZTjjxl7seDWsq+2teOm3juP/bx
r/3OL+S2SV2iOg102q3H7qhU08Z7qTM3yDZSyOOFxYUVdQbmiz2WIa9CU85tqmk1t9cwdSUczSJy
jQPBS6Rwzld1O3bGJgbHzAmtFdGU2vCqWUkamJG63nkKmRCiOxB6mMJbZO02Oh2krY6XaUgSl1g6
u1rdXVkXWqZjcFgZo6TFtm1dSY09almaiI2WMD9vDA9WnwF/qeDfMT5Gk7KRfSglCoCorRSE6zuH
nhOQ8TI4S7mNDxI+Bnqp+btV3PIzBIAlOYeuD1cANXuuBkHkFPcHDcmGLo/yjTN7rE4Ft33k+NbJ
hGM5whhEGbpyQwyuf1xsuR75Xpw8b1SwJwDSFTvRQAxs3Lmag4QrbKu4MDxjUr7lEr8dabYiSgZ7
94C4GQS0LAvRW7T5H8F+7ja99hlzR64ea+Ea+zxNrcsMTnqNeGhHyUWgNZvUXUfv1/0lNfxAnXWS
3XP1hPMhpxVNyU7Z8D9ypspRQbaPVk+IdRfEGxVY7W2/3frcfhBHG2R/Zejgvd8dxzRTVEvSh2+8
KWcgB1I1dOc1n3GETSDBFp9iilWoaKn5uURMH0vdYVG4saEW9E+C40IteMrdOx5vdt7vBr3hTgK9
8K0rcZeiCwu2BUlzkRRD3LpockfIE5PVwlfMhQXXTQu5CffXFY5VHaue2R0EL7bnG7THlHAGjPJX
D76FRiDV133bXxan1nCIZ5Ldr+8hS+Ah4Qus5Nbd2o3IUFWb61/WHHLEzn+C5Jqlt11Hn9iZQ+2x
rdz/zDQjxOZSB8w26G069ddFQUn7zZuyU51NBFPg8EOnDtG4F+DohsX/vQsJkO25MVg/+dcUTgqm
t5O6z+Kd4YiBWJfYZIydHt/L2LdD1wFswbdn/cyl2k6joUUZEniqdIA1f9OD7PsdkMMZ4a0+qVGe
B6b69EPHZOv6kgvpgdlQl1lvyNC+GQ2LMqk2v+QbrSZT9q18hUAZUk0uS5uGCv+KvBlenTE4vavg
rz2TVHR6BZphGTiIcN785NrmpwN3/xnQYJN7U4jOebIIMboZ/FvJ+vPeLBOYxomTzfxAEWCGYrGq
3DlSJHKCJilBLiysNrKJW+oaaM3V27aeAZptzneG1kgb9eWQhbvQLizEYPaoC6SIg78LGbR7pxkK
gzyBqSPvDL+r97HYhbZ8jPKvAl5/ZCB8zjsP7cFTlJWg6dP3mF7KiKaHI+Nkvv4D66je6MC4csUM
d8u6EOQaQNO+TYzMPLb2BDoUHjsFiB9v4cko2PqPlFr2EUaRfrefI526wbsTnb2FVzwXHX5Yj6Fx
PbtcFxYCQCJl6Rb/GXlh8OaznVGasy8SfsbHEZ9w5FjBgJtNMjx/MmqFznjuV1fwkncxYf5JqPak
9tWueAt2P7qR414l8mX2+ahEfR3Bc0Jn53Mxn4dIfDcOSXZNcx5Oq8rOHbqy6WIeIq3kcdrAmYFF
xgjFf9ak9gVzKPgBHhldoZ1MYcExhiLDI12Pa8kXfEDzEVRR5/ExreugSswfhUv6+4BMC4GIcFSk
Y+GJZHRIM8OhVus5fwO9G7R38F7r6gYe1GtFnReU2LJesImsKtElTQVUNiUx6IwLuEV4APlnmxC8
76aEv6O3qsEEqjGppnmu7cZLNUvEmCMZn1GJ7TD4wKqNOZJFzDZaY/cu5Hw2jop88ABElDXEZjMT
xLgs9ySMQznI9bOcb9YSUWGXmb1nsoYqVOJsGl+fDOL5BZDxX6HhIy68el3NzbRM9TbZleKPUpUw
mEE2LuvWx8Zcsdzqo2Ul2rO1dwWcwm1woxdER4uH4RZDD6H0VtiOa1cYzVxYD1N7Wcl6Tc+BFlEe
PqVv6FOQgrPRzDb1ENEGHGbVyiRY75+UvFpfIxOil7qhxe1d0H1XnDCB6ZEPSkr66Sv84Bb24g3A
AkhL4XFCzFtKmpSDGoUxI0GSuNoMlp8A20KsXyv++cn23FGY5NJ7lORjye9BS58bC/itGg48NpTh
grkFVJWr61wKiUJju27/CgTA3RV7ORk78KD+B2wwEM70FD8REDeegEZkESJk9pAqaBZmCyDX5Jva
5MSWJ4ZFLv/d0ZspIhgWpnO1HLc1btHoj4K+NnCHD2PL2g6CYRpsmZyIxbq5m+pDEjnm/T7ryEaL
Ndvhsj0gR6miyKZcahrpnv232KyC3jGO7oF0y3/s5zL1MsmZ8Gbt56w4XQrrYt6GFNcKIPWIEzA3
Qp7VPyB4O1oGpWuC443oh07QkF1zD48nDqoJbWxngAdGFcX+gNVXTInPh3VmPxgUdIN5zWnes7Fl
OzByWO3tFEujlhJU1LSAL+fpPbCJKgVL3cFD6QBWa/YI7F+vMGMlzEYO5t2L3nbVIHpSBp76VL2W
iQxfy+BtaKcHXNL1ja2twZI4wevuwS1Fswt2iqFl+um/qBV1hAAHlGWQ25xXr27NVLC23+DzSjfI
9pYy4Dxr5pnjX1zy9AEpetor0P+4LFj1O3bS0fi6oOkUgljh2npTLU+3dPIApIVEed7hhpGdN+sQ
LkYlg+ZFsg5UAhIbLmFpGuO7SY4rqrnQuu9dlghh4A24gdZeeGWTZUp5TYKsNpqpBz5k5Wcsbsnm
ReiH3tJFJCS41RhTJ0EDC6VqUely+ybjo5SyOzFcdZa8xh5mjicxXohrDjyEP6x7lfcMqJ+wWiqN
wzZOK8BQGLV9W5EKBLpjt1ip8cw+cOABV0YJi4g+HPwzy4IV006/v21QjYoRjh2oG1ThKBh1pZBB
vhgJJYxF2NLfVEaG5i3PQGBtMLLaLCZ4cKj/D5ebo3y7wi2XlxCe7jE4t8fiaQBemUtjWvxAP7Ny
vJ/zANIcYFcbI3ICwB5bxTI0v6hCP3syrPrPWqz3koUmUYhIpu080Z6pBRpT/bjrWqbdnhFxruVj
IWZKlOfw0zr5ZNrirH8Zo3+/YFIIvMQwZlMh+SiTYp4DsDZjTCR1rStE7j0HYhJu1RzN4XP424EZ
7JCvbplQ/zcjs38QLrPqwVmWrz+CUMekUD2R4jVnf32tH61OvepJa333VLHG3Xm/IPUkY7xFA/IL
gBU8MmykRa1kSEZuz+XjRn8nzOrW89rDZaNhVvpsRMSJDuCRIUqzs9LF+VDE07VSGy33gqSyY9Dk
KRQ0bBk9tNpMu1w5mBwHLn3yr426cxTGHVhEWydEPUjzGnYLaFiXJB6KIMoctKxUksNJ9ip1C13a
q13KpFPQP4ut3aV5wQ9ZjCNy7SpzylKLciGhFCfzCdnsqC38oIY+8VLkuGoiF5ionG7b61QqZMGN
mVMndmXAJi5u+WXaLIj9F8QNNABQemo7hsNYus5yYC5IdEC8mFtfiorZDb/b4SevPKnDgB4ymTQI
VIkPbGmvHJN2Z0C3PHfjS1vKmJrBUIDH1YSPdOFwqgh9oOuXJaWIjiZvQKaOia78cQs64WUZnrbK
KZVGY3bHrobkQg8/IyEYWFVAlB8gUwXpT7fIgumFwnr94PJxpviIJyo191kiYQpKzGNLq/aEsW78
Cfn+QiDh9i1YR03QPe90A/MIT3VIaS2BluWfOmehtt3pMmQxh57BH0RWfv8hqioMMCWmzqxpXxIT
tynmsye9YB+klRhy+tKBz6kqlVHVbMbj+wIJ1gCs7g2t+CzCXA1IULkNmKQlqv/MX5urMe94VaVV
Bf6ya0UzG0t13CNs/mCHU3l84GVGXo5e85Gd7dBjgzBAmP7QWz2zXHqBB+68mcPow8A2FN7Lunyd
NsJ8CWnewCkG+o4te5xU6Bf0ZllRRvtduioRwyMLpk+zBfAI+6h3MvEtgk7GuyVDDPRvVgFEG6JG
UaQsxWYUDjU2pYUjUA0e2n+QwoA2YsE9cZuRJRWubFFkyke6jE+cm/DnUqhXEs70ukYXiotZH5qm
D5J36CermYmX8aOrtEZ8z6kv027lDsB5+lT3TpGawZvarNvhQdfNRILPU8fqP2DLUy8vAcyBdTgW
l5f44HUR53dAqXErrhod72dsnD5mee0/LAH6gz53IQFb70vIXkF7EGdL4LQdo3Fsc3pxr5Xg3jqS
XTGoIAcgLOCy+DOQcF/GVGi3XFVgs+kCnxyQ3cZxBXT6ocFnTQi7CfkU0jWzxqpzZYt6Emn0Hotx
8ylhwUdn80oNQYImD/2x8Co115Ka+6J+ZUSEJh7peAuT7hY6lljjuR5O0ZWdp2WQvj+8B1HNHvyL
msbOYxm2vDWnN+JQs8Z8Ajtjxjit6AI/Bms5aekGx4dNAB3jisWgZKkcIpbwn1iSyYSvGXPN2Tz8
7w0ZNw8ZHTrFCXFArZppN2F6cw5Rps7o2oRcQkATJYS/h5Xvyb2mfd27yNu+JY7V+BSM4bJTUYmd
+lEjpB15SztgVvGAcp9oXwaQRz5sdjCoNSuOagMpLKkWtJCOXwdKpZMQOrWurHbHF8ZL9QSAiCWA
slp1kcOabVxFYvL83UDTESc6wGeVm8MEPvHKk0Vq3uIbYohFo/vEOAo5EFUYmE0Gl7Sg7FC9YQ09
CvGfDthGYluXa+O6dDFE8bAt8yYFhv0o5qb9ZPXm5+2qOUIsneoLyMlM5n9agKjlWGl5Wn1z96j+
+OQ89Z32RQHu1be/GrVJt6CNf9yw2ETGjME5Z08+HAJa4zIoAvkt84B5J3ZFZEpE/YpuZpcdwHSX
G+Wh0PMQkWGg2dnH9VaMNzik0RJC2PW09rPcXd/iTW7elyPUtfDjhWmtmJcHuog7jF+LGpJ1sc61
DkXzvwNPZ6GIYI40nMcf7Cx6HrYx2IyM1PY5z3EdA4oAewFhm0AHKbFIZWUrvHD/s8Iav8qU7LLq
HLEbOJtz6v9DgXgKUGV+/LixOssFvKl0bJ8S+A1Oh6yHSppUrh8bkoDCgcBz4SkudKthn9Fx+rhy
LzVMuCo6LXZM8OjjdPBjZXHtTcOJixuZdG8fdjW1Ks3+AJ2VctHQmq2wNXvUiCkLVnghC3KDBTv4
ESpvU8lBsyOzKIF2sfuWSKdTqdXWoI8viJwKP7E9tKcQP7jMWtV0uh92KuvWk/NSqxCGhth79HLD
ezTSQbJjhh/i4ZLUnv8T/N4J9QuqzaKScwSKC3OviDMJ8g0RMP0jQ9YHiIWnbtkUZPHsIqI4VFpl
+efSwq2PcKpO4P4uJ8PZiAY2dC+/+glGoeUz/fgPlfZ42ELqGv+MLdHypF0hws4CDmZ0E8saPKNI
jgXQcLu74OUXbRUBNE5sQ73i6k+7tup3O/UsWct0Crc7ZUhL1zpUcHfXNk///ixQnV/nvT/BRmtf
j+JbB1c88npNsFLjjZxH1egVazNSzQgCkpmmkJKFmaLBYaTq68CxrMEcpaxbrZBeEnb8oDU+Zb1s
kCuK/pnxMufNWS8f9JIKnH7OJECrhwT6FYZ5HSQ/RNb0RJUJoa+Muw+rcEDcUA9eh3sQRSRNowOb
zBBG6/41mB4SpFx4r3oK4Oy0zr+koLMDCXAmQMnHh/06BsWwhVHotwmhxyCVfvZ1AJMNUSD/pe6Y
glwnJGzqC4GFcHfjKq3bxcADG0lSlVNFYmACIurIzh/wyFBXiagahlQwGVMfoZCQ8/17dFbFffud
dvgX2n/2FoioP1QpAGVp75JU1U9VECga1ES52BtuTb0DcNypJoIJJj1fXkwHI7flifR/9d/TtcvO
Z6pre0wAO7+iOvk3Ik0hG767sOLxa8MHxFYcqIPl5nyTOavoXCevNMXezkDB3rWQrjaEAL76SNeU
acTkTiJ9MABV/MMRsSkp87XutPHaiRv3pTw8H3SnhxKmX11UNUey6IW5shx5K0ejxMlF6YRnZo+t
yv77Y7P50Egr4szyyPCo3L049x7XVr0uWBz46zHf9ExlQJ79L/dLGWnn7abr7obxBk2HrCnnQgPQ
Gr3BEVoIx8Y1fTLTJO3H/J+BKAFy1cvacB9KbN2/REFuOsuGkT8Mp0U6UbRTJ3jnVpOYh/cgatWU
nQmAeLXfNP/nf+oK3bcoIhcz6wHQwftzWhDBSoxAsYcpICsB26UN0DFrwSKDwIu3YvqDrZjbHzVV
JbDJjsqntgn3/7+6qXJf9oq/2j0BDe7sYTnm14ECrAmqYWyW12T+XG9UZ02xWd6UBctauw7kcgIl
h5MKvRjeikx5XedkKC3ovWcHRIxp6L6mhOfq32Tn0k4ltf1DHmuMJGAXOgh00MoRTWZgouUYtoSk
UkxUck+dId5P56lm3RoY+91ZcBthLXJVAj+Z9U5tS02CmDkCyHaAUTgo6tNkNOevgyfVLID3TdUX
NCnDbM+h55t7rESa9ESRGnQ3aJhGBaV30XTnMDx5In93zXkHxX3neHTTCqkr2GK7wTdI/T20Vp4m
Ojs0UZH9mMNGG6YcxMQ8VMBLftBcY6HQ+g0GBUNlm9FRjXd8wY7IoOMvQrhrfA1bkPyS/nPKAk2/
9U/zIAB/yGzR/B1efHWhLTSvIs+CxRoLNrgzlSCYWRhmxKMqrqpgYCm+AaSPmq1T/0ZIwZeEFnma
r8/XwZTFgrQoPd6EufT8zJk0CA+iLlzpzYyiqrVNgIY2tAO2lpI5xk09bF9KHJXLH0JgNsHlKu1o
Ka9XIHCBNzMCaZreBitrsWzWK764P4RtpHTwIKS3cDD2nhfB78e8TQBuPX79E8XNJmwcYWD29OLJ
IcQqq46VXLjB4UDdwg6eiTYXFVlmmMaTs3bPIIvb0YLdPOkr2btBQb2o2nF90YsnLQvrBUb1YSxT
0bx44oisOKkCiRCpPKX8VWn86wkaO4oDJUtchFs+8DcBT+JR7EgOlYXvQkPO+7ktbgcCd6D8k2Kx
FiHUObrnfJibILrP2XLQpPj/gvLSizANT6zFkv/vUtuhMwt7GCZAta7lcaPJblQ38WSPy9NdLTtm
KPVeWMxUx/l0DwQbPbTvYMI/1ZvfLS3Cndj5fVONEatznrxP6EPNhRMmnZ7nVDDvijwW6WTRC7xD
jfT38R/InPpVQ2Z50OMO093xZcdyxmQGNsv1d/uu0WKaEm+HF/nwJJzliDrWK6L33Jyrs/ACyLgC
/RSocr+yHIthQIezBEUJe+cpuOJTSd0e1bFYtDvwIO2r0Z3yIXQhqsif0mZnrcJiAGlgoRZtYVu7
UmXw7nn/pnQMmn3FN/StO0oM8pFJURHNTwsBDTTJ/8e0rTILtWwpxS5/NIPQt3HgRPFNg1v/0U/n
SNXD4G8fmcCOlGi0esUAXrG8KrDp/eiW7G+vlFPjMxFfqakmmefbBbbyVdC0wjCjteB3oOXcFOXu
KED0bJ8d4TPovaW2ltEXG0jTXW6JEZBcrBgCsu+tO6OikiKlb1J5VJWsFfSJXbQccYyXzsU1vhIu
8TRDbptKQ3k2annuAGNIevhiGYoBNr/QzMUHNs1nO2F5vd0+/+5u/3SEDOCOpbXbb3pP5AgVnPSC
Tf06gTUNXplPeW6lk3eUUxDGE2Bbo726TAN1afCCxP7KK14tgM+nkWo4f+ff0g0X+dAaGUm+Jx3Z
fsPwYh/fF7Kim6folifvKLcEVpzuHm+FlicBmuzGrA/w0jc2t1G/eZM0uc020I48y1BUNXA2D80O
eyF1wUNGLbto3HqveXqLlVxGGPhs6T7i/76cy4fZ2HJJ005rBylVVv+rcMEqEdXMW6VlpG6EbTra
BDbZRxkVPfZc1LqUVE4Nr4fXMxgkO7SyJup4pvy8qSMhoqJBJpidoXKnZ5Y66MVfj7QuDE+fq1Hv
ymN9uNTK9hgc6m13NlcYVMVIn24VsQIKdIu2T2f4730AGD7JlM2302xDiKne4zucTNrvRbfseXgy
mmTXWdsoFJn81bEOoyskSPREoQJe8t1LkTmASKr6DBO9lXOVR+/bankVzQLj8D4rSxEb3tSW25m/
a433VPOosa5rgqZVIZpWQde7u1vYQa3T487vPC1T+wyELiC05tlXkU/53hUSafp7ZzRGEDm9GAxX
Py61ajdA7F+SQUBB42qhW484Q4qUT271GkV+7B0y5aLd573KDDl3ux3cP1c0DL4piPXcepGj52YK
55r/QUDA9J6baU5syGWNg+LvoPX82vwDNgtaVOZNbhnb+uc9FUiunF+dk001UvKsxoa9N65ckc0J
VZjNQCF1+dYQJ9RAJUyJrvz5dYMj6Nxpa+rIctNzicqp4UQQsddRD3fy9ABhHXb3ulLKOJmx3HB2
gxYr1Iec6V/mexzyr2Opzysvd/Fz+gwos2J2CIks39Rq8GyPHt3CYOvUUeHYLc35tEW9WiJzEA1a
WdHoUZUffn8y+UxTs/Ma3qf3yuxCiWKkUjMXUhHlOWRvjaYmbUB1mlsSSFZuvj3jQ6u3JuxXtysL
TYVyRMa1OE4zfzoA+P6Y6QmGNf0G3GobdY37bKJfz+Q5yoFcKn6NbtII1kz8w2lFJO1yGtXAbjVu
qX0JmJlrTQ2Y8T2MKlaRRvMQzCNsLITfN5MxmRiwOVq5Z229LiXqklPAuOxNXaomv5hMVJ6JH8Bo
JDjO7sUyhrcrsYf/c+e04YJftCOnA3VTYCiVS9ZYmJ8mtSmu40SS7eFwc+xzVvuX2/TDxnGh8eKH
FmfDGfTt/YuegGS+l5cS+OQKJhvkHYQD8AMV9bEfvgat3zf7RxKMRyJ5pfPEcfnUi/5rl/IyKFHB
7qWqAy6lczDhK4yWmuDNyakS7hp5t+2TVEOX+g2UGlkn/3Mj4cvlqQ+ZNfkTQt2dg+H2YlqrEK4j
8w0Jookuk7VgtrwvVt5CrJwzAAx0eZgTAgZl/pGKEl0779eESSbNf3Zt0FBdQ8MmkQDTqQwLTAzU
dFEEAid1i9neyitJu8E8/dVNmvKBaJbFm0qwvJObJ/7rooYBPZPl531v5uoOzAHvppkDTJBgV57R
HSfX1w8ePvW3ft/IRnD2fLwHKavPby77w+93roqLJHglUkg1U+HoMTQzsYHaDfbj4aTxzTh77kGL
6fsDFg4F/rp/d4SXmeVUcFPYQDPZZNmaXy/f8U5XY5U/9eGEimsAUtZ64LVBPtLLz7Jt3yimbXw1
sKvtxvDin36Ta/6ti2TtQClrldt42qHZoW377rsJU+Lu5roJXp0dXpmsKnOt2lsiAlWgFmvXClWD
VoIyGEbbs62y2qmCNFs8bcoy6KPuHntrtI/P3eDQOrufzhaM06mb8Z5aJh2azIeeaTAYK21GlmDg
zEW+Lk/GPytm62iOd0HhM+WSPIHcgC2oZ6cJDoJS7fqVEcLiTrUNcxVxWqwnvjtYWF2+QQthWZtq
RPaHNhoXgzEatCM+dUcoXJalev8TiyhVw7SKWxyRaNAt+vHuBKStCLYt
`protect end_protected

