

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gqDFw5NFAM6CTSTQpb6ewV0dkTDze+wC3QoGAxwxbjcNW9/DsOht+2F009+7g6jE2OnhGLtqTq+c
HspFg2GBAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OROCzcjj1wgCYlIqlabkGZopoXwccuhDPoDiFwbBlsbzl7flKX8tC5m+07o0XejIs9tQT70vCTz8
eor9UB573WqZyEwu6nS7RfReZTn9rXIEfFTmb5LNQYR53WQufFJWXVGGzbi12Azu0TUMNBykYjra
GCJvYkOLjulS+N02/QU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y306+4wGPVAAsHa7Tcr0Z+Y/dNy6G34dYeGbx7ATqkdiT3xoZwFMriTbyxCB/BNDpEEpWtR2x6B5
1geIXl7xRsYW2a/OzYZ1VgC14cIMMrlyvjd+Q0oeBhNwIf7zzOU0YeLe10Ln0VhNNlM9hG1yxJpm
PklN0o7dbe4z3qSMhzdrqG9CNO1AfE0zEYRDe4xK7ci9EcGBPeIBnjhSSGUwaUeKV6BzeVeTBH5k
pFfAdDfvgi3P1VwvurSSAL/VyrhWR7M2OhP7fekXRqEU99K00pFciI0NAEcJPUl8pbYtjc86ccu3
OmuQ0fZKcUeaRlPX6glqeiiehMLm/EPWzCdMgg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gSn/ibMO73s4UyV+DQBAOvPjnov0A3ONpbzDn5S1gDHbJc8laliw/uAOvABs0KKAN8Q7GKr5UYxh
qWYO6FhJPBG8V6RCU+sAaoeSnleJb/buC83HgJws4chUKE1EbA08UnkA2E57wCSfAlSkdEQl5xrl
E4NsCY7zrBmnjMH1Xu4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lI1FhNfWvnI088CMtuEIyHMeXPGNhtlppeaUXaQvRzrpC6F1bRvO696fznybaYq7K8VPJB0YyXVb
8oCJzTtV2jMI6KoF+McAzbvubpz0ru0XOCjjvcTsZJ3kGxHGUlKh6xdlB0Gez6kASJJe4GeTuEaI
VZNg+Q6ea8OLPKgQf7VICmBv1vM4svyVLDI/pSGiGOmfSMrfWDP60zo6tHpkaDS7uHEj2WN7lXT+
Q8c1SGnQvLeKyHV/kGG66fpNSvILAslBR0l5Xt1/csaBtahK2IV70dxaZkLZ2c3pylf+SxXTt7v2
CzVvxEgWwmwKjiuhBgmVM6qeL7+tokO6P+FlQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41056)
`protect data_block
Z9/k7vw0KfheuYlCQeXLeX7Uqft26wnR7ul5XRP/MZ1e0uN4ZsgEQKjx6WfbBTBffFQVIQMn1cqV
TZ/D0f9XwgrHLcPa9zxtgp//ZNOJTNkzAcGPXfR8yP9YsK6NurWEmSDty/b19hWIFZxpMaRSV7TL
/BWbGo/RLzFKs5Z9v82/iRCA0PDa5whvgfQf5nrdAp6MecNDd2OZC+kr7ilNUpuWBlAQmKDNW4VY
uGhEgspSjhsKtBgZVcgjkzYFg47CAy9RBE34wPQkCRbzdSGK7LYHMIyr8ujC8hsCUuVWUtFHGHYw
714k7oEORrN/76pOWja/Ibui3pV0sEdHeWNHE0rxZH+jblIFguhD0CX6wEZoLnlUMVreDWj9vItE
VdBd8VDMjV/SnMJ51BMsOiSoyl/9X/Y6yKU8J6lYZtaZtd4vGNlyfiUA6EZD99922wRYfPBJXkGO
K3Is3BvGnH/kuthMDpHRRbPYiol4wXTarQIIiQ5MSqMDvQJMSrNnmMFbuU/dWN5Se69ou4MIVFlh
CIXkMxd2R9+cCOEBREpJ6h+w2GaLnY++KP57NL0a8Z9o8MSBQ84iOIxWr9orTRUmwlQnNvlxWUiK
ShIdAISVHkRUft1jMVFZIgmdAq3QP9geoP7Cks184QmKmMidBOgfbdm57ea/gYj3iDW8AlBY2/id
LI2Kt5YmHYD5TA21E8fMIKlJixWbUTJr/V72fpnFn1VzGM6TnmB4qCecOaoQnW2mYF49zQA05Pzy
eDhZ/F14C9R5sHdeoTdLxxfrKGmyJ0e6xKO5+/yQJcFvMsC6Jjg0o7icX1rEibsFjtdsip1Pq7P4
6rMXkv3EU9CvVw5ZFER9tPzglk2UUnPExzj5kT9ntp1trNYJrE42izEtRffeqwUyLXXOW90XGsjr
LJMMjSRWV82AOAv+RewBf+SoFkr2K7YgjIv9PcleMmJAICVyCN8+DObHUjboOXdaUcKiTUMR8L5M
0CiqQqNCTp1MJt3dUAvLAPiM/ni+8wBoNe5hlBmb9ZuvVLja3RAuRNQIgAvoScvKqhRSEF8+V4WU
Yq2IZJ7oFYVWhlnJIQ4ZU04eKXqa4aUYpF3MZfo1KtJAMjXr9jBeNspiWvWjYasZHJ2X2Mk+V1OB
rTFYc+rpUfzX/wz8VzNlUu6e0tXdarP83No7rXaHvulIsfzzaCnDe7zBJxwMI3GcvjPRlkVxq0Bl
w7jnd8UTu5o2dQetKTvjgRK0eezyMyFQKYbuoFAE1HZ/b4fKRA2eGRKt+PNvR/Go3URgar4EyMOv
iVbZ8vvGWGez1xw5vEVGKAA7nqtbP3WmBcJ7vt9gwdB3lrh9VuSOCcHtcwfMCb2hEO+Y+aGgnVzK
3OnRhZiP4KJcBLc9E9nFsv3UMczgunDfQk+MCBt5cnhgsmjT5kObteIpGJgK36x67V++rBW4mDZm
gpT/6GUJclTlU/wxJA3OgYGwS3MVU/9Sm4QTbU1aqNS+pYV3YW8q/aVR+CPmjzQVpD+9QzTXz0/y
5zx0TPR7ceKU9mzXICGWeGUtGp+V3esahuCPADqIW1n3N5v9iPyDnU1izw7nMcKytcvg67gVHpbD
aAvgR42CFzNSMxLIxY1kJulxNNqsO53NPkTVy42F1E2mJWjVBAdwUmgmrsQ/AFjTyT7hqKt23sxi
ryXnvmSligh0SIqeXTYNGFpWfez5RcqMma0fg/DdMKaJSurPF1TuWZ9+Bf7FQG59OtQ+Oq9spa/m
Et2YuI9T81bk1OTbHinUClsPLsiKlwfcnjbCMM4/bnI7fdtYRq5KnMDXkGpzXaE26r5EIk0EaDF3
vMa2M06srr4z4UENd6gHkrxyq1FRHWEE9MEKpm+c7cVVPiSuheSlx/Vvy9dPzVaAj5biBSSCkksa
7D1sTF5PyTfdoYCc3wfNglivPWaT98RhfUzT7ZhPd/j5MF/6v3CLvpfCym75fmpyhb5tQyv+iGB2
qLv555TMtOcK8yZTp9D+xENM97T569nfGtQAWM/tJa4y5al4mT4ZoGFPUREaNiJ69n7E7PLnEYuK
/bMOL/Iaqmwi47Xaf5iqyjcEDH91E2ZYBN4ft2imte2dPDmSpoGdmhdCAWfOECLqjy9xZdb/J65O
WcfBbKnz5k+P+n9sQNRFrWdqHPgPKzTD56CywjZTgxWT4K1sl1Bl65VW4HWO2V0VeRbqiyNEyRlz
ninR00DdHk+iJgDhvmcy1GZ9e68Y15uMJkFuBnnUPCTMmSSKnG+338oGPft+CK1K1yLSpHOJyGRf
2bI1HJShVo6qsEYHOtlXsPNM5LiSJ9FWbgtlvAmh5g1tUwdCFrz0YO4m6S7822jgCl/XHlyF8xCq
DyQJFvFgWe7vMVebVwIBoQJKZ7WyKV2sv5v5I6vB8Qpwxk+CPlH19Eaagqe8YSW38fhXKeHjS2M8
mnuHCMynmWxpLLUQI172xt51up2sWZKJqHz1X+Eno9R5futvzWG2H7J11WvLglI4iag6Ij/ysy0d
gkmbCeqKmBE2MmL94k0NJnu4woaovKdeUtwKUkIksOOKRo75eJRuUFBGlkAWyC9AqWIM19asi5PB
igpf25dWyulvB3PmIHKQoegChAQf1iDpvgEYuhzH8uV99rmycSBuqtD3XzwT0CEyIKGCgMds1+7o
EQ1D7t8sNGyj+gqHefz/I6AsV1gIVC2VPpx1I2ZFZyuqMQ4b8AgfAM2djPBVwfuMCklxEZn5YtKy
gfNU6zHKQ478zUrvSkPBNWxTKZIDmEitC1f+1rL6JW8ZWiyq/Hrt51YTBGGwP7CP4XdGhXNAkZ9p
hgcQym3k27dceqf08/fMgSsGhYjgtjcg1GZgccMr/aRn6at4++CuU/f6uNN19m5XKmm9g5IMgYT7
3DIL1nczQOfKmw5SXLc2lTj6PWvQOtmcEX/QraHzEhnHeTQLmuG1lEXj5plRjmXL/NJoXBkxUiCI
1A+At3R7l3jynmINuSkk3oNFsr+no3zVbbiXbYo2BM2e2SqF7CtQTDx4zEXjVL3vDyYPdxX2gxzM
W++Fuw0y9u6iiQ8p3ucSLJlZCsJnfMwFH/JlVHXifzMP71alsoFYWfcWfI4myDJf8DlAASZzl0qW
HStYvVk2isbRvw5F2e7ZW/vtq99vH1zM6J2ULEORL3AEA5wtfhcmr/NrEQj8GGiKhZQKWDofWAnU
enUa1ehYlrA5hWvKmi1b/50FRUeAKVtDotP1sjhzbvy6tmisNKe1Twu0p8I/pGn+79b8akRzOiVk
eZSnhf+DswgLbXYS2rY9rFKokImZ9hH6gkU1sdR3DInVVYmkRlZzdtBqxb2nK09Z5hgZTD3p/qQ0
U2B2UgobxaKZ5at8BdGBbypDAC9tSZGgpLgYz4Y87BiA7Qfrep9/cLZ5cmyi40XwqorTxkPxb8CB
/9VGhD9Lt+A0fAe/nHuDl8JL8ftqeXMofAGN6vsB4GMsg2LkbG+82sTwP4OsDNI1bqg/4kVIi4CW
uDiwZkYC4YnEtiIwIqbdJyIRwMMT8w8YKRSOvybXLzVwvSylmJs4QuMg5kEHztXmOxhc7870xTIb
aCrpyP+bvveoNJ3HIvDVeCD23747DgpoKX5xj1ObEzttwp3Am1LCWaXMmD1wXLBp049XTNwi1S2Y
QoQiPM839hVvwFwSzXfvxD2cc/UamZ154B3Le9/5vaCvpv8d0LXzi0m589fpDHuBHIovrYXC6CfU
Dy/E/TMnQ70XCEMqEGwgmln+AURthX5VKlfFSRL0eayfwfIC+t4pTv9ymZilMwGN+qojvYsGeBou
NZI5OmCML84zi5iImvergK03pCt2ogujGz1LO0QhIvMyxhcGYc92breLJHHeYQQtF857vIKnWaJp
Z/zMG3osmz871rRrTYMARleISUuhAP85tyT2Zs0gjkUbPLWOISyMBUpoVSh5SUAO6RTCv7K9se1H
MfaToYUtD5qPojDe3aIPbqdDW9Cisv3LNDAoafhJ2XbYknaowkWK4Pkq21hpFxGWuPe8fvX8lsdg
Cb29HjWIIXMXLa7MUNvaKGx23bHt4MhKzkPwIVFHfDAcj7j6T/d+Tx07r/0vCMWbIyEudh5eQS3L
aQ83ktBoCVwcdURCSaxGlgXzF8QRn6rImrkC1lgYAzAGnISJhkOO4qrt4fuOmlZ5OdzATTHQGyEV
VQGauTeyGFlrZURyQ2HS9nx2z70dD9IFRY3UidwzP+sH3Ba/O4Nh4sOXJ0c3buS+PJzvGPk0fEoP
WRqd0oBEbulYmJFyEYv+K0jGxWLj79MThwqB2s4iB4W4LEt9HkcmoCs9WEzFbj56Urh+Wn2fRhUF
sq3rr3QYKQvn1MRb1zUo/mWZ0yWK7xcYrmqNmEwLojIUjBLwhsgHH11ZrTHx6hZS+Hx624P9e5sz
4joszAt65fRwLMIN+BD2BNM0rRtxg4z6Lj6EDkL6sQ0OSRlRjAdCGW2mo4MMOYt4NiJvJQx+yOkL
/GFleaXc+2Gn0sAaDEcmS1klfs3YOAHxJw+aEWZyh0wb6F8aZbjdWDnqUAZhaEW/qXpAX7mhTY0D
VTjU0y0DY1M6J1n7dGTTBpmTH6oSz4Z7EH6oP2zoAHY+p7B3jDzGgJkQxGMX32x/+X8C7V1f4GBG
0TOmqwlmg6SHND0gBk0+ToDol7SD9pA4RP8RrPxRkp31jcvjCZ/iSwM0y3GNt79NyqpFZ3MO8gP8
ZU6njZTVf8Iekmo3XmGWmb1SLOJZkJFfspMt9RD2wlzo97DCLbz+JLvuNhYgexcwyKirwAW+zKVI
GBYo/EU5DbI0CLlKE6IsFZnR8f3NVMGEjySRghyBuBALp33cYWXHiNL3iUJFiTcDAuyEA6z/6aNb
+oUXYyuH0jWrD9FnP+aBDtVGQRrxNp0xoPHV5HCYkzqc/oaT0cR6Gl7n2mK5ldg8qvUG3it6H2ef
VQ4K5c/HdAfB9pRfARUJ4fxtpUznMYmTEMsvE4GxQkkV2dG81dXgxO6khE/IfeFBZ2+kuJyZHHRQ
lw0KbT1oXWz3oWGh7xvA9sVQOZKB7FbwqObjDSGX29dFJx1VS/Moxt8JXiYKzkIVlGBi3xGZJsNs
XiYz6ZFP0Q+AuclSNSlD5b+LGRR9eKXokiyBWMMl/2KjG/8RiigrNmuqkHB6IgAg0gCs2knJl7it
20eaevPNLRqxK9yOAz4ohytaoOAh35+QoWm3g3PEEDHQ9Yzr4mTGDnkB1C0MBf0MPhgqCK0x32/N
67MEqb62Ln+Ih5WY2bCgqdlf+InKJn+OFryfv84sgXHV5pUX/p33etNJujkym0DrzhvYEx6o31Ua
olB1+LUjQYviR4nrJqdy18ZAYUuqFR40HyVq7yFeclEgbYipYRyRwXf82g9W2fUQCWTwpZ90bc5r
Y7LlcLzzBVF/Jf4dPKlbD/9fkeKWV5ss1kuoBkTfZdbIYqAC15lsjMRN377ozIy9mpg51c+Vx21v
XtCn/Dq10AiQmrCFaoYsICH2PkD5yDRObgHU5le3ioH9LxfQmjdZqcQcbfq7GwcR/Ydw5S8kVett
41Us1gBjRRQ3nEcM4TbY8g89HicD+OIsokT/MKLjcE4eiPcvoBBQXN+TZItw+Jh8f6GRSwJh7Q8/
lLlNyEUs42E5HU362lpP4a1c0iTPBdxEiFnZuhCgOLu8AF0QLs0/FE98WYtm/+mI35z83jlzbRNC
mT1pejXAbZbKNorQxsyX6mLNd7hvy3ro6VMGP3B0tPYsiYZB/mYJkZi39ST4aSMy0djo45QpkeGy
nvCHyCrFyrGDScEZ17Ce0B3ef1YMA0x+IEabjYCpmzwRgKilixqrvkTQPJbDQevUqlz12WZwLwCA
jzsb317D2LLEEMXsflLSAvMhHzBd2RF0dxyhSPrKG3ZroQefNPKaOu5d5cF/Z0TtaJMIyDyl3D33
OfB4AgDVyANvSIe07Uj6TO8Q8AWMOXXs+r/EH6Em//YOs2W2cyWsOY41/iazhnyUmQTEnOOJymmt
S7/XX+HTomKx+EMOkRwBDfSNmFWWBL/QSjb8F1DHwuqias6rEu3LEQnDhv08IwrvyzeoJcE/y2Dq
/4OHrC5hqzQrykk2kPedVvCBtqYjoze5WLC2IIlc8Gev7RGE2hfA0TIno+k058QxAJ/4LjrUZ9E3
cLb5cywrQC8iPw/KonWzsOsvDkXoWoN46NGN60Nmcl3KpStduoU0M//YspVhFo/rNMWlz2X9lxzU
5lyfnoQyCUgCAPnFwvMQ5PDuxGqon5GDR1+7bAUAOHO9/KKNvJx3FTvbwJrsSV+AG6+0/P9afM3a
9Gf80tW2ZAlERnGHd7QFyMA6zzlOwJJNs8vKqibeP3+axMB3mWcBwcOjGdt5ZVHhg3C9B1teG2Cl
Gh2zFNjPrMYINBY/fNplzpznQCS/E1nmZY159FTkfiax9WzibuLULRIiWOdRGlTPB2WWNXHempEU
6J/B1gZNYo3uIqWqQw6jEcZWXKFJ8MVGLUrNtwcknUgAORk7j7DzpNlibvO3smBJecDgjwfrRTDn
5g5rW9BHyOnwMx3OM/1xtEE/o4bwhmZOPI1pGpKBMf8zUku4XaqSFS9S7EMxytUsUoHQoMK3d5Fs
Xmgr1XJVj4bbbHQIoDjpdqMQUj5I6BlLvYT1mDjQVMzTsBAy0ognCF8zRMn9W5q7MWzeZLjBzhcS
bNUsEeFN6njvqSPS63BGEqrvEUp7R4bqYpFFeTUIjKVlS1A3OORLsfjO3lGGtYS55ajHHxsE2N61
KVt+BMdjULmgHG9t+AM6vTFIIDnzjlJqTok/NiCM4U3+MpQR2mXw0/1ZLXfa+ssAaCJznXeuXisN
EupUIdToSrxPx8EMiWQE+F/0PC/NLD5xjuouVXLqw8RA7DDJvm+ON2KD7q9XQ8Q4UllID9IJVecX
LvdrJAWWdt/4f915FhetOxSGuiFyhoQMvByUMtZRvYKjOvf2UCE4KMgopyVCfm8GOMQ8P/aCjuaF
sgq3bPo8hDeeg39qk+XQKVyKUtfh4RMuA4+K852RUXT+G/73CSnBydNL5CmZmGJSNcYR1RT5zjDL
qVpmD3kQNX6yUvlmNoU7//6p2bZywIGb7WHXDKXipuL+dXpCizUFQwpCH1Hj0fjL2zU2ZmzzkHHG
bXIG1L/sGLI2hcuyL73S91ex6PP14OfYd6Goz1pXRJfQdviEPM00S4+rsZQfjyX9tddJuSJmYGKk
7PuirmigvyxCsQBAgIMHnvrngGYoiSaKdbiQpiMLT5kVg9ejocRXzG2QQ9ioci2j5xvEyhgEjqoU
cB+CObGda5fN6I+8qN4dse6be0Ysy8NH84lXNdUoSqeODjlSsgWdTbKxwKAf6zoK91DakprI5/RA
YLv4IC6cpQYnz46xQmQt+pHSP67JukqjlzV4GHKLHC4z4lHVhq64982dq4J96YYthmI34ktveztT
nvozRGoLPJu6D28ykLBJ0jn2rojQilZLttKHkvk6gfcffjm4b48fEYZ+eKa39jyUznpx+rIf3goR
tDBsIyhQD8E07s6m2OPtUN6JObnm/6uwztHump+Wx0ru14kYLxYzz52oAM9FKQwxczN4B4Xm5AKZ
OoeWUdkhWROteUBZj0GkcOVdttGfkLYbbA3LrtqwD7FjvdccfeM5ZVPk4nzQQXsA3v6LZdxjiFIa
lKz+/ckFlvZGylPdva7itlbOjC1bTE1PMjNfnG4L5dw+sNuAc44HdCWlsIqLq5RXwtq9itlqMCi4
g10Ah47IqUoNG/qoOL6xgbcPdoy9eCxbdnbae9BdQWHDpA4zPXff2T4/f0ZOV543ToZyjOLE4U8Q
M1rfjrSe4plcI14lMQK5O9zhzG8TUhNQHkVQoq32s9pKxmnAdb+2+CHWxlPXkYOswBlJsEH4U/eI
vJq0jzgqk2gPEIfnSuVRuRE3NUCyX5fqbGiPQgwUUWhMSznfobIRmKjbFsJ01t3I/juqffCUF0yO
Hc9NylTB01kbj2hHZH+wR/OR+Q1FTZeKRadKA5CHB6ZNW9hSAfMPzZvLHc4VDbUU9/QHBGHoBEQH
bqvXFIcVtmd1kddGkCxjIBCaNiJQaWhMexMV05quAxpG57DNpmzY331x7YD78d/LvI9zzqoqPLCe
m9sgmxgNRmOVCOUP1T/KOC3PkQKHEDdcI/+ZhgMFqWHsE54rt0baWL5wDqlBfTkpF1rR/YCWqS8N
s1btAxSp+LF92liHvvDI/6GPAB0ZqDYcyDYBkfrVl6U51b7il+Ef2sLhwxNQgdUhgewSvImLaDaB
xgAnwFAIBw4tlWNRnVjA0zWYSBYcuzmdKLjNyVvKANzVU9D8NLkQknXkJkCk2T/IC96a4ZGe7d3v
0PbN5vBpGzdFpUhv+Uar7JIZco0+xTmQD9TyzvZT2kxAmokutRunf61iThj//V+o9WMD62PGIU8V
dne5NsInP52/+I3PM5tj8lP4Byw1MCUo5BKzIcbHknabeojTGzwYDdZpqHyIh1OMuzY30kob41qI
7NfV+fqI0EFho2+VGaMoKqZ/YxPuA3mNDSDrmWq8TDffN9HUheobBuW3Awa5on3TJDEqiJtnQPXw
R1y0enGpOJscBDWhtthvNPqqWIvVYuLFcF6Q1svckoFRjYphwjuMZFXvj4zbDL/Nk7m/xwHzvR6V
RA4yFe3GHr4l5ct3HxaPVzyja9jtxLPqgjPynmix50KmvWeJNU/yJA5aFcJNwnTvuV1b1G1deF1a
foK+Xn9gDQ64AY9EKWYnST81Tb0sYyCM0n9HFNZ14chc8yx/piKx/Kh+iFSPM8kJJFPDlvoDeX8A
93uDJfyyUnvpboqf4OIrIOB0t9fIy6h0DVWDkduBY0cBIDoNus/QXotefGPQi4+H4VDU+0Pf79gg
ivjmgCgiiMUOu6LeCecKRsRVGQqgcMALb33a+eutoivpmwV2UmhnnvZ6z9ODAJhOmhGYof5wi+1b
gP+2pjw9W36AMnWlmh3XHfAHpZ3Z4CooNKFGZk/G3fvOA0/dRP9zQ4djDT1AaymmrcClLguJtsm8
d7QvJn4X/vnfi1gcNtIYjJPtr9+4hwhTFLH9UsoyhsHWYyEb7SczTJKOCXuWOMGTae+/w1yS4eG3
EWiHSZUunXPfevV/IuzLQlroj25r81a8bJh+TcMGgAmM/wG5976yu2esr3gwnZyUFre7e9AgNEOm
1JO73dZkOpW1/nbewNTCM5HnhvWHvOSlqoCb9jfJzq1mHHUvcdJPCT0ePo7h0kF9pPwrFBMvmxON
GwmdUCxJ8rXLmf4LQ5Nz9xmYHroXAL1u4OuHpNu4jAHRwtB8ldX0R54Eclqw2CJATJqdWe5y6fST
GXIeaPZIE7PhH7bDAIPZ6G/S+4waX4coP7qUtDbRhiPy81ymGQasoAfBAgZ8CZove+IfGB5X/t62
0HPlJ8d917aF6lZTkWxCnq5fo+FSoj1AaD4lBeMAHuhj7zh3hl2tn5TnGV0z3SSuG5IQ8sLtBHcS
pWPfmpIDSXZxSEztSgBI0Z4aPN7YFpND9P5mhiKQv3XEF1QWPnrPp1o9CNBOnTHPX6tUYoA1RQKY
0YoD2jSkDX0/HZF86WxqgD/xYMBnhHmaVX3S7zrLrquRi7dlDS8vwq8PVcmrtWOFOkE9o/IZmtN8
xB8a/KZMx6NIPgTMRsbtALNmB5hrCZWYZHljJB7igxRB+YCA8lxKGG57Yu83uOF695oAWs39nZvy
j8u0gyFp+usYKBmnGQPAwvBNn9h3TAMbca2FAaDZyq6V9+Tz9Hb11uIZJqhhoE+aQZIJTdcLGHPT
647/b+/i8sT4rrhwdft72vkmL52rXji/0PgFWKKUQe/lO6L+Y36rjYwNJfCIp1RxVN5aHKQa6LnL
gELIIHQGFVKT3nqRAQkpS0mNRDbUoANhDfSyceb33dW5j5RfMHmo3QGMlTQRV182n9POLmnTO/l2
ERAmbu++UExhWDu0x+WbP6VwTb71rMJXnOo6QA7EAHaVENtHcHXHpp/C8+ibVoAsJ/Fu4osMvwu+
yDH0JQlMYgPOhhqsycp/uIO6RvCiG9pNhzR0yiu/57IXze51Z8iFoAIE2H9DIRwczvUAgkTBRWnn
XdX3w4RxeB1HOvFhVdgArzD/yUfZ/EEQHr4nRduc85bNKZt2fLzv8fp6m+L/3Ix/mssiYbd4YWcU
E2iaNOQaw5dcyxFJhwUWcbrK6vtuQu6rwREW61TCQP1iYqGx5zaolAz16JKIxjW4fcvEeOEp0X+u
SC+X32xSEsqHCX1j+tUpMmaXCbhLBBJwRKkbpVctiq3n+EtNp8SjhoJDOdJcX0EMt8WIHWhiiMRA
JPHofgoQj+C+yDhXRyH/1xmZXCk1qw+HGWkFbhaLjsfghCi/Of3HW+4n6RF9ADHaH4N950rhsTHJ
zYW7W1euosJFW251urrAaiz+laop/DlTOLoK37LhRM8eGQLgGQR9V+bM3Gz9mPfWBVuwm0iB9Eud
CBxHUUBRSZXO/+zyDN9LP1M8eyvYEPQU71wg50a1B3rCjQZgkZwEWW3Rr4Ca8w/AHqOjpAObTkJK
wKe56iujxFx2SfZPEBUAatDbgWKsvj2aPP4h53+P8ZUcwzvjFOZg+WQ1e1q5hbjhPNTtsnpnNfZz
d7XoqNXk/D5aqKx109xoHoJQHoOGFjPoo7ul7Qd/Hw2+YZVn5NAi4gu4oxDZFY/dzsREjlxyDx12
KeOEmd38s4BmoRjaQkv5kYDQaekI4zJ5tG/WX2RF3APkE8CDPnDFUFhpFVcrpKhqTWrdEmaghW3l
cJUkcFd9LKpWAzbmHgvXAdwsQ8RH/GC/GlH0QNub+063iSN2u928U2Xkq2bBzLEoLeGA3ydoHMZu
UlM1dZPTHURn4D5lAiGm+v0zfFC9PsD+OGGwaR2AtUdwbR1bG9VGpMEeFZ/RZmSnD61Bm+vAAAiV
t8pbF83ZY0SIQ64MKtpQcT2vbve0/YfzvgDBZPFyXFhm3fPTgaEKur8cqtr6x3oBowBZ9xlEszY1
CdxCMy4GY3YhlMUYZd2JEtfUftt6ssleKQvUa26WrDriwLeGK8WMlO6TJyM2/+4Tlj0YENigbbGZ
TrdrVR1LfNIfzHHfyzogX1OvM13qo4U8VOyRb3mgt+sJI2yWtNwUNdWKYaLLlz2LecrxAqSMKX5a
eyYR/3uDzYsXOHgtOhZk+0CeX6HpKE9VSGwo4Z1XlfvE2Eps2pTMjSS5F3GEfpXN71g1yLTPkXvx
CIyc7tHYI5UF0cx90IqwftAF9v1Pypj2J0koAMahMIhiXKRv0rnJJVU9COejC+wuoivnrLZGNSQn
tKLLAm+Eejg2LHdJXT7gvk267ExHovukHt6oBD8kdFRt+cYcUB9pxLYlDaoarC/vZ5I5RUuTQiIx
eWKCfCnQnA7SQN6bb9LRt1mzLt/ksQiydiuwem3WNpXTxX/uVtewDV8uDEK6RlvtVVSkK+e/0qCt
m09OydVZtL0msT4qi0px5a5+/85KZ6rHZ3En7KbndU53QmpYhWXPGzRO6NulSGWRVh9flxsQ5epC
j2FpyYvU4Pnz98pKOc2ApLtIiXuDRR8sHadrdCPx9I4aS00KT8WBbjDEHWl0wYNAwdzF+T/d6QYU
h0g9M9Cye03FLeIb8/55MaJiq4NCBTEEOUHyg+0S8AQ61bxXE16QJwkKrzGLbHR0J1aU7RiSGkCE
uXngEunjihcKWuQZBcq9X1S5c+k9WWSadUa/JsdIMzbWwktoA2Qxm+aXl0SziYBFi46zsBpPE/fi
4OYxFZEH/DkeU8c0Cw2i21MSTxarweJiLHzDeSWN+iqB8rI2IpOqsOrQftMtcc6nQxX5VVpmnA8P
ZFroW1FCjr9luwvBpA6yfpEPEg45IQRb7ptgJtQyEFyJ3tHPhtwnWxt96rz5FPZuzgfsO76G6TMv
9yznUPA2cjmehcmpBqzEB9nRH6n9l74R1U02vo6QcTwOplPbXrBIggN8aNfafajYwC7E44CGjwMW
IoB3SuBr/xiF36aAqjKChLkAAgqpAmbmedz0+Eunfe5OXy4DK3ns0fILR54f4O//U57ZH9y5ZT0b
MgTabzV/KizUxsQEdekMCxs9VrQltUKrrAw9emGo9OlJT2p0l3FDsex5bNeN03EiRk1g7zvD6Fq9
0i9tsF+GQqu+QaLRU0N1hDwtMgaoOuDVz7jX5AXsF38PNauJt1JCZgOrfzXUQxo3hJgpacZvR/Jp
zvNWwuKl4LAhndNVlFxwnZZfavNT9eOXVRYCuoaNiXvBFNYhND69ZoFjQovqOOiXDvl5Xct7UpRU
P2XkYJZ59v3hYTH5Jw21ACgcqMVBCkmJRArq6XtrMn0+xEVsMXY7FR/uMDcFgHS+XjdOhCV7+562
x9749oN7fEpGM0PO9HZv6d428nruJqCp6IC/bty4ACmxVZcZinGZCFvILEURnEXcGymc2WW/MJE8
oLWcvoca3SH5B2aiPDfinm4woaM9up0Xpc+2rmVk7u4vYRUDHcNno7xyd1dw1NYJ3hysDepVqjyt
I0tF4VBJ7IKqwnmtx8qXAMmkvDOV+uXLA1kMWprM9zpqeVyX2u6A8M2DtcHvH7CBSJMriMT+6DHJ
1qE8WPlK19xsfxFClT8Tl5/hvbIa3NIU+0tuA5QltS0s1kjKXAT+RDvJUrwKqIFU2ksYoQxu+7Bx
Wmnppo30yKS/w8fG2v7pMGzs9zBkKlFSRQqfaTZT4q9FcI726nuHQ1S7rcmyUL8xTZEWP4AvPl4k
Fu/SOPRHdEaTP8/XkVfYoOuFudpLsA0+gB09iURMHSQnNBwpG/gxwo/XLVPXEs4nXCa0/RZ3JxIW
XdX9H3pTiO9HwW9A2GNajBEB40JrpXMouSHJYbE9mGqkO8TT0p3y4vH1qXDxEbKsZpADnMxQb/Vr
lt+90OXSJhVBoULzIYIA4icJ7ele/JZNVWtF38AhN9j3eUT9O9ukq6ZBCr9jtlPiOBK6SOq+UmsZ
8r2OGDGf7lfXM1BGpXUunYURhCvBx32FahlqPxXbn/ZeExFLSEn9wTO100OWoAo8YAjzciC064A7
pK+1yCSKNQVcnAUrmlnInppVRqW5sVcJE0bJQYGGWYxm02Nme5ClR+QPV2jj62941n8Pa7sP7g4A
DID1a8owMraLaBvQVOhNiiXYX5HQKgwGKbFiXU0MCtZzzmQSGjsX26frbACzVsOfyez+hMkEv96x
IPTE0xTxLwHisLTLlSzk/yhCIF6sL/QDeHvHs0qKSyUyjhR8QlvHnKdMVhyyFzzpGm4wKsDZ5Zm5
sspuAXR1OoCuwkT7CSqq4J+aSCzhFqJ0/U5DfJ/bgv05R0DEXuf7+j+EIukEo2jnR4DdzqbH5pPW
OhTyf6iA5K4rX/foyU5PqNhlRY9XalqAMi6PrzwnHplUJJFeMgRcyE59UZ7hSGSDMC8yP9BK3uZ3
pjQXcbN1k7S11qDmextw4e48IjdRwx7bVHQbqr2EWrtQY0zFt9u7Iqw4FLL8JUpiJMCz8yabUGmC
znTZss3cqRcE+uceXeYc9WSElN2oLXC9l48/CfyD4fA7P4W6PCwkn4Rvw3RoPTiUOSqNrN9k1ahU
AgmnHmepgVeF2VcmmkvDPMZCtgYxZPYBu5cPRVJZ0YTouZyQozDyat/Jym+iREPhr/Y0b7O/NIop
8fgFpRISZkmY0j+K2eA5GRxmAFaUKSOIWxQ2T2WxBjIZ17VuwInVxbxh2FyDpyTcp9BH1WwrgyZ4
DavDH5OKboey41xjBIM51PCqmNvCx/lswS0IKQ1jjcbD1WYFvQuqtHPYezpcIe2C8g9h/XxKIyia
4KRPTULeV7G389UNPSH38YsjizEAFpv9485OvGymN7f/YpQ4sEaoMlfmQ8lW/KVMqDwJEthTaPFG
TV8JXKsFqlsxh3pCpdXLjw8ce8MzBTX84ufgjXuQc+8nZfsx62rK3T7UetIGD8Rq8vqTTTazwPup
HqJ2d2XViMX48W57ssiXGtZ/SmM/Fr0Ejw9oVyLwdK2KkuKL7Tu2RqA4APeRx0gxv5NNQ+JcWtvR
D2Kq8BQJUOsgOUJtTAhfHdxDbQ/PT2cSdqr9PWwL1eMjOLf5qZf7IVDvGXPNilNTo8l7xZKN/nsO
aM4+RRdqHfKHMpn6UMO9bTzujT7I10jvRC+QjTtO6CipJ2lx8fPYSbvfTTOR3FP7g6lY/jWJ7weP
YitTP6WN4rfxmuu2C/2+5Pd1MV1ckQdqZnSUsa58x/bk7UM5OWoDNwLXLnh7n/n/KO4brcpdqGk1
pqac+nEiqv7B9prkGmzoSOQeqFP2RTbA/dukpQfunGrJ5+yXQ63XVZXA26TAdYf19honlWwNJhh+
9EQgrmWgqfhZDnQHW7pn2lDMZV51iWR0uqOP81+ERN5t4+ZtAllooj5BcLxVB8o5UEXnXsazBFbc
DrHoBgcYpXOUG9lgWR3iOSnUYpiZylJ2JM14KulRos5mxjAaZG+SNNOMiRlw0bu4IR3TnCKnJuVw
skpxT7rkTWzzvHm7LKhWBPv6NhLhq1BfDR2zavmNKvGtZEi5tlEDoTb/qguavQ2p34vOmk1FYiL1
DV0gJWSfLjAVa8skP7U0HIMNLyaXZnwoj1qX8yTJ7nlRWzf8Drybn1ofHQRkX+Mg1ZoSHFvwHTfX
7t69asumPCKiL/1u5V7BN98dFTTJt1n3TY4VOb/SxZC3Dg5EI/97wu2iut1eZEZBSGATGXtQJBbI
vDkVlwtixqaoML3ZpzCtKHxUCYRMbU948WpOjP7QqKyuf88/BCpz5KXgP8F3WazGqSupyOR0VM7O
1qQ0WzX4JVUjfkTyVIL3+XacOQM7sfmTBEzpy0szDwzsZJJ+5WlR57JCXQ5Ml3bQQroHGeCRS1kr
cC6ined7Jd3Rg0q+vDloixI+BO6+t2munmzwCtizsI6/fSKAiu4xa0bLIFLUrJpnGSijivQyJcRe
NJV7irZhRcIpXztDOwcK8KRyyRcNLUPfXnm2bZ1rryaNiy7jEcS1alm+02Pc5xupJbIQ1mF4ooJC
t+oKXrRXdiC7v9WNoxgNOHWsXvOX9rlB9SwufKQ5EZGk1kS6ya8byVGAUwfr33ScNadW15Pbll6G
1IQbVRoqCZ5ugQ1EIDLdy48u85u099TU1p4wfiIzjGJibPO44TUPQaXoBykvjIMoNEsxJE0nJsaR
v+QNcH5qvAFel/wVRH4E9mwjn2WMClAE+QndOod+cuVqnWrrABJsF20IBnZsN+uPWKPBHwhMTtl3
nMH03iBPibWSZV5euhgHWNBjd02OFg68lWE12k8wKHs9FOhAt9YyNQMRy1x/iRtf0WW/dS7OnevF
1Ij+QujqqkbArofL5sDPhECHE+aLvyQ3DIkfWDliAgqpqC8xuGOl8HeQYGnZ5TrogkH4nmxSCL/m
vUflLuzg1r+Z/TT+CS8kkmyk91dA8BFyGfJ2NwKGTHJ+1MJs7Ze/nqGpB8ixBECJW3SBZ+3UXlKA
cdNbMcv9o3VURdRhbHV5gzXpkE4ZJh8hgiXCL9Qsh1REViMLfxesqKaAz8QYv95FolTa90AH8qMX
NZtWFO+A/vdszXgdO9SJExiggLR32HrD/g/M84JyAqx5PNfKQjL2g6aLJ9jbPB6cM1qln2kAxjxz
/kO8ssYRcZquM9EFOab+/dqMk2r8uJPZwiF6WEdm30JLG7997ZWLHkwLeLhEK7ei5ria19/HVyCR
/hhZVb49zIw9UtToN/gvjko8cn0reN0Q5CVg+ymIhpCcHHUp3uKBhWETSYeU8D3T3vxRG57lQpwG
gS8RFUvmWmIOfdurTrHGKr1LGT6kkovIQoIT9rvl/bBvVJYZOAmJba6eI5w9n8rNmGotLM5TTOBu
+zDHsZx4XYFof0SYW3FS+tlrZCWRxuIsiqIxUj1euM/4dK8hYzUfIfq+NdTZLr6npqw5fTlKzkDD
4iKzTn+5DfiCjYvmHoUMlnWiwnijPosSHki64qZhfgnqi7SNAfklrZsQgqPpIZviAsmDmaa5LL4q
7Yll+FveD7P9oKgfA+U8kpgUsmmbfSNxNZHfUr5f3Ul+FChzS/FIxRgbAXleRE+ZeKKAoC3Zwz+l
7ZRdJ2YisHXozGANWLcaDAqHxjeLdkVh+Sjnxkv4TeKGTxRwA4KHz7ZxpgVnQRz3i36TOnwsVtH+
O6H+3+3s3w3YYeXjXk/dMTTD4eo4IEgo9y8ILW+isgC/1qHkI0wSIfkQdp96O6CXK5SffcA2jSY9
CeId81Bmd76rxj0LwCe8yOOIOKAwv4xbuA7j7JDt+X3TtitWagGZAFt7nJFUCCnF/6M11fJQWfEF
4vzq/qoJK4RgRgQzI0awQvoq9HSwOOxHrAeW9Rn4jO4EqAiUvM4JaDRwi0KG9bqLMOatXSWt5BZp
iQ5V5jYC0Jx2zdJe2SXc9PjT8NRqX3OaENMp4p0nDZK6dH/tIfwn08L0JIeMNfW5enkF9A+7mBA9
vgWECj7fLSFGmGzfzyFU3drLJLU90359jjsiquncX0b/+n2KK5O0umVyzGv+Zj6YuN6MNMEhwDQA
xS1T7lu4hDFCVfBK/GIyjSOIh53EGiDs+KXQE2NbQNCEAknM15qlKXcQBFNEt0GGzSK38vFER0oR
UvcMbgaqBHbJqPkVH1+BgC7Uc+R2zvQ/IygBJorGGQy2lEK0EsS8gLUahchyV6WuLB5QeRm1OLa2
6yf8Dk7GRkrTMLxkdQS4dhvSlqMYnX9pg2MYCsQGTo0YPjGO2DpRMI6AMOvN3Zh0VK76zs+hYY8g
y3ZvlEB1zDf0OLGFbLvh28wnyzWMSkZIn12tHwe+hlC8cim5k7kJnDX6E/yA8DG1M8jvGvrDzlnF
GPieczq7nCH6IYtBbOvO0RvoBn4OIymF7kDToD7ranpcLhpJR3uZIPqjMZhipPmX6+TO3J8FPSEB
TlG1Q7wJ/HuAK0ELAOuOkcvjXJ3A4SI3miKmDITPMsdaO50Op9Cg115zwWwGNds5zEbyA3ee9OHR
ARuL1N2j6oMGGMcelKWyfYFhPMkI6W/ce947nhHpeO9g/5tAerXZ31KZHeV3QLminO2D8rKs2DkN
yRYCvfr6m5UDr5pgimtsBpduEMynZTMffiMtampX9APMnwqTwTlJzdOnyoAPq5XlCzHE6wYSB7uw
hxv8JuA0Scse2jtKacVvACZEY69UG57MndwUEKhnVtoMsktfKwAKHyKOB0TBCOSuQ4bP76kizgAs
0FVMG1gEpIep5GN3l6zdjgo0fWP7psP3sUtHvCf/DmasjpZ/uO6gh/ZO+UHsrIecfN+327s+yt9w
HWkJ49zEKs061+ZmnOAKT1bSAx0FjbB2MzeilDclFRc94eQT/6LJY5VgOmJt1p8z/i7CwXx0uaK0
VyZT/WQKUCo3D1jkA1dvV5BrzeGL8eBIqd1ZnCvSwg3qMY64FKcPTs66ApG82ouy9n+/qJoyFjW1
CDKHmdVf0SQRjentnUd9rtFahRKPYlsG+QMPdV1nxcYCV5IoVSSa+nqRRrrrbx607YS3+CnmgJ/m
5pM1cnu0IYfbOEyjWho4b+X4hxP6PV6+Hb/53rB3NyeLAGYx6DIXZtSKGMc3PpaiMyT1McJ3Uu/X
XQdVAIOuXOeo2GFkjbEGyRnZJjvPejsdipqVMuCS8BttalEDkJiGJmIPzVVHzxbyCKPWFXI6vE67
9z23UxARoXLRnoe//8VDzJPm5c9qkSo19WDffF36utgMyZqCD5UdO+/jItZwgJvE5X69RpX7vZ4J
36A5VtRCtWj6aUHB4kZy3xMpfWScQYITtBuO/PwrWCjXsws945V5myRqZqrbG6UwHxNfOI/x8wY2
V8FepRGBK5d+VO/+FEqbpMxrf2NEEoiSwtnl/jDueL5VECUdc/le9r2yn8DbPArENVKjabGt4db9
PKDU8i0n+J07fAlHRYWsSMRGDdOsPUJXc/YZvr/sV/0lPAGwcQ6W5mX01tdGZP7Jv6KG8DZH4Joa
nDBQTCXzzsgL3lG3AxtRbJJyFN+HF7dTU9QZP9H+B7r7OPQUniknk+T/pK14fzQj42DLz5XJw+Jp
1qkQySXJWiza/yOaPc6uYu1q+nUp21Mr2fV8EX88blOiO6dxxqgNI9rlyfEeFpQRPnLFHRq0rNY9
3aAl+SsfyOoVpa1VnRWOzFcpdcuFw6TgkROWuc1ZDNPuUzumpY/xzcXRUnP1GxCtDRMCPI3/Q8DG
bBwXA4/eSD/x5nP78UuyaOU9qp9EYQQLVenPoFy2/7ohNFaBHqPzAT80B4hjkojUXKlbWLp8f7rx
BB/MBID3JsrAFTKCCBILJkiqEA0v9WvpdjjR9HG6PRmSUarKoYpTLuzjt+oEolkmJaKeUDhCR3pT
jCnq/Hhrc21z+OSzD0TwUIJJmfxRfi62F0lQl8jw6cc6+TPXG4z0xIp4CHRX/nM1oYxgOTjqM/yf
vExDvSAp06mVOP7e1xpv/lg9eENfWXqAlPt+LbKH7IbLFx/WUtUOC/bosQ/q5WD2baK7oT26MYZq
bsEZsRvRBj/PmAukG1cM5TrGYqJ8rzy2bTNYd3oBpykzddYeAes8cvwMNGc9/UkDuk15iKjFfcE4
TZD94NxmbWZMfW81vbC0QIDpPoNWYeqmXoLGnWWFuNScTMIZdvWHvUpBA1UZ33o5ty1P+qVniON7
K9poyeW+hkIktWrTdWFTMZ9AzlUssQY/5p579o+n2qDgquVIbG/tZZu51j+0wK8S/uoRK59g5K8b
dNbuTcUlnMr1MI3goDN5H6RnIMlhNav8bqqhlXeT1yxFztnFKlUvhDoMqyGj0VH/qCuPTU47B1ML
ZxVgmJGyVreC4QDlm+TvnwCwcCZbK1A2CKDT+n46tVK4SQss2wq3L9ASqN7xt5tyQIB0ZfMx6l54
8jlgjQX4WAgSL/cx7klQHlI36cuqiM++pUi+oVTzM6GUk7Qh+oEtYwVJ7HrxTz8Bb30A47TObqL+
L+lfL+JuDZr1aIxr6ZMCcQVJ75IY8htjaDRDEPZDfCgKiBY3ewE9DlYitj7wN4Kkg8ni1ZU4TyJ3
1G9HK4rKL+ymPb8uLZ70X6s16Z3gDabLA1lYD2tUxmhfi8EZDs8KXh1dFd+HRkScS3MjNt/Q1XJJ
dro1zvINnm6otyfbrbYm3rCOTzN43yMLD2O3pX4nGtMn73lGG4A8A/Om0cPVth50jaxgaVSqI3uQ
2IPLxwupFVJkbWrdyT/+azhnxLK04S0KHCQFl/9sFmIcqd73bJzN4fdYl6inEVpkHrMFTdLZJWEX
3a+IdckNOFJ50egp/QffixVW69v6ZtFeenKrWvT8xwpCgTtNmkRZ9H6WZHRVuy3pdqUCPtzWM4KO
nCTJNRgOG59NoX0YGUiiHVxus62Kv6zPBcsgTUXWq1GR3zO2rq/FerhZ83xsKoa3bIZiiwA5oUvs
oqCa8XjovJzXqMHeCSXjGRhTVOKVZFm1qtkfJxysqYoi3c+6W8ufBS1UZNwbvDPS+npFk/v/3ZeI
XVZw18Br2zcIUY4EFXNmWyZ/iK3Qmri6Lu4dVS+faOeMd3BETjg3cXvkcQuL4rCI8gCorAPKhDiq
51gePyJQktZ90iJIV1zqXTZ2mpqhg/46qRRjBsBCUdm9OdAb8Qw7fALrQn8h+ojBswbSEBvyZ+jW
1Ad2TwrZHLVCx7P9dICd/ZCBSEl1JuOi3dDdANlOc3abOdR0zdaDH+MnvrYjHUKnmq32ccWvDpEu
/5I0vrLp2S5FOVAyPgqyTHeiDqBle75cVszkZ5ILKyujsBvX1pl85GdCnAvtUrV99woR5cd9BosS
K3shn6ujwvIf9HoFjZPkdp0YpsCXGTWFxNAkXjfRHupeEVMPewOrDV4O0eKQlnVFfHLUag4G/s9r
GOHky4vf7SPPZh3ckdA8eOLpWEekh8ld4kBM+Vsq3yzIVwnnnmcxY0aRxo/GygBOSpfla8EjOHtL
niKAe0IoJKP2ilUTChhaosF/aPqjLrwKPUAYo0FdFcF8zfNsgqwTQ7Tff0r9D0wK2FBxxQ1FRhPi
Z7smMRNJwrx1dvr+y+w4MDccO6fkf1Rf5WERjYblq6i1nQULeqhZI3k9x7SLQiL50HBoN+wJeTCO
dp6sg29wXjyEb1Szd9tVE5HC0DeZJ8v5Ofr151ghvNrZUdJd0UQhC3/ULFtB9nLelFXjwNaDAKTm
beyK1bPU37d6LkzCF7FimQkMxqI3Sh1NI93zoh/H3+neHsW7eVa+22yWPlkM8F8+ubVuIrxV7Rv0
9dCO0jE5jnSf0+0velEO/vYdwG0ilyIl7DFf7UJUpzf2QM2qpxNh6TKmXchli3sncLiy+i8mPjGm
C4Mxgck/Q1Zciu2Vn/6AU3fyEIBwsq8RxeUM0JnEvEyk/zwv3zVtB9qBYmIlWg2o1Zq+pJ31ovjo
L21kI6IBZSFoFAMTlqKQg5qqFRVJbmsdYJdm/yDEHRgZ7fBGJJ1LsLRWWCPCuNOb5v2tU3z5M1uJ
PKmenAdSRUp9Oolf7754vFYrh0+ofUo+LJlwSBOYj4+zDiwrDBEuOh1W4Ey5XKhPLmUxrukY9CFA
BEiJk6Q9kl0Cwv8ZVUS1y/GGLvBJiWiqKxIMFPTYRzfS/9uSnp+smmGQVWwg+fvKIj2fOdEpoXfP
l2vbCuRKClGvDOlxWJ9gVby4gZFiatb/WUFXbr9/Y7guE4Y+M70mtIsBiM23++8OYO2M2+CKKTxI
4IrJiTFD48on0VgvLsAK36jcWLxcv9CeBYoFyCxSLOaQk3dFnPIpRjuFAk5Udme8Y29Cm6Ec0lBR
YNMjaH/ftaxWXvU7N8MuUP/BXzdtYUqnvzuZV6WDsQSA9s+Q8h6P9wOuTtVuac5tNkJsVHRcxpwp
BiL4MNlzp+hlMnS3ppGpN8Ger00Eu8TtdisGBAShGSjGNnQc7Y+G6TzUup56RDKEVJJ9FvTNW2PT
eWSj128P+WMeQiLgK91RTe7TWyXwQX9EfALKjPStBwWTTu0122fEbCkZsU+f8r/1EWkXf4XWXM31
aZkbKr3Om5EcGOu1HCV90udc2qbTjlcFUFneinaO7ymAeyqLflmNhMjJmWqBX7Suvs7ufft+4AIK
kgnyLlRFRfD8cKA/fbHFy8co2HZTQM8P2P2VkKWK9SaWo6ctKbo1YrBqPDhIwHpoQaWlTUS/Gqdu
40296VABtnOAz+f8S/f6P091dVCslTeXVuz/+ydTgEYHe0s7FvYiSyY/uQSyFRSB0mWGyuvbBn5h
h3A8dPrYyYI5vjK3yrjBEQ+chj74uPLJjUOAHmW5GVIQuwPi1qvz71hweSGdiQcqXkbF+ONackn9
WlKdEWmhExjENpXVN5lDRfNYQqjhWBjdwrkXwa3Sk0DxEmZhnmverkZVN8DQ1b91RZ8+g6mGOZVv
7ZerBWUnd4Wq//2bdc32kccwR5VBmpgKxayc8jj+ZwXOXamB0HD2sBAS59YBF3Wx2dshtDir4tlT
Yvdo2+Kf5NeQs36uusOUOe1XXzS1CMkoTnlR9sv5/rLCIt8K2q2KY3sA7mFLqa9NI2uxvRUrdiLg
jWvoKLrc9pVJqpjUXGuFFZ6q/VqBpTjeiRHP2HSh+/S5mDWFWcTq1IDB4BBBhLPuMiw353qEyd16
vTihG0GibV+KYps91RDUIqRepIsgqvKHQPX1NzdxKJVSTDQ5j6o5CXYVXuetRHsjVhA4czWjxlrf
wa9SHpMZ9gOcfPtK1tsdn5Ec92jGF5kW7GEsyMh6yzYWzyiwSz4+h58RFwy84qtTarjIoGZANY+B
rnCbTJKSGswLusOmEMtS+HEFvCy9eC+00sYwUHV3QatfrRoKOJi1K9n2tIQPy4H9j6gC2D27hW5P
waADSN14oTVJ+OKsC+g5p2yTW09313lCShlW4OyvFRyu0dfV7707ooV/MgMK+LzhFts6DEXmjM35
usEhD7s10z2GKEGl/lImCHh/EdXGHxzqyQcrlNm1TL4g4HUSKBB5MORZcnG886QjtU/zAAdOTPHD
03po6i/7cqFklhv7KpJ2rpmUZkrPhJHhu2BgUUbzyApSTz/zZf46nOJCzyvTpi+uB36vpcGg6VME
dIMBmO33SoDcRq1pnLT3gQjGQI0z/Mv8UTnyPBgfZqO2u/ip5Xtc1juUtilsH923bG0X7Y0rH2iG
lGmKn27bvIF6+rSP095Hfo9tCTeDYC3b8oD/Y0c3klAJM2MCfsTKnSHAGKm7G+sNlmtiJHriKDfi
OOaryz2nMXeaem1ES3neVnD+WlYgYxuZK+Q1NdumvjT/p1nRyyzIJIx6FH1jIrZxuabp6OcUbode
1Uu8eL8k/SYu2v4KHUBfld5ykUvvGtXv4nJT+Y8a5AG0v5sjz8L5zsj3AR9vznGmDHB3SAAUziJ0
hTItWaA94gJ++ho3JeraU5x/VXZ7ylG1z1Dckd9bmlzooO0VgWvn2srx3bkIvCKHlU678OnbXLR3
eeUYAycmiYFQXremhfPUwdtbM8pi7Ymu9TF4L2BwR5Qo/vt/DDFnYgcDgf3Hk4huheJkNdQcgij/
Mb5/1ZeYHPx3lj/r8+v3fBjfORDPkCs/ePl3eyb5TNohqsNbpwR+IIufwwrUUYDEBEFOw23XAZof
n3WaHAlQ0J0YiYPmfFlVlC56PJbNoS4LegiDP4Zm7TQjA8myKOdJLysHTkwv0v6yXud2DJ2c0zw+
BrQX6NgJCsCRAExe663OZzeJA7IU6tCjz1X4hTBRqS/TWBbAU/DX4sJTBavAvShpFpECeOtvXrJ3
bIuqo0AabXY/arrBjSDH9vv2pjALe28oIsmmzB6QjhCBlGu9sMfBRq5nCI+XZcbNXwc9FDn6jvl8
iDKGH8GCLdTt6rZSbVEV46QWY2vvDcR+YlL02THDzPEBVnlbtj47bFnwMVK0NH75GaJkwRq90x/Q
4KuxWQCGSm9DntbTd9YMti1zokFePW27D+mPpRU4kCcfZDmr1foE6oqOarIR93bKvJD0OTsSdNMY
veuf60pl/MGf5Bez3PaggOPGxc3GMiCiD7hRP8Mw5aeDMrgx+49RVX8+jCgH4FVxMhwPc+mKl0N5
LYLHHcDYUr9wlvTE1SKnRVI6ripTQGxsiRNCpkoISK9gkY93YNj1f3q6dE0dPVQ+uPatcu/IL5Q3
GiEZzX6OqwQqZ0fBkZn2ZqN/p0sgOM7DrY4QDqDS5gOBSJOpXoo4LcetxLjztAmokGIgqrpsf40J
ZUUWTVs13hDctBKzP7MGfok2t4pyzu2Ty4n/EphInndPK1Q/sbLylmIwhysS0UEILzYhFX5zV+4c
Yiff9syhtaa216A31gpWHYYHuV8IrMKi6H1ueIAR5gocuBT+M7+8JYYE2Z16hJCHO2fZHbCnlhIy
rI9cHpocGeqbZcxHNhXyJvNInw/Vm9MHW45FQ8PioEpo25ATXko5/AGK1auBuybQJn5Ud+rxSkWd
olb3NZGO59xrIlsoyKaP/wQenyJ/g8RT0WmLEHV+STh7h8SYMazmNDrdpJuUjLf4P2QjRssfJGdK
DbTG4J7QPtDe/ZKKJ5UFS6MHlGAcCe5vNcBShi6piUExd1Z/TffHF31EWJgIBnigSm/oy0bGumvy
n62abXWJ2UmYLx7cuixqnsKQmVHL3wv8tHN1fR6SC2hrXEACHNHfXnPZSIkgFYLo+rDgO0B/8Jo9
K/FIh76ki7kGq8dM1DO7qgN+ky26BDD5euaVnQh94rWmkTkJIrzmqnO7teB9SQqaLoHX3LvE/9Ju
jLzHIKBUW92SWJpeRd28EmskS1216Aqt2FQGp4MsUY9LtLlM6D57Nk6J550tJSPv14h/6ea1C4e0
XkDyFAIrfXyWSwiqtEO8RdHAAhn11c7OWftZ2PBgGxmowwbyiFw6s9UoEUb1r29o55E141YzmuOy
Mq0fslwE4iNlxzYCvwVFZMc7Ej4o9zdjhJzyU1Xs5J0loBYZb+GwiPu81OPQyDIUGKcONkWuJ75O
PL48kBZ4w6ZS4/sFJ3rqcl2n6zfL+r5jonqvj4Vb1nDYsVw/1ktA70XCsFW4HaPtxc5YT+izNhVF
VN/aC8KV8uCPyOkVpvSbhn0bdyebC937fxeR6Kv9SjxcedSYgnHl42+TG7UbRtf9RfAahXwnPGhZ
cAJbiwJzngQ+5iDBn5EPFqhFetq0/QUGdVxtaLP5PBk8l+XTM1yWMNcxEt62ZOeK68HiEdC+5mK/
P+28Azjps7ob9p7/dP6e69mEfnXbiBIAUAskUJCD0GxR048xHmQ1CGkBM6PZJt/+yw8ZLygzCLCi
3KXfSOo2763oCIN9UZDQ1qnJgVnqKSc6+lGs941EZwFrTD9kKilTga1Y34vxsbutPThjo5wiXUin
xzF+UsrBng764TIijCqILacQuXGnEVs6tnJYxGs8MmaBJMLnNVOoM9upWRbvlhHvQQn85eYEPzwt
8x8vxniioOyJRNh9WkQ1NkB6cB6MmGqtgn/+/5bp2nxSBK1dcDSMT/qQ5PNbcnnD4B9PEQ4gqdET
pU6aVC4sQaFrUgmHyOCdQHizIwo7x4RIUsLN16fM+HCUGUqKHYW7gebAw7EkNFTIyazkdhksb3+w
GGObVYnZxz57Wu3jS/k5o7RyZSv0rQjQGuUoC73UmgJpJcOncOccJ0pCgubF+esoNPX7pC390jLR
NnIlY07kZkCBt5p4ZAxcBf9AVoMWf0RH/A21MffPI+tyl2Cd3bb4jdbwKnekUlcLlZ46/8jatkUB
OWX96C2cyKzSymHyGBpB21v8Z5AmPIi8I8JR4EVR0JTfvyzhxjGOzaBHlAdSsp8LrG9kq5fE1eQ0
K71KAawoVuaZuYGvUK1xCCTPpV4tnROOl1Fbg6TZAOLv0Kw+8HuzKziAmorxhlCTd5rzxUDFMIu7
QtHiStkdFnS78ke2BMwW34H+tn5xtgMgXmUKr0SspKF2L8KWN/rLzOVyD6O4/C/o6UFm8frBw18C
LmOzptyQ2G2yTStWzGgGwD/dRHvF/1+6gYJ4iZdu4gQuzoAJRJ43aqU/F+9uNbK/CaF/IENgOpn0
oSTEQTH2tIXCx1f8EsCiEpAJ5jaMttKA/NJmEgC+pE08UPEPtv4g/FujUKXwZkBfO3MFG6I08ADn
UgajTz2dSKnzIuzfjvZGXUHYu8xcmcn4fMZHIi9QUhmjPTHmJc4TAngavbDNKySS7UCXEbnS5fey
02F5GXoAGE/mZeGoGac1rPb8moUaZKzXoexbqcpY4aWtD2lroHM56wZf65XyjDQssQ3gUeR7qZIa
pKArAZ9PRpWWt81Hyy/olr5pcK6viGPMw/GXcp1fRuDkeDnHJDKodrSMvKRHQl4YMeRgBXc4cB5x
DWskAZt4nVgNIv2xy2XZX0b0fbKnKk8qVT1Wap6Z6qUKe6VDyJUCHPKD4eBlu0izWVf1hBIt76q8
AEkzpfo9F0jhCljTqw6qNN/1bqfbTFmrbLc2WlG3ogCbyG3Z8hhGxoxFokoXzBQ2cBjVIkMSDmia
6yq1XqQ+SR7OQYHANryHFCIsS0bh0Bro/mVSFF7reP7aS6sIX0ni+ZyEg4NsBHgRMWpjZRj85/WO
HK6bHyoTRh92xiGenKnejlQ+5/fCAryjGQ6D6ZyH8SSOhsMOnRxa3fPGzBabDCXyUpCoxTymZhom
CW7cheZz6KxZDCJebJ0KyZHZjmOnAceCmLXD3GrkA7dn+KIjA0T1LGBpTethilBXcomJPOyZ42ly
Fpzyb6rQ+/c00T4xaaMxTT3L36AmT4APasYowkYnEtGGeqeimW1p5a9zKvpveLI8gMz178dq444o
wj553F/z5FzhbW4g3LnJ0om+YwQdiYr0cLfCd2o8HbFRg8t6FW/nH3Y2ErXBBJOnnA+0YWRyxbGP
9MblU85I/OvZx/LMcddTm4VSOB+aGb/IY6k3MMgfQlmrOMj9kLIIb4xm/OAAHGgHIYKJNfG6Z6C+
E3V3ZpXwabB9TbhWiUNlVg9wqhfs9a1G6TynDptC0B7shOunoN/yHvKkF2XwIGy4AeCU7VVANhRj
hyRrQkyRyxWDMX6mFuhOIMTuSDC0fm9K97LgpPBy4l32f1CNSKGMdW0SF/i31SnLDE/GTm5MyIva
Hvt1L/YFS1m+9asK5qYJaJ29Um2SmGvY6vzDo/Ivh8Yl9zeEeLaMe7PpVhsh8YZDpOklfF7x/yyD
66tq0kgHAJcYY6TnNM8432u6aI8Ge+RYlVgLDy2wmIRJsIu2lYfygzBItkjcLIlnr0H9zLmrmyDG
lKzIsiDhwhzdOn+W1ZglxDQXsJ7d/uSabbDIEhjihA321XaV38Z1ilkVH6qR+vG5aFRdjSjjrprV
xxFCsP8RqiyS6T4YE+aO33GKAkYI8rvJN5uhjQzELaKHvzvkyugMrQeaV+hiEvEY4pmnHaoLfLU0
RLyt8laJtVpvzjHTXxPi9TZPvD0t1UHTJcHDCHEhIhnSIRQoDl+sqDrf3OOuauoi6aW32rgZcf81
rTzejjp6z6LqM0nCNgM/GqW0g5tKuNHRR9fM07elNzSV1LdORmSpT21XDaOkvHZTakJrF0Y4/9rf
m8EBOVtCQ3bDZ+Kd3EIT+09DPqDBr09Ukx0GPZ4goNN/ydgfifrrsVcNGBf9naVqSbTwqHAsDAgt
lXvJgz1QLLLayEfpZxG0tH1r5PR5mfvv4MGYDYPQLlJvFZri13/PR3IGFkFxDsAnGDSAedSIyH+a
4qZemhnjEJQfv6/sgYIQfIrjtHlQYYiafCgRYZVsz1TbAE6XQNzHlXDCX4l3/4n3mPu33qmE0XEw
KhF88K6Np/4qiGBztpkSgeUMd6TWbjYMevRY1DcplUUx3ZbivSxUyC/h19Ve7z0WgHF0ujGDWWMz
gyT1Vzrhk/q5abqatcsLZy/Vqw6PviNwVl5PevGhdOwWfC8LRpnuwgVoh95/SqzNWa0u7/OpKwAE
ctsvJlyhuzOaSOjtJNDqKaikXvXkkeFsAjWNPgtvUeqHNFI2NhmgQmAvLuC8vo7sL5U87pnkMH0X
qktnPeREdcfrF7G67raxJ+Tih+tncGMnbgZ39F2OD47ZfOAja7AKvbc1sjmK6hpF8hxtvNVZoUzM
+ABRdpB1MntCgh/QGfDagFxFKfXuvbQvxAeCZOP/FRyR6BrkQcD4MYIlsRBT5F5lYXSibXnNL8u2
EhUFjcOirxCr9HFwxpgPy0bductO90+UKfs+jigROdAyc+MX7oE5AMHlgQULioj+K/sucA6kYcxv
kZ0pQIrgc8NtsmDLs3oet7kDeNg/l7a48oiaCk/8nAEjooPvIXsfNzTt/r2ME5H8Vx5drGWqaNlU
xwqXs+gi5Q7UKDnpcQLXtnwFJoNUWlHu1V4Ozsgx7hG63CtLMgfbMoFwpdJcLMPbwP24Hc+fgtdQ
K/UFgeWrhvLTVyYOVuCTRsRXQxOkiLUFZFhEqCER8powyF5MbDgxTcIAB9Xdp4Rsz81nC6A4ru7T
MmmoK0AHK1WAQa+hLmgiTm1Z8Nvsjua/9LOH+Mb+NeKI6G60GgtAYz9bjHlKIkP3HqOVWGYkghOy
1upWMZSxApOaj5WXFqXupKy9Rt2ZYStU6pkBNP9yjkSVgEaJVdHMmWJdhkvdXIOsAmphG0rh4YBh
vghzhqjewQ8Ymo5fYZzlaJsUpK4n4IsLu2up/GgBf+FGPVAjhh/6DqsZiAxcEMR8KNt8SdYs+hat
Yu9FWwLHGFiZz9kdruPx2AM7/fxZEcPOaHNXRMPT7c79uDrhHRxhQEb1DZW0QLZNmNBbtf3ZXAdu
quK5dMLwMfOzbz/oQcsk9T42t+sQIuuiBtAUKHOGkBbC2kGMQA8Nw5GWNPp9IBsWRDndCQWH5uGV
Yvnb8TBd8zOvEOqyd5pll/1BVZ2hNbmvYKMmYeRdpEzFLRYA8FJOtTWaeq6tvc/fkdEMEyv50b3V
BVVKSK28Fju2yzNDyYj9Nyu7/3kxn42i0KSQGu3/VuCLFc8uCtQYpBtk442oYftpsV/ZcPyYVPg2
AffyqYnIyRnPbhFvH1xZ1w/ell54DSRZbD95KUye/4DUNcIX9qLDrjcPHM3sb6Jj0yavSUTOVqpP
zGaFvFOc/7SlwgBXjddDYTJRWdepmCLGbO2wJTigNtLyEhCsfqwqyXeVjARB7l+zbi9zcIT+KiYv
slWGijyKG/CbzSsU4bLaQDW0vJ6J9OYSYpAM9FRtCJWmRMXwwu1zk333bulnzHMo9rO2xwkLbEoY
eElrTtFh8ghE5Zmkq7NDiAjRgbotQhC9zMzRh2fWEIwGFwczBuDzPu2NRjWIRNyH/j3C0alGoE7L
7jE536a+X+6Wxbj/ZQ/jj3cgNbZqfUwocB8/LnRfKDUyVYWLdla/toDNfvuJQl11zXNAcilE+8XD
6xKEtqsQBn2KcfxLc2GnFpN9qjhx87/t348UgxsfOk81bweC7QvQrIIkbWrYwZMDdbK8Q8WGtjsA
kZYd/89qr1ItmlON4grEbORH7JKY/iCmJPtc2CdR2JahRF7xiDAv+354nFFYEYNLCOTus0ufRIv8
y3vQbGBUMpknqxWJYwUYqBFxmrRqTW50RzoF+liZr/T1DsA6osccJfW8aV+IBR7oxmx2D0tKaWKQ
3WvbLDf6r7otDdX8sisNyxpGltCtXfe6muksonou8eryNFdQGG7kVaV35soXg+MtlDBFT3gSEWRX
KVs2idBnOafrnGGQ1Yh6Ei/ViW6Dxq7dI1gvnUUrmW9gCy1MJRHXw//Nn86yCO24u6xS59KRCPIV
gK1/4XYHFJvhLT+3IrVZgzcm4D553BdtlHBIEn7ONQDopBanrZL+P6FN7bOGTKYJf2NPc2SrMmJg
Yz/HOI7/QtOQs86pLv/38izIaHa342VUntLozvFhbz8NG0uXM8gLZxHL5fs3OJhMcrL9YSx7q1z2
y6H/d4ij63cHlFkjzHbktOpR2Bdkyu+wH8DFMxzgDZmFzRt16goi9ZcG4TR4kVtWNBlRzi/6gdfo
c4BNSwOOySJHwLQptWkQxpW+JqUgI/9l2ZBBstedvNZsEaqRDwftdFDvXuOjrQ/cpCgA7bt6U7tK
j4/+XYHfkPKlnlLaTYebdA7CA6wc7qHz27+rU4AkUc0o5P2bQkM7fsG2S+Se1eJX6m+rQmmQjZCq
LVzopQbbp9sNDRLPbDYxcRU7pif4opyxyCmZHNJ5xQwIeKZ6yw/UwZVZRgJrlqhNkHdfwvmHzom1
jgnCD4GYRPqOB3mY/4w7kTgKMCGHe8Xx1hjywZ4om/DBXgO2GDs/S+sxhJmefzi74/cqNjtjY8wQ
aBEO+I5fpeHkeeZ+LNtSctCWKEzhq/9/bK1ylzzxHsqXHM+VAR//SMgso2tcRgGiZvKuNmRsvGKV
wjzTTVV45BrcpNDPrfDQXl9nQDxVArzB4YaelNDnwLq7348pV73vjqhvvyOd4t9ZsrLQNqHDdK6I
Z2p+BtJ+ZH0cxNGJrolJvEKdgv6jKNUYPmSW4QLQGd/pACmEBA6A8Wr4qlyc/fzjuQSWb6IjVxZm
z9I3+NdYKcBIG87rWxJyajKBGbf8Czcxky23K+rfTWlDcmR9pAb8xtPbMVsgLXh7cFbfDw9/ZOAT
tx7hK8iDJIuedK4kfuReBfT/ecGq8tZtlhtZCOetNWI1QLCTbpqX3eWfwKd1Bq2+INSdMMPhg/7O
Ew7EM3N8pcvpRiPtHvfcskyXOBvoQpe1P8eWJcOrhOoWKB2l37r5pguq8MUTQRmHy6325X628vRq
ikdoi/X3kwgMpqpMaET1fn+RHHXu558yibuW+ES9g6O5UyBCd8aZDbGpLn43N8NbL1iLyuFljtrZ
Qsv8CnrK5FcK48sUKNMSOjSIlaHiwAOW0x6ARs8FsnNQsN1ckHtpT6ZHTBGZzPjBvMgrzT/HIaAz
c+yOZDlyEGZsbRmck3VK57sV7G8FxLow0ex8QG/HGcsFQQmImUGKkQ/QN8ToHThINTvKjeqyWdK0
3JsCjAE6aStaJGDuVZvEUUWL+sbiLLfczmNAdq/o9rxGzeXIAXf8PjBXoIK5EXJVl140zOldNW4d
Cx0RAHiHzc9QHNPi+aYly6b5rH5qiYMTmIKeOqa1rNIDT50xELBjqMMscCaVimhxhsGND7XNsYVK
xJDEt6nTdn4WvHuPr2uPqYwp6qnPalvhqxubyCDgLkVi0qvSAQ432sg2UW2rjLLirR2rc1CEVbF3
4oPaMB3YcCMEQmgYbGM6rGduloQopCKBZ1Syr2k+FPfhQUUQCKFc3/TK7ZtCc7paEVTl2QMuyoa2
VNpsHUsBAai7DlXLzCRrZsJz79l8eF8GIDb6LD8jtNSi3qv82xQw2UJgk0wdXz5EPCZLFeOK1XVT
ZFzwexL4CSdqqMSEt+B6IqB+4YzvJrhTt5gS3vxI+Nrrt6os7/zOKwTbbqZ7qeRQpiNzsDRjRVrx
99voDUd2bKeQN2ttPG6I7YtEne/+3TYAiYax+7wv9Lkt5YrGJNO0rLvaF4XuzcmkjErxCZYNM1Z2
GktCU2pNbQReQPlkQYIU3FNkBkk7YXs5vTH4lABFHYZq9jQvwFIovSYM4xoGNj/2ocfebPkIy2uW
pV2eux0l7O6hGc+PrkofSKnYxPoR1ERwX43/V49ZCfNOPEQtNH9fy6nwPDgfqBBK48cRv7AZoeaK
BP96clkzSS4NgCy2oFFiCngzdENQ4Rxlvkl6oIs66/UYoAX2Vj7+xRmo6OnCNCPt2UbXdz8FKNNM
qeBHx8gyCN4S/UCjdb8FKOIvvTrhIXZ8IGiT46ZltaJb2Sn3dp0S1FQwI8gpSGe0O5a0Ha/OwgLG
Qk6O6nPXFCRLhyskiYYirbQz9JN899w9S+ILNuXEGu3brpeZ3wAlvvfvW4Oatz6BYzoRTQs3jr0/
vmvhEdzFZXL8f6VlTEZnSmGxZXkn8Y11O6bWB5ODHa7p+Mr0UwpEnvG6+u0CWeFXd2Q2to5/jnzl
jvmr1p8Pa84NyvJu7IYy9+nQNaVHfFTdsPboYkjw54c3Zu85ZW/3mh9JQUx0GAP1Yg+vAyVeBGlg
2S80va8juBVAuBaQZIJP93hxxTnmis6+x2INVOteQxRpBdEfo3i1dcaglQhCiFC5pwvvS2Q0KNLt
6qW7VPw1lXLAQbQOgbHCgeBmytRonjtNyerm66yiUmVpTHs99JRQCe/rTS0oNIXM51fV/QHXzvTo
TjwP5zUV64L8obl71Wo4C0fYY1eJHyIMO8pYqK/GCim0FEZ+PDJUYpxJRoUdvasg2gz6ywGcoFtZ
cwYs4II0ORqBfRtsjOMtti+0OML1WkqpV2jUVx9nMw8+PYFQBtzHdjHmWAHfXcIEBOfwCoYKLpoT
czAZRR1Al8/xs+eUjA2UN/IZcGCBV43h09V+yYFAtrc6QTWXgQQNVsINc+rOGJ4XZ4Tv1LqeU1w3
J1w+/H7xDt1uWjfaOA45hWrHTpSnYTn//giJMBAq55V/3Gl9KL+m4mInVUz3oOHEhHudkOvp6OIZ
YMu6GKg23nA1jCrKnlEp5eW7qk0+C4sMNrxm+VJ33sD12SkwNWfnhbaynnmqO5G8XZkeoIFoM2Tc
zgW41naV1QJ5SsSyWrsXR5ge3JGqNzoDSMhKNiZo6pYYi36UWXO9zCbwOFV6Zl19DYdjQlwX5/6c
kuJa58VlqcSqYvFW/bsgzwM3Xbr1viPwENYI2NtYVgcIueVmZDxhtwIlH2mmqME6awWBBW8ZuGOH
5vFk1BYS557djpWCvFJb7Dhv7Q7F9dAAX7eeTnaI319rg4JRCohXccs6jd2L3enLAh3aGY4w9PdK
aTVX+4dW28Nwl0b2RD/siLlr6h75P8EgiNuoU1A4wLe76zcNSmt91tn+JAd2uBOcGWXLqqBaye+4
0QguYw2WpY3GBC9kxsPJ/LgAw9wNZZncASBJNNJq9Gd+KFNR0oUheGNTxnxkPe7eInoIxrI0Qhv9
cN1yFdGKOW7JCDwlAJKwzvrpyzqNoDhYb+A+L3numxnuIzkr+UKEUp6PQorTBR+lvHe/gRh948bS
Uo9vEeFjSJSG98f7qBPotqwjxmyA/JtbJNHvcfkqmEyhITnivsIUhc2n1xViUHn45akH5pzI7F0M
sahbsOo8Dm62EKsAsHEoYvN2ab4jsZuO+bJwXFXBNTesQpNA4XYu+nB/h6BX0Gb9LtOlFGwNR6jI
eCZINZMxlsqg4/+mYgBkb3hjeP+IMCfEHTmKAX4hlmGwgtyONIcI7GtfDSuErRhKzaiYIR0en4+o
bGybx2XrxD/c26ujvAANoPHSzjj2C+oUPUMR7uZveYsQCrmixMZcEY3iY8G9S7VJFl3HYBBNrYHB
UG9YKMUHp0v2EN9l2Q03rOLUway2J5mlGfIi8HwbN5AejiHQwwohQQz2md6+rVTtTV6lQWcHbdY1
xgN7j2FtKF3xNanEvoNNAaugkHz5+o1vt9wzSndv1+HC/cTdDkZxTFvO1OT0FZj38tkVwns4DoVq
HONLrnKyOoLI+8Plxji4SC/YzgQHWQ8umAfFa3cVn6bZlF1p60lkmMMcY2NiP5Kjbj35EZ48a58g
tWxQEseAof5/1BpWJsHZ7Z4AOdDPvrtt8iZ2JBaRtYC+2mYFLu1egNOLlMFrJ0SON77GXUw96t0I
JCWMo/erSvhXFweoZ7RS1y6uqDO76y1VTWgC/We1srcvUqGzruK4gBx1muu/CbF7rntLbM1FZXK5
yrRtE/aUPVjE3pv1VS+C6envxwFWXUEyUNC+zIYVMODn2I9zbccrjP7yY4JtnC8gjX2M6zI9yMdG
QuAuqqPdR3X4/pKAPvBeTppYz0sLP7a4NPOYtGpc+VSRDCEPUzHSR18pebnR0c0/egzkwXAFwk+/
pC27FTth7ieEvwmk5rF2ArkZQdlffeGeqDohii6OSrRv4F3d0RaAWDTfSu+5dbX4wvyXhISY9LHf
jywld3+O6MYjzWLrzrHEd2NUBflS4GhRuSYMmW9sgR644pzJZOovL0ZgHeiGym4t0u/1Nq0c0ZG+
HlHay53JyEhSy1gfxXcp4X95WKHuPsGXdOOW4fIhNx8FJ0NzgCb+72XT84euzNP85GZcIIbKZySp
Z1U+Bc+bESoE7LmRJLKwUJ9CGlhKnP0FDFq3XwDyWLb/T/qHoFKI/xEZvTUJAXRm8PO33lALchVY
lVhAI9Daq4zqome13U4ffUVN402ontjDsifT794mpueqdDRjmEor3YLQwvZJ/RuPbJKdg9bpccwG
WN/SUQmtSEydVhw0t6F2f3h8ITTgtYGmvkJcM9gX9B8zzh33QYzCNMSOawQ/e4+OiGSE40uFaX3L
UYdknc+uiTcgErAizyILYpkVwvmk+4smnQHWSm+V0eMyww8yq2+uBdZz1WhbHdnt/ePes0oJA3ga
L3LvUUJbgcIxoFQ/QmWY+3Em1hjH6xmrJj3PhnkqUbsrx7ugbyTH7C+fngjidCwh+NlNx7KgWL7G
CwDKsI0APPMbeZb7MEdFkXvOiULRGycrHintsCq8jIR0Je5R6mefNjtXScFsDsJPq0e9w7M2FF9o
a4Qpy5vqjES606F3SglO8yB9OzABLUTK6+IuJCCyJFx4T/0C1snLvKNVxDBZWHY6ggKfbOX8qN6l
OHbcr2RPDp2HIkYXi0zVKqgU2mxCpad7vGob4btTqxvYATY1ACBu6VX5EKgv52t3gwMm8+aolP8B
jPtut6kQOqgOIE4Shv3qswsJez0igrpoDGqNh5VB4Odbx9YPLON8bdwNQQWWjal67CCQXq/kVWCM
91/X2X+OZjNnw8PmukWwCpW3613blm9O7Raq4n13MJ4F66sCZNlXjywLI9AG14vWYL/dLPsm6OF1
W7AMT+sY8QnFlBsCfK+i25MZn7KzMFfXRT/dFh+EU4yxWk07XhRQHnzFr7EV4RwjNCx5eMkc7gx2
5blgAEpXkGNblpPRKiOKca1BOevS/WxhKvMKJ0RM33opStyL8+EfC7aO509gw8lqtZzirhGeB3Aq
a6KZGfhYXqo+cpDWkDZLA1QUsp2twS9pC4cMq3qojs8OHy572Sf7IRTgKmail2nc3y1SbA4R+Vgg
jHY+58XkCU/OmE5PotjvVok4zVTvO81xVtZ7m71HhG8DCKIchQffXOZg6FgwcpHnJwxjvBV9keZb
DU0zVXqnad1s51nprfIL+/N3dabYjvqwmwD35S11/R0uBOe63PKXerlFYmY7fyotQlGiGFJRCwuJ
rfjyvUq82nLRiDfq/ftWrCo9Yq0amBYPif3iM5MEKjbCBuOXmUdzdP4XBT+xrWgBv7F5wH53cJUv
4jEOS9QcQAdpT0IZUzBzxYa5gLDc3J0izHEa1taJgM7glzHnzvEqQOKznDAnKD843sWIGGkyril4
85QNpy2Mu4+7CJJ33p9BAix/3rkP70SiIbptgINn/s8KzjmBeVr8GYVi3kdUHoVcsOzGQogw9Cqq
Vxchpx5KPiRBA4vMElA7o7lKWXJC/GsOcdH1P/u1sizE0kSVgK52k+MB3v1WxxL3OjLTMLJ2qLgO
cEJZWjVnmnI5nHusr7nIfJOqcBK3U3cQwKptEASHWoD0fbCKUUGEOCI2rgFHgswsg4x4ZX7mOi+U
ULoBpmyQnsmR2DFNJn1YAeB+EnVYhsKic/+Vi9OERCfo7/eXNm86rFZ9vNVHdgDDHB+JKjv791bN
8iM6GdakOFCTGyk11/hiRwsVYG3DX8Q7FAlSEEBDBxTo11wHOerpvwvb+X1W94mN95VZ0p+dsp6w
QGjMh5w3tIclm+qI/pqiom+RifqOu61PJ4g5gYFhybNkLXPMAkg5uOa6WX9xsWWLBlKJtQM/pHlt
aKvKPEqfrAt4y2ACzbOvzFgmI+t1IaKoB06vGouvc0jJNUN5aDMjdQzp99g614/XQtnesl26mizI
KG4DR6Sej971sxbOtz1xyaVDHZHkF/zj3H2DmcXiauEFimmEbgAftQseR14e8cNa8LUiuNlo6gjP
0ekf+RYc0SIPluM7/PQwB1KAWmbK5xgZx0gsSGOLSxosiUnQ5vLdrwCaGnc8lbkVU4K+va3CRFmf
Qh7Cilk2Z9icrD/4ef4RgdAT0AkU+P+FPxFRd++Wba+iWzSNsQ4Zs7r64kF5NH+To672rpjPhjtE
Ufgws98T2FLbha7Snn/MgN4wzM2XbwE9x+jQmAjxn8CdFVE5zkdX5GwIUTmz0uHIBUsbgUmuw4xA
4h54xbhAI8l8ZdHGI8MtD88sayRtlLleZxIIpc9Z5yg7vcWge9kwAADPasT+QfrUByjRwfIBs3NB
DYXqUNEtGx1gbRe3IuK1ofdGgF3HcoTuM6PysXYqiU0gQhnNAORnnYRiL4pb6yMXehNkoAFYjHZU
tIAOyoLKtNnBkoLAjtpP81omALx5OHiT87BtwmFkfuSvqgXJX1EVv7tw73dmMz+1XGfOi39lsLmB
XKy/2hH9DD6rZMSBx4KTLYMqfm4y2bSuSZDDDZKqJp0+xUQg87RFMhUGlxU7Wn/4T8FhToJ0tI6M
U8YNuEzuaONbn04arbRATVWT20E1z9fDJHbauVWgjIzCEDEdH7xjveQa9rdvbJvShdsiYubFUoqO
cWh+ZWLvkFf7g/Gvnpa0P0GVPNjvZwXOKSiWikBKOCD90vcNTxc2VE04NEeBoG5GgRDI15xvoXja
NmFIPE6Ib1G6dvwTyoGWFNJjL+cbyacYyS/m+v18KIZj9HMpGhwf2l7g0fVwu2Cw2kVTbYY8se7Q
L41knEAgMdJgkg1KxziQ7BTvF0FF8HAJsALuxBAWWId1KHD0N0wgc3TqajiCLd3Lk3yDorBnJuko
c8EHDWJA8WFq8Ae5fQKDPLBCIiE+JdjrC0TEeyzGFnI7meRLom3LAPcpQi5g05u+PpuJgdKZ3qyZ
DZ6ru7O/qLOSdpVRZK1+G8FE8Tn010WYImOQ6Zhi72c0ey4ZTtzSEjnRMKuR9q8buXTY7DXVdoYU
tULKgm4EhlrIe6nBQnsGSDD2NpD378HjH/9XHD+ft3kcH6IFmkpTYlmJ2WvyQAQQT7sQxQxUJNis
DlsiTH5MJjLIM2caAeBwF9CwPgFEJf+AAcvzB/9WFEEPyMi76PWXqG0bF/f6sWwa+mMCz/OP6MIN
NtZZZB4Fn9ampt9pmly8oLJuFl1At1O7CmRdMljy3Rs5uVJIE+E2zB06WITj0Bbp5fCS9rv0QkuH
WWDbB2QcClkQCt9HjfSeyLxroOeRGrg3JQVaQfDvMI1bJysF2RjjrigiEVoejeNgbOLkkethbZxj
7ZWC5lq4zVb22nLxGK+fAT36nhXyumDJ7MVHnNCYyyOjKUGEIGebL8/EAIeRPM5BV/5P0EQpG10v
y65LDWkB/nP7uZgGoI1xD5O8eMSXlap7Svmnm14OFNGPkLMP3aL0vyfCLt7VIgDe1HdfKlPRGbFT
1UVTGdQxFNr1trzdwBhCF9cV7r3B8JYbtOUaM7yyzbSI0XqwJXIbsIAXjkW3rCjoqDFFjBynelOe
zye6q2ZlNmOzTwb9QruQQ0jFfJhDR76tLN4RC3WKRPQHMv+45qkv9OYBgkZBlWgVm8RqmtjkwGCm
R06W7TvGLO+IvRQwZFhBXLyByYGEscDCOMYCzEIBhGFMsr7tl9Z89x/epaAMwnIWfdy9WQ0eUCvw
BKgbD+mdKv9GdxVnegU6isQHY9gdZ9zNoW9aNHf8vDuNeFlOtZitbkuOjv7T9c4UtZjuYIAHt83q
7anJ5Asp1nXpgclizyEbqiOuI32CxxI4T46wptM7tSn6/ewy6MRve9s0J8R5lbpYEK5Qe53AbyMy
mS6FfY48Yd8lY1Qwnnab1UBkkj4IlTWRvVzHebLQbavGSgp11ZKxtw27taKwU1S26tIISGLDXhbg
Np6VxEMuoTd1ro/OMsTh3uq+2kDUQN7yOH/KR1lu8SeSmYeQ7J2wanTWtaNZy7NpW+Vuni26KGdd
qsBrbmiMMOZ6rwG9R2Zh6kkkdGJTPKdKJIfrE1DmST2ifv4q5Oa8fqLL5LuxI0UqR+zodjqhYKWY
I5azO3pdP/m/NtlgLASB2iUHUOeCMr7Fql0hVh6BoSD9MQ0ROiEEZ61GOLcNVaHEtO7ykpe0COa7
v4ylIQ+Y2t5vsvPpgHyMATjkO3SrWBSu94bk8gGWDLaXnSaFf5+J0vF3+ND/zi+kJ2eMY9kGOqw3
rL55mhAb/7aJ9wn7hMpP+6ez5K09BqlGgCCz3j8a31LTy9LTSV5qzZwkx5HKBw6JrndMLavw3m9A
uykcsNz/tqDyIc04xqoUfKlRv+iMHY6tnobe4LTRx4VCZtkvnWy2ooTvsqVsg8Fvcbhfq5Ad+qn3
pRS2QO74sDSJWeVTyCRcPT9jM7wDOIhLzDzLpf2IQWb7PtrpoMWraLtGb6KOL4uvhL3/56tEHEU1
2EHg9Q/4MxDAKYU/tZhNklUPS27QvvUnYXM8jGALLrtTvgr1zX4EFdDNbJymoq90k/cDTQPZ0/kv
CpgjnjLbqLNM2HpnPJiCPdH89VTnW4aD3hP25hVzCLVlpbfeL943R9SxfOvsekO3/BNaKpcvwztc
wWpcZa9vVY+/EPoipkbLQOu6RrlnC71QA9vQzw4dguCfKgP356gbXRHuUR4hFJAWJX9Tnw1IHr/Y
+EHjzwuCco7itCCR7whR2H1fgac+3IItZk5/083J9vGOUTHFob8POUqLceH9qCGrd/1aUizVlv3I
EIlA8U40a1BGW8HMUgPb9MgRV+fxf9mn2Pv0g3ofCRTbAZSG7MA9IRyBafzF3yy5fNY4bPHATGSK
gaxh37w1Pj1N0Q50eQwNFOk8wV0r5j3IywGIEHGG/YPgbanm1hAzzNGbm/yJHvuezGLaSKDOIfAe
SwL8Fe7SNrfIM9I7aNeMCoqcYi62UkmqeND2fvoYTjO+kA6v1ulHmYMuAZCTPxtIoWHFFSAHaNUF
LpiuaPX+noCl+22uD4Xj1jhAFnD0eHM4KOPIirn06QOjkd+KtBrJ82BwlFsFplxrVkeT49NTuf4g
BcT28k3TTBVaWqPDCj7GnH77d1qu7qGiJek5AY5haWOVlpneJIZhbuiqLRvb2gGc9y4CDSdB62J7
QC6Gb7DzYKIbq2xx6Jn2DXPin9NgWXZ88ISLCnOZo6t6lzOPU6PIMMofwO9b2fG4Fa8gYeLTqHKH
sYHN+3rjFzXd57u/hgLo5uxZ26gjILKWICHpYtxLvJ0R5wsTNXfgENrorWDGw2JQux9FXoVZ+VsZ
gMFSqasMQNet39OmnobOdoQcIOtcrb55zFDUdoy2je7oeGm5DSaTLmV/LTE2ZpFJcPle28SkD9wK
Mc2cUnBqM0BlGzi6Gt0lECE6Fl5c7yOM+SU4Mp7ijJTB4tph7fRB+4fhTQIg6pH+1qpG2I5y1LAE
aDs/M7OgNaxoANL9PiE8EJIcTqtl86QscrYIAIRXrya0lcE4SfZOx6jIelnQccFeyI+I33PB4abS
RBV3sSCPzQVqjqXFVkJ7InrNgGuvC0e0Tys/AZn/7tPoenxy5K4IMX2K8ERjALFkXpKlV3uwMAds
S4YzNU2m70gMswaomOlMV5y53Cu8/NkpXxydshaKm9/5EM7yeE8dXC7887/4UPDWfm/ZhoPVs883
Prn9lezCLAK3+fCTfLafl4ZZDC5xnW0T+F+mXikdYgVWR9Fd0p10t3i1GSdFIcp7s3of1VDT0vbk
NNajgI4bbWe4+r4fA00bfeykO90EkRghb3C9onxdjxtf2H1ho9Zf0fe8g6Zi+3tB9kBc1VL5vz0Q
Wi8+w4pTWhuaOIfZJvkHDbVAyC61pSNQsjHj4yCtr3MYJDhaI6jGjtJdRS5AWfjYVJKTPo5VpsN/
zuvwkuJD9xXY9FpTFMBauSeqdkOf43n1A5VtTux+bLQJZLV/E99kNnpeJwFMHwF4KKDhnTO8GZ2+
8azZ+JWH/H/Jlm7ypCy5AFj7eirM7HGo6o/smJg8IEKdSghjBgvCKgcy2FeszO1gcvqzPJcIgBQg
4kfGSIOmei+xK79ROQ0HvyWBtHX8YuTyAan78viD0l0GIi1U6HbMZM32VgtJRSjdmxnGYzoS+shP
nCIlcrAxDTMKAkntGVRdcpRKD8lacHV3ooUmJaRZFLESIpasOUF1+0JwJ+3uAS9/wzvqJA/CepB2
1AkFyr70bTGQjcW8aN6pF2se602Xc74pP1oJuhE+umlTII3mAbEHAve0qND9YmDlW1m/32+lbuNF
27J1RZ0C9igWBygn6utMo+5iu8xlHP6KZVvsCd/DAi/iRivFXZD0uU9fsVWPRhVJ0/xDxWacLLDv
MJgHzbM3UDZode/ydU3DeAdxi21bjhoTSeZTV3anXmmMVjckxFs3gEtN3XLosoCl9I+KD7ukez8K
jidT2QOLcM7NHJIjq2dMawgg6b1Aw4q8hzMT/Qf95O7PmiSP240bUYJaOlQtSke6h5YaaPoaD7Nd
dU0GzRLE1hXsyUH+HnIoKKBBiDtQH3GpF9EATEScBUSwuPJxV/d4EpHrm0qwugE3FICXZbtSvzns
ADhu9aM+3PRVO3fzDBQMVsaj1ljjt8VsUhlanYvi2yeoY0Rgu1wjyuW9z3t+w+GNrIEmn+E4qGL0
EG/qKYu5JlHCxgeFCmZnQNzoFYP+Y9l6aBHZ4y9DZ2PHl9HnCpIil7yhf/zVUY6p7wDb795u/tuG
qm6h1FfCl+6x1k5yZlMYOgFD4oTEkO58qFA7jmPxOSCTIsyrXs+FpYtvJrxtMnjtj0EL3A0hVjaR
v+eEpyGGct5pT8ctLMAXkb2sfkL4d7WUoWbKkSETX+JYFct17nGwAuqSlxF+iX+9Lfm2hEKzdV99
SBiwOcMTUxpxzNnLACAKojD19AWkutpx1POAlpQ7CtyPmpItdEHmov0L7zvZ13ZKL7aO5uXs+iIZ
C65MWze5xF+Y4KWEnP2ko85PcJvY34r9z5QE7dTR5syHZU+AsDZDRUhAHDUVf7MM00wxNYZvHUcY
yB7frhoKHEVaLONbBMg3OdBy140qsIxxSK8E8piu3dXtHEnqH5fRzv+gD2kNxBLq/DrH91Q0HTo0
Jtctlsebc9FzYhZHrJiFny5KDjMWg1JzFIyrFkrmYy/GJlqKkC50PDgQ2BTCmd7d5K/171pxrNy/
6V3kvJy+Ccq5zXkD6Bp1/6LzISsqGYZhqRy4tIfeRIpfS4T2GKtWw7ZFTx/Ixb5pmRw4ALlPWRk6
XZ9x4CidEHg+Ht74OxeTWxuqOZ+vMN5sbqSBdOO9tcuSmm7uJ/iQ96IFGcKyBjgPzlh4BwoyVw5w
ZIWISTgMv65CEUNf7NHPdWimWyIFJZSAmCmaUUa6uD8a2BjVCHq6jnkHfgIMTrDS1EDOMFyJJ6hY
rmMXjcKI8kpyr3PBe3jyNiIzolcpLi6WA1CbM5kwUZfeFu/PSPE1GsXfzB1+kPIbxQqPtmjdjj4O
sMDRE5Fn+ZIy81i+z3shI5lA0lXOXAiG5k1HR74Ru30dXMVIQI4sVxoSIvPMkKl4CeXAXWaz6ba/
r60KdXu9BqafUs1sbi8T/oisdRY1LKdL0YkEqAu/8ZPomhfjS5XaZ2+sWMR283L1x0FtEdT13qTK
DUv4VpBsyHITohbKruF/a/ZiAnNwtSWBTAPoKBFFvpJNMLGJFAO8yGoVWgcSrgFPmZ/WrlKswJyj
4Dsz444n5f2aJNi2F4sZNiHuby2nqZO8XJcCq1R4Hexx2NaxS15Y3YDBuDfy63K2CQIbGb2OHL+4
MddjV8o5IfUI+2MVu6RecUmQh6jdPxK0nS8T17nqgym/ZloRkAnQzNj+OP/JRrsFHyIuaYtfdoml
UPFeyU+GfUEo7tgk4bfXTLhLo3xofC1GS3JlyUkWhdKLBpvTpjx30C1PYHtTteHqf+ZA4xNNPSJe
GxIVJlxQTN5HFaZi7FbkXSBndij+wC7gVXXtumHwjuR71vlTY5nLZd2fpof/RRiQfBxZEuqhrLxX
g4ZcDhfxUhd+sGIZix6Mx7ma4SkzfL5oz3rYuoLOWmMHat5v5PmrRgc3DfUhXINynI/LwCsdsqbp
cCad1jax56kPTNaVxPOK2kLLfRc8OsfTPGJcifPbTYSFoWYa3BNjGg04esFDZGEJxIchePiFJQD/
7pab66fLfzaOoC3qMkpF38MOpqFCSE6Jc4txS5UEw9RRBmKa4jNo56zBUKBNcpEeF46ZcgVm/+qV
CYof36fTotGCSm6BcJIDZVVKL6Dot/ByV7ZQRvdj42PNgLIma3BbJN6A5BEXQ/dzpFqenPEVw7es
7dqyV6EpFtIw+dMt+Cgp5XJ/MvNBg0OJgYQG/4lT/ZT0fe2CTGaq3W8yzJe2VdvyEHygpWdDezqI
fxwcueUadT7fP69qvWpAhOH4SEXSIcsSNVHJ7Agd2b3Vq6vvbg9fgni6gzSpNeWVOcxZp/uzUc9v
UL4KJS7yqBbau4hxxZ49SoJm5T0JHzDz525pMKuw3tcE+XLPwpkMYBNhAPVnT0WIDPz5nzCihs53
nLWLMwyFDm1k7qs+eVnQfdSXx7bJBN4nmBKJsybfdEr3RQh4VjapwwOmSviVI0eWUIaAOV7wtE8w
gF4LGDUawNgMsO1HhRnBp2FAbtYVT/sXhPFG/g1cuebxkuqE8m/eXDHMVYEo+AAL75MPiCmxkg/d
8Lh03/AaOiGG8ERAbYUupKCFh8kPFJekETFK8TapvjQwt8ZhQGQWys8867hoi4c3z6IPyty3JhfN
N4WE1eDSCHOw6e9mB44TXv1vxkFg67FglDK4pyipU3XmcrGKqHtWukWPKbW2itkeGIgy2ywyTl5h
EzA8vH7PMYG54wioOUaLW4aJ10rJhSbxBPkxxq0UmNM5//qxyL9cr3OzJX8XCD0RhtXNbdLWy3Ai
zfDo2TRRmfqPWf1z1oyS1jcDwPa/KUhFlPPDwBDMistJ/S6Kis0asbdCbYq/xHWZO9XlO2r1tRGE
nenFxDiguvtwUIM0uIof4uH9KRjbXgtXbqSH2kZYgWYwl8/LZmHLIlQUMBo3aPqTnAX/KqbpUJ/D
U2asHETz0r2BcFCn3EOvts2fJ9GD/IG2XL1OwPd1wXXf0VvhYGMfUlw80PSt8YS+Xbs49LDTOPtF
k5km4YCWUpR2fhGXJtvS3sRrcWo2hxlLsGoJM/iJqU0+6U6t8os5VDrQ7hsHxhloU3DgVqruQAGT
f+xeLaDJXEflsIKKDZBGUdN6mqpi5F3aoJO+4rEaxxJAE29CYYVn95rwnz2Cv5tFupM9B/N5kf/I
x70ym7Y7cxSJm3KDR8JPC32L99L3fE24QlI3eJsL1pbwd8doje2JOngTbDJXumMCpj/WA5/KLXmb
7Z1abqqapuOxdki2zqlttI9kYkdFIzf0ZjtJRaX3j+Ni58w4eVmSCv8Xht0SIhfMZ/TCu1qLQ4NV
G02Mf3AaUYG1GN86FTwNY7oLJF8uPrS0giusmI6161Ce0WhzqegKGkvfjmDuY4UE1v3NVD0qbYhG
5xpBr7hQjTbkMvDq4bIn3pOAaqNXVqwKGX+NemLuwQSIQ2Vagkgz8yzTMv8Q+KK4XAU0R3WOMiIO
eEEnKJoJbPAHBlkUx4PJyCeZi3pDGf4oRWBV9slBqJHDHfTu+Kv86ysvwc6giYrbzwd55BZuzS08
0NGvHij62L2NMoFKTj5q44ry8Yz66N/6xk/Q7tDPQ6AkZHLYk+hjHK7/O53iap9NbGvaYBWBF9Fj
QvzhoB+JRX3NBpokCCitKev7Ujbvp4W0Yl+56MG/LPs12AgTHpkGU1mWo1CNBtZzbWc3MhOiVZPP
NuhM9CpL3SwdvTqO+fTXeYqln5ILz9DYXlmXqfUDGvtW7B7cFlLyRr0dTQUr/CBhEo48GIumQ3k3
QUMiT0Fpzo5f7blCKTFfwnIaE7Tacr13lUpL7N90N65kx+0/p3r3P6eRe03kFe5hvJEF9dMy8bfB
DEX3xQPWZSvoAHHerTciVDBGX4cX5QUGQFqJPKwqlkM2IVaf7ExOZbHeYUw3hkVpYrNuP3PG/jKI
EnIJPX7Y7Hzb6yveK8ANkKy+KqkCV/OKTwbgFNlKJgDmeIMw1oJK14td8WM8qASiRQfMdESBJbA/
FOnqOoHeknvzbQLvp4n3dAa0I+OLaIstmFgwW8xggKYiIIKabFzQnleY4N27sjAQbOlhasS85lgM
AA3BhzSKlbAIdUHlnJ6N7PkUy9tT36z1ckh09ejv0OE5B6KOj4yh8oNjsk/JR52n0ll1q3dlrhPl
oHSv7O5Qy8A1+AdkZHDdgylGX8sm1mvMO+AnARQD9pEVOxJ9hgjZPBhxED2aDZsPfLaY4EREayXl
O9YZMF2xHr7SYk95Y0FwqJ/WQhUKxOlBTnWVi3v9uGY6IHXpztBHZ88Gb1l85JAaJfJQhFL1VkLi
bDoGUqrIEPHogF6vEY4XJT5IwjSTY2E7w4j49BEKh1UtxGVQ7Z2zgJFySoxo0S+nCBNIQ5xXnRn/
GnZFTo6tuN2dFWnE+5gL0PbBODFcEFdX9//hEJzZ1lqQjJLv6cJWN5iQDaCefiYbsekza7ofl2X+
Ow0ul4E7YbxETUzkTuRiXSO8gsugzCUWQpcHM0bJlGH8OzmwbRxiIDTi4jotsjLqAxwzhSHeCC2K
aIDe2jGJS/n87Jlf5GFr9geF52LYZYPCCEwNRe8OdQ+kQi/BxJRX0zmM79TndQgoQL2Iupvk9Qlr
e757VLYNC0hNMDS1ZXnzE8kzRPlmEUocYbFGa1ms/H7etJ/p/uARMT1wkhdKj+M/4mD6OY/zjWtz
i8af4doOwaLH0ZdYQf2Rc6kiriC6/1KcGHTonQm2IUrgcXK28eDxBcFB7w/FWNGSzSZTFpu8sxI/
WvGcN1vf+nke2khtfxZM02oSC/jnPVdleT4snsjRTOUjrwHylH8A/JTkuC7RxAl66Y2tDy1hLL3h
Q+L9FZWH+zYMS3oviOfuueyKl+01WIsh7nz5UFX9v/4uXj2f/QC/Qz/k6gospnVvd+EAFopVfVxe
KGMRVS3+cMRS0HMwymR7iiqHpLQ4UbRM4rlz9j8FuQ3tpx4RmLoNYwd1u64weh8tZNJ8xXFFjZQm
a5SXf1m2E+H2KPqIH9JGemLVsPN+uUUpYhN+FrvGzdjvZPNHzy4/4VEEMCNOLcugcQMaoPaC5cyE
JDP+7A//k2BX8A3guWSO0vmG0g/A/XYBImQOzwksZXZ2v+yYamIHNFF1gURImWKfsX4AAx526wj0
mYkkdSSloV0qX/oyruA0PFObbXSQlJZUYBTNKWWQmkc2KVJcTCd6U/X0flEj23S4FYtwROVrjIbz
qB747UXSQKFQ99GYj3QPAUFrGT3tByQ5GznmPGVAOZ/JkREFiDrTQk3g4sz3LmlVDe5Dveqzh9KP
nQuYfSecve4rl20nyAdsaWkSOQ0d0UxTWJCX/w54kR+k4F9HfcIlsVdXqaAlv2I3SEnZjROtVlB3
lRjZ9Fg63qS3gNTj82F3vHvPOFsLehguIaL0LGjda/lLGTKT3ula/AsOn9H+GTXQ9iX4BZQlDLZB
vFRl+giJE76RJ7NCMWDRS0jiOJ8CsuZZnrz3iWeOeBZnJgi0ryfVlc2The1lbPQpVdiY+KX9wZA2
XDOVCMiYlruOsCMPRZpmplEa4shomr8JQ02tJRW1hDc8C9S0YyN9Q2CWyj5uq8uRa3uj1kiVeYL7
R0z80qNrBlZOFCGXtFV9jgp8uexUYZ+J82SWZn0/knI774x7uyt92OPq36sGAEqIKbKJGMPSqJzp
VzjpAz3hCITYy+RuHnZGRnl1j59f+y6UjsfxOkF8g7quj1bwfMArRNTXI3Mjv2RtV4YDCAuUMsUm
uogffSbhc7TF4b5L8y/LjroMtTwrhzYmj3KpgYc5DF3GJiddxu3+HF7s5q69KZDyViVxEU4uRZCz
tnX7lTAqlQH3sC0e4cTarfd8RRnk5luBAeltvykwJV3S2e1vDG8s+Z1z/1YZKxm3rUvxT+TCHzZV
1TbJ0NvXLT3gXgojjqAPBZ7nnVsyZ9BSWgSIlS002qW3cA7rMT9tF22K6UjYNTNs4GTroT5mpNrR
UrsMBfIwoBHcUHjPzSSXcNm1R9Ihp8RF2vBa9+QY+MDkty4CzgObSQ9Q8iNExXXpNLyVjFeoYuHz
KqEWSxOTW2wJxMVHpSEe45mQAqNGO+8OyVdeMk8AxRdjUI63wl6H5Xvi6YrYViAiExB199uXEiNs
4Ut34p+MT+2l2DQdL3vbMR/amTf1ThyWwSpp1gWsFSWfAxTDM4p4YT1ZbBGBx3HL6WucUxNV0Awh
NEjgVR3b85iEl4+C18j4AT40zmMLSs+hT1mOm2k2mydeRV2PDX9i0SVrbOVvNYnfSquEcyJKp3jJ
eK5lYWo58pOJfJXGTT52f9cSDjN/XcNgvkWc28ONIDVbkSv5r+zO2o2ukStpFrf3AbGoDhgYHkcN
4qk4FZrDHWZ6E8rDfHNM0WF/XVOyDeN7dggfubOt+VeC2jnClyffibyZP9Dj1NiKShQGIefhiD2F
ApQ4RuFOhPQgfNtwqB+6hQwBhL6ri4fzbYMKHCn8ja58EYYVrorZ3qb36pjOhg1OqchtCJEYldT4
xb1W91KDTgYdVt+sh+gv4x7z0awv8MZNt5kqIQfEGW9HJXI2j87XKZCZFHdVNDLVmk8XM1IfjWfi
6xetqMUwyAtBUvXNsYMzpnIdmmlDYKTwQDrQcjQNITdL6N0hYImY2xGMQWyF+13cvsUHyLTzVBly
0xOdGBTLKw5sXu8uL4V/mIwvd0hDCsL7vQ3xKjPc2R+oE8sLXG2l+eeYPmEWgI517U/UrkgTfBIL
nT4kLKDSsOoKxCHkDEuSYspHt/CcSw2pFdsvy8HOomiqsSeLxiYdowA9OS/4BHGpnfHQjpl63TUV
JkXcLFSwBzcz1kSoBCrwwbBIvQJHo6IrHQOlVvUt8QpIzgCxxN8bwPnEwCPOLQX04osAboWcxaRL
PeRqSjktJ2xD+SXR11m30N7rb04YkZH2M/0fAy/8MS4EdoAyKUJftPPiLYwN5a/AsNO8UMU1uCyC
XeQKLIIVqjPQnVB3YL9KzyE3ST5iSNrkaum2AdOZD1u3yT5S5A5BB0fiEpSwnaLLYGc1FFgcH3YB
OIbel67ln3wB9o8x1Hv5SDUR0JKNFVXRdx6VGPiAwZlQbA1u3GpMkxXa24Qeymn/QGBYIINZ3oQX
GyYrIicnc7VusDcrx0bT/9QFs2zDVC2YpYk52NGUYqQBc5wuXCe2tup/Ghv0M5ka3W6YQXRfeBVZ
GURhYmIY6y7hziDn3pCxFjiqb8ZEPCDsumfxG6mXkq6LuCwiM954hAV2chj50+dqFoDT344L+DPf
8Gp3lz+LxvZ1qnuzlqE/QAkJCMO1/V3iTJmA3ofzExZ93Pln0ufI+/plEW5hYnlOPJwsHblSsXzC
GpPWq0nXrvPyCZvNUnDKZooqMIuJuC3uZJbhR5nU2QFn7SJzaR4oVQyhX06HQjE8vmY1FRfbTMjY
MZ1NpSd6RW9IM7Hv/T5CaFwh91vCzXvZMOLonlcA40beYxey9l+osu8hGGQbgBG5uQeilUp8q+Cn
35H2zq3RW3zGgj3HX+C+pRgQjcGZ7qrCh7eJxXcKrU2Eqf200LIYmc6VJ0XuY+n2wH+4ZJf2UjSQ
0ZUIwUFCXCWpk6mi7IxSxLExYwOZUx2oeDUV7UVS4Bkw4JFssihXB4nmH4mg4MjpK0bKBsVIp6U1
21WVamoxNMcji2Cviu0hyzDw4/CCOOWHppcdN7cH8B3O8Fxu40stE63r7Yl6Whbl7nrwoUU+S3ZD
NCiKu1RtXa7/RhbEUfbrPDi2FctCBfJNXCMrI+FVfucQGkllgIzlJi9BArFGxF5/etg97Ratfmbu
mD1qVIN5r4yHBEY/CmP5vJYgiSnTZwoEaYyogMCU35m/4y9KWsr2JsTisglhXvp6YaqXQ23LrdOE
4Q7fkizKekNoshjbVbrNz7uc09KbRK9yOk8JdyFKeP8DGRLO3yw1d4BC4vORA6HHVIvMePq1qBsV
fv78mCEwApp3qrnPBGwBQRgNfdVyjWcIyYx4ZFPvP4pr2aKg/iyN+roW76P4I9xTEslbDsa5Ip3k
Iir3jowK+D0AcSeYGvBwx//fUrR31QAGwppv1uXFMhyA/drVOQg6hQj7lfMPM+KNUuXsODhajVGp
QVwlshQ28cawEgS8NnSE66kaGG3zipCzcOFJOOOI5Ya7BRUfwOe2RtlDFaFU7sg0O4y738GyPMgz
5tu6w2ywE9Mo6hvQ54HCywdXu8GaGnZeSQoEWV9KXIw6CVQ/rwoFGvM7PVOYR/lwYmWEuj9TGGdL
xPLGCvwGq3s+trU69I7gtyz0ssHqo0XJuDRHr+7TZhJXY5qqM+BOBY6iUwOiEJsPZ83+aD0bjsEm
lRzVhIvgZ3GHDC0ULoqNqOEO75qHTmRWyDwuKu2FJlDAcaqA7Fdr9DX1bqroW+QhS2a87pedGg8h
LXrmxGGWpDdaeXGZumW0veDR00GadunVi+egJW/Oc9YVEj3t809Jnq3K9hG43CS0kMaUEQfmC9Ry
baz57FEkgq3W8Pq4wOtmHnjMwivycEllhYe9ZOZ36TaM3W8JkU8dAOsnd7Z9I19ExF5nUuLH5BAU
Na9FhaEKJdIBnHAreSCfWXw/68ICLscTwbwzR39UOFI3eDmWNDv6SuJLUW3KqglpQYRgTVpFAXzT
Hl5yEja2Xs67JwGM15XC3a4VFCltaCSa+XeKgomb5d7990I/S2MgFBviJNNCcz0KpgeWISIWcVC9
S/HGMbNfrxEmhQ16f5jj0PkdbKW/n84gAJiJ3dc7kk39VrM+xHfG+6RD45q8Z7gVLfG79A1+C6qj
J8F8DarR/LgHrAC9aNxxZO0yFRXKXiSl5FGp5ktpfY5fGk+WF4NOpCVWj9sh9s2Vp85rUurU6fiW
+P7C7sgE9YAy0NYP6If7VKn6r2wcK1h9xI/eNIB/rYaaMuypstDCzopAVTM8g2apxFikQ25MHY2E
vof9KMlrXszVsb4u2XFviEAWeS9AfqqZ3KftDEVzmrjXg5c4VdDpuTPgQebGrFsgYDlyiRfs6Wwz
5X7damVdvYoOodSyD6wtFQ2aZMVKjoePkyF/yHqG9uogkHquoYzsge5QYHLanK3LIlsFgb+QHUGS
zcXJYgetQJd8ad7tPT/m1YyoVNGEmmeBzzWxqFD6iZJm74neJnV0SnFD0VP3PjbFrudmgQMEqkM1
YtMak9Bo/dvxpxGLWDYd39EIih5co/OfZfnp+xeNdUjp6dBxzv/NjH5s/CBI5MdzIElNaB3Y//te
hLq2VvkoUfwkTwQf1GEU1QahkRUMVpWtODEDjU4/7515IpAVDjjSSLmjdtCAiRS6+rskU1ANcsIv
+VFYXWBq9HkFPnFUsWJJ6Kafh/Rn0VPz5uqkLcGhJcChmU5oqfgn+V4HUnvUtJt0+gAZY40o1ZWn
bneEQY6lDmlFSkHeJxaQ+OpSSa5Zeb83UIV7bJ9RypbGEv7prD4Wd7oTXypKM8U1SGMgAlpnGnbN
GXpbvwdelQNdpq/8QmjTOfT/g1e5FtVjc2QEhEeLIzKzEMsR4pHBNwWqDTU3xM6CTvrOS5w3wQF+
E3yMn7im/bDZfBiSSfoypJPVo8t/bGCIZk/NrPWYaEn2u52vinhcuyAxGVRoetr8mci+UB8AsA02
CCOCgFb4FjnQnOxU5eSnd6U1wGywhBw4oduy1KYz9Uy/fRpUtNXSiemkTVPF5IgajlyTs6WW0o3H
0ZN0JQka9yKOWJbOLUPH4otVN50Ogx6nDfs4ZoXCKug973uad2UdKyAbLI0m1ZG2/R7DRL6GjePi
bmz6JwqwnvoXv3X2ZAIY0TCXN7/oO9eKmd+TVwMm/+Q+WD3EghTQcg34Amr0HnAXkXx8ZvmrY6Lo
GLD2FXm9qZmdlhLbOM4c1PpLli1rpnoUZGvmJkErDGCYbob+UJmonZjVoxD6UwKEB+2wAapjIPX3
p1yLo300sy09iBBqjd/WsB0YKKnDNcohcmgpLg+scCZUusl2EtCtoVTeQiGijgDbkcBBDdtk8ZAM
veKHIuu3I9C6fkYORmAuamquQmU69uyfIlIZlMtS/on+xxgIdiOuR/BSPw1yDevm5lSN4kfO5Y+R
CpvlWCHW8eAYhnN+2GRWm6E/vornHhFZb6Ms3lyPRAy/5XQtGNh70zO2T683Hd9rQxI2J8EQtSyE
n3CrcOsx7N4NjKa8P7VI1IQg5Kzse4xllb9AEA0mFr8MbKr4WSRk1yVdPxCa5mnvWT3LMoanbI5I
dLEvxsXghdB/dgE62Kq21wP4lNS5mUn5F7FwRKlscdbskXe3DX105/p4wCrDJ8TKupvxcZg6WclM
qtet01iH8Keqke7hm5wWR3FIJia2E4cCBARUWuPjNstZK+bBrazOMoQb/H0+Rscxcne4ShlNZbz4
30RySui/9aNQkg4IOShTe9WouI0FQvKRLu7cX5YSS9ZXsgqoHsnZMBwZeVOaZXx9Dv+O/CUCNYe5
wKKVxZlnJguQOdn/3a5o8rh+Y9mwenAFp2pCJ2yMKfB1L5Wh4/ZlGXatyv//BjMWXCkTCWebEDdr
mrZHvhvw0d0vAbtWOI6KL/+cQH+d1eyHRdwkI4rCnBiTD+LIsOzyNyMXkm7B07Ahu89X2wu5mBcQ
YOY2UnbXMFiPnlQzp9FtFtSISchRrznoJ7yLrUmoauNwViqB69unKJSH7JLZA+OZkzjRZFAtrulS
1hNNamaFv3Nq4PtIl0b3njuJ1mhu45vvgnzMDKT7jFV820oMrfjH6VeKmqUbJQ1dTzVVRwxy49f3
/H+4ktIh7cVe33ALJDe5SklpSMwkrcMw+9PdWrk8IvfAPGrSbtvn2kZFaqkSiQl11oZ2YJor54f0
N/KJVZcByaW6pAVzDViJwrpFLe0lUQrkQMO7itqdEmb3iDmiTLQ1zHxDCDjb13tops9Mdg9jZlhx
5DRaLoa7sBQKJWYLztS/bLDXTNbG7jsnsXLheC63ldI5eORC31aZdFOdXgZM/GsNVHfieMkoUBHe
qmeUvAI9Fxy1K6KotwCtSclEo0G61cLQ4seJnz7C0+DRyHad9r/5ORzx1mLwGxUDU4wIrTCnvGku
JSHiI2aq4zkGSrbyxK1uvY9UVhlT8xyd90MnXFcyznP5+c0UkUvgkmuv48eS4lM/6L0pILV0689r
aMoqRSAGQB7e6QiUZ4jLmJMz0AJZ1qN2FYVM9w6kkCT8FS47lvNm/mGY6adHPp8aPp4qaaojka3S
rkefj9WZsSFm2W+6cnr8slcVdqH2GMPjUM91E6gH1GHfRVHhkN1J0DSGQq8oR5D/HRUNtsx9IF0o
tS0jtmlh8CmcRnwKbVbN4SDY+emuqK/X0Vt8ynBgX6jPdc9WDqa5olub/g4kfWMXWDHe4Uiqm2dO
FIalmymcfQZybl7u22RrMKtIkbK75e0405QxadJwOx95IiR5xB27unrBSSP7cX5J7Dir4tg5zz2I
ZVwjOxE95KK1zu1eF4U+lnJpZ3PHeV6PzEBVWtCDOHFadDPFRU6XZvz4Eim7OrfIuR0nSZPQnHW8
pQNp+GNe5lTiGAO5QXrqg72C4RAp+QRUel4nu2M94F3X0gIwtudblzb+0Oc/OrSfd3f8F3LX2D2i
IqE2wB1SCjr2V4mxyzCNYMjnq84+l4+jot41/Z8RKcDjq93GnF7qeP18PH7veu6kk8sQddBeYfjO
PCdDWMom13Xeqen/JVWtzNoOJ77+iawU7bFP5SO2TFH77jqtwhrEqR1zqaffgHxsYJaHd/i5BNvz
CmED2ATLc1iabUhF19OR20Rv/By9j3Dbnic5yLP5nldmnJh3LclypYxJb+pjbHkTaTOebmJBl3Sr
x1xCXooqsqTLIWlXgUiLjAXMem5u2aYTmarJsIPKoV+mb3cEmy5P2vtl1xxI7q3CxN4wioirwVw6
4JMXe9XG1+RzWVek9dB5JXJhbb3pgTxozEK5YzM6k05Ih7eDBg8qyTnfvuizke40AT7bFpB18M96
ylZZyotkyxjf4NrDGL2wZ3Lfr7vAlBSlk4iErZXZt/J2XwcTXdh+gAKNfvPa3l7uGB+bVd/XtkIG
3FC5l0qh3H+ZA+K1BdW8Gf3GMfEaVjSP8ewOvBgV0cW7foOUOwMRvtXpgVMaZyDInzxcsjrmPIH9
49E/FkP0L46R1e91JI6pp+gK+YBmQgIT/VFqNMwH9wrpb3rhyc6gKprGiSRQRpbAMhiGhQ6ROuUe
Nsu7uazReXj8rdfdbtK8vQaSvKZ/0Zln926CVFDagtxp4WvmS5JRxA+zcdhI6mxT9+P+RlgGyYgK
8mHf3NscMDsI4/wRDxnHunuoAEvLn/qub7WwDmXutxXszDr0FZGIjZ9KMVxd+Qz739APGXOBv2nm
GHi4XjazzbNNAbgbjjlajNuztcQgQofkoq1GAl3wKDS8uEyydKhjChfK9YSLTDDNEfRhEJmfY6Cj
uDv5rxtaFdo+APSa/pbCzPZm4PbixcSnlijiA8dkuAfzqSMN6M0vVpAJpSVY3orPUgr2r5tQ7Wk2
Acv2FhpDSnNYyXnfriaTiQ4J2HRfjrqd67GAoxCXsee6A8dJLS6frunYzc82Jtyw18jehWrmtsz7
bP5lhcwWDDFbbBI5mxt+1eDfYQ16Ve7E+2Pis3/PVKJ0f+VTQ3by86CCaN6nFH8fR5g66jIW8b0P
5WmFSDBy80kfzmenCO5umQQPmTvejDiqZ5UgyXtbQG8C2j+XWxf/dzSDY4SbUn+3uEdwDU1gX4xs
wyJ5NVanqLEOi6fJtmY0gbm069AkyE+/iRvnSqYf+SHdoFUopExq45FPtQ8AxEThg+SOwDEXIBrf
DirEIGhQfV6bNUGaMDt+SABd6LwZW2/ajZutJuZk5k7rwC7KARjzYQ7kT4RDYjYeA6uTUrZn9mt2
vgXQB8+6j/O39rZO7k4Zoyu5v5ahmev/DZ/ratmnYQprInyyzzvLIDFmXNM9+FYUrxZtBjx77/vJ
mLI5LukUi4FmWTxxcfiHNqqyGlmx0eE5g5vzDv9YgHryRKURBCp+4aVTjZGanrvgWpkZLB4atMg2
4QDN90rGNCG+HbmYkTWLQNpYz3UfyHRhl0l4tm8PTXdhacKQJ0f1F4YThiA5vcferS1K4bA9EKJU
gEJ70baVAMITaChS16MEHcohM1viQtrUmh1DfbbJv4Pwebwp5qQbD5XYPR1J7NFoiuPMxZkO3hcq
CdI1xnLtmxH4UrJScqtECptC+J15GBNKN37HMFEPNSC2BG7Sa4IeowAM2Fagz4TSAcW/veU9VzSy
5DlrQYoJBbjO+XhBJC4gYcl0Qj9GvxOEF7cj1QeG1cJImpWP+fujD2kV8LhUABozrpHCr58yZDlB
+PwMHS+Wom3hgUTXEHmO0nm9Nqo/3ghkYrtBVstjgMoWiHOq1huLActc5C4hEsz245KeSBWszUwg
ZG9hupZx8yEbnCi3HYWl0wirjh9jby9mQyCRsili8Iz+ev7UzCrEJJ6QM92XMoDMT9ukdT5kzHUm
XL3dIeZxH6RnWxc+syc8oZA1Mp0qwmbWkNrFxEgtRZqnv+EBzAfe/cvN3nc4471hNC4wVphD6Cck
0DR/wrLZ1lqC5xNje/hGexqroCuWpmfFD8k/N/pIMOHhuMrv/M0rqJ+4L2Qh8BB6DReljChPkaOc
JCjkS8jM8ymVkNQ9L2zweK+DkXQUDk/OCyQ+MTjLjlpdthcP1DwJt3vVQqJDAbBQrZVR00VkaVDM
tVHpjdJ+H9euupN7OCXNN5C3z0pihzI6+2mgM3WMahDcC5WgKsnOSelwb97bXy3OB4gXSeaPtJ73
fOiC1iMvqg2fz2pfnQeuGVsz/iWwWPd6Dv9PsXhHCWAxWHLN87J80igyYE2NczrLii/E95FTSe9g
x0u2gm+bFmtGAd1R3jV9Glv8etLGflT4CxwpXQGAl/kqGgIktwElJmlVmmCDlQmxK3V78HSHCYT6
VseElLfja/y/olv0atqa/mt83P/5HpsODd/n1qbAibu3WgNi1CMfV0tsRPZajEwwZwm8S7Z6V1E4
0JOWoXsZZ8U3mf4ZrHqwDjv3zHWJFHH5cULKUSsoYbU0pNHILMYSC+MQydTtXseDks4T3S7EPddC
vYmZTG74eGfsYUdBwTwLbdRJc/0tSpszIzUSJ3QKUTF3k4a6lWnz82gxXhFj3dQO1QbmmGi0Mlc8
Qmt5Bej7v16WjW07VvLIPO6gbuFU/TvwL4MJDoKQmG37Cl2Myx3bpCHWoMOiokUa08D2LlhIU6uV
9OmLvMBpGPnlprEF9iOYl0MyVYoa6YAM3nj/qyji1G8BKW1v256Ss/qOHnqI5OCeJuW84ty8ahuZ
8UbEz98s5nnf4RROI4T4G6U2+D6zm9MQfmCojfjYgpRsBYVhbJe5rGYj5yz9h5Iv8HqzDKtMB6o/
mgrUzV7y51sXg62jI3lpRMri95RUqgfLNr6OXUI9STs6WJSzb9Qqo4aL9D6sdACN1CbZ8x0iNimW
mXEbUpErYxFu+Eb/REGbBuzFM6B0i0ULIgkfUXgIhZwyoDlIaK1n75im9pTptOfgbkOmWII0KlnF
FzNTwA9lBKqTr7hjIHlEV7Afc6hU0inno9kbdyxGEtpGoU+8rvGk9ngBjwIusYZjxOsJSQ3RjKY9
HISF2RWFlVpw2NLGMBqa9702oTWOvrON4gUgv536vSJF+/4ULkE+pmTlrAhIhEnx8EYYKfuJASXs
tj58ObKo1mBrCh86hZa9uFlS5Ksr8b/hRQC9IWD4fTH7keHwHBQjbRHAAXs4e2Y3+Z/kpo3gYKsZ
bJv4WGF4W+FpffoB6cpo1NDNTFCXW0mE+KU5B85wUiAgaKXR/+C2Q6/aF1U+Sbu+fF2+DeTaPwVz
PSDQREtE9vkyNz3bw1GV/+s+4kk9VeTw2kvOW9qm0VETkeRh2SppYW6tOMPjxm6/cfQyMW6BDJIQ
fdaDNGqjL/xRDavPf5KD/+YVw7vZKu6zfmnG8DVdVsyJH0XERb7Qy5uEy1hBieiEb+uUqY4nMdbV
AXdTPUHwajFyh5oAiWKvgRpq0xC5fEYWEdMD9EFeI70APvB0Hf5EEHl0IVCSBmdZM1zYIQouJyJv
RdI/1TGU9sEg0F2spcqDwCr0lWligwyjE+vR43hPG5SAPASAgDw9rjJzHo35Jo2+XtUS5uOwS5TB
8kNFQEdTLlD4WhNM0cfyHwoo8jQi1mjqSRGdi901OkE2okBnUWRLPJtt3kKEGQMJWPB3xfXee8iH
A2YjLc+ZnFqIHx78kePczUH7O8kzdPNANECH2GCNjnBl03vLeE6AXhm1OyWd1F15zFOB9fLuMgZC
WHgSFH6zSUKykSQlQ/n89+0o0A86d/rJkGIXQe29vlA8GNo+fwwdcFq4o3JwZiu1x+htFt8LiqMV
hn5gXWEEa/N/TxxVeNwvUjBWMmfK2kFrqK/VDup8l2ikfc6C7Hih0iJpWJFH+F2+9C7eSdgHW4zp
sED4UTfjjGXuHNOblNjSi5oxOydlrIcNJAs99ZE42fo7S+NaNdkpHw0ytaV7m5HEPV8lPagLmyXx
d1TdPTcQMSM/wDEwYoxCJg==
`protect end_protected

