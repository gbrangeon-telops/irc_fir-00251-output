

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eRz+leRSRPpou0Iyb6bnhB8hg9kPbBirrzFUAdKqw/be3+N8ZrhDizYaLfXqnwxlgZsSWJCzRfM7
HvMw/rTLhw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rl74r1iJC/bnSjzA+Rx4NZe56NnmjoVRFzUux12uAkwgT++rVuZ0cWQxVSY31Gff9TGn02lNxavo
U1xWF81U2u/Zi0XY7ZHmbpbdUEdpSv9huiEIrpuLuTgWjBSUwsGYqRxHLx1vq4vioRXFlAhPk9JA
iYodwxjKI7YbbZElfVA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lO1ylq105LQ/xiJNZcB3fPTy1RngsQ3yQ/KJ6FM1qs+SoXmUQjQaEb6hJLPAypYN8r4VdJAzSC/U
5nFe27DWNjEKmiIleROkH20okne+9N7+PhPIZQnib521U3SV/ecBImKKPYRpHhAeqE7OE/DzQFWx
10ISqR1I6WBii4R8gkz5k4dkFHhiTU6fgkIHLUXXclJrpQ6fHHlk7MPcpQDjK7bXjIiQ81qfpVmp
P5Kh8wiY7VppUj33GlIcYsNio8GAIV3e0kBKLoX73uDqdvJ/2zBzKOZoDd0As7C4AHF8YSixL0MC
djalIDRCSOBX8Rd9h057rIe8ZIXNMu/BHoKk/g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aJoUzTg4Ju9hNY+ZPcuNUmGg+rCD8aivgSTst8VRB5/g9QHuzghA24ad2z08gxWDFeIOT/HFgT6H
g4nDsyLlbHK2gxUijkJ6ORkRfGOxb8UwHTzLEIRJ5zmkHtJXYM250JOsiukrgEDT40HqdtSgre6O
kXXliGFm9MU0LwRby+I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ca/+TaSll/KHF7mIE37XMZRKDQpSdluwuJA9x/CRPHNmOrubSxRKoPtbXlxVM6ehE2hXp6yB6qBf
Fup9ZI873BFwgulDsuQHuOSUPGo4bBHwDnNbSi/4G2je8uxqj4KeP/bv0RKunNMT/FTascQdDh6n
SVSARZi75+ElUvhBfAjPHB+yugMvSxDk7TRPn1RomvNtW1CJTL51/PQt26FoAtnxmwYDcU5wo8WT
ATzZmP4jq9ClSvjXHkf/VnlLenBFunDj22Ef6vdvxByXWMZrDdZyqqIvDvktra69BBPdtD2LNyW1
FCI6v17qDRdmShLAB1bJHs4PPkDtQbDOwcgx6g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5040)
`protect data_block
HkblEnvGvLY8iROl0hW/Fx9ykLwuXP+pqo9EfNtoshoJAkNBqU+F4za/GdIJwcI/GUiEQh+L+FhG
yLpc6T1x7z6hH7qS0KseSY26i97BCCirElRv0Sh5WQKYGD73UAzWtHpKrsW/SahyHCSBMSAPRIJT
HKHGmlARXMXaZPxoWkAg1FkZc2aiM2wK4JybVurCcB9HOOA/3rhw5rkD4AitShg22PGpuzbnepMN
ynhcVhgOxdUkSgUrOR2t6lmg/Xvi6da1RQHqiuZx7sY+8uQbP3xIBgw1Jj1Qe61bXQibykLeqjBP
+1sbtv84IkrdIU50MC4vnYGWt2mkTk+Q88iVAzVvNP+69LTPPGbK5aueR4YqoxQPp49KOVA906XF
9qc8CnUOAcBD/+YkEuO16My8EC07yhx4Lf0mhyYPqk38QhCzPvu/tsVjQ9KflXGkgqwz2mgoW+oA
/vDImdqX2mfNN+/KXcjV0rAnmRbZsI1U3+iZE/imQqTHvFDWO+D2mwYARsGhSKjDMQ1czAr9lonG
K2ZHmRS/GNL6z9PcKYjZgqxPyHJLcb42xhZo/fNi9kj/vgkFY15zvWQMLTdpHhX8kOVFuCoT1mjT
9l9/rcyHq5TaRcv7vueYPMaqEUzn0hLn8fNqAhapNjuvmz2HVEN0fsOrYSJFF0wxh5rlFVKjeiMD
fQOfqESNkRXrc7//NPfHVpl+NrIAzJSYK++bDhgRO5yLIWGdDSjzrLFjJ+QwY91NKZsLuoWjafJ1
mmKdxFXLLMx5yotBVsoeYAJTxqDeVNa9KqXS49ouJ0ay8GnXl5zNe2WhnAvngWOM6eH7GH2CFl6T
rq8GNXODuJT4X8fYnj4GYceCSe6ZKRXRAzK99gmS+C3U8+UTQ5A1lFH+ZSCOJNISujztx6JAXkb9
FoDI/hoTitL9JszZ9ERxx84Y8iWvQyZXP7Wh7mtMUMsuLtuJbV3YuyHysaaVZUMwNJ1hvtTxgGif
NyAWWaE1GPHejEeXz5Yq0ZSUHVbbe3zh0iPlolwmxJiX52Ml2nUOGzm/lFYEG0lAPZj3/hGxRXCi
sklVfgjppjwDETPtRlda08R9gnFu7Ef33TJn863wsxnM8RfJT+vF1GtGFl/MJnNLTqWgtF4+iEQ2
IQdkXBn72LPoqV/5r0rm/GS0KBy2NxiwiiXfZ3LUZG/WqVnuCBQrTMPmHkHjsofaxJRuEyxGb5BQ
+InMEoT0wI43IIvLiF+KaTMK4/zR9GGs/k94Oal7g1TZU7snGwi9bRxa2lvwf0UtL5xT9uwtaxG+
1FxQJyEVBs3WWNAMkh2QqvrjfdQ2nRkt5lj8BNeQzMCE9F140XUBg2t116knD0R2DFD27xc6Tr5b
83oyd6KxKA8gb6+NremVw/2p3qBWG/Zjuz5DOzvlKq1q2BoJCXhwaO1XomUajVa0HacBvdgqGpDt
s65BeCPmG6IxbM891G2L8DlWusoXuKIRBpezTJCyT5wFRxw+GGp6inMR2p1XHiqTO+fHrLyKPAqm
ECmJGUNbIzBlnYIp7KX+wVaxLDkLPDBlJzxWyt4HdzN1H43iciAq6XgNlWfavRaHBWfrOruqOSrc
HVIN1TvIq1r2AVK+OKGVxf/mg83gpjwBIhtKGDFyaRCNwL3mZHfoqkPX6Q7ZpkTk4OEH+RDHRgfr
+a/ijnwYf0jCHOU5KdbTHeC5uUOUgFth4r8Chr6ZKMiZJw6ztvQTalnrbuKGqC1l8FfVhJXqUs1i
5SYhEK2SgfaTQ42xfLHu/sQzLqfvBHgT9cICvzAt6915JlGltY+LfB8GvrK1DTXVFI4kmbSH4kxv
yRzWZl43J2WYSceNdMxRurwX9cYOAKa/KT79W8PGINFVK/G3EMLmzsbWRasWxg36fgoU3MmbB7sh
x5dtyKaaEWN4rfrLCWodV62x+wZWgiJklFz3CeiCo2XHI4Z4hyViTlz6ep4sknx73Rs7DykYsUoC
YJMAK6kWya89zX4EhCJvUjozuv4xgcz76D8NfpSylmTw6tmbUktmgGD05k+hTufbUZp2o/NmaciL
VU5Es7Da7tubaN93KcICgEo8LSY5NYqSmeNSdam7LcSOj5j56cPp2xXqTs74o9FGmmDPzntfZnhd
Xgk8EWOpAs6yiyV6yYTmgP5AhlAI6rBlaemHhLZ+FONx+OzCwo01ngR+EYZ/6gqnCxeP1fVrGQAo
hyyy8R+P5hZu535WhAWp3T8YEX+KoBfQ5diu3jc7YneA1cKwxT9F77yWyOzi9k4HwcJZTcfRTc8k
3ts+6PNGySmXsXVywAk2EBJ70CU9LcwlOPaxylXljxRs286SbxRV782PPeivs7xcoZiMdAzykoMV
A6QY4QOMAdwBKy6LAoWdwvMzTAOlpYy/mgpqogYqPCCBm7Vj1iBjfIcEIEnbqmaPjtjDvzYqsXKr
Zv80fV91GKmYTYNThs6hfFLlhtu/8JBPeo12bj/XPB6ZPi+Keg8s7ztWSDXF1bzbs7S2QyzEW12w
aGeNAP6q3iMmYxYD59RFCPkW+vtkYeshinITxpuLN/rYKYjkCf08KpLrpzf4jEBDUanaq67LuDXK
aVZG5EqTqrJYnbE5PaG5EocQ7U8oOdkVoET45LmjFnc/5wJ5eoLPQwRiWDzaTq1c9fJNIFqYoZjh
TxLbSZ0R9eRdR6Q/gVlYNr3iEmRVHNlYvRkn5uXNS2drlgVbGyb7GynMxi1O3JRpf6s32Ah/Zkrs
cpaMgXX1TVN+QBPn6AV7CBNx7oe26WDP9gqc5UFUeUf6eGQ0IQUZX7rbcP40YazSIzT/bTAjh8Ty
Twvnj30xz+o0hbpfpM3cmUsYekkitNy8y0EdY5TF9mvZ0vlbLsdRZff2FOv+2ze9JX+aSlIblwUV
lFzvKJ4vEUFqRy/I+PmZCtEZGumX8FPOVOD8lvCnrI8Z0CGVSgoo8qIPZubc0/cnu9Xk0I7WcU6S
FKcH+/zSfFadpF1fjIXboPOXRMlm6bjugoxnaCNrcSr7BhiG0YZy1c0XVYaX+mwDxChraoAp+ne0
bfCPsXbvzS3461I0leDHQ3gtq1Jvzcer6NGSdB8Hw698CA1JQbIqUJGxr6+9gy+L5fM66Lm+pAks
Q8bMqCwXGU+xbreALIilWpC/VXYeuubwdOZi15/mfv4PKya6AMEQtVZqBGEKYpIwUJdYrlJuMelp
lTHNVfvcYoO2tHE9S9hva7LhNJNF+WpRqr8sFvpI/4zPiPSUhJHk1hNfxvkBllWVXtc6BmKn36Fx
AkAJGFrocKr/pZktBuGTXb2myGuClNVCS1o5gvLGzbZ9Z0YMrHNhdOANqkYz38uiYlOketgyzDZ4
sJLJFBIXoqsWVn9pCiFwFzSOVWL3jMknfXiNI3tHlbBQqJiezZAOmHcwT+Z09eMQi/LBDxJk14C2
jY4YbbkwSXQgWj22dJXUjKd1sXOLPkAhEovcPezV9jL3lx3kKBkRCuAG1np7f85ZDkn9v2huNie8
Z6LcP39DifcoZdIhcpADb08+nZbQGEIAsgvmdUi7xlJvmxLrUsm5SC4SB0mTulyfBrXc3pz4ktQ4
ANKOdNTInC4eviaPmzRXMTm6bNN6yN7/EqHYaKv0r7tSo5lp0BTr0e1C0eD1wxaT5/CQsQMO/v4L
DYdVVExCKON+YHJluq0ri1YNFyP4RO6a5ZqdfnckK+XdLNbx3wpfjR8z3hq2UX+TOo4p8y73SSWI
of+BM26QpQJN0ikwY7yZDa8C4R4guOGP0+DryXVvF0XfFqXIjJL0oJyM1XYABQbUss1HZBXNUO93
fbg2nkB08Uh8SRoBKA1/mZI2Jl2OxqknYFnqB+aWFWC3VkN0fhkjY380szqbfR0xCiqUayALTNrN
+zlRSq3tbHUSKy6qeyEavIm89RmSD6H1x6+t8fWNyqrYUH3PrdSpKkdXGGHK9DsI6k5iiAcgAd6y
neOsuKhAPFmXAf+uWOYHg+/DLneh+7PbL2bYUyU4wtWaSBjx451ajHNlP2uznX/FaFi2w2Lu0vBj
nHmGT2fuJw7cLCAhUFP8HIqLzTMee2YelYipjzcw8xML5n0sR6BfNg/ILZSnm7+Mo7ZqwFKCuYlz
+/j16gBPVPomyqQVxAKCwwafELpctIl+9tJ60dtdvZBhuaiPyrGLBnj8XhzF8ivMyirJ1Wzb8hhc
pd8C6G42S+8YXATe9QvSFcFiWe3k7mkgylfULo5jaadIjPO5Iin55nSC8UVItWPo8maFK4DmHW/J
/fFNA+7SGN3hHHDvlFObRmVAg7osTNY0wKueHDAEZPNstG+2N3LI0nTap9eXxWiQ7OvSAvlocU1o
pDKeldmIcNX07j09VrwW37ZJHTwxEjL7TqxkQUJ19McLjFNDYRMoxPkfDDbngJZHd1mC2byMpGlw
uR7kSTOtgefbwAti4jNdzmWwVOH7KrjCd9HTsKsrrFugutsHqKHaHqJew11FhNEhlxCVh1fCJERr
yJWSIu0ADlGr9kj0R3Jq+B1sKAqZSVArHdH7bHNVnu0zEDV37Oj5/T1/wqQ3+T0ecgrunHUFGfkP
p6JdB7pf1b+L7aMblyVKKs8x5iO5WkwPoz6dkntzZUCoQScKeSnXpWpP7kCdX9HDkAJcZI4LgX7L
IZTb74Uo65hfX5U4ijZpIx8Vo+63ZiOmvwb12gfyPwG3lYaTlvfLPf6My1yIFA9AHdAfCC7vzNKv
mblXkscplf3U6CL2+2ISAlhoPQi3293d5FYTQoKP/9t9afFZprhntkppyJj86wGuHD0r19FGJCrG
JbwqWazI/CyJ1Rh9iiY8fCmgxC6RKwlcMJm7on5BHOSg94m9rsHku62wXkcM32liFc27sQtfop3o
UsIJIDq+DsqoVwxCTgHtEgv+2Jth6UKV5sJQXVqV29U/OV3g08zWMmC/CWApqc1f47l+rdxcQKG2
qcgIzXjhgY5ItP5ZI0Lu/b3mrJAn/lunNYO+fO2rhNRxo98mAfJ0OfkkEcHV8csNRfy0oAogGNR7
tAV75WmfPSH7CGYpN/L+X9CCJJwaTgENrjJai+XIdB5XfffoJXsAe2jdWB4IrA87DeqKWp7kKzfP
WGa3CS/8cvP7QZtHXXvtv9WeY71jmzXugCO6yDmfSchegjMVcJ+mKX95EAsMZGYnywUxFccQPvDw
vq6KRihb9zqkMc1EhNVBnUuvwSoC/sP9RzWoBlhvKUQlROTEFHlGUKk4bvljh2MywO2eRLIqqSTy
sfpmhVgpnZqIjm8ZbDjV3UCg4RWyhA1qi2SziNFX8NImqKkwIHWVtYl+oGFMMCRRhRF9bWkMQG2l
5Kiw8bQ9MYWOpu6Go0KbYdCxqEer+3wnxhpTu7QGmnBM2NHYbO1+dMYMN+buvRgVGTx/oTWw6M0g
DImf6ONgYsAFJV7Vj0LgwM9GUJo/1o66eyEB4ezGb+38uuOUBRqU58J1VSIe+Mu+GZFpma5q2tfq
idblzNEDHvqw5eEKLK/VutlzURSiwcNHTF2U2MhY5f3taHGdh8l7E8YcWEGHpldX93SJfi949MCu
3Ld3MPWvJO/dhBCwnpqsLZKngS9mP5vE/QirqYLSye7I3kYkc5H5xcFZQhgGiPtzkGAUmVjaP091
g4TQSKayPpgkqK7quX1w3BZ3Xymj1ycFYd6ng9/O861zQPxtAAGJjcNO/QFw0xG4HYxgewz2yWCM
cL8uEMbJ8CnME4VDWni5VYwOYqfr1pV6jQYMhxqLfuUyXDnN4dtFSsD97Yiy0wE2SpkEdOQSskAt
0LJyjNKfNQDvjMTiAqygxD/ScLCrpqJi+MUJulX8xjgSdMhMreMs0uQrnL4hNEYnS037pHvEhf7B
seqY77DVByMcktIAwULMyw8WZODxX9Qtf8Syfn+3e7Zm/UcmOwwUSp4ZGeTvbBvtWhPTjKvGmUyH
6JvrF3QgTPODYkPNFp54De4iRCfSu8ZAqTKLv2q7AcaMga8oQiqbtYGER56gcwC81NoC72HCFIPU
OJLtH01Ez9sq93CqFTs+qJQZL21Gq8yxQD8DzsdxprSq9WtqG/FiBsFUTo1o1FSJfPGxyivYDwOe
QLCMeq/Fd8T0G4VWWCgSwJLz+6uCfTEUf+QxDm6C2F92eMbeaOXbjJbSEURslK1RRI+IYNkrKU3q
BRiD0WjMB+w9SfnpyLLQUEdnACn/kpFDnrFCMsjM1ApE5rTfZljkNi7EaGBIabRE1ghJIRr22Lvx
H2HGaFQJZkBCa/K7raC1HUvD+5Pqx1NbgaxlF5c7YmsLZMYuPpuuqQYgDmz0Kob3zKAcuI11iZJI
142G/QzGYMD6nilnZvQlUOKCEcd2NTzzqAFePyqZpJ5nbPDRFYunXzGfCrL/pue20O+H8Ln2LAqo
IseslFuinE3hTXL5WnqrexE5MvW1cj7P/Op6ufG+sCntOYuHRq/gCh2JnXXJYVi1Kc4XnEGHSm9y
W+RyZQb0nh0yNo5LYCv+bAaocap6mG6NyAaLnwfDzEPEuPc0Eb3Ox/ZLVo+iLDs+4kGHWdyMV1N2
rzU+ShzQ+up3aOi7OvPZTWfyI+VQl6OaSg3NPta1SQvrP6JSie0ZuhmGPIm+TngbyP2YUJHdOlXy
1ItskyiUMBUHHyByXwbvCh4viMAQiAQH2VIJHlloAG5SxiLNa5j4dMQlz72omlMkQxyoqAaRwsXc
O9ngzYaU3YbG/oSZ1EMrRhE9lqaf1KUW
`protect end_protected

