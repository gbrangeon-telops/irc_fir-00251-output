

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mwxNacl66MFUVIMc1Encct2aHZOcb2pREujQa4vWHOpoY4Ryx1q0qOlrkehqJnJB6VdIGpRZ75ar
fafQO/Fcyg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WTY81lfpic8wiNg2xUTFY/9pIQI3CKsiY3j1Z19a6adif1iCy2STS25TLTe/dZhZiWj1W1FKdbVN
mTJAkstRD1IiixRw4XPUhHS0kg8DebELiBmCxBLwbMicqplV5b6X9QbZ+d65v5AnURtcySKvK9fO
g9n8up28DiiTZN5JTCs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wSJmxWNG9Vaz0hV3ma6xxbW6Q/tt4VebLF5ALUnEWrb0oMwD9MOvKTVg9bgiL2D83XqOs88TpeXX
Ifg7m/wa0qnVENMQDpzrbdsY0X541kchr6nHO22IjxAZU0y34IzPOD4wlt/LkBIeRhuE2oOUmiUB
mj42HGuDYM+OLJ75MJFObfMegkawW+dQ5MXJZAvaZb3Gdq+Nc//x1D0rUYdDzCYkIE6Z7scW8Wik
/MJTbyzmOPOK9ZoDJMjaYzyR5QyLAdSzLEdKbGH7TxDHRl54Q3XCa50pfJuN0PstSuaixGzvKQtH
Tl8qJKpy3o7KeFGSzvILj3NDt+zm7na/fYnOyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TWs0qYIcIilONYk/cz99Kwd1RIRPFnNZwYyu+ici+iMJ2JCkq8jieFKJjspKJpdZ8Nc8B4CnG4qj
aN9KKPyGY83yGWxxRkXLLk1fDABMFcSV/QWTMe6VkTZV7rSzb+eWC79VK61VEPbjbvhhwl9UlHat
EKGcZET/5AsZpsdS5rY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J9Mi5TzDBer7RNgnQmNNaMr/oObsCpVjypskaWXDXbsUL9Tz8WTWA1k8rjWfCv9Dmq2LFoNWohyz
5PixLjvzdMk+0EAtGJRSdyjvZnuW2bmu6ekaURxk6HvWMfHmukxtVO9c/su/PcWlhTBaWmQfDEOk
MXt2eXdYnsY9DHX2xUQnYdQty3UwLIiL21L3I3SO1yyv2PefA4p4KfovFGDUvBPco1deVqNYRLx4
GphEA4vKS+OANoIaExoVeJSpvDGH50O+wbHahIOE11SE2zucQ8cWichU4yUJXYALRvrOZArC8ClG
ouWj0ts+fBWmUc+Q65XK9XqQ174/nPdN3w6Fsg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38784)
`protect data_block
e1whfMM14J07py8FuEEh2OOw09gZhV/rdsg2GCcVpXEp1dbFDuZaVs/xgM67AMssCjATQNlVW8Vd
PKhtckebMcrQBmwOkbwCDt33kDaVV1TIcp2pVrwMrBnbQ5ADKB9M2KtCKPKSOKp1JVTUyeEK2dF9
c1AFWsLZ4shSchwGPJbHVzPcnAto+8PZCGxowXZEpp28KCX2YHyH4tSuhUuDza1HMyKxQgSx43jn
ikGycQINa/cbSNqPhVjzPitHAoIes4BgwvkkZC+2yX8VybCgv1Vo6a+nu3Q7zh4qH7FEHAtlZpB/
OeKKRymjox/y3KKuQyf98kjNlv9DafFzFIKt+AmqbidZL1CHe01rwJECkzpfedOqxmQAGGhxHkzn
cnD2YgTVqqc0l5gTbCdMZZ1ck692zUXTs7DtSPBydA8Vl8QO1kkGy+44g0MSE4NYltKYk3XsrCXD
4Gq9PUzXHzFX87bEgH/Yr2RrjKyNLWaS7fqZ1MY0Y1ovCbg7RFDX+HQEUKMvSmdNk2Pn87ltnDXC
GhWhUUkmdRZ7RzkIploSKPQBu17WR5zcTuphFNR5esvY82ulGIGTQj7gYTS54/XeQnp9Eem7ajsR
67z+jYGIC43PCD6dZ9m0kV6QWsd1v7eeoU51r2xIO4EitSiHdNLLWWMZj4b9tNtygoTzwrZbTlvS
HBzUkWskxpWMSttIJcqjmC5oi+boiURfyTjlkJWZOc6pKnArwzcJycVTVEjCsWNGoTC4WKe6wEZ4
bjh5EVlA2qXEUrD8IyBbJigMD3X3IXlK1gfs2kGJnmvjlBL8CxxYGoEg3oMzbGWb5IHkbSTazBP1
8T4WX5liwNV2OLSpKIaLCJp/SaaK3UJgvdR9QV33bdmvOSsfYhBPRpuOclCqLM7nu2RLN+LEWO4t
sxYUJ1mkhQaL2Co/XKDcSAZzaTohPs96mOjtZc+bB4pM5DV029bt6lwq5ZIhSkXS7s83FANfcTgl
RHWQs8LNYTug/MwVPmwJoif1U9JvNKOBqkbD5o5rUPFP39aP+XsxDX2kuj6oLHfY7+D12dJTQtUh
qii0mmJ4ss//pepdtTGtJN1dVgQOuBA6sWWxA5fx2uQIJUUgw3uwl4+6bmggBavOP/x7v6OjC36A
gA8eKcGZ2iW3WUc5gTPtyEjrDA+S+9uOSWMRVD4eOJndGDBOTUXKS/pZW32nIlFVfvhMTPDOcM93
u6pMSxacIhv1iVIbaOKzEHvQupTPeJwv4uz+UGeTwPUxKzRvX965W7zp5oyEMzg9NTZMGVyOnKXy
HbGKlKC0/x2LqzdWZBmTCifXaLQOAahsrBcc4mutD8J1fA7oaHOte6IYeSKs1Z3SItH1MSwxy+uu
s9lVjyAo5cPk/CK98EaPbdHBE4epArot3UlCU/T0lB0IlteltDDJ+vtNnFwaQLuIIOac6X0tCn+x
T4Kp096J40CQhMcAppDdCcNqEeqQ3EZqE8dLXz0oRSz2KZQMkk8jeN8mDEOU/Ow2Gl0ammhNMzFC
tCzlGIMgpWQ1iwiWVku4TyD46nT7fzVZHU1o8GA5VYpDzM9QxHyTGuQwAbjgzD/Y9VS/xShMgi4/
RXlrc96ysnxeXIkn8b7Uq2Xx676C29dgbe1xnW7+sxMtdgXSYT109fJ+bCwOu4iMZ6K3rLAPDTWI
5E4/UC5f5vJbVHyt/1x/wyAqyueQ8szkavwZbhGEcYY/fXzA9NT+Yb4U8f8EM5Q9CZ8Ry8eo2Fea
Oozv/a4okrHRlTOVcsBYFAgSsZsUfLnhBHci/B4+g7WMKBK2ArOiYQ/ixIS1wWTO6Lroy7RXDEtw
ws9indEOAe7COoO7fgyD9KEGjCdeuLOSxYD8JBxGxm7B9KgdW0vDDYeQU0AEZBjdRZ5YxRZh9CPs
njOwH/3cVVediIWv3gL2BP1+eCfHJ0Z0guSGC0psROMFsKYbKVegvJU4tghiPYJxfvlmqIMskL6A
2syM0+5adLptSy9JEb2zkAgaaNDxTANtFT0f/Jmtt2zgDnUNq+4fRAxkFlX7wFEDbHd4ChN+8amw
9HLQ61enQbmHIzwQDk/jC3Kx0XiFjXAeKyyv71hWpysFRruBqgvGQlwHdQ6d9MsTKttYpe1V3Azh
wYiaSId3EVGu6LNktMmnIzEGLpSLnfYPp5sSaAnxMd1/w3mU1Gzm46bcqN7jEDIvsX3/TuV/G5o/
fEDs4UeGPhM3lrNBET45V2IgjyFkzkMSPQ0zXLckm0nRiPkTTdocwMO7agKqQ3qo0njk/YjAF1oN
Ce7akvPrIoYpFDq8J8zw8OUV+mMgeUfuJWV49VoNgFE4oITHLHuXIgbLkt9TgmJOPTlE44uXms8P
yBLMdmzgPWJBMw57IFgi8N17fQGr8dEY7KMVm0QnGuSIjD90QeUFjpHQn+hnmg5pg5MkPElao/tv
DPwbQZYABbwgvYrRONpfnbEkQHmi6uBT6ZaxMp4fjk4tJh+0EEjJVgF9fYhMvahkb76dT6llDPt3
A0fYzZrzqXTLeDITVJrppwmDkJxDKyrKj/hnGSnh+07SFYV4a1nu+K3nQG4WjWJSHqF911AUnzd7
xxc3r8l9vswKpBncBo9/JlmNhlUIo6zR1C7nYRMsdfeR4ediuuxQXLxT8E0hNMubk88FE3Pfdr0x
Tyi4wshxOuH0kenyRsigjnksRnCTTmUtl+IHmbDzWuO16ycwFnsZww7OtMqrxqwBDH1e+/BaYCX3
ekemPWpYjwPdbpahTLLF8beVWlZ+Th4+hPMkp2zmKqkEP1BO90IoQXjyzrFo5Qu8zNVRCaW/Utk9
ody9R2NL/E5PMdbqA5G8bA/e/EIzcJD7XOjObX/CI6Jon6+yrnKPbABxTxx49d5qK4TcG1fXC5Vh
s0QVFEt603ifjwDxNvlZ9hNuxWbEX079KMJ2VcDe2f8W9CvCagMS+shec3UuSgKq2E8ugQWIxjDP
EnJrSTpiggDj5TPbMGfjfB+9wevclFKY1NAlSXoyBN5zTlyyr7MEjR6VXw17ILDBnw5mHvnR3Mtv
Im4keRDOd3STXVg7bKqH+SVW7gjQrP3HtHJz9BQd6/b+wTlSqR8q9FJ7Cs+7+Sy+0/cBzy1rGKXB
OkyZQx2+EIMhra2ne1whUcXUMD/P4mS+uQjfPV5vVVAfAe7HCQJUyEl83bK1rZEHetShz3DbEVfT
sdxAosDecaXk+N8dS0b3QCl4bVIW1KxKpr1akJMKJRBjrVtrWt0UNsZyulWDNGVk/vW1wamX32Wy
jkDfW6+ItrVwUvPgggzJDBNMZZUUJV5hkwSdpHt0LrsFz827MDkhk3ECbn8Oys0Wf63Uvk0OmHMs
rvHioWqEcEIlMyL5UzCOCDQ9/hiLKXTlqd9mBDLUavzC/xK8WgIIbXcdjK48s9NcqIIyXSfAr/v3
zZxK2Qu5J8jaHTL/JsmZsSoXKDniNXgUhF4e3qKRzv7kJbmfreg/2rqhFUhW1fK5CFf8AGmNcDBC
QfwnalAZNLM5j9nyaYmONOQ2b1ZkantuOCz53NNIwyQ32aCfefr1jvaLPU9Tx1bROJgdm3zbI3Vu
Ra2DHH26a24n/coWyBuJoT+O4WoM1uDZ4eKywAhsgPUqm8vXJJ6uvlWSMBDPtWvaC1Bf2eoJsXPb
blXrP3agY9EWgso4LYkL4usZB958cOau0AkcxRx8DCIwpyVU3qT7OlKfheoPWrIcWQKJPXAOYx44
Ms9Lz6cMPsqL17jmHisWR+sw2uSvGnQV/PR50ahr+8mAB6GrTrKy/1Ft4icQu59caE41tMsi2t90
AmgsfEPneBSoiG02bc1ZheiafqvFwR6GjYqi1zLZz6GOvd3cDitkLKLCFCceCOXWa+P/EBJQnlF1
ZXY/GrTcriwb9V39X7bYyMez346NR99ImsuNLU1WcT8Me9xt6U23AYYWMOR7UfCOJrM8MEUyAUi0
zMEYWstHO5nP04zX6T6svmRM8t6DfDlipv57rXfyQO05EPRLodvelk9TmYPibHWkDFwYOfIIwBQE
yMmNsvncHHpUo/5I99JTrzLAM/o18xhJuyXKCSLkd8jPQFJPsMU5qMbnHfNKu8Ard53Vbb9JgRb8
Lr7xElSPhLDSNrQZi4goKCOYERRluX90ydoNEGPlTZboDntcdYyHLz3ka5fLCI+h9RXeAnmHv+pK
oDYBEtCElwNwwGrEIBPHIkx1wQi+C2yDNgjIx/Iq80rN3KC6uklcgSOigNryjJGmhHeni+Hx5Lm9
N6dico8/+gRxX1V42Dy2x9jyHlaz3gw8i8QAIDdXcS5G2HW6/dcQkLrP4AAMn9C/PQz+hDF7Bffn
o9cQReyoR1qF8wzMwowg3rAMHYRWxGvkcMTSqQliMxKt7norD4A3mVFsbqByH0DQX2j5SQNPtgBw
/1bZL1xRXL7NwopRc4ypRVVwEYJQj7Y1kM+nxxFOykbVZzVV525VHEfMUBXst7dBC7SrnxSkL6tJ
Vx9qp9asEm+U9OZNJKvo2rHSm1gVe2DZln7kABWFW3pJo4MSe1gJAmMDbow7GJuLY+gTVt76FiUd
ciTiQ1/sakq+aIakaG2VQy9i6W01Rbp/EM4nSotJ3tQUVTsGO7M/0gVKxaExGiPOLKfuIcWFIUgC
zvYBgFWJshRLYiK0BNMLG/33VI2DNhAenICHjJKFAqueJMjVJrF6ctnYloLNNl6PUWz5SIWl2eJF
Iu30pUROl+F4ap+Qqxcti89/sYP9UYL3XApPo7TWmShj9PAnTmXyRAdcn/AL5Mbmhqbpl3v791Cu
ZQ5cDBsNhdqsTiA42mUQJ/uwve6iZXDB1TGK2zXVcjE6B0DRhGDU7xlVOqeluk8dwU2oHKqnIEAg
xjl6T4jtmGzu8j96R7zEEFMfOWRIe0ixGRhgtbeahC4WwejauEOXXd5CFwVM0vv5e8LeelaswoFC
6HF7+C4Tvi4GgPo0uMCt731xiMqRfSq9ugk7FuLI6gBfU/7n74cGHAxUdw19F/5Nqjc+V4rQKOAc
4ci02fom2BbkUWz7+3cPH6rdqnClO8ZdyT5/ahvtq+e+sgQabxnuvhbSMw41wy0guk/dWkqTdJim
pFKQ1fBzRz6xXEYJ1xAn+d/Hc1g0IAw88lspPsFgUQKKu+yQjgeeN9edGgzjg0CEy7p6Jn1+Pj4S
lJbKjHMf0JcwAK0CrLBvuNY3YBhDZc+HX3rfeBczSnftTJIJW9xranBs4+0q8sWqpzT813Vw2ULF
5vuF7Da+Sp4ssY5wunA/yFJhjFsXa75Xrm7H2A1mg8fye8Btkls1HHr4PPEr3JXnjmUuHVLXUDFa
GR2qCmvREp+1IEVhtD1sQK5YcLfM5kPuKCtMKfOj4ZFE9HUFUiv0Y9OqlAM18posQgti+IFr00a3
CgYaku0wauq8oTvgBmNpB7cVgFjqntcqX+iox9Tvgnnpt734ogFc4d+BIEHyBqlSPHOXx3TUa4OU
xybkFhW2/GEokjkudKg5qJzCn4XK28OtOkHXuM+8kO9QlOAHpqR5gANmVeGVelVlwpBQGLd7lkLN
Y+ARQQ6oqbxlFfT/RwLDkB2e+RfiqEeKpUbhqwj0WQyIeyWSL2ZyiuqC34reEvaNtm9QdjfIFOIm
SO7bpuH4LBv6+lH6vgRiN4teEU2d/ReA6omJZkP2D62/rHEqyCKAObeXIMYE4NysoRN3uNx/3jyu
qngIXcSjnRxmiA629jo0ZmDcwyjkDLo0U47oY0OwDcQoWPQ6lN09nd81lvkFOcbpdQehSKSKHeuV
5JUWnRdMKqxoxDWExFQxaDGxN9iKeuo7sdgIAit1kBYPKIbv+7o0oWnBPXvfVHAiAeKvqk0kNLdt
rZqlE2ARloEmq26IjFOzTdkQTuOzInvZaXFI1S9bO76evZbSxOUfayjP8vcuobAROausC9qPqwVu
xTz0+age2JZh6EusmELm2v+ZzMADVu2Vu9hXZmfQELcKXBozbYlD9wv0AV0kjEpIaMzoykkN7rx8
2P/y6bQxFE1H3JiL00X9cvMNYzt4/xHdiIjYzNVsscyIdUv+Ge9MOou+hy6OL3NYL3SrOeQFVRr2
rTFunoC7D9clGlkNcYeaL1k9hJmb6hMpmDF4OZRe5A60TOl4Hrhoq10MXEkj1AkS+JAMLOWYCqjt
IfHGsdgQ2OO5hCzMty/ELBem4gB0r0oQIeiW0yaAcFVpMAawVBcxLkUdrbXdgbAqqiSKM1KnBTGf
J4FP234pLIwkQD4MQ/JlEhub2RBhEkgOGwOwpJ/lz70RZaY2L6Uco7gfpeUulgXnOPESrb9BlFqb
LjJdpTCDfbbyk5kykPASS9VLzQfp37V/D0dK6qesFgFdeSPpBaICPxG741Mcfn7j7bpWcz2wMFfS
B5sxZfnNU8NH5BI5ONufCX3vwbYu1dOhMohls+GLWCDnraHxScjfHidUzGz0Ux5HeOdgmELc7V+7
cKw9qTf7VnZJpbk9deBHfxFiD8gobrLL4WLwE8sB12JvJopv9GTCUyOY1EI+Zx3YpNzRZzfVOaxj
JZZ/ns9COz9C/t8nkRhO8r50+57gi+W9vOKl3e9Nx0sNrIZVSNH5BF/DNVxoBFcCD8XmeSD/r++h
qEIczZSRvBETwx0QhhXWmauJ21+ZLll+vltpYQoTdUDk6+WDQrVKkx4sjrVh9idWAU72G5U1UE+l
fikXExmbKoXdbmnYIR9PA1X3vRuXywryye+yw4vz9pNvlx2c+CGbvJTHe3gBJ5Mqj3KGVYHnE0RC
wUy9FT2WyR39eTWWdXfPJk6I0BgWSeW+dF7Y7TxSWuX8GYjH6IhWYiIt7xM7vx4zAVmMwKRBy1AV
jVN1IKudJCnW4YXw+ZMfO6ZCpp9Ehry76/+kEaUU2MQ3Di8URpspGtHSTlYcXOEX3Pkul6y269NW
Nh9JPto3VvdIz+YuYr4PejUZPQopsbsxyN5b3wCgGLlkcOocb8dIRSOxUHGttJtSFlkVB3k3//BZ
WQKZ3rs3tvhDCUTC+hlqUUoPI2BV7tu3twqf+JSbdaa1IPkYWTRYdOujH64o7S6gGBYRoM7paR4j
McApwwmwOC3vVTb0RHcqvG5hvpXjVvxQNi1cOoZsytOIblmissHWV6SzW8/31qzJkcdaCCFQXrZX
JecXdpEoIXFWYHyo8Ell7Wtj65JBFDIPO0ynWTrx3lZJZ4viEB8NLNvjvbWFeNhXXPbBeD7w4WD4
qKf4zNsiBbO4jHc8P4k0IEYKDdXHgjNGLPFcZvYvoUAKHKEQVkukwYgHDjXINr27NCdwR7Ku3NZU
Tax///X95ZZBOs+PZ248b9e0AO+338pmqr3d7RFetZ005fe71MR112hc4PjEPiUrV83JyzpFZ8vn
ZRzJxm6x0N+VUxrsWvQE3E0ptj1Bmp1EXCF30BAvj78jC7u7k4QUdDYIlGvbNTOkDoi7MgJ0LzAN
f+WTmH9uNG6i8EilbfQ9VHD2AM/uUIyBR+rMH5DTQzIaIiadO8OaZ0GAassLsgAUvqfbyYEICUA7
afWHXa+EGuVMJKZ6B2g5oQXgHuAuQ7h/MJnhbf6G+pR4qAaTbFddkAeufqKDyZGHMavdx/KtOgbk
LZ6tbBsQgT0d50NwHkjBavNk5dGwOKCNTWkGbtxFGs2VoUBd0NdLVmzhu9FGVCChzo/t7r8j63tr
JEr4pfSIHDtX5fPV2ilApT24EaJl6MHrdReZ+qH8G0f9PSCfNCfKkgDTjBlifcFcN66G1VZSzLVs
0S0+m3o6VH063NrtddCTvSCtnvPdktCUQvNzWp6fi4ayVR9ig1RgBrBBmDbkH1amMO9JLSOrBy0A
otvrO1ovoMZxkp09LoK0TCdrBtrmy9NKfj0xkHrklJOvtgrXBxVlc61Du/ABWu0Tmtbh2vPvqWyq
DrwoOsMyquRhVdbs1jNgebRxQ7BPJwoJ+YFdiajcHEdgXg5FKC4y4Au7CV1EqtKOkC/cKLSEngvJ
75hnLI+lQBica9bu+AsKsXl0WPM7ClBQ8Mw3/AaV1JmOQ4uSBP2Z8w9wHHvnEJOmL0Q7vioYGjNg
/v0jZteZnqT0NtpNqDXLcYx+cVCINTl9rwTnHeIv1UAVQA1QLIvynlu/aYs3J2NwA6Owaz6Wb7YA
D+FgJtiomBEsCLvfqyf/p3j55x8F3j46ITP6nKrtAhaQz9F/y1YhOulW7rd8XfMU3l5Ub/0GaMsX
MKmEcfUalDrD1qcEEUX9oH/C23ib/6ZcvgHFAk+cTFZHAnhkumr03cn344uQ+HCvWRPL6m+VLGH6
vS9pSxTmCj8dl5O5O/esZIDEVpCnRaB4vrF6Ob9k/nn413U3xXo/dMkjboWzkrLcu34gH+/Wqqj6
uTAab8fG5ARCRrZ/rfL8+61Mv9Sj8/BXH+3S5kqRAhGrZm09T6MXkZzqpe0Lbyp8r8XqyW0FtqTV
6WR5Z6u00/I1F7vqqNvs9CxF0cnYxCfD4kXPoAU3XsL03TPlkw/7ACES62LRgbyWVOxFOWFRtd68
KQTtl+b3YmWdKXaB1MuGYgDBBBK7FUFdWrS7nxHAAlKaYyei5KxqTRGDHl7nOmq0epVvkay1XPdi
qyCG1nwI5z/NexFf6rgtN+mCzV0JWkhIHZhD5Bu/8dEBsdhajtzrUDbwYetxwYvUDUcf69ajL/jZ
e0rcQRu1pCOKxXjPT/YCDEj+WUDKhL3HyPJNU5Oy7leDxDrW5EwaL90pdGB8WMN1l8GMAZMH1im/
BZJL6oZIiA4RDewFA1aGIQyV6Xuse2jhaj/7g89N3gwqEog462N9LZ171SEj+MbRggSng0juAa5F
trxVe7EQ9T1CwRLzovXlHUKZfgfOaQReZit6zcTOYVcQVD2O6v4akSva3zjvFt121l++q8IY0LCA
L3PEdHrbBmdvverxg0cwf477jkiVKuzQ3idvc9yv9f8MVQq28Rn5+coOXaeO4aIt8rO5doTmcIPw
T2l1Vr3D16Jaja+/YQPt0Lv7+JckvlVngjP84FpOlxH7QGthCIp8VrqxU4OGPEHbxh9465YqC1YU
xRj9W9fM9BC/H6r4EMmC/ES7xDjq5BeZ8voKcwbPZgSJp+wUwPG2NONG7zk6y1ngKTFCp3hWUvxB
P8+L/LH25Q0Pwt9VAwZfk4mN8yBAj23atFXsWT1uarsLk5yS9DCQ/AA6k2CVrWWhAfSJJJUOOU54
QID1xdz6IP3P/RH/t9RMd4bpfaZMhVUmvQkLH1pJOErT6WAe4mpPEQze9m9AD6Tuf9/51xij8IQc
+XmUh0EpknqWENySaZqvfHE/S2T4Jwag2MwVj0LK8VTvu764nssdDZLJtjAJQa/Sr6Eao2hmFDqT
3VUJCkL4HCCPbumVKxN0+DSQdbj2lJc2xFiRLIle3aHqm8J6bCPO5KauW6YTOk8JLCZoNjhnrEHU
4t30IF3/Uj/cg1m6IVAxsbLdLUrJ8WtgYUAVhursP/FQgKPMqNNFttd8P/FfyjbEJHQQmltzCk4g
lTvKZLvufw6piplB6td8nSZYMmz9xUw9NvExnbz5MFSjFCfjcM0cgMJ+KGCrJ2w9NTwxzmgMHTSK
lE1ZG1/LfCx2xr61EqWe30HbNv5Srlo5kWqr4yuKLft8s8HWlMGv7zaVV4p2uRPE1ygLVoTrtOCb
mgKPrCBgZ5pdZ4Fw8/1fNtP3Kja3XnmGWWLJlRqqJaaw7Bt6AhLpUIgJCf0cdwPAk5sc3CDRVyns
LRGrTn35bSE1D8uii7KqKkAbOUcC/UBjqVYkkQBeaw9ulbtx4Erkxca9aV/pxY/5TEW6WYDCrQpB
zoKDwG5LoitQxaVhvmzhifWp4a8X/yaBW0Npq5qJBInhjbR+Ej1PCJeJooY3fNHGO7PBthPtny+9
v2O+FaVK4PmiZjkbc9t3FvJ1S0UJA5rnA01ZoRRGnF0XqqT9ZEU/yv4OZ3mkfid4G00r2Z3CDyDx
17A8q3MD9pGrikVMxCKmqwjGE6eblB9iqQTBY5U34xM6vs4pckO9NPdFa7yfCVOHLAPUJP6f6DrZ
TclXZ2OM0amJ1CxrZwvhFCukF3KAoI1rQjsUq6sm4FNyxxdtWzlEv/ctNDgMVmePA4RUSMc7n8cg
Gm/wypq6c2ch/D7RoMC/WQtery3U+E9N25En4RLk88+jXL7v1LpY4DtXD4ETDKd503FGjO1S1YO8
Yaba6KEg8EVwgFHHMj9mG7keCujWssj8uftTYgdbd/XsOf/7v8sfiIXO1XkougjENar4UjsgRuEo
eJTQ2ZvfxIWyrYCmgH2ickciqWC0e3l160kk4YqhTkD5xPb3ydb1AbygKn5H19caANeVlXRITFpO
3kxX5WnPI6NM7k9MqVHxWSOG4fs71D+Y44Er9F+9LnrTLTVGxIUAsdDjnr+5bdblGJIVqi5Jm9FO
AckB/LFrLNbjJppXEFf5xdPbssI7HGQ6lCaIRQU/q1QsWoeFBzh759eK+zSJMcfPpvogxM+JLHFl
Ba6KNO65FhaLmQYl1XwEttSR0mNdUdT5SJuT8LlojK98xnom4WLn1ZqNOYthNL23242KhGBUDSfO
C0ooQ1De2ADgo3acCqck7ictOvMzRHB8s5at0duZhB185fgy17QUz5bMdxGnJdOJ4jtZ21QBvyZV
zmQ9tt+LOV/Vq3DKiGNBnTeqDfMw9Fb2W3Zu4nJ2OYR1eAusDlYbNufj3Qut3KAl3/JNaSS4/uvL
pEii9dUGG62YLngR7zjkF6zqXcDCZrCDd7KUqLYCddRqZZeBqqCwN7HX3bxvjIBe/9K2zVqcWOR8
WpWqExG5PnROCxmLmkdoFn4/ZFLakuQffS7lhoEbr/0F2vgtggkz603suPeCdGXfkcTtZRrTWNm6
MISVvsC5g+r+PY7dq3mwQJ5QhwtBKEOlaSVtgdLd4Nkvicee5l0kjqwJXnnnMFe+tbXpOVaf2rGc
RsRIL+9XkioXQ8yLM2tG1m1R91lfrd2j067ukReNUigklLem4lP/YEPSNatyxTvrU9vwNOvJ9lxs
yx44ww4tADVaouCICrINBNS4t5bSlVikbAIXD27T2XWNgSCOxSatW0kuQC/SRZoElqdCJoo5S4Mh
t2ILqxfwQFqqbDcFlrBPoMluIBwYOvO7yWJqGykaSyPesM/EXm05VTC8UNL+5kYh6MQNa/lgZTMS
+8vrDRQg+ebxoU5pWbwxwF9o+wuo2LZy2xeuqc2ge45j8jREPqKILK67KcNJBnOfLTLgE8yktYIT
mCiGSPBk7YIdaz8Snlvlt8oDy5D4+UfXeERCZhuT9HtJ1ULiA8ZPt0YnCe20FIQbvS0qk5CY5uQB
hp6G0fbc2raxGX9QEvU056kgvPA5i68s9ME17bUt6DNCyMRNCDqVTApJWP12BCiKNrPVQiP1VvPS
WPssKQf19XORIp8jsJFbCNSRnFxxPQg3tsphNbTPewBdO42uup39ae6dFtxUt0NF4dhppNLO+c/w
bXmh/0ik59x+gZQ1zJSV790ri3+TCNADKX3qoNQAS80yc9o9qpGj55Avnj6/SUXa5Uml0OrqJXrO
VjWoCBKFTybVmX2Ho3rWCYfPAOBPsIIyLqvYERtet/rY8CGHXhr6sT4KnDhmm0PDAv3ypNIOgtCH
bFQHclD/8at3eEOVmego432BiUtubT6CsKgeuenPRkKQejaS3xxBysreRN8TNtO7YxAsdhquGUIS
d5k04axpvQ0T9hn2OLaj0v8tqzSzASZTgcHQrdgiSEfPK318mcRcGsJ1WC+WvXLo/n54jT8AXimp
44t5nFE59/Z3Pyg4G8BMlAZZOKzu4UZ527as72LJahPM6aAzgbA4L1IM/ijGjhbiNMMnmQc66HUe
JmcASYs7whHb4frS8QCH1+qQsX8b8RqsKDa2kD1QfOiPf3UqS2P5m1t1VWjDsIbeIrvhF3AUTJrC
K5Ep0Ad0Hdv3exM+L2glLEBL6I+TKqeckEHt4uf1kcDvzpV6VKhiB8nzUtlxBIepNdDo7x6t4z66
qmV9ifM3MvKK46ZUoDaCPnLv4LSnBwsRZwl+QpGuKksLSJqS5Nq8JzcMbfQCBQa2/B3HzHtTBCfR
1EB5XQ6a0/uNuXhRyYGn1so6VSnLYXcu2oIN+lAgQG+/mLVYM6E/wuBIErNNw9QPAU3Mv3tQoptY
VL8LCDzt2/3SzvHrF2ZkftzX0N3BCDlkQ2pIr1/c30eAZGy671Nq0whgtEC5QAcXoJC1Claz+mJb
XWcmQEkUmxz9y19lJDk+/jUTuK/YWKjME+OEifEZEn8Zx50gUAahqKF997Bv0K4SlGGlhZu679dr
MOxjMKce6RNsWSy7VKqY0CGSnVu4JYqSgttAyv7td38HqfN/HKw7r3ng3QzjmyiXdOwUhyQWDLZz
DY1GEE61GdLPs7lzP7ipxJHw2SLjjdr/PAWW4UY/UU3NmtKI0YS3DNIN6yDxlfZmIZ9TBRIQy/hW
91/UEwWORFw25lnOpdJDBMrjcTYLONVN/QzCRs2x4Dy9xnsF+xMfucgQahRJIvtsPJ+yWuWVq0ze
HbkHS9SrPH0LanjKSYYnpt16HaB0nJAG+8D1ydFWsbf420BlfkiJS3shwksl5+68ah19ARawn0BF
ybgBiF8007buR3IUOjQggtfUjjsbUj1xWSQaNt+z2PnIRO2x+PN2dEutki/k0jNpJlkSHJ7U57Eq
NORdhXh6bmzHIorPecp2jZ98To1wogJ25vY1k5tiZinTcnXRgfGG6QOGNwifbwUO/iELjLVBS5nN
V/D4U/hj6vlxS1Vi1QHF/6Ige5svAYiyH/fnM1mLYTA6uOmQQFKfENmH04BZ7r5bt1CK0PmLPeHT
tPNKEmpbw1Q6dFS9UQp6A1zZeO1bwhq4IyHUElPPdsYX0i6VCYkeswyfGUuvv1nQeAsdozuUzmkz
mQlBRA45bVOVIPZ95IJRoJKD/GaOoyYwb6yj58rptwjGAjTVU+mEFMNylEtESVjdIgXicXBybjbh
TQNcdi00pPV94YpbrWgFsFuhN5fYFtTeyFnykD/Mi03oQ0Iwq6wTwCwE7f1iRHM4rJGOSAeob5Dt
q+Bus7muWFy+L8siqxZraop5M5QGixLqMAXFTQooBxoYRIvmLU0q/QcfqO5YfaJC7Tan4e3KALov
MXAXs0icVd6h/5EyiJ68idode5PVxfN2A8zz3kjGur2mARtrwQlBXQmLgjA43W/LP1iGtW1oy9iL
jLQF18Dbzix+e/xHlGsym02kMNdcl5gSiYa+WTcRLVZ8cp/8lzXKwBQlaLcGvbRblZQJZwz4GxnK
r5zVVlFj4HFKs0dMVlTUmew4Xwz8oLLX3NpVejv+AHcBhrNAt0k2DaDVgQ77jpxG/Y8E9c7LBj0u
+XaAfL56wtlpiUj1x9z3Jdc/9kez7HrnNeQ6SzJCisE3iJMFYK4XFmmr1kIgG0mYT7IuJLJ9Lhqr
4thokFvWLpRMAcXYRJWWGOVrRf3Iz438xvhdKgRoiT8V5Fin1r8ZUJFcTK1Iu+6fpIE97HSrAPTZ
r6xG+xkdmfZF2r2Pq3hZemEV+Gw5tA3zlN0BbfTEEN/ZhH3HMZ24VFnx8bHtlZDOtRft90A7eGCP
Ch4OjHtLLm4Jo60OHH045Rqdmrofigq09cXoBxQSY5qUhSw+lj/IVnY9VW3jn1O3uhKaXAP3Xix8
pyiFDZr7TkD8KNIqIxR8YqedBhqvzZmijxzCglUxE4xTO8fOBaGMHLrvrvy8Ryr75oc8+sRMHY6I
QXD3Bvt5BjDCfSstjJIykKUpQHpD3RXTKUu23i+BUjXEYoXFGp9IB1E5dlL+5tDBQ0s1renL0piq
tl4tku+Tn0E5tN004B5/9BJ3y8MsSXpR9kOOOKdo8vqKO66bXJNjMBZyKeVDsTM0C1t3u7KtTUXR
w5ux6cVMn5hRwDcp4OrL+ed5xWhZjXwMdGmXwBwLmiTh/LrLFPUTA2vnWJOFm/rB6GZP7OmuLIx9
aSdaRwTKKJXuPKfQDpX+3cYa7GaePg4M5y2LMbLg0srRJDOmxxFZGqPr/ZVpUEhC31n5rAVujUbY
FLErQ3nb6yLwY5sOyj7AJtktUwgpS4yMp4u+8JJRkXjkYml4UVyvhD2EpAba4LeqrSd+1ZxAUu/a
7ISL25HVrNABNk6DyK6GqAJj7jd+oKPC3Xb5l28gJjf/gK+cCuBRHr64/fq/fsNKJe16TWPjK/I9
gg0PhGuucL7zqUXw68NzBQjgroboZc8ORglv8fHLK+ddVURyCoXe3M4yj+ozKCpf3m0uWs2F9cLr
py2hFyK70L6F4YVhJwo4Sgr9w6yA5bWhk6A/mGQfwgqiOMCoIjy2muXendI6/BF8pSAarNrLAaA+
FJMUreVyFm/X7clHrT7Wlf+myMg2F7czeD38YYelvZZ1STh3EOKoLdUYkc7wWKERhfJD895YQZxa
nxbC0l2Y0OSKrb86R7KZu4jMIMkGrUpfcc2DQ9/M4oLxKYjz+1v+jTUVyFPE3+ThZNwT+bnlP5Wh
P84mqe7YlAeVU4q4IGWGjIxJDYBdo8AklGX6H6cmAYK4ri8Ku3yBXSRYSepLZmH/ap2+LisKjZT1
t1Sv7e5P0kK8KtSCQnBbLH/p0nq42mDj1BF4R9DB+MM64hi3WkOYYaps4SaBBPonI+FRzxhAzeqK
Nd3sWEg5OO4LkE/WVMWsg3HO8Vjh16Q+2oLXNkZIaiRsE2HJTR7xzYOv0oMaDsYX4AT/xGcFZxyG
0Le+7K5jMwQo3Fz7uu4lA+k4CB5Dxu1aB+miQeFOXHR80srXLRCCr2Y4PRhd14LiM2qO098SPIH/
l9zyORCjooqWCjldkH4QzXaLsHnvMtWzRZaGrfXdUlPCjNTFy3kzQQg0tipB+Zi2peXRXx3uyaw/
0owhKO5O4QbhOOlQQw45tMZooEYQyIYymexhidDsRQK8KZPUNGneZbehHhDxbUksshZUoo8zNV7H
YBlcihodeE6Lv3qZl39H8/hBMvcueOhCOjsT0IuIaVP+C9mVU3aWWlmTrEggcYvUolg9GyEPyoQR
b1NsA5E6nUhdtrJ/dBlCTQL6oVb8LCSRB512/owW1qGHcdwIoPQ9rWhMaA/Z1Sf5NF3l+z0rUcSN
AfFZI/JJbYfQ+Sa1I7oy4mmVZHAaANm0mZuQgih5hYYAIpVS1Duq5xs0AX4etnCm7f3llUFtht/l
Jh7pqBay5r2pUvzn832a5GKtbmCs8DvX/r8oRWJvf2Q1t2hrMx76vynNlXhpnBc2E71i4n78v5rz
IgUpY4OcBVxgXxyTMJ33wYpC4i7lCP+tksCJc56bjgAv/H1xpYJZpH5aC/S3nFOfWQH/b4DckxxY
vbHyHdtjQla3I2dBTfn9aItcKStaNSFTeVqS4Q3xiftm7DrrL+LvFuhLMKM9WSEIh1RK5lvGZy2c
TzlanvJhOxI/KTGzjiZHFehmdhOAVXNZPMjx619FZk8hlvgqE8muO1RlC76OHL5SEpIrt8KgG6Up
gVe3/kRQ+thNrrjEdirPK5rYpoQ5gIiSFAR4JUxOag5ZlA8LJjABYhZWvinIjKXbKxsjUCWRDykF
/hqGr+4a697DVj+ns8bu+yAb5FR3Q7YJpwfudXAV7eC57U+7mX0KB924ivlDX/W09urpBpWKlj/b
JL8+1n25ZVb28y6yKOvIEif1z5AnWIx6M+WtsTfvOK3ledwoT8u4/Y0oteQf2+FwbcfnJNgvW1De
RDiZDGYdjvpDS6ZjPuliaoQ4NOHf1aWtI3dylI+wNeWDWxQXMdujrSAp/kkjT6g5WC45LTCyM5SU
1nIl7iZaHsP1vLTUX4rQaojcRnt1czqN6eAqBPfLM9+pIAe8KeCP8igGj59uivP7Iz5eTPWmi68B
ZYKesCb3moCTtzCXjhf1SOjNcAi4ly3NSei4QET02AiZGPsKGGytg0b+MDa584WE7/RcVJVIJydz
93Qs30a/vinXnJgOwdJzIzpImfPZ/2gHCYqJrsBjk3ZTrp6Sw/QGGyELuQ6mExT8+cssd/DbJcQ5
9EIfdX1FhwsMOEH6a6YCikWHRvNUeirXMnx3vdGvZHRtwdOJ6IvMEb4wsJQ6oB+oO0RDBGeWCTGQ
FitiKT6TM07IF5zrnazIl3R90onLlCaVS7fS6O+36Ae6i0Utn/3EtXgi9DIWkvTUhBtulF2li48L
SBeM7xb9lkhBVs/6WXb3+5WjzdQ9zFx9OW0/xDYx94OVtwt2BUuRxYoHnokgtrY7JUk6nzOXwR6U
7WznB2hJvhhzrZaNRLE5ayGyKeK++r6nmw1rJH7+mmt5A7VMH4V8k/9kCy3ExQiDJmqO/YZxZhY/
MlxwEoqZop7fwpPxs0FRS7YRploMM3V29pp2kF9vHhpvxsIWFB6kfeila3C/38OLPs6zbvgqoU1r
hzuk/t/kk5zIqT2jaA1CK6Cb/jTNp7gYDg8+5oMU6Gx02iXevbw2o4t0+sbhgBO27EcVgf3OxXN+
+TUuB43hbu5U1L2S3Bzm39X097Az9kZJbQGhAXx8jsjVKOvFSqWN8XfHbMsxuxZpWy0EGlHxWDe9
D6v+jWfw7W99H10HwNgq5Z8d3fU6ycqaN/mwhjHTvM1a1NrwxKFvGTR6YltabEFJvxK2QnsMrpye
/g8KHH7syoWr59hErlkW7wmHPkHOnsDK3gsCEKo15H30H7hZT5/dkserZhweVFU9YaylqMGTaAOm
+PK6q6tvyPstJLq4gtE/Z6Xm+8hknZqVWdE3Pqjp/4NtUmn0wWoLFU8LLtkOpmCBpfHoaBCxzEv6
5hkIjhvC9FDv+CfquaCX4AVAIuYfrKVjHVJV+AW/rv6UukLBx1eDULhooChPeWT2pJlhuXVVnWkI
HxBfZElmLIzsZTCgYfKVcRIHxdFEwaox3MBKRkDtlgW7Foy5mrBt81I2j2LFBcUKZmJyOJaP0BMw
cE9dyx7Nws+KPz/Cs9GqZVcy/vy+bjTOodAlDMVa95//jV3ra0rSJmeqsL7HkfAW0Mq90Du13p94
/4pU9ck6ABvTqJeJEBuhvWfMjN7l6mdKgFsb6hutnkfGkcmhpTWhwlRRn4KdnOJ4FVuH8wyFHUKC
p3DtqTsJA2pkb0RboJSubXk1MVczId6u+7ry8btKMnyC+TpAAOWk+vr3oaAxsR27YEEy/tASIw9c
QU3K4wejjoiIDxHNS7wQCS7A5KotBSkYT3Di1+2DCgvB2p4GDrtALUSkWu2UnR4MwwNEmJ7AsTaD
f+G/knGJLNM3GE1LsbE5jITAhNVe/jq4XT0ccSB/cjy/TiMLzAKaR2lNuPu/7BDsAAvczKN+7AAN
PXS4Wt/lbnWIWWcwDWWzaWzxF7FG/XcAF1EEJSA5HC3X0a4txbTqK8AY8xruNzi5jYtgXY3JMQQt
NEv5Y0Wdch0mcgDdsdR4XhDLbgQHSbTkwOdvAJ67krqVcfIwyEz9R9XuwyySEqg8As61JTqo5QST
cm4VzJlwre19pP07Qzdfcf6y5dEsmv8ZHD4IgqTem7pwp0+jRxVxDp4fRlQpaD5c4q2bT41YuhPh
Yg/LKA2A/FbMYA2R7in5DviAJ3aGEtlJA5E+3A1SQ94oLelL3SdSBAuC1lpQX8XaPQ8GjBAriXcZ
dxSk51dNpq4MsSYE+XPHBu/LpdbmqHAV6wbIJywp2Xt5As0NM1+vnWDhTUiHS2HysTulIeQV09Cq
nmj6hrIq0Lg8Uj/K3Xs7X+hKmRqauaDl93T10UJhcpTVmDXirNdu4PExklzSZdWncRtHloejTkPP
f4Dx0GT4e72SEV0xJbpooQNxeK+H61/2jvxGEoe1s5Uujv0VDCAoWBvarv7vpv4X+QB1nKd639D3
Tiqx5xrRaXjIYlL0/NJx9x0LcpXuAn6r/GA5cEGy4AbCBv3eyAZsysEMt72E9Nz0sxUponBwVn1v
4CT/dvB+4WPNjD57cYkDckXLblizdpM+7WHwIsTUSoyfwyo9f28KiPdikZ5nZhu+JJbHBW9M0FQ4
M0okSkslNFFspM6GJ6rCe277NXZ3kSIdrIIO39KT238ZpkWqTJZVH7jBukbVKvYFCxiRccyTqSNP
QJzFRc8X+54RYFb7Pya9lbWpN3TU/SMM6/fcjlZE7b6zQH0shQIvOk8PuiQpE3i45SsyXDkk6M0E
VUPwLfTw0CgFmzd524wes+kxSaDPFbwPXDFxc8bbWcJYlYgzvBhbtzkH/1IuKcXccavwJzYixmO9
m+btwYAWNq2TL9qNzEyWxmQVXd/aoKeTcGjDA1aWg01a/Jx2HTtodXGMnaEBciobj/M13ZE8BPmh
lAjGmp5hW6Ie/5GEmExDd56Y6nICtkiE0kK7C3MKSPwsZq/G/3kgnpRscEtp4Q8n4l/VMO7TZiOq
HZsWmx4PIhjktA5ggiWD5cvQTb6kINtI7T3DLT90v+CKGc0RbeLu4gzoZZ4TOlmliVgVRytxSdux
mrNmQDjv4QyTRUD+dRD9wd0M7fP8xr9WodVtU24FlnReoLfefGAZz5ARo0OoBH+DbcT67SVY3OCw
Re51P8A400oVdS+jUxV7lrQEhnxlILj4B/X/JHfBBHNCt+3ZzDM/pbx5/HDlyGiUwhR+D0ntwZRx
ROZwOpqjb8uc+zCNJN+3B+6fxOHOQxCRzgPa2iVXRifBiRx2C/nPD2hG91fGnJ2lUOisQUcCFz9t
BmYGW4PHSnCILqp5DJ/hOn/PHYUQCq3PTaCGomzgPzS485tmUi/IzZe/cz6MEWtkpGkdw4t2K+9U
5uU72xb+MOzjgc4eepmIr/hWM7AQiW/CdT0oKgGzkoyGBEVJVXnGPI7IHQXYDW6OUbUkwtvzszJU
zWl9ybgNcCGww1lqvjzUzh5asZxgj0Xb+TOusVJry3lPeduF8p9VG2Hfj4Ehmg4jKGXjDMJhwg/p
zi4DAh9bMam+L0OQTEDQROenurxplZJz58Ykta3WLADjjScwFAw+lva8TYzuKLfPWW5Ci7DP18XR
7i2A8FUvmJp3xo/Eu9fBG6co5ToWOhuUKQF5634jVpKJh2YOOVw2cZLiEWQGf5+kzDo6JG2nVmsZ
7KaiKMy+D9rQH2YTmkDK3h6RcYR03Bz3ZeYo+2ArrSAwaLHn1JKss7S587Gxm9hOJELL0PTfogE+
5iA/bWIPxRb47zI0RBYliBqd2oBIMZNtHDUlFDWzn8q8WAv+Q5cpBHpRSdOoYe7FN4PckMU/+Mmr
VjP+gPg3K87/y2q3LDwQF13Oi7qxHY4UiOLd7sVyS5PcelWwDCpGP8IPS/6KqxG17CKRBKRlrou0
qxWFfoLLFPMBM6Cdvt8O7ry5it+p7xRuAzJ+Xn/Qbjvo7MhVAlC1p/qnaIAlHJQc011mxCtvUm/i
ZrSddmXeyejYm+Y2mTK5/KLPj3ysXIGWtEm/iO6SjCslNZAhfPpYl+aKC2b7DmyA9UWCpNWvKw9J
WZfzyVsjVimmTSGJ1yTEBTf5uYDKTc78J6Rvw/g+goqBG2Mr4Hl6SCDej5Y+FzBLcaB03PWpprZN
yZJ/Zk6e1Y3u+c7d+QChrBWK0jCyWHeMSFYGNGV+mgMyJFNZ3R/AOJ4iJBC/JeYdL96AJDRSXOhU
Ae7TdsZRNXQOn2QnEFVJSPZ8pw+MJNVY5EyZwmGZOZyVk+QygUTXO+7hNGdGsH76/XQKiPPbljcd
lZFOQ9ZqA8EZWAiXTzwlykTRLyak7fzF4wcjMiPo0+3Qfwyvi3OJT/kirSxRJ99yCledNeY5AIzl
wgHZ8tizpreAIPBmaJMpcXlY1x3Ak67eSr3K0s8ziED7LreAYkSpTh4Tr6m/sIeH932tUg8MAVik
nzDKbJCIM4OJJstaWkhoJH6JnXPWPDfM1imVcMbBm7QDOMjpgzwfOaiiyLYt085Q45hc8PbMGC7O
g6+IQtEtgCmMTCKTqk8h28oNa2VXg4HGFfK8FirPh4LrXB3blM5mE9JGpJ3yAdgy1H7wMO+gPTOd
ex6CuTHxY+cNUezyna0ynCE2R3rIIclsgEcR7YuVFzbsvAGH8hbmMsguIKRyD5Y+wQQd1sk75SCr
Pskr9z9ITIIuSGqr5sYN36Gr9rUEXeNcLs7Jrdj6DUknfplbbQxsikvyfVhBA918eEFE55p/Y7hV
KvUlr2sUvI/ItiQ0S2lV5RPnDZ+cpuv8weRtJXuHJc+D6pGSIastCAAYBWKdnMZULpFVG/wpb0x3
liU8qW84i/zTberUDuyvOa2ow1wE0jaUNFYCfbEBwKqA4reHKv2sVTAGCYszf06k2X9E6xwzTIEh
E3xIMcY+7oK/jKSzOx5NSRZtY5F+GjfQDGHDf+GIkebSDk9OfycBlGfX48hovdqcY4j5Q/JwmtCv
MB6MJaJuODo5TgaXk33vYgy4sX3qIiFmjKuKk8LSORGK95q77IaYKiFxTqz/bhicj/7c44McM+NY
Kofhqy8fhfsMJzRAyGBLC80DuTTo+QQEuYC1eTz9oC9jY6IFl1rL9uLKJvKPD6aSBgIgPE/rLfv0
NAzLpV1kor20ZJ7iJOd/hqB3vMQe6ixsO257pIEtB3KdsEPAPRYL/3choZvXUnyG4oWBEO4I+tKp
qovwwXUMRRY8jn9O28xFG4PIgQvSyxYnZBrzVbgAYwA0FwyPuz9LaT9zLBYCIcPg1Wp0OpO1+kzn
cXyOTqMI6VDPCwuXbACIsPAj+iMpRgm+TQqrLFZxHAMYuGMfJx5sM7M0lsljq846/5y4mcA6lSyo
NSD+1avez2yvUmiu2oZcNuawdUF04jtQSR0qVsoG8XQJ9x2LNx6im9bzLXVwPU0Hs1fVDOMgg7Ju
1dsuAOhIRzsR6CSuakBthvmNthJ06+jGR5xo2JUtriMc8owzPdpoJXb5WkKjU69yCjJIMM5vaXXN
zZgwxyJggWvK8kCGpz4lnrH47LfjggNdxvrYyGdu/z5z8dsPPDexmVUDeWCP/QDveEoCjcrne5D6
1F0NZynz7Ci6XNdBVfsJJ24ixCRyg7bauoc8XbByQuSkShtIVDjAMObXrFPVVRXE5YfMMb+I/r1u
v7LkNwsWCr2dz7y8GpkQoh2clIolA4XmZ/J+hNP7oWJhiKULoZ8ceKJfWOyE/iBr5ifjhDYcQ3hN
QLnmXJ9MoTcGZ6TND3UTIa/i+TQd7bhiDA8k1cDQ4K1qyVvn3B/jfIxaeK5SkMCXQMlEageMhx/H
lM7GgSzTY8kY953qSHZQsPqneH0oPvfBPblaajxmBC/+WsdDh1gCEL0WZrGdQIwi2z9wb0fpjbCy
2dsFuwta4l15NeW5ci3VajfFQ+Am4YJtPJWeIWl5CdQdAQqzsx6Ouf0s7szd+h7ALhSveABJH9VL
PKpiAhkeRf9Y6mvFO780ANcIvTiRTYLouSZqr8OVfapfYJAGoUIKNusMz8fBtKUJoJNPPTl/07y3
9yQ2WlDNFpk0u5Cqc91ucUXjdeLhI/9yoT8LkIDwNUtHH70Xq4Fz43D54a/LAHcx6u/pOakhDD/8
OVnv2Kk3I9Ifwf08Z2QaOqiR8/dAbCrttyFnKEjTV7AnfQYVi+rctmLDTlHQsXwvGObvFUXGHSxM
kmP3jN1co9vPC6HfA7Put5+Yf8QFPS03O9GCJ50TGCTE8Ic6sqZfqjhHiNNj5yjH1Dp2Z5RoKtEi
LOP0HWqpqhKnRr3HG8jpyiixelytDSkUfx6K3rg2J9EjRTdBp/Jsu1J9pdEcgtIUT+F2htWpmlIQ
6XYELXa8ApfI0ELMV6VPsKFYOS0qiea0K5mKyyFfWkugJsL2aCIxu5dOwOoVuBIOpenPspXtjYAh
j82WpMe6e0fgLievE+m+R5UKFEB9vgNUGsRE+CdkovZWePAu7q8KBqDO8TOjyRvlfHIPR+l0ZgVH
VIqPfzTEnhWcPs7Lj6XFtgvuUkCUiVu1X5Kg1bskPDWnPQSDioge1oTMNNz2jq5pRnxAo3QofQaI
C3URks68fvhO/mRN+J06Flz4wdm0J0g7wH8fads5a4PIjlLKdd2+DGn2Xa8EGQqeXSfNXLlKgJlM
eXpYIYmRdEKX8SA4pYaE7XDtxX6YgbnMvjEQMZA1hNJ4nw3v7fK3dXn/aLmy/fAK3HIWqHLvBpnB
SBLLvXrAv+kvCAQjdYEQsscEk12E/qlD1mKkvTfSZs5F0dTt70E30IUILUju6BiAc7hMMisK2B3s
54QT042QhYubM3qvBlpOJAosxBm94SlMt71pBQueKzPCGRVdBt6ZaBI2LRfkeNR3LswTpKWUw6Ul
/5coKrwVamfYlljwovPMqyXEvNZsAEzjBlT2AlblaRC6CAGKQ6vStryQ/XlP7Hpc+FBwHgHHmcdR
ftvlB5GtsuVBjxIAaqL5z9iabLgDCLptdkNx4+MWVlbofflK66qnNX40S0ww+Ga6hjDuPzC6yelI
S5KvwtoVrIJM8a4WCn0yoedtTQJ4TiTQQx2mOyVOHtvOgIZjpi5aJz/AVo+WUAn5ZP1gs68ndG7o
QZ2DBap6z6aYw50gtnS/aCuuB8DAsSPXudUlpzRCh63ddjVOaI4ZtAmJYVnYCEbcSV6LvuGQ/60z
VwASPlCSA6EYBR2ZxoNB+aQl6310QS0dJmgm8dUk2mzHQ3Bkqk5dCxk636stMt1ouQNueXJLa/dn
sNyjVUqxS3TWWQ6d9caQC6RcIKPgbSPvk9pePSYNbm5QydKpKYeO4//2yD9HBaSzqVikRj21a63c
AoVkMQ9A8TrhOtoucUVLpkJdyWN85IagPp5v+us2q6Va7WobGkaQnm9PalOXvcNvmiC+r9p2ct3p
7EZHSk9K1NQR0AagsibZ4We+pOwmdnz1dAi4Vc62sgrLiCcaW/YqLvprCV0MnkYh2rixQ4fGYLB6
n9wAGOtbPUxlR8BccpNa/1JW4Aaer8fqlmI3fWTZztpWqWbQ2vqbRX98sav4bV1CzpFGCvs2gbML
SnUC5Fiee86Ikd4bN9uDzjWG+kBml6HA65MpMGaRxBEb/HRSgX1fMGkFVObqjHetl3k6Rri9VJxH
dNx3nlFQE+c5KFg2qbkwpUtUpRlDeCkFS0cXCHcnMhIdCeKWfh9sUID07D/RHHXlDa36pFrFfFPP
8fFqxRHDyQiRYGoXFdQV+hWwd0/mHPx9BKZiyJOEmBQgDWrua3WdC9wlLVyyCYl5sTTS0E/Byaf2
ePbo2dq6KBwOZZx8ibMcqlWiyyRkSbFtUbpuLhQgkTlsBtATGy4vYuI0UDw2a7FNq/lmq1WtmKNR
FuUKGW9f1qbDoU6KJSQ6n5BDIWRLtFcLwDOreg5V4lcsVi1eXlKPeBDlYmTZub2LgaJ7mdgPPa+i
Acx3pTkoDY3MAUfBp0QhXhOSjiE3jSjq3F9UbYGlgXPtGjSwwoh2RCeotrYAVYGRgxckHKOU4Wmx
yl6wOtoAtHn6PHd+Q573AlDOqH17Kov8TTakCFOXQe8gOB9AAWpMjTyLQ6TdIvoknFMxOabr+kNz
PAvdpteS+6AFGDtm+xP1F80U80j3blM3A8Z0FWjlo+HJO26v5zuHYu3xER5T5wlvjcyL5x1gGiuW
J/ScqL0tdPx479PdBXDW92VDWija4VhxSpre1/eR7aE7FJ67sd9jegajIiuHLLJ7vr4oRw+P9cxv
kv3V0BU2ROXavovSnQybAbcI4OWHp6xX7DI1j9NcvRUxNVTFDjn5O56T+qfkT/CdnrRp+Hpi54ti
arTN5X0WCc6y3OlgYZ43K8cVtOouiu+Jls/EmpE/l9qzuy2jOCGOrMGlwhOH+KTrDRzIvkCS2qAc
LtDIzkgrudWZ/1N7ZwlhDOk/azoRpXdudO3ar4jr18cJRU30B+HkU16+E5UazdvMIY+R67+v5JVp
dnmt53IUhnFp46s4nAMc7tDB4nfHZdsRbHf4URLnez5x5qPTHrw/Y7Vfobfe8lPOqKTcLNZdtKWE
Z0QWt0SVkBl5SOHFkJY3R1lbN4xKLj5Os7nv3FzpXsb06N+2xGovfj2rEc3QCGqdhklwfYzsvrkt
XPE0ahqLM2D6vwjaEB+ln8k0zI1RjIwppBJJzEGpskT61Kqp48M4fmG2Nch8+WhrTOFLKeRSNA2J
sEtkHCp7DpibrYzUvpXXD/4bR69/4jvXhKvrZ21f/LQhUvUFbMKdkI7EWEvn7+V+Gh/yiSlH/I0w
lhCs/s4/LikE5K5V08Tib26I5UZ4jXgAS/JpFVoxmS1zOL2j64a4XH4QMdTOdUqGuPlbRPRNHjjS
EUxFzgXqimNZ5pCX97cTK5KInyw1F6Q5Wfr/LsmPhiNZWCONyCFIFqJj0uw0OJ3+7tI9lo07NubI
9iMLMCI1fAxM0po9N2UqGm1r65/JxPtLpL+qeT3ew7V/wxqSkQGuNj2Il2p9uCYiofao08SkExMY
mmWRm5LKc915utA+4K/Ea+9WjdlXqa89/5VkmSqArvDyYYUF/D5DFjkqQbAaN+jacoNnd83cpiJr
1JTIeWQm5O8eDhJzixUFxITfKR3gChkZdAgyU/VPAf+nyG4QcFpiucSNlBsN3bft94cOfNRYNdlL
3Uo0TGIrVo/RKo74CdxkcF8uEZOXWFsSCWMLagVa97UhkFSwqMxsqMWwjPszCD/jYLtq42AlivUj
TZ/KbOyEpK+NWeImJ5h3kKCuEAUXpMmEN4kd4uXnab7NHEn2MYvJMKBnt3xMrBMxEiaeprHfG8Ye
A8Z/E0TirzDZ4NTzPOhHTHgZk0hzgB4v9FkNKNoXgroQbrlTwMUzvsrPMRHys10x9vwhag9Fr60d
1LrMgTjuMYkdjSVW5O+U32hzHv6orYKWMnXcp/D96warHT+eLjCfSvBPdlKarThQstJ6T7uPq2Un
J32flbHqbF/v7f52NkFv12CI+BESIJ0PH4aU35anJgwaD2H2gLpF+1CeoD8rfQnKCHt1i2o6P6R0
pW+ZwjQXhZia3LgXxGPsooNTdbg1DlqrjCARxCB7EUMB4c6Z1+5jDE1b4wGsfynavLQ1DmAxmr7x
RFiziDpgQ0/3Dtft1oIIPzL4y780Kij45XyECiq4//uLJSaW22F3Iv/8npro4y7XxHwiwptlROfx
bzpLqY6dadcUW5W6Ge7SZMxvheFtI/SPXWJ8loYqytMfqnrr1Le+vMu53zvCwBuW5fcw/BqZDVaQ
q4Rjceiym5gIB0ysZHyiXvv2utjJbX8RmDxvM/YW3CciboarzjamhZbO6HYtEQOLi6gfquwRypev
RE9pYJaHO3e4Sz4Qrmv/EHvfk01tI1B47zmm1uYJPJAMlmUj1gdnfJ9RlTn/IPNJ1VOYlUuDaiow
AWOeh1a7r2DirGS6SyQUiRKxdydq/g36YuYcbid/q6XSoWZzQ+328oEVlPnaovhGPhypel+000bk
/uFGIQ6Qi7w3eF1YznABWOmstE2+ePRW+UxN0FjLgiMlWylr4rnXjYEFHKuw7Y9WDzQoFHdyXW+O
YyOSO70EeeotkXYxwVRckxpfX10ATkllqxYIqWw1s2lwdsMO6A8ctdwrxEUWhvItmdHK/M1gk8bI
MoSkw96LgNZHHg3g0z9SFU13MexoTz5Z401E1J65/Hpp/fdVzq/kV/4hK+wp2wqJvsGsowerUNIQ
BOQNIUiWEnw58GavNTOOGbUvRd+b5XvA9DubcR4smvuWGl1nKZc7yCZcBto31p2ctOxfAOt1EKDS
tQ3OWeurJLDlf6D202zual7JXbkFZpCJ7sS+xugsaDowkjgwMtKxOc4DPxUM3BiGuFiLblocSN5m
B74d6pYjPV4GzLYBJ1Yzb3GwinQjCgsrqbMRwxSsG0hfQJ6mlhcBh9aTyUoU8VoKtyGeXK08aQLP
LUs3nRGV+zqq43JbOpz+IU8lOS0PQwABXjE8bKDD1LA84571jsH5yvjNnmGwdsBRG5DlFN0cD8AY
Am3/ukcV2A4zVsGtgOvFk5OiYYmCpfTAswO1nIV70MIDoEi6rPuy6nHKeTTDA1pro+cJL+fGYeTy
YJsk8kHnAeL5quEVy4G9+Rqonle3gWAwSOdfOD9M5gyE9uSwsveESFUz4NClyDV0Fbg7u0vaa4A8
CSCp9QKclI2ks5InIaTAQeylIk5uZpUQUec7AJIF49d+V3kti0cFo1wBfGc2e3xY6ZYAcZPVpdqa
JWjl8K0xUbnS0YZ58Yzyy34aL8XbY+hojRsyD9fFwg8XPOkapnaRgtQ4JwXSeWGSeqU+/6/B0KkK
Kq46TTKUs4SikLR8XZxJFzIZkapzQiaDAstlDrr01wevDx6nppzC/GexQs47KodWoYuvHMSZHv0s
Q8AHsOJ23yr6LIdFUuTmf3m0XtNgnm9PMonnuUCVsVcdNQMeiUaJoHx2cKw0dorbZtqbWCUcLjo2
zHhpZH8bnSyRIaASxrEbaZIVf9ViTD60Q4kkBMzVx4B/zPzVYGfXnG5PlGZrKpn7FZU1unMHkQjo
vNKvVbzXsZ4luMPuxAOp0ZXdh1fPjX21485R+lMio8J0hUoApRGw3fwxADfRjb+nB0ufODUkCaxi
oxQM6ogfRMiSedcccXBv5vJiX/J25ZbDsSlkpR7B/u2Bi19dMbZXI46VshQD4M2NrJ04uB7MQjPc
qNKradx8yOsOe36RQjhWV6KQhcoYpcYzFz2cFMLXcmO6dQ6+2ANejC+dQNIzzi86GGxAaxZKzZSr
e878HtGmkIaVNhFAIY2nxCDTnuSawFelHY8T8QDTHD7nKPdoNYW+wpzl1YbJEonCB3IaxZ28i5WO
qu865nKzKPCAgPF+EG0g84bfGsYKOtUpXMrTz/uKRoDiYjLexZemAZHZECHDA050IdmsEvWfaoZ0
guv3qaVW5BuHFjV1knwilEtf74LaTO2fDFS5Ox4j7CgkxC1z6QStKgNhzSPyaNgz6ESj9Jg4NpK1
A8H0fTn5xU8m45jcZ1KDgQH5VmcBchCYDMvDcW0AVa1Bgkgs5/wgrmNDPn6QdEk4hepq9aNnQJ4g
a/sOsC4Hqb5YlxXvqt6zLczvKvJZbaV0cOi4HdG1J6UtIs9dxnK39BuVu4MRogDwlzGpmnrdCXvW
ZHVDxEZDlHHg9XRNtFYzgTOBKti3JkNulwYM9kCx6GcvI8ejuwYXX/aEjJlDCWszbdtpNfaGEHu2
28I7euxqexrYKz3fJZm/6BviyXddhCNrMmLnhgRagfS2dqxWDAWn+PEKOXw21F99ZySiayXZB78U
ZKskHZWpGcGy19xgUYrWpHTgCDZV4m9w/oeCkkfJZjFkYg/KZ3X5EMTRq4uYfXrmzTRPVoTYPRbi
3rywwzM92AWc3/JvAOGZYYAeTybe6CxCGdAijwE19KZJrmIcS+jMqLi5lc1bejvSyiKA0BRK9PCL
uYn1CYXReouPJlBL7Q5qwl8QEaaAD96zwhzyQG1Ry0kPjZSPKLX3NYIwsVzGORJyfUYIl8HG2xIT
Rz7VZs/u5uSg9eXQB9bBoyGtzYE5I6jmNRSqNrTre28unp42aPVL5IJ2fA3DIfxN1litX2CIxNvK
qdB8RVBpxGo+ujT8mc1UZUqAH2k0reUXbaXnFiNZokH7edZAZnpu/5plZn1KQh0GNY/IXVAdOF83
xgyWtipHgiAgNAuVs9qDp+X5q1Dn7bpqNUD0M/KJmfXFLfvGCsVmPjK0tQhOTGaCohWCDrlLoaKm
EPsHyMVEv8qBlASSKAcVH23EIP+PKNUOqn5a3ZfkstlLCGBPDip8vLV1p9IYWRd2fPK5sdUZudiv
YUnX6sIMSisJuqY8oWxfjtTu9bIQ4R+Ri5EXqmsTnpUbczWQorCtY2crDfKjV4hGDSmGBcHFQ/vd
02x7t8D8jdo0QeW5BwY4Xt53EBxEWwDMXBkIGLc/3uRsSsgVZxmFE7ItsSRnx0tVUTSSZhhUexPn
/L/A2mHBhi1xRxersegQVIpOkJeERyYty0az8PmWzfWChIWyAt7g31V+dT8K9efzsRW2rV4rAEBX
eHN2NA8ZS0LYsHq6JAOXbnXqib05Cq0/R/fVgo6TAyaSCo7uhjWtV7H71RdOONUdZneawt6OY7Jb
9o/HfJGEV0NmKth869d7eApNqs3TYpM/VGe2/VllFTg9jW6GVQjAPmfgz/3po0LDOq9XEcB9NVo0
bEjr+KXzejPv6EC21mvo54UUDxXhEk7Pt23gN/EXM0X6ft2Z6Lkc/C7JvNml9V/fVY+Ms3qpgtFo
R2ViPHsdGaV43dcWb/a2R46859FOks1B4SLBaVdDG7Q4D2YFwbgLwSsYd0BahZBUOnH2MeIokfA3
psuRjTeY7xN6OnylEPKj0khoceuYHNRpaeleLtOXiFFb7GXVy4girQ8wnyDECzbnncVA49G4C98P
qW1ME0v83Mex/0jrxbhUOnkfUzmjtn9fL/Tn0616A+QRPoZJYRKvtZsbB9N6MGZKBzG6inuJR354
Q6o91pcPB28SLOY/IVwIabNM+XJIIuQEPpJISM9hrI4+yGePPZTp2Kqi12IJXqq5JPzUhUGxWHU2
Is0cmQ0vzVjmB5pg3dEmHn4XzffDq+66oJvC7HsThUf2Sb9bg5vA7D9/95z2InBI3kJ7SXVgTb+y
Lce0fvgI36F6IyrzPzLUqvsOKtcq6I98wswrfL9SPYZorfuM9HwT42Q0JYLArV9A6bObmjiT+06R
teA/fKki6KFVcGhw/UtQvHFQpprvc26TWOGdJyjJpTQqnSFbBj9V2+5wbB0D5Dg124GfJvTPy+gh
IMz5GTp11axQ14YMemFT+ubX5lQ8dDME/Vs36CTkpnywux99EWuVCvfKDBnaJN56/T3PllHnrz7m
rvEEyvYEEIzO6+fdBmgiS+QP/XbY1+LV7ljjbOKM39uFUa74VHvFoTxBWiuQsbSxN4TDmTRSLq5q
4IJAyDq04lJrfLFWMiazvMTrAEvkWbb8FPSWdNECRioVwaSe9Fpo9kjdiEGkZ2aSDLkg4iiJE9xf
WyiXSomAZnwbWG4WYVdtmLPOuSjW3dbEmgYjgUnUsJnhwTCGQjL5ER7DoNECR5bfEu794IIRWDQa
kZ8XzBLpKw1RrkWJJT4HSzLLi1zFyYmkcCqrnMpysCjL+UZ5eRMhingpX+n6kSMtTuNf0XX2qOU7
FXbf3dOcvHWe0fkK4QLJBlwDuoSGXMbLRbniu2uiU7O/19kQxjqihiJA3wD+kRLWRQGp4d2hW87Z
Be9GWl1gbiA41CqJQOZ2vpZrrejelreX29TZgaMd5y4NxkOOLBbtOnysAI97qPO+qTGUU8RSN9wJ
q3/de+b92ENb5sYmb+JXo0HJ2BVvF0ejuSjXappS72apqezz/y+B9wpdFuQhkzyAJLABgT7vkKps
6810tmC/qjz7JxYbiVYyL/8n6Mlf4/aBBzzDJuBlCGHqdBqfjnV1P+GHHmaBjyqvaz7EgvaZ/Bpi
rnw4Mj3CXFCFM5EBs0f6knxYZfwz4dG0JNCysQepHY25QeBFSDgg8wuAQ0vpIK28jVNsP9DAyfwz
BlaE4QctlMqtb62lBbSUJhHwcjxGxbNBjkYk0GV1bADnQrVJD4zCOjYvK+quLI4F+wEtVOTJ5w9c
1ayVyIfRmJnOCwSEDBb6V9prYe3T3a7fTWOUBdQxfhE5jV8Yh9WpMpIpAfn76g+J3TyC3WkYDhFc
wnIMt5CTt+ON1UAF9qtThDh5fbRFJ+GheDPxewHqe1TI1oy+0Ka9IOy2aYbDdtZd8E4kW9zyv4jO
f7vQImlA+6A/9/YTgTCwW+5DMJja5GJKupy2d7eqikz9LRYWZNKk/B6ycsEIYHpRPVTyQhlxGTj1
vLZjtlRsmV3w+RhRwD0p1lTozYn/UFU8IjvlDUg/DEdfV9lAjMGADhorpfDkcLvDfb3yJKPi8Rl5
cziP4NjZXVgjONuKp3HV2+Bka6YJHwkRLdDMXgvchRwTL0RhxRRiuhEdKWFbW4Ck0SxSqIkt2k5u
6hQtjz9AIhcd5/rbY30210ZdOqJ6x+69KfsFiVTPn42amNtr24OQFracdHAkwdiDgEQaffcs0tLZ
LYVL4G9a8lWyLudVk21VsBSg6Cd24tCHZFhLGx8BDKbG0/TSaSEby/fRL2emeIzOQb+Xthe+WSa4
EFDUATwvEKcO8EaSBr+Zl6QqPvRRbbSQr5/qyhz66xgdZD4LKXPIfbGyTkqc9yu118MAXi0wwhKQ
oPN7SSPEfO5oIIB8Q/5ogtUgCzPc0q8V4I5RQWS8pOsQYKdv09XJlF6jto14czg9Z/6dlNpv+8wR
bQaMMWxFYhrskVVcIjNXrtuKSbwY2MJgyRxN2bWVhX2rHldkF4ZPK9rjryBYgPteUrCTGuAXg/f4
bUptipZtcPJ73/LsK4+6J1kHOt2H0x9EVV3+LIGlB0Ppvg0rPxE1jY20NkJ3O8hb4bZybYba3H7r
5Z2eUw69GZoFKEWdjO5lQNDNf/jrbLtuLgOQzja/xcEyN9SFrJQv1vxCgQ2L5xY9FMPYGxgGJy9a
rG+gnVDJE6kzxtyBpRS/Rhgz/+N2AWCChA57ZHkqio4AqoaeypMGXQlduihNLQaWvIgTBfZs9vrL
uLAFs29AuJxnGK+JIPXJ9BXdbaCdPMWeN4aVO6jtddan/PNvcCLzhEivb8epGmMPMS+YjRsJU7N7
3pqMrrPKB368vwV/za0hrdcTouZsvLHB0k9lCyPHkCOQWKyore5VPjTPsi2tfSFCN9Gg+c4s8+Sy
fPvpvUinEJGh4AIoGa0p4Z2r7G9QL9TzeEDVIXGn+f5RuZZqThak7HnHP627OYNjLsRwgyVtsPS1
o5lI7a8p3Y/o24+CV3phjpg64ffxglY8Wi0dKTHF5RMPyreYd1SohSXD3lMkCwa3cEdju3px/5aV
10Pe0xjI8HWsvxfK+oW9CeJRvtetxOBRDHs/csmxlSnwRPkfqmFGsIbDR4pUdr1DJLV9QAlbH62C
KqUACPWSmsVhAT7CKmAwbkSLSL/HRRv4vkkJ3FzenBcA3nB2tepww9K4vJhJOQXqr8qRwHixsYFJ
8opUMW4MBvV69w35wIAYNddR5mxab0DimSverJwKOUnJSxQR5KpDII8M5DgISrBxOBNEQj8HntyW
L1OZ3nAiztj68O9w7bL+D1PgLx1AVJTw44Os53t8o9RmT9SFps96KfNpPSYVERa6ej/BIbC+Llfy
5Oam5ORQvCfLhO7qZoNIGY6D0HBbWfWvtqgTakkEPqjDAvTpBO36W29Ak6Ri2MFNOka9zvjkVryU
lgKtSk47fDXU/JtjYypqolKRtCu4Rowb87JCnUvfIDVCcC4uDhEDYLPaa7Tb54A545XwlQ3epSxR
25NEvsdYr8c22y3QKIEE0ZJTobnCNRXIAHJvVCas8ddX+3qcwaD8fIhWfwZacYxDlSx6i7NWlgNQ
ksJP8+FxhgXcoTw8QJtCn+Kge5Ckeqll81JPRDI2PEE3enGiD8qwL2oYM16WJuSSzp4P40fuSdqJ
01YNxIcDhvuko0MapnfBPcZlBs3H97HuRBht+EhzDDHNb4F9+4XrZCR4WtVfhY4eVZpKE5qj6VlA
UbtVVL+rRjYYW7VMs3mRmQ1szXUVSsAH6Z5PMdyis1OHaiioGzKn01YsxfDPehQWVFfRqzqk8KyC
9QtyH5GBGYLzQwi21sLBIJSZIiIjXEkOs1jumQ3kLIe1liOBuVjFecWsldeSSxvYIC1gOIcG/Ypl
eIRe7PLUznrIkwkcoLe+iyiiYppUqlWlVqUz5Radd3TYRQFqSi17P5GxwwOYyTPz1mrHYrdhoBVd
+L7xLFIbmKio5GcDdhgdSTMViVJvDQndi1mX1xig9ASoHPTpf9c18vDPZoGqWs62vBqRq/WhmiRd
k0h1Ub92zPfglA6nlae4BloFOtpxoPT9BY/oSYDQW0ouGA4IczsrCS8/3spZvYUgzV3Cvzs/8eyD
yCc1sQuEb+mtOk49kFLOUGmSuCMX04vL6S2GeZtVVeRiaGf8BpRr6dEEIaTfW7AoB99/rRxjnEuG
gSQZDqTd0jFW2J7HyJUBvRsB+rGVRlBPO4LOM5vtahD1VHkfNoBVLVLdI73fCM0hKZDCkKwnovF1
qbCrYv9Z2Hd6sXzIrL6pWbDmC3suxy3SXjpdfC/VVQayZtI085mj3bCOPdN6Roq7TkVI0Ev9V3br
BRqWd3XA4Z/HYjoC9m9qL8ktk8whK1jXAUeLfRTcVBgTLfHJRhMzZknnopRKvpdbjQD9oQ1OVeVV
9hVjnqy6oAuRM4ceAS50GatluOJ+qZ3N/hxgBumCBP5i98I+MrmG/JuBjiRiGNmpcz4aJYIHAAHc
Tlm/LCRCr5Q+c628Sk0yF4mfuR4F5W+IRhuVzWLVSKmZxI3JzqyuaQcIRM8CnAC0MUwwBK9h1fNR
2rYkDE+uraDDHYk+lwZl2dQit04vhcnuvBAO9I78F80gDGbWh4TY7A+yrvua8myPt9F85gElaXeG
hdP8aq9BZLHlZnCxU55f81OFCRzdwY5oOvw3lL/7u6kahAheO6xpldbv+P0WOXTH+6QPMUqAijmY
c3iW5rHR8vKtL/uh3E64lZP1wKKc4GZqkgCS/PuQLxv8GWCdxsCqMnd6+/BHHMRB4iu145qQlrDM
uo98F2gVakpJ1pP/h87U96OYudx8OOKaOvktu3R3zeVjqiugaNvup0OxvysSgJaebKUYfK5n9tL5
76tmgAzrxd8dy7sm0CUyC4A9D3gowEimTdTym2dsBi00oYqWgu+aICEm/ZBO/zHo2VkiZm4tYNEe
Ns3yWx1YIc8LHOGCwRf32yBs7zGfCIWqfQzvM9e3M5dXefuM6Sy/tmglcGuOVHUE83w1U9sJYhun
/dl9LsKi3PwAh67b1GoKGMU8mNXo5MJNqpQGjVdPKzLmFLheDmqWaRyC3QJs0zCejup+lbmfDNmJ
2yyQsRlEshWSCd01RM2y3u614OhWtWoOFuh8Umzq7L5WshtZDFWYLIGf47/GqQFJYJDNRzI7qCww
99msP7xaJIZYpM9To5ka6PkRu5MVcahc6nsxoxn3tbxOmLSecn2QqAuYrsxrUHJeHi/7DVzQl4JV
XdZVewJySc6p4bxUg8u5W0cq8EKMc9tv3h1eA2whHaqm18BcD03SzBXNL89A2oecRrwL2iAE+lAo
MKvvWSUZ/jjqmJZd0n4lm0oMH4/DSIr8HGYQbbw88bUGpyAJtVeS6texJ3X2hXOjYpWvyfzJj1H0
nqZPwOC+cVgS827qEqggpdiNe9aG9pt8p22kvgXh04tHkkwfYgHfNrWBwKKAGY9Bp9M5Lg8XAy3U
Fkap7aMuhBDZuRXXUrr1pQvHRj66W1Spx/IJEjjNSkyOF9qGSGtDiCPTcEitJlhUFT5G8+q65ckV
aZuBgJ7uYdn64qPqWmCKbUXjz5tBT3uUgNkJe/88HK4zVCew83RzYGHxODi+TQw/a5C6ArWtZwYZ
RwmGDtPWRthk6t32+LJhZtmQYKIXWEVyUceW5pOiN5YJp4uMsNaldupMPIIWghmBFnahdzZjdHiL
Tlwbhd+Re2C9Ol72iTPeTPDaZ52fm1j1zeURoaBvPw4kpMfhbnz7XAD0zPU6y2wlQ08B3n7wRb68
XUzYpnpc+yR2BISC8YaVBSWBAMQ67bBHdHQiUtzDMjzqWqOD6zMhDXMiYanZPeDuXUW5PoqMRGS2
UNifV1Pmg7N8VwkiQpvIJ2/YJeH0gAUKQ31q5dMKZvjin27PB1Enw9s48SKelD7VrURlwdD8XPpM
yXn4w5CUsG1Rdl5hP2N2jX+3JDEx7p5bxKjdsNmYCuzY32Um8ZWN5DUQk/RX8fWBcooK53BOQ9dx
ymidje2rjsWGjGSnmogJemfuavhftflMyrQV06EOeHwJVH2x51Yhf+xAlbQBNT4B90eDIINFIo99
3hZHLS74juLC2LtGeoZqyrS9DbRthrTK7TINPoZEUPb7Zs01sBt+UHfIpTje0d2AUgzJ9ljsJvJY
bg/8f1tgQ71dTsCCfQJZ8W9HTX7eb2WnITljz/xY1fR5YHly1V6NHfRIzf5js4LwuavKEEBm6/Ly
4LkpHyb2OQTSDJDvR06yPnXiFY76LTxf1MeRF8UtHYlUJc31vN57OktFiOQOu+EfHe9obGSlgQ5p
+nfjpmX32xvzRQ82jWWcbvebq6LZfYVb5ALUZATG/4Gg0s9vKklBh8hevZo8G3XA385BOT3k8Caz
ZdWdrEJOdC3Pvey2OZl2E3WiCoalkA3e6lbotWexG19cqZdLKOfzGNjmQi1eSlgBWePxrHImzQvE
S2vUk4f7VOvJ0Ze7g34d14HkuIJvw7hS61LWk4ToK/6wjEQIUSGHOWCZh54DsjTmg0hIvnJNxS0y
93E1RcTfmNFKQ9tcLdf0hZx/x+EsAcsYhcfD5T0kVocCzrmwu3Wv/aSMUyfpe7nGDSd2T0QjtszB
v75c0NSKFH7PKyHJTwb81TWcOSq79a12iyASD053WelwD1vLGGGH0Ryz0R32n7a9shTzweRWWKTY
rqBZdv5EItURrh1/nUpRHFlchEpdk39IuE9UbtQCYOAdz3KY+IhCk+d6RuGph7LKQiW5SO1+AIO3
IUqHvMZRJ4CBk5tiwvF8PHTiFngtVN0nap6E9765fnkcl+5Jl7QvZFi904LqvthF0o8z6D/wVdXz
nHqIxrscZ/8Sm3qr+WMCnfvcsW+pPlw0NAny/YNCOozky1l7DA+CAUVeCQpxEz0FfqV0xr97IHDA
bA8hXjWKhqqU04uUAI0u7GP3uc8RCSTJTKM+s08H7GPdrsIlBf1RZ9/KNFDlWqe7iMTcDF28SqK+
SdQgttyydCb0i7pn6XrXFaaKur0rWaA9M3TH8oqzPG0mIfAX2zeZjQkSfUrEwtPqxPpDWGHcv5li
9BMPLccx1RKDD8w2KlkqzGfn6dB+GRf+/JPNztJw89RbyXTRtkDVU1w2qE9/Q/rXPKxrT2YDr4Yd
PowLrngXwUDGBWN10MlSw20PSSFDbQ0nPM5VTLvpNwPQ6rID/hyrx7qk003XIx19NYIX0TOJEjXW
umnb/AYKKKrpPdzqyUm5sCeIvXNFii6jnvT2c3CKZjYt0cKO93oNqZ5kC8BwbHFNgELREbeQhyCZ
YLExDJqFu3BFoHECwkc46lspDtBO6hJ/lThdqLDp8lSki5DHKw58Y+QyUGeHXaed/o3UAmoo69ED
TBZy4SWz+tQo8SALKf8wZY1NOxeBHSd1fvBZ1sDqi9fortsKD47HEnJEL/qPbLIGLO8vZ2cQUfiC
GLBYvFhSOaipSfNmZotJl38mB0fODdN296Ofx1z/iPrKfaM8ntfEUv7QvzM5Wmi4JcjMyX12elPa
XZoFs/BgbcK4pHsA1mOTSIv7tYEZLwvMO45bAiDtrlpJQ5t6wK72JhPzyfVYKQvVisdlz3XEisGt
uRFwoFCCJph1+R+P1lHf7jeyvw6Ypru8OYdLxx0M7qVAiRVrmNnmLZ4zYNT2lDUSRQrXVnrXYKKQ
KaGD8PIE8fIrAvSeHsEN+qXVLHG9fvRHcdOhEfiiQWLlivjfMc6ZIg5Gmc2M0KiqE43Id0CJ27Tk
SrdPX6M8QviBoVPNDrvtPVYdSZkmZSr7cpYRIa+ijG4PkRsk5sG3qSgTK+5k3jj8Db6ShGg9/sVL
uzHq33irEthfchzZ/LrZ0yS0BKW3LzdGkGurx4acCk4IJFP6OV+Dg4yZiYRU15TE7UllV4zY1X20
3r+dXFxuqyRrxqXRt3vd0mGq5n03Cn+ZqMBNp9UKyTzScfeYnj3ZzDYDGnLw7gDY6UKJWqxdAbbx
+yAgM/cYCuUoiUcJ1Yf8RIx3U44DLK72yL6FZOo9ygM2yoH5NlGrvQkCJzINha1kk4I6QhJeX4Q6
Spr6geRFcelNhNiGse+53aLzM3G8z+wCYHEyO6eUu3NSuyxY8CkbI38uulYJYDetL2f+PoaWV/kA
B2VOse/PwD8u//qS4svjnkfEdFaXhqioSnH+v2gHiF5LQTpQE/w14MQiDLXZIaqf6d/AnGbVW3Sf
9laFIpFH22N0KLCr1r6/7j+OBzuhCtc35KcbVPOIpjpKrdRvdccoJ2BCNhEHZ1lmBjnqB0HCxoct
Mm7tPRE61Hefz59/uD+0WwEEPKW4ooTl7ggS2vhGXCF7t+DmcFA4Ooj/v1BmCTRXs8kdUWxQii9i
wu1gBfEXH2UVoTSb5HuAlxhNcfAuYlcgl+YrJ4YranH8GiSxjhf6WHrLvewjGvtSBpwStJnseHoT
GmV3j9Y+mGmdZlM/pwH3AfTIlLdD/BzL5J6DEM7mccliwGYMAZo/y4SbNQw4v1AlsHKIAL9r1ge2
9nBcaRFqZ0fmdkqWhf1D633wd0dIX0MEqyz/ieYgPtxiwV3h5HUPO0P+He9Z1f4G84jXo2PfHm0m
EQMzJ2SG3MvMh5V8Y2qTMpPymvPv2SLku+L478bemBkf+oiOE6LzJ64AKi0ePHJAFgQBPwIlmRTj
c7RPAIA4luiSKlETlr12b6Z14ns6Q+QvT3J9GtEZKw0mj7wG9Rx9DiEtNIRXp/aK668KyHEd/hKu
uUFV0OEJVpppJVIgH67GWoMr5koftqI4u+GOEqfB3wb0o1uzyl5LZ71bLxL05xCS7Idr/6fhA9cu
w2KZUTJhdgCObufjlslQiFH34tg5ptHndr358vp7QBX6bZPG0IClRd0mNFCLONRWQvny/qjKL5OL
oGLmlLsah0Q9Uak7p9BmR/nGDYZMQfZS+npxwyxSMDJOipgNYimIKE+kq36wKnYqRrsl7TRu5l/A
6a+dGuRFkfCyx2SeC6Mlni8km8LL2U1JYPOQfj2nQezOybVKuzCO95qi0OTYa9yDFd9VyG1xb3GF
z2b2bXb6wDDVmxUZdMzhqDzII2AaRS/tWVZ1VAU1Y97lL+wW9a7SzgqTYHotAO/qxjqq9wqIozcK
ggYBzbnpnXXWez+YCY78YygRWfhPp9bypQ4plQv4ZoiaVxSZU/bdUT6z3hA/5CvKHVKE5Mvj5qLv
1Steh/uKG2mpTnwbbuAKs7xDSSJRwRNze1b6HLjzOTfybtd/us0g6ZGDqU6k/bvjEfuPtkdnH7G6
Rp4hjcs5dCWkJv2gJRs5PbUX31lvM2ajm76G04y7Jcx7tfmYyUeskDYgpHWTOLZ3tRb2fZI42ul7
LOSVrtS18OTlLDi9iNOEmtH3gc5uLWcLT3BmceL50t5DfHYJFHPhCoWTk6uTrc5x2NhjZKWj/Eg1
8awTOoYKKrEIJk1QiXqqiR1wD4xZh5d2It9pi1mxAu0OWo3sGU56v2tKsfON1E2iep9gLybP7pYq
Q99l9PFtWf5OMNfe2T2GU35ihSMA6fCaC7jL5ISLeKt4ec1/fkdwdviC/XVyEDCPR0JZoVM0oOU+
MZIjeWGWwbKJh42rDR6XT5/WGXKyURdjAgHAugYUaABtJbHkh+xP8m54myX7DpSpOjUJL7kLrVtL
HC/5JisonkV9P6FdATD4yyaVwMuR4ltRxUp+Y5P5lfviD0Q8K6f5M4l4Q+yJMV0GjA6vGVvx8UHP
4XNiXnZAFLMbiQAH33aiWPWW19rMzyBaGeVNGSx4eu+fyimYHYNbennyZqOmd8DIFL7GrJLt+z/o
h0cgjO/VcIWjMZT07n18Q8k5QLcPqODCLXtlNvU5CdLo2at0ycoQm7tX1NRo1hxBhH62H1yrFIDg
hby6sdF0CYbNdfI2EOTgQD+cHu1GRTf97BBUHkfYV2PLV6YkUvhaCkXzBurbDGR4IuzI71APR+bH
Zdv1UlBdgJ76OJih93zbotfL2gqj2bp9mTZLwlHIeMlliwKtmV3ezky3NAYIy2cQhwNlCg517rW6
tg1aPz/EBMU55ljoUDLQDTizEsvzUXJThAQzq6yrS4PFMJXsMwb1K/VJ72GFz5PWoAOTM7EcP23G
sHaX0kVnKynUvR/qGqBbrYXmXA9e0/ljwS9y3YL80PyN7TOrIVr3WyySrRPSMXtSM9YuyfS9yYcU
NRbNBt8JaZkRZ4EM3sbNNMThJ7dBNbop/Gu1cNadHQ00hmS9LVtYApxd3NpnGaby5kyoPHu+r6Qi
rdoeiYMhFDA28q8yF1lg4lHel2wQj4GTeArq2NxrVJPz/+BwqBNyPxFeyVPeagwTgj7eXp4AHJs7
fVxYTBOQfei/sd4K9mSWSt3FDAk1u9jp56SLBegTJXmW6IYF0uA7l+kntckYNPam9U3ACahwo7rO
OtV/RPnauVOLc3xhsLmfxTwyXU2KkO8xvHf3J7R41f14WY/637cPvGdDqEE3TEwU45noXzWQtPPT
qRNqHemGFgWXKwjXdrQ+BYCu3kaozybq8nSFR45PN3BojHmp/Agol/X/+uUmlBY6pDqjhSh21cso
Vgv5IqFIqk6OdX/88zM6RbyPYaaeXt0JvHb4kWOuRPgF5PrLHmi7B/8DEGulye/NdQdt9nF63oEx
eVfV01pqpj0rP9c3CIe6n3ow+BNhwkdafvbftqLQO4NLppbt6WKrnu9Oulx/di4wmVxUxSvKOXNd
A4oZXr/bM85HyiDsLcW+9jI71FVNpAErSDAg+sVvGX6Tu7wkhVQ1YV7f1cvQu7dH7VxwjqpexKCd
zT1Ijzc1FQ7u2FDdeka3dy8+CfEl0Qgnt5eTeTNdSvKsyMjCaVzAe62qD3GrLc6WbX9neUoVwt7W
+ZcG6ZItqAusy7I/Eur1R6ShFLRGfexmcRwc8KQ4496Xg1ifoL/GMHYBAtbDI6DH3lqNhOwukMYc
itJVKsWiVimkoiup2ALAIJEV+WSXqrK9Wc82LhTYV8/G1ruS4pnfZdT0kEfPmAwBLBblJa/QMuvW
fsHpFft2XEgV1u/OeYfsuyPgeHjsm37mDcNQygEf9pG9efiG+MjFBZKEjYMNta/UKGj4qw6iSwgG
AoYwGhcQUwKxcFdSSr9fiEi4raDgtPkQCQyIurHJF3E2b4A4EhKCm+skn5Lb5+PXzmR6TCy9+dAR
9C0pFOc2LqeKDpscaVaXN5zcCQf/G7Nh9Jl3Abj+ICyGAbHm3QYVTQyU4iC5kvjKmEgS8m1xuoDe
6dWVKr1FoBV+iw8u3ZlFtVyWIDUgrn8z+zzF+Pixd3xekoc4IRmcQZCxk8RE/rcv5Hn0Srhf0EDx
3sV2MAUE+D/awlDKhEK6pmYFn1rBpl7dFxLHCBupCMISX/f5ciQLQqD5+0EHAf00uotaHiqFXa5o
o5bmO3HfoShzrWnJD2N6zcgtMr0Wj3hyfjGEK1aJaolbTNTG/IZej8nkTCE2pz71/2Q02aNjtVqK
5eNO3XehKxzysjPnpg0/ZNy4tR0uKXsuEdlwqApjR52JD4tCtMdjKqM43VFBd1kd7iZgr4S8cite
LrH1hWpAzOklQnm7+dVqoBsHi2/EU/mSTUF4o9rqtTgnLdaiAUJf75AgCab1kTgyfNaYgiHXTv8s
GoSS3kmU/McSHvrljq0GYKP1Xhl/j/K+SYwcC1K88q86eC82QNc+m7RJgEl9PF4T3GjCLf2gL7Sz
fxzjkoRzd0zHT71SMxqnlTEgCSbpZV2/7P9FfqQuZmkqom+cfkanW25Cmp5QA/ToeQ866rHU2S7L
19+Sh/afNEkZbmOtiqk7ZCnCuVQpmMgmYg7rqJwL32aWgXrKhQZWWeQ7q5WjwZByxPdWt7Dzeiqj
WAR8kjUQAyyCd7F1Ce1fhLs/7eKzzIRcSGBxRSLp3seemC9wsztZPo1MoAN0u5oNK1+4xb+Fd1Bj
k4cqJ9NcLR0jm2B5kiP/uhhtYOZ1AqdvhydHYuDZD4si3GBNO+fPMUgJ60K5ai3Vytli7urT/TBs
5dpd62/p4As9aJTexeSzG5qgjC8UGZ1HVxcrJmurYKCSnTeKb44Ps/7AJIbqvWUeuNw7dV8Le8vJ
7JpCLEJVjIlicHL7m/iwq2IBYNUQIXg/fbh2ssnTJJnnjtVI5OhAh9yqrRNwmnLbhL/k+F1lwlwX
FtZ+MDpPzsRCiYnlwTYcabO0Mv1lKLkLVR7tS2Tu3lt5cfPUEhW3JZnhN8r8HQ+ZppX8xJRgOz26
NIEDoZL/fWdO5nAcCvtkFftHUXNDc1rpD9llVrQhJlZcNBqRR7liT4vC3VjIj2kPvTrf1OXXbQ+H
GzwtKR4JTtkTFG+NaxrUeZG2GrlqUQl37L/JZULt8XRl5A8KiJHGv3kucHUd4aOFT20pWRWqcow1
tJbufYtrTgrrSdLd5N++eBXZezdsxf4m0qojeUHMalkBNlVbGUUn1n2Qck7e+V6hC9NtrgKj7GXO
e018INhGaKjOQK3gYkT5knwLm8QbNWiqzTIGgBq/iIUnCoLQghmx5ZneEctZrtZCv8myUl8o75kF
g5Ot0t51Y1eSvbk5LA96yTvT2n/hBR/42uAqAu8OxXE51urqimE7kDl24RCpsM5ycG9CHRTOMkaR
/vOxWSle/goYSWa12N55/Ks3+fnJPBPGRpRTBpQttOZoByEpatvc+BJ8c5rKBtI/OtXI4aAHEwlS
2ljfaNkheJZQVsplV99flDr8kOOYY976HxV7GOdVFMDAVoIdAmV02KyOJM60Wv2r9nr0ATpznE/I
99H6b7f86S32HZTHNCZxUjV7U3QWfEJajy4GDWC6WdmurktmwHYwANSWjhVmWbUeI3rAH+NfKyhj
js2ytGGRrITRZSPaZsX27ZveotPrj2M/mO730tY9niv9eLPmEevMpuTRaKFTxfvWw0EQnvvYWDx9
y3K87vOK5Ot7kGkunn258Qal+e+ZBLaZOqEujyAQPi58WJYfTet9YKX2+6dNixFbvA3Czxc+xSw0
jfOUbZ/uzrpJn3CPC1R4J8XO/zZE7QC7aLg4qGYAPCGUzTkobEnH11v5ZjVnCdh4xCZHad+TBfpE
KZkRmoOaXDQZKH5woiD1wHY8np1xOVmbXr400JuEBlyaKamSlEPO68OdA5uUzw4zRdxN0b1CMNck
Zn5kQ7qvSN5l/BVV9RpGdWNjtGXXCBV7LLrAG3M2lWC2LnCVhzOZpp0vSKRNZ8i/gLBEVLtdunXv
53M5ml4RCVJARRmKHI4Rsob3By140Go0o6TI0y4sUZL7ZzqfJd5Wm4/xdFLzzWUD2ljVObFlAjH2
xMttOtCRLypUZ6ujNbD9Va+cGpLSe+vB/MnNmI/QsW7Zfsb8Q1o6NOmLJzabqAegG7GYIqYS6ZUf
p4ZyMHuSs2E/fo+Yx9bQmLLr7+q1EMtVmh2Zv4XWyEuAnnTUMogrRfbBEqPRaML4KZzUNF5m2K+v
YIAAzYzanvcUR9qxRVB9es9iJhOud74HYcip6hOhu7ENknFScs4u3fvCg6HWkiuW6zqyGQ3qxapk
0dmXU6O/CmLsogneh6AssZJrvGrlYqgfpyHh2RHDlDS15ccHpa3d9GQhfcH+vn3TiYYFVEuff1PO
NBwzKmdJUeT8O+PeMVDYpG5oQVpMSFdu4Q9BNUl72NfSTOroD+Yf0mJ9NqLbgwjOTmtAH1XEL4sH
hV39Hg6YhQzz1bRabN0M6bchemwoucx4Or/oX/5Nq8o3AepbNGmHsuwtXv8FUkVOFNgwZOUDpXhU
s29ALAf7CwEGsQOeq9mIpEdsZwqZP04Njxzqv/HKQPU5555h8T2fZ1O7Wl9PxjP4hYKQdyWpSAwu
T7OujVq7T5rKYUA6+coTEshNZSebRjwMkeDuXlhHxahBc78awYiCOSOn2Hehgais2BU42D7ggPbD
x8mNeLOObohszwf0zsa4K50V9ohIzs0nf2pxbZ8WQUUMAcPFDDsKCK0att4uP5lKEBgeY50+uJdM
qRYIzunvB7aMAah9+GLLIiikJ4LdhkYvKkbpSC6djQdLxW1m3hjAOnp2a//v/WD5t4ThlYO3xD5m
mPdMp7egSPGZ3AS+dmq1PrRIPunaFRO35GCqQ9N6OnNj7MBKAMX6rd8mySa1Us9m5dFKALaYWFY4
lFjfGO9A9v1pXfUjTwWAmPDQwNuNf848enrYJEV8SBd9zUs53PHLBFYiYkrN6SJsfQ4RUt+D3Xr2
MOdVJBXSkWkMX0mOZ1d6XsOEwwRxJWyYJq7orFjYVJVjbmFKVAbGFTvDCxZZJdjrNdnGRunUa0jR
6YV8nbtMUy93+iKKAr5lB6fuV1mAgIrYt5382WU/e+mcafd3Up5TP+xR57aTjTEKzMCwNgbZkb6D
a+3H0NKsfPZXpTwawUo14oh5TboNoYaG/6ULHiYXEOvDUTjCKc0Vu1bUTvjkehAekPNR23mFHn+X
hzpIshemmMsKmrcuaJRMJVsmRXmtoEdRPGBLdolfm73SrdR71E/5GIqUK15JjdBABhhESD+ZMnWR
oChTTPupXqhjdJTzRt3P0h+SVSUg9mhKyiep8sb/5fLX3456a14TZeVCWCepO3blJgwJ6bcUTCRZ
7k3L5J6Fs61lGAwzXXVSWXZvhMYEk4mCG2l7xY6I9yUInxnuSfntvFfUzqfdOZlgikHqcqIW+xCK
ParcRdgULjf5Z3me6ALFifQJnvcMz2IJULyT19W9bL/xFpnej0qesPS3n5Y4HvU36sceIznn0p0Y
GKpu1z48Egd/cbr5Vl5YdbtZ7uBk9xNJq2izpEGQtyQh0DSFSQtsUaJ6bNHnveKvATvZXsWZvhgb
fBEF/oNW8frPckMAYHQT7bnzD9KDnRSAzL2GDTNqEkW2OmMqiahVIvu2QYW2YYnKEXriHLhxRvEl
Wr2mfrqYmy9csMh95pci5LWiQMV/utvaxQRnrE3NbFo3CpWcpIm3pGMXELS3HFAvWApv66oB1DTC
NHIuaGP6HDDW9AtpEOJOfBnSGhCpQmlR0u6mSRxlQN/rRRJiJd6MGYzQNBmL1cN9MbY8MMH+C8SQ
6bYNfDjaRTLDkwrsKYSbCH1GSY4i5QCAS4kJ9ToRvyjjYiNRM5Scy0dyzp7u8TCb+bQczEMG3Iww
Q2T7gqLEwrcD832FGMxXjTvRp0tt3va5J9ZBVSNKDJ3KMxT7gEsvDUO2r4sFKSEfqx31lZxGhHGd
6PLyr8xqiLpVKUflq/GUBRrFoibPn9sAGEw8I/lNHdrqqoZUiu2HfjJPhjVn5Yp0rb9SAhqf7tTQ
AUgFbq263UkpJTxLTJYCrXrmI4ufgG8Yfbu2vYCjgA6RhNoNUZQ+o1ciKRLqarqAxNdFsRN3s6G6
wYYvtmbKtInjCFMJdMYBVUhdf70Jb0/+bXSibgNt6Dn1BpCuIKzWp/GvYHvI4t9i9jyuVyJQGQv4
Bj1eZC74g22Hl9+EUQfLwh7zN1lO0RNql6LRLd54MUFQI5809ftItfZPNiYXCn8NLdAnPZaM6xRj
9PWE2QBjjy0Hc8bVy3nm+RGa78q6C/0LU8fxKBQYji7yHOu6EQANOy6HACECerT0TooEVwLne2BY
/VMGJqWo33gEo8mLi/PASX2Njhq4Aplpi5msNROnxCa4pIjHf5lSDB2cXysGKHnBEABidd0AaHpd
ZCA0/M4Wz9JL5k6ug0ydZs9DkOOHpAGKbaB4RQ7CQYqm/FEa4neeV8VYxkLgaWKa7p4wacPDjcxS
niOSX+A//y2DqS2tHL5ENuuuXVLj78l43H5xAD716BEHbCdJDRt2tioAfeKKwKr8CdZyqHdhv2qK
SX5ZRCoDRuZo9O5Y+PjUWTNUXhJomrN1IZ3kM7JjSGX/hYEcA0aXixVKr22VIlYk1oaAOoc4wwsl
lLd39P7HU90izqpKZV35TOtIVrGRbGjMWh4W/Ivhqjh3vt+LHZ43BjOfssnCzRrskyjrWe9VCjuP
A0XFgBSfFy2C8gsQ4kBwhcGt6HcMuKyGphw7s7QM89+umiiKfkGVR077MdYvopjYZ2+LL8nBQxDZ
tFjPRWAKkm7ZBh8SuJdsO021r2gbkpZp5QWPsdCsfJWrBqHqANcJKNACTdOcr/ICXhMFAHyEnPdJ
ErYGjKdrmsDs3NrO9MXPuMUf3AzCNcZPr3Jmpl49uPFFBIjosqetqlASe9fA4kDGeJtW1U0Iwy6B
ZOAe1mGPnrGnsjNOp2RxYpTaE9YPlv+frPLbEinwcqgH5UJZlMJrTroIrAgKlW4aqzEeeoPAsv4U
VouhYma/mg7sM3Sf+wYqn6nhRADYVd3na/tw9YmSWp2MvHVRPnrydy+aAVEuXdl1TlWx7AhOht/6
evTJ1iYpAC0tegkiVPBGVBEs9Vyx8LIVnKuXQM2/yzuiRjF1/BPoYErubYodZ7aeupMgUY3rgY8o
mo1MjD7vEoWZpMlRt8hiW3eJv7bBDgk7UtKqzzvBnhdOXAfh/qWOz8u4FalcLc3UU3fCZLA0+XCh
e5EDf0y1qB+RcWlwQ3V03huTWgZNSiMgebqrbsD75qxOpLjfBtahKolcpg6iZDB7JVidgGMrNnQj
O3nt7YEP+EBJTOiylS0nINHNFNHS73pR2T5Wraf9nJTUOTtSX+sUFnyg0nx/VRzi2SrBi7lDoFnk
m2QW/+D8uGJjoiVn8D42llAG8pyDc+51CFZ3gM2tijKy9CW2yi8TTCIJJuu7Vre0SInnzyHZZ2eq
6dh/6G5xyZxMbE5XY4PPx9+XbMoEFotDIMil3pnxH84qxz5ETeygCB/mx9E095BufkwlRredfnhR
7+0ehMmg10AdgGtnhp062Fg4euh6nefmnI/xbNqiJ/GpJSxDFCowJClksyGSSSiaQiDJqIXgyBe7
eJjqfFrmQO0XM53KLNcAcKIntQ06M5yd2M/5DvzkbvevuioT4PgulE7QuaszyitoexMhpreAupc2
Cah00mwjQ25Ak64ngvBYc9/Js2NCmiL5PsJU0iuNtRcxT6mWbfCZDP6X65KBrqzi3/FYdQzdc9Xf
aECbD9W5s6/DT1uXwUFZ07w4auWkv6hvvL1MCMaWXFl9r2ofQlWFJg7vFkbWlhYwX0bak1YhWSns
3qBBrDeh6RXKNiEBr2aiuyT5pqNqKrQvHV33mccfDbvCUH9bNtLDYWi7cYoZSPpVhWKJBMegvjNV
RT8yqM06Cejpv37UXE1gy2cI9yBHuAG1Lo4RcrM63g/fbRmTU4kSQkbFw/byog3v+2+Sm7aEEkBq
QVKy4YRe+ervV66h9KMsCsTToQtpMyXr5G7ok1Tp+0RTwhzDHtyz1QD8Wr6OqKh9muoX7r5D/WBq
EWvduCQ8Fhpjb28FyHiXSoV78YCphs5R9Ustt/JrQ+na5vrwqP0aRPz6c3TzKHKdPdX7XceMjen9
GGCIa4vIL5YerKY3b9+IUzkcwOphsC6uN4NhVS/uWCkfQiBWlfIGcTOFt6O3Zym1qbmvqTj3kypB
xRMoqN/wKPinUd5XCynkWOAMYXvjst07JvKXAChk3EOuVgemNXNo+lZ0I4fQrotMYazZAj3ImNUK
0SE/NkmZBA1UCXOZAOZsfYDIySxEU0Kb4LAmf61rucoTW5zGaoEZfOQgjUw7dmu544gENp293SV0
ez/R+keSU8AiSJRpTkQyyKyuWyzpeXSA8c3HhiBeRRMOWASoUqZpwEG0AfzGGQzUmuL28vpd9TBi
HBhKlEiINuQFF56jQ6FQ5PXgm1xNdC0KUGr8TElJLCZejTMF6foGmIsnc+PIO/nU71hnv7wkZmqJ
c8b1Ru74btK7DfljqfOnNlQkEKc7dcu/WD5SNPgbig0ChPHAPbgLj8eIsmomgx1KQ2EUD9mHpgjo
8Q0+x+NTHvsC6pMNnN+6uzvXsyQKRpKhOGAEEQOE8sY8vQJTTKn/jzLN7RX+oe8eYEgyGUH0Gjin
Ke26DjeTGuIfaYDkoIrrtqeZISEYkX5VH3Kq3q0d7C2VbaX0cJh5JsLnXT34fEo38CbawDXRt5XV
1JJwBPrZBdKFs09TdjRYCWcVXaPz2M/njDZqQ5LGA69tLyaaQ2vpg9BZ7ALVkO8xs8MwfScJeEsJ
MRmyD+Dx4DPc3EW/mGNuSgx/lMyDfsFLRD/F6gSAF5EeRzMpLT2Z20r4F5eKvg/Vxb0askMH64kY
7cd86G47tNiTDKfekf83TmWZmWETkbpUccTOzCff0vYacgEDLdSWuOPMms75bsTBdRvl4Ie9IkY9
wwNqYdxt1Ivycm73jZYB3l8KPZyrf9ciXx42ZvUY+3DJxxAwF8x7hhlsgy2xJyI0hLW9RBj+dAKg
tydLQ2ixPyHw/ZCc3VcjHOskYioc9iIyaaFTUev3erOCUeks7wZJvUCuV/MZglYw1bd3exmKZFYI
wvqQVQXTvi/f1/ykPY+PpxqkCUROU2p5aeuBNvis7+yY7DGPbx71jG91frjBnM2fBtxmvSp16Hbq
waqLOzryuScQmL0NV1qB74frGFMwawOQWTbsqdAHzBD19tuE/zY76lc3wcxZ2Y6zlP021qR8yQ6V
2Fi+hvim6BhOeL+fIYTC2lBj3Q5JakOaqvsc27Th6Vam7zsDlppUzJQkk0gRrmo5spTz6styWzkZ
DDDgnClG3YKeCjIRbBKJM3PZrztcfAxrpuSrmpAG+IntB+W1hXN8v+9R3NL2UKsyHyO4qNrYmyyH
1xkc6OAyjpDj4v8+ucxyLExb3Zyd+Eg1rc/+PwohtpLkxbKn6UQfte0tEPinbvv3NbO3imGeyrry
fNf6lTe4tG5ZGsAwyKi55JzDGHMrjENRDs+C/aD5b1QDomPlWUxTCVqaKfebFFGFD400xZ1N+UaU
mJWtQbgNP6xcYIGZCZgeG1Qk3K6x+IvO8vmELqXEC72g7pZL1Ab6D7SzOTwOQICp/+0IucoLPO/h
oos0TrjjNk8JRCIPeavNIpB4vAcnVg+3TquKZLL7jwcuwpaPZAPcMzpAMtCf+eugVs0AccYDJf35
hoFldrC7j9rX5zJdb2DIcFrvhvZD1jsqz5Y8xT4HNBmpTshosuQWsi51M26iGpdY8OttKfSxJnpR
LQAEB3IJpznk2YZVxh1tRqENLxiV3eH6FcMsJsqHntiwOVexjXZnu/60s1CPU0FCEUHFmCC+IOoM
oooMO1RGrZU6UH71DjBdiu70/dip2b7YT0nrSkKgn3430Po2V7sK3wTWDDSJNW4qw8UYXPpxxvJ5
OqlvgeVwv4CQMXFsPL6KYqPjQYYtIQC85hEUYRhJEFRJaT2GiIpUgsGDB6hWHhsacNrSe5998dri
ZnbMs5Gw330UlQf5D0yUbDxQpLH5IH4Ax7KeKe9ocqeqD8WBGYFrYCs7ebyfcmeGNpMsj5tXrl66
IV7yAw6a+YGNjjMlKadfcOT2Lh/tWKxu+Q2VsawVvMI8Dtzjp5sOv+9bGpwkQZrsFB2aocOqv+ng
bGjHKicdL6Jmb55gdb61tSQ4XzOzruh/kvFX87/uCYt9RuSXHDqW2vBjRQhMdNkDRgtTS/Eu+93+
YlYVrst9aHOacIJqw+CUSyKX+Y1EdJT1thqGV/y+AT9w885uzRcFv1+zXwecNL0iaGOO/yG08XKK
3oJ+bOXpCsRsWR4v0Oj2cxWdHsp+QZ4oSy0Di4LGY3z47nJq3bgbykdt78XMFRRK9rWdACJhvdOb
E/VNHu3jjPskQhczLJG9S9pwwaz8TosJuJz63o7qGcd6s8s1v/8LvqYG5o3zJOJZYAyWQrJkcKic
eGAAf8b/qTsESLNYIhgek3fDXgWhexpMlkPj6fhZpyGTUvSkKxQkJjQTJXP4kIftPTMui+eX3Q02
v7ccojhHJbZvFisFrpTrbiRo/guqIv2+ykVH76ToDUj9Sb0kqMdG0GEBaXnXbAaJDRS/MNxPTbhG
lMLYIXN0km+Vkq+3/VeywUA8145lJV4LvNoiEk7HH+uityj6RdpFxjtD1eR2y67TA4yHLY3y6c0n
WxwTfYCw9CD9r81lXb64ukOGfgsHbP6xaMSO8aXm5lOn1VgL02NshZ5q64qnzBO4dgS2vGiz/3+G
i4ibo2Vui5BfURWenZmeogwCA+rNVqnv8k5XKH1KMdfp1zn5LLYdTIIm1o8PmL/wkjUOMDDsMfQm
f1a4up1iXY1tAausWNpROtKNlnI/x9nmWcZHL7LfgInZL1lbl6CdAGkwqifVFlrXrjL0NNMB71D/
z0k297NOTpaBte3zzIzJwoWODJlnCwQZYRgdmjjnq7QpR+Mix97Z18e5wlC3Kimbc70jSrbtDwPb
V9//W6AwpZOZc7qp+RKB5tzWzjqSFIsjnUzcaa8jtyXoCY3ZM4/w6LHDSJZ1MiPZ8BF0phmXztAM
QzmLtG91bGIkMqrerE6GbQNg/s3thC5CS1KF+zsAvtiM2nlFPAx0cuuiO4VEo97ZjxXungVEEkMp
SEX3TcSL/z6dNnGBVlzu7yhizYNgE8Fu3XF2Sm2e78sS+CntBZDJKfim9pe+0Inh5sR3PJnJgpg6
lKpJFhW36ExeTJGllYrrLgArtuGYc/FsXkid3w5E//0PNtj6esapZJsc/aQ8ZjFooTHfBr/lVj3H
K5vwJuPvHNsMqWbH9HFExJFel5EZ9acCoyUoYGoNShWRNYdumApxp6II1lqFDFBelIGEVFaJoz0x
PawtuoHiVMZFyciySadQpvz1I+Gc0bKnzbinht4kGgguc0jCOHW2tOXrhJFCDDjbNvyw2DvNA7uQ
BlK2oHhd8GI/LQtxUIiwUtUHwftuVz9vX8JG+nVOmwgJbGzFalAYyaa+gDsAIbOJYBP992EvomEv
dZjYXsIES/UdehjEB1Jmtk15AgBmz5+PWZnZkf5JD7EkwJZddg6hgX4+Rs2YQJMwemPzGCNYvwyR
/zqMp2qInK+JpnR+4Ejhed8MNJLRp2eK7jyVAiRuLzXqLEYRoT85AbZodsB8iHIvjEhEfQgVzbP+
lNiUHgYTz8nfTyYh9NVaRGPHzXAsOhLMvp68h6Aq019N6T79qKbzxzV4WgywuX+Z3Si6MpFLVLgb
pCI3Og2cNA0AefWaneXYYLEkzk7wnOG7vbIzUla+J60z64N/ddqbG7tXaX+xhOHIlvWiRu01oEdj
jj/47XEM5CFt0j6vxAaYmFw7j0m+LeOVbPX86pG7XkneAn9LTJnM1DXG8ViCg/AETMyPXIyyI7yk
R8pU0TG1U3br2vwLCVNaRZSg8YL+JQxIIKJyva8V6/KNNl3JrtvxSx47XJ3LxqUvyvKlN6ezgGDP
w5lMXVraZnblXo5UTp1EJzH7SGuusLmkJLSKp3wph34XBH2FNzEYnjsztJtD0KYzmoRlNLskeKy8
lWdxNMXoT0cAnkO15A/v2Aqi9e+KnmqLwtsvlWngNeUY2YtyW41bBxgLzBOlNA6LhANClqi9YGR1
qBxQE9WNV31lsWBgd/G/QxBlGemzFOtDRwL/KOVJR8IWoYd6cGtk+qnWgsXclGYmSGFFnSs9BFVQ
bQGOG2gxH/FpX+5XHp239mmGAfWtdD0F8ibVchEX+5J83r81+M5C05YIaV7EVZ5CaSe0baKhWJi7
+cHL+VtjEz50VLMQdHRsfdjMrmG/n3V0ekA3YEkYepWc/mbVmHBWcallrXspU9ZsrFvoxR6uK4Ak
BL0LGNrf2+unWsKvt6AffR9JMxwFEe0pcfP2Y0HcnISzbtURdT9M0dH2iJl7rTaN+ARFw+y3x/nX
+2lD6eYpTKA2Sjq6y2GONTE7771Cp7uP3JY/f1p869NS3pJTRu6xaaw2dBER+W93aWQJr1Y6i76j
Bt5a2KLsb98mxxDY1mqIx4GIAz/3wmLKb6NOcI97Fhwj+hZwn32AnBNWXtyU23m1QttrA3T1K7Q5
+HJTMoVOrQFagXhojKDSmFLmhGTy5WI0gbd99+mudXrlbxafPcl2zhyLL8OiBOvQykZfxCYpxpnY
l42sAl4ccdB8ZkHsznG6FE7hyVF0CsZlOrsKUXKkev8bicMduyq39KPFuySFkyPklwvVo/8Ygzo4
Ps0F3zJ3s7k2H+tyOWYGhiMzuo1Bj7cTfNj+8H3EIG/XHdUxmL6gaeOsK/I0q275EBzGiCtpoYEq
2lLK06B/FpLItTHV03kvxrPslBSzsDIpcXqpZTTQPxMpqqKgPywEINl0/WxXNRgIQe/Lf1PVlsXR
6bt2QxeLOh8RaGna7L1R+fbkYcmopreMWFLPJSGTB/0nAb2/Pclt7awCKpw8bT8GW5TZw/XdLsuw
woThQmCW1xqplaPAZeJzaYdzM6SuE2zI34l/J4mKUj1V3/4ZX897y0NAwZS+Dy1FfS6R5Hf4Jrqw
KK+f4Z1u6PYRT4gG9oZoWOMOl4h6UuCM6F940uBEaLstZumuqCFc0X/eT0K/+q121othZB+FRyno
YVOuwDOIz2WGCpeuILfKbv5Mx/zCsiaSdrCntvG/mcAJ6W+WjdbNIU9oY6UspCJxgBi+k6yjIkga
L0Iw4vaFazK/slob0egyOEiTEdY0alQZs5whoUs6D3kiuQJrRAZtoNct47Bz1xG6kVzpSYsap9pA
8tOdmEpiseQTZMYH9wJUgY2aX9EFddbmsrYANbgXjFQuv3RVVHJvy/G3dmokWVJjrPzH02EJpcbk
d0LFwHPhHxRXkkrsi6m6dVwYhdy7dmiJhCr2JbLiEQdFRQmdPUUS/qkvqmJrTld3h9E1wAj5PkfX
2JSahnJcNudAttSxdLBwhH8DDbKmqKMZqDhxQWp4UxYJ/55YBS2yzCUJZn563EHvARe1CPqEFFvC
4haWdcE/1RAG5VvooZh5PtMmZCGhTkqwqjwTmbFA4TfbgrvUuizygAseeUpAbpFCMPo5Bey3cwZ2
yplXG8Qo1uFTLX2+XQHPIUhJw2x4bOsiMFsyeexPtm7gbcoL7F1meROmo46Z3FYNXoHf0KmieqUU
vG3qa1BO9KH+yyYmprkUwmJe/2vWJmDMFzpw5Qua+Ui0aWrv7K+NlcabxpOj5xDzrUDcvaX9FX1F
SgyU7HRnpMdi94LLuaXrkQyQ5XrSqI0cD1q9kxJ5kZBehkQsQbb2Yojt5iq87lscEkRVNdL4hueC
ikD+0OtazbuNaL0MB4gK57M0VASLK7kcBgACjWOcVRwqsUMAe4DhfMlpPrNKYYm/5xBWqEglHUYf
K4xgCfdLDbI+hj+GXk7lf7xAWMtroyPd4cneupkP6Xln4R9PYjhIRpDZeJRFe8T5E2eJI/U8td+b
J/OsXQmnmYnlZiuNZ6CALSnaRhsJgmHOUuNyHHFTVclXyyrjvPBDeNyhMbsD8JzAmpxtLMHLCDl1
f+n4iz9yCpIaYkpye/xUL16uVyjqQShBi3pVGCdG90pt8Q3lGXkxm9H2ur/DOIyrzj2kLSVdz6IJ
U65HibSVGpmbyIMOrWXmzGAjROH3MsNwF58U/13vByipAqCNTpqczLfvGuWwYKN7t1wMhDYgLSsX
EtN4J9q3eE/eAgY1MIcT82aNQ7nGmTffWxWAF0/tkMSsUY1+TMk7ct27h94kbQUFyo60zc46GIFC
pJ88ff/Wupy+C2vqlR+wpra+NHcOy85vXZoS8RXAghVRCYkqUJXKQTO9Y1Fo0L88wtlRQ05BU3Zh
zqK8omVZIhTw5jRpTkQi4M0JSoEDgRo8AK/oGdCB1NX6VQQ92K7oxXQd1aU3D4bgvgUNZODQdelP
opTkUe8VXv1YCMi0xX7bNF4wbhX9MB8KtpZ5H16Ql4LH39ij/N+bBIaU4UCDvnoRBeDXXN7OqKno
OvHs/wFThHlluEpOZH8TM6hAPtnn+uDeiylxRD7EUp3pepfLKgr4GDEnUQD92sFgc/XEppsLYXyf
TgNZiPxA6Pt9F2qdF+BTjt4vCSoYay7m
`protect end_protected

