

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DiIoz1dwiCymBJ2I1DU3O4UDdOCD1IYbLUI0voLUvMCBbKM/4INC61S/TdKSOoUevx63V7g+6/mZ
lHiHKW9CUA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o/flwcKffhg09UZzkz7gv/qZXGXaahpZlLeLvCPnGMHOV0tl8mkXW6lQBADTMwmBGUm7XZoObamg
kh0wsLz7sz0k84YCYY3YnDkU0s6XZ4yFdgj38M8k6+BTgeZETPuk8RfxBp2vQOv9zQhlLgklCWqU
H5aMJF7gqYDH9lzMxcc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3XDlc/RrM6J+fMEvhngyPf44nazd8NnlO+9fuAyN3g8+0X5quo1/68MLGc1czSBp+H9Wyu2aBKOJ
b7lFkbCJ13UBsZfTOKvBryDWOFa6KdkhYbTVSV9dfXRZ8PoouPNER1m+r+jF8e7EermzCIExWInF
5NIain6XV3z5eFAoF9+1wNHgh2DL91NQvcMqUhxodAC4EBuf80hcej88xks12032BecjB+B/gAMW
Fju2sqB0/mqHcdt7IfTqsGyFva1zLX5LMPhiF5YeiK1qj1zrDwFPgvhslJ9mmgozdcxNrfEp6yGo
skXdLgGuFnqjmzVIe1RLirf5OErXnL/7fcq65g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DYSqibotPAlt8I7+ZHxqG1W8t0MXnDrQyejnExd2/xGgdjHg+z1O251s8cO1MsyRynExFZebXN71
+rcOQqj1RiIoWzG/7+iJR/rcMh398jmqlJyWLU5IbIHCNoZyFsPrWxh/+WMiLYcvsaCPV1/bb8z+
2IY6rcDkaBrqk/EwYjE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
otEsDJz/b2bcmmVLOLfSwi5yawHEPe/YwdeYC6bj4QnDnh7iDtRlCB8Vxsd5V0BfHeL/WYjoeQM4
255fcpmsdbIm804UqNFTD5E3bD+pXsp5hjDUkd5BI6UEMxrdFYZ33Vo2q6da9Kuh+R1oMK735BRX
27ixqS9zhC9yoKM5h3EFDD4lGv1ah7oo8vFXQVvAoHLV46fz+yTbcdnzjY0CBY6ZcHBHkW/tXesi
gSqE+UJ05pdgmjP4NMP/1EbWm0c/tA0kZtZOMcSt52FHS77tvDYPPfsmt8s4x48hzc87BHtAtJLb
p2k4Bl3eRbmVYlntF4Wojcy6kk0ClpBDQDcHyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 32608)
`protect data_block
xeM38aAw1nA24Sd55RMrJk71lbzwnTUCqs5L8LBRw+sgxE0OHzo3oDx/3JHEex0xgNT9tOmeOypZ
siwpT4TzTpDtcNbhCa3O930pFrFLTrPVRYbjqi9c03SyGjdW8uO8oJEzhWpAo0eZZXwgsoEzXdc4
vt9d8y/yJ+KdBOWZ/ksxs1hgJV7Kz3tqJUTeXltUDKWeCUZkiG8d4gkueG8bzRHcP3K/u+0ruzNM
9UwAhfrbJRI5haJxgRJAsCSnrPGvPI48xS7seUKOn4TzZpteBKE/QOGTymA7sQ+epPDcVL809Fk/
n2tmcs0zlPhktx8AjQlVTjakgK9N1aIQC6gBADmma+FvF8gvQvhksL9vtGeKZOKKft2VRGXzXr9G
uUWRB3A8duvKHDTe50VfhtCe8n+TwmZFoX7xPUQfme7vBNcYjK/i4djG9TObxJgAfFs3Im59wXYR
MouDcCjoTBRlXppyuKhVu/3Z17aAJ8n+0wMu5DOEPNx7oX1590PiEgbF9y1UHL/8uIBqEu/9AJUq
33iNO5lIeNfWmxd4M4rCGMbQb1K6eLixPWcYAGTRGrT9mBK3AA5PJx89JfgJ+AtXYLq5Wnp8A93l
1tMaepAPY6wSceai5ipVxymW9ldWb5aDfcwvKe1FNISLSAnhzahDi/x0UlA/ysxe7Iq3Q2uPeHfP
4sht4odjbTTzTRS1+GmoS+sq+QGBTierRWO4Crv2XHw1KykR1rhqbNePorLLAZfpv7/sKuzliVok
CXc27j/NSVMHWnkdwYMFRPlOxchJJnyYwi1zNaenOVfMD0QPJt8AtBrX80QI+sGkjWRH79t0FLtU
NoVbBu8Va+md8Gb0ynVBZq+h+4iLzOIFlkfmUj/QnPDY6kERI9VbDHlGhIMG07Y49jzCsSp4eBUR
n7CZeEA+1s1Grjlth6zzEAbZAWo7nBY3NmAXwRATZO0I3pko2PfPU6NayPu2lSLZrX6Gjz2DnmdB
1ySn1pp4Dr7gjX7oLNO7qnINaZ14hQOoMxcPZ2VRqnZGzMlw/3yT41MQ2lTbvsHNHEkwdzN7knXV
o9D2cMHWUEw8TrhwSryYRTsZ1GScrCTRgiMRyNqKzs9YsUVE8W+7DXYLrFibDFC73VSX1L8FEFn9
y5dQFYSJ3BAYdwEimaHRUrNUTzSj1JADak7zu9XelXFOVXMKis2zJy7kBFYvmTHtbiud9gXiWEd4
w2FsLFK5QcGhbvdv+GXNc2esYcMkhJ2mSrNinCdq20mNFef/z72yQuZKs+Nuj7SCFwZMdJMRyJC9
4PKNgN6u9f0VCUCdUQN061pIQJtD4AGb1xhCLBwAU+QyJ/FEShq/nJegvq3ba/AD4tX0a4nuyWbg
bTXVI/ya9W4TWilDlWYWojYnAKoo8tpHd+SllS4XgUziojWDJ455aVv5KLhkI4sS6q8OBAxPfzWl
iBYwz7nDyOqo2guS7ByySywlbbIx8l/AVgSTO5amOL9HbthayfujgVpUXDswRx4Pn0PyDY9zXOGG
K4rnsROzMGff4utXrDP7Xvtsq0bPfa38o/qa+XZwIOKdMxM1TgEOphE9vakWBQItgxyPPXVLcV4v
IlqrJdBjS56O62776SOKxhk5IBwvcUr4/BBZGYZC2JL13lqbFD6oMgE7lB+AzUC+5KcoQjvOVkmR
eudHDyFBeencCFhZEgxuyRc7NtuFTUO2o1HBIX63L8a72P3t+axUL/5jBO0+glM9V5GkeV+wphYK
ohj5yf4Et6yaSz6Ef7EVi4fLbYzxb9U6G9v8dX7hhG2gNcam7GD0BfbkIFkaeVMNq63hQ27Z8+Ep
r1Je7BkshPGKUTQ6xLHFcc2awcR5T1V2oKsD09sEEewrNt3qVLVl13041VD8P3w9KGbvoj8zYPzi
QrlDlahDUdVfiB5GW2n5SjADYKrz403W5yHY6u/LZziY+m9Zn6wUyPhP+xfyoeIEh4+EEtgefUeZ
JqDBFLVzcGbam1fB24cd9IqBjrHexO2K4iKN04jk/aZz6gIToLTbmBNC0HhwFDR+pVbB+BnSQK0F
nYiMv1tUSh9JzcnfmzNVXXEbx9cMC9QBjfs0sQxzaW+n2WiovovhaMDV4ZB6Vwvg1ysxDoW0Y9p7
+pIyNdjXcjf6qMKXq3QJsvsWGrWoiV1kHfxNkAkJxSgkGiAiyEdP2jCsPzj4CDip5Ceplw2Wa+Ia
CC08l3UpsilrnvDFXC9qLm/Qixz67QexhEEicfS4pzutbpPgnVu7fK9HRY4a+Z2mCcNRysc1pR8y
4foxTg/DddZ1VlhtkGwqhoRjpYeSd288i+naNhFPZBmD/VUFWPygUwTgP5DWd2ct4lSTZ+ZUsu5+
gWLdVPUBe6Xp55nGqS80ekqwu+eHKkP2xNQxrC3vJpFIBoTMGeMnp+eHFHbxAF6pxYWWvbkGGZyt
gHd/1NSK3LPMFcbX5/pzdAxsM0++jPkpSj1e4Wf13pqwx62tpv6X3AN+W/N6xHCUrcLajjRNB6GV
kRueDU7AQv9Zqe6KzE/GqhEC+5gkwpBMmy0uZYhKW6d5yUY8JFe00Gn76jbChQchICSWnupiC5Ai
cVuMEB0xG7ohFdszu15Fbv4/q2N19uy7wP4Qbib27COkZIeYT1amjMWOadWsvnNO5d4qd49TRS4y
zoSGNTgyWm/6kaSUFh8+YD6g5zKzCT4q6MG4NNEHD3gVZd1mDZRQHXOifhFJoeEmblfiJtjVDj8f
MNIrHwHEEIe2Av9Vv2HO5pDmzwW4QKZc5YTvXPt0TGhicZv50kzmtnQghqTg5KvWalQLYfPR/Fr/
EZ7PD43wf+zOGSivC/qoUyMStzeAZTSKZZH80P1+22CChn0L9U0rvNcUceBaJxchiBwb4tQMQvvS
xdH5RvUI7Jf3HV9Mvrmz1jxnwyRqe1qo+VYQzAg5fY/tJZ/VaX9vHVXQJ1TFmyY7YpeNrHGgs1RJ
vfDjF6TaddE60CH4uk8T9vucz3B1Sa1gwKR1kveLYGSI0FASezn6R1WCz68WH4s1lOWZbtwO7rID
Ii5ogQtgfOibQ2mZsPypsj+DAL5m8NG5sKoBQoL2DA7rHPD202qXnKNpi0uU09aOZ95XvCl2ybe1
Z7x5nl7QgWm0R4bBlzOe6AY4hun96+lylcOfXy4NAVD6XSFwz2dMHOjZ7ghNnENLasTqf2ultJZK
IaM8PdEujeyBfXYql0ldq6Y2CIWapmlDP4ChN5gbwcSagJ4JkY9IyZxpIJ4TChIRqjZhqSE/iFHY
XaYxnQrxOYaS9EIbJl0NgDCT+hhUX0boQ1ht2KPrlK5+7rynCr7+8IkshppTI9ZQMYtqEcjD1wVj
STQXtuj73GJ03BqnXX74jNZkupzK4aI9UW8hp3KMx23krCX+Rfx5nc5XYgqztznF5E/MFQ0AGxuq
I9WpG1OVr67w0OlqiirIAuRc1fH/XBjc1RsbDDrJfeIRxZqrP5CwEiQtbxrj7pghQGoXVTyH/e47
gKqdDy4roNvuSJxI9C0GEcvK9hDa3KrqDS1YmsIivnIfP+BWJrMIkbLKo5C60mcBpC3u0wbfN4Xx
AZZHdUFoB48WQyAjtW++F02mIBcZGnm+AtbQkVTSCb/f348jwqaxi5Z5VtlvTnQKPlMkz6m41Ha+
k5G4tmAIaYGRId7QH9ecAE5+h8ePFdlUX4NQ54gXQqCZBJaZwFWcMe9MCEdSOP2S8/qJztGX0jnJ
mIurZX6XF5fgl3XzOUCfZO6ot053rCf0HM5e9Xvuii8t0+xbAUacsq9rdTD1AL31zyrSm9wUDiQ6
1HuUm+XIVsvHTYCttrcbnAk5lCext7nyGMVIfvnvnwXLpcv/i5QH1BaoU0nb5M4C3x8uF+JwRl28
ZemTzDxUH0m/9fOw2BMKCpd84W9pvX/gsRnG1YE9Cts7TVLjFi4HRFe/r4VEP9pwabUFVrl9AILM
xnjdvddfOglQKmMHD2iMtXrTuTsZPDz/7HIPF/C1oy+Hg7hgNzJDrSl/1BVVy4tQVs0fZqdgfrOQ
VFjdBhpM3Pq9GwRy7kY4UGIpjCd6wY1le5ysuO1daKNBf+BYB0Wtq8vpdDaeZNv7Br5b/NUY6K3B
ccuNxww3P2QQgPjwQie7xBAmIJcgm+fEu0tTJKBw/ajmeDuQMH933wrGMnMNUxGmwsgY0C1SquLZ
RqGKvd0uP/AHKzAq7deebYqSnkYO3EiyMryADNQDfq/d1PBGWueETzZLj7a6UvxpRvf5/RVHGOoy
CWNCV6LEcEnpWn8h26WTvW4C/tHkMUkMezCTUOZRga+eWXxJ+EOhvAzQkDkIksRPztfvYQ8Gmj9M
bJ1kQEP/0F1JJsj2gvFVt+64CV7WiJ4KRWMayceP2wGa0kwa35gtut1SniULDuCvi3jYl0mlQT81
7/hg6inEwrJU14vkItiSgHZvk9IF8qJlnedT9AYp2Qeqe4UMckJNtKpu1nQHFwJHZiQ0dRu3BI4G
0NS+fjdl6O9BxO066FAx10SkrbqroscI5605lcLpc7WH6hZU72UwmDYcxYuzrD4848xk6wZJD6H6
Qlm9ks5lrHsm0nVMjRtzsoKW+ALuNMlOSR3RFVxOV5LYcgQEl/0upCplXxbbawszVHhy5Mxi6+ev
j+0wuM8GnfeFSUOYFdv5wlUeuQgVCIXFFz8xo0ouTQZFeK3gobuBy68pjAhzooiBgTI1d/WOTfqY
U9enY/nDBwsYKtiJFG/VoUGyTD42lv3IzyMq5MH1mQKAoJSF4cT+TLohtqjCuEJ88ZwUe/j/YTCZ
CZ65g+jjjOFLlc+ruCfXgv7zjKbi0JZd5f1CZZCLqr6LPgAd+GGTJ74c/4Yxc2M1TiiaqYzJtzpU
T5iJuAMpYlmp8N4BHkmlMLYE+BSSi9/9kgrRXi4W/WK1B+F39v592zlC1CRzKd/n4F0FBTZ4Mb28
cC8Jyyy47h5BEEC8Q23o8VIUwGsidGhlY5a009eX5zp2nOTTGNjVO9guMZNIExPZEEjeFWAoQUUm
ajXwBFtOuwRiLgEVQDtQ1SVKCAr43gcc/WfMji2VLAQkbF7TOmeldDu0wUGSxVP+YiFumYi9mnGG
bOVI4nopDOE4/Mzgr2K/VzSyMEEvIQ7QjDZR3QMzA8CthU+/+h+4koV6PlQdHhl5af4THyApxyX/
JxYQN+csWLrxggeMhkHFoyJOghGDWLo7hLvtejtTRhukKieWqOTN+X0paXfG6zMK2ryfB+h1ly7N
QrqtNr7HVtVX6jX9MwnJCWomd5t/V8s05SJLdz5NRYNOZ8vDGRURFsGRlx4WNIIWJuq8246KEHCS
/dTlTy72XVkTkw4RvCl/ycFkE7MqbGSJsc05isha4ONcBnAD3HUl4DydtvQOF5yp6j2dyhpkneOZ
5/b36tVhEH99qu+7+0dXHoFA51l8WAfF/nI/k4XJ6yEMrvUGoguUJZVmMVho/RsaIeymsxH47vKa
aGjf/nn1SiNdda3M+SvgW4sj0fNGrBqPIPtsZ2hhKgI73oKpuEHnPJtwmlUSUXo/TMWg4BYusYEx
oGtJanBKFH3MI1luqCP8P3z+6jtIMQcGllo2jeWzWE9I3yC74j9geZBs4pr/HwCocfoM+1nxuufA
CA1xP1onpXviZbbEIxnWIHzUNAvyMpq3QLH0T+u4AztBxuG6RFsfZcXcuGoUNpRmL8+9GiO+tGKu
g48C6zgmHYYBNVm0QAp9nfJJXob2c09+1oqL6z//S8yIemnQgjrH3eY5z8NinCRiGZdrSt/5G3/c
ZJTl2UQIyD+pbSJgMlnCWLs7zUD74iNm11UVs0LQegKEs1z1pDn9llh+CN8fyWFe/m5VlWle0WdV
PMC0WcKYSpOBDT5FtkeGNcEYo+hC7wBCpzTyUIV+/NfLt5MkqVTgqHQJB4d0DzlDTme/xbcrvrCe
prYQ+hlJdkSseonnObl8kXtyqSEvzgpJ22bUVadeHaVdV8bibZtsipNrDPyrkUgVk+gY2nxTURFl
lQIxZfuoT+z28j24IGPRdo/TrkZQ8zsEjGUKPtjYDjLyx9b4UHTW448G5eXvaINhJuLn1hdnZUFY
UacQ98w10LHu6MFC1dwKG4QktRh5JGC4gy+xN7t95iQY+YbUlwzepaXH9SgjVQzHpKpGHJ2XUPwj
T9i5IWYeHGFAheKSUKOKXoOwscQq2S2oVXIh1matz0z9vLgXd57wAFPIy/HMo8WPGUgJhtFl3uX4
muyLIMYqLPgdtB809SqvAKPH5kNZVlF5sWVff2XmHUT7HtDDUi+qpzrLZVxuyh8Vd3y0MWo5pABC
BkcgmdM4YHKGpFOgll3KKaH0M4qb7rXiEhoSCHQW+93rMNqRiZHXIVk6z6MeN5JKMRRGV2lo8GFX
X+3Ng48JzNlqj4VPn37tcxHwRbqoYLrtgNwROpzbtt2FyXMbISrKAh4y5HOCjNY90OR+HEPtI400
cezAdaHCiMjbPHDkmGn1SVlCJvM8KZUM/SJhlDlObmK5gjR061dw2lnF52ATyBy36XjEAn4YAOPK
RRJ3uNjqO9M6f5T5YKWq7r9S7CCl00jpDROzC0DriFkb1PGn3DQxiP8d8i5cKPrOgcF7gJ1uVpOg
dge0MoSrA14B6vkJT6WJugwN4ADnqTOs3hcwp2hIJxbQxqB79tjLMsEaqYT9lQ/gZEhwJkKb8u6e
RYf39DfvOG3R93nNMggjPyTVnwur83XB2nHBITRm/5Ijhi3cMtUktKM0CCEZ/VTEdx7aZswI0SH7
gCGXy7YxzurcAo3QPd9dlqtFnyX406LDT9PJsJTuMV2lT29lOOfJnGC5JCM0Hr7ftjEqQGx8LDBF
du6SinkYxigGu45o/vh6dY7rhCD3uJiPCbOT7CSfgcwD2v7m/XthEZz/iRu7b0ldn3oMtQKSdpGk
vFITiUlRn4uGkkFzaqdQcWl/F5TP/zMZl4S9oeHXT5O0GJXIt+y1h9+C5kBIuM2Kx4Dg8OstYH/H
OqHeqatWyq+E3jqtPZe5qygXfHlCX9/kuxAIBArO/8aSxG3gYFmhuFGi4re1DnhMdPeHsbVcUnFl
tZdjYgsX7I28QlbB/yQUWEmj6x8v4jLIXI4f9+sTz1RZz1HBgVXe4dnMWmtgD1dgSZxdk4Br4mXX
2cP63HspU07jozjCs81viJ+8pzuoXQ8fs6ZiA+HORY6BMghPvsnpC/nXyqVq/nvG+FJhrwioPIss
t87e/M8Ud4IUKIi1xKfipzloGatfOveDURNemq/zrGsKf90fPHRSs2O7sTZf06J8hhxFAmgyXGko
p8tUlozOW3paNnCeqcmpDWzT1A1RFB6IYRPKsWdI+dS/pjoU0PutjqpkbeVAjHKoMyf1rlM1grsd
wMHG4zVIBvTtlaWQTPg1SX7rR3JRAvEJcXytl6bgVx45BUElvWz2xltdQmChUKhP2N3dd1Yodx4Z
3bZwFKhWwqH+8sn5A5tCA1ICZStPGBDGy/R30j3H9j+5cMl6OqOp9N0yIUTft0dhEeZzWzQvs4/x
5UqavnvfMN46BaNeHMKhmnJzSxGSJ5GDnSER/TG490J8UdC9Dha9FCc0gjAvJgCGHiJK1viXWQsk
uGysHhYvn2hAKiLxWICXaHT8G9m4kJg/WlnjIEDPQV+wEJGt8+p2RGA9xuVvWR+ZOcEnt7gdeVr3
Pi5h4UuNXkqfOaW/iXY3MZDFSHkU0nYWBk6oYNlUD64BLIA+eX4OTCig9Ss4bxrI4JFbVVqjeS/5
rVTdwZGjOYBlEwy3g2qI+WQaGdQEO1Yx+DNoD5pbsRl7f5ALsGBpaW/a8LNeT+boAvVeImp+uAlX
MBMN+RAlXks49ufrxqLB5rBwS3ZzEyUNQrubujTTGXSLDzYzLXEvp6sKynloDhmJYKlwMn7qy5Nj
Rm1ZMNIeFw7Ck2uaogMkbcp9zY3ienZGF3joBbp/d4F7WRFiuTOdHq1tbzRuyTTSnBJc6/qiApg0
H/D10Nb/Og1PuBe4KaIBeZgcjHx9/Te9WJZ4qDL71GSTOGgX08zonhoa3Zpw1wU0AYyJ2hJB0BoF
Wzn9bA1K21HJgkGFASE+xWGtzMtU4oUykRv76PBijZtWUZQHGsCU0eqpBRGQFagpHGo3cmi1peAW
fwdwpygLWb9Xe3YaHfkWX0L3CCC4LW40wwx9TJ4+yP6jY/QcoVUO1d55GgsGl8pB+mx0WfcaVb1m
0vagtB3Fz2ua4205B40BVWDpZYh/eDn3Mx5wS3lrddltOgQB0RwC1Ks+skKeulhBEiOEs6lFALM7
qhJMjjZZUygbOn1VUpY74OkUbx8UPx7MA7RScip3uSuE1a9YozmIvpLsSn0lAVZ1BPKBh+KgwR6J
3d5wEdX3Lf6+aq3x10Vt6jcAFgiCGAVGlOMUnHI3WmaXXfFJOV1Y3IJotLEJweu5yXUto1F9YIhd
K78BepSlnZHhAOmuH7cFzrnb6BQShpr5c9zVpUMdfyWuaSSrj8EWMkuyc204W5fcuxCGCWlGnu8v
/x5E0ekPdbulQHxzGIHmTSlU2+MeLaH6L3OVfxH5/WqbCPdpwvC+xd8oOCT4O4oT8u4RBP91IX0u
GgY7ckFxuIcIIea7mBbRBoijIh+m6w6/LXh8sjiekQi7O21ZJksE+rXXDhHGv43PDS3LqhI9c9ow
tEjJmLBB+F9MG//IPH7j67R6BqTPknFdumDpfsborYuIvpew1ciz7JREDP+ijlpw8zJ/+MvpzCIy
owBeiNF01HbtUap4d7o4bdmwm0AJxHNnz7u389E2bHDvItVS6NKTjf37PlNK0QKDFSMrW13gf3Ym
dCq8opFX21q9sPE9SzbyPmNXbSOEahkavep62feI3FWduwXX2OYvKcLSnsZzLME5kBVfHIrB7aPm
SjYW2nQnYU88avNGGVacbxymRyuHaAWrF6K8bjonl3o42VfY2IU5Upm+aaxVM2Vs7Ycw3NPaFfWb
ntXjgmB77UbScOUWlqEZAjac4vB4wzVzz3ydbwEvPBCL+ezRuE+4sa6VOuf2VdgLGUGI/Enomn7k
9Zj7D4I2cvzDUlv7rDv2rLsy4ZKPMZL7xhOElHcluye8QJiCBDS2NoaHasx1P0IjFPoNzvmCSkYg
1vSgf+XfMvF7ekyqxUEg31EYqD6aYgOzL6GE2GU5d2/xfCltYR/Re2CbdlaOXZKvb0EGWvO2JD9y
ikCx+KiU7RFqa71ZjXxlXGwUFrbypdqAJNj5kd5PVYKejJOzjnhqQlIO9rAvWKNu5pu4fLSqZ2Qt
9rgG+iWlnDQ97VNVZbAbl1lVDg3YUtCwaYusCgQfGTHcr1GXp+Ryjoz0HK0R0t/FsHux2Ft3GJvM
RlKyVSYjN3xPAMr4SIoY7yCLOvsxGo1nMNPZQo29wtn1J7tB1c7Tj0sNzkgbjmktWV4iqMnex0a8
1ocfg24+tAb5bFVQCbfk9OlkG6l554MhAiTteqKCzVrW1PtRduKZLtQyHHIPT1RfUQhm3pPsKQDc
dca5vcSc0ScdrDrVU6/zxtRq5i8R2dp2mQom9qaRAZl5/PuSIwUFFHTibj0YSEwDWXn+T8yjYykT
tJdj+sO28QSPDV6Z7rCDyZqcHr0m5o4vKrz+R7Zx8Yw2RJkegg+/YMuIwiXoYL1blxmkCk2dRsX1
U2+16OYBnAnLbkf/5+TqvLnjrTlAMjmhdnBvIu7tsuBHVqZo3kWTwJEqAWPkqWhDnD/cM3K04U8w
wDrsdXygqARtHtpK9MCYYfvp5KTcqazXJSv7FX+3bgxhL0GP+Hv87XCzUQzxXG118Y4HawKk52ff
dRHaICjh2gTtJlFZslGfnZcDKk2hORMgo6JLaK+80flMpky1BoIXThiaETh8ZqPNJA4cv/BP5u4G
VkMuRqJ0pKJx4twdH8bLGJuhOkwRjCLunVRkksqTrRKrrAOtzegpNvJjQk5C+5WWd4d8zouneR4x
5P2VwSm/mJkMb5AhytjJ3UHtpzVFbrBvVZRjdbX256qrO3T7tYb8QfTSY3MjuIbyCsRSmt0NH3MZ
Dy3DyuSnw3I2p/lIHeM9htRdEfFO9KCsXz78z3wGoJ5r0NWPI7QaTQE97Zexd7ApItjvmSvNW8Od
IlMxmfmcxEwikb3cDJrAFn9IxbpE5DoH4FPqx6BAmp8C0aisukIxUV8B5vTASAhQyKzG1TY5fTD8
CtJi+itL/srDJkmOcfipTsjGIXBr6ANKjod8xqIrx0N5JnmXJY/YtrCCMGUhW5TqEegbxZ5k2HW5
ombL7Aa41tmF052f73zvJpL5XfdItmxiw0R9U+0K9CH9NhX80O8hstktBg2+sDY2Cbwf6SXGeJLC
8xuIh0Q4/IyvZ7pJVUfPLOjopNuU3sDZz0HDgP6PHf9ojVtNCW5LWKze91TDjb3O2kQcdcaH9Sb/
HViXI/rCk2h+9CrS1rDy6dTVrZpC2vIszJ78eLwWy95pCaT7NNZAaNP1BbB2hz00axO1dxi2/qB3
6ulsYwFzezzCJGj0w0fp+WSRSWiKFlUAKYmbRHVPnP8+9lBLqRNliit4fpqKHRJWKS16cYCISp74
3O/PzYC1UsDQuD8/udUzvQkT7W1+ddW9xFeaCvF/9++vMd1PWGbF0WD6wuBISoBv74L3ZOMG6GcE
+rO6vIcNG6v6WO9RSFjpnLL8QpsREFJl7b19A5q5xUQMpG+hqZqAIcQtUeTb8igf98qtGKZGJ3LT
7vse7QJw3sks96atf0w4sjGNOns2wiwRMPfiW1/+nCEJOwa59Rud1da8LeBC3VnEwjnMPRkE5e3F
5wkUHSvhRLP+1o2x25fdKOzPB5NZy908+YgO78NpG/kMYzz6Wr/gKavfra2uZg+ZExvjkIiTuuoY
d4YeoKG2CLeotDSKebaDrZrwCf4UM2m7oJvR8YtMs39lVlsAwO1OTn8WCgLi9zTgn00o3vLKPdpG
sqq1rorgd023R2KqWbiRGdQ3gkZHIx1RDingpfxPHM0VhWWy4rFBzt7wpwkyUIgsxFI7+hhBeNNx
gsRtzzjkBfN5LE+wII/ClCleYJwYDIkHTn7/ZsDHGMiCnpkCQcsjMb6zkOIbfyN+nALTTDATEZya
xJRDwKFaIn5DsTRHRAh7PPAIUQmVX3Vhpp9IlIRXQOndFTP0rqeBTg82WJRINje7oXzm1hP9SCUB
JQ+MOO4szwyyfU53KRKpeR0xJ2RWK/CECkqCJibrhjdHkr7UiEjqbJCzJwY6TPWP/v1l1RbIGKzK
zSpc5L/V03rFVQN/iPKUigzsWPqlSFb4yY8F6qmuzgLb4s2NDVMuIVA9+y00BYd7vVxRbhGCa+N8
Ai2NRqrND2mYOoq0PW6XEs3UrpoaOt9zptcetPZgNoAjb4uMGtSznMlsO4WNhJ30vE2WYpGyq8wm
w1Q4xrJXBZv3sdj6hYJCWX/AVioGQCNZ7+YaCkj89yBdKHFOsCukJQnggyQnzQLeVlEKfLOgPOjk
VSHeR1k6lnGQfK0cDGEjYGGapAC9A2qg34luwjLYErq/FWq/OYXfG/uW9Y171GeIp3tGP0WjNLEZ
GMIt/g9HrfFfudSF53NptDIDlf9lPk+nrmFQpUH2WHff3TCEIDZqW5/KkdRLa7SC/71+VqU1Fsk+
qQ0CmWA8NUVQOHUPXho81esiA70Sb3Wyt3KN/Bruznld9R4nVcg4+y7aaoTGAc+pLO/CnugqhuHs
37E2GV66x/SqxXlPI5tOA82uFZRUwHEEJ2K5Ux0S6d2E3rU4UbA940kIZ0580lwSBBe4R83tDoLf
SPURwP59JjdlMtzy0QwxnoYFmGxH/jnK54yHGj6sNZrefV/wckT0nD5H9OupYLsCqPxTbO/8qkOz
ldsqSqbSeIDLPHMDP0voVdYAs4MecGMkdgKKZVyJU8f6JTZaimBFysXoPJ7zpzHvByiKIfqf5TPh
kiNxp6VgVJnhGbojkNdXA8fCKZT5BKagkGF0Uw7uQf9/sCbLqKJUNvHKkUssWqKMOKnxFezkrXtI
BPFE4xY90smLPC34boIQr2rXN3Al9FdOlJorJ0HdbziGDpbUn9wBhK93H/Tdm+0Ir2g/qCIHujcd
9iZqxU0M5oxYjoexqLmAT1SFbkRzNIHDUSaVFb0EeKh+SUltMc9ncb5jhsoHsG0c6CL0uBu8ozBD
t7GQRxJsd84q4egshaz0Sh0ayUyUz7UiM8TKSAhnxnVex/QJ1B0UzuMeDB+rvlnBGwehUQywanB2
pTNhzpoJvLJfsQgpC9fqGHzQqirgD+tHBMtVqfRr6vWIdvnVK9LoRHLGTbWlmOhaiQWhnD03xdvA
e7PL/pjB3/XPGIeG5ueC6a+yinUReJGxLVwXRLm+ptzbNdL61VkA2QMo+0iascxWJviZaRcVV7mu
2TBpXEiabSrQ38Il2V6lXn2nvyRdI1+r6QYZI3xxYL4xBYtWUW5L5oxPBl8doDX5Oyv4tRuiIPkm
PCF2pHj9ScgPHUJTWLbWlE2HV9o2t6QuUznbpouwqgW6a0y0zIiiSH2TLag++J2j6rcJbUlwDb74
8kfRHeKYuqrmarRaDYtc/PxD+xDdm1HVNz0YKkylcP+jsE8uNv02yKbo0V0MPLzEncHdtSR41Ck1
APB0x6tmjcrSCUZV0UyazvNCr8JnzZLp+Xszb3xd0PluW7F920//FJqPLWY5VGF8I49mntpLBvmm
m6tJbS35g5lxYT8lpm6s+f/SLaGbA+R6bwaVBHav6n6ZNEUzKGxBDRr6WBzj8gy6FrtFee87Et5f
mCy00w07kuICLELGMMbOI7ENfJp9VM8xQcxQH/7ZkIgeub3oPl/Ms/teoW/LyuoEj5uf6IVGBI3o
prJwGbHgExP5XvgHQsvO6Cv+vWhk6Its5QF28GuP3mUSDjvuz8PMzyBdBvTRK2Ck1QvjowaxtDC/
dYTDtKftgdc2OVGZXHN0mSuS2k9uUFUMWwIHb+OLn3hbH9jckk2ivfoWS7FA7lx2GtsidrWwkKfH
OZaqGXE6JbgZDbm8WQC8JwuA66U9nUyfPERf6U0tdClJMEhYpxdxC0dLpGVB0E83LiTvve4XK5AP
bnKo8WbSq1cJ+K4SG/oZZYHphSeKF5jzrHdjRW3gHo7+JtyreT5dkOhRao5YzqHVykxdKkEY7U5T
nQ+PXtYBQ+k8vfENsgS04/hIyhGOq7tIK/Scw4uFoWtQGzNBxQSRh4s9NTp5YeCWKEPvSVdfNXO7
CT9QWmsf9DwqShYy8V4Gc9v4TjT3G+c/cNCB1/q5QAKTWg8h8oaXZATIb3zh+hfsPRY3zjIGTDwW
ZcJ42Va99+93mQK2MuFisFTOJVdgmMh50wKbJDn/yIMVA/yawQrNwQj5ZL0jiO3I8wCANQl/5+lR
EC+vv9Y8AU5AXg9vaZRKpDiYxxlqbMzz1I4alQ2Ve31fdjLbigkCzmZgHd1Rf0kaaZFGM7v6A0ru
8M9DhOTsTQLmOzFrRRYP+oCnYAffv4rZJWO0/dZjsoOkwZO5a3Qm1wtM22ezrHHaNSKhu0kXkkc7
DC7pT/YOvb2Zcwk2jviWyzSVRcge8PWqs1S7Er7Z2OF//zG9KLdOICvWKNVRUFDpLRfm44g/asiC
vHbXLI/XD3fEwvaNl58hcmqqfJ0qWw1DNZpvUYOrF+MHMnz9oTZhKsVZoDrA7Ueb9diP25IBmzkR
wPTnmFWJH0+LPwDJ7XFrX3T+qQlrFzonirvhZ7aH08kPhXG3mtbV86ePHAxQThVqaZcd1iAIpGFv
VndsvPid3ii5Gta1iOdY65h8ECkvL4IRqk7t+os3suTtDDrZF+Z45crnFzNrFriWsr41RZaSUbOo
Wxv9xD8DQ+6AKImvRo7v6hsVNWn3a3NxGl6OWxyanr6Fl7d9Kzx/ej87SGdGyt6ZVHaLjmhTaTDZ
e2LD12eGxwqHYy/3mvR7DfVvsZ3mZiCN7x1gYB5oItC6s3ec5IPa8ji7QDYcyC2bYWVb4zqtRO55
hy68RD7wSqGaaWmmCAqTaXFmAdYuZCXFRmM1ueqQvcJOOtVyKnlB4eS0uYLhn0seYhhRXxHIoBio
ROT4lBUWkfyiZ4SCNsF8wyMNt1y3Buj0bdd+k+Z0AbR8bFcBB76WUF7iR56STGpyzQ7i87jDfnKZ
F0Xs4OiwYv7FFWX6VIJFQz/53CHDUMTbgzOfhV9+WmGeHLr//hdnBnn6iqDsj3KMdPy1ewEC8San
jQvaPcpwSVpnM1UQ5qWY8q6uFZ+6n/HRj3ZPVcxewwi3Yt54O21YGe+h58vCoJAr0Ct2q4MnLbR7
Aj1efmYyyqJrvQVel7OkAi/2XS8TRQ8YE1TyP3ufgGdYyczjIA34CVyjs7bHVeB5fZir2r5jxHwH
g++m6MzSbGd0a9DDRs5MFU5IAWh60V8srNou2KZmkdU9MwtakoBYoc1hKMw6uIzcapr5fVw+vt/M
DHjmEHWz7ltU5m4V4nnnW50xAT1PDYrHsnWOD/TjjPyFqsBZrFzfNQJ9yRVTHgkeAgnyVD8ii/Qk
mJgg45L30qZElCHPztd9lo20+2tZ4dNt8HEq5kIMpNZ2lEhocPA21AbqyGU8TxoXv8CbeQEoqgpN
G0QSsqIURqrxi7AAioOMHde7Rkw2KIcYJJY4ZWHd86k1Mls93SRrPOx7xiTSSrk4YhPJQrwfOTe7
QER1iszbX28t9K1x6Ctiu3OsPkzAvpAmgQ2TpY4g54whqHOj/vp7mujmknh12cBjoSe2/Dvcd3ma
c0SGOzWl1dwBj5zVVPNIRzqqcdi7TYthPl+DoaaxOLzyZaXx8iIzfjLrNY+ll3mfswuKJ2PcEwic
MwOnKrmjZkYE+UKmd2OwxKOtQB0I1NkZijYN+mwnOT5KaeBGZdmLtvgPs4b36L+87Wv/LXY1zZo5
459/+zEQR5MrJheiZPJIWjYf+k35fn+r07vwbTJxalizy7B/00D7EbzZGNzPC5dgYAob8stWX/ee
exsdgovPHVCgLcXqH6mYkZo96s4d10PMsBFTSYTaa3B4ZWUBdIh0a8yIv9RhnoYj1QmaU5PB5VFn
Hi/KYR48c+bVNipucCDTLiJGUgOyAyEZA8faJLmXrQC/MTQh6rceEb38m1II8Std9OVm5pqyHF/d
kAFkl8n6DMsZiPbhdmPJK4PdLhwn1U+xshqf3QGheGf147A/vyHaj0RIJAo51Em2sz50oWALk0ti
Ymv6mQOn1w6EcBiw6OoEq5nhCb7rluWojXrui56ioYMEziJr9ipuTGEso2M6l2yDGcG7tALBCm29
o+HKKwKXW4LF6v1MFN+R9axz6woQ32L9kY7KQK/i225IZNc9mnhzbXJJC0FS2zNc7JYJ1whdv5ai
2LvY7oEVwl0Ou2Rc7HXamdyFUVpNge9g5LtTUs/fF/cDtwZ77ywZCi4Z1RHG20n1GMdXO6mtG3MY
cDZ2i4VcNtKtx3yIlp8YMGJwndPliIyabOkieHWD6ieGD44ggAAqo/YmIlqgJlvUgejGQXMSq430
srxYaLgRulDTsy2dmenVKolpbP60tRD4JEIfCPajtsSu4zz5HQbbmqkDJI/tuMgJL7WpHicLF0Ly
JQSSHy9zvtx+rAfmg2dcfkZ9PPYEBBo88xV22PwwdZRqfNC5L/r2PWP0tSorIpuohsdbD9rw33T/
ets6aHghCSbC53Ngetx4Wwlcyklz1aej0+bR4Xd2eueDzI6KsoEuaTbF4QarQJE+DnAom5szzLQ7
rgsj+Rhl+OTzIPrDAOtxh+r8YKS9mIt8gt3P/RJqLu+oyi91/ilhgvGLvew4wvirg+vdGvEFhxhU
f0VyYYwEhaLR+yefeoWs46AeCZbZ7Au/d2WLdqDXf9zulik9MRhZSZUrupyx7puinbHIH5k+s4Vr
eqVDXfghLPQ2UZGtIywHBvKYvF/XV4ri/i9yjohxyc1ot0szAPyVeXZ79lLYAVjhpPnYMO3CKTcR
N0R2s89hMOPIdS6zwZM/48NDyTqJdSm/I7RUGQrhH+yE8od4xWUo7LeQNz8Ln3rOpUMMh9Yflpf3
WFf3XGCvbZG0eX3ul6Rkt3a4dZN8eOaTjN9TUml2xCt9e7t7Nm4Kl9Mk8DTh+gIy0Mf20b7NKnjG
mmdxYROCR2bJc9gPjreRE/kND+fgKmJqYp8A8Pdgx7r3Y3KdIfiKpMVJ2Nvg1tH6YvZds4xnxQaS
x+430GhdaWA7qHMDZX1dfybdNFFtNL6NNropJwcPOkiaVf3TYAPcwAdy13SA3wEP/QxjGYmNoc+D
rOUroH+bzwbegXSrgr8EQBQXwQZYGnbsvD+r3hJeYEFfapnDftwegeQAzCOEUlRyZ2PH6IkLvkxh
Kf0LSD32qqOZkS0+DcRJaWpeHNrG8+ZAlHoSwx28CN7ova8NcNHKlBwUCCl2fHQoP+ZzwozD5Odd
ekuDxTyqj0TZPq9us2MPnXY/ldnJrjIL1dxiylXRVsKfXVxmKQ78L9TwIgjcSrl5tDJovi+wip8r
igHjMztRBPQlwdt2fR7lxfJ4mgpcfMwPLKloUsznXavpcEWDgD5TX4xukeuOc9XBCQt0DQwJAw5z
JMYQGA1lj0MQxiPp5XOQHdIyrz4dTA4mwPe/L9PMi8HhPVmlRZkCgOwPsfMCzeVhBfZ742bSkFS8
zOstqZIfo6zBf/rKg6VrvWMM2+2GAEa1D2YTvRa18n2xyfwzAmm3wFDHhNcHXYfTQDx1qHZ70Cd7
eXbVZo02Z+uG8bmBOtPoGwmSZMgmEdlxaBG/zk6it9QfNgv8hay5k02LMGSxpF+kwTR0FYE6UluG
Pnrt2DihndQiSbmIQ0PwMG1hY1eGxMsZ2RU2ra9Sgo+BVFtc+DRSfiVoKZndPOIQObjNGFYPXrj7
pQ/OXMusbEyS5fNIz92YWrFipfUDn9ShMN6SZTfvPtPwKtCWQKcCNuVyzEmqFnidchfuqQUlZ6Gn
wICGobgvoSitSKx6A2Auo8VGowO1NEGkMIZUZ9lzf2zw6QcYUPmLWnmJlbnlNXPJ4UDoV7t81HYQ
pe7akQzckPSi+mfllK2JTvEEPrv12Oht2oEFhLzP6WBrtbYYinBZjvspQStKH3geYYUtYL1IorPd
F8JzBcm+XUbKS0V/4rEKc/mWzs9N6ligHke955Ky6X5z3p4K/30eLN1BQEML8SWDcsO6pT+x9w8B
Izkrw94w4+//2rNRiZenHd64nGdBHpX0pvRmx29AntgYi0qXVqDtG86aS0Y2oeWxV0e8U9N1hhb+
jaxQ+s9n08QNOISeN08ICdfs7+o2ClalD88ZxjtlkpAKYv1vjN34rnF7CyOQg/o5KluhZNDRWw8I
WeR9OzCsOMEQdD0TrZYCFikyVEp6JwWs9BPTpO5iMjhntIJ+6JbVRLGXi6u7MKDgleVajfj0HlXg
S5MZAqpz5gYbjI9gW/eVrc9h5wysQScMbcfWwsWeURzGcelRFFbfLRCk8q7ENtayGykG7vg22Thc
vwdK3UqRE1YjRczuuRYs/ZbI8lvMzlhLfrnUSwgmZKnHIinpwtzO3LjkyOGj4+/Njs/0rmt9lyNB
JG752nURLc+jBkqIlX0z/HiLkclZTpbhFrxzB6PJ7F98YlNNqAW1dIZJ27j6jTDXyno9CZhkYBwD
cWKEbPXQa2ifh8bdiMYbRUw9yFkmj7hU+LdV26GG7eredRRQL7K6OFPh0A5cFB6LL7nIhxO3xwX0
rtG9upBwOiAwN7sjbZC9n6NWSrjBsRm1NMAQSeMcgurO5GPlmI2GPse3fhAiKb1nBLXyGuK+/CUD
L9JvA3qbAFZyYbaKkZzx/w8SF1KCt5kUgZZBU5063BYzaXeAvrbDCQ7zSdtfDlfq31jb1KdBsdWs
te30QvHPwic/tILtovmMSfYvoh9u2645PYIPIu7BUA+lKl4yx9qoVRlXhE/b7zIPRNjv5L24fcyS
NXNM24DBxHeP1OgIU49ezNkqKNcTOYQkgi1TACtS8wnkps6kZuV36YM97c0dLFdQ38lUol5EOkha
EQb8eaRLIbz5JS+so2QYI5OhpkS6tcVaRKU/7oC3zg/kmDM9o5N7TXlWNz24drPmshiitgwUGicg
95Kg0RVwUeE9KYlZ8oi5f4f2A54ZlYk5nWdpINVAxqRFrrx8PfsiVTL+rdFS/3Q8WQae0q6OYAuq
yqLxk7qge/Ndt2OXZ4gQDUFXzKs18Ho1k49XHS4jnxqLP2p6q4XCxxe4ReFM+eO+9Bvd9TSqeRqi
d86pKvgF5H98AYQuJLVlavHFh+pjTlymFr4yzJMC38pHUDbHlwWXK2A5OO7yVQ8kIOHgJ4Z/es29
vZoigKWnAb9QLI3VG3x00nsO01PN0Pg17rq0DLmEyN8plBGYDkRbjxlxFHLhS5groLAXy+1amYnP
IJwCDSz0IBYtJED0D5ITb+BPJiZ0w8hyTSsNTX+goEEd6hns0YvLnCFIuWj6Fu7o5NJx/D2RtgLO
8UkxohiQLNtJwFvThg+tFZYx/EiMRaupVWsxz0sVRrBWS7s3DuS9CtnKw6DHoNGKmbfoU8i+S/LD
0LccBtkWyiy9U4p/Gd93hBeomrvk8LhAeItkHVdl6fyQh7C9NrPh+5xO14tui22+Db7QmHSh2wgg
Pg5jyGAJicUwb6kin3wQYs600EXWm2aVaIft48n/BCzGA0k9urFHVCyNRR8Y00TEKM7ceJBt5qRW
72qZU9r4QQgBZIoKOai7o8VOI6EIS4LvoSpxjjTdwrAEqDEZnESKhyUhjT+Hk0fd3c9PI4V541gT
hVFhM1DTEn87ELkR2t4505Ghb1AH/trv8wIsLprE8jvjLnyAwTno8hJQWxIbv8emiBUKzsl3LGIr
HAqGZHxyPXXFOsLPDr1vtM8b79dW5k9slkA+xYg2dNgttPCLw/66VKXHdCulUoLwc/vyue+fPVys
7YWUZMBaMJd7snHZI8fnRyF9UQzge5W94lXopHpqp+aINfJ3r5AeAIVk9j2cbTvd7WrP2q/8VPex
/DL6ScdoKDHW8FPfwCgI2pfbx7Vbv9VM+sVORWfSg16jgyph8Q2WmnGpHWS2pdLd7tdDP9IqP66l
BNP/djOE6SdLBIxYdJFzgfiVgQ5QOd/0+1TAHN99cEXCtToLgEMIO3wBdZwSAx9GGoPrBjerKTIY
oD+vgoupDaFzFPodbKvYOcz5Tbr4oLFw+eKH/I6aiMIbEQkatXCZ9oNc93CPBduRDchWmKMbfUnV
4qqXHGEsrGr/QPjBM3ZB93cqwVq54tDRuVrxVPhHPAd/SlLhKj28DU+xAy+tgx7+GBTRGUvtoGjS
A1O9rV+2ScU6bvETptniUS0sp6iLhxF2G53ZPYsfX4mIMElulwhxyIZL4iuX7gDOuDvdSb+lu+AB
ICRaZ8rwksu8uHoJrNnJtdoLj2Ek2XZ2tf/GWv3Db96zaRErVnq7ZjGpgH+keoYP/+iCsQMNzNBA
qfp2t7La0tHG2V95XWsSJFVko8jgsr9KsaS52tfIqlMShj4BFgOn7WV/HIzhZukBjLw40qDtNTTO
M5WwzE7S41h0HVHZa6m8+vVH55Nul9HRWLWfWuA3B0u5qLaAt3aqWz23Dy8fdMyQVIBbaCHSyol0
313AOTpSJnU10H8mXYqp3N9JAMF2Dzyih3bMSXK07peRZkri+yl1qomTaAjBD+gFr+y2KeE+Jo2s
bMxlyy+dy8ZeFEHC3+rvvmr3fFlKrrrW00jlXx33hAFj8j6nQaxbXjCUTGjFoYllHtY6sFaCYS5h
nQ9gSW1vGu6NfC4Ii0jN+Fsqf5JnQKKTwfhq99JKXowvGf4aQsZHQSUOzYw/RuyHnIqD4b8R3qSU
IsC192T6DCwLp7jD1UHxbk9cSHAoBOLu+WpDDTgaiW6OmOwbJAL/HR3Ao/OAnuCGVwRhhxPDNgu5
+wVCyyL7154ofMqseBedMqsGESkOlHXYTBVtpivR8xHRtC38K1nfbctwpS385ejnOauerN0mhw+G
0X5vyRx8HS2CXleYTYmP0MC8qFPyI1eqn6+Y22DpQbVrV0OgS2dOrIxDDIQudPrJXxjFmMx6lrcs
yenwhzPyGWhJVsSG6HbW+hZ4tIQ5+yS1lKVoXtQn8mKwo6D5901LeE7zTSGUEBysTof8+4Q+tuLa
0oP1r1Zz6fFFz/lnPsKFtZ2FadOia3DuTUraiAxsxLeoUmWSq7U6NldjW8AKUh0ZmMFLT3qJIyuT
YnQHkKFgsmR9JyNNnKR4Guwmg86FSYYFDaMzR+PYDFb6UdfzQFLDKjJYja2TOGHWF28UH+NT823N
6dogYPZrE6BBqakFAbc8AKzDtpqJIEZX7NC/+Ow5Ie1IF9hEDkXzoX/KomegmgtmBA3LJyJPS6ra
/U0MJFdZmkoWuDNaakav3nIytgiliWGxs7cT/eiaJq63Dl9E0TSiplQEXutoJ0uQK57FUBg/+a1z
Rj9f0inhcdTE5nGaWvJ+y1mWRcemjL+FRnVZxYIowcIxEKXEn9qMaOjn13T0+gEmQaKNPoHONLhx
sKrvWqShUKc2G0+OD54d6t5wotjLVK4KYWWpEdFZzsLSD2eCNeNQIZrvzzo2vzYoFXGoXoYxkXy/
3nmDx5TMgyeB0iuA+lcPtT/vyuWAivHHAX2xAPB0ArAXELd5+NB2ilBpnXSK1S4EAJvrunp1uJJj
+rf0fWmmIWSPzNjrv+vEpNKLHwcO4HrvtFJ1oguPKFq2cTVRctrwD+ujscPe3L8ljxRAqkXt/R+i
d9AbWb4A5vo67ywcNUhd6xke1E/0AOm9lZKC8kVjlU6gmYQ726lIzk+0VoK083fYNnnoE2xMxxn7
HvWxQHFLcGnEpTBYZYJuxpL1RSAVaj6tNpzrzPQi6DBOzp2grzDXACNuRFMrIEBTqDZetyFQXEw6
72zN1lxZEKtDPN6favzIyIOiK0cy94lcecSK9ef8r2ggZXf13hGMyooT/YzgODbPH9R+TYRQUcaI
PzafB4HbMe82X+dXAmr+iOhdkPGQzlWKPl6Tr5E5TpCtXZBiAQ3dekoTr6Odz8tk623V1MNQhvh4
AKF32n4ZwPepWRIp/kg8upFtQYhsEr9fr/mML/aZK1DcG+oWTXo+7GxCw77m+VMoTkGUO57Ck8lx
5Gou++nSTwfKjaVcjlzwtuNmQiv2ZdNNu/HFcdSwrnesErbjO1PlTw2Ry4y6fewQ6Liy75qqtx2D
jX0XK4Ta1e5x4KrMUoOj/1/AxMWZruCV9P1rRONRp3PlAMv3WdaaO+JQsafx/8JtIt1f15RfHt8W
PqvXx8xelg6nIbaeY0KxjBfUn3lorCriDU/rn35CLdwsAoLw1d75N8f2OKkwzFn0G3I5/SYkPxqC
a8LAI1JuZ2uPtmHiUq1osQw1uO5WUGHyILQpco6uorPnQEWy1Cmzuc/APaupFCYhG236eFCSnXiF
IkTWuWxWgAxTmFlBA01iivtvxp9roH5sFem3Abv3NlIZFGda3IWXV7u9S57nuPKIxAxd3cuuu2de
aMk4eOMJNE+/Aa/p9lFZa7JmyyQvo727wGwk+bkmM8GbNF2vpu3fsC9G38gGGe3u3YcJ1d34drDS
BEaOV5ridcg9F523lCJeFTA6/Gdb1ZamayL/LtA9tFdf7ZIHIcAzD6KdFW34HEvep2JZ+fX+zQ3+
OZ6D+egALl7DsKXMjzEowisHtDJjcocPhF+M4d05e7zT5G7um7ycB2a7ky7IoSSb9cCtblwMAXKr
1xBOaFeal4Mz46P08NlFoWOe1VrQsxv/ZNleV1shKIpOlbK3U+xIrN+QQd4DZJ7VOc3X6NA9Un4j
EAGyfqRRb8gxV+egH6xHLuygvBNRsJ/fcSi3uXyvRC8naTv8dwp1r029TVHBimLnXK4WGH4clFlc
hyrdPDT3XCCXzilJXQlRzTGVJ1gXuMOKwrIOdE8KWfyyEA0dEElvXfAsYy0oQlDFZO/DuM96NhD6
F4Tt6bAwzg+Fh74rJT74eXdoNLspbbI8aHDk0e0bEQD56M14EUeGBpjdKlkXF0kLsUJdO4OCVjnW
ie+Giweo4MTZSTpGj9wBRDwUbTIT7CEV2WZjTwCTlJUsI8hH5H5JG7TbTs66Nf8rNddX3QoudLT7
GbZvOyDXMw2ca6zlHgrPCHsTntzQ5aBtLnUnf+Ixjwg96R/RYVpy/vZZIw1DOFjcz/TATkZpj+2K
Vl9Cgunrs/PXEJD/RjzknGJnolFjxG2HauVFn0N9SYP9lrGRT7FSdRzBJPDsKMoc+H8pPWmF/Fbd
sXwKqKRU3suHWhKuF98h9mYs3DMbP+hqB853E+ecilyXpzwRmRBMx7EdjrTmV/nZatoJf0cLOMIA
l6VgiDTSPwOVHNsj9akbl4hf3DBTIcY1WwLEKe5ALw1/JxHXBxK8MdMq1DkzZXzMFahA4eSLJ3LA
zEND0LVvsqIT02ogVoIkoiHx6pXcRY9Bf5wg7iZXhh6ElJRPo/Fq1A5JQNu1z5TXdqbYQ+hwZ8UZ
UlYXyU4elK87t3vpoUk3nd5AKKkF9QzxxuozzbeFocwDOTM8vylvCzDbbQtRAWT8k/qmy1hoZsrH
r+s+EfrwWtjPpJozqQI9/moCNTglexK4hujp2qpvOssMfaZh5RLXGdZ8bJavOMuKgOoygcuO6H7/
e117CHUguO7y2PfcgI4jBqqgFInfHB84r/KDTaRUni9USx7gDbkcv9WC/Qp/1ZQ9QYHeYUDSLZkm
N8Y7h9ZrRgRiNfUizZN4PrcfdD4KouabaLH4r8jBadj5c60cpN0zY5lEWvrzAu8fTSZ34FXPKrYq
ghlJWsuf2RdzW2LwzfE0WLyGlCSJrZd/ljxScJyTL/298CzNo/1QNETkt2ov7dV5Cmn9FK8/THee
Tk1AZR3E+USGoh0rtDr53P8yFnyni8aLOOtjrgdTAk83r9kQulYIbnPaH35MfuKzCNrejV2h8dpZ
Bfhpr5Lh3IG4S60nat5kqH+tiVXqYrvD/rEn4V/EgWMaqSo0KwtcfkjncG2kkNkdSjK5zbieSHcP
GgYtHttBehVlBmOodfj8YLinhhsuh3jFlTN/VUXZUwIJtTEWb59+4C2s5EXcZvxB+cQ65rLa7ZIJ
eHigmg7RSyr4RA3rUsyH8m7LxSLLnJh+AfWIe+tG7ka9HahWvJS/Iy1uFiZF/wVlmAzZw3fcx6wy
y5yFpcl/OenDgIITsqhBL6A04Pd0ByiEJYwzeI32VkfT1SxpFs4cEhebg5ITXsxIIXr6UW1i/UCw
34XiPuECRQxYOAw9QbpcN+pXAXmpWawTiLS+xcilpXYAG+drAvz14xUYvxjiO3jOkFMSnuVrJ2Pn
76TkmOju0Dkk2K3Eu7/qfesYLhvVwyasihwgJfRYxAMgM6eF8PexiC6uPMW5GAWp5aa+apmrGBnh
doE17AwKGZbYehISH2UD0RYePumI75mmp/hhQEUqGYZpOhYK03d8jc6og660wJkJNxSKLBqALwL6
l64ZhsniH0ca8p0gk6nt6rzJeJzZ+shrpg3pX60j2x14qfuZk2EagzwbXcEcZlD0wa/dqGuRO1bn
Y2tjPyQv53UT98pN62Rk3V7DtvYK3l/+PTixFVPzIILn+YVhdbMLk/T9LFtoJa3ArMuL5jk7QAYd
UTBWPGp+w53zMfBvvMWRHVweDD8rvLNI2iwk1UKrZ8kJ6OOttmU6jbz/kElMauXYDI8H7OIGfyyD
It9/U9ETDgq77wA1Rh4APFIQdBmm/EhVqwHqX8Z5Jz2dqklV9obdH6Y36B1VF/ddq59wxNSXCHAl
X3C63F8q1X+UGUn/PkmEu96k2I2NPLyB79l+9JOsV9d2ohCbo3yVULDdVFB54Jx5O6qZcsV05lqE
IDZZR8b6XbnwG+T/BIXTd1ZfgBxSv+lYIT5aM7zt/HhqJIwQuyGhhjyNdr+rCYQ5RnARS0K7XQ44
nq8pQev8SCDZ5gTYaRfwoq9AUIVqD5+gJArLYH9B5tuhmG1VlBTSWV6BIEboMDuvfl0L/ft2/uS5
zrktHV1n9Ap42MeRskgeZPJDy1evPB4uhTE7XILKrHYERc+u/burhCaVnLoinuxbQyN0bd2HI4GJ
OXrYCPqSoQJYqKVWlc33UyCwOjtQCIJQdyZ6Ey5jKj0djge5ccCvzlNVKFBIxoONIyZ/5Qtd1w1Q
p7RL7XgjbKC8h2r2WVaMp2ba0flBcjz+i92Lagh//PZ1L02N57qbSlw1mzJc1T0TIt2ExpGC7fJT
hdEva8dJ9tr3S9NGpllQxnXhYNMapqbtrdGuTU0BDQ7lM6OOTEOTqbEEqLofPp8sdCXag9yTH0sH
eFEJRRSonQ0+Zfg/8/50uQL/23ehWMNK7yyzdygwDieUstkLr75SNUTQg62Yj8SU2wMbi8AFc/vP
KaalCCUzmSbEQZIw8EYzlUaUFbuvwFi1CoeZAv5bhKC7/wp8YWHNQEvfr/QQQyAWp+ngW9++3q4i
TlddWGLUKPFlHpEsC0hppUDgMmIXeqe5Ffxuq5zcK8qaqFOnTDhyg27zE/MOV7Ws5UANiNw5HYmY
Cg8qDMqZUK7ruyRUpMAM+hgCVKIyAo/sZfph7IPGqFyeiiFcT5rSsXt+9eDaGGZnJerJ1PRnt1nW
NZzjXi91NLXBXqAcFtBXixiaau0yC53bw4ZZhyDw2UFMrX2w4UmvnHkUX0Zr9W98r9R7iwtzSt10
LJBNrvt8lG/mX86JWPkTpahGbWUStTg6lMVdGSgX+1x3oj06m17/Xiv4XPT/UtQ2uMtIh7QWTNHe
dWdXGXj70hJYO+TwNwd3Lzk+YHp3moaKntOS/aSDksRt0uv/XX3bqtY/iIhOF7CIz70c8/8h7uGQ
C9JevDZLZRnUi0sZyOEtII5J6zJn3rI3GMkHtB3Exf7aWxeWnGUiTXwD5LpyvmaXOHo2mJZagPLu
55pRrmdWCT8kZgsGdBipLGZnsoDArDm6HC+kGWy4ijuuh8vAR1mN4jfQWAIbKk5CpJJ5UaSvyeCP
XPPZ9OF37N8fJZqUFi/Z4RMEqLiUh6NwZlIfy60y0/umF3HRaN0LjZnspBGPQUsfXtYgjxEV2Frc
UomQO90w/fgRX++HNXCPbWVVpob0RdqN5/zirN2hebMheFogP6fuaHFKZWEdBWk1YBdbNd3Vp02Q
UrxSS+NQKUVUxIijmdUF3G55/Sw2XbTwtddjgttIAhiV/vA2lZmyhk28JQgmUZZycYctaHCfQwxR
XX4tmTi4nUZrYijwfW0k3AXk9AGNKDjEyCHttmPmlKqAwqcEJI+y0NGKENNVAQJWSa43MKSVyTql
x0/88E0SGi/37sS5O0m4uukaeLM3NJatnV5INSfW3WwiUK+Xe2ms1/TAZQfj5j4g5/xhzRBhO6D1
Dn7pvuCYksZ2sehZlN5BDdhIYISNXUtCC0RfQ6UM9AuoccL24BnTZx1MeXVGCgkvh7d2KOLKA9rQ
xtUC83fxdf/9rybK+xKJLQEt20Xc50PjBXUbG0A15NXsz9jtnONrGOX51YIHkHoQnkFzBEhg4uPc
oNmlWQMLUd649kjR/bTFlQHFsHDlwxYNkdIJHg9mWGoEOLfIANuP7n6+OHtQ90xB0LFe2eKExo8n
chjBa3KQ54ljdkw4RsWc0TvZEJOSURvCKlP2RkHi78APTZwW2w+jIuQpBx35ji670fGOE1cE0Ohb
Q6cadm+pd1eFlgA7cGgL9FfyegdNYayVw+P5Dqureqpbf7RIq1qMIm8X8gHT8c8xgKIBfJouUn7y
CfrE6/2ZDvJFuoGmc3dipoJoZxS3R2mtw8tMnV+L+zbRrIhEnzWHIEUJzQwZd+6wOWkhDJeqjRqv
yTQTVUbNfIZRCXFSBgSK7MflW0NWgLRPxZggQIK86+8CPwyt0D3XtZhbuct9ciWvHHgfka/q0I5S
sbwZCxerf8RlUfkNb79uaQGn06zCQh5Emy9Mdsw8OgVCP7EIR/REZ2RQDrIBCygDjbS7ckvdmMTH
mlmUalJyF0ptzS9R1T0LCsGpaU+xScVqkqYaplnM0Le01GdAkl2g12kOFIL/KbLIESWG/tFtQezo
nPo8NQvWCsfH8OaEubb2pTwV5A96z8olBwZwSOgH0RalHRXB1QkiDRBI6PdxCd3VILY0SY3mph4H
waF8aKULB9T6RUDZTG/QNMDjzGLOwTyya1Fl0X43Jt6eJ5QegWwT74fEs8BHL5k0kfkCZuwD5l+X
TggiZJiRT01TuT3hIB7wfbtFSPTWhcHquN992RwwFSeQ1eGqhXcLtsNEKFYw9AMw11fRymRrpy15
hAoWY6ZWDM+Yh0HC2bbMHmEjbfuffJuUl7K81yOek/C0xDWjj4Yo4JslN2d5Zuukf5U43KSshKJw
mUan56Y6LREubg6sEe6zwNMbCg1Q4PR1yPMQ/hVPloPRKTM8nxKHoX+13GjV8UfqeQg1Dk9zFG2e
PHfNtcy1nE/BqIydRmNqhAIuslq/ERF17WVHVhV3hcsLeMG1Mp9tB1DZ0u0isv3rthGqCHS+zoyi
gTtMLXJJWXZ7lNc/ZustbR/zOeq3+2s+eE/zOqiR10iVkQ7Gy+m8T04/puqCbLsWC9CsXS2FUlge
/IOtVXVBTDXpr3VEKCPeeBdtzn63jIKJHcmXTKOUyoDLSqYKJOo3sEpc3zr3YmXs8JVPQKhXJqkt
ZwCK0uTeccGSkRjCbVEMuy1oDa5qs4bDnpjTLsQyLETrGkTNDyCPoQ0N3wmydbtpfFvpstnuIg3B
UX32GrLQuSxnA5SyWb7grfbCFVS0LREOMSVGi57+TBYikg02BPS629+GqPAQAdr4/qBtCsJXPubX
lCQgND+j48IQjEpNsQeJGqeiYqlYSX4iGaBp8nMSM/JgZ+MB3sNfoqp4nzkAxax1D1o6te9FxLoU
/kys26ojSQekwfxjhtqDWgw7gV5A0kml2aaAktTzHCAfznooh8RFcS7vWLYsZsS2ezLrVJp9uxVn
9g3CDWIVHBWsGUGyMmNsEunMudPq80FVI3ogrtkUUUTwqCzW4hyal+IE2+VxL9APwAMeOkkqAStS
r07MebSbhGhypmFDpjtZrbXz/7hoM7N/GYvi05FG80LDGtKoHmXymMoN389pMd9NICRPzrGgxLZe
aosy4kaSO454egYmSjie4tH6z1ZFhSj6tdEq+NdmNkPnPga0k/7aXChdF12kWYMb0Ra4lOInH78e
R0C2KGCHvzfCszsyYigUuOQpO0JgoSAmzhN4z/dh/Lt8QnfPtZSkdh5lSnHbqPD50GEGwr/N+Ff7
ZpjJ/BN4o3lqgYGJUay0CxcOCyYCCQjwGeiV1QbK5r4ji3e29rHI0n6Dt616rPLLjNABGVD/VO67
3/MW4iJ2WQ/FvYwNMmb3E7h0EcFK9zguD4OZ98Y+jpvgyUOtgLEVljhJQVkieRnw9SEND8cdey2Z
ZgXpz4a0KE6SJfI4u+6fPN8ToZUx+br6GdKo87i2t54It9SMjZGSUi1K9eCzySQg2GoPUoItLvdf
dvNB3uAcZCrwEO5sMBhJiU6GIRO5liqoBON8nPDi9Wn+PDR4m8B6hEUyLcsEK2UPTdAg29+mQXB7
u6+IAARLXD3KHnV0zs9LDV1SBONeXaILkHL41PZptfqFjAqG3SPEjsc9WvpA1HcuFiGNTBkUVnVw
ezWsQpF6TO/CtVDGefCGSb153tQOEII/I0Oadr9O8qgEGjgLZzx//VngFHWRSwSaG47bLaFbXkk0
pl9fj9RpdWl/PNTEimZisFnb5NH+r2GjYLM24k4qWBc5HGe+4tDeeck2fVIGPkr4Dwksv02IjiSf
qhuZJCLFmMOmQzrwuwlXqBiEErO9wzXque+MzzduQIfP0i6hky6l68CrEard5KNRcZvkNcr4JtSU
N5jlUWMwQoESV8b//BwpBEyBUxBHKUD6j4mXuvZrPoSA5Gqy482Gp1Bn5My1VdNbEedgSHvK4VNk
gpFrw2ByBrWI6goF9RDh3EvTs3k1vnL1H73EjUyWGmNLDaflSvHGJhDqAu21poliQDumetnfaTZB
GUPzto7viNONlUH9IvaRlWhLsc0omWZ2GZ6BtR8z5C8g324IUbM6Fm7i2nar6OOddZjT9qsMZKll
IczDZYtnUoy+hlIptnxjAhlgC1FCNkUGL9r+fLX6Ud9uf0TZG38O9vYnixw8c0ZYvwCDNluG9XYR
Bg4Dqrd06/jCUxclkxZWxiACfAv14rOHfcBRdmc7cFfbYohTQ/HDoYNUxiR95hCN2kFMgAAb7BQb
S6XxltSG0fU/Ubee6GL2ivxsom+StG3CwaDxI5+xzsv5KycMf0rs8R8PDOB5qOtCTaviXyiBkAwP
VR3vGqtl7fVpgj7llLMrIf3ryEGvVtEf4bnfdQ3yirZ9mwf1vFoaiIC6oFyMWTSQU5y4t+uPvZTI
TG0AW68a6QMf9bvs2XTQ0226c1eh/lUViKZolwhUz3dFE84fPUAJAzGDQuymtww0hdSD2kajerkl
oVWwkHoViDISilxqmYMgdmfFjKr4jAVz2RC4xWsmk+IUKKGTmgoMCJPpfbDbGBR+E36I7h+cFSkK
IHW50LB8KDMJQ8drndbyKFmBccYDd4PVTQT1hhLHzzU4RmxDncjvTlyybVyDMymvMjPle1aKFYXc
mssTYYvLE4E79zg15BszUn60tjqooce1OiWZrJHPb2aRqR1vQNrNMS51LJng1YAyo97UguQ78wR/
ghpPZWeZvIABVxc1YQj5kHxPE6b7+f/bT/lwyXxd8imaGC57RbdVT8NbLp1vCVS+DNGnpVbRiE5x
OimyOONJXpL9ldr/RRlJ2OlQE3DE5EOkTk3i97LxH1feU4oVu3Ar5YdeuGqHdZ4ZRD9rsZOmGNM9
tubf/jlZVgolSpFMU0SNT4mbdrMGhSpZPhE9ADCOLndanSMljYpA1yK7KgTvBjKS8ZqXsyK30O+p
smKUcHeyVz59ADUSGwa7xFMA3ASQoQIXwK9IZAlZhyIBDy3LcF7GIsF3i+3YvxXaaFGViokKIHbd
KT/1VEPigJQTA249Ks3dsMXIe4FAeaktfzP6u7daPxciI3lzZRH3lAKhhy9JNAlYQTVX4HnHxDml
Zgtc9LjgdfrDumDTkoEPvHyxFWUYMDCH62ry0ig5lfAw0BwLL2z3dMxd29cYb3nXFH/hIKBvFSvz
CBmmMqri6BTfTne79/SuejVnMDzXDVkRbA3W3a/NlPcrChIZ8SsNvh1OWVySL3tEyc3Sk/09R8eO
RwVhR06TSmutc5LRWwrIrVXdxVtoE6o6zxGHQkK6zCtMHy4UypwRFSyaUsRW34e0DRK7f8eUWzG3
EgQaePymJ9gsF+ztd/AO9cgOM97xy/mP/Tn3uQVWx7s/f3mP+Gum/6PrF8oY4ARE74xifGtT0zJ/
7+HI2L9nlOOhFPOU0ql1gCe/J9YkTvHidztqZf45c3SowuIiOXQZSmPrI1bC2ZjN838QK3yVyNUR
PZ66zXiLQFCXt78r2Pu2NJvULWJY95IbCMFhyq1w2ZAKnD0Zr9MreiRGrKsMprhkR44XlSt6jsu6
whV48IVPFEWJUS1jzRfMl4vo+uh/EzkzmyB1m1BIzyrYYZbt5t14G5teipvsK3bmrofCV0/m/LhP
fpzzt6UpL9ulrEZsP/QcRxL6dtUCiVLvnWUG0Ig2FIRtQD1gIyVZuLz/vsVul6wm9hkfC1+ocsXh
yFLJok9CYqBVpSRJauYkc7NbbEotBVdcUDV0m3rGc+WH4fHhp0CWy6DNbM5umAwRhoiTRSuKPtoH
ZTRUYrdm9gbyQPOXwi4JsBQ5veocX3WPPv+SpTdNCxMpcUPASxpnpnc12fhosfKdD8HJ67SdxE/L
xXBw5fy+087yZvqV/iN6d1JLOyZS4lE3f3io6rNUeZhQ/aWfkn8rd+xLg2RDhNo+PGnPCbC4cGvE
DIPsHeTVoMABXtB60swyXNKneJbnVytetwlGgl+dMSXsS2H+hmorAzvCKSlJujBZ47hNbyceIsLT
JxhPoxZY0WR80L5BkQum9XvEvdhiqBQScitI7VO1KGMRaaLY6mXfRxpVZxNVOObVHR8DKi966/5h
eArC6t3t7hRLIQ80zWQ6Ws21+BxRrWJ6hyKN6/4Zva0LAq4wKBoLfLcMKVETCnJLVi3d0j2uQ6HB
vlJGJF1jMmjX6o6AfO+E79kQ0EnTLTMus7TtQuPgp6LaPCXLJvMKp43rbq+8Jf1MAVHkCNXjep3U
2nS/Qq9h741Rp4pYf6SKbpVa6sHOW/4twrkW6kIfrLuM8GbWc2y6GpWHn9XHiojUF7YRQc8osewK
4CdkSlFAU3VrHxbRxhSw9RXgrljCrxBEFWDfWGTZ1O0c6llzCRQsHTaNNl3uPJUG+OYPjTqNfAwz
G5wGif1m4VXV9i0GVy5KoBowjoi2ZmwZmfGA4hw7skPPyBYIAmsUZ77Radr/qmYV34aIhaGONlJB
PZIgYmB43clNS6keQMinjfBWCOBw5dJdKOLzt8wF2irqplL9DY7CqdnP2S1Q3jZWZo4IDQEgucME
uY5EZ71f53CZTV5bAuSVmAhCi5o6YzWrlkbcih1uYasYbqxxHgH2DJ+Q2+2luJnbjCcizBi7SwsB
phZQfgDhQOPMFYCXe/pW80sl2nSd9VHWoixMOHy5FeEvkaMtlv28SGgqOtycaHM2t0BNnhJtRMsG
efEtkRRJkxw2jOggUHb+Cu+Xrc0BGQaLuO4V0g96tXzjWazc8xybFskgrwJLXWVORRks/xJ5et+y
gEk4QEnpMRFCyA2aT4KeaD7W0zc/i5QS49RN4aknxQRz0qp6Yf5CWBeimh8vBF9rFZ74jz7uue0Z
WVr0D1sXNBPobMRsge+nVBlTgyeAuFOoP/XFx4YSdeqAAxF9rZP7hn21689FxZTNJ9R/n+fLiT5C
u+D7ox6w2gUPqOMgRidFMp3zwHg6wBbgeyqA1RsY6DFSzYL4zGsekRAO3d49YQPCN93RZZurNFJg
VzsNjyQzUND6fT+2Mq2uUXUgRhh2/ykgcnfkGPtjHm56GmZs2Zao/GzhicVFdK7w+i2dZxPHRJzj
MXSxpLgv2UtrKrTqR6T1UEuEHs8JPUe7Qe3f2jtzgQ1BoCLE1io4HQpKc6c//KXhfgcwiK9SqHCs
viqN3Qlfx9hXXIgb7C5yFVoa6mWxO38OROGOS2myb9rKGCx0M9X/Ag7ecb3QqIpBru3bZhTdFRgb
sf2lMEb6oFKDXyT7Sl7Yoer5dSoph5zadfF7D1GPhBok4GQq1OqVtHzLnGXpXMZsLgJiusbzxINt
EYzzzDJyxcaykzWrSonjx9vKzDsscghmRKOJw2eQNd/YwKHmgoPuSK02EjinziEKlOsIpwMrBLVy
4A9vxNNARfsv6qn9wEBc8MTD9rWLtfD8qP+CScphMCrmmxOwyd7P2Ucv88AN247zkUIl49NsVfg/
O0nPKobZeJMld2WiBfTtJQqSC1AG8rTwQTUn+ZF8mP2tQ6094jXCNVpUWuE059so9fz0R27j+RES
z5YynLlcjCGWRF9tyYp+6d98D42dOkSAuCvycio7X/SYYkZTVJsilaeOuvOs0+KAjPsn5ltXhCrv
eFXCHIOYbeuv/Cc36PpedCHnxUnxBiygnbgtxp3Y9+caMivxgPnq2o2Qx5gzrjpRyz5jwXTWYkpw
YIc4LJqolIYWW84UDpoHi6k3mAnAa5+ANyFcsRMdvq6LpxrvxAJ1eCp9sKOwuxMcs5fugVxeJR3a
DOji/YORZNpoGlFs1EzN1dXisVBWGZIOJAzThFsR+HOWfucAHssPgRn6PXeaIjyFVTsc2pC+gU2X
XscHQCHnIZzrZpOMSqXhWhg7tHlDBc+Qyeox1HJcAAhPsUitGyJxH3EvuUGsanCqbFTHlDjcG69r
kdfkELKnrv03tKGGK/OPmnwB77yOG8VmX7uPwyw+1F1l9zwGfe6gJNcCJOtlsEypevi5gC5pj4jZ
OP76SdnQWkaY87s5SFnKu/nlr/oxh/xQ3XmUB7UJ3s8zCzJG7e/O1pWcB3CBvuvbhuyOOMxsTE9W
4qFvJY6bOsPGIgZp6H9AOFRdahZQhGBxN7NlS8515UZQ4gnJaVUNxS4PkEG3p8vM6wffVRcB2ktQ
Ww8MfX7qtoth1i21hWCbD1HIX3iTBZKqP48H8MSRKTScYqXpo1mWo/Df07CvrLjH6OuGJJi5Ox/j
K7qGRnxXHWM56XgWcy54OY2zZAkhTBesWKiBQcssRTL42mPifmXYAN3pJzHXau+RcBPVz5uNnX77
KfoUh0P6c7SXYjSovnoDdMqmfrFiQgng0CHHIhZL/j6to3JsQdYTV9y0ZKTlgE0hp9p68b8kcqd6
2/1GU6YmZTLXzNJ0MqL9zOVMI7Jte8CY2JzUJxuQMdgElz9zsmttP8qe0A9GmbO0Yacg5cJYvHIU
n1m9kjI0lQ14q4z3LAMi6igKH8rd9/QHGP3ZmlvqWiWzJKMDdBBzQeY/3y1+nPCXQYwydlKXZIU+
/ZDZmKZ3j5ulpdAix2XMNs/SFkpnY5CMPmCO56qT8qmmdvlvqp6gVZgQe4q8NTet/Oh12POPFZWK
8oldoAAD9NeHsoN4VN09LDzMorxBQAUh8TYJes9grMXC+KZZdFPk44IAmJLGswvCz0FxOOYsv8hV
6cAXbtwfYmnbBLCySyT66hsdikvwv94TVnFl/yqixEy1ROIVWJWvAanLhzKF+ulEQdve1cM/8UNl
nl3yjk1f9OE+p8zz5r+ZpUwMco15cy993kmE7B1D6UighvCPwrIqWFwgfPIBbbWCkYECkZM+TA3g
bhruoMxqt9WuWY2zY9rzNaDZHTQJGa1rMjcsPqSHQBcJGKg/wcqlto5HFI0pBbteD4AG5il1X623
OpKZI7/O42O7uSKTbbkLSe2bNf1CbDATPeIRpOOc9ctnF0LFmG8zqj12/frhHJ7UOJbs+rfA0n43
VerCJwJ77XWvNUVSJWq2n6m5qeQgWJpIztyzBME+ZesLURahrMJWKHVSucSj0vIS7/7fcO1UdCzT
c+oZoSR9GEjfy05mhDPLp7J9Snsqrsa6e44xIg7fEKzDodTsXFNjYTFvZvrAkho9jnQHx6oMFsOS
UmWmvZimKOqhZxEg1MDGlFtz/uSZClQeO4FsC1lhgbMFLngox+KEVrbefwln+IPfCyIOmhEAjxuY
d434TSTqx4Qf3y1oRG3bd2Xyj+NVMCZyR6BqoWdCk/wIvUlfxo0AYLy3PYpA76TT4syKb0UjSfoW
qwKgwlOEhQztug9ZpPKYIYKmlA01RPhZcuH6GW6od10Y7XtMlNyxNtI8MTIPLo8HkofjA/cRkmT2
n7U62y7Apsr8DPjEPHHyOqug1Fit3iktlmp7Zp/+RZOqZEzZjQeic9rW4fj+C4qEtSJ+Zc84rbCW
UMEWC5GOb6miMLX7F0BA7S8TVqAn/BEfJLcnS0oVpo5Yke4UJGKV/u0I5LGuzndMqYaxInbAJrpR
1kIYjiuW2j/9GTj5+dEkKzBd7wqSBUHfb+aVXLUjxewfK0Dbaoob70dEDpgMenMma1wHNdEiN30q
QudA/T2SQLgk2wbMpuWylYHE5KohnLNmaxieVSzsIcBgP1Ylj5ViX4VsFIAsUGzk1Z8WtSP9xbkZ
HdQsyTwtcMNGRNwRKDquM2Swd2hkJ8lJnyiRMt9R90DSfCwk5t0VbDYXGjNDDRVHFViS9STjOAzq
8wJePUZluMdQjRCsSKPJjgUMWmhsPmvAyvNySuQ5bE6Yv+7iovjIxwnqDwmEvJ2UG+yhj1aKGFwH
LoWXt7Y8yLTcCsVA6tTwmbDpCeyQYnrn0Ye5KgpxRulyxFNQnn/a3k4yAGXCJiMT3UPEzRrQHt35
ljatGaYU+t3oVmK2anqbco284VRziAwKMTQHxP2QyjjXPh5zI6BLBqeyIBPB6Qw35B3dFVdnNF/A
EXA/BUO5meE5G8xeNtXMdNDggJ9uxAZAvSy5XzXK1sXrzw5D/DNdfpDDDoa3eMyIc4zOtIncAISQ
bgeRJIbIBYVCCqpgWQwuPujL5F4OsrpjCpHrxsdrDF0DPLAF0KKUY5CB+IKbhefhEauDd6rRJxPW
R7GaxTaeswFELOGu7/XDzkoi5nnp9vcTmJUuRTRJuxqNQ8EAVg25066Oelj3wbNSXZYQR70RqdGF
S4YZszLOnC7FnjUZYeydhFgMlIoli0wnU9+pe/iXOCDnfczXF8RPrzSjUbpXjUUjgXV01bPsL47Y
0Wn3vv5eCImSRtGafPCCJievbzVRjJhVYEoULSL8pLuzepWm1u/fBdlWM/tPDteOLEdzt+nOuj4U
z6IR6fVqDLlk+J5akh4tjIIGzA+3/spDHn7Lh+ywKHZ+p8Dn45xfXv4+e53TrMd3PbcOx+52HJxr
LjO0ypeP/aw1oSGYPwzrM8G/S+MUgEEZP4BaWUH1ZAmycSasL9n2KDg060OV0mfQWppW5P9jD5pr
567p4TwwokntApD3CL2K6/q0bR+TT50a9se8HEtwcONByGOErWu1U8ticPC/ihHv9qkWkpf6AsCZ
QcQSNdZkaOwC0DJcUqQbADv5wu8GWpL9iFhrdmJugxUfIbXZkwSlkb7OEKMiZVmPANIcpnBDo0JN
vSa7AuvnM1t9Abkc1f4phHmL4XqUJ/FuakZlJrGOdEahyns7E9G7jpXirrrhjDZFqSq9RLjsoQP0
LtTl/coL5OtVwGSgkrzP3mB6Qlc4n8XeqTrQ++pnOJhXm8Yc9WO96G8rRlJEstJ9HAQFkbW8Wl2z
wbcYDVxCewseMGxgqOeFvIwLt7mqPXd+ofqb7MnXTT1Yxf9ohjtDoKIxTzs5sckaWCnhTBrz9xWC
TCjKUYkyaw6CYkwHTgFYuF0oiMH2djoR0pqYzdt2ZCRYiIbYo0Ptv1eTm7DsaLFL25X31RsBHZQR
dEt7qFOvf12X66Q2Td8XZ/8uk9+tJbJhgecGNgYhvTtXcMlXeQ7QDJtcSAWdVPKk9hfgFgdcjc8y
S4MBeJRQ0GyKqki+OwWEqMhICuJYnIRXs8KzkWIVip+viCcTe10gU874qNvjWpf4aKl0QhK3tPNg
PYwP0YNK+FDpr46MZMBm4A9BDb8KfntWhjIOoguxaPBKfHlhNgUmC9Fr9SIrSqVQTcv3zLBUdjW+
M/Iq0mWW3cR70QsGzg5dBInZxVBbuYxm4LUrhGgcAms+VWO5kQHIL7jdIrmmSYdPskIyqsuta27w
ixY/BVOa3831XZ1ncnwcwGzoxRe/zHcBUTNwqSXYorTQjgkafCgQqFtNX3dshpUmhPjw0Qx0y0ix
T8dXUf6DSPr11xw2mcNc2Qg/KbWi+d/AitnjTWO91ryF3zp2piKIIM4QPsZv2wK3QW4m24KfSr13
2zmqiUr+PaPgi4Jt/Rz94VRPJDTvLO5+wlQbtBLcqLcScNBMYX2GuD1tSazvIo31SI+G6rK9fPHz
UpBgNxZFf9TBCxdoq/SSK4hl0Ct3EuU9FwOOFvRMRL4iLxo1qRj+0M4yfNJ3OlZR9xNQkNJ1GPgR
VD9JzC9oswnEvvo7wek5ULBJtAshv4RzKcRZISTDq56Xe1S+8vUhhjoQT70rnKG11M6y/Vq+eTWr
EpEEBr8Oh/pcdj0JTThQ7jFPfjr7HN+4ueouIJDoG3olxclbOEELsXH6xEP8cNAG5oYryQvqQOap
UTw6mhIb8PciINJq08khQU8f0l5zUPJp19AVo7d2vwUw5VezvG5KjCsYNk7bIkasVju/f30ShoGt
zKY0CovpFwAFHKJXE/9Dkq97WlP4+RhcQnB7pVxbwd5V7Hgeyu7dMbLc/s0vA22brXt3HkzS6uxk
8xXBBojPJsGEamwmx4m4Cdy4N4c2zMFkuADNFoL6kgP/YUFVFAolGbr3laZEronArfc1KcWkzCvZ
xN5DJ0wZnsYc6fu5HzAbdjlCaPE1iDIi8HhjijsEbduvxWsMI9rwaG1m91hIisqY1En/WZ6G4oh9
d+XTalMS1yx3sxPXqqYGFsxoS6Rn6YjyBg1J2mVLhmZxyzQTB/gO+IQlmktji12/CAtb+bu03kHM
W2JT8sPW+FuE7hMBbLW0sQRWwkW7LFeQO1AeaJ5myoB+oIjf6lep5fNsHdG7W5cMMa6p7gviJWNi
wxoF0qkiQkBSHnfKuvauYJvbUEsupgVGsLArY62Krs9zQU7KiUY0GDKQLm6hgI8GT3z7uQA+hzox
/sm1kBP11jIXp7eh8XEpu5AfOxzK3RJ/jZpi/Mqwjzhq0LxLBQ2c0Hxh4L3uWBwbQBKUFndqYDPY
kyIH6av3wORUiSToTmLI7z13EEUx5FlyfUOkSwoe6iE0QCpHZNmkSA2E2Zt3BMUNriEgXYEgfUgl
ioo7UaDdF2T0GHtsoNN5G9ISzq2C+e/fwduUoou/aPJJQD/fixNI8gArAcjw99PAYxZAXKltHSTL
N0DqXY9E12T7vGclQ7XT45jV2b44mN70h4vzFwpNIzFFeJCDOS6d9zm5UEPgu6iyjeFsLzkI0SXM
wQ6xX4voSbaARHR73HbH2OtJco87+q4Mjv7RrM/RKw5MnXY9MjpfiD/vT5BmpaIbL73E1DuZWrBp
tUwSnvFqR85O1A8NxA6T3xQQxXhxg8zwb/JlNsTnaSyBapVn7tqr/Ds6saoN6JJsVNSleL9n38Ex
zjYXt46Kt3oJoxeUwG8d2GZXtA2fszwKMhiG4HrT5bpuAv3iBLGgPr0B4cD4e8RHbgDwf+Cw4oU0
+lklPpGESauI2QyMkeZwCMwPLNRv8evanGpLieOltv6KHsb8P/pCaG+lBEj5YPfwO3rr6tH697R5
ktknIqMoiluMqdtRrSc+VmTF2Zug5obemiX3qpNs7TtUTI1XebmuPlQ4tUS5DbFHp3M56nbFwcsu
WT3YB/7+zjUMwf3Xjq87FH+mLiPFLlXZa+e/XeS1ZCuNOiRly6IRcbFuFQctOtA4OwqqRTAoYI4U
CTXDY1TlL5f4+AeSS+1AfWZQNZG8LT27SGf+v9uh/1uT/9eKsHY0NEeMeoDxq4kdCJXuIZUrd/hW
h9voFlgLYwPCWv7bmIf1XJF9/Bk5TmF6uEjaOJBz+ccFOYyO0rYCxDibsoJNI4IXeF307dDmkyEZ
vUrT3UAwqJl60kKSqhVHIxaIQQBXcJa9EZwXZtaGxdbmIQKs+oA+ut35u066MD86herXrZkLSAyb
U7p4SgChFIe9CCM1OjbIAdNNs2Qe7W75MT1+B/rdBs6KbdEzg4EZNv/ONn94OkJ9l6MwdLX90Hki
FgUDQQwujJodRE6pggs/ky47GA/Ddj8cPMbXWlsHc5ooxhJjfVChQL0JAyMdevRShMT6O2cUwbWi
x6D25HSyKidmuEfZ3JbBFvTXhssDYHSHP4NKCvXMc7+HAcpJAJaNiIdCquyXBA5oRdcDOPdnz4VI
TAmyECc4Orhwj4HjdYcO1rt1gl1xsBoYxXDLrL848T1v805u1/9HVoRNU66JAu+wVR9VEnsa2Xt/
BH7X8jW+ONyZ1zIO+4rrpQ8TQsIIx/0FrIzZAsZn8kzJiKNivX1t52qMGVqYppM7LI7NVz+ljiTR
qd+wfCJiKIiiIa/Kj2qbMCyEplPH/tBC8f8GhIlUSOkg2OHx6Jy/4fQVJ1MjXu6hFGhsbeU0Okv+
Uncm+dsiwS8HqGKIaBS7Rib6W1V1OXUN07o8Mm2WjSWLStZahCLHMycWkcajiLGBJ1S5OX6GbwDS
Gn5EpoVIh8luFmWo3qtVrPH9mYnNfZre3Dczfdvu2iSzJgvmcCCIJZTVj3R6woJZP1IlZ6v4W7k1
mkVwp0BuVn9Vw3qd39Xu5ZG7DNy7sxcKx3hgkgbI1j8ecGTN9jXqSzjHOkL/YUTPKmZEU/FbXx0r
rpk1i6pvt3Zrg2NRWe9xTErjxoMXn/P1GwfC2GTODjmPhTHD0ocTJBpTMfQ8D4BNIPIMISNT0WJc
DYH+6wOsWc7CBISii6F7FlNthwpTZ1Th3Ue7VaYu132oUZF/+SAr2dEJJJYxY1t8PuvBbKcEPwxI
gXCM7gJYkBp36q+dtB4WYcTfHI7isuk7hHmEquX70lJ33PWbsGtwTvM8dNeCUnqOh7poiyw7d3PK
ToI5dFDuOKLhDsI1KiYbOAkfsGGZ6Ixhq+xmMXFzO33MdLsLyU/ZeHSCWvMOODBOiR+gfFNKuGod
kCGlE2fTph+oas//Kei2eXLw4DyMurWmBpsg0CNwb3mOOsIZ1XLsQKnsQh20TIZivnTg9VjATA2m
/OMBpMeqQNbpVTQtFNi28Lvz62sLzOcL11zWngrLili3w4fsflso15fgUkJQ30ilI8uFV5W6YEVv
WCZBEvuHgtqcRxctbT+3leynt4IGK3WoX4POCrh97q8Couz36QiRwk+1/JWLjN8tC910l3ySbk39
bWv3zcPMCF7lSN047t1DMl9yutlJmiBxT7hMTBxM/HPkuQLuJ5wlKQtshbGkuQNdrEWJm7AzRgdx
GVo7rANhvpWYd0/g8bmQzjCbxj/dB1lwUDbXhVQObnQqM1BXstfIIHL7XNHGjP7jhkzJv7+TTM6p
wRUIcyPfNdFMd1kxd8B/W3yzLrBBzvNoJUD2fJ5uMeuJkCRYGtb1v9G25LSoyAJO8BSZrZCl/46A
NbXrup5LxV2TIq0YpdpBuG6a2QF7kwjJNpJWOnRiCu43F4SYy71bA/DjASG6dOJ7Tja4yw4iDy2f
/uPnNMwstxTdjnB+Dzw3lvBH1NQYgmrdlEvqTq/GY70ruyIxfoKs5BJE2EyihJWqdv87paAlWhR5
93gHOh5x3rBtr0Sr9JahVmYrz0mG8mT58avcTVBZ3MVKzbg5xtoTx0enK3KCEOmKvjwimBEucyYc
orpMnO9JGKb6idozHHcS2Fl7sTm7cLvkvHL3XL6+gGbJ2gGYH6oElrxlh+31chgZzMmVW2w2NUSy
ex++GZ99h6ezmmLf8VTVBzixg6WlQreE9VNRKrJlLzxitsL2tvvilIJYECocJoo0KQ/coc4fryq4
LcpRQAxNvCufY85iRgmB52gxBBSXHwax3RCqaiwx087QGqeteSOA0mfmodYkAylDO0QCAJgZ87iy
qbi5Gz1zr6Buy9VXu79gwXypLNtXU4OhKlR3zAVRZasY7oGN2kVPFBjUgx0GrUsP0bFpUIPrTGSl
2OyaSbSNBYHE6oeiaIrFXObcMRs7KhmB/eQFRdjjr5FArTJEIg8Stl97UtTZl3Q9Q/UxwOrtUGK9
IIZOlqu/rXIdBcsKzldc3fdUBWN7QIAPyRDpYKEysqFJZImOjHjuPEiDn3gg5ovQfbED7VCwiSrd
DcvHNJXd8ko7U8QfeRP2R5RljkXI6KHRLicPhPS/PnBe+6dPY+NKwa5b8vQ5Di8JS3DErS09AKp7
KIfoyYt2aUe9SkRKOOZ6BYGrK5DEnnuDOvdFa5OFIa3/lvPJmqJ4XM365To8eg10lkc2utwymjIm
IR4QlC9GmOlFTDYIY1BBcCG8f/G1qbmdBEjzxcwou6ILNEOkeFFMd9ft3cdP/aCYLYNgsbeQG66s
ga2VS/XBgrwejcjJVID2Z7kPNpxPvqwC6sBOua/czVrglv13AwJWcHYBt/8nB/6611l0/rlWOCK5
pEkioForYJWzdT+pKfqiCGleRV/xQS3kW2eT2Xot7JGlUlKR2haQsQwGIlRJiKGDepop+Ww6XcFz
FOBatjdETNFyYP1oxisjxFRDmpmDEaUbWe0LEl+/X+qrK9kVIp/g+HJtfgrs2gxWNuxOBXCPZdyd
1V0sYxYoXh4cFA/p9Kg9AjWOeF7n/5NccZbMKbj2/tV9RPzsHX94KI5fWcBM8Jn2Kulxj9sNYt30
Fzu7Hr0Ekjdad3RL2S9K34vHQUa+SXztXypungZY1J5y8faKPvs5dnjvaf5Jl4ZB3Ljz4eqRDMNK
KZE2V/b2gZ8AjXM+sfGrPO5dCs3QHXI/YusVVZJhYxdONoa5ko9b5gYurDQcz1CJnw1J1OksNc8x
2jTdxkUsdIS9pkuWGXWj9nMpnvETis1pDCdGUNuglIBrg/jdgvuatNC6jkvy0+z0FloYGIKeJWlW
csC6E4asCyL0oM7y1/g47LYkNa+hDnkvCvbrR44h83N59KWtaTfmGD9HgGTyiAMMDLIIyDtOBPIo
FOqAspxzzGK+eAVNsKE+EjCK5LK6URNV964XrK7f6CI8qSEYvKbSaI+qqIXvkddxy28pEVN66kqq
x7u4RZNqg1bpFA6XXEtYxm3r+M46HHpkhFOT47DE3moDqsqzH0lJRMy67OdoXQHEkBYHUHklyiAs
J0G3GtGEnnYgzL4TgVbqac+84vMIjf0OPpOhE6P2EtSyjJZ+KrWbDzqcsKu/hzDyGsM6Q8Hg7QDs
28mkb0O8ROgERhIFFG0eoayuTAaNnSi/0g9UDwosH3LSEj2ZaoRnYAR3qP6gGYJElPB1E/IhyFgd
Bdg/sqo3sM9gfQL+Mdzh+P3gxQ/dGM3GRM53zJnrPN51+iGyk+wpRABQ10gRYNOv+epuwi4JXA8a
rJ12NSErKxKz6dDE+tXjwlHbZclBX/2jgYzqB7/8eUKJtEaYQdCm5V4mkXwf/TdrVuEq5eM70d1T
adtWFFBM4yFBrUQ65fuzHlDzQOh8FO6XkkOHOzbybIHIeRL1hfOUAvb31i8ogzm6Hrwkn1H2DrNF
m4MAM3RGUc3cMKgIbFuLPyGf/7xWKI4+Vk0QYwDy4eicUI5OsdLqkygTA32/OeHrDR5efWCplbx8
Q78GowC+VUUw+P8zFIk0rR9OWa4PiYtizVJyBiyGo8tPnv2oWI7ZlrdfGhffSIKUPW1wvt0KZBCg
bNjG+5NaZo24EP7CnPyfojIymfSO99xDiGkj/RbEBm8mTPGDPkxQdrQ4UMr3Q4JyF3v/Gh39h8KR
F2m8qvhmZ4t7PBElilensL03gCDErRLHUg1oP9xjHX1msRuR4mNvlqPsc2X68jetGYGarY0oQQVM
GDFbnEbUCsY/XpYuVXv5hhYdL9vGm5Glljm7wGm7KNbvZtiqk6Udt025dREQFPHJuz96QKVZABMX
licKzZ0zuv1Oct1YxriEvbiPfOaevSnGOjmANZj5Chu0oTGBgB1g28ciZcCh5WLikkSxOEi8V1tn
30HwU/DSYkM+l4zU5yduLZv+I6aWNkBgxXyScBeNMsKi5GjI75bSLOlI8CWMobXDLvTdDCq+9hUI
LVGZaxXVsG//4u5s774tFG8BQBHD0y/7UJQw0Y/rnGzENXoV1gpCopKZLZCX++VDgyAbTLb8W72W
M/BH3PzPii+Q6dBUMUvN37oSj6QGTfscbrHSCiLX0m+m9T6bUQTV11bPoOZ271pWDZkruojRWL23
/PEiWPo1z4GeGDlMdtEvRQMAK4C9JnwD4uww14NMIZY/qzVSlRSkTTACsd56csOvimGXXtgBY3WD
KpY4A0HPyGet2/YaaJ7x5enMHVumMZh65uTIx126MhIFndLDXrKk0t77Yap9+/z8AaqIWoMdYKL9
4+nsRA5J4qyLUQ1wgBMX1W8LXw4qAjd0sTtxroZ+9XQOC8BcGy20Prz9us3mGqavzccprLQSHN9Y
2Xn6E//Abr5qZPSAm0SXJnnwtCo7osMXhEQlnnnyW3LlNTGF9xV0NPraZFlX/TyYHNqtLAGCbdYb
B4Qt5q6cbaWd/ViwKl8QeHAZDVE7rXpBBrQEcCR6I8fst6+/Gwg2u9eilroX0gW/EMbax3I8QDnZ
CtyYNauEZFK3YaN8sFLB7d8G8/glZdc5G7JIxmOgato+fYDEX44hkDGeqXUyDmCO6bfyYZA0tgml
eIdx60uaJJYnvspg8PsUecWOXOJNeOpKmRRNqQJx0Sj82PtuHtiKTWZgBeQBnJ7QZ+ND2T0BtW+x
OY7KADFtkqCN8GYioTE+J/Qlb6akVzPgJceFXieleVKvTgdyxiGXU+AqxRupkjU7dub3h5eVutuO
FLR/9IVm6y7hOPNEb4G509bpS6e0ywNIEk5gepSIQycOPw43CNxXE+Fxssi+GCMljK35QAVFsYip
qLyLw448/nj/e7Wc3/0xXQT+J1esrwMdGfBD6eFfSyz3uXPDqJlNBfB7hwLjx0VuwtIXfAhLPzUA
kxTNlKARZy7tDOjRkwWi/B9T2tB/O5SfaxsnbrQUpFj7uNTrQujo7jbBDwmy4RjKrlb/kbQwEepq
ZijrKVu4QzgK2l5Hax8ZQTNRIfc/u2ordAaJHOUq8g+GSHqDD3tuZkZpWap80sAw8lhu7bmm+Efr
l80KFk6+JpLerfQsidNqOx2Xk/A/WJN05iwxYI93LCCUqqDWbcoDRF4PxMLWbNnAzzmky08C+AMW
Vm4h1rM4srqeL4nexiSGIkcrerhNtE7FmZ8nas1ZGiB1gZF3j0lJvuTj9qEIjes0snipnp5X6oh9
lVHqsSzp5edo7YLBulKvPeJmNnyAMgvTUJQbPO47HZvQ4wVe233lUUZnMgCPlLqE1sIen+hI9Zh/
HDGTUhy1JeJLKhVNM0laCaf/ytrTQWdvwwWMEsQpTkQ7+ogBfh8Ly3eAXBE6sgkpMRXlqy4coJqm
cAWBkpROuE7g9cJFQOpMeEx+eDdKF03dMORxrSuWFNnWxzUd86xz5Q/MCzXvoR7nwR2FkoXxxdXQ
cXj4N61ZhepVDBePlkBpgtoQV7sktaNEXcxgKRSSTqDMt3WNsqjeT5XpWeMOY0pZn/hzxEhd6iW9
PO7nMMaD21+cmpaPGpU5AleNMB+QeEojayT5G+PhjyKtkEQzZOR/FNmC4kdDliMBi7oDtojXgtbg
aB9DPba9wHRGEaYTf9uKyOXr8wjRl3uWOPpck8ScuyDoxQu+2TVYAafs9Sd8slqpd9Va9rPYj5vf
5ZyIQ8F+LLzvm7AhvaYNXtCAU/ZeEnMMN2TrXx6zIS0tVJKM8XBrO4tmXXCwWTkDwS2juu9i/sK0
8oDkSPBz9MPw2LXS1SLz74guadAxQ3PeNvNbFoZ4jSaFLi2cQ2k5+PCh2p0W3jOZRG6oCUd6+z9g
Sh0HxH0m2ro43ACZ2Z5xhD3e/gf39afI+/Ca6A7JrwF5egMvUUC29JqoK1Z5oEmyZU8RRF5c8mnb
6x27zefXloS/1jMirS0ZBUhzGuE09j6EPIAyPcGWvyRG4sSPEAjz1qgTxlPwF4OBGU6ASNU/D/6B
kQZoc7CSpgQ7KEXe/WCx0akaQLxfyfWpehAQnJb6k/ghcHOJ5zbBRoCUFcH2Wqii/hk9gn9Sd7/8
3izjrzATElyZl+7xSyL882LyBIUQPKNpMajT/ULbXcV0v9J2CI/fkfZ1ar6o5hNaczdlxTKNHB4a
7Sp3sQWdLKUJUiHOXOoCIIqpiiZiuMtCWnvgHCrWPM3LLkd8W0TKSU941DI2yjTKN8NmbGjndWaT
O+LLww==
`protect end_protected

