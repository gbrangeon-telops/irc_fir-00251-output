

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
q/LTCQu22IewzFL2xoALv0V8R0cS+n3ZGOXTlz6zO0tHpf0bhYU3nG7YhbNw5H8bMFnHmKPTo6eG
UeGsZXmzfA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RYLOlBm3BPRhwpOnNgJH4Vt0qZdXkt6+qKeUVOFaD4rlCQUegbI8dSeedwyfmRhRBYYfcasAbBQY
SHt4NDprJvJn/h7vAd6X1UjRiIi8OF1s+lR2yqR+Y5n/Ai+CRx+BajVy1wGHxdjiCnM87Cq2Hq6s
UytlPbN46pRkluJe6NI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5Onxh89dWZfdY8AMW/MOzaZUaP+doVdup9B0riUkkwljU4WHOna1/K734H9kkMqSDTQ9ivkZIsmH
DErXjPeoJcAWqHloB9UX56vG6J+JtHhxXpnFa4rDUsDzFadXGZZrXqt/NJt/7/nP2AP1p1qeKRkq
ksYRHunueBYG/B5LuPR00cTpoZaaCYuJroh/pzkerIy/CPNX1RAKt047HCKtvFBXH7wuqo/yaUyk
Xkrxw2AQ0ggYgz1hK0KOdWT2JckcbGgVwPsik+mchcvmPUBKx8qFAnef+ZSGsUTy+3gjDznrQOsF
sJM7rKdsAjU5OLq3k8BWR36ur9hbMdk+lvFEHA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fe81XuZ9RrG7wwwI46b8GZQ5C9RFsRlLr0EzhGvkV3ZMeUUoQPwYfJl6GHoj+GDA9GnY0KeJe84A
xt/fhvb4h1DNhpVnvsOo41gu13r2msE3kvHyK8en6IodL/Mdh8CmalY/a7ZhDb0W+KP7rEAgisED
MHKHkmm4OWbTY9lIJCQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JHuY2RJ1GBIZ6g9aWOE7BqrGN8uQypqLnY0uHGFvCX6msmuceGWWswz4xbJBwz2/gb4ZfVDTzfAB
RXiuZlDm1B8txxWQYaxO0lZYlxtzCU/lUn47fRBxEhyn9Yc5lQx2oW3B/G9c81S8zCONQlmapnrX
y4OR/jDZXLz2wxMs0tkWUSXHisAbuRctLOTsTUfqMDUsJS1g+TDQCDpUDXL43sWg1LCRd7wDn0um
3q29OwHxtysopGOz0DxmTcK07ZEEnSJS89piniLxLQC53j2zOhAk7sCb4iRKccCVkkeasTjlcMTi
rJCab5WZRXi1gu1yWZ5s8tCfrKbGVSZTS8p+pg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57216)
`protect data_block
2Z8ZLgIEEeNcuvjtu8y29BZR8NPx6LZwNxw3UyZcg4M6SPVL0P0RT1jgMm6+OA5Is6RpR2GSwnHB
rLTOe9fGWu80YdWTraTS2jXeqElYrVTdhGJP0GTX+KPXz8zm0OHr5ci0FZSuOWYYjFrlceinPyDS
BkzMtDm9W2GMXdOvPZ+fSmOFjXLBDYfcntpk/djL/er5NcuyVpAc/yFd09PpEBq0aKVpCj9aSkLE
vYlSv4QknLlBJuzf0rx5wPZi+QUDZwx8YX+ZWzGbDnk9khATKcLLRTOp5R3fShXW0wEjsjnw/STd
KSkKkm+azLzYgDE6YlkPXprTLKzgU/lV8huGbt1cruzXNV6kKPgHhH9jG75GAQ2eD303eHBmb59N
WObIs7jNIApyUong4EaPsKb33L9ddo94h/Yw7HuxLwmaLh260hZzTCjDyZ7zwMu0qY9ds8cQvUEp
vReOMiNW5pizsS16raURUIBOxoGeOEw3rfBK3G8v2UuVT5kwHLFW6y2T4Gaf3E/CZWlcX/URcc7G
sDFJnLLoLUm9I4J2tEJNkqo67a9oROM8f5ClpSG9Yir4yHqbI/L4BJBsbZdLa4zsLmMFHLXQMg3F
LJf+6q8d7Nzdjs5E6f2Hdg+uwDHFTaVOcu60Zx6ANCUkDrivbu4UVwhclfESxOeRzkKhSrjjwFtm
1utRXW1oPSEo34VwS2jORHvLIyfQX6aCLpyIAo+iFJFnIWOdDUnVFEmu60+vyCJwh655M+Gcz6cI
aIbZx0KLs0Ml3Y9KD4PQNimzsLDdmR0TflD84baLf9evVSZEHTrKk59C/H/lybNZw/61XLbB1MY3
KUPJ/omehOos/AUl1Ykpo3hKC7Y0fGUCuzyYBOBw6YmxGq9NZN3rfFC0bMraohIIOr5aQ/aBHFNj
Qwpwphhzq974GtFf3TJIwGuI8zTuDK2x3MNZHCw/dCeqm/2mw/+zvQhgvNnheId7/8xWlP+yvLbD
uPtHX8CpEAaLjoOaVOG5o6KPKRLIHoZi3V+n9yfpvrOpBtvGGgR06vaCzhx5TdQzO0T3qDhy8JWy
dJ/gLVcuws+2R4iD3Z2+C7YCnjhGPaz3+m9AXfWuoaSVoujERWY3zbduj97Vbz4q/X2kC9yikfun
CDZbrpgQmIu+vfQ/V5yupiHq0cHibMhWcbmzn6MDauV6lC1j4ALyewniGymIUU4AEoljgRspX6oD
Ccb9PVNl+vLhVH3SJrb09IlBzYHLOgaZj3dsX+yj9YGEFxx7QSxe0V0d2CQmTwzv4wNim6gEEIJx
PsWhZjyJEMV1BjV3cBTP6wu4ktvGsh4liVnBas32l6qWab224S4J9JgmQ9PyjwlG60UCeUlbkRmu
RGhTIoZkuglTczvnnegH4lIS1elXKerL8B8HsL/yTowqmN5Iu0LrmIe1LR6F5SGTzmzO2chqYytM
40zaizpFct1X8+SPXY5EvOG1CL+wDRlq9gafafoUi4kxXXrAwWL0mga4maBgjlgJDQJbtKYhzVnD
NFEoV966oi9qFVzi0WEEPnNKL8WQIHvg8BdU0qVQbj5GTevWeuF5OrvuNxd715FkW+jICN+sJk1h
YhzmolZaLB8ZflkAAJKbIKSqRDTBSVkCVyhDlmEI2rjvWwfOhJAaSliujpi93E+QkWuIlu1QhRit
P/LdU0+FoArfsFvTwObGWKC9aOLEOYBHUVswyc4sPVgSLXKhQ+BSsdvkVh3Z3su6ALytmQKLGaIG
sBdB/ZtvZbXilJqb45UfHrugnEzypWCd/iyTRWYCSWGPqlACGOGQKJBeSsTRmPmnDVmwERIIXYo1
9KT/tabKQmoj7SFf4kwz5n2rr2GpWg5ljOW+826Vz9rf1G00LgtGl25MY7HFSIxBr6OEteMjz4yT
TPU17mHJXjNjn9zHSr2BBhL44WQ3AsLU4GdARE2kbTMi23XMbBZJ0FXcG4AbLIuTs0SJIYRa3Oew
4NDJDNXvFxTuika6ZN+BZsLqwS10umXePrfKkg2hbdQ6coRZVwBh0j7yNqpH7tcnmE44/DivPz/h
sp6NIC+dMs1shBIU7lrkvwzTqWcQD44PB0VrrUCb/T2m/hu/IJ2K7YoStlkXysUKBBH5ojFG8uHX
G2kkDtgZ7v8E16V4kqBE5ZffkXrvTxu+DrY/MLI7BuLkpgGvIHu2CGtHfYR0Xh9nLO0U8CdS+LXU
nwfox8XNOQf05PTLKp69TQxaXDg4sIl/yBk2ggk9eYivuoGMIJRpUf66/VY/pr4ipq1JIAwB4nLW
9vW1Jo7cfF7QSFaCUSjWYSoCUVGx1AfQKuhDdpC/IW3a/N8U8V72MPeqEoh1VA2Mnzu2XNRDhC5B
p5WwC1v2fEYCvOSFq/KYx8ZkwM8g1diKprX4KJBrrhzxLroO44poEtm7ASLS33qA4I/IGtcp11ev
Y2hOgDp5pB7bNqMNmif5cFCQFXFLTOsXi969qQHl+2yP5zB39DCXmh4OVUc9jbkqinj1II/KcJlG
29C9iGfYgMt3KuTbFvzhuVGUNaOFdXG0S253jDn7w8jLOdTTXQ18wpiPY1kaN7jMtbahxvsUkE+d
NDtkI/7IV9Tnp8YtwTIdQJaLfTWxaVkaqWzoorW/KYWLWUXRMCtkmL5TixXg45ef+vkON4hL64+I
nhycU74jQBiEqfM8rFOsY6CoNqUIcHI4NdFMi03/Xe2GZP+vTYxrK0Yc0s3CLujFj816wYOy2Eko
ZZt934nYaIDh/rPPvn02W7k8zQaPlsjn1vg22NcXyVEncgt0EA7CNgf3q/PeD34q4S2IYYgzIcmK
it6KalCBgzfvJ8oWLVd0/ZraTp6+q4pN8OEZjCgoFhrt5BkT+yXfU/nkJCqP2D0hjIM1meGzOdj8
g9rohdBcxn3G6lN6VQ9F80ruLU6gq7T3CIKcfl1DUWcfWPoTkIF74CyLrdHG4GTm6/PbD+Nx9Rt7
/AzwkLtIHCEX26r/qRwhy7fv7LC54N94+OYO8gzoyictyfMnsc/gbnnyWQa26heDxsLNDCteJc8f
iVJQM6snBmjzvKDrmVZ7frS9qGwbkB5lNkAOpzCoZZjFHZ2TE3i3dhNKQNmF6Uwhfs0I6SMTPurc
y2Aeunil9KoT5kmrwKYWWrue01quguWK8wKMKbvc9UOn8xkiYuy+bVXZO1G8WAYC4exbYIoDTp4h
KGza/QxNC9Y6kTMSwlO6iBAdNEcOjpGSB3eP1WLdplOAju3pxHULFmYKKnBkgK9p2didKf26sTep
t4C+mxji2Csstv7gI1U8ygHAHALOthyeHDgh2Vo1vFXOE7mYmo1wjKMzrNjno5FRr5RFz+85MiDg
/F3X0JNrYExEInfL6Us1jJ9yXTL+KivTIXNlU9zkVIL89r/NUr7iUqUUOKJsCHOCmxGoMxzQrPaO
U8ADYE1LHSggVfRTb4QAbCC2emwhOxRf6rfkyL/QeKD41fWiGZ0l4zWcQP2K9c1uYembPweVcIc1
+1ylZ00fLd8db4ht9WOiqB2bXPrf+04cMfP00MfgoHqhGnlQHHZozZWfCjFfGq8gUt3+wZyLC6+U
op0BIB+R0oiZQXW+39MXmn+17JUHuBO84hGfe/+7VOOC6PgefNMtcoPgaS04imzBMQDFlrqQON/A
gnNssde5cwHVLX4TtmKt9HZkL61NLzGmgg5DPPN0gIU3CkXtCggogGCKSQWkSkdUi8aIWFxzEHZ0
CjtcARI2vFk6JtElo5zNYcD7zAZpcZx6FtnOSMBsN0bcrDlddZ8etdDHt8qrJFNgyM7kW8qgPLKN
AoEW0y/6WF4oxZYOqsnp15votPdMgVH1O8zgnV9K7MfMystdvFmlrmVbRluG8paGqt5fJipzdiDv
C5KPsOmkY9ubVg+LfBVOMoxFSXYHqNacX+NDewtAMk2Xrm9nHPH6YGrPfWFUUbKsYf0hXEeb84iT
gJ8XNrAXex98XyB1PS1Ppaq2Up6CQnN06av6/sMRPOxNa6T2HiDbbDf/3txQ7eHJJIG8m/ymXDKC
fAAqPKZPiqhVMprBpJ532V36OJTklkzPPK2NyUTZ9ylv1yXMWpdE5RzQbv6urDtvLnT9TNKavjwB
1kYbOApLKcmWvbesZC5/RNnMiPoLfN4Fb87RFD3hpJZRLNmYZkVidy75IPJcm0rrcCYrpM/E0HhN
PFAoER3h5lU+qAqqs8Wtxw6StYuWZc3xLbUApUS7b1mDjVhbUDvLhM1PAfyMrj7F0RJxCSwarAZM
x5kZpDruD0mccA8+E1i1Emy9SJU5Cxp7yV4To1qOa1Uynyu8wImqVZqraK75CjpAcCZhBdpE8ttY
NXbmWZAGkQ95hotmPfB37akj1Wa48oMqQ70W+y+NdI2lDn+Hp1WlXyD+eDN2N3Mc94TGvIbI+aq3
4rMGvFoOIKFZnV+ITYAj2HHIGRWFZKoSbEo4a4GQk4nqSYGnCjA9fVuuH6k4mh/GkXDTPty88kV5
XdNp6dvSH4MHYOrkd/xTk0zFrbraAP1ladSxml3NfexXbJICej/2KfOT3Ii8aa4ltcu7TL8VuPIW
tQ+2hhishLXVktZyD9FLCAcLwhgQg9zrClw0oh2lm70umPELtaS8d8bWjsHe+oF8l8b5IJves+gF
buHTLudaTZTLG79LQTWfKAZVnZ8bT/RswLOcL1/kvU9WKu+FmzlZh5BhIxJIBLlTtlhUQ8YTruL3
FS7t9+EmNJqblzs1Bs6TjrgbJHmNojQEA11Pply3apjkmx2q6co3jFO1mpXXOJ4MgtYfuTKdJSTs
ekdqCtPnjqW8Rm/JmvI/I2P8fyJlOHAPLwu/ebnxipEIaWDxizTnm9pksDtpN+ZP185jx0hkLSxW
4aT9PuCoT3OSdiRsHOZ4IOUIEdXYuUPidPNyWU8lCwAYuLXNzXwJPRZaW00EeqNc5/Pq8ZrbS4q+
j19i3Mb+/cLnASZK7Q7G7cK74eWgPT5LbXkibqz1oT3MmdFms+Hgez6Zu1ndkq+t686b2c4aN/YJ
3JQc1mZuy6VE/n66eVu3BNw4xBdvjNiIrMXPKBJFUXfSfpEdtbFWDTCQLVoZT2gdXL26N8YoiKZG
zsWZwhBauQSfJLQw4PzQ0freMr7f0eyqfBH+8+DqTFQDC2uoVuj2zNZ72hMW4y8/7qjzsKKG6A6J
8JmehgfisODpC0dzzQyWSeaVnlYzoMNHVxV5ZVT+rRbgrkG2AzoVGpiXUFDJjp0tyzZfXy5NgWse
90/Q2VDxB2J7ZV0EHzkoLkCv4ffNKYPXk6/FH+3qNO5boQg4L2vvrUr6D7oYeovwf+ABglKdJs8i
g/gb7lpSnjEDnCa6YrD+g9YMRVxTOANiTA+7+++IUnAB86IMBTSg2UPMY2Avh8QWCjQ0O4GEY28b
K4LTRfDsSEiz8F87FvNm3N6iLtkHfMXpDO5I+gFU86cZTzVDAdqVq/sVQW39f5QBo5m+LomLU5My
LSd4uG3MVFdwEZo/TBEOAG1Svtgkzjx8fSinCuj1BupDdKZRQXrxolY6kYOBbl3MP2GRJbGXfczz
fXp7g6rqGNW6xKusGgCZdAFlyD55pG//npxr0iiVBUZufKL9T3WsVKQjUH3rrK1aCWa21Aj6eWgC
egPbB+Fykek4hXPSSwXB2WUjvNrlc/dDFV+EuNHjIjX9m4VninkqZpl88iXLivpxkYvsOV29Squ+
yfR87tYfwZRWog/a+k8blfmnnVXiQA3I/9De6TrFQmXMB2g9FkNaFnZzS6JZlSP/WtwbcLAXtfSK
T3G2WUssJIVu0z+zrvKchxP3JUbIvvIvspoaDMN7NXWIdn+83Qa8F+RayusPsc3Otd+Udqw2XGtY
msVTQPTYi/hIftvcXW4R65MQYrNTc/FmKESpGMK3vIfJLwTtLqbzi+q2ed1ekCPkbOlhu7ImPdvt
YGE4vesmR5U6jz0JsgprM3Kuwe5eQhH5lO48T86aKuRrtSFdvlREuskdx8040MaLlTY99G38BXaK
4UC/jA3WONsPV5yHFQYlgI4Nsd15m6lROkbwcg3nPEpeQHnJKcm3dvO92FbSaaeelGrDbk2iSm0s
tPl57WVZtf2mQXr07RJD3DjKrWXRRx+IIeCHmXQujtXIK+gaqUb/3GoDQb1kbD/18ULxCYyJbxVq
vGeaNh2zNvMumHCprx8nKkCe47vSyP2v6x5FBrDyRbMzWMQIZyf6sLa/59bFc6Pn0jCxRtIDpFvh
HXaXEfQzuwcDc3FKLlIAHlZXKJecuvFjSrXBAHTni0o9JQhRRWVknSQZtkTrzsPGjJLCUd2ViiL6
J2vbH22fq7lOQJEWyPNIWae2jBNbs+gLjQHEeWvONxXpTJuPwZuN22OeP1ya5kBHT3emIThAoVot
npLgYzhxGo269+vjhyQk7OG5jdIp8FitbGg8INSFwjfthh3Id0Yr12gyT/0rIJsl3qO65BrezD54
8h+z41hLepvymogvbF6z/QnjS2dgtrg9rQPeXkciBy/L2hZ0t7xqj5OEQUHH9zv2VWyF0orMXfE8
SwKX7cR2oK3sjpkJO5o3scrtV1b5pzn4tuDaVKt4esQXTW+qwTQO0iG3+ln7fgLXkNH6o+DOKHmO
NbuUt0Cq03iX3EJAM0+502qsmZ2KNmts0kFXjyrltMc2xjEAh1OyB04PsAz2VcC2eOEzG/wCffRC
tcu3i8nsIuet/RpQ4geUKTW7aLVK8Yz+50Zt8toa8i751C0ixgncIScC7hDutIWZOiy2nIseFUyi
Hg1YWR/eukbg1G+ww/FusiBMw/JrStu2vOtYN+fk738/kVrftEejlBFk7A50NCaQmUxIEcITt3Ii
A68EY8f42+cXanx0uE3s0qjTws95CGwyLlskeT7MoPdVYxu6vBkkJUrgn92jE8poBCPN/UN4ylrW
xdEUpZ8cISkye2bAJJp0X/CL3FR6aupnzlHJKgHFamC3v+9t9IO0nXA2DGKg4FutOihnlGLjmcov
Zs/5UNI+xbkserKAoFAeRYLV1UfZwmFqMJekyMxNYGgDesVcdeyh7i71eVrHgeMEBAmQl+EDb4st
8wYTpnT7xzvvojihRKBrLq+ZsSBEJ6si5i2EhQh/cm6R/qJ/3oGPPiVQV/BQH7jld2wLOufotug4
M+xJFKqbuynxzZFNgB4Hsut7QE+txwFFco/aMfvhvYScQA+R0g4N5BZeCqysagB5lsskCyQgSdE/
oOITPuVBr7yQSRHphKrc0u28Smak7j49Lw4xHRMSJD7JNvJcPe9Iq5f7iojD05tLPozbGMozzd6m
ubuMrYDxjZvSsftgTtdzOH1bF1mAz/83J1mmREBof1nUzee4+lWffjBX4nNnBK1fkHrNLoPPhYKX
ZQozlCw7sLD4GGmeF6VJD50sAqBOojC9AKRst3hFcAvzXUP8NbRIb7MJ/Tuj1KC5cM24xzNJFKp2
I8VLCxT6ek6US176ynKArs7voosZZIPzFA4gyFAOeagExqvCpHb6vVsufCEXrBWwl1IQC0YRV/l8
Kx77h9d1IZIroimP+gAX0GGAdKjploAl43Bd63yNYmqcyNOSuZ+AvmM6pSZO5f/EAJzqe3+q3e3e
sXhbY9WjOf0gxTicU4sD2rQyJjy+K6HmqLHRdaaDtUl1ql5iLhj9wCzhbQZb1rRQDsfWHhH1CwWW
sCYUROSgCKYsRlu9Luc9tBWzgE11m+g9g2ZgEAh3RUuA1Mj9cpOSfwUvuqymUP7rJfIPVt11PRRq
rgn5mqmVB0gK629Kh4SiX6MzlhFm6o/RKqFagFxySA9XxvNTbOOG2X4yRN08vjO9JuJcxW03l82O
R5prT+M9CexH190/sV51sZ/DXldccQ5/z6Y7HeUEQWHjwjgfI4P9nl1Sz4enlizXdpZLzFPu5BUG
uon0jbm67ZI6okNylXhJXHL1wZEa4q78jgirw70P2xncX0bKBXTXro3rHMPW5xqHH4AC8ZBm7At8
4nPYGYmgjPqnXEgD9oVUGcH+7tmzmXRXxICaF49pCtslVSk6kLlz4fJ5NfckvA/J4amR39n4nEXk
2dV/6KFpXnqFasKCiIDNzr+lGrmTW9dM5dAf2z78s1enhmA6Iov7AnzdkoRJ/dJxhs8x9iyZNg/k
nZh1XAzT8Y6wNafN/QX0rDUcXpToWiIOXQtZS1AZ8DagOoxGwEGzVxXAzDcbMbGmRUAeF0CrSBfJ
qtGoliBq9KO5RJQ+ePkfrbOJnpbC9znfz0EknlRUpcOLPvOKIbMW51WYSDJiNZp1UoK4544EzMmE
0fsiA9xwpiAd7g5dLh4AmXSAeeOx0j4ghW7/QEi/jEXE6bBj5z4hIiayk34WypGReO+AoTeRvlLf
FQvueNfaBeoNS+NJ6rH0WEso63JLDLFlYpZH1k3276LL2BNl8MovOU6z4DFj61pAoaqY/ezo/MU5
qeIHdJSTXqJqgePvrCgevjN6JFLMhGOXLirmTIFzWkl5Rw7xuDCnrLqpfCdvaQou3wbd639RJR54
N7Og0fhJYg6YQw7tErvwMVCdPqHAX7giWWnrMbFgq/V+8Vpb4dMxvTDv44wG3UnvhIc12TyA6btQ
eJIGYJs/FlkXgj1hbMAfqybANpaZ7VWIPvGVIjqJBed41MN7UwqyrxSQnSv5MHPzyi3EdbZSH0FU
XtaEbPu712y7ri1lnYGC4ETia99lECc3oWi7LFGvwmSOjy0NZsXEIWw3BwuWdHAIq/FE5GMD4mas
UsrqAi8Rdmw+fEH9J+X7d2Q1jSvM22N+3dpVB3Bg/zGkoLQxUdbswDiGbE0H48uBbNySCP4z1UGC
5O2tA0ZqI5vzQCBV6k1OX+rCRNAdptheMsUqOM0CckMT9QdAzEVPggycmKspl8lA7gyJLEu8lJwY
gaKZmbWg4bVkmeXrTpDv3MqfThT6yeCI4EYuCupC2/kYzlEbmaFB9NmQUwMz/6FBPnh8i5P3zjML
IPFqOzQWcwMAcl7Yp3zOpjIYuLE4KFXPriJa1VSiBu88bZr7JltPnIU+gaA2nygUrgXyO/KS6lVy
WmGtNHWV0Jxk16QoW3fqLbK07wfpgARuoaaMAJXbUngq+LqsKk7FCVSGpWSOKA6oKEvhXIUXoNJd
CXXOSM5L2IMsgly7ihaskO2saAHcdtpUL8MIKFiwOBaQu0y1ihWGfp5SMmTVrm2a9Ru5gk+Jv28o
2Ajjf1Tlr85xo6cTNNrfG0lXLQkIz4tMkK6PrKbI/Z7umUjaS3UPN28AV7Loany0wjUBRMoS4tYY
/MwwD6j0DzZ0WCDbE5oC2fvG5GH859jxGKXFGcpZcaZ7BgR5GqTQf+NjnXL1mI07n2ic6evFmtlk
gM/BSU5JRVayjULh6kWldObu3Bg+/7xkR57MPV7hpfV+4uqoCnMe+Hz8VB0QNsfi5dpaqT2MyKGU
hQyA/Ot0qsvHcCyeIjq3/iXlD/BzB0gdQxc9ge6kdgNQkZfWTl7ECWmbyG6P32Xrfua9zPoxGH4D
sS3VDV2ueafIirWwyqPp8UxVYCijCSjWB8EUcJQYuVPLHWpMrnvQwLdfTghovY8zWNfI7WEWI/iv
cu9QcFF2FH5CK08hj42C6YUGlY0j7DR/iLNlqNcmFwlJPNf0xBWPVHw0xhbBqFTpHzCyQGBbWXoD
CxT8CHqmntQaIorr6jBSVR9ayjiUxTSheoV6poNCdLX2XQH6njc3bjKhoZINIzE+wUdQyOswN6vW
Rb3fKu16t143AIyRTmHrLXkgJwfzRQ6UfCGcpJUHeh1ARaVmglneAURDgVUvjS9nqC2JQGZfSMAX
w53RqyTsT9P635IJJ9dgYdrhRIh1aE/L56eNT+J8QqHKysJNKb5+KR82YSEUI9KyLMDtSoPnLONh
QlDWAKJaqGI8fnSescdkGeDYVZUbKzzzJkpQKXKUY9xEG4l3Dy/d5o2Ow8I+KFVFi/tlsRVeJ/IL
geV+fbCnXhHSl2MNN17t8tOFBLH8wDOxUZ02Gu0nPCMOOm1Ux1Mv01QhxXR0aC/U4BpmgHWYkWwY
jv3eGgi77G9SxG8TJQ5hCBjwyjI1AvcWNeEY5l28e0VSFnvSpzP57CxOLtsYNsGsZLkapcs2g27g
vxbkGRNvdyhX3SleH/ClHooRBmLdjOUnBShb9C4V4GR/wGrjsZCR4xpsWun04m1sg2JfcsCZtTlr
7QWE56TTHyLJ8zuBtZzq2zqpGjdSWGHTMaIN8fPRL2GkFHprHet1MOg9304jWX+MwRw1EU86LjW2
hERQStjbIFZ0AvfL0KzKEQDlWsj2MpgRkdy/bsG/483GxLH5BRhsCXO0cCWM2x/pQ0hbHPT/PQdh
AD3kbrz26fLESlvJUcXyq1L/FwTw/j/l6V+RGT+Ehu4z43BTmfaY0LTo1ZOF6swrBVaw46VAJyad
7CiR0++RmJz3Zcbv3ly6EIk1PBUfLMDkRXv29j3h/Nz4aTyvkZr8Y0H3cuc30FTkxOaBUB6k/p+J
1d5ZBlD1mOlBeeh1OzLNguWhmm3YYn2WO50Lk9opCfSpQ9m9poUPPPoLfEhBWMNmQvcG5065Q8YD
uCck/zeJjXs675DOaMqYwqwok8UrQkHvhkgzQsq7tgL08W6zxx54XBDwlBQYo08qAuBS2sXTEUBO
A+ARnQwsBSXgBUeTMMozsX3UyT3FTP74mAv+ibLXyiYU4/Avp+5Pbv0GnEVJjHvOanXSD+IcXwVZ
zfzxRryCRUGM2SoNj+fEXKxls7Wm2mcAEjeyXgwpFCRva4k25VVV1LcH4dnhJA2P3EQk6BKXq36+
TPWcAiAO7brpnJp4e+9jYHoczWVpoRF9yd3T35Vk3ac84ayeakrpiDca48sPjrPJnauwnelVrmld
gT7KLzIbF4VrBIQW53cranXf7pnO+68UjkZRTjXD2+AXWjxXu2e95w14UaI8W5jGtcgexioMf/a5
FcjoHcB4r9qM/cu7FveKItSz+U9OzGMRXNpo27Lf8NjDTjasELBn4T727s9nk9rfwlAN75+jnLkC
NT/LsWVWAmQguTEFQXgAaniL7tKvnT7kiJfvfalKtcBa6DDCITxoOI+PEpeH9lO2ewooiJ2RjQDu
neYwqoStsM7h9xPOeMj/NCwR4tMwjmnvo0I5TTU84VXGetgF2t1xgIjTBx79L7qeANv9LVU/FPrB
kDN2PU33ve4n7sof5nkTe8wKfx5ToAXSueHNd8pf33FPPPxe/7T0cNRjE1/7Oq5cF3dT6ye7U05p
mhKtuLLkKAoYiQtn1TlaGHlKOEzNtUJFUXO5lX6vnQmBXmsj40JV9+ww3f+UkzPFUh1B3qhwmUdW
l7id/aSlwgD2kZd1qKFO6Nofbaz0QzIJhU6HYxIMOTR/TwlNSoPpbNSZoXYiOgzfEb1mH21CkGDX
8bBiZvqzWtFCP/229g0nJMUyeSRrCE8TMRvG0E9N2KnmvHOYmfkRPetiKVX9YKV3WCsxXOdmag8S
+DT0T7WKfi6exopmBswel3rEYJ1SYgXrMcpkzve5gOa06Px69tTnzMk9LEL/3z+T3EuzlZ1bKeyv
k4UM/4FQ1ckVpNkmVK7KpLGoKX2PxGncV0ueP46chS+Rot766v2vWgXe7g2ugetGwslDmoytbPZd
vZYF57DsCCxCcmH703QZjmx97u5E5Vwvk84hPFJHtnxkExc6syOe4sWdxLA8Hjf1IERoUFzbe3ay
ZIevNfJGCouxQYiZ9RXJWAXe883WMnlgbH0KHmsSGC+CHNx+gt9lDGS3BxUIobpLVHHmQBgdjSCa
dTrVYyDLxOF+7yTWTbx7wEDEZF8czwJGQmLgGbqJhs5LxMNduxmBcwdPkUK5NOznejIMBSrh4MG4
ghAu4hxZm5q95dkeT9kcjqHsJdoOLWfxmAd5sBDlUL/WHtsfBoPTOFsFKmBefZGUSeDmwmPZ8Tfv
1F2ASKwOtsSEdAdaADrGlpPiMO2s4CGHwL2wd7oUQGAAQBP5RRQyMLXqJ3HHOSMtMB4WywusS2lo
P7xQcH/1/a+qxFdfqmadMSGXYnoxbBd/fm3TDItldWljSClCi66sST844x1M/PgWHEOJAzG+8MQC
9w0TLRx2i12+1PLPxAtRbbbtbtmeLLp4bCpO37hbQJF4jW0+hgWLBzFp15jxTjgFG5975UdeHQJl
+cj3Ys2hd297SzxOUorO8pFIGGwymtxPqVk0UwPcHa6sfH7gChgGp+V2KcJnva82wdENYMu9iJiG
E5vCSPtq2hDmnVLQL203GsmWGg7FQzridjndrQ0Fu14frqgmK9zpoYCzcgIqnYT7KoYFyE0bNpEG
3su6o2YvON6epvv8fb93KB9WxcW0302tguGcWr2S9ojZ6vA8tpUJi8OJpiVZFUUx1tbhC2ZE77CI
WaylNTIOZkDSPasVpxU7oqn1bZ2BPt3K0VsfRMq7WuOvrUqFqFsDa1MyApvzDQs/vvZZqvghOlQr
vDUsL0OnSnfxWP7SQG+xdoHEgxUaPfZRFNB0Vsh0Cv6OPARGkGqZHlW/ClYNAHvQBs8wdeHtXuKW
Sy8qRTuYJzwCqNpBL/5MQuHXm1y//NDjGuzjdx84meHxnvsv2Hti83dmEZCwPlivwFYDUKTMa3wE
3Qlhc7DZsVdZ+bE0PJ9JC7zg8KYVGUx4VCkVIWTQeQjOBw4M06dNX4m3PPHOvJFVe/0+kEpGK5k1
0YjVfA4wC5Y7cS7C1yKJH8xnJe5oXfSAmrmTGFD5ji7rU58IN6TNYJrQMdhDmJKKEFDlY3u5/+jJ
61ZMdMD+E6pR00mbQ68jevv42krq3l9e6WuJ0rWXtL0IUsziFepyGsMqotemb1kAhP78HJrFVI3A
BP1loEJbxxa2Ve/E4VSpmU9R5FsdminhqqjEXrUIeBQd3Ig6XSgqLR2AfYuWcZPGrTqboj6Gmgqj
7MkAXcm3/A5ppCcmjE0ofkYJXUIYVY9C3y/GlyJRvSzgQeirSxMo8/WmMY7qJXciScdyDudyVFb5
dDSOW5xOL0lLg2NAz043etuCII764Dt5vdIdWkRO2glVTZDO6FTcD/UsmecHhDA0qq+ocuFU8JnN
UhhNAmwQEaUxpmZUuxWd4FT8tmEQBZqcmPrTqXLyimJU+YnlljbVhLLzi55dPw6aQnVve3XKHExh
GWram3WrTqkIYsslgSJWJZQAfRr/lIj1vhf6iRFrNZ46GF5XldMmLWvhVAZwjs2l2QJ6JELMb0vk
n7AZlvpUILnM8uiJXxUYaVLsON96rqW/02M7fFYZLvPhessQxQmfae/AXxEpS1OGXHNBypAVk/GH
3QaPAU60O0wEeP9ETFMP9580gV3A1cJGRbvpiYno0kNkoz7ONScNHNL0zT/1ei5kbTo+pVb65BQK
lpXwAtwSmu7nVW/GoPQiYZQHkXI+uJZcrf0xO9sI6zpav7TqmaacccRgvQEiZ27trYagwMzDKV09
YHtldKo383CD7ggm1ZHXHYB9akTMDmL10+ooQafDo7yoUohsfM8d0NpIiHNkotF8q2x8P2aAKtpZ
V8YTh78fBxqJ9Ev4MwJLIx+0/OPItQnz76seTo0D1i02Wfnsa6EndOzicMDq5DkkV1TfzGo5v8uS
YgHZfrnh8YZQOIKBBjeCJosHcQW1B4J/XD6wBw2DO6bqjpyiwSRj5HJdoP2D8dXQSBR45x4GuizI
ExzOBGAAhDJj3fAOSK4oklBEvG1upqlrA/wGkL7jFl5RtRWdnQgxP2BqfgeC0giYrFq6qHc83Ll/
3yrDFvYSEXL4YEIiMqmqbZSKM4HWlpTId/VQUwbtSUcFK6F6yeeRyBH48ItDwYc5mi4T1Zf5PKtV
Dh1bf6gl+GFMt1UkkHGOk74s7nYvtLbs1gQnlLouNb9Kp8k0TLFYpSGUzQKzdWS0YlpR1HqqWMYH
2t0GUNbepjg3q2N1SL09pYhqMGdKSpdG6lSCvILjYCXPlOIYbLDImliclB5Nps0tDfO0N3dLvNUO
3HCOPgLZMtYnP2O69raXRxEffqEbIX4Uygo8JJgaODdurF4K+Aa6fwLp15nol9et9eJOHnatdiWW
V5EdPNUxHJGrMzta3EYAER9Yv08s741ri4IMXR+m5Eog3NMIvnPSjfsBmE9zrlYmaYTcPH/W9aNU
hJxaZRAdFLSi4HFlOb768SMCOxR4RaIfMCbx4HUDBc9NwQ9EazzRG/QqQ22zOWjouXKi5rSSC3YX
zAvpX2lzin4JjgNWm60RRcfO9OSGGti/xwj8zkGQN4fn9tFIC70umoiVSKNvPhq/Ei16ksk37Wr0
L5toOGoFzSxuGRBAUxo2I5yeuGsoz6K09KIPKJHFmzJvMhiISeT+aK6HeUnNhL+m3HnYUKOQ2dls
19P81nUdp/0QZM2TssNkS8CW3zkdcnpOlClpyWKeRpYt770enT6upJGlttkyx4OigD8cIFnRQuVQ
mbvyBxPjIRTNYZBYTHg74oHWcE6h2ykPhRbIGX6iIVh4+QklqMt4jHgvah5Q+TCaV6xLJmB11Rmp
/NvtceZn6RiNS8GXtAH+du2iULDIBN64EovBpCXFcqEkrLscWFAMSlCg4jToIfvBODyQlOpbFCUq
EOC1C9NDVf7Nf3pG+qQmeAIHGT+fUDgivrtGu55EyOZw68gAjeUYpQIjgbH52Y/2B15I3M3SfibW
pgPa3phD3ogJFRci+U8A40mLovj8W2TTRDVFhWYUbuT9DCQuD/uDy97qyfyhLMBN8KLetJ5AG4IY
5PX3IG7XSht//CKpoh+UnZdR/0lzDykphbUoenv/Cvxra2PSjEwAJvic3lvj8rfbJRGG3dg9XaQa
mNmVTCSUG9dwig3IOBEiD69VHhX78pNZZs8znCrwaYmF8KY5od0A3Vo2Ppr5/0SMRKzaOOlVKmDr
fUTOL5Xg3o6xQzeyCbW6/l1ayRlXyRjLEhBirNE82PeblhXIW9eKRmFEx1sXBNwnwldDJ3igL3w5
ClAqGFzsjgUH11uLAZosJcZTsoc0G6DimEcKApRRld5ouwhMhskdJKTXdzWg7Ssyj7AGojqXHL1g
cYxfmNbzkTDmmznJL2+IcLpwG/GOTvUWGIk5pSSGvTeUsefNCYBGtKbKaHJWSfHguI9sWA3RMo5O
1guUQSwgeB4mYtO7Ta/s5pqyOu2vmfP3Yfxr8vPK8+hPSj8+2okz1Ta8Rq125QizQ+cCHXFAXAjz
/JD85rCgkRGVrcGdv+hINSz363rBFMWcA5mRNMWqu76p/E7toHFE5CvDOpcMPWXTkACEGvCLsoaH
oBWydSjnISC4NNAUUP9PoG4C+fkAVdujP0YuksOWTMxvKLOCXn7iscitRN7Fd/y0uwq27pQoq8Jk
nuEzNJxYO/SdvH8iEMBMB1ZyrwwKaJEabs59k0HLLGlBKzGTmvK0PZR7+RX83V53DlkFvLNXxQnO
fiCPTPOyPIAjtpf7AmgyGDV/JxAMxdDbsqcSqElbSnp9iUykTUPm+i61bhjcgQjtzifymEL22Rw5
Nr5zJ1d0OX1k/qZtFSGL7CMuYekznbPcgj+XIKoWlaUgR0oTNvK1saP4P0IZi1oxdmNrOpBOaJEq
8zn1VCaAPE+3vGI9Oh6yqGy7p7OAk3/X83lToCHT0Th4Mw3390n9WuMjNBnuXJBIwWwzTEKkcQfv
apVVEqgdhmzTKSu5CUh9FwG1hBN1Aj2kjCsK50yEbXwsJHN7XtZ2+YewDJ7vrvwQCRwuxgNqspON
P0GjUpJ7Q2VjBZpY4zM3Td5hUS4BBnGUYQxjaOn3cKE2ohtUsLrHsipFXB87oJxfFfwmkahZUPQM
qfVbHxfA5EHK+OYN314S7LgM2Q/B/R13JxzRyjEdQNWEmr+4g2NG9B5uTUy1At/z7rQMhDLB/p3h
iK4j+guF0F/v+chkNQzKZNv+LNM0lKX1sSsBIdzIemtVW886uYvTxswM95bEZB6NAdBLLyPmTgWb
aalULzU1iN6s1uLmW0YpqIocYQTBS+muO4dkm8+Fjr0xqBjS9NY30v8zqByoGSknApotFC8lCkX1
05S2UBYVV0A5z1bIXdKSGrPn1SMV8EYolbdA70+ULU/+WvYMaRTFA0H6Dbx0T47jveAutFHM6uCT
UQB8WC+KWXIgeaY09TOcXQJCbGXJ2X2iWS5dhQqlB4aAfcrzEIHH/MwxMGqhU84Xanckw9BOTmwO
jagv8q72Z+G+N8u/18cTIWrQ19r9/bKXlNoloGpiu4Yd8U26ZoaVeWk2N2wtk07aKLzb/IKXwExQ
e+YSjOTOqH0xsk8U5t1txuOnFHpy2lp+cIG+ii8RZCmHWviLbn8GOl9/gLmgy7xXAyFNPKyRT2Pn
uuuFL1RnNOEzqD/448pFtGoW8BmL0XDp7z1uCJlWyJAC9o2W1122Mi5OVNz6IL4YraXecjusd6gL
CFbJFzo70pHzlI/YLEX42wIieq6PrW2lrA/KV2ePXYAvYHtYI94PxticPzfo1WB+GLnPzabwrwgy
CVMF23g6GJr/Ee4eGd8ZlxaSsnx2xhGsFJe626pMihZUMeIjg6RAJ4wYRWB+PfqWEgBbjMNboV3s
yYBXNEuKW0kKoPEX79siiEnBRSWl+NvLG0S17tT1T//BohC/qoQTSdfoLLQEaC0VqbS6rUFFWBuO
p/u0dQyk7PNBIa+SjKkbGtInDWyipYeWFPjCLoLz9l1JBqVOJlXsDZpLCp0rYDbDpLKhc6+mLmfS
JoBqPAdE4NbLXoaB/D59Jk/5dbHE0BCwbupCwEWbvbDjZxBrpCkPXPzZKIC0SSITBFfnTBwXQPbE
24cTpFE247TL1yZKfj3XWiX8vMg4h5XM4TpqNsDmahtoWtTSGXcHQgqi/dSDQ9+GX1mRFCQS2VRI
JxY3s1fq0ScZEuiO0NI2LelpNeiDURgDv6KmVXZQDVRt3Y61eqKHR7DujcUSeHSNcEjTGpxEkxh0
N4/MaT3VDbrnRfV+XVN6KIU/ADQARigm9QrhiCKrhfCdaoP1TcBP/EECYLoDB9hKTHqi6uFeIz51
KVQ5hUGQNNBw9ElxsixqpFpDJR+RRx0F3hySPn69hOqDek5m1VrKaADkaTqxA+ny/4Y8kb6TNOPe
mCuaFgrW32eiBWWYrc0tD7H1prnHWKX64vFgO28UdmK3k9dAOjv7a4jcG9GpQiYN+l106bGlZIM3
5ZEvrcWt0errF9/DlckHzV+lPHpODSfSxmfzmHNFz6HDhq0n7KJrpeq5LhvxUH0f42ynBBO1EQgH
IGdPJQ/Pvfpa8GnOGmnyMGx8Ug/3Rja7rpS70yI24QIjmPMlK1wyl+7SFT7KsrEVeo4yDV1I+a9j
k1lbzDWrKrQDsYDVlDC+j7Kd++7fisfGKuTRYguXthqVcgVT56R8jg7r/QrCyBmXb1fT78ACquiY
zdo5DBkvrBsCu78Du+5uXSySdxhJdy0FhLxYQx8fWlRymq41RiZCOF+jPLLVI5e0IRkcfAnmQ8zX
DvNv2+oQJoBdzmidsCUkRshF8CN6XTEWNiNSZJir+GN5uE8P6K59iwo+Qke2XbDTnuG7lsh5wG4h
826vnWHMlZzqujH5gOZlg+8LcrQNDxRC0FzXR0bpvOeg0uz5CmTWFL9fOe9nyDxJIJueA/S3lwoB
Qo2Vq/jIXtYgYkDGkR+fEMsUdDRjFpSVye8LuC6DD1sXvMyQA9IY8KHVYHmdOeyB7iD6GzhQHPKG
1G1yVTfJzu65O4TNkvaESnpm7BaKfRwx1T1k+1cDDLOoXzlO5BkEfpR3nQSk1CRdyqn0O8C2EO7O
ptBzLacOb4QTojAeK2p9hFDsON5B1r4P7o8beOo44B41zt1HnYJgcosBhZCs4OfM0aGjx4tEZuRB
K0/F29mZkdvb02634a1OJ27n7Jq+L4gnkfCR39WdR3Fj0UjfaDDDc/kfJ9sg81vpHPFVIgdLyD61
kuWH00ybUKxRZXX4qzFVo9BbZ+mMSSJ81CixSUKlw9AaoMwcA6KuS1HxVs7jw//Rr8m2+6s6zv43
CeBxumosq/ZxCJPbpw6xkbItOefQamPnO8FYCFuWocLm73rUVWRv8acd4UXEzDJ7Ep2pE6vt4Dsj
qS8GlbJaSr9X6wvLWXl8Vdm075PV4aERx7l14ZeLqamFfwfoiwyy5M1XK1P0JDH8vGeBIA79CmCa
LpFoZCVfOkUDuo1I9MRIq0lGCzw4zm5aTx1ZsjmG8Tm1famrgXiNoT+xlJmuN6Y7kUS48EIYk7TL
mUOQF2NBhcZXqU+rFtn7nrYzUYAfOBsywkRAq85o1Ik/KFowz6iaz2XdIMMmZccoNjryev66qY5V
w1pMyyRYxchD2+0xJnATDe6twgxNuiAkyOK+pcoihWTrEX/UfMzQbjIakuYa/8c1+iVsiMCtl+rl
qc/M+aOpCZQZ8A2rr0u0nVfXQZcTaHPG5x5mDHqUI9zBApn9rAmir5CmkeLNyA28xocBjW/zRsEk
iaMaaZ3h5miVhnk4FkgACVyHgOCl5/RK9zy0AOyqgZB8+GNg6d973Zl5ffivghw3hY1NRyIxIdav
uIg36V598lEgrIHEfCKlMyMi3jzNhlV/yHDExdbJyrVAVS/KFCU5lN48f7lpil4dG5Qkd+s2jGFG
tJy5DTxqJNkNIvKztN9xM6y28kfsdY8gdq1oCv7lNNnbSJYs5wPbDapAi5wMNnbuII4qoDYrt266
knsr2xVkNmvr/H6zv1PgA+vZjj95Llb4nuzy0WBBZ8guab8mOgBuIEfhx9mlR0Us7O6eWmAOdLD8
rbUYqc+IQ93aDqjoChxrDk7UstMA7Slhh1v230BrhIiiYoD5c3v5V4ftNuUVuqTiT8oYxhw7ou86
3jzua2nVqHBWXXp5FS+if/L5C8A//NTX2h7Ki4bvUGtC49hdPDg6bejmWUcRSyYa5e9MjSFy4H4A
eUpESAPbi4JxRY6ICAWFd27VcUJ6vmj3MfCnPQZqHJ9njmJMLQg23tfojgYYYxpc1f43QrWtpf8N
XtjRbsuuBdU3rJicfUqI30b5BfdYZg9FkL+I0dblgRuj6+8qY/266I4h2WHUroNhDtpLPMB8e+oz
9g69iAV0zxMFBvtQ4ZmvCGjzHblpfT4jL1VKe0HpMTbFWpobNC0luRwRAdrC9MByh2ltHHkw/JaR
nBJY8K9Gh4zd/3xisQaQj6ine14dSBR0sAWqX8FCt+VSOcFOLpRR/jGtXw/cBYiroG/KPSWWZNBe
ostuhgyPnVn5mkaipZOvLpS/RVVJsMi1pEWYzkaDg9M6OTqVKryzjzoAxepnNn2C57/TFmkmqJCY
Ce+EaNdXxG489MwzMjc1SfPyP7U45ZAICSgmRwkH6OfNPLhLEMGZPpLRgYGCOXsXLaVD0uOTd8SX
29tVnA9Obqq3wrCxlgxlBGg2YlEbRpds3qT1BmDBaY6VmqyoVOC6KsYvN8uZD96Y+eofNVDf6JNE
nRDKXQuoDGYD6PdZlyZLCom5FkKKLeICXNnNRpHTSZQY6pSVLiVale0GLElejJsyMePznjsSjw0V
HRxwjGp8w5YftE8iTSpNruGKJI3UnVhstbz3oPhEoYvAQCrQruZ4yLKVTn954BFoI17i5joghgU2
MgNhva6PkXjYQXRwpclhTlWDdDZLx8ckefKsY9aRa/Wu+47dq1IvCvjHVrfWEvE82TH20QD9iUTW
AWZXfzbOzkZ47h+t+meCeFdobdSsSBLTiUVmQM91b7wehHo7RwH2GExBkscEn8oLsReu89mjwP4p
ZnSVQI0lq9Rp5Q2y1YUtNdc2cvUAYGeJPCXiARYo99VUOV+75ROG/jQ/YZcRjEx+Dqzg3yNyLdj0
mzblydUd48knoAggExKVLNUKcuqGf3tlnQKPhSyebDnxGoOChiwX8Hy6D5kKUbCt4EOMTn7tkonP
I85T9+vWnJo5Sw465BVZsm+qQTqkTl9gL1bX9kwNLdDMrKC7lP7KwjKhBVDErCqozUCv44M0aOEn
CYxDDZy1YvyX0o8RU1N881gZzwjzzkVg4pH/TWDJqD2HUpmgivP/xDnre1h40qfgczxjbr50A01R
8qSWjmnMWuaJLKTYI5Uy+cZgcI4xeYrR+Bw5eSo1PfBADMtccSDrCWcbOjmHbfByCoi0mx+2Fj5p
Rf4OqvrXcWX4vrzRnNUJDECawijni/EzftQg56nHmMdC9bqFTtcEL7QyGJ5sgQ+HagLqAqpZf3rz
D8KAip0nnXbSjnVA78xX4ZYNavknOHYhMm4tNOqCxxzmyTlgGSWy3M2Vq+4XvOn8bp6Mg/po7j8v
VwMg2KslzVwCsG7r8J73nFnFnffFo1b48PJV6M97MyP5Ie0RXd4ScTJwbskEPYzqV4up8G2/rrwr
6k54imwSkNRFLMpEZ0qlkM5+00eHpQKib9JpMhlodqLgU11oCCiImlcO6py1FspZkNN2QLpT41vc
q6L6iozB8XBfxZvuNcc8cyzE/mt+GRLaNxlOz01p7sxHwqZEas9UgKUrc9LbTWBaFXikvX+y0MAu
7t3fqQ/kSCFOcSmXTL/3GMna6ZezvGEnRTz5GKopP/jVnHiGyhqkm+h5DbaYfKFwQCxFgRF1Ypf0
U/UZ/hZwmpKixAUMyjUduYeQFsVHLICo6PQhDMZAM1b6qewQy3xhSPTAKlrB4yZP4rC8DZUXkZsk
uAesFXvo6bRpDgFMp8+ZxHzb3CJAuHSTHQCumtBP8D5P1pkhhBIEhAloQFGWos63Ue5honWWB8mO
nppVb4l0BkKks1CMuVHlubaOGnRXdp3aQKUmZx+D5mejZjBmq/0WEeS+dLHuQTqsE/hk9ZbNIs+8
UFFgTRBpwS87IitMiaeqmeFJW6Sj4yzW1T92jQtV6gZtu+A4n70PqMAW+l9wKIiNwERnpt+6a5US
kKlwm5E0hQM5XMgAXyDbGEkOqWSgetfvYtUIIq6dttcfisPao3GAsGk3ZEN4gNCyjOkABHfDLRTg
wza5zSGHkAVNaf6S607OWRJPv5dwWUEWaCgfjft/s8te0MeA41DGlF5RiOUIHQHggbwBU8PxU78w
7p7fTQLmZPmqxYxfdpd4Fvc8vlzJBZca3Laz0SHztZZDjZQKkYd2bvuJk5Bw2rL9hy3YAtOZN+QM
4we3vvvshMV8qYuEDMz4mJs5WH3uRGCvsrhw0v6y8GEVZB6dli5RZ6Qm1yZDlxz1Bb0g7rJQ0vo2
fe/98EVI4pq9PespqqkMM4z6FSdy2KsEhV4E3xDMbOYAom3QEIsLESW88VYzl8hmx11fZoRmjJWI
IC/9cEJOjGwAIPb9YpgEbX7ZLv4M2ecFC0MJU5432T2wqdBh5kwQVOsdk+94YFcL5kxP+UTqLs30
rridsoHQEgcOgbpg6zAM3Xg+m5Ub40aTxOeVwVSkj694H4HxnOyCki0/US4PsXMAxCSQcjOsSPx7
xvo/9sOqSWTBW+lH2u0RTS9+ABV125MZ41ZdnJ2TaY+oGHdAqNkd9TOfwPMkrU13BlY7giexH0RO
P3n0JPmA2777hdGsUI1/3cPVtbQkAGrC2helI6axbwLf2VlFlk/dwhF2xHwCCYxQqqhDNuGYym9B
8C9bA3frcF6cLGMGgVjk3Hw4ES49T438tI1u6uMTXN2T3sH4dzOJyqZQQ9908PWAr2kWTDKdjbb3
WdSP4UjRb7vduiBoIh4fNBjufpvf1ay46MIOvlKPpIUJnXS8K2CrwnZNT7/VRswp3iBLwXEwhFyH
vLxHN9BbKFNm3K1ejOZVGoczII6Zt//Mg017hhbia3ROVdXNOoyR8W2AHGfmX/+KDWuqrub+/4Ar
6ECmwsQaoJDB9iJtl2e0q2YNiwKRDUVMK0Jm5XfsoIJiO30wttQoqJ0yyxjxpLGrD6gIoFHcSeiq
a2jyvw0g3vU+QxVuupao9Nhx9/0uvpvy1us26wJwKjMJ4rJgm+MR8Q0BKjvkRXxtrvPmXbqziMAf
VzaXd1LjOUVNp8QvHhfQgF5saqhNEbg6pRQyBe4M/lGy6Mqz5+X+4Zya1NskXe7yh+iWqo0NpIw/
N4AiFgYOLHjFBglhbHOyk6SyJ3qoqt5zH5rXEI7G9FI3ySAgyMP1DQl1I+uISAEg25wuwQluYjnm
30DMwMa9w7q4wM/NGBS/fIxWGCx7IUyWL2DsxwrT0Acjfttlnzv2OAOXyYCGO3bUTw9Dz4e7vTwR
LWOr+JILbs75LHhrlYSd0stRhT1arfLccxlwxGYqMsPvjuQzzjx8EzxBTfIt7puEe7NVE5KeKM2r
N+o0Jy/+P71ylvtJNi6qOf474g3bmxYnzpmJlWGhR/WfKZtSr4TxFEzImm7lowf5eTwdl8dXnt0M
zRuMdGRgY2c+WvJpOM/izWLiBf+04JH1fLnGozd0QH98JClcU326wh+L1nlxwXVbBi5XxYG5zCyY
T1Vr/fqC8FEXTWmX4LeNq6tV6oAHxngBHD0PB6jrWikk+wG+d3hqzlkHwqjvFqrGu7DsHm4+GLbK
bpiCsbtRw7sZrpaXOkBzcMicmFODz7hTNttFBh6kaxT4eFg3Av8TdeIyrgmXB20tfB7tVPoaCdcL
rF6v193JfOuKnsUuXgMWli+Hr+i1rPvnJ0a0Hun+i9FZAAZTlsf/GW1BTNAmVQUw7xPWhx0LvLP8
FOqaaHFTFPW4sUM+IecCOUWdi2MjKcFvpEJlBAb/laBk62mxr16fNrlCSuABXGqGLVzEeuPo+c+I
Fp4drCPkV+WMXz/o8duh89iAHBhzZxYyXdJJPXzv/SyrN/lYm4tJKr+TSV10MXHAbh4jZGVWMPQS
9M1lZKfbyoTSMsUkHOo6mOoDewxwvbK3tr7tx/cG7T8WugeDUpAWLZnVJDS7pjYB4zKMcQCZ3jw+
gm5/aOgqWec5GATEkXUYg/KK7NOOcWqN2Bqr58GmMScva9oURDhqyGzg0p+F9esVXymqGaL6k5El
xXUjmR8PrRPoIijDcUnZV4w/mtsfl/Y1jgFp0kcFvVIghQZLS0BZXgPAhj3HI5zZ2p0q42WnODef
VBx8ElmHn5qzP/J1GLO7+vjEWbaKOQTnzDqjUU74/6ky9M1t9CYTvKqQn+k0ppErBEVQceoEVXBA
YWovqD2BOMlMKgL5Z6z5X1fyw+Jo2QfFIUACbywh9+QosKMekoOAYUhHMBSCkVNe89uiCeSxoc5Y
nETtUb2LMbrCE7eXCVesXESArNS1vh52SrgM12qzdQyD3fRt0C1HJWUA1qq48jg6Wj+oR540ck5U
ZwlDTd/5uzF79ehV0Dl5ZzZwMvwPDLa32tk1zTG2LDMrzriOu+GLbyX9Tro/N6g54sJX58d+TGS0
aOZyrrEzz6qq5uiNkz9WGRfms+xBtaBA5jD99vpZhV0bk0k9e7uttdBZiUKNPcU/ZQ1sxvpa5kL2
C63nur+i09rXrkErf6FWfhbwzP3BRKhNOI8TfGsB69DWYG5DxYmgHbCEflVXuVscFglpRlPpg4xo
otePJ4SO5Hg/7qU7DmMgtW/emasrCvrDPzMGdw626Ng7noZa/oMR8AbhxDUHcXUELIXXRnfo699Z
zevqzgoSvA/RyyLUNtMJ9/l0Plm22DO648NKqq1FLrOroQT5SUyDFurOIgyCC471MiKEAkfnXnZy
Grfd0dfNVy4XXPB4V6CfsfbAEkLuv26QBBTYKrVCSfR27t69zQbcgIgpaXBnwiMv4AX5uLF33IyP
FWPJGnnUUtFuGgf06/47r9OWXn8lIIr6KzmMMgUVmQRzuhxB0uxhMpbfKMsdM2wpF3FWaymqzfWK
D5w35ogMkX3Y7QzbSMyS0bV/LusGgQi4oaAgOYOiAZWXiCSWRWUZrTsplATWDwZnicZaH9TfZrZU
RqFbA8dnuXHjHA4tJcVrsaJShccpzQ8hwe5mwTQYYmBkRaAX7cm7hB5S14pLzWYxzDid0XthUBiN
TN+wNzsAZK8L0M75Wgh3moJfakmD2pSj43nrrOYm1hb0DpwWp+RPqZHZXIo+oCcp78Kw5M3iqX6s
v5oqmeP/RuPBd7c/rrDeuCw/XffEwHTPfZeZDMJN+XMhHXE9VXFs8ETNuCkPA9XMqYEXzCngmJ1o
y1Hmf7t468iGmEST+Lrpp10KKiiQb7n4DXp03MeXMl2m2NCQWfq7vUKkwL+H6GorGjjd3D7TBOnr
SPgKTQRvPY0L69ZndzPXT9Rfb476vao/9VCAfbgECMy7B3rVFIq4toxagv4uqNChl2h/Ir2EM7yA
oaUC4j7SHdRH6np++EHohYGyPCdJrQfwZN2pDBHsQC9MH6MDIuHH3pr54l3fPkMIx0Kv74vFaObU
l/NRfuZqk1Vz+VQGs8DLR6AyKtfBLCTT8HYD1/Or2hfCQij6L0ecaRAySLQd6MNmcfESgVg61tWn
5BWmAE+c5qK4IJg5S5Y6Z3rOqkLeSy1lRe/rLJHmdAhSphqaOIcBcRa2K8MapIuL3a0Np9OT0ciG
qgSw6pZxkboJ1PZNkH9SIPKPvDJR0/RASf+lCuPmBY8CSuhjUa0u+TBm6ITnxMpvuDXx0l93aoHR
Q0VfQCJLpUfHTuO8z9okAYjeivGkjO32iJlE4P7eZU8CcSeGg4gB4DzEccIPATAgzcmQlM2OEbBb
LQeDuuEwTmmr/9EFNrvmFJZGahmdW10IyXpKlJVlVvoM8MqnblVXYvLWb9dzrfODFWBGEiSm8od/
mSSaFAUp1IzRQVF29l1ZGyMYPEPEO2h5bOlAFxY/BfuQ2WvBlLRrZFZv3DxTJdnwmEBqVt75IMhN
pbloJFlNj1Rd1B0msRaJUrMPQACvuKHorPMsevG4hjsrcFmUy8TPU0TUYX7fOZAz0IKpc0z16npf
yDNIZHBPw7J2/khnnes08saHZ7ZcEI5XN5LPHqZyWjRn9x9iw42j3P+CbFQE3ZabTGRtyn4M8Wvg
pe5DxicI/GH4mcvBRRabjy6jRUV+Asmkf+6pwQiSiw53TJcrqxRJowua1d/dOtGLO6z97W1hAgPg
e5kpGsaDoW66wkDQ7LQHDjJZvw57pq4c7eATimc9bRlC/wOSWhulwHeqwu0UZsty4FHv+b/DoDgv
LyrVpVUMAfYuNXam0IHe4MPMPldw+T971h3IhkYKrkhyxrGLuIQzzdn12UH932WiAdpey0nt5QEz
nTnSAcULdJhB8Oaho2NvRxF576yEyegIUaGTp2Vo8Wq19TR7hS6VtjYJMXYacdhnqFc+GrWvnwHZ
9o5Bzklii259ubJLO+cuNnf8SDnj2Sshjfc0ICNl9oQ4ZM/KWQa5uHbDbtSxKaKSb3F9xz2Nf36o
aTtOIELSj6Mw07KpMY4dbwp1Eb8i+SOTB6qfRdEmHqdLh/MaOQ51p5GSs0aHH+PZ5msW70MFv34p
hC182VD157y2tdEG2VYttZX8ggPzeepgET+T54uf7/Qes8BITBVXtEtPqawtgaq39jjAiGcHno6B
5vmJ8n2Fi2pjM7geIX4pCbxXQWAdoac5u6n/rXtSTnNEBE+wX3RZD4JmrmgBttS1Vx3MqqL4Znzv
jg+oimpCP91pxKfVUD1daqm8TOJu7HIMxbCwABtMd/C8/BI5mQu2lHfMHaLOE1e+KYZxs43g0Sez
OrAA0BC3c47FiXh6Vr+nfEi5qCo7BZxrFiN9IhpqkwB/Jfp5MS9UzKDwZ9KeQnbzo2p4a8VlDUbE
NGyIUFgqcJ2jUceDBj57JLmcLQLVgku8fU6+v0jFITxj3mO/cF4M1JyyLcuitkU/wRXBp+IAWkXF
FPz2wIRO1tLQQn64b1/LRqtM1JpyxwmXHM9y96JOPQixAsWT+9Jw8JLxq9wmGPDz7jDD5ZgDRmnT
1BfMVSZhiy1G4qMXr665mIytgPsBfxcMxj805rKPQnkFM/f3csK7dgwKm88bWBAtT342HThx9Hr4
PtDatT4hXpcLBVBFkf4VSM0ZQ+SOEFZMAFmKJtWFZLFpbBk4zocaMDuaNQBQt97Xf65f8p3HzpQq
G9NkM5uZMLytbegPebuZc6gyvq2zip7KxJRFgKSnOdBgmNnSdSfHw/VslEkS2voqj254Hd1sVZBr
VtS/lRX1NVi6kG4gaKiMQXusX5pdnHt7ymjq2HseTRSgxEB7z2HSXvXchE1lb6RE07gZERcCdKds
2AN2lWdH4YHBAB6cnSohb2fp+KEv7LamAkmA3NET6flV09+KieFXDWcpABoVyPNlGiXcdmfD+91s
M55DWBb7NXpvv+638IX+ExUSVPDkVLQB3YjI31EWRfEHlebAUNtaYkBHdwULzq2IysKxEI30UfTt
SafpDpn/k0+N33ot/9rjQQkW1v64yWt9JC5BtU359QM6Z2IkO5VWe6shCPrXKFZRSbTKFplcmA/p
LGs/OP4bstxa2tidKeE1+jqKJb4fH3EgmVQdJ3fIVr7bF3wyeDnYxQeN9RtpAafutdWd0GKccYgf
kQbwMjDmUI9+8UyDbQPjwo5tgSbiNDWuE3wPv5jQSuhFkxrL/0lv+EX2x8WtflH7Rcwng5Uf02Ek
WLu/oTSBVHX4PfN5nEcXJ8bVjvnWwVQcDbPOk+HjGGS1YShmWQ2NhiKjq+2SW4rDylOhTlkmL9OB
jUzOj+lv7ICSMTJ5hqWqNPDq4I3yJF8FZuaR5r0LPYnMGzgnXQWLyxLced4CfZB0yUydDNUjVdBo
w2r6s0KThwOycAkl8MeIo4/1d459p+rrNhVim+JlobnmczUHSlhYyKZIgv4SSXLeLOoVz3IVtY3I
ldvxkwQvuxVaZHfudFECoFTpfWldfmFc3l3JqTxkhNF2EQ/KeiqlXR5nT2W1zOJFNfLbEkA7v3fm
S+PM9BGq19h2WP47kgSa9wvx9jxh+5vqchmcLflIkzl0gDVQ1AF3XBRudT/HyqFZKGk24hNbwQW5
aM/tXHIJAcCoUVlKs9oI6uPsHuttVE35oDvk9L4gwydZm0Xi3a3fctlFWKfgPaByF6wmGqYr5aKA
MxDOxk8pFZ0QjJSPBAup9QEQ5deCbeCf8gY4lGMuc031EeeYHAulVO2e9FeQaCFad0ycswtddrqK
BAao/A11VGcScQ1ASXAXyMvSO1Lc9YY5SW++CGzFVkk9iCtvqG+hxfUAmTs210GvKK9z6H1NgBwB
FZSuPCzUuk/t41dg9BGo9qAxiWDzv1YDfQj9n800wjlfy+1LiXDQ5z99vXcfs/57QuxWXQgu3zwf
sTbh+zAyooHTHU76qSE0sMeCSyjE4VlaR4+MWcdXNlzE4CAn0RYcy3bHC3izO6/VndR0sdEYJeVb
uVzkf6/+K/yfw/lm/NjxMPGIre+QhBxc4XZwo3iSQ3bgTfUCVkCky8vPMiT7NNP+t9iInGuj851l
8pLRSlZxa5D+2eHSbQtSqTdJFM+WiRVTsdlPA1gkaAaHvOpuu2ysYEDiAeFz0tIvGEK8sHiuwj0d
iSKrMfVP0rlKbNZEpoh6d4iT+5FHo1P4CtiCd20xue4XELAM1lx93eD5x3xelRni7Lv8BnVgTJVX
cy8hJBNMHLjr1jHxIgUcy5IfIFPftQVhqqws+wz5Hj2eweMjkxa0cO/SZ0Jc37lWNTVeFQn1tSN3
s3wfP6VUyhYiOXo+4a00DZVH6H3SkPDlkVjosvDOD0LDAif3PjRGy+B3QD39e7L5l/OfOASclog/
+fccR3D9SlwQTS7hXpKHicsunnEmjSeeQloFCewxKJ9A2O3yumJBPEpPjo+aqRYQtcAAGfYaa7Tx
s8a21BpkJkApuFa2SO1W7pVCsJi/fcEdiuzaWyMJ9kD6oDWH6AaVt+EId1Rz1wYvAzm8uBBL2zc3
M8jY3qab8FCa7cl00s4zGM4nCzUKraS2k3fH4K0hm35+Z4C1DwJJAcSZu62MXtcpb32LPq53j8FS
XtQ6ULiF/oHN6VOhtOQ2UOEtTo+7BKQEIpcuUBRWErJYJ3xjtH9ODUHye0rExx3YexSDT9d0Utxg
mXw/5S9f3ZEUhRaAf5/1yC9oWUI8ALTfgG74X2zHy0r43HduuZAAwh5t9EzAeVuDCLAmwFCn444y
nIPvajRNLGkprA+u0QSjSAOdXJuV2Raryh4sHjMAxna1iBKDdA3pEtMIuJeT/NCNGDWryM8MkMz4
prT19eXQgMCak6FFWbQyPlqgwmDFskfVYa+Hc/6KG1dI7XZxC6Ng7+uVc0bkzMqIgP30Spcz+uKf
FNgoVGYjU5AirZXN0QtkQxh6NkrgLXQEJORPs7Xn5u+9OVhTRX0RHGJhAgO13li1itlUf7xCxdQk
TMvtyXUYDR4hgRYrLX8r70Dv+SxUca5ntLSL7AbA6hwF5w9FFuHcYXkT5ZaPKzxf05L6e2wPVZMq
u0HH4za5gv+3PqoEXtd8xpf/7JJsqvb+YsC1GqpWEM7DQmMme2YhF98LTSXpOrlXfBdADzWsTDvR
28oQqyiS3Rwc+NPyIg7SL+Z/p/COTNYgwhcaNlVFvPDoDYXi8UBEPidRhyJPTvPlG504y3M6LRwz
uWolwjRJMTBATLDDMpR0leGwa1NXCM0obI3wIlXRr4MVBDYFp1RrexrnQNPjH7vHUWia7VkT1qD8
oc7PipyPPKP9YQBS7CxBVYrFCGYrnINofHtcst87O+KDo6sFfSR1fi06SMW/XTmq+28djaZbacPV
VaMijcLnssXFymzru47DPosolWHv1rMebZnAXMwoIUzIAhJpTmdpFuUTF4ykBaBbpM1ppIgOICXo
gEbWp7KhTBajXziP1auX1vxZpgvrr427Xpc/Q8x/Eas4ds4rCb+xKEoi900wjec7VlkH0ukH259J
9KYgDDF8bh/DxQ8YmGptRmkDwk9IMYo5WkhUlo9/2VXHgj0wcgDf6XQImBbXKPqnwUKSy3+1IafQ
7Xg5naHggIPa9amZE95NiCEa6XRAMWwla9w8FfdGj9HxkTeDDRTNOttJFrQRpamh25T0tEmeefdm
y5NaXKW2qltsyrcEmLNKCveWyGExpv9IdHF7nf/7M2cLURZlrhP9C57sxQXXmbg0Vx/gdKwrgfEG
ElfQUTK4cfY/b58aT+md8/W7a6Xg5elylnU3mONT2tLTvHY7s9wtG0N63+HnAtusxJZEPZTMSprh
4QjLD0mam3aonHr7e3vKM0jkMpZoZ2XCFV6VWIqv4ieX8djGe62szu+5YcIye1kSOD6jG/6XJD66
yxmXjlHtSPE1WiLZQz1bnZe8+CBlfqNTbAnJbOkKXpFPryU15zugc+d1ASeVCDIUYjn+Oibbd3Qp
yKp43MC+FOlr2Pqrz1vvDvZairVvH7xvIrl8VUSJ0lRsVdHb6dSyLvAvlLazfl2l3aBT76z6cYrN
fbTJKdlesKl1gFcZHJauemUCiQm15ns6Raqgq9Y5Kzd7QdiZfZ4dUWiqccko5zZ58DBmTfeEox9O
2joX5Ele3ugY4wwXAcv5tHTZovzBPwPy9oZJJxc79Bqb8hEs83ZfCXrHy7cB1y9CIqQgTju6T0Zq
J20XoPmJIjPD6jjBMUDewbsGgURxqKtV08c4UljkpZ6tSkrGUVZZFk0tkuJCBq364rlW6txpuMwO
U4UyKEVeifQqSOSq0ZqvA3V1U+RCTR75P51zL4Hz7MSayaGD25a5+qyuKzfQKcJom1UAh7YTioYo
F6dnZUvjo5Mv/kGmC7oJepG99b+gZmFEcjj2uJcaZkH24xR5nqEz4Aw6MwXRl27DmEa0iTmT8geC
5GwNNFoMEpbpovNRGBl2h9+olAiVhNuBM5TPTng6QzGQuNSajprCL+fDXuT8FqeDXb4CMnVhcjXU
FNkRT+W0ZZVc7kgBSioR0ooPSFvGohRIkE1aBTizpN0+YDPnbEaUG8G+QpCpHfLz60wytgv+0zyt
vvLzdnFx6mfh0nVoZX+0e3z79IfRSxprcb0SnNpD3xXRCi/izF073MXfEnzfxsNO0dY4WQquzfyZ
yTSoivMK+NUZ/FoTDDnRdB4LoG0ga6+NQDITeLIIFbo6CAQuLlp4kBsPZLb8hOMJckgUpXo3N7ju
GEx3HTHPAwnNX9+sHurj1cexiIUGcWirnYRhbClEtB/7lpIn2GN1QAU1o3AfW9RVq+l+REBllWpQ
dygkCU2dQj+T4kmuM/iRqVYqOAbv49Ca6L3HMxmGTWNSy7nsuOOh5Qp2N1zcY08TPA13qgYcfAFO
DlifpdGBFroPLW9sq65G1UdTYM6I2geNBXltKo1vmvctXk3cHAsmG6pHBP0Yedi9ZSHxZsfbZlbG
1p49jp1Ps+YmC3qovxJRy//33A1GhfD/KK4MjLCemMl0bhvPrNsP3W+I+RPgL6gWvyIBsdbfUL4K
K/+GuhzUF2af29TOLOXIlAdyBsT2YYIROs0WVGX/Rk4XrkOF1rZb51RolXPW1Ao+e/bvg+5/8kUi
AbmxNUP6Q3sX9F9oKbxZsLzCc7Cv6Y7mFB+BSmvFPtGIhrOc54GwYlq6STM1IrX/WnRVGT54XdFe
duLcyzoRBUE6INEwVJxDIdRXJ8DrQLOr0eTJYX2oBlHld7dfhMjiUSXQZynagGxOXoyiVy54Cg3w
umr2EupCfd9DbTQahMIMXJ/zE9oOcn1LfHmAIINAQNrJoxkAcGT3kw0I7iKS77V8dDOHLvJpQ5x8
7w8nG0bjqx1tUaSLotrUV3pq5vPLzABwyyIEHygN9DSzlQbWCC4EjUWvZFXOjSHscbIaZyTl+1RE
pr2PLgwkPoZjR3jKsmQfgLJaR+LyobNmMM4FYH+N3tbBAHj0uRlTXZDzePyrcAQbgcDtD8EzpPmF
20GfwLjLINMkyMV6yW2z1kEwtLNKYOdnEs8SRneACzQeoPotTY6ss+1T1KjCwXa4arAb0Desj8Ow
GFUQoF6ATz3CCMHJg7el8Ft/M13SP9BVaMPREmEhlm/BlHSBpFLF0ko7KIx3rIQeAhoFnQaE6l1X
DcIadmZlXGw2+JkpGJeBRv4+wn08nwQCu55VBTT0WR1Z36jiBNeWnilA3TgTHWKSkB3QSnIOOZv7
u/Pmn3QkBr3h539ZQS3/49Wdu5QwF2voHHLUdu6xbLT9Sppr+S6F0UP4j+Kk8vr9Zt5qtj85jiOe
OM10Jdw9BNjt9mqWhWEfoz/0zNkmKEzBV6YfN46wuXDq7j9M8jZa+PBSgi4xByOooc6Rg9Q5QDHW
oDRldt5VHLxGdpjEQPwXRv6HrRBCnA2AWoTOg+Suml/cd4EJicJdAQwbV92tz3SNL8GKCrZKRY4c
kTDoux/WENeusXnH4QN5xhP7T54ZUstNw7JUpA9Wrfk9MjgkYlteUjhkKcJ+T1zA4XuzRR2njscZ
wqUI4MZLvJNYHAMz3ZUTNsdtjrhEgX/Q3WsazX65lzVTk0oMa6PLSqYhVrACx3GvmiZFZxhP0kwE
B5Y7/bKV1+bu8+l2wH2TWlBOIJzj+HuD9Xy2cEvE+BCzgAyrXd3gbZ1Eks3wpFdvJgTjmsbEBRug
c1O9zNAkmK8SHQsVVhQYdumyea08lJDnk9OIHfyys/OLWawLZoy793XF39y+OoiT0HH71faen9rJ
vXv58F+nWriC9hSurYpEPMjrtmIaLso5vFvbwUTvQeJfXkKERGsirn3GNBkbygJtfM+K/1WKaV80
Cq08NCOKEhy9XcqHOljVZ5tDtPyJLxVlsHAjNapCvJQuPCIEZooWFSobCLrye7D9AQNfuSYwqmDI
gFogtWwFR6gRN11RhyyFyu3ySKpu2M2wUGBxnn6Ny3cT07Gn++bWXS3W34Pt9XRv9XPXjwoC3fbZ
/51TQGj+TunstS9CyffnBhEGRcBTlwHlyqE664Zim+3LSwmT75iAiDtAx1UIk5tsbl/GDfbPv7xQ
Hv61Kc2qpsjHZxJtzI/p7XS9NYjN4BmQlu5ZMJH/sn8TypM6v0mJ71PA7ff3rVHxapVvyNGnRW16
8+Xz6t17nuX/okXv/n8IaoSiSsLUMt/hrY7sLCNMsevm8NvE4Wd8Irzm9KUFyLkZLSzd4TqgKpXJ
CzQbA/smsQiiMmOpeO8MddZ4lT0qzaDhRHkxCPgef4VZF1MN1cYs5D2QpejS8/025IrR5w3AJ1qX
+M7AzyTmChpZCY6WlcWxheA6ARSereChM4+qzMF29Z8kOdF/i9TyvIzkeoEwAI4m26rJ9mkDdBgo
IuA5N1ktQf0FARA5yOhwTeKl9AucHnUERekm/whwjk81Bj4Xdr2AolrQ+jLqe7qmehofvMABHqGk
XlkNkrgiBjik5z+8ZvuuV0KDMSFln4AqIbsFsJeuzSmP132H8JnFcA6usttSCkctDM4O5UgvctRo
tGX8SdQAUVaPR9njcU6oaZK3xhQPI9XtnJiqPf3wQKd8uZi/UEMIfap0SoXAWbRvvI5f2hRyODmk
1TwrkQ4Rb5zVwo3jLRuB027CMunMvXM7XARSv0z5rqJUGewpoZLwX4tJWXNqLXBIzkNYwfdQAuAH
kJbvBCUloNoClZqGQFB5nzalgiPQ8LI+VXe7g4seFx6ffqZjwcKFHKc7APMX0yBDfLUQiGSvSYSn
vcsKiJ/NHGTlSwN0X8GNeSVHgONF/ptiLo4JwMRZew5e11LBDQUSsmKNZ4Jis4NG8HLqjVdeTBTU
Wl8T7fywBcJL9lWaDsTnIjSsDCS9pdIY7HYow8U0LVmUXrDvmC2MW50/LiDuWTXYv8NEKwsKcH6p
NJaSpT4sZhNppvISzxu/5ZHjC4kwmvg/5t2ZcP4wuRAEPH+oab/kGoQR8uZjvlVdsCNG7mT59gJI
AwfQ5foPivYNVJpATIg1l1gmRtARA0hgM8QH/cvwv3Whffz2lvC0CvNphjCfV7jO8RKSqEWBw6MU
2DCbTiuLBuiYiQ9op2F6uaESz2hvKwJe+oPZWyJJvEyz0XmTrSfqg26+UUj1fBbZNAsQnFKNckFj
dQgaeOVIEqD3qi2lzR/ra4xBaEK8aSX19VYe/r+qvron3usKpgoIRSbNnp2RuSI+0LaWO+B9hWrj
dqsDo1nejJ81WNQAk/HM44EgsvijFGGJ0Ap/ZDLYdrU+Ho61UWqbgp6wUTK7taGH3AoBdkjVH5ee
kRf5dQHWnp2BQbeEdRC/ZRVnzPLzV0OSEZ6KCsVC20fdy+uZ/EMWkjJjWkxjxSLSDl5fDlF0vQ8M
lopBjgku/tqwhRKxiWuHe0IlqpZ0gvvRFx3y8N2dgVCMiuy5IM7rGpQWUwHeSvHGUZapd/xAUS+h
fAhOfxuYEiiEccWSzaNBOI8j/aWVUELGv5tU/U1CpuW6YqVthD53kHmNIPcbDlW5xGMjvu5UcAHP
ZWrqHYlOibi7jjQUZ9sGy8X8QBaxZ56a00N7741vE/WaSOulJGNMHh2ZuCtocy8+IjY7E7rwc2sr
0qJwhHQl/9nyO4dutaQ2AEiOm5utfTovvd4aTPy5rDC1jh78PICh0upAaz6xiiG8f5h8+KgN9sZ2
rYg8qTkkviLW6QIkgeZLDjRNxiyu5AnWj6ETwAf6p1fNyGCb+CdqVOHQfpwlsjneMcTYGFSc5llc
rjeL6wBJClhBD0Fh6WQ6O8wxZG+aAuxrLR39Y7kSLbUIyUGJOblE640LrSbSnp76iJ9qon1srrZi
8IuDcPu/fxe3V+0g5wQwN181bthEXHXVXSiFETYr4zvhuav6WmvZgbYui5HE/tz2SsKrY8LRut8E
Hqp7TpquN3OYU3nKe0zF/tOZPPDinAosIb78bPzFapsr2ntCc58e5UCH52FR8dMncHr2ycmOmHd4
Tc9n4DO5qcofxdpdgrzLfLNOk38cbpJysBmvv5VPAltUOQ0k6mGE83/hH3pg9WnV1aKe9BXetg6A
0LtLb2Yecglgy1yK1ODey5ScKRprYHy59sGy1jqIYe/hUtR0sxHOnzA6o1xrzeBEpDUrePgHe6Et
vgYIYSFomIliVJ/THQbtQFDTi8VS+s5tQ2e+x/0VOt09IVigeruCFL2eLgKCCccZrxPC5C2ZdfBe
8p6lDBmLCU1Uk3gWuKuI6FleZ/n7LlBtXh6Y3677rKMfjjvBhT8T8mLpO2/uKLRX+tR0wH177nDc
z2JmZKhFZkufoQeLg+uLo68YmSZgitOaXy6jYCxhGfJ0Clx5kdO1rXkMCtriMaXJUEt/FInPxoT5
JWONQ5iky4y7cP/CWmtqiVCJR8UmljUIYNmCPhU1CGCQGuW6iQfY2ewuQQXkpBwrOheRmLlHo4KV
Po/TjLhGQxfLJuBw5R4H81kbsqHVTVgtQv4EkytSWjI/bL1ICeUVGtlw0Nn2WkRHLTpkR/zDpCRx
3S7Zr3IAABwT1kf+tCzSeichNQ3PEP8NMH0akRR3U3BYAQFq6oxjiHufhjIvx4PIgZZelfY3m2/n
s2VmVv7aphkj6waSpJAq55Vv55h3vEmZZeDGLdFhVTG1N0TARxhPCcXF9NzXbQObyP0MwAXyrsOJ
PBqWwG2jHV2HLvkke9nCLLRgBQZw7zlzFwdX/905I0V27mJPGQMqxg9O/FfqDswyR9mpK46UPJLZ
L34kDQRI1I7sTSFxd7bJGRySXjfE375AjKAEySPQ32WOb5fUa+rWR58arcMLYnPTWyz97kXDAt7D
vXH1XSRi8SRMh1c/s/myuktRFylJUQHHM0mpn7nt4aYXRLsogpCI62Z3R1aWE1zwzQSQyDIuZd5Z
L3hNcKKBqFAU4R7MFdNCHsIcqLK9he9DN3faEmgeOTQuCAe8vup3Z/8tX7IkmaEZwbo+k3O6hllW
+fsRFPct4KYFNf2iqcxAgU/tuV0Cj11YwevOT1KeYwbr5PiKgFQ/l7UhllRPP5N418HikT0PBk7I
g+lryVPFcNIfUZ3B8N3NgUCvvvkUsIDWvonJaKqZgn3fHqhvGsYcQUzKIKGB1cf8+k7mV+mC7Apo
GuSHvM77l+kCDPTcRHAvSdwRR7uRWJlUzx6k4nBpc22VcclcXAjl7l07f4bZGN35SQpgR0sxlKlo
WACeTpoUUF+MMmZtqjAcEdiA7YL3ltE7/RLJqRqTlJd8Y2HVVXp93T7bUY3OYL8tC4M3miQMFIse
aJ4r4VrjPQ7Q1herghzG714rgE+f2AnWfJTgTSYT639R9NjmFgjZgHPurwjpa4WOn6lEUe6EkzV8
cuOCtyY4qBjbAJV/E8uUyL67neMIk9p60G3hqyqNi9z/h+HRNZaPVaavqyAugP6v9VOrLn3FQn3e
qNj96vIMCuaj7i2vuPSM6t/FENRS29t58b8t4kAsIZVm5ZyQPblRGzqVzBq0q7IPGyblSay5gJkT
SVKjPVrMLuzJQfP/jPnel4TdEGNYu+hdg2DbG4S1Z/SDC+9nUvnsDqpKUFSNa5C6D9M+YYFlq5n6
x6wcCYVxkUz8x9CnaOnhSN+qLZ3Y0CQDfdPaTzrm+iDo7kF9D2SBX279EYKxVYYWInkwkaMeDER5
hTvImUXRI0MuSPJZ4LTfeyZ3t1F9jwh4G2I5l/ReNn1ZFhvf4tKQqIg0Ts2lv1IYqLlmFeACDBFo
Ls14qqBT643EVhSFy1uu6c288IQyRUBbgC+VrC71hQeJ8UCW35CWqQLv20zYtqly5nEy0/zpUOgp
tOikJoXYcbkx3MEk3vvc/2rrQv1igN2W3S1lKCwy704UuHGlG740+pSFeB/iNIuPxkCve75pkwJ3
cg7eOqKYWmCxAqa5vlnaXqzMnp/py3phrFmnndCd/NkEJBvYnxLURsj5gGSR4J5OPNQ7GdIk3xp/
aoQyWoeFszSyKNMaH6ZsiVmXb4WluZLTwiW5+m2FOHjj79oD2ut7pr1RVrMJFoS6WHOGU2i0T2KU
/nhfSgZcU3Tups86dYoiVVJt6tbwv04fq1Ap2nwdDrsVX+dIF5h33bRyHR+Zk2RkVt1EB2Vb2ZbJ
ZJJVaOeQyKu559qPVh2EwuscbVd41MxtImq4QlCkGUq3hrxB/HE0H7ZYqbtvyXFS1InWpNd+TP/E
JYbHEkfHXhNeTjrsh1E33bk1LIpE4lgKqzoHgN87QFj7oERDO5s55WL3/uTeaJukmO3NG95aDFAb
JYRDIErkkPhs6dhfzNBVQmD3exBNhrGgkGR8k/5UyyyPkHgHneizAJdkRicbzuvr3UbL/tXkwqMB
PsIhURyg6BXAvDachqz+Aw3+hCUMSSPg1g09IfWEX5kT/UIBZeVx58RYlzd02xmxe/kGKzs9PaJp
x3auKxGtdWVlj1fsKcJaZo+zj6E8w/8Bxsieu7YJt3gB/8QDt7y3ufxPBiqfHf58l3cQFxROco05
ezeoptlqr6Gf7VDUluoNqFcC0yD47GLQYjO6e5tI9+tDskTMNICP2TMP05heQZpmgC/MvVS07lmd
10ADOnaeGnfKvLCHxK5QR/S7pNeOjZWxPG5IlZluAfNbELOzwPUPuW8rva074OsXscra47dATp6E
a/KBS6JMqXDmEItWSr0hdTb7Gc9rKuON4trel2kApCslhr30qik2237aAsR9pNB5vjmp1PX4omk5
NAvTKN+VmeUrNz3LK8lp2MbifGHBVfaVeFST8qwdB4X4R57LnMLBYoLEgQDvA15PKsoasGqb8s1q
WTsdfzNkkxt5T+AB+5gbuJYgXDf1vGcv5I/pkVe53LosVUrbV+JK1xs2GN00hODTzWisA28eQwqg
VY4XBC4Wfa2GpNJkVPldsgfa+f2YSK1xjRmq3/Lq/HA+uJrtdQtjXquCS+nrYuhER48m7RixfsIy
BRWqQvFgBiIZeCYQ0c5bzZLgVTJxMBOezYz7+qqUrpFug9pIoTaZqJA00KcOoKqjM7lap5ghIE/i
czRPR892+Xbuqpq06yjdFPFmsuAj5UcFSHLeDUacrWEOm83hb5WWwlSjXQnRpRb8kPbtFTFvxEX1
YQMiI8saKCtNR9iOsNUzW1l9azzK9VPaIFNtlI3TX+00TAj57G9LuX+LNMNleWqd+xRn0d7JSD+H
mKKDfqeZgQU16rRddiIU3X5UT9pwbdx4Tu+CCoubHOQ+HrcoK29r2U7jwYavydjE3uCFNMfzOlJf
UO5+aGexT+0TdLBCdjGo0Q85nz/E7cBp1EkljAbsY4wGL5ZXbMGEZuM0GI/MHlA6IAQfA9+x7/Ew
dQAzVgGaOt58ixQkxVPacsbReEvULJcJlZmCuFr63jd4TX8H8lQ1pRjQ8oh2JJApm86BF1SpBUNt
SMcmwtA/AudL+kRkrOIlpW032qHRlgWn+gluqsGYvTIWexL+/ugDWVIKn6/Ofx2cTdmJT54G/8Py
Mlt5IwiSgxmQKux6WVAyZ8bi0l6X3LC6zJgAeQ2qJ9nhrxbRcdj3Iei6GfDIe/EniluM6OKsmnPv
Kdx1hnyDiNu0OaDBW0pSJ78kxWje5KwXxYnZvzBjK0rkiz8mSUHo4inEj97m7S+69BoYPUtfYAdi
FUOMNpmCuTVcyZJuQ2o7fyHbtBB/khJbed7eMLxtj7D8aQgRtmsjs0iXocpCba1Lb1cUbpSCW20K
3DNymbp1LIH4Laq5HKERwLSlaHhXmiP9K0HrBaRoSzq8tvGGC85qSrDef01IlBzx4G4KaxU/w7zI
6EpHhO51f/b10ZfrQAhJpJi+YX9Nf3MC6VSIU7OOKiOsR0E8IbXwWRniiHPjeVMGMqMJ70wH72Bg
UW9JyaJyHppLNXiHG1/ad1/jOXRKnDCYN/F8Q72vezqkG5zjU8KslDWy0Xj8k+qEmS6/MFHjuFvP
z1Dt0Sf+uzXYviZ5TZ5STDKHKlCi9mNsBnyUgSJICiGtzSmq7N+EvPf+b3L8AuoFdT+PVhd7qi8V
DRfcItj6y7Vtvk3uo5YDSkRe3px06vn0Yv2IJQ8kk3mRa9RiHLCRHlcX/7dsx9en3/gMMv/cDx1c
Gcb/wpCw/rG4h1+RKwCGdIYT/NaG1+ujZHBSBWzAb6ju6EYeCgpkUpYU8lubU7kZ488H1NeQrQlc
UFCLQ0i7NUz79WxYhZvs2M31njOKIlxiMMXtG7Bsew88Ji8vCxuiCf/IYm4hBQn6cdD5XY5bcGek
Lzg0Asa6jeS6HzsZUCM5y+90ZeFLcekq4fbBH6QI3lNNjfivHJZfQqSRM4pHpXSBHuDFVPBREnq3
XVD6Zog3U/2l734CAad3sWkrgVdm8CIG7a2tSycm2e2gAH4aQaGpvCRaQyB7Kk8rnBqwBqu4b4rI
gDZvuEmF5eDqeZBVMyVbmfkM6f+9ubBFp5ks5BqM0dTVO7CPcoNoQX5DG+E0+25bbxbydi1dGOyT
IB0OoYaDq3H0tuQ7uBHatmTExmbjOdNueFbAqtlQgMM5Ilr5o2Q+HHoorlLz5eglHeQ5QG0AXhmG
ZQd2wREGJj8y7cQLbA3OcWSs5A8PGeFhdvCgQqZ5H3JHDUNISRpBF9UbMcmYCNovx4j56IZdTcoI
Zq7EqaEdsP0xoUOybcTXy0HzKEv+YbGCfbZDJqcGl0leqSQ1MOqk6amfQ7MYQpOPXBSY4HX4cs19
PMqD1UsGSx4zEia78UsnBtnTv+/i02PSpXhMo9HB2t0tuZMBCn9X5J3cWfWX1mlGFeXrKMNId+rY
O/WcuN1QhRNQribkGnh7Rv/L+IU/NvGwr2O9zuRCUCdferS5aHAh1PXTTnI9E11KSy4lDHgkbCTZ
Yztf96KefRi4V8N/rDC9uCK7bVRH9ZJFkta3HIDPPQcfjN6fuxrlPSat3pbR4loQZQd0nn9u9E4d
k/jndOcO393ZUFQaTYuk9pni9Kvm0W/gjhNQ/pXNPi8EYYiUIel9t+gaYPNdUmVx0az/p4N7lT+k
1FJfm+v6lxnOg1tzz6aYRADniope8ecyXdZ7bNOqSfxi1WApq87KtImWqMZcGD6P9OO/yIDiAFnN
ioVnwCPMosT7NqLtWxhtTVQp69tGiih3W2x1+hFsSbUMfK+RHPiAzvNGBShUyD9HpHpydb6uHdIp
87kbxHAvGQETIEKIeeWjW4DiHYrOg63HxIulsUnYNagS8bYlfo7GPYLgk7nsnImuLprELFEWe4N5
2YKtOUZwXeV4ib3guRk8jMqVwaLEgtarusgghHM4NuQ6qIdrCEMJkj5NSgnjCqJEBzYfaQJMqpwj
+DRgdtC4H4J1tUdo6m509QXQdxgoskPD8tqV8ylC5rb60gI6pLPzkrgNhu1I/4LcXHx1j3r90pzT
JVB/Q8QKCYbvdBwUqHbu2q23lnNkSMb9hhxuWNo86S2Lnb2tDAGn4u1a6Ty9eE1j7+DYlq5L4tUy
jxZwEvWp+YHcNywoukkA/GVAabl65ef7/JeVkEclHxye67GWouA8ewGtyaX3hu4v7x+Msa4dfq4b
hNm+OkFBXzVOhY4FweUeXJHC1BR5fCuLumsv7D2oYfDQa+QAIyCiz1sF8E+KmxP/OqlIrrFLUXxw
Ux65kBl/UiTQyXfbux5YZJZtzL3pMpTQ/X9SRXpemrcQmtxISVmcXGl13xVBB0anGCY3SY0QXTpN
+4fPdIA7b0tqiKfcRDdDa3a0Fg0OycbZflJXyF+zXL+JeErqWmw+FHbwho/hZgamEnH4TKV8+mvu
s3MIWF32sOLZLpGB5fkiNcD70AYMb80RVn8WpNaJyQ/k6m77PQCPcnaDLFeOyHODFtJB+yHfGnOP
zB7uHC9LvmeuGz4yKExzBjFNXDsED8+Wv+fd6j5ZnBelEASCcfXxkcUtJuioqhQuiK2FLPUiSSNZ
Hb1oUaplbJiNsUtIJmK9neK6F5R2d2rgb4Kbdt06jrY3sqTr1r3+n8AikgDLNFl6IoAxGwOn2O+6
OJz6QTpmI14cotVEZRnLxNvkUQSkKKPzkuSP91SJ/qUegLcXdB7yZzf6wxZ60EI3kICvxpnpxRQr
ItAfqTPwOtZOsGA35963n52ByzjN9t+wXx09IL3yeFG52E4lggSF7VWe3snj3mQudpND0WfO9FKJ
flQzExm4VMRQgv7zwUlNPuQvyVSszNz0gJvQsSU2Hmu27AoaoFFPVQKIgGOwTa6hpSJnnALt3BkI
3MY9pwPmdkgahlvAvlDotVsfClpy24lhbTzOO5VSy7DKm/+TprRCDH3mT9K/Pjoi94XDj/6n99Jy
N4JuYlq7nww7Uac03Ctd7oS3EqbGgIyyecqpiMWeg17pos69D++to6JBg7L50V0JSDQ4UsOxeVN2
RLvuY2DfbS2o/OoSDm6Q5VK8d1Tn1UXgTKKNkWYLIbzObQv7QpEzz9maNQFlIffzdKuA/oO710dY
t/+q+DD0qd3dwh9KFtvdASKxBkWVRqeU9UQK+E8hvgRrwUmiC8m/c/bVF6isXl8yJanzpwrmr2qE
iXU/ugxO41eUVUfrrkhT/wq33FmDlDLvBaoIB5k4Uc0YViKgZtu9ZeSC01zdudPBqr0IjsjjPoEh
7mZD15Ba8B7ovhPCs96uAbGsKnwSsY8soCGPCGzbsEXCjg+Es9H5qti9yGS/ZHSVOqQ/zVlVLud9
kS4jy954mz+jqCv+wKqC8Thw5nFjXDDps8UTcwUTb4S7g2ptLCKS0w4XkPbRb9YJklfVH4Q6DY6T
jt79Pznqgdt1VSl24qBOx5Hms9ljebYx4G41QeP4Jsdv3wLF/9Qa3MV9yknheLnnUK67NFnLnhD+
kqRy+DQIly+mF9v4KvFA9UtJUmR5B+MN104E2Usam1/4fiyQvxPtJesJKVPOjBh0SZxox3hsuexd
CT7J+HWWkLSff6OVCr8MZhulrPWny3QB86VmXGHg2Adrl7uaFOvPwMLM4ZG9agVT+niM5DiAMf5k
IYmo0o529TWL75k4T7XoTaXWSEbiIFnW5Z7sMw8pADaFk0Ld4zWQzOi57yz6769/pESLyF8lWytC
h3P76CQh5sZuCiCnXH4ayLcwMPNM8jXDz4bM59E0AbPJ0a3USbSTkZONdTyeppS70lpqjRCxugzU
r3pdivwZAttzobHZMVbBN9fhXHEHaXb2ttiRy60cGhmgQEeQdZPuFw35zCfVa6riYYOuCmET0vu5
OtgFDwMb2W+pWaMWHa9DPQf2x8UTBvalqbswoMT0Fd/DN1y8LBgo65eKY3kRKY5hJuwezsjGqFDT
qIw8gMprxXmOHB79FVhgZO7x6/yb6odiPfN36/jWdcbcpcu4kYfYCODGvx/LrVcbwuY/foBRFKot
muZKdFfj0OCeK23582BRq5/cDmCJ5OEAXcPJDX1wWCYi89ifbiGK3l07eeHngZ2cUCNo0zxJ71CP
2TgL6zJihyLhTqhWrGouDA7vHjCtQexu1CdJiDlQz7jLCI0Sl9ht4kYV3HCz3XH7Tk/6qcFTf3/u
SxKmwnbyT3RKQM3DbX01X01B7uGfuF2/ckBz9cQq4FRCAgrobUpGWCZkC/zGUadQINaKiytgFn/Z
wc1/cH9EDHxc2lQNvxPU7VmvmuW7iyd90mrvQNC4kRf6SiLaqDZvLD9B1u7aa3NR41wtJwHnMDNq
14F4fYYVUQaqAmxBd9rHFo2xdGng8oDgwhVqRt88qgFj9nS2Jnhe+Ogcw2IpeMi769rTr5aV7RMY
gJ3K+xQ2UH80QNCllrH26GZe3u5k8+BCiPtTZzlA3e8tj3clyIJtCkQmHkbvXm3JgTeiTZrRaXI3
M1FxflOlkxfeNmQdGjUpFWUJ+0P4w5lLtMxxGcwySV2khQOQsESpzrXSGnxUSGimMBg7PfvMCdIs
bg2b/jq/EE/pufM8bbcDXFvhA72DlR7b9gvYW9wi7DcyUzECjlIvtpSMTLKWR+PBL4bSBMsBcnEC
78LWCv2azoTkmVlA7OpYd71KbWsme9V0WDND+yzj3KBWoYPOCCBQ9yQFU9UZw4aDI9FG/tNfDPjN
o4HJPLuiRCLCrKLxEnZKLv68YMC769yuicH63XN2lAjKq5Yx86837FJc2rpROPrRmAsgZaO2s99d
HrWfxm0A+lSbfUhjPv6b+tA66B7VjfgDIt74F0Z5jCYerAVIadeDMQ1ziLbKI6SAjGaLnZWKLSOU
MwS3FbaAIGVus9/xHwr1JNn7xia288UrQ744b8u9xBtcQ2D5Qb1dFxitNiFtkogs5YT3P0fKtZGm
Ub3DC+orgbtgVqSFibvWsfyv9VExfA7MSn9z05QRCUa/eg2LnCQOe9oce5lNvnx/WKU01AA9TfNq
qt/GDMwLNvW2wc7u7aupNovC+JYQC2L1YA/9Ju61oQevTXxUaeTP3Bg4RTC320IoVXUzDdSZzfq/
M73f8+LYBDyYOPtKSITlV/R/qpGNpJQc6DpvzBaT1IsfGWdDK+hFyFMs8G+1hsmzMA7bnsEA8YlP
9WdzEaFYBgxQ5VhNyzGzIfAMazXmUM++IG+5tHanrySM4GG9c1B8OoP26cD9V0RRahGUnxxJ8GyE
pgqhNTAyseJJ3RaYp7V4QMTd0C4jLrOTh7fjpxlqzNmfsDCzOusHuMYwRH2WSxS7+w4rE/RAeme3
kK2Df6WecEG0gaGefYocgPhutuzxrlTkhyJfsRgqCfT4WDvHv8pen1EkFWH8H7Sl5oHaLF6el/y3
EZcOovVQ6ZOnBI8wY0yg8+4pMwwyey+TXDVcoyV6gdbmXMVojDCF+akSqzOjRaoviIsExwhN4d5M
XoYLu65C1m1CKgSghKvKNHS0McFqVq+m+QiG6nywvf70qF7II9qg3VVv6ZCN2KrkvxX2HWMXgHLh
J3Bh0aeTbaMm3xtWzQWG3JZVC7C8vho1B9IE3xl3jhZleQS51j+YGTDVWyJHRPDC9edPJaacCBuM
n/2YAcbANqf/k2bDWgsW9sw4iTUfTiDHA7B2rTi2DUx8/SL+mRyPXcsPzKuDKTnxZLRSSHezJRAz
G7jTSr5Y05/Nc0kqKT+8c+fqHYegt19SvxOyY63AtZ+9jsgvHEpARo+4brlx0dSr15ML2MlkfjOy
Uc1XkTztx9xeTe3r6XTmg4ak6aUeCCrJYsb8iiu5PcV8t/+oajV0zfBbTT+zigOKnc/FZ/Fzl21s
QdoWqozlxNOupILPzhZzcP9mstUQuDxbxPGuM/7mCsWqrZf/89U5x1F3DpYHwbPo1hHP2sWkxT5L
6bymIQNBH4QFzHc2ESelxazvXQWkgqSz+o8gEO7e6FwFESOpho7NXkriaxEp4PgOvgI8n4e0LJEI
oXFmTvBUiAYfWMMAHg4jatmjgeVR5j+SacZCEZ/VEc30riNTInLZ98JhZ4zBvc82645WGoSnyu6b
I0pfdHqKe2waOmlmoxEDzSon9NKLlCLl4gKp8/wDgacBS3WUyohTdMU1AcO6kcBG2GZsWN+tyLFP
Wuz3tGWD+HCA8AMVZpFeCvy/MyRty/xIrEpqEj6mdcsp6ugRTfBt0mvR5OOZ78ThFndSNYDAeyJb
eQI1fqKpNvs1EkCcs2Q+59lPgUIg85PU+mdZnTNIoHau7neXzlMgHbrvhnBmv9nlrUzNHrTUGDm5
GOo9fDgcli8Wx+NV6ny6fgjSqfNXJsBNzIj17j5lbeN47P6+Zw+KSaxHlIdZkU7m4SCohpDEcUtz
OjJL0VMtZRovwwTvbc7LJ906ZjdTbj4qwT56qHxGzb6HQ2+ntEdKdVO60SMAVuVIOJ4fD/+99Paa
+aFNIqyYnQjVbbliriLUSRjf62wyo2fwgCYQxx2Ly3E3gH4bIBT4Y0bKsT0V/USH4OfsfT3Oabrg
FwWrCyLcglyu3shaau6fjak04Cnyjr2K0Vf213ZtZgAnRzYt851h4uoVAnea7IcBZT3iTy3camU+
dn/hexHpd7fR+Sf+Vqwo6sy4+yfWj7e6KJJgm85lHrhNOLk2dffBMeQfESsLiJdv7cSNlKD6eL3c
Bhfzw5vGrHv9832v7BApttEsTu/yrJVc/W0vUA1AJ2SiWC8xHekUL3/wrjQ/OJ3+c0Wshw46biXE
irRcBf2PSaFL8+isrkkkDdy/z1jrvVWYnJsglihi2oV6GdH/G6f4mrJM37RxO+/HocPhsgZ7FvdA
gj1rdUCC2gPMvnx9fXpyqD2+vnvd5BAz771Xf7KQLd+7fcJjAW9nyqDOX8BQPBQjWflLDNg4mJ1H
96dV3Pf8fk4lPwpjQbvGtS6uAVBkQqnhykw+k2C6ABplGMrKrVe7kXW96K0z+sVNdyO1q+TRjxSX
kvdtsMmBPqu1t0kHzYgdjeDYMs0rn35+BcDA/FPF/ovSinCjdYg61etYRc3jqyqpr914Vnt/47DE
IAY2IeGxzfqHcvc003auY/7YIkcMfUq+SDdXhRGNCtWnZhw3EOg1oaTc2TtZKTMqBXS2x0xNreWe
/HgX0I+JnEacWC1fkdXvjCRWLzWk/yiaaO09/DWInV6hJhmatopgUsSuvx4CfXXD1DIuz3ak6a+h
GCUqIo/na2vLCRamYVW/wXuRvtgzI3B4pv9ArWAE20g4HNHuVla7DJMEAn6Uqo1ouQnF5IcN0PX6
q64ZjHcskbJq+xgTRR/hC/DQKUgGW0kx3jodT6ofIr2xV85A0qiq7HsymqwUCEdtxPRe1ihvPz92
2cA8acn2CkZ4hKH5mNd9u4Mok0kDxcfh9cQeKppm/aToNyVto2sB6pa1wwcqMxJMFarDNBDHbZ52
vsjcdW3RtagBFRF+JqlpLoRDfP/XlwrGhSWDGK0vU2xHFlpl6IIEQSLSjNKIa7UXupISaqCzfA4M
hsicCv/ADCHQs3OnTnFrQx2jRcMr1I9Wuw1TAs1vXW7uSFUlRszTHvCPBPWe5weKgVag2b4XF92V
ygE9+fLgXOvFFLTSJIf6aEsxNejk8EzFFoWt/b3UKqDvhvy0aKQLDqUS3AGUAD5EWjZnXbV0F/Q1
/U/Mr+xStUjCiRAdXOqQmYXgCR6yMfMXVY8r8QafGSmlQh1WKmE3K557Yk/QegsJf7maPCHDFVxu
ovcOCwYIK6sD/ivVfoW8SeEH5eUOZ0cVI5jhhRMjfHd82wDU0b9oaEmd3QN/6Qrtrq65Wnhti9tC
4i1OLFMfqGdAGQcvlDCOKUIqNI/6657EsdlIseoDZe+7DevKE07WZVCE3jRXc2+cHEd3Xj/LTBfW
HVrri9OH89HoVd45KUXDhnscsFBd8fNSaMe/YTym11BIqmOd9+siBDvCL5Zqv05TUnlz1Xa0MraV
IniajW1B+S5EPA70eT/cjebPLjQ33x3yBZ/fZCC3vnvq8x/OCgP+98EE9cPnpDxxIvAkyPI6lIYR
IRI5IJvc8lIR3SjK1f8w9sXAKwX8md3sKSE6Gp9LUaV/tsK4I+iluatm+bOZaz5xyKRTcWYKK3Dl
/zIhcw/eHQ1ZsfQieklJS7zKHcS6RXtLyI7KRWENuIQWXha+MOF1FZgroso2ybL1xx4Nzb2PEFtq
tz3JL5FDQOiWwKafxcmZ9KnXBOy/zGadARlq2ShVSqE8RD2F55ZBYmqdUu84VncnZAj5L0MT+B5R
he+p06Xh18Er1iQHV01Nbp3IABxiPbmm8XgpAnnt92h3x9Zs/ojQsfOLvjgvEziSRZf5I2lNLzsQ
MPJIUgeBxw8Mz2AB30x8h8mbPkP3RHU2/8c8VFi1s6+K88PCkl0asXjYv7oRBXZsYp+l2TlzXbcZ
mT6l+2eBtnkzFwsTG12bIeSYDuuf6eclOkK5SKIIP9ukuXa6s/et8UCG8NP1n3inRA4Q/8aiywXW
TJI4zMyWYecgeNt6IS3gQsSBqdTPpBWImqwEtQbP0XcTIckjCkDpENUPmw+iRI3qsBSsOJVtVcDf
K/bf2hQPxYjQRV5VV1/+38zoNLbwvVhfOKclw91ve/EXa7fFCWfz4WuqTLMcfJJG7tl9UXBo1F3u
R0MrJlXYoi2Vq1k2cWzH6jK8/n1sigOBha7m77v1Ca4/lwBlAsAJlJw5mZL/VF2f3EmQBwsHegDI
NqoXLeyV1f7Mo8za/iTzaVuseIDWdO8SyzgvnN1SC8kifgK51iBJ0e+3d00uQFk0H4trdG8alIwL
szvwXJF8lufmxBygecTlrydOQDVU5vOAw1AA8pxz0/ZBl3fzlo9VesaAX+yDtSH7MMRwZJWi5OsE
IDeKErs8AQc71GynIk2B1VmWZ+AGluhtEE7tqfbJITnoEefJpsDdZJuK4i293c9nhqUgUCw9fpsl
uY1v+OyAqHseLZaydh5Mg9FJIFBP6IKQRqnxK4tf0AsQg08IpC+h/DSa2FlJNunXlPcPQICdsSpI
h2IGHg6xGAYPd0fGpU/57R0J4yRkS+rgfbkY4E4kQCMl487FwquQYmgUHvF71r0Yybj5a4a1mmeS
VDHGWD/GPcJgApvwA7Z6FRuhHwi1mwwhk6sxtFzPZfGzCc+0HcqTrOaY6UcGuZfdGmD1ThDVD/1J
F376QcMuZ/xOZ+qy4KVfOtmKCP+Z7i9tWJ2eWOguYeWfeYAZkYISmpBnW7NVNcf0PGD+FMAWjeLt
N+FueUDcxTtO0q+EYNbZFHu1BYzqAwjV8dW+jYI4JlJ3ju8WA8wSd1sDXxsISkI5Rmy0b2GTPOiD
TzDdK1Z2JpaUBnCBxlniAUUA2kiaRvzpZnW1MPTRljn+mWJESN8fZqHawO+10EPjiS9m0T3UtSG6
VL9uf+AxqlYMm/trOghhH5rXOEPLAI4Rf8IryPdJ9hAPN3LsmPA+zuHCZWa8ZJgQIb4hYwXl1wS3
t/Fo876/rjyoX3urq9yESBQQWrOznKEinJ1NPO0xmu/M0pPxOnuwtjHpGC8Yb7gfZ+wCAwHMW0Wx
qP0Mh0xbuCXlAPjpdyh/65DMGCYtilER/zC3b1ggAt6VIb4Vlk2iL9rmeaef+GP3NwiTNAGaqlA7
ijG0JB/9fpwQE7TL0zQXA1enNOD9utZgYqKD3bqAiObiaOfki1YHbhwOHKM0vkJ1qX2CitzFVqlG
0f47rPuRUxuafuDZeKGqlNMxPlyEcApE0ZdkOoI/4ybZW/Yx0ZBI9BxiisIDP0GC5So9bkbCskPO
+BOUqI64CUOAx/XslsoYBBIRnaUXd4bXKBfvGBjHv6tdT5cWh9ld2o9iLh5BdkE6b2D37PvHmRNk
/TJX5JAJMIRoDvIXGuBXO+BmjHoPEWXYRAuh27ANjSio/bmWV9cQhyvRnm6AnXzrIC5yeRj1vwq0
HJ28zabwEWA++GDRc0EE3tfQa3zlGOzDwa4kTatzr0GMRzoreH77OV6XlzjYVWrl/Xjd0co73tOg
AXwG10XSbZakAPpeSdnQm9H87N3wt/Ochk6oMM2hFBiFWLzmRdcAO+pzmJ1mfceTNs4aBSkM/NF5
nb2hZwVI2SoRVUuHtfqAc0K5AHg96G8KiJJ6tTo8fFIqywXWHl5yZHmHcZfHQcKK7riLzyP1x/u9
81xoLyi7COrCl+dBLuIAfIWzS6tQRcHo2ueo4q9JlWh/OSAM4/9BcwUkBBVzsgOJdLH3Zcoq75Z+
6TnyGQ2DVW4upuN0uLclb26ild/Va1jYy3QpZ6tzmy8EMWZ97wq6E+P0R4WMtIewg89H+nyuxYyz
HEjdS+kSNIuhi/J1yq2o2DO7czlFkrJnQ0u2l85LvbLG+Dp9nfm0/gTi3y30TkNlae+BJdn+0o05
LKhspwto6n6lf+iRtFyBA0jhcLo5x/AyODBHO7sGMv2iEwyME0Bq1244iMExDS7uR/NP06VhcAwY
crn74PzSajrAhFre9xe3GGUSZcG2nQciCFdn60QlmwCSVQwGQO+HD6vyDueMUVFzJBXQwlQpEyw2
4FpEevrSN5UrLfUHTt3ILksHw6Piu+0P+wJkWyxh/uCb7ltHV6NH7phoklscPq8avrBgIgbLNt8v
w/3hVzNErXATHbBGumpEACvw9/jlM/wj4EdKlyLljC6h0goFCEngvtHwInbWq1Wzlg1v26dbPnJ0
af0na1CE9iy/1Y3TFs2ucH+PQ5YT9Qe/R9AM6rOHEW85LzPhf6NACRYb3onW8wFv/5ZQaUZQdwuH
zDy6e/2szo3xNAaT8ezFUZdRFmf+/btllDhiMB+/xcUogvuHWPfVE5Jtmt5AhzgI7/BxvDu3FiVR
WaKA0W1Csf3BXn3ZUmJ1Y7Py0JRVV1fk42a9jj2ITxUVgcnYxK/aj3g82xaarhjyYJgmL71HwM0W
lZc7onGCyePiLJGC5PW9XURID8gfdqMZp0LlaaihHJr3jIv+cOUnbNfKKp6e8GbE5FopGEd8kjUw
TXKO2szisgytRofEg+NoIF3xoOKOBmIPn6OYChYIEOi0HDTkW22F6LmI0XHgLJcp811YypKDG88p
SUyFKTU+mJhGyqa3d9zSSYs8y2/dZzKq42ALpu4kOJo7kCTcYHnMF+SlPEjUF1878X+N12QqEZXb
OqOjpEz2U4MW6HCDiWO6oz7oMqDbockP9Zw47RSWNwXdka+Uzdp/5mInyd0zsimjKEt1efzozKX8
qLPEoYH826dHYi54qdvY3xfHvD0ttcr8IHjY9ig+IgW73pa7TdTFZ0rhegr+ZTdyJDJxOc4+6FME
cdBdBAFFwxQHgu9RVWm+SzplimByWPQybRmzKP96H74UHU3cmwMboaxhHxUIUhqaPQ4WrO2oENP0
NovgEWDIpkEM9PSIx9uHLM61lsJj8mm0fFMzTQLPNAaQneYoP91ryS+ZWP9AEBcrh+FJIQTR0+zM
DVZVbsAU8Fg2HehlcrMkPS59/S2M7BYAum9ajqxY13kz8y7uxESifU5tvDMTsyfgh53NrXyr7Je9
uJR96engM7yIdjuzUkXi4q/prT2Sx+t1QFfNOGz1yI0fNnn/KYQMb3FLmdJFTzEKAOH6e7THMtVx
kGRuMiCiiqujmNKlnx2KU3KSMMUxkIGtq90gZQ+uR3J6pNB3FMULTjPDtWp+GDIIWdt3s0ICv0kI
GBroNl4P1Y/OuGXKQG1dqgDp+HNxqgSs6+KKnVNq68kGLveu5a4ZcQa8yfeSxETQMimziYKMF8TV
zM16W1sSbSDF0LYPC87VAk9nZUL3+YTDX5PKzLAVYmvLsofiBZwsCfgyNe4lTMyYnMz3zz2rsQXq
ypHNbIBSU59DO1d+iCol2TAb6XwrUUK6DilscL7x/5gIDxBZNSB65stI6XmR7HQQZG73lByuloDI
gPR81HztWLaC0pTD0maR42oEfruJXWVTdbC9uUjHBbEaawQkwpzSg/WAi86p+04+vFkPcL4q9MFN
4Fl8+uTpNoHDZhvRdTfJkJrp4LyuVOMhHANDn5C534qz/cSndBTmmKB2Ev8x5wGb08nGhE1YHZ+d
TvuR0+xJYloR+oHOa8wQOcUbKY/tCsS49FTswIU01uLsxXeAtvQeYsBw/jRZBR66q8reBXllF/tG
oFKhWqR8aXGwSnHrn7mHsjOYTw8OniDrVN5w0a4+X03PlPFoe0oUpNLKVsC2ow5Qm+E9dK6oFFkM
mxp8mihxvHw4VJhqss/nd/luY6q+ymO6eFDUoHWpG6Y2jL5lflEjXPOqiFwgDRaCQXBtAtnJvSqE
Lwef7bkJ7iIMM/zKL5I/w2pW8geWzbVzzaDaLlKb59N/5tnroM5zgSe8yImKmD6Zs3OWQWDEyAkW
ly7hN14U6+2DGeEyDii9K5vpdk8H+a+BU/PW/dx+Ii/TcuvobTg5S/MA1JNZfqbA0qh8OQdzow8z
GIfJVPgUuNEoJNwZCQJ7Op2SejxHuCcZawZYBSUXgJ5xjyUZLArm8EI2mloHff9T98qakQZhV8TG
rRRp76iYCT/o5xw7BwjofdZdB8VV67BVGHuvXjrrBoT3ntyLLy1Qnk7Q7wLawYHSPYh0Bt3HzcF+
3w+aC7ioUms3ENYTkNWorw2ETZCM+5/4mXcPfjvxcAiUUxkWCTZtARHDx3TxWFKYj0SEtk0Xp/jt
WOXWPwV1R8UdPVoLN4Erh7/K/RXt9XO1i3Io0c4G7BVABiRaqIYzHD1G6JYhcXTvaNV5CZHV81J4
Vd8RBZfDJKsUNludLHMSwg88bn4Xf4D8jThXUY1Ga6bD3HZx+QMh7nois+abGJ5Zvvx8DOUcn3rj
ZE7Ku7YRrRoIugg7WckDHYrhRbx5ySI3/o1HWGyIL/cnASnAn4QGQM9CQLR6OE8204ZVSYK1YrEX
GcfwwkTghe9y8Fn54rsJLZStZVDhLesvwPnv2TxRG+SZhqNspXrIIz0qO7NWjPoZ9qrAgmnCxkzx
863jXofUdz8gX3/DUb4jFI+my8Z91jN2fY5+b4UWCrwIh2/iZj7awcKEiLgxyJx99AFqSBonR+XI
foajMwOESRIpzvvdBTFTyFE/fSIjM4GCrZPwwKurM60/0uyiEtS+RrqbJm8nLMpKo0IHbZomYRg0
LF3SFSnto8rktiMtXQ3pibhNlbG1ROTHYlKxKGmDYpnhNzeWJflki6c83iS4yywZ8CP6aUCJVvZ0
oqDiZxPstXeJWEt8vyjchC8O12x+YERobMjngwTuggMoJ9rd1AaSOTqDshqa+lWayXsKqiQhGh/u
L2RScBx2Ju0qehl6n/ht4+Mdzt8dGnFAuS/DOBkU8hjusAcCl63XpSHijLb1UpBwddirZsTSnMNN
0671OlqXoDnAT+qZlFcq3dQwfYm6DaoxsbCpI7lEnarYP5faSmwO25zl3y8LhD9Iw6bBV20fXFBE
IMsMSmSvAMcfdiyWJ3Ib+x4/GfaXdlu7P5pqtmN/+L6DOe2YvgK9N1HxakCQVrMDIcOtRNTbsyyh
6IfufvGF8oRqR3MnnImwwNJ1PYsOuyt/Mg07+oaSDhs71g2doi7VZ88nJViG86/4jTsex+ZG2Rnt
L68MiR2F8z4Va7zAcE/2I+dUASftuwCH18Bj2bm/3E0W1QoasH5qKhSPqOnMo49mOEVZ7UK+iJs+
mncsJUm0vwivr5W7UGSm3CWt4lPgTjWGK2f18JLO8g2D/tnR54LyaIklEeiPQ/mMxprdetm0GiIL
9CIWD8IQsp7AgrLLJj8ULlPungCxDMYBQ0cY1qqdEjgp9952Jwa1zvWIGiFrLEIBSSqAKp6kA6+R
2ShSZMgZyG6MEmKvqZVwD67KnuAfGObF6VLBXgHZzVThAz5zUybHA7s7UrTRc4tmfoTHcY8DDafY
AX19PDnBKnWCpo2eW3JlnSazaU74ZPnEL1U++vjl75OsaQfXkfCFGm8LzwLjljPESd1ry0ljHF4s
DGU4L73xUZCwxIOK5zR0vxUMZWgmzu6gVYCLKv0v3OKDFTdu2txNPHfuNEhF88ZEsspRcabVqOX0
W3ACnN2OYTBVnCDATWYbim7QsLEUETvYXTvdp9FeF9czgZXA4HHmDru5LHaVLvmqDENCpwSrPk8H
nl4ziRazxllQyQ5dZumVs0/NiSO2lWVJ0Zwe0dyBSGP4Yq2PKUKhkVBs8qQiw8WQ3tansc/+0W6A
Ft2lcoicnsNif3x0gUKdqPj8auV5OhHxmJr05dx7mTH/2NlPmo9BrbT/s8ovoO1RRVBXwUO1p/TB
wArOHqR+veY46HaIZFxADZQN+T5r7OCSsn0w6Te7Q6DYpRNNmcEaWIro3uYdqxB2sfSpDFpt7/lb
h9OqSsyI/+T8/5mRS/LOWZokYI2N0k8HohGP4eDVT58I2PZvDlsg7QYVq6+LugXt3EvY7ipOtPvy
RgPXo0cWJLOGilJurdWawVJD06rMPS6uae+73veUktGlYFyD4clTT37KUQlpgQdJE7TzS5fF+MhA
q3+V8jicm8Sn8jkkJOBDpK6MefqPEgFQGIH9ho4UxpRnykp09BVe+J+LRhJt+/JXLV5Umbdz1nzB
KWahms94iDf8PPeIHMWJ5dVcqxG+JY6cAlWV2Mu++4pxnxOBM8Bd51rUNSVKMAwGEtYvqTk52xPJ
dcIIr5VC5Beo2eOP8fyNPzPKF6T4A7gDcpkbcpKmRKgPPNcHT58p03eZLPiYttoZo3xdQEjXIBKe
jhI3rtMV/HAP+2xFcfD2NjMRW+TrNYaPVnOMJzA8lPgkBu7M/9iDSR86SOTu5Cyq1Ohp0PWmWBlK
RLJ8IzmTfMtqhTjmJCsX8yA2Zfn2n1wxoeZHXMEuk+CQtcJ0gDQIhlryIsagJDmAjFRDvnZl1fFj
W7MAiVxu6R4P+HReYQ1fD/sWdVB4V+L4pIysRr1LrAogW9X4UeYOy2aObcfwM2O1ZAqPjzxPeFan
4gTZn31FF9wLl1zNW9K2PIKoFfPbH5InSO1B9KOCQjd0UM03DqlhSVV54UddNP7ysA3jdDXHiGXD
gy44dXBdh5X78tw2vSkI9EsPbh9emFGyeaSPyp8cqhVAa04lIvlUANbe1eGjCUpB6I1f3yJ60D4V
rP03uRYPKmA4CY0l8sW/88oB05Lj1me854lLo8w061Bvni5fhv82561TO9razfD6BtvMcdL8hJK+
gXaaPKUE0CVRYmDMVrpNLWROx6FXDqSbryUYS84bKmzRxBqp0tDrRKZCnKwF4DZ5sjAbt2Mc5Nzh
KN/rsBnaWsU5bWbD8Y4XznHbf+v4pniDQQNayJRKK5rfDipoDQ1q/3I23WGVjAj8eCcbEx0grRvZ
Y/UQ0JH8I57208ljoBkGLBXFKYJj7dxaycQbiVP5RtIY2Mv2j2IiFa6IFT7BvE4LEfMT3SYEBWYM
7tcny//k5T4We38LngMOwFPtVHwO0BxaTvfixWMmx6WcI4rqdgwz0STCuEbOaCWjzejxcEmWiD8g
FT1fFLW4rjORzRV9jmE0PCyzV+q2dddGB8IlUrs5oD7dxaI4uRY/53PtLzgFOMu1SK/fhRW/XRTC
jr+WxXw72rauzUrxmjhxlVyxbBZOvr8+7Nf8qYIfnJWdyE2zN76R5gfx35jgoWX9TiMOZvvLnN6y
XG7iyiC3Q4Xob3zguOEvOrcyuVdPSAaN1NkmqIHFhbH2H4rLo/GV3FrEvvTNzW1OgVwLEev6DK+k
WopL9rbWqs/AcrFRO1ups8teIsGNT/F8cg3Ly7k+G7R0GnVrZugZFIjo03do5FoC6dLSTCkqLkm1
RYZLKa3dJYP8nhAcFroHceJEEABNvsK6pXgTC29NZ02vnL1kdtdZ5vdwrIl/NcB4612Ols62C8pv
Yg7+sIyuJND8Q6DL+umIZxNkEqwFb+8irbo4e0qKgGlW2c7pBW4rXGPOZck6f/z1GO85Zc2vkrUq
OT2/BxuYg6OIV+iqKoMtBIfgPb/g+U47T6lRIzdaw8jIcCcqEMZUdo95R3lDsD9kSYivsgK/AvDN
n64F9AEpT6PdCgtLoAebizhMqrGkcbC1wiXtM/99L6h+3HygCnvGwxMZmkJK+plRFVc3dUitz8P3
D+GOhFmkFr6bV3u3uZvCs23zBBLD8TRXYQfZUP5P5KFZ+Z8nXdDXFkNs31cjZUp3f/jS4U3yy+0Y
4HWo3iQfxpuXApGnr+iHQ+RlugE4pKkP9N/60lvreYQht08e/S7oPHW00sCaFvbNmTG8NM/pXpqX
v1qZ1d9zy8tQOKRYm1dTQVgID+FuDe0oTLUwfRUlqJ2kNsUH9BsqguEKOwsahbVBtki8YyUonYZn
+KJ8ohrklvnW0u9hrnoNBu1Zeh07HyHzZGrpfPiiVBXLS3jFjJYubtIfCFSLnCQkT4WKU8+mmAHD
HxsZI/ROB1WuIOiq+NNKxrlqiGjb6HO3SPgfr2qWM7zqN6SvvuQmnVlUuBwJCaWYtj3RKR3Vdbk4
2CW2EDXWOxw0WqKhEUYF6D5j7OOGiwzA0y1QKJ8iQELYmfRItu1t9cjrM+SK3GZbpxVHdD/x7f9R
xMQ7MnexeNBizBANWMzW8tNycBT5RdDETdtZ3oQrdiw0OXtxqhv9KpQ9KJu73cokOF1zTSOIMh5m
slqk8dbT1ltSve1ujXYzMXEwo3hPPrF8DsKrKxG5kTZSA2shgxkDw6FUFEGQehe9hMqmdtoJzCDe
Ingmp+bDtW9EP5Rv8yT89o7QL8zgdwm9PCh+N2tHmUDrQtAseRSRNkXcKLTddFtCKsOW3m1LP+nH
DrX8Dzn48wdhl7Z+1hLPQpnZjpfJpnM4ZBp+CqQ8nzob6G4ZO1/WFrC40sJ6CDkgPSfFCMfyDa/4
kHo2qMH00f3gMnU5uegrRaY0g9I/e0SdepazJG5lKImCpPP9ElRym/6wEd2R1IC/HXqiYFU5oK1c
vkwQn4ctnO1SeUJEcKdE+gV3QF3/JYzEHRvoUc5QiKYrNJMmVwpwgaX/LfjXYQuVMhiukMMsHM8a
wHr16lDB4685c6+AVdY0HsF60kv2Qs9wAPjKaotl/DAkGpDxtn9pBJEHH8C8qhR7clUMylgzXe3T
6gRC5fVqMmmCouMUqqKeUlhG0Bfl+xVo4STuBhO0GQpdhMlJb/IIzwdosKw1WD+0ZLxpwsZrf/bF
qHWLqNgAz5erK1w3Miuxz1baFJ0gSZM7ONs6az7Vntt1joUbVuHvLufBjivkFm9pMAaQnLRfV98J
BUjH7aoUVM2zfp1cl+46jnWuh1xJqa938CC8s1E7HAd1RZtVmKLUfSKJbuOBtmgWk6opvr3aW+V4
335A3z0srUcmEhWC0jLoy/D27DA6OfsUxEY4K++wBEklYlyOdoAmrZWP5/f+P/nqeD7G/IH6dcge
1WZaNWAR7SD2fuiUyDtPCiKylonS0t4PnfJGpJWmO/ZvPqpDp7jdLOzZibQzjqshjBkuNxl2ffn2
Cpij5a2xBYYSzqmxEpxhmRClVv8vkfF3uT2/jaOMWo8WuU2KBwXK6vCivJnBs2MTBLcliB4bWQhG
8aa8UNf7RtcwWOKR/XI3xSlOdQFLrlyzANf7CjKz0Fohwd+mP4JUA1mqvTiGL+XGMSXbBamvlr1c
RLAyBqOaePwCS6Kwg7Cjfc8KBF7LokqCSpHQdNjCLE6QUCor6UdaI6LZa4OiZ5SGAVG5etTojNdN
5VQhhn3ZOA1DNoAqpR0OZ32r4Ie0zTUh9WZS9qX89j4KRGB6bPAG6w88y+A0dmmb/2o9FpXVWHr1
o6NWE9K9WFH/hZDfi4nwWG7BmLWmGm3txMlWWqueAnqMQa3bdjd2bUSY11mlMhWHVkQuui4Vsd7h
Xmr7hYC5IEdT/5XWxFK0uvPM3rPSh7TwGX55bPO0HPnNWw3LfskGPPc4WT8IBm9NTdk71Arfjqle
glcJti/rLTRgjPYAvC1hpIelUmzIuVULwviDaYi1ZJj2xTIcu+a6ZjDVp8j/d/QyQ61K3uLoT/iK
ItbSg4g1Oh2nzzW3OtcLE9z9GcYkzAmgustddSpTH9yDXOGEJnGCcvSMGllNW5i6zvPNTxNB5B0Q
QalnLzQ8uHoFMUMiWeYy3voDYc1VhL61TjJaZwe2mFiFnCVlLz9PPE1SgbpYmq91oXtxq7m7daDl
FepcOJKDLH/bDrSYA0/iOwuol3OdsDJLNAeRhTCkPOlwOP7zRcXpbUTeaiZ7kegHpX+Tfpeha9Br
fzhZFOsH99ZHRJmardg8Rmgt2WYpAUqNImXaQ6S3NQKNh3IcjNxzl/nPCtSC1uivIp4bPvoJAGFO
jmoaAerdMhVq5dfOaDaUGZcmdpANeWH6Osy0LOdbKZK9gmPJYSs5cLmyf85Fqjdu33dQZFDVzE0Z
letuvuldvleeF8CBvn1khgw2BFO2HIPHUqzV+34SQQMJdsb45xtc//oF2XhnvPTyFWcYtKMcbivi
Xtwom/vwkWFFxAlAUE0HQDAL1JZ/rYWIDIPesh+KKld+U3PpPUhGqz9w+7nLa1irJjeyFigD+a1U
hRJcoSGTe76x1J80qD18xAHpjH3seDr30KrctuAQADZbOmvpTI0KjVWKtBvvR7o5Mb8ZPigEUIoL
7CRyzNWkc/QdK5xYNHIhClBROE+FUE8lNHJbIkCK8Oj7T9qkF472DioaT/oT99HCf/7jFMsqh3d/
yync95IOPSWrJrKBgoxk7tWAm8Yrz96jYq/a2A7GpTjgrcaAEQjvbrErlAFEeNIGEftVvqC4x0za
MDzQ80K2AmXM/I7ZTq2mbtvFNvN//JALS9ivS1pCHlf3pzDbFcrWr+jTS/Vl8xdLAydlLRru+ZPW
/YUYqenBFoRo3LjDlVfN3PPP+jw2oIfuC7T+02ZXeNmCiryW/xFVQtDZYusOD/8VjuD6/jgWY4ey
yb6suCooLH6UAZDiggT1qUF7FuTxdVAfekweotDkN7ciiOhOoAephUNe21z6aC2riGX/7IZSw1iU
TLg3UmE8dGqYigKxUZDQlJBuYPhmOylRngYm+h/HZOAyc98nY6q65TFPla2Dqgf0virjlsKIXrY2
9DiweWRxCLFaFEdJjypA8qTmvnAvOuZCmr2N3mDe+KWcHLCgqIDSvtMD+ZjIiRsyZcpXho7naRVE
hLnZK27dcrYPbAA1G5OmGmU09ayyUasdZRBjjagQ/ce+JyWc8g6OB0gt04mwBWcK9B96SJFCNhZc
ENUxufdht87S7WllMWZxp9nJv4FeMWOpAlIFhrWep5Kl51n/yg+TLTKbNUZVotBV0PVEP8LEfp9d
vIjygHVLyy0uw59blDK6+v4yEakqfQ8vq0myK3TL+RaPprDJJoEdcdJNIVjVA3x1TZOehlAQ5TBc
k3UarWJ2U6sJX8NuxC899wct5M/l4CKO2UaRzuTXwL5Q32IMY9a4xYZKj3PiDat4w+y2IDT63CVR
FaVqZH2H6nBhwS9cFJ2FIgwTadDB2zH0e9lEIyymI8vVDIT50Ln4HkFtkSMOGxgwxrDwhdWRWGRr
VhXpPbEav5F2bSv8L7d7D+t4Ifu12so++dGwlOSJfnhdpmGjBj/pVdKvKQFI5cbacxztG55sGEtJ
p2jSZnPHqIx+LqyFgox/Z+6MrbLOBqabIH+WBLNWk0PWEa5uZbeeU/PVY6XM59FG2NOcakiUu4D7
EXWMmuwPvCDQKOGnhlVse85shnnr8Jke9XNHR6NiKCfb8JDvP7VEQZAGWHTNrOhiP0i4MNnr/xZD
I3AXaFLGDbRhzAQAd4TavttbAQH/Q2d9DLsy3f/95KRqNeKV5lthhW66GU78aykuN3ozr17m8oKf
p31Wq/n3L0DgU+YPgZJC3yK2Nmy15M3Jo7OJ7r9FkLqSgsKt5jNNKlTiQKwsM+yFKJXRncvsha94
mswqnJQemUSGtXRZgnRtD4ghzfJaQWp5DfNWCClfVj/cPOwaIzEQstjqQnOoSgVMoCj9aXNYKqzM
L2HsgiFR8hmpSikuA44qr4+OEK5GqltM9sJwMJeEotuQB93Gh4OgeBxATr8mIQ57Q3U1BQjtSdmw
gBFgyEt4bRUJJ2VMTCopmMb/myrT9yRYYDuKwxEbbiDSZWDqsVA3qoazDqCshpg9SnKUD6VXOw/0
hsCAPMfQ/bP9CahhWDpYsqvdGQmxrh5JobGKLp/tNU/527D+X0LB9m7rWerDXcFI3aAc6cN/qovv
8PaaXL+0leDqNG0JcmPKobJfBsjFk/tCi7xUSJSJ7fPnkpNOoEdPWJgSXXUR62GY2oVtuKU9VSX5
8GHRQqDjVGpEeqzr0W2ODSti2bxUWzTuiK8rBj7aTzfV7oLZkGTD9eqapGkR/SGmDkmHj4pOLRP3
fULGYNDtFMq1NhUmyBrXPFJcmXL9fhK6XiUq4SfawD0XGzpkbNScnbWTrSLWa+OAmYvn9nqptfKh
nXzmc9qiLUUKBBE5Uz9lIirrbN8aLAuSXxB1RTQhls0v4yMR5L7TUyCSCgYpEQEktec+Iv7/kogh
Nrx5v+NvjSjDIE1LZBt0hlqkOG8nlX5o+k8At67m1HP4mYeYCv0sZc0Mqv2ziLZpGvvZ1ybPdXhK
GeeZDC3XtNBBjDSh3KNehGoS+kEC2rFEkHNiQu0wjVFWhLtpdcfUHwWIgrIP2aR/J3VlGyy/HQgq
ULOVBpwAPGwFi8WYdGUOqI/4vqUWsruw7tLg30rsaNtYmsu32FV8gCxpJvkhmLAlUl2lhzWn1zpm
xtECtGICAUB+CRoKsYbPYo9MZWJN9K9KyDYHMrPpDs1dgCXhZUbcAuLawhPscni9QzNuLQ+QMa3r
dFBGDxZkn5cHlNfWNlwGYXzpWSPHADi2aivj0f+q9d4Znn4UhMVRAI7JOHYutGc3WqTu30FKH/AO
Iha/sgd9A+DoCQ3qG4yTQPq7lDcHaoC5xBaooxIxgytG+jZi/F1HxFn9vOR2eicGAyz4U0Ssu54d
tl8R6cYX6Hhq5zdnmLyS01n95lwlkdTiaj00yf+H8GdZuWNTSnJ98elquNuoP5h2BuRlsfd+M8Yf
byD/hkBplZWr0wXfMjsIYH9gw1gR4FEB1MEvE9pJL42bJO11tDdPb0YuWQexq5bOsFRhP7mDXFbC
tv9luhJ9MSfLkuXzLApd+8tKhOZGgXaKtnB7iIP2MQ5N5gPSD4OlicqQ3QyEHrJgT22olwI1BtGs
T07hejM9hV3ifTljklDhPvGlQpu8d9P6tumB+VLaOj8PCvk9lnQau7oeWbnec60R6fLVWuEXtn4p
ZuZuAEHM1MrjIiyerun+/h1fgTorwH+UWOvPS7XZG3HjkRv4+qM5zRQi0O4qy7l1vWwctLcN4/xj
vIrmn/LBtPmgkI+tQ30qzdBx5laM+ohUp42aPhDNGnWVSlJygedOLCI5XMRJTDXTS58k+kW6odXr
9qKlz6TCqgx0jGVstN60WnaIrfYQ+7k408AIFqFMhtfcgG9HJ7CgdVQz1jqkR6yOjNWROUj9+snm
wddq6Wbh4mGa2xDVRJnSIrwIkMiswUSEWK4DKEssfnRIeK3IWB0ERfopl5WsR3ZyQw7I2yvsAtmq
MC9680hQGTpGTWkA0UsKDnhClanvF9xmz6Iw5eilTELptoVkaCVaFTlG923G0rE+AjIAqKPx1+HK
4uTLapMFL88E/5cQOuGhzww2YRNg4IpLsAOO1bTzGqNjtB1MFQfF89cFLJV2vkWFusAz17rBk2zM
m7LduhFDgpEu0Zd4gK3S7X07h1LxGClK54jRFEgMFYvoC7dDKVUQ8y5IA5JpOt2jSSj6GcX4Aly8
OszNXngDlr8IQINj4Ql64/rZNNt5KBm908wRZd1LMW5e7Ua/jues7FhsYNIuAJkqQLXAAR4PCjD1
YUn6Wm8mOJxUZkYfoKTHkyQszZv9dH8XMNyXURcZ5xmJ10o6xyNLETrhnmEWJzA0LQejvIjgLWzz
rO38k28n8h3GXpR05HbLPldqAvYfDCgwibd2AOvYVN4wZf3NZLsjBUe8k36ZwKZN/Bmc2j7e5FTj
zshjU8NbsLTTUv04vb/vuyrDUXbpYnIZ73K4iXDtS0bIyv9PxzEmrO4kcG262OEN8x/HF8qVYwOZ
kpIC4tGtKeLOwWRs9OE0aJSW3PLMYgOIN2RT1UDdTz7AByYCurp41uAWAf8CwqyhPMnI7nrfH2Yz
8hH6oEqb1Ojw9nqF90irFeCsUPhNrGDu4UD6OMzMMejO2q2zfT9zki8moMFTrg/S1sSS3GY+J2nh
gFoMbv/yCJ2q4PzcDyRZv34asZ3StAXKrYpjmafnsOAud87X0JFDQx5D+pJY3ZfAVkpoZb3P6aCl
MEPjgWCu/28GyJSWg96Kwt60XJ+z61LHs9L1/c7JtSn8l2XIQ7hTn6uZfUB9fLr2eiVhGmTCvzvf
3gZboKK+ad6ryGKGWrxGCUI6ZCFYb5CE8VcF+0FWaIayHv/Wjx4/x2aiXUwi6rXWBig1JlDj8657
covJdk2cJM7XMFw3qN+KSB2vArm7cW0mpjJdG+VSDIBaCZUnAAwCcBqEQwk2tC3anTwbH4+G/QJj
f9Qq3GvolXs6tF2lT1oyHHBzKuR/ypX4nQqo8RlRTMpGp4hR9Q32qv8vBmJ2/dN4xDICuLGBWubC
jlWbzWzzcU9ewi8Dqph6ci+vlER1ZCAV37gmwqSuQiOWe8VCU+1OJ53CfylMUpMqskls/Nylw7rC
xH7rVNxtU910iTvwzltK1qdsBVfonC/YouYVQj0Qlq3NxO1pPYv4YyTddfVALqdJIck4uC+O3oWx
KUlzbCfV/ZaC0mEcEW4zA3sCpfiXobcNu8SGBvXxtiIX+BtSM7lj4OQPXhYPHYeT9PLO/unG+4oN
kN1Z3m3IrpGi166Z7tTB8rFV3g51CxkndRDwYyC4sYcT3paINvdFGMPGkBP3iEcexIGB9Th3WPEb
20VAVA0L9C6mV8JBhnak943vltUTVLW9KH96dfr7mZmSQIS+IbkAFhlvNiz9xr1imvabnqSE6qch
luepn/yyIrzcI1WBbGFfwIiPduZz1vXz3Yw8ZEJnFEbA0wjMJQAVf1OV9D6pKiflQpJwmbiA/ala
/rVXRVWCPwEC33Zm+n/D8FGYiO+Qi3e7RHd9qrlPxONl04pvEkq+i2UhJoCy/5QgyrQEXRBxGuEs
JQRU1kyU2UAOP48JT6LRUt9iEFVZNSEJ3ZzHNzXns+3S5GyZpCWnLWxC2Ftb8CbPD99GvaGlG88i
//YxwSBmGdzRVVQy2o5WSDp9ocRSAo/ienOythPyjhtj7k42OqhZSgf9WgnxEMHJA/JcBMk9bX52
HgC+bjVjjRgk9gQFdvAFl10N8miZ+YAcM6ol3bJTpxiPT6Q5EAaxZPFj754/+OO+BVn6oWC6wa6s
Y47qQHWJxY5dMNaDaAZUIL0/4zBetvr/ZvMyJCgD88qhYKtj05/S+gv8vDhR1p0fWhVwcX3A5Iod
VWn1a7fTaRG2jyaGP4NabvMRoNWwnPbRSP7VLvFbHFpyMVlvjx7toXg2mnQIEPpdALWNFuJJwr0z
icEAiHsNXjzctIVRGpFdxZZ9T7fwn0Lhb1AvxwwEymVrpS5dH+N5hFSBv2rXViEzkoknib/SboK0
pgg9/MzPrDgpNiGhryIQOhSLCe03wIzTg0HNFa/6sr7wbCrzcTDKjCPn1AS72m9K6HcRmP/B5NNr
x08FJVb72HoXK6YlkaFqqZM/X7B/MX3IbXufRGTCIjJq2Lx0O9xL28GBGS8MsxvCZD3Xr18fKvPE
Pb/zPKrBUP5rXcKtlS22xbs/cBRdHHz8LxX3J9fHI3BfRW388N3FnbbfZw9xc8kM4YID8sz3bCI8
geRNwIvPA2pmUEDN0U6Z4kzbWZqtShCekH1sUdjDhcEpbFVMFcGpRkq0fMMRs7n3kXKFRgcPKslS
knn/4gabGztSaOAciLgScfXgSKbX08M/u9vY5Icw65fW3dX45ewJ0CGwIjYLBm6h4IIFURUpDWSb
/QIRtsaHwX/tZj9v/cL/5geCZT4rYZCPNX7sclsv+oh9boOhozbwT/vJDFpjhgf3ygVHdsBWYiRF
h9KZ7mY4M86bd8QiRgelRHNwtbTQCsmeai1ggNtpEXlAGiCh/dJDy2H7b36+DZitAX25S8dsq/H7
YE8ZCyegm4SArJbx4Q606p92pbOrVBHPTjn3RMavxjG1ooCca+FMuyMYXdx06XTY1cVBqWgMnAux
2SPfQvg59QWvifGPXGCKL++gUzOsa3gJkCE9AbuHI42T/eKjU1Ve0uHk64K64Sa8HFayZv4fBora
3c5TT9pM5KJ1o4h1v0zP7TBgFKihoo+IGVCwiHbF1q5EpUrgp/iiQQs6K0ecQePGBeBYvJ52Kkqw
wyJCH60EcG6F96LCbL7Tn8KtS9LVeu1dLQBzN2kkpgodezFVq6BdiBs3g7pnq9Bw4Ec9AyLdIXPU
mDlZ0OfMfCxReE/Tm0eeNwof2mplD68/pD6nfoHDjK8cRkj3oNXSpqhdqczDXyE8CB1TDSqIYObZ
Z3VpfhChT/hozLPSJGfytrC1BG8oMDjD6sYABsNNCK/J7kTFLsLrWzwBTFc4V7YJECjoKMAbO8h8
w0eK1/24/EvXhX9Tek/ynLTBdqzWIEZK0EnR0K6x+36T7wXwwUXBURbvJEU+IA/5+DJ5aMSTHlCp
5aSKCVchRkO2WmzuI9adzW7PlumXeRw3fN1MZTSdlNXbNdRvsGaXMlfciRpw4hyGTH0t0BdZ4bxG
N9TsxDWEncnrzQuOU4YKTKJ+HmYyv8uKmeHKve2xoADoogNdYRw271dpA34ULk41VlI2Oyd1Ru3I
oAt/lrRLvl5rIR/3X9VYIygZo2/NJLWW6gh7oWQTxCr7kVt5IeHNpXcK2/Oiw3Wxi5B7MJb5ZjzV
X4Bjrgnm0eNWByfVEKhPq7moT+3+IGBC+h8Y8tcdMrgL0ehhX6OOXLdt2/0MFHWkxQNcjMwHedkk
txbI2hA3k9R1MdWn3NrQMmR5zOzgYOChzOcLrajbppPUMwUCZxzqNjvuMHr/JnIl7j8XXy+FNWrd
i8w+9w05hG0jKrIONL8xLUPyumOP5BJio74q/0uLgU/yxeNiDtxA6GHzUz+65lOw1XMywzuo8MDL
D27KRZzTM+lNo4oWbRJ/qD1lhAg8pz8i6eq9wRi51UAmKb08H4UidHB8ixgjROi8NdeY0An/crQ2
FCOxOQA0oPurnXNjAsc8goGmvXIMEYFr51WVOQtyetBkfoDaDhj9qqEgTmxBPfaikx15TnhTHCQA
7lYNeFRh1DyfBZJEBRLxM4kXhcaK8UgkicS8e031SIdXPZQP/CMpyX/az2WsXL1L7xuRH2Yh7VAA
9IDveojvzY2EWYsYbwroSvGNFV8D6LqPSE908Qa6iEaq5dmVRi0en+jP9/zuNmj2bJd4sJyrDkyX
TpBB4Mc/pOkZzhHTTMc5s5c39o7bdOT0SCmS0FUCKet5QO6Ism/X0RVJ3mPanhSJW8dpDHrKFhXm
Vf8dHledTvSBgSYVaqdMbjltA8vyTy73sam9UBjwSl19TvTxV4VMYYm/2PUnhZaS89eMyBqvlSer
mAaHwQ8B89vGrDO+jquc+Ovn+yRwfCroKqHBHikW/xdFpvWahuBa4RQchpvpeEnRIh3jh5O+9IvM
rDXcuOUFQwiEpYXFJECJQQGW6/QmLY7J3Th6TyTILWLLz+iu9M5yKZUM/+4s/rulaXO4YZhdZFsQ
Ohq/ZhUtRraq4zOe5hemu9itsVG0uuTZOmPybm9Rju6wfDlEVg+QfNELOXtXnGn04MkhF7MajdQA
NTlQCKSJ7TE8mes2T/k0DjEyaoXDpzAcF8dPS04WcEZGKPXqPQ/sIbBTJlB9EN2ZRPIZcSErfZpV
3aDm7kvJoH9K+xSTJfuf3086fgCmeNmZEgW89jD2MT9NW2rcctyTy1dnZHIiP1FWA2ZzcqbE0bYD
LdCRml/+fPqW9AhWoSTtLCg0zBaWxBQlwR5xEZB5sJwoLGqWq6jBlOWKlqZNSEPsOpLEGpQtFFED
2AV1VrlMsNUSgwTWCpUhrKMENcNwVEEjE9sLxY4pIHIsnSznKJoMVxzSQ/BCD70VDfodmGezs1IH
8fa4YpAvWEwLuEVc+MdD3Pc8tnHh5DM0pULjwryazH6rMJrWOgGSyMp5thM1IbZijDYRFAGPwpgb
wEcS88VSg4fSuXUNPlGKZGghR0cu+dg5ji1SPiUJW7pF/2EHa3Wdq3t8tPAGvpzBty2wRWfZ/7Qg
i6NIE/VbYTNcq12AqpXZZnRHRmV6i0DPwcPwLQGh0wtk/vO9k3XEI3FqwWmhaPT1YetgSOa9/IFA
G1jn0KXzl3HVZCrXW0HUo5yBbpJgxoeAw4JlwfIkO0BCQt/MD5HBvOhdxTMIkAeUyH8YFnl08h1K
0impL54bbkaFvIrJrOsg0nDH7HC7ca+r88ro5fBzR8S/zEwidV7Dab5DG2ymcTntHWG8Ij1Mhdov
GRwlz6XflNEekayKTucQM6GSnvByez5SQs8yxZ83hQ/nqte3d3I4KCk2HqwlM2AjMlrts9XZw5/l
H+5iF1stsUtbLAkfCHZ/qjueafbuhqR+VOmVPulbRCsQmiEdU0PkEUjlNNgL2LIKnpZYBbgOwl4Q
8ACov71zIOW/U+VB4n5rfOJ50MNpQaN74Ks+FNQaH+YOsIbI+K+h3CLvnV2IDKWxfMbACCze3l18
YO/2PF+08rod1HG1liilM1reDQrCs0xrIiBJROXQ2nJQOdV3bu7NWtqek/vCneh3NE+LnE0oPqmx
BViR9gx0+37wF4WklZ55Ti2G0bEhfp1/FRWbCAcVyzLn2EoQhmoYJiC7/jC87R1k3WrataCLNvDN
R6seaNxjXoTO5auI6uye5D/CX1DaH3/Ux5Typ1xUWciV3/eNMk03e+0ZkDfd9xxzyHWfbpUjZja3
0yj4Nu+syB378sa/oAjFU1zPddrSLCDflOfceMqCH7I8X03j1m6r2LM95byBjWfgVWXHTIzFpDXx
B4H8BOtP06owTG7w5RIZftlNZTyvT+qe5Ua7FmytlqL0qsUkFSCJJwZj7jhgnQ+brTq19KNBwChg
d/0/3QDPS3d6zOxo5Vni5tO58H+dE7hrFJqUl1uM2yc9f8g3ISW+lIe5mgjaTGBObB0trSm0mqUg
Mi96RITHk7tHGLcesSJEOMdlU1Gp9qKN+18YljfvYjkKTn3NvBeyICSflpDXdFsS+DTmBzVxoekr
tl16GN5dEqrSlQ7myHdCHKUdcwOx5DvF+rlLb2F42wasbC/sHInWkscdvCCAIHZMrGScBMYz/aLn
iINDAWMQNQdtkqXL+H/5tX7iZdg3E3iDt+rm0DInOrbr5b4H/5u4JarqrZzwlPkEko3d/WLrbPdk
UodE4yWUnJbflZ5owFQkFi5xgPtM90t64aPQeKW9HcmST/RHEQceV2mDZu4vFqooJQy1pMLmJKMr
e0jm/oBCZ3y6BtqUgplpXkeF8W7IQJcVe64c1eyco0OT4NwmmExJvr/Q8Z7n1ZtngsPjM6u9tZ8R
TadKiddECl+PbjC78L63Ioqg3xYkQP0H/ycg5NPjpy7zs1PHaVufyG5AT/ew0Yg1w0IydImYMhW+
AShLicHaVAbPbR8Xroc5ODUra82g0YulUMf44T1SXZsLn5zY6EsqBjCfEF2OCjZetmapnNMlEaxk
vEpbEZfZo20ex6P4nwoJSgpANoS5bSyuj3l0AoioAnwuCWmuKno+vjta8rlx3aSfOdiBwhhr8XEx
1fykyp9TzvLFhjq5hgojlQxMl0KxHHWNbYn9H3aqBnPTmHf5bSDUltqknKwFjqRWSGkBw1bM8qQk
AViLJpdv5WuP6xagj2vAx4je4U6FazGkgMHm7SYsTzqyKEtOjR0JSu/qEhngbax9TGtS8HuyiI29
okPAfvgmOy13iiwPk+InayATa9RRqZZOEgQB677lUa3yp85bd0WOBMucVQckJohzTDh/pFj8nbK1
UYJIqMsZH/UNEw6dZ9U82Nr297VorrJltRGblXfLXNUFpPgRVOv+8a+nq8DstAU1PbOMkxkK/MiZ
J+IsBxONt0S5YX56FAjK08TDb53rqmrAPvkO5RHq2mhdbczcXUofd0sRW7T+cI81aq3fxzmj4OXp
AxNwdYZTQtybAmBXK9zY0D3S13m3HT/63Pbi4rDqQGtf/yTTw/ls5gU9sjzT2AyMCnHNwip8lXMy
sOPdWOx+ZRQIIXNgVM/qSz2fXQQaUYpvUeXm3MAHXWfPkt+9xfpEr0WuHGdX2ycU9ZAvr0uKEYq1
E+Tzcznelztk7YVbmLdf0jT8CCi4jXogEkK5HdS0eZQE6BgwFPN+VoCm5yLVTnWS4Mh1e/Zy3UyE
T5ejRiMta8aoimeuN3ng/thvpT3VbZqz0gG21TrIjLQyO03k9Dy50cV/Yq0eO8iFmebvzfH23SKt
zf/1OVuydHxEUWVqSR430GYVZdA603uzR1JaPgc3B1JKaVwUuOroanBRteJ1b5Qm2QcTkHPGc9M6
jflS6mpoQIMiRQA9yYWeGYfhlOP6WKse0n+10XeWn+z4XVaxvnsSqrBreVq7YRq+obWfDx7GXrnM
aKO0xyuQfjkJbigo+8hgZFG4tZYuXMGzmaD+WHqqUAjEehJRj/5oXryjnu24lSc1voxK/TAUeJzJ
iCiGV08TY1Er8n+KoZC1Eeinb5VKySUQtzbeTkV5UrS03jLvopu5TxkAO6lnvYec5pmq7wqtukx2
rXGo9XfGTl9gTc4TbiufyH0arZjgJ31mcRrdpcBkDGxOgzKDlnNHGL5R3YmyAqewa5YfSYQ7MAHv
QSEb8yYi1b0CyxiAC5Se8lklOAI7ggHhLmbbRr0bS17e9aXcvRk8lqycKHQphwGjqyJ11kibhGbz
56h9TArUFx9QRd2j3kAvXfWEBTnK8asbnENiRq4vAQm9xPiPs6DQ4Q5K+IqFthOyVr8j8l9sIyn6
COeH/H52w2muzRrz7BYpQ1J4CVXLzEGD9uer00OUUmOXYONQqLEm0+VW7M2+WlCSq3YENooojn7v
s51pkOix9cEkearUq8LI7O8xI4NV5w15dFCxvdPoguSll8BqtkCZNixYNH+TvvNizpT130AyPlbE
L3J0Iiprmi9bnF+R9p4bwraA603ivEHTl9JqmVpefHwwYsnYivwPCmcLm1MetvmN8ADXtGNB+16S
WbWJY0xZ62M3lybQmb3yB+2eiRw0Upysxsn35eEW5BYLMtoyTpRQBD+PTWIyWCpZxyu2SJFDVLSF
CqUO8I5XxEC7jmSfHBV8mJ8BLgbwjmEgCPJ1XiH9nh7Vre2yggls+a8C2vCbjK7NJuPj/EMEBWif
C6i21dVYVtMzQc7pSDgnKRSpPbf5p7O0/1yaFQENMKQvg9+dIOtLeQvqMrsXGkI9Vp1vbp/vNlOO
q3cAYKuwIGzQQ19zXIGzPMC+dFRLvDfCU0aMISXu75uSD6o4eIWUpomUKfnlSOiSd3XuOEnGp2PS
2dxfVHEmv/Jc2b+ttp6iVM0BTwuojpllF1W24h9A3qvEND6+obDU4L6R8hdzgUvP9ma3wp9+nTBH
hh4hDX2N5M9Hc4YW6ct+MSH+YGBiXQW+sNi5Fu0I+Xv6MA4O5+RhkwzKIOJ5TYE/sNHqmfRxRMgA
eAKMLzR4NoVU27GPZwuWpB5qo0vOANnIf3xL8M6u3m5w/msCnOE4ukyaGdQN5HTyfLftXUgVWsXl
PB1fnEMtm0nGrwrdJw/ez7gjiy8gpV/d8i7vsRjAys18CwqG7K6ZhejImLV9wDdE+C+ilyHM0iPN
aTByxQwxXXaot1zYNg7/hVb0gwaT5HPsYpeTb1zTrXK+dBcAIeAhHCn06q2b7SRoUMFyAzNsia3V
w04JXiEZ3L0CDcOUkfEYc/vxjiL+GigRLCzuBOhTNejFkPUFeFoi+s+03pZDcWehqFgeHJOVIaWO
Lf687xwu8PSuV86o88z0qSJuNhskF4b/J1GUmf4zso2ULXa2K41cupkijoJSrVn0JvbSMNnUjf+/
OoqdL+wrv8QTYwPsy7G7B4rOn4KA5H608AdiCoDWPvPXp1hPWfnHFeVPKYWdZYEthGZ4bJOh/hel
7nnDrz5sr3VxQBKS0t8Xl56z71F+iLP2j8fA/oDD52QAw8qSQSKkL+xjWqjT62Vd2pyz3gsBp+k5
RLoFf7JfyMolRl1vKPRAkWriTlsVbrKgfRP/Z8WPGo/Sh/kAg8eYgdqviT0JnBgZRa0DFIx+56pX
LEvyAWm79b56TSfVR0rkoN+oUYFMZLJXbdrLqX1hULsgeyCSb2ZJ5RJ3vhHTpnSj2dQN0yE6rX1n
/DH8EnQzJV146WD/+dtKD+C9DEYzn5ihjvuDdBIz6CjnI1bemQp7pQou3X/RQTDvTY3Vc7jHQyp9
46vNa5QSkbSEp2yAer9O5joftBHgeaERMP8mEfVeE1b36wxjlkH1O8RXSuWxpUgJmMR/P69epYLX
c4eovf9t+MvC5kPwwCyH1mYv53irOpUTSbgIvwIhWMEDiBjC0Z8rYOOHgiCjZLgZujxl6swb2Xjz
HLTE1/xm+9y5t9xonsGOV3s0+05o8b1FzapsbyBx/hvXnTuVKEtthzLUHec6+HMQsOVB3sSvp351
H2UcD7rpmonH5xAZn14emONpcDD5OItm14ZXEtZBgrtDoBPGAjGPyVbc1lNPh12TnrpEPDqVdEy4
ju+A7nSDDRmRbU2PvuQnuZ/ck0mMwVGHshh91dAMy4YPKZPSKDur4LG6qQHnHfgObMD/dyjVOqyR
BVjBbhNIfmbMTCfry09FWFfyga5yUikPoqde1Nyn6EawR9bWgxJU9Qa0A4qS8dyD0q5j4tJzQ5AT
pQFG+gZZi8HF2wCz6PBzoFmRoqrd1fDh+oNfDTuqDomkvrYK4u1Zo562UWVSKoJCVnLWTHvbioso
RPpe5Num+ZMqFhk4l6uTgi9KxziEDPbLU45J0eDmum3osVJDfMlSX6eVrrlHL9q1hPuixkLeQjiP
/Brfzl9UmKn25yY16yQgehaoEuxB3QQaUyADxNsmYmKEwo8oXZb1mPT0rNnalmwOvZlOTCiNqNmP
XQOjMGW8JhJvl6G3NmTa4KsULrugC4Tp/OqMnJxtTn4f/YBBLtQTV6xK0d9xtjoO5fXx+1ou/oTA
5aOSskYS+5rlUvPPvnsxf8OTzewq+1JRKdF17hViVsDr0J27BOTGmuF54iZJBtblDR5NReHaPL8m
Ewu6m1Za4mRhFcoQ0E+/l4fmdvgVVMtNEjS0L0AQ9/ryd1sjk7RprD7i+3ni8kK9S3ZR2DuU2Jwx
6XRyMPxWJPNgJ3egiWyx6XaHy7cocjCLVl/GeevPv2rWezYLPWaAccgOHCqcM9i/FjMdkjhFdDSq
d6CszrPpxRbNcQF83pdK3cq+97R5zrYpHbgWQvhxVCYLK1dvhbqqWiYOE/ZEwf9sc4RvNouFe7tG
2GPPAX77wW6se5G14eGnnthbAFkDbYXz5JQslmVbKpE+i9CD+R47w3sm0MT8iObPFYaj+Brz2Oct
1kQPk9GbGk8Y+0swssyt1pZE95kPlfKLDSOgH3I2MfbHqDllQRxwZmU2uQimmjqMeAwJl918qKzR
GDzuGwIg9FpVqELuwmlA0AICGP2nMomnMLdGQnVexQNkYeBjcV+Nuuln0yOJSOZzei6ogPXka3SO
Y1JZjPMBiz2oVNcTRe+U6RXcfMTgU1MI22fhWDMCsD2R5jZRA/5OUivw8GJmx7UKsXt3VjlAwye4
Vu5Q+2rHx0+s8MMp+UD7/I48wGkxrpsuizjNTxRFnknb4FVvki91Tma9EDXgymT7LM7REq9PzP4c
dHCX+bT1omsF+DImyOd1GxQZatjrJAukrXBNG08b313o2nuc0sY44AfFmfaExWhQn7TNbETsWX9G
HuV99j8fFFB7/1FBX4ibrjvD1vaBbBRceQGDNYpe38Hb41IkX2VYog+GOHiCo9JQNoVZsWwedKqP
hnWaaTd7hCDQyaPwNlBKYgZ0ib4eHICOALb5ISpKxkV/gOs8vGDnbdKsSEVdy/MdYpT8HFVJUU/W
BMfu9xD2LLgSsowcNNNBAxvogJmAjSgzzYNhAXRe6XLHK+btFjOwRbq/YplRYaV/ojHdlox2syRL
Fj7PFe8IjpJJMVkAoUjcHgfH8nQgHTDdGysAwOA5Az37PpEnWSDagK+KNMfd/HrR+Qp0rkzD0QLC
1xww/Cv2YQzJRPW12owzFb0i1FkChJLb/tHHXKnyV3VO0i0tyQadhErAZQWSWwU3ivECe//CbFFu
zR6MBmq80oCUdo9oreujLviGE8ECmLuOKhgW0SCo6ON0ihkIfkY0S+McQIxs4o6+gGD6tju8ldmT
kd08iEOoYObQPkEXzvz/wojcFMEl+Ms8DS1cV9emljcsMpze5kC7UA1sAVvEZT3ztNrife2vbrJS
/yRXLImahsxJh8sUKlSrHKsKiyOnYrm5O08UEm3ZvKJqUGZ47FylP0UPvTy1C+D+fwlwyf9o4BEi
KpupyN/vR6AoP8C7JV4/ytFnxpw8LbDb0VplPkpgCbVxxeo9wEb3FzWrUVaoMf1z5ailCNQbkUfH
uiwMRQTo88+pAengqaQS0ZE/1Fl/mKqPH0xvc4z8fPZ5MfAH2klLcT2a811KKH7fCCSODr1yewn9
QRRv8oYlaiJolKLlTmH9jBXxSfU8PgNX6l//16ZXpQ+Z/Rj2dwk5x3EhqhGVT6ia15JAWpRq1AVc
zZvgTOhzssfhmBR8aIOryBqifFCaElGMC9eRfRxDgJMZ5545hrZwo6C+/BGvEtkKFsMv7jZLKBFQ
neFXZfcFIaEGNZfrg8oMl/pS+JKo0VCBi4xKnwlCQ100SkNMgbnoQY0w7dZe0HhjZVvWhIXo6zqX
x6CmxL4nFOlmQYpcDgpdPkx4ornX7/XE2n3OvOwuQ7U00jbSnhPRVlOmNQ8G7vc1p1z8bGkTEs+n
J+VLYteGV5A6XSByS0vkqNSP1p786/i0qvhx4AD/IfJQF/PEI0u+cfHNbNJTv9ro5dHv3gwEAgsB
WdPs/GGAZ55H2UKK0QVb6943LgMx07Em4PyVMeWkT4dQnDeQsC+dTYRlU5G3yY0mtdJAKsq+Jkyi
tvtsOw2kOnTUxzOpBhG4BRm1pU0w9ykp42KIl1tO7xt3y//VeO/++U2BabhH+7u7KJrnt0TGyK5c
jgiK/2XLiqH8KDDrG+Uj6rk3eWavQjrrl5nzw5T2f99vuR1uIN+i8UE3LTcaTYrAEH0v37JX4xeG
m9IM64sXWnw7a1rI54wno7NTTshO0eV2fwfFITWPjJv9snMrLjrlolC0hcrbFwpjEXG736XN2qI3
ZeFgWSC8NXdmgj5NEAoBtXeZCS77YU3WJ0rz045K/sPLDokbuaeHqY2imgN/1q6hdKxMVsce99co
r9eEz+4P9MXb/4IyQaOs93JZLvegUYmP1MN48h83BNOOHhCvxExz5wLdmUsX0EADcdFDw/7NxEzO
MdQmqUPg+Wy3IzbOswMnFGbheyBzPe8/kCeZPy3jqHn7sIU7KibmS0NBswAQ7MdtgzUg61vrggB7
zc+sbNQyhk8f6V0F2AQljGyLGjhYL3vlcQkrKl7ymp9eDZ6cHJujJWcD3rwDazUtiendT7LDCB+l
TxbvFdlatdmItzHKsWgeQ8Fzt4h9xMfsBrKZaZs8/NnbTXu2Qc5EgQv5qEgnpBvqFol8O0UxMI/A
GyyszMxvm04vDtgtxXWG66xyP5TCOcImzDtKzrDURiuaWmFVC/VDl/5E3Eyx0zDpyvk2gl+DD568
iwxY9HTDHiOxhvMKnSwkajeRqAAqiD69lMyWQSv72ikTnfu2+AteGjEw7qgAf9cOu/QC2e2Hapwv
QmieVTqAziFeCLruobnqwQUeTFeIjiCJzyvsgdqvarP/6o8Eh+7Ef6j1/1Kuww2OjWOwVukMqfCR
MiUc045gqmHLClXjQTPhu9E/8aSvp0fp33agcZpfH3aZNjZ6l6yl5h6M/7MNC9jzcOB3Y2mdK/x1
Zndc/0WfEnC0e+ygzITDFfkoXY9gPCcaUzcgJ+V61b70OiPioNeJIQ74uKFc5QXuGwGhY4VssCs4
YHiljaKXEncYv3Eczrv05yBQnJtB0EHafcqx259RNcYTL11qvyP2Wv36SghieZhGIrZQ40E9oW1Q
Hz2l7LU7HuG17kacdLYgad+13TSfWsl1rnXZmc4Fp3aDtqdt6Nrf0F6X6M2i/TPqEMw+LR8J+4Hn
jrYzVdBLniA9qPxLIrVP7XRo/Qs5oSlaunJDIPzEluQkvf66QERgruzJcfJwAYO/SvB9J3csoieF
+PWU4cdN4AJT2a4vtBFi3h2BXeIgO7tpE/DQS7FcMPbgPNnU84eNupmYnOx/XsFxA6wrrZolbUHI
oKFix20OlVtnyjNGfkkx863nieZLsIUDXgohpOp8/zbW6Iek0i9tZQ9ZkJQLsptSHXJXrYNQoS/h
NRavC9JGvyoA2oDZstx8hw+R4HUf3QxCke2Gkx9mlpHeVWYd5MfJreRKjzy9OHq0WQSWF/0PbW4m
FIrDIb/gmqXptm4lUzKNVXgSGixbkm/0tAZezvw2erQxlu4tDjEte05n1SvmhJZbwpMVREAkNqmS
mikXqd5LMMfxwmtxnhVWLXZLoaj51nz0rPQvdekCkpeN8ywqvyKtccMQhjnSHUhR1WRNkn2HXeUX
aKjAGcLrskismvmBUAMUVVHej0U7L66n4OrVvpXbjCwNSkP3IZZ7/OYoqxJ3fI6Gqp3OIEa9p9ej
zWrSA8RLZzImFx6RSjHD1QoIkEvIujcgLwQh3BO172qEAn8Id3auqooNsXuO6kPS852fzaQuadAl
FEapaxtQxr0LVOsr8YZhcETyhsu6xNKAlT1MpcIcrVCVjS8PM41Yw8UbOS7KHK26RknwbqWN9/vH
hi1hlqdas/Qz93Foxz7n+0NVLczKD/EYWRmC5awSyQNRyZF6h05LpPZaxVhStJCYomZNIUdQbm36
YI7ahmz6eeH0WePStsFHhjq0KHLN8SXodppP9jj9x5HHLIsCZxMxTUmqRiCTV9zUeTRXCl6udndg
+dlDlj75rYFlhAykEINJezwLAyH6pvysBpEMBblFsOkyn9vzGXSfdi6Pcmao6Tne5zwxJ1HJPOci
bxN2nPAyuGL3lhUZ3Q+OqE2iHWGXt8hpR3M6nNtV2Q6KZJvqZj1OBJQBNJ2U11CgI+6SjGHTYld0
iGF7bML/XecgZVjLig4szUo5FWV06rapQlioCgipAhyp4mS56uVFs3ikFm18YRS8kFInfyoP2tjd
7Ob410haBCnrdEpMJETM5DqyxfhsR0dOhkIDcl5P0IMukKYHWZNaG40HhkUCe0UB5xfgTc1o3c13
m+BKwwWX2uobtS22awWflbMJWPVKtcvvQ6ZdmmYEFs3dOKjy6fVjYGMa8onKKsECU0yguIZ7UY6F
7jQt6gUS3gVJe1ZF7DXKp4anliKk1GAFLRxSdcaNRByC47e05atC5bxLSDmXOlVSKWEiHyYBshtB
ZydzisKrttjFE1ITpj+3xx+PbdVvb0Pp3PsgT6UmAzFSr71BvjtjNwGumYgcM1HhoB69JknezhwK
ze6LSRLhYZW0DuLlzs7XwawubzZCGABuGoRi+lpC2eXiYj0kwyBKn8gQiNFrprsShO7jJebtMQGp
RKABZYxb5yj+7QcnJnsysfSgiJO97q4cLarUVUXxYlnU5FKrOcosFbak1CxvnRbNa+OdjXp7Ejs4
KFhnuv1tPjD7JSjKKzJPv4S55mm9MncaLDgMoYYdAAI12Y9b648K1vLPwKRQgJrdhHxgW+cHlaFH
6DhWuCwYwDSMiGdUWXgkkZWU7EiAllbFwZQe8dQZ36Zn0rmi1IXbc4Lk4HdUQwfWt5jdnsS1ITBN
v+hW64igWjLe0hNcnFjsLtr17FxJLqy1CZM1Q+G/W8mEk/emrvtv+fh0zP1gqzKh6DVjHUzF1IUl
AkW3l6P+w/2Y9WWfoeNmK8HSzHjmghp/GUuVV5sourOS3sms5oe5E7Ylry1ZUFV1/4d0c4VPxnd/
QOqoZFPHGbiEvp5/XyoYNjkIbFHnxhiFvkOuSsb0atfPaGoDK9OgZ6iBYg7KhkxSj7m/xfToew4U
FXgZx759JN3RIPRi4kBlmS5NVVApwFUr4oWLxy6i1dDjoK+EMESB5TcxMJ6QX4QBZ0e1/Lm59HUn
xA0iuuMmGFKh2wUvhNZjfHdmaiPmjSEIBnE4BFwns5kLPEzkzz0AjYshd6RErIFn9lHyHM5wCoDi
ZcFc3EZsuQ+vApWb+Xe7eXGijisM2wgU846BEzlGPrfrB4qujF8JuFqsilofmiZiSX41eLmLRdus
M9u21o6mg9Qu5FDZYBbNRU6op2VXRhzFnhaha429Q7jkxK9UHDDogW1bp80Bs9Ybojy6nGCyHXdE
Q+x6BExxC60e7aQzZsRd1nV9RCuFek8Q+gaHTW76zee0GMvO3KckvjpoaQ0uj93YzQRuG2YA182f
VXnyZHveBfJ5zzpiUTeWHsQvtj8Zsv985cKMjCm52p6WRxepAlRArKEGtTlSPXrH7UZJppCmrBCa
5bC2n9H+jkImE6zUk0ql6YUc0Ybr3hHpgnCP8mDBGwhdQhRvQ2JMUx4SOipqfbCwHeL7Ja2bJX7H
m/ShjxwHhh9RhhXmq3ztlLUIjlf5manew9tlT0D27swrujywocfrKemCrNrM2c6q642Z/YhAj4cL
nhqOuisG7SXWTvoFHhfe1xVIhs3XkjZOWCDld2HWlXgN1JMOTWfw9ln9xxEkeeN+1eSHE2FMzQNb
QcZduZplu4iC57EXk3TpGVrmZIFfXmduYDnk0yIzst3bWHgsJ/++az3UU/f/dcURbaEug37BDDrc
Nfx7vcgVOT2QT9FiDVarLRdya2kaC0Jog8x2h5Hh4jOCvnGbQ9pb8SUoIQECbj2LbVl5ccMqxGpe
aNDJm3K3LiIJ3dnQiAfMjSPb4Q7qXL9LpG0OUJlOgi+oslPALjvDw8V/NxSmASHRSHYc5CfBIgy3
TEr7WOqQXtxORKdVFTwGINPPEKLeaqnfrwfruJ8Q1gI5hkzpoe2jacVMFveNkpFnIZDnpqi3jU2X
EBz4DLGgIzSmWHWeAaaSmOGaQVX9nWfLJ5UIoZJr8XWm2EaXxXSQGBm3N1aHGB8bT4Z6/eU/hz6N
vxm5x/PifYru3tOqECRVlVpz9/1nGpCjGZnOBqe8IOrGKGkFO7gmi/1qk1g+WBmjbC7LSV8byM8X
di+e4WTyvNCN2ThxuOMXxQrKzOJ3TbIi7yJYun4HjLj/2r58X+KO7RSwMp7XwbFmn0U962XO7QIL
IU1aLfVITR/yBkzlAUqJj2acjXBda1h26iXV+ZVUvgEWXDfcYhlLzpat121xoRrIjxft9K+7MQPu
zQaIZ9fXJgVsSYVTmG1vLt2D+i2kG5gtJ4nb7MZOMBRxzxFT3FAOg+hYfZJ0rl1BffPUmeHsNSM3
crYNW1n7XFnk3GGFTGupL61R15yiVkqEGCEdYfL0k+sAMi4Q1J0nUO5+dFzt9Teb7f/zzHGeHKqM
8nF8T/Pva0q62+cS1eUnm1GgB0o+bsu3LM689fDskPtc7rDuZeWYuP9i8A0R7L9FJlEXN7LOXO9Z
sO7NZzRV6p43QTSrpZkxxC9yERxvXiN3y+d9y3xhmNslTjOIepN8A6rmX8pk6wZlNEh+2gLuJVGP
DfEf9G1J8T7ovfKVZKPwVFXtX9BSirr0rRcyZ0kW12qKOhQ6uwJXABaZzGTIUDNp/bTyME8k0wpy
O2jlSKL+Vfgs688wSBndFNugb62onI8x5J+Yfr+NQIN9wjqef4Ov4YJEjZT7X+TzUGAKQCrT62IG
uJrdZ9k1ofe6pMuefq/Df7ZFsRBThbJJVtuQ6K/VXDZbu2NS2N+F7Hf66cOw6AkzqAmcwWBMwp+E
WO3mcvu7OypqIDUDJbAtzOVYpGNg9P+7FIkaWVgwYEw1K/YB/W6CU21m3Pt0gK5EXIHsKblaRoUJ
1dgQwA/b9Zc0MdeiAXOuMKr3FH62rLy+Z8LBVIinZw3FqnXnGo6CQh5tRJHcsFa9InM+EzLBNryS
NX9LzYfDAJwc33LKRkkhXyarVG1MN9BmPq3ZSnKHa0bw+wgooNOkJ/+HP33lhL/MWp8hgD49hsGD
5fbMmBis4hyOO3EjLiNLIFJrsdYT53puDon8axDVtF4KgvddJcQ6q46nZzhPXgmz/HyStmNoI+F3
a/MBKbkN9Q1V32j7xoRfoHnFECrkOr6ZZyEn/P43tcZtrtr1rd8efbtVLXSbRgEyR0LQlC4BNy91
Fqpjjrk3WWpy0zZ6+bDhAVWGx1d7b1e+DKJhOFwLRxEvK8ijpvOPphaSu/NoN5NR8UnJpWXY1CEM
vCO90LbdTB5nKoFDZt7hFgSmovMlTrDV+9NiY2QlDuvkOi0E8drA/yWuF1uhRFOO62q3g0U80Bsx
1deaXtU0xwwr3E2U4inMPozY/+eUflDR1aq+YwxIyaprSBgpC7x3tztqsBZXKxFJhkR66k2ULHdP
Ysf8gFf9MrktwOjJmD4MT6Mz1lR3Pa06OHVBqKgMqF5AEdvipzOk6KbIjcKFMtCRJh0HcKeriDwK
ETg3Rfzfe5Ov26YFIBJM8ZZHSxVDe87FfpykcERIWstzy+TNtqI+mlLZWspl2kPqE1zlvVlwKwOf
3EVnBneQbB1kzsUMKpKhOemCBA6RSjFfzwISmgTCKBQWOhnww4I0eiItsU3/kERvYcJFm+ZJ1kFk
kGvj8FUmVjIlz7rHhOswXYsDS33C/Lh8+s/WfHJCN+V6Fx2/dGx9fPCpWeV3eVGe6AsBoO3Kre9X
CJbofcUxmcPpy6PRJJCeWKCBsx7+y8N0Q+8dDQKpzGRBSh/kOdMh9PjFg0/OS6CrSjDA8JV4NUCP
wSJriK5UR1cFt/KAR78fvpuvIopNaMAGZPPZ70/TmWh5wge1dhVwAsCDXVuvhhW1BYaCNySInS/A
oX9M+40jEdZoQPZXgvAL9QjYAyvt0RqFB7JeuAamC4/0crfKWGA5Bfh6mCHQ
`protect end_protected

