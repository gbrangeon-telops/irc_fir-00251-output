

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XHCjR0nUvMBgM1clzO9mSr8YEx9qhDtoXdaphp+J1JlsC9lSFtsV1/eTy/jaNsyBimTHmHB4CLra
VqfCr1I3uA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ebEJK3bmI2t+WsBGbhWIt2XB+F+QW56z7Xo7/vGiNjxPbaq48cjkY2KIIwhppzuYFDUdRDxp9Iva
RlWujqNPGUrxJ1F5Pa0zN6dEMkhKPrWWxZpAFto5e5cB6DM88tJus2O1hLy9PRfKWKn8u2fBqIhs
zvXwIEX3Rz7kU3GI+Wg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oZLpbXnbPC0EfiuqzOyPqmT4FdlvB20VtdO3P1fZux3uAWynrmGeEUk81RKG8dIjeHdSPnugG+6c
jKeGIJZZbH6MRScqnz2QBuupQkeYWE+dCLOq6/P5LV7F5481QZZ3bx28u0vHGlRYhLiMW8KnJ8Xs
JLZ2IP5YULE4cFTCCV3WAM+IdulnwSP3p8oyM0uQffeAJkOTKR9dl0lslKFBplzuTZ7EnXSmYYXA
x4iYEfwbmUZvdla6dJXCCjtKnKqL5vI4L1nHOaep2f0bW/K78py/TJVV+vsvE7+Fi81aNwDFBE3d
V+IzN5VNKD8wM+OpLL9AD+xsAbJ5JCLz2sqFWg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YaruXmtmo/2yQOaZLp6UQc/TTak5F2uchK3/c4SsORqNnQQMwFmjpORZM2++MrgqzkHH5KHH+0SE
PP+ha/JFKIuufLvaAIVDYgMKSDFaxIIvD/8aIAhw7TgTE10+TXTruuPFiw9U65VaBnD/nSEGkP+6
2M+aqBTG/2UNkEELi0I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SWJkuOmi8gVneMbAS0rfK4gI+24fr/0jQv+b5sUWbuvKyCco423EdTDwW7ROH+M/MaGP2QTzNz1B
sh1p0mypy290KKaGmvaZfJU7NOmSNGAsA7Eq3zQGPHDW45/4GXnri5xLLNnybO7r0Ndv34V/fxH0
f64f4NRroCys3EmRDJeCh0D+WDA98E/EHP+OtfmYOGeO+CDzxS2m3FIcGKs7pkeR5dgt+S6srqxz
96yb5/UwV2cpnC9ULYZHZVQa9WYc/XM+Dk71YUYpaEFd7osc9zT0azChQq+XAkJsqukhufRg3dQK
YVPZotO8blEly5GYlPFGnRW13eEh9DRYsb0pSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13296)
`protect data_block
zQrCc9SxNFAM6oP3g3w5kGzDjJIwesXKvkxT4jontLrfnTYD73X2hGftI+uI8G9M0Hc6T/mifyS7
1w3bMRTq7utQcpavu7Bb2uq6VVj11wvv1Z/5cQ1sASnY54DXxNUPSJ5FL3lxR6YYNJGwNdRfDpDC
DlbMdgjlu/G+eZU3wnSNEqsCVVv+Pophp+1CeKOpixs1e1uVNqaHuCBM32vWXKlk1cWcfLSbCfBq
H+gy4bwOPkLwT84kF2KY6FP7mxnoqmaZn1n2Vy/VqgOCE7K7+/e7+BO9WM46H9xW1h9viJtSQvN0
FYuA7S/jlEbnrEG6q6HKv87Ivjd12r+5+a2J+nvfTrcZEjZXdgeQd9ey8jFr43RQOXn7LwqFYrUc
0V5cN3QLMxGZCnCX8VbgZa4xerRyqCBKk+VMdER4eD1Vyr3oQJawyjWHJmWqNLOMOMkEBvS8TeOw
GHxrIZCiwbuiqlVueVVnvIuDwdSZU7Px5ullyQaMNzdY2hxmX6u1+3SZkoMEIRy1onXxBw65mhXw
aMFa2Q0x/sEvl+Po2K6wfo6tfuGvfNRwvL1o8aasXr1g46srxZZ6Wck0b2gK2lVaO/LOY0aDeMGq
apcr2s09qGh0HR2DtVFksRVX+O+egkxcYgOgPimXIHuaOIhXqds1zWSEPBwr5fHELo+4YK9k4TLe
WfRHg8ryx9rYmZdSZz/fuMerOakdXbD7H4R7Hf4E/Ls0x9kg5ZTkfuDKb3gTu5/q4TP4IqcHoaU9
VmEVfpS2zaah32VGK8pJ87brQZwbeqe2N0ZLi6TumyDWVTVvbbeD11XB98H2rFN5KSaBKpwhl3wt
liyR0gQyXMHJ0q2E0R+vZT9roZJQ5J8U8lmU4YnQuyXupQs20wcT1Ad1mgUxfC3lYbjI9DrG++NL
p7cJxR+/mr3+bwrgLf2lLoLFxRDluqFtjM/957+Fze9nM7CDUGFyjeJxmR5POcn4WK6SPXkJ4MUf
UtcraqanBvVHya4TlzdA5jRrKufCmpQ98SMx6uCVzdrmGkMyWsaCQlJIuQnw2mEFIgdzkxuiQAfR
WI4AI6VCU+wm4vlS75xZeuRfoYTOrLwzX6it55eahI0/m9ND1PJfaxBxcjIk9EEzZ+IUM6TjqsW3
QJOr97KTmsTpWmuLzxsNxzez5cUg8zQnQVqN7CF07ywDvoaS3cHhkpiHEy6DO73K+vZDRgAUnIjh
2szPxcwKf5LDxQF9XtKziqJBbQfxjxpvUx2vOe+dk9wL4apSwzsWE5ASPy6J9KblYt9zRSKWUJik
dhsJPjL/xusHBmszrcCHoj4CUQqNwYA4olTfhRbpzxWIA9x8Zuw9BAMLfTbEi6/dkMnN3pl/4oim
aQ7jO3aDZ4JDLHokQ4oi+g8s9I3TrkH+0/VMMdBiEOG8WV5fFeUucYgaazQ5eGuVE5fAaS1C2JQV
mhWSbAdvf/OxDR7KQUcIkydbH9EV6q9Mc0VrjF15THwt11R1bL6ZgjXbSswvdQRpfmSAtQ+rbLM4
PqJN/yXqTB/NMe8Y8jgfsB9SYrgB4lA1F5LS/PZkPrMXg3ceEClSejBECC7gVKlbxovv9KVo2ORK
w0AVQpagwIWsmgkiZhtPdZMSKvx4ttq4iJYQrNXowLjw+yGPRrtUFYu4f5ne5z0McGU5B+/+cSl2
P93NOBFSFHH5qZXO121LB61EY3H5/JMskjXOWlhV6ROdUARRmqeR6q6Q/YVomlgYYDHCKzGVSPXy
mzaKs5evLGed8VsBaybOJPOs6qHEgLJC1ClhFHl9G3NI8W1Ie+hIP7deAXav9dgkjjtVkA/JUOh/
cOBIiixbsjxxZ3Zt8+zqYCLUHehT2t2KqC4eRJEicn1DBMfZKRIY82KnBFeSWfWtQPcX2gRi5GAK
xVeyh++KNKOCh9W61A/2NWfU6+wZLyrL6AlKZx9SjEhlPa9nloOLY7JIE6t6civxSVvMIQAXoxhM
Z5nysX4/011O7m5MkyB3ve5oV227i2vgSjKhnMT7C4S9W2w3FBlF04Yr7In6TwPD3o8MnHIY4zPQ
mQcg8XuqSeAuCgqVUInPfTINtA0sDzEcsMjxUMrpb6BGIEDr9KdK96GzJ2SoJuoItJ+pXY+Inrvy
fDy2NxDB1sNnFR47ehX74aTfj3jbUJQ5zz2aTSyU+Kfo2CiX7RKcERUayzoiw2v75LMA0nKPUSzD
n+FY1WbtLtLnDB1cTJeVBwCDfqbxDoWNyc8TPCnLmPvHqeZQN1XtUX6lxlXideSGT4cVCWnF7fwC
4VbKax31Xrk7wyA9IgdZWFJoN1HkP2OKIJNz0KYrXjxpwY3hNi++Yu5VnFl191U1MBLA8eVjPI2V
h+bv+l/lSiBA/Dzp4vgktler2trm6sQUuqw/bvXUdHjoJRXG9/EFGrSnXACD7UJEODUYWK4xlvgN
Sx5tgN306zdGSEZVLox8AuHobqZqnliyiV0wwiHGyoe3gkS4DzfrRULGwKZKFDp668UFu8lvrY5P
+yw0jbJG+Fe8tkFy889Vag+ngWyCwWeALsUTMm9C7cXr3HxmMZncqxUh3WSmObBUy1xkoKBC7o+L
uF5I5LxUIbjmTiZESbpYAlNsYIhQ9tjiwmeOQeyoUMLfM5jMpc5GTVdenAf3RnyaWNK79yl9zS4b
BloPqS+7I+KEV682Gtjn2/Rt7GwWAeudj9Ekqg8qFzy5fvIAvaYAMoV3cO/MY/snjLNc27aMVgJK
AJKWshz4yzwVI9sUmV/fHTP9Yz/Us0sZCanjx2XbimcTXwSd8tyVEncVviV7wYFGThQbHCLQ+RW5
n1pPc9QttJ5nf0yr/jN3e9us+IXR/UZ2FS1PwP4NJzv4LMNw0J2+QYNE8QVdsTqhhtzx2L5uqBFf
jqz0KfwHeJwpDifjjtGvJa8m4LXwNb9eCgnrZMFA+oNZoia3A8H652tG71Gfd7zgup/1BVrOwtcv
IFsGfr6Gbkk2qxl/RkKnlEXcQnB1JQkmE20QQilrtrirrCsSHCDHFggFKZe2p6xvdLTIkzDEL83l
TUDNiCLdB5PM7vuFPv5+dvK7cj0PIOaZQyianuUYmywDqS+ZC121T2bF8gPGhE4MI1am4XrAqIOk
LntldOqr5FQDWbIKDzjqMg+pEOPnER742vVspIgzYtrQBJW5GgCXIFXEm7l5j2QsNGVXEOOhpaJI
/mr59a+XMAFcp1I+hl+kHrHoJ3ymETIEEBXpF8ODUdFZxm+TwuOw+xD9A27TsQb/cy8jgEhYjRbi
SySaIIXrXSHeJoZijII15SQjkac2bPL1rmt84Q6Wd3M+Ug71+XewmUWyuXeJ44tQu85EbcSzF1WJ
uwfMpNxfJuy/T3Jo4R7UECK53TlJep9Pc51soTVskZeT4u+s/wppz+C2YU+ODNEIU2aGhFGBeUoJ
u/5qwveMlXZPw/2fzoSHXO315mq6rA1POJxwz4xLMJDx2dYTPIR6j/x7Gla2glUeS48KlgAyC1a6
GBpgLNfFO7mpRlU+cD+JGuiRSnZmX++tLFwE0/T1JhmxPwGPvfLrqDXQ2F5DvSsBduaLbGVxPOua
cLElBupwEqLq40uxkD4bgoHAYwp78anr2JfHas7JgZBa0o4VVDK6pibiWbenR12TGTDyK1najTwW
OKE6B20Vi6kE/7H0+8Jbn/pWO8ONF2L4syqRFlbqLDmxP4DJPjH09KDyy9TiEEjD/GxnQRFz+kMV
JiqSt/Djl/cipg3siJKleYvmEmCO/rOqMUYy7/ZTNEcN07sDbdjXsbAX2s1Zu2cOj88RffdmUwHD
ndRTx1TygkxPo8VzXE/r/50wJ53QMZS9qpSbHUQ5FlI5k1q3YBNl16YKEnLhF1EAmkOqYZE0TzEF
JMaMVlFZiZATwZUH675Li4xWxSu5cvlPa1DJzFbZRPs2FKTLYcYN0aylhkaBdP7iMu0w6dzFquEc
vnZ/H13374qTCfHP7jsCDrqUZhBpgkKddk47LzCxpuljorgGY7YNgPVnsXjvOUm9mjyajaEgwOUg
OOup/SrxL7GG7Y1/uQ2Xiwdztks44vylfpS679o66c5Kx3elmvsAXSjB4ei0+Qp+lHcMm8xCAx62
Pd+avrnfdhXjvsry3ZjieHTiCfsIdadRp71+bJlWr7AzM+OLpt5eThaRt8Dou39aAI+f6n1m4n43
wQ2FruGhjIw4N+f7p07rwfeDMdF5OEW3Csme4IOKsUDPOl0w+yvlQeKJZtEHqPkc5vR77LhK3t5M
nQ4QbiGLTrRmH3c3htHt9EUz0/spql/93XRWQQYJCyMk5dX7o7O5pFLg8antR8sbtSKTYixS5H6n
1UnBOgUABWum4EqsvdA3bAtGWhvyeYJURE778zOgPnjmQ+clVVxG1nNYeX0CHma2T3Me3N9uE0Sq
d8vJ4zS/qt2rVCMeIL7+pXZqPKxHAI4r2aPKZd70VDVZPW11Zu9qsdOedtxgp4KYoreNdGU1hxW2
rddvOvWxQwUuINwuH6Og3iDkYxaRwbHGRY08HNJkmV7bAunbKYKXzGJek+K2ShQ2WUCVZCtrh8Jv
Eaak9dXXErdytaheDAdngRNFWbSYiT/aHpe9raCTq/wtQwzX7dyfvb76ZpCozZDewwAZmVjGG//T
TTl8oWhzTRuuMjWWvYqwLtNdN46U42hSMt49A/e9iT6jsxwl/0Q4k0/E/Y4mWeVWFY+amY0kyZCz
KfPDEsbqanRqdK6o+VC7TTvetdQocaac35aydimNv7tKjZulforiX32SB76QoHe7NjxgVao4eeev
91tavxMCfn61tLc0LOgG7gGGJpKVG51t0ljPcATbXqGtacvL0RdD/Rrgp0/JlIeuRAu2uEOolyQl
0xqjNPLZK7WKvEXlRkKwIJQyB+MLpdrl4JmNFJGVYjKS2B5Y758hN7a6CG1J5Dq7/gNnylKHe2T3
qXfAoiDMhBZ5qrZPXd5QVssg5GBUR6YRCzyU3tWFjQKTKXcQoTXoUEyyOkM/aMDoZoxODX83XGF/
IQ1BhqVgJyAlUOW0rfigNx+CcvbQG4gtH2L6f5El0KWZeiAbB8newC7k/VMKdl3armblKm8o2UDX
mXZ+bXD2XIxyefblztQfuhG+/UHUI7Ny03bPuYjeDU3qlrYjTn+gH5nXtcTkMnc8zMYu5sNO1Qu/
o+UigvogLvPT9TZ+cqiSv4W65ShE2qIWw6mplrtKk7hi8+mdbyvVf+iBpbnC+UZ9NZkohZepWB3W
DgpocS3mUb+VxZhAiMk+xxU8amIzx1/aVaAkSvqUmbb+LIHZBAmcd+NzGTTjN10SewNZpfO3xDCw
hK7jn38QiAYgKOErV7L4FAZetHv7kYpjKJ3iXrVUYdABQ+zoIxKJ0wWgcxOhxwFsTNGctj/HqZYZ
staR6tDTrukzNRaWSRKumbt+IlKzTKd3MUksAdRqkkoHxyY7kaWl+ZguAm6TBCZdTpkT7sfpHUPz
bKXZkZ72rOc40e+oUWw1CfP2dZ+WjItDcK5/f0KK/1zkEm04kKC5ED0JZF3yWiQrBc03H82QTNQx
xwNptV4Puy9Bu67UarINubfR+UwqJ9Ff2mNo06NNo8/lMKqNzOFESv0X6mF18itG6DVO/kWOVpnh
DQAYQWDsZirW8Gqg469yOCMXOGhSCvvxQvo0/dZ1uGn2N19qhjoM3Jso7/jJ+4CacQPcQBXlYrL7
7+83JfHLcVydPZS7Z8O8j9ZNE+mUSTHcQfJONMkuW8dCcsuvET99JOnUZBpUx4pjPQZnfkcy3a5x
G7uweG+Zc5kQX0tMXDuYZTYJ9z9hLFnzCBCPS2C2J8KIsE1son3bw/x1EUxRey5TD0bWEqOOUFsg
xBThMCDf21KzuoscPy/J8iWnPeKR7b1yIF5qGzxmuD81+iFbcilVqRPDE9JHqiDvVVTCZEwNvJ1p
e8ynBoy1lbbUUuLuPpXY54YfWnaq3DFNfDUtbvHpvwgI/CplcOtBvs/kGJimINAcizIayVm8b3mN
4Vs+uXHWdTL0MPolp2XWPekRbhQVdk5HXBJTnjIkEP+nptae/uGiDOP3atOG/zUwEemJHaxGWROp
zLAvQrL/M8i8twQToN2LAd+p4HA8vGqqttGj5CJto2EkrAiQWo0jS+hINbHAS4N78t45Nqe+NruH
QC+r5jnvc/xOpQeQnefvUOUvPjpje8IBcJakYIiudv35QSQcozEjgOOHbRHfmFHpYvcIpg64QOjs
c8Hj0+PstDyTOEo6DA2pWxHZW9zKn6OPAG8dybwPSUUY33YiWsraXXZ2t3RFpJnssmctwUWEnMCB
XqIXwXyWJHnXM7B5kxGDQtXLxMNpxFqBYuPvlJV/Nz/SpM1j7LuKZSB5v9KsvHn7fIJC6Z0K80rC
coDnhWcAuU5YuBpQ69EuiwZZqzWIxj0hGrUXhY07HJw7PFEC2Iom2poXPe042/nSOYZUCJUQM4wz
DPZfol8iKyi1KTRpoJJKC8xSxd/tB7aaQZOWBHZavb3en0DAKVS3MzrgBaL/t7+TWrHlec3oEyXx
RSO6+5zm8Z4iswg8PJfyUI8sreQpok1Abm2oC8R/y0Y0KIvwjipRGySwXpHbpl0DF09YJRXF634X
1v+7bD88rWASGQ5h3NzoPTy+9OPWQKVQC/JSC5rOVmkK4BlQ5HQbgTzo0dMt+gzPYyK1EtULH6NJ
gDRbNR8HMuETD1Sumidd+kkDTU7OeJ4kyDsJDVnqHYx4IWBZDacAc/Bu5UPH2gBEhHOej0tDnM+y
TBheBfdZUjPvfkI9mDvS0Ik6M0Tt7KzwaCJbOmXvj61HrLAt30bizEYP5pwivtoiyuZ7ToDoCqmL
lKKzy9XOfMnSsBrn+o15HuEE7IGZMgP0yZpWN44/sRy2Or1MdSNPp64mJ5BbqQPxebB+aWTYhga6
S3tQvRer+NJLIeHUKcA8KkYUt6PsST7ErrMJZIbQTUzm4uropur8QXC1mRFsssKpSE8tykhBSQEW
oxYE5Ir/1dNwQzj2DOpXDlMXe3BauEZiRnb/+2/SWoFaTPYD1JQ7EhzVEwFuEuHNMUUOS0Y5etFu
vo5bDPT1ObDngxYFD1ac8n687Ip9HRhfuRa9+khoB8kfUYvT5rHvzgaaMuhi01787zkN98b6EPGo
FnO1F0/GmDEGWNVLhm2+oEAs08bMmHnslytBUUVVssGB3u3LKkQpm8JGDlnLCzkpb2l8ImdQtskT
WkT7odmsr7M688Gz5L1Kf+7XD+tkYtIcoUsJgbjO+BQL37OrN7F89nlI9FWqDmQxC1RRJz47zTZL
hV0maqseGRb9NOwbY3W0ZHVt9cA2yVqstlQfIrWQ322ZUSpcgMqEWalESvNAi1ymn7+01buH4Gm5
0MB2aDFQBVD/TJFBaMwJ8K4E4vhqTJwbFsx3oFrlBU/mVb38zNgHOrJ9FIapducI8wL5qtNCQNgT
WGBjgWEjePgtDMinIen1bvdHoRVoa3DMOaCjorkf92sBdOHUC5i664UzTOlRgcXspeevfWXka5FY
q/GeDylF1yRbUYEliD0aDTAMiQPpxVBocL1sraKuW6TKoMg8CVZcs1/Mr9RwVw1AhwX1Fe5Yz9Wq
a9Twm3Pz8ZvCGc1beG4yvAShIfVp0EAJcX+X3ezkSyWZEqDBAr8ypg7WuACYnz0K2cloMoQsqfge
jqfSAsbe/iKP9fdXkVhFhxDZ3woADUwz4RaB2p3rZw81vqaDOXBwW+UbZn3XOelO3LwQ22uwAVzQ
8V2GnRvGgmRXtDxoAKmqVtdhBwea7B3OyTYJpIxc36NB3juADmO6fgdwK/9HOaqgoHTyT5hvA0G+
v47kZ28IVEw1zs3XDwGzn9f0m72tyTzmN2pKNpkdSK5DkNvr81GqIRQt7WtPAmjd1MpHh/Cug9IW
FZYop1HYFuk1L1WqCoJuIJeIDx2Sb3xM2XbhUfQ9tq94VbahmfQDxuRpY3gu3Bd5Zb571C4zdGc1
ztO4IaWYc6IrrMEvRYzl9TuOjF9j+PHFWw8HJw5mQI7p35oSjDca/pVNqNFmyAtj6N1ody/Ytx6h
WVsJlLnw+MmLhso6k0BC9sgc6xLvdGTy7La88ieFZr89BxBQNvuMF8ZVwPR8KJhPJQpQy5DaGCdd
ATzvlIdUOEZpeHzZZcKS58KP406nkEQ8Skhs0EKj05fpSk1T+E1r/X8toPsOS0SspEgFDtEx4af7
CxT8QB+O3yiSVAP2h5EUH9n4aToVHoSrvMcn0m+uFd86q1IHHLfFxqYJsP8invX21+aZb0sfCd2l
6pMGkYfAGZWwOYW1baimRxTipx0QoMdrWQwzZVQyqbi/2k8CvRdZnKEHHgnt7rN0R9CqWfA3FWC/
T3+BmH3Ajipn1Gm9FCeZnonTk2ydxPIdrNZuixQjSj/3JCDjv/iyyRTBa+00s1GO95boFCpLoNrG
HgAx7xvCmqZ/CpKsR1OuNevpEfEALhC1SdMhcBlIehHzgadnDfULScdEU4EiicIMac8ZoLnUiV5b
MdX5YA342ZB04QmypQht9wuMGsb0f4J5LtC59WOpuBPFC20YeFQzOBNVwI+MbBzv4Cz+VrE80J6m
906RFrdUXc2J9o5DaTaMBvbqRBduN2Wg8rN6rD7JArCk6RC1XVOl9rRO0+X/4trzr7Rt9nY8fUJk
BLUHP1yZM3PxUu7uLJdMD8L1vqCuF/P73W1TuGu7PX/10JvBihWDmEKt9o0SCb4zwjPg2XSTZjgB
dM2LRJnik3RuMxaI+lerTAakNu7cuAXKvhQC67c2K35W4xkPcXYyLTo0NFtBAOUETDlSP3xDIfbI
2d16ieVuopuk3j4fGCOfpzBIMf2SbJ1EqgSTwW+YrMyADa9yIKm5yxwZ+vEnyJn9F8eEiJN1Ds85
jIIWYH65i9yrlZ/Dpriy4huUQpWvJPrEXyPf19+hPjofdEwq7Z2+HRLL026bc3owgq2CC+YNl8ka
E2QrQq3hUq83HR5Q+BwdnDYevrBdwL3aYqO6TQmTn2fVNMb3HSDv4Z/v3ERT6TvEucxShTK8bjJY
3TTA0JGuTvzEVlma2IS+qbIneVvyFTmuzq0NHoY/EO7vnPm2YJ3HIhtv5YXIVC05s+V5eYnBEs25
AOPj2hwG66kgFABsvrgxbEBsO8HfAJHwoXgFzBZjRk4JPzgDg3LSp7v1eyRyeVoDrwDYzhHUos1N
KXiUkjawR1HZ5OLev4f8OS/jrLviTApTFKVGKdufo/8e378Z1DjbOUruq4EB02LjF/cZ089+GwsG
PBG7i7LyFm2ddzrvQeV2tMBgRwGon00XHyIp44XjhDz0O8qywZTbhWsSFlHbxVV0N3vNjb7xvRYH
g+jrNTQmCVabqYyfNQ8A0nO9MTy63cDo6nGNbv65ZK7G3PMcnwpLTowsSCIhzIeI9xB2qHmO5B/b
OqiFhligSvFkpkvoCB7OKb7vpMl7SFuWDr5zua/HJEjQSH3kkVDN274vOFiK0m84QJeN4UzbZUSh
tZ6B2dqeRSLFvjY0kz+aucjxsboYSHcF5S/5mt7PGIYh9ssKyDMentUToqEBQp/mweIzmlupQP2n
m4FYdbNAe7r8Xgmr7p1135j132643Q+3zxOqDpDxaw/j4xP9fiL2Wg3gjlkvCrxL+YG19CX8MBAW
1T0GWmQCi+uLYqDEIyS8+qVEmWJanHusWPmv0q6yMkPzTXLU8LTh21h7nKe7Xtqz8t2x/WoXETFl
N/b7aDcvo6f4nUu/yYlyyang4fhIsIEJg23Gk7JjIoVoQywJM+G+d+PePpVenGR8LHHDTwcrsFbb
StB8YUoTjStVltl9x5c12bKVEuHhEy/KjYjFGGC/GQDHeHuV7hioS5RGC8SyrED6OFzntLXdM4+/
BrTXT637uj7/7FEL4SZnjc0tcL/XdLHvumX4RosfD+nWaf+Tqh3zg2vu5SBDlFDL6nsS97C9lLSr
FlnMOLif5eu/b0Uzapz/ZkeD48Ze00KJBlfOg786PEYh30xLZ/G6jWAkFfSxk984ItFMmk/elufk
S/HZMhduN+mthFvhKrcFtABYMB2QP/LjbXlmvl6+LCHZxOmxe7lhGIHbkh3e0sy6aTlyACP31y+M
dLYAyIk78WJcsec6C1DkyiUu77QN8axw5YuD8ynInrEYUOInQs1Oxxs5KhCrRZq3RkSoHtSlJ6r3
zCgICBhYfvw2CqTFb4BJULYbq3/648p2W64Lo2f5/+9Sx1JLlQxJOfhW+iyg17xtuGibzuri0qQB
09QwFtic9FKPvTieOo90WqPjcrpzAUNsKHw0lrHVk2dHYnp+VjE7Sj0eueTxhrsJf+1zKdYGMXFr
W5RK5YOUVG2RWY7E3rddclBgYcFnlI2TsAJ4dYCMpv+OxQT2CmZsHy0MWLiAbJfssQLxQjCi8jgY
Dy9926vWPl5Picq3R8tj2HNL/tZU8jtiVXMT9bk9tMccPBYfgc6NnHxic4iaZuz5bDQXCUzA/XSw
56S2rmMT5DqKKgjQ2830oIfEila3ZTF+wNgRB5t1pRQ/r1K0iF88kOv339MOOzwSNoij4f7awgQU
S3QR0LsnB/7BWCAnP9z54fVQ9TtVF9fQsV7H+vmLb8hmooNZ9yWZtzcUyTPOi3RHMIbtI5B8ZMZX
XEWgnT+H6fZJ3cVoFg3bBHjeW0nQFEzv4QEjkQmiRLZplUgTfEZZ84w/uIxZtt2v0Ba6xQmAaQU0
Jqh87t1Gf8XmeteEtZtd9vjChOHAN8ix1MIDjFpirQL66tjjMUfDwK2Whjvr3En9LMosmsuOHrtM
NJQsAbV+OVGZEW041+l0gGuoAYe3QyS+wS5g87evlUZylrs9Skw8J7yGRAhLBsq9ZvgxAMt29t5P
6m8G4rNIpMaC8oSapATB4ketdb18oYIYFgKMhQ6cZ9SfGGYC35iQR2aY9Qkm7qvx1GIuSt6pt2CJ
H+vtBO0c/C1UlzzE/te+6u2WAOWp5y8LT6bFl0AXTDdOfJYUP72AuaQvfV0uCJisie0fjCKB8eLV
392y+ddtpYNBMCZXMpwD/3vRpvYx4dWMywF3jHX4r4NT7mLW+hkPHZDt8LW7pRrLttT4MIAFjKRX
A+dqm00e4POIajCitD4FkB8IDWE4H9ckNPiy2pPcecEyqYX8JNjl6T5WTJilGmdnN3sMAcXkzaac
Nc20QoEF7IDxbSafzidtlHVesCktHzlUezCYqs+Nc5SfUHsF/LiZYghYkLAQeMzEVqnxUkZHDDNN
3xhlOXVsm0xQR1LwPqCHXpEYBgDbRir0o4KddAEFgGOx7XOwIgbcwk8FZzJZM0ThAC5lFppTqEtH
aGSbcH3AxnyvQDqOyLGbBv8BWQki5pMTjlHqlO5wCMqFglgalayjj78bD0pthXV0OhYi504yEI7V
CAXVGaX9sRV9zBGQ9EMdXPL7huNpIdo69IvTjgZJELhkoW66L2tYQzqEsSHVcLrPiwuPJWW+PiON
x4gioNVk6HpnPWyq9v4z6lKu9BHx8IRK8WDj6ffi7BvwXvqWaoA4lj9ZGyXiAM+KhzVtsVQnXsrl
Tc9NFF3YxNBHDJQZMFZgK47S+RWVNADcKngXeeIXzVuFCvLNaU9S0atxY8AuKopPSmqxdP1qkq/s
Av4ooK2sn0GGb5b23S89J7nB9wWNd2MbTJe5EoI6iq1DlW1/G5ZgEba5S/lydhV8S7Q5bQfWKv2G
DnvPafDpgzXDJRyKa0zu2q2l6oEMe91XKEbGP9lxGf89k9y99VJIWxilYMg7uVAKw11PIMgnHKdH
c9LqP+0a1ldnjyARZvnPXrtAaIJ2W/jJu+wLTDsvvzDQrNdusTGrbGY7OfPRnxECJz6fRMgu7HJR
nJoi/fE08oy8puX8DntQU20f4EPnSAnOYpo0K1dThJXtqYMKYQ6ALLK/7XRT7ruQdlXrOSfdb/25
HKDLXzujeLnDl//zbZKZ44KCuKFV0zuWvsl2kyq434JR7KlKwOS9zABBKp+Zivinwuj0pIX0lNcz
P79M68ENd5ZYTmm65aMYsxpB8i1B3wcB88R0MCtPtLZxrWN42JPic/Zf+aZINSvIuNzvK9+0kaDj
gAr6on4OmwQgiEaMS8WxhTcCIL68eYyuaOLXMgJl9yIVQFQYUTo5npE6pE1G32G0sYLFLZqysh5b
7jEFs4kylN0iLjivv/TlTlmfi0mXlIPwJCv5zGwA5gJFkvPBjuBw0F2Rb7MMcD6m/CfnTtqhPCmH
2fpxGuASte4UzMsWHiSIyZT2xYiO08N2avWnth1uAw46oyz4s3Ru0JZQBJyG4IGqDWHMjc2ZvXyY
t17LZr0cnG1mmjPh94uYYfEQYT8mZAD82/Wa4v9ULRRiXqOKYtX7jEhfjsAC34Po23MtC393BRGF
GFjH4ed5VcSseonCnWrGFu7aIh0hx23lGGxmldDJzYoiELv37uWJsOffEQpmM3LyqP/WOq0w/O4K
hQHMnbw6/SkiIb3cPfGLnHuh93b9pglxL+2ZLki9HXvofS0o/05/+w18hIakQB65ciTIMx99w3Nl
XQmvx9jdhXu/QV84dOQh7PfwIXx6E2n63VDeFaO6QU1yK2v0TXWNVb/A4X2R/DGhIS1T6B0qLzJI
s6uoNnKlzq3g7EpIRKfQSEmlNPf+zyceZAHAs/YvX8myg5yBzpLoMScMLkFazeURICCMGHuup9pl
R3mgNX0vezpADjmTutCAvt1OBWiPUS0SCa9WhWJJFbeIbi2kPQxuI60++/Xj4+Hl/j9YsmO6M7fz
JLwODZ62/SDLADeZnH/86GyWpEgvVg1PqDyB/9n3glMPDMV5CFGrR7f4MJZCHgcdvgMPt0cu3tOH
EG8hNcT1q5li5fg7LaYG6mWr035rW2Bk30YjXIXLvMcg+3rj+VN49AvNNORH523Bcbt8MbCNk16d
EjNAfrnRDwNjg2rlNM6MNs1hz+EMJh0aGabq3QRzwbm6BqHPtI+hX/swTRBmiuKGvA6xidpzfu1R
8xsHlO8gZB8J8Naqxw0Z+uX7UtsXCsvAad+dACJCurUFfetbN+8p6+1ndbEzS2MTY+D4pv/uYei4
dy+biZw0uZSe2+pSJh4+ZAq41Nl8fNIg3TATWrHq+HON/SLHbld/BSDjHN9P/YH6EqWDwpo3HwIB
JZhBKm5AqEC1RBH4TBV6x8NsJS6+NpiP79JWwARIGUfTGvZwDlXKm6m/1vOqQgM+0sXX8g3gZmti
Yoxq7pFK90tWBHHLLMKfGX9qpuv+5qjH7Z6Hk856uv8wzWqGc0S/sTFfQNTeSq0Tia3mG0oR4UL3
zNo2UAzv2i9PEW4CvpJkn6+KV/qvsVYz/llt1kKBQNn4tbPvR/8sMBK0DqCZkH+A3ybPZ1h9kKpC
ZnhcLbAanPMx4LhWF04RtSBmioSuhSA6ufGynOnQw0ij4JkpXgcbMb83O9kTWvTzyucDleDyjzCe
/w6WefUphLvJMC7v3Sj/wjfqI8BeXVGDRFpSkZHJCrlYmVQJDtFmIZPEPg5KmHyXdM5pJ2quyVne
bPKYDnvKP79LzvhwmzAYdAZjndGYpQ3WuwCdgrlTmjsB7fdNe0Nf+n5fY99Hfhx2spXmlOgNHygF
6g+EMmZ6cZfGIa/dfApOXmLhwgj7bNqoy2dDLELhnkzBZm+1uG3QNb9eQDooeSYJGbvwBb0qmyGs
Xcsvoxfy3eu2vwd+ummpDfz3p0A4puCznAOoCGr97QZ11c4McuwONrM0vxIXWNWywJ7Lf9KXzDKm
3TOfUxgW0oBz208e0e9eRgeQ1D6Ti1geFq5FQU4g6U/TB8nD8W6BR7dGBk5PZ5UzTP/FPtqWLj8W
xQWs3iGX881+Ze9WGL8ZY4Z7MN8obC/LvyKnC8QGSAf6KiKHG5VwOEYnUI4Kxfr3FTeOMse2+QLe
8H1nSu6aR1FfgZ3BIidR+xX/lzUn3JpsiOKYIDnT261+WBol+xUxTJaehhMx1ECeAnzi6N2aHXlL
e0OYk4Bh9bISkcAod69DXl8ZlqDpst8UUKi+88hqY/h8VrmMpf+udoGiPTjO80lvIPLoszk6jFyk
141ZZ+/zCeeP3EAjASz+SNXpeLe3C00aC5LC6JognGXRPG6cS7Yuwj+Ro8ow2yHH4VLg7GjLUoQG
lr3PRY9gwLLZuZpCqinGpu8Ox1OVoZAWCg6YbOlbE1rQ2ahJD2aNGxj2UO8SMfyTMzNzcjSTKU9c
cpCfPBlNOmwXXZ/eCStr93BGVJRJfjryVKGAoeBEhOAEnP/BtB+bj2zUTK+WLZz5pl9lNzscMQBY
OeEIK+2dDrewUBO/ETCG2CwasHfdN5EkZgGGvIRyCeLopOJRs5TuiLYsJ9SjWEn4DGPh9bn5S0tb
ctnWB1SWAMPc/kqdQW4EajvunNy2PYcFLfO4ZRz2r9RylVHK67GnTN17DQ1N1Z+cpSPF/QRs0l8A
27eUoE4Lx7/p4c2ik1vvT16QSQtJnSKXDA8owPOinmvdGm3NoRG6CdfJcMaEt6w8dTzYP0wjPKh9
i8cjAwUV92zJU8v1n4CrNf1VMCsgTYA8S73vBrtGwsk8b4pQl8+1vP5y2SsRNtyn0E3o77Nk6uPs
uJ20CTm4VZ4v/obcHgbceipmAePVisjG0mn4UUF06fT43b/Hc4c4qN5KrA0stIP9LYm2FQDIkCrH
QjdpOUs2tUiSv+xahXSTByD93SgNn/djut+YG+pNuQ6S6jsZWgy0SWLuJxcUVhENXmHC+5AzENi1
+ds97hG4DCUT0q7medLwui5/tClL60HYVL5xjPnKeXxFzeTNdT+jOSTvCZVDO9WxOOfOOFtydKxO
iQO7hh3wf5BS9LCXRvHFVHHuwIj6rQ0/HHUmVpHovvThO24DUCRoLijcbkDFchQ/9vegw3a/VAN5
kJJvYdrJgt8hq5gb0Pjho8k8JfBbXJ2GPZkoXhu9VSkOMj448iT/9fGTgeb7VsM9lLsSIqxqJmtu
I66/OEM1lSepl5r6lI2171IrG064YLqu+hbvPxXZhlrCTnz9d55fJMoDd9C45pOEw+xCICqLOsCl
3RR8mvWX7ngM1UOCW3pq4s08CFh+94cYow6LuFdyhHW0rCiWXeXk1HPKDS2olXGRofxs0OOm7l+c
LS4ARYrqirMHzM2Va+K7v/kTSvhvVZ78LKQZNjc+FA/lNv2XqUSnAsiYrUy5FEFEa5a+NiRLJcut
B7Vwc5wLhEpmA+csdS2EMDIBBT/juQPCxsk5ZqRncuCqn9MIdmTdOwSMQ/81xnexSf1+yGnQ9tmV
QZNmVA9WpEF27mHTodRdJckZQPYq+zVRvsMYLgzHNlBXHWrI4t4dFdhes13TMtDW/nNn+Rpt1mfD
GPqU80vLD0XVM4xVbuV5rKGm4wEMUgN7gu71em1rC7rQEIaalGqRVDU0QvlLZeAid7cn3h6SfTL/
zWcXvJJMBpXs44teoH+Ittt2ifyzPg44I7eRYkwZblKSXmzHcE62182spDbIdEZh0pFGbdoJMx/7
RriNQe++U9SH5EjzXZSL0pVCoTHNYY8c1I2Nlr2oQz9gTwAb7KCqoiH2D4jmbSgbrDZDGGJZavS0
w+TEbfSduJTVW13H46fNg3iqZplXdtNyVEdPNDkyYm7bPCbnqcjtM1xnrqpMsQO3BWvdJhKe3hyg
CPb2m3MaeZvKO2YRue5++mKq6GEJJogLwT6kW+8IY7NI3Yn0J82z9MdNSdH+VJYpjACcDK9aUgIf
QnDKLRrC+z+zt/p4JTNFPjzWWXMMMBsj7n9TGQ/nFyrqwyU3H8ab28+XPHAPrMX3MZH96/yfs/4F
UeaQ+i+wa8RRICKK3kE4JZJnq6FIpJ4vB0xiRd/sJwZIzpm2eAmxIKZSJWrCgDAbJu3aWu5DKe9b
2lrXtzwQmcVkjG5sfNPO+iFzSHruMriyxhiDPoLIWJiOwG2HEsW6V4t9XTMqDJmMkh/Wstrf1V7T
vhxhUv61p7Rw5c8HLQCQnabYIfJniTFcrhbe9JiIPGYn6WUlbIsfuyJq3380c6eKMRWLP4/sRHdr
0E4slyH1zMHZ2Da5gQ5oM51IYHxrY7R7LwTArE1C/keo0/IjdkXtP5GxfOtWz56Hi6MWR49GQ/he
IUs86v7FW7B1ToTRploExljYStq812RnseSjeRwMrp0Co62/6zmu2Xmwrcbsm6er8KLZpU+6wh+f
DpdJCkMUyozMybKSl3EcujiladcFF4zNLxwKj/dxMcjkq9kZt0h6YgajN/QRFRHOEYvZQXDtoFOP
yNyy0iy6giD/Q+oUbA9+JE1O6C+y0cX4OnOcY/JXorOleuKfThaMM6sHIoK0V9Fxj5ntl0JinHEI
rOBlwjRLBp2vl60DVLIJ3lFdVv5TTFn5v9y6rgsqoEsPnYM2hnwuuZ1vSrVyS3YtSyQhBrJPLW+t
R1LyZi63c+3OypRfkdGij75vqCygr744CpF/lq4O8T1Jo/ITlhiLNJzNha3+gOi6fs3U++XIMvxk
sjUK25Rm5Q/yIwJJ9yLNRl6WeHixcTj+lCvrhOEUxDawrDu6UkAe3oWBgCFT+QQ5UwBMowAF9nFE
NJod5WuyIT0IUKmq6RhZZjaeLK6Y39GP1LygLlAB9EF0hOC3Vd4DUl6GYsRBpRvM+1J6i1DAs57q
e8clpQD7xnQwV3eMGM1+txlwdLmKRdoeumeK6gz66ACP1mLryqnXzUNoRy5cz93UyEGzZXnJGj/L
frH2ilYuAoYzT4b8j8TSah9OWNxYev1qv36ckR3yDw77LsB18BkXdQKZYGDlYWAcDJ8flQcDhtck
AMNceWLW7DNzvR2gdLve3NBs9wnceg3d+zRoKJl8ozcxe9y0tsMYilWqAjR3VipS74sCw1cOi0mo
r4Tr/Rc99NtYYOT1uwWm0kvJXzBRWsaR1S1BIBeJ4zrbKcXYaV4sZda3JCZT4ZGWaXzhW8VlGuja
IIky12i04mYnUx0HrPnDkohpjASok5QDrW/tVzouPHc9v3dtbKu3IbFNEIOcYfZLG7xj43GWMTI5
BexPydLxcYvIzbtxv0EfG3uMj23zzka7qqhgXqwdnhERMWFNZL8xWq24oxjCMySZPTE9vPkt0tEz
kR+7XrE11anZOyhTMfRBWWwoWhUyOJnyYTs+EOs5tSUHKXBM7y2qUdP5a1iy/IimSWyVmBRNV++r
jXZB9KBDjVDXJTH5E+jZKeMlrU8ub5lthik6I0OegPEJzf8Y58F7Ea3TJ2e0gxQVJ/E3rAdhy5Uw
6t0u1To2T18pVk/KNUChGxLLe9znj4SSU89mwb4Wmb+xmiOS760ymrZvUMuTCi6B7o4HMaKphXbD
XaqppWqsQqBSMHXG0XAjQqRUJ/y8viUTVxY/XwCBQv/WAKu92TpbJi2ewhgL9ajmmjWeY7zu9r/X
ZjmrqxtHKrc0yiYd68IpYb9xYgB3fxQfgpnboXyBalTlZhpd8pvxNTvXKcRd/S+acj2Z29H+oDPK
x925MojlWYCyexcQUeCAXZ62rzmpvTDeSkdvRBKUIUCEQv8dBRAMnLr+voh4h4DdmjRvIjAj8MNi
yWPxGJHT/gCYYXqQOooLcRlO9SPGaW2Ytx6tBY6mIHBwhaldy0HUntArwd+ep6ZQDm3Bs1pOeYQn
KDu1Y9qHpTSx7xXtBtw/KCiy+GvYquWOBqgnRAKT4hBmNfmLzw2L8E6OErgJiKQEj8X5kqHuxTXX
uJ7vFfM2MhoN/YOzyMeG
`protect end_protected

