

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Qn7IteVsnZ/mdHCLR8tB/KgmTn8ijcYuBtDLGh2oUVKuF3qoFWhv7eC1IOCXLirwb60qousghfg7
0xqsSbRyrA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VgzxfdCZunpPyUwqbYGeC3ulpMsK7w2LNEgFOrFKGlFGTp9v30dyUA7MsiKFgCrzzKT+VrIPwMvw
QxU3GQIE0b38WJ5xx5bDenrFuj9fMfRnJLJFcG2V0iBV/hYdVoEecQkZyqCPVfkUdjfKW2nQQ9vE
YSgHM9qDx8fLqyQ6zAA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1ig4g7vOmzvtScDRtVb+tZEnSyg+feSk/Z8usEB/u9AljT40pDkFhR2JxLDYn3XXgfKo9dhNCFm0
whMJYjKNylxxgSFkNtQwR2XIg0BWg/XJdnzmvhE+MtmxAUvbHjuEhgVFiobIjRufLvFlBirtf174
Rb6IlMY8DFzGP8TNtNYlVuQtzXS4NvjPSDwmxdLLBUryIvh8XgTaS4XKcRx4c9SU8usSs2eZmKp1
PQzsFR6KYhbJsoU+KNdgC0qr7WxKSf9E11HFfNp3O241b9T36xgfVJMNzGcu/ZHXpRemcPttjJFK
GMln0o/DwR0gidlS+JLK6pgrPDgP5/6nmLlP6Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yE7rDdP/qWpLchJqOpJirpc1zOl8T978Yfk6G9kBcFGYD0r+ZC5agvccz99iMwduJEgIxwFmjnzG
7g7dI8mK6Rjj6eLbQ31Mhsmq+p5Y7KQTNM1pfCzFCw+oJzuBbgsBggo35NClB7Hfb8DM7OriNRWJ
U8K86UkzA2Prba4TIBs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BN9F+vWJYtgfrzbWbiAE08ecWOdWyzeeA+i0U6sGshkhExwtl0R/3hfy5ttqQZECat07SJZlP3jh
V4CCuSQw513kvIfiNR1n8KZK1ODiyg59gOwmz19wCVgWfDfnfDXmgYxf+0derYmc4F2n9+pXRhDQ
enznNCCvV1TM+SbAXbMWWC77ZJDkWposT7aeuix0KzNLkoMsiFOvzPJVJxWsxkGPtD/xLXraVjuo
/R9zbJjLpYz0T/O/R4G6FwuMiIZFlEBmhA8YI04Xnb8Of0h/udsHa/BIz80Zs9KgMYw1jOPT6P6u
7aYcNrAi7eu92a51ZSDtMllbDqQBzVGgrUZg9A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15376)
`protect data_block
jCREVWLUDWABSoV7Nl6ye2LDHsCC+rZaEtV8+8xcE/4yQzlhhP8MK4Xke+icWHOjsVminsNGUtwm
4nHwpv+N9wnzW6B2uxvzeHR80dxRpVfW8x2DS2/3hpY7uL/lWFu1otY6M2tEkNDXsdZh11pXuPGA
f1kSW6WVO09UM/ZDNt4/+/U/RK7wPepcb/zIbhy1Putp55LhqVFQzed5y/OGolj0ymdHrE2hRORi
eoGkxBkUuRwHAqqUk60vx83p4/qPusZxkV/6l3BGL9ZQmPvkOq9LbHaYHj13SGoVY+xI601Y/HAI
8K8RTnRvaTMfoZYBV0VEYdkqMQLotSy92sBEiXgDCkMDcDFxX5lqE9vun0pKXdQ5cdKUfTypLw9O
qfaj+YAIN/aBM7g60uClTJizWAiyXQyG6+PblO0acFoyQk8moMzTf566uEWrN0XxYKmz1pnCzFZx
HMxLASE0h4EnWzIeTia3WOpGwvKrxycRXly4Slz+UbdvvIXyjqrt5q6rCkERmpSTlwpRbRfpCNW2
O3wJObDYjJ4lIZKOBe+TKc5FkWKR7ghOkKaW4JewJOM4GsyTOa5+WvEil3R9/0sBbV9+9a9v2gqz
C0eJvCxd3zlUeBvFUbiv6lDgsB8prVDCV7CzRkrcN1IGIIPlTxbyDVzJXhzoYb7jmksw7xzRV606
Mtrh28KSLk5ZmVXNSO9DhM5f4UONYUmjxiGdeG886+cKy+9HlfKJrFCZ/3+Uz3GbBcOkxrgHTBSS
th894X76mL54+/+rgoGR5fq49UKPycfLBhrq4vOsgbkc+AU/K6RCO3eMs0QtBnvZBABCFg64GWm3
SoYh8s+MCVGG6a8b9rzjBerJuwyeJGEeT9dI2s4sqxJLP3mwyigVSsyrH4hPgdw1yZ8FXskCzspg
Z17YAiRb4eJuNpw5gtrjCNhOa08bYsHUw8aIzLj62lYvYHShZvxcUEzIi4a8QbsSN9I923SfsrW9
Kny93zQC186aDu7N32FZkKKrFkW5Q6NdlT/CAf5uoSur1e9PgEY19BVAekG66yoeFhLSs8CTgs2l
PCrSWwRoO30g99dW3Z/vZ9Zasv7eMgWBhtL1KoXvmx3oxkeJYT813p+65oq/Z10cFp5Wj9sZZKQE
aklXRaVBXFKGHBVYMPYXItwOsEUyP9g+kx4AopoumnWxTA5yngz5qAbEBekZLvxa+87Kh/XzET9x
FS3w1HKqGKAIi1ezxEiSq5EyEXXy14gJdBYgBdfsb9qUFBGgCjCjBQo7pE+1nAi0uTl8gyVnah0Q
DmrDjI9lh42hAhudwxTPJib09jRA4+TptMl7wPKg9mWOxOWZ0hW3pgs4EMMQ+mEKq8GM/JwmEH7q
9qfcdutBp5bTK2/W7mgLGkIqXklpehb0SIFzhuuOwIvcpzfBf/1LZBOU5Gl1EiHnf0MHjSGfAbvi
/InARMXYrH6bylUEan3H1m8wmXKW6qoZ49nEgUqPdEcf/zIrSHOrkj6j4S3UmoSp7bcr3mTzHatI
OQ5bmUeOmhvb2kc5X7vbMp3SvgrPG0JiwKmN3GCyuBQ2hcCQ0fMS6Qcc/8SYOfvxcPHb/olv72GF
XGAKz3zfcUUhneoQ9582pXH0kI4Ng2blnceAq6vFZSgNV563xUySelwQCHzElwYuClJmAjug0Ber
+XosUB7FlqufRdQEchm5TxDQxps80ABoJ/1Iy55JxUl6ZEiGuJSRktuldQa1rQyvw9ICl+8CQbcP
w8GpzjA+XcBpRiDJ1qrk49dh+3eMqp4IA8qgdLFkzxg5YZZMjcvdoZe6DPAXJppm3kjDEQdwjXzY
tYw03ssffhZDH6vyIxEjABGUzvaiEkbhrpEII1CRe+yqVlphmcpWrTX327c7jA1KWy2DiAxzvDQZ
qiD74NHXh3o9mCD6Gib1ZlQ65o6iJsiWksOftlMwadKRHyIh+R/wnx/x8upiKnksxfgkvN6/pWb5
6oq+Ht5fcoMJHW7U9ChVxjvzYk202MV4IM3gzIPR0F/A7h2txo34sBAUbCCIRGFI9+H165O1oE/Z
824GVbUpQPBo60//w0OR0QpCpWe/j40fYZ8Nl5NnII5tam6mxLZSB116n4nRWciJ+IcrSjVXq8aM
QI/gunMlK+zHDBC5PtLWuKr9OZiX/awrEmCl+Y2H72gmkoBIeiolNqJdGIh4rgOH8Og2wdHOv1EY
8VOuU4eivmfdvaof4seohDNc7dag6+ejsgc3kA+BHMy+DilqxJuqZXCjS8AdKR1kCtFH7Mt4Bk0U
bJGSJQHnSzM+u9kTOOMwYVFxISRqMQCV6lqwpNg73qSd8MLgiY/yj+gzVKnHN73U/4Ib3BQbORvE
mMOFSdUujk7h7NQYWlbCgA7SPSXFI4BbaI6KCRDWkcWXlEw4LPcCQj0Z8LmaTBEWycknnKoeJoXY
14rL4KDGP/ZJMWdF/M/PbAzpOHZnK6yXg299kOHfhxNLWBIj2ZxHYTQ0QTZprbME0CGFWougxMzU
CNkRx/qFCheuRbbI0jfoPc01T51qJdUF4cNQ2GCcHpySZhZko3IazjgVx78NRuKra9P3XFtXkP8v
YBimVvlvhRPpccmXRVPl0gm4pmRE9KbQ1inKxju7sy4D2E6KPfDGNWrkOT1CVvpq/ePYjTaAb61C
xNdOYdDL4TykIKKcy6eX276xYsySe7tBTSBCYcXWLgCirSx0nNIsH2M/l//RDWQEdUikwZo7u7MN
Bb4nbRHsZuFSLxZz0Sl/7W8LJE3cBFdHZE5+X8V6D4dvD3ewIgCG0lNfq6IlpLGTrNZ/qhYhASWO
i1i1WmTG4Qk1Mygh6+O5TBGgpgMjNEPgPlv6+WB+l+PEjTbn5gwHpKsTrFetuA7XMiI0fpTELlU9
KGPPd+5b2XQn5Q8eaPypaZ9p+nOTl5ANGv0u3+sDVo5GR9qZiRkvceNe0sgEXyJmomQukXXQUx1x
/mU4ui+Tf+XjEHNT/bPKp3m5JEvx1JaJI+FIz5d4ppMKOspRPM9eNq2qvez6HV9qR5jPB6nthxcf
MYJBQnC/j70NAmQjfPeIxBkdFzUlrgGPOWZ1Sa/3ftbRHJFVxSv1EJNKSk4ITIZSjToeKSJSzsPL
BDmBfw90WuPjof6YfSs5VEVUWflfcfxVtSuHGN7c0AffAAHd252Q61QLE1/NN/yiYLVQ/BURYVgt
TjEFM2e8ux9lAHCpmCpLmLhYmesheYPyoY/2Swt2M36Bv60JHBzpbELIzdYdWKQX5t3IMaLbAjbm
sOEl87+Uc6VamNiSqzqRUIpk1nThMwWM6mueVvG93bJeZszoSABflCZCTkB36oXCsCsMOw8xKpSg
dTVgCH9H0Hivg+GWEhgPZjqFQFChdW/oRrlfnQfJQckJ59g3ccdhCXTYULvfqUJ+9q92Doc7MX/r
o0L/zT7sIUyntq6aPQkSfQaatGvbnvf2V+H1j6I15+ElZM/cLye/kOSfeB/QM8qngdEW49iXAiU5
xXoBJokzT6UCq7lBKgLA9bp4O83WclpZ1a5WBoE9O/TMyOD6ORl2FBIONgCqf7rZhIeeWmUfQvja
aKQZuAhX0Yn3zwqTP2hntsxUh1MJrNHpLwq2dlBeUYB1L768H+Mr20f/9ht2+NG5DhdUwM1AUVST
3zyvtuKdyE6zQgqQlqHzmwJAMsOEhHDU1EClDJDWXcizhr3QdTbsypEya51fOyHMxtNwnwo1QQ8i
U0s05ziKJK0dEgL+mkluI+xmISo6xNs7z2KQP9jbafaSIv9JSks5X7OoFBxUf/QNJJcRB1DmM2cO
ehDrRIWjxTcSlmi/Dgco9e/aR106S7++5xtiCMHI+HApUIe6aXhayIODCn/LrTn2SysOMHK1aQ8C
h8YJX9OdH1t6J8olVi9jIwLlvRVVECdk21m6YBm0351q+uz14D5pg/USv60WKliz7lXep2lrRA6E
OjkDPJv3QwVHnlHnTXUeER5Uf863gZu7LJlq0obdZIjpxLbLT8QeineY/6unF1JwUicP0OlfWYAn
F9DX1s4bd49J0u2GcHvwDiziMabDsZ1xWf2Rj1Uw3jgtACvse+nK/uGX+qa+BH4IziKQwxWunkZt
pm1LgkR3jfyjkO+Wisg/TgroZTkg/r4INAYZbGkCL1bQ59XDqzSL4xYfcCdRgj6yvNnnxMcdIYKU
/kSn/KUnfzGeEmX/PrXfTGk63gEi7ze8DqzeFXdEG6kFJsILWoqyJnh/SAshrG6XAGUb8jghC9jL
fY+X36S8jgnqb6UFWV9Qo65fSSpekhFyp61bNJqGuofqblfIZlkj1P/UYzoD+NRCbg77V39yfHhs
S7xC2pMR8CkD/TWzsCF1DY7fpjNbmCDw6zp4G5CIWhqEmFPURrfdt7ldCNHGGvnVI/sTN8B+eK0p
OvN2mDVQdmzFUEztbkVUCRS3H2dNAiy2RMbcnrMX58UX5hVKl55xs9TPKRjj7FfMfYQ2hPmrI1DR
ftbTiqLWEt9YA3GAJStgYIAt1AlBrYgF1Xl/g7diD0Yj71ZaOnXUEdlwkRu/XzsGt7Siz/yijlcu
KRAUhUpeItR35V8Vimp9Ndk8lSlEsXo5Zp4aHQftJYNuSjcpj5KLxhmIpUzsHB7bZNhINZZFVjKa
zl1Lp65D+nH+M+PDc6lGXKSuBR8GgbotcsgREjxS7kL3M8RyLqA4Wdx5TnsDu4q6r1/+FlJBx3CD
0PSGYf+7cqbufXv1yQjydFFEuxIAD5Dozswdc/X12auE4PS7W74DlQBawhgGDhUDF15BdBRuN71v
0N+O6lU/oRgUpA5yBQUtCpubBMdR9Kl90oKUy1AaDvHHtDOw3ppVvRJ1mg+ewRKPR563Jc16pGtq
b9GFPb6KaohYD984zj4nyVeKOVe+SG9gbAcqWXD20O9+PX7NDZMFeQmH8WEKZvzmJWXlVaUBmSIQ
yM0fKkmJHT7o1VYqhdrGGSLK7vnmq554ZocFamo/Nou2h/Ob4c/LRAoKk378WDKT7VoHnLa/TVZM
nBHpXcYeoaOrCgOsEqrMQn5eOI/kXN7M4HozeN+nKK4Pig++g4bZ5hla/FiyGTh9myvEmoYoSrLu
3tqxukLF9pXt48XHjKzImsUdN6cbphdDo/qkMejqTgEX18ULKZqo9lihAZ5+WGE5HdC4dRWsZy/G
wXuN4+lUIbHROmi+f5hy8Yf9/lIEdBn4/PAi5255N/oDvWPgS3/Lsf1F66MjVSOpQpp6KzCkwPh6
MK4ohzw2NF7YyZxEssfGohC4sTMSsIXhn3aUvMy3fo0hUZu8UbFF9e5KcL3UFKyaON8lx8Axz+h/
aPiBYASCdCPbIRHWvX4xhz00Wlo9bNoDPIcIXuZM6O+0BpG/+Bqzs+bEoQtuLVDK3sIA/qmE5nST
R/bDHSEyGAevIZfrD9Qtp2B9A0XlbySTicyit3r3eLrbm8gKHgINSSOsyhbC8dJJvQOm04pQKpdY
vEUtXsZpNp6q1wdgl/xd/LV+zkAz0mQ+eM4KzQ8rYk1gJr0t7NV+aDuQDMoAVYLRkzejZaMG9Sxm
5db9kTXcuwqywxp1+cIomm1rZXLokiDBD7UBKQMPDsSXgk6sdyOs1/IIi/avE071Tus1VHlpIiSL
6SJ/3AHuip1sQC6FgZkmr6EfQSYebOefnwv3bAvOvcI8cwTRpcEJCt5qM94cP1jlGmjU31iG+p0G
sy8YWwDuSDy5ZXQULllsHRr68tGt4AcZBGnkmp2Kh/FtpCUeXwUgQ+ka4bB9s8Ukihk6NdRNJsnA
dwZmoBYo17XrYkga+GJMrQBx8K1m4VHip12Ep6sEX5cyyB5gIcQmzP1hpetWUVbLMdDPqwgV6Wsl
ZbGR87WmZgTYgskhFkuJmSdJmGAY7p3ZE+PIU0QIwnF32XNvxMzcptiR4leOo5OGR/O+HR5v1FT7
N4bJNQFEc/iVoMyAdD9TrPehqO6YyDuANpFC9zJEVan/5b3yemZJdy0AHF438+c/DOu86FZMsPSH
fa9MYUnMjEBcJr7sQSQpRKjLciWklLUlp9ANkJoxgfnl6QTr2hUsQBiJWKeitEL2RlTtdLpZBuHg
Y5cXFeUsXp7nL27Uh/VmpPU45rkCzN7Ws53ZswHf7bktIvclyjJ/XmmHkKzRJ3aklmL19kcV5Cs/
tw2y97cg+b+a40t6wvcrodgBl1xOfxVw1gG43hr2B2CbnG2y4JQmspOKpYEl1IIUA8pDA8tIMfmu
FSFrz/EHs4oKX7wrflcSXYTCma/mXDSkzZPjyyv0zeRL0sVnGE9ORNjA2M3qLfXaKoPEyE/m50nX
IZLy/RYoTLhzJ3gv026jrgCvW4Md74G81oQAEJWihIKVNcOf7uX2cliC+gPABdezJxABD2CMO443
HcJT4naLLKAMojArHMVdRdNkXNWLj4+WylwOUKreZMNKDCRikQ5NiGuFMXWUSidnEhEogZRB1Z6A
1USq4Ee/cwayhCUTm+tRve/2oHguBpluE6h7KGOqly34hJbiKzyzXVbvgMAhfpB5j1hyR59W74l2
NjWTXGyX9r84t+0/2YVXnDGOy3gwfAhp9IMtkzd23Py33fYKc1s+LvnZtqoFD9ptYaqYVBUUv/7F
GAkzXNTSlLKuCKwVKBI5uIMr+YXop/rU8b6s2iKGNy893V6aF51ntV/K1nmmDMLCpAsnWoZsxPRx
qdg7aeUDAO4Yvpz6XeFY1/wVdPX8b3QR9QtnurECTWMaazTUg7K33VUryknUR8BvLMPOadJJIYtg
LA/3MBY+8VmGYflfdc+AndKFYnU8kiyaJYcj5fTL1Bv9PCkbG7FHpFQz3jVSbFbajHb0zWANOu2s
X5wh0QNluXRN8wYg8TBDLYIUjd0F7ao4WAXToTk26y3hIQ8kxK0Ga0ySLgn7Dr4trK4DQ8PkAXJs
uxeu9NeczqBg/jyc7nA9XFJ5PmY23VLCEOm2meLJeoENxGGLX7LuvxWXdvCeXEHuyyOc1x+rh+Uj
/QW3d1hYoWwpkOqErt9gF5kMvmrd7XzxjzVBj2MDKY2H0cQkkPh91O0LzKFo8QUVWn8RUOFxkDO9
5jzLOEcJ+5ZmL4hggS8JddHGyVWQwWEtyBY42akdvRH2PTmfjD4MECUnXMu+pv1ox0MtP0rZF00K
LGxzInqT/VwLJhV3mQc2bq7/g2EeQDfAGNeMN9Cmr6C1WexV8VpOAXHrpv61LorqJ4YZzsGLP8s2
vRZRyX//T917BxhWLcUizC3bvemF6tcvsydIj9eCIGKUOqZsdwlyBeSOK8RGrhqraePQpMhQmKn0
jBpU2r3EB4kLwIPjbsP/LlAVD4lNBl6xKS4MeZ2LocfVkMM857K4m9HIIFgqp3xYx9m+/WWD4yB9
yu4S8nWkQ/+CVmkavm74lF2ZL9Wi/cqW0BepsEljenIDih5QBz5tN+S+58Sa6ON2M40QL6xZev46
mB+HyF1jYGoJqoDMjaBDCFyf/MVFZRF+EsMcuEyei3LywQkDQIIDnS4/yOyHgtHeKjuR07ZV6AAa
bnJE6NsCQk0fmZMhn8alNjhGfa+hSr13flDgfQ72JaZgwmATqA+rFOG1xnJcVxajYNC4SJYEzrE2
dQQzbFz5Pf5u4uwA2JhGBdXRvmbKQCUt8ivViM3eEoNWKNP3FtrSaBR4kt7T0pkjypuVVQ1/w+Fm
7TMoumBEau5Wmtkodx5mfZ+0RTdeZCzaZEe5SSQk7wXAggcSlRjBgkDeAAoEJEjuwkHUyrSJQdL5
AbltylR2NZCoRFNWwfi9UYodcAicaDUDsWEwChPzCaEBZikqhY5+ByxokyaUy0SnSntghLCxKSwU
ROp/E5Hbporu2AbsDJ5rNXiPAX60xVJzMnIpgloCR74Emr6pYsVV9fhbVdik6x+zNzDOBCBBfOk4
a6eXXJbk63/+bhPrLtgGcWB4Eq8bv1JIearTwh1LhGwaBC+EOjhWId4u2COgVrFJD1I+0aVgHtb5
2eYxM4yvK+quWut3pq+glpyTigFygDrUf7mjZGM5ykA5nxk0sD3VjmSRM8AIhc2VxYW9Y5wqByxs
XjlT2HUTHLhuUIVRQA9c7UnkYEQo7YHGFkAt0G4SGThygdqbtkwNnsxOZKWan8LAprBhCDJZUc+6
dG1HRReqwPSuxwdCxewSeHCBquxP8fX7suFeXBapwKJ0AlGPO+Do/c+qrikKGVUvWiOqPCQTGCOs
diwn/SxyGhyxDpTEHcdXW16vbKy31o7UfSaqWK/hbWopZN/PY7ZMJyg82Z/DPpJhjLHmZdFXDG1h
5IaeQGdfxq3heNCeL0TO4UmIVHHWeqf2fMernYTed0KuqntpcK7B6GaW0cH3zp9jEVVtqBcCAYXZ
Ib0xN9jN+9ylGYd4u3e7HRXtVOrddyDWuvsyfXcfSpQsINpzcu7NcpYZUVBL32vFlwYLQ9eDdSzG
ECK4eYgWOH6iXxH1x/sxX6zKCSbOJiOKvdCqAwkf5EXiWAOk8hRXQagHaZaOaWt6W2YxfKOF+kOp
/yC1iN7od9+3OoLsC+yk7F3h0KRpPu5pBbFPnPtb0gT/bjOJKUKDrMFBFz2rzI8NEsAhy5fjdaVp
VVORaIJqLl2C2J76KGLv+k4CPuDJo4/NlriPoQxy/Fkee2So4e4nV5QDDrOYZAK/TNSoL+OtmIfc
LdjIQJNIqXkval4HEDcAF60GuayuI6LLRP/sEkvVqiF+xeeDyQQ5zxEb+l+TLRQTZ/lvpZYUDgwB
rb5EMuPM0W/OKVLTt9Q7rN3ER6Vct31GY3JSdJ2JIxMveL7jPhPOyWRNztHfnh/inG5Eh3NFYZbM
fIxrAabROlwW6NNpEE3yKQ75QVvNdxVrxC0S306m4t0rUGQs6DkyRpTACQm+ap3eP+q7/2VEvRT9
cvNuKEAZ32dM34CUrSi6snEpz9VY+RzPH6QX2KIo4pvpV18A4uLjVPHxalgoipN2muVnx7Wa6fHD
jxGQzIMLx7ZUDdM20f6L6XITuPcR35E0OEMENaxNlYmtZddnGgqK8KbiDIc+i9vj8mbfbcfYIL0x
fYQieUU6c0Lop72ZyBs3WusaW2VhVpS2FHbqojg7yiFdZpDNuUCKyzdlladxhJW2s/5TV0yF0Kt2
FRQP2yoH9tC/rvyVq7Ie0vp9mtUiIFJh7BPVNC8S7FwlIdLLM98mutMLLtCb2j7katAotmxEX9Zg
WK6fo9KVr7LiVfddEqW8AR53NH3mMjtq5eEXg4sa4M25fxtIg7aVqimUdcY4zR07qpBfE5wCRTlU
14xv3o/FqnnkjKbIqbBx59GTUGRm5ElZTVOZW2gpgZeJrK/jn8wBecU6W5lDioHOzXwEBDvWO53C
DHmxdVK043ga/acUhErxw+CjtsEAfZ6cwlAGUFwfTIfUaCdPSv107DCJxl7Nv9ttwYfWB2pxj3Jj
m5FCeccgb8txMNkQA0bUQ8pSWRg7ZduB8t/UwLy8XFDLN3iv+TWP5d0cXlB7xLl966ukhNFRSTw7
IYLIn+FSRjoj2zzeQJapvdSkerZ1G7ADJTQAt0zObQCsZ1kusjAtnw92b2dTQgO95/gaSSnIbU+k
nbhJjcqoMyr5E3mUy8eONhYiuzlC7CVO4RB5WmP/JaYzgk/dYa7JITtvpdDTs6rSjAIIdVqIFw47
u0kISL+E+ZT3xqn3RrvvhC4qFLLuHpeY9NO3HYhHdoOcD9bqh7SGLtowu/ACOnTomewQtXDKeH4R
5cd+k1HcIDRXf3TWg8W5UPjQCeB5FuI1wPbVtAPSFgm/mX4Fnb+AfAUQ+lCIhLQnzSHGtGDP0iVl
MmPsdUMbvbldcJSSLNjrTP/Jm+snRPtEgv28ZzVOvYEl8d7HzguE4/LbuqfAqd68pi3NttelMrKI
AihQzQdNUUCbENYZzNUGkpp12Y6VwzdicsqiByDtqgl8O3pImZWJGwscVdmw6gA3lL13hXjbALWn
cv+ATpqdCz2sxxqdVf7VNLcCRrvNNTIYmOY+iBqpZjKi6NePS8eySwjIZ7mQPltegS5YZSQCq2kz
OLRFkQwHuo1bgNI0mp7tLaZfsK5G6+5dEoZO894jSuRUvzBkXhqTxb3hvgQkf+r6+dcNTNbXrmT3
5NBw887GSthyhBGCnHoeQgN8vvKjEacTwPHahLeGI7fhU4WazLIq2GKS4k77HZiSQIebjQjNcH5m
B4yLO17oaXWpDcXufmZzzhDt1iyCamOUKAk1/O3awDqtBv9fuKXJ9FAeeeFFgmlxqFPKy2b6z6l2
50n/HunYuEU5L1ALFROWTyL/JbG+/D0IMoXVWmQCf9l5DZF0EhasjbfjHQrdKAdlPkB1Lj1/rRyW
A5lfjMpYmqGqWodmkIO+Ugw4e3oKvbYjt/4JJJQoyuqHFJt+oCpfm4mVRtvgQuOW7Jh8TYS8uSn7
rrsvCnS+7dBidfi5MW1kkktAwpBWrcFV0ry8r9Xjp64UoXXBPdDRCaYWvIh/HGrlugxn4G0OIfFZ
eAPUL7vGYLbgLHnMKSAaFPI1Jb9fNEmzu+diuiEE+5HYpFjwCwQF90M6jlvIZT0ZMOLuyqXt+0dx
dhQvw9jYMnvklncY+cF3kkmVkaY47m8S0G/m8EXTO+j1PL3FJTqOuN3xIiCtTOjR0HWlh4zabCB/
QwkmhXn31LeVS+4Riwr9HoWa6gTgkGyk1Xkyum54zBqMamqXMXvrhfFdapM9WiYW+zI7bh7AhE1C
jdNTp8YyWjnL9csloJb7mgqbhPTBFyrNkvXrMQVY8bilPBEqOCPxbLLciiQ0NA5Qj3xEYfF8TXDo
xzvUM8n/BFQSXnwhiTnqqgLoEVLXZNx+0IgcnzVLoQ5obxtcnoeCgQFl0F+awGtTra5wj+F6lW8m
97Zygwmjah2BWASBYrjyjQhaqgjoostA9fzRXD6KumzsTcMyYWc6dWWqxqxICiPodOdRRttDaYKN
GOXdEzdsQWrXIdMvKJRjsIb8FP/L0JFmDCE7APeBVG2lyI3uF/JWxwSbjU61D4pWdKCsPme/5E+E
JzIjCCU6CdXd0U6J0prfw4utsDDuB8qo7HOct4q1S47NLhg3u1VzUwt13Cxx9U846PYpjNbdwHk6
UgR3CaGSQ7JfeaVoxbxJAdZ/mhQ8rPS2vK8VqYUE3z2tlzXl8g3s2PssyEvy41kmiyQdD23WgXIZ
YWdOtlYb5vRmWOVsRTztBdfRocNd1ncwyCHTOtsn73nIxaF3pfwQaNT285CGQhslVhCSPQUllrKT
xeHHJ+1RS/koFDlp5hYFWMOukWLmFfmlu6rHQpMzdpS6777w82h3Z633mai/+kUZj1FiB49aS0tz
jNFLUjn2C4/Na3aKaBGFHJfU4hlAhrhROdb3hQU8HbNqv514tWDGkRaT78V4/JMa0oOtz2eDg4LO
NePtZ1nCf+ZNuC2oF1QEGDFkbd6cI2yGc8yQ6W0wpXJ6QcigPIeRSBO0OUsXoI+JmivFsRxF1j5b
fEZ3379b27zDCYrnzbFlcPxdHaaiQeSxhKXTnLrviytWyhOZXqVMjFYEMiXz3ZbeUyzTxILV2kw7
jDKkd9njoHQ5511VtnprMTmRbTnzUSq89IdXVzNQCD5r3NoICUqy2ycrQTu0NJSrP6xvrPIklIlG
xpzWidbsiEdCKicCPMKdawkr/KSbYtLQ4w/Fgav87xRXc5hTKjwaHQq4tqPYygLZyaNXPzLFXjNi
3GkgF6IAGzGsyezbJvu6BM4Oj975kSakK3nBdgc6ELNNXk8Lhp5VXZJJORSPXkNhjQT/WzQhn4v7
aO6YP7cJ3JWb63jiRbonji1QYPKdnEgaLFJOKNYpd+Sxzq69sMY3DVH1U0LqvrCbFWJWaBwK2un4
9c9SmxjRfFPYlssSRLkvJPOg1KiwdENyJwXDUh+Rq0SURUIlzK5ej+IQsqsN2sGzATO5cjgJDra3
m+CXOU3JJE96vbzS8JRGuCPOCVKmVdWLS0W0bUeqXmUylZtypO5bWGphzq+TurnTH2JyLERLQOXk
0sBrsozVJODOHH5K6prU711IfCOiigs7VU4zf+KC2WOlI26cxYr6P8Vjm6m1yAWwyDyaF9w1313t
vDVOuExIKgKh31Eth35dAeFn/lr/EDtVHzk0160lkRReoLoUDVdWn3Btex7yJfLze+ZGbU3E0pL+
bIU9AZMOzgFntmkRVgt+bLPg+WRQQyqVcMWTfVM3DPCEFxmURlKQOJxnCmbDm6j/tvDAw7ajB3VD
UFfKmCSbMChZQU/UOCeJ1TQQEggd/UWiuH7UwzPabGd3xjRoECqLuARn3CxYnunZrfbkSN5VEVLb
vOgFPtCS7hjrblv75WLOqajWGNNMtoa6U9gpaIacVhXuv33qW+OTa1hDfx6Sk/NMCLyc6dOPtmt9
3fIaZw2qlBpHFEHTeUMlQ+NiV8YdvnLt+1hAAUNHzwdi6Nx4WFWqCB78zvbuETER/UF/M0K7sofW
//nUrr8Opvykj/2X/+60ibEkzc5VJGmLsSnu8DJP5njQCDDEiLuLNkkhxn/2c9yUmEUZEWHIUOGz
CBHkV98s8GVr2Xo7pz0qJcHzxAQEYj9eAku2OoKPQB2IRY/JD1PVL57+ktfncy8Jbe+gnT/vCqxu
KL8Hshc5uzJa6JP4qgOqtmGTzb094YizV8E3o/nuMCiaUU0lGCWbleRNbNkCJvDMCQYRoNKRFKE8
01ZmCBnJS4wNXirYLwuEWxfbu7RA15cJVftpXTi0J+8BViAJf39CwBP+eApDYx93Jvfypd3BDMo4
dZIi5W6WvsKszIaGJDDrq7d9as4/DXYY/i2n9VzWIv93TsXNJtyu2rIfyGnkAyIToPlKmm2XIYoJ
DDlJ8jZomX65LSL8Tz9299AUbJCrdr9VpbGM2o7pYau+VYK4lB2MNdv9VI3s+TOXFAC/zavGndj+
pfCWY6T0WxQssv++qv16OWOQe3iD0yU5v7cOaN3KYgp24wn4nW8bI/3h2S5SFhiX+HWtPYteOcfW
H1i+o7D3ovZSBaiSghz2WUbMnDtznn9yP8bhqwNnDLysAzXYMYcNeBFZUfeUWZEVHo3n1z+f/MIV
DM8ldV8wetCRf4zkftlYD3SjXZTwdaErDe/IrimAyNImZ6RZmex26tR6USce6GYIRXsR91wrJMqY
HkJNDfiai5efxusBsjUf/6axJV1EeeppC+AxMr+2765LNSGnfqgMUGBCUtCGfLFGKj1dqGQgKM8c
BMfSuo/CFkr1KxIvTo3zqZ6rAWU4QfzUAjgb8P4RDNnGgBZKgGyzX87CmArs7jAjU3j4+f7TraVY
Cx0Kz+IL/lIhBHD/+xMoFmynOIUZmnHTaCHwveST5v7fmj0etyp9ifcRc1hUvR9D0nZ/IGyUCs0Y
vC2kS9QZXuuOUr2swaQsnz7e0Gm1fRLRssQO58853tfHDln/DqFSqFYFzgNNE0rQ1IHdpj0PEgiw
r9YeaxWhOnJG2TcBED+kN+ASUFcQ4s3yk9M+y2iGA110SIM9Ljt+Svj0tZ99+011qnIis4WiAnuF
hTtdR7paiSluNCjoFMc2Ym6d4msl1afpR1z5mfd2AFCjegT1F5b7e94e1A+DkowWlYoLKVEmJtfy
z3vqT2g2cOv0HSJc9uu2JsqZIafgGEQn5zWRJgjBGXVP/KYA2txWQfjm7/dBfyPquDKTCOwOjriX
BpVI2iCT+RDJNkBEnxIiJwbk+yqIjytZdaJNOQxGyN3FYGO+TNAiFZBfaNjHnAuSXu9dVFQWeYjT
d01sW2k2hyyR+ZlVLXfjeuDm1IHtij2fr2lbLuwtqM20aYb45Jxpfqnrb2diu64pTiEG2lLoBKLB
xLap18Qz8sVlIcjsUaqBn3c54bWFF0xCkNuBpL9vaMP0GClvgeTjOlbirBMKPV0CouJak4Z4M4/b
iPT45LBFU4X4cKh58j7EMbrlBhfQMQtSySU4MGPnkvda8zSRtpb5vT0WITz1gDv/nyTaNZasuzzs
h7Mj7GiQdqOPNabSNMJwkIJfpeJPpjIGZBc0y6XLlKlCS9z+Fm6DFANzUNkryXefCHME1VjzTZdR
7TIGzQTHGbGVGrfv1+Jg4Sb+T6t5Z49RHSVDp3aQKBH3pm1nj6t/fqo92oGF9702KyZNOxSxobww
wJr69tsT+Acg5+RerPAlxBJf2ZahC/6aWnU/MXG+9h/jpkgUdVvP5B2IeuaHFfSu5v5WF3PBoLo2
FTLU+JiIPztQk2NBrzMq/9gzWu/X73hyOgM0+LK2GF5H0ih4B+OJXxIBZ0uCdHjUEbXdFmnpANtK
ZDF/ghtgY4m0KhECJX5j5uX4XvBVzg79XNN6E8sUl4KBAnqPv8XeW3nyQ/OpyxXLbJP5aUPV6GqS
CDLwv1o0eUct5uv9e+nXTbM7DX/ksSwwFVZTJNn+/5x8fcy3lFbACMjpHDwOmNtU60ngWfVPZXYI
YutucnB1rhr3p4W+z1Cx3g83cXrst5H0Z7pFx7Gj+RZ7i3dPxbpE717kM9yHuCoox06I0CGaLEF4
FPdSuiGSZIgLq+oZccxMnZr76yIsCfHg1uqnpe4wmMoj4TkzV68qV8aUcvKVXh43BLEEO5L3U6T1
mvwWfRCmoQV+Covh0zGw659KZ7LmBRDK5xjG3VTmffXhb9+yEWjYXAGYuYCzk8EIc3+G8DDobpap
hXvLzY/xS0yMk1mtCR2KXc6zz/tSHUVMnHapmYdTVprEcoAr8BcBY+zdZYXqai9dqNsQKcPmvtz+
JFk8nw8VrBVsd+nPdZgND2uHJqVkOaEBoKpTv9v+1NBXnyT4AY8FJoo93MTGUN9uc1vcZNoARrHq
77GXoSdzA++gmeaDiZUxjbIGaU7phZT5kW6teiUgxSky7Ju0YC+q8e+nc7Pxl9QXr3NRRCvMB5Gd
VgQ0UvT+hzFbFBrSuW9xgjGMtQpaWbvbuSfpYy4Uad2wg6atAjgr3Ee1Gi6bS+sZjNUOTZGutu2d
IcvuwFU56c0X2THLO64lqELApVgZIsaU3YG4yJ6HibGNVq876xjKVDfXP3oYX4S/HSHlCC5LCAEi
h5rPahbNGfTrNCctdPrNAj1Uji/aTlKdeTnFbZIlhDLbFFahV8tJu3+ygVwOybUurcEE9YtQpEGf
F17kbz0LcWPrJkZ9AtXr6G/DcMYS+onM2kmpavWMXpHzm0zLP/AdDkLRgy0i+BlL/+IEBg/3bAAU
9R3abGo2Y7iZs1QclWG+4WakDB4tuG92E0PQOS4b62XxmfGffBAT91TJA3cIGKMiZjI6kWAKPH+T
FJuXiSBEY2BCYoIazKgh9qGyJMV0MMg81BLBGb5tMHR0WIWFTaFsZloinXzlL+YIRKQNEc4IsgeY
JjKxbXAFRSOyBonuh3dLr5MM9mKRuJ4BpO9razq0PQSS8QT1WLAHPgKEItnNbLXDd3tUFGirNmqJ
GKEIO0tVrq0sk+UfwQOOdfdgS0sT8RYEL8K028RAWiAD8HW2mi6U5eVYzYb58fPqPmh0FUf5Cc3N
alEtDa2chSsBhixZDamECzhg1sIC7C/S+SVv3mx5hmJbpbO03svSnVpjTD5vBxZQgAqtIhF+fEUA
TqsZKw3OeGjaS2Jqh9Q0gpmugt5y048v6yZI4aDEMbqShmYNc+9aNK6HadHFhCM1k2Lr317ZAt7G
H2KrpHz2mSxaXSEVDFs/rhGIrExplQOrFa67GhClDOboMOuY+Fvz4v9pYBilrmGTan1LUdzvCQBL
6MVfVdZsaIO1/7OmU93KpeqToSuH9Jaj5xzmxpIpDDFRpwQSOgkw38UD221lkt7bbh1kbcQ7nhoL
h+ahHzeEiAHAkwLM3EktZA5AoKq0ukFKjHRv+8Hu6kdSyCkRduKbf/UljKggynZcaGhQWGNXYTFi
asdLv+FjBBZAklksh3vsZNWcBQZhS2P27C/CMrNMaykGSRm9vKVAPGDf6Q9stIQ7lv1ljcBeZZlX
lXUfZt9Ce7g9joo/4bvzJF08pbO0YucV3QvWeRtpP/OEjhVDCZ9F0qo3agWm9gNwfR01DPQAz9K1
MayDl4TbEIwPy+nr62zvwmENahx+Zrskm/wY8s59iTh4/NYWAvOgtMW7gutOEMz2STMXo7qgzKI5
vQGCzeih+gxCg1kZaXSCjEkmJOCohDzuFOfc5swKiN4H6b+hTauhRUaoc6WZjWFpg/GCztTyd9wE
qjyzUCkyBbB0u5fEDXJIMPEVlqjcOlep1Ef2J32yc4hljkbzil8y6pJEb4TfOpJn6hip0Rdv5UnA
nJbOfYOCKfwT3/SuEYzk1yIh+XAUrmYfXbKt5+3ZqSuXFmamtgRJs1LDA5JKcPmvt2h+sBPUL6PK
CkoDk/lW4mbgMLwqxFDdrfhqEXAVnnL2XEm2qcvUfbEIiD12QGce4XXK7DtQlQPGA2JxulosCG3I
JwGJO4zf4YHfx6Onj4gae/pGcS2B2FmfQEbupwvWjhQYMmV7CTnbwCR8FbCnnPiRNca0bwUnsYMC
JjdJa/CxXn+Jp6tc45Rf10xJlaVn1y06Px92EGZv2PqLBThV1ldbUQMoAxllB+3nWceqiUOl2xUg
kBkBogVQcYfWBA+7jR1nH0vu6NVzk1Ysb3Eosdhd3G3R51j0Jx6wiDGZGUUqg9vbr66gjEf8ayQ4
G017EyMebcm6OEX6I0N0YDrU1xrainY1LVVeekjN/nwx+WyK/NZeKdvy75Wg9Reo38IK8VYI5PpD
6JCA31l0V1/5KHpmwZZxwDC9S3n+AY6TMcq6yhif2vZ3YcLc7ulEEaRpWJOVa3S/ujqZZ5tHWSO2
gxM3MNgKEYqqoWYnFGBSWFEhrQwcYEw7iJrO6e0azFGr5V5m+yAR8bWsFnceB7IMw+zHjWEHTuL1
pSUWznzoOICuQ5VgP9MX6mhtBjRjYe/6Y/xCodw0QIjJZjOFFCjvRUbvZ4DRsYH9Ndo9iDBYQ/Hg
uQpi2i2IIX0vN/1eqIOdEqpojT3zYrpCTeZJV4AGDdbDR8yEqQK7sCF06jY5BBZjr3F9YVFmyXgo
QvBj4ISMsN/u9KRVEUPgE9kbVyc9ndnUMZ02Zn0mI5fhV9zyoOswKHzEDJL2D1tJckjWT7P99V0Z
6ZIkhAKjylqjF46cxlGqgdG/4SFP9HF2DT0qbp8VqbdCqiOAeyhlQBF0CO3lbTdKv031cJgjKk7d
htdy2/8qNTF2aKffzKkb/jsGMd5JRsfV46t3YksOH6AqXN1ngeGA8pqjhOB1O48rQNLm7BV/aU2T
67/43mn9NDxgYC8u48QcTd3thcg69K/nfQ9hUC33uH5lEMxknzV/e5IDql8zRtL6dcp3L7Ezxyni
2+dYjgyi/HGCbNXMXIV/fTr/QiKcAIOYrOA6OxCRrmTkxnLnHEX5J5rS66SJz6okhoY0hFuQeHpZ
LVkmZUiyAh0pXn+lkvoLty9o0r4u8AqTK+Px+cz3gJVcT4dj8YWC35RwDNNFCmFFketzcfbViE3W
nVoFxEW3wwlfa+/e8W5Y9OtA/NQSaWGmPSnS1NguyOre/lrJbRiRh8MJsgl566TvczynD634v8HW
01YJSIRNgA9t9yBC5ldH1XZ4t8ATK9ZoxJmr61u49+rj46TSY9EQLuwMEwtEQVPmHAmRVvwiV5ww
/lXdo+FlpEpjgYVGj9lOvTmJXUcMlQlkwOCp3E7Kzjl5uH6lS8LaW1V2BTvQZyGTjP5eIaN72LMv
Tms3xTyEFPLv7OSUVMFRFKM6p7sH1PA9r97T7ed0bRh3lvD444F1zo0CLU/uTn0kLXVHRKClW7Bi
YwONNeFWpEDYl8o3sXby9MTxYwd9fGxCJpaC6bg31ucz2tcEIwKW7PIj9+z+7aw0MiYbPRXXj3Eb
zlAyEOcZ7T3cD0o2acd/K/lIBWeIbEJxnmg2COBugDcEGDA2MZuP6nVT7NeGI9jn2PY3WKBjWrIc
HU6VpI0u16dReKQaRF261v5svhzOtYbbnxIJOR9L7rwmxZEDSmw0Ftv5oTj2hxusJiguSRTQktiA
b61kMP2UCVgU7WRK0UIdjV8Mrqc5tYy+MXFmkl5OUaXaLhHM/ve+jDqsSNAIjUGgqqzyHcoQx78V
PIgQo8kheampHM3M9gdomB1vZpQ5gHpzksppWgaPORYICO62JjLdo55Yi2t1l9/KpOvLwhhFNkhW
8lib3Czmify+Fkn75meMSh8umcJQX5W1DfC8fhNAXyvXLQOOkl1aUdxEk3HpZB6i/9Xxhw6dvDN0
Grir+NRroNRt8cy4ShII29+za0GJZQyf0pKMYWyqyGj8/T0JTMiIw8xHsYFjuCr6+z9Ucto/i++y
QuCgW5inFGFZQSaxi8wRD9r6LAsRliD6G6tWI8s703NB49LnxtaI+QeJY39UMd9LuLRbNSW9LHBW
Ffj0iBD4wDejRT8O1Klhq+0cw/PjAeVTxtRxCIeXhLbRq4gZWQt1imeKDIKMqOKDotWVSotprdl0
gj98YuvZae9FolvomXfH9tIa7ynS23p3lPmCBKpo7kRVpnc3IOyhYHMUFBg7J/5fJJokZ7+CUhe1
8yWhOq4NbrozROWJh0v0WnCqotcYRbkuiZ9XQj/rFfvmgV7MpWFmTf+0uh4SmnpjeHG8p5mc5xgN
37Xn0ne2L9bdk0iWJraGtrEmIrsoMaEVnOtTfxNm06QxBRj8vdW9nYWKtqAiOtQN5jT6jG6FXOW9
hhPtCZYoWMxYh4SNYwgVvtGuuEFkSjKj1/o3zLPTmH5/hxxcl38Q38T5Nj8cCA0eXJDwz0zxWAS8
FjQ/jM1SeEjNj7Wc16DlJY660vdt5gAUhTR8j8LDEEzjUKPo6KhAc34UFEFvL/BeoJe0oaoUavOX
TTj0bynvI3wWbvLKofP+xQ9ks3X7f1YIHRsuBreyvD/Zn7lZ9wKgjCnbOSekEmy8Vf11oSSC6fxY
xUyYIJ5bNypvlCNXPeywi3DmQwRP07kiN2s52dxRnbJXnYsZKYnnJRJ9yo75T2+R/95yoqzngmCR
52WSnb390FdFcvNwe2Z1SIzsd/0wkj/VqJlnpRwxG7jGXHy/c2N0ugIdSXD1Yl+mpMbQEwEFU3RX
uViycis5pKTzu7C3ogxFIievQc64W5GeOpURp9sbNw9ucx5ntgxr+C9rpZJqFl0aKnFYoMMc0+j4
040EcjFbY6WuAoozWcyd7Iym2oe7y81FQDjnGzgJyrQLFbjMIFLxfillbR3XsUIPFzkLoeeiTlm1
Xi6n4eKDGJKE4xmJYkx+x4mNx1O0hSAk61XSpQVIsJUjL0yIuKy5liXEdEQvMkKQ64aW/PkHtLoT
90ykMoj0wb6HAJIO+Qwpl7vINS+KAphL04IMTd0MsLk6xgmkSePZB64fvdzvnKKubLfU3/APSddy
0cGo2GlEpVHLHmURzecC2vpuYuDFiyIgeeAYk8cIKrbEAFutE2XZhYim5nERYK9zR3S8jXNU+baV
c6Zo7OKGs4tlvTipvTlhEp4BSne0WAgkX3y2Xo2GMnBknznL2lVOKIy6ABQI6kz1JfkwIE5HD7QD
ylNqEC10qypi4ld0kwvWPr8W0ngMSAlBwicSCyWezqD463VAMut2Z4ZP+G6LyiRM/K2foxqu7G9X
ESaB6ceXPdnG/yZjoCWTPUAVbQkRSTEbUS6vzAPJcMLwdbecSNNuojFB+34ZgD8PmqfEwnj7CGLA
YNsiMHpljapfTnVXsrTyRMaar7U4aPNf+2Hg9ghly7tjqd2jMZxFc767qKvNXov+J3JuffLAFiti
ue+yKtfClDdozMSt0jIlF96zvmX0adkBJaunX9HfhGQGnCpYyP5f72jEhSs4vWdAFUcvIu4MvdJ1
bEQA4JlVNYXmXwOn/uJZi4dJzhEG7VibPxWdPQCnYYWwWM6ooF0wXYIfCyki/WBXyzCGAlAR+0NV
0OAwM/jElRIAdPGhPHn4kWCuYJFoMwbPC2D6vfGj+ggnSygKuShTcqVN9cZ4Xb9Lu0STAhM9LNU7
Bu9AIKkqjcIcqAXWZNqdnob9J70EFeUmUvJLzwj1j05928DxBJlEopGF+hW3qu5/KCZetPnRWglV
MbVs1bztV0mDW/GQFVMB5/DQsiplkHlsdh91KA/SG0ymJ56gy5bsuzuuhIUssr3V7tiDo5elk36b
5664wdhOyA8VvyhZgECnv6BscVv20h1OBY2aWPuvR8w8xfifLGJ9l9lk8DoflOT+6uZ7ON5WN6Is
Rviziq5giy6aAFRzmuiBcUcUkwW0bWfLf8mECSYrZJeW5KljX738W96ApvNxNYS2OBqJ9QVPZvcH
S+RkSFwKEExpUNmNC3sX8ECqdYmmojmCs0nIwTM14eW2UdSAd6nYOJrEQ+0yrTJKy1o3OHi9Z5dT
PpoJstUFxSlbvuyV51aDDLuQuTYZg9p0LjhB1HiiQGDl1ivdw7XMcdbCbGO8gHj+YWq/s8op+l36
pbcuWCf2v5DvhUaRLL7c93VqxKyA5zYrTC2Wm1dluEixoxpFyOjblO4vkQ==
`protect end_protected

