

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kNSODHF2BA8phv8L5aZNyOOK56HCcQ5lgKBxF8hcTzwkWRF6WnOKZaH0cAk+oZsvi02J9SlLLySq
oKFSyBG2Dw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
df+BuhfNWqGLyuHwX48C4kdWet0FAm6osy35ZO6nvLm9LeYvgiC7d+QWQpEp/leK8jaqvimQleVB
qNUNsNTBZzVm+VZnT/+N9fzr+Kn5brl7DACKZQsJ/J0EK++GrIymGQB1+7LWFg6RjvqxHctXSERU
pIxXjKUtzcqAwrR0kd8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j4klfuw/RrSoDKuTiN/Si4GPF3r+1zWV61wAeT879HAyso4ajbQGVJETjBzL4XBayVtdsViewbVc
n3EWjppKn7DU95ziVUsafFQrG5PCVJ8TPZUJisZwRf1u8N8ojLSjd7Gi7vpDvGySyTXx9aoOQ69U
XzJmTqPAeaivz/FLFyjHWzMuc078i+06EYa3j0uxrNsDH6/IL5syM3QcJV3812LlPGSBhRN9Wynk
J5AcITSvkzy/dqcKICGyxp5ubBr16BEoG7l6F/VEXvTJm/kJnHW75YZ8OAQ3I6icKjHkLZysnDlK
KEU2K5X/pkwYnpID2ogdwsEuEQr/xxo42oEmKw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AG9C2Ti5ZMi5neBsWpJ1qwXbrUaWpaRO8Qn1fL70JVZk4SiqmPlFkL5Hz8GrFfE4eBlngUFZoung
TTZ2IeyMWjxhdHHDVda6+BqJtPiX+FBQnaCzRd4VBLDnB8KUn52eheU5F9XtqqkHq+oJV3U19TRZ
Rq+NhUtknFhYrHlVXfM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TuUXpu2xk+duDJnZONHfYiEzeCuzIA9y6Ut5Y0LAE72Cfiq+aIEHs4lmSaypPxj5+E8SKfd42Iqd
iKQPBy7GWczcAr4hdHMLEortigKfhxQvyiAB00CsQyuj949i0l26Eh+7iirhYh907kSXNLc4JeDy
uXkHZzsX9mKBsIZLMO2TtO0R4ECsHQbqo/hSpi0B8kY4ucdqtZfLpEsAJ7G3XH1L+CD4o7on7UAz
BPPpoVV+VIZR6heT9EgSZTHhg3uYl38G0Ezv8g8s1cbXnSuowx0B9mx89vkctBzRxFOLnzsFdBr8
DIKQCrHZfdOhrNHz4ZkgOrKjCDpwEkMA4ATVfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26464)
`protect data_block
xntCppVDDu1qeLm+OI9e6Be0/AGxhgx/zfyBGGn7sPSR9JGo0JOmnpklyg1yGTg7zyDCcaB0pVGQ
TmU6GppDmknBq75ropUQiu9+P1BaKNXwy/412C67NmNwNx+FyNFzRoV99W3KS3Md2RXVmGTd3A3S
M4/+GKZJBTB4vDHCyYK480KL/5ZeCGlCo1eAqJ8t3ya4AX/t1nKb5zubDaTxjqXOyQ4T05ciY4hT
JG8K7heW6yYWCEVZuxugjS47IaUhKc7rzY0129fTRvdOezVkQIH+rOlXdGDJgsFkQi2hJ4UKm4Vy
zwoNAkBf9lR5cg3xkD+xTDwemEEoX9RlH2KRTBXn6E182B6rvHyKNtvHEGZDeQbGQBYksLosFHxv
nHyhalIgSCBkVDWGm7UD76Wz2ymuw4bQhhh8hKizbJ1cb1UKZxiVc5bYJvWWuGcgt9kUwmw3N+LA
iNptWtVElUvIyo2ZqUFAmgXkwMeHQIaayUbIZzmm+iqe+QchWPT2XRYNcIsT7ZH9OyX4iFeh26Iu
ZL/JtRkzChQr0wWm+TmXYc2vC+hXDzr6d1k0x/ozf9yV+3AzWkq1HvJy9pz4cAP37AdEWgySrY/Y
0M+lPkuJS6o7ho6wjg+hAgmpm5biLCG/wOa2ckIXFnQbZ2db/X2X7YFH78l9SvsMGQNzJp3advfB
cOlctkkg6oMj883cCSRzbbC+w/Ib71vMuI8BY+GcrzCxN+v22f4LUjt1TwW8TIZnPdc8qkkUbm+C
KuM8RqHa/jzbwL1gdHnCWI6xNUox3N40qGhLu3t4G6SGmCZaYMonQgeYnGM7kAopRRl/lS6czFXN
lUdKYeGXoddhLBQQzly3bFdn7ZlQNd4qCSD0hP0JB3Ajw7aEJfTF7NXdBgdK/QzwPph7W6/dM1I3
N2JOeCVwQEWyg7vYZS0/D/r3XZ+IPisfUSL6LTRGHEYw3tJ73wOnGpn5Zt38NeBSg+URVu2JuiGD
gJpCB7zo2AAv37urA2FSeXz9ile/xJfFum7fa76bQb6M1bclkMIwGIzIxyIxVTB3czh11eBVP9Ws
U9ooJ1z3KDl+zjltho9w2iKeAEQNoKQBZLwiz7M3WJlBldjb8TD6Ew4bTbqgiet3hhsz7bzWq8ic
1sFyTsTm1+5hzjAV48MLcJiNgysOf3mtkAw5snJ/7Wqx3ypUdok4XJfEM8J+HaDzV2SRnb26al/o
d3zLz0ERTSzcXQpd7DEWh/p/7Q06mnroyQ9Nya8MTXrrKJTpM1CWkIPYGpL5stpV/r+n10+rbEJH
rJcYk243NrcPflEH2AAMQ7eDBHtcGu6fF9tTf4N6DCMnucxc1Uf033oHYKDpqramz4ggEuyKGvI/
9g/HaL5WJcA4ZVQeEjG1F72RxV4Yb7mBFi2H73G6cNkjamXeoIYZCmmG4bQFd7vYROcgBjLSHXK5
qXi8W6lKHLJMMQGPERBcXFDxlTRfVXpJ5UHC3VpkGlaouqhk6LC4KL6lhBcNs+7oabv2ymF8Cmxj
p5VJQpNTvJqJUVLLKcllZ5OxqFg1XINwyEYhZ/8p8t6e4zaiU2W2Xn67CKWjiO7WzIEWPsy2r0zd
08u+q7RBnKDsfmPw/3ER38VuyLC1gSUdN1CwR/Nn0y8U2sdX2ddQoLhrhqrnMSVO2Fg5CJhmi6jG
mjO+FRa4rlQG1jUdV1aNwBXwda+C90VZSEOsgipuRy5iPVhCcfehrVBVwQxWLcnWJEfC0jJBd/5r
zWDTTSed2yaUKfiF1rIfJi/8jIyB1OofDpDyBjAkgBs06xd9z98whJP5Ol41PBHVePALF8rktyjk
ArTY5gxNLanzrlGAXyCYGw4hL/PemYluJ40dKGJa0x0V0P/WT7dNVrMoQOtlp+DPXU9hsmNbrky4
UujTsDVHQ8zECKihL1F08CqTZx92MGAmVKLGCEfc950zHCLGu3N1+6sSIgC4ucMT9/aZlYUs/9oy
vC9n0MVsR0T9Dw8MRMQ2Vno6fY7Q5KqJpl3MZLkGmaSLrM+9aZERHiRHnHHRiZvtiC66bTMQu4BV
1LE53QZ4v+p+hb6WTKmSd6f22o3WxVpae8t/jTJcW/ue+/V7U5fB2f6P7DIzg7S3Krt7QHdhgTZz
ypdwX8PRuuBrg1UyCyCCyld76kR3A31kocnjAglUJMi923FXK68Z59Xd96kQJ3qg2ZEXX9IZljsU
QpYFhb+pE4RdHaKy0yh3MSIflrVvoGfmBs3he2ziYLOWlIml7Gc1ba9jSa6Ul+r8pG7c6V13/HfL
NSmh8y4EMRS7hvXKB4jTn9zQdXYL8RLGiNkLqEgRcxWjh7+VzWTcRZ0Zt/fMiJmUKAhi443ta4JH
uNPKnP361hhH3x5NE7fQPTvB3Mnh2SHp8fVUW4t9Y3p8wXjTA/XH/oi7lK5z9kGiFBU4nac+55TA
9qNAEgQO1qC2cd9Yli2aJGuBQFouACtqHGjp1OA07hvvkLIhDQCepEpCMEV5ojUIngX36LwsjBrw
DGM/eRvThzsSlageQxsR1SFK/+BT5OtfVA59GrzSvKs30npT1x2vb6zMQX0oWsrzB9LrAquOKeZM
CgbLFFtssR1yQ+76XP9L/Ax3aGIYED/WGCy2ORt6g5Uw12bNO0OyfMY+7Emmp0MwiXvVD5eKxiZi
HQ7roVe/jkNvFH5svDKT4Jwtq6tose4gRxRCXMLNDFD+MpK8rFYpBAq7iSCjGkFs9nUix7xLpci3
YUcQZD6mUAhYGYakaLgpUt+ZEzfX8w4O4AP88Ab/V32wHVrIzkrVkR5sNCw1536C5Zs09klTDe88
cHgqfnXk9T2ddzlnj8mNQcYfyemo1bWJzK3t8hFhTQg8GPuRt40e1NnPYA5S7A9RITaSxNjuwk/a
HhjuSlc4IRGcHnsCviEqeTFF6rVi9hCXZ0qik07mIDAGcDDivYsDfi0Rlvj4Ug4oruq85IlxCdox
zSqqsguik+yEXzjcOjRF/L52G0LQHKHXEbMDEW1IV/+DyvpkeQl3JLU1utJBf8kKwBP3+gYcO7Za
WLBg1fcw9ve7JDy4avhz9WJZGQg67UaLMqtABbiLHcDnFMOsmf8kWOzbdkFSQc24aIfcw0aX818j
tOWIFT1p7kfr6p8EXf42k7xmuUhTa/ahd+Sprx8GYhNs56OjqAqipRghyTJbAtsd3drbKEGodqfA
eZ117txWfKNn71iULzjfZSz6UR/4m+LUJl/2JaKD/r0HPWivUxUh0BHXMsJ/x4Mtn4Z2znNhtCtD
pDVAINr3GIbSiLkjzqsdib8iM50BWQfJHQyI2sijq/LXBi88EAJbpUQ3v4adViU5DMSgCG1I20nA
Vu398j+22IbmDByzexTnW12LWggO+k8mDmRpsjB+H/mOR9xJepfER3vhlfqPUSHgNwpEPr9UWGFE
4NfqVdkBZzdU1dbT5yderoKWgbzQrp33Xu+f3FY/zb4H4id+v/WD8zKVt8wjRJ4R5Sku/d9RsYma
jR8pXgWkZECpMF5lzeGpVNt4tm77AOkr1rvSRW1zHI0eiZ4/imdrv3zfS7cVYZ5AxZiETx1Jd4aU
97yeK0DEFPj/trx8y2csTSxo3Q17x+Gni7vIMbRtKU65AxqxiafdG0xLZewM26gQjHByIz/zV9on
E9Oj9ASEKN++yehG7Ei+IBX4/oszrl8Z5Jn3SnstlfpbnrG5j8sXINZTOBRbzEJtuftmWAUVfewr
7uvLD5EVpV80A/4qq8m8YuwtK8dJIYT6MZLHnAsTvbMhZdKVM2BQQNagMvWw60cGVW/MVRFBWawL
71B1bZ+UeCO8TOlgcksaaT3tk/orAZctXMM+BZ38clJe2C+2ZXzVIpTldzQzr7VvqqmYLTBFPioT
2o24V2jCoygUV4d+T59GjUJlyk/dTpG6upUFzroAmcv7CZb6AhT7eeN4cuiot8LxabMysu5u/TPB
rkZr5yddTMmpYbnY/gRIFZ6a1qqMt1HSWJcz/JvFVZwH2lQ2LHFBPWRhbL2o62sjN3sNmjxpOCoP
XOQTrUpDmTi+WNeIl1pra5qFJrk5PFsfqetQg7gtsG88GPtJaoFdsprUk8VP7h3uZqTJHYOIvmdh
NUUr3yO8td/JW3IGYIpZh43zGAh/NlU72XQgZaK2J4Z4mmB8dnqP1ls0QN7Xko/1yxvq14Dbx1VU
6FuiMKGtfn2LXXuZMevoTF0FMsOx8/+mWGm9UamL0k5+gNX4ueWQ153WL18oKSfoh6e3wHXtrUpr
qu+hUpTpMFVXxYcshQtYxJnzagJ+DZCzwSmHB5kSYeVrL1lJRVpCbajz/fquTo1NQmYMAfDQ7+u7
OUoSuuYQobVLiFT84rwGGvEcLKdG+NXRhLtfghPdugoT4RiKHgSBeGKxg4JFLIVj5mcoiiu1hn91
EJ2Ym3EythwPwomvvahnXzrmcDZSoMaiwZeU9tdPJn+l9ILFxq7BBXact8ZpjJt1SM0waCZm5WdH
iJ/22gE8/H1ZprZU9qjMYJECCitcZe5Pk+/oqBJ1ALNl6KglNdluHNzZrkuRylfLgebjhuldVANo
8kxkcJ5yG6EpLx8ODXUjPEGkILChf0u5bdfXGzu1kSD8de07bPRgBuU7QSQwU9kbyPJ7sb0BrtCt
G6zOZj2GKEY0KO9r3g9gMMfFfJvYlvgR8GvxqJ/j3eAB9GRlElv5COmM1wPO++xuiaTpJhGwQwdy
hVQn2U+/vNpKPGf8cyJ81WGsMBNog9i1ONw/u0i3+nZwa6VEpLZSPY43JLCsBhZAKH6RBMbjE4YS
B+64RArAaBnnl1N0xcbMVZxKNUGxGcioZNg7Ic4YhJVPXFmZTujaceHICCU+RHKxbRU0/Hy91Zor
zAbhUJsTWEggIjibut0wgTQ2IGA5slxMoIpWxGBFuAFAclJxhCpkyfAEdjq2Ve0NLQxN6qA2yl6o
vs5vFc+JBYbDOZk80cj2CnOk+HlfPP9fCRUqDeUke81sHl2SBGope0VGWwY51FFFv+VyYiqxnSHi
8BULqUWybjow+GD7Sie+jkMAiG+GI8lyC6cduvpujIzPLNwIigtmZIimlGmnbpWRApEAZlrV/TNS
1F9VY7EpOnor9lnhlHkZoGTXdbKzH8iZOAyIPtDSLjZRDowflvX4otnBLNvTi3wCNh6Jp3o44rbk
V6VOp4PLGsrma7mpfcNKrHt5sf0GGwoATQp5FLynBY8MitiuTflESgSM4YKnv7DN2kFQ76L0xpPB
JvdHkIHjujaNTo7Eqlg0N4ndMUztb8l8u9eYufHmcxD0vRxMslrDCWGgsORGmxLOQTVK6XJMOBs1
F8rfcjxpXidxy2FGSjjZkNgBbikdOqD/7mjx+nEJe2+PTKwyWj2pZZFo6uuFrr3RrcqfHhD4o1+e
pdfIhrn8MPRbeBfAUyp54qwZmhF4AlklqHYU7ImP+kmXGsx8RoaRDm1nGLf2vjpo0TlMgOqFHW8/
Uet8wK4lg16B3Id3SDMFC+DgEdwfmpzG6FjNsTMVlo/CJdV9YIXMRPQ9hzZ9qipdkC/ALZ5VzYiH
iTWAW00WVXsz6YXvZ0m88ioDMUairfNoHGkiVmXAoZCBcyeHMRLA0IohMbCa7zD6b4HeV4ijfxQe
rOLmpUCaQyP9LQy/82ZbaZ219PLnd0Q+NA5f0xF6tq72GyrJnAL03T+OoAIN42XclxWc5zKyWZy3
TUznWjT1DUVOiZImpIIZBqLU6eSRsk9rgUoYl+WYw5jGSNwcBcVJ/pSadWT6888ydBFYQZS5Lp6Q
x17rFBvmv2DODH4S0ICJGG8arXF8+zFdj/c35UeIBNSxqzpLoNvna3g8vIhlrteboAcuVkA+Pt20
aTHLc8NsHIO4skpI5y+CcvR+7rFtQGpAFIHZSSxsyTNVF4AdyTW5SP4s7zLf9dzOYxaq8ayxqrFL
qsD2vrDOc+IByp6XQNvp4ptSyEC2JQlcIKl0QSxnMKAcesWQwJU0qEu79Gs2+A67VRLYmhGwIry1
CJ4Vxdjl+MnBjdsE0b+s+94XQCjUbPNUHpbpyVF7XkZDhQJojsjqaQPGnqBnclJj6VuI3+mF/PGx
VGNQAvlmmkutO5j35ZrbC1G71IKca57qr7Y30XByB+sMaeLsXNPvB5qlfaO+W4a9bI5M19BOJXZi
ux2i1uK+0OFZ7GyP3BYwo0DZmqeDIMUeviioZfU8YKaGtLebRVsTIKH2pt6xrlISlxLtOYTo3pJh
vkVCHBx1lORQRIIip6ofLZruIRk2RDI+rE3Gi6fpZ+Gy9a7Ka+6c6ApEiWgNXDm2ZogaaT+wahac
ndXV7MQqeKostdVtul0bHNCuFcmeBB4X5Wjta9L5uQmglkJHLIhaIvspjLN4A6wMcnoYMbvhqkCS
+0mD1Wa3qgZ5UKX22Q+O2auzo0fd9sN6kiKrFpFvz4cp2an4ppWnlnEgSdq5VIEk2WMthgAwBwk7
qFNNaSZHFBytJO1jcMcC1zggcl74hWamJayD0LB4yFkTQ3p/XonQSTq804pUCI0dBM3vukjBmFGc
8k877CT8obmRwIOOjQ10tk+Blh27ns6thxxD3Xrwgfn+S/tGh94MF43kNoh8JinN050/IGQYsCYb
uHyQ1UTTlwoaqSaHQQzLWiyCNv91XOkXFp2HbJyA9WLULeMAw6Hjaw2YV7CGiNoMTqEbi0hbudTX
+oPX0E3kq2w5FuxIWWE6zP+/CJqq57YMV3V8CyOZHA8Ahsy0e4Y6QVCXgWwkd8ObTUQuDCpGVxgU
tKK3qPGXwamnYb/T5e9ARHqdghI4uQxiBrXbvFxkISWTy+7A7G92vwhVUX3A1a3ko0fcM/vyzh8O
oPTHjoAZHzAkfP+sI7bPT3yvwyAzlIJY+NQHw9OaZ06Etr97kZf9QjNjKgh+7uhWZ3aJ94BJlAd8
xMeu9PPt8qQmmr8GG7X3c2CnG6k0uC0z+KTxogzhZHsUADTVxIBqtrdKKlJLudNdAVcP6P+f174V
fRG4Ahqj1R5E+wQh+Et3fOsyM5UjEdOc7hIFxc8ermGshpLpwyVDH490k2WderBvaBIw2LKnRoiN
2f49Jinagn0wupwLYxpRsD1dKA60C6gxMDCNBg7BIzNOo09pZP7YQL9D3nPoT9KLiaThX84PC5qu
/YQzeVMju3q/dcnE5e+pCy8gECHKYWO8uU3LVvXKF8EPTlp4ncDK3su1QUqG2a+XCfS5LFa8eIII
CjCrWyur/55uSibzcFQhCadRTsFBowf4ZFoFmEtPgRHSccTdupy1lEvCh8iz/CbF/EaOEw8gpvad
zViuUAk3o1pIUdxzrOdlskMnN75FF7PTHZvLOFsQAdHGOetySVxjrZ3R4zjDZGuTjw75XS9D3Y8h
SliLAeBM9nA/5DVZbu5jdyJzAvkPoPywMs3y+JG8N1HJOIyYIgm7RPVu3vPgU48BiWOwNgtP0tcn
QCAQGxdvjkQCSwsCFsVdlpTYi70HetLE8kDZLRnuQy359VVr5KFytPpkPRge5uNIYG6c2Ylgj5v1
7eQFiEmyGtPTUrCkGu5ti1x8DQkXGZohI94yIE5VHTbsJb1tXwc2I3BxOGvc7eHOywVlKHh1Cbjj
b+OMXLEQT5rIZ1MttlWvQQUq3xmh2NfB8ZDMXHUSQE7hNKjcudge8Ew1KOLNljuCJHQiOSOa4A8K
8ySrj8rwC4MR33Mgr0Xt36URxLB7eXNHyPFBbunLAShlgHExAYiBe0yVTHpLvuCaOibNscSZffUS
H1V+TgQnmJp8z+NJTU+2Bed0ogVV6npZxT+Ld8CqBdD2u4U4HZ3khzMjPZCa0Cl9tfoSPxq5mno9
CN1Xq9YYcWerGi2LaZ/Eo9U+L+4NrdVKtSv7HATgf5CZKTUTI9j8GA7WcHnGHRajOc2jxoIRmn/0
/scG47GYAL9x20hgdw6w4qsOTp8GdC8AnLNp+YnLo1EKNsjivFhcxDxqY5T7Tolp78BDaQbgyOQe
2JNh5etfAA3Acz8RcQ68TyYDH6X7W0sDPC14uwNrFApOw+BBR0zuSbRGjENPmCaiC10IYpvuSjdO
Y4s/3uowGaBSnl1oBvx1r/+/hksRs0sdNH58VZADqlHKdgnT5e9D0KjAYvRMYsngZ6qEtA7c9dsO
ZDFI8s0fbdcWjokmPOTEn6O4uaCG6YdiHIK0wWBmGo//dX7X9j+OEpRF0XD3IYp/3w0al+IoSojJ
FrIqZhR+alCy3cWjzliLywZE4O5Y1BPwsuyy2ViX+7omzUU/U9OJzEw7Qg58gTT9L6RJwiEnl0ue
27FnAlFQ3qqlb+1E7VMkfGdKawlKY+XYxfUiUWDCRIBgSKrertq/oFCjgnVZ8VYi4tk9yDZLOodV
+7tyu5IjOJVFpAbd+lkSy3KWS/mL+wZ6Y2oKNkPVLN1iN7mPTNUxLzCgCi/h1OeVsB+6h+bgj7z4
5zL/mOq14n6lGHb3Ub7Rp5J3UO9jDBj5IYekxJYzi87sA0hqOiu1kVPsrDHdQbCgUmFp8HtUEd6L
lWPUsTqsg6i+HR+GCuxT+W5vScFFCbu+1AyoC/mHqyAvlplEXQF/9uDrXfyv1d5P+S75f8Qz+4q1
X25VbefxDYdsgkbuod93EnePrYCpt1D2VgATWuCRSNpg9UkeDUw1SdP3sYQWNZo99tBNHTgPLSa7
Az94queuwQhpZevzB9C3x+obiljq3x+Q3n4Drk2C68VxQ85hNZpSaD1GIxbY9/NYe5vMTGtHGACd
bFPdp7/cVI58K8liAuUcvFqFdHkZEpXXvh3ZQieFY73OYOTQ9Ayhwi01Amho36YqEJGl+60wmJVL
vpwZk5vWcBhaq9Kr48RicVqpLNyd9q0drsx5ypn5+0cvrMgIYjQYtJfuz0iBVVpZN6u1mUfwabMf
ni2liup01/fhkEHCcxK0FVjKkG34+aLqZR4J0R+HNxkwJ1LQwWP45FiU9sz8VB9VsegZQMsihqos
ifPSILC4LLKLrfzVmXmU5fgyk8eQ9PIOqyeLDJBTrcTYJonl6yr37gvY8cbf1eDbzdB2YJZ9mVAT
aXJMAQzX2hfDfR7vqUZI9KUbNKYQkslOoUPHKHxKDKp2p3IDDrE2kPUTkwNvJkejozqibK2An7Hl
ej0nFYY5r7UhN3OcL2iYdNHTRahVgTV0VJJyYFY7pRv9oXxozAIXyBr8ApWtwRajLoKaccKbvC2F
7OZ0mGXXrQhyg4bWQBvQCfJjixVg9UOG7VyB2DLsN649TDAL8H59PZJjSEGOPAWFQ2VjMrIK3sQ4
ayFA2bt5Q77Uds8LE/xc1wVgejbHUi/TcRThepMfKLhvQUSoxMMD+AjgqYkjQEDVX1nUqD3VCxUW
u3AngOOHBbjDMVU2auNxfe5UAGowQ4jvX8QUIdakTT/faVWurqMmL1Z4A2xu7E28oVjOuVKLKgba
BQCMywZlId6LYsyfbN59lKEP20cIpQ6gglM66sgQgpZh4aHCu0kr88GtCOpwxQaJb1mO652ttbiX
I6QH7MOfEVy422esDhpmEevIPaW51yq6EgFJ1hXp/Gg1sn/iodVvLByay01qopjlTUR+7HKuIAhe
ADyAyE0c5QrlIxXV4G5cRQWNqQwWwn44OBw/GPV4JhJXj7UElIPi/Qb0sKBsZlXCqJJ8ioIFWQma
qmlQDMjrQ9szx23xB3YOazTvl3S0QCU/CSoMXesLGf6uuTuIBfdAXxXYJxUR7xXSk8KX6vdaG5p4
DmDQjxVV21gS7Q3iEitUzhu1JKdpuxmXFpC7mZYxX5al4NLxCFssIsfPMFX2fsI4EEsbS7W8X4qc
+MtNBTstJCP3r3qBa5gbXBwAitArxGo33vcg90g2hcbIGcz92KCy4QdMxttuqrmhK2JXqWwYt55c
f5HSlVhOcJ0qmqAtRnDUQrDV5UTw+jsyIboA+aI9Ac6/0e/u8e8svwVwoAdCNApLlGV4+66UbKe+
fdjjGSlvtB98YlJdYFJkmmAFbe/r4daZYSeDTR0Ds3JAh9dlheW+rr15Ag6nngHWqjlcKsLEYnC8
JLVEeTuDEAirYPoVYypvcl2LAyVFQnIgRz5qFzwABO9TXqrz/kKe1vf63lMg0agxbMUMLJ2PVUfj
YoSLS2kS1B9BWLY6sZutvYovRkD7Jye3WQkuSSkXPBH5H+Lyzaz24FCpTozb2etezuMpWDvQwi9O
q4F2cHVYGFmZgYCqF8dkCRi946xGY8igSVL4aFbZfbuInsmhWnmNKVQcBd7q/MunvFAcE9y12JxY
/03t/GgfkMAm8ae3ixoKKU0sCU+K+HczX2p+9YLFoR3gb1SF9gHCQsId9+PtAtPEw5RmJvovJ+v8
ogt5zK6seHAtSdSPAc3jH0gKr8TTN9s9ro/vbFtJpH2AJ0nXFxNKKVoqauiMy2pAzt4ywfcJWlZJ
szNg2rBmQAzIm4b61jJyLbCArCzgDMNYnDtYc8S/5SMrfMOpC48GfgiU/E8RrC8jqxJr9L+QO+yt
WyiAVE4+r+vQsxYgmPllwN2qfjtjNniogJ6mnu4h3TlHl9Bs6NYfx1ro81H8nZr7aWC6nA+LP8tA
jIfvke8OLd85GSnJmAUmCdhbJsDWZo5a4JlwKSZgLB4zpikQ9BenhSCyvUUvJQEQufO14FoJe5ik
KdLCWxJCPn5HDq3Vp2DtpTB6qHvHtty6uuu+2V4SgaULTDbc7/S4rPhlu3uFZRasjRtQrY9AhXMf
OFkxfTmM/8Vps9D97c/Vc2pk3Bo3P7aht8FDXmsaGVfC+8NM1qKJeltkeosA84ugfU52mDn09uxc
rlltqOPkKaAhE4PQVfS7mrbs2XNk4Zu8tAv8o9Ycx5SICymMBxee+XcaVCkksKdNdFH44j2U3InO
rhor09Yj4dNMReSJtXC0kWBa3WQQ92HjAWKi23swGZaQwywwFMiElNZr0UmjR/Ynt0wcKPypY/KT
qdtfl6xrRor6W0+H2q0t6ltTFk9z0ORRjCq+hk4xv8TPhOQWUx7EQZXlK3Srj5xoXXMXrPQ1kLYN
RamNQi1QYfjd4+QhKc09N6FvsHuq3KidgGcYsftPzXths+ZcnQFHNr2gp1FLKwyrXTvMbGcoWPFE
y1Uh0iTRoqsh+lGSjB1qCBF+tyriXRvj0BaihdKUcKdMJIrWqEWuxzqH3iUA7xXa+eKTF/Z20BO3
Jr0LDDLEhtF8fwTYSjlMd2QHaob+Vxmg6+RBGTE21+sZuwKfWDo/DstpE8EGvRDpgpdIAqfLvsZb
nMy6hkN+MCyov0z1ozqFbs6co1N9z3uSCAn9Fg4diH81ZTLX1pUmMv0HLNbyHzsNzUDhSJbWem0u
dwCooOkbw/AtQZ06eJiTQQqBO40niSxDD4KsuD3ifU20xd5tJLcC4STOw8ZRMNPXwrnHJSw/JMt4
F58K/Das+2+HvcBGgk2Ksod3XLrHSxTX9Dzry9X6atfZgT65ChEeVlNIpjCQ5uU3/Q5hrr+oaUID
ZHEly8dhyB1Ihy3m8OsDUyI7mh0raxCPvFMOJ0IXhrbyNYiciU3Rkl+Y/7sCuG11OhohmB9fA0m0
sDwbstCvwX1B9mMuUV2dGNYEG7K4LNs7LAjupIuF2MGQIPSUfVeDY5bO89wwVq2kltCUAOZZSjSc
NrblbcAVVmtgNc3qqG/LCKSY2cqssJjKJeEvdK1P3lAPoa8RDuQilG/bzcwYoBraf+LaEHh60J1S
D7s8pkvcjoT2l78dnIXUVTTc3WmLKHZAfBeu2PkZ4KZ9m8j6+1D0GaMa2a7MBb5/fugp7HDpuBwu
de9xtqbpWUmd7xuwOxgO32rwDRIzBg4bt/aKT06MKyPoUL5HEtyNZNLhwAw8ar70qO62dWwKFt24
ZNirOJUplEnrFR5cKiRhcEdluGQIHSei8vXeYW/Pb+sP6HTwJDGVUuksv4O64cATf/GaenbKOHyV
9ArjV7XmKeWNEm/QzNp1z1faAt6T9b9hgPiX9epeEV2jTjRRbN9ksGW50XjLVQq3QOAp0Aq2doDv
JTuh3zUxp/Usddn7HOjk63enygTLj0/OmBNnwEDTFO57i5L21ZimOROTIScQfB2po0YPreYJb4uf
O7X9ttGDofwKH5tMfx0ygnQ0E4CR1/IWT9wMPWZWkdN1iUYFCgpAFzeb2pMEzAmMQvJSbyPINou3
1HaQfFJaO8Hk1ytFKX727a7W/e7fOSl9p8grvuKV6kQN4miSi9ey8TYU4ieW+4odGHP6o1QEFGMQ
fS3JSnYPl0q3qkIHlJQLqlnclaExBe4D/w/zbyZ2J/WtUv1HG8mvE58pE/F052Y9TiBQ8k0Oz4p3
djILqSGKmzClA0nDQtileXarkt6PMjeiT3Q9cROQvNsuyKLT1cJ0L/XNXkHbU3m2Fi8bT9N97gxC
xlhNL2zqOcOeZ1FFvrnFvbWUgMVsNu2irApNeqInQCcrB2sy2Ivu//5S6GJrLjSewxtpft9kgq0U
3dfAOkUd9q5MLFerrNJ4WbbiPQ+GtUrYdtR/nsidhX9G10aEJAT79YRPBJCgjBHCSz+Twf2yyeNA
e2/vZmYz13C42GfB8h6w/FAW6iH8u1hsSFPT0fgSXqucM/e0TSwq/ZBmmqXuNMbDK7q/60DhSTLx
1T0iahWOI8d+ghpb8pSiWe8fp/8pN+okuuSEbH4+nm9JpNgj93BBxGvxzAQeW5vpRlQdmCLh0iPK
np4F90xjAAFwHYf+L39b+gHLO6jKkyVtstgCJ6Ht8ns8cl4A/2QEAypHgXdIenKJzqJlOzo6eAXv
WgmYLNuZqcBfG0lE6tWdtV4s0Xx2zUM2FZu4CCzpzlvVepIgsnx8kwb30IljrfHxIVebtSRndUoH
sqsDl0tJHpUrsitDArbIgEPwsiHaY2J6KoQ5tsJZ7dnLL3eBi5dbeXjwSIq7YDsjOC3nzE5YRLzV
CpdG0SUN8HYEU1vxEzLm5xfXJBYoyEHxzqOPULQ2zseFTj4jaY+Jeno9reytmHfGutWyE0T6g1iY
rMcfxQcL6nXYVQO9s+yM0TQ85Malv8HN4ewbgKn/o+JPRlTHArvzsuZnBofoIa7AUMs+5LiTZcYj
wMw9tMlhk91o7TRpez8/QWWEZ4u4TmfO5hL/nCPKPmYibR48mPC3ZR10A+hgsWn9CdeL6uK7F7bO
idWvQpk/eiEpqVPz+BwGVeXkIaTXq7o44paPvl4/Z6jpX6MvIj9tswBor0m2SZDJhcMsXb4Ix7z9
us6+VJHkXpXHEDYeoHMLllMMRJaUiBYn6TtkjV8ENemnFL1iFZX2sAkwOEVXcU2wc9kzZmNUBlnP
x0gxmAck55G92+W+hYYrNVY9n0AsZWS+17woOl0aiNdvJk5gMUYTIlSyb85rRsHG36RikF6GtG/H
KmPgPNZR7JwkUaUzg6zvZPNQigdM2r5Qn+nAptRAil++TCZiGyelTtc7vRMTgXfWTc+1bdMRFlYQ
zGBIifbMaHksBpvLNQkqwWLZsVh8g6rR4z9CgghjZXOASspOhdk3SG+AFqoHF5EwPKR0zIgY8DD+
IAdDOiYE1JNFUnxfuUbAs/382kFE1JUL/Jch+gpjpx3wuQxTj2U8761UMkYprXaxI6icQtVYsHsh
/qOna6Hx1y9vgWlJyniBUdO0gqupsdjERlLbiZDldezXC6LOcfr4HE2w+IVIenOv7VBJYmuUHBx3
43I7A4EkaUyXHFzQFhl3iQkDjlvQaoKRd3uee0DxRaTovpk9PkWq0Bw2ki/MYzHqr+LZOyFJ5Nyj
OWiCWgSAzEI57S5pRjIHDSl7qL++hv+rOAGTl9D01Su86H7qN5Bw9ZBh13H39j127DDETAu+hdgN
QVVWjKtKIdnAv8WS32Lg1pyOO/RdDGDnhKPQFFTVAgQD8o9eUuhsGV2LuAbWYzDgqC6kZN1fBznH
+fnZuPHowvuGH0Lkgf8LZKGNk2uKy5cPh11aQFyNsD12D4DI2bGfzgevUB9DNbp8ReXDbpKYLySJ
hujB+8N3O8vno1pc/gBYAw8VXcE7RcgB/c5moWyLeEOkuJbHN73ELR8TOFbpyzovaCkTyuHZoS8k
/hKu9MdREjZHW/Fz0KHseTi6M2te+/uuB/Ap7Z35KegsAcY+R55IReAYE4hJY5zi1lpBL2K+HORf
vAr7ZoGk9y5yMXfMioGnHYK6G66/rxN9ZM6HJ/r6eUc6P7DvXyWy32C5uonlSt4SsSQjOepx69D5
mheUs8ppBusaby05be7K/SGNe8efDzgRrfNbLQXLzquLbVsaQW478zehKhy9zjj3ifoW/8gxN0G/
f0DXSkUziEHfIu0Ix6GNHakvMnmfRoxFixu49R1eJzHfTYPRItvMZtGkAHyS/bJwbQrXqMdYvIjr
dZgp9MKiTVah337hcHjSgY3gBLRdiqJ/ZLfzpmdEdxQE7UTE4amtjfHtucUHVp5ee5K4HwHVNnrm
Iq/tLG8+sFFpCyGwJ1rJTmBzugedHDRpYc1Hnc2pVGJ0sHA6dI5TzmlLCYW7NkPqwZmDEvPuRdEb
PFcqnROm7q11dA12kiHqf1gj5z3RRGiDNn7HpTwGTMx9FFD3QQR5aMJD0h1IxmvVJkb3iic+ch0E
oAK5OHA9BaBmY1GSPNmIqopKgxtr+vK0KgwkYD9QBno7UwYU4X9E/+pShW+j7zx7Inu8hXpLbKRG
ngAzvca9vuIRoDgCTsq/uSTEBHQbkxr+GJ2wyozEU8cYwgTUfZPD5EK+CPb9a1unvRI3txdsAkb5
eDqtYGlH1q6MYGjUNidBF0RO61u1UUuTDiCQSjPiuqG04XScghJ+d2Qgu75uKdByJuXrsDtHkKEu
qAY1MiOIJcl7XHrPXcmBtOmGC5A7AP8kO6IAJif/Pj7V0A1Az2hRmwLzp5Aj9UbYam0WTkbZ4+he
I9c3UFHbig7Vc6SVoQch+nMM9dN12yCrJIBnQy7GOwsoC0W5D1r/dym8NkRlDi0fccfNQd9nRiXG
8O92PYnSx2QIFMPJbK7fBm0MNpXIczBfvYR1zaA+eiKHQQcBDNd5PuMnubLRJYbdVVfHZrC58rKy
1UrQsDhiyeOrHBejSRnQ/Z1ehLrNlCDl3mXCAsx8TOfZVNHZdFL6NtkXk2D7Ie7Wb+UGxpF58/+m
5/JuL65YbibjH4BeOytvfTYpzhUq8aP4oNBbDv53YzZqoXp2nouOsbY5l7BU/fCmTdu/0kb2z4z6
QoEF3ZZ67Ij3QPYHIxwgBP4ol3Wl004k2vT0oJgY+CmftKpxaEDzNuXYhVSZepqbYErcUR20l1Z2
ezTtRzc0EhY0z5nQPydg9jp6Pn1sXKD6gD1gcCRKDuT9BwdWNK9ytHvt1bE9Y9d/soh2AE2VP+h3
gAX7B602DxWO16U3YBClOOkl5JVfpNG1t2Mc6bODukdGGS7rraEvQwYwBd/Z/rIxBssHpe3g0ypI
oh1nrzE92mmHWp+Ce9K9C6nSIs/d9wZXNG/28QsFYLJFLLfbVqwC1XUqVxEBORwkgBCwHZ3qLFIf
sLcITqMVmdnZNAtEY9FvIPWoTzwU9HlphNm/M5tvsAfAgVaxs2FC9qyKYVSu4h2rNB/4gfVn9ttn
LrZn+DoWYoNrKmpN1n0e7NtBHd9RbFLVbCVYmXbFymhaO6XJM1T9sG8FbuIqlYgTD7v+wL53vzUD
r6tjsxgbdwkGFzgPvKblGVsiqOVQeSV571lV5cp3dX6LaYtSevruQGd+CrazV5lw+OzdDRUSHlHK
XudXPKqlC8vJYCOF9aU0AP95X1sTV5OEFf0ER2LjhD42l80joql3tEx4aF6sh6rN9BUf0iSRp/3W
RKVNsQb5RZe0YKyh0tHjblEOqobT4X+K+EPFX6xFcj3GagrUpHONfh0K7nPvYhlSVdc8nfesP1Zm
uea+6JxsCJ4+is314LD6UtJZ3GuZn3cv7ygSqEECYcvIGfIrHk54nrMmuawglUVDevZTtasypNiN
qYrfsJZ/Oj9GFzEEt5WluNkUXkmL093tgoVg/NGvJD3I59npY9t82MgOJH6VMzP9ENiYUeW3/mey
ORclRyJaG9VMPGJBvmE6sqCOUO6A44MLTwgIUgDtNnqVshOhTPpVzMXS8czeyhKsvA0HnghYyoFs
x+S+XZtrI1UYcJ6JBhyAVyoPfiD7vniJAeMCzNUg0LV4jY+Ed3Q/iKKCwP8t0rMtZdYvZIlnTHDA
A+Z/TM8q2HWFE8EF50Pks09Dqr0mJsREIyQguDQ1GiqQVXSdBae7Qp6hmACyQjo2+ZdShmEXIRmQ
aWsEGtDoZjH6SDS1UbX4gMRs320Ij6FLpXQ/KPKdG1gAezNEHka0GHzGBPrwADfBf0CIoiqfu6Sp
1rD41BicRJzRsaADQnDB3EpNUZZyHAOytTXl/faq0lsVK+7yNQsCX4vJfn+5g7FlciV0k+Y5xxzM
DhzqofVo0Fp/yauRWA1AZiyipXckQcap0AmI0hdIvdVpIj+AdBF43MlydFzRFzQsnCNcYJVo+AXY
w9HDMqBvm5cUjShNmXr66EPtYUs6ge2C711rhG1NrdIPTapiTd3xlyVex6EemWsZV6T6iguvQkaB
dFfakq1SqprFNUECSEk2+kZ3qmWh/1jdtcKcGVrlj0czLF2/tCnonMbNpqrOpGLURMwcJrBG0WdW
iZAivAbtn0FBAkiObvv0Q7o0V18/caSvLRRsckcRdhgyFWrFiWS31/0mMdDJ1xlKndvd1ZLzHUws
fAiJSJeUIyTYIs0eLzCbDhj8JcH0vf5PkuAAgPLUaYKqVM4/foq3Zl2n0HWNpg9Xg6UAgqtn1twF
OkPjqZ8mipF9i+Z8O9AvgMqDgT7ztElSoDCiHbmw4+NfCdJZvJOXx82SYJTbj7JhdHOoQh0fneCL
ylQuclM4etcvZJ7THuwhIAEisOeKRKceQO6i5yHkc1v+0HCS4R6kdBz//DONNwWW8N3duYPc7C8o
e3YL1gbSMVcNsEAlK5bvOEkQkO7+/9hOGxwCNeXkE9v+XhtIZ8JWGbWszZl3CzMyoInWh6ipKFfo
LoaVFB9VMaa1KA+WW6JdlRT1l6HX+SedZq1f6GbQzwNavPul32PxBs4cSt5dmRnBjqpMu4XLi1NZ
ATSknlEpB9O7jdYMEb6QV5Xnc4tkm8eC0jJZhHGi7Tebeo0qkD6w5MpMdCI/XJWhpxNIOAus0h59
MRdF/mQ5GaKXqjdY5UzTUr30H1KzrwYi4ct2aq6rzBh8+x/euDlhcIffQOjftSLH8R8qvrKjwUqY
ytO2+j6j4jV+XREBm2KHfjPfQKEGT9zc+WZ6vLTkRwkQ5LxPPllPq9cKaj7xbfQlKPGxaX926zB1
S27QC9Ea7w5gsNeDv70mvIyC7EXqnhAqchwcxLtJCKIMfbXJeVRZKTKH+dRLKdn1d9oWUMk+pA4q
R7wpTLNWEYu482bUXQ6jIddNDgqMVGHMDPKRrmr/4XTvJnWNxubvXwON0Vh2eq2JOqeNFkwlZT47
ZD8/adfdnNiisLu5sbM6kUkC6KXcXZQuKRvmr3S5iRVqKhxRAoDcK+lQ+7/XG+nRRm1lm9wMwsFp
U1pkyvMJxPI5DQcDX8+R6kiL/WaDGJ17elEuGxXwhzlmwr2DD0OvxmPsZu2AVsauxM+IBKRbhnPE
/zsQBJkPxHGhGC1qm4bxVRDTfPpl01hDMbQDrEX7a8/18pIedWC2Xv4CsfnZHgt0XocFfpFn6lXS
sbBhrwo16ZpRsc9C8ztjHglcxMYBhK+4J3vN9ZLIyKxzX4GzpbveZHqcBPph+tVO1Rm6OI6ssTWR
lihvjd4lZOokeXbh6QYRsY+7iya4n1s5UqoIDSB+9SvrPG3HqxodFMYNd7+4pCrJHHblutBsUGqb
2bfQuCLLY5Scw1lIMxZ50GWh2emMsE+vQLtivXY37kzl6chZaARIKFhxNDSyh0JVOzvbKeoWRAXz
wZQkBL6MsKixO/6cai2EWEeGhuPeWF4Np4DS+m4ruFae3Vgfkjc+kRVhdAQ3i1+NmTzaMLRye1yT
YyG2pwpSlYqaX+zGHxVyjoIojmINluXXNjr8QRNHXWKtHBTGYsnrE/erxmyqbrWY1uJ1HwnYlUSU
sQ5fuGtEFlBl1ABcIpoHG5+6p84f1Cvzrp4A8YPdfHxveWtjhjq+RvHwuo2jeCaczbyx8poMjgj7
ARH1O4hNfG5xN5iKLCnLbU56Re4rQ0Y0mY/oXihm3A2HlXGwZ+J9xY/fezBF5HqzgiJKRI6TigEm
ycGdM4yNdBrjGZq6WpkujC7hLs8bA021cyXb7KgpLXjF6lD9jTfB8mAKV/Quf6baBkDrrrE7O+oc
x7pHjza3x4JcAwappZ8coDc9GADFr8sZDUv0NLbl+r1xCl0aSsATC5VpX7CnowNWvL0bcbRVRGp1
xZea3avRbE6tVfWYI68UiTLzkbc7+GB3MrPtgNCsAgLmyTZp7jXNo6BsGmbGTLNTroADgCEHZp8/
0EgjKTh5tH/a2VsBjWNWOwHJSkvrHjVsl+sUwMUNvUFPbcxqXQEGZyeGbMz3rVEIjNIpgf/EWkaa
Jl87DIe60BV8VgYSUabMNj5/Yzm3rCjJzoPYyjdSVY2lgjRt4DnEhRLUhDwrru/+CDNQTjcQ6VAf
bWXUurwA5gS4vDcwe9phLycAfjI7EJUADsSmwUfXVnP+J4i2t10LGMFhrELMHo2WhzMGdSq+P3xk
VLp82mmwaTE0LdiAB966ppXf4D0IeoTN2hAe04asQtoQmwcmttqCV9elf96VleN+Iz6Zz8ztgqpf
y5xfMXrm3mria18R7umaC8YSUhVg/hZiN2PeSosrLG8w1MsZwgVNIvnGWu+iihO0EJqjbeIwCwcq
Cn/muXPOFFjd639e196i9AzvV4MB/6w2HHiPNWROVGhq8/GhlzeFU4o7OkYjgSR2GsLuuh9bTgNl
5vIIDdnD581BkahDjOnPWilx9eKvrgq6VJu2yD+w4u/x5nHRT7/1xj6lOkmr2eRBgR8ftQu1bNgV
DF9pvUqweV3WORXgbNwt0lzc38CuN+oTGvRoVVULtVhS0v4ldMmJ29s+53WdPb5GRgvKdfy0hZQX
qKrtZyD5cBbRyxnEJcwj7CfoXrQWxwPqIAkoSevHDevNlvcTLWzqc/kOk/QfzQv7lretqwfpBW51
0KI0JFSOz+SNe+Z2KrW57zcEo5xSKFMzxUIGZTniA2Kl3xn4uJyn0a6q/FCwm002JBIx51H8oMOc
fEsZuSwXX8PnV6/wMYxqBgu1dgVdXV2K9JWZvYP4IdsKIWgvmx0Ecaj06UGyPOT/fgyTYDdqNmlM
hzHVdbofY6uGcG/sUrae4UF6R80yb1YR9uoZhRQlGsUjhqKOUdcvFpUusveaDSlnW+66TP1zmL57
x6QVJiisP2+K7c6z+boieE4QwoGPDbkgaAU0i9eF2bh2BEg1wcy1xX02HGBvFnnBQ2/j1D9H5Z9U
oTxKmWqXh/N2Q9vU19/TqZ3+rTrmWA7LmPbIP5iaTd75ygVpUctCIB3VinPSrYebJkmJYTh+TFzV
4snVymyU0ROL66UCcYdTMsgPCHEOO2gYkuLjSng8lFLSYeiMBEx7pcUc75Xoa5eiVhtBAESeXmuy
ll2aQv7vD57g87q4k2bmKm8RWCs81sb+DNNyMB3Hfo0wAnKuRImplQ0hU95qnY+/zM4nuQp3sUi3
RnYQkKP8ts5nrowZR1ihDGUV+E+9ztyTSJtKA+oWSGdGaubkUtiKOPP5hXp7c5u+0urDJF6q4b3P
RELYMQQEgrHH1E13AxLvdI1QQL957xjPNfJ//h8v8f69hdRforQ7xXBVcXqDEf+fbeLWBE1m/avR
C4fCbuPnepGZ3ZWTlnETOpCK/B+FYjEq2X11K4l6A9l4GMOhK18562MjvLDLO7DHUYdaHmVnfkij
DzxHmpCkxBwGIO4y8et8i1OS1MDVFDSnleOYHu8yH8EK1b+xRP7F0jRXMz/6bqS/v+tKIUhJDupq
0XVUpfdV0sJwvgDcagbuwtQPmwiK/r+DyAVqHdKW9q84MwlFSFMcfK97waHM+z9BvU7Q4cZSXl1a
p+T5HTwbJgXY3x6LC/2388SFkrpRzaKeFoVLQwT1sDVi7p2PCbLvoO2HQRawcv2D6ioT4EYbHMc1
r90vCNMM/dSWuU19j89jcBbDmwRga8rrvXKeJQrAoPVZNg95j26qESZTpTcNB6xS/v8dqA6vQZyT
yDToQwzTEvGGGCTUQFFRLRcZkNd/+g8/2CUk44/NTDoQKwrz05OPS4mX23fnc16Zema7u8G50SnK
b3veLOBE38+4tRRFLHy/ICxsUxZS924lZMIo83x4VL0ozQlHtxp4Tp5TwARNu04OJTNG4XqYuxXB
fj39DHlvKeoylkEZj2E4kgsTTM98AYsfUwQwS0WNzGzQgJfh7fsThPSCKmQ9LGtCpQhF+ZuHGrsn
aS0Vn/P+SwppFEU8MICxCaPLccqNEXtLX2aUGpwoztmW3yd0bci48DiqZywu7SCEjsxpqOegEpaf
rox/PBXgzIItWC0k8ah8Xgv55QQwlYpLEhyJGXZsf/BnED8dnGM23DADPjdkOi10Y26cLJKXftev
PRUpL7vId5kYamSEtZNLGY6de7w+oTcgSBcxAGzdm8wb49vYDwzAG1Amqv1TClRCYmOm0KZv8/RC
7/uHqt7Ghnkx9tP9/tGvhELX7Bi11Vx0AqsIELrYw8bhO8BNNJrvwfPxl9BEY16ggaZ+BVjbaMXv
PUSfe3qsQKdi7EFbGgZwkceLPix+C7adw5w/e8Dv6PndoASAxsd17tjNabQSkeFBVEWoyCLuoZbS
VruvO/TvA1Hov6QojaGRNhI8LVqSbh8cQKmbnhz9x+F7INmdmOVWzkmXiQCFj37AsGsxarq0PPW3
5tebYt/o9iCRNGWGwp/VTEvwkyrNTqDKJFMD9STjk2Kh4V++OXtoiNS+pdvCRcvDXQ6ZB0JEWm4S
ba50Hb1/Mgv7m6JP1amofUuXmYSn6z0J2c6iiHjdd3KuhTSfRK7iH7Aco5XVLHHZ+gBB1kVPT3X3
0j0Wwo+XLOy0I3w++yqe/eC3LbbiG0Pjt+xORDM0hyB3M0JZ1y6E28x47Y4ijsKf+EBe8OTzp/lt
zFgHByF6AvzbF9ZJN31OvkGeTN7Apgx8vEWlQWDrXozYLSiJ2QQoL/Ic7bgELeSiuhHCggYdWHgC
T/ptEGZ/gchrevz9rf+dLAh4GYtp+BeWr73wwE7XvoN6km+LsOv7be7wIiN4xclDkzDIugfhm1cz
XaImWy5geQIvdQDXpmsMr8v1yh0fnelpFZcR/9EZfjb9gB6yshP5otpO9HGnXJaN8WWzBLI3XSsy
g6zpqkUJAIpU7xhUbrSOBQFPCKq2vhnLAarGyTVJUGootzW4Wfg19Id5TQitHHDE31r87PUwGsSz
2rCoVg0/LXN35sWJnYsahgEVxqES4jD92LtkYYTUUOrICYS+PwwLxeO822BiPebS5zVE6Mpq6IEf
efqc8T3O8Yb1mbH9CvISEUctgeUL4gfi/+7PqkL5XA4Y3EmhsUO2LtBDtU9rryQmGo6pFfGW3e32
mR0Jy1bDJ4+IB/LtsobbkVeVhqcisGEwxGPa26s2Xj6SMRp+w95HufdVFt/bEqNpreOm4tsyxtK3
Rz5JbBtXwvuo8yi/F/IIZpB4lFPZqiXY+r9icsax4O5mXUrK66X3V+a4eoCqv2RKiIFx4JrRE49Z
Cx1h8GBE+sc/MNdIKKOqWWfNSG3Pf/OpXsyQHrm2mTn44q5LNZQBOywahoJUNMdVmucK3UI2bACb
LuwldXx0i3f+m/WkHCOnMJ4Epe3OWByBogKR3q7p91RikSipoLADF/NUZLnzzHYHoPyr/7wKuPlD
QNdEzK/Qlb0kPoNlDiXs9jx5R1ST1OeoPuVtPspEeJvPsnaCKX5pcDlmA/FRvId3Qv0DFsDpahyR
3SkyBegXQzdN40/tTorcqomnREw2jODfLVw9/UT0tNAUL8Gwbiag5c+emVcS9ii/ySwgT8SLROYO
ABt4ap7Z4dizWQyK0ZsGBSj+b3xChhpnvqVFdSwKxlu3+Ksl0dyrekytTJwdR2YCl7me3XjH9Su/
z6TuP/86926RyiJEreq4Cpxmvq07LjFtdl1OC9ZLU1HINd1rPEYMxzqUBWV+OQhFggeOqkNd0ihU
byUL95xATb2eZWgj5z+ycrWlQE5hMPIfRreqVUbOLbglNYsDR35Jg9IAlt31VSR74RFzJVoBHZks
NoYRe7EkoZMA54GKfHCvSahQxG7cKkqh6R8r+g3FC9znceT5goPQ9ZuTNqy7Vu9GECtJYmXfInQV
kMHy+ViarjiJmLMj/4JUNLReduvn6GApBqKxczrDxJsDIOuudwvwCe+ckriGsgds0yGNbFo9VOTI
J40Cq1k4/znBXGzKZrev/MEssB7thy+4/Ry+2ASgQoLpckdfXdJtrEwR3136md6vK6Ff5ZyAKPHq
03llTNk1/iKP6EyvWqOzFPBB8cBCgKJPzP21bEpDf37I4FXdY10GbG11zlA8fr/NtesdDJdlTLvO
tU4pHyQ5AHunDNVFf0vqfvrjeTHFUxR6r+qUViHEPS0kyodfxdff7eBvqJ7dab9s1vhjv1ZSNIyj
8y4yLsoplcO7/25FckYpf87wp7hkXckmROEHCPzjyM6DJx9THIR7TtqMml+0u7zTU/ARsmcuOUJI
mztQ5u8HUKw0MFfpL4Dn0dGutejImcfSqK5AOSe0By8CccenSX92EE91L29MNohKcj5KS9TIs+Uf
52A2lBy5kgU7ZbdHGkpSoJupq1/8yzTsjUz6wxzUKYOOAAZEC5WDsPKmVySlh3vsX3ZkU3zgzB3z
8p0jneQhylH3mcWns/YM3u90WLKPnbhJS6WlfUKQEGkuzcSAKcwlyW+9AYekTbXhgrO4Vyz9Xfey
OhpBRdSUsDc117BMZM/fPd3BiTMWI0oRKzcrNuxsy2iHSgkfjg9fA41sNvHeqWMDqAnkia3uC2gx
pZLNhxPHkWTbF3Ph2FugEVUmVwM+UFiGGuedeQfPW8L8i1l5bB22AYf18gPe5FCD0q2xwFsVx6ch
VNFfe0Ie7HDIESB+cxVsD52sISP976YY9Ew/OLXBx88YyZYbCahHUbcsmLw2vZoTV+gZWzRPu8Tq
SkvxqdBidn5f1KmRzWZkIcZO6yAKUc06bIAKEE2NZ1PQe/x5M4tsIklNFCZI0KFjB4nOGVSZIAGR
EbHcbNCoOExJkHMIkEjFL+PDulTK9r2JRw7ouPDawdgiWoD/HIM9uWxJjTpaZCvkedNhrlZQmDnK
6jUD093Fr9Flpt4rkfHe77GI8MX0zt/GzPm9wJ5E+BLrWHZH7b0+GTgLHitLrInnU1bw/nay3bnO
B46nb3rXMmlDL5V/iJuFXAO6lD57l2Sfj5l2vHH4vt5vlDfaf4HWOIcLvM6NeESrPqqN1RrOQFhN
W/6lkyNNXNNVsf2lrIYOIcvjGtib6g8q8RaZiG63tw5agb7BUM491QAuK9rqZM4txenDZ6kvV+nr
AhA8JJxanc5rVCO/cekgaE2mWXYWjECCEwtox75jDd+Hx+DFRLsUkwpdmIrQQJ0RSqF4BtW6qltE
cv8jrI1esa4YUqF9p/LgAWF7QZ9CzxO5ssXc5fb2znhef1Z/xtMlDvWtH9jLIPzy1S1B35WrQoWn
YpVqdMZpqzFphCvqfdp4Cm9ZRzcF8IoVz+L9D8D/2foiphnkzkgzpR++KRvSc6UoHFi0Izg4T58/
U6KSlh7XgWI7ddkRq1AXBd/4izBBz3rI9klwHUDVsSGMuYPclvdvHTzh8znOoV+7Q2Y5COndd2iU
fWPYHBCcjdFC3eJKG05+ZS84inP0tskiKGnRkCDRk3+89QkomHG6+ippC60uRHWjQXrlDwQvaN06
J3kv5dg1Kyo/Z9p6WSCpj5ojgNGa6SlNE08ExjXV4d0zQE8ngvtZKFSalNChTpaa8v6akyHods31
5zp2HAvgjR3ewBQPZp4/lY1Xh9p8jOzJf/fzQuQkvHpCb+EUY10YR2Ih7HTdotiBLO4vDHKZCRZc
rJiCcXqgVg5pqzUZg7R3S6SzI8mCqoIHv2nKMra5JHYjin4TIICgVoopMOTukT18C3Y94fAdHuwd
6uafl0dEWuHSsbDek0BN/5rrIOhuynjyNrkIuPVPYID0e23Ow3gR6g3dcfthVa3J8mLezvlCg35L
5i5LeZF4VYZyRkCwLT53hPSyvxhy8BJLd+oyd+neD2wCuUVEvFcABF1Rpnu+XqqXGAbqLNdTP21B
qJ2zWlBv/ZqgFwuGSx6paRUp7jLf9Ivd9grqtHAawHytNUgOuGCCM9O1+lBf6RRYRHSGU6sNcxO6
ITHMw/YlKwVn3cdgNPkri/mDgBG/GnVo3b9/KWQ4zCef9QHCVqILu9l46yA0f4Rw0PsMq0aYx+I+
XyB6CABx8K7xbP8dtLblM2dUwGylmvK//tNNqIWIvLrzbpesRT7qBI5g/LJlzq/mfQkLLeP45zpR
Nr4fXbUEpQwZXd9sBWirPTrouHbpda7BFyGP1MrVAJ7mzfOaZfoHeZnQ9givZvHsym2yh1qc/VX/
uVJbFCFuAEOPEHi3C/kr+a3w6h2xkmC3oPCXFQnPSaNimYIHHzbnUxBvxvEzsSR7L+aNMl/9hIH+
GR/UQE6LZIge8W5np5yeUJXB+peRslt389GecxG57f76J4yd5uSFNOGqjgzG4jojLUXitfBcA7qK
IyclNbOlG6xYHbQ9/rnnzTVf0hwt5759SyYHnlmtj2sJSzIQxJhOO9DyUempUY+Ly1VKdwF7akAs
XkRLQ42t0wa3fr69rWPv4jfZuVkVJBZ57qUTEOFE9pYrBNXAs3pG5BMiCaQgwMlRksNpAQf/PNhg
pRHlXvfDzpa41lbFkqmpQs7pqrzSt2vLgpArb6uVowghi1LSArx3RXI4YI4wjB6cDSL9Kyl4/OT1
rmr/QkG5DL+qKUm3WG0C4Jv2ussZ0TG8oQBde6/slJcFDkGkToGyj3lEOcEObadGKB0iaddJGh7u
vwXxPpu3ZtD4CW/5dDvFop3J7cABDgqSkY4eG9gQJukoacwCnBmyNxHa0U2cccX+ZkACvqlmEz8n
nBythKaNSw0e1x9hDgVAbMftqsc6uvgN6kaYLqWwNFz04OXsTOSL1stHQYodU22OHBacqdDA6Ped
/75t6eFs8LX4tS1fmuV7cxip2ziCQStL9UP6Bt9BN+5oZWmGSg2bI7N/aw2QLTQBkKh5OP6ToAR7
0faE5hwOA73OsNHm8SzJwpwSCgpPXaQ5TYVY7iiF4caJXXwvYHiAzbTXAyoGC57/KKdL9r9jEW3w
tEDK3gnjNP8iwFrldkujwMOaleFo1WLC+myiY+2o7T/ptS6/lYeSApVoz9RhtWCqrISVmVYgC7YQ
ffyxrLuYUyPA4EFwSyBP9zlhgzFwCvwdwaZoSJbsaFLAxCBdVO6jGxRaosaJCN0KFL9/JEB5zTGC
pEXxxqQG3xA8c7meJYa2JsPpemrYHJqZPkkJCHdtHDJVMbv3QExKYYWwgikYVf5kaPij+1FZND/y
qlqBYAAvJXQ17fh3wo0kPhBr3BIDl+AYVoEZROBaTyRMaRx6TnrfJZ8bS+8bxHxzA0ZIC5nPK2e2
HoYu0m/dxFE/uMEQgGNDVQrDX/h09WgE/QjhMyNBTRLPxQiQGiTyWgJPDdcaELMhrxXeth4evJuU
qErysTBV0D8ANss8yusDk+PmmZdKDz1+IO0soamYt8/eriREJwJI06tsxVxNhQn/ZX42/XE/TIYe
8xQxsrg3B50QMJCnpZHxjtkc6nKoHws2Vc4Xm7Cyj35Y+p1BokRI4H2HDXvdyXGu4K3/sNSNiK57
dpxC1ePvKBAJdNcKYlqVdqxCPuxVGLjbZtigFtLOGb9Sl3Igt9AIlW3plQbBvD37/wet8j+AE28E
KKJ34WQnDV2ZB+6Go5aPEFycttUWfgAXHHxyfqP/WaqwB+TyOAMl/2t1lf8X1TWnvSxQMUf1cMBg
fsNRmMOXKfwKnvouSdXWPcyR0I5Bv69j+Vym4ncv1T+PRBEqIiAI4UyvAtZNVaJErT4IJMF1ztNE
+svU37LIWLc9Am2VVTj4Y3kgTc9FpG4DayPzatdF6rU1nKp5EePYK1ejBA24IcbzuH7IPq88OYJq
Ci9DsHlVnaDU/LpWHDxexBtHZOdlMD7gef7H2X7HoMiSNNawYLhnIFim+0R2K1g2e9wvoFlatc60
7hP7CX0yH1mCEXZGGlK25256uoQ4IipTHefFHl30MbBYHp39INRoNx3PdZSa3Qu8G3evAsEkKXpS
IyPkwG56Rm8fTc2lWjwjWrT/6JNnktpiJEAQo0782/7GrZAkRZQZg0wM2NYGvMCQO0DoUFPc2YfJ
h/tFlLMXYceR+RsNX615ThjHY6eIA/qQSq/n0+b2XJoSZ31iLM+q2jW55BdWTXXJV/9uKePouy9G
pVKr9zXWaIdGIqofVWK/eYAtrH4FGOu39Ape3jFvAngMBdCEMidCFOzQPaFd35Wvl876sog1SLkV
3TZxmq4KF6Fh6B3cMgkDR0xguHPrM/ic0qgJXqbygAua2yuBl2ojF8/e9U1hSpY/6Wb5pqdJGbtk
0rZKEfCbDAd0EjgCTZWpbkMPQSQynt0rdZAKNzEDWKAXH/vQyVYARJf4NWs1vcSIb6pt67Y4re2H
L7nhtXtgp+Ctz/xMB4Bo2ZGATpw5Aib41qU5ULav9VeE2Va/cbfTO964Vo9MDws0NLjar4rb5mD8
W8d+GFfeVgz4xS+4wjgEArDKnkZTuFxOYhItDca5DHkEMJGB/ZP9+DWgU3TcOM2ht21p6hLhIFpa
h013BoI9+/jGY81DsQ4owsVEzKNrEeUxozkkfuQ/eI4kD1KZhhkg2ErDvjsm4MCn0g1S9mJp4KtZ
Q28Dv21hCsCpRTYZNpFnbNR05UsRLnl/OIyM9hzdj1ZuGcxVKEsVTyls6P8z2s/Y5C2Nzyrmh8pu
5+raSDafMuR9wRjJFhFJCSC4IGK6PqhfRv0ZmKp2JkAsH3x2M/U/3CNSOUqpUTMgZTYOMNdnDUNr
l3uMFLalS++JBNNxynOGzBjJB2kuYvd9SdqERkrDJwXP5vPhj1a5OOS1OcWSk5sxbS9m6wJGRiQC
ynL87nURqoGRi4Vn28SCk9gDUWBrKaidQGIRIlGbqlgsdENf6M0+DlpN36HBc+err2ax5J210ePH
K/fWiG3ENUHKGPEDklv4ZHvKpq5LfkFkaJ4fcbxJLR5LE69/SYHnnfvFMEfgt3s17wo2KsjoWjhT
+l2cygrifTpEBjn95QPlFoHDkzcZH2wOiZJfu01TPHNktUaDKjr7rJb/4UjgXiNbPW5UjxPhros6
UW4H2Zo3qmY/KIcJ4ahiqnAPCAJ19WBq6uvdn9ohQdOrVk0RKyNYzp+PEck9MSTOTJRusZsF9AVv
dDeO3qFtZ6pVMspxTCqnkegIlLxXjPt/zVpNNPSonw35Zi1zSkXUlEyRG0Pb3mbZfdLEZXeITbwf
Ft0xRUi314nzpucx7m4z5WmjSnWNMkgCo8jYM7i2yaUye36pta3J0sFViMPSg4V9BjsT4sapnf7N
bNHh0U6brRspFb/P57hyiiVdvso9bl9Fq/aRsoiGlp8XWugM0hKunUDTxIWkZj5n73dkPBMj2IwV
HpKPZKrOKbI8cd7+CP5p5hdKfqMSJGoUE1E2NSsdIumhfvVdMtL2eP/f683xZL6LToVbfsECSaow
sY+6UqAeAQYDPGgCuIquUUZ0q38ZE1EuJnxIGPELdVF/XIbS7jhES7iHHU8xgdQblqruzCHRD1sx
bmvBn67m+D7cbVO89k1SYrUhhyJg2wpV8uSQ4Yg3zXj9/yeovi2KIfUFTPSyP4FRW57NcN7x6ZZh
1IWmchrRjbXw0TjxR2mYjKBO3Bhwjse+kAPhVgM26PspuDg4zjRgSX62E0+bptKX0uLe5md83EBd
rEWkXHIS/kF0ka+XJai8Z8soTgfJpUAOoPQGKureJA5ZIRI5LGasH5X5bLt809Lj29Rffl//LJaO
3FxAznp4+6whXfVR8UAOJ3DCp7tywvWods/vB4tZKOuu29NCaIwvAoo8Y+6LTpJTXUp4KpvqBBYq
UNrp8HBUN62cWzbQ3t9DPbkBd/6SfCda1f6cv9RHPxGuDdl03GpLJrO7TIoINB1Iu4GPEciu2krv
Z4N/eIcod4jmQAUVKDYfp70cY4VDGGSlaUrMosd02wXIEokEQehg2Px6xjdx3J1j8UQS8hpvaFO6
UVebkBwvEgg5mabCSiOkwSOtQQehC4jx7eQ/HGotKOXYK+gvWpUedeUuvQ3AO1bKLywZIoU+8njY
/F3SsCjGKG3TLtBSxcU9XKFT+/SlDk6lJVxj7f3HeBXjNhZBNmgknjZ1ciWECV2EwVP+bgPcyQPK
mga2Qc2gmj3+dS45WfJUAG6FifqUcB3Z8ZW1p9PLieDiKqk7SVeKHZOcNgbsT/EoNk8wDiB8jqB3
Vs9CjYiAPSY/itjt/eEl69/P40qm+Jf4p8ojksJKMfIwEGHQEqnMGu7tJQJ0H/bhgfFgTqvwh2V1
kIsG9wL1gshxhWjROOw+Ky+zqoSWvttRMIZ9gQF/xIeTl49ghyz2uAnJFLiOQX1bHYcpka2ht7Y+
EKGir1N0+s+TH7ObjJXvPmP8ILKHvErcEqLCVGrhHr8g8ZxSkvknM+Z03kLGarjqarF/JgNyydhW
rlPPfmqmfEwRpbSR9ylptJkfxbzUCrk+g2aFcdtmfgbpwDnLuiPxHRAI18J3Wv4E/UMkp8ATNxbg
0f8Ogm4EatkYqtYV9lTWsMOzex2p57IQcBZ7C03iV7+yTpb3cnhLOHA3X+2Lrezysz3t8jXtg4Ue
2GPrkwflc82T6kMPAJgCXl0GGwzY1WMg78UxldC966XuKgaOdEkOWageFS32TF5L4u6r+/oMa5IK
/QORAz4+dMu2P+FTsTQKTOIpCIa7ioiQlJJLziRfOYn2+evaArxh2UIdlg7DPk70pSX959mVoCXD
um8R3XwaG1bW+eDLY4b4Mm0xCs0sEWaRR0+hTpx1nJ20L0FCX+WLyBXzJXIScmE1E4+01zlav/NP
z3i20f4VehJ5flahCRD0bjAycHnmIQPPbZ6aoChYVv4LgXpUvECC0HNkyUHIygoXpb+Lt7Tgoqyh
63YhDRAygF24pgzg3cr+StzQHxNJGNF2S8T2aambYp1wlNH4erY9zFvxELr4w5rTinQ5JjWG6sdw
SqwXfxa0pDZbEfB0HOE+DoMrc6egr33U9W8Eq8tJylDh0Gi/3nhrbaF3kFZSyByZVy4q5IQWX+Qp
k67pLMCxSQcJokF5QXXw/tmp0gYkieMWTY07pUNgmYEgBHnxK5j1+l/boZK2dHD4Lc6P9V6SUuj7
zUlZGMotznxOvUz5oscvR6KPTAG8kVVjsMsdEjGcU3w2BEkxcSNnZVRJAHCsSBb3Kf26glQmS9QD
csgdojk4FF9J3J+x33xpDEeG1SGKGgbqcNSWLF8A6pJfvpRfKqR1Y+qLoNOYv1wWRDQKUkeYEVib
adbvhzJOTxIS9RUDjRkkRpyuXCyKPBJxqu26tKSMRj/Dw00tkbFy602kAIpUGlhn3PD7xLG/V3oN
Ve7S+J2+PKrorYROU7z7hO6W6Zp4XOo8t7PJwuWELSrtMcOLK22/g9NzTzbzitHm7G8z6VedCADO
boCY4MSYqHy+8uGJG6RbnVQdFCtL2MjOsPEZBS8VwjjBIFZHCjVitBlG9pcYZCCk4ozJWCXbNot/
fVU28cic1ABU+sAljafT4FNfDpCg86TIL11OF1gjV0MepwHy82suhR2YlPdd3nwETDI+kvFvRhm0
Re0ncyxtUmdExgSUCVA4MfP0qw+ayr9v8aODirxM8MOVT7VJ5SG2hCLZe2rqK1g2r/W6c2l8oAxa
38boTmtbIRkDr/aKYQXQAFZ/YM9pOT6fJ3l6zIQ/IKV+XZ8feACdxksag0truc2Z6Pl+FuPSHgtT
ub/vcwjhdQ9png8Tsi3x5/sUCgvEitq3hMdoEvl931xPd+VMG6Ar3TWhEGRy6y+E2FprvHG6nb4d
/4wc94EYqorSwsOsYLLU0B5dJMTHxWtmQTcH8jv2PgZZT/j9up1rUaGyPA6OqdMKMY99Rg1L/kkQ
vaDaiwPoqPfmZO2xI8UDOAlMVa22Jo+i1XBQaWiwOcmJgzChgxyvj+dxAqIsmq/LeOYHi5k/xt5Z
jyrjSX5EExs4sBWqaxY5GGM13D3enXozuqY/aT7Q+NT9izpKCyIXuktDZr+GczWzBcGWweQamNOx
nnPIRK63AoPzBuV4e+vg5jnAok8aw6m+96uzcu2ZygzDFdLloDcVQaBnt4huOHUTJsMPwX8fzhH0
/lDZTZXe2v+Qo8m7AxT/1SXr1FxH9zeYTuaWXmx3BQibSXXaXamVtuZjDaXLQicitNDMIC4cxlT/
+ZfrfAc90r2U/OyZgDLKD2dbnLbIlEhyayHkeXsdz9m12S6V+UtX8VPanff3frgUXL7k77gszYj0
fLUmb2KLVY7NuAVvtEB0BivVVJUjUBiNHU+1/oAu6lqay6If3mGsDCFe/7KaQ6Qz6Ybqj826NIp4
nQAUitTTTtFzG+kvIVIZZJS/geUAdBa3diDYYGhJj+1yNSNbzQ2j0gIee1trP952z3rBkPfTtGac
hNzken2n/hNfBD1F9SBBrw+G5UNNzVUjINQDdLXjbiEX3VE+9zOsZEdED9dts8qYtvwyFtGwbrYD
gQx+RUCapEQnc0KCkHVQTCbCngowlBnXbnDfSU1vQ7DbY8FVHwd37yYKRdHQv+9OWZcC7x862RjV
gEL/Du/ri7F1oK8VqzrKGpfG3fNQQpX+vbA9E0UJ14xLQr6JQ/eb7GgpfJ2hIDNtiOzKTUVlZOKC
kUo6oRETQJfqAmLCqaJd+MHXjGiNmRoVyslslyloBBW3Kxucw2R4noILaLwf2ngsyqVdDVBf083w
FpwHP4mLvnz7amZWbSoUuEeW3QEWoKhaa3erE2jU9nYySqgS49CuV2C7sczux5s4qQCHlqCQMx/K
EEC26h/S1Hpf12hIsim9gpYXocMiLH7AQEOXRF0RAZGJvsteDSSFl++Jqbf5sh18Jmwmtql9t30m
VobDhtmkSOYix/DWytLkKK3knitgl2DfXZdwO42KBJpEhwWWgs+44WpNMI/rNE9x0KrA82TieGCE
mc9J5NXl0ehTdJGUoJd93Wnpi1ilg24/WphElfvbTHA2yitdGcpWOS1DJyNWddfUL35QuQpGPGk/
WIOvxlzQymjNTmMr5fw7xi2JJvddTR2h6OxVjR8KDlQactk1PXnqvPAc578QaYPZHmLzwO0gkMn/
UNeMjEwV7KkajqYPRAF9rTmNIX/Em4JCWyElNPp5V0Zwybq4pITUdSh0wJxxCgZna//DZSRqicXz
uAwlusifFUhgj3hM+yP5JPxv+Gnv655hffynjinRXeFCQHB7GpSM9ZH4XQEZHTLHHz6RpmidHhTE
wlY7nq4bu0hAJ1MecWluHp2S0Ja/AYZzA3r9BtdkzXZzky5DrGAix1LazEMkGrSKSs1f9D31qTC9
ZG1m21uP7kukgR31jri8ApxOsmoOefoZhhsIrVJ0qYqiKSSRZxq1/Qzsb4NWgKQjMjqdFq2ft5mb
Zb5gTVM4AWmnW69/4vy6zWA8hPtRPTGbh1G+Dl4qFcKG2MQOh8YgYnxhCP+0IlH9qjcFYb5wevao
ycvaGgn7JHxFiA0j8TuPt2HKXqZmS/lbIbqL6K9DQVVsV0y4nfRAiZzJuE/m3ir9d+RH+zFdacol
SsM4dCHpNnUuFWKgpLT15MdHriCO3dMs9hTFipOed1eU26zyMWjbDe8ysf6CppSQibzOKtrLm2eH
4I10kxGDuOA3IqUxbY7GUDwAipemWEsCu6Dt/+E5ETfac/mmhIcBnsJ1RyY7FYae2BbslsUWvx/a
exd235+IypwAydIDx2kyrx0jA4fKeELyhGOnWcItcsk+WgicHBdMEwzuywvCXZhPpCq1R0GH8Qz/
j+4RoEm4cjF8RWuukFGlGp7dB94u8V6GTMqIWZZI+Jim07uOClQV8DPtoci84MqDFdep06R31+Ua
pYAy0mDPFSuyxbk7Efw8Un+lhsJEtR9FV7RVCGV3u3yMZYRjZ16B0vt1wV5+Py8kR0fm2AfteJRp
Z8KVDPt59zZdEEobaqlAfMwAWhDi6wIhDGLCqodn6syyg9p5qg45IdE0xNEwGgks5f8Wgc9eAGtP
M0H367bJk9PoB6W1ED3dSqIx/JkV8Na4mWskbWjpfxMNYg5SwVbG4CX/+zYYZeZixhZNdwP1mg2b
/czCwv/VMaiElFgpUYa5pP4bjjAldxR5quTIEycrICWjFHVzKe4qpNcGN9cejdCbM7KdVb7NWGKW
vcRLgzcyhSpOaxAijnokNccTY/Hu3dHAjsOxU7PSnz/usGpyg8zY0mWJkCZCl9FF78CvecUXdW2/
anBHT7B9UTe/XGdiSXLgktaasZaGn8xoxAnCiwR+jw+uWv69oLLjIXKZbZS87ksAu5cbqd1vwN+s
7Jj+Q3R4DyNt413QTMUbEIzN2qqYwZXjxNTSLMFnQ9srXXj+OunIlZsPYa9qIEexPsJKZYrrYsd6
yqrqnqYKKavZp6FZ5A4t1GdDSxtIhT8CV7B9xBM/p8DR3Y2ceMkusCnELGJoTUs8tFkOJFe681xx
5zBWNpYnpr3g5cd7asScjePj015uBVwH7by786XGMrWJjOC0fyumaeTkgLq7XNqRM5YCZcl8Lywm
hIzU46KJLuGWmE0uliTfuoVb5Yj6Nkj8iO9s3sCewpSq1Qwapkr59H2Di7Yn8hssTrNla2eejghg
0lLkkwM5Dx19XnKO6UyyWbGzoiAT93fHRGx/tUbqVbMeq1hjiZ15+MDk2jyNL+sCBfAEnzY3RDyL
a/k2QqkXYdt9vxFN4ZlBG+6yiIEDTMLeIjMamfjIIUR/ZLA04bkn3APdMLq2wPFXrBO9MJWza93O
DNiljA/ToMGSI64WnZKPBTNT2GbZddyKh/ldAQRgWI9Wu5RUynYNA2NtWgr5XzXKVl8a6UcN1NG9
saKuEpzygkK0vZYJrg5rJLC7cLmNtaQZGSIqC4NomiQvvwTWTVWkzq/W+C2CCYSiKROBQ1D3ZXFk
Z8wOAnX9wwQ2y7zYUoAXoThkqrgD+siOsP5fWFXuBuHFr4KpbDXgIKampNuPyp3MDjMed2rYpO+f
cNjN4t+EJ6hagen49WukCtt+b5kfZhmcRL7uJ8tIFjXxTlrPRav9P8p9QN6xLUbqdSFEeQR2vCQF
ItAcylVXT9gYX635cvEk5JSgn4Rw5v+92Gq4XqsUfEmniDjDCI70IO8SPnWA/10KfJX6bPcp9ho4
dqXfbo329ZaxH6sSWET8hqOMCTuiMJGXOIA2u6OtZpIPkfTIwRQrXMyJeOPLiKOtqxSYEUbbM0QW
Oi3E3DbN18vMdi7HSp2Wv45VsSrxOzVDwqu1cEkwvFtzq2trxWZx0LmxgvAuEBFqCoKfNtnUlGlT
IRPHboe0Fp0d3EKb/EBs2RMdopyCw8LZWtyyxK8pzISoJNiIunD9iO5dg8xaqscfC6iF6qtxQ1yQ
aVYBVfEK602LXsxX2tSYtPkuFvFlhOGezFUG3lYKTVlxIO33Fc9Fr8bS5Rfs4Bzq/kMhwRJ0K6os
XqXcapnMOv210adMcrB1Gt/OCt2at3q+PbzCfbV0seWL6HvMTIRjqm+2cc1AX3T3muvDoXmv/MZm
eOTifwun9H9kxvQixRv0iMPU78hEvQDRKoxwaEJcko4gAZBwzsCY7BBPYTPreUIaJ/qILEE627xx
evn/CHmwBXh9SR/EtBmrVXUq6x7TDAh4LJbQU9BUbOhubbgOT5JjhkarhwTMle5XQynQwas1ntgA
LlkCy3gF0yxeDOyqSHd6j1IFUIF6JPxQLsFVWtbU2jdQkVGggnsJZcLNkDC1fWTtx6He544uoXeq
EGC/JTPAIWQpKXXtSHH52U3egXK0qaMzOaoHhKyN5ShYYtyZGukus+RkCfuGSrpcWQtm68dLPXNr
gC2l6Mjls1dLxNCOX6+AmUdl40Piz5Vx/pyrOvmZQh4K/iWcltdG1whafQx9q1NIS3vGjh7p+Pl0
LJ/+ZfYgRiH7xG8cv/7hcO69/y+OODEuxAhE4QmLH/Z19+MZomSVUpqfans8vpfjbpRx62n3lpGO
3p9HnnEHSoumBoRCUHMKXZLQhiFCResn9ow8Ik8t8Mrq0XrKVEiVDqJFwyeRI0SlKcxRXnLMjg/Q
EW2bOKQqpkPjX704Z7Sd9qt4Ui2JN8gU1drmQAs6sDwlvWOsTTjlLFQrcMUu+joiLK+dR2QMPIPI
Eu2ivrvZlMXpNoN75uBdB6V8cu/dyCEPgZinuL3ZSTKD/MhldvSkIgNGvrfdXmkpSdeLdpzG+e57
HqP8gIUeNG499Ham1hLKODr0nejm9vGtDBp17mbF7Q9SOkvCrWsbDha6J8vrYQwdzdC6i4H91SvE
vc09j4Oe3oZ/JDsLjSVyLAp8VLz3VxjNcmwiDouziIUxfbDw+2emXKdCxFGho4LXDA/7l1+vRUBh
PdaDpx6A4Qs/BkxTDgfBYuQcqeiDpmrMXF7XjlL0YpyLGJvEy+QOAAsg1R+Vo7hx90kRMfcpyrGF
VMAd2Lm2nKaLUv7h/VuEBhLaua0GESmWKTaXmi4b6d4dK9YEPxHLhs10yqdWDuZ+ESZErKp3ku1n
uTWj5XnFMYw5PiUmZvi2k5B3+8vYCUt+cbh/fGj34T11qa04Gw+/oGonzOgvWh6Peq+A2hqBPWM2
vbAiMnlfNc1fW6cFmpoYvbzM0uXtmvfJJfl3zPP+qjVpORkfFPp9BbbkG/MfLbnk0BgFboShVg5f
P1/iPgStTRuUAnDzghb6tK6b/EvyRH5fH+7sIAUBFo5+ejIBvEM8n6hF9g7Rp6cs/TPuHwo+m7qK
7tuoNKHAidcujyhTFpL93hFEbSZgVNFfkgbweEjj/UM9Twh1SuTxjOizGo33dPnmye1S4q736gAJ
b5HAwxPjO9OwdSFsJ0PKcosRZy+u3FNLn0onzaqZH48LY0wYOoy4ZxZijYCeFCFafVsxwg78Vrk9
gYGHlf+3FrtyFyOgxuvRyg==
`protect end_protected

