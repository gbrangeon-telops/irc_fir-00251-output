

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MPaacDM0TWg8wcifAVW4jEGylx4PKrqc4CLboKEk0r6t7KyfUnirQwQAphZDsR83L059CNEzB4wD
M8AKmBfOkw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XUT3zAfEi3anHP5UZ9Q64SRw1RnMtcFX7nJsXqsc+jcNnlmbg5PdhmwV7UaFs/PrWKFdgim7UZCy
o9NtHbXd3iHyUEXXZiWfkC6NC5Dndoi/rfKSxw5AtxtcCSaJ3/cb/i40IG38fEOD0mldCmJ0WOZD
xOW9J2aHwV12uWmmUBs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5hB2z6qFvCHrfde+xOJHAAm9Y4Zd5X0rYu4ngUzTSYyHrr6WAc0PuLxe2Zog3gNAv7DFoV1y/Y4U
F6T4flnTjzAqIUvyAW8+maZzCAeWDi8VgmeKHRbLydt/JWB9Ri7GcOoofnS5/hxq8wRCMMkoHbQF
kNzxfXz2j2QXU8RR6+E7pvqcJkK5H/P2HIhS88SnGwppr+eD2lVT18h0s/QB43BH12kpY1JIkQU4
LOR3Ej9QoPTxmx24xAodMjc6qGME333306vLcWETw7evLQ7fHCoyGS8qVr9xvwEOuA+HtAnx7p26
Z/azE34tKzoImCmpb36r638Bv/NLBk+b7agF9w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n2iw7CqdgxuZ5kdEH+pm9NjU5keAcvOSKkOt8pim3KzIVtdYby3hWhnEsC/F1aUQ3kkgfoeHTv/o
nwfMP+AVXxDoH7hATDu0iX0A8s8avaGhFp6novk5xXzwMVnGP5Rbk3GwwADpRNWqzKN80je+JhyS
o3J4z9hQTmce/KBAfWo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sR/mTVuOveJs41YLuqwkxNe6mc/KV56Pt/6c0cIYmcRhmwLHOU3+/VfoPpEClea5ISswKcgmSmEA
91cZp5XMe9E1MxpJldN5YBxK+3XVJrpKIG8b4LM2yC+ZTp/81AZ6CpAKQXOcZAota3bpWOVB7WQt
kPn3pALJ48nc4gaIOk2j5GO0g6BLITkCLwe8Z4XOzYZAEaEB+5dJ58Q/7AbNKHr5UdGO2UVVG5Oo
7GIt9ETizL/sKscnCI3CshbxwDQPtnh9/CAQY2Ci2Oqc2ptOmylUrV0jpazJ/ulKvyLMe7D7sjb1
BOUUkYAI7NZU4AkYW+pW9jcllm96HEkuSjkTDQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50560)
`protect data_block
I5BVF6CLhXVg13EehYknDaonWuprp8Wqg5T1Xw/z3mHU6SfnkyvEfFyO4nceM5QwKUYEumww8OLI
xx+PDSdNREPUNIm1Wj7/+0z5AYOTbAX6eFzJa+Qhqf4GSJ/ssUEaHamzurZUajiUwKcL12AnM4yH
3ZVacR7VVIdFffZQvus7NNei9E/l8e+77JDvF+fHK8vgNPEyW9i+Pd3tGRP7QYgGSDs2bX7N2+uJ
+fPhFqMkgrDTa3tDT8bOGmXYE+fSb/tcWDCZ9BcHrdNREYKTdCUgDXO7usBHFtqPSSBP7DDWxmZh
Ka8cSxC46xPXH4GCYIWU4W/8Vhgx9AA8ZP96apDSur94yyQSfIA1GGhj+O8MVKlY/jFym1Ifktzc
MCNZ2DEUILZ6lqXbC7ABg3/Yslg2kRmADVsP2O7PEyEZcBsf5ble8Z4qDD8w3eBeKp0aIn2l0fFc
efkHZjMiZxwB2Pf2+kR+RFHa7FMLm23tU4kj7AgwojX2qiUFQTrH4WnV+e+O1EDP1itKMaOdG2my
WQXoGUW4rxXHDfD6d5cxkFXp80PcppVvuRihlLkWhTi9VpBebrB8/RohC14VvxaqOlS+Cdq9eDJg
zNJ+RJ4X4GsAXDKFxdSu3dqbhUQJuNpvCO8pLitVOhcP5+x6eLYLNLwWJyq04Sgtaldt2ESi2xYT
xZ6mUTlFleoWJmE1/BVufe9PRlUD7xOw0gdRUV5elsdie4FiBtUASYjuVeJb9mpirUG+cSOe9Be8
y0eyiZ5CBULrR2lloa8BfaKP349pmb+w2mSYIDhbwYBrJPj3OCu9vttNxrFsi0XtIulsLv7wcP/7
C/dISBxciPAFFDbuyYwkN6PvS3jmgyhnMx8dZxFF0SGMzNnJ+TGeVvE/EuDRI0xUNOJRZiRko64s
NTMvq+FtEICe57g0O8E8XJJGISFrCwZoU/SllNzGPEhGVqnfbpZiMMeBxT/eVO1+l9d7RNvDLQzF
R1T6+MCI7Qff+0uteY/EZwsAje4QPSLa521Ov6G1TIc/AMWfeCFdwFi4w53+8DOsHZxq6A8jPmnJ
pKBxQb6YTG2QMJFfGo61oy+zl+Au9I3BSOkfMbgo0gcvWeOgGsE34GPb/wvb5L6P1WLZfvRV32Zr
908EMPQm3jTxLr0KVAtolrJUTnJ50j1gtYZE0gmkY569eUEiFSXjEiSlWz7nZ8Rafj4eK2I2MJoT
SSZrimxOoej0WObksrh/p5wB1dhI1QGJ8qH9j0Ayb93jsrvZbzdFTF/aRJBAmuTCH1Y7ldSsAZ2r
Y+ObJv90PdMRYdZzWvIXZAxyQ/BfTew6UhWRHWpLdYxtuxKR9B/7bjkmgAUbZ2lxpicMNZALhoXT
fKK61EO7IVHIViZl6vwBwRgasi5OmiQOU+jDsAVH36PSbjQPDec2Vc+xmb4fAfsuCVp7cNNbNK3t
7Q371WTsjB4EtMkq0rYsG+7J1igMtJvEMkIv8f3N3Wev6Ym3722rMVNPj0TgGrUckz+Pfo+LF4MH
2weIyyfoGe2wZcup5unhI18JwLU2pyYXF8ga87GCgDrecjqg85bIrQM/l00gMKcBMGMTqqIi/oiR
3xvC28HdfnDwjcomRaJeuWAHyLdV2qbuaRjhxRtRYsWNHPGtr+AJL4dJoKJ92CpVZN1qf+k+oCwc
9zQiA+1Y1deqwN/xaLFPLfCZuPWtDRBR2Cuh8iGIXFJGLLIU7oNf/3cEDppX0xkNMRTYoN1Owlju
iy1DI8I1PQlnmNLg8Rhnq+C2c1bbqjHPrck0kCfhsZvT98W0+Aq8cNfYX9OJ4u8NXKSDfqnB9grT
LNMpJqhxXFOPlsMFOqsgT9beF2KUlM8IXXdLA2nKqs1ETSqS6wMqd3468HkkBSx05OfmcaihGoA7
sCC+Dv1/MSMF3a6HrfsMi85pyKo0qmefjB8fWEnKR6EvTUmfy6c0Kgr/MtBT5Sdlbn0aFcAYbqVQ
+/fWJ0EdXaGCiTgrBSEt+UyJl645sQO5AisA8hXRUBEzRBEKBU/N8DGU9YQNZBmBj6BTFZ/XcUGf
XSMjWgs/ouIbg8gV8gk41KrHu33YF+2QFsjzA9s+cfBkQbb6objRFxT9WctDnPq3hCpvqyFFLe1B
tLzXZrWu/3sEnb/95cweG5gpfSeZTcq7miRjRo3Js7Fj/uXnOPIplTzxMroRyIj47JKvQdI2wQlw
7Zvb3Vd427BTHuLF5oaJZe4PSzYtx7/BTkjhW6o3GbEQchLllCte9Rmb/7aDjlXUkk3gNFU3SPTd
RyzLuhSujoXDfE7sSVoSCRlC6fCmotUU2isLZ77nnfY0xSpexmvhQQ0TKJp/SHUeqGnQ5yXfEXsR
J1BolDRmfzLl+OrVEFfhdmpQzG+RXoW06sg6HAv5EAfVX4RmGlx64tyRkQS59ZUw8FxSSSQVUaKL
LuZCgfIQJhji88Cbbe6TiFSTiVazdG6M1gT2ohBQFx4wesk2odxnlwdLll09IzR2k+tMFhlivYZ3
KZgfa491X3RAcwt9j/Z8TEry6TkSjPIs3LAxezPined/r38ONAHUJi7w4pLN8trvRrs0Cj9l+j6/
g4aXg+QSOcH8Ci7c6aaMur613d7G3sO1lMcYidusDghfBzEpMvnF6iNNhl23QaKHvJN1kDTx18sq
A7QpDRRNmdiszYY2ySXcAJvCIMXb77hEC4uCS7GVrbgeDSLZZNtL9qhychTZtDqXWkOHDYmVDIhT
YIONp4rGzYjBNDU7jkWOgQQC5mDmEPVZ8Z9b7qNFIgWTr8gq7umESaCvkv0+3sNOoUbMHOTBqqJk
oS0abTS4p6tb2oC7tgaUWgAR18gGeEct21eOm+O3GEcly9MhM5Vy81sviX52yqv2miK7Bg7bRuhe
l74m+iiA8blg1dJ/NXc3DLtDXTCz9jDaEJ+bej6xxHafz/dBOePaJ7sc26Yyq08sMxRMfAkN240W
ieFjYoNC3moD8XUGsOIQn9qHanywFnL8jV5NxYaKDkHWf1imMykgULYvjocwa+CZNz+zqaFlZWVX
yczF+9FAbZ9xWpvQUTIR/jy0Dm8Ymbk3Eq1PpS4ZSHuh6xchiOsEFdFQfOXyMJbmCXPuCJzz9Ozv
PClv7sCE3pWZUj6xQPuIBpAIEZAF1boQahf4mXJ+z8G3QH1E9C1QPH+MwAPJCQ7MRvs/6g0rt4FG
rKl0ZkGvlOsJmq63mMtDui2tNTauq1VgIeBmDheo1whckTn2D940aqkMRRTl42atRsEUJDcqYK7Y
IoQZ+JPobiyddJ3uAtYBhrvetHPoaZKKumDWRPOdUqONmyGr/hsMsPg8Rq3moe5E6M9NK5yeu8AG
+g9DsJDGwTFL2jNxi6RDNFm24Vyi3hJNb3DqifgKljOsH6HgEVffGMAm6s3u87bYEs7uTdVfoRYO
zZsaGINM8D3HYDDogt7BHZ9jJLTCu0lygG3Wi5MNlaYr6SN9q3f4gZEvT6ldNVopbVAujweEnZes
gJfD3ICCSMO1G7+mciwjaL5oLM9QKYPKR52iu6mIRW8aqUXkQps3PcRYDD3FqRW38bRJfkkMJSYv
V2EDWmji2FuqMAuO2pVKPhhwIIha2tYj1f6CNnRhW0bAydxGG7oTisZDRNkF14EW+N86ES72DYSK
wtCDW5sTknayFWtoZRoNZteW0OKSnNKq/XGBPcGF7hV8dNJNEyaaNabWcPmoZ5Xpksfal7+SKqRW
EqYUVN/QxmrqkuFIHR8QqpFyO6CKzFXzAe5e/VO/MU4MBFPXpMgYVoTE4xe8dtCuTv0unJ6LIc8V
Dla2b0dNE5rHYgjTYinqsX9DBahrtbsKdISjB8K7Z0mtQDI24la5PhPv7KpngrbPbHXEUrrW+v1x
JSPpUV47fqzXDsl16nQ3ZIBTc0bEoL2N+XKy5JOyqY/tg7IrMrYE98jbwo2MWHyHZknnFc/8LQwa
HdR9WzzJaaYHJd0LnRGtAkUsuBLPY8sOupa/zPRztIwcyYWaUhXAIJ8NtXkp9ieiODm6oNYFOBxU
+49/pnDI87peTB9JL96eUU2zmrte+woNihJSrIEwwzx9R4EIZ/fdkcwmagi190n/zeSZCbZpsdWd
FeyyOHCTsqN+KUt8Ge52BdyYikc1qtzdakupgyrVdggyX/d1g1iLqcCeg0qMydVim0quLU1zxK81
9mShd+CHOnSxLlx2cN0V5or3z4wSkKdKQWVODC1XSYX9XCZkpCJKFK7IbebofXhOfZAIIqSQ5wA2
+Gxz2RkJyw/J0cVHxa5kU0mOQpKnk7q06pFmsuEtlOZ0u0HlFuJt+l1nWf4tI7vjxQOpVdCPLJkJ
zic24HTxHmbcQ+9esKXEl8rgSwjHuzwnqKbB2Bwh69Mc9uBFakJa9FIMM6CQ+ieW4tvrggrK9SWQ
bP2cJGzKUhx9v65Cw2vzqhmz/VrHtOnKA7J02+gbqa03hSZWhUmastUDUzzN1FoHKih5J6gxZy49
0Aauk9h6b5gefZx/qcBuf7S/EutJgmOrbR5QFm+w1ybehQebUQZNtyAlDLWt2hsfyriK3K4HXk0l
K7mLqTFyrj3ZXaXMxdXQtsGFVaFQ3XtvJljs2KXi5nC7VF9GJ63rb2PSQWLCjL2BTK9Czf1U1HjL
XTooYiYYsulsiA0YhpXDToi9k3bRlpZ1WSEZ5XEH1Dn120imSjEZlntRGUkyC2bAXzi9FWAd2QDU
g/X7Z5oGSYPqASyx4+BmpAcFm8QvLIGesi9f5VwAFeyQsAzSkzn4qtGBJV7tCOWVvfcggjSQrbwG
xORK2P/o3oGcgK9oFiDUI+w5K5pwzCKdw1F+8T9tMTh3udwafXjT4xnQjqU+521XL/RxhZz1RTym
0lsSxjT4zZMS5xwN4g91zGJIhdueprZy4Swua8yegLAO0OpUnFz55zSGcoNNMhoz7osjP/InPqRD
ZQ3oq7zapfxolPNrk6PXyib2qNst+8IL1mP6LMl8aGSYzxWXe6lzAoaKfcsCnDuJ3ifPXKzDiiRG
Ke917OiZIcuaeVdWGb6G0KUjKhf6RbvGUMjSzl46srRIZ9W0Ju8l9I/wor5gV3byIKgioYttrdFQ
Ut3suFXlIYBj6US4GCNiE+7NAFDQ1cHxfhKl+3r4m5fI7Dk+fEUEAuvrcqqjaGmVwl8qtQ6R023b
kk4rL+rXqHbn7YCcksV0sixVrBUFhw7PKAZhvgeEPWWOhzRapYscyXv034+cuVwd23A0ZgGc4Nc2
mpo9aliELVqQ7RQapRl/mxoOSva8BSDLelxK1tVONqTtGcWrYs5hcYkZsVoQOFKOGjtJk6NxAKtq
hwjoZD82JC5iWalbOmQJmjqKZsnuwX55vcGFmRbcLk4rChNn5BcP78UrvHsAWU4zAM72a0xEVl8j
XsTcEDCyAzfCVdBGR0rY+xxKDc7fVbgQuY3S1SlWdZZ7NKKIIJucQARi/nnxgD0XODrUfGP98QCl
DEuaU6CUr/Emv8qqNs2JNzFZmkMM2GTQWKs9php/XLZYaBPGt5a3IGI177YxG521MgOcJxqQ9lqh
Rm+gfhPmRTj/0KTwOmIYnORTZTa7I2LUJ6ZQVm28+DGyFN3VAL4ny3hHWFKzhJW4H+0PAkRQChND
/17j9AlPNOSzI6rztkMbhHLVsAfP+e2T4tKBrdl2zOzFH1j4SbyWqreDoiwoUsccLw/OJjCgOIQd
68GaWHDG49RrtIBfEvXLnXjVdVqZAMy4x/PYQ+sdPRZULgxKXkZcjGhEsnMHQ73fvTz2c4i01P1n
Zua/LYLQ8dxtV2c77nDf4Nmy5qNb8LEBtGqjzDbx1Zmf/GBcSjw7aS9+bIDccnuzyQ3gS1iWJ8mY
Ni22YrOzn1EcwYImaaMza5l5bRgnSVzNRXg2gV6dox8StTK/hSAfHB3nx6Gwue9YoZ8qXmCm9eqp
Kc9j8Vxwg2BOt9pxGd7KEtRDH7ruaTf+n15Wl/bi03yb3CL/bXoB2wynp2EhRzGeHy25uDWrkjZF
aX5h/cQQsnOYlAHszB7nPxKnCtEIYYnEEn0/eNIuNuWXwT9QcqFXgLrgD9P4Bp9F6hXvGZPEcoVA
pF28HWEwt7Mhspd0HQkmnFOROO/uqQa0H0b//TerkhxR3lSj/Zha05YpGM9MZsRlKbcldBrFqdFs
ecpkLgxKa3loVwb50XrCy0Ku/xnWdlNYm6qGyS7XKtQSzJTYXM5rfGCYebsi7POAqCQF3wzdnZ/9
cUq7v4txk6jbEmNQXc0Ov+D+S6JP7FnFW75i8AQCXhvzGctBzSBDPAyl0+dxD6ZMbyajc1fBCWXR
uBY+e4r9W3AhiIiB796fFoTB+kHN9xLg1eodYwbaN9rY6BHjuPXpgMB+Ud4Jy6IlhgG3StZAWRuB
41L8apyJn7V4VUJ6kLbQwMY6/0wGdYWoDa0TsM6rPIpnUGDOzHFHd4uLYIGegUjXt0tptAOx9mK2
jgIWZOzeYnhJ+e0IZBc1863KZL0SpXwZOveUbVNX8sYruJG0QwN50trBYmcuJVMagnSUp4EI71d9
nh5Km7kbQ5E75EssMgV+O0MO5v25e7C4dJ7H00ZyVztgAitPj3DgYfxoKuAxsUvqThfzgZnP1LTX
L5Qa1vTtqjAO5kF0ikvXzrtJyJf0dI68tfOGQAWpp/GltNaksk9i2T1ivhYvIvWYTjDOVg7Hp48m
abnfhtg4VMCJU1sCEiJIX7G3+SETzZSGf/EmyAxGXxJhv5SM+M4QCufvuYO2saxlEWC3l9r7Gf4N
pVgxlS5yA0HuHDOMLQlnwai1m4MkMy38SkV5kHQtJf1HjPny+1UYfWvt003oxUBJoD2pYZ2VBn3z
rVCSPcBXwhu4U38sgjV6+0Zj9GxI7g68/ZKE20uVucMUe2HassD9D5WgDeo9rRKLIOhYpqyoGYn0
zWnk671khKcz/oktxDyOxGLsZwo0KdthK3dBTc27yuQYjFFL2b5iPgRGKQt3jxJpARpYsDAhlWoO
XUV6mOzJxq+kVYNx83x2KO9YlVL7qQ/Eg9mMmpjUuhepTPgrClJQBsT07n/feMNJvUfaYitgEbUc
oTeB1FLrQmxbhB42dnCaDJ4XSe17ontL3xT9d7BCWkjbXgywSY24XIbi56AUuXvGZDdmA0yTR3At
a9qKaxA4i5CSOZ7PX3sXUYa8AqyD+2RzMGlwhZP3+LNctqDHLFEWGz0+v1MNTfuE96dym5MV+tbe
AMb9Bg3w2YjMaH791rkyPtwlfzPNZdVdqjFdcIxO2sOjsxPfArYopbjdckg5Qe2oTA2LOhjzl7J1
KrjfkH+trSKU8s5kiY0o4wb6aUwpbp+zNlS7wHQ3egRpTYHRLitmGOHgpbtgqmHOu7RwPFC4Pu9n
5SW6FoDuGkC6GUtwWlInNPOTbieR6qRjgxrs8QsEw2wuv4wfayDro/119ID4j0tws6MhPtjp9eKp
F+LanlcL7b/pD+wUDCS1H52eDK1l0Ts8G2hRPK158CL2ipnWTPKsknf8CeZ5AQ0M/AWCxbqGAgpQ
e/A0eDy9UO1esbCiUGM3gOyLBGRGGAN85bDgQHz5ZUB0WbmxS9ioiQg/tEJ2/xHxAnbgwRTqkWx0
tJZlhl2oWbZLQtbl3hFSkTl2eQlkdIjmJksSQrR2dMcibmuxKLDKMV49HkvK7jnbma/O5jFDqjby
F7IL8jtJigoK0dkBq7Mluz0JlYy2hXdDukH5rzNtCVhZOHXw4Qsb3g+MBymxXw6DDjHHr9ssw22S
uV+OKgzQltuDqwKPVzLlnrMuTxluPvSJy+Iy3ofCObIy3vkMTC4M4FuVk++eAQnvMvbGl/l22I/n
CbT9TLHA9DUXFSb3T/0X5E8DSH2kdz6urxyamCSBMPIUEy8+V+bNxqZBVekH5f9H9BlZeKG900GQ
JYm5lFKxeTv5x1iafD1nV2xZvWeEQ8FU4jjp0xrV2CoV8t2eHzsXJPvlCNIYVxwVSt4qQE3T/xQ8
+lZqOJ4W/TmcvcKJ1OWoT6PP2Ig9L+d3AwERjZNSrF5bwaSXPJl/S+PgTX7+Me1fhdOgzXwGg/cV
dL8Nkh7jU2BKt2hb4U0NTsGCy0X1vbPNSH+DGfVv0/eUp5aCW8jjPDLAFiuw8Dacmsbkg7mkEBMf
KygPx5J+ZTizAOz42Tc7HtGYTCDmRVLn9W0dltk2c2m+KrRfbwvitiP4BZuP5tSpgPM1UpuVJvGj
DEJ/+j9h/vABQoZKxSi3Vu1DHzLIwT89EiW2uMot8LqF65Ut7ClZh7aw2ILate2doSO8E11g9WRv
2Dnw8riK5GcWJjkhC7SEjRkF5lvBJOaETDNPDoVqoayakugzV8ULiJ7nkdvvns4FK9P7ZIB8w4lL
0s9qkb2/gIZxdsLo4TDavne/kwRkFuqjuLFGtCOB2PyrYZOTRXJeXr54QfI8nOs1uAti1kCy71am
6zFf85EXBXc7GYZ22SZsO6H+rIif32qIqyvWgV6D8UAgc8KJwfrvc0mO9Rim76MBz0yjQN/oVsy+
kgYlRojgQSrqRiLba4RqGXwqJ9raw5v/SAz6TW7b4vYuWiyWvQzCLpPj2A9go7f9vjDtZ8t+loLp
0WsjyqWZ78aeB94Z/N/UNnyOJd/UepQofLoc55lBz0EutVnp6163s5p5iqhhfRi+h+u9ppZJ90/P
+HnuUs7lyuu/wx50Sow+jAJCbfKZDRqquvflfyCjwRqHAf9CyKms+kPbiuNX0jtGjrxgslUcSzGi
+4/3yh3bC4219kVCVS8oqeGqycV5VlZjX/xFjfvM3j3aEsVfDbj8bryZ30Clj/sl18eFBC7hSlnv
GW4FdSBWhW73jtrEve9XjaFT4y5amHDhPSFLQgDcmHoiTorptN9/IZUmvCj0npmYbY+JGP9Rbfs/
dcX2lXz6s0VlVSGIQY7o59RA8jx+YcIM0iMcWj4ChZTzmtXrWi2JQ+E35jeionPIxJucrn9QQhSe
fXFXHXLhtZ+948N3poydI9a9nJmsG1lOx9v88MkHlyXFuSyjNNY+8igtUrSHGlfYtvS/RjlGeUSP
kI+Pmaqn8NvqbGZ36nLZjIxwOH08UKRnFKa1O7Tq9I3ZtkW0DWiUND6dK5g4i2zB4YyTewvKdvjq
gbbT6ftviIrYsZMwsyVqMYmW3K1qG8YSQT5coIZ0n6KVa2hyz7gmhqtglrxVlpmP9zBvQcwH7Ood
0yyjnaj/Csj8vgZJOkIzuP/Yiw9OKvvGlyQE2Xl9038zX4NOUZX7xSdqgJBj1dIArPUJHKYWk2up
oLcpbSNXFkGjHv7t8cZpWIzbRcpqr7pkvD2E9MHgxsTv1lU2+Q6rz9elELTeKZYj/lVgvAQ7dqOy
zOUPhZ+NphmCfCUZP8gW5qGNWF/F3vHN3k65303y+W0D/ez4XMmyILewvGTsSu6tkBMJeZVjnbgw
xQbi7WqHk4rt0V8Hhf9fRP1x27d6IxAwa88sosxWUDqa9koI6NNV9SDqvghSh3V/IBbOsv+bshfc
sRaoA7VMsFW3Fn7in0KSHSB9MyH+Al+v4eHkglFKhjd71+4dYQFnw12lDtZ2gSr54IwC+kgFc2KK
4WgglaDFXmEfCKJd4sKsAvC/79Ma9ATG8TztuJIrL0qsVtltpWQktubqbiEfn9ZIaoEBBIpUm32d
brK9MpvU2HHcuF0/nMFHQRAXBzCt1ri7SG0cHIo7fY8cdGTRo4RCcJkykQ+Vm1JIMbmQLdTdgoxM
GBQlZVXeHX9Aw33eRgsshIKVjY2zpFH1h9uQUjufDXhFifZuf5g6dhWOj0RPPVSFnt8w20V03L8I
0QCOBY8Iavq2SmaAnCryispT0BWW1CPtdnbly9g89eLtTsemqJURyu/MPam8xVCUUwmR1Q1ZG348
7744UzbZbtqyvS2LQnW/cWLu7t2Ulj79423z0a+/FdhX1I7HOFXPeYQICve1EkmmsxSM/SrEoBA2
7eg5tTQ/pHl8nD1CNXgTsyvFrII9bqqVK2EheJ2drb88dWMu9jGo6lUp/16sEC+MX9n/fkKwHFlh
LLib8YAQyIRN8lnZlHQgtjX5IDblaOSMZAFeyuSueizmjnxOaxgKVBDirdl+wlbNMBB3lWw2k2nG
HfbzUiFB8QM1MRoqePOejocsJMdpJdb8abXsSVfTs59HxX3KsG67h3M0BR3JRWf9IgIHIpX65jVV
+VMu3pqS9lhgq3pKtQWcnkUzLgm6ExXnDv+zrY7Hrxzw8DRKzZyKzFQAmpGX2ZbhdEjnDZgpJGBE
NlGyw3BkG5lbI9BGJIyR0Rns6JzcBp4ZERgwTp0u1+5XlZbLS4qG1JywR3ihgITAoo1iWOLooc+5
5sdDbrM9wzxJY6H3XMTpnDO1pj25g+mwaRgU3GwLxB3iE/YLTb+NUU3wSN0lHiFpO28+b47GMjfR
wYwFZNXOmQTTSrXyhamxhA1Kf7L4W3kLEN+UW5YIDcLJLGTElPYExBI6yC6FA/yodHDDhqPfS4en
Zr+ygeqk0FkpUu2TW/0hMi6IyJjQUP8RmxJXYYtj18ky6QlezPtZQceAnmxSlMjkbgWfBRz7g2KO
YvczHI6elM/U89i/KUXma6TCmHSY8tsuPkitjodW6P8JiX4wKm1VOaUQjYROix+9O7Bg/tRuyg9E
WsLTxG0ey2XgJkJK53WAZ093BgHrOhN2fUn19ZCZtswC+xrRD/fdl0jvsC63ZVEvEZJkH0bzxQBu
wlYy0saQ6i4qx1m5PWfnT8XhFm1onQCauprazN0ZjkPBYE2Cimp2wnv4z5xUeYEmq4B+IxIRQMgt
j4DnOCC9KzJR0LcvZ8mfD1LcqV+UYFcG9BLBNrBEVzz1MIy6fsV3vUwjAajaJQyW5b6M8m/iQSWV
Gr3GT1euVlsd4e3bhtVF2kjI6k8UzaqxBvc2Hj8LqcQ4GfOlCOHjGw4/x7hC92ayVdSzQIBpThLH
pYXRIFE5uioY792RgNjFxjn0IK5Exs7yQBvFi4vWK7ELODPjm/SH0gCVevU8WF7bkeT/oPBPHgA0
lFH5Gq24QyB3zEsbiMG1M5iouxE8M0yJOPT1x5StuccleHK+BpuWE2ksaalXktxpa2fTOiZIoJh3
5o8wnghcChDA0mn2u+iXSjvAc7xpCBPXwulyc96169rf0JBQauuNKrwbRdCn2mxRkHsk/N73ib0G
eppGLwR1K6LnZLeu0zFzMoZBZhtdawHwU+DaKRCtEIGVoVl6I/ZQPQ00qGQ/6zqJdYCg0nY5m3rt
EFQm3XEImnSBTSmosyDvidPSa750qFYj8acwDKi58LzzhmteufsKbql/ECO1XIGmyAulgomO/WX4
tsBRnlxB41IZ42hYMmae4oCpQr1XzRiPV89DglRpIdvUbyNm+2BCEzoUDx/wyjlyjpKMhXABazYJ
a7XkvB4ehtSRvTlPpHIFDu+EYky6KHFp2cwZTFRpmXKHq3JZGcMCPNJhC+Ip+OZ9vSJbKa6Gg+Ut
hncsHejxLLJTkpO4CzJghie6ybuwNG+UERUKNliFcb2xtohaZCL/+6K8zTti2q7Ufr/NFs3iOxYp
eAvyafRo1NtXXvbYkH6DTLy1NMWiIzqUjhScl1TiqBVuv7t+pG5pUZz9hF6P7yfrJyeDMcSB7lzZ
RuM3Ivle5GvW66r8K0p/9obAKyvqiLg91HwPgjJkfBM4iuvHfjjyBw9EIdy1LVvHJcvFVwqC3vY5
052V9u2SNZxmWYFwVyIKpElTsqOVZE0tcb8e4NVYig+bzMLEG79pexsSJzb9h0nFvJ8biGzVRAH4
lPu/B2Jgl+ohdOClUamf9mLTBieNNjBaGDyc9tkX+LFekMOP2BdK/R0tHCrf3WWbKW+QFxRdNA/w
+hjFmFPMX7Kg2bkyrShHudEiR95YEUHcIjvI0iRGWOOl9UMuDpcyKwz5Kd7qLd4y7yhrpF8cEL5d
1u/l1kmzmAw9OYtnFtgwBnwGeWcM0sP8Aj733i4aMUMqftaXV4vC/T0DgR9pcHUhKNFbUPr+xkNP
Tbkj0M1N1pWUXaBGXh8OY/MQ8dzNgXEHYLfsximcJut4x4W+4AyjJopA92/vKcur78yVmo0Wf5C1
jzVwQItj0R4PpIGbpk9X+0SvnGsflpylf9nyQM/Boh5AUfFWZMWju4NZ/yzWj1JdziFpUII5ndga
iQu680t/BtW9y2MS8Q8L2fuekr2pCnNn2XffbhfJjCQgAEvRg7LGOGkMWNutPjVE6ey3Ou9o3Qi8
5TO7P84ZEuhU0oiM0APJmzuiyakHN1MNFvI9gtegBN7M7Olt0dMBwEbgsGMpV4mdva5JuT8HoGSw
QoeONsLaIbr8sLVCEAwPM+Nfw531H+wqkQtvO6Ny4QUtNDPzbbeCjaTM1oSdTa6ikIj0gxxkLJ3C
DIIWQ6DuJejtbOp391B2zhmFzV7le5YWWNZmt4fYAneXLSJT7I/TTJR2G7M4KAZFRIPXNb+dBkqR
hHEngpVnzEP2TEab7xa96ZmUuPUrojPPQdxY5mi4dGN4a0B29rZJdEYX3iYBNphlSgZRPiGjSa97
DhIRyqcPhDC8RZBEWpS4hkMrBsmuRubcJJufPhwZxDewSFPfrcsy6KHpojHF3Cb6jyJpGPJlvtt9
XGAO8VgIumn4de4zo+eJlayGGcm9mlfa4UoCVjaAocxp++kBfLYGkHWDkn/lYakkd43vmGNC+e0p
HfumcCMuv32eG5Brbq9XFBEKJ3GxhMvJFUyB/C37BY0/3/elJbGvFaveikjWNT9mwVMk0pRs8CM9
lFDobhq9e+GkIgWjD9r+TOHRE8H6hFyImI4JN21L3WqSaNV8jUgBd9YxoWLPMmBYUh7QQAJzE0K/
/2Up9JzFG01Z/s48PF7C7SPGHjTQ2OnSkt1sE8fL+5rxHuk01wsLMlqrN1uMCH0qleIfBxOHBHj5
NCqhyoJXBBZJf+4jMKTZBpk3JN4HJrXVZ/0dmkVuhMRuFg6IfSyKuGBe7Dp8MGxvYubvxFcHKV6U
mV0/kN4w25U2cHVUgLDK9QUungAf2pUfY4+6MFrLtgEJkwBv1UMkWq6hewVJX1Ei2i1wLu4I06Fh
/Pe3hVDb7Q4E6Gmu7gBD1K3rYWflaI/WRi+Kjpj/bK6wFLosFxEDGQmFjDXXweBXjmCCaEAihClN
I/sGXis2tbCkDbp/4dXPUMaIvVev8z1PW7AyCmlcyam74RWtoQSFGyboEXd0o2LPBxPNGLOGKv90
+iPaZ9BomAkt/muYyMM8R9/OMvLi+AiS71m/iICTFE6UxcUjxT8HXa009Dbtad/XE9NUoZjglTRc
V+kRVZS5HM1d0DRkVg4ENirkUQ7E8u5tWzvetxgJdlmJ8Y/Ws1luVc0E712xYsD0KuTX5CFx9ur1
B/5ew1xV2ls67CXMdP2sPGkKPOPRU1i89BkgDkLcrvH6c6j5WCRtBHH2X0xKtfObotcVsxWG/vZm
3CUtU/Io+Crz9iizCoDpHRhFfeX/0Q0ymhnKG3F12NwXTnzW7t0cZdGqAeiKcIjcWOhGShk9bS4v
v+hl8Mww+Bo7hm8kR3XvasZULP5ZTCtzwYxUYjkGOnrkjROo5Fg7dlk9cGjFO1YqPplBgCIjIBXM
XerGEOoB8ztDsL0z/ZveaG6l2ywLIg7qvn8EI/WIxaA0o2y9vZvAfpT4ri8WwZrXh5YrK9BR+AeJ
XxVVcZh/rcHKuw4QCKbJiUTu3kUeDGyUaQDsJB+CFR1LkQuAKlN122zfO4TaS2HPOGXMfGi3AOBn
mc9YHBsm5yAHbyLFmTotaZN6uq1xTI5yuG8EpEJy5byMBew0Tk24IDyxuMNAf4gSLoZaV+ZjE9Po
Vt0shJE0Jnfh7UNp51bJgw9Oeahj4rmo+PEmqGNYFoaLho0omKWtFDGU6KEiXOSpOIyXVIsGohA4
leDik8Y2Y4M3DFzKuUrEtXbe7ICwcnpKY0sBFMH3Qt3uBidfgttAOeyPqziFfTOwcDkGwvKP8Bb+
yIigRam+DgSgYD3BP7th7quMQwHUKwjkgDwAvxQTrSg3yKZlmubvsnuKtIM0Am2Z6Otr4+qUzlpp
MNqGu0kn5PqHlZLgHyYPjebgicwWDa0O63SGTkOMndoS9u6A+vss8aXwAs6WsIpUdfMrKIU+2GkB
c5uWrY0TvNftdbFQ4J50+upQ2+HUhlWXdNft1UDkFXYbQCSV0C43x8mlayJiWqeOahMJ64fojCcu
L9bpbmdVmqe/fhL1XScwGWgHrTE8dto0G2Dv5Wn68EZCkPn6dyY+8uDFnP0GJbAtc+W6Ye7XPvKM
X9ObA5Y1l6r2Qz+mNFkaPZ4gYXWbW52vPJeYt93Xvg/fgtK/unoEBwJ+PvVZG/DK8wy1gpxEhUrs
eoPnMfYfjLngdo64JVlQr73p3b146dbveegD3zViMX1p3m5avEeP33wpPelzJyb5UClvA+6CKWPu
jTUCkveGdQxXvZD4pDO/tc5gji5MwDpG9kGYQgyjuO9pwhKJ/UUqGSTB2yAtNHlaReWbLakHm3Zy
2Kv26Pua15mUiMtu/bhSM+4pdA05r8EZzLG38ZsywMCn2l86xiakUhZmOLuzyXWHxxY2knhByL8P
dHefHsrKxl/54p77rDPxu4T/WVXZZedqlTKeS/aV9WGywVGhEO5etnv5rZN5/iEThCuxvMC9sPZK
N4SulCCK+oeHC0oW0CwM8B/Z0Obm/tuyCE3NgQatd8qyNBDES7UMIMuSo7ebKvQObVtYh6KRN4NM
S4+ln2tqO1+uPdWg5DzLaf7qoFHEuuHSG+YYopkusTNXbS/x46CdpLlK4ROTkhuisLfOQTwzrqpC
Jaqich4PoLSaw3LoAxGKEk8516T7KjX5pWA70iCzGJEyHpjq4T8a14GOc9dnjmI0AuNP46JR3CJm
FUyr2nSI4NkAdZ/19xwS0lCF2e68+rOiPd4g5DjfmMoNDb2WR4dO2g4c/fuXuqvlWBi0sqg/b04/
VtFdOz8O//NbUVV2yXgr+xFsTfttbAV7SibML6zKkbgTT/oq4/maO4yzIRrhWenPfhAhRMufZ0q+
sBh0PxDZ5Vh9gpAjHryEfQ4BPm2yX/3D3ifm20itw+j3JH/5augbfof/aPzFXoRrqff/yTcwBX/Y
eW5nxQ0mt8NnZteY9QG6nSPlQ8fS+TwRFsL5vXBCkFLdE4e2CQYIWnGD5Hx1OuMFUeNRTiM53rGm
L/fP6UFIV9TNbHAQZboXj8SvTjFSEKqYsfDvIOt/VRSLiWuVd9TE9ryWrdDDe++17NUyITKCxBul
VJgflsfW7dFI04751/4lJdNQjb8NRlx+PDBv04mTSCOWkiXQFJjm/mi3GpviT2xp86GTobI98Onr
7IoElQ0J1NQng9kVxzlFzVh4SIIxgALKlob7N4ZlIhSxPSQ/tpUE5IKChJhr4Ax0TlSweVLDTNd2
NgI8VBLkTuK3ba/nVHQoqcz9qnt9r4Bb5+gE0jn7y18Il/dhiP+wkkSkwpci/T4ceOzx2J1TwdaY
2XrjyrUqoCOGxlHao2CBDhDVFXRAe73n/8BpFA3Aa0JClTMdYqJ/l8nSLNT/pzYIGhCmH9eEkYM2
j2wEMIVuzkteO5jJLBzB66hobiSkpWAQSLKu8fcnIXjy4OJK3PNIYe1ENA5cY4eGYh9U1sjrUTAd
e0zGVw1gXdX3oNUCJ7Is8nN0nQnHIXNYvlLPEbQVhC9PBeX4c2wV0OopJtK2XGZi+LHRSTXuMQEV
DmepvfM1b7jtAz2gPaY4X6zYbbLMi+7h1hNTvilnOm4X1LpAQMBW2nwB9m8azeYeHgwZP67oia6r
Ay1zz8Q53YsLNC3cUomE2fTM4bXIkd2gNCfg0a44e1RAdMoXzIk+28P0w3ZyeVNf3wJ2iqmuIBJk
NT77wDySXQKyjU2Vt+vfAABpBCAE7iCz8ap6n3APTqIV6pCVnU655nr0JJa1pyaqG66JuUjsvEAx
wkbHCxLgaep4OtR5pdNYnkO3QgdCV3u3te2OKOy21qBE8N/EZFxm2E3gNJwPvh7njnrri7mbNTP6
XRfwJOlIXZk2SwqxJlkNVPo9Vp4D6GSmQbaSzZ5NIlg/Vp1MAV9Nx75391zJNlmkwjdblf+adXk9
TnpLCbPh6mcTVp9YjUQSxf4GZkLHa1j+kqnVfvaPw/wkp+ZJ8o2y9QQ6DXt/QwU3stOLG/8jKJyt
WcQv+gnR8FsaaOyh5ruLo6vAG8rUOzq848G7ohqea9BjYOYpBHD+lfeUgys3uTmMhUrcUUjIR65w
+IXjIMe4Yq4imnnhKfI+9f/Rmr2vZYvA5EqlZkT2yqGv7zJXkWu1lrrAUrZcIWTifAP56fyAcdnz
LA2Pmpf0WmjVQPfb10foz/NHKH9Ml11/JQn9Au8rFYyJUgoMkzckslIdEHYt63gWYOB/WYFLgQHx
IrQ/ZZIiucICcPynjVVXRyCisx8+7uR6CBq6Bfb0uVBVwkJVTcr/NqrKpVeIeHljwtX5ypYtWz6Z
8SLdlae8hX2imlIqUC6qQFVavbrxBGzqQCjJvtn8Vs6XPDSLJEL+jqf+KD0yZ9UyiPKPzoHoZzXj
LfOQWXc9q87A4ZZhw20ua0V2USrY9y+E7Gpe/rbf04I5oZXiX6/RmYl3C1/l/tl6IzUzQfhzDUdZ
SMvj22h7BCdz3oo5bJeRyj/jrqTGQdRnepDmUdRapDKKsb2JsU3I/DL4pRrNu9HKKqndoYE1enBQ
4uZ97PuU7GdzPTwJXnCARiYui0iv5Tes2UAKoYq+E3ktG7MJkqRS4m2ZJSr9j09Dd7rguQWmulrs
rZMGDk5b1RASiY6WwDj/ApO0gKfNG/JrLNGd4r8xbzllunVtM9B4qFzM5ifN6Ln9+PutkxxYNmJH
DOQKokj4qvjYRgU4ASzUCSsdriKPhlQJQ7GmNBe4KGysPXZ20uU/DJoCO+hGqb45Qq8SHtzLCZoU
32/VyYe19gahkRMDZQ7phMtFamkytVZtcdkKChvUKhUqFBdt3Dr3bEm6UYMDUMpYO9KQas+KUctm
lXEPZPhO4wNszRfLzRXRPCQIsmFYuhkd6EeLSXyntAkLL7gH2BrEyVyzEhE2eixAD9vz1DE5LZI9
mbod7rFWvmAo3uP1FLoj4Kd/uK/X09e5DAanMdQiocog9yWaeiYrvqYfYj9M8keWUttl4bFadz6k
zFFLLxeOKqJGLHLxi+asG0JPmuaRr0/iHoTZiI5OIK7N+gCKvtxGsCWkflUrA75FhGv4KluPg8qd
IiKGJ3qlisHRGU88r/f0nTrH//pjjBeptJoXLpMMi+VEseK6jHJz5RDg5WpM0OFD0pYWmaM+PLvy
VbcTfy0pWLTxulo2H4QvZCqxaXkTSQtVy2vCchqMIlZZE1OXUzlV+GFXn0eOPoYJU+8Tr4Tpur50
99+WT8koLN3fVk901rK2hZd0nr5tMsWd/TI3V6Gzle1pwQJVLJsxQ+dkIt+pRsfd8sKCaJ4xuRzC
aBAhM5TbXr9u6vnw+aMPdNDEcaUPh9wj4BjXEXJ1fDGmWS9xv61EBnO0r205+BbR84DLA9ADlayj
Os3/C+kd2fZVCJbscncURUz9fGBMdUHmFs9BkJIzDL4Y1ubbCnaipESK06ozTEHr/GzZlEFMamo4
3F6w+bzP1zrop+wERFz5umd9ncISQ6t7kbQ9b0nnhI5eRUMNKnZhHjqwDltWitHba4QK+yS5D9rs
SD8yxIeEHhAhsf5s0OD9Tu4pC8/SeNtoG4HBkoyE7Bp0LwFBe7Kc4CW9Sa4AL0dn1YETzYZlppaG
yBQsQo5bwrRgFmHx7RmDnHGnGmVw0lDvUn3ZA3emPlNqp7Nt86AZ/nsOiiK61OAhH1n4Kvfa3pKZ
pgv6GMLlegAJRdJKPgX4ptzRi9x+D5odZ+4QW3EGWTWASvn5gIQfV4CHZgmJAjrCdM9Zyp/tAUSJ
z96nsJSTFtdUr5K9EDwhF0/XlVNRFtFDJyBNPpq+Okzyd7gtB7v66RDnxQVcDVPBwEtDmF9crTWO
T2VunD2JUrsUV41tABJ41KDzP8E6KStPOfB/HAxm9mNPMJgLRlX7EtEeS648o+Tyqcy8fc0DmPOn
rKxi2jpCQ8yG222fRCxsC3U82TwW5Uo7Jpb/aGU5FbNoAm+0I0FVL4fOYsoumBa2sSKDXS7vEpmE
oprhLqGa2eRLc0K6Za8l7RuK8hnKmjZfQ9+7/soPvQ5diTA/WY8ndRXgLr948I9RVYg31SM4aU7r
kbcXr9DfpNPiv5m83PumlR1U5rRVyjjhWU8q+qOkqPFuUZ97V1k30pHZI0Sor4H66btalVhUt3Bh
D9KTTrl3G2PezkyRipP1tBiQdo8dAFy34WCft0Fzkju+1AaFJJmtBzFex1XnRDawb+o4hzM6fPuz
ZIRD3THQI13pCdMqozXHHO6ABQjbJKwbre9lrmTNBaDLjAjFzvWYCuqvqodBOFlByr9ukW8Mvci9
ppJGdDieP7slb3TtFedohLzCem48HegFIg2eZizT2tAOC50htjitFhZ1e9PzKFFRZC3ytRGguwrg
PE9rZmt0IlfPPAHV1ocbmviQCSfmz6Ptdfpgy9ZixdpmpPX6oTuEdEeNj13HH5yR50fp1Pz8yLKr
a2tUh1UZ9INPecDe2BXYESj8ORcIa7VLys06aoQ7JYm83Hsb+k7CCup0ntZZVOZ+46AoyPS7om3x
VCJQqef3lll6wFlD4d6JwdzNbTBupLukBhpzImnJntE0Q7/ZryKZ4MHsCVy0ED1JGFSMCTn9TMYD
yThclRxvFw356ofQFCkez9ZmEPxFr2GfNm1rR2uVVIqDOksjpb6w8v40FvE/LUqnwdlqBCrmVdDw
wysj1kGvuyjD+nME4WPbdo9dHdw3qAmjLW3Zo1p/bmnDqdVLlUVc7CTx5qQLXTrtIuySERGAVNz8
rJuq0oTSPMDFMP8PCWN1lmF6ZO7MV9RrHkYy7FDpohqVom7eJYafJoKg9AOhJnpkgldxpPxftd7z
KVJ2nMi9qIZxW5ZGcbUBz5rZKyYJiND3INVvnBv4ilYy9eMQsTUan4QeuK11oAhcI0xRrFUwHufp
vO7k62Xz176gH8ObpbAOeXk5vTVWXr1BSQq4SLjabSmQURTEXunsQpsLhMUm7C9yw7ateAuw9nns
zeLYpL3upOjqHiaYPcyaZ8bm4GYUJfTVU7We7I0sQVKOkV+uZfvoYOktDXey75rt0hWvCjzCwJe2
v4hA6ajHfxmEneNgGFN9obu79wxBFvv1C3FF3avSu5O/WS+/fS1b4SCz8ppuGyj7qg/zNNddOpAy
ejT7BexNPrU6Z8TZYiY1diLBSQjyxTKpn7NE1nmNIvS9HgKC/9BtDMUSc0TIIfrbXiMmqjms3AQ6
Pg9Mz8nckJmLdLbIQ+c6C/FScC/PDNZlSrsiqv3D3eoYLK1YEzbjuj4SKS9+7zN0TmuzPv8ebMUG
AkpdX8kndsG7AaS1BgEnGNDGQJKjPht8PnxOxtLXPgijYVJshjwTPGH0UnpS5cfwL0AyAHX5fdaR
o4w46T/9PcuOEea1Ri4mCDJwZI6XMJpJoKi04obsd4X3r94m82e0DgtxrqHUzbyTXTomp67HuxZK
9WB+X/smQRSCIUqhQhCXJyYluJBTBZUjwwS37feBTWfELv2qIYyfJExiJrl7ftiq8KGAixJC3qgF
1NKjWgdiLV3lwNCnyPqVmFxTJ+Ap9qhB1V+xVjihUEeKWHvjfagy0OuL+bXKrbTrUO716+pwkC3m
NjUrXCw8t9kDoTmhHA0uQ3E3SdksCUZhj05m/YVWwzVEeH8HijPrPSgapQFXNDN82lz47DLk41qp
Mgn9GRh5308smjfR0Sf/LCRZw7XimW87tyMHsqUePzJgs4i/nzKhdyUgLFP+PA0wGlg3e6homafm
JlDw3W3nb4GQ9FYfIENAC/Ek+KzFtCZ6N3F110C+L9Z7wVPLtO/KL3kZYCWZ3vyfCONp+tJsRdqj
W7O4Pl8Wa+CR4Gtau/8/FgHaZVKXDX3N8hXCfQF5WROV/t5uz8Fz2c3pZoAjI5Q+1uEEwf1etDPJ
//bG/eKDKae7Hw8o8gCzqcceasfU0BG2zXe5zi9gCrs4qrOq6bq7a4UghkpHBwU4cGGjD62qTwBn
I+acs4E9hytEvnKQ4X4uoLmWJHYwrc9Pj7KYGmXR/J7qe2kuODBwWOqLqjXsqmbBWEUYsDb+LDPG
aZ74jCtKwibYE03+Y18NMvPlFA6bB6dbdROQi6Ev3BA54FU5Ke6aWnpveXVzjArVgfbhH+2mdsNn
l3ljxFHaw+YchriV990ZfPuNdrx0nPSM2Lzmv5NuoD5sQ4rEqwY5sEildvSwKqI43q5KeJkFPUPm
n68S86sAInCZD1ApMOjiNOQQq7zoxZAkgSu9Q7YYTqtnPzyx4OcebHkRPkQKJ4llOsGxzBqz4Uaz
7Xekt9qekT60iV5ulDyChRXg1hHpxbJFL8bL9TfGJ54SYrqp2o3PXPQs+cPhMS/QkiwR9w3S3E7X
AVdS4bwDt2/KRlY3f6MyjWMEqI1T3r++fiFRhSMOtFjA38uGGUJsBtL7G+G6j4Lc3K7V4w+UIymk
tw5cejR9f/4O7iwsPUUKvoomnhB5A7cDLvOkxuqpbAAvh+e7ztPll9zm2X99VgelsS0wtmJ2F/9U
hApuNu+FXFyQxfdbEvLWiLNBEHCh7A4FIXFV5JRJmSHk+tRde4WJdn5OypP5KsABtAlQxDZvOABL
PV0bkXrWyGBRHNwsLeam1mo3xOEoBgJp3pFifBMoxCE5XnzVxbPMCl3VRd6Cli/Fk5LrYdiKEs5T
nVndRvW7mvRxSNPkwMd5Y+fzajV1R5fcGLeZZA80RnQ9FA2iOnE4iNdAe7Va6WXNX+TYiuP+o/0/
qVmXaHSVdWbl6Xwar4Kpcc+0h0jExl3DSq372Kco8EmeUGfycyXb8YY67RsyNsc6rKw/e+amiQ+1
groLt4SWMk+3IDZ9EK06SxDk1F51hMV+OJl2kIDcuZsphj5Yz9lhxJrRvhzBFEYF+k0nllangTqI
A4QfWWNcLlherAZHtGUdY64TIQt5OQZIV1ViDIaMu1NNg2z9GP3y+L9ywE2MDECHoR5TZNf9/CHE
/CweeFPMVGI4nPNXa/HazAMqBjGx6SMPjx+3Lda8ZPXYhPWjI/wnplQTsLqPXhLJ2FW1OQ/8HweU
nXVsJWx1eYRdR4WQ47ioM3lx3sDkUy98HqnqdeKRSSrHohO5H2EgjzjkONWrH5A2xbgCflnrBh1+
xTLmAKjRZtTXdWR0SrSLxWBhc6kLVRP1rEouw5vOYTC1lVhKttxAdtv5iu+lfcUdq0wGE03uKqCj
9YbxsUjBynpmwKX3HjzvoE0JC7t+d+6RYo44Ffri5xFCOwDP31cM+lrTtLOv8U2+6XmIQe95Ip+g
h/g+wjg+EDiCGDkdYDvW/eTz8Y7gTlxjXpmjbKXdboyy5MKbI4I5izC7k/F3HBxdG2C+dAdh8vFa
o7/+p8qWR345BZGr7S6Enz4J1KgGweJ9c9vHjKe3hcNhODgdYSgt8dQokz17u3J03dlMZJOc7mcy
lyOUbMlNvovq+42YOnwkR5aXknlDd2rXUrDyp1X8EnfgKc8Iimsn10cQRlU0rA8jmBKrHCAo19r3
FMAozdkC3WYU7sdhOWI8VK1w6k+2O1kMg1GOmYGEc1mIMpwWKrr3v4a4UzdPqy4kIs3BWpB/JsOJ
vXT6WjdBqAFyQrhLNGIZV0o/F4q7uG4CqepLLs800PT2bkrMhTqaG0RZW2PnJHLmmY8YraRahxyF
DRf7jONIupLT14JLOWsPfIbhMpYbd+baOMaAE2kHYfQ5NgoroQdJ2IgSrRPdJONIb7uPbwVkjuZ1
6ZYBpqUAOlmx+4qH1yaoa4A/VK4tu3539hy4PAqcAOtWmimMc5SPxwSQGNzggpydArB85O5pejYi
oDM+vXkETjDEksUKv6ZbwLIvvTENkiIAyjgTnB8zepIqr1gXZW/JKMzX08kaLhPrjJKTpk1oNDSy
DNlsGCNg+YLnYFfWEJR41niMwQXTbPOFXPdMwLLwfiiA9ZJU19vz/iipH5iUhX2LUH4ao3MNa1tj
Je6uH0vjfety9TQjumOAt28ZTje1JeeYQTVvUOfCHiNZRSacaIQkjp03PF50MjtYAh9hE8OtDqiH
aaj/DLV4OkrIg9i9IW9i5JFHZ6qBZjh+r1D4u2GSmlhm9fYhhXQgdk8BtRypgkJXGJRwClGyXsaP
+t4w5iDE3hso+uvh7pBfsEBEwxzYLxhDkDTUm66Bi5w/MicGjeWqTPVTLwijtMOC9eIjZAm+UfIz
DuNRUsTLmpdf8FdIr0GPX9jmbilTwc4QCW1uySayvyVhKLEjNPasIH2eWlU9JvaYxJc/X4DlYT0D
A8DLT3KGc8PswoBb0SC4Rnyzd8I0dMB9X/khhACidV4uqlmqrTHcHPFggg9gU38XsMnXfvuEKMdC
kKerdJ4lgaB1+/pgo5zmkskw73X3nmZnIvTyZGJGGjvQ68jcSy1bdg0iN5b0fQiCZOLQJLxtq1fJ
Dw40i0YYB8DftYZk6ECieXOyM9yGiexjPHgnfN39axh0zTRxD0jWLcrvnBKSTIg9r1s4jHKi/QYl
oC+L8E2+3nColjBZwIRuHFBeM2iDAH0Ndb8wryqD13HuAED5aaLpiRtx58J0v+0hIPF0WA8RDWiH
Z9BFzvnIeDH3Dw0bTfcz+EGNobyuJwU5ydjM5m3povwGqmiii0ePSnVDLnLFCiHZ/tIEkreMZ1Bi
b8DEB1xDJNMIAuFGGLKE0o6y8rTw6ZWjqlKieae3mdTj+TLOgd6OEs+ERETs1HZ8QMHI2NUArm4H
K60bOB03JvS0TYPx62Y2p/1jg0ErPaAg9FekUaC7rraV3eI+yIs7yhYIKOumOI7ML1bjh4Dfwf74
DVMPtvBKlzXnzdkoMKB3uZWYtP5uw00VNZ/rikSbjQQJUZLHUJZOtvTTnaAjkf3ATDyL4UAClYOu
OXqNAyAI0/5PGzz3TQ9QgTk/0Sihor/vvtXs1OlH+bxd6XVAZzHONesYdpKjrya602JS7pnHWPX6
jHJysdPK8RFw7hNhJoQXvsS3lSZ1q0NKNvdY+vrJ7qZPM0LwP0yNs9ChGJ3OhsNY4nTnmM/euwyT
jFsAelabB4v+BOkMBNvyZOcjs570Qy7QHej3FhtQxvs62HaOvDFSJf24PGiJoZXBqHUIVOI/CDWP
FaRgaAlZ+/xhBG8fYdibUJKEplrVmNxTLn2AhT57TbHV/JWK4zSZf1yaSqcaKMM5PvagCuIPMdfX
4wF8YXsSGIVMfpvbLLxNk2hGijiZlBRaUMuYKWZWc5BgpS8qtMBNO/V17wtiyIPuoSNsb35RDus1
dkBgO0soSQFdo8PbcMBViHN3R9MD89L/VgLAH/tBACgdweeXHk8TVaLAguNBvEjFLH9E/bllslx/
R3SDeRIu58teUFnv8UfHzhjAz5BT2hUkm2jfEEduaciKoCVFv+2ja5HxEF2gSrSHfhY/nXIbpB6F
FamCRLQfQKwTBp5V0ZVbi97WNg0wqkxH0Mbd5ZLmmnSFKf8dovJzN+lkI6jmP1YsWWa1iUaNxeiO
lXevZG3xLWLIpa1hRR/cugsJt9lSHzO/PyAB4ILaMANwN2Jhy1etCaBiD1X7IkaX3Q0teUGo/TzZ
xN2JaSHrUiCzNHle/ySVeJJY6itkXvsoogWauFYGtJMQuv3zXizVynomxhNiDZctecQpUn0HHsTd
DK56Hx6J4D9VKcHigIvxKgBXxfnCQqLmtJJ81ZmxmIvLBOtNJ/ivDRspeE5I08SrZtTByxbRV26q
lUhcluS+qqB1VScCntOkLBS/p5VochLcXbXaP3G5Q2uVs2vZY41mhj+kLRobCLHVQYkSOWx0MnV4
SvW9qs5W9LAY6VwIg5Ncpz03ZMLH+4bFZgD3NxFxJStjP383UpgxaXAuLofB2gXHrY0ZRlDkrUSH
8rQ2VJVS2zplxUHnHvw0G0acMgttOpFEgC2xnaTGCZnmiXhsRTCYRY56eI4jeP5gYD2l9XcPK5N/
pxW+M9uM7tQ0I3matEKG+n8C2bpkDWrwdyPjj0Tp2LVH4ynECjF+vMWvZEWUmgWrg6Frc4rNnG2E
qKMfJBwB5Bx2ATiVY1AJUztkMKXv0tnwhO5mHyVpUPNgtjuFTMcZG5WBOls2WEMH5Xq6/lWdglvV
2tpaYhYgs4nAUc49ApNTjq5OfCAMgSvoUSDJzgKZW54EHabbqIA+KRZGmPN+oSTQe4PlmWF56/nF
i1vOVfOSKjQF1SFO+D29z5yVksHpc1LvafrZ2KRR4A+jhSgASUzeIgH7TO1iSBMZf2rquFuViaug
ZW+CzMoUx4K8d+hLoIbQ6XbUM9E0X6tpjH5zXSAzQXgyCGJBA7tTLmiAM1A8Ym1CNX4yUQAi+l0Q
L9zV0mqMtXt5jBS07/7bksFWWVYvOABiz7b0HB0+ubwz3tDJXPx4T97G1L12iSn9Mc3rhaVnklB/
vXPTKqXvLO+7WFcaxX7WWdM2TVjKgPj2IvpMvVYryfitKok8WOJvWN+J0kefQn6W6wMOtxUsGc9P
qcyHtEUusbSq1gbTj7fbKGaMhKwqPJ05CiN055Lnqm+j003fJJML5Q9IDKN1xxfsbkpaEU3BxbQZ
i8f+hCrSHaYPD04bGz4nP5kVmueZKtxWHpIYLduZbrsD65bMUNagu5PmcICWZ15Y1OS70rVWX4iZ
/4hdkwrLi0dS1Jp7l9/IWOqdZ0vzTad6D7jMufVmxXWOocovsUPXESICKQ+GOMXwxYEVfAV54B3p
ulVu+vL/Fn2z4x0p655egrmcgw2FRG17LWwusbWBUrRyZ9r4JfLREc5xubWsgT+my7Hazl/CGZTe
wEf7PhUlw2X73kxvTuo4bQk88oLWY1w7oofVThx6qPNVgwZ1HkeeFoGeIF2a/ei+llvNumrayG0Z
84Vpx6THjjv4ePPGKjtF1m2Xu+ebWj7JXhjEAEgUsc/jxaSgLrSXyGOxyoytCsccxdcJFoUeYxla
pJjNrgX3IYwZeUU6LiCGdHuHbG3LR4U7P+L+rLZfEsfwQqiDhieG6Vu/ZLZk8lgbnU0UzagUVPVS
GMR/Orb+mCJ2Gg1e6SdGlQWW//c+mqtEiTCNOH35jdyeZ/CsT62/Vi9+swgindeDOXg7cwR3sZNs
eb1hDl98H1kK4f3ULRPNMEqIsO69UDi0JcRc+vrKVuy5xFoVe/pqbStrE7GPx1h+e5/ed4iV1S56
A4DhHWI/5Td7vqd0kmUiqOY26h4KOD5nWNOPUD3heYGmKg0tBBk+LeUuoK/qylWdc2+lEFMpXvIK
aT3ZlLsAkP4r9G1bv+Y/VZC6uXeFAPMAgrCCOSgl8K5teU3Ns0b6PsSqRzmDraSDaLQLrEXyK0kf
f2F0+/JlXoFclNdxzl2Je7sLq1/oEdKwoEQhgWqlwS37IgzMS0pHk38UYNzv9pI9XPGYqWwwtktN
5FkzVpNf9yK2B9/X+0KY8lnEVZ65Q3pnpYnCTWelzz+wm1WBMtZDeSkE33QHCAEdlsdwsYLS+8lg
3ourpSLLldXR4Eo9WuUxjpnWdJ/q6J8kHcppsOTpmLIQwLreUHxFkNMqFRU0KszGTCq/ULTfjFAl
FiEiIoTRjyPugv8UwFuwu+FxAtMu98PRxVLnetoOAfKCHasPdsghwbhN7nFHIt9eCBbRlt9QHowX
c2qBbBsAVxVhCeAb8OVO10ngnq69xLJcVHXwS3SXMu2Bzvxvs8MpfPP9WqyONHfU2dRRTeTV9Q6h
8wNcH7owo7i5FEqvAEEhzGgNiCtDbEpBuJsAWkbO3F2U+UWKG/QYFMFKFEDkfwV4AjSbQ/66yZPf
af6M7c+ysgGG38WWXwxkCspms+VGlFrWYqMGUSwJdhYRaqY7qzDSp9zQuCXp9E78nb4E+M8WIvoD
AqavUP2omfazTPEMOAHo2xZM9vU3foVnK8a9aGFDFXaVEVWko1sO1omHrDi16K7YmkVVIWIszRux
BToyNmYN13zvYq8K8eQmvhNBZs7dU05EJTatHLvTig259J68mus13htqwiYxWi2Yuq/cTerknJ99
+BBc+WGvR75ETNkLnGelDtnGljvmibIFALKxUBGfBD2kV0w615ROiXVi3Gs/zNcOKWeHgQoHT8eE
sRi10cKvpT+xg5nDcih5+kVjFCKwG805th7rHqyqf/98GXFcfXLv75mGZG/bOzd1UyACXVCMtFfz
i6qQ66aF8nlj9KHS1XGuvh2BUu/kV6YJ2tDkJJet/Qk23Ng3dWd1Wm+MwS2Qbq/TW8a2LWDAdqLQ
y+t347tesbW97vPNcEC8qxUS/DCWJNAdOXOAgFobV4ka2KZBr8Sok2/ekRKJChUcZmOkP7leo5+c
s6+EZsD2WybwMz1zqaO568NYNTn4096KLtibLD0FACJh+pXYyc19BSNAKfdvTnbQp7V8LenjEzIv
yG/prDc6UqXdZ9/V8xFySIEln8wA1SJCtF8eeAH9RGFWXCcuPA+xML0/2/BI5pPSshWUfxbS7imX
Xw3i0q9LK5g3aqC5FA5Y2Ktj2x7yz3//PN4YJ0kNu7sjpDLHso//kx42r8/64sVQ76z+88SIGLYR
2bjdo+02/FpBAUHqKBmq9PG60XomtcZP6i+Ms3iSBFDug5eem0gGY7X7Sb9eKd2prj8wLoWKvVil
slwppc0fLO+yUS7Egm3tELmXP5q5kX8CW3F2QGbdSoHz5hsz0XQyZ74GotC7ovN9v6BLItkQRbao
6AGHP/+t1yc5lzXIYCAMcPwk1UDX5gc2hcfOritRAyq/HdMo3gJmaAWumLZt4+Fo8M9e0t2i2UTf
yPvXha7r3dB8ijZCVePi/cCo2rH1KDudtlIgjD+vCsG48Uw/P5LbktBzv1YQy0e8j8ai+IAx8BwE
dW/VyeObJHS68MUb3fWEBOYTc8CgQd64664XMipyq9d4J7k5P2WkCSzZ0dwLEi++h42pUNXyRBAE
MEZ6FP84mGBNPIIJAIf3EULhd4Lnk2JdbFPFPbCTLBvmbrKnGW8vslGhmRctXcE3E7xVwpq+3B4C
TP4hciuOP88U1dJRYE9wAs8yQptyRcor/dxzBkR6qN4sC8lThPrcZnIuUiDmG/vFFOxqjH8YCRKz
onLfbUXSG/R2NfxztuCw169djCIY4A4Ja8bPHZCskoYSyCAGNT44RvsscCyIUNA2nZuFnpG+RjdM
aP4FWdsuE1UofBObbaqXawf5LEW6J0aOvBzjIMwoyGbdshmeR2mfms+msCQZySZ5Ezgz3925YkJC
ZEoqUYsM1d+krU2+ia2oFj1g0OCJ7NlBjQL96pEO12stZ6DEm/CoGEfP/JiPHZW/V9kUFg1mVTDI
anZHfOULEXZyO7keH07fsIoIfPFbp7s1N8ZA9kmE3ctwSU+AFUJiw8HL30DLnFG3nUEvzYG0Wp8z
Bwro7y2pJsvMcD08zDANY0xQpQ1RinZuVCxSBNgEihsZYMxTi9lyR78QUh3q+ZZTP2OZYYoX0Diy
M3RX0oWqz9bgXyrANVrTwmtoTHSV8NMeV8mq3Q2Ps/gg075A9MgqD21zI71mPG3MRwucn81Q+cKn
yHhYOPCpWL05CK6/3ON8rbm+1SRft3GKctIES5b5hoq4PQaINSA+RosxfA37Afgw2mUPsOY268gC
ShnnNMEsExasHCIvCntJ1X4OXwHvm0UrjXr30HhW5AtqtFkBitjBpTPrzCEV9eOwG7VbKUqH5cO3
WXDU3sziFG93b+2Q2znusYZkKuNmDo1h3BoaZ3u8qVhR/MJXRn1L6hs80/xya0KGWshLWXlzuF1J
a1u1HxhfyWOCvFFTl2/wImmqlv6CBwRFE6Hx0TWyqNltMvCeKohqScZuFJA8mXbvzG/K54hyGhOl
rENJOAP+D9C5F59BfKmVHm4K0/KwqFKx81bdMwL7TaP8h/Eqk3k+vEh1KJRLICqcbE5FZcXFwlPx
myZZHfLS01g8OZxZkmvAkhICQz/Pvr+adcjc1AYi3QzZsqNcogZQyhAtVGznWnlRMp+rKxDtJl+1
Rh7dKRWiX53zPV71uOJckwTQZbMj3kd7LfTjlv6Di41+QeA7/9M8QgJXxlnzEoxXfxGVuKlgMvPu
l5RZsIgcAr1RRETxRVydRJtO3HuANUukM8rlHf2760P/SrJFCQxZkotK0nVMec8rqc9BS7iod03t
LhSq36RCSLPzBe5urpkwctlZ7eI5hTYjnFuhGbJqXu5fAExLU9pKUxq6RR+59xYk93z7fgN8UE2m
Irs/E6UfdJGABN1YL94DmMTgrCSlOwyjHEhHm4B2fGCBJ5Ve5/iFYpD39ynGMJXhXG/BlA7wdnQ6
F9mc25+MGZPkUWOrzFzi4NFTjMyrrIyqUtzuQwA+TUrVWouvuOUe6UxdpCdrowYURndmPE5aVk7J
nZJNMwIsQlidZMF9yh2oHwN2KgEuGLWgx4WTUyjLh3oPrBjqhD21YNE5c/k82cFECntMQgqrQqwg
ozk2Zw8E8QMuBfuQt7Ryq1WU1XJbLa44NeWUdOdMneI7W0edIA290HnLiqc4TNb6aAIpRUMx+LGg
9TOoOUBWWuHazAeiCInWFYXRTTplCiy1OqegNtDH3a7ek15ERGI/auBy6LqIj9YTDB1G6kvIjpL3
jihiRGgrVilJUuBLxzPbTHP8WViIzYoG9xZXVx+8+KEL5029jmtrXQ1/bmDR1jGw878yRSgwmvjF
QujqlVtvNLSIvQ4Kki5YQMeW6flooupwC2aZauapAQXxydODqXt9Ijx9yKh5WxQTUMA7G4TeUeOf
zaTPnRhFHZO5PJyo7r1qfzHrAk3t3ph+14/df+n742ZTJecvtKYRnKveliAsVGORL0qAUHV41SuV
tmXQ2Dg6sAPhtY1EWdmyuPZrZp5/GnGtxzBBGki1Gea1KctT51u0e5bJLdObKwVxm81zT4DDWWyb
EOdpAgOwmDlpZGQa8MIUpyh8m3Zcxk0MOfmFLykBfmUL+xs48CyaJLLCbbK2y0xKHeJh7GwxkSGM
AucuZ9GAOtBHviXcA31EbYmwUd4anbD94hNLz75EbeSt8kQo1X8JGyAYo4YV8vKvnGM+MIfaiyBI
PpnM8D8veKs7m2oGtmhqOXL/DnjKY8yuaH0de0QHNMDir5FZkBTeFPjldR6MpkbfOfM1hiXNF/ob
fEAbG9jHBE0xEa6sS7qRts6bG+f+u8mX0H/1pdqWL7OBW2zJmbtzvteThmmqSqGOJ5p3bw3F+fzO
04W69iFqQLS7vuLNOu1FE+Yyr4bPKGEL/0oKQZajitXubgKZXHPoVqiUqdNs7oZlWrGPzxgo8Q44
BSDOUwhdtEEdyeZqUrYI3zAf5bFjdg5qSI1PJHv7ECBthaqXAw1sTXMrNzwGXpQhy5OelAUkhCa6
OY6Sdols4w4zKMyILlgz4a0vee+vc9a9whz1HHRWw9nr7sF+0NLfZxJkzcUvXtMjAd9FU9rrF6Q2
Jux5Ba+oys1mv4DhP/rXq6T5WYetPLBTu84peme8BJN4Sku5XzbtoKswUBOO+ZjOazgv+dDGtytR
NxvtyPjM6khgH47gUa6Oroe3mY8ZXmPRZfClj1E5pNakdeQS0vyDmm0c050qjO0lDIJAk/XuZl8n
1E0d+MytEQSXZN+HBY8+Zf8E/yMb+fBn50VN75Th/QbahKPBhz4uoGRaE/BUM4isFYrS7qy84AQk
PslTSIPXHsO5sbOnMF+Cgb6RkNKktak/DAEtRpGJk9dSfvCpczT/P2q6yzOXfi6XX1DHrZTTkR4K
NnoQFfTO3LodK5vNBq/ZdgOGIKLdRkVcIHTUCaUzrvL+z6eCCXnFE3YBaOdv28IfWdgL/3n+xR0+
t8AfbMAkjl7BF/T0Mvu7ssZDiEsnuQ6W1SgDhTd2zdqmaPUZiu/2RCmjIGEgKQNzWoLF/aQ2Me7C
B+kibpZUisO/jXTx4DqM2oFuFgudHXV/jgXetEGSGf0UiGbKwx7TGaK0vbqFyribhLa9kZ9Pb89G
DaSUGSNqd2W8bqm+ENbJC2GPEmbhJGXRwH2pC430H547owGrgQjt6M9r1uDjSHzoJv/zyL/e84WG
W8UBDOx/tX/8eOlvPzbUC5jMEqpiabE/MHmsN5htG0LeN3wgIuS26cbrLPuRJ5Sdr2QcFce+m3ub
3FAFPtxEV375uD8i/YvQ6OaWrqvbitrkNj04ZMZRzpzc39cLHlUsGpLiJ5vXpl+S6op8N5/d4RFt
vCN+aJwiMj/NNO0XVxk1EjwU5qevW+buH2Nzf9mt1QWnaAOT2eKBpGTjpFH5vFnEH5rx3rTNfw0w
UlcEcqMFiGBeqEYkFO2/Q8TN5WgdL/gVIL0kSMO7Cvfobzi+V3yMEjThzFBP+T2bmJdKVyohyvvj
LgdPQbro67gzpnFB3ZHADsZPXGnFqJd6k2qZ1U7k8yESByO7BZxA9wOLEJuGKjGVv2iiBykgsz5N
vkorlKdmRKNkApy3AHRpjbMDmsQsPcBRu91ei+Vw1w0XBBpkigZebH8ZRYnAymO5vFnbTCpzTsMv
2gYwmHCLRYi7vNYoHw2YQtLvIrm4lsE924afixtJcZe1EBkAIrfPFZ0jcs4O2njYsMrhyD8Pm/kH
HwfKqUWuaktLYwr4QJIFqYgGk++52bT9mw/kCAtajog+j7PyvcednpUB9PTjDd0VhYviMNnMrGYo
DVv4ZxfVQ0SCSvnv+WmDwuBBx5G4jLxKc756mHW6feON6uDhB5Pvwm4LRnQc1vUkVOcd7n36VCLH
fgypVU2UYuw+0zxQbSjEid4wufY6EJF08HY8k4p/JkUPWT0JEwS73kpEQDD32nOYgjU4Zv71Naxz
wUbQ/inBBC3x/TntkvtkL4r4X10Vx/Tqf+23N6J3slv8b//9cFV5vAsrjFlNohcSySFXihsXlhcc
t9sCfyESbO1Ylq2HK+y7ajojf00rlxjPni979wSt96edo9YW1N9U8wGuSZKa5kvDq61RdrOjdJ65
p1ZajQMXmfAjNKxQU1RNs3A2SRrbnu6niJxjPZGoPx3kGM8vkFaTlfIVJq4OKirmdumOqUg0HLbi
mBAZI4OHbCmp0tV9h16HBjIEk2U44viFAZ4ZKuMIwP/Xfkj5sTEORKOdQC04oKCh5BeC1/3xoZK/
6HxDDr389leVDDUhRBxr7++ZZpoRxArLvjIIbT02DXFiIxHWNyRJRsSUqjJtWiGpUIbDx10D9Zfj
Yjsg5xpirfc4FY+2mpZnpusZzAxcji/pKB3hgFRQEYaJAMzBVJU9XfuUWApJJbO4p3WqImf0Cggm
hO9gO1felvLVuxarrCP9FoKL0oVl6irpx/IzSMWOTf0xs5hMh89ZM+NNqkBmk9mcDrhJKt0fXt+s
Ng16JFFwLnEhsHsDCj+3oakc2nUskg5XP46cHv/aNFAu1+dctURvHY7tnAmbBBTxZ0r7vDGFjWfy
iM8kcjrVQtpZE3kYpDa2ucJV7IMznD7JeandsB9V5X73m6tGqzQZSgWGDE86dBBu3btBZfrgWQVj
APTCabkwR5xWfyl8r2DwRaLEYWVOYtIEuL/sK8GjG4Fwq9NV2INbzlpVeDdP/ytky6W72tMYTlVG
AG3W++AWovncQeYQ2Iex480bvstKtRtHjyvifxF8LxMBU6f3222Zddg2pzh0idWK2fQ75YeIFI+5
GfzzT6woz1j/tI2D0lqNz8axWqy0Liqf3v+CX+dBKojLTXVrWQy9R0qt2qNa5s9075AwGJZUAPjc
48MkM5csquSn5JcBEz4s+NHz9HUW1zhR8pPzUKnO+VAXdV2/1lDIC5pMslkDNGUbZXf8YWqFae/K
6ywfIT8HDEN1pDKcGOK0EDybSiMGOAmRlIdKBUPl4AFdmG++L9aKJyZeKPHZ9/wX9Lf/6O/wLJS8
P4Z7dWCL9BOdioNCafpY9ue3GCqzu/UkTsY91RXyAzlVtFATeAcCMHi5ecQLar4g0AQ3mY1sv1Sb
WdRBP7chZlRVW1GM43dJwOPxBczGo1jU67egnv6yOwxCyTz9mQXD+tH1JPD5vCv8FYBDUIsA9hLK
8KhHiKVjgHCin+E1Gs/vHlHLnA2YrL6MTcUwbBhGV6bmAySgSIw1jZrPGwfsKS+8eTyr4fkyD/Pk
kNwaiLg33IVU7ncx9erCeuvKHxmHiP17oL6ds+Vat+90j1e89LaiHSOcE/ctU6WRpXxWd/wee+QN
tTGaIbYuJjUBsAcCaiDrb8QaZuGKL4bZx1TtmEyA5EhjorczPJNJYGnbq9u+yWlwMv3GU1y+y5Ui
8gcRoAvQXX8QVxkdIyTg/cXdYIyJ9/v9TfawLtBjRe+DIa4au1niU6E2iECFN4N/ae5Y/vTzYFB4
dkuZMqasEl4rMeup/uZyIQEgjt+aUNno7BYCldJHkhZZEoZXmt1C7ATxby57jVmvAPi6NOdjH5Ir
2FJwe54LdFnY9dycTWRqcBSFaj8E+kckgjQlChXrS4Vu4DhA0KeOsOrapQoZttoYv7kszThR2rMl
LL0eNZasyq7iUOZ6SVx5VyvRbQ6SBRUt92uqRxAemvL17zsqtw1o6UM3Ww3zH5zpZ1lK6xVpjf00
XWy+yCQtMiK4eG2TH9jeUZnNbAiI3kXup1ZIInMCaFPZcxo8yBEaDp5p4JdwMKCIG6HD9SymkdCa
HL0hENgVGc1QQyKKHuNEpSa7nIzVvvAYTaj8LDssReStS5/UcIF2jDRyvzetQ0QEiv/oFVIJ34gp
n6npOBQr22nIK/snRkc2cDZtfr7UhhVOemdZVy1gcDQI+yOHfvPdvDsI8+MwLRCpKpO3iWE/4Jo9
f34uOY6nQKv9c4MwOZOVpTamPyt03S7Dj/dvwrujHUwwku+zqRFUaUJOlZh5Re31cCCU7uBYt16w
UkHg0vnVMm6MqDi/3+65J6sS5uQEkud1JE5Tc+MNDoozfJmlbJFPj2zEDp2lHkxDuLUgrGcrftv4
9gt3ukMh2rcUSW7tRYI33tuSMcPOaPp9NAHt4nTch1Pd5z0jjGImGkqyXj3pobPxp0vsksDJjzY6
QbsmV4M91VItyuUY+tWhzrrmNEYmsdm9/9/GXi7x+BFbCMMRZigvAm3JtPP4tOA26Q+FWDEoC+bv
16eAGtBxECzoqJnWlA8s14kkF7Nx4FV7oY0/mZ/MWjo3J7u2DCnPWJOkbPDZFr0ggmi9asA4JBpc
QJFyBBHLhiIzWei44ZQ/2AFfkhDvQqv60VD/AvouLt4EgzfIP1joJp0NRqjeVKgNTRpl1PzMT+aj
QCQUD/EGsjYFyAZk+IiDzRRDJE2U+lSQdHA8Kk3WR3YcAx06BpS6CJP52EmegWi0ACHBJYQmxVcT
IYE/4J9ztn6qWDQyWaMLcLOWAAgmu8xC/376X6uzRyFitOvwOFtVt7HZhUTXvDFUP3SyIqc4bWiC
v8u5It6Vxl2IS2ixF+TcvbsaqCHJJjrHhYtLJJG16rCXWOvWCsZSZbpFLSoyelOf+3Zon3FjB8ys
dpp9miMCdkQCxgAiSupCFl3Sh98Ho2oVFVCmJGQwywS9TG7h+FnKSuvyw7r10dNPn7nt1TyAh4fw
wwePfz4HVlce2S9z02c1+W7nJ5YudZSKxDf8nAgA0Fdn1Xx638qWeuwfM+/8rW+TQCyiWsJuhyfr
TBrvsNhgjvqfFzmiEculwUu0/MDZdMVg+/R1W3B5NMkjXALjb/1jbudK2QEnt8lOWjcb8SL6l5Nz
TH0gGnTW0CBBnfOgCTSFX0jT6fjJsXH6mgnPw/pe9SPi2Qcbc310++7qrWiO9lLwtoLCCQ3vIstk
WAGVEtC+nM372KHxKc2vepVAr4TdrI8okUwKtxcnBWvRovySP1f9Jvp6hRjBC2pYVvwej5h1Ttxb
5A4PgDhTb+ygu71CuYLjxY4aip4N/xOrL/IzbXi84JweaZVpQQO89O/NcidzzH73nBikUZ4xAOxj
G961It+F8PDq7iRxtYiz5G7FscgjLF2Xlp4U/AqP/1tbxMhpA6+TyIB7PTn+KS5LbS0pBotgQl/n
qHxb39bVfNUNNg2kk1/oB8aCnnQoRpxYFQnHGJja3EK9obAogvaTwtQrXPQn7wNA59JJ4tvycr9n
yO4nlu3THXU6u/454Vda1DqIcO3YAdlwWN9jjQLpiWY8fkuN3zFSUNEJdc93pDpbCavkT6+HzDGa
EUhhqBFfzi5IhqX+aeD+Y/TJtzZFSqd/2PN3vt1qp8dUacCk4dthvECjrQDFxWCBrPv5GVR1dm+9
WxEc4eT7vv8hiNfn8CqHn+jaVB3Dh/JZAYznBFVFeBQWdMZKnqd87eXaqV35GIBXAbssLLMOpI/V
/aRZe+epF6cWxjop+Lfiy/EJXoCanqu15LMmXnavZL59sEqvK9drPohEADX3PdYR6MhLggqPZOam
tv2h6bzCffjtM7XQ6Os/yTyZJ48CJk1yMlRQYyaCAfgjO2ZV4amDN/4KBW5SVxCEzscpR10RusNV
Q3s/VZhvPW/xJcWRFXM45O9VqhMEit3ea0djfM5DLzRCPz/VkXMv1Gv2M5QTvpV8l5y0FWr7tFqR
HfMxZy66SUtQ0CKxYcCPWaz72DDltI50IRlxuPBMEUoy+hkgNdtVHptfzJcUunjyYJGg4Or5APYI
BFyNFAaPIgZmUViCgRiaojMrDG7OCt6ruQVuV5m/MOqlL7Nr6eL8qlp8qMqweJnpGzZeOpE4v13r
0yj8v+ZT50ygb75HDRuvFmewwYJjfSDlM6ecJhh064j8fWdRZtDmZaN3p2HzLoY8iP2FQ2cpnI0W
hRR5hlQWZ79XsL1ELnJpe3FNXQQNxQIzMEcRcNkZ0GgHt7hFxZaOPyGCHXzg6YYsDGQFYD+VnjHT
5WnWNFdp/PmOoYc8/Ubf7fJqF4hfMQJ5MngpQRxk25PBRfo+9lEojdWIMmr6+TGMd02nQKo2X/Tb
h8q+Vbnj1m9kumIjsLGlxN3GlnLv1fR5vtUIBULTU8fNZQuYNAhq9Cslaeh7GBKbEJbn4X0dSFi5
KXkxfCvoLgVA/WfAois5tl5ntqKAZKa0hEh0v7BSiEuALdHpklzQrELTd/YmtGv9SqHx5GS1IfBk
El42el83ZMFG2xdTaqIgvJaJ9QuBEcD6pJ11b1T0QXLasD10y1t763USBQf8Y5jxmcMvMcdyMq0U
bho+FsZtON4ADn0esWrhrOezwRt60bxR4KzhagdYlnZptyUdrwOX4+I09at2pOOpXqKbVU1rp//i
9M4h4QmqqFt1XepIcvjPGiHLYpngqWa+QNtvCEc4n+MezrNkjOwlIplqhRl//ViLc2iXeX5IgyzL
u0vgWVbueEnM13Drm3ARprHwkkmC9d+jK1/aFDJwuXWCaCPdiPNpPeaxMNhENhpZpusGPfM42uhf
Nik/hFaQShCy9gygAutIsVDQd7kr900wpJelVoql9MS7dx0yaazdEI31KEItHHxUl1zrjhIrXGRY
1N/RwkgDSwu57cFKan4nqw/LuvMYtxMljlc6wel8APRmKWsAUKPmc82Kx6K+uo/3RrzpWNTsEFdF
2oaB4uA2Mqx1fv9wjoJYk+yJWsAFTk3eFJ6GxxFmvDBpYD8Pr43BCjSfSoWXQ9XonVDIlr1ydRpb
P+KSWIt8T9ZBO41Q0WvWEoLIVyI1YvnkKU6NFXNtIfotzlyHjF0LlLe6ZrW+/7xcBCQFUZRWP0Nw
PDoYJAf/hBdl7rKKyqS+BWqTHyGBG7gXVUCuTyVNhIJ50aCwA2KdteaVL3/9c6OXHiSFy69hot1B
JZR5vgZaktZ36MiNmdd8NgLWrlWvklBQQPP7I47i84l+oh2/de0PL2dGz0JPu0x1ZsD8YXymBhX1
wxZiL2Z+d/4BMKp4l/KcqhC/lGv0RqV1A/XZZyWvNKj6YGFRc9tDoHTAjxF1WQFQZcEVPTyg4i31
D6QZ/NoiGEkitZIrszGpbb8oul21sZ45RgLqygx1IYnm1uQtu8gm0sR9VAGVdDndUEjgE5+ovm07
gHBhOx2GPKvddhqs2tMubeXF6/5KBXh8vThxpBXJWoTY01MfX6FeoSZv1whSoRsYo8MciFK9F0Su
XNa++FwksGE3KcjrbSu272OJXFzZ0tYbztrpMwZ7rKmJMjX4iJ0Texhv0C4cBXzA2a4Dab8zf4z4
FXg13xD6GAaK45eOhuDxGs0tXWoBLxIK6BmsgLYd+OIHohW8r583FSUoDuB2Q0PMUtAdu1Dv9c6l
uqS3mSOyVLLceCn1I6n0yLwtskT3m2XqALeMZPcG6UhPHKfq+tZ1yKCGbnnT++XrqoNNIEtaL1Nc
cB7d5MnNPZsd94C9llzis+wKCo/u++BHQTRms5alrMIbUgU0RwnD44qNpVsY0XXWM6ryYGto2yet
D8O5ZHsp7GPbB/AZha7j82fU4560xGBJaCHCCmRkA+nfBElsX1MT02RqIjpt9zQlxmzYOxYF0PyT
pH+03NcOPfv4RVUHD9BWOh1l9b5Ojb5qbNHbqZ0rh9TMMMLAAO3D37T5PmPiQU6BJYmmBGWH8dfF
lTtJukOWGAqtOe/miU7euIUlQUST0qN89OtppJwp1BnkSstPsTzz3eqPmBDYa+GvtlCZtcRdthuR
zXzGK99rrpeFYQB7dbuH0P3OPce3NSCiM0LJNd9/WV6DXUG0MMScoOsZwHloBFVhCAifqyQ+0mUO
poIArsj7vyFvDrL2oswaUBsbaWdTzhclp0rPv5d9Mlv2UyOnkq6Z87NNzg9xdX0B9M8meqZ+pQJ6
yPRIoNqNaSAgX710sLdRaiIIcdOWUhYYWFQl3sVyUHvI8Bpz2cJK8ejQ0f1zekHsot94dvIrlQz4
Or9uAeAebE0rPrjC2Z5zGFbeGioaDcTAbFqvQW1rV5bWZfFowgW6nuIWLVYa9m1Yhc+fXMPLdh2L
LT/wMjy4fo5Vv4vd1bY8g3oKKes6qixt/Kh+V0zWTSvqany43wps0/AL3Xm7s/dG1AOxTEZ/A6gc
ZYLW/6vwrlm5KUTYN3W9AQQY+ByFA1DYPYaTlqgCZtOHzIPzJKHccR7tQN2iNHXsMM7py3J4ZzpD
vG5FFEyJM5FPxKeq+p+g90EeOptOd+c//gnWOAfiHtn9YrBKEMPSZhv8ljjTIjBH1WesoPmaKytQ
vhw3gBvY3LSNfCsdtAp1O8w8QUAtntJ54U39niS5uiqMHQzcZK/S0tUB6doBgmaH/YB8X1G9Zeab
fsbolsmrfxVhx1/j9RMC3gWnyfYW2Zw/VTj+lF2v+EAJamipNT/q4dUKZ8xzNyJqNYkUzJoTvigP
+kg9qbc8IlWyp/LWvcWG+TrOIHBlMIXW40mkpQcj73XUBSmLeIt+phabnDbVV4F33eTFrIYlyuUg
hFLUbvfdPz7AmQTq1S2ihk1AthFoVUYxieCU6MB3dFDuFUGZqoLTU3msZwXEfUSM0B+VMLcaGblT
edm7N5T7G8Zuo8N1UtyE3Sa8C32dZUxt+A31MmykM9ovgitDcp9HTQF+mE2OVZpiYSmFDFwVpt1D
dUb4i1vtSbo3h0SIOTfLeS+GBBbI7wrIRRQfxlvXahdn7jlDGbtY6gqlXU+cYt1Xi4KPXAfkM46j
yh1R5SiihFU5cGKQ85HvFQ1CJDtLRG5VHUEgqCIJGAAmPNd7mq308PJ5XRXWjSryyVA4CzmlVNy8
ki3adtxN3DA998jBZiQ13uWYUqwrcyFHabO7v+jQV02ovyZMOrMuAjW7qR4diOsi8MaQkBrl3xfm
Umj1/eHIQ6FZWExi89v9mQzZ2/Ab6R1uDK6v90bYqwmf9yBO4iSHTqeJd6oM3sJ/QEw37O/+kqjP
Wf1SOTYBo0jVbVTeXWqHOjMpOZCmkKf9epcYP55/qRiVW/g5RjVuZA0dig3PQ7Tos5Mx1A7sAp7/
/xxqQDNjDMzNLGExSmZXY4zxj4A9IZZ37+ZqEgHJgfziWUbh6RIQYCffxVPUuTSF6OEBQhKHBokW
+G3aqXoL8F3MT0zx6zhD5LkbSUifOH3kQWKK5VDoqHtG2ILTxsQqmC4txVQxKAPb8RKscfR9zJ9y
TvjuYBCc3ZullFOELTn+IWNqXsEYmYxbvgAWkHmk+N/SxmEiZq+blYjkaoEvvTv+AcKVcERaP8W3
z0OeO4I4u2+S5HAKwQFcVsizt891KZ0bGGlTitO+Y6OvPQANTqdV099WAmVa95kdZ82V5Doy0JwR
SzYPVJWs5y4azS23Br9RS+xzKozGTJVAQWDZ7J/cCebWeaYWIZQqzGb9MT3XvL+HbW1rY4g3lG8U
pTNtTWZZ5yWmVuY8muEh+JsDWUFJ/ahW9evJilo5JxOQTAKKJOYqQJDAJ7skNWkzWuvq6vigLqc3
ae0mX1Um2aP+us7Vv6Stve4Bqr6Ko0Eazw1qGNqBS/TkKG3IKs0Z+1d7eqsOMhUcXk2BcEVLtnjk
pIdrD5PkBwOIHAYonx0/mGQGy4P1/LSDG+o3sJmjL3gvBarm4Z5rOQsn4+nErHdyCDgRiHhMc8mT
llG0JQvcncwfuwE628pUCmu50CPCzoMyY8aD98tLXCEAFWfHLDa4y8Pasuio9RfJXq69S6Cq/3+o
EpOUzO4RlQjdMpX7eSQXeKmtQQOABkq0dVgkf0qazZGz19R9wBKYQYuguS/kVgcuqhUIghZlzXcO
rIsd/lSYOPVWDE8FDjWYvNsexjR2zFMBv+1m7z7+qQrXDANwWSfVg/8lT+VQildYA5j74mGzw/yu
kx6pWqYF0HIN3Z4yYa4F4vjRqY7bq29icm+6b6LVuq9YrCWB0LP5yDPV/mXQVjikdL7CSXfshU54
25WdDqpaAeRbUyTVOVC9Ja2XJXm9HfeQ2JsoIzYS6jYEZyhzuIymMW5pgwr2H6bfiInEruxcEXyu
yBJx4s5esCD7OPwEDTLUdDIAo4JdB2wOUzih/ZlTge93Clbv6h2c4fkHicf7AXWJ8LVpl2yDlIch
z9x1K3KAiUvFCrspkHQQCtH0aa6/dGZP/or/yauwdRqk072IVs6k92vQk5KaDrRHoBztE9kNzt2b
FsB6f8pzKLrzYMjbVOsgi55qB1EJM+ostjYwI63JkrSy1QV3Hv464kP5sjaRu87PZ46u6WPEb2Pa
PQ8jBr2kAXjJ+X2vPuBS28g2NXsHoQTDrQNYKWvZrAqLgAKakh+4/4I1fm0VmO0f7niOax3BLygH
YsylgCNQotojzl4A+ndakScGkAEPXdy8TwpbSMESBG7MOqIBVIU8LxT1zgqSBGZlQire1DQ+A0RO
0Yr7Qjwmm9TZKKWbIj0f8vV5VXZI9w5s/wGuLGeq3mFKPzapYad6vGNYA2c0NwwETvgpAbvut1+L
VO+/0A/a5W1T98PBGV3XOEg4mcViPGHpHMcUu7yB7/DCapQXYA2drYq/LS8A9o7PHLhPHdR99Lys
jUHDyiE+CKgP3YFOVerLYihh+F/IKBuqF255sVjV2fgOpTaQjsiWy88Ta5n5EDlkxoHdYTb0cXCW
WrRwyj9nlFAoCvs3QS5lcgo2DfFn1zuTsAgAgf92OC7FUKJqZPVyocM9T2C/KHj7SxfKfgaYpEBw
K6ejm38VgoDIdwn/iNN3cyEx45+6DpbOT56R2/MjMKa+0BI2GiPhxdCnnefikTyaTE7qofv9bq3J
TdIT/hPOzQzH72pNj/ujeB/OocGC25Dbva3CvvsjuZrPS6WXhtz72j44uPSJZGpXlLocvZ88dx54
m6qST/mbJs9NObpSQ49vPN5xDCr4jp0pCcfJVKxBfim6+vlwHpmvGMkWXg44ZX+cO/Y2Ed8ghNJH
7RSgZVc7wlHBTq+ThQRa1+KPXt55pn1r8em1EHmEb/mr0wE1NgkZpIAFns9gnv4/KX/lQNw8PO5l
nOql77D3SGNZ5ZQukLAkx21n/IPhzhCCS0PIIE0bBq2hcT3g6CmCJYbD51muZSuwxCzh5W/+oqCT
8KvSaIAuZc9h5Jjy2odVDam+0DPbsxteyp+9yPVw4VbuPuqYvZCpN5s1cwggkH47BPmPDSdE5kML
zWDEU1V1ugJGpHKXLQu65M+2Ui0d2Y/0zDH1csoZ7uzSwRwDDuroOG6D5ALjw78lJ/3j6DLnVQXM
WrZ4f1L5k+oH3aH5M5nB5nMx31IW3HBlN0aHimyDDL3TD4rXzNGLWN/6JPOsQLQuSAoe/MQtqedF
sTB85Jse0RLek+PSs+H1jKnC3H9MR/Y8+53Ygmn1OVOLMKUq+557oALicrg/LM7EVBa7PiokwwDX
UQ9qmLN4PnQrs7ZWUTW3jszxbFKkL+XWUiCVOnQA0GUkobOzSCPCZ+W9d+sKIAOH/nv48/y4cX0e
CYAMfaFkb+ehs1iII/ozDBjBoVrhQARestQlpzRkke5917LfswlWX4wOzFkdPrdnMWg5kZEWXy0h
XahIALj+5og+Wjb9jsOBId/VH1wyeqevy2qJO2XWl1KKVkPXSTv+yct0FgtsIZpbnMtiodhgKJ+B
jQtzzEXLY6uXhhbAagR6+IOVmids9vypa2vCS3u1QgEFe7anHiOqxBLBE1eWtuL7gdMLYJCcMj1E
oh5nzZy/GwvAPC2587UDexm8RDe8AHXNmytcUEdeLKq9BoK5wfeJXOc7Mo5AwJmaL+hirPCUR08b
fNntLrRX26OD4tsKIhn6YMeevop4mbmH73qeSN9xuHTtNfu2ElhK1xX0y2yi+5yMUbI+kNgOPjp7
iE2qUFKC8Q+FhWNDi27dSRDsZsKX+R87J2pVuJGlcMO4Rgmr3FV26nP5+hBY3QRBx6VxRTKoS24W
w6F+HJwimHD+zOKq+affJcoGKXdaEjcNByKhjHfl3K0BPKOzRgATnqtFrF74IOcUCh35jkFw4GHC
+dw9/QmwPQGwWOqr1Ix4eV/amDmsGwyes9mfpcxIeqyIgUJMunyru+n9GrfGlM+es7Iqw781PL3Y
eVkhQWrukbXMx261U0CMibimXI+vwiucJdncdzfu1Q8r7ToZ5Chhu3XLmKk5aqVXQPSIN3C4lDoP
uPzZPDlCyBruO79VymNIs7FsCiK/GwDkDBU2kBq1Lcw5VkzvNfZs/jbbhIjZc3/CUXipFubraYIM
2lOHjp4P7OAzjEqfZSc4zw+yJzRKkrCulILnoUiKz8U3pE7G3TFUhc7elzBrMeBHjEUYhSQvX+88
xAHEBRfkkTBTv6bmmv9kNgYpNfq8R4ZW5gTH6nuR4aT6PanzrU0VMeWOou0uAptiD0kTw/rpcUIz
WX3T513TJHFBZAMpMlMDijHMyNdXsaA6FSJy86USLRagUhldLVGsz9wcu8xNPpa47e7PO9pyXeDg
PPDE4kdbMN9JQ0b7NhE6ikw5K9hSjq9JrItheGx3YLGh9x71HRX55KGb9agzb15IzWk2FSk2YJRx
1EJQDxQlApz6UlrDl1+RJDzBf3ZSd6RL7gVP1mB7zO6uqCIRK6mffF6hUkVn6oYMC1p88p+ZrB1u
wZc8X3MiWx7WvXiZn8NwvQnnvXXLlJCU0oIo50Q/7jWUO1mCXh/L+NVDRnfcww/mQJfMFydwhsrv
Bd0LqjBdkAA68VID2/dqjpsIsI9gif3n9mqkAzyn7hgKunYVdCP5be1H5DCaoDfGs25I1n7Mr7qs
++tR0Nq6IpK6yviQwbBIET82+hG8sgQ5tle4qGNXkw3Z10sYm8vwELtkUZ3VUycQd6vV+QA+WPpA
+mBBAkWRYxQy8kZf5ElePeJ1z/LIRZp/2yYUtbfUUYpr8UfP+a8FYRIPxDnJxK2Xs+tFEWdhHg9k
GMHGM2nEOmO6p0kTyjQD/IGbZg+LjmhrEqNkvv6f7rVYSC+j0bUNTIuImcpif5av5ctLVnmUe/Hx
SI300TDmbeoJ7qoTrUxoHP6H1TzgtphAyz8Z917hhNSYqR6rxuMBB9lCs2NC33aZEg3Jh99f12z7
PZbc7lg74Qjnugwl1nA5lyco8XrZ9xhKy4Tq7bblI7ozQgqyWvhnDRQv2Iiic+yw0Ul1S29Ri7Nc
gqBnSS8dRTE2FobB1EoCguE+fhoWpRqznFFdqhNo8aO7X8iOfEsHuEGvvUXLl3GGqosgoFLpmwQu
Qb0LxOw3qu3MW7Ip6A99gXHEHYEvDBlbv4jniLgYjUP2p7pZ4MkCz5mxp9poE5/4Xxnm1xTFV8ti
2Pg1tdz35QQmLAmfdGjR/XyVkd/UktujfsUeTUIhXiQEo5eFKnZk2nYO4wkZGJqE6egHitVNsI3t
r2+OYzdy2I2xWaUDDbiSmr6D8cdRxt3K1QHBxBMzVUSYwAUrE8CIN0w6eg5ASiUSYRm74x6jA0ko
g9v5OSolgV9OmbpASCV+8GYP7huaqgoSm5GhoVpqMM87XsQKAVqs7FygOFUdsi0Ckm4X/bMeBmwX
VE/8pFUgIsesugo6nkAlSPaLHD9XSnW0RZom0QJ9b7YmUixTi9+MkhLpUFWIAcLx1jz9lYJQGKbK
h2UvVISOFBW2XK3Zjx3QDhWrpfjLW2mlHSH6fekSA4r2ygSACqYpPysSRH529LUvNmVCrw3tkyaL
X56n+Koy4vJXYiQjHZo58aTSoe4v4nAqPeH83/vvwh2TR8GyMrBC8ucA78+XdVNTB36zHA30J2l1
droI7Ozn4aHiFP2dMoI7dFbu0g+Sorjm5qduTbr34aFi+gEZULZK3lzUXvx4MrCxupp8O2LQ6cUe
wehuZkXJKH1xsm3dyg1i3UjgvCrT4BGgE9jYmVH13P9HAMYZlDiAklzyMaFTefq+d/RSBSGNWwW9
KTarGCcfseU3fBqRCdJgLMF8qHHTtAZryDvieF79gt0osf459g3WQqWMe7azQ8DZuhPsnklkHOtI
/NHvU7hiDo0ytQ4s4CDa+SI6CMpJx3v8mIvrNrejUO1T4NC7lfS5cg/bh/O427dc9vPFJvkk59dy
KnIWEG2n3FzzqQ2/9UvwnevsC0TtieeuVoITiD9BQwVa5lDpicL6uteseFL0qjUfWTq0TuHD+V0L
DPd2YfpA6l3Z1jdUkph4Dlzd85Nkzerkq9GQLsPk0zuiEekBRXjxXDZU9KAar4utxXN6hVqKOS2G
1VLZKTtk9iFAMmOTakwM2nkXXRll7+uA7sSBg3886RSXgbSRWIEqvcgiqum3qwgY+RWx2Y/tmctJ
Nr7ke77wULi6CXODuNSnDd3fnApBpzuW4sk9Jz+PuWJ+0E3OtVA1/yFg1bnI6T29DZTE+XuXfFkV
EZb9D0sY90FBwg7dpi5o7fQXMQ5v2AiyH99rNC+j4/7e553AmWp0yrSzk0eicVrVuX49lw/3EzdQ
oGcs6lfnnowVKtNCX+WR/US8akMOt6zu1KW3KfwDvufKzIDjignO6klg6MqashLghYiCbBV8DcBt
GDa7Xh5y2UQKTjNkCXI4M8zvrVu3DSjjJcrfvmOlvodZtkBsd8KW4/MppwCSptQlWGVYV3pZe2Wr
x6pXfdxtinQTvGbTHevH7ZvyhkI3QCtCiba96TNR5E+/ReSXE1YOoarHVhnGLD62k2lWOF6/Ul5r
+IjHMra8/EDiFQUIM1vksCgMikcuCXh/Tipgtgdr7YItHRPzj1mWJK23E/khZzcndQ+CrlU2ZmwZ
J1DJ2lpHTLNtj77j+ADYHQGn4qgxAgr8pSAzGUxBI9ZQEwL4O11XP0ABYrc+mzonDFiDhDRFngcZ
/sPZzDWCCGZiZpkvTdlICZxAlbWidINcS3FiNrOsrNti4qiDPwoTVnZ99BUOZFq5o6L+gVsQoClg
HHbC1GUn6TY6D2DUdBr37aKf7Ee6QnSdOwwPl+DRRwiAgd2kml3Hp+n4I4zeikPKv/d1a749Zh8z
N1E01ktLYzoyg0Pq1edLghGmjHVf8Stspm9efk86Q+Qi5US3MS3LCQtkqBa337c4VwJfcYyIbq26
VzuwNcgX8Y2beHtZm05WHdGAdvpd5q3Z++tXUqM3J9uh97vaZH5gQOPq6VcmSfuOrtQAx2cBZjjJ
WnrOJCt2owUJOtdIDJYvlYsQmtGLNLUH0cjR8Gb5K4shDYzSKzadfmH80fjhDyzRezFoI+O+au2b
WSX7SnlvhufLMw3oqLT84ZZW6lxckPD0M0E8og9m6lWt/MN3lJQm4tLfNTwq4OEgUHEZpSKr8q87
UeYOl9XKcgwNvWc05fHWTLX6/6n5HN9+XEtCdbL1w5+vHesuyh/M1EwVY3k1FrLyBk3fMV4jfX7D
NhEsQTXikVteOromCog9Vj6TNjggHPy+QiLv3Xa8qvwZ3+rvBqrGm8xVbWfzkLcTk25rFokwFsnD
eRw9n3DuEKn/t79y3pwKqPDiEY9JuaWURst2pzUQP/UixalCDOTCr2/xW+Zo00ou/kiykvt4XyGf
qQT2koyVXztNMKWlAPCKAFoevxfIiGULBMq8syjZi/a0Rz6iqbvYcUsIfowINzDR881aQMn7cOjt
cxV9Y0Dld/6ZKTYw58ZMpmvr0KZcZaYlQk/jghm65TRwwcKWZiSwRRFDJS3x9bq+KgVNFIcnBJ9y
Jzzs1BzX4Yz6M5laqLpKA4jc+NiYhoZncYsz61M5xxRhnz+cGKFeXNJfdi+scKToKXu60NQE/Sjl
7sSFBvFTig2FCvRfhMH0VpNSAtWXizS/XR9gwXaasXur7qIoH3BIyx24hbt68BJ0YuZckzqTBV50
crCcQUPHqfBwNGY+KgF7oVlo5VOaCDqXjuyfiZgHVFN0IwFnFLfCASskCOBqbt2n4riaR1G33tXu
5AB1s6LJD2mY2AW9zqirCsPjBFcs63mVLqTq8TqrJaiX7Hx/s2mA30bVtblmTCspx7g8oOvegA1/
x6kFEg2Ma7BdtxQ4hGdUq8ieatkSH8S6h0ppwu4id0IYL1LdLjNcgGiOB0vpACGsuK7oxJ2i3r9j
E43hnd1idffp/YudQRXyE2N98i/N3b1QFWXhdttkmeZB03tj4Zt10Y9oFr8xmWZw1N1aZbPKYl01
1VqeLoM0I9HBOivGBNmw0A6J56y2ML1YqxjG3U61AJWIwTCdQuYDBn1lt59UTrZ2z1URKb4G0/++
WdetUP3h94phd9w4CLDa060AK044CNIG1uBBaCOTU1GeatI54OriaUq/7G7vdup8yhYAbIYwklRr
i75vc16dHl80MKVF8OBAcYXb+ZsrdeQgOWAX7CEKUPxIVDCq05uNH6GQUNAboCNTppQ32RS10kDd
22SSAlbQHqybX0JIr8YtmW5RtQpJgKUyFJ8j+n0LcFpwqI5FWw8d5qv9DsQ10BwQgrZ/86gIO8BT
QngfcPmtiCGxI5/aZLPCFf15ynomAbDMJyLJuZzp71lPWKZGeLXj0LlQh6YpFy1ENj5+MAA9S+tj
tI5iIs0gitliCz9JpbrLU4YmOz16phCWZqZTv/p2Wn9wp3fFI7doDG4hwTP7pChJmfu0ohvYz28e
fWbm88y/K6CF2Fm5eSKqS/Cp65iPp9YF1A/fld3n1t+MsHQ9BoCC+bh+RxYDRKhcXHaq9AL4S5Bh
mhQ7o3JoPfdE4+0W/h+kcka1DsBFD3L+tI6+GlI0gGX615F9oMtWoP2KaMz98kd0TLsJXZnk6V1V
cDR9kc47j7Mj62X1H3eU6RnBjkpt4jFbae4SMowIt0+KxXLNhcq4pbMuvpywqwa4wcGK0/TCsLJW
Fct8Zhc07JsyTMDnbHDUEsIe6ecIeaU56LwCuVRygWXfkburp4svBR+00PsnzeFzH4jnm7vdtoSt
ilW1O2kZEZAC2xneg5UL1Qejp+AEn1lHaqCNMtSYqnsYTodacYO733GUxHgQKY1Z5zY1CdqE7tfY
MwY0O8uDsCm6MPDANK1BAuSCeO4GIbIQ3mLWGMfOU3KODwlc3Js0Jl/4cyTilmoTTXgJELMGAt++
dC5KMWGFAnxxRpZrILoyeB5NAJdTP2OWsf+gfW+bk1CNjyVYmDUpvzmFQSjiaSswnuaTWC5N7lqh
72mpkf5TxwimsZ5j+oaAwDHKDN4UUfBmsfrjZqx4mbr7oDHzoV4NIOctp6p8f9XWMetdpCM28UBc
St7nm14nPDZ9JFA0tp13hqA4wYNp7XQplcLssU2VHrIF+kheSbBkAlCXkVeWnZwOw68mzqiWjAYq
00HCrIFFpk+H7rf0C4ccakezIM0uBVLvTKWaBT/Ha7/C8z5HGX4LoQ+nPfoR7EFun9DaLjsiBbvS
BGGKWOZFXC9UKbGFTFcJEPdp+PZXkT2veB7Y9FOHnO0kiBJe0NzTugSdYAxy7vRGIVisOxCzFNGG
8YnclmCtoHGkmumKi5j32hRf3sFl5Vzj0J1PAk4AG+ftMpasI9X8+fRx0StSCDA11HxhW/hhDiV/
0tUTnvFsLk13AN1qN5HUxcDF5dWnemQ5tYWJS6UZg1vO84QD3I+ertEuAfNkK1TQKxDBRFMAoP9T
hsOqbXwFvF7XyO/+ApoT0ubKs6EUTnYMXNEXm1fWI1SMwbtdGqDbd5NxAiLmkKABhmBI5Qkkx4RI
yhoqvZGDp55Ephl/CrnyWWQM1/Bz+0NHLw5DxR+aWAvTEWfgUFWk/9eh/OCiksLWEn02MRGtruMo
FRBLvx8scGkthuRuSzOKPVDgYs006ns06ccxvZ70rkI4zkT9aK9Hb/g505BTTg/FvhZPwU3eUeAw
nIU7g7Lp0MHfzbP2aXnMa65rZ4UVjY4fpEyMl3Xt1I1nZeIQN8qaFhW121wUreWdic3wBiV/LEjA
cCUwIJuqSt1tDq2FLSbRCksxo2DkqYX7DeYQTfwSK6UQ32ddc6ukPm/d7LYSMNKa+QfkNHnCH64q
4F2k4jOM00qUaUi6re5+2u22WeuuRdEyOcF/Xigp9OL0G0LTJ1Sw+U3Kb1SyzHp3ubR6IGzb7k3L
1R8XXX3lqZeMY3BiWzXAtkoibEdR6VuZ2WwS5Ngifj5OCoNZd/ACo0XJYEZOlFONUwPC9pG76xml
Yq/i2UpoChOueb6eY69PTPhu+jwSaOVs5n/QeibCv092j8HB7lLVneOnDHbNcOPViWMmhDX7F2zv
MtuyIXiCjaynII2ezrDcS7UZoWpjpWBxO+qNdFWs/mekuOz3uonwBmhYwBOv+OFRA2Q3zTrMtGH6
2Zgl2a5DAdjdFrXwLA365Gz/P75la1Rm2R5WD8OYsx9bJMugkwKToUboZhRG99YE+njX2BX+CM7B
yKX/drQ6Yel5ATyL8qDswxsEKi62DV8yrNhXNuBhQv7nQrI+YhJaDoDNwzIYEiyMQ1eRkq6zYM8A
wGNTomJ7pFDNP2FB/a8FhMEAiSs1AnQvXJN2KrYjCjJyBuJa/BYiFXVDZCirl7nVoiYpdBBc32Wo
mU3sKyKdhKz+LzfjhbAbWE7hTsl2/skipukHvm/unitY4YHReFUjEAG2TKNHSy9miONVgK5jhqMm
1ShwqEbrpClN2KqR3j8zXzAkH7vWOmkjeT6OH5PNwRsIXgH0LpUbnGZt3jtLs5T2L89KDsgcKnJr
TbrN/lNmKSX8MoX8wbxylvW2sz10mYlpDKuP6IIqG4HdB5OApmp6aA/miD4I28OQeEVnqO0qVGvG
1h6FCqVtFNR/KObNQ+xFFR0eRbE/VSxAzcVEpi0ZOi15eRUP1hn1AfBydnngAZm18k6WweTHFL3y
BRKjVaY1uWpldgD/lVld5vZO6RGgUyHnahPCcfIRrXuFvnwhU//f3aDNQuX3nHZAIWQiJ3HoAaCz
BD1qff+27AZltvAaCT1wlkynaXBfHjRySg5uwPIzAIVhFojSB35aNyWHF7o2VHZEGe2M+CO7pSOY
V5YBx+Rajzf+WTkQtycJ+yiMPneO+mz7/mJUfDGXlCxnAcce6pVasWmDxLkZjqdv03QTuyP352s3
qJySVRkeJMFuCtHwyHjmiCxYMp2V3xo6NRHRl5JukMs+whsCSYXIW1Ec0mQp120Y7TJjm8HqkAVN
HO/FBhUrzI2YI8I+epwJfkKF9wabUwEJ8V0tVGWlbr8RIHZevLpftgMY3XSmOWK7pkXlNjNbg3bk
0QG/hHYmIR/OEyALQM0Hplin8g44ai+OskyShAo7sJVGL+VtBha04M/8WtCyCXQX3dQTggbdFuQx
LCmpvPSp6y264G7a2sJzzDA2YUM8zZyDmHBXRsD5dfQ3//PccZT+Se9nmcmgF5Ol7DbFrgdwXSDP
qEMuFeU3Vd8+BVoVJQKWFrzjVxouPvdBbzUEa/2VYbZrErn0AlFoZUtR8PwWMA2HQH6mYxK3zss+
aUO39+Q/neVKWdR4FvPGZcJzlITu6NJuZSmsHhuG7E0x3hL04lZ9otEJYeqXh2ovX3KOTSJ7fuyf
2NpvrrNwjl+ibZaRpGoSVvt7MwbkexgXgxvrw6yVyh3vL0RgzuW5wZgja6LBF+ipdtjQDZHLd1R5
lKwLc2MqHPvvLSz6jqqCV0DOoxRwjzCNOf0XoYTPvThOu7vwCvrvslfTC+23NCViVduPr+V0NBE4
ih74Kn2PaKrDCCnOFx0UVuNivBEGZ1uXhnst+aKSSsqZUgKUJRIaqByT6fIXfNlDu8D6kwhGOilS
WXD5TXqOhICGfXTkkzaoqfQBDYUtuffB9eBGMf/L1pHWPhRl2edTulJBfYsbDEMo3jXKV1bstTsj
xeAkcBnQvmx0us22k5ur2buaNRVKYnUoP6ZnJznBAud8iiDNq0tVo6ZQfdVVOhrSki2trTxNaTgq
7dL8f6VpJbd9Uv+uCptT8B1OdQgW+sFsUbHrXfMcYQ1802j4EfDvtQLM9pJF5CzqVxrZ+TBfHSu7
l0Vx89kHUwAfykibQwLaSF0NMZmYBMd7X73CG6gBZUQdY6zdURJ9WY8BxFeQ3u/d0OJbVlFs1zCf
k5P/jME+qwReIZtaDtIaqp36A/3uPslE74MLGglq523kCtuyogecFamfX97+xuC7PhA1ghbnAt0e
v89YvIupAafr2YthkmsGcMKjnuCqMmOlGm/uHabpXvOXfZys5nLAdnBaaEz0sRcZ5VaXYoB3Ei+g
3fpMdp/PldZX3hA00MI/Ttub38ncJrfCHv9C/jOQTlIVnvEeiKQ6d+F5teBelHC6F9xWu43fYTf4
ay8mAYcsWkXBC9/sSC5T8rhJBPXTVr4ljzyS2K0tis2NJBFCIA46XLItiHkhvasO2fsZBkDeFu1K
4UKvCp7RwINnVd/xlLMTGPz+fjX+LJAyxHfZOXY55ENMp+7DLD78TQKnKLepX7seYwDzPDLJOk73
VS+doVboQBfLmSmljIvD8m19l+oh+IAj5onZJU8fZv8K+EcW3PbF9Z6h+/GyW4yuGynxMKbO6177
cMSlms0aTQsiweIlK0n/JEZfzVV3Gmwu46G1TQHQEpmTNGTo0y7rrrl5FnWGRtDgqTqMXuNyarlh
Q1q6X1NmfcRWuZQ9GzyWF6rQNDZZF6iCVbZpRoVlFOhpsAyT4ky9BHuf6tVlWTUB8M44QMY/Ryxz
MekQ9dfnXgkUHRQVHhtOPsgitZS6XIpTnVMj9PHPy8mcIIZSTvg4EvrP0aH3dghgOwDYQDRqWlu/
ay0UXgWstJXJa3WJUGBW3uoyFiwoq1Z2mA3MH72z10hFEmeRab5j5q1LVjCM6Uas4N4E7A36BxiE
Awz/CAR6F7bLKgOOQIqOlOKhQaZ4G1e/1XAgJkh82PfgP0BInDg9Wn6asONTidHeIUd4GhU9Wn/m
o5mT7jWN9e2ouCcLxUs4Jqr31C4YGOtk+D927IHnAnH05YgLPgs2LuryPaRGR7/3fut+4+s+aAkz
ppb+gO+wTreT6T3W/hW27pCbG80loYZ3e0dZ03cUwxSSc/xKbU0Y1PRqeoMqxOQSkiCD5CaUXI4N
98CdODcPFNmEXG+FSZAu/nD8SVXjCbbBmwvEDqbU54awVTx2PmECCxy6R4HaPEUyJGSPBfwO5bPK
C6WYaBLg3uANaChYXuRa4CA5Gx8keg+k79Mk+t4brCEIu/16LOnVlVjpbhY+ejjC2/FFpLUgkOSc
J3nCSbwu0ZaeaVGcwmWdoE9Oh5knRGCkEUHXucvqKcFbJRzb72FNDNPK06KisqRgBfoofa1lYuLs
tjyyR5HVVjHj8Y8Sfo7nIX5EQSnKe3olnPQ4VZkirfFno7PAQcX25lE80tjRLl8LMr96qm8vtFaa
BsAG72f6sedw9fuSpNnr0B3Jl6O4KR52Gs10OyFmvl17M9CgBb0qKk/pTTexhe1Fk+AnXyUy0fa2
4hKnImMhwTBsknf2kDnWZiwpHvzDr91W9wcrnK9gB0NHiR4klgAnovPvGK2UTl0qQ606dA4a9HiK
S714YKQNzJV1e1elDQYH85rDlEgUKigSVIGoFXE/Dj2dM8++dtj7i8nMnoud66vW36VOiv0o6bSz
1iz3birp/VROgUfHp1cOR2AFNZ0z5cAyMO0DC4q3zmfko1fcn/ybK06hvlNlN0ZrESyxiNDIrnx+
y8YSRvWboFU/2OKacrRDtoybk5usGZL/TcyT1EQAULGkBDtLjhb6QA9GfgIXkz5d3F52uX3qZD1I
/1s4o59UlgzLraxd8G1p83OESh5PFvt4roEqQ4DKC30REnEaQpAXblcXYQk0QjetwoB8PD1DN+XE
FVOEliZyy9OJEq/1hf1lQi3BmoNt114b8cHeNNU3ujVi5gBnHrrVTiPi7mPJBoSzxs1s6BDyFgrN
Erq5v5Lg1LvyVpg9pBWaxago4Y6nYAss+BDQ5R3KMyQJQfM9favB118aWdKw9kXmn7Ge5Q/VBoM2
w/PHJjZtskupfPO4ej1g6jOk5um0Ikhpjd10Gza8yWVRSs/p5QG2d4rIDf5EhAh2wTMkLRZou2od
tjFAVJ4Vy7e95A3OiyNOA85WBprXb/mjoItg/Hh2c1uzJa5FLvqiPigPZU3XMKybekWwFNMF1XoZ
tp60X1HDfrcGbS7uvoI+CGKS7yGT3eM9lzjN00nY+OxTeJ/BQDIZEoI3WCj9TGws3HXmNXu3r1+b
N4+1bV2CyI2oeewQk+wKQW/akW7zuhaECtg4jJ3rEwOhzR9W6evdedYSeamU/jnLnJabT0DA0nUl
UveaGZX+O9GpchQDrHMH+AGoT7ykIn2h8of3CpDsSsyGx+aBJRIdF4vw/SrdCUpGcERJ8egGgE7U
oxlhltXKaFXTKP9nF3P8njEwLCD2ljFBv23DrAQZ5OPkgPuumDOiDkk1KoK9rnSwX7yRa1JBelRk
8uU6tVU9ZRrrNkMT/cPRXjFg7RX22xdYJ1OSqZEE277cOK3LPCc6QIQeB/r8B9LQxsCctR2rvi9R
BoGsHrrEM0uE+l5Vx2YY8S2RF8sMUTBq1lbTsV9E8u2NuidqGtBTfX8VOKtAFUwhq8YNu6Fjm1JG
G2HJUIWerMRZnv5itd80sfR9zaACkkjEKTd1eJyf2DPkB5LDv+bDg7P1mG6AUA17yH+opR3crXC6
nCLbRvyz+gA+VAi9rZJBhq2RSNn/UXWJDFUxDxcZLCikcumwqisVCHxophuZ1uiXEFKLb3vQJbVp
Uot/iBIZ3TeLYluEfolyU1bAXtUAt9taO6KzkCE95vRFpgJFFV7EbGQ9NR3zDmpm7uIfMT3DiT2w
tEUHYPRoDmhRvAFQju9fyQ5vaxJ+kC4+dQAd85ceS3FhK1naeAg7sORqjYmjzutQIq1nemCoHhso
+ywKfnldlGvcVPykCmchqaWFTiyo/5jGpoGqmrgT/07hx9n/4fIUDpAR7BRoKXAN3xL3TOSeOmRg
imuslAk/pTctaftwYsha37LI/Swpa7LWCWdvgloSs1Q0O8ssKYNApZtzW0bN3B2LTvWKCDBbRNjK
HtNERxGb8+telzhiZdWI2iD4+/xYXqQALLKhR+uFFEks4DMDQJj6/Pyj6E/dAl95G/0LP6ZWVdHX
qjZtGwBsriE6UIt3yN5S+RqUKDVEepS/jDfGcp790A3n2ENlrb+Rh749TyALlFepgRbRstrZmj3j
gtRw+z1YmgrCVNYxq2NjHrGGm44pc1fE8l5PJDASjedA2liqQL5VhENdsjpvnTifJL4InRxYsTnF
TXjsx5ovfH9Js+lYeZOF2sJgw65qArQO0Da6Ys2xX6f2uxxh7WywrXLht+EeKznsQTvHhQjkmhlT
omhIa/kQQvEeJWtqemxSdIHepJttlECzzfUPi42w2mmG6Q7ZrywoHSMBohrjVwo6u/oi4oho7jF4
Tg4Y3Z3VNaoPdgFc88/TBdprxK9Q2Kq5P73dGmUaPEsxTORKQzUFbwKmG5N3FEVheQeR25LLmoN/
eyXKjL0LWWbLkwaaII9NIybu8MvnsFuaYNYkN3KFT1fKPF8wuprocKa0McPU9tMRgWtIH4hPx4IX
W+6q3nJXHp0NlIIFaVczA4NbM7V8Vk3ksHzCy67lfkG05Y4pVCmF0xuZ8OQ11dBb6Cg/oN6arr5Z
RKJxrKQsd0qMJv3n9Lg2Ly527DKGV45Sy/dsP57wEkkz4zxqeAqjgX1mm85NnlfmTsOhCTkE920M
n0AzEtzdVf9yrFQgZwrBR23kXeNeEIohYWFkK8y3ryTRguR53a/nTCbD/zEAPzxjdAclLXum82/w
ehjMFVKJMZCpdJARHnfEv4TjY22aXWg4fd4yX43MIgGri34mpR57oBNGwNq4PdG7erX17i5QR2zG
vvrrvQN7/oSDLtp/hyUDOnDjY3PNGaWKtRtkOHvgmV4QJgCqjmjGGpMkv09PhpIObq9CaQ5tg56R
qwEgibVz9ARrmY6Xe2UNbehato4lxADLex6ZZYdmbJuyFZwI+zuFjDPLyCM316g4QxoxhaopiPl5
PGLHO4quVDW8WSzKmunsxXyZmjcw0ID8mfLq2mmeyUD2yC7mTZfTXEwpKVEqLpz+J9e+OzB4qXLb
nH2/0AXXHl9yil/s16msY/O0jHyYmnPYg+cjmDt4i9xRMRWHjEftDZpzG7vdX2yZzHEOruqqdbzt
AqRrTI0HFVqcB+8TQ06ccVUnCFhzyytvAm9Vqz6UCE7lm8W1nGLqOCl35fHptfOpbUt+WnML+rWc
yzikFqaxtp/fguofStScA6v7bSy+urUoUwUXcCrZiO0AKFMBIclqUA4xY0NaTsyvkeJnIH+dTAK9
nlEW+8ORGg6LssGW62RQOI4cQH1ksszhjYu6wqv/RtidY6/ezWwErErgH8MSL6Im+F+noSuPHGej
1I28bBjdSHTXmBaUTZw53h3hHg0jL5tPcsHCFezd5N3QYsQ0XFx+PrXOd3Z/GlCMZwAGePRYsoch
pbegAvAYhVWOIL2ASqVKQvdNqPwSImGDruGQ7Z/QkgH4a8Y3YqWPwjfmtoYz+MCvxMeMlfi4sHfZ
FuYA3bhYH5Sn6oLYdlrq844ZtzTUaStpQ4hql9751Jj2m6dzAveD1RM8V+m54P7LuVERN1bbEekH
OC6B+Z6pQXxHlSRLN/PwNeNhlNypbpfUnPDS8jWI97A0309hh3XcR2b088Eqi29XI4T3BEyWCUPW
jBfjOl2e/rFj23bK6b9/evYpGTK/9hYPpAft6wg/tmUHP6PbMhRHTejxhq+H5YCuL2PeSyyigbZy
f4OC3IIg8whQbhJPV20DnjYwV+uWbRTqRzvLp9pxVkICjRVoGS7VZS0k+rTcKq5Tnh2S+ALNU871
s44yicTvQinDzz/keGHUBBTDkKTYhwy+2WwY7jgrth9FZGxqMnEFZhjTNnVF9A1geW2npsdzBcxx
+4NnPbfbdHl9GlECXFne9k0ABhe70rsD4M2l5TKDS/dwqXQiGBZrv8sdjRT6ckhvE+uAUCEqvm2+
DOQgXd+e5CdRDIfwAyTsY3iqPD32Uqm24xTuYTGKVz4rI55aoaE061lAagudYLlrpdKJO9TCF8df
AiJgVMEriyzUyyVqGaf+iIOdL3nTuaidqZoP6I7W+vXCcT/agBgzlPAV+abFqJ0rN+wEC92hCXJb
kK/q+ivZKl6rVb6+yZeQ8LVxr7U2EokJ2XdAyh07WLzSx/S3VvSJ6gQnW+PxGf+BjYkOUpUu1xxM
pzQutxbAI3uXVMvcRyfFff9RQEMhaLpyAcknXt/S+xNDe4hY87pmSESyznpLJLXfyHXOyVpJlf6r
yjEEu1YfKMuDupLSReAjHO2CFn38V6Tk6erbu1wWoDRcRtTSXnwaf1gTgng37EI3LvWJhNfIP2md
EH+5lbZGEnyEuqaqrc5SQFvpRZgn9Bs14WSIPDWIcczI703tHcXy0sReCLCIzjUiPhEriUudiqEV
leemem17JKlFMnpYWFdwHH11/cp96pt5YjsOb7XAKJAL/H6dMTKs7bfULqYG0ChJR3BLR99u9Y0P
5xJU1BWrUesZzCfL3okdAUcnA446cla250QQNF0+S/E/pXZCTaMYJ17bjzKHpL7Nh9Fg7eqYdyXe
otDHUSTIdgHWnsZTdSfHAPWpE2vE3lxgVqHQD8/Qxo+JYyUAGuexNpNbfo77Xx0zxbWzhDtYmIQ4
mNF906KZLk0W1QNcVPj4cF006HqMELOOsXlEpTkl/Iu4xW1ttLOGNx28iXbskkm7zUofeiH9TS89
6GMnJbvV1OfkwUVJnR01kGW2LPtqAlE1h3PShVzh8DhWY1iqpPvjUbWeuRzRK5ijL7DHVVYQR7No
kNDGxFTaq0zz/hbVPfo9xBcZ4nZUYWc0S9l9wKiV42mcSVbh48hLk3ywP+Zds/Jzejb6fDE5YZu/
I567jZPWl/veo55YWaMpvXRo35f0SFV+Qrv6nviQuU7O1tQeHXzSBVi4pSpRcmXZMaiy6bzqrVPF
hWv73J42czfvoQ8bykiHJNxqt6zTC6jWGWRL49QS/UgGMIjQ7tG69HDJskY/eYfuXgovxqYRl9ZI
Vv3UNt6TvVfOldGm3KC8wDoyg3+FfnyhT+cA/6BiN7XdkFW2do6OzwWTb+NI2Lo+wLZ3iLAp/+fM
sE+HgBv9PMn3lzV/Grhscn/3PkFDG8L2wjOnBXtKqT7S9yemfOplRzSsbq8HuxJ/8DZpOnDGEV1b
UtaGoy01J0k+UkhJ96/FogSC/5X228Bh564QE3gXJi0WWo2LRdYQYWo/5NdoIh4ru0mt+/8/hJVK
gz8L3+SHCn3TGWW7MD7p7NAU4AmUBW2wE0maWVeCMxMGSXtWvOIA0/87TARh/K90Sjf4Syeg4PDh
KwoTgQItS6b6gowW3ayi/BX6nKZXD2Wye6lLJgFcqiIIxcJkRYJxzGEn5mazbxb3XCLg65xwucl5
nDWkNDp8EMXMTOxtbTz4gDmBd3ryQ9zAqkIoWF7PKC2LzK0MzyTMAmlPTvhPIik03GxgDQYb1IBf
+RkDtPsssT8fi7pv93CLgzc2Lu42SYC0iXHUff58zMgZdiIqjx/UW2CVR6pc8vzQZ8VOVYPOIxBg
+Ja3KTPteH2R6IRJXS5ZE/yG3/HqwB9rSsK/2oFPmB3x2Tj9JvHikdN6sCYLSIaTt+tDLsZnBCcC
sLeshpivOVpR/QZ7vj+CsbursrJG6VLQUsDjqVNOqvnlMDTDAnRAmKcX7e2iypzqRIaxEC9OZ5nh
z8aoyEAWZQeMgsZ1w2ilmktVIxuRdFvZe0m9qUh2pZWTzjEnA94r/qqRopEAgKjoCRV71Fu+NIMX
VQUdF+inzC9TptzBLPc3HON91zMTiP2T3llYmLdsNPl9oDrrYdjDB5LmCtTQt+bnStr3eihumDnh
vv+d9gFkR8EdCrgnJMZkWqaUMgGsS5caXXV/bE6RUJM0KJGgIWIZbbPiaENRfN7lKPCLF8w7bCoL
ES7QiO7m6KVJiTOJPeHFp7m2xVR4pTVb+L1fmdqUsuUjSfTvVIcWeWhyswGwTmicGVHp9hmxM9hQ
CPI9+hiGyGvqzXStRS7yTsnLKblrxrgRYs02p1WvosmM8OvzAT5L6qtyyzs4fE5+X+qui+qTYVy4
Hpo7drSqJJpSezLvUsQ0tjTE7thbTZQWvhyXiOLuh5vh92sNHlfX6JPIKZKaStKQSgbVT0pHK8Lf
8hazgu6gzbMguomQsEyD+FVfOuVOduYwhD9SNdsWycJb7NTSSCR38iLusK99LN4QsYv2VttJRtoJ
x2gGQObHPBKEvQKi8RjKP6WOZwUwY+XhqOuGyglr+FrSwKhf203yfYaIgR52/Xj90O8NqAwZebRg
MgNMKsUB9k4g7+wFDy1/QceQcqM+hdAhDkSnc1Qbgq/FTlZ5b4NAR/SXprPypUJD4SWKiDrnjty5
glsk9A650G/Ri4m+H5K82z+Ub4dreL19xDeX+R2GcAwZxFuxNPpl2u1xze8Jk3bhF9YbaYaISzyi
35vBAs4FE9rjwPyL142OkqynOVmBZ7yaLIYFbl+v+EToHSt4MeEQE8y8sVwM5jqnAGz2P0cccVkn
SPpnGJEIo9DHBmtUU86/luGnpdjjZAaqxcQMdnL9vTkM4uEVPj1g70CIiqc6fBxD5Gl9e14daVJJ
UvnUxAyTkOhYyh0INeVmG99EQQRo9sWy7E0V3xy7IlF/tZb7k+MCLhlmNy8+PtBdGJozkkYqkY/O
pnXWLlN4FmR+8kQXFPyl3aqQ9NpSk4e5aJk45nue1sitEIAQ58UfT1c3MlrPMnK/cUUhsc/6YZR1
i20twpl4gXc+pyMrft9GKibYO8GxuVkDs6JTcflTXCcEbcOz1o+Nc/xQBJt1m0d9WjfhENuS3Nqp
J1/ZWRm99vR6/rosKcPOXTTvlOOFWZ4j1j54jCU0NeUDSoeQHRJHhOVcAeOI2aukaxI/8n5NKFv9
H43zdytLfSPV+6WmOPtZThj9aylEWGRM72UjHDTDziGutXLl3IwK4SpeyGLdmepQbOoYGYuN4PsW
hsYGKAjwtzlpeFYoFc4LTDt8TMUT+F6RC3ZrXbWCsEVHWlyOtHjnTmLW4Eel7EbymwI9zdQvIjS7
as+K9fdl1kqlVban/5NHy85eXKHcFBgR4Bz8i2cjYYjAyM4j+T5z4yuPON/d8xV4WIH6O9nHNo6h
yJG380uqAn/qeFsI29Y19dL0A6A5iWQrvvNzJnbtvJocdjmNTZ9SENm01pXhefajWgUhBlLP4LUe
6SXCp0YVEbQk6CGKb3I730gK2EBBvxudT2+i3zO6AgssXORbYoMlyGPVLy02UNYD8Ck7mxyIYR1p
t0bxt/wvE0OidywDhEPHqbevM79mZIbyift+1Nm4HWUwhOtdFrdIkB34k9713vZPVSJz0eOgLDig
WX+fHUU0yWazf1H0Pk9ShxqJjQueABHUwFHLWeQwxCRq0Df2WOpNs18e2fLnFiQ87VfOcTl0cnob
hZZjn0FLUvXPG7p1FkdDK8u/dCvVKqbs5MXJPYYrlrLwLs098lWkOyBD2a5xfEYILw/0fEKajfeJ
soyLf0DHZ1zYr+4jQ2UHC8VXsu7xRTbS+S26jxivDEHuMj9PkKKo4rBo7vzTYyJMXbAZvAn4q1Ky
Dcdy6SCTOro6bXAE/Cyp+hgGOPssw23oUiGB+HC+M4fX4zW8F1g71BSUpf5QgrpWaPdoXUI+t1gt
NzFR8unRCdeq/Eg6NCG+vemCobsGpR0dxK7c459PJYs+RbK0XAHhMJGRFbj7HRmRzJiyU6iJgkrz
6O1EZZPzTmVLPhT6B1drSzsX7LrVs1yTJW+CnsItMACwTmARfhW6wkJS6V8bOn2Zc1k6LZH42p2e
aT8wcjRZB5N3UghbyO7xWZ8m7hr3Fk51rTyeVUkUVhhZiOykRw5BAsIEjEBzv73Tz/VuAsTDbzY6
b3PGz7Iph4WyT+5JAta/3kinEpF5gqYUBgrXR6lTmXXicREdMGt/eCP741mojtAWMpYvsY2oGPzA
8S2U2NMaFU1CyF90UteUwekT0M1Xaqz0+RMJErrStIaHOWPAHM6rFoJJv7odjnKjRq3kt5IobALT
FJ53EIewDPe/DLZUt0bcxnPfkr3sCkiZ81s34wtS8LDCjwuBqUrv728WgJbHOKgHtonN45ogoI52
redo7B9Bk0tSpMYXHNkyT1mUJ3xoNsBoelI+MtYLyuSK5XK4gJCBPiyKzH4OwhHjUv3gKTl6DpG3
acgtbB31Fpce62Syfw3ZdZTOtMZIyUaoKtz+eA3wt4Om2Ht2HdnrY0e4zVMeW30Pxc/gWr9mtmXU
6rQy5VniZIqKVPU8eFgiRi+CX1aAOz7srjj1bFpVKeW8X9rv14pWgSa+mwc+RRSy2/4jafA5eu3/
ZhTzglzK7hAu5FqHMYt6SdGOgXIt5jVxeX+s0RBMngruTqDgXzXdBT+8PhiBIQ8atQUCBK04COUH
3w9Q1qanGytvkQeK5VbUsjdyOrW/tOd2g1nk4t9y+jzh/QnK7X+SxC5vqyOXdFQwfRWULprxeVZm
DZ+qAlvWvMOMCrX/ksOUKXGMIQ6CXK+4fRX6ZHcxPOUqu1IknRrsr2/XgKY6zP2AJxOK4rWzko2v
zVKb3pYkZGnmKTFci32Lmrr14jgrE6uY0tg30lx37N2jmmrJ89wedgwitQRYlRyHQQkzVhQokapI
aC5nVJWq8zvqgi7VlD9mt/DyHwdjImvW4YmBsnSCYt+/JG+mJSaCQnyvEhH9q+Ih1l2630z0w99z
ns+zCoV2UwklkhV6ZBcsSLs1gB4+YcdDBfhG0Wa7SdIkGlKSEJM2rZbnilVO57mgTXqeMUIiimw/
g8rYvm776bUK5zUYF1ECReMERfElf++nxMwfq1ku/tYJ6fEoDOBuu+uhBBNyphZlyVJmCRKXLzOs
fZmTpHdPWMe/4g+kPi7CMW+d53g51PdVX6O1l4jMZfhYk0xpDf1M95pINJjz+L66fTSL8wP7EB43
ALbuOjd42HQgdl8anULEeFUGHA2Mr1W0uHXKMsLIlmdA/JbLcBkEvSZkaR3uviXd6c+97K5S6Atv
VRO37vNnci/eKum/dcrC3+VyILrRB51K2kYsa+7nXRtY6vX/yv9CCO1tmi6EKAIxLTEiAsji1goe
VN0UMCfJtPt22v5f62X03c/lSKLhXg4jQ+gDCiSHQDPpDE9PfJVKoLiHL3hoBZBKQ8my0HYGoMHm
JxpySqZMg+cTX6IVLqCPT+I4VvyyJN//l2o28ja1jsKBoZsMOcGSdPc0wAKjZ08VvX/Lvakwpnu6
b5f1cYt2749iTrcNAO56rQC7upX2CXyMgjsg08uoarRJLwpsN+q07HRocZUSH4iyj5YkDXSlfEwv
G5kxuDq7iGwjIiCbct5lxt2o6HjyJ5wS0XElCSWam5Sm498fZa967YVo1kVsSMGcFVwxNl8Szoe4
udix9XSiiHZXevp/bmjn0xPZw2Twl4gfDFo1bGyNRHaC8oZntkJ29ZAFOYDFve1uH63qaUuGbPts
BDExwn0cPpt/59/IaF3pQrPpoQR2KiFbDUeSJk/fsZp6dJtvCOsIO3p58EJD+w6IaolzVcu4O91E
cct/GSjzmMISdCp6EOIH/DrVkomxzqZlQKadtq35zTd6rln+FZX7r5zk6wZXiV5aVAPUO+P6V5Gl
7Ntq50h/vTyjQxXn9+lRo3694c4X+57pAsXKkLpjtdoGGVjdyEUMn0J1nkg6BNoPyzyNapqTRSad
3QBJ2SCCikKcXH3PlImpNxKf1A8zrLJ+KQcEFvOHEyTXYj4i3LTRhvsphWb8gJSPNfG4/3qx6Kn5
HuxXtz01l50IJ+ZNCEW4loa0+q2FqQ+ewo/QPODgMG/9DXleGOD5MAhfkgtr1bc4fd7m/9J1Hz/G
H92g7iqTje3fefqa1lc5cITJ+CKdyVUgkcFz452zhjr9XbilhaarA1H936eN0xeKvjc2UsbAwvqA
A/jV3UlH9WTDS1oX7vLDI2GMQzwHNvvMU4k3LPEro3r1TV90yPM8/3BRuxVF6gMGxhFD/DIRIqSm
9cl/VV4ukhQjV21N8pM+I9nS01NvYd2gy9aPNZKHnWsLTR8Et/uXQwNd+56eqvMzHzSTXZ03hV2S
2b/H6rW4yb0j3VbKmOlfo8K8D7dPUDcI3dZzbQZpQXrwqINd0PqDypxK4Xxt6HbKpsnlAchOLm5g
IuY8pLJ4PvARUx0VHKU+qhopi2Vv+NItczQTgaEUvbEguEeZqzYw6tvGkTEzM3D77zAVWbUi4f1z
pcBO5y1oUKd//cSIfuLB4G1eleSmNYs8VLbUoqMgjwdfiA3+Atg53B0fMflD1T7XY8hxUZUfMMZI
R4G5aqViDRIY+FI/+7jwzkmUDC4PzjvrJFmofOnAGWz277i4/Pg9K6iUWHWkP5KnsxIYULK6SQOw
2Q+Rv7SU6k8H0qsBj75sgnBS+99Q+/phNoCZv7VmvoD9xX+Bgz4Nykri3pc8ygjbGXdh48nxKmWj
3+6JemJO/JJEmOKvTcp5GZSperlbkI3OFUDWM1XFvuxl9bZg/lS5JbLooaSg6i+MVLMuIVqHvzXZ
IYGJRFJ4lRKKSCk/3XGSxmlHmc2zWh95dg7yzwo5s5DAtef0R2kbwJJOVPRsN3NChtd1DNiRRues
PpN7kr/t6J2X8X0XnlOKloMR6JhHsQlOueS+uH3AT8HFQ+XygDIVYfQ/xeAdiHxtXHBmSvaX/9x8
WVgHrIh0lhQeKxN6KoLClX7vaAerKFDHOCFpqXZOTStb2foiyLbScg3aLkIJH79LjgwOqqZjXD5Y
bMHMBxWdtSu9VOfaGt73r3xJFJypGa/nuYuz6oQTCc2XawIzvpeySg/8Gbxa3z4o+QBDWxof9mev
SP2Vbs095g5z9lez9cr2GLrKQiSPUQ9cOUP6vn1L3bZToi2vis0xPLlNU0mV3/XWo1MVYCv43Q3+
3r5RUI6yRlsFERPiO0TaBGF+N2F8Un4rGn42KOpflceRX8yhDK7gEOLPUL9ShZoreE+S7eGRD3CY
n2jr88O5DlChVfsHnB2WE+oSqYntv9x1bT+HPJpqhMZmZmAXhSvkuaqWLrKq2GsGZrp8xu9RVKb0
n0JMfgL1OEjwN8xSBHIg/8yjLnlzCNj4ssF/YyHssIfNyQ7GFWmvqsqpJChI3ZaL4TO4r0pbg9b3
/IogiwwjcXNeQIHfG+OO1T/a0t8PPVyVcDG2SrHTp4srNOEhIqQ5Gg7JUBm9uG0ufqqFx1RaRE0e
q/DPD9TAp7wDjjOI1HtwbnmJDB5GbEBQ8WU7OluXeUx43Lj3AuG1FYejleuTnjsON6FhMP/D1uyt
lRCpQJHkd7+l3r05PLoHNYaH56EZ5LUoyDRrSLzcuVMcDPqnXhWCUu3x2/lLgDsOlOALXuv9nole
6wS8cDtwO8dJipGG4TWvSgKFrCnW5/sgTkZ4hl7xpbVO0Fi3sKzhIGEd1hXGEqw3spYzO2PH1I3c
BNMUXjdC3aehnmBCNGP3yUkWzDHFWu0N7fvNal4Uqqm9qOHHDj3PQaWofT+bMDgvNQMDRHAcTqMm
JU9ZgMwDfKM0eCksKuQbM6WIlVXMAFnT3f10rCii0ZLxuZFKLhjrM9vZLwZIkuE2ZlqHV4R7e/tb
HnN4373Z1aKdLbNTmvpzKw32ACNNaEftbp1miYHcsiNngRyFJbux9QmLUyZTqISZ+KgQIBqdCaPv
z5M2xxOAuIgTsE3oPNJGquCi2eAy/NTjfYJNrRRfOBA3cE4WkZCSFZ8AA3cAUkGBRiHhRsfy93B3
Q8mjIseWyDrlBsOcTszcnhp2Iq4awQFzlibGCTel4OFBO5fokkRfkGwDjgW2cD58jW+bcOboqk6m
DiENWCBZNDDycMh05PdDMkgxMz8SblV84ZTvS1xcEUy7ZskZoWAUzWDRzzveFjydyNivpN87b997
mFRPHczdkaWKb97HR0AwEBa1J+eXn2QqbVMpqYRMNBKS6GFKapvOfgBVcESTbw81/2GOZvwKpn7I
Jjis68AQ4fLIdEcHB2RAxdmUK59xZ8NvndFmmFOyWk8Uh4j96kLBzHMsC/eX+WiDcszKNsfXxr7z
OfI7pPiJ8uIQOz4SmT3gSCZiw5IqrTZfVGJtOeU9+cwQfdYBCvpKnppOJyOfi3DfodJjfSj8Q/Us
Re8zIMGRSrw9izLgFSpa7lerJYcqeEwX8uXHVHfRi/i+qBgae4LPqAMXWy5Agy7RTYtM0zWrR/zy
WpZYT0o11nAWMgyuIMnyICFsykyDKUUF+2R5hTtFHUrDagCgnzgWwEn9z6mKMz9AwnMX0p+n0LSF
CLoIZL21b6QLFifLOT5rTtm+wEC6gr4t8FfcYmEn4h5TorMYDJj/rkFKYPnm2ygvtHCmZFfK/cMr
kz78+Jf+s4x4la42HgvKNEU+2WyqckaTjowtIyMY/IwfkUNOIVyipQEsKUdN9XjkeMcmhOsnQbmv
Mo4YLqr96iPFVIb+ROvG0+n5iujvUtEtYLSXY77hNgtgfNqzrheiIL9Gn2MubdTixFdQp7rJBEe9
C42qZkayLu8pgIY94MycMPzuhR9pAZnAbyGiNGZa2Xqj5RZbaQvBKr0d5zya4cgKf9Lwn6AnNqbe
W3GaD74aj+3zJs3hoOTHSP/DX1KfvPlswExm9dNSOz6W7hJ/RzV74OlDqiqblEqi/e9xJILSPsXi
huajvNu63TP4vNqI3x6qtkmYDQmQ9jDemy9bc/pzfd4JHhQmWURSszuKiTerUz6ZnYg6qscbgFOJ
U3MApesGtbNLPWTevSo7r5vMeybbPY9cTf9ZShFs5+suHi/SM+7Ei895IsbiyIN2X6lmPr5WtDXy
6LFsDWG0owyO+gPWy67EcmmFHqS40N0kMVe1gqI3VDy3hCRqv9fJNSYGm/AkW1XIvYOKR/acv8vN
8zi9TdStKRNNs/2/OyCdx9PCjd9LYoAYFuCOj032soWoyR2KydaVNJGUmcnwOlm+x87whES9Sd/R
klPiFq0xnFKhwUq/XPhcoWUa24fBeBZ99gOByHimHatq72slsR9g/V8Spb/aisa5CW/xRlLHhM0X
uzpKAI5azSLvoKtvfRFEtFv9mR7t/TnEgclyZFYQ5XUxPhk/Ktoh5hiVqtThIRbBjPYIlLYwi0YW
ZWPEJQA6w6LxiUM9HPK7Xc5Rb0oitjlellZb6yGlpQTSZmAWCWyETW0QArSMTfACXOV0wJBZ5VOb
jSj6v/OgO7d/Ya6ONqUaRtc+reVIeVZtIlsqb8x2nJJ8tBc48pJp5hTWOWfxsGrhBHyLfH7WuKfx
sPEnVVvngke07kTfl5oBO2vL6AVkh/loowVRxpfkhYDHDCV6wQygYYgRbnh/rILvHn+Ce+IDrCwm
VXJ9JrkDHUanjVgbozF1asae3yPN4tj0dHfNtW8EcgH6L8+FMMoyis49Fdqmp0xPVPrneqWJyjQ6
qn9mO34Lei9K0ur7EYMIVGRWvcSQ9SqvQac2QOu0YpCjxTro6ogjbVoi/aqDNvIHxcEq1tQK8jD3
luYYQZhSGfPE1P5vxm6dcF3DRlJm61vIQ3o+553PQNc+WWwkYBDij7h7gZcRUOKEcWMGVqPtZeOi
YxHWM0XTJrK4QlABUpjkE+BVmjxUTY7rzvMSRCmK+bQXTaajhR/vMSB8Pt4DlQuNLPm1xeXiRfM5
wl2BQSTLrpmU/BUQ7XOx2VSRRKgx+RT0M4YRds5Kp7eIZQp37HLc8PN+Ermbbf4dgdJn8N8bA/Lm
TXmPyT1Lq50oIKxcrEvXDM1JglNvXNHl7cbZKuRfSQr8e/fmN6K1D/FvJ6sZNvR0g1VvXa+qx8aT
uYkCd77DrhwGdtGgvUQ7/r280ixSp21C6zxtQp5z7GaOb9sboSvQvJmtso5v49eJShXCVyGxImUN
cww/rGcSRLRBxUXLlBIoQA1Y4uvkWgDcryTN4x8rLlDn3JZYZ+CH/ZW6DwrUOJ5WrjZOBsKPMgtJ
7R9rl7ObCRXyMH+8L0P3RIrP7Z7UK6W5UAL60bDvUlSQ7PepPjWMkEv9phGb4Qy5P00fHJ+PKe91
GvPBkuOIEXAGeuAI3hjs6IO5KWPZUrNuqSxz+eE4UIpAm64FnrDsTX8NeJXrB0xRyoGjHeL4VAMp
Ye7UdC7ULIkCPWx5MBWmWI4B1rtIoTpRa8LymHFkp3jupnIxllPG0j9eP6k585PvlA+Mf5Xc8ayl
L1DeIOauxI8pjiZqlljZ8J2+SoPxIdgj2uD/J+DkNh7fESukZo/DYJ4i9ikxP1xHGMrkSgs9w+jQ
+ZmskyvWthn/4c8uk74JPO3kZkXv82h+Ox3wY0Yq8+zIfS+ox+fMoz14Vt5TqFRdTXniRrtSWAdV
CojUwRbgAZWO+KGAdNlmeR+iLv90GnkUFpE98qifoAXO+14sY0itPpOfeadnElWj4hbf9vLyxoiR
zTfWHy7JZbBlYF+OCSSmekyI6+65nBJl7RBYODk7cPgVkkU0VumfSLm7F1WTkW9MUvwE1KcTsd0+
QE12HpwFw73Z6rym9wk1qjj/i7Exc3BcjB1ouLIgB96YBjG643BQ6gb8/aBV4GFkzbRn/8a4lYt4
kaLpu7n1+bBRrrZppdOYvkdFhg5vzOa3EL3Ou+3pk87eaaXajucrmTc3jNz6qdpjVUZYwssk2/3g
VmW409sTK3ILeQrfWrwsx1y1NzXxtYXe8YCHTofXndV/OenHeYR0I1VAY8fzBn3BLQFmjgPMwahy
OstlLTC4Qc6LLupp8MogjejVxNNN9IBedB30rnYHqcvpwJlR5h//ZSJi9im5wmpVJFHh2VZimlYM
fBsKlqyrErbNsBXgs4MDh27VbWG6K2wtz6JYcgWBYo5ZPIbtIvXXl84eTmeALsirZCzNlAGLHNJs
iXIHF6L8pfACiwDq0wpT2qW/uX2WKSXktjy0D2UVB5EUu9lIWdC7HPN+hKX95nNcKHzwF9t3aSXz
+LfDb9lJtJxrvF/FRQTxB1NxOo461EebeF/NupWzSZxrSTxfuemvNnlIMVj8M20xq5+qzgmtXLp9
mtipgIhZxhtWyNBlHg4MXnwQd6O1H5fGflBgUahMXTpO/mIrsFccXkZViglX2/FrrJZ9tM1z96S/
65oljzf3jqPnK/CjrI2TAhGtEO5s1xvBMQfMi2TCtneITch90sr8jXcylI9frWdZkcWyTTStsNXs
FpIfxENk2wmfG9GYBdwBFgMSUAbpxyvXsWaBOPpNyzeeUTghm+IxljXxAJQwsWQoDGW3SLD6djYh
HxefkI+0mRO8ddWuld906YjVYPs/jXiUj54W7RGd5q5Bdv8YMOciKQr2vNiiUziCCbhI8dkkbgB+
8MrFSS3cjtlPb7yqXa63y8dfc3vNpw9pl8lU3p19z9pgqSI3bZeMmEZg2JDlI5yfyobqFlNptYVg
ydBJronPULkzJWwwfowrNGVgXHcQ/kWuBF9zDN8ftxOo5hH3/RF+8ecvDQ1Ik1OYojjchrhelGui
bOCH8uhDycGicMulPtusZv1EwVGsOCmZvlLW52r4wMoeYNix9rfgO8OuBN5hC2QcRhbOHUhoEWPF
c6tZKBNZz2VHz//ihvoARzZ2wlb60SYODA4ntF7b2EFi57xfPG8eTldh9VXv7HcasRlh1R8meF+l
lJi4sCXYaBKtPk6ZoxevED5jGckTVDjI5TBazo3Zzdr3ydb1kytkmRg1rVFGOY5jGPp0mpBnBMp2
wSU5XunHZpX9JF7fT6ZKauT9kfg08iu6ZSVA/JqJykcw3kn+klxsVe+pI+dgM3Xsnt00HpgzQbzX
C5R/UmRB1C/s1GsS0zt4UVuETwgHWYtcoTNTHwx/Ia5/RlrSbahuVYCAIbypydmGBWoXr5GV3Hie
3JMeHhZybGuD22YKFWODt8I0n2lgyXtR7fb+hPWETW5JluUEuC8/iLzXlVMg/290pCR9q/cc43CS
ovffdm2FtduNBL8JgLGUKK0eUzg5v1lOy/LXMi7IpRK7CZx/B29/emDPyw+sqUosULTUvV8w6TM7
NAhNCowaUTR262oOL5EKQ0y5pMjQY+vdu4X9uL1P3QfK/M5zSO0B0G/uMtcH4RwHI90fWrDGu8NA
VL2Vk/8SK7Gc74x8rxTJH47MjLJx6q+FSq76Ai4hojit/Wl+s1abIJwtssoC7urRu6uXerxZQFmo
C4W1wBHfYJSWPAqQnhYz7QfzvfJ7mof9iu4fM2srXRvs81hZKJtTMlmy3kQZuQs9HC4YkX1eVQTY
8VkYyESlG9TFSgMUFB7u9sI98L4/9HjZwlfwekklYQ0UEJ/n7HEZ5YPoH11y/wmXNm3EQG+2qxpL
NM6CC49QSJRNF/3gGDKSCWPIdKFb1k67SoP+pSXy5JgsYgoLWiAeCDzu9O/zhpdUPDVK5+AEvQ7A
zC340nn4ylXfvBOai/gQpwOgXvRTlOEmVp0WVwfcTz/CGhZvstCpKsC22BLSolGuhAOLgbSnraqW
tRyq/t5O9eRVJtCYn6HKoz28KvPErPIAirbru65gLhAt6/8ttpIkhXimWai8gvpITIBAgJJdd+w0
V3T77nBqYl5+5SXJ2oWeQk8xlmUODMGK1GIgZYWqLaXto/WrYxXQhM87Hovz2LdPTAE6+S1zjJrV
6OGb83NcHGc/sonXMeT0lCRU0OHehSlydf5PwmiuR4+/H/LnvCxDjsEQl0nVayM+E4SX6rY56Q/6
tSe9hwd50iTq5jRYwo7tcbmis/L9Ze5SmY+tVSVcUFg93wCS7dLeqlcNUvi6yOBJGh3V9MFzc/Hr
P9O4CMUCDWYn/KY0/pPZQd5DMOqOKFOZbmR3O2+X6PIxrpBjdtdKB1qViur59wNu3/LqhLh39upC
Dhh1UJykuyzPu3kZA/ogdOWC5e4ulBhPH6xtEBlC9Lb+5vkkXySx38hv3BndPaRi0HMASx8iNi/x
8tm9cRY5xu0PyQAeh7il0ypbuYyozVvAAVF7ExgMcj9gqc1BBFOrUhs6MWV+wegx8PX8c2cQgHPg
7H1PzErKLhR/a6ZDWngKuFQoCfmAhuw2Qr7NTnzPJcllUs1uUdeX+FHd3M24IMJXD5NEionx7zAA
+i3zrW5wT357iw/2mUYIsfA4VyFQ0oYpi36cdNAKkZXQcchxy9QmBBzI55CIqG+lDC++G3Hjkn5c
pDS7OAwBHESicskJ5qLYM5kojzNHBpyxI5TXyRrmeXrBE9+1NE+6ljgIe2cHnEK6gqoiNS2oCc5z
QJvvTlCHbDZzMaA5cOBauNVxFAJ7rezpXTNzdpH8NEOhwUuve/Eaz2XF273ETi/fTw2EWLPQ6ghr
Zieu1xgdbSL8944f+Tyj0J2FNlaJwAo1GFfyErnfrDV8BL9QF4sigbx5ImC4/x+4wO2brSZvbu2q
cX7TR2fep57RlHrj3Zs0jtV5Ce7clSTgaIi5zag13aNjZ3VwqZkLOuyUMnWEDTdJfivVdKwAN4TM
Gw==
`protect end_protected

