

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LQ2vJKYKktoZrCpK4juRqJANqbtQy3/ocOY3ZqWcaeltVJ85vibXAMA5tlVvS0pp5GAf58wutyGk
pEVV5Zv68g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oMuoQxHU8xamO4YIRqVhC5y86VVKXTIB4hGEIvLUCrdkutaN+fgAx1w1DFW4AV5UF4/dcrqjOzkY
K71n5sVp1APv9EcDNy4SK12rfM6JNEmec1W0js2v54algVfB410d4rZG0ryxf2jOEEtG3y1R1uZT
docKTvmf8ciwTam2vyk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RwKTb0xAeUUC/Zlh40ZbRUmoUjB02ejSjmyrw31uw3LFcwmpLfrEGeQFx9W8nBY5yWIBOz4idUaq
fc3pMxhJHFC7jCdnh3Y8hC14pp9rspO1hZLfCOxHKu7GOhZZlRDfFJE9YTYvNMQlQ719mBEfy5DV
yB6StZ3JnfaWR9muuKfjZivHmkGfCe6IBabrX2L7+LYnKKp4Bj89EkuYxLdjSsxwwHL5yBSzQWsD
f3NymUlojWqzg7COUuAovEX4Cr2S0yo+Zr9C4jJ43pknI50nQ+b7CaiUKqbCSj+K5CzuK/dZ/FYE
aO9kMeHqHP3vuIYIBhuz7gnYm8SB2OlUmalvFg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yN6ERKfUqtxcEaZPhTWcKmh6+v/ubkhs44a1yogYIxw8eK2NURIBs5ApjPyj6y69SFt7ufKFYnlE
zs+yxTyZOIDjE0iu1eOyuLmYVN1yfs8OFxlynJLngPXQyLVxs9254patixjWMGwWk4PkkE6mKJuY
ZOkdptcpF67u2/mYpXY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t5IcFW6UoqOUfYz1GOxoQECi+9Dv8vBS33YPIONcGWTXCbnB+Rky6dyYF4Y8M27ZqAdkRtAsKEP1
XbHsYeeN9tcVjnhsAEW+ZxZyVmGkxa8lAjUHEo6bSWwd4akFKgw3xIpbktgKgaV0fLwj4wfHvTcJ
XEKHWYqSYc/CYMdUUlUPXn3ng5DzustWIyUHmy7pVesXYKHPGiFba8n7HX/7Kf+2y3k3y0XUfQRM
e1vWugHsLB14SmtA740nmVJ5TRRb/gYA8FobWc86Rp4qtvRHvVvYBe1XopHUWeY1WEaPGutqYtgU
FjBA3NC9aJ03W8dZxVcVFZhyW8E1aSZwJp996w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1517888)
`protect data_block
ChTtjPu//dibE7Xb5Ro/YbULlAfORZqyTk5Z6kfhGSFTLaZn4K3X01rDv3WmyAXtM5k3Psr0ZTIV
WJdFVRaZSnj4fjQP9/J8dAJgwvf5Euu3alCd0D6CGZkepxg0uAKj6Foj/F6bopldTxMVfB9BUipr
5ijUBKBIB5cjzucNPrs3wQzKHywZ1AslKVZCLRY7blgCezTiQoWtCo8K43G5cVNzN4aUIiiAo1v3
TQwOzvfGJalb8mktfLWvxxH2ijthgrKPY3Ej9F1OL2olEfVuYbR85kjgabrLaRtG79X7xlJfZgoF
84/l1i7Lwn5w5oF6aS9Vvi2ECPlC+RFpOHvRynAIknJo9GZ2aqarhFcTTVPDxZQ/JCWCzh7+pro7
0plnuvCFVb7QDH5Uhh+IvTL8NKysArpZdRX59J6CrtYwAGjW4QBRXZFM2h6rA63xwm1+FkKtECL2
ZmW5DZwO7iDuC3FukoImyQerQFTNXq0zspEaa6/lA1i6smJp7xvxSxPrA94wOVyP9cawemLoPAAd
t0lDjnSogmrUdXMFOQ4wFXu8Pji5mhTQl6hPQ6AovuNl3mK/08KdLHfM/WjziXTx5fhVkKjFZCeL
WAMMwxUldn3Ov4NVDBG6tLCEPRSmAAI6XmrJ50uuYEUfQ0JFVK8f8wnF8BmrAJvv6veUizLLBDl7
jTTA+FZ92DzqRlIxrRJRvFNcKnolhM1CIEdyJPW3P5KumGfup9vQVGfu6Viq2ZUGxpFR/n/De2Du
YoRYVwS1+yjukrGm9Vu77gLnUxynYi+KG1bN39BRDAKGkB3ghSwbzMq8etBzSEI7IzZTpAnx32em
jRKXMLw+rYTxog/BOc+9OqPqKBPUbHyc5rIMIlk2jA1GU9OTYrMP/k3HFGzujq+X0WNgbm/9pUhL
5UrfWXh0VFUoQ4QsX3U+2SqOmgq9NPuS5HyraT6eFz7sZq9+IQmCnb0RJAPpQOxU83oylyzZ4UPk
vBCwigVTmJoGAru7C/lJEoCmAxYKkT47G67hFFdJ+j95pXDBetlIPkWIJ8UrUn1G94gHxHzKQWWk
UT4EzPr7/BdgH+j1I/m8arlT13Xg0z1Qi+5SKEzCwVvi2GpHdDn5hpfiXKf8qAWlrd1ONJxN/Z6I
19NsZYoNrzMlSwhf9sPd+WIGzBVguPfwcjt6lfgLbzziN3M5LSXEYLeJQPuWk++esBEY7laTUrwX
iSOYHqhU8EQcVsuokpNOjdbzku7iQwCubHyWwQGunn68hERuQDWzfdwSS0+Wn5s94KR9ocilSWb2
dJ9URnULH43B4ESUmpG80gYSqLKrxDBfEQAbQNdrxOm7Fe6H4Gr9/GLbcFriG8CkxbtH2mBLmvYp
WTWnRXk8kPvMuqpPaHz7JJhDGibk4znKmbIQGvwnobnpus7TT0qFHP1OV8cw411n9u+iWGAVtGu/
UbliRmpUztilcy22q//jbuirsAyXs2KPJvBEP9YM17lrgHt2Zpxzyv3Cf2LgpEQ8wFlwhiX7yAnJ
JwHhs9xClNmd/VyNfsALg04xTPVNRBA7mSS2VvT+O2UQMMGkDNOtf21aPTOH37phHn8BniEBjK6o
VIkNj373emkoLsH2mVqTHxpnl48J6rEZ/K5x+G4yxYFoQkN1FVxSbHARoQHs3ZaaXBgpWazdZHVt
CrJydiOGH8U44jzj7I33Agxkr63VEikut3anz6CGSU1ehInFCeTEkcl6yhTAKjBnX14S9ctQ51lI
oLe5k5GRgjZGDonlauIfym9zUGymAyCGCJGZ7r31hoEUu/Xgz/n1H/n5e70j+kfz4VA6RS4UDoYp
3yHGjDYqHwAgFpk1GYPLX2xR8wfVV0XFo6jpWkscmlmjb9S5pKumrLjh/wCIBD1Q3kLzrlAe4+Dr
0KiJ5dc985cf6pNXGhNV6j6nu8yhZOAUL9IXg9mrLTISCtODfe+2a6cGSZCEw2+XRVGtU+lehQ2L
7jwOyoCrj1P8jVN8iYvBUdyy0yQvpSXAMKbgwR/Z7JckqSWa78rpFBNCUnFgLd3kq3MfdbL+KcWN
CNFrPDK80KtQNpg0wlEWReAGX/TVf2OQVjrTFulO0dgHbk6b9flAXgjJlbXhbMgONE2PhyZ1hqAj
dbzfBVkdSY+04Ep29dXk/R//SID1t0H1sij8tUP5NC6i9bhkRSrodsaR8dQrRiaJsuGVZQeAoeNC
rOiKPfe6tz/QI6sIDZ9RfuJoZYlBz9GMcIx0P/1186Uk2d5s11ODdJ1AObCGAov1rFJFf81zgCa+
asqKaV1DclugGW0cRezzmmkVbFEUYDTUDM4br5mxi+jYCbCMdGjyThwj14maCRt/rsrmPeOqe4iq
swYALDlvXUCzu7GpmU6Xxelccq2OMDtqMU3EGKCF+mMPIenZ4i53KeM/iXYCWCQQtYCl2ljhAd1G
TbRobOHpM3EigPTFTVNZ5XB3mBshPKs3lSI3abnX72nnGftDQWu7+RmQQL6Ev2zYB8nAy1oQydrX
73Hr0tbalO3jSbEeB5Z6qC76FL2wTli5wDzIkmVh1jsvICODQxcL24R0lZ715/nOjfGSZZCZsd49
wxvEGtNoo3XRgBSjO9bIB/rbc6jIIjlnCvuewjb0nV+SFb6iCLluQu4VYQPMJCC4oNkwjL3wcsxI
A3sFkNifZsOodbAkHuz1LIvc2rlOkKTTxgjuv/9npY7Tlso63gUJolm1sPu7zFPbJiSSXKR0Rplg
Z1N4fW8hCQSb3iTwtkqV4WhLBeLop0hr30U4FhzOI82WiXG2bO+WD8xrZDvqRzJpVRZPv66U45v0
6COgTdXk6ZilgteXB8sTnvWBcZwGWJgmfAijOnFjiN7yqeKgOCMCrP2WI5rVLGsgBrZxhXAe55r7
WWMevaoDcF7HmeqcnztXUtA0BbLRHY6AbKNubkZUoPGmus5W7Gl+azp1ECbFTY74Dg1DuFtgDcJS
yD5aE7gm5WRzFquYamLZGw1oUXNcCcL5021k0MoGQYwcB/6RYav14Ebse/6eBv3ykYxOXByNlQ7L
b72+8OWtrDC+ZiX0Vxm5ZIrEDztpECcChYCnXokQG06zGv++qcl8IkJ5DIF8NlzhyJUAshEaxRAH
dQGRThVvsczYLg3vCUnq5gHJOk2YOec/PWZzeHxmvWX0EpVjsje8jsqcQR9b3K9uPeJ28+HJ+z5O
aLxAvJMQrcUhzL5rWoMyW39V/G5Lsg6sF2g6HeEcB2NAmBZZnvrSsF3oq/FioMqj2KFfw2/i/+hc
7dKwcFRk8gs68o+cpiLor0bncn6HeM08Kbjx4Czeqnq+3WpyZmWUTvR3itTkgv81a2YRugwAhK86
L9S04/aJURDGUDpusIMEumbZj+oVsoP5U9qKbhK1NYn1JS3h7kIuXDZQ37mQoN5mCPTJj+Fkr+73
vqcZVe9OwecH/l+dwL5EmA6jewm7+kJdwUu3Bu0mSphiSQIk4aC7l62nxEBSf+Kk+IMgCs5KmO/l
49MQDpqM+00R6iTWgWdo9fqX5PkH+2BfkIkhxps2kLgb+gJ5GmVlfU++27Nu/9wMYNXLqML0OULz
4VjDIWN40GTEWExjedgsbVSNEdeIz+tpzC3kFWXENRmlkDnfgiYUFMaHHGDZjgFES+tH+smbkJzj
ymUEOIaEfhO1VBZDsPa8eRWa8XghVCxFPicj1l7gmg6Q12UJC0XOm4hUczrjHkJKCI+Nv4iU3tgC
My042vF4h1wRM63TzLUPfnWUTSQtDnexILXvYbGKN2BDilc3VVvrXuEjp/+ezc11GRUwU0W6Cf9X
KM/gXHa1KFaMn4HYoZGQvV19MK/ne9Y8YVyuZIDvYrTvA97Lbq5mhWlq30Fll3OZwfRKF2BGenBw
RkrFfkO+U7KDdxncF+DICAawrx7ZOEhr7zOZj5iDRlAinG2GHraUHu5TTbhD8tDfqRayG5A5QB6s
JIYtgCOYANaC57yGvHtqOf67kH8sPJJa3wziJj13Lw24xE1sEyikPffkpCFpVsw7lWVIeVLBT1R7
9LaLZ46GapJwTq0cgdt77iWgc/N4DAkVuPK7SmOe4FgRzOKafBmHbgYTei3T6Z5wfrMMqZIc6/ac
VI1q4i8oTFGeUOtySPDQaGqk6s+4zOp9/5YG3SG8fJaUvHXrMqYqIjBTn6J9eSiM7kx+HWDphbWM
9qP9F/gAqJEY9Yz8gomhvEeAgWMcEqFGR2iSUwg2DftQyi4pLzhgvSY29MBYL7DKIi8Mr1MUai2Q
tLf52//EgQ8lunoz4JkN+vfHcN/fiACs/ErrtBeYi2Koc/vFJyR2TikQl6Uj65B3Cdp1RY0F4D81
wXzQjj9YP4SMIIvFOITsU1hn5ngeyDWvZP3Eu6sjDOUTQce321FehCTYg6BpzUkPpn2JC+DxxkY4
Ss/G3Ay2fh+WDADO6sVGR799QzefIuVgZQ10/Tswugj8eklSkb27AkLMBh5wcb34+ivkkHp6gevi
o88//Ukz3PTeEAYwr2fpNLAFQednqNkoMHmSxNdq1w35Lzj8i+DHqkatGWnTspAd02exDoNe9ISI
52VbmaO9zEcp0jnelrHIW3k/LLt1bv4dU2HuuShPgNZ7LcmXhD7fLsO77RTb5cP4Pl8enGC5gC4R
6+wxzhzIvadg6uhhqpcCzkolkrO5ercGGSFqRS/J77O8GsYL9YaxVPpmW0bUPOJsJsAWqyvoZDw0
C2GJ13vU07QcSjlXgkdSP942pMgFaTuA9/ncRVwAMKptbzFobeKC+A9O1xt3DqvNXlsWqw4/N1GA
XwGKX5u5cAGgcR0BxhAR3Y5l5lUMd7S4CI7/SCb7latf0P5tnJa0oMtXBEVHov2Avh/UJvNT9E5F
qj5V+RQJ7NrDzwtduOgc9WYoJ2UpIdhcJuHkH9qqi2JObLeyr5i/ueHIynTLY8iVJwmNcceskiO/
GENkw6RCpxrU4UyLRAbWQBIrhL0zkAJrvsAm9ygAnHdHz+Qwvze3iY4ZdoUVTsqZ7PJTtseqwELn
/9Fcm+fjzZkI+jLdD3xcntPRaEgsXLWF/L+WTgeW0Jmc9uzzf4g2FSKgIyuZC5CJeh0botj6Momi
ilAKuOamy7sX0BhIzTQ25o4o/7qbbcpsbAvxMhPl3rVWeLMq/yDqzZeMFfRozQVxESlj3WU6dXin
L6ySQBAyEn0gFNo7Hln4J6DUZ8EtaWZh+J7JDsDFtyHxspcXQJkcFDCBh0MKRrFPWEAjLjOHXdnD
gxmMMjkE27x3non19ouekveFkSXaSFtPEkEI+i9k3ICer8F5iAMWp3wBd7gm4Mzaq4kiGZhBm3Me
mOlOluUf36QXNEX1LJKfnLJZxCJQoUghnLMbuCGU1GWqMd+l1kvkKHjYQpB6Yi+nI3+pNZ6aNbp3
F4zQlzYRV07Mbyr4fwCfULXxc1HAKFQlfaflC8m5jPbrtf61QU97kYGuw2MjqMsnx2edaLs0+tMv
w4dOyc++nNmHx2RBc0g1MCSSZTosyCqzLvT2k8oxEBTfM+kHJFWN9ARe1Mkk5M1VofzllTZB+1pR
ThjwAcjp0eDG6fjF+06f2SHIxF+PSwWpGKiUsEKAi+ytkZY7ApYZ2bq7zO7jIgpuWGPGTRNroeyu
sCxkZPUWHeRlqwC3j4FF0Xw+Cqd9GJqxOpaTQazSLx463a430/vbEfl6MnOp/frnY8CKPx0r1gfH
+uHHBsuZ0N/91t/86AJAMdxvrAvTH5W5avzV2vcOgj90mMBiyn3f0aOGD8yrSLWBuj8MTw/tyKAR
3Q2VkGq6KiMEADjvWeSfBPaYioZiHudkraBbiefUbuTCKetzPSC5K0AsiXjcvwlWJe4lRV8TeOTJ
R4cGC2qyjJY4DHJMFSqpLKbTPmzZ/syjepNWXOEyPrah0725a+JDgOdltEreXYLfutddjs3k/0f4
WsxrZN/N1PCO19w/sVwVgCIxYBtZfLypOjUrjEQXXY3gwFoOcpjYf21NR/Mq32+MRMiMS+YAPUTf
K7GzZQxlbDxMFy8tU9Kfi5HksHj0+1eRF7+lrJwSV7UsSUL59i/Ey8As1UF0qh7DCSJvUB+gwhe3
qhhardnV7pAU63Y9TJiWrwDFjlFskRdxTG8Rx4N28aHastuP3eT26syO5H+d9ScEFho+T8wPy5my
fl7RnRrYfTKCFJLXlru78EaMR1GCYpDWGKdavDTEvuOvgtb1/bKQfc4iNXGoSca5iJVj8U9rP+qY
P9H16uZRopMx5URungtKBUR9Wy9cd3n8HbsLbFjhfz5g/aMJ2BqJBGN4y7RTmFad7B7LRG0n02oy
CByzrBbnslLi9+xtu+zTO37vHx+1MZqn0TMz3W5a+6E3vnVHYvVcDe68aUWH6GvK2uG8bkcOjYWR
I1SGi0K/bFxoc+zMmkPluwD9focD/6ZI1g6Vqi7mMmUAAX5sdTePGOxkpa1vqKZgWIbcKhgyeRz3
4IT3XZ3hDqNZY/vEHzanhfLQgCD/bqL/DjCGBPjkCyC+lgbIyssJeOlsRmDkBPaFnvtbgX6LGgqt
HyWPt/iu0XddzNsY7OaAh06SGlGD04yyZEaviWqjjhM0Kof5LvpFhQ53PVFvxWvlGfPa6B6hFOGQ
dD//osqtUrMoGg2a5WwEdnF6gL1ZYtDHWfnpxEhoCji1N8aJBQLAUt1DGCehKOjlJ/uCtzpoJ0Yt
DIOS24BOwx8AfLlaRmmvt+wdDI/mflSPAMycVciL4L9YEzA2+LZINR8wpakCP3Jbq2+CFsJbdOvd
8hcnwKpeeRXWwt8cIJyrfn1ekoRyo12QJrhyJQ8uuk74Go40k4mii4RWgkArUcZYLlhum0A3udzL
nCm5P/re7gNJ9EdS4lSPYtnFzD63ZZ3tY7ghbuSmT48PChlRaUhEvAR09euZlyzuYYxHvJxJyfG2
Z7gcVCs2ZGtZIGuqRBB81XmQsl/ID7QjQYol0Xd1xtky8sf8De1A2EXOGYtKIOWPC8YRS1b4d76X
51AVrnLUMHYwn67ry0z7ybvmvGIMhbb1ojDUBzsqwdzIWOBS/VNLxQGvN2clEtcWSs35qgwygPUS
CXbJOsfXNDwuw/ExKqe/XxlNdK7vxZ1R1Ssi/xv4oIvwsOjs6tq8ntgYueIUWwIo8jyBV4dh0mu3
+lwtQVZwN3y3O7mRDgG523mSVFRNMD7MPPSG2Z+oXUEJNjn2i3cJS6ZiPaYqDDoTVosFir5L1008
SE6UR8JZbrTLmA6iKNluhl2UfZ/J7DVget263r8/fSkm8VrOyqg1yL/frE/3U1sTVkAFtjUxc+oK
oaL5eSAUSbm3M58EMpY7/0uFMKlQ97/TQtjWaRvqVUcg80SBDZbvQkhYxucgpwhfgZVoRQxJ6PYa
5GoBHhUPBpn5Pa7hWJV2rH3+/1cSXs1fNTp+PBkxxGBrhUqWDEqHK41qisQnuPyXxLwHweg0K/i3
bfF+xRsbj6Fwh8vymrTcDYqKOz87+HQGocXRcQNOR/oFX1G4pR/yWXwYCDHmRn+uDbR8FAoymaBE
P0jj8eAPXDBIQQ2jKeucpggzHh5xdDN1db+LBd7p1R1NqUF+CXpUZlgVHbQmYShhln0Yi52iLSVD
QL5I36gpmGZi9aAmaD7783VjN8oREDSCwHX2HS6zA1i+fp1l/tXtTQ0wKgTvhZkYseGRtQglIToi
cyl9bjLBCjKjeRxMG8yBQGSEHxET/oFjDn0mWf9Uzftz230VpeDY2RFXfq9tY6gtfviOIU7lYel1
VBz2rmd4VCn0GLIfSMC6vo072S86xSOXssH1whlxHPCgjzM9BcKkNFxXszYfVk6FTI0xNkha5kek
ziG500LUXWFoj685JbwCCpk+FSX8Yv04fR6UCfH/v/X7QtBBqRk6xGMAPlFjuUSk+Exxukx3tnrP
yJxYQ2mqBq1IAi0pheiUuly2xVGCgolRWU2zPaTfh6qMe5Ckbe5kEu5WTJQCv2KZFZA/V41GvO/I
bSkR9tpC2LskvPUy7byRaTHMxBI+23X7ZA460jMDuYI4zRXE+nYV3vC/pUWGGsF3ZnCw/zMDR2nk
esGBwvUpYmbtftnFtRUq+QhyPvTz1Y7wBdGHv5AowTlzC1YSafzJCVabjJulUCSjNnjZai1wlnVU
jAipamadLG5d/MRk1le+9YkRY1BQc8P7j5kYAheWFhdSVmpKyYJFSlKkkr/8oY6SV7Pcszmqs89+
HJapk0V2m7Wb3cot+4Sj6LfkpHE0AUxk9JTIoTnbIS2Onpkjh3phba5sx4co642IGYlogCzuXO7g
IO4ZTlNxUnQ3tyvec/+vjDxHdxxr5KdNkNjUEqY5FIwfQBxRB+bMuJexbbdOmuVw6EMLzZZTR1Bw
djbr5lwd8OrpDfXBToTEPFcEPq4LtT7aTAC/vC2hSdAdJN84jLRVvH+uvUtaOMotMhtAFLSPyCFP
+kGYBUOpML3G7J997y25iYZYgQ/LnSU72Is17uyIqoZXiQEpWRqraKOJImuHClTcrkTuYFZxOWi5
y/V7+Kf/efFebC+78m+daaRzNsz4C7X0rUkWe4FkL1ik0UBii1wNKJmId8IskSwkSXxm9loyDCGj
YTAKCTX+z2yUfmoxrWqNVzSMJ97KWKJP+HIMMknIPbhZaPgGer7xPMbwr0dYZJD/rbMwnhSjRY0J
eplmXULKzM9cCOhIkRK+p1VJtDge3WjEF9dsdzd0qqK1R+ffANk22I5kc0m9tu/aPjjr3EIAc5Ie
9VE6e/0eQI9K+D2TuQJJKFji76LjA3XsJJYbOKXaT5R2tnlRKWHS4k/FztTr1YPeO3XAIVWnW5TG
ZHr6cAjEAVIJo5TWHeOx6jRZ80JFlwNsKkU/+U2rU8+Wf9cgXRo323Yqb1PA5JKRjgM7S9YiUrVz
qrPJpwKNTmrf0sZRfb1zOMNc71xk+wjbVkz8H4VZOiVVw0DNBOFfnJfZVEW0A2DVrexn5aN0gXRs
z8fFQsNxoYe22ADcjQ+JNA2s2nuYyPAW6xrmoit6LTn02NdLvxMtuN7OvjV9OfFA2RaBv3uIlloU
PsMZ2emRNskhO9jCKIUb9XdIEZbf/kymP6viLB1Tz1enS1Js1dvJBbdyp2ZTEyWgkBtCCehN3fGP
u2zME+Pildn+Opcc4zlmCkdR7uhUs4enIlo7cRi/Cwd37jiQ9hABgA6gpLzyLQWcO/L0XaHVIpBo
8R4a8sjhKt2FbxVUxHx4JMVls32fMTfquas0xd/nwaPP3NxZzEet5nHkTUBfXZkBb0Mevl9jc1AQ
U9Cu+JxrTrXfqLAMQ8RsWvo9eRfF/iQmXJ7Fm8oLDGT/ViA8WWW0Uqv4I4z9lNuNZoPiVvDc0HFL
ad95eiTxlrqreJQx+AcdbvI1pZ/V0dAzZdbpDaf/Dpov/dL5HTfTVHtffaET98lqFneh+TpLR17o
nbof7UKekO+p3zUkpToWuXNLikB/kCqwStwu3W6EfNMtpBvLDqY/OkaR4JvtscPr6teHwTpldnCC
4Sh4OI/MYswPlvZKJO2QZw2AXhAAfIUUpVJfHx2l7VDlb4IgcriEaaEONk/BX23y2j61uF4LH1fM
FtO3sbjeTQlSDT90csENsO7F9Be5aZWxOkoZPKD/mOuwfvNia35PWaq7yLmtBtQCM7XK4f8k2KB5
BJl96D7hpL2jVxzjcm1rcO1ObEKpeAXpjYgAak+JdRHc860HPdc4CTyFI+Q/W9GQuUS2MvvCh7j5
xjX3AFFMtgijcSHIUr9+1ib++a4Tz9Wzb9WT42PvHH22hEnG7J4P8UW6y9XhTLTYXctbJqk5EDcD
xuI+sjKoTfTX1nPxqSsAyZu35bOeilmzFkJ+kHdoJz1I486YhC2gXktkSOfKlcEPmuOomU/j+wVD
ShgN5Bj7vp1VX5v7p+FeC4qzRdHwM/UPR8AIu3N9oVKSMKpO06zeej3a/W4wAGFu/jl0AsDJK0/+
L85tXvSaFi/drzNjbHyIPPxQ0+mq+tASto8HfNp9Rql1pakVF/5EBSVB2pWMNprZLnx1XDQMe7d9
q3FR5LJEVvaYghdlwGr3dTRC3DDHIMc9Ulgf4SQZ3/ApYEyHjfhbniRIuRbKFpOwn5PcEzFrN+l1
QIV0px53Ku+M4nmjFhqhxIZSoqk5N6zj5td2SQU3LPD5fRPyXebnzSJCuQL3GYDcicPPZLPbu8P0
5mu9Y7/Te5MnQ5hLpAJSPq0feukeEvskYQitl46fukEhDmyolDN36vR25hFvnPFXbOIGzJ6/0bR0
ikIOOxtLCLba6M9FUziQxB4m9p+cL/mRrvReal8hs7XuSTy68rmr9/jX6lxFTxYUN/CAAG6fJzN5
JLWfM/sDa3IXzGlIImp7QelNdXc/u7GQ9pLGTpikL9Z5S1loUVdTb+n4fTl9S3cq0YopPKKQEi/7
zk15xFPBPdbuWZ1Xn/9aycvMMGuzCp596eX1yTgObyljb98bPdeHFbtCDoAZrNh8ynvkQl3aJ4ks
t3oOSo5lCpYWeMjSLPM+SXtaQhOR85l2XkZskGJyhfNSBf4b1iKlrQSoeWZenHXQaxNNdIxZDLDY
a6o/mzPYuvYZjTQ4ri5/OBBbXuF6rQM9pJWPXcxqM5oGfwWHbwHtcYu7D0yF7jnpzh7bJ4TErOzO
4HS9t7kcbhG/4sM9YMcvvTCU6gklabgEArECQDtW6w+pSIIYTWmH4YY3zgsbqm3UmvJADtHIo5+v
YouZ+zkvgqCo4K8d/ek2nt/c7eFvXHAu6Eg7VGGVuefBzrz18SeXbKURlzzEF1LMjelqe2GvQ1Iq
NYY8zy0Uq3RVMk6LanilI3yv3esBcYz7z//11fwpxJ2z5HHkL6W8+BsMWwp+75uN0R6ZDHQz6nYx
m9bn+JATOfkN/Kh9COA7Fxuo5+eFt97CDCEvHmx4FtDrx5vk+cPPkVVyyVyUS+0+har8IIC+/u5E
u7uZOWnEiNlT5rGQbUjt7GEOMcks2wH1QxTvY0LKyzs6NkFDi/wWLr1H5nDagGEWrSg6pLRu04P2
34GgrunnL6TC4yTL7LcOpfDZrcWm8v288k6bBiy4Xm9lhePN9ZX79rKl4Umwg+cTQyG+JA7fPMiD
KAGOEBsfChwhoB5VYKGvN88gSbISCKeAguzjJcEjQAS/eiCG6toksnJ4jWYtjigL7b9U/aYwlJyW
pdZEHsBQuKfEkYgX5Oju7HYab9bdHPr4inhDWKoT3/hvoxSGFm8+Pt6mcbdyYo9Crpohg6Ta0gYU
vifeHawTN8jLGgLatQxhL4pEM8KDVq5P0UkRgRk6FnmVi+WFWUIt39Zg2q8cl9WV7l6tyIUNG6zy
q6yUOkzDbjORZfNKSU1szs9kMvjMBlBkg4esfYjgPL5nIAZF/7M6OakXAHIlM2+0y+BXKRlhYC+V
FT/KqTeNq19XzKp4BuGtE5xIPCXlH/RrGOArVFfusDfGAv/bSJ18KY/cYIrEeaU0VUzhE6iP67d1
+y+DDcGJ+phZBidrL1s8CmHQNNG3b76AA9SMjK91J6dilmlhME6a/zHAoJ0YuP/7BLdFLKSbnTTu
5g2BRhL8bpEjhbsxby9bxDRkkRyZnPdVelavnyN0k28w3JkFhrogWfLRQxgXD1tuzBuNpn64QH7k
V8AXjmMQKCZfOd235qzROVS29ZNCTmILE9VYR8DvFpvVL4PYHkxH+CdPzVwO56mGwc2LmOY4+F+U
3haWSOtaI8dm0z1tpp9UlCF/ZFQ18LMBfJwviLBkNr4OPBFVmi4HCseMxERi3xyp2yvHKHj0/WIQ
OVjKqJgDQGlz9zuwULOpKlTlfKRI28zM3rfgh5uosDDrDz2FPMdfFfBDbXZ3UOWHlgOQFOZOLfDH
2RLZ9j2mCeWvh6/1zCmEE5dXSgZ6MmxssGNDX/rYJed3iaA7Nr2VjANRzctnvMiluM2AtuOf9XvO
Lt0/UDl6x0mbQXEB5mVlsS3sG2zxvwmDesSqExbnYooElaMJYcEX8DGxqwH/WARaW4WdDneqaS8O
NjIT8ICWPzUCI3lmtUNROQMO7jb096vgAK0xeSnM6Cud7QwBKWoMh8lRdE7TDku5QGnYvnB1KsPS
PK+0rMVs8+nNjBhMsZTvHRFLdXAjhZ0xXW/FCJJA8KMW5rf8cH4aZvpls2Az1gg9GOFXISHpwSI3
zmDY4yp8o1jwBb0rnuLtJ9a0fpYCmr8w38CHkiV2bunK4wM11JaVe5hUJeDh9mJZPe9cMUTIRG6J
XZQHs6A6S0OxguiJvbt/xJlR2zwhwY+hJNoR+ksqaFY2RMsFSXUxNB7OIaNIUkomC9on7Nia+JBd
aUOJBbazN2pKJw40gh+uGwSVG5fgM8PzUxtFdK6byMJxau2P6nwzRtAUUV+tgDPymYQYk01+NcBW
h/9gPUGWjO8ceFqd6h98ifkdLBNQb70g8qtzN0+Iy/vjFkDHnKqpaZVBBMpCL78SW0EIT4jD8lt7
vZbmzfWkqYlaGTKCeLDizN8Ewpzt0lrTSiB1Cw+r7/EBl6TGjGZ4Hp/HYVZ5EoX4e2RPzDEFwpIg
jp/CY/+WiTAKEhIaf2AfDzRVsfY3Yhfx/Kt/sxwUtsjG1rKcdRNUzvfY2TQXaqXudNlVK6zBp+l2
Sw84CG6jwhEbPbPxw5jAIHndIY/0+iBtTdCCiLuFw2XhyOPz24gQ8mKyuSQg3OekhSpe1i7232bQ
e7E2gm5bt9GW0SOv7oF0lsrEsBnopaVlWeVbcIbVIof5fundqMlgSw7xgDAGoMlZz22DFqThiZx4
NEl5Sq3mJjqjGn10eEw2xK/sw5ZVewYYm5mSnjtJmaEvgIWe4sIheulC/cCW1rOMfrnnTCTFQpYu
MUkTOoks7z1EwHu1O2oeHLBXyyZzN+n2BxVojYAuNyOOig37mLOEziCq3CyWyoOVCPry2YAPPHCm
thlgmAYUrs3J/fKp/NRH/haGxKcqaBimjrrcq7VDJ7uYi/MTIKPYg0mgt7kH8R7Xu9QG3G0fQHH5
8S8t7ZPeDLLEEHzAIsJhis7evdhEFsR+e0FWAGu6GqDly5dvih952bqcJl66tx/EirXiU8id6kRL
kzD1gtNXW9xbPRvAsD6RGo8rSwqfIsEMD95OyKkCkEfUnliP6s/0LvbIfzWc/KYoj+pBo/LwvEoK
t3w7H1LqDXkVt9YfTtoZlZyosyW3lGGncAR2XpeApoAKykiYUN1PUjnDlRUC9HBQtNbwA1IlQ7mB
jlHc/vo9pcA1MUgKf8OVPwVQ56gNNnhK5b1PtY9K0eHMNRLTBuQ/ghvHAJ/pN/Hy6o9i+EjUeTdd
rmsDLG+Mb76ipWWeCIAorCFWEcWZS1lCQUF/Aersyvbj8DaonhHd2fbh9Z3rbUuZcPdVKCZGMCiq
/A39W/aCHT2jcj00o5PpqmhpL6yPQTidHf8SO3gN9iEjx8h7Y5agFCMRZs9+7J/tQ3sIJHfCQobd
m2oGrqfaR2XZtQwhk2yyuh/KR2rBvEYXC9m0HsE5P6E/0M6Qp1XsK3mu0NxdNhXsMNXEuIJqdYfT
nZFKjU9B24nU01iXtgCvNcmfQmdtMb0fdNm8tz+XYnqIunYClFpipQtG/Qp8ZamnB2kN4mU+VXov
ajtosSFRPSmI/xqF3e63oYNrMIkqf0OexK9fsKHLd68d5rAmi3dmabIxw1ZUcy7R+DWMMprWvU96
F5d5P5yKldM9Ls+2PcUbTfBaTInTv6WiIMnJHChZr/9vO2kQIWSusewH1cogyMdjtcNMjT54Yin1
aGJYnaakTDpiIiUVKUypm7XxODlGNwqpEte9T97hjuksG++TfJGKpb59JxSyqEOqivjSZGoGZXyG
M2uziYzc98PCS0KQDiqkIlwOaslxyLQeGB+dTituJkyYOPZviipGcd48r3JDu5hTr/kUlTNZalqe
szcKNL6NB78mjVFcxrdo9Dk5TuWS0uslnH7ViqVcY4rkgoSmmHR/BGEkDsc3SpkLcyPFRRHEylHx
folvtcCaM5pXjl9Z5T61hrBJCwT6KmqTDgIwYh/O2o+kjxyw4san0q1l6cH+L9e2VJU04h5+0ssw
isEcrxywyJl4UEkM2Fb7Mwn4tjgZXKP6lV5KxRv00ri80g2f53JgNhQQwDsW91paJDr30UfKhFe7
TEP0C10/3bP2xD/Oyos0Ru5zMJQx/Z/CyH9vHgN9XBQbzm+cB5Hy4uKIBz0UTjrVAsCOqTsvgMc0
p6TQGt5uCoaW/pXXvZGA6QplX9qFwOsu5Mwczl/PSeqp3+/Hq6LJ4jTo+LEVTA5LXHCimVzsFw1u
moKKuQEwh8YTgic4iY8gE6tzLTh5t1xCeExSQcZRqd1eHaeH6NNgJfkybkn/TjeezwQSz9yZBUr9
zgDStIztaDPFnHB+0yjQVTZ/hevsMBfRnVxGRt/Ex83dIRUhrzux/TNUPdZzQ+3mzquqafU8OIv5
YmzWzFTpU7Z8jgwhjF3NhOA0HbU/IWB+no4cjxtP6K4jg7TYrqAMfBcwhneLj0rfjC472DVL7Z3R
tsz+w27ONyNuji84QPgQc+W0M8SOOA3KlbOZDiu7N3KaTSHFGxQI8WCdq5D6JxLxnmsitWSNT0SK
94JIZVvpuc5oLoHO84OZF1Yer9TdVq1J2v5gjjCQM9aL5se1rIo+7wEL0N4xjgimx2rTrxEuLQ36
EIbNhTF84vDbEwNVIrRfa6YAZufREPMzsgg8I/I5gEuilPOtf6rYdT5oufL3+Nl9fVBa8pbsqf+5
MIwiSUhe8CxWUMP8XjxQ/lCa1QjP45nxoOhusXWdO9ZPq5NZ+wLYsCDxQEMmbiSmbm01SYLabWv+
FSvqB16wflop4RN/w122G1qq9SF/IEFSgwlhTQ7+o3z/dKKdE5GDOZ+TuWr6y4vqJ00d5pUG8HN5
SMzKVqfnN7LacMJcx0LtQjuREDDlKY8uv70rTEDmXMQCruKUTRJJGtXCuB/q+0cJ/yobfn6XzaY5
jG8nthkqXmk4K5ull96IKhzBzTE13GjIeaTsrGOOgA9D/fu3a9djKAzzx4qge2mOynl6qEbOTdKA
uIkrjJ/lpvCydoxgOQdRsLdUkFJgYu/WjQTKKfMW9LaIsRIZYDhIEtoQYD1LlWt4eaNy7RwnFc1f
KInoR2J53KTU1A7ucg65fCty+GKSEeoxENvb8ycXoYPJUbMteLjT0JoRJ0u/Ou3W2PRUaY0CXfo0
BwgJAoTb8rDWw48nSDkmlusVT988vWRWnWjObsCmgagHLUwu/y/mCEbmVPBwMttgYw+gXOE1FvDN
X5N13F2RCmpUD8GSOEjwRyRktLGX0JzB2v/U+8KmaO2w4YFUUwBtXJzJze9kGjXOjMh+KhZsUgTX
pC6dLrz29YPgknFtGf4oySG7CZELoE6lCbuy7qxPnBgWizCmq2munaTD/aLU2Ai6fGseNAGpTCiF
NvCtlvou+YEST7liSlHujBMhmYjgCRTS4nB/pNkH2y4Xb9qSkzBSr8ABMQWrXUTb8DaROyUPy4YM
nO5a6e0SHgZhh0oT34DUZQDglUgjqFC3eJ8JJRWHeCfCm+wJGHZ4PbQ64OIf08v06ObrY2rpBAog
EfNFsOh9XN43/nw+FIdCCD9aAcqCYMy4PB/uUq+yxpLlub0JoamkBQDShNmf8NLd7LXOwSQn8n+Q
Q1AwU5fhLQihoYlcmC5RlnkjvbowJdSND8tGOCqvRC8+H1EB88OoSAHKGbK59KH75kEDpjStX8NC
h2mfpvIZE9ABCvslrMbuehJLfAriZ9Qnw5XnyNFriqjYR6p9wnMyHj+ke+L74v4qaqIw1AQnr27Q
6LbKdzeKrRVj/LnEokVnsEkQ/sqmw3XLKdrKZj5FNG7ucaACcefHnV9B98aB9vPDsN8OnuYzxrtB
agm729sdMtgi7SpZ7YRztwDav6NvqanZEtJl67yYs1LzI4Mtuc8sH2QpRs27ux0/Y+REpzD2lvgN
MQ2jgkRcHAAsvAk4qWbFFaQXyAPtWF3HK2g+6shk06l5+2JIISWx2B3P7oCv+6uVmnJXCPF3O57a
o5eu2b1x/uS0xfA2GrFwlfM1COupfYzV1QeDBEJOAmai0hJC/qK1JTV5VtxChp5RGbscgcJi2Tiy
xH4J42loZj7Jube1qLX0QnWAv0r1cPq/2ayq7QvTr8Q+fni6Ia6Ri+g6M5+aLCmxscf9y5S1zsIr
AWj107ikXsXuLQbOmG7tkikUetL7Jfhe8E64DIGzkS3UW47escRD8hlMUXhR4YGPMGtZ+9dQ94mI
rKd58PJjG5bgiqre7brTXIErrd8B/3S+ecNcox93Hc+mtuzmVJT6ZZwWnYIJpzcx9PXAzMxONUaU
Hft4urKaKvQuqlzGDikVcaCgxsaNRygIwpBMNPeXN2SkUdVPDX8ijS9uo4Edl7W5otwNRpjTvHLy
YqWw7gmDM/dZlr5zFVDQfJVUa8wxX0PVFWohipVDvckDPSXfO89hizxWFWdh+g1vP7kD8t6SzUmT
JZYlckamw9WMIUoT7sINsQ211T36SMa09sT1ZAOOINcBaQdez49cF/okEu0Fs8j+ybo1d5A3R+Ru
d/9NRa+rdq2VtH0UY4pCKO1CCTLwjdsE3yiYBUN9T+GGmp/VBTIRGAPbOVYnXidNMkqzOCt1bQzX
BfzuvUf0xb+wuDTN4Z3kPO+mf1T0p8siDNTNT2goTE700z8N+1wTLsAQdCUAZTPYt/i4P9EBEmXY
j4wPYFKVFuZBGn9nznUKXznBQn2RaKfmaxH4cP2a27qMAh4IVbns2gKcHjmyzC7BFbeB5ng3d1Vi
25Tk/ycnxORhpVh1//0iAIEmNy/3TGJ4a2zSG4URfE85Oq/LXq5ujvKvEWdCHh0aYRGfu8Gp8r1N
5GpeFpSBRWxlzDOS1bIn5N6kn50zDTklVFDBJTjPQ8qzglCJCQSzTDkegFSgV4vBKU0C2WgM2aDG
+MpuVCZyJurrqSkC8ZYeLCKKgZLHEktvJt+kCKaNf8dL35TCmOm2IXazKwOqPCuavprt3/7zAB4h
EUzJVxANBb30E5F/9mXPS2omnAtggl1nkpud60+vWSzeZ3x7B0RdR9MH09omxl777ZK77Bqj4gUt
lfRzFZVkWwhpsblG1bEP39L6uuBK/m4m7A6iisuqylUclinxYPZjO60UDHwgRUPiQaK5hQSOzKNi
xZH0gdVxzE1DNs/iHLBtikcYnTD8l2ak8mnyUSMs8D/w6SfO4i1m3OxVu5zquD7g9hGHlbzqNi3N
z2FP8ElWljX4Bz8QedaUMRhcpGdM1RBl6gh3Uxn/27qkh97KI/F/qJmzKGKbaWzSiHvwOk7luOwu
aQVkT5GilGhgykebpCivf2ZZI8P6k81DZJoFauASJ2TwAm+vREIbBXjM4rp/TKV5Sox7cgJFB9Ka
PhbT8DO+t97Bu8SC54iQslGOXPxAVv7tRiHHGSfEH77jYyFuq5KRfWeZaRlQbESRS34FzSs+77sF
1KniaeJE2m+AAjUOw4r6cAODo1sb7FG96i13xYYMiA9fMKClrIdxIivAjvgrJyeo3O2aIm0TTuSa
QUuJu9tSe+qfV+xwkP1K2T04FqypmL7oPsd3jfG0Z1T+aP/Wb0MIGSRFAzkmZk3spa5XsDqRWXuu
tmDbbqQGiBd6n/cwHYYvJmVwu5XrvVI/OcG826sg90pxfLXaYOHh9InXlROv/CKE0SO5tudvel4p
+Bq6xaXrzjVLXi4Xszpbwd7lneIuUpIIoHGfZN3pyt7JepfCZ2wLH4/tsTqCFQNqEZCFShj2h7Au
21Q9ISmmoViDM2kY03pM2QUKG1ghHhxcsfDatjShL+tv/phC1/QZgEzceJr2ZVfCZVXy7LRv1CY1
bB46mQFhjFu0I9dkz0wsPZPmeHK8dVkLvGKU8ieVujhpupSY4nxWCahxIhBS9gHWUYWHGuXUMwgt
ga+ZOTEhYpIDe4zTPv8x6+WEf7zJIsjCHeoHbH2Krstm76sYEIHX90ca2wXOI7vPNEzswG9zw7Gl
9cHNjwsb1qQQaloK4UvMhGwzvw1wjK6WOM54//3tyo0oIE4BHapAejKXQl2NF8D9w69YnY89kL56
SIMqr9YImgQyGo7odrtiIcBK78DGl1PzQGUGVA+Px6dXd7jFfzLuDxgLyD10g63nArVkXYirbqPJ
CAIATn4Z8torYvaqa0dke6e8vBAsgGZlH1O/rAJ6YQzPhHJN3gZ2m1TQ9UTa6jdffe96K/IWjd4x
+2jeeG/3XLqyr8rMhoiI0fleCX8i9OsH8XvGSNN4vCHfTYFGa1FjPPV77kQl707NfBZTLGoQJi8j
YXqx52G29jOQ/3z19ySs6h005m4G34YbTvrBGB/VeJ7070HxMh9zIC13odqPmf10zk6UYDQscVxG
mgdKcxdiM4XnV5Lm3kb+71HlhM84UgPN2gQ9GVTbWybduU+D9ninC9s2lLUw9bVmhXLWNZvelyZn
gcz7bGL+jIXRX+dZCZ7+OSRSZ6pBDXTeq/76Y4g6csLXagonJM6+6ccFwKVexRI/szj/TlQAJIFk
GFV6tbja8YYFUrYwhnOafK3uZG789lKx4dy/2Kyw7yHFsVHIhQN6wD0A1wNvRC8WNaBkpT8z7cnq
WK5hdFXxu+wR2FWyVof3WRfjivENeXE9EpRcgJWAowZ5bK5xH4LBgzg+Zv7p+P3Pbl9EUiA2XjUY
n7JDzsGT04FjWe4hifkdGZ9WoBIzgZ86YvwZlEYWXqg8AaIvS8+VmB4IH+gAb+v/FGVwJEKAThnL
btmUmOkCRLQn1DtKO6GPKDah0Mrt7+b7VprVzl9jEsEUT0iiuebsEmRDr4wa1ypVIHV/l8xMD3zA
tgLiothNODdWUyg/Xh+SyquphSPWKHvBP8g08AuQmfm7hBREDq/H4Pa/atvoBSFAzUKEansix/ar
ELyNzeYPc4/joETo9t02phDTo1NkAUgQSsgnz8UTyHBdfO610wbwEV3sgQQ8l58XEl1slyBKB0p3
jxIGI0LbI3K5WYQsBsVptmO07Fkw1kZr5o86Qt6E0ix9CXZHPH/ylbeVg+n17s8fTnunPRbLGpeD
HoNJX13WyfBAvXGjsVEs+HOH5sNlSSSZBnZp7MkqxxiZ13Ofoq35Bh10ZoGiaj9XmUe8VicYzKEL
jdStQDLohpUzsMLHanKHzLuk3Y8Wt0mrRdJLiWED/IofQMc9Vma8J5FYvakCA4Y+kmZdtQlvddYu
9hTCgvV59lF2rVoVu/iFe6Hst2vJKLU91wR+/HmHMjUOR2WHpL2ZRu6ixkDnZFGBXDn2qjz3r2Uq
qI1sywcjcRQlkBWeBgM+nlHy5BfiUV3lcP25qlpoqowoOyVdDYCTNVimnrAMscn6qKw4pKfFDRUs
tLU1/kzejwEVO1PzbGZ9goBdxoEay/Flzp61m5hhTq7cjY815L7osLVW6UMw1zri9aNvqJmAuoQP
qRlIYJb/W2thcPvLBfY+boN+RHX/CVqWPVuvTSWkbwlQYCgW74NC9/iFWYFq9ytgdYhF+7MK63Nz
L290F4TB9zXAnd15GL6G62PzsIk8UWf/WdU4YHq3TRhmub9Xn2lC7CB+KN7mgH1m4dTRsQGRAFNY
uQGjab+nd5nR3Zsgyv0Lb+E7Fp474CLTZBaoZTZDCTtTo/tfy0TsxJeFOesKTUEnYdIrJ29CBLDy
sn0aBQ4m7PY7fUC3NoAfni3DnVc++IccrPOtw/iJz5IuO/C9OfA3ezBEmFWv1D9yOq/T0PS4YDvu
xYNf7VtHvi1hbERZrTSL07yozRrsrpRyOUPR2+Z02KKAY1bDqodQ/Eh947ORlSBVFLOQI0+ooMfB
uJ3Wxl+x+vOvMh1yjgkVC5x8jWOCdblJ1Nzsu19ntHy4oCnNGIQEX2d2EMlkCogq87ytBcZZORpw
JCi+f/QpXfsIc3u+1J3tjzwO02lD0I3WJIEzc+rjxL1cjp1EDnNo1aRuv5320UNwCh7+2HqrxS3s
gtnhq8Q65bhkXQJWgDg2LTGU5txKv3ej0cDDkqTT6Nmge58jqT5Cq41+EHMM3w86rdd27opbNy7H
iZ2bYpkJXKRGWmHAJc+n7l2ljzC0gPe9CnW693vzamcW2AB3jWdELuoXnHBLQBmxdn1vQqN9zUHu
oQ1V15zwgdQ15hGfvNL731slkWv8NX89i/5i8BTF1nZHGNwyp1Pmw989dVBaN3WLZdK4wlpO3hNG
4VPcevJunctmMbkymMV9Eq/iqBJeExIC7jNK2DNb4PTf9ob4K+kvBZJIzgVlHObk0Vm4oDjP1HKN
3/YSD9iRj3iY/dRQZ4HkqrM38RIwjQaKzPpSyaomlVJHsBWjoVIXTzQm8kRULehjC2C5ClBeQ+5e
P0YLRAxIG5rW50zH4UwEcP4E2eOfO/B6cRDSS08YW+TEgLGceaQzltp+lKq6f/DN7erhqhH5ytzg
F+AMppFK+KwAq8GNatkcQBWVq2PXFpu1n10ibisxNrU1DJINj6HXa0yfjk65NwxpRg+yl25bVEeL
wYtHzkKCKFFpQglknzsnWebjdT/6XoJr9hosV6aW32W1jS2fYkbeFAF5767Rf7C70oIaqRPHa6uN
fZLJpWFeluQ7WY/M/DV4UjczF6FtJcChFdxSb4O6c4pAOmC4MoFXTB8Dwd+fRbjkPT6DtAQ6AvQa
CeFn5dTfl2MUninTNJiU4wpHIJuR2I2J5Fly9rLcubHycXBJP73alAR7k3mfZGeaTTgjrRRZ1JB4
YmySChXV0qs9T7ZPzWj4L64N01HiTICsLDGV8tnVbcuIXNL9DQAmjubHIsJen8yaUPl87uHSN0n8
k2zoc8jk4DZDJ6QSNOttjs8XNxCq0la6pwwzWoLuDzJjJ5b3MjEwMy1SGoJKRwSN8jiQM0LGQeU2
9oRGkEXnkeYvj0hari716ZDVhqhRLQGgxXiNkf6JAnQe6neNQS87NDUubp+hnRqFReUaOgyR97H5
ird0BU28rdaAHiwfeJHOgVZpVV2C7qAqNti8Q6t7J/XZ/IH/VgvtSigo8ugqbyBwSWtVj0s+REdB
/4GHDFihroXqoIdIww1IaL7p2KGcVEafc/9z15IQ2iux3NaviMlgnN7S/LNEkoWEDHbJvHIihcOq
+4TRbPe17otST/JWZV6KjRAphlpWVP0Uyr9jFf08NkJRx0yasYQvYcgYNtnjkAnKRHA4hBY5XocZ
cCBwf7nvYswjbbmb80P26GegJ4wxHnjWaD7lEtHIlv6GQYJ1CVPmZTzrm6cT2/j+wTrLosfXqVan
tXnm1Z9R+wtA4smHTPlvX/KkxR6bsf9MwUmJOVQwoLe1DYOpNwMUGHR9VSt/NjSFdYDCEJMDPkdi
Iv8aaZZwPsXdfk09WMe1V8lVOKhFNTGjqtudgY+G1OSZPgmn6y5gj+Gv2SuA+bzrEMUh2uPFl1Lp
hiDxlKk+Qp0psa2/H+3/sWqY6tSKJQ2WvwwqMzaQ4rNutnaLgmemGj5K0rFO9xhgTZwTlVOJ6ISX
gARP/psFHxWGx2HSACsx8oANeCN9ZERG/Kzpkj1izblW+opO6OmDxmkpQBDl+JEaYG0KRlKYjKpQ
4l7WowJZl8+Gz9IBoqensb6tBmwfRyRbqXxq8ZYzjtf+bIBHLviRDIUzCk4ZUQ5ZDAFlPSt+aSqX
UOSiUwk6PoqDcrOymzLy++cObVWkrzCiueNXUX2CYnCTArH86NAbwFBCmbzlEO7p9lZVAWuNX8/0
fJjYTLKLAzbHUK3PvD1ABHsi2NIQruMpb9NzjpWx4iECdKCXrOlmrcRWzXWrb+bax4tlU7cq45bh
GOxSXjrqxfjqmvPCv3TtSZJNi7oVtlwC2bejP6kye0NR8xDgulnE/7Mw02iBXjObPIClNMIHF5ea
pKQ2yzT4ADtkC59Qds4pyydsTk9R5vEqlf0JEXLYF25K/LkzsrJmac5j6DO+7NwaPXcUJw0IFnvx
Aq+nYbAl9XT/yGTbbV+KIAn3zt1ttUfi8IOG6okj6b+BxmQoavQ4XFbSsZx1GhDr9BRucxNJHXKR
OUjg5hzB+GbHqJWjvKDO1BxIzBZnqmN77HCh9Mq1Zw6VbWoM5ETOecWgdlPqTmldIPbHkpdDvTG1
vsnno+FMVX4Ga7Xw1Ccl5aqQP9KMBGT4pDX6ljgpgHTfGElLvVufFAIWE/66T+5rQeA1KZUiwB40
t68KeRsPFeAlFS7iO/PEsDP9gPyYcla3u8gksc27x7P/HmcCTYntkifAtMbpK6WEdr4YpNx1/oks
A+eo4qS5didaPXYu1rYDjTyfY2jYoeT4EYebEHGAjpNlYYA3tiLIG5umO07Dr3n588pN5JfKGGDt
E9MJ50IkIrQZdb1pfCupUQ2vDtI3hoqWAQN95xprjhHZgZUzeygdO6JPvZU/8oo6pqzeW+ehkB4F
75oAHrPHx4G4skVYGjvaKrJeQUByht+Bxb+W32+R61rjMjemjyzAgVnQ16bFHxWAl5L924TVLXrH
0rqSrOFFmYObJaEydRjIAPbUiiBy+vj/OVgh4yMe7QyUE1NBD1LvhNWMLUN6ASl+7Qb05+xSqla9
VCwpoHV9ClCOGREKOu7d1X5tucjvvcfu13+aNJ5o1zZqWKpxc1t2YBG7NaRPPCLYKrnEO5/pJBK5
i/gv8cOXLJiP4xcuNDQNWVD6R+de9zOMr3uwT6FuOCfvBrvvYGv9LyrecCfMW7JH8DnZhxKekbW2
/Y0Bvdb/Ho65NMPJlWaEAuKblrVwXIcMx+4kYtp6Y31X9m++kSV59kySff0AYxjqPfX1FFE4sRlY
+MYXRiUgiA9yNIBSvkgjajgXGUKwri+TxAz5Gs+iJZamzpsNuP6YzawH5r1pDrHJyYSs+X85/oH/
pP/xOLSsDUwjFGYhAD/e4Z42Fn182gHLHH4QcjTL6SdD1aSi3UPn2SuGPLpIsGGOswwAp8utfz4a
832qv8JKq3gLyo+ZHYKExDHUOoi8ZOEmGF96fdvg0a+LtIGqEWzd41HwM742iil7uZnPlk7Tnn6D
QA/LYh62WJkHUL3YxkwsG2IiuGpy6xFkXr09pxuBVkldBJVu7TwKgLryVvSIHploro+CxM2H/417
BoV7qJu6+eWwtCDXpjVntdqEg+nV0YPTB0aFDR8unSLURfOYEzpoanIqEbG+BgWt2I7MOazn5lLN
Q60JuU9WyouRvEJb8I4L9U8wQxTe6F5ameMsVEB+OAsJjrTUCOh/eGsG3HUjsI/2WUBTMjSXwj3N
JUtcT/EOkGv0Gb4XETWW0xHrasopDoT0s7sqjjFfg3odq+CHJcKPsQ790ixQYd46pFFk6LzhmESh
+efg5ITIQu8YaMw2tWOH/2Wq4x4bgMuVHHNqhtcwoPQTOSZEoajWmbd6Lt430ZiMP9L1cyuD5GrH
TyRBT+CiZlroXUJin10rtKjOrT7RSrAi+7voorAP/vwoC4iIRxheLW15O4U3wFuXfr7cAfLG5OEa
b/Cu7IQeHRkjxuW9Wcub6TbuESv2Q/i/C6+nEPa7tJqmySYaRrbNpZUuqjMVA01NlLTPaWNavvhR
m3aEURC6WSvlmOxdOPefFY6fJR+RaCL1nqn+fj9jTWoEY+ZrswIJD5Gcunpug16WDvIZUrFIQ/yl
hEzuvGs3hUDxb+n6KBIrMCmRHH3yKdxS2GSrFRkMr0PxbOud/FzNCuITMPceJapz49Cbmkg9sRyN
rLgPu53wU2s3BjWuzQSPSwxPeoCvlm0PQLv4wyJtalil1Mo2Nvfpd/z8eTMDWzLigf3AJC0dUV43
FLMJUbfabEY7S9t2UXcz2+IbZH/OPwwjkr8/AFIa1hF9F/mymbDdrOPa/QI/XJsXAeBwSuNmfiTc
DPn+dhRq1PvcpZUE5UVv60TUvO6hnOFeF/aqBn9XbVLFcN+7lpQnRO6Lb1V7hpiz33+d4g2uGIk6
WlwBA44qfDLXcVjB+iscMVRkYe3nLXiNC+0T4F73QZ+mHmqzqepzWbl8LykFu2/Vmq2knvmwH/d2
F/hWM4UmZwR3HZK2eN4CK2KkkMaJXzfl6ZVtssYHkpDqpIdqMnSerJ9caU6kiI+6VmirwgJ6U8e0
UAfF6e3NXeWD4JS+QqOP1Qm9O1v0cYGqIfjSaD/RQaMpyfd0Izc6EX0WR1ja0G0EIY/MzRAa/SBI
PFL0vI1P0v5Jxu1NSfk7zXIcRRfJTY6y/MhpzuWl8HYInniydol1Qc4HjTD1h1ajnpd46Bch4UTR
ekPnlAYZyrH50VM4yQV3ihze6F5aBNNhzZ8kYDww0Z38MYS8eUWfIBBc2VeAfTzsMCJpdxT0cFHF
e4R8RboGntDJxyzy6p6TbCYQwpnOZO+LQgI/RSM+FuUTHixJefkKhh+F7ACJ+tdp9g+JXeEJ+ihL
3a/9wtrbQ4b8prswmah+4u4MbNX/YvsPQHKMIoehRxHJl+ZlzLuzuhp1hX91A/Welm4nMPtuFAtZ
TZica6IZEjOeoihG2fTO3hmZZfwjNBBE9bzPiw7u0FWYroTBoVrdbmpbdHuIXJqgoKNFNZMT6uEr
w8wrJ5pt4nzi+Aca76812fH82V4GZ0LzpxZ/pi4Qb6VmzS1nqvF1N4YqCK8Y4WSiAHThdp0D49Ir
WqiPN+wg8vXm4gkmslpCcDcKkkPYufLodfj/ZmrrmZkURs4eE994TxieDh+nMZloCph7rY72gYdh
4fKo6fFeyG0H9JO/VTmDAkSYAp3yG5Nxs6cWp8HA+3Hse+XpKksV78D9PIRlVHSeJ/j8nWHtiJUi
f6rxGu09G7L2hQiFteqVkM89sqFayED0TbwzK9HE3tLnn9PcL2M2Syflx5tYav9GhXcuNjpn+U6A
D1TyltP+RB0tG0RhZT+Ie+HU3WiuLWsSWVDTLEWLVszbi8rMNI/ZxGNF0dTu3CbIIMikc+v3LPZt
Z1a5iI+3Bqfcnz5QZa27WMRjjLPXSDzdsI4+ODW8l7mbjZAh4Nb05zkKMBkaC/YyJN6nRE7QP7tv
SBintGr+uWcyFaHt1in5xvREY4vK6baM/PoXUdk9JfH/y+CJEq9RlQGghqOfbEky5qDObc7ytgtf
5PRYddiO2NBvZI/p+OZQgZJzAm5Gm9ouzVfTigA+cc3fPdXCRNUoKv8MZg+P4vqBJrU6hpytofvZ
geRDICsSXqZfyD8HLh0hj8jkxQm/SCShVC8z62v6L7Mi1I59T3X7DW0ERE2srgvmLCz1ODPeZY4J
FkLjerpr5zuSI5aWVk1tnV8MP0Az9UqW0ZldcthnvtKQfj7trVB4xS1Lwakj8RwcTkHiVZVI6azx
9cQVwxr7JU9QDGbxeJ/xS7FfOIFvqSxFL0vslU+ykp+aDuNlZCfbYoUQP/IoQARb/ElI2GpzcvGQ
soIwe1GoAmWhdExYcoIhLMme23dHOH3f2APhi7ReyBMCtmt0r5FcJWFb0Sucn3ZH20ZQL1I7I94y
JBCC6duLgfO6Hns5/FpLTR4wVNC8FZ1fCtDR2MjE2KFrE3XBFTBiWmQrunjjWMyojvvhJUJD+jZK
LIkHbXOzyDQarW9M8omgKIk+YEkmN+XBOTfj/l+cuPRnR9NTRnkobsW41QQnaGuQkflMWB+s2lPA
MJiqt9rf6olayHEABVVvy6YeyGHpg9EVcmrdWqhmiI6JqIlP1RbULjvNbzUsv1wdBdWVkLLma5H0
AumaXMdvnyNYpY8FP37rQhGhG6jqldq3vOm/VYDdMcpMh7WdKSEoTN8LcPN3YFe8cIJve7Za/CzS
L3mvxzQvcY39ALZOQFdfKmTuiDBS15GHNwZp9EL6LumX54xfweLdOC0cTAQC7tuFrdQybXhOCLFh
LY5I0PgcovM920uhO2GHUT2UxPpCywZEeHNn/36k8wi0ZIRAWXDIYCO4+9cSC7eH14P4zEZx1lUS
2DdLhQOa8xp6flUZ+kb2ILpK22Y1PP+HOLGbdjJA7AvYazvEEffZG2BRwtuQFV2vB+2vK7atf8c0
Lvd6ViTe+hB3WeyT+sI11xo7mkwQZFOS/DWH37f/wSOmQM+W6kYoIl8C7uIZiVC4lJKPAWeraR5O
e1ZXA+u03Uo5M7IuBtUMGOxa7wiX+wJLR2x7tT7aYA7sJLifnOa44KksqiT4obhcIMNkTVdjTb04
HdQK4l5pA+rsX1SPD1Ggw5AQxCx5ZYOUcO9lbeRDg9oO2CWaXCGndQVTSBr7H1aLjsGB60anBfQL
9EkwYSqN73xHScRJ+f7NhZyhLrTpxdjWnCuxMS3/8YW5/8i6QXVU8IMEXWMl48C5rcnj+eZSKilx
DJuiUfw3zJ7cnK5qLMNTtpMtbsDiTKEz/JDaBHeLNHt+xs/V4RhnUt+JK2SUtcInoeD84wBj50vZ
lBZoJ/0Tog1UQevaFyOE2d5gzamhwtwUJSnuk41iomsUYF5Q1VyO9Bnuw8LfRk9KsXBAsjxImnm/
v9j6RJ7rWX+Ma8cHtv+MeJvzdqilPzUYL69OPHfJfMUUip3MUEkCKyWVdEjCTCSaZRfy9S+HdZZU
LFlQH8Kg35CJ0PLKcLJDT6HyzaSwh2wvZ56wbyqJQsp3485GwuLUMIlEc6s5vAQ+lv1QF5/7RDzF
9GYnjaqBr+puUdbWRmdk2F/zJhVxzcxwVEWgKuC6Wt1Rh7fguz98rKWMEfTguglidGAXcUAoZuiJ
M4j/uZs2uF6aQKA7DaJES651bCpFwoYQxGxKpqkG/+pfcGH60M5io8oB38aezpKEe23GrggYQzOK
p0ztNMPGIfF9ebQQtHzOKC4uj2wJstyjnPhHDDxCeZPgc967rU/eOS/axFZxSx+MsxY+zBQS1DZi
reMO0T66cHEsUtmC3XvYxmSEqBQhU7sRkwC3EGbOzeRnyxGFNMKodq5+yfSoLfQjxjhw/HJl62/r
cG6p39aYLy/G6PY2tqDouijt1asZYWGinKz6KR6tatCwsFz4Qb8whn+b/Yc5cXnwOGAQrS3sO9aP
vgi6erfjUtVc/XxFwqRH+Bm0M83Pgw6Xr85Ast3VSon3IcKLVaDbZZsIIY47Q9GFiT1BEjXEMxK/
obOs5sxfDLXetZxFFcS4uqE31N643eITAXxCrjE+rKd/J4qwwqSbRvkuPMhaLk8uKe9wq6MiVkiP
Xy9MEhe2fEHfOU/N+CV+ynRFTfGJ4RSwzacBiQ0e/6+EQUuLTnXp29fXIofygUX9jnxvCGBy8VQv
64+Ow7ki/WV9LeNtNqH/UXy4GZwfgGWy63ldZZbW1N+IkW+BIRcgcRYinEclAOGjRCbt32Ok7nq0
O8nf2WGKVT0InGJlTGbnK2hDysEZ1d91gYp19Pzld/G1AMrAwcRSy9HivfNPFiJR8I+XOwohDwnA
OMjEQSmXp55OpkB09mHY5VEY1Zv4xMONoZlO4LYI+dwHAbOeBI2LsQb1rJ4rhq1ADMoKpnia61v4
7UudvbJ0m84ohtH1Ub6dbY9qipVD8hHOp17UboLmovPgEvzLO+XrJHO5rwAJcVfC9veLDVUXuve0
zUw9GPGpL/8N+tOh15iNOeuMrAp5ZB49fOl+vSTwyCASiVgn/75C2CJESUFT4OWBkMyhlqPB1si7
UWBq1vjRIqaH+0T4HgRvCNNz8ScUE4ltz+jBMZnkCC6w+oF0QOZgbnp338FsRbu0VMIfK+gubsgG
0I2pQC2WQzlG16XzSKlMbGCg5f9bKvvVwtFjx7aQRanekb7Dhy8xm5e0t572V2lPEtCNhfArl0SM
4Z+2aMh9S+qS4AvDhnXNlSKthti9Eb+QIqYP/4DX1ei2lYwnmYLh47imK++hBephxC7M1c/GYYz4
C1DXWakElDPfdSCUUfUmAqdbMpjpv0KNJZSP2+7y0AgkqKS1Xc7sSYnsBzN2P4UgAmJbf6hYJZ4X
VcTgPGrZLg1LhiBuF8jWGVT2HZV7jXO46xyuBZL7JkNyBd/0LUN8X2DsJlVXFTTqkBU3/h7rHHdr
NT69JTkQ2+4r3RXM0dBZFRpFwhXDPgdyNr+GUsVde5tossK69FPHr/kqKtASEZeDqPiZUYSl4eVI
RYQI3eB7/U7ji2TBQu8x1+F08mFctn4DeVJryGIOsRgniejPrxlcX3u6JyYzoKZT8q6/zrpXSru1
851sNDTBJE+kEyOgscT25uObNqBcFQmeGb6G3w4evahe9domynDDs5QF/UuKfk8nLEZMeJPxgjKG
cOkp+joyPIPQlKNbTuLNQFDCtK5+GIxPhCCwN6MvchJT41Z4J30zkYr77zA/471NeJorI/WWXbM0
eBSrP4/meYq2nV4TBginMOqWX09sd4gfd7BL5lCpFEFWTmC2W5leqRi7IS5e2gYJRliZsaSAruPH
oViWPnqK1lqF9Mc/AWiCOaeJ5PtYh1AEADLUDEm5u2DY/VCcyAxQGUDc9OoZ+qF6P2crMsZvv+Cf
ndATnIRyBYiOm61XbBJFsEJcEKBsmM0RLVDI2fDhI6rpiGHYHtNpz7RaxRFR0z77lZ48FgloooPa
bPBRRCmaUH+l2o2Qf2wbe/nhEsktiGBg0DXn54r7jIRWD2uWezVFnY8ztmE7rqPD1DUpKR3U9Eih
5aSyirKj8PzOwzHofbb2iTyowAjP9VKEn3QU20mNo7Ydv6PRen4vFxEkMRsdtQiHiHJJ/DzmwimT
aLQxgWPd41kH1tqPRM1G+8wrxLLo+wawvrgfiNtcsAWjdlu+khEnK88ys2I5ZU6QmT3Qc7DoeNnw
ObXuTQ/zKzLjtz74SBDUHfUDXHoev+vFsXSE7qqifHJ5A6lIYVKb88nzTTwVYHDLBcDIykSh3/36
mDvMQ+RPgpClmdGb6zpJ8mw9LvAlOr1mqachIYEzAVUJYkVXrrI9DYvu2kGGMSr1j/KRTmeGiqdH
HzgEb4x9yVKs1q2Wb2bCE6I8TWJc1bbTpL5XtgpDzCTONhIGncQzrim+MZQSzdRidIItyZ4fabVe
RIgSheVL2mTwpdmV3jEUzsfJ3lpWxo2CcizyebslrR0gNQFGpYghGKr85y67e8ZAlWpkRQ0K2vHc
TMgb+31VthDlxll9+59fKF+35Bo+kv2GULFbPMjuQ9SMFBTz2h6xrnh4N0+2LAGyDPYYTKjig7V9
ZOJ7dfGasfDrSXtnDKLq+vAfecNqmuQIaCXTXmfq+vAQJAd+SsDq990UJaGFLVtJYROwZh7PRWZS
Q0Xa/p3bwwSgN4H12NVAg19a6nKT+EmliTxenqdyNJkbxzV/21bqHsR5rSltjVVrR/WHPSBU6zy6
TeQ7KRmaWKZ40HqIqAxTmehhWyrtdCNkkQ/LR4LN+xxV1pLUVyoBVHoVHz+TTj8HfNorYvLOc/Ir
WXRtsK4tunkUtQKyKBsP3pexes1mfWWJfD1Nsi+7krDSqsXwCmWkDvhdLBVp85npe1BtGlYSoB6a
HElfpY7QIxi3f8s8DfoPdC8llldHikOqUyRWrrN+95EMI/bqLKyLQpFslWJZ6W3VivkhX27OdzWY
8ZGXDi9DGpqS9Sxy70FuUV1asDQgHR9h82wYLr6VOgTj5oJhIuDsbCdjkWghYpSayM85Oz7gDqgg
6pN1NXFXh3aMdY9+uoSU1XhZRCjmgPM7ANzWBZTszDfckpuvhTDQkRg8HvgPxE/KTpKLmYV43bG+
WTDw/+UhWn4TD1FQAmI4pH98zUS4XC7QgervI70SolNM5XGmshLpZplwCT4WDJRRjZFxlk3L5U0t
HkwWSuFc+BsZx18W9jl4kaIHdz1HXaxx+3TiYBlf+Y4IsgDVHBzTBBLWcyLZ0WwAxGRjZGz7mb0C
/m9tm4bdPgMB0X15rirz42uEjhWzsCdu5Ht1SX8gNSiAh95KZIUTarAiV9ZPadqvtmbm4JWUyCeo
/wVmheVeIIN7dUBp3Yf4+YbHwH4ystExctwSG9tlgjU6n44zCe1y5lhi6UAd6ODWBzkah4ObMKvB
SaUn7gyIflzaiNqttFK/rRDxABzHwuNTeMvN2KVarKMDk2y4Nr4kaQc7GaouyWZYiUzAQbK38XmW
x9pBx+8MyS2G6p/H1yrmss8Dl0LTKTw/44YtakVE/mEdjc1TwAscsZ+FRO1AdflyfwLIyQ9/3sBq
h+BDqduMzHusya8+wEz6dy26m0juXFWZWOv8+UCR8LAUVX3t2gO9FUqE3vL8Nl38DKxkWF0/w2EN
RE9FJhOKgylD9SYUo5fTaz4cG1ioKQNhf4h2PGrodjYTAGCdh3iY6FjeRuNQQfmK/tYaLrFtdgeS
X0P1pDjSIm5vWDbbZ8RYbkZ+JMf7+hSIXQzQv9RaPkIPwP1Yej/Y5YIE2CMB5pBMY189JcxDSAxF
anfVY9Ge5bPriLOieWm0AQ1PssxqjHahIKxg8DukhKhGEuvwfgdT4Cwpu4U2N9SOSWkff/MyoMC6
Ilz2Ga2LFFyljbeuRneE4Eq4WUBJUad6e3Qs2tqBYA5TXf9zI//VGqOY8kiEOQGu+wI52fcEp+dP
fM3LMBowr0Vxu+pCWcudlv1UyEaE2s3X1fsFufR36jzlObbSP5HeyHm3XTd3DAlqSB34VYMzoz04
wkAMM4QsAlXRK27FXbNJkTgXyJC3RfDZFibZXsEBm4B9gvgFNySrj0aetrQdtDi/h2DKatIyIIy/
3Ahs6/WvwacsRHriKcKkErPi16j5V93xWR13xTRQqgt55BEkRDhAboIh7Zw+M+/YVDWEKQfLMsJt
45SabZ8dum1eXEn1WdWOoLEaoeQ/ef2aYk8YNtCEEkB0Y07yNk8+hkeJSMAQkrtnV5p7lpYtdw67
YYxpQhJgGakEhBJGbANlwx1jlxCRYO8NKH7If9jr0irXZy9N4UCqPQ/dZn9w9zjJHSsd6h8ax4dI
KQBxqeXY2HtiShCCiwzum/Vc9S8xMOzACtlszDtusx1t/y/LSMC7XIfcQqxL8Bp5brDAxHzoNgKb
Fue85N71K/yCM2oF7zxnnR6avegNlDCD9RdY62Td6si6J6ZdCT21tH6qU68OTD9EBkDzwrKv8EO+
KxXgUFikbVaGZXTUG7I0DMGxUBDkwVKRz0hn39j5D89xsMof8BPgK5TMEyaxpjZLZbtKPSV30Q+g
GEipGPgKoo4NT1kfZu/aAV1OeJV79ErHv0donZ4GKEUaQNHyiw3F0T7i84l7zcl76f9yB7sSYtym
Q5enJKvIyUc0fWPXPNMrbC+xoLdlPjGmQbct80Rsu4bBnn8D1QeYPnA7SEzjUEJgGy5H2vwnSc3p
YJR2qjkp+wcxiJVWA53it8d8rsiuIGNOZmMtlO3ur+PrR9155OCYHK0JBN0ck3T4dfB6xtHg6jOe
uoTqKxh6Bb+XnjtZPmDWHXpobo30hiNY7KEq/Ck5o3WMcPaYzDNrkx0DjE8NlTZWcVBGNOL5ZVT0
d0YezV6aE2I7rCzRO91pYBwzx7qKgLXn+QVXoeda5rnPEDa+R5tQI/XKyfpONaKsLBZj+nEioXu2
F84EDRHd4pr7isfRBudh9mJ2RL5YCCCV3asdGaFchIxcmlRBbgi7yg7ildVcPuxlJSfHbgDn3QHC
X4b4Pp7ambGMHxf8mWCThnnZvWg8bbQRXZtPSC8h/eG43XvyGCzUWfQgHDNu5ksYGwXBQGo3SvnM
fHTUO2w9bTptHldWs++9bIfBtWcLaKCsjosS1/mka2f18sPJJpzuu0kkUh/F8UiBgDpOs6Igj4i2
S7J3XlLl/VYUDB/sEvexIvFITIIPaMW59fjra8HY/4Sd7z7tSkoaJRNaB/He3hZl1Egkgu8CNdUB
Z8xNg6kRV2q+otB/XnSN98YC+LYR5tvuy0roDjjIitBS476iBqF5gSI1t41Ux/oWyJ3Fjg6nVgVs
RShY4lqPBivmYXeXAuj77LPIvqsK7/5TuGhoFfNVly55/Grc4aMBbbmoaC4ejoVShtHcc3Zt163w
ldPbUn+vRxsYf/mcIQiz1B+tYWAXWx2rR/ULaCLY37ujhRoyxGj29ovunxO37T7hdzweuHntPfa0
TAeG3P2d1XuVcfJDLWKPI1nO1C037VdX41X28smD2R30s2vHeJsvXZFhTmIVao2BBobPhLPXGq/b
F8zilP9Aa/GZYl6htYeTOfDCduaXVoVoWlgomLPOYZKESKs2bHgjxgbYiF6vNKTggddCQ4ly6NHv
FtSTG7zcalu/D6sSDe3AxWEQ2iJtreDJHq4UzjfchKS+qTl1KnICRRbEWeCu8uP5jRFSWYMtHRpn
+oz2FynfkBcoWCdXfwEHWD9XxoGD1a5pijFzo0Gtq/8Hr3/9t1LFyz0Legp2BVl75B0YZnlWm68N
j2dP84lRLkcx3R0tHKVpWzhBMmaEYOWsNC4vw1+A8wSO8l5+0EYLUWZf0yg5f4hSU883ksy3qjnX
PvSnmlLtp7I4MyOk3wfO/wkfYymDCikjgz/n7cBY7FKXBHbOLkrHfOxrAnH0Nvv+f6/e4gldqiev
Zlxegva92Vm6ph05LgvDyYRdrys/AZeWe3Le9bEKfyXIIZvJdnu+VZ9gH9ujnqItzklMdOwmsHhi
ZkXDXUAfTR0vfeYTDPCMYLG710FKyl7KAQdqySc/vqMY2uQmoGZp9lnKcxfnF+GdE1dtep8gfapN
2E9qO8gG5L+JTaiTWyoo9SG8sKP9SenCeblTjLxuk53vyw4Dlv2QoiP8IA7euR7NfU5NKGM7jKuw
kYBzUVvYSwpEcrHeOe2r+8JzMSXSNkY+PsX+XvOQ499HdiMKSFW1VbYPChAVBsWpkwoeSIfBoAKd
y4HlS9rcvCoyTrTpjYsbmMCi3ZUeEJvWVRAg2BhX1qJ/d2FxHlNraPm9/qboPVkWCCcVwIYGeBW9
NEAe5kgv0XvjTVytiK4nAOKu8Et3s41GIR+S/D2cnT9ZUOZdDtV3xIBwRBKjPp9zSyU7DY5lFCFo
DbRW1S51YpQw4xITQODUo2ozxBVPxMxr0rwzEmtc/L06FhLpmAKxfqQ7cR+KJQH69BvgjXflcl9M
YE7wFaIMZscz5FK0IR4a390JVDh14Oa+mQIjZXAVTegZKiskh1kIxzP71YqrxFNgDP5PKV10bk4T
j4fyIGwT+v8a/Qn3U7c+1jlCvPaCJ4L30maHG6Z3Ut9wDl7gJfkPjhcobugH2DhqISWKBK3DJ1+N
tgCkDd9ejA7BCmDc5rXNTKn0ZlPFnMKuD9TQ8AI2dKmBIyQ8g0xcquxVvId7swp0kn4ShL2ADD+Y
Dx0hrseABttcE8STAsj9h87vpRDRsPD3d2jzebE4qJWwYwcewWtpQvDk/U3Upu4ohTbvA3GFcDnG
jq4YWbfoYlaYZOdV0jdC/6iXG79dDqod/M8THLhgPKtOxgVIkPyfLt/ekfrAzEdelXvZ8ax5DPpZ
P9Bo0DYhjZiCaDyc6v1X2aDUzq0T5hLG+uipoX4vvxTD8vS/V5c5mlofCRhNvDy0fOXJ8J3w36ND
SPYo1pDT7KL5dI+wAGhDwP3wWj5pBmde8x4xds3G+Pi9FLmxiBx36ganLcy50Bjd8DL+EcjpNn+H
msnQpIFx2MES+EslUflY2hvOEn/+nH1zQ242ArfSBzTktHHFjof59NpvHmjJXZLxqIxLRRLSwqtI
GXHDc08hdC6q5VWKf4Dhsrt5hE3ovH1M+tq3XWT+D4J2X3q8zwRoxZFFG7okSxjlO4sPugicH4kE
BUP4WBv4mRtybbxRM4gaKzmne3ZFmA7gm3ghyZgVa6WfF83bC30DNbsJFOn2MzEGHC9jHlL1ikie
NYyhfTcP+auu1Kky3ZLEDjop38yalPhgt/5SrExXHOzI89DklZb1W0gqOs5a638i9nOP678GMTIB
5JdBbMym7VdKmN41WRM9sM69nsV2DU5j6yCOYnkyzbL8gEV0BtM8CzFYrPsczOPV9dGkHC+pR6uR
FtA3ott6ytNm1tvyefFhd6mLTg9NNMl/2Uw1Gwgc7gbqJ8hqecsVj/DOJbwMAuWTv1R0Zj/Td00c
z91DkjoyHrWCnTFzTDk0YXDVXSe19kIkx6x00a7eNOu8xWvZ2WCc1ujmayi0es1/MmMbMJ82J4fV
JziJ406NvvWYe/scOfIn6zWn/hfGHaarrluVnVFe7qbdLScIEv7/w9SwdtjApBCuxikEcEXIx6Kb
M7LOAB3daqiMsgGkspmOIA4BTj7jDWtTulvZqyI5Dy7/isClduKqHcfDVKi37xH9NNbXEI28imyU
sOHeRIthq3zNmAcb2vLIEL6SeT+MmS0EuKI/yy47FXd4C0Tq0z42MFMhmSZoxDh84uTHqpdm+FRq
q0OYOq0WUoVl/OzA1MV0iDK296t8Un0Bvz5Gld/qQNc5RR5RMdF5pkDDHrlL32NcbcW+fjFdjiAm
uMTa6WybojbPhzeSmZmxUN/DYo01vyv60ylUD8C5sQIv2+6AnQgKv2iH3QDHbqVLJQ2YtsNDlPT6
+RQyMyh74NgazHkGyAbSEas0FNBEiengMluZVMw2iCKLbk34xpCOmyvkDlRoeW/nMuw+YEiY69pF
y25AV51kuJMxZdM8EHrO9mbi7FAqC2wQNreNSWNX5dNz2vbnzzYqzDyr4bvJUyMvFZSH0RGQhs26
4anPpGTddSB7sEVOvdLrprSc+YT1ZGO9xpwE3YOD9k62bMugu9KakFnkoFOunyu4ALlWPRzalKbX
x6bhgf7T2PqUwo5UTrP8ciaO0ti4i3vCme1JQOsu/bLRy29TviyJlUasbSUgSbShi5iwT7PyV4o+
17UFuPJKgORyRxbTPPCHiZbBFG6zb5pzWdCKvxnIDdZQLLsX0PSQ0ysrg1iXM/onJj+QHbonCp/e
Zgi5dIsG/ZDJrLrT6tKVXp0646ppHL7i8SU8RnwtXjH7VIIQj3e2SJ74Fqy0EGwmsTKwTQFMlDLe
WPmRK3yuQsCLwJIdwngUE5GUdS8/c8HELwr7ZmHlBg3L8Sm+PKm2JXWc0nYYQQ/tpRC8RnT/0jzv
rAEFaWgzcc8VB23aSKKnmJNsTwd4vYhaUiP38FNKphcefj2zmmnMFHdHHfGlJkbaPF4ECNm8+TnX
Iato6RY2nbTlbn5V4t2dacQevpqJPFZbqruvfjVTwaBEtsVHczXKJc/DRy6V8Ct6IDhWKvcRm2x8
QFJQDuooCZYZkqZcjs5Ynsvv6oNKr7nKRRM5QkD/SmCF1iPtikiWppj4IHaX6lIxnomyKD2vO9Y1
xqWLlFnv/0eesAuEXxPjrc5Hnq7kQFEh56L9vZeBqRieely4z7tbTaEzbH33jIhzeJFE9vQXCqFP
3wf42yCmFCCsM9UVD/ZD6vD+1cADH/hY5OmU0o53G1npHDo2JZV8fRg35tczkIVDAyEdiN1CeNF0
rlb1DpxZdLiPmyKXzWdM0DYVGJpnFDIWOX3AwGQGRCDYBUApzJ9ApavprnUAPPMH0XR/sJJqghXq
SNx+wxg41aBQg5BrKoH1CbXImwSFRSvOv5t4/eHux7MSzqPgR/EBsXbvWFH9PPK24GhUKvFePOwp
ISLSgrrwsV+mud3VVACOP7vyKuB0rS/AHQSPw8Re9HuoyVaPSPQUnnk47uftKDy+3g8fkH5NyRYj
Cfc4WV2T5c2LPf9cWElT4djMKuzggIHpMj+H7qmiXF8wu5gRsqn+1Ffa38dIkYqt1npl2kbnsWVq
kwwZg6lnBqkL9jD/2hYk8AqRxvOU7VviacNAhe95HflxtCV0VZxK3aNLkgz8PWAWmcbFS/+IcAaz
9Honp5EuCMrHFe0UNmiR0zPNQoArYfQrI3L/5pk+ofKkixaBpj1ACjyt0FS5Ox0y61yT3hylTNuY
fe2sX4sqUgepSX6nftM1Ewv8fzhQ6H1KMoNNr51Vt6HXS9QPsGhfUOiUBlYb7OjtDAScvZQ2QZY1
w0XulE3vHxD7/LVh2aLOod3MnMcbtXDL1IBrTbjVrIjrA8IizO6VwrMeQZnIgn1HGa27bz0QdPpX
OKJngMXxk/VJqejcXWl9hGWW/p70GiXsUxlZuDZxlqy+EoS9+F76iHERZGe1L3+KxZJk19+g+USG
SHY5mpZYe/Eataml747tyZIhDWT4WGIS96Q68K++6ZLWSqI9Pj257yYo2O4RDOnCM4VPZuZS4PQd
y0p0MizDOw9saInN6+wY2Oh6FiRgK2j/04dMzjFAJgIDZTgAQvmh2czhU/1C3/W9TVFtOp81B0zm
7F/8jEcDot7kxneh/LwzvilA6CTEto+j51ocjX2SKjvU1AFN4tPArjoU9hCFoJ94014qaY9g8l2L
RdZWRSA40jYlq8/2LrSN/tztlhquVwSO4F9vb0WxlYwGMsOMJ7D54I+nh6vSnXFphhkOBzvaA/+a
BohR1phhd8+mHimGIpOcxBh4XcEmtnaAhf448lx8hT5aRSI3r/pERUOU184xkIKmBy9Tt4AI6+S4
VZGD465d2zX8DTL9Y/LahrQeo3+baLBD31OZPl+5izGBhSpRPaXTfagt8nQiStgIXoUcYArbNnFP
LZjf/YlK0aEJBq5iVgmvdbeYTih8v/gTNuoj8UydzM0xTelxrF2RJaeePl7hpmsEJs0uk3cwz2LC
WqXJGvTqtWch4a9LLu5ZqxkmW9h0UiALEGgzOjNVdDevibDubCDNKRz9vSdCXtDUsoo979ehvPPU
SnZSFo3I2Vn+PnsdT9pXN5F6yNvml5QckWGmYDzVRU0vAl8RIdYryCQPqSwEFkXhC22EcfiPQN9u
pc6DQKWX3aOTsEJGL7dXkVtwhNnPzwTHuz/v9OO70oi45wpk/LAopxYPWlIpog7gyDcduEq+Xzyc
ngR5heGt7KOoX4M2r9G82XjNzX5pa7MlAiIM8tS440s1Wlt0/Iuuw5WZvtKEWb2FdzytvCOxB11W
YI/5cUiciehi0R1eWGO4pxGfF3JX/B522eiGrGxKV+KzyDTBZXrDGQlZ7TpdwleTFiIKeNqMe8kI
NLph8ofsIqMuQewJ13TndRF4jDbUqFSgWSCvTTyYfCZoyqj/dDLtzHtUWkAIP5yRRsdQaiSjMn+5
9NZrF/Gjwbxu1D7nQOVFTn79z0sZlobmqKuEpIibjtaCBRoTYWVHF7+Doasml76Ny0LBn5QQ2VnQ
IacnWEEmlkkWhfnzEMPDFT9iClkSZTcFQGh+BhurrRl0ugawfYnXlao1Vw3Bq+lGj1736RkXRxtK
vz5Ghw5cs3lfn85SQZv98Oa/Ld/CG3YT2I3N0ov3Tj2A6MKshrs3eC6E2lUh1X/WPRtffgXoJAjR
NrfJnb8hSF5Yxuei/8ZMUUh/w5LafxT7D243ZcbH2WkfXd/cufHtbS1RHAeHabBlTRGYL7lhxLry
/XcOhKracq/7zCFOOraJH9bbIBk/seeamiLIwo57eaGZVDC4GiOiULX627lfadlgTrMFC3AKzfaB
GysNoFpGo9WHiSMXMu1KWe/cS5xiQ35JGlMwADeZMfk4TziJAC7tINcGqrHA8pOtbrhVTKGZNrbv
iZTbB3nfQH8+QWWIJSq1md3vmTmfUwpxaQgHefZfXhkS+kvMN0K8XH756BOHnaJlnESFlxkTOhj7
vGiXeHn/BZ1Cbh+eEh2m4REdqy2xccb/91rmllmip3m+UY8LuRO1HB8f2WpeTfvSft5dj5/na92k
kDXJuCkApA+/ByN74zx17wxaFQzo4wL7jGRh7ef9EWm4aU+hW8DyAjroBdYiLgDq4MMJqhB9YYWM
BRonjeZAt9QtnSYNvlIKZAEzRToaT19rhjuavLVzMObXzVovKqrPXtpxFChIcmrHngpLdJnFb2Zc
pf5fuHMkfKlgKXUrzz06UayGezoZVdcUmoL67ZGnpgjlDd7WcOkI4tJPQc2rQd53tr2qxm54R+Sp
/8ngLRfRdI3JfHG0tAVZrnZGLw3eZZEe6qCo2Hyn90S+CfzhDBpeqNtartTC5ZI/V1zl8Zaovyu9
QiwVGSNsRqUvmc+YdsuHnP6E+ZaIi9oQtqGbc+BTPx0gHrSIMiGf8QNm1eq8Gou7zfNtBRBwvSpO
Ht8ou3mc0B6C8qfTQmUb1kXk+KfJnSpdXAlMtxKta9wALz3hdvkZFSTTKBQE/dITS9xvgeJ9q3PN
xxmp4yePdJWRw047YMRYnYf/P0ccxFSJnYlgQP1/pqzWekiTq6rJgok48hf2qNF7gThtwM7gy74a
v8s7jtPQKysJzrRPSwY8SVZa3n78P4ZNuLwirlh8xhfyWFqH5eR/OL7PbTM8sjehKh6hday5K6fR
0SU9cbHLvYWxlLbj/Lpm3hglRgcCztykp0SQOqMR4Dg3D9aBLhNo2Mi883VqGCqSsAQKK2MqO7Vk
KfrYStybfW+md4SwKdwyEbgQf9dTnOcesQ1c77iSeKDakaRsFkgs9PRQCzhn4ScCO8KhktpZFAuI
xgeX4oZbyhlyvdK6VGJWQr0W/Ieu/ipaEyKD24M330/hzlxRz+IHqhiR1yAbVzSFgdYati4uvQ8B
HTZ5nWY9tH7NEOb6lqHnrhaT8D226TErHvSvGaSdhZz2/lXVYsC7b0owD0U1la2Gr75SHHsArvBP
md0fa1v3WH7hmR+dMopDBxsDxPtI6qqamX2A96/tlmcn8XHdWyC0UVVArBDSQw0Kz3m0b+BEvlMv
W+Vq8mOnSbd6bvfsmuFonBW2741utDVMyU58FV9Zf5ctdpRKZNMK9Qz/Wpd/JP7l5dP6zQT+te+z
lCS9nd/RzKu+fpEk3V+LTfA4aXYmE6R9PZoEpSG/cgLnTsmVSC0Q8Hx+E05I8PrbWnI5HozypkHA
QRFWAnQmZustZXQSFYw+53Ayx8F7K7Q7pOHtlKrVVxl3752Tp8bTt83GosnUOg8UcJaSTKCHNWtA
LO0XY67xTdgI0uHOmN1JNw9c59YToDaYNYGCEX7EMty1FAlXqaoA54kiNlHBEjnCUCBwEmuixO2/
JbIyihp5NkcfMLJencxK9pqNTrKB2m6ICYCm8H2QSWCeMdzVnui1kZDvQv3D5V6+lP88OVXV3Ol4
K0T8Vh/DwX4EpvQUGdXBTxUylSqLyU6yRlSQfXV73QemMTZ+SgPkFsTTY0O4KMS7m6Sbe2O1Scka
887a8FYJNdYhGZBkjTvhS7nIxkiHEfJJ3ZuCqCftF3WWJaEkVC/rf2+hlU/PxG9L3NOxH43XS6BV
kB36GwFDnMwqadzyZRNlYEMB0f0t2DO0vpRH5DQzc/LhIcdeF7EXRcfOhUHsK7tBdO6Tz6No5efx
BcFVhmTNGVmOHiZCD9d094YAsE6s7nJSkWpj600izaebZoLKRMKcBE9Yv5Vd/MUozvYsKaj3Ym+B
yOH7R5Wq2QGL145cgIWKq0KTbItMMCqebm8cy5yNTfsAdvzNfzSU/CFHLyLa4Wuto2SZRoE+El+F
1RRPg/rQx1mtxYQagxFvozQKV8V54TKeAOO2/weEpZbV54G7agm5hP3E30WFvH+cARKVnPTWv4Pu
lZsqoUaB+7pPeJUZI6i0x0ATTmOB9V7/rcOOlKZyMkYKPFDq304tB2Cqz8OKXVBc87fjIXeK9Uk/
3kUJAmwfNu+vLLbKKFfUooU9N2EkMCPIl2WFvpSnDeqpmXObe5xq4JKvNd8WR5RRTZDgeKcTpton
9PtKof7pnwjdtTxsPHabbHDhSmlBhfbJUXgIfxJDFAgCM5qsPuiEwySMd4Vpy0mC8q7O4df6gQgA
T2+KoAUibLrX6z7TLSpZpzqSIg4wqLTbPY2PysNpdeRcCoKeiRs9IYANwvpx6SWRv5MNugzSeBIM
vJivtHbv7U8ermD0vjPoV9+FIveXKWBfchzUfk0o2SQV6ERDRDxKIXsyslDF8u49eE3WFo6wkrBZ
nyMnjaAq/sFImpGbFHkE8O5RBpOuruIVaAZk5JNU07YNqcCAMnu8nTZvhindzNwfzDVzubF4lMqq
qlPwAU2qaPdZBFJL2QKCwLJ3hpKVQt6EJZX9ibnFZCnF6avHQcpH6M48cLOnP5g/vYsNWqFkTw0A
VjOLbDP2Mevh0PFI/BxxBzj1IbyVkthwIMs/5g0azu/1xAk+EXRhZlImFYcD8P5mqd0gUTpZNgCt
1JRgLyJPX/12dJsgYRDgGvbTWUhuXjyJbrQhMoWpHW+8id0NWzQ1mOsF4zxk9t0iHulg/wqvt7PJ
XXBf/G/NZrFvKoPBJdWbSVJOfdgk2AaLHCphpwz7z+V7cijcEFH9ah7bLMvg7hl0LLu0qd7csbG3
L7KDnz3Ocpxn+gbwIhBKkkHGeLTOhwZlZKRGt6GZsCU42FdhZFHksUK5R++Md9aEPUZGsbN/mj4b
cvgo/dzRxlgAJ4rZKLHM17pSXjjVJNIWcSTjzjRjGgjXAkgEBt5S2xleN7wOgP6fayYOG/jsw2+c
lzmZWPFz8/pKd+7qOMmDwqxoMw/p9AzDxgOUjbEN9gkecBrQHsNVo+qUZ0Lgp12UFeP4+/Iv784a
j8+hFeMbG1mzcwP+jDCHKWXnaFvQLtu8WwlG7515eZvdiM3JbDyzaUYor0ySP4E2uSpfLOPJu7Ir
OEG00tsnQLIluuBxb+JqCm6oS88uGh9cACjPSKB/R4Q4ikfmhxXQ6nlXHVghZVZ6v6lAd0QyKg/o
hlF/Bps9Hi6TZSO81XoEPUYuRAlzMUoRiKxvp83q8O9YN+7B7+smoydPyTkc+KcbRsandIiPm7uV
QJGti2Riseu6w19i6PAFnRyJAV8gQSTdYHYfsnEwnwKpDu9A390OsawRictyR0NUYzy3mwtDMX77
02oVwSlMXABSWFAkmathlF+hXvC+9ESiiA0RVY+qZ2SqNuemUwyqzNJQkaXcRSZoghr6EQtNzSSt
BXpqu403I3jhkUBzgO+2bG8JGKKaikV2U2or2np7TD7SQsraPqlhaQK5IxlG2qzIVBljAD6bR7ko
c9pn3og40eryWLSxpcThAEG2ocMT1KJnbfvEDU5Jb8l7i9dSacloFzIUoLs8WXNdXK6KaQ9p6b3y
iVK8CAACWhR51KDNhnTKoMAZt4SEycpkSoRqtLqYJY6j3TEdWjQr5ppgSF7G7BgG7hEWAxODSa4O
17N8ILGD4CJpIwXh5I1f/zYs03oRdPklACnHJ4MdXjcYYx4CqmSY9Ny3e1snW2I2wsqKDZ8IGQf+
lKrIlQU6f8X2Elybkr29DiDPAgA3KRsO2FQTDMcsaw0E3cMCpYTe6vKNN3bsnKnO1iP11U4VQlXD
780PMcnKMthPuF80/Z4E399ltYKZMDSHwDKGOT7rZkQV5wCVQsDX/amuOdxdmefXcMIbkQ+1Qic3
JQUjVe6CpKla6nBgPHrDXB2b+aHIJR5AkRaazmS1SohQM1faQVfYooCVYF0eooDsebt8CH9KjCwE
rKLTG2Lh3HY4GGUlhtxsO65bqxzOq4jmhlQSOTPVYGY+SHFo9DHx7WJqXvP4fd50gz3MEluzwMrS
y04qQSqKAQ09lv0a4le+PuQIMSUYQiqAfSfyoyXMSFxMX9gbbiahtItNPZYZfhRptzgy9aIInTQW
bU52PoHVnjuha6KB+4eZ/OovHsBPngM0vQ66U7H+JyCgibxw4MALiMY+2Jp2yZtembKAej1NaeD8
eWjuQTn+aiTs/By8m64qcT2DxpcB4TTPwVhwS350PmxgFsOW8bYI2EJEiP2nLB1pHljw/KyRXVtq
fH0mloc4Y70UyOWF6drKSLOhACBTbOag3JmxAzM0Bg54ljecB8onWXTPSOyCNDUZwbmeLlvPwtO5
UcDtkfImUoGnuyGiEJHrHC85K/FyFDg+pIZKWz1u6ztPVP25a3riRdG6oxWHmvMxzNPhjEb6oZmi
nyyT462p8l4YaH4DaReULHfmIlI+qbpVoIaOOdvbaWm9AjTY31/8llyA8BmQC55UujNM7h49VayY
zLPOr2lrDSLAglbx842Wp+O+/Oa5HkasfcRZr79H9jiS9EyG85LbTKg284nBSroZXChGX4rJTK1D
TzgQs9j5MvhIavePdQGJh37Hpj7r0EoEVMySIVkjzmVMQNZxgU6NP5gYBuqlEgXDjvKKema5j4hs
Wc8jyX35n3STgICrss6H4Lo8Ox06xaUjirDprUeXezdZxdh70pYK9bXrKY167l7WdFP5taTtuU08
PBIWxJrL92goUsv+OTz61rTacj2chgGm5WYwMZ00bD3mAFCSAiEdgfOEryN2YPYMnhN1RbOmO+AY
l15pHS6K8CzrCzPicJhh1Ff0yamJ+MhHVVHn37meNYszFjn+oWAOlsm7d5Xcwv52z3Mj3PqVjxzB
u21+NF6nOGxd4QUkrQzrGoS0xuV5RQQYqMo+rdivwv0kESoLpX/2vNDDRyyGmFkU2WLVkuRqRqMP
yAl3uflkwL2/4LtqZAXHdYeWh8D7NZrEE61m0S1R5UhVw82ocZajMP7TiUb2ETw8WlttueCRbpC2
0i/yzmnPWCiu8GjE57OAGqPfAQJ54sGzWZXatqm5/EefmdmUPqcXeIuLjCsZlD3C1AXG8sOxhgKT
aKjVcOnRRCAAx26Z/7mLFp4+memCMVgxlXxqHaVG55fhJmrRsYSbFM9FVWkvzepJAfQ0qw/1LJvs
z95O1TDo/9FQUXQi4z2NlWvp3W+2EM1YAZQ4zLokzRbxPMNyJlWDnlbVRnNZlbQTNM0OJhjDsN+9
8pb035G8ebRXz36yqKfSbpE+mZkkd3IwfIf5ZrpJ4G+Ugh+nj4uGJ3gTX1o15hSmNAH4V4vjKBF/
kYbvKwrC2EHVu+k6cVTQyHWhDkCaJDRgvqIZ2hNukIqf1ROc4Rcj7WO+fs7WujkuMvuPN09BFHD1
RdQoPrtysRxICWZi5BizZcu297Ikpg1SJwAxGDHJcOIchuf2Lu6MXCgGoxIbCIPt08VFCPc/C2Xu
YCY1KoZLjg/5V0LsrrIBvxCkc0I5dEMREAUVxT5AGtCN5Mmz+jW8JkEfXT0Ikq7aXxaZ4yQxvLs4
Vf0EBFTTxgdZuIEW5bVxGXQlpcOGtCz76QX6iQSWLL2XZBTz3uC/IX041SpP9zTTHHv1K4+1EtDw
21Ygo/1Bd0t8c8aAUzG2N4xDLL/ifoZIIc5g5TAFSQEabLSQF7iJxCMpTHf+uRqwybvC1QH0+cKY
nSGiyzy7dE7ozqB4+EgiareburrHguFuo+cjgddiIyMV4CLikZrq4A8zpo/8pgG9s7n6d01/NnUS
TEgedSgMt5lcpPUnNLVs4hztqNHUQm5tmT0FhCaGkna04JOQeB7veLpYURa5/aZ+ndLV+FKELPF7
hk5251edbREpVjTxGpjYvljuBE1EzO0aJ8x/yUVlnjM0++rktecAtRYE1agRPKe28ERaH7frBnJU
fvlo93cklMxs/Tt9jwMG9wDHGjMrKMqS3q67mFE2NouUzEbnO1l3pwhNAssC6WkYmTs2SGLJOe/N
gWmYsiRICsHzboSK4HGHz0rKMRRD9Wlkum34ucr4MJyPqeeyCx757rnluXgUDPJGMp//Vahm4ukv
Itfh2K3QtZKzv2NvOCc/lNuaqpSBQ8b2axGK4ncw6hO+/AsXXkn1yZPgkQYQxJr2YyNmNIPKwZ76
lVHQKzOuvwbnXin4BqF/DqQt72Qm23yS3JWRFSZKBzeUVKBA6f6IsYhQlaGTc+qprM5ow/w/G/Vv
Q38tjcgjwZgQ47YV2pvoKTC4w37vulASkfhieT6J9PEJvIZU6wTSeYCOLANUPWlaevF/JRE/S0JS
f8uArCljCamZmXjrweSSoZQjL9tNsAp8CezxmOpoTlRgbJ8vjg3PwaTiVwimF0TckI5z3Hcxc+e3
s6sqPwqOPqog+KwzoGEi5cxlh383zdJycbCLJO9YxPCfT/HlVmYXkzC3eCFQSMSeoW0PqrduMtVv
J8NtKzA7jAovtJlKm4BWY4AHYPmpa0mgE14haBzBKv89A3WWIkJ8rTU4sgTteND+wxHMTe1pSh25
fKimF5d3txJ3J71MZG/60qTfPxhZSBQz5BfcFxTBPKxTe/ZP7c4lQ9ypuEdOWqZvxbK3zbf+O5BH
xLQeA8uLOfUjKIvbys9rhYzEZ4qUzzsToO24kN7a4FXftKsU2LYcyqpCShvu2bAWt3piyWSaLdMd
X+tOKuuCMRhcNoAJ8Zekfv8ZqKzsbjqMC73/9+nlN0lLSB5J0MXb5K8qKAuUuRwydM5fNopmg8lB
JMgNmZ0cqFbDQnJQ7VWs74qFWEm8MZJwKSlCz8+Ux7rl1B7qu9WPQW7igD/O0VAEWwzmCMivCrNm
ZizeU0qVZR8WKlCOrO/+HJjbeCjNgT/JW7M0bD8p4legt0NrPleWViBam4DLkzgOKhKIPZaGGkfJ
qHBj5RIgSHoq1AwgANlUFnBRhsd9PY7jnygmzZqbH8Ihmnsaoga2s+DGwqVLC5fDT5xXWu5XrS13
JsdE9uTiErpiS/0vw8nL2k1bsQ+nNK6WaX7aLuZIByXpyG6kdJVqqvoyg/B6rtduqitsX6sQ4bw+
kyeJqN3Z/pX9SHwm56X1Pe48vOC4ZMBVRrSzfdbvZhM74HsopA3BAeQ9q7Fl63ADrGTIjVIUiiYm
jlVY7ZdVIa3udBdrlXOXhLnJAiaIRbY7c5NhEob8P2CZa1OWJdjWrDMFXcPvgbBWaCTN4TMcCZ0+
0VId/aaTBmyHWCgUDYJDxA5RPCp4QcRNxb7sQ6QT9eYWYu6ip8LfRWa+a90iFEUk+NjGPAEJ+drY
O3/W1pJjT5s0V7lw5drzEL3SqUaHzNWXfSdSzdPECbFP5amCxUaZQlyXe4mzg5xQK2PDMfs2vDUU
7f3/GJWJn0DPwWtM4ma+7oXeH1PpgQUpNdyY5UoFtA3foSUnDBnxXF/jELw4U3z0/nsnvxEXBv7u
QKj95GmKbBTpw7LCcbnnoKoi7rME3RuyNHttI2EowUQjLn+6qE8QpahkYvgvRVQqzECMkw5P18ZB
p5D2C2CoDDVQSe09aTXAc6oGM2VkzY5sY4O00XcNxPwhQjMAz39H9J51lyEd4aDOpZBx4vip3W5r
gL8RGS49DzegwvVJJXzsvO5Funv8a/QSi7HXlfzyhqQ314CGpHXG8+mvGgLTC3zgWrZhNydOqf0I
KO2KkiabW4V6vgnPbfFSL9Tt2B71Pn6qWCqRTmsjjFAgQMaAtMfy4gXg7NlHjSDsao6UwyQn7xBL
/uRhDuCLpZpLPlqQFIvHk/9P+m+q7OZGSkmRX+4n3BkjPDrowRg63tNZ3jWDD7PzymuszlBYSTAX
QP22S4TDCzCysIFN734/3sFrpHNGjOpWT8bkf+DAMKQAJAEXyxQMeG5ZBow/sIfw9j/JjjGjzOwW
nr6oUmx53FIYIQTdgfvVGJH+8pce9Qjvi8tB4TAlgiFG5v2oWz+hfKKyVMriJQQfxGYde+/LjT4t
/Cnfoi85aHBGl6pvyNeRgLGdpSm6VYpG8kgsOkhjGK5SIpE5O8xcKC1w4HIeNosRPSfDwzcMDcI2
ZjoBnmZf/AdeV6SxfC+3KqNKl4l5sg7CD6/ChdJGLyJ/llCbn1DrDJGHQgRlEAztgdsVkoSrDnCl
MB8bMjw+jQDsRV/UQyPkKVtxN185ho70AkynX+nIcTT8OFawxdmW/f1vMole9g43US8Dox4NO0ki
N4gYnffLhnka0escsPftQwpZv67FMaqkq9kpKTKweovtCtZVTM3d5BnUXHt537ovyKI63FOxizDI
q4EC4YUcDOO47UUG1cbEMKyS9CGaO5UFbyaCa0IIeSTifeXlD34VFFTjPlHRT23xqSafKaNXNHBL
uVEeQE8Ha4+cGi3DH3y7dligxYHvZcme3frCBcnrHxkwxn5n+ZUXBO8XYlDj/eSKJyaYGZdj4TzD
3siNoFZldEQTbRrR1K2Sz2sCjv6MrEmddbIECkk1r1OiyoIFRGNlTAfLSELC7LTIw36JHWdb2Yft
91oKp6DcvFycnrAYtuwcR5QPlykiccD7o4RDCYNiWI33r2xuu0hkEBVDKOYzxvRFjjSB1ck9wr4G
JwLLaEqaZefQEuIEjwlzNgvgTzO/PrM3aeiG3sq7/bQcYEkJUFhbrn6OYE4risvVfINTjxg8jyds
jVhHqvNr1UkpQpuTaPBzhdcVvj4mQZATH3paGtOuW8ucu00NyWIp/zM3LiVrUxdCRtUF65XigNjD
HUA6/87xeZsSXeYjuA4pcy5dPQcMW2nkFHmAiOacbhqkspOI6Ndoo4U8THXKLoMzmA9Zlkmu9Wpx
5wY+eYTSjOf6UJTkdXBK62nPOmYueVn9deirQyqsYI03O3yYD61rYp8C0vVhjO/GgA6u+iTvLdtF
0l0pvUyD0pNvtA4gJObCPbup9TuurssXj2Eg2IjKrsS22N+n/Somroy+vguKtsgIS0dIIKzh+dTK
44dvo/xPf7QXMxKmeadB2wAW/dS9geqjFQbDGXw2DvYvdeGpSdAWwxPvy2hzo9j1GB4Wad8forAQ
FXQvW0rYZHg9XVHgKbYa9eNkuQPcgt6QVtWMfFWMcueY5npiKKJym9A80vdp2doQI03/IaMXECmA
jsITJ7tK8JA9rwBirM0DGF1stphqXVY35RTwkHEgvQcMLTSeN4qZUv0L33A1is0Qebf5QiZvnbR9
SRAcASIv9MdjwwPpfAdI3zyYpN9fz0SsBbSc+lLDcUkm6VQdJmzI8bqxAYSwkz5arRKFIE8QLZt4
2mNlu7w3Io0JtavaRju5SgoMcbXIgmtSFNF2AjP6zk8iCklyNSb0tW5vHG+DoJ5DOcKY+axmn3+g
z6+I9tN0/lOKbO/nCM9Gp1iIiBJtbDAYtbCQKc+F6uC8GWuh/cO0KyZoO7I84DUgI6SoGvlw9J2F
pj+MhsMgW49NXjMUw3o0ECCvhsZXLTSWTGp4bGSTFJMxAwf6SJD9wctpfTjbFVNJtdmnlfaRsa0H
Kp93O/pKorjOaCfgXrMQl4JzUuCqhwOESz0ugGy6d3FsCzZFyk1xB6Ujm1rPzxa2fDjwptpHYlsE
vhqm9Xfq5IyKJDDfa/3x9ky6sccxpuLrzYwSDyHwb6xAs946wjOQp6j8i9ksN0nDvHpXnPwgOqaN
O6VuQpVLKq4+BTTgt5h6ECtaxQc5YL6fBTTIPa0VWcosQzmms39tD7hLwTjJyTN6yIxAbHAD23MZ
ph/zQj2sPEQkwF4VGF2VGPVB6k0eVgoX12ciq0e0UNFhMs1xApAxdsb/OAlPaTPnED/gFwZG4TvJ
Ndj/s/MZmYTWGe0xiSBgN29tF291rKZd7k5urk4JbzYNwcVsmnl9jD+kuTNzh9uahpTm5SnqrlaD
sB9uAiqurtVEf+t9hJCCv59hhw248kGkfDXNpYIPC5pU/s9lxJ1ItIsCeDyCDq/z7C0QGF+ti1Js
hMckF/EZhSECZ4XlzivlQdi0Qu+Nl+1zyzuV+sb9qPqO0cCfqyfLeDM3HRxc1fFEyzVigC1UW/wk
jH9IWY2yvWaDQO5NvEnKCEgJU4M+q/fH7s6y11zjVL0RnoW+2qht2nhgjJ7HcriCk1LCe0j6SaW5
9AoIgmThrGYl4Gdnyea1iUqrvR/sZsa+4Gfg6xmnk23+Z58Q88lOKtYQyekjw7fUBYY9GQUgMevP
NU+dSt7Jo/3dP5VpxZO9/v6Hn70abHzV3Jb0uOTNHdijydyXvrCZFn7WcrI3s33kUbq77FdEjigF
XtVO1sd5YyOQPB+mZVtuhZPtKLBffA+PFSoU/7xpgxnF+RuWCzqKYmjahBuQPivPvmrsS8NR9uxy
mSiDrLhoUzazmgNXfu6hdOB53JPvtEJPAXshvk9TJcg3ON+tCnGm94Z6lia3w1tUfH+AQb+x9Xb6
N/qPzo6vdzZJpIWI0RX00oA6gG292v4rG06vLwMWa5h+U0eZR7h9hmG1ToD9i9fWmqtmE1778nVJ
SyKu0KLBMxfPnUwUuHIQDMcNbUUSt77tMIHm1d7oiXljMnJuBGZhmZRQzwbC4v1DGBlTE+dCHgLc
Im4i1H+Z8TL9oatgB/JkUfQrouf5dNy1aBT056SpR+hFR9gi9kAf2Q8xbuPe5V4e59rb1ByEm9Hh
li9fjNoTNLAKGQwO2YXCr7GN8JMvkuC6Kb0mzpKEI8SPHbb9/+oir4mji1J6I2YC04XMe1i7G41/
8M+Ag+gvM+BrvxFQ4HGtcqUe7ZFmi7IlSHMQ1bF2IXRNE5iWrzPIMDApmGDJg+Nh6A+ScCaGhcA/
B8T2dd5uNkyIyCDa17HYPWUfYux2b1SXhpGlA9twR5a0/6sMK4597riRVExbjXiyUTmnXgpAQ7Zr
jDJh5OPYgiWrZU7AHArv1fp7mUUk7UIWSgBLGzIUlu9Xv7xwmff/B2U6cYu1mPGuTYbtXl6kFMMx
R+VsoWsLgjZPg9L2ruJjIUfiBBCgNU10NsJn2Fd17BukO1qREKCAod3j76NqcObr7zvzPstSt7MK
avQA7WGQPlyRynq1ZQVyuZtAqKCZFplWR8brl4kqpmrfc3dC/9Urt06NJoN1yxCzYa3AETbPg60i
Ggyu121pFI79PveN2HnXcZtmI+mYRCvZf8KmIKkyHffrSJWvNjdc6DJhrg5jvYBvd+ftnfZwr4e5
lk+Iv6wdey/YHupU8yLxgS7stsu/9DxnPF8a69IkfyDRbTNAKSLqgFYm7Hi2Aax99z2K/R85o7cp
v8vZNmcPtnoh7xXoLuA6ePAsMtLI5wX6wY5IZXhUci1xPIIyFOTb6FHOpkboT1VH/8xYHn/y2YL1
7LVGACmGxawVeEWJOkQEGqE0sLXoSfjIO65+Ck9ldRm9QrzBqCHh2QR5DrleHAX7QNirZLLffnp2
yZ3AEWHaV2uDM3UmfKaIp3nn5x6M36DrZ3vUeL+a8GK/9POqb4bb8vSJWj3Sx2F+nnDhK8CFuOb4
q57S1w3Vq1Y/BhKKuqED9C/zHve35VEKU/WzXpNWxK/RARDIGGe7Kib6rU5upPdH7l4/k61eYAw3
20P4nn6XDHBA3FDi+qamboVvMIgFYFCza3UBQXmkpT+p1QOZJxt8009ph2k0T4s035kYh5EQ2NTw
NNEGRxqH97LL/bL92a5CIEBIOeWIUUoaSbjWHDKjaMdHjMd4VT1EG91rVgA71ELNaqWm+4XMTFFV
XlmECswd0BckBXimP2RG+ZpnZYxLEMTJkryQdPumC1eI5Xz+BBoFFoZSFFraLPrQKPSmN3s7SZXM
q56c+HCz/tKjNHAzO0EaArvwL+pglrb9bCKgIhW6cVw4UMDrUyRy6GBXiBOdqEzhK0B+rSoJMYnw
9tnMPp0b8uFdnJpomiKpo1/3D8pOvJyQo8w3VPeWq+F4fHBPQqgmOp+eABsvJudWRxaMCQdBWVNb
y8A2A9JNE9tMtaiCLgykZAFYkoyaeY5wYWjYIv9OUqxYigju9MDoDHkBrxKT5mEC7bR1h6Edyt8O
y4smmvaq36/zSkj/5UBRSVdDDWHe2teypaBhZQZtqg1drvBKlbrEqby9DY1ejbz8ikJX16Xsco3C
MHKzZYm8LWlUyGAvk776UwvbfJO7hkUozjzDIN/aZj8kGHKHzDT/3W2KshWNghlEemQocN1dVZ0R
gCSHqmOWApCw+UJImexHxV2fkJAgBJ2oyZXZiU9E6CERk9ceF8Ip0YbzKGQNsdYqZcQGg1xlc6al
omNxYlUWe44Yvblw3WUbFxq+Pd/PAq116yfajLWmpN/6FIx5gk0iyfThGX3ql5WryEz1NGA6Ch6M
SMKSPuE1/Oeo29uTvHCKTT5E1aJSCnCpARfpHsNUFCNcBb6Xjytjn9SKgR0GZkkiK/3e6V3zrr2C
LGaPmbI/dEx2fJfAHuV7mQ2Yc5hHlVOCr+c/9YUHC/JWfgCsb2p5J8LzIV2q86Me73A3vHOEegiC
MxAZDVHTeaVCdXkdMUfiK+kcm7n64MR2wOGiEHNGo5XaguQLv1wdJ6YJGyZ7Q7UdRUA6d18SV1/p
+3pSEI0VoPaybt3ii8Kax5Sh7wkfE91u/Swi8cNmSqwMMYOHcG0jIXTwUIIp+AoH8CI3lDpzqIB0
/ZUEgqD6ZHZ6FpGm2aL6yPRhqVdh3AXxHyubiGVygwYvUrsfCwNrsyCztusN2K4fNpHUvch/0fyA
b3Eg8Ww9MIGjppUvOUOAdHFRmbvqZ5OVOketL9POwga1DqYn9kl0CZR+kkuwHc5kmCY23P+MCHuF
pwrCiGv4m4mJRPJx9ayKXF0g5Vp+iLh9dym8pBuaGT+HzMB6Qd4CWCBoIycs/ovbTzs6F+Hz/MHW
hOUxYARkpG48RrzUEtueWmajbbk5khxRhYkVYndfOYr3MmfR5kmqjhaNRYTv67NFDCCiQOpvsgq5
ZUglxC14fmFMpLXBQOa04crXUFMSzO07aaMLZtvFHcZKWzlvwiPHltMzpt25dQ/XlMMrcF0nNHOe
wVt2bV59z5MIqCuqlV9/JZ4o5J2p+kRC51dBQA6VsGDixT5QLeCR4HU/C13TokzmuWp8x2jUEIUZ
HYqJyqXOduqRjE4dNRlSU6EY/hhxYXnvvzvzRHhuFnHPayjqpsQEzUKdfb1UOydAkK6lgwmMHdr1
KJIEzcHoBjEdLBb90Nd5uKPDEIoVoSrnjVcvwTPw8L+VKwyTrJIxFxipYnBsckucUn8wqYcLWBwl
3rUlLRlvLmB8oculkkq7BwGs36WGn3MFpJcdD0BGklYbX8XQHf/UwJh4exB8YpRqyKDtsmhIYaNn
3bnHckQ4T/9HXHXRpNVjMgI6UvEcPvjIaUtjX27sKZBRz+G6hFiEk1bSuuHAII1ZGotz+AnMriwQ
wJazKNCEm3QeAlBr1FoPse0J8q7f0rz+Q/7zf/D9fGiXtkdAjNl22naST+eXaUERdrCxckcefrVk
jqO5+NvcS4zSfv+8sgVvTUQWwUkBqaGftDHdB7pgXnf98XAtFakyBuqKVQNV7rYx4fByKzWOuisp
3J2rRjJW+SJmIUjqo66iC6RCgAyfI5hcwyg9wGFIJQJKHYO+ZczRQubTZs57UAT/RgoTvZcXIWWX
ekCsyKvy4p4BTzcHO9BIyI001KJj5hXqfeMYGoxz9QPkb+9/hb0eHWdftYJLY9GTB6pvUZErFhcE
Z9+cVMiH+x6t0ngNz79mPV+qVNIk6Cyga+2cIYUHdy85rhn2qBSaKREL8or3mWJLU8bk9Ahz5Kvr
Z6YSNHYT7egeQUBMrPnL7sVTaiJa2DtX50eSRF6l/r/SR9M7+yOXhcTip4yfb0/ewKc8ZXE6dmle
IbnqKVcttJlZntWQFAuSRxmDjsJoI60tEgjoyz54cSY2CccrJ4xvJ2Jg4tsubAsjo7AVwXFl+KsH
6QjziKYAWzit8oDGLL/a4z4RIOGdusowLrXeIP2P1rE8KVsdNGh6I/hEzCPzmEmgWekCzVJt0FAD
7KhXvIlpNHGhSIU5OI5eb/DWKYpZOOkb7YYm5KWwRLOjDl02GwHp8sx3Ucows/FPiC1T2Uynte5L
h3M8TeO/rj9qxRTFo2cynnyeTNQevaSRi/srReZvquxPXCro7DqlEzylZ6levJtcuvCE7A+9W78Z
pwnNObFIqn6kM+B98mp0RuhNcRuZZfnFRpKXVwnmHVBq40c8aAYlltgUS7TxM2BDB+WkJlSIoa1d
+mCAwBsmVZpHZ1RU6HC27je0Wri4d5VNxynDEMThX8hOysw/DY02Hwe6/dgamd8akFwebYm8HFHx
AapgBot8c5AzbxfCkR0t+Xo3hAPCicUJ/4MKl42k96V5Oj+VmojHKDzlo6kz8SmQ2PyZkOhIzJII
63WQKGpSBUd8HRixnsM3dBoW/6hzkWf4gwzr2U0EsdAwn/BVWpP5OVXEm1RyuhgtS+aesueX0ps1
UZXRe3mpIR8oX5psP6D+jvObC0+lFlUdRNd5K6FuU7h0hwnxadr8+DyZW0wzC8dCQK08I3XTSEM+
ZrR3yOa3Om/OlxSIhJkKvYMIQFcv5v1j7Ba3fytX68u2KVKh/D0/6Ne3AiRpHvcZu8fVZgnSsfQC
nnQm86H7MTrgmjkkjrNDXbBfV6xdvuQy7hHtOYKDkmqQ4mrDgMfVA0UyQNYDzkoE2aa8Ycjs7Kej
NPEkpsr+IGl+FuRaVB1rIuEvaKaLygcF0RhyHd/qaAqrPe7hpFs51hGCyStshvjh0k4SEGyknG4Y
Br8GfHqWmPM5rcwzhPDRkuxiau+kHPfvDfWcbwRucZhG4NoVOVqRwwJhPegwIUOho7XmeAFqfYnj
RkgT2thOOL1tln2ZYyJoASe6MT4IX2jCf8CxUSoKnQpnb+6Tw/gaPiJGOD4HcE40Eh3+o4SJrtnS
56j7LjpkJjDVtXmfVlmq3kbYtpde7pkntDNCiysyZ9foaZQsqJNzUa2d8ckbO3HbZvrPOIM/uSWv
IprwikIZz6whgY1AQViPnwVTs778owWaQv4sm5RLPSb3sNfcWUlLGLg/YLEZ0EmXjzvkERxaPOXS
uFz5A/D/lFSrDbFi2O0/NkqutsWDfxwg98gUTe3dB1JK1mb7Wx4eztEBWkVzn3vwBPq/y5WA/5If
sueoque8E42cfNLGpV4bzEcsgxgIbyWQHt1EinQ45jbKyfx+UhmziS+jRcF4DJlDGQExeeo9CKdg
7mOQq6MocbEzG8s46V3grCaTcaK63XHC9BffqAsUY5grpSRJUKTSC7Pz84s7Ww1qrgO0q7o9Aq58
tl08/HiJ85mrr217GxBBH9Jp+Hzsyxf0HcwG5Gn92j55g5qhdZdhEvFTrtu6MHL13RjpxRTGwD5H
4Q+0t0+kroJNg/om6Spw63ohhU2OpF41psxFFigx4gFVAgzrJbmbktRkHEaJK8ZU2YSYxOGbMSDV
Epw+oRfiFjhd/GkgUh0Vfe1FJJ34RacW3UlkvFufXtTPQZdkS0hPVwNR/SrxOjtKsJ93o2oB3XGT
v/scEj40p4fJUZAX8FfmmNgvAbf3xD+xPgAIe3D4k/4kmNhJwP/061EfOdbt8+r6Q6M7u3pzvXca
XVKdiMsp4QRQFI/rfAgGZxO//OGnmDK+z+pLpYfoPj42FqfNzxWn4Mum5IDGtH4cqxzUBNe+sd4j
w/j80UpRPCVab8xVOTdSyWBaoGW/KtQsnsROYYb+cutW/WoYwM16+t6dDW6clQuWnL5lYRtHh6Xl
pK8++v2cFzrGJWdjOD94O8vpgJIhLHzYnLnt7UNzlIRNnNWD1jnTJ3zIQHp65l4EQj2RLf42ihpT
cn7Qs4lfM+vPSZWHekvaAz9lW7FErtPlyqYmtqfhxFJmA9juh3Ylyf4xNVdDRzQg4QKW3fbJCKJd
WAW4uehBMQr76eO8vAGybcKko8782ZRoyjfIQ1zjBK4POor27pnWV/d0/ZUqiFI/SXpJQAJmihHZ
mE8rUFOoNi0bNJAyYDbGn8movKVLXCK4T+iUcGXMWYuxB5YOcSctTmtReUeE1sKL1a9iiSQjujB8
J+zC6GV50+mAM5mk9Vy/rhcOMyRkXvlqmfH1E+0/7VUh6o3eYqaa6W8vewCvraplxnHl6MIgHDt4
5rd3RhawbQ2EdNSvDz0gtVhNWTDCDkM3RG6PLHs4rNO/V7PD5DtRYiywp4JZC4WiGW/6eVpIHQnh
ZjbUGXYCXJCQ0gWmYHQdIHzZQktRaA/tHuwUV4FdUQpiFqlOJcq3zNePBlFixEfj1csdJk/mjlTE
6sG89oYltS9L3nJ/Q+gPzGgr7QRMfqUGQEcV/yqMOoP2yHg8El3gp+miJl6iL+blkpvMDrgNQFyj
Uav9UfsFtvMNJ1qCTi7gKw7x1sHb1flkc7uNTYgwEr0C39gCUaCc0p8nyjHTBWe3MxypSO168GHg
ofbF+NKO+XEh/Rql4kN/jhKrkfAFxkUr4LvKKXwNzdufNCg5n+tcoRsPWhgMUnW2k7eKSv2XRPD5
qLKcJmthdfnLLbhg537YRXFKx77BLH7FeddB59XDRHvNVD+sMfjPU7GpSDaUch0mDgebDtfkMNpA
wMaTXVgA/2lBL648I2dG5vAFrZJ1M3OvUK0vdljCWikdmwdsRcYU6HcnldO5Pu9fjb5fgQyJPaJV
TFTqLFvX6NwR6ulMZEyXiZgw+UbA+0a+6CViSwOkQIcHidqR6td6oIew7AOvnLR3RzxEQ3UFWv5M
cXU8uwboa7eU7N8r0soIcluc7xk4R2lnBi2xLg5ytSBwnBXIsS161+uut0V67fhbYVj1+prajtpo
OJYspUz0p0qw49HC5xa7AR62R6uReFYlK+aFIiWoBbaV7rQsQvUYuq8dPMdIURGDw/GRM433H6fH
kp69wJp19j4+cdgJVnYuLx1o4MS0QmT+NWBmoTvat8215TdK/p7U9xVacZ+X3cmsXaAr1SvVORHQ
rkTnA8v+lGiRsSJ6jpJPoJFduZmoaAPzHGR2l5lfj+r8Yjnf17oaAJ2cqYFkNUtl2hfa1WGj2oe8
hRVUTfUhBn8w20E1ol4CzNALlPD1NYU+zJMT+A5fXluLKGJgTZmBPZ9J1P5EBPq9PFnY6qHtEkmD
kdp1qq3HrLqaSzwnORYrFhNXQpvgZ3uEf+PF8idW6IIQrmt/U5FWVZTEy9+V0MGcGcegHa5QKf5v
Ci76JHGfbxyx3xMHLeAC0ui/NdDvSJpYsYEKBWkTnkntyla0m2opszV2FM606eiUEYaEiak7o279
/uNASj7uE3XdvYWl3DqPT7Zk0eqomVpKB5E9iuHG7pbpZdEIEoiXVfZD0QRjXR9QASmJxfSzGInw
Qhbk5a7WZw/KS+irG0h4RJx+v5bcArtDCMpCEU12hVqsJS3NBFYCq6wu3QAZ8vrcYHVEHEAzeyMJ
cHDZThH43nxknf6TqOOUV+l03Q+I1Zk+seWmMJWFsLNjKAwRkyr1JgC00Wjw/m/ufo8iGx2hnY+t
/uylqQDJf4qNw2bPoSD72/bLVZV8e+a5D1NWAxGfqhAHnifsEoSsTjF05i7Ez7VGVxdX51P/OG1Q
nzbtU7WUczWqb6HBZYi9ShBNQ53orp7P7aX7q0XX0mjB9UIbpkeA4i8Tr++BMIPg6yioYPeUcotI
TXYTXbS8N0F4pKubNOQuLBMqxObtL5hvD58NgAFdieJkMPEk+eVZj51OXwfF1zs7mU0cgONe5y4Z
2vvFRY7kWyYSC15F5KDzbI7522eTQLWErIHnVS5iS5RNW9N7sub9MR4w2Panlg2wDhxdYKGcsa6P
PwWJy3dqZUx1LHoiP3Ye5Pyn6RRWibsWWZX4ieJDBQSIh0o7rqUDtdhTmAg8OeOWl7wSU/d3wmaX
2oJqMuwormvhfVny87Y16Gg7cAUFYT+SUTIJf3zdXgcuds82kwghHn7gdiyNhkvwfKNznOQD9YEh
A7NBgdTq7tGmKh4gQtyOUzXj2WPWpOSWB7LF1RaLBkR0BvwoIq31QzTlyP0ETfCdTfUwQcHurftV
1kPGdJHvt2R2fwaABIZus+4JfwDMPggk1stk6gn/Ndbhpl01erpbUgMny4MxZHxHKoiIa0Jnt7t2
zBU5kCcUtpixJ8rFhu/HpY5oIDR96nprRMtdK6UZ/pfyGDB7UNABKf4r0KH0qpXcoYGATintd3Uf
AYtiK854LcMfT/RLlC/bSVFcNWiuSAn0vV8ZgtE223Kbq5nSF3rMxPJ7/YpKruRUEtwy5TkmoFsX
pVIhiQatX6rajLoqbRXBxLYlu4nRe3mT5QQf4MHiddeBqPs9CMJztK+bvLT4sHhN0gYJn8tdQzmD
7rC4ZYeviUzFj+C1wIUQmvgBsDKlhmxw9geifQeUEoUNcE1UkRauwRX78QAVxHJM11Aqn2Tq4h4b
6iK0/Ub0uTKTrBlXazPD67hk9fpA0Lw3OnXldq1AsGaMC0wNdpXM47JelEgLrFiUkmcdEMh1yw+K
oJRSxDp1nCh+l0N6khX4v4oQWFuRHdpgSQGn6bg867DmYig/K6ES9QUsqhxF9x5Lor7aFl7l78EZ
LrVhjUO7WcBS6u6K7MXAGP+mzFPTMnR5LvXgPx8yLJwlCfcoKaDZVayPKEMY9klwC+uex0rQZmGL
tTrD1k0AcakcCxsJe7PWkcE+1xIKNxC7K/lStK4SP/00lWlKalE6l4W4DbOpLx/d8mz8XSxTAgRz
Wa6VqADj+8aFZKnlmYGPhOhCCFsPOJPl8IuBhUen7wXW5WoE+kKk4AvQkjuLkMnLGDlViEMINuBC
KlxqsMv7VWToat1/vgx0/DuXH/1Czk5PkkU5hnwMZdq6FY1EXjcHqMff+aO8p36UZHptdNrzwvH/
dPo/LMt/q5S07BKZBb8iMypztGCcbtehha0f/2Yfdg4WfVkKP5RKV2lIWB9586ciduoVdfaScgJ9
SR7MyI+wrShJ1+yLeqJh+7FK/emHJ46DeabhCEc5xNMCDJ8D3GHQ7UIm/RzOG9gjuE08lK+PbKSb
Yd28ALAIuN9q38+G8UWdSh+tiIp215zA1nlhLcBkDRz9BZ4pL4OQBIYPTI6riW8yP8wDluwQVlLB
JryX4Mz0upplJYyU+/8KjNhaLrpvzjOL2DTxiqVlMOMpML4akNgLvONr2uOJL3cfN5vusp+0TtwE
rLBe/Rx+00mOAi2FaNdZCP6xBPzbCY1TCsCl0jYcbJatQpeN40KI7iTsQKErG9M0auQ6tbsTUIbK
7KCjCkZKBgAnyKcfriP9aPVxdqySRx4K0E0HhiS/BUN5wEZAEymgZWYwvn2PA31ZFh3q/AUZhH2p
zC1mrvM715GJnZtaYHY8bn8M+OZgdS2R7kHyYbInRdVN8VyKu8nCdhaLBiVtZrQ+cBdrJOQdsfxD
8Feke+w7QvQVDrM3Jy/KOYwCBs26/jbZ5rPo52rOc1TWgWR7UzrShGlWc57VQJ00+dFNm64gwKCt
kUOCmAC8VcqWxU9Mw1a9BXYfKytGqqVJp6iWokqa4mRd//46MR7lzcurkoQzd1Iadm5J21MIrvAX
+XEsGP8qLuhIHqpzwvRaPoSENRXB8kHpWvEXh4pZQPuoYd9sPQTaTrcSLUQjKXzRm7RGaXRlLeLr
X9C2y6Bub9HFLDkbtPieouH5JJqA4DKmMRkyAYEXmjMfs1QASuhDwF5gwdE6LZz70FbFe2HIv+Vq
LmUzehlnVLrka+sIUsc3YMzLx9fJucUp1FNtARFODTjKyURTmqE5iPB/cfUX28cccvrjxOZenGFM
/1UGl1H1JSrK9VE9heFa17Z1Pndhy4A397IhDb23TVh9d/xtoezwKWjJ87Lb0XIHzxo5atCnz2AV
xfCIQE2TGq0ocKQ21kCBOqMU5nTu0gv+KuaYEuLv4SdiQBQDGnUfXAdppaUKwxy8kmfJvQrYTR8c
buVZdvPzS9PkIza0oOySHCOBZUb3OVkllLy/naSaZ9leXgdbIzfBuvwXTMHmoWiYgy4PR1xYqyrS
Z+mUpuTkr90f+60/53r/Q9G5dTfWCai7oKxFYULwZn3005Z0PNIoURImzf77vq0hkFENtMZ7EZSR
HqWpIVcoGuLkOtpDncBNzTagGIEze1QXE1bfWgBtGcVa1t778A/xIu+w6VkcjpDsciQ9yhnlfT6X
6pT5iTFjMPqpTRh3zQLTwh7IRvgh236FMPUJTRKxlwor1EXlgMf0IgKfh559hw+/SsAh3H+pl2id
gsEV6LfZjW5meB51Ou6sBFldE01rhwBhE/KsAyxBUGzdrKZbnEM3eVuXseVOybNz7ywiDCmFZTeF
ITO0tGTI3MWmB4yeG7FIjstZh21CqR3icHXcV1bgyRPX16duyt7hOG1SeWxgIcknDHXyL+DN383B
U3mdVf4dr703HuC2ggKIlZOVM5hceBbqZRC6J5j0Fba6Bc6NBXY5LLLHU4vI542MLa/VFQo2zPCe
qVsm3DxdZ5vbxdivFhu02crWkUq1MR5Gh4+dGl3SS7ncbI8IuqKxfMfcAeUXydZn2E9VsplmGyyK
ebHVw0yvnTYktq7prnB/bzpEI3cQISN4XC29b309voApFW/GNdwKkSUGAmegX72j+HMj/yWgTMxO
kgcp0MCz3eePosyfi0L7BZkXAlBRV6S42xK/AV8Ti35Pkn1vmGXYvmK9fm/S4mMvQjDHEEOWwqHi
hCnFyhKawbQqStesrbscPuuphhGRIFgzlT/SagRWl4V8Xo6qqjKaTz2tx67JQ5pC92EFmstzkZYP
20vn2813AHVws41BMwhNnL9I2MHLJ1ejsbjqsxm0m46rQ9tABdZiOPyOIf5VJ81KCOfhDRbJa9f8
i4/BpjYS1LsnTsyWe1LeXLWreSS/l2tgp3q1CwRdyeLrZyU9l2bM75ke3vcK4OOSrGVAjEJZq/Fy
sovSX/Fy0qgmk1e333Z+kPL9+M1ytN1buFXtuBPRSVgagbdseKXdgvEdpf3fkmnphktxZY1jVcFB
g2xJu/guJaeUSN6cg/6lWDDTNPzMZeOMN4W+Kiv4+ic3p1B494rhXITaFIvZoeZOhb8tvecmXGID
CB/tajzFA7S5Q/htacPysBjMfzSFTiisMtKZkx0o2jvoy67GXnysTMfHU+m/F0Eec+h+5dFxPmvP
in8E5H4UyjTUx3TRtaWif6MpPUGSo/r5r4tuK84Y5Jwq/g2UdPMDepZnB+U2ZCdfxMqGY+iP8omD
pSD9Ce2lt6AjZpAxgnPPd4Zc4AT1iNuUSb3xmcL3H1dvzMUBQ2gNrqAcMFTni1VnMYu4Mz463k+k
GH+e85XO8/4J2N1iLf/w7w7FP0eduaEF1gYWrgAG0EaSPNabiDUz8qBjc6USlvX2E+o8IcItGM9k
aLCakZxpk749gc24khe8W4BUwBE0VcocvlI95y8ezmz0bB1Y2vgP5KMAU/Wc7j0vcIibpRaRGE09
FeVC3XIeCI6U/e7h6j7FpxMACWsRr26rp0V0hmAVVWLyDmarv9knVMxfdRJgb3aHZpF/H6WSntZa
5sNb987mqtdXItnaBRXo2TmTq0NYnHJYEaJhzeiE0JDsbSWBX/vWBP+cdeW8b/S0gHr69mfImHeX
2htkFHR9/QYbDd7KQaRAv46bPs/Fs01IhupUJpSZsTu7vvTZQoMDONl9YgUYfKvOgUox86IiSAmM
bCtXu0czQW1aNcaz/Z8F4GT3lztOWhzfnstae/pWqzlkUsNrEhYP8fcnI4L79oPLtywtsWjvEpNE
ndZtvvzdYZNbtivrSzelqy8Ma7JxdHXp2o36pK974+c0bLpTX08Gtsml7TnUUqs1y7vZ25tVTqnw
i1JSEcB3YaiD6rFyLlH3UJmzBrS4rTpf2u3YthCK6IKaKmrxuT0ER7LEpXE1vRHSncC5HzPWCTYh
mhHzm5MLnUvPEQywjkO0cCJVwFUCxBt7pq1NRYKKiFxwYpgAtF+zd/Z9mUn4hayJp4mkmXwnXai0
bPjT5zeifBtHSHIIMr+Wa+oZfXtwFV5w+91jK87AuJPOndT6XxZQzqpL+AZ0x4iYF53pWyu/O3F7
Pd/Cvh4G3cuIn8ijEf5jVjSFaQDJwimgiXAFzZE7NgT95Aks41lnSnM7feuN4R/9duYevZTo+PF8
kXJ41/7jprkzHRi37y0XwdNlSbDPvajF8yFI8d07wiJnFn/pHrObueRGFqgfn8lZvLH0HwbKY0CW
jL/j/8dStRnAnivA3SWRkCvXomwhQW6TqQU1QpF05LFPruynHRImJN5C3RjAV6wAUdt6gpfKM0pO
0MQIvRY9wLrq4TaXBr6w0FCSQoyCCGLVrn1BAwvZMZO2pOod4CGhwBtdtQAYsWyXFUumywZp2XRn
ggXOjZVuBqz36rqDnUPhhgvU1JgCmGXtuTDwgKcqwbkk20FlQGpc0RggOudOrEGjh1W5iXDulAtz
veyww9d+heQsL66hTBd0FOyETwyj48v28wI01e+djusX6cNwMItm0kKtLzBhoSxkELdRD48i1AJr
/jRJ0L3NU6gbw20KgZzJCinEAINQLmM7aSL+a16BlZuS+Ymg8gSB9qpwZ/ZzU9HBF+KyEoStgVVV
flmkeQ+cgt765s1wqI42BT/2yTiXB0fnUhtgJdiQE83GZQNKS9wXopsn6ccHp+b556oS5Q5JFvTA
zqWmuhEo4VDQE2B7mum6YSsctaiKXC5kLguYhN0CKPQlGYUStbndYt4yBHMwcsFMXdrM7YRMTq9k
XpMp5RXRfOdO4I+g7otGSuS/xGmHnE/ux73h5U+sQyAZPVjNhMVVFEbQAS5B3Kn36tsQu46dKF2V
Ziv4ISnD4sokiE88C+qjjjApqEfQX7ITx5s5eRdRvjfqD7D6P40IiJoi+U23pyVbj+ACDYUoS4rh
/ANcOyur1wG5KuFhfttuz6In94NxRC8pGRtZrCKlAjVxi8C0sUNO3XmUxXUfVnAQfIjMMiMX5G1W
EVCtLXhd+w6wlROsU4SGwvJL3Yp/OIAByx0qvF4Xve8sW4wd/pxUaOoCsH8T0Yvx1bnfZ3QjJTY6
DKJ3kSphXHc0JLrOE7Xw+SLH0xNI78YQVcEXfh34gN/YZXzzMC+vfKpZvTzMe4cvDeMHNh3Kh2VN
EtNynu1fXNgn7JEpL2CMV425aHGrHtjGMyJ/PZ0roOEp6fyoB+SwekqLRjWImacUFCRVt7NmZm0a
85cTE7dbG03uUvAtHZVYa5S65d0Mcx+Ob1BxiG+4GhAy+coE8VJRx+ZzY/zTpHOuIXWSWhlDxGiq
BmvFQd284CveXkqbAZLFwQqCwolM4qzgza2TpLG6koTBxLJhG+S5F818+bmQYhS/z9uCJajNiTQE
eRXD064p0or9QXKY5/IhWwxxg5N89gCn7lhn5cACWbRvOFsxRGJfn+9o8vH04SYQcNlX/LRPIthS
WcQOCbeNrZb10Zq+b6bTUhcwsMzwpGCK4E90GfcwMCUEXCIk1B5TP/rmWQbUK2VkeMDSRFq0RM9K
yZHOkhjl/c7+Oa7agNwsqOmqM7506whVWTzptvWYNTUPCKHVD5L42RWfdAzB6XhRybH4AfQ1TLY3
hgl2JyQ1UZGcRaJ4rQGG7FtMZtOMswOM0TJKHhefLixgAdObOsqSBdjMrkQBCgdh640DKkvH8/PQ
Aw7vZPZiPx70uRxxEkN47cc5xyaf+Wx7hVlE46gahHwkU1N/yvDQkDPI3RiOPgBM9GOpLROtXnYG
kCV2Zkn+k74Rms2By8qbvjP6WCSP9+Y33dt7DRkvEga5Y21UiIpxd127AP8KLNetBPdn3EMvPiuS
pKXs1wqLE+UQ0U3NTmr63fGfnC6GV+vEbjK2zUI/bC0XXAQxVxfxD3h1euCpMIVP7F1jfmDgdkpR
0anWO3SfGrOQnzHJ2+cOrKcAXfPo/EQ2CSlSI+OYtDmEz/j+o5rvLiOESAUfw0Cw/kR+nOiPAecT
CarT7rul/9FehEGq5Epl7JvGaelvT5V8Fnl7WZcQcYdWGa0lWLac3Lp+i0E7YGXzsb6MT2y0PwuK
aJXdkW74pEBiS0I5aZ+h3zw+4UanbxVmfaz6o8NRsw/ZTdQTPdQKpW9RyiT3VDg7c40vwByEj3Zr
ANPRq6aM6G+pigiXyGhjVJWu3uTd7KRKD8GcF95SJepMPM2YSaNkL++4eaV96/CDQR/HJZE4+BJu
9xTVGvQjc42799MQk6rExz6uJdXma8+2gqSWo5EB9QrFQH3hrDHLVo7DF9C3Q8zMsmhRcwzJgkEF
ewVs7TzkFYGyBAQ4op608ozj7jQ3HodI8WzljIegMm8g1OvFoWP8GcT5Q+0kaw+BjcTB3fwaMRwO
nAaUmnUDAeA7D0CsR/GNlKfbapViGeueMdNyLbvzbNluvytw5jYYJIS2Uhn7fNO/PzseAzmZc8LY
0PxS1U/Cz2XyhhhZpFPF5wu+i64QC2e/WQ7BfuhTVWyNhzNXl1RC0CCDrGAgJ8p+snSi3KVBpZuI
4u0ZyVqSO/Tlk29Vczqz37IQ6BFsv9MFRZnpYb3yTSvYAIDkQjqqJ0dqI1g8T6gsCgpV8xcvRxt3
FT72REG9rJoZ0GSoYs2y5XgY22WzObHQ3CwXWTg5Q/jMVB7/8xXvVLRPjy/rMwE+qSheXjmwl+7G
IrJJ6Eac6jg2bNklQ9WS96iHMIWq45stwQFN5YCbllnSDJ64LAwhEtwqOjJMMB7mSXTKo7GwHgVz
d7mPBB2tTKdFKihi6aCFwiNivBp3M4gwOsWqE80QPrEs094JPjIg4KI1Ql1Yr/EL4fSQ9wRe07VR
ICMpxYzgilvO4fLokQqq6n2hFvWHI0evL2v1i/+nKFgWVu/9eqyOB/x58snm2aXTHK+yKviH03V3
MvZKCUn5+keDRdM+EaNLZwITUni2HOwoFTWycTkYtF6kOeYDsydW9yxPdLyf2gVMcGxlUHLX3wZv
q6RXMeEid2/OBJLx5fFwqk9uHEQI7ChvEUZwypHzCpHG6bj8vBpwiH8UPcZ4fPMjg1M9epAsxe0D
we+VFUudo0EG3DBYj7MBxcDWpAshqK/+ZO18En2Vd9Eb5gdnbNepUAvaei4TOhZkOV6j4z7+jeCo
fzuyWuP2r/iAyaJn9j2HmXKj/dBAqwpuFf3d3W8OnVR1OhinobqM83AOvXiNlEaCl7iHXkt2djLi
I6/19hm2rCyX8YjXBkFCc7Z4mixNuJumhEVgb2NpSoTPLvkDQapLKkdx0dvdxtJc6p5y9iqv1417
vWjwPR1YtRPZTsukW0RHtTulO+x6aYVOzar0vw9FTJ8YheIcPotH2YQXPzJtRgzowJAZPt5UaIgQ
MHM+Xt0uXfWYqHXQZs0LE05JkEIvR6xzIU3DPaHaxfelNvJJ0d71ZcLwNO21vQ8GHZ8CPdNQ+/Y4
T+Ly3P51UODSMh/LXQZfHEVKAxuzVucP7P2yVLp3kEqHunlyzHP7j7r9DPdX8CEo++jb4cC+/VbZ
3S9vProXBMoqUV6+4jHN9jP3Xh2Wr5vjKloI/qjSSBHIN8olL/YsfQa8U+YcEnixg+7OguAPQVMe
XR+qqVFS6AFBvJV847KuuWumMuxLechfKl1jVUM43uIHlVZcOzrqruE4yFniTw0ldksIUKXGeR3I
cHc30w4MYbn4J7gSfubTlNFVUcOJjkLuewOyKHp8iybeVpMF7RZ4I9udHW6UneLKpD+AM7eVl5rI
Nsdu6zbpghbLNoxwbbT7vqQyXQBzpbslYHQlEk4Nnq+51DerUqd920tglRnK60Ww2idSsUFveZAu
88hZRAzM6z+/r5IVvzCSZ/nXq0DELOXAvBJC1OJYesc5uGbahmviqfo+9j0yJX/oHTPP89lt6KFj
gIOUlSICpdbQa8PyzMd96IE37ej6aBNxWaN2d9vsYKcLXfv6rJ9M1XEKm0spWxKGTLZBuEMEHTde
dHIdWzxDTqhG0vksCYTx92REWQ+7loadO07SET5E0RRa4agnGEGOXB1aFi/c2FlRgjIbKNedkPiV
QNzoVcohFXodv6q/C2TO+m0TTCdQKym98JwzgGykt3iyNkZI83iQtY9+PJ3IbL8aLvhiDuoLdKZ4
UF9EOZMS3x37je6VcQgsc4y9vAMZvuU/EWw369HTnOdoo1i4EBrHMUo2L0AlGIdL9DzsfMobQPBc
zGHUL4I3xgXJNREXWm+zfTSi25piZZu6OsqwVfHVSqVLFtQ16FgzS5qowoy0P+YXanX0Q8b7wKSW
EP1k3DrNsnRTq1DxHnLIBa7bg+BY16Kkkl5R+nEMjq0pUDv0oF3BLtetKZ3YYVxAVAthkn+Z7lm0
NnDf9iV14Axj/I+/3eQaEGtNr6POvcJBwrK0dLEayJuR/+KmvBdHZjqlTsY375vvW4LSZaaa3Skt
+IUsjrHkHZF1bHuMhYjr4LRdSY8j/ecY7M+wS08IA+YuJ9bI8ukSpvyBZl9605z4nuazob6iZJso
Ee8MyLKsS9QoqiVAdUQAo2DLbHMcqKKLpU4Ik9QLhTnBwaa28mAAUSccuD0idJOMJHZ1BtyBnvlf
cROTtH2V1NhdVTjZ62kd182iASO3UIzkeucEgVz/o8MLFiiA3u4l3uFohNZ6PKBs0s0EfTokVcBg
hNueF/+qtLei+bKuNMzdLkj6MyjQ8rSs0/WqIEv//0E04q+oMeC2932feHch9cwslyPNE6TkqvJp
ld14d+Y26FuiTXQtDhbpuJTuvKj21RpiU31g82BavQ2AITue39e03Zn3KV2wnOglRZ3uWc8nPWdR
NTaO1tW8bDTj/bik1t/Gq10zMmMtY5PDz64i7jVmMmC41a+YMJXxlQ5Ti6nQft9b/ueqKzNDwL3y
Jv0eCbC3PpY2lesvZrKc5DHb6wiSwNZ92caO1uUrqwM8kGFHH2ppu3MQ4eWjL6ubXwQDp0ZYaVjb
+lJyFCeW9DS/vL1gLRHc9ib76PZUTuRT9zL4Yp84kREaDr7zHMJ67/2agvW76JDsoetn68OnRK89
KN6OIuxDWfTMMKdPUP/dIQR1dT02/VYm31+vV1HyPtEjn2pYub6TFYMgtyu9iScI7ho+wo4QxUc6
oLxhgZX+vVRPGDXR3Ennw7e8eCBGH8vsUtP1h5KLwO4tiQblZXKVRQP9LaCFo7NUcxDiW8X6K5ms
1MCICLuZoXsiNh5LWvkKaWu98i9xcPf6ie7+wf5y76U+boCzk0pDt0PqPdOeTn2b6RYeXgOfbtnv
EEu5kfulz5oftwgokhOkc/d5X+7CrYnnrHQTEaWnGr1D7qUqy3M8aLggqu4d/onzbJto2LjMIQrX
15EhonC/Icah16aAmlpY9qn6kMcBrDAz5gDzqbSkbBKGfaAI+Hi1yVLxbCBvWOeKkMTE7mvj9hDk
qIx0UzBK1sknMKBIxC1V+KmhIQjC/BqVbf20ThxWm6+m3e8IoF7D7G2Kewk0Uf+On4jtClHIVudM
Do33dWpnOE4Tgd+mUI43oo5zA7A21HqIHfkK0N6Rsv7UbAeEncv/+3PfRoCOb/IwcD34XL2s8nrU
Zj4qBnXWhLHGZgoBV7oRJGF4A0eKgUR8haiyqf/t+0obMarlYsnB8wIy0pFgYAgWi4LYvpdi0L5F
NLMi1fBrxgZrjkYqna/DcsFySv4qSeWdoGQ1U2RpKJdzTQO42J5wOzBj2Qv4tmnFPJ0oJF2mP9gL
xuKrjgF3WID5Gqw/+6/QHZG/K5NsQCJ5EV7WVETwKsOUYasAwU+hIG6zOtHDYUxLtUGAvAUo9/G6
zeEen+ILLI3BxJOpYuB48Z1WYJOEmIe125nmBYRGyD2fXMLr8RRAxlHjytYDmCxXqXcL2niNAfQe
wNah3n6KApWscCgsc0LQnDXX5jBxy4gbuIauLCriNhf7rM5vX1I/R5zLiK+C47+o4hx4AYWbFIp0
akn3100v2JVz5y4FgWp82PYoLGnCi4VZUc+2OcTrjb9CvM7t6OOlRD62azoBsiuFsddHrwAgn0Yk
okk81zGsfIJtp2WaQ/+n7+bTfXtsXvbW4+qn81txJ13TLqR24i4b1kMwBtUaMeuqrFbwXFmUktJZ
dmbPeM9rwvpG0tblqa28bCsRTINVRY990eMbdCtY/xEyxmO1aqN8GvAm2Tjx8fHSf+fbTCLyIJ4l
TQVozY6JlRanAiQJQZgkcvDqMwiX55yCHcltgCmM0vZuMlrq4gLHWN/hDd0g0OzF4RR1usGX2niJ
oxWmcUPkve9ZwFAvXKpAQOGZHIf1wGAdwxbrKMR/T/grj9Anbn+wJfNthRJbcidhWUcLBMuwGF7W
ClEDfz8isRwJReeNUwS1nwyMF4eFlNf1+XprCa80HRjZMqE34Bn86BgPFV4rChi3/3uOUCXFkLAl
sca9TVNdqbheF287laKVuTMyO8YtS9RT1mx/UmX46WbkdUX8kRYqLeJ5UlE7YvNUp9RpOCu+hwUa
Mai8h4t1fg3S+l5H0TQ7s4XaUdnzvqAUwCAV36VE56098F3VpQHgLhfUnyVXFvsxqU4yiyrizu08
7OFI9EjhBK84Ldoo52XjeHcEyrXmTne9zMXNaJ+MZuLolD7bQROby6F97mi8Ztg7yjP1630Ua9nX
kNHDUVgp/Y+KOlIX+b4fHNGdFmH2d0wEYDD2iumlaNdEVEQKc2m5dm+nQkK1cZX1FqVmkx7N2zZV
8Dj2edUZ8mXGRyhNY9Bx/cmtKEBiCmS+FH5q0S8v3r/4bd3RutggzJyDYki22NdE6X9kKcdnWgy5
nG78nWRYiX4PbSZu7/FrJTnUNsFOcxHiMkYz0Hjrpj8acps9UubSShM+2ScysHsPWt6c2J25dIYm
Q1wEQQbOk2CacdXcf+zwyVyf+mUQ4nZ3P6X9Cep5QwZXVmue9UQHvE7J4ZiTyLpKBYYhlo2Amlor
+eAmGxf5PaptXq6NTBMSk0yLsVO0WOyMrBIOR5Vo0ufTRNBZzIg7k702Lp0AcO/Rpuh1UFlWkyWi
Q5dTwvcSE7Zorwo+zWYZb6VB4xvJE+4oBDQTYsDImEwNdz9yM0LNXxa0NMJopG4K2Pi/eIizZAVW
FBPBmdh2eTQ36LtPxi0T82XzxaALiAKxF9spY2Vvdi5iiRGbH/PrneFPwm7eF0gGiE24cpDMbjf9
KrPoKC+by4vA/idqI+ZmqqTdRMVs7HiaAUxDcpQezEAEigqI5oV4d8IMekiUSMc+f81oj6Gg/5Uv
TTF4eg19EnYqsRH/Zfmz/2mQIe1lpBUuUMfp10kwXetZfbA9KBIstdqt9aTSdhY798W4p6U7vQY8
XTppOo/aMJTihrJjQP/KI1TA6y3SKGJmU1R2OwdnklFoXaWW48IeClFIZDGAgl77ejzUH3cmEu7I
QaLtHJiZLFcLxcKZ/YxOOAN17HIMeDid6nDMSjvhmxG+bZzEdqdcU+ceY/Z8A1WrTKZwf3VecHw5
rbjBP4wqnZpe7swCyqqjbPdZchgkHmWODXBkKN8Pj0PU56OVOXC/suWrfq+7CS4Udkifspgypzya
kyqdc7DDMv7Xxr0IUwpyo/vW1J1wVQoJ9C05cDuadF3zhL4f3343MKiDiQSqOuIEGPjQu+J39izY
gHPTegUCGc1uUHdoFA4uKwUNNmbn6FOWINYvqcdU618/bAAZ/oC554HX21UJltXRr7GQumjOdt6o
mRMjI5O6eBzw2JygwaMAG8LuWUnFTlQC4IUy7Ycy2a+tnoEAuk5SnVzeuM2SnC9JkRvijC7Wsu1j
jDoUhGp8fYjL41rQNPfRBJbYCKLkfiMstNDTxcc5QhgNrznRKrjXhbBY4xWjih9JNYEIF/FJAYjC
PDSM/3AdJ+nTdI3syzKgWmiuteFsBZKC34QTo6hxe4qo61mVoGsdySzvFfM2TLrUacIWrf5jdu+x
IWdgJdjKO1ZEuZaBq/3DIYpEq9qqMzh1n24sw/wBE2OoR6wM7PTm19Uxq77eTqZEKWAFcMcjeQ4f
jHa++EbI2wmLHaZtMpuMhrxsmj53GF9qToifdyNwXNXmaE50a46tncDFrcQ5uJSm/uxk4jn8RG+/
ZaEYemfXd48+sfE4iEz3VHWzuQ91CIoL26Ay3bWZ9MYca0PVjP2izG6tDATlJhr3MfPoCi+AGTru
6Idy8vg9nVo6rKDqzZ2HxaBsGp7EWohrZsx8z2uctGCJZR4qUJlsORtLx6NejI/HDhOrCJ6IJIxq
GUgpbjVvUxz+nUUmf+dwwFpM3ChtEHAt4p/jZUmmJ2rjBsGye6SI7Ngym4P8SLnwaD/udT4Oj8sU
WDOqoARPTBYebU6Bs2PLuWTnWQwY+tyScWhcUnXpU7tKjoejX7xTWcWvrq3HeWLBUA1syciMEnoz
vGq7NTVNoh/8ZVyI0+De4XUGUHlupFPmmbkaEVK5UMlLqvD3VZKD+tYNNH0pJr9llytgPSb1/ICy
5APM6jZgg2+5OgO+m9BcC5rOndTvmq6XFXXYcFlcr0gzELOHJmioUlro2F1gwbTW6xFGyAObLlWy
AVRiO9BYzQycMSGcd9Dk15gRAuBw+gVHJoHKhYcptMo/tVEctmWeiHTJly5AxxkLAaGGaNt1lJRX
IvcnHOhpg0lUYx2jBElBj/J6c4X6wTGp65ng4LBGiraJ3HKhfIMguB4P5jUqnyTloYeLMZrevnhi
x/N8eu2JUwUTsEzXareGt2Ak75ZzBcyFaMI5rE4niN4utjwa6r+1igapqlmDDRbH/AQCUmSgTmlj
FHthg8923EujDOmjAzAzZ2pF9K8bwwioKaFqH47QKeEIZwrKW8oVeZDFuDHxmzOE1R+BrHk16wDZ
DkDd5TbkDagmTceqhsXNW/LEXyMhVzZOwDWrHcc7/TTmBBQHHBBEvhgzoVhQ9PPuR2OEzNKNsYKI
eKCo3kkzBpQ4G7n2uKKC1LH0BsZB4XGPf6ht6c/IUiNzZJjlDUXQcfipzA+N4fkxh55aeCgl9W8F
iKalejvT47Zp3odQtnsDdO2DNXyBkNfNAxGpx4x5aiuYuFbCJlBqV+9X8KFGx6cn8uA/RityWp20
tvXt7DKDr3i8tGl8rBdukxbpAtCdp24F9oVucVOLstXEY3qFq01DrKjtBcDDObzPI8QK+o0KXKz6
86oLhN4anTzcqxF1jeWF/vsmQGBRKz+qiWN//WHYza47n8+jAmVIfksu3d11Kn54qNZyRel58r9Q
Yd3PtxdKw5oXj9TVdeg/iHh1IqEhhTGGYintgem2yHV2YbAYznuPr0kG4eDhaWinfCrDJUIbAq1a
/1K7CFmajiTsoJBt7FUIGmC5JrYhDTCCJk70jqSIUiQIS4Tmz3wEKnnu+YAYQ0NOUlt/1ULRbFMs
ZexBHxQmg0YzA8920Zdi6MT15MiHT4Aaj08zyiMbohu9+SS2IL2/1qIJf+ZC931MgEsspQhhUaNn
jqC26Hwvc+I+XH8SwwpwJOAwsUqtuURSvqmGR+U1nhl89qgcOXI5ujL8AKWc17q4UedK67fCtUP8
RCqw+c3Zs6Ol7XJR7lnM4w1hioRFnstrQlzV2RmWN5soaTq/aQdwGvzO8cFZSH6DrF4OpqQq8QC9
43IzoMrZj0uzA6E+DrB5R3cIONNteKkQSXCYnhnVccq2rF7sUGh2JOJ4L1FsnGl696UXOcM3ZEGV
ao26x/jCHzKWt+EN1MfJ5a4mNd9B5tdgXBPdXX92nOnEmyqmAwRlrarMlmqzNtNbixfcsr75GJv8
n+nMx/Jte3HVXsTcd0Qxy9BptD6o7XSO1mbsrR9bcG7DDL51g+kFLG9M0xqVPuB2z+82d5pKtW8G
xsFfeOr0+FC5n3qrVGfvoR85fS47se29eNrFpzURfPuEULnC2WJpqv3NPd4PCPoH5TJ71ILvRB8t
aOpDXws+t5e1XLF1Ctk5UAv+72FUOHcE3bMgOS/Uzv1n/GoRlso4A6/75uTUZ5TCQMJgXUtIOOIs
R79n3bdSq1Gy9kZZqSuWTnzazyXQXK1yTRlwG9ewKKDh6jvRYjzCvuD9FxpAmNU8tyP/p5DH+1YW
ZWBNO176sUjWFqCsr9Iu8sUlUX9LIxfFZMb5r7Yj2rf9mnjFjHoHKnk96MAF1nItD6NxnIIyR3xJ
NWWaaldt2NAPdOVFpJKjDmJdvE+ZbpydpfIHVYLoTNnVXv3AoT6tOLsTYXNB+8kYeoq6aKU8XRLH
eKl/g4xJuJGUBUxkBHBQBaWZJKv+P7lRpoq+WaWXaMoJF9XXLQxLLMHxLahL+Xcl36DNTJBtdrbF
hmpy7CKWW0qoSJbSnwzmtpb+sd2q4mf6FXefIacAiN6iwHRuo4XEXqH0U7DAciIF8q7Xu0UrpUhl
03zDxtsmG0/z5r6E62B7z2Y8ZDamrRZV10NayNoOVlr1TvJ4T3ZlQef1O070QrAheo0lOENWdhh8
+rwvJKuIM3ri6vkgNq4P8APhf4mENePdT6v3QQoMUakIf5Yts6ZTFXZbPMLFUVFFdwlQ1BGP/orb
pUyFGusjk0fH8xF6g8/1UZP49jC1fUKiwdsw43laqq4asPz/CjxOu/SMKkZT6kz3Z4sPu7AxlRO2
xkTltTNOq7iAR9NZ08HZrHTqnu3fm0XfOJxP/jDFBoBZBXmKQOw+rNjEiLWOzrXHGZ1R2tcEcrWA
EMx5YMiVOSLiYWrwlXWakvaIIcDpKn4TaPSKGYheO0G5pvMjMGxv5ia4suUx5POcaz0EA1vCvd8Q
peeictREgrPTTbDAqS5sFNzCTqnJYIOhqjm8ZnKFzXN/RVClqYdJfUtnTjYM2OEiXJjdQ7QtNoej
zliHIT44W2Logy2/SNir/5O8lzgwOVmHo2bUfwagZBEYsun9ZCVh9yUWLXhVQ3i55Jb/Dttn4Oow
RQ/FvjjYRXGp6dIsfszoduoz71OqzPnoc+0Yjs2FUCVad+05TMebFT7RWJs2f/gKu2CfrQWn33ba
E8jLr8F+uH3Ge5d1YfbazcUagMF+H0KosSFd9npirEyF5oHW07gMBZTe37HsPEwp0m8xRKBPXHZz
Jl7WOVB8Y3OrrEsOumG7rJHc3BF1A0rKwyJ/GAh3WtBrPe8VfWpqg1+dawVnR8S8c7at+qc7XyTH
E95BRDC7vteFuLnk4n1fEH2ElKIFVaCledHSqwOPbcxPV29G3n4uMMZgMUzTKDyvxJaL1GkO6YPo
3dcqnVPGO9dblJsDGlYWry43zPNSzhBUi+j+7iv3/6fiTJTGCp3yVX2gaEEKUU24bhUITQvHJcxW
x8uHacNGfaYFIAVLe+jG5tHPXtgd+mMtJTBOLLwPDPrT56u94W2O2RGRFCbOTo4q/1E7GbdrrA1W
N54PqsvQhzCMOPrvFMUSBMfgzYv6a2yG3j/Nj/KVG84WWsjXS+ZiPrPgxkTO/YLM7Ri4JG6xdKYg
qCn1DpHupNznihP8nkJyqz3NpKtxMUpyStiBCKiYMaebHlI9IThYafkUw7H2M+ctJ8wfwZqwq3q+
pPYw5312p6gGsL5WVBOBVRTMFQYm08pIY4qvQw1/6FtgL0l8oyxxj1ilVYvNz8rukjDqgtDGKJK5
8E6MO9Hw8pWnHOY3OUBRmBz4ihZ48CS/sBczD1PTs+rPiLsUgOCq+MyZ9djVd0J8lMDO8DWwZmrM
gy3TkepeqDEb2ogQBZf2nznmOScmoI1kVLdUoRWug717BYdllNLxpR8kQ0ls5Jgq7avTxcDzQ6vR
RN95xBiqPQjiG8AFsIq7ZtwCNkUD4v1qvSBPrAa32uOdSzPsc69OU9cWSYdF+rZHTru/tzLaJgBx
/QeFEZZk9APt3zZWdHJXLQSgO87uDS8mvOaK+l8u21Y4j9kxxTwIiNfzypwE2Jr1MzGWJ2AqJUTc
lFmTBnuIhwllS/Wy1Z3nFhffi/lCMCmwEyLRAKim9aLMhhbLfkPE/gdp2/mMSMOXT0QYtq4PFrd4
tb/PJbxu1EJmLC36VtM7lIBW9KCBif4SSpWqliIyh+9StfNlWKAiPMdYGzKNgcrmfxdyqQILUZW4
gU8zvwtlRvkEjsM5dBqMM+ytxeV7WpVg/SjmZr+4ZTVDTBVjbm2MzZ1ibN8EXQapY9SpusNdp7Za
BjuVfjx4MG2KsQJMbPW2ZjkLt/jgrfr97so85x6XuY14XZ36EcnDBXo8wyiE/MnqPExiQPd2pJ93
Pe5NxL9ny+vbFSYh+2KVaKw49UTU50XV4oQ6drRlJ1bsaobwhbr4FR4ytqsNzbaqYWK2zbZluIMF
jQAqXNXj23xl6mlumrhmDFNSXruppcn5GPE2CfkeGjEEMPfzeoBusLj0VG3Gqiq0zMUu4ZzFi6Ie
0RC121eYuDO58GOGLKBmr5FY3EBcj0HgRCOIElSPXPi0p5HXTDJF8ZYjTbQTPBXGEEp+hlypxcDc
K0ID1MXFDX+2XOL9an6hxbbe8PzCc3ZnQjzbHvfMiY0+icqmz48sE4ewzOUtQ94mYYg5mYsUxaLz
cjSG+rwEHFlUSVMkDH/q+bViMj6T2gE1y4Gxa1TVu72xVkAo9ek6gpSranLsNbqxB9fvDvFt3sms
JrBlGivyp3cHPrv6n1xHU3iuV1NZkMwlwXQ9rJwJaX5ZKxpP4/EARDPf+b7dom9nV+ksyCAGnw+C
VwWZu59LrP/XloUCh/prBLc/Vr0mdyEAFUcMLOGD6L0kuIGqA/T4EePOAvJRiUhp83Av3hBC6J0V
Y4N6yBpc7jr6dbMQjsWtksEnDOeHis/oLOzBea990+SAVWAMawEaqqM2qEdNrP6jeSphXeCJyNrm
h7qzU6/wHiP9y5H8PXSBbm2VLP7pZqZJsFH1vnN2EwSqAMZST8qlEc/3BJu+gaX5YKa4I7NDVwDg
GTox12EErTO6qU7pIDLG4dtANX8+d7Hoq6Rhdp3l+H9X6c2gvCwMUwMwk3wej2GAorQq7iKyO+p1
XFbphRDPkRFVbjkkS2eVKM94yIP2M8PUXY8FR0MTba8veeP37ke2z86EyglmOe2Lmb1BBufP4n40
ckrF3q5SJBfLB0TocpHSIEtqsHnpVePt+rhYgvXaNq9ZhVmDL20vi/ta7CagMdXkpH4qXxp05AVq
CTHmnu59ekb1D/Ha7M+FmE7mOSAtYrlKIb1aRrTgq2/9bT321O/VhoaoJC44R1vDTKSMFmWEHbjD
V1PCdSyBRzVAVWSuh+DYaCsURX+cvS/J0wZAU3rtgNI2kqPpZy2mtlbAPi0wGscvN9pbZDe9wHoX
LSKyjYVgi6Uq3iOFfVZfbqojaUqPl2EBs1TWCZeii0ZYHu8nzPZQWv4NX9WVNSOJP9ME7JRgpg/F
C7KPFCRSAVgaB79Ge/4G+T26o5Ko2cOOlqQa5KlVqxpV9mPwnNAcMEaUh/70J2aT0lWk9ynIMvJG
IbIK2vJ6V1DCmziWi9NNgCHsixvu6ker02nJgS/qiWMgNhnaSDKqrnSXHAuaTVATtYdVy9h006Sr
XI7+tghM6ZDdC2El/5MlZNZQuuN3I1AvnKIBcipNYa8K5chYiccAS+DYfJ7Wc2F+dsYATVVda5xJ
eMsr7mmHX9zBJ11FniDU9q1ID2Kr7YYqtdac8AqTr7AamQab2u7CpuHglV7RB1beiJOUsb1RzO+p
V9efsxDeY8T39IEuttROjMDhfoHqG0vzZ48MsBcGLdgjgz+3HXj7zopjC2Xvjd/5eFd4e4LrRDiE
QX9fkbuy1HoP3qKiXnj9xDo5bs9EGm3dAbPbuB57bmaPRm0wBqzUpg5O5V+CrOyRjtm9b7UxGIcP
HJkntDvZWbSWS5yyZj4Um6WiQOQVlIqAPIKL39wraZkojbHNvWYoiH0N3chds7pvngfsWzIhp0mK
ngrHcpwsWX0zAEMN7dLnw4j+8jNbPsZUnWdrJ/xH3+igcJghUAVVIPsjS52Kil/c/kbPlFXY9bCj
26JFQXaOd5/j2zEV0/hfcvDHH6s1Wrs0+J2DsUt0/fjcSYSWOwpa2ifK2UuFoeEOZtKUoTlVRHa9
JF5vW21/D/8fe4qAZiiTsOvzOHyNHou36EEsJytg4hSUHbDa7Z9ekMExrlZ+v/xky5G+HMJmvrF3
W9ofrJNRJ1XzTXe8vdh0Ji2/bMyuHbaavrTxPWRYm0oJKPzWVUR0GRXRK+S5nGXeaFr3IDkjALN9
WRbnr48hayM1Qd3VN+ZNdfJbxw6z1syK1Ejzueb8DSlP+iHZj8YtSMmhzxJzm2yTFwZ/ocEcip3w
F847H1lKH7egNNsNijrwis7Of3Aqtf5pKADMt5s2qPF6TW1o3pMh8uraN0ivAPs+DqjfFWnPtmFo
G2uDPd8obojRLcTx5TXBxQ74emQ7cTrhxpbRHrXAc2rJQBmuGveJQdCBmpRZ+q5OIEO/bCs3b9O1
ZoBbdWxH/5HtDAWJENWmSM0fDjyBPGFvwIVPD3KfywMjRiMR6419eLWbarr+SWU9Tu6XJ1wK81k4
6/KgBwHdWa+nuCoLMkZKv3AyWrAgm2/8u4InbafZEcE9LDOdYksn5xbMOV7czTkkb7uMvCrV/JMc
9nC4aIJ+g8UGNABSw5uCRM5A4qkKHgxk7zEDMYf89Opv9mDRhEQYx08xpKXq0V7unsuKwdOcVTTH
mMilUmhL6+dc4Ui2XIPav8bTtULnohgjCr4e9Q0ZVi/1P1EUU1TI8PvKCF/J0KbQrNapR59Ve4c2
wAP2/tT1sdLkjQuAAWqNNIW6RXUCpfd3oxfCooGy9E9vPG8bxDDAAfYtLC/R8nRg+5Ym21NyQO4P
yszidrBUfDfDUPUNHpJlWxgnrrrK8/YEVQ/aCSJjPOV2855o6z0AoEMs3XdXnA16rwy3KBvLt6Pv
GOTp2eAhRcxKH9w6HzYjYVM2Xrz6kE1hEXHFUAyvY1hieTq3dMgaFOLhmwoLC6p/k83I04ubJDIF
3YV/4zGRj2NaG/Y6GK1efRnKvjzxI8lbOaOejplT8MxX51gtuBGkqpvYYMr4YeTDoegxH4OLrvKQ
vTVs2KtKQYyjFyhmBfjQE7FQuK15RATa4oM2/z4hIr1bB59IZ0FYIIvebIs3bnneOi689mzB91kX
39YYrJZMKV3uVcgxPVSNI4Z3kc6uLbRBkaTzxJdbvuqNflNo2sqZ26ewgISoAnhLxQXO+gIMmx1R
3yQ0mg4A1rHe9u2FWgANDPGlfAYktFZ0ADEnw8+M9v/jHQB0cYNv9aq4FRrByce+TRqrIh0n84td
BuCO+KYVHYf2EvSJ808gkn9AQ8EkLpd53YZaiWQy/G/0lGlKG17x6fwz6pTueCvDCb3wo6G1lm/z
YshbmFmkvYd6Kd6Ip+fdWujW93XA76K7HbVJAZPbVLJke01E6aptTwPGWbErE2qG7ZyuVLtNjxWy
Xog4VlSH9LcK35A2Jaihyg4WQV+QJeP4RN+jbBSEpytrozgr7QRIPyvUxRHE40q5AAyGf1EAUQkZ
PGvFW4C7cTp19ssfIQHo0vCv4B+QPQMWmwEuP/OPzCRKZa/u720xgkmXxyyOytw9U9ma/uNc1rwq
9xtUp4NU2PkBa1uxhAqwWuAVO2KhCHglUKBhHKnHl+QGveo02ciuEtirJrnjZvCa3C2wumjcHwAq
hu2VcmQqqWFhTSPbmXlmDW5LYFsfg/5y4qpmsUXmFdNx2wIaK3cAQg48KcrAu19rU6VTKPRf3LMQ
XwJdOhQS4pv5ydaWx2Djrizrl3hKzHbhtTHwbmdefYjrY5lGpBGEg5PTJwQsUQ8uWDchBNLOCG7z
wZYxWBVMFMzP4bBFnteYdAash57nJsHt+WLsroE+SdH55dPh8sLCf0FSuWRkGUWLoTuQOi1QAXK1
LJdUUQJmvscK/16YOl4XngTjqtjdHg589ybyMhCGZUekgAUSptNBpuJvV9Zvx6B03iNZ+pPcySdg
pKMlh/ElvartvL97YtAJGI9z6TMWU5ruUlYqUe4ubf9nVGpGSOWYgNdX2+3Zi9EiZB7mB+c4yBk8
QlB2dCeObaNb/ryKGWvJ1cj+9N+BoDUYfQiTQxpi6CN4lel3fbqMUkOBgfEpnR+ueHH7C1HaJ9Oy
cGVjq8qRWxd9A/82/+4WjK92UAWRCm3CzMnhd6+Wny4QExCyzmeNzZ14ffk0nZ+Ejzni6mjaUX7X
LqRnXSKLNHX+wtsnU5wGpMzsCnSTziAgR9vicN98XI4myCHaaxszcpiJ1WSutk5ci79XWKt4IO3r
beXHRQqrXKUERQdEnXghFp8k1f0A5NQDma+Ss2t6aHWxRR4/VskIcmC2H3k9eq+Y9rS31zqpvBUb
rCGVV9PdDAjuEkK+JiwkHnaV1O6vYBcfmkbiqE9C9nOgglAIRiwv4/E8mH6p1s8ZRA5nELGQdLl2
O0kyWqFQEB8khhFx6UGzutNcVbZt8RZqIqG1/wktJ4kZHregK5MzCWRSWJ6xfPQx6p9pwMmICo/Z
cp3z9yZggw3xFs8ZK5v977BElG6Ry8UU1E1AuSFQUGg2oIol3z4bKlEE1AL3Mecvb+kX5EaI2h/0
IiijvfJ759+6/3+KEwQzfRnmvaOMwAds950WCPYt479joiGI2WeQhZT12U9j2haGDbJeZamZKVZ+
XmnJ9dHBgKnaNy+liWS6G8X60fDVqKrEza1pLR+Q4LJs3maAmIhaAbLx6WF65W1sMcjMPmlrUgri
z5AySR8D+vW0u2Urf4chtrD71lzWhXGjgmTEqvMb8FhyuS8YVCJEOdoYl+RoW/kBhql9wMSV9Qvh
mrdXvLlGoqeXkdoUYcou9wMNXO2ztjMrwU7f1GLjU/ePWRXbEYsgtH2R8qpYVC+E+1wI4RyQ3XWk
TIN97Zp0U0YRc45haBFogKffhc42xPjWP7Wfu/CohExMo+l7LvkUk6nrGUY+3Ro8LmXDwCJJX2Uu
v2peeIOASgmD6ER+3m5O3yfMap5pfo0w0GNHxl340saRxUEUUAxfU2A4NtFbTHdiPYBTIXOk/Kc7
fvKAk9D5sPwUMcWXAymp/o+l9gX3EMHTcScRRswoJJ79XGDXjpKzl8j9cSDOHTqXP7+IgTQoWiL1
i0mmKDJjRcVoTCNi0Om89eMHk7kxVhRx+Uy3vNkyOQyLqUWwpge9CoLjlKoESsv0M9moNzmbLWSF
16dem+0bOYqcJxw6zT0vw+yS5MQfDNEgItCVotvfVQdgRjPRQwhdbvRxC5OslgqfV5kTbJg1raxe
kAbwUh5j2eNcnUSk6YZXsr3rqFgMv35405y276jGMSCv1Db8MWHFD9ZSzzBxhhn+JwabnKupHEh4
/GUB/WrFlWKX6aCcqM7OGC10vFDahwlCf0PUSNhhSqHHv+OVfGtvyYlqwSKbBLuiGpvctivjcKSS
jYNeGL9qlvTZ0e4D+rGtOxHWDm1ECdQhVo56SE8hQ7DpwUNrdLvTN3L4EeoH7n1woZV4a5ULeLVP
PLvIhgTpY3K4py/U9+UtTxVsFWOJ8lk+tYkaRtp13Mu6XQqoPuw9cXV8EyNuNJ3NzK5VO6m21znF
TE2a/O+O1Rfw2DS9N6hd4dyHafe0ep2sMaW5aJ3I6bcstO6hYvMMvPB69u8K360MV0fWCuDJASuw
WsDTZ3fm1OnEtFyelCusw87lRLrVPtb6eyNjfgQ9KX8uAI1N3b8MNgTUPPwWDG9GHA1f7ARuc1fC
eGtwbwJDNHuuFI8c1gE9kto8BkqgwVq1tzChyJT6ntjVpYpdo04segfIHdg0YObZEUDx7UQHDqfC
ZB71xX4ty+QYHKRNSpc5I1RLzTHk6kk6MzdEXLlMzQJN+s88KMOkElBQwCwXiz5T9xa+bjgitP9Q
nFFeisOnV+SgSl9ANkwAYDp6knoxrmujUbLnR2h+vxCpvhiwtM7DneUOa6ZslIOmsYSg0KwCidD0
LdmtFwzJ0/p+AQxQ3K1/4HbjAl0wdNpsHBFXIFZDs3lc/UX738sOoUQFdHNdRVKWAplwo9Dd/b9z
XceWFk2LKKe+JDwnoeYtxzjUrZTbJa23uVApYYm+reylQvipJ1mAKZVdosuJZCLC3Ks+qA5BuJeL
zS3j9mQRpo54TC/TMJVlYIJaRzVaxCzT0CLgDlLbRvHoEPbwccPu4ttxrazz4TV4g8UjYECLdIE0
dzd39SNBag6dIiSWvqiJxRtwQPIlesBA7f+kWpxsjKhkb7BRf2nMnBYGAqw8Xg2yZDMVbkpo3HPx
Ag4muEHAKv0Ze5K7yqnT1dQQgNxO+iZrtnTuIuVf6oRC2/85bBPrttHrq6k3SCeJFcQmAlggBBtD
i78BRJnwYPHqoyhJEpyzYIXpVKTg12627xE53ngEBPGDNRezhVWUANEVaEKukeoIpXJ0QKTM+rmH
VQ3HOT9cWhbpRpk+6XQQ9Xq8St9URr9id9ent/hdYbKExpXFNztjQycBT1UhYA5HM4/wGRR2r0xi
rwscoOjCDJ90ycgnSg7y+qAGMsguTTfkw+5puh310LWuPUVZfXS3tvdF5r7kN2bHtrcCa2Ov/Y2D
ZBvtVrcCvMK0WAz6L/gUFx+umHDYi0uH6eNauYYCOh8x9t5p9WJbR9ezFG0/VMvks9ACtOBm4TBi
UwbHkCldgCh5geXTckC8l90cS7Eju4aMv1R661fvcQAcZqrsiETn0/wwupXjRS6qWfrkMWnfeGTq
mK0Mv2QfqhKmE+77f5ae/jJhq4o4DQ+J1vB4t1GajMRyJbxZuF7uJYpnTW1J7yNv0BGe1fajq3ch
QUXnVwOcWaho3sjylFWit7JTZJsPv6/rjyuNEwIilhPOgHM/5TMxEr1B2JOATHRO0V/APPa3JeAd
7FyX98vuakg6vsiFZIj7YUsO9L956+P3/cGSKAx5Kgx2HsuKu2XBL3NTTavAgtC5Rf2BY14FOxtl
QpcAc+ZfxT47jOJdURvfPmFClYixAdGkEtXI3q7/8pdsyIf192C4IV+qqGscfd2b90YGAB1y7rX0
jd15imBpj8mzfb9art3FA2NlrMUAQOVurJBvcbzHpwD6YoH8xd2fpyEVML2CStq/wR5Q4Y2e93qD
3kgPJqVx5imaE5JPgLQ69O6HvIP5XIs8lhOm9VZcxuRFTZlaovc8iti8SqpY8oDCM++LJ84AperZ
Bi/VBsrWjYAq3PfukhSU7COu5WGoFaWjKtHgScfetOkCjBwPK2V6UarjFz++GjLkzu2GSoPu5Xbk
i9+el9u/xnhbL5dU7cVXaLRfgYfS+YhegpUURqjAePD4urLNXNYwARaUzA+gbHRpGGafwmdUVbWG
6QS8TaLFzX+yCcVV9hGMohJl19bKYVA8BW2EIgrbhKjHnOebM3ezExQVYKum7SibSQvu9Oc9/3GQ
VBk4VQfcB67Ibq88/RmwafMGOUfgnYJa4EWvIrmx6DqAZ8kCtN0bsdJAs161RZ8yUfoJN6YFNflP
OO6ehd6ysNYEwoItsqJhRJiBTYx1rDD3LmqUJq+5c7tquRvKumcY0SSLFiaZdkxQCFsnnTV6yoft
QzUNZlXIdAarMUMbIGpucjrgfsgskcKo7KFyjmNcohQxZNh5U1c2/ecsD79+vSNo541EQ8KZOtSY
K/xBzq304fr7/deLGGbahKd+bKKMQCZKzrmzDCSe7d7MvNilVmTUi/8W2Q+Sj2r8CeqL2dm+ircj
4KFavFxTBP+3XUNYQQuPMbB82mH83o4dBiD/QOuKKfRfguvwI6Spg6eV2e4KkjQESAHH8x/rUhsq
VKpyZSh7x9XnIqlu9O7nk3vihiL+4uE88Hrq+U1581AXq9ePzBvNw+e0DQeKwYTKN/GlWHkWj36/
6P0RPorKr26PxKdb2NsRk647mhSK1xwGmX1UncecdIUkwjjVj1GSx2wZv8RwE5O2pYMIWMeBIDDX
jvD63AQ2vKktiO2nZKoeQAL1nquGy8zHstecU7EjSDjFWWdA6WH6aw8rkPnRoqjQeoudN6W+c0zv
mTzTqRPFaNZB0sEDuZkid8JgBWMlwmmtZn7BLnu4NCi7JugaucxzUYqyQX8D2dlw1JhRCA/qOWWj
0mwwcbJcWgsRIibxtKv2JBubDXkIW1tZfacPusV+XVo0jxeHLpCh7NSO3GZ3xUcsd5GqQ/hv4wQs
9P5zgd4kVWOld63JUyPES4OXTkRDZcmkwxwjFT2VgS7UXiG6xxxLesiD61WTTQau2nDJAjpI9OMa
ILtNd9VEluinyIsQ5psZEV5/VcNtnyWtMgJJgkQTJ/gGTF57CfSM5cCBvhZZVkET+ClqMrkackgI
8ahOIyKJjZglEoBHYKruMN6T39C6ZdmNrk3r/yUez7G5KjckZsJpy03Wy+nxnrcYFqMRVtFEJ4jB
3kXWe/e6OV1pLJFLrNXasxO9VK0Op8j6uJMwY8R/ornV0hnFG/lweAXBTZMiBVSaw0uRlxKDC1mA
L8YAD4Zj/ft9Js5uJjRunZrzHDjcXZ5jYWcywljLg8YVeQg4c0oL4d2DX5NFuzxGkGSPYetZyn6D
wU0CPxsD7MUB1JSI88NpfCwIBB4u07ZyHrsomImynWJfiPMfxBoD/r+1+Itphu5cAKZMk59EcnKG
bCjbLtxOa3nnayKrGGvCgE0ANpYn2anqkjQ+OwvP20msyGxEAmjIsp1RZtyIbAAXF6Y0udT0lF6t
uxQUmeseHSfyKWFknGtLSEUCLZ3bpwi7rU5Wlst+k2HpNBjWsNlELbv5fX/idZOnUnSd6lUG0V4d
oo1mbTJx3I3FUWCk3hCddxkWHCeUwj9CAyqKCP0gTFS3N7X8f9LZQeC1vEdXIcrxYRta89MSnu+F
IkrMUiUJ60VBjnrkZFu2eJ6aDcFb2xyK0O7B6ZIijQg0Hz6adacWarJ0PgpqWp5wCEjp7SyHhMUX
Ij3kbRKWnJJ+rmm34kbqKxH7mrzMDSQe+jF0S7O6qKvFow57u+vNLLEPD60nFinc3nOWEY1TlDrx
HX54+6nez3ueJcIOcZcFOtosC3L4SvItLrXbN5Xxwyx7Y6VOrnFQB0t5/HzpyUcdmrC/BXtEkwPK
z+0PXIQq0T0Wtm269bQsgso0uN1KM7KlBdaXNj1GojXdocDL6Eyrb8XXGv6ppHWCKnYTE6WhOTS2
FEcld2REzaX1XaIPhgVOgnEEF/KHCHvchNv9iCebmQhf34CLJKqTjqXJPOEnH0VY5Sspgn7FZXrn
DPXAuDU3my7Aw4vs9GeADKe3SB//fG2HPWxSkaOkBR1RGsLfwV5saDJCBO0k3qol9rQis1tXEjpA
iBK5Dsy/cMJezJVEXM4HQuqYEid7+Cq0Zbbne1zYdpjWc+HTqToua+sARMhDU5bCVUXWRG+1RFLw
Qu5W6Czh+N2k3nX7kDUQ6ls7KyoUnOEi5cywpROjZf/9O6Z3f5ZMKxRjWWbS7OctQIiHYqhqWFt0
zNLGjPlZSgCADICafvDujxBG3aZcCDOD4bFeFZdkqvGenB7Nn6z11ubJI8U5tkYaKctfLzcSavKD
k/j012MWn/LZRvBvr7LXivDRVjvxB2OSlojc7sTH1lRnGz0CboT5A29y0YYDeVp406/R7tI5bb8l
gD7+OAY955DSLnPVS52tJpu0eFs04ixe3e+akydMo92aO7SLQgDzlhsoOAVkQGD3aIhqqjoWVt7S
eblYwwkecweNLdTsgysug4sq78ch9SMp8N6772a0EyFpfVWUrujgWpl9Z8ZmLvVxHW9HnF+HkJ4E
MXu1oVPrVnYs/BDI4IlK3l2yX++EBwCA/9lDrIau5SL3Ml3lOUdw1Itgpevx8nACGtLmu4PQg2AY
GTH3cCrhOp806jJizmWFtq5s2qWsBUMJArwfA8yBkIEEHnHPmf6wM426qWdZal+24V+sm4pwDr7b
VY3HPq8Rr67ULfOY7j936WXbbVCLo5SXueVtCQ7WZMlVp0ididT6N6oerKsILQWkxjBFHdHzSdFC
54WjcaSn59uFVVieoKkqnT1y8wwr243Krz72WoM+pODHKqT697dC2KlFLQ4obtVY6B+HDnv6FvoF
KcTRoL78kEnKDS3vKZ1oUogtB8s6NKg/MyCCqHyAjWFvmnfUlXhE2BU9bkkJMNBP+xwyYATVAc+D
WoW1QQc7TLZOlnB12QSkIqvQuzlF64r1AfgbaKCJqFqAG2ZtFoLzqI94OJQ3aAaK3vRQIb0fjjjx
99ppoFyvbZiDq2CISDMtd4k4w4csalIImXb6A36ulKmIvtfwpQpylati31+COJZq9mOU4EZZtWrG
r93+gnU6Izw8sVVZi1JYX3NTRBuFiAL0OI1pqBBKg1X3B56K8R2+DH467LOEC5yV5KIhQBxGajez
2pvOwjKvZQI+7NTc+Emxgir2+zlGmlonhUzaDmFcJKUnL1BYZcBMxUrNlioVFM1YsrhNqPh9vJY0
Lc+dvl9CWoWASGyLbdjOZRmUGGtIUMJXkhaV+1wM4zr9OVs9lkAbw5EaZ1tWoSOQvQ0XGnOFHY0q
ArEiuPOKDdTC5QkmeBnbnjOgH2vt8GM8m2fXoSZqmY7ozA18B8DUnPnY2agWTPaAiiGQ4CUP4Vhk
o43YlCxbkr32KVxRBfX1Nex5JkYOgyLrH+qW9N5Jn9eOo/8Ww6aTj7U4waUpoNTIydvyN/+frWxc
Ktyjnu5WxdmuOSV9wKo5MoZBRBLAAbce/NMA9i++KoC8L892A1rQek2MsBXtARYDS1LyPDdr/6kx
ufvh6ysTT6pks2vT8RuY1/4XuUdfhMYaSf/GzypFV405rvlMAgwoLVGLAvjKeILlyfTW/WgeX6uZ
vftr664kMSxYU9WcSJqzmNq+zA0GlUqmQjUpAhMEs4Wyh0rgU6dfhpuGyV96a4map58FRkynt/KM
CZtWjUVO77BdndGXxr8esXerO2TflmemKFd1m170kYZNR6llsmetRkYkZA69B+GY51KZUhD0bJPP
cL7G8LfB0UuO9lYGTP1R19nmEobbDgMwpgnpcYIPZB9OGAxCjYy427Cnz9UAZpk+Hx2WHrk7u97A
YpZSraL/0kqlQ6iiwtqtXH6HH320+C+osqbw1ktDMtpBvGIM2czpb+1Bu9n0F+6VOyzw4+waQk6+
6RZET44J4IYqSRkqbu6HveFMhQ6ZUZflmNWcS2Td2NtvRlZQ0QBWtrhsGkz39S1ETrcH3+qVliSl
BYcim7gcoHVNuq+takYoISSgoEojHsR+rUSi086FEB4sujy7mxFahsaUh43JhZzYeesBxvWhnGs3
VQlvIanECqe+mRYBA6uXxmQGLEpbdxi79W0KYCbi+SaW13I9fxaGlXKY9uibHZJEA2BjfSMOQyDS
vyY0+yhncEZdDHLXOXTxaWrT0aHwPBD51wMe02HEjpuAMJ0MBA/GMf0+/dQdYvGOqSEoHlZLnzSq
fp3JqLM6Mh+gc4Zo3XYaent3sBJIrkheZi/MVPQOt8Yujj3+j3ZzjQiaEBB29+YXHCM3Poe0usF+
rDsT/Kpv/Kq/tXY2K2NQPZ+RW3BVW9kAM61kDZRQ24a/yoPRnpmEiiuV0M5BhsrSIdUjXTNiDalH
CzBm5EjCKiTtzHSEdscpO9rNbCPr6yDG8L5q8hV1j/NHValdC2AImKN7c3XnFeiHBP4XxUdaP0zB
FpwYCSLYJ8il+whe+tjS/wEVe04U0RUNygBNf33esLfYDYdeEfLMBFs/oPWrUg0h1OUuSokDlVRd
GVOFzLLsllgrdm0hml2yJFhwLh9XZ3+6BPRXfXYnAuW3OV8Vdb0qCxwFBTWAGo681YD3ckUGY19A
/D4gyc2eamVqLM2FCbGycLw/l1V/J+Mci5AY6augFLN4+GgjzA6r/27DFuwwGMKP/A4YvFxdZHp5
jGquCC3MtQrTJHW59toccct79RXlbumlOqEjqnPCwJR4eheT+TP4KuYfhr3xAT7Cj4FFt8UTA3dk
vJ/bdU9Kde7EPSFJBapucmxeFwtKP0l1OzTs+9KNFkE19Yic2Wa/dkiBPouVN0yegGaxD7m9nei7
k8UBZRp6NPUQegio22GBo+urskbU4nMgOwj5aadBT7zIQZPHooKYHUod64Z3Mwf8Xq1T3ayIOhjd
nHOHVSg1SBcBhp+OVOKDartQ2V4eQBdKGhFyJPFual+5DElSYBHyxO6vKElhdUI7U7SlqjU0Et0t
5DEZ5XcYukCzdMFtS67pI9O8htB1f4DSCVfifQ3uQV8W2R2XiaiVa2AsErdjZ8yYpyB0t0qQaB1s
bYXp/V9M+RCuPoG/7S5j+7YjjMlYj3/aRX8gC4aoq+EKtxpMlHLsK2Zgk5Tei8oJdD6lbGs5OW9E
iBYfAHjNMCaewx58J8nBZrMoIJsVuDbxa1ni66g4BMPJVjjMaU5U8iRmxU3dc+pQ9aBP+4tv+Nex
47akXmAHmbGq2T+9jL41sYcfo/s/yV6MFDuOEbqtONX7nOK4Fq0qRIsPWuLMm2hXctC5Gn2uVMOU
GhpCap7dDTeQQYg2WcR75A01j8Cyw5R7PUZhfG3th1EMIAFaHbKPuApO5JMLF2vvZ4KhKGDCD0EI
qSYdS12y+m4ay/HZPvC6VYc3T0a+v4w2NrnlMQ6HobYHpqu3Vj7Sn/06sM2g2E6TRFDNu6n2HWqk
2eG6uNQNZ9v/HkYY+c26LHOM0c/FR3SajwOyeeYWRo5qeT308De0ZA2hkJu7KArEPH0BLvQ763J3
mEIpDipPlZ9PKN+9pD699CS6Hdk28NaqndoLzjZXfc9npQF4wPBPFD979PNfgoQqs4vQ6mElnXbY
Opjt8FVzwzv/EmhtQOQ55UeS4QD8gJ5ShmXeTf6ZgVkk4lyYgi5KFHhgRq8pEK4ovP5q9zRPwBHR
zltzkNJDI3R5cVp1stSiIuHiYnNm1+mgy/vtYR7CkNWhyDgcI5G5L7sgXaEhUU7bGMnKnIS7Nwqu
0x/3bm+h1wrgKDmtUIgOG1VXzZQPjpraw1Dhpu20jsxRG9ivgCkyuALkaP5iE61XG7mWDdRpmcrP
Lf+t6W3FKgQ2lQQgkyYPh0quyQA+8LXMu30a2LveCHRAZnbocW/vCTvKHxujTuTdIIyO6Nut4xT9
qgjbZjGyB+nSnMTI33UY1thplFo58dWduay6VjvVLH3tz80FfDK6qZSd1qATHJDHQ5LJSOHaoMrs
9N1qMhZ3a/csRU2sOIZajuac4mcG8pHF24PSGHJpfy1Mj+LOVBtbD8Rd+72UhjrPY86VTyC8Hzbw
7zEKmOCljjTDk6vq9vzgMKXEeOrx6gkNHT6X/0oxPe8EjdJ1mw6nDMwzZE5zXEwjWEf8OebHFLoR
qzdMT2228GW8QAUeDnTLGzu3l0ssj8Q7QEihU9XKSMy0yoveYsq4RNOwmvU1WqB4GYkOeumd9mvv
hi/6kYqFW+DtsC2HqvQu2aEVpycRoe0GGW80j4i4aavqmWyVKPkAMtHmEk49HSun3u9bpl0MVjCs
B1eK8hb7lG9OIGCZse6UzAEDCjhE781Dle8buGQuIPrVPRITLcLw8RPX5dfXovdQnsXEbKCnhdWH
1uIP3QCP8sKVlSTocmoEm1TVgdajRnASZFgwBxHmfpEF477wr9zwUYqDeOw9+hb7aMGzfavL8ZSB
RKSimKVt15dfjCyZoX+zcjAwwGDR3aOcCijukODx4EFqF1rvTGDW+mMVxwclbD4XPY5Nj7euVnLF
s6RXWKSZs4oOKVCF9WEoBwqPvqehJ20dWF5XrGxqxPKBWwHhLlgSlfWonCErClgjEgSo+srsCYQt
UubC7ZxVR2e20SStR9ZfwMbynEM3olSj/Zknck3TBhvrztUeyuiSWtGlGnvM6nVmpef/QZ3EdPGe
mC/PkU6+F8RfMlQSev+YxMmHuKSJCR03MAqZ+FFR3tpASTJzDgWU1jgomHm75jAQu4v0QkfHSR+J
n8FRDKOHRTDlKtXAPhK82rxICJpUGym8MYuzBDw6JhzkjQeYc00aRvSVLWYOPg8JjUzmSfLCsVjE
nz4k/nTlMelWj8wzUaUfbUh1pCfl6HlgYnORiVowY/JP/WdFJfMfLQ1niGeS3UeGw3YEI9cVcf3R
/YF7a+T3A9ErPSRCd9Q1cusp0SZFR/upB7AxnFxEIU+hcl5mKuPg2r7Repbe9FmH155+IcJViKxe
esgeSuRThUHsDztn7TaHWPj9XpOGgYaWDpvuyVNZCB2L9FYneSguSV71NqBsmbz/S2by7sYkGRxm
9YbN4X9VxeGb5scKitdNrUW2hX4XU4f4P9hb/DYFB5iK4evORA/2LldiTcTGWGdlj8NIhKRvXtFU
hogVqXXgHQCfq+090McebxJb62GJ8g8e0tfM+ZKWJEGee85/1inLmbM2zNfQCQQHTzQK0ewQi2fo
E3YsLf3MSCkx5BfWE2fmi+fywCOHY2kOXfEMvmdcASHC9QZbinrk12PI1JlFsJji8x9BbbC8NBje
WWRG0AugCB/jobujoYzowvPTyAQkkznKBCoWkOagXsmwlx5iGMfdpx9ZsveKE+v0loWUrzx4RENg
moBpObseIhU/lmKWbttMKNeA1lATkUWOKc0W5JIKKGXhydfmyUmsvjbTMvX4RvpMyBv+rtrE8efm
IrrqR7NBQv/FuXfSBxUTGZs4d4UN0VjRIagrySmf8ZBuIhQ5FZDjR4QLjAiGPNtgnKuRctuSwjbx
BomZw9ge5XC/7S1XJjHKr2Nwc/gxDiV0RX7VwPX7lvhoWxvP6Fn3hi+CKZ8rg8JRWZyAbyzEdFLr
AUIVxi5UoUKmLIX027IMxw/aDZdPJ7LXgWWQKFss+EFTnRGHhaWAwAsk1VLmHLSCosf/O3PpXonl
rkLnTCiUaNofvqeMnoYoz0lxCkNcQvE1amunorO/7MD5YluGeCa1hUSCqgbHvo8ye3u6vsRw42MR
Ntzt0fQZdnblcWHgPRYRn4UEBahGpfBAZBmg1bJ5anOqMLK5sCX2VDR5TghCmLkMrSmRFY0shax/
D1WABBKyFE0abQpa5k5ep6EXi4E+5DThOzU1FZczUygR0YLVJbl9Qd8q1s9SP74qOyE7Gh+5PAcp
PdUWRhp2SNvK+EB/4LVMhLb9cb1ime4FY9Fn8mr0pj0iuv36s8AX2c+ZrTyTmwHQ2yWcMGtkAXQP
13soSQUZcxdIrJ1OyUNk4p6xAPvtjOoH2a//rVt8tSCy8DqHtwMDZhfKt3lAQ4y7n2CXwn08FAci
jVGeItUBjxYyLfVcxL9Pz8PCa9teZppH05y4GeN1tTIb1A+yI9vvFYjtOwtXD10wVQDZ9mSb2D88
nxwhohVDSpI5tlnJW3IhCsvGkMul86C3nebU1QoyShoOMRu+NSHus4cHvG9Tu4wbU2y2Z5pfn0U1
Ij8MPhe0vy9LiX2nD/AgYEK9HreWwm/m/wR0CtgBq/SKLmZQzfz42KMslvINzQW+vT9PEtBta8Jz
QnATdH1An8so5z9U3UpM8zG25uXlnSZypIyNZ+SsPb6PJ1qQGaS3Y4RzrjjJR/NGFA5/r8JU3/Su
QOBwku170zMmf2hw7+tKTqz6N7w9oyHsvTZSj2g3TYEqVnjuptw+gDMOsP/jdnDs1+CLwJ38WsfC
rsSezXkT7BOe7sg6RqlHqFhOO06G4TyRFo9myiT06tLHTkmtY95HuwaI3fdo83y9SCK1TQTGazV2
potqhK6DHMZa6BzawOuKXZkXsa8tVhwuP+zTEVpHQM7/QSyQjPab2nlOn0El75SFfq8froQZJNpK
1n37XXQw+BNUSIqg+h9mXGXM16QG9m0ExrJYEex46odS30asAnyB0tqOYCaRGGf8ckrF7cyIYdvl
Rq7NpRYtmxg8i6ItghSulT5pA+zR86bIfMzm3176oowR1KZ9a580koJNcbzbFWwVyQD1HsV5Ai+B
dmWRw0G1Lti2+PC9tppP+lpSSuK3n4g/uvJ2UXtklc5V5uL+Y0twEwZNOt6cFc2qeokg4qgNINVX
S5ddHCqoV17+8NWTlugbWZVEn/Jh1SRw0ZAeHn1n3FlTuzh+8Dg4ihiG8QsBAbM/ScOFB5Lbvufg
7+MC+3ysoBlHQgjVMXC25cPC8D4sYQB8353sFOQg0VT6P2d4KFslCyPAwaov+A3caG0q/RUkuqBn
f6mmTlyT8NClnkv8OTvP1zdC9PEV2L1fZhDgnx6nGPIsnX+nSDxQwiaorjHa99NevhUETWrxswfM
fk3bryh29DomklUh7JHDbkIG3yLuBKdzBDp+8ndm+IxVmPN50Up/OzLQ02U+Ftas7knWC6YBpFN8
An7cEPFzaeEucv7XSBdRDEMgAKNG6Q1/kRrPd6WV90jiPRW87Lr4/aeD3324FQndCsLaue6zZ00c
y8t2y4dGK+3SUoQ601nMyfyGpCsoSlbpN+iHAZ3SvTMxlmbRtQWagGwCNlUTko3kmeozzSO7/oQh
tlXfx4d5E6CVw2LhV9fJP10Vu8qW20J0ND2DJpobbIooVl+9OPtMfeuaYtwtdCCwfvARaCsc4X7F
FuC7t01MN6kQbRN/6t+xLTwGy1utUtw2vi2MjUgXRbwf+2xkgu23ZitVZyFFBKt8FQzzmccQ/qWa
k3Kjg7xjZD5ODdzKwogZAy+pynW23Th0vE7u0JTYi/y9YEFo3oZuAy3CW2LM0EcffWgrCEbU0ZnZ
uIeKmTP7Mltf+V5zThjN2WrdipmZFMpKL71e/Js6PYS3CCnKDwDz8HnnM4CIEfC5DaIQHNql+ARb
e+lgA9BtOZA8s/T/59a40TF5LDKBCQBjoG6rHLDJmvR3XBSoHXkzq7Z3xwew1La3SPXOZWgvl0nk
N4Wy6eHALL0kN17Y40K0Sp9/nwENsGcvo49XyVq9j9rwU6YnMRsB9YkXU0GDMiFQg6UTpAYt0PhH
NcYYXd+FkVceqRYt+1Y2MbEkEVvPBaPrNiAbchzXS7+ZgfwzGtsWq4wZY9qfM1VoMz+yMOoOdxgy
gig+WjJFOmN0mwq4ldjFHMEVSDIHkdvSrfSE+QcozBvPKr3+510Jbkk1S8nqPumC0dYmOV1aahH+
ENXT8sPunUm73BZCf0sNE6+zOUaorEr4zPnVsD/8y55NmZetQSRTeR8060fw4xuNEBLL3UiwMViq
wsR8ugnu98JyV3YwEtQt5sn5qScLlMQrtYGixaTT5kcIf8jejz1OnzJsatarY69FllqBUQXe1vzN
FCSZV63/gt/Gf1I8cffANVUv7W6V2pRWjPcMK0MeYbXHXSYfL0W2Em5q6RhdklMzYjEsyb6ukqrv
Koy2uWygr3CzzkDIBt7eASmTebauPKtapaT54gWLBHO2uogVIWRX/MK7+gQtRpgg7ZsNDI8unfxK
yscUVMzS5g9gmYQmG1Bz9lth8pLYHWHi6HYjjw91dVOC5Hv91SoH3ILZkrPbs9y+DGWUN+E/CQ4C
W4B4xnMrKuivWKLITMPsA45XODksBfLJGhIvPhJ6bjiG7z3AeIAZjBeBu4mGiqmCnzx++hRfaW26
SmZ0nPoRe5YXrWUvSNDFdXvQJUVQb8FHCjMHMElWM9O43O0l7rmyVu6ZVEAbcNewjJHRnF5iQv1p
A4+JKC+lWCLPSXxlhacVxrqKWtq6E9/gciW/4BWcmH03H8Xc+oox7mqFa8gIlMKhK00cudeekaTC
b3EQnxiBPsyTtqZVJ5twKcpQOMNsDOLcPF4ccHOldQLkA3h0Ep7rytwIZ0y34Aq4QnlEoS4N8hTA
oD4wKCkFXdPdo1DGa4D5c64fBMcwAox+sL7KjWYmQCwqr6g4lo+BkoLWNrky4zN170EA2T6dpNyA
I3rQSUVyZlc7xfmsGzviQxtKFwYjhopRLhpYIdS9r2r+jLv+8gVjIHLb2QQWqHNk5wgjsENWmwmE
44lj1TaVs2oohFux4zwIUWee4sjr9SMBClPeTsyqDMkZQjX9jC7M/i2zM0YRLmRu4/5CTVFCQkPa
GDpfiw0krAUkrfDKsTcdVrZwvybqF0nLT/iaFqss+K9mHMrLEAEE5QUn+1/Kypag6T006R8xQE5/
VM3ITTSevSgnQFx3h9RaNISSTwXfaKOcX0aaGFaHPON0fO2fb+TDC0On475YYuwjVLeQiiFwezPH
TouqQ9P9YpwsI/GGmQV9to7r9f7iFUBRdLKYadxAXPO/+iu3XQJOF12jeaDHydfzkaNCF4GmniOA
uKYKB+vK73Frg6feub8pbTHv5OBDT4IJMD2tTiQqz0LPVabVwWETruZX7+FRwo30aDvTWS1PARTb
CtVX20SC1JGRpUAKwBMtm5S2m7EwTHOwE6ANRGp4JC37T2J4uGlpPOyCKiwPXTiknBAys/bXIvgn
Xzwf4ea+5PWEjLGdBvXRuA3/K5AxtOi5lf45rwgsic/nJFGp6VEbaA/OY1Ly3wmr8Vsi0UUegJO8
btOuXL7a1/eYGn9L0YIsFZI3yo7NjrCfE8NOfN17sIwaErSUMPa3Ew1gxpG48m7kqUfK8Rzl2pcH
g8DVnHuEvWJX9U9nFYAbjEQ4BzrvuMWxEj57thoTi4iaxP+J9LBClyopSflhlpudVV9R0gSgRMHc
VwIBEM4IIeS9un3auDxQHMfFPUyo0KARUthLOeFj95weZrvOCRupfrzKR31gU2Z8H5pUWzdUFIGa
o72ByqWY3sC3iMgGggCSg/9d7fvmBE7CeGBaG8C5Rd36yzdwFhrxmueimUE0MiDRNdYfTZ0IGwqy
plMIstNmbsQARNnRepvKg3qs8Ho0Lc3CubgoCLkdFK7oILHvYxqFC7tPnayMlWOutneupyqK6o+7
boaUuyNyPXKmEIqG58ttbg8344TGogFE0hbIPo7D84brDj5BYQvykib4iLnIkIuGr0Q3t0KgSEDM
tcVEJrkSRFv1T3qG5jY6EQImSyP86BxAcW6RfuSpcIgeUhuKW5VyuXtjdSGnioZQS2rT3R5JiF1k
hiGRNE6vOQj6WHo/c/4zgACrwF3SqJ2I7YyENSQkUaQoF2ttnwnWPgUtzQ1I563WWtXduQ1fYYV6
J80bU1snLGc41Wjg5+p1K7Gcks2fcaYmqzVpykQnvHwZ6DvvOGYK5nXi0seb1U8xP0OamXauufuT
SE5sRhyNxHpzOhM8fAQBfgrqyIp1WDeIfHgTpElKLOEg41Mp+xCL/vLdfwF0OyUmqiwxI0CdS2ug
oavjosbIkQHJbyLPNGkcamRx3mmc5EipYKJskZ9K4UlEFil0J1lyd2mdbSUFs2o43sTDgqefjB/Z
FG/UWL+USIJjYmhEb0jLWjurbQh7gVItHkmBqDiIN4slkSDW7eBzm9WugiqeYtFap2TTx6MhayC+
mscjcLJdlNxYhOsCOHUb352ODwH8CsPSZ5xBlBwpl6Vd2nx0VK654FxWz0/+mSiONm9LY23mUIGL
ESBhYzCPq+aSgcEUmmzFqPdrgKXEcGSeJf14FsvqTMlzHewMWszXnxLp2q5I1zt4uGKtNJ/pGoxG
JrCCTzy/JIFa554bjawl8+XwioRhSrTTVkuUynrnulEJiopyPZ7txUgbGe4vqTCd0mqpzBYZLNQ9
F8Os2z44DgSZ3QtExeKKIZ4UkEH4yaLDQywsHizTerYFBjKADqvaOFay0tGiVAUEkv64MzbPzBY3
hdGe7GGY0pNWFAYnLwS7CfiUiYODzuy9Uw9X3fKdVWiej3Z+xNGnF1BKd2gufhJE/5HRTzE6DobY
6rdXV2umHxsm119U+/IAxdA8A8knTsXBUt+1+qWepMtre/d5GP6mfMXtL6ECX5IfA7q7zBLvZF4q
8p9754HEUtDCizWa/Z65//5KnpWrbsN7oXPKDiIlG+4UKIsRKXrSDOS0Q6+IrRYFtCQ6cdrhQ9nf
WoWgncd06ASBLajuFtER0LDZPu5aR/AHVUNtN9PWLIGvz9Tw/R+P2DB5rUAyO28PtOE9KwKbk15o
uFyr/uljWfLTdFmzLfgUG2h++LcYSnHmljSSxW5Zjhsp3GwxjT2W/0sTmzd4EpQPq6kYAOKEvRwd
/BXg+Je4O+nQ8YDg8eoV20DWkbuyELC4G1XZ9BAb7t5RMwDjHhngqT6TRUod2Ju4FDUOgdn8hC2s
SToWaSjKFM3mytZlt9Eas7OCcffoex2aGL2u6mjRVrfXVkZw0E1zG09TRgyCcFxym0dR9UVNXKrj
3cmf+eraDOs+YbwT9KqHioRmcgXVGEnGZsNJcNJ2RYA62hSd+XhNfHDOlHHEAsD8VsaFR0/wXOtR
nY9ewZhUGGNTRuW000GE/u2I5PWmrJ96KhooOP1Rc+27qUgVDx54HLJp6DNxlEoqEBReh0qcKpzr
L24m9S0VX7yFPKeu1c2DpQ6bTjTh4W5PTs6EcA4vqAPBf+4f1Xd999OsmUEcPZm6dY0hoO2tKLZO
KlSvFpsKOh8uxsZcpdPvjf4dgUFJPhJsCIji4aKrgdb8Wv42ZqEazQ+IErecfyXnecFty03QtFuQ
fqfSVKL8KrwzZ4WFMb1hxCxqHYEzOrA9ZZmyaJUWR4Skd6eKGTcKV/GHsF088gKPx+4DoC6wnXk6
c+rJDVqyLqOT6cZHdtQlMQJU4zs90gIK2Ltu7BdcVlUlpT7KoNEqPgCGc6gzQ7yVXx7aTqgP+1rx
bhWoPYsSPpVNqKoG/LLgKZQUP/0bnuclXiZEwgNZuOB/VLjqU0/EGYN/bdn8R+ZSGgp5cdABq17R
20YTZM3RTZp2H203b/MZbO3QxjvqPBTUaGfUFHaRgjuJCtXAoiiYn3exZRYWzzMDwc3Csl9YyqoM
ZtZiqja4JENyj+RDqAntQnJGM2YOAl5NB75Tv/bBOhCVxXYTiz0hEz+kkrr8YYwfCfsahpHjgSKn
wfv7AVeJ8gY2AcClZGkXxIdm40SnSCkGcpP0YV7ic05p5AbIp2zcgb9H/0CZPa6TQs26Ok+QtDDB
C0+sR8Pwq1gyMOjcOt59NO2q3UgXNbxOw7jPPPEwbH6IB9YdIi++MluOEUeqE4leg1jwwx9WTJCQ
tZsLRngXPx/k6w18oMTEz3veyAi8dTWsp6E05z+TyS4UmwGZOodD9mIO/9SndzSPm7JOJRpBKr0/
OhmjqX3u8SL4cQBFNtpgZTk4ZsetDpDHZ8eAwjvJEng2lUMKrcZgILcHSZmYierbGfi6vniHLlRt
Hr3RHPK0KpuUax9rWoUqwCDDieFHrThrYT/+3zav/YYmto9Dn9ls4OnRGuMq1eNbhm5XQhXFk3mz
Aduuf5IKplIz5GFkEMsl0bfc/kG6Jun/zlAF9fWArzytPgXzGDWOU1iJ2SdUdDhDmSETRj+1Cq+5
iqdjd2EoEvqIXJXLd94gUrcX3ZEG26ToEhWw3btlOmTLWx7xp9OnZ5az7pltFWJfjayEfEHkSTps
myRMT+fFctyVkPejCiBneYe/6vgV28izyw+gHXHw6L6sELaUtoCvDZTy57JDEI9dUwNQUTP+JiXY
uQ84GW4edbqj0s24NCFCrSRMpRqgTprFSakTWV8NuXrXx6U34xWLkGtwOo1eSY+An2uzE1oRp8W2
L2o7ob8qMX8gBNdTN3ngMv55EfryBK4NnhkLaO2r35R+EhFGwBsbNI6mGx9hMwrV6SiTTgy2H43W
M1fYZ9sS+Wd90C/0cxrAoafJA1QoTdzdSfa+HTkjMbF4vuvrYTDbLXpazoAYclsxKI2WRxcOaNPg
sUa40GGvorxSIieHj+m3uKo5cq+0xg6CWz05nGoO+f8mQcx6rAFAbq/6JKtpuxfne4cxYUrODcXC
1p7Ikb5bXdfcJmjbpmgtQokkwLOKlXW/Xqgla6H1sPUGWM22fLVaJp/JzwTa2Tx+ZgfXAnD5xDx0
4bCZWGL/G3h8udCzffE1dX7xiuIWnITBNITqtFewqc5R2Fs6xaIXsFKQdvC61ZMZWVWvk7eXtX3J
GKmqsppBmlOW2cQ/zSCRyhASZmKLwCGzWem1Z2L6CCdTqvP2gk6RPibGsFcp5LuEgFR+zh7kbxIB
GQsin6TVHILCdnx4ngwcDpbyXbJTr2VdG7HlBQslCgZje1rqwOz2gpXytaIVj60aO2hhRqOtUK6x
4nLLfglYXGY1eZvvV26tNMy2yM0RREj9CZj+dZEMPIRog/Lwu/rh0GWQkKxhJOHsv+fNmOwSfFwj
zlvN2Wacfx4SaDXHXIDQi2VzzIJX1j6qmwSmTJrkY0DB2Fh23kVx4zJd0Nspu6QNGo/aKMDH7rmT
RzP4CgBokqbFBl3HauuY4E2GjSVUUlwpxmRqGPUX8OhNRj8QuiT+CM3gBoizhxGkeZa/dotr0/lF
X74tGeXyONY+vNjgI1HDne+vknaBZwnchYhJ/3bVbSBp31YiYLpwDg4rI+oaLp+ITXWbRdffIXMr
8wX5o+fThurWzEtoPbLXHjqh4AchkejXSCntILKCaA6qMZ5XDaQLAimVQ6mNEXzaEkX5cQSiiJEA
GEFebh++cSyS7sOBWEtBP3bYIj2y3zccLHD1mX/r9PM4X16e33o2knW+D2Gq+GeMlPkm5J9k1tBw
0tvoZHe6eMNuQofh0091FfxO/6lqCBwoOYEL+LhozzdN0GLSR8d5k6D9nMVEaXF1d2pMrWWOUzIE
MzczNTZMDwVFeUDJjPl5hWA06WtI0b8MxFSYfEJkjBRaw33W9C0Dv+epo1q8+UFrIua2CGUGvLt9
FX1bL6bR0Q74D4It6KNFP++BTmpOXz3mN7N67/mFq2jGSn7PNY0PL9swgggTbFqIq86GsJc4PA1x
xqmbF8+ELiOeZn2TEJjfZlwlPnQ/LILmYUOTWnD6PnDGsRXFQLk//qrkMARsLzCV17xFrlpvZCcG
zIT3gjiZ5cgb9A5YdLvWm20kpLa5995V2rEpXWqEq3MSSxkIK3YdWdEJXfw4kX7vcHNY2c1r259v
x6MDkrc/UPKRV20mPXg9FjgFMBBZnmkLZ1J8T6kJQ1BawYW47BcdxKG4wdxpN9Xgts/x579Au0mK
reXhCSwo/3IobyrFA0ir8zTCYiv2N8LdknAmRY9jqX0qImHrucFnuE7JsRldbj5S9NTpu5WX8JYm
zu2wmKvLQ7hdm8xwssmtN1/cr1Bh7o+ya4Ur+sBkTE3VS8Ile/aWLvYbzZ/aNroD1eWuvyhjWBdg
m0siv9AV0ATJaCCDCxYkvUG4M//imDYlMBIHRB9PrdmwUGaz+AsvpHHklMad3F9o722gyNqdPQ/q
SiMsPmcpdUszNw+0F5mmwFlIXPadiyehEHPq7I+nm1/7yI/+I771l/WgpNa36hBzXtdLbwqri8d2
u8XfIDMey9O/CEMibnWl+N+Ah71NiwsOeeulSAXEA3435krprE4FtO9p9fpggcqLfi1AgFnwLkPo
blrf5wCqU/RgQkLYkHXIVXJxxocPvwXp9zDzAmXxz9AQMbBfHhwx7se6Ge0fGAx5pdj3ndxK2ukg
FHEs9CASCTclv5EwnUjegI7i9Xd9Do/pwzulpTJvTj40U/lVVcYSxQHfaPws+K6iQ1GzFG6+Tec1
i0ssaqZQ6OuUeU4GH9Z1zTDcGpKp4kgG7tlDd4NMX7JfDk/2ME86+8wFuIwLQHVwldY0lY6i3oku
qbIE5MJROG5nB37/KN7JhVkZlGHyWJlhP9IjBjx5hDjSLBgIiBDo4AI1YeAvJgTyKUNbUCanb2ez
dFW1fgrrFrHFzOf+tCaGFOW0UqkmUEkMtr9iCIT05tlar35a5WO1oDR1Yee5ATC+wctsPOeN1/ob
BdmQbvXKMyEK5IxRHyQGy3VmASvgR971ng+jJOYlK+ovRn+AHdPBGXDvZxBxZ/fiCA5clqGengfT
+oqpjOvBTmWJmFZWCcISv2d/LLNcqCzRyC6S9pqJ5SlP+ybKzPBkFz26OD1+H4ZqjA21IbZu93YO
zIkIIBtdHnPy95ZcYbs0KkhrHoU7yMnDtb+V2NLICg3486JM8d11U/Dv6tQxiak8Iq9jEbqW0rmP
wgvA7XPI7WHETzetOH/WiaLsQU0CRndeOa8eyFQtzQjTKY8K+j1HRU8yoq4EBo3kN+DmlYAPplRC
kX75H9DZTPFmI71+mHw+T3rEtoLJlPU9vdrzTPSHqhGgTmXJU+f3vMJN09P7k3ArQ7gD+/u5Bk20
E9sIufHoyXwsE9/zyWhASTOcQqb52Dgcepnnd/7uTs2clqGq3fg7Nr6juTtrngMnmECGee7/f3ug
4ntsOUAIC3GQOP5Cui3ky9EDt4J/UV3cq85G/12cY0/03VlN0vELUFlmoezIMV4bwiZizeGZ/XOI
xD7IMO74088kvGSzlm7kRo0Ut+2T+mY0DNguYCTsdfez/I7VERHlS0zElfLwkdPc86yCw4yDOcaL
9mHjhRu727+xUXTJQeW1ELxbW1lkTfdj/SeFKn1/SL1uJg4NuvE2TkISppcK2HzRFt0UQ73c2n6W
DE1BKuY7yxXK6eTzc+mMWACd9Q16TGw6lCtsPrY94FflGKMLkqJs/IGoyPDNkbRoiDagBuD5Fle1
bf6GPBnf8g3NrB9HCzBWIS8NRVn6b+orw77OgPSPKTpa4vv8pEwQL5iaVp0UOB67/6zMdthRl6tJ
DKh1m96M+1xCp2c6WlP1mnSKCb/I+vGq8bqynyXCUDN7u0qRGovJliGM4KHk5oRcOFZA1S5uVLPj
CleizZZVPEJSORFvA8jt0mE7mi9oTy5FIJrG0rwHWjoPLhgUs5JA/vVvaVODvdAoSJ7VNOjXfVAP
Szghm1uWMRmuJl6D9QQFB/DZRRBf1FrHKgH7Ee+stDgsQOBoatfcTqEEA/roTZrtfah9qFjpM9UK
m1uo1F6cD8ToPU99eLrKELPTLdLo4nlrQe3Dqi05SS5+VeO8QTIoEJIHe6TPSIRGaqDf2Z8ZWl8Y
BsOwPD6oX/D/PIZBj5jzqh1AYooYnw1UHXDfdM/JNZWGhuH+Vzev9Ar7mZp+rTPhkaeBK0EViXOB
6+2M8Sl+OiSEq7cDYJtHHSzx70s7UEXEssYNkz22Sz/53jvjdPo9tRfB9a6SBaMabyCQ7WqRmQKi
EZTYujNz7/RRfbmC+iSVGt5YDEF1RNimUugVSwA8BozYdTSg4O2qgdIxLVP2cG4kupxRgEtXjwJ2
n+3fYTiQab1ITU0rfP1UiChTT8g+UbVb3TZKo27SiMHXyfhIajN+99SVg7gvvsY77UjsPVkRCDlG
uWY9D5HSmxKHxH9VB5ItLkg3884zMSFVctaNSbno29RCeEn0rqVMdPmHC88Aqy6jsnuunieKKfgm
GzhlfYPSKey1n+qUm/jbQ3Aq3bQp3wbI/M8vl/51Wfh04bycdHVIXGR7xkeaJFstzmOO8BtZddQI
pi+tUl2KhDMgjwHYS11wmfHbHB6QQt2xHG4wB25+5pOpUL6GE9xTfzFD1GJs7wavqKzWU39zM/CK
w9wO4aeKqviGGcL1SIN9TBbQkf1XJf5Tghw9P8mAA/WYPXJ5vqCOX7UysdE/G/6yiBx5xkzrL1SK
Op2cLfvY03uTDDl33bJAkyQyBGgKvekqjXS9On6yC4MMMr355wkpNKtJG1XY0g6yd8/qHKazpWv4
GFjGjgpnBvvDTWzmTL1OGgR+VSrqpsu40hYbadkSxcLPgzhheAcdpPAlECHTTHjmnmjV+AWAtXXB
8MSovvvbYFaoiHLMryQ6Ck3ZXNJpLFgsBhS1BqVL6rOK+oCgdGwTzbWZhd8xlCEmb3VARhcNaF8O
k4tAtBg3PqaHZiwT3iqKt1vYoeV7bZcezwS5kA4mjMfjQfHYLuu2yryZcPnyiTvNMJ7c7AmxXqx3
DgG/8pbsa+7HPSDIhg5wC9ESebgCs4D9vml73FCsJ8hg4ar2+z5L6ZdTKiVJ/LAHxGKa+WKndjUf
gA81Ajc7msUWWGcbUTwgA1jM0QLyxNz2GxBFiSC0atcFa+vujXQch0WqnR5FbktCWiBcOY3cBfgE
3BjLLEEJawPxEihPyCQQ8e0M23d4xzEE3XgxJjiFTUAy6zAjWohC6TvkUAjCE69mPgfhaW/LgAld
zv9oP+IzoB6VESIHpC3DFBjuD/Ctu7VpDmUpkNjqpGP0Xhjr2uNwfYk4co9passW7TFazwdu5axd
8Q3Hkhp3F9jAi/Avd2u2gUPHROokbLb8JkODdb+W3YDXZAYCySdElut3j0k/A28rtMUlrQtJMkWu
4f2/X60qotuS4TxDsiGsy6nAexvttx3px1zI231SeofERI15vDdaxi5lndGQACqneUYyX24Sj7YM
L6Y5S2fkT1xCd/Oe/GjHbbOjyrDeYpaUM4Gal3m9CT61T+K3iUpAk151qj5YyA2B74slsflwzY0z
toZOsayW8hv5Y6sYU+0tfKZYCk3nmUSY+IeBwYGeJqvdxpEl+hTMq76kka91uxcJJcdInt4TMDp3
0sTnIjBHK1WpXLmKmCVJ2LHCcsNV4FmHKmJ2w0oDh09liFi+aBDNs3jGx3vUgL4XSeYVuBu8twCr
Q10cm2OGnsrDdqaSnzlZSBJzEyZ8J6z8A6qMPjiFEED+taX9c42O0tr3rTLSacHnUfn9s3eDYMwr
XCmwfNm541VDEVsf1vAi8DL47+sSg/3+nrxBBQwRngAXhw6fP8IieASmXBMBzJzmTo66r++6rqlq
WhloV/RcLvk/0LFXPQ6cjQHoxelpK2OAAtkZkjtl8SzJWJU1BecmYrHrPhAInaMD+xI9nt4CPAXN
zJbagXt9IkPbkgm1u4+TY3dM9PondpbkZrQzAN6AblfKf+IUpAlkSPkkOUKlStY6SlKDoCC4u3Y8
ogBnxR9Mj3hCm5wPCpLYlTPekrUAhuaRmYtbp0VWe67HBmUn3HEtxlc6+y7361Fr68CefSy7KJq0
LpMuF3FCWFYvyP10lSLnFMHu9TVLDNUbnyf5k8Fvi5ScV8TyjCq5qB4SI+EIjMS6N9xPibU5tKIc
AWcAyx3ZAe5U8Q6K6TtMqTOPTMJR18CYkQGdq5dBuBUrGbtuROvYgtQRW4EbzzjJcaQNDOGxT1xc
bNyWs6Ikj2qbfxFB2vxQ0cQldO9JsmP0MHPGTh1II01Adb4qlBgx61cRBFLlspqpj7z3QEUBkIEZ
LY5ERDfYNYEn8eAzFD9TGlJQdAaL80VD6/tLQJvdbwkq24N4SBRUPurhOoVOjxXfFTy5FL6ApvFX
Fh22++FVJgnxp6Lmpn3Md4dlyUw8Mp6LPpFrSjJNVoLn2E3lJ8QXYFHa7ZKnQH6LF62U/HI/3Hot
2umIDKwPfhtKmnaJ/4/d1lnltSNexFXgN6bKp7qBHTZQGtVChx5mlgVfKH0HEuZW3BFGfQbkKkJN
74J+4j50KQ8DWRcw3nMq6l+FvNSZxxyEzkb6gZzDE9S2KXzmq4mhNxMD7tFWcaQNU2K98bSpX7pz
vxP5XoHSGuo9bVYqEjhhv1gZLXeqIhkx+Lm0G/E1PLDBjYboGCS30Dt4u/KA759NjN7FBDxSBkO3
FocSxKvFEsuo+X7hcGpNaafHKocbpbIvVgaE3UpkLnUlSZMhNYlZ2YKqGrUVZDfrCUUyHnqlu7co
fYwgRDxRoPHKVDQIDDBnWCLZm9+AeIWQ7oPNrVPojJPy7zQ/l6MrQbM/RmfSg9aPFf90Ihb+/VAg
ZCHNANwOnhr6VwHKpM8IRKHOFK0sRwLIn5s+BuyZesl4l3fDbs7qS2hcWVgZGXPkqPhq3rAKj7hR
u8rc+KHbGhSXI7xlp5V6ZIH4F5nL5zyudpIM3BUc+rB4bfdJ5kV6kSmfW0oxFFHyMVV4Zk1K1f5z
xHA1XJB/8eJMuQwJL5iXZDMkczQfp6T+GI8QlheKgCovgC9hxbY5x3aPN7DAAhoxsx+EPu9AUNqq
zGd179qYb6yuHtxLonz38N5AvBj8r1uUHQPAC1GNo8ewvuf/qE3DllbZWZcJ96ecN01pwOwUSNzA
tQc0J6RRz9snw9APSb/PJ6/4oLYEzGdK2GjS0Zz4Rk/MHwg4jXIVZ0opv4URMUbVHt0s5pedmFhZ
7cbN6Vgvx3CJ1Ur3Ao2FN/o4fs6Je4kNMO8F9d7PDGUH32ewK2O8ZuOfH6SBVRP6b/3CSbXcNkAJ
Vze+Ya0MVqqJwg9FXgtWMnizVcFGZsVN7A+NPepZk7tMQUQhj76OXz6mfsCGejG0frTvbjN3eRSS
UC1DoNXXz9Z/NIpgoOYbWEmaY78bzs+glm46cFD0pCMBcscPwiyC2Mk7uU66FTbK6ixn0zE+VzlJ
8rJJ2Qwx7EMkCQv5TSO6KxSckT2hTRGDK1TyTwvJO2Zcy8GAcO91WHDlBt5U0zZG+sT+8Vg+Q2z2
5uIvnPnWU+TD7jBCNN70k0m8luUtnyGQcIrMXvTXiNbmma10puFTHhoKzs1i1i5/A7HQrCiMMfvK
sXiXnxsemK7JxDyYY6bXLRlczR4DKXs9+8WewHqRoQJhVL1SIZiR7hwOx71bd9NksphyrwjNVJde
W+2TxaT9MHB5RSPMyBccpEMVlnSokqtemUBeo6UnTNHwkKrMK8rqp8ZWCy0iX4zQ0zNXAXFk38X3
js1y6/7thD/OlQwhwP4wBOMgk7af6qjfx+cczCqN9zUDqJOuc+oPCPWv/AmXSdAXW6MSLXyayssT
zbBLxnFyCx3P3ec5u6gb/PPYZCdNsoxGUa/4bibr9QN8KIXyN1OuMhS136HPBbmBncIuXTXksIKN
ynIE80g60YbKLnVmaOqrD/eVIjRAib4DPYwcOL2hubyxh2Sm/oT4oul4IaxwTMmekrz2NxaOVFRU
IG9uD+9nW8gKkUUXs5RMt4f3hAFRyCjkjRwZ3MAVHxzm2AgwBeR5F+iqsz0HxLWm6ph+d9D1cwrF
ihoLdH3Jwp6VuDEqnExqpzMSTs8u56TyNWUhkm8O5Kwh2L/9wngNoYwTnr+ThVfiQDzL2wJLWoxr
Z1WYAmzxNvA/FpW9e1uJSjr5DJ+gYygptxDG5HbPBv3eOUSZXQmc6q0k3evKF+CmI034lG+Ta8dQ
MEnOOi3iE7o0SpKSMwdue76rVqE0qtB8nL3yJo9wDt3Y8EdzKvK4uGkMjLigEstDydJ2eB4zmZL6
ZbZi3vSA4ouI+YWumcdnaiLrOvrWfmhs+P2/euEdwydxut7aEr65Mk1DPgMskiI1AjYvxMNJJrvo
GqcEqtGyPboVZUPoyI9KdJV/mMRYgmsstnzU5+yNjj60SocFE0gNzDonodVRJGV6GUN11vs2vEFo
NTzojSJ0+U/PdF3EmQAQOO4vRCvZ7fAqgt3K+lcQpwbQtfC/tjhIOv+rRLEcEfCS5RrN8q86eZZK
KDof63BlJ0H1IEePPNlVsIbay+BO13PRsmmD4sXeMm9yDOx0FvLerTog6Ck/UVHURRtpyeqrM89r
HLb50YKNViqii/CCmYorE6E0kazYtGJAD/07la64Gw/ZlK1K03YGxKqAfckPrdmspNHjLmyVqXAF
syb3V481n+GMisAySHi0TcxBoMMoEr9cDUZYqJE2PrQOpEDwZRIUD3Ris5c6VQuaU2NYSFu/4SV8
vuFxV8ILomB9Cjft/YhTZO1g/9jyVHIi4CU0HRuMluEtma8lzzwUwRJxKGPKZV1HL6hDBQhyzN+i
nPinGcYxlP98mf9uOOR2YkVSoTSrfoIe4afaK/jCSE9cqN67wcGUxwgVV92KGQWopgnCxbBWr01l
QQGuDoeaZSy/E6j/1XBPGU5uw7PAIP9YedSi6jr7Df59mSEvxFARWxJj2yOsWVExnnlQtU70MnlS
sWFUEHPZon9VGm7wa/7V4+tHaGkHCvaT8DlCsqbdYdKSoMawVDevOjtpIdvR3GPk9ptIl8UbiE9h
kHqIrr443AAt2XFmaPJ1kgWId6xGd2MZNzeJmieKhfKFkU6MF9cI4D+Se9p5kRNlXwmqAN8XLSm2
biHEv/yff5NC9PuyXD5YAeOVj5rwGAm+bLLvcLXps6tE9kWJmdQnSnN8KIn1zHtC7ckC/xMUofW8
UwVbx26MB4vei96wyCEdhwkAJiuXUyYFfyGs3WkcZ16xB3AxpFhxI844K9AASVsvPZvprvtKWned
RAG4P21LXCGwriXqIUgMzbNOTfz3E0D57UzdRPBH/cmdvIO0iFjDdm6UbZEja3D90I5cvxkCnude
y9gxF2i+dm7cv30XjiZQ3qP5Z2etEdtttMjh8WTPYkiPSU0KuwRPinn2bZBbMGQQVKaHTYM/k/7D
NhK3Nc2htKPPnxfrz+X5RYvmWxpkQ/i+lVZ8cswJ117AyFvI5b1c4ilx97iMEBfAUUbncYeV2aPO
gmMf+qnflm5tvBgf3YSNyYigXtd0vClbpRQmW18Z2IIInoRamCUsbPNtJdzPTx/p30Adp2s085kC
W58BqJUI0nxDboj4jAuDDSuoSuMfbvR1a4Cdl2A8/VW1qe0A7Ui3eFEmMC1TPmbLnAIbvfr9rjma
TQp3CukTk09UmDxpLAFIE2BKBYpvAAOSQQWxS8FmH46B7ZwCHY4EXqQ/IiyDdqUnzHwPnPz8KWYe
0cR8tPC4XZefIE4vKQBNdr6WufhFGpur5fG9QHbYcOvt+UImj9mg+4njEAvXc6bHl128tsch7Lba
SdMAsvhYlRUnY4AsjruIMlc0TLknR3KHYnpHOYHq8K0wNSDs1BT7W/lHyMQX7NYV5oLNefHlJsYt
Crx26C9DNInwtWQVKHPdl6QbEWkiGkr/fCUIO9T8BcwHtf8VORLUwOOA3n5jFut7/7INeBihIY7P
Mfzx/bD64NXJFumjvaTXRFHmDEXtmxj1+uuhVEjx5JIKRSld36fKFf1uKxDn0sbZz3D9LRvC7Y5V
ymmN9TrNOg/5bFo6bMOWe+8pgRvidKbxazoGvVJxjaFDoZjPHxnvKAlNazEQDY2TnhsADtAq+6Pu
iwcO9CQKOm/w7cRIOvfSxdIQD8bZCPqEGxO9MW+eCZgi8wDFdjQGHOwnD0Hsdl8+K7C/Wteg5z7x
O/YW+FGe4V8O5uAI/IgDyQUMY02mN48C/Ji0rBtZDGwLPOLYLGFKCgCIO53UQ26c1aZvulwOSWsH
mIxIqysXLk6Yoie0Ag3aLE2j9n2I8hixB6jgJqnwdt1W06m9hzSVvqjJjyU1RJl3CAYfXnEWtpSQ
N/QNveoGLgiEexWCXT4Kyp08D1zw1l1V5ryIwSefhCviaOb8cRH9vbLBN/S2Zla4W411PAzJDFnl
zMmcqWb0u72ANVGKORPD86DnoVwRFRP4MD5P4tIzq+OnfrsTP+AVV6VvDQ27ONjth8eVD7/WvbZs
A4GBoFmJJsCjYbpPQLaeM+iDiVDgUoRaw7arUyQSDcjszFJUYHpoW3FxStzUv0Ya/MLuxy4g3yHK
uEGSMrvD2+NnondKVoAMjDApAyxWEQR+ARG3ZGFg/tEQvqPJZqqLX21sbJfQh+tMtrEm50GbI9hU
uxifOmLFiKO3qS+0cCk7K2nmcurBPfuGHoic9KjuFiBhiAap5ivk9pliaBJwUkgRLauuanZBoQ3P
1fW5Cw5tzpvUuP+X52I5IDCUnMtQGHZ6LRiqag3IlwXYWSjGQpjtlvFUMN379qCOyzJtY4LG9ux2
N/mi3WysX2SsOn57BeA+rn1P5/VH7jK8caZP7wkeVxjEboi54MVO26mMvHCjkqLK1TO/mVhcu7om
c6EC99ol1bfSNH2n68iAko4cJG7XCoObJmC7+wiab081FtecLTTpdeqrktT4k3Q5ZjVlXxJpe3jV
qNDyvDJderNhKr2cXjWQV+qkAJWV5FBGev9Ef7hSiqRiIquEtc7gxgAjpGJQJZvY1C8Gj/tm+de4
YvLtUhiWL/BYakTuI/H1pZeAx5EjlnGetqTNVw9uNMuKzDhbI3tBVnTdANorzH9X2V9RhJ6tZWnh
tPBzrFclGfbxHRoa6BoQsFUYdZjc/AXtSBFaBWp4nX81MnIYp2uaTm0ZnDEZy86rrxKwJKtMl9iN
MSsKQ/D1uKxPnpqhaRezgANBVNatCwNOlMv0X7PZru+E5XT5+EvU7B1IJddcsWdBomey62hsQ4N8
4UnIAf2slToOI5V0c8Dnu9dvtCMZG0zyfZBRzLLS8Cv8yhWhNGHhis84I5iGJB/Cshqv0nyTCRSQ
pgNe7Z20BJui8t8k7iXG7lXw26dSqAgRG8ZQX0ZBjeaa2kykwwwOa4vpoFhPu4bCqpm6eA5v1jNF
N/Rar82+U0JpOlOUq2xBE++DqllPY3xjCDl+SP2k9dSHUUehrgt/iUr/Us7D4eGlgVin8m2WFawD
/n1U7AMTRqKTQw/numP08har/VSpp/dJx6J4cUV9NiYBGWsyzPwGUiTHA5TPlLrGjyAfsgSSfkyr
PhYQQbV4NXziG8avK9k63PjRi6/oGnE0Im3+u4EdjBmGUiB+y2+U26NHiCEaPuFRayXVeQDsfCNf
evK8P7TWp8bEM/5C7Z1WyRyxbzEEJbylaV5Ecr0CfNu3eRpFWxGZv3WDbF4fuvDuGc+hIzeUoBQf
/iCmNOKx6i5wh0klN0yOkjCmvQxU8eYM7xMOVIq0/u3rcRMs7W7+nhgtZAOXVzLKbP36izdwhMw7
hilWY5Hgk0kdRvmkgz2TuJJUoZlVr/8LoXWjadBs4faOqFaOqAj1RTAC9hsoE6r8al4nwljeyXFU
aVkmXCD+yjSVBug/eQ8rM7FGJS8IKb0OyjXP5SxxBvB6Oj4E95b4TjpQQPkbV7y/4igKKO8rg877
NmnYSfmkfh2N97ExFyEI8ayqJnpYUwJtFOkYOKcmGjs81GH6YWLMK6OhLwYUk7cmtz7LXiQEE6h/
Z54/pOI2riSGTA9AFUT0Y15YAOjn8S8DXpr44CK6Egz6C7MVlMMsZfsyxcX7agvDhcNdegvWQ7XW
PQeSLch5RcMQu3feNThzSbu87QGae45Gup1R23umzQZ6FzG7STCr2q2HwmZLpm9hPibrW0HvK9Ha
0Ip4YnNXo8AQQbqL4+WrlLH2glR7j4PaC5eXzOgRZabDN/PaT7xtu6H9tHIdSOZQ7pO7+J91LENi
9dgQ4jWj6gJdyRdJk1BrvRXTy2HHVnOBtzaSLIftCduyVoey3GoCexYdbHcBoKYFsQvM1Ktp5Dcx
cX5x6aI9ssZLrydTS5xxV14wZpNchkpTipH4vdherzs1KwFcYprjpBCmKlbW2XEmrAByJXvlRBje
ThO4Ggc+zo2oISM3bJ03bPRLhC5MX0iVVFuu39B03+76ZiY7x5FhYMScBhKbXOu9ZbK12dMzg3L+
0kXIdnn6nxVjGvfM0h+OaRdr8InxDE/G8EEgUYiAzu0SzVa/gs5Wy9D9aW265hLCWAjk9Na/V/1a
IgTP7NhnipUVjbJfPNbVAME4iv5CHBQ1IJR46lnspTB/JpCHlFWxZ/aXaTVbpvgikYoPuniAU3Rl
cYi07vrhvBSPzaCM6hWNichDX8H/YTJJGqoA6fWYmpfD8ei25JcQaej6QW8gCfonaEmAuab3fq0J
uaoj3nGsq7BaasV4IltvLx79hZXSvjlfUhq42a9O6DxhE5uKkKA/vVsNt80YulkXeiOS1kC1AYfp
lB8StgEz7aRSclKm7vQ4kFVvJ+/ip5eEyPDy0Z63GfYNtHc9Kqly+SdQxqyonkTGLRWklHvRnzOS
2JZaGydH8MJRyO5hLZ4oAxlDr+Tqt0lhIfXC/ZAd3rg8YIzqma2aKsBc0kwv1LGefyBWXuEl7D3R
jlAeg0yA3HwLsdQcFNWyIRplGXBnKTtBXwAecnZybYwWtp7PchoK2NF3FC1txREOSvabVjDzXKf9
SS5LZyPCqp5MVVYialT9lQ5Hl2bKN3x7c0atSV31QgLTy+AtwGcVglpuoWgJApXvU/DPKOZnZRTp
QjGtniXXnmeD7lb7mCRuKc7gqWGH2uTA2GOXfWCHyELa0qfLlK9L/FGmENhqCjy88yhv6q0UDaKJ
tFek1b81HRPnWw/Xm+MpZKLKb2JKmL9epqhCIHF6LKHPe7TM4PFt5g0LWrG7zX9aneqDCl04y7Ew
ec7e4bLMVvY4UdXVs2e+Wn7niYkuGjeBvnkfB2Hl2uv+gU3vwSA3tM5AjqJRVi20dFfsPpbUJm4E
/IIdBsBM4/4OHRtRFqv54ykR1KCsm64D9z43DEk/iOAqRzz/OIEJhHEoEX9/f18BDaOVxr+XH6iu
5gyGj2qzgrUjPWxlgUUpSFkE6dyIq+6eEnqiqGidCdSrYk1w7VxqPaCihnruDCqwidIv0+GqWHN1
ZhSZC1HUJSelpQWenSvZEbyJHbfw98CMILacBvuKLLR5IpRm+t3spRLrc987jC96wFjlV5KSReuR
0qC3FXQgOZzoNQVAiGXnp+cdsrb6YZmEuUUTX0f9015tOUmQMDz6htYSL55vdUMzT2nWWn+qiRz5
WzJ03US/KInMCgdzdMWYUZXJipMN3OD4G6F7M3GFAzO1ILvzGIySPTvCTHB75+AXR3qwYBFcruWX
mxGEYq+cHdg5VmxYtKafMbCxpp+3n4jEKlC3Vd6Z8Ia3qzO2eL0XZupKj7poClUCSPCAPv/6i8gw
t694R0TSQV51uIr44rC+58lPoJE7CTPSSQrC5gzEDgYsMWXBOJZArhl49OjI4L9/j+9z5suRsPpz
2ITKbexE6qbUEaID4Z69X7AaLzWGC8SrNrRjdWlRkD40ho4xhr+J3Pygq3wRFVTi+PcLtShDhzLS
cVvjVX0HuVSvLx+TIvM+m4IGFFOXtk5ESQ4XIrIqYHZezotMc2GdDoKiVhPKaiEfVSIcbv2lDYC2
/M+9ge6TKm8y0WE03xZnvYvQNk5DmTcBkUP8U3fTsP3jOjZkElSY2ny4YlN4XU9JiAfjruahUlU7
HUEn1kfbfToeQS+aPQRyxViyo6Az+EDmLUxA7LEeIO1osE5MFkWbCrXqy8bpMgZ7B0UPFSJdirGj
bkRtAxOpIdR081LvB0umQdAXnA0q64CeV4cYK+61JHygPdA7nbQpQ9V24YP55hXvEimCzZwE0LJY
VGS9dn2j5cGVF/2mIKgyCUXUMy/97qsCw7KJ48tbMLLczAdWIe36G3GlDph3xGzs1/RKef8Gblpf
aQIKWtrJRyaHzIpyVfYP8wecf8dmxesTn6iwADPs/ES9ALByhMqStnVvoobr4loLZSJ32DRdzLit
on+ditmhobsqsNzHoCqE2Vd8kUfL+qzfjn+PBZxT3aYCVNOYLcxN3cfmlE22I8FZppLv89AHPCma
d6CueqzwRK0F7LOUkcDoj8LleGM17zYiiH3HTmJLtTjnN2WWVWul7kw+ozjPa+/KAQc3VcEZVU/6
i7FST/9HmatT01GeYHPRa6PP61YXsnyLCSs70Ekf+BRIEfeDB4L5jTU0aGVk8O7548jeGrCO0CQs
TudGnkw5+SByOMAfE7q74+XHXgId3Msno7VKBglwWBc8LJIpw1zEJ5uUSSLTCo7XE64BtkR5zl8C
LeMO+zsP2/PyOnNM22dw6tmLAvMarTOXfW7tmSy+acaM5yLA5RwFTpkTB03IL2hRQje2NTUzTf/+
KuA0dcWudBLCpNi2GoHEUOm5/3gLtI4qyr0d6ScOtUklcv0S3Vq79VALF2/su/9SLE76qYdLU6nm
8pmZw6STdTUY/7m24TV9c2cDiPFl+/sWnCeSS8gqZIM4xlq3G8vGj29313gznLt9j+0a9+yNvqFE
J5JTFm+d5wHpsCnKdkG2YtwWJaYtVfR9CcsghifI4mtMdAN0zvD+1zCdHqlbUCLFwV1G6ekVsIwP
+hSJdSR9CB6b2KHQ4Od8y8yHIqaYkAUXu9zuS2y7cc8SlMfuDLovytF84qc87tfbu4ApOb4klgGn
A/Atyi45gBoaDzocleAUy4u4TG0wXKOQpYG8slGMn1R+rQrlt6t3gjKezSunOedXhTaoMJ+ikBf7
UaOk3SGcYhMlbu1XsKH+RfKpCr5OYcwTGx8XARCsCANafR05nDCRIDelp5walmCsrOBw4UggkA1Q
lfjcCfa8AWgupGuVhCynGSVuQQip/ZcYSd05Z3dYvTHB+ebSl3tF+nZWS8zP4rF4dMxS7NCYd8OI
aq12HI5Ct5vybsxztgB55CzRGTpFzK+er5uNlVI3e3drZWdEGe4fXZ0bAK0is8qRYBwVZF6jQ7Yu
yquB2vIaA3svn5kdEeZXY5tYn0dMnRyc+foput2WuTMawmoHUmBo+AZzrLOhSSc0qm6IyzM8Dt7U
Zz3ImFaCVkr2aXg/smYCFz/ARcfMgtX7z0nwMKf/ZFybL5GTcQSJo/g3whavWqRp23YPRFmw/6xh
/TzENHcl+onFg2vUSvK6lfcqjtCo5BFuhxYbVyd9hjDHE/xmq6k0TOnLJOHLioq9Y+QRWoEQXI9B
JLkFlD3PapsEXiCz2UOTUMK3u0IUfShlm308VvGnzZzsJIv4UPJsmTAYUwYQi4//iWeEXuJ5WCCN
wYpbs5BZXFrJssf7oxqiX08a0gooKgABjwS6osbiZyTU1BpAZ+2WijTbsB1cmoubyRqToipWlW/l
7NXoxHsCKcEYdE3cIJycyKIOMCsyaZ1SDP9H259yI6yHkCEEt75SNXjUy5n9PyYMwkNW4HEz3T/a
X+tJxITcfUhLcjgCx2SYq4qRZyvi/+UDnvyx6mAYq5EEEet5LSVaRZ78hIP/QSWl3QQEizBIQham
3R8K7W7IS2p7r1nF7Z9P7QLxwIg2axiRAuIs0jIBwp03RzS1NWDkLkuyD3kTs3oCmtuqNUazyYA/
y6b9eAxtD6Jq0z04uMEczqeF3jw8CgOAhi0F8eMy6EQfdpZZdURQZKoskhGLkGVm/74QgPx6BUJl
San9V83bfAaMbiShhREF0B5KivpQ6hKAbtTv8fcNASqzMilFw3rC5i2v00CsfydQTfq6dBEMjuz2
a3xt/wvdemcGlthvg/iHBsuwV2PLrCCmMpA7LX0p2sl4BVDHmc3scYGvwi+6/sEuKWAH7bdlH3Uw
rK8dMirOBLu1Juj+dpEy8Y55hTYg9Zvyl3IY4TTRzQWN0jXg1I4WPyMqdxv9W7qht9R/zbQHRO8a
ZpAAq2yCLp6/YyXwvs+6U87paEse7gIqSJqUlcsyAAB6DxjedYRG0NtjaUXolTRk1ZFeQQZpfPPX
WiJmDdDvyQZJgCINSaUSwOvoNRRML+b9x7ehcji5h82Q0d1TFU0+eWpqBibEmi6rJm/eCODG5E8Z
+8cFcL0IoLQG8Ee3qVGHWP5iCIa0tcOqqSEANlYpqlNV8UdPti0/PvxLxE8613vgnp4HUYtFoDdL
qInpL/O7VDQu3yiZlF60xCaUNWfYSP42ggPI7Hse6tbjEiu8McBblQa6BC+FFDsEZFzY7YHecdD4
L6RsAmkZA3YyhgmPozyQ3yz4Dg1goTSeTFOl7byeh6WYNhQ3N4Tse2HY620CcbPPQgdSA7mEYGSj
86QWSR+Z9repEkiWkHTUn5A2PN7zsDBG8UYTlfaDmSxFOibWK0avqhNo2xGKmMj0YJK2wEAME1OV
diEzupA7Xro4Mk6gGEHJrY135r4fUzMyA6pg4tRSqZba00WhBa6RdZB4nmccQM0NON65Hbzo6Fup
GShmbyJayrUl7t1qzLH3EXWZJP8mugY7+dUlmYzfE9+HYfrmZU4aIb2ogD8ynFtLrgN4AgGksHsX
lKze5NsQ6dh+1oSAPZ4+8jAwDd5SYiaBByYeWl5G2XxHW39kpo/U++C2dkIndJq3fakwrGE3FlWl
tKnmNAEkKYzV6dGdDr4JwQ+2Xv3hVLW+686h0aqesyFkdWl42roBXsVPr2IgqjMVpe2rm6EktqJ2
8iF0ui/lUUq+s+A0Sp6twQ7QmXhMtwwWikkSXPGCPeBG9o6CXciRxs1lxSrZDd05XfbwjyjhxdjT
YC+U7IXK/hjxPPtJ1z+2Vs6Y9V/NU6BuElMPO8S6ZKhlB2KkVNtn4cLg+bsbUO5d7Cj5tITKyYG5
ABZ4f/C7qgakD2wgS2J9TLrpBuKmSRbwJmSk7v2XZZEKR7tfo1yC9VP9MXix8ftYtsus5lQAQShR
wNptZCpeKlC8Fz39njMj4h0xlk7eEqkif1aDWgHBjiSILfmL/n4bI0ZoPEJi0WLTHZEujYXs9+ss
PTQ1ym2iQ6arsy1D1mbOM98xl5so8qXC98+Li4ZOlayycuULfeCCv5fy0ekTRwozqmaBBVQoxnh0
f/HTxti9WEk7FdY69zRX9OUY0giXFBQDWScJ/4gdMXeqpG6cJ2CmN6qBJrHBDBj5VrfIjkxtxRVS
nTJKSGIwXnUOaXvJmPttt6xyrAo4EBHqqqFE57d9fF8UqQbCmI+fYeW8bGEJeW/j7Zb3xJDLMeEv
JRZ09Q7rIkIruMVXYNoHZYVmGbVGwIdtqY17BY0VWjIQDw/sUs9p0cBjBM24L0WCbTe6kCJBPoB5
cGy/OnqQtyNXJ+not3JIav/bjSpyPcd6dcpE3ljDJple87w+kcEIz3PEILcSQmwUOrhXQeeSK1Z1
2GqhdlfTu+bjxDwofcE6gBF1ikGlhPMoffsK5DMWT058aSdBiM8Q/NxaboNtppBDgTQMxwTu0HsV
DdNN7WxVYj5nU4sOGfXeuld56KuC4Eo2NcJnT4FjDoFFXfs64DhOxLsqMnLk7YXSvKXR7ZYmzvE0
z7no/ENhK16msHg/chZdjxxOb6rxqIQknEVhCeWytvnyxbCSgPeNiEpn0LwA6w5+lEWZ1bLuiPwD
JwadbMn8VDh8r//78raA5Ll2HH429l1nlWFLdTMAjAaVr3BbIORILo6bwVywyeQoLBYfXgVfZuXn
J2WoWhytSFNC9zZGvr2ZAlaHMlI52NJ13xdJzvCbJCw9PPtGS/Ssn4cd5rs1QZ5pplJLBrpLUEiJ
Q/QZVP4oDKxHbxfpzll43IVOlJCyZdkg4J+lefuuPgxpyKTtUweioyEcLC9nQGCADMxjiZFNa5L6
jF9jmZwGyCA6rMI8IkyRRxXpaeYhWY5epLYEJFK5VbYV2uu/31new4TEme2wTCtvDkt8O8HGbUKJ
lJdTOhBt2lVBVZ9RYMirsmmjzP/zV7eTRi410pkoKTSZKaHGf0a5H4IVe+zj9qisOhiRxfWwd2AD
JHvCiwLL10e8EbVADRRmDMz1xthY/eZMBPpWQDBx+8AZCcRu+ZEEG6ofp2/miHov/SU6Q3cyZEdq
CUQedvPKY3tW4E9Mu9HR2HOm1VQwmi+YwN/WDvAC3WKAdQgoauocq3jnniyEpne24hQI+sA9dYAX
SEJ3MMRwn0B5gk1nwgQYNpnJAL8atmpMkTzLUZxhod5SeCZ3RBeI4tUhi4ps6KuJ5krxe7pw0rG1
Oyy72MFKUvr9JkV+MOwn8o7r5/dHn8W0dj/h4TfZ+kWP6AlCvaB7rVRbaihG31VKmCc3iJu4wacm
SLc0uDEOs3J1XkTz8YvtKa5fz/ftAKQyE/szUYu/uOIHveN7puPVOgrGcq7S7sq9FRDkgPY8eK3J
Jl79jU8ULu4gPa7sQRWD3VtIgggixb9PJZvi8Cv1P4WBdC23v5198QO/O7FaDlqSi8CTN+5nAVAN
CNtEssCcULymke9sOBIzaJb1u5GRUXREM9rtoloytsxUWb+6iLZB5hoHNx/5uLEIWBTUrnvTYGew
K9oaRmWQgi05Ea8eUsYZp4BXggQB90C3rJo5hSUiHDq/HJR+zhXfwV4ichQKBXJPUtyYPueO2s2g
5MpRZbBpO5Hm8Zhk7nk3aTri8Dizk9r2h9xT6AYhbBhOMj2rUctaWA3jtNKN8vaC5Sp596f/WKKG
+5xXICG84GG2wUhktjglxwIMSUkIE8AZen5hCk9xEY9iqIV8e3HO3cgilSRw4nt0wd4gF+eMGMGM
LaUvsiygUw/1B8p89odnKOuwY+bhHvSyBG2KES68Wpup4HoyOjpWncgLko9oeBW1QEuGearhgXFf
bR6JMdZV2hn4sw8YwKptkSuLM7vu09efg4FGqdD+1SNtfpFNriUFDz8ezEnsg1FD3zK0XTx4YwBI
AeJFMoA6mXP8GDYILf19s5UFurGUHHgakzzaTfN/6qvVLry5cB9nwX2hUCZA5dDesJNhvXOE3SBL
8kmofsFVvqY8PMfAEYc6M/ohkzN4K+nwYjvR9k6ExqivAyZDsutkadoYx0c3T7jaED5DqUJnKVLT
tX4/5MLGuBaEGPWA1hrmQ/FPkBDLpGelMW9HXYa6vUdx5UOf/Rdm/AQcQ5kX/Z1xz/M/Mmz+f2S6
355CFr9QibJ2ixBFr8xP9r8khUSNS+oOD0M5rifWX+5zl+9byQAdn2XH5RWW/UINx4ZfuJWp9AKQ
epa1vUp6K2ejxwafvmXK7C4InjNrc3NA5JZVMz2DxlryND5IKCyr90FU9Iy35joq0YD2jbE+LYuM
lIB8ULf7u92okxAjkrEtX6ZWU75G8oxnp7pR5M/yhM264ybVrgqSbS0sojDtL9unv+9p9V4T/wOR
ZiN6Tnfk7Bd7sDx07Q2ssefnCABhE4/eFDityDV62E9mOFV37eMRj232CoP0TCaiyb7+tW7tTpFV
RmjZRY94kBordxJtptilCaxXQAZDmbCqAeo8I3VgffUfxPM4Bl/a9JtC5EXXx/YEbf7RXU42NGrz
OwKHJmiAB6uCccnDu8lFoU4CbR4FlUT+hhCGRZmOj12zu+5Hj5Pa4jC6jq6yHECrH6jF4teXyaGQ
+ITHvxAt+t7G26uu8cjRtzXHMIAe0oc68xQJoEoVYL8mKSGB6rrWvS0xyeCQymxkPP3A08mPWCL/
vnOwK9+0m+o9uNGIVqgXEgZO2Xve1CNbiJx/r4Ika5/L9ASihoS0MJpf35gzSDS/l598a74moL1M
YTi8bsG8pGS5LqfJab1oZi1btPSwhGVjXXZ2z4+DoaDEPcOdvJaJK5lVcXzjSFfzGLQ4KYbJFMeJ
zkyWSCgs+eNApKQVRub6hMPaEB2LcFxrpnG+uDxHVVYEcS7e4BtEySDjZN3MoZ2B9PDfyNmNhosT
RD5mXooAWSjOnxmFvP6K9n6ngCZigf1F1hwbO3tP5InpP2aR3aJVtkh/oUBlOy3PYFKx33dUVl3+
lhnuaMVoHQvaG///4CZgInBtJoTWzotBgiXC6QN6l/psErLSXwaS55zdSCWgy5bqTwDlZzk4sw8h
JGTd1yfFjCrBP5HnpH9vho9QizC5aI+R0LcImN/kVxmLhBROwPVyg4glgEuoA7vroNCEaOMFQRW4
dT0rHVS/qOrnTghse6HHtHAmJF9uwOAggb++mLbAQf07xh4oyHW9tHpxeSv5FX9kIs1dc6RhDS3Z
P8E5IDZMc6hKUpjJt4teCHtX4unGwN+GkqjIciEZMg71eKTCn+pXPzh5ldl2T5+hJxiTZ0qBWQIk
8l64URi2mkwsGfF688+OIelrnGPvliolcU8elTcawO3AmTzQCJfxR3rJGp2QibnJVxltoOf76srv
G6ABlLE64B9KsYNuLmj81YPPgIZmiLzRZbmOiO/f6RQoLKQLF1IPYtXLOaoEgv86qgsS9C6Q2WEK
1sZVMajAh/x+690hwEulOL/Pa8Bne0yBeiSaNu5tgJCW2ewW+tI/DB5tu8zzO5Fj4uzPa9L904mp
+B8qqsVFWishqesHDgrRLdkyhWP9BgrmfiAjTwQABjdwP/4P/sku8X8B0vKM/XO99PmsD/DXKs8F
V4Ux7bHWoWw190geFBM2Fep3fnP7gqWXk2sg4mVSmDRs3MTHNtPDnVKIYK40uoaikyq4huo/g8KR
9vM/3LjXSBc4PIvORBsN/JwTc5FBHOIyJbFlH0LOfgiosRFFzNlswPTlLFp54b7nkgHiqMNaBGgR
/yVERsUwf3hinwW3EXKcfxQl3XjgWTHob/oTVtr54r/KSn0qzycWQTgpsASmbwZ0uBtmV5FPZLF9
s/0ByVP3SkareiCmW9XkyFuzMw4Kw9e6VLu44PISusjeD0WNiPT6iu9WXu7dPoJ7xBakVna9roLt
KDmByqDxHnPbIeGUcUik371+fuz/kRzDONPkwF1wXcwa6qzMA1KLqgiZnu1GTZtgUVgoXDyaFJGO
gdEgDZNjjzL8bTNKB+xm8jn1eCnulp6DDt3ZksEn1l2LnHtqMa735MCeLCwm40heSILV/kMfL1HC
sT+afw0tlBqnY3VyvmdAc6c35ODV+nHl0CPyRkvoaq2MRFWNB7/AFOz5eiY0rS8I7rd+7QHsOh7Y
FEbqBn3B6teSudVuOUqT6JM/ZUey1WYRV8jTaXvz7C/UGJzJJcncbfwyvMK9KKXI9671UB8CAZV5
vn/Dr1lKVqfe/lICK8cxbcszvWGUBKpT/tkxCIh6eSwrpOVqsJNvTdS79Ltc9q06wpVNBiHHtAKV
zBADY4IT/CfzyEUstrGZAs+8efz4W2bvD9yqfKmc3lSrxI4RyKzph5Ik34Dfg8wuKmk18ugjvq6a
Z6PtG7PnqqppTEtnqcAuCImJRf09d5kh5uM5bXvUk09Y0La8jc0R/VIwjVryrl3KF3xTNDja5FkM
zHYHE+4ufHzCZS06RAmM38UiJ5nbBE+2e/tG0BsS3IPBI4Pon3yN7Ehqb9c4LUwWKfbgas1Y1xsB
/Z57oce/xtTy8BsgAo0Y+mv/4KvK63eOi9qow4SBDId4wPVOi71rJGKonl/APUBDRg3Vwig6n4rM
CIz5E2OPtUvDXdHdHIPXYRDBc2nIrGUVYhMdJMYF9OOT015+z0DsMa16toHu5IsSqza9XCFcY1GD
oCAIXDcJv86vM0wfWFxP2dcIBoYUYYhyASEzW2UzMrebNN5TFh1jGT16EU9xA2MSxyvEvl53b6XM
8WpeJl/onwuaZiTKGvUnw15hqLYsVv+eKTHU9YJv+0B0gq3iH85nCHP2wAATExMjp02QYUWrwcL0
5LvB5L6MGUNkV0di/FBAH98Q1AOuPHS1XzuAP3y4+7nSuVMoTwUl31bbTX2JnoOKcXUHHcv7SLmK
enc65r/ureI6JaIKSYDyTUV6AQD/PLeG6bN1+WP34aNd8u6I0R7VZDx99/aHjuEDsxqOobFt0btY
RAeMM7ngBga3401tXe2HA3JkKXBsE/SZL8YPc5O0+N+W8igPW4bmF++88kP5hLtxMVMHIW9lgl+X
GRjMdjdeDbhNiyJlVb9C0KP/aLlPYxhQ0SscEn/A3/qyothp7huMUrN1yiWLyI5Y22TQ4WzntMpM
//po8rxsKSZBtdb2KRxd6H9k/JyN7thgAkqfi9p+sKJxS7OxHRYWjfkMNjS6G4i7/RfTPDU8YFC6
U4xbdlsa8eLGb3AAtfc1fpPFu9eErPDkeaQJpemortf6TMyZ9hsl6V8nBgs/4VCBhNLpwonuYVja
GH9v828JqrcJhiJOL5D2t+WgBdXDvLEi/bRqWsb5RWd3dVTJLYu8X6IUyM1Sfw3v+jaeG5Ka3Heb
ToDPf2+4M0U64WJsFlG4tlKaVH84WQOWOU+jJFRhNOf/pAuoBnduBq9QX67bCCCc4ttFWot232OD
/swfwcOUb6oIxFWyLNozYarDpbSoRWMUhLiDfxVwBeGxYc+fFTp2D2gc3gqE1wRdMuH2sb1COCfR
zrtu/r4PO8oTCXJD1qVd1AfB1pwn4fD1Dar2lI0IaMEKmS7DuBvslxYlboX3XwNIRoP6dyl6tAFk
SDmVw9Ok8ApgcW3uEofc8qtP7M+VZ9ccMWyhanpT7k+UrHN+GQuBf6p+wy1gydye7zMk5aXmisWw
yxCn/KklLUA0jNrdeq1aaXmprzJ9xp40xAVEgrs2x8rCz6ipWAj/sr9XGpZri3R0lWiaOqsufXp0
kEtOXXw+halz/ymzH/9AxfZUggdjQlEDtZZ51P8YI2FpOxq1+lI9QlFd/90PAkokXlu+KPBtev/Z
Io8xyJW1nA7AS6i2yZxOi0UAXipcCKXa9US+6BYJnDmlQZh8+tDcCYjBtsehtPs02z+vzamX/Jrn
HXRNZk7QlrWVsKGbIa1bNVPMKHxJH6AWmUsHkSh6h5M4EdOsGzclCNoJL+VDEr79xHytEnZ5fOvA
no7fDULvTvQMRbYIICP5Zman1x6H/tyxxR+A5DuF77y8tWkJJyo4OBegOK2opYIIo+VVDEf3Z+YU
VhqeBMV7wdyRDTh4NhlEPEjcT7kMHhEv3TkKUTlk10T+BuBXJ5UhG0gQVVmUCE++9IrsE9ZVU80T
yrMv3rqzNVmfOX4A6GIElhrJEGpbXJ+1IQrHjUxyfuKKUrSv0RSKiQHmk9jzmqfAs3OUvS0T8fTj
8f3lUMRc1IDNbBEC7ZOGS34ewd/hhqVb9uTMKI/zLUaVqYLwjqvzbDu2svGlSEqPxIVce2BdY8VR
EQ/qcPdxKK5IExhHIb/RLAvh7SySeY5/2izn4xMlZCipJL9b5mKbJnOOSDpk3VHaWRNGDKgdJgjw
TEBwyPfmO41fwXpRpkPArIMzN3oUgiFLvk8727dmtPZXdks75Kmd7gWaNiGB79l2jMKWUD/Fn7B7
KSsBE9rhfnNW6y8FIGYtGpJ7MRH+B9gsa8aPs0JHnU7URobrWpCYz/nXfiucJL8w5txH3O3PH2E+
Rk5jSB9QlJbCF2EVOiT/JQv3kEgBZ3Epx5BKbdsm1zubyLr2KXrtUWZrV1JfBlTrEcd9Q1TWcSsr
3Eeid4vIi5gSu3w2IRHVZZr3Pczrh9SxDI+A+qcOkSiIGKa8zmTW5CRPU1A++shhkMvVJeyOcysm
LopdEi6V+TUMOlN1WxvBaNCA7/Q4hMa1n2gyHPPoQ1zNRTDLON4SEEZoZrN8jGSAUQehTqJyCl9w
hJ0REJAh0o87DuW9Ly870B4yThUVlLUVTE/XOy8F5Cbei1y4lJel3lY/fhz34oKUyjshTYqKR4+E
b/0NT6nY7v7ibbDFQVdoPz2JSSOwwrFn042I9kRNskMsrgwUqWadVLT3KEPCEMZeSuLd3f8RTcw2
o4HacP7JIJFoIsZJFABw22brRB5aqYurb3eWDKCLrqb9yeupJ1MRiHwE+ZCW9EZ2xMmk93mbEha4
pLT5Pi/kYHoxSTbshiC0NaAPdAVbWHv+h5fvxwmlN/3LmzVL/JfYhXnyDzlRe9Dqt6pksqfxonV7
R6hu8ObPOEc22bv4ZYRxNLSnFlWZscrcDZpg0sOVPwcA8HawT13LZ0irCpRkHg4cNTZAkv6IAruu
J2PlxB0eQ/tXwk4xf3VcqbZBDqdtLS04SP3HhpOvvLcO4Bkb+U7p8vMxlLjXI1OyRaIwOtkcfuku
aEoDt2SF9MENh7R8mhZllm64V7/njnWlhLAPW0Wpp8k+8Oi8AiTVjDWT6YGCHIkDpuUMQEwJ7QOG
YhQI2L+y8rhtXcdDBDza0C64gZdPfGRjrJp9Xns/WP8Pfv6RHpw62O6LSUx4TNkTovbfb1KQ4Kq2
QwmKk3ZgqklcPabmrzSjujQjhH0USMA99dqkispN3AgrWbfxvV5bS7ZcCq/xTgiwxf4QcamF2rdq
0EX2zzCPnAHF/DE8yCeQLYccewNsCwszMcB4TW/77tudipWz4gbBKY4GIYlpjcTLhfjfXTO/Hwjp
8q65GJmXhN+6VvQUsJGjPlWO3uqtQJDmgxzwZMRlfEHt/b4tmXTz66MJ6CmCCVcNyf3nd8Ha4/ZS
xVLYeIqyNytC1OllVuY77U9clf8gayVC37VzFVOb8LdCZMiTbMScQj19wykX4HGx3EA8h7uhexsl
oizbyHjUxi6DUjjsKexjz++NJ8kZecDS6u1M7CJ9+RyknkY5gUVZtmEcY3rmXo9FHN4RMRZOIJCW
jdrrPbBlOnG3bb1M23UtGt5LeyDH2e3iTrYmuArqoLEsk0UcooIJby6bR2s3DuR5o/H3TSeogzSc
8sho8NjVwHwvcSrwO71/PFeLUoFVVsivN2VBlJ6l5YReVL8lYQL0/LuWD++5mYB+6bNsOpBVWT1R
z6eOzKPf57m2rTiI27XHMRUkGv+2TXoMf3i8dSJ5hM/IsKHCgVBwxoqdQ/RwGNpv39u5K+bEnGT6
hj3Jma/rEOzB8Q9MrDA+eB4IYmHDwa+h72j7VuWl+lVSR9c4O5RBBzIUZXThorc7R6DFXyvbsayY
IuONLotPLlEcWAe16dIiT10LoxmsiBfW9fPXtBwRrDqgLst+p8FSHPVaH0y+yIFBAz8Jk8EpBNkf
2BqBPVSuEnKaNatoP6Y3gg/z1tnHPMNapjDdYk6jc9IPcLDrXAGW7hfl+b7PjPBRRze0zpOw6xhP
u87N3J2zNd/o9uh8m2UgyRia+gZ7JzlbSYgiJ+vtibwVTo4Bf/VT+48dkBsbHFvWBRDNbCtvNNhP
mjewjG6Oc6hyu8lTU2QoN9VKQvWnop7QmgGYCkf46V5l9Q2W3GAKbN4XeVRzVA85slq8+rYFvoF2
McYhQr0XUWy4efhKIs6t7V4TYXebTBblRmLTrcLr3VoSMNpzEiOjGB92N8q04hMAo8AnRyagfwxL
/X8mmyOrzrA/1cMbMOo9Q6gk5D/Eev6PmiNlLP0mZXrsgm8riRRvZXRLnvBcltl/EFzX5hnvc9he
bYv9uxYg142Mav1QmV5tEF7QcZRLLuDvG5bPQF21c9SzA5b9/irv7na6nWhYGlxQugUvns38MZ46
0mib1Ao+zP/dTyUJlpxqvF51T5qOM6PrnDBrJmOIUAlkcJmVWKl6Eca5vqCouxEyuhtBOdLnNd3l
6OfHBjwQIwje2/CbkwODBvYFs6gGGvq3uMtC9kTbCEjaxczihqf1G+Ohj0qnLvUm44bAbRQrIf0n
udt7eSGIYvixaoGkNwQLgxWLRV4OGks3HCZxMRbZk/pFQOj4DpCUQS62RDYVc4CqNmnCoWevqV/2
vElDyjaSk30734OxjiTJ5f3Uq/V9OG7inzeFVKSzk+EOZigZK6YyE7QESAcfDKbe6eym1UoGL3dQ
3fYqVoGwWcQx7Q44SFS4bcGoUlVbWvjFKTOsgu2m4OAwG0ehnSnHIJtXRg3QYUNika+Xz6VkMNMk
tMP7cdkV6M1CQfGX+yQtRVHbfonGnFuigwHZVcSvspq4dOXc3jCN7zz0UnfOykiiwk6geAbswFm6
2H/cB/Ca/Scs6pW8J+HKft3Xv1bMLb4VQLxBBCTL9BomtHEX/iTkvrqb/xYrvnkrr6LaxqzmnB2y
gGw7S2o1PQbKpOgImSORfThzBfZJMYPIJjpmuYvhJQnvrUbZo3DMbOshW7mEc5hYBsHUI88f/Qks
W3kKvwZzpaqDC4v+UB9sOdbQddk4KRvz/C8e29YfBm3kzkPSR7haxh1EiyppF3kkrnxotYIHJ0iX
QqOSzGf6q7GpRWBrHMjWErqULekg/2wCtL4bMQXFaFsLParjeMltpb/98nxV3+TmUjADRAcoC9MN
R9ZZNTHUxKsGHv7v/KjKncuAbsrtF2WRR9/oeLtz207DK3tsnm6EhRDvIZVhEiUFHDdT4QdMbt4O
tVqM6/s27Fxbab7C8HjJ6m8f3tvkzMKvz23KeY85GwT/xA8YsGvmEtJDUOgRKI4Q3oemmuAD71oe
yeHDtT+tXYxOlITGjomw52/Ms/VCYBlRzxYn9fbH45zq5zAkpJir46h4tCrl4eYlABJFPv8xDFLN
F76Tydne7P0wkI80dQIHD5k0QOMOfG8gXx4JVRo/zffYK5YsDNJ3ARld8vwBZfrBvNMklbMwOo0y
tq6o2u/UqbKOosirP68rMLZat35u6OgywxemJ1BeB04AX1XovGCretAaqRn5K+MuKNx0Z1j+x8mN
jTDxamgGpYZmNOlk8Q2pY2ILEDJlmhIu+O+uiksnLKuXX1b+bgkrbFbQHa9T0K2n2OMl+KG0Bf5Q
5K7jFoOGXGY4yuWQ7lzxHVkZkreh/R8D6qbeVpznr9Uh877T6eLnZBccdlfEUGnqY8u72gPcPhmY
VqXSnaWDsGIGSxPEgrwWw3b6k0jrYyciKgVqURys+Tx6lFqinvDYa4sk8zQsQqKZrey3T/HN3Eie
PiuBsVyaHb+ISbmHSrVIF0qIQkOFlA+GE9PyB1qS7ustev1VxkKmPnf1XguyY4nmbT2qVC53MQKR
ESOhQGlEFq96OR7C0xat0X/RB/YxL4T1UTOjZVmjR4mxWOllIlxxfWq+7LiK911piph4JLPVx/En
p3jlz7hZyHdLKj3Tuzg+3bdfwuprvH4f+FlamMuKk9WtrRiWb4DoCc1+Ffnibo5tKuviw92hlssv
jeq+lIgrntwX4cNMXCpo3EBFtwQtkP7DoOWa8Pw2HiQ9jEjLtn00OsbciDwqtdlRFmf3tVvXdlkE
U3X/gww+eJHjUfRMmJ/+k6EHiwCdDbrYQlL3OeMRy/a4eRU7uf4cue7VqWwEy9Q1hoyGZ4t8k0CB
Y+l36pJ01DDU1DfAUw1vR5ks+rB7JXbZ7y6oZOmXdrDFZxwORHFi9st9acWV0H4nA6S7pHJQ9VPX
Fie1c7qwV7dwajVwspoA3Ko5o5vjbqXN9LDm4tx5l10M2FO3vmhATsX7eUkXuHe0QsxhPBll3y03
Zlk1UL0QtoplwgSTKf11zOrtbAqcp1Ay5xyYUqXKygqte/Y0jW7n+QviOPHypSfZ5ZT7onIkd4b7
5y87/c7iY2BFT85Di2P4Fn+dMhmY2eNHua4RoDrbeooQW40qxA8La7ypz65tXsh94We+90OLjgB2
4cI7LROUqFvpi6y8Tku04d/VI/wDj2uxAxEgvJdiOrM8uOxA/1KZZBXAhy6OQmaUzDGsSqAMyDJG
KOt0NhvZcWUMDUTebRCGPtR8147lZmWM1846wVyVEjHgop/+QOSoBwddriv0Hd6e/PnlhzbencIH
ZaRP09xlC919Aw2ejbYQ/SPJxBx9dk5qsw2Aj69dzsT04+ekAOQFhXSsiQPDaR/KnhoW1hK8FMfl
rWpBy40rXBfQ8pGgq5WtcOu1jtXK42RcOt0hVSkKSFilQxbnuXPCUWYhGhfwSDMjKy1nfzqj1sLr
IW9s9w5fDBsJN7wkqhm+3FA85O89OOrbUeOgyKExtCw8RmAlX8/zBToARlSOTabZDhMg9eErgYbz
Wk7Uuu5vrYsotZiyOXKyd2Z+uJycX2GZ360Xm18bMJl5Pn3ZN/3fOEiJnWc82F8ucsPte8S+MjTw
qzazFHrahnyipBbR+eUvZGYfL2WUvegXVf53UTS17sORUPDuIxH0blumod0q3FXRURWk2XCu7yXc
1SjuvDcE98/vnpGqg2Ga5aS7Gb7uSF8ZiaGUqTS7nGdOh+2AR7sW/RP0toE4zCKnv6pI0RejjB3L
Ynhhy6FFjKz1tz/+WuL+9hKSpRT7HAlC0qnAhPG62GUqQ6VXDuq2qBi8a/MisFT18wnRVgKtQm8E
vfXVzbUoDEFpLAkdwltsBB3lSArweg1tC58/7BafBPhEk5GcChLcz+HgVMSA8Ju2umYDb/MkZta2
Kjj5188/18QAIe9ADgVAVKbJ4Z6ySTfZUXEkNebxtnhEz34AdMRH1MeZgZn6OmV4kp9JZcnqfXtu
l+4qPXMGa53KJwLtppB4ym7NxP3iaYYwSDtnjcgxtbR+0Qjsi/ivGw3yBYI+dTRXQtradcDU09+f
nDXEc2Ywcoe6thpJ9HRqm1lujv/L1XaVoOeJDonn9gBs3xK3Ltg1JEtpt4q/Bjw11TlJRsaQl911
ZjA4Gogj9a8QOcF2Q2ZI1/8zEB4RGjI74aKBGcN5rWPZLgN6F1KR/zyJBvmnRA65ohz1zzWcWoQJ
nmIt0JDbbOjzQIEqzvysd65SJ/nJiVe8My+QePyCrVoPxI5R6W22DrboWPiK5SPrUTNNxYjJ2fC/
JYJfpUYfcu2DqyfROin9MetLHlRytAwKWQTKLuUHYWupOOOvgu3UvhIVjpUAo6cYWRgiosde3d/X
tJxNNb4Hoca+rZwcVdKJtKHrCJUaygM+wVjYT7n75+Xm99yQPjkPFJ5isubVUjx42RsFrCpAGgCr
AqRR+pYu9iDE68w8GlNzplooyjPypCokRHA8xmYCP9YkULnjBAa6PAU7klb8E8YHVrs9LiU+CA2j
hUDIU6l3FpRLWpYJlnIZdYro8X0yuj7pjDda43zZ5WCWD5qO51v0eyReRTgJmS3+mub5fnhsiqkO
be73WYrg6B67iiY/LkpUt7wCj9FASM9N+7aZV82HDOtxbj7GvnCsoYZdhOhIAERhMTJ0tuUx8LnM
3WXEh12gwyHbro+P50TydEa5V5EGAfC/6CD1fIvpVQgFngQ4mKIcl6A/msMS5acGo0BhgKdIL7/a
s8MZKEF0HuabCmwwHJohBTfmXKSSnEB4KZ0xMHxTwLxc2uHLZO9/NnW9YTKobLdCD1jkL1GWbWmo
b6O6meBlHv39x9KUVylfpELvmOY3boYoBGwMoQ9DjwoeUSh12NkwfbV9KwjGIDvbRfLnHgjv8U+J
aF7blS4FQ/ZoVH5PMBscLvlp27+CAdEclNgGisez/VldJoPaw8Sh5gaDeP0UpSDBz2xZPvxwqlut
kSq94pRAiaxVgMU1DIugxyp33weOBx/Vv211sVztY5+RfmbhIRRe0eGVDEymw77Cte5c604LMgDn
c7VY6Qd8q+DhFcy1T3Sho2XcGqj3Ga0GJWdW9U85yCbOTzW+HyYx6KoBQOCt4SPhpvw4sh1qeHLh
4+/JBPzgysX9bzso8wxdZzkd7zgjhSHBYLlZA2fVt/P6SpoR02dP96fktFIjL0eh97x3XAtXEZXN
TSAHLwoXXMH4IhVWRfm7W7Yth987VFpkVlngxA4VyaZkbw5Ei7sa2MMek7+kr56pYJYd5aZjliCs
AwxLPyoKqwvXu8EnVsf1sb9L13seCg2rm8dE9qtwcRXcAiS9U6Am8VfwQqUjGQ0pKOeM1XGNaIoN
V89N4XJxIToXThh6H480jcYE6J/9p0EgpQpUAzXgKXcIM3rJq5KvCBuW3bmHb3la9PkWENzo1Jq2
AIJMEF6EVrlKxUkeNmkh/wojqUuCsGQI8s9zMZWo2Mb1HGe9PZPRXp4J9HdkwDL3quI5CTDMWjzQ
1z/IkuBbsyxm0V080XX2Ba4YvCfe8uj7qXOZG33cKPlIclUO9T0yUhu5gOCgNveaOkAoe+efUgAG
2w76VcOLYs1dgZpO2tb+fY+ckI9hq3kn9spOtpRQPFyt+WHvsB7Kn7YU5HBq03AtpPQHlN8Boiii
a1q9NdTtYy2wjU9xlRv9WFbbjdcwkcVh129bPq4F5RJb6f/7UV2VFeW77bmdEfGmNS7DtAd/w9hy
P47gPtv5mH1XavqpukwuqHC3daEnKWZCqBY3KVXRFA869Faivta+Ti8YVVvN/gClmQI5rfylTurv
O9VOrlcEAe3HWz69e/YBSgZjVabzQdlIyHSmMExJseTgZg29CJeUrn1KvAqU7i2mNLqr/sOdZK0c
fRoYYYJtQJ3qhOvf0SkIBPdcJ3rpV7hZmYUoZNuIdP7LavIgKopxIuFzEoPvfUR/Uv4t8Izj+Swp
OIcB8YP0PcoX4lB4JEZFNJDxQZOosCzRBqrtQKHkzC1OALRsRc4+XSKiHFwQ9Bf28ZKAGUWcrFeH
UvyE62CHSuz6k0FcerC/7k0tGiJQ92dcnSFBtAszS7iNjiVjA7trx6R/zGNmtFMxXyg/pa61B49y
nKvgauJmP+CG8HB1JBB1wPqz0wqOymN/G6l3wvfpSp3cI5NODJjETUg3LU9k/OajSqanEV8eYx2Y
d2Ueq7tE+Vnm2JBRPWh34PV4ijNFKAAXeBa8OIGOW+Dh5+nMqgmYEgxYDK2zp/lDumbmXMSfvdIU
sQPyUASAyHDQv3ZHlf8Yaj5phtHrp6Q+YpID/qW/RALBcTD2kBQlkY1N6/ZNr4S+hThQFehpDMbX
LmeCG70j9k/s1HADqbqgI6pPlWtMaaRbszLSN7Ck1DtBv0a7x/QMm5+sJ4gDVL7OJYc4b/yECpk4
Iov+z7JfCt2OjmT2jfgA7JkOMZdVebWBUH0mrBKyV5CgnIiL5kT8yv/+71Z/fsMnLMMg+AaB9StO
cYPEDCP5bqAz2HBwIlFqqHsf8gyq1lEsi4oks6vfjLEouTDnKBpLsS8nkX1QSlsPZXbrBFuQkT7o
1uEoSfiIZ5W/a2mI/a2JnGXg15LwY9eyx3SXbcJC0edfBYJPthunh9parJfl8zAY7cQjUyvZ8MY1
+VJUk9crmYcLZO2MI+2f1x0FeBftmu1pAcMiLau6D6Z8ZDgAwjcx4E6cHT2CbxbFijZvZHLph2H2
Y6M0w5sPM6RZfht/wSQFgD2/JmdbrCI7hDON8anqIWJ8UK5WuPVAGf9mtimkX5ew8kEyWqrZwQZs
IK5JVJgyYl1OTjnn4pF2KLLHXAmri3m8MLWZVbC/4r/NBPttwo9H6e+kDGNawbZKnCXuXZxepgA6
9Ay5McmkyeldOAJddKDBAoKkfEKqL935AXXYDtpysIG0I1wdZjxDHuoGyOnGD+GmgT+sI2bT0Ra8
ydSf66jgAdvENXn+hzVXsPiPuc3aOSyP8vioc+Eq570mrPbe7E+fWllx4dLGbw7ohGZWwOTLOQUD
J2k+CiUP/IE1BljM4t8ynQZllBXcaV6UuLJvxq/zT4uTfQxpUknvCj6ovnmQP4YODUCgrvFYI4Bx
CAlrC7ygV7/RSVrA+SgTzmfEy1Ow7/cGPqQlav6duop/zuiB4G4JzzGem4nshl9ZIdIEZFCC2TXb
iGJL/kCNbnf04CWK/X+fn2eazFmj0ZWibsx9/+CEwoy+WupkfSJ8hcE3u700Cckuud2Ov1BkJ+cg
lzxMm96r4CRbCDegs9WXvL1JTCJQS+8IuZc5KiiMH3S5NBE7UrrWntBHDoafo6rm4OsKworw9l9W
2XcTEZymkq7udFj57a1h212+EMjgtds3xYqPFaCcbtXNUtux7P8HH1QoLAhgfGygotSNIsZVxoU2
SyVQ1EapHSiFVSB1aTqEUaBz+yZNqdgELrEFqR9NSaMEuTFvRRo7RtvOMugAKgG2TfwVnh3EnPc6
pl8cnOvBcOhQrjvSPW9oAw9miLthP+D8aXXEvsTX8HEygV1dgZSoD9zAKHhuD++q0F2n3Afvg9cg
ulwtWv4uWlZX65bOzKO9OFY82Z7641zORI7K9JN1B3SH5WS49nKRH2saxByQkyXmJwolKhZKgIOp
V/JJJKoLnaQ+DE2nTyRYVuW/UC4ixcEY5eKFyLLnOpHSKU3pYkDBfIOnu255cdBNlG8YZTzBD+0i
uEPd7uV4oOEF0c3uZ/9zfVp0Xo4ZDrfleqa0s6YiBeut7QxyUtxX5OoYrG6k4CJHXklYCi0Xs5Wc
sRRrirwDEahXxv9Vf+8nvLg8mHtgju2EdcFOf1IPtJ93hbz3QAzso9k4kk1wbA6bdAF3ZgWBVn9L
gbrdNbtcN5l/1wVA/W3LOLVb1nr2KdmeuIAxG5GJM88PLZ1+IYFFehrg2y3OLIpjpQuOmZV5JPzy
jaPrHqXZMfPnR+lICob4sqQ05ma+M8gqw91MJShj1/uJySEnGjNODr4UYC2HTOYbFFeRgMqhMpjK
pLpGIvFgxSnIA98NNvsTkDdSN6cON+HRxyqqDcq/wN2aD+OImmDaDU96hSCFvHqCg6wKnpODu5uv
x7oqg5OvdPhLur3pkycQ1JHAkGM/AvIdIvd6lrE3GQvHQi+mJMy5yzAQ5K37jeTHRmaKlMvX/OIM
fOJdki8L8dyx2DjWcrJ66ot0n84aV6A+j6ppiEj6OW1DFiURhE+tW4Ja3qWtTzqukRBvWLUfHB51
6gIsjtJcI0LqeqnIu51M4LMVHdxbJ+pISfMWD4gsDN1+waatKWu0DKRAZ7qkyz7bYX0/HPfaci64
yv2Hkv4nTI9L7/LgrIKUFERiRc44v5l9EeOgX5HhtMwTds3c9kdVKgQDrRCqtGK8YkWvod1F0izO
RBUj731jAW6B89Q8xfRaTwMazKhfSypZRr1xDRGgvAQ/AiKL0f3E/ssE/gc0t9ujdjLF305PSgRX
sp9/CjCKXbHNvAjI4ws4BTRYLNKQSUyOuphtqzEfBy8DuBlDgLWD6Qixqe8BI9uNFPW4vHNMioWR
glwu4sm4o6t1Y0r/B/yDy2Lebhp9EcgkA8CQV7en1yDWzbKvVDmF0ad/SnYOs3RLJfs03SYLHeO7
+8V81Cql67QuB8BOpgAiJBE5G18j2qhgDp4KTPRMdNw2i7V5Kb4Z+kVdKQYUEDattfzy3d5t9ncH
ZLpBLeAF0zoHWOwL0fJBTeeecbWMPICaT9L3CaD7kdsd18QSGW/L19C0s5lZSgG0Vsa3Rq/vvRjH
M7QINg5mQqGqfYFhap3R8SYSfzUseCQQaCql8Mp2aqFGoER0WXAoIurw914Cd+JLZr5eOZgHKO3s
jvqOS3lBCG16OLz2wv9ig1MMjdtcpXD/5igcpXJ4pJonB+X4mANCmZD0/WhMu3PdWIU+c4O/z8EB
eGHyeIhxgc781wxpkfhBclJRvVTG01vl8kICE1NiebOumWwUYFDhHvQuor6zJKITjIpHQKyfx/wC
Zxfimj3V48f0gBpX1fRS/FJzW33vlS2uyD4dUlnak9Lm6d2M5X15aRI3iJyp0jqVRtmY/5nuInV4
u8RqklM1EcpNOz/n2JgHRzBwOm9URG25pk7xhmQgM4isxX5bxkX/ln6pZ98k6W+e1M+EQ/zWBT2W
9T5zcyje4sVEa/ymg3g44ytPwAXJK/qx3iMJ6J8hj50UI/nvPcpLmzAdQn9OutBun7AdZKbsEQca
3xfdqQ3XqRaplkGgpOTxL28uBTcGaTwTGShaPm0Z7SlIRzi4usMn3zGXjbjfn8C1OLfc2AdcqXcv
EjVkvyVq2+5/Fo63dfnacUnd1YCJo/UlsBzfxBESYyCgnMILGtWYRRFGWxLiu9lwqVQQRCoLR/+J
e/iyeHfx6WaxmHxOAjVWMx6cckqMEflkVlz3NwaVLVRKpfRh9DApql+loKsrDd/7aKym5um9Hnb6
BHu/3BkFF739aM7T+FOXelMrMC6htmh/a66s6zjcLJWxelnr06h9r6xRAwyyaaHila7K+JvfspDF
LwfbfBWzuu41cc6rWPjSau4EwOEbfT0f9SzUzt2svaNjTGxxDUQvf1vVXB6CLVKo24ZZxlKMKJ6w
KgFOKVliTMd0702VzgQl+rE9TvS7VO31lnO/YtBFs4IoXKcNRs7Tx7VXyXcxqbZnhdXiZzh0cIxj
bAliPA924LRLULiythDYxgVFQdU8CpSFiuhN9rrsVFdR9i2iDsr28irah6pP9vErfwy0/Mxhkffc
9TAf6cZE0gC5F75Z9RnkFK21XesJBr734+ksL+W49+Yf1eW5TD8XjcTBUR4+dAxL+snQByEm0NDz
Ke+30d4OMeXGeDXCDEZeXk5M7YdnHbqPNcbOBGsH98tIvZJHxocz5yD3OlCXQwg6EnVMMWPmntac
pz8+KuaoLs1+t3gh6PV0LvxcaplU8mG48jIuldxOJXlEG1aTq46AYziNEJklZb87Q7OUwYf9ASvc
W66lUtqFANfWvD6T+9/1zLxCvp45shvW1keK1ac8Y60todlh0tFRUpFdHZh2F7KiRKdf89i9oAzV
FnDEQzx9ahpfwSj8uKKfO0e3od6+OXqyaVILtWmAN+31hXeUmc4/1YY27E4206FLc68pNjKsmKy3
1bpOZPHlRq3872L/2UAS72XPoLl9zvqYtpaPrXaO8weKSiVvUx0Pi0/Ti8uniX7wjwQf7TVqPK6x
kY5X+mSzeJ8idz57KK3/G4oh4djNLtstwwgg6yjAIbu6lycjAj5J6G5W2Fmaj5o6a4LByaXhvMEL
l5Twcp8ExWc11jzXR3h88dweXe9gRsJzpa/n4etsChCm748cnKW9O1YeaqKRsCYQnSC1EIvv69ia
7cE8wwJBfv62CagcdBD6BvOsrKZcw3Bjcj7iGqXMoZor+mP/XpfCV9s7ZQwLgqTtAu3qFZtrl5RM
NtDOWtn1OpSkCZ19Gh7Y+eqi2/4Wlwf8ThTvIQph5q+detbxLv6kTygU/KK12Sx4nD21O8IISd8c
FtOxdlorqUjFWxPgQQgH2lwQ5vJej7ckehwreqcTtiX45uLqlgYXaabJ+KAym0Kv7mUc1uI5mF5k
uSoJyfnsuhEVV2Sc4K4vHXJGCkxPXpmk8GSFj0NskDRMSE59vUca8Xt2NyY4xpX1W8Azor0rpYcr
ioSP6MHc2YG0DXahXdAAl0JXziYRGGhEmzZJvgohKjolOnImCBjLFIoJhalQoHHUQF2R66zX0epE
fMkbjR490wluDhzwsNHe8eOQ5l//dhHelH2jU9EmxZ8qENuMuMunKYoB/M2SLgnYjiPzf8GesDQ6
VeykXm8zyXFIM/yj0YGEy7+Vh8c8DAHkkLZ1k3g7hJFRPFUFGlpwam1Dd9dJBG3XXqQbivudGvQU
iiSE63Lzo+KMx5+K23p3c7N1+0l/Ih2tlAQI8ps32l6WzYVSNovF5/gepDBn8IZ+jpPAfPKAV7sC
IaGbESHtcdgd6KHZMSd1YMFYTmuhoP4yupOptpDtqyG/Xscg9Vvo3unZmKd6uHNj+5QqR/9l+MR1
HVxSb8tqDueAx2atr/qRQTMD9MbC3Fkjn9sOxxnYVl1fRRLp7Fl3bfUHCuhGhy1atO/I4L1IU29p
lOvvFnnx0kKAa4es50hjk9H26fAXm9o+pLXEj8EJKUixjXY07ZfPONOSgN8B4tK81Gh0oVIfFGWR
oNI2gZUCgqFD0WP/WJ2gpDZkhgY2Pkg9c5xK582JBkg2u7saqZlRf5ih9eqItqA7Fd114nkGvLDW
4AGPt+5IJoWOwytS8I+kcVgJb2o7tfHUCR9afNL9FnzCA/eHzCtmjR959MRWm+S+25D3HVI8Leb5
ryNBXuqGMcc9fR4Q8E+4N4NHLbyEYpXkDtDWLkBYSosfNWUGVhy4xZhD3TjQqKXgg8uGtOSY/7Bk
yW4LrHDQJfNKJEzQG1Z6WkuuBK7jZPzCRAGCkso2bDMJQSs+taxBXgRsnFlLQtaVHUogg7iUsAK5
zZhiPECepguERHoy5fn9y2byU1EgEFNa10dAzB8fVsYnEeJ7/pNArtYRvjZ+1fF2bv12l0g00vhO
YHMpt43n2ryWPYgPmI2bjVAdrPPgugiqABhYo8nkiUzWp1p0FwPNfvsFjA86bx77otw/j88kHnfr
84WYGpDGHv+EZq0K8ujd76DlGinJfMnpL5udKE+7IGvvgaFsw870Bsctsit6HtcDVw9syUna1HFB
/Knd1uV4PEs6FPl835xLgLhYNAx5zeCWANOGhHq5i/dRL8GDa3p7iUFdP/+v7I8ooWAzH6WBSbY4
F/RFxtGKJxFTbjmOME1Qk0rKV/cnFeBFR5Nrm1yDqNIyjTHWnsDQys5P4vP1WEOSwpC1hy/+cJeg
mJcd+RV0UKUPSZxDpdqqQEzh5j1qpYUltWyXWwyhrggneo37FzDGpN3eaG+FMVg69SGllw+sLNBI
dSQIlOZgXlCbIfYEyWkOafxu/enaAvWNoEG4vBzg/R62vE2mPCLo754cwRT4B/pBdPZiujgolqBN
+p8m/YoCL5VPsoGK7hCQrkiLd26d6lQ3N7WxaNG7BAjiIOhnJinBfAvgu95niYuis9MDxPTPRox3
aKjUKOnU2uebZdNNLECXt9812V4HfRX8nhG1vV+T+EJlAe3cjxaabinMHxkelhp+rsfKId1OUeM7
4QTJxP9yXGY/hL8HwKWXQGhmG7aVnhKaW04Hhop5L66L8PO5AQDGu3odIoIw7loXH1WWIjIWWCNn
h6/Xn+zqa4VgZ3syo8CqAMeoriKiAl8Q5oNXXdSmc1DEwYhUmwInyOg4r7RT+ZWnnOH3SnLHLBSB
xWYXXjMoH8A2iF7jC8lEtWhrunPTlBJeEEbl3ban7VHoNcG8cmkbiMUGeTf1dVcLItOSM/Xta/Nh
oK8O8fcNMb+XvKB60sjQEFhGLbbOMraIZwJFID8GESqJMhYkO7n2++LSxXJaHibNcQ9BGcRNFm7q
/Vj+uNObzwusOxhNKh0epIpoM+jSkzyKHyOiuWwFCNgmh6QCiy/29D85YYMvugQZznB8W2ur5Mju
RcV7t21lAsmmDqf/367rW4dzSWUs3AmeSQSDzl4Q0f01J/eMDc/BRMQEGRrsFMHquDQsMX3XYo/Z
CCIcKyT6wFetFMcBwhlutpuHWSC9fvhkca8xaVoc9QxN1iMo5GcsVNYA9sPjceaCN3Nj/UXI88Or
C88qOFUQNBxDoftT5dUHZhh7eaTgrTnTkjC2gwkYbN87ubj4KWy05YyRgrVlr3Oi8GfvBw5uPk6y
27kaP+cS/N3KXqGzZUflM+CahwIbEH2rfuqdY8rQe0R529IdUYZlK0i9Ya0ezxiK5pcf7UaNQH5G
YzGanKs2fO920aIidi3gLxd/fH9C0mjxDNfdKM5mubzylEz9IxiMahzyTfPbdxiRl7ChyfVnfSdg
2NX/mVLSKzXtRDpdJPfwoQB3f9I6+pdRmDmU4fgJUw0ohuEQZiTWdhO1leGoDL25zsde5Nv/PJZ7
kBrptWDQMBroKYJvciaf6B2TcjAIBceW9CYaVPEH2/3XsaqL+5fNnaZL9HK/V+bghgrJSAOkAa2F
KeNGD8ONLkpSY81Ib+8zd9jML4qUs3lDP5FkOzuc+0yN4WhTC6Kts9qT/q7rqZCQMd3dO3ZQ+a/Y
a21J9gRynvL9TefpYnF4ONpWpAmFS4VXHzls2KjbHC9b6ecEwF6xeAlDIs8UzY0x1E7odICd7+j1
1hrRWp+H/qSwN4edWcV6uZs5ohCE47ACGGNLQAPDuCMyXlopsfITQkyOA+0PoH6Fyz+gyRSD63nB
h/igWh2PTa+eCQzK/wI4WR5k5LuS2K6Xinxf3BECDRBO+AY60GilPZxBPvyufdZBqP9RijxIxUbn
9CECm0ptCluvS3NHUk96+QyJXLZHD+GGRsmrwieNOZVUdRDJOn8bDcHNphQ0L/iw8yFuyXa5+XmH
NB/lKS89ltpjKWJxk1awWjO6I8gMEMmaP3ISvcJl7jWl/Qw1C5QhMTsudqp5A8y4f6nirwfJSmBb
xlyJfRcx8+yqIYR6kFzI0CO2CdGrUzIamPnxkVZvxUBiVg6jlkRigxTPW64vOMhhcGVoUat/zU1d
yeIN7/2Dbq7wHXOnr0b3nxFV3u8VvM7x4uL0PLj/45mAzpC/a2exDrBY9G36p0JcE3xXTcRHPmqC
PBUFlfPgXNuO+meyuV3iXouCDdE3cuM5Mj1JgiQ7BSX/FtxW90Wkze4B0i9t9Pvpvgrb3g3N1w6w
lk0JJG3eWSBB1C2ZJKWtr8g7TQWNpuRPmJHhVK8dZA2FZq/k8vQppFc1d/G5pccgBSUBehu15wjf
zWf58sHycWwJgGHM26oNnkcOlzcDs8wkj3xIKAS2r4ykUroKlEaagq4Ij6e+OhjtZ3zW3bLz1vwf
SL/MaKchtWBKmqDd6AJpvD/iMocnF2Iauq5z79/UDEQeOpkQAxtMWS/1/BA0nZ/sm/nEGOL7751O
IvlSslfUZK9BT5cRuoHBh46VgflmvXGtdKwbOWVuk6Ive8BZBxS+HuNWR5zNvukvMJiw34mWaTzc
p9n6PXs9ySUu33C7doFVhJQKgC0o4K0kF73UT8OCXOKioElqX/FqViwm4NFlEZrklm8RbH7+bCnQ
llGFD1JA/BXd0Tw9jqAfF4YgywE/yEVdCxPOSWIxvd7BKAAvJ6PRf5wBkLSKHDqPtKA3Y1H9u8wM
7lR7jvQfelFNvdt0NBba41exb91yFM4iE8PFQHo9/xU42r8p6a6TUkURB1dHYxpPbC/QZ+vi3hr7
NCWuo0S8Bk0lMEhdJ87AXw3xfyUJUeMol4iVp911a6VdGiO7W+DZufiVO3oPfDH56MAckh+pVeZn
nmWKioef363wpot74oD09rVDQJ9nkhPEeb9YATPJOaeaYbR8kQq0ktKN/rg+gbOumSMeZhLfA5nz
mGA0lZaydLwtEGi+41xq5mzDDiC21/v0hmPBn9ZfOuoNVFAPqU2HloDRfft5NcTwPrQwfaRqrEX5
SlARvp1Xuvh7CsGVyFheBko+kLpgHBbCLOsm8AMPprWtCVtokrEedxkKKRG9ba8wYaWHQ7LJw9FD
hes3zPUsOeVqwGRen8xr//r1LyiAirs8p66aVGgtS1l/KsCgGTzR+72PREq9RK7ZDdk1Ub2XPCmX
D/e3W6XPFILXqPP9u2ul58u1Vn/fNnK4bnDyYp7juuDwYgFLISxjz0GlQMouqe+IkNi7E0/RlFOq
VIXyxv0U/Kk72MEowlF+P53cIVdhMF4HjGdKTJjWETuQ3tz3G/2CrTPtcZ5at7BFO/OfAtY/oYBV
ssEB/xo+5sHUL5mmMd28/N6gvtbq7XOC+p8/bZnh/3CEl1De7NActr4eAH+sdFsOgZDcn4A+XMNX
9z7GmC3961GggcaHwc04ktjDUoj6bKekmDtSBRw+/YTN4TsU0Zxs9/9T8jl+32H94wxZ/mxtth1V
ik9GFWV4rISLL3sCzNPUARd3OnnuDZChHOxWBW+/2ZE0aaMR1O2L8EggJZX86MjXzgeEl0TiAMyp
yMtZB7+7y4dRwOIqpWm+55DHeV+7kxIpQZtI+1NdxFu1skOt98AkisqKqrTQCRCfJ+38TAKMJQTf
cPME6FcEJGTnigiv7FJLDedGBbwAubVlGPfoBshw/w4ZbD8G6jdfh+lle8ktY52mZGDXPHjfW9Gi
uFGevwrQm8USXNTPvlszGB2mNXyNbkWvdAtqVstJnkhNEBHV4upaZuY+xW0VAVvQlOIiSwXTi1uk
EvVmSv9K5kVDI15AfXL0VOlsM086pvJDgYUJJox7xaz9FXnUo80rkzDXP1GOOURzVTwse8cb36KL
m9go0uvIy6Cx3v4AV/+UOhKxkvrY4FAw905Y1Kljl9x+f+kJHpNN9NkzNO2FqCVqaVwTJHU9LRRb
y77tlxMiaXX6Wj6lpep4So+xJS27g1EIiiaEYtuZNEUWKOppdnQiz9QWg6z1aEutOPzTOWHx+jqo
YqsxZHRHPAax4FtHWdWVSvmye/42WYHEe4vspb1XTRS/eTqzpCKR7VC67T/ANffXKBt5SnYlXFAM
mhAC8i1kCrDwCqahRGInfpXzxLDkHo4XnSSSTe52N9utp/jay2yN70K3PgzmU4n6gIFSrywyUhWV
+ZMTL4+R0nnaqLv9iKLeiYrjIgI4SL+kMs4TfgKnm7n971mVCUTUGt+DnocCjl7v6ZCdAbEorPbL
xKOF/lTKgCADAaDY+tLDHvGAkSJ17MHJUzp6sMeyB6unly8VLwOuiFBQR+tAhe5Z9caJyK82ZEm9
HVeWvsNsLyk6kmnH/be2rEgPLABBZes0Gh2swpgvvmCYHF0XNw4PB0EQgNVHNn1l5nG7wqF/B70S
8mxHuqakUlgUbRKVXa3DL+0Y8X2n4PO/giPztRWW2Sf1rLhTqc37j3ihC/gEhtvxeoCqNPaRo5XT
qacjcaJkNtEjtiN5r2OMls1zxHPb+Oo5ldBLKG/JR+7q66oA6/V1HQuTR9bL28XjW5Z63RWdz60h
13Ml8+23oyOyPIgahjuLCsKZAg87TEpQ5igL2WedQGygHB/QO9EOgtSTg+Eech5dDPr1heEg9sqU
pnPTqwnDeBv89T2kVH3UQDkenwx9WaaJ4O7a/gSKI+S3nsKdqrb/TQZ9oBzib6jd9cyt5Ed4cV9L
MUIq7DE3ph0O/nBqWd+eclzqR9OM5CMNrcJ+pWZ9F5c308RI45331kzAlKJZov+4MY1KcyLHfPIU
yn7quIO3ey/iZxAHrlXnLOkdMFRFNegu1hZDmpAWthQ3GWpRyuxdEkkWr9Zue7UWnKJApzx5bNgX
U8wbA3bbIKDaqmVvA70k6t0/lykDLQRy+dXmyjMqYgNkTCDV762oHtVRWTEiFvrUUpM2BFWmn4ps
stzoSy1LqzYqHf3XPJT8xtjiKptEUON75/0v5ToDxnMXgNIDGhdD4MHao+RNU3PBaBjSRcxAxAkL
+JAiC19rZtrAaHf2546MoN0yOhDWZ9DFhg5akwmY9VqudSgTTfwuB4xXSU4j/0Oauf0FKJBLigwv
eHyCUKo3jiqxSsmU3yoqKixoAectQE+JkkFHtvY8yTm2OtEQ8PTnNGOzfXlxB3WtWiJWo9efehOt
TtnETYJVYAZS7gb50u7xs/YWmGy3jV4SO9F/dUpLKJJxtTeK7jSEQNVn7mGpWRtSlPSWw0bNR+kU
34aFhOByx7l+sN0CZy+WadwjFQsWFUZhzZQ2j6eNsQTixL8/piwOGXrMGbZ/g+YNkDK6muIFJS9z
H9rPIIUBVahKZ1f8AbVKdKzk8PMwOdNRor2fc58cmAB/vHg6OSNl8lpBEXa8HjiDWSiFY3oSQUtW
Q84Demme3hdu7Ncw+NyOre/68Xf0CHrY5HPG7rFKp5e9Yw3gke/LSMz7Ao7TWsVE3VMLNhjCAKmF
HlRTBQu+6OBcRUKCk1pi80wT7wC3drjvPpHjEUBomFIgQWV8d/Jlyo4jF9xGeLkOkHDBvENMPAQ8
3o9Im2a3n06TZkZhAGoZP0uBPeKf34jgzMrsMxZeP9MnwKR8pvQb9Q7iZyJeXGgDQrSpyY/n2iDI
TOKgHxrg6IGS03CPJnhjKcdEm2rvltssXx8bM96FN4CYZkdhOJnpOn2dhkxkA1RHcKqppK64OjhG
ZsIRdjz8h8Tp2rTUVe3I9zYx4l7/gRnKg9v0JHV+InLt8SRoM2jGhuWS6QxZLlxwXo/eU1aPowNb
Re+uNyeuLDiCzF4PmtREAes1tr0sxdZNmxpSnj4iszFhIJYEW7DAV+/AWgkpfQrFB0rOuCqFCKSq
qV9beM8jttbXwIhsWhKQugDKm+zETlwlY+GKS8+9QK7okxnvEHfW0JaRk0M/60nFLCJTSttcfT8x
+w86GEvgA24AyZ+ljf9JoVo6VH/VHOIP++Eo9Wbxm0FmCvRtzuFN1Vkultxew27+KHVjnJNa1mAA
swzZPeMkETgk8r4Vn3FDO7hP/nyyju3UMzNKY4Ra2a2DwOOMFmXYXtlNjZ797/88c2kQav7rxPnh
tC8SPKeC+7l3JP1D5Zzi8L8nGt+2TEtHRnpYFxfo8iqpMIwQse6UgoxHeuDe4EO7kh1O28G+lZ7U
qA/MYfKWf6kqU3qdefYEXPpgSnM5PkuqilZkjIbJTyPTtqx2s+T7/UMCvTzJKk8raJhLQQvLYuWd
hZ5LJ4bk+MoWebrDDQoFt743x5eojPdTW8NdK261D2WBohC6jFPwFHYj0/Lsz4YJGwIDLF3BP8mc
4wyNq6GpALLbd+7fkndoKh2qc6qO0lA8VLoXs9s4inLo/iasyjli0gIQneCEERUSuyqZDYh1OlNd
FeBDLHpp9RyoWX2SQmd/hWIis6Ffr/94lwu7VdISY6dWWirnpjiDbofvZ69iTtpokNmdQBp+EBlw
lqVI0KkZvFPhglJ7jcaMlv9Tx539uDJdGi7AK9VgJOZIoXmoULq8k0jrdrDlr2Y7zk0nKDyJe9Nu
cw1Z4t1O4CYz2PbkwIxd6vo8Ymzo+xGjbPQmmq6SSdaoLlukxDvmYOqAm1X6Dm1Tj7YAfuMrh7YO
oH/5A7IPdogwiDcNbzofk79gXLVM4ZeeT5qJezulpelLfkre/XTHtE0V1Y9Pl9Ccy+5XXF3eOf6g
FVmXiuecAeKc0GYQEFdWPSqfaIfYIF0pbTTpaXmIcMG+c7YAZmozIJN+wKkJkWGoA4JYcRXhsf7w
7dnruHQpDmDCTgtRVwtzhYgRj9BLHp2ogRI+/Y3Yq+l9GP+GHOidmo0nXzTSh8Y12o//PSvsMzLy
2wpUXYu77YSaPNc4NJVQ9qBudoNiihTZfB+zWu0zprwAUmhkWgdtDWE/7F/DgIr3M6jMKByUCSMC
+oV2dRfhmfxykt+Q8hBRrRQuEC7I5c+uOPvHzXFI9uQWeGJubyGETJitTYuTctiqvmi5cQNL+7vi
Egxrvr0jP4nyAz/MpubvpCCbL4jrNKKz/IeljFleglA+IS4AMnK29yGAmNLKEF+iqbU9T1iZ2wuM
/SaybsbIG/6c6wwkHYnXxk7X7osEmxo6vVyUxszyhRKB/fe7FJzAT7WmXFu1ynnBsoQk85vEzCA9
CoLKh2IFRxWF+ggBySYo8/zLxIY6HNUZPOU7dFh4iQs2Ryd00AskSZvtOC24kHtRfqDpqd4B6NgH
ECbH8fXBhTKBXPZ1Cs91MpQkvh8gFTBD2JNdrgRpLoMXTvC/3knU3jmgHN/mERZ2I60ZqMRZZ/yM
X5DKTDg+Ck/5f25rYqqLE1A3AuglpEMifTVSacbOIjDWK+l7nC1FoBaGRlvsSvZp8zLjWCcriluE
5xq3zvg0KcFGoC27ViWWMdGE0G4T7+lfmAZg3CqTnCDerxRJ9n/sX6HEL0Pq+ro3TgYOBapoHRIN
VMvKjKJsW3JIYmtIR1YaGpyQT8tpC17jp2YwU7edaQxiazjwVYgc+d61UxmfjwNuU551fu6WLR97
o+b2yRq7LGGfsP2pgzDxiw4aVTpxb9zz355Q0RBp+ZVCkZazfTb+MSCmssxNJH5j4izm/kOj/801
dcw+TIVawC99Fs43jLmUgv7KNiYfmQelMtT54BOEGsyfkpC4fVVK7WoFLSkRPOZ/1mOZ027UnVk4
zHnA7jhMrAWjOkH89bPRmP5ZL/7DqYImam/UtvBCAR8SivPW2LxIPIczCe7UNocCyP0IfTShbPKK
cnYSIYyfOEiO/lByaa553EBr+0CD4BYShhblBg46V4b44k37un/T3O4J02Z4hmcg0WO0KK34N4Vp
snN3n0eU/ndfldcQiKl0CXNKJndswdgvGMvWOGdDD/wvSTvCLMdx8LoVMWHsxtIG+qNpLOOgiRYv
ePg7/swV6wGT0PfEqapFvRCYGEBhT3julDryJhHSdVRl1lltMxjyQAiVs5qe2sjfkxNReen/cq2o
7QDx2H8Lct2bnY5GYdRrGLqwZckSBwjV/8wHbhkwnKZDHnX+g6lNRCQ2TgNjHiJd77HOTupm2wq+
OJuA6M3Yl/3mO7JZ5MHh7qhZGbyWKXQJrPYiOXxqG9gEoCF/iFDKOVCAr3ruQKZTTMuwSwbj+Qbu
VuIRfBAD/4S0a7db1AFy64i0Ncm+J1Qad3P7Q+l3v64OCAYldyP7P7E6rlqC3iChIX7e2yU5xlNT
QkgTGpT1bK4BiKJgxhyA32IhPprLtmCbees9SNsnixKpVc3Sft8X1fjPyc2u86n4oRsnF4IWGE0o
CLy2d4X7kSHIMWNilHNtYsNThdVV6m4G84mfznzYKKxEW7EoLiYq1cXNbAqhiNk4EkLZQc3LdPlS
ENwEm5SabrpHbl7enV+0z34pdBaRXvNEmiBJ3lBNY/Pcn5WIuYSzhlRXBDvngFSLMAPIjo+iJFCt
7b6R+l4vZC1h9Ikotqsih0cpd9YdnfXp98cwGa+a1IVllPK8ChFe9mtwqMq71fu9F2HxUds2qvwZ
VFje6uRIHWxOozemlbhXZ+NO88GX7ihQDST0LP8IbVHPL6DYOFNmL6Qm4WOC8d8jPbNG4u139Els
qtDT9442qfwt5rv9ElZyZvFEjGFrS6wGM3kdTCMlfjNl6Kc26BGfwDX198dwx6EMRkebuEAzSHPp
eGKV8SFL0anQDhZQIskT1oA0eAUwLirZFDwcJrB55dcYtOtvKxga7D2vccTCA6wrJlYuRnpXknKh
vpJdxl4YNtjCh07mwpaOZn6/hvpG3i41B/gPg0tuBY8vpZCc+VhfyjJeySqxFD9sZg5cNSua7eun
1bQKV2KuVL6H+IJjLo4B0TyIs91qoSwNIra1VDNtYrIt4IT8ZAiLZ0xiTVU5SSfHUUFrC5fczfqF
uYEGQWDQdMvg4YTJ/2ccP1OZDHU+UpRtX7wyhcmeNjo2EBcOoVkCEabtXiL0ESrxAscZGGy2tgf4
Bp+he7Ooz0J+dW0+rFIuN6K5CLe2buAZMD+xsUOI8NLtqaOBrTXaMenDE5lEGZx6onIMZRwYPP1v
ipFRSm1fDHdEPo3iqbbCKG4zpl+rjupO2CRN2B+VDrpyrf3ZhZXeY5yK9PN+SYbplum/fbSi0Y0L
WMjgfyISYtwCS+wea85XAPfojtGEXgSJcojKdLdmx6QNMAIU4lrm+E9YBaq3xCFo4VJ9HB8fRZfh
6i4hXf5JSZKzji+zCpOkjrDDNsY3E6IwWmtVJstuWpYwJMoCNjudd7x0Q1RWaC250LKxgtJ9K2LS
25sT/rgj2a0RwSXBBVF2/jOOjhckUtrrt1fx1h2ro05Ad/HPyeZ6GJkTobit8ndmz0FOi881uw4T
XShY61ekYL/jbXruB2r1Ymee4x5qDfmXnlNeyoqtCScEWDumuOVFHTgqnLccoW27ZrtU8PeZyIEu
tq2KVUyiPFD2mBTOUQKb8ebMErgMO6DSSQB8GSW6I9twYA+tQ4XHlp0kTxwq3sW/l8OyRsx/8xva
T6EvvvtFl4ZE/vPoe4mBzNZ6MtVnvrtr5CjnCc2OU/lSQHRUu8j+vkfE2WMAS/1CyzEVnnt+S+3V
MbBY+afWlCaedw1/9tVUlToZXM3GslIYrdfr45mrY3O6xzWHU3Q+nLJFWPcZuf0f3RZH5lbUMbHn
LvYfdxiSw+BLRKPU/nJillAdB0HtXIVxmh62aIhN5ZlLKpw4ffiL/G8yK50RUtkeJ52Gqdx9Mj8I
IZYgDfi/i3iGBjCOsmQw7s8r86gJUibQUtt9oyV7Lw5bkn/ASAYhIdYWsCszCzdHHT5h9lo0hmhq
bkE7XWuskRlQMwc2jE0FKsFZoluOAeKYjxXAc7WMyLCUcZVMUbTF9lX6115DQV98lh7QeebUIaVf
/IG+nFKCk3xvRNt6DZasu9lbXRqAXXOAzi2gYf0tbFhwcRAkiDcJcnPYEjYRaZEg/wYHOOjpALV2
8Zbm6QLRlb3oVy+8RTP+jPLRxqJQkbYOiBdQKUOYfdH7OABmBAm39jo/Mf8Xl8wHysevxASf9kBv
VYL1s2mCw32wnE4RixrAyTBz9bANnr/WusuRc4/uQZ4LA3Rn2FYJ9CkY3fnIZLFoorB9WpGIohNG
TfLpgBjlJTwrtvZHsVWZo5CFcrUDl9ojZMbor0s4qf8bmDuT3unQVCYsRMAfBYJScaFfEo/4cii4
YzBxz10fXRI2q3GEb7dI3y/ym/T+Zbp6QRdR8DQOnb++CE8xyfujInAiHYSqiYoLp6XBhXx2YEtA
Vq+3tAXWFSJfVC1JuV2Z/nsl/Q9u7FQGhVX2r05S7IvW7XKFMnEH8LdA+M4HI1o2F5EMEGGRb8Nm
fREfX63S76LXaOPzFVLw2zbdhuOcCS4ZdTykcUBDadfopa5n1NvJfSeI0mMWmQzwAQ+3383SioDN
ilEYsZgP1fa2LE6sAXgS/2PPleFWCD1Ro2D2vEVcb6OOHtsvKLP8kBalCcm6sBVVqUQSdoBupHRx
KCfQB4KU2qsPGqsbJyQgObYXtl1wq36IegsekYIt772YirOu3TCM0oqiKSvnMPsEon331tX+OFYC
5X7vC+0fpNdzcJvVppqzBeq/N26LVcRMswkDNEayciJ0+yDb6jitUhUJWbg4YmBiTbYE+mVI/DnR
TVj65umBchHKRzgSG7ZmyZ+427zlpgAVBPy5IcluJjWJTJxFDfVs+9Ub87EjqFCRcFH/oo2A3DyF
AVEh+/Q0HTi8z/JHpHD/rKQKFReqpc4/MKGD2t+NTs99hk/oO81kRK6j+8yg0Y/oyIvHdVIokQsY
fYaAGCm/egBWDDa8fOa+Xmm0CtmroleGPxqxqbBL6/g5d/SxHEnFE1PXM7sncbXvi/5DItyuvzmM
Ihi3oyci5kwjdUhoG0I0NYnKh69yKdxsXFIeqgAh2He4MsQ4RzQzgrS3xy3TXIbUka7dgR4ruB2G
mX+vS7QgoXchB2x1d4mme9dybZ0nsCeo/d/KtfyyLTrhiYgPz6+2vDxtgWCKjaZ4xo/8h3p7XTH5
pZekUoWzmo5gxGVOJIah7SxZSjDWZItUx7TSvZ/UZg03YHOqwFiPBhTIEv7vZ3aIlBJ30FtSHFpF
fFuF406bcnlkBfChljE/i8YYGXaZaRzM7pLj9shaaUv1Bz1rK1lkv2f2J/AD+og33TOj1x4a2BKH
wQXbHdGU1gvEMnyN9Nn2KjAC4rMIvDkfCRaV3DazVi+XdBxQxIqsS1sy7OBgVKfEGNpt+0kgyQOj
NUjAclV7x6MTJ38gJ0jb+E6Uf0YojXfcy9qkBcFxnP3U41H8oK9YLM/bYitPgkjq09yGo8SYBkoM
x+rKP82HB1zuQIy/fH9kMG7n8PAs4TuJExx9qhEHVD2cDjGkb+llQ3GK2Kuz70k4GpDySABJ/sss
EXblYK0mVXaowYvoQa32x0Ys7cd6y/sG3t2v10GvHUq9invWlTZJ+TX+L/AxG4I3O6dB6XH2+nht
5GXHbZw+u4pE/jTR2prlr3752QXIEaV0ZPO4mN1IEAF+mtmHMi2fqF3RV8/EHXNS2S00NSbjtl/1
GcKB1N3rEN1tkmpnIAL/c1Zr5RlyJHZkmRs3AzpyuwxXJJMDm0tNQ0CtV140njyJGyUMg5TuBDfw
YJCC0yEsF8KrPiCm/NQJp1TdPPsgul5dLISxxCTI/56jO3qjOT9/Ui6P5ElAa2VJGa8N5mHbyyjz
ugoSbX4ksFrioeGuTFfl/zs4DgCjobyHthn7HDBfTgyuGbnYIT6ud8xxdgb72/M3YYe+jkNNS8wk
e3Yu4ZOzMPuQheAL2tXZE86IxzL92XDX1KMLwLcJ/upAegsB0SbedSsWmnG5f/L+CbpmDveVH7UY
dAjxMTILpF0g8QrePE1N0KPyTtZswJdzR7RHPTt0BkuFTzgueZU/nzy5eutVge7UFRCpq1epKULJ
f9idcAkXEgO9rzNq1GVBYCPwXaX/JMUfzUk/1f+3s4Vn1jSJFDXwvR39AcsGcYjJi+LyRoZk0uhb
uXhFb5RfqgmRYNjPO9ZShZmZpiDX0FioRTuBODpEDvBpwqK6Hd9rWCVdh2If1dj0uy4UBd5MnNkq
BErBOg+b0cPSFbWIzxOq/oBB95KG7HfLTrdN/dgt9ZaLK92pOdAWIXGD99FtQItjbTu+P1J4qLKz
6EUaRM/pBVgGoieMXHG8A345oCFrF6SufAIek0g+ajlv5j0pONctkKBcYajvXAu+daBylC43oTwJ
76UgVIRcYAI47+r/QG4V9xQg4An0U+qldKJEAuuiOJ/s2wCiLFtonfCNSoc4c6UwZnL6ybuqqYBS
92c651Fnao72abiW7WJHSKQvrtrHP2hbD92GHLuWhENrrgW9PYsj6w+0Kly0vak90wPE6wEefpNm
OQg4gSUj8nDHQYScagTM0DhOyub9xKclugdkMMvkrPtJ4rtjLrW6nqudLO+HZzYazLJ46FniH2UY
Ux0httH/FA0WOhJCb3rh7tAf2Xn+5EeNr/fM5e0rTBbw7MeR8P2DjH7A4O6bdk2wAGlPjkHGhGTt
oz/jPJHmIK8XC+hu9WfRCBRYzYff5G9BqVcftBwoRZWGLzfEREqgmZF8GCTyxL1I5IxD0bQDhmS5
+5OwEYqN5pW6Wfl/au3l5lkwpkQyeotg33TGHbUHJOAl58an/gbXdCdkE2aJ8G+6EsTzJcXEf895
wfMzguwJPIhx77sKvVDwzVlmJEpQLk2UkJHddqEHXYHo4PXpSptdKF4mzIWOFcOM4f29xEcCxPgg
5xzgl78hOxGVZ/gn3pCmWYecw/wgMaTm7htl8g5zCBQ+d3QnIz7vJm+wyHRxvmXFth8mptuFx++j
pTL3yuTICN7lasyTVxaxoxmFK+gN8lP+SUmIW+bTia4OBg+l7t2OJF7ZbdX0ZeLPDINMHQGBju65
slGYuhIVDPRR/cZ85Gga+yGBHcUrXq4BOuET3eGboIsgHRtMQZn4lia8juHbVVnZt3Y51gkKAkzL
eFiTE33+6W5nN014MCzugvprAjVfG9t8p3s01mZ2irVmqI1zR1RL/+sBQOW3SQtCamx/OyQoWGjV
NK6Seer31iD/wxyNb4gpEoyCpRx1nrvKsrpePkJLhWS5jiHarjTgcZCzFir/mPt+iOwtx6pIrbDN
eH1MzXiRP5hRiTSul2ctz+sm/2GllN278iUD9nKpWOsHefi31sv+zT/3trVZ6X/cWYcHpuloQZxf
QfJO2Mx2rzaqE1qfCztFF8WLQ95WzNjjZx2UUly2g7yj4SJXFIsaQQCVZVy39vnCwqpNG7F/PWhb
rwuE+h2ilrsjUSsACqtWsrUWTJAqg6qcFXiPi562bXoIqYyKSizKce52QA51FSl6IYdvdSU36KtT
F753uzBcFU5xI/iap2kXsopdJ4Y33R8Dp9/dosm8ycXcOqA0awD1219yecZ51e2NRXfQruvu43jF
37xeb/I+NMDHKNYBL/w4PyRyc1FJ82Xr78Tuk5WfM0aONzMwiS5fxUB7C/PydmAufjgPWCxntnFL
wdF6o98j0Q8igA02vgrBTHN/5PiErkm3VYoNLguHf9u+gF6yt7zo0O6PyYvef99T/XiNYslIKLTA
MPI38ZvDllc4Vw/cQruj0DM+36MZ2G3h32zaDOvR0E3NAICuHIztIKiDCH4zrCUelj0CtyTpLfAm
HhodC8OcZDFjvqKf7vgd5iBsZHaaKSCjWu4xqvEjbkD7fb6Zm72dW4hqbeg/CNyyA118PT5vJ3Ek
RqHzaA1KfvvZHidqs1igVOj6ZEodvY2FyeaxBZ4IUe+cBkBP7JCQ7XYG+G46kzb0STnj/LnY1ge7
OmPJPqobEDMM9Yd1jbXo0XCs/XhN47zYvP2kJMceA5lSki7BLsW4BifAnewzlqyxU/+pQt81mFfz
4VMSg8bDnjO/7UaRwuCEeA7j44EO7jhqsTbwXlpDPASPlBiWFL9khC3D4nt7peQhDzyI8HiRnXdL
N/ORCDNmZJplnrMyslnFBnrxVb3PpXGTx848vVTO5JqKN1b9jp43KrNBirR7KH3Sd8h2GxTl7gun
gciqy5vZ2BoYHIDH1wlWQ6i3kOVjr+olPJEALu7pzWAvuAHRS20aXxsszZ9ov2zxzCF52yXkIZBI
qxQ2ab+yXFYR8QE0mGrrNOZdZdP6JZpXiHlYXvi91vcwAYmmfnebWa4dMoSQf9mGjA1YZqg0KklO
VLjvBR7ZUDmvee8lXMFznEUGJZAJo9mwW5StuwcFyEd9T46CYPAD70Sfi1WmcC74ZZed09NTaWR6
LI3Sh54xAELeFsoRovUyeCIg2JfttZsM813d6+ccAE8I+zs7GPBuTz94t81co8b1PrwVqhXuD4/Q
XV5WYUSJtGeJsbnbduXrA7BhJh05X3VKfMZIxEM7Xrer75M7XO3pb5tlJtTkF5CFy9DwZGEWeEXB
y8xlIitPaoPLZsECiS0XZKxJvwgkkICKoSzhxg4DSSj9m4LaDXOT0M5Mz4fxB8+UEBl87pYY+BMf
f688puScee25BUamhDi/YdyahLAENhL5sDhnQ/g2SuBn5DirSVplR1i66wRfv0mgj3x7Ibd3UScN
L0qDJ+76aZLsR/j/hwFdtUvef4zaKmxdHTDRgCzpLsutekSM+D470kZwcOnCFIdvRFdBizqGjBiN
wrnfRP4FmqLSp7dL98DBoVo2UXFfTr8WexKkuLTdG2Or2okZLupGenYrJAij9Fo5MW+IuXs1DHxB
Au3QYtwwcF4Q2wK1v7l2RvvmjChiKi84dpu43WIX7T6SZ66vk5DbL28AGAzgBRUTd5TttldTTb5q
hgjCymQEkM8Yapazkysk1DwahwIo5ELCsQLGD62xHRZU9JnQSAi/mxZh+Bcs4rhqkRbuv2811WM9
0M54QwFA95y6XGyfxkXwQ1E8VjB8zY1ara1NSxCUYLeNNZIGAbiR7Ce6ysW1lpaGqc5hMFJf1Eod
gJyh8IoehiZfxMnypw24WcMrtnFPQNEfSL1wTUt1aq+f3l6W6cTVCtZJ/Wox1qabCr0CT5Pprosh
gffFT5jlEZoGAOafwyMoYoUrEsbHkM0jR8Y5FWnJXc1q90qJJmpg6O4j1JfBitrkLZT4feQ+1oQL
Zlx2u43Sl2WtziQOd7zlOJ8Oeaaz1jgQqB36urgREFA4ZLzGondQ8VfCLflPlExoy3Tr6KscK3KD
4XXeRd9SRB48OqW9vu475FoVxzrfsavRbl8Vwfjrb/oXefJrDSesar5h0NR18eVGWY1QBFETowwL
xVcL9XBcgn3gnoaMkLBgHz24PiT7Lg6qKXjYRQUheTjijkTAUrYzHIC3ZWVTiKKbgHo2zxsNxcYi
GUxd1gfcKADcBOArYc2LcZcA/cJ7UUWHlRMj7kfWTLbat/BexAjYHZmUFLX5oUxEjISbVhDlrWkI
RbvFuizfI7w0DBnGRpAxNZm00HMyjQHVG+nimhSgbBoB4Q9/rnngicnqUVlpO0haS8/z0YCs3cUB
7w2Q2g8TU8sXZM7ux1f/JcHvsa07a9NorKbatcYA3Zzsb8gY7/PoyDVOT49U8vrF/eVqwRmM1nsL
R9ZXXsz6qar70fy1A2HnMJ4Wf6rC4iUtTJ2lMzyWv17VJRoSyUBHsOOl5WlWuZjmwyd6uJNN3DzO
izpyknxmuiO3ZSp/YOiVkEoXBXPwRRWaGTcwP7fgplABA6qbrgjKv5RyE3DQS+KjIFI0DCDsLxRZ
VpQ2L7QtL6S3OBCDsGPmc59FF6yFz1Iv7Kh2iUEoGqswGZrrybcFsx0Odit64N1/VJkcavLr6eD4
AR/YArf/b8Vu8YE0i/vU6btxWqV6tzzVslFeojOpwe8smVpRMwnh4PbccDkpJ9Hzwn8q4/tJlN/4
Q7jPweLpTsNlD+3qg+Vg/rKi+jQJUGN9mb3bWZ66uHTDkSD776jnh0J+U2oH6kdjWmJhHM0jR+4A
XoTNiTxCrvHi9uO2NTdSC/INM4rqinYkzodk3U7iXrVSW8r0bdKYQcmxaZcmzQZeBhBzMWKU5J/3
oc7oivhXQjc3a6LzpjiyoAco4IJ6YwEMddmwRkPl41dbL8g8SLoOxrEvxLobcu2o8vQlYxnl1CIB
Ad/AhnFYRBfwlu/h66GKHbhf368lAO14JUh6Ie1bk7hX87tzqRXvDK6UpEvrgXAerdOIWPa4OUkR
FjpNRR73TNEN2LfVyEdbpQE3MacKA6zn16261avaH2wssygMXFkgDMe9B9Fhm+e4pD1hOcDhfRHb
uU/Jk//F7WriFct37cgnCbPtkM/FEjQergLatD5++Kmdna2nPs9HRm7bHzPNPR1yE/zY5CBCav6V
cA8sY1Z8rFyHMC/gXhwoOtp0tgrAQ5FpjO83h/hqADbtlDp/QARQvGPqhWjJj7V27/2uYC38jLEd
Mgpjkg3VIvjYHFAJK/9n8lVUl0R/NLCm3NK36LDjOInLwRtlsUp0JlP/iLbP3mx/m/to4lSVnbPM
nvu/L1SuL6bijUM3HGpS1UZT4XV0C1R+a/AduELZwiroxkSm/6i41mlSJUBmZAROCd4ht2E3POjm
wLfy+j62RIftpakEeOIKkGfiV9f2MbM9y06zPG+qZJIEIqwCkizrzu2bWKFZGMuLvJKupLdhdlcC
XnFeYzFvSX4YTenesJmR04rX8NXXFQKku4I1xQPgZlVKrgnrj7RbxjNlSy5vV5oZr9IW7I1J8T1G
qeyx9utoEqX4hNVlV3FUFuW3m60C+Wg1R5RSjLFozaOiDzF6pdpnr5vbUOeY/l2yENxfGEC16TPS
PRi1gBztyGLGLUVQ3YYHVedkfMxsTYOs3qmeQid3+XWMxR85tUh/oAitk+CPh15d+HPFuqeB9DnE
5PQl2EL7VRatHfl9btzcVIdCcEIE7GmeUhIY7XnbybuAILCRiY4cjfjG+LRxuef10drsQArccrEU
esPjylXlx5RV1infXA3uScwEz/ZqFJk8AXgRDbiB43a35jeOiiwSEnFen/dAkG/AtlIcckYjHpZ9
oKQIq84pePKQBYBfBMEh6oT8yPKYMoVLAsvkhqDAgS+fe7riAPghBfsDfExGjdJrEDWj+0QTUIqD
M8PjBKWzfrHPEt/d92xecxBrYUhH+aXpYNri7m9yV/d/XUvj/cOGAqbS8yiaijUMWpEChEyC+SFW
cNvMgD8vJq0FWfrxCQ1+LbLzvZqE4ccJGHubqeOKnxyjiTMomK3AVWH918AdfXrOBnBedwUeym5k
T/QWNXYVHWyCzTm/ZPWOVPjgJf7B+LnP8VhHxqpiUwTjebAI+SwwxLhfdr4cMr8S/ydR0r5pZBP9
IzyqAEb7VQgq8/pwkLMm3t8tzQhEKy3atKfppRZlqKb1HROlGAhZVd/6OELdciuhTF/3EAL4mQFa
8BuHBKfI1hjnzbEq1TA+3DX4pbdtyETCDhIPD9zXaI9Zv6ywNfVJopmezPmxlLB6l24h3jE3rIlS
IBU5i6zAVOrpZorj523S78ubLs7vCDP2b6gn40lhJEgfVjyzILCJx+FcNwDhAL2phfE10Jk2K3T0
fsMgtRLgG/n7y+ZtEF92C2GK+67I7f9gNEm/1Pn+SBTF3k8fT2JBTwJCIOFyifjm9tIWmwTL4doI
enUnkABruEOJLLs7iD8AYRngqwWgMcJKDpyXZ7P7KGaOKegxKI1FJX3rwCVdB55WX7mkSKb0kUA0
iMibsQ4aow2i+ZCPVVcsw/bmtGlSkCxddOZx6Oy1oZfrlg09yyCg4xtLQ0+cpZHZSe2pApbE+iXT
bFXOlAdVdVZS3Rb2B+J6nqYmrHvNLvwbvz5eKu+6dVPE4YWKCNFS0HhHiO+R/9YsIYnqp09X0wWA
ZjKeioj8w6HeUZ8zysimo6ppb/P7pWX9yNU25bKTqY30Lf6oDW9E+6jitOvcUKNc7IicrSHLOmUR
JvcyIr+///qkFWd4poTlf8oZCWlyBTIQAMaOTK1Z8h6KEeD8iiajgeDeZ47NlX5GZAV/sm/CquCm
XyqrXj8xzmMPrQUGYK2H+9CSTAu4hn4JgWvkkv3eANadbwhPtD/meSpuW8J0VqaK02d/egjppc4V
oWv96ccA3/VsyuHl4pWoLgn2mWldbpkC0QVEqX9/hCaIAlWky/LHmKJfREZ+nBSe0AL5WB9BxRHB
SNYZdZAlAa0Y3HhLJ0/UgNOa7IykP6Z2iTtbZ7EWFOXBn5CA+PA/QHF2hyFDEDzFyeAMGXb9Wlzy
URAmybQ0GjfB64go6h3hU6hcmaNLQOG1neaBgEK7m99k0Iiyn9UGASlW19xq1QlykXefVN8jW/+w
/Ct17btBiZ+g4Wo9vvCWIgPP2CM/nuH+ejYao7L5sJMMVPLSkwPH48mp9JfAbdOFawxdiPiI3Nde
3pIzu9KSmMyp7ZCoItZLE6EGLDOA3GwmTZO0L8dePk2wmaPN9S2fY5siU+UP9sfQIDm3bHopmngn
VildGPWmtrWNRIHcWBrGooVo62s3wT4jpkq1enbDHf2fBIGXwTAHBONdO+XGpqzw7kjUpISscxWI
ZdJawja64wJjBPf2FRcEXmJWSKy9V7eswhSBx/2DUsMseyoigdaNXC1KQSYerxMPVzleyQ7m6HiA
hhiyQmuhG51aOpdoQSCRqHbH1yIkBRADXuLL4y8dh2CFgKCR1l5bCcIwQAk1yAdooAYoyGJSS2p7
YVh/fHjcGxN5HrFdV2SPB0biYmUvotq//HwTA5x9TCECKN3c7D+MuAL1e9ptm7Bxt4MzxIVQrhTv
WLiJj+NU3JtC3n5slE0FmK2XyrmT+dLORu8wZr8gN+OOUK1ye3C+RJLmDQjSOFRSarelret1ac1W
fS1BxZHFFRQEp3bMKQD9/PJegVSlum9RaY8429Jbla+J3/fizIwselwCtwdCNAENYFi0p3vuyFgp
TnMlkK7lSWqHyO3yTf0duJWHgLiJrZtxKfUH8YF1PGyJA3SApNobjJw5iZJuf29imkmoe25j2acd
bJP7lgo8Gftc06iTvjExdAlsHP4wby3YGcxLBX41amagHCOZYVPdy5jW9fWoO5GoVm1LV8IPqxO5
tMhrZAPCbfWa4wDE5gj/TXxqs4zwN+rEiXskkAx2ILoq4bEAnX6ASfl6TnTEqVhg34ZgeabPpH1a
UyVvcyBvl1EZRhY7Gy5/9hmkFZfVPCzKNjNT0IjMkuoBDHzx+qT9EhRRnZZ6BvY4UwpQILFGJOhz
OpXYYmK9WnLJPDCMfGAAZWOWwcPL9kCyNBysXDThJ7m04MAbGI0HexyuZ1/Hqe04LruNZ01PceVB
l5rSD3Goo+QrmoSxzPn/GOvRxZA9Ux6Mlc38+mYNEfNd5lkkjmqqm/NHrT4ID8P/Bd6k5PPWGBZk
DEp0/hy3LOUg49bebSw2vbHXwhXEl8lfJKXI5YmOjFbEAaViYFPNmaSSD/tiU8HBWKhg7lRT2ikB
GNIe/GzsNVm2ZqqcfXmowwIsGvCWVbwNbS/oMypCwE3P1c0GoJkv/OVlTKImtVSqaIMG7KJ9SqLF
ofsb+/Y0RncIcJ5TxEbe8CBLKCE2Stp1+vP22+qZcx+OSKWKhU/is6AHVV5rPR4BeggXFecQzd5Z
pSh+PBQydU8wK19PSzi21+N5AYG4lJsGm5SvIVjrw9ZGI/pEHAZ+qE+0IuYvNRyhriilPssKiybj
DN0y+D+G1buYHIZKT5fXCSnK5an9glsIUMMMQdWLSTRY1VJSjz5GOSVUQs7IxlaFyyokUVJux+iF
oCzXVxjlefD9wPERYfphscGJ0P2goqIHzaiPIBzZhtZ5tGv+3BakUg1q8plL2+c2+CnFy+yrd5eT
Ppy7U+p3tdCCOy0kM+NPOxfsttktREJF3Eqz5UKU8EXAojR3RCed2w7tV+604+877UgZgK/YgMcT
ehIn6qy97mHl9HkrUG9jWYFWSmEjKVNG2k74qCTPqaivKvi87NB9PxUrWA8cT2P/8Ej0Dd6FLIBp
gipfM29NZVAesdoN040tkJj4x+oVzyBO40Dw81XjbXs2Uc2iL7c9+/KqR6/Tv7520v1SykW2ljc0
PUGpjPO8v7/PhE6SpMMA0LMIKH99SB2BvgfmxiAmT3crdyj7a8NnxfUckKAwTcY9B9T0cHVPNmY5
aHiAMnOgPWFufe+L7Bo1MkibHWv9xGkJb0//ICLugCFNbXTCyl4sREB8QmRqerRLG706P7gapCHZ
XOH3zC9a7Q0DQZaMkUFOZRFj9ovbkQlre43yPGyjhsOaom3tPraNuIwWDsMcw7WIWlV+Z7jhoIlp
BVZL4u7+OjvI4OkbUf39RArZSprY9Nj4wRuaVugnFU1CQxrZMJYEv4zvfVcFL3xYgLVOGDzKmDHq
PB7p6rnIz+K5hMMlSBEslhsVYNB6f2804hIyOcNmcGs5vGTwpgys2s3BK+KcyReRqDztKQIUKf16
ylV74Yjb/WQy7K5DJEw7BckveiVMwkIlSrzDeHNBxLDFv3T3+zangzLbl9JoKw/9VrQGlVFgH9Wy
Y/gGFQeT1hz3r8eG3Av4tpoCgeblL6q/nsBpPrrsicOeSjeg5qh06uBIrSxWGrAN+76EYmdJQpkw
v9xeEokb2FtGt2oLSbwbf//07UuOJk6yT/EyihSQ+YheHfkyp+zJcNicbQ4dQPOSj49fOg/Ull3T
z5dRobARIgqBnWjSoEqySsx82a6260MqImdtyJ7D5oc6zy+PYDC93FySo/Ate9Rr45wcABau6fxu
1VlbBhgpqLGedVjZ4VAavhlaBfitpDrDIa8gmTEeq2T/ODnhmT4KUPyQKxC/YmlzM5lFB8i/5MZq
LQzioEg2nuiBOG/xeV1JJfamD4YrsY4brpoIe4yupQtsdqxDsrcbRXKbSQOg3SQBt8j4jHymWoVI
EYRx0Sh2a4HjqWHJAZYN37y0ZM73OLY78v0SRtkih/bHImJ3z0Sq/qFx3pJ6dF4OyQzcysyVIEPW
z4AR22jb/ouTnfNIRP4abQJiayZ/+ap2aKBsiDxsMntbKuaqyl+uymLdQuJAGiH/pxF/5/7JegG4
6szIbzOOCD46OUTFuf3UiCywGuUb+zIDBK/dFFvzRHieoczrd61bzOch67F7g+s36wfdWPA5xXzT
VGtu8PwJbS4pxh09HMYHQslh7D7ocisPfsBu+CNJNnn+mgkMOaK40yuagI3h5pn5GHe1QMaRZIU9
FaDbLTs+Vjmz/8v3ZqYpZZ6xLYc9tCaAeXfOIJGlZti19vRNi8jZalwxXG7AAcPBTFbebu1EKYKO
RdDEz+/PdBUXqOiU4AKpfORPUVRzKLCOf2lh/WwlmySmkzz3pqOuoycN+UEooxq20yyGXujgPj4e
br1lq7Iz4BJVPzTlNFnUmWlX4yiAKGGdN/qNpFOVyi5acPI/hTz+HuW2CZ3vZ1byN/MBetVmScY+
S3CIH+iMAG9Ex39i2OpmshWVTqqPZc4kMqdP47/jICuUkmywIHkWIHiOu+MlJpyXEWTBT8mjdQZN
3yRRgX4m2IX8IlEmKyO6zmChmlefUH+kQcABmXM/YDX9kTC81aQ922+rDTvQYcXEz8PQwI2YaKbF
AsPAUOP90GzgCGRmi4hzk38g6mtOBdzjHe0MKfY85xybZQjNlRynnSdEpR+Npzu34KWzX1VGrQuT
t4HptAjdGUvTk1wM3mUBe1BOA9vQjpJkBGd7/JHZDGb43Bd4Yycd23gMYhXjhTZplzSNCBTYyrWz
I9roFcXZvJeA9SWamwHATRtmwuwSJWJcil+rgfPolrlM1VWqK+n/g/ipXZBC1xk/mwCuKABqars3
Y5OKNLjrUCxYtpsSq2xyvc8y7GyyJK4AcAIpEuOyf3ZWVXHIqqkQioMMeCVk+ji9PLkZdVnp6qti
jtDUKdJn3JNjkepV8gdtqLlqLu2t6YmlMeSAtEOA7QmOiK/1YUl4LELv3eOoZBnBhc6il854mmtQ
Sz2kb72zHtYXp689M6W9rexLJh/Z6D31zMmtppXvLlF3QDoqPYxIIzMdsuTt1XQinLL12y0mx9bv
m9XQ6gq5cggOiuRyWPBEuXnBAqS5Vvz4OZFq7y7nDkIBs0lGcYTnrY3RERYXTnJ7pRxcsNCoKkLq
x5O7ZEZTBdb6paryTSLknSF3a36cvmTyXQLer9v6c+bO52JbyqxSZdLB7uljs52OvpiDTtNJUJsT
IptffSkvn0gtRCzHk5rUYVQnsQXiVZI8qshs9nmen6b1jFoLhlGUXsnQ5H1LJEpy1lISpFLrLrnp
6DYfEFU1CuTGL5cZBIgO/Sr0zzBKwl6dyJlvvs4MQr8jCu5+UnR/syDn8nqbHvHO+n2i1P+TboWz
i9V1oOEh6iCwqaSqwWCu4reVJa/VPSomt+39ObsWvjWr8x7IMAX6STuM+x2/C/1j5DNvUuyaQmSn
KhNvr6RPPJRaNu6spdOPf/XthgmBTTcVPPS0tvhD9VVIRjFJDrj50l4sfc59P9JSgonPaC3xijrr
GHRCbBC+FYuSeMNWYU3TyuACOPbmNKG7uUrTtYUWTVCRu7pzuTEb+jizkAvVJxWO14BnIUC6EimX
7lSQF1oKGpeEipqia2QpYjePaQbZOkfUbCQMpMfpItLrkWwREWJMbF8U83CWeByixYAlr4a3wRSB
/r3hZ4A1A4IfSWl6HLE91d8yBIqe9q9PUavz60MIgVhIZV85QtOS8WKDHMGVnNzERgoOG7ieEKIc
OE8Fnz3NGyoORtYEbQeYJ+G0bULCyAGwD/TwcJdeJbw8wfmpkgqEHDtCpWElrYjyPjiJPBgNOctH
Wn85Bdh4zUGFRokPokqTB6dYGIFWqJh3IMZ8LRMM8azIYl06bgtNOD7J5BsC4nFA67quL6G45iDL
BSu35a7pyXQC4BKjDrLqo9b3pUF/U6NIbN/nLsDHqwv0DetsGjwWjOx9fRVsmZSr6UWOK71Lkgp7
c7pJluTUB86FX0C8y9L+AB/TelFLoP71EPqT2JPXrLKh7MmYnSEs8p6cvUOBqwvnMovPAQLPBhQy
1dJnohs1SmTXbHg5bQAGjF6uYf1kZFh8DlIe/OqO9YRli3R5ftV7A1GajXjVJlqh4j/pzf7BHXbR
LOpcADONBiWCHr+PK2y2Y2Dvqr1Utc2TxZaVUzL0VGA5jiDH5Py8MTWjg/SrYTgKHyPggkB7cP7d
KfeRbyotwS+J1mF/pZHcO/ahhogBbPbxyuHUGkNZWhIQARvSAlzne83hh6F2rvHjsiW6XSdPZJ9j
AFT8krlwhnyTrOoeamzYXaMri/rXRUHWLl1x1mUTuCxTK7CFCjvV7pngXn4FGV1BfLXuQZlQjvU0
q8Fr5V3KLs+vMMZH+HPvPIZXh2+fvoe+6HT89rZ0eRKIez8Noj6j2jlvMToestziCBWcWOXTGyXC
WwsCCGi6Ts5SiiNmT4i2WfF38WHVUmh7ABWocdo4lKV4jBHqYAlR8gXsmfZpv5lcNx6XiBbHzamN
4OwCk+Q0rUKp2foDSWEvYmx+RPodwC0ECJJNPNfDd8RnmrYi4isvQ2IilcDgfwWOmU4UhpAJc407
GnaTcMKjpB5VuD0Y88oBjrCFo3+MZ96HNMXnvhu8kbVsBo+Vv16ysesZ8TeTDlCXtJLR2py4kdGl
lgCzrLZ22vSeWGsSeERnGc3D+Mx7PLOE7ybdDN1NVBZak6OAUsXFbjUCy5f7NTcUa5837+ezr/JZ
DzzIkhgQxJ1DElCm5FZluj5AYbBuFX8aq0CPXSFbTqVFnE0HjBL4/D9lZF6on+NZ3BTI3u9IdVIE
kXaNNSgQLovfhjoLElWF7AHw0ow4e4hscr8XCe1zTI4Zwz6C02yAgm6Z8fnufXlwmDwOR6SwaVCS
/7XImtlHLDwtmfcLdBO7/6sCRHv7XQVflr+1eg5WlEz2VV3v+dhTgkDO5gC3ISiSdm93pVs1E8pd
UFlFT4pXK1XtL/hdRKIqrpYWaDARwbLSxGapX7v1QhuLn8JfItAs2JoGLOKyRLM2tYdyrsZE9t3h
zlK3VtCdnBanCZZy6m8cTt2YL0BgNozhQDPx5pgZJXbsODjJNavzffzJnobYOwdyp/Bbz2QVHrH4
PGTUnRSAKo/C/JrRRq83MlGWdKjfySZnasia7HeKGzGKFqKiGxTORodGFDaYp99Y6JKbKB3SuyFN
L+G/qx8yo91wEDcCO7VMAxiR0QX2zHneoaYxEOBYTo7y0F42tLmzdM7tTAW/k9Ca3DG+cEavRMQO
3L8U2oIGxeN5/YAjjltUMNGfiI8+0eF6FG8c0cpCdZo8/BJ2LBa0hJWHgXmL1NkCuaTXyhO+0Y1O
ILQXT7kO1A9pdkoPogDbDhxnSnOTdLVLzGmMHQIHR+w9PFeqIkZ11UPxGs3+eFs1Ezzd8XdMvf+u
6fQst0Qy9seW6qD4yeTKIv3p9dZRaZkkB2Hh9/ZIYAyrNclXGSRtvYARk47tuBM+QWqqXp7g4/IN
1SBGDshatgKV5Rl4QSc91wQfco3udC+n+mBhRAEvKuG6DuR9BSThouifCqkAtFUew0oL27q2ZTol
ggyWAXhXPEWGCDq2G/o948UGLHwGWTFd/r1dzfS6wsGPzlzXnn1sCjBjcVEtRNCOPLSj2yGURHqH
wCnqGjc1NUiE6h83Z4wCb/jJJ/4CEKGJhtEjKye1wshq7TRDYVYO5sZYtDlOOTp8vekFrxV5cSL5
MoxMDDle4b3GxS7cDYUiXnTAQjB8gfCERAQR8xabl13qLmG2hzVGsfBG5t80ZC5ary3RSg7INyTr
GHXEAigdlGzAWMHzd+xH+8331lVg6K9klMpZ78msB8Fif1b1MoVy7F9SdDhAcFNeKbEnrermi7V8
nUa8j6iy0UjJP+oxBaxHGhNytK6p2UiLXlXuYxJTdwf058xC77ibwNI3pNyjZcOqSkgzCqgFHX8P
em5rlvKbN4QV7ki7AVjTdnXCPWzS07r+XCiQS3waEULaqbrAzvHtByPsI3r6WE7Q4WsnR+0xnzt8
23KREKfCtHZmFcHjLdQ8uhyom/sn4JeQuaBiwFosa/9irInrbCWIwUC7qt3wCGAk6f1oesFsjx03
/NOfPXWXYOJ8/DzjI8suSj6hrXF1oocpNOi6rLzZThRnluNXU7Y7KURM5I6uZaYBJR3iQkZNMcQw
fQNxKzsQdiL0xBGKZz5JWHFPTMNZ9MZPjTWjxNGwA2FOMD4/o6whesOkp/KPo9wwgON896NVJN4b
sacVpPpIPmJwSf9Lt644DuHo4tBKxC0vSdwCpkVLSKbGVnCGwJwG/wFk38NGv0/vKJlVQe55WhwZ
5xRM6WKY3wFTa9/SwfeCLsYsHCQJKURjZqWdGJOiBqzvLdcaHQdmmhZq9eFzzTnhdJjG2Zsyh1+R
V+PZpaiis53NnTvgouMwmJOOc7+pcSMVFv5B3gBv4081NVMzPibpMES4hRDreKUofPBMfbY4QIbl
wVnGrAItfKRZmaGb3YPDX1CAVkNOMes8Au5V9Au/tALgTRGh9cM8q7c3ZL7xEbV4U2L/BzJfwn4D
6hf+9ZSWgca1padpWUUw91vKgudDpb8mpNkKgloRa2hXO9+GVflw9TL3RecY2y/aRdh7UkbAebRA
hE02xV4o8PaR+COHglju6HDRl7sxRW/bAQLw58l8DF0Q1nKHUIezIdzyKX550qyBUX0bO7G5fYsL
PGbxJsoGSfZIJrFIB4MJ7A14SuQmHVTXJRx6rcx19VSqiChlLCNOpU95plYIT3SUAMyutU/mA7qA
SWlgZ9d8fgW09cQ+kCvSyyqkueq4Txh6cqq/XlymN7dyXGod4bSgiQ2fnLPE1BPWC8d4vkdN31A4
5IevIDw61mMzIolLePJ/gle0gmOon7YarqpJ9PM6Fn1+YfgIBbgrzS0Dkw9hZWkFxugJmcNnEJCQ
j1uq9py6EHYqH1BOETXfbwAWKuObDbSLE8CWGqi2xbOjBtUqqnUYS7PkJiG1cuU4RUcIY6WHu1F1
HXD7zCr9HC0qfk5EnkM/ludkn/xSLAD5KtP/U9QEbPH6WK5TFIML+F/3jdwxSF7aWau7sHiEzvc/
vBquJFD0R/Qr0+ZMzW2o6yMk55V5oiSjA6+QJsHYCgo42daPcIRi+UaJBVrPkO93JlKe8E0I/R+Z
LtpN19AX3lKoV1WEkfnKZHXUVCC01agcnm7jVn8TOx2ht9Uck0IzgwXk7Nk/DXWcMkDE78uAX2KK
BmZB4H1LV0jBSfI6ORpgcr9V1D5YmW2QZpPA73iHVifk11zLA/QVrs/SH23Et8jM6wGQdGb8dDVD
/tEb+Ket1ZJkpp3+LfZCxlZcwVMCYy1W00eMCuItNheOE+tVezlVmbK8w5wdMlq0Nv5Ub0zcUm70
wIGR4WUwAGm4EnwiHw+pKKGzvoBoeAqfZ1l0hfhg/qLvRVbQtN7ZhPE6j6UV4PHHjqk5o+nnb8Fq
7KBxF005Qt8NbHs8gOboc9BlShO3ycoQwAJwnKKWBNWai0nBeI3pq0E9u5CIGvo1VzSt2QBBpnNN
aosaaT5DFoEbF267CIC/OKICastgIF5QotbCqhWzmAZ6cUVjSIxUirRbINsiYVqB086+Hv3cD6Oi
vY3CQuzQRljrvMDL8eVIDLpd6/bA73+LqbJH0xlnE+uX2PiXyAZzfnyOKJrGalna/sGd6Gj4JPXo
VCVRqbLSFdF4JPsoo2/0sPDKLZXgMl0xlEi9YyDwMnsIcc1mEG1A8Ga9ENmYSIeWi/0fmBAiQ+5O
wgBtOGGnnHEO7NUzpAmh2bSQtL3n7M1Df5vrNOMCcYZfaQ9QkOFQAXKoW0jMDjFWd+CKeUO42ZUX
2hMYrfeWqEA1z7wSymYTuoFAOTeZBa5LDAc9TkhuzdWFPE/KG9dwUM5l/2R1qvhD3bsS8qO/fzkU
6yS12pGDcvuZ+iMnGIkyn4zQhcMRQ7F/VlNOkD5YXzC9qw7w7pmBxEVpLU/vb9GCj0ojhfb6jMpm
MRENbLXmRFP1oTbcGrmftgusu1X6kScYig9u4GJ3r3yBou4Dx5lY5QPl/PjsaFNcEqYHkB2tpbQQ
JBwrnYATHx68DLm7qi1YXyiI6gZnI2sI7aBr3GyLWR303Mm1bIBBXd4lFLXCUGgVK+0KCEG+aij3
JxaEDZ4Trj30AWBHmjGDJpZYSz58rwAsaoACl6whTsdNsB8QlAk9SzOdC6oMuMR+axYeAOBHEAxk
Ds8uQLChp7vFe5qOqNyzL8LZfNsZhnftQ009CLZK5hE626M5CGzh7zvRLJlpU5utEP/ic6riPl7q
k3iCeziX57Ql+Vq9/t6cAAJpmQUSAkEvM/ldwERofnGpusPTUSq0lHgx4J3mjYuDjkksvK0wH6uZ
RWqAuGsQH/OtmwiLL0UoOLwxLpuXANPKBz0n5ROtiAAjSklNvs87ZjE+lRxAeIzBKxtZWHITuaRF
WzprwLdQsNzUBVsmWCpUY3OBwnRNCQ3juV+Xvcdm7Zb8Cp9lcRKMwbgA3rMSZRksbPebyf1wa+8J
MpkaA8cAZYtkbFQPTcMC+5QyPRwN0m3cuTLOwcJyOcMKNoTZRm/KOFtKE5Z7MqFpoumi2as3KPW0
Jcsnb/b3DnDvG4LrP2/B4NFtBXSisnMkfe0UModGqFa/wQvux3aVe+xUmDAfUJD2h2Q6qY/lMH5/
hCgX5CvyISTUkBTHKspmG+2sD6mZ9+4dHsANxcx5qjukJVI5PkaUFobxkYNvjR/VGc0ZSwKzeBEl
K5mW/9y6U1yQT01946yxz1c1pON5N4QmUfD0BnYaJjcxmqAryPlpyVh82/jlTekMfIPj0kiDtUQz
mwfpMGU4e5pDI3/LlBRX9AwwEreDv0crgZoIimGN8qGNIMkI3xYHh3f+0iuSq6ym/JamyQbOYLZF
8jO3k3trYw3GxbXW1BaDKJvJJSlNnlfhmZf2K8mFC/0Xq2b4mLOP8Vbj9LGix/NKNkV6MlAVWja/
JLeSzUP8pvpRghkClKTnpUQBKLiaNhtd8cEPaEqsZJ5FTpduVYC5hSUkWlnYB4Efvgp++BmPv+uY
3YwgYikK33tPyE9IaKwOqivt0ws5L0wIJvzA0goOwomfThy3vKhIa3JgF1kj0YzTvWzoytMyhvSh
CruXGY3061Od+wk0lpNk5X997q8ZqGTq0Dn5FWT99j8JGvNN/14N8nPaIQnfIkfUPL8K1DwCdKNd
OhXQcVfCjhkJUSYutw6jYhcC2UzOnCNdqODXM1DxPaA76RhiorJ0nd2YM3jVYgOYVrzXmStPsQ8E
bZRFlq4VtpySwH4Y7MVj8/Me3Q450HZKvvIP4lQq5XVAogQz4fZfOqE49dyh66hwavLl1GqtR3MZ
bD2dGJMrT8+jkhp61fe95jJsc96RxN0W4ggMQDJL82c7S/i+ZEtREZEeYfsXUgU5UE6lvduciNmK
NFLv9hjOdI7WCdEXYpYtgw8YBHsJQsv04v6D2zvzhz/IJoAB289eVx++9zcmB5AFuZslDCls2EC+
d78SJK7bPKghRStVO6I3tXZ7x67fh2Y+rCpQLnofALSdTYZ0L2X+RHjQRr4A1/aQoOZ8rPQO/zPz
0bR1SDeQiM0ZGh2iTJQ5y4pciDjsA0PdBVyu06l0Mb4AXftrcfh1XiAUvtoOdCr9r/PP4F0iBsIH
kUQR7rV66rApZnfCRFrew70/SVGQtZrRIxyUlOdE/MSsVhw6+/b+Kd5DwtheWSOzlyoPJfOaz/9o
x1SDP04WYR7St1ON9q6LgAMgOXxtCKgc2Cpx8i5vk7qij9vKpJ+UI1SgpmA1RpH/XGDzoHUozjo0
CBM05waQojRYztlCVwIw4wlEoKmchWlabVntR80qhH1r7wcr+RqpqedPP4Baa0rUFxOncLcHKNnk
s5BnbyD0S1fCtvVtjnGd+jHjTfh7leis81FbdWGbeiNGnFwGmoM9mWE8xpSLz7n04HEukCw/xxYj
Oywf4U2KAcIo4QtyaIl5UD5xwcUtPdHZxqOxWN11WiBRj8jlnqYwNu5R16R/yW6rLyOqcK9PIbCS
vh9iZ8evU6kdXjk1bco25elKoO57zIdx+o5EMxvVwkxNh6sUmRabEDlqJiQc/bGDy0DGjFqeeXa1
EKCrjHgZXJGqjvdTZsOEiyzEbWIgdP09Qr52pjZtSmYX1XDKxdsPaz0Mymcj22m76Au8WEc+YlF2
wmGeBJllhop0O2m/rme6i4bci6rJ5TTUNG5Ped2tSOZj3lxuYSSclN83d+XJ/8gJu+ovthxfqx/P
XWwELxhZM3kcSDtj5IE7V8YqIRSylfP9e/4qCaV/Tuzsj3iVZq4Y8PR44Hmykl4k/yGj1gdl5VwB
pcIFi7jFFd2mDW1OpnvGDJLRZqzltPdsyTfGVsXSy3S4WTXPbNp3H4zeqE9JgjC3C1hj7LpPH5UU
ur7KM3WihDSLUmxmFxfZKEIaLWS++cXnpg2HdaGZZ6zpNn8oyVUzys92iiA2+xVsgMEhNW/ASkjF
yTi5BBbO5hAf4D8OJ3yRFWnCefHbYZWues/GVI8Q+eeTR8QvukrQvF4zpW3JcCZKISdpP8i/6ojH
Ayiz11X6kHeEoyfhowhs/d69O7CM8NYjN/TQsg6As7RoiXRWcp4mjwz7e16VBYDOBUXf5sM3vNT/
0m4aD5sZ69dN2rQ9+6WLpQn+F8IV2CdoGUxruHV7yKSBnCnxl0J7PuCgW56zFtoocl5knfnvCZ9K
AE8oUhVcLUQePgsk4xqsAtBTKD5XF5HH6ChggywTb7YKyXyfw1cwBE/uQYga57Kol7o+UTDqviUL
Zef8q5BWnfNSsGJi9G8NeQVJLuHyyYkqV1ym8SiVNlV9310bMCEEz/A1CwKmC6xuZQbccKZ2Y01q
zKXWT20uDomUOFEhL3yrW/nkoF09Wt9JjZmm+EyBvhAhDP6pja7XepRT6AOW5DHu3uPU8tsDNJmm
6erPtsbmpkElK+tOPS658YCJbRcTMG3EMPsAHnYI0qFYUXaciQrR68pOW2h0ic+UTuP0HIbJtmhv
pdO6TU8cCKR1CnsrdfSdo5FMSPLplO2z1KA73XcXxWR68fXxPI4L6X71/6DNjvHr3wytfwV5ndvD
PrLBssisWsq/X2mOPnjQDx8bHb1mOW3fwILdbGN8UBeBxBSVxAEMaO3vzgg1vHauzHVPRHRpIMl3
DohSSbUIaRj9bzGDHyMiS2bHuNvvWyHNyH5Yy4Ceh6lWimFdiPdpgBAJn/VOtUd0ICjyQeqzlORs
fY1i5ZNUmHK+0rPwQhDgtHHSaneYwxEhTtzBiJBNUIC4RVYddvHYJrTYAfVVSsmmhpYiJ1z1DUdQ
OdwVpDo4CrpxmG5jOtVkBSB64+dcw6lBE6woXDrmMfHePTsIbY/ytIGNhfh/QjnxUHhspDOZyRCK
IqKct6wLhqFTI4fMSjRNepSAT4lkM/rVp/9IhOOI8bb1zR/47FvNwssXVAPSLUfAHZ1v1Z/kkrj0
UsOZSPVs6XeCd3frHow4oniMsXxhufGHR5jQm0i9Dgk7kN9hqD6dUNE9HxkULtdkO9rqgTNoc5To
jXMlP9wbhCqRbHr23PEGWeUmzsbrCeXUVMZkq/ZB0fFeS6dgAK19OdGxi1yY5g0FsifVo8bkK6UK
fHQp9FXo75cPfw5fPLUYONegK1wc8IsH1h1ZOuS4lOFekWF4/T14dNLNiXmHQC8mS5eHeVQ2vOGV
MCdKoyL5IV8l9eFqaKclf556mWeOnhNRmv8EfdeIenK+D44dqbhLE3+2YB2dZ2rLh4XQMJpFDicj
KIOdpiF6LExXHxIAjkC2DBn2o4UdByQ8s7bnwDIHisccp2FKNFqxdYuVa6/tnZjr4br7IwOhhioB
XJXtIr66A8mW/v76nFySNWb1kxm+E89NYGHwHc5Jkb4j6BFTUpSsB0CtdboRmqma83ZbDEwjRk4W
0nMpVlS7K6WCwpZ6NfSrflL+uRcsk1oocvjvCrYhwJ++24Iffz7/qba0p2xl/2e7OnuPBKIxiMTt
xF0N2qWgajD+WNoCiGxRGgY5+tVGSBRgRzgdwdn9gPf05q/C0h3ckazMTcJneiPxO2L9PAxhtyIJ
dD3ppZfKiVPMTJSKUOdHh1L0ki+TbIXJ2I8mBhQGZuzF0qfLEyrdVSyC/3R8xGeSAGRk+bILNIqi
FppfnL84tkPrSpU7fkUZ0UxjORnW0fjwtoP66OgrZLYiMtb6hbJa6jy7lGeb6bjiDawB6Ob+7uCG
XrG1ye1EOo0fshfy+zpJ5vYp8KqFr/QyNf4i5cgevB5sI4F6Xmv8cU9928WkW4eWQNyzQLH3qkKQ
qCQQiKkpGuu9XHqVSlnFhzhLUF+hvX8cE5k/TesfxM3k/V0CPbrb0BwZectPpBrOph/dbnwTbc1R
CTTgBEU5oqHL9P2tPMNlZOHpI3BEfM21GPyPpdWR5q+RZDemt5jC9SZ0cFLnkHHnp3Li36d+wIcC
1ZmeVgha2om9RH+Bf4pV/RPWzc1mJHodu1KNSpzCqQsPcAWO1WuYhxqN8MoYHo1gL5Hgs9DkPz6C
aZZmKDJhE9gcAdV8bRzPALQ2IFU8X6uGqi5PP8gB4z/SEgxi1Dri4fP6iOotxu00BWwrzHlpUv9b
Zpeiz2Odq0ukRUfPEkx+VZ+k9IJM1RvwxS1Dl2xQ1kXgUJ3GPAKq5JzH8owJg8YORvqTztsZWAUo
FruK3x/gMP62xtMArmlOKuJpbZJuW2r5mBKo1A5FesFfxRRdcJxNCNq1q3oUbF+27e6LYJfA2OA3
9jvTY9ZFISyAziWK0T1Znp0FDCfRb/ZsLawFrGeA5q4afQ3Lt88zhJkezbxXUMQsEASv09N2CE/0
yczpiSlW3EgUlXRt8cH273oZIGPGYxuepDIwpREicrg0UXwO4i/w1QUTymfixSwHsd6En/Rn/84R
PRNFEUzRdXZ6S9Nf5Q1+Rd1wcrQzaP8122uAM/3XB9rmwVaogVzHyexJvZsMfugP+h8QskDT5LW3
iySnwnZsWVnS6ox2k3D6yGqmWYtslEkutJDSnxyTPyOHXMM2Hr6e35ofnmCk4Db0rKVQ7VjP55fZ
zvPCJ5rQkDKihVYnraXiyjK3ZWd2wu01FnwlYah1KbvNk6GxJs37D/x707nXyjk8s3jGLWSPVQ5t
nUS9LvmR3fZUyjWSoy1UyiMrHcyW7xNiR6eGBNQnFvgbCosCP0zNaMG8ZCQ0/UlfGyrokBkk4Ukl
50mppHzHnC/jRO15vj0AXV+8sXDpI8vqgyosPPKxCvZPm3OTo01A8t+r4966TjN70PXEwbinA3mv
BKAFoXcE7X7/+WjqevqhF4fUqsjXIZLciUuqYwWjOFzeO/fx5Ij7yQBaIihKoKCOeJBrc+uFZRBB
VFRvAs4FZ61RTeeum013GtGMcFCk8vBHUeKMv62eS41yes1SRx+Amy5eGV9Fvh+NnFzZWk1ZIiVh
nu7hLBYe8cuUajKuP0PXq4qQdgHJ3tZUMp+9NBuPNMciFfIwpy2JofssiMTTsmYa4LS5pA2LAv3r
3nipW1yAOm0shOr9OlUsoVGc4GX/4x5vICkLc6QzdVF3MfHZK/m+O2m+jy/mHtbHcLh7j0zxp2uM
Qli+gVZ4PNNDUQ1mR9abkZGfxBmk42RwvRrNF8sF+Ittjw7Err/JlHVsYA1CBjYXt9ic+/+tVYBW
HQICcKjPbscD+eOo/t55K4557avyLlxLf9Pu4Gpw/LXMaZ1DKMHZNN/ugTPZ5KrYApaJCaCMJEG1
UNYKe94Xhysk3i7E2JhBmtXqOHhhwMZLpHhRqAO3yJYPj/COVAl/Abx3030TbiPdE4nEuV9l4pI+
QTXNvpG2PhZrIqTilX58U1L0uYN51svq0LQqmyHboOUQcb85Aj7t+uQtelWlQz4RlStxBNOaLuic
rlzpxnkLUPGiJA0sN45OK0uM8pFJMRlhjIx7yUdeahEVeiautAUymGXrdJ6PMjBINv2fN2amlzx7
uo6qCjIdMYUTRwFtG6ZU1Q6NJXEuKn5/U6WGVTjbbm9KgAZn8wVYP8lFn0Uz4GfjJ2O90k22ev11
eKUTDaHTo9sqMftBZCYSqOzS6+m5xzOblyY0V3gL7g76nG51T26rAo/f0rwqQyhUEoAVC9lsfe7T
R9934oOgJAoUNk8ydwt7+bIipqHS6dLClPX1y81Da4geo4cWoniipEtwaWkmj8ZdBpczw11Q5P9e
pVxbeA5/GvL5u1wnph35kT4uyQXk3M8ICvFDR9Fr/cYpi9AL5nstutkSPFWHtJ0cvq2+ZD3MtCwU
aF0v18n63Q9ve5Fp6O1og8UWK/aVEdbS6EIVWiz1yqePM5AMgUPBh5/xRGCdY3j0KP3VYNctY8Cz
chaogLH7GMa8xHfXPhIvjgw66gthMWDtMNk5PsxMV0lPHqiT3qsqKKZT0k5Q7MI/AxE5JDYX3Ayc
gwiWSFn9Kkj8u49RWiYy+c5jZbW8T1/Q/w/z7efPkobLBucTO68+440oI6Vi0yt3y1w6WlqzwiU/
76sMNqUphFYKD/gfIbPjYGMgXQrTrMgmaSgfMNgCkvPi6FpmiYy1FcrpaERaTs8GwRTnWw0NAhn1
v4CdH8xylOoBteG1P0XLMTY4cxgAYc3LOZOu+DyqekvPZbf6WTiWPmvqfmJS7OMJpLFfekK9I50d
8P42jUx4/ub/8xlwNTp1c8pJgJnjSf2RpU+P2bKE3GOQLNctoThETNZCRcLDtnR5r07eO5mtEI82
hPC2kC2SVtGc9E58I2zSXtwenOchEtzaENVKVql/zkFDd+J6DmGMzrVoxGyD6zfqMKjuJq+DeMKj
RjLAdX3cLOGx9faf6w+12j0/+LW4zoy7y6WvKEYLwusKwks/0e5KnudmcL+35Z+Yfjz7xmfpXbJA
lmVzr24IKXM93fT57tBpEJiqZYDCiOSDEtItExIzUGK7YJ50ARxdpbh6ciByDcMOMnSDYrkQYt7q
3RxftLESup4wbH6RbyJCcexgEUp4ADEU2fcWpOXf7v+nDNpy5UCtY9rAadgbf8wCQGEVLXhP9PuB
aTw7pkWykvOtSJ/DGESvjhMNQEOGFvA/eBUVu3DqlkeL0Mz+cCdL8gNK6Qro2ojT2ncUaGis8dgo
xrIc1CB3SOHUM4uM7I4CpJ3X+D7sV3bAxXXWGSkqDWprCINSJ/tXXw91zXuImydKJi1Pc5xdLcZm
nEaXMphDstyqrjjacSbGyHytjmwKHEHuismXwy+XYOKRlTJ9cMi2dd4bC6mXcQSZo3dm/3G5xm6A
+8f1Y+fWBBpYBi4oZGFPRwnt8OS8HZCT9Pxwla8iko6y1DP3L51oxgxvGMetZjCKVHyvbN3DvCeb
IbSTJVRGNfp8bl4NYOjMO/Z8tSV1di9MfCpqPi7ll2TDZUmmMEsyHgDvSk9Jdks0VU26x2hDEqL3
zxr3DQwPEkySo9zBke6Gq3WWeFhN/Tdbgip1AokkD4ONNOgL56XfxPCDKjFwBPrgTOhueuS/QMzV
d9Qi50EAFK045Dwbz9uJ8QQ+V1MynokEOa7/JHocViFZJoSkAk09aUmfDfC/b1IUnQYE5b7NNUSG
tv5sus5QW784u4ZUEhGZpFa+qExg2s3fjtFeRMA0nHYDUORlKlcO0IEQwvyA8SzT5XlDI0eS/uFy
qounjPgS0d97CRyud5dM1jZ35Q91jxecKjr5bKgGN1EU4lTKnDoDXc/fYQtl0OYNb/lTL5N3O9+8
we9MeE9FwEQFhP74DnCqoAC7zu4DUa1OTGcIHbuqM1vwk8ft3eDJ1POks/q3X9Zqj8qO9uj+KQkg
CR03rxd+o0GmVLarmEjbRwAI89ym/ZLUOemlZcf/kXu0s5G1wZSsmoIU6QyeeiryG/UphhY9crzP
lVuW4gvBfJKu8XCDbTxtKLM3IoXPb/H3lcXnr7zXeK7Qvy9Tx6BcnFKnVdjzI/aK35NQQUcTeUma
nZalJwc7ebcXt6J5aKTipJAqFdGjiIAKALJPxsQXOCkH4EgmSj62GP5UZEsF2/MRazvINq8QEKW6
rhMCW3JTtupXBrpG3ZMgGkGVtL1lIK/Dyc/6b3tlGObgBi7pDimerFOvHX6jJMg19lNABqRgIjPg
TDfCfPMs1RdjvKmLBySUMF7LDKEy76Nz4uWqY0Acr1VJKzuFOAguG0geD6WPBHN02830bF0fKtWt
iIdD/HqVlwlu20oRK0kUXurrZJkuW4QyKnOzUEAroQhQv6ny/rfDyAo02CXAlirsmJsXBoTt5o0k
C7PeMiDSnWk0X1j+nw9Y5IQZpqufOoIjBX1Ylm4r5eAIS9l4AG27YEVHjE+2/RZ0BM2CqcQk44W/
YaRK3PxbzOJY4XGdzYGWs454EDg7I7+m6D2Jy7ctnT1/aXxlKNhr6sPvSgVu2VB3O/GnBUtjCxTj
kl523YtuHTh8y8zFUOGEj5iFtqVM2/BWXGbmaOzJJLbQZyWwmwhe46YjUiHf9ND9qLor7QMbwbFo
a3iUSq0QKqpV+IBkDfrS9ZSjV/j/Ltevf2IYPftEmsmlO66tUrIyB+1ccCK9E+91QdHB+VH//ChX
3W7YIR8wjlfipVIq7tbH7tSaa6ujVrjkCq6ysh3MkG6xmzq+CQBcsctQjzWMnZv4kGLTxhHoncEM
dnXeo3mEFRRBMQNPLFjYjp9oJyCSb3/a4waN3dJSyq+F46lWqEhhJemz/9mKG8Z4/Bofi3n0PgEM
L6tfh9b9U5XiL3SX6MKJvfcfgRc51M+HAif024h3Bt+l5IKXuno1UgxWBDLZxLCYRryOU78dedql
ZlQC7AiFAmOdqO3iWXGfMeLBJwUqqUEfyygvEg0Oh9xHcYunS0yPtC6iQhM3xQMn5EH6CRetpgXH
0gEKvtAe0onxkZHRov5Dky7qLvzre8VQOINAVVFYHGBNHiEDUSXkfkwgsR1Y0kB084WXiLFXjm8W
WVfZMbH99mTAbnuVrxJDvl+GoA2KbEu1TG6sHwaZS9b7iOFcZt3PpXHRh3Tw/lCLHRIZInAYsjDI
1woAoXj7cVjq4LjpC96ZsGiesJ0y/4N0a/TjYw7/J+5X+bEm9Ui3Ow45yWk8e9ga8EWH360NS7TX
qicWAnCxW9olplsStRTeysyXhOZf0rKB5wpHuUyjAFZZpFOx/V+9xoYbNmgKoaPQaDZiuGJkkRTO
Ye517F2HwmAUThuCr8aTjqS+1bEJWVYAHrQdGHZcyGz3XFsPf7w4CCEJ4smPuWPP9/8zvVtzZj0K
CIbJ1jj+Uv+3uE+nOyw/33twKyCpYLxn8lXD+d/pE7GaB+XkH7F2HzlMZ0kQEWD8G/gRTv6q0qG5
IX+aZc0TQuKrQjnClRAEPyJLx2oo3vXHpxvlaQfTR2Ij0VxBOr2V+4DTPTm3vxe+cpqFk/XZWTDd
oUwTtWXFEgYnRD8PIJhMrVTGT6AM8dRnjumrQT/hDEJB7fSD53rsXMAcp/CjQEt3NLCuzeYp6Wy5
r/EEf6vgbR2p+7T9d5NTwnhDzcbMkew3l6v62HdyFvS+dbuZbSYrHfXu/GvSexhDY16zn52a46b6
cBla9DErasgE1sk+YgKiuW4YvUAMXEU6rghmlJDrY2D75gX4NaLRygh8yCILugW9BuSAWkL2hybk
OYUY9gkjPkOTzH7oo+8HnSw0IQaZSARou7X6g1+SLWFWfCeua7gul5DJS3s8ufHBRh9nWvM7cTkJ
nC4EGiEH22SQLB/lf65TmnlJlRs8qeI+8jeAwaQO8y+9uRGnHwoeSxyOPhxmuQxRdYkf33vxRN9o
GzhYFE//89zmDhebT2q5fe3bLaCesLRyNU1KEM7bRvqH0bJcE/0AoR0AuCwZB0jfH3K+5UkwbhzS
MMQzi3FlzaGqKNM/uBX9dn77Mqzw3vH4hvsSS7T4H+vSSUmlhPVevVYlukvvZbdHPk5GJdmPpjMB
I8nGLg7LBeqmqTq/BvOCLsjMbsgOxsXRDhW6CHWBWiWjJxUzYUIMWVHy/D2xZqgwqEr/Z68wKVAt
JN+3Z9gwfHO/4iq/Nwbk7B8TT0BGlHio6uKAcGXuDfAY2SefEbxGaEzyoURhBoOp10yvJbmRM5R8
br+3Sdn3ux+p96eQtJQmgk1Ojof8Z3UQyucNBulZN78ealP3VEK3GVz9T+sU/ehgKKoMBFlo0/PL
0HVFyyRjUJUpmEXQGSdVylNbCKDDguFcnogfLPsNzV4IEhf8YIf8FWjyLd/zsLH9erSo3atJhHiD
hMp+8tOdV0PKfmZKeXXi8h71dsW1qqOiocd4nrqDkj6kRfyBGW3Q6lDr1paOQZjPYzzZIl19Iuke
W4XSHPFox8jgPiywVHHQIIeR/5zFO0eMuL+nqn70f3G34sJZHJM0SYPD0CkeyKrYKKPjORh5aD6S
FqRhxhftK09SZ1iSH0BB3/2maXbJeqsZ5IxU6QyJygBGTBYwef2K5l7XAFtW+YiLvgCWacSYsC3S
BN++bg+5b1J2Nm10UT7F6yRZHkUBFkUZdcPiv0LuFqstFWHgOzAHW5Y5/8v++WwIctLrCWtA8LBk
8oSNG051B7gcPPSplE769qYWvQr4R5u1vqzYe3yesK6a1VoS8ac0ox1UFAGMOlqqVe1DtQJYgCB1
W56FhgZMNTmmMDCfNvJ8xvJmQ5OUqIAWDTdUnKYLysA9IbNiklZy0D7wW94/b5dN1nBblxo5p+PN
8RqO/Gk+h4tK58uyBH0eBMoNLGowwMdxrethZ2ee1chPEdbvd60gOqAdwTI0gvDIjZM/PWvMH42N
T6G1dlRekaZmNl5o5kvT/NuLyfqpdH8jOVpqGzL6gphCk6eyW/LZ28U8Wjc1GugABT43qZmDOXHv
6jc4v8LBVo2NiSFM+Yg22keYE0qh22U3odW1nhmt9aOAKgt3bYsvtDttqg9ORhNB0jlBBjg4qLBC
bvB6Bvqw2g5sMnvnjPxVB7CPxP+xVisxA2uwQanJuWPCWpUP/EWKrmqCjz1Yk5S7bzrlNrKT2JBv
PBM0o73tp32sbF+TgjuMZ+Nrp0ciSPuCjR9324cJZhNtivhjW9HanCFVeBG8P9MD6XXZAq8XOQQh
7uwfB1d9C6lvI+tLTfYgzQFiU/9eS8Rqm7EY3wM2sVCuFf3BvD2r8xUL4s6Yrm//sdjitMyT6Yf8
JvH+MMqV/DzeUapqO86thWIEKSnvUEJxlTTbundUdT/eCe3zatBvQKVaPe2H9YXAgEeKPU9cUIXD
KGukrjLPg6yxMBD2hMKFcCpBna/6cRgJBnQD4rd95b2nOU4Rf5M2+CvccjIQ2dlROY3L0UNG9ch8
h78D3PlyUqA+wcQLEhLujIN5fWOArYZonKS+rQyxbJTz8OzPJZuEHzTt1tuIAdO+jyuGBL2b7GEO
0fSso0GYKB1xL6Xf+/y/Rjmuxj7NqC/fmQhPYnjkkFHIerfkTkCFa3ait6zeL/4rzqa8vZ9bVlzZ
IYHiU9M04N2OdQ5mmgNtD2apKIKBfqQf3SrDgQ2oEOynYB6rVIfG8w2fPAfJ0TTCelYDRDzeKJQj
lTUJ+OXVOWHPz3SI04XRkK8np9fCCtZ1XXOBaX1BLOI2VYSL/oO7mzV2Nb9zc56clQTmIQGTfGbR
JEwmIn8VURbH8k+nmMcGfj5HdhUUl0UwCsqD/x7rpHtaL5DPJCeujF+JodVDaqOh74FetX2vjgXI
oYXgvKg9DpjHCXWow2HZHk5Jo4pkzTg3/FL79Ba28AkoHCQsaUPggGhoyf8md9D0hqsS69mQnZ9t
d+5abkk3IXZOueNBtCfrJjd9bEFZIYxwDjoEGy9x2JTe78JrVyshPD13JEfTI84PR+qZX7/FHKGS
UiqKMQTMU/89BHjirb3+2N4JoQE2uIYkM17u8FVP1tMVBicIquwSCXzuYtLfRqgeTu1kb+8UkMzM
MlE83vF62CC2WnQSwsj7OCFG2XY0vb+EZSZ6ra0mhFBdp5rbVA3mi+JlFF6lJsLbqImJmmIQ8HMI
ekmP48PXUJtAeu7fiRPOtriafGyl24o2QIhmfdrSDHCnOIXIYOREGbO+dgIk6CoU9a7HMoiCXUfW
gzOBztJWIXy1cODqVlhyhjtGmAOSUfAdV4fX5tzA5kUJDHqcAtaanorfR0FDjgQoc3OTKSL2jlQZ
QUmN7Q0D4IQY7Wtu1YflsmGx2KZjpbRJgUFRVp8lwSsnH+xNULMuL6C9N0Wl9gAN6EZzdSGgFzQ3
h5p485GeS8mbVVKCugzsuEjmhAa5NCb0/zq0+czK3MQfkf30hXQhufwaKPccqGrAZuU+NgtAkerF
0x4K0XBC70n3t/E8I6V1nNZR1/OMudiDZrN2dUU3QrfImuwfGRGOo2fd+Xjaq+2cwu6MPq2xpvB9
5aewJ5yUeGsiQjQJ7HQh+Rwi6YZhycDE/ltQPYZHOSwqLZN0bZZtMrMKah+7fnmQ45i10Z81GggQ
Jqq98EMNrlWMPzb3EQyp5KQ0itlW+vYGFKOTmFHpQa90OmZIog7D5l3lO/juNJ69+xGP2wJsivdL
mA97hKGgOQ8VbD+T1Uf0GLXkl5ploiYoYC3JcBI+Z80j+Bm5ossm7UC6a1iB1M5OivHMyKI2ACwd
quMWF/E+xS94LZcWXlrg+mvc//sKrPmg4i0MI4x/B6/eudGBc1jsOkgF5jszJODpgPeRpHSN/mxV
LZG1SppuGlecamLgKdu17vuLjCjr5mZ59U1VoZV6QN+Jy07zh99OU+b4GuKUn8iJAgLKS2/nqmgV
SlfIhl83HOOshepS6dcXTSA7XrVv/KReojdqlf7TKJXqA/Y8xk1vdVsIuqfTx7c6NHOrzXCF+8En
at330KI36RncsaUDr+ic4kI079BzvtKlKdHWcoO6M9rvpjGIDcbEj+mCNZd762IIvT6b6EWal249
jjIoaZtWar+UHOvWFUIBOQH23TvH4xCfIRq2Zwt3sf+eFwej5SCDeZgXrEMYBD4aOnyK7fcN+FVx
kx4hZC+QYAFRIH0rxzcuCCNeysWXkGsCyT24fmmvFfFvTrI3d8hhFjakVFY+isf5GjkZpRIJsr+e
m0PGdHUe40VHgzUjw/oDavzbmfKNL1Sjgt9R6BGOaIbgBgCeLWcpGknsVJVl/mCbamgJRb1QiHDE
+yUPVQuFrijruwdHh0FbPYWSYxT0NrJbWETS3f9fNeyvBK+0hszY5pVYz16CKjpYDgjR/eyAENeR
K9MKqNp0V6tfEaMP5IZfcbiz7g2HstwHXE9UbvrO79U69XSB9Ba7zcaJ/NgkR6NmkFPQsdwi2OGO
cBPVwmZyaJyx7iqwughig8RSp+iwfAZvqHRGn70DGR9LngMrkYWykV0YzvoJrZi/GLQ1a1tGAOmK
gZwMRTfwu2GX0mmsOGO8Nab3XCoTF3mFrjzYjI62hzUph8A70pAZBjWegtDgI6h2nStHRza2IDq8
U0OvkyEOH/8FSYOJ6z3pxV+wJ1FJKfnFVcl4X3Wf1+YgAokHsKKsXZr0Ln5VAZCt7vaycZIrdBCS
LSIVnV9TrhHK2SByciccr9tiNnhCmAYJaZ4vMxT+jKXKMnP1fP7tDgCxL6E8Gu8lLFbGv+nt+y7e
tlKC7qux6/s4dYwR6eimdTo0uxonIzmvruZe+hbSfVMbYfojaBU3uUwPhLOFyEqx7wNpGu5e4+kn
VqDe1vy/TfS/D0aaNK6rSW2542iPGwNP5S5xawftwvsGBkpISuiJObkr17aggoi3FWy57KpXp8dE
WZg6ZTG2L6hW4HLGz9LpFnlUKpyZW/DVD4F37z21PeUS3MafqC8a24lYPEpEFnAPSuCCXXhYoizW
6SQC0CkQBDAKbl8Wi2YUkeI0VahIp2lycmH1kZbTdWDXpsBAgQXPZuSLTGKywP8H9wmGiwyyV3mo
cIJCzMIeS1f6htCJeZ5b/I6BRAc7YlF6hy7i+rdeIzEWCsKulkupdNcknX76yUPksebLCnSitOQ0
kXQVsc3raZnyVCGRJDCsQQGIWDz/SawFsNcHjBnGI129gmyLX5qGsqzcxwQ2E19+Ta/k0sUlOqRj
WjNjGq0w771wERPbibovGkZaAeesHtL0WFDhXwaly9xbp+sgeTYxhfh3ZdT2PMngs2Ei2vhuceIK
q5+K0uqyQDZIzJOTpeDhOoLJf2r++Y1FShjYz5+q22UIm1zdfkYqwxOSA2MxjufeyDQinnGvtBpZ
XfOnKNCJ6URRIlKE+8RmDKx24DOP6ha89orLKWxLS+lwnJipwSO0VpXocwVqGwEH012Isrj6rHWu
ki/TOYBAGRRKTUxfIyI5ufGDc82q7WXtnxw5SS0GgKO/QZQ0W1r6QaB5Cc67E1xkN1zWRRjpJHGQ
+aeKxBGwd5TL1o95OcZ9yZJDT9N9gdhCQU2CkcQ7myPNbNO8S/vynF8EsYxp6GO5vaF9ldNSzqzA
UTIoF8nUuEW+0wTif9PpBw8lyhf07pMqO+3zgthznM+tvGGpXTnVvqFJCz+ISa6LnXWGe8q8WBSY
6kmQ2iaGdQB6v8fHTib3ldWjcQc/0YfIpnTJZLnSYoNgnnS1I3REMZNZYjFrAamYfx5NQrZLlAoR
D44Y5k1HicAo/8YMcVDpLKp1SG+VoQT3CxeLNQz92AwuaUPYArTF8othIrrCX0HwSKQnotNoZH9+
JowVIkM2d0a1uD9BpMGdpuHlT66FRCE057jfTIrjF99U1qLymbSF6RJ2DdiN3QiMdFqBKJ1ttA1i
9zjiB4HPex4NCwWD4ZvnlzLOADwmLNugn2F+uqPXLdzVgUMXYnAgZ6tN1nh2UBdkEkAOmtBHpvCW
oPUl+bSHGB2GaCg3G0els2sidQVyx1Jy52PDnTI9HNjCZDZNh6laljSGLOqISvqJNMPrlg/7dUT1
pH/NJ/NBaG1LY3TE+9f7so5gqYUmu7cD4MPupTtWnmZ8nkVOftFqdmojO8Bq4TFWzpOVWt6SlLTN
mWp9pY+GPvIaavEPgc7I8XxxK5T+KTeHiP+zI5EMEP5BSjcAvYCsFLNa97llmtXuN3G/TNZc9Ulc
QXbRyO2QqdUbeh6DiVCVRq8m8ZtPcdqUSH1PDRbuPtBPMWtfAzN1n5RNKVdJSd/1rBvtGN4dYFS4
B1MkG5LmJGIYsuGWfyIy5nUNFnUwOehueEOMwJsAYUgZ/hGMPEAfnfrB+7FVGuxgSEm2o8pTghiA
Xl7Gs0q0R5NQZYYETGNY16bzDFPSt9WbUJ4fsBq17tGbjOUjnIB2DhDy0ltEhGeBc4B28yjjmtEU
n0jrtXShhi+cpQXE2N0FMH4FAWyHZJXardPGV3+KYl6gfqto9H2ejkgUpLY76vODlKaXHk6oOLfX
VBQw3WnWA2DltmBHrCgVr4kB3XETUcdH3SwWEQ8j1uaI7rjXWaZPT5qb7O17lsCB1cQCv5C0Rvj5
0mXwUXOMrTaNpaAmXlxLX+JhTYsfVek5GAqDvYgslFiVOo7R9RKi+7agEKZhRpfvwTtguDohK5f/
MLDzndmCwQWrRmD87WXKp3nDHN9YVkqzFTh/ebuJvNmpIqcP+ZYje9R+VaRNux3l99AJx66T83TY
7E3UnRnSKgl7GysL3t9USZJ7ALweVR4LVS5tXVFxOgnBuRXKo6ZOoZf59ESoGQA342lS4v8guRSV
DdB3CBKjNd95NfZTqxWCOhLMPMPuGdOhADrN4u14j1rSuHYW9xR/8Bl5N50hk3qwK5GOBZNT2Khl
IvuVy0njL2S8Ee2CzgjcFbRV4k5hQ+sNk9weShlzQ4hYiUCdgXyHaqSoKUxAXW2T6cERP5Pan1bs
EPELEFmHY55cv/Lex5TDgfFO0LNgJZmBc6N5OMgXOCy/UT/H5mc9JWoLTymCNJUybUMu8o9XzrnT
dqhuql5bfLUGzbFBSgMNc1U8lFdv1TVbPsCkE71vE93KrXq2DcjwzpXQMvD9cgqmrkF6TsL9/x1V
B4f2WOdq2PIlC1FToRj62kvN08RSECyi21wF9gXtF5bObvFefcitV8DYmKBxo9imCRQF+j1/A/hT
1Ll/I0chNWIq6Ta9HEa7iaJxYVWurzfA2eC2jbXwTY4I1KyxgHYg0/SUC/SPnOoDm7IHNpd0geGR
0hzNrEMBKeoOWN3HrcY430MuHCtmpgF1eRc5xoVENOcpHcHvWuWdJDJS2R9AJPCzX2L35+KVdhXN
DZcM6c+x3QQqOzFaAbxCO+vPdY3neDFW3VJuven7hY260In5QMVRycUKfGwJGH3NK+lRjBn8odaV
eNXnJ2tesVmOHMdlkBv+BBVCDULLCNvxEph20AdPAW7KFtOQz3/DBZTwwPjVz61+c9MI31t2yWoc
rbLpEXBH+VyBx0YNgt6a7+Kq6e1Zy4kBaB8B0x3PDYpF9GvhM2X54dl0KBZT1AnnrQ7wSWidBz0R
LNF4a8KQXfrw8TNS28U1ySIZ8fKqkO8TEF8MUHJB2mUhPlNVGWCURx4u5QRWdLUo764ZrHgLVA/G
w0gz3i82JIEXbYyfqSIWjPPg1DRWzfCU9cMYXi2f93ffjginQllGi6elRMGCvRageogZWKoRoW5n
YbduE+3+pmgsXlVs2SbcSXUlqsM1ycKjebLV5qerro63w3/FPGICFRwSSF9OwvmYyCv4TRCKMb6S
KleJY1rLeCceUtjY42p/TkgfSerrS1PdT10Gv3ifol7pkitOjJt20gYpnnemv1Fa/b5Yik/8CGYu
Z1dCChqNyKADkoskfkHQGtQOdQ4/MHxcNZdURDfpzA8NVget1nhFzlDeBMqDxcJhquF1F2opakFc
tcgfEOJgXTJTWaCKp1yglDl6J/bT/JAXaIsAKdmejzsPDxwZeXC40YLoZ5z/jA9r7m4ZXTiOxnLX
yPxTQzCSjgugaj5gzWfZtRu6Eu7YFAjDpcbUC37zWjst18iWoMrWX523hjtq+HrSdnp3MLyKuZVs
Bn15tCCYxWQQ0+AGgxPdfes2iF34UisHbqKUMiAZU8v0mL9PS3oRko6ciUGM6CGR7PuO14aR7bEC
BCPiWWrdC4/s66QgYZWbLY6DWJHLQ7fzQC0Z4jmYK9ufeLhzuEG/GrKidHxHbO8VAvKXOqmO+noG
bdHrhJ91X6Bbg5zk6BzzAZgiNVr4Yqy2Ks4SqRPPF0vi8EkxveZaLlwjRpHntevmFlWTr5sB9IzS
IJ/RK/8DQgm3q8z+N55UrXz/MqmsgoCEZvejgKmqC80FCCz5zL4zeVFHBdPg+hM01t/E6rW9NKlg
/gFIfUi0+XfEV5k3ZNpdQUt9CSEVtBsD8i2eKTZly159hNr/Y2iqzRqQnQ66Lxje7dy45scA+QTE
Gn7+wlQzuRtTweBC8fAn0FHuR3bSY4AQqaGI7akBfOWOEgdAQ9Z/viix2u4j7uH+XAHUOmSiDMCY
jL82BopvX0RuYknYd9S60A7GFJfl5CCWTUBP4Fld4olNWllv7n0acuiUjRfblJ7Uj8KP9lpwnThY
XRJNQ8lJlrJncDy0ERAXVo+vcS3WM/1IeftzBpYUZkND6Inteidwx5fAPZCCvIkZaMv2lJuGoK3o
9GF5Dfug5K4R1e+QIUnTV8lZmON+ZT5isIqTWR2cmWS6d5Vywo1o1WQ2FwxXnSEG3+24T4fDTP+L
JgqjnKVbwikmhTBIK6u/6q3VIxTorOe3bTizJzmA/pPfn1ha+NP6nqDk7KQcBGUSOQ2AlvISzG9u
sreJs0GDk4QdXwe27nQwi2+6pZ+5J5endhX+vxgo3peGfHnVFgfGFOaKQf4Lb6CgieKhtxIw86b3
l6deknNGru4WIjVMFAHi+khJd9U888QW/aRVra7lRvARJrQg1VpsO3OKlQzi+iWiaIiV2B6Y5qdE
7Lj6Vb9lpTIJbRiNNhR722q1M9oduVZwjdkIspZT0XdOBik0GM+f2gs86Ah/rxvbUezXvkW3z6b3
7/9t+PX2SDj8M1X0ulcsONIEQwBJWdtGLSOctn+aTLoMlDt+2j9LuUnsn6Q0w9zWMfekaOqrUzEw
ht9gf1LVwsHpF+sqmIBVJAvq1mfliy/WG5Xp3RTmVv+fkJYcDKIv/kMi9F4TVBAfEyXKhps4N8dB
ey7cZBto3KCIbGwnr4PQHfTS30vH5MSTFt9G8oeltdbTt1Wszn2S89DlxPYUJI2WEvSElSlfV3/+
6RMFxPYHAmycaI4MXrVOtz3ROgb6cRfwbiMkwXBozs/U82HqK52FE3xDT5B4J9+A6BhnAOWWirFu
ehqhSKTy6uMWPt6eAb698hST0SImzO9bxmv0yDP0j88fbkIvWUFixQNjdmpksd655WjyFu9cYkqP
WtJx+HdcdxvExg0XjFfYNjhlVJ3MtOBy2euugk92qA4OiIN+lZiFiDa7ER1BfAzsOv4QfnKmcqTX
EIL/ZpvltxB6d1V33AVmqPjs+PZM/lQ9WJ81KWLOTDKr60QX+xTJyO2q19HzSsiC056RIJ64l+cU
Row/W5CF8Kyeptd6jpgCgwWiUbZuAnk3zEIymVTR2pYAv6WPsWaFiV+zBdGg/u58Q9TrJXwvlZqT
UU3b7F5GQMkW568oxtE4UQ6tX1Qn3+nDMcFpaYnHbPpdhpo3qWWz/k9e8zTv6fGy0GbaetLwDEkS
AkxEeMsLKXgz5+Z8mknpjUkVavEc+eJwqBb5YvNsM7X+EB2sPfGKXPiBvSX7pA5tC89HSbrgp/h4
kquVcnVki9HCXUmWOSg5AF40loTblsHZdr+f1OHuAvrhoVNC1cXBEKYdie5xXs3wDm+CjeXw1FsY
ffJ6wejA21MUAzZ2uamiM5J7JAKjAcQeGSbKyUo9gXn2z4ntvO/Ywsli0oFXxJRp+eh0NrPeSSOr
hR9gTm4gZb4f8Umni81ftGCCp/nAmZm5cXF/P5RFPPlgvubUJCEgEw6Uz0+Cy+iZK/H1SGXE5Za6
rjm4jOji4OeTVDjUtpvjEpXmwUxj1JjAspXf47FNLI99BAO2bwHEFwuQq8LIhTWHipfjQ2QGR981
ykDpUZXJPsjnX/VEmrlybHwbO2GvaiFk3GAGRma68zoEO++uCnM6W2v3jCS0wZf7mJKp6pN60gum
HJ/SXrQJwKvCpYqZFdJmje1nkXaNKd4iAahUijRbhorS7JZ2llsUFih4jO+yYh5G6ZtNLFkJIkH2
3aBcXBQAo0Ic4a7/GEa21Vd3P005S9AESZECFP0yTB6ky5/eslHlWxWqeDPbVQ0txcfLS8DURS1H
QFSSXZ3XicVDYS8SmYYCQHtV8OBhF/U1it6o9QPu14jmAm1tybrCNZcS0Klld3NIRGJZ1o7jYro7
HaO4krtVk3xM6UwW2u1zvVTRTpZhzMCqI6jkIyT1HDLdSJbTwkh5f81WmBrZPtZKJI4e5h10bXfC
FFWstqZfxTgbSa/0zN3f5+bI23sgmnjFYVlMN7ABbRIT2jWDbxaHnHz3tEJSxPB9S7IkPrjxIfqR
GDRRaRjOFAI3ycTfD0JR8Q4sFRnPY0Tgei87TlDk7n7YBdNDbiBbfH2UgPx7CxUuizoX065yMREW
uMNfMxoyCo6FVy89KnLsteUiDkLahb7oM/pfqPanAlRRS1Y1yU7ExKL+FpLAWSXAAA7Btz/dnZ8O
6cnWOdma/GFYmGPEL5IYADkASowSyxN8zxCPQZhFZezzGo5HDesmuESaSMr2YX4wA7bdAleKLqYv
ikqqpd0eHUrA2VR5i93390DRmI3HX8ORG/XruSR6VyKNIHyNlKtU6mVsgh7L5kawnOvHSRH3EbX1
gCQkQOYqzvfdThZ7xBUmjvQOUTbN6mLlWHkrIq/rO4BWJqp1PHBWN3XkDKKm3GYRpfe7UyR9KUcr
mevSfRlLDW1lKWn6VKewozrNTIPuFlwQsUDChjzKIQAIy7YZd3IWu30BWDprJWkoOKG9cDSzFE07
eDL9V8CrfEgVtJS3egdN5wbULdDHjv5zVEhri1Ma3dNjh9U18yqWVXFfxzCDIKz78/VL8rXFVW+g
2zAbEpz4ivQEjt5CBhr4BqjLakzAauYjg57PlrhufvEvyp7zyvN7R21xdryRk/Nz+0OcJ+83q7Et
zFeQLge8axNesU3HaZnfl0HOHFTNgkbl1a5fJeZLWEjM2oRlH7AKD5q25ysqwwOHbF4uZ22SSvGy
k0/7wbvlflfolZSvE7eOtTnIRvNH4oXw4RkaMpv9tc8ebk+lWN7UoxRnk8+QfXSz2B/XtUQQY684
Ukh57XWeBzd9z29yv5eZy6ZCc55ZXvOLCs1Coe0AI5ASLaspFBFJ7eZWBUqF6l1aSdPHqfkSbXFf
rEtRnfQRYGP7OXGhfMwKf03taaXYU/EniDp3d15XFak3H6vi4PvxmDwAoTylCf74yTHix8PRw3S9
tWJ+6Tvmj0Zyc35dpwkpsPrKSbz1mAp0+29lyQiGMxbyWVxc/UL76yGiCA5SEzv6c4D1FQQca6eD
+3bvP70ixDVPYvRqYwQm0U8TbGMCMdNNIeymE7SOBQ4dHQRNecUFA8IMqFzSqIQmA2rqnrYwahXP
BKL9VQFkggWDFTAO/VwUQm2zhJYkX55910Jpo2UpbgD4LPyjef8MIKJFvX4fRJl71tqKZoa/cQj1
9q6xGmpckwtBt+k0nrtWTkIIPgYyDSj88lvYsHKzf52B5NOp8N4zfzwLtXcPQ2D/vXoHhVXDqcN1
q7E95rOrqmSHKhwtHnhBTrYAC8e6MvNjnJr+ln8VLYsAL4XU2pA6NZ/F1fceGOrjVhR9KDnSbcwr
XwES6XzrzsdPNUbZxdHSqbV+kqX/xIbPVU1VdMR5VpXLhyooXgVTNqLFUcVB91Hty/HXSRGIivus
aiCI+7oLheItzdLsEOo2n5KAvi9gqOEw0P6rcXdN1Y6Krfa6OQhSE26Plxv3XCeW5RF9CQ6nNh6Y
aFGKC2+FywI8tJ6gOQAwQahmuj8JngugmADsZ3ALSWQu+TmpUg9//Ay8aaM74OnXpRO3azpBTqTr
8QzPVP6TwlM7CAGMHwCYWJCEiJl+xK2KpjHKhu2UMtqJ1wz7HfavCWS9jxm5A0vSXBv5YBLfcrkp
Vjkytlby4RIVz6j2RkjAXj7NSB15+rgspFkBE1AhYQD7GBCfk6DBSwRG3q0LSpvkdeYSNQ9p3UIo
dLXtV5AO0x8Elqufafz5lVb3qDFahQmAiFDekElB8dTv7Hi0FIMorhf6xPBmn9Aw8pXwLlod4gvk
J9lUWkxDi/eC/s0c/u6bI9KL1JhlEh6n6D42yWRUiOurrkMUfb3zH9ITzMFRuVj7JrJRFuA/H0+k
U3P2o6LEytMsVSCkq1hsc7Elp7q03qpV0yHk1LLZciM7nRLm9KwIKCdVXfHsYGqdnB6plzp03L7w
uCchoIr9bCiG6al6HT1WNxeIhrNqGO/iaDcpPHFCbDisKzBoQSJ+Z+9ejivbA4HftgufPuA0dQwg
QGTn9FaoRD6fe5Gic78CDNIL9cH72ZbLXZIQkFfO3+JqC9xMVts+Rl4HOPvVhMGhCt1DnrO9oxTw
6k+Asj5FapFrVnYD5lHH1DDWvK2p28LKKxYxshMMaXhZAD443mOZ/REjcA6blD8Jt+rFQH0CoCCb
29RMPTcYzFSRKdnFs0MdhMmtmxhSKfl6QwAXg0cEqJ5fTq1wBnz323RDhld4gPQSUTkSrQIeOOU4
tQXYiKpEuXN3tTWCd0oCRNm4vJdqyGRi44/PWgANehrVI3ydOg6xxLE6Pqftspc/6SR2qWzzY8ir
HrEQnvQJYqSru8YrYjNWY7ONdPCYRFIYFde0BjKdsW74lFFUPmvceJIBrJkBvpdPc5Ztts+AyjO8
SZlL5NfWt42LWIJXM55f4GAz45pVUFG3iK+0aZEbdiyOnJLSKJJpLGY7AMCKg52SbK4wcCWDnSoX
d/yS0RIIkdf+nRr7LBnzoqJLdfHs7dtqrnJIxPiajqWM7fbmO6WYXxrwgPCeAL/NHpSbWvJws3DD
75/yXC6VR+hyDYuS0ozUpCIZ5LTVBYXBUp011Fak9ni49k0MfJ/3yT+vYRAxmGSgEmH39If3EeK2
ucgQ/oKDPzdMNOaz08VUABB3cimX1mPhhbXKRlFI2N4u+OeX/MxGyX8PzZWPXIsQb1eQkzm15b5e
z4RlpHPk95ujZrTBNBqY+ruskFu9/rhUigeTMpR+38oFal5OZN/GSFPdiG2xcfHwWPKnhaYzqOM8
h0EEw2gK2mawjkhIIZ8/UaIr7/2rQIjXwnKZIz/vGr2d39GwN6NI+3erbJvH0PTKGiqb3ctvTOVo
qVkYOUtfozx59mEmIjk5vuzry//AbveXLUKFAIPFP6o6ejjdhBvhaC9KXFwNR8m+mcFZqqUZLzZZ
YoJ1OX6pbwstevqhZnTx2MCC5Q45/+eQxhXSO2AL5D2S8m2SqzSvgeuu/kaB7NNx1qZXCMQKkKga
ZUONX98Vi+b919faXIOVLBjDQiN8hlzKTnHmaFKywAd5ynw+hchYo6nlaESEpJy4JMwU0/cnkai6
Jw7omnzxK5zwYgER8tDenR1ufbmqZmX0iLel2DByW9c3k962HYfFKQ0dmuVTexqpwbPof6AaSuhP
mr88mNuHYWm/IQvMeQ1hELKbLoWmKSRZKiYWDDJDFs6BftetiawP1JScmUjIUzwdtimCU+DbyZIN
+L80s26xtA5Vw/gcW67c8qddN68wI12y1J7bvrhSD37SDtRFSO2jW36cFX6zwem/8K7jQsAUqX4k
vwL8Citvo6nq/GwbStg7HZfcYLqv4qjWxsLhZlo75okUdvC5hbZ40Mex2NovbtiIKND5tYEF+8F+
5ZuD78mbUrHDOkEwh7Ce3/tzuIMyPtQzvXrEyW+KWqvZnzgMRRC38KL2D7J+GTIRmUo9+fGcyHCJ
Hni5EEzxbeU4PiwsFMBqgnxBFodg5uZ+7R7Q20TIEPllDWaGW3J3llnwQrXXEfIgKxbN5QDkN/x0
OAgHGsQusUbFmLaEzzNQynDp5gmgEIyZRGfymOvbCSdeurrZdKfLfIBgALw14rvDgBqVJL6gHgRo
Q7AGKrUCFXo/IW2pPj3ZnVlM9cqELst39YabNv4OcpnPP2cJVoP5y14lz/rTsdJ5JVt5MirchTJU
9fvO76H/zdYafHdndgIM/NTBNuEka7uatHTi99WQ9mMGa4+ON8Bp9dXVmZsyX+oDHRiO/b1aWLAI
ZjjzZrz3037SDS7H9TerdmBgmAK/CKYiq6+4oYVtjGlGTvr4u9M4F9h+ZnAdzhGOrJT6eUjD0Fsa
wBUxZvXh4OUBhBitbj8zlm8N+YPrUxM+6WrOscEnj1sEejydDcrHFkiDlfZG+QkpKW3XBNFjpcvL
vEcjUdxTEkFZ2K7+aerd7BoeHbxqw5UXyVXBwB2a54oW4u8Z+1V/UwH7j61iweXP9d+lCcQ4EYRK
p+CKBMc26USRAbBBfskO7IbgtYT+fzCEiCi53QhPg7KJwKyKQIi2+xiAioHwOVvf16R8LzUBHjPg
Dhbjk1N260KD4rpQq9Tmb7rB17ix+NhET66NJjV15fP5+cAiSquS+ZzxOJ2FsIzr82B1EVX2SdNX
LtPIczVzDCaSLzVCgCdhOKxIBOwQPVcTmzRJHX3UDQXeud76Uv75WVT2mMXMKljZN83sFYbeTWyp
QxyaUEREn0Usef+UnXxAawiaZcGYT5XXvQmh8p4pjsiQaJUQGqo3hSmhM1Y6mtOM4J288ByoqE1h
6rNDgwSd0/KRu4egJhnxw5IwguDXSP80NbNeYAmu0HFM6UAQZZgt5oln27Eb2SHRNPa7I496jbXZ
pvAwRUeOOgF+npYRbqvBl/mkoSaaV3LI/PAGmds8xSJ2izhbb/Wx7IdlpaOy+vaHGbLZgfh8P0xi
5Azoc/qul5zHwgLXVBgE5nM2LxD/Tmna/gFfp9AoG//aKyXZbpJjTE7iAig0u/MGRs4e7nIQMpRq
XqoagjANf6hYXJ4Y1rTZfayDo57r7dcqfPdE0TjzXw4/Lpcvm97uG6KhiZOxZeu+VKvT/RbmbqZb
lSsPzZN1e3joXxcV5XqzOppzJGls/U1jKAW2DLw1WMEpPeojZV851hrNLe+Bdl7ze7DyGUkqdExR
WlhfW5l3WVe1HW5dTHlrt09gUT9k1SiwKHATRzfypR+1d4sGFxRZy506oKN2zCKaj7mg9P6Lz39V
VrPnlXjnsg12KUVq+YEaqqnt8Wrp7tA2TYpx8UFmTyhCYCjO10Du7dwcCdeIckWR9YmPgAtO9oIh
Qhua/3+q4gm3Q+r5jRIZfSvz7CFEaL5jUKo3/ih1vTiRqbKMEWB6MgsNaDHy++1YUpF1ObzcMIDJ
mZLm0Hmb8WIFYL7gtTkoQjixToiX5+3pRMcuBKHCF9OKFD3gV6zI5WvhY/cCvv0r0CXOH0vzhFkm
J+AC/dIMRmGoG9fu4uFfeFEUg+Udedt+FLmVoFxUc01Xim7m3zXMQuAZ9rbeAMRGPxSdXws7yOMa
GuHo7tmQchHO0tV6qXjckiSe1p/6vtOLh3sLbFGhGPEoLomTHesCNTJoz4dS6pdVj1LGZ65Ee2WS
KUgewAv0lboIicyP7cWKTcCLD80+jFJfmVqzSagFDnKa9+av/nHfc0EgfzyXZixLAMYpSaooKaEQ
cwQX+cxK3lWuQwOYbTZUdN7U/nfgK4Eo2m1tWvlGp05iuKa1dhUY0+w3sJSulTUbrFyKkb2UOHZX
y0f01TGhBnjQ9QXH8AYjqB2D85+zY2gGpgxBV0Rm9z8odOI3Bm0XuVyxVh92ieEZYMUIiBZhlRMy
e8KXJ8iSrzw1JZCKQ3xpr3Ys3npGAt9FK9DrTRoUnKjYqZvZOROLbunkTmKQ7M4gNXKYiEPeMP27
1Ijszz3N8HCVOLbDALrNaPOOdyU3tiF1shvdpzYZKClkqBPXBB1FJ0CKmD6R9AhmtQqadlvuCKyd
HqM/MpeWYG71ydPASykTrXnSPhFPKVS/u/APBbJi9QeQ0yd/MuYUqddQuhCNeWDiiQ68/GWaarny
2dgi8G5F3HIb638aLeeqNQ9KRc6xtkp9Jvb+PPlxpyOMOWMb3ETx6J8sAdO49mad3X02Y3D/AV8z
1vXBHND9bAguUltOrkZvBGeXOuSU7ERf7fObR9PNUFmkyRmi/PbPdg873WuHrrM5XMWSOJJjCNLb
PF+g3eO6zJPibGag/7C3RrHgtiWgvN1DO2hVmH4QwZk+BtP5QgwA6q3eh/iQSmdGtO9lScjvlUw3
OtkBQtArlcFqOcZXylnKYtRrQyFPFMfZ7oy97feYj/kXfJjMlYAArlxq3VpYl7vtOJtKS4L0ZiTk
KhoNCp2bb/FCx5FqQAA4tcyxXot1VRnLgZ2jCyUhPDfg2kNUN0CNuCaINEFcTVOcpCF7/IU61NiA
M1dQC7clAXw/Pk2o+HB6CMzQ9UH6YBg6xJ99n59M3wc6JDkj43/jJmzOkvCX602sbFLZ5Z6ii+Ze
FIFmSAvzDjgHcC5IlZgeylDNwZUWsmOWWE4ZnXWMttkiaktlmJmn2hLMYK+xW+kBCDLMfHJ37rpP
MiUDrcOYZkQDbsLyM2PA/udv588c9Oje/EAWP7Kme9jj4HRSA2qXNJ1eHGorqT66KEbMoqjLQ99E
xqkckxMCRN7IQjYMSfirPOEMAacFPntuucDbPQ2K0izI5RTiEn2JnGVMwa/1x8HPOB70ZttHbPv7
5Nv1gD1unAOU+loIY0t5rDqCPij1TLaLqUNWgdjRztvJHA2dUK0RzQfcCPxYUaU0x8mh2xtDxAVL
p1XG+NcmegrXD+mNwBDpqyqsdEfATF+71TDyX6VltBRfl8h+tkxysoc3N8u/CWlHjzUQOmRPN23b
nOdY9qiQm46v8M1MSIdqyG7NXt6wD++TSSKevuf9ijjtcvmSnaZ0g9CLZTmpBNlcFsLQzb4Q4Ky+
mjOyvYUhUGAZVvQYYYsckyuyjvdsBfYpmHfU8ludgLjLRTvl1mQgvEiNDtgK1DvsoIuavQ8ZGT+l
D6h3Ve0myUJr2v6AjXv3YeNqik+3LfZHzpgC9Mu+CkghbVLobbC8QRh2iP1P2EhwDSKpsDrQNmd4
gauT4ZUGqiVnOLTjF1ajnBSYngHe7SloQfkK7jQ0c9umhYr/++hYlbXsIdgk8tFEgMA8tU8dphN5
HNToMERAgMNaS2MjUo3PXwloju1+GBUaXou/0h7RYokWzSNDSHYdEK607ZlnNw720htWQjn2v941
rp6WIDJYRr+1LigVHu2+MInKhQbCXOxD6KD5refsJ4eDKtHnkX902eLR9ZG/2Bm6oVmTBNqHDTy2
pdxs0i88Fwk8tIUn1O7fZ3Jn4n5EcQggMbAS9luBXr6KxuLL1UlUbD3c0/+f2KE4ks4A/S5G4hSs
e0gguzRYuPuHF5pkyAeZgZaeRwT/CdpDLFdghUliCzZZelYw0h+l7QK7rGoN5MAwvNmDPtRoeTOZ
F/EvMQqI+YU+kTICJCm1YLMm6E9YDyCsic0nmRL5c+b5B4wRK+Liwsi06ahrdLlIfslTBBuzd427
tiHc6L6D5dfs4jl5MEgDm+Xje3yYSSyJqXvDXmbaAkIBWYdIiPm+HZJRzuGyniTgrTxvCDESAdjo
PaymXXCswkaSYBLgGIM8O1wPQNpKgEWzhPCp29yyZC/Dxc5D4AYxsnkj0AXkKQb5iWIlApDdar7C
jjQvhakmDn30QTq3aOiRqbQ8luXMEfX/xXxshJHLHtZQ/NVT7IDD9uOv44AKXNdOC+2PtjxykSbd
pcT7lG/3ENWewa9e6uQvTAGE7s8AbeY8uwA3pKXmIC2hBBP+yfBCpCaP+h5EGXb4cffXBB+Yo9Dx
71Lwsybth/WWodN5eSeMZlFkV5GNwpgK0wKC2XbibfWFAdurle6CvrER/Whj3TFwSwHA5c6SN4oB
jsjxuDxG0rthF2hl8B5RAblWWodQz676JOEOeQHouxrnP42bZgvSyl5OkkafS0oH9PiPkN64+YPq
bYNoeomf/GuLu94nTv0vpiYMsWDzgSBABmY4d6rbmp9I//lCSvOwzPONkHVgPtAH03NEjs77x2TX
Gcs0Vq1QV8h62yGNTsV4/VwWipMDr4gUUFYbkoLn9jzG9D+p7oTPuuNtdvR/pQZEZLxg3GtRAsB1
sGSz43VezwQeHSSpYIwWSSW1H9tOYhPWnH08b4Vn8mpbawZgXA0uu7PzwxE8pIWGURQFElaqEazQ
7ZiX9X1IBlA1x96zPUHcOIrZIS/mFSrGJEkxPlwfHv1WlECCtQjRrLB6es/7kq2Ig7FxKk5SeQsw
X/NG3rOKwu6uVI1o/AZq5llElMxbwdu+XBJqOfUca+Cw+U7ur7CCaLisuuqqH7CsXf1WNzx2V6Xw
wU9M3DVI414m/ktzcIch/yBGkQLARUgZX1hQxk8PVPapMD+cBTtqLEin03z205UTcGHkHQIAagqK
DYmQLI42acO09d7aK+lIIF3jGh6K/dgoMwITMOLrRMThNukweesWceSv2lkXW6TGXZh4IyJeaHjv
ktVBwttNlrTnaTFKQgFfCEtasXB5cdrxIDxiuvIxOeoV4GoQFBBQRJLn1VUKKaivuEPb2wgbA1kF
9pSssefCKrBZQt0wgIiWYrbSLCZM26AtXxi1XUZ8sOkya0ngGrtDoiPFkTpRpxidED3sToKNar0+
cwEzNGeroz7cOXlq8+H/rMoOzDiDUB5dOetRszHlEDoCz6qm9u+hlely5hm+LhdsqQXuZm7AfxO6
hGV1rPmDrPta65mblGjcrs7+MgqtQnU3E0mtR7x3CgzRvyTOoBBjdCgyu6lpqEl6G8JRpg73R7an
ZWLrQfh3GW3uq3KrwglgNIz9GtewOAkNTa+VIzZVVi0nbtaDaf1VHyPRznN6LrDXB2axSCmmF6kG
EMkM6eLZk4qSLGu/KbpyHkvLV1N6NpZz1oJ/kGaMkrOK+NDe1hth0JWPraZDhhWj0rOiOMJ0Cv9K
0/aBji2i9FaE0BIA8NR46NowGvf9ENn16E/3hX4NVwryeOImmdRooRoSq2udBiD4fVZdKK1f2C/z
IOa0S8HL9CZkKU5uJes0Ene5OHgzlbKDUDl6XTONYfV3+DCcji1pQeVg4t5ffUns0RVY4R045SOA
p06+XgA4s40USkFAqAsTrfyO3gq9zKGWQmp6NVM+3hmk64rJ9jgLPZoFBnfftNr9nZ4mdHzS1F0G
7SQ9PxZQMjTO+o9kgR7R4WcMQAATRcOFuLQPr/lrELQnB0eEkic8cBgVi7Ibp3AqULCEYHoMZKSR
Mk3jj9qqmWP78hxEuDZEoj/9e6P6PHaG6+9ejSKNsENWWMFecvsJVzj2MMcwjiIUDNDlc1gv1UIc
v8CiVWh36Havv/m0ZphKIk83qaVCMBHUGDiO7/lFcqrIi7Am1g1sHnHaYkXRxyQ2Zcq2hqFYgHuy
IvZ6O/+4pqBMQNsvdVCoICzWwtVzmnLX/PleiWlIdjQrMCBCwpz6PXqNMEO82VUGki21zBgN6qP2
6bZYt5/776wZzgSmKSxI+oeb01nfSf5GNoOKS0YqCR1oVWCvhSzUixAgt+Qs2v4WD6QCNlOnm1VL
1eSmM+cULNnnSsns9P/ykXSqXgZeR7sAsJzgg6hNDrf6cqg1jXIdCrjwxZHdJI5i7h0q9OD6D8lJ
tvfbLGwjCE5DoA3km80s7T6V2gZCDvh1kiYXAYW9SIZvC5vahBT8ePJfoiYAGNvHOWoa6tjTz9aU
c7yYq+aq3d4tJbfC/83TZZ5rvThE/JeNiYGb86rRfsqPzMeP5S+0IVyFpv2bwsWHOyEtAa9ZRKRZ
IOhA10JkU+kt2ZgwzOZ485QGAH9gV9TI1iZRkOK8xxmPANFnRthwB8z39mv2ysYCzPlOmehqZ/xk
Nr8JNQ73amk9op+m9Z1Y6ClK9fobM+goizALBJDVkpIEvMPbSpe2ltI8g8rVTUrNA8AGRvOWXIYu
wUX58GfHP1+XIXH6XDCTa0U1Rh+OpdB7osWWWokXiYigBYADWQTz6A9XOKKmqQDO3/Cv2SQlDgBx
gMWjgwfDpi/r45ijo4Mb3k2gGi5FfN7aidPXe/jZgPQxPL1fy+QN1s/oVPZLGQnhoQYSDjjRjVAZ
Lhr7CEym0r/NLm7yxH0hGIQPqk1+gfWsK9aGBqh+lJf72ssrG5mp35Nni5u5/NqlfUpnIPS/JHEF
2QimPtysHJT4SDq7f3MQhDgghTRePZFcbtgwCzMo4XYHgm5zqLyyYzkP7mfGUEmAu4ba6l3OHAZ7
YVHXJFSp2ehMwNFUM6/0/tVh4q3bczbeIIflVHb8XPNAQE232kPJjY3XANeCTTbgRkTNstl9uKnf
VDgKQR5V+k5c87YUCivXRXIETAKz/M3z97nZ4EDjZ9PHxcudrnOjeMa5RBv65S0erekziMfdVGQ8
ORmPRSbkQZO0+n9/thQcaGlxzjXkwcMwd1355own5kf8p4aHJSJUewpiqw0Tw56/FJlYUCnwtq83
d9N0aqx1yvwq9AxAbrzLG0PQVTl9PMCDxbedHxnUvOPJp6BP0il8tvZbFFnJ2NnIMr/4e+dE+RxE
0QIQn/X4/2Hlsx9mzKB+mzwsthlG2uB8OkpwVXg4RhZagJzGbb5MszrY3VkpjDPSwo9AEIF2GRRc
eZb4yEgQkaMTmIkiuYouabcyH9ivQi81DteNbha+w28L/iVQkm9zD46NGdXuyjmBmSzQYvcdFTAA
XKpsxWGusO8AXiO5aE5lIVCvSd2nhFQjR3Kt9ZZbYrhhnU/Z8J8XPLBKbm4b9oZaqUj5eMhNw0vn
Zp3XIZTnAARNGEKztpkD5nV3kCtaTGP/sOWwMicMWav9TlSNldZv0KFYmMIeUlMPvT6mNfemjym4
8Z96jzDVdkU2GAfmTE0vJw1YWFZjnlnYWjGx987ejto+gA3AVF5HsTMb8XU07IZl1V6bykvf+Yh8
b8KFHgePRG0vFMFuIRHnYFFz+DqAN367qeCQbOOpOjoehaiVqeWy3vEFmo8wCQ2MNoUxMaOXF6zM
ei3FLsHN/Ce1mLrzK0w8qwca6rOvxJTvW694LHmtZC8hYyecFnZJf4Jbi8X+6vuuoPKJc5lHKFcp
7+LCADbGXFaUsdOmbztUYe1KOFcWbXO1nddWubhac4IEX8j/f/r9POLJsBOdcGNw1GC0o7veQ8KI
x6EvnBJOu6Bt+2h+XxqkmF9JswEuJFojMcLvH9IgHFrxfEhNHScljBSnMyDEXkaXet4mzW1Ni3ye
TbyFYQGwDcGDsyRQ96FMslTASHYTgMNy8GseIimjvfaPxQFvSnyJ9cU60qJg5uPAq9X20YGhQZKj
MCR3VmZHzHfj9F2y84zBAZymrBJciWZOmwAJk+sboqHr9DKQ/82fCXp739eUH0UFG26kDc+kHNq4
PMszpDMQwKup4vSfkbGikHAMZANYcVBEMf8QY1HCOF4KTcJfXtYGLLvywxUIi8XJyxc49nzasfBQ
o2wi3AS3wnFRZM0N/vjmR7BTg/mEt+WxKaoKCYCBgA06z4QyVaxJh5XZB2eG6w1FvWBrw/65teVy
/atN7Xp+lwzhalN9eeL473AHT8uZDQsBmnDB8KBN0ep2GYjFKbY8x13+4MYMXeg/jU029fAC2xJ/
OYw1mvg91ozCqOMky2LFNwjJRa8lqvTKZ19et83LnoV/Se9I4cwEReTiYiEIY9YgmuWWrebSXMGv
xDcCof7c6msSMjFNYIq9m2ygGjBi/XG3lQywdEZf/Kc8Juyg4WSwPNCgi3IjSQdekD8L1wzqdJwN
qlZgHZ+Ol56+3KoJs5Mf3UpDpz5auopKQREe6r8XJl7IqyGmf7a/ImJL/xElCDn/DA4v2HAnF7Ym
1mHvp7cW0Mv6sIcTS++GBNshNf8YOPoHqzkiJP8wS/uV8YSWmzKhIT1EsyqFpJ9qFM3jaN1mVy9X
YFvH2KAd8HJMOjpLWDQRatLjzyRoVKgumaRgxSOIwkxUJr7LYqSgRdfZZIr5NJcd4UdygCTM3uWL
r4PcsR8l/aLrKi06x/Qm/nPtYCsL63XcWJzlrAINd7v4Gkr+5zHGq4SoDOBXRZYDigzWZ+EaE3yT
N7ALmslTb9Y3fyoWaYRXSxOarT1a5ezkR961JCKkbXQOtV09d1Ufj3dgZqscOEhnuYZ10DaYkkW0
MK/Z1GrPSKEFloHN1IUnYkGHpjNKZvw7Ljg71Q0c8Hi8PBNDUzwo0IoMA0mLEMS4y/Pu4aJOo5AQ
8gPLySbeaMppbO5duYID1HqmLo00Y89jjeUAY+j0f8rIgieaP+ORsVci7HM9YkVV0YHuGky0sZ3B
Nb4FmgCONWMz3EjXpg0vPj0hJs1H/c4TaXtuwh0p93Q7O7AK4uGwwPUDzZNoMcpqkONc/1GfSp6R
MUWiJjiLuiCH5LX9jFVWg36ErWe9DWz8omVzEE2cXVf2ZOxbAx0h6cNdXooOqcA9KraBALNlWGJ5
Bd2FFle4eJAKc+LYY4V14cDZvZ1ulpX41vRlLziEBZMmQGb8n2uazTKPjhQzmvocNVu7f7hx165x
2VsruOMpi5JME64P94k5kTgvDlNi1lLDZfHwoURzoEFqCoVze532SQnZQVPzAcgwWKwD9aF16J+f
9xLvy+UnPCWCEbPVp6H0PGci6hCWCpkXHVwNGRzeAdrBLAYEPJ2kGl8xeYdK4tfgYwnXMGb8/mGv
URUYSfbrX8X1d7oeiwb5iQAlmWqMDubchmvg6TKoWKo7HPuvniam/uUdAN+25QfeZZmpJNS6nC/A
15g9c94Ewjflx4nQuGDTRVXHbgISZhVj69T9KpYKcHUgkCX3mL3oRKWfgastd7360f5v2j1GlHs7
6MrR1s1GN9qm2pHtstczC7UJ6Y/ucBlI5KXuNdCdKlnsfK2sBd+r97lZnSThzfNpWhYvhF4M6rI5
KAqGt/neS7g27yoNFjAO5s0/4ank5HgSa0uxH7n/bFmaIyW+RaSA4jNpstgbTiNqh0odW57lNTOX
dtTZ1sAauqa0BEEYkZVMZ1QMsM/VJwYo7YrJfgpHCgvwWQfO2b5snkT1aHw25GoxUgYkFOWvJGm7
g7fRT6hcdgx1Xydj+Gs/fl+4aaMakY0f52yFRUfIkrh5hHihh7tba3KR8kL2Cg6b91N1nvAmME9K
+5esipUEwdvTPeHZkoGtxK/hWmPEKTogqTV+VzNzKSXIMdNOoTMNr3ajR8KMJRSO9CqWtkB+JzNd
u7W9/RuqdMszsTkhH+B1IaKbbUPLUzL9RFpPJ9A6PSPjCPBjZWRPpOfY6yNKkXulkqO58MHwYdcc
Wi1p32z4729ALHfY03P/j25ykQEwUAh56DAQGJvBPBsdXGtZEN0GP8mKGzC0rg89NQJTWj3JW8O+
eJmESUVx0JX1ZnlLAfBQLkhBmw7gTkQ0zDEI44VQfuX6tz/M4wy5W4jCzlov64/80TUZxNityQBz
zZBOwkYLzKVDrmnOL6ehulALPnU+JGfgxd/KYO457Fc/bGPqyFXFZAGf8/ppXCAW8NsyAqgyCOPT
UCn93Fht2hCq3yIThzN+BMDN/9kUTvLxKKwauo7TufMDNKEyhfSlZp7liBj4Kh1r1yqnD9JErQSX
4P5kubFlliATE5KWQgtwJI6D92vXMahH6w4QAZQv6shymxpCwEDyvgbiy4yF8dV+JeP6OS/xDNHj
3smQJF8Jlb/ZYBPfBAnrUUFQmrDApze4ysryisdYlRz6Gngg+LADtlhlVnlchw5RpeYmW/IBEJ0x
8unMuyHO2ii98mYLzcQhewQGGUv4aQI3sy8yODPP2VdER0J+KqkGKL+QDc1mCGo4BGwxzF/U5Kly
MKC6S3ElfvkS7EZMeXYpI14b/CGmYXpCKBGVWJXBzG1KrEoyEYyYfTFBlQBaqbq787HEDDn8LYtj
jGGVKq31xN4pMMo21WbTQj93dzTgyG2gekkI1yawjd5BzxuW9eHSo4lz1ZMIk0b6vIRmhVq74xQR
Wu93ohFcgev6QZ912qec6fS8eN50/ZQS4VkSvvqriLLQTqVuedwUlXpvIuUSJ8E7JGplxEtlDsLr
RLJ4oCgXzQtMR3L6ix8woINnh6qmdS4G6xpPiuRz1YVqa1WtmrQME3Lj86j42+7Cxxj5102TKgtc
a3atkVdxcOmeKVXiy0IDL5KemfWz/JC2T12IpKQePx7aHNxSHScYWMFMD2oa614s9Lc41wi8Xcmw
Ia7YyE85hkr60eYrnZAS2I7G561hy0qSWjNZwZ0bW/GDYCBzXMmR67VGLG3kMExM5gfmQaSf8Skp
rY1M03bue80lDJQi1B0kBJ39lZ9DkHIhI1lO0YoPPOlZhdwGRnJBzRBPkA/TpoQY9mSccBZOKRxo
NR4i/gvFwAHLGOEjyFsWxhB0+GK7+6Yld8Ct0GkLhF+d0JHSLPCnBbMeYqtrm1kuic6nkyKVM/Cu
tzDhkyL/qKcBx+CNxnBCZomehdrSaUBXu+jt7dJWxAsRgIHoHwhgB5ma6+3U5+a1kUV/kkTV05dE
tspG84gVJ8nvFLm+1LrHLQvtrcFqFnm9gjm5l+FF1DtmBmT5EJrFbo+HhcO9USXfLMwPVujA8wkp
qIHq4lAGy3/qA/ZDRQgX6yFRdXw5YHf/j+Ley2LCjs3oRqEmuwquhHxvwIavv2haPmM/Nlpv6Q8Z
Ocw9mM6iwdaYUzr/cNlPEoSFHuE3dTE4h8VsEY2VoPShh9y1F4ARQ4EbgTu4uLJ19pfpDdyDCTYH
LTUpgQNk8/QlUYDM7/G7kyxZDSF4HIeEhHRoqJo3MR35aU5ZgEAcVVnk+YHlinAxrnC4uOjr9Apz
4ooHiSj5WXDjhSF6ofsWDmbFf9uBB4NgxIu1XGrGeJ5lcT8P+HKIEdqVbeMrNnYHXQQuaHD6aDPf
P86iH+FBc1fp790Fz8+ZkafzDSkbvtZsaV49zJswMUgSZcobQYQ/H6RCbHGSkk3tK+k1EaAH7Q8C
NDKyBi9IMVCmup1NX9po4hi0OBLvvm31AmVJvuWOVc6SEsbVVfVIcywLr9/6OtNtyYeLSnlysfLN
bhNgH6g+9O6rfgfAijSXWMRHUJG9ppjoKCz+4pPr5jvHXY1wuK/eiqQO6Sdjo7vZHQ3HUs5gUbhf
woNPJObdiymBx8mqCStUropR3wbEynx/trw/uJGxGdCHWYDDvcD4D7B5KHfijg6mgZAcNxrDd+us
v8Gj2NlPzEWwQOooDcpPvUU14VnjECWORws4frOpep4GkZ0ffmWxTqboZ3HylI9rG5NcpLwa3tDH
tWgatY67oWH8pG137eggobQGJTDpTWJLT++L6sLww8wUkVmABSqFMALHTq5MAiwuTOcim7ADzNhg
3afabhcyeih3V9Kyu6bDVhPsLJNT9qcio3N3PPTMkY8lD/Kjwhpku20tn0nwIq0FWQMIzVygujor
a0S78bzfNajNyNWNAZk6tFbAo47ShqkHCk6oGMpnC1anXTAyWvY5nuTYGy50Jc2VzCqJOAuyeTVR
FSm9WDiWGivJr8Jyu/7SMaNwWdGZvWh3530YEKKHMi1hVZGaDtPUYZMMBxyItMSH3HAybg3YSTjp
PGVx9xCgkiA4e4GEXwf9+QLrVZTdb23bkk/brYVmqOLalIC/RPhgNANZXCk6bdWLi4b7C6/BehUo
cy9yxkOm3ReCesqb5Kq3UIQRuVdweHEGixs33F7P1GenqvJCtns7iNmsh/Gvz8LCWu+T8oRdkJz2
eneE2w7im8mad8uKYOVvgP3pi8d018Q1uwk92J7nLABf5WW1+r0Iq7wn0kIdDkvm+b8nhYt23VNc
k/KyklZxAgq5PaUFR3C9r6/8jDwgS0ibcH7wHkWZE00BrTWCN2KxvuvFGdFVyMgMEfUOvaBVTxJs
HIk6pVdxomYVtWKs1ttm49kqbtPc+cYSJmYsjGOnd0Cyq9m3BLGLNIAeFN4HmM2eqGPV7kzSBsiV
wtmLhA2Ow5BxuO0J6M+lVHFCnGTU51084t421r6CQz7jfrtJPhUynLET2WkaCN2v3Gg2ePYM4JSf
BSAqD+3LfZOwuD29c8FdCUisjzsXOhDUJ6Xy6Ll7F1w7BxQGfDiFdiT5yO9U6NQcWKh4KKv5UAY8
78tV0Q7aRV5OQGDEReQdlB5W9UCQ349Le4OzB50g37uLL1TOiYvRUBdty49oqdH2wYOxaTHMM4LP
LNwXrCi1S1riXxmrqmGAhvLa5cjsHBbqrzhiDbvFeIW5fJn/uMOmGfPlb++KhZsV7X6AlQ9uiFwY
OiJhX0kiF2DkLCNWHbKvXM0Ems1V47a1MsI1Vkgv3cyTOfeuIP/vb4zcCBSBxgzB7Hq/VmiKTDzt
9jeSGko9skfj6CcN0oiunapIYKXP+SxUx/uH9SV9SoqKASoP7qWrY4yMKkp/2hXPCjMh9rt44ynl
87WcoLoVY65O7fLHnoobJj2BZSs0ilRaBnSi2S871cMNHBj/AJhmoyBLWKHuR6MZ/igdl6wq9zL7
QvQ9bpiwyaICv15S159jEOSaBNLZG/t/BINdiag6Gno4KDlDEe/9Z1nFF07DQxt9HKuZD3C24/1G
UXTD2YLprXQBPZ61uAUu5roYbUBZ8dZpNAXW97tBit1bz8rVxmx93N2yeyPCR0xqnlLfQ61GQDic
gVPiHKO/HMokEWJuEPZkzvmXfd8FerEDYvlX40hr8R8SedNNOD1DbeJGz2rhcRpgDyF/shg9zoZe
QVLXrj6QIgNksO62Y2agOgS3FI2e/fB4HCgce7NjvhSeWs91ZsKZnu6zJPZkJK29czfAtu+lEjpF
ZfDX3hoZ/kq+qoNFzoImJhI90MmXD7OnQjY7GxHKm6WA0wtrpC8V6RyQRKO8qg6H5+mDQs25VGZE
4FHfyd34TyTZAVf3WalASs7U7dDmdVgZgQTWzBm6+Zv7kZyh7Kiz1PTA0yj1HblKmELBvOWi4nj9
GPbthP8fHXaeMKRXhzQH3U8ftJ3NsZBRd9rahCBW0bctTGQ2d2qtfMuawvAmcJEEXT45QPicTagw
paZ/Bbwg4IY6xfafqQp4CGKNXjduhw342RMEBWawta12G1LEuUYRYTtZWx/UabIW6toL4BncDNte
oLLq2WraXKYYqBtQfUMjMvbrLG0mahKrwseHPwZMplv7SAIFsBKMtoqJOhNW5QyFCJDXr4sJlfAq
5ExTa9PGrPxncrj0FrCfNxw7UhitMyExTT6bQhWwZR0YXKM3CLTHSB02Ok+UmCaHvjNJkNKgLIdc
HWnckVQl7644SeijAXDGrFPpQDSjeSsO2ruiABl0iIW1XT1KyNQ4xi4a7oZ+FcIF/aBr3G32Vs5x
Cps9tE46f9BGxrdDO38NtJOa1xBWX9DUlc4ERXDAA1uMfNySVErYZXDNoikrxGaHBVLrQRrVmAYh
JJ9mtEz7CpYrDTesJixE1b63EzakwrJYp28mPGRL10Ik2cdPLSWcP83C4eBoy8PqLlobJckcltr6
bZOn2des31J3j3FBwVFjUHou6ll6895d9Vvujy30cwU3n/IVS15HK1v4RMZNZuLLhxyMGA1YHgy5
qEcqb2nK0SsJnNwUZv60X8L0aEe+y6PEGx8tWhtw1i8J5CXyAuxMrYBcZEgb/l8p7p+kHE951l/2
qXz7Nfw/UdxPpqAKEG/W8HtHNCFD2SoWv2bixiX/P/RdQTSfA6rdRwz5WXo/aniG9ur3xHsXfBu4
MSporJ1XLwwQPHnvr1IqRnZ/b89HIvZnDSNaXeb6JPxOycptkvcLGzuVCN6//u1haITy2GA6hZiw
HenhK2rR8hMdlbC6UWtqpRo11F/2cMi7OPZ0s+R4UOB4jp/UnGNCQJajB2sef4Pf6Fyeimo7/irQ
0QXOxNqTuahPI24xsJ9EQ/KvBZTaLZpQNUazpXuugUAusx8U4DdXIb41QLNYbJo5CrRv6V+0BscZ
kgogIFgmrlPwqy9mdFjjaR4N7G/Ri3m+wWaiPdeEL3czXdTmh9lcBAASsg9EquIATM254mZ3wNy6
peu/j1CyEZ2vIZlJb0U1cvzeBx6hjfvwG2uSBKFuUfEiuJpcaJc7LnAJf3aM5AgpvnNBZd5p7mO9
BOykdmcq+WWZcYIlYVEgkmKepkhc6WXEgJgLBrGZmtucXMTYMzrFy4VXsqCAbPcmsG9rDFwYnoNk
P4nRjsAD9wmQwNuzZJ8N8EaLMVrDS88HxFN8gu8t/Z+O2ERRD8Q5u56oaGaXHcCe62DO3dmMDEnj
Bza0VPRqDCH4qJExqZbZaLcLCNgkg97YU+b5m0eKk/ZlJGC1U93XdXXCwr8+EZ20JAfHSU89GaLS
2Zjs5Fg2tAfXfdQieycuLezHIauzlEbNmo1vWtIeriGLK7nFxajbLe0HCIybfofxIhFPiMojpI5H
c8WX9TwqZyIEIHNO30J+FVX6mrlmTXfTcck2gnARnAZ7rBQs7zlv1VKuISjYURgv0sTPXWvWWtCC
kkxmfPCRUHaGkNOvYUdT4J8kkEz0f1hp5r7oFtVfW70C4Y755w750AHPrKgDqKHdconS0SskKiJp
P13X//zuwkn79zfck23UjLKaLgHlIkyWhtQbmMzgvh1CGzUHE9bRcxDzulG1Bl/jJybwNyAFR+dA
BH+1RFh1SEtO7pg/3zWOvhLEHLFItTxcoILZuV2s1Sf0/tVANld6IErQNOrTwu48+4Vuc1r2N1PQ
JIcNAmWpLPCLJ+mJ1q24LcIiYv87mhs7qELUC5Vh3Ugtoy21m/L0Kpu3A4ax4TtQcez0xUhvzRN0
jcQ1kudmcA5SB23ZrTajA/7NDntaCnMxRr38bgc642FN/jNOtd3QwjxmkmXc/NXacL+RahPKOafM
BLoi/44oh7AbGTBHUYYkZHIJyC3XJY85BK1eHoC52Tu4D6F8Nsl+hTtmAuC5lzcbwCBEANL0ytky
7c0RgCmb78/Nr/ujyXB+VtM+nsg4Ugt1ZOZVYU7iTKcgfg4cGAK+AyCLorzABKNjgLhNbynEQIjX
jPMm6yCGOEYXbykN/b68Z4LLxlnIffag7r4gTjYocUe91sZx3/jbVclY9GCY5Gju+tZ1NrVSlQmT
Jhi34RCEK3ygJ4LYKgTiLzWny1ZnGYNIBMoL1k4tTlj0bzFOZDGR1T4aNEeozF0jy6K/2UNxV5gw
rRelm0nuA1MBMIZ8VtK8zJS4JxvgO1U9+/X4h0UUUktRE7t7oPBsvAVYpFbZhE5iwvYi13E9T5oc
+RaIqnbrYSW+iYXT/IOoy4Y16OSUVZ52bzFx50H026Z44YFUMCv/nrZ7hfifhI9IQO07mDjuJiiC
cRXITr6XsrHJ7RSjTZKIyBFLtUxmAK5McKazuD3vXouHwNl5Dv2cvDW57zi/NJLXPlkdpvug5jGN
qcDF3/zNprlRpbjnqENc67stE6MfCfdshPLoKU50M+m3ExZqO1zQyP1V+Pu1QLZfezWP2jGJDTuE
iGJ/xzCE5BHIP2ORYuMgcag2pNd4IjH42Hbh6f8zLFjwGZQ/sb1k/DMm0xJ29aTPYAs5YmWbOKWB
1PcCpT/k/IxSV9wWMOT6kBLfokPa0o+IHrzsMtgSmmuy3EPrTdTXUcYyAbhEGcDOcdeOgZvsVBhS
EP8G7lnLzaKQUs7A7LjF9IMl9vOaL9aZeWmV8+f7wXEeoPQhHbI4kuDRBD+4YZzZC0YgNY1EEyQO
2F4UK9enDoSEtBmI6FNMUtIGNvkPfuF+AJIROLBHjjTfro5shYiUKPQCsPqhgOrEgE6u9G2fymAV
RYJMQtP+nMZAETIf7LoYRrn1Iz4pptQp+BDc57eULch2QuSWQdINEYrbi//vVnjjbzOawktB6/S+
RkaeDhoUplUafh7kf/EehSkNjAW/1NJXv5OOw2JNfPD0/Er5EHPLYDEFuZ0S0yQuKOkjWZNvqTN8
4Iv2rZJX9lmXczSSADKFWQHRWUVtgfelNqLmidqF2J7ETssWp04I/EN1On4Uk7PIN2h9UbNvoTBG
b9NAd/0RUFSdbK7cbDw4lovE4POq/NH13ehZioj7Z5cvIdbKnobfyY1JZJ6ov9bZ9Yi0UGm8z5Nb
plrStZufYG24/rrD0gGDGDLlT0a9zkXPPsE5nmY/5c9h2XhIUj9vSjoS/mmad3PSvZrMQMyj0clj
r3cCO4ypoDkq4cEvDnYiY4huZtjdpuMrUgWsF2025qylX2XQkws4V5NZZHt1QR7TpUiXkAgTd/os
IUqf8YboNYUO4qQaaxKCk6wKmt30PXTpO5IjRSMXwprliYYB38dKPfguc7eQfif2MNLKgywa2bQI
htm+p9wfYIr1CnSgdIk9wKHWZ3zveXQFF0eF94SJhig5iBhaKNjzTTFNRx2dciCk63/OzseD5+GG
mcDtboCdOGPHMDtB0RYJbi4XTOojR7ebriv4mQYGTdRcG7KqRa6PLGfIbKyZZHXqjMp8sNQQmCJy
2IIqr8pO35XL9iFNoGZA5VoKrcVSyaZ6r28F3uAkfBy37byvinwJOwzq9mdaiqd8S+E0UVETDVpQ
4QMoPH+V9fYf0FtIEX1f8/y86xRnCJxab4awtUWEoNblCYHgjZUsKVW+Z0S5DWGMDNzodyKZZvNT
4rZ4gywdkVKkU+GDKlWP48XTKNNom7j7+3EplUzLUNUyu9N5Ifyqf4AbJjuDE2m+TPpzSKCLDLyX
yvAwcPwjnE517noFy7kWBD3jkXip3Zkska+HhnW9dYDdSf1QCL3bNj1mTAuFcKo8XoxxOintgTgs
FwFTMF9U99hRGogjROX/3ahYvoIM2WS+vA7jxoUvu0LiKoZt6A/TxienMbHxurBBN9svmuIdj/2r
5bu4ucDL2rSo4NF87wa/iJ2D1RWjyY6zdNvDOMTNiFrnBQMd7VNy859hdtVLcju7BFCFvsac45F1
rztPfxJg29rZyK7f+Cq0NP3n4tNp40vRNRZm0AICRpQQyo4kFk0f/Zb3XuIP5ZyHbo0CTHysIbLd
ymFqhneP5KaKK9jtv/6FrTHPwtvsI626DFIEPg1CDkEYFy8PdYGe/HADLtcunecVqyu1+Y3RPO3g
ShOvKTvfBB9QyLz36TzPAaT6Al98thmA2NwFCVyaflxwyT9fD8nWWbA2dSepUHxWOYRF+cTloe5W
ClLcjFqWjWUCk4C0sREv+dXRnJYkO9Z8upMZ5tc0HRnCXOcSB+2q+zXZfAYcSbKojpER0LCJVFV6
GixCjkXB5ad/G64FwPPiSSgWUxefI3cXmigBE0bwkuTsLDgus+5bOu2necynwHdulNV5Kw7xurot
8KD9YukCUyOor8n5SuYDI1ej9OyrVc5Zc8axe1Gu9dVx2DUkFHOhCPmX4HqQAcb/oOYa+LQuL+R3
Eaa5E/iVZ6g2Fc3QZizYVmnbPnUwJudII7PFu0TwXezdGPk3okEberSjsGxRBoB6ayWOxB+l8N9a
dpYMb9lnwSXw/WxJAzPtDJ/AOxbZNaRKCNVqGq3LgZ2KRTSbYnJH9R4x9LG1l5JNCxmSLH4CGEog
whUkvw3pvLQ+AP9c5nVBCsArB0F3uIStrEHqnRl++Y5iBfEwSm4iHS/vMdp5LuMDQsoa4jhJYKfP
6MiTlrR/Q3uxQViFVlOCHVplN/YsgmQw9PfQRNBp/e6sPJ4S124d5eZWsxx00x+HjjP3BOHiKrLW
FyvzmLoCLrM6ZCV44fK6xaTPPVOATM3PbR2xYU42SvlV1FXjoWdbQeyI6qzZy+SnG33uQhX4yirC
+nfzkdg3spsYtUtXCc8vH9zAY/1g8BZMTAcQUKluOrr7iuxFB/iPUD2aR6dBDlXzk9NHHBNOSAuE
HMgE3CnYXTGMVq9G+Bf1077Kp5vqjX5YkcBiz3wKRRfhOg19Hv1xFp45twhJInSoV2aC+w0WUoY1
sjXseU6vbqluHkkXIhSdMyDa8qWU1LY8jjrxJAq3+mjilsp/6A/dJN5VYQcDzLKaEhll2fgIpiim
qsL63zfi72NvtpBLG4chK33VBBGW+aGJMZjg15XRzX2yyhdPLBJ9O2E7eFxAfmHpYJsv89Ei0GTN
LAa/nuEqUE/UioY22QDPuIQaUgYjcHi9QCfq7qJPxnHHdtiZ3M1vladWfhUTYrcJyLfgj9rIDlA1
UMHwTb9aFEIZuTsEMFyFwZ9JKa4Yg2HkwqZUZM+FMSKltiCW1Jzldc2+umU4Np+KtLzlI3JKyv4g
Z6ZAPJ+FJYks9Qr9UfcjlfdAzsXnm2Hgitx2rwuU2KcFwn7AcFAlx7/1dCHzZjATaNzLltUwGRdQ
/rdxdW92ue6kev8tQoqqOjKubgXNzk3Xtb5v22u+nS6VsiksXanVtyivwtle6akACfBneJyTkXof
nMvuytVpi2bUA6DA5L0kDKh9ithWxiFhmp3Ou45NKKFlI5FJt7+c3zvMyKA2X9gWzoFCgbIUMbLJ
oX8kmYrpvcRvUQ8dYXWZ6poGIYeTwL23kCEWVX46nPbukxpng+jlU+fnS6PWidYQP8ATx1wBwv+R
ffix1KTxmDtmJuzCfXw+188YlFfOzwKJYuaDD2wYtAKHzqgtUfbSnOorBc63Le+N+e2W3PP6ING5
tntjd23vOV53Avh5HIp9Tiu0PnJKLg35cUPHXFuEgXUucpl02VIF7K4q6nmzUccRFHQ4F8vtfIY+
dvIa3dnV2VIPXuSPyrSrSIBuNT6f4ktL1AadAUQQ+7si5qbMhz5DO8NjuaCmPGrayVqqznLnBWrS
Mlea/2DecA8RPKtgif+p35Wo1zojyTVAH7VGE0BasdCkzrg5Nj/iDZP+3LV21++wxQmLWViuFjIu
E/F8uAFwp1NdL5T1eFF7+2X6PnvvFiFSWWnD9oSo1vcIBUUiwgOQ5YUQ/Ow/mygjnEeU/j//7vob
rfvb3UB0Q4yV5L+l15+8tWp7MRbRpazy/GGsFo6QF9YKGR8aQYXhWrnKWuMO5ijSC+e3LdJ+3HZv
hEzxEHSR+qg/I7zQzjM4zgWq44glQWRlf2Sb5EMomC/i8hzR1xNpfrfOekCDdrYL66Cd9F5L/eot
2pEz8es0gNhR+2ibJkXpspsFzy6V9RilqUhKpoKWqC0iNjvVkj9SkYnB7/KX0X3GI8Tp7L0rj0Ro
5Y7LBDFkaQVhQI9K6cvpo3L1zyD+55xUBt758CK0OP8uXnye887sjtlufBtkrDs3GtaPUMpkeQj5
rD73nAr0BP6Q1WWxZ41ViwPT7XLXQpTOy9c2wqsu2eaY8gaTOP9zcvmW5GWfx9JEsWnJGyUhZO+L
k2NWSH601qFfOHOD7Pvn//ovGVlxfNRm4GXPi87rA5d5xeqpdlFXSpmDD5YHexXaFPL47LIQb9px
6vWq3LICUATubcqtGsqy7vnEhZI93jPcpjIiaTETCLDEtmmLVsCxeLpEVVVW7vRQzbKY/CfUtPoG
UZjHjLzO187s2/s09L6u0PQNtLJToiu10+HXAYLkrYA1aH9zZg6qqdcnr7EQplYLqX9Uf8fqI/qF
qHp7L/tCyXsQIl+yjme8TDSLG0zL20C7+2lc8TaGYJ1ScI9Kr3WljiUQ7sBr4XuYzNHQKy+pQhXe
QGajvb/RQE593c73ZhNhBMg24CRRLw10T4UmtWsNm1NPGU52nTli0i2WSoQT6x2rHZMoNCJD51K8
SYwUvRsRyRA8n8mvkgahsye/LkjzqLwm25RptM+m2S11k1XskaTnEx+cikjt5SY8NJMnAhsI4ryI
KosN2mofQOQDN/JeyE6K4awSivywonrq71ZS3PVX0JOTGEWBrp4kyX+8d9XhbzbqQ+DrZRSiw64M
IRzzcA79HxqGjELC9mAEpmg9RuprSyjhn+H7NhDbKEnU0LiJG0hV6nt+DXKFYGsUGDFYxduvo2q1
ZhnLxxYTaKkL4HgCtibCAWo+zNzqzgSbMKnotK9dqNFard4lsNEl/Mvm2LREh1U0+Nb5sb1WWch4
myWe+jL1HyYLY82nSJ+2vCCRvocwbpOudojgdqNBymkQho7KQP7dBv+jw3/XzMpmo5X/WfJ2odDw
8MLKPvtnlxfGN2t88HwyujDMI9QsjExkH7wSTnSq5ApdJPkvStr1YF7hoCfG6g8CuQeAA29treim
FMr4NETT1oCfpUcm/KtvCaUT2lv0fIIJQkBR8JNbo447hRjZw/li9hxrte3mA5D16J+J0UMgH/2z
WOnTTbm/QVrZPe0lBDMN769J/puGoHCrd+VaSIIwEAgnEG3f5x9we3haNwZYzr037Owv8W0AZxry
1IJJRz3LulbclavhsdPWc8N3FQNZuLHJexKzv7Xv6KM8h0Y4KreION0ACVpu7uRyLJ2yEJ5Tue5w
buRxIvyYLqLbIsJGtQgmE/TmOHYiph965rUNf7iTmoJ/wznfOYKDqajWZdZdQjfjWlS64HfDFafu
5eqeYlLSnNoF/H7Q5HiQwpYcNpV7l5BYsE9UOenDg9EzUtuyy1UMKMJVhLYx+nXolT/Pq3auSiaw
cDAHcSmKDED5t6QoDS95VU+qmNnRMuPL6XaTE9RI0CPiFhMTjp4TOndZ/pY7SmVCv2H1nFbksYXT
ytkW1kiIn0fXMygJ4qVONgG3hQ5gPBfmZzrsrK05IwnBY+8AQ/+z+ikqx+YCMyksASADcMJtzMzq
Lpo7DJP9ddQ4nREjTpD6eQgEBv2LhLr1GXcxF59Ja3yPrOdGCvnqOT4ZWOIfv7N6tHiQ+K31/zR7
3FOn5MzmPN7Kr6AOpVd+/64wGLnUDLVNrMBswgcbaL/qD6OhU2DtlvylfJAnZs1xdzJJX5k9Lu4f
DNbrmJetNPDQqGfJboDbAAFcRrzLrRMPpd7iYIaLFeFx2H63HsDvUwSE+H9c7yHeIulEiS9TVqYA
xbbyFeXsdd8YQGJH+NOhiq/xvVsBgzXkVXAPlVCkEO0bEA4EfNKXUrMNeabT+oG5shqu842ZN3Um
WXxntTNyDG4a+jGdQBRAtRDUscFCfLWVCuwvA+xUdb/HMhpsif7D/hF9tkmCK5ekiBcKZn654wyT
LkD7JCDSFm50C0GQtPu4f1YJpCtsml2OoTvpBMs+g1rBDbRlnLkQcNoWJbcMQ6DMfeXEG9WuZ+Nu
vh+MqjmDsuvsnOsVZ1xzXnuNmPuAYRCJ6GrgFWFDqjGD7Sr/CxcW8R8pLJPOBgCLKXCCbe4CEGJT
pSMrPb33MIAidJdlg0glPOh17Jw7FBiwifLkSnjcxq/lLdqIMPxJ9onC1lm//x5R4X0by2YXDZF/
c09rnhUD7a7eiitLjXXeWtlaTESFlHVhatLldapD7bIfPoFTyqpeSuy30XWRZ120lYx8oy/EGHF2
wigAZEdLtlrNzxd+r8ddvFXS2pLLf7tmtr9H4BkQnT3E4/QcSAXvmW7p19K9I4u7OlUwn/soCRBu
HyU8cCdaB490G8eQwxmEkyBkFNw+QuOGTtxhQd1jK0ywfxgdEgjCCxonrV0vr+fPAEqw8k+2ix4+
RLCKssXUYyPmnh7uzPJq12859Rb2gbzGdPW2KmMj4d3xcfJLkRLS+nA6vTpdvBolVj2Q6RpW49H+
Wrq2+FpSbLK+dyUL0IodPJKeYsgJQ+JTvOVjDIFNUfEQ57CNtOSs/sBbCsF2ZJC5DcYjy1czk+2P
bQRv0MCYmJlIJqzIs1vW+1yke8NpPwTWfuwWkcHW5YjYvoF3sJISP0YAqoc/tfO5FZyCpayoVdFZ
rRUJPRI/KWLWGaJ/OrY3Gh4rplEXM03TERcLJ1gzW2Bd1Z6KoqoVa4xm4YKde/4KK4Yiu6vUS2S9
2lrP8AltSsMnozHQUhEf64HCdau00Lb428ybCSHulr+IBtBAPuBYWiTCFYYxlNXrPfQPzUbYcng5
ECqBOKJPdBD84BpfSgXFlTLi/qwMSoJfMTLqx4yxiZIkjmeiARadlV5mq0yWTmofyxHhoLIB6W7g
pbm90m9WvSo5Ipa8c/c20a+M58fST6Q9KTDjrt3Id7I3KqQlOSlLs0Pg4LkMa7ia/J6yc0cH8gWm
NiHAMMfKaKtpOx97Jtqzkgho9r3dTCIVo55EC2ro7vf3fUkvGrJaa3v/Jf7AHsK6beXo+S6I6nSi
HLcCE609nViiJ9+L+LXK6sb+y0ZntuogdT13Zf0dlyPdM6G+aqr4AfJJ4CcdRlcXgZitpRs9+tP+
GrkJdmPwkzVZ9oA6X7Co+l/ZGYGOhBqJOrCWUVjcd9+SU8YFPAfhOGXGui/ECfsnoGrv7CNExo8g
QpiXsIR0hLEBPu6G5KQy8+PO30J+aqGlgBlWDm1ya75O4RSiViDhLfrz/HTvT/fxKQhqVhPOPwvN
Toaq7itQLUSDg8pOIX50VzZE1d5nojmaZLqfQ/InbHzk2SiYOq8pOOr9+5jFSAfVCuM8DxC2SWIy
lJL/ZbaXt3WLT407Gjvi9YSIxL3ZmfVRDvpzOO5xNj0e1SGhdbPHvA2RUxN9cbGYwThtNzE7WP1q
jtgPixziL4PebVbR6UaGprs03Nmb7UqqUbQi3X7/AsGAnjoTL7olT2c6JUTfb9MkOXYflyezfP1P
pvrIDYH1RSWERieVC08vB3UE5KQZFNeYGu2vrA7bFL4CJ/HturR0aqUqU8BsdsuUqF8pZ8Mx+jOD
Bh2MdWrWXtLuWpVoU7BQzbM213D1/uESefCaWaDR14pCUgeKja8qnycnGE6kxYPsHLL77Ya9K7eo
vLkhSReW5Xtytktb65WZax+9ORiPD2S0+bSAOoJot8AksYX2Z+KsdAedjUR6UW+7KRYKGbi2ZQgn
mJBPmzDHJCjL/mC11w5kiC6D4e/yQKr+WgDgcpEhTJAUNMv4Y3u07OeGPEanKuxWp0ultpSsO9Qh
BUqNzQX8tZsDTWjcKaByxAL5V6if/oYhYZhypifB2EL6jcA2m6WZciXUDeRLjU/yKsDMUFEO0toV
s5kVEzXVOXD1GPcmOTApKO0w3uB+XsS0YSn9dIPe/6iEIc+wminKqDPHuC2TvgJkewAKEvAgZ40K
yWOnzkcHfWWAu0jV40vAJ0Fjk3pHBSn3w+qfIUvtvCaYPdVcCAd7jlrn5P5yz/8YuFPU4dmpy2MX
aMsda0LruYd1WuvBLw/uvDXjEGYb6zgWn8vNeuX2alubuNoxuYfLVm0qnCRYMflTN6aRHCrb584e
jIczwfGtJzUk06DwmlDD8CHlaynafF/lzzIHoSJzz2LKYyiUeLdPzipvKKyy10BLimccazTy6VG/
7A8iGHAdxki0mBLOR3gvXkz/SyXEcwvYAKKZo/5xL6VBpVbApMxd+DHKmQJ1ehC+u79wJp2J3BnS
1PmwWDXrpMUdTYkUQbHDY9BTa1cp6cl2ocF7K97QlitRdiC4vijcpcYX1igUVfs4lTKBHIEPfyf4
8oOJfF3x3OOpROLsus9kfLwHdVymv12DGwD8CVTehlNmIVP3UQnxdk9Tchpe7jq651yWObj7a7rw
lG6pNameYs2ojNCGrgOElvqdOfDHwK/xwi1I+Xr608Mj9zJDMbeh14YVVU8f2QT/X6WGEMP+b0xm
w12igSZ0rNEAqo9X4X3w3q9LU8McIy6rDn2kHOAGjRey2Eb268F9pZ2LiPSWi87sygXQxuIw5Vuy
CbUuD0G6n12OmKtNvmG5CADzrDfbl9L/rcCE7ach5M3t9Hw96Tv30b3nyjIend7Yx6tBytZvN8SP
biW+0XSB1JbnxzPXXdONa1IIhx9Yy2kBsKYbzUg+9zubPoYOJ4MWaxuXIY64P3a0PKaAJi2ohlDI
F2O13WFbGSRrpmU26fm/EfBCB+VRYnkU+AeLYSMlxL1mEtAfwNDXprysTUPNqJCu8DobbZMokczq
lg5Eou5CLwyLVmzoQUQO+tFaMkaPV0qsFyOANS51YJAV6WQLXSbroj4IPgWPF61CkvFRO1cXeuyi
jSDV/zrv1dKX+qrnZFucmj5XzWX+us7B3WkK9Q/qKwgnp74in5dulcbv2E/lh1fIA+lf5y+dPVup
cxZ+LgrTmYsO2eJQKgbS4uGGTnbWR9j4iJGDz/jVdZ2wwvDCuzYvoVD6Q8L3QftOlJ73uKNtX+JF
/QbYGNTLVKO2hdB6/Vw1kykLlSjuy5h1vI9ojMJsGJu78kM26ACCFEtnn5NIgK5vAVLayYZ5cEDI
uSwDizV4UNf4+vHiFOsk8zh0pZFhkODOwWslYlUrHN4SROJWgb7MtnGg+3yLMRVYu/h+J1EbhR5I
9bzdlSHPLaJjYt83hlE2z084JxSzkfXbm6YKw/y0xhnz66ivyGFFPcJx3Wf4CBtd9Rw7ktYLAz6t
IAp7GiGEto1qeGO/qmyLjmwlcPWKC4PMfmOEK6hATdMVB/FlJYwOelQP3Cv1Y0zxPM6V4JZhzGlv
O0qjZAq0HWRb9UtcgOmY8FkqIOHb7DALkbcQRjr6Wyg0EA3J+vZK4KAMMuzSPsX/No+ojfeOGOIJ
O33YYmQ+duutk0kEp7z1rwymZsdYJitYZsJAM0626z7wpYrlwlykcWsMldQw8TlE31n1Ny+1hqqN
7Saor9BJQB54K3xSkrVj/qs+Gg0A5dT0EvHCySXwxLPokRqzjy2ZJhMo6AzYCtHyL+JWTsgxm30D
YguoCQ5lHSD8WA5UyCw2fT9BKbjMGtQNGxdoE8E8yt0sRgOhKCLus8TAwnL28f9B2AJxj7YYrc8a
j21H2HhmQJt1IpvXw/idxMVjyX43ZKGU1APezgcGABHe0e8FSyYGE31w2JyYjLAGWGv/Ix2YSoxe
ES9eBkwhWZkfMkIAeeqCR56xQBOGxD9GnxahAf7x/HkcHs3Z2ZEG6EnwZT+4INjeBGWXYBbVpr+X
ezNV3nubEpAjUdLOnR2n5k6rpj4xYLv+hVHWDd0okXv0FvcrnD2DxgoGauSCBRuus7WbOfEDL/IB
Atf/Y9qJQc6PE6/zMf+NLK8vjpvH/brFKK99B6NmUjSrFFgkA5UkjqUOf6UQz4DOmDmqcSlVGhSl
yItNCGikME5utj9Tn4La5ggTRfy6UkGbqSXGHEQs7E2e043jdIJLpuC9Se6+3jUrQ8+4U4UIBZ15
0mVhphRjJZkOz7ChPgBeAhBoCdKm7/MLOaSfnJkE3k8Q13Y1wOumXIwiVyBO7+SQ8vZmp+V3KETz
sHdNtGSeuLGC0p5vWyoUxB12vYCsIcSEQu87rQUqbYS2zDXtgQdp9Kqu66xCucs9jocRi8GmJkaJ
fUlfCvfjjdsUkvMBMeauQd2XFjZ7vOV/i1rOS/aS8OZLZjLd9KD+zd9dotgWsajYMRKkFpogQh68
tQzHW7qhaTP56+fL/apbqE71LxLyh+bMCYWWuJpR0TabUgnl3w1p6go9fCjN2PheHjHv2PeYIttj
PlFbHc4yB9dZQnCzG/YYIwgHTQg4TrpRHKfKiUVaRncQkBwRGP9e74WkuETeTiRvg4xarNSlIffe
i2KzoTK+7ABomH1VKDodfA3JOop2nxPGOQLikBdUJZapKJNvEathFEqbMkOlvqdPW4YjCFBZ7IEj
BR3Sl2PDOcI5b55SdA5NI92ztio+QP7uRO4swOCFVlKVHYsjl6nkl64nFTaXu7OLWnOX7W6FkxPu
bhlszHMy+ybxazLgHzZwq8uxNeguAi3AVjnbPrmHqzThxqx3w0j+7zWL+DOO+ztPAn6jmC+5BxwZ
zeC1fVXzJRbb5fIsDR6RYg7OQhcj5+NeBdPUwDsIT8ABSllHqhCA+zWHoRVSv2bDI0PnZJJPfdRa
AKBtm2u33Zccy9LdCBN8LIG41735hpOW8JhIyDeoY4rU19eWpTYGg3+0X9JIJSLkUyGFZOMD4hG5
vzQbm1PkVkjUGC0bZ1NmE911yiQGK9nKMFaIKPvvNGQxVKWTTJ6y5qBnApOOyLTG5wVlNmFeRmwJ
fgOra0EiDifTTMashiyE0cORjfQ0qjKjPwypIIWpE1Lar3W8jQa1ut0NGdTxYfilOULu7r1zCQIE
M0Hq2yII/MAwjpSWluWZ9snTh9WtyTFoJiMY21QAFva3p6vVB4AVE4T3Za+dh1azaOZH/q5zAAp2
9RZSU5CoE6A25INTm9/b0nB9pgoCH+zJ9fpVwN9hP0VHkLewEbVVJGipj/6yqh28nr/wN5OzzRnO
t/2Tf4wEVY29YpieyFPhozgtDilq2F+zSggyVR9GDTTp/KrcRmvU95Djxw8wtN3tyr1G2UXBK13B
dOkqTPbUhWTqsLuyHALsx7SaHQ3A+tuixcEI8EKNQAq6oyTrxfZPDJ6NYfr6p1qAiQUFUdeQ+C5a
L1gGAj6w8lcoKfZtPvf3SDHsoY7hU2987j0A3F+RnlxaS0xF2tKH4ColFGH6ZyH1UFMyW5jndTqv
RNTtQnjr7ushM9wpb2+nbYprB0pw7g0mzjrReD1E27gB+9M57HqpdjKYa34jAHalxAMTiUiFGvSV
/bwxGqMZpfk6XNpqOL1P+ps2dRrYIvXLivZlRJcuBm1CFmA4uC8ZvSAtn5iiztDeHs/oFV0YqFY4
ydj7bAMBah5gH9xqVFw3PXCf/VQagK9UtjOt/qWZq4DvOiNtOr0Ae5iZ0GuPnmXLNzG6mOvwQ7dg
AAXaNYqR73V0YWJeV3iSfMaUufg6ksP7gVzNwWYRckmhK0LpzmKDxCTPrFxWGQQ4BQye2nJjxBXC
hwLM4NnwIiYcUAO7FX7dMCnKtcXT9hBgWOugJHNDiSwuj8K5qhP/q85bhS4L3sTWim6dm/qxs7yr
rwkbCvCLqGQo0X9rH5afdhNJFB1yJfFoKJ3KYYWSBc3/rK4+ZtQuO2wgovkbbLCEqcy56vld/1Ks
osjY6gxeuz8otUwINyE7gkP6qZKFCTNImKm5J2V9FqtiW5UrGRGqP4XBlBujxglkQFBKeVoeczPJ
6YUH58MiHBZBOPhuXgByUF8HqixT5TcFRO9eNynXVlg3jAiFKcpHu9rNCD6UHrsc07a424M5nnbE
6QxVlKNipNhCiYtFmV+V8nm4dE+k11Rc+CyA2/Q9xlhdzil5H6hBMkFJLYO+HuLpXCl2DI5xsF9s
bqDtAPdocEQtPG1slqhtX/NiOlzHHVPR+HuyTVG4KAJWhvhyIl6X/sO8+CxixWBz9pc2LTxvLa6K
1nCRSqF8TRro0wYPvFSVy86+mbjjPLSAyTGbX7aP7j3OE1z9YvOGAmdnKRPytoYCFUDjqtXfQM0B
KJpQqtH4dMI4JFkaEGNo8hqscUxydd3Y85+HH+d0tnZg2+ThaDR91wosyYYyTe51xe++YuhiKXUr
LK9BYFuMOJJnD2hhzJWWS1vffJxsNRH2p06uO7IrqL3Q4QyTI+oQ5Z0UlRpAgDU4/vn13swV2Yfm
KqNNmSJudecMyNNdvyfPnnhZ0r9Gj8OPUd0XUxMxTV0m+5+YnObqffZImv9kTORkdpV4e8fnITlP
qkKprahEjxvmqwdZWVBNBjwVWGVDktlZW+mKhQTzUty3ICAQ2LTN26T7dH0yICBPwJt3Te06RBYC
TMhO5AR+Vylh05tOioyLA7WQLLw21BLpLkyV2bx47JNOhE6Ai/SjlfJZHFvVXjmZ53YdmDNXOjUf
cf21gfxFTEwUk48LE0ARGQUBETsV7QZPTIrMNGwNxL87yJRNAWSOh4SLTa0taCNQk3KYQxwwlnlZ
GbYr/cI7396niMhoiK0zs0kKhKPO+uo+VnFjwuoI/7U8dU5Tg8u/gjvCdxb16kpEJ+nwSzN1c5KN
uCZGiQR9VEUiikeJ2ji0U7xaC+AkZrVyC4DlYDDLlC7tTquC9BtmUIobAStoKmD1ZeG7At4x2CVQ
/e+UHIEoI09khrBdicAy5J3H8wSabz+++dXvnsJB592Q14lVLM3y+DfpCn8q7iBLgA+XFSy2jS9g
77mpFMhq3uqco2/iXLqy1IZ/gYPDL+vIQC16IHsf8cAU/1I4d9U4H+k5bWAuO8F4ehXkef2UKADJ
RhYIlpIy6gzJx4EyZKf4kveBsVgXYHTBZ61J2ammG9Nlx6FNVsNUZRc2dGWFe8nxMNinwcNgDX/z
U/6XgzJbdaVeZgGM4KGzqj3tCYzUIz8sMfi6cGZvyhm1kV1qm6IKJnhutDMkmVkj2WZYKQrTfYkn
dBEyaxkb86NOxtA1HVpuVTESkhfQVEYr4jgzydZ1B10eaQ1Fj5TahbIJY3fBiCp3Peh7kNCne2JS
iA9OvXreSY4bXCX2eDHXhWvzDKBUo+rSxU1Fakuk2YPGzMNblvcw6Jt/P2ZqYomn0foaMvZehkWL
/qreLgP+bNPN3Vh5Wg9F7LK7gRTPV0MkoWiG4ZbxxcdxkwPIcZmSyVjfVHAb9fFNM7Uc083MAGuA
+bvDRMOH5kYroR7D7vOukbJNRIefJ/0X6wlPYCsVMjLRRZi5Ule4RTDSC14tW0JC/Gs9mJeelYNc
73evi0BQqsV0OfuqYOuRuPoeoKUolDjuQm6wV6H9EZ9YC2QIQfW1hh555I5FnKMbdbiyui2F3z+C
nEqjRVRi1/iVcYUiKOJYbhJv/2Y7WE0Fb73sWF5ZZL6L1hHNtdU+RE0CfXPEYZRroWYpIeQBvLam
PiOMd8ZLotr94dnb7as+sZPLdh2bcGjNtVJCCQHF4hl1LL7ktm6FtwhsQ76aXI93u9LcWDAKO2ub
1Wev9MgDXmTkmsWRHwTarEe/9mAY0i1VQBHmO2QXFbB8Vg7wH6sR00PwrWxuTsJc9ckIpV2tolfw
a/uCZBXPLGucAHdwvE6kV5xqpWloVZEYT0BWj0TntCSDQf+OoWwzJsKpKaHnVWWal5zNePpBLtBm
Kr0kEvH1pE2Kp5y3IFnb3g3zP3cB8kOAI+dhW44p3U0Sm+7Qfdt9shSpaBEMSJ8mPoFd5eZnndIc
j7t9eSwsIjCseFnw0kIPmvSLOdA8kbCZfqpcpPK93gJJqEsLabXC3QByopyaoPa/kmzoiGcIMkda
yg6k0CHdJpMlaywvRm3Uo899GYGFlR80hIoNsEjH9vw6SB2+mXp+NwsHrAZMXt+qjV0dSfAig6wM
oijzWbuq8IWOukTDY8Rawr38jqmjkApny+3/ZnziLgBpJk9wiBMqomXuOHW05kVOsTeaZRTGCMGc
rDUJmlMOUOT4RYx5APB4fG0fSrOQkYI8Jb4Inrkd5ZXuKSvZ9l3yk+WPjff5L0QYitcq+hDyUayE
f4F1YKrOv7nzF5cZvd9gK/cqbsHd8OSc6PzQf6hZ24ZshkbkAtoYpzMLpVzAN0DTIPvMV8Y8e9Ne
VFf6vgmTmFfjW9onuBnPfrWh2MhTdjfkUGb9PfiklzFNGuKOaY2qUIoqOPw5xVZMaGwdjvOJCOJ+
rS5r84xE4svDhRtFrn9pw3IOghBQRoN2+N/LsFj2H8zikkge18o5CYTqv+EhGWIcnsr3wZIwGyDW
H4Pv7UIyCW5JuDXISAVJh/HbKUpt0ypu7orwRKIugU/GquDwgXwX3lHYbJWdD+1/+peZmRD9Td9L
F5QSwXvNAEoUvtcZ0TQqF0xw86GuqJvIMlf4+bqJGSUy5KF3h0TxvSD1CuwUH40DBT5puknwZKTh
F/8A4BhV0yr/JJGxl6JZudgzXOZ3sCHOP7Bl2OolRtxMk9zf70c220iDRtdK+3YqeZ0iK54qs86V
vLdN12qM8IqoIHmR4papTSFRChVMKgUwUNFioCF7gBbru3GD8zvcpihV8v9//2BnXTnhA2gnSadB
bz4+cCw5bqsykuSmYs5f/L8tIebNCzPPwCnDDrTYAZigrdFLw6+SUxBNbsKRug10rYVpE/8SCxPK
zrVXpnOluh8sv2qbxbiaod4A78Wo7fp53lHkZiJVSY9ynDzh4lAvCY8Ai2LZV2WcaDttuL/Nom/B
kHdODlx7tIdNRpOjMPAVZ8dHTEWIdZqVIclwfqK0KpaHwAN3AWBa1fgYU3YwPmR+YSrfrK9pvPys
SZfjUxp1aIlwEc3BChq6MmCWhVLtlVh9fq7xUrpDAEAXRwtFbot/jg4JO22F9tUrkUCf8ro/MpZ5
tSJKpG1Og+hQojc/uw4xTWMjOrpDeuhi9d8lCOx8Z8SNmSkzsDkc4Y8Y4kVDyUoLBGkWId0NYy+s
XtcoYsDYI5rDzqTTc5Y/udWSbU1gBDY3Fr5vw06z5zWOjpndbbDu6FviN7yD7hfNnK8JGkwqNxar
fPEXu8v1mezuvLxbLya+O0VxAi9V0j8gy+D0jHxBCFOuzikuDXa0rHGuKoGei8pGPc/sTFJFiSO2
tqTQs01E0ULQkM8pB80NkwJ2yLw9va/qvB9udMF5fa5XPgb/F5p7eTVkMujuE8dCWxS1Rnls1HB/
0bvjF+HhQNP02ZMupnvUyhza4fny27AktduwwPqliKDVBmkczaqwJ/v/1uhoDxlJCQx+43g7+iPB
aeiRPJzhgsqG7Gw8fTjyIyEcxbBkRZt6qHAO30bD6RkfeTLMVw2K9Z7ZLmoFuNQYZIZAhBRkAZIU
B4D+Bt4X+IQ6Il7VWuLLC+ZRWETsigm45cirGBx1ExQKY0j5RPrq7wBQhq867VyP8D11sZnMg6P2
AcrmY0xd1B3uHwR35k27O4lfdaweUwIocqMNmf5iX3wLBUe+lIB1vdO12h/PtfYN0RY0SJOdHvih
LarZxnEQIuIc4A/s0cc7jAT6ZznunIHb81eKr6n6bNzIawg7o2BVmmx944HGxCsYM7zK+pC6exed
Xfq28Valg1wgaIwLJ/STcLx+L+knLU+WW/bqDm6DB605TcNs3DHNZ10NeaQLeaNC1HNYMni1zUe4
9qm6weJSm/bD/9PkrvBk1P5vt3XVHXySm7DTw5lACJIzmYlu2nLs46fY+LGYcMmK+5x9ct1JsLbh
QBcA3fm8gtvhauT16mquQo3GwYNVoz31HqeNUHpcL+HKK/vy/4CKJhDIAj5FYxfFe2hHzxzNByIr
w6x4aOPW4wBg5cp3q0LYDnujCktJHi4KlHAWw7gVwt5O4Agnr5JlEmNF2uWoV8fOleAmIHuYI8DB
+wafxLKkdwPj31sJsepu383BjyE1tmIUItgpVuyXGayyGJX6zmgq7301JeVjbQ3xIMWqiRmPYy0X
zyxlXi+yyihPE/cX2vNMeao4VAo2oz/Mjlz5e5z2xuhOCz0tmObeiAVFQEKzgrz1+hEWXHrpXZtz
IRnxuZzg84+kAFnXUFCeyMHODtc5baWhq8TaYtc26Iky8ZrQxzAbj3cnPd1p+B7Vl4Sa5IcW9LFc
AGzmwHMRkrgiC+OUt2wJPWrIjB/ekMzNh/P+Ly3qnsqXIViqJp7GYXvnf8oXv2qTbRkBYpZgw/KV
wNgrR5pIE2X2oNYNZ/i0P2erE5jMrqUWjE7bOUw9b8T5JhNEqHtsSVtygkwQ3WCUi4MiIjmj57AZ
d50rc/m86AlFmx+DfGw2NVcZ5zEIAd3GUdW2dtpollJKudvBDBR3cWmirnkPJYGjO11SGhMAjWzQ
GoTOZNT8LOhRhjKTZzesBQo+5F1gDrwsKo6DVUv5r9UEk9RzQBLfSSng+l2+X02xOhJwtH/TgEpS
/iAuFOGuABWCeVV/+uMhjKmMhY/I4mUmZ5gxmYDeX/e7e7VyWJqYt4zgRPSVMqeNnMSTgWSXoolP
Rg7KinFRok4MLo1ruHkaO0EwEFazbi3YDPiwruunA9FPRfFN4SZ3UYMtS3yLhs5JS4YrG/N0xDN6
5qMpC5TAbWwO/sflkLjxdAOjwOr7CwGKsn6AQtWf1Vw7BTGPTh853IJfD3EBSqJEm0C2wGireFHZ
jM0xHJvRgFAOM03qbaN6ydFQ9AtArQkbmdaj1HEl/kid+B//J9Kt+X24K0qb6BzUuGFtPCBEmksB
/1AKjDV45/HHbHl1PoOpSP73JYxBKC0ubf4fa7VRIQWYB328uRS8OhbiPdUpAYuEHLF6pZb+UFlf
qGnMymVJT9qhGtzeoECPQySkuDv2SaIuaYmZ1n32cBj2MUDM3iiWtvwvV0un1tU/csOgd0PWxEIn
WGrO9g48Ug+O7UW3JDDekb5Y0k6cOBVFgH33kBW+Y0xtBHe23okE/W4+CTYrC69LOA5wM5iBkDxw
o1kjY9z/kGEMqU1tT7eL7yLfy1cXpFLBo6dNL9osHgvHC4IHcaMrXF/iclukraubTw0lZf4qzLse
+HRzqUz81/m+CxQI7rKhRohEjPYXlVaNdf15VUwteYfrKlQ7BQTuGunq9oXKhFnKRjtDLTo4SuZI
su30lBbueuEVfEtNpEDPS4fCHe+d33DwOJwsLaQT03P8oH95DxD5sgXcNqN6CLxtEls+xzPaKfqi
IRsM6bOrIRwLeTJH/l7kDFqONgXscYExRY7aJmDDZ6ejyMUBJ3E/TrOqqw6SR8zC1ellTMgii12T
FwlIW4iCwVj0qqopA98qhhix+MMhguxDx8/Tfc7CSRHe1lAFPQkGPaztm+tuUhWxiOlMoLn65X/T
qVmRGAH3ckuYgAlYDGZaZzal40KRhlEJEzNeYD6IZ/SZ01nQuHsgt45ug2D67Nw1qKs3HV6qxKjT
rL7O9eGQ6G1h3xQiNcraDtZjs1kKyHMN09fE2RA6qfGFQtxYttj4ZG3fVqxetfTqfOE6FhT39coZ
iTro/qGEEqt05Wl+FJh9RWpPg4A7eXb7Ea69mhgmoEQpOo2KuSkMrDLYZaDI94CLtmbVofot3CMV
Mt/ICUDZkIXDQfQMg1eRqLG4K9YbBUb73yFvZ5nOXK1jDOsUUgxLIBF6tZwv0/y6frSy7EXSmdis
pQO7HtR0lEglul08bHzI5HGJ5MM7Gfqw/oT/QbJRUGA0m3SH4j2m3lyiKD2pefxsRIwlbY0nL0i9
+xzY21gnbxK4CDePKb4oGiw11bPBoPO/r8OoFPqhtaf38RH+6ezC1yDdbffcBmMOgNVQ6BXQwIFP
ArcC6yR3iCh6NGAWhC8pyMgXezD95Mim622lYxUSZG93v2qQM0bXoeg4CMMCMgzumAbusXAaE7wr
VMKx2IsPtfnG3jyQ4T2DpWTlUS2bh+5LoMTfZTSunU1+MadKxINdKFxvQ7RI89OMe/1o5u+KYo/n
4/XVJrpJjGY3X8349ivQyNRTa/2R8aVgjSyzxeMpjyJFBYbE6IKLwiw3K3y4eTNoavJiwf/TDCLh
Wh+nD6lpjx3FrZsBrvyln8LRHRoYM12tYQxmMpylgcTKwjAZycU5aK9UUATt/zioWvJ36b3h7bZN
7k3X0qK0YoEEGoe4mju9TDor4uPeYxUPzsvHZ9Y0eIvXF7579Daavb55ypCQl/v+r0TvMgWZAJhj
auHFhY0zloMrgk3AvHXOTMvqx8p2LG6VCQBWXk6U0hi22MGmya6YvbCdd5WhO0JsPxT/PKpAKV37
/wjhgIC9n67Z/X4JAMpKljNd00QUvG2oWFs4LRJjzOc6DbPlrvkBWBQ+n3aRRM0XS1W+JbEKovKp
/6upDlRsSzlHOV9n8HOktnrL480zzKz3eYmNy7azEX1NhzJGXVJRafqhpbkoo/P6SIzr/kCWpveS
3K8CIdexRjht4bh8Vs+nqEgjF33+EololLhmHxbB26vK2cTVgi3+2n3H84HYi0p/cAo6/nblL+HX
wPo+ePh8O3u2R4VzwZ/l871+6Z7x8q4ZxO9r2rRi4K0FDm+yXk7MbWexk6H4weliKUky8T1kgMSy
EgXd4sVHa6xmRXSTiSf09Sb7Csx/AAX26ha/Z5yJbdA60qJvwHc2PXsuQnWl+CUbUBf0QC55uSHR
kDRfGUHsw0CRzkO+FkzEZN7tUIKUOZ39bPuABGB9IOVuN6Dh1zIA5O6ikGS+NaPyuTPw1V/TaZQd
2i1gvIW9iL/QsMNuCPfrcdH0rKma7smX/fgdW8DbnO4jvTbdf6zCBSw0O/kU18DfjUvqZlR9Rqmz
OF9nmGPdhYc7Ork1JicVBcNGvR8nzPYH3PefcpduUTMUITUxM5f49S9ECdxrPhIzjtNIgGotaN+j
RUpo7K0MHQZoAX/JT+xhdYe+WI3ximRtRYIXK5rLu3XQii2pd0nsodrmnu46zhNb5L/V4Rhcrkke
7VFY+plVPn5afUyok+z+IfzIhWvObAEdYmfA9n/kxDU98SC2epccVm9kM/FwcC0IZoAsvQC3XO4L
4J4iXvnN6r6Ds2zBO8I62p2TpWWmJvw2xv1nHWgl1uC4z8gl8ZUiTzsuCbqxQu2izgM7EWuE99s0
n4fe7wHAUyTpIjLvsPIqoUpzbkBRYNXp+LNG2O1zq5Zf8jAjqSkryecHEUOe/bAprq7+WkvYQKxX
tu447Jv1aH8ZXwYcIo/EOa5TDpFjdfAipSjwLfup+qQ1ZvP7c6LoqhtzVoQko6bonA96uChamkyd
LRyvP5dbuE6if1TQpez+ysHUj9E7s0K0D9CSTB/55Tye0JFVFUFp6BDsGRf43q2OxXDNx+1E2IHJ
9+uGJsMKFkV+0kC5Zh7DgBdyXu49IYu2uGopiKzknIOCZ3tLWVvLXf6qwkqzn1Xyt9k97z+ZYgWk
l1CvMEeX+aNB74X4gTG/nlgqznyntoPlP7+V9TRwwNwUpljiVFrYaAxB+F7pNbzZDW6Ssfw6a4gp
nKvO33n+usiDkKo17aLreaFuBM0VAlCK+RaCg1irOhWPY1Eb2q9meOysAYZZ5IJ2jH8ymhWinmfb
N5USBqile3KXxY8r2UiENYBHoOvmz3v7vbKdEtH0SfUirbOFcIZeAMMeBv5BXRh4LnYY0I5bt+4D
cxhMUv1hVj/qINaWk7THIl4Hjp4DlsaoSBLXuzUp78PcFyI5JYREhxB+pK3ttefOitHZf4V8F5EF
b1zwp6GBng9Wqd8kBbr4/PbTihKNO8M6Uqh77SjEzVrCXA7qrnnKnu6hJUJ0NHBGbkxQYAwLxFAj
s4i24W1IqWj2SHnon1qF47o9NRAdoOcYDYRSmhW6QJC8YXa3+g8okjtyICJyRtC9l05IgZVElDTJ
rLP2I8GGihCE9SwTZSw000kn8qhuIRCQ4GXhY8EhpWi9jNdwEfdh0ExMnaCXDORQ/UlHNivSrQcP
Tc8nC/QEsRj05hmftGypnuHyl78NnYQ/Q1JnlZW5wMEFtOTXBaOr0ukcudgH0oeDCVl/KhVgOOQS
UfFRPSnprgCEok6Dt5k39bVYcIA8OazmLcRyoUQyCa52YScATxGWLJ5raNusL1Et4fOw7mrUxM+s
O+wY5Nr9tU7BgHVqy5ichvq/p17vffrvOP1Qa8+oFn/fafpdqarfPnE4Pde4oufbJDIhFRTdLKWQ
rZNuPswW40DKIZFn8tN1/A+U+dMvDAoDa/EGZ6lu4m6njsKmMah9gUtrmkkicY1bWcJugG8DCVeA
5kSZBZtq2i8/sr5FavGcw9fSb7BHqsgu2zZnZSTNa8wa9qW6zeEQfRSkzXAAI3+dZ5Dl+cajBDAS
Wi9HcIOD7xDuMBQCxwj1/zxe4JFplojMKRtFHm9VWHsDR9bmvoVLFPW/KpmYWQuK68GZDAxh9WRI
3PF2iegS9fiIhx5OefjAxTL8lYzLpBp+KMYjFp3J0JX0l+N9PuvnzIjakY7BFKfVcmkF4NN5SZn/
eqjVjIuWQIMDqksDZdLaPJs8TPjdKQv/leBXgLROwd/hJlhHgbz+Zoj8XY5u+lmw80qZJAseYI9P
K0HXp0C28gA40AmkBkWZW2bfsqVxKBsUcdvBE20RMe83jgxh/ZvqXidPE0AGyCPzrAmldaD3hw6c
JszAnOzGu1T3LWwbmNzaKr1WMu/XepPmILeQjGnMVL43aDodvofSPY1lc0EleoIzeaRG83UWGGTL
fFkr9/nguQdkI82aeP15x54N29e6MfQmBegzN6NvFUpXVZfYBD/ub1ovb8KJFU0mocH3SztljABR
9+ySgdggTuL0s7YGohWjZNe/dX7IasotHwE05R9yi6v+PClS+HM1hFmtKCc+m42F7L8nm5DLlB0g
x/ssTgH1KnFDEiFXlnoXQfCOquzbRKgcmulqmIAlZmNERWVnoCiGJmDQNp3FslW3dSutemKLI1FZ
05u+E8hmWTDDOMq1Aok0cXWcLX1pFfz2Fq19a5w2EFj30+mknEkabHZPbMG1YsKe5849wIy6So+o
H6qI1irkkPv5oHC8mQLiQSbwuvK037DFz6yKVlKC+Yk1pGFfSB1QIZ+BCGTAtsb4t8167HfNT0sT
9Y6Klu86dru3bM+5lYWu9fQyOC4/19BPWjZkOQIT5S1Cmw33SJzhTQYu++ITw86OIQL1xb4BZapE
gfxuqYIIPaX4y7XVR2dM1xr8lgivpwhW0PjkDoUoDI+nWnivYWZFL5qJb8wJgzJD39d3ZruGOzlE
QOnOihFXOR5a+BX8KASZZwu53zLfZmhz4D5+B4cl/XKej9l5HGuu4LkF3x4+dSIADh1DsYV1fGAC
1QCJ1OJkpEOTkXUuNmd94CrXnSpRbAaxcAxj6ssxFD3AlNQN4aLZ95cAPdaNnmaqVH00gTWOSmAo
FuWGQejwIRw3QzhrlYLbgHNiqQ27gUsaieFpFyT1y3gHLqQjLHmUC8H0l/7ee+jb+734aldZvBsJ
Sa0bQGqjrpvLYbHM4UoMBBGRgLVaFZ4dsB7rO0MVT/qXMSUTG051Br8zW9k1E9PfIWVjW9GqyIWR
PoHUCHrn6rqT3aE8u9hPnOmGzTw1yyYIhuilxjepY5x4nMhjrK0/XA79kP4/aYSd6QlmXphi82sZ
vjRWM6GC8HhJ14+J9xExxE+8WHk6ioy3Owp+qrrHGXSajMrDHlR6xe/5Q8eiEEVes287sxUIrkzZ
6rGVCvzBX9SsGwq6PgGZvIR/LIjgWJKRjoNU8gyD0h1GjJ+Z3UUDL6qOwmW7uWsrX848ETiL7gfr
u70sX27P6cAlVL6XAU9ykPoniX4bihTF4oSI8GSPGcLIRQKg9cRR/tMwqPrYp/zRukRnpRHhtsPv
Hea9FHMM0wUdLIlRR3pOSWFeipAaihMwZmn5DPC48peFmWnvvvD2Yqs/eXzjGqKP/ymlwpRkTN/c
l23EyeNwBvGhh4yhkxmZFb8BEd33+X6glwsUj1uECQpxmQvMiwt0swXcuHNnySyFg44ASqet2d3L
Id6GuLFLA9T2iB4Fbr1N9fjO1UYvNOvmHYBOBtGLA2C49CXNudnMUT4y/CoitKF+SoDg27KGeFs/
7Vbhh60KXqUmH55OxSUoWb4JmzXrIhT11oAk5HbN6aMPtEIJ9UZ3vUfGv5atGW0BpS6gCIsojIZT
qq5u6Cm34vO4VzDR0EeMLP/UEWw2UbyUAj8o/TfzMf211QCT2R6Lf0ethQXA1ZfQ++eQQ/WksuNU
GrG7i+upwuMRkN0qtbzov1+BsaJqlBUG3Gya7Q6YF7oHOT7tJ3EVW+sRMP3V+lAvzNrtY/9Z9M44
+PFljNMSA9kAMsg7i1uG/qWmGqUUzhSoHAEw5G01YOrRWCba7PU6/8ef7HPtubwXWq1ziklEsFBT
2LybI/zxOnLUzK60vkvFOVRqp5Uq2aYokpEZfSj9mrx9v01FIg49IWFN5TVuimuLSur8R32RCeTK
RPFtm5DvzOpiIUr/SLd7xmferBxDGfV93cY1GIS5RCU8AAIEgeoRHRGQy4BIE3NmTZP06mb52QEB
TCtJnSEA3uFi1pWoAiLuUhl+BqxlsJX0kFTX2VNkZcywgb8337HiPXaqGRi2141k/uGezCj1ryDC
Zi1f/0dZ0uO1EX22hEgvO0BZXBywUUzYxWltvgBN2uAAQIsDYNCn+nwt+x15J7Yf8pNKQqXGqdbW
UXeBGjNOrwCOqtPLZSIpuALW8VPO3WgvK4a+Onr+rg264OI8MKDR8bmE665tkVs/mHFQz1WRRh5U
hWfVaSi2UUNGi6vRzj/RQIfpBAGv6e49d3s/gEww7YXfjEQ0VdXlQVvWAfpDxqYC+zm3+LOqinru
zN9v4rxrEtkXyztUYUJRPbXYoEXrKW6vNpbfi55PcCUzfuy4Nm0tTtq9JH5OkGL0KiMOTMPKaMPk
fPRgil7jMe8POaFsJeRifMZRxOB45V0cLIdQFBW/Ze06FWf1suOn+15EvNbL7A2jIproYkedD3ry
YYSJucB4PmpnZV/60TNHX3H3wJWpso+vNA0FKMleBVhaXIQ6zE+NffyjPBEZWgBcOwPpSjonJDah
gKfegbAccWYnxL8M5bosnC6Tep++QSTOfXeXNGX7LolOgaqelhkdxs0iTU6Bn815by+4vyioQ1Dq
9R8JRrKvzS6EwKxL683HDPDfTIcpCUL69uuFb+oarfrfq/i6Wd+B+v+EPmFHU89TkG7L6YLlWMmp
yLN2OKw7W2hrhHMAo7wE7JeAL+yH3W30D74kTwzR/Pl9bQHKFhkQrsxmZxChVGt2EQLwHpa3gHxI
qlloh/hoIMFkmVFxt9KFTTR9eByx44Yo6Ii69aCIi7jOCkf3FNQHoQozy49R3rdLs7oslatmAhGq
wD3CDGbKGjscfY9hRzfj5FJUlfzOlp6A7r4pKsI36ZZosTD+5en1dShw2Gt+FA4cwFdfwVsUKPdl
MOflV6hwQMQfN0pNrxTAARwsmLwTq556J6p8L7+E5ldfTzKm1VWizw1ETtI3TwTA+sczfcyjle2Z
plxajG/DSI8WPsi0zqcfbJAFPiMTNFKkVFizY63rNA4C8TnVitnSo+gS3QKUgd1S1osBZEyJfVvV
4yRoKliPpUEOza1CPBUh4eqPFHxIXAZrfFwE/aDKYjX4/qev9vVk/M7P6w5c8AsT4ii5fCtAqXMe
cWe5xRoBv88CyObCnK7z1/wlb3y8G1fSS4kepybRWb+TSe/VIuoSmtqkwX5vmxPW6bpHS8fQ+mAz
Hxf8JZ3o+kq75W/Z0SW9PuEDsMneLYQQDXD21JKT7awrjqYSCP/uASovJ/wK0Fdt+UnX8xar7n58
zFi/Zi9jC1O9brx409JZiEdKJZtZo2kCgrN9SJ/4kqbggQeZprSO2oyaewiaHi3tBpFb8aS4L+Wj
3Lj4sRVRp8LaxtJzz07jZY/L9JUBngHKaENymnd8DBZsiLInVnKKAjhA1mQHsCdgaSWrNQrJQDqu
PfFHNSLCRp5167SZePGVRil/l0voiBPQhVzVuBFvm1I2zvYA9L6V8bN4gdinr6tQaSTYRTMYr+cl
VMJvSh9FZ342t0al0/QPWUSTQg6GsM0UnrCr1Q3qBmlNUQRNtspZmnGso4rU+iCx2kKL+On7Cvo2
e2Av7RX44Igz8BnxF8+9AAQrl4yHMwzf/nlNd3iayBQTk8DwSC9dNb286h8j746FlAKo74tAjnUC
ioA6IgC2T1WE4hPbenZIKma3hkVoH7azz+1xnJhdKXEz1eG+metN3+vSX9xbFpXookw+p+U9YSMA
IMZet3kjyuE9I91Ctg79iqYX4XYhimflZuJw0cWTZ0oMGQMjcSW6kJ44LpPzsjWcF97yv8qGNWge
x0QfdGpezaIAN1GGj9gjvja15Fm2KfuNUO9JOFGHE3eX/jefTWkaY5P2I0I0kI56zbbEyxizRduv
SdX3AQJij2fvMUXbpkKUBIBsow3UtzbPqnNbYYAcI4Vu79Z6M9+FQAEurA5H+9jvKnVx2PVV5AYG
r3dJlxpyQ52w8M53ZmwSBfZuR8OeTzyYqPUjx0EbT62p8jdxgYlCIiIzkdOLGIsaFo67fmC3+OBl
pzA/9KUwmJUCg4ireW5YRjdewFiAflBMuT16wppWMsc5KJsoCBmOfHgKdYC2fqEPx2pKCDsI8Xar
SOZiYb2sYulKKBY8jY714cDtTLiIh1Cb8FUFBIH38X/6r5Un0lnmx7M7PyZRsI1XEHCxbFB9WrLr
3iQnJq/pOTEsS+QiSOY3/yGzjvh976e9K/NXqMV+NkFyeJk2E/N6YIQ9LAAUVEGsLK9w6TZAyL+2
4RpytmtK/l9teD6X4fpZgwvdVEt0+LJRN0NpKp98vRdAWJgrRguVUpwazm5keAOowbaKdHdWBLvl
D5x6KSTRqmIsNXqlKyyhLJFYFxUcq3QmeN6GpfIOTvsnaXL9+ytyIfdTi3abMZAv52aHv59u48ph
OKhceX5YhXU53aLfS8lFDeKKG6EgEabx96RNSLpwIoVysBW5zNt02xh8WVW5XZFxjJci0ri7dMVr
5dCSIpUde/Eg5To1TGbbG8G1IQ8vxYrbyaXl9Ojw5TyFRRWDewJA8hWpWAxtN9gPiIAM35BVVPQN
y5gTlTx4rCUvmSZ9YWgwi3wD4g1FsDNDvdk/MnPyn5+CdIQ1nLLxD87SExNDCktfQH7Xp9Isf3H8
7e8+c610j6iNcAyKKpdyyjGdPhquN4z5AC9VHbQ1uox/jmBnK1yA9J+IAW+RLTXgWUg+V5DlZVck
DIuqiviKiLz2XFXKiyJ3g6dxH5J8CA7g7Q8Oocexz4n6fqfwesyOoSzhIWF9YZQmodFqU3dCAiMH
GhCrbwNjlU/out+BKsGxew/21D/NrqgTlUFF4rF4kPmGkhvXFiKSxtg+wfye9wRFXBrNJEJmgupk
zW75cdn3uEs4HCvHtF0lfuj2EEDgISv+T2K4lC4ms58YRmYiznTyGMAKcEzJAeBqmzeV0eXvlJZ/
CcO54+8kCQCnZXxMZPGQog2VfXwbHniAc0LGDYDNWh/OxDuD1h0Hqmb391z3cFwp+cBLJSV4Ngn4
JtJiLvXgkolw6Uq5cqMQ8jvMoP9pdrFupihAHb8MRKxaxLURY4e5EEZSuI0ClIVSCvxR75/OmsI+
T/kskSPl/oIwa1TRtSbpzWQUvbNPn7Nm6tDSYX/BbJClDK3JVirZaUeMaRl1h2NL/rOyZB+ovBtZ
dOpnzRw8LtPFWNecI0Bsb2rQ4rBhcy23tfRG9sd9+8DfI6l934DkOx8F47nP+oByIwt+xWPqLKuf
3UtA5ofLh1qZI2DHx+grIZ3PP0HPBVH4YDgPpuSFEdHKGkgomeDFTLF7tQsQK2B6YIMo8mL0S3/f
CmUohA44SDmFvkB5ph/UCDa8MidS5+L2gKp8rsQqwLzFEkWif5SRtscp38z3M5HRcbG9eFVivp8f
0BuwliI3kSAUyXHILnXaBY7TTV9fde0mFHk0Htn8yb49iBO5+8ib8UQZr0a1PQ2V7lqkgx1WKaOi
4a0VqszHsPCn+ghmvfkUk91S+v80fSdffzHBOumniEwlDe4g5ljFLXaaptUbU4b+va8xAV4CNoW1
z3gzRDPsnnUvwKwRbdxpT0mBBt/YegQolIyWVQpErSxP2Db0ZcCvLLIcn8xUZATdjrAOROuliaQZ
hx82lO2PZNnTXj7WYBa3mWtjVNzr859dm+2wfozJBa7fm7bIObCHSvBWAR3gZ2xOXimu70gzvoAZ
Df2PQubjIbH0tYK5c8FHeRkQB/ITc9vgVNaIIERvAozVS82cuNWBEwHMwExaNdyC45wda8CPtFTZ
L15x1fToYQEW1Ril9v03TW0tKbkmgN+DlZcy1JC9SD9FdPqCjLAEwmPeTmn5ZURznEmcEQ7OZO94
HGZnM2/ut2iCf4862oUQ88rD0LecVL6hw0MZiCS2i+PjtdqXrjKjmfBE1EPADtgnf3obL66kZ/hN
LqSwWOJmBo/tNW71VVcksl5n9MlwZ8Q1yKKPLLtOrERbdj3uhy1DugAmtz71HNd9+yssowbGeIgX
r3dwUVQIR+LI1tAM0Nfg3yELtY1iPgJ7jAIawfNvhNoUbt3z+ze4lFePo+J4LC2ZfgOuerjOSh5l
6NB567+WwugbCpZq2AqcG29gnWpBjsrQo/t7uBL9OOEDkuFO13KXjV0jzXAn61TSNWLLt1P5j9xw
C6yYHEWZ59J80m8js+Xa5lC31kbaCXJheYmjMY2jEVZBFx0Ldx6yqEpDNlTc2RZQ8h+dSLhwGK7K
letnXwCtqa7tX/BkSiBAOAgBAtE15HAyulpAeSEXMiYEC9QtntRg+neqN42Qaz8NBkGLqH4z5N5/
72PudysfiFZfJkhTp5XfS5iSYqmT6U1yT4RMvmsBm0KeC7PBkIoNm7fXaqcQ/gJLXjICA0hUH8zu
bCJGwivW7OhztVRWPddg08AhMMDRzg7DMASQ/bbOO0SM0JFgangiwGKKyK/FyVT0v7+KWynZHmRd
Ok+nTXq3/zNcBhKXayKgh7LmqnitB/ZBwMuaq7uiZBqMC4k4O9Uq/kvGDqh82iF436m77L4/0b3m
BnoKesm1dovEvlGjJAvn/LWEjmP/JVlYGCV4AgcUbKjO3l2J26bCjtwzL96Gd3Dhqo2f4451ZdYg
rQYsoygfm/K7YMckGUoYBSxo1le8GgMG2T6O6A8AGg9fSaIZijnU30Kb9irm7r1X+PPESSimyEdf
0ktyS3qUi7kFHN8SkieCJynS9lw2zYJv4uV1lV3ZWQxvnG5NkI/xkJcQKGnoM+zbAr/cLnB83Fr7
jcEW34AGGzpEtdHuoU0z2R3M4qvhMF9JFPh+IZm7dLecHycRgTYRJQb9qmYb3safm5l2EC8DG6Zq
Nzb2ZIBauKuD/LpilLL51DPLpNN57oHrW+9mZFBKbLpWW3tcJzIza649MhPtWhLElcAYAdFREn6Q
vXUgFG8ZmymtvUIdUUgz252PiLUf8rq+WgmpMQV4DR2WHcG1VvWtb5oEIvN4dLipAqgr0hdg3ALj
WbnZWwss4cFFu6RQ6B5hygHOOAaUgumu87yV/z9vPht77GalWni5V+SJwRJOCO+mV7QUC9305/gX
Yee9jEsEESYODdQxlXC8P506MZQdbvC6iZlWHoG8xUFcoKTBmqQls7/fqGzh30BU/4XKPIS0aGw6
ZBFN+n7t35LpxQRnHzrX4Pr6UqlR36Xp4uV14mW2lbrffdUmGAVZ/j3PJ8YqSqKH2KEx1AsqD7cJ
9wFKZZpIZqHHwiem+aAdWjHs4IXe+FLHkakGi24UW9s4dEBPPHEuYCGADE06HhgPySw4eDo0MFQy
DujWNsC0xAtkQEyj4ZZaCVIJEyJogLXWob5YdSKI+lsHw0N+yoKQG7t/qWS8LqkKNDXpBeXD3pg8
AqxtxeAWWaPDi/F9KidU6MoC3/GnKBEew4BmKtzzg5LH1j01sdOP+6XzJhSTCbj2GhLhjnA8cGIg
JNEvh3hHv+Wll8nbopnDJYOMZ+dhWb5G0f0ZioKgpA4cOuGdTtFOr0Fdps/XLC2K/HqMoGwAkY0K
BVeLM8UR4dsquL/5zBj/CvNeEqBPd1UQflZbTpsGX6NGOwh/VhdAKozRosIGYwpoiQ/nXddsrQNH
qlyvPL+MEBgf3vLPemQD/agq7llp1Tn0H+UQakgUZC1w/nUWk+aqZZaJvhOmuqzTqtL2a5pxL73W
0CGHyv+BRhZ0YLxhFfO1RNav1FT7T/IClquqJE9OWl17NyCXx1VxzhKaIliHXF86YnAPWaJhX2uK
IGOTRwMb9bMcgMbvK0179bpnOCbqCkJqX1iydP/wfM0YgjtAG+EvQgEytm35mN7s7r8eYIoZC4Ig
1zzbRcXUXxTjYkBvMEKV347vvKhMgj/YCbentrUwnLPoKPX5K9ATxItletpHnIEp6FagKIACYMs+
u6zF70Y1m47lwR+Oful4hdYZ9Dellx/q+1fxgQrKqIQjhcu9FsRPQP1bFo9dhG30ScT5PCkKAQDN
9G/Iqrqco6DAlR3R+5UevPRzVBA6onBzKYVX4cNQy7RcglvadsHzBIWRGazcYrdHmHz+VegSFuUP
1wfyre0gslQs00hZLHRFysCfrCQl9VRlIwQkxX8nMRjCyDU9uiYMclOP0SPHiLzZ1tLLhs5PMzES
gp/6wbTkxODxnQu5xDMPobWZXXtT6KHysOf9j6zEGRz4ovGtKCX24R0CCK5PKI+ZvlpmPWakQu7+
9mFwy4j7ev++yUJz5Ia/+6gkAEELxwyG8r6aQA+5YPGwATrM3LCFoSun4oENCCujdPUO1RBvUntC
YmIaSoooz6H96Y9jh6BhOVWx2IkuPJhG+ZTTfhVXdhJW91Imz8pq4bsna2CNkzI9PE1eKyxgjS57
phIdGyw2e+Ej1ICU5qiiWcV/GMrUyhG7LR9O2nxYs7XjYAHYgkukzxoPh2/+DxggeAJuPEvYFgM7
49paAMqD2H6rMjZL/Bm5pYMUMTBUwASTh16YSW260smzZkjzwOsqkaMwPIpwhzvrHCynOoWvjmWD
xmIQKWDuPg9/+PQM4V40FCq2APC5yAK7h4OOdBed6570QmQAjpA5xLFalGRUeEu1c+ihwiUbk/Gs
Xtq8WooGoBzCWFhiAJDaCiAo4cM3aZGXLLC/P0xrwf6eT29t3wt7LrHKM8g+j7xVzO+36S0tGVuB
WX3I3ZLP/Qaj788yx23epCUtCXHMe5M8xiUKYCIknsGfBNHY+GzXFTEtVlV+qRrv/1jEaDpIRwGZ
QTBi98+QYPwsbLjh2toGqNO9n8hl7Zdz1GCfe/JkSLeacSNR/5DO1HE4AFboxKCErYACxlEFlWbH
e55A0gxHcXBvzU8rs9YsF8u1SUHdh0YVueQ5PGMiEwkM7Z0mfpXh8zzEhmCEQKfywSieEJySm6hu
B90h1RH4CRh2jCEr84PXjOA9AFI5zL9AROPh1FH9H3NdfKWy/xEUozXymx38jQOwUJYxWNJJgK/G
gh93ZdNJ+VZgMjmNw0yzrA5AWruDWfZ1Y1IB42ZsAbh8lsxXGSdY7O+nOw4ymiRCKigM7W774WfF
2q1SkRB1lzQoD4qnlE4nYz6Tn/1NhYAiuNb8q51cyk73WGDqGYj+TyRJYxH59xOge6yZIn89TuSb
p8d1cMYcjdRzH8LvTGTzctIYAtVrxWobgYLziOf6rTS/7fxgNQAQeo2D+3OSfEUqtqrjZusqQBm5
Z6pXiulRCRc/EhsRQBSZhAexO2SrFJrYO8pnkEP6lgLEIkjFalJ5pYEms3qzWB7QvqEM8pOtIfzW
2bsPQ1A8ZBNSOPxVD/E7C5b+n31qnP9DnuQFfEoIR4RqxTLEo04cveHvxPNBtZnLxJdCLRuQyDAA
ABFx7Wp/RYl90mUHEEa1olp7dE7bIwv2x3y+i62vYSE5f206iFldAb6jFh6kH0PgOUJTNouDdwK5
+HAkBK8ESHmLjYlyO/SJ39uDniKvQaQ1RelnmP8WiBI15iedJTMrRX/SJjBqA97QbP4jWXDHeu98
ptGjww+FfwuMSzIFhxz347dtPPndHFZrxqSySNSrBOr/kyGA4ddhghxONptXxdatRNUHx+g9toVG
bWhMauFmd4P0h7GhyDo8YLRY0x1AydMufjypp/VetefFmehQDixDJsrgWeLxR08yH/YtzVksFqIv
NnTUXS7ObKsFUny1LHagxwzGImFc9Fnn4T+8GpTvmv7ZF001vP95GcfWLUujrVOD6HGEOisGM5Ae
r29OuzpUBpCt86pQ8aHu5Z0fE3l/qSDJ7ggmCk7Hlao7Omq9GxpRQJQwV2MWltwwm4OBxaOdDkDA
DvylIrxnMpaH1I4tS+cz4tkBafJHmaC33b/yJ8OnafuK8S7luTPBkUy8Fgz0W2PlBpYV8zyNbK48
c01ZkU75LX3A8ZkzX217wB4RHx7ca4VdAhr1MF8UTB7K0+aOUVofiwXzyn3p2Nd+UvCiSsP2HS0y
NU2MHBpIoPW22JlprA15As2g/OrJF/c8Tn2419097K0X+hRskM+1ckMwCpiqK/PIDdgjRWMuGBoo
zekCNJxEELuDNVOHXSrOU6muVAHO9CI/SK9PKmt1nbSMsspIHG7Ak4VDES8rpeMnfBCeS4G+sRPP
EaLlsoetLz2Fj4i5WI9q+icc3E276SqOdNCM51ht1wYmJPMNI0+V00MkM7Al/tAAZoeNGZUj7ENM
8R+sqKgm5+Q4btpya8676c6EXFXIUl3KjBlSQzGMhFn8sLRFPKdAAnT2e2gFo0h1hJvNBOk6W8zX
nMRHrgrs30RN+gCTdpH9OidvT6Wz2Wu3sNs4UeD+VlmUv0oowVZJ+Wg2OuwcsVVebQy6by/mkOaf
dPzc1Xfa0bm6UbUhP+a7NLBaQeGb1CfltzFEKJ8PHgnB1eF2grNYxaFLxD1EgixI2tCUHXC5BFQy
jLAo9alm25Z/H9/HGlVp04CGhdxG5TmSlFnZNFk5x6+Y9Z0e6dcJi/KhVQHGKhfjB8vvlwWvG26r
a9B/aIkeYRecgsle0MitBuBcaHEy44VDGakJ83nIjrQJ2NwSCzRpJ3okPbtGPEeEkaWb5o0p8E7K
Rxi58BMy8XqB3s/S/PJl/9yydNK6SGxfLDO6e8e83xM1inrJSC+suvLfjDegcJQohpfK4GdbcRgh
HS4OXdwiKpEFZlT3Y4XcmwlFu+C+G2Jd6+xCipqvgpD2NZOW3FuEYOFz0jNmTRowbHl/H6uUqUYz
YYv1qPmQMGdFduid/XnX4wcvQwKH3zrTkuuu7SMN1bURQFd/F37K2URU5rKUD4YfpyKo5K9iRFyF
SV+7fiF1YRaxZUxjB9+Cxy5Iggd97tw/mDxsPBguK1LObOwkVMnmqsTVquoLdo+gpoj2hmP7d+DD
RZD8lr0p1FJA2aAxwLqgSF7qQoLKkTsUQVp3tZTTNSbeuWjZAcaLeqTpimZKDY/IeZ6R3Y7g6l1N
uxJuuMPK6Nh7yq19oe02UOJyPyoD115TNxExbvE+AC7U5ROWMaRAzxZWvk7zlMQdrzJCoAlbFAvz
SfZNzcHLT2mtDkOHMJ+4Y08Uy9paVnOSBJMY3xUWrePlSpnxCqGB+54oXRGCPTyzsCJBNk8BjNmN
NeSlI5flwikqpkDd9D2rxcpraAgC5ROl9k8Cy7rpGNvS33YXEWUKhPgCkK63rmDc4oTAeKAeP9dR
/DE1wuoe3iGI3oF87hIWwiAVX+gyQpcAu2nqQctOG3zmWmevbso3BsSLYOsIp+YT4uaU8aToJBgz
JpSvJm5JJbW+QbsRtnZkhpKbIYLcUcGQXEVtH0eCYGpY6pe98GHtSo+u7fs8uPvXucjel6SWKag8
WoVeMLxfSyOpA3LzId+MwBGGiWapC8fxYo9GHQBXkLoXe6Db06CFgsi/eaHBQlnn8zQnBl5YuI32
Tfqs7jUHIRPXQCEsA+6PCtB1CR4Nq119CwzhjIt9LPzeo3aPclmVM19qYqMprur7227L+IapKoI+
klmiZ9eEse92loxihpJLXfgp0oflAUkfArHpN92zVnaAHGpffXYzpVLuvYPhH78iqRrahZ5zGukI
LdNHti00l3vXxuOdjNuHYdbvjPKPBsxO+ItHTxvPFvYVNTCUHOOCaOk1d2u9ntlUDBKsHpyXW1Qu
DOlP8XuPn4FVpu7/HpqSwJxUNfae35C7tgC2IAKItwB028BF70wNtF3ou6qc9Ro+fze4Zn/MhJ5+
TM0E4AYKj3irKVkh6ipc571i0n5u5UecgJRpebB3y0fq4kj4RImnTspEjgbqgi7O0+UT/JynW3U1
L6TSfwPkitFx62DjPkwfYYkIPZfF7B9tMOXA2pgb23GEucWxgSQPNaVwAoFrNEoAvmIpO99aeKCo
qB0B5puhRl1DoCLiEXzgo4yD4fTQAQGW6rAKRK3vMIGsl2J0YawiGph2SW+nsojo9TdWtGnnX2b9
hjml6bZ0L7ROfEL1uYl2YWBLDBTpouGUDa7m9Jb6nCkv7swLHuoR02RmDzP09vQxME5ejgFJRJH8
xlU47kGzBv5ggyTciePi2DTo/rBReebeeaPP4kIi72J/UOsntRiK9JTwACMi2QY+PKScPXpq2Rl9
l92Q6qZytwjDP7WqvxxGjJ8k4lKQmsACzY+0r+n9PsfJazFE++3Ip/vS3bpmy1HpxXMLRt4YM11o
BxiQ5lQLWpy/7khEwwiyvFJkWOrjg8xua/n5BBJ83M/PyCe77qmGTYbBxUasJ0TaN9YtF+FiTT3R
mk/fayqcG+K/4ifzmGXDd8l4uLEyKRuAMXJQHT757Cz+jl4l1W63mtYTdp9AbG+1uwLbyYw5sx9H
2khuUj8sAnukdOwI4t+HM8SlQ9qC3nUgrqRx5nzCch/oTJ0C/zqZdGIeWkbLLrUQv/8W0nhNfqVa
xEQ55iTCdjsxVSQfc5armIkPXXBJ8xkYXXni/vFfjIGXBWEBlLAki0bIJiI6798PiHV1I8aq4aMe
bU4+lpkKULfQv5YQDvHAMrQzidV6mK0N/zsyx5upydVnCGA0rwC8sNwxzYNVNqwgkaLKbzeq3JR4
NCZ3jn1tY/c3C40r6TXrIxl4//RKXmN81lu/V5oB8K0G+DEholNjUeWZVaBD6CWCEtRy3BMbbuDS
T99+WDdIE+CVFzIwZIgjUa8OMFWNFmdkEd1rwVtJfovZVtfjE0R55qn8Aa0FzeqGyImzGpd+/6Yy
WKOAvDpPHEQ64OvLx/LaOQOLK+v7NQa/y8p/J5fof7WTpbQ4a6p+h/R+oTZFrcNXEklmH6MWnE2e
POVKP/hFSQm0FuGJzvLpjvoNbEyoWseDg7PQ7otTLTnxTz4+mFH00mfIcPbc1F/7RZPMC7+3r+fP
bM44fjK50J0q9QKxAMTC/V+oj5IfPRjWWJ597Gu4nowzrfJfk1fGEgdsi6BQ6xRbJYeNbOw/KJsr
6DrDF60/1zTeTjTx19mPr57ien5+pzZBFV2d5O+DI0Kqtp0pv/9RoKCCNk0w9kHh9EleJVdDjwWh
LO256/aSX9VAbihevX5zNRKEWcT+cVgB2ECyIL0dLp/D9Lkm+O/DMbL8pxE8aKdn0EerWY7Ibs7T
MDc1pdK3NUyZQDp0Qz3dlg9+6+v3ZEO5CGra0+5HMZgJDM7B7EiEbvJ+Bht9Qi482f0UUiyiWKli
f6fuNsq7eZIBpfOzOlai9a2xA2vAdTFIa1vJTsjcI5rnYIYEzN1VXPPCgK3ADcyTrTpZV8ccYfv5
byHh3xTNdmIK1/jkRXu51c/rziJiSsy/AbikEV6eT9uP/Ca7awJHRBO3X9t9VJTAG5iKPMjYBzus
PXV9le6SI4IHhPnhFyZzrDy6vVvDm3Urx6LxzzEiyvkypO8Dn+OYZnLXKew/rLXAL3emElPz+Wsz
/y8EHD21Xd4t/ntU3A371j0fMSR05veg2eQNo44GjtQI6WV4xR/saFX88+a5P9czHyYk92kl/Wcc
CMJYKRbODKwEkge2QQ88MyYW7Uug/HcSPRVDaBr8EJfMEtXb4TRDovT1Nab7QrUjEfwl0pF0Iroo
LbAZaOUtvoMzz/JBOmV5C/AARPL15ryrNNLjOUZ94NDvgUmagYWHpFq2pPVkDHFHQj4d2XgsMeFT
zigXSCPWJQrqmR5Qje53dyqcN8Wum9zoTLtaNgktc4f1rd63f4vDMTRfAliSVgqkgUf+nDGZCiDI
LSFJ0cgPBiMeAcGWSPdIz+aj+p9k0CARdn8M0+H4FURsZRhzVMzdrSGIviNclH2v477JNiUXYF72
Q8ZlO4zsBh8cWdN9Gs51tn55qgugrCa9+p9mFWEH+YFwBbXATpN2djiyfw285xTSP4uvxjauzWWR
b6uS6bI2CR3gY1NIkzI9QDSVsVUAN++IgdZP19Q11bqZyJ2sROJFsuUSOKXHPldcBkLcbXVhdg3k
8OEK46mt0O+9rLWCjR+MvPTEHF9xMGU8DqzFYKIgV5ucSsC7mpn7CJvXIc0K8vRtPvhOmj9Nkvqt
3SiIIqx6cwNaeAU9ZiT8cHNlvq2RGhmfgDClStYTLqXUtZdPftJVOKwesxbjPEhLdRDWs90Nd6/C
HmqH5SBL3xouuBGpJiUbBsQeO1ksE2mX+wr1xdqLSbiRQrqpktQ3Jgk//hU9UP8FdBvh86EYg1B1
JflL/olZAIBD0b2hxIKWP1QgJGWwVDS5zXqqf52IkkhNpYnEWOxuc50QDUeRzfkweF+yNfb4Bn46
HYxNsqet8UBgX/QfhKUPvHqgEXSQL39whhF1n4HtUGCgM1dm5B9Kd/XKoZN27uL+qMjeFeufyxnT
3OzJsSLggp+sJMqvvyxdbm8CAXrxWzPRksqGe526x0+tdlCcsNhhTpWPLHAd8N5cSJ+NvdH82Hta
8yoSLgIEXVUaPKHqszCyxb4ta+oTmMm3FDTV3LUpwaATC6rB+5f2t2oFgBoHgsdXfyhbml3ztMl4
0DCuiTrrKQ71v7zY+siGJtEWjo9aRlcs9xJ5l3+M7jqR817GdaZMRVTr26/amm2tOxGaMUfauoZb
uf9DPIn/5Ya8NilFigGEnczqB/FLRmHg3bLyiDqdtQLeUFplj2TCs8rz4whnSWf0m3uUnlU3AZZO
n6wWOnkNhoM+a+6Zb6Pehh6qGzpBls86ic5C4/0b9CtLuqDTDy62hQfaM43WgEIiG1hJ/TgM2OzY
EskASzU4b7fY/lB+/4CuBelHC76aoMLVg57igNqDa6MDnJhW2/aN+G7WiZzvbRnIwnGKCcPDw6oa
X2LtMimKb5MV5LCH//aA5+EamkhjiewbiLR4niBCq10mekKJ934ToSoPAudJ1qYdE4IeDV0OEDxL
ClCv7/p3kYl4Tus/FvdWBrxtytDtQItyj7Sqg3Rnx5HrcN6FMeDV5JrDXIWUlUXz+dSmgczx6EB6
xVFNQ4K2EtPNWaphBop9hrr2MHJj1YXrSIqd1GUkP9vFkUwLy8Z4gnE7ClbPCBHCUgaikikXZcSp
9+MGzJoBbEmOorKno7A4K3JLeFWUtdoiK1CnB8I6jTsUqTLmT0NQYtxOzJDhqwGQf4X0T+azfNId
gPaEN4N3UdPc129QXmVgOKOl2HbtnzDT0ve0Vc/01TJKmLtggTPF8TqI9GSlQ9snxdcf9hqWDmNV
I5PyAmsAgYBQbzxqNrzyF2gzWdPjYO2saysDHe6vhB5jGnniS5BX7Sv3LvucrTTQUV8l8VmioPhK
MJwZLhm0NXAWfchmTIeH9Y0vH4QH/azYySVCKWEaXz7c2CnmkDGJU3CEnouuEXA4psA7j1C66dpm
uyjuDLLLw+tMAt5a9d25z7KKIclzgmCkJqcqh/TI5wI52dESoN4vqegvw7RKQEDIgJVw2VF+H//4
03SVv4HbdsE96h/HYEtB4xd8g5JjxNb1eYGgV9Uou0PlDoYefs8euq2KakWSx2UHqvA8LPmNIri9
Bu1g0Dr7Q2mgA1CKzZswsN0uRx82lYF9wFS0mTQK6eNgFCzCaXdv2i22tfQfYRoIQSJPzvvnMhlr
KWxLjdKWwodqo9wfxhr90cph3cO+wAdIZ1iATT5OPU6Mhk8N1/xqe6b+uPL4ych/2AZg3DfaH1o+
Qk3plowNhe1yHR8I4SYwMXsB9ZiC8zOEEhCptp6rA6x0r9oRP0kK3CGygKGufOGS0DAIKQFiFp5D
ccLur5LxmyFNWuCIFC02BvTbTUx51+NhH3QNXHDqKJ0nLZChaNxMd+gPttYQeu5TOZhDdnv1AxH4
jCNph+iwR3gOyzmb5nNseJ0v+bBCHpHULWvjBVRK/4Gdeg3dcFYJViieb3QZ2cbfz4GrKY+COUYB
lhssVsAXxYzKcdYEokINqipMA3CKV49MCIMF7rVQFgVWiuRE2kCd2ujiM1yMEGV6z8YBUFXznJEJ
Na7IF3h9P6EjnkxPTwtb0dSVVfk+I45qrHZWmAHBMIyodQYZx3mQ+BgbjYkcVDy5Bi3XJcRvV32Z
3H1V/jo13Pc1tlQO3+NqtbG9rZD7L50mWMQnl5SFlzCLME6Y3uqx1uW/PcB4qFxfpWAt+GFcUT90
fmzU/3+qj9E8andpNNbLiK7EjuQCLM0BMuSnxQ/cdLS6m46vJgl6HqIFEtoWieRw8Ub4aMdPOsso
WjWyy/+h+c0y3Onc17ik/+aJksgUzu4nUBszeiM8DTg81ZJVKqOObr8BPST/QBQKHDpxPT7VMRBp
Zq65rMUuVK/MEJId5zApSdJQKONSqgvUH4JQsfGbuBNA+KNyiGHV4gV7lYH9bFuYHUMudwAQAWjE
c1aMjT6Zdh+5dH6lNKaToY2tAkIWdNM8ZpuCf83Vn5T16mG1fguxOo1DsmyQpyxJPcDV0uq4y1RE
nMm+uQmEbaVt0J4a5+wP8MkWJVt4LqL8pLp6rUbee+XN8LTcPYHElYjxQrCZJr2OwM63hhlORmEQ
worxVxnbK3xD6EhRkfCJKAUn4F4cKyAcodI2VZzaYmgNyi+oBxCJ5tRbwnEUpTYthowmXQFzXedg
u8/AUlt5ggTET0L5v5XOfjL54DvQWRrMGDOI1Af4vteAxFh9ZBQR8ls+AKgJIoRjQso3Ny7pShc4
37V/2bejCRCHxvoFmDkYGDlL0muZXxz81R3YfPI65lEuKWKH4B4I/4Nq7JiwTCLPug6uL+3mmHHH
C2fwNjC4PA3UbpCeiz1TD1uTvjytcltlQXzYxFFjVVGHZ5jIjw0jY5YYukM8lAruUo3PtX50ZX0t
HOABeOHOeFPDF0yjxxUlQcjO5TUD/cS3Q6sO/rPq6DM+kxibMKkMVxxILUInUdA0T6rGhU3COJkQ
ckhW1bII6RlJ2Q/XDXtX1jXy8F1P0FD6aeRPZJwaUm5iCczPB4KGqSkh1OjoBRLk+MTubkwTm355
4sr3hDUu7CJJ93nojg3O5dQ7rxoqKckR6uZkNjgi1L5V0loqb4tFcoHWuIrkL8wJ0ZylUgF5Mnsm
3Qs2bdlWroS/UN8gR0Aycsj9yTERdAgyMYwB23/53pvI8qn139s1SRqTfQrjSltMEEKHqJtjYJTD
V150dnLCCtN4N25a1UbGIyK2fr0gamglVp830u3xIynUTT+bshUNi+UYbK/0DTHs0bHzpA+ZJ6vG
RAKwtnIYpIL8HDz7wcJWWKLN+Yu12/67vsKpA8jUyBq83QPgbVnsP4fq+o5/T0ux9xLD2qjdeNUc
5OcYlafVR4SNDwC+xZsRShMOpaOb3D19dwrOagRMIWUdq+53YZKN2S+KmwXvp6kPPA8YSD4WnEBb
gaetbpgfblErF0qaKQQ8okxJfR/nV+Tj0twoQIzx8bkRhSP38/Fjm87CFTDYhq1zQDIHfV9h5uUc
5CD+hzPwsZ7RWPc5OhJG1ric0OJmxrPa3/zKur0YDCFx4qAyI+OymuZ+rEBwbPNQUMVb7xluo5eb
eT+Efd3SPbhMwq8g8RTZHUjup8o2qsQhuPLS+ROIyB7eRPHMpi5UShmWAASOdhTg9VxpZxIZVrfZ
a+cjqpiX/igU3+evXrJj7AAyf8aNexRBDc1VUOfGKonA23ykKa6ngdDb4v/5KWhlqKYyYp31031w
xdanCooPR/BaxBBP8acMMkM0OoN9vsSPsww3DXPD9LqisBPubs7IrfAFp52HRwRlmkoxGSK8/zqM
k+I2W9X9qa2MD6RDA8jLfus1x3PccqO6FGiaTqFRv9tl+O9d2upug9ZukAfjqs9TntPuSA+YQAFB
W9i4XDSEPoLKTweneg1Gmr023Rv+uc7xPYnCOhnSjupCrMl8jdAK+XWXJC9lHRNYYWtjw+OwxB72
4VqLXA/yr+qkJRd8fpAFogz3q4/gSc/Y3Gdm0OeE1TldLjVLDD3Me2rSUTrt5C8cy9UBkfK1sNTO
aaTfPYbS1vkQT4roS8BHpjAt8ryVIoKlZ9kUC8lvbXJYUwg36xV4/CpxnLo1WJ0LeYi1gC2hgM/S
lXuAv8V0YBPwbNJ9LznMvC1/SKFyXPxhJwBkjM0DB1bpsYShbPMT9YbC/M81Z5Q2IOKpPftqFH+I
ErITYoyPd995D1iJoULHfckYdlzGmmIKSMq6kf+Y4J2WmQDCyMSb1VNbWwomNjKIfYM52+g/g67G
5p6vIdAgRqJCRoB9SFwP4tbymHXpLSe8VRpQTYRdD0JAlfdu+NS5kmAwOdq4YbM4AUzNZjfO6KYH
ngrHOPBmwzigv/5/6OWp6GTTgfOfY+sgbFFF1GlJK51ukOydQgXE9yppUvN4TOyT95ecoEOmsS/H
AqBhb7rp++EyB0bWlsRgK/wkuW5afOrF3OknptjeNXj1QG+GDnkn5ArKiuuMiKeCRtiTm0EbB892
kfTKIEShB1Qi9U8JM9cU+DxNAsVPEoFWn2z+7H2dBiwdqzXbOjDRQ7lGt7B72841X5lxegHTSado
+GmaftqIt5qKHsMHahWzgklB4rB7+XsrSyj07Dl0qJSvEZFowbm7U6NbYJOylqJzRLzGSWowFg99
VPd2C0HMA8ADR6Mdqo04ZiEEK2AtfB8NIWd7sHBJjFSprWdPo+VYIsbuxDTpWUslTXIts/1MiLV9
XFK4dBTFvq553ONcJ2iyCZvQ/jK3Vsr1YkUU6MpiU0EiamP1M8hXhyjAdvGCrBZL+iENN/SPriLU
QtJPk6vUtVeADBdDf8L0Rf7FrKzKlB1TtQiQiuesMims6AnjkwpifQ2IaGU2VWiHDBr77g59UbOr
yIugmoIqECznRTDkxoV2WCdHxm9iNdNU2JOyxckuL32+Uba1I0U3L1I43WoOICj8qOFBl/NCjPoM
uyLN2LZZ42QCXRgUs89irVueElhNqy/LDkyKqBJukalUtjUx3bLu0vtXpnACiIT+kZGlMwgTAF3b
yutsXFJg3j0OCPu40MGP0OtO6PMCrvU7vVUtdB8/+e8DZXh0YhdNVXJEZrPIbqjQozvvzMV6Xtmf
88LF6KoK369G6H3BmXebggjgwiS+DE0RlRfe87xhiddp7+WZiH+Mjs2ujxlBuvPXLJyg5ZhkNBE2
SpAoAfAjcQ9grQvGCD+2NyDHjsaGo3jScp9wWwa2RYu1D+JCgb70Z4eUzp4QmAmOMUosTJRCntf8
4OZhrXVPhHBCWIyDxYemIf2P7XBsM94xoejSk/KwOPDp2VCTO+kNmxeqiQL6sx3TyO1YVLj5DY9I
hbgq8k8KrjSoiZNjPI3VzBNiqloNctMCciNJwxpBBmNyffHFExty6MjB7tXAVaw7S2CGiMnX+zpM
RsHc2B+D8WxJnOFXotMlp0oDzGY2XI/0SYtyMimwUnBl4GNTLhUkOQ7Oolx2CheXZF/A+/lDkP6z
8LkIKpv1CXuXTdsvR1dLCVHtIRjzHCYRqhMn/g1VQo1xB9mNWKV7QCjNLGp4yiVVXEqcOkMgzdu4
Kfo4Af0iR7QdUUF62X/B8pvhPlQljajL2Ocr/wqWRXU9qIQLVR8zC06DBeoqda8q3bqwA/whlOIg
Tgo8Zzuvp7ZpbryxLLgM9A2n9+tG7ogukub/PPALszOuOjfd8KfMqfruZbvlBCBUb3N5SN8dHV0/
7nMBDmfyQUksNAnNIV9ZR9yuOPnCKVVii0Ka9T4/G+cJ1O2qXW3YKDjWfNdcrtQ7nre+nMhEB0FV
Sn9JUEdzYEK/EKGcMNp6mbSxb8Ob0TtZJbMkuJVbTPf0BDWwdptEa/zNG2UpMSnEPLNfWZWYmFa1
ZobG8V6S3Snr9484a3uNAqL2gMFynRZHBqRHfhT+rwbq+vCq/Gk/COQal15Ix06fYlTPEoO6e3Ri
EY6SNhcyD81AQYHSMRq8ie9bq1BrKHg+75MBgYkHmcQBEljixFEcDl/XGt2bOSVmYtNslNNL6TDA
x0YueAcrBibWtpg8hfaCf0gr+gMU99FS+5hTAiNFVicYh7f/OIymNaQa8XOF28z2v0vxQlc56BrX
euUQKDV6o35EWP2/x5AO7E5hZnm4JT/sxXnHp6XsUMMlm2X57XPk00OCfjCSEC7MYvxnF8pDkqmu
BPtRdzEwNPpagXdasvQlI/ORlQq12PuwKHAo9JaCb90HSJZAeAmzv1agPVIvAwgHeNd9Rl9kSR16
UvoA3pFbd8u+Ye17h1ebKiJPAjR77pbHccsd6HX7gPDes7IeADJ7Dr4eOd0wGCaFl2yzC/b1CeXH
Qq7xH7eq8vpZtkeSW2OBTNifih3Pn7C25aMeIPUYS0JFxbiROh8cM1gxQlLPGyTxScyJVRje4FS1
+00Z7Skz/29BUR+EfLvKmv3p+kCLaPQA52bi/u577oFg08AGylQxUTgbm/rWJc6HA2fUwYQqITUV
rDOlZzVgBC/5vukhESHC31IS4tQ9HbMsVkyxq7fd0oMrcbagwJllday45p6pBk1xhC4Hl8pMFhHR
aB5ujQz+CaQsBq0SdM/0DHq4ZInO54ADZ9mt7yh0KfDZXPnScjJg2Wq0755OvlJ8MatUvQ3jAXi7
jZ5zkS+hEAu8ewxD4GQ51v+zr2n4MqgoxoQgv9QOVwhVrjGpB+SHP+ah4oM/9ZqCwMQH+Epg3+Y2
Y683Z680i8xPPofbRFyRSULmNtQOA6+6piZ54iJ7EeQqOKROOA9le1cFYgB6H5f/CMYMKZh9fE/m
U+TonEcUy+P2WVaIuzQb9m+01KChcx1filVsSizBsi4ryQCB3I9YiZvVVM8GrqEpR5G9Ec93dlQc
dgDz1HZjIkmX8ZhzAjyN94v6uuCknsHT9VpDoXL5v/S7Sh7z0DuNQaRCE1PkdnA0XbGYZ5TtGmSa
SPh6ymr24ascWbFFFKWr/PlUDLmf5z1BbTc7vayBxpmSaIi+ApqA3tV2G7f+K5gLa35NbQhC+60X
fqVjuBKlDAD9uyQYgAxG4MXeF/vgto4KYFH3jfQrDUSLO3aXDby62rqt0AR7u/eVAX1XP3xZu9hK
9Sejz3nEuzL4dqA6LvGlb5g6xoLI0j7n2ObLH6/xrpGCy6i9E4uE4mAGz4vpmKqi1fyngbocu0Bm
V5GObesPxY27HORSUN+cgSY5JcXnZA36Z/U9rLEvdQoyr6qbCv1Qw7crrDMnENG/o+QxvXvFfgSp
Q/1jt1ZydUuTi911cWhrBeCQ9Ghshlf6Y/aC1aH6VTqWjKe+1OD7QP7DZmmRIwpO4ipqAjsb4rP2
dHlwKYVzCAMN67ABtnRkZQjTvemLQqvhmTqiganYj3p+hE1doPoN0bw1//CKtiquOdMh+3GpkNss
KTpNQEKpEiyhQgVHbg0256B3XqVHnKbv4Sdmy47RYxP0mmU8TJech08T7WIIizDuC7rxOqHK4RlR
8vn+HaAP1wG2e76zH0iob6rz+HfYtZPZWzVThRH8ds9WddgIMUHsBXoikbKWud/AwTeB8iZ5Icrz
LIICV2cq+ntfPwhztljFCgzE6ucXQL0KYz4VM07i7kbIU81U2iYERvAzoyueNZqfGnl6ucttrv8Z
ATWnVWflyqirHgn5u4eQB707LqF8C4y69PxGrWi78RPykNW9dN82rcpjBqEYf/CVaE50wgP6JKp4
s+W3MT9L0EN94d/JbDu70RPMbrU402xinhcTOZMLfYjxYnwy51bJG1m1+me4uObd2z3LNHB376ir
wSJmUVn0cvmKSh8xNxCcoNUdl83NqfEshTlZc78kNSlhNUxcDcA7L0Yw7VNSlHTBSxAp8Ez4aIPO
ZWPRwwHmgY3MDFxiaCY/aGZ4GJdMeYg1/ROjlSqYbkbo9c2ytq9SLHOrj0/xkxgAC2iZSoLTRP4r
UxB+ASVP1iJuAINq+Ft8DrH5CR23d4KXCaqjQpCbGBkCEAtKoXXMpvI843pamaSRLEPZQuw4qSwZ
xH9F/AV7oCtz5xn+Z623aDrPVn6AqugW46k+wAfkAwHmf5ZkZfK8m787QGwlRsOVuU4Rs36Ez2lB
EicJP50Ey1sfp0+bwGEc0izhmcux+o2Uft9ukAsi5qOT8/HLO+QvcbRj8nRVbqtKx9Ufvo4sh7Q9
dttdPVGAvLi23rk7eyWm2HoaFC4pOx+/+R7YviQw6bPkRc5z2Kdr6mRlEYldnh06GMnymP+h5H9S
se+XPCA21TytT6fftcJOkf2otpFBp1yR/CiZL3SSc3iq4YZLpxno9sHOrQYJqKmqlqWDyMyvEMAz
IleVQ+Hxx968WBO8MKt7PMuiiLuMOvUcEvQWm6F2ktXhiFGAM5vJZIcG3UObDg7s4MmMWXAsrV08
uXSKaEYxpThDXeD5ChInvEUP41hgclnhey03UHGH40ABtSXrlZpmfzahxDP1uI/cwFyTfLLMuaQ5
bNWJkB5IXKdfMaSKstSAjUjfuT9wqIt57tnw0QQlgrAR1CpzJdcWc41+k9PUoXvTTjHr3//p2fN0
U3C1SqyQ8TVc0H8JrYyL7JCmQHecOGcIOYeRwbshpTcCMAd/yIxdUMcCg9G/+2GJI0OAw3sKEgzu
T2R2fmGi7BCd8tBJ67WLtQ4FXCcI2drpHnHPgs0uVGH3FibBpr2BP3ZlFEcnm4r+XvLwPYc5PBct
sV47vHFChnhJKQ0mwQMoC2gHbYN/yVyn1AeAczCFLsiLIiAyvNspIvIb5Y/RiUgCOKXviX6aMvfT
KPwyfWTQmzObqRI0wd7N5sI3ihB5iYQ2p44X1qikISw+0n4zyGiv3tOhWhncw5e2CTBEE4fntJgl
aEXpfrkfVmX+CHMM5MRU38ZfNcWfytDmz7gqRa0tz/SX1WTWssfklBxOiqkBPn81ZoNg04qMxxnW
q+dNYc5k0kkPM8oNs4dkF9tpdqr+uQFRSJZD85p0HNIjdh9eDjwBwwUvYRPBAtjEtAs15YoWe0sK
5seBG+/TdVFwhrXjr569oxJaFtX4y7UY/53juZW3PaGc54NVXTZSvr98lnbPwFrNH/faYJsyKc10
mUSKaQZBh1/cSEXBe5EOVuXB++ELQdxBhNQbn/Oj4bsCV+UH4/DyOcjRIcBJayStw3nlcIGHxGOP
x4zVpk8H7pEI+SfeqM15WZOheRDJUpCqb1cktUEBL/cmTILO2OqmXw/hY3vgK0e/wvcdEPMtc4AD
XZCugJI7pKI5tfLGKsqi54uIAqFy5KO9Oia9j7IspJAzTMhbPqP9eJHIcApViDvsNlhkVzE/qUWK
JomZaJiZsC346onl5YzGG2CIcge2xO4wKUPrOMIUss3VFdGxp0fA15vBiIcdnWbgMwbQdZMTUPwz
K31UckkBc078vWo1hZWZbTIhpc0Ya6GVYiuAgV/oYwX49dqYB53GbeDacB2ZPyjA2jfPaRGmMIGx
/UBytLHV8xlPxaesriQfveMprTYsWcIc3A5ED0iFvsTuMUtBQrVK5dht4fHTKY2vyy+VF/bnXI4d
35mT3UXOcIZNhQI0lpzvZgsr33oC0DfL8h9raRhFMlkB+SQySSNSUeV/JyscM58NyjP5jW6hnaxM
8H6sUn0KlIensokTbFaMSSr/UrvHxinUtRC/dco1FIUMg8zggx6z/oCGD3ZtZBIbUQtOwRyIfrQD
L88nAiQ5uuwX87ukoawweZxKOezK5h4+FYX+w6N0tOqxaS/rMLkuOYrXHmnv7bmGMexoVrG1QEe5
G0KXSxz+hsJglUV8SClfGizpqC6phajIhzqAMZ2Usr5zIFw43eo+dRHEUHN9n7Zo+bp1xlNAwg+F
M0IYSqSuwf1JTU/7QUF+JEcHlVf0rN7QQrveMulqtEhSi4LEqJrsmCjQHGb4NwKVEgmsft/Uz1Wt
UwBZFKEOS33uuT7z0cDXKOw/yFrAm8Y9JeG0Z4faHSXsXcIEKz+O3W5Oxvc5WfYzUo4hjDnudCn0
DxL/F6S/jfHoQvS4OoeKxjaB4lhDRfcrcm/eo/lpwU5sFlrWnbP/ej2Np1NMminY9j3c7Q4E2l+s
nmzyx9X55q1NPmF8QI8rU7DOPVue918XJH3b9piOcyTT4aF0q3E6+R2y4VGHgfZ/XHCkc/jprcQL
2BY2q67q+DO7wckYtDSaHeiq1BgCfHPkQoVRscrJIjwZfFIM0PJa0HdM6FX3iAM5J0knJtYZTDVb
QDiShwdji0BHMZMXOTGFDNJCjX5wCjdChF7NKyszzbnPykR58vcQHeku9HZfxiHBAC2Lq/l+J1fi
079P/y3O12FLJQ9kB409cJWCmKKLDf7Pf4qUW6F8yQQqadezCF9JaFhUl3paNcw4ErJ+YoJ/+35b
OG9VYfhFd/NBvwU8lQ23wwAiOpISX+T9hm2l1DvM4FTAX4zZqoPV9ilqXO03GWLPODWvJCn/5vAr
C+Np+2YnbPyjPgFYvtx5wcch3QBcCKCe/WzM2AXFzVJ4egxe4kODI/us+kPi1RRsHOnqOZz73cHn
i8eaNWc9XwuP1uUuBjMb7hVxVbLkG4npMKxZ4gysHxeoH44e6oyRK/xP0hULI+H9VTJs1KYlVpBY
X7eXBWHyuMnjVr+XT9ijJneHw3hG9rJGl2a+1RTL+WUYAEIIf6OjarP7eiaQvHejzTwU4juETY9M
0Hw665Zi5E+iueL/qr7btpqkBEQZnQ38m3/vC1eQQ3uw1l8vWtPnV4hWtH8cHPvdjLmFryrXxIgC
dRn/4PHqn7Vn32LiXwtNXPxAXE5vRpk/9PMhL17EtLoQyEhzS4p8Rc0dklvWwxhyYxLfL0MQCVOZ
NtX8NzhkrBEVZ6U/OUurtYRUXGe9yjtPNH7+eWSAagqna0JqQ3NMuVh7BIOQ/bz2xbpp8vwm1T/N
RKo5vd/Tbb57QAB+7fBGtye8xZ34MYjQ2x/m1MmOavq3TQiMy06zF7pP44LmKPd/EYhWFakZ/Ip0
J+kM8MgvD3D8LD+RnMf0u7RjrG3cRHuFICdrcPOchstK6425XIdC52O71c6oTZAKmxky5rnjTqy0
1sSvfU0QrE80+rkcAZhq8XhnUQGDqFhu9EXVRik8myUlMUMN21SUQY6H3f6fiMIWPEPeLaB551Ff
xsG3KPQiHWDHNhJ2xcc13GUBKy8VMf4I/8wRu5OeB0b5/XqLIJqEjjc9tyBrVhplHQeSY53WMx9j
HOetRkG3J+GcIpYfNAnkF1aysQzo0uez+PitXkMZJ/uemwVNFOuSpF9R3aK9GI4zwcLiK+93V6Km
+rahxBMPO0mMTpcT/SjnYitvUi+ztm8Io/245RHL07EgnBoKbI30shVyctZMcqxGoohPjy5hjtTY
mZj3A74+ta+KWeQ62OaICJtypcaMSDXdZBs2+HZS57xYZlBpXHweOxJ0lmnNtCBR2gmCGlgB2Ll8
vS0WLoNcICsIh9OrRX2nRNDnGnPd4SaQTPD9Sb+6pvP0ZomGF0SfnRlWdtfRRGw3kEa7yDNZjTZP
sIhMmRgszSDCxc1xTrPr6jnrBKVISYXuqyUSKH34nOmC/ad3NKQCw8m/c3oOeQRb7lLeCY+8emaY
065i8/C6jf8VEd/WVpCTgU7mjNWWHkTKaFa0ADT7Fa+Qn32l/kbLYz68hkErbIvVz8XGUL+tQ9bJ
GxhOoTEWpg3r47ijBQyKcqS1awbQRaAsmIkRQhRwQR4zjobt9VcUc/N3x6IGFfBiThNjvfndBpbE
3Irkc/Iwf1/FG7vzApK3yNS2OlUgitoWb4oxuD4VPGwhY7E4IDeS78Uq8iYwHDxOinCLJwC+HHf1
joI9DqQSxBZsvIRjuc9v2H3q6oeY0N5S5v+o3XtaLPcATQfYp0mF0ddLqQ+yo2gq3vFqBpHAbtL1
qeXauYDCC9XDNcAlNIE5Ss00b1cfoUGdGBid+jmT98/MKfur6d28cszcQUoTg3F8YFp4rN6rBefn
JFNW2LPg8ZvZ84UPBa0S7sjJEpSqF7rVr4du6s1o0KoDzexJUdrBxvnAci83AGZc7nleoIbxcbAb
nZSb5FDzXLz81XZdG4qvE6STGYLZog+vgOSSQUqM8H6c45ez8RcSRN1bjXfFosW/zeUL3rEGVbqV
asKOtfiiHQcoxERKLs6NSRB3AHZkGnqFNfhq9TiPMmR8r327eFLeS/3PL7xxWPawyvG+tSovpGV6
X4A+hdZOhhlInk0JPbpWSMONzLC69tlbGwekzE/ZevYwgJl4mtK71n1sDkrfvD0MC8sYlQqQ/d4f
vYaZwqLTu33YLLsMPmwsY+IKC8wbekIr6V1J+cufLdmEjlfwMgf6gKGAauYJdIMNj7oIQIg4JkNk
23hxOkEFspUw0qsPNdAAKIYYAUPyilXEa826wVH2TYQBFwYE5vJGTxi4/Fq7ydtxVSLnRE3hHAbR
hWipZxB/2IohEnprJPyIb2ki5D3RVl1Xmhq8NGNBG6gNX+qVWOjuq3iNgafsQqzA4I4eK9apaS1M
ZiWH1ZFBB63kW2Pz8xbR86NCC3O+0Td9lbNJN8D4+i1J+lQAnt3FHk2A0u+3HKVV2myB9DaHVQi0
JvRvzdKq+c30HJNaG5ieHlpvBNAoqhQcrRoxDm9mc51AInscuhPUUU/mtb1vcsJYtENzrb3R4dSF
cJ1BjUQt7nkoIHq9Zp83X51Sc+4BYdd3a6wSyX3LNfM8IWqQ3TCFrXJnSPLUGmYAM6N3bnYccDfp
SkJzZ9MtmNskNbxukld9KmOA7uAdtJuKbJGdPy4/gcqZT8Sktp6A12bOGzPsY2lujeRu5vlb7P2X
L49qrb7AuKZlu2xTB9GgRAsRKhECR+7ylMv2BQWz85uEcS1UNHYDtVgoIkPAAF5fXavCa4oAyTMA
Is9H5rryydjOIi+YL5/XOLA3DP1CWjWpgjRfljIfb1nQbz4WLPCmHYyvIScNUcTYBrKErdTjJVbk
NvqhByUKr6cHno2iFVpAo15NGTz8z57+FyqOiOdN2S9GHQZkY6B1sTMy/NgA5ow+fmWdURW2NUBe
OQ/Ld7x+d68nOJrxCGYloHJtSu1boQ/ECSXuFy2bZpFxyGqlECQY9+WGWuurNsQNgc0SdzGGX0I1
ahrxD3edPhMneSqvhRTGtqtV+hJGHAj6nWxMG73HKsnSmJ7M69jczUgswZ1bAYsEPddx9AyIlL0m
DDP0axJsYVGFxGY81y9wbksAPbwt8I09RLfY0P7OCXZhqgr/o34rznMb3LyVgkgag8FwtQ9ww22s
EeDyH52gtFz1f/rBXKBBfAMucSngdWQaTM0Iu2yGduGY4IUI8CgtDGcVPtxRVFH7uZ5coTdZhFSP
H59MbX0m6zlXrp7WG1l1O5RTu/ANhwxe8egm50RtmBNty8ry9rCht9JEb1+aJyMrCqGlYc7J7xHh
fQVx3dFl5KATNWFq9ll3DYIqwPDEoFtiKToG48tuGEBnakkuyyKEeqrb2rLerS9Ftm3znxQQkizV
QVjXgEHlHUzVXJBxJvp568RWD2f/T+cs8W3vHGVBbQp1/bWJ6l6HjNEkbbdKtATKASSM04KLSplw
3mIcfoJpd2Ter3v9vzEaitX7AqFqmjfHyLAr9ZdCidRg+uTTlBSE+kkhjgIdkuKBqEn1i30aJEXy
MBgkSvWQVr2rL9ygdQsr98g6rSxM19UtHFKiUC26tt8jBtiVCVBBlcqvvH+pjmz7bzwfIAiZ7riz
gaYi2uDzCAwC4eoQ74HtKbFGHhn+xje5r0gR5ikuHOC5pz2miw0w3MRrBXNPM+v8a1RjuwjBhzxN
9aWLFyj7LGYIk1C++hXQPYBKQL5ZvoydzTZdsh8CvflZDvdwnD/QlKf10v4y9hhKNqweGla9+/Vw
LVpLR68RDk7tbEyaO2lnGQ3LQwsHDczm4ZT4ZULzoAVird/ThjFkvpXaq2FsFpqwB2xlXEYZkEQs
Qf9Sdd9UfciLFrsgHbA9vFgNUKp6W1papTjC3RVmyxSXU/Da91fUoW6F8JK5fZ2rzLP9Exd3QoAv
Fsc/GtQrLtd13yW0X6N2TYyMz1HiZ86i1MU/Gad6CF5UkZ8iiMg/wym875onrwI2zSahqJQvY4Mr
SjXeJcQiYbmvaSQdpihgxE2dlLbkuYy2xKwP+I7ucdfCmQ9tIUEkuCbsb8hPmoRKqiD/23fV8CWu
cNWJkKSvr/5efTk1JgTd9AVW0ooC+RoYnrWE18VpQ5cbBx8rdyIA5sD8fzE1oyzL7YUjXgIg14K/
NRkMqdhXnhdE9/KPqac0z6E94YQULIyV7XH60gvLe4h2i1vDzAEhdjTDZiwl76+zg6+BLAPRhbqB
rK4Ci/Zh/mB5gAeHEC7ZISOsAlIBsLenPRgkktI/CVCi6RWITnv4mIjPRbtCPK+5b1AyIdXWcNwv
toMiju1YPBZ365PfIEAzJ/CyaySstzeFv9Eb78oCJ0zV9SLv7RLGIuYo2FDPQmgb+oX5p4XdSRbS
/YoNBF/EDTk1f7LKrWUOqwW5S/rODD7ceNt57NByu28xyE200YJb9EVHWVUKaDdW3lo9DAIedopC
8gywI3HcoWVj849tEzQa6x2VgrihlNDtu2VwW1kwbzfCzRquCMB8KB+nhirurSuBwk92cNrxnJWq
Mu8RYVsztI4DmwEyKAIYfZ7FfJBP7xBFzAW8cKDFSAGa6l49jqCu2DEn/ocHwdtEH3bdciaVIDHA
K68WUvZynCCRuCfGKSdceo1V3dYCBDdq7R/sOdx9aS8h/GV9Uxsu+RRFJhSa8hWMzBIzM98kRpPK
21YgaGHdz6UPZrkvNQR8PU5H2sE4ZOXZHGQoXIg5LyAPXpu76Vqas/3mjUVz8qmLTQPjYL+0Z2hR
2gSfzwKM7yBeAsmElIRwxyidHGWbh5yz2oL2D2XTQsO2fc9mX3r0nZRmKVzQqbn+q+tupmZQMTa3
lYaNe2XOoKTXA477zANHz6blD85T8zfIRhHkIQ9fLrGQKsmX2bC8eWIKyZ9e/3yD497UnWDBMkHu
J3hUOnPW9TtOiPQYCT7wkutINVmND9xoTQsveHnW7ooFPD+M1FhuHu6skJwjDoNfCvA5oQOj6d9O
//zoOHuenDA1yYU6WzSgFG+V8HRJkUTB/Nf17rV/J7l7EMkuTUDBE8X+MzU+KCiiyhATa67NL7Bk
tKgBrrEdZmhcroS5qTON06R2pyG5i9YM0VF5vP+jl7wZ449csTko0BsljJhHS4WyM5DID6/1BBTW
q+14fJKEwh9q5o2M3PrA1PuoXVW2PSEkrXaPEXxIwhkZCVypZkD/98kPWWs0q/LGq8jtQyuAgaGL
8l5sxaNMVmNWcS9VvjPwlU9XbuQkQKhrzz/iBrigKCwyyCskcJysxlcDBH2p1mVzIkCSKW3dN8SQ
LY8Zg0LoTv8b+dZoy2UAVmDURpF/zxTmsfmS0aJUEZdaHoXgdIFHQtrUpWNVnT18dEebt7MTplv3
KuldagnuojSoNgwMYg0zrYYTkGvsgGQZsbNbbRJqqBZG/UytOa32945kxJ8F1ca6L6Cd5TV2P3CF
vQU8fdqrF9xWet54ig1vKAz2haKweMwApcMY0IYKtczV26dw8hdalIVCiJheoDoyOI0uUzArvwpZ
AvKIfJUTLBAHnIVYW3u3kRy6g59+HI4xh+vBGSvyU+OifO9+PzogTtwAD4JFiXo+kAe7QUHZz2yL
pY3X0HufiT2YkEjEQdPlwpjE08KlaGWFkc7v3ya16ZsKn6fiWQHkg9RsNOQZ0qHjYfzUQiaeH03h
xKxnlyxLH6Z/JGvdW8GFgNMaZpCnXErFG5kr2OmUvqxcasHTDeN2v44OkGRyWnij1jHCrM0mLlC4
3Eai1xYkqtefclR20seoC6fGeg+my8f83zxIZk62wV2KfcAXkJuM/qFd8UDT9YnjdSO9x8aPLkzp
0eCNaM5hgcJzWMfX6sDTyXgTUdyIuvn9WbUaPxg76jw0IK5OIYPxsHyr4A+891mPxVHL5Vs5Hhnj
AnGE37tZMz0THtzxT7hCpaa2LQYZkFBLaUSn//cej2O0rIIdWiyPx+FIY9f4+vx+8FjHTBJoWzUO
SpYNu71Qv1GkJ9kHXDuw6t7nyXbl1jMclic5NGqkcRq71M5+CTGBBOwdiNgeVrAdvIk37X5WnY1A
B969ICBWqfAIOhaFSmvdLhV/TaBKBa8Bke2EDoLBarxhqLoBjYc1U4Hy3k1/5XcYktdh1uh9nfNd
odoKKCDAtX5u4oSve/cNgQk4piCnL5s1hW+D4g148yPqsdEA9aM+MvX20iQgtghDIyKpT1Ys1eUH
OWf3eKEEqYt//3oPJecBYB/SziFYR1WpzUG9Wtrizs+6BB1k9xIhyt+GBD9ZzdTm78XuxZ7qQ4Ud
2Se8ZR+D2s/UNKWu0e3HeYQretvrszbwmUQMLQVvvxx2vwPlYlDfc/tLvFDVzkqx/Q8JqUXWFZhT
SxejE/MVoQTJmw0cqKCdRzuUBD5cWZc5ShBg3u4MvnEYdZbecynujnAI6j6mzhSiMt32OqAOueX0
8fq8oK6C1HuCjNhJUGZmWEMpz9ra4nLlTJAXYDt4l59UMXsMZqdJzAGiQgll7YaOKV8vXEfVegkB
URKiMr6/ECIgau/TmGZUziAVjtd5dRObLPiReuAj1pyPP/qN0HC4VJ1+sN9RbxHphI5IH7ihzr8u
ql0d31VPG9SkjurYV2XyBevYKJTfWUakW9JIkgtUXzEemr8EkEKaU0BCuT0+79ojG7JE9Q0nSl6W
7HZL3K6k/41QqyJ21aVqg45QyyqGJHAqPfKC1totWo9CXRkwdW2R0/YyZlNL90VO7NF9yzDYKEKJ
Rjo6lDRKtPVNNK9nkfXMf9z/keUaZzQbq5eIHVgAF/BaDQIvtoGswAm/sIcuMkM5jDGOj5mvH/NR
MSuonyKI6hVIkDXAoV6Q+G/Cmax8x5z5lDxHmgtZYyijmA/W+ozve5vzUL7RrNI//+K8ju9snKFL
sGxc4z1hvxJmXDhkyKOn1LV9n2r2YJuN/1Ipbq3/PONwCFFvt/SCU/c4hbboS9bm6EaXChcUgjz0
+dSu22qz/WRAbtfTWBZa1zhx1N2XU8a2/HRCfVDs0RBepVpQxtczZPHlf+8OfFi1dPMC5/v1NTUp
ZdacUs/luZDOQen+nA7qmlgyK4jy7aKF9OtAnzAulD32vxVnq7ogBDy1T96+ifvrrCNJoDKt1yJR
lX3tVHdqX63BvbwHAUhKL0r9Fo300brqbrk/5qISqa61pvpI0qk8wsj48j+CiHvm3WKohiDg+irS
mRyMCFRfHHtiFL/BdROvAVRpJroRF0SqHsrJi9maGgvr+UA3A/mgGDDI6K2nEpmer9eFnLrc5Fqy
W2w1BcbqruTP30Hj0nBzaHhSrWJhRA4AO4/6DPvgER3ic30beTzvGaPosLmPohdfoSjUXi/Da1NA
K1ohfkGfuSqNLueCSv5xX8D2K8CbKJQgRlztHxKw4b6SyPTNjNSbuYlVZXC9GqfaUnRLSrrufhCV
r9GgWTLOMrgUtRPnYOHwairw8S8isasYRxzozHzH6zBjAHeq+BxLUj7+wqfSATWj5YTJML8IFrjK
lM8mM034VjoNoeAB0zBNqmVxl5242aRNkN6CyL/BGXMtP0iFjmOoVd4lAHs05kd8lqPI9z20Pqg1
4DUL/v34i2iRNcZj+2mOa+7Hg+ajNZtDQhKhLYAzXZ0kS0n/LP14nR5uREas/8YRi0uaRgXmxLYZ
1VSyg2judzBoKjUgpzCzW3BwFt+Ir/dLC2tn14VOqC0qxBpAeEGkF8b0ZuEYIfvN9A+ZiWXC7XVY
KYGEv+ySmh/2XK7ugnpat6TsOIJ9tIbB6GRIU19YBU/ccC8Cc7NQ9bHeAaDZWy8BYmxwInwCeWtX
ecXt/NvCsii7q5DbfS6sxIuiM9q74lGGuaBSuTpxAh2UjE331KD6PlVcW885FXCwns2KHIJJKHbk
dAC41gdJWW5npsmjVRIzgQ0m50Ut1OrnVfsMZcPf+Uoz0w70K5BApsPPIHtgboRknOyTnKNVuxIP
ciI9Yin3KfYN8kcrc+O6WoIHTdIt9FpGmCGiejh/GBAL9zIyBGD8ErMAeEQngl4CH1DwK95+f6lD
XjRYPhiGCmw+G3H8YgEPjHOAmn8eX2CdX/F4Qx8eVYQj1C45ahFzg8/wiCdBZ7zIsoCjBemhUlZw
Sy/3O5su+WQ18bjHO+L0cE4XCDgJjCIbptC6/NAeYWX2elyg+LjyKJ2kRVf3cvCERGWR4ot1LLZV
pay7P8qwX+W2qWGTjIfAINgRhuvd8J8vkY0XN01sjeOUD2kBnSl4gc/LraRx5cXbkrwZx7lgH1nd
a/hpMKO35q56LBpNmykb37B/s5eiB75CozWLFWK7o824m9GVYo5Uf0ABUK4EV2FqyusOZUyX69Yj
9NU3567B24GOe1w9D2EpVIlu8IYCsuHfvM+CNe8evLldterozbpX+GoZIpc7H4lxdAXgINfdytAT
vKhrBhztVe0p+kFD6xvBOwslq8exFS3dwSpIjP4BoCs6EamYiIIhwIOPA1NdtRgyYfwo/6SzC+qE
lC8S/fYipiSKacOoY1pOSu8n+X/MOUvpEGezNnUhC3Moiqd6ABVXGqm727zz1DB99qavv/bJYTOV
JmYKRDn+aDerA9MRdEytouE0VwZDH7RzrDsz2WGsArfWM1jca5Q4VARcElxVWHzeUGp52sESV7Cv
ZkqlfkBZOkbD8rdNVS928/N8A+K94vweMQHfJL1//7KM835eZS9ESp2R5pGfCCBciTuTRCbO+Mfo
C0Abb2dRuCU92cVYqGx3cy83+iSykfDscbtloVR53ZydrekpX6TOZHTlqV/+o0h4JQvhQzuQ2DUg
v50iTPr/rbEZh6p7y/f8zxlwz8lZvx5DN5Yc3G4hCu6Ry9IlPMe8Obf0FdscUfzMCkowuYCPqcp6
PWkusB9WMhqVrTDNIFiPY2av4St1crZUpl0eeE2YhGtquiwm8COcNT54CrWGiNtoLu1yDL2g0JcM
XAn3gpaqp/niw28e8arEcUwoCjKaG1FhfDuK2RFn6JTpyJ4wSOaQ+mHtdCrEwpNV8hEVXj39ih+m
17IYY+9l9biOtSQq7pwtVnuLovaTA6ZdEDEn9s6efxVz4gSazcX5+cuLADdvaxKvSwLFx2yBmFRh
G1jSSF/Mi8V3aOzojj6LJ8KIBy4xd4qOqrbXdBdXn624Myk497PsRzs5kX5U1D6OrQoFNZ3VRhpp
wM8T7jxIfXDv50arhvHguB2qpqj3L0ONg97GoAffQdlKquG1PHP46myfe0EyyuhOF6xGjNo+akDe
UL9NwVeSrwdkp1cLD4PV2FT1Q2/ZVnRbDhEUZI8sX/FMtSKnBwSnXao/6+urb2bFUJnYACNW+CEn
NxooWMlt2f4jK1BwdjxMkcqPlIHPdH/KVqx0dG9SnqxYZc6eSj4UWCEDiH/vMVW7T0lCP0Pn0stP
p35p91sp9Hwk78LoutPNhxAlmxjluedmhLZlznzmatAelK0HyRFf8CcMr93ppPANes4AdUsjSNz1
GCOM6IdYK/dDVtj3gvxd/Wjj6YPY2Z+Q6BJoOw72Z8MKtTIScel3TvyDNTLYr6DGRXpsWMg7gPpy
3Vppj4XpLqqFSciM53uewIx6JxQuqZK6TPreVrQ4zweBNQ2cZTqGIzCAZ2jgmzXULi6Hymwj+44J
Gjt7Gfm6dzRUI9McqXT91zpitUk1RetRBPBO3+Nat/Hr3hfWM/smm9sMxF2aWq7F5yIj48kswb3F
0ukR3ZCz0VPYAuKyMlnxklJNlLCsEfG6HbtwyCrUz8I0ee8BWmowlKsSMjFJ1BDA482aoCW7rLaE
6zeEzwxtwSvjjkBSFTkwmdTj68LFk5Q4hE8ntV6MfqWuS0YG+XuVZDlHiVRiBr+UHWUG3eJDUkOX
KXNrdHJvYxFCS57HBRMYLTtznfslzxJLH0G3b8a45cStzr9VtE09AElH6bj1LUXalsjAVBM3VXX2
gQ4mEnqv7cYLmO4cLTbU0H5bxYqP+XLpWe0Wxzp+s7EvGceW60ZluVb3ZBjANf4VtAKdvTKiG3yA
6EsbkMMlKq/4p2mJoyDLrEWlI5eL8cVBV+zN7sclanijnoOUhpZ/uyFAaGfQwl8lW/19hwy0NV8+
wQtbHJNg8ZGj0EOIcSaMya5jSgxPUZSpLnszueupTRYeEMm/NORIbHkucZVhpTC5B3/arQthKw+y
qSkOX3umqcLm8RVYcFQXtFMzTKpBTGwuDsAo9PUDKLTw7A7+i6iW7DT+QlMi0ahij56HCjzJQpDd
mzTzm8GAFjRkr3MdDufO96vOvCeJamrFHEPyyZyAS8C9yqEVNVQfXmjtz5a13btAGaV0jHj14JIS
3iLaCHpPhFS6TD1hmGrQ0GkLLBL820JMgKg1lLP2ExoQ3m+umLGewBTa+4lvDOadE9YoGtVLxCiY
J5Xi1gEd2wvse6mpwhS6RAR23PFw7WcU4AN7B+kXtRYJetBnA0PIlWJrXspwQpe5uFZXeJoYJeCq
Vf/ibTRsgNenbqkk8DVsZlJIN9wEAfThUKhzwlQMJFvyqPR4PNiuBgDegbBUdKJjWLtF7f52WY6i
Oz2BZtPHHnEpVIQhmz3gZ5iR6E06NYaUVxr9iavKSh7Wb25HfgmVUfr/dCDIQUfQxenohBtQZd2P
z3kkLFNn7QO3mpjRQ3HFZk/4VO+a6h0/S3NH7Nw/venw1zYoZVUtXUUv30MrsLzceRF+kaRd6H/S
kW9Rtw7JNFOjhM3JXhziWjOP9G7HEl+FjzerRPaOpv4XNcvZs6tR96qLvCVw6O43rSMGIOFpe608
1pCyFdKmDfnjXoloGyMagPbhSNYsNSEuu7ByzXPY1Ruw9C5dz+e/2VtEhA4JhLCh37lkQPLhfGZC
zTwEDqh4KnKLU9wVjykbevD+fe5dUkiomx16BNTIy+sWyJw0BXzRGPcihdHcCPAQ/vCawIJn5ZgE
6TYryJoflFk7ZKIhk8Euy7PulWx2bnAocBEPrSIhc585FnTGzkoX7ZpgoVXXvMJxiOjq2Dz0pgIu
nCzi+1F3ZtO3mFzONDIzt/mlfpgNmP9X/wVwn7BmagS9L3xdnpPswlIsIwEOKolm3Mwg9uCjOn9u
rVVlXuColpTScGzK/dfLdSqfPO9gCIsdXSVDvVlodNKG10WExNDlh5aLZCkK6Cl5eevfjQI5iHSj
rRaeA3ywLDLAoiYtXhtBiFNGwcf1kdXOF+CBkKzo6PjMyIe4FvBuXDV8OFdZkucBWgogFL23BF1i
DUNKM2aZZ00QXBMuucX+Ua9Z+siUXTj4QW/dM82bi4iatZPnhYsr+cNiUUtno9O8l6JwGI9NZUwi
WYudEbubK+xo6FafPq+Z/Mf680J0f++mTl7LSW7YHrC3tTmCgC0SMKdtpaD26cx09004EfLs9e19
puqj+0yt2223hmdkohZyqLRJ65IB4n6rURT1OgPp4hq7H7dkNC4TW6Bk0mLVCE8YThZkc+YRNTal
PdzuCTymT8tCWaRefYpBql0QnAGzpDCnLFNQI1iM62xTZ8bx2tMbLBxFSQOPwAN4RyL3vyxAeFqV
4omj4MdoFbmpswXOXTRacm8B21oTTvbX+5CBv0zWwbnzsjYHU0xX0Z1UCfUf9OVtMEy/JDip4uS8
YHQeSPGY2NQFEKRKtVm38U3kYfrc1Q6/ooSgM9UbrXsKomblPQAdockchZmvpnCzq05l2XdGIs+H
nyFtvUAGC43WBSXFExRU1PknAPwuv/0afewXf8INs+loqlf7aexrkxDh5VB8Giot9QQuCnw3ji6F
/aRPgDmVV5KLYnmeXNKTw/TYRyEu56lR5GIBkHKORoav5pOwIGABauQrbFcaBv8wABrCBLj2CLr7
e+VwVsWQw0UvrjHm7+bYRktfLMGcJ0eHN/Z62Wyo9cQp91HW4asCspFovZUIIsf4uwgcR4CnAJAT
AjjhGJgLy95fh0Vvwl8xuJtosTxnHYw8QFkKJ7oM44ZhOgQm9aM3dNv0JnaT/BZ0HBoEjUHs45ie
yNGXln9ZoKjw8eK6rpeSp1Br5lRa8Rdv498pFBYNita7kQ5vcEV6pfECezXIOnDI5UlTzJGZ4hPj
QECM1OCvz/vpGGeup2QkC2/z/vvuKBWkkPUb8n09Y30s11uSYDm85UTmPhYLEELTQ4HMxqLqSvp4
z8VY9f42zJSgVv6ucX8CBpS3kxO1U0NGHm67N84WGzg6OPCccrrolitd38rZgosRCVtjX12k36go
X5HEkwUVNcUI9YDsiDAFh3aP9YVS06B/xMB+5iUpIA7PRg6TV+ZArCkgXGVq0pTNZ49wIqpzzW0K
ILnoLVlhH7oLU9gXj0U14NtEYD51tugMqNxXenfolBIKYLeita5UY6LffZL8MZIiz0DefZPkqpfk
18J65OCjZfj3YROe31AKYnB2gHva+/XApRTH0kyYW1TDUQpRcBLvmE/0ZFo692mHazA3tBN+v9vq
ZdLBHjaN/xXThxc2dEa0LHHLEGjjtNwnOhM+2dqbCqhVwfosWFp2im1kh8C/CasgKnJsMEvqQrFE
ouf+iry7Rdm5L0WHhvUGeoQtO+M6/Kx6eKJZ21YRcCNgMlaCCcDqTdBg9Z/rX/6conPRMbG8RZLb
o84Vu9UI9gltATrzg0ou56KqKKRRphO7Nzl1k69flZXoNugB646tzqdko0RhXngSBaQX0A8GNgI1
uD0+jzrUxv8zAIku4+OmK/nimim400HRWhptoNRdaKlwyOesGW42EQNDbE/eIXtaQ7wT4W0VvdUd
d2H0k2M3WntFu1bixzsLIqApF8s1GGMqo5fquTKoI/vv2sqRZ7awCX41H+MOJ4epEDhw45MXS2z3
iekRMvdZU9eJQcU+Xli16AY2v38Gni+k43DjDt5I8ZWz+UO+amfBlCOwoUAqjoBQWKODso5OnzgC
Us/slOkahjZZrMFVYF5lS3wi8mvgNZuae1wGRuIGxs6WL0afZvuPCaqydEWoWhbe/DPkcCRmbFZm
QjvA19S203nECHZymhYId8dwcyxP5GkzuuOQpXsOh9xCfDJOwxaGL+yeF2Og4ICWnF0AEtyR7yvE
jnof5kgfufaLo0AaRvVGooCQkT0wKm91wJcGuAvvAqzqVN8mYuZZA4Tn/OfPoaCySb0mUXDk8RXw
J7ThzC9gtzkpysDT8e580ko1hRmOkzcUn4FLNYW5Ii95W8DbocQcRZSlOrmBPbpRSmiY9v2pTk8f
pYSVNxJ9r3Ht6yV9D+3pVa7JmZ+scOMYlgYFpj9C9cq+HZ7bdMkL6tfNjklQLrqz36zzDcNgs11n
hfRfdhO4SQ4dBrgSkB1hEUknU390dXDBbuOLo8JpvF7RYantdJIy8yZrSbItmZQQa3meCvd9e/pE
MZzsPZOvOX5xGkTqzT4d74IKXRjApelOistWJaPiykGKEt1PNEG+8oOVUm0nxl3rbQiBMBdn60S/
iISUzCaImcUu/GdFTDfAQ9/GgzNPZu/3fVN/ZU+OPhArlmKLEEajVAX68Q/qy5E0/qvRJTPkar1q
O5OlR3QJsigAEMH3Vcv1bwC9WdfJNAVJRCbFNwfUZL8CUMzm6oCF1fbeOAhKeNZF39iLhm9r9G88
7IkGUnK9J9fE6Sgd1EE5YEsqTrx9rzP44tXnaSn7/Hxth2WKfqL2o7YhM1CndnOwsyBQdTY9k5G+
GOy77/EB4J6OEJDoOBTKuQr3LeIQi5xiaz9Vb6G7ZhYo/ikTSnOCgnaMuPy3ZnkoPcf+lkNqNWaH
bF4rp42OhexFx8rIL4gWQ5NAGd9lHxMueeMIgp1SrWjvrOYAlxhcEO4O002xuf63xMhllLUWg27F
J1mVXJGogggQdaiyFZ3CzazABT3M5QLfPXILD0JLlc3yuEawrHu8RMmlfH4jcx5cFq5zDw3ODWym
ZtutyK/sEK2Ouq2J6Y5f9i9q75u7qB96oOdOIRmJHhf7UpZfepq6WVlvmo2LK/47Fv8qmMmf/jHY
Me09qp4eezrCvAm+aicTWs7vjAtWUHFWWco567U4HxExljcgcOYgMBblgcjB/1XIjezj2rqMnPSy
GjXEhudWaiJEquOhqyWDL2k30HbvW/mVXucanc1XtU9YrvBjdpX0rWBO2BeGyLwvpEboNVUBK0kj
wF4USjJrCnLJm6So0P0WrF1kbGOMdLy6MdBpYndrG18oUTPNQvw21LRqyh/T/3vcdWobJIF0JEnj
aBPKI8F+hnxO36wERGayoUWIRXXBOlunJBZu+UVFPzsqPiYI9UFPA+301IGhF7Pznie/ADXVs+cQ
GvYJb4vgEDT3XCIXyOn54myIaq/r9kjlVUVG7S18JG6IlpAUWcIZEeLpuIdj04onnhC/lt3ajExh
L+id0PhMhXkw5lM09k9bnzEgHzhwZl6LiCZ8oNjXWI5HJPpsmg5F23K3S1UTo2I8s8qFJGvgvnsK
x6QTbcU1TowkXxpw2RDTNcsEqsrhSPGLq7VlL3LEUSoI41mq8f8aPcGCAUL9mhuFiOuxA6Yzw4Hx
SGfQSBtjfMk4RFWexu0EMT8S3N0X7GJA0B08QdNnUW66NylzniF/AtYgDA6dSJL7dwn4DA2oEAgR
eJaJ/RkJ44/4upDkyNFsG4HtReOCY45FAvJXT+PrNzgbiJOH+IsyRNB2S07yazXVc2Wl/Nz4Twin
+HfzuKdrNGcUC7T2+dAIm51QRyf1PAjxkNsWirpeAeO5dLF6GovkTB6cOH/NdQTXDNzgM+hXJnW0
9jnEgsVCGyA7I26juw/zen9aHgD5CFrEqOkzvNdiR21Ag4CjoShVZYGtULg6s0zS76CbF1vDDhFp
EAx/J4OwpSi6cH5FEGlZVKMQ9P5piV7TAhcbich1lsGK80+vZTc/qmutCT1Z7L/xcRuRkvZK8n3k
F5/0o2ho1a48bOb2QbU7bHaHpqKpD2y2ndCaDSKiAx8l3fJNn/gGwG3tFDbqo5PyYyjIPDhOBo/5
u4oPYRkEIZR5fu0wddOsUVv9tcJGpLPQYjWr+WYFt8MNPqybZUJ/7NaeqTM0HQSpDXcnA/ieZvUL
kq6aZdrhoDMhgPPEjSxqXTLXmeD6g7KOcoHrlfOyq0LkOKZsK00DCzplZIZJetzZhrWFMW1v50Hs
IiqZpYhES7y6obAlWJVhVMpzc013O20hCY0qeRbWN4tUcsq0+PtuRzVe1ecC+SYbAJzv7hhFPlCd
pBozlwyxuKZipEJrS0VaxLw2kkRDBpHAzfvQQpYhagzDSNqmdkv6T0WbQ+6kyNhYi+A0CpZquIc/
L+kjDYyNCb5dtH+m4SdfoK+sty6643l5HurPKjs7/WP7mF3EgcSK8x1RoaOQyY+0Ew56Ij7vBlVz
kjbnub4MgMnqlWIrmvmsW7yPIkEPGjBEo09/dFm0Nw2Wn3ppCQhR+rSJdAfjAPhtQx60d1qGl/Q9
tYFJKoIWeOuLmo6qTpLEGhhEHxmaXQBKwMAz3emEXGUeVMHJeIH6aclaArExDHKRxQ3+pdeEB/NW
NScI5bQOBd2HCB8ljfYZbTSJqK2oABc3CE8vQ6yA4doZOq3wwRHJM4UiX9HoVz5A6d3Nzp7B14RR
Fv2bnPditr6AwscEzWGK2Kp1sYPk/1rdE6sNqZPCEjFaKp2eiv6oGHUFmxtgKdBlFes36zrExf8k
WgSSwE0HSNvqZm35yH79WAaOalQMn7o+JWVf37yYfmnRFNlSPHJJdQ0ozzSnOGO6vI6Nc/yWfxeE
njjnRTGso/D7SxxbQOROoAA1Bh6ssJG4iB6Y28edSUp+eMfvdfp2Xq2invWabcyFLGpjMH3tb0YH
lQXDyoUgjTClDs2S/t8mPkZI/ORdUHArOE1e/DfsqHWwgEPZLilS0i/3Jh6AcJJg17USSXGjplSx
pcRQjGESLK2pKfAtqKyoxW8xyG/2V0w+XLtixV+6ewWcywpUMlH+bDIR0U2zAwL0e1St2QIy+ELC
hWcTOrgTX0U+J9QFfpeuZVnTHaGeek7GveDZhInA0CFfiu1TjcOUNdg0tacTFmBo3xeD+D6cZj1k
3+kEW+r50qwsF+zvdZi29rGCdjCkSxodAK0YsJfr5pR5Rqd+bx0i2Fr6Kg/DRLjQU0bjvqxbTJEp
jalbAzOz6ecMcGq+GannQ4Wf/X68Bo8ZzgmFDelLBuiN0Brv1Lnh4JBdyfLGKSLWXjXXm0VdWdRD
4MgLT8WoDCXyvLl4cY75Y64LnVxpJ1eKX8FXPXB5qRGGllfEFMvOqV3TeudmpK6vKt1sv631LHU1
ABsFa6KbfmlqaO0e/K0CNX3eimAHvZO9yyAmzEunUAR3Xxzgpf3BQ/TEvoLlTk9bGq/qGtxm0jXz
ezeQpL16B2IlVTMgeESQG4UDTQt9uG+2GLKFacrAVmH4Yw20krZMKOshT+B79kUOuHi51rSL9DVg
c3fCQ78gpd4IqY0dQp90hPUeV9/wC9okx9Om5AaqLpOfS7UpcDabTJdAVg7/niFTFKOKWxEQxVFN
QOzeZ3p1NjrMnKAkAABNESRN+2mdT73qXuZFW+wKbg0HmNQMMcN2/xxPbrQPP3oekVZ8YpjlpXnN
xF8FybG2UN2hOmdmS6LasjgFFedP1RbYBggIIaU5x5UqZH/akHEDiIQVxOeMKAPH6p9babfsqUM6
FrSJwxO3aZAhRH/c3K1HOBwGxyVtpdJRxSO0Co+heH04aJwGs6SUV3cDkI4DziwlCZFZZQDbfH3l
PjxUJ0X47W/h9F9dVHU6VRxYHLevx2szK3Y4F6cAp7QcCFkGklEo5tRuA0u5aX3oVBCLFIp5gguK
uEUKkGkqNiU32ebxEYdAjlpOuM3B6yXSWYooYIVKxcYsuXQIecJl/nXj8hxvvOMX4vwwjPfJgHvd
7gIhuiyO+0A/HQZDTljhHufGA1btGQQSQHY9QMR8EJZI+/cbk5FpBuUjSzu/78eQh8KKVUboNqYG
98xjxE2SMINvfTWie7ZTr9c8WGS8Fj0kTWddTF4ilni4e1/sui8EIb5TQHFYyJrgAwgKP/SstEuC
lU+z3mksbqGXqFMOk+guqGJy97KTa1/c0ZHAzr4ug07M/bTpFE1s8A4qt06QVqYtxAJFD0eJx/SP
actdXWQ4Fvqe4WX60JhBMn+ZCT6rNNGBOxDTqUbAtuEW8j2FJpwbMiU0y0fz/yh0SOa/7h9ojXsP
PRbnVgAVrVkZEZgoA3W/nsUnOc9XTKRltL1aU0tbgtc4TZT1OodnEOdsf1i5W9hBckvoc9X+lfq8
oxcktGzuG2i9m7Cm0U6sf4m058d4/BXgy96WiAoXSIPx6mVujKlpW+/21g866828O1C9+prG4Lvy
kq/em8zhVPB4+ib+nJxNwePehiQuFwIcn5uRNUkgdvIYfNS6+loSDeGr296a0SHuZxl2yn18cZBU
MJ8Tro8Tg7fdQrP36xN/Hly5h9qG/8sO4mN8Qa/wfD8O8lHJ2NXY4Mfg4eYNLIn+xfmKLAjG1HB6
l0GvQ7hHoZnzmCBNHJTjQf1VwWUkiDx/CMe5Kr+b4/kNjfvzmerXzkE3yVzsHja/8r2p6XPoD2EM
3hwVJdyA224GOcHr6bUOB5STcLLxjoh3+vkCMLM1fIYy2TUhyii11i0FLSd6e+AoMnRqhlLlypWC
rd/5U6JGFRZOw1GrWTsHK4APaHznQ/a5R4AZ1JVbVAw2FqhS8ZZ6nTD3LlHiw6gXv1qQybXrjeSQ
tL8R5m4/4B/qZozmzssy836QQ1BeUDfuOshl0sFsGJkaIBQylh1vPYjhNRQw7uUrmYpwqXQIK8tB
LAXaQPy7UKAG/G48bWi2PRLuL3NqdnCj6+Cw/NiaQqAW4J0xPvxdMYRgLXj5nNojpPzypB/87hrD
TFYpACk806sLWZVuCWH/JLJ5kqEJbnXQGREZj/rd5q8WS5ulujh0fwxmr//FzPMfLRjWIV73BNRz
UauTOG26UC1rpxcpqT4N5Bhv8w1XESbLdx9FlsocqgD57XjYs08rXkpJ49wAv2rdDOl6WTij38sV
nj4QutUoTRaMN3xr8JQhq4w1mR9GbJHhxPveG4fgRZcO36gcsc/3uy5XRXTnlHs7FVPTn0iIaZN/
GsHYTedXGi69cDMKsVG/siyduBZu26I60p69btrGnpXx1qGAidFnkOODH3byuayOBy6lyWGAgc+5
4Kk0usMv2+hvJP6uc26aJzyuTPV6fElhlme4Yw7TXCqLYGsgkcwZi0EKVIQHpn68x5gOk2XbmC8R
G/2c0vq5LGM2aAU/0M+0z6r9Ae0Ed4jPCLF7p7jKPEvqj8Kwl4DTwmJWPp5QlvgCFrLw4zgeWIUg
InsykIwSzSM3dmtupJjPSnS9nSmHJljxG1im79kukG+mITvnO1XuvfJd+l2CIy0H7L0jJ4YjIuDj
F4IbUC9rDmnZLNKe4m6RzCjHxaTdJamQnHmZvYW5cxdpDMh4o0A08lCycbKXPhO4BfacP2cxXkTb
ajvTdcqSiaoB5C1Z9UoUqklUMgu8FdpBRA8JwZfhC0joe8wam8oOZx3F1/EUiwUjwFFGYeDvHIxv
E2GS0cCjHfAdTqz5zxpZjZBWFK1UgUXdA7rJ3blPkkidkncwGc6XYWmsrD9fE+Ml5b6exJUo9THV
JKkYOZNwUgUNgudDMZy72vlKGcDXIZe+xbLYnF4uvxemB6kT83/cOdi6MBJ8x95sZS2qGJpbzNVv
r4w/emjLz42h4v2fZjPX8XilTTEIGRP+5UpuN/jwr8SCCL424yRHnZcMXMZeq2+A0tT2TcNJuo1s
DGpWguooYmzlbDyz7wIOEGSUfCp1jggZ0HjHHoVFHm2bm2Zk3LHgPOE46Uv36VlD/G9a8w8Og+V8
GzU0mq6Hx0EzC9iOt6u9uHdjES1FtCkGLCwEn2gGXO+uMvrSCVOcJb+VDbJVRoQqFORFQbQqnMWx
I/yygo/7QX1gJdD5NorIM9M4Y68pRVjDhtaUgC5NseRRYg+hFY5i/X5rvXH4hw1DZoBR7nw4OGcz
dVLseH4/yvEwnisBoE8XhFucSzrwV4EKyB/ZHQKRkYAVnoe4NrDghAIq+7xrM/CyA6ti+Xnhs4U3
vCVVh0CwPW2TSbFQhIdiBjJsXcCKLhb5gjzEwQ0vdLnciNdnjYu7gSamaj2KZ3NgMK8loTRMrgmC
0YakIN/jtVIQ/AWw8j3XONm8wyo2JGSG7Tqgqj5eBUV/zotr0faaF0gsWu22NibGwTZmSpLXTj71
vMrlCDKUAHtYNe9DW9eJP1GxiSFKBbIl8Mh+2dNKAQ9OjNKggo6oR4lKCicYbutGeMM2qpGJmh4p
1Xcsik7hxVwWvqgwuGj0yXgnrHytdLGU4Yr8lYXaItn7cEyBGcAj5umrGFURfUmUOUwYk5OKOy9U
TeeFS0eQVn1y1HCmwptnXT2ozTp+f+H+C/lrzOznJ6mzpHbCIqEZx12cIHRco5nh2z5Y1y2rZifN
h7k69FR39GEE8IAMNgHG9vbHb2h6ezLR8/QveOccmicfxgT9F6GZhDLTVV7SChy0POPQ9LXB6UeW
qPJFfCqICxWcAPXkbkkCoHHwqxA8DZBG5IjY39tvfVgdM5PmzmKi6mFaYG3uvBZSoFLx/iBGVUmI
NgGQvnsHRvegGNEL635TwcGfeUfIEGRy7iPU+QYtSOxnroMjoY/6EitkPfBFeA9qzURI+GudjDEw
OEmbTC3RCnlbwb8pjZRljbwpr5pxv9oVZBAv5RqxlPfs2ecmIZKqohGh8oOnabRbYRAWO2kiOkPt
MEJ7Tr3Ih7Hd/duQXzknX/QGFH3gi7GMx/oucZoIVom6ylwWuE3i0H4J/PHdQqkktGCmsoO5+STp
Sb0rWV6xvCZ/RayqzXgRIt4gUWMiYPiXcmYDYFFpYQj8a1b7k6qbjBkYaF7tWBtgA4Mf4IEFt4Su
zavXX62qVQqoLhBGUVFi6eFe5G9VqvnJPqj03EWkR1dQ2awbZYMPKieJY0wlPyJYgjqD5DPpYE2X
3xOFpMG8jtTXLrCYoP/aqRsbkUmRYYYhTjts/McJUnhpXpdW9wdxXMcQ09TPoIOcVqsGFfVj8POV
Gcj7lgQwXzDCI9gt60pedsEV27uBhNNqF7JolQI3fJ1mQfoffTYHw4qdSpC5Co3dQbzwjkOxyh1U
TPGtLGpDS2ZfadUV77HE4Df9WVjFXjiGv94ozmvulOSUKoFIaWUD/SQ9SmFRoEvQcnrVHdMp4/1a
4UuMx0QLifSKeJnUg7DsQCJRLKmhygvyO4UPmGJlvC/8VgmAghKcIX5JJ0/Zd6gCmLwnCEjbM6ZP
5YGkWSZNZxgW7EGgwATQV+WtZPCqifrqNGeyYLMHOIIV13wrq1ae2zWR/aAW86nqmr4tRQu1PuCx
ANaXjT7FMBLFRl7tn3F/j/xIaD90LBRGqpiTdCXu5fHlNwTvsHtv2e36B/4qgz12yxiNwgf7TAgo
bKpoEaasiTFM4vUKheA2+5cFRUN/Kod/5yt45L4viT2UpPif1gbscmoFGPBO6s9FoyHmHS7bRtPh
hl2MM0uUMPAcXS7B44gd+IGzSlWCzsz3mJt4qcsW/85L/3OrnwBBscXtRWLwk7ZTas27NqxbJUM6
7RGlXtb1PFbC5uc5AJSp1dQ/wwhaJovsLUg1BJPnxCIv+MT+cJit5lRB8LTcKMee8Xf+aDwQIXrq
lrTNDtc2B60PtcuWKoaXWXdEcyw9QMO9EJv6at95hqg3WW77ZX+xRyMTJyKjSm32rRcjhInC6SGw
9rTsIyO1ocr0yRqOH/yP9MdQWO9gKrhP7K4t511BN6/efWItSp4meQ9Wk/CjHk5dt93y61CPhjyW
galEluNrsV01xn5WTHmg37tETRtUIxBuYqqm/W3L2pW1ZSbO4+xHwpDEG7lSznh+iYp2VCHkp1/1
LgbuUyPmvNSeMrWC3uwsiQTcjc9/u72TTay7UyN+lRFw57AZvvRzjKRGdnGFJo9957a5wGZjJ0lu
i6mg4qg/dWJao1gLGW/QB3pXb6rw6UVSPmgq6N5XRrH3I4GSmZk9ruUF7dTZ3l1qGbJpdJRKvtWS
eDtDL/3oTnnhDm1OkI1YcqWvnq53zvmNLW5eNJJTFK9Agz21KFaHG6uxVD7JHM22Y5DL/8c4m/zz
IYrsT9AXP/j1V2xhk4iHD3IBmeNcrw6eaDoUTQ8eUp9s8MQtdoYgxVZsM6EoKfErvBWVHBHC5eAq
N1z50uDj/BbW39sMQJz7DBo/24R4GAapC8upgHsPKYzz7/luDzT9ZRpcF+Wks9ZoAHt6Mq7BELoK
wDODLtGnDYm75TZD4fftPDl2uZ7vXDpRXzW2Rf3Q7nHQwvtBIcPqD6IWIlWdm9LMsXHdDdZpLUDV
2Wh5YulrsayHOL2u+1aHOfxJYBE0SwXLaKsqD0/xdCb4FHkx6jjD9z5Ypu/H9oVksN8ojNajqcEW
wO7q8sUirb5J/6UBH70XCabNHQRBA50tnba1F9i2t7v0ZwmZdHHNJzCQHOWisJNtwJ3dBd8wK/OY
avw7HpjUYy6uSQYThY0w9E80jNftiIr5PO4ICcH1aZbGevWQNYMrNG7h7XSpFnqvbB33X9RlARRm
Snx8xee8BE5OuRAS4Y+V1GZuzrh5BtcnwMAbFlGz/WxFufr/VpUasTR+XAsDZrlt5Law/A+g0267
ZJpjNDsViR/1bXpdybaG6XXJ8v8wOMxYdjPcJAr+9PoachEjnQWVT6vpYDkAIFQNmBUmf9Eqq32s
XtOUl25yl38y3gPxMY/LvgC5gHVpj0J3aDqlYhDd2tFOVHmcfHB2z7z44yQpA+VjxG4EJq3SOBxi
uPnwpoSv9B4Vkx03yQZD1d8CMbfiwNUztfdt9DP8QFTFddfCWmZCMrY/hyZ7/IilA5GETMh1mMjT
6mpaAEp5xxTn+Fc55FXvW/oNnRcvOFnP2uUn3odv3aSxJ5o02sZ+KHpH7IrplD+9PixJVnAHTXQG
0XdVyhw5Cufwd5e94gIjmyZED/E84FAK/FAvb14HBwvj1eWVdJaNnkRo/pPuhTFrhfT4Xuxj8C/6
uYp86JFjsZ9SLgQPFZfZvJw3+luMp90S9lR5tI3O40ediQJUcFB43noAwI1xF6jAI153kb4F0Tmx
VVcJ8m7t2FLmEcB5+NvCaEx0yByajol6R2zYL/KyHW9aVbEpenwsDhSz5iQd77lHh1Jmbs0aKRCn
K/hszmqvmOdaDEAF5k8wtPx2+wWFj+W775Ng/6NO/pPSoJ5CubOtBPWoBs1hh1jGqnX8z7lO/gmr
wqG38ALDk8yDORnYn0hco21j+F4QCtM4RhSw3OKdMGJV1u3RWEtyv3OHcSzar/yathiX9LaOSdGH
uWXJl25orcR6haASiuRG4HPUGONgvQ6JyT6z1s+xAVG8iAN3HU4X5SUvJkLhLhXUYltslFWZCaA/
I8zlI9MUDgTJhtIRNymJbY4NiLHRJQ3LAykDDDjS14XvoN92XtVCALxUD3dFa0kMwzpExZQHlq8e
cHa8P9XkTduZ/54FVG6qNqu8vxULsovyJl4Bor6Iv5DOhQ45vfKaG6SC7A5+DybUVBqIJnsxa+q3
BjuG+Kcj54wlZbahy5usjeNO/O4iImPUCK2xiEaq/pRs40ai7ZQnTnEjAXgnlZ6vjbyPL3ZrVjwV
XTwHDZre6Z/nM8l2OZ4Qr+q77Ou0Wyjgn4/DLvKO2GdhU7I5nEktpRRrko9pKYRhC5x7H9QsjDdH
39qexLOza0NjzFSVj5cnCpr3DEKbwRGcetFX1Wj0Wsj7nCzzTkUVfuMmwiZBtTlw/8XkpeXkdvMM
s8v3mFdcdPQ/ZfifxmqE5WvySAW0eaSNp3PFd5pMNff2kMtaZ8iuwWP0+EzHgodkrM6DhDV+5B3K
cB53IKh24hLO8vlnuYN3VAs3Sf5q4ImNWSefvWWNYCemTVOMiYTbL+eViKH4AUQHfVTetxcvcF7s
jPjnLXCShsT54W/8L79Gi+bbGi2xXGWg5RM/RK8le7DoJBBo1vRhYtfLca6PAmE4eoS8AoSWQFC8
J8hKK6SYxkzG8If+FhZcm3z5PEYUpB1xlPh2hJuaYl0nFH7Kuc5MT+oEpHX34LXVm/h9NO+eXfDS
ZhubYaeb8JqjimIJw4Y1JCgpjFMX3PikG6ApDWRhoW6chZo7L8T36/VmMaEB0rmH3gLPnRvk0bgd
fK3DGUiR/CMqj4iNKBsijm5s1WyXRdynUgfkb5MvHxy0wOCG1ktg+BXJjJLDwkyTh3A20xbJ+Q+p
Ok4oR39IspCdBVSrYqaDeoTsGRYAjIAOOY6cwN7xKm7GG6sWBh/ZCBxjbuUxp44oT+ma8bx0FbMW
Z0LEPMv75873887dRdIwtMrPXgkGENeFrDuVoMEcsR2wausjr4s6opvUJTfvmMQ+xsISsMDUrglL
Hfgz7CNubH3K0IQ+E78w9r8EbSuJLZErJ/05x4WA2KxCyFutNbq6gRzp9ngQZEUbSSyTTh39fiUS
omrMjPUtOllWUHXjiDHw6kxqKpXf2CW1uDH2MNWUKOp+ia5uBQ2/2qasQ/rDA0f0EXP+JKq3jBXH
ElnorFiMozhuTBBLDv1HpyViWzBfOfarmRZy1wXU0PKjGhyKUK2ozaNLbtOllBcZAY5vudVIXiPS
I0NmlzdkNHX3Y30k81rZT4jU8Qu2f1yyCUP9w5GulfuSL8ByVjQ+1T7NcAPg9LvBLh28/XjZC0hv
Cq8rIby5aovqlDt856O3iTNC6Yf8ZlRu/fOmpJF1AsXqJt2Bm4X7qGKkz30okUcKDY+ng+dvFjGz
Dx4DBgGusHbCj165WLEX76/2cjsMcNiQx/3qiXR6ohV7wpW4YV1DGfFC+OSPQ+oNKUBrSXgP+LnF
5d5di7m7ihvK9bOY1YSIu/0J+taRF2oe345o7gnr3M5TKYvezse/7HOeQDePBW3j407hdcXprP4+
kBtRH9GUUiEfdn53WkGzvW3sAPjgApJ3TecV6h3rscvP47D0XC4rSD5lpmD/9Lqxa7X1PD++lRot
QB+ov2n00td8tiL2JLTO2Iz3oo7Mfo4fnwpt45T8GMFo3DrD7wpFKBc5lVUvoNrgzuEw25m/u5MR
OLXCuxYwxPUvpDKWwedjXsC6EESrmUkFcV85n2tXvzpR5aJZUX6BnrURCiHvYj2xJO6coJrTlHMu
WQuSjtR128Jdq7utiXgsHhPvKTOj8DutPYyEjR56oCld/fXh2I/RMPtCZikqU59zcQ60iUvH516x
+DiHnXJFODWoG2XxyV/kKWAjs5HfrybVfoBGiVUqLQAQwaWD3vomz9h5MO2lFMundYM7eyVSvcGA
jVpAGra7J6fBDMtdr5k54DF0qYYZtWg6IHla0/JpnWLC/zkuRpW/RVb381bhSF2nDawhIMm82RU2
W+qQqwgEf5425Iwti+U8Y4hamgMUowPEbPWh3tmNBUA7WLd0cpA4B6QEkJ0KG0lWaPGJmmZs9p/G
TJaM7koBN/XG4bmm9Ws/c1PbM5of7EmYUekF07xtcPombKhNGg15B6UoEAhizbbsxHPaC2FZJp8D
Rd5eUcjxj749n1ZKkfpV3FpcP1HjbOVKv1izl0FBO3gjbR8i4rj2JOHIKVQUStopALo/O/sNQfv3
HAe0QzIPT+QB60caGGBDM9Kg3qaBd+ra//DeMilxk7VloALOgkXqZGUCk9DDpRPv1zJEy1VjSfIe
dpMgGwMXHpQgnEqtqOqnSpTSOkfwTyXoGCO1Wvq5ByWVTNuRldsTh4VYyJqRg5uuwtqLiPETlGpq
O8KXn0x2m1NyiQ/oSkufTBmneMpqDzew1MPmzSQ7o/vOOsxRT7UxA8mtxxynPLMyWOBBXptuPbyr
sm1dPwrvI5hfgdn6vISPnoR6cYBw0kOWUJ8YZd61S7B8L3964siuwYVgVDp5+aRhhz1GSMgeDB13
UH3yjRFMK86+35AkR67me5w8o/xIi1H+coYy7aeMer4VPzZNMpwTcgcisg0l82bpVf/G0x1pGa8d
haGZ5/QvVgTy4dShQj+fPZzTbWfxC79EfFfyjATSr/K75XVCUfAk0bXR55190tSFGV1on2YmrTc/
yLCpW0P+N2NQ1cuCMcQVeXfE+vAbX8dxMy5DMFUipgdVFIbeBUK0POwbmliPPcbGF7Zl1G4hkDFM
DUE1/YmuGHuMd3pD5jVS6E2f30rbL0Mz9YCuYOO+jwZerIqv9zxbRXXA9FHMKBg2SdGczEBc85EN
xJzdoCqqFLhMk0Bz1J7VGsWVwsIXfNHP1ZfynjedGDyd+HlYDspA9USbpLsMrrGz+DDtRMCMdERq
Zob6+P4x6FS8LMJmf0l1yExp0IAax+poXuAiJkINQNQYLNSzNdYW3ogO9ZqkVMwvz0inygsK89hs
0vYZGIg2FXuadAF27hfa8Jd2C539G6hrwOp6ruD28ojpSHETeNKmu0m+VVVSK0E7kxVE2l/fIz3G
ypcQNlv2rQKDLCwa8m0KdTaWGhL3Rkje5In7vXWs7RSaMosjdRo3+ZEQONznBs6Re9mWV5NEgjBm
FFKr5Vc4N7XQ/PkpqbrI+8SgDpgHZpCVCbufVxutBBRBlipY2W0HbUjn14d0Zc1ANxUAyRGfqdtK
o3dqm5OmwlZAVOMqOxQdrZr1nke1iJruaBQqZ8aOPON/jUz+F+0g4QK9QwSsH0aq+vKlEkE5OVvd
ODoVL/VazsX3Ggu9YWlVhDhJZACIuPtz/m/EDkpuRkcZgUOA4jYPBvC/KqtW+j1ACrl+rf/Q/y+L
S5QtSWxV9yDq2N4Yw7Hwybdj4yzjNc/yRfOYmS5KZXbrx1cuymFwTFxvTkiBfUZyMe+qPkaVbPUg
v2YNB4MNPvLE0FJ0ub4tNQe0Lm8mtRnN8OBfdHxnGuymq1rqdR/8t8vOeYM1rXgfETCD3+/JH2pd
F5+NuMMlcqhSNxtT9H3GYyP7q4fE9y5WoWPTQdh/9BKNI6EQJoqCZzC9UNYAll9rDvP8y/+OAx22
eLuEuKCVHD9vRDKwVmRMSs9gWJ6zdjs2Su2YcgOvXZ32a4rwWZnaK6gEqszuDpiItitsm6D6PJLf
tQAbb46mgH/fvKMdlokvtQXGVZ6wALXIe6a7FUq13psI7kgLVsxFG+AGrouJ9FMOJOxd9nUmwh1Z
l+elzBgLSfAeD2D6ivDzjwhKD6lkwR/p/FcApUkWrDhzaumDkPP/DSTZmxkW7E/0aosLTXvtCvYA
8cbf0XSYyqZiW+hq/ZSL9FB2J4AdeCWgHo8c07seP6Mnjq56zknum7l3JJtwrwzvodNA84aSkpgL
D7jFTqJ0OHqNx9Vl9k+IEbNk3rLGdA1tE+pjPkuK30kcSUO++kgJblAz3xt2zPIMG+2TdPTtOzg3
kysayGVYTYQflu3x/TSaz4SW0KZD5KJxq2KQQScgL8kzxJiSSz+mfQS4X/VyI140+lX/VWHzkIpM
lad5MdLlWMNmfWlvFgWKTK2lEJEUX/meQM5qKN9LPPGCMOY6PM6fTSJEirAmRW7UGM0Wwhf71sLk
kFA8VeBhswhQEDO81vQa9fpzPA1N/xuoEQj6cz8pEcKFx9hHizN/dTtKSPp7l6EFwiWdyUE6h97Q
XH6RSQt88KCy1g5rXPAQ7UhLfFz9peooT1MCf32DNYR5wV4Sv8PtLQE6U5sCUlqL3sFAElZmN5pb
6TZSQ3StOJ4uBMpd92AWJEQsa1YJY212rPIzkNlarAKXUaVoS4asbxi2KKMX/8SlZ+Ku0AVnLZb2
j6x/0glmJ1Yguh4teKfUsuWObm7dtQt46DVDhSXQWSQeUuq/O/rRLX+fuxKIsJ6S/8N/tHCfHPdi
Yey+8xm1H/xQi2PL3LAU4SGPsYdPeDPraZDYafUiyy3eYNoj8q34O0yaco5dezO0FhqPAK3R6J2x
3qJFA0Mhw+Tbf0y2LMY8yOWGlodncYy1+ND6IOwB2sPQNsKGfu1PjjvitHAF1OGBHBUoOn8S1EP0
ZLGi6bCIIpFx0B0WX6koq35u6jr36/sxypH673H8ajaF6okQoscrmqtLuLpjlH4UMPt6qKZyOQkH
a2fslej+Xdr9kf0VY2z+rZo5LRaBprgUlT9LcWJBHy22zGFz5+HswSmhgZ+fE0MsupkQ/zlt3TRH
OkA2FXkMEqF215DSMyWwCfPmW8XHzo7O0+ZyOafkn6EuW0ShcZ9snQFaWNAiNqJpJhsmNwzbVOwX
l3HLC7bUYAhG+bpCFu3HpzEIf4ksUrSXnL8jcfBMGara8ZycjlQFCWYinVjeqve06OH1864qD4xj
wKoDIHMASWOk6CO7BGj31tNFfJ/xSdBPGFxnahMAzT39tHJBVL0MT1id4ysz4tA0kJSlQC2GA2++
Y6zMmGnv+bR/vL56uaSmczef8IWTBjxp3+KOnlZ5CtkFJTI8ROb8A83fWh46ssGfyz9aHy1hwT/A
yzqbyMkUusX9sNN36+KUO0y/VD96h6HXvK5MRY2+BN6P6XhM1CnRwMa+ky0MJY0dyH5BtTJ/eWKR
v0ashPcjxkhYmkkttON6K55OohkYr1tGn4tFddncBAgdn1nE1q15IDJdL9rxS+RJ+v5ZM4s+sA0/
BV3HJuGvq/yj2HI+km1vG7HKKC+xAoGTe0hKfqUTk9TIQNwKoUMf4pUevBacOFta56Cyt36HEW4o
kdLPZtiS3mCANQuzVuhHovYMZi6qtD4U2awndbHQxpTlqJ7AAFumFk/ZrDfrpiSdBfygC658F0R1
G5souMI0tN13v4Z0FtUFlqPTiRxsPNYQjO75ttE0cuqeBRMki8HJv7FHIpgWYfv4vbgfvzWudsqA
mOLVptcLfen/zxm9DrsFDrp2nfMKRGxY8cpB1TCR/9xW/KDSa7v8GOPk6K8B4kdQUftbPUEelDDX
LQdJQA/6r1S44dun89mQv9jK1za+ILN0gumRzCl4YM0Rq/wlD0r2jahbDQHyTD7k7PRK8gpNG2hE
pUZUmNopCJ3GbFaxBPYMEoO3TmQzzqkrm1Z9YPJGxXjt4acPmKbQX/y3ku4D3VHWELrJHO2mnmp8
TMWXxbIIkEiGFkyWF7FJnw7Eu7WxB+jYIO2kA/7mmxOeTbPeH6sL+IGgpEa1PqAEjsFEVzDl0N91
Skb5oPFhqBCcoRBU4BGNREVhjdSILP4QzyKvTnXUduJ2GBir1XjV9AOGqi8Z5AQc8Y0GvMaTZIXW
PoKWyP3g/TAmg8cnSs8S28ozDyuGeZe1jSGm6KwUqwdgXzjTKE2BkBWP6L5xBzdqS0zXuHuZs04z
Ak83VGo4fZMixFTshR79XgRiBYMIRI9YBrtEiGiDcRycDbsweunJLZ37oRXTWLe5e1mOKBP2wDQM
tjJCmC9GKY6xfn/LMkXBc63KQIYKxiUauBLfCZBN2+vbl4q08bAID6BteeZbsEezHOH4bENZYk+t
ouaSnHUNHOYUQ4/jd58igqb34WTIC43dFj36UcJ8dqKGbJMuQFOghFdyWsKQrSMgQdqZLVpz1TEB
ZTHpxN1IuvPLI/iZVn6O2a5TjPTKhtKF2pe7j15YybijJHbgzsmp/LhK4RDlDJyTs5KMDDlUN4nd
qUxed10q8VegNLXS7oSMPz59HaWphz/QB33DgwKJUeK9bfAR2H9SsSEB1XYNQw9QAyCpyvej391J
JcQE5mNLKq3T9azoMnsGJ89YLJmqPctuuwuugmFATsodqLc4aSK4+h8PtAwO8lYp8cs5s8o/xjvv
baQKWXy6nSJMokCYg2+F44ZXiwsU3Pd7cybhBi3kJbuuoEWAem7C8ATc1XUxH0/WvcK1JqqJ25Hr
/GsXUYYyGmT1kWytlE4H4qwVBXuuXygJmqIxc/30A5yrZjbMJFTetqIxllyY/91TLJdyTmJ3E/uV
iY+cIvA1DW2Y6qcumUms/W/BhYTw+JSw31jxe5W2PvQ5taWgr9mj9zvblSNGwLgg3agKGiZcv3YO
JgGJMwPfvOTcRaQN0O8yd7KPcUARgFMJD6BSmuRLa56d6DgL/yVK3Rx3IBDCQ8zbmQXNwa/+ZkG0
8hyOP7Cs6yIrAYwwYJAc84QtmgAFAyxrMhuOpleP+YiJoVbIKWSpueDF1Y19fVo5IUhRMUKE3JKK
gRwMiOfIk0HVK8KvAN2v+9s7P5pTv3Djy/Kuce9JOv1RAnzVY8YB9DVF3336xq/Dmtani3wcDy36
L0CLHnfkzaT2i3N6OOLoR7F/WrxdyEzv8YLg1aSFfmMqWai1jZ1t0D9Z2P8stFgHyvu0n6q1FZj0
jiUHDUQqjhKC4uHQ5e3RDLd01pnZIVAEus5ApfVDz/knKHVAwsxy+ooSVOx6s7A1uopSq8Dc5bun
XKj/uaZBF8t3aaBKqPTX5KPKaa08aW9/oy9rjhwxZph3w4rRqrgPy5fhNJlDX7MgkAQE/gohlaMX
tgQKKr3cnA1YVQ78CfVwl1P3louho8RbsVX1cCLYEUHC9x+b4yLc0RYDxKS+wfD4nvnTaZOrSWob
daKvKliikXQP2jYmWLQCoarfmRuAe5CcGde7BTKvBN3Ukb9HfxqWjHFKTbXpWG3B5evRsIOtJ88k
U6iTl5qfyB9g37M3PbQ9UJjBgozLSdhQtfGtwmAS4yCGtzPpcUcLPT7IIgjyz7hZxpJwfvE13pL+
xnboh0qA7alSm5MofLxbwtT5C7Qiklccf0Fwj5zw0bPMcL3H4ZqTUdx//ciepPJCXzufhKUpsHz/
N9MBF3e6zZDWGAY1pmVn+6UmklAi14sYzAIOA3Ka2szJOLVpOKifZI0jM80kurScB4Tm7hWu/6mr
ENIJYLG2gKWXXhiDukuOHOzpuHDtZswbTlzcAzFmqsvjaPxg9VOxKsXRsqVu7SdfK46cOFxqXneb
8eXpBbavgLGNTSlVgSCXOAej63piqcg+6gIEiQFYVxBIAsqUCshicoKu+XvCWiRq+oqcZAiCLuL2
CleY2PR8t7LMSAIzwnFM2cwuQWhLiU0tWRWiyN38ZQF4YaiPPX7jkYOmR/NoVspRUD8xTmLPJyhb
/SojIDZK4v/KwaW9q3hmfmXd9sZBHxVt1l8ui6TQc24A66+G8jj9JiPee+VGMGgFgLMKepM7GDWU
zBJ92eKZKbuXIi9ocjdilYvp5CZbjMj/ft0TKBKDgSGeI7I+cKsfm0oRWwY8nGRQX4yzGcD94h6W
Ugt7sc+YOm7WmLQvFRl3b8DEdUwTD8ttsuGRMXvJ2vOc/jiaKAYpoz52U9cQRNEaperwIVNJma5C
3JVBwl2TKDUmS/f+opoHp8ACUaMYKrhPMPa+nTLrc8TyTrNHE6cviEhxMfNth6oR3kleRtU4FiVZ
GAVD0EJU4Jvl7sz7VJSeklQ279rDv56dL0lRpTnkSIdiJvoKmhbI1RMIhECJjWm1Z/Ru7AQ5Q+rD
wsQPXuWdYGZLZXLqUoOqRgwNYLUz13eKxVzIfL5fGcMZ/z7ZmC3Irka2Uebu1xXn668vQ93Dm58E
0MF4EU6HLa8cry+gdhgGAOJHIb8LjGFgKQ76cZle5oK1Hzue1q7NBzfK6QXTmnQyNyLKprb+WPnv
qr+vvCwybRTRH3JAVFGsprZeCHEy9OEWaSMFdXXgeM8JwrB/Hpve3tghxN8bb/zuQjwjCqXXqNFm
eYA/tw+kqY2QZ96riSWgi9Xyw1n2izxUH9gWPkWNH4FozW3V1u/6h6WFeYI3hKeCAcP5DvUcnpks
jz2WN/a2NPv1J/IvaXd7HiDuMxKv5ttA+27Cqs5rrn8ola4aX5GMkloZsbsFMGgl5SdqjOIYmREs
SHwNtFJqoJOTPMFMtTzMCkQOmFMBNF3ekdcH1B8I7LHPVoanii+qDIrkaVhnUNeB0iZxUmhr0i9+
mbxZtJSl9rDQmuvI76JBHhFM69R9IC7UMeeb1WfQnR+5d9FY0SrqUhj+3Aei9ImFXCEh5XSATnqv
C36DVCYZWKaaEFdUGPMiC2I3kYaXV6vwSeIMz9ZXqbVxkH2lN0Bib/suqWXipQAcqNuAtjn6RvoA
Nh/imk+L91ZWwlTbHlcwQmQfVtweFuo0FaOwZEaN4hqnvM8zv6SbqxGBdDHS/tP0wD2TOO3XIPQ5
f4vDIEN5/JOCwCnHJ/aZ2SVOf/kPoRyW9EEO7lIM8F1mCLhLxGdH+cUBbuysv42E52HPZnyW0D63
y2NH28WiY7X8yZJF2tGlEUJo6rLn+aqNRHHM62udlOFqU0ChSS821N9hp4/23RPNYGSVoIwkxu+v
A+Hl24lJMKvbFyk9zH5vL4kRma+gnwwojjjqCDRx44bG6HRP966lu/EyZDDe1sEfHyJeOV0AcAx3
b7UM8n1N3sviGuXST3bBqi/9FjZNaPZ7CMui2L3sjtOSSbMYbhZUtm3OraYsi+LRPjdfucQgCO/K
RdFWwscAvfny0Jg+FDNQ0ddIeZz1fvVk4QCDr12ZisH6cVEtbpvaF4z+3wrgMG4gTsPT4PyK6X5v
U8/xlZDqqnU4OO9PmIeEHWEexSbMYFrlU8Qjqa9vAs0lSj9J4qv3rNRCLd/f7ygMuU4kw/48GFVG
oy+y0c/4o3CZecLlS0fB9Bq/cjydEl/9FwmF+NYElisbk/ilbWjIvOA3I6p87ZFeQCoXIz+IAPqw
7QeYNwVNeM3CAiUU7x5z6xXuq5uUPMLdLv5CvPQFowVZ7OcIhdLyesh+uQLKVKDzaphVZPrjpG/p
712dNYjOCGy8uUqwZd844S1JHFyZg2+Zn5t88j++2xOcj4/EeVM4Ax8GgorrOAq+6kFjrqc37+kn
WGX07EJOaBSx8EeZBJrufnMhkMPj3xHyMuzvVhgNUQVd0mDDpyQ3+qXvDl9lTVl5I5SISzHCg467
xjhzVCA/1ya2Isu5NPdHB9iGD26DmS2C71fsWqT9iJR0FkUc48xvvKHbPSjS07u/37h4EdfsyKW8
ls8NqzQ/UX+uBNYgFHfJcdtUvGkqBaIK46xpXSMGLgsVKDwRvccbwUkZLeC9uyJcdgrpTd43+fvy
JCHqQXtyJ8H8q0hn0YocKtx6iH3FeVnBAOAINzun7BiyTi6dze6rJpYqrS091JNnECbaWmLEULfn
7u92SUwbkbMVZJuEbwZcohuXeteB6KcMZvALhnx6rrKAiplW+FTlfWna91K3Vy+6ahGnmRBLYutR
ghcXrsQfx58S0M0FVxjLd+UxHh3kYo9B8lqdKTciFuilQh/Mbl9Mlc2Rz0+5fWVcHO2mpbOfhIAr
9Xfhm4y6CsYFcAZG/7Wb8oZiPN49n9eoQW5g/HUVLSPCPfbhRJrQyybIT9A0Pc76GdKmov1RzAfG
8CHZ6Z6z2t+PsO5S9d3nt3Q1ZcPsGoyijgCtIQjFceu1ED36fRGsO28ajwXbQDvfh4iIYpF/IWcv
wiH9aacwna0SrvjDGdMJR/sCNvOTkTI8zUFAbfyGp2g1HkZhI8Qjpvq5tFOERj9YpVRnpS+KVcmR
tSOPkN/diYOYr82yWoFEngJ9JdzQlCLN0G7NTKnilhgqsY6hS8kQbiSc7XXK2OdQZfdhAzAVpYjO
dRw7ChsodC0AvZkbCcR9MvP6/n1k8y/i2kxEpWEozURht90CrPoQgf718tp1KaDrqnXgLHPoQrWi
7FB7H06+gNHZKJ3LALvV+e9ctD30rsQ0bVuio63x74QXa+31ZUvW0N5uf4YRdLmPjciaWeKO5ybZ
5mfXnlWoVqF7qbIoErYYbt4vQuYfmTSJ9SLBzxfYuhsTfq4KyF+PMpePNRBJQqIAXcK+Pc1VDlyg
BGeWBo4WNPGxrTqm7uNRdlpqQeXT9fP6q+EjR5SAuhOz3APvRDKx2thtGGDPRHpt9UVBjw/LpMqE
q+vB7yo9gy47lT6foNC0FunZkW312kWNuTVaIFcrHWwuE60V+siSEqPcnHDZmfTIm+5lYgzrM1Ys
yox6GX5M7NtoZ9YjK4yu4E9hGfAc5/8tHPnUgNqL7xh2c3Meg9RZexmNp0UXkPQV8kAfniY/VBlA
2cm4MbW2ECdomUogt6wjT+FWpic/vjei1L8wmRNvr+uNJnK8Ta1NRPbynWI5a3zYMC4IslaIDF3H
J/OWQ2vRD7flgkhYHWzfDB0MYB2FYmiHintTscd66lHRwQHIojCOH/k0fsnsG0/0rmxBAIaM99mc
p46Ll/eZ15v1cThEt6sSNzwgY9f+6rElDLR/JKq1NkJplDPHL+vfe8xKo0vuOTjTzaIDmdnzySyY
10WeMzX1EHTazxWmDxpfTF2fMHRztd++/GlvqpqLxg1CKbGNlFFLGBqpZfzkIpNYCtqPSMCIIwBz
YoogkdGACmkFD+NlILtONHNkD+ZXO3K4MbwTFg/vlOxFwQOdC1Gw0bnXmHQeE7P1zBQVbb4E5fBq
FHCfDJTBQ4pv5cnipJnEf5Pg8uauAkVHo89F+NZyT0x3iQJjeYHwAzOmvw6NSGz5NHkMAHJB/6oz
ZXZMWNihGf3GQ0R6nritHFAjd9fwvDXEu3oRTFW1/R/zPwtd5/WzR62PJrK4v53h6wZXRJrOJ5Pz
wYdqUVLr/tb7F1o94sFH9bJRandIFeRsg2Mur2FK0+5/YDuvIa6XeLkEo7Kw07VTxvjA4aF2MOZ/
8vT2EPRT9qzI/zZFNV8KjskZK5s37NCfNrIJ7JmRqM5OlhZu/fIU7DGaqJkYH027TrEpxtV2y7p4
r4juAarXovORmzeLNt/ytsgn1AItbXrQ9MP+lUKt+PkC7kThpe4FKf/VMKC8eImxgWchD8HeZ0YN
DC9ysQY6Y257p/ks/EXGOizHNLV4QQ+yXX9byycN3PcPf1lKLgrz7XVFB1i7/XJ1iTykh2OLYsmt
7tfMEnar0muQYOP+BGeScShR7JE2ZooAmcs2FFPApoV5NX6mlGMgsnAf+1B1V/XiXcMvPtoBcqyH
I90aFuujYhJ7A8RJLCVCeBPUqrXIA2N5i8Hm3PDDtwkkD9Gm115beGmg7rlCMtEzJYmU2sjEx2CF
vIGY5i199YQDQivYUx9+bNkFDuEVmsFXMgPeetB/c79MWjhIltZ+5tdJaAUD+ImPn9+3BLKxEtMD
ocKY+2G7aOsLvk3yLqy2Xk2zV3/nUJTAbv0P70Q8ch444hlR/1e7InrKbJbYCyLqsVRrqzvR4ZhC
MNF7UAdro2BP2v1PdfN4UILyxcdIWY5cy5hLzw7Bnk1wLELC7yzDcXuWLuUK2j61HidkoHtvMD4y
kMyVcTvLLkJkBHfxPuvYHFMvQjhtKN1+2zl5UG5wMtwTTZaBaK0UVC44esbnIQHXIOBM68utRsUP
wDc4yLnrWJdBoTTML4/WrmpRFRBjmCWRoufexo7AYVf87sOVP8IhzSKmTOOwXAWxngRRE5kog8nM
S8KUaKOk0pBPC+ktkRp62b4viqqosGLMzfp8jgZ1R55v1JcI5aJRWHec1vniUDguJ0xfoKbjC6Ri
cyLwwEIapdqpUIr2M3UXb71wk9JdPgyFEEwr5+OpFAkb9AwUVr3g4d50Sm8zSrr/FN9AI9TsGy0b
GIu5i9ZGqV+a7yV/iqyugwpZr1vi0MpPU6fJdhqx8u+1Q24zyiDmO/kxvd3hVAzMWMAFm10Em+5J
6gExyGZuYQL+xVeRfboNHsAp9TOU2caQgRvhrAqq/FcZRpT1rmi2bl4JDJB/DaN+Lt1V8zXPi116
7IZ4JnY0WXM3yOklW8bWfmnnFKGyzr8ztbw34Ow8T1ZYhqoT6Y+npMzCIjw5hhn3idV042orIF71
KIuIxi3vwxTHkoAwWPkVYUIAzfUyvEBfkD957vOaEZxrqN5Q5noMO9fI3wW+qSN4OpfGgSQYazXO
QxZ4IKb2nrJhD9EjLmkjB4iPP35TPrVqiovFn+mswbBQtq4U7gXxuwUHybjESwwsMpz/2dmzcpYw
YKOirIRdvF6SlHSrGJQ77UxcIMijJcd/nvqlaqIYXiDKPt2CzABACQoSDKij00KT5s9ravxbBiv2
hxg4adKQFHK2RtBh2+XxrSnEr62NLRKLMhiF68XoLbQTpi5UzR1GG+oNItBfsK//OgnPqqE8h9TB
jTo356c3yIAV7MIR7kfYrPTSoxwwHIulA3tfgmyX/bGKArM1XfooQJbzzJ5AOAYpsb/nC901cW99
yfepjSL0muaV9Uxd1F/xlBDMl9gi1s0/zoz13nstJ0KMx89kgjjaPPvBjQGfPDkwSc3SGky8wkcE
SL/9cHTRd1vbkwWUtGmB9192mzbaubRgX2D074zZDzlpaDc8jXFc6C1t1BTOomr3ckMIinBQnYLX
Yw3KhJePgVaeZvbMHbpJ2HAaBm5Du0JuapSUdWlI+TN0LGPSLsliPgV5vZwlL4SaorBB8FU3182J
+dCrFxZ6zjlI7FAudPUGWpjmriSJOLLuVgzovdgQXynw/mtxgEKyc/R8fgdNNkMJ54LthEFeSarh
4VVWn5uHylHKNNFbsMnH6rUbeJXVcM77NI12erWKhP+fcmBQJ5igvhBsUalNDDE74Axzw1VDh55Q
/Jxu7NkWcgdgvJl//GG4vnlErvMVb3GQlfGZ3Lgbydj1xL4G3F7dnoMjPUErmN4ndKVhFqEdUOms
xwSSgdg34sNGoDHHvSq2vq2ItvvvwBYKnbPsS8PKuf5aMWHuXeZuZkhWVH8aJIWhNxbdbtUKbHYQ
ZV/3l8lU0c5KTaRAKpYLte1DnguZrrXmm/6xgRqA7GzIrcbnAhoMtYZli9oMI9+cslhWCXm2kwbb
+nDo4+JC4pei+x0BecFxGdPUZMDg7liHo33XhJRAQroQeedtwM6kqNBjn4mw7P3/ojPhCXDoRsIj
OwcTHBKqlebBlTeJo52f3yTG4OapC2c2FVRO91JWZDem0S+I6nlzBRPMxF1B+rox22HjrKgUCl3K
M8pJsy9jXdfN+eF7l6Ew8Y5BVBsPrxL605wkgpXHOL8yAgqG4Thu7h65Aauu3w9k06Wh12di7Zz9
k+9FfFxQN+1/KvZaKKh2t1pAAotQbwZRBc35pMEYEtQA+CMorGF3wWahBq2+gRxkBsCZguuHv9O4
diasNPk+/6WCIPMjirxsGaldyIaMlpsEbGjFOR0tQiYsuJR5fFoOg0AmyDY1HhQJhd5CTljcYwiI
NKQn2Z56xyyRCxVGZphucx2/7CzPa7GKNkgUEMYbtXiRMQ7Pn8KW/z2bU3CwYzt3umU9D1MpcrHV
nwwNy8PP/AyBlKATnzUmyqJyTT4qISo0W6B875JA4hFCaF4p8W0X7B/6o+cBsG3mtxeHjIHTZ+oh
B/B6ug7fhPOLMF3GDSBf+LcMYydgJZ+Vs+GCCeuIQCjOH7fhDtk50yJv6lxfiI1bjLGPhCju5aAP
gbh/QcE0FoIssMDB4nti3ukSqESCUGIOdBmBGWljU03LDffhGfRh5BCHLJZ7ZQ15P0Adza0wSIrt
zCEfbCKRKHyjT44KxT0VrF1GFAV3CKgdSJwSSiYp/ldBKQJ9DqrZ92vqlJtPb4b1S6cXtRtTVw6K
Cdf9rGr6uzpUKCBmWPTIpdsyVoCHK0Lf9W71EbrEf2VtVGVFDq0GUwL+gocHUFBGqjukwS7ZpoH9
idzi7m212If/B/03zfUjKsX1THx386VArsnWYzIGW4yD1mo4HIbWtviPVqLjq0PotVQt4ov9ZWVU
nelZINbrosjMvkxMoTXdUjCPBVrynd91bnOcv1GjqTV/RvIzJrNOVTXhy7/6EWQ7dP4FzfAjvYM0
wOnl+ExZNE08+i6Hgmw51XV5IROIh+/+wzsOnF+dLHbVbzGSjuF9tlIU2oQfz0K3n/5jhwgF/Ujf
mJ2aJDScI66LyRSkxu/xtrBymiOuJ9NpiqsXtK4Q5s2tixJMwpHG/ZHooRAIPt0CGL9Na98msUN6
m9i5dYQntxnH6nEZboz1lqm/ahkEpriaOhaiH2YNRQRBFdqP/4n8AINLr66nJcEM2O90iOR18rwG
2g9LfzmWab/kfqeyorphnmVMkfp2ht2x6GlT8Xm3B15c3c8gyQ+9ijoOEnpu6e4IhBSoeNTh1DPt
p1x4RE0jJ1lOnIXQ2hH6RhrqYsaDD9Zk0RIxEEAlWecPvjlEaTigj2oFbWFSy67UnBP1xhZ5dF1O
Anm5xkE6CgRE2Wk9sKxQBW4gWkFvkoZwltg5inQu6wmhMclBvDivZ8gTafQc+LVwNtp1y7AiyXUg
JKHfS24eWhd6sd41laauDbj4xUQ0aMHbtfu6PtAcaVgQw8o9TWsuMz6zCXoheN+XRxwaCfoCzZVb
DhwTP/C2xGuVlaJOcgx3PisMHVWVMCgmAAHUChwLODcDjKpIwJEixE9L33t13LAllQ/bZ99Z2EIJ
DCsk0QbizwhO0XMJWGeGk7utB7O8yBrVZF81fUoyyXUKzcJJufwveZmTLZmknsBoeNcdclpRCOlY
Y1f+L0qdbFd1JD+cgA0valbYM0bLlu7+eJ2n72KnX79aBNdCrVU16e6ZzZlvlOKsX3tUhpLR/Bem
XK049YSCz4+iijjHpMaWamO/nk0UztcqpnLsfu6kj0IAr0NVrxqAYwZtF+wAYZzzL81cyKoQVF18
exQySJtses+HfSTB1D6iYJ90E8UTmOShpVBCVnf2GAs4E4o4mYgX6iUAZw68rFWcBj6gjM9Xzcb8
VpYORarzbkL/QobKmcs/AZ4J3HCR+Gca+ovZ5xUeijy7uFKu6qlYHjrC6x9Y7h3ta9PDKREbttFM
UUNH6h1TAeM+CR9NUtSTRjMhhSAotm18x5jOE3T4/odfxBSznkOggTaHuMWtk/M6REKencDXCJXP
xK9OFybzNgbq0uRjLxkPh55l9S0ZIqw/fPNuUiMaii4UWSFNK0VU7cnCoEy4hna6vYaoektgOSW7
yRbYqwqOZ7qTruJ8Yheh33uuGN4ZOuPlLDyXBK+SgV0E7QRckKaaxkr+HKgtE0BcwUXmgplxzP0V
pulHJYCZMnHaVzpMnJIQCwBmbIvqbr1tTsA8k5wlHlk8t3eDEa2sR4iUEKCHx1JIb/RhveyEK4k1
3jV9KiBwUDd3yc9m+9CtRfW/CdaeHj6LemUyEfBPYpu89JXAXvnWn3hj3HvJ1gzqCb4Ay/rFRx2a
EmUZ4MqT1TvQM/iIfhHQaszzkS1GBB7UfVCfg8geWmIcyr3j8dhHx6z+vh5t0jcEnQ4qCrPt7KGM
3TtgKyhkbE0OUbeUgmGNYFunMcefPQ3kI+JvTxmLavezmUEtZHWfepHLe26Z8E6BQdmgjSt4KXJ0
bR4icUA/9YhYTYs5u9k+Rg3+hFCNeUiepL1WfIpDn8u7HUSgq+HUVwB/0j4j+ZlQtzq+dG+FVMRE
P0BwcguTPDv15s39tSJKUO2/Wn5Vpsxi9VYXaok9entXyRNOjYurfw2BTZJx5Vu7+ovyQ76dW/z/
ZhDImrnS+yiASTMO/0zshDMAWoYRT9CzPYcMBbj3dERbTVXTNuwOSgj72AnJ7sMzELqm4DPn06H+
nUgfE8ZIre2rtQe3kFl4jOfSmbZ9cq50fbEKkhRFSI6BnuxUgM3JjRciP8Sk1jYTiS1yPtZed6cy
n1SeDE/xxSFtGOQ6HO2EHNPME603Q9lV3r1CDnjvTXzESKjuBKCq4oe3tz2UEXDIdA+V1KJEoCw8
FtHXTSq9mdROkiKQCjZtq40dYI0TDSZzmNvi59FlOih5mCjf2a3uJLiUkp5KuXCwyvVgd2/Twwj7
L9rtIyqu4X/vUkdWhhX14r5NvZSGEsgy27bWqE0VoLPqunT61NQTioXbbXeKEMeGbI57K2dokiFR
d+UDBsYZD0abIMUzevIkx5D+t45V9dTq+vSzGKvyiq438Xhpc3J3wQhsKuJhENBbsbtngDczVxEP
BS1BU+Q/PffR51bXbMCuXjcIB52olfzSAl7ndOH3uE6CYpA7LvSCFzp+UKFkCaH60WOQzaKGxPN+
4LOyIHiu20wBt36GZl3gLkgi+C8S2d9Jc/ODTcx1QJ6WucGpHFjkaDKaf+JbO6R201M2GtRtn2Lk
QSUb1JYfKJt13Zb6SYWF3KjU4RyFm/eo8DEGyFKRbcciWFBQ1bXi2XSHsdZ4eg7XonUfOgYuqnTI
OpZwJwZjpXagVBWXaiuQEXPrgosTrAkM0COoBS61v3zSJqAxUUmkMG4r9HKH8lYRqGIIoeiKDgST
euqEo6hkHWaoz3KNh0Dy8OeSeSujg6UsZl7RZw9zajh1DlekdaeTh3+DCiSvbB4/sfzpzREhK8MP
LZWSnvB3gFhGQYUHx3zAfYGbKIPn+ttb0fAokeNC61DeLTnu/mhShzIKFZnfDl+oaVifG6XIUB9Y
cmG60Sr79VJTPe+VacMhzEZcuJYoYCjWxxeCKCdu0UDvZ8Wpq5Y2IY/JLGqKkwmxtvNF9nfKu3CX
3zVC4XjMoKR2oMBwQHHFfeByI52uFe/0ifYywKVceIuBU4xRgkKQP1dlqTQWB7eEjiI1TsfhKi/Q
4EiKXe5Zq8CLRCKn+cxfe/GCW8QRH2eNZQU3qeUO+WqwTUa1cq3zcFpiTHtU3lq7Ps9H9CPds6Uk
MB+MPviaU4omN9XxMybwwT4nczuSGOVkZ6WAVMV9phagYTdeFHto5zSP+1lq0bMYzV0l61QxyAtS
m/liHFMrH5DjjoLXfGpgydQZp2rK4fXON0f8McUBM9ETWWxH7jRCi6loHYkp1UtRqKZytnQxMRy6
Gc0d++1dHIiX5PLwEWM71viGL4y7qN5u1c3ab2TEZlaqek9J4T6XpYRxGxb9BYKdNRUhyD0I+qPp
2nW4suo/MXAnIEHSvjScinfV13xMOkFfRgWNsyaAQPQVIZos14JEsX2VC7siLKBWExEbKszHaeek
MZ+uD4YRH+Zz7ITNaLdR8goJQuZcfEpUZdHkMgqAEwxN6momnU0O80P5ka74JumvT4UQyve00LLH
s9cPGK3DxNMp/KpjK3uQUOwndcwIs9KKw9C5BOh4LqjOSKDvSuNZOxQZgZTJN6+7Ia6mS4zxgY9M
j553CNe2d7xDRxLKulU8D1EhA6beT8+6fJfoi1DyEfCaai3Uv5VUDBwv+jXnOiatRP2Qs2YE2opb
DzH00wKxs5qZ8J0iC1MeG77R8WNsWoPj6y1EtJ2php/Vpe3zKTGOh7BB1adtVriiC0RYNAGqDz3G
LW8qrWCazcjmhIVc19PV6bq4Og7gBuDrilcisapnxokbBxP2GbpOvIzD5/KZhjpKzbi8N/yBWzXt
4FoXgdItXRkJP0FYCI7TWpyEt0FpZkI3K5HIg/KiIY4jE/mv6iVgxzNtc2CwE+8dXnnhWAaWAhN/
fJC6RIxaRnPNyqVuBRs0aVCKkeuwscC4ExuAznEKISzsq0LMaStBxuC9LuWNCvbcjlPFYEXVrQvx
BzsKno53BXAOGznx6neBBbRyPWUeYTzeY+Nv+mtFH7BPs6eVgSIyjpMFyd9+bO95ciEwrPeGkoqZ
uCT0VXBiEwor+4h8lLtJXSSWpQdXaJJwc7hEyyLXbRAvW+ih5iL8X5ymfTBVTPFpF1VgQk4q4A3G
IdF6zetUqhgiDc8kVGqW1sr4izmNsTyU9KIPcQbmfaFa+4pt7HSs4ShsrpNAM03nscFsqpdcmChV
2gZl7z1jpHxY/Mkmrku0+GigGootke42rAyoc0Q8z0Gt/nglsKHLN9XZpX5DMLBcE4CU/2IQj9zK
X9D8i2tX1RDW+W9EO092r26bgyg1d8IpVteujw5tS1+oFQ4lgylZ1cWgMuVxwAs3QnL7O7TB2pcN
F3CJAjY8qU5dbXVuNnccmu5fhHbydA0jv+J2eHkKDIoLMSOmEsk0ZTJC84pA0p1+VZv+C6u+Pdfx
cawGyYw5bIGE9s0SJYwGcaEvcbc1BhgCSxxCrGk/sv8rB978Rw85l9oUbJNkU2ANaeOH8jl4B91+
X8sF+efKlYNnNrehtfXrxWEWKeonKaBdcQ+L2+/1K/4tCpeiyIBpifVdkRu8/5n0+JDOPpRWXJ5o
OHvZCxJ2Awk1ew2dkxpSNEyezJnipMDND6wZIxjgv/RXOs1NBX4cDWOCFbg3KA4CxQrJJd5xRa4Z
6U7uCchiqlBGIpi/+7wVJ+7Fl47LJl4RxxRpcqdUg/HITvgG8SFOhK+MnmzCxEBFtO2ly/KHuhoT
/ltr4lOLb/QTMnGLUflCdDxBsWpiIF4NfrVVI992zIj/DL/upmWYtxsXi+t4WhOCJU2xUfe5v1Bs
iDZi2WnHNjTQESysMxpnYvTPKiw0boMiJfmUALvVTy1QgKozJ8olUc07aGUIHnvB20QQv1SncmC0
/N+HJdxcjZMuSAOMgflgEP8Vu8mdUaQ8iJAPwYYy2hXuGCxkbgiSi6BF9N1GoU0QNXGPG26BiNLm
3m2M6JzTyd0UJ33CddGT0H4YO00I55/gSqudBG36eHdVwMR8LEetPydzeLUFOAAqevtqzL7N7am6
0qUmE8oAPGpj/UfmqxGuEsr7Y1HkLWviwt2TI8xFFUTBUqA0ZaypWHG3pgFHAVkz3frn/P+qhBW2
5t8qwlLeowrXrILjpyRbWdq16XFu/CRJLWk2r8j3RyMPYB5ztrQ/OdhRkEwIVBdS3uLYEmrXsSk7
iH8Sbb+vkuPtMXUqMq7n72rXFjYo+MTXPtaOIwhgQtrP82UCeKwuSzjrndIP9ogOkmJMbYvhqI6W
SEdjzXoAtyZ4oWfGhYLQwY6YssI3QmAGHdYiC5UrxaG//FSmCGXLg8TkTTwizAiZYRyQJ0IMRJ79
Eh+062EwGbg4frfrUPq6SYBOcyghBvDa+Ks4JuDcsKZqm7DU+9ItZ6fA1+SrM7q06xSBMK2tzx1S
HZnRk1UTliYSmO1KA21Z8KitXWd1IIRvUjMNj05+OwLk5RUOt1HxThrWBBghiLz/iGCYjjwEUxih
Ng4K8D/5VYAT2Kka3AYB10wCfF5K5El7SY695tGCMd3GtOUd9l0e+KVmur181qMqh7MWBJ7XQK6J
o3L+HyzBYHvXkMZx/rSGsGYWasC7DHdMzcTatpI1rOWDe2vv5nxKZPl9gYzmwBM5KSHr5yhSwrR3
DZrAM7RS5OXR4o1oatHucGiQek+9rlLuS6nFL4+3ZpEogn3dyeEGubQYdlhPmLMLQS041/P/8dqs
H1oS5y0Hx+51sRSU0T9jHLwH4hI2MPvZnUbc9v83W3akZpyn1OdjL0rA0zw9t/+PxZ1WXKbw9gnr
gfCiY03ujQSWDr7mBRR8XUg2gAQ9OFPB5MPOA0Du/PPL/itiiciWIwlo/2ovbxhWwrIGsL7z5oNX
X+qw+j0GXPUrAr2Dvc5ZuXUZP2h4zh7qiL9OQVR5ZdFYBpy1MSqGJ9BdmoupfT9R9/XjKwGw/Wb4
9S8j9AC2Vs8zc27Jh03KDVUsmfPAcU19uVHGMxnQVpdzXtIpi+o2DKF/4V40FxK95ZP41CfJga0J
Z8wA5KCKj6y4kpTvoSOmybJ3pADIbhBQJmpbUjNMdtmkNcQIKE/gbkS4Wj4rs8Fvh7Nh8/jiZWtQ
QXWlIldxfFuim7jbOVoKbyw3N5FAvx4b+FNVErbk6TPdr2w9aZ4rxTIn8O8E96rClvfJ/UtyNE3b
2d5IBKVrHoDgXS4L3thKSU5A2xjq63seqKYSePsmNzx6+VY9Tm77LUIsf67QJ5e8Cu1MO6Q18G+d
KQTDDSQ9Py8otuVltREQ0dzN5L7ynIMbTyVq9/DxyKS0O4yyrkwcs7XVUi2TtgAtvKuDe4YZr0Mj
8Jk+OYTUoA/Mu4N6wci469lVQ32IYghv19oUzhgO+oThLFskJz2Bf56cjK/DLb0SZRf5SjFvB/rP
LMu0RX9nKv83vTYTgkV09Ye0TCY9Lb4KEJ05D9qmBoP8Xl4Wf0ViF+8BZFw7b+G0QxltXQlKxyWe
P9ZKYl/xhT7w3AbPdn3WNoqQHPDnulviTkG1MK0Kd5ZKEvFV0VliqTNX+38Y+hEreCj1HUymWLtj
G9jImfECzN5IDS/knOsbNrxNmHTKrggY6hOHX4Q1xpkOltn1ikt3DzNpM/NOw37+ySxWP35V7G8Z
vlnmQY/bOCHBrO78swVpLLhAQJifOP22tDn0LVMI9OCwHUlpmF304EhaQSq5qlEgWdsf9uj5nJmq
5m8ySYW0Yra0KK87H7eKoEgBRMf1BCGR+a1Ya3D2TZD38M99Kc32BVl3B0KC6Td2CmGFEb1A94/n
xMFQhuoErrUYaOoDzb+W+VkmNHz2SaE/JSp1oXbJWNKt2IsEei5BHF5ttP5VVwMh8ds7ZDZeULB5
MMSLgB7ZGwrQdQyx1C+OgnEoWWgRF59SR6811isvW3AURNgjiguwc7emL4Tepy4Yu/PZA8fxijhl
cBe5BXmP7/kOO3o2DwrQ5EJ1IolmgHsuRlfE/XdQB4WYFGOLd1gN/NJQ4b96OE+kzyEx/H4mgSic
d2vJxWD+j13rwDfYN0X6Fml7qfIsld9xM+sDPm9PNmA1UZmgumxM2WhRdJMJPPxFZAmSFyZDQSJ8
00z/Kww4xpeq3Dmnxg8DkLkC8bhu4r2p6HBz/2XQjiBhmA6ArgcopNo8svAW2WquWrkZkBCRYvE/
l30xGpU3gKDSUMiI3pqqAf6boPZbMT4JGbmkO5wifIYUqzk9OFMaZkVe8sCKAmgOvmlPFqw3R826
XX9CYCpuvgmpJm0SzaLAtmSQY8iOw3eHnqutccupT7C0rjYeUuG0UOt7Ws18LkPPyeYrHpL2EDnO
xtymPY98RfYCZR5a50kWibSWHgIJUWynsYGYe5NF/771xG2M1/O4wVXAczTi1c0xDSkARDh4yMFD
m2Zj1YbTAtrZ/aMcWeXdseWaWV37I7q3pNybJANwELCt/IFvH/aeYs2UheDOfU+0XaYsP9F2ueqv
f6rV7JBzcavBEoFzQiv4gnY/GWIXcfEtlOW7wMNVrbgfUAz42As7KYANjBMBH4zNwsyU+E6TTSwM
/ZnRvD8og6O+Lv0RXcOy+V73cXMyHN/KMSbdrdFcmQErKqFaKa6I2a0zUUqwGbq/vlGf3OlntuRa
U0zsclpWdgvOhYP+AplTTx5z1TrgCe7NUQsxyXEy2BCLJPGEvtlpa1en3ED4jtAGXeyn7TK8gvHR
C5sIZ7BZwyF5n7tgJTWu+1/vCd+Tt3rDTRSTxp4D7ENW2fnaoUNVQFOmPxuE/RetjzZvK7i0zIj8
3cWppmN078VYKfmMpXoJgSSxCpZqpN1PXbGMnI4rdSSUXHniaWSkJOJFtsSct3O8x55/ZgOKx2EH
1ujIahKZSQZ3GeCIgNKv4rHcUHRiB0tMlMJpSDY5B3XCeh9MGve1xyS2X+55rBxJaTqv9ng5XPRr
/aqOmVzBheLDUZc86fQpuMi6BPTqeZIZSpmrJkhtPZySlCAM5RNHPHXkQShISUrN3u9QHs3gWPpb
eL4l8tFeAZPKgRj7aGPRPIPrr8Dz2BMeSvS7HuF0zKIZV4aoHbQFHpScOqeZenNyRXGMcgTM4+QM
uGSeDnlmZTG/gYw+vdp4eKYLXxusJ3sGIAUN6386oSgt6eRe8lJc+4FSr+TXCBo73g50/+oABuME
tiYjdlf4OAr9jH0hh6WM40JR61hdb05QEYJOYep0sdYWr59uoZxWJNPtlORxILlQwkMmXtnfw7oV
r1d3rOR2wA1vtaOIJqo/AahtW4KbE8sJlRJWVnaqHq1Q2uOmqPw6i+uBFixPKdQE619tKNCdroKV
9j99xhuu4426nPYMhmy6oOKP6VM4szCpj05qleyom1EcIyuAOKD2Yh3isqr4phmf5dHceLPz3AJK
YE3BvmloBeqRg1IjqqNrjFw5X2pQjy6xYzM3Af8TiFZS1KF+dAqxl4gaGtOFm9Jb6Xa1t+BU1pWz
jsLNujRKEMXDNEqIhLv/uOmBLe8SGuCCL5g3lCBJcAqPmalqx79q3DCQpuPBUjBXyUdjgAcyh66E
NljwrzAHPrUgoxy79++2j23VN+FkrRmkx6O9PFznIhNQTJMfGnS7auXiceF/qvCU9ttl3hvqv7tu
RBa1sJjNXnojWJzFcN3PPLSUO0xGIAYQ0Cb1N6JC+aVU9knog75PXFZeCSIAJq4H83Nt7F+ScVyC
vveeUk1ZhSAkAQP+i+QtBA9K0qt4FP9ju3a5BvemCUikvoSDldDq+jwpyBOgV13mG98M04yZJEzV
6s5G6gvARYY4KxYyybLlnaDhFzvaKr03FdpFfHAmhkA3I6Q6NxEFyI+7pk3siL7m+7ZnBYmN19MT
sVcWothIpFLw0BRJYCmmbMPINYbbei0iLvFc6cjuGBbzWF8mQtlMZMwAGGTgWPhNqgAkv1QYGoXM
yJNRWT5Cv0T1hIx8uWa+gEsMynfSr03FMD20c8q56uNJZWftJQ6ESzb053LjgJk0mwWLPMGG5r/5
HV0wDT16xLeVT1vccMZosZqL9MIpqMQMo6k7B2uUFFM6TLB4C9B+zSD2AD9wH7gnMn82DIn2qrKX
KBuUAFL4up/8gK7TgQZDOYDdZ4dbb8QbDONGqzqOLkwJ5DyDuvQ6F1S+r9n9S/ul1pALxfy4+/5p
8WjmMl+r3Y0Olk1ucqpzwktnvgeGh6e9wNenU8D/fSGiwVSUgnlbJiWVEVM574wMo72FTORvIfqY
9L2zhr602nEV0yeNjFVRmyG+eSkACRuwxD8dXFzz8sEOk9C1YboxdUr3dMuwBUdtkzlUvRY1trCl
FdvJCO+EeGNvOZ9/UdhFbgqPVTS66LUG3Y5sRDOhyoHT+fi5WIIOR0UZk9mGchSkLWk9vI+WwKJ+
l7umvE7LniMAVb4P88HBxh1/Qr8cA4JeufbSzWwEmyEWDgc1yPrzB8bzAC5rwL2D3/xNQl3lH1DK
xGu5rdPek+PPBAAPfsa/qVuC70G1ZOVmOVnsJ3HL957/lzf5NsVmmRWbKYAnttNL5bzEk38YC90J
LG1XhwPTsUxu0SdZvFVQAs2pswlf1ybfRV1KISW+mKr41rlphgIlr3jBI6NoRHVPTCWOnhqu+LEX
jZVOoonhj+2dNDY1NdI7M6aTyO7GSv8AXi+BHfzCzTTRul2bpVgz5NiA78ehjmDCK/vGByfh7ZIr
nMQpKF1ey9KiN08TbVYyhg/djg40t1RNQk7oyG6rf3ldOohecIK+afEN8x742JhhxuQM3JEczGG/
VPmDCYpH30gnF4PKt6rjLtuzjNkirBehOZWD33Qb3Gxmb4b9kUpPBuukwwnZfIRKPNX1+1Jy5ALo
pkvZj/m75EhWKoKF6iamFHlKrQ9ubHx+m5/JWyfw3AQ07nCXyeA820Q/3QwcQg65uBjzYIDb+CS5
8/9JBMuVNMw5PRuAWKEwvyvu21ldy4meiCo+5jNtAcZH0kdwlZPwadusXAZeAehkM44oaC3vGDwy
gucT3RJXEzcN7kWkvEiAYAGcZcjqvYM3F2xK48gOzqsNgxv5tiRTITys1DaSmOSc00POql9mL/Wn
IlQ+35vMmTZyQsfKaO0PRiJlpcAe7WHfotzC4065yYS4SVmKG9xrzAURyV+FfZozS3RhYMNQs1mM
sl3KXm679Y+LzwT4Wr139BvQhwE5MJlY+UxO3waqf9sevBFGfWiDuadhCASQogbaUP5zoUl4IUov
LpVlHd2VeXsDcuk4rzNV4mRKdbDvIOXR4xhJT9sigw2HcwS2CLhOIb9CCMtF0RRmsgAcVD0q7keQ
98sJtHuhTp3bHbKVWTSLOFkV+VWifA3dg8n+nXKl3nxYPLwCYGCtGpI9g1E0y6rhWRZlkzfc4V/g
rwdz3g3ZvDxxUGsrDysE+rcOyb5vsdnAHz4gbnZuDRQ37ic6S03sIjh0610r3ej93IquPn41Xz9O
29yz+fM1YVnEy7gJAB4WeJHBOUO7OaG77sdK0ICjWAZqQN2i+0m3DMNsO1/xsKjskIrWdeYbNIGi
1H1ZX/plXl1CK24/iC+K4rwjUZ1BROeNv7TVQ7E851BglnJzo+hm5vgHNYWUe8ivPRePGA7fsF3g
s2YmzsmXUWQCgD0k/cr2PzoAa1r2c3VwubZEPEtNUEuMJkLTthZP2I+CHwsuk6tT4g5zUkfP5ayw
qhuRAwyDcfTR0BAg1kvfZHW7ehKt7QI0LQiDzXI6ErjpTG8GBBDo3xMZKG8WpfCey8LM7G5e0LOA
GEbLUPAKP76iR6xIYtzWYDZZYqLVGDrmsVgzdqUcWZx4w9EZo57mrzxjgofWtJfMYIJz9fcE2/aN
Xz7ejcELibdNNg/y2KdxS/o+P7uZIxpipsWkuCWsSBhWjqqHiRsXqjeq4xeSwfzgu6btUZpf024N
0LW3HsD4XRFmx3l2N60xAVvXYqLTJO/KVobnh94QmtM3fQodnLY9RiKgMPNF7z6hdD+2SMmFuq2z
Hxms3spZ/jEkxJ6XnbVYp+i6b0ITJtv025loHMBcJGYMjg1CWsgZj2Mz2JdLGZAfg/lUTnzpX151
ATLt+au/322heU0hLu1Cw7Pe/cKNG96OQEwd21/WW6nO9KpsT+LHQ7KYnAnxSxJnyOeR+iluobGG
NMfEQM8VwgHBytmCa1aHoRKbJNj04/3TzJ6F3xQyoHeSfDHePZaGBrdSjgZ2rWwU0ylswKhxQrEi
NiZq6gJ3u5bG2xAsbjr1ftuxvFJoVn1sg5hmaivV5JsoWstmrbtUrHSYIzfgtBqUDpk1rgzmfrTT
YrzXSXNHlOxu12N9aQQgHdZLkITPRStKl/FtODYgU79mn+mSTWBP+pNJrAzHwc7NJCL+ARy81uaR
JNB0GONeN4jpkk5eVSYfOss2Vdi7FO5AOXzWvgaiT+uSEJWcqNiagA4ZQfYb8lwtUL0Hs0yvtj5o
QMg+LKDaLfPuaFA07w6/SodXm5/cTocSwWV295fzG22tDbMrvsuTh6ehv8Zu/PLzDhqyA7RpyPHz
yWr7P7mIOapArWPCe63mXqEID4SA97emx9exn1ZvzngNga+Fm8bDQ1ir8KjLTFw09EEjVcIfWxvs
FNHslu/fn5IMLWzuroYz4u2W0p6FtPbjtLob8v9m8EyhxT7vc6GCjbdeugCKXrmkWncmsD512Y1w
UdprYrrL4H7qA0cUQwhGOt2ikoZ8gHRyStS+U1qpMV8N0Z7Jynf+hMFKMu5sySbGntp8KXdCaBJp
CAaXSDHXysg8pxSdaNvsED9bHicL+fVnyUpG50+aYIkRqjBzfjoifg9RElm+6of+R3cPBbMtjrCv
5CB1JV250RsaEopXFtApg0Kz/8LIeikGFLHEkZ6cCZ3lerkIxpfEC+RNJLN3U+GX3btlJl0L+nb2
l0G7y5MT4Hzbo0RmhZMGmMJYyr1EG6ztkZbNPP+FcsagEapTKpFX5jglUSozUsowrA5b9qMiaLwd
dEIkMUXZzj6k5QveJOtS74absvSWxEDavi/Eq2rWBfsk72Ko8RktgohvtfqlaD6xAjSmYDRVLnhc
NCl+0GEeJNbgiSMpYf4BXus9q2lLu1QzbQPgHp386A3wUtLhDeZczKY17mYIbZbtmcAyCoVAzw4G
DFTtTXaExw5HqnZgE+ByW1Hlud4bmUd5h8SPttU1d8bCXf9itvWpmCHtu7EGhh7DNnDVfG0paTEt
Fe4OYvoRoUEF3LuLxcgiULmusVBF6+WXUf2mAiVaTg0G6s/xvqf/ma8v2qh0PlFdzOOzXxcOoyrF
kbsTkR1tcR+XITp5i6JW4jT4hpIn8Iprm8/+ZQSYF36UdArmJj5rvp4b4yPgYSdsCsBvRBPJgPYv
b6ie2A/pAQEipA90cjhARk9npuzg0MORV6c1xLaaxWZ2NjbR700xhZc/tN6ZQO9NuOT/FC6SEQ/h
QQj0JainqcU+cwT8Z7g87cscHPE7XaqGVokUgsow3M1oX7swofYyy/IloK0imoCtTU3TpYMZ7nlZ
ozx52C8f3YQ9+PqADaTzhV9tG6ibivbZdVRgI9rT/QaM0hV7cp7IrKITRILaxnsNGrNP41l0/V8s
7WXjcRy1GvsaqXyCySYb3tyJz/Sk5823mxGFd9uM1MLwSNeDBr6UlQBwt4Qg+1brpmwsXau5I2Cq
Q6SrJOW7NMGgHRQ1t9orVMOa8YRnnZPCovW66U19sLRhesYOBrK1H8/CH7WECKhdO/nnOarBXwDn
8Yt6MTmtJlbVMlDjfzE32Ud93EuHo81+7Excon/47L4u/ec6tSv2R7j7Md3LG72UNUo4EBAykKd1
mV93mb5eUWRcSCqb8dRnvLy4IoBUhcbOXe2BYZySCEJjGsYSX8PcUtAzs/QjQBNubpvFpS0qhdaq
kdVAS36B8SWGXXGYKsSePrVUIXOo5H4tUzugaxyU49Pi505QHCaoW7/cDV9TLv0GLTCv4z4wXNZm
rtKbeyvR7J+Pk/mpxj4jAPaGdGWWNFg2zE94oc07NMqW5zazUBu+8HjbgB7OqpVoW4qqT0W5QIuJ
Yekz4GYWGz+o75VpLty7GoIc2svD2GJgzIT+3U1tZ0cj0vl1s4mg9V/LaRGgz2pjgvyYiYy9gmZ8
4WYBIVXdjaQMtrHoNsmmDWqfRntG59M45JAJkrJN5mjiUbSUzc7BrUVgM3yynKHuGEHRYZcR93ny
Iqf1wkP+F6Zc1P7wJCBEONXlJdgX7lMqIC4Rn8lgD/OzEI7rjPLe+DLhFmOGc/xTY9cINulQWAOm
0zwE2zfwQH0XRj8c0RMjTpLBECREb9BorNR0Wqx3YBt16XDc9bnpP6l08L2Fo0uzOhqc3TrQXnaQ
9wexh53ujf5gyL5yt4tT33leJZ5+iExOaoB6WIRckVxyB8T9vGWTmLAbjA/5RNLgcRphN+amPZ27
8oGtGZKd7jN7FeMnfi17z7+aEk+3cYNAQTvMDH4YQOIyOeiAeT/fo5koo4xR3ixrZEoST8Zpohj4
Xdz+xINs+jcFSCHNypREG1Vqe6Z5CQ1f+aSjPEIy/xfLOnw4AOa2TJKm2EPDnQY31Djt1BJludqS
7ELGU/gMT0q0UCYKlDIxQuovIhyMI3jWJ58E5vf8M0fDPghP6OtrOc+oR6Go7waoqfhcdVYuAdAS
TSpLKe+dATOHMSRVmMeraRRZKWUS3asQxMIxFae9co3UfphMCfi/UXFDdO1L9spMd6Ir3IwoYDIC
A8lhvRcQgEvtlIDKuL85ePTGcCx+b8jurwKDpVHEDp/31OCaPz2fNgO5NS+3jjUuqYn76oj6UEFU
AqVdU6rzfntegn3mBpguR/XQsMR9twOjqbT58NpcCE9hT1++G+HKJIMulVluWSJCaPHGw+hfeZFA
HSboeQEKNeCpK9+JM8n16esqTrCkZaZd+R2Ovo0mrOEvI4vMg57pK5ahY5QBxPYdI6zXz+R0LaL6
1oToT83sqiqA1WYEd54KaEOIXK/I3aywKhJCujbyYUDfEWwTsveHULQfSfUyaPXg1/HxK8ayu8po
mcqUM/BO7KKa+ULT6waEier6PJeyKsQInyuXw+/NMGOOI8x5CEOVNN/Hdid/pQvvJaqA+Vk9LeSG
iLPYy2joxj11rhvmKRnX94TSSBe4eX8FokF0vweQe4LKjTm5aV8GAvLZ1s6PEKICfbY6liHopPHi
XROvjmFRcffzpbbSQEmk0KLLudV2FWQ0HxRMzh649XviB4hBHSvX5Vx9RGJajIQQbbrZYo47G9aP
AWKHqu10lTr5Y10Ey7efgS7kkY2TVsIQOzrcDg83rzXTptm1hVlk4axROeiVMC/NLepOLujADpgj
fZn82uLzVLTiFwXIQPJh+9AjjSgIZREXdVodCO8HvQHlB8K86Mu9wMSuQhiI5DRJ8uNZECxW/GyL
vctV5k3UQEPPkIpbMl54iGqrmu4tRUi+vGo8fg15liPWDDkU/Bq+q+MASNpVSUPdlk7eQ1VdnFeI
SEYSLC72xNFyI4SQJ4xLNiWIZSReGFP/jvHRqUgDXCWwCfqbblyIvpFd/4kph6CEw/M14vGdn4QZ
KVpWNfDKwyRp7WUpq32kJ9W89xkmOieJ9qbOBn6bMghyHkHHyiGFTQXFnriyGMH0qkjHJ6Uu9xmt
/yUcN9AD1WmImv2rfw7c2U6Bf6FKH8NyAxRAGxD8fQuIeiMg3caCEysYKFRxufTSf8eiw9y7f1JP
J9+mESI+hq9+T3mJxyhwyt5H08f4fGuqapkUIW/NkvHFlLGsJEGiM/erzB65FhuVMDqB5+b066Yd
tAvmGD/3eCgvxIhfq8jWT80ro5mABqU3ZGOYN6JaS8NxDSFkRojI5uintpBVSgKhnnR2E9NuKZHO
fVfynxuyLC6xcM9aV6ABokCdB3GEGVNhOtc8VMbLd4e911Oq2KMnG3/+f5LtikUV76ugZud6T8jp
SQBv7YcE5/DYxWz+eEhBBaWx6XSEHiex2j4JNM0gy82dgtra5cyrFAU4amRh5yFxjQt34bqggcgt
Ws/TlAo91rexmWV9ADg6M0EVrJF+3UWuNxmI2Dp/JgAyTw9EPJhp4bzooPIuIzJ0CYTN0X0LgD1U
cWxr4G0QTfsVjDGt0ue/6GkTB+Arc13j1Xp1tM7rAf/WikOIT12v7FVvWrGeV9T3jITHrfQQzrR+
hvRTJbwqMtjKzhNRjRh7MHVWXWju+4wcA7tmYMlhKKIvYA6fwCCkRkVLNDvUVxkBFgVgff/vGHxj
sq8DYlWxJ8u6zUDaYGRRNSL2JZ9ecqD7Z0upzO+iGMFDVfa57zsGv23SkR90Vf8Sk7zNXazppu1V
/s93h/ushy9VhRQz1U4tgYE2X9qnAHgXtZWng9EZnpKSs0zj1dRg7mf0Z93fAiLQlYdbM7geGAm0
FAswGIaPCKwjq5YnP3CyN5rNTbopRRN1NjKH+4nSbgOoLhf4ZtmDQ/mj2usIIOyyiLd15yc+jsRd
3TCecLW3YrN80V52mo6+Nzd7G2RcSpBxGUnjiBxCL+qNnrTxDVpNQl/ZPBXLBM+naHC1e4cDaoIo
6oOirz1wE0gz6hPeAnGdqNmpSspBoxtjk+Ik4/rh+H8qjwzMdgd4nXwjkQLb+aRwibV2zGI8Faya
Yyd5k3g7DloyNwpmmX2JJWM6qWfwboXh30ipbsMivZmtg8arB4yWesUxIItazPzYG558hevr/p1P
3UHGslNHyKtvn+WDE27ls6eZh0maEQbcW2+bNUNw9LaIux/LBamRMv9y5fGUE6qYtyklrxREpYxA
kryG4Y2tpsik+jExlqa5yT2qWBYVJjEsmdTmnIuKV0YRwR1ELExhqMhFny0qgHMpONX0QkqY7AJz
3B6O36S16xNsBYUKkIEStcToQyUtRyobfcrsNbQeg4JkrEP56/HtIRwlxQ7Xn72pJgKNBFsm9E6U
ZZRHDrkKMTy7nzt4jcWs5pm10HEnhtnj5fpJ3rw1r/16aNnUkD514fX4Ssra7LKuY+ejkZGQpG6U
NHIsF47ArfHigsuQzuxcnLMJzGffJVNGRGlnyK3fimP59abpe2oseDntvHQUT8U2ZweXzfB01cgn
wp96SrhlZ6GXGcjEz7/dN0pJ2YHbuShWQSTy7by+dn70Wh6n/1besl/CNAtUHnucgEs2jysYyAlJ
RT/OkzneRyL3n13UcJ8GJwCSstqrHC46P50q1p2I4Zsf22/wJ7LI4wohqt5mcQhgHcJE28KNdiD/
I74MAjeMm9tWRkGY0jV3nC7XPdq0+xK7a69qLdCTd4vipyVOYL/Nh9DveSOF3EI2odRT619z+lxc
rxHF3hwpghOy/Wq6Or7iRIiUiJHccQjujrzp443OEDQN/7gHjM8vydJfpliMB3HGW4JILcDlHUPt
wBvD/8+SyoieHiQyuDSfYRVrYruXfDaCJN0HkoL0qzoxOCMbViQmT2ePK0N+l/1XJOpEjtrqLxXC
99QBMfd6WnY9bCsRe9HJZjti9N0ShUvLyeFiG8L+MNkjb5DUF+ESAoQTDBbRSwAjqTDb3gMxgOqy
HCUlNorM/iCVDlE9iH/mXU91jQPeKCjafVBSxr2MS1H5wIeWSTbyHTyE3vR75eur9GMZ/exH9eYK
b3qiSAWiLLjQjSu/mJ+SYdkAGNf0s5Mdb47BvcrJqJBbBc5kXJLqLbDDVX3l35JQoj5nNapFv6VD
SKVt7XnAPj0SQg8rm3IC5c8ewCIdVFN3a+R6vhr1nS7NREZ7zywGoCAftqKzRkNWV9j8vK7UOOWZ
0a0m/UwW9C8vz6BIdqgQWeT0hmPWKwNySlgHYWbJbAAKf4OwZH+hhRQ5qvCrJaSeM14uA76vgAGs
bprP3pRK1Wx1OM9P7lpOXdxfF7DZnLm+H8T9beajYCbfVpgc4w2yz8814aqdeBkpbpsqFYiqMvPE
oMpiMTlcQxuwqrJ4YuuCvAk1//F9ZQb7sBHkisYNIKSeC4o3p+oUnXosNthPGMFZZoe1UgbpJl7I
L8VuDT/oDW3HOIsgD/f51QYp4XSC5X7lShUQrks7ZnNpLK37RNh1F/MBPlBZn6e+8TNiCY/6Zb10
7jtAfTtlWOt53fPvl9mhXL17xSXJIpzZ5PH5fJBajM6p5JdLHiTrwXr1zHnQWITIdcVYoRn+8wUL
UZWEFO+xQWYOuQXiNf5Vqo/I5NQE23hcqG8ix22h84BbGrzuEGE0rW4zH3eXYNTwkqNjKwJpqO3n
5lsrQjwrkeJR1L5whZZFP+u9IhR2hsKX/ss5uzdTiEXvWJHZddoRjYOh6BNDs2DqOpmuX0temKcz
MdiKFfi+1Y0BI5OAO/ANg3Yyytd6d4l1+/0RzFc0FliIHnByIgoXKi1hsxJFHN+acLe/xC/apTBV
G+V2Sr1yzgMeZyc8NlbB5hyiLZU7mVamWmIJhMSsDxqbnpGqOJB1yJc1BPnh4U1lbzGKts+sS/BM
4jrk2nRY2f2k9nWZWQYJTjtPYwX2PE7F3UM83d8ld7XlQMfr+EmtOLzqlW7UpUuBcWJBU5ZNfkIv
BCkbF3PdE4iqNr9zWela8+asUbzsCYpk6sI94Ufx1GmSLy9iQ0xd6h3GJ/laGcNHb+X0AcMu7Xr6
PxEBk1MYa2mcQKsOOM50kh1HlwWFAqJF6vq1IN2dMlyJtPd+eyyFnnEPdiO7vW9YLqoq66oowIF/
KfRXD7qrnFOg7Xf2GYpkm75HxXTsVnO2w/7bDrO5Zya9gWuIrn6hWtzE7ftrCkk4ONXaPbzhvYdt
qt1cAkizFhc2jx3FdyQYdWiQrmsVgo7nPbQCS7TpubH2tI+Lzgc32AwbLpiJ8Y/vL+FYbFEcoiX5
sLbrsFXgc2X0eleiwB2Uayo7kaaN3OL++o7Ly6s2XVx65gDGJnJz27h3vhJS2MgyAYkdxl4u7tO8
tgkEd39TMPz50ZX1VSuFDdJvPvRpMnH2PR9GALS7AGEIm2D1LfpnICw3YPAaGfaUYuTIm8zLskH/
x2hYRLUCApcbyyck9aEZ844AASNEeOqhGIRJk1UtU2gE6P1L1wzERXiIYjiH+Ufjdl7yvIas3xlo
5J6lQc1C5+WZsR2zHSpuKT/qYNeNU1zw6cj6g24cAghU0TnQZYrviJJPVm1aA7xWfBOl/A0lqosD
YV10fT4W04Z+Q4xe4TYzLoM4DHsCqRPbeB6PbyvSHr08ftnXMmlOt9w9wrfc40w5m4O+xHQ7fk1L
r8nuAjnrPuyEnRJuGFUehXFuZrOAvowyzZS3GX9QKc9hnI830DWU9aeh2LtF+a0RM+sGS4golqLE
gErM2Ac1WLgIzgspmmKxGT8mks7La+Lz5MACVatKYOcTUlxGa7FrbvuF5KA/eHH/hUA2Y4f5Ovk7
S+GNAFXtoKVYLmdU7hgruF+ktTUD9kaaF5KsZdKjzYZr6FZqbLZA8tihO3bymkucG1hmk2daL7Va
f0GGSJ9WKOWjnRDC9I31Hw5k/c5DqMaXB//NrOTimYhnTaJ78ewUbf1A8leIDwEPTycjnzMts5Zg
V9Y/g8Zn1SNquXdVd7G3sqRMpZHC+WjgOzjV77t0WlMuk4AUzENCf2u5AoYG+1GFu+0AjKSaYmax
qdjT9TmQvi3Kh2bldxhjdKe736eaz9Py5uvrrB2AxSwmIpsdUZTB4R1aR9SZM9GWPSMw/SpC5i+V
pAzLggUus6Ok15+7bY0+PHLoE5/eAiJMYA4Cg+oSStX7Y0wzyr4aftdlCf/y9a7MwNgrMEj+mxiU
fPv1k2Rp1Tx8Nl95epIQLxodFD/uIr94xD/fm8Y2nCECC6TkrCYBmf+3SipbP60xUielDtKbNW1N
nWt+EaPggQYeB/NLCcopT4IuSfxUvBmAJQn6vTcIpcGl6bnyKNdGorqrrqrZEXFTxmaa17ijlbnR
ri+pCaog8Skk4YdwEfFMnikzZ0FAnM0VNqaxSwy4ReZDXRNKGJGeFji4rvyVY34CW8LAuwWbw3I3
nx9hjr0MdtDyUkj5bPrnJxmJd5A1JHB56PEGYqbx/CgLg8mI3ErZ3qVa3Fm++9qni+2IHJgK2twe
NqpU/OQiwwv+zEpCvjNG5sqkgMrCeQkAAFwZKL+W1t06QHfscwYcDWymxScr93o3LmNv0Mr4x47i
IL/Du2fiW/FJ2sRba9TErEXjOD/u4B9vh6Xhw/yOCQ2h2UIhOptqdWHF2XrQYOXBZB1KCbm8qHA7
tkqwq80XC/QxKNVqZSVKqfrB57Puqz+606M6JcoxpgxA1NnJuW4rsnz9/MP17nKD/bLi5z4uYJW5
hCsOmvqFe9yxDovXChS1QMw9Ea5vzlMVOeASLci+27OBm4DAGGOdUtewS43vFcQM0Cfsg7bU3g9H
CPw0xGmFa6O1m4BT1SKvoFI8Es0FrlilApSDNvI5FIIT5KISYBlS9SCgB7B0PLLi5slBXyvCMV/K
KeD3xqI4OPlpzCRsnq56Uwx+QvZ/cGIiHtL2+VZUAf5V01hSXYPz1RqXjdhgeOynNTQ/ZZdYsTN+
JPKCMkh32F2xvg6TJvytONJ/mOnkuIX35Jc1jgE3TfhMltj7noEY3nMiP6P7taMppRP+bMRFKObk
FWb1je7CV7elsH4trkx9WQpL89H2foCGIY7CPBEytbC6rQJm+/5A76wnQKQ8epgCpdhdyRd6dxnQ
l7fHgRhos+vMFFtxRs8yStAv5D4L6Gqd2hRJeNKv3+tkr0onySebvQG1u2Zh6/5c3bAzflGuVK3P
f9bHrhMOXhtgDFt0Q0iJDBw1I3hbLlIRI9NQNcOjXX47YbV9ruuZbSYNOL+o8OxAhtuZUQVjMUP6
kwPtvrr7jMOwAv0SjfoCQ1hbom8hZ2gYcAELU92zEF+mOn2P350p4nu0qkL+IJixi6yeYg68cVEY
RtC6foIYz1lA84yuIAH5yfirzW1S4+bdr0wNXdsm7RQUb3f2HUcaoeW5AuGWTa9efuGh0geBcywp
Ja4J775gokUm86oJnMLcLjnB2n0IRlkvxqy8PqLv0EqvNpqctrUTa1LLUYvqFLR3C+xu3njwept1
eSe6KxyadULM0VSnYqIhCdkdvxMe2ukXRgIqS0QUzBEG5+Z9yQpWu9NTmoJLley4J9x28TVc0nl7
A1CAN77OOlMSPp9aeWPyaUuvTchuElBZl7/XEiuTdNT94w9QNPLw2qkN/dgZNtsRD/jcj+HFb9vz
EhJBM7/ENU29kqqJLVzrTEM5XQcCwpYVbNtdPbKWsCIUumIHTrIJtWgBIH4fhWDi4nDTFFuTmF7A
FSRVhpvzOBX4DzfYEDZ32N23TOHgdPD2pJToxL/MjhcMM3Q3XhVAw50Oni/YODO21ZpA+F8ZZqbs
uwDveczH3Bon2ixlk7nUUjIuiHKJoR/tVjwwBMwCn19MnI1NUcMcAfVF6IMDRcJaNPcfWhkUY7gp
TFV9ybCcpGTg4GNfvIp4VgMZD5FbBB3bCj0AytciaXxLnPsip0nLa+16DtEw5KSh7F0YAEaO0Z3z
B0yl+wr0JWREIcrLonLQmH2wiDTJdjnpgch+POdPOnBBB1jZhbqdiGFggd0aDsKoHzcEna08lL0C
wI0H49gSs2UfYMnnc/qPP/Ty+YCLCrNGJoh91bDQpZFpoO2ioU54i72UIj7Cc67t7oDJlSuJIEqb
OjdxuHZaSu1oaoZjGLcnWqAlFW/wmjJMX20iLgIIzIV6aMkUBAWrUQL1JJn6HSthI7afBN0JsYr2
uyKnw8lizSWsFRIx5NAcCVuwcDmudsUr7Z0MvWZYxf95pRUAFiEVQ1FO9OlPbHNOtCceUoGikMNM
FtZCc5As5UNGUC8lDl8sq4qDri0mfGe+AjETTpb/NldsxMi6Pu91zNNNJzMXIpaBaDgkJr/ZsWYI
dyEwVd56/VHqti/hnQSefub3x0CJYtC1rDUe2apJ8bNUQwPkVtKGFeQZLhRUI1wFzBbfnKD019f/
MbPqM3W7H/UiSpYcnRdzm9pRrgQ9fYJ1tLdD/bvYl8nuISakDDH9kUQd4c5Hfmcp3jIkoU+STVgW
+lRv1f1BhaR+I/Oagy9e4JipmGCrwrb37fzlGorOXXt+64P07Yl+TrxCHeVRCHBv31Y4ESjmSsu9
d8IM+gzvPw38t81MgEZYDqlTNmTW+GbH9EiuI3DYEd5TFz9kAT7VIdF2b8HAJIjYqAWLnV7tii7h
dt52PWv6hFjm4fKNSGy1XyzPnZD70UtuZ/aCv+klxqs9wd8elRVj/EBR6PwjeuPeHE05F/uVSz2B
UHNywREarGNm5MQJQTey1bNb7N93ChtOEiKbHcNN65l7nkJsw/Pkb5XttMiCfQA/K/HmHOITbArr
2UddDM8a/r4BhMPm71SRlkb8iTZKtCaOaWnGGxvQB3K+fmQdAcz4zvsxziYoLprxf2XfwgfT+AiE
PRKpo50q91BjVEIyZYSkb03Lmvknmpn98xKgE2AQU8vwR40OWz2SFpdFG2c7LTjd0cF7TRRjChsq
u5X/IJlp9IaOTwsgnbMWkxN/ddY6iW8Uiin2mhShrBj4HpDGflnxd4eWrCUVUVc6YN1DWgYyvOQP
RW2vXx7IFc16pnzxgPN/TLLx+G7k+5L5h3p+YIcXAvM3g0udLXm5yd0fSWBhYH4OTP7mGJwTJXZT
q+QrHbUkHiEQF/XWUAvPFmzjcxOGjZHqUHLsPKfn1nAHhtn4jmUpg2gdjqWaNCvowD4tajGiR+3o
x3uVbszCgm6FQKe56rHTW6ieTyIhPwr/L7pn4ws9gFnAh6FY0GpYMep3BiCtW8FfCIemHTnTKTGJ
K/n0YQnsen4afvpPguJsxht28YpPo0RLIVFtBKxHmklGbULLnaxgyJwnTTJVhH9KtHj0k4i4nXNx
81Jk08EaEdd2jfkriiPsLUNM4ktfJoi7aBWUvSCVlyK2C0MQ1+5cKnLqTKU8Lh2gff9UsdD0Ng50
JdcGm0aQxSNzCuT7E9lEQD3cByH4oizfEky4wenzZf0vi1G5MUYtPm0a12XX1w7qGMyyzaoA8dlY
/DvrwRxVwMSvJbviLX1l+r8s+dCToGFWsr/6XlRcNwivnehiIfG4AWh/r/j97y5yCKnXZONogEEn
ExUGLUyOIEnEfHzb8N60A3bCFIP7EnBljIZ+x0ryQCQHcFO8SsDrvQuBXXrmkLE1EnzDn/UMIyIN
ZOhIPzTF4ZYWOcjK5a4vEZzsBvl/8yUrKaG49rlwGrtJlOtNirTraFRjFfR1kWgDiT3/GdHh5Lg6
Hg6Q38HHgUFeRJ7ziDehfKYWkCCtazE8QNJ4bWDmpoSPOZKjTVSvDk7D0JgoVh4XrEB9UXLJbgCC
ZVUOl1ms75gFJaW7iv7H8Y8y1gIkICpn4udFHOdKOE1cQjCRN2kgwl4XckhqatXQRvqYNCOjchYU
jdftZx5w1mJodoYCrIsvjYnUXGKla47K8FcaLN3kbkN1QhO+f4cRJft/ICafFbWjKj0A1FzHayTc
/jaX9s4gylWOEge/LEcO+h/+z+BEkZUYVopMjRLxdKIirL/KORM1aksLGfn3mpgx7235cphd4Zf8
9mhIJMnYTyZU64SmsmpotR7ci0gCORMmB8/Cpb01Ami/SI8bhprgbak4lBHbEriIiHlryXKWMf05
RdDDVmxVoxXDy5npTJWd80hjE6yMPSPnpEtx0vHRPgzr6UjWkuqueWM/dBaK11ZlNk+xF5+oPqQK
uWlqvzHyA+2BSPH97aKMFi42CacF9ZsePl/NR77THY8Su1Vk1cGmETlOwJA4wwMgOCeWMAzZkCst
kgpPtk9zIdQeMK97EFUIZ8AG+M6dZre+qw+LWrK5mv4fARJ0a92DXg9qBCUdhYo9EBsgZvQ/lyLQ
PCDTGohBq5vh7kycNNxAfkw0CQTcy7FXVpb1MRv/lyJjVKcuuDrW+4RmJTMQ14iK2nPBNg9lxVUJ
GL3NsqV8vW/uj00G5UQe9pcyliDosD6iuiHlOjeDZVNQoCavPuV0MB5pItQbu/bAYKdmAP1+iudc
NNiAQBjVVojVvhpanhwO0TQpU/cj2/5WelQwJnsgNbDbapw4f1Ze9AMGTbrMWPd+gXl1d/rby3DV
nc18M72TzroCx2NMZFP4L045RZRI9RtaSlThJvsu+wxQ7qdv7wROQ3zLsUDHhnd3MJYBwUUDgp9H
b1PfqZ1ol/jYICIRuaHEAkOVPD6BqzaSrDiq52i1zxx6kUQAxVMy2ijkSm++3Y5mMV1UaTbFoBdq
XozFoSG2bAvfAnIBc56KDp/R0e6cee2+Lx3Msod6PsXYW925t8McANGc4IKLpjvqfYHm/RTMitpU
pGE/Pp+NTxIUSWbxRyx9pMgHEFlVH3WCEZH24aj7MrdJN3Klgc6jNhwsbyjXf9H4S612siSXCWCF
JWdMSWuXlet6fL7yJD78Xw52BGHwLkwXzgSgbbRAwFcft38/c671VTRMyDZd8OLT1PjuYs/stnig
XpuetpXF2ddwBUv8gOjZOZux3BcCRUB43p9eTnx8sDJWRanqJZq+3ijzlNNMLtUmjJHdXreixYBF
JK65tdhZB6+EXv5zYW0UFjuGyZiEPcNZohoYNu0fE7Zs5kJNsFh8exq7BmjOo7LlJ+5PJAE6PhJj
SyX14gPcYwYKozu68DCc5+T6DezfLj50h1wXqWAGKUJQKZqrR217st9LLxK+O1gL3jCdf164y02R
hvVCF1H2xAQcMEpTLTAaOLlBqqKhXtALPnpGkW/BY4dRR3jPQn0Huce3ig7PpIN+3wivUGJNauDZ
cbZz2C4Dz3UosMN6z5RvcUlVE83ha6zu+fA0ccbRFxZ6W+WyBaOCVf+XdJK5Q8j1DBA7df5TboHI
3k8XU6POXZRDTlzq1kyDPIu2luFZHNe0j3+X4rd1/gfU/BbtCSRKEK3aMAyVtrlgQWyCrNzy7eRU
s6gMp6Ve/Cns53v3niUJwakEE8v3A531Fwkzm489dCgf8c7xup377YkeOl9BT1nc+P5HiJTZRXxj
VXsJO6ohgpgSTxlMnWvVerA2QtzIvKaOdkCOIcxxrZRPf/F474QfONsJc0FIAyg8gpRJf5Mxc7ZM
DV2/d8IynDHOMJagM2rL3P7LBzH5fM5SALhmPbJvcsuGjJEvZYfLo9u2clzjt/K8cLe7bRntBu7b
K3CyqCBywuvt4SEpyBV/3g6e8SId5E+6vsZGxcUsKOafr9f5+TjaJmwB+4DXF9CCn6x9iRcV5aKo
ZH14Oh3K+7qaWdch3NALmPIKjJe04uvunuwXoUc7KkWRwdaBx2cFPXUgyWR85Ud1P/s+3v2Y7Mgz
BfL31EZO9+04ExtQ7FrUvU3BtnaOprfd99MS+BeUckzDhE5ybQmW6cfT/qp/X6+AAL5Gc/C3ff7t
xjW3FxH+hFqTx93uVi7+bSgfZ5s/SCkfO351t6yD9VPYktOxDf7F9ZpmJv3l9O87I5FeIg6M6i1D
L/+7YZPkx1vuJH6V2I7WRyS/6jZmrO/k0xK62VNuYcHuR/L4aHIt8H9cT2tZNmOiKrkJCyZAYqpK
xfS6/O4EWfNIio+qGu8AB/CjCPgm6bLuAJwipDyE9usSpILxOieCqh7VpBLhQ5FXemp7gbqScWRK
D30ztuU0hP480fIlYlanwSd4dnC65nbmwnJJxpO/CUIpY/tLhw4fhNtFMRY3Utvouhr6qN8OXW3y
R/DXUE7BZslxGjOMbkDW99g94RUG9Q5MZH9PMAaS6kA3+EHQgAk64uHNzlsBjo3ugIVZA/Ny915n
7ivN7z7omWp8mnu6Khi8n53kW20VIYwdd5MasFc1QA1HsHQw8R82mvPzA2aCi5b03lv5ySxEi30Q
/xkcTP/pUuYN3DO/IcgwlzFJBzKIwGVkDZBOYi7mqbZtosFXWOXjNtOl6ak44j8NsLgwA4Q8kQgr
F06rtF1yelIGXNWMk4fb8MFZC/5dI46Itoxgmk7EZ9UnB5vYi1o7BFY4Am4sXClLmdh4Oxum/lVa
Ho0imWc/tPGBxHL+8MR5qy5zw3fdDY4R4bWA96VtqlRaxmZVcbu2CPjaJA4b756T8dm+3QWDX/v/
c2xOmk6ZP4EgmUOz5hL3VwA17FQ679Q0nY1Z90ndmsyPTT4+BJNX0vJFw+7fdU76yeK4oS88zLiO
x0/Q3KApPVCAvjWR/hLLv3kAcQUCVWNEJ9uBAqiNm7cG/Cdgx9qXy2nqbhcm8vZCJq/Ka4RzgUln
fZhOyTQy4CGlKSmyJ2ct+eUQxaYSmfyaTwIOR6fnVwMbdIF5PBg+OwKcrzfyHF3NGMvfjFlfTaaN
JExn4EAXO2o4gg+AlNG9psNuwjEhgazIsZ59xOLTsVUBw7mD/qWqnOsju4FhUvJHk1q60EK5LVGa
HGlqnMj7vxokNuLuNGJQ3NHPckLo1kEOtFXSjiA5Ay8owhLOJOCipceZQTrTUSvAvyhyP3ePzlde
GiBU4X8QEdDfe6ka4kQUO9anwG8EFjV7om4t5O1sX5/fk6vC1es8GB/1MffoBHNfG7V3ih5Luz/b
/W4e+6V/56Zt9R/2ezt7aCtgSjaolZSmGY+RomKM+BIg6KjFgzJzHkdiqhBwxVqihlQWlMKws8SY
bUgv+2duOMl7QY+ShWY4FQRdwu3MJNp1ltOtPyIhG9sqAuUftB5xy/IDmEaX5s/pCcjpNRqWmCSa
1VOzUWpVMwI09zyOY7uzIJTj1UZQSV2+UDr2BowOSjsYdWdsHpFfJoc6UHQ6jLVuhJeBhio5pKAC
dKet0+qBSsEze5ahwjtLAdSKQ87kVYwNcHVCl00Yy6i1pVXeTUOqssWRqAa+/kAQavTxv4ZtGcVZ
JSH2VtSvkH+MHwQd2k7RJdPBMLqXhDppNd1UIqf0LR2AHMpcD7SDsGG+gOpkQN7R09ELZ1UGPRWj
U20b/893GKKY6R6nPLnUOXRcL0iIQ8tEjipa0Go2+MgnyNiUyvaZnU+uFbp/1Zib2CaAOidL2Ukb
hMKpn7gjwbKrwrWs5QUSC2FvQhgpOqQFYdOk/asAVKCuC/zumuczi9enxWibbgmbHkozgPTSzMKn
Usnevuj+wpkfls/DOsFD/5mUdvPhZisGv6+y9Hg3Slrrr/i+pmh4jkVRfRXIsUtVtxk+c3xY0k/k
qMEFtof6IIBQaobIn6+iQNV7sjWOCaIwXx6yyXak/CXGkKRL26iofVfi2WChs1L9M6kIzyLdd8fM
2GHYcInGDyPRu7YoFozol8qmkHOF9uvP0KFFBhl9FsszZTDCBlU3Bq18OyETd7KE3vLhuvdaU6vC
lyassA5QAJqNHOW7Je70iuqAaMZ+F2n1zbMxfQQ7fJ60g8pgDYI7RTNiTDwskv0U9MC6TMg2tlK4
j8qZMXWBxxtDCfEJEdXZncO1m3uKqZ4kfR0p+23DFsT25l++fGalFQXOsA4kqjDRVyCaTa4hX3wh
bDlVKQ8h8VUQlYt6ocB7VBAQQiCxl9s7oSdGB1emMYQIsInxoZNyk4TL4kfFelAH542fHs1objaV
Vn6FQl89LMLKt8Kf6PuxU6Lx1d61lFYtmRv4LtRor+7REbNXNgkeWs7rPoPWOmCzXd1w9X3AAwzH
jrkyLvvX4ayPj1STcU0spr5jLwrDWj/QRUKUM1yiMqMmZ4cXAMFUC+TW0Y4e4YchBPrloIfQkeUh
6chtxKwPqje5j9B3jm+BDdZ/EVy+hJlNaQSV3BVv7XnJB8ZkO+omNS5HzhkYjgIMsEfHZHLjvFdH
CCt8jU0FwhU6oHDGKQrSxwZUO6rIZZnbNDUt5gspgqZyVfhizldfGsQ6Us0ehYGZPogUpXdTBSBj
P0NTCEefFuLUCejDb+AICkESeYdymLswDt+kchOXz4gTTpUXmPDP1MGMj8O+/pIYZQPydBhhYKDv
7oZHVdnGoItyAQ/IXVnN0ThbsbnwP1pnkWXRAkynNTM/sXdu8Y07sbwBql1umuVRqz2HVFp9NIR2
1o2ktrOZoM/u0I+yS0CYEtaNYsz0BxGXM6Onm5ZrkEDug9iwdMMYmKeSSTCFZzAHSB80YbD8/IYe
HFjYhvJCLsul9G0H/JkhIOytif6tTYNLzWQ2qNKlnGQTRi1m+LraOPcsvn/IVcBJhvRGpm0JMp6u
v9nL5Aa/9jDefXo/E2dpVPhvG/QGDLGNy/gOJRV+gUJBmudr/l0gDgw9Q56kdhmgcNxpGmS7yLf0
xi76muPofC4apFlOGi8IpK/fZHWTRW8Y47ueOFmBt8dMVoUywhjHI/dV27hCodrPuu8xXtrz7v+r
xKeB/ZB7RAGOjfdv5CtyjJvZqRENsBZfshVqFAip1xKp4UG5WkPNIRs7eGVhDwp+57K+w8PGiX8f
T68oP7k2k46nv+BfHgBCsSawZlQuQ01mUSTS8TrN01tS0Ld/Kv9W5KC/ORjv+RfeIgSm8BSjnzUG
Z78Pm+w3uLEhjNhBefJT/XzYKgxQopJeRBXV1VNUnWOWzijZAweLuA5XDXQOaagIx4Wj7bBLHccw
BrQyazBVtu3s3dlICA0G7a0c/vcOv1Yrs0/omEODUrc4AlNTfRdL2qoGiOcEKalGKWQwXJ822U5U
j0uTm7dQZF49UPSVI4znOYRuxz8cIo9yfGM/IfycdD3p+eCq4QR6HaWQu6/yV4Nlst94IEZbk8H+
nlkaO7eplJWujdQR0W2rJylMLtEhEC32picMyZ+stQC5n3Sc8qenoNS7ez0mbkUBeCIW+bnfk4FU
RyZqU+vh+QWEvPnwGRsy2VMb80Bnw7IIldtkVyF78D3W1E5pVf0DSDEnmfAvIASoZNqrp4lb2tNA
LmYN+NuplMpqkFI8YSK5+fWYKAdrRe5L0ZOlIi7/dAy3t5qY3MWw9UkLntWBikmuQoWLdnb+Bld9
lz/ptX/ZYS1GjpOcdJz2ZRRPbk0NHhvE8h/35T1EOespoUFWZPBBX5l90YA5kq7FE11F1Za3TnNY
OlzY3HlEuliZTulOM0XfZ8z78DzZDrssXyTMNG7L+OxdWdogjQ81ldpnKrgoupRgAnenVo0tmXNg
wFGdz5UN+YzjTzG3RTGQz/6Z9zmFTK72nI0glpFfkWKdGEE2AyWwVYV1PYFrPyjl1J0oGHgbwm9c
rMq2NoW/phXcW55rz7kx43wZWIzlKmDDg3++WEXYLDZERAojNqB6j0iHiqV1666bN8UvmXFECcuZ
RYlAT4SW8K3cjpJkJkaiYAH5IyZoumgUvXssmVWciqMKuMuw+VayV4kivKd2DlnJcPxSMnAnMXel
+w4NDOsjAqQ34Vi6JjSUGb86IugE+YjBKupy5pqLQXk9CT0OZ70wIFM65DWCeIUxtVR47qL1uN1R
wgHPi+SSn71ZiNqdzIQB1Rm8GWxdVF4BFP5vK0vd5s9amjgbPlM11E3iV16n1sfL69VW6Aq/4Ywq
DorPX/K1BFg4y62yl7Bu+/455UH7w8pqnDDKJ0dxVH6PtwJ345FM7NuP5OCxk/aGGxGPin5s0zz6
W97lOGnfYTlqYhuM5BlgRW+eM9SkOFT8t5AHpigh9bTkIqckhY+9JLDIh1PBpEizyupUEEWYqmh1
JC5qJtnJFpreV47R7rfWXJM8o55HjQPDKktOBVZmfifr2EQjh62anF2SLzBYBehfhNtRE3udHx9L
kluhzXagMGG2Q22ckliBi/wLBruziRGsETXgfo6k6E4/FU16b71HffweIVk2l/IN3XMIMIo3Py9x
ZeMe+T9pb8km0+94a5qQlfTwQHgWx3JyI6mPwQLKeal5Yf8VMZl5UO4kpkA8DKf01txpSOoUIuUm
EaDpG51crgS8Ki6//ctqJqFnZhjzGkoaJ8L5PfTKp7CX6Rk/OM4Gl5qPV/MNM8klSTdaVLvBLb9G
DqdcrAyHYqLHQEcm3r6y/x5ZebrGyyMxrivsnNnERpWnFx2jlJQcSR2/QeP6O4bq7+FsHFhg5x0n
4hRYsYUPTLVLeYNY5Krco2FzGtcw//oyPNUH4prFlN2q3uv33PNPkAVRz2RnBqDFQ+xxTsmuCBsx
sLnxVPj2zql0Ez8HhecTBQY1BqL1Ugd/8wt8CDlZ5ePcz3Ld8tHdU4z3ut9p0iVetUDaMmD2mKpm
1oPLmfZN0kr4Nxbk4RFYX8/08lfvu7bqIG1YNm4pdrc1tBf9elTY/7MZAHxA9h7E5mu//SDZmgja
41o8acPK4M8B8U4FRrhTGd9LlhRSpAxlkA7Lbye4qJnUljer7mrtF7etm+FGLRd46PHuurl5uBg4
qVz6V0MtC46CUmXld8Ph8IQPH+hx6UKOWTgzLiygtBFM0uli0Y4eju5agmHL1qcBb8YOo+ZRTJE9
xDigVgFl8Lztql/geWT+EUn+F7n8d30an74Kry8+O33m0JDANdj36GhrkuI/BzgROxjpyIDobsJi
SmjoaDaCGh12TVKj6EmhF+6Zs5wh/RxPJKJ2hxAZgE1A3eM7NVK1GYf/4AKdfN6aoo2JX8gKS8vC
idQ9r3Gs3ir1PFdur9fTDy5KR+hTO8t+p8cBpcWRAt/cGOQ4GGeRYuak6C3jNYr33/eZFYlz9Ga9
pbx6U4/vJv+4weXME6fmY4ywJnzrtFQ2zr7M9y5mRyEuSs7cnwdSZorLeDU3+MyOB5OyAQ7Yeilv
ttm+w47lZAwu/WlckWvtgmq6HCmkbLbP+YZQBoZNwd2548SZPgyoHRXE/J887WZzGkSSQj+gvsYP
iNxPORvrbG3/AIpdISykXbjXjURWaSuamjo4519Ng2ThoKlT214PfVEPw7E6QfXoorNcpxejzGCK
iR7ho2xy85QX8oVnSifPyicuo5M9mu30Bi6R6GxPmbOc8buc+Mb+Y1lRkyvBNs/Y6qrr2hqiQ3nr
pFeucZiCeB95pGsHTfqszZDSdHPXmFSn2Svv6bZAF58PvCAsQLCVv0DM7SDNL28CIeYrHty9Rx/U
DMFmFpEFdKNSw+npWI8OR/3bHaGTTvq0FQXLVxEmKZsQ+ve8iu6T6TVnbRTGBLxD1tsAyO2fJb+u
V7QY+Kp+LsDIEs+qVcOwLhKgcAiO3PBZV8BEscXdABSPbd/AABjaTIhfDi0Zz0Mbv4SLvAnEK5ix
Yytih755DIymRt39pFwLNQoFcBiPwbOcTZ+Clrk/90qI6zvGStBzXMKAB4PMYOdcOC8MTGN83+vY
NXg1e4NKipGps/7TcSPTY4cX0GRHcGb+MymTUtmrtkWUwMVS/d3PkitOYa8XCIDe+slYWEhzIsDG
DNz+X6y/mBMN8OmBQ724wOodTvfRhm+EEBjXa9WEMR7JxsUv2Weq2g3YzYphDbT2sm9NsE2D87cv
uS98V/KE1PcxcbsSPzrNtBkJVHeq57VA52i76xuvcjV9mAl4jnJusLhKXFmti7MJoNV4lAkz8FkG
+g2tbeqMeOQxiDRl8S3s4ANUCrDNmoi/s6EzT9QHVL1u4xVWk3olaRPoB3BEdn63bVy+VGjLQ7QF
2LuyEg+eDgH92vE8CdZyvgmN/rWmWY/jn7Os0dh0kmSlx2KcT7MZWWhJiVA9mjvzgrVeE9RKzuoq
52b9m/5L8r8WnJ/NEQg9ihuFLODiFQ+xS38jAoK0rypvFOsJrG78Y3kfsC3Rps9NA/WXtkpbayMU
DoLH7KFiU0/wckb8HP0uyBSNp4K75xf0f2GhvTj8ijAZfy1v0X9vpMHnYP2R86lpgFJQUWRpdZzF
OvWoZTVp2lcaUrOUnuDUHKWcg1jM9hD6vpCv8csm+Td/aPUrmzpmY/l1ItmHN6Z+wRiLNz+lA9Wo
PmxTYshocXbEFLtl3vtzQiKGoqa+8P/oT79G1WbxsawZv8Dhg5aV5xRK9esLMMrkSLucZpI2C1wt
MtRwmldApoRBbjCiZTXHyjq+gStm+FWzYjede88ewNhRnyUUxHpXg6mBzpXyrt/Xa/u3Z3riVS+Q
MVv+LAcsIG+Yyt0GXcb/9IK8x6yPvPdVvzRdKXhKqgklTe/MdnOj6IogSjwsmkGMkT8hjsWGKLQh
gXtbTdzHM8dzS3dt7BCXdLTDbvhyPArB8gm4bxYVVrlFNR67fFZutxfy4t8jHWDES1yk4jNYtscy
lG+kH3EJZB1pgZ4I6VVGr3AtInxdyhZTLLC6CufZTzVtnG1TLene1I5YRVVcICqZcBw12FVCpiEY
1IgQ1H0CPZVzlvVWuGG1gQKB8GlQoqURI2irsWCKg1rZQ4Q86+0zhzf1tJeFlM9GzwOwztVTte2J
C3u1lYz13OszrO6bPGcQsydYUjtVESM/iQokhxNyLGGNn8QuvkA0uDL9z52JLc6+V+McTfkyU568
UnqPmVxFDSd+chlX5MABqhioB9vcRjeCuzVqPJQEqx1sLfGenN9aB042LtQbvQA8bfs37syxO+Cb
nrf83ADXPQIG2XWrkmL9nuIRhmlPc61btX1B7PorakhpO+KIo18YXiryt9BlSeBgYPGO2jeB4saH
hed/+SCpNob2IZH3S9uEpkQnf+JXOn/J7Baok1Vw19mcolWyRTHnqHWNyPFpQIyJq1dDYK+DuhH+
5mB/xMnuibWzXZTwvLRupw8I2hBwA/bcUmBljbkj5DMyrf2dEXTfEQHTVUd6VsXgit01hBvM+/XW
47Yi+nDmPiV0CDZx3DLzSiHdm63Xa4uEEHlq6whvwAGqY61kpQSWIbCBAp705iN4j7uFmUq8v0bk
1y096GcadlrXo7PH7MNUv82IGwX6fvLEllWUfHNiOpjHyG6mCFuTMXQ40KlvCuPrQK05uFyekqYV
vnVwgMHqh+lB8TkoEBw92+iKwjUrWRsbNQTxhn98/MrnyooY/kt3eprPRd631Bt6Q2E6eRwXiHYk
9OwMMwPL2bIjdyGmNTlEg3ZkCBwbvVW7IHOuIJUZldYqTGqbKnXAUylrDD2z6Bg04jseGcj/6KJ4
/XPJ8QzvTXBJCpqBiziNRIuBg2UhZnoBG/VUh4oJvnH6a8McqAjBv8WuoXYVUi2TrBjBZw7A0L2R
ILIXah/dPAtR0FuD/aQcjNkiIHzWvCBIhjlZ6lb3sUBR87GQAjDNklXG2m59VfPEdkdkhSFek0dR
u3npzpcuQmO+2U2tRQ/eu88rsjmJST999VjwCLCSRq8RDFR+87n0JXeWQcuE1O+/4bl520NcoFvd
d3M8aRm2MPjnKoYYuCljnEtGLI2SU3tPJPxdvouqVoRNOaVE5YoKiytCPREPvpHk6VWN8MEG9NwY
/BU8sfbCrQBcvPI8hsbtz812geSVlJo0ZBP+ChOw+PYpEPEaVHStDWeIqWu6x4XbcTdjNbv+8MHo
ZrjY9cYJaEaHx8ykF3AX3OU3UtPQlqT6x/PbKaLs8d0v7FWSzsLlw9mIpT/lmHQHDHQbiZKSPDjN
zVj61Wvhg3R4KK3BZ0hM5J7zwNYva5HvcAa1yBI5grLYppRS7WeyCHMLqw1dnIBYOSzJ9V5XW7Hg
izUtH4wywVSS8zwTpspxJ3slVbF2ciBldGUoTHvfgbcXscwFc7aCNfq9BwlegLckosbZkXN5tJJM
6ITp0M5rD0nIr2qW4Bgem9dfCslYEycJkVRZDN6eG4a/wX3x8vqLbak4quzVVUOQhJUOp+ilMgL7
P3JbTo3b9/edaomEJZFRYybMztOaIkNWF8jurh0zFnpQhsbDPY4LF4uz7MUd3HWz7R0umGL3yOw+
1V/B16fp/qu5AHbw8GyTz1H30wOmkBON7bVB/VpjwpgLDtZ/HCdoIZ3chR/LJX76nbz/r2CVlw1X
gz/c7rfGtMI54sIiRv2E79meNVRc6kV82QOKSdPmE58sUtTLsLnnN7by5sB2zkLdn5DbxqWN77Q5
XtsiIJdkjZ+YIXKvpYEAFPJVL5vUcsy3IBBH1GSxaaSvz7Ypf16YX7tVfb8pOLYx3ujoQs64ScVC
QJ9x2YZqPyA7ltkWaw0gNjJk7lx4o3zi2+1FySx7xuS2MceVCwmUe3UU0YbUAy9Ln1eD5BTKfq+D
evT8c3Dpsx0b/4r2rzJH1OsVRNe9MmMXMkOj/PzJH7+UAMtNK7NePcakHklPS6/UXtgktMlWsPD0
j/KqvscIStOGJxd7F1WD9WnwWvBbnCF6kfh+p8jtlS4reIZk5/EJUDzGPBtnqdZFb+dlS83nVJLQ
Do4gYZU9zxhSzLsks/MGxL/jo8ydL7FjLFOqeUMrYuFt8xkETX2HKULDn65yLStCRm8maJSCFw7n
ZaJRCVlLpbrQ8c6Gbd5zf3CclshzfVVqBbqPWHmfT51JGnIsqALY8T2ladWs3+si9nNlK/cq/ii7
UBbor8YdciN9DkVzbZ1M6cP9YxxE3rv9ruk5x4Zg6bymxPYU/BRiDXqCZmd6VLkFVaqu3b1PaNUF
CqA889dpL00kEHPEUyR6IssolIXBl5JwYlIXIW/PmFOnowIcP3zbYR6D91GVvcxEg/sHKcEXS/yK
5QE8vUVPRNxfMs3cAs3A/jOMrlA08ECVw8lp7I3h2xtrsC5IbJ9YXVqNanIRdCznTWbIHLMZGRvv
8VjIYKftjzmBd9Z4g63GI8/Wfnxj4QNHlYj1bsCTHV05suZeBu7rtsLW+0pTtY2pq7ukfTPqxkTY
hb8ZdG7ulEz6qvO0xOSOGlvkALsVRncVci+2qNtnVZCAcTEJx1kVQPsybS48WdkBM7nKCvImmAYz
cW1PjjgzX9TsYzx+DQ8EqxJ5ACfbuR3x97AgWd/o2eZ7HrMcWQsA6/L2S2YckN1k1lfc0+UzWJxj
XFzI9NpNfvPcaQgPOKJIkDQ79YYhAECKDeFuYD9V03ACgxKtOrHhvGfGE9ime7kOlK0RILMTGhbV
3+RnU2WjpeqFmck+LaIwRdnD67+Mlgemn2+at0ZvdctV3CQAU8CLxuNFJvPYz75TFt8w5eCxRAdN
sHKB2DzknEkps+UNTanFt+53hM0+10y4cN0+qGxiMYZ+wIUAsWOhRM2nidOsmamZekGEX32WCpqY
23mUxGmrbf+bsZXvTuevYzPir3tSkQoCFlL0GolkpwworTRCeNnIBR9y4PPQK+Sm7atSsl1PjwoC
Z/664KRs8RyL273fusBSKhGDw2yohfm/1GW3zWudnwngoFchTOJ/64R0t3yLYQ0QoilZ+PmwLYGE
KJsCjpVP7qrUwGDVf2i76qMV4ZMndEuQrOpRgGmYC5E8FCTlvivmBkvOqKsUagsE9Jan+gUI0sFP
I/oAUbf/nk9tV1PGwVwjyqO9l4jMtpsti92gaglcY/nNqjWPjUCjS+e8ytwRy+kFABClyBSypS8v
TkQbTG8kbPg2sQViRKscGZW35zwdoqnoQmvuwOxMHlgS4lkMYOYAJ+jdSVOd9y8NV9vOtJFlig3B
r3+piWk+6Bb17/4DuSPsAzK2wsZonl5CLPR1MHbJXR5SsyoOyXrgGnyIooM9NBOVYTqKY7v+zRZv
eAOf2QeW6sjFEJSR7rIp4eHLVLQ0wcKsSwDTUGAyuRPbrxVhA7wm1kESAJQj9ECcPRAK+tAWeVHN
DrBEcZzYr6AG7OulH0ANDr1liqpzJnZJShKc/I/gguHjm4ui5KxZsYXvtS2MV1VgdmJx39O8qFdU
tPL/E/ErTikbmIcXAyHWn1Uggb337HNc9L5zr8L2mwwojDogbKfknTi1ZyF0w0h0U1MuCQNZmwSa
SD9Mb5EdtXXXc399c2iiLqws8bcQ4tNCyBTAtvHOSOXtmTJiiwGt9+ot3DZ2nGgyWsiXIH1PrJm8
uLXMoVCsH6zePDB+PQgihmAdIvwHrH8V6gNvvOhCnPs5nF8HOvxKpA+5QlejGu+B6rlyyStYeqaw
G3fxVkYp6cNJi9/wSziHiPqRTreS+ywY4a8ayu2xLPITmTmTcTvLC1n5BiEu/nYnnLS6U6e7CWrX
Q7h0HOsIEbOMNLd4G7ekm0EqOUBNlc1yGYrydJPdByN4ik4AVJciKTTIRTTvZCbAFQ8Oz/LZdbo9
ifUjPU5MAbmNW1WJiz7ofu/zpWX0RHIUP7aQ+zcWY9gWn56VU9Uq3YCYLF8XOglPuYbNuSgyAK4R
Au2fNDXRkwasV6HMxa4byrTWqcDnSfcBRpU2eQIyb5YDDEE5j1DBzn/58pGbQ141AaXlxWmJcvMq
wrVx7vZY5tXAyWo3D8iiQ+FhuJ3JYPpRCMrlifiTCeg+mUmrvvTI1fJDgPtRWKR1wiSrSv5Omho3
gnheLpI4HSnauO7XqIGNe4a0DODN0QRSAQS1Oeq1EEZre74bKVHOCohNWc/9x+0bLqPW8B7VgWS6
ax9ac9ehaT78EBTtPuhVo+9H7M+RKrNsWdLIH9S79WcVR9JjaOyAcaCxrNK7uzpjYvrFdqT5Iq9x
DyJM9lqfrqR5zPv/hN0s4Jl7EL4zkpjE7xkjnO1p94YHYkeGMn2ixiLLc69Mp16mWk/C42f8oAwP
IarzYV4OCic7rstq6RrGGsvuIvLuTcWq/UVriLKiOAXwOGY/Gkv8knCM/PehWbDFlAB5RALPn7Ge
mG8pUZFMFj8I10lTjIezuv0tJeT3tNCN+XO3aIh3IdbUDOqA2KS5SA3JXFmDWnMpC3x+piZsgi0X
DjlOVt8hzIMJQLsVuLcRfVHIc917LFhElSDpOl/8cXemrwqJnCPaXxOWXPL6XUwtzc74fZkE7J3w
UMNVDm359hdqw8qHaTqvI5xgRV8qcrersLgA93hmjvsVNCmRATzkTWOaqzI+45kL8Dyi6Y7dJtt2
t0UHuGG197Gn7cJ1o8fkgKOx2h7yOhzwstdAW9ldGkigqZAOoXyyl4CRIGCWK1EyDzH7Wqg8FPUP
zDsoTdwS/3LffyBtrvmz7TBX43WDVRTQI/mP8NABXLuQ5TZu1yJLg1FoSpTGY8mHywFeG8Nro6eh
hHhmeiHUjdfihn35o06mfeZ6KeK3/D0oCNs7m38a+n2+watwxWksTeGrJcO8JbePYGgaAd7CRZJg
iQTqS30UyMH1c9dGoKMnptXtqxQ4B/Bag/Vif1RQQozfWv9AERWDNEo7bIIB+CpyaE1/2JD+1Wjy
UyIzcyqM1v27UqVihvV1AKJRbwBGmWmVFIVXYIpvfAeDSCKOgPhTlwKSW8toh+MRK6e/qoziams7
uQM/88xLaR8tnZF61OXw85IqK9FncIjK5nU6xXvXpz+ir536qwpTMUVfG7X80u5fNTuta/9ipWyC
fYJzoO6JTzRAsmtesFRKJCmyO/jPKmIu+tDi/u2mttL0eiR7p5XDH+K8KAUi/qpk1YXfJGs04RKk
D2IllDXglkOUJM8mMMLQsNXh3MUL7q1yUJQiTsJc6z8F+n9tbVflURQ4fP59nqk+0NKD8wjoOUsX
qyKmX2siZdoGPOlc/HIQ+Bl/bqJsYn0AfcXj3x5b+MlA+1d2Cw6ERnQ1ke/splY1aGEqi84MG/FY
ljdZmTC4ifdYbhXopLYndJdAh3Tvikrgpongty5hkZ/vifwYrT+AVmyjlmlaGQ1n5IIKv4AaV7dw
1+X7AKOgSeNa0Q89NaRw8cIys8aJdG03azmxmIOWRHxXAOECgS/IU0mQRdu/EAPy/nHJybvgkgHU
c1RAmcCq+9+oYRGFwkXXnHid5fkpn3FLCUmbmI2kH6Nx0BohJgaynwX7CEaH+PLSXFQtxws1qiJw
s+0YcNad0eN1hCRMRtG5q68L2OEc+zYH+YYVYc3f3uwg16eXteVJFVNz2wfBN/guHK9+nRnwgTUB
VTccs8GchtvsFzGeS0yfZGnPFu52D3aJlKSRg86VjqlKdrSh0grSwY4ERIiJjsO113Hvpr87uJz9
pUwB4Ocr2bLyAyan4vMlpd2omho5qbJ71llR4Ku5kMaDtCXpS6eTYfBVZWI9hklAruU8mnLaAMZy
o7p5f37nVbTvbqt53x95cf4s7/Q94iCIFgAlZLzkDe5IRPyw2vdLQBXFZCRW7RpOsr0cDDAcI8fg
0i8rN6a0evRwBJaoMfN74tQUonkKXEl7HxFbD68iR8URzVMIXBlO3PVg8fvYMbaVEe2LJsXtY6OY
CxWhWzFDmNy1fqUnCMfo3zwAP/RKxWcIgbwcYOKsStwSNBIdhNe31/OnikpNJaYxUQNkW5AvG2ln
2dd+J6BNHk3sIKJBj1ShODzS7Cus5q0rhC882hrzMBK6hkTn/96M4IjgVzvY+sPL4KWxWyPxYA0+
qaPaubOLeQr8jpC2+Mcu/VGsgA3FE2tni53h8tg68uPBf/s22eYOupP0zMYByWTGkbKFNLvQGQFE
UUzzpP92Vi/qqOLgfVCszlR7X0VtktUvq/FrCgMo5ee6yuHQkRZS/shMFTVnTMGW33axs4nUX9CJ
lGRMA6aoZA0VHLi80YheqQ9YiwixcKcsBDLKWCYiZdVWOlzidXt9vKJ1l1D8IVMmj62XvFdJQsO3
l0FzM/0Ku4HrKReOsMip4oUf3SxQ7Z9MYyjReru8BUgNpQUx4gj3RJ+B84xfTWq0kxdHrPOmnwTj
9MEbaEl3l4jvrGLhOkAruAIucYTMWJqTQyBEzwD+CK9BD/7NxS0LeNsP2JKCSSi+uUv+NL/BUpKl
osBcT9a0uGBthKztqt0jtwRbs0y+bibOk+d44rWWDq/N+xwdTwfU3cDmCfKr4j9hlkBiwP3gyh58
UMBG9CVjKJpQvrNfPuesnzer6tsCB8+/PE8RRyA3L31TooRrEYcDiBktatCnoa7E0ZxCbcK6Il/X
h3d76597v/UGYZ5r8jg3PvEfTQOdEHmxBU1g/mqzrgtmiVYR2hg7X++ASEofgMeQeRLKmOI5qxPk
Lye+v0Yux5T5+x1gx3fc7RCTJRqfZQayyQuEHveGDSinFte1sAoNRkOGCSw2xBW1bhhdp27ZT9+W
z+zG0maDHmneq0pT7WO2T5KBB8OXAW/J7J+NqA1P70ye0QFwQOYJe7Y2YZsALL9g+ABSRc/8SN2t
ZAhO+V96pCbzm+V+7zPIZTAMn+AVtw0tzy1nYhKlCVtOAe0TAd2d3o3HItclnjAYuLO20zwij3mm
pILm1flidhdyLqCqLl4u2dcL9OoChQ7Rmj4+nBzD6oiGzWtrVdazX1otZJaXR7rom4uyQAySR6sf
sau7L7h7pWbpO+tmURc33DOpqRhb9CDEa6nDljEBAhQxmQX2Z6u7xXQDTdZ81ltkzZSewCxQxeE6
djkfWG0YCn5T/KmozoRXyj7B3mMNA/Gua77WVklHpeXHBquvKkJMmq5ngeB9z7O7CSvtgP1CK/j/
pnA+BQapy3RSTNmc9MuYT7dNdHYPggmzHlgKkmxcvqpTFukBjry4paHfVvVUNSXxVDb6h6VNDElR
oNO5S0OiyzLtLWATZ6P9dk7WD0hLyBir0sDXxkQuiIExHIg6+oNC8A2d/t4/mLmH4AbAOv7GFLgQ
J/Zd2sCMnTGOc8O0jT2EIcN/vexLYpuU55P5jCwR30rxibBJ7HS+wMFWZPZCiFV3NOwgsOjDl7zw
XDKq0GcdTBvg/aEWRIzC+LO6vnDaZWf0IqLk4B6n2ZjqH+QkCmHHtStKBbdj2LXmhO817hBZEeaC
RP4A+2271TNeZa7ZT1kKyXFBeqYM9B5kq+DPHQIR53P19BRCWZm1946cOXAK1rqtrcoph5skrjmV
HmJptWqy4H/znzFTjIE5anQEnIRHuT/+PXpVaMTOKbSctzrCuJYJstT2fGcu5xIzkqL2CRZVqwEJ
K/Aym5Vp5PRQUVPf5YG2da1AxBN6ulS4pDUpW4cCcLZ1Unb+i4W52iAnkquomTuvxxrTBwrmKxbg
W+Uq6BH3mfTBqNby8vylQWq1u7ADWt9MXwQNhFNvSelFakpj/qLYGrpZoYd1mYFLdXOp+CFK6DJW
sE1u7i3IQTpbBy1L9DhwCKV3xIb47Wk/SjYv4ZG843ARIK2rV5n3Y99crTIz7LMgJMn+NaiyQM8d
p1FUcjbzI8+KONb5z4atrX9K9BGJhmb9GP9pLqowcK+fe6OL/Wkj7mz071htLlPI4R/FzBybfwcr
1Ylv0/HO93D6YSSjn2qL3RwK2pr0N/mPx5IT9H23lZVOL78zayvyIFdveUjLJo4tjt6I6OoReJJ5
V+zDsB71NLuisHwxVuK5G+bD9ulYIxuG1KY5lqApC3RC7A6vN9wz2IOI6LvCUPioAG6R/92RRj6K
HVrAwWPD8WeUrIPcaZErRHzClXvfvqqq077nGrwSHw9H63VPdEXyQ3PNfywAN9aXouVx5pqeA0uv
w2hU2sNTIz1ZZKipV7vBJyitunteDpDpNY6DytMXGilaqSKuumwfPqvJGqsjYcN3brU3UoLXG7kN
gSK3hDOkhJ4gDGosKeStW6nAI7pviWV6bXmpBj7voupVbR6zeVNXeAac5k/J9qQhjAnG3/Bg9jQT
Xh//39AG1guy6e/MAnufhkbSs0twY+Klu2YdOCQP6Y8JQ5XUg60Ph9tOKxA6aJIitiZq6d3Pps90
D2AE3d3nGsN/tz1aGQ4L5yToHOJMarI+40ISUOwniqIRirHNLAugxEF3n/02FFMNEtaufvXv8FKz
DYjainzBY92MGsnZwEqV/kM8baPFTiPqkgj+pjoLYa0h9RtxZucT0TCWliwvXRJSuTBuDTv/MCIt
9Xyx7IEeL03C85UEluws/lk2OaMhYo/vDr5GYkZmeEtMfnTqXzEtXM2lITeJzruy+ygAL5HsOvVl
0yFj4ALS/vgpjTT6AKNog9EVI1KQaaCuOXMeZZGb+dGFoM7qVlzegHNbX4oikIGZIfFclqJ69mvo
KqII5E5kglnW4431vzLsy4gArbPlI08lOodfq3gbrK0dGE55elstj6bOkuYso239SZjT5FqiE+R8
PBqtO4CZLtBEDIPnQYJCltdz7JEpVZN9LTk+FlDZM/uSdi+1BewYklb8cQmQGJDm/nTPegQ/gWn2
a/DDLrf0m/IMdR7xGkW9SR1R0M08M9bYuCq3S05+BXz5WiKzVVW8G6N0T+K9aexoSMuXPGwos33l
k7VSph+/AqqEiK2yZZjzvmOlZ5OLrjAW/54OQPxXbd/vHnZFChJv1ov0S7UKWPEti8wyiiZdFaWK
bMB9vbLSYWesfiWBWgDqCX6kRCi37p7o5OEX6Tyw118WUSa8zxebZtf4y6xWOvJ9SjZNEF+wwRnH
wvdZPa2MP+ONADA9dhG9JsE4sv7Pxe5EvI20rRotMuilmGOOqrMpfjji4JE63s4cGD55KQoXQbeU
gP5NcznJzQBSXRjg4IuZ3oF5xwJwO9GnNNT0/VKi7fBix20PWbRL9Bbf19amiUXLh16ODWmeCPPe
5l5mQVhyqtdIMik+vMaX8T7vqHT4/aAKotIqhB1sTZXD+3Ls2f26K0Q+zCg6rSYiAzYEB2SuFhj4
p3gzeJrMEkmSjjk8Xxkr/MzJ/SXv2x6pA7huyqVdlYoYknls+vahKeJTwl0BTKCag+o4u3BL5fO8
wwxELv0pJ0rq2VdUOZDWRTfUP4tU/nCw77c2KDER1GQ5B9J8k662FE25f/bsyhn0uygaJZPFAaOK
1KDVEUVLSzbKr84A8jewL6kONbxtXNopT+HnwuGr33ITw6gW1t+gbFrWaaJnP6z6FOb65CJL+OnT
vZ+nTyc+G6dHngx4h/XhYgwBprJFC32C0y1LaKP1qC3BI2VmIEjUF/N+hLIJFNR5jLtGSdt/IaD6
cmckG49kVzvn60v0DiCaWZXWh4SUQDkxyP+I+clsHdWu2a2VTjsfnvUtulHI/E8B0ZNRQkJYnpeK
TxdThSpwh41Lfq9WWzIuEN4OPVMmtAPr5cMjCzaHI2MoN1oom+8bYcCuRDJicQghTBkNUKEzDoR3
XwyQmdQ8Oruv30HUbkxf+Cm219XI40IHZqDMFlHr15f7kQhh0buaWHpBooyX3Y+2sdr+vV01IAkw
4NSbtg8iEkvZPXBOTlCSMaEONrOmm9UjXXQJB6uJ+nudW/CaytO572ObuX9yt6OkP6zVPS56bjdD
gxczqA5z7NJAsgMyHD0daTbWtFdaIdBg5Ptuaa+xNjNp7tDWEntHAtg54Os/kaGCsXLrr1dH3xzE
XW/e2Hw845fcUZOCTAyczL5i5IJN2MTuJvbLEOvidTfyOOm0tgiCVnSkq28bv5XMfQ3WIhlCz+AP
fg6JAeV+YQ1Gm3XwxJptxUPW1+iSQ5CCbsZ4qOJS2VWcgrhk/CsU19purWn9aLHRgmB3ZXv4BQN+
9ucRpqnIAVwhIy5Gfc8Py7iG5otfzbAAsM3+cr4zXdNnUhqxdyqMMy/yIUV7KwQi1jI3B366h/zX
WU+VG2HeY3qvRwdLOPD6IrRHzX6IMQpPI4itO8U57cPKoLTO9WcoYWE8HHWKNhMyFhSxic7xJpMY
6o3XFkHJ0AAahkn6T2eOkFwtANQsd1RW3XjlCXAlpbP3qtZ0zmVQm6h7X9huFK7NIGe5Y0UVeuuL
gfexv9s74p9i0VFPOfnNZ8ie/OOSqpb4z+CxoDS2yZzbCAhm2LHv2YzKvuAbA+itc7Uoo+u50miy
C2hFgqbfAT9lPwedwN1gvIROMRZlAcXuu+7pPr2w2iTvAgbAlzCl316YVIuI/dhqEF7eDHxl51mO
lJ8xw73LSD98oPuEtqKQiL5DtvrLZibfNO2MGfJBdzN7Sqzfc2y3j/ofgoA+B0s0mAw4Mzr70JYP
mhC1JOUy+j61OFDKRNT0ACJv9GtFwcsgujO5C6fQZeVmPAU3eDIAfAy7be5VHERRvj4bD0K/B2ed
z8ZMqdr5xrQfWYAVPc0wBxqXFPMVr/9YEbQTZ/kcBjyVmUUtj73hTsCtdvJlVBFJEZRzpzDgAZkm
5vEYP9sESmtzEGeAy3Owu4UOdX6V+fJB0lFU6WJwsulj/xT3pVtyw+kpkgCymyXaXvkOGjpAaAtJ
CxMj5yFC2itiXmMhEWS0rwjBY/OCeujI2WVRaQZudHszm+0ahCift5HTt/nidnLoktDN2QRm4JZB
pWRGzFN7yrD8yfs5a+IqBPxNNg1Tfvq1ScdrkNdpX1g0ZqBNFlSLg/UvPpozYLph9g5VZYaFC6Vi
bof6ZDgYI+JTPYJZy7vkqrCN6buu70dZ4f/7QhMYLGH6/9ypKRPTPq7D16KKsTM6/XDcwjSkDp2C
uQao8n0i0VsTLaaTzix5DxbYfRlhVtbZw+xwu36ncJtsdRpKi8+KCNAuN5kO0AxiZSMeuNCt0ij/
yiY1E9rNVbSWkuaOkfFZ3Iv2n6Gp1lAYSdpo0cdLXJVZEzjKCrNtrF5Lh8KPYeuRdNK4p0pXfkYG
Nu2G4ghFgsyFdwOWGJaUymvMzcQmp/QsCjDmfYHSwq90J0ct0wXb1Q1KbQNb0QuXu5LbmRJAqoNv
7R7XqTAsHO8E6kxJVuCJQx17cBuuYlglNiYzbUFq+bOWIDV9WyAB2i3Sx4ffNuvvGhXEXQK+dYhE
A+q4Ezx5EKr84C9/kPgzwE55EiIh2dhdaU2ZFpcB/bcbWnMAMoGQKXft9AhV/CqUoQk8ZW92hIaz
dVMPwlL6E4gOGd2vDvkUc+GtWHrQZE3B30zqnOdiHJrvZVnXmjnR0XiJ1rCUjM67PGqTeLb5cbrg
/wQK1bzsHWlNnD4FTCwlsZ4AkJvMWZQtvCKmy/fKqJgvD2nQO7isB043EY1oeUtwRkWO7p0I8Ngq
80O1gmDuV2y2sbWo35iz5MneeMx41UcDmSxlD7wmzsSWy3MpV03P46hyW79htXS/U68AZNFBIXiQ
bdcyzgYpcWGxd8RrKISo+jnTGpCzHga7lhmiZlLp8RMIOg6Uj/bP6W4RJcBNeTDxXypJCRi01bA1
frkODy9yk8PSJy+QuFNKkFemYdLTXErpskMPiojrbFUKSTV8IQaQWmS0ugVJjNWZtdotkHIKgy7D
dcwSktH0V+R8QyD56QF64K1ZA4bN8vPoIsQG6gL+1CXNzIka7JTEEaMqYMtzRPc5TTJTpAOLObRI
BC5dGd/fCweEF1QLea4ZnEs4OHpzxrfZ9yJ6x+6OLnk1Z0CKE840lmjLAtdy+tGAdTKXheeMFppa
hbnV4+V8pEdaWFl/dJ78aq4zmUkLla66Ore60YkheGsbpS3+csrN/fSDcU7cQ2zotWo/pwZmYQKw
PVgBSRC2DNyOCdUSypOSuOaORFQIx0SNxCpLquMdKCRfqY9aUdltqaEFsckESzK2rvbgZq+dGr7I
risHtGdYqXQS7YzOnFH8SviMbC84XvEGRjEaEKAUPAaOI/kWtiFFBkfjokfMWBW2S2cYnd8wRW9A
bQQDovZFiAEDcHOBqdYKCOgvpn/uqjV9RTV29nYBnpcd5OsMnfxa73ECNtlkz/FOHB0rcP/JVTHN
3SJ7bzbdhgY2KBW00pojAZd9wCtqyKRqH9FXY5YEwBkN2Pbx5d2SuHKA/HnV0cNYR3siqk9fMbNH
uNYvdw8H+VBR2WJ0gdVE/ekDkjwTq1VvKALV9wn3GCndyOebdpvFwiIXg+vLCYftmxVW5oztU8q0
F1f1EyLGrPfL/bvsRLJgTVHr3cLs7GyuSiJRrQ+XdJuEJvV/0xt9NAl7ezzszz1Owva+Ggf22QTo
tpitAEiFaOWDoyQRWjO3oB0Kvo/qFzj6B/bBXuqwmixFz53sCRS5SMs8RsvnbYgCBuaSuhCDZQRL
q/j5dBOpfCayeeO6xO9JyN6t4YcC6FgT+HqXZlskEmngvDJSgH/cqY63g1EQ5zK03DL9Z3IoIOt9
6GNtSTJpkVjH40eSWtWQXXJeMECaX9/fs8DovP4UsezP1afErva1z+lRO5fYd5GPlTqCUU+GK6gC
jMTSNjpuoFsLAecY8u3RBNEQWlPvqj+ainghjapm6uJpw0nI449EWTILxqosKVxC3wSQzMM0VdiI
IT/00oth0t7Bar0AEJOIMT5Mk6ASbQfEMoe/tM5ealV2LFkR1uaLYTt7G+ba1bhg/CFKalJNtfOJ
EOhaFgNcmX7uL0uTmOzMfvXH3BClucWCSmkelpNeZjxnagyPmTle8ZC9EvtK4TWdGDJneg/9ylE/
iBvKaaSekRKSQ62ZjTUOx2IelJBMMZCEfPAo1XXaiZIid8ByD6h2iOddh7L0PUsl8JUh1nve/p34
5EpbX31B0PLvUVFFlwtESVGah5ZWFtcvIuiOpBSCgW/v6YdcdgkoFWz0MvOpPGhuZSU+xQ07VVAp
XyJYcJgje85big2tMTeifGsv0OT0oGKr4jGS8dM4nJWouNnvVxhtTPN9YxlLwpifQsZQBfuq45xx
3ON5TsnNFJAfblwK7CSfKm46oZZmiomHKBOSahY4LG8S9OoC+TlJraBIOFHM2QtE0NckHJTzUnIg
ZUzBPmzIcbyFwKiYTqbvcwkEliPFBIVofflenRUrnx4RZcMZE1gwI1gS2jZnUPxmU7+lfh5LNULz
Pz85VsYIW+B0sYs7C8ojYeVKj8MK4KPtzWh9l8XnocU8uaIQwsNrHOvTJVSlDmwet2X8kq7uzp5e
JzrHO3cPxzhKuiWmTdBtIAMJluGThYiwLx8uhMLJnMNjUvS4uPOuwu/9VA76BAGRdkcuF3kFk0CR
adZzgBntdH/KTc1lWha8j6S3kLrsfeJv5RG8Bi2Q8B0mo99bqJ1eIMizBR9zwgpw+XUbCIwTk0v2
80WeoUmpfiaJ+EM/sN4WkAccxzskWHeXYctNtCiUiTE2v39wfzqmJ02FenX4vwbjqzfwWSx390bt
cHN5P3wJxqC5ifbI/RuBeuGcZyFQSFFm5s2aFlZLvCxhbeWjvoUImHyF3B4bIk5AeykF/Y3E/eEh
70tAxWxUEYxGGyE+9sDYWxapxdvk754LJuOJlk9hbvtSMYUKKlc4Cjw2X6sHrqg50LcUZL+teWk7
DRZngUjU9IlKtaTTbFuUQmQDIibD6YLg87B69PFDfdWR7R0J7ZmffUHSXvrCr/YCZsGDJ9yYy2Os
emCTVfW/jc/3hJHveJ39+pd7O2Q1ES/8m1hr3QY9caUXFCG16AytsyRvFVgkTMW2AExMAGLAkA69
Gxum2GFoXm5QmuHCMWdtmcGQyA9dKQLUQ51lRoKhn1KOk56gYZedPgooUedyD7ce5ZGrjag6+tEQ
iDlRik7MgHIMR/FS4kV8EvphewB0mynRH3FQKr3RIanWuCYdpQozo+c4GREDwwrBpAqVguuOcqbm
WPKKViGldb9wUMOiotbTVDjtwSHLF9392BeQ2XfHuQ0RXcA0aPkAeylj61a/Qcoko6SSCf7rbYFX
4V8caTnD4cGfz5AhrApzGaVEU4MdU9ZNKiJx/Xf3/IvEb1rGeQS2dSMoVTDCNgQQgrwawz705lMb
HzNJ76imzt5pgzBJR4juw5Vm2UlYoscKj6wycQ0V8qAw7Ba5IhtzZl8U1MhbdSl+dIDJb51Z8y8r
WvUbMboOHxvD/VnUjW5np7TIqbXNGCkFansRKVeVAS+iRUL/fDRmzE+ZtPoX7jiGgGoeUGylzDss
K/LEeKomPu8mYu3gKzwdmspKQ+7axyLtalkn4DoILxcwH4gtVAUHnz9QSkmpFOJefqCsNMjpIizI
hE3mZfDZ+i76CxRZaTnKekl86HgY5B1OaZmeXHwEyT2hO3OZoHNYaVOP0QXk3GLL1AynsiINZwrx
MxPTQJFckq0bQUxbZYS7g1izs33h45/+EXE9SZX7DuQxZEBmQmoGsoDOCKmM7xFNy1E945jnz1hT
htuL2AvGlMcm5x26MSidhqWhacbTbjBq6OcHPvjN8EEjvEwN/Dm6WC7qpijS6Fpzj5zZj5zk5rWU
W+pbYQH6+OSH8z4cCK7ippsh2kz5rT1VdqA6tknjWmtfyPQbplswjei6tIoDn61wfRqk2OOGr+cm
SAAre1RF6or8BH5F4IlHLQ9AzP7tZUG1QoUS1UK9ILz3vmzsJdirHK6JQ4FPNL3HiBzdE4/bCkOy
Hmyh9iSydgw4L1NIYLY9BmLWJ9mptmdCYPdKMekKHt8PYFl2zFegJsnmBp2afxP8GmauM4t26v5p
DshfAVSpWSyEehhs3La7vPfNTXIloKArrW1lkah+KKrWK/y0hS+kK7yy9agX3llN55swYZRinLpa
AoIDhACHgG9JS0UuhltaVsHgtj8biREyEpXLDkuZ8epTyhE8pRNyHJ13vOtK7hErHBfitPTYUlFF
zbJEYmrxQGxigBmSmKrogx8mzdv3NXKG2VmJHYcecUumf0rvCRZdsosz9CP27cueK/jWFvVw4tb8
NS+uAV0ekaufSgutaIbpFDwLm0c3Bo/RCkW0FtdckxP1l39y5mLvnToEOOeLfXaE5V9CEbf5T7AX
b+ojbtFM7riC89nZZL+qdb/8iBWtFhHf1/gOA81cSwq44RYG4CwZgL+1awMdPNFjI3Gj2y33LPv/
O5ld5GrdvU1Lciqto6HI85soLlxNHKhDraMQ6ZtmCs16wyq9i19tp0+p0b5F5jenPKoudw4ExAhH
UzQK7dIdQK5SarbXZ2TnD7a3BcjpIiuq3thlWfKflDDOZNakFPcXlosqfhTvMhk5bsYFaJ52ncqA
4HiECAgdQHi+6zNuL06FZ7mbeCvzONacy6OrL/tyOcxKKY1/tCD2t5uYikp8u3Z8mQCuJ3iLciAu
ZqqIaxBEsDvAdZ7+K/EUjEjBkkKr9poLFHwwMLHQLPohm9AHR7a0Tgtz8pFeKDa39F470qsRHr24
r8/cCsRo9pneaQ9kwZlZO3gjTQSb5hgcWgGACJGsaxr25SiH8ucBR3Xzf389nSnkG9KA2baPwW8v
bnAszLOCAumlULRveDiGSGMBwrM9B1GURO475k/ZPjXZiG+ctcL/xOnhnyRLSUvigCWxvuXj7FIn
cQT0kbquynonvEa37euqp62q4sCbkNfZmrzMpM7t7emMbTtQgXxCg3ZjRG5Lf3kc5mEspFcMjJc2
H6EIqX3rtkncb44Oab+uzNGtCuFiY/qj66MJyBCFDT3yT//ceI7B/2cHySl6e5wEPTr7jRMILDGs
gqZ919cFGXAEITArpkHljbriosd4niSxf49uZuqzLeeyhUxwDpFwMnbIGxt1AuXpP/EVpOXkyyWX
34WTW6MmjEbD+79UUFLbAjxFfppd2z1r23T6clQXWf4K2gzBHjICEBqb4vDLIoS0bGe143Q5r/Qk
gIxfegSJAJ46lhQiGAJ1qykfsZtK2iiTQs7Dn/IYrqrKI9N39iqH8uHf2WVGi/wWHXaNe8uccxjr
MZlBsYIJ5Thq1EgHVuibtpQKKQ4z9+sC1tYB0cSgQxP+EsOBvUIUZ2zIDnJ6sXUc3nOpZXxOIRv9
fZgNRo5tdLE7IJ+Eeth8ElQHyqZWaM3Qp9umai6Vn4YBVpDVFMGdSzx9y8okVMKh2/7Bqz0F8yOn
9j75hAvXo3DK8Gf/cTW5vGp15ChtIOyExdQoillgReJ0XWo8i1RVcZJGkmi7up0i6WXqwHEJ67f9
fgS5zmO6vWl2WfIGwlvgVFSD5dxRQRuwvaJK5grfKsY1e6q4QMeTHEbWhOSp6BNZtEa6udSEPt9j
90DHGk/R+Hk50eHyMUCcYXp2/eh6lMSbVrXODwZhrKc/V2llDiuTjrj8p2g2ECVg88rY2Nlzgdgl
L/kP0jXcrTpt5hj9sr9wzT47yvmKFMmrWO3Dzesv2nE+66L7f8a6nGZtUEB6X0hau5YFc7BRLieU
5t3WzQ7NK7z9YJpCH31b+1VbLL+C3ze47q0tZH52NEjZyuz2imEGHmQYDrSryIL0lX+ll7NS1FED
tUdQo4f7RuhLhVfu9IJoCv4160oF0/GZy/PagnDhDrSFbB/tbDRssOtMf25MpZ8VsAt5zVUDRQwJ
G7sHxmdMOZVE3A7IlCX7uBOQJWoVZyO/9MCg27kTrAkIPUhl2futnodNxtmb7n+QPIxCzzaDQHMv
l8g18p5bXz48fqAZzVQmVdVs/3w6GrtJ3hjb3NPiLhs0tuw5UI7HskfJUwy9EPVnbFUNe+EQD5MR
rlGVl1TXMBsceF4wOax8kuefK5MFPbHao/VLLxP/vE977hNG13aSrapWse3aZbXe9WdL/ythgwt+
NJ6ueS3wQ4WfWShdv8Eej7JNgDghtYuQFbHtdD+9MKSsuZTJZSARok+1n7gsiRzrm0ar+Qk2G1lq
a7scXju0MrN85rAG38EmSE8Bka7vWv8eTh/ST7hopl0oxd8K8lkaTcITGGp52b88N12N2APwbCuP
QrYDa9bHA1MToVfKb8204pmI2TtaiCHHtlQ959KF/6UyzYilkW2xKIjrpQQpzSFFYgavLiOq/GDm
4zvivrJb5QVAuBymLmTMaleoufrQvNzw7qSpg6507vlwH+36zWWdY3ofX9Len7ZC1prX68PdaFWN
r9vu1VvdDbLR88I8KGQEc5xLSFq2liEwPie/FFYBRGMPWTHXBLHtJ77CsWqW7D7wsPsb/gQikPTL
nv5AwlZNYd0VmtR73ylM3hRdWl7RbBvZ4Q9utF16rtvNjjdzYFVPuF5p6EXO2NRnRV1ZF0Vk/p0p
R+Vd1ad+CBnzj8fZCi03nLn9+aee83mPiA/7feJESuTySQu5OMwdgiXULzbI+kWBevmj1xnXcuU+
187pdDac0OEP7UMD2TryNXN3zV39bXCKGP/qXdS9ll+U+YKLm0/zAochaE3L9UmXAJXtZPRjOsp9
hR1z1KvmbnqDlufszTQT0mdBOTnpOX9JwmoEkL2Nvtl+6DM+njOwexuPUFPRzyAYRlYNCONVRU+y
WQJqEc0zbUPtQAgZFesHv9jn6lJl0J3v/5S5wwfBPxC0n3ulLRH8ZZZWbGuYwh5vcGa3TMV3Mywa
43oaMv+WBqd1U25yFBq9DrqW0fdlvMuNcWAr46xox/4iVxbOXWG6hV5bM0AssM9FHc+HfKRMDfK7
yWz4AwqzQyZ3ZGwm+Qf3l471iJXnKCPDFD9xdwLW1Xx8laDHqJEaxYFwVDItscQKUqZjNhzhKUZD
NU4KnLAC2UBYzCknFzDq3Y4gzM4PKXLLpln+Y7EiNCKoGXrwg6XkTeppp1LpFMpHpJrbCQ7nMqSO
lXAEIGmOwZoVjZVfW+i5XgIXGpWXAN0JZs9wh8POXEM/zxJIf0IlzfOngXeXL+IwvF0RRYZm7ouT
FpoMmVqizof33iY8rvfNT8icsbfsyXHdYQNQZRt9gUCL5a+seruOwYD6vveu7vtPPaG8CHe4m+I7
vbfU3Cc8Xh/OAK68GkqgDExnBjP6IFvopjLk57nZSY1DSlSwj6Y0tykJpPiYYpmn/RYx1gYj0ahy
nJQ+VlgpLS0bte/9M8UwTYVyADXVotN/Fo5oelAzXmOKVflvv/3Hs/pdn70TO54/T+ZWdxFpfHMJ
rCNS2/Q3GHQszPbzy4irFsbN11NcdfVc53hun3MYkeVphwM8sv1TpUc14gcpKQNhwgoCAx0tZy8R
RUaDfeqJ08jMfCeNg/nX9JfT5ltBemyt5cX/Yzi4vnwkQRjgEcE3Xy1aQEXeqUS0jLmsonRQd7jQ
iy+dOhUDuVgme0qb0aXdq3eZr+3j4GHzsSGehObGzk/gPWgplT8+ytKj4JBHhn80a9yXpyRmvr/O
ZmF0Gse9DkAtzqgkqlOcf78+WNOonSIBcPU54MPNcK484ZqsFE0pAda5fcV/F/9QuL3HRyZxo6yA
Zottnu9+i/Gv96msNmNYH3LAesjtTpclPTNlMzFFjI033ASEzD7YSVOPgBlM4CB/fGbg50xSyGd6
CZReoi/kJ3pxQb843TSEa138N10kPl/6ipSUUfjyCEXCnpMFPibt6P9dz7KV4CMr9xhd+0x46w+4
1/EUMFLSVjQoPo9BoZY1SO7u/diLhAmnDHDTv5kIS86DXjzP5pi9rWraFwxNUKzJKy2/CbptLLS9
0bDuGs86H2b9Vq5F6Q0ivSl21iy7nQBDF7VNQrRiqI7FlK9baeQw/b9MqWw0firSTcjwadbpmBDC
aj6rq4nJjGeaN4eKdW5Ha7c5XYlVP//U/OebwI5I4LyhkblDhXau98tpp/v/rwJMnZGdRWcIw+7C
NpBIKnxFZ5k1z2Yvotkvfqktp00sJ9PeE+PQqFSjNE8b5UDbJNUuLgBfZ9hgbGHMR8X6zHRx3O+K
HAP1/aP2GEDI5HGhX7+Y6RjHqWQ5fw7XP8b+rZs9nLtpP4Pk80RnAxTWydMWl8g/TztGoex060/o
QUWst/ChaVZmhcsyHupj7eOTJMLFFaQyNMmduPVSnD4IOCfGw7oE92izREgAXovGjjGm3MF5VsUC
5uQ3Sd4sMDNG3NESgcj1/viVVJBWWw5mzqAhwIL0n07m3j5Ir710YLyZuuPVdBMPlbX6SkvgxIMo
/3AssgaRCc61kw7HBGKD1QdGP0YwLNtrYWHSjPLjd6XC7aV/1dODue75M+w7enetTmIV546jsWfT
LyZTvFmm56/f3mWUmnpImLFUOzhIdCgVGmZ7ItCtTWVVBPaTfCYtNAscDAI/PqDTCJLpc49r+2O+
HArPcBeMwi3hVc5bTuzlBU5uSrJPx453Kz4Z0Un0vrv3oA4bv3hjLPLxFfg+yE4oc9HHYyYC8Vmc
NffDv6zqjLJaKp1PowWc7yEXC013fJpX6e1+4a49rrheGDxo/RY2i6ex8WuWNniKopv5Fr8ndRL1
g3eZ/3SBnvu9jKLRnPCPbf5+9CL2r+P31LW5PAMYUjkSzmRLEqqmf32L7DzQ4f9JtOZj/v7ypOwd
2oOyL6W5oOc+lIXLiNBM5vbzqVLp35UGbsdi+RkQys0NNPNyyrzeixXKC8Q3WavAXUaq5Nw5xANo
cmmWzyA7X8iC+E9euRc7y1XtV7fqN/LO5c+L2civyC4aVw7i8wqTluVeR2EPU01Ll8MfpAct/8Ch
0kDvMGIBs2wk89VwMeL2r5CKOKXERQ/KJzR5+oFGvbl4lz8wKibAOKuQNYwGoM3KACfUeYRkq7We
sxyqMZhejB72U0gyYF+Z92EMx8P9w4N+FbymEDjCR5GuRh8g5QQ59s1acznIa0Sp/UhfEeltlVRy
C8Owd7mldFN8EyH7ERcz5NItmw/D6UnvGa4FgZ34VSJVT8J18Q0oL5Zu2nd/Efnz49zuA7o3gegU
XDcMQ2StscrhYZrjHoi2fNcQO6+W8Gg14JeiSEuO7jjIeKwKoZHsYjZTVN5MVo4LF9inOVuHKx/5
q9/MySLICR7zb0EQX0sRxDHSY8AN58dpBPoM0yxjgAbl5FaOa7FfyeV/yqw3sLf+ZBJEoeHNppUO
cHfGvuKDMjcwzf2IUjvoL08bFbpxqg5X4xHeOL0d/WukCOHcpGejGw+Y9/qmOCDT1NhE+wgTTKcJ
D+ZdLL9uyeSVq8A6cE9eZGPXYmhkKExXOtBSH7NDQsZ+5B15PSA+374lmh87490+qvr6b/wCcAz2
hKy3VPrqGzj9RvufmsNs2ORBe6zaZajIFBGbdxLMyDY89SBi/mSUeZvxUx92DekLCnFU+WYxAYAL
RkMWxwOZAWrLrojo8V9ClwDq0d4q2F05LY3mE+aAat6jkyEAe3f25PJzNAqW915p/9eraw/CR4HW
/RZ7+KU8oPDKHo+no+i6ELMSQPisPUO8kpoWCLkWq6fIvolSZ0SYyiCNNh+2q59vvA4G/L74+Wfi
w1WYYaGU1PQUcEMMSCcvcuVXWmWdzjhQN54cqWXnUGjILlkOZrr2VvnFhtehd3gcJWyfx34TD2MF
xTLBNd8oXH6ZnEFiZ09wu5rOUKlNPEOo3idtaE6TF1ZgzXV5QFcXn8zAwqgO3fD7Qt9R3w2GEndy
DFBYMt5GkoQCOmO1Yv4nMwaRKzJVC8WmKoQDWjaUOz2GP/BTcenMAlYIvdEAquRCaLyKJHBlQNy9
cE9h3iLARsK0BLagkfMtbQG3bzQkkJVmqiV6TWJnPdT7PxiDxFG/ueTbBr0uFc7Cy1gxyZXqxi2p
BWQLiXUvQLT6Tb+0GavPr8+mOtrv9NYtkGgGWvwe7YIs3e1RP14dYGk24ftiXnWCp6J81O20NQCQ
5EMGFw6bAVL+V32Ae6NKkRR40V51NSJ2qUoZoDM3V2wsVDorTKfEOqsz9lMRwqKn3todrvWovYLh
wLSagwOCH1COWwTOdJt4o4APqgycH1Cg5jtAttFe3xdYFU/5GclTFiDvQdrLTM1465NOaPjdnXh7
UTmeqEecxkFnIR1Kq2mTn0j8DOAWH4ErCDB8Ki+x2V01GZSUFqiZebnXkJi+ybbjy+7T0eKkAvPh
VvBAkYAVrAl2j1t7I6yuX8Cxbf+rB8v7sRZI8mDgliHOQkdwkgaXSeKwuv2V4lOW4EnhX5pHAtII
H+mGaMADDBzZnVNN+f6bcMs9tLHcUOdbdqvTaYd2FVrsoZDguFFk/aspUK3fKVPkR29QPOzF9jVV
KGzgdAZuMKJDzUTROFO9sIZ2rACARydQ+qncAt57KUVzceFL8DNc5/u8n03ADmwFAVlGldEj66FD
RJICWeCw0y3Ic6Qa1qX0dMNS9bmUBFAm03saZCWqtryUcUhRhTckZuZGZuKZNcIdbuZqBQ3rvopN
kWoMg6zV/DbdhtPZ/5omi3cPkId1N62uuKAhLw8bwwC3Nx7ZU79L1pSqvvYsXpy8dLcZREp4b/Dk
qsMHRjPKYrs1TszABmkqgUwBp0rQmgWxIBXUogfkw1l+V1V9gQbunT2ElpNBdK7HaEMpNR3pSdIK
DPeoWIIYBR+4D1fTizTsi17oCsjcGy1FRR8KxbiKeOiEYPtq7AcAgjTU9XuIVMSmpzpQ4JTb0hf8
VGPzCXkPzKJwjuty8swnWUuYoyUqp7P6HIIvfkWzDHgljVNPH3wIKKxBVwRjttfbkwdHJZR8uKCn
vLCeIo+b3OdrLqhfomqojiT5IM8zPxF5O3iDzpn3rJzMlFNVbqktd2/2xgWkqlgd99HSmCb20DD0
R4CqEYuLa0F5dJU0PfMgoDyUIaNS+sEyzdZVoqKEaNccnNdo7bKkQr1QUHsvoHZwoCEX57YlKkwN
h4rAQziKfHMI0lR3unGFCToOKbBz5OhTgUb8c7NlE7M8OKROe4zilJkTVJ1EqgnLEME5bXRLxD9f
CUd621xksCoHNjOvilGAB1PFPpVZf8bQ0kqVLLXJPiixlYpEdYTfC/uMuCyYI1G/CffjSf0YWxxv
XVyAfsyqwYS0HyDlWw9G4TeKKMNnGrlu+vMkLR6u+p7PbfDhUipwX+b5Fu10tS/qfKZByr8POhtM
41v//f7GT0+P6RX6d0N1KKQIKHu8i3ZWWe2SdEA6xUhTafwJu2zzouHvlDSBmBgXdBXIGP9xBCoH
+qgvA1nXikKAlDs3LUjcKrmB6166amTnOUaz/37nGeL+XoXJjjLHfDViQYieJkoED1LcueHrQPnl
pYA7VXfXGzqd7NDfwuoZ1OBp4W5yaz95hZVbxzNK100hNcF/Np5fJtzzHGS3Z1W+z5sE0tlXJuwe
IoYYSVEhZ0FeAobmAZwlEK2FgIPkkKiNQBurRn53VwyijZBz2aAHGbRBjfVyMfRAlUCalsNR1VYQ
i2EhaFsTKRKh51XSvv4LBrqfIcN5FvDh5H4m8wtDfB1U5FXP47mu8p5kPZWIIpfNmxlGwE2XdFdM
unctE1NWrzzwnWvEcL0y00DLf1TtaapYe9JfA255tytKrMvpv0QCU1EjPBqwNAoy6icMyUKTViHI
tSClhp8KlQTGP9o2KsKhXFLgmntt4cI4dn2Lc+/kPN1WFoiUwb+rtzZYup8ik08M1sxTMqXt2L+V
q66sGMXxK6AqHmzqtASf/gXt1NGwoQ4LtcuUPuQyNMmm5EcsHKG6jTyFE2pHrBgWsfcTiDaec0Qs
/HgX018DtGLAjFugCOBeWHUB49EMBS04c3UzqjbyUPcuIIySbkTkdJ4nOWJ4/q6t7zfFiv3CcIeG
XY9OsC1eDl1/jvE0CJBViZCVxPmJnEC1S/CP57sZQSC2ThWnWU7cwzvfSBNgCyNyjHwisZ/u0A8J
q8TQDgnFDSw2zQSDj43o5RncXgWDc9mAK9rhxO+hiJ1dmv34oy+UAAADQryweWBgzKcnlkngRyb5
g6f+MEKucDpyuX+44spdAuUHjJ68hFamVYI8NZHdORHrOcaqGAXUTucdH9OGCQsjheRVK4YAuYtv
edSN0FgVUc295Y3Y47EUOfetUpBMCFn3RhhSEcknECcFp6TMFnerTmRWSrBL177edFCcxC/LuY2P
L/ezcQ2q32QpNdjKhpGnDsile4ZeiR2pK/xt96kVcVOE1ysypbKLktnuBokacsuoeA9GMHYBIEGP
chkWx6puzPgFuBYJ0aZbXUVHTKid/D/4Ajs6j/iz9QNprNCLDcS45pbMIAxSI0uVCvlDkqjfqXWP
hYWu2Bq5vcpkBh8d/d96csYFdUkcuD2gUSsHShW34BJAeC+zO1jItr62JiJn7rrN5okaNVt5IU59
BTiIfeC7PAMk5gE9JeB2MkgqHJBDB+vJLOWGhAfe7N3Cv6/ILWNfBBdIDw8s7naLIzppDOs1F1i/
TgaH6qWxUImq4wB8IbsrZKlHvp1Y63x93YWunDS9E/NcvqykZW70NMRdk0GvZ/ZnpTaOtQo4tEtI
5ZkszrFvZit4wGmReqVXjAXeo46aWqBBA44nsYZK7NwLEQbDBeB7DYudSErmk8uAmv9s4DYnVeyN
zle+EpU4OFfK0GWXaouMrKsbPc7EnNo9MoC1BqcdcYJ6J24MEHBN40JT9mlknmJFptmtO+4ACs7b
bhL9qNdIQbD6OK2BrQbQjtcJ0j3TCxuyn48UCFPx4T/DTLidanHljv5YM2LYIUvtbH/A5V7RrV5g
CKBltAk8ZlcMZvlHDmnE8pVoDUSnWluYfFCyqpiVGQPKIl7oMqFmLGvjUNeZ9sh1gu2rPF1VeU8r
duG5ZY2IiWOtQtKa9LFJclNYAdjXrXijm37l5sY6TTLm/i61zF07iO/SN8VYzd0wPTgZ3OuPB626
EffDCjzw9oCLgtl5RpmSiYQkMejfh8hb4NoXvts9pUIKMEmUjxozV/qeN0SP2cdLScrHFNKn4Eiz
x8KpNBIMEuhVOkedQs+x5L7Y4iNLAj6hT4iYLMu777AtYA+uBMA+1V0ujtZaE5uDhXzPwzAm2P2L
9y+GgEmETdlm3MPjBuxF961gfDxanOIGkkVzNcxw6R7zDm+REnAj9Jw3M6zRWTsrZYsT1OLTuX5F
jhHrmWGCF+6oNmsspNfTDVpuLI9k7PwPG88RQrBXNw3j3/ki57d4XjBfrG+z4q+uCOjWACZyoy7Z
vF6I1ZjkHqGxkwZbptnlAj03fQ5Np1MKuXDHZZsP4J64H0W1DJui17b/pihXgn0OeO9j8zix8ahP
ukconaBPYMBfYqDFyTaTefFWx19ARYZ5TKCshsYnV9kuTQT94KOHoVeP5BhdU86VvhHKJ8uUOGFL
rZ6JQkair7MKgqnGnc2PINMaTIqJbDNt0niTWsDQNq1svb5ADCxzca3cWhi9xPtxhsgKUZiD4oaj
m3tx197dXtcbJBLCfIkea8g3bbysYFkW3IrdRym4oX2nioP1UUnirZttgVJ/M9JRGP06v89+dFOr
lmD3X+OKqaKQxK43Iodx+4pGyQADujBmpGR5jUno8YARrHLzi2FB1R+V7jL4RNY8l7AgCsIf33Bp
D3EpStjMsVVxFGjY6RzZoPou7qUiDzuVf7CTzwpwU/5x/cZgD0v6Qjs64NpMFAPK6CvaDIaoljXC
fM1Unv0ornYru2fkfSKhEZxacYsZnTQe07LBjtp5GYWrvYvQyT+CbKMzVVYRKCZJOHv/O+JNIXSV
m8Jz7fPEhwEODKAvQ4p0y1kRve/IjodZsimDp/0UqrS2jMpFJboH5qsalGiQpe+UNRwB/LS2u+gL
W0bofIFiQ04loUJ5yUpidplPh37eJO17R3PyhTYA7bHX3zwfOtWnO/mqr1ggJjtQOvH4Ubld0Xzd
cgdM9zisnW4LCtty3bXWV2FjL3y/3lb0/OZoM12ANcw+8CPvI1lcPwJtYKyc30swJWCXVIdrGTHz
gznIro3OLgY7noBYrPhGYZb4f+4/MVrDbwTNFeEPvZo4SMN72HCS0d7SU3ufWHXkejvV3KH50a1O
dSloGHDEOqbauI/xq3IWTpUCUCi1laCsnTBxVfco+LvFDuMBgfn91YwcS3XeZ3UZdL0wKqL2SoD/
PhwDPJn+Umk++OrQWPgzzusG7n9EOvqy3RDl4Nne6Gyid8Akfln6fuG4KncFw318vBIH9H3NPW6n
xqTDBVFZiMbNs2YPc4Ep0dMqgQmdTkFiWj6xyAfaER8/mYqFTz0SODkK9A6/PNy7rHqVFNhWKgEc
BdPBuyPyes8WSJCLU8Q6CtHAXc+uE3rN2Axg8rvdnjfHRHDiAkAsWuIHO5cUscr9Ga1n/Ez73WFv
N3UsRCtn+iKIp0xQSSI38bK3KoVu34dvV4OxaCPgyNdydtlaEXaVdwR1GK4la3vIJJNxYRs9LImb
NRIKR+WilwfmJg/my/gu85SeYtZ0RZSk9S4+egxmu8WZuojOMX9dbdo73jiAEFdASnPbQkifmlbv
aJor0sLwYDySotFkN6ZemQxsWksMvQA38AzEpSI1QZJYL4YbXjAK+Op6h4mt+8Ws/MyDVMxxOhDz
GuVS1tX7FNw++uuAQBq4KkrY0GMHMApz1EvklNU1R4r7XejEHRqulEfyYU0mdRM6jM7g3bqwFr4Y
A4kx6mEEajQGUA9AVJ6uMlkDbzzjzuTrKKqfc/RR5e2bXPwbTVLuA3pdpAZV0xWNtwTkyVP3OkiF
OpaGU3zA3VCoxbYlRDMOHO3sLjPS811JXOogVSebF5vRvS5drphm0SxfqYTKXQdTShBoQNFRii8a
IlHMerKrzN50B2llDCZXAQ7KceSWmF9WHSE3F44ewl0w45YxGWp0TNc6R8YwWg+YamvxIn4OaeQt
B/ebKS3XG71w9dQ9bydPFckyFULnw+uiXLLGC8Ug5D6aOtC6fbQuV2TottAbTN1OVk/qYEDPKPql
FnjWIwMg+zOefmjSsEt2xBKGKLNDrwVzZnp4yh8qgF/BReQBEM+lzdexpfN0SyvX+f4Ee7A/gSIB
O0HYENvwO4GpnDIlpwTLM2gVB2vZu4zsQLr+xfkfqo2LKU2oZr4AK8HYF3aNiZP8lQldXuI8ffAM
CIBlF7v/XnE988M1ij9kJJtVkkNB9XC/1/UZrpkyqyOfli/zdse76tEI//k7EzvrfRkR7JmAq7nV
XoNfA2R+SzArjWJNLwBjB9CnSqCtI8OAPMzLuX9gHkJ5l5ddPhLs3aURwa3nxuMvZnOqarLa4NSY
zFaZxTPxTVnJet2MNQZXJTzh8XmpobL0enVOw2lypwYq0qpDFHBl5qCkvWlxZvJ77+jt71PaJd6H
lW09zXk6Ndd7YC7+d0CTZoTH3bmFdqO0MN3+BdilO1kqkpjZKwTOiT9fLRpejXRrSnuDJP7bKj1D
RXoLWSt2RavaQmo1xLf9qgyJPHu0TgNfPE6xDC+qwrZv5I3RG7qy7uqy6Ols08A33eWia1darIm4
pKDOR9aQDzAlrjUjppa8mc+MjjvRFLCvZsolmNj5nZ0IAZP2mj7oSRPK6ffgObXlQibcptVJXS8Y
u+mxKud4SIvwbAx++TyH52998DVavMki+sPkOqCoqev2SVj8ptlGvXfzE0vvzI+qOeJ+JPKdSp+y
GdCxUu8B4m7kLHZ+YgYCuw9dxksOaL+Q6E6p0cemeWwTLASXbc88PeWwuB/q8P7tNZyKjPdUOBab
UISDXijpKX5d9zQuOEBraxC7OByQNJrwS2fLvzayOAY6FI3s98Hg8cKXVodLwTVu2qTctPbAqrXL
cgIKgjUkk+P5XU45Lc8KA77LNRSfifBxTyqdqpJgokztnrgTEX/Gexccunu4bXy6C64LNrK/0T4K
IAMhisvWUtFBJL4wtq3ZgB3IP8KrhT/NI6U9iQpL9pKjaQZeTOv4NoNXWYasUGPkYveqPy7UEifZ
Xbaab/DkpJFnYMCymlSmL6fw6V48aDt9N86pGKtf+GMIu7FjqsU2r9G3wXh/vnOVHYG6ami4aZ3e
eAPBbxMbsVQmnWiZLqjjalRU+AoQ4qDl9Bf+FluMHO3eb0OqyPcmfGesNj4K7dGEKWLA0TbNycsZ
xANWoXbtD30o6AOwPVdJbhx/zDEjlJv7+tEKOE7RECgiJpGXhfSoMLi2ZGxQS27PYt4Rc+VedRFv
gEwxjqWx8shMlnYFFnvPEuDih5YMCJu0DBZPYYk0VUAhO800ZF62Qotii2+5wkZ0XE/+/C/m3jfp
jflrNKNu3XpFTn6DGDbGzdRdH8ztJpCkpVTnTLxWkq07wVJsATBLusr0JuHzeI7f6vvvw5/MUyfa
FHP1RAMDw7pRCS6E+QQaoj3azgd4mzUU0PvP5AgzfhK+ziNouiM5kvjuKh2UJ/JQ7cHXH8AHmiCN
WWk8pD9y34a3QOKoZ/cJzq96YjaWvZh8FtgHm+6W9LJENjmttgVzI3x3xnGbGBkPu5DW9tnM+K2Y
35izVyWDMq30dZRpfY//svdccvQ3udlI1/FyHIWayBWUwH3V+KoAsXtggOHiB7D+/lRG2d1it+rp
Ztk8O1q9eLAgICwMH1hvRU4dB3ZjPnaWmVy5moId2Rni8qGlq7pUCCanG+2QAkpv4gYvzKCuO5dP
Ixv+QFhge5V786CWC3Za4Bi2ZaGCIw3r7jCv286mPHsXW5DQS9cFbs4Nhqb3zLHt7j6iFZFKyvFP
ZoWPIfRFJoyTzt56h38xv6P/p28ZmPCD4aXkG/J8U/+kHCpq3gmS438yhCkIwPBM/E+Dp4n8t+ay
aZR1TSGEcKOS/1Hz2wFd4no6z5Bgl1aNAFiCH4lDJaAkeDnRUEhuFlplX3eJdSawb4jutriNvKN4
lHL90WgvMg8UPAZdivMVmn7lNuMkjRhCbOUNLS8V6lw56o8wH9ANXDIlLEUp3vwindnFH0jn1CUi
JQ0t65ig7IOVYlDS3dqlIWICdSmgHJLQGJIc6wmrFzQWHofuaGP72pT8P0FrKR8Xacj2cCzFDH93
o9Lq5GxCxE/JgIuCLr+OjhUvf+oXZ6QOIktf0CIA60pW5zk4KekWcq+u/W98fF3PHnZ025164n9l
h5KrFGF65GstffYpICwUx5Cq/EvONP2ZuS3Egv9+iLDlLR6JJGsZuJrnj+dmXNVcsTgEP+jWVLem
Ie1R+QEzv+0o3olt0dmAOn/LH4G6xVo4owkU90AGhP2hu4PBFFZPW3mu0gxk8O1fUNUwz8Z+5CX3
ZhQx56b0ZxeyAgNNwankQ6e2Jx3t/XjRJyIF3e3MhOKJdL5cLPc1WbJINQVcqGcuyoNJgYv34XYU
jw5Epf2RK3ii6uRBIB2VMeTLKhHQqQ3jrrU9N65uEsarsVHGBHFC6ijEyWzb4m9gErkz0NUbg+Ty
Y38b0FygPNiAbqeX+NbGGH/B5mGW8YQHROOUYaIKP169jNi96cDZhJ+ivItIbU3qLFYGyp0CgoY/
Gu+hbCrmZrXQBNaT3uGwTijGwuytjeFxNFP34FcqhEG5TnvrXRdRSOAmQSErW8eRZf/REfE33HXO
J1SIfI3uGr44WcD1FvmNrtMhjcJZ7e9g8lKP2XMqzElHe9PyGC6tWLp6hv9gsZIStBU0bXY+AF2k
4jrOCcaBV5bfCkior4+bOVOH1OrYg5Xywl6HWmXGeIlIl0awCJEXynur7PXDLtHgW7WhnX+5qOZx
69lG3GltTuM0buxsvlCxa/eY/OZs8aItetjXvtGcVk/dZ9CWCnTfjWUnS27wE1QspirO5EuXM70F
oUuOPdI842LGh77H5HrKZkqukG/DGnXyejzoqthA3UpIQxfI/PBAM1lz/5WlAG6g4JTbmL9hM9of
eTLNSI06xwN7NGM/pbMM4NV0Etiw8YPyjk/ASysCKzVZsq4Sz2laNnd8VOu2mXhb2HdLLQ6o9y8y
Y2+HVLQl6wWYTMLJp/vlJpyaSGnntyOs+QAqjAHMUp2thVcQZMFwaL75xBnR3E9hC9XOycWUeJk2
QTDvwmYSfotyCBAC0AodaeumMxNVZow+IgfYUs/9nXrY9ilI7dwe7vxI0nBnHJE5UIZ4hDWLXFam
195RnqnYSJ7hxyTYcqo8v5pdgBzFvWrzlcfcAXZAFY1J0M4nTRZH81wvLQevwdkQEZ4iplNBvnxb
GdQNBwZ7ysLOFzWeuMf8HevuatKQ1AJIDWZihc+o+mW5eZWSsZEGAm/YJNjGoPKAewUluZnxZGPG
vGH0OHE4Dmi7SGiScJGGpnOy8V2ZWgGG4xLSwAqLipKz3qBYQRY3sJeMEpfQiKgoJAzsFys0Kins
3Hswfps20xE8oh606smNR4km0byyjfXS8IP0D+2LK4i8oSI7XV7b2uluO9SEwBJL53kUH4twM7hC
kyavajcEtxPVg2hKF8dbQUB+Er/A5cy3GWmV4vs7SlzIkUi2W1hnBswd2NgMCTTFM+bi4yGzcQaV
lV090t7dByI2xpMbm2mn9FKgqBJIfvpWZUw2GWrBe+RNG+VIt7IJdG1pINTjL/GZ9s9caBEjhvzZ
QysdDxcP6TqyLjQpsE99SLejkViSp1eH52NcYJxILFiqlf7shkWZDDHnRnJPo028hQh4yzqD4lxn
Pgpz41w1utF+bVkszv0egmwSXy6jEvBow7mvt45PWoNus4GTYoWowkjuN6Y28pInaKc//5eFBQb6
KCZYVT1/zrvNatji4LVKqFDvwduMe40DLPgpqWoj9Qh0GJsaAfQSxTOXlP6pk6jt8zyccQNa6Web
iDDdEBr+No7WCpmzgEtwYTZr+HoTiNz6s/OENl93hWrnk+tK3oQYnNQsNIj5BSEk8Vtoi3ffxche
NfkcROzGWjfgn1rsjIyF7BJt8HnhNVJ0V3Uu4ldKA+JRX3GTwxn068fefgnNbFNgY0UyWFcx20ib
mr37Obe1VzqMsTF+0xT8h3NXKM8Rh6IjQkSBK9lg5KmfVm+hDeGXNg9+Mc518BnV1GRqrsJby6jj
5CYtdLZTv6W8QhOXfOVeePY0psdDR3LuUDPj/va/diZu+0aasH0uK/64S36oSdYY/yG28Res6jot
/omyVOh1HIaEZg/J3No+twCi/hg4co22nSIHKzznd4CbvaCznYai8oWF/JSxTWy6vNZVvFVuEgrH
LX9tHHvuy0shosXEKMho9KN/kfpJmldI4yQen8XgqXiA5y8rRPGE63boLKFp6HD57UBz6auuawQO
kW5jyla7gKHhEnabI3hJ4l38SoMFdlCckF8IydNDUViwRfWZAyF27/PyfUL9a5VcVlIpnDy6LiBy
mJRM8pNggpAsZuHsqZPysWFpL+Epljh55vkWR2Mfn7YuF1VUnNdbbiRi8h3I5zW/Zyz4Bfn+ou+7
MZywF9VaGcV7vKnd8HcgfQ5VSPIJcefATFA92I8/F/KrBpYWnzBmm5Jrf7iQd0jSDQz5TJOPAYeL
FTmXBKGj+WK7B4ZohFkil0SVWLH+W0LWm/qgT8qqVRYbRH1Cq7XAUyiXovUC8+QrUIgkQZBEQhRm
3VMO0D+/oHFbpSHSAgtPM3jO3IO9svkgKPBkjCr9qFSPUxz1ZJN2VX7BNMtdAAQD/G1GFcFAaATi
lSbLuspSPTpf2Ec1FwPiVjnXRslIiC8wglHQ6UDPrVEU9aoAS/Z53jUEQ8Dekoon7PjDKEalLDCP
PyOMqPRMYeDDQqxH25M3+/8LupVU19VfXiRanom+V3b+HGB3Sy7pk+p4KojNUzvdKG9SFuHFWcdP
UF/Lzp7wG99vTrtZodFYz8QK8B842PVdTF6EEwrUXwXHAMCX60bQvIZIIee1LnvJkko1bHTXrvtj
T5gx7xs8l7zKAm7JtE5G+3wWkFO5eZG3QSvxcoKILQqY84z70y8gPBqEq1j9IpjWSLklVQhhU/wu
IBi0ej1wukvWcnjVGI/bhpPV4gaBhCGG3UCJZGn65OgLjFCb+V0MMvtpb/vf7UOIdQfO7L/trBxi
A4EXPjr7mF/a7EVc4w+ckn5vtw47v8wlNQL0X6FKh+W6BmSL/D7PEti+OG+5hi8QF7n2Reb76tsN
7vB7VHtbFqQD25fZevRDSyRt1hZbZGXI0zTlH4/begRBM6QCdxm+YtF2XmwBKfklXFBfrO76WKwe
4KsFXGR4cUzfQxSbq2XIuXPsO/ej3g47k3ggFaiLA+sQYET2BupsHEww3H2SaO+j58fpClTMMKyx
i3udzbf8hDBBbDXTNj0Q5nXmVlgYOJW9Cyok5QIObeuwKOsBkUp/XtLNA2FtUMk35swpMOrseSq5
uIAQ6vZv9hB5a5r5/XE7Mse/MelqyeWAO8xNZF3YUdLLtLLvjsDIb5kw9xZQw5QSebxUcS+Ve8Oc
jdDl/J37PJGSZBT+JcAUsuNWio4AtXelmvL8JVAv9Ygz4xh/BOJWqid4OzAoSCuc9XkDGxCTRJua
NmKMlJbsA2ii0F0eADFHgJHT7XVhG2/LY/1FVk6AlipfVVZU68ObA+CYb6IXPiD9+7k8fdRDvShZ
bWtXPkve4x+TKsQv5MYMMHHabCjXWpV7tqUVcoJIm2DBwUtn9qEsii8ddexsmXp4zBgUZR++OYLJ
psKfS7wel1UCF5dyRVH2hYJtL2v3KR6B46AV9W8DoxH/Ki+2sdCdSECYRvHdOuWgBM2GGrsKZCY7
XqG9ElF6iqEpG0df7CTAR7PMUbmTqpAhyBczcji37SGYHSIDsJ1EXW9SG32B9wCnn9/vCSrCyZ3v
rV8YJbSc+RhCO+sc4qKdw2osh3tjZMaGo/DyK++XZ2TYZvOKA6psF1x1O4ygEO5E7Il27WcMqT7g
THiE/t5UW2aEpEwn6Yt6+idK+zENmjRWvOKL1Y8cpJj/wJjs1S2e3J6F4TmtZHJLK0/rwUr8Eq9r
tzEAliW02iMoSiuu63ryJ7kmL3YkA1scsXJzwqnpyKJfuOzdP5o2yYzirKd6/RC368g8pSjDHXgM
MVj9kiFNq6SExiSBL9uAS8il8IHkfeHTmYGoWE05bobn7Q1u9VY1o8vurlpHVOnNqTpYzT1K8sFn
gPY9v0mZHIXHpP0VYKLF2jU1udvZlwypjL+/07CSqyqVyCzo+6Bcjptgp9Mrzp8euW/1n+jzR1YC
Awm89mD3CyntJgY/V+3T2AgETk/ELr9T3YqLDcxW7899wrTRE9R0PkhC2jkDeznACq0LbwH4VYt2
l63kQ5aTIAYV//UfG6LgyB62LzmWWvKruMCJsqQ0jbwU+p5nFSNgmZjFqC105vQM8bkoliplivsx
CFrUYX8YeZl1dHcmYOE88p7WCIF5aNdO4jgykMotdBzxjzRLGkLeGKAWaoJ+9S82xbS0e4sDdEdJ
Os94Ur8RwTj8JFiYGdmRHyK0mpObbTvnji5GRcBRRhmerIQcIorJHPBqFaDLOxjbdRZtTn6EQ5tc
UsGiyaAutTSHopZKt0euAat9SQ7kJFzK7uyPmR8utph/mwdzsseOCZZ1c6cFhvI21ypfNSonwB4M
4cnWa5jwZmsWA5i98FjOwbiYMtROmFAs+q1m20n9BKP6l4ZuC1UwL8B9mQjBW+8D5uZqhnpPHWSJ
TQXV/jJoYuBf995sXwJvYPCLzDWEnhFOIzZygQBAZMG5pr85RA4LjAYz1S8RD1OOa6eJ7kAzuvD5
cuFaOc1/3AdwhhmdK5TdJkyyf1kDw6R7f0fB3WWooDBvYYV5mJypQYRcd4oV81nc0nO2v7YuaH0e
scBvtDeF+MjOJQ9rEK+6noHJuHjV1P+WchZ7t4NdS3i76ePhCylJyWvCMmRv8mkQN/udRs2OgG+N
1kOP8VAp5vz9Y8+78UoWdHUUMZT32kK815JKaARdFYg/faZ10iBaWZgYA+WE9pgvwbRW8kICfu9m
jqqUuqRc0UYN61cWVNXTdZrYfJHQ8d0Yw5SgqyrQNo6jKntVojCUZSsl2KR0zcpraF6LSujf55FX
SGzX7SzH9Mhr2SqZRn7rOZy56Wo+zZMFrBjthEwQSID4FKrCEXyCb/UfVqvEesHPcYJqdKJEQSBG
lip8093pAuhnmC1AMTECGogZMu3zrdnUbGQ7z3HKRSUeDH9JyfaOgQUSXLj4AJ0CvM06fd/PE/XP
5kZ52suS6995KL/p5GqmcKelI8PevA0ZxsRhO0g9BMmZf2EYZu/ubYLjUYZ1uqj+4I8iboOJDmB2
xaol07guhjTxn/qJP+v/77PSls8bF/O9CAC4GsdG+fpAITq5lUeOljDpGFlDhq16/aepD6xSDU4f
/FMhRyL25B71OrX1x1314TdyABf9+HSTB3nwrYc5reH95euTXpWTMHfU/eSbR3piRrGWGHkq0F5S
38OE9rBlKUf2becUFuv9YLeE+aA16I+otxp0Dzpk9L/u3lTsqUYQg54n1RFEw6B2eEjlL9AGaoKQ
7Lhs5MqlYkgmQoExmT+hEI3uoQ6pKiatgr8GMD5V0x3ldv1SQzgdNAX95GBkAceYAtAamIOkWsac
OimHSq+i4z6pul/dB2t+daISNJhk6fbHxEVdRkaOBWtkJ2V+FvdGFLjdKHArQXLVDmKTz7kVDpTp
QrAoYBKSVmgV15cIHsNX/vsGHcSQc+8dHOsAhCm2RSc4XNXCDYKHR5Zzau4CfFR5m5/YEGanplDv
LVRl89LFpxl4smxyEZr0KktMPbQn1h7i1FGzjySXhXJeCL9//gReNuWkDxa/h8XkyUqTEwkXl5rS
TTgTg3mJ12YW7gCQgNcRsmWXxEHtJxpbuD+l23TyxsVL06z8fgkzEnXpS1DBpKEsGr4QRHjK8btA
rbfbJnIslj1t21vv/ulRhPzi8v5EP5k2QRkZCndJufFLVFoQHqJY8wmRXyEXQcfNqjx1EL8l09yl
hbAm1rFTTvpDOKIR8MH4HaNBginF2LDn+kAz5bVbQDBE15RfTu6CUgqJZJdbCcaJN1pwT3vEVKUx
YZVn4SBnSczsPvpcoFVn1XPtKGzLBTdWiJeK12ojzu4ycrjwaKw/Ht5DMaH74HBIYpQSNYEiNZW2
slWy/9CZrhsMIeh9L7cE1X5c+I0TpLkXrynM78n4NA6rRHTU98YEN7/8jYRzvFteaiP65owfrM28
qPhUHqPpDejiY1F7Ac7yInqjPuqIkDZd1wnuUHqMTs3HzJehsGrgz+A8qTbd/4y0S5sV4rDsDeOL
6ovJ0W5NpOCucLt1IG/1ZtbbpdNZZtwQFTviAqVSyK8JFdCDDZL7LgnnyioI1R/EYXdvG2hLn5dg
dhFqx3OZJKgv9l6LfypMibvt3x7fxDAenyhGFya5vacKkR0QD70UP99Y3AKxbIzEBewctwBY87r1
gLzYCqBgR2WX9KxsR5aXi3u4bSUPP0N9S6xXfCNZ9vNlEd69L6HWcqcUVYPeRPW3tMdd7Alz1GwP
Rm5JasVkRkk4e0oX8mtarrOk5/CRENmzIRcRE2ZQswrYCuqwo0nIQbY+BmQhybwtZiP3S32Nz/Qq
30NGZpUcKdfN1f69d9SLNIksX6sj9ckeDqrobC6btbMjh82y7BCvKs9cEUEvL4melzao0e1Z88Q9
JJO/fwBzwj7NWdDlKpm+FKKeZ3QbJZ2mfEYVxE8DohIiFD2JuoUDijwgyFNpGm4+9VM48NLIaPlo
4rOaVHzjjzTOR8LipO+uPWY+1C+yjEd6tnolEox02SfN+5PBJkDTsh9X4HoaK2qqrFpyb1JZhEv6
Hf6HhJMZOuqnuyqv0fIR3FTbnG9EzB+cui/A0mSSs0vXeXWh6HSVspj+vvHrinnakHfGl5I++H+/
ghC+3xTg3mbNDdq+3wiCXaD91J9RBl8NZ2vaCmiqjOuNjHpYXSj/vzWM5Zt3gWcfFl678LMPDoBR
4cBLFb1OhkAod4NyZuJ5DC1Xu1ZoW9IInyll6md8sK64aKDfukmzQnIJCDNIteYv59x6+vBGCkyi
QlPPraO/9Qjb+A0RwK5Fy2mWvzkH+WhxytF6Dwq6/AVHq9PpsAk9VM9757ZNqYGBps6pFfARfPXW
titlUbsxxpkXP9VYyUx0StHoXHIenipzbxaW96bmoHMi3/IedPGVXzud1zSx3Vwp3opnMREWKoAK
Ry5wQvQFKvD+U6hU/PaNPfQjzbeLW4sWg2kOjBrsK13R02hWEAE4e1kU3/y/hJfC2hxZNBnekWDA
gZvGyd8Ic3vpxbkk7f3xUBbZSgdbCgD8wxRctI+XkUcDKjijjyF0sn0ydW6ua6zzYVOyGeZBhWZQ
/B/L2HWEZ+Vm1BKnMx3qy7G2VNe8kO/SlinvgvNLzMYS/ttu4V58jI15DYhrCjOrqXbke08hlzd9
n/CGxuqaniQbl+88K1pU6vmELQTQFlDL7iZMEXPufYKnwUiU4AqTG/mjBS8lkCU/If4CESBz8IVP
8G42z+nD6j5LRy9WwxVvJm5nqRzWXRVD1oQ6QnJSFGKp25DWLasSYcHTgi8j9rkHYOJQHA4TxLbZ
gBN3vrfAc8kZsr3oKJv8VFDGggC7An49Rd5xSYkZDxeAlJ3G2Y9QH4HK552Nwpw0UzMHuLnYtdea
t0qFkDsP+MK9wm8+zmE0dLaKd/CamvHMULbVrJ8VTKcrQbdXsF8YFwXPmXw3zJDXcUdVPDqA8eEg
4BG0tZ3QeVxCD8F4AQylHooEdp+T6ubRUMcp+UQirAX3JkRZFBo3bwLm8SyeVp2fYM0unvjCwtyh
qbIQJg3TnfnVqA0+CZoVV1A1/4FURQztZd/ufH5OlSGaqofoNpPzNwPGIrtyeT8Gr/qtU/IS6ptt
Pqey1NVRfeUOSQa7i8oBN5I41nUiy1M1CnIl3II7z92Ff27S/7VQJt9Lva62CtgkLAtVMZLKJHsQ
aWZVGi6UEDl2knntQ4sLmhZjfanpgmmgAqCzwSc+kOHMdr15fRqLhSoIsKHBPaHcceX5EO3boJbt
tqPHX0Ej3DjLNhiK4VpXjzMMDjqnbnMMw4LOor7JT+g01KWcP/DqCjlduo2v6KBBY79+QeB7Tz1h
t1qmN4Rc1+porL21v/veQAHbTJ+HBp54sXiruU/4EBmQTuk/wmtjUqvWaVaqEUIMiVrfGRsWfrz0
5j/8FhFRLyyRBh5xjVG0rwYbdtInKmJLGv4znhOJIYTEj2pGRWgr5EzZd5KYqSQ5kl4CZIcMjLWw
WAitsCXnF5xiZB1MPAmBVa+cDE+qE7HnzQPOV4Qrbn3+SbzOIuRykrBcnZ1D2GAum6WGF2/UAuzP
p6ylxzATCV2/lVpBmGxtQiYdqvOoIJXlKqzVqLXU9GQjoTDGx0TzYJ+VHZ4t6xTy4Jpb3hBy9ghN
SV02ysn7uvZNfZjtua45mYbPlSvfBVPZhe4n5sHuMgk9q+lVoK169RkYTrHLUC4FbakDEywVBjtS
rAL8bfFC60wUU1gGSuRy4v2/cxjJLmNZnSaoNteaWRj8cgbJ/Cby8qK3veIfK1VdxjKDxHZlBabP
052TZNHdPR9TEXFvFlMPk14hZOpjCBQ0urHOWIwaZh4U/jloEb6VGPZ8T+vyTnvlBRQX2JCy2IdM
2RPlsPpwP6mXEvsVE486n1oaxHa0tDO/24P/Q1H7JBIIeJUkUVFP3Sc2iM+igcttlP1EHQrawr3O
PDfyjw8gi+/7NSBO67CMiDrzF3HIN4NpVkyxxCLxabRmcDJlLQX4rij7nXuzhhizj/zZmojubmIi
kMrQEQ9uUkXHv0gyM65uWgL2pSGVXRHggCn/iM0hrb2WGZ2fj1k1EsA9cPnj7mDW5nOtCIOcthUj
UWxRbV84egojG/65ratit2Q0DFP6wjHyUU5dqclKAWKh+3JUFkrwkvWZgiXN10tnWDzbyetVzF6g
vRL52qBl8YTaHpDK0WGDwE2x68N7MdUF53uWU14+w4pag3LNQ91siSObHMcLjx331vfNpAMJzg78
UznriKy4Drz+eOirAc8o/Bd9Gp+xfHX4zj65EgGaIfLeCuu+8yFpdBa0TX1gPH8PYGexBG7R4GWk
CfYSEaMZJBI81WnAY0Qv5/8r3E1T2b4Y4UaywFMTlDp0yLl6TeauohF+fDroVIM0fBSsz4Vui2vi
p0eKNdwxV7m7XAhxou9cTEK8Tokt2+RNra4RJF7gG4ycuZbd/j9yrmzrwoRg/aDiSC3eI/mgJ9PX
IConoCT8nEc2beDr10Ctg+Nn/2LjdHW4NG8GGsgcuC0sLHp1jyiyUhrXOrXCueO7KGwDttOqpZBn
iZ3DaWFc/gdFFDgzs1sZfiQzMI1tMqh8V1z7AocJPUIn+lGMz3dPHA5g8h5TIJUVtdq9ZUgkRXQD
cVvu5v082IDemuLU+xhCe7O9UVMfAEEESRthwrxgb6RSI6JnzXFGnJtLiJUyBavBpJwOqLrI8ZxZ
Fxl4AhVGFL/HZ8lUW5vgCJzSHezOWE6P0qsex/1bXY6M1ll0pwWCIYwoP7K/NXXmjIvoHAjTTBIi
pw+AsU8UJ3g3L0i3WZV0Gm09LyT9OW8GAGKZQWM+sIkGRCA/UNGfyv62YPrSOuaP7jTIdxHepwmy
NgVvlw5NtcLbmGUaiWApX5Y6N9TvZRk6EVJGDGThN9BIalMeo2CizVwtcSmGYKEviikEb7tpLPNI
2LJu5X3c8CBphr5U48i5f/ygJITTyJL0ybJciYJQ4l4zP9hlsRgg5m1+0XuzTHoTKjflPLZbKxmw
4SxAbmwcH08PeHvi0ZlsBr5bfeyLj8MPFed8HcEyUgiBxppbKyI3EmKwka+duNhKOofPOgj9TJ7O
HkOg9e/76aktM2tnVNaEvHfG27xgbvhOrtAFbKQYku7S7G0KnAM3lP6gFHwCryz7/O15eC9xxHz2
YBXIm5q5kRePMvkI5j3RmBmoq7PRPY0p12qi0RIvmUX/pfJpxApG0Ga8J2fKiqEfIyk1V0O3ABQz
EkNEUhwKOQjTJFrTbaHdGg0DyQP2bU8Q8mBOq5CVv93jPCkSqgKq/fKcbF4n3G2wZZ0Z/PUXBkJL
tQ6adK9DisJ11/P3FGc72iYwgvwrNVTdezfh8xeID4iZTObMEePsjT4eMHQ41XFerrbxTi9gmC8q
Y0NLqu//wg9awH+brjyu0/66/2e68bmkaFIEOhjpmNv8Zv8XIM+NadjYpciNC03n4Od00c41cTzD
8GTbQQGNES8i66OLSsqa0gcJ5Fi1grXhPGmMaxTjcBE2UfP9hQTbdvs3Vfu+sgi95jbesEKPDy9T
ZMFtppvYos4ZqbQ3dBpdnZrs2hkKgigNfMI5YC/8USUp7vfIqgfMOYlK6FPkEcgFzS9imykG+8sh
Og609l63LF4D5Rl0l5Z4cS8vZLEul9FJ/FZOkIKqkwa3ZWKX00Lb0scw2aSzpcjqZvYtrz4SxUkG
vYwTfUUFy5sZ9YTARSLaQJuLK7dkgXz/siBmltfUsDw9wkDTrMOqe38rEsK1UVpGyXkngTUhRHle
7dqfRTJAsaKOqvg0uS5qOmW/lb2ALiynJSFMxToENorKZyr+VYIDY7VQQ7EXmf+PlhMOkZxdE8fm
JrWE8MNUu+rLHxhLHOSynEQ9fiG7WJQOqYV7OSV62xQtUpi5wUMZgn4IoAukoUZjB33MI8wI1fBL
wVLMVRe9lc+EkN+gp5QUKGi4zonzDbhKcgBJX1JScyzGClrfmKM0L6LqmKaSVxmXtDHRYgJW+Agh
i0/qxpaE0fIqilcKPSQ4KxvDZk8FHm4Wj4XGkSI5/TgLo13WziidGbuT4gmg4DhlCdCddUmOSQTp
6CPbtmaUggsAGKmxTWbV+NhORQYQshJYEOT25giBmEIOnxZTVh/tmMUINEOBd1Wn1nLBD7RPUCS2
uuL3lsPgG12B3Odvf9iaZzeGJ5vOJ3LGge7tjZkxpiqjpy8jkouxQKNT+3B6lxoiwFN2SeIx5LTP
Z/F7WUCtV5/xm4v1I+AyikCI0MINyK7kqLeaRFXnWH2Bv4ZSBWC8SXTn5evfCeBQBF9m5qbbHM8/
plQJZ1hx+72bQ0jrrQlg9g+ZvXOHfWhuuMjV5E5yGziWj1hAv4bIbJGkU3E+oyQ0tSmAG+/obNPP
qmEo2v6zNQPob+PvNmWRVU5EYMeM+8+lfzw/Yp8DPII4idohy8/M4FJ5iKB1V4UQaRDs++8YPs0W
zN9gtrBu9U8GXq3wOGqBV9y2I839VD4GLEtVA3Z8Cu2uLDVzng1PVAAlhzR0LpHfGRc6X2EFaKH2
JQIhAX1pa3Wardw9WQ9sUbqU55AwAVtgQeajZ65epFCN5GiKPe/lwsTIPRLktL+5oWQRbjaSE+Ne
gnLjM0ijoE1spJxmlSOVWsHKSyo3hQJ291KvZCLYgt9ZQx8yzZiG9LBgzZbfFVtk/0wDP3St1iL4
K10sp4AVwL/64jixeEEpRAq6AyFupvXSqjoi+aQiOZtQAtUqbf1QC75S468uFcQn61j8Tt6eDq4l
+T8cfG20M6cOuTzQ0DvNBlzujaNkDo32jse7XfeIzY7cR0TV1m1BF+bZWhGOIEDibtUhFTMSo/sS
jTRLRXQw1PuWnkeme6B402vwh0Ot/dpCyQsHW/wmsqGBfOh5ePnLEUfPAaUvP41W1SVK7C1Kqf2U
9xz+JEbvzww1hzHeU+ROno/9VwjwZdaKYHa8WjSihiShh5Q/nGE1u2oYR4MOeMe287sCiCT0fdbF
VkN1MfRecmCUxeLOyGObMoitTfWTLNRFq7Hfp/iREbYZHDQTlOBemhKGARYcgjcymzQrYMHhDSKf
nmXGFeF7lw7AlSarLCc5jf5nkNB5dIM/qvz0kByfYjca0WLo65Av/lPP1boZaBCyIHN87f6T+O8h
w52GW9ofvNGsML4Z6GzN6X+wwG5xQ56OFTPOiz0JyUqUkfKX4JWijZYhwj2xfUWzh6BLt3prEqBp
ml6r6AcltCsZn/pOvXrRPUXsTKY0aIu8Mqiq5vx2Jn2I5J2CWAZGpediakSThIpzLNyIt0MVf+aL
cfWeS6dQBtjd+503e6SxGCayWVqHDYIi++R7KuNMpNJnop34yjb2RVdIbXk3VoPEHaEg5jfMrUm1
7M4X1JWfld5MqN+dJBzo+5QHO1SPMki/aio5EllJLHMT1WTe/MiYJpYfxQUpMQlM3IfK77b/VNXd
CU8bT22P6iZTg2o8jDmCvkraAEqCmjvrvwpa6J1VNFDTulGnIzkr0pnBN6SogiKhg7Hdn75oiqgw
t9TfSPXN00qMxfSOzN0CvFklx2J3EVHuC9CaOoJhdAU1cfaJROmrbWMQJJfQkCp2/q3AoKovqJVW
S6PZUvwYZfSZvb2rnLL80DsWBwPzj1G3B1BbJg0cywFf/XS53SeBr2f372NRfSPB/Oz2ND4GwTlL
lK7Tpsb6UKNsQxI+gNN4Fbi/VlGWGWhk3h0m5kSDx/gWs1uh5ltDi6EwsV8M7AsHOHdZEMwkNZ6F
w9B+FxOOoIqOhIE0nA/0ZOLbDoIAtdjBfl4O5c3qgSmHIYnKBXoM2Z58kWRg1/4mIZtHpz8NI44n
aMRKdyjYV3tfoBS3L9YicHD+FT0mIc0dJXNdqTikGjIt+f+Gl5l9339fSzJ2cr9iDSvWkc46dm4M
DpcGgQFO+4zf0rj70TQJIbn3n/kVznfLEC8EbA8LSpBi/eavEh6quDRPoJdoUya7qyblcLXpjnUz
nyuDA68MgyFGqLw4b589NGDIYeOLWW75fcFN1MkAiV+UEOtYjKp9Sd3o/TV2prKrg7YBegaGt9sN
eCqCVlQPF2LJ3EbKlshjhyeFeUvBjGQkR7xg6clboKhHs1hql5/WLYuas7Qgxgzj/CZb0/JUPCbf
NFZoWwHeQJhj99u0+N68/Ehn4RrBwaHAZ3wLokJ0BAqmSOMG+0HSiuDixwAZzacKBmbP+74447l5
MrsM2hd7R4q8smcXpe9yS5jfya+MND4962UVRpE7+ekBrgX1RabyqJ5yhQWXjI15+35NoLmsRv37
ZF8e0n+qpgtNSfldpK4fJM91INHMewc2QQhrUTE8167LBKgDqzlnlsRkf0/SBR4pwN6RyXkeaHCH
/FnV8Z5/d1/e01BsoItX3ylnUl+kT//2eBl/dpXiVGA6gAbW8NzUi+UajIz1q6svk61GUKQqiME1
Ngbp7zuDXkVKyT4aS6WNGRANVOvIiB0SwtnJH/Bbhk5yGLcc1rwa51f7JcVUFPZoc2mLW9DVU2AN
7VzjZXga2a0oubP9XWrPf47dSh1JD6b6z1WNzdQ2nRf5UV+lKycne7DMuf9J3R55SpKS9FWLSot/
eQqA5PjM5Ai3NDEgqUJfD/iNidIq04tT8vrsvbJmcrMzuBWrrxlF7y3qHTkz1XK0/i1p/bPXhZvj
olN0a++LfLcWuli+1SwYkF0JMVE1b1mqpK2ClW637t8bjkeUSc8K1IlwlamaraFM1uESBKeQ8r1K
TCaOT6ezYd6p8bzZfAwZm9P/D8YiV2sCb5LB5HOLy7a3jIhJsLgI7v6CAwiUGf+D5PuYliSnOyt/
f933WSr2HF/28FV7bkh+ZDy6sc8KnasBHkA+MKqSG4599R6cy5MuivuHGnb/2pmkPkmHXPXWud+s
PExf255SmwlOPMR94nxRtzwCHInqJ/FH7YpWCzjKWB8dB+1JjHp0MaXCwT9zEcz1VqswsaW2ZWMW
5R2zB03pVquqTtFAiDNHTJsn2x2TNLn4XGqqmtLxAR4x9l/uP6WOor6qoiuyWjursNtL4B3EPmiN
oNLnkbgfVDvRSk+AoxjVj8C6VtnnIvWN7tSS11sFau346DIeOyQruQXMm1fi5Wg3FtZ6DbC5pyW1
6udH1ZUa+qDsVPpXSMv0QJYrGsivcA5aI36XneiGTf7mvDzIGCEe31mZ+OzrMjQZ+tICb2aXjMRp
jGU62rvyknf4D/Gq4rWE1f4TiqDF3MNpz+Z3y5Lnv7LQ5W1ZeID+G7CKmekCJMx8Jo/0VZHVrS3W
hKJlFnCgIVo2iNAA5WUJWSrlOYLZ+CVxdPVRV0lX+Az5HYE8P2V7cMx1k8Ts7PxHmMqsdT5EX4BY
pnJj480BiuplIhaWu7887Yz4ECCzcD/oQJotqf3x6wQ/8indyrkuewSSYGdBTtTwSQoXCCoTX+JA
ATGtJOH1kJcYTeNTOiurtAQoJWZ5yCOtZtNCrmEYNkrBVizCTLw/Gv0PZQMD1w7ItYa5iccS0Tua
wAETv/akUDFr136noVELmLKuOtn7LAImYJ8wemW2j07A3je7JeDMCu2dzxbKX1BI6tPHULKO672D
X3MmNSCZ8iLqTbxMBLT1KYynu/dX97IhDRHdQbajeVYbiZmlluLfjW6QsL+1j9WJbGbEqWyRaaoV
F9cb4CmobK4eKqyKeUoRclFwsoS78J1cpKm2gDpnEpJP6JX3JELW9eeYjEpUKgKUSg4dJa2Mt8Rm
rseu/d1kueLNQX8l/h8VVJiMhcd8aUOX3cp4TsrbNGJNas3Ht+QbDMHC9zBPq1e3ZuNTLTR1jJSC
JMOzDHU1sDAgs0aHZU1oIGmm2032fyK4+98p91UhUO0Oo1ZW4dgqfyY5WXTaOfwR/GP3iyRdf/FF
rFeje9/cnuSVmgq5990ebKfSJnTWBLBHrlicPqJlCsT4hZEM5ccsRpYon3u+0ZKKqyB0FxELUtwA
4bHz294R/esx/ePw8ynvgV/3kUp5Y/zqq7w2+5lYjMDQFniwwkJsea27eljk7mqUwEPbuRqzk99y
kcH221zCf5IM+YMKqW8HwiaKmbuQbKwDHRo+9kSsKQ5YdF/dYA5aBLn7VXC0rxcbH3jCGzKbnNgb
ulSN0rvNCINPp1ovKNM4yGv7tZzahY5bwpVS1jq7UEg4eaEvwIiaMRkpPDaIzmUpnU/ycIHGx8i/
noY8V38llfdC0mlV+3PjMaF4BuastYWU7gPH48C5NrmW7G0WSyvA5POwNUTDl87Iqv3Zzroyi626
zJZIMZ8jAlnVwfF16ikJ+ZtAFLvTdxIYo3V1w9K0pyO54TBFyu/kA2JXPKWdqG0MT+5ILRTSI24p
AC+5F0E9xo0GdAXiUEhap1ISt72/tM7dykyD5OxEvVaDeuZ3KJQNe5HacSjXHGQis9NeAYMvDKro
+U8dvRvYru1P+WtuxUCjPUPeWpUALKnuIW3OgwXAE1oKfQUThV3enoh3OZ2BxpitMW3A8Dmbpi/0
fBxZ08ccaOpRgEPfoouqZjLWqmZ1y949RdEcSZDG0BG76+MBhePmTfJDtzJXNlsrdJe4FDoMaBXo
mjjca8IaQFj4Tw4FHoBA7emAVbhnW131j3Fqe/qJZ3nHavJVcutqOmUyIgvyQovgtfIG+Rxxk75V
I8S7P6mJLN/aCHvaVQc1cPKL1NgRfR1fZuz+FMBvkmCdHV0HF/p2wQ9d0npUtOZkAgImN9Hz+NT/
CkjwojSPftNOxHzmPMRuTTi/GCA7hWbj4gxZWkY1vpi2kn7DCskm4sX563xMwEJa2uqrxd8FBZN5
JJYX7eBFaAryqjUMJzhC7z6NzUIf7/YHfOi7pp21h3gZ2v8jgZaeDp9h1Rdg/91qXzU/clG5a2Tg
GaWr96/QLy4S9Zi72yl9mqfqkjhUObtYNZVy/vf/YJrdUHtE5A/tITmBPXJM5eeP4YvLVbzjay1B
KxZmR81sNHWPMpVIuxLDxZh3T6lKB1GlixBvzGKlb6vLLvJd0kaB6aLd5GVVrQfDo3u0hSpRugky
nB0ZZ4Feem1/r0FBvn3DfXda0Qs74QrAeJbuQ7Khu+EdQbJyY0u1I898V9X5TjTZPAjY1JE2X2VB
atMjc+Sntz8nEcdjg4nXvZ8uA7teZiHbU14bcONka6zhfKj1Qytz4G6W2fS38OzBo9I72mG1+91n
Gxv831qhDQ8ZQ+qUO+6O6k0Yu17sI8N2lVO0/RIRNZxOgnsfPhYtRU1aKl+mi4r8+ljzuyWmitVB
b1LdYNponuEaH4QjGSVKwtBrVGMh+erElsCEgm/zD/KotXmlmhzV9gbSI83ITpLMQJBfOw4YJV1d
lJVrGdHIT9H+dPZM2ZlKMyW+k5cEfJ1GXv2wGVciDNKmjMmZ8zxwmB0kaIhFMmcratF4SzHajMl0
4SY0oLgn/M7jSpxE//mlHhVVb/yZqnnByRz/H0XhDYFscuPyy5seE7rhlK5u++xVzcnzdEcx4ZkM
gon23Hka8m42e1RlAJZVQ4zs+TQrW5yVo9io1qpEWqxIStxZYKh45fcJb5uekbxsqhf3xkR+7o9m
gitpjQcU/N8QnBhGzIkZx4rJ5nQ/rz/dIetMccPGIZEMe1kpZg4uqNh1vgbCG7ZnmH357faYLZBi
eT/KUWfQJ9iHVxI3waVxEuKV3imROCP0mrLYOUueTAXJpqrlALMMn7HHlkYJPviDQO/65JmwuHeA
40fJi0ECXWG670dN3nhLry78bBzoGJzucuawehtydgUmKlrBOHR4F8plvYfFmUYgAVXdOwJ7ZPrK
uAbCTHjBVA4p0J32SzgVpmNYabcosOSNVJhaHr24KJPe4vhlNTASo+BP7SHyVVNx7a39/Nr7BX3A
9CRdPJNYSvkrxJY7FDk3qqxp3zxUzvCFnjTmemnxog7nHYVBcym4oLw41rRH6U68v4ue0xH5r1yc
r3qtHsX/mhVGPGn3eV3x0G9F/UdEMz3FJzTEpbliIkjdNaYvkxlocprMtu7GT8nf2EXnANtbj3cD
dcCPlqDqq9LWixlVm6S3Lx61kKqqizP7ivX2IVwJSQOUWvhEP9YHVhvJvG7MdbjfcdD2YPrvdVn5
XfjoieNyyTQTXiy9CZS4vPQRDNi3WZjplO0j4huSSMGlWgCKEq4fT4xykyZMLsmAG7g1oi4DGaMk
yOjw9cxNxLTC6j+z5dyO/I0sjgCpmpl13ONrjQX9Td03U4/MY2LZziidMR/31N5tM+FfvjmpD06F
eWaKMkTn8+D2G6xt3ugFI91IhQj4BF/wx8MbdJ2bi6++ZxpplCOCoj0ICUs/pRdVcqWFeXXvjB5K
W1TZJ7UXz/GdCYTvzhV8yXmhwIjiMHICLJRTOpRbPHpPAixi5sYeKf9hxKNSTq80Wfpcf6xP+muk
oO7PXwa+tNkAMKAAUjiiaJEUIWDGQ2y8cgUuuWY3zWAvtoFIWC1gcCGZ4xnVbEzrYyBkrjZllLRF
TvV24AVY7u8S+q+TkSbG2NVqKgpgeUqoDWuYbwYPZ76qmnvqQUS4RtYCISRU6BKdyFymNF01Pik+
KH1A542YCA0FnF5e71JNuAKM+5a7SefmuLtBEB7RT46Rc1WtgrpKaHTldJkABOBl3J2EQoGW87nK
x3TFPcMLcJhLGkwmEKMNoCMuoaZ6ip/RstPZPLBfH/g27NDAjU6tWfRjA6MoVeKYPywIHCqwxJgl
Rf7yl3qrwvH4RBeyxb3stv+nyHNLpCQvGKfVJDXupZIaP8fvTmod6mpL5yPVu6vmx42O5/ICn5N9
9Db/Uc+b0Ii02Ju6Lza/whkQmIE6q+CBQ6P6FwnZXBRZ8z2eCs2q61LfJfqKa07sEN9A7N0gqtQw
HaY7I+I6I3sKAxkfms5jBWmE74YkZbsTDKXLppXqjdsrAwVcrZgPJpIBBwzxpL2r6/zMirFwLTAF
AExQO1B1t4mQpM8b7mF2dOzXqupo5itz9i98QC2lnlcLzyJ3fSVW2ImqCkkvwayR23o8PdA8zedM
JqXR02CMBf/8/BU+FHh+IdSsP3o3Uiks4cZhX7xYxQ4MJ5pvGoovhPJmzmlCSiUKUoTIwouuth42
Z1NBUi7xaYXlk491arkGivwz1AAbcG5vNN14VseIfFQxJFS5D25/O1oPvT+ldGiQDuZXWfJIbdll
n7KTggaBOuIjQ7116dbIDwmgSXnzZHqeaD9j1oiJqtBEKNm3h/LCiLd5vg5hjLsW15sPCkOKHGmo
DjSyhzdNXD60zCWQ0Kr1TNL5Q9fC/1j9U9JO8FTfPLD6/bzkaO2evmO1rlSLCQ8axwH94rUPRYVr
ZCQBvtQyHr0cJIggdafEc0kw3wThO9XGFPCOTlG875QrnSLeklrtL73quEqSk4YJf2AYX6tEASG2
sGqmM6XX7SC4Q+/QwCH/ZZdOCfA0ws/ODy0m4fAMhgxkvnStWBxlxeCcWz8c5xAlzSyH80I9dHXH
cAKp/6Z29uWmMcnbC3VYszmge59OZVV7TgmIH39BIXca9TriAu4gpDWy4p/Ql0Ct+gC+JKU3Pzf1
sfHiPyj/dH3WoFblAhkHOIG8OKgPje/gjxLHMXNhWOxSYkab2A8/2ksRohlfzsKNUqrU3vzRmp2O
hUEOO3I0i15gh3+0tpAdutr/eY+AdL6IVMIEFMfPnVoSX2fE988+IJRSzFH7gDzJhn410GcFUtgJ
PEz6bYslFuxC0S+ktDVwsLe/z0X8jo7Fwx10ynzWtdVgKZZl2EGiTupeFR/0JC2i7u5GvLr08UVW
ghToPnsX8sJZPH2AydXu4fg8quPOfMTPPDkTK/8utXBEuSesJXr+D5bdT6ON8ROzgm6mtruROZ42
64z1yTQAlNBWMKVd74fmlTv7YHcCiiJIy2/prOfRFGafK4ewMDM55J3fKlP9n00tCPWKXDxgIZkm
dzRwIYmkABoEoyhfGj4kdnlmTGqTBcWfOquvajsC82b7riGME9IfEZMFxDbBNUWHzecMbe4g3ReC
vTK/+rYqBie1itSSNFKK5IymTTGSNorHM/5PH49/UjP4uXR7/2VA7R/iXfDHddqID3fAkH12G/Xa
D80CGtBlOFwrJKXytRWQ5pK/2oz43yrdEx9gd6/4b9VLmWzvziEf+CbyeoseB+IvMDH5v43CnsxT
EhzLhF62xA7JUgsHJZCIGvdUjBkYMiTrD5tZeyKwmToaGYoORXCVFaFPz/hJGbfo0lbGqtvnZfFo
HQzwJXqm+e/GwlGZ4d4Xl7O92OHC4f6xMlvrgJHxgDO/KeOO0gTrLcT2UldSFmOZOxw8c+57SK0F
7uGgzoBNfv59spZ5tXdugac+p6acm2UcsDaXCqbyjaLmPSa/8uDR+MGC0mqvfhoSzw5t5MmCNLDY
DR0+fgwhuEUkhU0u7Qs9tTeS00cqEdOqHXq5Ujej8AjiBYID/GvNq8mK87yLfcdBP6MrYUeaE03X
Y/TOLFNKbyU1ejaPl2PGjYGFXADEy3NQmwOyuDILTKcMc4Cjd83EsQ/Q8uDGkdvgXbd89HvQ6IE2
hkWOtbBezFOS6+vhqJqf4e0d2tF57i9vfnh2919n88dl+u2SqcXGN1A7YAN3Us1C9aCWfhrC4+VI
mt2Ys3xIgGjGCyUpheCP+FldLGTxMwDU3rJOx+iRbEWLRxhkzR+kbRnZwZJ2WnRJaGurHM932rNM
OrqQ2yRaj5Aub7RWTw/AM1uFpjHRsgjk6eeC3jyq5P9RW/vR8/ExLGUY8BlSCgYGL2HoVOwmClPE
uwy8jm+CycWCvCKBJ3zeDeCBA6mkW4iiXHjD5bRimjXx53Lj4WvohOv0qKbAnkPUd6vAS/pyfQ8O
ErtRKthCbLW4tXLwIA6H7pSriX1G6l7asaYROLkkaNCD6NIp2dofl2aUAlCXDTtQuuvUtE+AcLDa
Opf6pCas+zA6x5rqvb935mPumNgrWU1io1RK6ik80J8Tz+SYU8hvheAClouai0vtY1M/siPmAPkp
AbDS5kBmpp1lqow9EWS6BRJiQI/OCQeoSLh/4sJrPLJojecjwmjOUBPo9f5KVEdUMyU9b1oPT+bv
nLj0toixnakfHh4sHuWJ1Dlb5AqOlj3V3i6NXZ4SxXn3Mzo85TwMhriC4DwbpsUsGxUh4BAfSne+
0Z7IpoaefpM2RbxiIhE+nvfS4NWddprDDkhoBuq8HXeLIsk0Il7eKhvExkSxQiMKWVTyu3h1wQi6
noAd2s+dXUthbQVRpdWN8KfqNCr5ze7KOT5A/BLgWPt8Uh1vFPwqNIjC0GyDypUbofr/MG09+gCV
SSIc0hgwAw2NoCHdE14+iKgxLaaIizPbbrN7+nelErWvpWNgvuPUtHWjWAk2GRmklijSGAJi3Zam
wGnMjRcLuuiqePczbBrN1kw2+A2Q3n3KNl22dXk+a3ik2OzDpqTxgrvSe/I8nV4UWTiqTgBw5bIb
JRFjJBqlAHn/P6dVCAT1xFdcIsXxgvjEldcIqDCrDhaxaWf+1cFpAKJfZ2cfxNH19iABeKpnVEsd
AsNlrQgglwMJSZyQtn9F2530ppzOQGC/YFYIcRFBUs5jWMwfzIyYX8VPQfIQPffumucHucTvyada
EVz9M8x+oVR+6lFHIe6VKWx5pxASnXWQww8QJuauNZJoGtaCvHr3UQP4BrpxgYn/E5Ez++6dmn6g
Gnik1gpZRlHUoaThKsP4nzq+93aFrxoebXuej7THHyJxUWRALo9mdIqkU9CgKWGG69PmktKKtRCu
ZzOHyc8Z3bsMFGwt8FdPSOO9M/nDVSKf1fYdlXKeS6YMfYjJj5fRJgSXwhoDalYRE5Zb70xT0P+Y
6nCDpYK1Yyftg1QXU5J70mP77bXRIBTsaCZYmPBU6v0C6DcUhLVXYkkx/zd1L9jyfMxAZ/rqeU81
UK0sXv3y3QYOaGeiroggKk7yTsxSvNL78QjMf59IfCVRzDBU+j8czh1MOcQp3TdXvre55NMsCn+w
oYngjAKbR1VQ9seu0Q8Env7y2VYZifmMlYYNpQCIaGvxQlDtsqOpEiNeH9gOQw/BNC8SgVlYyY9E
KaQSUg25IZOvK2CCulyaBzgmXUznFDjT+Bj48Q+y/LSo5iTBiqdt2MTH6EAEavcD92lBPfitW0YZ
Eyh72JdZs+KIxOgpkC8TkV4ktZhaEw0tz8FaephqAGOx3zpNz3UtOpSqKDgCVzuIpYxYTaTuMXNJ
A3sxKVWLAobIwTFxx7f4pZxgK2aAOK2adjxkcRRf9w9Nr2qcIstop9r1ylsJDqr5b26XhoE6ioyP
Jm6jcfLXotzYXAPrEhO5+Jr041bJ+9hh591KnrnAexm3+dfU29lg8gGbuRT4j3pFV6HpxiQDNfM5
svwXQcOtg+TrEj2zHkXtHOdOeqhibSGIjs3Q4dwxHYvn4VDoPbEWfrVQM3m5K3juyou+ghRbPF/K
J4EqEZrThXoqLQCS+FzxbmKy04qMqrKzfOfdpaKdRmbtszzY1oqVK4QpudvVTeFqqEXWT3OZhNUf
nFfzjyoJ/TwCONLxQxBkx63Y32oBXQMmtOgzldxs1ZG2vgEPwryitOnqFuorq3WQO91qpUT5zyct
uZQNx4QaSf/jpS4P2eJ16/jP3b2nu7MNN5wFPbyBmuIcgEloO1uqPurfe3Uds3z0XNjHZJTTlysc
H8NZbljQ8S0owlXruzX5gUQwkCOzKPhFesooUOoCFrTWHcfeaccpek1Rf9W5VTKFIb7e4eMROxAw
9AFXitFqfqUlZ5FtHMN978etDcBSTpr8GZz5dKImFWqAJc5JwJeWg0B92TxfEt6ro8mftNVWqMLG
MVeXhSBpFNiScCzXUqUoxx2E3pvuWQOYGceMBTqFlzsYTMrULp+G7sVxLsVWBsxTRmci+IDn0TKi
9ILy58hxpVbv4neI7FuS7sNBdJrr5bJBQVizJXVuhqAYzNf9y2ULyW+mW/irfKd8OpejYaQWoZhn
kHsTDBbi1aBhPXA+mjEtGw19CKY2Q54Fx0rcIiv3+2gvUCv9+3Aq5LLln9e4sbq9Jl+QGNb6PRAl
FB0R3kbxqurENFFJUhQQjEeDH4BkaFtxR9ZtMOOjCemt7Eak3aC8XSQB7GahIyvB2XLXiT3uYC77
RWl5TyPn/2rk1tMnSGlb38+8u0SCNoRP32gFRxbVZDnNFga1vS16IjX8YPn21oqgyr+OO7QrxVVa
4f9FJ5MwPfH0aFnFis71aCw1hgSS6V0p3VgtfH6UuVAd4EouHOtZLJHHuSBbdFhgX9fZqZH3dkjb
hcpu55V8A8fojYt84Ysro6lEGDJTlApojQ0X0wma/z9eG/0Ynrhy2SYmQRYeHFrOWz8fNq1wjfas
BR2sgYU5Qy+gmdswcyiNs3dPM/gf02XnQirdq77rNNwM9jTNH+3cT/I+kZAMhb9as14a7i29brJG
gJWtb2DG8ACNvGXCVK9MVe/U3QKrkg4etCBGF53ER1xU6d/vkp0qNRfYbt3J5sf6bWUtBqzNUD+c
sGkIUgzFSA4MANN/WzXtf9gUQkEWaa+wXUneitI4dl0Pj5pYZLeej38kgj6QEu3pnt4ZrSvImjJ8
oEbPHKq6ZQfOlkoTszjYskYq+0/mtg2X4SARE8Fyed3WBwfysM+H1bFXSgwVxABG7isX4iFZz2PV
0YHlFsX8vDC0lqS2xe+uFuy0nDNR2hL/fASJ48CgaDukk+0nTKeqwQLbjDSCcee1cX42eLGPcQgw
pkSsiKkf6I+lE3PIEw9sPg63yu/0uHJ/+fTqPjI9LjI4ztGAZ5lw1VzyiF4IIqJCtpiCvAZ7xP22
ZsMwkHGJHb9pHz6GFT0gKMukb26kO7g0nPx1dANz3/6ByTBfoa3qQwxkl6Ha6eGbK5RLo94dSeMC
qyXBuPEzrWpOg7HubCosvQGnyBf0QPuVNNWWYquJKniPFXJMnXIXJjfKLMf8V6kGAlxQyWtkbHqi
Om7tMIIv9O7Xevwd9XjGIl00VpClCUgEuZE5X2H9kY8FtuRaqp2DhP/5pPg0WOxKnm6413ho+Foy
x2U6bea3TXwwgKR7arfNAAVASu2ctrG6fyKAF1uzo3JHewTo9jl+zmAFupz3EvIN6CPSC8RRM4I/
VF2Lq9/p3cwOr/ZYXhd8+uXohanYdzhvj12se9e1EBp12dpbXKIW51/2qGSfPwoeQtO7Ar8f6kM1
cRpCCx9JIBPqtnz8CT2E5jd3Gh7udHwdXRB6mNT5kes8iSht+LgLR9xbG08jM0uSRGd4vFBnwj4N
jUh5tkqucD+kFPLALPZ5nQurGUsy6WNG+Wgg622E0gms5+dIIyM2bBXNeZmMeVrnfj6cUr9M8acQ
vrShQ+Tw3sgf1Gxn2EMJT0fsdCnQnEe/ZTB5ZyruzWF9ooX5MPhcR19YS7mvviB6Do39m1MERB7L
mNMS/AAKis2xwdt357Mb8Cle6sbfSFKJqN3wr/5mY20HHcLqlRVEqPabO5yu2dfQ/9fNUWSqMxsH
jmntSYh8RVOmkaN3kgOpfRrJr97hhE/DoQV2gCwPcpAD654oo+tqX46lWVv5lme4/bfvqXheToAF
YveXu51sfwWI1qhvdxPzDC9dKKf/PbUCYK1Nd0KLWSegavXJZX6T5PlKjFZU7Ob+Dah3iCOTQ1cp
QF3+eH0I1dJH/tUPu9jGtvRI0Qo9gNSNhjDbVEQf2Q+CfvUhqmSGrDRojabNrCfIN56vvE17wtX8
H1eWhH+aNveGOMgogYX9HgzMCuvc66Fzf+zoJUXQV4p9VnJx1iuH1DnR8VKpV6Yce754dxpHqE09
ED/vatXqjH4Ra7UKEuP8jCnlv/kSAvehl0YbWiHwrePqtJph8Hg07/7qleLse00KpIVt6GVEO9YN
dq5RWr0izu8Ouj7EORmMa8jO5042T7e6phpTVgsgWXtCSDFkUGn8x8Y3nq+XaOEQyNJSqHmlz7Wf
t9CrL2yC133ue9Dh5/uCJeCu73tfrH/VVYTeWxvsvxqCb4dByfIGgXvXpdFqGKKUE+Y/CmK5DOc3
O3/hKfxnEUgkx4ZJYPUJW9TlF0CtSlnTIBBbz0uTzXp6W4dbrZGUrcEY5auChwAXxMCgJ3J6+Gte
+WFlnjyXoTobvdPtwKVPvJE1HOR+q8I5jp6oZ18Y3R2uElTv1HT/E4MnjOO0mQkSswmeace/R13f
MTEaeCQmhlPOd78DJa0TUqb4QCWlZpq7sCGmdyEthZrorD/FAUo7s9NRdYKGNkoLBTNRDVF40A8U
QZq8AozC5L7Nb76xxEK4swB3hAAfB2uzyQrdqZNx6cTpfPl6GGLxpAvtdBfjVW4Z3sZocv7s26Sr
AiBLxYMu97f8B2xd/lvMwJZLAh9sfrL7Ba4b4U9+Ir4YUERR7bRm9DwYfO76fyAGQncNqjAv4cEk
X3vup6bTIX/44p3+4886d4au9pxPr77x4zuIgPFPX2xPBAY7sUmQeqngD53809NXDA6IGlBOoQCZ
7rHAp9UHXLfDG4l6rMYvC6ZIbjrMnO7ryzOxAAIMHDHZhazGPPmy4uP4UyAIs1DxEqa1LAyFeqi9
ufw/lgeq+FMiBNiRhDvp37fqtixiW+yuRGtLlD0xZaMD3hkgNJ6Q3YKRHTZDc+6bW898bYokWzUD
QpX9qeZ1JDAnKXTAtwO5wUVV3gr+CgYNMszLlExvOQHwWqtDUx8le1ZsUZxS7Q18OJH1qNpNg2K+
AFKG4MrvTA7cuOwHBRUzCzgLt3psuQihHE/tLouUb6tvcbX7osomO5Xbf1w+U90VYZxd9SiQKeYW
1hrzaTThri25Ot49TP/QAYMQpNfvmRryuPCm9Yk2PnkqC/G7LHT3AxAJH2UfZ7xQ6cyTHo31hQau
/oXrtVgueqH/0pKo3SB31rq9xnxWTaCO99rErPJyf0AB4nqVDMDgIBHDqkUPm5msj8kQSzloPV54
l6Zj7QaM07Rwr5XghVYpmIFJJ73qW9su5k385lsIARctDseC7OjIuNnHnjmvhe4DP17rDmNPpR+S
Siu/WLiMqCtkeVAZOoo5Z75ZhSvHVDQxEmGzd+yQL3Yq0GqOCu1R613Ydv+0V1EAbpMVrBkJT/T0
fq+Han4eH+oUJ8gcggUNbRrBUzYOJ2q238IWzneiTvc71z4Lh1Oe8li70l9tM09jHVvcIcasJZsF
UiZd5l4pYJtlR43/TRCKpQdjQP2cxvBRjQFFyKbJgdKDqLoO9Tz50Doo//lQIHWm2Q/Jq6Qq4BfG
wtxia5eC5D9kqvQh/RhMHy7cdg5tQVWgzz29ZfsecqrQ6aL1z6KVQdAeZYkPOfqOQWSUUEgHouun
D+OWr5r3Opqe26WfcxIdTL0e3EJX/oa64buMBhQzwpXkb0/HRIVHiEF8t04nJy0jvzOZl9LyXE1w
/T7LTnyf6dzDGQ9rqn7HZSYa3YxXn0O4fFXC3lYX0UadDcbhfEb2JUiYKoVLSAEOdHkKGBRKNG31
VmQLzRbR7u8laF4cQJBRYQPsrPeuU4OBKhN1A9uvuvQI+7cWlKAgEycwfCcAcswGm+5r5QYGmJl3
asuOGuxelbMCVzuG47nxtpRg3Xag2e1ghP8+zlVoT3Y+BHx5Uh5LSvGYGd11OkfRaEqxKOkqRA/y
lBwZkgi2eDr3pOfcEzph/kKshhYsxi5ItGNVd5MYVvRXQnfbsRxlaJkh3Rjv8FJqtWuQbH08jw71
7v8ZiYnZ2FLE/WLqkrs9rAotd8HclbTDJg2cssxPTA+YiTR6633C7jEGtBerN1dkyOMk2JcHlcAU
h/8YBQBw9b+PcpMFu2n3ClttjhaUbD/4tOvQebxJyGR0SLAE2dPFTEeM7hApOinOyeYfEZwnc79v
eQjZqugSGijayGX0JYOEiNksPVEyJv4tWfRMcdnixsW+9hKaGvDnL/pvV5bAyWWvqQyEZC/1trrw
2us7tusRpR7ZsQj5+tPLoRZlXzwUrIhkpE1HKqY4yDz4lxsVoPW5TAVM7eE+dVf3RS5Z5uNgEwO8
5m1qzCAPb6RY9P1ueG80x9bxQ9roS4SzpunkUqJhX6xPc0YXnpDRhOJ+J0jBUKFNcbGw7KsnObqU
xgqI2JW44KNvN0dW0WOWhPwBPQ8uJ6jB/24V9qDcXaZPRBGMAFdcfqmT10rIcWC5mbkMmaQjWhiX
JnwfOSgv097wCzd/doEO6Iv/j834TLFAoeKFrzcHO6VB+9Yo6SVipMUUMSO9UpHSxBXwJwejfh1/
muUYj9y1nHxJ84yLlmxkwgdSp8RG/qfDS7139GW3zCt0BnllLsU160y+q8T3JoXH8awjd5pYaE61
0nT6hCoI43Si2MUOMVQ4aei2I9Y58inqDlXQ5O0Dh0bgnnkmpCwiPNL+QP0qG7hk1UQLGYFngzWC
XBvOCXW44jb5JvDTWw9IeW7VikJE3sYMlPzFvOCDfWpnTxpIHAi0ibVWMbHcddFSMVXe1kkT1I8l
nMYURv4VaFYmmPliz+Hl2Sf2dByHtUeQmXMH0989Qw8EZb6+tzfoB+VwHAfqWzF8Utk76XUznLdp
GRIq3hApc+w/11YowtAzmE5EJBXVhHhWlqG+C2l3HzN+xo5JhPjEpPz7eqjBAMptJAcm9StP0JmY
71ANGgMUy0bQVTnQUHY7onOD0Kd2nrORBdeS3OuUfFpLihrbO+fpDHOaRtDutkHtGTT5HHP6YENv
+8d2UGTSmtJjnPCClop3ddLeQWD3prnPSctOKJNhxUelziH/j2t4gygcKhbDcEs8PKbh+S7wBBBf
tBPXJfCUFynLOLT0XOMKhqqLocUrj5dPj0ePWi4TqK6JguQSMTqu9FrwvZuwPVSnFxq3Glt9bcqx
Wio62bBYZ9U2KC1U/cdtvAq6XHW98eTPhT7Cp+nMKV2o+ZbWikqgXJ6io7D9FxQQMpcoSb9Ww3pZ
0HQ/dYIAV+P+lVHIwkjkdzcAKBtU5Dw+ZtrU/pbnpvSNzF1eR4Pwn36MSDijc/T9AmcEua/94wAj
V3zOlw+owtrqLswF4Qn4zm/Ly3Jy17YyLgE7x5qS/8XTpUaJ3avH5zNMsHZFWuQWHrDJW8QlaaG4
7WXR03GwYR7Rc87zQj5Ew9JRnCjsBNkYYRxw1NSSc3yHEZoYsPvdjUrh+WN7tGPWM5QG5i8sG1p5
+UzVzJksOn7wUZP0yGuQ1ZYT9nWH6sIT0NvGNvH45zjBu5bpJPoDHzx6gRe1+RwneBFQ1yG+W/Xi
ZsWJ845PyTzOpR7mPkrZ1TDtblif6CkwjZ1vIl6GRziuH8rbkegULyF2fy2rJqqoS1vfTl7ar7t2
yO/BHiKyVyMlQiO98bPm2ck9U2VxX6Wy2BPOSJZJ+/zx6Mr0fe+KxKGBL4kEfSI5qGs3E9QSZZ6y
WZ8VAqId6sikMf1BUYh+Lk7FakiYt4hviXhBmG1ORsYCtIVKjGkKD91/iuCamcRWXn5uNK5eFRYt
xscEa7NJCDRR6936JWSqTeZHLDTUL+HGz8KbisWKxseIUuraJooDTD97UyZfStQi74NmaBaxVOnU
SZzKvfL36v5tMe5i3jwrDl2i+kmWSAlSRVbT+StaQ2EckWcP0Y1TBtwge98zmVe0U4y6XLfluaZ9
wlli4lHz8GjTvvNDdsngUfaicpVKMiMFLynid1FcQYknxm4FaQLvonJNmWQ30xvrZxzENbjuQow8
iXpYa1sreHfzuJqIMKLoK9Nilb8L0mIb77LW6gRo3McwMvq0ZWxc1cC8HTE91FF+YX5HZuX+jD/2
ODSIUvb8mgp6y3nWqI/bStglbQDRIs4GAFLjFlAABJA9FGnHz8U9QAUZNxGqVA5RadwWlVF2Xtxu
Li1uVoq3EjOv8YPdm1BLcW2lUpI6NUOL3F/8Hotu5P5KRTxmoQGCGwu/At1KchHkTqOG0HhTU87m
yDR+s7FfTfRv4cnj/j6Jz3Yj75/4BLVcR8bo8kMKapN+xCfPboabkWY7y6BnivTN/Qnm7yjJsOur
ts3rl/EvYZlBwpPXvHLIlyETV/C+YjhYbPHDHAt+52bANR37QfbQ/z/PTHa2tfholc0uvwkt4I7Y
GznaliQYKbUQvz6JhyyOZFhRNNiYleIy3HxvKUtq7F3Y0ueMiLlpAWTCFp6OPY1wW8hYHdAU7C62
Jhv9cQ1Clk+A2Rox01wZwYdI7bKqLzdIkVXoeNcwbIYe6QpaTKAzu3evppoY3e9rt82t51O6qfbd
zsspBrUH6Lq2de2YhNVWGhW2v/ETDRuGn3b4ELkCdE8yR1unYtTwLlOSn5ufyxqjrxVvlbYiCj1+
tqnEJrx8qicnoU9Luvz9faBTI5Y3B7OQbWNzvwMEE1HoeS04B0xTOipMST8YoEqB2lNLcdn/q0yd
Xh3gmMTKyRTIqBmo2HmVWOfUSCDhVTgi3VjSZsu/E3KKrdDLZRMcvu/dl2ucWvvSao8esK5UA6Ly
UvfSKL3FB164bO/LZl2fYi9gjRUn6U07vlF/0cxJRZBM0m7nhTpLmSPJDjMkB9OfJwQym7xDnrrT
OD4wwx/Q3WBDbJzhU0xBXz7nJKhXLwjk9MpbEJGJS5QblPMOc/FnoaA+upuzzu3CB9UF+4V2mfEy
rTuKolu0m7xrUW3YzCHHcrrNr0F3eeWlULSzsncwjUzl7GLuCjDwK6wG94HjwJgEw+Zvb7jnnC2r
OOmYGKrnv/FLtCC2alTKjd0/OXl3plpMBuVYWI6kTsoEfGvJIJOr4xOVkcbSdyfj7G4uDnf9o1Ut
f9jl3ITiiVK2TnucpGwwU3xqFAFsVqVmqZC+iGSdloPWsW1gl8ZqwVGvuUUAKwhwqBWnlJ5vzpLF
G/Ff829RI+K5J1amIep8g43MejsOmgTwcDW6qkwri9FQf4OX24ZSrSU9Rxz4UiJlapPz5222kIwz
uqGpG+b4GF+HKutT06AOo3Ta+BvzRd50lyXJflnZkGOFQieZ5+CC3cWt4YmFT2cIJ9O0dDK0o3rx
hK8+0bfKSrJU7/PebP0W9e4CGGfz3Tv2IFaubWTFedhKUf1gVgWRsRNhSXTZ3BU4lXKwLIzgrYar
Hbe6jIjeKx5fhmahu4wyBWQHhF/iY5CuM1c39pgy5R0XHW84JRoqD3StSORdxhTOo83iMyQAw2EW
N4fgR0WVZaeKGT5yOvn2mpcTiCTkKXOeBZ4Px7wTC3bOc0XrsNGQUlyY2lm3IL1Cmg15/V2fz8wX
dfAX5JZEi2LW+d/ePysSW7Y9TtvNUSiVwVlv33ZZZ8vN/ppTUF7loDukGjehZ4V2agenyuYdwQfq
HQ1j/sicjcCmsNiEF8JAqECnmy8UuN/jzrJzOieHWnVLzXzqbAfmkpNAa3uI3LA2GPbgU20QHOKE
D1h9wbQeuJJ9grOs2U+kIxJcJDUMH4OQ/jCVBvxy5Nvxqfw8JpQOQ4mePfqKW+BzyjnMS/EHYX4M
mfGQmk0U6tau2YOfNF2XBABJOZiCJzPtFa+xnASGiXzKX0Rzt0H7uK8ernImNEtTtqvLcoc2SYGj
lFnqrB+M7sYoVCoGbkvcCp3tWPAfj9wISlvIImmJ7DedOzLo2Ib43mLbWl98LfwGa4BHMjQpvCDW
W6djPkJFtXXpNtaMs6/gxizb0JWP4+P1eXjwT+lOiCNbonf7iX22lqFTfdingDRXzWPJknArPg7L
CLApX7sa3gCDi6cmptpBGiLPJ9bl872KxF+rwbTQC74VgKWBi17YnLRwvpiv0H0PEsJW2i1Qe3Wg
l1jvD5Nj9E8DQqQcpxcQvT/6bK9WNu1dai13fP4O7tQlPz4dkpTqV3hqiKjVtr8t8HxeiqziCVJL
9RkDWgh5VPC0q09greHzN7qJ5Rv7FdfK/T7AXXXnUMciVhV3z7v+pbQllAoUsQ67UkwNy10cMukN
UJcEMOVLZKtgi6Z0vIHCaYlvY+OlKt1liSF1j4wS6Hc8FlAZRB5maomyeS7USTvg3mUgc1Y82EUH
JkGeC/K8YXgaRl0kv4viNab9mOuT74VPnQ+b8a31EqVLjDcKPlkdIKX2NCLgp9fSlQwipYmjFm9B
8tdkAuL3jO8JfLq3nKnqjhrUwJNxyi7Q+NSnmVZcBulL0ICs9LX50hBBq7fJp/E7ik2N00Dk9UEh
fz5k25Kzs9v70OCIOQerDcsFDmPskqK+UkC5Uq2nxshrt6GsCcOiDebM589pL+7oyVRCSCE1Urvq
xd81yy9cbplkS6Mbt0PeFuvYQGEOMwalkB/PQVu2uCwY6yG7IJ6finYh8/iobXt5VEOvjEQsDvEB
63uJfl1j0kFENjV1fRde5XQO+okrHBFVRJ6apW3hm69ojGw5ZJUn5spq3TFrfiPTFJCfkX2YSeXX
WkWMyI9y3rG5jhygxVx3TCC+sePa4ZqEitRQL9gz8W/Cli5uMvsv7URmzTmggCt5mRZWsBeR+Wwd
MeS4UreG1JxgCRe7w85BCV8HhDwnGJeMf0BpKqp701EqtCTo8Pc4iE670TYzqxFa0KThTUTvFeat
tWiKrt9Si7B1V6z47vnsGexqMTPDzk1fggyQV6kl3Z0QJSaEL7fCe1tEqq/mkN/Qo3VOae5akkv7
qGRnmATKYDM3mvYuO6vj/TaR0aLibukdsbA5KCYX4U+PC44/nZEnVTNS8KUzIRP78z41MQFB3P06
Nz5oGlKMdHBHypfDDBJe3MxIY6a7frSITU6ExTv1SdbmY5Bw9Q03cCug64P6lKpONCeYXMlqOKLB
CaV+FwmtHYbJBRuiiDxSRFItzEY+ruV+dljAULgfqM3b3TpPN5P5wyVDpbPmlQSz5zmYQOof8w+A
/ceW/4TYB6SW+m6kUEpvTXrLRyhN6oomTnQZgU/7sr9h2k++jG9caAvR8AA9z9ysprOLjxWgTiCb
hLYsAvG1BM6/EpGQXAzf9tSs6Ud9zMNuWKC5P5gayDbuYyOh/DLsjKZfxaeXl+xRQEsoHOGH0dPB
I56vhA9fOLlJwLNqbw0MBQ2icH4P2leBNBxw5+JDgSvJnB2LPVBPSs6S3WrS4I/URsBg5TCu7qmr
eJ+ngI+ABW8k9bCHAeBTT1xYG58DHtIvEw4SUJ0W9VgtQPwzW42CQUARUywiEHVn9gon/Cs6VdNA
zAQik5QtVoIuu1QLHWszCsk1F0cVRaxhXBrv5T/nurGCQP0+X3Ue+ZUefnYYBcJAKWPexUNBpOMo
KsKe2hMPgYG6MbUJCdA/uT+4S69QSszeHewBImZgbDYTsHPJ/WkNoHOGMDZag4Kxyj8BoGQ8xeW1
ZI0KclZdmNadjUUgmUbsVh1rarzxeh8ptAEwVSZGGtT6L/nrDNREjZfMpXNGhxchy91zUx8yGhPP
bg/kNEpyMPnQAj+zuxtwoVvpqKRtbmHQ5Ta/pdaKoW4ybmMIdwbDP9xBWP5Q0cGMN3g5gKnqSsq5
uixfDczi/waMP1PFJNujmG/+wJXJS9JYCOMoqa0gz3nUpHI1EEE6d6MEcSj7r72Sr/hCfv07JYba
aEPQnfj4B8HuDW+hKf6liOMWqzR0czctS+7i+wh/AOlYQiP7LqciSfQbEvNMB/NM6RWXqTaCfdr3
oir9UqA8aEXpwiaXIssEV46GqnzR76qAPMXNXKnWqkIdj4ar6nyDx3fnfpBldW7RAOYPuBv16B59
iN7pgtmgANguJ4LE+xbpoJIOf2cM6I1QcKUABgKtb2gmxNT8Vb+fS3VL77zbLlBtnLVbta2MoeNZ
/cfl82MLaLoZTUw2LCrRgU+/XMcMXBn5V0gFaEZAYVP0mAGiz7HHQBld+2IINcxLwBeKAuZc2gIs
A2F7VQHN7dm+b1jObPbeUQee7Q/J9aHXi6vGQnBhfRxfj0VpilWai7zBJZQmHbHaZnZQdPTQr9cD
hjl6AylHAwTIQKZmUhfi3RVf5wmmHhhX2gQ9YVYrbFoYtyKbrDTMSu2MmpMVoO36gV8oSEFMNtje
mGega82mwyyJPOKuduZDxOc9Hu8QacLblQCk0jtSGrREnbSmi/bYmz/26r+zT4skpRN41LP/yJ+U
UMjvom71HfIRkkl5Nz/8XQ0Tu3tzu7hnb352oivhZRkurs9kmrIOKLbKLLtx8zG6Kfa0fjHYzkiv
fPfHQAxgNMKgxMSq2DJVp0tYNlzXZttt6beB1A8IXclFDnR7nPLns8dTcZdH+Ynvp5k66H8ru8sl
t65V/vs5lKVqwCoC3eHsEE3KEbkhomOYq9J4nbloeCqFTSJ7+sxDdkju3WxWK2fNAcDFdHb0cTcS
SM6rt9t5tm5XoRn2HH/la8a40xwBriHORDQ8/cskXIBrQbce/GhUiWrfBZcyVrCFFmZ+V1gmFpFm
JwAm5wmjK9y5Hn0ePeAQUe/hvWpOy52wxFiK+CavMrC9KrxjqmlqBekfG3e1O/yubMS4/zRQPRbe
5B/mBsATP6sIQ8+g89fLqHJtbIJl5tI/D6LLofL1G7BgaRUnWNaOnRZBMAMxoFMN8BicCuT4PCMb
EzC1jlNJW2rRTc+9Cgg713l0ylzQjMyfj1zg8/8v9ehpTLUY1hjJPQwhWgw0Ak6i8TnU24CDB/Ra
009bxrK6PyrY60U7tjrlm3PtfTSLCo6930oF6bjAohwxMdARQ4gyCdRx8y5fIRXEXNqkVDVa9EOv
XTG1gPSNljg0tvIStXW+X3IkCzT13q7mzBkxh1eX/ifcvrgE4KgQKTLHL+ohSNjlogLRvz/aRH0T
jrxZ2wcstPJMUNE7HRyaE9FhOhFa3Vhh/hQZ+SNaG/IJv2rxE4FZW1VhLLp4QhI3olKzvdfVYFXj
16wC4DmaZy+92PFhmiFzktSRpLerdg4ulGZoBzs5QSruoFmcaHkLqos0GmzqIE6kux32iVVRyAtY
AHDivg/FSqhwPL4S+C9rlsKIUyLjcxMgyV910qoXW40asgyriZn3rH2Z3KCUT8/46Lq4VD9sujtX
cISRVVqeZ2fF9xc4LOYHPs0Lcq9Fk1+4rD53nrHoqoTFgXHlE562dDdUcvPcZyh40Z9DdmNi5APY
buT+FpUd+AmoFUskDaOldFdJPxYL/bey4IkNOKKOqlG/y9/7vXQq0I2yzHCCTv88iN7BIQafiEkf
zx1DRS5thzFf55lxMTjIkSaY+Iq11dATfJanrsMbvCY/GrKrVXlCTWaBPTa4rbs0Kyj9NL53gYH8
5qsauhzwRuNzbONbtGeXJxlWcRK/sCCbtcas1gxLNGIFXqaGEictBQHj+I9ddoqTmt+oC1vXWR7c
ZiNPT8dz3an2l4sYzDqJ830jJai/jqgFJZ1OmiwVwvHvDTYBwIhQuo2SdyrqFRX23NbMn/7uMBW4
5QLrtV5mefD5dLj/uV8zyh4d1qv80tctwGqxD/a70utGns/+JR4UPvhPAJbgNVKDyB9qcxDhenpL
4EFkjqapwTWfDC+Bn2NNJDTCdyBbFYHMyL2u3FmNCmjWClahV9WZVd66xT4CzPnL6hPQKsAJaTPf
b5b8Ti03IKhvu7lTCrLm9/rq9suwaY4xkFpQP9avbGr+S3PAYS4ze3lPHC9dP3WkUUOvLQXwzkH4
sSiZb7Z9SkBjqUfEDvFaKuX6znCCbX0D4fMf6FD6t021oyj2y5diBVUZJ2/Nidt1QL4+wkht7m2D
QSVOiTZnmx07NWdTvX9Q+NET52Gzy7qaTs4RXuvKqDWDWgeACqQpwyWbfWR2vhm2r3HzoMGzkfyD
pkNHJGO64X+1DZTy6FYpqp8/6Xn3NARBX7bNgXPI+t16P7ZpEDr2LyrB4/24E5Ic67U7Nx57EHoT
lSL0pqdJZqy+OlSKQVjAGPyGrlEMEjIhTDrP5XJ9B4oQNwnK71Rpz15KmAHqBwQff1MZAr50lctv
EBeuJslHrJU2uhBiheodTBG4dPavbZWjK1InEC5IV6tA6jNvp7wbeQg2KWc5d9hNE6hiy9JaVeLz
LjVovzZk3SDAajdegj7Hf7GANXBpsX6wHgDb4Q0OGlNKsKLKk9/7ykhCcUAsh28Yu4zI0LiaVd5d
hUtCoO3BGYA2Ren+ko2FWLkm8toxi8eZz9QyEKCxlvs4a7r46MN+eNP6Q+xmwmd83QngCesE13i7
qiKXQpMNP3dMorKXoiYG4Bc0HqEmW+3QLYBiUuuXZeOgL3hnOvJcE9wKFj38fvPAyMXarf7/DV3I
mlxLaEULt90kuzCqGdjeSXMwJGXdVf1+TftxzTbAzQyy0LKO1xjmbgOblcoAfH+RG4lEo4/UDVg2
sN2nrOyDDcsA2xBTPN8wE4wx/SzU4bBnvz0hwgvXXDnnpUMztZD/XeGL7E3PLCMaL3pAZV++0VKm
hViD8csbLrFSCs8fix9uS/3rJeHw+/Yf9FuF2fS/iC5sgt4v1KV4mlGgwPjRrHAvX2Bt2B2vuo9H
WmmIPGvKFblmTMTkQu1c4AkNqrY7WDaPEKOaBRWhx/A/LtLx5W+v+RmCkCEmE+jikKz6K/sI1ZTK
nOYgEJFoV6q9iVgw3lqFOlcbIKNJC5jN8s3UJ6VipcHU96pqcToirNpp7FRaBLDxtEPXhQQfUQ6O
mSg06mRR6Ya98I7si9ttDmhatfyRtH7lzrpLajSQd75Do8xX7c7RPOb75csxBHo2sznH2oNEAKlR
k7CwXRGc93zXz7BtAZxBZy42QxNFkwF6QkxLPNxka4gdTGnndaaMDGHm4ww6dqMKY0Ce516Z2EhT
XKZfoY86CIewRqQpSMZ53lo/jXWkD6Q1CtA0nN4kr9N2YW4163UqRbPc71G68YaB7xwrKXT26iUS
7LPtY5qCNn0LZkVM8t/3U36DPXzacCfNgEqwWpRESwPltav621PyVA5hWge9QpQlHLTV4SpjfTtI
c7tS79lfanS24oZ/mms0WyFtF9y38LaBctMVQqfnrJoocROmHtQrk5KE+fwJfPmflsrOGC3jcwRg
2hG+wcg9FFUIx1t/srFI3ICT1t1XtZ3DR4RaooHJsBuqwG1/daI16bQZ+wCpaSv6VuzR9xapWnQm
wXFq28LpYFCFSixw4tY2bMbYgLXz0ijHx40fnEVX0SfRqCYvaLvuiyx00IQFiUM/64/4aqMt9tdO
9jG1rizFaCTMsgznUvfj29KqL7NP3YGhjY896kgr2VC3oUHlym0ZlIeVSarlXbtngmOGmO1uyvTs
g1Vm2yQ4y+bSNNRqRMI6hqrFRvqwp/WmyfSSi4cCoPApDhxBCYD4b9CQmcUFcRcxzTF5TzTsvHEo
iueC8mGWT9nNByLIdkE1eq3rAN1LKFiuLQ/xjCrbTnhsHobyplvuZk/wdm4B4/VIvwRZLsfoT5gu
eoTU5a0bg8v4VZvUF2V5xJIDt7exbbXnWZceCyjE2t+mgIIo9F9gjyMkfNRwJtgwufpe3AIi9EL7
j28nCWtn0Slasfxo6YBgTaEg3kZy1UWvUiIJZbId/VfyfQrPMyD29mNudPnjs1mhpSTxpuzNsdXH
SrGNFIJ9DZNDPdNwJGq0TdhuKURFcIn+8gvy3ATXMr9hBWYEP1edwa8OjGvbvNDbIiZPa7KNXbL/
CmPtPXJlb51NLV3a0rncLzh0rBLXZWTjfYhoNLxW+xe0w9wLZWW+flMOaRWjUQNqLqU859cv50si
uvJDRBSBqucm7ETcvrWFtRxVSAk1YFvp6n0hHO8xOpGtCdeYmknoufiGtsMRqFbXsoUi7PRz5Wf2
nltfalGgpud0YRcs4WAonlDXnSN6vq+SMiPoYiWfS3pWe6OXUWGtSix01SGLfT3hEQxMMezGLAHw
ww1knaJ+WBlfFJjv0QLUBVLqTxSjecT005bnxG8dzzLOoVLg8NCxTv9sorTvdGizY76BfXrY6rR0
HQGOk9ylTmFboa06DM0LcJ5vb35wVnLQpoSsr0dB2GCPsM2Z9QlS7bKzq2Nt7SscKEV4mYOeE0Xc
1ObAXHKe98qIS1uvy8Kn7DijkgJT7IuU5vvNsv7ZB9Pa+S3Fp2T0H8NBliRiRCqe5vL/su578ngJ
y5gbtPLRBnTXqwqxAjQQxZ6zkLlcztSgw5y/8P1XWAcC9Cejl+pI0rH2OnmXd7oDoz1r9ws6dpQD
ALwFF+kWFm9EFB4F45DRlgL/zlMIwTl66TQ1e6oFvGQAQv6ABacEKmjtIfU/f69wyFQcKk7GCeuY
7gDXRoa2kI7pGB4Lc+jf0iDeVoyBdQHnZbJJfkU8fa3qUp/b5RFN/C65Mrokw8n8GYzkTivBOCua
nOGwzMj9XS2msHV8CM72gVuCSW/IE60/0G2qAx1hPopO4BVswLJWfCBTcvwmX3fSPQ+UUR3cGZ4C
Ea8tuNvJWD9wbXoATD8W2gSOFlrrE5imDEnWjMU4IIWdixPSt7t9DThJ8sv99D9eYtQsuMpXdER3
MAeo+h722Z9dw5YwGP/QIHx+azyaNK9N4mztS1E3DjHLxKqBGvyBDOtD8EziwRUiNG4Qavcpq5Q6
9w1CR8r/3qxLZNS5QRwHJ0S7Boq73yh9yqYDngInkL5In2uLYyY81PntrXdqCCEbFDi3q9ptbJJB
UgwbGj9So632hKxxJ0f/TOXq0ZMJ1OxezhMGVNiX5M9kyw+JRmOv3N/5iGbtuVOpT0yQSdMv+F7c
GD2f3sxNljeWMuCduH0W7o3UXP4RFdYaByCBWrLzVmmJc2sSl0hUvulKoB+znW6bVwNvYqTfpF1R
nQy6i5elE4MCQv6qPDhkKGU0e8BNJrsgezaBaaZzbVArc0z5r+i0tiU/1oDqqXnq9xfsMxbxzUGJ
CplugzyEzcCVOAZifyyGTkjBwOAAM2hRgNxXTgXxuLNfsJTS/uRpCW96du0VnmtkSBzMAx7/ECCY
PxUKkeuUelbZ4yCGNYxKnSS+l0MPvmLIWW6qTC7l4pfVc416D4rCnnW/hK1qBGu80QVBNvUTULGe
lM4K7bb0BpRgR7Jvh5mKkrLIbxXKHTlJa+GAd31NJQud4yNUvMueG7a+SUNvOKIPxxzBcaGM07CG
G80XS1IA+XeQszojc58M20sc47AzwToLH9yA0nXmVmqDPr+h5q6QsfzzX+0yA0RB4207fjrSc90m
38eKan/OfhhGne3kmYcGsATK4c1wPv66Evu6fYFk/dR9Ylf9b5qg/n356fxhPxyb7xV47DXrCuIv
R4U/VcX2E2q8q0/YAAjbFLjc5MnFQN1uWahwHGOG97Nl0JDk4mCiT1EcMfhZ74HxsnnDVVocmsBt
RRChnzz3l5ylid66kjIcjjJIE/QCVkX9/c1ikIQyPozHdxDYfg9YU18eCc/t2FcEYwWsqKAojsDv
4YI2HECpWWQ81NNXY17iYwXc169jCq3ab8BEEey44mk0RTIZ2KbamLQfnotAbPbjup9o3idZU49f
me+kL0+ZmkhyhNdwvKA2S5r3QbZT7R69YHpjy7/P6621rhLB28LPbgYp8CZgJWEoNU1sop3RWjfQ
l83JKlH7C6TfDUbCG0eSykCaBzLI1lV4sQmaAvfhbSc+FSgkJI3QtnqaqSrL+otUGg/u3ifG7kDY
tD2wI2CAdSjLjxtopb3tEZZBYwonq4wlumQS7QvcdhgY8x5uEL/oJRIRtIN8go0auMM4VQI+d0Q1
H/vLtz0N+dAEUD9Ddn34vWDurw47TJNL99/91/lFAd04wyKdUpgKWbtf9v9Sn4nAg8AF1ABBPFLG
hURIgxMZng6H05+RwYw2IBIsaqMFzWkwfqDHT694+FqmAUzvXqr2ZhJt+ybSOKpucCdPGqzcfYRq
rRY09DgWSjl/6aTj+RgDoTiEB4hS+ooTNp6inIVfi39ErYYsKH6DnCRylyqQihbqal1TXDNYqXTe
miZnXPNDm3TwaVV/I2ff2wQNVRiMqF/GgzKL73MxgfXfXyrA3RIvEyufenQGbqjd/CXwhftzHLcs
gsK+xOu/rMh6LEwixP9ci3LvCRM1jpu1WuxikVv72NZeHVbp+dkaKOfz+3N9QLAQDtXrp4Ris2vg
VfeyBPrcpkppXIy/7+JfntyxwrK/bjiegtuGc5HGFtFyvqciaDsbLKtPz0hMOfplPoFysWZATsD9
OFBtBogPA555jDLz5+478uCcDyUeNfmh2tTF7Gu4GQPKNwAJF+rLtvWEjykrQJIH/rUFca66c5G3
rbVqOEFAa5idsPNLN3KqDqeqKrfi3HVg18EkL6+Qg+CdtmOgSGltwkXjlizznNUii7sSMQy7AcQP
KjGQI7H55Ms3iRgFBlnKYe/meV4fH4vex/q/H1v1vSxu1cqHo+lJWOEF29P/82iEvdcNcmj8Dt4J
u+vhZtlMXbeRn8pTmdq98nmCNGJe7RjDjBdYdepFJqI5LTvDdniLIbEN2D93tJFGe7ocgDOgeknN
N3f/gk9rzhnOhiN5dv8he9VOBGbVRBIl8+8J478T8PNmWqaoROgUbs5YuuG/mdOdrRpJlVwMQUE6
vp8pZ2Hq9xupGbUgBWW1TgA4G+jBLkQF9RIaAAm7H/l5oldfa5YtwVQwA6arvEw1ohHy4Wx/FRKA
6Ivwm+kbRGaT61zLZql0Mb6c0TYkUJEv91kGMM58rxi6H2gQhhAEVvejJb1N9x10i/8GdGsj9mV+
75CN5H/M5thQN0/lUE+7sITmfx32HBodVLbM3pR4myt9dymDilcXnVLVfBXFWnbCr2+SukGAg9Ps
xuTHWkOwog51Tu1XNuc/XO14Z06bI/Sp23Sfq4rmNEqgqcbTnst9VWBvBaZTYws8Pg4UtbtX1g0Q
EKEqfOv8mN9YJwxv4WX8fZaYdHxHX58fI9qkSLwxVqHODz3BIl/odwxMXtK8j4tvZX3G8rn58dGx
cipiOwtHetQO6rYhlKC1tqOg6w53FpOYsQ7LdT31kG2vqCwb4PvVsKpJwB9r1MASArL2fAmJpL0b
h7epWxDvmJfdQ3HKDp8SgW0vHZBMgAt4Yp3OozI84Mq88LfvzPePoIHbd85OtcdPZPa93AR0Jt4Q
gdw1z2O7gwAf/6JeUnxoDL/+/gAWoL5BRtLzc9G8Ts9+pweRHiSqukMeoxgYOEVGSyLyAShXxo7B
0z/0/iKA1t9y1+c249dapX6Gf19D99uMSMgZ2RTG0f3NAjVV1X+R1dzWeic5Cz62f8pXruTFbSqi
mSiAzB7SCXUxPwl0fXwlMeayL3ZlxnK8IZELGKZzU7S3IZhtCFo/QKeg9JXbkMVy77CYBv6Ed44v
9RCUzHBrdVQq7QsGYp9kwg5yOvTg8X8OXoqTVm7l7gT2+2KblgN/fyEmNQkiSWgvOxkGLAkjE7YZ
nbevTN0fr8dV0DGeGpJ0XnhKV9d9mxGYa3xB6q6o51xE+mf14yLln+2jduFvRvNwY6N6WE83cgr1
tCXYtPhDnxo8vJbDt09CyAhEWL3I7eLuDxAaZyVpcJRkg/jDllpldgg259T5zM/0lr+UBGRlbBJm
rxWPBoLFK782K1xH0nodk/DU4x5HKhIPEqG2miCh3uDDrAGIo+NYl5HGPE3XzTmoyeh7ThrkZf1a
YiAJ4BSHU1wJ1kDc7+DBHjs87TY8H48JRQ8ooBangtjS22rWPUbVBufp0eMzWB0PU2x2dkh5+Z5z
tTY9jNOUvwjbwQGAY4D/UJUBMAJb1DpARgBPs/RlUXy3Tt257K4X/mrihPKwp0FX8ZX5wiWxQj6h
6zIrZ4DRPqSYEi2gsL/wVFQ3lU5oT+ZgkltRVbiME4FqAjNjdXhgXNBiIDOGGg4PeQPEOMmzv5DS
Bri7YYsRyWCpcvmz8Xm8e0JPBDtLZpHZm+F22KO4MRDT/G3n8t65z564ByP26jTuRbYWaWnBT8/X
ellGln+PhFrIIzjvQ6DNBYsNdzwdHQA4q+8kAL4c5WtOQlfbLW1e4EdmVchkGkZGViWUm9D6G1O1
7R4taGSkfaHBdEIeS3L4QvqNyngrlaOL2yXU4CogSqRfcE2OfBVD0ut7bVgKOqB1KNlG671YCZ7s
w7BnH1xSuSiR73rM7LFIeZ10yHYT1jhv2HadN+39sXMq+cKygMy2DsgKmcve58PD/bnEf3sCNSv8
Kls8reSTdZbnjjjbrmJzKrtzT+B5Um8uhQh5ez8IcCf/2oCBpGsm0XegETNwv+cFcrgLddHcJmWi
Vfnekuev5x8XDKx+3ubopajF+mcBtp4ZjfhKADZ95ipuN68h9t9/UxUo1LbV0iNLccCHiSAyTbYs
4d8h5CGll/r18l0fJrbetxwLrZtbcue/5H1jAuf/bJ1zCwefDkZo6wxaE6NsMn+/ry8Af2BGaF6Q
C65VEz8WEM3NbN+LT84VeLvmtcsfdK1ZP0V+/MYZNPq+WZuDk69V8qhnOamYw/n4SHKNL1z/3eG6
m7oA0bYv6AHuBmQnKjd8k7ehu0tHcIZoq0Wich5OSo/dMJvS8ZPcab/gFNIbVknT1iTNjqqbsHQk
WC4i5l7nq2xVWDdOdPSgBPlwKNe0eRcQZfePAlEHBsv/3+cmU4w6ws2EqYc9gGYLipM8JlTjfWPd
c4Me+KWx85um2DWvYmqGulNjtGeQc2KMFUIwJgaAK8HofhCIcxnwnH495w4Xi04KUfAKiTtW8XYy
tkWpdofr5nM6VjePN4Coc1t30WSXA+HRjQxTZ3cQbQ4blJWgA54mnsEXXhtGfO4IQUVishilROgW
4FexHMhn/uZU2aFlBR+kQ+aSvERLB3ZfD97wh5YE+PFfiQhKxJvqtWP+JcyUGpvJdsW6d82B9uLz
h0LQ8oWKgJzQVhYgLxW+aASPGqV8GQCvy+h/uPVArsc0xZL4nHDnSdmHmzm7KhahgwR1Zea5XC+t
gYbd76TDwvFTQio6TPf4B9TMo4zscaAQBChmNnuUfZOZF3ZvICN9f4+2bZFPRjBXSl+8ITWGw6Uv
RPqXBzSRjAj8zSWdU7IT/lO01ZqHuDhS92Syq2oddYGPZHEmvHYHDOEj2fVJMN5m6N+W7pF+1US8
TRyWFXV3RzHz/SvzHK3Rcd0mcanf2XZ9WIvcIeuArFRQJTCj486ybR7/YlaSCQ+qtlspER3w+eJn
3pkBEba7VmEd31f/diNk0FUgY8jYeX3tjU5EWs7hYWG1Nttxku8dUVc4nXn9/9nczkSeXmWEqMxL
RKY3O7AveCRAsUwZxYER16zQsWOvHh+reAzdiw3lbyv0E+VHEXturc2mFrB9O3P5lOwlVU7Yu+jf
wAgQuzdKgkIMQE1HdT/srbICEoVoXzY8GNuAh57puJtbBKPn3E8AULGsRZqgo64HNCt+ljyyCf5y
8fH0YOswnxk+YUHcaGaNTfUHe/93+6sLOrUQVVRMXNkXNaItLy4VjaUOdMHmWfSn1Ezfv6ZyyfSQ
NwcLM6hHmY50xZVx8Lo0KNJ76ReGgu+mAwJNSTajnkZOBFdhsY7G5hDQSSmQADMIocsTukN/rhHj
3J6mIzcHFT20j2UX1bokHCVNwHbi95SV7L/c1NsBp0cuQq7Rlf8x+ut+UoGRXG/uIc71waFkumgz
bxrEGkgQwNpZoc1tSrFJc0cqQqrzpkZ2VF9iYgxxs0R1obb3R4zZgAAsha/xHg/QaROGnLz9YqPM
em2XMpqH2ZCdSVe/oLWVKDA0whznDQfjvK4zZDi+WXN+XASn2CiFK6NxFEK30pZhGrqNw4S8yGHp
sVU6MnJCh/Cas0X6z9Lg6Q75pDQ7YFhM+pcWm6/xZ2wu0CRv2R6hpdfO0tzJoPg/WjfpehwfTJ7a
USb9QWAGHLZ2L7FfOYVQWIoUtV3nJ+5uM+XU3pcXk8nY79HpzPrS+E9QjtaVM1TeUWN5aO2hORoM
vc9fK3FQV7+VxUBKHBwcdobf16Hf7/4/yNpBtVgaKTrxR1dzw/Luom4yeUMe/y57bmsngkUO4VkP
KsxUtHX7BeqylLljp1vMAHTrWeMDyMOcjbUyfdJoTSmGWuoqulb2aGcwe5HkHkChrBYE3AKUqx18
6Z1ZSdFzHzm68izwB6yu7W9QeGhQ7T2EWJLZRu6iro5coimyDMD1FboVfJymZRZiuL/yxKKbgUSt
muM7PgAGdvm547phh3Y2GVgwEcY7+fW4G+7Ji0McoCxe1xkRB1YprtWPnQcJj/eSsNzmFaYViu16
8+Dlrt7nO+V9poybPpnx4qHMcM5NHgM19AfeeyffZc+5aSPh5MuhMnNrMxWYakevCITkUsFyUXG7
cfQfu1hnvf9cCZt+35Ln62sk0ykpFeaZzLdQDf+1E9zQXAfI51XS8pOc1RlU5lJI3CG7zYPD47G4
lGP07VYJDEt97kgtFZo/k1s98Okq28FYQoCv3xkbgXHu8lOHTR8Qc8IHlYOFHUWtvSZsI4ng/ysZ
+Fj3tj8qjUYGYmZKfDbkruuwt7jjc3Xcagd5UBkTfq0hH+iw7NmXN9vzUA5UQB/3nNtuzo2jI0lV
e9tvrIzdmQk4ina3G+3yyqovbj1PKKbmyehnB+4JVVu9vTw3i5ShAeR0Q95DP5t20l2KxyRHABbA
4eXn4oLy3OV3bn0h1uhMmbKYICRBxpRuzDHuOXV8ZhEyAaWH2i3ZkJQrPB9sJvrR4wdS801AGiep
qsy4Myum2XvIADHGnDYgcWqQuwDtlj6sLVLJdbLU7c09JXI3LyCb/AcDxog9qfNbha9gYdXCsLMP
QhZ5ZluVj5NXTb48Y2BHzuNCPhiI+ALrVz+/NLA2c8ioAASjEDpGAhcnG9bP1GhUShWADEKO3pYI
rpK/EHyasPestFR/IrVQfCdnILlnqOva8g6lUbG7geeuErR/kKrIbTUvWhJJg1BgyFimEeMokzWH
WCbZL+AfiJ0RrI7Lq+mKhucWwA++734QhwC8SUz07Yz3B0ct0hgmdz4J1rSqHKtVLGnP0w9fCpNO
SBDbMTp+iRkmRx4q7aQBKgCdynwy1Mxs/x3QQdLM5hD4dYohCNVf7fCJ9asGY5Kv8RB3HjuH04hF
uiLabhtrRzR64M8khMJDLNBAD65Zg1hZAIG3aXCWvRY01dAPuH91IDRnhOZ43R/ZPK8DW+SQcCgg
4NkFIHjrNTcxFV8CPolR7fiS42pfxJcuhtR18KbdyQ8miC4yt35X1Xq9WJMfZulNatg8htgSiIs4
5oi7LGM1GiZsH1NHN4d3VXopWqKMyiTrfWwos+codOIHzT1fKZSpZ+oKCP+6ug2RA+KMAW2EWzx/
IL4532R1Hy7uZqAA/uQyGvh+mmp/1c49+Erxr0q5+fdPEFDx7L6NcGyNj0XYm1QyaMlLJY4NKefc
YlImPVVcPWmaICekoSG5XQc8R+i27+QlNU1EQXOion3V+YpBeyJPZLMxbTswb93alDQbCJ44sJVO
jEL567X2RM3Wj+Yo6LQmoqgoPmQLItsmOMOE6Y2FK7eqpGKnRiOjauyRB24mOwZjvrKp7L/6ST2/
plV3TeMdp2ZXLvIiHkKE9Qll1VkzOLGyA+8RXudMvjoorptHdrrGc5CPuxVPXpr21QL5B8E2WgG0
pd2IYw78kACZ/KAKQz857P7E4zOBNbWDimo0BRgmaFbq+LzZ7zUMQapOgeDUsnfLGT5Ozqy50u64
k0dNPhkPgXbV4ZstEG2EmlGnKSBxOeZWSLxPVvOjykbsHjW7pJvfEP6ftkc97zonOJFwdSWxtZJe
TMd0o9/pZof8C7vwqpulT6+R6aOHfFDmPg5F7IRRhk16DS08BFUlS+kW9OsUlVVghWMkoE8kMlZm
cgbKIVzAOmCQOoAM/Jct9O2PY9nDZU2GQriLAgCLouqlnwAyZN3pew8S9hkotLKxMJhosAso875/
R6iYKaK6wUaPSPV2cW7IPIw78p6BFIpH1IiKIPmYuoiUwxHbG6HLuNVzfdfezM4X73VyhsqIFpJa
9IolQLFZTPPCFhSMV9DHs2Um9I1P3cy+R9uolqRUJ8M4R43jXtXJq8dPzwqdyNEyODrvzjVg6iN9
0panQ5Cu5vx3eUqD/USSZPcThVh7p8T+CpyIOEKReUEi4nv7BT5+GQeMjcOUp9HrU0S8h4oMxT9L
YJ5ZuVDeXo5RXuONBMUQHpjow75DROQatm7SKTGXtV1wOqkYZGjtqdGdJCbnCAzShu88jknxoHUx
us2RzTD83Stiw5sD0iAJez3h6l+qj/1PPQDpv0dVYAvTzds7bZFkq00lPlTcfX1cDKEuevOxaUom
pH7sEyapaMckI+jRW6zhb+mXM7n4r4yLCi8Fu+ZOC0tQ1F/zFrTDomQqxa9qI/lCee74VqTzIV4y
tnvMpvfbxeU4wzdFrVZTtnDqIX9e9erS4kKXSqMv6cuGI+kQEwZmyhZ1thUOUQGGhzZG8ak9Ungq
SOo6QVjAKLfpvYUeBjUz1KgVLas+L2LGUwLY67pCDcKPAMKRHQTBx4sqSxG2UwC3blZi8IXyo+ne
FxD22ufC/EHw152GaF2eN4R2jR3UvU1dAvulFQGLZBX3zKHScsHQ+iE4YLDGgK0E9DHfUMxYLiWa
JjhXTbJRt+MbMgRIyAkar8uQTTBxJE00A9fj03lZYb9inxtgIbs7kMGunkA9AWHV2J19YB4vho5k
MS2SxXsPDp09gdcFjOm690XYTjTGAgHuZFcuuuJoqzf3DpBev0PUWVoKzRY6yXjaNaMYl15dnNWS
DvnwRSHKkPbSkWBxW+UAFi5JOZ8c9gVtg2V3HgxTJUl1SmkflrglsVd3a0E4cKd8UUwieORvcQNs
O3Kn42FWfHiNzB9vhW6AMmrW+Vw7NuKHdKMDJ9j+xbAJhSIJS6mhu6ZoIjAJgrlXnlLQgm4V43Tv
c8VU/u7dGIj/7T2Bz+YQek1YmBG6MgEuN2w8SbbnqRHERfFEx54U02/jUHRP0/FRZL3oK/XjFcgv
zLdA8Ray/VEZHoWJzeXWtqQG3PoFpvICDtc7ZRV3dmCzoMLT0Q/2ocOhv8gUeaHLbZwHzE5OPTNp
1ZtKQGHRcnjGpBblrC9b1QVdQLou72h2ePwKLjk1D6v1xpTk1dtAvK92EL8gSj7v5yx2rz39ZwAC
V+VTROzrki/CflUBrlG8EGZuUAtn0QazugzaULLHn09SLlwNw02lNuyiUGk8uv+UsMXUIjPHHlyQ
6yRoQmqDpXaXLEGbpAM3RfyruBZlwttRhwknqx+8vUDLV4yZocP0VPTO4AxBQBg0k8KFm+8FI3QN
9gVBWgWO+NzoA0EINmY9HT/3AA/P2r+aXnug6EMh/sNM3RrgHV6mhDNO98ej7LFf2LcGaFMY1dAH
6eie/TZvx8ImthY46GLGmjlHpUkNabQifiW65g0OH65/12vL5GUzXrJcVeZP88P3wDihzmVO9D8k
LSyphF95UdzBJUpad+mEx62KaQ0nFydGK99eqEjwt/G3mudiZuNZE8ruMtXXwDDA5dWjYwJqpUFx
Wg7BVjpwRieMKh8Bavj1igugOL82ZXaPeVyhC/26b+z/aJCE1jCLcvktMAbbmdDT88jJGfBCRt1p
R0rRdIRKM1/Nu6moo9uPpo+ngp2CRAoNhPvZfcC6jqXo19EBmEbUgpnqn3ednygCz9dKI4pJ6i2q
5lYOyYWs49qa6zcuJBMJu/lWXwqBQF5KTskreEMUFxpX36zXovkSpvYWkx9BN/XFgbz+XQKqaWDj
TqaCyibmhNwFE3CFAns2osyndaBkc8V0Ka4VVBdPlj4C7rps4LnVSvAKDck9rwo95ztobG/LcqX5
vQ2LwdMhZ9AQHPVDYFpoF2HL4uk/8eZOGuTyjspaZMolhxtmRbArlSFUuZkO6HghwhY7eBC7usCf
CpSbIYBFrzL19h6gXN7pwJYE1R/2NHKSBblA3uetcf5Htt9AmNTcK1WhtODyqztmYdjmnDHMCE7/
Sc2o5Gm3G7UCSzlFTmqvgYDX471PjVY+AkAECrksENOrcstQKQm4Lv+HMdEcJMK4BqZ4SV2h7Crz
Rk5YwhwJ8GiFqxVADxR1nyR00h9wMORpzuaN9tkOx1WlRNdPrXuHCFnhIsRSsSk459w1a3CSa8Ej
aPA8I7g+FMNQaFoFPRsliJ1l0Tt6PYoN/f/PpiSZ2UmMzadYPzhOGxxl+N34/o8IeUvXYpl5m8VF
oX25ZQfVD1MJtW06i7tumP7NfOh2qfSuzPCZMRpR5OLEZ4VrCcSR1kd2G3F/COfLInV/zTi454BB
OpXJNqXyr9O3A0LPcBUzLY0uXNPAvQDxzlyRtURfmk4LgC5GEikjTLiwV19yfkTs5rMfF+CarH5n
zfQk29yj+G+eSxnTBGFXFUG2x3QKQwIIVhiMv0Jav2QWzZcrD2T/5383/upnR5D13ym96/Xz7Q5P
1D42dN73h2GImYvKIG37LuPxPaAvxs3EBFJiwR0BHxEqkZiXNH3HglqTkgmDoWTGwKIZ7vWZzp8w
gzP3gqGInbPscV+6AVJoj1OQpG5TbLR29GRxVbpDkXnJ9DJUiwphrrnegRQKFYJkiXiIh4Mcp12W
ssYU4SZHfycyFIBQMFCOmQcgRy3+ryxfWqDcnymvT0eFJCqRXaDe+DsFi9HgMgUQ/TTHUZ4WpH0u
hMs2UKvZlD6eY/Cjkic+1znDLNuBtAdygRDNAV3Egyv0DWwQm2YdikVTn0Phu47k0zPBq8UXl5hs
6LAwzaSXwPQRIVaTsZOqWhhMytb5KWzkeF+AyW6f3YWIqPAC1hx7eAClI+wA7Lj/4FazesXE6GhL
uYmL6dY5kUpmD+8FJA/qlenPQSWQAB+xKtVR765wBZk5cOVJfvgWiBEEaG4F6Y42CkF6/2E/tarF
bD+tKCeboykUYVWeJi42wxyYo32WwhvfrBO6SRTdiOX2ZaV6iGWQbxcfmb76ad9D32TCAT3S/vC3
arV/iqin0ZF7S1QT9cr5xPSgU/M6Yyd/IcFdkCR3YtY4ZmKOv5KjVi/NHspVzg4Fmafoi0cigE4t
w4XmLMN6Mgwd7gDjg+NcfM+cXaZuh0qUXNtNIDqgN6Ek34ygqVrp9KfyDjkBCQXzDhYJO/2m610K
11PKEfN3Tr560ptTMiESEx0Fbi40qKQyz/jccIuXbLQhmtHsDCF8RwJG3kgdYLXppdD1B9aedPQb
DHM5y67k+c2HvuL5RvDOamKlxmtzt5BK3elf+JGAGcLs2ssj8VTNdAIpSCKe7FEr8VeiqNzFBMri
5Ay7Bp10e4sxdq0ID1/WQ1uOYNglqUP1XANumhC2cJT8EAAvERwWIx+Mgb6VVcpbO9O9pGjM5KMu
N8fFPJc4pFhW0YW2sg51vZbAl0ybTiqJRfLXtpzGEs2RH4xoeUqQQADZueffgAkASL5zwcXCu8zt
WodGJ0APxWoNKNj/WkZ6SE02S9CkPLh219gQc4MFYegBjlpV5l76C9gcoWWdTgbgwlMDEY1VeP1E
D57s5ZLj30dvbwnTOXPcVekRBEzfsiqfj7uO7z0c11jGrqjMrtc//4SYKAp7b3o4mJrLAMXdm2gG
k7Tl2Z3Dr3KjQNGJ6yi2qY6L+RaJIIJWfnpyDnqnhx/Zc7mQBTjy/pwb54O2LuAr3HFezs4cByi2
axDHoCULXD+DYQYps/VlVjtppouCT2L4U6kLMMxiyBnzL5eT8hto0Js4H8chc+/88eedVqAn87fR
lrneys4K7fU6szPdk/kTsv9dghoWJM2zsP1RAE7x4P7/me3enTSZaP1bc21zmSaqupEl7TIUpg+r
3UinfB4jySzHw0PmAdmpW4BPq/KXBJa4bizM/97GvsTCzttnqCUjP4taX2duNvniaqNu6Jr51lts
kU6DhW+7odH86P6iyN7fK/B+Tr2wBIJB1UjQjrQhKn0ZqEgqzrPQ3tAT3ytXhL3HuiiBaeX+oZPc
t1/nAw8/ByU5OpMkCe8zb6lINIQb59IsrFIR4gzAJyGBkvumqJi8wOJBCDBEXprR0868+gqZ8L5M
vSG0lF0wIwp8PDPeUnfoJd99YF/jbYQDkUSCDf5YKPr1zroZqIZLl8Pt4kpZCHfXwY7Sayl5uBQD
6xMdkVWPuquifrQCNVLmAMu1Pg2HgdaVJhrUtN7rbUI+wml2jxGJsWLiB/YoNHhH/5nkNY0XtuZM
XuMveS55pfvB04nnGkzEyyedyakDlOMj+azapIki2XdzleQ+ftafwMBNI4EypnFrCyLh57dg5Prm
H0JCrOi8Mpr/RzE9sH9DPRir9OwVj0Hy5oK56QDRearz+B+WTcNRkRvIiLYMHJCuOnBJl+G3vi/r
iZxuLYD6Fj/54rLi+61ZWIicGS5+sUe7QJvbPzjPLBufFFfg1lYIdFFtqtLxK6XWSW6cyOJdcUN3
Guycyu0IqjsmTdZoBvp92hExKcJ4/A+08StYG7pNl0qZZEJGiVV3khnfOSvPE2eq8XgKVox9Ibuv
o02fpoC4iC7IWlu5IGY2j2Oc5AEGz4fQBeiQ0NWHEGfNOAVT4ZsNOZMb/pGKhsvqzrocuzatD8wE
DCTgzW8LlUTA46qY+6FMd6ntFfhupl2Gz2OOfHTep5u9I9QMwfU57A/S3vr+PwDYUL+jrUt5V6N+
NPJGztIRdI6d5DPls2rzrIKz2VqaNUZLAH4cdYwqHxX/eh+9emRKrMe17TNQDgBWh/iq7PdU8U86
1zxXTpnNoVMZkjcNkHJOf3b7YWMX6JB7VSwuBoDxqFGJmwXnojWbvO7nWmBodRb0wIokG8mU0PMv
hObw+A2I4HVlzrq2UEmL6obYoNw6gmolkElLhR9r4pIIfBm5dtgVksTPVDQ5Syj/zmBuhX5ptjnP
tvU4CHREJp86A6y7rP4wCMXVXIueb6XNMpwI1C86ci5het5gotSYyITAHulqThmsZeCd5u7Y2zhg
6n9pHtPO9yK1RTfRzzPEMdn94RS7+5BU1Bqer7irgm1mzTn2ntZwThpVXdT5eK8ghyxoSbxrr1w4
wKeXzYkKTnXzdxtNDPdJiMoQKLrwb90NJhiU8WO1QosgXi7Q7knXh7AoIRwEgRtbWTack03k2PLt
uX/EFlHFCDmOqeKAVZ9KbfetZ6X8qBYqnn4UsB5Q71qxx100gpqvDNdk541RwiFwZyJek0SZY9Rw
FXPLpEcaKjU7sm6mk9saZoblhXd7VSqgGvGqCizhGklXqlZJESCnXBZWdmttzYiasDro5abE4lzj
k5AHm7xQRmrGkC10HFFCyIiGdlcfCK7ZtBFkc5uKk1usexmc0C7W77B8fAxMirQzTGbCwcJzYacj
RPFtKS72CYcmgO1dIJUwd/h8cq04uQwT51hKU9lZii286zkrc+U4Y7BKDIWHZ56tEOs9fQXPY9W+
oSfv6iNQSzOVcoCOTbMpArqpqIu5FIKx9PmH+oa1tXswnzeL/RokYC2BoMKRKquFH4S+5EHTuPei
HGJRfajTwGBbLzFwLQ7a0QfabaunsdSbSjs/rYt9TKEYt4fs6DnuuA90SB+BbjPttIjPPEy1MhEn
KugjfAhu8abpPlLqi7GiC3RdeIP2WIUEi4CepILF/dsDumBv7KPhSWIsfGWuutF3BD80bk7EtYbz
PN5truUAFVPmyjHlab1t5Y/AtHc9ZRUIVfar/FTwhVKWOjQqEhhRC7ruO+haJqUbwsBfActfNF2z
PuQ/SMD4fmSSUF7xAwZoVxm3axOC7qwz9xF8SUzIIoDZpG/FcIHS5coxvxm6N1ohopLOGSwtilET
Ji5nECbv71WkWqLFqZsBDMfSX/4vz6EunfXuycGJilS5pwkGE513wymSHgH6DfnwMcHAdSwD0a2P
Lz1bhklrfKb/Derke832Z/S54srERsGQcRsS5QbTJMrL+Je8pRgX9k4D188R/EoOGvts0PAqtG3c
q2HxVNwbtngkdO6lDkWeTuaHFE9Ut1uAZaFIlvrtI808rDVcp1TDiFS7MsiNrpDqQtxsuC116/BY
FXDCDo3p8tMnWfreO+9Vlu6rNsBGkwWQMzTu/lwRNemOcGfePXhCOynNv5mPlq8QVhecDJXf8c3d
OfVsDleEDdPRF/JtV/yblryG1gCMtAYzbgTvi7q1kE4CErkzvHOUI5/qAJNtWlihdL2zyGcwXocm
D9a7ozdR+e3FPpPWHYXAIe9SVVgBAyNpQmc1uX6ClpFsEpyRfxpL+Q19PY6mritqbvEOTt9KbkHi
dKjWmZCbCZ6KRwMRvy7iHWu57RGl2mR7Hi+tzQFYCRTEeb01uHPQY1YeKPiEFM+WQzaNvwPqtTDT
PYulTuO1r6Rco8Cu0JDU6qpr7RfzPIcy9cjyEIs8MYxdeOtCGGuh/Le3eCPIeqcGbHs693OM+e3C
u1OxoRIMmAnBKwyUNEVo6YMmiX2QtMatFHjsYr/ib3qLrzm45n6dyk5IM/TsPWLl6PPnXlysx/oW
xhB+nkV1diT2Kt8MqII5L84xLbT7h5ztrXp1toC0gf1KMEAIKlqOjN1UPA8IY5y1JIetFf9J9Jq3
EhAe7ldvRCAs5sfrF6QkDCaZbhVOGnaw64ep0OHzILJN0XTETlber0U839a2S+Bbz12mMmOSlt2m
RafkYnh3RyntwWL2dC9N1WR/GwnNv+L+3+xoBKKGTVAbOmHPkS3NKqSt62vNmD2OU0zqCM2wQqWY
sYcOvsKdZTFwPro0OvN4yGYWOCV6cypal1mF0JmJWuVlbqT2EryE4NCNNsONuEIgokse+2DzfdY7
t6pJcwhm6d0ITtKA4VozZiZUy8tZKtBJNJggzUY/LRQYX1TEnJ5xWODbXvMlPHGEzyF6VJM2m9L6
7kI20Lsu+eXiFdiJJpRwtWunamas3h1WgBcpUSBwluBWwlyXNmup/UVdoHrNs6IJkQksLBq920J6
Hyva0/a3uH38gJGbEhbY4Bysmj2p+VGeHMQ0iF47SdZySvvYB9QWzbDUmL43EWRjc2T3HQWeyEWO
ETOMYMeA+95pexpPOPySFsuH93vhm6ROXptXjmmyGpcKljuNi+OJyaVggaOGZK5JA3TWnivOnqz5
z/ONqWf7wUsjV3WJ+x8jJPVPXXbop2WVSWOCxraXW5Gm/3lWRypHW7G90Leh0KXAG9y9Fa7gJmWw
tirDq9aHvvIr94VfxthP6XxADPR0LIRp4UMNPyVwIz3XHCmIAqnN69PXuXiu5BvSMrZzZIQxvtMn
JR0VThTfvqbK1dTY90w98s5Apiu7SH9Rd11wwLIpO8zHKG942z0Ksu6bmKKA40dR99xg3jszTDXx
KA6iGPX6vDz1Pb6hJoN1qf/sDvaoA9EpH3AzsQ3/lVD8OPBYMfAYSrtZb7bH28nfMpjKSGgmbBif
f/xzStJLblhfJQawD9SiQrncYiCWKf4u63J5eIrTEA7NUIWGrx1viyFXSKowo7Bp5Tto6LVcPdk+
bXcrwF4ZwByUstHFCrVy9XBdyQGwM4QUvBxTqT8VVk264tljJC4Bu03r/1TdOMov6grWgdFviHrf
f1MaW3n/uEyVHZv/OeqBRTIJot+zhE36KV2Dqc5KFeWYJdhRF3qKRlekxHzf30SQHfcYcqP6VfNl
nVWJlHe3lmfFhNQn83LeVNvBJdx/4vSYoxi0cCRvTTnf0iJfv5NtC2o2cF6TbmAGXgRkNVaumDWv
7bbybPYUs8L6vN/eueKkiqNCGQwdStVZbWrTsuRT9pz9yyTRVcLEKD8+3Nu6FV+Y7wYeJVuv/hoS
KAHBxyAYifWzQcOutuw41of2BI99/usKd9+ewrgcwXpJUD1JgBLS6hSreHZb208JvjsGXD8weWzr
FimubL2VnX9QN9058AGQHJM0AJ26FBUptMBgX2Y047Tlw0lW34UWd+ERuXG3I+oCYTixHu0HQiji
JFlmw9Ibrnl616mMxECrRu4ZeIQaZ0G81kypxQfgPIcn5aEB9WmFEUn4VkIQ4e1V2LBxZMKxpnTj
sEyEAc5XB8oSlgX3FWHxKbZmsYpGaD9DkJ5h0jZfcmXIz0qUQZ9IM4483sC+8GYQkeQAB0ickl+T
F5exaqwQ9fpHhXAvcFP5zNis+vyHyDtCiVU6Mc3is6c8fFBTfNrZ7WYPuGQVaj5AEtAS0NrLtMNQ
TwGcLS89rU2/AlSwtyIQW0z/xISpK1fziJhMjPIvPExuBWH8pQC7grQo9jyAneVHGRVTsiVYR8Nb
//26iQIBMM8nCkxxCwzRoQdRibaDQdwgXo1JG/EB32Jv70f8E1a+ABUAXBpdXG1UFFwXthh/Itq4
87QDMOg0OxWVTpuuwOj1kRqiZJPewN+JmS1nfDqJeAR8KncnGw43zzEyXuPa997F7MiugNNg9MzW
+2SGHAQ1E0lNr2H2ayFzifrkht8kT1JSacPU53BbN4u1jaQCXW4p5ymWEibihkROyNk2Eui/Z4gE
vDWzjmB3ihu7At8PvyotsNvD7lN9REdvFjcsunNRv1nvGXGN2XHTvVWFYcjGGK3k9r9fKvCz8qZp
KSoHARKzqvhu0TLYgcI6CIG8f8xN/HxxLJQ2l2LUKRnhBZnx+KKAJDE8quq25IuPXaXOYZNdSgnl
ShmPnEh6K0RaekX2IF6zAwQsvl9PXG28EEFj1ywrE9HSSiSrWDOjzjRhZotqczyQyOuYuWinioBr
8g14bTHRwTlycAUnN8fk2mOP0FSj//012mU398q9TWaxXhFYWVDLWvg45bwSy4L6V88fPnBBF63r
gH2LnKkOsxWYm4aiNZ1CdgezSD2k3v8HyRMQ82xv3XFYoRteHy7BplLcsQIAr7qj4l2gViH9cIhu
R78ZqFRZL7mTddyJIuhgmlGf1gR6fUmo/mq0e4pYAPNByUB0XoYPiP30z1czd/nl+K5ABgkND/ma
OC1kZJ4MaBHZS/UfHSXCp8LZC7NYZKMoxf84eZ1SSAXzIBSor6OzDiWE8Pv/63zU8DHdWmdsT+Dm
p87ulfGqJQKK/6zWdREeJaXVsqSX0b3SRFajoLcxWTM+DP6xYeIIGrBqR5A9DlbunCTu/Jy+zrLn
sWUICCZXYmaDbMJr+bfnMMHDoCvhyzlfehoVMIt6IE4ttJSlErzmbQMV1snFpvwwpgoFQg43MYaP
yvYqer5AcrdoYGDbO4YAiTuo5BTi7ELOHqTv4g3J2GsEy0TabDs7bsf6Fb05jEIylYmn/HIIbWSY
YrhgLCNZmQYYrrUjLDhlfAOkhEu5C9JAEJbsw++MwFWy5AiJToImAuHDJGD5lnoYv2wDlbsJYlnV
j7SQTVTFhgFECzNdXiKyYTj2OABim4x1WonD2iBvwjXwUIX6Crnt0g8pCBut7r4JGcSs01wS18P6
mo9SbDorHe96eZQHPSPNqzS7Wc4ZN3mTAEGjpA89pr/ayO9R0GaLfBEG9dOiUHZgOGWiIwgyIn7/
BcFBSqz2kbn41+YybGNAmKNixdSaha5E+tsbQgHyKI1N/puFWvNr88ATjobti1vk3YMTg2i6MjFA
T8lgVPSCqRw1nL0+V/FS5YHwZgA7vGaVgALlrURdQFxlsS33CsoMkmk5cMGm/9c5pE8Sdv+VzXEw
zy1VF3f34VxdjPS4DT10AFuNcVac6F79oLzN2By6zK8syGuNSIXZU4LNYK48zByPsGGIGC4Jdq9j
rpSuZ+7990JTPD0oIZJaGs78gTc6pcM6//8WgWVu9IFWj4n8BqSyaJE1EnjgIVNSVMz3T2KWDGKK
83dYhx8FjdkRZdtbQd3rUl5d1chCH/Q2GT+Jn7WOszQk4cvsg2BkvhI1jWt7oi69OHt7LLP6m4tb
JZXWlIspLu8KZ9fRhM7g6ElNwL8F5+UWbIVz/WMZsJF+Ai/45oajKsBwsrBOEcQk2uWTf4lHGnUo
dDqZdEIooW28XVyuVuyQqsAgur6Nb/jN2YVhU5JQ9aXOwdMqAf3eemRMG0oGgnGvySUPsIkkynP0
bgbCJy/olEQrGY7XfUPzspR20rVWgzmpwcNR8VvcY4gXvgF3UHiHtcE2tWSgxB6Wv+0B+T598/qS
UpHqbhdVGUH9gTEECZ9xcVqg7RIsB31TdNjt1v/QPKdRsei9ovOI0r0hAqk68LZCs7zHNz4GXlAT
5n1sYY0G+SBGVP2bwlDorj9R8KCWzqCKyY4tUJZnskK1UbXZ1ttylsctjhUv++bPKuC/fM+2Qlcm
0D2PwBaoCzMebJh6h8ihMKIz5YfbuRdDeekmGQv7raKLVkgblLhzBAUBTJufyxFwiXYSW2C0aCBv
F+rY837rXARZ5oTnZt5/CaSG3YQ1evYX7TkfzooaqAT1sn9SXA1tY2gyJHhpDzOYCJXYe72P3K4W
WY+amtT7GcWI1k9iGk7oUZRxvY8GQygNjQZ23fcBG7S/QysScLgFVq89uTU64tRNn0fzc4f2NO/1
TwoAKX1AhAraHxpjZ1vduEtLP2Y7GcJIAsL527i6irANJpMJPv3G73hxkhcFL6ZGU8fmnUiu7L80
RaqE28Ecf3q0gZgyjihpmkRJgzB1aJw62XDykHSZh89KQEmkZ8LnamsfhoVqvRmOi+T/MK16sEbQ
774ye3Y/fyXu//TpO3ZsUJp06UsqDu1+RxXXPC6EfwIZj8cmvOP5O8xbfNOvmjPA2ui4USk6Di2C
/V5VZPB9kq0ECooEWGv0xB4nd1hdVQO5dxbg+RDWMAGWq7jKG+xFAICz+97sw17l36Mn1tyILDU6
Y5k/ROQCFQJLo1zKVi0flneWEAeKwPoTMlF1aFZe2nAmofFTGKBHCrBqjOkiGyyTJ73WCDgsWEGs
AeDrCkLp2trDE0YtXD0rjJrmHCQKTpzu7gii1OVgzGjy4xUdAOsRscuGVmVc/sdzNuzgyHJ76ELk
ma7kpAcXjA5/9cASEWeWUXX70tMbQPvHsEFb4z9Il50q13ob8QcJNGkqXfgFcRKieIgxjOO2y5dR
lw+Obv8yX1LEIWkI/3e52LxldAsFYP5dEl7dzK6Nv5Zdpj+9mYy21m6B9QyvKjxin//zMoPwk/ZU
lWJcUeumC4mh4gzdrPvIrSa5q6MVmEljw0R5QfVln0q6J/XcNSISkWqIa5d34WJAuCAoJ2ycPTgp
hgpGZ7Tc4jHNyWxkDiz+nwvMlFFdbWj5xQKMl+1pmC2GzmAfIZub0HGkkEpdirGAL9TJADAkELq6
tpT7G6Mn6gPO6QdmZbOx5yY8fFV5UkDMBHXRbzuc1TZ6Fsq4YiuWPkHvrx92B7R3Uo8yUEI9OFq5
xhxmQcDZpLzON9zYHBL7oLbwNoRhUU2VKjknx0YJ+1E4Zifm2WRVQmrj6ZnpuP3wXTWMYJtAjCYu
96qd1sSscT+26EPYmDscypLIN2qTELkqh7n1ckfTpLeHxW1Gcc29zFoNU90RHMzRAoaoLC4i0gea
OfAyxEbD/RqSR7bdMoLy1+9fqFhJtMO2lGtQ9xLS2Wclt+0kli7Z62t4Qk8lfs5BMcnWH8kf2cxr
QGxZS4Saw3U33irthbN5LkA0b3NipMDhF8K6Ok5tRtTQDLxRQZxUepzcmCFLHa31a7vgjo51xjhR
w2+CPTzz/2MNt87dm6kAGJ2CRWBARwXa9HCcwYo4/ZkPeqVdlv9kwjtQorQJCT6D0hGBRweJS3Xt
aJiuy5j1jZBBexuY0XirXWRty7TPw44zUw95STJOYczfCcsHwFY0La/cuFhPbRd2EifehaMdFuqe
XcLCYiitmY/YQuxA1kGN5k5v7w02UI+wCvHOBlRr2jktWTtfYithP77nhlS6I3TitfWND41Bj0tR
+DaZFdDwVEipEUbBzbncaOa8T2KzxvTGB8JkRp7FBmHsKBspPi11HpWftWtpdh/frk+xl7sDLTOP
hrHg13b3SHB8ffGMLx0xlqw6Gr47+aZ+OsdSdkTxG14J/+uyHSd39lDQMBiIz6Jc0FFlDbvdzgH1
sBkzfI813zRimwS7hjtUkf4DAe9f6eDXB33E+5kdOkyqTMa72Vv7GpLXsjp9BMDYvLdQDFifvCQn
RWxJDCwiwDbA5SEP1CAop5WhKURggDLRAJLlWicJTmr2RoC8mSm3/5jz48VwiH2zbQXCxH+nspci
6gZIyZC2dGKTkiUzJ7hst0LP4YaMSLoH3mjevteUzDHBOgXVtYrLktZshQMnmfS8iDMQsYTzqnxc
x31LE296pOGA03kXlCoth2ToMTwHOsJA4+hwcugt7uxSICNhS4uOqA8yriFYNeMCcvzTPAbgDBBJ
J9GIrkZDTSkgTogOUH2kcPLeQn3W3Rbq4BTiUS7galCT4eLgIHNbMjwBkHcrtT9iVyHB8am7bvnL
Q/pNCNzpoOAXLWiEAaOfqeWfpI0B4lDXoZqvwWHLMwgS2+4UVTT2ykoVJi7tAONg0lupqu+M3nw7
dCpJrQmUI/rZDjE58LoPJPzhLjyI+DM0T9xJcssDggel4TU9EMg98ulMefuoSIpo6/5fwaqlTnx+
G4ogDfu9zH5JMXNoHWYOB4CKkWz5T3b6ksb3M/R6qpJvVm7Im9gQgA3op+Qy/KgHWq3GCU/ojTUK
bEN4MEsNcqmpwWV8Nqvv4jmk8349baovPcXOMwSURmhVd3VOM8D0QChph4Fqpx3Rb+DPB9b4Ohfy
/JkiMnMbHYtEVDhCHbltXmUiVufyRFNjUeBBG/vPvl56wdLY26S2rrjbm00wGOl6xemIdZFz0AFO
ac+tlGH2zdEI0yHEYi8Joy6ODhJbchDQWN64x280rVAWtOybKU8YJPwuN2Dm/Bf9dOUfgD0w7wOz
ttzKHYhAb1X0NcwhcCiAhFOh453hcq3uMcw4uyX7gk6znTM/TrmJlz6M2SlvH/nuDUkOKIOrp5B3
nYTDEw6bYbLzhy4cOcI8ah7icRmyP5Ps0sMTmzU7SFY3TixAzORKl0s+n1rUutBkbnUPJImilIpO
fklSAyTskT+xwNnMKe4wickpX1Z4hNAsxgSJGCu7mIxd9MJ+1auFPfMcu6BL08Hh4yzJZVTqnzSa
IQ/wNGVxRPLJyOiKu+5wfAa9/xQVFoseHyCFbC632O5xVu4rKPnIAC6Xk3pTolY5QGUiJRxVLMou
iyUOC9hrLvBGd5kSv131mNwOrBHmqQ6zqO/0Z9TxNmHK0bVNtV2LszAsFEVM5GabPMPsIY69Z25A
koG1sF+SB/rpkRPwwrQ9ElvcYv8O4deMhV8pblcrk/LwSGHsilF8FUV9nMdyd66o7iw1vJn3G/0+
ksJQkWLSrDNNdHRzdSm0xFy4YlO7aziMVXGJUdbKusPwK+0rPxmzTLJh8HMpotgCR3QW9jkfC9vS
yjatFCzrb7ujHZwJMHikkRefXLQvQtuXdUsiR+64WrNP9OQmQzNmuFwKOibF2jxyTQZUtqFjcGV9
qkZv23WllQcySCcxYG/Uz98RwtbwT1WbIM8Q93354mO5t/W99NJlK3oyzAEEV2Eq7fHBug2TCJpB
1STSSi1q40o0G6eD+abav2GeAyMYRxKyVbMBB1v9BrlaVnSVc94zXkGx8gmbD3yRwYxPelhl1T6B
vgio3+Q/hruyLCzjuSxClYZR9FYYKas423Tlx8XoJ/BH75u3tPbMyPaPO7tk5hU92F7WPTiAZRMw
W3DwvjEyF+CwJSrygKgoPIXblDY/CySWPBDtigJ9S2n89cyBJsn8VV4oPvjHqqZLxOmW843Dru0r
9s7CGjsOs/7txU9YOl1hCUE3YT1FECqDfkyxpudsDO/5EZWggZeLDVlMlPJxN+yV0YJjMQX0kYLR
VNDhh1HHfCKPZ4ekAnjh+bRrdtFkAINtUXH0e/0uWP+0l7KrnszfGo5JqEJQmIAQFcLwpRc5W5Yq
W7rWVJCCAZS7/Sbx5y0YJSogY3nopPqdbDgMrvTpdCqYVfU6nOQERep0W+hMwBwBlkbKimhIW6iO
LlyNcPk70IfpUDo6tcGSB6uO0dsf4wERxTg7IQaIZ7LsOw/LgazY6Z35mtLM6V4suxSO4031krPe
85gEh1Vhwsva3De2r+Rv0rYB08Nl4BDJs/lM/b7n1C9s2ZfOU+63Delj7hMYQfZW4rqAQb7kAc38
d+mUahYjKQEmpp2bNLa7jMNCy9gdsQI7/pOoTtSvVfQWCBBeQ37+PeG4x7Ob/4IvMyn3fXPdKLvf
Bp0QNt07OoAlQ6IpvKqsyHdg4ntGpS/MaJL7VfBnEelqEBwM5Tmvkb3vj4rExVhMJlIcKo2P3UZu
+a2LVKHvVSn0n7N1TopNxrTFgvrI2MKT1kh1VGidVH4BtqUvVEPHFBY7d7l/rKz8ei63bHg332Kh
l+T2H3lPm+b5u6JsoGNcl+b1adXT4nZGjHFlucQitGGVQpiZFKW7CHlA5TbACGHSj4oCTgcj7opM
MSKem5Yg8qTwpGXTFQF0h3v1nS/6OWsmBuvxFAW5EKbvGyrvs2WlbV9DPAYSeZt9mRuRkzqac44v
8qzF8/38+9dLAJtOV/+it18GGfrjyW6eKD8qioWCjuqgnuB0xRdhKciSDhPwPX/QXkb/UwS7/jmG
j/vb7f06FpKY1DjKDecDJ3ZxGTykHZ0La8l8jXedW1LJy5JzwUI0HxyayOGkfJDm/qF3SH7uK+pE
qoVBQ9IdCCJFM/ZdBFXsqKQ37MxPF91ekgDKgBywKMZr7qbqpduT/VlxR6K4U3/21JM1Om4aDMyn
S9lwYp4UWwMv37YxIdvdugGg/V1Uqcv/AYAuauOA+tu7ZDm8y+tMLTXFfE2zn/8J5eVVDLI9h6LP
wqKGPQ2bcYvNgjKi/qyCJT6DemkvuxBx2SeMeDLEMgtOYM3BAftMFJEQL9RKblqFqZfeYVK5Ll+L
TFUf7qWl9nAJIKvqwxQXEtBzHq3woXvJiIDNGnnHWsptaQYiHd26bPs1ykvnxsiMUHneOSC4FHb0
zzOCWwAcLmxqrm6STCyEV51w8zMl4OLwUrqaJWIb49eif3nv/05WXPoZl7V+3PxEJtkC41BBrLpx
aqb3rLXd0Ssd8RoHE7uYRSnH87Jl6XCoOaLV3cWx+ayY61P6Kw9NmEooyVtXy0HoVlLZt2iy9pwS
1VmTDFmFJn/wodu76+RwErmlc3vgtFO7JT9nFwVoTOIn6Gw37A4JHlgNUusskGJRt8QfITuZw8Pp
74hxrmZCO4DOuIfU2Ni5I2Jxb3U9n7pasy8eP+ST3ySzpAEE+Xzt8i7gs3qcmKV05DBKCBwGMF8g
88NRs62yIV7l/qXgr1fGY7rfOMho+5UqhiGclsMpSzKUK8E6CuSjagFtXJkbOnNprSxNt288pFad
B7ZyHCVp+bI2yTDK7/n73mSWrQm4a+RZZ09Xv6iq3+JeDjUtxBXfK3E03T2S3Y8KCBR7FwibXj0x
61bg5/X7FdZKWCSam2W1gLk5UkWf4ofLJYPOcRVqaND3Upc6POw8ziSVM6IQQ9XvEQVpb7J4/1hD
tpTKI1jlJv3F3CHaGsxiNxny1kmP3zNXMnhRfiaZHQtm1BfHNCMn59JG0p3MT8F/EQ27lEZdXIrz
OI7u2Dicz9ZnQaWouG6TK8rlxWcEGo/UPzM1SSBgZz1Q07IQD0QtaDMqky1bcSghoYftOEnnnHrz
zb+IofKZA4S+phiKDAK69x4Tp4NgHOkGiQsB8TbFJXVkQYPIUJS29bd1bem0AkJKBjj1rR+4V6Rx
OoGl6LOJbw2/nBiCOBE+sZ62R4fNUxdUFNNYbwaUgf+Q/v1C0swDQwEI1UpzbTiCdT03JdgjfFzQ
R8D9b/Y+7zpIZVmoA5EJbIztgbVqnvXSLGFgHsKt7rEm6/34ryP3KqH42wAuU9P4VqEDj8A0oZ/F
u91GmbanJEK13lkhQjD5FlyufbBBc5747VzEHbcdHkSdR1iTjJBqSjk7SeSmrX98XMsr4gVsgUlL
DgamyHOS7a83sgQSkRGq1ly6D6cs1cTyx+owAGMP26FHaBzX1IhJ+iu/K1Pu4BenLKLuDcNWsA0j
c469/xiZB3QEUVtAfx7rldvjtmCqEb4R3/8vybGi2jRnLJCtWRGeDDhQM7FMgxSDYRDIgvbzH+AQ
CUQCeao32edIS6ASHQQs9sdZOp3OkwPMAKLxijeIjXyLuCxT8zcXFKhz4T3wC5dFhOeV0MnPei3U
b7oegzUKxBztn5Kh7VMzjxDfqLky58Fizb40c6rRnXv5t95ZfJmHTUWr1fXhhexLsbPJXEOwvMBO
zRhn2nq6hEN4aApflyaSkOG7eY1OO+wbb776NZ/DN85wHbhwwOR2E1A66+QdCsD6yGzpH98xTJad
4QmhqdoOnYJda51+I0fGkDie+u7rn+tspX8kKmRh9IL9k7zcINz4r6CRfp7CXi1K027X05narVQz
fpCAZvI5nR2BDi4s2wxfeL/pQ9SEXZGNtp4ZkGscEpPe6PQ1akxZRcQimR18UZrk2FP/Ed6pWZHa
2UmPhwtsGiPEviA6YH9v5cSXRcObS513WIzulKpru0oK76Zpna/yGKBQbuCKLcFAizL5dvV/lRF6
476hOouAPQNQZ9WUaPHW6h3sY7IkjcchiM80RsyF2PZlhHvfon4zCx07+opHW9tGlBtvKW7DEoxW
ET7cnhjlL/Pgye0cUSWyGrzotUpaO6WAbcie9703rtPMWfVfzjsQvpGjShyE1xsHThAD023rMwT5
DfHnJ3Q9luGH8nxcr2pePZvWc8uiWg2BmqPpDS6fqWxgNCXWSWRgmnM1WRM9iRnSdclREA4waFy6
H68UwebbkvV1/2cT++r+bwhJ1tkvKtzyYLKqt3UpLcxHrkyOERs5Xnhe/M/9u7ZAoVNnmDhOe9RR
IXopPQpwCyGV/ga5HlScqsje1XOvSkvsvESd0pzFH0czJH7Mxig8xK0H3H6JQq1Ab8XY5AVXAFGQ
5LA2fDMC5Jw6BLZ4ghMUvw2XjH9OazD+tbsZWEH3bbzjk3zHB33rcDURKvG4wYi549xPOo8S3Pnt
ZokcaLb4eg8vn6owMa4NdZSp6v92uueEDS27bdIP+8a0djWapkbbawjpoGzZfRVsRHqIoFIB/Ify
YLXit+WCFMpXGjdv69VM8FzGIvjZYDcyKCUJjEq9sVuzT219peP+NtToXGSpQrhClEserPbaHtyZ
XClNGZIs50+QmYDbggZALEKbCu0p+6gw9fHmiJZdvTIXpVdKsEkCRhIBAc6RDB1x8n0QBjh/qbce
Y4+iE5DnPY3zsviOBuuwQusLxGz0CRTbdwk4MoHjOFZhaIpzw1y+4ZFPa9Io4DQjWK014+giSRNn
Yaz1aD1o7C7axyhALfDmOZqVdxg2RQ2GmVci3ZKiVQjyQp/sv8amY4u6JKFNrfdrzpWeZQrcOrGT
Y1Lcblplr3YKWncIMSCoTz4BGMfvYkS+qVxcs6eUWv8iVRzYC8KGAwzpgB49HT8I2UtEVpmWNEPU
91TcFcOMe1eDMiKaTnTETOfsGVJE3zloihxzewlaqjbfrCCjs7EDXKwc31aWfXAs3cQ50qXg1QPU
hydiRjZBSLbcIRSwh7NyQGkrexh5c7/Ew1+X2BNeJaXh9giFtmSrQdUjb5scdT6FglnSF402h5o+
j4q2iI4LIYoQ+f3bdn1X6dmOT82C8PBrNIqwt/9fp9csn9YLChHtaosaisnDF5AXOBfnC50WZMol
K3YubrZvOYZCJ63treK3RENs97dW8Fk65zhEn0PbnITE1K9MasDamdYZ2KWcoT9diP+ZMXTE32YA
vou+uOF6id6nHxo1UkiElfIM6HLJgzNhZoabrlfqN9MomE5YHcpo0II/TAenSWCm4z92B7JG4bt5
/mB9+pBJWq+F3eHTkAO0tfLl29j9VZVrZcYtYfrD8B6QJ5n4Abxjkjf8IzGQwD6xXjJz5pYNp00V
/DicTH00VMwjlcZNrqCBGjAgqnhxhUiK7Bvg8lPeTtts+ngbJh2kIGtcx/RWTXVyO4bO6MdxEWuC
sKjbFDHG5H8UuenOLK3GudOum5oKO6xHURqvcw0YhqTbf3FgXnGyB7kVuAxl/HD5A5OTcVT+hzhl
fchjmfLdH9HrKRgXIAUe3P3mw9e1AJwDYakQIfMUVgS5vZFjOMQufpGQia9E5q0kHEE82ZBPaO0k
9Rij1cAPJQKQIVcuOYXyFP3ZUJORqugQYPAZc56921OfhyFnWUC8wlAWZhfmmfqviGyc+0d5xMKq
NxizvDsq77b9TJdMMRT0QVgaVqqUqeT/79ozO1+SdqRrq3MvRId4IzL5ln0f71Zrom+g4OCM9sKc
1UqMVsofzBvGTkjlUn8aEnngZTY2kQbeoCmw4sjm2gZLFdYoNFW+msb3yXLhMp+i0GCElcENEy5a
TdCk2SkjulWZG4UV85f8APtswXMXXRMNWXi2ruY7oAuHwlifM1jSS5jpI92IVvdFPPUzAGC0bwUV
MIMM2WcEhv8zQA3/sxnPozubhRNcQ/vAr8LXSuQfBxXzIBpOD0jFD5m20AEBSw1tt/CkfQ6iwlV8
/9+VqfOqJYOF9kaEbe/Zc8Z2NuCnWcS5NYRA/xlUim0YPZv06mG+aLZeYhv2g6s/RS2ap3u8g1u0
Lm5v6WV2vAX6HGgR7IO/Y46fr/5NaJgl4p8+1WmbC6wMXbgHTlvtqii4bvYFCssPNK7XsCJO7bY8
Jwjf/+TWoRrmdApBTwlqtdhniuPHuqdiJqyxnqjfHTqRs+e06dzRBHJN0RPzaMDk0NPQVDSUshtV
sVmqcKWDOLdaUtOSSrJ4nK2pvAk3YNSN+J77IpKbu0d5w21jUO5TNlOmtB4iQNpolxh9a4sFBVDI
9kh0l45YwJW1hhp2lqXGGNN6XNAbIYwFVctJJd4vJjUjseEWbJLH8uONHPvljRBWfrdNRfoXAj8l
rlWnVGBM56azYwJMh1Ao8Gb2A6xHxMsbsploJYbFlv+UI94myST0Ve+CPtfXSclJf9KwXCIkaepY
HsqXEUKjdCHh16Pco9FFdOqAoN4mKa2NmvHyLtgBEjFwusDHP+5rP6/hZ9Kgw6vYYDdOkzvMAslQ
89wGKQyf4gBZLctmEmu4ELmFY9DN3Lksy95KmgtFkmR0SsV2U6LuHlVhvgCghZiUzBZmrUWA+Kvr
DRmGQWQjv4kWattwrFR3/ighW7u52EhaMRmZA8pvHK2i7Pya2RsORSh5OukEYZ5Q3ad0ibjlXV1Q
cWIV1qhEkmzHVQOzXjEGSnTdEgcLnSSfHpnAU5r2/UbrjGaJa0Cb8jl1dnLjTuhdA+LHsWKmQAxz
oPYqpapKfBsP/02fHrb0Fw1Qwpkz/IdWz3XV3jkps7s2bnOV+bd/pne98GK10l/+MKoUd/4Hw1S8
PKinkDCLDKpn5CH1hsdwrwq4IDpFuIBvWtkBRRWpwZN0c8YpTzfuWLltEwQiWzUnpKKn6g5bNI9Q
YI2ZX2JM+Fw9InpeTM7tMaUDWhE+ZW90l3uCfGHFnRSbJfALBFVPMM+I6TMJPP9Uh1W1KfwPfKqv
dBX4RECoMxcunGI82WMLVrxnxYmM6mcROHM20uL2lFM08QTjTZMbhGhA9qOSvRj7kH/Kc5AG5EMT
soldPJfJLQ7qRnMtw/2iIT62+T7DxGtP/NGJlcCLSdrJ9OUUgawyFCCOa2o1YfnMiv4QvVpo0y5C
OcapDU1ePR3VCKVvtTuOs/APIuxWDjN87OA6AeoVKWjWzXNyPh/YvM0wnSCAXz1dOqfwf9K4KJQf
lMTLRlnggGlOBOI6TcgywuHj/NDWFh0KdYjOocGRn6RdeV2xgIXnvZnhM/2a9Pxqe3MSfRC4P8V7
VwpxDW2XVoa0pleEJF+5JrkTSpwud87BUUla9d/6ZqHQlTvxjldH4I+wMBkfTAzGsA66HhdSC4cJ
EFFB4ToMmYVOaskj2s/v/qSa+L3GjZ+JcPTPjFRnNETDjvmBaODjulqu5vxy4b2ZzEN/2A61GrGz
QbotfmWIjWYC4ZfYzmYYZRhx2tZxc7JD4OF4VxvYuYzM/G2zr4mu7yguh2oZNfq1mgb0f9uSrh6T
5Ph8pP2qFqggsiaijdE3uVPHNphZ3O0OcHreA2mjZUgRSG2XEKXfn3JUbfRmjPExvVtWgR6+uxlT
s2InKeMmFE8OfYWfS5cHreL9MNY4h7iTsMqSqlk4twWHn/5ATVAPcxTzpVn4s5t0fgeEBsrKIQj8
sNGtuuzmkJG2oQirhcuh4C8kx/AuO0MuRA8SKW7jCUoBAW5Yy9PsZ5fK32Cm99oGtqbTQIpmpg4j
qmTDdXIwLvHJMDQxW48i4zJv4VJ+/uyrlOQK4R+TT/zHBVSw9RrJ+MR+K9VRoEgcvRdWp/zFc3xD
thnoOaGuQZ5fWlqeA4z/wMnYJnNEob15la0n/fyGx/gq7G0KoH/tfQPsqJ6UATyRgFZjPazv6L9e
JjCz6TB7KFiiVwfxwB8F8Sxwqr/6OgX9g9N93UUOI2d63MLYRMoK8YngUldV4rqq6H6QlZDoHqYx
gmtM18XXa9/xGPyFMYmDrSJjm/B5YYxMNICCqxjq6Zg/mQV27a9pFD6mRP1IPhMIzWNqqtgSZBr2
SAaYuXsCx2fQdGA4zaM3IBj2nTxHNWaIK+J60KPutT29tCvSYz2VwJN6tr2ThKGdiNaCGVDOFvUq
mOVMbEbFqqsCQ/E5Bg+XmF2GR3F0EODEp28WYwne5JozBKTNCa8VLLailHx2U6oFX96/HEK5WzrB
0SMtgO99i5KVO0yDnvlkXgk1Wd0diAVDMgPlJ9+qUrZIJqGHJrRsCiP7nwdKGrNA4LHvbnZgpfpS
5ARcqHEUrvdw6WsXZ/7+w7mCI9aidUs2Gq7ZlU+XCd7JRb862tBcMEidPCKCPz1EXj9y84JVzE2L
prkZosH/VDpt8mI6Kf++2LSvi3+wxnVH0QtCFjZs4HAgCX+uAfBaitlztGH8pJENfEGSENTIKF8+
H2fBSmzbYDCyrP2K05bRSMksu94G52cmYkOiWB375J3OLKEMc9XbF9tfyPrf3qxwM7SIkleki/cZ
kLEhSVd4hUI4Mw1wrQW1WoZZFwAdgdMuqIFIY3+jGoEjCn5oxcmrGoxgx/VHaeY269PyOfl4kg9b
ChnuklsB5f4CiT7ChdQ3EqqorckWPINg8TaxQLW9o0BU0z0Cocs56vFstUZUq0A3YKjefxWvrIkG
yK8jqTKvpcO5JqW1m54zH3L1TmyLmuRIT/9z6Qwk2m8SdlNdzc92zfw7+KBE/TN+7ZEwKQtFmYLc
mU24kd63d4xh/c5n9YZXkct82tAslj7eVPL0VgePlefjK+5f0NhRVn9B4FI3JzBDlB32jGQaM2QL
9hRXa8DqhTz6q7DmBTwGLCEL0RE74I64Dw5nGXs8uOrJEdCQPE6TGRSdXSBSMnHVSZkLvKlmhSvb
VysJoPotCkHs0627FYHHLLlrONl/vsrWiUdNQa5MUuIVY9aikN778Pqq/v4PIMsNIPeHcb3APZYJ
l6RQjPaeOEZqZ1zVTaX0SlDv/3+bdJ/VyfL9of3dc47KhuKBgIcJM6PSYLGoT2Kw2oKCQssXwVR8
y2+1quVVmphhnDonlo+MEU1ek/sykhItu8UzlhQ9ysO5ngu1qcqaDdRV1rGIcbr1fKqWr3W+AOTB
LHX+FsvoGCvizsZ0ttPGuMkUvVePFc/AwopJPlR/G9X344GWUU4xZRqTycnn4Esl9YZMhjfMqkVQ
NQMx3XBTJ3Cx2XZ0upUQW2yRJJUfRrUYHpSMRggXjUs6ceiZ0awS10KSFxFfwOuQ3CkbGAb3Kjby
5eG8HiXF0X8b1YRQgh791VoVnRklQBDsy75ZNfeDbr8hhBd/9dC2CuBLmiPhFccXnyegFFirS2nl
vLubT4BeuX4P+Ndyux3eyV902HQ68cWoQskmzmupgrFRMd8H6Cv74ZXaUvqSXpdVdvxaPLwoqTR6
qwREcLHaIuE37UnONa5b9Lm35NbI7RK+ITkxx0LDtHSh7/AtyCtsZKKV2lPAOUPYEthR2zpihZPN
ju2dfFqRHw2AkQ7pVzFyfx6DbczxX+/y661k9yCTJz8GFGAfVCuX7zV9GWuBVk61+I13lZJuP6S4
rcZhWOUPZzoVQh7WtbtMbO03HtO8u4r24O44+Mrq/lDBXy6fUcMMALpArhX0oQuE/KnMwIkQlS5V
q1pTPmze5qtCmQUFyC6ymBZZ/JICW2FRjU4stm7j3eNhiplW3KHw7slZius+GMS7zYWcdJ4tuHvE
zO+YgrcYBcGQR78w04Bsy961T+gYB/5vsn5loa4i1uI+VkHHcDB/WxnNcqYMs3KbfK+lJXN7UCwT
vV8D68PrxKaWm+V9Q8HnqFPLcCBVa/RvUjAWdRi5gCV43xCQpd78Zf8yu2lfBARsPj+TsdRw5Jgu
ObYDeDmHdhEXtIUCilgMZrqIAsOmyOxcf9lXqI3Xs0qN3fckSuh08BJh7dURxrEMIoc8iQ1ESc+c
CC0KbFwDC7iVAjCfM2hoAYlWjIYWkF0yXk7gOi9o7hj2GiOq1AZ8nMvUGPSkrEQzdIv6jR+NpbnC
ByJr3SVmiKCgtVcCdn5oH7Xy9RNl3x19hHnwDVvggoDQnj6ASrDv78NvPLx4fQVaeAYuQsffI3o4
Zdxwwhi8sP6ujOz5Gk0y2t9xHTmM3i0TFcba3j7Dkld8vKW2RGdkpTY9VgFqhart2W1pWo+3MJdP
rBd80fVkFzbE0wfrnZek5isrtd/KEI4YMA3Wl9BZy7AYVBkd1aZe+M4jgThC/T2V1cZpAeqTshq6
EKlmrqwKUWu0TgPmiYWtJyRLkzPjRIxDhQMAM4sJBC3OzMQORZTgD4Et1vRkt4SqCns2F17WHuZE
0GaMOvbzLddXB45TOjk3EwH1kmlX+0gOemgJ25pw0MdJ8thgEXnJUUNf78BPaRCEYwFPp2Yw004R
tJVBJ3ZEv7PIXZU6armEW5fdYGhBbWGQyZas+r/CsYlDx7fJWYC+b+3NtEovnDDWfTy5dwA5RILn
Uj1tqlytNKzdQ+v5sZv+UsNLmdY085HG7tNULmShM/xrgzDAB/fBHa7rGSjIueXSN9iuAk8LRUW4
qB0Fh0SVziQcvolYwJJrR+4CATMutyxXcmC07m2pVSIDajkZzw1EyF7y8UkaliRt3UzvgY8CGyvD
SQUc9YAC+4UKGsVpIU9M8Ecj4cAJLWlaOHd7lyeKAm+xQWMy4uya8X04zOnBCPtQZg3rqddQ+/q8
VD8h4kalu57/ST2bFY4/i/WjST1NH/iCHX9WzaV7pDW8Vaeb4T3X10qiLhxanG3aqi9RIwCKJqix
7GXlMKtcaU2QYk43vBH/nZuDulLG6v6W2CTjhpgR9Cj9EbEb/hdQ2E0UCuGqo/Iu13GT1PPtpSoe
jRXV17kaMyUH3KltDmrLVYURWleblkIdl3lJd7M4eMwcHQ0hXVAcsjGxmUrgaWjEW7NLfLpZWNT1
5/CjU7GLv1U9D8V5QOOagEmRQxuxo3EEoSSlSJCw6OjnGjZFHgc8/kMnKbZkz8jrsm6LNYSv15vy
zvNofyTOMQIYe58/kABHZGKlolFpoJyPl0A/qFeMs18OvceGpLIQmA5056GZ48bi/vvp0p5NMhwU
Dwe2WcJrJO5wbTZePDnLxa9YLduhhMMkPVFo6q/BhP+x4MXf19tuJ/oHtYfD4xMeiukYdRBp6wb4
ScjK5EQPtOkZ05/19PoYcwBxwtc9v+S3DxeBk7SYviGaXfZMCWSqEMwzAXvvvaMZ6jYhvGKRIUeb
+lYNgMwKWUUoy3VBrV5AlvNdJD2FrF2aiZL1y8Tj0N7kOC5w5qy2YzMTuCFe9zQL6szp4H4hkMPf
sIGlowVGshDqexjPyoSrDemLQSSLzBsaU1GR5fFUo/qhLQbMWWAwRePTpMK++toI892H03yLpTr2
A7CLY/xHspgVUz4IXNlr1BDevcYiOdx+luAk1+T1v5zrWENX9+EK0c45aPdJbPeQb/w4VfzBo18r
jyEW0r1qji++JCmBctFPM9sXHB8dhqfd0Il8uOV6h2iTpZvND79UHQso7+IvUggOVjjgce3HAKsF
hnnT2fz4eoNe9E6e5YYkYPI71vNPtv7l1zM/g1D3V50pBjQ+1JlWBugZgQb88Md5KgNDN1e5RNsJ
CfYeoug6R8I4w0ifdg2bEi3AVo24fhKdFIrBXC1zEB5+9ez71G55DVcDw0MT3KxjRqUsHhb7a1AA
hGyJ40/PkqNA4u/dN7w/hwAgxEEtwbXjCsD8snHVzklBMWfduuYbzVzMl95+iKCPDeOVt86nyw9G
Bg0IA36rc/O/rWHoRxcjUzxv69WcHlv0whIgG9NM6eYUQYS6JuHLKM24Qn6yM3skDTpp0BZTBgUM
r1Euoa+5bL1iwmnNqjAltbRZ9gGjqABxrFRvfpW24jPTOYotC3SMJUI89XbNKLIF9zlRuea9QB9u
esRjiYvRKeDb5KykNOBzeL9JXej9bCfzkMsZkdFYFcSnyqv2+lA5byTlsupYlfBtdAVtIV7o5ERi
HMUjMiyVLHltihSFGwlIXXNgjpk3xxR+GTBfmzBX9kz9Jf9m5Zn7LAul4hH0rH5caSi+Cg5p99/1
JR6qaaOQSCwYWTIXAb/QYqapXuuaAdwwc0CmhusG+Cb2qinSF2V0LpYABOoEP94/1+9goSZhhPvg
Zgkt2pl5CgHYMOlr3WR4L5Us1AWdXbNYJ2c89Jt8VigtHtABfRo1LCxYq/Sbqh5AqqXuhC8uwHih
RIP3IlRJq2Lrzfm/RmUY46ClZikxs2ZWwGi2LvI9uQn6OU35QGEu7/2GCPM/pqsfMxk8oNvWCWTS
Ur2RQzadtG3l5jBh/QUIYlAXTD7j8RcsSmdhDiFKw7q0dOaXSI7Fyc7FomtL5mTzWkEpHLoSKlNG
JTIUbFDKls9Kzu6sVcVYsjktFn0JZjDGSSER2h2W9MR6IdfP38bhPeN8BbHM94T9+FfK6FkJRfz/
Eu94Q0HIKczS60EVozRq+R6MqF7D7A6Nq0FUH4ZCOZSt4gT1CePhn9uJvdY6YQMxJ9IRlytyMz4X
DvMpvdLvsQ/gVBg4DYZkf27kTjAVFqyD/2yIKBUcJDa9msEyo5Xd6CGe/rh4si9ovFViwy6v7xB3
2st2pnosuQWl6HI/VWDjxryrZInKgDDfKve2TDAeAhzJHH56FwaMuN6C1tiG/+OP5C33TLoskpTp
uQhfB7nTXls+C+nHZuUebwcHT3RaHc3DtfYh+kAwxiPVugIIOFZD/5hizlvMiJWUlwuqOKrqlseL
miTn6ieFsM08jYwJMMuVtdOxe2plePJGr9qnHL+K2RxIlEvr18d9te/YyDJ2silIbhPLoVrne52v
hpk2CEkPpPDkofLndFFelgkBg18IprLJvisxWYcfpWEwueC7LfmIKJwXJrbAzCHTagF7mso5E2kQ
/u7ppvZC6k3kgNbFps9GuJo79NLxA/w3jXseWyOPmqCIRb8f/n4yp26SHbKgCA4rkhMtc2Rc9AZs
owOTCbEddzELwubzHRPCT+gJbt1WNYv/UtpuXe2cRSi2JKRkCuoz8zW63GQ0cQrfzhQO3R9HFTts
pwKqJm28I5ITm/mUqz03NCmGi/PW6NYquu0iRMo2jOFGq/KJUWjeEe0aUJEWeT3SalGjgUaWKPVP
HZGUbUrontK9sqpSQ8rbVMRBYV1Ql5qaAEDs6A37f3XJDRnnTPIWw3k6x+FFvAJrhd4vhZb1CvFo
Nfdpqp175ExBzFXmCa6vjnz8VO7vHBhceMqv77W0poqBIIa95iHZlP6KQX2ZwkFDRLSzQG9T0E4f
SsoiIYKT6HIz/9PtUBQQbeAhPrKZYiuMPH+0joCEZXN5l1YOByC+pKY6iCCUOYWHyXysCUXxJ05Q
IFnH1FVibYD1eShTiW4/lDKvnWczUXtEeZhD7SFIEm8PWTkE8ClsFviMIMDiXh0c+RIJ+VLJhNtt
6JmWvpdU02xLOE6EkuCOWddPYy4YOmeRAaw9uGToo5wsTTEBtygNOCawQfjXGB5ICjnnCGyBClhl
SS3BuwHvdV/+4fWbR4GYaE3RQYzmC9VowWeWLGOFyeSm+PU3iX+O67J0IEmmRwKvLd+GWc7NRayq
xFs7rezz5AJmLcCejfl3M2NdSFWaIuvjJcLwgBIP05myR+ak6HFUIYRt7V9GmYZ/fjx/4MYg2iYu
w28RCvwAr3Kw4oqvznkF9MZtnqiR7kPSfdllvX45CMXIr8WO4oOPry5dY9bcv6IXj9p1SCIE/9sn
DemVWJws0RjnzwOTTmY2Klkc/Kw5keK7wYcXQazUcNHhyjaaSk98eniVb5GjG/TIrPna/dQAhFfh
EEOTvsTj9MbeQJmVVhjCG+znnWY1Jilb/Y6sAwprexUatbVmrWCGvJR1/dBlE106MNDDh0AHAHDQ
4DgaXgioKUhMugzMAiBx6Q2492MOU53sMWB2H3kzuCO2hRr1kyTBOIiT1KWQkhr9BgiN7pIpSbsj
v/MAmZE+EYzU7oLKixgp2VVLWELXP77EtPpNe7n4Tc5FbFL2HsEyEMenQNV4Z9aN0hCDHowPcJIb
FVKHY8ik6vGOWDdmDObBiDdXPewXxY2wNPANk2uD1MjS/7NzYmSLEhugyP/+lkgUksNgSu4vPvzH
wlE1uEwZvCqThn37W74ksCquOaqdE9rxjEk+5HQqheU2YNhgzn8mLomJooKQEmDCjFomz2kzWAqm
Vgn/3kxvcLOpYsNyrvt1nhL4w0rRlYjOvho5aUSVvcSacBOUFgSZKvapOyv+plU63DqfcpyVvn5v
CrSRudkhcAWxO9LzTk7rqiJh+zgyoSAUjU0OSo3fT++gfsvjYKE0C9RlS7TAB5qWufTAEIUiPzZN
vNt9pEl4YikBZ/wHE3xBsRtpGpOJFHDmX7yl5EKTXZPUapJuentGDNsWFtUSwUVUtoPNZXeSRXcf
0n8PNCVbLNF/EvwV3o0m/BXPe0cxthjW/RY5UO9BCczSpf0lACxgQe+UILIj9lb/avR2gksl0Ys1
Ap07+xprBKy2ulIG6XOJs72ymDVfZglzq860oXTi8yhnd7d6ETnQ60rWIL3+VYcKlJiH05aLDZQI
kDjQNXedji9Ijr6gKvJQlBZZtbj2duCIMRHVFUHuwK7jMfZZogChDeBg2ogKocB8pLRjcZzRp0s0
9eN+aUi/hyF0/Ia4dnZXgp1uj8R+4mlixEWZQhpN/XeGJ2omB+Ew6W8/Tdui84CKMKfbsnT6gDj2
r89wWyOor0Ea2XYHLr9NuEYxD2xqK57XNiL3vOel2J/ykHMMmEvc9n/i67m3AFy9N5oQt4LWEGZ3
wbVPHY1FHqH1zdHRZCzYRVz4aQ8Dugicc2I2wMHYRj6g/w+yUcpXIijQuJBSRfOV+91d7NwVHlgs
o+BQXhIR3renFcMNtj3TedUZ+39b+EgDDigTmbUInlxP31PVJjeArKCNjnqvk3rKuL/9eKIJZ26G
8mTLiuO61Kt8LzUm+yxuEtE6V+WA0yQ81ldE2UQ9q7zD5dK72BzZaOovBNNEkWKgeZbcEKmz60U2
DKg6c6G751fwJIA9TQIeuO+ZsgAg8z/wLfRIzQZvBA4xAKtZTDh1nxiiXCYF8au4NVYt84vYIThW
lrhw/AUGyXkrPezjg2POxps10qJGb8U9s4swwAfiSRIba6v65nX2wyP/x3n4viGZHQVfEXsvyVWi
cTT9IYghZyuGPI/+2c4rXtnPfD/RyswtHQQ0Nkn4MdnakQyXKpJhYeyLetiv8sZUxs8AJhbuyJ2l
0LGDYp6lFfUeJ7x6mUW/GOizXzIaBwN9lx0zjjJnbY+Pxmz/3uRWCyo31guk/Y2knMABwlmLgWhP
wnCg5u3H+Ev7sjwM9+wui0wQ7rXmt4W0zHdjWa23+IOIJG2CTkNfA89UxCLSiUzEtL5fd7ocaZw3
sDEj4U+rXPaXddn0hulfGUg1NQ8/bDpamZZe+x7TOGnAQYXBE+9jGL9mMuMB+FkUA8lt2sxOqOnz
6zXoieduVDJm922t2BAym949c0T7S3EcwsliBsPJDFmytktryJVhLk3FjmT+K+i9raKBr+4zEfVg
nAVtrFV4qwGk6LimkSEPaCozh6iPfJ2J2/oGB5NOH2qD1h8FLMZWoi7/dZslA2K7aSZY95H2uE3T
IamgC/ZE5r9IEBkhdUvTwPQQd7UXHU2AS3m142ZxvG3zQEybsATcxy6EvbY+sJ4cp9K9kBmPMuQT
F4/7WIePzMEv6jHRSbieFsMgs1RfxUyLRfxMOkf0A72qdHmKUIn3NUyZo3h9/jO8b9rKEON1b85R
FgcStwJOv84PKSkP7CL2wGnXLpc1kYqsQrBBNSfyVUdIq470ATUe1r71M6IqMqvp1uoz+1a6yYBM
G8bIFTdl+U9rcPDFyksMtyP9YXHDTRsWLC0hg5l9KsCqd5S+TrnF9FXjVD/wf3n9ElKKSusLfowY
fIcxMMiyJClbAzirvK88MQLtBz8p4ct+EHyzPKL3XQdnxjyVwhlgnps21WIVpC17Eylytu7SjuB7
0IwfnRbycj9LxnL/AYLu4upDRe+ZW1/yAR/xIVFkkuAClizI+GnnWNAc0L2vRp2+nB3l+GjPBG7s
cxu/+lLODzcylRiym09RW5ic0Qejc1kSSng3OvwfdVYk9XFXkzBy3Hwk1Km6Jw/rM69VpNf+P53V
gjLQ5nrjJ81iHRmxpSzPzNykW3/5nhrzGEk5/WVG5GV6yDBtYpScvpkhAoWwEX9uNHlaDa4mCmvW
vspwBCYzLBKxM2i13Nq79rD6q2wFH8/TrPQzW49u52pF90TIrzzB0nUmWlLMh9qoNJGOAXQ6rbcP
wFJGa/R+ZxFi3qj4di2zAQJqY9TLybW1vP7xskYP96hvHdQKXt0Q7E/x81gpLHF7udBYZpv1p0dG
NK/vnN/IL1ZBWpaW9iIF/Gyg0I3og1sA8m+lAhSb3S6z5MIC4C47pE9Ad0mfj3wyjfBfUmJVMD9A
5NfGX+XvsauWoWVb6bjLIcwqexvdhRclEGlWywVCoo7FhM+oYHjhMyP0D/Sa1UaQLYhIoKiPMZyn
SD68CIzkIlmg1ZPkOMmN2pkHINjEW+BJXbPdYbiLg1y73zs75El4hrLKhb4QSMUOlHL+g+BVXPOk
OudIvfnw4yQVxOOScLbMvVGDVmKKlrtwrGgutIA06HdotDg2ow7GmY6Iv3TchgFHn0/UvDkceUd0
6ghdmzCpaJivGG6O93BA1WgSqN8kEahs818+YB1MOZZ6XP7Mz9n/rZalKouclb3HQKXASun/H+bd
p+cXbK//ADnVn/VBVbr6pQH6/6SMWJygo5qppD5zJu/kqeE747CC2cXsrG1PJUs+U87fmcOmKTP4
zuI9rD4oGR7lGvs/RhBRrWvFr+8LvndfDtkVVNWLObBfnXAPyynAtOUa6IvL+o07TkAyDi7+ooOl
gRBHbo01moHsfxPy61vqASqau0+rj4Z/EMbEI8uN8JkKMBGyNfOnwEVnkO+5LDv2RuEzodo903KX
av0bxILYoGtb8tCNxo9o1/D0EjcM06W797XdkzfcrzNy+Go+PEkyZHDmyHtdBHXLkJc8/hRGvFC9
kwtnK2bScxaJC+CJWeFjVFJGvswE60SNoU0WD6WApZZYDQTz8UNC7FjsmB8HyJq53/3yjLUG9Tae
symOlB6aBZA9JAYIkla9XRshn4odsFLKsVcOLzYF6/H8kg9/FxBN4aW4P6vCCaG523g5RdJiXdEK
xtDtxqxQRpbx2qdFlQCyMrb3kLy3kPZ6Xu4f+R3BFkz1WBZgFtudJ0kQYPedd0XNvlAkcPA8FoVY
uHBT8dnrlmXuB6iRZAcw0SKeJEe5TNozI8h+bQysXm/aIIAPpakqVHRxrGyQXBkqtzjJG4d41Grn
5RGtSrmP7qPhvsKYr+XvK+ohq0QbPoglpUIsiV9P5DmCfdTK6MYSyGlFrAMxnADll38YICS6D1yj
bln4VP7rgGihNoBZywNAZfZkj7590m+HVqFR03eez64uMZMPD02pM090nwxDUUkY+D1u2C/I4cMy
9Esf9YYG4wBBaeykmLiMnqULfqBAciphNe/5fX7+ijx+8YE5kteHnr0es5Gb6e0nJL46du1TP8Se
XNUBxbY4UZgqLUCCpze1HlwwORJfzbszna2l3v8z6ETnOlc4WYDcOGflDbOH3VoxNeIm8pZcss1M
f2IUkpmo/lCJswcYPPAVVFlo4TSo1fgpv3fKEmaPlQ/55Vw3q52Idpy7hOrWm0XAubImcfSIJi0R
KsChRVroHurSUZpWgrVzkAIr/2QsXRdv7zUegUSMlJ6oq3LgH/yTfAHUlP2UqsJO5jfmGzNguZuP
P+ipAT5/1j8tLahmXQDiHkw7u15jhacjsSKxHUQOa5crYhR+ITvE2svwH9iwGrQVnhOf3T5rjRBR
saFDY8A3dSf32J47AjJN7OXCvZy2b3j/0EZZ4rXAF7yG5tGUmJUrhyRmCPvprW263wuX9FEfTpmx
QHpey7Ry70z0xFhjIiHTlxmTK+vpIDdDkzkRl2aZskEwwn6uNjyH7kqzOms/5vklaLYyqUtO4Q0X
ti3+KFkLTtACEGBKa7lUGcFy2JbTf1j2aJaoLgHo4mKDGmrynl9LrgJbnVUMGvixDshMUR8BVo7F
wWqXs/r0gWQSjHiGRG+z+0N6KypfUevP0/NKOtnA63xA4+o1fYjH/0PW4uB3xdiSijGFe0ugToG9
YA4OWWAfNltHav8pvE4WwfyRwyB5WCabail0MR1Ylqs8YNzQ7qsRuQU8Zu3syj3oms1X0U5ul5xX
4k4yW/9+A4/4GUV4TX39JWqk8X+N1jhRj3IUXsiKCFO2oHeUJtZ9/E2zPM4poFyleS5M+r95w9RT
jO9WvjDOfEysYB0PUFe/N9+L+HKYpZFGp+xvx/PShFqGYZdMpkUd4Ve28DUins68sX1n5kbbIMhy
1+0N2r50B7wXGgNa5zxOnnZJIhPeXixiQdzNUK0+kEGqFP8qBVyhXuGjFW2H2lI2g519NLRcuDrx
p9wKD0xWeocgg7yaDidRiqb6wDZdCOr0Ddh0SgU6JG9088YJTN7t79p9K/4vODypw1BVaARcdej2
SOnK/s/vK6CjZbvC7juy1GnKQC2JECSGXKPxpF/zPLMJ68YxeThYT8SUbNF7aDdulBeNm17PFAMO
E+f5vQKBokgXFr2CPd95WUfU16HvMxFt968kAkredFUXzgjc8FBXy/hf9Z2SW3q7nxTZArnk6Ul0
3xRZwMTN6Y6jEDFDlRIKJUbfSTajb351as9Ha2lh107pYeJkZU9/mFEepQh5PpKBH4S6y3P9gIU8
e4WsjEDm4cs/cjOA7ISY3GBRAeev8N5fXYP4oTQzT1KRO9j6P8e6UnyTapA2I/ebbHpG+qKDtbZL
MIc6MhkmqMBIDOIO0yzjPvDzLcwsa0fUBXVa0f+vzx3taux0Pt4Yl/KKz/tazGW21Umb+k3nSJP5
tJ7sVYjQ9nZv21MUcOgSAvNc6yTWa0vlngAQZCxgLgWRiKWHmgk/1V57SLuzBxSuLyeTBJG1NOpg
pvc++6g4NRrFtVaOQjKPsrSXu78w+os0HMo4ihKOUnkjprcI03UolBug2F66pxiFIxEApKYbbBlJ
0vA4i5r5Wjiam61JA99ZfssxqqJcU+cah/HlT/FnOYcW4RLeBSz7mlwanp6iWp/fCuM7LRlpgDSG
Oc3eZV02wfbkvZ2+zEuTrc8IgXquMdQU8vhWy8IDweHVjkykHsLqoD3/lyj/pasJgJZyRuXtk8dD
zBxIn32lbj6HpZ8KYb0gwEqpL2RJSejPd6sV72LLmL6M46gZTzFpX7A/AVNFAVZpEtGXz5MvaQmE
p/po55KE6TAYocRF0a3Y/xE0J/ITniZu5KpunMVB13V1SgzFfkcThvBXOvsm4bH/QN5e7FfMYFRS
lFVCAluB1WLqN0JbY2b4wxbqiDIXJoy78rGz5syb1rTsFalVzazns8xGTGzoclKRxvcjmoSuG0Y8
5tpQGtE76i3juQ4uCRQzOr8KQ1d4wqVHyzCuLytpLRxG9XIIYjsanNgkfYxvMuaXqWwKwM5G6+Lq
eJBFoLSH7Zntg4QN40jCeBEeS4mgapBYDHMmvK31xrfCPX+psD6nvno1Tf4skQSyu8OuJlHyNFR2
l+xC5sq/k53XuE2QcqwjEMmk5xf24NZ53vW8g/fzY1IxvEyo+U578mu/70fSX071D+VhnEwZSC1t
979dITzUHGric/83LIh5oE+04IJqlZJVwPudXlQO9cthHSSmsf5FkQdSR4TXhXRU+n7Y5ySsOpTY
qNMsKH9+PvbIukIiTbWfOPlkqK7LZ2/0fXkTYV5XJlMM7IOo/bVCRvS6ix8uNgmQw0FxSNGNn88A
UJO7iYbq+YJ+xMEFVkz75ukntjcNaOro3Jxhuu8+vLEjhjK1DvTZxrExLgXHZqZnvyeaPhvIBkHv
T3n6JLs4+7LzWseKlBtXPWKjECC4PNq5tqRRDTmzEIJPB93MTJe5jYY/gV2OSFMcmQolPohUVZqU
x/Oi9WscLzyEA6vmBZQiFbINUpi+9pH3NLGA4bnFoipsBj3ud5MyEqwyNOaH9j5FsTx0qUwojxWz
HgHJuEJPUHM0EjXeq+SMJCIl9YmtuN08fc0liPmA+WwOb9u7Ct3C7Eni18BM2DbF+mybVFUVdBwT
K+141wUQrZnl63a3wXQQV73PjdLJkJ+2sOqSS+F23mkrowmDDWHjxod77+J2omqeEfEdhoBE297S
7gc+1p6twaFtdOMD2U+QQXHjCt7s/VQHHdhYtBhXixziAGRnM+BB1/v/HnmFwlf7j4cE+T2D9wb9
2EjhlUms9GkJj/P3S6VWWK0sDBapbzzKNtg0Loy0Y0vBQbJH8pXTxAcytFMZdFwAYj2MsjCctNHi
HGD819tOHGTjKYWbO23qbcQedxf+Za5NMDF11qyQFWgUQqyYAmBRjYtastTFxrIiRegOxUZ5yv74
p6WZSTKIrpHz9vlbBfDmcg6kndYOTplNcJBxaq/vjHvh3PgyRN1IWtOLkVUquU5oODhYBajPfIJ7
nEtSKUdSgiv68SweFsT72r3ackLcEGwGlMrY+8CMezC+JKrhFDmq6PK0Y+PedINxginmA89XbBkz
E7bccslpDcNo0QoTCbOGyUDbO8lOhnWbGNA5hur2zoMQFPd8jjKv/bAUgjYC8Sl37EP8FSaefK0i
6W877YqaFTq2WDZy2HzHKRamBX6tiQVO/4bMqTjvU1Bp24H6Ce49IsDTB9VbvM3lBXfCP8kfw5jx
epRD86bT52SMIfVJz5jb/h0SjyvPrGH8KoDt0z7KGZl6gcRooCGiC+uwxNE3uv6bFYan4YdaQzmG
toWzAG8P6vUYsKnbtovfX6BrEmnJ4ynEKINMM3+NnfNXXhlmh2wY8LXu+cDlxrUaIv1SRyas/IGD
JEqBuSWqTQ5IvRpMXvvY04hvtXbYLHcYloZFgBWUrgIRLsuX/ZBmi3wvsCFyInayjfFtJITiB6aT
MkA7IhbhTZz/+xctU5ab4GT/iEJBd/+1tnzQRngE15YADwq7WRWKmYfLmYsTEoaHmlflR02V8FDy
5Bdz4kGd13kOnqFJ2bDK1MOoFaOpq8Jjn3Im/smPg9tQHs0nQQPTbQ4sBqSeG5dIsTC9VgZ8E/2p
qA5iR8OXlJzxVLLf4fH/2wAmI/PIkQtSCCnMEmKjrULdA+gl+7kzaqwEGcQ4XaTxaisZtlUw4HLA
UleUk8z+G2kw5clQPZwv3T0lDBS8ZUI2YrT1fIxJYIXUAblQGvbuoVTaZQi5KW8BkYXIyjPRUKrb
ZvLTRD3+p0hq/PXyykzDIweXw1mdft+HgCTpj/HFd2i4Q4aYneBApdCjy3KQxDlliWgLMWO/FkU9
+xIEVWqdw0WAHdUk4QC3ch+VzMA7/clMU9nSJwYAtSif68xzqDBjL7Su4zQYujVeHlmaLIEF7yd0
+6VgYtV0IyWTzFaEjojpVFwcTG0C7XjVLwM7Cmz/lta3VQ4gvytdrEUmyImx4YsOwZy9eSjntmxX
BUkKv37k/KvasG7wL+hrNlP33yM0aMmjmSwuvTqCd7RV2Y2AiZl59cSY1boslfbuZLWECJjF586W
pvvsvNHMBk9Td8u6LooxDJxw+rC+RpGFVvRzzVEcut6F3n9L9UxTP7QWwkyZepG1xo/mWFby0fd6
xZhwDMaJXnD5h6/EOksO8R8wRdEKmI6mrzzC8hJu0Md5LZQ71swrHt+PSioWJLfsnu0zwogDEo+0
4wZNh4N27CFBw4e+sXPH86rmLklDYEdO/x2iDdxHBCO8mo86hM6XyQAVTlNJHGEWroM2NmA7lWfa
Z3kneuNqSyDw0szNpHVX6K2V4SK1vGzW/dKG5X46FZcpRAj5jDbyvnTd1O9UA1Wyt2xN+4oSzZKA
HGsyVU5mxeHhaxHfy1vu3Y2yBXnHc3S2EmFLuJSpvlTvkP3kYwTshq4cT9vw5aFrIgDcylDX4l73
XDixYxbTt8y2BDhMd2irgDkjKCh8VRek44deDx8D9NsIIQD72sc78eiZAnVOgh7yXbNQIJHtsvE8
hRUVfQTs2foNufv3FQY/J/DOLeGcVf6MvKcsEdghu8Ur3gIfyQNEYAaMZ/txJDz1OaaZEmiXXOiC
pws9t89mV4j6vTba3gX6SCNE89haOkEn3In51QCJ1AD15ZEXkrCa5qI5l7mJzFAA6pkoh1WFp3fs
oCgCV0tBpXnMwfaW9OUJjcgNnYckUNHpHGmoGibLWNW9KyEmbIyEbNBOkO8xk9e964JTOz6DxmHf
Dx52Y9MZhLtnRbMb1a0P1uvwGLDBV40R8tz79uSTM+Kn8DlL9tns6FlrL2/ZsaJgXwSolWef9DK+
NXjolDS4dqAickeUCe6xDXsgf8VZ+PetDYnGhHuGKlOdJJ8v0Bi1gxmRoeOAUvHk/NuJ3M1mUb8Y
4LKyYKLT6eRGbzPBB1CsSOqQyV/7koV8uxXy5wsReGnKfu/bo6Z5ays2CrzfdZZ318/rPnbMVgzH
bdPJhD/xHocSA1/bsM+v6/A6R7ggb/FNKJ1Q4/FkqCfSBtSxZpWhRrtgMl8ZkUxBR56BGRzyNih/
1gqSSWt/q6W4lCw+MIvNB5aDh3tjqWJvx/vm+J2szh1OKVCGf1eJTTKhVFvxa8/IRkyB2JF7YMwC
lYFMEyGxPQqDEn/xohzohLEuUcXY7HOhrRmxRxCsk3grV+RSl1qQDSxOEPzs7LRJXuFFaK6+0GaO
KSrpI8UNbtjEGY/k8HGS81MKy+5iIzPWRlZW4JNU97Feg81Ci3n1f7ksgmmcZVS9mpXNzq71ercW
TNa1vfR77z/1Jrbn739zGkk9mN/jnfY4jmzmUq+dbpblMDY/p+djr32n9pgqp89O9GHHw55vFqy7
r6oGYBb7mVbwcloVNu6Kuk8OvVRSfLpfYonVkY4gjm4n+KzdOWC/l/p90FdNz7Smm3Sy3TAr/aTE
HEeJIJBAjihHsTYE1IbtSsXKpQFDIzywLsRFEToz6G1cLbHunY3qDt+mfyoRretchdxsPsWsssFp
/OtBzFiw+OsE3eNdONEyGmOq4Gmq8pXmk4OU1PfCA/uqbQjJyf0CwF1oiY5RAan7DDPoI/sj0ZE6
gAfoRF2bMHAzm9x2zM8nySDrFm6hodxa3URgh6NPgiILMNbe4ZaNTroq0NwLPNQGgYHEBzZoizGm
e55MHOLQlAJNCwV2US5CzxZciGJjp41LFVZtO7s47+hfsiCWWmOK4mgMTS1obl0gFN1/S9yUXH1B
GgAX7Qwn2TsxbIEoh4O2+wwnTjXRXDne8gO5ExavK0G/vkA4a8vgFUzl+0k8PmrXiUUJeg2y5c/m
/M8yLoak8K9lLCNLF7kdiCsJS+NigHcblI2JZDyvrcFshU6MBxZsZNIsJ952gCmbUglc23Dv/iWd
b9Abc/i7ihAVsC2OX9bTrZ4d81i3qpIYxwk9/jJrzLtFW2KBdrWt4Hs4k2V5Z8dfJppcfBcMOdvk
TfOefXkEcm6Iz3lDHBNKUUwx9+rXid1qcdONYI4MGY6Me0d5ppmciJ0nAn9NSimUqO0EAkWw3pVH
5QcoI3fCXeouzr46Qsl5rHn3Co604ADFt4i3TFs1VGFlVTBdNVzTvOfdlN4Br/Q+J2NJn6GXcD/J
I34nu68J7WSeKJRiNhIb8nhV9hMBqJkZYUx6QrQkKXS4TadMqKBAkCEiHJcpem4Kpd8kmUL23UpF
bwePDw+0/HPWaZHg8QDey9BkolQZNIfFb4HYas/GDvNoyqaUu0dli7w7pryx4xS9Lx9gK3GgZJeK
uNUIfR7rPt4eoKGJemujtCVOW4YgpVjM567uywkbc3VaLIMbb7kHchPRGmtV55nGYrnT9ym9nDug
KDR4w8QxOVRlW/jbvXjThkxPqx6APzd0f3p2LfYnE4xlLeXSyp+8eCUqw0ZGiD2Vhvo9jfmP0FWL
UV+Nk/wZZK0XT3yMlIrHA1leS7DDyIYufk/sUdMssxLOXOrpsbqqcP7QtMrcDCbNSjj6ZDONtWvJ
fq0neYFxBeI2++XID9iI9C6kNfgc9q/dkh/zPEKsOcCduGjH8GDYVZBWozqqkWN4BFfOUUH2be7E
rtJWBKkPjEBl7nUucsuPmZcz/DPWq364dSajuGI4J0hJ9wmoS9MOI7Y64E0rYsLIeWdMnL4YEXzP
/Uydz/avF0UbPhvR5/cBDdyKlMn2W0vrybiNAp3UjEh7fWUp3dcSxfm/pVCjmO5vOaBBxQSBvKpM
vNldGHGhzIQVvpJp5G1dn4ZhH60RNmAtY2cZUEEWxenyK60pMqzFGpTPHab0MHjKp06HLWt1O0q2
eQ6HbabpuI8Z/W7g0q70cc9S+Xz+SphgsPsw68EjcUqUJe0CLTgYXdaAlpct+tYXepakdQReBUrr
/4qa/HH3x5otxSYzi/j8c0wgLVugsel1cevDE70WWCNg32ewm5RNVMe6iwyEDSXrKaaNVFn3THh4
GsZNElT6foo7yBgqeAlyWoWluc+fRSiO8nwpoTQemmcyr3wRvjjFb3vxKlx5VDehjybbJZo+/N/1
5IYFINY4Q6Jh+AcayX9ZrFa2H4BYqD+dYjTofl98bZx+WV6TTBBrD/w91vCjrmoGN81piv8J5kao
18ZNZQ7KhBVbUk6pBZWbuTg7EdRReqA3nA/0rjwjcenVE2889yRHOyzFrd+5velP4+sDCloiZc+R
fXUVIw+xrmH6PR4xOXA2j0G6/I0v36EVme1WluvnRiPJfG+baWjZG4MLxD/3rLk1PDy1ykHF5uhX
YCZouRHAIDPky72cX1UPz5m3OXnb4bqmr7Xl0m6X8Xra8xuaJecljR73rAdJeyqe43oUxCsBFmEY
tQILfTHw5ZdHYHEd5b4vcoM3xRzUtXmu7BUGaa5wultCjcEUqjQKafB8m4sloQ8kolXBrCAs34xj
WLH/HZX0WhF6vfzvmYLtEyH9uDeVDfdmtJgNbtWX1k5QXJYsekKw9C5WbyXyxBVp/CF1O3HJi6A3
qTiQvlUQXX1pw80R5e5thOneH9gDZTm9G4WZWvClQ9xJxirfjvxsKZMSMkLJh05CrDsMoo2OOoFT
QG4uk6/nGxIDR1IFgRvk3VQMUzk+xYjS45PTY9wmAxsKZcSikfNntZueMGw2ZyDj04n7c+uAOOLT
2a6KesPRCEL435YB1BVw6n/0kUyoeY23LY9VveWqRaKXBSftolIx+b22T7JO6AuZ/oF8xtoj/USN
vSfYZYduUdbbZ6EuqDB7WflTRyFE8GgJYFfqWDd2PcOpTdW3ZkRTfKm5+FVTmWUVqzQ6Knx18gMn
ZFD0lg9cGRXl7JUQeWUn0WCGnYtrHa9NAgjAZd9GinvySzgK0Yv0bWCm3MsvQxeSRN8M+LG5znjK
yaSLSG24vDq2vkuG2KDy1bL10QjgazfcaHtp/RL5BGKx/JXqCTqY8Ho5BXCnyV08mR3Ubf8TfReH
tXRRvNPxM8V/G2lOksMbN4W2IFkfPKqOHbDh/ynBgeHFFCVk4GESyTMeHg+FYvGXJyUwW+RXMM3Q
N9RXed4kS+0XsVjawU8aT7R4RqqGO+VtuJrCoXI2G41LpDmr5waxT8iKuDL36lvVUEE5YR9ODQCJ
NHyWT/uP+rW/ZRXFZ53PYNtj7k5Lx6MOpELXwZdFq+l8DVzRkkkv9+fvWNdbJjw0LjXR9yMJpAbq
o/ihRLCgbm9N2L29oOBmH8ElQUS5VWkGmVEtbfe0xleM7HBzRC0r8bzbOt92la6Odez/2FNFxmMa
HzX2GWlcPuojLoJl56iSGlg7N6ETz4wY2nEQmaNAiG8ol24yvKM5V5IcpAoMSRIKQHf/tp4NwWlK
SyyEZVz/Vm9DpUkWvH58QSbA6p6sAm+9ZqVzO4EM15TPYIHUI7t2NRaY6FjzGYqsbZneCZwfzPYD
Fihy8SJ8GVqtXPaNdFB1GVEIC0pf+PwYNty2WIeFVgfharqaGOEV8865aVDtTkLhQPbyh67zTlki
e1h75PAte6oPImocmbdecYl5y6vErNrpLI4rjvPTNJpdjj1k2+CPcBy71A1OBVPZfxxPSihZltg4
onkfrYwQa24T+ahAzlpda+MusnP57yQIG2WsLVJ2J0rBq0VT5XCA4S1/b4rRfSx6fkLppiI4f4bV
fT5Zv+OlU0RQi7BSyCEyUvhQ3/ppar6aWyU60bovGpxYgF1IyMncND3nfKq7v9A7fyxLgscr2qcB
PkvgkGyvXJ3Mn2JJNvs7HgaCqAnowO5558CzKnE2uldJk7/8XgIkU6v7ZIKNxWrMGCmfXsyaC7vl
GgfpjC4Fhm+/EBRDbSRG+qxgjXWrquu+VhpipvtMfN/lIwdvGcGGQgcJGZz0ot7dJ+qaSW3Kr8az
IEEkzZ53NKA8RkkN2vbKRk9zc5b9HIaRSIYOwzFVY2uoMJDGAGHiYa8zzN0mpPmQdiV6GuX24K49
Cvr4HrxvOTEuVo8UPMxtbq/wf73Mdu5DSig/lX2lOwowpLqrv2tIT/WbOaqJUmFQst5X2QDiuNlX
IBdaoKDK6iD5YbSaORQ5A9Hs/4v//P1pXwa4uvUG1Bygq3c7snJ6FjjHwevgjrHCMfJWDmeXTlXS
MCzhjy5ajgtG3Soltn4EY0MQueGjaYZnREWxTW9XJhlXgbx6wruDMsMeMWkucm1t5Eygkv+lxy8j
BpnkpBYgvyQiC9Od4N3wBHonJfsIAWiue/kXQHRsE5hu3YHSTf45/B6kPMarJB3o7v6jCAP+EOcU
bJPc3URPpzHXPMHlpDZaJyvu2te8XyvCsTFtpnkPPaExN1AkS00d9oth05NjKqz8CnavYE8P8VNn
855JnGxLH2qVRy/4vY3biyskAFMWQjwP3gm+qycx+pCEGyByarNjfr+Z1IkEDOf5ko0X+7NIIkgO
g/zqEFv69UUUKSUF+AHFp0Nuayt6+O0N7F0RblQMWddjtm/CwUGM/qYHpch/IYLdwOG3Rimn2loY
1ycdkmMeSSYTNuvdi3ior8PtqdCh1NtucAy/QrsiE2wRsXOL6K3GN7/nmbynEZ/ZCepvnTAcD5Ez
UYFbKz9xctmQkFB8sDyB3bBbVvKRzr9WQ7tVDlIA76lMlkuNRDSSCOg8PsaYK1KXWExLQH0unAQu
5g9SXcJLUR7ai7DN39DJvPkSKQXw6nEZe+wOJ2MxmKtHFz3i6H1B1uvJHSXJMv5C02aEdDwq4n9Z
OJICnREEaVENQqQOHBvyXODXorFyWh0ir2LqQJ4LinD/wbPvHotet37cmp3yvf7NIWTgoXeLplnZ
H+wYt7PwIBnquFcq35nEATyOLoPSiY/Hk8nTadNl1kDkDF9sn/e5tDlruCAv91sq8vxMq9UnKlBq
DycV+vdI90l3t1DyHrYDJlTfIGt72kNy1TUaBfa+hcz9aLhXNbRzBrg39kP3oUSZN4O8Oc560zIs
YUpTpF8XQ0ePAUcHdByM0va4v64H9A17g6FiLsoEqojazjwNrotzCGnpFIQDMwWVfrFNSLPMcko/
Mp0jhACQDp1JisZ4raOgWb4g/TN7weJ5IPwY/3JnpBaLIMVdrlzQJSE1qiSRf6cfMCnbUSXC6VKz
MetDZ5QnEmgEIyUiUPQp/GfnIzFkBmAUbEW5jVptAMk02IFLIR/2fv+M7IeyoW/c+vdMiCci0PEO
dpDulq+qnIeiR7syQAMCHw9F0Rmba0LUT1uOLiNur6gabbPjA+k14uPb2/h2G8uHo8pnjxHyOR2+
gj+SpTGMIbqZwJeaQD91xLJBgFPLrv3eDSlDsXJgg73p2Cvh6uv33bStKAf4E5S/jKSy7YAdNq4g
Api/h/Gi9GbXAGXCFLBDWG3jBC++9C0dO5OBfI30TKDdHBXuB9mQ+zS5/4z2YU2z4wsnvUyQBhU9
hyZHEuRf4vch1oG1eEaD1VdLacGYDNqR8B5fDCeyykirmUvlgcfYBUFUTKra7RmG7FjUkrO5eUUE
QdCzZa7rUkf+Wi7aVlpqNjw4apnfToopQFMejrVniUmMzInkP8pROy7yfYxHv5nv9uDS5H4FF0s/
jipOjavfnapOXgH/2aUCltgR2wBkFyCU9ZNVOZL7L4SDIEp1X/QAddP93BmXyGD0wMC/1q4zuNNE
zv+9D0o2xJi8hHg39FI3tq+MPYHZNKtfOv10reiiq9aHeEkzdF+7EyIC5AeHxHHNIwD6liQLrbze
MZrDukb/VwrU9S2D1ma1s+ihXvxvPKAO0ZqO3xep4JTirFcP6DRTNs7SI7b+sg7azm3C1K1IG1cr
WEn6wPPhN+zVLaToWQTIKX5+/0LAIRbmENmumeoaPUsG/5FH0L2l74FiezQgEcEaJFUnWydvsE2o
s0or1J0VcyKlF0t10NW//Ssips1jYOc1A6x+XaDMu4s6uBBWpJZP7cSx9523QE1LDVBdBapycl4G
AZ0oZFT20CMOOm0EnTlgT5UW8etm6KSqg+ZwVfPfa4MougTwa9FKO/S/Loh+n/0ZudlfP5qU6brr
cCbwOBUiv3FZQJ7uMkievXCPNmXcf7fqnZGVGbJcUJ20rkuiD42YW1VfxaEXcEWwMEDroZc13AmU
a2IMwo/Y4HFmVMGJ8Gg77yqC9LyIJdgHkQ0B6DsHrcYYFP7d4adyKYtkie9/2dwfCojduY4fY70V
Z3kBxIgTPGGrc2IEc4EfnCTZjHrW7fdh6Epvjb6nOx4/sVyqBNbxTL7LWvD11KJMeXgJGEbCn+Vu
pf1vyitCnOXIs/Hv5IDR/0v7RdP/UrHibuslHKhFyMlYBWAyshOB327ZCFlr/87WFB+NBLVw9WxP
2UO5J4o9w6xem1SgIhn4qv4rk19otBP80+UaOZo/0Azx5Dk4SQPgbMlBFCjkLG2q8iiSpd6pg00j
Yjnao3AW204auGqaZGFHPqYRTdw+F/+e4EFJYM+W0+hqWzSBDODEJKrCxzjwgv4wN+k7h1Zn/jic
0e6LqzF3OP2eUjp08472YyptXSFz17UUnZDprCons9wieiBg7hkt7XLciZBjxUKlGWdL+ttV9PbY
E6P0ZQ8F+dzCfcs2pW6Qgqhz80S2YFevspamwNaOHFAr+3yLgcXjU5Lwo6hWsN6gMxExnLWNIQ2B
4UPgDGGRjNWlCu6yFtr2z3dC3M+pnx3EcfhBUOP61Hzvn0nMz8UgAlfu/U7ojY0FOxPx+ESccBpL
Sfs5x30TRKD7a0EbvYKIBoKWvv8/MVeY/vteePoeZbIntb5W/90hN+s2ZWV1GIXPbmLOXNmWa7lW
CAlHWwzfT46DqjYXh9zKl2JH1/uGNPBdTmvGxkyKgnTzgxNtqQ/CteW6ZoUw42CLu+ymK+pU2JK9
7cs+zACa/Sz+JGlolrZ4eOHZ1Tadc40TLhbZTcfXyLqFQ2WOn/vJZfBJHFaCj4PEA6HHQYa1nRz9
TwJV9tdW2xXzYkvAqlZ45f1emixJ0SvUyzrktGHITuUElEhJaPRCu+u8XbPh5rQJ09H2AqZZRcr1
x1d7VH2TE6Tr7bCeAdDtCtEwchI15OspMWSwj8dNmtY67ZWBJdUJckij47BaKLmFzX3i9QKnd0FV
fYqKio5RK+HXa+kOYYATX3B9RZCldXRwUpmZVe87jewfHVFNNpv5GA8ZLDdlB5TmtfPHlaIWTE+y
20JdiJs+DWnJiOi5O45ycOkoEnvWGzDZ/Aj2jIg0tSO+Y1aFIosbggTIyBJfnZ3c2QQPBZfW+Daq
iaZXYk5ZO+D+/RvAs54Me2qzq+9jjq1gcwcSsHXitw7pwJmtR0eC3xiSzPG1NxOl65s4pUhxlPLE
37z1fBrbVQnwoykfTMWUNqMqo92s6UR3gn26kjw1a/tktvN+6EWbxayms5/2CG0IkUVZewRJ/meP
kwvQRqWzyOBhgF1U/JviQXZbDnprTuCATfnKKQsGjNdIHxTRIq9uDzRaWchc4mqFfYtyIL7L8BdQ
nbYxEy0YbA8WbcqKa2uM667DPZ9K8OosvIoAiHYXT9f3iOukKsgZukLoploA0rpNSm2Q4XOv91oZ
GyuY60ac4l5rWdegZAUWxlfGkg9kDxL6jdZAu5P3+Nfw8a+YtMX9HVfrzTQD1nA8ybBqDhnyd+ot
LwUCqy9UMXBh3v78a+eKZW7e5GbxZlZmbqmge+fLjc6vHtzPLpynBjKly7QK/u1YqMel34us2F1+
GRzidzkgej19UmmzMuwC3mnioLB2/ntLRIuUHmtkEFtBxYvwfJNbfoAsY2cDTE1fnZtVWDBmLYsW
Rx/+56gGrd6taDXbpO2SsGVYyhMAIN6HfiFPu79+q72GMP+oZrC+0LunacKZCWJ3Ow9QX3wCZQ56
Y1QoIPxYwLHsnZkahbiJaPZ8HMHf97bEIP45MvjAXC0Eq11PtflEye7781hzpvDRkxITEAwyF2Ct
+Fvj88s0kI1XgLiid1UElbJW86TQpW0gFgmzHeMXdUa/p9F7zMQQZPBKYrKZ6gO0X8fOKWhFhWBF
0VCjem4OlSDML9z2b4rWwhc/WAam1YWqmOIJNKl1/d7kPxzCICVlYDDLgABTKJ5UZYcwlaEBfqYB
rT60ribpm0v1uu2O1lHns9WSSr01pSWaDZVP+XEDRsjSV7+CF6Gn1OS4tjX1tkBl3Z9hrycpjeoL
r3FhtqzLND1REXo/oowUTAXGOnq7v/Wu8ox/BM/nz+wXlzAPY51ZEYCReHELPZK7Sf6iQSrEGgzw
Qm8uH+QSrQwW3jKmRhqbSct32P4Dw1mQuCHzGWYLc7bQMJDujzfrR4DrhYGBblzT7JqtRdVdusPN
5VFmwljT+j9gTjBJLl7GUP/asAS4UYWdDFDVT9wYN8IpfPmfaR90yua31BdK9qPYgTN99Qy5wrcS
IDxG/edIDZ04AmBbT2zo/COscGx1isUEyNjwxNI6D4gKJCoSTwoXYRTdcr6vNP9Y9KozkG75IpG3
jLiwKQ7KAX+/+2rlM16EN72MRiXxEQsJ63p8cxSP1XLbuwdtMQORTLyrq2o2byPDWeRWyoipw3eg
VZEr36GB9y7ExU4fyZMWntjUULmcOnTzEHZh/bxmXsJ2PSSXGWIClQtOgYLtDEkmgF05R0StZaol
DRyaeoDB1QkIBudyC2NTbwo14YiecQ7eyjO0bt06EloAIXa4uJxY0UTuYpYx+B1KvGgbQf3Q2p3f
R3NyLTU1sPSKNwOR0MPD384AWR7vusBW0iBwmJzsm1rNGgqtWwZIsimFn4p1F36OOrTVnu0Nu4Nx
jIokRaleA1lvo0OTksf3/PT39uC1naqedoa/0RDeJSKpNxSoFzYU6tpEJd1bqYA8DrUZIsvvQTZb
YKeXVi2QgkkNu0lKACv/4n/FWaDzi3MTqbN2yCRzrnCSxrLNUwlQXs49MOMOOqvCkDZE8vf2WIue
FoVSDdyd90i4AcwK/gjW/iioh0nANX1mANbX7pMYTqgMBxMajdFnQOVfDoZQrjFjUbLGeuPMvIpR
GaSATf8nfgpWFwh7BPvGPqQ2AsNYXSwU0r8ngp6MKDE2BVYpaUgZ+m4sN1q0Vh52fZLQ9cptQ23P
0eEcBH6I8OJX9brcKBtvEvPvEy+sBPaHXQnsJ6vHoMTIiARGweeqYguEsrlp+TbEvZEbVolgRDJx
6QjDl4+VtXepyJFJIOkK4qV9TxlyqJsphjB7FX/zcZ+vNDEuFsT6kLBXshO6QWGdUZF+bPqUMY4V
BNeLpQw50cLQ1NjlO0L8LVKQH5NZq6K6VX6q99/cRZlxpzSY5ssADgkYYWCI0Wxd5Tjhpj4nz2yP
OP5uAPVZYRBXC3/ppumQrV4T2A+yz6gcynbiouTITp2XG1i0p1OAA2X3nat6tEjyrm27453aClA0
df4Aeh8Y5KdDqlX0JJ6+QbrDlqHuMfXqz3dADBqkNmk23ukD9mlwtgXk/qqBs3uG0W3hpOKcsLMm
sNDd1k3+KUDv8/+KDnwp/XvVCqv68QWGhNVzqT/jjDP1TwEpec67MrFNC3lrTXhRb23R0PIQNDGX
G+1B2CPsnk4527sEjWVtbpVjArBh4p4dbdrxeraDoZ87mgj1tBYxpOI9LBUoqhVD2quyMwm84he5
Tsyhe6Tg9rKlJu8MZguFK6IG0T4iJzYSYC87eq8cYgHhzg8tfXBMP1HHXxs/YpBIR91kmRPOP3K/
B14hze9URKOvNUVgzH3g32qhURB/SB+a3KHTNCLl8nhePFHK14iqCS0wSMkkDWmYHc6zoBddJyq8
roJSNPIKEphZDimjM6ofnvSn67R5tQIRa+PfVMmI+Lf1XarR8fDHnikw2r8LgeqAxjFn4hwLj/2C
nIi5pyKyCVhN2s8XJM7Q6WQM8k1soFdWDa4G7k7cbkwRP3t/8Jdg9JgN0K9eR4Ybs11IV7AT7Frp
C6yNdAh/ChIsKZfpufVs1q/sIAHPl8MDMxXilmCy5nBaTj404Ffv7+CH9GjgjuOMmZn3ul88m94V
bq9TlPz3rJ19hWkKbEcx63eU+8h9GJuoGEqy+ocbFYQvcmB4f0rTg8t2RKiVJdBEpofS/fGw637I
rGv+RkNcMNZvFfI1Gv6a7VRit73VkGB6Y+uDUAqz3ltJp3if+dack6zYrt2aPUcPGFLF/DaIjrNu
QRjfo9eKlDtHrnb7aqlUn7oV1aLRh58QaHYSmRvp+wZOvdViC93/Iw4jCu/RrZPHdocEcMzLV1DF
FbFZr2w1ZUD5yAN5baKC/dXqTMRz6goFmprxrAOOzH8bnCRd7kSbdPw6nyeP3BDKU8N+/Apf+qEA
xQN2yV1m3J41NZ7P7ccIRHPCl8EYlcGsYdmSMEDh+6KP3c+fpMrT04dvwJKliUu6YaJB+ljMGmOa
o3OfdIHXX3jCPAEr6mbJ2mqa1RDo675iLhSESdPTOi/TU/6tVaer/uOjLJ3WsYICKQ4HqAKMn9je
zj9tz+BP6T/Mz3/ZyxRqM/k2GTXvEHEGN1RD9z7o6MQFdnLY1cvmB1Eq/vBAS1QpeF6egHi56wOt
CDKzoupidFXjm5qhhWyuAWz/wKaPu3RhNRLsieiINdhIte6HsFY837QiFajsgjzVJ2G27zrBSBfR
u3YL+9kjL+4Ue7ZczDhEHpVHKfwbetagGhXnOWJiYyCInKwyg3q/SR9a0tiD0OsNPnZJ3p2Chg0d
X3Irn7lVHPQ8r6wIVqz7XtWSeeYmHpENN/4cIZsrUqv8p+jFdqthTT6jlDc5m6ehl58nfafTsfm+
lS8J5R5xV5UQbVvkCoUlf1XPJ5hGbVmkap8ip4zgIkUXmC4QP/p5GiCK2GosU+hfMpGbbNmKHOaz
n0fLIRnPS8iPt/vdNRmbUeVMougjyvsXQSKpTGQUnzilOPVullq8nALyrJUTBw9mHQpr1vP2gfWD
0dGSUQ6xBTSVK7Px/9LkV3ZZUZUJgKgDxivU5EkQ+nkBX+x8gji/NttUhN9j9GAEL8ilIU7nkW9M
z4V8JCjX998UZatDCU/Cr9StiI5lMZJ8okU2409msg/IS+8fRo4TFzYtxhKC+1kLG2zWmk/1hf0b
DtZ99U7KXWuoPhgRKZqZGq2kLbPvTWmxh9OJCelgXqrwjx9Nt6fT/UDmj1DHCY2rS7jCVGBVmfMc
JOSuMUWJ1ZqaSVVZkU0Yr9otsBvjDZ8XxKNHfqNkdftOEyagd/movUv1hviUyur74kOcKXXQJ02r
cFALZ9aVY6SQ31xBFXE2QqZ52Ow9eJkaf+NfeMUsdo8ggokg2cROw7h/F+eloq7PUrCOtv2t0U4X
TtdFhmaEt+HP93D+qGFa0I8TDGAatASt5bPaBjivdW4/jtlGaA7/nUaeb+pu4ZNhjv9VEcv8hBUg
SfsDECrXgeJTqFarxUsrcwoGvpdTIsS+dYCT/YC3jvnWOpuA+lzY+40L/kSwb6EqDeEer5X5rrDt
MrHZY060lM3AL/WHOGeil2VuBx3suSlNkt9vhJbi+2V+KK6xG247vzNxsMJNAWICVJUZmDxWG53N
qI5Ch50r9ytF0oVqYxaN+yRpXTxBBPoDfg9bEiX5+rKxCb6lKuhiWtVTejYL9xg68p2W1lRXw2S0
2bAyMkiAo64/0IwkPduZvz+PeBkXaTL03wl1/2w0PDDu1eZR5UrkzuY5K2HMAYbyWFR9Mr4kDO5K
cTd+kVZS/++1xkTok+4Y3vqLu6scB9LRZ8kvPtTrhiIe8CCH+0gzrrFvZaOiW10YNnT2Pua+UNPY
zVs6JKjlb7rn4xNW556Ay1UuWtt8bc/a8EQuQQRdpfw6UOjn6weZ3aqQt8an4tSXg2bn8zsmNdVS
4U/BVKVfKx8kVOXR9IxzzQjXykxr6ZlPYSFoL41K30dVNznOmlVK1BA1ZBHnnrikn+cK5Vtpc1p7
LkQwpMc3ZCo6/UCORcDlZlAV5VRON1cfDKrZaRXgJEPqfvZrmDXfzATZ3Z7FP4Vut6MXULx3Fxxd
rHwKnlxWbYQytGa2HenO9XCUNB4cFmSI5wuECpzl3rPaPGds6Q074f0snDbIuvII/FemXw6QxDsY
yM0X+0bmakvq9NqvnOq48X3cbLC+uzhpirtZL5DGPY+tdWciKfiJ/DURmuuaNLhf28CzdM9ZMwzB
o08iCWkgyea9aAGMJrE7bQH+Vhjxc8oZv1fZioSqtbXHvV+qOC9PTfQPP58MQ2jetR82qpxje2Yu
bE6gIaBEj9uOqGe9CB72s+E7sdvHmeL++ShoVd4ulmvCecC5qhLew2y6CXiMXHeYVpnbSh7UzdaV
a72wvp3xXey1XeeOSbOUZZ3VxoYFQuLQBLHQfNlZETdoGM34jb+Yh7UM7m3GM7dyZszoGjwJ8/yW
lLOcO4t+ycVKLWeb7d/bn4kiTjhQxFQANSH8VyQwzLXoWUKLJ5u0cPMVFBGtWP0mRd2kTBeU0RR5
bFW7LgBLIOEd4SN3Xna3fOz+G42aGOpQWPG4ZV3zKAApco+9CizmV/NTbWM+eVgX5CdY8YJoFYw3
9v/dzum1aF4tOFo2nabAgdhpE6QZxbCREKmwr3FitMCMxI6UbMhAaNs7wmPVvkDM0m+h5XfSrnEv
jeduAqZfEfl4DCsjRPCXmBBAADLuojkNUYVebFsbxg4pJi1Ghc9V95Ngv5Ct9VjOiMpYY09P1Ess
rnAuIB4ADwY0Bh3AtQTGZhGBpeKkr+qQ8/GaNj4d0lSG3YwY8d7cQTxthX1var62JPYnBDZA2I7/
W4yo0iWN4lkY/Ey51q970lj9tT+YH8AE3NFAXcbSIVL7PwlAsPs2uW9ysNXvy+LF2InBuhK3KlwF
eyloCg7gMrWl35iLhdTgqHKXhFZX6zTj7anfHKZvgElO51GbbypDONkK9qZbY9uiRuS02ZWnJAkE
2DI2Ty0KROY7kfxAmsfCHV8Aws/uNfYpYROoqsV0heVbUmXcYIfRvhZH2mBZUJB1mYpH8fD32Ybz
3wM3UL23oeWUMdGFUfANvCgFWW9m7C3IAgp3rW6wrpkEU527V5tzDNI+iqeLDa03Kb0C2rXXK9/I
OnKaP3kSQKKH3ePeLQ62jpzgk1ccpjtjwfkskfQREAoMrM5eOa2vAHi1KjDyG8XCqC8cS78bm1uy
y+e2uM5NHfZnzD0J+ihTGGmvedkS3IU9RT8PQ9LJ8TKPu5/MpZs1C7Nx9xlovGIdC4TCe2KiMBMz
UpbkSQlK2LJG7OG2QMVm8VgYlJC1zyfFcf2rPdCEN5DPLGXTiwjBX50Vj+Epf6yP0n/dOKacq6lA
ItShdehlhO5Ejw+9/1qcBqUKHnDcwQHg48XUMe8kxLzjwO6pEE7JwO35bMNjbMjNBkPUG4b6K/VV
0x4Y9DLzNAehskG9VTP7ZqvHaaFUWUVOgvC1YmWh2Ni6fTlIIOicvWx0dRYDS5m8SbqY0JJXHCAW
WSkJFrEHUKWN1eDxs1IgxIjjAqe/x/LQ8g6ezWl20+hHveEXpJY6fXcaDSOmEsGx0baY8czf3R3R
LShP/qx6mMOudCm/85f9PYAP22iOWL8YmcWyUN6UFlQiSuRWO08g4HKbuoC32F+R6SCGuIrwLrTw
hDGITQAgRpyBpqOg0OtqWJ5//ILjz66dq9uVgPiYobRdcs49rwJ34Hylq/CrQgNhAZrOM+buIuI6
jGNx+Q3vDuPLEpmjR+z8J+7guU54g0nNA/tVEKPNogQ4Zvvy1BunR94AduWgx5hyK+4yuTzAmy+5
t9kdwNtIn9CIZUFTmWgXnc6NByfvnezfMgyIBNoflMLh8STfH3EZU0DgKTitG6yt293fd2ip0/Ft
lGPDEzDVRb2BNTUA9Vou+t35Qj5/NCDN4GCeEF6Yn+CXxG4JFS9q+OtilBxQh9mCmywAHEaSs1L3
BzutGgOo378IZqkTKrAfzYmzFVEXUHZpPVq2xmFGudZTNiTYN2LVh6r6frLLW5aJoY4Y3VKMeIMT
3S6C+a9rRWwLpLHOpq+ys5pTOemDZT/A8LSKHZ/KYPRr0CxxAXRtU8IpnRMpwiZzr4rthl6A4Isl
yqs7IvX7YqGkGbGRHcMFUnrRtVuogPrbHI2X5DcDtTmbNVTLs/zU7kY9J6RQrr7zL0+zUBe8TP4Y
Fi8V1wu0jymrZmXdkxjCGiCRWtlcT4cICtvVNe5qARp0HVv3DlXvcIw0F1e0rKu2CKJk8xTZrxMr
PX65tcgJ84kvY2SGlFzWdzh9QWsVw5uku8jLdotx9R6EGoWgHzThaArSiM3Njgq4nSwc/yrfyqpI
Wh9XM8RI8eI7S0KdtTMXfWFtWHvRlbfZGZDNelZMgrWd9pxeOKWBZAy4klIGOm+RTo8UKEKMC+YZ
gL0zgN+yeI3V35msbl4yv9eIgCRcXU3uhxh0bIWQDU1Oo3d92XFCvaT+VxnIO6z2Gr2uuNIzMr+I
PWAFveDjvn1sn/kMdPhS7useg7AL6C+3KY7dnLbP6Ngd+BgVjVj8Fo35sI0sgGTNHYZtBT90pOTb
zx1UKFHeHeaKkjwU2NHzUh3AQ8y6ae/yTnL8vQAco9FvN0TpEOY2+Lz4dh+LUnkbXvZuI66J9WyH
7qWozFwOG9F4WhqGa55QnCmTVowcVQYSW6iGcdqFRWh1Rm36mRaqmRuT9iIbHs+sLTzyCcBG6qob
7PZZi02vNlGefidssDqhqcwLxETGiT+tJSIXZEC0GsjFSr7yKqD48weoiuXhzlzY6hDEQeOA9oZb
D1963KtviEakyf3RAB4+5bbCAETQYRtO/ep1IbWIsjle+wMmpPpZeuZGaeow+Kw26fXDe119D//w
PDlaTR+hesNPu1X9EX8W/8aVjtfu/QmqpukYasMBUaeblE7vgXiPGilktHXBascXlCAmhXb/ggAW
NDeMMK9pnK73QsxGTw1ImpBchPFL+0LOqpMhT7dgAVbbmOtQbsSgrwRRU/wP3DQhfP7ECPCxIo8y
2+Li8WhWh3KxBStqds0KbDTAHfTnjd7dTlh3vNOsuDB1hzsj31quG9pwKkKoqWtapnFxatRoRMAM
Y1HqjKPFs4OdeT0cgCaRrXHLEhftgZ9wBkCay1k1i4G3s6TQWcLqhzsl4O+xwAYPlXAXY1J6xBZj
RQ2BQqCAti9mgzyKdYzztPOvZ0WajJb+ZBbiCs0gk7PU59fpJdkvGpHk6XsAQ29hpQQx64QBmD7y
AGjcAaA0v9v1BXm3CfDpWzDMklNDTeMaPb1c1xLqhG79YvOn60H72hhueLqYcQJpqQfnq20MerAP
b+LXN3MEGrsVexYcxFQvnBviXWKsLJMknWhy0B0rZWGX/1gdg36K4n0tQB6TSDmJxaZNS8OK5gT/
dMMnf4vbnJtHc37AbXSn15jlVwrwEICSWOjBgBMZiHIaXBQOZmiUUBrtxMCMYMmf6MXpz+Kpd3GG
lorvHoIo1mACGTlRGYKPq9VE8v2R/yI2UhXZU8Qi3u2X8flSRaH+qzYno2Juk9jSUZK4AftKnqMj
cgtR5FfURTnmH5ydpJKOHLVSoh+B1ZHcEfe6uVnNCB1PIRny4vn+5UnD+bSo1Xv3Jpn3eoCJA2yL
GmzIkB3sGJKkGk8fYAJDEKbOFgkQ9XXhI+S3iMsn0XF+TzczO03+M4EpIFbvjomeXa5AXYZ1xLEJ
L84VWlqcNP59rHD2GHwchvnVClKtBVAcE/XdEveCBFrYlIoibeJm64goOCYqjVvCbOqNWJQ3mHRc
sBRn609eGWFK+c+ggjt5GFTYyyEAxeJ7j9Xu6fRE7W7lBpvEubL8+qPmbejiyqH4Yl4vVoTXsFVa
fDZkcLLl5+869Bu0Wbf/ytsHEBPTJ7NxSwEjvNg3hP4g8LVSkWMjVxtgI9sTZhweSflY/z5ZDxSW
uKa7803VBNcgPvnuOseZs0AVWccU2FubslEmu6w09uXvBwEBEgXhMECG9bf6ibwqSnNeofem1Dta
kCLUc/zc0qJn7+Oi5z///g1k17TrnxcMgm0L7x7D/HyseFhw5lTrNc0snidtn4OGX4kzhLJv6cHe
QxHpm3mAPxoKh7gRcdEx9shrq5rfRwvV/xAMl3JzbMUaRcjoQ8GZGyDtIudAOZF2Z4735IweQkXK
gsaGlbGAcKtYwiwBZDMmmFirDvtb5mVUzlRUp0xo1Y59blh2Z+g6GQL9U8m3GeNzoc6BjadUGors
wJ05P0nyQ9qUGVXq1ZKBmBJ7JGFldkVB+JFXZMjxGJS25KxyqFhnXSbtf1K9s6OBy/EyO5Vh1Z7o
kZWzfb+UrrmVPUm55scnQTlQ0zPHtM6X9BO3EWOk6agWFX4DoTVYtZMq2EViVBNOAKs2c+Gdjrml
SMjfPcGuOTnny0xE3pIFfX+LPyUDaOmanOYGLvEQaquWi/b25TgbC4eYVfM65Yud3tOSNxZnMGVi
aKqzFfnSe/ZPjbKAce0Skpo88ZHqKo+feVq3l1css3dACoIXjR/1PtCzUT1bUZt7wPKa7V3MiHJg
+eEn2WbiZIlksB3rAILGvyjAc4Mdn1LFLrFqC00Sja4JxVu3jcX09s/G8L2+uzuQfky2qN4GFHpT
Ox9lQGWj/TUrWwrZESY1qVjD7x4agq8SppAQEM6da3xagw6n8svSvJNTOrZ6RFlmuUOKW41IBeNN
YcDrLNvAIFY7RgvefNSTV4HcDrLY9CBRHCDdqqQJzIouCETGcNKxD+OpIsVZxFteHV5NnFADCA7f
XOJl43tmPDqzHvw7buZng503jOW/PI4mtILCUj0UKzSXgkPMTyoQuUFc5iqso1dFzCO81CeJn7e5
KQMkyx+0UWsxDoG63B/9atpo/eTBsxCoSgatvhP6EsAWsjNvI+aPCKXesHdbrn6xPsiJq8tUDgeF
QWucmRfKHV/z3IWsiZu/LG7pL4jm+9AfQqIAzLyMGn7a5hqZ8KOlx7fWik4+iW3d1vG6hJHeRQqZ
xIw5TwCRTb9zvJwfi7jMmBDe1pyHk3ajg5TMzc2ACdkdhNHqqlqYUlYRniL0T+d8vgia27WIrC7I
7UJld50UoeJEzo4HUrsUAup6M/7Ue1kjpVe47x3wn3WrwXTih5k0ThztPGiuqz+PCV4Uo3gh41Za
Nk7FrOZujkBXlnIF1xeISmRznY58m3C5bmxKgfMKVGXoRGKv8MKND66r1cEuP98atJEJwwrwW77y
nrsQ3cGeI45g7tu0DNWc4fykAX0KpFdv+eC9OSbdO6a2TdltjgQfaZ4Ly/P0bbHNpefZFMDDuPUi
LLKA3MtMe2PL7T2r3ngUgTmTYOv12UIxEszAM7H36nxGjxja0l4veZ0d9uLxW0Ach0YBiB5tCJLp
4d/uwq+TCOCitYiP9b9fIVCovbD3iWA63xqgVyVJ+tRSs9UxcwT9S0or3GU646qA9QBuxajm0KPJ
5NfJFw7BRVNUjvR513N4LziStL2T/l0PKc8nJFmaLGk1TLcnOExjh+xm0ZPXE021uVKFhWB8VLgB
A/dq5d0N+vEkH1T6iLgjNxU4BW2dtwtBlloBZrIEsObTXhKTLnzbigwr8m/C0sn4lZNJ7qTJwf4t
2vvatWK4u1YMqncaJP9lCFyM6bMGlQAte6av1TgEA3fYr88+gJAJfwKIeQCYAvIb2xqCguwER5qq
MkRslZQ81eTQII0B8NwHlRjAWfSoH4wc+Zn7WVB2YKTIh8tiRMJom0TtWqdKbDKbNPDff8+P4GWR
iSrhryM9Poo1oI+ek0yhRAEbzmlolrGa9C3zAM6/XachxbdzoduSt5Bju94aKElDn+5ksXz1c36S
SS5x9iQuZz93PaeIZN/wtjKGCphP1usH7DoLWH6bcFak0+kkRvL1e9XgUqULIw+q0YrnTtMgqJ9B
lWPouCfTpqRFKCvON27NtK0zqF/hNgJkm49gRZTOQUukf7U85r3dWuasOr/lmmeWXjYreQ7ssYzu
Z8jPCyougWfbUrSfv53SUcdd93TFA7Vm2kQC5gCFEn6txRKRXnpXTbo0OXq46NINjcM2wR9GNfto
0RjfGiJLJTfCJ0e/EBGTOwp1QfhpanGIjdHEXvLKDrFpFnOdeWl3k1v6dm4e9Knz1DeknsqCX5u8
9tE90j902F743rjElQERIpzk79VBIe1NgZafHYGDqcICYzICcWlldaqqpqyn9y0gSqlkh1K6Bu7c
oCv+tw+qr4q0oqKZ8Yv2BsBHoHjzLnSzqPVGku0vjeGfKwK1LchtqHwPLtQ456eCCC0Vb2WYi/28
G47WU8uKwEZKM6pqP3QAb17k3mNrsYZVD5W/kZTGNBi3pjS4NavxanGUx0eiHAuZk/5Kpwu2Q2Pr
xN96bqinz9j65hUcjoAlBn3fsTJUo7KVw+N0T+sb7WF3yI+q6QdAnVV2TfhiRApJi9PKc5dirhPv
N2Yr2Hn0BQrK2mpn2b0uBD6GSmPDmW6pYYSWgzLu9SsgqVrGcsFf/eouaRSOFzEl1bVKH7PQpGNy
/YidBw/TA+aS7Hru5RrkUNLEuACqSe0K9VtXCIb8l64JwaJzYnQcuFIQMkLKIjLfS1Tj5KNjeFBX
gAUgufC42NCs8wXPzno7k//wORjM790jJarqzkXFu9uDJm+JETP+OBJX0RvlLSTOmocIi/zY6Nyg
J5yvejrIcXifvt26tl3q0XOw0Zp3N9TVEYQzAjq5U2+1xD9XE4GKQ0/wQM5m3fmSRHzu1haNRFZ4
4AEEGxd7XIzpmCVeHA7TRjJmnFwaM2NRDCEYk5+QaGwv1O/h1/4p5F1t4gUmXrzG2UeSN9p8cDPo
sGqMMuDQZh3RtrlDLdEInSBTnto+FaKQlMtqdsG49MCMJ83jSRjpOgZ5k+R1kkecqLaB4yHSbJ8J
65Nqw5tIUip/IXK3j0LmmZRzXH40W83vl8gzD/ytcji+gD1KKnQy89seGjhGFkrTmlMNHBQNcoqE
Qr0+eyHcwvk7//cHyBfIFucEHOfuD0p5n40oYDBv6szzb+OM8fPRyDLG7NMChnJ5ndXa0O25fNy0
OUmvlkSE8AUssroMiRIJFGdEJ7g0/BHKPJ4JrDUHbh4aAbf3IpaBBmgrhJaoh1wkxwzhFr/4Euro
kH0SA50SkUmFl/NRYIYC+7d47KzRF5qL7WT214WGLQH0ch8CQVLcSyIZnuVn37CBClfKAJ49bB2m
RcY4/K5o9o5lBaq1kB/294v8ITBX8mdzDC1VkQPUM/NCLfPGjEDkP+I2QwxqweqqgWpb+/ftxHHo
ygn0UfQQsAqIU1mx2qYeNzGu+AyfNf2aJkAnQFEpfTru9VnAEXkxPpU6RVL0Ilifo/rlI0dCdIgD
eUGnleYl5aZ7oTtHZMYnwC42njgZNsBROEpPCUjhGJuudeHRU9tfmWTqRHGo10tM9R2mXCU1QiBN
YqnPhmQvUr6v5CvnIQbCKw5lfo9vAKEoEMGAjqeYNOq/6wTf8mZrWVnjeIs+wnFX7XqdBH2ecLPZ
zRAYX/+GYjUfoYJHJI60kTQGYJk3Pzw+cFumImefC3IQWKMHvQwisS9rOFBya0ylmSoEqmyjjMl+
6GVkqif9AJe7M7m9lq5H1tDIYBcgic1aXh8X6zGVa1aTtxIJzvMPBb4BGtOSrSA4j1JutqNk0dME
B+6SGvVdfXedG+9Qz86fNRWO2lEDWUM6kQfuAG5xl3ILfT5PvDv4Euk3MxrO/uMvwmJz02z+qCwd
/fh2Bh0OWyqax9w+s28dujZrYpfpvrFWlkQMe6l+DtXjDtT/gAu6bKWpuLNQduYuhAoP+ylxo9NI
JVZBzfqteKG4CDvNJ+tDRhuusU41B5cf5RBpK8ZfzxqsAghB/vWIfz1HfUJg3vJ4AY4RAIgATjO4
ebQYjM9qUXcbszX7sCCwELvPw9qNWaHYi1VQctciB83kEugzIU5XZMCZbC6KO0FHz8RJTfX+ifiP
zGYDQRGkBGizq36QPL0UL6rKRCfJPCskPPyqOdM8a6n4BZUAkIIgwB3kiwSsTntp2bMTgM66UNLC
cM2MqWCvIN+mXm50lwESRi48sCWBM7lIh0N4MGMdGTMBzNELfKooaD+T20tMRWtXwCpUZDt7VLMV
Idji8sdRxuIW00dvntbho0KEhejLBKXW/pw+g4fv5gxBltNED9demgj3Rwe6ACqE0O5goL6KEai5
vxsV7x40YHXuUUWnMUA8pox/oFt36ih766CP8VvY7aHWp39SrFQeYvrexZnN48fnBVXHgy1sTUvF
w8QkMKylC6bdHG/j7wNaDswhCXTruZWSZXNc1v9UHss5X8oDGe7Ycb7gyE1ijZMwG63zyHEPP0yV
NwU9yaMGE1H5n7NdAwxAPXOVmhFFD1nb/9NvORu1M6SiIsEKGo3eZuc86AC5b5VrUR9xJ4SKuR5b
njjEUefrs1UnD3asCpOvJg6Vh90RGR1HI0f+ZtfeEnHH1UvC7ciYe9i0UX7KNgyB6Gm1BWHkixI6
LoRtDPriBU9RIEhE2g6d1XeHhIRs+UEPbf91VgFzmTqsgH+s/41FbUmRX/9DU3HroqVoUlAhIpFf
QO/b/LbkWi59hvgSgug/wOXRA+IJsdw4u6H9/shQfKDMFx+yQrRruV7KCa3AOHrHdJtI7tipgFTI
zt/0Vf0d+KPWGW/Qc42R9Tu6w/h0SIIv9ST9qEO8vL9A89jCe33SvJFbExdfrquVlABWikDKfdaw
fBqDQSKOjaAAJpsP8q6sHm9niMdyV4587/zpZ33iytYJ6ErfM6bW1bavlZ9EMwZkqpmuQ1DO6wWt
ibn1rPDArSI0fMA1tHssO32/V4AEy+KOBkA+9PKFa1aS44+nn8cDQMtw4CkeEs5las86py70Ftjg
STjBSBIj9mtDDwRYSRqhKX4Xrq2Xrq7Q0GmnQDq0EGQPoD7JW0rCdp1LRoGz6N0XlvUGtJaeEoGr
PAiq2gCqi46qaxEhs32d3Vs5Xlnl2BKxerHP+mcgDepQFhMVW69c0dgUFuJzFt1yvH7QuDRUnEuk
pCiA/j7vVtyj+W2opu4dB7FrwMR00GcBnzT4tgVgk+/Mpvr/Em4qxPEX+Jn1RATcpNQoXZ+OkUPx
eDctEfwOtcxJ0aDGaViXSU0y+X1lQLSAOKb/OAIHiDL4TYQ1zjTFo59zq4Zo+s51jHsAh6pW06m4
k2QiPzCkg+JiC5P8SQMeaRlKtVqY3slrEzm97sUMq7gwV9HtYQf7rY9hpHOHLyGmpC/PhRz9BEy+
CiRqsV7b796r3q5doCLf/RCipfG8ZMGgKHOQPIuYFqgH62EGR5Ge71WiuiHEDtKR11U8Fnrt7Iv3
LdctG1wj0TFijp7DONu/4IqiaEIghUV9tFP01vFgGjiPM3LbnRToM/epX+a25o4nolJoib0+khCi
4D4eEh6gKTpL7et3E1J6H5giqk4W3oREr4K+k0BlDXFjx5866kt5b7hoS/sozZcmU0S3A/7ePflv
qdjNqpjeureVKiH8jcBUxsJSbWI8vMyixN02D2SLptf9841F0ALFWoOgkCDw9hpey+j8Doc0pcQC
1GBsl2Wz9pJSWCSRMNHkAcD9SHp9C6fIV9BEQPqF1NfObmxNKRstm9tWsl8MzquXPZ7G3szzTL1R
CcQq5rHrvwxzH05uTAOeJOBGnknaUI3HEK4JbwFUxj/VKrnntFLPc5dxRI8ZBPzcIx9jl2yaI2jX
e9QYK627Kq0ofpGp9yGqM2ymO87jlDHnZIgnhdHyWhbYf1+SbAxHJ9lZNPj6OfMmb8fH9WTdpTRo
ZRsNIH6tKqW+2xb9LJNfAqCgzXoh7iUjYMWuA5QREpfphkIo/93YLm4jfninGUoiIPQIt+p8FLEs
OFYV3FKCmljb6xq93jyqPxhdo0njfdJM7CMqesvSdrT89VOD5mLauKaqnDSC988jDdHOFwe5wJN3
HBa9zD8mc9XgKSxwOSkNCwzLyPlxqfNki7VJM30cjM8nIzEwXQHKIfMvGnhv4gynw54mGx1hg9G+
VuWeUy1mFVYet9FHmwio5B0eiEZPpCdl4saU+1SbpbTsvk25p5Sp6lVjPALh65mieTJkBkQ7jS/4
yTXHFX91dDSwjm8sqvka5DtnOvxJD2DHjWyGQjfuUU7+Bzu31rjRAH7Zp6bEUeX2/DtsO+ZxwARn
yzZwmaU+WU1tj7ILBdIRVaOTR8Cn9Koz/mq53fWtzJQgYVSvHvO2TYqeT0aGGUJMx6F5fooAWgom
WW6xkw+CLc/aQ1FZymQ76kfpQ/HQhyg2sabSLIZFhcOxRD0BEaqFAvHJQ1G0H63A0HE3Qnw04LME
sQUzX6Ru+fO1+VxA4YqunSWoCGG/PjESRVOLUeUYWbDqFTg1Eq/vM4kG+LlVY1amsSpPQPpG40In
KgqNi7L3x4WLgllSnIkQxsTLzL5kj2UVUjsbkInJ7be2Gb1jQpsLj3eX22gr4BheryV+KhaP6yjk
or1q5ovqqRRDWW6vhuKw06S0Ka3PpswWlOJkuqgVBuAE0BbT1GvxoXWrleAleoJcBkru9OUV9rNV
dRFKY/SNE5T/dTLZ+T1fbcX66BlnyO1qvJJJN0PFIkH2SMfxbP5XerN3cxDEmJnBpdvkjLZuVLCr
2U9NE41UF7dI7j2cjdFOZLuBumnsEo2rWZYvmURnwNC11Na2YetsROLuQlAYo7E3b362vofulP/F
aFqB+3N9EHZjgrFkOM1z7QXt6jYK0kHQDaatkhUfVw0bJ/mssi/R+4gVJYfl0CfiYYYDqDoG2B5j
iMqsv+oKb+f8JaociXvgAu6kb/HZj7LwfPUI3MPvN9OwkiRVR7SsSEyBgabEA6gwsovYl74t/zK8
HLqKf0J+9opCQok8o0157Oogfpj3wgU9ZFsHJcVoD8S9x7xBJ3HtptNUI4ess5xrO9Jod2at51/z
jRZVq6hXyMIQ16WWFlASXfi0dVbTtP+LRlGWOlj+rKjGflgQ73UI3MRdT/NeBT7OD523mbPLRJQR
NToQMAzJEHT6RAA7vH3FYpk3b6JAwuMnunEstpoEHWHkQubLVShCfXlMdFZBJNbh92nQeXUzGxuJ
odV4O9kO/nxeP9kupBzWC8bxCCRA8CxX7GF/APgfF1jQ77QV/1wortoVVOMBjis6I97x/t7EZ7mW
2KhwOUEnTLZintH58FPvGd9yEr4AyMmJEiQpRR62ij/419/OIxx3qivbzSpK1alU5tNXQcVDLaDp
Eua2Pn3vCtKBdQMMIsPNTCQmox6YvverxZnyyNMBejUulLIfydHE0RKwRWUoMK8O8MjOU5kXOl55
9/gF7fGVgEDjVux5PWHG5hoeHXc2V+DrSZvVIDw/dn2EoxZNdvBfaSlI8pro3XfFMPSV6CjTXXeS
YG/c6omn2CvOhh/+fYfjNRcfVXlB23PnGx5WiNZ9Cfcq97h5JYLDjyQIBiZGMTgiAiaEjIQAcyUo
1RCw6R+kSei+ZDmc+ZAN6cRxx9LSx8Oa/QqafFEqFBKed41iGSWAWq1TuHwsPcjayuoCsYFnvmoq
nPfmry+DJfCwDPPQWufD6VTZW+nw+heyXHnzLBXT14CfPML+vRW//Xe1nY2wfIrHr76/u1RRt9WI
JOrUXjUffFXGwium0QKbHNz8FZ2Pz7Mss8NF1M7IWeJnj3EK+S7lJghJjJHDZcq+M0Tely8lJwp4
DO4YsLUXSnEQ0tz4szNBGwrsuxVPDOgwbtpMXokkyxxlwA48n7ikWeohlR4ZvuRnPbol0F0SdXBj
6xwWjLIXB+qD16WVVzudmSgSWNZ2k0qMel8GnpEsOynyMi6whpSvlR3bawZgwLj2nvmTx7AYknkx
ngsBLg0ybmVXTEFDux5/kaZkt8PMXaMdiLHIGxFYgEgODNwTmxS1VulletdCUjZLG50/qqSeQiM4
qZNd/8qGO6KzLPHeIZWOcs946f8aV9btdnTE74dmP27DncdxpOD3/l1FW9u6pSY8sEhmaJIzWwLW
9lkY1IhLDcAYebshdWlL5+Vn/HsPXDO5Gr8P70fsSEcwkYA2uYsjR0KjykBSWFQK6K8xMzsBg9dM
LvkIGXCE2QQpZeYCVzFHzid/c5+W1X12Iu8xGKJRKn25u0FZLVXbjzeOAEdVvgHngqImp1XZpVgP
6bC9Rp0vAx+6onTg+UEvYABVZlvHIpqBXuw+jb+nvSujJ1KgRtMgnZ5V3Uq4zDuYvQr4thBD7n99
dCEJlHhYcXIpip7WcMYx+V0H5Om9sHYEp8hT7SrMELOnuYzqAuvemloU2PSFVWHE+UOZk9OHtoZl
Pn4Pv8QH9z3C0HDh1xMPE2QerbFKBXu8akza+rYSmaSY2o6PmiPjxFzsZ1th1fMNZz21h6zovdwg
Ip+gesPa+IXvJBpMMJBWNQ2Oaz+UL9medjKsM8kpDJuNmlFL1SUHEEMT+3P0A0gME6F3/uIUu4zr
2eLixSos+R0adSAdvA5IORYAe2Op95+v/EYaVpQhvYEm63KS5VgmwIBY2Bfm+7JiYb7eug4Rz5C6
DUDvGQeU5tnulv6Jk+fIzO7WaKmfVFGfIk81My/TPxAqs/ZTl5d/lx6V33GUQq/JVd0qkUEslh35
dsnCNaXEezc44kJQ2HyIiqXUTw4ZvE8vtUVBwpjbdhQuPTFGiaVt79RTl4hHrJxGwS0ilrAKUCLt
VqD3s0Lgoe74NbschicDuctOkip0zo6reMUv7xMSD/p1+bqxL9+dU3FvVnnXmrsFCYDNg0BOhh9e
Ce5hp0JovlpaEpTmG4/1yeNrVuxt9M3m0ip3ACaPf/V52oN0lv6m7d9zwwOMcl++yf3u6+Aj2k+Y
W6ZEy7GWHsOKgtvjs0pISH0Qdo5ARBFfwcOgEFDkzdpYnsAboFj0ro3uIojzolJZcRcntukSHzCH
B545PJ5/PneOpjOtNE7HtvmkLM8MMWtoAexIZXnI+kZYFrZd/qmestxBFfTlzkWtQdlLeu/CPfje
6VQxSnOuYCkhEGC4SQWiwAM7s5jc26myfMaYMf6R9Us7Ar88Rhx//4vzcOvt3/f7Pww5dZ2GlOO7
B/px7SCRat73HXeJ8mcHkvDRFhRHibsMcbTN6rGQgP24MdbxuN4BhUddk673ydvArQCjw155QirE
fRhaJ8yNoFZ73awVMFaWIEBh7CHcNUXnfuJT0iMuGkmDwccFW8Lx1WI7q2xIeFhgQAMGzuxIGL4s
BbF3pJ13EdjjEkm/xkhJGahBSaBplO+qUL/CsRuJiA/HnaaZXDT/8nZ+QgrBQQGTtoHH0lVKiT8Q
GStPfkIdUSQ28o0yHpYybXDBcsRxkYQwTAniASed52keCL9uywnasc7XcYLBP5wflnEWc8/fqUGI
FJx3V2Iybl0T/Gxh8PGeXtuGoVRowHDhH5UByDKbdpMM5iDrCxvAPLoeWU9PtRl3PUO3rd+pbALM
Def92wLNukK70GKdTmMiwDEbfpljI5oU+baZdNHYkunerAVGuj0vWH78TqntbRBBAZyfJJaEFbT8
0qwJx3eAOaJdBJMWZiZ8zCRYtEKxPwKwRxuMiONifXSCMbYwDQVk12JpDaP0rQXmFASfe9zYIs4v
8mgJtaiU8sktU8cHpd8vT10XdO91zjwdisPGM7lUWuV1NAhua8WDz6DcnN+880bk8IaJjh7+nBNM
mqiKnEQBTWjgDNWBlJEcXa0nx/CX+1UkYfK7p4Pu9k0D98oy6dqSErHIqlyrbYy9XytRAKB+tQ2H
yle/zJWNkdQcAT5WTDeRPUZ/ZWHHqRnRnYaDblluX3LkZLHTNeWJfNufoWJKuuqwX7VUrW2FyoUK
rk5O7JAThe0w2y1a/lcmAIXI3Wj9vvNmfKMTNXy9aujMNilKd5HuTlRCebJert7Ssw1rXc3V6Qj8
TDXUA39El43Bjd0qgjgJFrn1SFRyyggTUm/N0bDCbx52fsawgCuSmKGpcMxd9HLAbROi3l/+dsak
oGY0gZN3W88cRQ5hY6HzLagpDIJTCX0qASyk/dRezChngTHqkFjh4Oc5tOz+UU3WdJ1Ju58WquLa
YCt5cgHot+3Zmin8baIj/AU1gvshkLcb9ECo/UNZrc3+VSdwTm/HirEw7kWJqxdXnAvGBRnyu6yZ
KjBctvYBdb/bQ+kpA3VcPRkVHq5ek0Ng26BGodfz3v7ULzluPkId7c2o1GYRncMSa/is8LCpqUFm
4h0JARghoU4Q8xH5qnDXz9NXgwi57OinS0mU0sTF63X+KWi3EnJFq/wUK4End+1llCS78lhyzXkN
AuWyhYDJLdIr3tKelGA6KNdGlKdaiKuvTIgJGnF4uyEkHNnUTi0Ggxe4OdcJciHPjNoEs/napMXZ
UL/YTlMLuiq4YKGIdX7gjbVp6MVR7qHSTlqiJE+RTCfBapVRfGO/tp4fUeV0/toVzJfbRCtixnDv
Q/IsN7Ifk+oVG0TEwr5tlK11b/Q+dsP2a3yJltqbI+nQqu9K3zG9edg1DkFEsJsP8pnxj04jk77e
cqDz21NZGrkbjjYtOa47Iu0+R74uLXS3zx9O+6XU6oewHg+Ro+Ws5WWIiUgR6sEqK5/jQa005k20
aGhaC8GfvBHLaghAgnItQHzqcx9VnovEzAC2kXl5x/KAIWI0xwXeOT4dCg17RQ6GGqkaf2DVYGRJ
VeKB2GmUKIIrExROeX0x5xFUGcJxjIP+LE46BIIuxae0McEnPbmB5KwzBiuu+znQyWx84K1L+2mm
wXMKVt4CCcjczZqi8zP5zrEUbDcTz76VTLk3AT6ml7Ci2g7QxKZshJuC0IGUI2KJ2DSOdnns9Bs1
4DV4cOhujENEDtWHD9v2NjXlwdKQrvmMHx8a/aShlAFoiXAh9Bdh6SipDdVOmeugOzTaAQC2whFF
SzYhA1MRZm3Eg7XfgXuv4uBqUX2Sx8Sik0unf5QhJpuqVGGDkxryWopQBkj9j7/jLf0vANEKVNDW
ObWiYLqP2QTg1V1H68YDIAkS7HF2LrvWKDUxmzW0giVuSv+MNeLcB8OtBVpikr1ErTMbRdvpXaIr
StQ8Nyf4ScimrsPQXa1YHj0DgZNQ/4IX+zhAnBRJCweaKKW2YXEuVagpdDg7mgUSKjF6yUcYz3XV
GhnLbde46B6eQNbdvgVUME0419weZK6wSSOfOHAswTTqhK+MozVUhm6jke4TK7wbf2APpWgadM1L
7Ogz/yOQclgdeWD39aCLJbvLeFary1vpPQKb2VxL5Bc0l9j+BXJ0wklRrx52xq3vTDxzLIBWOa2P
ad7DLUOPKGx4CKo3p7mURhbhjgdEpDdynWvgKV2eKFItprf46PJ0GhoKlO7tS/n2uDLqaiGEQlCu
cqiyY7jjbNlN8MtIyQH/BBa9NEKJru/xs5MpFFaR8grGKtGxmPi2NndC6K9INdSwZBlka1ex6k2K
CRsncSt85LzSbMQ+YreIP0XabJOnLJA4RnKGgeDnEWUhtauuIkWdJ9AOU3l3p7u81NwvX1uG9xZU
JFsw0ZVqsNC5Tnse6imr3hwqQKTVd4gxNixRUiUIDOmjjw9/wcj1SOI8xOc7VXpeQ/x46y63yCbo
RSN3al7em6VI3X9qfuT6mNQgkAKWDvd2TzdMWUrqls9szeejdKUU5o0TvbV0aGWyQ4rkD70KRPqk
1D0U8SNSkejniLcPt7VJ9AJvJGWMgkqj/u4yDDYu8sdUDuNc+dowh+0FYxyQBh7jt+Ucx5tdCOoX
kr6pUiD955BNzZh971JTG0KudBBOIpanHBLa1aRJ4d9oiYcRwMD9Rmhx94VlpFVkcs30hXehu9vP
9iiBSkcCqJNtTqdEJv0dO5yU626qGmFki9MMzcynrf/qXQ6NsrY0NJpRrInbMCyqVmKb2/9JtfCn
RhrCGY18hyItfb+Ag/th1jBd3XXbzlnX6dszdZ6t8VW5FvK4qjbumcos+9DLdLPpGwEDPsMXGOFU
CxmVUtYzdd2u8Bt5WgAlZ7zlKFDFnBU1n2XDVcKnbakeXI+Nb9dkuIArleQZgjuoXxhpyomupr0B
FSWI9yb5y9TSD35czwSUcdjwbXoR5kgtUZPb6pmyFZNaVSfqDsSXbdBuGNaaVXYn/2P6a3XWZzZr
9GCd0BEo1hgk9LJoLbPoj5lPVDWe0yMzG3OK5pR4Ig5IPLV/vFMIqz7oBmLg0j1gRx47xiB/Ion6
ko3gpYnveTwwVmASAwKuevwBAMTXaXmtymRbssOznnk8FjKwBjf44fc5ferSjidL6p0uuWx9D3CJ
x8rlZUN2ho8wWm+lm7P5Eq7hEC8WRGUs5kbE7bQLUJo74840UJcM0ZvHHhyo6YYLd3Wj4SoNXnIM
f9bWV1c0vCS51TgUPfqsmquH9r2MapjCTgf8O2dPpbOcfHBj51XrdtaxlQyvaaj/Ts6QVcQe0xqL
VGSb8OhemQAhiYblzI0dYiwH9q3rlphuRkUzx4Kkiju71Ylew25MleXFAG2Fg/SLaibrC7IFJ4Ub
9nDRCAdtjzRke5Zy/Wu4bh7yh6sf5wEKStrExnCYoUINsO6ftiMBGbDbW0LV/CxUOOfEWu7YN5Op
U82i3rf5u8ClDuJ3tBRPYSqxGzOMxzLlnlYBZkTCcALw0syVqc04PSY/CukNYPJ8NT+clDKM6Dog
qaC8R6xJ8jVL7GV+mF6NvsCtPZji9woNM2ueJozJ8g01ks4rNAEVF3vfB7xhsU7n/NOiXUY92CKe
1cpza0sPeZbJi6PZ5qb6I5+mqU95JIUP/5ciQkdr5OQvPfI6TR1jAUfAM0JcZ+4luSBtk+iCGexs
BqThgstQWDlqWh3iy8uqKAjQ7pL6+rni1kkOCPMHIpGmUcBDZLJhnpzMRi+twNreflJwlbbq/rwV
YDng6q0S7rJtmoPZB+jolFxKA8FZj+AMA8kxlFtjS7PrO1RK8oriiXPW4fPQV0YvnBfKooKbExJw
OOwHRnE6d4UZSZa0eGTEue/3AePCDFiMe8eIU3Ja6W6mLDgrFv2o4A2BHQu5+WLzstyPXCwhBs91
1u3OlzsQYvHwjG8Z5Hg6ipYZ6ZErwMyY9Dn2BWlgbE6asjDyfe4UMAB7PCZbEd7XftunGMpxOUcc
Wv1KOw18Cpg46kbiDvDAh4pKG1eGCtWfh8Ju6ABdEweNyiviQ6wbQKrm8EkzuTs5F+6xJpo9SGMT
fXNZzKPIPGHgtQv5frh9qP3MEvmgGoDGDcTOyqAoflqYEDnR1H+y5geOlbCdO3cPXqtDYCA7B77L
V2Vcuo93virpMgwxlF6n5kUf4pvtDBBFZCq0M94/EyNnLaCepmTz9fmCfGOOWS0+Rs3u3e+Z1Y42
eQtDIkFxjlyiZubJocaOCXSPeQNtQsjjArfkp2iQhRGIP7MmACu8jXW8Oe8bZV13k/wDI46eZ9M3
GJD+HlwbgPmaGZH1wZ7BTw5PrjMneuO3pQXbsyLltih02Q7mavgbz+TdZzUwhyYp4XSSaS7QVhF3
cT3dlMzI8sFYiOpTY0ifWWmO6Qzbjq2Seihb2m5GQRgJZn6JPzsta1irsratsxiDaLI4vSApRMYN
rCIkZz0uKsZV4gmiZRInMu8paeAo1I/WPeqM9PenCoNX7Rauj2GsLoWDxKDoBcjZZ6qEB4elFb6L
CZxDtF/dpTgE1/1Vewb8LrLulipetgPwnsIkbmUrq2Pcos9YAvu2qNyElTA7RmcM+Ad/6PIO3MAE
MvEtJFd37qRiJ/DnjPJiDXrmkjx2cxX29q6zPz+amKhOIoESqwnTe2ngLpjekODcpaP5U5aiOcmG
v3IaVrDstzLtGCo8NTilq0ukIbUlt32+PH3eQhQalne0JH8r3KG39c75cfzGcqyCXudnXihs8l53
krGUswqFqrPFn12M18xZQq7/kp9aT60dZoN0MU2+EWJkvb/f63zNVtAkIGdCnjsAfjrBhEDxpwZx
WDF7AjRJrJsQHCIdNhap749b0I49gPxAF0rr0YLc9KpvdVF3OWXlyWAwb+sxYpA+Z7nXVHxxhkNr
8IBhwnFt+vBewjWSEMhD5YoO56m2Bt5s+KOTgv9OmnxxRbzS9XDLKltUarsxAkQc8M75vy412XIQ
zlVxbks9SLBeXQcxKlY8uBbVCyrF+d7Mclgb92P978mJ5mprl0azdrxjEmDaPPGK75d+w/HN/Cqr
1+8PWrySc9Fl5CaNzo+k6W/Esn9Mqyr3zXJEm5+T31TBD06NvwW92cl4+P+bNJ9t82zcB9VaaDQW
vRkMH+UHa+AvwTy6dd270MQ/vWsZHKdPsZS/LF8KJLbdrFCQJUFCYrFjcy0l+6lwfPJoU+Kb8adr
nnuIX6BfyiGYxJe0jFcg99oEFcAitlw/15vRPd50VoeBYbbLFTKL8xHMy3Md1AOKHwT824ZiQkIL
pp0SDG5qepyo1l4MPoeTWShqxc8uZWckDcdH6DQbi7h7PcBNIfh8/73+rEEdv3EYnz+vMdhtltXJ
4XTRKi/KUmy9qA0+6b8fvH7SJWmAQlX/yBgIYEa2ru8wVIVIADHAGK2RNMV2VGCrRrdBbK4zRE4k
XIbJF6v++Fnz+BgSpRseQTO3WdbxXBf3MAkdf4lBneBoSKzVfwWSOEazQiB3m2kTR7tQ351iS2e8
m+HwBrPKdLtHMwYmkAp5WpAhq/3fsmxOufwyCQw24YJVmE/EfiVk9HPp2UzL1oO2h/lLUU3e5D9O
8mMySkJ0ruK1Ve0K8HbU6Yufr2rV6FSaK6Rl13LWmvUfn7Yt6myFwgvYUtmEakyuBFxzoeI/K7lS
uhUoqnBRsIGgVvmPdaq6DTJLWSCAiW/Yhap2mwO/arzLWvFzrELnl70G4XWqJ/J0NERiqL0Pefif
YsxRra623YuX0+dv9rKoI5rxDZ6FORWKxorATHDaGNY92ipK0GkBHTDVL9ihyazJ4zaXQ4h8i4LP
cR8Lp8MJpppUhLOwe75hgmJwdln6dqXjDK4JSU/UcCJqeldVmZaCtu/Qpj/4JcwBxIuxEsA+VZXx
gRW/dXVsObUjukRNSPrv2K6BXxyLtESdLxp32BBILcTCC88/IzAgrtCDk5CqoE/2V2X9Ag5PlUTz
GeZEH5txmgmJl0FUvrXeWIhX43bcGYtwHp7LNueC1FGWc0u6+9xZ7wRZh9fuomffQeGwnDYCR1q/
S+jWydNGeTVOsWlxARBRD8yFwPNvzudqyb92zgbMACwKCaXVEfpfHIcRR4oLQWimPjUKWtYR2AVN
x8Dsu8UDlY22XM7/bJI9eXb49JhnPdkl/KNBEosBbPZj9+PmTl1AKL3y6Qsr1zI8e5UWbhmH7hjq
0hCzCUlyr1PRHFOVLrAg1879VMlB3G0yGr8CdVAuWuxBm9OjhjyrzEFPALHyegU8KN/J3TNw+kgv
rhcntv1sANWQOgE+dx96Yn6b+PQRfAOlko8Im5aXZjEfwPhht3tNfbCJAV9AEzN9t0LNVjZX19zu
ctGAeb8c1Uw2gVgJYqa/W4k5wDAnXjZ2ByNj+HID72qHq/0q4vHxY1S622Tcsd5KxyeLMP8Ce20c
h8W9qIG+sjkABq6qX5cxVp+cvj0hfdJMpRmBaqfZIghsJl/RSp9TLnBWRVi3WNM4i2DQRwz2bFme
1wHnDrKFyFQm1BtxlxrcTa71/tyVkq5r2zEjyFne0+IRVzveCl3Pfn03Mkob8EWt7F2MfHmLA0nb
uNKpjlrFgSdtHt9P+Jp9gtRXu7MqaeyUXd732clR9CFFO9KkpoX5/iBrWmOpyCyJdTh49K2DzJVn
3QMTABGGklZVgOwt9AlvlD6Rn/RKnNrQhRX/02Cfwg1mWXaHqQZzHVZ9YHYv77ZlC2Gaok5cxnpx
II0i2Vo9QLkxuzst508gfCeHdg+kMMsTb0i/AN2OVPCf/i/1wu4bvK7WvZowK175nZF/FGtrjSaf
n9H/2TRp//VdWW0FBGsiRvVaashRfqnRXZiRea3IVykxESK/JjakcVEQhrYFZOtSQAfxeJIguwBG
BbbyEs87nB5rOR9ZTRBZj3AdiWZMjZSyuHk2WxovoIleoQ0fnHdHTcPjiKesXjwUJHLmrObLIiZV
kWqW3QUAkxch/JKMBd3MHOSXGatzH3cmfYWqlkRoCwQByn/ULFnX4UFxeyxbn7CCYuqYGUV8o7oP
1OQAihaHzTc+frAgUimiG94XGuGKMeRiK+IIk4ZQzUcC+ndEJJz1bRAy8lviaGrqr0/J0YkuDU5V
P8WlT6dBkSiZqvelpAg0xkSgQEnHkpTurTZLs/VLV4MmccvDklm08yd0QcogRv1G7a9C/wxh2Ig1
usRE6zFLSVD8YxjxxgSN2LB/HfGdxvzHY1e0ydRU3AZVt6QykOkPhhqHUmkqC2/jvfN3g82OZC2M
u8IaQwSWY/EH5IT0z1SrVK33QUZBtfw6yEtA3XlCz4+UyxkJ/M4CRrWRIQA03lBGZl/Sgejg0GbS
83VI8aj8FmJOHdbke5oHShaFINd/6NjSSQLFi6CNSQKB4LM66w3JCM2nreqDpVUrGZxkPg0pKS3D
9adhWy/ruzquM1TQys1FfKuY38alFewhWvrawiWg/5QmzcyRSmwXdXSxZzD/qT/G5x50gw52wA/L
cyaA2kdelrDRBH+yfrBVYheEe2ZNE/f7h2tKWkjIxgUarL2VKkRPOvnfOT1Ol0y81E83zChVxIoj
HNsBqfIceEb2OhgvO5yofqGaKZ+CifCDnHMAi54saNI8vnyuTlPGvT3V7IyXG3Zh/cDheTqLBIw7
J0SH71dMPnikRd+Mb7ZqyE9B9JzDKo6oTJCvene1o8DtwemWnf2a1053ScASsnAAmW9s7JFVs3B6
NsukGJHYGhWuS+epnKfXt7t1OI9ThRctqn9U7/lz85nkMr8W3OZUykTEeb/H8BkQGEUSz8Pr6obT
5+7ibJXPQ4qBv0xtYlB+VBtpJEyGi66b3VivlanqzC3nDsPbF9Ul+Jqt3CblS199hf9peKuxK3Kb
kJFalsGB7f4+VM5ZfsIO+arSKNVDAw2ijkJcy3bvRvNIK48B1w9yL3NEmtm4KtkC5FTtBkfk3LxN
EUd2W5t2eCLU/pFzhmT360675cS8C2IKo2SNg+ARK2e1ZeZvHm0g1yRQ2vyMvacxW0uF5ooIO4Nw
cSqKs1ZfGBJs8V8tNuV8f2k4pefRSqagXb0WLePOi/m+rv8OyxWXCp0IxzpMq1+Nq00y4ZFCzcBo
GWHx87iqt5kK+tmSeufJrLES8pXfqOaMxom/S1ByQ0788zhDsUVgYDVNY0DsNFQr6AYgz7bMYSOY
bJlYJaavcbu3xi/dRIC2jFYp/Qrv3A+OqL9NJmA9wRjkrKrJqS1BJJPEqWomnpH5HpSR7Nr1DNnN
HMItrAvCD42cSvZmIIBBnxan6PtzSftqcupaQiILUxcaIqsBIg4jy1tbkfQpZUCnxdmb0ud+7dMt
gpv8Pjhj6Gl+l1cUgQL9e03NUAgKrDqAShYo2X9TA8dfDQr8eKC73bX0itC7F0FKGIx4s8UyjsBG
IGjThWIizICO2VGPQcfqNQzS/A0iGJLNAoJ0abSdn5kmi68EDMR2Nwu1i4qLmhwYa1iTEMI5j/vY
hg+K8eTFx81D3fn1mK9257RJiUuJWVuPMDP40iexSrW+e+FYoJpd1Vs/TyIFKH0Yeyvhe8pFmERL
lSYELaWWy+QjaZM3OIj7rhREWWLi+oRz5kZDB4w6bO9s2JfL6KZNhUD6M6TyxwWkc0f2TOb+GWsE
CMWgPbZOoTGCj24Ylm96vzEIO3OWZ/vmNUUjV4LWRfoM2DOj0QAwa7kfRD7nCQJ3DvOfJkmAKq69
oszPB8cXVjIqrr90b1jvhXLljONAmlDMQrkfhdHfR0Bet4FrkbJa8TdR2I6wBs2qmytdK8/S+6/b
0f5Ls/cR+pZWOEeQc9konqZEiqwCOGrSGKWhbDm1MEEXGuiKv0vVlHYGr3K4wDaRW8/JULL/bR2C
zzDMxglmiUySmBbzV2Sh4uAKHJhjzKLUYM5VNS5yPTspEH7XO40yO+8ZWyRVR+rVvqMPCKuBr9LO
aIZaYlq4c94jiJ0aJohGvILXVsuQozH+tWLxB4p+Q1F6msVMkPaHhZSC8ILu9ZZ/HeEI8Ca4EoUK
Se1ZFftU3UKYwV95qb0XuB2wFNQwOSAUVARXYzxlI67HfsOkpAFc8WU+zgvqjblO0nCXkY8VI6AG
ITQtO21gI7hY1SlRYB4vCsb7brxk/BCTeOZC2WjioTdHu09rq31TW98nyKR4Dar/t6+RvPb1Azvb
sMGfQ8ap2BjZX/RhJeTYgH+3Rv2FvdkptKOjhme31VX5K87waljppqQKPrUY/rDdU2JkdyGbxkFO
XI1JDUioy0dTR2q+jPTZcZ+PjicjXphAj6HGS+gz4qWi7G/hFQjrmITapfBx+Unje+pbU3FJk5J8
wUy+Z06z86Hphs8j+lQhV5YFaDVUrolMn8Pht9ExOnpeqQgi0jBbRLPBPk3TdZNSOPnJiKvzNNB8
kf4uMxUDCw/1UaGT1wYZJXAlWJo2FS0k5LlYVDpEoLIeIEVSSV2qNt66bh4pOzCdjv57G0VHHBvo
AEjUb7qIlCkBvp8oQJVPiZW1qeyjJBiIQ2zMGwCUbWeFDia9dnmYvvtg1aeAZmnSYtQI0Qw0be8P
Cl7L0iPcOKCojlbJFvKmwbdwvEqeqOKb0FcKfVMNARVDwI+yVnXvldsFadGOEPfIYQRlzoKw6xll
D5teG97MNAv1upAT2lg5WZzZu4Bvc+RF+zJio02Si0mrvwbNhOOUrq4fF4gPtExGJPw4YcvNKEr6
A3WsGaGCtqjqmnBwCu9CiJbeXKJLvYzcqmPo6d/CY1vRnGieMCFq9jha3+RChUjFg10zx9tNejKI
nZDVOQCXbJVmt1ypkGaSrnwtXcBcemg/jvD4qR606EpzuhJIOiWeJ043xLVUFpOF1KYJjIdOGasc
ZXL7fXQyXMywSZPz1u2nqANmkyq3pP34HDpK/bizxdTEAyOr0zPfsfpRtsCAiLsa9KJgYZ0l1j99
Pr+l4yBNIZLPERlrs2THIRV88Zy/ggUqabWXBIuD13xVmT6PHpWfQrB3S9CRfRx37Q264152kl4A
oYWlZYBVdm9y9D1Hp87F4FQ+tyRkVxy9WWQE2z3XYHulOObF7zaB/ePj2u6RzbWuUK9pNoAUwFoH
mG5ennqlii5XxCXczWDT584HHEDLVvwZtkkRqPQx6DUgvhmMniXKKlQrhzy758BFoBTAR6a9BZNz
+KocpreAJBxmQ8ORk2T9iknzW6r1ogVbx9+PpKE1Je1DXCZZtW4zlf11+gCO2vB3/hBsksN+kM9+
QZjPNYWlgWN1T/flklLe9my/ylS31dmh/SugyHKv0GYR+qsoQYVgwB1arHdK0yjvB/ycq5AejzNO
w5xGrRycHQ8Tz6XQ1iwjHaW6wVk+/16LdCERF8SdyaJNJqqMcBVpZdQQRy/lbEADOi/i+v0bKx/3
g9ZuAONdBkzeJHkYtdrHcFv+fKTPIbkjOMm17KTCqUMdcbqOMVlfEsyqGVtrkbcmgEawU9GL1wlK
WAYggjcJZTnbdHVCdQUI0foOYDKn0+talUd0boev2MFWkhG6kPU9Ud0eJg8J4pjwJCk/qDA5jXoj
mI4CgLUdvNayuUfsV65jYpLrxt8G6AnThz7stwv0dTISpjcveWPOiDkqtvvJKVHZ6rcSat1PKrag
Gn7sFTSC2ZwDFreCHmKwtCKPhWk9uwHXdfIp9zAfD+oFdHTiK2TwKeW3/p5U3e7Ty1bMqIg5aiKr
KJsGJTudr/NoNFHjThISY8vBSbFqkCcVbG834ATzgC+Yn95UaoSEFNKTWI9wg9GE6HQXj2j9ZYXH
OGoYHPJnPhhQEHp4WN8GKJses/ZTMmUGAJHHWiWEuwpVeKm8xi5xqgnm29eJM7j7aGwkS3BKQPDI
H0elYyYiehm0IvgfKiBydxkVTNDmALo3Jo1yAX2K0H/Kji8qt4EPLsGH+Cg/Qvr6e+fnDxEtUbnf
v49WrtHO19adWkks95crZHcKeFWHXUx47L6x4h7WTtgoI2woklwuetfYLFvx8S+PYldEmWHPKBls
WSOYn4qmlUhZATUySzTlN3i+u3xbxlkan5sC1MbRFWPUTWi5OSSoHtiEoRD1oNsQ6HRVSLQrp87G
F4ZnzHLjbnDGZJnlTr8LUSoSojQZJflB7i8UMixXiA1pEpNyx4iCLPuj2ldZw5FriEHa3fOYTKPt
7i8KNGwW51AT3mbw8Nhf+mqI9vxWmzClyVuo2ceHAU1XRiV3D4/WEgG1TZ7eJfOu6nONkjBn/p2H
yVJB3Kn1iytgFoszgnFbZTgw8Qpns8cGX8UwJbyPBJF22PSC2RFjgP8t6uCSEkGTCu0rZTTrx3YR
fYT31mAxW3AnioclIjJ9xGkhXXQMv2LnQljpCPnanqldEWCC4ixwUZJHpi47i6H6Ydmtaxlb34wa
kxRmwhCdna8wbhxMMl2+M1gBG7YuK4OADw/LePfoWGAYv8ncZeKHcio8i52SrxwUfbg8clITLQGp
qWa5dj5kKllDWUyrD27dYMIzUrxlOoXhRF6+MgnE16/sJcGH9YfzYf7qF51MqOfPtL31e1SE9eZe
wfat1YnStPL8rfI8UUr7XDgfcFdO0jvFgUTZ9mHeF+fBCLNJb3s38ZYnx8uh1Qa0ikFTYQu5fQIM
9C5EGU273sDSUVifj8zR3rZimf2OtdGKMeCBZydlyffx/oSbD6RAUpmjct3hQu/WqcHy2bChcg60
KQZABuocwDGV3xfQVcWx2y3fiadbSF2jGuPFfn7Rep3TTdZqGZE6Lqxf4wAjeILwG6JWpoKEmDHp
K0M0YNEa44UIjHKiSta3ffXe1MvDUa01BccvxOQZKjT8XltgKisP6yxrL9qL4FHg5H+UBV/+Y2xC
448mQuqMR8fov3ddHJNRGLylahZ6qfdeVWKKXxGbpRd5CZUcgb9eB1oT1fhx9pCtTqpafzl70WLc
pBl0JdU9P6tEHlyYPDoWX/Ke9U1YKVCKjoNgA/at43V5sPHDHotrjwmbjJlPPMCK/juO6hCiUDIL
pQbhuATVZXgWppKQds2bfJgs1crY+n0unZAZaWkw6f0B45u+T8cmwunUcC/rkYahVm7NGoBbe9ma
NA4bK3rWOugBCjLZfB7kpIzDDCrucrI25fjrOyOYugKu+dGJReohliPbDz7GJEXUx88xJHrt9d02
aqfOeSNZRWeArx9ax4aN98fH0RF8aea+30XmKObZXceZfsHhVhk4QkGQwjpU1mh8fRx83UltxbVB
eLmk3/yonpcm9I1fdfIkZAdooXfoKoDip5TZZOtYB8j+dYUAihOm27ZZLRgMWzsrpv9OT2qAAojS
2AXCF2/3uH/iB54e0ZgONAxoVGFKTIPm/3b8lG0fgD/ialFCAN5lHqcfZARMU4oFoL8qfGCSUeaa
dunjg4OTHeaK6x1UP+cqElgcq/SPyXduM0zeGvWgAJ8H9ORBZNoeDVcfFJmzvwqN2VvgI77oUoFn
uTW/4z60h09nCctd3XFiYghpebOgOhukG+RaEIxkDptsriMJT4DGHJpqwE1bQUlLqxszKzsx4dDO
tHVOttBZMqjINnU175BwZA++2kyXlnqO2B3/nnYfVvUkYbL3ZdFHCt0AHLkKkYD/gtPymuQ8cOS3
/dcPFZpUGs6ScDPmuDY5JSWzV9JORw3SE7OJz1iMK9TBthqFkp7Uj8EDGMU6basqRKO3umgK4wF5
kmkWtq0S6hympU2xUdYk50tBZHFr3pkQ+fp5YqQS1nHRkyF7vDcFdRASpy6c/h/Ry7OnniBSQLwY
AWeVKCrPsK8yLqhzQrwhtS+EWTBgY5azKBLyJP4GfrXuNeJlg2NS/97YTMx+6Rf5OPP6eFHD+q5s
pi+VGHM/5FSvw9ptTSVg82WniN77ymLx1SDc0Jk2DNKsUeDKeyCp00mWKACYZe9DwPBv1aZl/7Xm
55o32TM6HB8c0Xo0F4lNespgDtsrHcnZuDiZZLaOa6KwNcvjxKEs/989+7DWsgKuHEMyCPkqI2z0
M5aSSWyQAheUIUdcqtFY5bZ+auQ9qZXuKz8d3TNBe2q56vc2OFRfmLKkRvLe5+5DWR96g3nDJ0oC
3VlB2wZMIgqQhrtW7k1ep0gpiyRUtURDKHNr+XtXNsc2/BfUMS+NuyZuJDdBHCQw07TkTQFekmNa
/h2uTRs32TtgSfqioaJBeSsNecUxopttc/Mxt+sgjvR2cj2bR2cp73GIEte8eStq4UBMcTnUEOgH
Ht34ECiVrRfHYAxZslVedEAqH8+3Q+zhExZ9O/F4psU9y4Shh+T/1dnp87dONnByD9o0HT/kE++g
wrWY8BQ634XnMnA/o44+W9ucp4IkcZkmfvleC8CbWMMR3V+MlFa8NlcSTRqNKr+Q4EeKzvbAWAVZ
4iirp7Va9rFe9L5yB/TS8RElB82uAjV5OY/A0PnvpHLHTVW+/QStf3+h3SkVESxwDt7t624zqFUc
tk3TXXu+sJ4DvtIqWy5UjhfTapWpE9+O+3X5SLbSc21sI3/UJqLUzrcPD+BTveXsAeTsCsHOBwFU
NwM5j5LPpxVEbXBMQnQ96tsZwVFSAIrYATuyKeMIqZqHpas9p5u5r+1OUo1f9GoZdQxqNa3eiIbb
d3UXQRRjjQhLB15bPheyQDGQ2nVVzyRelxvuxYraqCud933HUetphs6i9dPYYB6owOul6Eevm9uu
wUW/uUrDmEi1KMZvEx0wLgmf/evqKYt1rMsES7ten+6hZNcV1MHTaimdRpPx1did0Pqo2h4L1v9m
mCaG4q1tPUQtj7SriboTbnSHYdTj1b9zw4Npf/hQtm7ZsW/IyGrcnuVp7Dn8MQZaK7h7rN4e5ci6
YklhgxCnyes9I93ZMUN4oDeLvnIgEzCZOhrwXnY3WCpzCII8Mh1p2seY4p9ISeF5gzQtpuD9NCi5
jgGSL6EbVBISOLYX8tG4VkVLvj3gO9BROJWtSvBGyzMqQI4p7Lanz4de0Q9+Mmljfe91VqzEKwiO
UgoXNsGdj1KR0ni9cT4dqfSf5w4oLwpG56ArduKnsdyPtSDzyFluCVbLH1DvD6IfXS407jnBuU0V
RxpEOwDKNjwcUQPJ7jPOLP1zFJQ4+WX/n26Vk5Jq/y1PmH1Qa8fukrO0c9Z+P47KfNp537YnOxKb
f+PUQqqocrXn4dY9XAnnYl4VAptavUHUJG5451eKXe6pmJcLyEkFwibHYCBiQmlPQEySayWRcA9u
RwJfLNIXgzjs0l8ScPBfasM+dDMyNs+ud0mjkcYKmmunZptQ8GUDP0Imupr6hTsil/rRBcWQ0igO
MP6S3k7t2qxwp4w+Ef5sndrfKoEzoIuAuZF3GGDxyjbMxGkMBbF8MWVZkMmyCqnsPMUliNRiX3kr
KJmN9rQsEYvfv8LTiNhdxu7yzZVnah8OfODMeg8yRC7zGFBUHXUHrbypKBBDo5TBzG5/6dJL/+h8
l32MzGfqamhdNL9t6QZRnpI+eQeBe3yiZRWxUKKSMabWRHWFPshIR75fwgnqvh/DXqKKRKfOYEts
qcJay5t74XWnqemPC+bd2VsC+FtVymVyRi6dc+iNkyHpbWzGFPJbbz2QJYhdCPWwwGqpTNhezMSr
KfW02hUpFSjUKOPHKMsSQbsXHDdVv7fMpSZ02dNBoqQWBOXIQHEhzQGHO/+1ZXguslMelmUU24lX
K3cui0WAPne75C2HtZDTFdFZ1XgMe91PaxJLPDS9k2LywEcP5rIchFd/L1gl6lXV02wfVBedx0ZF
O0zc0sgGdfHUeq+76pfyTtuXkLH1DnKWBAAJoRwKdJeWGb3PNc6iBHJ58++o+prRkHWLXaUoT9ku
zEWls+ifkdjQWb26IvAm1vX4aixvy65HXRbVO5RnmefjbChxjDUPScjVBCYLDpDT0ObHtq5YdjQZ
Nwg+igVTo93TtbG2HicBnr4BDpqHbsaFJmcyHMg1gy13nRQbbt08LsCAdOhBUOKcW6I8KwKcFsBx
WJwxbuTG5l9JAHb0thzQF4s/7NqFJxj8vUZhYCXlSgoOaaW07W9VM62dbjoATU04atjL/JRxLRBA
dvp+g8IZvSjhCtjK0sDlWeeEEBf4Am9ARBiZEPJd+T+zi+8ipDZ0nRs4fAVY5HhR4itfdwiMh0ma
9DLEuvd0TcdXSdmSBy8+FYpal5TcoTSjVz5Tv/GTuZ8Gdc0ZcxiC01R2dVBBM+mnpXJckRVnfczb
1Fg8dxvW9PkQIjlw6iSvc69BypPCNgItVMmN7FGBbdKgnP9j5sJ08mS6zCrL7lTUVN30ElYllwo0
AOvMEEpiq+erCiC+Yy3Tny7wSL6Cy2qPvLUmC9J/CMBJl8/ncik4xywEW+oLJwnSZnd2vwGVQ+83
yFg2H1Jw4XlWGgRwCNKDX+SG3qCk7L1Z6fG1CCS8s9zblbG2COQecioguOARpJ7115bUwCjVDVv7
iwjzFzErwVfZ0jWKsFS/pdgbWnkWJrKSf9EePK7voZwbUJERGy2lHziZlpB5yEelLmuhKOkeOMdN
241gJA7rNyVw+dpJfsZz8FG6CjdiLvwjRcbEAwZtaI4xfkU4KW4LJwrozciiTMdoMZEhR/jWG8lI
/lLbmRT5vOQzy514GvxinaeaL7WvzxQ4QzBs+jTr7lDrkmplJSB8FOHSKEWRh9FLPEWPWHsgJHFB
HSLPnN5laYKWx4QsK8c/CcA5DWiL8Ko2PfP7yiP69TMgAKZbNHAQ425ycFtx7uCxX9+go2w5tIGK
zncyEeWUjaDwGIqF6C02gA6wDRHbX5OWpKzZpPXQye7fgxY2df20wl9v4EF2NdoA7V+iJwLN3Srs
a2J7evjQ5zBBFgIs/nWvQSZBpqXap2bZ5ZwRj5nFQLYugeKKE6uqvZX+1TgK57rLqSJxiTXzox8D
UIoxcsdxNhrI6hsc1DXJmiM5Wn95mKXymQvun5HgsF5ttaFwxSZD2qfW425W/n9rf/mA0+iFzq4A
5EtUCaWAgMm8otmRXymvOJlshG79+EmK9ImkTfpb21LzIAIj1rfgYkPh70mWINK5HH0sjMBcwQ40
uKtu2z5X8sI7cvPNlRKl5QKrXEeG+IdppmkZYEdOEQ8ooh2m43DTe23rp9VQ2S0+mXBIRvUfiOX6
yDuxqg3ULQ7tK++hvSKYikNytSKno2SQM30orv3wPrTUc2imxAVRNKVRG+BOLMMyw9Zkrk3JlKj3
tk4pQ+XHelso80pM0XLd5fxIQALC1upY8gHkgxS0bB2hnP7A8emc7z+jjgY3O/wnZk81AknPyJDn
S4VHirEBHaj9CfEkQkmtd8kdMDRWNHfp2+WK3ytlD07O8Xbf2pvHajMq5oSFQGPTVWlIDPDTlEZx
nLtYitu5LSqI0N0bJ72/bjtqq6Wn9j5Mcvxcdj1Y1DJIVVLVJ6bHT6ORYJ+espKDh1eqYMSFUPNP
z1jFRPWDBnrV30MnrsAHRvUEddbZOKxxAN9Z3G17D5++TwC5sxBO2Oc0f7Bju/lwH9rydVGbQNpX
48H/++MHNoXp1lT9CSDx7H0mRzZyVKUK03iqvAefZklO4LWY9NBytcB1dJPEsPLe/dZqVkDOpmEt
8GVDIKwgUlq+dMsA6q5Lx6olQsfOA/Zh3lZ/6kqkuIYfCmQX8b7MTeNuE9zhlKwmRSG5t7mULwpM
DmAqijSO7O/SszQakIv4EQvKpKKFUWV0zAXJMDgrSMF/nFDQl9qX0j2DHekMj1cAvkEaX4SWdWjS
MENRCLc79FbAQD/Cn+5347kJ2cWdvuiiHzbLA6wa2v5NEwu836bWvo73x3NgQwPA6swpM0SrdoXh
HNpVd7vCRqbYjhs1IEWG94e3sm6TEuUXM8ekfHN2pxi6guqEiQkAR3j6+Qr9ah/YieNCFdvKfFEM
L5LcTZpVtuBtEyBfiYV6BIFRDHrsD9UxkiQLu0OSSELwVVezVS6b5YTkmEi3s16cfSSOVmUaxQKX
SZwuBGBX4IyxY1FMqTOUxaniDrzhJ+TK2Xu6Ave7rUqGrCDUGnfVN+lsKlIKkh/aDz32nALfT0Jz
yYtm4KNfK7hRvwGyF+yKbK6B56Gm3qu7BhMq3x9RqzhpYn4lI0xcI3F0q1axzqKhn6q7woJu0GcG
Zt/T/te7TWjhZN9/ix1NOgJjroBEPGwYl0gOzlaVxBE4aP0ekMJ+iza1DBezrCE6lHQnZnIiwKfu
XOuapToZhsLJMiwWeab0JYZEQ049gMgxbLySO2WvZd9PvbGwg9D1FdVAlRCQKz5v1aRmdu5DtCxW
PRls+T8cx7aQIkg6bkMXgAWQvltlhDsRWqB6VkQMQUgzzNjTsI4+1xr7CzWI2p0t+U1AW/4DQtV/
2mfsTYCtYOJlv1Ds5PnKEjdRpzeVuWIIeUTQyMdwRk1hDtFruqTsRpUcc3lwF6YPP6ytjAMIGOMM
3pmbDKVIz1cxlLNnWNNRCXo/cJS/50ZtEje4Tlf/P4jg9JTsVRAeeTgGchxKhDAE7vz79cBl+CdV
nU7BlF60UhyZOIzoMF//NC3qak5wN3iel96vtINeSRmG5YSifIK6GDdDC14tM5lB04ZP+f7B9k2v
UVH1O2mAbj/pf9snD0ZRueiETpFylCDKZzbQUu5bvoQqom4GmJWDjto0cGikW+zd9BFk7D7SrdBP
4mHKkdD7qrxiPByMQIFqhoSG7ghImmdHfsWT4ur3aGnpHGWCDx/ORaDheHwYLu7eL9PIZDN/nx66
t338+oFDxHGR+TGc7WlyF5nxsGF1e/ciaDofnFpyvF0qpz+Gqe36JUB5FPCrMC9s7llXsQZpj7Sz
Y1BW7DjQqr7UJSTRJWNRVoz1+VritcCOVTXmLdp8NlUiOCvPx3ihKnot/sQqKokeU2k9Y+f1wcbn
H0gDuhBs6pPBHii0OKozf6nG0CF3VXYtcd2bYTvSTGolVPnAaXTiaMl1HjZv9L5c4BlLH9vriJVu
GUH/wu7vAvU5LaP7BHQk0gAK0lJ5U5cbRH10bpvu4fYYlaW4oXyDtOjooV8PO2bES03ZEt6OaOIM
YyG76/pL4gaXTjrixiCzwhSxhh2ti1ULpdGP7Gmyaiu+Dmw4nYDHTbG1TyL4hdd2JVzCeCHvFlMY
J/qB7g13vLmiGEnOHqchKp9zC1GvrRs4bTi8y5T2bOLaDuP7JIasi7OKwhRxp/OjxcCcUujUpP0o
SAKAULGLFlKKRWZ6ZxibSXV5lM9zHwGerkna++ezdzJYy03B+cA7R6pAiSuhQ7IaLc4dK6WIC4ss
e3aM55QECgCR7qUt/YmzmY2DHWw0wXc2o6UX8ZsXL+GcZY7R3kMU0nq7z4IDT5otnESBaOAAf5JG
8n8SXUKrf7d0/7dBLmMxDCaDU+hKj8qYem7VmqbWwf75qhoQru4e/4+yN+wUiHJUMloGNIa7IA9J
4gJJWIhIndFhHcuqgoaExFqRXti4LvX27PwdDoVv4PiRCQ2uqhZJ+fT0okJXRaXb0ieUtjgXXGbs
eKA46b0hQ9lF+Sz4S7BhtUpzwvBGOH/jnWUvsIfvwDH8tReweWEKcfL4rGfW9Gl2E/BehUOdCePY
5u2dh4ItcGQ6PUEs6Rt1nyI7L/PvSXOGlKqtceX2032vQI03WPbUImOWvlafq0N72FVvSTraoP6v
aMemcu+m6JUh4Q28uQ1m3IoLFNARwCAq6YvmkOsfsjg09MG9uzcdUg2qfapfJiUedV11g7bBd1LI
qrmvGgCIqq+iMUYoXMGd3NVh/tLKjTW3nYlmZYce/FSeZsw9Df0IkKvayHeL/Z/dyM1JmlVp2gNd
R6jyeGr4CelGML/EjnZxLRT33krXbLTe9wAkSg2NT2tYZR6FLddU7gmtEWJqISCfJNvRe74Y6Gbu
zomBFekEn4h0S4aQIpaXTNVT/3qCdJ8m2oNkU+OOTGduwqQxpR2Cq8dt9Wx7Czjpwyt+pIk1VNtC
xe8v/p8R0hK552ZK1C2x24Ns99t6YOAKVg+Zm9cWA1IOkJuV4x2wVV/w3fvSB/f9t4GHWKSpQWcN
JstLYKpp80T7e+BlBmSx2EL4vJQOgWCt1pTOOIt2VPND8gR1G3hv2BRbj9Y51ogz1HNWVoQm7/fs
1Rhjr0EpYk92/+ZMW4RMXAtuIrWvQk1tLY2QqOS/ZE9eBCZl5lFMc/VqxF89z+bQpqA4noA8V6A9
/PaGa6+yfFR8gbYUd2Ev2KFVnFEKvqKVVUdtsXQ/Zr1mEYB9nz1clDjUDlW5L3Pq8g8TOCuIbfrN
471hI/jDZ+4UGcQr1qVM6T9Gy3J4hoENQhOtb8Ow4WldvM93UrlXRNNWnZhYGAMHKX2QJJxDCTUE
f6cWyJNt7j99qrxhY+N0Ydp2pDfM7Mws3ns19ICkS8XmGc11T7MO4DHPf4wio4lJYwKIZNrucjn2
hcaUVwA0Qitt1HZv4oo/CSvRUWw6TsY2J+LgF7FYVUwA0ntum670wxCrCU/phrT2g0RqyTbZQ3L+
WuoGUImzHnhc3nuT0vKxfamEDykIV7bS1mwwX3AjQs0fqfvfNqtOHTM4CY9TQEXS4Kd/4aqUsrZQ
6fgV9Dj+7QrzYAsDm8VT8enc2tzOVY0QPGflYmgRr2nvO1Xe/tW7bRh42ze+v1y8FSYBYhSvsJNK
IdfObW6CDae/dEhd6N8ILtfuarfGY6UNTEzOZfWkjX4km4kyTaIQDoonMp3lbRSbaBBSXn4QTOKF
sK+4v7UN7itTuWunr35gE40oDWaZvBTH5ZHvuwiFljWnRDhs4tCaauRJBEQ2xNqT4Qcl8TA+yHF4
xjTan4PgBhbfKmvYGmFPLE/UiAntIEBJ8iTYMu0VxNdspXwmzjNpQWr9+vugJYCvOeQsT9osq3LA
YRZYQKjllNhjKMMAoo24mRDCyLnrkyd0nkUbTdr1QA/femSEPPuKt5wuppfwS7d6Zt/M7HoibliX
EV2cYIRPfGXa/o4skanROL3TbKuHRA/VJzRCu7Pm/k8GXuZIejEB8dRgCXs02YXA+aNIGihNvipo
Xy+gs4tJqBVB39seU7vQ03VxbNTWO+pPPXuLz7dk2AD6QU3+F6bSfLijKtUGjo4rpPORTBteJoAF
G7hRygelKpJWBCl4pgx+2Tf+qDxaukUEL8Y8jtEN9DIf4Uks2qnD1UVU43luo84AkfjVztF2E0wa
BdM3Ohi090+go5gkwJvcpqCUPOANmOKnw4IG/tyAgpQq6gMf9ZoRJd/LYVnxBXP/1FYuwckfgSs3
uouk1Zp1/k8WM+9gnm7VBbd2yU6V49NrnB1Qn2nvNvtemjc1nFKteNF24xKTyMPAgfFsTq6hM6jJ
b6Hhxlu/bQpZrAmaPdfFsMdI8Y3UMjK7fJYsX6C6kaG1fdedr2g5GQm8DpznpuPC/coZ7r67zUTk
pwlG9ZZPPG4nW/oqXU3sCX0xx1slp2FtZj21eDGZmIHF8PBsKTMl/by6ya0JhV1rrnQEr8s/9AnC
8K2OYTVRTkK7bCoKLXOnpONvVGRWy2OLnGpYgw2KvWxL5RL7EmyBQPSjba/QcFaCggt3Sgt0NnFs
ZQe0FTTsI+PcaAjvFUO4tQj6rbbFPt62uLK5RV3eb2VtoVthblxf3VJrnKT/an2G4+cllQPKDkdG
XhhRLwh1FCCSdvcpw8FnMOHRDGnX3agAbqz8doLv4HjgP8yVvkRUH63f7m008DtxB6n27DpZWteE
q5SQSfq1+K8iUElwRI5I0E1OvLPfDpXqEJ8iTnoRNbq365esH6YgmoC7gxrIYlg30g2XFllKpVpz
9hvaeWD58e8RPgi4ssd/I1VmTIS9NsILwYT9Y9KUzS3qaQ57/AxSbKPX1ZMAAUv5zN+8RyG22vb+
OVfGOKwYQrMjOC0WVgpVHMFe3dYkqJSXAMgi8Ke8Ybtj19WFANecLOOdS1Zo+t1Rn3McL+3cBG5b
ejTircsqvjDrVg2PT5ppiMhItOHlAFs2e9LWrLb9ZM0N/jRCGxRoM6pigM+khmuU/hhqADRRHyA7
e4btQfxXoMTJmFEfGCrUiIE0KcExSO9LafOFKToiwqCD4n0VI7iiXqCl398aTqaFB20nAI4vgSEo
FClQtByLTL1+ItRk3nX93MTD7laJypy+Zyiy8LZcAlhX5SoGP8i8iymbsgA2g0QE167EtacH0vts
vN0mipBipxWAXmkT3V7d4sj5KWh1MpmoussbRYbu5aWSFovCRu25wRvwhjMcrqJy8p1Q06U5diyl
r7PRRDU5u61Dz3pUHj/sa730c2C43MzxKhnseXqpbdBG2EpgvjoV4F0lH0U5O9RDs9VV16mA4WU8
x+Z4xIUZABBxfKLYcfRcyMEmKogpLmQeBfjlnlu9ldajfL6eHlcrh4pqiOpw9MiLKhDV2+MDyueZ
28MT83IV5AY6GSE7TFODTrizfKHgW/+hbb0RSHKu4z6FDN9OBCzFhGpfFL3rs533c8lLAmtoU9Bo
r9uBeqWzY2XoI/ih+a6BX8RDbD6Fn5TGjiND5ES993bJN+h0zenfLv5krC95NM3M4d5vVSWMWpry
BJ47rhpcer2TBY/ni/l0UKwz8mDzyadarAvZGo3oi8kUl3vrVt5d8PczpMy566iFoNtLrQsLwtoL
+GLQQSLBRA0xYH2/kwt78+1i/9uE3IfM+HyYsU51mgTahYUeJKFq3neo9LEOMGWp3Fqy+EcfDdEk
AmVf9eqcqU7jNeLIpR0HWNQupvyojL2cq86b7G8jxYor/X421GN9ro5OeCLqb1bor1BN+ink7ifY
iru1xU3xcrgAZN30ua7giQPKxon2KgFJVbpTS9ms3dbOmRmq//p94/ElKxtAygWT0YXgpAhf8I1U
GOPNMm1Y9x6EpHJTk12qiraYlrmhXBgdULmGY+3Fg4HsrLBeEOJP8MLAOWNvRUbldMmtvdqIkItl
CFIzJYVojicTAqGLpmgluoLTL3+oi5UPYJQ3x8GOooDIo0OCPIxywIGji6cshkX+zAS5bZAWGQoe
K0wyeyU9Nuh/oJVU0fb1Q6K9/bd/rY+173mZnH2JeDUH+V4UoUadNbIWVv3b34009H7ULEOvGYJR
BCQ456pruTAm7DCv6NeTzc21WGtd9bHTm27FafX1fgvHyvDI6l5H8wzvP/6ZnpRlD4DvzUnf/EAu
fVzEh1UZ347k9DMEYwmIBo1OBteBTthFUHERgxgPqj301t4Wqjq4L5jyhyQ1L+7Q4lS1R/TThysX
r0ofrWvEnIlD5B2pkuQv0IML3Ltg0GvPrwf3w8eeDFfpP8RLis+mUlF1y1fR2DS/9sPb1szAOGSG
hBi6s3YPpKFGvrpFpCadOS/5Jjt+mLss4y+/3sX6Yi5HbQdHerKowXPQLuq47ijt3njVBSusM1Rk
mUrXVK3i+z8jwpqhKNSXk56lBI7WVIyAIJ3CUa3LJKGZAATCRFWtAmbULPpL3s0cMB3UizjnrnIV
S8TibVvFY4y2jKZPC3vjtnKEuGgl+8z3Ls2k3DSIkzmS6IYl+cNTJ2H8YMaE++apXjGEStStfp5P
ngC6TwhCLfS4B2me3wNOs1BaM5M+SOasSFm/CYA/S6T7xxoFQybBk2UwO6WNjQ26pUYBmSwQad7Y
l5p+NKOy42t6CNGox10pVPRSabEyiT3afMOnwBmWv2ifrKBysv2IL1EdYfatZ5fg4H7P/6ra1fRT
qIucqLMYWdq4KbNMsqUOS1VFeiljtz6Y8VhBmYdmV2ezkXvsP5/7OSE+hg8ZuPw5CrYU7uK3+94m
p5A/j/Gia+2pIge2DtmLE4Pl6ISkV3jnbxYO1o4T/7fLHcm0/bWjaFq6hTX+rAWuCvyB98fCKl7Y
pngpWxz3DcS4A5wIfX0tIksrv6OUGq3MXm9EIt/Nq6576zaJcQqZxGS3ZrBkGN3jEXipbV8fj62b
a70TMatKWHOFUEcsrxisYUDmRt6Y5nL8qnylooK1kiQ1GcioI/IkAofQV7rzGTZNMH0ri05l0Ljp
3R77TE5tAMpKzTGMXfPHzIC4wJeFW9z17N74cNrFFl82JusKj94+QgVFc3LSfjBr1a1E0X8n/wgc
3/p4rfSMEcCVM0bQypf34slW86KLFKOnJrvVos+22Hsg9v3wXGS047JxZUgm9Skg8iGp4flF8lYb
UCYmekFomwT1LRZLLSeusKtHZHDh5sni7halpO/muXNS+8ATIy7kPfu64/a5DsXhy8sWkSNTQSZZ
DoiLskAQwKCa/dy4KKo3AMWSHaty3evpnIJZ9+jAvUmuF5zIZCJV1tn2juNVfv7BYkkCfYCh9QfH
VjgDTjXqalFKUwmkR/sga6VCCEOfnmdBSypR79/bMquZhPkTaN+Vmg3e5pZDLSQPqfhSzWA+gzvv
kY/OiEqA0xdlQGW/MHjP0VqbvCtWXZFlvkEh/Rpl4CldlgOf8UDKAx3VuQhi3x/yMzZgaYlNJZwe
rAHb8sCTBInGJ5arZ5QqWOTkTRqwVHUssRikbmS735pVMFXV9ZPndNw3RRkFn5rZljzB2OuBe3Fg
6+029rUJPMbtC35P7aW9KqWxXlox+N6V4XDe8+HtW/FWsuM3oWQjw4doRzghsNOsO41qA9972TzQ
ncDf/25c0KpbGb4jac/4OKlLJpgV3hFOkSy2gug9Ai0wEPgc3HTpGrKSmhFzDpgWw6bAGSnh9H3S
3gApPe2DMoevipClFNYs5zwTIAcvGezk3+Esq4uV55SHi4dAMzCoU9hUrL8xRw/4xX/zY0QhaY+h
GLWgstnSdR6smgqUAyEA9YFqEWdrJ8oxMUKy03GdxLNO0wrzZrnk//KBFCsqJdeYtugn5xv1CkQp
Mz5JZj/evatYQJvGOxO2PxwbQ0M620l0/Ov5Yk3PV6wlO9gnLmMLEcvr21GQbSm8JZY5I/a6P++C
HBhibJ/FTA0JnhPopKdzOCGZx5TVA16nMPpmlBZ6+h+g77NYMYQFjNuK+sV4MT5Aj4juWLBoNwAV
KPC2WGPx/ripOEAzOUstKbUAxphZXDhMXtx47RBXCdYbCeJFK2n7TKB9sx8N6pAyBgXe8w7v9DQ5
spGoTFXzvaT2Zgll2VAkhHzI5nTHUYVuPcHvVQ3oMb8R2YrPC2jnprezG1vvLyMKgw7p4xJvl9dT
/3Tm53mgpNjUdh2w+xBvXFBV64+wxPc/+kKvhN59cE0S73qsa1VrCec58jQ0ZcwHXRScumh8Q+XZ
+Hd2L+xZ8q0nKZ8V449rq+Rk5y3CSkCxZinyT71je5nf6EEHaixiB49pycjFSMb/25H8i1CPmr6E
B8cpBYNwgJ6u0ez07KSuhzPcSc8qKZU/ceNyQQSurwte2UQL1Nsnmto+2IB0PtRoW8Hd364aAxbC
hFausl8FPFbZ0du7/OsUGCKfHfUryzirw+UfQeLM68oUqkXlPxDzK8kXwp4wPNklWc47XVpLU+9Q
UppSkvOeePyXCdddE53PSiVaypbZja2OHqWfjPI/ScW0PDAT/rvdgxasEcvpWafSIF0/RojRozh/
4FN499Ubz0B2t9d4D0Fl+zBaogepvf18nj2btkD7pVSRufkqGnaT1ple0Zye1ZnSw6wtXmaQpXeo
wQrLHAC8GJgb9doO22k9Ku/185jImLZRTa3jMTb/OPMU9a3z6C90iKZftzugc3hqFzyuEva8vbiY
x0Ngzq/FRe0P1pp+SMpAksvdxJSIrSB0xJXgNkm9dLJe5GaO9pte4eh539/IXubaqhPiOo9bYbzD
BPbycd87ZO0QPKlW3ioCL5la4hhAVcqUPJtCzpC6EYSQCN9wRXdGOnQMA+8UynzdeStAXiBlcZpN
m7so5K7K5saO36wluLCduf4KmFDapia63V4mVbWyBr/YmYY4qz8VnPQ9oibwb5PtZOrhdufNUhjp
/UkF9AOB6Yf4DXJtDhqgPqTJtz2ZUmzgh9zpMUVHd4KjtxGLZUFJhcd1CRvMLUXQmp6xsAmhW+gR
J9I0rsWvKqPgtA4f342T17nJzsMk5Sn45yBSjWz/qAKNbItvyVzpeQ+oV0dsjnppoxTC5R3HfLPh
iuooLEGMCA35+q5I5ur4b5V81V4vuVzBQSifleRKgMMUPpD/SgIbIdOUNGw5WusdtGFr6A8OjqTC
ZuoPJqU6Pc3ZOir/QsAn+nOnS5KAsRfYVeG1cGVbgTEwUofCnNA5EwXu1lh0WAj6eE2ccf24gts/
G+Uv2A23k6decSID/TX/QkYxAiN5EmhNVynKFJTOd7opSSYi7mGuQMPzXwosAYM042hwxL2V5Yp2
+pZbjm8fxMX2+cLxmj7Nxf5pxfK2ugNlnYeHhn0sdtnDRqrm0E8FZ1mVDgw2uZfx3dmvj5I+JuNg
bnmFJxJ48Z4/f28RToxQqLynYwxUc8mlZDkrU/hClZpoe7qV63qYfsbFZQCCay1tQYIAVmhL+/T+
KF8Z7vE/x6LkYNW+LwQJ8c+QuO9tpIDplqnOrVa3lLf38KJIBM7dOuY+F7GbynARGIiD+Mz5zlY3
V0Wb6dcbeqVZQL3e/AU4otawBqYM9Ok8EEobk9NreS1g93bxySKrZV7/FYcN0tKWmTPHNsY82ya5
HI2bQFwtrTlvSx8wXC3FDDQXPes8yWf1axgPCmUujQWMP5oSpkVlLdcPaWrSAGSXcN2Ccyv9HLg/
aMT9izFIyXIGxuUzlZQRvb5m/MUkk01Do5ZZ4zyqf3TDt1E6e4V1KZtXfYRSgYrIJhy7nQorD+sr
rdlxndc9siKS9HRmfpKdWkHfu40cSmds4bH00wGsg+o0TQhZeOcTSbO1PzHdKZpg7AvFoairoorI
ctRSucdY1dFeJ1nGswhe7fJOQz8slGMqUQIUnbQjnLJ93pJw4rfV3DX9UoSKRo/p1oYNUYxdmxm9
ds7GIfY0mI+x71Ui+MNqmCdZ1WVxuQkR+SopmZLW+X6kvZTN5JfgvoD0SgedT1L76egW0gVLujCN
lpl3zsa8pEF4rGT1aaDhM+8r4ykHOS/tta5e0RKqE6Yl90K/3eo9bCR9dBcEvRH4ClXCoazDYwoW
s4bfXplirhK9FWjVl6ycdTxbChNfeO0+zm766L9t92yICXePAISUf3TyLEmFO0VO9r148TMKziji
JvVkHrS+LKNxfpZAMKMawquObARi+KWNbC18mfdTOeEUFnkNeNoJZaFHWIyQaOxCUP+ax5u21xIJ
frgZRkYnuRE6x2Z6OYjj7k/z2xRulZOjyT2m2gijjIuQMwz2xjaw/Vsgu3hIL+LHfF8CkxKl+alv
Zy3ItPABAc3oqMS5Jx2nUlgkfbs8y0ZBU69ToEcoZ8nm219yhfPiaz1GlAbA/k99Y0REhDSCBtTI
CA2fJ5BrTc+mp+JKRV12xeTKYWEzwkVcheGprYaRHIyj1Q/PhUzFl1RDWlBO6XI8lzgUN+oqvyx6
9CJuZ5xsUOH/pwhkkEto8vrklhYdmNpjh5f2pcA/UeCokLJsHPkfQIhz9hWLnVpme8dGQCPYbAit
520yHavvP1QFN6prdoMVDLxBC178sCFOmMilPxrTJQ2wpJJ3KWzhRRpl0UvHbmb2l17C2y3n27jU
IUwg2tkCCReE9ux09Aoc1Je1Vz9US6sfjsgnud8qzcooKqZmymn0PcvdWjFPv2kGElays5TgxIlr
ua9/cjR/dRs8KsuITUWPSVQ89drOz72YkzX5mQRHDM7gyigk9qcEtzcRMV6cn+UNnAu7a73A+KtO
oeQFuXQ1qL/IufApBtoXqooYqia5n79foKodJCHo8nAlQ/p7MGRRPaZ+gKFwl2IrEeqx0QsVuGjy
u4IOftirNYke1ias/Fx98tpxoTs7u9w3ghULrQWMn34lSpMGQkEdm5UOG67PB2k2XaBzfHCJyLwp
8KsPvCcMCn4HzCEtkBPuErW+GBiBT9VC0zk1YXmgxd9Oa86rpqsMQ3XRAT8CnTd7FhLCoXlxv+jo
T92xkDGHrV9kHXurEweM1SaJvEqWn4ISWJ7bg82y46MS77Xtl0f83MqMucw3EQd3mtXD0BduFfNB
EEjho0t4ATyRLSltM7Eo3SyVJAYRtW+aJq6BIym9u/cn7p/PkTjDXGbWjoftFryjJG8WZaECaglG
jU7pPjXliYBRVW7+Dgj4y+/Dzz2flyYMJ6HvzF7QRMZBLRxMbznFMiLZB5rJGRErgGuDxE0vdxNk
U9V/NoPrF8v+YaodFGB6vFextX6GtrnQPOY/LFW9EvIOovwOfSqZJ2tVReXoGMTaiwAL0b+Fcf1e
kels0oAeGA6P3La29rOpV5eIaIpOCfNi3O5E7lNGQtyfrlcfGpLd+C9rrP+Awrl36DahQvaf6tHH
pJSnNWWG26VEbQUkOIUo0d2cle0lKLF5puSDgfOnECwRiXHG96kMPW30RxWWNMfCU+A+FwwLyDLZ
R9IMVzPD5hy0gjoj37O+znQzMPgFfO54NH1EPXKmIugBR7FRvAV4D6QuQn0NUjaBPZnmYkGDAVL1
07NZ995Zr03juqdD81zXD6Litrou9IwAoAE67ebq54NVvQESUQC5kecU/eTWNfhrbVbqtZhiMMub
hwp8+xZlACZyPw3hTwAFa1NIXrNUuVxJTzOVpQiGsxTvl9/8kcwqxplgUCReB0FWIxrXox7M3KtF
ZolccLjH71vXHqMN+cNXxl6FjTsrP6+079zoa9lfLXHD2hPa7WkpIYsRyYHdIbBrZ801wtBGLHty
jSH66FMEdM846rR0R5ODr7rcbZPTx/tv+pjHJG4WVqwEbIhMw7mrmkoVbyF5WZGO0ztkFqTsiwx7
Hll75D5rEJRr0pM/niVZFVzlI2WMFs9eE/VsR7q95DzxUAkvVHotWZhtMeNrL0ZDI5cUXbEN+dyV
NjsLzwT0zp3b4UUu3CkVOGukjp4TDDe73VtU56PZ9lcTeIm+nhKw0yb4BvF1t1WstEG45dIqh/BV
jKLQqr82oOXBYPxkYC70woSkLvo7efVdNgluK9ctClEez6bnffVx7Xq3FigiklwGszQhda1HDHZG
/IP5ovaqaDpN+g78aoBPymG5v6iGXNZLbXT7/Wg549OvD0u7Njz/3r/1OBULvRk6G5IMM3Dzdogr
oD7xWlgzATYCPUlHUpMob40eH+L2sxcnoB70sbkZc8hQLsEesBIdVkASl+ctguxVTo/eADGPxlhL
d/WMOxhulI0oz52kqCp8rpqlf3NQc5Ntv1aD+p3FgSbjgXg44VJtesJi2XntW/0NAvtTz0UBrx+c
SdngG6TBArsZIByE9f/NW3B8qz7f3CFpmIWsNz/SOff5VKHZqAfCjH9CRsexxugunAcVvlTqp55C
PNKnkZGQDyNs9zuSvN0zSir62bbmJ5uFjtzoJw7XIlFhvsVvVeelIHg0+OWCwfiCzliymxKeiFy3
/K61nqBi1qtf+bgPs+/PCW6oiVM0EdPzTGqVqKr1+sIbtwCJr0JMIGCEppgqkIJuxkshK/8Rjvyr
mDtpkJggrHwA3hW58mPx1B4kTFwPAKpqPyN1A7Ewk8hqWe8sWSTgTUwv0WxnPlawND6ylFiGWCY4
kI7MnQvXUrkfoADNtiNkOoVpOY+bdTTzMaZUCfZUD5VAAWacdRGKjl3j7cpQfUGgcsDWCsj+RkCn
S8QGby7ATrDI40afr2e/fUNHKGestslmU4hx3hisZcjKmvv35iBKgLxyHssnbBatdO8JgbbuseaA
1cKAhxiYJl1IJ6FbpPXGwfcl09CWUziRTUj1b/vZU0CJ0YD7Gumb7pOicG5PYXonY1oC6G115WRq
ZUFDOqgIWkRkLsG1iqIxcQWqmOcL4w72PnSGm1tZprx+j/qmIx575ef2h2qkJYWT9eyd60uySFlh
0PoH1pnDQu4LMgKYlg4/Vm2c4RXCs+zLcHce3W7Ew2/0SRuZFoZvBw9IxYeC/ZY6WXFa4cpcDxZO
s3bY1BPfK3g0kpGNaOgHZqLOlq2UMjShVDYtYJRp7CNS7Ua+yNQdeALQFl6b6N604QFyoZzOkmlU
fXGDgp8dmZ+5aVC7C7ElEfWCF1frCrjgLSTb/+GKlO9oSK8SWmxZLOj3R7aHKZCsQRcIU8KE3UXx
CrjEYvA+bk7EdGXSSX01oyn8EY0YRUEbiyRGW0N0bJpoUDAVsOriRv+uV5Qc8lu010dB1T12Phcd
nm/Hz5H0/LrlgJDru6gH62Rk9JriERbimZSkU56kMavh+gV38Nxx1NF3hHaJV6L3hgnnTKK03ADn
J75reU5QNwgbnxMaxw3zkjhkRNB5zki7K1F/+b+aUyk0L0ctRdTe83O2INWMnaS/yjTiPDOQCuEX
39TjV3IpzqlPdiC0/z1V6zbBKKnFgX4kD10Efkdx7bvw1zHdkp6a7y5zJ6024JhcxUal5z9NjIDm
FucSHwRARmt0aXbKpdJ8RMo/OBC/iTnmq0PCn+eV+xVQesmytgUNwPw+sehNU7KXNyQ0xR32dZia
pGz9OT1Rr5ierkj/MU4vK+fmEs8WSY+z0aMErERVZ3czjZw9bVFtdOrOzk2jeWlDhReJ/nCkAXia
G2Oi90lPpP9Z/F4RF6YXlHORFk91nOpPvNAtuYtRuaLmAg8NXEijfpShghxafh+F62wEV6XtDC9c
vdILQ5ZTAMdv6rQFkQK1Dp2JOTxk9J8aY+T3sDOuol7iWsjxt6xcLANkUq0GlomnaJVQ55MsHFBj
hprTZGhcoChXpcmiJIwjPXp15eGe2EvUKR5zm7fwEjQyVm9ZceIAop3NVDgYWze9m3rxQMvVaKXO
ApLYVz6tiTs39pnfYSwCBuIg2AqrkB9BSCuoh59Wmho2XgXiH8t8sNP4yhUG64b20hCEt86RIb7J
rz8xI4/Vpour+yQejHne4scbkHXkdA6di5cCyGW6H+40phGjAcTA0hqZfd1aA+i18CmQfNu4MDdy
WjM7gwl7oriiFRH6Z8Ck8gMjwag+jG0DHkkTxDzUFxqnp8IOYsFrMS1Ppuh1D9GmKc7GR2/PjWRx
syXzDmdfmTp1kDbEfudb5ti8/KAokLMkivstdZptNqSDqedIDp76y5OQiHJmHbSjijyI+yEU2Ui+
5m8GyaBkUWve6QhHeEV76lIheO00mzYIXMa+dhkUcgjtcWvFGbExN49O8iIz85t3a9Q3/Yh3z7Wf
MW/z1jFscNo1nEtvbK2YZeXqsLKhQiufCdeueA5DvXi+knOtNksZ28cpJsV9+XLTGzSK37WDCUfq
18Yl9GcdYvKaHF9RrPPIkMxSqCQGvnufP1WX5nvEzczX4AyIMnaHTxHbw/FuQrvcbAXYMb4ZvH0L
LK+aNRqDQZ/HDmNgf96alNv0TWWqTnm4IQ0+ieFtBYQDyj+1JKOXxF3RfAG4ICI3goA7ltT6yoFQ
pClc2G+6WttTQ+yHNOAL5z7bUzaSK1H4WjUvUe1hL457X5cw5mtAJKUOhpmzWQcND71Qji5FUrHH
ZNZSsHVcZUa6FW3RYa6WQGYpRzug8QdBXh3Arbz1OTyav7Wrt6f4A9vYXD69PeKy+sJCvdInO0Ug
uZ6g+obxlsuTVKwpHUibloyJJlfJ//xq6+UMhbKeUQSEtGYBzTTlFFWTuIZ3lojzkExzDy0xTU4/
4jhixx0CbemHAPEHfeNh0lnj5SXkb1/q5HDR3oFmqp1m7h+eH2GIBxMM1s/inBvsqRiEUUC0c2Dn
D/eLSb69Yo73bpUTe5bTQU9mio8Tysqu5A3KjpRrbpm+YNireFKPZ0w8ty8IDdwK5kW8rzwOB5RK
mdreb9ll876w3k7QXxhlMcEasBohhqfd7FKzgDtupmD6LeaYCH97mbiBQlUYDkC5yGpBKsCZk3B3
7Oj29x3NykflhmDjKA1cUeKKWIXZhEk83thMs2qRI2aNC496oIQxkwBN8DukgfHVUmbOhrwLcbLz
1opOSBccD9i6pZHwroIWGAZihwKelQmYs3OmhL6cyd1l2ctCbmWuwR2bGxwSu8Np6kp20vRitASu
WgnUiOzJzRMFZE+s4Zq49tl2wjD2HNuidloLSu9KotEbz3fib+bcpXMpvO7WMWZj5+8xEidNEVst
tkm+xlP6LYvFbD+1ic/Xa/wztVRfmA235Mv3A0A9TI2NUglfZ28RYDeQYNs7HPy0RE+BVfpwPkYb
/0PUGTADEVDhwwn4xozuYed5XKg1L76i8NyzDNl7kLdQoORw5VbMUS2Eelb7rZNlXyI9zp5AiE8p
DFpOLIfrUS954+CYucqFU5boHwssv0CPYqZbitne0NCqhH1BGsY6+WauVb9DplvoIAJroQyf8eD7
pY9TjrBp+hGCR/VLBeBlF77bEjnc9P0QCArSNHT19t/0LfaJ3abFZDaRibjRCIb4jCezntqskQS+
Qv7KezrQs86j8xXZAF4iMYCPmR1p/wiHPIRy6C4kENpuFtqausYAdae9e60M6e/vdeaX4EPIX65R
kha73r8q3dNQhm9kYwnMQK6DrE+y/YxO0ceqep35d8R2i1txMeEaD3VUXDl3bwXg0OftHxieKLpS
pJL8WiVhzom4NHub0LVQdU7bZRwJNFRJMkEGFnBuQ20ohvqDAFNG0HCZn4N4popON2jS4hw1yz23
gHHNgA9Iveb9RbWjfxlyckJO58XdatMmLj5Re1VYE2bpfMT/fF+7BBT3M3cuv2E5NQKl5//IafSZ
hk+PXcNjgengWMV1MB0IjfhIthAjl7FoGHR7WaVA7K4hs5Ag6UoqeVNJmlT2/ICrYcFFyLeJeckv
gd79aiJK3uBHA2yJ82opuYaIRxDVC6woOouUrAXMnaL3aci1ve+haRaj6fPKuqe6AjefdUKzG3vj
jV8aLWx7uwbBhPbbaGoCr6ChYHbH6BFordQpCcteNqLOPBlXs/QK0Yc2iCiP3J7bjMxnL1xFik50
maQAFC9rd1veU0ypVfZs4aQzpOj3UDSRxCnz6GhJG6zGshiLQamu+o0tNZwmm49X07yTB+vnltGm
J/At3nJBqPHoCJL/h28Lsl6lb4AnmBrNeuK6053b+TPgP76gCT9P1HKWURezFUzeXAaI06Id66MV
2R/fwIUehibanVh3oitDGxtip2UaG0qNCjSddKsaCKO76Q3A+0y2g3a08U9FnsPMma8hi9DRQNjs
fmuqHb6Qor1el84z1/r7SstloU/QLFCFSD6FmlII+ZtGEFHcywQVv/fsP8DQ0FkvCX2Zwe5wcbvK
yjWW4QhaF5lAQk8inTuT4FCg2SZGKgmYMuaMR9w7se3ex2RVUYjrjMKgFKWuECzJu1kyPSsj9iXw
WILXQG+YiY2leGUZs/1YKwLdLGizcuAP47MjdOsEvbE0E0qPbODdwK2bftUSl/v2NxIZeIusOS9D
66C8JSz7Ef6C/bBxh7OAR2bFVqvylNzv1QzmUECK/IsLSB7QxU8a5P3uXvqGIEfUJdt7aIQ8+x83
LgXt67GxIdf6HDtIPI5Jfkh/FBLkvxkTzvhTbTM8gkiaVBjmX/EHiuo+lbyxpgynULj/thz3T3BP
HbTx3N7z6BtCWSTe/Xkrg429Vmm/5TJX5WCcaUumnv+D9ukplX7VV/bvCs66aqCIkKMvkK56NLcN
EZ6LZs9SV52WcQWooAuVdaSe1fdHolyRBhXGKre34SgVE6zkHTlxcK3sXI2FVQ5MHLnPw3GNZnRa
1Cv0lGLeIZKck/LoxcbqPiCnyoUVrXZINM6fJhoxn0/GCMDPOUw5JKpmNsbosi84rEyolq2xL2/l
Gny8Yl1Rd+nKhFC4o0YQmXXH93rVV4FCjWeYMVfs8frlSioy+x2J4nHmwEP+sWStY+lRHZy6MNYD
fprVpNCcx9DFa4FNc1cAoaSGH/1hhhhrPzwLxdyzjb46CZTjcrmub2+6FP95bwbcFhqTEPFoV+GX
zn3KEj0GEw7ryOJOvpc6tBncvCfJ15qLwcjRTHNQs1nH2zLSTzE/vXA3b9ApJ8YDk272NKa4/7CI
X7MliRxMEFTk4JZo9KR8VbylTedGpvpbQ9t2jo22gFPb4+0897jtzFj7NEjxR58n/8I9WXLTuquC
I5kKz4R8/lVhxX1KByJ87aoT+tuTRXXW3oDJBCx5sF58Ssux7RMF8bZ60r9gxjVJ6xSclnqRUmVW
rgbIlRkalT3YH4foDd8Ho9SIMXv0fWuacfHaUSY90m8n9POjz+E88+N9hp9AnAidni6W8agFXCdb
MsH1u4ixY0tU5izuvAvWycbsxbZcq3y5vBMiyPzrn9PlwEqs1puPyUPadA9qS/INxqL/5dkKGFur
DbBqvu6JcMh41F32osglFmW7L8YI4sHRWvRl4sTyYi95qMPEZ5d1MSQfm/V2b1R9hzKwq2WNobNM
zABF+TnlS9Bt+6UMXsY0dd2Op/JSSvuTQVTdOzfwTX1KcFcdDX+fFbWh0vW7LHygFRUATvrLPyne
DJ5okj74BAAslut80ayhj81MWlEJ+i2ajSfVb+thwJvt/A6bxVnRJ7Y5VcTZz5kKnEaUXbcntRvm
FLzSsL0sbACbm+UcsNBT6VwrzkclVjHLjfla9l5nTwDEcHSkM5DQkUFfxhXzkvHQ+wQ0J2L8W222
cqWjFqaS+Xqn7PPc3/n+4N4TKb+148oO/mIZy+NM9A6jFqQDvP5NfQortUU2Wv/AanyJ8nn/RMND
7G3VINgbVsYQL3PEGBtNNnkg2ikhopv8hPI2XAvdHR1iLP6yZch+rtaJrfNCPHUk/MJ/ua5mg0Ap
iB1C5Il9R7s0UEup/FjKLBI4j0f8eme2KbvGPCL3C5wyjBavd8B+y77VSOYo4bOX2btLkvFw75rJ
dnTg79CAGlIwNmDNiL2YdwkxR5JI5GReGCtHYmlpzXZcUaNjVMF07uecvLo0LyBqb3SmP4ewHs76
ZXAeVDZJQrvLl5f7LJDF7poe1k8MAhyLRFkU2vu9zFYvuPrxR+nOoiFLojCxkoqSK+KUkX0FcNpQ
KC8qB3gzW8oAxP7qWN5dhOU/5O9/ndA61dSD0l0m843I5hOma0CNTT+DnM0eLkFBC4dUaUJqQZAl
+rKW012eczQJRyiXXxxHFGIKWXoqq65Iyb6yzjwNSJRqL9N7bxJ+jxvgJgX9Xba8px18sFOfruSb
e+XAtW1Gd8l+keKIM9A1Tzz/x1+nJs0t/gjoJhYbDnIRjixmyggZkhqyOlm/isTFWxA3br9ScCoQ
qgI4jy5hVlEeeUEBTYY/1sqZ6TwQjC76LkJz5rccCzz6h8u3ZLaUHs9zb23VTXw97yo2P5tYl4Au
nLAJGiuZwSHkYsJBP/1WvrpP/bU/JsKer9KTGrOEtlnxy1ynq9K2vcD6C5gr23dAffKNrJNMYisd
qyApf8JMSua5T5fwL4smqBMzCH1aIy6Vx6GhLOwO3WeEsKsnPouTJKWM04FYlJCoBqvhH3mKVgPQ
7sOKjuvJCL6xQqK3blINI1d4ciEJYLuVk4DLYQgFU5JE5yXEBocHjAlsABynF38/Mg22GMmHJg4K
cCJ3doCSroQ4hf9A8rYP13eLyzrJZZlHyCyhlTyAsvgF13TUyWgMjYaMg6VbpcC5CQ+fs5Kv0hsh
pOzrsvd1c2d0C16z4e0hHlGRVh9C/Y9/zYtg7YbCk+d+vo/U1ZdsxRnoJtyVEl0x4u48P4cWMhD7
XQKoWWWSZT3BUI/C7rmoHckf3fZbo+5ZiIzOeLHYgblMyIj/u/8nmU/nV7hoy9W3yKnfuz7ttEgg
oKceogE/Ng888mCbgLM325MXKyabY0exAvMBWfq4Hq21hY3ThVcJEzjhq1L/XCTplk8aaFKVU/uB
UbNMeFs242eX9QPT5ikmzmKxaEeVBG0TMBLWn36w4255uTJqwBCAFAD4RCqDVx24YHjJfKlsF2cP
zUYb0wpMZkk6mjyOVWAgqxF81V1VVRqxLjgw1qdVCR0QNrGjUxQzRAsXamwAHeCUVCMzEMmZzSb4
wG8ZtMXUrxcgWvVLo5bKIg0FPJYVOVcJG6fgTZgq7NY0t1BJOAxTjhaUYRnBH8uGowPxy36XS0V5
XRWwkx1wKJZ9tvAqPK1DFV3TIzz4DZSjzAvTdl3tiH9iMaSEg/7T6RuJhzXaiXsW/t/eLV8IRGQK
nHwWjKfJkT/y8YHBbOSsiQvLc+6G8vdba5TkRGpHZ7otDNAZmkTh54NkdV3GlLZnzFarD9957nzA
Gix5IaB+gFaQGoTrCTNbQsKdeYs5UmsmtYSotBN7YchqZiRPMCu7EObEv5Ox4o+Hae382JIzcHNA
IbkUK0U89qhzKubFUm3rtXumeBi07F2YBav5yMcFUdYxuLhJoWvCEHMRC2Oh6pkVB5sDOvu05RmI
Ktl+HUqpr6zmPiHkWPNnji1+ct+vYLfykQNyhxNYliQML8wGGvrihm4/LnRX3hrgjpUNClVXqqRs
9ntvIJpuCi2nJAh2LQ+2WmEEnAyzHi0uAqwIxNMRH8zMU2qXU7b9FmV9MSq55rOx7NV4v6dmimQB
nrbCjvTOvUw0pbq3VCjgOM166zWBKV3uExbUJMXObpuCzdJdmaC7hkBzK15yEm1oSgXqERd59oqr
LXNRKWPRdbnR3z/ZmGTgsnY/pn1sI9onN2O7auRflSdqIuNwuxBNycd0HSCxHUE2DpSzIklYOp5v
VYudjMMedkSZjpocKBYbvq8s9baOdNt3LgA9eDKZDuy1gs/Tz9nWIqjuWGT6YrU7CMZTU+dZT4Kr
v2cg0fzUchuhZEqMvbuDR1p4BTocU69DjIvDtzuUR2/0qL8HcUOk9n6EAJ6otddHITi1/6jeF+Xi
m+ZiVAfP6vUAi3WgS5MAJW2mOuGAiqUihyoTsEq89QyPt3oeZkC3Cu/T9w4l/LLD3y1J2exuNbs7
1fRQK+7xZx18bkulzrcl3wQkH1f9xoDXI/V9cIL2ium/Z348YuGhgDlUaTZAu+aunsYilQJ6tZ9X
nfdN0CFizkc6IngF2znVNCwEj1PJNyWgROpZoRw0HVuS/ry+8cIeWz9LECXSCuLz5KDX+gnIQ9Vm
AQC1ol346k0AvEbkhIAx+EGA03A38DTHEb/fvwRJJaKamcgtGgEG9ecGRgtw/JiaxeQceSHfP+y+
SJBQIRUSdN7VGFICJtil0vvGDONNq1Svt57OXqFQVpQGL9Q2Muprk3C/XYTvtPzs6OjweAefNVIf
hoQ91xcEgtivehOfRjk1SA4MtUWqtczo5H4TK2wVT5NRk9Hz9XsJn6Ms8hR54wVP56NEsLyYTaP+
M1j7vLbFR24kEUFe8CjGPd92ppfeQOsmdY7IUTVsFnW61uJFVhzVWpHsZhxJ3U4vJVIemJNdZ6av
cwq2XIo8dAqTEcpCp6MrVxOMcLXzMQDUYBBmVqJSuljejd2XsIKW6twzj45y0iHRG+28HV00P74b
vqxj2DVVVLPKBWVKoo1/xOq14PAqZ+l6yCCbLGtXmX7cCzPLtfsQxrVxWdl4qbyZsIp/R1g408Oo
9hst0BZasFrNHiqfQsMpkvMKDgT8yaf7/Wub72vqeFM076onSQPMIZyxc1bajtMTn2a90rsURNoJ
bHqLE8/IapTM2SxlG8HiMRmkiA+hn/SqLyi2enBz4ssEIv8g/GSHMDtBnW+ljTFmJA96jpTqfTWT
x4CbWFemhEg1Pr8YYMlug2i5zMDAhPx45F2ARNg+Ec8qKxcMoCNX5gOIckPm6G1OXtLFCHsv21J7
HqIRQvTEc4f5AZxeyyTRmkmXRECYv8StoLP8R66P+rZhO/z9ViY15TfGPBaOlUDyD3c5vRhxxrcl
OkloO2chTafjZN7ait574qKAszsm5xGTGQ/cSCaGJeFgvEVhtCzIUW8GMzGPoQ7/zQFcgfK0I8lo
kkYpgaizcVK9C4HuT6KwF7R4aH0NRq8iR7dgO6mDClUMBNPFNy6xXpKHSj+fFn3Q5AWIS8rbbJAd
exagtRWIbQD+uzx8640By0GyWJ7tJD+YHLLx4Zaoa8q3M7/wKAVl1Lym4CCJCMVSncghGZc87OSF
1dysbIS4H0BoGGmFbVQH+29e91tFdmCxiND74TDHiy31AkuD6iYViuHrUvJ7hEcZ7o8K5RhzLGBL
st3w/B8bVvcAlnWmK60WeWgM9pY0dGXRNFDvzzlkqlXGCQ/WYA7bE0dp9pbGXgBQ1liJrQi+D58z
IMZbVQRaBt8dupjTphyfDgU6HfvWkroebcpNlk608sJBQPGedcqKISOMSKCoozVEbAIvU+OYENXv
4Uv2dz34n+Qz/jRI0a2517AtOZ1LRW25DB2jS91kIlHgkIRYVc7I3yvOc8NEwUYQI3u70L7Qi216
4xN7wt3mXbrCzecG/+JLNZUn9+Tb9kprSrLR+mwWLQZvEy10aHGX3bOxFCimAmUoMqTY56kaC08C
qmXYkZLC+u93x5QJY4aGIaSM4D77eqhxksSQ7T2UubE4ut1DfsG1s+yK1/DinS0PHpgraol+kJ+u
6cf9MnDQUqQIPHn8IkZqm8WaOEKr7Dpkbr4tu689aNk9EhHD3NqR8k0jHV9ng1gbhwC1yh+RYX2t
/slS3bADM0vQ2G95bOvb8gxdIsrhfxIJSuM7BDKO1Ke/s0rTpjNSyizW05iYOZRgV+KwDe7pb+95
yf64S3m9ntAUE7B7uL0MY7nNnh6zx3+f4SH46bpD7qUi8bB+SSHvmYQUP0M0mypcL1b1kcrtJ1aA
OZLxoTR0DMVXZMLoWLwUdn+EdhLxb3g/RabdNVvGsOo0VUstqdO071DQ0E3ACQ6CDQeeYzF6XYIr
MT7d+4b+xYTNtbusbTNXN3Cqfj8spHWTUQIxpw1mvupvS2yrQL5sSLAmUV46rsiSPa+lFaVL3SMP
lTr7H9xo4aOWtbV4pJPRaAYPFxzb4gQVY9OMH61kYBAKIvpfB0Be6Q5aQt49IEN5StZXt90uJmyO
+8lzhPY/dc3k54MKZUVG5a3i1LpdbkDyRk5SRuN/s6OCWRPTVZFmday5pzXHFD6UfWLwslV/Qxhz
hzB+AK8/OoaIua1mpeMRryeVlbcazuk6ip02/1a0OyHhE1zkiPsl7pg2iSn0ZaE5eYO/7z8zQmUU
DDiVVG/otXed1VnZ/l6e35jCAkcguARQJUnUKXJOknTSHkcaSodTGILEbvZP8xtK5KxeDtwaLYPS
c2Bnkr5pq68+33yolR4jdTKQcfy+/YNrFD4pIYb9Bbeal2Ryr2/a/0w+/2jPZwgiqHoyZEll1zZU
we1HmXqM2+O/2zMB+kSSTEd2ZH0Vp9jmHYlke3vvsFSUMZSPKKPYXCHZ55h4jP8x8UWudK3isVQA
M3DLn08kJEdgMecHx3w+Gw/Z3UBhwSNSa+OYk5oBAWYJV9gshqf6roSzX7430aNQTrxYUtEpc5/B
aggj6UrcqUY7piz3gcMsZOaHUIwDT71M4u0H2c6PuczQzWGechatIR3JaMI2+Sg5dwmO+VNYbdjI
khfyHJ+Je3Ibtv2Y2M/HT2m6yPIIprr8QDqe70eMs2zxyIm8gdLX6TZ8GY53aYsY5b8j69FkCaD5
9Qf0bzPm5/VH4O8ECZQ2jS+g3tToWIH+PcuOdQa7IBfASuQXZ/zry7MrqWKsAq199igxA3WT23di
uAkyjDuIfwwnc9oGVdPH0NCR1aITA92rqs57mStE7PRw2+UONH95VFE/VkHz/6BJuB1X5zYzk8xY
M0Q3/xa0N4kQ1f1Wtntn81CmcR7WbixNZOInQOTwPXKlu0zpOljwOZy0WehhgfACBdJke0sLvl8n
03LhQkcCnvWOM7szLQKDs6nrxEC7h/juW7zVEIG6593V0g6BjDAnGpvDnhs0b9eu2nu8QIN0ESBM
e60bvBUif1M/TyARKdkXsMAtvW9M87Pt3hezlLfBJTo6TNwdmLHLkv6DB2zeqh9tLdVm3N5mpzVU
dB7rj93EJzhX9OkT/ctFdiRMNjpC1fZWk+W/ZsjW/R4ye+g0TBY81rfCzekldGalVQ48Idhvhp3d
l4Ua/ijXfUFzBTTHzLDXdPrLSwKCVbcNLkNIiF0h1VK3hpXxpN71M+GHHR96cLxY3nPPhNfeVc3U
AwyqxkKWGRoUfbNjDMUQaoRh7ENcyl5Z0PAb0eS8qz1OalCPovLj0qQ8IMBr0G4n9lO9fMrNQ7a2
Sa8VrOK4qDdb0sXR0iT0VA/X/gnODZUrcKjocAMXJ56rHm4mfqLHyUxvob3IQKfQjldliFjFxcNr
B1YqIsGl930hu4gUKDocVb9RNUCmLIPmI6bCHL2WjDsHO54Bv479bUC/bk5uXfgz7/EaO7ftKR7T
m2Wq5c4wGxJkbsS/UG1zp8EDarrV3LxLLdGFNcVawHoS88dLU/ovsVLbuIi/aZ4j2i/uMBeSkppX
a86RorQbxeL1ITKiCGCunUaBlRfFWTh1/oPDbTIbllWud5LcpghXpYWtFmBu8UAoDoDVslG3PMel
q92KNrJjUBY1FYO1QLPb+Q4FXs3W00nb/C16OmihrhbKz/t3rgjtbeit7hSTNH4Xh9gD7fF0Nqh0
ee2IxJAQghyZXWewqqjb9b6pMNXtvYxYtrRXO/FqV6dkKBe2GGUf3vfZiicC/lIyPnpDDsR38pdP
iaJ6is6c1E/4gcLm0VDBXqFNQ2ywZbfa3G5xDxw+QrvRub8J2qsENHZnKX/siFhDNCBKjmiBBTZM
nlnbV6b11t69UaDeAhsXUWVTSSDQxaPISO4FsLgXDIe7JpirknIJ6LZi8v3vg3tg5eDGzIdLiIxZ
u2TJjayd6r0QdKRvDEnJHMrtEvkFb47YhrPEn/phh6XECxLF2FopHV2yzXqMOzGFanc/Ecue4RfW
SJ7YDMKvsIeDuzr6ebP04PYM+gKQbYTgIRZZBWqufK+ZeiXeBJLRUyfmvySNQtrs2CpaCjJq5hzF
8cl+Es7QBbWUxvB3wgKROlSKrOpATNTZyaFrS7XSpfL24RpN8hIP2C+/bwrXzcVVMu6oQ1UlLr4E
hAnAEb65jQPmcxesIsu/0RiyL+gh4EWCLkQPQXXse3rKXl2GVww5dUyyR9lKcGbPOf6+lC+ihn1J
eCEzo3W7Xqzk7sFp1B2P8wCi9TXjxJYR3UlFeLrcAEVpvKkj0EjB0r7J6XGiEjPuHnZxWgzWFYxC
KwmZYcji1aWeGN7NdfO5bKG9M5ixo+8jGOe2slrdeJQV+RSBzXVzd9cwwRJOKptIAAFAeChK4XbP
WSIDBLiINn5WSCT6M1XJuSmSkU/SIqW9KeBPmm/0oTelMCKXAXDpqoVFd8zPdUKPwhRp43OoQtZr
U4oxpgSb0S8zH42TVSkmPBK8uZkPAMiO8ly3hCPxo2oK6xMT2qi7dodiDKfY1h5i4Ri5QMxnyo1A
zeZLUDkZXlUXNc9lECfme7nK9b5wdp5Kv/QOT3056hlK7PuMhxetWmi5wT9gnLbm31gQ3wYwTupW
mq3PH16q2b3jkSQPJ8AtjIjexaDmi19Oh44l0TFz+GTCO2eP7IR9m0mLTPbeAQYGGeIIx/w/mR49
ZKwcippowZu38u+kpzRZx4iDL8noZjkaLS0kWsVAvIyib9mDEGOWKGC9PMtWEh1YltM2pyCy/3Oo
x/blPJTaEc4hsi5IEICOr26Nvaad/hyHLYrIs1H7KNog/JiZMBmAqq8OIqsYmlQTZFnaN1ws8beP
DkGGiL4Dg0qvHxivyr5utF7wgH754itG8G06dLnpGIYEWcMNTrViWa94LX1gsSwzcvj2sbVcOZ1y
58D8cDNxLZHVUIYaieRW2r2MuL3Nvml8zAXfN+mBBVaA2qOTGjJoWNITv1ad23y7u4gBztXxB1CN
HYWC5ZlVaJTLuHlvYNpIzJuv0vUmd6LMyjP9bVbQBf5wTRJl1PSXtuOf6WYrAfmBSKbXUVnm+ikX
1iui+lrSKLxpNrgSD1/+yXwN1oTJu8/PgA0TJujmebCBhLO7iBY1bepuqGyYtIMxjJkurib2Zez+
UVthF4DN6EXklyVkx12G6xOSOjOHC8tP9zJzewnzjcSiDuE7MmB4u4y5QogHJjo6AD1YYzooPRQe
rqwTvjfrHXd3B9bv5TIkri9cCNYwr2jTcY4V298dHbejAxTNZgg0qKqxpbFWf9HOt4O+hbydnyKA
/z+wy8TGgz7UOF0eYF9e/WE9F3QwnOwwJZQvwEUNwJV1j72S+vBA6ZXEz15m/LEHj/n+UTByk1Vv
RCpFfE1R/VyfpNsbWcErKCqxAip6W0p1cuzO+j8kC8Pk7Q3to/HbhQkeQPBvzIFJW1OZdQJfwCBD
y4+9Bck5gpNsQY3xhmlZ8e8RQmoK7EhzXnNC0wUdWA9MaCWD2WApXpRKROGmt8PzIosJh6W/+cOu
knLqAQchz5svu6b0GHJFiEmtjAcyWfpdjWDPiJvAZUJ2FMwtepS48tU+g4Vi5BQ+Q8s6gklfROQ3
X3WtddUaczsy9RGw7RjFlZWMgIK7WFHyQ127fCOyzf+ezgbwXvVUN1DL2eEu4PVcDN3L/OzZK93M
8vWp7tC43Zz9q4bu/onA5/qncpUow4hpLgKtOLeY/dN85yS3iH7xWq370DYu2yfoGPJ97piep7cI
SRav1swEIqUuRDr3FWjsFUuT4BNZL0m2ryCb+hOkXCFmwveDQskGCFLiIB3gmDTFm/WViVTUj954
MRFsFmbYo5sTypYmPkThTcrgW8tqE5b0DzXJru/DCqYEqygb/v6gQxHm57Wt3nA6Yp7oX2YygTqD
x6Gko0XvaiyUiYxRMd8h9K3eDJaAN+2r+ALRbrC06LP1dQMTwmXJsRiyAbu+g7OFZzca+T2Q5q/Q
59OKUdUQLrjcQP70zDadm9Mfc6FnOTq8rTa8F87FBDwGVWj1Mj6yG0HHgS1mspzmS4ylC7qwIB+K
ZXRiv/a0WIXZNkoxbCjDjy7egsQAXFicoCPMT+urYYmyB6iJcXujhHa8QEnINLwZstPH4qsV9PAP
RaJvsSKmVOsGoeEM+yrJ1wPYr5ZI/9IT7c/egBXQ6enDKYX4BMyb/n6c+xUExEz78N5ToE5zLbnM
a8H6/9orNrdmVq4kWlGNI+Ha63fI8XWLN44T88Z9YI4/0ydKD17x2Oi5I7VuDI8NJzaXfPnl5Qmv
UDjT4CxglJCMeM0cRHDU0/xjRehV6tsdgLAJPWtAAt7iQ1TfZrDHUIWdII3aFmcOL+mszfvaaf6T
n/35m85rzqo+nfX/UyMfwM/G3yDZjZcXpAmrAXYMZl/eRdhJvxC6ZnXPJkf2xio167+LLY8jw0rS
IZhM330zlIhkggYyFHs7POgnmaqvlDQwEiDEUmOp1+EJeolb690EJB03yY48O/0D86uqzneL7z/D
etGjl2l2Z7ez40s8GqcfuTKPNjWi1dTOOkwa903vUrxxAxBwq3Zy6WUwozNlNUxHUuN4REmD/ZZT
q3EasxjZqB7MOYXBWaT0kUUZKn8My+hSx2UUJw4+3MulD9uRf9Kxv1Y4Pb+dFuxcfTHsgQ92cgJW
tNQjP2UsDorW9nv1S1QIrYNod20MtPYPidnQ2X7cZuyljvae9znNn0GYsY3v+LgCsqAy21WpW1kT
SuprMqlR5vhMXMT/3L9q32+98bLwpI4/xDdFsMh6goF8LKctNvGLG7O7+7L7zmItyDpTWgDuHQXy
T/rR/Dbm4oY+Xyn4b0eUbMpLxQ5ai+7OxVBEYpVMKubnF1gWfEKKuxBVY6HpNAOmwda9uZ7D/6mh
LGuH3ec6up1v9/x/54WB4cenV5+FdhrfFxThXWPqR+AaqOG4taiuvsd/3dRvakHMzlOtQc5wuTe+
rsaUjn+3dNy1M3tjN7fgWZIkf7cqRDh/xOuVNrUcrxfIuXKlOXfXDjGa4XFwJt3cG9nrUKuzn0If
X6JvIZ96q41VAErxofaC4L3vxDZI7z23fdY1kgb8Ys6GdUACQon1kGFOtWOzqY85LUaCEmtvktU8
xeyVhyKdIJ88drnS14GijJLfWDeb/tEg7cHekpKr+OK0hb7bPaujZo3qIVMiWDA5zm7DzmnV61kW
eaXENU2Ijc8JM/IIKBMvxt0ZJ3C1NngprsLWZi1EktT58Ff4BJXvcYyByZydz4MfETAf9WkCnCVa
ipYbuNupqvNqirq3wg2zVZAmV4Dxott4fW8xXYFT0+zZ8Rd28c1m23ko3xFY/Fy0Gp5xbLN7x+Xn
3NEp7BA9k6GNTpvwx7SEUY0nlA3ajtdXlhxOHsfMcRapybE53PZCjzPIBy8Xn/hzi/lE0769MR3s
PJjinnbCT8pG9tXED9yQiLZ92ey0+RqQ36bZP0lmSZ4kE+2WUF7CYHvFmnsv1uspdD1c2Htfd/0W
r0/hcWexsO0vCPs7DvftEx8u+UOWMvUPiVmK9VBfwMMugGAGd9NuzqDuwoJoTMQ+NlJIaEpNO5Cu
ArG64yQe/Toog+tOktM8uozC/iWeuHGV2uJ4IFpGmfBZ7MI+rHd3r1NxUeltc104VHrxlot/A8pN
xOwQm4qUFoWrI7CNjnxRSZua4J2XIRerd/1eDDK5f7v0Dk5PBRzZPzg4FXFEQxMTdyig3df/RKyr
hkm2fdBA4cNJJ0jTrfbpqYTYE6oD8NW5HSm/nwxgYgBtuxPUxG0RV8DpSLPCJltpUWhx3zLkL/sS
l7t1rr4FCpdW2KUPXg6PSLF55hHT3BXly/St8HecpNPSsQlBL6Bcxk86wlJOnpV3UwiJR9YKZmt/
hpjUybXvGdVxZ1K2nQV47e1RPuOCAvXuX1miBmP2Kdm6ZtsetBZEjEXf1Zjih2LsJ+g+c19gW6nl
pqFL4yEEHzfn/HTEir01sA1ORr2VECPQuoDpWWEqvJhHgsr1kvF5Z2vWoRCIUtnj5jacBzxW0va/
dEwH3Liac1VlUS1XrXLZvBVJrTMoBi5ueS3aKmaTWG+qKo2c3hQWIq0wb3jvlEjBnCq75LmRe7aD
vunlexkQ5CId6fRGZEiUfJ4Dagn36r7Iqw4JpCmZziV6SgaiwxFATcQnA6yDMtoYaWb7Hb4U5x9N
WizcEDKg7JIgrbCQd6mgbt2zwqZdn+ESF2/Vla2rDmcpsFyiXwDRLSaWnB2+hX2GKzKQU4GKbb5Q
f4Qpbrioqu0GBHRZElU8r4qD0doqMFFakB9w1jjUNMqFveQF6YvFVyNhwWKB9clM36ZnBs8mi3K+
m0qJ5nx99/HIlJU1IvM9/i2+TwTFk+ZzvIWuBEEFSJ9l5IaqwbPP/L/GJIxNEalaVCMNPc7XuYqT
r9sm4+6cvBRsiXnOSDS2mAEnNIV9tFi+xNNIZN2iTx+aHRBlYp0rbM3Kc30EjzG+oGTNu8ro0rjk
WJzOqyVSjCgmvCmWXjhIwl39y9Fb3qy8btGWTA2SRLSfpcBgvkv/nAKnUKsIMAnpTdLjI1wl+wQB
3Al1tDAh7a42sY9onZ9+ySlqwz/gQlF5AYJhOYkqdtYHW8ea/dl4+6Cx/uowDR/DFcHZSN7VpJfa
nMqNGBwg9HXvX82U5++/5+N9whk4qAKsJjR6yzDt6KmB8vkh7H94hkb7J6FrDO9EUDHipOuLr8b5
Bu/U/XMqUI7yjvHR8Lx4owihMU52ExxsnQpdVbxGX+rP5ZIStq+s+JMpflgaNoG31MSj9b621hLt
WOs1fTSh0lPo9GVtoIJGCqj3YHRBLEaZbAlIezHgcGAvoDmfCIWWTlYa7+esYdeR83Bhck+olinZ
gN2REmMR9A6YcykFxjEFI7KBoZ9PM1lfzjXYLJo8W5hfEtzTm0nLieaT4Z4dyOXl7fnWlyJQ7k/q
MOSzQ0FC06X7cIcuSfDgLW2tx1PrPykHYNUOCkisehN7i4q+3a/5ynzbae3nveGaL4FXkMdWOj9l
p757LvszLD+39VzFZBGX023zx+vsdg1MMEvFAMDdFL5WTki77v63xIMrYTd/1ZtS4aihbjeJDZFu
ljOPqrWw2M8dRxU2zr2Om1WBw/vqwL3Rumn/KEtYrDMV/RGQmwAsU8yFRoYqm+JdpGVpvwVTiR4y
RC7bhgT7ffG9K7lsI0JDG+lfCG8FzHofyHZVIIJLSh20qcVwX5bTgUWLJRrKWXkKoo0pVhfL5mzM
yuRFjfWtkfVAXLf/Md91lsEQsrlaahbyYQR0I4KEDEpUyNIqcOWwd1t4kxR3GZBwYOjDWVqPq9Bd
zGp3tq87YBxCNts+RA+r4gbwoUhd4yKsNUvOu4fOn5ekYCx12AkNHNqeH/lGnNdblfeuBQ/qnH8w
YOGTj/t9jY6Z77pwFxsIkNJ63Jxfz5kBQtjpwKJIC8W62UDfBAW8+5FT+L9Jy77sa4TKrEA8dqe3
hOWWtr+o+PNPF14Tm6mqyRY7lZHNxV0rUaNGx/fRSIreun4q94a8o1vLOfLWSDIhLuGm4qqTWyvo
qJ3GdSDA071fRgphw9COYbFdPGvZQrHTvpoOcSQKvLsToNALbKYlm4gKVhBg3X0t+GLCsxnaCnCY
JDVPiGMSxwOiu0CZuMyk9kg/J6PP/RzCjPtINW0qGpJ1l2fZpQlEcfmgq/VAKEQ1MgpYZUTVQBD+
nLdryZ14YSDwUplqlzXvRD/MG9gigOBrZdyWSpXPYAXSQHUZGC7d4GqYs2PfucbgUfqHiXdSKn7p
jIght0UKW6XEuBjzbcB74ZnsG+K6vZqcgNrYkdiBo1xDVeaLWIIlImkATpNAv97vDU5wjJGcQiPw
2w5t5CErrxMCR+KXVOE8jEj+TFTE4R7PYR/p2euWmUC4Iea4XrOhR65r3FTuZ5oBrLxaLXWrYhb0
fSWqNPoSx0AMpct2bznMpa0HFUG+K2MIjOowEZ2aw5AX2QucIcRmbtLLDG3M939AhsHRksTTH7QC
6hY+0Gsv3AgadfeEfsZo8XX/K9B1BJUuUnOprD7QCzQICXeBr3IaTyKyph6nvE8mPd/SrWcCSqiY
eXuP2+fnaYMfnYMzusc+UJGlf1Oowlx94Ddx1lVOl0HdmF2kGoGwjGDunk5FhJ6e6uYCDEua8lEk
3CDu7wzrvi19KoKBIYOUeYKkKe2EKPOyRtGCRGopj0IhRvXKZ0Yh6Zl5cGZqePcp7lu5VFXIaGTH
aGRs0Kb/CD0xsv9TYe41RINBfqmGEi2kSyQimzTnBiYymOEdfqz0dINF7xhyuZsd0/32Q8P6a+2E
vX2gW8UOz93Nqw1ejLGnsUBDscuxf9A75FHg+FuzQiCawlQZqMD0dEHa3HwwOM5UjZlbVDJ12i4I
Lx25WSfXxswWnNdr/XsLU5AqD4wgrIpPjKcKeiUDiFXB93RsRcqpTCeVkJA5O57LEqRfZu9n2SmZ
f6JZLFN1+A7RheBMlxOyLdlxxbZmMynW9omMTKNZSO9qW1cn8GHkqa8UcYH4MSq1NFksuNRq6pVB
s7B8f6QYEH9pkmDDVIIxaNpswDlsk/4KcGYnH9LqmgCT97vo5N8ytncpKpt1FI067KjXCAY+t7eC
8YZ7WIqpFN7a1CwcdVoHvTEnle7+amAPVmcLOANf1LUgLCCZ0HN1aC2QPoYdGdIjDK7mPXTAXySr
jbUsBP33z08pGyuqfKDiGlIpgsO6G2rFhKe/fQbYqlNH88UR4OJdpw+Bc6GCtVZzIL/a7kcMrc/x
/AcaoW69JSz3D8mGpC9xwJbPAoEJawITICDcDWqgNvZQ84Z+aSp05y6hhLIk8kI2HvKGQ12Si7J6
LLl4nPnQ/ziJR7Owvx8tqrEc4SwRNgt5z/QAlmhg8hGZc+AqvhD71IMDxhcK1xma06MjScV05peL
qeTEaGutoVSo1Tqi/KX0XQdnzUVgxHccojqF7NcSGfGO1JVAb0cr9sgK7W18LF1ducVVtpVjEF0o
qWcXK55GMmsATujMJJo5DVStgDyXA9cacVuL57tWdV6z1xjMpH1RRscExhZGoZhZeWrCgfIc8e2Z
cT7Wcs3dPJWjdn0hkZifaVJeKXod9b0vjLJnh5XfWDMRisSkRh5VRb1wYW5BOLkA9NCKfVWf7VOv
gI+Vlm13PqSIRxN7UqDogVt9nxp77mXBSsWGzcFCZoNKmyjC5s36QLQL0A1JVrO3rmdUbH04qgsb
B6/4L4deCxmBmefQD7iqXpCGpcIsFFqEq41YcbRTFxwT0rgQgrnWHj36pFNO0AUADw8bJsefvK9t
fMfajc5Y2pvehl5N+8q8suGY9CNfp1F/6QI+S+Ohb3+JxXnDbTL0iCgNxIdZvIBBOpSe6Nocvdur
1sZJhgh9/dXLh0LmVzKJCNQEbmSXKOgAGwLlodqoWCtRnmyD/Rr7humctOwW8i+R/TNC2jEUpLBR
AJb3wYrVNT5/KQUF0K/W3TvE3XAD2srJHw4CQNqb1HtO4i//Jjns4et8eHDn2AshoP5jZpJbvXdD
XNhKGA5pIOBnjh/5oio3S7/KQCR6Sn3Oa16lzicOX/okcIk8WnHxRZhUyhIuzVZD+hxYsmfVKb+4
VXMmxOjk17AMoSxn9Svm7A+kZa1sAOa3OKkc/JrS8+QtXTG0XjpK68SjfmHkWMabUCRdDCaNLnro
Be3V7ALf94ptXEW8dlQ213KUpXD4eY1nsFMGiv2qwPoGs5SFpv8/oQiepRBNYE5wlI+zlSTlNHa6
HPoTir4jOz4Bl4NqZQoQbZp62RpYyzKK+aMC9cvUVOAmMzMg4TRjswyGs33Cv/EXI5xNlfsNUEFF
hR2ZFcwlL8t/y5whzlY0Hp/lBuFzP91IwlBgRU7G+M6mT48Z/en0ghxPnyH6sQygphAzKUYQAXaU
JslNY4oV/XDla+qeCpU8fFmqS5Mr89v9jx7ROV7gLaVdMzNYSC784If3BJUGqCozbInQNAvmfDB/
ubsjPh04tIGkkt3z/bWPsKfb52rnQBGOPM9PutoqFI7xO4iqvCLpC8DGJca941rLchFdy7xNsuUt
8IYWB9DzEe5l2Xqg8cngs8BYQor9YcFTLpnUoCwgmiPYh7EC0iz9UJZgNJu35NJ5JJ2g4DXACvEP
43qYZo4rI1fdurLP7phC6o3HAE4z5GfJY6EuH4p5RaHOnb3dqzG0j6P4UMskIuVa/RA/7Ic8AyYU
oyArc45X7vK429ZbrHb0yOArM8yVS1gnGf3x+8SzwUU2Bfu7XJHT0CBYH0/s517xlABPYGbWu3nY
RzSTXxQvDvGs2ihIod9jCa3IHzXgfh1Ww5Ipj22bgy4QVE0vOIpYnEA19CVyyc81qnuoYzzTwmv/
Gh0Fv4KD3jZakjSa1UNRIAxQh25oZ1ghTNKrGqmaw814HH+3vixIKvDnyg4FoUH8+KYRJZoH50ar
eDVRvRdvqX/jn8Qvx+ZZDucKj6WQ7q2QmRRwBNfgAEiNnhMxVZOCofRTFoYWF4tmB8jx6JuHyfZW
GzZ0LE/BtykEt+6eFS8JYriIOrf64Aw8qHiAXV+VFuKxnzhDxUHLQCZZj961MbxauYdrlgq7x+eI
0ZOJ8S+TUsTzuY2dK5NUlBhCYM1vWkCxuQNIs13SGPUkpRxfzVcBKIxH1Zs6i7WPoFNurHaOJnO+
61avvCe+TySdAuL+b607niR0wvowM2gnoWoYDt1sy0hSwF1E4cEk8/rZZN+mKhnHOViK6uJvTAb/
cqLRPSQG6Qh4z/Ur100tFCsuVwmgN/8l+08lNROQknLAixvxHVrL0NVlCEJL6BmC5ubLOBj01gSW
2JH9WNXCF5LE5MfKct70TXMp94WWFnCygeuApXLw1xjJGn2URobXw+q1WY0RpijSCEUz2lGo7dRa
o9TLc1UFM6bMpUdtx734Fr760VcT+9os2g+Pi0oHfV+OzK2zziKeNFV6AvdROhD2vFSKwWk+csRd
J4Ez4pnZS9dm2PKIaAwNeWl2CKDPTHenV80of22L51mXwYAIJrmG5xS92NKJslHmURL9UhUQWVqx
DRpaapPNHV40QKpJgrnoC1v3nA7VwgEVx3esurpwRLD+V0Xdo0JQMraUDoU/g7oHHs0L7LUaqbsh
wF/6g0LMjVDnJTyeiEYONbOBRNvRV13pG6nmwd0Q0XVEw01ccVWtBvhWZNtmXOq7hHbE9JI4149V
qGNMMAZ9KTpx8lJw9wXaTRael7mbrOOYgbpbzkXrLFYLj5GQRVMdIssW+6SkQSmZuFBDIw38vfzA
fObXBl7reL2veYPFW4VNI0FF8pnlUM6TzkVLeez342kHNZ2FVNXaYLiNszPVJgDdOSwW2DY25DMq
UJzlZyp6+Vgfe3buTxGbEFRGTW8WRKAyxH+R1Gb4Epy3lDHExtqQapqJPDYGVbrC95kXqnfmsQ41
Pe3nYlaosVJ73C+Oui8H1nsm7Q4wsLMUe0jJadv09KKd5DBm/2bdhlGbil7Yuy4bvs0MqwWRDzwM
xx0byFWKW+J+VwsHdhtCvdELXEZZDjJFMjnFlzUCozQjlCZXzqnD9z+oJ7Q0Wc6LWcdKeTT3hKSl
6rVpNBL5vOl/zL8P8nHmRZb2jX6yjtfsT3GDrivN4Uv1XuL2+M2UsvQe+Wl4mTKxEaMIKWRIEfT8
1tnqqOIvH74vzfb7asLMqWqnvlUjXSrw738lmtaVY3zTnSMN5NHDACB37GKH3C+3KN9+WM5DXpQv
i66iiuYKVKnNiWoMP9/C7urtGt5/KRSxUFzdYqBXE3sqCfBqqF+1c2u7laobNEUjjlUsVMfnP3SI
cSWl5onuOBFhBDRw/RQcwwg8hv40BjaKVyz0ZPtMi3doo2shA3lnA5m88qhGBmwwWjNiZDcUq3Oy
UEmkqdXmD5Ix6i6yrCWxR/lkcTx9axnjq0zan1oJ2XthXcieTYYPr5ooUOSWwmLNVB4rpJ83Wamb
gGp4EDwdqo5UtAUuukaBoD+unQqhkO0BEcKrA1w4Wz7n0FFCz0jxIhZLpWS8jFLIZEJXrGsSU/1s
Epfc/QiRpJv3IXUyht++sl4b2eRVCem+ZVjJ1yuT0OPK7lsqEONnZYmKv2c78mTon6jaCPIhhyLn
0SCNEdWEw2x/4nGUWCo8VIn6UY3V/aRn60QCDVz2shscNsR0aiAhN8huIYuMoMtZppj4MmaslWmG
qJPXp0bnUaKPn4sNsvtUZB/Pk2Xfu1Et1JP0hMyY2vWx2rQfQmccPfMcf+JI21Of8WKYHGvEkvxv
CkQal3mn21NzxgQrkgSxxP8kdkYmaBF/X2M4hqFGisuHgzyybPzhHek/Qawqr1ruqTGAzmPHIlvf
kODSuuu4u2j638F+8+DuIzIXogAZItQo+KvVjb8RNzP+u47cyG4oCXk6Ds4Iq4rBXirpYFtTy35b
wE1ftvC4KhmcnUZbgX0BNJ/TcevOQptzvo7xn+hEY/Q3MY8s+2SKzXniOVdQTJT5eXRBEvMMYksy
oN0Z/qDEDmrx9Fb3kHXDrsmNl35JPvZEVY+ywkgMQ61UyYwSyKL59chbVfkgDCxn6iVFo7l0gW+z
6/SYfSDYenHo4ILnk5gPJozbsOSxotjGkrds1Z+Ec+TtWINXb7GbWGYZOrbbHB2wbFJ8pbnnJPxb
5pczRIEFfwnPDcdiyBXrq5rP76iSOfU+smgSYkARx04jxLkeSUuVhL7/gKMrrxAsl0msUU5yk/Vi
SCWHp9q6CzRZLsOrkbfZoNO/Pt6NRKvQpV4cP+KMiaF70zXITpZINGGlQnK5rlOXH1UdFQfGP2vQ
cPrf25eI90uhoJE1642zB76HRHz+nbYYGE1suTc9S5JRBQCA58VlnODyjfAMy9TPwSqkJ2jc6rMl
JXV7HBO4o8dxtu9grFKfdYLCTCypNwI9Yp1jSMEPFRf/3SfoYjUjhnV7TXoqY93xFWINH+ENHCVk
d4K2Bbfk2bEdjbIXe9nKn/cVjD3ESfVR44QN/DKUQ7pvndG4iQqS20iXoyhxFu88NA+NsZced5UE
e0JYD6D1Kf1gpDYEZBNwK1KlE33hxm6YrSiQuhClt3uMo+rXiW+42TYMol5culWm2+zelr1eqgWS
TCrsTRr5aukx1Gaxbf9yFpGACu65M9n5HlC28D4K32nAJ23ZgJXEVSZgnFTz7SwtKOHvLLP+y91Q
QOk2mfG86tXYh6PsrRgjnE3fAZIn8VckqGp6/Vr8nKy9Dwd86PuISOPh/4GXzoPc2aZtMtXxpiLp
gshBuRBZRQc+kU6KQ2v7Dql98DOUlKGs34edrOD7wTPqOLfdqvNAbfW9HSAjeSgE1NQvAUexzjP4
zn2EK1k6gPTrX8ctT7iCD8xsqJn2OSe/IMWjnlZOu6BlHmcSte/JUM0q1T2tDr3dExo2USGZrudZ
ypJx0RaXuQyquA658MMt+P+WTNL0G3V3RwsecAIqJHYEYMCYc5X/VCpmT4piUmLspyWHLvNfr3O7
e5+Qt9tWEpVfNXPL980pLIjwBrh2cY24I+dgCom//EqYTfmXioAjtvzOUllTz9HVh51WjvITB2Ci
AfZ+1fGGBTs9yMxzazzobO9caJ5kiGVMWJkmSHylCF50p+ozRGaNrQdbclGzfuZG6buDXe2wfYTv
WZbhkREOq/7wRorKGCges1q6wgcV7znVToE+Qq399DY3SiDWdOpLKvSmSViVCfWbvlrhI0SlvUW3
b8xEGbRpzjHXjIT3uZqDvdUd3kYXK2tuap3Y9POEaV/sDTWrMu5FyUp18S2jZ5akHaaRfiKgEA5u
T8fwnyhe8Mt7GkemBI8v4GmGxSvcpFoI5F861DTdeY0qd2VTMDkKokGGji0FSzy+frjcMoaZFOBg
XA+khWfDOJKhMDclx89ZyxnUTRiypAg/zbHJDGXKjLkP7A+jXaHFF86y4gCHLQDjyCCvTncKRZAh
NrF3hhdJ7RdWuqrSQUo0NEOId8DDQVH662GfU0FpSYA9zZIscWkC/IpTn9zaC3aKnvoU32j2aLji
pPFlPyl1AU+pCtH2HVtS+FiRqkjbk3YBQw9q+KQyQUNktTZ0HGF5nlPlP7RQHqBK4oYQTE09uCUe
l+RLqHG5zr50Ny0Abec0BbN3AIxpxU3gTupyM9CkHzgZ2xzuJLWOqH5/V97KQiwKB97FTYQvmfxg
nK8qkHePHRO+n/5H0L9LKQS1W9KGxaPkLm0U7RLmP++SC2d7VCy1i1aMRzAzh60UIPuL01CD8buN
9TZZRgFwrzVQEq/nnL7MJQrYaiEWc5ccrpMCeUT+OMPoPPtlVLsoRM3ZFhArdBPkIhKCv7GYh7ve
K5hoclfzoHsCauxcZDu3vJa6VCnLzaw+zCVTU+WVnqaAb4BT0QBxljxpuRGd/Qzq/YIf/4oIVKOL
az5H0p4FLsuUQRVD51pTWPAwyUVXgy0hjgdlvlBByKa23MbU5X3WNoLEPuinO7AFToIyEstOjfJ4
N08aMdYpm/rKwl/zbzU0sMjUMITrlfWQbK3ctU7r2OKXH57YgXgt+fdFVaSFGqlS2uhQB5317io8
mmlvb4dfa0wbAJIK+h8GVa/AKpVt8gbSIMkBbeWntRGw/SbrISuSwfZryBxd1XB8mTap2I40kX+e
S5GhApOi0O99QY5kDSmAMwJjYBCwjTp7yeUS2cns4hu5/tXWnVXSGi81Fo5BtB3An+6314Yq/RAe
GjwaLA+LAKPOSMAlwcvbnAIt75YsmyrkwslmUxH4zxgfX2JvDDqZoXW9Mr2CvHhojNXXKDq8R9xM
2FBkyP5YniD6ilX0qfAfwhDO8dTwjwVP0oWXL5BdMH8W2msg5dCFuNL9y9dsAO96P+PpffskhCsw
TkG89QqoNNkkHZzRv5k7qBPqOF8yp+TaHgMFTYlWC3UqZ8C0Xuf6O3UX0VtVUEMDmZzTGjCCT3L1
8eZTqwMDetmTWpCAQ7D2PLmUJ04gZIG8e4fQdUVnhflk41GMC+p2YbOqXDvNN5Ti4Fzl2HlWdDZg
whO+DfaHgSlK2LcDE+2vUQ/RLZ35b2+W2OlkgDDxByNNcisAvgYl7+phhDNv8g4TWhN9xJcio3DH
L1J8vG9qN3njZkZz20+7VtzZpdLZMj5FYH2W2x+v4HFVuROvQX9tbvrCrdDpIRKGcFJkPepRy8zA
vLrm/Ihf/TFeuNLXECEbtdyA3U2dOd2IhvSGFzlDFMvl3gmWrhTjTMRrHezilcaSZuq68E1aYrq8
fKlmbpTfSOBQ3I9p6x9E0zOqEMkNMIelBMWUw4QA8JroAwgyyIaawgQNcotimRXNghhZo7V+Uet9
qEs49j0bWsSuLdQx+50PAfF4nrYDYWy5Ju1ngWY+uAMN3AM6b2TN393yv7ux/eaxBulCjMHh02ag
SxF20AQg+HM/WAcJxKRmitt2yIxSY+FnZqN5HDzXkESTetk+cif9CGQYtS4BFYwSbDBigFk4Gzoj
W8kK2GhA1+LxuNmut48W6MEiFknno8/styiZ9t5u6EdyfKPtUu93jhKfMSpjOIM/QAoAqJegew9H
ZHnCtSupWao8QdJ2vVhXPgmbaU1IyXS+/YWr5n36xYV9yPii1id30Ezr7afD7dGE3dzOiy2BYH4Q
be4fiLkenJYst39mpMGqf1kuuZ8Pm7luinoEhCMbrdSlwvqzdBBLpppIQ2qw6Xm6deKVa14Eobwm
LzgGNRiA0Ya+HCcIn/MkpE4q+vNfLqWlnWpzERW14dxcotIC2P0rr4IqAIT0X4ccI7VhbYrA0PlQ
5+S+eMeR/aN7DActrtWGAr4KamK76z7Hgz1eVoaZEtsFEbOlTUY4M2ZC2/XjjXNqcGm6gucM+hj0
PxFbBFRnuRB+qWzfUjdcG7JIHJQqHPYPIjEtOmybOj12UJhkqorHcBuOFhcOEuK73/ziqAPj7t0H
q5K+66nS/a7fMUD74FM6fhsn0ml+Eq/wkDa6RCi8z4dFMbl97RpGpvqyHg7TWx1EbUPkury1gHT+
WK/fv5mi1VEsiohypvOqS0px0OeJ9zjwzaWkvwdOVlU7HsFUH9mUsnDCSDXYwEFxIoXQlUrRm9Ps
OtrAppV8UgvBXdbTFTbEBWf4RBYZ9vgu+IKHCOsqvoSB8sRW+3TwL3aD1NEAQtQ3wfeuR58s+oV6
TBMUE4cJ7DMSTjQ+CUs9/kvBhjWTiU4mtmVznot7ktt3+G1ICxCzHnwAkFzEaCDhm2r6a7/VSVv0
GR4eb1VEhFOYZtfTdICAAgMdZKGwcBRvVGIWL1Etj0ASQz7EWOhtpCfnit0Qp6nW5GjYxaJgy+GB
d1BX9MXC9Rvo+/tY9J2wE24/cRgK6CUL97KBVGcqIUP2bZAzP3mQ1SEfi2UgiuZyEOwjvbDsbZoE
YTeWcEhyszkFJ8t/a84SNHGwaIptbmJnNDSHBAnARKh50u6AqV1i6x6hwFciQT3AIuy5SSzEWgzp
4oWiRo/Y9IYZJD8VBrxBnwCqEi85mcJgf/gnGT7fYXoIcTYHlRswFEEbs4lcfSYTmsQfOnqfJa10
T/i70WiMXAbJiHl9RCkf8gMccEKPeMAs0QwopCf9BhgUg1Rsfj/Gn4Iv7EZkKLC8aCV8s+zQYJRf
ThlQBicw+3sfwlTf07FZ+lwBomA/766EZHOMaX8iIlBIpMxULfjr4D8ChlOV8H65yycMfsVkSO22
BdpBy19pxqwYJGSCROb76Fy539OSYPR0ADOZPYIt/sot6fz0aeAQzrZC1V9K/cNopATopfKwGI/S
Hkjb0xtz0iuyp4VezGx81erftVUanmw/v2aUrrXAAXi4BeCYGE5Xdh3vQoGqOxN3t9tGA/cO1Lex
1FbOFtJKSufqSVFSXM5ooV25362n+wuo7IX3FVuHLh7fouQiwED48nzA0CD8AC4vWr2q1AcIy7Kb
rANGWFO4ua7/n4dAxCUgVKps61R+aQI7fxlOmgga0w7vPHACJYTYqSOLkgvYHbX4iWNS76lKLc8N
E/QX8pr5eSxLVKLk2Qkohf4HbEWTkG76MAYUcBSU3lZBlXk0SAaiAvflRufqHYPJoF7hrv/yA74P
IlpsHNnLDHWqOLSutnmkSHuxlaOiWRpWT14vqvJojsgZ3VW79OaJPJvuDhgPCCbXn5cbm7l5UgQ4
PDrZc0HiKMWh0yd3tT72gOqKfvox2PWk4TGt5eTuNbRzRlqTXDs6g+EsuGWFhQDkjAd90Nr6JGjo
pp79RRDvYym9OfiQB0f+j2ulkTANPAB92N75rWDgrrDosudmKHXvlt/SpiMm/a/5CM0A4ez3YtAR
Nfw1xa3igqzEM2RcCkpv+l/v67aKZpSURrSaYA1cPHvDBZkVSpw7NFFLYF/zpJabD15E8UbBKg21
aQ71/RK9JCRNUuh3oIJ/VlpTapmtTP/efSnksoRa4DVrVs4mGyejXefpRcJAHp47BWDVqGUwmYT7
gX5dqiRtUEhq4vkMW+sHvmLmg1utNA6iwYNXI/ulthsLWiYmVHfTsTL87vKzqS3ufOLzROe0NmvC
HMKtwrXRTS83I+pA1annXeYXKidoMrzAdcKcWkbzUDKiEWiQBVLdWIqQDDxdyGsH3EXLXkwv6cHC
x+z+b+aWqAipdI+CAKBeSakULdwWHiMFkzs/8o4JiQ52oP9/U0Aso/WhavyZRVeFrudPmeU1F+hK
xDWZ6nx3yGXe1qX1gaKvhKHa4/ZOUFkqEml6Ms0itYhcM0zdeSOaamlCcfV5ExxCAmTWrpv/r6Sv
FM0aSMteegwgnuGWfK6QfkyHgPdsciGVJ3OPlgzW0fP0uifeDrjqrzNpEsiY8Tg8m4915T4NA7OL
tC9K4fOwPwfBiTQNdTB1d9fXFLUD6xDuRMsV5Ues82QvMVao1aLurqVgp9DsbnMyJops80PLeuRU
Jh1fs5RPi/AxitFKtKf6DR1H2kVIduOjzRXxX4cGZhfuHOdNwKBepuI8mUOAOSwL9hRMiTEjM2gr
eLfpVpTKz0qZQaFEyRb3qCdl67zBbSvaEkgJjImHf6K7J4c0j8To3nMNq+MRh85mEJrGxBBuwwVP
9FSR8PypJkDEgg7MtBCtroyEL9eLWduKmISPhxGLZBSycHc+vROcBPVO29mtmLLqaVwZ+pZ81BG9
Zev8BUYrEYAqOZ/kq9m4VaPciN/fFLFrh+9ebO4vXHMEoUGPaJ9M/z5NLAxuPdskkgGErBq0ruyq
Lpg6ykp5nCXFSldP9aTorG5MNL4z0cz2g+Ps4GSQux6rWX79Y8L2NeVosjw0S/E7jfcODP1uRJyg
36/+4EwiIxkWb4x44JDyRcaDD4IPvgIEc6SNmDpZ6KFIuSOYlJKZyJqwYtzOsGH55AtzTa/jhdvH
EwwBUOrlH2Ko9yn0ZcVV+wj+yfzR1FemnCDj+tJyVtq/g+pN9CDjPVCmNZ+3cPEXkCRMwNPLDr5W
vhmox9vRCiwcEf2REpVZ7VO28TgWUQ7IHhDzNeL5WSFrMI9Jz2SKQWGuVzuAY0W44asDQVF/CVFR
3iM4bKeQuMBR3XChz43OEdRw4vjfT+5085imbJ8oMEDj4sVQwrJ/bj/bH93fwdgYL1NTpqv/zUfV
nIylxWYyIG396qRNgT2G+aLCVy1jBkLvqmEo1zausll/8LKAi/MoPxrIe9xfQiJHWlGTUbrId8L2
LCYflTmFkSUicW8/vsp5CKFHIJbNTv17nJSy85r/IDvbpPVJC6WugxbQYdBWEcmMXmpA9X7vFGj0
APhh4byUDtGFsuQ/HiJkafar1DCrTcyIsHK5tntCYmS7rXQDusWit2MQjqLF4v61cSYVteCFcJvB
OI545a3LXPV7CltHc+VBuUnVOpaZPVteh+lrxpQ/t0y94+ZIizJVt9CxLSbZdzpWunvOJ+eqRc/S
XClOaib5sciqkpXoPJ7HklX7bNQT2CR/F5SC8ZRGFrbu9RtCUtLZu/qGlarTSgo9Bhyv3gS/3RVs
Ms+iFygSi9697zIO/boHHA2JabyQi+PHGA3zkJGuwcIco52veUyE/4+xE+jz1jnGyETKzkbOoqmV
mLAcMf5aZajUacflHHGbQPgT7HbCRxTn8aKan8bzMjYJiTskDpRFL0ONiHW7s2rf61BrspgRzRzL
DJT+JHyUA0iBkqSPdqPI3IbSxqz5qn1oM+esBLEs2nUNcySjZHXL3GhK21v403op1q1j/ZUuc37o
ELqHfHsz2s+hQe1bZOk4q5gD+q2ZCo+7docfbB/3QjlM8ZbWZjBFKYMc20Ed/oAqZWsPrBEXNJbS
7RYKhs+iqAjRitY1j8TZp1rUcOxPDG8pKYZCNstL1SfsEJ/zQgXMRai33P/s+WlEM0S+rzlaZJ6E
oRFFMGzLZ1xCnUsD9o7WjZ8mcsEbgRx74NWRqgW23I+NSWfQD4gdGtTOY+69mQmg2B7j6IXlrG/t
bxcRIQaWBnQUwY9Ishld93l2IFAytN7yHBX3z9g7Ayw3PhmiSSpxmv7p9zNTMYml4gkacSIbX/ak
E07Uyt5tgaWifRydBBM1s7jD1TAUnn1huE6PuiFXd2KFjLwDZ1nvuixItRMZVheccthdVsU5IxNz
cGyatmonyoXTFN3yt/QLuWuGABVAxwdxW2KPXDhiSASRkOXtiRwFbNSLKdIwPc/x5bXFj4VoJUyL
GNdykFg6GM9/rsy9KvHUXamaCg4JyeFjptwmb0+Mi+rSUGueh/fAw+4CRMmlwB7+txwPJ1ncXCZH
r0wz3z1KpVTBwliR8kpufRtt2Q9SirzWnCE9Jm/Bq4MiJgFu5iLEa/n4TmbJLp/1khTC1BeHaT4/
fBx0O8GlbNjYwUzC6Khryag0amuvy6IYRUm9N0OaDgwYapiQNUrOk2SR7WkspUEFhzcIsmxT2t1k
IEmfs/D9PlWv/JtikS//Yza2oFRoUKtoFr9q1infmdK0owDBDMBUyI6LuxS33ilOBqGAY3VE2g7J
p9V4Hv3uo0ri7tU4IPczDej6x+OhcRtIlF85hUFlFXQVLSJ3XNNsLdQ7/hDm+NUfrqbXYI1VTbPT
l5pG+2ovVUQfz2O1DYDI1LCMFiqvYkqKOG8cdALmE9RFH39ad2ML+I3yWtjFOUvBXTMo+JFNYIC6
jc32o7o1ya3kxEwlofXD0v+B2iPbnokShtxh7tchHInCYjfjK/115ITfQReeQOwiVuydvBRFRZGU
7U7LUbN+3nnAExWTROgIQdjeJgYV2PCWmDKg3I9U6zg3UdgKi0k+40kaOfERKP2l1jzga0b3aL2A
3iJWzNOFXl3ZOvG1xZei9icT3aLLxYLuVfpjyDz+dHSwt4leDCxHNa1q7X0cPp2FQrwBr+PGYLCr
x6cFO2GzaFTSG93fF0/qN/mOPa8ofUn/2egQV1vZHjBx/GtX1GQAj7PBeJbxaUARbmm2achA0+mL
P/aNPV/UyfhfgOrME/UnI+GlrUNGvPIR8bBZFRDDulZVux/qIFUSk5pa3FPeg7m5644uet96Tl7U
QpSv0vnRDXVbecchg2slrNLzui6cKcDsdvXUtEesDXExFymRik/wJsZlFZ4eBOxdPrCuBA29Hkwm
3Z2I3X1zyl7RkZa3KTogrjfn9JGCC4MDxJO68NHuFyoOOxKBlAqsqvLl0/pDlNgOT0gs1h+j//46
2Z4riPy7H3G0eMxLuaDY6mYzQHKJRts1sKAue82ZK5y4wRbfZgjQeALx38XklTurG66yTt4+kw8r
3hrQgIj6p+Jy6HrkOVB5U45XS3tvwObYhCf6EMfPSTUzX0UdzfRkHSukVB5EWftVp9s/JbaI2g7/
VVSMGcX5pAEXMxgTN0jFF9iR/3FfnzbNIIE92BWK5b/vEzsRyxYgfhpLTMpb44oVYMrEaLklq1cl
AZmGYSnfKV1CgCQxjE2ZgPKuQpicGf2+S4Z6lLJ6fGTa0jHncA0ouG6iJ/YjuYfjwviftvWIewSw
fNepvEnwi9ORQbR+gC2w7D13KEWKrz/zwhup9B8Mfq3/hshAvy++muHUSP6yp5Jc5BocgyHb0bA2
JI0x+OuW6jXDDc7n+DyI6YWGhJc6qYeC3pzD83RFErHqLwWRyrQziSly8mlikF4sX5fH+FPBoi4d
0+iWsjZZpHskHFZYaXIBItH9141n8sJvp9YBTtJQMp3/v2u96pXE40wWItfCZq8uWxTBcqfnTLv9
Ski5vWshspirQYDaEnOOODIhUB76u9jGmKb2hB7HaY0G8WebwGrdKHvQsPZ0qDn62RfSk6+9wnMA
QKQI9d/873x3n7/Toobu4KMhylkA9uD8Al59gIqxspPzhEdqvW8xHDdNox/KGp0IH0c7Gpj+ax5L
koR2qAA9GfFbTSXjestJG2bCuPonN4ukeey+RWRDe9HC/WjjFlGoteBLlNZsX8VzK9Vt5cvv3In7
TD7NASb8Mc8YmZR8gTDFwheil0SZdByRjqW19rEwWRFTyvuoCI8xXO6s/7cGML9UWYIhqwwzBN4I
XpOFDIwT1O3N/KU2PnuIAJ+hdjn14h9tAMsUAinjpHdjjbZkwCqpX7e/fL759RBfJyJXtsb//432
jSgfESZUFSDx+0ELuh4vjeyKEB7m1D/cBZkF7cUrWML6+2N1cmtmR4shx2VJyLnI0zLHUd3JiXiR
VgFoXysBNXFA/hnk3Hqiz+rvSOW2BGvkO3p+E2SA4ckJ3r+1NU5DGgy8v25c+aEWWcTZvxgvlEOZ
Y48QbB0UhCOig3s4zw4um76vA5dRfKfKd/mbTlDVD+xJRbzKThRui3JFkmdAtG4oDxKkkMqf2tP0
nC8/REa/zh+rdS+euNb+M6yxsUgEQds2wa2mMPzY9Zgd83DMioGurysz/QZvQGwwIZ2wYFCNMH4B
gMKAfEHO5pXxQBzUgxvFiqYkaWLgcXQT0rBs+WowvzssZZLzEMSxYJHErPN1L92PPtiFdo7XEeNE
zAYv+F00G0fI1cTCZwM7YRYSmd/FHlhOA4eUc3EM7Syx2ARqeaYlxslnGYJaUN106AAUrmaRcAwJ
NPfMyrsEEmi8kYkZV8xzxfJHAgBNK1+/L15HE5Eb9ffHM2jEkwESYwFbMkXYz/tX/GXun0eSILRY
L2qKjDtT3OyKp4uZ4pqPUwIlrL3FGPibZfJEz8I8cJP/8W/iB0MoAf+ljqMGB0Qs6M6j1IGVEfLw
DQ9PVTNJMv/ZvQCOFmv50nD+RG9caWbAbFz0d5z0/fdLnZvV8TqO4tJiUXElfl+eAy0mBWi6/9bC
jaNpnhPS5lPHvE5gN7zcXb+BXPOmMoDkHSt7KXYzDMs5WQwR1xC83grYqfDEihqSRHdVCac6cstu
K5MDAIoqmEQo45mA2/8pPJaYwRGOBRE/OdAntvKK+WPNsUxIMAhSGGFPNl4d7mCH7XOlBSFC2qBA
FmtwLJgs1Lkk15F9pAEWvkhEPWySGJdF80WOL1Tj1h2oGEandxZUQo5d5opCnzy9e3DZXGS8KWVt
n+d6rpxZhdsLguLB7okc/ICO00ya5XDpVsKTIjVkV2lK3LtmsWmWT925T+RwFAX7CzYagFNkPISc
QUFFferShKHfnTA06a/7v5/9YZSgnxdKi+iF2QcgVbpTyamyEOzwEGVdXI8fZxvFoDm+gn8qM/yp
X/ZzYDNvGTsz/DSq2yHZLJJRQS4cAd8Wc44ZexZMq39daVlst3SrjeveZdRf/iUHh1lz9bANkNwT
pUBQ2Kg5xygwsHjjn47c4OuisgyM0R3Q7NzsIYZjzZoJ3pHkvhmUh0LrN9nrveui1CufszzuopL4
mbiYVLzrysXEXUQf9MfZ2brcgXu8thcqaYJazWpvxObJZaZ1mkMyDDdliH9Wga3OeyE5NQjoQTTp
Dx2+aJnKqauspnxN1T7ukSqvHxzTFUw0U8MLR0H+ZNZ5u97fftTjwEUW7SLcHPfv63WIPsvzaqhL
jr3HBY/ksfkx1wquO8HsBuxFZEZJMOR0RpF3LM6tDZbt+Bxzte4+B7C6AWBGeQn3h1aeKZDXkUbQ
eKEwhbRxQssPccRSV9/1rd+5mnIxo5Qyh13N8hIN9sd8Wp5/qcbJW5Jf/gXIsEOnof9yr8QA704n
hqIRzYhpMhnbvVqt4f417e0+Khl/N5F/SnUJc+DgkOf+MmHhEPXHJQQrPmEJbjqnWK6beVjwCUUy
IqgYXzOVSTeY+HoN5SCEpBMVGI2dkqadUicSCcSk7XoNQewW8phFaR7sjHaSyp5ooHKpZ0I3nJDu
jIwJ7Lq4+CR2yj5YkI7n+Qr3DzxTgT4gkvy3gz+3uCejrvdzjNa1iz1oirm4BL3mwT62WtAeXQod
bKBT+ILroEB/P21y6MFROmCDng+uZQg2Y6PWBvqW9zzSCmZr7JtGmSvjryee5BNQ0jVhp7M4T6LR
CQArwuIIG7Kw3q+lKPYyRcLdmZFdoPyW4MFY1ILtAcEqGgu9W6rdDbF0EwuZu8y8u65OtDG1Vjg9
mKt2r69/uGPdK8HncGE1AqmyBv+ISEDyazEkBqdSgohhcZoChBmW1VEsNWWAM1hxpM6d+CiR1exd
wE3ncvOZCuTyiLC+Q/OOwr362j6rCvV+SstSZFyv9d+s6pZgdLUxc1p8Dyh9teEpef/cG0ebuTb1
jA6IYpDSi4jY9tYftKopX6Rq6GWneqTP27eQ/18tovG6I09b786xGowSbNZyEkWOo5eP6EbQ3h74
Q8wWJT+MfK8KYHH2IgfuiW+t/Mj0QU0LxljgGL14ldhbGUG4XIlbRM4tm2rU2ruPaPPcJsn2KbQF
fzlhD77YDq6lhX5WIw0iVV14ZJyFHeWlYhnIovSlugWs88DOVt+830Hc9N3Q9dLVfY0Ws8K1Qcje
jxSWzo5rweKpdegF92rt7y0aFz2NhTVKGDqUbhAn/D4FF6tVJNFbGgkFP8cCDzYHiOvETCCTMl0h
TsWLk8l8IWvxmRSFNPfZcfYgE7AbdLCKeUtp9/Pq3Ys5gNdWIQGQ65/r5eHPvb4JqocZU4LmR7oS
dOO31+xRtvCy9COcgz7lVfYMu+xF2K6lROJleIFslP3bavOoN52Rlw9GlMIcNyMdtGksPJej57dd
PoCwWYXEN8iez8tCfV7gwXT+xIQz9y0mUASsDdJZh9F/5/9BI9YYyudsRGUxuFpkP29Q1CbVEFNi
R4zpgbirXbmcA8qWSOAMqUNJi0UTNGrFdxpFCBZm/EtyC+rkpFbIQM+UFPUBQ6M3nf/3QEFfj2We
w5zuhoIkNrzgGyf9kT3aDDxLap1I7HzqV9A+OnoyZW3xbtV+rHKRkTE++8YTnkR5eolO4xxwDZFA
YNX9iIXTHPwF7hFX0bXdqIjsFff7Y0fkzbSU2987CbwNzcuad9HTMswvRrWLYCdY/fBBg+TCNdEV
bkPfl0V/ymQMYZlZ49S9SMK4Vo+5FsFwW3jLpWRiW+v0i4dCMbSwTOgiVrb4ogKnZ+hAk27S4SX5
gmDaBUwNVcrQYTSyafYHjkt6hOPV8OBueN8fC03MqxZj8KezscVYS/wqJtukaQzGLwAH6FXeHDGq
gaG66RxTUtVAaLY727bYQ8ELO4w1MJ6jL7p8kNmnc1OJJTtrciRHqueqc1kI6NNyQJTqgMuWlPJl
wQQe6R/gviRBgZD+F8NSJD8XL8fJdqBBusbps/LRDx3QEV9iFyIZuD7As+H5hxDMrMdhsOdCJiVm
f9+ow5M+y9KR2Seuxt39rkSzGFJWcIDOfAWmI9KcFK3iofgCENcFRy/b2PfKiNQUY4rfeO7jbf+j
1lmxsrSnxV3pfEafwqQ6XWf/ZhqeI98Cc6NqIBDh7NwZD8xw4UdV644g3cQRlKBhDzE0/anhKRsg
gfRbZiq4+pykL9rWuiVZFiSOVZfXyqR/NHDyDEJuvoqhpM1SnkacmYK0rh1BbsanbwbwekKKmtyB
/yaggxuje3suWJ7M/xXnHu5CI5k4FKU4RQYAFi3n4FH2XQvwVaJ2rsRhhTojthkO9IrY9UpyCY8B
x+XqaC8Q+zGl3PYzp3kf63IrYw1V3TSYuxegwdC7AJWUC2PRuE7879Yeh1unspAJo2ZM4d7xgZ2N
EoFqQesnLFy77lbCPX50Ztr5fi8plKoSlAvT+05R0sz6MYmZhsBIhwIoMIXEIPw8VtAOc9hhjbCq
JE/8xwsEMCKcc5Q069GDFNKqUrfe2PKdqw3gGfjYsVSZ03vGOA4Z57v1fdNY45DtNfxcNLQbM3AT
rr1l6RbaTtKl6/rlL7/GZhMKjyCmuvBeZMm2JuqwuNNHiYAFjkwRHVpxyJcTH5b9P1RrGhoOUf3W
PIjB6tQx1EQcWl/QlWPGNGKO/8Q/RRTAu5FfCzH/ZPgvZcvVyQg4yE4qTn6EAkin2Ey54YhKTegY
+HcG4fygrA0kt4JIUH4XcNkvy4/PS9PWyWmCdqEIyXyg4Sw557V246/lkbQf90OfNJO0cJ0KOluY
ueN43Q5U6jZWB3RnkOHgnS6ZBmq6b3UG3kgDFki/dDtG6M5pJu5EG7bFjeMlICHHpHJXX0N5e+re
1J1uAhd+N6Wa1z2G/nj1KUwWizQ6RDYbvWNud9ISbujA4T1OOZTll1X52MpDjKhJjQF6o20Nck+x
ZhFDj1MP70tdvErcL1nGHDu5q2ttHhGDp2vUrrwvS3moSgYTCK94ihyP3Q3xSvUmKV6LL5voWif/
qbzZnnQ5TtQOnvbRiEyufBZnSfnuQYsxIxaN8k/5ZPYGIiElfbLjX1VhtdX78vNBaBAKz0yJHPK+
SlA6FAkH5PLlL7OqrKFhwUQD0ep0p2uy7oxy93wufhIWtJ6krMk3l6OchUqre6kZDVlwI/BL5mQc
ZUz53AE6l8qGNQSAHumQmHQf6pctUAocMitz8Vg9lCaUzoUm6pKI+S0FKfNKPrySCYLCPxlSGMc+
NB+FdU4exUCWpvdAcF1YviJWtjAMEz6v4klaF9E6I6wOn1kKWVrIZo8Nj7d7Bu2CEK4R5BndVOpX
PDbt3qbUmNyjOCpqY4XfvQHAeNDciGQ94phvPEGizal6RILi5Mb7PM3+Z6be1cgeUHopjkPol6wZ
XbF9ugSs416u1YbMoA8FqSXFJkFBCq64zvjVFJtTttYCKIV6+tVs+e+GWq11ie5b0o1if0JEpQR7
69OOMpgrJxConcV8MsbCkKG/hofVzxh0Cr1yTUZrvL+yJYMCkgjpQ8KDwgQy5LqZ4cV1xc9VMyCk
jK4zKOcIN+PNSRr0RfzJP7liSlKrzmOa165YcCWfzJyCyVy5PRvSsFZtPf0u07LAlFxLGQLvK1yY
7jG9obpGieNcLrjVLXDq7m4bc2aCRZIfkUz/bd+IUEe4XUC1v+TTAbI7VFBmR9/Wrybd2My+k42M
V2RGSYYWLeuhd6+rf/NPkSpev5ryC+D/nzMMdP2senI0duWl/kdeAn0Ddi3N7kY1Ulf3QcVYEp2n
LAmwz16LnmX7Z5BvbVvKSJOk1EqnFJ8hrDojuMRvjNmWokG9bA/vplXglUOFT4+u7hl52ZJ3XHEV
wBRFjtRD9PJjh/v7YE0T2iHup2sw6CDWa2AUVNIG8oD1xXDTyFhz4eTkbqdNpuuYb6JDY0MHADKT
j8kNMp6K7Fp5J7O3TXMmoIhwk90H25KiLPMfshM8MgZZ0D0W2P/91W7Tkij2Yf9LSlwYNfv6A2tM
CtjISX1N4bzV2cXlxNy5LCCos81yLwFJ3Gv1Tm7oiM3yormajpJxkpfaCS6V86YcZDpNIdsvbBf7
pvxlXVuJxXsIFreOguJKeL5pqtnIt3haZ00X5ZxpKgL+EzCxb2Elvo685sLIHgn5sN811BCt9vwj
kdWCAG9p+ujqbjMCPNg5oaakncJqbWCdh3gkOcZMuQcY+fSEk5xbm+2BuhJWhjr+JLBxcqKMuaFk
ZUcKZVvuf7cTgFmpEKxrAvEZtg4R3EBTqixXLpCYWDfZwaTOzowkeZ4Gw16AYjf6BtAB2uZh2ySW
5zjDtxQlQebtjkDGesgsWAbk1rMcx0quw2ZkODjbSvF9H2K65bhLhmOTOnDtlN9sAg3a6IKacIRx
7pbcyG8sdNAGT75JLZHAiKKCPZKPlm+ibwICLpFdQH+bZDo1gl6ldD1K1I+ZKw2u7Yk9UWkQ2p39
7xXXVmAbWydq1B6b+8FcY2Dx/e00Rb/NFx0/6NZaq3xNEV05nNRVQYuPC9dE0qonrKGRk+jDUa/b
0uftlzexKTicQOUxI0PRWKiEO3UNfjWgUr299r6ouIyIWnaSQPnr9/EC8ml5wDBX3YBFrQJOP0nN
wsAdK5JAnS9W+xjeEFSam3ipRCpactqULDmhG/7xzAuyvOEWGYCsIDMPM2W+cjOPKZZp4Dgr08rX
WsiayNBtrb1dHMtgM3NoNrz9059ybOfyxMctVs3qZIRrwgUHdE1Luxo68pIUth0augV/IsrGGL/f
EiS+0KrdXFVKuwbK2K4DMU5ZkTo+6xjrWarRGfwyY+7YiShHTVxWsZxjznKY0/Vll2uEwsyOq7qb
YhNmNZGm7CBTtwODlwc5pnCQDGKuhNOWYwWpciW8eiKzjOrfoAhz1nmqZXKOq4lGegdZEzsVv3xl
2V8VuqFu5nEQD+FyL5wcVTwuDsqlmEBngeGyzlAY2gNEWMx6i0tbs9gRxFvodZ9lknQhLp24APHv
0kPzOw3gap2W8eD5ePbuDE7Ucrl0DLHplULqVwOPZWdLW2GuRG2AKtiCGfgOEVfI47cMz/ITZtfX
yDS6DqJWXcTJEy0tWqwRSfDA9jOk+MDUK+captmD0bGn/pRxTRlQvG+Xp5QrsibBlhSfP7dHpUdN
1UXzUuyrkoij09ZI7/TBBlGgWtC0JY8znc1csOoaU2+ezb7XG/RsDuSHHMd+ntOrc+KaycxMvDoX
xMhCBPiJ/4EjLK5zsj2u8AriOp5SwaWef1MQWjSg2LC9TXxVJtMfWPNbbf/rCTQIhscWFXgwjORN
jDl8tRZaL2D1dgntkW2J6ryGgig24q4uilFwZ5S7XaCrE8hRR3OjBd3nVfM7b/CPnV+rsxg7H075
CWTc4gxKWhU00hJhQFNFSpj3tHJJCgjXhC2Nn9VNGnuXrDRGoXSeneNGKcSovoSOayAUrIM5PMma
OLJpRiinvD0UKRBL2tIKwF0p7EQxwBBdJf44m12Jgxowlg2zZOwUqwxm7pt8tvJa9RQdY9JQgRrO
/ccxFubUFi9uHSDIJg5r4ye92fGxoDBnzYMnTkiifqQQBUAknGkMbOHoLQJ+X1I/LHkzLvouUGrg
prYrxDCkXi27TFzHMpx+tT4XRiu3STv1F6vjOlF2VzFZG/VLurHA2i8c5hFTD6ciQza8e4Ej1Wy9
WSnXmprRvZ+zB3177r3AKUDvCGDI8q4uEPEmRShGptwjgHO+TYqQ3XwSOSLDrdbPz1q4O7Ik3iTH
YpuOf+jaBELez6TREDDyfPNq0+LmR4pQ5OJ8hzm4b7Tp8k913r6ZxWeT+pOEku2d/TW2XlxaMCLl
toFQuJTnOyO6vAB4qOXCZ0UPXuPWzZ057+cYxROyoQjoSkaMJwhd8BEJmmPZr2TkKSstRlho0ynu
W2qo7pYiEEtEW2dZJXZenvUmG0TVRztw8W7/Oj0S4CPj7/cC5B4eqV8YUakqDHa1zPkETHchE3zT
pl1Gp12NSpkchFw1znCw+mh7KDZ0GMhCfS6oHDAZmNZS3WjNbHOIZ6FB9XccgfcbYLLmEPmyim6q
CbD5N1eG5f6/3UTTy/aCtklZ3dGXtyDyy0zFzHBk8q2v1H3QgmPNQRoGxXnTRC1nQB9vcJinMa6F
U7AlnIh6LZme8wlp2qimFrX5+scSPJttSL7kJtfms7RxuTYEa03zv5DN1gyR3FINtutzbnPAM2FD
cESmkJQBLzOg8HwBXi3VmJrSIeNTYf5Y5fxvZ5OhJimNyvFb2LBNKVvXzyCwcVyak0jf53cKl3ch
CLt+uBQfwglY4OuybTrClBz5IFJB6kaJEwa3VXY1rgvvanOw/EFSgtXvYwtZ9hb1DHsapTlg+8oZ
c8DJs6qWTAnYggnqsHTmVoGAfF7hKn4edlGDsywToiuA+ToBfx+BQvvtQSj4USifIgafg2e9mRqO
iApbmBNnsB/qVnPUzIHCH0mXApeC6sjCuh1MnnQWVCwc5d5eYtpeiS/wWhd/4BgVBoTfABy93dnf
508h5DMlJX8i+IffSKO16K75merrqx4/6Nu7gUQOZ3ESnNPxWXKIngu2sW61WgSSnPFZ+qagFHsV
YH4P+4EC2EeHY4scNv+Lhfb+OSQZPMXLzp7G0bPsNmF2ilybOv1pyxUS0qr9WBQiTm36SVobNsRu
Tpe+enrn8GUTq1ILh4IRXOBgHg1/Qx0eCJVqSXTR/DukMx3GbOAUIuzXpPBf339EtzQIGGNOQRSZ
URBKX1zeRlczF7nprbRCb+j8BVOuxNPe2oTSAeShJl7ZckZUh4Fqo9WDc1Xs+SZK5CXZy2U3nE8w
QMk3Mid5xZbEttO3IUxPG0XrWnq1033g6qBGtuNjbJ7RzXWrPV2+svipOAKF4KJbM8NVFiZTNCLJ
ox8XIT5JUMlo2LAaDjgwXwOUXjswbVHl2CN2ir1lJTageyiFAoA/5g0gzLNTGj6w300h3aijBOjY
lmMOqtJA8544sssfd66Tw3EvWU3oYXkFqq7C/qM264OWnbxnAqZJjiZvmfCj9hD+t3TNaamKXwoK
VUKYiABd3ChLTcEdnhmP6KTjzR367FqCzbWA/D/2Qf7tCaUxSTEVE78AFLjPKbHQF+8wAJk5vpge
G83rOUzgLSfLpNqji+0yzMBRZF1tMcEqEoYt2dHxmSwPe/TSVwhRgZw5etQb0T3nQDEBwdAMXRJt
SCGkUYyo7EQlkk43eStxbhRE0hgQ3I0W8A8LdEFT/gaNFVneNmCL1yyScj0+lRTa+Aa1E+RzAyh8
M0yW+r8Pz0HCS/3mkJ3YssoKC15ZW7ceGwl7Gbz+MPAqDiP3V0Y45ElvQ14S4fBm86SgiCARSPK/
mMw6lXpXcjdTFSJ9ij4LM/ckLu/zqV+sqD8/Wf39Rkq3Fg/jweQHn+tzqaiPpVmK9I2CY7Kg3Mgn
4aKb/qOzUB9l1JmSy3cz3uCv+qWbXu0/tJoIv8kgLgb45beITyqPo9E9OW3N8PeUA+RnTzw/SvNS
BHzazd+tRipG5+UkvJ5Mf//SxAuC1QlqhwRanMqYQkbH9jJG1St09xzdDuEbRqUxBdmg4nxZ9Xw8
P3lcDN4w2PLxLMs/iiZCn5Qb550sR/PPm0/CNu+OEyo2IWUFFBmCzXPTrYrJQ3WSl3kTyiF4z4AE
fnO1NB0Tnl1xpQywOeiKJa6JJbd3/4+pXYmjs9Mxaj5egeizzljgrUGgbImONH20Wk1dOKBjU5Lz
Ydnl/763YXrjb4ndAxj6L8n5BF7naZ0m3LlpUXbkuVe2FHz0l3TH6f+hp4Cu9XL6NZ9R4GWOPmQ9
NQDVR6dJo7iGbBRplHl+AAbQk7nhkJEeImT4f7bue0pWY6KGWrrYnuJ1eQEp4lwgtcoGdn1+fzyo
m4sw9rKoj0bEjnsPnjRIU3pZB5eyLxw502/4sRVVHD4WM4vcjruBW9uUDzgm5uaLLctUCek2d254
oDkKP+KPztgNuA1qwRUCIpg19v3yCvPUXmCNC9pq1OHcDdLFdL06cq4Nhaac0wauLBA+snm8osDY
7xR48zwdd/BGT1+WEZ+TSy2SC1hv2G2J2IFeMHt6cly8F2XCjzsV5JQp6ZdKYKdRxrtgfuiIewaS
TkhffGXdZ07FPGl07688lOLkmpkSwRhzfuEW3Otkjh9ekGIPL/o9Xw3RtVQd5C8z11AP9vx6Zur9
oBY2tnEhSN8qhzVJUMMGII3TLqMBUFQ5ha40qdrUP1Yh9J/TzUr3pPc5VJs8Th94SeFFoj0zYNLL
aes0+ZxIFhu4Hh/dV2FBRBmoRCSlBE+jHobM+b0gQ4VWFPD8Sbe7tQCPdjQiKntVbpRULRf9yaKy
ub+jwFFza6yskuQlSI+pBPsNxUEo9UqHM2xQsFcLApcYtRnVrg29g4ej70C979ZP+zQBRttJw6P7
nywJXuyOGdfQrAVpaHYVD/tNamL3q4XLpi0ALC21LGBI69XsJ5uzRsgXyD1CfyCpHsbf0EVVPpVF
v6m1W+5IZ4WQYtQ8ROmtwJ1ytW+ud4N3tOn2LwDmffAGZZ5618XanznFLon6GeCyvPHdK6QERNa5
peiu3PCDeUS0udt4czTY5obeVLkVVPRJm4HuC4FjogzsdjGwF69XhOiVQM+zklq0XKHLmPlQe3Fk
KRyiwwN7DgGrEnqjcRiNZam8bnICOy0b4+2Zop6YYn00zIqhM0n3nMjONe4+pBlnYbETLzK38iSS
I71bKCcQ1sKQv2VeAYiL0cxtU7Skrweup5fC5ENh/Q29OjIV3391MH6WX6Qw9/OYjoqDiTIlH/kC
/y/IQ+HG0m5drkofwz2p6cq/Yj+iDrbjmkSRiUwpNH7c1S7/e/XYGdGTw8u6ciwzL/cELMdJNmpi
wb5YQveS6FVUHf+x+vueTPCjlktrBmNHIR8kSWQKMbk4XF9sRkscIhItrDX1nXs2ek9xAf/RAKdL
boQ5EDmN1sJXA/zCW/DBjIxi4KtyK1290MaRsVFT+EzAE22bWayQjCj1n65fwKYLqlT9p0wluc03
w30ywcYjjZTeWq4k11vjz3jiFhpVAQOAcr/d1RtCKwexdoAshmBuugmZPmusQ8xMlP/zH1oHj4GW
B3+iFnsQY4PXb43FlR+FVeJloBG3mu1UH4Ai/Tnooo1FkuJHXaQx6YFhm4tktnGaAbkHNtRrHPk1
lRaDT80bhkuh4D29njOieEfBZpGiIASiMVEreCHOd8U7WvVWmvm0fY47xxLa2MhzWs2mxBdaOV9T
Qaeqi4yVSUSWqf1htQjv6qwI4fc6ITYVtTtXChv0KdbZXQuk7MZ9VJNnyR5Oht+h3Mwy9kLs+Ozm
tiL7IFpCekSkJUX7jdrC70mUl9rpyfF664PyQa6HKOtCxkJ1p6Ifbi8CXspBC01rrSb8WRZ2egDA
MakSZZ8ry4rK+e92cekqZOfkPtVOukmJkl5LYVpWSl1MpZdL67OLBwQtBTid5mPca2KGJTYV7QIR
4PWudLqkHRKttjOA0Sl7Lftdoh0NzHKQV5q+lFtKWbfQLVT7HHwIdJJ09kc9w2rRfcoGN4ctxiOE
QA6CuoB0/VLC9z2zDwVQl27sZl9ytx2ZvkdKLlyADaKaJrfHITooe0SL9y49hyXzc30pB1tJgERP
eTACmNzlCEBEBXRWrYF1gAwQBQ/FE0LMtPEAToPpLmEO3++nl9FZ58YJ3jaXEqJSU02P/C5JKnpT
n563TZfdMUmKX9lWvPSGKNseJYLb6ww9oma6yvh0tWh75CF5yGDra6Ak/rJIi+7MO1ZAqeZWsQBe
9ac7SKtpUhWypOPKstxq2H4kbsRuW/Dz7bezNljjFiRott8vQU9sPRN7/LKcNmkJHr1Pv090mfFB
4H8/lj7wIIv3tZkv/MwVsXZyfk4r44qOCxR6tIP6fa3OlkClUFneLwx1m547/j9/ntEFrBIU1a2p
GB+4CRumYcSzod2KuD9FM1BDrWWSrVbUibQXKBAcfPMh4wVBL83H5Eb9a5x8V6dUVILad3rRJ25e
RAivLGQDKLTsdQbf0ghqlfV6SR49+PDTP22BMpG6MgQm/DoFwW44QxgYYnIC4+3N+gzBy8hgrHHt
SyxeeH0xF46gICvXRRt4s+RNgrBlbY+Xl8YKnoYNgbOccJ9WuizNswEixrsl7TTisNzyslGNJpg3
eqaPe5RwpIMPTKVJ5WVWXWbUC8qHmSGVMl7z2UhZDqkBq9WjS0dc16CL2JYL0YCQ6yKmv+Ci8Qc6
V/lcZDZF9nxrJqrI88F+PO8u9evTbyBrP5hmROkt0E84WmlgxfAKzHBO0XSdOxwTjhPe0Aks8a0E
+zHsiMgWHz9fYV9Xy7q+uSARwxIXkamaLiRnkFMtYo8MFsYdAvz4lN4tr7xUIrlXlBRk+HiWPWIe
soPVtOHbm8JoEtCoZEMwtaPW9YoEO5msLSYBdOr50kZnqhJiNOXiLZz+5GPHLOaDcFdMTU962gXO
OBbtFI4raY9vwtWCzunY5jwYp/2vF22SPtUVE/iMQ73p48HOEMKE9fsj4et8mxkVVlooMY0L83qK
PkvMm2C2hsGIDhf99RZGoTTT/JdxIrcFIhdlK6njIFmqXcW5UsaF8N5NdmMaCB8m8+J2hfj5wTW8
uf3k20lKkIiKRJa7YtQHLbqK9Njx8mJ5VcxnZ5wE22u8ETmTuX5sf1ax0gGXok/pNmSKqrOsSnEX
GCWrlquYBdfCGvVnA+ZbqMZVMcp/WfjGGpdhzbn6ml2m44blWNbRfSlf+N/dX207r/OkzV4Xp/OQ
fN0KNWu36s7hgib7X7Q+r8NtPuFtP3hkmFhzfbJ491Pz97H08USLtAwgSV72a5j6/2m23gXo1dg7
uKrcz3moAa3xh2XwBm05yyvVfNCBp89N0zDh0ga6RvIaQGKMelV24ePWVwUWTwYnKTA8xPs4CQ30
icdJVdYqQbzzfC72AIoRkBXT7Md4a4WY0VSl6E508O+rWUrHqZYesYleGg6McJu2e0zkIQD4CGNr
p1SetdqWh2USyRA2ieAixpKI4luj+uBKQk3oZKcTaogLbgDVOuTeiJaT0Op0NKwXSOkaBxusU9Kl
sDioMuXO00fgrhyV9PZrUSKD3o30cP12tUcwTuJ4ksCPoM2VAFMK12dmagJbgy3yEDWl5eZaMUJm
GxR8/6lxxXLywcQNe3i5B3kp6xYXHYe5nG8lkhBFU8FOjvQ1O/Gq/N7LsEH37hvCaMvomgDBFwZd
v6Pzls2tSruBrAfQkq+1kNp4TL7lGuLT2CVirFZJQO0SxJmfHCidQ6CQN8eVtp1rVrxuXR3Af9Vx
8QCT3UFdsEuIT6in1Ox3T8cvTzNl8bwY4Yk9LRqli9u7irGxgCha8Nnq9qN6EpnfQzMGAcuwrkKJ
apwNK59ADDjvFOdU/t6FCnsabwqvJZihSyeFU+WAFsbcMDS/RvgaQU86JIsrB/cC54UbsaBE+R3f
95NlAB+UAqZpEnrc3nWHvJtTXhUgLhcZghybFkqUXJFm4ENdIJtNpRNEM1YNSXF+Z/4lO5G+7guB
uRAIaBe5r+L0yqXUtxkrM3c5Ev3uLVgdpm7uuh12aVDpWdizijE09nxKoKt9cSKpUx8Vsr3ukp6+
CGBN/np02OX4DQaBWi3OfPtval/QyFKXjGPtJT1UvMnT/4MqPhn3yMHyCuGWTNFcr4D3XYfTpw0Z
G5HgCu/KaUkifXs6Dd5eeG1PX+HMXTgGy+K+9noQJo69F/m5ETOheCAso8trIjqlUPnhsL3IJRNB
5NZyefc0ARC3f8xwrYtICJfRdjxHTnaYyWwzPMIesbFjMGomKhDyiU+N31MIAwGmk1Ne0Dw3ZRTq
G6s64r4ttQGyF/MsvhL8HDHRg40LkrTNPU1TB3HdbkIG/TFUQA+bUVF6V1EBKb76lBdVPMGJJaif
tEImWwa46Vf7AiQdJyP55o0IcE40pj4gBDlb73AMoaoB4Cwgmk48FjXmpcBPKv8FWaqz3b1f9joQ
C7JMVhg9+fPodiEeub0kwbsWv0OyCT7mlVCcKmnWSFc9ADNN7Usufjgao1A9No6AaS9VM+oFaaom
vYIxVFMLESMYUlCCvuK/6wkTChEyBBjgDNfpe4/o9QkiFKvnxdHeJYCzjwzj5k7vQBm2vzLm0UIB
F70VQTYQ8Apkv43yMsPNA6mPald4SohVq7lvdbgMmzJvM3P8WcrUzYJADUfTPHegZ2TRCCrWz0d5
kihD7nYHnBt5zEkfSxAWEE7edzEx4aMbiOsjHWq/2LpDMm4TPRQSTM7GNZ1ReZj8Q5QY4jxrHfJb
xE5aYbFzc77DO30NmYJ75Ip6F4HI7ZopjMjZuwP9Y1aILMFFSP+TF2lrIgRN/agFtBXIYF0f9IVi
XdQ+fung3YWRschfoQDYzoRgD6AEealW8PsBkiZHFoiyJFxT7AVeDI6qZMROCHZ31GL3mrMk1d6a
dnG9nE/X5ueN1urcC4MUruDmeQKfSmGiF09q9g90WERPXH7imPhnQgpSQs3VFjfm/oX7bFhhzTiB
9yobEibP+/YH90A362rjaIhFfsWd0z5pkkOv8wiEiXyPoWrFjORDw7ehhPvyV6QVq9jHaqvUzsx7
B4+JNrLtCAIstLs52OMR3zXsbZtkpduAzTpz7gRd1owz2+j4lO0xk5VIaNmDD6uAOvt/JtwON1XS
svrUtGt1WQ7fd2BXnmmZw73EFbXB378XracMcEAMUWGdyS/Ki1wq38AFCjT5H3yiBzg1t9ejeIFR
y5uvgRrfIjCW7xTXjKTaSKC9EeHfMy71LBmZWyXTdJr4aKjX2o03lTIMmnbBFgQ4CIAv4rWpjeYw
RXC3PYisTdiEMUyXyr/zLx0thFPSPnR8LLRYUz1cDpH1TZ6LsajAcTXPFXJxacgxqpv4ZxZfpyG4
pmV6i0IA6ar1Zo4npX/vJc8uAu6BwIQ2+HkLI4ekDVGyKHAfMAku6dYR30cr1MNXh9kivCTxAHsb
5qBo9ksl4I6NRensIJevoHLaoTVY9Z8ymXPSSVdlkA9bLIk/lsOPvxQU2p9TSDhwQQHtgsw4wGqw
3WAKNytkk0FSsKckIUynfx8Cr+22QB7q2Tit9KrqmB2sH6C2vZE8SP3kTPYSJunkwGFAwJ4ya0Cc
mpkj/LA+VPfcbp4ej4HfHYlKHC39puAyc/VfnWV7vSVrbRNyR30bMr6CbK31n7HKkKqYydEAtBwa
fiqXk3dBlLqzSPRIDDoNdulcK2cwsfqWycFVQ7gHDpHE9UUBMjDMsMc89+WU9UlKICIMvr46WCc1
RZDT9ZoJZe6HGUkTBMWoD8YGmLKslEUuerku3pcp1+zfNRLZCrbAoi5rCd5XlKX9sl+CpXJr7Vze
9mdrX0sOCII/F0Hv/kNOZo0l2GNSCsU89Aw/mixjRe+I2EglmkKmG9aG/cSa1W1b0/G0pZ9B9A04
IASjDK0oOzVd9izbjn0VUkn3dLIoafV5mJ9ZSd75VEqDzUl6GwEo/+QAnM2QRAl+mlBsSbJ/7QE8
ztFTnltY69CtgiYiPPk7bz0JPNYhQ2kvNDCkrt+EKdkR8RTzc2iG1W7JZq4mmI2EMGFuhINUQkeh
ZymoGO3OQtB9QfjJNz4mZt/5aKJOIjHqWqbKrMsU/2lXWjqo2/9r5xKl7+F7OihGan9Vh/4uuCH3
yvV/WU2ITnB5/9ySTL7wPGM5Gu6cBVOQKBj5vNMzDDO1RC3bTeNjFdWjH+hvskzFvjoWpjVelgIw
BoHmnW+C85l7aFWjdxGraHYPBY2z7cWAdDzpCVSazWBcQHe6y3E7FfoVkrZTgB/x6+ThkL3oEJkS
6SjnRRyeSgi0FogkxZ51+6NhjkGjt/4nkjfOPE1gWTll00dIqLCS/C+qWZeSVeqs5C/ZGQdDmtmb
pAOQgonrGXvDLsxFVS2Q9dl/yz/hAWN258aYa2rVUXXjVd9P+jjD48iyslVDKJ8dNQE/SUAioKpF
LJMLW799cBdf61o5E7nk3CJnjYvAVPx2BAoepilxllyuySDIMAqOCURxTzGogig8Qt26pXblZZ/E
mD5jNCTbX5HL0c+sJMKpk8dHmNIdlSeqfJFuIBvH4yh4xxrCkNj8DDERqBIm+zuaUtQDXxHA0ROv
l2ZaZpFXy96hoCEHUknSHgytpb11cEsG6sVIonMDMXtDwH5QGTd8g/bGyXOxiSf2Bj6i9V1iI9mD
vwWe9UG0CBwhWsCx9ka6SYQwb2d0+uGUyVsJ4xZBdqsJE2Omgn7W4RLo2CYe+KVpR5FLRQV0yyrz
U0ydRR1ft/+JU7zE/BMDBW3va2ZHrjhdmXh1R+Us6L5AvZsbUAPvgM2HAEcEuUOdM/of0zWWm3+8
koqTfAl1o5xAFfR6btkSAFPMnokhOUkZJj/vTIGdKUzLeOGPdHQa2sE032bJ541dRtEVJK82uiFA
LcCXHwB+DSWpjoG0UVidzCgaQJoz8Y5V2j44KXyaD+OtnmA+1lZgDunES0Wtlf8q/K5c7K95MV9O
3aIuYU+Lu9knu6vzfYSqiYXHVh1Zj2vmPdbKHttMUL+7355E6Bm1OiEIqZVcFr/wQsVqStEAc2pd
cL1nREGdtZdVxL8Me+/qiXglplrSqsCeGLHW2zsHp2/eLaYpCoRL0fQDLirvpC+wVfW2kQpuCb1T
I3cho88VAaafwVTrFX1TyTNcbWH10sYj7LKgSkHtUrEe1uuWlxHXvezrMfujNtbGHS7wgM2pOvr7
bnPQJPJD18SHOZ0hmywlg/r3zwVj92QUFcRRUr+3fRVfVG+VA8KJfuIHW7bYSG/FMmb69gdNJKmJ
wXza6D7JuAvM6o2vAeLMEmHVwjGVt/gSQEeJ6sAdwgLNYjy/t/8nhRr6HsbQhOD9tkbBQZKlrv8N
95Sem10a3zyGUlW/KDf4nthg+Jy8nUxh59/aKQrAQ7MTK56D5r2lrinNlzyPCqukZG6W7QG98OaZ
cYlT4ZxPDNfXy/YqQOvWc3ddvq80B2sp39z2og78wC/wrIk44ntK+OGrQX4Jou8UV6a0zCavO9yY
W66amImNPe0C6UiL7AI1A8tACgUie/dSsZ8RZ0y5yNMaVP0LtE76llLL9BEbwZqiNLkJ2rWJNz1W
2P0lTJr6PWGgvGYANPSA53LX1AamzHAG6z0fY3YzT9ffvv15qewtFmWsgVrG41LkDf+mUKFyeDeC
+hvXjrYJyTMHiSYzLt9ZWCzZZ9QR/c9J81DeFgQjkrtE0YRGpuDR5t+t0ygfz6OiU19Rpe9Yg+K2
dwB1M15TfZPauf8XNNtNqOw/eVKK/NtNr2g6++MHDysZTjBolmV9uA2nRlL5kMPyfsTfOWRphypu
TdurlvpJ24W5EqiqJXfPgQKWQOY4CVunmkMziOMf8Bwx0iWA8hMZ4TIXLrMZoHXGJXZ5v1hXwwsO
awukDeWl7MV0SZ3j8OTxBvuFfLqE6SaGx92YQqyxdUJBQWGheQNC1ktCX+IVMWY8ckwmM48QLtKD
7ovfg0uXRJx+f6xU4BEWrmBjq4FYc06r8Z/zY29JlvYkcOV2n2Fz0hrtKFGuUTV7/RFwvrtdGmEJ
/G0qHnyiHIdXTSWt8Yogdla9Oy2mCZ6SjNa8yAQbvqGDZJFjRH1Rckzpb32XhULWtPSJgW5Tmj3V
w5FGtxU6HWK+Dr0k16otM5l4OC/+BZnGUhkr5AXexxaM+DWcok1kVtTtyO6Q0BI2VwG8OTss7Xnp
O4a069SsfS+35s6f9HZ7Vr3nvVPulLRozcpLP/Vms1MxblcHPqooKEVlKKoi30vpExQf0EOSHbsM
wN/T0n1G5+HSbbM+DZTjl5NPGSQjoG/6YPuyIJkI0HMc0RftXC1mVYxUCEqnQp2Ifbh6vW06SWKq
ien44LGyOrwUKG5A7NRrDBgKo5UQoebf6J0mNxNTqdwf/Mw91si3nCw9TMKWmti8QbgJG5FsJOh+
FeFeldZu3sq/bLMs/rDrPZDm9IyfM9a3LqF84KkrTH7cko0U4DcCyuvbtQlfZg69IF8YcV0jeO2x
HAb1vrwmuaUEbLCR/JqJ272f1dgSyuQ8pKhQquLXAQS22cTaUsXzqQs6qPA7PUyenr0+DqHa3GL6
NcDZC1rTe0bZPn+zVCe1/rzmGwRo91pauXN6ECr8MO80dz75QF10PDwtfBUzOQevffnTjo0I5rXG
JarhlpLnc6CPTIAfzQqRaLo52Q3N+6g+x2ZRIvz1kY5reBoTeU9lG0DIHJYc3ewuez9mq1MGjjZH
sh9h0z+NMvCSzGRkfl80ZEg63dIrbV4dkrSOlDA8rFBEVmHRnS5ySPnchIepBea5100HCH6s3Gzr
CY6d5HsCqutvWQvzAHuebrnHLnMdOKWHtjqgVi5tgeuhrV5xiXstOG6X4McCYEf/aGJixT+/RyQw
G6vCDaf7LESr+BK2fqiATlM1F4o4y545lkeZUPMbu+jrGaGoUheogyG3pHci7tguJfCOCO5BHjP/
HTQxE861r1xXlSPmDYEGnXb5zZRATx2nrSRGrpmg6Am4N5xW5g701Ad3bCmUV/F7i+UaUKXv/D80
Jatm7EP2eDCkxd30F12QsgBNFKX/8NgiqjGWIbkLKQT3lXziSbHuKOLsO2sNNaAp1V4rMe2nSPc3
BG3AOreCEOrvz5OtPn1cxd42Td5MsnuHer5dJ9TeK82gg7KEgOGCY6Jma3fX0y0U52R4u3viyTfQ
jhUGVrMh2ngz0SRBfbDV9s0USezjEXbFzcHrnyfMx2zgU3jUCYNCe1ZFjEb+8dOe1Abm8qHrOEoQ
Ay42rXY57lL/sqmicgLF4f+AGYfYRinwfy5cu0IL49MijnxSwWNdWWpNxx5wC2jdmjgjgpkfvMwP
KjhBaFNU8Y0buYLkpsxG3mPrmaXLW3UDSz5jn+JYpMwEn8niq1TuTLjyRUmxM2k4Jc8N0XAIkO+Z
fqwy+4vqqX89gbaX/FRlZ4r6kZfxWyPhHngQA+Dd3nPLx3tpEPjrEmXEIx2KvAatOtmaySArZYuu
wQ6SyfG+PKG6YWVcVCz64Y6U37lVRVOgzX0jbuXxo6lkV8oO7E0BYvVgZR01gyni6lBykIpVGrmx
VqSYeQlWIxipsYbISdZuvg8FVskLlMbqx9dhaYG3JCPOBj70GEOC0h0X2js1+CQZb4DirlwzmoRa
C/T66yJLN2Iw2KY1YRYPPoXpQDr9otcnqYl7C1NDVthWuLd0iZurtS1BOyaJHgGOmqdl7f3NprJG
kvCtjSZXXL6fs7H1CIDIqU1WSsxlH9inZGz3BPRjsypsF7yoh00IiJzuOH1Xj4FKTXINgKWM94JX
KkyP5KS491I0owFYSXZukbN770kUeeVSRvDwmW0YR5m7NbEtLV8/u1JgPMK4Ee2arKRVfzXiAbv9
woiXm5yd1dalJT2ULYxvB0LksYUkTD1RmHfvOPEK0hrq0ZsjFyDukN5tAbraZC91SNIHj2mHP5hm
HJ/GczBTPet/ewYb0m1C4lPjhnsmoTkH2rd/4/u7OBA/3Bs/V83DA5G40qGnwBN2Iy99vYdtUjw+
4T8v5Vcwkg/RA7zlLau9Z2EmqDxlH0XESQxBfWgCgrTM8HUSX0qvYYdbEQFq86vmW9i73mgxpfz/
f80cPg0flJHONq4Xnai+ZN8pqavVu8FlQvDlHKlPGIY4B7BoEqiIgSoDTB0xtTGwDEjTTBjThpbp
au61laWg5Lwj9malwydIQ6EZBuzqwojz6uS4G1MkYFT5tG6RnUSeSZU4VBOUcG5nuTMijPHjo/Jq
KlGlkVbL7UpvUqnPqDWP2MooQLgYvd4roTcIgaNkCN52KqLoCvqYGApAo2EeXUr6I9p8VUKnLXj2
i478Gd3NhD53CRKJfNAFKOmGziYEOUwDbxJEOVBQ3LWE8goGtdlUjKJZnFIGLlJX41Vw9kUG1cli
uP1uGaPVEPnVo5wj0E5BTJQT8XnTnpg4EXRL2k3L1embce8fT20l8mWsrZ+Y/GPgczBhpBU3GlUy
wlsPCArDHqhvgS2g5+kOOZ7GKCPoZg0em1r85JikSanHjrtScmtR9qF9wW4GZRcyTU/VOrMEEppS
5zrA6cpsI3vcVpeVDbg+oJqiDUJ4iuNtq9LG2OTFXL1ZvRDnGP61Z20oh2Tl9CFuDJEH9X9ZU48k
CoXasFxi1wtHI1qxSs6Lfu3n8zAMQL8Bqym44MUWLN+pCZu9DXcFAWTLF6qiQNRT+cJIjIiD1ccX
TqiUWYI64427yT4yN/QD8yK6axINA5Md02wk873o+JYKPFOyWd0lJCO/X9qRqt29qNxMaszytijv
ByKRNwEzDuWwlTLGSkuLpQcQUm7HKfUTGzuwtn4y8k1k/xfDtB6VGHkFvslnzakHvSeddoGvgWf4
kRiXDlLsDv8+1j0v33pxeHoNcFBj4wQX82xgVO+ltFNNEm5Lsf8FFDkAUwSIXG0XXdZoDRWm6Chg
Dt31+KqAC06Hg8A4PZiYHqz3zF7Flbll5GCvHBKXkZSQHVLrPYxuFoNkHUE3mL7eoNOs8Hm6tuD4
HcrUVUoaY3b3TsM1qMDz+52M1s7QXxR7hBhqISrTRRhqr3SjogtSYDE3cLP1O/p5kWVAWoVG0iDq
+LVfhaDUOC6L6emYTQneZEf4pPHb5lj7HJvzDPtv1YI4JU63jS5x54GsalKZWjHurfq4hTSn+FFY
hALb3DDWCaApkIRwjtn49IUFaCMmypWwgC/v82lXshqVeMbEcZdcE/0R+yZaBCQtYFoEz3Gsdona
9jeKId/dFuvx5xzTjnit1ozd5fludaTaXvd5FqoHAi1whIC3fykKckqMjFIH8bibbOMrRJffMuHQ
By1TvDyG42XXyUCX+dw/t37w4fCcFjO0weMmr39GgGhDCPfmq+F1+Et6Su3stGhDABuLb0LDaDvE
kGaLJsoeoctlo8SqO9wKcAiDTaLRxn9MgWgrU2j+hrgQhcX9oUpcsFHJH4V9b6zlHRqmTGESSXJ3
iGzBC0cCLEoZ+ihaY+LWrknBctpdm/I5cFppV1jc7nzNXy8AWQ/DvE5nRIItmc2VAankhOtc56Vc
QXfje73pT038GZI6BJbfWBTFo3FJVsTZ9dIXEZphviNUT8XP5a/9IP4Uxu+gCnnbiNvVvH0DUezx
T00GRxshJA4GOF9fjtXRUkKdWiTJ4eL7VXIT1wM7OzS4JuROgod6wBgcHq6Ysq0l6mW8UGavPxMi
aNbCwBETpvL0FE6CF3KvT53D/79NjEw2N8v4iPGjd3NekipokSanxEbcJ4kFMyrd0+07W+gHhwdR
C0GNnyXpWtkv9a5pwLsygP2E+wG1vV8HiixRPta4e98w/UNkzQUuIT+sGt8oHAXCO6RPJk2x1fkx
lbJfruS8joGevVpZuxDESO2DFYCTC9YzhMF9u6psaeDn79Nz1R3BtdkVfPxitCsHEHSAV4zbbqO1
IhEXsvo41ha7nxKQ3qVgNXZ/YTkGUm8LwATIbfazypk7z68dD+5ZE3gU4ctk+mdx97apf39Fy0KK
VBNV69pi7hFcC17dQFbH9OC3M1cKcLJ4X0KKcpPw5TSE4JY4L+KX56QfIivqYwLrGeuR3yc5+Q1q
p4OpFD7QL4P2Xurlr+FNR6DstwAYVOXZTizib9KqxG7cO12x6mVAwD9jvjF6OZaoIFl1hNlMDdS7
qMmqJZtBgT825szzMKZS8EhxL6GZ+c/S0fCPjFF6noltQ2a/ETz4Y3Ih5dvZEiqj75FES/oYZgRf
fWH/fKnY8DfD2sVTiyTQGRVldciqbW0oLDqACApslD+heXJfCer20SNOcHGfyti2lTBnb8R+IzVp
YHCGHB+0amml0Kbowxu/x9qXmc956RwCswyYjtkgfSMfF2U6DMlHAO9qSWrVz6N2hhba5qeKthP9
orowYnO9/lnxFhgVt3qsNBxvE8gCDMUzGr6Y1+J6yI5Xjy7jQ6fPkLq6IeWmo3byMMWlnCFJDHBC
OaOVo+EccgbA6UHgEUuMN9o1YoaI5ZJ3snzA0Arkd+5Lneh+9zzQCmasHWszTGleRYd9o7XxI4lQ
kmfRWk0ZYtNMWMZLgyUOqkkly/EsCkZa8Nq6cz7mWS9Jo36gbk54E7k+Jj/3JlucaqQTWrKum1+a
isiZLMc/XLIzmxiPl0ygi7o/b6lbo5GUtmerzhofCjPjyMToOy1D86xKXf6W+mdidnozAuNXAJOk
kmeHx/JAJX6wY0uyN3E4ehjR08c9jkrpdgqgthqyLXRykXBUfUBinHWcMsdp0711XnY4oTAoYYry
O8mGgFIC63NRMRgdBiQ609P5IhgMEWrwje6aYrhkljwRWdn5cdaffooj3PBgFQ4EbCc9TJ802DFm
uZvGCDHobGXx7TLBeMP2efMqo1jwZv3yZk6ITwxtFpYd/KUfQzou2owXAa+dniD4fq0urKff92KH
3nVPdji+X+5U7MShZhRv8VPuY7Pj0INN+jv/XQb2jReIzuxhqCIeXdB+si5Pp0w7xUl17Jqf+bXw
AMu4xxIjK89UyKsigblihoJhtquTZ82W4698+gkRICcmqPwCKgQefcQXhdEqWir3T79ON1oRTIMF
51YPxD0aG94tCZTLucJ+fHehovKTriVQ+vZbp/jNwpS5jqENAozzPyzd1rAaPtuQ2c+hl6KkiZQe
+nZ1zG5gvJtS55AXlCxgIgSB6QHfktEqPV4Bdr6FUmewlVo94efyN9VyyCX0W3fPjmH8xmDQXoR9
rkYKtFBU4RBkLDRZBF5qL61CujfYPSNFQDp5OsA59mQyLMhKpxH6k/IhzEm6yqJebsGSJmDa5JZp
6snKd/11XGkm1AbNtWr5cdLz20G+thXlIcyaO9at5367YhvXa+0NQEFp+P+ZR8mBpvkzQataf9tJ
SZKWo8hDg/qtpcILu0LkqRWyVnzfrvMy7Yfp56/0SAspBE4l5/GGQ5lZ4JUUe3msFNF0IgcUuk+B
XURkUdIXaw6nihQlncl+0PAYTUQsPAcwz0DCM+iIFpsu1gmaydOyUdxRyzxQeEJB1QmsaYM79DE0
0RjiQeCCgNL/sykiXuCV/l3O9XZncQNGPUG41ljbwZt0IBZSO39kmv9XQMvYkpIojGgW1LZUjMov
DBnYchwzvvM0jYJ/buz1xWHkbO0aQRyKKRTejABYL6h27BpO0QR9Ma9cZ7qCkbZOmYaDajNJoRBv
F7NDVx/xASXmLhKbfh5PLwucFIxgi2J5FFpe5rCzWJqXncZe2Fz6kwuDvawjD5WhUKp1/hMaJLYm
R2zCov8RE3Q3jfc9JNvZiPD6ufolz08vvf53BRm8vOZU2/aK6+1QJyvI8Ys4PW4DGv5sF/DPPER+
V63ASvGspiG+YL5e2MuTCMchnz6BqqbtzrJgou4N0yzhpLrWnbFFXTsSprPEwKQfcMaNqpIxC5NU
U7/LUsXeQ+ETNYIOm3FkgpBCAuaUBsJebm45uX36BAgS2qM1/+88KPRQD5NTCS/d5DSXe+IIIt4H
pxlyhcCW5Zjjfsf2pQuIEfYJDBSar6xg3UFug0C2rmUCWDe3hy+GmVjYVn3n4QL7LqXs3zOLwqJl
hXMwxqUtvejKwjL7tKwx+okfDydYf2/I+wXN93dh31/7x4DDQNjH5vv4fjG+j5PgoewCOYop7vGt
o8hC66gK+jtMQE3Od9Z/+GOikOU81wS5tpo1kxJBiAeuNOoo7nxZj8CYmOLqP+SgdtHVPme0uP4e
GQWzgHookqFDiMzXAnpVXEgh91DU/QvE50+cBh4G6uigcYmPdWFV2gpuOfjqFkyxGqA3MdybM5N+
W/z97LbK0dMwrlYtqwt699OAhTVBVBrFLmai9CW3BSLZShC0bfOMbb4lFlcSfiIGxjiI+MXg5+8k
w023uvsja9Q2bET/KHDEap9WluU4ql4xV9FLQyKVwym50MqVlnndzFR7tbXGG6yilIOiPU+4wVKg
rtr7xTmVDu8ihJDCZyP1RhwrBSYzaRkgOpl33OF7X6EAJDSwBRicjbuaKeQaqwWCG8b1IL6FTly8
g6mb4iukZe33bGZ1QmyQ5sejvgfghFgjndrzm4jz5ehuFK2WneR6w82aQBwgd1h5kK87HXKAFrq+
ZYx3FYuZ1Vzx5VUchLQa7CJs2NqkWLmUDNWcfQxCqbBbIiRSnG8ScVPhBAtWaYsJ6k+XZjT2iyq4
iuQfwD08jfh3rFUICvYwrYrYXskZtoodX4XKT20bJLC9DhB5lwBczt6ypXymrsSdTt1jDX+Zxgdp
uCeGa4VN0b1+3Eg38ztilLla4P0Gtl8xYPT5AOXlniFxJIcp9WAvJjq2By0znzAUCjxJ5E+rfq1U
lsZEHViMUJ9lwTaDN5xUeb7vh0d9WrjTU4c539Kz6M0N+DcxG80D95wa25zYMTbPzcBXPEPrNDil
jlNCwjoQe9LZGqGlcExF/tdI87ZRGsy3Vgco9I8nx2F2o97MjxG7CVVhPTSmot6E/IZ9sGYjTL7e
9uc/D/IWN9VJAM+HABBcX/I4CftwDVVYOzatWDwviqqQHCbQJkpsa2RTUYOldgrP5cKmJ/l+4pZL
vWaEg6Ta5RfaIXV2e6z5ZQZdkVd8NlRMbhAIK7qxB0hP9ZJdE/5+wxPAUMAh1jKnBRPG4tCTGHx+
8+uW8DXMDj0vMLvJitk4DqCsY7qehnx+HyNq74W0kpUAxfQ9wOhK43jBtEqRjAMEjp5G/aq0LdgH
j2GSnzvqWbrC09yxOAiUzfzlnHmDL8NdtAwDllGj29wO69mObYQsc11UF2noHXqJB5Uv0FlsEmWq
yVmIjUBTrk4BzOY0tpIePoRuYnOCe9IYZLvQnyMQXIf5IizxE6rxOWctUly3c8XDHpfHC5XO1HJp
p3VpnvU4H+BKSABNXr9b1XZy1Rt55n6TPzUo7pdwxlZ/yk01ZhvUZr/xggdbSHSs4lzdKVdbxvZh
Xtm3zWeyyICHnrDHIQ9EOfvU89mazTYyACfLeryG8EbP2pkSwpeKUtdRDmdYBrbenwKsKi7mZrHN
nVwY4zxwUdo1Uua5ox7N2AGQHr9FJwrO3hC7M5oLJ+QPcp26v1PvbhBylMMmLFBDvLPIzY66hApB
YKI+b4wvD52075bR+RTNZ4EPWc8+rLPEO3inDLLKBeHNUk5x3NNBloa+m20Oh7+kFpAYwe7YJrSl
6QEVuZl4G1D4uz+ao5O7P4yF8AgprGHvUG/EtwRrU/nHiZq9agpQd8Tn7mHBHTWq4rhpRd67GPS3
jOY5PoOrS0+oKydQtKLV8NiPen9Y9l75ViUUoBF4XKj/XixU1fnzhC8lba/b/Dg3cNKahYgeY4vO
ARHZWOcRWh2sggi/eExk+nGv8FdSX/Keq3nQAHXPSG3SknoTfvc8hDYnBPdUwB+MIEjipiWaGISW
EKT8tnz6jlDRAvw7eGEkoWxVeJ11aPh3cCk1HviLjaju/1SeJR9253bpxEqN/GeYIk+aYKAey29Q
b0W4swhBrMsT8BmTz9ILfla3z92ZxH5fJ9XdlLuAgxZKmtivTJxwL+K0K98XQv2X1pvlaLnk9jyU
xW0WMY2t2eUcUEUiBt9t4s6YdXtx/F8wctV5kHsEhC0pQMzZgUb+o4VVfeyyqBGQFX6rFNt80plX
XlJtg9DZ81D9Qo7oi2hvghRDH74wjgixN+JBmGnR7mbZY9PtmrzIkIxqF4CZxTKo/+EqdxergRMU
zYlr4jSYFQxufLVneYbXmsIdWt830M1qLpvPCiuakSGMwIjyb/AsQAXlBo9ouRkdJfMzP/OY6u9Y
SQNXIBe3furJ6F0cSfpGiQvHengxDnFILsvnUxl0tS1iD3SI62PHcSQcLAHXVpxSLOD//cFBoplH
gqET9b08l27EKeTERVkR1rjWtubUnO/0FzkKyimaL6T4jSKTvEi7HQDmrjHVWODtoUvPkbWd7+V5
37XPBH7uKAXgerpNbiBIyAkZlrjpVJU6WR7P3elQmgEX3i7CowkbIQFZJ/TX3/tGP9BsNMVL8bMS
l2imDPAUKpSggp0jufrItj02wEl8x/yfQV8D49eEx+h10C0Af0AquEPv/3+qpfPSHOJaE3wjpz3m
hrVSOTmnl2bTInyYDVY8veFB////UPx/3WVW3yc5Xob93fZFrShDf0p33I4ZHxCIXDH+/Mq28FUP
hSI2K8F5OkPE+vJ+5L4NWQ5+G6gH/RBx3DNdLcMPHmzlsPiYbaQ5OmyzIRw4L33FSFcDZ7nTxsg2
mKciEBSVqYNrqeijgQe/l2vPdwpGWE2PZwc3aTMy1RnLOh+McA2wvfrQ3keYoPovBqEgnOHc8EUg
m8r3/HAbVYLyRkhZTwDJjhqHaCFomwaerM3q2qmDXxaYOMLldrgHJZzIwdoguyw4D3NSNVjmqFfD
thWthc0J5UhfuAUF27pdrO+3/eL0oMq9WfjEzu4amki+k+4cq8B+Rslv2qiPbpI+AfFcU62l4GM0
8+nthxk8oHGZsx0VpqengEcO9KsoxMsZwwUr9aQGSdFZzHPcaANfAMtSL4ZUCtTJEqP8ufuHmt+h
K68Rg0HcqRs2mbSk+enNKPata43sTAEg313OJtD41XWTn9FE9B7ziImHo5wztkQyoVg0kFlOi4qU
rzI5LqBD3Mt5ylEDJWW/TtavWhZF6Sy9Gt2tNZPSoht12H7b0crLS0ZVDbP1N4qfQugEdNGQ2PGV
lo1Rb1wneV+9ZqcJr9tuVZDTjwVadZhPMd7gcnD53RiVzKbrxe1J0vhR79YfeLoZ+xHRdWiivZwK
i1UhpzEl0CypbL6licHaPI/GaZ6PY+4FJdjHD6DndhHMG8zMWb/IiqtvHMPBZ7hTEtAURFzSrqQz
6PMuXi/yHLPr+kEMAWqInY6+nlH/0xlvfh07tUQde5XeslzM5kn1Uhl4oPbpVMRrzHqDyLVdbncY
56bPdnLM+fIgfy0o8MXFILIwKIuceNFCATJcd4dQj+yIf6isnZ2PPR/694BvJunzfEkgU5XY5wrQ
fO0AVjFWOwkzVkWKLfTqYNg1C2Cbr8ySwbjqlODhWGGYlSBHWH52CUW3L34Yzyc7g6g/vfd6IoVJ
a+nN5Mkw+Qtqgy6zYgtgiEyY3XYy3GxsU9eLYpoyP003a9nQLWb8JjBtV5fqSKpgAVdfrp02podW
3ya+Hbmrk6NGaqTtzQQRjMCuTa0hpry/iem5wEts3bkU5d5QqRTHxWQOhV1G33h5cwlbvycseWWO
cgLPgr8R9DE2ouY0N2rTuFvVYXqeb81k6cqy5B6sTW2LWyyYsWnnfuCEK7NHCJtm2OAr0KgEOuzf
/P5FyPI6CGS+wLon8F3A+6u984JQaBcVjSxx4/csxlsyUI0nUnCtEQgySeAxAUjfnhNepMVcyQlh
EXmIhju4mo1S1kmhStKYlsgp18qxrgkgnBDdAeD5iXxd/Mncs8IMouekX8e6tDWYOfDDKakS/O4Z
VASACdkK6SbyIkitZRBXdx0ZXPR+nfYZsq4QY59HeSGpDc5ZcUTF/VZfTbpgRDWklIfpVVSdYgh/
54LyHJcQCSd37gkhrru74EXgBa105O3GK42eT9hdAOLr0kp47JUxSUQfZG9r4o/AhX9RwloR5DUX
HW1Mehq5pm6+msCCe3sADWxr+KkK/c6pxNQdE1uEjkgAUBmAAYMz8u1DyvjF+UWowvHCr7nfDL5F
LaQ3em7ZdFge6MR4tKk5pDoJAWM4ljHSXXMx0YZRDbox+37O1hjGvn6SgsnvwNkbhv9Gb/C3T8U0
wDvPq81tzomsNzgmKeDYalb8nuQdkUK+CUXZ1TXYd/Q2zOELoycTUxaLc72bMccEBfNy7mv+zFKJ
Hw1kGjWK0givwQIRog9msOCf2CByEEaX3LfXQ4UZTU6gP0FR/rPuMczeHKkjQNi53tvGE4gdnK7D
zP5pQ7bD22Xb7tQ84LuxqgFQsWzsIbSedM38Oaxnva71wMEcRKo7pILPIT8N1cELmv4b2NupiCSi
Soh8Dxwvg8AUGdObpJ1gNrnt0ZxXTcjl2GfQaVFMHDNcsAalieeXxOJDcJrQN8L4CcoQQSJy4DfU
tRdaH7dYutkTvr6Ws81Mxaq7ju3vEJ3EyGvfiOzmb5cchYg0sfJF7OPhaY12hekdFu9zsEi1KMZ6
XmngssHKElzOiWrpNGP/VMhaI3pFP2BAtfxL+M5krgB+Lwt4BZ+DzTpXVOe8SG2t7jgis6WLkm6e
bxLT4bTG2guqLicoUuCfYcWMQy+guOp3qSGgm2A6Bs9ztGPfOdCvTsrVzRBoRGT7jJNWUgnufjrM
1BSLDCHDa+GAvRJOkKnCGrO/Z78zfEy3z2Epi5tYe+koonIbMLv0RNb5N0L48ZA7Zol2ZxW0efxz
cMKY81aWg8AQilIfjhC5jxmLl4qMGdRfvli+Ib2PWn3VX5GzLKy5Q7ryq3LqV5C7KBXlp/+qiH++
PmSaeP/Ul4k6iYxEnCJA8LKGvdfm8VbXOka9POT1qTG+Qp9Hn7xAeJfScfDSJx+MbVsfAzdtbSRK
Xg0059j1Icsm44/HEQlZ8Pf4Rl6bShX6/6eQLZuGd9K+VTg95Ne5VCsjUSZ0gee1AvMXdzo9QZfu
78GkQDlwOatheJDQd2GbZKyF8qLt5WBShL9UqAKKc6S/2YNwSfB0S6vMI3EeBX5hfIbzwbO/OkqB
OVs60kiwUKOgU/rJ0u2ui5XzrXmBO6cygLHnoNaL/Aqt5PR56rw0Th3JXNUKGBAGBV299++W7sA/
gzlcMzvKvepoHtpGznZUwAZdpqeYZwWlLwaxSpyPVtjwWZFsr9ButPtabz0HyK7Tf0sdbXpRkn60
KnFIT7E6mzIiKTxMk5hgpcXON/vD8An4Pm6dFEkM2783YRgyEGekmGGd3wakgdK58DK+XqYBD2w6
O6zB/7a+fXooY/cG7YlLUIu34d2jL1l8S39v0UNk7cbmJr1azedKewFqwU2a669vg2ceVohuBi/m
krZvQpnmNGrrI7GXGqfhAOyqRTwsPz09xNrsrWR1kri9sr+o278SnN3JovsxIzdpK+Nb9ZsMgHIX
7hVAKnyWpLSuyRaoTr3FtqZCr8xco3EheouKrfMRsWZf6+aUUKVU5Z+YBg1CT0V6ecFK2G4e9ow2
98SFaRJFEwdeyCd8iqlbeCdoIqjMRKTWyxMjB8MeIHiurgLHIztH0KIYE7+0ImkEFoB8eAgnZtSQ
mc7n1wPevBM/BJk0ldT3BMRbMuhgExhTvi3jXCWynwiibTkwANtgxSo3SnwozLkQjAQo6IuHzR4F
KO2tPLZDa0Ix/u8wvFaqXgMqN9e7kc/cgR3ClGkJqQO7LSlbMO+ywkeYZRCfGEMkUy1Fjne4cIlr
OgCWiB60mEnAxN1NI8lolSVe2XzeTIJ3PG3qtXiXKAYoipaT4FQBRyhXXQaCAHkQrpYxcD0+jbdt
M3cBKUrme2O5H8A8sMhAN/9slke5n24yeUVvVBLKD++ciehpupGLp0NWSJ+ZJUBgEyjE94RcQK4w
fHhhfLpQot+oBXv+v+ygqGv1lhjrs5cGR5S77gn9sz4Z/WdbfCTYrXEQgBhhI/AB0G8Tdq3hdkST
9nc9COK8Th40FfnRgek2AIVbYJdkUyaQwDN4xKvbAWCqb5/k+lpnRB4EPGrn37fyVDFW1eRU2UBO
b8dzgJLKozUss3pB8ciU0AttG1gQSIEthiAujy2LBNXwfLgc8x0oBqYC+ayixKlJ/whqaqmbK2Va
bo4N/+yi90xZyJrkHQ3dWZPm4t5c9284YnEB8X8i/rZV2nCPa9jWAclGvtYt9/WUmbSXZeRod7hn
GJ+JGuC0a9Jao0SaoXwZaxlvQ1Lq+RNYm29Pn3TsruCTUDQF3Pg7ebTfRf4myETwLRuy5xY9G2YX
SBZEcvsubjhF/M5RKzQg2W81tNMj+qqOZTLBu2N25Cj8s783zBg5nogR87eLhiWdyn8TAAkk9mi9
FK69O0U68PjubmzA+UdWr7TXr0Yc4B12rUpw/AhvUwj0YhxFeuhFHhB4u4Q5O1jr0entonaG/sih
iP+K+lBeNqdVdh4xkkjyPhBN1wM4oqPmX1tsShhE0Iy5KZdbDPiGVJV0vxJVU40NaGKsJ9VX4xZs
LpBxo+iwNrdwtXgL2x7M5eo26XW3Mtx/vtkjX+wFTWb+C15vfhL5ly5r8dFga0Fxx+nXkG8FVXm8
MyeOroA1Pai6F9zLwyopuK8k+vsOxqfAuH9RBSXBY1vPkF+vlvOw5r/pLwzQgGW+v/9Z//kTjHl+
23JfHZHfuMiw9vpV9YIP0qGx3QiUU1xm6AwoOPpC/jFl3F914IL5tLcEByx09udwbsssYCwy45R8
yifRg8xffPim5g7mw5T4NJWeVAXDO+gePr8F6aJfOfZrQzWNNi3S2DV16+Y7PAo68u1vrJzgNBhg
B9OLNY8URU1AM61DmKD1dP16VhW0yxRDdJ3GHoZhQUZvwNUKyDm67CQOyzReO34s7QLqxRpTKgQm
IDTYacSExL3MC1zaKMWRz6gvj9+6EJAiyZhGbsCwIXkIowiSLkk1grcM0nUT2Akybgq6YopMpiI+
vVxytYAyIqdlfm4raED+06nsgyNSvjodjD0tGTJtK48fJRmjcEm8KlYkl2x2uASEbdY0LSIp7C4r
jvWHm7C+DlCoXDZKT9rf4jTV+dTkzyyrtlS9QImQUOQhw9U+I6I89qsts1n8qP68Od7Ld/oJLtVx
7aYj6GFSgXOpYY4WMv4VHzNO3Av9qDkLbEgev5CrJ0H792vX0k/y1xcW6obgT9WWU6sFVlxVIhMM
kMG1khLAovEay0EyhMm4D7aK+hfByz7ZG+79iR1lnAEKTMGyiuK3dNb4Ve80qxMDNFGKbf+b1Ct2
GWO+eWmZj/fwq7CRCeg2c7VwCz77mBBjIj2/r6HfBTtJfwb1G2Mx709fC3DNeXrhvf1OyRaaGhgf
CxxSSQVwzp1pTaueY4Ritr+MU/lcPeVe+RjPvpvs/5tGucRwn3TBSoO7rWJxBGRF1l3o0gnleZ/I
9r3NmyTDkUkPNN7v6vAIFQ1Vqcn0A9rj2Spt/K59md7O7OGE8eCzG98qyoPGTJXlqr2KjmNTIQ6m
ZA1Xt83zQGeZXWOkE7EdGrQ8CiuG+RduPeD9gnXNV8h4brnIwVwfe3KSRQCU0l5Io1x1UCqbhHUK
MAIWBYg2lLSb2U24gzVV9Dihu7rbMNnBL0tlA1Sql0+d0e87skiYVIt6WLBjbk/rreOjCT6HrYtK
r8gYne9/gexHhEOewPUpzyd08Ew2cZ6bNwYEQQRkI/kCSiPI78Kg6WmEx8yal7koZ3bC73WES9ee
/2lcG0tcDhWk8IlP4FilPKa0c23tZOVTEx0aTNjzHSDrdm2wBBOGYYZC05NUMtxFNjQF6bNNCCn1
6chehDjBCfwgsbHipPcD915BKS3fWMkcWs42r6d10oZ0l18YxDXNaOpdc+KZvZ6WVY3mqZez2Tzf
BROfZtcSQGC8wt7gG6xwOkRN3GxMDU+OkmhawPaDwRfrm4GhzFWKGvvnG22hVliUhvQZyhaZtBfi
D4sdvkwg17EGy4o7mzqpzSaHMtUASfSmfYOglsYyJNcqh8fHnQuoIPRm7O5Ub3MLx+zysliCVA7n
SZbPGsKw1CrXzCeKWTAxeOhdj7JDZebA4/Ea1NM4VYeBS0iictYub7ZjIGeDfRmAWhhvgBU0UoBr
gxCvDBOOIsdCIazrwr2hIK7SgifsP7ovE9NYCIf0esiMzf4+yvrTjPrwbd60JSC7sHcYYZKQ8WQG
fTfzqqm+Y8z8FATEruuR5b7ym2qrqwyqOkPoHTdVDRQQST5JVja3Vyl+Qcs9cafLCBjPCQCLHfY2
A8loBHeKvJCJH56rG0mxng+3FQYhvvDRkZW9NmHhwqryGBvUNxp/+NGzpiPuN3OSR69G80VtQLFq
sZRQHrP7j9wsfLA2VdZ5qnvN3wbNGCn+wYSz8J7WXx0UiI7rWmcjn+wJD7YUx0z6cN/zE8Vo/ZrC
qrl/SBzuQu4f7xXegDWFTsIOzke68QxLPvUhM8ixJDGYK2nLJjGLI5Fg+jQlSMUnJYmF55ANgBn6
HpAE26iKNSyRebpqs7SNNPEfZyHafNymU5HIqWhcXeJu+/4aJGBGgwa4VILy1jXn8Obu3fDifTL2
OhsFCjidZXXm0FOvbuSIbBvzLXuGCxl8245DpEjYCH4GXcX/8pa/WK/G4oGnH1hcjfOxd6mpHf+w
z8wFMX6mu4P6wpO+JwTAomF+fKiCkjDPDJD2D8fBYVc9koE75p+3MESVx4oQeq6kUymWgSWq6LxS
AjvUS309IvKWVDijlVMHbydOUh+sH9GXT2BgyPIR8dS1YqoY9l2lOe+7Ldi6LiwwKIMCbLhzKlyU
vhT77h428tjHhR6vQDB0daNq8lUAF7yfqbxzosiup2B4sAIM+6rciVvoYG+HKc7X/BL62EhOLqQa
zKsB2JmhU3Yb2ySyEJeo9DaLmJ24DR2zDQkX+H5JGnL7pPdvRJz9RK3R+xT0d16FiC7HGXheswON
E0b+tCZ/iUrtLXiBVeGxinXyc4HCugweO1aqqrpuf9vE6ueh4KfhlcaRIuWw+RCAXzQAcx75mGsI
yJ8HqMre63XAjk5JoQ50wDn38T8FpBGlTSR9kmQbxNVH9esrmkMxSbBI3UgEaRGq3duRAB6diIhD
KwvrhAPVzPmm9vyPt87fPMilnw/2l5VwnFKF5VpVsxTARG2oNpGqVYark+K924B7YpvHcWtZAuzp
96oLPawgghuxQFuB5I9EhgbTnDNhL/WFk1U/Ubw5GrjwMSFnhPyPg7ZEnCwgl87Q1anTcBCulmvB
oZWiDT+gSmCPicxtHVuQ7sTZqEDiU7TcXNAFe2DHr5nfBJ2rN1cscLlHEM7AeM4Jkssvrm5CfKNw
deW878iu8+uTmlOvucH62F42Y852rZuomh19yy9LKG1kCRza6UDDnmC5sDs12Qfvr2aj/zozGtEi
VUYCkP9+Zq18I+VqhgOOHBjznLOxfCR274MB776WTdmuIi9ud8hwaFfU1hzCQO3uEUy7yPLmzFpU
NJlcmJWhPnddU97F+GHjqxTi20mhsrcgCebtB3Aq6JicXtXXQnupElnCqS+tYwyZmH/lUe7IrV0z
QCzyztf6j5VR+xNCsvKH/eGYX71H1tPphgoKe+yE4HBF5ZlkYzlhb0D2g31tl55RgpFhacIHGmTg
afkBZFXg+7RPTRI3ehARvW5ZCBU8FP5hj/wOrVesR5Vm4xbAz9Cj8vD81HDFZuFtWvSieEXvyLD5
tvt6JQAWSxy09xG4PJvvg6P8v8zADUDGxoA17KW5nVrtP/rdhD5rsKmWWDS+G+WjkPr8rsYhPoHz
cO3fHptVKErIlSeSRU3e+RBgL7nIMdgo9NcCjTh+OOc3YuFiN/wGjhCKtGBaOrNK398OHKd0faix
32MFmNm+mEhR2Hk7t9clYAfOKtE/g871zBmU1LiFntxa88/ICRd8l+qLekMhLS85GIsUOO+6zwJ8
l0mbWyQpBZvkL+ezhNeKD2aOsJrf6ZSmd+sVLpebxHtaL1iS5PyMdBsv0ZLgRLrXH1vPK+tuoTMn
J0Fo5HE/oTe+mKleKtqVVkl0UIw4L0ZWKTFrYJz53MYL1CTavBlaePVV7vK0TEUoWqqutZwPgTXQ
YNUiS+5O9JaxANtpp4oOICZajuR1faXLVbwmrsLrHyfo4ER+P/eft92YO1AJdAYqPzkci8MsMdXW
eUe+ByjLzzNHg7aOlmcRG2L7liFSR1Oyc+PErbKUW4fr4/QiLZ9dIXniD8oCGDiTYYVcz6LSMkdE
RJJp8qroZBmCQR+sztlETy5rP/RBCGaMUoGmvuBjjhSwuUZdIlXsa9KhVoPL0UoUpjecquIa6z0O
nBT76y20HZ0FA2DivVNpfmWbW76cae8W6ZKCt5E3EOZUCfia+s2zAWmJgMq53Asm1BTKn9iZ+V+b
KJX1JIU/SwuhTvqCentrLa6BM8leIVIiqsA/GUdZsxojEbquZ2CW9McCH0E2qfVG6U1wdW+gbTdy
99zdkVNrtz38mjPNVKc91kmLlnVFpLvfqRXtI2H5a5YlCDJa53ub+kaUDrOjCAvwy/UKzOY539Wj
/3gjV45kt/mSP6Vt6aMa29TzNhxSINc4XIfwl+Mw+k4/L74Ukn5kwmP6ieMEnbxE98V5oywLZpiX
e1EDA3Svy6gJ+7mZozHlZoCsQGPKnSxEohC8I/xfVCjOyQMk6Hx/LIfi9CZmobA9APsYIGBEu+30
1LUdhfTI5SY2OAFsQ0Ck+X6MYT27Y/1j7FemnMf2EVTC2dUPu3h+yYNJ0sCfU/QmVW/R3NeORvXp
Wz1mRtLWfqJCCCVMQHfE8xc9tz18hTvNJuln72b6KFh4TwKQQgJdM+dDIL/D5pj5vdvOZthfGc3X
eC+tYmer3sc2RDLTcEQnALFthPnwAvOvrjsf8EIdwjWbqr72oFwdVNxEJhDGw0xx2z4qjYs+yKvz
1qFJP/YGA8gFV6nKGjR7L+Dtbd71lFiq3QgfufWE0Yjvy0U+hDpuGCiwWBP68y3IMqyEkwwIsvaO
3WnzCbNag17j5iuZ8VAPMy3HKqlRAyxlU6o0i2sKEW2UNdFAKzcCVKnUhSopB5aSofe0ipNihAQ6
MVbdSLmy5ZkUlryxOpOFyIK5UUKo36UmfKsDtemo/L7ssm1hCWIS06I8S9PHpOnJy6To90saSNL3
pYrmBIVpuBy0dl+JP2AW5sEBiqZkdgLwLgAtrCI1exzxP+rvVW3O9t0NjPx1/h4mAg1pcHqB/hBe
9siQpc7QjSJ8r2nboSo2K9Eb43PLKeBupN06hXTAGmk1aVgpMws4pdi4B5rPe5O3gZCxX+XTjFI9
aS+KmOr6vvXNQtGBw4B2DHJd+um+306z32lP037YShY7U3q/ExAz+Cjegb+gmStwnL5VGS+AtaDJ
Vm8fPdfpiLg0IUbor/twpn5RFRjH+VhW34Tc4c2YdzvzoDblMW0D1CezWLPwH9T+DmG0/ls3U1YU
lr+vu3LkXLaELTQsRT+XMAvq83icL0AKxS2ZfDPmpYtkjuu1qbxJdeub/89JRQU9Nc30HW4p3arY
zXaL4q3z33PbMzNQQ8/h5pRWzm0KU10BIZnVqRgnTX5HEJYE9ZCxelONpQmgj6ahYGzoE3obgUW3
hIhXXHOPJmyBqHT9Llrk4gNaovq3ST8EzEGRSwBbZJqUdQkGrytK+YKjA2H67yAM3/r1nWea9j8E
kkypZUZ9W2Sg9BVVtwp9qFWwdpeIcuGhZ5OAoZ1OlJDx//bSJfppCTBcvxU1GLXIHMgdqQBy6FdR
lJXTJc90l7QcgZ4yUEpnSCItRoRt9YtLZ5uy4sK+fDlhtjLufAz6YTdF8wG8medfTr20UcTli8Px
+4WLcCy66RvaOB3XubrszX3qeMSUAv1Ff74W+BwwFerizD/tRmm1Cbvav8DBch/MzIZ0isRdKYYD
FE2vSuVofNMZ1TCy/FXcXyh7uAD4x0XoOYE1TAtiLIr6Rc6ushzsSBsy9FfavAY0gJDtYzsW5Df+
/Iv7mTLDYcVoHk9Oz+rq0csBW2BLThQXCsbE0zx4PcU6E+d/n/oKUpW7dqbFyn8/BwKHwPlGEqup
kAexqBF7eqehUhCAm9SSkaJ7Eo4fOYU3tnVIK6xPwxsrlzyRXNewHutDiFCdRg55zlnMnZglusce
czaLx3y29dos9WNkds43qF3dTSSmgM8fZVL8btVIQqWbnPi5t9z13qoCd7LMeEABOJYTSxzZUiKZ
RAJVLv/Cae0FwXgoD2efRfioxfrAn11h7UL4tAIiLeEfZ7aPY6bxjxiCX1UxAzlsgZBnplcO+0rW
aPWczICNLHKzHpXj4y+owlAPlkpKX70nGu2B9zuzAwz30JbkgVaP5Vmc/QLv3eArn89TJcymBCF8
QAXF4QR57yAeE4kmO+PsXrybv2aAbevol8ZpgcsjzzyVd7KaMiCdWVKou0ugo6F2YxhKoObzCCh9
Zmg9GvK2bI7m3IzRQXDXs47mPfrPTFJGOgjBGnHNvgeKrXWVWlKNyEwZwMUsk1rgY0RYlTa7/FU3
IvOtY4KJCl8+AcwKBjYklVRgE8XkTfwQ21HcbCUn2QH8lhDHkFnMDkzSyC8V6CNhrIJX+pboCdN9
1kkxmai0DrrTp/7ipDl23UefiBYvFnmchmi7tOHysj+c6UO37xPJeQdUoISSDTj2Qb442Nxz5B9D
+xaqXuh5zaIhTwa5T0XVxB8ZZjd97b49ELB0Lgd+tH9yFaY24Ez4GgXeILZ2H9h3y+SedxjUQe/U
jkwR+Ow6bDR1iBxahSR9Azb0vebPsaaOuf1jhaXPgHFKMcmkROgPHYhmPbrszVtodn6Q26kHUOh8
GQWvzJEZshdhcmUoM5jkNENt9hb9M7+n0nx7x6OvToigXKgEGkn3LNK7a3IRyElZ/ezP2u+4Lh2o
3hRDg4LozWL5RHElGfcsPHyiK3HQMmLJjNyr39zNwd9E2xoOWz68J7cWLb4auexcfXjlcPajOGlK
iv4SK8U1Xx+zc9Beq+wgn1wOFdXw9BoE3yQZxuXCd3M3TGU+ilap3h9yL23zpUmecX7aN6vq72oZ
gzhUhD18+3ra4qEZ9wPNcJYQfvyfwBVLwv/sy0aoP8bKceB/U6YTUqCletWn2KM0sSelbg/8QZZT
iN8tek0injQMVWtnBnLb0ozvgEzEqPT7rZO/YImDacOUAAjJMRU/KqELktLrq3PhgNBFAbV4+LbE
LL3lHVKdbJIFqhhZ9VcVlNDFRXZfYuMCMlWJteWMZ4nk5+rBsWuqg2rb9tN8pwEtKEnE9SglJjui
1jqDshmCeG5BdGFsmdJf+C1AyljD7tGSM+99Ked3GiXfPoJvx0d4nAk8Pcr+EMO8HYxkq2Ru6czB
W46yy2+bjUvDaJbtNKC80xrZLayRc/e/TXM+r84KWz1Og4ffHVsQU5H8sg5a0R4b5TnoeqZY7m5j
5XInhmLvTQN+r3n/GAGPv3FUL7h6tEnES6SldkB1fxKifVb3KkeGXihXA7a11ckCUEpeRmszl4kf
hCcPU7Q6F4otXmuFDpp9Lzkub6yeUzIByIPJEKcKRU8OSabBYSTWucNvLvb5WgPBYvg/bVfIiw0F
TmMNAKXSF9EAMeIR8GQ/dLFRavEwf3HVH1LdNZu6MO88ynoTPG3TSKZdFHRDSAGsLwEn6AkBrdPp
l868sQvRcid5mp7U2T7iQrcdFs+K2AZthZWAkhO+gOkkuBm/VgOOddct5bQs7o0j/p+12RWlMHYY
Sk3/u5VNJ8ID/s8F0GTNwj+p7M8ww1zlsub0czHe8Hpw44Q3KbpiGucLgVyGddETrRykBrT9bs51
7z6dBAT7u/Re8JzLkRRYmMV8n18aI4756bb5abl8epiRFaqaFqz5fgZ/rY5NGVI++bdwDryfVjEJ
2hvy6xhKI6kGPiempPPiI8DL7IbaYo+F89z25gu1gACPyhEmUVwgm0ebjBVfGffo7dJ7syC1tY21
/0e69gAakPMaiI0HRMId+hKWv0b3xPNGh6yUY/LY95/POT1vQksoQOTGVhKRJ14PJ/qE/9Z8frrZ
0jc6N208Cax5xPb4Lmo3pbJ52K9ACROLzdvwG8YR0409sVZFo2dJPP+lAmXLzjITfZWxxW90hQ9F
PS3kMyIiUo5X0xa1NKQ3C5BckxMwKxHvwLovcJ8IImLnNOjzB3Ad6qM43S4NNrg7rlMoPslj1LVe
dgt8/oRPwDstj8JvrR64kTFn9195KZAsflrDHQMmAK5PCEA/vjz4sjwQrQBpQUjKf8vbLflNaYBk
64d7QxyMZnF/qvkXQ1pwxJKS7JWGdIyNh5zD8Jg85PVzB33BigLOXLmuLmfwnS8kgpdCKtH0nEli
e1Vk+DE6Mg6bO282DZdNByupZRj2dFwHCOqhJUzoc72BrpQoBTRbr4o6PqDOJyG8yZahOX1WY+XC
n0lkxyNHJ2a4j3xZKxBQ5WAUumfd+8P9GTCDrQW7UKr1HhcY9V1rnLaWo4lNWXPc9gFXcA88UtuA
3YtZb8M+mDD7cE8Na+YK4kesf16cJULQR5kclMNmAQuxlZIHYUcIJMqNAdSgAiDMYXkf706QPvi/
nXfsMbeINlXUUmCsbn5kN/hPAhBmkw/tLOgwocJc6HX2JfSEimrzjtOJER3KIbbpcf0M3RCFBhxS
t2H97cqWO4fkqph22pGt+XXVMsWSsE7FW5crsJdDRPmUGVzjh/jj1Glw012k4X+HliRfW4JC4NFf
Tgxdbu51+DmcnbHeO3TWGCSDDSLWByLWcuJqjscvt5S6TLo58hVz7IqVzVfjTzjbBEF8PddDSa+M
slZqoelzHnNXT+QrCTxUnUAUOVAGwWt7gbnwAan4FDqOvNabjOtLFwXL2EP6KerubNxNBWAfIAqa
m8oRUov2Rarujh89CEVkaMF2P3x1vFRY/duXYv5JvRYrcBywSmX+HIBP5beae/Uh1fdFEKZxI4IL
ZCzIzToM+M+hMpZ4KE6V2o+djHtkglczUNZuk1WdFGHVAk+58MQ/useG8G5JTVHPKVJK+Imji/49
4fPvrjsCH/nTxeyT1kB4AIb1dyWDoIyuodhyQoMv/6hw/yiPDXXHERSMxefz4/T7deKFtK1tPLcE
eM1SFnJ3JUTfheOJofR1vxAzlBTDf/Rsma0vHsJfys4ZysAtSfBhh2IojJ6TpJ861sWHLJVawZX0
iTm9Kp+0E81j8nsV7PdfWrkwQGTf5oIxYuYjxUdUoZflfWnlexncQylh3FFfU9S/76pZA+VEHWrZ
FQOTOzgTbj0eKZwHFiHpXYM94l3iOuQGoZ9PolklDsz067V/e8ke3nNZXSWoctDpcThXQQSl0p+k
GtSKJzYOnnZPmfJ6yQRxguIxfnmefoT7ZnQhHOStvhK8bpZ3aPnQvuH2x46FC7HrHpRix0xhC9qY
xAkVhYZf8RRrdZEutTvngRJcsHdbJESP7cg4nKe/0eG1KomL6BgZV3YqXdOwrIbqNi53o4cEIE2N
5NAnyedViKeIZIzDywSiOlftHhd/n55MhxajT2BX8BPPxtlZ01BkxbzAC+5tCfxLrd6wUnKaKPCS
6PFlzQdttfxPi848Am6oQ4A5IvPGCS8M2Ghk5pJ+nPUQ5/Z+a1+b0HbkuDyA+l0qmME70DcvI6aY
iF7aSu+Z1MU/+zohXlyWTmiBCpoGU8sLagJTqVJFAoNc/QDxXio/eDSUJ9ZXLMA/G4/yATvSB7Xh
xh+RdaqH+F1GaGoLQaahuyCZeTg7GpICy4xhDIQNsSYfUKIhVkPeAzXaB7kHdbA/+XVvdAJrKXap
Qr/xMvcKA9ykGqgHSaYzGkCYw+Yrt0amB3ITVY3E1SbwdN+/kRKIeNJ04E3NP4iEosvaXUo3dj0d
Buovk8ZwD0YcnGlEZBT0EHsNMw3TGOb/KzfEmPnRq7FmZEkCdxdPVzKsXy0KUk6xAO+U59cRP3g0
8Nj31LGG2ofcX/WUox0tBV2olfCY0rVESOHt6Xq0Jgs9FY1NbBWsoXphEEOejo3kAgz88K1LVqhK
UyPeFO1TbIN0szsQ7DTIbNtKuxdO3qbb6/50Ub6c2LP87H0nYP0GlXsg1ylfgGGp85P/biCiTarb
iwFcFs5mG2ocjnZnLjXC2+6Ro15/HUGFs0keYijey/ryCSn39x6uAg4mmCp5JsCI1XIvYN66uiMQ
3E7m/mUzMFK8VTdcyqkaYyARWuuko1n8qUK5+H+if2grjw+qwkcIa/QorO8ZvrXxh1iAz+ouRAi2
zhmFcvHf+SJD/WWRU9yCt248tY+6FKbu/u9q783+PglnIwknCjZ8egmmxpS+go+U0i09rOi/5HVl
zN2fQlJT6c9Nu85wmzlMxYoyTygRpz+E0MFPZ0FctOAwQrmbYSVdMK2zySpXVHKOdR7IlN+nvR2q
75TsSkCALADrLW/X2vHSqSQv8YzmqSP5Lokkq0Iel9skK4Eqy5LH4SNxLL7YsuOT+KIKyiK7R4ye
zf4r/pYJLLF96PN5kEK5Ycr6XpmoEKG2HRbtWg9dM7mOI4+m9lx8raIL9z/LkBwqHeKDCp4kr1Ce
TCCO9L4loqixH5bNsmsIw3DLr29OLJVzHkH+Usb8PLjTNM/CqeeI6w82yqwddXOthgRcXvuGGhn4
2uDYJfCE+OqQrA8Gbg3gOnoHMJRNEs8GQBvV9MVxcbdOWUHBQiRwmQnM4MjRfmTfFPuF2fRjtrGZ
KHtdz72lsJwKOBCybzBa14Aj2Xm1I9y0ZAhicTLrH9Ry3QOLx4owZ8JzxtD1DrUObr/gxdaMQc8N
AY1vnPAcsJT2RJBDdKUW36uEpnEbdZJjtq77vbnDI1d4r5lfOAzoLyznnMDsTQO47G5lBiuvvkun
Eeew2Qe+yA89CLFy7eCHlaO/yrOCHBxKcr99ZfnPgG1Xs7RbHxYGsdJ72M2xHRbBlBltYI9voIn6
Buoqs0BYdbqDAiKdu+kALx8tIIfJvX6B6sSXg50fYPGQrkPgXnlO7LoT+C0oQi07Th142ktdRnsQ
pShwFffTjZSqN6cFtvqXE8WHuIb/m8rCsOSpQK8Iqul6/5s1QjKNNROzF9hoOSiiAtJsO1BMRmVt
v9so0gnSLpxDAvz3QJIuZD+YWMSLD3KcvkiBw88GEpdre4OmQPceHLdQr8lMqcB9DPra649ptFds
eUwM5oDgrNY3n0/QxgSkgyOGd07O42wxDJfPISJUaSg9YWx6vT/I5PpIKizJnAurSPBy91fBKoDr
ETvJZ7Lc8l/xnD4aOxeqDmYg2FTQm210uQrkNZN7diUkCudQcOQH/+ZvFmrFkEUkqd0i8Z3YgRzT
PIqcCSqxPHgd5DhK7ltJMmG4uhc0RRrc7RnvkVEePM4xP3z32Y+GDgUkLoK77joMzePNdfqGHWeb
5CVM8l0fjaO38u4Cdax3JGCI6SjIynEtgdFMvbdWAe+kypqJCGh07n/Dnh/tcjH250yHqt5hEKO7
3rY6x9jE7b6X5QGVLhKz50t3teqixsOg07fcCTBh4Ni8nspbtt4QGoiid8iNFY1IQj4aSOLnVhbm
e0lX4vo+0k8oGUfBq1OIJOXflJ7QsM5nevDbnurnIqzxcOl47KmgGHYaqSvEVWtTFZTA6N+5GkHp
wfLWF4Y7dVMTHIHlPJMQEa4nkAXbltqRsD5K80+YQQ4kzcMg7et1myvhdciBNVTcE7zLN3O5Qecd
nlelokKUDxMsOB8bA9lKyDUcL36in3WpJXTHU9o4ulJyveYBKv4fnAqL+/b7+hmDWBwewancoxJg
XUHxeUzgxtcGMnJlYwJxomF6ZPgEKQuE9dUAm9oCMUoYNT3JFF3AabNn5AQvhE83Kl6z78g+MRqg
d4UTvj0EcHPotjflQYwdm5EzNCjsIy9SqnPiDnyQ7GYpODPP1qrgisJhftsFCzx9LXNDFTDEe3xP
kRiwTg4Gcll/j5mfZJqNRrQemfkesxmLU0DITLB09stvnKbuF8fSrIv1ibrh9y9JWJMXHt8ovSYk
95q4glISqFEPDZclZBpgJ3rzzM+tBdNUTt2X27PIhOGi92nZoUKa7YNzxFJ0FDOgNRCr1xdHmNO2
QwLv3mxQhhxpJwFOC8VDtoyzhPY/wAVqoFTgqaoYmOeZOPBih9twgf+aRJxwdhkynAeLU7xwVYAw
kUiyvRWtLtIyXTPrrVnIaC/oTbYg6p8CeveHQQcAfwTOR65gk7ACiwULmEbASf8ZC44514wJxTrS
rR/8saXq5WdEXRqhSac7Qk/BIoU+amQ0NIG343vivfZfKfHdKgMJZlc7p7Q6K8T5SIqrgUn+bgR7
HdmI1eKHX2DsaznvazKp9As1Xua6u5G/id6SVXIq7c7IhAY4H85zee41lcXqbw1CMtE4whh7MA6M
H2UoogSAV1EiXvSnq/2g3dqpwgwVo+JnA2Bni/VSrir9E+WNMIOPcr38yEv1BprwCZA+JwyRXKfY
wYA2a3UviP724UUzMLebSDY9tob0hYt/DsEIiRuIMx/dyJ+fmLhS/lZa78jdSlEoOoBZbgqLt5Nq
eDHxngIytKMs9PdvsqXiiYEn/i1qZnGpuj4hOVP7HJ4zk63AoYMNBmKChTzntfKI0p4ODvsnIKdx
xL/dncysYMBj+0BK7maZ1g6AOK1SLlovJqKaGH+VK8pSicSHB4/rzGsZyH+ssyycWspxuftDbmmC
/jYVZwsMAslvvTX0YKzcPgIfGm1M8doCwxXYs67bTuUhmm5KtLqtN2NoAoh4+c4LTxjxXqNAqBGB
M32AkNYPVdkNmN8xlXlQ+YQtE7orNn1jjdo86WqZFOPHrqzs2Eh7bUqgQdH1AckNJKhJdCbWLAkq
grvpHTHxQBbl8m8LhIPfzpMftwwzE5aDSaS6mAGznsucNKEtmlWGYkn/dacKzaw71kdABPP8QFck
9TnViii+I59O8tO6MRDKJyB6VPLYVRjdEtB8X8wepmMbhBMXL+X4fq+uPUiih1DPVKCsixs4NRSH
r1XHPCMqDeXUkFt//AH9y0tLLrg9kS53wnbIQlLUGVl4wdwVZe76qCDhHSwhzWSWMYmPD3IyLSUW
JTtHtXeA4RToWX7HWwF772I+BOG4SvFv0K0Ax0V4W05cPfrG+UMYHmkc89m8JrtuJfuXXFM5HQin
oQLf4NobNmldUinvef6dbUzVeSvLMmfPJnumjUHmwNVsWKTfHobrRCe0w6gqtRhs06wIZHpS1gTn
bDfR/RqK8LaDTT4u6TfFfu/TcFRQUioF6U+npw34Qt83PiRj4sOESdLhWtOnVsH4WtRNmYtsur5e
GvrPkWxaJ+bSS3FGwfp7nxZk7TvIWhGr52b4io7fVMGqMG4xFyr2x68LDXfvqfrHALIjwWsT4dwe
iBRY2sM9psdG6+26CppvZHnEO58mZZf6D3YIpT9KelUqITH2zJiBzg9Veu+t3fTbuF6aOYnh34ad
zmJsLMFz9AUWIMPxNOYrHBducpJU0t52EfznDd5iv2r5VHKjhZkzImlEz9HYLrONvV9EuP9cvoMQ
WO46gl3/c/sl0DvXctFjW2RPoFOwKTT3GQUf+mw/255eMOxHh+yV31VCzgnkJ55iHEiUr11VSNcD
ekUt4VLgUSc7S/Ai+3VnG4Fe0tkUGsMt6G1hagnwQALQQO+6S2NBtsJNHITESKVF4tq2ImpuH5L+
mLFGnex/fF2IFobdbdemGdwIJhTlbQjyfl1PClfv26cbyO1tU1oXFXMkv8KLNDmflRf9k3JMwXgG
avk1QP+yJ1zHX2GCL79Cd85ToBnfbR0DfSvCdbzf86ZB/LgZWRH/LyphntXuZZP3tcw1c1gOWQ2i
IhGWUEI2CaD8XpSprAcMtlT6yBjd4yppAYtstPxDj+pf4U9E+xAdMRz0FrpNTB3yQckv/vfVfdQE
fsuUAoksVWC92/J9N63oa21QpsncmJGNBRrpxbdofFpMiZdmAzuqYsji2zya+Gb7sBGCjITrXttD
4pOcS3Dg22b8ahEEgdhqoEBdIBk19Ea0lwAUCcw7fvJVQIEiTQyPOc6bGLKpxwerjzFcN8GGoJZY
8FCKLRqg8RbJToe/2yhaHYLf/+5AKIc8EpWs4js2JZolReJOVaulzODVuN4J+H3FqilYz3h+j0o4
ylaimbF+d4Mpnn0vNiitfGDJWl3DNWkCt741m1jSawxzSsRAEJpk8XODpsCG5w50Yz0NDBDpSfWG
uY1fuJ+Jzx7U/1F1nlLH9Y0ShEVt7BYkwGsgl/H0HpjZ/GWNKHoHJm+LhrxLtucVix+SU9AeRkMr
EYoMQ033RDKk75pe8yRDs/dm8hrZ00R0FeRcpCvjgpsudrKtPbGM/rK3WLuhlrWV+hS4Qdk3fY9a
ofFAhaSuUf9VqU/jUvCQwT/NmKSVlrDKFvv4YrJcLbXtVzyXqB43dKnlX2gg7KusC0VX3XbQ9OMS
7VBq9fi2Aa5VTxTHsHae6pxbaqAB+NlDYnll5bkxhRPVGQgGBM3ZmSsWWd9anqk7twiuzlYwJtcT
8qZsbThtfaJjBAoqzwNDD5rCn/I5iahB0kQ2re5vjOHhbbAx1ASDjQpq5Y5YolOV0l/SLbF/ppfc
JvZ+kYiZ9LkYlIF2pw7UaxDm0Yl5+n1jji/OiScJtydNclh+lTUdyV9KHFz7aSO4BMNOTYvX44M9
ogbdqAQkMkf6PrKxxQCc2Vt7OOkyfheXraeBysaSJWe5b9ewhYe/QbyBBGkcAeT0TbD3JH4tlh5Z
70BuSl+s6jfPpz4jjovvb3YdNM5ISuTsY3ADkV5DO0RPKQfTtDyHoENJ61McqWFTZ2zkiwqNk6tk
JoEDWyr7miSlI7q0wQIaekVIIcsWltkbWUJpUnJ/QOJmzM+jStLSl/569twZgKyVto+QsgP6Rd6S
DHxWMgVOrNf5gs++8PFZnBXIU80S5Ir+8ZoMhBlte6d8MenpYc/98NFzvN6+lMeF5oOcNPJluAwJ
2qujRrGFqx6bK+gUwxe0HTzwyn87wY1UxATGOH2jWbzO2VlFLHtDFNYghOFiLuANXX4Xee6s4iVM
OrTbjJEZvS8DRvFVJYYWmtdFkMGu4lIyKJLraWFgdighvHVGub2qKuyxJrw86849+kbRPpAppYeB
Zb4KJbddLRonqiCEzhdhC75j1JTPBiDGMp6MnOXDz8EWC58lfF/rUg6nRea71ouToGitn9CbdEyx
SpqSOsuLv4QUSwVKuDx647HavINAAddiP2EmGmcBLhCq8cpYLNisA4YilFJzyM/6t70A5fJSTnMg
Hf6CRqDZ+XPZltUPrJNJHd8k+Moo46PqNZDfRw7oXD+5jhZ0n0oh8gsVp/ollrhTzUUFECF4oh16
hEMTw+voziqu6yTCGhqNYEq5lQMHs4NWQdb+ZjEY6g3/gbitjo1q0oAJNP2qkPBHOuYBE5Wnk4Rk
qnsUuYSmsyCzHGw6ZU7B8/PRY/VIpErmQqDU2GIPNsu1J/K6NjVbCxnaQwBLCytob82nMRUva6r+
+kcZr4qtpdG36nXp5IjJ0OWHdUl4mGNeaGVo8u+4PviS0mHjiWvojT5epYvpSwOrAVf+4Bf5Q0qn
7yUpwWZs094O9TtUm+pEOt9S4ublMlnTHM+VbZcRSOzUcehptaTBWly1T+iKeWO0JXV2GI6XANf/
QI9veUekNY2LZASxJaid9l64gdyUYmeacRSXRS4G3ifaaJmdRQiE200goVQxelUNMuX6tZHsOvS1
P5K+2GEp65+SH8niIkSZKi2isztdUplQqYRBUQ5I8sGMEkEN0oJ5A6JhGuQcRHV6RY65TGTYXxNu
4FAEiiaKXD6hUiM1zpzJ88Z+cyRmHIkIaOhQwxRT4bhC+ZSf0lL4x5MDlHSYmxQwbosLl2kbpfnk
OR7yYtMI4SGoCRXlwQqmwilhV71uHP9uAeA4o2/VXk28wgksPr+HJOS1ZN60nsPgwXz4VHMTDXYm
M/t+q+D2chUTbUj3/1P4JHxaUzFnup59yfqcgK0fPWrpLGF/Txq5a846SGMZSZsgD/nz0LZdsK9e
iOdZcwxnoxF3zqv1U8Z52WV5iVKggLpoQVzlcs2mH6xPdh5jiuxXggUl+oPBmAIZC6hIbWfvAo+j
CmX9YBItwr4DaJ069YZDRKNfKGLGVKqsJ1z8jMgShgeXziXCIi12et9rV4zW9MuINtuB0+0anF1K
OnWbvWA+c6JpRp3Z8OAZxqUoSEpZ5dE3fuDBsd7pn5pXFMR7LQ2ZVcsc/k3xGNs4kP5TG5B2JHcy
VLe5iMi1wkhFCocZBf6MQRI27Mbuv4pAqHz0QehAZrEnV5eATKMt6pqY/DyoWyX+x7wKHcbvJJfS
QP8Cgd+G9uywYq/CLIQZU6Np50Q1L9PMjli0n+KtQ1COTx+CtVLIo5TYDuFIaLSBa4zTYEuc5xBx
V4vaCzvZSuDCpDfghVupdozRm9AhCDFRU+pAeRYv+8P+xlEBOidCv9OZTWDlHqmlOYkRmtEm4cRt
9z9gO8su1VKhmQ60BAf/8BQS6nCOKi6b9O0poViey2IaBx6q6xWfzRfNeMEhu3BpqwP8mdykmy4e
+12QKTk/vUrHhHSAbpNsKC6EUUHixT3K/91IuUE414oJcn1HoOrgjPiufEqq6KbbSpY+6drJXMy+
4BgKxIxzYvatd5f535L+wtFwPhS8sDl32W2/3yHnCgh+j3XB3aCwFuo4bK2iDi81wx2EjXHiZtel
XBBZHJKuFvOZBjCZOO8dlXxfx5SeT07AnS9gSY6wqNI7G3TAb50cW7nWbOapmfDVc2K872rGH7j3
axV2MQo4HDoJotcGhZsacGvehzahiWZsDK2zRKVjNTzunIfEgstUtTmIUnNzO3Ods9m9/pCY8ao0
zQdLW39T8xR2DBKy+O/9emA+obrCOTs6ihEE6cFmV6kprMH62GWk2tM9+S4xCjBoajWtXCtqFSfO
EYdjiYR9GiS7TzkCOUC++BvrmhmhU2lLxRJBEF5/28jt0ezZFH/cJcAPwnC0MaGDGztSU9MEm16w
I4PQB1jP99pe56n7mnDveqkrvBK01PDvxG6UQuPmX9lZEOUWNztslFmARXHfPCvnDs4Bi8K9fiDX
L5zCLjr5zzXHiPhRzJlEZHliLQFnV0PcDJkBREI/9CCiTPYpZZev+Dss50e98DXfYJO4rTwdP/QL
3SSUjPDcCGoeDBhwfpFr/mkBmdV40gwruKjaThv0+8WXbcXN+6sB7xccHgR7J/aq/WKFIPyeAw93
RzbZ6mIa6KV8OFP857rUfkrreNu5IHZ5pUqqE0VOXMQt1Kty6g6TLPHhkfldlO1dgt0JUbl9r63W
Yxl1NIaIGg0nMZnhH26noxLMM+tVVXr1FCS42DWtwXpaWgy3XG5eLLN8vMe2k0RW7vQZwWj8gSnj
iyT93PJWlr0AggRTUb8qEGZY45haHwVU7+t9P3HZU198WMo/9h/oVjqmEs1lTi7f0TeC3srC7bhh
E3sL3Ua6YZkFinI7GsZR/5k4J98LiBF3By1FsMLmkvkNME30GRb7+Fdfuj+afVwetom7phzqsyxj
MOn7eNBS/z2omK/eHYvtQDKuxlfyAoxfCrb+wYEWWXzf8p2Nh2HrfEIdWT5xRla6/QiTTuqdTYsz
/TG33KbFlrTfTbmvYQ6LqTCCvfyUcfeRmfgq1swvpm0tNEdqSAwMTCRrIOMDvNjL+L7/FWQIDh4c
c3g8RDdy0yNTcjWTHOFlAzC1hwOXpLmLwu4pF2NRE5vpzYxfaE0kuh+A0+FCOTiWMogl9ggnigtb
TpOsfJ9yTuTpsOTk95xHVK12d7fu8flp4XtPIONwTfC6lHIlm53pBDMG2F3iwFDVjZ6JsRb5murc
H53bL6glnAtjIMmUHChT+QjtLsnU1IKxB126SDDXpLmmsZaZLYBIciOeHxIFzOTnZhFWtkvq1KRx
P0x6+cT6aog98nT/ed0GOAR3/UXxVacwXnLMoVh6vBoCqmQ7rZQND3YOsRAFom86hDqr3v7dBQUt
WGKG5+PHhdHt56/qB4poGCZq1C60OLQOBXaLZIAxZTGkVkkKx0vKfvUphkf+htvKIiOsTmvm5txy
5s7bNL4ZBZ7YWVHpGa3cjP6nch5o0ivn5SjGdbf03+XO79/VLUMpVGbncJWwY0JRc9xMrx4QE4HX
YEHUV88Isqc54smHuSj44RyIsbwGeUlBWOwMnlPobJFRLkw0Vw7js3+Pyesu0kTNbmU84wBcNRHX
E+fswHXjQ96EO5iwtIoLuBn7ddScPz/zVXFXMo9YiVfr9Wmcliq2sboEp7OR/rqbSpLIRW7+sW21
P9jMrjTUe8ANz1/zWcuxyilQpbAp9sNMQLPFvv/k1RygXCJ+etbNwgCm169CziWUYQo6S7c3LZfx
B5lMorCShkhAnG1hN5ou4IP2fDIJ2hSUZBJEoa5wvMUULvst4wxHL9OI+N/ZjCpWu2Ti/a9WaL99
Vt583aJOd2YMGLNo4CF5TNhyMjM2XUkzB9IMVHwaTaJNNA0pT3bGx520UErioA4eAkKfggodoTsr
fdLimy82YT85CYjgxpUgTHGoZY6qXoavScp1uBITdILd/xEhIFIECPa/k+WIX/XBkX/Cw7RDRsMd
RHT0G6vyW7Fv1kFphYvwTrY3ZBteRWYee+qEMF7D+avmSrQtdwciE9HFt34jOKX5RCElJPMMP4ko
85rOS5MmS3HiU3AkBqsiB2m+nBGZuhQaCSvV7gJHHyu0FqFa/cqcbPcpzZjWJfzdfLI/37Tb+BVG
CM9/Bagwu4tRF7Lq4VfYHkJ06jnjoXxZaODfTuSgrDslNMQs/bH/hctxZYb5PVESvJpHZuHIlxoL
sLZr3AeKjLih72UsYOwa9jhqji09SQpOg37fx+8qdC586zkK5Nd+ZQzMHTCCNhYqIWXxPMllT9to
f24p1VC7+DPES7M5fpGIMs+IUxb2jS6TyjBkvrR5uM7eSxAMn44RogBwhLViJJNfuoeYXE8XHp3S
ym9SwhCyfK56UrvpOWkXfUhpPdsi9W2+RUwSzMbxQtKSShJK42XS/BrA8h1zNZfDES+QX3ommeXb
BrhoKn09r07f8qsO9UyE0Th0FC47w7OH01fBeE7LcSxNNYxIXmUiHzY3OShoeYdh/QEC3CzU6x0w
qcdWXkohBHXi95xapOcdp2ER3orlVHgbZKZwc5KPUfrA+FSMp39BfnNFE6WM/Wq91aePsZxEDyAj
+jWNYT8mAn4ktgsGGkLCjz4PLJdFyn0Bwl/+l3MaQxxs37/icYs8mg0TbYDYbVuQGauIgOpJTOvL
zbYrFlSD/9s9UfrRx+ULIr+mt2LTT6M8B/lawC1K06AC9eovHzyVDd8CA5hSDMbYV4iv1bs+e2aY
W8AYSpz+V7UuqskVpMYCKv5dsj0+2Efa9PRIzJA4eGRlVMrSger0qIH7wQOiidoHZMjmpdBcGgjE
t5SqZXJqx98ji+OG02gwbJFefDHa8nJBHcG+XrOADFVr9c3SP1vcpDntzMm/11CilYLqb8405ikR
AWBcn3gmM1W1kPR1FLZwCf3VT2hIJjR3q1VGvA5tDoOoI/DRgZlzFFqx2Q0TKvWGx45aR3fTYTMZ
6BIKaN9uzrEvUhWxFG5sxRQTnrEs1JXrtnPe++hBh4R474BHqliq8dmkRGPHIu42EGlNg3ob8SBs
FJi131TFo0DGa84Fc21kkHpK20ekJ05oGMw47HI5aKzbym5nsN/wQIwn+0Lok0LdE8mF55mYJ+xJ
qIVyZDwu1s9WgOI32OlkW6PW8UsJbq3zeO/sglPTTzQwKglk5jenrMEiEF6DP5tYoqLfgRjjkJ3i
BMjzNdKD4sydBAl7dwO1ODmmYEZ+IuaaC4yuXlDYRkH2AdggafYr+9/WpEdEaIkXIvR0335x/xGF
w6nmYWwXjw1B8OXIZaYNe/gQSAgEjPF3bRxf2pk6pohWcMXureXWSBOBrFkEvhphpsuMUnXti+Nn
wRFrNZlMuYIpgYwGDfForoOYm2ZnSndJB5d43uDVTro8vQ2cY3UJpJlSzuI+18P9QEECEwRKrE3q
LDItNOxDSS8FPM+iI5ksej+opV0Aihb+9lU2KM2ysfog0HbV71efbx2mHSH/gUfAeWtMZMIFw+29
ulz/QHE2SeHeTqEl0QVU4x55qH/CjClYhcC7DxHbGWKIDV2MLDPDuaj7jgGGqPrm38401HkUl8FD
ZZqEsnYTtS6/7KO4tEmDtrf74GcbZElSIF5BK4wmv0J3kuXTTVJ3zk2Dxhasf9m9NRGeYl0frOYS
NFUuFqD2mDkGc5YOragQKJhtOrFB8/zUaJ5gMbjwOdIZqffXBSYzlFHunxRfaoAObKSHLNx0usl+
qdT2p5wrTrq29631zbWCrMXKa7EkzIxTwjylgK7UdN2SNvzc7lxVTTgsYs6QSF5NzTqWpGedbpEp
MfOVttPq7XRrc5uJNO6nZB4et/Z6M1/7f7SdDqPZ6J4GRUkrglQtH9y04+nbGFh30ClelwF4c+ER
uUBE0h2bEOjSLe79n72hUD+IQRSkj5IS4Oq38w9E3acrn+zvivH9g+QTQC0i/xWh7gpSz2hoZGeL
2Q4PHevyC6Hpu9Tgt7eSKM+WXFeLYxn3Mft71WB8+2LgVGclmX5lQ44SD9i++boSY24Rg74ZPlk1
viQCtzg0koGN3ymrbADOFc5AOP0NwAwOS1tQnyg+UZcZbVsaapq6XLMXtVpVTRoCD2uVYMNdd1mD
rmks2ENw+ghjbqnebmUxY0gSq7yaLFYg68cQ1452LOU2QhLUKtXQzIAqwut6L3SPMIsw/gDi2bjU
OZkWqTmWFH4bnaxMjznOHY2kxLy86b164+utSzuAkbTp3nyTEnlwpFBOE46ptiyGNSg/Qp3qvcvK
17qkk1T1vkJ1SFCTjrk9I3f6R3fRiEmLjeKkY4KNFy/hVcHUUXdRtXtq72bff4M+i81q3JFq8Dp5
/9sAzfbyR5jKQz9ZwSV7pIDkkhOIgHF6qITAoEnzzl9ovq/aMdAlYpcFsH4QnpgYg8FfCSJQ6a1G
/I6lWfI1Fq1v3ExHTWz758H4wdQxWj8fgnKoMOOBOEmcMXm/eSadX18y+09G1wAt6ToDsc712aaA
47JWcsF3+RiCbSne1MIl9ACbGXvXRTtM2efA6odNeFNnPc3r/+dLlByA+IXXkL269LjjrcoRJFml
kr3teMIx5AvleUKwskOB0PY2ub3UJeKs2zusSlsI8MfoTFZC5tF9P1HE283fJbl756DnbePvfqBk
gA62Clk4C2AwsFIF5lSkc4a/jSUcS2aWV5Kh/xqLR/GTL77dLuaGx07fgZv/pOE4/PuAHMs8ybdr
uxwXfXnDn8MZgThMd2LtJCP6osX+CGXRaCKCe0VIbnwJLVZtEYPvX6NC4xEsuJjssuWUUvZsUM47
85qw2/xINB+TaT4muG5lgjNzkaQAu+y7Enufb5IeA7MU1RO+kpRegJjiZDxdtzGx1nySGCNeeCwg
UjWNR8/n99k4vj4NamnxnNYwovG2K0bheKP2TKvB1hQgj50Fbaenfu92ARmKVdtqhMS1zyJboCdc
UjHcpDJXbbZxa8y6WgFl/nHd88wA8cK4O1yGcsnnbZxwfDAJylBQ54cJYt+H975wfQ3pdiH59G0W
UO4XKECVOYNp92N+nGH43oNjc/wkeQVwwbn+4EqVCpQ4ruUV7M6Nytrg2CCfz07SezKZ6ctl6Gia
pZ5yaYs6YmZikPUuHtDTh2xwlKYxUQz7YxPRPQP6CZoXy+fKR7DABjaIezKsTXDGIPLw6o5KuDRK
i+0B8d+9yJ0P+rjFuHMKOPvqWPcPaQr+LW0ZTgmNQHbMZdv/JRmqeJAnd8qfnizTiYlrmdZ4F7LV
Gy0Vp2p4oPMAamaXPqgqxW1Lp5RJsOmRplZqyvGi7kQsKQ9J0i5BRDCyIB7M5Rg2OWmRfWiJ7MB1
yb1fLhHkRkuB4YIaY3guSDP0DkutPgLlicPlrn2etuzCD8Cb3bWUWWlMTxlWe3mR7whp95beqyLz
zwCFMPOEkBEHik10OWuCJtRwf6FrpPVATzDd9FcJ5tu/AQy+r3gU1EkHyvA8KZGTET56aFH2bdl+
sVjct1usAQ1Ab5Q7yvVObJByxqA0KV3iDcsU6TPGGZwYAcp2gg+AeUoYht1+suLFOMiFa9LLZYsc
ttvH1HBY+74zgaCGISyGfTbIsHBl6KCYo/HWfu2uQcyep+znIsj60pXk135Lpd4IHuyHO2qer628
QkL+hWW1epgvI5g/dbAEmThu5puLYy4W6z7p9rGU+qph0DcQlByY6so1Yo++cHcrwAF05kQeBmHw
ZDb1rS/MCmOeF/N5H36clSGinNTwKWu+UhXzSTEmlHHrp38zb24zaDOEPC8Kgs9DoVIHWKs/niLU
xzYe9JR31QjhZrK0SfYcxtg4Wz9R8nIRp7ZTbsClVjOwBy8+VceInmCC/WW+D9aJXumPBYZbVgXH
gazyo1NMDhi8BzaHfrImm2XzYOoYcwfDIos3Q5Z5wkzuKwtvnZUtRrnnbBZUGqfXCmY9clgDVfIR
i1Mbri8PXF+vwE1WOqopRHyu1I/Yp+c7mZFF5jRWoC4HlZnQP9NLAFF62+2J9nPC4n5p7weN2yK5
KJo8Jfrb/65u/99t1qRJXQE/If8LqS/n9DX0mr57HSulc6oKp9yPjvz2ITW+D33naR0g1nU2PK8G
qkHGP3NwLmyVnK4s0yQkcDGbj4A9UDmU9/ZNPxF1fYcMODyDXDpyDaomu3pUPumRAyzqdysGsWiZ
xc/YIxnjhrMespPm3Zan4ocvwoA9ijNVikRc25l7ofYJqNI/jT4/pvIL9RhfZ1+jJGWai+c6iWcT
04rfep6w0X+N8797CuGg81OT4GpXTkfJ6qUJYo+Kdy1/RLzCFBM0BXlwCkQhnREOE4JUJO56AktD
VrOxGhqYiWQKX+diPi1XoCPCEs+NjNvkkOw4t/g0BIbqCnVPDtCn5CwcwiLDnqaFIugIMJmZn4b9
0j/qLMbfyoWZvAjBBaYMIwmnrZhb2CF6IUTfwJJC1UArOsBSZRlNPzNk8i5FxWNbplfN3pjwaC8H
K7HinAsTi2Tzf5sS6UWZNSEgAnSNMqihzhCKiJR5Ww8EWaFzEDEkYDZ4uYYWHD0M8aO/4hGEvU4g
hfWN+RTKjV2xG9haG9tybTZ16pDhZFwl9BX695Z3XCWb5MlXy1UFxLGDVFjVFHetCzX/XF2E48uH
5H7bdFYugWPPn6k97Z/p70icaGSIdt7mtzoT7hWZMhiwosfHutaqGNhJhHGPUEcdbNgpBCL9XCsA
6xFzr4iPOBhHgmP5GmgZ2YZ0lEO8BSovK83LiPtusu4aqHHOKLFW1wCOHBDPFAlB/JLFcBQ/Q5z4
qcF+8yfYQKAdwCgpr1gsr7im2YRbLrO+ueGlZyHQFERp0QvTSKYtPZ8Yz5O6v0M3ZwjkIlplzoc0
6FEBDrhn8Qp+FngF34HyVGahFKx0QHdeWc+YfgGysyJGVbWffG/BBZLPHHIv0m1x34BtQologRMd
w5kjKWlPZQZuq8BkWPExzcWCfMlqkV21UZhCMVGak/zuOfgtPcOYxVOEmcvmq2tYQaUi3FeFPHLD
3bnya87aj9ukpN9R3j6SfyUkkv7Zr7LiDtTdJy3HL0DjdDfu8shlV77Z7yfLQx6VFs6jhf5nWoa/
OOn6tvhV4BQqHDCM2LLkr/rQ9IuWL9H5snb9lIrfS/PEoPR2xWCqSjbcgDMnO4D9JaJR54Tv7o5e
7KyTm7WCWCPwOQqQGKYkDbKk7GN3urFU3QhkgvUWmVHp6LigZu+9K/6pvV4xWO+wYssLnAvwN7ie
5L4gf/Fb3XQYhgqWdM+oF7dmD7H8huZPt6cu6fwA59L9Rk27D0XUgmrqed0d1XREEYLRu6U9YoM8
ug9tswWT5dSYoXczhwmO07PK6s4lR5Z1rxOxSJiP3F3M0GRLUOKbPwyoz+CaGpgWmvFq1TBH1rd3
O/PBjdElPNBAqE7zgJdMB/um7U9zajU7B6u0kAMOlyjedAl7K59vZLyVWNMP+FBGxNGfB0ZNVzYU
IXb4o8xf31mZSQY121UunBJtJXIRUy55gzq/2K2QeHfvlB2ru32UCQRZO8ON5W3RX36UxHrmh8jX
W2hU1tjZVq49Dhad1vyuerY4LcNzuLH3nQTX/c1O7jGqera1MhbdG0AHHbH3uf4bgM1TYoWpGfGn
xoAYBHo5dLQt1k134tLy/j9hlSaZ9y9592Yk/4G1dTKCettDAwpjne5sKGh5qjoqWplqnkoxh2lq
QDZ/7PATTRP33G5np5GU3nNZF1Jql/gQ1NK/xl1lLsDkDGXTEBqHijQEjFxke4v6+pPkB1cDEt6M
/w8XkZgqWq26f51B3y8D2cU3ABnpgCaOF6HLiUqs9p9EI1nY3cnwi7PQJOP3BeTRhIABXz93iHo8
4MvKJoqFeswqDIoNkdVDB8yk7AIfL+DjFFPAPlQYZjDxCw3ZwcUMPcI7KCfTLQ74IiMjq+KdF+F+
YGuLitBLL/6ONXybPjF4Lfiqbf564IfAXnzlTkyZKOkxC/jrs5bpj7dGAEg0WhQtH0fBQfaKlOW6
k1gZ1h5e7yJNUsQbJlw/6i8R6MFf0BvmT0sEbLteWTbwfu7+ERe+9MrU4ewSfgL/vxLtrknP6duN
7k3GQp2yikf7SRI9JTrXLWY2VO+Kek4CpMc6qSfVubO+Pt3OOrc7D3WJ+7pp0PFV2Nispka9xfa9
VCF3okuDVMIxBF8FX2t8zl/Jbx7yX3wSrRRkApLZr11ht12hiKdklFSVSzEa7wMmujipje8YpgTR
UHip82t8mi0aEcu5IdJ2dE0i0OuDMXQEIwN/zlRT7aeFRjT9vQRJkRJ1VnWaltxYhC5yQ1aN+nZr
/JzW8P3QCCRExC15wAucPAxDKpbf09twua6cnzQY13iDl1HgQkR321mwyY5BfWE/AUYAl02lmJq0
AxJmXLAbUjJT2VwGgaY2euKkT/mkoyX87dB9YFW+QufyTv2jokioXFQ23TlFHx8mEIs1wKjgBvjF
IXcDdDSfTSLeMmNEneQCdc5LHvDFG2LfLgVaeU3wrbX5VaKPir6YzlpWZV9zrIcvlCts33fR37Uf
m9kn5of6EImnjqZTwMKBIf69C8EpL+c5NbI+5RJGGDcOrekQLvBzY34rQ0KHzG5GhaW9kyuxU1k2
P+mAzLVF7eNy0YJVQqiqANHS4bwFzokf5GThEcPA/zQpBMa60XlgPfKHN0PrMkLRyGhwaxWyauwf
TM2Wxtc1zspyADF1Lmx4Dx+bKqenptN3c+fu8QivrfSxguc9PpSFjNxjztlqEkt+A9DBQWno5ZSh
pwITePx0aaFahlA1xEk+U039LxQaPZNXyRKp7qY1rhA+ptQvwPPz3oib3OKZpVBB7DXWWzB8ycJv
OkUb2+kN4Hc3JDtbd1e+pLMwilTYD6MY7vsITYNmkJBzx3jcDC0rFMNBV1bzPI3tPRfhsEvGFx4Z
M+/6lxdubtfy63fySBo3y3Q/By5snCL28CVPrrNJWc/KUGhnb7cWWYAzcoMvLtsk5CAE7tUHJxrW
FVjSrf5po1NbeF6vKdvw2Hemr3YANgvTFVXMFoDSzjGxxkUePytp0YyMxgmuIbCG+5e3rQuXVa+0
P3Zq/HvLGQYmmZbs7LXVtmrlBW8bve6qmCcVXxfbxVf0icPPK2zoMsyeTAQ9qU549EIIGurscccp
75yqn4K0v+Mrf9MleGtzbbbGTIhKo2YJZqbysmwVnqwMKfXr3i0zQ5oX3sGRYqB/101L5Hb8WG/j
KU84kBJ8jd6/KOcMlJonQaysXEyipFC3hkAbWjWF24VGW8AEk8oDEWW+3tqSJ7HsKlp6tUhAZMbD
tIrGVKqzX4y1BBRwUJ7mtPiw+PWPEjd7K+CCq5h1J0HDrbCByd7TpRa5//qvw7gN5ls1MbyxExQ7
j2tDT3TllGMWcB6s2HAgLMyd/oJx0K2reISeWX3TcpsizJL5X07v2AL2bX/nBgbuC8LI9gRSMoFW
nEGtUb3six3n5nZQKIsfwuZWy5qFnr35lU7EF+rfquMsvQlNX0bSONqf7rnghU3xfCweFS4/+CVW
9DhSW72B2gkN8ZpuNTws/AQTIbUzVSI5N+L9RJe7+EXfVGShBoaX/l/UyLnQ4eGbDnicVrO5xc7E
zHg8z+Ht4RjH4XkWFN3S3g9AfO+uozG93ENc37c3YsaPCAjUxMrBAYOTUalU34rUIyl2VLAHGer/
t+e5beTt69A1SPp2Gb8HaQZhO9hZuxzaJkNamNiic+PyBrzFxCXQ1TMgluppG/naNHs8rOgBXgV/
FRTt6fvDAD10B4HUuoutFeoVZ0DZ45/gVJbcPQvya96ijlo/EwTgW0qIUX5FySnkC8vwiAEKcK8I
2q84roFvpwdo+GRS00GKUteGWwIrXsbXBLQ72XX6havuL6dDusgyHsqfJy7yzLCPANS4TiExjjkW
/2YAoKl2m34J6dOLdfbHfA/rPD8n+PEBQmeZwnTYkymecBheQnk2kI0J66slo12Mvr76ldUM7TQf
xiEpRM+e8yiP5Xmmp3fdKvHfZGe7Mlsyr7uG3lLXdeHHPEcb2VeE7A/eAr+LPc2SRLcjCVgJ1cT5
B7s5oeHJCx6jrBKW+HYN/V3Y6Mo64UKVLXKvNjwaoukDOGbQAXG8D4XSVvrrd/63LsvjWtZHAlaB
S+SMDa9LypE0d7tzJUEyrBHxaWoKdMy7Qp6Dh+KWQMq41ofDKXQjHQL1FgdovSB+JB636qEIbtrH
Jh9UXgrY93dIWsafKS56Na+A/I/CEt8ll6GQZa4KMnKUPRtRZFWuIJ40+IK6A97YAXzYmkWA57uE
pYQXaD3KPNYQ4zTzOarU1+TKBoqv7K2ilbStRPiS3E96/px9ub4VP45QU7fOuiBoqsQq2wkhZtA4
4XmJNqlmwvyxwSWDfrt1cdIrjZVs6vIT2sMu/DG2Fp4LxmQ7U6hx9K5wJf1C7YViUu6XRSD+iNrK
3mzkchG1gUe9hQ0ktiulK8LZlR3Uq0OwprGQ1jgR2c18eNxB4F11DbbYyuCHM9/LEo/lu7V+45CS
O37SVRHurSbVPgdIiilF6He7NKIuZGrZgDiPp6hOf869LrqCVse9/IHpFCt7YIFkKNSZq3if0cnM
Pjm5RHXib3f+J2MXkF9+cOMfKvuVYeglIRg7jrNL1RAcHSDPvclSGMZq9G141wIms5jSGXPiUA4E
1s2l1r16KQIk2oB5GmKsX2zdSCyb7k5KIQfLbLeV7LpfhWleMQQXo9Ap0+r7cEQ3e1xUcxhjErHh
LbJSLILooyPTRrgrEWAcB3Rr9lxdHes7oZf9P3ucOEKJ1Pz4qoZSSDkMUZIsrQCLMPg9oE+xyFf7
yUtt2uRC/lDbiVDv/JPNxbxjjdEN7cFPjoS9C3kugMrqZzjHjgFqC7o8ydpm1tVKSVar/r9NT6kV
HVs/JCI386zWrpwt7XbmAqJJZwREeiox8oyo1MiwWzh6+V5fy1iC3H+ocPgzFEW+Xk/Pde3942wf
I1N38PzMAtc2iMPalv1LmRyZWZCYwV3a7MWPeX0YyXh45SwJo2MyAKvDg6Fvo9ygLG8CWzhqzAly
u6nDqskPz9HKfXPTofvPfOAVrYgGGSfeWqifeVYRR+Wz5X08Jp3aEfyMTcpA1Sd2FciamV11VTie
c9qITAiSChg1ph19vO/6a/IoLix/kASe815UkoUFaikPbaq2QXa69stWZGoomrWUWElOZLO50Hiu
fsVm9Dj/sdAPhfLYxZkwqfVuT59hmuqaxeirnnnGN9r7R75dDTWgjU/pFZxM6jLLbpDosOx6Dblt
DuK/K0iq/MxBqFrLExg02Coa/BSpE4fDejJGckSoT5MULpADSPuH3/xWBqZ5XvNsKiROrHQ7/Z/P
UA1QhtL2Y78odbjGokqbaqnOBTvYVX0i/4bRzSZacyJnijvr7iYif9Ima+ehBtiJoxAJC76p/w3g
muw+CYvslgmbOrJaIw0i/n7lVouwCTipTgGE7v+0KxpCk9qM2uZW7lK3ju9qK7lDebTNE6yORq1g
eGvzAd2j88fsyYLMWdXvJo2O99pxt1CvxdXVBYGZTBn3OGixK+GlZikH47DWxBXf3LrGLGYgpco3
SD9MAUElxc+jQpDgBfh4C6mQHB5qYlIngRCnXKr7IvIKoA/nM/8KDjJZJjrJOEnmEnhmcYq0uetj
6Zz9LMHchMPakK2lCEnq0l3Kg09vJ2EHG2z8X9KO9XJh3uNyUB1I9g/dT95A1XUp6qZQldbwWEAe
bzMAmUU940tDcmj23P15PQ0poMwd5jr1/LsaILYMCf3yIoq60vA93uZXAV3btB+B3u8S1DE4v+Yj
1mcBQ2diXcnBcOV9SezCiXdfEvCmdfqf4cKgC0V/9+Qwj80vlNkncCec82nzreYmpzx7QotsO0cR
gjIeasYZIj9YttmMjKRor0R8bPXycw6P8uRlODmRAZKevOHkAu+Js5Bcx1nWGMG7kdJ8YuGJrotF
xBhLQe56XyqFHBHfOQt4n7FEy1FDfXZ73KNXwuuVpfMJhQzeuDZrwnEGRvevWhZ1PnC47bvPcI/K
wMX2beMpWKAQVudJWNrNNDGmalwtu8ID/1Fi4By5qw/C7kSE0/hSnNmQCcx2b6kZcWD0ZIYd+wTE
i9BAklRB6p/Yk9lLLMuLmeb/4tPr6rtlTy5lhWF/hc/T28OA2yrBpUH7gI//FwyTIP71Kc0KTEys
vYhQNNLQW2TaErrXihaR5bALZ8W/ip1PNTRWZw+Cl7hQqsNHy6TD8pvUbN0f8qmvDyOevPh/N805
cFWwuZqYazVToNxk90gy5Xq83LDejwiXHbGaK0ekloD0swHbp0DEvxqu7oeHEY4nuL380oJYcQJv
yMQd6HWnPMPvXN74utDLOelEw+Ub4BqR8spcL4rwENXowA5+Qav9+IE43ep0vLN2Oo7CaVTpC8eH
Glezf/O0SREkP/3/F6lvd192vX9oxwAUuuFhiCQeEAX1kDkFpo4oi+YuWCdcW341Mwuh/vhwZ6G6
Ckgr8AzxgFEgkVlO4VQYgvrJ9q1PnjK4gRoMwGFkxGymN2ZFHIQiVetsfYkkKAzF8o3o1pPkYDq0
2uYgDmf2dNYVL+4/4CkoSX2WuzxCQn8NDqRvhSFUhPf/OBHfmzZY2Cn8g/adBP/h5HkDVzEQ31bt
pxrXDgopOj/y4AScAotDHzQn+2USJXvcJ9AHa5gfvQL9BZKU094rrOWUHasl2Lqxes6NUfhO4fht
HOGjcwonPyV6SxhjAWUofJcvUBdk2VxufkB44mAsAHwa71z6lBlQO6Tc8T3F/cGUE3qcfqhupJ59
COmESwAWOmokzDC5ite1HKeJhJYKEpvL33JSmcg8UBOYygl6brRZtfPTqq81B1FbysOPOpz9djYg
QaTATKH8OD2RfRV06aLnhjsNqn+HZcZ3NIficcmTguQAs9sxrack0u3QsglZYHyH8otw5LckVvxY
l6jJ95LrFuLyTjVb/BPkqs+o9+pCs0wSWNLpHsxif5XQYcluRUnvQKgm1nyv5ti6ygoMhF3Mv5a5
sX+esyhvW5EJ+c/Yps53yOldQ+g9NiIX0dHMhqwsjVBi8/phHXdffENfGrbffEyWU3c+Oufr17vy
2Ea9qGR7OtVnkn2apNZUGtPn7Bggla/IVGiOrr9aEV9RKuDg2hJp8voJGSV70B7pE/4LL4DRs44I
iAK9TYzSytMmUoYIwUdeKUxcOkIHPfyJi8q3pBPTNI/Y06jwrgQcWE6pmopZZUc8BuOKx+4roFBw
E7C3GED9zxG84a5MO321ACq8mRT/IKesB68R5K2CzqN7SXcvHVGqXG2NGMcfbZXOqLTbU8SoJYuu
tkmh0VMIU5jFTdI+qdjlSR6IjGJVoq5Xfdbygak1RzW1MmwIar1sKYdzkPu3MoPwJ+d4gkipTRxc
VkiS5K8gG4MF22hnTjOxwfmUNhKqb4EG3lVk8EsBshq6bCmZAoXn5K+nJN08DJlLQN0wwpOYyC4l
F5d+rOymVGMSuy6GTw6JNatmNLm7Ds97hziv7C1O9nflVvDsKhARQIe+XodRcI6vKVbMMxzHX1KW
KPzhc4kfKswjCLB01wNGXYsSlTZc+0NI+Zk3CMrTVGLx4iT1zE6RiV1fnRkpXrZUDxVDVcybnBAb
UEentMT62DOvA0OlQiIc1sGEqWLEMeO5S/Kq4xfx5tV3CTI3ryqrmdMXlj5AnVgNLDrU+Un6xO9d
WFqYstRSbSY1LY3aYRC7UNc0VY1o9YJImb786qpUtyw/io9Xuyk3cTXc7eVNXqsLQba8S88aSbbI
yNmOCqxdPRmN20pggIXIFvW8En6SEtAdEB+4Rk+n9+YQonTIoJvUre/Tnr5vg1+57kH6DGGmzOti
yD2eTtL6zZunDi5/YpDM52Ti8S/b4zcrnpIS4SCSZ2YoRNtLLFhqrYBbSdtOWlVEE8oBeUb4h+/F
mafwMvn72W7saC1QJjsXaEt6bPQQA1hjqSCW4PgRemf//nU9WPj0DExYsoUpnalOSC+WpLaTqLz3
RV+J88olNtO1g6rklFdi4BHH8yzcV0K+9et4CpB4WjtVCWwmRugMIIC1IHCUBflO0TGUzGlKg+Yl
jScJ8XK/rbQ6UkcaS63E+Db6XdM5/l16oBL2EqcMmN/SrWp1d4okTaUws+b0lHCAWUyOH5xYhx49
vUpZaQ6PSU0X2+oeOXSNOZc9FXwM18doyWWI+Y3Uf8x71LAjnFgVnuFhXwgrQOJwC4CVsrnol01p
1i7t3mQ2A7yKSvVobJI3HUD87gy/NwfQVX1VJvvk8T4DaxIMbAWnHZ6T0PQEoLAqcnhi9ILcLVAK
99yjd13pspWgoob1c8RU6lhXmhlqpbYSKFa8NtoEDZ1y5oWeaynoAa8MytAVjbQ2qKWdFTTPvPGd
V7yZxNWVrPKBVYpgrW9hvUi/XwscOQd5VTCDxKtDBoFff2z/tx98VPAo+RcYSB1gx7Jxyls4Fxj2
N/om0qpc0mawIaJO5aXCjNSLZD6hXN+CX9t/D976L+fw1DF9+h5rBq7Bwq+s09UU93hReOfO6aFh
XH1huAxb5TapzqUL/sFrJce570hwUlqfwNrbCSmJTK5Mlk9K7uh1whDnbIMHdgQMZITootEQKPhd
x9+R7GxVT5+XAM9bm3clWGVAlCFRP8DmzCwr+ul9uT9SqaA5PG19zsY2gT+RdM5hZAcFpgsLL8+w
2UEFq45LjEaButMta8tr/YSDuQxcUzHZO/i09oRM+yNfHNdUQfqiA+1rWd7ZhVcfJfEvGLQtsCr4
dUsfbMEgOY5EmtbKiHH6zKNLMofDJe/4Rq5GONK1EqyzM1gphemu/uWXxL52hqe1GHtU3hbTz98T
JSx5tDEv7FSz2s7kwEz8A6MHoro2+zyBLTd1QZXSy8XsG39LG26fP8tqxg42upne7LLj+VmlaADl
6W6XQkjzFV/6bHYTsbvApY9SD3oRIyGdiEaRTszDe/ymwEqOL/mm9oo0SBAu3SzyyeI9ZrR5ZOyf
aP+IOOiJLwfrkP00cxhBEGuxAFuCQlrDhe2XIyYWzIIAVDUqIPWE0e70RrY7gMC2aDrFBL790ICG
T11yDUk4ooKm31DMRTGYfy/2VnZm8daBv7q3vhbQsYz8PsDeBqm8lYff0yfr1c0L3Tb+f6A6xJ0h
oeOF1TJLzdHFuOHAjOrOoK1vduSsEEblDx9t6323B9pn0b29L5LXDougpLQsy9dOLL7Im3FBMr7s
uPhHCMJ981zTEhMcRwaZFV5y0gTIaNrQDyNUiTJIvHRGsVpu1MpNZdcTqb+Va5njYT538DuaJV3z
v0KWp9XYc+Wyxq5I7iKb1R74QWoQ2xfSfipkatHLYghcoU7iHQPzE4uaDkMhEtf0rS5C+HCJXz9D
V1Fx11weBJmRqgTDO76uTIqJnRW3d06GaHmuGz+0pj2J6TvUIwdfRNznHOziFPeCZ6K4DEpX65/q
WugDP6q0/O75fyV/h470DJuSVK6SyQRICjL4Of1MJiTNODUBwgL5PyK919PXCR3jeNumbMNEMx3n
C+u8p3a9p6MJRwKwqujlCs5ISmV2V1q8DdoP95mH0zCtZiT5Jv6ev0k7uvx9s7wrMKcAe7DLlmaL
sf8Pp9Z2/wdsMj3FKvZ0dDPFRjmjZsECnV5i3EW9L8jBs4z51i5Rki3YPmZqJoxy6O1+DLOuclPo
sxGF/DhKUpiEeqWjnE+JWD4HmnqbbrSdE2n6UyrMZbbWbOXfMH/v04qXPCqbWkUGrRIfbYyOJoKR
ghtcdvEdeKjh9q/wiD8fuidXidPiTVjHmBfYpqviAJXOLBxHJ/dYQ+E3eYLS6G1xe9PhKAwj0g/e
Hg9cr9y2/mPlRKbrfCd4n/GWr/yEoD/kakWeeWmdPjlg+Wv0RjNC8TnNKhOYH+BZHzZ/ltwk2epq
YUX2UUgwEjHlc+2343JKrZH36LhXzz4DL8YK6c0qHO5fzv92m4b/93BKMPbYGn4TCKkiHuKIHHtR
fnwRNULJUd5zvGqm7npWvXKmq2YD9F4o8ow8ff/+0cRgZ7mquDf6UoOjFA9F9/kzeQLgeaOhCCBb
x6MKe9t4Re2KuA/sEUS2o03wK3eDNevtpK8leYFRtBeMA1rVpiK/wfBn64nGtTXpdFfufouH6wWU
NAymesqse9YA0VAOZltBOazhs7WiaMNoeIJz4aRCdjI70w93oNM6MLKSxofS165ABOs9FpsxzDL+
/Tqc/gGKLYO/0Om8ZdjwDmIeYAVTpr/BGaqqtAg/rN16hFLjG8VS7cnK73WsBihDWNGeSCrvek/A
lmsVo4Fszh8Xt8kIELLUYKd3roIHm/uJmISm3sTgRj3Xc2SXG5Jrs5bfai3M17E4g73/HwHa2uP1
Du9PdWLDEHdTuoYGwGlbOt43z1hNdN1mSWd+iFTe5uSHkjecZuQEfqSaHUTjP+y/adAHFIZXa99T
ArmNt2gdjrScZjVjGo7arH3MMaCzdXkLU0KVfI+5NweGAclhhTv3zhHOECJbFHCaKtXmLfWctvnC
9hV2L3VH3Vaj0j/pixF3hgkNTANBP/XTYlvJU5XFmJAFWO+kHmLdT0j5CGfjvcYRShusA2uWzyaT
A5JgaJfadJpCN8ewLtDF7W8c/d3Pk4FIyadW2AP9Q/UU1RWTcsHpKcd0ynivcWA3wdvPXnfu/7bQ
2MLJVd7JLECtby9oCMBeIM54xpeKXK4A7ev369tt12UpebbqAFwYvihxDDTxJmoy8NVg2WsL+Web
MBDYVux+w//F/MI3GkU4OCIzqoPBtsenLMGPuotytH/RDbnlH73RQgPTxoal58a2/6hEilnBCPEp
8uNftmD3X3NQLGxLjFDvk61Uw9HSUznngeKstuTWEGrEobi5kDUhLKQDps5YR/Y/E9tyP3hufWR1
NUXVKm5i7NzXXNZqD3Ib778kK7BnDy+z8Aoh4ixmccfz1kpago/zjSnmbQsmIda/KRUCpYHoWrDy
31nlTxiAySUgu3uj9vf4ABrvqZg643QatsGlrPfkldmWd54YW9InK1yhsojgjunB8BClrEBU5G4X
0cQ21NMwuDGXY084E/JcDL07Z5huhysVN84QAoqiP4TBK4UOZaYMB11b63Y8lv/DU/0qyuMaaCW0
5/4byRrbPMJM2wvY8mLHtonJT8mzFgSrBdMhBv0DR99tBHdTmKP2YHRWQcUQnVHolG7v+HKiJtg2
o8FJPhwnvskHVaxoHQT2f3495sCbZT53cBpUojBy+ZbdpZkUQITbAS1/GrF/n8cHoTllv9wjLCZQ
8VSEXuo1riODX8fx1FAFQB0XWoO9+3NGM8ZK8S1fEFllomlZW/SkQb6yduhpCRBmHjZnSxi2/Mwo
Ul4RLKSiP4qKtrih/YoFveaXfVmDFT4Vs6cZRXY+6nD2yv2nyDy5Eel/6C0qh2U90MntAu3AhVp6
9NSWmj96gKHgCeb9LyghVpyDEg4yDkWsjKsfEstzjNEYb+UCm8G8zxijyP/9CHKnL8X9ohlXkV7f
1OwokMEB6WnY9zu2X+RySnlu+UKJyGrUnEJqq5rEkvLUK3LuyOdMCSCF0G7haCi5GgKAnB5iY8uK
+IBAmg2kGYFjMKiWf6pcrEuKxtNU21YSIs0NpUQvxz0iKEByPqcXl1B5hbBunh2UUsRfMKUIl1jK
lkOr1mEnyeKKeGC8I4TvB+MUU6XLmB1Z3z4Nk1tiUoUPdsZS2k63KJ7v9+KP1GavpbLxmduU/XUl
A8wntcF3ITABvOLb8oLeH5AG01W9wtPjB4rUsP+gyRu0YTYxsWwpQDUxNt78XtFUtJUY1bi6g2WN
umYQaRvMO8opZOHDMBdVgQFQ7HUI2g9wt6TPGZjb2RhoJQ5YKgBXKMXgdwCdYNdRT9f1dOcsI/jA
3RdCdFpPRHaI9jLQZUAfdqq+nXMxHu6PNP8P/sWp5dbYookOzhqEy20m9MEL7oIKnFyP+UTVzE5e
OJvXUL8ogM/n1bPd4S+X2Wh4QHeTxWULJumesPy5m9uqDACP6dJu4FVL4hkPYBu37JP5DgUByJB7
jv5QUppgfvRlzC/sNA2nvGWaOFAcbO5ojZGB6uGxXFkxlOBFPJkoRUG4OFkGAS+Gu5tP7ktWfAZk
d/KmbEom+KTnoy1wX5XcJIrigdkcWsp5uCCC6Sh5PuEfjy5wLLzmavLEhB3XsYkj71+zWuXXBVOG
BpH/DnSbbHX5TmYI78Zl5POyw2b/eILJRkeuRooHqYESLg0c5UX09v9hTqLRhtPhVNOubDZEXLp6
bFs7xatHHsS5urb62izx+Fqulew+Sx5dj68SYCdd3oOB8ZVx+oV0Ue/tDOO+Z5U/bp3pnHp+8Ulr
UPPQoNuUonSYtcTfGKFXzOgbBnd/6HPPMUA0ZIlV+7QttPxt/MlcoMjvfUhKpqQHH79evMMsdj1g
8EltXfYmlJDh05oBL52goqS0wnZca3Fp1y46al6MEv5hWLzAZJnnIOKHCKz4i/6DXKdC5LX/mXNT
lmxS5GIf90sxGW1JYP6M8K0xT8xPTpEC/f1oqBMpIuekqmiZUGjkk1JQm+C4CzkOXFwL1m0c0m6t
5+dfx2cyn9XYbNMu2C80ImqGbiS/0JVz46TSg5C8Aoic68vIdJtyRM6WYgZNU9YzuWerQHbSeAO5
bChqm61b3qxHHzzROpr+Vd02CNzsi8pZIhhBm/HEzVKePDO8SGFKLWl8ITRq2bonkL9LWxc9OwGR
R3r92F6oXhok29B7KruZY132sFLVdOacmB1Bf30iO5J4A04D5oIpPk+j7PWXHnJIf7CuV3dwrODe
aKzOsFDOs7qMYw2XuQNfgipyoQlQ4leIvL9vwC/iuslDVmC+LDHZnW2yygRV6VYQuR8Pr4S2rOJg
QSfkYZqCx2sNWUdqd7tVLMSlIhYFCGOzy9g+tp0b5VsCD8R35t44PyDSS9Z9plGvzT8tIvUEiSFk
gBzNI4xZYL59sHvdkCYk+Q86wE4vu9SnN7dsR4moeYKH+cGxK44HvRfZyengzaVsMdJge9lcsA4T
Fwjys89B7cY8dRqVSpK7KFWGzcV4b0zVaN7Xo+ozX0ZJyUezmIOuKvHjHSBALzzKW1o08D+ljB9w
H134wYKIEOljV36knjjx2z74lkBaT24YvqHKWBliuMqkJR23601NsfhNK70AKc1OeYjrzcBajPFW
ky8epZRdoUj4FayBoH9ZTTToRpnaAG7Sw/b51G2xz0OiJ4hWjsza+llDRaaMi3aPwSOVZiF6M4R8
7GSl6nMzHQBFf5OO6zxMNCPpisoQGjzq1LtWs8in6g3VCUHquzUBj2D4FArDTBYx8mCar6NhYvR7
eXiS8nNPzUJZ1bd72XeevVHUwKOEjYviENMUIs7OmFfVR59KcvP9dPhVAf40776+U6/Wos23ncdO
ld2aFGZc2xxZ73fWwKXPik8ccN8aW+8omFmgTkB8yD4lXFKqgaV4IeQ5KUk15l/iAIaNB1uNtqWW
60Mf2tJIYdgmWO0c2CQRZs9OXVzp8Vt1Cfdg7L2d3yCYNfBdVDf5EQO5AxpjU5c6nQDqoL5Cx4kn
HKkc7bb61pMPx6okm33uH9FxwdKqXf/YXHlqDnAU6iVwMqrkeyLzYPKdOGj74dS4321AGdaNwqxU
Gpt/8/nPodhHzhArU+z8ORpeP26A+k6lrT1+AjK0AyAzOrNL2/U8Zt+8wqtM8zJHAMhHsOqv/35X
S0K1qxx1jGTZVT6Av5vHhbfr9unmAI9bncxQdlEoflnPHfvWZIYBK+oXXfulZVjEEJs6ztLUwodj
zKTcMhrDdil6jcpy2/ObLNUxQJvIPiFPt5ec1oGD0rjNr0LiNbi8M/2I3Kv7q1WNMuMCF0BOU6RO
SzpOuqQVQ1rquHl+9FYPWd9KMDLlXqLVV1FViukQge0eRXljjci9Nq5Rn23PO0z80XZJzjjLDW1L
SHSKAGvkahncIOswkz0mi4LXNtKCuT8ay9SLExWYHXAXQfdcw8kA4u7KDYsEgo8s8rdOmhjIBFOR
U5RV2LdklUzaeSYf1h5/SfUwYLMhJ/08vWG8AdU5XSNMc2lOBdKmsI0scrFZrMCrhPRiPeq5OIS7
VVd7WPU5imed0eBqtIvdmtPxHJXHb5Nsp6UXfeBQztmH5WPIGTHGtVrVd0xJB76jPLdapTxYOy27
QSCZrtijvDuot4ZVXvcKU6Z8hqCbwD/MfEGthVZJ6aKzO5dh18Bc5FWnarSWQZCZzb+z+ctKpAxa
eiBVdX9mgjzf6jMrTU4ftbxY4p39i5NBXDGRYbY0poaH9xDv3cCFdYv70uCzllqE5+L15OJV9Owf
IR0i5QPgmO9UnI++AeuhZPT5TKFfDLHj5z1Ih43vYT4lY1Bjmkk5/FAKUd5T0lwshm0E5tAElnqI
zPKD5bDdtZg0fMxvP2EuJnODeqkwidDRwUkEV3eBHTyHoJzZ3XDAuC33Gtg1kYcx0sMxDVo6AB9A
CzRNItMt8FV/vSdx8clQ8IJE95eAuaCXzKPpm2MjVU/wzH3TLTjv5/NA2lx3gvS6hKH53ZGzGS91
r9oizIC4X0uZFlzYjFBJHnnwKAHxEt94HXJ/tEzeEsx3/32tTyhjwZi6pWCkzKPlALaK/4F9PbUK
HbfdegHlungap921Z/Bu5PndMq1TDB8Lv415kOd38KA1cbYBcSFL2HF4q/rWrvFQtwLfE55VOR8S
il26kne0qQR0vNSZsrpdgnwHlvo0Fj+1ObbsciJUmdUqIjLLtnGcexWFHJ58nInuBlUedDSfd8F/
8C7Pio2Z0tkFDuUMm2V8L/ZaSXEiKoUgPYjTxusVIRWuEHGX0YFJETQICGwnTMTc0LhMHWijwf13
U1CnvMZaJbedSZHdtud1MoXiyfbFntq9NZAsdK7V6hhtkctlBmJgKbpDmOU6AoVPM8QMMGfRpXdp
ijob1Cj+MRzon23LnGBG/ijhI8ADCeUDnnIdzl5tuehRAH8+UX635k01uLhoBRkbWSxTG9LNtEan
nFR+PymQfD1Q9/9EIkzWF3YcuyXEgE4sve3CyYw+B0sYqDF5nE/yI/ODgL3JOq+6r9JmMU3SFfZD
69nKkGpwKm62RAUuND7AtmXTpkHG3wAaSMj4+BRV8PgpaubvLRigC4mnBPHP3K0mlyn5+m8VWQ6E
fyxmS6kUPbtg8E7EHmx9Cc0sW0syMRiRpasuY9dt+1T8S8tA/tAo/vqxPJUx7br1dGNBH7y4223F
G2o/ewwoutkAwvGFW5XXMdGj3aAVdkWfGJS0RUVRSLoZc/wbsYDPf7WnSqt7za3YTVs35Li5+v8Q
ZhT/go0JkdaWaZPPOfnplXa14dexGfyDPD436jum6dxw68hcvjLFY+TgoLYw+doBFMJ7JCiepzNE
3mdy9M3ZIsyMo1thQIOol5ceWlLS7jKlUPjf97IcAgQhYiCXRxAyw9ibuqpMSTR3PVs5+0C9zOiN
KCD/SKlkQBbV96poe8i2poATROaWjIjcQNaZBqMkOGIQ0gKAuzdbScfh3wcRbt8PgKaSIch0zFTx
Ed2hVYtc8fZ9W3QFhCVr/t/gPC34qKnPH27uQ757YSDwwrxAhLqdu/6SMXdibNabHLAwBJIQK8op
XFf2Klpbg1indPzDctGvJ+A8kRMy8+GATX/JkKfD9tdo2OcOEht8rMFY5Afi/hOkAZB528nlNqyP
LhcjFhU11UZcivVRJnehvBBb/ptyeVN57RcZ6hObHkNHqj3Zqg3cVRB+h+XGFIKF+CaGOofs2kaq
UwmE//MN8fBPF371wXmEOhtpPI7gubF6IXGEs/+480ClILl47g2paNNLHr6YN9IV/duercEItFDD
v3gtBcUM6QIdw2ZwxAHFWg5hRjR+a1wH/Ht1fWwYV8XYmjx2XDcVInHrjiD7H2Y9f/jF39pDHfY0
Wq3ePSvxcvDu3cyGScewmfZs/4CaPkAo+IyzaSKVHPqreBdv4y00VpN/vmm+laGTLX928SDkBmxV
vlpDL3jbYEQW2Jcxnup7mKTzIXigjm9M8pG046n6aKUNyKJgEOTU6eLv2yywJWRu9WyFNgxNbB4p
kT7tjR3jZ7eh2IMK1hCs5AnLWUvIMYTHi2GVD0t1oirHhNQFivmfqveETM3m6ZJg/kmFsQRxTyTN
6cp+E7TQBzGO6OLfFStN8oPJ3D4PrR1WXXPQr2wOlrdiyznj9VwmhEeGKe+wVwghMygCK1tEEBQS
iD8m3A7yZghstkiURGN5XQavLgSuRcu0Lm6GBYYd9xCf/XDsuVFHNoV+XI1W9KInRj5ylb3YiZP4
o90L1zwheLq4IJ+v7C1U9ASmuWIOHPoo/3CXVGWwQr2PXBDE5ijFDtHwHZU85m9u4vpCL+GvB8bP
MXdaEy3TfcLsu+/+I1L0lyb49kqkDqmWAPvvqfZsLNw3j090JueH1kHY8Si7Y5RfY2PbSzcrZRT9
wPZ1Q0HQLv7gZ0kIKmJiBImjqFNNnVd2j6ycZTyvJo6CrWTQ3OJp0yG/WEwPuaIOacJsETiD2e5+
aSoVl4q0kOspp9HluHeD/+hKIQ3UUnJGwd/OrUKDLFLguAYaRHwMS3lw9TiIHfSfH8hkBqwjH+a8
6+kaC/6EYbSMYHxLz1Ne3y4cYa/ppLprrbu1EN63hbPSIimpSAgigcwVteyknzRFsUbGj5dHYhBd
RPvOovxswVPfXG/8dtqaeamjFYHQJbtfDRVXdVpUnWNEZvJlZubaI3Pl3OdS262KzO/rT8CEdnGu
hrUxaRXaez7fh5J2ITbZE+sbcS6yKRWS7pJneltFbJvtCFPUVsfKV8lbtaudZ1Wp336vur3UTrCF
EVKpA2rYL+T+0FCC8mSmi2mNY2yI5ZtUOLGQYLRVsK7HKMHUCat3fZlpyI/HpCi9vN35D5wJIdj7
M1tc/6ZKNjlBZ93QGx5pKB93DHzA3x4GgSWoV2tlhSjZ7qpYuNTKLQOa46l1HGcv5FRGbntmnsJh
NW7if6ie7KX3Ty0cCUtT2Pb+s/CO6TYc3idt48hQabCAbAv78dkb53nXLQuxBrYGriIqohFp0+Zb
Vf8BBQLjY5Eaf3r7kzHqyzBoENJxGSLOsUO+ed0zPLw+aSu97YasTwPwkzwhyN3P+S95cL93yoiC
nOLCNXsEc+5W3XfghgzQvjlhW5VKJ/v3T7RB9nZzdYUEf95Pf1LGYClghtnHLQYFsJwmgwID4TQC
V16w3dekEJXleEjNl6Pf49UWzxzqmTJ29KcB0TzWTcWG5tTtvRHNJB+7v2MNuWfz+f/xNJARLLrQ
K0DMUwYfdqh/3YVBDIsnJ+btq93cpdPtGRYhXu18PmulELoU/cBdJJQCcbiosdFML5e+r8fKdZsS
q1i8zDrWKvQIscmqyXpnE/uBP8TkS8LWwPHm5xOkVAWUMC3D3ZQEyQrdOc9xpKfRp9TUf5vP0Caz
Vk4ln0PGOphEcSsb60XHUPa+5NiYTt4bXALaggjDVDUg28Tm3u8PQlO3BTyeApXqd2Jgd11VYOO2
6LjqT55DPHgLg1O71A4mVHiPV8mde7ykkmqSYzdPvRqA0rFtmnqu5sVrX10Ar9SbvwEycfn0D3jy
OwlFYnyKLbu7E3X9YVc7CNiFUncHJE3F1Sq5pCOZVF2vsNoCeyZgFiadsppfXjljgF7zDffFtbtp
SilY/GgAnt3a0eWr4dzHCDzFwylfb9N9+1zVAgHCe9QIzPjuoV96FNkUHCj75iqJ2a7KLGmjQIzS
ABGeougxm9w69js4cQstgkBKIqKGxYlpUw6pXEMr0HBVdlBzLapTEz44ke5pkLEKkIPiBSVEzTsg
iuwLB8N0WKEUxEj9k4FXUHNHlNlxfC7NiftFfI+H1uU55LmuwWAShEYCVY7cNi/pYjc+FGRH8SkB
wo8dpq5cqLKKTISDX/PPxgHR4q4Qasphaeb31oKB9+XkWiDKBx3TELClM7gCqhJplyfyUOdZOhRF
eUFc56skSogjsH9XypJ4fiaZGYr+MYdYUISnst1F3xuY/tNWshslgiuceGf6ZjFaaxCegSfBLdiR
+qOW4YWHKs75uC4973O+mXMcOmgSFm/q3wWpSqUVAWYpY7eKMgzonLQfDVh0DNkOdNNfsDKPcjkc
GIuWfwpvNWj68lOjoMT0RXySbxjnonRSpBoVaLZfhCfEtkUPS/8IEbZbtNmxjfqxdcXMxUNh3zdy
NYWPMIWDElaBSn8XTeakvEDwUSTHAkqX8pwuidp1W5FMXb9krqoRIkjXn9Owwyy3asnhJZEuB9VZ
AsoN46CDtGNo+CdoeN9YhnqaMNmyf8oVdwKctbfkV4C7u6Pnv1/S1DLKfh4G3ethAkc3XY+Pr4JB
1bF9nJI4Rx/w5qo2u3B2cBONY99AwFTLWMwinwxC90stcd6+fCaM0fKzJYI+I/93SQX0z1hOgn4C
XDdeoXZDYNqgFL+nXacnZ2C2ch0KkNm6fYlLsuVxgf9XQDHUQtdtcOkpx4s0lTygwEtwAE1vvQg/
RWae9FMcDYiQdvfwMO7einp1pEoat2EzKIY0ihsTcSnrxO5Ow7s82EAo55xLpChqrmCLfyhpQwYl
mCCNRJzluJ2mx6SItlhCXWjFbfQ3gkpR4UR3ajnFJP5i2XeAUkWAY0drudlNHXcXMstRL461JTzM
eLGjM/339EiZgfK0yW5N7jaHeXdCFafbfpjqFMC0tuIGj6D8dusd08326jqG+M0LDUNmp9D+YTVv
wjlZ48uJ7+xK4AbRTzvKEGz1aAeRTD7FOaSDcnTka/9UuGPKS2uZAy8RIufvn093cyBlVkHpSR7d
0w2jtczJYc1ruM1DANLzRrpC2wree3D4+txG32lACXZivv0iDSbZvf7FiXed5dneybIsqIa/VuSl
wGni6NKbEwmLosxAq1NfMsfoM0mx8UVdOGIdi9MgtAu8sZM6gr3jTOf7ovR40ktx8MIY12mduDwW
xH3fZZVP3u63ate4V/lt9+PdQfJ6jN/BAxaWVUPyik3WaBko3iCFVXErKtfp5G+gerbTqVS7EzW/
8jQb5Myse7qRWXB599XrReXYwMMII7N0djkIuBMiB0A5xvXRZxpp+NJ1PVIYhz4jMJbZNInXK554
dbUIQja9pH37atatyZJuBt7Lpd4ntMLAwv1G9TEkS49tU8THYM/Q2pGCNX4gn7QPjpQhPJaexk2h
akEyzbcZDI+dgSkeR9L9P11Bx4EtuqL34BgrpRRJX03H15jjYFLKqHSU9eRkEIOXlC1Zri/u1Ldr
md9ktEHkSLptxd1TRsSLU9hPWwvkMdMpeQOJ2k8V/wzLo95WHqd6LYaZLrTyx/mqx7jJpqAsx4CD
c6ybrijOfTali5guIMuWYDnpxKi4oHtPP6yGsDSuHev2ravOmnN4D9YrUBqWYMPJe14hY/btgljN
TBEokTnFtIVVnxFwGWGxkA/Nq+nIBitc6LeVBXFtn92umilOyZC9plmg5JAhrhLmUoBq2RMs/ZeV
+cjkVAVDE3Fcn35N9dGiiK0wnvYx4LbhA5xIk5hUHjPwXu+dOd0MLz20k7dVIzGIy7u2SGmFHNwT
eR8DkcYQAPAJTLmjZ9Ibm1ZgEeueJAgesJzxVvS3Bn0otIo+VlvhS0BOsZo/oysdZpufK+A2Z/89
YdIS5+XK26vp/KbWLoiO8h5Kdigo1oCecZRVG9rFmhzMj7DpRzKES7fzOGbVSZbz020MH/qttX/I
w8KsJpTULBrk8ors0PpFG2myghV0kzylzQZTq8yPAaZpigxGVCV7BscBhiAaFRzy3ZidUeB8yjZQ
oUVLjHM2UAmTwIHYApyMgd+OS6udVGQwVqnNJL9WO2n4Ypl1gIM1FVJ5U/aEEPKCSD8NGYuNDIC7
w2xy6yKQSzTWbsvE9vR8Ge7v0gRlXjE6kCgwjcd+NlH0UV6A/x37erz3RtPoi7+yfv7nooDBd2+A
AiuPkI6Pu28XoeSMq6tdHwP+KMHxQAng3FaDqaFpjCCTjd5smwpEktN2FNdUPjiWQogFXoJHuyLL
yuxB0lwGYewxhMmQp+jLy4oBT5lEeH5KGNrVqrPsKL8v9cV0PGY0n/0WPrDtcQQlRBE9RnOKM63m
Dr0LCu4MpF17uAU2rLf7W9NqHQ+AajDlkgZASExU1DbtJo668n2OLNI40l9vqpLfeotNBFn5X2MH
1aeED4rEJNKeCszJaDuXKdf5EK25WQ66MbTDBRX21O6O+ZvgtCv+B6weWr7TD0ihx6FES5qlSIyW
TyVX4eGc8j57zfALt4jBz9cIt8dfcXfOF+CbqsH0zki76+6CfCGa5W4dB/etfEgaRBSrUCREOlaN
g7Z8Eyg6xdEn66NpNM8ACvAMQx/atdArBWqVf8w3ixVYmkwbOgjBwui4Loo22W52CIATeI9CFO3Z
3OUyzRaGIKdnzRjzjXgXVwritcPVK//VXB54Aq67VdWqDy8Z8/XUOfYG/xvulXi9Zs2k00au04xT
RwuAxmKLWsV2mMgE0HQtQKFo3ky/HrkxPTKxEtMBsdGtkZ/nb954mC0D7oeWXgilgE30iZEON78P
YgxukWQe+mD6L1pslG3mC6L47yErR13XxvDqw7OTCPCYD1xJb1SpJVW3COsmoOlk20d80rAZjg2L
SKPlkGWgC29b9Bv//XmxzENngmnFIKf539rCdqsz4FDYL34IABxQqr/7n2Wd2kE7eFdM18ROnYUI
jiNKy2pYiKhJIl4OGuCu5znP/VZJF3YVc/iHzBMwKgKVEpqa8FhihRkJFB0Fnih2UgG1ElZGfCKd
e+polvpHDI/9YL83m0n4XmTzxXq5e1szUZnEXdtCMIyvi4saSodvtdyc7eEFQjWhPKSmR8+S+I8R
wGhP0zpfuwzvMXCs3MsRQk+zGjL+fiicee9ffQ6SQD9mN4nVXNihF6oL0xvvKGrnu4iNeSpvzMnd
bW4k44SSibZayAIYpgeKe2qAPwF0S5c/vTAF5xyRWKeXfpGF9xman5SOVVBGWRiqwpecBZASQFZX
3RrrkKTukwBNd7kAn2bsAlP4DAscYGfun5kFzpa7fXMctmDyKlDjxOeM+wf52ELPIntCiQwqlHbC
uKSWJdaUyOCemyJmHJd7tODPKFklV//06f2P3KgEpw5+CAWseJafkrAehYiW/ZnIZJxhZ+D5tGsU
H7Qj1NeoOvIfgwFbKobnLREwFp0Pvx9VlXyW+TbNz4GkMati0zbEG8j+PlBi57ZNuUqMl6GU6Dec
IJ9hTSwqLrPvKHKPZaGgWOcAPQLMdLoAhZLz989pdnQNI+AzqejSvyHZFqNXSpFAHoSjj324rjGI
C4jX6rnKjLy9OV4OaH+78Csp7/9jJ59L8nr49EGefz51QtjcCDR8iWPUo61WZHAjGZbETLdZyGxq
xjkGwrvKxv1mFf0f+rzipzM+JQPcV4nAVKHm2HacvXxenTWxukdnH+mX0Z6AS8UKradN9krUCqHK
YFnCallu65e1ebCSzMfyARxzZJFl9JONNAB5YgPgFbJ1L+uluGjeRDA2sIApeU/9DT3jPvNszsn3
I9t956OnKaSvmHbijwwGmznoMNcLmXkAjw0ES+HhxGx4pWwaIzKHwoTD2khbhw6yUOWTL+pLONqD
5PP5+6Yk6/4Zf6H6YC83mMVilVBlQO8AxZDf8+QYeu4CJLNqMD1kNyLy8hyAHc1e9wz804N8xHBz
zaTEt/HdINyLouSKup97Hw/xkE1hxIfPxyq5oE3h4v2Fw2oF4PYSHqYOJF1v/5NEG8Qi8Kaq2BU5
dI4mvgMfXrjjBkayxyJc64fB2huRoEeRdkqnQu47Sz/thAaIAZShkoWnQ6hrEajM2FdSIL6bmKCr
eaJQjnGSYdlZUOeb0/LUtor/Ww/m+2SyookOwAFIe50lKKZ1R7M67s+NEp+wzMGRzqi23JY+6uMa
jUgMbImqy2/8KlWVn4ThfQ2CKxhXUkWYVBfsrZELjEl30+5El88lKFayFIwc+ku6K6S7a9ZRo5CH
5yWsoe9xaldpHIvDXRlGQkRtCvq0/sNSam3u+fkYh3Tow9SKZI00icXM3Dnl9k8CmwVLv2ZjhBMO
0angVq1LU5hsfjGq2LrLCKreGq2PVUbQRiLxIvv1xVrCcjNjDZnSjqZ2F7gM3vQ7ZV2Lyd+KV7/L
ifNU7/i5xsDn57AEXNrFWrxhAcpgmu9PZUcbuhF6d81zdQNvdiTEhJROZverDE7xzhnsTrjteLJ3
jlvmTaThADzBhPJHviQa0/yJ+pHn2FdlNZU/Y0u84zTPRDaBFvQvvtm0KXNLBAhGzTRHcr7xi97b
eYwY1RzEgubPNZcNH+uiBT9lkOI3JvP8pQA4VzxPPdVFEQHlKDDoAYKpsENavi5UEFI7/PVPkEuQ
n+rDHA3moteqbgkUsWie+ZSU3rascfnYSiDLEf+kJmvvYvRYyn7EejeifC40PODCcN4qliFxvbMg
y6mALEFfq3Iyi1rfGT6hY6xSlxo3YIZzCMKkrjjZ6UkZX6AhzusJVuR5VE/Tx3T8hcnGS6OUIUmi
Q7c5K+9vT5KXwTIrdxk9FIE/OHLeBOlnITL2IWFEq8pQcThz5oTISgc6BgNky7hjrAkJu2EIfWvw
B0KHIjK9A5ClIrx6ZLoj3pidSQmKbGTgZ/uVQAMcGc5BXrKrFChV1YnjqwxqloQyae/h6aUSQs4x
OB+kObKH3mVifqXs0MPWZiaz/6I5fDKeP+KJKkOFtJSPaSsnnCmm0S8bnnQOjG4nvB20vvw1hmvV
Vkzw40+hAYWO7qIYwPI3M8CBvwloxGZ0MyI98Nz6tSDZeOg3NHNlNOEz5MRz6CWXx4ShFK0tCjv4
U7nNL4R6OH9nwvgqMstrpl9Fma7Ts4xdSP8C2EqUlX3D9yJoxYqEIRPCFii+Yc8C6gQFGmMAUXuG
DiH9ycSPW4TMNjKjuJBlEvAkO01WDczDk43yiwY1cNNmLebDqdmbNoLZm79hGXci9J8+MqLaZnrf
h60S3MOMj6Y658KaX9962vORo5gprAPLaUrswxLx5wdOBMregyofIHdIaV5BYAiX3SdwK67lZDJF
eAtSVa8Ww6ouLiGsbsOhY8bizBu/36wPhAcCQOvI0tXqZHvlXlJjxNfB5MFwNB2Y8zmaIV7BUzoK
Jz+I+U2s0BAk1oDfv4oUDHU47QDwsVCrXssZzVLLiJndPkZbTGICEC5q/xw70Z6pNTe1JyFD69VW
8/hI03u15qBlURP2qTMm55V6LFClZXvWQyRetYwwgzZ+lo4BWAqdN9byk07R6Pp46U90QdkGEOT6
HWXRIQRGFKJdOB1LQWneaac2g+iCyMVASMQ+278XN7F8iYgbHGGKW69VV1owtL6CFvoDFrsUxCGQ
6EMRxl7mE4xwNm2IAkN/iYalAyaRUhtkY45rG19cm0eAKhkAnykbGGYwYQlCj8QEyjIy7NkQJJhe
qpltVhQViWNk1xD9TJt40B2P+kPHeR3o3N+euERN4qbCh/XzW1hUr+Ptk1DKIfcb/+6TYZNC0Rhk
BoUxd2Q9zsHKBg4XU8Qv2jOZtX9WkXw66NgLbKj2PEDym5usPTxAqjPdzGdY1Z3mhCOFVb0SdYgw
IL3ETglSIhHl408Iw49uVB4cH9l7itOGAEUkOOcHzOAy4d5GSwsRG9lvKHRubK6VwnPqLvqxT5ju
SMq6oxK34ClbH79m2UKTJ/IJbK+/XO/A4jHVZyY/DheAZi+2AcHT/ZlwcgJRV843LW2Jchujn7UW
YUQFsyaWfY1HmBD8vVrlKO50KzyIUMs6U5sc5IivTb6z9FaRAIJHMBg9u6A17/ZVZja//XBddqq4
2bYVjdCkCJs5Xb8hmd3PwKdkIZ1+JRY5hDkslhtKd2jZI8906H75w85iqCT94lWPRD0IiDGYfZhg
Whv79cbhOHGLeYgFlNfdW31jqE9pNDVnUQRbBrfflB85PZX9Agr6Nm//3rBw6CwEpUE5CF3+wzDr
QExP3SL2aJykOhJwj2AqVofhmJO6CpGYGKLrUchydF4bGB2AcPfcyn6Xu4i9qZLM16CHO/S15UAf
KxI+ZwA3c8GVARVMprnpVSZLiVwSitCer1ETlFoZMsyWs0LagyFYs7j+MDu2chMUz2I9qxqkWRb3
NyKojukGGrnGWm1+eQhG0cN4efmYAGlX2JIMALCy6Ba1cNoKUoMgd+YhHwG2kaJH8C/0RBkTarkw
jEuIhHFFy2hPL6DavkETa77MZ3lYzViixsFfS42nyPruJXgIf8tztz7Q3Db7flESjgEucjp9BSL/
DDKoL5JXX9gBAzJJKIbqOoqYYrOUjXecai9YAHpn2h3hO+HPojyM84MhrNSBLnRDGOBoG5WBylOP
NdTpUlFfQDHgGUgPUY9teaAaRNkHd9fbmOthTObj1++kTfW7r8QwEg1woEsvIn/YhWX5t0iRUD8m
Dn7gePGjr2v5FdLisD78KIwuLcrzpZe0UjkkYMA+UYgLMBwu2RMWyc6TXrHi0PWPJ7AwuQpFIWxH
pCwLtDlV9p3WmsFFyguhKMiNCoajAHNydPMXP7+wGIZ4oLM7ShG7K+vCSFyUpmkJL1leiDitFpeQ
YKNV/UrVLJaYrPjNWhLlZLd6pOKfTP05rl0MWx6rTaj6WBXVQdTaZ8RvPHDWe+Ch4SQE+TNJnych
CSRxXw7xOa111sOqkQwjSsGYQm4xIh2/eZ0yGLHqPaLMiGw/x3OES1XaN472jo/LS0jztPcDIWGJ
j8SZ7UN0qDS427fNYp135vnAMqCgwKSHynLg5lbdh2q5KdVxNZTUC1CDt76btj22ujRV8Tu3q6QV
Pb5cwSEj0LQXSRHaOsBf6qMXSmkPAxLHr+ntTDNmR5rjVAHnj28w4CnMYlC3jOyZAquBCfln7BGl
xUNkC6z4sLo+2PdxRVRFsLsULbQHk7+KRHuIgrbzGUVq+TdmS+5xMt2XGRrZKxU7MZ6CVsHX+rCD
loGIT6gj2LcMx4C0lwfE6aO5g3ZCdb5VH19Hy0wZG6KAIveb2jl8dvpWPo9zUynF7bfrsXpjteXZ
IXnjOdUCEJtpiDQW09loSrtOoCV4AXGNmvEaYb/1WA3S+KMGV4ZYfIY6kYg0C5wUy1vnRCcnT75p
ik1/Dul6EgjR00aJ1EsPAJv+Zf9Gm1y7wbKxMLMmAuiqABFgg0lXs5sMxwLfEsuTmvew0A51Y4N5
DaE3VVpWIiIjrIwpTqWv61RMPKhyK3Cm+fH1+dYJLPmX/EBEczMdUB88vL/NrxoHL/guYccTSYwC
mQfY9ZQxi8jMmHHfFbRuyyKNGXBprpHsR32aYzJ3t+e3/opuQp8WYQAXsaAagy/5MEKSAQFssKDm
hZFCkSa4X2xXUbjXfpxTZ6KekDoplF65LMqrVnlHV17hH3qejdtOoL2BVgmSqXFCffr13xE9APqr
b7oFZsrdbHoW0dr5g4Wy3Tynu1LOKHpUWMIgkSdtwhMd4FNdvARM1Fm9w/RWRuT+AvGH8hjRm9sa
A53AcBsrQZwBocUkai6Uk+4wCnSMPMiR1rWPyE+NHu2hQfofFMcJTZmZbMcON8yE+MGThb03C7Xd
ab9mWc+rVqi4LlmeLWc3E2+2m+Et5YSsU2QGFZwR9PVom8ijdj9FKO9pP1ywfG2PF/0F9h80VOfj
IglNGl6Nx91TjFGfFJdny3INuuihh+bHW3QWSrO37NlcY6ML2/9YQfYlMehWNE5EWE2nStCtjmk1
JU5+6Nw7cVXeDcuCz69d+kYwC+bMD4iTr9GQ7U3lmZBBFKY2LFkSHi+SS8VsNyPCNhoSWjOnm6hB
o2HVXqt4MKJQSdOzuVDpIe3WupJtFdL7LdaOBs8WS8NmPCXaNSuWGWo82AhcymBnmYcylFBQZpq0
vEqH2ZgvGQiwAc7jp5U3B2MKBC0zqvYP6ke1FWLG19+SMRDXv+Sv0q1+LZWG6Jb5ms6xjt6CLgvb
X2yaZj+LFepkTR20Q1XKVfLKe11ZfKDYabzkoJ37Jw0qXZ1fJfids7/RNVu5RLdh0a5E7eQRcBDw
GLBsJacITJ2yheY9QqV+E4D5o10nvCEQ1r9SvjM0naVm9Gy7X9/u0kv6KacRb3f0yBQR1j9TIRXZ
bftEB2oZrIZRozMjFlP/5kgapHO7m7ajirW636KQkYXLhVeXYn8pVps2lblTmARP6NyiBTqoGEOu
WzU1ZTiHH0ercMISjYVOfldB7UfZn6uhxo9yFbxCiTkGDgrgt0v5PE3YheLD5kTYPdC7os0BVBol
LHHIOAYWAEBor5OfDWddtaxvV/FUM/TbNyCT/RP8MnlYfDfTu0zksXgZAYzQvNq97T3LRSv1YSBP
CL4fAohSx+5MuioRii0srjeZbzJ2AKVSEz0xggPNg3glc30S0wlCwtU0lRtpoMQ28v8SwsxcUe1i
5EcERbFn3CgHy/Cxot1dKdMLgBDEkbKvPLuMmu/pUOqhH/+8RNz9V6f90WWzOHlf6umeE/qyBbNe
nwkkV9oHV41Rnr0RYTG72vEdw26/mssPusiEnQU+sXWfcmOB45t59XT48bDelWd3yFxK5EQKqVmw
cLfAWAAr0jac7BH2Gg8AuSOS/NFbNy6vQSXcvL3u4dERhEdgtVdm4nrOszAG2bqYirzjhU2sMrIr
w4hz82nnekjZdnXu1N7oBqWlzGrsADHRcVB+kljj9mbkqi+rHi6FXNPTc+k1u713gH/ygDiPCyNR
SGy7L53q8Kj0IbIxsNWE1ncsKi5sTSmRzpn+rqMRx/e3Kg9xPb5WVbpkzvPpI+KLlkDLcYKanOU9
aMrAvKyTFUAakpNRuengik9BoL933JWZ0npWzTFVoC+p9s6gdSzwg+hwGP2TvMr1L8S1Yk3nv8Vf
vAEJNIp8o0XrO5Z3CxiKCH2iRBZ5l04YttY+Ys5p517x49ZdoNvWKgPrEK/15uBUBfDw4hpw8/yK
gi7JYWHxol7jUtf3f49Tlt5yIeaEB1eLjge1vpO/u3uRCwNqqL+pNC5+zXAkLw8440dW6kbJL2DS
4I6lOR4IO+mpV9xtmhm+i+O8nC4bg/ZomXx+T/O5YQ86dJYufe0RRNqw1JEYX7TGA73oVd2PNR/X
9ntXPlbFrlzQCtbi2PsdgHsECp6OpyWXeVQhmTjIYo58tOxkQY0Hl0AE5wada/m8ioHKjveyj7PF
C+/hFHSiwrUD0wUMf5iEmc7Jn17k2PW+0vHBx6nu4IRnh2n3Vn68MMgtCCM51n1cDlAIe2UsfcjI
vlkIJohENIAsWHzeh3AvL6TSZIAAzWHSa84r3xxZYh5u9OXtW6YhFjTLRc6nHca7cLnLK6iS2KMt
xynVxMwpC4932JITbr295YDS78cTKpe06GlYNTk7MIRNZ8aYxV3dGzYf/hacyoEQlCTVaGFZc2hV
dsPs8pUrGewypZqPccDhiUTTsPFdNQVorc30EY4UE5+wIMx5nWRfgzPjqXXzLCxUu8E9JczleXus
w8jQzAQgPiKqtteXT23U7h0El2FuXT2ms2DJz5glXkj2NI+4PsSX8MDegB8o1Xxp1Ie1B1FoAkqz
v+KVVcsUFa3Evpp/Tk2bQjn6j9rD0Hq2iIDeGfaj+Wg08kTrx4A9I1hnDhH16zFAjrDYBnE09uAI
tXiDzzBSi0wL/cROnK0gK1cwz+DLVvutClKTAmqzcwWtayvtHKCpq0CYXq9KdFQQ4n3cV4UW4hLo
FBUBmQVRA2qV/oprycvk1LNmPbeT2G00PqAFASY0cQu4q3tGOQrczdhRL4W3wQSGAKFg7EQ5tcq9
8G5uq3jGNSqt8klVtESGjXcNOC6i7WwKmStAnjV4r6JrhZQDlOhSLf4lVrJsYPleVDqPbfIfVM8G
31D0cKF3NIkHChMbkXWfMgDKT2qiwtV4PVYuZ73ejf07mLZTsutuaj4jp7aqS7OZs3XvZR7klR3l
VHfST0tL0njMo6lMBB3dDsGJA1rxoii4TFpfUu5AXUJSd93hR21s15K2kit8BalfcCoVKGWrHEYg
yWQOG0mkqiu/Co63J4U4HubHOBpTGeZJoxR8kyQ5XPstLehNcg71nLNZ0+F//mSHs9KulfNQs12N
HguaRz6pG01J5PkfySoKWSDE2EXYxXSAornNSTZvRBNr04G/D36ss4GNwB4e+9jxPnIW+6KQAsp7
Rtghzl0hdnkjY01C9XBayu3QxltmWgEelzPAgmFxYzi4yJxWVf8+DnApFpAI1E4nGZLXWjJRLdIn
xIZLHvgmUI53LjhVj7rR7ipCdsVvf1W9JJN3i/Ir+hSR+RK8OwuQMoi126A7RoVRAH+mFCz4UWrC
CTNk5MWnE0jyUzBD6q+nUGfyNRZK9MFjMPxITa6f4+0Wti4cahp3E94Q3gX/6+2UcbcqKHX5pdbb
6mikMmW2STNqfu+dUOKfDT8u+zuDXF6b86xMHHH6Begq85nP7ibuXlnIm6OlOwy8Um1oBFNNWylr
cQ/VEGtcWA8VH+vp3RGTUxlWyk95Hv9rzHw+jgSCtuF9rbS7vahqCprQF48snFtANvNqiUvu4iuI
25Ij4Nyj9yV0fHa9D25J7jsdhhu6qErCcB8gmQwc2FpSbdK+/rsZAzGBwyGsBmwHhxDvDuJy3suP
/sTwSCZw84CsxdZvJr/p259eWmD0BAUzNgI+eYYmfxbSxVKNlwszAJAxEKTa6AOMg//yALp5YmdE
6qOXR12VMqI1LrvaxvPGDGL1TeXRk8Xgsi95eovhG1QnPqfjBdiBQs/l5EKAL0dN/4hbGutACSJK
kUK9pMW77Ol6kDYctDMJR36FiFy1Yr1Lyso1VDaYWI26KiaCe6KtAwXOpp9qooQWrvv+qPL2NJHJ
yjYmpFH8hlA+vDNCg/54EQToS9PNwiD0ntnmnDYzTn98Pa9GLgkr9TqAeHQvRCC2cZf5zi8QsfkV
z1AZYfHng/NebAASE/FV+6rLAUeV8z9rODo9Jz5/GKSk2IV/JeHOz+AmgnWweiaQPuomhGNYfErP
aK4uXTIEefBS4o2tN+nvGK9uLXqitgAo1K2B91F5KNivcj1ba4L4otmj4ed7TYqy3ofIwTEHP1tO
uWwzGyGT/Pf01BA20RC8UBj1ILcw949M9dX7T/OuGGyfGOdcmbaBqOqvADJR6a3JcuzU166ieFz8
mDDCZwXp1AOWsmIiYkfrdQMf3kpEeo8i4+4Z/Udk9w1WGzWiHJnV+XCIFBME64ncpyWhqNetJyDM
FTa9JmXvJc7Nrfsnlg+YL8z2i7gytfFZ7vH2FNHzy4+JRzJ7+W6IEdQjZZ+uhs9Z2WLRu6EmnZzU
fKQ+lQDY06QUTvdCYzl0Bh04zKds3mR5AJaVbHLJ762NW2qGMbtuyMUzVbgFl/xMGC6A4QaHqXNO
XgltuF1fH7m+K46bBpty2J0ojIajapaYNpw7eGn5ZgFGzw7aXv/g+Z08ewzMvTFMAkBcvRE+ORFG
14QOg5cQfdi0hZIqNNc7A0enM0Vzl4i4MVzt9tBi0soSX1Ka/BJlq5btbI1DQvW3wwa4hGzdMHil
778U+9MaunO7P0KI8JE9XcNNKcjs+7muDtd8c9+9VXS1VzgRebbwh+fw3BjYGioEVwOTV4gZc2it
x0P2XZXN8kW7n7+nVl4xBedtUuEXESca0EUJohQl12ZkK5DD6Rf13CGwFu5m5PLARo/+Gw2a6Ejy
Zna6B6h+9/im9VrTssLbggmmoFONB9uWjJEMJ+uFKYdGbKYRXh5WHm+Qry5u5xH4M/v8vpS54AFH
KG5THrIgaTfpWaaCiMV8OiEEdjctPVcq/63orXdSqkOGeqE6bbwKwss1yjYw4CQqWUk4NPiRge9A
ZSIXQiho3x9gVTRnn0zBYIyGNrWbHTKyn1hi5xDnvN6ci8iNDCXWqVt0OM+s5407kDnfWQH+O/8a
XlYzUIwh80DU/6+9KIyIIfNknb2+qEeh4AJFB9i7i97k4fanmwcnMbY0NPjGKlzI7u+S2XXQfztw
/0r+dC1pm5eb2UNIGx4FYPRNYFZgAghKHxOKVKcylAoiPnQlWb+UrLbxknDaqOAGTYW8fQHCNzY5
zq4S8IXs+UpoxtwP14DU3xdW/qVcFD4yj2YHOdqM3DGzhhaAJXmXN4E/cpbkbEpyjjoP67RDVMzM
+Sm/7d7LBDzcCCaY4zK7+OpFjoE21V8gaYwhUmzBMnkFeLl5S5Hg3olQba8nxTjudYep2/FxmnEv
qTrzdjBTJamK+JcRYfFz1x6zfq3vWgDcpTXaVHoC5UKTXffmVm+2djvNkMYEm5TEFsmZ/TUax2zN
CIKlHbOno/OoXbuLiZzvdh8RKtkrpXc6bSDb9oJ/exfxMEkHq6SwW9tPcaMWwkmATUeiZlzHz/2f
CAIdmwi+TzFu6YxCR+dvSimc3w5sxWMmBb0q14u95IL23xT8E2Bc2bt0ExCtDUckoTM2w0ZJoUsL
q/97NTvbR/CMS+OGCIcxIjRB9MKdeu4DEtxorGX5n/znnLXbeaKQAW09FhWyvLPWylSCIcLxMOkr
v4u6rTcHvKa3JvqPJ0f7P7mSALuYntFqYFMo4+TirIywHMIy/QK1nEhk/E24KIQQC6Mfu10a690E
hlr+vQMCBj65uaOFnu3pGTQYl6onHeNwAqbHFpIYyc3gHvUpNKk6FFyqv+NOuu3/vZI0D7xbnI6k
Q666R2GLEHAIGRigzBbA98l2IqOe4MwygONP2GUB+UrhKr1W+exY0gAdxAMGR8jsrkkc9DoiJG/t
bsqR4NBaLI91GA7nFPWJOKYZbTXiTrpEZFJ2gwtYc8aLEA3GOHkFw5WQSdbOp4+3kB32PEMqkZ7j
t1dOyhoh+SfpTCZKyu72OVJG2SDU5XqJLBctlkWz6LqUQ+ky532sYPtPr0jVHdesa/5XEEyX7O2m
aWJnch4sfhR6zwHACvkUnPVfp/ZrfVNHgL0cSNGCmOI8tmxpixlVJdPDECNc1t6xFcvoeFmJgFY0
h3Rfy9Hmhhb5PmHP7xupTZsnZ2eQa3cIL2NxBnN2y/VJAkPmk5hrP+aVOJZWW5K9SH0/yf7OZLBC
JgZo6011pstJA4qsYpddWOaK091CgwrWVORV1t2Q++dm/4ntcdRW3d9eaWp2PLZ0KuZCC8Ey6BKZ
DdQCBc5pu+i3+Crf5N3FU94Es9RlVyPyFoKmi+4rez8FlxetnBPoJhPm6JrwCLIWmYey0FcCYvrk
+Z/kXEhh2UR19kKhN36ZXqTLnvjdPUjy8NNTr5//XNtG3bMi96UZ9RjiH4CioDg8NGmwQxTFSe68
p2VC+SPESy3oU7nGYQ6/92Blc+mjoJ0yZf/Odr9V06xUx6bpaLEB8HpbkkhoEDW363FfPzrPFF2e
8RzENuzhrlGXqcKnRFif8ASOri7O0x2v5CKbapNzaqUXZhBEFoOmxfj0hAxDhe21/syMYGb3hJQb
Rz0JDSjCuYmgwjIV1jop/qYi3fC5wBLV1oEWUYUdoAED5Csn4kvhIx1qddcNHA/6T8xkrngSzOSu
7Oj0ykOmsZoRgpdYAzYPgqoQXcnuhtgltwHT/oFQP4HLh9eyDc2U34+8cYfPPMhGcoyPp6HREbyn
wSxsYzOrJqte/qMipdy3AtedMlXUTyCSpRvZulR/5j8mc1qJyG6DyFXY2rCo4sW2O8XI3dUp5UHi
PxuspE0lynMYH5JKuLeuD2RoKSavctS4ZXLXx8v2dnCyCBwB/97hrtauiPh5NKT4Kn2WSgY6aHta
lpqkvJSK3ee5/FBf25cAQmzbPHYgIRE20UBOb+MOmOlG4toUYSCkpZplP+KBRkYF/NSXBMeOW4Qi
174AtlkjiS0lqEI1TkyQLa/zewxtb5P4pgys/vtGz2KKkY5e/aAJqn2bTwHJGnPyo4UnoOV6AvBB
b5IYwtib5z22EY4gnUzEoedkfho2zLd5/x8Vcl+3vKMOxEEXRoKPoDDjyuztHjxGJB5w8mSPDG2B
H0NHPJTWnFdfffjWNC0NPYZaI50qABREUphqbkQLOEACAvy6AHuISV5eexlRhO7Nw4XNHBTp1LXm
HLaQHADcsJaR7BWdF7UvLUFJx7fJGHHAAEfWyB33EoYr060XqM+tzxNBfJHBrfHbFR7slmFexqDT
ESDJr8vJNZ6YEqlJyVdfzmrTgEo7IG7O5hNCuYN1JVw2tNPH7iBWSVuKKJF/puUDSs/uDZIka0S8
qm1ocEgVbzus4fcW1qyzXKyBXCRWaW5MgMs5sOK0pUvYebBf8ZUD7gTJsTSDAbCzHc9LksR/4JOX
G5IxG5jKH1jiFGi8sE9CNBlM5/zyRZDM3VUCNapLXrHQuPTfY5ykqat2/Trp3lt+TZLoa7pjPuCE
ztOb4HgszMVjad5bPB9o9selhN64m6M2mf9tyy2dosy4L1t4wcTjIvfuHrQNda4pPnaB6HsBB3AW
smKkgDc42fXG8cXp27Ry6vpSrvc03wssRpie2XMCmkj8dnkiYqKIJx/5PmL7HR8tuUsuBIcWYwS9
6VyHvmLBDV9Sj/vKBlCt+/RtQBaKQwnlrlml7l0HosXplcaKevWfhjrh8Ba/2EEvsWV+gfK2kH92
V+b0we0QHKrsY2vPUDE6SZ/PWfsoUCCOXN7fIkeUEUNz4VssVWi+/vXzrkAScN0xYCg/acC/DSjy
QbuFyex92YAhHrOv9bXsnsWiH06YEux/mKhkKeqNaORHQQE1yyZBME05I3UMxVLfN1Byl68yC0Z4
rRzXz9Xj9wQ8M8SwkvFpoPGcHycYOOrcGAHqIBFYnEiQvtM+uipQ0VcfCEeEpoFXsmLaeTpK1duS
Qne93i/ipj3O0tYgoVTFSHuIPfaQPuMgeo+Iytu/RudlUcYbJJPHziREzqzdJT1Lh0gvRrmUIb3q
n+5n9HmDMH9V6adJ+PNUH/GB8QQOYQ7HlJWw0Utsmerrka056Bjcd1RPv0AEfhysZehi6J/3WNdK
pW1a5rBPU9BpQZDcbtD5tc29AQRBWxLR4gjE0K065XDsnu8GagUJVNvO/fWWw8ly6kTq6ZGXE7wM
bTwFGAWwojVDCyIProrYoJLHLTSXI7OmhMzJsgdUt8TNysiIrtsZiHAaVRfFzGSifrEIJHfyRM8p
Vd9R/OmreWGiTMumuK+xM1jnb6pYBQ7LrUhK/QiFr36GuU5MH6ocgugo8O6RcK+yRFdsOQPizDoM
fTCb/wpSoKfDySfoXmZ3mkkR6LaoQ0a8m7bUUf7dIFdxnC2WdZAyW70N7mHS2CG5hnZuR2xWzSJV
DTus1XVRWYnZ0uWXLwCJBbyYIJ4GeICZx6CXL9jxM9nDROVC8Wrzjj7WuVTf6Kp7iR7ZbqPnJ+rU
M0ZT3FNIZqypzEtiktZ3ErUUqeNGegY/L/w5yItZJtCUGhic7Ncfp+51rjbnQ5mbQcDPsaef8sdH
qYtb167ewWcuXKAOHO8cxU/xYMZV61gMBu2LGSCVtn+Z0LAZ25zV8fkdvkYJgq6BoJPnRLeJ70Pr
XMeZPmOrCGahYBvnM+zSU2bnpK9gkleF9DBvmS2lvznqr1UKBM51aa5MKAe789y3scS0m0cLEqzO
3N1aF+MAzCV3UyhVKskpVTc7D7N5Mu4MvcoyfDDe5BevbWLtCIoMX9tGDGhmMjVh7tVzE7zCMNUo
IVkp/QpPmH0Krwqz1Fl4MO8Q5evimFHWpm0dqwI8+qz07AiTsLG2FYnl1/ITVF6vFfl5UuP3SpLW
74ormkIs+bX/XvC8oXDIttZYV0/CvhNqAY2efX6sNyIGwgL6KsCtNGCBNNB5sqXitjPOw9YHIJi/
PKAsP4RQNIfPJ8kpMQOPXcfqbf4rfILFQFQwWhVqj9Hfm+o3MINzn4CNPk5sXd9AGZADosBqnzCw
dStfBjHxXE/SM+EtTN2YHZrg78VCFI+p65EztPbggIZQ/gsyCplawaSvgLPJxrRvjc+uHcgLTvZF
nMgB530w5aSdgDRGFZR0cdYAB4ndn0cm2yW9FAQCS+CkxqbkfkD8wQ4dkXz2ZPQPMQc2FEHZ8Yhn
doO8gq6pBsr5TvoWDQsomNrJMCsdKtAz2KRIhNpcoXntFmosCN0DUHNC2vzErhI0NBGJns7BFCEL
3iyzZLukCBEQn6wrrOI3SCWhogra4tTYeS7v733r4mT8XavsZBRBlBhgxQMeAnbJ58GGe8wm9bEv
bnIqeNzZbdRSUHtnf4DNQNruw+1GoFWVqODDhHSKBusWyYRp24YCPJpAraBEmLTDXvnpoUf2U5+y
CbSHkb6iKGjfNGmkiX1SpJA3E9P0BIql14HOg5WIZkm15BKZt8QxybNlkqbkh5QZUsJeWFA3BgMK
SsiIkDcrYtnLuRF0adA0taZQ3oHpSAcZN0fwt2s3PKKv10L8GjSyFT8Hx5+/5DOxGuWQ9MNJ9Ypf
ViCOZTuRckJm5X6lJEJRR2z2r8uMPaDydqGGF+FmILXkOafX2Blpvp0vsOdRD8CjR1lLeQZX3Um+
i/Rh0WupqdbxFc4xvXZz+KS1OumOpsauaqAdHWzXwOg7hWKwPPsW9xMeK5juSMDQSFOVt2bEthGH
+sIF9LEUe+5QaoTFjEj+cWhShoKewt96dNsyITAJWempuUWrorGc04qxhb92uZBsgRUY9e2GU6gZ
bn1TczLMDPGZEShbpUzrWmbQTp5OsvYIY+EWf9ytKdGP/jzL3FfVCC1IvRu4Tep4FqKEpFiqpfHz
zq6n/KdzfGZ2r+7u72XaGiyIZy2pAqcqgojfORzTjIYFDK1c+qv8ptEAGMskMd5KHgf1G4j2wlvZ
eri9P82Heqw0c8JQ/TqXUEEFC2ZIcVQIIWNcjovQ2fX/AKV4MAqZbuRTgdK/IvlZQKjP4dPf8zsH
vsqKZeTZvL+SEjJfrJm+RXDmRbshIsUZwHT4RIrtIaBs3KpsI4Vmh0DE5i1bVnVs6wuuAomKMHmZ
t60WUeNEH9Kxh0IFZpfSP9HRipWz2GHmzq09im38eUty1rPJCelZjOra5A3X1wFeQD/d4ME3NfLn
6J1O8FktacsT6KNQGMQZrIwwntFjEncv+0zUf2u31nihOhvj2XaZjYcVAWud0/y17fx0mUE1VEAg
O9ySPZAnP0PGcQgrj9SnIFfchwt9mOQD3TX/1pTzZyDY03a7o1H1+Km5yJfm0LaSUVXzPfF4Mz0l
9yz/5d+b1k56DoSXHgNqABdN9bIhlaWiu3qGuTR3F4zcfmkuqqTQNC4ZdKk5uKsMlUuDRfxgsw9b
oerRoe2MSkHQv26Mrz0xNlEf25+PtuqHXisj1hZe6yVKFAh1wLN6aQwP9ZlnK+8OQpirhx2Phovz
xRAe2kLFE6750ysr0vqVY2xnDvkpnR3Nu+33Mh6KcRqSyhFZt7WJCy44cdbmXiyE3x1o05kvT7j7
8JbbTPoeoaAFrtStmmbsO2NmzGDBQTnlt6V5xx5NMcYXawyJuZWeivDnMdLYUEkrth/nDiX3B0Ey
ccD7vkESBLS2K0drrt3VZONxnQHD/B+MxQz6IhV8BsfUN+u5ZkeAFiby9TcHyRJYTIcvjzG1yMju
VPWJbVC+vYo/L0YJAjw/JLE4sitEJ4NB7KRuDpxveYmUD3wRylT1LTLZnWgd/6dTr1sBvsLKj6Gb
zYjk+Shv7yQysnhh6h4zQyO+9tMRwJinXg8yPZBwOZt8x12QGPG0BQLfXQewLiNPCfBniG+XcyAd
WqUuyKaOIEQYzL7PBW0doOGBd6eeTVN5MmYhs29bMPiTLWeu9uEx8w8TDVvV3/meCqz9/Qg1LD4T
xXY4hdDEOXolEHJvUe9c9stqQmd8XDTiZ00h8EzddAvQHipXadiY3YIs6Gf6fWrNGyMJV5UopeXT
Upu9N1SeaAj4etqtJp0KLzis+sgcc92h4SMVzvK1qODFe7B4JS0KBJcWkRYvQ29y1ZA7GiH4Yr4h
ZhxHlSVA7/AQNMKi+sX8GP0D4D+TsM9qPyUbpUfR9NRcq7W9sNmSNuhYIeTgXbXLqnhEOnkSPUI7
M+6pzg6tjrdd6RaWUUZMfouVXJtOebrhLs41skUhG2mfdfubkpcUpZ913Q+zoptGFQZjxrLe4TT2
KDk9OdSrz1IZow5jVsuUdYwlN7C3MbnMJzZFw+5EwxrMxhWo3vLM3dYIwykZHct5LDbzNoJO48fn
D8XfykXq8vTSngrIfA2MFLeB3lcR5GbHnuhTeuHsBpRBzyIuehSHK7Gs2fVhWmvFGvjIulnQ3Uf0
kqXyk4uVpqBWz9qUOMGpOunV+jaT/QJjSlUc7jKtEP6IeYHlVBYa2OtTEY4FXxSA/LpEg2WPqBKo
1IqC/vsyDCYlzCaBr8snj4A94246z2OTeGcpFm/uyIAgoKeFawYsabmLmQdt7f4mhwSqArODAx8V
mh/JxLSkr2xTCASPUdaRrX6O3CdyAH/Z1Qrhxretl+QT8Gwomu5CQyOG/1D93nqOEH7RQdnbwcg+
KHH5MBVKPoRoCkwB+6KWe85h1nbIeaA5palP1BzTBDi2aplkQA1N1Sp/6xKSONtKvffYdhfQDUyo
URl6darm8KGWFJLhSY4+JMkEVH19wbaywZLd7hztfwnYFhTn0vW9su3NP3bEhTsQIpeRnV2tGURk
ywIWz+6QVkKy4g/dxUEjseOMTGcMArsNc/IS9K+Xs/obGJAYgpSOlpIz+IpKY+WakWBGge9lJcDD
g0c77MTrIFZI6MOEOqbUdHu6TM7ocooho+0sjBsYF1JsyCRtD7MiCMjjysUHJMKnZPlUYineY3VQ
fPeQBOKWjtNePCaHjKyhdCnEY99DWUjqdoRhOnuzRPZQxqYPD9FMf1A4adIvhK5+6CZKNr/h02zp
36vhjp0AXnata7VTPhK/anbuQdGH7kaJf8sdUQ5FcIx3M/A1Dq/qy3D3T1N7KYpePbhLYy/ryZOa
+NMjbUc46QHMTWGj3IMIhtimuD+xNWdrQmGCNKVfCVstOhb6eWI7Sxd/AGQNrajR89p8EG6vI6IC
o9r3F1N0ASCtdRkliyyIYLx2nwGSacxJBZ57x+UGI7SjZOUe7WhOe6ShOd7bDHcEsjUXYOVKHtME
HyxQaouzmR7TpzNXW+rmzWQ4WtTTSEGvqUlP6luKTI0S5s91ajQ3kApgnwZGwLS3w/xk/nI458L0
RmvuUR0oUUl98RhLKeHSXB04VbllDsXoO5A2Q3qDLtindFRQ0pPXBgXNt/foTUWq72wNH7DVRXnL
P3h/DcHz1FQmTbgCUJt4PJW+0H6O0A4TXGUaac1gU2uNWI98a1/AafrEaZX6lzYt19ZXiSKnNdpj
24KPY2zDZffqJjWV+dSM/BI8zf66JJgqp52ksVaq2MMfpnc5TRjMtWVpcGQMw2KUf3jhFA6ugbo9
S/50Z53ojaOwp1fxdvPVHi65uVbXYi7C9JcZ/zB09wd1x/zKGP7qqxjGBlAS1nzt1MTsnZwFS4I4
cB4tQgR2xkozvym/KZ5197B8aCfZ3CVU+sW0nDDHbHga1bWKYAFjFqGxMeLM+u7CThQPY6CpIktM
kPzpzH9VW7ngGpkkNyfBVU2ba5VIAhoAWkJWM/a5NrVfaOE58tKE46HUolJjoCYdMxS3ASARkjBg
QR570kxnrVWVrnw51uPsUg0BLdb7bPR1QkYbZiQ6onOQOfme+3kmEbig26RP20V069GqUIGqcBRa
1aTYM10BnwM7vOn13sNzVkuaNNY5Vj4Jfr2xyu23NxWHdToaqCPDA0YpUWmpJRQV1CXtTUIeuf1U
w7d/6yMY0gmBtK/rx3crJwKo+N87fEwgPvsryL3EwcqFdTMgqN+bE4RQijYOOrcdF09RUXnS8xll
voy8/DlqGzmti+8Fja7ac08VNp14x+6xH82mg5ZqfVqoN4wX5BfWNwpAZ5oRCS1DgxVB8QiOXMwe
93/+psyelKTfgyeOC2w+xok/Ju/K3rnlkbYKX3sLBDPlpG/u4JBvZalYQ1AXVAlsI+8To/xVMWvV
beK4nDRDQKkzLPspFc4jwlMV3Hkg5LAkVWjc1i4icEC+zdl1KJ4/4ydu8BSbCTNxxSIwYhELLssa
2Dw+FOW30c7OQJTRscP63KnZDiYiblxFOFwgoTim0+Up04xGf5lc+QBZQc+lfOvTMxQNhsY+4aix
yA2b1yT39ZYjcUcJSX74CaAf29PEM1l98jB5CDlFCKbezEuYMk5jGj47Yfd076+JWqS82s/eU3q8
J05dfqQwwKZPQqMiSp6cDgjI/RX9+JUdyBnSfNpjQcfKv325fXZFAjHTtZHrP0z+7U3JazsZt9ws
TG8T7jwZjOdBdEY6XBckVjLQaDgXWs+o78zxs/ZAGJGAGqXS9rv+/Plndgr+ksr7xrJ/C72wOP7l
HtoWreAuBo6XpqEI92Rlg6FB1a79WH76Tt5sIwEtsMK+jSKMx5g9/+GHH+ThRNeDSt1QTalUuYyV
hxu9fLLRXO/UCi1wwLE5tV+T1hX8BEzEUEBEEIJTFdJXuY9AYEsDAYCxQj7NQaEE5lkg2YrpNh+H
77ew8AoonXwQKhgdHcKEUSzkBuNHTzSpApJhu9RPMM7r72UuL6y3lZDWqNjj01g8fE30mnO0ae8c
1YOJ/jIIuYDzEzCXlm8mkTpAVBoZOLlwq2w3E9rZrX9q3MgR+i/Xhonez1yz9MvFtpqQVHtR8mUm
PofjkFCeKhF4+0U7DYR5zyMn4NWsehhxsVCD3Iy0nlS4sp6qRRka5fzacIhyciD6ARfMO7/+HIRi
9+XmSwQpDlR016Gggu97YOpYbWjJdlx9OLIIaUS9ooDUNgzkLJtTkL/RFt3eW+IChfHgCvJfaZCu
3QRqZ7DxrRtlBeybpQuzDLmFxjWYNH0SA6i1eebe3dMaCdrGf7kpHJIkuT+xGh22Y8cBiiDHW9gx
iOEl30Rng6LOXp1Q9E6rIudSf0rJ/koucm5+GKT44P+/OzB+py5BV7CrQm8vtf6l1i4Y+dyuYYTW
BLgH8lKydTC9q40VTDe2N7B2pd/vc52kKl5brM/haKWem70zzqrtJb3D515TMjH7k1YQdNYqll1Z
5sdAWHDmoh7KRZZw7qjuHO+vtByqs8B9N3OnMF7uSnDoWmo1t9xfdmvaQBRpye9FJ9qz/auHhUpp
raUWv7x1OZgrkE6/s6INnrsyqKSHv1xFQGp2XnbNNcmuYCjOEj06c1/rzIBy+fnjJbMN9PREQ5kr
LeQuemJCgUubIbzHwXdA8j/CkJSvTYxSht/UzwRTeH/vc6EUu9mlF/3o/ElDipnJLk7jVmDYWy49
i2vREwine/yueTeAQyd9aMjIiblZzzWK7DG6pOrIptYSe27Q2fbDLmO+fSRfJezMXHLo30ebEOEw
6hNsJNhSw1RhzpWQH3j9hzl1v1+31QePnofyzMtjSyXJRZ78HPctGsjyOo7m28oYSS6KzZZhamSl
TX/4QkI16ocqoVEvTDvWtS+cwLz0TRIup2YRCRbNEbwqOKHo7BmLYGtDGpIHKMgicMcvRXQPQnGX
CF8RU84aYOJOT44hV4URmnrGofnYCTyda6mbX90cG6AkSLgHPRGhPRVC0hLyTPKX8ytCNF3JYryO
XNG8mkTbtxa/YsI4KuOxGdmL/byCaZcP3uKOlRHtbqVu9P3SlL/zWkrUVEih+A3NqLqjy533bcCC
/abhhOklfOwzSMJotKWyh7jIOHQifBO0/4Dp+HUpXy26Iasjl4yK1XEyvbOtW5xzViRNgDxyZ9yZ
/z/CO32thnzhIBVZOZHPy/as4fJa0X04uu5d63QCeq//QVIRzNyXXXplG8EiUPJzVAaG18nVU9Kw
4HVR72ahcjh6bDTQSyFdgusqy1VEtc8Jrcp8UKTRObjJwtjHAnKzhYEL8nieubRdSMXV2yPSbxlA
hJR3iL8fV5mLTZIS8yo1R/IuyBSTu0ozVBTF+h9qX/Jx2jduVvuvrY96KCtw4CPWfPi/+GiXWqL1
BkxdwGy3Dcph+XQ0sS1CD8J0oA6wIRb5SztCtb6MDsxqxh21ZDQIEC+IJ6bhNkn5u/qwNFq26v94
gnJ/K1l2FcDAHSsIy9OULlcxnK+r0i+RBujC0P73CuQbwvz9e3w/trnErjkfO5LDswl49p8xO4/A
dNGDgiy4vgm6S6ZqTQGiihbJH0NPXAEBFY/KnfDKJVbwANLB+rJc2WfKJ0BB+9Z+SKES0cmmWBjr
elf9ZgeBQkUZ4BPD+KceoWPwiN/3XopGHcCL3+kqh1aWXBkFhkMJH4Guw+sRkv74cGBtJEw/4KJs
4lAcZUvrqZXrU1DkTdIPljCDO8L4vZ7Jnk/zAb7N44WfKpgdAN1OVU+lTZ3S13RI3XUhIsUrhb7S
v9qVrv2s6bc3L3brzuLa9WOgEYEMvj1vN9g9r+r1AR7trWhglXvEr+1moRxfq2rSUadeAZ8nEU5e
nh68lCLa22M/To0TLErNrs7YWTglxEOh7eiulTVUpycNHBdyzQMXudnpCjm9gapObFyxeCIsEtfo
suN+3EljGZzTVzg6czMKAowYrcDg2YgzHGBKPQ8F3zJOxE/N5adibysDSUHAWBvuO5bzWrDxMOy0
ACpyNiyc4VHtcuBZwiUaCcTJL9m69lRkRdAVpXFw3RDsgPTglH+q2Hm2hzrZhfjxdFPXR3ehbQQG
XWFTsm7F1Unya1T71+jFUg2ASVeUebm/56zXSVKvDXid6EsobNEnry5XImW3TBLGTvZnO4IowBeB
6Uq6pMitRWjXCTB3lt2SqHA7xK0Mp9+5yYDacFAUV4+AU2LZ+cBWIR65w4H/VrKBJ4Wp8beVU4Pv
SB0j8SyXWZu6yFWv8CATPfMHMAk86Jk7szClCYZPgc5Rm355knF+JJ1bteeT5Y2DfukxspSq9fZS
2iS9uOT0nw64NYrPhn+bIUSFAa1RuqOoJHT64EJ2xtGHuqiXioVo0A0Xc3xEpVLp3/jMrGHZ0tWv
4BTaUxQEFo7QGxzZKZi2CzfauMLq4tU8b85AwPh7quj8qmVk6kNXGRZXO/IQ/GEqv/imRrhbcthD
+rPSEkxvVIAfIwzC1mCMmMP1oJ5p/evmP9EWkCGrZwkPLnqB8iIxll1++xMjIJihSui4ikK2d/XO
LmQCc+AhlGsaWsCt5eEArlckzMq9NAbwedDxOE1w2KB624OHPFz4bUvLYYE3RJNVNujIiOziMIWG
VBOSa3ZOZtxnfYJKsQvwVcoPUhx+Z0bJ6LL9MhYUcXYgZ70JAkRrRfFdDFBMkxzAZ4SYHFEB7hIi
wcmZ1fyvOaHrfq6bsYZ8PD03i7uhgiYT8LaBh6+egGNkS68BSQ/LUqoGfvkkHtRvjZRPrafInKCI
R3Ixwuob5SzF9TSdK3P8AiSgYOwc8tz0kVPbFDmXw2oMy5PsiQTz87XGzooE8UJ/RkPmXB6jr+iN
gnkjYEJoSg4FTl5eysp/mmqHX1vb3rKIEu0C5c3eF8xWV8Eq/GASQeqsyb8TP2zZkjNJB3h2+8w+
SwKjfeDel67HuzuwJmhgjgqTfoVcqzDUuh5KRRXwQv/9uJG12kFtWQWZ9Mx8Qmf7qbSUq40TBEuo
z+z0SWy5iQDzCypgiSYkhJDYMzysheNw6/07XttrOj2tBq7eBZANUfsPFUFvshoDTEgsTDmKa91G
IVhiLDu8rRQIQ+PdgJmLDMyUu2SZWUeds3I2a7nGQOYvDErlgDKNRrrUk7VDGnHAw9u1gLG1OtXU
c0ZHDc8Aiu+RbKLfzXHFpolnmHSLVqgaBQirjFcKBZuDK9o50KFYV+XG0cthPSpbtkCmHBgomzx1
Sn9vTMBu25dikEAZcFz12PvcFRJOWpEu0+5/RqoIkvAp72GiJj6NFH3jBFHuLomGph4KFskdXt5Q
eyueR97OuPEdI98Q4vdhMCqFVjla9auJfzHop7ihRtLh8acj9BSF3T6OVvoR2sACcQZ/MJ7Fge8M
eiyWuUc+Gyj5pu77w2nC0DSkGkrTJxPoQPBZpy/tqiI2mCE8Ux6vl2DQGicrBYJo4IBI+h04EEAS
K1xbvKV11kny7zjjqMxtTTJieMqz4xIwdbKiwQzaLb4LS+JnS5DEv36XUMPP+meV9IjMePGtboOJ
yF7sXU5Heq4xQzzMxzpwjpAr8KE+IVFM7lF/jnN81keq03c5E2YSuOkgAk60kTVlphHO5TkG+fu3
e6RKhZNZ6ODlf3F9ehGkWT8xbd94cJRxXEPCn/WqXva7brr7x+axAz/KxorQne5bMk5jRa3+1CnN
JWwtP9rZLD/1MA8ukkvhT17gHxmCuGk5v2L57k6nA+PM6bp/bnBwrMoUyNUYSNMw8PMK51HtF/nH
vp2c1+P5nUv4zcDDA4syVzWE8/jEfqjom+dmJmCruO+6Ng+TV594aIvnm+Cbj9tUdIDWN1xCXTJG
uD1GlJgtCqIN+JAvNYXlGVVixRgb2fer3AzoHlVbpkE6i1sbT24zPXUgGXXrK6Yd2rh0BLsALas9
87MNoxsaZKT4ZIbBk9CiHLe60k5J0IX6oo7LSMGrDrQMhWoz3+3Gr/0m/JLd8Ldp8NPl1kmJFsR9
F9ssU0oxgREaNLaS6q8+iv8lJSXKPfLRlXJO8Rr3MhrJbe0C2tfGw5WwGSJn0CD+VaApBT3DFW7W
t8bt329RCDNFmjYSjMoe3CMuxbde885+KraaQHYy9mQ0AordeTsQUorpfGrDiotk9zoue9b+n+vj
CycQflMq2pZu3LSO1lMIGrka28/2sQojtPA1usPboodtODnoZ02CCvP9PT7rghSFUy/XusNwD8l8
gn20KYl9t8v/sOiPypIHbn9EvdBQZdMZWxpTxUvxhTYLjnWFsSR6YSnBkehiolw7UjUHmfzfhz1a
jMIr4oHc7Ex8xXiKuDcTboeI3JZkeuLl+vqPEhHodZdJ4gYoq5dw3Fa5rEbsdHA07r38y1nF3znr
oIUYNYj39hpMvcBVPtB2k1bOFFnbTHKTibW15SoACEy00/BmBtiyrV2e/b71qidlb3Z3jL9Ts//7
GRnlSYs81nIx5mRwLZUoKHFOVTDjLswiwACgky9rXhAG7vZIHFquKaJJtrNwtY7S45bRu8cbf8J3
0yw9e6UYlbUBTD/nF3a9a3d9dujaHizeq2VBBVMRs8WF2KNTkwXJ0LnRvi9l7pYx28Pg0KSv25Ef
zcKBLT2w+pmeAueyVJrAJ0Hb+GafEEv/4WkN9Xwna1wlmxzJZfV8mFT1HKu+VvC3x2Or/1w8qGAt
lfaiz7lqdlUvDzQ0e+BERW+gM2kBYj51MZfOQbdsZwsO2a3mRnPZVdHq63dfd1T0zoWqENy0LiWM
wK3RjtBTpBvTmnCJcHHUxG2lP5O3y2cYwPfTGsemQXk/Ew5Ib1TIol6GjubNgwnwo0UHCBg/UM5M
NsccGcl2lSlbdSgjr+9p83dOHzJJ9RCisgEqt3f442ZuiV6ThJNpiRtQZeCS5COWNVL9mGoUOME8
/q8Dlr9snhOvP+QcnmdDL7dacdPeSGTjJqXFdt4kswXKjPFLK8roofPDOmLnLUmNdCQbUX0xxKJJ
VgjJlIsn7JOGHjRMdVCrz1l9qecZ+a7JsbHWcqsaHl6E6W2tjjxFgR8zEErwITHjSQwSSFQsjFNX
phOo8qF1KWzOinFqp+Beq7lLbJ3IAsX9Aay+eif2rUGPkXU8JX5FxeTTvLqs1sGBIXY2g5q4oToi
ihPY6snEkI8JyQOIqRDiKeSIv6iS5AabcbLaCDl0kEh7GaJrYRUZcPr7+rQ5JX9FVjayy825CI0s
LWVmx+mUYeG8xF+1IYadlVWjvztwe6D1EO74/Dcem2aSWN92dmyPA7A0s2s//2FIwkFwxtRkXz1D
fPcH3EM3czJRECrFoVySfYhIpv6iDKB0fBnZeMvaMyGuZxVDIUWtY0PyGzjdrQogSyDPaNE0Jee/
KMVuAXNkVsgQ1LzSZudOsvXjCAx8dKiO232hSXDGCMSSMSuiW+YERq9afudjkKAJ7ox6m7kwrPen
P2mKR3r/jz6mxMqmTBvJwRnW/16hgFeDqk1IEmBd0aeacDAlPi3IIZia98twWiOM+ULN3vgXBeOw
D9OI2QPZL4CDm6eoF3rkj4Tu4i17HkaUhIl4O8gwbKGqfmWxStbTsXH/1hS8cis20u5UrSV6Frxp
QcGK9+KDrhLd+iTZIQJEAE3jvLiGEEKSjANoVZifVV5D2t5OLc+rRNQUW42HKK8Uk4O+KznhPcCa
P/fyAYsYWLG18ewohxdoH5dQKzbpqsIn0Oe8NOO0A4RekpJxawkshwEynY/HMvIfWYMJloYuz/3S
9n4WzHdmTOP+jYF5rkb8ignFal+DV6PwpRdQkfSF/s5vqHPZ3AZSE43wn4C+XozzllkwA/E/7It5
YJrBG0nkEnj7ihRIlysf0TCLRgKk6sQkL34SfvkTZvgoR1N+LXn2YbDm/xjPvnXwbcRN4b5Mc+XP
xXvRKvJuAjFSwAcMZAq8fSV6rCLSCE346bpvNBr1qvVG834VHIyBfjQCXqPjQTCo7x8C94DBMFw2
lJYjMHapVsvoxF1puWH4hnu1uRrQMHw7iu6gQX9cBbzcVsKYzxOtwcsdVOUPCmNPhvlcH3nbmkro
C88lXmNxNd35AqwC+4jVHTDvlVYvPzLHQvnDuqjN1I6vT+O0s1iGb0iamnPVsJgKvnU5J+u5CTcs
FjnArIUAFOtMG2ywJgnmvUtNgQ5hH95y3zWtsQNOmnufqGTAcKpvrthmzJ8eve261P+85WqJ235j
4SfqepOMkuUTZ/drpzDw3ZP4WcoM58U3d9vc4MbTt6BBGqagp/HR8G+sgmQRVHDlE6avPXz6jpkt
7CxatzknZii+X7jwkFBCZE7yPWfEcJkPGCsJyPUqnBzYYHo0w/m8b8wRGnFiE5AocH3kIHB8N8TT
JGppbKT8EwRTkG1cKNzT2vNJKFtqlZo59FdyTYNHIvyonGuL031C14A4Czjg9bH2qA/gnIwDD/nV
MT6m1m+Sb8P3U8LIpzRS0gkiJSdj4V/wQSA/JZhDKUtTp4GRV3C2528yMuwlDVgeIbr/C0bmPlYQ
McO2CiL7YGiRJq2belwJKHCe1nVluTVEgGNfpvUYFi3e3KHiZDgeLbcwGveVOBamr5uQBVFoBaDb
CfPeDPdWU47KKMfV1Qprhg/s750zRzIVmASU7rsOh4fZyEfVICz8mBjzCvIfsxUaI+hVe1BsJYPs
Youzp8msJCXXspJoo4RfPqIt8nCgnSQZzLitOCoIGHJwLJnuDvotoR6SWbqcbw/p51pS4beeL4lN
yk8FUtR4cokMBO3ih4zTLIhmeDxM/Fjvmu8lS+r+WuafFYBLdGDzYTkMjlPJLWZmy4UAJ6R3hs7y
uvVV8XcEabEHYIiqp2sT7zS+LENfOJZroIQg51Q3NSapX+o5dAQtFUgCFlCwSMFX3amHeaBWXtxE
R9Y3lP0nwXf1kWMsOuNSRjo2sa5Na+PHYpToCuWUogGH0wOMoOeEXljENdKU0qlr9nygKFgGwow8
+paMQ2/bf3bsnUBn8ZDAfrVUc/Y9ArQfI0N3TTmRWn8iWkU4j/+2IM69ZLZKdvaHLKnTnkWOyShx
KJVKu2SF23izbZcbXmZypKORwSrZWRg6NJc23dFeP9lT9kgG4yw24yZA2FP1CH1vbV0o0PIUeFA0
AaUCw4t6cWyPuuPPY9bnhj4DX64TSmjWdWT6+U1slm4P9oj5RA/4HbJ3+8L8HUW46z2q0bcQS4Ng
hiBSgP3OF8O+VIjkaEqP+5klqKjCy3vIB27mBBxlpXb3cxk4owQRtdFQSaKLSL+Obvej7xhl0vzJ
Th0dG/6O+lDMdzVuZwH8zywa2CmuSv/G9vkLlUZeFttOuYO2HcKgkI9dOIrtdKKFvrjgWoCdMUQa
i5NfjRE+v5f4VtT4OfbsZKm6neNlDbyRUW1/P98+OXqmLaMZ5z442Lad1zhgJz27HnjoaWttZwiY
t9UNJcUaX3vIwooinMPiOLaTR7y/wqGwMFMP01avOD0S/YKjJgQQkDxwC81+yqAI4FJ8hs59x2W8
QKeoqbarvNIaVJcITgUz8nHtdkreJfRkGn7UCLBgBiHCwP7c7jvrU/rVEoQQ0PEO4jH2Uqagpa7d
nZKgxP6M5FT6/liK/p85ZUS4HEdUXP1YgCxyXzkvQrNedg2ph3OLm5+7LQfUYgWLLyzfuNYz8LUw
C5rvdqW+NegPD7AmhrFG81ozNHcUrH8p2XMBJA3+AawTvsrzJdPH8eCjvwbC4LA5XRNXBT3xo+JZ
5sM8f/vz2HJf1t44DGDEouNMXV4eqsRACuIb4xQHc1QB5GlnU0lzxT39D9YQJ82RaFmU1x6m3b/T
UBxXEcYrbVNg6SuFWlyuZYC37x9LdIUUL37LBH+YL1A1AMhpK8MbjEPT6fBT2p3jHYSKU22hLnbt
eX1/qiHXe4sSWjBmAleKr/IBAEvBW2IQWoSJ+D0bQ+zKkS8uYrflKQPyFiYKCoroCI3EPqBGtXcd
x0EA5iiizHQuRSNLNvY/CrxAlXiG1nvb0vvjxEGVWYWOPoYGu/efNgzr3+RAuP2EbBiWC+6GKq4P
4flMiFkn6htfXJ2wMrQgBCapxvEzoFmkmIyQCl8CVjC3wuiyOX8jXUGiW4ZioEunzkjDZrwhCl+a
exp7XObvmfcnR2skHltgE/TfM5lrAfFhSQbIckc4jIuYjN3cie7LUT4OJ95ebbaOMVh9N0aYPJps
NX977omhB0m4OGx9ig3fqYLDNa5NsaQXrHLNkqq77yPZaEVOYcgrNmzTE/h7uEZBs4gx/dZauJjf
hq9sNomWe7tFgGDXbrRQZrSLXmzE+XAOTOpCJRmdEc2f89vU0oQnVRGZ88PU3FiMmehwMrjTABH3
1mOwEONFkah8FAuKaTmcLgVZzA17EQM3alP7/QKC/jmfwk5EZZlaQMawxJrFZDgpKPLHCMmc7D31
t9aP/NnB5PalJIzcrrN4pEnmFLAHFjRSgAhwh7vckqDU41PUqLqEWXQ9TGWTzf6qo8Smg8XlgcDc
HKIPSR2Df6trzeXTiW2LNa0Sht/1QuYk+ZYGA21tha+5FMe15hvKhKWQEuUxZKPWB4jfGgwboeSL
0Ec/O3yQHeJ+uj7QMJb8IfHXUpdSLTFVUI4V6wNaMST/XssrHgveQhKBnBVXMb3A1HC6Vq8UtH07
fQe2USZ7Sbuj/SEymWwUKmgz8E/YlhqbnrnCrSFggjyQU33TeTIbwhEDC5n+98cLbVvb4Vd4rd+J
Rlb+KV8dklu81TSE1I8xXHfaaX+4SCAHWKQDrcL1M7Tt00xXqhK86kX8kC0eK8pouQMseCKoUl4P
ShdlwCMro5ZIMkfxYL7z0kReUhgjcr6ysZqKx+PHwaZyB5oj8bSYE9OirxYtZlZqooPxjnTWiKct
HYBsVT8hVCSeE3ousIOQrJLB6pqLltjolhsauExSOx+iJBH26Rwi5oTGCWRCMub3dWa4tXw7NKbY
Cp1SQn5Q3xEjwNVwCQ/gU65l/ZgVXEQwDaFmQ/xqDW5RIIGo6nNpwanXJUdhmZ9gc+SGsCN1GLrh
bScEvCc1mNXNAF6RR21reXaByqfudgaKNxPFoue3wnSueoMuRLH7YJJsqw3/qwzrsQt+sDh9acMH
oXzKe/zmFCp4G2dldkQEJw/3W0VVsvlwW5wIXMd6K1pBkZ0erbwYmzbuzD/htdv5B0Sz3ebpl+GC
lxnSiiGgwoi+frzNnn9kbI6NWSF+cuYi4uHZUkTfqKLqUysZmM4ru74tNTIwDlA7SxagpA+Ka/aK
APaFh1OBijzZFu+P1CjIwcOj8gquEYF6oQ7bZS/0RgGdkfaojw8/XxMtsp65JHI9Yc7F087ayF6q
uQyaU+etmkV2pPlfTKDzcTCYKlljILaKuW4qg9b2SQgTf4lZIQaANJ5skv/QjwVqSHsGocdkB8w3
GxLMyZYpVSl/GjcyByLgH/LIOqA92CKjmL0BCEl3ryfnPor8Ru5IN/kXhyfhLidtlERcs0l12MvP
glQetOT501U/Qm6JXakfJKPqL1+pGuxqqCY5dZVD+NBVZXF75ex5LkXDIEPWmolrnLbSXXz3Uj+d
53jkouOTHPYKMtxwX5jb3HDJQvB6p5ILQtwFuW7rqtec65mI1j4sIHy5BMCnFnPmSEt1CXBoERh1
coCNQPB1VVbh+zEBoEkChnAbcDK9as0KNPCNOGDoSTY5zKcUdiu/tbsoOp8gMfyQvjGBtO3itlTJ
OO6se/gEJolXbrf9BBzfAXaNpkk+zREZdapbBDFa5nGO4onarNHsBCW9iJMPgGBkNzLG8gAuflIi
h6ZK8FYzf+CN6mAGOcGeoYrywlD5LjOFik6V8Jon4j2V/BXro8WyjQZiaNiLpzOZkVCZudYkIfEq
8nwClmJXfaQfHV/DNUVVoeInoTQpfGoCeTeTElJV0FOANpNrB2URzPdmjw14vTTPaAm0dMZa6rhZ
s5N9p4kgF663HrwShiMU5Lst0NQsGwcUqnIGdWElPQ7d8u8IsPxgUveEiwaKLcilRwAP2+2d4O03
dORUPMVk6vUJEr9RwmLrhZqEbr2py4dI6cEu39YJ+/7dhFRg7OWHr8iY1lvRQPeTlcW6Jd3k/kLJ
ykzfcAe+A+C+U9bUCG9bAFZ5Q+t3X6rRysEBEk7uEpPELrbIXY4dcuB/Hc9KxNV0iEW5++DxVxJA
KSxScsr251Nh1+lkQl0o/a8Ri73GcCR2pVSRj/pW5ocpnB/HUJW5YU63ikDp8kQEdnjMT8nMrjwV
OsD8oYzPGMz3HLrGGsOIL+zUXJRhhe41anMDU5Owu0iKQbdgzJnSvtANyHmeFkibJQYNxXefSGO/
8VkwFvbMFWtF+n2Q5ESCKnr7ObMQOf0tTL/941yh9dxQBNa/yiILv9CeI0/h1VZD6psAT2sjcOj5
xlsIsjdgDARNqS0pxVyh869JdnKfpoEfJ1Cs4o6ywmBmOobtrqmgIO3wkjOfAYPKBmaLf8GPej3b
23cTtxj2jfoLiMPo/y1PHTuVjCM47MQ+admEPCt1bjRDZWYjRbmvLKk341ziz3T4hoG9FZ8A1uxg
SzT11sZVIIa+K0ehBME1bytxnil+B1lmcBRK7r9dxE3dVUer96lWx8peh3KpqdCBoxczdkPc/8V+
9cVNVlZHyu6sEKUaqIRpeKeNA4Bj9xBaL6FuNkTew+Xu14WQB+3ZYfBK8Dyd/Q5Ef1ANGIJf5P2T
QpGPOQiv3wMxML85R4CH0/SkqTCi1MZieiW/L8jRjr+Rm1AnnZKEGgeCYnS+aMKSGceLfZV7OYUL
FyuyEFh1PFuLuWRxJy0keEyod7GNZRuxGIEqZS8GtDjCJSpVb1ZiACL7VaX1Pq7pqKKg1XtiEVX8
mRTipNdqxOJuNaE1n8AzE++5DPIzNMJkfOVpO8ULgTcgDNbKOVZK0stlCQnDakwHz4XQSVMtV6XA
bsijDpCgAiSC/Uv/MQo7PEsqDJiciL/LSWZfQpFRZdN/V/HHtMmX7DL25lVYsb57U2QNFZaiEpfe
XCtRJnR8zGOrKzqvMjQSfNG5Xyj3lD4j+00domfdNfsXeDwUbNmjMyuvM18Wl7h2XQ3Ot8eONyxU
WtURy1KtatX9JyXFRWKMAdzDCPqv7TbULSBdiVHZI23g2gDas2fYd/aaZJACPReYiYqF5x/PPipN
9ycVUSfs6xEbF1Jtulb9Wa2NtMOoVCnOlPKSCNkWj6Oo183sP85OVcvc2k5BB6xTXI50cvBSzjn7
A96b94GlfxcWHoJnEcZw/lFkS1wb9zf7RoZHhTKjHEcOQUeQdy0PXND+bdUJPgea4zgYEKqp2r2q
rOWIvZjBoogh2tSlTa4z4mOKaNEQ8OrX9+g4/P8HSkj153sFf9aI5R1M/UO1h8TgzyKs8M+KF97a
28HvfEaXtPMPJYxfJIcOO51WIY8wbHVrMk7myBYgAgExsBbBwEa5MdQrjAK3wXU4B9jaCi2P5/kn
8gvO7L6BwLOAyOqHzmiZILrRVvZCsWADmG5E5ns4R8Og3hrLA35twH6rGz9x/LXQIcF+bBrAc1XU
vQ3oMVY8XIUie0y34VjQkv5QgEQ4E9F0XXDXUlMJb6iLagx7pBCIFXl7JTsPNtdTD65HDaQeLycW
Cz2LnVb3P5wlfpNhxDviW9j/Qs7yvMSQ+SxxuOb2brEWUqlmOMTyXX+xjU5XgqJAYD/hxKv+Mu9F
MaX6twsTGzj7okf46L8NUZT6LccZr4aidk29gA6J7N9kZJ8VvXHZ6DHuBY3GSZu4u3L5jPiUEJXn
Of/pfm2XjlYOMqh08eLzcEiLel7sLKNonx71y5p1gWbB6EHtpPOxdviGvAdG9xmx7NpFkAFcYAWx
ATI+kb3Mn56FDzyqnDUAwOZOeyJKIvPwxNGwdSlJ4axvqncWNAl2g3gi7DFXSKy3wFhh1dOaDnVr
EcfFKzVnVwVaWbDVEhQsCRgYFQrv/2aQ3o+WT8Gdv5PF1QvKFSeREsYN6g6tTZFMhUpH2R5t3O1t
SFomjObsGwQrwsKJh0eWLODoOZQbp2o0NUjTS2JvZmDFscGQRMzkBLTXYD0v6ZoidL4+wKLQGJAC
uOt0hofrJhls6mXxHmHFhuL99ms6mlOdIjvi6mbu/3HSsu0vin8jPrUPjrL4SVVRyDdPjPrlJ6ll
bghf2f+cLXHLSu9F2n+/nQAbAblh9qjgjIoAr6pXsp+KS+blmD5krTOnVwLDYi380jlrtYAKZOfM
mfyFGuKHnllFLcWrKtORrF/YfhMxI112Tlra5l5u/C2A2kMzUryFMejUh7vMYc+2cYKZCnzmMUxP
HBwAEEG92Ojyj8aF8OpzKRR7Bz94cyaKMmP9JqhOVzOag/JlVCn3uywPuZkHhxbR7/l5uGFUyJnT
PQhGL1a3B7BT1L9eadlDEa0Dva461H/2OzrfwfokdJE0zDfZ6fIy9/ZLVj7Q6DOTR14UGqw3AA5R
sGMSJkYYOA7kodPLxcxlPtoy9bEGUHwlJghA6f1RgHSOGiV4p4pup7YNNVvo8tzfIm3YwA8nvUIa
OP5olwtEWdIutstlvYl/CFZHyWRSb8x0pNGmjvTH5j8VgliYg9GQrMGRUzxAgrFXcyMw+ki44QO2
9vn1J57aVPTXjuf6OSaujH2pnHqFtDFXN4GjVKu0lkbzDXohdTOqccL8PmBvAvnxDUv0LHXV398k
q6ZD7Hzkt8hw6EZD+wto1QKAr6/cD1yXz51rObZbuuy+pktUTfc5IodP0SQNmLlS5AVNtKVuPYsT
fxA8piusNrHPAtqT/Mt9tKsNUWz5wkdCgoIBxvLvt/z1BsaESWChJBCS929m2/dQxqEDnh23kdXJ
SoivP/RdNhwuuck3ABo/hTwCJ73ZiyY6QwyTEHwq0+ZKDvP5Tn8mTwUndJUr9ZrfBPtoZMIxgJCd
wKTGMIzAHLEIB3KpXODVaTk9xKsyS5nogt8OasuGcbGDkvfsjP/GeRd2ngx906d+hKny+dei+HNl
TjtVAay+7wmEr2Ba4DiSh4tVD1XeV+5k/rgUSZ41mp948ouNkx+8+NkMLBlYTW8kUL/1pOxTkf4m
ZbeLEGxGnZltASCsDnJPHsqKZB+bugeVBBAN45rNbEN+PwOwhbwxmBJ2671P1hSNoaswvZhyq+eV
ELhz/v3jxr64he4Knax2Fktz0QfpMoRm+5P80vjiDZD6/yiQLsk8p+pnrH7h6dDMVoDpcnx0zLyu
BZ8znHvMCrjtH04qk5Mq5JEq1DZLXWW7sCe+erl6Zpw2OElmfZsV1iLCSPThgNCtNtGjWZu/qIKp
v8SkeY8ewJQMrBBm6L/qIKu4gfqMgGcPYhMTsb9ujv92BuqONwhSDwGoYDUOa7TaYNYOVtlbEBQC
YYWuOQsw4S8sg9/D2bqhtAc1eNWdrOlozwyd/52vjG9vE4ViCUe7N4+VTP8PQtBuo0iSaduanJwn
57CcHvONr2vRYByNAm7gmVEiTWZ0kzQj25nIitTUfexdCVUN422Sd6rNhyb2GLk0OeK+ZfJNA1LI
rgXrFtSLdS1rc9081Auv1JRUcZIXHhqDUAlar1E9arXOS5mE54SUWPjwHlKmvjPRAqM3QTvs7Y6B
YLoR2guMoGat8QYnhPATWWaNgC+4JZ360Il05RXCdI+kiMB2BM2PVNVFewMyrXIoDUoszdM9+YED
vfM3N+vhwU1wFu0pHfccwr3SDGpJKtf75woIalyicRsD11zpesKO7feihNWWSts4zefl87wtMhhf
7TBsB36dDxjf451TIWBar5pwbumDQHDJ6K/FHtI548nU566hyL/qRf/e6BkXqVZjj/dl299uyJ1J
GSmuOd9gEKaM/n5pjBvunvAwtPZt4Ei14j8EJR1TxtphRc1R8xesL5Dt3SigshPndpdTPJfoaBQV
nxzD/KMqH0f2MLHD5t/72+2pMdFUPR12w+8QcmRTGlf5DMztYixN1obHfpHONQWJBKXmSR3vH2Iw
vqESVugnkppkr5SD9kNlyMRC/pu5/vS754yjs4GWZG65i8OArIKbecxiA3vCuPnanMiN5tE5fQDv
TPHkZFOtAv21VC6kaWb7fWY4xqj/Wlr8I0SbTZugLnNChTByne7zTJXnooCyJ2a7AAQX57WSKC8Y
GOUqk0p3F81faJaxaO4zD4Xbhhz3SsoHfV2Fphip7UlLD3Aor6aeMj5CcgF7b49ZQyFxLUz2LsQ+
IctAQdOWjo3uXYs3HfI/IB30Mfe5t7DJAsZhCCJlzFoLg76m6jLLbiN8KSeWi9J/EgkNcOZoJhAW
5t3XOgSESI5AoLUY6W+eay4BySM6h4qkQ+9TvrTOMY2xlQhlgQncWSr6urCiwjNIVHRd/KK1l+Ug
FU6Wd42Qum1+TCRjEYwItYTvENnGia8njvyQy73thk8SFLUK4FV09iR7XYTrTIVbyNEz0qg0S2ai
2aQdrx6AQVYpL5mFRFLyM0R6RlnbHxHZzM1tdwKpoFMZPhkIycRhQkumvg6mWLZzBpQWhOWR/NRM
Qfeiawi8TuL1fjkCFRCXgzCGx3XDn6L2CQ7AaYiy3CrpAr9vv0qPFCK2MsEDUcEsg9CsSU5i9ZfH
y6xN0jHPoPzecb9RuEBk2d5qmDzY/BPGF5NsZpyTrIgy7WIqFUmbPg6M8GswEgAa2OZIEUfm5p6C
o6MDO3Sk1JIK/87TZ3xK4KVQHiI/xFo2yS901mnjhe6agj0zEv4ly0U1rCiDS0nUdRcfcI2ojowK
nQqIUXbNWCGjtEfQAxS09PW5jirKV1hdKZJRv7blb5Vafn0ClvNoHZwbKT/Lvy9m5+69dcpp09AF
SxXUXftBo4rSwxSPASHu3+a5eBTD9cP9r0tQ6rQgf8AvOhZjDidAOxHQeK+J+cDL9nnkOnVj0wHN
i9vT5XNlUq/fCjVKshDUPQtngY6brkcrL0S/cMAirsSDE/x14DmHH2MxafaYQ8pUp0BG5b1HEic0
cPx31iOigoK+TTfE6orNR9DOySpLPz6ocPIcEHuCeMUEA24xrUcIZlgIgNbCubp6LCzZwGIWMhBx
WYvUZlsKV0fyenlb+rjHy+9vBRScgTO1rxnFKPVhrLKVZ6EVjmlQT0JgW0YUPUsk1GYBEz77LTcR
itKEQgoVPmF/e8SEBMJbbSWQYIvxLsnFkT7iG4E62oTU2NTtmhj+aSpzancd9H07mxtZPhichCK6
hrJ1gBOu9fT0hjNiaqwj8hoz7U6qsRgSakQbsr6QyXbFKhPqinQDJkuAbiTDHjChg/o3nvXp1+sk
LzzDNNqNQuIJaiJmrv10nxJYXMIR51FEzn/XszoKF0M0Akl6okp3CdGMILX2BQfaK2OxbMqoSiAq
jmSxPwVpOLuwi53sb4VaKstsb5GrJ0XK1B/m+uTkGN6G5IhlzQxpL/O4Xt/9G+H4dADbpkc3V1gi
RvmmXRW+8kLOnE0uZNbI4I4QjprJq0+Lpn8jOp7+aWHla3QZssGNjgPeCgalKGCXp9tA/DiZsGgZ
00jGHDiP0s/0JGLOer8g6MGaDR7evyloDj2K3FJNnG6HCSj1o1J2AAEbeqwQxnP9ljrvbfaTTMdv
s7zgRapzbAeYdpN51wKCnCGOdqx4fqWWcz2Z41NoMMIzQY65RXi5IEKwkt8gAHoVHJwHRnICw5qI
/DjtFItlr4fpH96BEsA/RRNy+I4yWrcQ3Agr/Bd/GT0iNF4mSM3XfcKnjLEBgRKcG/p1TA5T4QBS
Rgo4EJsbzCxF5tIUxEDiOoAOjs7dSXmNl/eWAUO6ZhaAFgyTrIsHJMKZbmvmEgASXbPLNxDXXKVy
UezssieYI8R0dY2ns8c6ng7kvmHUKjevZdsUJPGHcDeOjLzuGzU2zF9nQl50SaZNkBeuaqUdOXav
kNxHopoV1hFh1gVs1oTAU+znShtTWFzxZIRUl8w8rTmh9N2kGn521H+IoQz9mmdlwJk4NlBncJQV
Natw/Pvj2KBySoa04geIUJYDSdrJ8CYtEU29xWBYHyLC4CYD9pDNtVhP/bohpmhDq120qJ3PU8mo
qsL0bMUqCGq3MavFtzmakY0t2cUb0n0EestiUJHgAA6iYEfQjtIpjIlhxi95gqo7Hr/jSFq8Ia9M
RebKptSCe5e6MOCV2D0Ck9j7RwR2QxxlQ2I3sCWWt47OZva6/5QP18nJT7QP2lqWuqr6RbxLC1Pn
mv+mgfj+DTwyzkRGg3Jsv/p7MKkpBv0jJFzL92tfJ6IQKpA5KV0mYu7pQGk76Uvk2ieO8mvn2qnr
ctVv1S/dNt+8oFw+zQplc3+wzboujW+iHoWz9X0b/MTFmN/uyOpcjUxGADJukE1widSj3BAUTGM6
M8T23m7b9BgMn0z2mvtpi4nrSOi+NWX2zNFk2CxgHeaKQf4TCLekrT1o/wy/sYCAQXURkJOjVXzn
xpv3h76RCa4riqOc14aNO23+c1pBD1cMHWM/G1NolsEZwCGneIHqad8VyZUVtgshLDbxxGKVG27U
1RbYk26tFrEtftcgPDAEsdlKYciGT190NcO4bfq+e9hIiCvkdtLTJCkTPBjgIxUoeoj2YvonLzwp
6Xw+maV85jbxB2p92phCKfcMB7i1jCABXH2FnRzB7KWW2eTZQNo4nujTemvoE0dgqCenpQHuJ8sw
zEmEJRAramnPjtcbcgcrDCb9NJPj3JdiGEveqdlA/8Bk/d7p+3msnqUJDYr9/OGm0ZtC03dNoCLY
AUCrOh2f8P/xU2M/ZX86CHe8ZOsi4dMg7So3dPtF1M+rJSU18y+C9cw2tfzMyYdvmIAUcPjZxBOr
NWWhunxUROxfR9Rf6c23/xxfATGNM5daef76/VkcH+k8OFMRkTHjbr7IQ5AjQcBLF83Kies6abC+
YME2B5CVTIoKsRdattJQBjrXHnhfETuNMTTbVwN+5k6OtHeoR9FJvHl2LpmHWN2WdkOUHKYLTkoc
TNoF/OxNaohOafcg3XkC4U1VJTsuB3OSh/GReF/bwNbxy/bDb74IeVx+WVJceqbfeu+W5u6Zej+Z
oNQGfTroASHOrS5S3pszrMR4/J0KCQh/L5KVrFMPEzYgqeIyK37j8kK9pvgiIfEp4ARuCTKc+Gju
46KD205815fVw37CGFqzGMRXt9qULlAEyYTyDXWw3jclrWm6kAZmKFAgighXQWIG7Aihp/q/4QfL
nPfIz9g7H5GvEwbzMkt/6q7bLirFTNhZHZuP36jSCpEzyUgLNnA+yIydY6B+THmF4lnTTZ2Fes3s
4cgukeWX/WwY3pYzVYA2ZX9WiLyRqk2X7LuJl+/PExk3/HGarOwfJ0b9Fwx7qFFPGTNK8ZxUmsLJ
8zfHdLGR9Uox0DKlW/LYYPK/VqrV52uEILGF20Wtu4/WHpPPOvKG0B4td9CrjW1dJ/QWaqWJPtuT
OElwn/zFMT2mqBWNnlU+8RMsLAcnZUqu4xsXLnmkJQ49dR4C+KN/lwwcv1EaBQjcmGqFoqsZV4Ti
Bcs6LDqNS3WyxwHWStLcak+x4uGZl28+lCmDI2anFkq7+xjd7pQ1Wew7P0YU3Ylu47ITmZSnpRgE
+djLs8RXL1EmqDalq8asY8E+J2wj6QWG5H0N7ztOmxh4EB49TQ3eu2fJflEYRC5Umo1hKU9EqZFg
mQ7/3E5uQB6rcU6Tv5XZTfBTeUrUMUN/YiK6EECUWODJYUTKi8gzEOLYFTZhdkaqymx0KY3mDvu0
Peeak77y9lC3WOT/y4TaJEpeXbqnYacZHvx+TyTpiLakxiwK15jaTpZKh5YjszZ2lALq8u41Y2W5
3n86fa/aX3pxSNu/u7zasA5cO02ep2GJjsAUq6dGyzepTZvZvV6N89KE8xVKp/il4Ky6VcWoKkJ0
pQUIWnMZxWIK4vrF/eIlVMaT4JJVNFVewUt5d8gP90Vnofe7d9SmSkbeMI1B/ajDInn6TNNVgZwr
E7OfpqYNoOCGJNeXiPJn5jL1L9jl3szeXUW2xP5z66F4wmY92nwat8ulU8SxNWetsYyO+OQaTQVR
YLkKkpm7FfIH+Ixhh+6nCvvylVgiN5dM9OccKVGIgdEYpnm1R/urLGDZljbD/t65Wb04JyUpCcQe
yjEnreI/168dJvzSkUxQ83dYsTtCdMJcZAm6+5LWrmsCb7tIKdw2RCSUPdNa0v4/tCMV6UcYMrQE
beRJrzqcuE82mfDThb/CHWRj2fSqgCy9TL9CXVgex4zHlmr1ng51LeHR8RvlBCHAzIJEREFJM9OG
zdj/0sqW7+TlMG6km9IHURU5i7r5FOAKChB8nc+tbWB4EEmEqxo+w1yggvSPjEVYFbJRWMWd3kMh
8uxzhg6k/JSWVyW1NJWH+e/L5/SaKQ1ZbfzC0Fv0R0g+1UZLUOn+LaFar0zIedeQ15Kw1mGLFP62
dhh49S+drn0Kia46Ml0zdNwI2S1TOKjADohwNmkQZF6URaIlN8m92QRoyloGyZRKb8r/qbMxCKsX
EP+3WClPVkbYEGFl17WPUh4zXlINw3pibKumuzss3N3gpahEmUbSTsXgS4wRHjbD88nk4vHwmUwP
z/mv1f13DJ7QoYKcSRrTi0kK+pQ65C7QI5FRexKYhZc2/6QDKmGR+mZBEFqDVytPVONmo6jZixZs
k2Bkpyvsf0MS7ETd65LJ/54f43/D3opYAL1NpdnVC0kzdDU3bQlAbk8yz1DwQAeztXF8vnl8IxsJ
gnhxVyaWAPfn58xQWiC30LEl6n329VTEw9bBLFmKazboCSxnc6VTo31MzDE8kOuAUWgfkE44jVMP
qne24j2dwVfMN5vVsJGhyVFlkTb7GckpGuluIoDeTIEjMmecX4Xbll9DATN65/t1mF6ElAROX6Is
G9e1uSx4CXjlrv5GeCidd6FW68/Z00cbWbFNS3G1idAfYQwuY5fJn8JDlQsFKPraN2N0hjx+Xv1X
zpzUYSWZ3jT7k/BNc/opl6jvqshSazK2javthL/dTMRPVamD3C7R2Xg/T7Zy/fesVLfgyBCXeB3q
jolpwgHWQTMdDaLXZ1Qnbb8Cm4xFyvBtrcCC7Sovs6ST5zAAAFIx4kilF6ja/P2EHZNDJGLWZKbD
gQsGUfuKlCYaY86vn0SM/0RUVgZ7mrM3D/m/DAWX6fJKqI83/P0drnrPTKQzu1p0XM060IKluBF6
aw7An1tjuTY0FhN8wUTaZMhxBkWHwkBMTpGIZGiOKceKEtD4L6UVrBOTjU+vwRQaVt8pkirTaLwd
7fcQV7dBHJYxQ2TR8b6wwN/ZbqqpuYuhYJlh3sv8WGuPPo9OOwrbZdvRvrBeRAXtKJB/zhNW3Fik
Yt3WaBiq1gte+lyIzpXJ62gDWDwKMcche1cWly4Ixa/ihS3UFEKe3WRcRgEX3BtZLrObYUYEFObX
58j2/4texzHuBNEPMIehSJ3KEvmmFDzmzsafrtkGMGdmdnIaaeI82tBXVr1u0lFq/P7Cv5Ubw8Kq
z0xdRUEzs11OTCXZ4nxcr4cXCu0u1LVdEBk2Lx5Z5fSHhI60G/wRavfksh5cOrFvZBBxkw6FN4bM
u2ZHsBqJs3rF4PL2+rjV8AhkTP0JQjk5RKmYZSc4ENfSUYZ2YOXnt0yPsb9Qi5b7Hb5OMLwet87G
UlsTLnstuyDH28mdB7eZ9ffj4oG8orAtsWpI3+OTo5RA4wRZrDa9x3XUXm5V0aQ4wUYGQeHkIeWo
y2GQaf95wT6SVFGJRGoPIvsGIbcKJyBBeG3YCK9ApIzm+ZDW4BIrNhO4q0E4uRFoLvUtyGl2j1Ks
/wh+CLj5faTmH0BiGwgWqhLe0FyrpLfdrodikZFUQLqqBPCYJWl+Z91D4YirNPAkTI8uelZ3coFa
9QoaurRx9EzGcVR6MiQSR9pXpIzAUXV9mVY24osR0IdZrLlEP0qMJvTUjsiQLEQlbGZCv1NalFBg
EE4l1uR69rsvQ6YGYJlEjLPTEP3nOJd5wNXDhiwl4K5jUv7dmnjQKojk5dmvn7Lu5FFPHYfpRD6b
xYfgsxowInwhHCE2JfBYpk1/2q5KQ4yoiBCrdRfCQiAZZRGuw5CRe1hSQDGCQHZE34p5fweEhX8H
BcId6PL3URA5xym8Xp0NzLUuDruiOIvyeaJWzNJhN3e8OEs5ccH9Qz87ZTIMP1XeU4SYvPZRtcbo
x5I7bL80C++nMwLgrSik30oUPO5fYfFCKZdYEoA4Oz9uSrgTXszrg5FoPP/uxc4wwgmo/hc/C/Ve
JKOsdgtNyzOrj/0d7S2i1HxSgZ/0VtrL4wdOojvGabhk5+36vz8qdBA3S5Uz25xbF7Pya0eWYltG
dRuo4swnhYwCZqqbfCeaIshVlCJKKcTvvKXcf4MrVDHwYxyTGr0K7faCpE4sQbRZuirlAknSw8j1
H80QszvfE8AMbKj7ss597XpX1dH4oFeveA4Pz8TUkfGXYIa3NifdSPCEAKE7IavV2nRgf2RcpEW9
GH+wvoszvCqLrHDhCi+O9KtS/erdswidvp1ohZZN8AIod7sNYZXhiqy3pSexNE0vuHYiOUfwWf87
QQ+PoBDc7/Qytyhg1G62TMaooiWf3O8+hzBH621Ud2jBoFuNpk7Pd7CmkbonQEHbV1pA30YMcoSa
7qhdqqyIlAlzlbBTnxumDzegRXaVBKqV295NP+9W65l+TXXc717KaKx5iBJDBmzEooiji42jQnDA
zadnd2wav4Z5rL9X1o/v64eBVTSvcMxujmW79Ub2sfv7iJNW1rteEUG6AeA/PSgL5+aMb4DuK8XP
FcKHnRd4F3QpP4cTcmpOzJpCZC5au9VdrWAl+Za5RlIRalyYB9iO9Wn+MLxbnxOXjPQsKvXW3xy7
GPo27mKILP4fuGmKXvRV4HFAYXs8E4mX71QxE/99zAhaGQcLeaTxQOBl5CUD9B5PyPgWdtw9Bt2v
D9oaDNlbr13/27g7rOMjst23m2X4UNntcv58nMOA+mXj5u7cqVGyqOj5YlzBZmA22e+XHdv4Wjh0
OEsKcFKdbHVhCJC6CtfLK+W50DlU85zJa98pYDAKcE3U77VtraOOZdqWESaPMJ1AhkPgrKeKOBNl
VL9abzsqH+UZKnKpTJ0atizGWXzad/kdbfAWpMkCwBoTO5B/xvbvfsABq38Y4D4vi57wmJ9mAdUN
3WPeRhxNwscQd8qmRTojkefMZscT8sGmKHBi5t+IwqFnYScrC3rYH+IgloktrBsG+yTkt9IbV6F7
1XcUTyQ2RLGmKx3E5Jm7pAltDWpN1uv386odK+ByaUdac5J+W3O60AFcnX77AveF7UPY94ZEorJ6
+272PB3lNy6XwmijE0Hcd6m2/XaIA1UWU/wu+pj559+q9F9pVNyRupMZ/aWKqIWB6OOrq8Cz4bPy
+QJTeXHDzmPSTq2LcLaBTwtbOF7LTP1urALioBfq5sVvDnF+p+i/qRuqIjBlNdOLVA+goClebnXY
oBSmow1ZSS/VwLK+tY19TIXSafR+MTFMeDoZW0AKOO4Ij/HedSWfjoolrmK25Jca+Kkc5iR9mDAY
L8xcGYtjLT0Mc3Q+ip7ALqmu0sElfYd9X9WgAgJ7nxImbso0x+OGvDTLL8jCDrxHOXtUTTnK30FG
cBR14f1bPNMyFtzw7QSi//eNykcznOXOn09Lwfie3BolFFPja7wX1re5kWAW6SV69f5hNBzwY+nR
dgFhmK+ZBo0M203CH/YmgRFs/QA2YtLRCXJr5SwwHw2/EAU2UE0wTe9kRKzAUMn2rwjqxpkN1EYp
N8PiK0nrg8ie8UMosgWsJCvU7htv/OyPQI/L23TSkWIAt6RUyjkB9oTU0AzKt7tNNeXRLBST/rcN
A4gAc/73Fh6/xr2hF6Q3U9mnQ8fNfgqxdnrzsY7xz+5xMah5Rr+j+e1kaqhJ0HMfpl7zcIM3Dr49
19C51tmGlVESXEI8xlMoiaYAP1L/GYFi/o3GMeQ5Cw+si/aEGtdNLifXOmtVMkAzF+PFS/H33/5B
vMpJz10Rc5KLIqfm3DiIRzeBr4EsWZ83rS2Jyqvdkx8BfoTw3cMtKvOaW4C9EG21DfJZR50AMi3H
7YtrN7zsEqRTZ/ub5jO7p3sxQAYNkSGPMUkOBzobH7MOvAko/3Zm31NZaZz0P/SGvpMQRX8JVTP5
yKpuVcJV+R6yZG5GTMyodAp9UiQscGTl/6ffUXVCnRDsxcxec8mSLBbgfVU0QQAwjtWLF5lr6SzP
Lmzpu5kOdCJXtXlopAGWWS1UKkwDxikoglLyNahBkdVtJCdf5gbgj07ZwPmHB7mLMxnWkSEmKift
mUTtAwYDcNHNRLdUN0dSe58ZiS3wgwh/oZLdxCLLyyZG1qQxgqJXnCUSXKKSYSwnSqzm5TzM2opP
7tfFD18Dgix9POri1xPguzS25Jo83HFVyH5L+sYRyIxLKYGts/ukIXS03MVm0yeZ3OFRvkmSRzev
bhaJErq58aOhgf64pFr1s1XxsdoP6FpuBVVgGXkLI4vuMuIhJCvrtpuruo1wNR+KQH2T3hXh5BbD
d0xDSmh3bSXglpV0AqLGkw7SBPXLiFcIab03hunXopHx2tOwYxQdwHJTD+xqknzKZLBrHsugoPDH
M+oDTQP5yFnkn2g3MM+cuyH5VJtaQznuvj8/k5ZBnHjMoSgqQEjRDsbVZPTY/CnEi1r0pJPLJW6a
FzTsJVGL5docaxuUGBKMLDq9iB57ouW5p4pk3r6qdx1x1Ad1c7SIMYeX81vvFs4G0oxFBEbjU11N
nqNTZvYYMS2EtUAMtBsfYYJ3T3Vw3W8EvT/ky94YVeV2Sv59muWQSrNqk9Cc/nX2m/mTKReXGPMc
00SR6DIZ3i5PyS7k7gg3ouGbHf33pHqXq9EyF8ju5NSG6eDuaagKFYPs8e+tvmny1RLpTD0YNqYo
jspBK5ZvgMLQLYhjjFV9nDWSRLCDCVrFtdIjooSvZmOMM2WnHWHYkl6rtoav1VmHX0BpJF2Uh52j
ZH+dJeL/3+uC6oMDY6/E4EWJK5WkpRqfJDrdQB4E/5AD5sYiiU4G2db8mbR7ewCZniK8A59akzfP
BxshLqd7WPu9FU5xkOF1jJ4lVCUBZGMXQ9H0cOvwzHobGNtF1sbOheFusCdwA8r945nFVju9HnW7
gUCMF/PJVOD92+Adt5S43H5fKz1a+m+HnuZuuYwUffXPM64k2M3HYGg6XLo+84s5Deq8OZPXumfg
VRWi7WthxFl6bEPt0yd7faGsfYaqU54wicyEIqUMqy/ZvsnEQkyMMgjbkMWN/oRlgI1WLyljqqzr
5lQwpItfnOJ2DWF9x8hR53xlbpkzpo9H9eCgi0lu4u80mNcR5v8uRMAedOf9kQkGQYWNXYhWefOC
abqbpg8EMLw9Ptz4onxt1EuMuZlHTy4IC5bIT3xIh8DY2XeWLqlvkdhhTsNQI7NR62kfZ8DxGlE0
jyYpm9mH7mElCtwjMoyCUpQtl9Hr6W6Zg1leG+rdfA4zX967PiTnKCxMsJZicrqFE+2NUe0FAdVi
DKALPWYXbU29F2ZNhJq07d1nunYLeZ9iHiqCgXHT1Gl8lG83R6+gY1uaC/QoeLCQVZ+rrGgqkeSn
+5AFpL2xpeJQWMWbFRUZ/1NBIKWTMa3rdRbOt8t4+LGtkhMqfdni9i329B0JR/wGrL0ZK4/GJ98y
JrVBTphTfsBnUMNYVgtsz+/N1ARSZHb0gwxuer+i9fQUGcHARJyMMRSVJKiUP94+6gZGSmWXVL+f
wDNLavRZLFCbCn9LE8OKo0slhqmg1M3Xz0NyohcvpHuapMRS4HLjBd4YeJQ8BEkYSH2kQOy8b2Na
gs62xVfBCcNvriWss5EUH1f7HdECfBrY6x5/PNIKWWZeCGezAvcQuBAnJmnT3IMiCNsT2p6qUKFc
7vjUgbfJ7m70QRh9vaYMtImb+vwzyui/TYUTFebC48jcc/CXLED/VxuL+Ct8J+ChqL3E3wPrvLN1
WBWK1OII9DgFmhxt9C8/mQpU0BLXeaJz7fn6GikmGmmMriHvSwCippAYBETFgy/ok3AZr8T6FwlU
RA1vASzNuoXBatEnPSLoMlKWcdXidsLbkkmYJgA0d1Kl/CgUhLLfFnAUzsf4is3a9ztGvqOZWvVV
wIMdYErjQ0y0uS3GGXLhrWcoKw4MWjWX5W4qPyLuT3O7kk/GDtPaRE9S77b+Gbqi7TAiRCIkgY5S
W4llYjcOFfITqvGmdKZGrJs2Di0jNAJIgNrCMJf9Dv7wPklMq2kejeAIR4mzbTw9L5LJNxlSO/W/
qNlPijjbhXywhvoGN/4uedayKunuCwrW62MbCGg/6w6Uy6pS8lVUNyasJqrMoXv2w4lAjeUQ8BcT
+oa16jLeav8vgKW8hTzOm8RzysFy0yfEqBex+28rSABj8Q0qVAc8X7hm3USanOiONwhj8UrdhNPe
+mtoV90b95CFOrhCvXTIj5b1QIwmRrEYFi4kiTrMQfjTwsO4Z9VYDvzZhG+7OUnTWmZAlCLNcyFd
qMBD9z1Pdf0uxEk/JVGnrzl0mFAT+cUhMr1Wr6SDVK/kvfK/R0FEfYja1F8pO9PQ+UhK7MZPRq/6
Ae2n5JrLZfhOh/Q0relhAv8jzfU2Rhkj5XNORQhzWGXHgW0MVc5ZcsWTFY7nveob/gEodS2q3lJZ
WandTB+cFWz1IZ8SotEkehCei3s4j8m+cmVdMLUcNM+aQQxSLpk4IUiwltXaew5+AwHY+Iw2zmLU
hoPHSPcWcV79lZvjz1+qTFRNYzO8JOxhOWPaZAApR90VhtxqSIHXcbDqzBJJxkRs5MbyLdAgEtY0
ob7W3/f8qzsWEU9oqzjYHG1bhtQ1xgLcMNOYI9WVwADqxgfGiC2MdekrSt5Mm1n+XrFiFehAUR8S
VsIi+LnDQwhmCz8JLqERInjQrFWk0eCi+YL+CZKuKWJAPMM/3PyP/fOitEtNqtbFoHM8EAflowc1
IJ4rQyd2cMUA6wosmym2mVpVhviBTbNwZh/XlC0TFcS4M/6XnMSKnubM7Djw8w9ZyR0HeovsaH5M
u5N8r2tvaZWC/D10O5BSK6NPPk5ttk1jz7LMJOJ/banXO57HO++4kpE79Sv7NyIA7twXWcCDdPxb
nj4i3oXIkuNxEvpLdAPYvJc7R57IbZtqY9c7fyO9UCGHOPmfH0BLV1rCyrOb7nucRR/9cVyYfeYs
h2abBocYyEdKFt6JOayCY174nTdSzUJe7yL2YKuYbfzIUUgB+0+PGd90K7bzZW48u6Fcs/0we8Dw
qa1N/nzSzAZE5yP0uaJzIfuH84fZ7mRWWSIzgIqm+c12DnhQAlNjK9T5ZFx5O4bIOTNLFq/S1YDy
YCsfPwoKdr3lcdFSDwiKl/jEvivLMItLt0XeTPe/ObuBfVmspjqCWuUlHDM670zNbeslfgHODPZ6
bPlYjIwyHNsI0II/b57Gy4S8idcpvUOjCcVjXDYfXi52qDbHPmyG0g9xJuW/yUMvbzNqm3d/+vV+
m86bw25i4tTSGUYHqPUVNKZ7cLVBxk2jQ/M1r23r1XlSxRqvXhNVf3KvLOIIWkwCAWEuw/o5qZbu
7LdbUDxlDEDQN8iAXdI7My6f9GVzZAeI2B7UOcfQeiuUHUK8nacyw1sy1sdLQIEqT94KwjCT0vDk
tSJMr+nd6o8VSRev/oBFkb59Ef/sv7vhoUXDt+PAOcwJwYCkYtxh5/ecGv8VLCcryndybjSvg4fs
XVfyX2LUrmwo/eziuhtY5cZdxkcqrWpygBlxKL4fpVptt+wFhvGhWeF24qEf528U56ZO6R7/RJjU
Mt1rv1vbpwf4GfdWtaeHUDmvJfklGrFG6bZYbdWSwmNiaTQfzFUF7S8xbKC1m8xM0jyFuvIFlzN5
yVF2k0P5t2j2LN84Uf/aTp6xvFzs7281cNOUUD5kf8rMUwpjXUUc8Dx1NahXnNinrowucAGfavQM
z4OJC2V8k/yVjXu5Ab4PdRt0LFbhUdN4Lq4GE8extK4NTC9Sdlxbl4Dxg92ZFcYT0qqnYoEt4dNe
qL/unOWb+DomJJyWBL4p/ocGRZTL5c0ImuhFXBo+ND2b5mrOVjTlRUgHg5q1VsOhFd+VC07x5ydV
Zp8+8Fphrx5AC4zWOfeDRjoWt3gdR3cw8rUn62gwS94L5zzCfw5ulBjvGrJ85iH6gQTgEHlXBSVR
C1G4hnsaUh6PdehpvE+fRndWkYA5qCP1N6edPiMSTE3d6QOJnX3wqdBWUPNZSuJkwbdoiXPyb+1L
Uv4FqT9koQRVuZ+D3UvYYmPXzpNYtRQ1hW8owEvw4B1TZnypI9QJdhFdrvdNB25Ksc+WilIGLXbu
fW1VNW+yzMXjW+YP5X3/WkME/hKW0lAVjFe1GJ3eQvCTpRhNf4/WJCyKXAP7R38JonmystJyC7j0
CPYTigkL/6mJoe0PXycprD/ziwGR1DyoYAkVKxYp7Sge7vjA1VjCCZpnnBMo2heRMItRdUHC56Q/
M7rX7cSj6SkMTWKhH1rUPv/63lLWwZp/Tf/99iH671tl4zLOK1fE35izwxir/S7K0vImUq2ose0C
UQ6GDQeuLg77KtVecL1mqDDwIitqaWlKQaFUsSv43Oh4UnbHCQv2tau9gjwCkyN+CT/ZpLfXfCLQ
k4nwBYAUX5fb2aJzJR0TJTx+EQaUEdrkKPMzpsv1DLuYbFMVEIOnc/A/k0Q0CNP5bll5NRjOgSNz
Q/t7CwCr+Qa8NrtDwUYkA6et6NP7D2pIm8B4IVH+P2JtacYLevOBzRElM6CVQdssJTmIm2D1KGma
nMCr5dxliR1eRaxa70IHtHWTmJ3QXzeW4qPNUQvJFmLyoplOkQME3pfOCw/AgzFlPIRpXy3MS7SJ
Ilc+/o/iE0dryBkMoTDrWry/QxBacjzvDryg9xUh2/SlyBwyDBHBAhPcSntQ6RUsuzzRYGWoUYD+
Pxqs6Y/3ZMPcBTP3OhzulDTrryil2/LwDbiAI5ha2aIDsq3Zn07O0FQHecRrkSR78q7cyTFJgbJm
xLOIIVznW+iMoqXirEgvpKEKabJjmrrZnsh9XdL5/L4qC9m4PxWLZK7XaFg3NXbrOUUwGDQpwice
kHPFHzq1AfacnMoiSAbeOVIZ84ft2XTvhqoK6mP87TGgnTlOwtkBSTwxPpzHARAW6qU09DWhunzD
Laxk0XZbeEqmBCWuGn0OiROQHRktSyfR/g1LXGZlIjLRUsOib9+TkOQwU4hA1KuIeJwVIY5uHM4y
tEzHpiNgzcMCMio8UeRiNJrDaHzf1PUmMgzWJP6CzlBTQX2zyBCjoFT3rb2YFL714wYXXrqIuQw2
D037JHamBs2Lgvjv+/hAjLZNTTrI40W952K2RtRp01GQMiskvNLPSjNIfv15O2i/Q64zpGHTmB1L
43WppbDxu11+/B2uR7g38jbE35YC3+d31pXeYLxj8yMjs79dx1vMbsCe/Dw0JBGXWP2PrbGRFWFj
l95FDN5vuoWmE6lb+NRb2QdvbwinF5ybuhbRnq4rej4LIwOCz+MMxmXPt9jXEiO3lYd+ZZRONxcI
8v59xoMRvS7AcUH1f7FMOl4r/3tShnpjCCPP/c7JsbWDfVMXzsFssf1O5cq4AAVSzC9J6zqpG+QN
fp9skss4h9ikWnhjxiHR/FKwFZUJDUTSqScsnvkJjSWJkn/2EvC0luw/E39AA5IFzRi/tllBBdAd
RdkEmmbJ5qJiyxn0nOlXmwMPAm6T8UKlsdvQRV4gEA8XRy4b0CNRn/bNyTlfzs2HAntUlDN9BvV9
z560iTJEu04A3l54xuSADpwiKU6IIWf5xCJdaiIljJVEVhTkfIFKJSHW4/9KCo+WydCJfJBXCviO
pqGlmnWmPOwQAigp8mL9CLOKD8M6fCL5gWMyDz32Ti1+WuQpfV92i4LCaUyA0hkkAefjkRJjSvuJ
rT8JYimu6kl7JYflyRawIWQb4zaC+94Q5X7eA6zeumnqin+2TpYbBNcZKZkP8WI1eOOMLEblOWlX
ApF4Pkb3dNNv9Uqzw4XDRz264or4cvTk3zZqNfrWoKT6cIQNfakGLfoAgYL2wd8+u1HbNAifQ7k/
fz+Tps65TufsUOKBhHeZ6SXcsUM+laKxnl0TOixYcYmyLk6W5fbdUOPNWmj2yrgUag776TGoHdqg
mPs1FAhwSsqN6X9wlUQFAov4iibCSvGhtZNoLoYM2sY5Opk9KwUvQkfYNgMidU6vwNQx+3rUldL/
vdiQC1NA9IL6t2itv701p2KjOmxrDCegsY7/wPc/WFb5mUUToHAG+PdFheShGcRxOgNr1ElpfkRP
8h+gVTXy3y3Uo/kRUj48f2qZbVUeLda8TzdB0Uwwi2hOSR0pRm6/RKHjZHXsvgjPTRRK5MDDyjhF
cKcCp4rrzv4ojwIDOw5OCgIfQaatk+9nQdrmCXc6TUJb+mhmmBqcd7AuxcNSxxzsDYhYUHkNGzHx
b0g8enBMo2dxLUQF4k0J+OIdFp6u/sqJSYHx5pGAR0gDpHo/nQwIW9Uj5nSwSZjRZKdcn8CFbN47
loBXdvFpXQ02c8Un66EHtL50HYgJlRxSiPKlft21lc+3kvzhrLHYJJympgMM4ZoC/THdu0Uan1N/
Lv0QBOe26bG09YLdI5e8b9/h2HZ1Lu/9WnC1lvf+UE4ps6nb9jMtxV2GkxCs5mhNaiMzw1dj6aYy
J+RQ4cbPQwk/W60G0yIGqsBBSAVyC2uASaiH6EYGY2rd1UCML2KtCzvpVZJ3o6RZ4Vlem+0WNlnk
WpODLM+AAtGGDRZmw+sNvnKlIbiLoeIqz+KUineDPsXWZOHCpC5+Gom9S7cnijcMsZ2OztdvH10e
gptGozOGiQ9NmQwQUhh4zx2v26A07H65thWXX6nUHOv7NQOHIwNRFS2ZJWwcBLKQT5JF1icH0Ci0
tQ84S2BdhzY2m1x/nvTBpq3sv3FD126Ji4C4ZJA2ZknuZF0ZFrLnnHKfE3K9aPnmIC/SJ9WVU2xe
lRgW/VQVvRLLoxRJLJx1dS8aiDLqDuyQr/aOGExNfFlnyCjOlnjcp97jTvAuor5SOLGEYq6gDhR+
h01MqX1F+0hjwEA66QzbawJJOP6HNyf7q60BS6lRbM9f+GdFUGGWL+AHSMajob/krUPHfcAWsbv3
YnZtBwkE3RM+F56XvH4llVMT01HnoCE48ySlDOpnCviMilzC4riWiMtC/cLEgnpMFHowjie9oAom
sQgqG3Joguj+dE6jhNG+tUvzoiR/vrcksl1bFp35QN5xrZPiAKCaQVRmmkue94lnThcUMZ3xeRhw
DQ88ESnAAWVoX3wfhXuFUYoxOHsAaTlQfbCKmLNeBK+Y6ToBatA9otqb3zpx025iF+s0qZ8zQmup
O46+YSjVrwHa4VTlqLF3OYRVFihoYtlM2HIf9YsOxkCv1HeGprnPSuw8Qf5nUtFQ5+uad71LjlLQ
Eax76IuDQXSdY4Kxa/XKVKfYtaOCLlzWMdBm0wQtMV7Kln6klSn2fYucOXBs15aqlBpdly2G1sKu
y3YXg9fXis/JD49GLieU5gnFdxKw7bcifloCcA45IV8RjQxQ1DTZiuTx/KvWlbBcZYqOHisqmWuJ
wj0lS9bT0tl+tjkHSv+MP6nsKiUuxcYREpnzHWm3ucvYl3h0jy4WTC6czVRQ9lb2bLP/YtEgrf22
iMHB5AulO9VYD9Ts4/HVOmT/IGb95frDAav+uWo4jTb+oDtktGEiEtPunj6lbOXy+sk8Y1h6WMpn
oS5l+ds+rpxt5lL6O2bbxbmrjU+sWFjpfg1e+IQbAWeRIxMbizg92xzXGNU5SsnMMYMXlo9SCvGp
yncI1IWmuarvEVVN9m0Wm0xjWY2o+pzfSJ+A5ZfiDK/8eR8koYIe1SWTZmh9Muj3Pv6OjjH1cpHq
KnMcxqUwuODtIp3Z7iSt7v6OEYFxBTOh+9ucWKynUuNKHqyAY5U1nUhdOcEz0t3rxDkOYd6UNP6J
pjRus/zo70Qyt/ULCw8bf4WsdJzBDDeWT6cith6+/kc+1m5rQE2jbD79gcvwrnlg4adXjY3VIZ66
goWJh1ZbZcJXoMmQ2Ngiz1qODtIy5anXuICE2x8bRTcNYls61grglY3Cp40bYM6CMIt9BWN+o2T7
SU+R/f/3IFRUZUhYwTZ5Je27Aw/7gB7GR+8gU5eLkvd7YgVfagioouX6zLefW95Kdl+qtZfc1PyF
Wv8nbZK3dGGDCxmAC3VzcG3POKO6qQFLgyjO4PPjnXtkiODxP7MYR/fMWVA+Ni6Q+xKuGz5jwacF
yAqRbPugcvN0aFEqs622hhdfUDxsr7PQ+9e/vdu+exCOo3TQFticwrSaQDE7S6iPmydy4GubO3D8
j0eyrJLLqVCTCUDM5xVDuVphKJuNpb+BRXsbHlsE4qHl70FfyjtklmA7LOggoJluYZDeeYQ+YkfU
jNuLKqNuK3F1m35SzFZVGPbx2wnJABoH7553p1t1GjEXZgn4sxiTHeA3PpOnBNck6kkE5aHMPcI3
R8gZLL0JVjYRy8bjD7E7/9S9kJn0h3QfIdrKxZ1PVlccm857lgNDqk5Wmy1SnE8db4NNl50fI2AW
Nyu6iYZpIXu0Tzs3Q5FFexkrck/4gmnc0HLHwH4AVw98inn2uvZzcPxGbhsXc6UpvOHDy8Qiyovv
D+exh27QlxnJTBboL4dlc5yfDav41yBuni62cNdECiDmx3XCKFlkkzCdGXDZc1vw7CjHbHRPKOfz
ROgYr1Lzzd/X+b8kyn6yEnFFQUp52BBNJcmV+VaHc7/AaYBlb5vS32JZoKu9kU5tVcbbOGaiA+gK
Zh6B1E0BeKOnTF+ASXATrb4RrlOVfDjr+uOgrrJ/4nSJTcIncVF8sQOF60KFEPhN9mMM+26XMaTg
uEGvaKaGeWBjthS5WuxNQCNN/Abjos7o3tvn87HYtxwTkL0y27RG2uglHFig8BxRdOm0qCS6Sw24
K3iDYo7AWM9CESuzYvGzfX718E+Xxwg2F5mQrtIRYBVjAlA/WRXpi+HNEgKbQvZy2CakAZ/dDrPK
fMdJF1T6U9hNVfdecdHdsDWStWxlSanZBqPtWtfyOG48OxtZdBCx6FQoMxiEL4/7u5g9FlzPTeId
zsQ6+hHicK7Oo1p61IENJnq75mtNb9t99Do4vQDkxU+pjS4i1sLM5CIsGWJ8pZmUckWnwMPdIqJw
ZgiL2y+aIMl3lw+jq8fpzvF9En+bbhD+/nV86BNRGSczlomF7By0gabQCT1ycYNyI4S00+/NHlTu
sY6mEXj5dkgHnlc95ooWqW9Df0bGEjUqpy7HIo7THkzlu3Fblhn1Is8VQWyEi2VffjAFOeX+VTUb
H8DEQWOrpA4NvfJ7d3XJO6/b5Q52VZ6fXxNFU6oNYn7bgi5BSzyJqbw3+9VSB537eL/1SoYuyPmw
91uJaFusT+n/odMqJhxKVUryD7ayMuoicVMFgM0jSjdjQjfz6slXE1pa4HNxAPFiaRQta3DlfuaD
oRp41BJzhhiLf3dpURa75OSpwXqETXHS5+KIZ7KlXODXfuIP2L9MvO4mxa2rtoA+rlcc/SwNF9F7
ZxPqWx49hzz/qcRyvbKNTat/flBXUPToSVE6M1M4wQZ9g/38rMkDI//PfK1+ybOyyUzY6Z5gYcQM
C/pZuCwdEezvf9SlUwdp1H4zFUvEZrWrg28oIUflPLTodJJcQ9b/cUcev26irbF7ZwLVEJz8Cmhn
oyuT81Ldhc4sgRgSpS4tTw3siyFdypeXgFAIvfeFJTG1ahIT+U8JI43YSCStBr84J2rt/0xwB+vl
/pJiZXIwQtbIgW1zQeZ03PilbWd/q2fvSEC7Iqd4j6xdDwjxrdeIETgBQvkZHW3//8VTiGecz9Yk
q5+SGpSLas4S9KEIfIVYPzAwKQ8MsfiRos6f+OyprclK6KsIlOu2b/s3SEhOHO2rzLmTklEZKrdn
1z/OfByOBIOoukwR1DPtCgZy3Aqo4GYA3gPZ75XrZv7MEdOjYDkrwx2WxRXr0v1yHokjN53CK9cx
jLG8+lOknL3keUKzzkeJt+nq09Hc+WDMjn1e5RDjZWW2CByxCpv+45gZjrEwDHvVGDjn7fsoaaxt
q24hXswGxrcoYq4jw7h2Tld42V04kyIDQfhpVR1GCeQ5QmkU5ZEjfTZB8zahLeXXpA6BkPCmBH6b
aHp3u3OyjnYr+y9YAKzztnW0LpLB4RQya0L3/Cve5t7WXSfIlBJyE85qvtSDJc6Z1b40Czak9axN
wGqnd8UHWmcaQjjJAsSCKhIavZIGD5VaXBjX1NjlGJntZj3elQYqpmfIlLiaEKqN0/7suVG8vScw
ILYlxSDE+R/3pLSA/VQEKopmPxvg4NCwgY4RQbajZQXb0Ux41e8jjStTUYahSVGZWhRMDGwUymDI
VQYxLfB3EW0s6TPVl2+aXh22kR/56x7ID1TIYgnzyHnlopGFF6uTcFCx0slZq7v8oQb3z0TmsKb/
uSSuUU3mGJfEXYTzQqjPJCyDirOMCU/FBlawX/0JrPfL48eFnsU2/jV5xfC/M6l5P0x6gHC4+d3U
SFSbJqfPqp2uqYDPdbcIBE8360+VDUOP8G1BK5LV/xu/doCv7zrNkUIvQtGze9R5gkR9IArirwXh
6YGsmtavYgItigKh/rRbzJQgF5W3sRNm+2vCMZA3bw6DrSruuhUvh0kshGkACv4xpQzk35vWHG2M
ewG1teaMpUps9yzqbl4fah7qAaGKq/h+aKhtGeJSf6ZLdExFFDzuXpYy4b9OUg6WqWryW6E0At9U
zCuXTqd/MoAJG/UuUrkgUO7lcPDpJubgJRU6aL1ai2w4mzlHwrOC1oOar6FkrDu4uJZWUzExCEQF
frDg1pzjCCeywzvKVQz3SmEMv7DNFD4ZNjPPVRjGTlHXoS9G/PJW1diCwm7BwWPw8Kv74a2ksyul
rOZEkBt/0X06F+/LoziRt1UB95csdN/S5EM91x2p8XCpw7k7Kmy02EcYXYfcTbfIUz5sIYb6ETtB
OYId2yFqfGSQGfBfFYzHG90rCIX6PoBjlDNxazWnneNGyb0rd7MGuVAYv/eOlTXZHcZyjqO36LdA
QqD1l6bhY//zYxYRx2oPDrLwMr7bAUz+CZUe86w5otNixu9P6lM0zdkAget0U4k2mas6Brx98j1j
SPjv/zg61bI5gXAlDfS6di2d1dchz58PtZe+Cz2+ddOJ5CW1eHiRe78V/5m7n7jOYCdicpLCuv5t
uUeTIj9nRAAgt2Ls9kcBkq2i8Pd6CXxmyHKGMPP385I2/fbRU4X/w079xkf0Zoj+D2m0/PaP4qI+
7qinu5WJ5fCtVSwfuSplZ2JmRZ6x0aOo0mUYFutVx1afq4WpAoDmpgRFfi4+KA8pusxhlgIKB8vH
DkaQn2vAo9fZyAZNDCf5XvpMN8GssnIKcxhqQwBQFNN6M7BqMusFc1pAe4kTB3BXSu2l/plGtoAS
IkgydaBpQ9xNIqRhvpFdu9JR0D58kZNIPLMuJxgs9LYBcxMxpXy11byS6bnua55UKJP8w71rjfPV
NToG1nzaBtzI8F0Idcb90iukMjvvF25eFzSiwgxWI7Oy3fmG8MKF9AdU0pnOfSvd904hRAp5HM97
0nooyZ20kqXP6NoErslI7qm8IWc66BMQmP1uHC6BAfF3kPQzDfPeTIDIryhrGYQw7HvOlQTe/PnA
byDo2wGlruOxUaL11fwjOtLFUn8wZZ4IX6bJcTvKMRieMUObi1pjn61mmxxbHKvZfgZbG0Zj/tjC
Q9B6z6C5QWHQTQi85/GiWkNirAr7NseTuV25+4DjnBbUg9eGy814JWFnKJPLjtcxjPKOsPGwY3qf
x8llbnxzhAuHtS/qsuTTw7f5lNZyoLaZZUaxFMwH32TGP1uTXqeWLO0n9pb1bZE/0Rq9lJcUca5c
ka56uw12dHCKVrHfw7I/FGQOexIjG/LdhYmfmR41opcaAWlhPmBKmZWGQDo86toPiagr5HZu7d20
fpCuiOGa4JcIFRmMKunvnFYA1X0hR9sxhRiwBpKcCYncXreM/GaTRY5ZUZLym4Mt2C/gkAS3lzve
LjDFS0WPzhyF268gEorUsYgDHV5ZAI+3S3GKVKUDzGL1M9etQJq7i3+bMOsBs/ak9WBKHU5vbimx
Rc1FueEIDaLiJkRkQDWiwhGMc/d8xNI558jkJarmjDVa2I+LZYCr1PZBvwY+bqWCMlQDUU+CgtZ1
5Fauk07LEji9JjNWCJOGkS7O/IK7GptDafUPCQntLR5IoACxYp/mqK7STWZPzeB4o+BlxbqYCIJX
jXIQVQd/SN3SY1kF6eSg+zeP6K//hFD5B8WWZUXLZadjndWthKz9n0gyDYHTesNolSPBUGIqsjIi
AoXurHHOjqar5HSgCL4D0hBX04+3wQDd/O/pD5alHLleiRHnXQCsR/eKRI4K1RHKb9JwRkfFbiD7
HHO273K0s/nJC4Y6UK9Hx+eUdgmigWaNRXFUZZY2VDtIK0CkpN6LtGmBI//CYy276Ec4Wv1KvwUd
xhTxC6XrEG9t9st74HLNsm+O4NIwR4uJUrpdT4DlHXL9bu6pDobhg9sRTQZmYLclEdFtIQrAqqwV
zCW0gvMsdl5ignsIEvyNJm30r80eOJpqlMLJE2hFd4s5iZm8nv5l2Q8KaTxfmoEvt16mTqlZY8gZ
Jm26PZaYYpgQN+d6OG83oDiMGcA5Nd3m2I8L64jRFjSdOH3/jgiEp4S0ltZ8ka/uxtl0Pom4EhQB
kPnTFmYtExpWyX7ZTjvxUjYWf/gNg82ccZDWd3wx7RS0pZOYtn0XVpBlasjV2yocCPwijvOv57K8
xGTdX0V4gPKgXGJagdJWZ7jbZRCWW7ZyCx8h5QKM0xHGCp3UURavnqkznq8vXJbAWtIyyiA+DdFU
sk0JIz7hwqffegLZtwEyxAJfYlLV5bg/7qGA84+IQN++32p8SUS//ZB0h0Oz7XsvCDg2qq6V2QHH
OUh9sPClmF+BAXVRyKIjhi+EvGvA/8G9b2XIx1ymjof1ObTXP1S9yNuDq1DTzLexLF5LHpcWkhnD
3EXxvtY588n9LoRpIQhBA6Y14g5t+nxxfmytQbJb7bmxp0f1iLT4Llrn+WSjQAjP9zHh9ZSm0P6a
LIHmkzZRkRMaIpxFBy5rvjXvSVsbLK5YmCAiUFy9ZiB94KLa8IPzTdwK4vxr8KoI71uDEntOvf9R
ukoJpK5uZWYgHXguz/JwPQsMjF6EUUGlRLpfkwEHbghHJ/T4ob6Ulo1ybUM7SqZmDGo8q+/NBaZU
as+I2TIHgD6t13+PjqhVlOW73HkMjrzVkSKstHUIZaJALgNUOg3EGETMxQApmlTHY6Un3bVxmYTi
5vqFsgAqED8/5InedTEx5Nw2HYueuftDaLqUoRf+8IYo4kLvSpUEXLcpuIicdSlMy0ljBjM3nQgG
spXdH+9C+S0sfpMjUwXa573jOrzx9Gsa+HFgy4mUKyoMWyXR32D+N0qFomJx8cULg0ypINC1HdUD
867NDPO2WPspvmKOb86YaughGz7Xz1xJGavgIhCtNM6Kp6nXMb5LN8HgMriDOPISAwiA2hBWUfoD
Fn9P6gT/mlK7NxcfRl3ntGxUn8UGsSbivgYtD7lS2o4Fl8by99E8nmmsoXT7A2kbqkJZuqpu+wcD
Do8qbpkhJQnnzbMMohupQ1CSjM2ad0tXwiiz/UTr2wLK7y3zZ8J77cGJyztcntt2ypReVbuQEi7q
KzXqTuxrCu9oYzBj4TuBxPBft59pjFBFOSh/EU1Ye3313eqMQPuf00HxAFSZqooR7Z5cXQEnKm3+
ys0kc2nUbyjbZPhtinobHzO2Y4DO/obIfKMQv13Gmr7KsNQ+V+Df3GuMlqbHaGoewJaWgaQBN6Qy
upXQVF4Y0G63ozaV4/gcfgTPvdCGV76+4No8ghuqhpEQ3SX2lOHLi1iKW7EfTRKIqfHFlQdKYXrc
GCWbrBcvjUbHuNSNV14DDSIQtNGpemy+hsuDBIP4EtrHp/TWrWKCL9Gw2Fr9ynxHEqZOCheAfy56
BSM7ni5UHjei4RMG3gIo4aj/+9rX5BAmjdpWR1KKyHHl0Mq54L3aQHwlDwsRIn5J7i+aYREVbKo8
VDnVH6+WWpnMGtWGUB0+vM9Vrd8h5UG9N1HTxhP63TR/O4HG2VOJJqxx94L6SAvOYktFC+66mtvp
UJcf139mNYD5Zje7uSSc+fX0PW+9R5Fi88KbJDO8zjatikYN/IVwhJygdDw2maKnkTnhTgxQKErL
JlaAfoi72lQaswGQex9IDbkhxdffBg9tYA4KcaVv04HcAtRLS/ryt3yQRcJkMYyDd+mf9ap0JXZl
hNHJpRgBder4CSp64NieBPral+dKoFwBQwp9CpT88ToaZavWi0atiCygMAs76TkSu3Pdd2k11pFY
ZFMyMkgv15C0/hOT5Hrdzg5VXhbhlyKNcbSfEY9rt4Wc7ZPNGKyYZ9eI+oC3UFxR4nWoVX+013YJ
HCWjRlsMnQ42scCt/mvDZ16mqNUaGpycYj3yJ4Nw+4mq5em/RIhxcyeLVamVfZmem7aU6nEBoWab
wWTWeNaV9yBf3Sd70F0c3aU9rMGMhRBN+PblNRCZGxZf/4vEjta9TkqfI+bv0pjCv9PTYEXTKyyn
FbbwzWTyJ736d235cZ+V3BJQ0ZCTJ9jNn7NvZKTHL6NIrVS0wRx+r0WYOX71pw30TqlreWM3N658
ezRvDBohJI8vxKYIz1W9bZnA8NTAqYrd/6EHPGdlQ8UDSxJpU6TjF2VtPE1VNQ5kANGfIXCSFn+g
A381e1G9oSXcTNyaEoMgB/A5lrblCEpqwRi5Q459/XDjt+K0oi4N67aSkJDD+G6gJAR2mZRp7nfX
k56xOxLLUfdd3+UX3qki693+8rTPwNIFAn7JCcudmJcosN3t49keiiHtVZyr1B+BFH9+HsrVlW17
mQgdV4E2k4lUxX9+4alpAqEElFgZJlE2BtikafdA5NXuX4LIdhtaRBQ0uen4wV5mLRqgQGlNIFMG
cWuOO+oh/EXE1kj+7112My2Zh+qvTxHxQf7SB4UIMchfO5RQNWvji+fSvIz4bOXs/wnrKFEjaY9L
RcIQcKGbvi+69Q58fn9DEuVt8L8YzAAIIaL3vRlIR3Euhoo8QCdTnV3K06MRUg0XMQIqbHcKGhUU
q2H0DuwrXoc7AkYdTMsNKyyrjz17GTon8SF8pNpb8rPubBPLWpGJS6/7PCCB9yINWCdQUCmFsz4q
ELcIy+WBZPShem0uebWuWlbalDr8oXGEhb3Ia6GiwIKGNSDULte/rf5e+HliwaCPjLeGkvtMXjJ0
koCVL7+7RXEZG4cXAsQAdoatKebQQ36nHvgEJk0yLMvyKwnRbaV6MN6rwfnr0QnzEanRVkqCxpy7
9tDTBfyoZ4mi9RO6u+RA6JIgTsAEKovPKHbp0NWrl9Rzm8UBOsohxYT83upHg8R0ErWfYZ7pLa2j
3s/aUQ3HLg/zIUPRYDKl9DfEtUyhYIYZdzxRbvWYhSu2x4XsMX0IJbIab54q6wEsRvOxHY4TvbRV
i3HJKj8W9N4jJLP/idbs0uccsZN0A4YhCvLDvd3kVS9Q0UmU3akAUx8es8ZAcwlrY8PcMBkjE1/4
H1LiNOgjQ/bWwZTJOOBdfp8JAo8kG++K0PIyTvYKjc2Qc7WxDvYC9txUXZsKtB1DGhhNrBjNfjNu
rs5yYImZOEEn5zBvcOcNjAjqVT4rUme3eIBP/mk3e+VndUKhf9mgWfLFJVDpihbq9oKNNph4pBS5
s/tg0t5mSyUsVakSzSYw81ALoWujv+WNCjyHoLs55m47d0C7EQ7Uqg3NunXoJMa4QtnMAg/8jE8o
+o5HkACv/DEPKSyG8GLS8JklMNOP8EqCQaOZGvn96D76Aq/2tiavUxmOJbyQFy96BQO9x5qIel2C
Xjho0RAmCjePBf0wf34xQM+zBveCVUyudiwWLTjLE7esiAa1tl5WENQ+3DSTT8a7KzFFViTKHDu0
rVeahOWsq7tsKsjhE2nam7Ff63ycQoAXpPqKtniHiaQxHKzI+rXDIESoF6AVFPul4zaBsqb1xp+E
Ud59+rmFHKXq7FJn6KEU23BOYkK9aW3HtxuaaroJ8ekAaxRQTNi6sKFPXE8cSW9ssPBtKXfC2mx0
z+pEJzVl0N8qi3OEZlixnRSADCjde8xY6lv+nzlIKdt3bUT5PzjZxMsDu5JVoPnK/YiDFVvYRgjX
0jif23goOq5v2n46he6wnXHQ43in6lFOlwXUZj2gnjaG+SmxA5udoKVaZ9GFvDCYXYHA6Os5G5u0
Icwf0pmOc3P2grXdkm1ZwdxKa8UI+j9pskHPnUlmoGlqx2lLkd5Rh6+a8Y/rYJFBet/tgba66Kej
l03QpeQ4C/f0XP31QHzKX8WIlM2aLxUb3Gu17og+HjMZJl8150cRdq0Z1Kym0Dm4BpUQlGG5xDgJ
5kICH3DEISxiF+gl0Si9NHfXBD1wKRKj6F05jEZ+y86GnmE9Y1IJVxmUvrYdQJz/1jiSD4DUfmS0
on8tV2Nx8qsLbC2QMT2DmnvQ2N3eGcpXm01XVn1U+nchms1knSW8YiSlDjom5idtVFzEWJiYEb4A
oO4SJe5KYPLZWYrYXyhvZFhjl3eFYUWHyhiOj6+K+jhHXovzKiN4F4RiF2F+1fpak7/gr89URLNU
lIKYm5yiEDs+xZdYBmiLL0qPtoxjwe/59+ar/7oxu0GRXC1IMv9wfQTrsMkPEFBQFx9kZfU/hmG5
ZYMhk9WXaJRKjZrAqPl5mTXYvi57MhA7YRnnMTKFMn/86NjhkOQJWpSslRiL9K4zV7xj61JRqdqC
rOkUSMfVUuUM9fMs/LjgU7P9RoH/2tnXIamY8h5yYYEAFzMRTnhTRV8VLfNOLxvsYZN0ccwbdlYq
tWpT+YBB8QxmtqezknqjPM1Rozn+BZFIc0KCGC5uwpcZbEAsfYX3RVDXBtGVFh7LPhnVjvUIUurj
RnBKwQQfV/AuS8DYFfKqg4ojKXtZTKpXTSwR2DQhRHDAsT19ORt9OpvaYoFRS8LVimrogSonXAFA
WP9r3fMbR+k3of7AUCYbcRmdAisP523Dcw6lejvTVRKzDH8FlnKEUcTAsdSr4zix0UaVp2z4aV4c
dB96bwxkAY+K2ayxhdJ3kBXdIcUJxIaiBT+augJn0DFsDc9SvDOCWDOTakEGdtq4aacX1AvCGUgh
UWI1ZeHdQfRnIFluhU57h+gcDoOcp8UTHe1FlEhuD5XYEijHB8G9nwFByf77gYEmm+MiRLzDVcnH
PdcX2vsAugrcWo4HEyNJP0zCI1MFuI7bRfx76WHWS64/eCToQhpWVyxNWN1ALPsU3b497e2/iJ6B
atrnJvmUM0Vq3y6HZBJlZeozlDRNAmjjwT/4iypn20G5keixfB+b8MbhQ7X6fBWzJU/Hmeb2Ul7g
vjh19bUHjdjchjOileFeI2bU1PHLh7O1iTOtjPSHEgCVOi9OaGJ12ESSwABlUEHxbPxwKEhIZO+C
a4GI/2RWpxWS4G1zpUQExfd/qlEgE28sa2YDeubMnRYT78Elt0sbVNi1sGF2R4QWQl3K2d1mEWIA
JNSBGn68+G5plYhv+15AQKsNdiZJoy2+s6g7SqRfBh9Ar+5z6oJYnkfRTCUPwgW1dy0Ctav2urju
1eHgRyD8snNbdpMk3/CCI5zJhjVSH9yKPRA7Day2VPq9GTufcjsDi31bMyhqi7lzhdsd5vW+PV++
1BBt5h+xMaPpgXWXe1znQolfOIMZjOlthpahuEnUWlZK3uaIUdLikXKqInoZdOgrZSqPe6rHEjZ8
KqUiTrnfBHQmrlaQc4zc9ZKDyMARoptDBLlLRMezXkq8R9P/GlTz41SBrQhL/MjUCfD92Yl2/Gin
xZMO1X0j6aqSycyvRh2CkIpl0ugITvl2Rs967+7dBniMwC5pv9vK77mEl8b+483wFERVQJJZY+JX
uM0KTwe7sMdLqg4JBIJwmoUwsnN6LYrmyTOt1EdRfBKio5BvKGpgfuCy649S8bflkIVVlJ9TuuzN
L1sGFNMn1zTZ7Q2qh1sZcPtGQajEaMWJmN9NNYLswlAV6KZF0uskHWbgfiFJjHTapzrtsyldMRqW
IFWyjayz9p1Jv5tj8ndDRxthdORC2yrmqOsr+DRMfjKga9vYV9txpS11X1kXX0PC3bSiye56qXmo
z+psdKVuGMO3yd/0Rt5F8JKiQ8wfWT5u3dsGdMpSKOM90jiAfDe2p6y9RFgtkVcBPA22rHywFa/e
LWUA0zUmu4QvB3sGhKpOVQVKWnlnZHhDvifgeI0SGt/c+7IJ+bWq+CMCJeVnfAPntUhvzpbM2FKR
DWApsQTmw8U6zK0U446pJrYwLPNRtH8KIu1cGcCwxPuUaFj4CdmaEYfIvb4AXVlOdGT5KXVZRa8O
lPTy/rOAT0dI7o6qc8YEM7gWocKduJwZ2F29yzcJjRk1G/mscKiiSdy3Ntz/ThAbAA7PT6+zndLn
LefOAMvXZ1qrdWY+XfH7M4TVtD3eA6WD0vtUaly6BGUeLad7hHzla9zOvIM9xoSPjUgNYUNb3Pf1
Ds3KbHNKYoPre8Nnqg+Gvz8443y2PDC+uISDj/2EFlnCBDKbzRMY1a4LgfPmON2Y8i5AtVvsJdPT
y6LET5BhMfh8+6kLQRtMU2hl4uZm0BXeorUwBZMbozvNMF7pFEJVyo8yQfru0PjjsZ9ctXwoyH84
BO9Jv+3pjcDfYerlxVSn60e3MErPgFk8XUypT//osmApRC9nOr4Mn+b2J5RlfiwcC110cXnftZWN
micBbl0P58rZfeR8aIXYw8qEYUAXdzF0RsR7LIjZEGmKgDomLUtNoqPIbtOgImw5f2dNL6A05GLt
qDFKW4Hp7uM6qqYvVtMHxjYvEXjYPskW/8CGYOgxu++46Xm0mBRNOdoIHHF5oNbyONqSQ7Dit13o
RcnauewugADADnC/Bxrb4gVy94QX7lTVaUImFBM6tFxL1Gpjyzz3lSl+cyZ0tDIyWCB9i7XHTQ3/
WjbxM2wJtzVqfxuN55lKPUSnHIv8lT6/kFCW0KnhJvvKh7LjVNJXXWc5AHU8qJrT8p37yDBaXEFq
m32WSF1p4qUf83hN+OGS9AjzDd0WSJvaoJxVPy3hQBjQU9AFDcd09jDkWeka27X+ddkUhFfnwMC6
vUyZoyxqE/nHJjK5vGOyXZEZLwmwwISbcNbGdwi4EuAd/b+L+tmuC0RsMkdbSypqxdl++iFz1TLQ
Uu0r8Y3vOoMoeWV69vaGuq4lW4TCELHolw3u5U1kmPK/ewz/jq3oaG8ShMdUGqOysZ9RqpJxXc9i
L6BozG2xy7e+imKgKjYi7V43ax0DZdd6J6uWLIkLiVM3WxMkBIUm/lnaHYUKug7BdEZKc/8f8hZ2
dX2aW1561MLZ3dE62Mur0/x7C7R5piVE9HYT/2K5Y+Ft6w+KP2sD2qqWaEV6FmrZE32GbdGNbssP
u6wIgVY5fHZ+Cdb11JOLVosuDKVytQ5C1++NDV5dxy6LORSUJszVcChJd4TRZxwVJLU/Kw3Aw7aw
4v78FnQvMR8c3ZUtp7V1wg4D0J0izfrIzmo0JtK6dq/timyrcbdqDUxe7bzRVIw1+G/pTEteQshL
fGfzpl3fyfeGkeyju2OJ+DmQ5J3/UIxdXiO/5k2NA4flE8Ip6QLxbcmzw2gwKOJdRkFDNBA9ikRT
IoQecKgcZ8F7LXiPRH7nB1hbnzvzlUucD/EljaZbOdfIA+diTm0kjrIc5+//+h9fOD/BqancEWU0
wxILy51AKQxqcVbiJ7G9VtqTeTdBf356KQHkL/9bHRezJxRsFp9VE+YUe+J3XfYX54z56ZaTN/xH
Cluel+jEYWElskjOeeVUaHsBH9JX5GW6zwsT1yQRXCAH/iI5TuFULb0Yznti948emjXwuNgz4AFN
UI95x977CWGcqsklwj4tTPDNOOgT3wgpHRslFiaqdRMBuKbFQnZi+bqHoYwErEOpBpCXDygLUxQ4
6f3+ECJzwZcMd24ONdw/8O0rzMMsEopk9+/t5odzfsGW6pZ5M/cKWeUh40mpvseM+3Xh0reYpT2r
UQZX9+KDOKt7IRaecUZ/3PqZkyLJidNUZJaRnZ/078Za3TaxR583YUBRg1f5zIdIGrB7pDFBOF7l
LUyHKqA+kIVNOkbtVTNx7dbvyL7JIYYqI2dzF+N5UCgxVSPzVe4Jp0c078yHmUE1yVzml5rG/Qhm
9Wmn6SRYDfYRG7ux52CG0vd5G27Mzx05hg3OtEVkGFL8cNsr3acIEjparmuAq2skZdQX6bG5uPvW
uHour2oe7oumlArZTgd5LxFB0MP97u32ZhP/FMxH/DEeUG25hUEmH7N18LXwStCjzu5OB99IH544
q+GzWC9toJ/R6sRmys3qHz3qMVTw+/0iLmxOyK6H/WsL7uOt+cTwNT2m1+9F9mTjQWufyd9x0Ao/
mvducz0tS7TinIDnWHtPF5OWqptgLwpNaIqwctehngzGt5E2X8y018ePHqyEB+IlbwBZPDT/M3rn
Ju3VvwKYzu+/ubevfj1ngxOlMi+J/wvH/+kEjZ/mhuxz5No0E8wI8txDJJlqb2Ty44rTg70B5zda
+QEBLqoFa6JLnNfsPbLwGGtedP1QPockQP7rw0CXtjDHwF4B54s0Fk32UAD6dp5/xvL4dIL5yybS
W3cxoAlqwubUXjql0qR1MYuL2bBY+po9Rm/KoqVcoDiOKcluSKmgaMoJrZmBcS5zM+kSUS7fQ8yk
pi9RPKFvTmrEBo40cCZO4KG7aMzvmIhIpXNZ6d6xNYiudheUwAi1qjIKF2ISYZL2ERu9HW9BMoRu
1Mh7crwXGT5Rl5QmYseY3J78lLrm/xtY5fyqr4g7FOYYYT0zNj5N4htBRAMOYw1fnvTymY6A1rK8
68qYJpZXoOkTWDx4fEbs32dWFtjZh3I4VUTg9WdOpvCkCypyHcgya1a9liXjk+LbcPB1iTeafDCY
ivArSYZCQUh/FmWhMtctNFgHtvGSwXfQ22PB+M4DwLwt7D3DhDO4C/SVQKpiu6hWONE5FsY7eOuH
naUB7MbJFs4Hh3oZkOb+Mdg5N79okyrjDNhpN7i4OS5fN4kiNeiPaP/TuRxmjxhslSnHhMAruRrd
nCpzW6jt9FQaAeCrudwK2Rq7EPBIAdVUHpT91lZRmzAxtgBV5jQNvAp9LOF7zvPRuUTPhyVGl4cF
v7iEWqgatW3EhtBxDae7B1EsXbmLeeZXx9/5DylP/EzgxUiyiEyZ8OnbuGf/HkKEj4J4Xbv8T6rc
TiwowwLzyoPujX4dI9oaNmRgQisQQb18Yugz7dHMnuLG8QQkI3gPv+MXG2B9vb2y8gOxCrndyBdI
GM/9BRAEjnOieVyYe5/w/3FY94o3XYAOqZwhwwp191HwVonP4eyWu6FUTM2reV2RLK9Q+dFAd5RD
9b28qjGBdhkrtEUU1MkM27qjyBacG8s2ZE9Uux0s+eKovKHQ9kOfaiP5PhzLqxpprBUwpST3plSM
wCZIDtJBfeMz60SjjZ/EXEgVBj17lQJ1ct6yUBLKg34MKkTDnc8AsoHNZZNHnHVVjd9lnKaH+j1x
HCG2VJs41/gtWBlk91M+dV4U4KEo3hTS7rOoejeVve0fYNyShMG0bwtkfLPvfg/pCfp4NrauxlTG
bEBwXxiqxqJRs/1gKta+b3Ulicee2wUhL8qgVpRDVRTn/3A/3A44K33RwCvcYIz1APuRLvPkbiGy
iP9zpUcSRAXx6rIpFQU3DUabFa47b1PrxFbY+vr4tRCHnZVrJp8cH7uwU+i7oxABx9i4wkenKkq9
Uv5TepwuUjrieYefIqjtHiXhk2paqpFtmNLR1kGI8pB3xh7HzwLAhLwzZcL4hl7tDgUJ+owxsk/a
tuQwA6l9a3RGeDMMO4TFBod610iqwyWF0YXM1VB7ee+jdylcH9PviXz0kvJTwub0c/jyqvT3AGC+
FWAUEjE+UyosfEJ7XHUBOiUEYkBpaFObpFsWRsdaue2e/RO2ogOLHvad+iPfPbJVdYAnN7rJ4VI1
uHKdT6BID+HyDTMNnr8VOhL8sI4W2uzS8QT+EBtwW7+umLDZqea3BzWFvboCMMfizSmybysdsHcd
6phRjHqzIecCMAeISdPDfsxkfPi7q4Kp1rCoW7GNKZBWzJk7O1CZPjPUVxWvBapBKH7KNTGLIGf7
OGTRl0KdvPdeRzuK81bRMfqnaw9Rcok9lXCZlLHwjC1ulLefTdgcwjYH24DIpqpyc7VOf9LMhdBJ
uu/aRDmoImP1YS9nBZ47GPeI9e0MMWZP26nPUvYPYx2R2/iPkkr2mhpnj/WMMJ70jiz9kESMzq6M
hFDk0XXF9oynpXuHjVHV3AMnN6OjGsm+bRiKysYUrPPk0TwxlLgk6dppeHwqycb4hliDL9TTyewc
gYOwqNPC+aU3/eWmSI8zslN3/9yCoE9GHsgsTp7RNpOn0Y201Q8aPJ/AKbJ9VvEw8gzkeJd6oxi4
Ba0WeASIpXSW/zImhgpiZkmHKTe7NtbeFnghsjm4lRLIt5UNWB1r2bobarPm9CLoHo1SEmH3wLTf
THhaEnXa3ruUArVEgqn09J0SGEFqNVUzoWP/cPMjpXdkMWHhQbF5HwtlJWksYXroUgl//PnWlcd8
S8NF0YAWGzYs2Dnzbt9VZlGxEaVQ+ocEyLy7qCk3Rmtr9ubFUusTMjzXbtW3DvBIhYNv1cDn2syh
+CZXX5Z5NgLbEWDiKvrUkwZhrUL3Uzt0m46taR+B60j+9EbWIEsDIJCCsg36jJoXi3nWjG3Dh5t6
nHHB93r4drj0kWd/VWNuZmdSzmZBG7/vwDTKSOf4wUo8HHfo2WhMwzTM/AKMxGO/4ywe88Tv4+wh
l6y2RfC/E17wumqErLBMHsZhfWJ/EARB/9ZFvdsOfIthxLfCSBXx1EsgCSet7711sGCYaappnD4x
9pzUaNDPbPQZvCdyTp6NNx2XPXa3Rk7MpClggfQNo2XwFjYFp8p+nm43skckMcVw/aXcW1nT/s3i
IGC1CNbjUa/7mG7CRWxE8BhI1PV8e31JD0BFPApD6BRdpw5PSp3arRvEtauv/1Wbu0hMVEve3xNw
zpb1L7nH8rt9FufnB+y3H5DxsXKBywiX+bwH4C8Vk2Z+jkWj1eQV71pTvSk+UdkmGzpoXYPGzdoH
fvlxqk92pyrC3/Tp4qQGljEOAiCcjXC6LJo1kjCXEVYJ/rVHBm2iOp1ciN9I0MJy3yz2VimrrFfx
HgBP9cLZL800PIitnAnnOhGn1lVAQyZM0OHY0+GqpFnl0ev3EI/byvbxgoKNUDSri0Lqn1GR6ksg
7Y/VpsDc21B6MRQRJ5UL7PoIJMaekSYO47H3KwA/fvQJgfcVNrGxjf+eVDQjNFLFxpMsW8vIO5pD
ieZO7zizIOWG1pUowGwzXWDTK4XRVj5gGhEcMNp4OUnflVopmsIkY6jkbdHkDMXajuzJEdJ+6nXE
MUrMGsEv5eHKsv/xbzUvsVZ0PC15KB9rnIkZwLHQMsz73MQNKFsU+lyDJY2Mf4bGVA49YO6ssXXH
OFjJHwbK5XIRvcQlJ97EXTIrU6gdVb2Nb9YGfPpI0uqTPx6uWVP+weAA+qTV50vIYRmJ/9OUF9+C
+HhORADW32vpgAac8/E2ZLS87fWefLlApWuocqlfHeSJ0R5b60dW4PXzy4NxLYpn66Eku2tK97HJ
uH/7FQPr3/7CXpo79pDpXt9OavbjXDSlhF3ndyTqsZQr/u8KTLPRLtUo5Qtk2CjTGSuFSOpNr1lZ
T25QRapM8C0EWY8OWvlPQz6p/NHvrcLvLTxz12meyxlc3PgJbPf2jwj4OWMV2madMqpE9UGHzV8N
X4eY5rH4cIKX/u5wtfX1+jUUNPnc5MGwYTipyfRgPPcw9IcfCvp/pHtZmGZxNFTWMRK8XpJQf/uP
CWL+abIwBBIEBuX2K9/dPFHcWYwgRmnZ/KBoI7lMDq7MiN1xDWuMxb+oyWZr9tE89xY4oMSK3P9y
UO03QLNg3FP4m4XynGyEylZcL1rFr9nP8vhxUL3vGq8Im/P+UY9ULCKmeaLWKThR7LUiEyjNRbGZ
X3AVT1lWevEyv2cDvpDp4+R6UmB3t6NB2/kEbODIbfal44OJmQGw/ped18Y4NbhfZ1sfTAbhVDzg
F+6F6tS4FGkfChYWTWhTh0dP88Go+cDsfDrtJsDVbASMhsRUhCEt9lSOztLzLYwT+p0Mplkr7DsS
JX/Irf0podeYg3XLVrhCi6Mah2RoPDwPOrPOJHj2TkoWXkixTFgu9txMJc+0TqbMINmK9xzun/7N
t+yC02IM0Uib/X4UwofxX7B1Yeklo2479is5xyBect8qbLjbfWqVnxTphIh5lebz2UEoWjB+liyB
L0hyuo8vFH27IRTBAWcX6b5V1voJQ9rA5n3DxMwHTbBPKUxzaRxkEs0SFs6V/NBPiMYPSl7p7eXe
2ZslIvAaKhWp58JeE8EWlTuyReWWGXXt1Yi1TGy0dpi7E3HVgThuPFEAd0rfD1Dt9AmdNmQontL3
5Ozep38Xuvcv4Mxg5Z1pWo+Wg9zxLd+mznN5FEYt0PKbzLTY64TbsDZm+r/myUrmsUb5y9FVKLoe
NquC/XXvqf6Jj/FELZgO/5ti9EZe27BTuc/7srAgDXip7XBPUf739k3lUD9P1/cOtPTHqJH1cnOJ
+ACJ0APUIGIO5FYCxF/RC54syV9E1d1NWMW9ysUpCgDBW1pEe3hG+1v0G6FXiFsMyGtej1OKAZng
1UMVCf1DAlJKTx6HS9LpNQsbW7V1tav816b/Wf/IjKW/FwdYQh+61Fz2/tvIyjPaCYPiAmls4rJT
JFDh+hzLrFM8lMYu4m3UYxwMRKMejP2Yi7/DBdSiwJL3c6tmjOpdzX04S7nJ8ras4n0Aa2JFTKe+
Pymr49N13d8K9vjKq5pJWCuak1KK3vHXBaPE9yO7a20cmJjmEgQaV89hgaCGsGNXOPcgtOgMcZOB
3WhJxmbpaXEYwZISBKPVR6nJyXXt4PEz+YP00lxWWeGpZ7RiY5hkuZhXQ7w7XeAOE1JsMcP/BH09
RfDvkpiYbnVqUuUSmieamMBKJYoiyAPjmJ3SsYxoCcc9NHI9FqFdxgrJ8dgevc1D/pObM1RShZBr
bky4R05CeOD4TOvTD//hCqjZ8zP3x2tJX4LVIsC3I4oScOS1U0/WnEKbRtJovcGvJDLHWW4zAGN2
Ngl/UcC997w+T9ib3sxQ97l5L5g61hEcb4KY2hgioEpSFQDZ9sqT2YZ7g58wxyVk/aqloMSueNHC
h3C3915yDDkf04cdhXjBeVjy+uWD4w2kdFvClDsx52o/3CIwdKSMTpazwWuqwtoMkvSTE+H93zi7
DKzLbF9MuL97cRSlicah5Ycsb1G0HnoTaSfNAGadLxhof9WM8R6NDFrLWESyKo1zcMCSfJbl+OGU
i0j5cK8E8ycp4NANetN6Hu7n+44wS3R8slXukTnoBq9+qdwCg76rk9FS23mG6axv1aKPrx/RsO8Z
ivbgKApjky3vUsev8quMDSkS9BU/d9BcLcCY+mXc12t6HPb+/PZiHKToJPGq2Vq4qrEOm/ouWFXT
d/BYDWEGIJS8Zp/a9l2lesr6MDRod/5KAiAXx0kp3KUuBj8uV8nOCZl+3nD1fBk/5EkeALaTGFaA
/NSMPjoNKIA9fUo3YI9UEQpQBSszKl755KHEKO55IbDwlHBzWaKCMe343ExbpzcjirFIi8pne0bN
b39CK1ityvnZUSK2icTs7YXTW5Sm1rGiZUfTw8iI+wENYqrNwSIiv/eWAZaoOmJ17lGCRmTVG3bc
5tysK8nV03JazTVKnFSryhNeUAtJXCkmeOtYSMdMo4gGh5LGaH2irEl17todQ7pIqimMi40G3QSa
DqSOAZXWuy1lo0xTeTbXO5RbmlLyD9Fa+rNl3eHDfAqEwnCmNOAdSQBc2rvAFyexi+R0jx+uqfux
i3eSyBuZWxfELFyp47XR/9ASQ8xu2trM4MmVHPUFSs3HbzLfKjSuW1FchtoIjtH8y7YQZf1XlR5t
nt3U9YWJLSOsyKwPOZkrlAqvg7t1lc+sF87/6RehQ4cfb8qrp4I0UdoTD1Dx9T1kHP0MT0FYt/2N
afUIx2tdzxfX3GLa1B3gDAe3Ay16QWTjUqnoLqCnL7NQLTDH7FRTsEfFr5Xg4FKiPsnNaSblWKlr
Hr/NQjhk7aUW5gMHWrpbdY3gm7U9OjRXWb7MDMq/obigRQsjlCwWGotABuq4mLpaPdBj+e85Ms5w
aJwMVn29PLQQp9AFhBzCU3KP12/RJiEsrw1/C7KQuqDOvxPRPIOKLmW836jWaznrk8EjyQDohmSH
MZbHbu7sE5AbIFZviFzSO1eHoQFC7fZ0h0HgrjFIolZzWtW7RCChr8PJz6p83BAxqRlCrg0OPj8o
9hqWP2PtqrrE9EVFgVRBDvjZ9qIIDElK+IVya0m57Q+rzVvv6Q0WY0sDx8qaeNZKVIX2ldY8JpYX
yXPxt8xEouRJwhniSB2TCPHS9SkVn8BqM2xWMAltTC0CKxcMEbxwbz6J7GMGn/bi06bmhmTumPMV
xzWKJ6THgLdIjDegAzzC1L9wHD6CCY1qeDv5BWTrkELhf6y5ttatVcFWT7YhtxkucfBEI0VnMvhf
vtBXluf9b2OUV0lrgvyR9T0D7m0qsF3m5MldorawSmu9DFYHY0nweVf0a4JoNOKQLJ6zy7YqmUbR
Hk0eKtXe5/AcV2ychKAXjVjH2dVsEiiz9ZIx6KCkQ7BEUh50+08Fm3v389SAcu1dbSVEgDPlOIss
HFVsIBUMdOuQhn6MLERZiBceIvUyQa1gi1K6dfeI7cxQ4WlXJ3VohfyxgleaGok3A6MW8ga5HljM
z/WKvT7QMdNb+ROBZROSAK6c+DtaoBsygVH8j14g6UGPzfy+5WzNuzzWCflK/eEAI7SiKyFSNNOy
zG3MFv51zDKtETMfL8rKc4BlEDwwD5XWZqKEjVyReHToUqIvF1benZAAg8WhQORex+BH6A+DCl9W
kt4YyXWUF99PCdfrAFoueb9xphBw04BSx8fmR5YZZePN2bvYN2ZE44sKKxVNKcRUpDLQ6h3Iwym+
29vtiabpHovSnBT2AS9GvqcWEYB7uFwgq3X9OHGDveWXTLXCQwrC/jcAfEoMSZQIsuX3FIfLIsA3
MI729acCBgrk6QEqA4B6eFNSGimKyl2N+O6poP9GcZtaOW9NV5cwLin6H4sb+Ri3KVTCHWbAqnW2
YBTInY8nuGJUYMDel4noz4BYe3TQY1PXluc1feqQTgUM2oMvgfeVLKOugDLD5muOxO8lRIYSLM9N
Hf332vjeXVnSg3YZk+nPNfzxBWLsd/d0Yf+pTuyAkeqIEhDOi1yJtAwc38zni6dKkA6DyAQuK8Xg
HUCAhUBRhGXTWiwyIInusEB01lX10Gx6elxWDPfHX0FVdVlR8eLDyznCIet02Ny8mmqbUgidoqQZ
NO+jNDDZI/j8ebAiulJjOqJFN4uPFLi8oefym4SIq3Ue1Udgig6z+nWHFwSwtZ4Gme3gSpvWz3sm
Svs3Zc6hBe9JqQd1k6AS4WGdp2eLTC195T+usIrVZDL825IkL9jbt/wKakx3QUjh+f881hg62hs7
PY4Y45z80MDYDK28Ms7ZTILO9CBZtUnDWo++YX0INa/SwFykzeOoDj/C8hqnIatKlHgm4LANhYtR
QbJLNm2oz2EYcnbDufxBXl2H3eP83mf6aRz1RM8zA+uCFzTQgIq7qlrmly7krExcce0mfIQvegWw
NWfgCMdycE1emLMjP6V3c/KWzhr4+OhqVIQaMU3SEIQ9jOmyPkrpn3E2w+iEKr8oFWI48OvPVNfE
s77LFCqDUfugYS3/o+bU0oe6whkvBxtTcObPY2kesOa7zocka7TNHTrVLb2gjiRorWYA4vJRdvii
UgKPZ9Q8W9Ojsxp4h/V7iYltp0Dd7nDVHZjGeBmlpYa8LLAQ6AHkDPc6Ek6+OeGTb2HQ1S3y0LTc
lnrTKdmFpaZPpS81L4230IxSJUul12KX8Nz/9aOoCgFOgT6ZzFsz8JtBIZ3cgCOF1JH6Aquzs356
eMvV+f38S5WxWB9YKCAeqcZ3Kxi0YS6ge9XQCvBElXpl6OeTbliZKomFGkLN/fysmN9srhRUFXnO
CI2RJ4b6u/HVDhCVkITHPgceGjnOMweDRlbM3Zo5LKOuT8nH3hksp52mnFIj/GYif0GxRARObzxo
JqeP/EIV+w7OaVtqHjBXtPH6BrbiL2brwV6OnTON5wLIaGZWa+BPXM0dXZU7qdx5Ze3YpFPA5j9B
lnviAa60ePBaREmiFcjAhPtSiXQEphi3hcOUGJADefdBfVXwZs2mcQrriP5ITo/byLBK0vn9DSCk
XbVs8IOU8iHtT8pU+40Ho5E4UGCHNDAl4wlQJ3UJrYAkXIR9+ERkrd3NvqZdN5Nn+Jf0KKXKYwRL
m6p8gDemORSXum79Lk+Q+qNuBVPCj1iZif6xpo5S40KH4CVq+QcYy7SHnG3trG6pAobKic9sGvtZ
yyYznkfKTUV4sQHlAlUwVygyrMKFcIEI3XPrn4Qa9gx94SCTfpZ8qwxqYMGEFsBPiKS2/8KvGr3R
2CEjdxRYBR2HOiJGfm1sFwWmibfcHd3e+OVaBGRGJj8BuFaGA9mc3UZdy/Dnnb4RtUFH0+Nhvb9H
XrKM3EXDtPpf/HjCBhAtGclUmntqLTVdxQItzE6JTcbR9wgHzl8jCPcjUh94iUuxcwVCO44qnOth
38WqPEu4NOXyJQeRMVHRtuYM2nfiXDpWS2v3F9uPNoSD9SH3sWk6Q/R6mQzSXCtCnOm5r4RnZVP7
45N0FIR3d3td9TyzNZnO8YmhklcquyEEuWRS08bfBYpOO/oxaEMzWK4Hz0/X3rnobUgx6HazjXQC
2f8TF6v1KytomBS+UteQTco6hgbC9FPg8akber+XXSzmwQoU2Z4wxIL9vix375P5tID5czem+ORo
vj7AU4xkJz3n0NMrG56kNdEu3k5LXFYc/xHnbtAtUJPIAoVnEDpuf8SZZX9Tm757d/WIm+pLRSTw
Ou4M3Rq25wsXyL0k/mr/cHjmXmVc84O4C9uxvcb5oAjaK+Dev7IS8g5hC67wv4rpgtI/RY9UeXLE
zLILHQMJ6I/kaQwkd4nLtuYEPkAumjPSBVTj/e2uYl0fM+XyGk1Sy0cvfmmbxv/CFZFn8nQmJJJv
m6t8yj512LxCjkj7w71xSAtvj91xg5KIlEM/uS5ayWKAnCBxEaR+NSORR0uYfIzWpPntm7MYuMQn
qLOyFK/PamCHgzbRm6ard4viAkFTvXApZ6y1u+fExmYUPcOnmxlJ31MezJryMzhr0WQd2/qBWVkk
Bbh0HkGPvamZl6SgST+YwBN9FQU2QOfSFOZeB3tFTb9fp+DmWExzvwbbKQzK35gtLkJzN+FWflZl
pkOGu8RnY3iQmH7T5lLhPCQEWADNWRcLdRV2dKunLGIJ6Wt9EAclzjqPgHzJzNYpf8ATDGEwgmMV
qmH9m9iIQJgaWAARk6DJiYMeheKJqAT2W8nmvpENp6tKJRYN8eReCVVvI2i1TlEnJfu1nVusytKK
xFPf4eaYT4tegsaEmr12M8UxD7XfZJL4GHa8xd5pjq154wZbqk3Tgml9Lflls3Wic0XVym2SAdLv
0rv0Yyc+g4eSGyJ7kCr9qsWbPgYNQXFbrJKHjr63fRNYUZdG96bh10jXDtoeFFlEr636/mJ+7wVP
9GjyBiz0xz5+VyMu8SIshIh8LzOj9l/X9Dp9msmqc0ZsdnucBaydTDS8yC3RhTnoj9bGnZxSd1NG
Gm1HZfXPKpDazVfX+/QHTwoOkurHgCLrwFfhvG8xCUMLsdfSxkSb2Ee00A7e0l9HfBD38sLbSOj/
Mg4om990W0a/XelQT2OhjfxnMMmYJmzID88KRwj6X02zJovqkhFTdKGekVpPv30AoaRFqQMVI0At
f5LBll/vR6bHcMTEWqyd1akGb8eHDiMS81b4miDAuCcaGd43OjNubEOowtbz/QscgCketknEaZUx
nlu6Wm48T/fwB7646EVvf6Ynph/i9oJSiF3DiUgCqkH2orpz/t6m0SnkZSU5uxYGqxKS3zlO0uL/
Y1xO/t1FtAhegtz5SFywahlzXLDCG+OYiQFqiDRBWT1iXXqSosAz9GdRLtXOA880jEvuXPzRGaeI
sN1m56lgrbZVwYgf2a8T8o6SpvxDumuhkOsrbOjYlLKvfh/IYjGQCapHJYTtTkMdx7+RQVTRuMrk
JQvo9TucvV5KNgM8k4TzIvp5JqorTaPoCMJiRnQjSsm3WO/QO9/uumQl4GbyXC2UQRPmAhRniGKC
0j3PpjapNV+Ng3tUzomu7fuGpu/ncXsJZJKbtc8CYRKdej7ZYVSe+eRkI/xPKYlxuR/wDYiFNHVD
KB9hubLrAWWxOIPK01E8L3FPnMFvwe5E4piG/1W92a5ZFKakJneuhUsgk65ZwcdSZmFMJwtfvQW8
GUCauKxdia8nN/ol3XxBh8yLrKsZGG1wsyUMy8Nxl9AupgFE1GbQn2qcXK8jV0Kry1EG2SxqNvwq
3JnxbThBNflc9Sh+11deSVvA+9DtgqKovXygCOeeYTa3RzMADM5wypd8IKpi86dhUVIXDQhvvGWB
mAXH55Pqc9Zz8lL2SQ+KZGzAYIxRzgs/zOg6bJcgN9rkTQw3GQgDo44tLKsuDoyd2BtVyrU8mXkz
vGxNDeTETKxhp5lzWHQkFRa6eUM+BM9Ft0GD8TUBH4cOUKoN9MGw799v0Ekrfk6KGrS8ehy7IIq2
pPjR4OY9/Q20pLneaP1VefbZFjarYdmDz2X8wFw9gQr5tCVYSeN8o9tHg6c9r03YTrMaKssGj7je
SDJRnKevARgLiUzPq35ekxZVlFu83SSYCsoqT1mf+S9BgxcuHc8A2wvITXVSDgv4MLvwOi6j4Ylo
mWfazBETpZoeJT7JTdQLqk+nmGHNCRaJPo71q3IS4KlmoqK8dOVA8cbYRjP53Tcd+SkNl77Ftuo1
ALRNyGLEgMvv1pYPdN6md+SNkNPt+eL5aupzhWHU6BH1Ki0qqez4aV6kvjmqH+fSerOORu2X0ZBe
8/TRj0kAXhQkBYRBmQH3oUg8hE6VJFOCyOEGA+vrzK3I6+3oj5g3NtOYRWTxtqbcmg4m6H7sB+t5
eqeC+mpTwSn/hxSxScl58Ag4wGTytB91+RFY/94rtRG4pGaEnkLa8wKohKlp6UbM9CqVPwzI/QTQ
WC+BmEZLALDnW7Ca4vi+7XITsQqh4z03rO4tS5qb060jH62Bx2zqpj2b+ljZCOXwFeVqGXLyJQJO
ZNOnkUSZRVzPTSiklzgnsr5HF2HFlrHR0vovA6uMyXF+vs4RPXyzfu/VDD0Fg0k2nA8af2aNnT8E
avaTeo30BwT9Ce+qSndTfjpJC8TQxqfz6w+Zc26nZ0pFFqC6e6Rgez91vrqI3rkO6AHBQDfKlJWd
HNEY4K1LFfquOET3kx7ZqVZnpDCHnEoeNNiGpSEPuliqmvUbj72nSt78gEctGw93rOFPrV8c5ynk
gE4IPBBaUjz6N0eghW7J2KBg/SrHFngwLAQexJlW4MK8vnNal207spRzCjIFNS/Ep+a8jAdp3d2q
uRDqftIsk7JJ/4PDme/uEWM4NGK0w94gLlsrmoNt8gdOazABhAOSiUN3cyf99bxO8m7iuL6Az9TC
cUgiTMVDWRqRYWwn0AsQAcrpf3EPrMgClvavg93emFTOlDW+D6/niVDjGtvhBepn92ZCnc0rVN5c
JW/B5rA6Mw/I5fGKN0gW7p20BaWzeQQFgjg8eC4BptxStJCAhHmzK7yA4p2Xxk+8vtX6/G8Tf0Pn
yHhDdcqVo7HOFvaJFFehIg7eCiocULsKn0ZfTV5OyEL4fZrbJed5avwNDSnfIxaXvpysCEI6xPFA
qDfb3l7vs7txqjgn5u3voTZdkHWdHesSAtd1Cik5lhAQCNwv2Ln6KLFN5C8X4dEyFyyc0aD4z2d8
po4+37EfKS2bVv9QKobuARqPQUQ7jG+2oqTH+ouz2YMyx1Hs8TJ98rGkFaxMe9Bo+lRRjv5Ba8N9
DKGHsxof+soWcOyu2tAErYmUOfx251chTZFupcbKzcLPaPzhy7DmUwJuPmivirNwf86AdWnlCEnY
zpwEdkAYmI2gbgvqrQS2dZ34LXi3NgvLSsG1/WAM/mkLOhgWhStFhB8GG3RZVqTGx6rNNtMHkFgB
fhEk49zIbEjv8zhj039MjYlXB3Rl7i10VCstiNzEYZ4V8H3WP3/QkmmZpprty9j1GIbMVqWxWakP
7QouhPNlQ01+Oxtp/7Gp8Cvc+5COEbjMlRV5yWpJeZrrLn41COT4DFLhpvv93RoCYFYA7yRTUKiZ
S8dD6J8WKKzZu6AaCd9G+BtJ4kPaAtZAAMZMY4/k9dvfYPo/zOnOoiHgfBENIlY4D8cgvYhDJ5EZ
DmpMn5Y0KKoUFJCGcc+h7mF80pwwiMb257iGCQl/2hqfQMXZcFaGL6FOrN2RCaG6lfLfjpcjLkBD
iFYeGgs9Ox2AWTLs+D7O14ZQBNV3vAWRArb8g/QAugXGfkntkabmYEuj5WuPN52IbgmCE6c8pITG
pJ6mgpT6gTqo/J73MoVdh+TfXgdij70mThCdYVt5NXS/dV4JnJmEk/PGstec4PFDWKay2YaaJ5LK
7/8D7GX/o63R0hxR7u9s0JcJx2om8fyTCBZn14valTA+18G6XJhkcfoLy2IgYPvKAUvYTwpJkcNM
lI8cARFiofDoL7VOlg4cdTcb0eWNFrO0e31QB/Dk3SNu09lXzvvTWDayuEWfgDWpa+FXnOIWhR+h
ynys6fWtStJHsRwEIqxjJpmNyJQJBvDXYkiAGlVad9XFbScdojlotU6j4HcWVhC8mder86Gc/jas
xJg/74JIsfZfH65Nj+tCB4QJayyznV2Q5sALL3J8PV3Z9FdNwPtjvqHbwczs4fdDyOpiaVDQ+KyJ
qG4d/r+gdAdA2eLxT8fzbPrDyIZJhBvtW09fl7S9QarD9D3dbMsIFaddm5xXXQdjsVhWoUtsgbuC
cw/CDLmSkmmRFLpeQcpGMOrhzmJbbIf++4kwYVwx4k62y9x9WKs+GUvrnQxCuF798sL5Kh+K/Hqg
mhBIEZt6nQbOkusAGqmv831pTc3VnWlXSj6lc7oiWHOLSPd9bY1Xev3Gmb8Yuvu3uA7XkuObmRSK
08sthLfSz49yHpJumFXVLhtCk0VSamw0f7drWs4Hlk+WQ5zURlVx+O77RC7RqEWtQwBCzWvuulyU
ll/rLHs0r9WVJb4pPCGKYel/Egfik9UXwA4KPxiWJEb8RmtwGJ59A96YwRdV8GiRfaZo16SaqEPl
uHK7/wfh3H1XaMoguEYFN2A1gW5WJIVArFxIuPln2T3loqRA6EKf7hGi8dlHVg6crBc01HjJV7Qa
ULR8tOST3glCo4Nmspk8XohHUe+5pgaevIKorqyfXt8Xgm1AcNmPFMUIKxQaipp8pR//I5KUfkUZ
xQ2wjEnSoxXKk7jIYq0uUxTr+nijM5EzVKbVKm9SdpjEKusARqw6/WgUvnpsVNzGsJffZISGVVpx
vHptGbaA0X//7EHw0bhFCF9YMxxQXo+2wdHyP/BVehtgP/hFY74uJpvW/2rObDFqdQjlqy7hH/Xh
hRCuo0e1fI0oM91hvAwNcspiLYd2jjE1nfF+R87ZXwya5v9W59k0m4XLLSas+BTOFeniIQ/EmrbR
265aPltOkn1TcAzAz17xcffAl50LBq59s39BwuqKZaQYTYX4FVYHxOjVMwuWfd+fYLMSV7v43wHj
kBrUjrkZFK/Y+/4bZh2vTc2S2khNheC30IIhr9+pJ3ZFnudIQ7rJYwpmLjSlmaQcGVUaVt3D0NnP
lkd8LsVqw2dP4/zhRurDTrOn0Ev0+Ei/2SlyQnp95aPD7wIS4OhGfVfm5K7YOfG0SDZaOgfMuI7h
n+phjM/ahPfHPw+bsmVVyGwTIwza/HM/zbyrU/lzSFPiRwLwBbvlwuOLf+VkIxqub61RMs5iT0Cu
hCWwrV14gS73RQmnRxK/YC6gThU+Ww7/cdH/KTLW7i3p3KD7P+JiFKNd1D5IAtWOn5MJXixiuh0I
OnO5lQ5ApXhP/m+rp6AsetNuaGNUeGrdm2HOkxjlhklI+D2EKy9F54MmA3KvN5LkQtuJRObhG7Pw
C9TTJYBo8pNMd6wHCtjcK7t+C7wPTv+SVZgICnYfHyNvTUbtbJBjx6MTpIvlQQslq1fb4y3pcOhs
0yXpD7mWkqAZa07vargQSzzgJ4sL6amNf4Dea5tjHb/etb5olkOJBFfvPGrqyFKYGZ/l6kpzdx3R
5H6RVIFp/cyhk7thmqNnf1gH5cjpgYsY7IbPyAqXzx5CUqNEkIgXnWQryj/0rWdkkpm2ys5SXqsI
5S4jIwJo56n2Qg129qKab5O346s/WNchDEwVFItQwjSo4jgd0e70X/vBXjfGWceeu6ttIgl5ysHm
tvJegQ5aG1yOyBGxGUm8HPZLHcv0H4U/zGBQJlL8D9pI1uGigXxt4ypIEggEHKtxLv2UTkw/wRt0
0HOlH2KZ3IWOwebMfGmM6v5lP5vdkRYtAX6WIH1gDyakdN6HFEgOwfbPOcysqjSlEwKsqiGjuPAA
G/GP5ReP/uqnJ9+bmcwqlYdBiFWj554ryPd9EJhjjY0p3QC1NbWsUscMhbxSvJfuxkeTfMWdgbu+
oC+5ZkhHMdir3dEk9Z1IAKq5NZx4Ffd+EyuJzjgI5FAxZuYaWsD/Z/DxRtFGXKV3EPhfyZFp1hmU
yrXUd05pAhfV3freS7wvlJJTzGC/EZWKDhkLOteEQIW4MtFDHmPWprDImfVVf66hmXxwfUZjkfha
t5IMLLpJCb0S3/FITHPJdso3zzn0lGqEQ3DccKY06wciYqGuncPneVF9wDTa1Bto97fbU3spA5Iu
+4wy5r0vY8NNG0plz2XH9FQxngoU2I9oBnAeIdWGHH0HCRKXOBILbkXZO2T+dJxD+u7lh+IObcBf
WYYaCt9Xw3PW9FnwA6vZIVdyVOW3OmQGCYy39DXTt/0Ur7sX1twZoYxum2KlBjK8VLJTqhL5Luch
qw/TKxtm7dE2+VJ/cvwiyAFSgdv3609lZrlXaP9EQHbNkSP2wRE9bcoLVHtnD06yN40WsJ/lNm4c
NZZ7fxOPnZqy2QEJMpU+blo91CWrvTC+4PSCCslQ7klgCxAxPAIMkdOqXgKWQGbEfSjVoKeuqDt6
Y60MSZci/XYB81R8wSi1N6DbLKtVg/nsy52SbgVSxxrOOBQVIcPO4ZrYu3YUo548UfS9oS9AvoiY
2pqYlwjX+EzeACiMz+4VmTRg3mYaSVljwl4MkGTDAUchix6iYA4FtR5eWTfV7SaVLZRWLsjU7trV
zgueKwbmVKTf0o+GfBg2f7UHL13hj3pq4SaJeyPVmmlNaS5ZfNq5jzEfvfFDPIBd0or/J62yWE1a
Odl9F+pRzbt0elXcY0ouT3j5/Q4nyj2b8OvYP8kOMw5AVTLTMN6DfAVZ1RSizDLzzrSwBkcvVKOI
i57DQDeX7mqv7jzerlRAKg4fPrSGeUs6yo3n7M1J/50W7/rp+f64K/oOCxuwjR67j4vkubexPK2y
myznmEOvtc7flLvkVDBeLnb9xicb5hYAGpDNWLDw+A9NjmoBdBKJ9kOuwPrU6GKv9ryW8jmsuDeb
NBqOdWV6J+x7rTYnY40tbb88MI2EW57Dn8QVdaRoQM4xmUukkX247+cGaGOegEf9UaYTO9wn5jTb
hb0oL1oWB/A+Hu8dzTFX8ft7nvoaVrl/P6hXCWJnEsSNiEK+VS7LKELAltzMHALUDxcPw49nvitZ
erPlBkFhIS8jcoOfQTW1mel4Iv6U1G8y72I4kjqzipO7HpVHLiYyysf2+Xdqr127hftReKb0P6UY
iDnkT9sibkeVpjwd+y9l/Vb3VGplOPSFn5k5XtsJIk2AVct37juO6gBaj/TgyLkBy9S+Z/ASIbXD
UfK5btrbqNhcQH1AsTdoQggeIT8vm7feYxRWiI5QChiw97EXV9La+3YCDm5ZUl/LaiYWIprxzGd3
ob/3UBb+CBhIp+tAv6lYvKgNwQkoj6LV535KmW6UZnNMd6WWSstY1FEUQ/A/P661y19fK7CVdvtJ
TqVMcG/7ynwJB4WQ4w3xMEej3elO6A1T9SOb0IGCDAik6rB1J6ObFVDKewfSxRJREWNSz6WNB3mK
18XMQlUSyUsbNnP+aA6rQFaxELH2BoDdbP9syTL9EQy6fy8nb7k97vmgF/CY5iscLKLkZco/HmQ+
qhy1IUlBdPmi1GBjjWHXewZy/cC5kZQlq3Fchik0UOnCUHBjdxj6VZSlQZGIrvuacK5Ru4MsezEd
DH3F66Zn4M8S1kHiClOYgLmovNfOLx5XPhhtzWFBs9Sy9H+G+1N9FCPW9Zuo1YfktFXn3vNl7XG1
kf6Yc2JQZI9SiH51vHjtajmZpgSlP2Wb0Ph5J8fNjIGayKEQO1FnGmUiFG8lsNhLjwDreVsEFcYk
sb5g0kKbDjKl0mE3nFfg0Knx1laDRkYxG6INEG4IRGn77MNVYcbF0m24P2bmdsFHcp9AGPH5axJs
F/jP7YQq1HxS47njWoWnX5KSqyC/CcvX5U/T5ovE4KXkgOqTnVb7YJR+3xD941FeQSt6+4E9ynXl
LFutvt5BY6Iu+f3XFnT4W3n/r63/TYfJwxs0uHPuUpat0CkPrxJjG+g0AWa+tu9mnl7GgItSTTbW
1WuTnvlKyh6fhKRyap2lMBv59w0MHcSx38WvukYdW6XMb55sfS55RkS0ViM9wtHmOaBF017+vgGH
+AeRurCYBi19SzjsIr3akXBOzOPrEoATbzzKJVSFxpGZHK4Qy4ZLq+xMKvPRnovlvVfsXJyKxxI1
fhsqyhiK/xco7W8Uy2mgdnJIjpA8hVbeTCcF4UYl0SeFYwPNYNTGZDdnCrVOJH9BWGw0zhBV4ooY
QRws+YP8SfsSRhvBk7n44UeCsvRX/3gQglW++rHEolmW/PAsCgUTXDGr1y5liVDNoKv2uOUb5AZc
PsqILwEDj8gQ7sSRGJkvz7mQ3x8eBMxb+FJqWKWOn9nqt7mn3h+QywxVTRZzm5YJKKVxo53XnSAW
xP/kn0xwls+fN0bPtyY0Oz3Aztwsh40cU2huSG3tjD4YMx5+xRM4gS58SrYNhHfv8dwWZKjsXXF8
GCqHIe/VxRm/mKuywHzKktkVkwualbnqkghxC/BcvHblbPQit29lcxpn9od+i9LfJc8LaYFZQSVI
1iZAEifbT3wSHcrTm6s3ny0PggzQXzd/q9dNshTEk3fOesORULq1/77u9DPFX4Sn4cSn7my2WoBW
jSs8sgAvQ13WlCAyJTKr+/Bbmn3duiTQP59VWBmXt1tjP12/5S2XgPeThK7CcKC34y1RYyu8QCTK
FUCQfXwCNSU6Kmaco4A/exP2M7r+8amvuGoG6G5iO6wWv4m4yu4FJj4g/bATz/qMTNNl/BXAwjak
hRm8ml4fr1E0qorTtMRx2bsro27crBDC6gGlNNYH3B35jYObmlzA8abhLqyVlRLV27LcWUOl0Jce
oZMoqA7dW4lZRYd3Usal8PF0jdWJADStHYBdskVx6u4mZz4E3EYOfQlbmt7u12G4xpkfrxkj1Jl5
l1x91XVH6SvHfwSaWUBjvJN453NrTiizYYYQoTIUnuo2bCUKl6NOvwb0mF7eBobpbJhGF9WuL8vV
mECLVKnRSJwc3kT961LjftEJZ6UjFzhQmqDJStfxNln4E4u/tIM1ye37LUijkXJNEw3aWldDtfIV
j+O9LWIBiuxUZdi1bwGuvMC/SU3xcoT0+xGwQvx1IJ/1s1ord3WBxi1tX+rAzSa9fwBLQTjuuN0K
porj85AYLhSnwkEFhEllsboIPV5Ac7jTE3PpEbq16AVtMXPbY8ktaKvswiCV2yz+m2c9/oq/OTSn
FJwiHDeDBykU6KIpZAJV2V0tIvC5eXjtqeSbN80a471waAuKetrl9e3O0A+F3O4Mao3vkYD8BW6C
Q657I3D434hSKlaOlTJPq4+t5mV+qgpBXeBhylSeGpxuzHUVLAf52sq54m3TmHbSepuSJKUgdwh2
kv5W54sKI4Z9tIzIOrPs9LdYytSJJ4K/10saxjsgR9ATViB+afjQpOWEOl1LHz1vi2SgmSlJsdlT
YZS7zpOG1jrB83dPEcVgmMqat2bWev9B8rh0iC4OjTkMkZM5U0Z2wZtYlW5TP16bpebKp124NuxC
bf9tRpsk18UsJDqxR8WmY7zUpi0mOfEE80zmV4hDFOzQzsZsDF/Vz/2RDANGP7HTKSc2mGvb8X6U
rAaOui0mqZ2UvbeYtiiiiGX2LzN+xB1SlUIhj/L29nLQUoGF7JSer0esH9OBelBfoY42GCajJoEK
hLJjQkAvD0qCZ++Qw9aXFOBiFPF4Skc37k6G0MGl92Ch54Vo52eipCuPs0JUrAv5KcjrOPcOxsNk
mnUEk3jP1BZbU3VKO4WJEFZOjzUyJXv7BO7qtNaTGoTCkLrIB5FwCXWYELJz3U83HB8DeTpOYwYR
UxrAPq9d4WG90mFjhkDr++8KO8F3jpR1oAouIF4keUIanwE5cQwp++kWh1X0rpu1uvHELdq4ThKl
r+yEIirKyWLIB4fuHXP8Jd3NXDoovVmnyI8R5guaUGi4TW4q5usMI6ci7vUP3JXel8P8mo5DbKBx
BNFZsErGVFuDv3EyOBX5sTXvIa2anLvwMfmnPzQ+OEnoKllckG68ELTh3awahQmDdnBUHDZtmfjT
H8DGu/sv1HD0X9YGGXoL5j7KtGVxviJS7opXWCHedWJRddK8uCfHviRy60JrsJPVd+KDmW8S4aWu
6Yct+BstOmRgVT+UBrIg3QGrPdX+mhNgWKkcL/L8GazXTEjrKygSA64E32R62AeyC9ThPBfr2NwH
5OgRZuVce647YoTYWBjTXan3uh//uA8mcRtyYDZ6dkZh11mMSveTtXRatwKCoE969HwYZiQCFbpp
7MFmDv1KeAhOL4I9DK8iIdy28bGnDJrFPaUibqoXFcuMHDxsvUkIuDJ+rraBtDmlrQiYUAd5kTQ1
UNjxtVjihPJMAigE/OG8Alj52lt4mGFuUi3YRubAwcTns9z+lpfwSQ8LZpoi2VqDmKThh+Xyo4Kh
EORF1h89hkgmFzEqkM4TjV0KoCK5T+lFoIco4t779HFGQL5fXEFT5tJRjann/ZhOgAyzZ22Jn0Oi
5MxlXN1iZ1n4+hPZwPHnIH9GzqfwEfOehiTHLX5qHf5z+1gg6+Re95XZpbIwsAS+1qT/T/DGID5y
SfP/OpIptEGnZhwqYDpYGwUeGeuL0IVYkwbpotIT2U7QgEq1yroBTIoykxlFhjxydn4Hdr232l2z
ExU+VolxpC9r4UxbN7HaWlcowphTVPzhTRmx2CivvEsUgwQoru3W+s7CeZ1DXbgYvU7H+1+n06eG
v07P0knQXy9YEhTLnsg1aZEiz/w7MbqJz7GcPRf6sQW0bFVniJKn8JcJvS0Zc01GPONPkn+26UpF
y5pGJe1xU4cTltygSprJjFqWA76Q7b3radtyZ0b8bh4dZMXoVnpEFOrF6oll3pRw3a3joOwcdqrA
YhvUREl4G+A8r07/Ijs8MTzj0I0+zMX6DMO0Kh+poWisIiBNutOkXHm9nLHMk0hCn1mYPJKM3Dqk
7AlBfcH+VHnKUsVX31Hs9s1RxAyCIQuQK9wN0Nx+o4ndOAlC6L+Zfy7KvUuvSyPtub91phcwGcVE
8V8S7iGJVgvCCHgoWzZNavmZI5TnoNt58cXbNIvOCZVMfc8Y6cZObSf+Ykbc2QcEbje1pmlN+bnd
minjvGASwMI8Ocf04X7GkZd6DlTtthUcSJSuEQlM2XBOJtC4sHOI4tKO1+C1+zJDpYulTkKQ2hov
jF8Sei6x3ScRm7fPmovx0fv4NkqqSbsifkzalnge2dlY+IcSCnPNT6yB+8kTpZdrS6TWNQKBH5AT
sbduAT46sMPQ2JPkE/WlvVwnc1u1F8CCaz7QF8O0R6no3k4IyzgHeJW0Oq9w+4zyV9zPJrv8Z4G2
SRdThH7zBeK0rPeiF1bzh/EuQllVC6RSGgLvJr0DDfhY4nn59sMQEnG5apg8iSjdi4b13jw5+s2j
Ou9mLWWbV08qACEkYCGEexJtqEa0V8RmUqUPHg0vAhERczfLw353mlp9nuXoFSANvmbN447yxGDI
gJjiylj1pIZGVNNXxkZtHJGggy24DmLd4WfHA4zh5xbVk6vZNrXaDaOhTYwkNXagrAjjXNUXhKNd
sm1te9YBMto1g9S32FZKYdaow4sTb+yluts/qzjLAYc9RmscZ5myBIe9x4wpjXCrk6HM3uvwrez9
lqvq5Jrl4jkEKU7gYYSTcCQzioMRzVH1EtrkTxDgj0YcotAZZUTtKuPMXvvjMr9pvfxP9jbRkpdI
syc7PqKGtaaql3qpPVOOYt/K3iuRUKm22+3J0ElI3jdZ8yXxOkPtk+6ep46hOg9rtl1LNPuxbIF4
Ww8+vj7jcVLrq3r+uld4JWiEQEg47adntbypQQQbqvFljJVm2HfT4Tv2i5R79b91nY+Mdk1cla/B
HF5Byk0GvhMsHVbIKXm1gB/VXfcusqjvMndbXsyAGt4NldsYDn9qY6MikA6eiiYD573QQjMzgY8O
r2DPvu8qoPmtT1VUgePmXpTRAH/l6P+ll47L+FN41Wt5it9SNS3ilwe+DrTl3biEhxBAz43Za/vG
5lB88+35em15yTvVJIhHUjR241ZGKjT/DmxhpANAOPTEVpT6D3j2FStKFuyHmtW8/gN6HKjN3Qoj
Hedhw9DPIP57pfGG23zPuknArz84lKKmxQ/dLfzghDaim0kPJ+wKH5Br7OWdflOIcLeltDco4zgQ
2dZzh4wJ5/ii1MoIw7kut5mQv6CyQFekgh805gSbNwTZPe5yevlAPue0sacCTF6qXEZ405T5Pafz
/vdiH2jbZxTs74lhz7oV8F9M8VxAWdNgn2k7nAyBAWS2YVkEBBAV1obZXhutpdDPyTSA4lYsynoE
Q+fbY+c5wd9PaiHEi3Ey9gEiK+yihmbZW8PhXMX4vgKW3+OQdABxbTK5u5aNuqvByzo8XLJSFxD4
RZbzPlsVv9RoKLA/xBJnlnxWPfGkqIDKPWdQqlCu7cOyGVJYZ5tRLhdIC02jxztZ3wjjOUlqcjYq
L15uf22GDQ/JEghdwJSu7xOCqGQLpfOCiMXs2sm4LBlvsHLsPraH8kknZrPYM3veNmVcG6/NvhSW
EbSkHyEbH7T0VFYUyiJfPGwgtmGOhbpME/Y9+VSUhNkNAKU1PpwSXznEvKjNFwR9gGUKheunGr1s
zDvj9WVmwBpTY19mHTVV/5hwHmGrbD3mgrlcLIeJp4PodFvLtCJYc+dkMXfa24xemabD2oWK5U5t
ulOuC/2KyWaUt5C9rlQ/DE2UQKqeP2HNVaQZdsp5aAzXag5MpoQwT9K7lnDBJn6lN4CVXlLzjiri
0DnLKwSZIwmER1ZvmwtrrXSSlpx/IrmrVAtY6sL5LMFavWkH1IBUJ/6Ea6sTBOpB/DQ/FWp/4G18
N5sYW6/axRybL4JONBJzfosW7+SfCEkB5f9C5y+oSPbBauOcfAeKwuUcJYGNi096fd6PTxJHLCAe
CwMjkv0TI+YttRGaYM4GO7Z5RoPG9MkXSqUOGodQpPcEXZvaO7HAQNiFIvYRADLHUy1DiLwuNV65
ExQhnaUVGQBxfBH7DDqLcJd3G+EyqCXvk/mTE1Y+f9vj4DalMbE3FpHdlHHaOxGwGJ468FoVHnEx
D3Fyil4Nsi23Vbm0RHU+sPtpgP7A2l2iXMCtcA7g9kndOOYhfmCbCDovekR/6R+dL1XO+pWr5/XM
qqUgO9pwFM1skGQB1BmA2ULFrSt9kO3xaER4Gv4vxJBhSZe8KUONkDys860Xs5P0nDcQYUGOpQht
8Cv92gIcE9aSbSEI7dAqUrO9mQ4hJ+KhTs28it6sTC2rHcizERoOt8jtPXqJ9zhmCc4JrUf/rfNR
Ni9oy9dpLtfj8NGl3PJIz2NJzP7gk2AooUEAHvs9gOSV2YbUW7FM9eFh2QL3w+uY2+ZPATJkxTx1
e81I5kCu+1FlEMjgyGcaPOAS42qRVmTftX/ZhlwlWvkoMHlpLNX0Cgf4hezqZXk6+TXk/9E08c3D
M6XOoEQuabE2bkbLzyQQS6/sYkh5YCzlgIxYxdpylcqKTXQB46zah6Meuqm30qWOeWbcFG06LOzU
V9iL8ePz3vfCYIeID00o7VMroQVeiGFRBBkNWolAoIjB0Bk3Pm72vdLTN7IeE5hiIuMdO5UmgyeK
VsoLyimV/1O9Q5ShWeHLa/oe1PBXWNClznAKn+o8js6AX8LwvEEZXCB/3SeV0WtuHE3TtOV0tf1J
9ghnkolvOdoDvBScN8mfF4/C8jwprmdXunRXVLyN8EJy5ZVgpzkeBn4HLijGuQ4V4RIp6HACoo/a
4f/ZoOKdoyfqTJPA4CSSnWS5k1WNDiyAGe2P/LrgUCyJ6EetDZxBmrEXbhp2g9DA6+zgsKe+myGj
vaAEQ53rWOjURKx0spHN4Szi9vKdMfl99IvsZ/lJnGG2D5MmUb6e87F3nZioNW7VChtoNPyyeGwK
vS6F0Wm0HLzGZu/flMW+HjDJuqeOqJ1p0l5KNTjsqtJlEduvSm9OOQXsh3/cJGMCBDAzoXaYUacV
s+5i4WRAnNbT0NCAnqXD1MCl4jwz69f1ZhQOVNaeRRvrKZzwiweIM0bEa1SMJH5kn/FYDNp0ZLYR
pR2iv2lNbZ9n0eqTsek1s3wq3mP0/n10TF+TJ6XscaghB7452s8pToyd8L6qR7LDWgIPKLW7yXhy
czXABJO5hlLPcWkvyWyDgGfGWApXlaYh3+Z7zIo2tllxgAtPR+AkJQuLuRhwEDYyn7E6BYA5Uxk2
eZsdS74gd5vkwVsLOAh9UN9pzlbJT3jUNhJF99tmcPJphIIB2vzbaKTxayxnxs3DYEVFYnqNMUem
LnQF6FJ5aNyeoOIEpkz1dGVgkokH8ZA38tB0hy4GzWJGCRAZOqrPeT9/Bvoeoonn55jI4K7Th1dA
8KISGsWLoMKTqMUZ9JVebr7QmepCIFfjEMvm4tGBTgoBOTrJK+00kwco3jW5Qc6+v6gB5QUXc8jQ
LIZxxUxFLGRRuEWxvUxIBoNmzacgeYVwzOweSHINdD/disS6vSoBoOgd3VWCjFSzlsSJY+sCBWFT
fd/Bd65nTj0e2ebS3tvBwrJG+rMS5p/ywx4UWnB62hKMcPCBDi8+bQMPDvKnn2fgeANycrxYQHwq
EI2Gl277yz4JaB2f4J5aQsXSlg1EhFZJAuOPeE3Kv5wG4IAS2yaQfLDNdbfIFmiN5rPIsIPaUgcf
xLs5CbMJbIE+9YjIcGBW720itLTE2iHfFU9rScAPys/128NNTEc1eKsXDIYUKJodV42tpfXU/aVW
lFAqxcJgnufA9A0Sim/siC+oCQGgqoUThdY1LYLgSSr4kiVjw5I/4OujX6qg1TRWrxRDdWzDVbQ5
OyIzqqWdoWA9U69hbH+o0Sge4JKph6maK5mZbwT2/EgKWzAz3Vs806UzZ8YzX0gU8zMDVjZbuCYW
whu26svEQObQaoSYZ0QscQl4//4DW7HxW3wGNROSeistwL31/DzYsJMqLUYTVSC5CUDJRnbUXDKT
Pksj9ygZ2cYidNg5JryZOQP+rmSkyzY/wSeyFwFj3JmHC8NtERK7/eSVHdLoS8buFMspuWx6w+gH
f+rexLcXFg79ChpJY0dWpz9Qnf5cbGXrvnm7TeHR63ZruPmQDafYb4JRyRx1GKF8jFC8Eht3qPbn
bCCMRW0tMQ//6+dZpImyL5FAxEjqtyeMNYyur1ng9i2PGF9b38gRwDypkx5xQXZD0k95CVCgjeAy
aMRN4WWLxh6hQghAg/nurYJsM2rDQ6kBl8IAmrqdPV/PFIYuDLEGbv6MjRS4DQN7H3cfCyvKsq+k
2bdC8QJpOUbJJU9j6P8R1530nIFnfJShIbOYu4afQmWB85DQq0RWZQxu83Q+/yXYFxvsWQy614F6
ZEawOkVBBzNfxM1FIYztSZMzVivdw5jZOVIMINw3P+z7ohJYiNKpFYlL/wSBFumgyBt9+0+Zvq9T
rPyFPex314pk7Gm4+YhBJzTQ2MCjy7J/qRhIyB5FLxaEcq75LqNPTtAQpARI8nXzvXX1tKphlQpD
NYs9E3jwmbc3JZO+E9e32eJnIlia7dBAwJFLWSlmcCCfQXt4W74gCBzP0mR4jD895haH3Z6p94UM
ZoawprvM0zRKr4QGstWsEoOVzHPvYuC7Z7Y4puxb4bRsDMyyhWSGqXRlZkdlBCNsYCz4+fmabj0L
7gmONWUbK0APb6GbO0dNvTiXnosfdULNBD+vVjTg8PXa9V59O0N7iJMig6MDFS5KKTP0qFN84K4D
suwQ29i8Qq5TQuqWP743tVmIlUzuLhgTXGuH4kzbcNbCGXeOVE+dbA8pY/7cixzM2Ekd2cGtzQuG
9va/tfRyRGNwQyc+LpJEZDQVm2Abv5qiMAA5iFKXjURdihyhjeqlG2DZPMbzsWMpyV9+fqLbDf3Q
Qv1H5ulj+s8Pg+a321nzFCq7uUZF7ByY5NvEdlWBGBTZsDaTHifRXtyIGpPfEtKgZWzdaVibhzkX
PcVAaDLYZaStezAT7Xg3WGTMptmThpsFeG+BY07/+tDcVTW/g27huuSRC/EvXJDDoYaWeEB6uNnd
6VRNvLO7RPOWAKPIBgUFwZMyLq4kqm97KvtpKJSa0/JQDLowwiBjVPq7GYiL1nI7l/eInXze9OzM
fYG5Vl5AE4xoQOkiifXg5aTHbMvGym7n7oBk0tGcAfIsn/mAoUOGGvaF5MrDx6C96TEhM497wR9L
E4V2wLAmF+/JXDkl0/ctKX8TlEfhfYAwYcLOFFtfBSnpotfkgsnLQS0jSHmkD1WlFBBQq5EAZ8md
5zSpmvsgeabcBFaTYQdoqalYyBnOpughGa99yn9F426rcrl/FArORSQYTPybn6it/GH40cyKJduu
GGjOkvRwZTcJ7uEF4jr1W8t+x4rYgAjmjjWWo9UcunzK5HahFzFdqGUVA6J+Wu8JgiVQsPZVC/e2
t+xD5y12L2D5pTOl4AaSTJdANI5ra1oPcVlJ3xPm5KDDNoUoPjte7ee9GqBzO8LpZVMpkZD7z/2h
FDXVzddxT9jHMY8m4vEBS7gPW+Ve2q2mqxMo8FikpZTKDVvs7iLXKftXjNIKjgO6u5JfwUTiif7x
xuLCrMIEkFqq09Ay6C3n42NglZQv5bGU9LVn29+kiz3vQyi4cEHltxkyyJwog1preVu4eRfeImxr
aUa0eq6FwxhD1KrqY3Ba901votv2z+EI9qdgIvPIpnojDs4e9+LK+aKQ8kDmMVtu3EUXdor4XCN9
3Wx+DXsrhtIn1SFps9XMzDO6rbfXDkjuaK3ZGcVn2agEC2XU8dkpttDk9A7emHvb8NQrZr2xu5Xa
I6nZz4GS1HveXgGD2X3ZrXowrkBeXLL++DREXAVYS8JoCVqG1F3hViTXmy4bNSHYkWjxbV2ENNqu
AdIFNDhyNnORrt0ev6DpucI4m07A/WmgtuXiqOIi6z9+5MjY8VhxzxMa7bUVjoDgkE92haGLpYtz
BeX68UwmGZzR8cGtyfO2hEmGqRyp6Hbn25MuLqQsskGrj+ON4kvyYuDVaYSaT/TugYoZ+rphdDcu
nJeiSPriE9U681scEyi411UPibuGvE57zAYvNMQon/ISxsKxjxl+yhjvBXbHIRQLo3C2JU5jRA/X
kGnq5ZiXqX9W1lFkxI7OZjCpyOW+3btUjdiW2y4unyTHTxcvZGi/67mtwuiDz5s3g+yEGV1tz2yq
lbmE22AEwTOjttEmb/dbitfnQvuZcKpgLZgwyuA0Z5k3Gfr306Yg/rbF0YGC/YyuEoOZXdZFyT44
iCxcNYKLEP3SbsSFbzad8o3yVLd/BxVAS3xmS05ZScat7AMxjPrg6J6TMEREMCArbX3qo6u9yrw9
IDWfujVoP8AKR3K5WbPY303sPG5yG3ZwiyK7AZd6devNpDZDWJOn33qMIBEtUsMJp6Np+GxZp9qR
eMSgbExZyw6D9nlL0S4SISRkJDaYbv2iX6y6Ft0Og7b7wCSZL8iaHhWV+9B0rgItU9Aq6orWP9XF
hK1Fgjw1bvv4VrE3n8Jguzv216fAkat58PDOdf2Mq+vzcuFjmEtCrvBlUekTJTsPnJzQbLAds63C
eqSCtYZG2uhmA6YhbKeL1KhLVfseskW+EGtMSGzSxkexMDAUv1wgJxGg1cItNaVYC6pmSV3y620k
uzL9JcV0ScGOx+aiOfZis3DPe41NIxBr+2QFiT09+zEbRgv1qCTDmV4hUJlGO7VmbpVCMU9CJ5c6
axZdeTukMc0GLHLovY4lLer5A09Dj+HjfUDy3hHcEQflAfrYAhJYRIJI0LoN3xRq6fqIpywONaZK
PLaK66hwaKLdWdwh7owPbQtMJGX1Pt0phurUsP/29dpormvfijY4GaE6niyltzp0gVbWDD1YnTQm
LJxDsbD7Aem8+HaxNM9XeBGgUCncX1lI8DGURYUxV+yc8wAY+iLnX60UhHp2H+YoQx8UyKN+aZVd
4m3eIm5zUJUVatot+D1LtAjVJIRibSVOQ/lULoNcFtM5b054BnbOlM/Dxahq1K0d2upI6xBXcCZB
gIXCblFg/a7ZJX7iLP5p1Tp1ZMVhBr1GTmdw3Q5wrtLgHVguI2/QTwKmKCDgkfOH1prNJeiXrJML
s6Iux5zAa/ZAekH4qWR6F64OJqNtbfH7qQpWjwiQ2pwtKNm0Enyx8OF5OKdNTfmzILKh83RuQkFl
InNwNh8maivujBwL5wvfP58kUxn1TSAgzzNVnc7NSViYAh8t/7W/Sgn9tWjV7Nz+YaMm2fr+y5eQ
R6QsRGZ/SCFBvwxb1Io8fG966WywpRGhmPbxv35pyUFbxy1w9Am+UIXFd6W1Jb8iJllU+u3O47d0
+fPImCAzF/zdXEfr4HwoKAydNe1bcXvDRXcbaYovoFNoEj6Tsf52XV9QgIq43XLPpjvGImQ3cYJI
pz2JZpOghL/psRI84YOoy/405ebIqV0IzcyMicubZiXMn1m8dC+FV8701sfO3Bomsc10/ZRn1ayL
cTbNpSV2+1eBExJM9Q37bss5rFtqgHu0JHJpQAvnA1qdGUPfocTmZw1f1uEOjXBV535anJQRvBDy
McU3KWN6iilqYEkMxhkxZRPd9xzs69EHZm430taZogqigAJYE5kXCCDsHS6tsBMRgmQeln3X4zB8
qLxd+FJe6LS0HqF24gRjc1ZjWv8Zd+0NKb72BjQ74/0VxkrfWl8oQcb0RiylFxIwAqEBqg8SgjAR
AlI3FKliwK2PcKg/sCPWmDfoMxsS8bwncTqp5T9USqd9p4eHcNy6NDR47bEOEsA2Tp26bSAz2EDg
RFPvIKyP5k2TXrVkPw94YZ9RcnfnGYei1OZpx31bZYBcN6bI5Oj03Dd/OjrHpRjle2WY9RbIbtsG
79WauCTWX54gWviO8/4l0vK1qiCSqxswopg9gDrt1LkCZ3kMLWyL3Ozy3S1e1sAQXneggnN8HCzb
aXa+ewnkxU9reK6K7ArtVv9i98pXDkkh3R+0jUooAtiaDlIlDW4ejluZGUPeexAwmQgYEJLAheo0
u24dYe5iyegzwtzrUrZow3eEimJRl7DCHR5z2iavoCe96zXr5Mb9SPui9sVQ5RXPbvaUwbGO/CXk
EUYyjTpLPyJFw7PB4+e1GGDe1lgEJYGWYhUupSQiScRsmdgca2mx97A1gas5CYcLCmYVkn0jUb2v
5EcRTjTXXp5l4rV7tYwnXgk5L3bvdfC78Pe02NB+MkpsIqLdiDaevhd18mBBqeKTTo9oY19FFJbc
zsxzhOtoOhAgeCo7p55yiYWwMUghDqBHy+AEnmYh/nCkEgOEIF83Gz3BYsLt9/sW2rW1fymct8g5
RvDgMvWR4uxMitySBxEtLNCa63/1R2l5PWX9+Qg2OjgzS+Hu0CuC4zeRrs1LPkY3kcxPdUE3cE3D
3e6+pAHsjWUlMl1EnyzO0oco6JucIKzVvERhOQlD2885H2tVOr6j8Ye5IWstXMTowCdgwtUptShM
1Du0rGzQ1pzOYzPIHDdv1bYgN99Vn1zfnlPGf4MhMoiqjQbmatgrxZw98AptSmpXXJwZNeo7l7ge
GxEfnWhFU1Fx6ZhDNjgG8zeu0Vy2VEE3a8FWx0P4dNMDvHRSJqf+/c1BWN/wghP4O+Jn14xYUdsW
rVeUrstNKeLJ9utGsdNsZR/wVgnF5znXemICXQNn/3N8+RgTYxKCXE2qJvOVgtBn53ZrS4D7PRIW
SqusM4Guj3qLQ5AxPPRinSOrsx/PCVbtRrfSV7DwC7L43AIl2aBvXf4DHF9wdRGRrt7VBiO1Yxz3
hSoNPVHEYjaHQQ70DQG+jWN4/j19I6HVYF/GGb4aGYcbRZ4dQda7Nwu8bdwg3E3SLJ5ltE014dgt
hzt1/gKJgic3Rc/pOZ3qWaNeFQ4HKpaFFqeJICCeALC4u86pwm26Yh0UxbkUl+6Zsc8usFjCtF1/
zJpw/5EbDzIxOyC9020RrKVHNdV1yAEPHJstomNL72hpoQMuO7vKf9Cf7dx7HHjTDdiN+Igwi2Nj
/8rzfl9T4j6hsTasRFpgPriMwL/yhDcamgLYDhliU8X5D/cw/HW9omLd2/XcKLGOnuOVV98fxNGB
OcA04KpXC1NlukqQ/BpvaZmbMM+U0R8x8DfyWLoZHITd/N7kD7zV4lItIYKI8gNit5udDvrHJ4aN
HgdLGfB2YowU65qlvgAgaikQHBQdaiNb/1jwzlu0ESNbPpUyMSZnvMv6HRVK7ntw0skBe4+VdHHi
dljCsAy8QugAV/wFiD+mhXpEYlJI1xH8dAsndtsXGObKjmCyzpib5QO2OkGW3WMhrv3WvwTniWtY
RWpKyFYuEtkWEI1TEBq4SXjZsYRZBaDTvemyJagPP4ilz3A4wLTVkJmaozG1UdVaLilgr5Zn4A1N
/JI3A30z198UREDmgiP2UoqoS6aNlP11fWaIUqsBh7cDzmeUpmVpwxiQWMSC3UFrv4OeKBCH48sj
bFpJI+EwOCvwkXXrRX79vQDP8428JUh0xAf31ybRkYg1C8k6N994J21+3cu/AUSu0lFMne7o+782
Xe+rIX+5vbU5rv4fX0IPiSn+ud+RfkZa+V9k8sGlQiKpHNLvfjDoHh3yImvXwQQpO0/otrisZAL9
Ul+bgUa8lh+dswtL9yg/b/W8kayPs664QEn2deVWn+uFVAh9Lr3wLGhaYwERnAOJ5XRAfgXrLUGk
WlZu3GmFSMMpjYVkVfAoOsowxpcs73FFZXkvWTtI9FLhrcfcmBfrCLh6i5+Bveg1Imcv9heyVuIX
wHrUnMmT8DJhARu5XmbFFxjC/BYp0M9nDGh1jW8iEkcylATRImm3bgdsgpLGq8XhS6l3YTn2i5MH
oF9xLtSElXpvMNc+/LftqsWHS09owcCgJZVB5s0YIyCyq9hfBSTcbq5yiAxBFmEIXcjf5oZE378e
Q612PnEJrgYbc4Pzf8ZKqDRjsb0WzeNVp0Ztjzm2GFpW4BQkuMIy7P2aluiS2AZTIUllnuddGmMN
KsQV9fdcbRdOKbr+SieJfxStbE+OrCIcEXJMrbXqM+1IzLphjWhm76AdwTHio+j1SQscSaXrFJMW
iX8BPmeMVskK3BONZyfJQyDDfgB3iKBrAZYqmxImSBK98WRkmFqq8Ef/0vfRT2yvqFwY5cQXjGoN
4UovxpGQHdZ6hi2MzMfbCBKCoZf6b/zHNCXWhTEKipzDrJBb31SF+HxLbrl6stzbWQOOo5MDy8g8
5ti/CgBt8tUJGtff4ZbYjPpfEur3hWlFkf7Gvi6y2w74mREMPTME3bk5tCdv4IVGHKEeNLdgMCLp
objHYOeOrjvjPgS11rJlbJqaSFQ6mFn56P9gmGq6+hnDY3UIY9oNn7PVQUG7MNdyZeiHHtc9RxiW
BgD8eHf0KEk32Isn46v4HJoYDIdbQLvmP1Tzr/C6/s3ppBFC4Yd8EksLEBXYpcG8kRZxWmmGF3D7
ymSAzO7e/qr0X7xda7wfvQnVlp3UJhgTRmQbQceg1ecnzahv1ajWa9+WITAyz+RRpG4s6oveRsNW
vm60v3mulsDkAsMJ1dN2Z9z7wfUvkuPJeM2cVBtzHsHtF/4MhRZwcOmF9QnGQFlzETc0whpzoMyQ
NiNyxxoW5Sv60o84BmOsgagTkJXrNSgENBEaL1cAOR4ojzq5rrYw5+Sph15rZQodYEcRi1ONgpWE
ZHqBJBT0vx8zv32Oc/aCbEDFQQrUR6EGp/wlCMnq1NiTBa+zG9RDVGtGv31s3m4lhy8ClPZZsc8y
X4LXRjLYy2ZErSKttyewAmNAa/W9MG2I0c5KQ2ZttTWNtoEeB7ddy4auaQal4/lq65vOWf9LQ0fL
AAiOfymskvpaqWbYZ1l0aukXetnZD5UAyR00YYyXDOgnRVLMrmaCIxda+6sK6cR58PReiOOuDprn
JeOSAi9C/bqN4iqb0s04DjsxM27DmCIM9nNOEpaXcd+ZtsO8v0JDD9vYq3ukfDzSWvGsAhDCi3uN
ePVxH/cnu0xGeNePuCdwuEZBbvHPfezFKZ3IQpWtdPo1Y7/hCi4r6+q3yFpOaHoFuCTSkZIcmb7B
WcybNLUz9OLWwngX/BVhbOx2M1Un4PJ3bUkGykwAOSCxz1Lo9C1QQE39PRWKG+07srfMTg9dlD0E
M7f2k1dVCltVtbhDFrgguVseT6C+jueif2mAHomg68ogkFPIyQLhZzylZTDGE4ZRcEU4sWfYSnD5
X9jUnoyWNrQJJtCy4N3Xfcn6lwQNCB4Kq3gEloYpDUX0A9BuQisT/Yt2WBM2mUvPVgGYeBLiDJZW
YMFQvJIcmFW+WwCWSHXpvh9zak6b/iEIE47Z717EYKX0wvp7MyaBm/QFBpc5AErHhMERC76ZMKyS
LkLAv9qKokRfhm70pzWUqoUndGTaDHaKwaQ6t8LlaA7az9rnVirn8SAGuzD87N8eofTIQItQCkM3
Zoh4GRGHkLPOItTKM807GscFaKejp+ebrr0/qWZA/vDSZ4i18fK+LDaj6KZ12hz6ekQmt5UNhFy8
+3wQiErp1L4PGSwodBvTIHegUBAUi+uCX+4p84aON3yRQxnrpezuvsTs96lI/Q/mhKAMOlCLVcgA
bl67kvC/uAyYN5kNA2XM6l1ylbigIa01YAYKdmHPzx5FMEQZkExiJuLwxmdQVqvagSsQ0adas1uZ
7bmsAkEn/lMLCSFGUf3s7wyUULcjXpMMIt7AOqpeJMidcw4uQ1xbQ3Xzuf63SityOwJbmSBQh1gV
1oTVcGoaoI8qyI+3mkUKG3yhFjBCrphcijMfGcMu/nDsfCMumaRXTxZwmwYRi0gb9TblkVKLRuHX
PAc86GjZN1ZrLERdyjLw6xfpN3XHjaZHreW7o7hUL32gu/sVRUDig3X4aq6XRkNQ3EBfdcxxSE72
ExhItIWitZn/AKroSbAYHHvzAz6JlG7AdqRY7+xQ1kBIZZyv2GjL6qj1Irpth+ACXM8gC+yqOIFx
f/BceljUICKjWedPeOJ1Rn6lGma0aUP+c4vDXQIx5aQIbl7dbvIk30N2OvCr6AWyjep6VnO86JCf
TfL4Ktp/NYzeXZIK1MmNLd1reVn/cUJoTytXZV1UOG9nYOWGEczuFxKuAaSvZu3hPyLjEwHNGL4h
33O1dUaWNv1fCBDpF/HsZvPLC11/qF/8K1xiUey5ilhWNaRClQU5M3MbX5wFMrKYwCWnO5NI1QFk
23Hs9JCeEmc8LhhF0c59eQxAK1qEoRnii8lYeE5Sh/vxXbcRgDKhPTemrLhFtGBKZP5NHYyXbHP/
fijY4xm3qL4C9I6RXB1BiX9XZrVx0OqcZsIpuCnIzSW2wc0rg3WyZdetY4Rh0O7PW/TXGCEemiTe
uxXQkDeUNPbPXmoaf2EF5virV65oSW/z8kaiH5zw+95laG7B6mQ0ZzZ8XKsm2CzQFR6Kee1R3F7a
lBIGm9OxAwsq1Jax113ezQzrkASATrvTtW0c6BJu7ucmWSjM6R3YGlw6m5FP4r4tZyd14oLiydkB
drUBHX7ntd/DGm00mmA6nUdc/9vzVHllwEcO2TLQyo4petns4mKKkac91gRB/KMIYeJxr1Tn6N6M
VS/NbcThovaddSvdKn/DpD/dZfjgIM2ozASg+mgaYkLW1L/gyeAZdMa3w2/xo0a+9w/WlU5VNOLz
Kvdjul7xlj26lfB/MVnhdRbSZS5kCEBGBFG/C5Cw9xtGaSLPpUk1njIx7CiWy13DDOVIPcZSYmce
Ev0jiJy745UqsO41HXdpqKDbqzS1UENWGS6KoufEtxuadxS4ZuEX1UN0QxSqz/lVyp8r6r/k2rho
bLZlM/vOvxzmBVYGfa/CRpkiXZj1BUMRcRQNtoKa+COU+YUgdk5cE0aV/9fgUBGAFkfrKTJltt5A
QCvPrf/Ulbzm27uORO0Wx4ivcFl4bSOCdqzqNS78+F6Sg2lsFf0bSfOSCFg4trzRI09dkT7awhcf
3ASKdnxQ1XhnfrdXd74dhcPamtJXeyZ/YniqxVZvWHkO6+nnuv5D2cUCjsG40AB9DP4uVJh65+wQ
LiLjNuuTMtXaXtHaiiXcOCoOR54Fe+tnXy7NCvXGxI6OTvA3Jv2aE9XkkL6BPNL6R3geeBndA6kI
YIgKwO5PemQtaLVqwoBdnPQWvjtGN8vxGj27tTeYDF8t59wAcasr0EQIXuNAlkHMOpPwUXvBsj4P
AT1n52XbOmG5CmUDgquxhMVIi4y0kIRpuX9sW7Df4U2gRYUeQROTd6LXZxhErJjwULiFosu3y5tL
DFkEfhp7POWRVmT/5gpZY8Tgvn5Ux4cT0ng0doZKqtzHO/bfM6KNgSxOlLyB2aT1vouMHoo5a96C
5irK+PLI0I2C0VDpYmK/D/DBs/7IqSSwAblCSBJ/Z0nal/fm9oJSGfRcRZ71VvQzZlZ3U91hbOaa
bJliC7RNBps1dhmzkrtmW/V8tMT4V4kj8HD00CIjaH2JhH6MHBifmlmBVZJsPcuooq82CDVI8pwl
jrRwG9zy2n3CGwJsbyYFnnycAgVseuwgFJHknAgUmizGhfWgtOPEQnY5HkXIw1EDjbNBynt7nrUs
HhTvmBv6oauU6Cvpa/FZsfXHrBknU5TY36Fla4fO5cjqWB31wDQRC3apVzesIxfBfHdt21mIxhAv
wjJqNGNgnaC7Y5ZeTG1g5vfWWjbtcGLPzioeeVBt3tho32D4h5E5bgGxWIFZweOEu25kaF8ap1eA
XX3zxEX991w15SeI9uqlkaBbATjBnlUmgXAzjcjt1R0JHLD2sRZOzAubwt6UHvTsQajMfn0JkeTx
aKlyM1+3VmzaYvoGwLvi1E1PrtM3F01ngK/simNgDK8oQlxyVSU6w8bBn9xeHrTvD3acCdhk3vRJ
JL55q5sCns7bWgxhkJI1B9IFCg482355nV3n+Xxm4D9BCh9ZAa5cXjl3KUMCz6WZZTOE+is9toiU
1DY7CYbo56Yobo9FLOGueIHCnTVcSgxT6DXhJeuIPxYkye38t3A9NXJIjpBd33kMI7Vld/ymXT3Z
W73Hk8vnHFI7NkyTnjeVFLmLZlSExqe1FFqNYQ2CJ8JkW6Dt6R5ekOz1qrrS0m6FgTxi0HqmxQau
G0N9CRn2soDinVP8ZyyS/NL3JZXgFrHGt89QadtmuoLRdJT8tRBI9gamVmaXCxdLLmdU6J5Jygjp
v16Btlp1B4co3uoyCiM9uT1zqx19RGpg3fSCFgC6qNmQKmrSgXy9b2bdkKlvegwqHcXGATBML8n0
BytpMJIyL1R2ORTt449gOVxBiNxzRtrItbpzdcd7zB3TzfnDhA7CoZqNVRPDCxcvz06Wf202sZ2P
z50DZwEewm4LsCFrL+pSzsJldopHTk+l5x6pr82lcgWwoRLrEIBCvA7za7g1raW+OomDlvA+ABNS
GjjsOJ9oAFMXTBt7j+Vt5vr7v9b8Oll86XHzD9oAd7rkOQz9jA0BzMHdtxuX8ewjV1oZtcLVSVIx
1hQ5iM1OurXXyOPEnlhxjE3RYCCZVP2DrcFNCb88GUL9iGVFSH1nm+4efwue3PNzb+p6A6euyw7m
zo37w1eL+AjVESkyTxzcm/mIk3NQpWLE0H3f0pac2JP/pU8AmdQXw4UGLZmvLIWlU4xjzmwhx84w
j6ntVaFmQJ9pR/JmM3g/5FapKc03UQgaR5nBftss0NVTWQ/9gdThl/Dd5mzjWK6zjQxsIXUWEYa8
muIOsqRh/H1gXy5GoBL1Qwl1gyycbduAlpJda9N1xeLbvzzqL4SPoQVYJwb89WhgZ110QmU7iQwa
Cb8DJkXDVqV3FihJj/bdSmZ5ZAN/mOnoPB5LghkQi4eFzSntBp2h4MZK1a8+WA90O/363ThYsWOz
MaX10Q8c1y4axnK8F/L4mPJ6Z+1MwVuRtshPalSV6ILACaNi85bhDn1w1L+fSr1rqR9nkY5mN/TK
TshdR/8LDKwEPa9QsQ9tQhnEc8S57HpHIFNuzpQGbBehzX52dB9xPyQSajPbnrGQn9a/GhJpeMhR
oNt1ee6rPr3BoKgb8HhC6sI7nn6gLP+GtbpO6END4AcZEY40HBCeAKEqZ+/oXr7ACx1jITD4jXsk
oMl8GuZiEhmdivbH4ogWtsxWPIWUen4eufxWqhLjjLrCfaz0oeN9fdd67qzm/7sB5cOZQtMKG5Ft
5+GQnqd8sWySsHZ4smwGMjGD02AHKS2rdpVt2ahKIaG6isgTEI3hi/fikoiU/Sm0kK0y+9y7IFyc
8yfuQMVvFwOzCcNGLLpOYjKo54CJunu0XRPDwpMSQA4R3ZQxcvDpGlR65uuJ5Gw/pbme3yW/HKj+
Kb0XT+AGfxO7UhuM1PRfoinwamxib7tizrqfcrmr9432tHyxLx3hJiyCk+ZEF+cewfcvjs7GpYnY
Z53V42pX/MGYDlVccEhNUbfvot2ebi7E667Uhg/qcTyzLDekyLmCXOk4H8rj1IV0VYiB72ZlKHoT
D7nBop0M95s9l5D9d+dWKPzvz+NSmSNfVYCvYc45tuZ+1tslkm/Y2tU6IkIOMJzpFfjnCHxVq+ZN
zoZsuFzNB5liOrlFj4kbDb/3i5rJ/xIlijKjXE6fpvywBPOsslSWz7bfKIlzD0nE7tjgNxtytYTf
wvBbCgpIPUbXlaPEgpSzANyficl9OUGeZNYYMFOMhZXovUISDeoLalqEJ4dGYZLriAKeS9m5zqSn
mWgnf3Ikm++d3TeHXAya/TsOqP22HoBvMAzFnvq2pU4PimNQDkn5dbLVcVBU/SRxltCUwyVml/f2
Pnz9Ugqcx9O9Q82aY7BjqTES1a2CT82+WULulR4UTjh+rp51ehaOpSmDuHB659SwmTgG8wvJ/EHL
ijPsy0Crtc9UXxAv30gXTOaVzM7Dk/Xq9+uLxia8oiVmk+0ZvEtqjLWfto7CVYqih5zG7sBQvFs4
RTxGVfl2BhwLMpe0TKlTObZuzdyUxDwXXer55FEvxNjB2CmPJTFyncPaH7muSchhKCIysnZ+y+7Q
T+KYx6l0G6P51aeuYGc6QEOcXL2TNz6qF2kz37NQISwI3lqu76E3xuBF27pgjyDeX9Rkeozl+z/l
DODgsYDS65FfZQ408Z5SPV2XlVrxqPc4mYWbSdsidwfk8B6G9lbeVVN5sLyNqzOlQMuMiMeO0bO5
C22VEkH0h16ofvAUSVAESBFrp+72Ar35rYQzHRguK0YD9SO9x0WMZz6PyyCVVNQ07arJB83B813v
HWEXdgX4OHagNpoUJiX9MTE/FUVTucbTwOmhX943ri657i0GwlH3s7vGoLW38ADq/C4ESlBfAMT4
MdwvdnLTAX/raEP+MfYvcsK7Fu5pg25OmkRS5iXT7ftSS6b6DRE9XC0xvTwbuETxKdaJSh7snwjH
T+WO4XlFlpZPyvo1Ic7gnTGyJPCro1jJTYklqratQTg7cCHOFS4C5k0XHG7JT81StnWLylJqAsUa
vDg3GjvJY2YBaq2LDveJudNomrz+CY00tKhHZldkR31ddt3De3LuccpCG1DKaFk37g7vJykUmTPF
a/ZwXgl3wD5PwEaBD7f1yWU6U1sJdvqv3M+Ye7/hwLkEzoPhG3ohVpkeiv5p9TFcgiMuDByNoiXb
I2PkmkmC8z5ozgGryHn6Ci/P3AC5ZXs1CEnzITdEN3yVun4W4CQXb5bfTzIh9t5QApvlVAVfapnE
DwBLWnaNsbOuKkIGTXgK1zswAIicV5g5dIayLyV0uBkcSmu+iUKfGsv76Sv9HbEPbekUrVi/RCQN
i4ECIKpfXQ0B2p50ayIrWu/Q6s2SzHWOsG5uiOByFPAY5wel47tKySKUFfROuZvgQincR9M6MWLT
CGYE87xggfiadWQvaIpc5blt1lmWrm7nU3xPhCPV87teK0Y+0Qfl5tYN/S7dg1Enq82qXGE5NPpy
ymphO/RiUCIVt5fv5kxF4XaVw7HriWQr0JiS7LCWUVZTFKyjxiH67SwRv6uNfksqRAVXA5KnbNFY
z/q1P8thybT8Jqx0+jZA3Zow/ZuCRI4LJB5h6msk/WWlh1Hn5ZsYISpDl5jDcVBO8Hhja+yoZTHf
rZxvjRyqFeu9OPPkzlZOcri40/1dbgZ/nE3iUjRkCUv9UbuRE1jQqscDZyHVCqQToppl1VVz8ABq
g1wDBucOVXyJdkeyz0g1uOBMrLhNRNRVCx1IK4pEr3r3RwM1EnkACYdwOMrzAAK17nN6hzFN3idU
GbIvVvzNlbu2ZVDG7wmTm4nH1/IMWoLuFc4Xxn1hXHa3/KEzKLYLAPGcLyhCZifZFodtuJFy/hVc
8JNhSyPErmj5PBvVyxrZP09/oN5fMe266YNaOHdpKtZWtgJgB4PqrAacXAyJU8k+fBvixEi0CJ6X
5FhMf8jZngWok1kKN7q39aMrI5SrX0EMxRTH6IZ48FRERA0kQefMl2Cwr/hg682Y4wBMYvyn+ac9
GeFUopogHuJCiHOMdfNCW+LlnIsZU3ssgCbLZNxt6YGtHKmx/qg7KP2DuRjzXRboHTYXxlent+n4
ujKzNs2RE/A37lKAYg8gE13CPm46GYFTfcmMQv1ELZtL9mPBJK8IcIr8J8ijIlbZDg3ZNQTWt1cZ
QcTAHj6IADvYTsIRorS/qe1sAhL1uhV2Nl8VTONuMRUBqbY805Btw3KasWGY/DvfQhyS8skTdteT
rCLSX9AlSvw70R8rIDRXGRE3takjL366Cas9dZr/4gmqC/EVbXyz5lUtbAsqbfv5QiFmcktt99Zn
aoPX+MZjc88Bg+qLNFTPrId0sbUPniH7M2++e4nxx5kwt9IjfzOKBmupud3RwPdqW9FX/DUaKgiB
xsoUEfavcUwzneLbJS5AmHAyc5/Yg2J4TkngS13QgkLQw2kg/jYlBH1+RT1CexZ2ehmwC8c6Pnh5
aREgRMwx/ubn+1SlnFlbnxk+yo/cdozNgQjEb7QaqVGOQqsKQKCFvIdC2sf6s32r0MpvUB/oBuZe
iR0ABlaTowGTjFtp6MUNNdINKwoi3sld0ORNvkeOmH0sSbP78oNrSEXlffgTJAvsw6RPOlN1o/oC
IZ+Jm7nUueBmil6cBowQlq6dFc0ss6Al/QoncKOOzXRjGwL9xXs62iwEZ77jQ4Csi78yGdjo+v2Y
NRStNk4L0kPg7BKYvdsimBpQ6ZN1JGqqfJsWQnGSfbaqd3MnK1H2Z3i/+UTwKmktf2YImL0ddUGD
PUhWpVEat+MFhi+gNKAYtRxzBZx4tx6w/BPy/b8r6EOMA6fGJZnrFZbCQWaf8Kr1lK0DIglKsyK5
la8c41FIc1jz9QdZcKnjQDJrELcp+cl6Ee7EDhuYjN2VwHd+AIH8Zxx6IceHi+e+p963LXxDaNe7
pCIuTUdJcOr8HWuq9IfBYBwG8vJnzci+/cmpbpuQJ1nhD7YOp9ySDKHJU7LFSuohliJs+NXPvddh
5ImH6QTcEENFmk91CRmbslnAvoPs6WSqTZmBPKD2ZbY20cRcn0m4mqk2qycjMZ5HP5LsCIRLmGZN
NtWyw1yGKnPBz2KJdcaObOVEGP1In1qY5NKUWSvdZjGaTbEs5UMyTuAB+nS44WXZgOAk3WKTxkzh
m69QA0DAANdqcEoxnh1JnuYZhz2Q6yynpsF33C569aWCeDb2pWpdBzMCotz2ejmgk1iQGRwmr8Ol
weISZCbk4dbBW4JDRVUgG1KGAXIiDWL2wV9hz1djTnAMb3UiVILP3oiMI+/4oIr3h+9odA1/hSfk
1iOuSbNiknCgDUCd4wVk6tASTjsR3H8Mo+Uq7nXsOHCCP+H8oy+HIXOdaUYOT3XHi4yc9NfCZcWE
CAwmzbtFW+J7nAknD4EU7H0Ytkn8PJRXiCXqSOls8dm3PwdFmWSxJFBPtwhhb1WZM+OCooeioWd/
6td4XOsq8cLZ/QE9ORTEdvooIFCmCvw/TKqkPU/mbv6QtafzQGt2EeD/T8O3Xz7hD5vvk1wHVZSZ
18c/c2e0DGvrHYB1Zx8sTGu+ajHRPhgoAU1p5kfO1W4SRebsUmpS8h6BBoxGb6omV/wy6eky507s
7V7YvNKDnYdmJHMj4NG2VEYevXn/D1pmaqv1LImh8zRP4aCoSTULAfsX0VEiTA1xfeVHaSuAwGue
SUdv4NMy8crnxuUEty/aJ2ngMhQ5h6PWmFG6uKyczEpeDYluwtyRo8V0a3m6nuR/jIcfeALQ1Qck
kdvlw4g2IoWRxBfPzazNh0tP/p4ftBF8ca7aSFN35KeSDUdmhrCvifTnw6DwsdTua0AHuU9DQsuv
k7zg+KjUhsjEqcabjPY+ImtmQXrobIJgEkxG14gRKQxHQ5h9e5i+iyFbDDFiudlxZlWHBx1ZcvYh
qdBbN5rIi2G4Hh7Lnfthy5/KsOuo1tCwmZzCxnRxDi+TzSTWZzjfMnLdRwq1+8SZznXC6gy3FgDR
4Z5Y4UQT2cuDI89aaOiBA3CaIyBtMMv7wlVKRlVYiyXVKBeJ/a32Vy+YO4lB6vFofvfPjrTavUu3
Pmr6/HtIipN5+PLoylrDt5ezTlZFyVauJJaaaDwdHBmRPTrUE2cd0iPFo0wilhnbAXLeL3LVibLP
qzn+LDC93sc7zSRSdvjde0QgG6dIqzYeSo0b3IVgDkhLHs8ORENkwmivxzbRQz6v4aMNzfU+ftMK
PNBr9mpKGuPeGz4z8wnM+S/p1YC0qRloOQOv/WeCqMW+JUhK/wtIspI7u5HyR3glFkunztddy+AA
u6i0ar2yM2lY8kjUR0FuTUNo1wFAZGGuFqK/VC1/hAy1xmO1oK3YrLx0Q7RIHZisoZVd47PnG16t
jKCt/hSx5veFbyOEyx6rG/ju73aFKeMZpqCZIZS7TBoTVGbYHDs78TUyjMnjZKgZSxQxQSBwPS35
n4ZyjvQjyYBqjTnLSNGkBvsXifhG0jNMnXm6enDkNwkL6fU/eGHl9ZjFKlFRIDrOj12ajqmzwOt5
aNCO9P5Z+AT2Xbrnl9UmTsz5DmdbU/6TSkqC8EakhqkqelnynShMC4uHFMcvzenh+3E3UclxInL3
kNZQ5t88ltVfE8LQJve+Jv8LH/9ptPlTxP+l9aokrBCQn6L+7mwxpyttOz9QxPmCJplblpPcv7XM
zJ0OMuXYyN5tlMLulqLkIKxkGjYKwhdC/ebi0yh7w9J3O8/BclaUhucJzrat23O6QK6CdfdDpLRf
ddYcyw7BHpHRDoY0S+qqVB0NULsHEPOKK4gb0y9gnR2n7u3Sd+D55yTFYdlADsHteYY3q4lvxRML
pVKpr19qitG9YUyZ/jqWldYrIioJacnHlC+EK8yTXdZ88QK/8SXedltpw9Tj8wu4sXFsoLMjXq2H
b42zWJe92UaZEEZtktfrkQ1DEfrlNhFV5Mjx8oGv+v9V0A9mioFtVfNcIgDmfTfeNVi505XqMcfj
2gCroA2+AShXBScn37lvlej07ijPsIKUxSJRdEZzHHoXiBD0YlCfOBg0wTpiGvdTTbUEdM96hlPf
B1d0/AmR/+AR6GxQf9boBjFpjAQJVnjpp2pEQaWLTMxQc7MJ7CYZy6gVbVepZxEJ7V70RSIa/F/B
/kMnd7kWYxm2f/LuiK1HuHWdFHaGFI5unu8+5p+6y7oI8Uk8S7elv+dzc1Ue+qHeGts+xQ7fbL8b
BiMnQwkLLCVOvIqPzQgCkT06LwZL8B4+ztahRLK/05kFZWnVgaCPgI93bPaoAc/56LzszScv6V3+
9GrcowkbFtpohHw503Pa/hX2DlzHXEVWjDvOUai2ytBQBzQkhVH5B7DUd7x8EQkU6Ip/nVt+DA4t
x+xKKfm3XTJoTKu7A5cjRJzb5E5vJFh3mTf4lXePIPpm8C/5+Upel7ZT1yOgiyj/kkLHHvTWSkK+
VygpevHqK4LUIPTr1zSST9GiKIAZr/6h655fICWrZZVo/1veaip/1YcdUYEOoH4b60IetIRAhxNL
XPd58fgCZ7eHha9iTMkE0JFHBbPDPl6WkpaMevgZRMFHqju8LqxYE7Ti+2ZgN6D0nbm2GGcJz3Ii
P1slduHkHQ0EojcyvyrBC7X4NMFy6N//BC+Kk4yF/RXcnv9pBw6WGneQ+mOsakZYKNrxKGgcOqc5
wbBRb6UqCDH0tS9AbOdDxIUnGJAIHvTEUwY/ZgQhwVgY+IY/S4R3Sy/E1i2HRq5Bu1u+WRT38ZAR
I7lPWd4bBoGW3zmWV9vLQjVgzGjj1yQMiVBLEmS6FJXF47YyU0RJrQIu1FlSjHNm9RDFMSS9IzWH
MYvfvvi9aTMOUkgzOp9CbwiPPCUeXDfPdL74X4mA4rE2Hmx2OY3xeTaqWH8v4/AzLmarPhOyr175
pE5lnnzOp5LsiH8YqzFYH2yTIkgA9FO94OFv4OYBzOrTquP/3HMxXHOBB8hHTaL9jlkeE8xnEDkc
E+dvzksgNvH9fOgurZ1U168keBNk2QaM9kVTacgP+0HumScur/VCz9o6545joRqOxXT0gSdj4eHY
+ZBXBws2Tb3TqkrfltjWWZeJWma1AXlQULmQIlO37NKMrLoJiQAvXC1rFlHJpVXVmeOYwKKf/AXF
KvX+1aiMHYd4ZVeop26/sE1uSX7oJ60INo/KBQAVfFPWNPvmQkSNOmTdcfhalo0TGQLgQazk/40O
gqarRrF64wDfK8yCeuoJjkcD4CjzhUSPaIWMk+I7wKkucFGROnHnodd+N+f351h4N9hAYjuc7sXb
F3cnfY1Ph/uBerUSBTO0FveJ5JwfkHS6m5TL8nvJULsOQOgeC95KO+GjISFEnoOqGECpHQsnK9nn
+rGMi1pVVPG5XSqr+U4Tmo16I+5wg4j1VGtsACjAMQzm/Yakl+CvkmkoaKklGU0uYPowlcCN6m9u
5sR9Qwx9VlGIBqgILhBDphNWfiXtmluJdD77DxoaSMN9yC4S8eGx0z37JlLC02PKudCAHYMGlxbL
v7LN1ZiCrVvKa6RwnSZLo8hkel5XZj5YdEN3KUPF+q4DwHMzyEmSS3qpCw/iRUAgnJ6euF8oh9Tf
k1QhnadaHmbpk2TGMiQViuRaEwW8K+eztuwH0OUxWUhBoD4YFEqn9AJySzbLQlsfFS9yJSRb2wU2
iY6jf/p3aJkioJvZgynJPHKF3ksyATwtpmcHjt72Qnwn4+OrMCRCgV3LvYyr4lL2BeZ0ABfCm+5E
7DO5eh+Qj0V0P8iJwRrZDjpz2CG9uDMH0BH0sALz7qXr4bulWWHU2KJ9QRHFROb4I2buFqX7pz4X
xPeIqQK/zGQyH90esYvHrzSa95IORCKndIxz6hfdOykniL4Xn5VF8FpQxUV7PGOTC3PYBg10v5bK
3fu1tuMvNWorL+idP/+G3cvcRIBK9UTHu0qvRwHkqV5/7OgtKKoAuO1WDr7pwTEB7E9jPNN0TIlD
IeKL58r/0idvIe/aXAWc5WxNfpsM8mIYWfxKa8dhYvu+4HHUw2hLWeqACaMCXHZsfSnQhpTaJEoC
73ZGylpml/OMJfwj4etwHBq5W8BLKo6KgzESJzIjp3lp7SiiG1r0oMRwQySc/IaOkgowfQIvty8B
dZ1TfUgDB7VG19niwlqJEAf8tUWeQXRdYRGYLyFEveEBcenlMZJiRi3FyepZIRWCSImG2nUJ05ld
KjE+dlPxGDEptw50SdUBoWIcrO9eFlM8nH9TvR+GPlASp0DOm+PeLbFqxDiIHftpKq03B4WF6TBQ
3fJOK3nhve45bBpOsbHvC9T2IVw8aJxQdtJ+/A9zx8N19HIIvvlOeFRRjthCHtu8/7Jjdz348ENu
3n8qRkuqB3z86IrwFHOyoqjsVaA/Gb03D9cpuJ1fzNXP1cVnwHitCIovDkq6Nc0adD+z0dPXMe8G
Pjy1r7Jek1G8AVuINaqyzKrZcwp8ZA92C6mJD5+elPrW8eZwRF00iIXROcX7qYOz7hFsi1mHqrLh
RuUwAXx+Kc8Xa491HWD7C99ksqPi3cU5ByqrA1JIS2Gk5sPW2eM1FDRn9egO7JGpsbObQXuiZ9Np
P2sHT9tKAy/s8d5lAPwsmUvSEMs4FyFVPlU+RYXT6gYesbltcqgU+MkLYxHGRXunu2HL5xmHS0Qt
DtIjjX1fmhkCLkEDT4Q+8LXCm/zkWMD02tnZvfpKDL0FgcRQP4GocPQFTMQw6KMakK3URDV6t4DE
gp+NYNYPky9kp3ohRSR8g3GunAw8ufsVrD5mw/aLs7o9egS5P+JwW9Gb7nua359V/zIfB0PBT6Ok
XPqqMD5SeOK5CSaa+b3zVrIzlpoFkroZKbkgSaelmQUirqRji4HtL/ukPFmoy4kppAXL6UV1+hoZ
lNMbeitkXhAs+LJHVv7Mz+ZZiXytg2rANpT+GOpWUW/Xr16tPuWFnVItWXATeZRpFmK4w1Jh7zUB
WB/DDuzl42IhEuKNmCFCHX9e1nMEAuOjB2GbUuyUiCtczlH1Qcn3WEPBe5T2+eAJ0V6cUKZMyJqo
8dr8UEniPLI13nyQw0fiMLyGIKADRHHdpX1t9cKrgzuujWN+XgEYSN39qFhj4SJ/k6Olt2H5z/Xw
KhG70ZHT7VIsl8k9hWPui729IN9UQ3bOc5jdBFwMghR0c8vvojtwSNb7V3aNl7pibQiT9/ugN+Ee
xSt4Hsm1inPL/smxVXqnw3NtsCYl4mtP0uJXwRIDA3RLLDFWNL3u4up/qpAgP2W3Ku4qSyb+vl2k
QAKkWWR4pr5/3K81MzvcpYU3aT5UHxJWEE8GvlAs9fzNrAQu0CyK/kSKL6Lz8JTcCs6PWYc60QMj
W65uE20ZCsektooZ5sMZ9msX83VBog9D0gbR8WXLftWH/r4lSAENf+7nTUiNHlpi2DYWUEKVONbe
chiJhTGbVWdCspsac4qrcI96+PrjbtHVoiH7h0roLrvgT2/OLU/JjMASNkAvTfMNbQ+eBsfoaxiv
9DHCv+EUpmq2d0Aj7ZC2niHHaVzOpbVlaSWTEa4h4Lvyos20qqRXDTveiGmtnOF/hw5eWQSYBhsW
rWAeuBYgu1RImf1JTyRVmRw/NsSRK9y+0STVRbCUqf7eA4WEL3kVJuupSTNxMi56uJ7ZFZg5rdbK
320d7A6YsjJ0uxdmOMn2oZAuKAUgjpXianZ4d61RkjQxDq1Fx+dJm1ivU1x1+KQ5zXkdFs2cHBmM
6YcyqnJnuakSDBie1pGexs6pBmtJst8d641RKQetPXumJhVPmwKNCLehkbNquSSst4fgg7eArlar
GloNWSRMFY3tvYT5ijw8woOiLCSYfp5a0cS30x27JxBD3GZOj/NVWo7yr5dVJV8R9J3GVnqoNRFl
PbIXQjiyj9cI9XU/hcr6iMXQxCm6QAxWAc8QcwRjH2VwcksHMkTuE5fRPPWEPfDhGOcsXsBtv3i2
LCckICq0X+uFRk82wpM6f9G7C6YqcdPjHrPErT/e8+i62DhUrWx7aQVeDlIGWIWhJ8lPQG1Tq68U
EYtQV6gUdG+ibvQOvnCvEFYyucYs7tHpXOVXTM1i3+3fpGxWJvRXJETRWf2w/ZJs+TtaQ0j4++d0
yOsrNoa9PYRMGLHkzFxaKwzkJcPFb7EyH6UHXWUpGkhMf/sgIslfCte/+oe4W43UkuVB4oE+xSo3
nAnAayI+mc21G2RLDq3avJztv7dIjMNe6kXKEMCWqkxOpD5OtbuuskFOkKRarYiUSFnm27C9z/Kt
UAcZ9YVmh6Uv3pbb03jjuyWvYX9kyIJWXxkcOY6JLQruHCHwzyBRurYvqTkFsRUg7J1G8B5eYqk+
J5OM/6rHQ+7ioPeZIQJltVVKz+CrUZE/EpQprSaTpbXISdeoez6MwtiOMeDdcAhFxJW4f7Ka1/bD
sGBa9JALE4CwAPe+FfYiCb1rR6qRcKB/E/95pG4TYmpHS1SmtXamTBcN0IZkrOxiASgtMkV8oOhE
COdfKlzceCwJi7qmPGTcPBXPYw/c5KM+haQ9z59onbT6JbdVpYu7Gjrna1j7TuNED7cd6d6uSe+W
3wGstjvmXZukCdf77S1USLsJxvQYCSggny+czz8GtfLfI/EhCSamzLlz9Ad6uQcLGGbmtzkQNCrS
M/bXyFzgrqSapSnAxkTZqAKPE63xSKAN1etpU1LebVQD1T532jKEMTaBSpuQs/iZmfIY3w6rOKjf
eMeNc5bB5zlsA8XqnB2UEvdajyIlEIoziRUj5VuSnOkV5IZdhSgZgRA43zop5CJ4YknPc5fj+DRr
HnT25ydI/3HH06WKowTk91MGKibu1LxoCvDCyhq3DEOBoN7lIWQmeHaQB7jginUdiVXNBskLVTnb
5BXQXyQ/RHeOzkcbGyA3K1FDdXQiPzNQyORwbIOUSXj9OTHbu1re0WZvact/WM0iLQ9d8Q9RgekT
aswPh97LK+ssVsYwaP+PVWzh0md7x3S6gARYhuojLObDS7UFrQ/jDrTUKcuMUgQh1VsOOPGmBkB/
/aYht9yWbNrg3QrUz2jJ1nonkMmDHVpFjGjg+6TmLk/9o5wNlLOxECKkIYGdFyab0jDYFIPV1DHE
6Cf3k6Vv701lRqcaQQCv+BBmkkFBHrOchFPtJuIL/oV2q56ljnXCffEYJ7Fd2K/lQLfoC0QrvpWe
8GJvAzMeZIEv1SXy9Aksi6mbgMFsAkDg6jLIeWmrbZ2DR5ybDd9uh4IsvuBwD4xBJ2H/LSNjAIQP
19Wt6BaNnm4sLWIZFc8a1ZruKnXbex6PrZJQJZYAQvpraaN77R5kEARRNlbCb3Q+NxGFBefFj/2j
roq615rBpANjAVj3LuedIMQlhL0pNecbptTlNrj63nT+dHWvKiHMxntuOo8gflXC3vwoTiIPlTXn
Zhw8m8K3Eo2trYKT747s+TiN6GfB4U+0Yt16kl1N4OSCBy8N6hoaHSbhxHAsiz3+fe0xHsvYixZu
/u1nF9SYV8WG2Z0MeTP7gZz+hi7/yGAgeZtd+BmGlYu6qHDUdUYzfP1GUVbbFRMgUUSqXEd6YGdI
CZZl6G9KA/g/cb19QYq+hF4WuP5DSbY17aIqRkLXH/CRbyddBJrUCkj5BwB3Jh5qX9iamnZuTyXw
dhoRc0nRUDl+/iWXhKAmuAmjFG1ed/bt2QArKPSF0sr0OxEpsmpbmFPT75t9W2xNSkDTSmuoRSX6
NSkGl5Ox6BarGdtEByWnxjPmoVX/1H/zBKeFqM9edhFA5rY159rEP6P24DJjzj876II/N6oEF+i8
jK7qbwdwe1ovqkkJf5DWGM6SzIdtcia/h/gM66F7HaiQZl9zGCJ2weptKnhQKiGtZYFgaBST/R9I
KXOLEHYxLOzq824bkDzIlhapr+fnIZjQkWuBIn1HvQWXIbIjsgpNz6LjaRf4rNn7ph49w13mm6lf
Zv8RmYoG++eU0CkCKtoCf2mXP8JrIa2nqGTLyRiytGDRsWPfWk10CaGNKjRGsWmgkv6AycIEfzVk
nF8o1tv7EWe30C+z8S3Bvd6MMfkXJk+7aw750f4LrRVMLECxv81yTEF8wpoN6+ajMdA01MR9P6Om
gMG3CyWzQCewXOeic0vgfbtcfQ9TLLrvG8V7hBHYQHZksYMFpN44VyLf/wRA0XRJzMRsjBaMgmHX
+3mla073YQbbdBsOc9K+7+eW/+1DJKraQh+E6wDSqtKwtV3YeFqbKw8V7OV26gbx1rJPnjWmeKsN
HD8MOhGtgmPJVtkZbLJqh0lDo6H1lKOJpapiNSZ62Qggax7UU09RhmrHgxUfKUpJH4Qj2iIM+e09
HI/iKpWdAJ7B9AsLczFClEgBPrIzhI5EziwT66Npol2eRoui2hw1r8JTiTOF6HUaf44DDjYbnk82
Dqvb+d4U7G1UKJ1uSil4T4HZvY5hghiDcZffwBDwRGdR2K3MQapX1lCAQ5XE+PWI+rqQK3idINet
J8pfmWtFVFaqmqzG5KqZ2dy8dCHaC7k8XQGSThHGE/jT2PwodsFHlGgPz9RDadDaIXrvOvak9CFU
WBrf/sRrFK9xubv9uhFvPHvWIyCyf+xULu77Pp+8hhfCAtln/KrfvUBNQWpcDB6XI7Ne3KuPnsVU
8gFF6iReM0hR26OZm0De7Ty0d65DWQLSCLPv7dTYzpUgnWwieitJfmU++KtbCivcpHLQWT9aCcvx
yw1HvGMFZIBJVUudRd+3IELZFIig+3UIuZjTiArBoxVTriUzn+QQwVsKdPlbRjlYDQLH3aIQcvBo
ZciF54iiZFpLsWtbV89NTk3dnWHA87V1A+3rebaBk5hoTJbsyvKNuHsd9DQ1BSwdUaioCpdcdhwh
1PbbkYX8tjrY9TYqVXBpRcfWmoT+x2xPTri5QKJxqpjxTCNzAkMrLuM6U6gcuI3S1W8x2Wu74zrM
MLcbf0BFs9j/wahI0SviRA7Lu98jz0oWYwhXKkjV0egnLPNA1gx+EOPK6el3FhoSXxa0svgRzDRP
GTkhC8jk+ppwP93Y36k8SOygXKx7vlxWzQ3h7FfFAXREvi0/+01c0/kg8voR5BR029FDGneS3n4o
ja3oLJx6yQlyBivZgmPQFYSx6tlclmaVMlqOctTi65SMc1NGdKWadZ9IwTIJfbrwrym9atIsJntM
jEyeTeOhUbQTp+grN7nIo18V01ovyOBosBcuHjdeqn5uzhrwkzUXm7QyV7heKejHuHNTFtVfewUN
/IkBplwWEYB49aCsXUo5F937RbXkfsymtFUu/DAFOvp0EyP+ajWoaQpaOvRhuvY2/Ak6hhK/PDEd
PNw6VQy0hDzamR7CYpi9t0IqU1mPrQK5haTWp3Aj/C3WOPTTL8VExBa7KSjGcqDIwnFFP2EG39mo
P9kaQGGQGmVOG8opOGdhB+rQSjD/rD3+ALf+8S+A1/6dIT6JtMx4Hzew310uEMqUmDj/khVAvJy1
mBxEzXXfb4Y87cMvMQN5QERO4x9Dih4QiK9nZMSbRqLrMNuNfoQdo0Wu9ReWzWA4/Tvx31CgL8Za
eKr/UTRRv9CSyPG+76EUghhy9xAhKLKI/tOUaL0Udp2PC48mW37e2/AYp4//MBSqwZyzaMVIPlOD
XWArgSIcQAMmNTFEXbM1byoSmVzGTHF7eYRT9VC+Etfl7QrKHsdV9CRIFhQSdNc4o6c/a5ZxUC7x
TqpBXqGFmbPNGgRlV0dkGO+bYCFeVEUqu4T06c77ecdQFqfnIo7WLW51whA2y4reHtcl5e3Uc/dC
VT78icAgsM3MP6JfLzTU3VljLs9qLMowYB/2pGUMlqLiGdK5QpFqqLfs5rVT7TgK8BD2rP7qN874
/+uXgjF9+ZrMpJ+l0b/n7CIlBw+Dv32YxG9OOcnWktkzu4wFkic3ueL+ntYt8Q7fT945nztTSE88
DbmAHphCm8bnNswJ6xMkrce50zXV9gh7WhPJKo6MCsypxm+VvXZQ5lOs64KFIIYLlXNRe2wywcQo
OIA6o5Io91gwcgux9u49GaqRuntMRzu5IGZwshpn2bO8aQuh2O08Q/2mHnY9GIYVNz+dUwBEtn5E
SwzZjCHq2SRO1DMV139pts7ZmbffMEl375VXVmDmUOLzcxWd5hfFZ65YPEGWnEJp/Ttg626RlwP+
eq5h7/6SG+eN3NakzHHXlOMmBGLwFgp6mXpcDS0PZ+IJ4kEdnjtH89j4SmxR2UGikgSEbJaySqGR
YU3LwgXwpvVDUHBJYf2jaxtZ5beXhanyxws6BY7JxBSjX2wpeU8EegmLOQN8YV1Ky2zXuLfHNFx6
HXMW3AKrYNCDRtEn7GCyBonetKS9Ts54RUAtEpPH8L8XFpKvhDl4QWK8rOq2fwLJ6YRgRFO26LnC
nxRCNnmQZRBz6FSVMGsjUs4AniBuJufhOCZ5+uaY6eDilndkvPPo4rDxRHU8wvn1+o6Z7sC3XK+x
YdjD7IUcYwIioIMtAimmFgpPN1G9wCEvqG0Z4B/paZsTD4Z3e3kbmOY9b+IBI4atQj6ZYmRH52Mp
AxGh3E8dnGgiOc2oWUqxXKdez1ZObXYU9jPnLqRJzhvlpMFF3DnBciw0Q02sah4JXvj57M1j3CQ3
yzO/s7e2AUn/U7qrXPnYTXkP+0al7POvgsYkCX6+ZOG1fONFX8/LWdIPTJ5XFJBuNlz8R+I5MfHc
Lg3kT/6PvgTOMiutLQzNu39iUABD9wfMi4dYlCunTZw8yGCGkGNxdqrruB6El3AIKX/B9VeCEZb1
mQDJF15H8X1hPI14cVB/ccZSXuDWgyFdhFmHFlrpc7J9EwqfW/9cazc4LBPBD3z5lhnMVP+SRqmg
W1Xgwyolea7c48e5SJVNo6x/iRGXoQdOYXxVuNe6RScSa33JNapNI+QGVND5XlCKRwagdR4xy5mS
NeoEQ/obN06Gh21TQ8amcaRmllHzDb7Tb2RPPw68IRwrm03zWlXJ8ctP4L/G6cxKE9e5LRau2vzH
rrY28N+jnZjfYGEVr6TSI1OJ/kxGbw2YuuDyLHECYYYVPSJO+Ku11MV2Q8FNoQ8gL13sXgAwkucc
Jlg634TYEDbc0JpPMbxy9O3fxlyq8Zx4cCjwbknBrgkFi6uihrEaabGT6r3fInIdvQI6V3lmQs+e
0wk8UqXTlIV3slCyhofEiF96WtloeKRXRKylBX7KTo4lVOGmukfONIkjZyFT8lp1Sq7ZZorltzbC
nKvAYMHF/Dcw0XlsXOSnJ0zf/pR16d80FaFuo+WTcyVSr0bkIq6UOQWBxK+9h9ypOvjvQJaD5BHm
rc7oDfZknDRXuwk81+r4QlHTCfokHyVguvmgFIxRJWQGq/nWhGCwmggKPykb8uMeSaeP7Tfk6bOT
8tgewCpiKoV5AnyzjmIADpwDnlu0fNsok6LDC5oYkGyJc+PEkkhAJ7tmEJnJ0G6iymLgOnP22Gwv
2bKHU8TWqT5X0Dun0xsHDyUbSGSEMmj0x52zXQXTxaz/CilO5qfzoiUQCLcyRK4K7hgECDDAHZoG
sfql93B6yYTxH33y12NTy0/laL7lZzKUb5R8OoJDdIXwNOvAFp1rCLp12QQJ/ASePLzLRg6M01J5
bWEegHESkAwpWkeZAV5elZaf+ftKpoxUUxJ5fSKalXr6JH2WdDK7E/tEq0zh5vnFOfZrK6K4VMcN
GpEq2hCiG6S4PW0ZpLe3GNMf4n6I0QDqDdyOV9LEB+N60HdCQQcuoc3dQFavihE8Y3UGLCkwoJWR
8w/lmcqX0SanYQkWd5qWHN1m0TYH6ltj80exDV+E10gWX8tdx4esNBlekZs4c388IRinCHssIjZj
OP0yAz9XKmAS7Lj3OcJGINKP0Tp+iDGTscOiytAS58wVFWiBnEaTSfjrjniTQQY+hSyIEM0fnRIf
ATwNu6YfjrOsSMrBbNIhqqVfdgveRwPj5FahO+vz25Jy/fKl3rcQ6HEjsRCkztScE8FElrHdos7X
1XJhCTfUcJTse0ARX5crQOExspjlyXC33XdGwkJwuNItFj0513ZkVCpD6CXsc8eKEowqYTKWmapK
N0DG7aJDzbbHQt81ahGvxadhA7idtzuz8Qz8wjc/nVAz/9yoj/RCy5kjLlMuafEy31Lc8sAIdQkL
8X6kS4hCc1x5Qc79snMGAkLAWt7sYKDKY8lflAcpvRhqcyN/xcrRIe2beH+GdBCqCokltnP4XMWJ
TOwDKFedBY+zp/1+XPtdAxveuTy9TYBZMyJZVtVSXlXicKRJSEPvjDHwpwjK4TeSTIQmaPyudz+Y
aJJnrvQeaC+1crj+Hkl4/T8NHDgfBIcjnVUpF7CHNVk6BVj5ZXeJow+f2jmSGKnp6Tf33oWI9qDj
Gvh5L2szYFOK4mrBgETdw2rYXwq0WrTqCUGYJP3Qc22QkF1kN4b3P9Jdfm8TL11EYbziFP84AvEs
V/A19TQs72ckHAgjHRltI1ILBDxqFxbfvSHbFEHBgkr3E7pFX7XZq8zwSIut6/r3IcLZBM04dCNK
4uZpmhE8gIT0fYAKs6REa2uIT+2AkBnbywYRD9ATxTS8N2jvNXtamT/FBhefBCLj3c117lBCVHa0
X+USq4RlGkeIYfR8YHD1qhsmnqrHhcWSZkTpvfjBrIbfaCKIWLhRzhhPomPUXop13nB5WTYjP9j7
7EYgN2gsTk4CgjK2JW+wPHgH4huuytXoI5u/95P9uEDS884GIxb4Snv6j1DKL9HTXS4zSecc/Zoi
2kU3L8ZVQWIPHaUPH/ShkQJLuQDYy0BM7ko6LxH5fdnblEYtdOuWIZzFJamNNlkUdMVujyastjEM
1e74PH7Sv+FQGObLaest92qmh3qXsRYG4moeqnc/EM+OepkqUqucq20sPLmiSrzH09aK0WbrZsom
ec7LyJhimWH3tC6kp6/tJXfGWWjyazHuPYHhfLRhk8z2a8gnpwfZUIHYysiDTeJcTmXX32GRid+k
rN+l92nM5F8BmgPLcuilkhXo7Lec0MAEYEO4NGWMQVTNqJUslCA/J+/0719UshggmhGhNvnBp65N
GVcYjmMQ2xoyyejqUoagb24Xc0+GLNpDeNSBFVI2mvkuGmGas7Rz9o6yh2dZY/aB6vbNXuT1vsog
rT9irLlcGJTMxQkbvxByJDLZtjLV+sIOoXcQgX1efKUbYxIrmfVMOKXiTHwNXkXYxYwf8nnV6moN
JLzREOtJ+j1h4d6Ki+DPbiv1eMmeWq7Yuf1EylwL7syWhZWROrsubPdtZxk2orkmmdHvQ1XSVZUZ
l170wF5Jgqb1+LTd5RBWnqH5qz9eYJII/4ceAylSHVrfkggLdRAFOV/mYM0UXK3T+2EOwj7EZ/Xd
55zy0IFLpOgkIOAjwUxi1LI9K0AfOFBJ00ZUX5xniy/an6Lip7NXCS1IQPebz3rcJIpKt3P93MoJ
Mx0xSsSlu8oe4h8jYvFpjspH3gTQJwthpKm0HuDBGa2rE21Bcdoh4VMaPEMlHBU/i75lvWiOXErS
uaiaG7P/ntQL9m7cEXzEHcypfRKhl6bgRsDDJ7TgSjGVH1vMjfsOwHnDcTqZyVDTjewOIyUntuLh
dDf7yxJRZpgtCbH4mzIJrjBE9npIAf4XU7cGPOG1vejdH+IKQrtmhEJ5YBZcv4hscF/yMVEnKuEG
OpjSKQ9EBDvAQ0Hdlz5ocpxJSubScsKZkNv0UOCvyoAQWCNnzReEF/A9B/VxmVVun5vIWLToBsMv
n4B/vCMrJ3277wCJcABNEjTGTDtiib47FeFaIm62ZWUenIF339oKKQcK56TSOwpYkasxxjeMkj5t
yH4ZcnRuVKO1SY4XTXT5FzfkcGye1Z8qzQME4BsHEPLBE6GIPk7k8BnbaDfIo/iQL+nvBmCEK98i
eAr0ACnn3Z7alEOUDuc9r2ZA4cS4AKlEVhM4/hi9VsCPv203FW/kJj75f5/yY4e4gpaBbJtwXLjv
rf0JBcbT2eUqtgy6fdArakHjwxQ2GEuWG+0oY/7nMdY9MoJ2FjyEM4n/0KJii8yI44d58RbvU+ao
+wUnUgmBfzkMkAFpJQ6SpgmRlFFDpAru2yisSWJr2OMNptZaTAnERsitqiBHD0efdDwAWvAKcT3O
qPJ+qU2GvERt9lzHIE+gvSGxmams6CcJyBJkFyEy07SN951HqZGhIwDE6+94H8V5g7tWc+Q4lbvq
HXiLO6PQq1MjmBv3bZs/2ucL3xKpizo9Cw62/8Y7vhu1QBGYl7fjDNOxhkc/T2aSdxxg/OR9Zua2
E2QgG0wYf6j5WyTww9wcGEU7VllLbaBmTRONPKVv4+NMYfAmmI70FzCq/ziV7Ppp2HABTMFNZK4t
/VBLBvFyQEmiCU4haETRlAa30iuSSC0XhmMQF4I7UdpoN9O1rOgl1UjbciOVXiaGmhvDgI3wQ1oZ
BCOSPRk/5PDljPoexs7rPlQyHhgnWIfPE1HCHDMiTv+j0hjuiOGDf8jr6mh3Gk1DU3G5ePPBP3Et
zzgMikazuTNFRC99ObZ3ZytWxaESHsyfJ7jbyYFxdRQLZtC22Hjo7JkqRJh/5eOq+1wP7isxRoW0
X5KmUa2ZKSAwpfeWS8Jhsty14QYAhy2oBRxviQEcdAK+CJGKC8LwifpQDjC9BMv2ODGHY2gLYwbb
ac0QBsm3mPWayfw8j7ui0/iL4h1N9HLErQEGb5cWGLd8YCFC/uT141nE+fUywsPQrNCtr28M8qXg
SyIzHC9pxEaIfLgTceQrKhZWRe2HoE3A4Y8MNmSsCIQo4fpGHZh1vpznTS/5Vc2q2xUwBQCahqJX
I1yQx/BQRMrHoeOvZgu7qQk69wHxvrNfTg2eMJ+SZ8l8PfMA7DCQEN5yP578vBHHPzK48VGhd5fW
RZ5Zqv6P9bocrDJSnIBnLX8WzGkgGsBOr5YFN7YElSbFFlJLGhiXxXvcLdjQMCBDOfBlXbEsvSrV
zlT1Rm3pdDuyczhdnqVgJmCeOMlPRWZbHDyhJT8icy5Nr6KM9GG9NYBVVF7///S0e0SQL6loCNDH
/BbFsm/xhqeVYp2zkcILtSsHyLxNaK//wNfAEVKpItv6BsKy/9EtbBstA6t4jkYwMx+6bDNW9Q76
sPVSb7fADfR6P3biy00mRgRE+63h/j+iFTyDgi4/xGrIUSoe6Zz2V9dg9STW4jfoYxVXaDxltGsx
MVAyUXINyrZuwZOlc4PduRoq1X/kZDBL2tfuc6ZTvWXci8oW0JxTzGyc+OUl9od9oaLkEgyVyJ0s
PxJ18y5TRgCQmKlFa5Vp7TH576bsrrHk8QrkOOwIVMLL/Uy3BJdK1B8dHlxKsuuxJpcq//jr1C1H
YFGiKELZUYzU5OC0F3b4p7j5S5PB8r6wDMvt4CK8MoNiE5W2Sp3/isyYp5b6gFHOUqpNxGA5Be6j
aDiSSMBV7vAdT18AEiLQJORQ3NH6cie5TMF5qFiFE9zE0eJEDzFL3ImGx36125L+Bs8v91+fLixS
4UjJHJ0DwpINKloG44udnMCF7248mt9epxtlW5kBkudE3RbPK56yMbYz3VYfbUdesA3EgHbNcZeq
fDnvxis1K99KbxgONTsmyY+XN/UcYIRCGG19eit8rZMvjbSoprVuEpf4sPTdF89MpX5Yf6dqfraf
PKesaIbpuk9PF0R55NU8nPdb8q1Q4S8syp42kVp9nX6slFLkwJoDM10ixtt+Mm2Uqxf9blwABYyc
SLmLcEfX6yV9U+ZbUyebR+LPcrIyDJr2KIR7lp2iQx2C7sPycnKUAmOqIf8jWL568WR5McvoDOEe
tF4lvo8AoySJlKeeV6HVR4z6u55d60picR/rizRiPDw5XcrIFoxFARGvQUqDhlFWnTTVkLrAikN6
u/Filk1bK9WU9q2/ZqQh4f9mk6nuXNSEdNfZgGZyjezbH0IsNkhGKznPJIVjLw9V0iV+hCVIj1DN
MQDgp4Tgsu4lXXH1txEoc4GHefxKUrlpQ35FbqvzaNcvf7gM8uXMtsAx3qWWXGbxQsh3R3rHng+F
S/KHd/zMXZOIxdkXIAk790yAxkN2WhD8vBJAToQ+KMfNlkqORCN5gCz7airGivxZu6iE7B80GoDX
fLER4KCzz6fs9h6TEenk+bsJ7Q2smm60yimNLsdq7NNiztezU2dmBx+WS3YF4c1hmdF6+HanjEJd
wJRyG+JGwmXinmFEU+3dSHtfO8KfDREVftZDQCEfzu66azqYlJHtOcHcYrd9bytKXhPhkHeg1gAn
b0fQszqyDO7fnzAD2tC87iLBczz7CtI15alWAVMSFB3d6seERfZD7o/tygVSWNhmlctOrj1CeoD4
oyufRtuPjHk4B3OkV6A9QaXlvhQlMXVtMzcJ6lscSnb4iVEiZ3otunUPWrNaI2hJ875ydGBax5CC
bosLuxcfrXa93C7wfskajvRGo4s5DHwnHm+F4dUU+67HpYRmSlBuoxZoQhl7DSN6wZYkNcA6Quja
s7tUrpEnmRLjIzG903mJQvZ2FPVvTwNpWmqtGDr1vpFHBKHSmpRRYKE6HUhHbxVyobJvwQSZ7Lw3
dhemoBv9xZjfiRecZLFug5+v3Hdx4RPUayYiJEIPril5uuH9ibn7WIFHSGh23qbQUjCfuLmw7yfQ
4Xps7gfOcKs9raVi4NokWjJmNeP7IPji9pm1+JCluIFRJ/Sx5jC4k1IcKNiS8UMx6B3JXGErYbJy
PjnaM+T0Q+a9eLDKhhVmzcQEqf9LAjVRklfEInXCpSt9D492AU0Br+hHVm1ijN1W1/EvjtlMn+jW
0PcutNOMezzJNLnQTsINUBIYlGkqw/FxknhRtmeTG7pSKSwgs04ks4SduPTghkSmimXGPi63sa8I
gDKdnFEVKpychjL5eCwrb/3euBWg5DwYV+CaoMm4k/xUykPUYrPapuutm0TWs95V8QhCuClT5kTM
FPt4q1oK7vFxtJPmtL9bBfoy4oqoUxwAhT+O8dUM610aLoB4PR9RfrydG9KMSr3kJlPyXM/M34Tt
KbolN+tYA8/As8U5INCuAQo659UW0Shhrvu0ElvGciTIeaj+WXTb6ov73p4yR5i5JSAvJhkyWFXU
YAN1MkXmzfHcxrPhnD6bGlReaeloGYOLvb8TDS/8mcDil07Ag/cdMhV/AqYguv1TfRfoisrFmjPI
T/muzniXXnk9xJeRxaXUVpcJ79aTbiuLGVUqbYldukL1R0GiwTqpoGpm/8g3lw0EAIs8pmP94nbx
9jYrABlhhM9aePhBnSafcXoJjPAOv7rZJIu/2FuUs/ms0V+nrznYmiSJ2V8Tmk0qjMLtNPZb+gYx
bNUO184NWOj3+PYoK/VSEFUT/kdP2PeqiQBMr1vf0I/XdLDskimax3bddtjrNKf8LgJ7MbYwN6Lk
4pwRTJB7kFoC00cxA9KdvGxI6OPr1aii1X3JI8cG7M9NNdH/evYLG0gKvnNX00d2LlSEre8H9Brz
g6c3ujBbp6xltWLYO/FF3CD4cSPqysPd/5fGNbe6XNS6zHc5jpAKdcOLJuRrv/2Fp2l8XDxXCOwc
/PizFH4Aj4tH5BGF1r0+XJOGXaw+Lgn3asuaJxKqwTdlg9m+IV86jDi0Ut8RxDNnXwV3JAVx4xhr
+Vt7ub1XiIDmCuTw9kk+KKolIA5e/xo7aiFDNek3wRGJ4+Fb0vYM+z2o3JMG6I+NSlR11T7GHY9k
opi/P2xa1cP+we4fz1v0fUBWE/TKnkiS9LJiJTFIVTYukEUkKWQ7ENmp2mEKNPfSEJPmnVKiF1FM
3l6HcjRd7INVVyuARA2EmxMQeyUyH9Pjbe6hSL2r1L7tc9LN+Km43lhluQn2iXN/+CehV/gsCPzG
/HbuZXt05L15+kn/5R+HEnslSnuiOMkjOcCSvWq7JqipdaPDCHlQI4kUEWsKjgb4FRPCnNaT/Khe
gFkPaSUAHrkKaOSNR0pi/6IB78uu+51L25TkUy1YwkRPsP7Z5W5zsWOfWfO05qntG3Gm4s/5Dm0j
b0iK6GWVMk9hRKpDZmqowFgO9ZloHuQ97tIU0O6qXRp6zOvaGeYvZSBjyeQNJzLza0LaCmgwt5wo
5Hdi110vQqO0t9zY+V5dQEfSq/tI0dADivNdHy/KHcqt2zrju+jm17M7NZt+oILaqTkkUDlOJEqR
qCDInxroxvXQ4b52WFVFJ2DdNL2RFhmiLTEi1dxrzGlDnfqc/wuJqoMFCBlKTLln8ObVv45Q1EPi
h9uAKJPgoX9+9C34+4kUBzGMYMEM6UihQGy2mehVGuZq8J152Dk//yCclSZCZ22//e7fmp2M7r2d
A3YDjxRT7v/Vy259cHt5jhV0x8jClKvPv6Klzq4bIOaNPTcAhawhL2I7y8EVF504xzqe3HewWF4g
mocKIs4RqUsRVnJgzc4dAWZrhOHOPOjOpliucQGHM1oM+jFpaqzukrhTuPt9EHNq1imYuSBbjq5E
PmdaoEpoSToDIqS0Sdy/6EXiW0sMpUcnbTmSxrRnqa1Ssf7aVl55V+rdH7xKJNZjKloUmxuJ0caJ
4bWET9sv8sNoObwisnmlOUTH/cuZrmSrMhVK4OtJdOQIk5+Xmw8zuCk2Z4DJx7ZwTaIvTxmBevf3
tDna5auzX+mLTnBB/niiiGEPyZoW56kx2VrCjIwZFlf1sjqb6pmZooVkFxJ7GRrcQHKLV1jJAlvP
kbfi3PRIfeFh0tZuGbDCsryS0SERk9vuEGVAA/toerf1FRtrEZQ6Z7eE5rfNybUmnmOObDBJoIoO
DlV4lyDin7IaThkGihSCYk9mV/97jnnDWmoqTXSxZ7X4cMquHR/ebsCmwCjekq1+Ub2/+VEIm4YD
mkEhfYDK8ixlD/wj2U4tf+58E+DMp+rjeeHehKtRg/nJg0/noHSPMdCZAHvqjvhDEEOMI2RMNPoa
jNtg6ghqXJLz43SN/2+pRpGa0v3wuH0MN5c0yBJfGipFyXDTbHZz+l8kowMsBh/rfLwcLyIbG+Gu
12Rqh3xOffkKeqc6Wr+K2igLR58+cgALkrt3+i+SAs4OIXkaYazhC8ubAd/1A0DyIAuUiAvMmORm
hcPIAKlfjjkpaRC1LJrmzsVRr3LTRyFjvHFKW0c6d5sKIzldxJMImd6aAnPWtcYUaEp5eKi0cZVF
va4INtEUqUxO99BxXuavUoIbDqCInitQJlcqDkfTRX5ti/ckYlDFev4bQhWMSSPPi6LnyfBNqbqd
ZivHWGNAgCSBja97J1HGYMcXWZY1tPFyUjRkuyprdrCMezT1QsiuhGuDKiGSAJMmSnse/aD48T3n
LLHOcI7JIB6VpTx8W3kmkmYyQHwqmE0LsxLo0N0AIyQuSmEB0w/9476mZVca6JlIa6Wv7HV+9BRI
1Q7BSwb5dApOn+cSTaHoHST8wl3pqG55rACQhwzROmM5LadAkRDQTzYWZFyHE29ITygfPZAlC/qR
9FZZA0Nr9S0WwW3dY4ydDems9T/KGfZvhGOOYEEpBs5G7Po/javfsaa0rwrFrcy1IwflBKoSiBau
K71T5Bo1mr7m0LqYYnx3hf4vPN5Jy+VQdEQLeHVzRxPHJP6MfhDNFscJf+VVTUz5ztuRSJw8jzsG
n/nrJ2FnAJDV8emkeXrXTjONFRZUvAQToqchXJWmNIpynuB8aUXcLhVJhHOusRw8xV7c8AFBOv4H
tQ//sDbrEGHKJo5C2Ou7GZr1OiFVrRhAQOwX4d795gZAoGpgx09vg6iEDkaU72QJjpCodU2XMAbI
NHB0wFrwPpm2Hws1Q0JfgbOd5sHxx3JiC3LvxE6MP9BOrTdZNzGu0l454oKyiZng8GF3mP5W0MP+
0Jl/mZNURyagAtvKqsl1gOfD+pU0rJOqKcdCiZVokYHg6hHK3fqVKfsWDwLqtQMLWVlG4kW8MeMF
brCzec8iZTsnW7grGbWcaNoAVBKkW3viGgwJ1IzvK/vmpvQm9sDmFallJNPdQsvF/l5sI8RIGnpc
btv4U++BrGtB81+7GQp9sd3P2n6xwGHIlIwW2Znu2yAUqcCUx8FroiX+A38C/MQVAsPMgxEeDf/I
845EZ88L2TiXKzrHod6TmN8bZyJ47XijuBMijaot6Y6iyW3/HI2H+Sx+1Zd4SxG3uKekjj+rv4oP
qBchDPLvTBF2L8P4+t59ggofHFmnisLa4VInkQRl3R7fP+GQE2wa/A7mZ+HiqePM1VnOuX66U/rO
0r8Onsf37026dOo4BeRRDj9YI8Ba6vBVgS6J4snBKgNI9qyVaSRSqeYpZOsK+WM/PiAbPzJlOmsU
q/mvIkmQNW3aXDtk7uPeXPxPdPQXFdBm1nbt6axhI3srjHFc4kzpqoZNHhV7LCEfgFV411IUYH1v
Nvej/ME3CtgbukYwRSmT8kyyf7RljOYw5pDxo5GXjliZswSzvGxMSX4i+bDcYR7Pv87M5tEPjHA2
ubc70yFK+VLWyiL923hny9VEz0k4ssZt6HZsBhtA2csvAxPEJx9N4AITR6YLYqWt0lVB6hcxffcE
/iLHMlMLXVhlpR/quUCa0vw0NCSUq4oOGGvMtnaTTete8mBL7zsyPQs1g5xqt9USH+j0r8ZcHJZa
QfLZnVNJNltlN7HsAPWmtcHDi8CB/j1rTpSZj5FEcq7NF9+AYcyU5SmyFZWocBuZw7agJ+OIVIQu
zLL+0RUsyGj1DCQo3uwRGIpRYSbOVniXeXJXmySH6OPlbXjxPASYp59tltRG1beN9HGREuLM8fUz
iSkijoANw9qLizhxF5+d36vXTxUlAsa3O8XVq69Fu+1OB1eW434skb5H+5OSG9QeK6jmrxGKhPSI
CTsUl93iEJrYdKccRYcX1rDrhh3rdTbod4Ja2su8lkFsiPWK8ADH2PvPB+Xc1kCSesKhzqqBOh9K
vYZIyk03N7LwAu6VbNLkrqVKFIVUTI6n9Sk0tFARjfS2mKs3klxsS6a0exzNEBY725nHawvM3I+r
XvEP/BHCNj0eg2IjzQ1PhOui4LfDVQZ7ctFHwx8IDx6vZgCgmzjLZ/qRLZNm7W/wBaw2cCWW0SRu
OiN5QjQW6V2UzxaouG7/rCvmvfM7XmyZfAlKjjXNExqX6HLacCguJamGfM/yreSgRTxXlevtdT7A
AqIOfDNp4bLVlNpXb8Z9OIgTJpKLwzyeFAHhA0+PgMDmQT2KYgd20A6I40s/+Ncaw1XCRkkzTuPN
1HSK2hQ5mUNPIgwxptpYh1nw1kxu3UmOhkWgjqnOUDG1Cl0FwAt84SO1tk6BIwG1CenFV09pg8Lf
YL6sSn7whqgPt1g2zh8vTUEbzj7mcaexuWUHWXYvLhSXnaOfNf3GCcl+dKIONZvd6prbUORw311Q
HPc4ZatN3q9gzmYd3bIP9HmTvHeI4D2rjJbDTi2CebsXRUCcuqbOcyiaEFzBbTCnXL1eloMxm/K7
pCPxr+LnokDThCOevicjQhPVNv94xCC2eeDdY5mUIHM0dfH3U5jjuE4BgFznr8Xopv6bCuo2lDBi
LkranYfM2Dan8NnAyNtyclwIeneOba+2dlR2/wxCeFWkwm7UbSSN9ZkAqDykK4bqa4DVzxMaL1tc
PsxLrTmm0A+VCVJdZInNg9Lel0dBO4+6uKpcp0y3wzPZFDIGCSV02yVsLPVL5JC14Tdm4g88Sfdm
QTRIClU+BLKUgp7YpMeLyU8ut3yFp4Xhbc2MuUSAhQ/xWdGv7dNWwp+MG3FFTl/1M6YFQmyyn3Rn
Pmm8kr/gYfEkYSwEoqq2YsOU6fAfS+dzJNpfWGukvPvA1qubnAFQLWHKIKdrV0FvUlUqCRgHnYwi
pgURVbcina+C6uF5EWR0PQ1KL4jllFHReh1Sf7h7pi5Fa8hYjR77XhL2oulpqqiZMRVhWMaQxcWC
6ev7cqwxseS8LRNhDlYBXPPDN+G7DS113HVm4kHJWkx5BuOXWI6nitB+te54UInX+d1QQ8hzIJZd
UhE4Sk6HUIHhpf95xgGdoLDJZAwq/FZjl/wOyB07mgFIdcN9qRtBYP/q76tgiSVLD/v50K3PETNq
scz1qk4GATfeuCFzt6UbcGVVeTkXTB43P9mtIezK07z+CHOEopAGp+t+aeg2vmktUE1pjJWKwIml
kzka//hbSCeq8xAnVDCQZxXtFlfqCpFOyuqgbGk5NW3XV4SiX25g1azOjPwMxKXKAlBahfm363ms
tZzwD0qtvgX7RXJyITBn7xs9h44H8rUINXhHVMgIuKe0mnGFKcgPcjJ3ZkbjLetHtLVwgJqsWkLm
39zWgS54xHEXjode7xylXVqjYrJjv1T3d88g1PXjCO1ffBHbz8Cr7K1e2h3Fi1732cGXxnGDaeUn
i65qTxkOV7C/WdjNqRhsinkfnY4fycJJc4OlPgu6dHMDMG/ThdamOXGZe17gOGZcYQZiUIOFrF6T
hyCTNGaTDbKB7GYd1Y6SIhPxWmIK0Q1jk/8i8V5a0qTWDTaJPR4k0qby/4AyglIyg1eFt4OfjYbZ
5WsUBKxe6QpysiTtCBnmyZPY/yuAPcI2+Bzzp5cLZKNsnby3qrKRuMLFiQ5MA2moDLTNBTWr+v0v
Q/lAugjkdJV6swpnTILDgIC+H1P8b2QLXIN+JNHHYBtKtWDD8ZmCtUusrpsAnXNHjZdkdaE96US0
epZM4IDUN3MQ7IM5n4kIUM3Qj3NlyXgSITeFz4naq834d+MDrURSwKl7CLPE4X62uorI5cVhRREs
gU4AsIhIafKsgHJdCL6X8WdVutCl1z+Ni0XZgjAaIzTmwnWQJmTqDGtQOXyVTCxISPpD8IN7geea
gXtAoryKtcIwV2mwfwCtIrKJU1Zx0vUQNxLkTo/1LD/H3JFK+r17EjNICHRRXhCww6hEhM2o9+Ws
UMWDI3zykvrOm7wKtavE81g5BzrzoLsPKX+CzyLerQGeQ5UV23NrXRlpEwsB7krs4Ga5J6f0Fb31
DEdu4GoCTEmqfg1oInVP0QFmASy3bWkMifuZgjnNiIs+WqVwCM5OlMdgDfACF+jbjJCcHbHgKntM
6MZ4fOcPT80n5aEFs5rAMo18hOfF2krGdcJuPXg+YqYq8hKL9yfqJymnGW16o4oOjbNaMnliEIUc
JpaXEOB629pN8bof7tAUjJm+RrXwXs6ouphMaom79CkPQp+Jd+mTu7+Q4rGtAlyTEJfOgKeaVUWg
UUkWHc0zlykcABv0WA8bEmN/cNsFXiVHXA8/bVbsb/bnFfLbT138MF5RDLA+C04x5pxrZgyno5Ad
1kgPOjb9ajkiWj6MDpF/b2y+vANx86TfmdHsLx6dDq2+wQhCVr8bZaTUNbKyS38IAo/AytAuYBc8
EDDaCLNlBfjeJnJGLGZZozChvt28b1xccLFQXzRxxhI7arWfwWbpwjpv//QurMqJs0nZa4MnX3Zy
OSaVxtV+uMHHAlIGtwLLKFhHlzQrnmRe354zyWsRod3pOz/V3YjmR4T9gtATBPeKtrv43TWjo8YU
KeR8Nc0Mh/FOh2UJSRRqIFQf83RymUnx40TjldgbV2ZTFwfXdUgaWEGUShhr3c/bV6fC6mXdq9lr
Zv4eNTJhZlViGPHrpTbXLPWJW5dMFblHvYM51WJh1lFHQURAEllGaCJTmQLZF3W7+Cbh4C1/jmK0
WeuQpLzpcrDGw0t1wtPj9LqvatIHuqC+xomj6xVeL+GzdpimZdB5FTfoERJOGADl1Z2T65c8iddp
uQZZAfNbpz6ORn1co+39l7lKyDHHYGqhj+yiz1gFud/V/70+FiFczYelwkmfRfhVaaD1XF13HEWF
I4a7T+xjcQ3gO7542dssj/bhCxLwpzbt4WVJFbSt5AD3fkyz8LrqcW/JSgTksrYfxSoClpg0VlLW
8oxcjgga//dR1/UwpxJnQN4Y1aAp9y99R6/9nxye5ZhzIodloDbZ2Ut5Omh7DDDge6WLZWqB35Eo
NrpEkqxYqm2LC5a3EkymGwoDiON1UZgTArf+0djwrQSqNnNWfDw/pEyk7jbPq9J/jyjFe/+v8kS0
D4o3LfMW3ZswGusxty8byhgVjnXBNluYH+CSqJkVPj4GQAZ4D9ogv/cf/UMbCNKnidNW7Xxw4TrP
p05aWuMjw1lhlcQTCO7jsHsQkHkXc0WEnBmUnYXV8iH2D5z3OAkEy7DgzKWcSipvmBuWqxmRd+uL
KQ5Mwrdn69X44VoxAqp+9ut2KGwbcqHEQtfewEybAtcq3ZM3CCzeG3g3ow/ulvnEsercbokHEJEw
kXulmVRc09eutNttoEZJHEzJ+2WO463oS9kJZaT7/0J9VfjpVX/DHWpG6xnhW8qskpHFb1T62xwA
C1D/LzYHQyMow3BNIhlMlLGGL9aaChstTLQU5EUFy2upW3PgKRepH7mZrZXIlWVuLsRsK0mUmXAH
S+lCLT7TNvEMXQj1xyZL2nnndsfVHJwOUh2Se6mu1ZUihM/bULHovE+O9yYCkoAtxjVnn1pt8WPP
WL8o5H5QTM/snfaaWhWc0H8Vc7sm0e+J9r/9D9hQI87PBzUGnsq0FWlrxfCQxLDVDMynZrjBJmtP
0czax6ob0MgjiaLgRKGavF3y1MggbROWnX4AcRRxX7JLc2xQZjSo2J3cQ3CkktaWOW+c0bqf4UeA
F19NLH0fRRX/l1uZaZ/ZqcLnDLZ+75H8p/zsh4gThrG35tcmTDz/pWyxat6x/KMRBWPz/JVSmIvM
2xVr40CTQu9Fr542PkNtWhvJrCTHsxurQFdcyqwuehA1nctxnk2eVHsicc4zY1we+Oe2PveTj2Ry
bMWj8Wts8EbTMxxdXOgLorSVfcSPVzYU96xH1Hd3x0OY+o7KJ+sUrjU3WQj3ZB9OgGlq0Eo+b9Sw
WzqzPAwnMUVzCwImAEYEQ7GxuBsmMRdD1qLeZuYLRA9TchmpaKoNPVKbA0bksAFfvtMoCiMJbsXx
8zz/G2+0tzA12G70B0lsr1hkyKB3iuMtGAIxX/BHFLw669qrswX6A0YEIqIgQuCao3gdEHA+pNzj
PdVm5y5YlFsWY5O6l3//5f9b+emgSQ+1NgJhZZxoo0jMhm3ZdChopfRooL3UGNorFnyL+bxNxvg7
IiqUC+lRoVgJfxbz5+YTp8SA6FWRJjUl72GlX/P+udEEtIobvSy3yu2ShPfUYtORfVWTud1K3IcW
QbftkvmSi4ATEaUkXrrRssPcc72nEafqtj6odmTNn7N2KPy8PexGTrM2rO7dUV8+JOSqaeqh1/6w
s4+7N6HXlInyXN7PpDgQ4iuxJVnp+IuCC6bpAO8vrBlSRyCEuFRVnY6VbvhKGhmvDBYMEeZQk8ct
rA81cl4LLBZw/hjjhMy1+Yr5fSBEhexrUM1mo8KX8XIv4zx5IpVmsKK236Xr6KDtSY9QzSg1cxo0
0XPGlZGZLGXrJTn0X7K8v3FZ/0uxg4xBu8jVYbytiJIMuP6N6a0EV59w5jJG0cJAiBBY6MvUejAV
vR/GYVCU2+PkKOUYTIcgyse8pAoblQ5F+QvA5NrmjN5Rd9BrjOd19qwq8Wq792QPVylHOAeCDfb4
KlSspmFMeCvdORvx4iv/iBkGorPFInV8umSZ5NiFzj2tnj72VKXVaHV17oOIUUJCe5ZOHh0QfM7j
MS54peU3FSyEpbOOyn5EXot3QABov6uSW+jwbjYly0py9bl/UA+aWbE1mT+UskkAkT8ZW0AOHx0O
MLLBfnDLQNxMK9LYqbQ+/USoja5zin0fowzKudusQZhCSAzq2kGYgdH4HmEuHStruvnHipNTglKd
9zpqsZ+prqKKGuyTMEhnnjGO0MqOLmf2mfyp1b7uFs15K19HKG3mhCFTQoHewPAWdS/qpYvewQ77
IrYVAyqwn2nwjthh6bD/NWNxSGI3zb2zPqLVVMCGNFu7sdBMZJxNC8vd35Z1qyFAhkcCT2+inz3n
crE7Ff1xg6Ud1fooD609SIEmKmsA/gyXFPVTgAFq6E/zVwJQV82jZbU8Wo1Y3xrpaRGHiWwnzSKo
0bNECw7PScaSaEWc6ZEX8COEAXGa2h34Vuz9tzcTtijKdFtMavI7bJPvD/OSeBnCx1HzLljZ7Z1H
2uDj0YaoJzhGp41NfBaYZjYsWUb4pzVnPqGadc+kc19A1Q+BEMqytdXgbJz70OfgNCNOG18tntx8
C02BwHLRnP4DEJ8xfzStM03ZEYTTc3GoTlD4d5kXnzte2hQPLMwQPWeGrztErTDSoAJKPzEHEPUQ
77DRtV8M/K72AP1gfsa56bXgid22dI3w3gvLlG3iV/ow2dDNEWHh4/YMuM4vcmYfGwlQhqhCUAad
tIIYvwCS3CWbrUHy4m5WwEk+OR8EqA8XwDmmC5v4dFIHbBYKsiR9A/rKQQDICtF9nrIhhwUGVMYU
V7J2Q2itimtmB8VHuTziN/AhCYUATZX1LlYf+G0KvccaMsS+Q/TZP33bJbdxofH3ELHy4w/B7ZQG
+YBVyUVPAnzidi2GTtSpQCGKf2JapBbq11RcD4vz2YIusRWaae5OWgCm39jBGYV9jH7AgXLQiaO1
w21xWJ2HC3eCmaiGYcGGI5bG4/JTCBBTG7+YAytfCp0OikXFsbeW5PNZQU1E8cO47jzT+BD/6Jbl
5nXYchMeqdr/qoqSUONPQCk/ELB1tPqpdOz1OhOz8WCYMJO388w9tpPOyXJEBvqZiKbyUU7knxHE
PA9iB9aUmVzbaeqai1AFjYDHYrixCuY45eHc2zF74lppU1GDN1AvqX+d8LbS4j+Ae0FLM4SM4aCn
3I+I77QR316EBZwHO+8tvn8uEKGXgVdw5LZAAAEuOVY+NhtCJxoURwXB1D/tYLPq1Qbk0ODyxuRg
P1R3Xc9lVjyjcGwmP9Nxr8Vz81CvGCJH2BSXp7+kRQuf05rI9BDeLqfJB8zMVl+mkJwvB9Ex7ua1
Jbr6koBTiDSzhM9YlDNcbXB8hQsL7TBVdXrtiJBnlVQ4j9Uy1ocJHkgT3pJE85nAjEeTkCLN4wCw
wRn0mx8suNFvxZgc/4dn13d7vzqz9ok8zCWfkegJc5c6KShHnIKfxQSpRnPKxpvojoQD1fUYk7RA
9UQbwZC0B8gyy4jnY4N5qkHqFBQ8kwHmaW+43zIJW9LqkCWPruOdc70+q69rGzneJf5IBLe31Emm
PcdaL9B9lWtWoKVsJyt3tFz/x/l4Ic+tvN1GA3/WvQd3z4Ik8SfwUuOR135LSpodCcHFcJLrpEda
0dc+AsYMEM5UAQDp9HhO1r84Ux6MYVMlnLGlVSgsd16fPPiUmtygZ3X3wdtE3ezF4bahCTDO9UAc
RZcqFV6RjjNydyb4Lclq4MIRgq94xj3E/pXVzZPVjEHOEOWGJCnVZ7luYWH04FUd6ZSVesFmEHZn
mrXrKx9b4dfmnq1mHyKNQgFCvl+Jedf0vWs6vfy7DNnUXNCFxtfHcKovQFYhj+A7fB6Vhjpwd5At
r3GTSpMK8FgBlB4XqDjRVBApwE80Pxg+7x6wynuIh5q6E79CGXbLj1KVW9LEFe0BclHABUEF7BcK
A2RQrD/jlDp4jTAplHXaCWwB12xRZO5QTNA5RniteY8rpzReCrQZG9xgVmDJRseWJK8dA0jnx1tK
H30v1K215wihhnfeREoyiVQkKb99NfScBUkofIbjL0YqK7k07hTBozyu+rFIAuqKuwEON0G33Zyy
rS1TfF5kc9Xwf/WSkf0CEyAlwY0pcosDkRdShH64QBcDOFaUXTy0cG6bHWKlWquEKKPRSPooRv+I
KgRu9oqejOjLdkU2unjq5NF4rTXtGs+ODcAkmpuTPfk2cVXqR/HFmWNc3m4xNslOmXt0T3lfC0py
BvvSRjn4cQHOPLwGejnoN/O5uG9syyAJFXaKWKxMC/1GOC0j0GO4lWgtkbZtEyT7l31ck6usUYn5
qUsYK4ryoQm79timd1C8DgpSYtHXiQ7OYSg/7Z4nMb7IlptCPj2G5zahD/OXKEqq0RwxxKHCSAeU
bakcvwzrr/umx+7G8BtHOC3ytDDJzysobJAJw1Jv+QGpli8TRQd8e4GB0v6Wh7KdIa/f/hzUelV3
IpsI8qzh9cEghTbnB5f0DKVGJ15usvkAnnkrMPwK5Y+s66HH/CloajW3S/9nu5+tMNVPSP214Tkf
J3frJh25kMEuB5B3ALWm+08KXRHqSVO5DLZydpM/liaWZ2FzWldiXGxbX6W4B26sOrjdeoyQM3l4
x/l48wK1foHgxQCv3Zikl8a7FOAhc52jO3yrhnAVfBBfaysWJrciqBjBD+LXMtfa2piM69t1tk4b
BKJ8BzvlOGRehnvyEXp/hr/M5nqgfG3gzPc5AcS1GsCw7jf9CO9GOnZtxxIajglipkVbVrOymsqq
c3R/kSlKqLlf6rIXbAtZ/+0LtJCe3kP/anirmSsucPjpOpq8P5v4t1dyx3skLMgZNWAv416pc5h3
oY1uEwMbL2EFewWlqYjFZ1/WNf9N3hqv7hoDi2hTE93Pz9CgksupKwWVKH1L6hjUF7zPoBLxIx7l
0OyPkyTfCWGe+MljwJ9xOOhb4iNbgaowX6zWeNf4C/wR9dRXbNQhYXMPRGky/fpC2FgKWYKM0/NY
yX1fsUOMRJGYCgFL4nkzqJKq3f8mPP/a2NAAqVx2gHAAfTtGoF1EBXk9X3o8OD0Dix1DJdKNh01D
4uvtqoF0joS+fzO2C5gKvJc7nLNceZn3acgjfeKNiHr8cN1bGRaEa4Ih223k8TSbsJNclKdgFC2B
lV+eK1ThCbb5tMdK+gwl7XA3wuQ0kfhx14Ij0nucXA6YQ2uGFohvcEwOY+6b1pIexYSxRiwEcl+I
xsJC+Y8hnDJ9zfhN6TYRu+sfJ9MlfQW6nCbQ17Gw8LmDhcNaYHZqfcLxEOh1NDcdayiNVPYUT1RS
j+ybUyLyBc3+4CNWF76zTE/EwnfpcsPFH2WdihM5YyMkMCEkliWeq58Lf7qIqR7AJfOoQRE92JFF
mDRa9Ds60p55KTIe9hVMP0Ody+VB/2pSCeN6y0d2xCaGRFHSmn5cdQuMU2nwNsomHbTpw738nn/U
u4gFAvI23orCXkFEN+2ttRZ4I3bK19S2hpBJIksJsc2QD/c00ErU6k3oBIFi9Q7uGXGfbQonR4mo
7U2eK0bZvxuaG9dhjBspkJYwrxg++ZgggmmY1BccjWr/Ev8yzFYcZ2MVLsqJgZvLmoZelOfdtILZ
U+EDjaxUBAJOCibFxDbhZfKLDoJ8ZV4eQiL+7+BSR0pF5hv1qUUrDo0v22LL8+d4YEW/dcrxInRG
OV3Xc5jAYeOqeAemJbghsosql83tBu0Fcqq/fYYYMWD9403XPOMJK3oouPOa28IjyfNQosB0gdeX
MECZzfRWE4K7C2KKlkW801nO1CIcbjd66sO872oEb6uGMtTih6xayfSLcKAn3NNf5J2aNJuEPEwg
TOaURi4qolQzoRxHTMc47rhtGR43N8yX+TCIQyPZmowTWwbXHod8V481bftRWbNd73u0cjko3SG5
1IFLRQVTgUaNUopCBYVwbiZW7N8lCeoLTcN00RSh0G1MgkYjlK6YRNoUKPo+K0l1Ki1Vg3nIEZv0
yr14MCUI/R/WWD1hky12w1XtBKjLZwNuk3y6pO3MA0NOh4TzP5s4k+zgMrFKJID9l6pCjHn3Ub17
hXUmfA15qCs0fHKzvXHYMM+ZMwptUQnOSgdp+6TgSvVibPfT8qv48c42Mjy1t08ouVGz4ejtu9BE
nG7YAnDLM31NFGnoV7UooUDrKaIxuSJHUAl43PhbFnfadsmiZ/61mfP71hSKS3DBLiP0boOD8+Ps
Ae/V3Dhb9y2HWkav9u/kNvLMWK9gbEkUD9xOt+VU6xoPKIZ5ohRH01Hai+VHODn+aIRqzYceC4FN
6eOUTkFcg2bdyBgVdEI/k3JEeNmNWlYR59ujBbDR5nCVUOgITbEFK5XBsnN2hnGWwiLHibOFnnKi
gB9Vb+1neaoY1Nt9PJal7T1Nvqy1DDRvg7SfVRqccDoD5uSKBbB5KQd3IOSMrJDRaLrObtJkW9EY
lkroptEjy1N7upDNwczrrU+tz4iFCjUiqRdPAEb8qxtPjThceusPjrwoU0VYPqk9P3GPRrBnVyNW
/O8MAb0f2MQfYIz3XqduHYhX6tDhKIjBshwE5Zr87eKfyCqG1+MLzsvRauEryTwJxU1WgS+v8SMh
eKNDitu7k9uJb2OI23hIWr+5O8yGdARwFKYvbwpDuDSo2t0I4cs5062enl2zOpa1O2h/rcPvnqdP
K99fiNssy3pm+fAoWKz2NTyBO+DeVvAx49aX/e13lDKXjOI29WBXLHmrVCrTgIy/AdEx2IX4Ftfe
JWXPT2nqiNl+ijsoVuTwCJJsb2rkw+jOXS8inSXfjL0CCswPdnRHH9GPggIb+gy7cjknVqAfEVTe
rUy9D7WBm9668+6Yjs7gCXx8XvgX18s0PfhhwBb0wK+kuYndyXvX8oHQf0nD9oFdhcBBhE8layVT
9xaAGUHDJQihm+vafA9I5vtp7I4GG6bUb0DfU5sMAsaIIv3xz/z/lwpK4Zh/RUENn3ClwGaI4FSC
CMIVLEP5UkHpJ12RYg5AN0kciOlwsV/zznltoNTYLhGttiT9sjrlFNTHhsgkau6q1tuetMI0zNWF
A3QH6jCBxJ5qME5S1Xt3AcTmOlGPH27VSdFFg6FX7BG7Hb73jZre/4pMM9WMOZ3/7fZs97AED2dN
aOyFyQLkP/4ZzNMD8KN2VhhQoi7LRTNlbWra1YikCzWsxpD7O4UXdUjp5W7Ctqz8Dsu3MRUwNK0x
yy19i2vd3S94Z2ly924Y0d+aW5aXbP6ecc4eA4PceyDtLegjzoIR6VuYm1DhQ+QXapy6l0OjSsDz
RDtoOlnMkPyBzD6QpH/hGMTQoSPVA5hPPmygwSexpbs2dxMOFW42DEfY1P/nfCF8j2nRltr0ZAIB
oX7aOShNwrgNx5bk+WuJlsSTi5kVk8x5PpYbTfbuIf+ymvJWtSXGSEZSsBMNmivd8uBwL62HH846
ynZjdVDp5Ocb4UWZi6PZkTiEubon7EhMXkO42zD0dNmkTFEBIM3OUuDtqek+/eB/urxNAwA9E0KQ
DyZkF3o2MpsPpuCibFcc8MON2zBLgYo+BbInEnCvbmaTUnUDN8XQxq4cpbDyFSqWrgp9/ckE9DFH
aeeqOsiq+J3It/JQ9YYzrTPEBjFl916LLcJ7cFbOkDdIB5z2E8ROTgP0eV9bgCoHpNYY/uNKiNdv
apvWDx9icAkkEzE0dMIbAArCs0iGLPKJi+CLxlJqKN/O6/0IkUI2cNWTAuRPmQSq+qRDZVxRjfal
RpgvaGvw+uncZt1SvGKIUi6tSwxDhVcLZ/j7Lx+ol8lAME0SbPNwf8egN8zaOnrpQSMrwUQKgCmE
gxCTAvYPWxVK4R9ON8e3I2yZJGVJWIwKNKY4H3Rp1bXQvfGCE6sgPxr7Y3juI7f9Q2zhZ3a9zxUT
lmPxA75ulZapTExOH31e57/u+bif4AcaifwghUHTqWH8a/qv7IRHFREs9lHviFgB0ZKig79dNsrN
s4LulRZOS1xAHwPFp2OMRXruRoORfqLKgXyu2gw63imvnUzxexkWiAR/9a3H/ILuux4r3Um/7oCg
uSZB1RuTy0jS4RNKnTCsWKJ5PRu0yJ+AmSuCJQej7qfK398JiHZz04B3NgoFbO6S58VbDFqNibdR
t1vvPGplhHnnUyEI/6sGigXzXDpLF46YmKCfNYhtpyksS6LpFJBijmk9wjJ24AR3/vMiDZCMw9Gb
nYO69OIU6ID5YT/h4j/l3V9yW6AjeBjdah0syVB3lNlQT97sApaBI8V4TNhetSBZSCXj8DNp+by1
HJh1jykI5UyIhdOS591duDKDUKpUizFSg9V3EuWssr9UE6DYAmSnP32TZ3fOt9U70oZxsQgW1126
XNl8hTLqeKU2h3tst8YfEUydCiGTCGB4/8s1ybpEv4htuRfc8TfQ+7q6Tbbk8F0XyUQjMkplMpg4
ca6jEJrsJeeuFySxAudSdbO8t2T46+GUiy9Y/5xEIUdI8YLnNtIIsV3rEV17Sm4PmrdDnLlvOv+W
aLxkXpI3J14UG380JYP+2MbJcgC+B5IIyk93nrX8wPuBECSgDNZ/hFazRSn6AZ8oLYcng/xbGc/f
g17GJfsAkVI4ex2VyxemkaQZJqlsI9YlczoamqVNVLgLmSFICVqIRRlxUuPlQIquBmgjhVNkHI5Q
LcSaVGqDdzZFJPUgkIPan8fnPaCC6aSJEG1ja7D8IRs7ISLmYvEL/ihJRkiELcHo1XqkAkwzj7vP
iIJp6yQE0HeHEVLFsyuEYTVNOA1q3C67tbm9yvPblT0xq8l3oEQFprGobyxPN2ypJT77cYJYJJFQ
osUIwv3Ap+M4r5HvuTmNyWhmgt46YHXyxKXPuzRrdvZzWU+Wh5HQER2X84n2KNloSmf5cXGGbFmg
rdKZ9bpW7tHemunSh2D+Lfxo02e6xvtMHd0wzIdsnIkDc50dpLmtk2egJ4sRpCl8vaNcgFBNeGKu
UL2kBevIP9fQQz3oYYb80nEdecpZo3WBvBpV67u8A96Rh8o+J6XbAwUfXg71BR4S6k392qJVhp5M
uveYVIqzH00tWsGJPIBzgRs3qRSuTso0p2EOej0wILn7Qna/GJR2VEBC+r2vkjNPBrlXLoiDtHhq
S66O2qzKAj1FJY6s0YLGxuEpG+/9GnRn/4pwBSDyPfrN4n0OVQPWYFl+tNvSLl+5YNviw25XB9Ak
TilB39ZUcvZXcWOqgyjh6ejyOzaK5EBNXW5hAT7A6i5SpgCBbd6EA+o8d2Bue7N07E3BNugTJN+9
wnIowJ7bCivgMojb96TnkEqCZVp2mY3HxKpA8pJStpTzJcSHVT9Piku1HMRz+0uaXuIX8oYnKw1A
GHOujROelHSmzzBhBSJ5SVQLZfW6U6HJw0CvTs08Szy+VDKNnrWdCfpmUCZkPIVjLmkbnCtVRnio
WdgfSQeFT+KOKrkIAHRKyPGakxE+QkQZF65VbrVeZeMib3g2cSbW943c0cVGw/OyOes73NQOS4r4
Yt0xHAOMpVQWS/2dpFUxcs4/ioKKzlYFMvSqjeZ5ErjBa3vI6tF9h1SNbHtoHXt89C2+7XWZQPAL
H25B/WhvLgz8p1lsYe/uifOlDHh9+F9HkznOI4Hve1L9Zs/wggVIUTCBXxulha02OtyEUKZPicv8
PzmJSuUt3CLUl7T8cVKJaPF+YutyKIBDtnV89hfDFopVgCH8w7gT4Byx3vho3TGiHxxnT8+6xvPw
zAWsiGr2ljgKBhBkvelHCFTZojqXjrLlHxexler7M80M34dnxNoKMnUWofMePFdM4vBmzD6qKYTZ
tJnn1THGmKSEp2L00oDtzIFxXouYCYkW8SXGyxapAWv6TkTfsGcEDym7QGjSVNRzW6TJkm74EUyP
fCHPuxrqMi0hNTyk60OtcNiIWis1QSvaWI4oh12jlsaeUNw2LEBoLr1wzmEeUZ11D7q78zTKxM68
atb+sG4A/KczrYvFshR9eWJl7+5M5cPN52HSLbca1MSjMnnDsYGLOKEIeUSGDVi6laUjZsYW0n5q
HKHU1HXTikoXJrX9xz4dz+NZZRrA4gLVPbw025fUIZPotTQgcNDigDlcexnjOzRu0QXnj90piwOn
ee0COweITfRApmNwMixB0fA7AOezoue0FJLHQI8UjKjWiwcmUtdrK8DPugRzZtDzwpWi5e0hkWTP
YSsUKDTEqD1R2nIVMUOh6B9CNgtrvB7AvrziyAfYNNQhqtoMYFAGYJA4uQvGtoUvmcbqB6Uqroh0
/vWukUwgtdzuhFUBbW4ooumEtjs8kIMyg8xmbF0GNhN7k24Ejzl4QoaygesJsFa4oJJZ8fC97hSv
q4u6rO2EwbOrZqHrbjPx5Q5mdHf4ORfjRcL9riDeDvDTJ5W+kDKC4LG07DY9yMRa6K5Ls5+QOhVb
1wtt6+0wQZOEpwuCzC47C05Dotjm9Tg+oyxt7xuLp6vUrt5IrB5mDZUb56a5yTrmWayoDoLN6ZUp
cDP3BE9ScaS4NwqsM+e5pY+fuXeIu393PeUyufLGr9tomBAxJdFrnfl/jtp8+9f/m7xLo3IF2h8Y
e+wxnMgRje6I6lxdKTShFTUn3NxGDNZhWyN8VhersmQUmKEgWe6XrMCJEpdgQ5RV8LWTgtkPNBmA
tDfXVimI1n+HX5L13G4dJ8S9bXcjYGG/37vUzVvGhQVOT65gF0N8oYppgwtIu9KQGpqBxkEKqwS6
rUExNF3OxaRadqoBMVjcw1QNTrnEw2MSu9R9UGaJaUDyjAO2045O4u3xlEZXekS4vABiDPY2ql/W
YsQiejclycmpHaIS92kyk9UMxu8gjqupe7aPBWx98cwd4fz8TVsfXZgI1kEP161bIMDR40RxVTes
gHnQRFY1HDXL8UDjMTn2LJKnKHsOOOSTKk0IocGIieom0IJA8jG/TtC1lVys5v9OIYlbnuvUbVJd
uf/rtZxEoRz01XHHnb6CC3377WOHTwzQ5FpE/2unS8hJ7hhwQwfmYuB2Ds+Najcwrc8dPdnjWvLr
AEhnLKF+fzmCgw3uqMOEQmUjTv4M31wAOy/2P88YL7znC7o1ate+DyVzmyau3cPocHOvHJZVHbVU
lhLCV5Uu3X4fJ5wdisbYp3L29HZY8XBH3Mk+eFU8v6YtP7r5FOImZSdlcnKUeOGDs515FjB4n1df
vbwjOY2INh7cZmxyWDgyyixJYl4R+Eq7pCNNnVrjqdxyfKIJmRwKiTzWM/oQfaBhar6+knKsjXrc
Q5i7c3EegyB0O4RC+ZjXmw5/ynVarvKwGw+RYN97mVXo0Nj5B1UwWtkY3uVhZXPkFBUlV/iWsHp1
y3v9dGQNafJ6bFm4EamZV+qu0E97xirS3M0XZXEKVoVVyCxfswTigYWP2nWUWPYOyRERLHV3Parw
7Uizc/pxJSONpOq8YR8aJZ3Xp/Qyh+DtXN/ESA11GxRgiW+2iqL99sF+94HKRdxsfUVGRuZ0QaNu
rzfVGrJ2OC2Fe1zITLJdQbZOedjBqAEV3X/lvUdaQ9xxUb7E9//FpkH28CrrulHm7W6N3c3XIyW5
U0OiEGc+Mnl0xLbbwWQPOvpHd4UqdBH1VYI8EIFUEx3bZ7uIjR2dlxGRCrGKkUUIssDX4EbRO+gq
7lkoZ3q1bvyoXZtkCFW2J3JviDHHHV62vd5SAOV+0hReNaYO6RRsZuMgwa7a1sOLON0V+LpcJjP6
qoeaUJyWrvxb3qaxIJJeFyZrvLwOoavOr3ZubbvtaJ2l1d4snQNJJ/6ogQ/qld48Fr7YzuZSe7bJ
MNrYFtN6AKQxXKmr9ItDlP75AjKCj25DIeFbZm1Bb1RQzdy6V9OBebNKzsTErEAqR2wTNSLbXlSh
a7nLKtq/Rxk9CdrtlhkQfxRh2WXWbCaVNa53tJo6DDZFItEuEGK0F6wYHfUdBPGt9mpZt9DwLrL4
uv0rwhPaV+vTmTLJD8qSm5QDaOP+i1BRVF/4bEvWIr0WZNrFLeuM5dTKtwhThSnu4BeZkcoqg6PQ
lu9/m20eQOsJd5QT4DOv1JHWBq0wEpkQJFGWUL2wRj0zvAFS2wh2YKwe2OoliHLJ4iJCd7tzqwS4
GRqv6IINqNuutK1GfynDw2gM420JDoPt/tkz2LAdoQnSVqvGTA+cIMI5Q6hoUp0Ze9BSSh/VPlBr
y/XJIiKUrHRq8zX+RhbjPABtNOxbLD8JMeJzpTElluVwojFVJHbvVstQxJ2I4WLEG8+P3ks+dFtH
ymC1p5IJYZ2th8NE4lCmrJmOF5AG1fMucS+1506bILFkpOZ7tQS+Lyvz9Qtp3svPTdu/6Mcp6Pj/
ywBbhjT45EJHugtRJ0wPnWlqTOHrkPd5QeRm1/ul7A5tS5tddKVHLloeDYgDpb6lTW0GbFPPMyb2
w7stEoVNi/k2NccqZLAm6XdLjW85f1zpegrKw+JR7Ko8NBScU7lv38/6bGuH8xvcnYxnTDHk8VX0
N+W4T5/Jn98Cpnj2ni6Jh4hkiwKbO8QGVgJTM8wdxLO+yit0EDFCl9pqVkdEP2PBrKQCDd9/5VuK
oNHW23iavRC9SpSOFxzv+KuYXoEhhwD/253v2p7HRfTo0NF4pjxG4A5bYcpSwb/eJTJ1CrWxccTT
t+tNqEMB2j97tAwe1kj8vZWL/DbSzdiu/5qb904b++uIELa8SZwsg1RjOBdIop9UEhCZbM3gj84b
hLq0klNYvGyc9k73WBqw0lKfdkhsqlrAmjAdSDTrxYbIiFfMxUSrx0TcbxR+wwf1HStBEDJ/HKz9
ELjQXt0WiiQE95QDpc3YIfqwdJnOsEwQGB0xMj6VKW/4/L7YuB6bUBN9wZfekVppowp3oq2GJK3C
mjyUYb/BIAF4+hh2O07mk2EMrAJcz8IZ83gIC1o0oujEJHKQHBWecc8oDfa5lOf8EdmTcElC0xlj
1Euog2mwsxZP8FiFojxNrUFecB00GNY1ZV407IJbI4e0ufo9Sd5YKPj7Q5TBPV2bHIUGfp+0+qVF
3WAg4WwkqYiPVM2Jhv9foT/wKBu7CQoO5dpyA8aRciWuSCWs0cOkXqEQLX2rr3nNhvF6+FtMnsRC
0tnRAChvqIwavFIkc+W63E/8BLNqljvX3AtCRYnYYUWpYpJquT8SUX9HBPEYSqrnMzesayGcnC5Y
X2lts5lcko7uw2O4Bh3GUskp+xKzDNcSGQcDvqvHkkUMu7s3bZLnhPs6LyySyXKWEf7id2+BxxC+
/cZgieIW1/1yUDZsaDxS4a8LJ8zMjkBM9drtqTnKf68F8YDynO5gAlizfDFN6TD5i7Me1nM8E8/q
wpMFaYscMr0wzCC6DKmJUnwv1yZVWHjf3wRrj8uGpLRh+DoFSp73uz6iTRL9VFnazqy6ag3lRiWL
Rtw8Z1Y33Bph7HN/QYYSV8+vuRxxcuY2N8xFGUYkw8Fu315LSkcHQ7Jnari6hsle2Ufbab+D3EC5
FxlYly9+PEfbZtUPuzs1nJpO+9UxJjFUlPnjkVgTS8H97TXsqlsWpgeVlRDUB1dFFVkxFBh9paMZ
URZDGav07dw9kgSkmxfEWlV26ll/OyBfnWn+tkNQX3toiieFSCleL+zHjuMkZdXvgL4wvPro3YG7
Zsh+iiTInTr5txfw4SlMKxL4UmsbwvzwmYRPfDcxovYD7lcj4XxSTlTVsWBWy1i0D5XsdbP5qZSF
MMeNgZDUFoqTlhxXtVFK8OA2qL+O9L/mKZI6FKUwk7pgz3rqpwcr3eDaZTYnk6JgZfCpAd6gBSlQ
xFRRHtVM1np4rjXBKz210j9EgxRgVH+Xktqef/gtnSoGqYN+GcFlDA4w1G/ZB4xdF0K4iWcOFAqg
OvJEtti6UAdumQJKd4y5iAF0Q8s8eNEMIcCRPGa7EFkINPgsoon8Dj+UARTTYbmBiol1FoV581W6
/NiY8KMoOf50GmG+cngxO307myu3sJyJq6v/95Yj9y3wBnCFKQPJp9pNk8GOwk9w2RY90PesM0Yt
R7roY53bMudTpGvMYvuqBrzyDqtqwn2WK3y9gJAlGU2x3xwmBoOTnbudmfV4kAfYvMoz9jQ590+d
CUiWhtbSLa2VczdQDFzY6YY1R5Tt0mJftuShC4hEo58Gnfjd3qmnDIfQuWnJa6dOxYu+wJG2jecs
BG9f7gfxJv8GNg+iYTap9aCZPw7v1QRNfsXvdqhjqjmPUwlcV/+WqOT09kQH7EhAhoKrCIeoU1gE
h71FiuYoTm0f+RrSzbh6KEvkmb+CHBqPZa8xgpumk/jEh9U53QJ8Byb1bjYPiV/nRKdM+k53vsdg
3oZ1Nmx2Vi+onMRwpwm+iwH226zyc7UGbpAtIqbZ+VJJOLguoo9TAwNM1VWRRldA29OfyLFdYT7z
K8LGgJMUbgi6wF/eFRX3lXEIhOKOhtJIQkaQoaMpLWK7j1PjpwGnQD87fWH2H2IbmtcmSRow2MMq
riG+VfWTQJdtk1b3TT9ryU+28CTzbdxwkWrhKS9RB1WV5Zf6Xu187RbXJVxyOp2qQciO6xggfPax
EyuObx+vrkbLLM2cKNIRAqGGrBjpmsvQij5SIJfNzdYFW3WOCTXj6Dc7puS9/kDFgkeWyhnTHEgQ
EEJwCYhcXpUALhsuKvLfYXktKGj9/oxUQWq5Q2TSdPAVC3x+2PRYZacuJovUso39j+MzUBXuDeem
YOTGdASeUSpIAUHg1tuIaoz8fr89ccIYQLvRuVlAdZb1JiGhOXGyfAM2XlLSPKr6MqJMWgAdfN8g
FMCA60hoaw5o/GwdFGjJbc4A37tvESlpPC3kvnsWYizRsCbqg4WBOwCFBrb2ypSbdrxwh9xV87xG
4l81Xjpakjx0qY2PUj5CbIh3H6SlF27N5iL9IGFNV4P/Rrlp40qg2bwfRZxlFHXmwlTLJ076WGRo
yqKeed+p80ZEEaNI/zec3ItjgJ9+MQTraE94lRDcdvsnLHAJi0yVD5/xpDyAWZhk+n9dCV2WG8eO
RGIGXYCqTjPaSQPKTIBqocHMZlkL/Rp2LTyH/OJIrHHonlHuaxCqejZe2FV0KGFDXvrhBQT3nKvV
khEspN2WDZM3DuYHBWQT1GLMVB63C+lnmTirka3o8QHjW4JDXwqiFjsOsQVpQeKY8pO/y9j5+VV8
qWFYiRSAd8lvhMDO7Uieu3ALWnZvnQya25Zz16u1Mbbc6zlCfJQq16hQY4ilO4bA4JkipEER67kL
2JX7rbFnv9w5mSXFfvgfT0JOG5dYJHYuM3OBfei/yDERmspooMDFlmONfeWfFweUyRs+xpHeieEE
TvYqsLjq82M3ZurCuxduArZIlKV2kkPfHEZHsntEY2qITJEk6ZvdhKh34WurXAn2M5ZH4gFYd6tL
IdWnQJuhkxIg/n6jQzGjlqsLddGEE4s7ULrmaRijNMH1UQTYZ6GTM4noJaRcqihI96RUm4tntvp/
EWpW6rD2vNAXUlLoNufbyBL60wNEqBiAXVOxQ5wwVe4mfp8xJUu7RswQ9qVHE4j9vHF6qeUcGo9t
Dj1gKC1PFYkIwdFI0JhaJpEoxYaFBnu1ZVSUxsnHHTTAAyd3iiOAw7FCWRtWqhDc/wmkZ1894qmv
/IDzE+nGSHUu1W3qj6kwaxYDfGGiHSoS71g9oQSEqJDIXVNvsRBw4zqlKHMHa5RFW2CpK+rcaTpy
1Tkg0IZO60z68wQSOW3co8kA8ay01uGsgSHu5mZmkh+ww1hqnjiXIswcGYR01OSRJ86WrIzAagGk
0rqVd4IgjrxJNGcGuKVN/OwCb8iarkmSVwMrzFaamCheLvAzOTayk5+bnB7VGcoHivlVa5G32z8y
3c6k65qwLIQuLAI+lNvfqK2Mtt8G0VOT3fZY+0Z3xidcQwhBrdTH4DHU8lcpQ2O5IoLgqm8+Eh+/
14cv5zCqjEomZatkuDBuzjTlZT9rJkYVb5faf5Obb8IeRBLqM1hcE6bbaspFiS7NfwcxKkw6QI/h
ccdS5a1y22sHkF589ujA2Spn4Htir15ThV79w3pSwhJWfSqit4F0YOKbrpEWi4h2AoDNGWVZkrvB
tT+J+7rZL9o3JgegrDC21bHStlzPjPC8pa7vA34kEhAcWy9vuOZ5YlTXwYLAUiKF8COKKWVuOl+8
7pViFbEGnOb8aDrswl6AhZXkL1zvKK+wPbVUum7hIYIzuEaGbbYhucJoQ0EbcOk3OFiBQA42Cx1Y
AZkZEQKJ2Sc9+uNTKxkQtBFDbD0pR9XpkgvpFCQHYmqDRKsO7hBCx6Jpmawj/1cw9Lc7GZhGybmP
VPYr/9hIls42pd+j2te8kWDiCtCWEvAeDHc3mfSU6kl++rT8XDVuL5FaJWF8y/XQQ9B7vF5jgcy5
roCVb0GJlD9sQs9CtkDJgwcpoBHL/EiGOkxNuzeT9kNm1xINI2xca+CxoIfkTC25mMCR5ay1uR4R
gONFm0BG4MDauEFUebRlqhK+rq4D4tI3WhjxGtnBc6yDT9FDPGUFazfqiG3Ux3XbabiZ4cIyHFfu
OmzLlA16B9XerGgBt9RsyYWP+R9lHlM7A2fK5Axoio/BAVLuHUaydhyY/QOoIEQJQJyJvWlZJ4rG
u2kde51ONYIaqlSZ/gTbOFeSgCFi7V25hX/6lK72HaQEfukL48sv9NT9OiuJL4F6yosDOrdmfcWp
V43Lsx4zUj/JJgohJZjF39jyTvkNsPtbKxPXCHz9ONcyoYd9figMY4VgMpdtjc1BbpETW5DyBQJq
Tce7+GlzQ3H9INhZDa9d0QVvCANEAyNVhkofOZs6xMe4IngK0pW8PiG43BZCraxlSD0tWW8tK2pQ
n8DR8zXowZq3gz5KY9O4/AZdFnAg5noiHvlCGKTu1A4vhnaFVIcKmxCZzwDYDEMSUezMlxTXlEyx
iEl6re54mmyCC4d+wsiXUyH5OdOmo1VW2Rd+OAoPsDOdW7/jWe0Z8C1f5zOW6w3pOoxYeQ51EprS
LljWEvjp5WUpjJnwmcTGFvRRJz8PV5nkoQXD/+zlf5aDv0AfOR4cbF4B+Lzz7dKVaIpKs8iG4LZc
uCQDqqQ9xiNcR89YiqkKG76YciLAqax6yXpxpVqiWi9bHmAERlFZxK60nn8alleNreX90ry/Cema
bwqqSvVp9toip3l/FhMMRAZfMh9znC/wKvZbA6Y1vNUyKQCJhZEJcEq1DLymZ9lODMbGq5kd7r34
qFdwo/pLqddoZwRXkWGceScj7VVYGaamFQXOFc/rk9uvWsOFbYM1bHHKWNbtWNL2k5vEfKpij9MW
QkGtk7pO3kzkZoa4VdehkznuUAzujyva2Ej37MrXKmIKabuUMR8+UunMshhwy4UFXHE7sDF+Hi1s
LM2ildjCgc094fIVGGqbCpPOeLoqVHpHh7fXGhmZ7Rb3vIgfecVh5B1g2B+Q21ZbDPoHpQTD/Ts7
tr9QzTCALGdVJoBN6+vYWyCLtRSRrGFosGV4olaaX5uyIjTe8N5t4oKblllrxzNRa9xAa5un2mVi
Gf6TbujlX7xnao1GhpYYelnobrcQzKtOSCPIJWhlMmmVThUhyEiTIitIl7ZQbg2/JkwswEVF6nKL
CA2jJMuTbr2CpfUsqsjdQ3ciq4CSa1ULhDDsFpcoPtQ7sLGneh9M2P0Lobc0r6h08mfOO7R9ZJxs
XxaKMAQQwCyaGRRiaXOGiQk9wbKRr7HCODWlMKXCGRP99Zy0BMZqmj7Zg6CCg8MMlxvcacqOyU38
xR8ot+4t9tzXjW5PyWwM8VXS1GfBL0lXaDnuULtsu/poQo1TDs5VLk75U9xENvzYLVT5DaHudaKp
f5B4WH8wteIl/WaSbF9bk+11lf9atrFTei0f3lFQauyLNoLmpNqumTC0LReWsNPvLJNBWcPw8tgl
RMOqWsPayTWy9dZRpRHIiAD2tbCUuBWf6Fg1QC9VTNDqwOdwlNRxCcfyZvGoPzpbBtG3cuaohSHW
x0kdyfh4uQAFzUJtqdJ1Kvbc14Wq2j173vhd2XOCTXsm85+gaO2el96p/9hEdJDjhmqjEkplR45g
ybxUTUDOuJ8LSCAtmgR+V+YOzoY6gy9GKbX2CdoKbdYwHNZZQX2ZaP97MC/uazeK7GGLD/qYi1gR
uMPx+a9XnapQRRqugji8BDt9B2f0vFHl+2clqcNOaG/ts+nVjlmQq1MUki61j+t1ZXWPsr9nx1vY
URu2vbM91B1V1ab2LD3XcDb9DkcWQmQjKwO7gb3aId29Znj7b0RO6Z91qThWNjHwFntFcopn/TqF
qz6N2YL8ybL1mYWo6MO3YBLeKFVyIrLs7dFXcVKa4MMuUB5weXlSvqst71XO2Bym2hkyo8F0QCbq
Fwsd7r3pHumMxk97TxqsqQpKJ9GIlcODoz8tj8bwarb7+fG/rcXA9N4R5bQXmslQ2AFTYF/8jOIQ
I/e3DNnPhJUrWUpwerXymlqrZIWfqXHQfkVRLkYUWS7JNYHHOb4jk0NgKak9t00494lPYthHqAyL
+dBCqJkSnx6AE7kDRwoeX9YMkHt0fTJV1/wfEIjvpvFUe6ZWvt3AtFcR4TbuXyP5+PaYXzjv5vFW
D3J8tom309H/+PXIKLCHI/iMw5VoBPRFFkTa8hOnKFbaxO0NmRddInR47FJw/lVOcAoQaL31sQVB
yK0cwdcAL6zgsuEY9sTytwMbdaH56U4hzfC6AP4kFmxzGdAgrMh2bcecg3B3hdCdkyIS47LR7P4W
cGa2+lJXQBEuSxkkwOSQ90Q91ezriAFZncYoz6wqXtC57Q8E1sQr7KmOpszPqa8mr4D9eltkR4Ql
fHE+MUjMEXK+6XmKDCVTYZComIfVVPhEDnphCG8l58e8eEOkUeV96y5bSd1B4NQ0ZiDQQNL8Cgv3
B8U9xgFgz0gx1lQG7W44XRi9vQG20UlOamNthRQOI7B7DlKXEqpqh/lOIPbAGmUe0Q1iEtpxGr49
Cn/5zM/gbLK2Yg0xO77nyNuEIDQQPdTevDGAQgBK6CHeegokUO7rjX2BLBiIRi3vjQwYp+70Hubo
fl2xrqaWzovimL8FAiR2SWP+yzup+8GL+fO2Chti7W2Ga34Mmk9dT1zWYpZ96wM2+6bb2C70TdL0
LKcLRUdLxlH6WqCdgFInF1ApWNT6UCjzMXYfNYA3g6P5E09wAv3dHUk/0VkDSN9+t5u8PCps+jPs
eS/JBy4Lgft8zztT2lesaPHAmZQXUCSSHgHsYCGZk6naRq1lQOt6t/Y1LlAEJRicG2UkdWWyUuWV
690JZ6bnyj48JM6oXiHlWRg8tsbQOQb080ox3NXcg8y090i83bLzCebmb86znCcgvqbF9FlpPY2w
IuddMTroZg/T51V+bpGCt30tQGuVZk6G2ZsK0Aa9/FfARPqYVBo94RHRKrdwRjmJiLBndE+hXsNl
E8oQ/5HUp5rAwulzh5FbiBW4KQf95emYl10kPK4ve36OqA+M3sq4Bbnz1bnvm2ExJ1VFqC8c+WEu
7ZMnLeXtOY2hW9jWSNe/89S8u2GFOuD/3YPVpcySgV2iZkpu1nYdMpnBIIUUSsnY1YAKJ+YtXpwY
1W8vQqmPq/Hq60ZKDgYAwdt8Ctx2aJqxkP+3gSTAwdfV8wzCjMYTsEiI177Xnsvrq51APVM09snJ
7xH/+jmrNfkYZPfGLLB2CV3tx2wYWltEWjDxIyzSbRnqPsHs+LEn2fxmlg/+lnNx45iDDiUhd4LA
tYtHXxLi49pPOq9jpM7jBGN6IG5W9cB5dZvyvVf8I1Ywdxko+KB2LiIZpRowkn0bXGH8l8vTc+zr
1hdB9OeGcrwdYIEuTnWB/e6YsOx+6qziYzwg4htuf94WD487b9M8JT6jfenUwdOkpS8h/1BBrmLd
1CdrM+i4vE0U5XFWd8kyaQfcYsNghWleydNwIUAe4gskGH1KmCrzAmN3Xdtymqg+3o+w9rz2QLsC
PKvc3NMrv1iaM48WmAmeHrfG1YYpkCZy9MTun2C2b0UXWKNtuH2/cLjZ3Q/pd2/JNYtCxlnBXSaV
obxnHBcDJ09KjxkRXw7NxyOh9fDlzux+kJaQGMVp2fRbPOJYhKIV4lQUc7SgqPK3+og/l914S97W
9LhQORIughBv6EJa4/qxqnYJz+xB5AS0oBOaXm9bTzd35GX4MqBOc3tb3/uV139ieoN7b8taPYLj
JShvTKjBnOE79mEBc80UgvLj280k1IX+2BlQ8uVUy0zHUrrqQZx/enXoAVeKneOhsBbKNEt6fXLz
ByOKNcoq0JVxFS7K60O9M8GPQzf5VBwUd6lb29/FbLk7mph+kEI+xFNdRPW4Te7WORAfY1Vj6m/l
LQ/D2IPne6WksSGtOHGP0i0/BTUoQZ9qxnQE6DTJNXyqPcRzY7k5CwyuHxWaCScr0wHGklUOM6kV
KAqlxkAHuturIPXh/EwntH6wmyK6pyoLEbekcK3kG/RPCxcJqGMM9Y0O+hk0oHby2C5B7a+Hz0SR
0rupeVvj9hH2qLy94Kg5tQx+Xp8fPbeg99G4pCsrDyifuL718jjVHUEA3ibKHhzhclpyKTHBWwpp
L+hdlXVFMq4VoFtoI0OXxJfUz838wjK70ntaIdPkPfuYQzCiH/jFZKdLaMom32bjPwuFvtzVnAfY
7zPps1PJSNlxYLQRVMu+qf51gD/8cGG0NnQcI9MLLzH5EvsjQi5FqhRzvmcVDWebQ/9RizFms2uG
ucn5KK/AYxqQHk3yp8XK7wP8CAo3JFKacwWIB1N3roKdnEXuyPXGF+j65D1pubvbDyGhFhzZBfpq
PClGBxGI0UtVgIpV10COe1TALKgObewVGX8zqjWxhS1ywijyMzUDTAufQS3kQ9qOtC/3hs/dosMa
XEDXrAOz5O7YdhW/NcOu2VLqyuV4KSWccs3PAPJppJ5/KlvRICdwA8pk/FsAUBgupL/nG1Ohmy0N
9SehBuh8ou/coRDX03425I/trKz/xQk5Tc7lAzo0BbxroCKt8OgVEXQnNUYo/vFqXXRIg5+8C6eV
M2UuIVEBrg1qejv6UBVxk6Aa9wWH5oxT4VdrT1zNLlqUZYxjrKu9cvnrVLBkQFqbIR2+T6ncmO2H
9EeXYq7PmHM6y6XYtA2OTdyaRRe10p5waFvbcRbQxZAO0K9AMOqUAPqSVNl5F5kC8UKNeRK4OdJ3
n2jwYr7PzzXa9V/rlPAocF7VyNjZYq0exrCaOfOq9+41bGbakmXurEShRucnbfl2doyIVP8jgDEX
rpC1MZvUzex2ef4YFEZeLcq7yX8r8lQxsd0S/8btNDoNd2kyDGtZ/jyPtgeAisH2mejqli80O29R
vSmrOUjKic4njYIydPQYJTUnM1DCjZMeewbkpBCveRJ7pvES/V0RAtJ31BLoYMUBVZbNpSMLSCJZ
jHgNChFDRuiGuq46QfI2HQbndvOJueOY2VOLEIjvVPfLCfWQEpPomXJ7485Db6yPJOJrcyH6pW3m
Tz6BeyYekZFc/+MJKU4WJny4BB7xSx+RIAKKKdSO74kCGpwGSE6S2ACH5FdAWFFwcSkBcZlKENlv
OgEFKHH2lVH/T8q6IgFS28KF4866huRFMmQ0OSPmDDjTmb6CymSu6pMwueY76FdL4hPu4N0jwQur
lNhxLvlJmLmyp8qUqviAI7bs+wNZEIlrLqa16XTNztcV0p0kgcQhczdHH2ukNNdkNb+cYqrdv42g
UI/RYeBqAp9MkhNGmYumR6aTTTJKLEfoMF7Wtn7z3zWFWZbgBoCNC1MLnAfS98998ii+S/CfjSGT
9gzi7typoOnAMac1g+c3bUrVmU7eXCrT+6WeUttmox7g8DKqj8j35iy+8Uvkqqmp93I4cs4QTGda
CDzK6rXWVe22hq9FbV9RLHVEKtljowD2mWED6evg3iVst35lp9wzGpQQq/aNYzmiHsetSPuVFL2a
Jq1YWSgTIV6TNWzDq56ckhY3NSXGqX7kXjlt0PcqQzuEmX0FQ4usgtBye5y24y7SoAuacJlYa2aw
uku5JqAuMPD+w1BCx9xcDL+s3G/huR2epoII3havgHYqlUTUyJwvw4XRfv0wRvQl1MRc3qLtKH1e
in+7con99e1L+RRDUqlEg41pOcSNPeUoP/e7tkhW9P+TBNyUmpZODttT5z/j5Fc+Lbaayqp5rldh
6w3dU2ifRKX3MyEblZwbC25Zst2WnCHKaRdXTUwkWL1E+OIXGyhP1fSRcTBoyUfWoFY/MHXNj3p1
Vi4jePB3L7fKI9rOUS4+NBqKqww0H7IyHXe5H2PFVHyhDot3APDZk3EfLTHdxUc62TO22/AOrWHQ
FaqT6f2QYd1mWaYWYpmouAhEmGsfh+Q5RspkcTqTqAAi6GAtvds+UjEG1CwJOYvqAikNNZ5vnl9e
D/6R3dV3vvqZprpudBNDKjQirXFpHQQmDcyL1bkQfVjVUEMFSlB/wXmxtx/txVfN2m4XZKRnFR3H
7u/7LBbCD2Cfok0Yx3xhVQRkkvIH4wvTIhKldp5bDhCV+h+TQ4NnjafXIjGUtt+t4AoWWM2qlZt/
26CQWGn3qAnEMpf6i/l6uOAyMAMAozFzfnUhPHmdPS8KqUrUZKm7bb2QfMay5fLF0QRqqXAyX+jK
1kMwen8b+t4dDWHT9UjINCwnSci2qN2csDKf2msQYp0oOEjWYxe7ExZCyuM5m0vN4rB3jaRj978B
k2dRQVPRykzBXVzWj9mfLOUCF6PGLHPfX0KAc3PtN1p51z/9CIbm6M+O64Z+9ksiTURsgSk7iDEZ
jNuwffgYcRwg746LFJ4cPaF75Cc8/aA2Vo91efs+1N347oViwCLUjiES6FGPHX3siiPYc77rrGij
iuUrFrXR8uLF6+pqhsxBPK9KjjaCoetpAcjtqrYyP7wOZMhYmeWP3lvYmZr/AhgE4dn9IXev1oEX
YEP44YUpJ1zVDsep+oA/Aetc7sHLILJh8JY6MJDBrJu4d843HDyq+CQ5CmPCHAKxCNnMYQ40JpY3
vU/p2h8U+nZUOC/r3DsVhOeN7PJBk90s/xXD48v1sVoiUTLEOiBfFcayu3q7q4R3xn3A9A0P1PGl
zMTY72toTDJOL1BrSx/zy/je92PthYxQGJf1QBENbeY0hlFEFnuKjTaEF7HBg1NmfZ2jP6l563N1
FXblZgPNE337WkQ0MhU8tV+QGi7QzqJ5MufykYqZn5XCXPr0+IK3iL8SIYHhD1C3GI5zX1jPRrob
jKUkj1xl0TS3Bm8Zpkm4fOubHjq6cnOQ/9ybtvb9Ah9ESVDEoUicbMZUvEL04jNuc8AbYTcoJHRa
X7ii2ADkZ+GQAykT/EUO6EfZsG7dWIX+j+VYl7XmVQYmmlV1YiJ1XWsmRU1NnrNy8Ex79q4dwd/m
xY4ST2urx0MwobK5Oy/KDZHLwD+FarfaySW9yqQY5jbW1VCHoobL0eX+iReCJDSH/0pgL8NgB/tq
476Zug6318dL8q+kyuuEqAY9HQnJb2Zf4/9oO37Vt1Q67ky0AnIKZIIFJEVxEgmCoBLKI6S4cVe1
c3DMwVBCpC0m8KfWQbYr9cRDlatlynxKmbsfUs58aLsnqtKT7FgBoJfxD2Y2mZCPG+cy55Ft3vT5
JC996sPt+IUujhukaPKTz5Z62Np5MZEBAXLHIvGRNahH7MZyoKcOgQnAq5rVGQh0EIwnUgjlvBRS
tyJPtzLvJDSKsFA0SjGYkyJlJ6vKqPzFnMaBewAJQKohT6lQA1EFiPIEASP1Sp7PcXrGeWZRElYn
ha/NeiKoFodr0TZF0eGqmKomN2S+s+mmYkOlmtYE5TCPzbhQDSrun1pv+wUEQH64w2gKxSxAN5EP
FEOEWCJtprIAxLngDdrsHGFvZSFeBud0+i0zBS7cxIZs8isaALteiTtcql//Scd2VZxiNQeHp+04
RY+HMSuNbYELvIh3mixYZ0sqRYIlOlXkFNWO1nXKgTiNOywbuCLXsgSkCySh67yX0O3zsK1yEwsb
UNIInRP3gT7sI33lyehtttrjGMQjOmbkHA8zLjMApMcj10koi5TI/mGJJnYFZa9b7TOIGj38MhMG
T3lhyohwmBxV775Psdnkxzp69slbEgD4f9BdWGSC3kTPsO8vei2hM1b6YkzI0Y2jVujejCx4KRAV
ngMPfYhEFIqDbKRN2ItQrIA3XtL1F9pOQFNHiF2n4ewA8BpySJbLT/mNNHJdE58BZ51G3bHr8K+Y
IqzYnD0Zpz401AtNK2lJh7YzjF65A/pJTexoqYFQ+XKxXebNVCBwIyJ43HgDIyj2BmOquFpjXqR+
VAKkUeAnCwbaQfdBmxGA2aaRDphnrYv52K7r/ZDg8NF0GpOSIsfMCdYnIu959NG2EEYO/AiMk9zN
HCiylB9943yfKfs03OeQOQ0nd1ZpNkhJAtxLOB/2aQnh2IuyHlMqvGfogqOi0RZPIo2Wus7SWlzV
UvYSONgq/ZRBMimovt0jK0xdqAtPvNee11BukPmoEL+hm8ie3m8z3ia38+2740Ubo/2F6dd2Rf40
Ws9Ut3etFtzAQ8cNqMzfRvwCYNPInQiWS1+1vFNjrnQiFt9gpRp4srVlQ4Tskwgl1Yrz2irPH2Dx
7T6lrr8iMGBSwHr9NO+xBQKMeF8DxSxlncB7ESLCgDCMymtDOXmdRL9tKKl5pojn7SohLi4cdbzn
mAOz9N5OeehBIcB768XWz54CPIwOxA45pj+V5Xc6C2nVmgmWdgTlEvk4r4dwrxXAN+pW2YNqrVp0
/aV00rtSS7nURAedyclpjOkSSIPQvFlkqJo3YQaMJHLpuLH8y38ekYz0t9owswiq93++rkbMxcan
gJpo6VCrUkRYKg6blPdxBZW+WGP9+Gohn3v/xD783ARqUbusK+izAQePrm1Xlkl+5pMkMdh3VVU7
5Yhtjh6m9TZPdp5Xtph782FYXIEXM0syZQuzSyqD3vaCmlWBlMbNCD+v8+NsBBhC0rGpnUV5B+7A
4+tESfHeAV7kPRDBjkQJB5/sJxAq1mp6EE2BwKAiJtIzI7MA17LsXWzfytZmLRGpQzk5h02sFnUo
FKSBJMy+uRa89t6vpRd8rORhlTEMLQ6Smaix1FOqpNK+bz5XnWuswIfVYwGfJPsvkPkuq04UiWAK
7rvSlsIvXm4Tk2QnyBBiitIoZKIgBkeU/tJMfTd0JEBashQNRvZyvUs5OYDxJkHZwm42vGOFHFAO
pBCKSHRiKy12YSvJAOeqp8jbK1rMRpqZOEkV5hWFDQDV61bkPHdsEIJ1Z3562PIZZS26kxkazHq2
ibqZVfzelQcPC6u4MCZ50DBamv+dxutL3yofzmUbEb6KJzcEg5wX8gpemsAHgbAV337OZoXhJFgh
K6cfdlPqv9Db0Zq2XW5KoOZqbQvNd8ZmT+1LvVoT/rAbDmVhwBCQh12+1sGw/3MTOdGUUaGOO3Bh
ZE3zyVw9ecU1C/obI4irFXAfP4uAwjUjusxIKyY0SVdZnZqWeklrwFcpu5VMi7bu47L6mqMwH0h1
bR7ysv8ZTqWIkn9BfgImI92KbSEWruSK9aPfQjEsjrkubWbAMvZ4Vs01nN26kjjCE8PAXi3Anftg
EiQdjXKZRb7KvchdQu3qKjmueIxKl0jKZZ5dGFs3yeVoWeLcUZv9Yg7/SHx6g7MV/DN+mndDuLi9
buem4TivnLDaYMTWDM6liC6MLWZ/QPMD/QXYHKRx9pv0rW1krsnz8D6QW/TAbh2iwyq2+bjrMFUj
N63/qfWhl5EZnaYZWUjZCxkJBYmSAgj/WV5whpI2/hn2NLk9tgVsWYAW6EvfDVmONf0xfX14KdY5
C7kpEfElAmLlfM+J6527Rt4Ti5hIrPVmYd7YhUvxkM6xzD+0xBJAWEImxwoYJ1+Mnr4fqgtcqXU2
lUpTh0raYCvWNktur+YNlg1gQP7WlrtkFM89jp7esJu/6SYY3ec5VQ6Q/B/6/EHnmRQnIChi7eln
TnVabbgAghTTMmZiA4UIL/xLtwenlM0Fs3cM9MZqf5EPyH00GQkw+GRMXGlmiGhBDua4atKrb6qL
otM33/JTj7O1WvJ0ikgqCBln3DCbi5SJL6cGiupLmetdPNjuInntQdckk8PpRWh+1IxJbMB6oo8z
4iZ2V7AQHCtfyHOF2D17QH/erjq9QlAoa8gCdxGwtjUd4dtNLTsO/z8JuO3WBdQxLQERxPtma4b3
ASQZa9sBFYnrtFRx0Y5Z0tjxkf2IXdNa8bCRd3dnHm3iw1azycp6A1t0B9+XvaWspB0yv/++9ibJ
ehlw7wBLHPKkuFQrk+rKh+qhExIgiM6SmQiW41rDDpVcIFs3GWjlnfbHp6IeteVsMatkVMGITkwe
knrr64tJoV7Mn5UsOZDuFCuXekgaPwddkEKvUC+Ft0FHLvViZ/3f7VC2JqXwPSYJmFqP7+ArDCel
i2V51IGRt4QxzrcY97BYcuZSB5+lZh4+mBAZvJjm8bR3QbAXL+bKAEZBEk7iD14LjO/akCwo+B8v
DP5p1ovC/oMghW3EuOdKWWDlfy2U7rsiBlt/dJe+e/EIFdnvafQg2mRhCrprXcQzGto0fvwldJRB
Cxwkr50pTRwmlDRVh/nXDd5DMGN6HhHX3K4OoT5vADUlZEDkIIObOFau2QCZiUGenEXRWnl1V+Ej
ASb2EFO9vNcFWb9aPJcmpny0f+Lt4Ad2/gHOH64Wm2SRKnjw6Sgyfl7TW5H1nQgsWRvhiU4j2sH7
NXc8yewhM2jgQJkfhERKw4W/IWdk2zqzvkepGDd3hufMPwDROOylA2u5y3RckHTK+VG8fScHd1h6
6APm7YyWJhWjPfAfFNnX0VCWwWvQpvhM7mCm+xzsSj2Aopdrw5T3vhV4HH72F3veen+m7xVFK0mn
h0/uXYB70DlmqKwRdY+WbiUxTsrs75mxC57eLWSD+8sjMjvEI8mSvrOkp2Kihkcw6KG5hRcXPtbH
S60bndsZFrAiReWUygCSFyVe1I+YTlxcUBjz0x/MkQM+rASNgMUQzyJT7OhAnWbcntMcTCSLYUGA
g3KR5GGHkWXt1n1ZwSqjdUF4CmGPAzq+XxxOTNpxEDacu3Xl0IWgBEDTodlImsJWsOFX7BeIU6ST
BzxPwZSZhLTnvBumKoGjhQ7TBGJ9ahl4f9nDA+a2ay1+8RGND8XL2zoBN0JSK9qKcC62s8oVUXVZ
q9FXJQS2Blm7n7tzMYb7rRRTXYkmeDaLkLvy8ZjiScVtf4umQrMvixrFlePsO5T5cMquEQs5CX+b
pBWuZFTSly5zKX/DiiaLnUtvBZBbvzl6Etm34PU6ePWuMq24/6+iQsP75ppAhUHILzzhTX7axjWd
m0TbgB/gJAoN7LvTYg+6yUXYkXbl5RT5gO8m6MHTQU2VmnPcuUQxa6+aFdKEIQBDAOf0H65Xxdqo
SI4t+RcS6/TKlrx6xgIxdeF2al4O+8TB7Grsh6U3o7Hje2BEfhOAESqXkmlxsOcAjULljo+WiA4k
RC4a2LB6AIFrN2/CnfywPtjGUHWkVIvTI7EMpwtTGyhOI5mf4VSPBmR1yF9cvRCzOHx4GfGnchFo
Z0UbosSOOYdo/PIpcAZzbc0J2k1bYag3aeWTdvDavsO+x4vI+3OXNFzjwdLCkzWikCGT5T/f/0ai
anXHhYQPVmOaKmM6f7tB7KsPBtbotE4EbeG2nhNe5grOPhPY01jPpWb8BAaRJ2x+FXSGWhs1uSez
TC3PoUfwhcQ3Iq5BOXxNOaPqou4fOKcFd08SEZ5GG4XdkMFHLqz34L8tb5TbTTPIT5iaihFvJHdm
y8+U30SnwrBnSUxAnYAfRGab+i5O0YTjj5+ykRK+OUrZkwoBWsJKYTu6i6UxeUvAhCsMl6/fkg1q
lXoKcpYLnoq4Dl93etTV0k7z6OUYOraWOXIoqmGbdnM/NtQL///j4qd7FBVTrb+B+gglXKnOEbbx
w0RAJm7imF1sljUuT0euPYF3Ne1+lWb0teccmxBXWHpqGBl0VI3G5a38Op5lto/mhowEuiY2i9y9
/Gjjz7wLwAEXR4iv8R3X5p9bId93aJG+NAGVjIrdUycjC19ZkEIV+l8BRav7fKbGWLVwC2RdiPmm
v95mvaI41/zMaLSwY94NQLfc4oHtfm5BQeWlj2gYU/lCsQfPtQ+gkrJWqAbkHlFxmCArhRAJbmie
qIMZaAlqn0r4Xz8LCuXMQUK3JYW6BpIqzDC22ilmeT4pKOi9fdlB4XlF5IJb4Jnlz1mSv7LEwJfU
ib7XcxK3hBy24BoIhgMa96ghTCQJ7fjwRyZerikBpQyYmRbEsyj3lmKAc48WZjmg91TAyKuCwX5D
oalExO9exS8+K5BNgTtM9Xs5PJlHV/UqdGeU9pswgspYTyFCXav6wWvsVsqvNozpPYtD2HVrnLKu
jScyNTMkOrwAnqboN9OfcN26nbyw0QOt4ajUmnVUzViBQduknhMOT2GsK/YK0/3m9HejLn5rLb3T
rTsy3gUsczv8JCxcHGUYtSYBonukrdHw7B4OUhMoa+ih+0wJ413XIpGwm+2Yd1ns/tsuTjYAumpc
DqBTlVJcJqMFzJ+HtZzyx0BhNltaxeEGeQhWnK3Xnn9RFDxa06DBYHHQdcmNYpuSLH3UW3hBFtR2
1vGyMA1XZ2FtvZ5sPPGdRaP8VjSfIzCslhiWxRbnVTcuu6LrG47rkD7S+RU3AbKSQZaRljf9UTe6
q/Rvg6kwAyR7A6eNIOWXh2DBOhJGmKpZaN/fq5NHW3Fri76y9Km+5497aWPuEGYxbhSyFDe121Kj
tSivj+rem7pqz/GsAF3Ygc24A3gWvZLr3BKsKVZRTmR88xt9+vvWpjWcwIvEBVbvQoV2FN9Duf60
OvInHIy2NhyrTe05Dk9zbo3ECZDgDl+CLaLO2dNvfZn6L3NJ597fu4Q1Ro0cyUa4gAdTu94b7O2T
l8KOVb/iiPhj6l5fl1yOzz2/2pBRgrBY3zdG+hAekhKnYiROpH87CzIAgbLl3cyHRhXbQspzOD4L
yy32yp0T4SW5/B/cNTzqdzMvBEqqSO8hiLJ8BuaNdAjxqQA3v4tjb5Em6StXng1NlkBMwA9SL4o8
zwdPkbZUXiNP25Akp5cFTWZaoGmxonsxvGPDMjLtjKf1NTY9uq+jK9XbIi3trOlwER94firzsguW
xLKcFNsM5MYtLU8vuevwEJuSvEgkcuBFnJNztcGfpc4CNmNt1FXZigUy9QA81Av+x7pkHszO/r5S
tx54uWQOvd2svwYOcW8lRjymzLZglTFhs+mmzQM+l0tMwsjvios0xs+rkpqXM7tMzndebCdSLMYp
G0VdTI6jO2VHAClZU0qb/UH6M/2i3i+WPrcyCZIHkL6rYp322a7cZSJ1r445vPph6OoalN6n7var
CiJiL6355ONd0xQeECFOULe0RMo+luXTU5E1yH4xm/OptgZREHeTRBXgUFShkdF/QOMZPtoitU/0
iwoAD0itQLGNZAORcB7EvfNPHcf19vDGuajlBPPaB4z8uNq7oTGxcJHQMZDYQ/3dr/6iLnHBzcwH
wrqqw8MygGoa5xS2VvqaL4c6yTZwrNZzZsNoLVjfI1A4m6CaByDmH9yirzfEW2iEqGgEIRd1Csgk
UnP00PixEouVRRNXwKb0igE4yRL5V0jsp5bVLxemIfbRrSJePRFlqoAU5U1Ov0S9BVhcmK3v5mmw
kPc1FwY51AsHOYi1y8RQoTbNKobu3ja07SQV2dED7S0LKPcc6NySpy2KE7CAnvW3u+sl/t1P+/pF
kPb/JI6YijTlflwmr/5vynw6EHbTPKM5oaRlARtpPlt+2bmZJWKDYZbH+Qrhfe7s2DBTU1sBgUe7
OZB1UUXvaEbE0aihHhFY12sNVBl26PvM6mseoQhf9aF3HNp/VxqLs3Wn4xcQyWH0SxYE+DvGe3hY
dVCPYXU1gDeC7oLpoBEwrPR8AkFrtP7WF1HWoq/hkXZET04tGf4W0FXx9Smg+zItFrBACD3hLGMj
Z/e4jriDD7iWaL/XjtxQ/clSpksSQQd5gGezyQ4KayQyrtwX5lhhmW1qxRyYsTcWsrDDfICJkj8w
wOidUVqL17Qcf/qsXZoQh2wJGxKvJm9FRMcBYi1BevNVFOl4zFKeHvIDyRmx+zMTtPC1q2DSxR1p
rFnDHXySHQuDsqBurJJBqQDVZEHDmG4lmUBLTdQQeBFf+A4YPjoBqa5IZK8D+hqzGR2GeHzptqYy
5QtiE8XjtcMpWRcExd+ZUyGAS46prbOHh/codVnLgjW2aK2mcWdAN9VQiEMBlfwEp+ItKBw8OSiO
f2awZvswHFciWLJ3raMv3/Y+wYP1Hav+nuOqX1YOQrfr3+fpTGTqQEvoDMBGUr7WbFzwH9qRh1Im
Ott+0Vjg3Cqm6wV+1wUeArwpzlQS5omNpdYMMbS1hatXWkWAU7lUf4eXos5iZMiHaV8v0B2wPjzm
WiMF+oP5I+gCLCrmq736eZBD33n2mUA1cN0zYf24RAD2x4f0EyWzPTe3deRLqZlo8Rx0HRFFdtHf
IrPGHDDl/fyATcmo5ZdZmQjva528MjHxFX8x3qhLltELvDpQEEREIaJgblJDju/ZOy4+mpuaAt4V
pMKXy10zC5yydLKJASvJHigdUHIE39JloULzGW8kwt0QNirT1mb+dUKkHIACjFJWP8yexdquutYQ
T34sah1Y1YJtbjDKolTejnouBulriqLYlVG/IA+yzCAYpEynVM4vU8kW+O71+w1FYiv2BHflmkFx
cHek8ogcywHDDwuoeoKdDbcnOuWgoES94ZRPBBLa5LtE31CwkZE5YnnGLT6I93xNY89k1Y1HZixG
lwulH3Ec98lsTDTsSl7/P1y5h4WIOL8xCDHmThyIMdYr7FO7boGRgHEz/7IzDnM1O/WCTpwELDa7
w1HqECcUz0oj/9aFkVUqpAXzI46p3Ksm7ovSNebwq0DoFD70xSqrHCZ8kuOF0lMEaEQ5jY0uGdb/
SQDkCt3XP39ND/v2chA3aTPnSHFu4mLzAI21LlWICqbqCBZnsNmmRU/Y5t65H05e8xmP2iff6YuC
ov/72+owJBlbQkPaARco+WonUUJv4+zGCko6DEbk1dV4RoLxBVK3ADNAFM9f649tL+yuV1Kq/l7d
YBdr1buL5VksLZ1bdxCsMmSDeHf4Qse0FlXBZ2OA70HBSf5YHtqeAUzX1V/Z/k7+oZo6u5Q1LwAl
oIHGYYi1ioaRasH7e+RwsbOnWhbLzcjLlkMpHdjVbrK78ezMAEhlyI2TcsvRFzyl6qfA/42NLkr9
VFhLy3plEGWEbqo0+d8LC9+Ixs4ESnYRXFtecZYZBz5QVf3SuglucjowOXH5+tBQmRPSeqjDkbab
/nla6UZ+9tvisVK4gn/29Y51pMQqHscRvnxWy6QA63DpaNx1HvY2D+ctjeFBhupez31fF+9JmG3F
Gpr5+lzct6NEcgvH7/u/zrP7gULrLuQiV9KM68bkJ6tgzaL+Wohyh19GKboApBRm5qulU7U6fMpJ
/P7kztHk+CHDaJyzce9wXAjlyilch5k+pwfkxoypHGfguo49od0Nl+Mbvh9hSFK1Jiu5uKM5xNvr
0UtoCM/+Yf1jUG6YbUjX5GmFVJ20YbIgb9Q1Gimu/GPJTiv+/nhTVymPLuARYB3cAzf/+zASm07F
fymoCZYABrWTd8HqRZhzCXWIueT+S9tCqiZLodvQQyUPoWNP8v/ne7y6ruewPt11V2GjyE+nMhAQ
OdEgoQy5Rj75ENFqOWBkiWNYXpOpGp9oYOLNw7+ohi6u0jkPB/CKaxeqpLCD17esD7n659bsrkbZ
jsBAuF4dB78kZ77o1v3DaVoBOfUjVy3SiVn446WAyZoS3q9XZMiqQCEPpTuloZtM7cLXbwmTjj4T
uxHp0QINGIM0qwcZCLwMk7Y1q1sX3p4HZG74+WNyzv+g7P0Kf3bk0GRqGzDAoPoLmhq7VvXcdk1L
eS7BvxXbhc21iASXEdGRtYAEEonYSPJL+w++Su32X4hd1PGmLUjMl7Mzzx2hQaTfmu1XJmnOxXKZ
YFL879uKcDAe5g69if4lFomJ4d+Tltn17GKg07/iddZyNgYmRndV4cwfHLwknITiGwFIfnYcqOtm
+6gCAbj1qNlp9GDsMzpenfsXTO0gzLKE05cauuCV/zKnyQ8AqEQlVOBlC3j9k295lQbKo6+cdRsf
HgK8xVa+NdEkHZ86/4J9kOwIjYdchThp5YZ69v02echxbfP8/upMxMitmP6qDiNXWAgJvsJIwhlu
f8dASZ+FMMl336j6Io7xf7dbCKv8wn2J05QZ1s0L0LaGTwz9JM+xHlr9EmBBc1NN3IEKqddBQCtt
ceTQ8z0m3ENa4fyzp0huQuUEK5r0l4DM5cSOfjVDbKAs9Y2ncrodHOKqYzlueTkxbeHshMNSB6nQ
cooabjLveZ6K6O/6bwWVtixatNy1Fem9xiMXiCu5CvJBhTYPPby2bs34YXmN58etcfSgcIJRV2bv
aAp/Y8yMdqOGgBAxQ22EjTvNraZemRl5Af0itOaukoX+TbrBDmPVtF1u+6+RHnX4suiFK5YrPf3h
x6e1Pm/J1jXsb+sAxtFUJmZenXXAY+KWT5rP9Grhn8fsdTO6PHr1w4Y1o3KSmaKo5DtTVNS/UdwG
PxeX0rSlS2WI1DyZ7L9tgCWqi3JF29KGPD8jvOK9FqmNl/4sDW+uJZCp28aio2q7XSx72VZt7bSz
+GhoBbmRGMTKAsX0LM5FHkXiWjJX9XDvsUdUqKxlxgitt3TbcBUNtJL6A2a2n5wSVjz4nZcca2gk
JwDerSbusC0rsnpUSD8bkEXKpgenfKrNYmMM7k2E0nqhgquztIPRqOQfm7eWrfe/kJI2Bzw2kKK8
Iip32yNKURxeRB3fvBG5Pk9rPM3RolaUYDKDe4ffAmr7BLEbedRqFqPJdgcKVwDnhGWCXlpHigb4
YUd+LzajrbuWY97GgvbVCIv34y+p6WPgWpBzoPGT/eeIMqiAjll/SAdGcp0yFRYQduSYPkkX+R+3
FJyrQ5rlSaf9jWSDAA7cHjqp7nlWZcIR2bqRL70zyXxYgNEhJCluxND0/6GK6qS/L6FSZGiPMjQM
UdQvP5tubP388LAPo4vvmP6pc0510WAGtDk7J+HAYN5T1qEohBO5zgidtCn6LO+8fMuhTYEaeAkW
HhWc0CJod6Gc0n9tFVHjVSderyFRKjf/JPB6xwxhFnJoyhSl2V8U8Ej+CrKcJK0V7HFFkinSK7uo
cBW7AmlNQZqkTy+YDQXMHVL6RbTasOKvvNK4m0nEpvyp3kw1winyktPlDQs0+XIJwkV+NIBtVrr5
1E6I2xa7Vaw8DWIleAQw2ZzUzsFAQiO8enma5jJ79ccCafXYqINrYnBVIVhTChQCeTSybVP9IDu0
rO5AQ/GN6YKgVsh2JHXF1FtrPQgR9Wckb9R90hICOY8RffyCZYQluaihLbPc+YD8vsgOK7RYiq+o
6heWgACLURz10dq5h3B/d2UcZxGUpUOK+CEsdffDVACQqhbpiLkERSkqZ9+pImGb9aNBs7wbUzHe
nz70HB4R6sqzN/cDnU7jKFFFx8Az/kJg4LaMFkhlsopGabvsJj8T8Tl9IiUgt+J010e3+bXmx0lW
CtN0U+gn7WFDy82Rh4Z2KpgeuDkeBjSQHb0EY6LOsly0/NDtUAbdm53zFzk2t6WeiWbm7jqbrz2O
1rB4F+kJWmpQPLN8aogv9FEF5ZNJTrKm7r0k1EFhoKHiAJs1UWUoWPeVMzLQu0lSG1IRlkIHMMfl
wz0c0c7UVx7P9rgWWhL3p/rx5pM1pQYPMN51ehINwIk4HaAxRVTXSNilTkr4OPlJSpM0OFLbfOcK
giSyT3ql1DQMq5bMyqwb1ke7eU8kfhdJT4rHZPlT766Sp6Q+G0QZYN9esfL03gbn361FxsoNnd/N
PVaTdXRB+LviVpyQxo/uUleALkcPGD8qGtB0X3FKaP5ijKWQNahonI2ninSOk5n4IDITkohKB2MH
yI4GaHNLiIDG/kuXGinMadpZYh9EK8S4UBux8pbAyiwudY4tYNzh4fTrRdKT8ZIvw1GNvfhfsb4L
y082f50g+ziQQUAzG26D8WK7y9Ulohb5GJhXA7EuD7wkWm6WovpqqMLsG8wiLwqE6XIXsMMyyTD+
o6qqANNisGVMwPiTq0xuVsS/J/dLQm3W8IwewTgNRM7UNOrTh3WMWoxlcHJ0RdhYj3gL+X3XM1sD
KpT3dD5tBVrobC+hhT99I5Wca80CX0LJ0/0OKdHx2lr42SMe+n9TR7sviOb5dDrziVk37nBzR+oc
WKCbcBm+jPHRN05yEHS1CgsJ0qcet3e7y1v/TjJZDTagRRSm+Ces3S/zKJ6Gkd1znxsSPAcADmlf
uXhGfrlfKjPi3eUdWbVg9tSfL291pWh6bab3Sn3miYU46wMVwpwO5W+inODBSXc3kdzCpz/+XS37
CRS3Gz0JCadyJgs42HFYPt3k4ngnS4AD1rwQlzsra1rc37ybUWuDOnm2VsMH+GBuWRt1v9VKAlDr
EGks0PszdM/AtdfsuGGwdUhxEIdsCMK1gAW/znqJhSCFEyOrJ9Cee++FztZP2/OMWBwL4gbd7K+d
zbFA4goALSVkgMH8w1NmiruV3p1KhlYmCdfjMpVJS+W9IGG9R74M5+A464UOku2Sg8b/8kxAuqWA
bm8ls8KedUSEAn7nuHQ6Eomv/+q+mxUpwwdvqBKwayMc6qLlwDoY7aS/wFOWrJn0iCo4K9WG44zb
gQJDiLGLaV55VNDtOV8L4bMIDqnHKVSXE02yoFH2J6vy8+Ahu48UXyJeXJOLNZTeeSq14gVpPXQ0
Deq8UBM41ExeRSS8Nwx1p3JfhpHuR3PxtyRqryzv31otHnCiF4I99HwCRf9wjWEbJBAZvxREb6QK
Ne/VgyZmrd53r9hw5J+XrwewQBkK8MxYR5B7Ac+4QYW+f2dBrexPEOpUPRVCNTwSpmempety2gDH
AGSoTTb1HbS8jpb3e6k/L2ox8rjhs1hHEmzmrSqEb78DnSSDZLwZEdMXP8vlEhKk5cwYZmdTGa3o
jxuZ804V1z1b26yPoJaIQOj3VVIm5eIkneTlzVQPFBJ3GpNoQlWnwr3FY4T+lc6709+mxsM1RNih
f+MQ5ag+ElUf9ZY6PNYdrLT/+nhSUIlmZDvnrY/76EpMxPUzsuTRO8iEGPB66bdD9pYlmik77gZy
cQfgfwMZwmpdmerbVbyIBKpM2GC8XzgXLJXc/avmVruQIjoXwiIa/SMqa/vkTkCmlcA07PKrwnm+
eGtPjRa2fCw6222ArYIWs4SAVWhVUMTmRu4aPFFqmxBMrAXsRVz2vZ1brSUbQdV4UIjhDM4F3ahk
0zf0ryvNHw5FY9c6tvns6kjdtJOk47ZmTAlgHLqyJ2Srb1Ib0lbSvx8BxjaEg5jMzDK4XceolUAk
BA461bcLEOykQ5fGC87E+ieNdPjWuyakA024XGdr0gWHFmE2voZasWlRCeHFpjYqSJSNGKK9pf+Z
ZLKcf0/xPS0goHwCEfd28+2/DZLpE7ubi9CWaA3PbZxk6HZYix3xwrot623r0yZxQFrYi1mEx3O4
fxgNVi/AwpOh5lX2mM6PKYxp6Uxqu6C2r6QH29jXvMsUGdr+T4nJamli8kXJt3UfZkblo36SVC2P
Wgd/LVG9kFPempk+xofvnrzh4d3xffdcP7UaqQBjHsCyih/p2wzE0Fah8m5QX7J9low9uIvriKEB
8R59Hha77HzT8VPrM///fCZ9L/EkQlKL3oCIbDPzVuy9gSLAgFo2vcJLtdkFN0nqtcTNn2a0DQSq
eDA8/Ve1vCANpeyh3Hn2gS6k2cpUwmTTk/1HDIlL5TwQcj3N+mx7RQHjSkXzRa1L9jCV9autUJ6i
efs9RVnf6l57Y6czwwd/v1+rNcLSwxxdt1Iz5gEtjJzJiA/q7BJqLv6IyT/NlPZ4d84lmXhkXOJp
/pSfdkwlAX2vPcUJbARY7kvHvq7wcIz1dTIQCwOrDn12Mhbg4lPXIXXSd7D+ciOxeULP5pXKPI2k
UL9lgnBxJ2sE0088I4T/E/SMe75ojeCrEPsx94xhNM8NcYL2xpv9F5HOdCBnV/69jSgHjf84tECh
h/ptNVi35ZKGfjad4HF1iINLnQmQp1AdPE0bwTPbMyFzZEVrrS+xEw0ZJUj2vh49UBIAm+x8Q8KB
sJgOyh+kgI/bfwX/vX6inz2Am9ECk2uJgFK5Oi39lZXDGwL6y+nC8ynDQIxiI1eRO0szc2mpLuLO
IEk4XPbHgyzNPtOzHr2LqbxRzZfWwIWXHdfQCsrDHq0C3Ntamds9GEXv9OjmGcGQfVNzi+fyhxHA
463ToT7JKwkhwC8w3jk15dPZ4L4DaKQRwjllVl2PbFJWjBdnOKJO7W8+UYeGh8vw11fBDrnKXuHi
iSkgJWoiz++eY/XMgWuUyDa/Db1TayLZVEZiv9kAW2L+ks1KxZF72GVEdNeEbVFIYIUeQfpFAibv
Sx7VpbJ4F6D92tBAgC7lctWeyd5zcHfmG5my6yDsc+H6PzwB76+XhPIRLrVq7Mz7UtZ2j3p/Ywlu
B/6cxG1N7D1m+6X2q8v7yWldVUNaDVmLstb4rQ9IfOy6cfOqmq6NZcDAe7MjJOB0RQI8t02boc9F
xp2W3JymOZRh62WXPwtWD07gG/zZk6Tt17CLpNNSXrSUKa0b6QV1XaTraTQy/yZmMh3MnjyURxo7
UsFwQhZXSW4HjpmI0YsIniqGcsAsvEhNZwvceoqz3ocyy0ehYptIA0JrxFKZ4UjBHgRpDSQ5Ikg/
LfJyDBQoCuMN3WeGiymdFNlXutKTmkMx2aWz9Kt0pMNMX7eUL2fS7oJaCk5AMZI2XINq4dXefXUz
rnjigGA6UhiMDwJIgr7W9/V4UyoR4E07RxVIkPq7Wvrwmj8wEXA89AyIFTllI/HrSImtVbsY1ckB
cF6+FphTSY8FItdnrGnACQpD0TBii0QDpsc8sSbg6/mG0AmbB1aDwwVmZL02B7uuZ4UnSpFjCmwf
y5pjIjoksv6ZA+itVJEmQWACcIAYeuxJutoTXVmC7rxpJ1n+BRt82gjZa0g3m/DQkw7P3/ePEmXA
A8hJWskiKQRAcNqrZPPdDp6nrvVNPqKgVyGygSbnJZXvADmpZgHj1cx1tJ2J4LDov9mq3QZHpcqj
89gBNqQDLAfjS4TL+hYgoK3msgdggmG6H19CRMqaz3I6NUwk9wck/QMdFohWq4kClx8dkRvpDiHk
9dYVfauyymwh4LyfTtIUsbAFqXFfjJN5vSTByiAnEdQHz7CFtQhxD4Mlro1ZkN/K+5szUUTvtDId
9xNC+x6FN7TBWA7ZOWhMyYi2UxaJ1MqRkAW4Fs7V0lE3I4F/s3MqCL6XYMJobV+JMK78Gd7uAySG
Jd53dP8+J/xSNSRda4TCIGdj5p357RoZEVwvqcR5nGFrPxa3NkG5rKTjhH7FPan42MEAawMVI19s
42eZzoO2dLOM4wGFoz5ZpBultywnErtJgHWWVj66vduU+a9kWnfIyeOIKVQ4/+1wlchevevPkB1i
uJf8VrpTk3tWpZVe6dC7jNPcT30rrhpHB5KhomPCVC9XOR4GM9fJ198Wtwyn7TwxctSw1lr5THXg
ydmzlXGoWhs2y9ms3zKUWwPcrUqxSUTciuGsYP3onHDUlbpkzkBJIjcZE6ZggruPq7FCfGyfv/Ul
CFV+KWZ1jZrpPnEYoXapId8t4PMj2FM3kFEj+DlAKnsZbHAwJIHRTVwrhyv12GQ3lndBpW3vHdYP
w7SjsJ6KA2Xu4tIBDOMVtnDm1VTgkonSgSrBGnYC8f7CQAbxqd0Fg5QNDgZKjGS2qSEtG87LSS2W
L8CW9mpT74EC3EoF1G4WLN2Icx0zagod6cyGVT7NyEXPGPFO/njTrAeQWd07REabFdgwu9xIXOcN
QeNpDCKmwkmbvJVb0V+ywnEpfjjPfdqS3Kd1Pg1vtxFsDoVtF46j3I6W98kWDI/y4wYtZ9eSoavs
60oGbNadSngVr/Fliu/Ec9l3+2V7LV4QBRjD0ViRgU98iLekn/asPVuCquKO6U5leKGVZUIAKbnv
LTHQ8WoUtzzld85ERyKcJKVk1TjX6ZI0J2lGn3B/9lucRxF2//HYye7wpQYctbAGaw7ZQR8u1WA1
dJFtC6ojC7fnHzvcw4OrNBkUra2/5pRFWhBDuG6p4okkU1LPNE1pb3Ry1U1BXRXoIExdvgHnAn2f
NxT1T+gQqj97d59DvekYfUe4gKkj3GCHn6TV+LUawqjOdyoeUg14zTghz9S5Fp10BcMqVbN7r956
BW89WU2Z2cxc2drLxL3YR5T+BZfLTjPlxBm4FipiP6UyuJv2z2WF4uUMRFnJUG+TFwtBEQi8BDXe
1VwXGjiLjnu0Jo3k05/oWj/umxGaRRI7vkATs1/aTB+bnRDBLxW/lXXvflA0t/U+iDlzC/JD/QjI
0mabnZyI8Rm92Y1vyMr1nQsrQU3PO0t2tK55mvWUnJGdmbYUHPb+Aq+l7cRgZJyLeTcattb7Wdcx
IP5X6Tc8fZ4iGGfgHqdbyxQ8AAmySvMuZuoBLbI2GC4Cu57dpD6IvUXs8gGqL9AooKUlm+Gn6kwR
+SRES9KYl2F7vP5cl4JATeT9m7ORmpekaEBJwoP4/mCifAiBnJn+ncUR31wDHeQESoyz3iN7xxP9
fXbEkYdE4+mHxp299f8Lw8QAQQ9yhdUIeFO4mstMW71DflLhx0Q7iBD9pifBqWFbMT36WWdHtaNZ
hzkpNZzt8ys/wTEoR4Qahj8EXFuGwUjZgElioeEQB//gJ+L5ESYa3W9gHRZ3vmuTiITNpQVFB+Mo
uHRLpoq2tR8uS9DUQEAJMPAIW+3GeE86cWHOLJDJen8BgyYAMv/tAp38b/IeQf5wjrXoKk+MiPuz
BDTjsOkCamviBMwfM8jBGTYMdukaBoTh4ZZsBowcKVwHDQ1+7M6O+xipXmIB5iAp/NwuyEqayf5Y
vW0/vkOtDdg2bU3GKU45gBKBSd3Luz6GjHadHOuIzl6f3ffivy8PnZDiw9gk3QW+WIVY5nncuKUj
HDyiVmOhgnBJuDKDKtE7XrwQNCSOKYbwBh3hb0IYSFNn/f9TShuK2V4ZCURbAqIu13k4NCaNTqKU
9fQqpcvGqkyqmj5gEHVuZ92BEWPEk36iMCrtYl8A6odrZN0S/HXYACG2DgaBbw8beCH0eNHxacZ2
Kj8TgiMwSQ4zf71x/VoBAhIqOTNo3voShm3o7HwISKqaQVc+/Yexd8d6Lc2FzYeG14H3EJcNDMpU
3N3lwbtNI8iTxYG3eMucM/oKpLkT9AbaGaShmIsG/5Goh1G3XPIqQJRz2zjkQpSTqbaE/go+RcJG
0DLw3cMeFlMMfZc4qqpedUAwY9UbE6CfMA6u/apqOfaStie/V41C+hCLA29/pzBXUvxU5XRMYExj
lPwH6FrFakWbWvWRf4SUKRjBE2jmrbZIZ8CU/WlGJoc+5ogpnvHOPJQqxk1PJQEZ25X+Ssg1TXZJ
Znk78sDmrM8nvTEw6tJEg+iA/CaCZB7sEG7z3KamgPZLZof1+Ea5fkicMWzgerC79yQz5QK4aCx0
ej1U6dNhaXJ15omGwjbyGrNNzNgE3gNz+hRmP0c2qmX4xL7VHDkaJQj7PDahlEtTJnwd7uU+QCZS
jv4iGVJLcL/VTdFrbmmFX1dsAufeQyY7P2Z4tMQ6qptM4xPnPxUTq1y6eIUQF+oUhg9CW9J0wmHp
ymcCNqOUYtE+3OX8K7xm6H8/4l0VmMeMCznW1JF54zPYi+FZa5xLQ6EdSgSC0jgHzYavwoxOfX6/
Ki84jt7uUMCU7hayAiSLoLxGjlUnDKhXsg9l2XCPSIb67whLKdWwbG1Z98KyV2rsexMHEdpJqsLu
NxLjC6PedZU+mRyL8hEjfMh7CkjiD5H+aR5kGlZNrBNGbziVVzYEqzKELHdOwtsEwfTgpFVsxbdQ
CUwaJ0N2SH3iBGcIYkfLnd+jSytJByY2/bs2tQNakrgVdXFjZ4tvMukxLCehjiOPd6vxpbbUOwq/
5YNpKwShz5HFqoPFkKUyUdiEqtTWk8A1/X/G8j/JlG6304gnukeM7YXP0qfsBgy+S+oyHBfBiLNt
Jqve77qwb+vIGoMIbTpDvlskGROZyiZyTcbo+YNrxQwPAU6Mw/Ts9S1VZwRyPgmb/HNg/vdIjXbv
7XxmfWNOXFTvWr5Qbp0hO6dkM5c/CdFhKIHRu4eKR1AwV0kqdKTdGsIzhTVd9kP0E9LPIrw1gcN8
dtkX7iE2djNC6sD4HWmEfmp7//jszDpzkyXZvOdbH4YvL+WB2z5X1WDG6RTf6uSSBDIveSSS6SmN
NK7bW9iiag7Ni6BdoBxlXrEYaH//PGmz9yijNrHX3TqbxPuC2XlXlzP45jgBYGofBIpqsPNxGAat
yxA2KMLlVmMeuo5um28z7cVPb/PiNiyz3dAr7Q7dW1hSIWwwXOXbV5ehj/OisYssljy/BrI2Mt/h
4bRsFT5ryI982KR1cpxzCzIhutEYYfQYbrr1aBejvi5uZfs5+90PFS70un8lm4XfE6Y/IOqHzJNI
vL6Da6N5t13lZe7jQnDKuG5eRuMYzGqOYVy34LsOPHEVbJQSQa8WbgpyII+p4PjWxPxcQmFXAZKn
kaPXEGLAfr4YGKcnwhucbtF6q3arK7+0r8tWFF+Mlmcvv1NCBw8SNggyAob/5sArKI4BsKAzejWZ
7DUgU3WRGR4LOQe6Hl+MagNewWSbYhATiLGqyLPhdtO4TC2aPOpLIoNc0qP68OL/x0E8hznB/Cqc
RelMG6xIxjD2FpR9UqdYzSiOvobp/El2H3n9YfnGkzcPv2Q7mKfv4XG9SZ1+3NBGWlP2EC7iSntw
4/J605fFwreFASfFqAEXSt0yIkNdoWhpblGIYWDP0ZGKOvGrfRleGhFU3YVeu+psHBhzc5QixOSS
7qa3H+7LizH3ZyggJ4Nt9SNcIk2KApgfPUiuN7dLeZgbzwK5wqG/cthe1nMQDmTImZlTcORZdGar
ceOpi62xpA6AfyRWfSiRcgtvKHUhg/oMklKTn5IcnK5+qL3cwHmplZBr7fkozZ9D+xfUlHtMw8KL
ou6i4nRFEjySbxCOQ2YEtY82+YimW0TB/jHj0HBG2f4CsqryNRcz8RaLVh3k/4R8EfeEUtCzyzc3
OLpy/8Z+GSZIzOJYKb7bUooX5FgsmAIMq3Xy4cE1IptOP8nLNl8EoZzZlmHr7FgQxKlmHy+2hQjp
kuwDX7k21yrmvnq4HrFUM6x7yHdutruw4q6Nkutp1dPwPneAL9n5jnrr+9+5EyYo3FqGB5LUsM8m
K50KA8ucyf5ObmXB72IZzLMEz70AMj9MIdpZegWVJdke7dsG3DXHH+Go3en0ArcL3V2BHjFdAAYj
4eOpGXMaqkpgjAaBhV7Pqc6PQUn215/Yc9/29INCxEu/jJbc4ScYknnt2qT4sDI3/OQMwrPej0nn
VSA9MxLiHF7Pf+aCWSya5TPo3aYNrqnPQCrH70UXJ1xCylI6AWQ0XK13um4vyN/a+DerY5dc3Id9
1QshQjRn5wVCWIr6yHUuuN8AHMfmvBbnEeq2wYQJOFAX+M36l5/N6ZbJMZ5Kh+G5wXRv9LucjIbA
md8tcX1wG8fEPGbfmoR9Vkl3ENtRqqaz44B6Ad5hcXcDfxlApHJ5C+haaHY/rvtq6TdO585PU1cs
Pt+GXQ4LU0USoaoCoSO+IWNr8bdyw+VR64iZdS3+qcKrko3vl/itLhuX5NwR2/iSDa2ko9tMp+I8
fh7R1uxu8WxePqZw5iT1QVVvqW5RZIhH/WY3CTQ21o97TfHzBkZU2nUTQZmNcApUse83hfc4M1Xm
5DnCfNMpEzNkS7y5vxpIWRiFQG/kb4e/PzQH18sfXWuukUjPew3LAX2sAFrBF2EwWTfeTpjKH6tA
b3Us6ebDeSX6+3lEr9UI7IsJVH1c9xNfJCeKmcLppDWk6lZT+h/ST0Q+5zBlHgpq4cljTEBLqhX0
cq9oSXKNziWXhDysIg3rGnsT/yokY+pPH1nRcNyP9Z335MfnjOvXRkAo8xAgV6GZXie6tlpgLyQK
XPwsHDG30VBU0rF55UYIR2RpBD9vnUOw56w66FVAGpWY55HvpCBVFk83sA/Je+jnrgilopbRUubU
LWJkURT2vG/FlHwP8M07qREoGuWo9vHRLsxBexN5g2EXrEnnNGbshxDrvXAXUth2lZkMi/d5qAkg
sjHUi1yJGSpeWChUg2PSOz8q0tF5P7HHRu4f7ZKW3L0+RU3rdIIMobzVbO3k1BvlDQn0iwPaGiKD
h0w5+mMpFmnApsXXCaKCYMnG+CNHlR/eTMgufdShG5XARkpVEcnwzXBnlVNtszXw09/zvtZyGCU7
0Lhk+0+PBbprfILKRhrk7fzLUxCrIAifuM7HL1pR3rl5Rq5MPrMdL1aYKMgk+biZLLm/ZrnveaZz
WK8pl3vN4mn7Mr3eCyuoXwvLMIMeZfyk7NsXWk/vvTBIt7Prp4k9ktpimNH5pHKxWqiwIWhtm27Q
1nQQpOwjoOuf6D0tc4qSXJzqPK6+RFUClzyBLBO55ziMBR7Ab8PyxHdyC0BsrStoRf/Zoye7lTgB
BxnmjyQsLWWytGykXxFVrlqrREdfrTbtk/Y15ZH6xQYmj6w2cVxdllfub02qOQXPq8fQPaAkjQd/
+SmkvwMEOZdAtj31Dsf+TMKHnTX8TpAjhXw8m7n23WXXWCeSC1ctZ0BKsEv2WbevthfgfUbxUw0+
KwE1wEjuDcfe1SZIlZvSb9iDUBtN7uE/kehuQLekgpjWMtCbTdx59VkKFcfQAqF2+QzezXNdcsyh
smfHrlTibnYr/YPpYjwjKtTgg1s0UHuCC6+lvyXDVrJ4alRAHlFwQvafMhsuo0G+/Uznj8z+vzSF
3tOgJqY0885/KdSJ4P7YNQ2UoCxxsIwVOIu+5D1PxEdIE9Y6A0PTa9/kkuCb56Mvr5EgH+ul7bnt
l6Nsu04oXa3BxlBOHiwWsxPYKyLEZAS485IlWV3pjTjhu/Otokct7BqKHr6G1B+GJgH4ExDK8zMP
z/3bQloqT0Ac0ITaA6PzUYkbuNZmti5/rALd3qnILBP7joww0NTXHhMQnBj4LsZjvKGGyt7YoM4V
eZ9F9/ePnSPea25jJhXwt7+jrucMGFIuGIAoOu6S83Db0O3/9fvDMEtH0KHxaiTkUeRABKTjksvL
rTimSyEZZJOkegWwrAyv9kfLMcazcIJqHa1MUALkiJvrdIT3fSiltiwDmk7UYXBTebz+D4QO9Nhs
29uEsC+FqJ+nwVdoWWZCOXihLdFzJJRg/An1xbc4yZgIWJigQe3uxv8T2RbUEaG3CMikJcdCavry
6e7kRM8KcqVFqMU7aZ/TJEh5BEFcUDMa/YETKIgLXKE7jdSbAknXi3qg0EMpaBDUBfsLVfY+YIuo
6c4OkfxDg0jPXPLELPCDrfJ+q6wdpwpCjFEy5KI3iLNO68CQywZ82qamNrPn9pZRLNAMSX28NR+0
X6pUUBr9S9wtv+qJ0cDF96j7r08MMJnfiTXDi/Z1ueUiPNs5zFZk3Py3lCmA+rpnkUeyrOWJP/sI
vq8XLphbfe0u5opQZBB5TziO35CLY8ZMMrDfzRJRwKFFuMsbuod2HpXBgvtID0e43aXFxyK1noXF
I7XgX07M/gYBWwDa1EJ0sz7tfRQvPyTnfxpJcdKclMF3J3PM0DOfF2B0qBWGh0NlacBOppj2tXdV
MGp+0J0I8To9VUj1YjvxtNuQ9sYeLxbSwyU9R1lUdE2YBZd5L5wlJH/cdN+S0jgmlBWUhz2pu+5y
lSQZorX2UROhFaH2694qNRp+DNorZHwdP22/aG0vZfxjMzkkVXBt8vFuQknoYYNj+RuXe5dgOShD
gmEbNZUPtKNnwklXiMK5Cm7OaWMPIoA1kfgpD1YEzcXHq6cICKCzRc1ugWpzeFrsozE8mIDd+P0U
8MXpITB8tA+UxwWZp5uVjsT4zcqLZuThglFA3oE+yiLyAKFH3c6kxnCcuKImjZ8NViPswTgT8Ays
vmd3kUKoCnBc9yLfEpdTy3BKMfUjqBj9s2RlQT7kng3KZiOROeu31cdOJLrCTbeKdjgHsDbKPR0k
pvPi2G+bfvVYKfWaDKWzucSNtemsBxjSAoVW9KjciX2FJL5110NobBEuE1rnqFoFr7kc/R7yYFRq
fpMve/x4k8RFzKHK1MTXhQL8MPnTNSgqE9ROd5qc8otd1bMc6D4WnltUPRa5WeCph9d72LlXODjU
2m1mdPH20LdOQuodo1GsKYztag+rNq/WAs1O5khPd++V90OntbZkf1i0i4NQWFkJPb66njfm0lJd
O8k7XrE/fr9aBhV0iI6xb8cDFsfZCEFKyLOTLRdVw2gMS6MfsJ60yG9k5GVdtRMx/GuJaxjyIEQM
f087naEaj39hmQEMjOhTyrnpnNZ16Kh2z4ucFF/hiw0KvBYOkfoA2PyBfjRuESBRJXvWRhNe89PP
ac3f0yKPIUc8VavzhRtFW2zKpm+WB4ontJepfX9YMktjawvadLCetwqV4KJjpMjhim1KMUUA/x87
7zd35Nylb8KIItI5gLvGYmCdnmWxGAAJFLLs6OVNZNQFeXrmCfxdPvbmi1gff1C4kZPOQg9RgDZb
3JOMhNkkJ12ZLjAAFCm3VSCFbXsFLjuX4xb7J8Uo1EpayfQdxULZOlWElV8tzI4+f19G8j/mslHz
pEs9B2DXjILrT+QlTUMQ2PGbFbLCVDkgmixRRavMGhm3LRArFHoqsQOImF6nb2xN4fzBy/9B1fg6
9psfwWlMgojYN9kCMMF0GtCX2EVOv715rkjawGHPHRUtk4yjWUPZa0ULHZn+A4NUxQp/7QshHe4t
J+Gxiotyofdo+KYeHtGVVSg5tMmPnv17gX2zWMshm33NbnaUvUqG1b2U7bhsBQVcBfIodkmfjBBO
0C1DDptIgFhkIc2+O11DiaNas0Egams6lmpGWHJeSTbXX7VpqyWN2sTp8XOTnCvekiE0CEUG7FDq
6MMHN4/pmsGlrERo5bzLu7zJ58TMupFouD0b7rpDfvKRtr5IpV32r2IoA6MDa42VFZ6B36f4TKIn
CCA0e7feSYoBmMwbPnH132G5Go0vnKuiMZ1zpj18sQWDbVMe/4y5BV3KEhHy97WiIj9Ypl7Ux7mg
eBNcJBBEASITFmpNp5Stay5QMf1c5JYtvKJehj56aU08R5gzl0RQkWprV3b93GWUVq7Ex5E1GHsx
vOiTla7WIxW0V9D969QX8sW6Ul28Y42DwPTg7C93qpF/guIthp+Vf79i0l1LsU/lN6MjSRvbEyVz
2LDDey7vD2ztseMUPHcPiRhaN9y8p8YgRyfMrvQdK4tJJvYqnCbtbHuckEb/ptUowe810T73gKXH
Gre1IweYkW5YnxdREU99QaYQlJ+TMnNtW6ueEYb9uxn8MBu5iYz9Bm5LAuFQWigb0ollnYgnjP3W
OKFOFzxxnFtj7PS/Ae47Mde+m5CvlFoDZmxdgHu5dZEkSnI0oSRTd+/toVcQpA0N8glT2T75JZB0
jIGYqeF2scAl5HmOLK2pDWQCEzVXd6NHUQNmTyc9LZz2WESsUwGA+C1nLNa/rcvvBwb4PZSb0Hbi
IiqkGANGqzonl1GfmEs7OcogOsqHqXetg/ZnTv0YOjhkNdIQgG8IKdmWRxdJJ3jzf7cwy3XZd+Rs
xRzKlgrQ9rZFcEUvjDWxP+eKT/8XKAfEn3OW1npfWR2fHKMEKD3M9T6TjV+Exx6Li6SSG9IzcMSe
jt7y9GuD1ld17P2Ij6xok5gVQeYfLXZ0+JjV8D95W5fRiGPQL+NwOAoN0wp27Eq4ocEYhFlL2vFG
KMJZ7gjKWny7/FeoDgXQfwp9h0vOkTOr/fKceXK6t9pm4i71i+7yoJLsLGPIcwABHQUjBfegAgQK
zmVt5rKTJCHEB4mxyRbFo6u84iDhjtA1fKz5wGl1zjldVPexRpeEM6xakbPHQ/2ycn/8xh2fsZKX
nIENw6ke7r19gaVhRvsm5V8zix0HxpuoOBmOsjq59OPIp5MIuzSYjccCeZUrFhho7Al2PZCT1BAN
61/gf7rE7Bxw+nQyI53qzG8P8O0E325wzhfVls1mFWwxlS5dUKz1zL1jMxWN8A12XqQi3E8ZKPfC
WRfZrj2Kiay2xUo+srxUsop5ZmyiRdxOt6ee0Xa6zbI3pTKccz3LLR6bMAByzdVri4NY95LdBLkM
1p2V1Hq+g9VWpcZMMdaipq0JBMBf1KhyxbHub1SkXuXrb6bmiRsVGyEPk/5zc5ovZ6qsEFyHIR+j
S7/aiKcN0aAUgiOYq88lBU6k8qQeqYnB5QaeVW4kisn65CEJGCa14em+ugCz5+w3x2UM5/FblyeS
3YMSDTG0PctNXlSAU/vGiofquzGEPZkHuTG2cJ4sVy4Ub4ast4c4PQ7i/gLY/IGoXEY5C3+OkewU
Bevw6c6QrQP9oJFkWdKfl2+fUpAeR5/ZYFHrv8+l6t9eOvLXFB2uNENQrO5KcPTwFEvmKknT8QZ3
EZQGTxDyW/4jGLn4s/r1vGbilwv4UB8wS4lcIiJ10/osuvY62SBJo8fayzMmHaXQQwJlx+zwOqzP
kPmth+XvLHQmXjSNNhbV1pZKk0S/tNAdPyyVKkAvlVD1pzPStZ90+WfiPOLw6rgOy42L+WA4cDPE
b4RyE24kYSyVQhRSHZHXZi4JV0hvL/5kDolwF8DZuhNPWQCpwAD51Zwv2zsFYd6pDGX88a7etcwM
deMTl2eqwJJh3/l/spvbllGH+i4n+eRkkm7e+xflFtauZkDSqZdEojPwdGQwt4+WBNQoMOImaSDr
E7x5dnScdBdSqjhMA86CZFRVUmwb66/7MJA/fWnt11xAjBS23ptXBto3b9zti7qtktyb6nY1rQ/y
7QB7TzDJ1kdkBdSMF3ZCE8w4053jzM+RVdxC3wnxYmYoeC1CPHrKc8ZsNaAB8xBnkW355rU89nj2
KiftW9qANpHb6RLmGhgYdjSRA3AkKHQs9jnrZh4DMXzFHWX6OaVpEA7oKrdpUtd6MYT+dbJhGcVS
axwzsD/5C4wNrl7If9KYrOGM7s38hzKUAsp27GwGq3G6Dm2kP0ZxuW3ZB3n/Y4O/REHeLvaBfOk7
KkdS30nB83G3kJSqRmXg5GmbRvmoR2fPG/4Z/HtwHIEdNJs7DYO5PocoZgla3v6hg+aKBbQkhn7w
qegicsscNVdtFLdkj+mEu4YuihaUpKvHZZ+dyuGvXjqAdveRPlp/+tgzhHhTkpBUF/NAb806COW3
5PhSUUe6jpjlw2NuzxVkcCBpAfTVSxY6TndY1YLG6nslfl1L/uYZzdOiMcaHzKkvq8aJR+4ni6/P
xfx27lVDBX9C9GQ7cjHVrgxhqv5RQicySq7wgQ2Y0RcSfGUgLn8LwEm74L+p6A9blHiki8CsabMQ
lzScQNnEzbdaTgWOMfcxDMqkigN0Sj6Dh/FkS/FemCzNDDQU5VpyBL2sfCYvwMKIAe+vu36sZVRW
GCLF3Gq+/GPGNQ/RLsYDgu37WQB2f0s9uuhIbZ26sp53aq7EISsOg7ML1uiBGJQjcOTvy/lUQL8Q
nGRQlPh81qK9Uf0/qnOs5SOgycFtqcwmemfZzfSST52SqzaySSxdh78QTGVQ7cbJpPXA3aydMBv5
GbIbckEHmLfP1SQPolgo8STMH4V1hGCM+R+zWOX9rQTTmsBoJVbXnz2me2uv+NSSJf06tS53i/lC
rDf8i/bMlnarJHZAtsYpVir/U+XyANDHLWs51Foatc7EgdRsjcIjOxvrISwe+eWSw9HPcgRXs7ef
HleLx5yc68y2PijdOXbuMMl7XbKaijdMpR7AOffuU2/NxrrurX5TUhhBFcwutcKev7Xatf9bNemj
cAwZooS8kDDXJK6CtgtDMfImgea0ThRJkqb3L4ps5aK6+s1BuOxcNMxclRKmymyIvqn7C4Sn4jL1
PyVw7mL4Wg33gpbY2l9tOQyD6YJr/No0WNBxL2/S81Nox7bt2HRU4Y2bBojEWaeVrbXBB/7iUbrF
F3rAxY7i6cvk/lWt8sHPXwY2WHiGnC8ijuXhc28wxyILTAzTewrcks0mFfCIZL00G5idqLFJ7okO
IZn2OITO1soc8h+Jy5T91QBuj3WB2cIInzvIIBt+s3H9n8/NARm7p+b0U5YTYXRksr53Xifpn69P
lZTjuaoJrQb9N33VTg8Yos2sOYyR6c8Lj3+6hwFS3mQUsfLO5ZrwJDYxqVNx0UbKjYRd1Ti3FlRT
0nHOz0bVsjwAfAmxxoIFbgODMjs6dt6jiqYffWPNF5XDwv3fapiwhF9hal4LlNN7v9xc2KkK6aE9
VrZVK4nwLqmici4AFJiQBccnXAKPRDAwcWtDSV+pWAEWC5JdPrDzpo3WKPK7dz7IRv67fCE7ycwh
djkaqBWJH4kkRNpdTvo338/o+vO6nZ2q2gPQRDKIzfM4chQG67PilZTmtrE8vN82QrYfWDygcH32
uA4g7kAe7tSRDnYeKgim4aVzvWNLx5LpS4CP51h+kAUaIyD096qDnSdVrjaG2haPYwsv9ZDje3b6
VrducqFgbDHvq0NzRIY0JwLNpxMfiNXzk/zRleulZ+huzE8GzpZVLc+qHWzsuu/F0toJa1qhz+d0
A+jhwq1r/qxAyA0/WV58TcPEpw6tMfwIzpGPULDjUPjiltu0KNcP2dIcBLWHZbAE4U3MQJgRcFgj
vae+zTeT4zSUjUs/FjcNFsss2taUhS+fvp2DSmrnURNxvUu5piHcE/zGLqdP8ll1rRgf+JIKkvLX
V3WsZxn+uurWWQLTFdeh7vV1MP510803ejLrtGp4fCo6UQgi1sPvfYPGC+ghN5WJ3zDH+QMK48BV
cv/Bh5KGs0YzI6iQV3wgor2QCJPAGJnSgsI0Ux68RTDyVevfBzDOXuS5NgdIt9Wr1QwmCR+MsaOg
iXYnml74xf5GvbR8HdgHNNUX3brumR6nke1vfV1iKe1fd3e2xT2F3GdkfzTam53vrZktUWrVrHju
J+DGdmR/GrnoMQ1dvd4/GxX8PXuB1xeEOgDDPOa1Fd9o1+DFlF6ajbMUZazB0Eib2f/QlP03C/Os
9/sArJERC+qICQUI5nvczwp2gAPb3bAQ831RtqF4JNYm3Z2uiGe9ySj0zm43C8k5r9rRoyCjbrDY
osAGBc0Wb5jx5JhpPAajELSrX3YEYOJe/eARxEYQGezmO7kXKE13iNXMDMfouR3IKMhbFk1cDAac
xTNToC7crwbEiYHsTY8T/d2rqu2ya/6jF1edzSiEy7KqUrPb6qTWJSEdopJhbEFkFT9kf+BvQmZC
WBm/o78/MSZakZXI4iqUH131saSeo8xGG87ILryvodCFQx5OtcBTtgQVl5K57GsuzcqbvQo400ub
OrAqt1oRr1PgY7VPhD9QT1/3/E9Jbd3/LHCuIktM84WTD1WkXN35eE77Cz3C31Fg+lvfNePtdoW6
XmIIScGPr7Q/XqOkWyNip83U+8JaPLz4ZSl0F6huBPl0X/XvKBGHMRcr+tUpy0XcaVk4ieLDAvHJ
vTFd3h7aYcVrpRntrW9tTDPmv/As1afDBkLDHsPg3DBBOoexL4kr64fHB4nqf82ulxiwvTXMjS6G
cSnHvmOosOztJtehKnJfFD9gTN/LFVuCx8C7/GeT9PaAqgwo51tDazyVXjEcI6an7Cz91IzpBA8t
KCMUYorNgos7ODnYEofYndq74SUay19UHohPcgCkSwVd1UVzFvYUVst/9E1NtvDZcic2GUGioSIb
lsrZqciiG0+LLTuoKADgO1FyVGQno3dy1nO2artZdauP5VgaahnXjsTGbjmzSJ2M71GDQSVgkECb
OJiu3bAsdZRW9GQMHL6mhJVcEMkG41wx+anofLmvuTyMldcLK/P2bToOX1X/ziC3I9xDTvdYGz3f
Yffdnyzdh3jx8c0mOFQUflJxlKi/FVeXprZPSbBY+SCj5yGB51cNWg2wSZMW/rMqdro+5ueTl/hA
LX+XLBUt1H2qM4d0q45LX6AdcdxydwQly1XH+Jtv1DxFao3EKXrmA8//ANO2mmjLJs4perP/43TA
xcipcn+P6wMslcPgt6liOypkroVAJmbiu8q2ywZ3D7KqognBS+sQKg4AlCUoMSM50icqdDpLvvW3
J8n7E3REQNs1hJZyyk8Sikfs3+6nDB3mb/2iqaLZgsoo/W1pIiTLu8IwWDPH9+9mKLemlsJbSJyj
ZsMxV1cjIMmyJXpsQncQc6TKAYJXnOFPCB19rwgQlQuVyZD+lkvlXftywaXu3V4jhHHR7A/oGi+z
iXbeiaq5j4uCkCY9bebVdYR5I03Uq3bzyvCYK3u9js9yV1XqyySrKEVf8W8yf3f2k0SQ0YUr7+PH
3uY3mwxnBHaCna5BJAklf5Auu7p8POpYplF/gW2S39hU5+GSddqW+igKmKnuDeF3aSPpEbykx2Gb
FD+TQTcTat6lrTCricp5/UIy6QcruSjITj/gbtMkmvxz+oinjijaqWqpM1VyHy71GGqd1NTMwHwy
IzmQSK3ruO3JHE+bts+h1MeruOHS3sgK6w0iU7VRjgrbQJO0rgkjRpBuIy0yQn0E0Yde1rjdjVSG
8+wQYxROnRnSGIMBHLGy5/7hMuGi887tG7+00YEOBZo4buYmbmazaqQX9OcQM9VhocGMnnbfUD1v
iY7vQx1ACLOCMU/BE+RlDKRVZ/hzMO1xGL5EOcJPA78g3doX2KXT+2KRjO8vZjIN3ErA6eACc2ZF
RD9A5C/N8KPy8YlsVWX1ASTwaNYzk6eYuoXN6/siOJShkTldNMZfEcndd1hneEWCwNj3Gg6JKGy0
3K6i1VrLac8VBGmbd81zNA6I7tOV5Xn6W1Hgnz4XCJJkmx8kYuZrIEKuwjOU8gAPJ5n83s6TZIAb
nakaPULjJnCgag8vz4bzCKzMrrWQ67MM79JU9uhQxMiFHMYu/UIEEJ24cjF2zc57SevXAAtG2uIr
PiqXzkp57YPekNlJt+HQ0bY/vTOclSudwA7Xy4txmEPLN9hpKY2+dXnLvLHs4ETawWnR+lCfyBBG
kqEwisrsBiEzZpYTHnxvtfxcdByRhi3exHg4lLcGfw1644qp3knwtxtVWzS075HPkKxdfp3WnFDf
91O72JHNN8aQPXE5aPxPWY1KO0vQpk/XaS9zvMrUH286un7sBcVWKjJX1nYBTbGsQKcikEVZ7bP6
9jQfDofNKeLZwcalPCdq2OrNxy2dJFvYzAgcYWRvDtg/+TOAXIiZjEwoOoFe0DQU7H/owKq/c1fh
2FA0h400GWvDMj9JxGoKGHSsIodxHHitcN1x2Td7t6SyTLGr8IgB9gEJ0j6SFVTvmnny+oeAva00
M25vm4t4qyftbcgk0YOaUT8Z/zQY5hs1wfgyNzNcqvK4aPRpdL8PmalF6lUj9ILH/qSRVDV/3dCz
3kgzxidFKntcs2j2RdB4YDoUDqtKAnlc9eOw5pN9s8poUITXFgGJpdfIsO5PvLI+bA9/NKc8n1vf
xR/6GZ4pyz/8TvuUPlzF2Yd7G4JBtTzapb8A5/iu321eu7Q1qilWhPT1Bz8V4OAiso9/d42To4pT
OSA/m4WuLVoBO3DaaVkM3LwrJmAxLYCrOW4/uJ0EuMLp2JtVtvfm499zEH8YA6f+Z68iFydJ9heW
psRJRwX5JEo9kjWtlDaAVzwwgfXtzcaB2P59/MGFY+CXxaue7NxTGnGYkzxKwszIU0gxqAtmw1Wf
IbJBg7MUW3g6zmJzD8sTKqH8fO6nXxeQk9tm3s8lWMiGWC8xij4IogUpUKif9QtRic04SKBoTo4Y
xtjKRaWGQ8dp8wJEFUiA1f0889v3yi0/zdCDh7+0hFfjfYbxyibCdtm7O+iYNC2ymIwcK8SoP0FH
v35MIm6oWFWI2ZFIvaCOGkEFXRYMLMwMIZlE4ecIS9lVceUp0bLCXnnRTuHhDGFqu2vKcN9oYz2I
LJ4qp3Lcw9HXDxyeCJoQZ8WfvTnrTle8JmryUjG+gNIq0Z/rCckZlD+BhKYsfhpdklvOoHYPg/z5
XvXiKTT4oSf/7TPbVaK1k0iIdm1fMM/VxiWTALxHLcSwSlGXsHDGjFv1W3ZQA41qse3uI9YW2oC4
h1FjUdHM9Ex44QHgLhYzrPAKJhXw/TYQ3GHrLCnMYrVXGlyFetmq0ToZ91GRwssFJlKD1QXlhQGU
LLkxFVLwtdddB39o8f4SXGQ6rWHhJyIufhwWebFW6b3RqAaWhOWpLCtK6mha0Ymk9asBEAsJk+RP
ajjl+imm+YaERcALOsIAlh4cN0i7Bv6Ir0rWhVv4ma4fVlXMJdAnhXFMqBYMg5pinOFsn/1fRtNx
r9wFgfPNg9UIaOjG1yoyf2ZQuAVTfwf/9l6BjvjOTn2B78HrZVFAhbUem5hadTdHVcJAM5UtoNfJ
4LU7fg5E4cSdw1gMPV/idr15gwpGpf90V9NF1bKLAuHwvjQABTQyVoEwKLOmr0tv5CGGP5Fo2YPN
6zl2BiMks7r5SdoOfrDjbBgbH3gAB7hg43267EuNMQ/N2lfEnTeHW+/XX7cgP7VGeLgS/aGEgAO9
/xK7HxAQ+1FvT52u3/Iv1Glsn5fdQuBSjoKGvY2ssrYz44xEIg4rK2Dcko8vJIMnHOFaCYZUeN9V
Anplbnh2syjuI7AiD6jR6lwptxUYWqsNhNRG3sQ+qlPEcA4w2AYP/J7Yo6Ip2q0bPZvR8NNHC3Gv
6QsCOX3hchW6O6FzbwzGS59UjzyBnMraIL33jRDg07NDTkFdKO1DUaWbVEqaxd6+0cb0t+97TOd3
TnDf1Ib/BL5Sj594Y6DMxGavKkCsdBnWYT5SyBQTT+1+JEJJDDCvm6rZ6DnOunXlaxteUg1Ywx5w
FeOjNiJ5Hr1JXTsyunlgcOKBAqvz2ru863uuPL7DADiVok2lx3yU7nijz/Fgf4ctjpQYRI47TaFi
tfrh5ff4ec8QokBvFSPL6JIsaozbIDms+rAyl/O+9QLiq1gVBk/eBvnQG7B6zbDHW7GUfPhWqYHl
uczpfc2nH4+P/IhX1jqyn0qdK4tnDRVa1AdOneq6eqwDBfUyAb2jbA5va58Eftt3b9Ppp5HNmlS5
vKlYTo/OuG+Nhy5Gg38/txEg2TJEojgR3YpH3v4n4vdY5ovpuCrRYFKlykSQ2yW342h9qPwMjREz
3w3UOkfrka/ATxFvXYnOJOlWYxnZyQh3t/Vj08VnU9ngaRzmR0bbk7pIYUD0CbDNges+r5GNJMQI
9UEL2LRdBd74UVh81igSEUrbURKDujbCmdHruMNtvJRI/4Zbj6p4MzoZfJR12sn+pUOs9rYJF9Eb
q1EwZCc4ktjwonRmyqc2UXmMqFkfUwd7D6lsu3IH0OYW8DYRJLot4jUPj0lF6xmkHSRFlh1CDWDR
+rBPiH6Hbw9JnbqvIpkHdmKDme6tAFrhcjMySo8tOhmjGgqYnL2ClbR7Ov4IPzj9P/+bNBH0pife
HLluHw/YuP7M4riercnl7hFr6BJPSlAZJ0oo0pXF7YCHJBMXgaNOFhAIZ4cn96eXZx1qnaTBRVBs
GBXDquq6/TWcHzSBX7+JCBr+IesR53v+gep8obdbC3Hbl0KZw4WGpYid5DL5uqv3TkeMHbXFYIJN
/DwoeiTdu+flRY6Bh2ApuDgbZCE66CHWNlrIN48LZyYgJncAlVnbfM3tvoxljB4UoKSern7laTcj
1wJEZfIrsby5d38glKmk0sXB+h8DHOY3N1TAso7H5zjKPxFLF+hCo4p/qQEBkc2fRkRyI20r6sPB
mtr0rd7PeKTDr5VGDwqOZr1YjioMAdLKL9Qr5OZYTwKVOszC72PCd5PNxIZq+DtZC/EJkWIVQzog
+rv0VMDQNZkMpkMGCTfhN0x1JMbsaImiJtT4qK7CHEDgIPHB/b3ewKnFP53M3b0p17vAaxHQOo6Q
hMy8k+zr8lrjX+JNHJWXeOrfq0wjvlFpwBQlHPYlQ7XU6/fTiwfpVlA30CWpHuwF/YrmprASryxX
Ezw3CyDKE5kEU1Ua+3uR2Tgn633C34xiozMYnywe03FXRPt05vD6OY55S+cGmfa3rEJte7WdcUi8
4KhKY+yF/WpsE3lprnsDmWSa1omCYA6AFM7PRkBRRP57n25tgkhG1spNGaZZVp08/LvTQzM/4efb
n4TSDcGyZFPnH0YPOMiG/nOUxLHEGcT4BM/S7hJDmQo0r/C9OXNruEkpMjYTSo+Xa4DXF7yvUDwj
wfR4t3c1CO3C4/RUieiKw4tqwvQDUWyNO8HHKHYYJO7N+ekIsP+bSESoZRoqZb7BQTdRR2KRIYoA
+Ba2p25nSAoLbPchOYmGlIk23Sfm9ECOZC7IgNoFKfN49axWP4c1CPBRFBrjQp6dKjOyZhtQ4m7D
ryV3EP6AhW2E5VZkHZ4cNoRfGS49IKnusc5a+HRM1+AnNPt7sLB6A5Zchkw7JS0kILnd1keSdGQb
vqkCGMuPslmGHo/Be/xBOKLY9L5wja5xVteqYi1dGrr2wfJgCv4K0SLsIWV8D9AJL5tmA2QcZ3ly
+t0/trp9aLNj6r9/RWIl+e57n7JX+KStH3qbWXoEjN9Af67UM7vOzsHJTdPyz0DiVgjpm0BZZVuG
WjNJFWakK39jDawRm/UD8PSQyn0d6g3P8S3fY5DDXS/1FgPhYgjIjVFY+Ni6eR2nphqWlOU3e9O6
v/0AScCjGTBhdhXRyBFwaGw9uzVo4R7dcafCXk1tgWwcAonbZ5QRrJG+bFxcNhZs/bwFnuG2uZGP
vLlWhfjQ3tE2n2+DLeL6s0houxRX8/9j4yYbDODADAialdW2Kwipu0V0qXfYYF3A5CpPrOlSh73f
Av+9aBDguN+OSF2DJFyOOx5rEikoI5yz5Cm+tErZXGb8aqqIDM591yw0SPF0ld8NQiBmn6BbV90g
DN+X7aWIvIdecXJWAA7yIiGPpuy6ugYSBYHodTBBjaWyUwpayEFkjOZieUESFJ/5fpqe4pdhpNc0
2Z7fAjTQgyp4PWjsh4O8BhndGul1Mm4D+RuesR2J7oyDRDwUkVDPQB0NK6diTaohZdLQ1mC8IGQu
NZSvLcjtFwaqelsG21UrmKa10VdoKBs/68d63FH6mIbcASP1MZSykaLq5Mia9vehlIoxPPTUYcmR
/89V0XDgQgWSjc8uRtPyauJhk2ZOdCAmmgOx3SvOWm2tK1gMWy+VtmtLBnwW8V0uZiKpWoJr3Wam
qWF5eZ65r+q3uvNkxCd+nda/4n+SIDtCFtROVuAhgkJHrZodUFRcur1DFmvagN1Xb0NQoZacBdsG
oh3xBBn0usaH5qCDrRmn3TiN9OU2kQqySkmRCCiqcmK+87Cvjda19H5tO7r0M09CwTM65xPC1+vV
Z7dnwLtYFEIe1K4vyZxGSehvrlaaAQYSxmaHHtJn0bi0zGS3TocuEhQqveWYcTOmDJ17lw30HRJB
kCDcU3ie04gdGkZBHw5Tp8bcL++cdpc/iHiGiWCGBOYXXfZHv9JyYlAOCLhRMpUYopGdAn1CSFjk
m4CGz6FuQMMYya0Z5r+9iVIJvghxQYqRNH26nsKELCb9PnN2AzjojmfzrzOy1VOE93zykcWFNHpF
ZkOa6VAX/TJrbNqUcoAwm2o+45F1kq04pvPFHyPaPlk/C2NAlbZ85VglIQEm/m3v8Vk2vbKnUezM
kBgLART22KVUMZrefr21K/kNx00Ap7xW7gu62mc4FRcOa3Egxq6XCQq4WY0z3Htf2OX4dm9kccuM
sSdEASsJMOTGRPmSkN94Z72qEE6bJ7srCMoR3jTcL5PkwfKQKZnuP5NVRNKM+CailEn6kK0KAzoz
OqbJ9Urx2g18dEdbdwdxW9GCg9sOm+bBlQUMslthKND75hp0dO3wrm4h2U0rMrPRTqvWeXfJZuUE
jTG7sEigueY4drn4tELLspvmmAUFSKlKHqnFBH72j/WjpqfB4WsueZsR55RbO8OicaNO87REi42K
gFBgmdWUeRh14/g3fc5XpSIeF7NhHn1Vc31AgMnlgODLjA/qZ0Zk6FnZ48fUlWYRFvQvZHjF5Dy4
ASwLaoiyC2gMsn1WGV2Jy3yx6pElyEH8ukYPpQe9aWLRVsYNz1eFmn8MavGq8zWOhMRlIYjtTE+4
4aPJq1nU95kteBftQ3HmVz4mIyOwMWwwmGha5G4S71R7+bkX1ogfDZy2Oj8JmI9ApxxectTB2mTM
jpFvIU6BVJqgDoTCqbQ0azUnMMqTBo4rOfnCFPJbYwlYs+8aVhwVKV8UxhdicVpiR8ML2yRdNib3
5GiUikgx5MvMmzEc4ML4cRVVBdvOB2b9gRZg/zvj8xO361u7V3lzGVgi09Rfh6aFx2bQAqoXU3hU
LNOvB8yT4PUAUYicoBDVjWDL4m+DICPPaWV7U8ONsYT5s1aJQthWlorYpz9Wb7NB8twzP5TCJS3N
AvqQ8qXh2ldc6quB/LFwg/+NBbHDZiDiFlObWyLyevImYkDQtd5a8vB04x0MU/TugU2oR2Eb4YcH
BwmIouoq9V8NpE7M+Ow5elaWHxo4YEEwPpmc4zJ7HlPHrglK1X0gHt8+8iNAuITV2t5mhTG4YffA
iovcuH8xHjJpCWn4xsHVcSLyJyVWmNh+qEmLuqYJxf4qQ9YBRVbyD8YKj/Vs+K2/Nd1CvS7O3hKV
TjunARDerVPrrvablOZ3OUp4SOq6axEwVKpPBDik+uVJ7kAkJT2P24IZSYvsrVM8cu57qFcfX62t
KU9X1DHb/wV1UiR9DalFKcpcLwQEMpHKrIelmTdZ8lEBqh6SErd3hrDIs0+tlLXrUoXjxPBKXQZu
Sg/YuMUalfAfiOgt8PBX3daCLmJGZL4AvFqbVwY+GdS+sNT7nu8wkSiXSNcYqoLekg5cKj3P7AP6
+gAjBMwShPnH+6OINMZ3tsHa0fAzytfeMQfmfZCFQMnmsJxJcDNmKY8Ix1cCZ58H3OE71OmHC++9
EP0usFGiB9ZDpZu7fTeDbv2oOo3HsVRq+vz0xn+qld6tBWIdhk31eaxcXwDfhhq/CxnxshWPYCVv
zCqOABCkTttFsuyYeyEuH13cI6QVQ+rb/OM1/wXCXpnW1GEQmDiKKuqQKWl7eTAM/3vSlfDrboy3
GKBpyCVTV4bWuQNyRYJnNRwEtSsyhpoE8TAn5h023EAaypKHHFX9FXTwUahLr49FLevZEYrIQG8x
RLaRVFxmnZcrk6tVKKH4/HmrrR/ek4IH/Ca2v9O2NdCTGfvDcf9xdP5y1eaeQj0V3+zWQdLm5zN8
lkXCtg+SSqfqAlGxL9lnVkke/xIcfwyawuOv/Krd7ZBBe9rPl34O5603uxiXLaHQqmt3DsHOkE6o
n83ipM0j4BYfy43bDK4VvEkDBGIo2P5i1RhbPJraqy6/t/Eg6JFrstnELxYOJrysdmPLHmJpWDcO
aNu86uSTN9LMyacaQhc6lPCL88LbSimItGMuQGntLwf4sGxD8beXL6/CcWfZ6DE8G09PFr8OFind
IBcJwu4eEwl89pm/f3aQZFeb+c0vO+5UEFuKLogROi1j3lT3NEw4Q47S3mXZwS2R4ZQUBIndF4cT
d+jcUKim9FB8eDyrC/OgsurnpxSyD3uCUB5tRb80qthQHe3xT3Ev5M38qpxZJ3VsHcznC2iVC1nO
7EAG1ZCrZ3kv7xo9EBMExtKu7FMXLFpVIjYdSFJx2jl7ps+zHR3/ledqxnApmkubpJanJOm6lw34
4hAtZ8fW/K2M79J5TeYj8g+z5h8Ma5cPuaCbQxJN681TdUCgzK3k9NaLiwoFUFSJ2Ornh5sgBapr
FhB9gSllaVHhjDzNlRXItKhBOIFbxeVh60cg/ACDPjCqRB63JcfCP3wP/cj709kDpmAf+KaRVOhp
V4q0mA/LwhKUEBKuFJ9XQvV943nnx7DnaUocNuJO5r0ABbbe9iAd0TLIRwtQHDjdsDCs0Xs8M3i2
RZY38yh1fh5DPUOpkqPpTIwHvJUoe/nXRxYUAwuJv4hy+VI/v2iY8/8mzCXckLEsPu6/WlOys+6v
6IfbQA4cDsyTxQG5kZAapRZkstGPClZWM75cz+VZbtuyxiM4JJYbjxoQ9jGUrEkqG70B4VgZ9o6t
AhrKOkqwNHpmPIgt+/eJUf02UoQCz/Igk6cSOqd4Sh4c7fezNEShNzzuY6fM1T2UGZhq/1cYg+Tf
KicD1iJzxxmYB7sxFJnfirzZNV1KalC/h/FdPf8BNJXE7QU2a/DyMCdksPRu3yOuURHkEYE/YkYW
BS7oqyXLEo8i6/6E+1EzxU0hkP74AnLAwnyXLGkyvuYbKF/mPuvYwYIqMhiBvkcApOX8UQ/s4FO0
s9oTXstLrEhqwv5m3X06OBcUHc5V7jRAWv6vVbrLeZCpdpg92wTZNLLwN8hU0E4SeiEi1jXo08o8
yQ2qUsYCfyxlbon3xcsdVhssll7zi0/mC734Ec7ncDVgtQUXKxvffQs68IFGI/TRQIQTl8pVwkTr
4IV+frkP+yl9g6RuuvY1DlyZczb/OvQfJEFZPkpJUKCZAO91cjwZyJyfxDKtuD8TiTVRopKJCAxb
j0p/33RAqqJeRLnPzqrISyS48kLbdD61CIcdQHy90dEVKxlSkH9ikpnZ42/hfqbeYZarxa3lzlXC
Ejlo3wFoRRdjBHINAiM9Av0jCMdy1+V+L+c+5EJIjiZprMQOEgnBuoamxnNCEUhDUSzIepRYoYbL
zCQYe96Pa3KMjMWQva+yAMgXd8KgwNygMhVOHVzEw177w0m+qG+oLaGke+w/tRec4Eto5Tzap1aw
l1kWFTHbfpzGaMbgUrRR4G9zFEXXeLHpzYClyLTCaTOWj2OKKEYmiYpxH7CyrrIhCpqovJzoxfjb
FGbO6NeTs3Ptpc6Gww6/Kqaz8SUxCQnt5FsJClHuzybLtxciKB366Ud77385WOqPsD1FEYjNJzLk
oysqoI5xvDVPVkwUdBJDZ/1Iuw5tCtfKH+dZoFKcqePbSkm07APWDIKteS9q1i4IX/x0I0cGMYKI
NcM16xNFFuOSDJyxoGpbisKTRzOmNjbCDIOc4xIrAuRVymZTpI8uLsyn5yMuzG7J42rZFsuRrzvd
PMisph/4vUtxXxJrKqfHzw3doZv2T3BeTEL+mXcRMtj7eHMXhQJKESfMuTbRUuIruE/i64DUbeWo
HSsPN6DvsaigRlOghbsrvUnyNYqRMZXr7rIi0E3g/4v4pisykffckZhfVWaGoag5RjM8p6Gww9Eb
K5m7r3pDyogQQHGILjk702tIa/q7RO32yLE+WuOueY2TwGogBmDEStRr6heNtIfE0p52WHxYv98Z
jWIaOALhhe5m41QJ2tHISvosq10kz74l6PuoVM51YI1cMuxMA4iqRkX590/+vyBVsygRItCTey0N
Agzt/L1iXUUXBiiwilDgOyo7ZM8PG/qYVcqssUr6ER89eO7zID0GMmTd3h2GxF7FQNvkFtTaeJjS
3qQ6nL0iJaBwaWDdWIakHQrHIMxvAoqsXKMZD//IoSi7RIZSZpoa5SycjKZKRQyRpUUO6uNA5uDf
l6mIFGXWTWYuPwoeUnROsKEGEfx80KY6YL94Mc5gHLmpECIZyhP2VjVMzoS2sAukESgxpkHNidC7
8Ub22j9pJXZbBAYgVLVC89KrEYvTLrZZ37HXjBrhw6qHLOOZxF43Wo7FXsZMcSbIeEkqJ57YiTzw
Y5SYE8LbWA2/ZXW1Rl0muLIMIWJUQ3qg0XRsDX7+UgIoJkXd4yWt2tvanerR7un4EytO+D8axxgf
JxfTYjlZcTt4xN+tt6Qwa07KrzGwSyqI3I72qcFKKHN8L4RPmJ+XCf9knjibcN+adVsq6F7VTN8L
VsRmJpplArEIq0zXGgdho3weCgjz8jXYQDD7+tEBMEgXWcNlNYENwvWYEuiwToPzwULNRjlNOufE
Y1ab5yX9gcziYCkP2AC1c/dVTrztGTHm+wpck9AR9iGBa38Qbfs4wVYxVvHADvqU1I3P3A8PP6Sb
BxBdls4E/KgJhihaWphbX3zxzS9VDpgDh1zVL1epc6EdLglh10D3PFJ2lgRZWtYvaK+3CdCpqzLP
GSSl3ZGz1GSXlH0IVyqxuwZYUSajo/2qg1VCGlDiE/LQfFiM74yXD0B3gLfdMAfjNSySKlWy+8KP
nKEWuBuO2tIEF4rUMafvX1TTexphgLxILa/T++nCMXsIq+V8JnmkgBuOHswXIku2guGjFLHcS60a
wV3rQuuQLQpVKmrcBQpru6BbeFsMnXwwvULHVXgPPdghzbae/eWN+BXes2qnRQGEWfcDhCGaRy21
CxXm+AOsrasbN4YZn2m1juTza2D+GjkB0E/ng5BiIvduuK9g4h/bUI6BF9mUYBw+j6s+0wAlXzSd
rrcqv+6mgeVXTRKiGhG3QRbM2GbdDsuWPT2H1FfdkGXt7w6EWvz8rzbA9n/nSRNodyuxr9ttI/d/
10PTDe3ibyYG0HQ6lml1QipKeeQ2r28PutJaNJ/w5yxnVBVQnnwM8HBzB76bg9AcOF/JZqPTwt90
U+Or0q+FEt/GfBuUQ6m1rfvjN21APIsIUpWs9d38kjaLyPYYrYWVSjuAAyUS/MDE00/kVYpRWwpc
OzyaTN/EonGDSoHD/OXdCmPmmYN95BdO8dkVCo4h9DrwEEBvFo06FRJRCvD3J7FKCbm/64Hdm0zY
v4DSU1O+EzPxtN5WnVAqgC3qtYC3uk6EIG55AYD5W5oKGJDkChXjhv4RY6pmmKjWKBvFJ0YhT5gE
d9WGVI+2IngGdSJ8Bm5Peuyk2uTK65y7uChTq9atM3VAXHxAw4ZdFgLxQAgKY/Uf8QgVD4JRydi8
zGiW0qp4yY4ZLqYEskHlS0cN8HG8OosnlkP3aQ9EivG70Y71lCUpNyq/VAVYCXh3jZC11IUKgS4V
Udc5JisdNhWgspzdzRJGKZI3KbAhKgjzgQu1StmC0jecDVaCYIxJf9ChlQqLXj/ewoKoVshxmJlA
zQ+9kGa3zE1ofwUHmR84b+eP40ROXXLAsWq+9mx0M1bNgfSVoOtv6NFBbvg211CKD+cRx4FT2hFL
exiylvnUzUdDgK7tKirV5oGavIv3RL/RaT7sRF/xxUWxjmh31b5/kYeVFc7yeYo4HUZDOgazEGsY
JW01Nw6ZoxqP6f29ub8zKe8wSSPH939DBVeK2a5BfAOPtFBAGQmjd1bai60u/MOeZwSDX1QmsQAm
dQZlrcqwwEAN2K8Rw0OvuPGOh7G0zfkKlOywteRR9lTeIzf//foWuO21bRIa1ARYdoZxhPnnBbNv
VOo/kw0xYF4/9+E74z9eOOrbcFb9VOFOr1hkKFjrnQ1zQhoSEHQMw8QVMz0AuHE3XuJc9Cgt3aKA
qcpuK/VBiZanxDmYgUCajFZOTGfC/8ttkw9NaZMjIUAt6HitHUxNQPr2uIeYpTbUR9NgR/bnbp00
JPdzxfmmUj3XVGRxvpzpa9CFM+mU3MazhdpQhr2B5exO1fsvmcFCR4Vk9bG+5W0IKVLgVaJmW17x
LY4CpfjLVu8DUFgaUiYoRwtEPS5B4xcCeSf0QLCvJbow/W3LGjkRJVtKSyDqrJOzIzeiOx53wXh9
xJasiWpSgTOVwDMnapSw8V5MbMnXIW2h4uI/YZPW4GFKPTNaS8SDRlaJqQzPgNqTaTy0h8ecBusb
dbppygolggdnteigCoONF3YmH4sRfTadqQ7F+FuEQ6KDNGRgqdmac01b0VeckWe+vezy/phjo1E1
id+IC2xEUK5t3zx+EFdqBZ9b+Zc4IGNRvUdSaXOTF7BFPu4e7XMHiWmnTcPbALMW2LhdQtdVwunk
2HxolldKIN5hHepIPzMdbsBpjPZfToeqm2xkxX/kCTja9SQGYxmC//Vfd07vhAT7MpRPHZYbSg3s
Q2u2CCXNorz4SsgjHJNhDj6wKXqJVNPp/VaTOywufk3lEXVexao5cIeIOUyma+BeipVElbpdgxvG
H5KAOMgCcDv1HOjbw3zG9MjgfUH4RdTYFlbqzZzLWQa+3HegsQBPeh8+RLewlWYC5lwhdogw9rjW
upIuDTT0m25a5VNGUcYfuDwlmYHUiAFZ2b3Jk02xLxwni5hNdu+NzHt3TnL1EmVfzZaGwy46WhyZ
CzrU31Rjw2XJj/N3o94FopV/SD6G+qvXZ254ZKJDYGXxbm9qbdoEkQKhBBXMAbwg1O0r9WrUdWKp
GQKpj8Q+iaGAWs/MbSh0yY3SdA4tKCSkCLkRmQ0M6Ij7EQS1jJQFV1LP4UL4t6Uez+GAunvRTja3
Q0f0RmqeXM9V67xD7DNW/ykPdYlrkrdTH6CJ8xnZieSM47JNiTo6R0dwAKKJjneNyHn/e0o8Cl2z
m5TS1knYQtt54U4sTRgOsZ3yZJ/T85OZ6HESFokr0GGeX0J5eD8mwoSRknaYJEs9tUMqsrmAIt87
NahdvrhUm6uUGCUqZ2pqVUFS82oPeNNiXcrg5aM4qxjZ9KT2wUpKESzjAkQnVppTk0As/QDpfpy2
Tkcv4ubIwiVHTkDfxzSDhVISvFFu/pscLEIm605Jxyvtj/Q18gwYddn4vLt/ydAYmpMxtxQFzw5K
fWynkbdKQNiaeu44E/rxTxj5rhWk1BtcPeVIZIM99rW5Sm8vniyO5hoSLndkhMDsPIlifaC+1Z94
PFeW+rObGQaiO/BLFOXvfjifwd0zl+uT3lvwrT2nEpIg0Pw4uJZktFepYIkijvPXgMhDxtmwvpXD
Qr05z5+whg2S0+XMB3YJdnehl4Z79NPjOOH9Q9VvhZH6QJpYCraVVicbiG9nJzoUxb7d7Zh7A6+8
PdLud97IOcHCcBxf4WEX7xKA65lggGqQu+n48btp1rLNwH4QLb1ENHvD86vPYFYSHMyJGFoTviJQ
c5IYhCAV+/UTcBCrmT90HJHYpZHcD47yYr1EIVvGyFzrFe69v2IigDMjuSmGYiyZCGLP/dmJbsvK
TLbeKugSZ6FOeM/xHZ5ZSgIqVOjEPBDPqiHLHaXfQY3BLukvquUTL9R+NF4vt1tOqn4wcltSpGHV
u5CnRn9Irg44MfrhIlWlPJ87VS51TgSvSfRcEAAMAuC/qf4yv2e1wxQwYotn1xz1Da7T8k+uN7M+
sym3ddvfGqonxRakHVr58D8+B8nIBLOK7IW4PNQeNW0Y9044RQv7R/SfR8Csyy8mo7m6sDem82dV
w8gOIG4/S/ZGsn24DK5kwPGZDJsN3hFtgnJqNr/I0rKenXHdMFVpKuoTiWcgeVnNqNJR9VEmNBTu
nC9y0CNxxGs55dN85XMIwzcANR65ydKeVI1UTz368LhT8Se8zvtGtdD7JDv7aJmoikPNdC11/uAO
uB270vKpr9c+TgFyEzZepvEQHIy4VImwlRwq/vaIa3Pm9mKwmqoASChFY8AU9rxJgoC0fo1K8v53
tYUcFDCbNh2Sl/JY5lQCRgku7srWLh2wbozWFd8yeg5rL9SO+O0rCdvTHuHztq4kh3guYKfgQ7qp
sm6+sYXW35jsAyGNS42g2jjkKi242XjQ47K53/rbUHW3FTBVh0VwowO6FPCwjxaapFcYrnRn8FDi
Q2JT5aAus15YMfBB/lHpnZuxFIA+TmwfW1HPgkUqmTK5ApDqDdES2j9IdDgOQZlqlVOXz7OxoKkL
aK1y4N8ak2cLvIqAye4K5HyHxTZPyWmtsFuLf7eN42ybyX4kkBI1PwuD7wEJAfLoItcJV0Kz167z
5Srh6HTjnQWAVkCtzBW+DyI7tbE7yTTCzZV3QF2tXGcocCke8cgzdAwHFslIithIYRTZoctnVeDe
olhgejZIeQmYHiNuX+E3bXYQ9EEw+XK9BKXoFV8uL3mZLJHvrE/G9aO7HfUjLfUwPpQOmVaWe9Kk
ryNnkFJE4GyvIaDUohuurqOqmZ3li53AsxBwx3MlI3boIn77FGHiJyU4zY6xQjYbxamEhtbqG8Je
v9xYFF7o1qt/YkYRut7LL87TymJAfGDFTj9jjXSBjWoa4dzKplxOZPoR9LlKVDALnZBLcE5HKVUp
m8nOuDkvnqq8ToBY4kLBA4Jq33juacGa2CoGpHSu0GPZM2ta8IZEDQWHsklq8OXjIe1Ad7+DbmCl
lLtK+BRltnNlj3KzMNCF2YXNRF5pz84TzbBz9m+J7MrCfQw1renEPw6rCAcFu9koDAttRFNDwHzj
WkYsN2HyhWwFu1i1jSSiLz+x58mYcDhzIRWfEOHt+B2edlHhwed/lqGFMnj8kKMUKDAuRlWtdb+y
BKBnZ3hTjnx6l4rWzFw3mRivNwIFatLKKq5361AdeEUqyZwaHL+zyvlMn8uV0sTMJzQft98cPq9g
P1SjEehyd1ttymbnOkmtDiNNFNU7GivrqSdDMykrxquokTVd1sGC59GkXo63QaCc8zXA2R/+vSP5
Bn+99ozrv5oYdYFS5wbYYwV0ejIdTEXeUPK0gJvd2MEvLrLpUrgKWjOPvs8P4q8TfBuUyckASrFH
8Mo12GKOrXyV30vo5Uh+s9H/vfuox+gazjBrQmg3IPBccXqKLwJmJSnT8yhJrbOQMFiZrxcyz437
v/svVRuP/hsvbEHHUtki/sKS01vjiEw/OrMUJ8gUIBZb/30SfwnT61c/pVWIHMvRXt9FyfFnFynC
UdMR6A8I2f8tmdNZfiotSQjC+m1To+R4XrMpTxg1KKD6Rh65IgKW87mtZL22z6gCUun//wWzGQ7t
xKkhcHxAi5fPlrDPI9w6Y+T+a9MuUjo+7Q9RLKsWlUIYBjQ5m2bUSbGSM7kgCRMopp2yZ5EU8W0Q
6Kc1u4+GzJKdwdFOPBu5VvzjYEXnT4n43iLx8369/5jd6ULvBaDkGJamg3M3BQ/xMQd5M266pk3q
geWpE6IrWpzDGxmQZm5zAOyB8/8pPsFi7EISqa1eTjVg5ELkSsAoCFvp36Wx7vrc5sKsLVfJxleN
uvQWbm06Aj68n3a25+ln/M3JxFyKIpJtT0B/3zzBCmBrTo9EO5aRdvNJWDYdAGHvOJ8hQifN8tHQ
qM37pXS2/a4So+r66LgxHjnyaF0p9KXpSYdu5DQwglBXvlGu7oRw8VqE/qKfdXITvoAFBB2eNJX+
HJFIi4Cakgx4Kdv3M4JQqfUhZRDIshkM2I7bbONy2dfPJ4aeaHCwbqEi1bcKxFwsodbAlt5ce/oR
9OIJYydKPzIe6kBjYc4yvpcqoIhBsNjE8zh6B/o2GlUKCIZYiiwXzSALjyWidPnWrY4WUMew7WtJ
QPkf778sTAioNq8aQAI74VpQSICDdb2GYEZxUcqMHNhFNBzMWybJYZXL7nl5c0C2BA0fVuilGGAI
8816sJhw65xXMSQdBfYDUSL0nkGKibWVkqCXk+Mb+koEi2GYv84QWpK4PUiczONHxkjdqAORkL+n
F/Th7rZuxUKlR7lrczAZQ22lcML4zaUdLcmT8EWw/0370pYOw/VJ+iu5u3VVVmHYhvGhhZfpiYLq
hgX0QPQNXN+jbQdv8w6dt4NW97CQnwRgPU26YuocndOqzqVGlYq0+TyTiChrH8CFc4iog/z2o5F+
xVOygZvaC153Aq5XrwNumvTPXlCs/YMqq/FkK5HHDNDhJux8YpTNsIBSJpqboh6yYQ4KInIkuZCY
aWB+Z6tqisLF5mJUaf5+jzg9FaNhruxoMBe7Lv9y5AMMf1YcBoOBC4vqB2Yy2tglyaLo7AK+t4CZ
mgH8e4snmAl5jrc57JW9juiXK1eGTJi/vow6h4m9SQi4L5qqBi5b+EaqHdlHdNPWsJsKbvjbdCou
z9JbC0DdOlYQD6nIkZ2HayT6r6fuTrKrf9WW1cJ4Pny88pYokOQUJjVnGPGp0hFKKSGNWq2Xqpr8
muh13VO1NPUSuzNnYFCxoSOVkaUvTo7qvxRw6JSqrs/XHVlw57XkqcccXFyPM/dBmPnER/DCCp68
Xmfm4o70gBo7p+yjgbZurNUyQBvpBzV/TPfelgdCIDcb69ksetm+pRkAWxp2yuJPR9fHIiw6erYC
ldoNWOCI09ll6n/k/jAB6GSlLo6nJI5lxIglEEd0Mhm78TAC6Zp9HeBSMKb8tAHyHXJnU9TYn+s1
M8CAN4eibirjs6Wdkv9vELgHEh72yNQvbENSjNNocH4z5kUsvGfDYvb/2JHCN+AbW7u0Z0p5GC//
AsjaU38W5iL/DHlnJGtOdxKTX8GOeMhbJQt0/rr1IB/tpUrV/1w2cSJwGbAUj7p1S8RNYW/iEzpS
TxWVZl1ZIUaWLwbr1yRHFzBijSz4yJa7ON5FY9KLHi1h4F98wXqaO9u1uv1ofCALJ5CVxgZ+V89T
CpsCcpxUSQpyc7Mk/Jnb1Ia7ad9KSFfYKzU5sTIlbICIev81O7iLUJlWr+xYUPnxLryyUbtCdSyw
tJ1fYxozUkVolKFXoHIi/z9MIkjKdBWS2JgQAiPQ/p+f+lIooIZM+tnV8yufptkxc3sisC4yygRY
GHBExP+gszglO+UTISIsAPIHR3nMhNf/gDSWhG5uiiUyycBJclSssxGIJV/51NC8wC2GdiOo37Bh
zUBOQaJA5akzGFqqiLsqjxmKlg/UTu5mTRcCvJ5Kxq9gsp5HhSdjmTA4NVw8FnBL5DpoUNGKpwhl
6ZeCj/to4P2yA2E6BynjcwN05eMv4PgsxMq9N94A9ZjnEjty+hqOySeTPltxXphXtxcqBJkGMugd
kV6U5UWfBQqHZv2a7bMmaShyJkOF7jcQ1ZYPchjfciRJnE1VyUnzay6iML+2RZt5+No65BmcMjzu
PtYS7AAa3JGr1UQSt3gyu50kTxOYhEH3uxim5j7A1yIfm62tLNYSnhB2ssHsU7687KnscKPw67lK
swC+I4WdutCT4ugp9W/0GlkGgET3Ptf7K9wauUp7hZa+KdrCHmGkUvkhQh55PhBjBlhZihosOXMy
441xJI/4JOM3SbxFLCoTj26EqXC/3VyRgXVAVcIH9KIprnm91LYlI7lFXuuGPqzr10d48bFS4xsn
OiWxPkAF7cv7DdOV8uh/NZO5PCLf/Zaqdy/Ix3EWUANAm9snCEVgydZgbjTpMv+AU0MEftGw5Wy5
ITB7RyZ35BA2Qd1OEgcuvTXuTB6PW9eaW818wHBGjtGtdsJCYju6fDrF7538UFgk6H4MvSsrtvUk
acD8dDg0UK5lOfWovynjhrShc+fwpaoQjxQdwceE9wFNuG6Sokt5ubWqUKBnvZ6TtuOuuoAY+pEa
vgbbX7+tE10Wx3e/e9iKNeRTFQTe+eZ9YvHjYcy2tgJULsrMlMr5oo0/VPWCvjrAhbtmBwUtkQ21
18qwdUsoOIJbRx1UtQKrQKdGiQVrPBZJKcv+5eN+IT3IXZoFU5Xyy0AQHRonBvsNJdrdfR8ucfqb
99orOq0N9mNNs46ZWv9oAeHIahbrRYmf7dpdvacgLSsQ9aZijUO3Kng3OdhAteyxXeZ0yw0wtnzr
ujZ4TczkJtXRFfiFdaVxsOs+w5TpXNE+2DcZwiVYYJsFZZdek0XYX0pXywfZFie6tJWbexieFgLN
IgHl5/WnvtgHoNXrSiBPbYtcWcvGn5Zz7CO6hVVGEJwoVVlu8asguDVEeL0UJA4gYl3hhM9YKk36
qj0wa/XoIf3hxwHnigks6vor129WKkMVFVBW+BP0YDZSV7IOBQ40hOI3lloRAJ3obLvkAaSCaDV+
j4QsjBdbqxOIfnc4KqSeqRM6zpH6kM9/QbHncFmt1OKxO5wtc8Ko6LxiarkiyDyrGwGIBJb7kxJv
IitftblMbCwp4awAjgPppTKQX0NmUsFz95i+t53jKKl6ZQejlTZtfYqcawAXs2uba8X+S5r98uwz
c8h+qAt5e9lPFK6rrb6tXBk5MUS7gQmsL1X2dVCTW1P2nwi9dhhleUVxeyhm+Zylr7TfiLnIWsw6
QuO914GYWwos3/Lmxy38ApQWSPa+86qcREJUivMQtWRNqZN1BgPLgUMk+eM8qtXxg/lPvn8rL4Rn
SRH48zRksItMDA9RnIDZDO0J6byl1rP9CcuE5BExi6jR5ldDGv/ywnd6PoQb0GPrbqeCeyEKVwG2
XbaMcGeAJ4eaOv39hHpFSaCSjmY7XGZG7DC/mNudFW55fz/OeCFBkN1wblrUgCzwTu+Nxk16A/CE
8b2WsHCoPBk/oOIwYLSupt7jnFZZo95KSuHU4cK79jLL0hLzkQ/aDliFdlJGTYFiqfm+qyt+WQ4h
5p7WdnY2zqYxo/F7yIgeTcihdq39z9WIfD/Acec8Mw8NeLgV4bEOvmsyb9Ia6wdGiJ2DkAfA9M3s
xBDXI1fw0z8ytkUSFkPUunNaU24IyQ483yqEcPZKCK26J6n4y0EIrrcmTfSfLRT3Dna0z+238LnR
r2xQQcjAkdcXE4tIlncuWFYy558bhBB/wA4j3aQeBIISu36qXTYLlT12ZVcmpPSGiTx2XBV7MR9w
LIp1SJD/Q+fHaQ0s+1c5z2JjKEdj3Bc1dlL84DERmfvzew/Q8J8MNtOT8+DrNsE9alMulPJyZtvy
kFO3YFHrMR5DkZ0/YNByV1iQQCZzHNN9NEe9AiD66wzjtqPzP9HgmVkwRjWjvs8zvJLpKjKRqN09
Ftv/edUZiUArRjk/gSth96vFDKTptDXOM03F2Eu5M749/8SWIRL8Z5atjrrnHy+KoAFpda8e0+C9
3P4NLI5LL3KgxFHweRbYYeGkPNY5exzOwCz5uiJno/iKHreyvwCX684K465GNZgEBqNATBM2K1Ux
9SAoOnA02L3eDK9nDPrPGhnEQNRt+ztsHfM68aNWDBTB2lUe9bIABWbkc7Sgs5RJ2ti44gtFsG6q
6yxRYyvhwP5j29k8eWdqJdzRyG0qWrOW8eS6SfDb3+P7ni/UlseItV9rlFQrphiM2bJtFfVedTGp
rC8tX75/fMudBD2k60OoTKHpj8fQY7+WE6xhZQ41vkfstHRakmtd0jPCjfNpWulwq9jJZQ/j6EA9
8u3N43AnLFTwyp4Vbx/ndiCc+6i4s5Jk7tEeqRpMZwa7gHFLvZflmtg2nu7gaIJwLdnMdYxxIz1A
jkMiKz3vtgtu+On3r5Q7KN3DUoyZOBua8/arL8aobzxtuDrlyrGFAv3GwbxeO77XJSHjWzrcX7Mq
SfEf5g8594R/mwDFHqrX6ZFoawLUvpwInq3470eMEkR8vNX0K+Vo/YPiKfOE6p9/tAqJnBp6t5mn
DhdyfbjhZZE4ITddb4xSGMoiVG6sT5f/bbkVYu7P3iTvbQiCcTpI4tUOJdRiClcxx2ibBuBs1zhi
WsTfpqaWPBBNbIGbepx2eDuKo8ugmipX1WtmpkCOtk6f9+f259heOo4Pcp2UO44XGR6RLX7Z9GUU
dH8WtKZXfGSy87a14CY8L/VEyfTy6f1MYHMG3AJ4ft9eCkrXq+M/mJZbuo3ZjrQc1PN/lQQFDEor
mi9pLNM0YBf/WGxrS8OPbCc0JipRq2QCFedJLBmc4bjsTRD4fuWt1xbu0uarnbyXKxlMAiKmKMI8
XXz0McHol+oqEqF6JmTZu0NKnD7rHG/BfBq8sdkbb3nukVE86LWK27BAXjrmthJl4/N0FiAPDcO/
fMVRcXRmiVv2YHxVI+Zyad3D6yJUpNpZbsw/2q6h7jfG9Jt4WX2S2W5QqaLpI9kl8lO3280SR1oS
wDNC2T2XeNzj58rvRfQs+Nn3uK2+pbxKDG/cw0hzLpQNmrVWD1HRWJ4j5do3hZILwY03Gxy7C/28
Iv5W3L7o/zX8++GkPSSXfaq8+4cykVwplNFiLzhOqWhflSKkNLvXxPwhZTmINicdQQgH/ijzA92U
icfjBJqEVLJ76q8NE6HwZtVGC8wihFgroTq0wEckyNOXi+uo9nOV+rLCGyCdZjMu0f+09VF9SezY
uR8CcgDAmhHNcnA/rA3S0vmmIB8r+qfERXK3bZuDnUoU5ab5HHAtH5IiGbOysyKYUaGZ6EPF4kNF
QCpyjc0db/5xbfqdxwvLbiITwcHMNUVEZmjf7P5IjhcdwQ0iLnZSvxLNiXGFnBYTu08T77CkzmbK
fsVvyFvV0TMBuolA2qGGeF0Vi9xR2cd7q4LAAPqfof6X+tyH3jjzEU8FXJDkmaNfbnJQQyeieb3p
loxgiOkYdNO4mtCKaBWBcj3qnHUxh6n37UhcyzS02Po/OD4DjFuQbK6+V5/2jBL73oQKF0lNOF+4
0b1po38dlUAEsnfn9QzVTXd6DVy2L0v2azG5vCdjGHw5IUWVmbNMDx0jiKnmJeDKd9KQCeT1oWIF
LmnuIv4klHsM8QCk7PI7pBjq0DRaS9PWCIcNK37U9dK7w5TPRVU42FIP6FBg+lOqATOOBaKJHph2
94ujeIV0IDnHWW/ukWHQU/bu6TAoFipLMPWhWjslaokp9YWXZHqs1X0VWA3rOGTFIB30rR0eXPmI
ceu+h0A38Z6iKVPJNwPifxKNlvUe/YQNsy8xrLPoGIzGNtcnvg7mnPEpGG+dK4jNQZeAZLYCwz0W
xU/gvtxDUvGITQia8CcBnUS58MvYm5fcYiMGXuHb7BNI6hVNeK7VtGpMv27vDgK9OYXWi7nbRTXK
MI4lM/NSBKW0lAAl6Ab35Uc/5s9Ob8xB+GhnNCMSw+TkMAA0dqx+/bvXr87moAh2Vy/4RYFU9L/D
DcvkCgyMp/qc1mt7nEDAFaCJn+gzxiuDAgfMtLrRSjs/6ClnowwIoDQiUgE/4kS0fiCwE930x//K
RBXhTMhPO+8vO/7ugyWvCghSwy3DRszzLfP76NQoXGrDkfcN9fvHBN1nd0NUBqgS3pIt+h2H/IaQ
eaH1odPqOu5HapxBGXar3UP1THSUDKdia+vq8M7JcGHidAxUdocz9+F7Jwx9JUXnggHYIIYN8ScH
YBTb/lOMXfkSK4XJgsCrLHssHV6GYs2fuEhpC0MHI6zp8NdqLiYPnccXO+A8ASe6PezH5rCydvw8
4Th7npKUfvTnu2IyML4VUMba3SakOAD1f34HFIfNgONtv/h7tIkiD2Fyn3IZktmEIJnVDICLCuFp
J0EuNLIAv6f6O0XKpLKsFjb7mhCzxtZjvxTkPNzGVAVFwFAxdMm3x6W+KsNpTQ8oAOBQmUQlJO19
E5Q/NMEUCZfIimaPF5Z9LKwwl9zhCEJwVSF6S6Bhhh47O+eiFZXASCjGJYvQcicdppvnn1OjgXoi
rDcx5RN/Qw5aASJ2PLDmHljnDzVqq5yAXoHxl7iaWte1DgUWyzRxDmQg7CHpYsGpp2Hw6Z7REvLV
VE4MWqBHlS0uja7ye+SPa4wMftG7V1ZJ72EtwdMdxHIyLRd2NbJijm0MmRePU1/hhmAf+ltMnrUX
DJz0zgjaw/Y2MqjAvJWP6H4PZhShGeuXyp3txvxvmnzMd9+4VJEIAvwq9Dt6IMisTDl+JDRRmb2c
5rc4C7uuBxJ8DfNPglLvShiXmHNU4ry2L61dH6JTEaotHMFRPLYpEAMyzDO4nEFviCzb1mg/dYWc
2DUaECwEBRROfAvkmagMWrpTjXw6bnXP16OC/VRJRtnlr4jgD3lh/sf4UuwKhtJ8wmUHvdxoxw5M
WhnjXIM+W0CRmpFGnhlnvXDx1uoRohGATo/bP1TyF0rdttyswjeDZFhnILYtdSUurY1qWPNDl1QE
ufzjmY/FSklY11PDCbQw0oUi/ssEKNIr9Zr5T7GAWM67XVQNtQl72fjjzraWXlDUqmm6/SOlgkQe
z6DorfSJt4PWQF0tQOibYg/OX+An6ieRfOHKHdMdw42+YPXm8FpJkwQl2hta1W+r1s+HIHhTCI2K
6kS8RrETNxRb9rIPloKzj8IbF9OOGhlujWb6qjkFlEo1SfPsPhfGcIWhiuCRgHyYbiZgVpNJk/Rm
ydewrWFjrQHxj6kYDE0B7cJb8BmVx42RjBO8gaR4DpSQsJiGeQ/me7GGpP773NgEbk+WhU3VdrP6
SEGWU06JKcN+XYZrwqn7Q2UA9Q1AGoyQqqTFHgGxnGcpOK6x5/B20tb6O2YzmpZtr3twcAqJz5dG
bxF8Q73EDv91yYIaHZC3oX17ECD7Vv/wQBjtlKTJy2tAUnD9zmr0sY/QOglzTTQE/pJGGimKGQEN
zDhvbLBqw4lTkBWg12OHmyXjIzo0payzwWI2DhsKIaThuK7SwPFZRmr8IryTsfzoIyx0uVI6HeCr
4XhigIhgHNefxV7daeQIJplwvS25IpJMpJA1V0CtOVOc2Pa73U5Zf2dLF7EmtEciv6ubBu09B7FV
U+NW9W/nHeGEH/DPZAXwOr5VUZwP85PTa480fGkRoAffhJm6Uf9L3sPKfwonfZ8ndg/3O3KG+LR7
enIRMdllmZzliT6jQLkEkjdQhgSLnXhlA0e9CPWb1mGKxVD/Eb6Qe0XdjgvgH+8z0whWqqZJOv3n
ZkdugdqMDMaw4TNpte+Q/IUCpCsZmLyxDaYyVcNokA1P3Qfn3GdGRPHeP4QUWFVfDrbXlClB3LQP
4/s8DqQmMdnUI0vuAmvlFe7cfOg28dz8zFo2PNhpebrCoFvPd+gR0ZdXww4hHOOlTsT1gH7a+jUM
NVNiscE/qcXr3ibNoZK/GFsOKU78qBwryGkSiCb+W+PCnnsMJAJIRG1XY2g0bb11PtCyRNGPj+lc
1BXFeeXIdutzsQB9mfjUiwtTTi99keONU26AKILiDaMtgWHcNz8zDzHVKDGvfJHxDaJ4yaldXfnw
I3naVekbf8F9PYDTTl4Uupc1BpVBGZ0/RMvb97qDF6yX6MOABjG0sTUfDIsm+ojf5CKF+NujeI//
4fM+cRyQoCQWLZOAaGS2lueMVkA7qfvxJ9+rey40LQz1jOAoHZFJG8MbSePBIb5vn3IxHyJYEONo
s/ThTuxZz6SHZKiJOEQUzWO6jnMj4Be6rORtw6Kvm6+2jE0ubexQx0Yy5QYBJUnEUq/6btkRdaOe
c7VaZenu7h8gh5Z8Ifnzm1ccjN4a/vQEnhQtDjmlRhNkyqyOfEZg7A+E3SJTWaEIbybykSSS9t85
GM9kvMndMLrGbXfpfGYRFCxzsvJ8lMBu4e4MzoCgF6d3KP48If4p1eGUKuU0v25W8F+DHEz542BF
BVfo4bTyPecIetdtVTIZ4GclK4RbJBdV7bZ9JvgFzUoSf5Z9KDdaKzYbFIk1RQv4O8NXLgd2TBAu
OVOwL3oxm2W5gE7kJF0ltOdKrGR+w8XXXfvfeBrIUGBmQqk8HxTnGkBBEUtK793wXSdu5gpGUUgW
vTVoeQ5QrXfJ+xwkmBe9hbVjt5fV3rkjpRgLTgulIbYAHn7KoXNMH0JIHlglwfvw4AGPsyzVLP8V
T8YPGhSEL64cHKl+4nz2ybFJAOKIKFhjxAUB5k2QTw99uKi1hTf6B+aWfnP4c1KypyzZEtziHB7I
Ap5T2P7pK1zQ1ZC9z65Qwcl+INuBkl8a64JOl27l9Oh2xknbRd2JC9LWMLMfzfkZZ5utJgrqp+kK
xE5rn27qS9d8m46b/HKIcGhyns6hhvpvHCeTdDfpHdDqb7eWiJwy0kOvuaMsA37CmyffavZd0lZC
B7b8E19zxsKVPjP9kFMawNffo+xj8ngO/sU0VW9x5y9okLycg+UZSBfOvAfw8KGU5vRgUrtp0Y0S
l60KLKV3fdbTmNT4zIQxiPUpkTAtPh5k/OEhPWDGIOp4Qts8fxdRctcN6mm7KLDBaPxRHi2D1363
KHNuPE+WEqlQMTLJ5EVTDr5j/bBoKRj5MlJetuNTamh7PEHfZONHsZQuIMT2m/oznUywwepxOpEG
g93oQli2EX+EjNoi3kAjcQTAhdjnvHInMB1gvAvb3RuqLX3BrR930xDKdNwj6M4iFpv70nXG9Oq1
BEb+nRULGfFZnYjBhXvaUfa4gqjAzTrijg9aFda3zqZE8Z84jvgMQmcRhcQRKK+4o3VI5gigQhrj
bVSpqakOPe/JIA7WpE/8XG6+3fy8y2XsVZ0xhrEMSdtldit6cuf1jQrueg/6nH/9EsVbU4cnRKN3
Hod5VTaZITcIQ93G3e/KR69bloiLW0NcrSmMWPzq6GJpTdC2BtJvNe0ZLCkQC0AOvSL6zISxy2lD
j8Qs809TcFHYLFO2XcqN2qFUNISXtlvKbZgqyJ0Q/yXcTYzOJxRHsR4p2E59m6jEb/exHZvnSKSy
PgsYsLU5VBsu1VJz3rp2HIfu9kMsUi9T/WTpc5zTzkUITzXDAGKet7OffDMO0bZwFndaLTZKo2yv
Nuq6ii78R8zq1bYccFXTvtRM3ki0bhAWp1ePOUp9gNCUv3tNOOfSG2+5Z/iBxRhPclqnCO7Au3c7
ceURAfFDwPJgEyykE1msv/7LzsHdwLf30/BuRMNEiBj7QAGT0TPN3LQKCVJBl1GcldqeBx5dWIzB
IP1VuO8jAlUGUHH/9fPIkgkfWbQUOdUUHD/2mChnfhDiiPOqDIOeKTRpJNeX0VBPnjO9jemsBQYb
U9lMR/xR7V+m9iIS6GdZckNWVrViRyPoM5LGEOawvjRHSlck+dJUpMJfAzb+VH+hj3v2se/pydcn
rQAf3mmG5pmzR8tyYMEwMKpfOCwegezC6aQe1qtqGD6xAMEGrVal4TjTUR90fyeeNqt9XiKa5F7Z
sw6UTgbJ1DBgi0plyUkxeGcBL8UfRb+xFPJDeOHT3l+dPR1XJKGoZzAGYfPSAJ4T9uShl5O6fDob
AwIrcJtIaZIuSgQ88JujkptjKKbqSCbOTH/L44p+OydsmBRNWRTklvutCywWnLVIaYuR+pJhfDZM
MpygF/roTYd8+Lo5/oWd3B3lnYqet83h5aQ3kcYQh46/q0hHmhwXPNfrWqkn+GL3RzNlsAUGhwVK
Er63dLlQ+8xrY/s7LF8H5sHSp7n7jYZeeC/dzG+l6835EWGPERQvaeQw6iIvqU6vq5Jwhns5RdG7
XelCKOV/JzOX2A/to4MpYV3bq2s3IjYO7hGaXmLZBkOnvnvpUfXpF72ansAYben4WG3LgF8VY823
tLV3vjOEBy6+wBSYGeQ8Yh/lNGsEpmxYR3xX8DVoKCPH4lDbE0W2Yz6qY4waA3BoWs0i0R9nf9So
rX7CuOYXGtZW5nlYZvwaj6gywQ9mRHgeReR9bKLlrqrZLJpbDHTRO4BNgByEwrqA8EfjdIZXFXQS
RdsDxM3AKJEcqnBQ/T85iIGqUzQL6JgtXyv/PhPzf13ZmEFdfT4rGpot2MyOMKzwZB7LJslOQFW8
jtPY2APy0ZzLf8o7S7Bhd9dN8jDvH4haqyV4qVbslqF89QYH8V6dU4O5hO4PAs8t2SLzExjAg4rc
wWSCMZF56eGzmlOVcK6kZFZBoNweJSwLVnlGllXHUHgeXZSnp0BbTePUPOus8acMMd+J+Gc9BA1j
oVAlbJVSo/DVxtIiXRcTqJe/cAbRgvBo/Ty/Vlgi+4aG3R87mz6NsKQ8uwjUsMGG7j0BzGgMTRlg
zU5HfeSty3I/xC/il1dxmTind5VAL/8tgrMIFJVWwWrlVGkv9QPjdjJTzcC0d/JqCb6olpdCGScy
RDBLxwKJWLx1DUjmlFqC28avrj3Z+1YJuS97TNJwJizGMpoLkJjK2I6lv6j5qA5Xts0ZnOqKxlEo
mxBGK/b9VWQ7xqjaQtqmAtHMzi7LK4icEmVeCcj41YThq3JdhUSqu0uOTjS0RSvDqyZ81wLM9vnH
biRAYJRzrUSMObazXHykMFQmkKspCYJdDLa7D02FmKI0rmxDVLDaqZD7rHUQdodgP7Nu1CSB51e9
RZ9HdaU7WyWRH6R8Tcbcfn/2XcZf85+oG/kFYiu6Um0yDqQ/uHoYqfmOcAR+A9y8pWsNVJlkEXqm
3ChFDBtPCtwn966WCMbX/r6z3k5xwJpbhN7n1BViPGnDpuzywSWEHnMWYgiugpvsneHqyziBPxvw
2bmn72S7e6tXgYSkL5mpYnvZUNTF/xmIbTc1KfYkpSMqGUsxGibmPKNA5ahppKhSjr61xTCGUydX
8pURDouGdewGCWUx9z7L3krKKqwjC/Z3OsiPlC69l3/9OtLDsxVg/UZ/IfQe5U75tIGgq9U94sgP
Af5an3Xwh+qp/z6O3jFJzn6hMoLiUHks7AiB/Z26+BvTe0meaNYhQ1PIsfROsAcOee640vfPzFI5
aTX7XJ5ZixPRtiGVpOefJ7yvHUls4T0V6OM3PTZ2rEqJkSQemsmw5GXTm+hvh5/s3EywEpKCyRS1
RvJ4QgHdLqtVIGjb+usNztmwh/KDuLM2b6SftUHlZREueBOxoz1HUJ/F8mZKgpsgpFNdvaVCvOA2
WqsDTe/yLTZJqhqMuFQjpH3AI/cxbw4Ex1ZHFvnmcdGaEjtHfX/gFRS1RMXukM7QgK3kQND34O5Y
U+bFELKDzkrjphkg6WtAJFz/GKbyPvZKUg8jI0D75QqSdbuttQbT0JZRh1NtmQkML8LeHW6+mwP7
tHXPqwutETx8kFPlB03pjy9O60+6z/9ObAjttORSfmpQe+EgE+Vw0DZyhNA+Xrr1r4tcTrAUGlRt
BlpNw5fLo/MqoMBZ39VAxhImmpuOdsWAteBJHP6rwldtoWc+3VbF0GJotibFwQtWG3wsZW8nWOCf
byRvqp2sVsdVFUZgdQp8Apb01aMNWjokPM4GIyCAe5lCxlXzqHLlolfVCcYF0I3+ZWpH4fbXUMVK
7Fxp/Muf8kBYZR0BTsclGIWsqz4fHvSSIUNmoS87/QKkJFsdxzfTArp/Y9oDxCnpGbh4zNcbtmbG
vJURYq0wCFHjg/w+AYEtk9qNqHG8WgjLVC0d14VSQZa8jEbZvyR/tGFRbiT+FinMeoAQtzWSd0bx
RH1Eqvqpyo+bLszH+AQqsLCC/IrnZ+TfbtpoLbJC3XbXl5I5iJe/dotBD7OBJ32WioEda9qZkdSn
R4+0Uf4482A/2kdR+f4yEZzKGAcqb3zRLCOdIdOO9jLOY1mxwiVcFsAHRcs3h7raRoC84yjgkkJJ
l60DoUvFyO7asLzrAawzvJfm15H30zifwwUJlXyKNTIJqBFnBeHz386PzSQsp+oAh3/pdYsX+gTP
I29dxJ+IrxRfaimf/fLWYqox4ycMF6VZAQTT/VuFLx9t0EG2ndmawSz0Ur/uHkrZmu5+Zb2lc3si
hPzPw7ElA1r4AN0C7dEchQ/zi2DFVEfQSOe9fVFFVeMlDHKRYFSVn18SaIcoWrjtTv7sPTmO0k4n
MUREvidSQ9Tz70yTjEehgV2QG/dH/Dm9UKs0Z8jNcBy3Lamj5rjj9FtSYoIlhKHKFV0B6OLAbX9C
7P6GF2cmmbjFJwyoCfxCzjqzQfGK1s5b4uaqgfLVm/kL+WMCoDI7uVUU5oLi5FhznK8aQyEfu/Z/
dJZ9T9fWlg/ul2ciEuDEUxHYqp7rnqzHRYRZPcFKNdQb9Td9UV20KF+8DjkEecgcrc80rD3W4uby
Nyil/XD219uX0iq3+TYuqaBZ0Q0Zc5+w/Hb2dkEax0xCnEXRyzir5rM6o8lExKZsIQ3zSVbov7Ck
ePNePRkaFwlJo+rL9eJWS0DoTbrQSB8oxqO3LJY8t5Fn3mriZ6OYim3k6GCI72ii/2d1tAUoqChN
JKynXyTw/Ote2JZyIFpnzM9Vz823De8vfDCw3c6iYmpnBtH4bt7vX6UtxqI+JnDrmgwP3+tjwT2T
J8FfMpbQQHXq+a8iMmQ1Uw5J3vbtHt/VzyYD8AwjmwrxPiH8+BCT7Nu3jq636SI5jlK2Sl0+rWVu
FvD2VucnlfC3t80JkR8BpQvVQOXmcwgZcBOV8lI52AilOU3dlXpqNMyn8yhFHtQU+LIDVh3sExuT
l+1l1daHob8mBNPPYWIDALA4kS7gqHqQ2JQdJF+0ghr9lQZYqkvTgBnna8QlY0LlwPBeSXH2vnCb
JMr2TvqYTFWTR6ooZu2NWgmLyfZFTgm5xVsIH0qvl7gO/YWuTOOl5Kt3W9dJiWHlqUbYcpNw5sII
aTVICghsPkBWb9KNWMixPB+ju0MQjYSLIfCuyIrlCt2iybPqAtpb4PUTBi8vxUuWlfflFdXVj4gg
XrgK0jVHtKjAwEmL0x08ff8QN9qM86bPOleokCcqHwZzap86qSkX5MykAq5DXtPEp9a078Zw8I1F
84pbo2tlxPm8WqDxsoFhz5FzI7V3QombipwetybTaQp7C/E3ywZJQifGkPpIT6ckD1nXj2tDoyHE
8x+YcyyP6p/3ZH8/F73GuvVSk0Pgq7aq7FtS3hTa6qz8ck1afRzwVQzR40MlClz5WJMub4DRirGQ
Hvd6vLE91phduOFfB6jRfSncqh7YgtS8QpJNoA+DLLAsd6PVrgXU8k+IJyc4Ryd/IZjVAeDuK9i2
9y3jCayMNb9HVwkn8v62+sGXvHnINevGyK8YLdGl/kcqfVIzKomjTTL/6c2G+mfcuhwXhjnkBZTg
MufkGNsoQ51+xf1qSYuo7ESTMCd7/+o+Hlf+rsRM49I/ky8w6dnv1r/VblABO/p8/88Swkn8W2NW
goaAVxAVMKG2AVAg81vhHYBmgkviJqqlVdiQWxxAfRwtBDp4W7KacqmakEPB+e9BhM5mULr+vUqR
QP9/1UDZaEHFXRZHrZ33IHpA8Zz53u6qQzMCPnd4Vc5gd7JUMfIhD6RVUNzTc36dkoItYpfhSBo7
tq8E+9w2S3KjmsVnqqWPebcuA7CawT3EUAdOPDQDdAYA6PxWwAvKhwquQGyN07AUb0IledKb8gKm
DMVlQKnQNmrn1/6cW5P6J1V1OOWmkoJSEnGIaSg2P2TVvoUr7haeqHmUxczO/nDwrRxg9akzysXq
w2NPKQA5/F4OBgyWexaRIysu6KpYXPhIkHYNclWPGqkc8T51AMegO2hiW2g3u7voSOZzdAmHKXbi
8ah2sio+8lIYhPcm66ZYNXpYfBLJujyTd8QtvB3egjmoGbYXI8OlaVaKJsi4V/BoGP5CjwLVWHNI
b5Sp29P1N8vNojrnbPeX2Gj+VJrD2jXwBwkl9q9bXQsOQw4f095fNdHoajFeCwbC4NGU1auQlG5t
b4NRlE6VqcZvI1aefVOZvIs7pqPvXOXO062+U/7oBcXcq1atrHmsyMTj1GwgXfvDVXbeCgxVoA0k
kZ8Dn4YyFMcCSPfjXle5q0ZBGYYLqsDmpAqMEMjb3NxxSNybewTFeikQNPofcDymuLwv3RYuvB3L
xLG5Z9jSfHT5MRv3Ezf6loHB1IzL3+nwGuawvisjdII7OaW3u7/AGhAUNQsvhDxfb2qzCD9j+icX
ZuyjWdsNAykM3epKuAGSt/NhtMlyHCtQ/n3hYr/mrIMHV3EyTeObc73CWIhOTty2Cu4T6PljQgm9
1F3bi8yhT8Vc+ofLqP0iCkUWJ6VqTi7U1Tomy+GO4sqdocGLV0COl+Gp+xj79A0rN/zaJpNjyFei
RwAn5LGNka0VJM0W3zDTEh9LGpatNmoPOlaG5NFMpiIMS46amf9559oSyKD/9wQmxlzv6igmwhfR
EF6352DF1F8Z1jYGnIg8sd0roBgkBSQEkgu40LWGOQw2R+fICEYtEs070xOJ7rTuGBXBXk0EAl/2
3FcHTYbP5fZi/RYCmQSl6JFRWIs1Aqu36UB/pY7uXGNLZ+2Ai8HfqBDr605XAMUl80WK2py61l3X
z1Oxnzeq12jYZ3w4VSns9pLfpewncVB3i4v3ldJCZA+usg+nbGeaXgPYBhuLJXaxpypAVOteQRu1
gDyywPTu2dJkYUMgwmvNSgA5bwh9WwPg/U9Xjx6ASxIkShiBbgXryN+anp5lM7cz6d6SA180soXn
Fxke8tBzkyuueJzi6ZLZgoLe5JTNSfBTRkDRtCcsXwqAIK3OtRejRVt1Fvoy/8sUMm6l6/eFn0wy
2ul0xyRGzSY0lMj2xa0XzaSnmRJ1IQMkKYZMFWp4gR6PkfrqHIcHwwmLp/fhb//B0RTxVHgOdl8j
Dxofl3utJBx9Xr7o8ZZQr/Zwt16ef2Nq2suKEXIwO/9NAFLrRUCAlH19RYNSeSAn4VxKEb9XyZvh
VFOvZP9/A+Ei8jojAlOQ+XpVPe+vUyc7Tc1kjfsJ5EtGOoATjd9mTbhIapdzwTOMcgm68dZWWf5k
QXt8rqD1VQ4d4W9DHf7gpjDAPpLLk1ZZx0YoTaEHJ0m+W1J7gjQw0XbxSrWzpMsMprleDGzktMGz
b4vSCfs4G1qmZjwUgfTaajhHDC8KqVVj0x669yaI02+hsJOACRgFlLa35Jjl9y3EFwQx8hU76mvu
igASK9oFQZGhbM8Bb33w3Woyme0z4faANzr3xUgBWJRvdr9x89YL9X7Jt678pO8N4qVwImd4LJ/x
x8mK2xN6csfcu/K9WUIutuSbHKKftCCXsSIWSjGMGdWljqvsXnQu1T7jN1vH5rCfThdxoREGN91X
DusiutztB6Ro1OM9udaZxSV/6Xy+pprOWwdIzuT897p9CPwk4tXAt+x9Ebv6VQAvbKLIQ3kULnTf
49/fRqbSGoozyD2UAnr/jbmFVNYbEOtFMvdWVtq0RDgc9nkWsd4ZuxcKEgVIAyYOneAixFEKhEkp
3sujy3tPKp6uXU6eSq1uqzJCKR9QS7CaHDtY9+KSwFAZl1MRwY2U8aggOQhjm1j3X6sjybYKok6N
lWj6rHpT5nqUG+tlBztA10jF1HRYaUSMFVbgemGWozOA1WYUZFudYUVLImWKcC/uoNraXVTtSc+V
sjcjbqzZd3I0fMsM6De+4BshL2CEzsjS1shqo8nylcvpaoWvTvyUoMOhaNXUAgtTgWGL25uFbQlZ
gAOKRz9LltGKLzFDG1gB4PHpSmtC3is8SPgLXVYV5XIgX3NKBNgAduTb0ae1677BelSUkgo3Mlsy
xgCIAN3mYU5MTDHe87tbW+Wd19koSBWiL1T1lw9X2F+yQVvmpfm8XhsOrS5CO21xO925VmZ3HlFQ
ZmoPJRbYspCaqWCiiwc5aGYYb/ZvXr6CxWGQ/e54Ye/6cNKy9CKFOB0WkTEPb0rdhF66nZBPtkUE
wX35yzH1MGHDQFcfIodOepMzTwuXSbMz9u0BElET9jbx8I+M306fzgUu8vAIe8NJUNPTiTbCQsCb
efh123ZU6UeoYnp1sHoEC7AgC/2ogC/KuDWvYt8O5aNDSrZKeca5TEZMVCX0sKn/pQyVV48VhvPH
C1I5v3hG8v4Bgz6gzrZzhnLjUGuP2ZQlTCdmiUi7TY1xLytKVPMX9ak9wcHQ/wMyuus794tDkaaA
L9a3sw08RwbdJzWESCcjHhubKb8xzN56C90/EyKWHMsXZwkUTeX6DDpsEwWbCuAJrcRejh3uhj34
S7cY03pzsbteUbkx12WOnONsdwpjcEJUDHUDhmhomgxoWgcaYU3wUHCemIIhhIJisUpHNiwqLs5s
UyakZOa42oTG+tKikZbR0p9Y5igpvGEzcgW9UTx4A+rIsndFG+5bGhN2j3Ytt7RP2HXvVLqIuKJQ
QpMARIZI2mWhm13MhWAZTqOsGCbsrFZyobo82IQd21GdkPFjoJ6VkuzFDVjxT1iLvJrqSCLTvZta
d1HqH/EAvrPvAAibfVviRP7FMvvcycfPNI0DCPFqaPxJ9OWic3VwlkipYLJKH7ZlxT6ZRgQgkt74
axTLZ4autyBEsM7UUTzAC6hMvynAnDq95S+tnMtNPlBWrFPXMk3mr9MJjYhn16kJ9u1y1qkmWMH9
DaZw2CmtmFF5BeLpCg+GKLtCrXAMK8OdB1MmuF1JicuXUWpy1jPC6CqIRdpjuYN9YB1XTFhzDR59
bROWJrpQIMgJau26qIMqOty6pT6cI7sSwHwO1w2vIAdT8d67RYy7FFROvpFtPB4bGeB21qUHwAf7
q2H5fTbumZrvsWER2yz8A18V8kOeE+Ad1gEjcCc+wAWmszVLE5O5WpKm9e2KWVKM3vFN3udu42Xv
MlHIp+HsOJ8N+o4lC72I5oPx37n3akhgVHiC7r1hOmiTL/TLAITE/gkLv11whPb+E3t9exVK4oYE
u/kyD8VKQCfg5TyE0BH37d+rTEUZp+kabjS3JGm5IFu1sAfsAqF7TJz7wAKnQ6clZiNkGqt+Ivmb
LZvvi/Zex1CEr6nJJtk3zDW1HgK7HDMO6MOs/V7l+wIjInPxd0ejqOijBfDfpXvNuV9z45g+8k4b
M/dxpt6NsWPsGS/rGVtJWroWy5TaSg2D996+P7y4iMDUvJzUIKUx7yopl+XLkVO6VOnsaKhjrUA2
Pssrvb9537KEM12xwt0arqMweFM2NzVc8Fa6Nbx3LyQKxHCGPNwJ1GIPESkwAqrIPmja6E82WcHV
IQGdr97ghnUyX5iXznluRWK1k67EJz9mpnHZffcv3C2ypL41Q0+oZBVvs+s2HbEWRKRrZja0EY+a
w3MLY9+vD5RIBJVzNJXU24B9SEtj1NALsA8e3idCj5vYd6oAIs2C9Iu02dgG4p1LlkNpMkAWx3XT
I+D7NCbS+mhiodgtzuQRPMg+YWNpv4rc5ZpCRGs98FxMJKvzuyw7xB+zhy33A+YkL2FpqE7SK+qq
My4ieyJPCimpMHq2eJjbEQKo6jW8r/Tgu4bSmkwZB3L9qNtsCFu4E/3nwTQGJXAwzjLSnx8cp+oj
xgvQe7xNoIwj0FOziLS5AB7DRzF7LgE+mmxxHUdW+sSfq2L805thxykYDoPti+xTMiXCm2llAZ2K
sgJqzbtGRklbZGoIMJvcUHdYmHgbU5om9Yt6KyZkLB79D4rA2g9skMx9fo+H4G+yQHLsMYvRtlTU
EGjt6l86idWhQcM574nLES4KMVB+AfNYnmsr3uXSEdIj+rpc8X/lcxSIDPtsBDv6jXJnSRjbsNB3
fn6M8QxLVuSCrxq1XHreDYNKMc8P8v+VUyuHJaqwnqwLPSKQxgeB8VITXzNxWypupDDCv8xwhgSY
+AeZfYUlc6E8PA7k97V7suwi5ZHAzcM6/CWNHRte8pAC1jQu0tbJnTrn1R1gnIJ804QCeYcjeFK6
zg1T5pDFteZo6plKTFpgeNj8TOiiXrsKFFYUi29iNFKcfv5F+yHd0CDUtFJ/DmJqxJXo8sJnJM0r
gbmM7OXmG7P9SF7fLB8Xd7Er483bx+k2i7T8GjUZvOA0UIV5gY/E03WFgxosEEIqMWQ+2ZVxCbay
w+457UTi15gzX1B9ee7zZEGYJI9SmszVUYqqTS4+nOjBZqPG7J0Q4X+7nGXbltpPeCz9C4bjiYWe
KUAQkpG/og5d/p/5Gk37ylcrpOEIQyKUfpTHtDr9hq0PcvJiq6HVvvrzPitVeVh5vx40ZWXkztBc
X2m/i0Au7hSzemzOQvu/Zm7ox28jl7MAxJ1TYliPLfwLl3PJmih+ipCwgh93Bjk1r0+hFIPzDVzd
G/ys/MQprPMI8LhmGyNtmiEDhEkam7tMq8i0w9t2cwp41GhVtnjxTZxMlBkUGEYn04gGJXCkyDJX
6fSrWuTeiNLqk5QEA0G4dDQjagwiNDvw1Ogqjd0FXMSPiRWGNLJlfiB0ux0m903q1ut3y6L3iQUO
MUifbmOELJ32/02+2/4FTEGy8KD7nM40QPHRQogOxbQIIkGYFLNc7/MYrqdzBR5BJFKa96SMyRQc
iciDsQZfN+Pl9IkHsHoK8DEC7gQ565C3ZwmAxEQXRSEtxowk91ikPagqBBL9/f71Zf21E9x3UNAy
C03saWEIaDI7JKAQGWCek9WyWA+XojmLyW+j903yweYYn1ZTiQ0QD821Q2t0XQJM032rjPQy4N0i
vQxalHcJznQoVT7HbkQxrvsMlrgpqGUp+k+wLBB51qL+2wNxbl/gS8QdeKpq2PBgMVkbV1H9PZ1i
D1V35AwTCGt8LuOJDaeG+llNLHiTFnkZNqRkNT9OYHSnz/7l0Ev6W2qt3EAVS7ZgmKY1bTO/nR5S
0KhM6yXKNrlM6n8aXY2UC5TmetwnojRJJ+xB6VnbALe02CPZL4xJ9c8KSYvLas1Z/JPcY3KwcaWa
GbCIEUp0FhZeL/F/86wqqrC2d4W/v7a435lmBqmlJKEMK0tOp/MOwTr5IeB8yOWRXln2Qgir3D0A
3amo09bX/NkaXg6NvfzTJv3lepqFVCv4FFzFildW8jjcOw3SXxHSZ7UyxGtrAGQrIPQtPeFJZ50Q
UDD7tOxJclnguMN0PNOS42YjqDjQNY/RZMd6kMHgVYyBygWgPUN+XxhQHLro8oV/b8duGsQOHOS1
Y8xl9grnXQL4T5c0j8R6bFoW9ItFNo3h7Q4xE813Avx/sb78z8ZuqMS31ls0bITZcFmrTq0D0qHI
5DoHDlSs1fp2QIZ6fcLqyYT2l0V8Zy23UC76ww6jDDUWkedNaxAk+RkKUteEJ8OQPE51S44GU6pp
g6DQT0/O5/hTTAWxR1YuWRnzma2o7n1zb7sSKzRgpNlN7XQ8aSxahKXLGApU85BpsOTDGvTna/5g
McbHfkoGukSANc7+H2hv9ewO7cc1ogw25ShaIaHXivKdhXRGqSOJoDSKgfZIU1DtVlGIzQdBNJmD
fy7da/8JnPhGS+BcQHazKo+nzUgyFII+tltzvD8Jpiob5Wn9e5hR7CCyU8mRdebOkD0tjh5Ltc6o
Ye5OofY3qtUyYZSd5OBeIWdqhqx9urnnrdRPQIa1JJW1Pk1zYTim/TO8BggaqhT0sVWnxAIWn73a
/Xv/FrVkb8lU1Ptz/fC4yP1G6CHIsEzXkF5aQZpFSwILcYwT6vsgAlqX679fOODs8lsHhv8Dombr
JF3SWC3IJ+N8KMU3RO0UXjgfEUXBeC6offOj9ksuDFZnXW14Vq64/AdxDmjk2u91FaWC7g+AgO0I
G/Vv6iHJxY7rymJW3rQJ+EWgnw/1KqjJTOf9uNCmy0hUY2fbGkJ9Sjf0gyOGNmRGn48ZxAQcIA2S
NMaasKCH8kEu1BTUIAB/leXFYbvl2ZFXlv6wzq3EKG0y9CgOKDvtN3pvWjKtiQNjNEmamoF6Lp5g
pguwFQnOmNzZkYl1CouwuJXTNNtLGScTPp7Em1jIR03AEdTa9bj/fSCz5DyWSu7e38Pxl2VGuAWs
Ge6/cvFrAKJ+qs7Eg2ehnG+l7SM14jKdMtim09/8kJheangDsiOpqVnW++zoCK5RK8h/mXL5llGs
b4u5PV22aD6p5CvqBJ94npAiBnAWrgtQ7RHtFCl95lgmOQDyk09v3V2OofA2IDuFG38YbOAEYQae
qIY+CAbWQUj31rNcEWksP3h1bVNwZNx1bR5oh5v2FV/AEjcfP7ojNcVgift0gweJ2eHD+ZnKkfjk
hLcVOeIhyQKmBlu4EiuCo01V501ppSoYP8GJByFCetssERpHpgjONbaaqcWXIFibqMm/PNVr16TY
7j+qis6QLQfZq6mwh69z/AnOmRyBuO0/AjAh4DnwfaWFulZonbHlGBj7jEDkoetASKcMiYyglee/
DLOck4lDCUSvt9J/mA4t1PopOlkmyHbRD2PUO5nfCD9tnAabDkPrSLUffoVNCxJSOkPaDBPn5jS3
QVH4ulQ8FPfocrJUIuOQWKeWKlCRStIUFlmpeRTr3le3rjgq7TMpNJGOat6dYg91o439SoKXg05L
gLpYSKyz0k8JulWKF7yolX5dDS7e9Fx1g2trs+oXrfcqi9EXrVn+HrKsXhx+TLTCiZPROtPVomOP
oY3oxXwineQZmj5r17VGriSr1r2eTduGEqy/auWHDAv4wVjELhdUvswbErqdV9sxylEXT+6ZI3sY
+f4KQybt5vjO91RwsEUc9PNnAGyTTrlVvf+BlwThk4YCaR3y9AvPdmwdlpH689TT2TaPU9vXYHfs
KjIkV1metRYnDIKJfJUnpghoeYI6gLIIcjcJbKotEwuIySSUgcbRLhLbyTAIracsQgmvCfzwaz+X
igdkCKWsj7FHIJj/WAi3OZbObS4omFtqyR5sjMD5hOsoAmYkDwIidwdnOtDLhsdQU/oW8221y4L1
dzdSTLoPE17L6gNH6hZIStkxHVedFzXzMQrM7KC2lSfH0J+xvff23kbmh3rsHp0/rGoX1wZIK/ol
rgfGmvUTtmH1IwWLOQWC+4asPXQBpdiHWh7ANuEKazmLKoJUtIrtebnwPjD/+HQgIPSyrZ2XMTpg
LpR2Uyk2Yln9kq2/Gdbv29LQNZhwvkZFIQ48h9OFIdu7cXAaLULB3dqRUBuZnrOYFwtEKT4MuMWX
4aDZrLf3eIX+AzvjDxkjx3a+jLdiBvMgWBqhDnVbPOShAmLOrspm9XaWh/VHTYSQwuF6pDrmmU7h
q2+egnCZTowIXgcoDY7s2Ht/jaP9vzedpQ0HGJJj+Ir/rT1cP4keu3GU2/2ZyAL3fq2XYhzA+MfL
nIhFHaZPEGxvtBoM5lRntemPP7gt1CAMybGLESraP8Rcfd/OWgxEtr2w3mNR+tkAaLS6ZF3UqR4T
eAvlB9NYui8XomTsk/lzdniJBTTUBy57Qh42z2Ckzp79u43egyW8cmDzINlFzzb/aNFcBJdPedou
zch3SfcwSKM7EyT0JcU46QkIn/IdAIvFou23P7b1ygqT/vFZNieb4wFsIJDqIPaUmW+2Yz1NQjcl
TwB0bnfiHL5utyDhSpf3gOLhb6YXLhwB4AZvauDiXkz7nKWMfo78AaZ2NL8oZrkhnwrEKfxAbOiX
UxjUEuHAuhcAwnwHYwvw3F1RJMkV+vmN0Xf6ahJ/6D8xqy0C4Fxxf0WWJO5gPo6x7r7r4XVgGtx0
sORhnwOW2DGHHWiJOyt+2x6z6Cz8MANV/1DiYcUXFCuax/cGjfgKwgxA1llYfMOI3dxz+Hc6GD6F
2OxgvBjqrF2yHy1AO76V1wUIpOG6TzkkTl6Xb0L8jHqx6+CXoiHRV5xNC+36emDJq+OWeqbETa0j
PJHi8MmSXbQR3nTHW7sSzScU12+cn8k156p8nY5s1ZsIhEjFKd9eQtbhnTYXqLDYFLrmAOPC7JZe
ij1pUpQSjZPiyEM75ps/irARE9jT798CnK+sYrX9vzBEpMYEz1QqiXfPvCqPILzJjvN2jAND1no/
ha3ruBgAjvtRFCLn5d9IarC7JKpKPA/duKhBiMjMNAqAuedvIi48X7XasGqLMWeouIHb9MKixVPM
RaK2ai9HjvaavT+iFF6I3DbLa6nbELecdSPc6eUM7uH/IRnKWMPB/Z098IAQrm1Lhk1gQyNvB0HB
HIV1NZ42oWilfioXZ/CWEHlD48V4N0n5Fs05b54fcuRTon1VXxt2MDs85/bcs8LdpBRDsObYU6F5
+FMr5VYBt5dv7tLBZ/apiCBufLSoQL9OFFyp0Yskbmfi9bMuS8gHQfa5Rt2Mh1Mlz4r6Dfkon3YM
MXtHR+8gdHdzNzXc6n8q556jmrP6dhmfQ3vvqC9Zp3tgqM/Mk0xe1UWaWpYKpDHaDNj9wR/pabu/
w0mpywQjmlhL/JwZIonUOJD9eHGnRF/9PuwNz1LKgkzNrcwogu9gRZBeBQ2sTy/NLDBlfYI1mRAP
kD5Rk3IciTeym1DSiovwm/yILYMzSt9JZ644RyXhPEeFK6ghz7LxR61bTg16amKtI+qsd7W1RJXv
3RW2hYRaBdRUlyqFmSvxDdc9mx8BisuVs4QiUh5xYt0Tz8iQncohTr9P1OFru8AoVTbAGOEfjJg+
QPm39jh5FKfCc81/gJcwTHhJ1g4Ix0BZw18VUr52g1Gj4jKl98+R9HyyE2+wCvLUA+0Js15ydP6W
NJJXrrIoGhWf15iSxwt1CBz+ouRH4R0702TMC3CJyPBGvAY7z82KldVSW5zlRf/pSs6Mx20qR5Zd
qkFNOtHDwCart/CiyVOWSmFrvqCO6+po897ZMaVPwg+M98D+HmHS/CKB6/teXG0M74yXo/8w6XYu
8X26/4Fhmfvy5d/1+xQROT/N3FkLyPBd9AjzCvH48fyyu2Y+UWOIVckmyl3LsuRxJvtH0R2SVK77
XFYOQxt5KhmFf3j9ACApJXN8jgFVU6fJLpl+1gZ1Rqjgof7jx1QgfiZfe2ZrpoaDd8+2fi/CR+pd
KzT6R9BGz5sNyWIg8e5mJCS4eQfZLt88pz91bHmTSdxuqhUUWA+f7838KzT2y3XPqG6AmcmbYp+j
hVgw9zc+jhXbKqSQVZCRm0OPt7HesAYFf/q15cXQixvkIdWPu3osJeyoOdAfQlrlN5x335yIFPRn
b5eBQgTAyT4ETg4g8xwEltARrlN8PP5RDMbujBYbfkOukqTWUJkfVOvCmPj5bMd2mRDFpJgYZpIb
KNWFQOQG6b3fKO+eYYAkn8/LnYfKq38lD2PwlzdhweB/fSLcuYgSwtcFtyCN+c6LwjC3gEJjTaHa
sUGwdqrRzTpVQLMVQEDzDaWcVXrj3+yMqBunWg0MRarVvvJOdwdOettXJBphFbmKB+0CqCx/DdxZ
jOditR8tJhfP2ZE44kvfZ3fAUvdK4lz4R6dqgmm6Lwpf8l1Z+SyIZl5UXRvQCJgpW/4Lk7GDZHTq
R1/yAzhvGrazHPlcbMXssJHLDK4ZQr5eZhM723GMm0gQcEJdP//Ao0uNypfmlfBQ9WLajaf8gKnO
ZFasl0gbiHHBFUBe1KKp3or5DVg24+oiZPdK7dxjrcrIf0rmdHf/AWh7fJ4j2GrsIwpuOn6gHYfV
QLmVItmgKvQdLboH1BX5yb/MrfOxHElvTAZXZ6mnT5JXfFscs2NUH+waTP9jbEoKzU8X7EeLl0nu
Y2VzUp2odUocWL/MboDte/hF9pvn1/on6iITb0NQ63HCxp7BGePtXpu1xevpF1BJ/PhqY8mXm+/T
N+RCXiERjMIUoKl6V3C54Zbf0dpf+avl1UbnW/fHFXXY+2xrstT43uzuPuD5IDkciysqovGK1AjC
GhpKcQislwmZKcrjMS6SheCyLcNo4Gbk/vYOJIR5pFk2hSgQJ++Ra0WZKN9HHxM1GcyWIEjkM9h/
11kzxExLqOdrDP2AiIE0XRlYNYDwFqm2ePy+lFMTuZeKD9qgFRnfNo+uxVXNZjXVWT0iRRyol5cY
/xiC7FWGhwMQSoeaUlrsFeDrw/mDcgS+AeD+n51+rp0bQtXTwwmmRLyMJ66M8gdD6wxUtfoBEwjO
FBZ8ztyt+rXssT0oFUCBuVN7nRTt06FbD/Iod6ZyWIh5bnSXeMA71PfUtWb9mVHs1fUnGsAAp0W0
7Ia4oq1h1If8eYok0DCIr9R1Tyj/eFX3jxriZySEDr1/1tAiLR/47yAzo4/So6xBfnjG3Gm644/p
j+x0a0AYDYIPgSh1iaYA48z//SFKgFNSqpzyPogkX1hVvkzwkCo6eCwD6U08VtkR6s3tmTWo1oxY
iSd2Z/nHBzr8h3EUIBOtHruo5OVyr4JgxdPoiyqSzOZDAukE/GspmWydBlXx7j8CfzjRMzowFOas
csqIMgs4Y1kVbA3V+YwiDkCcMUesJ4qDn3pqcOKvoSMJE7AedGoTIsYzd/T8VOQa3r9uHmDKoVlN
3ePz+mAQpxuVhyeF3tm5UXZFX+SI+ZjIzzmZSo1NiAxk4sIfXcJg5tw6CS6239MQoXR17Cs94n6+
I1/iltFVFN9gBb8J37q0Mvvu/JWB5D8H1CvQ6Yt2w23d5NroS8AFmFQfr11CbdEGYagcm5/L81yn
UWYB6b5wjRPQATKlrld6vzHNRUPdqPnQHo6yyxOK9mQfhmtHyixs8RkCX7hkWCcO7T98OfP4Fets
VIxObb3lM2xCG/Mc2TJrvbuN3AHcpAXlPkrklwBGt3aTOvcLuVTTo6FAA7kMyIbeS6HVtiPGysDs
WbcKxJbYpI3CCGLe5VKoR1kbEu/vDo0yBhFeAvl0TFvYB/xTeaHJ1waSyIGqLoXlGA/ZFvVB+EAh
B8NwcPRfg/2Hx50jZD+iwOTzWmA6FWEPh/XwYl9eno2OcpKBPnVFFT96wM4YUpktLvypJRSRC1Vq
bGnDFvzQAatom96yGApIURE4I4wlHLQlVlKbNfLv4Cm4nrkRQ5/CYyv3sdlwQwHr6zUBfRMjQhoy
YEl1ZLj15Z2jfCvQqAhcZ8MkP/JbXEvODPIzPbLaF1I2EDCxfYGedFP78g9vqroRtB2UZHtew7ub
BuU+2TmJ1mmGLrz4CT/SvKyS2DXgIWeN0lspnloRS7yA5O59O73W+4cd/OxjLOjhP9PB+A84KFos
yvyuKPQVazVy8d+3TdmhoVaQ5av15WfiPakuHct1MCNhnfn/wZ1dvAHkSoQKKTbO6SaLfjugXHVW
lk489KjG6XcWb8oBGCkW9KceDRnCFQ+k6YUZ9rBj7+sgPTe4yHVp6ktcrr2T786tYsKSR1UXMk8q
LtxISQz+z/qJFsGDQP2VP5kN7KyO+lXbUbMQbNZSnTzJWr1w7cMhvpJ3ugrBxH4rfdsgzifZgbHq
2KvM1uvlSQ44Kk3BBGTYOLEaWgDXpKGRWOsNE69GhvHMe+aEyLkdbGDqIn+6fPIRCt8hJsa4ki6P
CEFp7ZRG3/ZU+76J+rOhCIfaNqeKlr1PNk7uH2xFC3LCG9UAeDKsqLoeMAl2jB13uxQ6NxX83a2S
zx56jeRPp7msiIpHXJpDsRDDeNC9SsRkL8X4B3sMUzdQ2VuGYhPUGXroqouezMnC5+DwTtguNZWw
LU2XGTFp8mPDCH2hYP8JJAf6x8c9qKI/EhXsosPE1p0FHtstNfieZzCkhW/NuiTOSuvqJ2GjFcuo
F5djoBR9k6XSGeBRIMH4OvUioJ/pseZ3fJffD7zkT8KeZslttnrIUiALZZYrJOxdc1NU/0eMAzK3
/U8JUrlAsjU2RySmyh7QYtDP5mazLfz97tGISVvPMEIwUDUYv10t1SZOas5vG1buL0Nv7fG+zzMM
HMuo2HdVAlg6i8KbHHwNcTOCp3qdLcSCja0M35/1z7XpfQKFYUEA68TyYQJxQGGjUU67qzJdtvLD
da4e6bLuNt0mjmEOjofRyh4EKGfbxCVj5LuTW+h/nNWidY8TlmOu2mqDbJlQGkjDNaKSVdTDrvnB
iAQ7Sbtfze1nXdZnpGueWJUKq4KcK/djtf4wLrOHsKf78+2jaqrtHkcTg3m1DqD0h15zb0YSL7wV
J+vic39wy97M+xI5fRH2oSqxmtBPILI5zPfa7GaTbmNBf6OEsZo7CaM03NryCrPbiIXmhWVWT8D2
7B/szy3vuXuJVilQ8qB3gdoe0LnP62fBIFygEeuVZxaLXHBstNlU4GAVypNkVZ7fdcKg/QTMaAkN
di52pJJjjtwDrwoha+jfporUuRS9PxRPCz5+co8y/xz/pythTcx9/Vp/7iDhyOMZopjyYdkth2/1
D+4FDxeoiCgSCL4ETLBxeAHku4aIugDCz2H0xqzDxik/WJtDfsWocBbUWBr90wnMY9uwdScxhvVU
BYxRNj1lsph2h/YZKlFiTFv7Tq1wSyqSObOLyUPjGCIawp11a7GLeDdymXBZ3LMLY6qyf5Gm34ta
tldBFYKtfhZQyVeZYfXHGDkfOHitYKaRXuI6T4eS/K0rDSHD9whgXRbe7IGx5dvT47LUjfpp3Mp7
A/BzpvNQbPIs2jCYFgVgtfTl9kkIuvvHk3sElIgwybxEybDPUAAXKoGQPFhGGHosVTwdFtZ+2u4e
6JNzOL8xoCvrRSAF9wu1jGjaQ+XOUeg+Nq9lbhDwtXc12aL9iDpybnVTBLFcsp7DYpvvxyBuMini
aM/2OHF094mpm9pQLR482b3BnmF+69of7+/Qy603Ujut2D/1Ff7ThrzZYEKvqpOKTnvFZwLcrrLw
p7AtGdXQHVf9hcCvgutfc39RQ8Arpuvgcr9oWCii2gmrbicM7eDczTAwOGV8JbDCw1cM9a+WvEQk
1X8HsW/eGCybQk9Q+kSWwk4lo6Qgr/+Hx9OE8J7vgMGQ0Era14aadCALZXm9BHv2pPT2JBDKoG9E
ltuHUioI2vd2bJR5XDTOmQLtrYzQ4wBHd7aQPDdcJjRkLSUUEHeLQ6adwkbUuGB+KXPBuWv2FPZA
BNli+fI1N+sGEd6AjWBdoRaLE9A6LJ1VQ533DxtxH3ykODbBKFW+JiyO1Ruz0kdUfwr6g0neWdqt
HVWu4jOl62xV8Uqksl2VinRsDR0QlUuJqt7Vo1O+or/ydBf/RgPNnG5n81cypgyxsxLxVNYqQCF2
BTChQ2OjPvxLLf47i+bexeBXLwZRjV2OxrqF5+NGCdW6oW08WfZqZ9AaqYg/j2GFyTho420eYRot
h4SAaYCHXqxI2JtcL8wGYTNPTDD+GPQSeqI35aDQhjzguAONNQ6l3vra5mWhmlLpa6ySggrqw8Nr
paSYCtsqItunmiLaCFrlgJoA0fEmnRfhyyF4RS5Vc2XvdeNSDG6QnJfKi4rD9pyfaiLNRO4tx4s5
rCR+O5G7D3prxoD+1mG7qnyuPYvFRfgomgDgvsnr7ynfQ3YZXckqYSTaRYo8pjWh5XAkfhhEI1ts
qoRUBBu5JaYCFOeZJp4IsXJ0F70fujHJIR9CMFnU2+ZxBCJl1ktIN1fnFyKIvoy+aHVQ0XFfxFhD
8iOOi2B8YUKho4Hr+WpsU5AoCIV9utC15hHJLbOUY4KJ/qeW0uSqLSLz9Pe1s40lHJ9VjhiPDAIA
e6zkrPixUOHiVagWVv+GGMDFeCVWNg3ntYI3CaFh6+ZNZ9ZPYNVUoqRAVAv6jNeVgLaXdZt2/79y
qm8UppC+ZDhD6/vpJywRo7TctKorp9N5ACInwDmoGNXbh0AMcanypVJYEg+55udK7nxXGgzNyt5V
+ysu9UDPbk49HkzQCHsZjjGl1fnYULlEi0oQQKK2Stqy3495r2ll1lmjzpjwz6b19ELvDbTBrQvQ
R77f7pel+y9GgavuWIfLVHFbYQBGZRFfq/tEnjvsqcRN8Gl8OCG89RuMHiuwN3Ux1P9IdzM1gtIn
NynqpkDoxXDh3fRrHcpRt6Ur+ovBvpOPfagDvCM9Ya/yXi+rvH6tKLrE4vw0UINLETTmFuWEIqT7
h4l/bAR8P4BeiBuHAzMcA9lfb2bDEHP14vjnQ+Nvcb/mTLHXU1Ei3bouv0bCutZ9l7iiURA47HG+
8JlNgmbVGd6jP5wPV096Sc10mhBpJtr6gbzQhJVYTRMOxtJo2JbIOMVlOm+rGycxEtSbXF5znyml
Rec/VaM3D8OZw8Hpe1UXXOnenc85Ett9ab1jfKEtUtsw6/S7pXjyzcoFj231ZEYxQUASLqzfA/as
yBqK43XX/mzX86jb+IhptZCeslfO67+PIUJ8EI42az8Enj+EQ9RRZQDgmBlo+K9F2byv1+kHMXQp
n/1D4S+Ya4+gPngA0LlHlCBdBMisdgE0WAHJRsuhCTGHVKrGblqYrgY7eBLQ+IKjDMldhMemQzuT
X8250QkUUnVX3pNynOztMn87JyjOAvcIL1ZWb0685M49eqi0rPNvn9cNpmwVZ9UNyCh0M/Uf22GS
GJQLKPedMEkLeiHfgUE47NkVkyzogym0pXQ8qD8Vflp50r6WGXXJZph3MWTBR6x+LG7icEJedEpr
t2Gn5o645Id/tVW5sMByasMCcLlKL6ba4fPdeDS0UeW8TvfEyzu1HLcKsgxxBejYPM1wta3r+m5y
ztKyWHWxXCQoA8ZN5bZNF8NVZM1XyTYC1aNm14Jvbg2+1sxdp17Dg1xiMHzk74ChWzMX2bzbqJ+T
mosRQMnX/f8FZL804j4v1q8aK+EfCkaB+hgzddm5SRfX7ryEDdl5olIGlJv3/6AZrFlZuyHOki3U
hfIjJJtiABJ2r0vJ7BwcX9euXcIzQTRXnkoEpmQsH8p3y9I9cmMv2/HFTZyds+HG+I1zChf5s/Lh
SP8Db/Tck4H1p8BjolfO+w7RDJcoIWb1CvuPFnx7dIE14Vipfo6BkmYSDApt9WRJp/rUweVrODfx
VNoznG2IVSbDFeV2Z/AOlM12aOx7GsF1Z+fgc5/cJmmvHXVNu9CtZZFp16CHDwLBdbWCPr3/4QUl
Wjhg6Xl+QuqTqpFfDsNeWbUoENbrHfaEuTiGj38Osgi7MlmmvX7QmJt4q9O0lPSjBWq5J/qj5VuF
sMgxzhcNLvP42fwzRrXdq25I9DysTWC/7bRXQTgjmyDfqI8kF5tBJeLX889FD5wJP1p02PFvXp07
/uDl+VWnpqFdiqw+jnqt4Y/D1j15zPnKI6PJOmyNlkCketYNDiSl4CJ+Hy8FRB7xusqEyTqx6Bzu
5csPTrPa5DVdf9kjKL7hC7PsrkwYHTZvZ9ygvTllQ7LyWnRAS5vGZ2UvNrqnIaCT9ignIeo++Ze/
liw2rsnMQ8J1w/QUO59yus9yF39MZEbpjk/4vVD/hK+IJk64SuWmbmlykHKVn8UFIntlVM6fcKFh
cZ6m4Oq9ubJVLI8+5tPycKDTTi2bAIEeDOSZwG1gIdF12KUZlB0gSyBV0ROyf105jjp9n//pOpIr
MJt6cp/XtevJmh9w8pX9b1DDWYF+q1pjo/NdyolV3CwHIyKp8suA17lFkFCCuetfurItCU5FD5iu
+qouQ845jAdhXvpdG0kiEjdIKrsnAY9z5rI7KEouQ9mmKw8s9LCt6o30b40Ey4fWwt/glLpzEpxv
gv58ezC6H0NATGPM3XQC3LL9ytysQv4tS6qGlWxZxnDhOJbq79WKcjZfS0VdMf17c3Np5BUhW5ux
pwq+ydRuYylqG0P+w+lhfS1Y9SHMz6XTjuzU1biv/Kk1pyt9w4Pv0GJ+khuYq7EL4mbONbe4n8T9
nHkcVNIi4Tul2KYkQ4RyoA8lJwcIuPy46gZmBYrL8JzTV/+NkouejGyZ4nMj2ftUE9aHpFi+8zH7
9+hgPYaBAdlZKhaknsPoyhZEYAEuGzRsXQTuEmx4JNKc+TZBXGY85wgc3zpe9IYdTsiE/Ss/+gCe
c+hvfR6AoViYceosb9sG3WMyhZfMHGqGeFgYjeg5a4PiPzru1GTTHbvBIGuonnVp5VCejcjlmhAW
9dp+wN+qDh9R+Y96CXInzAYZFTXZE3nBB7DQcNrSMZAsTxqoShF+28RmhOJQF3UkMNa5iYlPsQBE
DqWyQq2dimqbcSVPAr6sk3SsfOqvf3EOyEUganqIKwEhor7Smbu+VrWvBhhe2mz2PH3fvYTLLLAr
bYnME6diT3omBMd09CAaesPiivI1EOfJFxpaV57S5/W62JSlyiGWz4Eq5mVByc88Pz+iom1McBQW
IyFPQ6pBAjkO0U+Mtt48NqrnNs9ShUKzbNE79ZEq/tcgBpH9EpIhaD/iouMdOZoBIXYEms9PqdPh
PJofPUV9XffOtENd/rYnqRd5vmCR9Zk8cNtXCXKZCjxzlpaNixb2jCzR1yDmuCOPnpRPWGhSRuUm
GfNtItZZA2ZPPCth2HuExEr90Jou5+b+yaIwukzimO4I422TteoL8b0wlWVpfKHUG+Oh66bHqCAE
G0zpd1h5RIq4f2Wr2EG9EmeXu+z7uTQRSwFnIJsMmiftSXSxuBY+QCmRZC97NJsHWCtYfe5Gu/nc
WYvNixSSrQS6CsVHM2UWlCqfI9ETCjWcBlTyhZlhHM/r9VELklTTiBRPQVJIDdJUtdhMm5CPFw1q
7nBsB3dG7oKdY8ZjMzYK4VcfOlbsyCtAJLwowmXvGsR8P3fsbI8LomcPbY5E1VFe5S/ee/piD0Sb
tD4JqDXSB2CSpzw9mDfsMCecSl9sy0ElYCeMix3DHjfbLKFjxfQem951b/qS5ruCynTMQhby5wKQ
YZbkDXOP10N3YW009L+ZEs7MterfuaInTxQJkpe9vz7+P+0Qc771LUscU5MXtCiS8j0xvpgB8ph0
7aOrDiflhUO33j+wdw8xEFjQAcTuIXxufQGTbbUGs33h6B2nPXlPlqETGL1UCcvdwcfUWGkvxxO/
MIBS3KtXpf0jxwUvEZAxI9jw1DLax04lW7AIwdnd5UNi4OEV6a/W7ahOrIk7ns4P2Y+EFdIy7XJb
ZjwLVfel+wAEGrJKCRKBdVDQeIchYQ8BhtlE+w2T8QO45c0erd4w/PH18aF/VVsf+qcfGtBnhH1/
WBsdt/wetAjZy5cfDVHetpGssDAY+N4L8rU9oMWRxBIMg0Or+yIaMAcGiY6+DaM2Yyu7lGeIIIes
rWFjZ4JjLSX6tJBkf5Lh4nUWfN17fFlTa0yalqRAPvLv621kZGAb+paMuyDshW1ueZjkHZewgVME
CGyBIo7rpTNNZWcmVKgBSh4V9CjkFJiGbzdUQO7CBzLhwHtnOW7m82N336yNUcYKxoUI3oaf3Gro
iagRX1Y2/c62hQgCr/X0QcqLD8B2KJ1JYfwEUYr+S9vn7YhYbg/DRBHCyhjzwjmdEnrynrGjg9XS
oHancJL0VMqbp0BSyW7R8M7yAIaR5CMzt60Rz15OgqDfxBwzGem6nf3ZGPXg7nT5FnuKYYYAByiF
QKKZSwrS/a/A5EcrfOliLW9KTL4BDB/TgakcOqBtKlsclJhUhhPSbJUiDnRXHxO01SsdstXYhSDd
9djjkF+ETk03M2/q4nY4CKi4L4P8ISAhOFBPN783yn7DwyEZYlQD8vpp5Znp0tRCEw6LxvlfWGkc
RggXZPGBO/KoqWPy8DnNfDnjkOHDn50/BsvYh9zfqFlrCaUxRFP/3CjJbNeI8BwU4TldcDOSUpAS
QvgyNhNfh/+goKBF5yj8glxVyVckqFaoq3KZtaGuaWlo9n5N08mQsTmYqPLya9w6NU5JD5rfCDVO
vVcTMdp17F5f+SN1OO8KDEN/5JRob0WsMCCvMYKCiOtADrr3j8t+zrY8qLMfuVlsu+0vERg6pTwD
NedgR6IfqHGasIOrqYIRk6XXoe3kGlw37X8137QuDJRGwjkrzk1LO7BU0rJWeu5Mp5WHptiZ2Dt7
nGHzVU6QStsZ6Cfcr6fQSquTMBsSMhTRKWRPOSTudIP0T9nkdHeSjhV6XoS5rmbJHJ6ypwLjyu19
fs+FWjguK+NCeAqlbk/TqCVsEJXWYkNAQqdSriPEgHW/6n7qgAyqsG/dptVAJrYbhQXD2Z/46Qsy
UCVkdxzxJWUgYAHz8A2u3njSeuiFgSwqxOtEomU1K9HcDlgwQCi67Yd105dHl227RA1jJu4Tez3D
JIdvX51EkT+n4LUyVzT+dvmTDKxETj23f4rFSdAPg4MiqljYo74wzgcJWRlicl01IToT2l7rvH07
cLH1W4clcbSA0VZbHuj5FWgditWhVZIDpEZkVMpvK6y2guwJ+V/xeYq7TDfxV2ncWRiTDBZPQTqJ
Q2X0cnDIvA9SQs3ygN3gr7jOpdp7TT2UDM6oxqDUwvlpp4xohNr09gWkaMelO+Y1x1dHKJP8xo8A
SWDSzocV3cnxDkswNJmoSDEldfZLf4p+vZdPLMt8uPkJ0KkMHLumbzXO7kjcAWm+CIJYr5Ijr+go
pb0XRhk4M/32ze51j8dmZ++OT+o1CkL5jx4weqVasfh3WJgpNUtGttF2FZujTWhyyjkFGGUyS2Ze
f9TxaqxubXE0IkurZpwM0nb4n8n8V/jciIJ3lvXxxgKUSB3d0sFV3nKhxXwQg2abNmss/P0wvim1
Pv5dRwm/UbYwAyVhaT2xLYYyL21eJvgg01rVFqynUog8hm+aFOY/5E0j67BsS7ehXuMZVoDdCimH
S7BgcDB1YcZrYpLgD1Q6yrV1HcozswmD+aYvNxi1Ew4PugiiUtUPbtV754WUnn0YMRVyEBt5LABI
hQgXnnAHlt6mdG6kTm+apqijhGPqd/5khktv+ZJJvzmzGWWYvT1ZBWy3xRst7471ixgZkrtCr7Sc
0xFjn4Sm3H9EjG+dYqXkmmVlFfg2Pj/tjzoI30UrCPyBBGZxPMRBQmrlOx/1XAT5vg/nKqF7uVZ4
HynsrNNoUup9xSJv5RiT+yx3Xe6pRkucO7P05gzCMQJILGMlhMuJKfj3brKIpVtik2tjxNMbW7p7
9nclzlMwU1S9MOOAY8vVxljhaffx3htGdhGi8d39iGJbCPhndPMQWGdketkRS2Q39MuDZjpQmKMe
/j7kRV1g7tJzSoFDHpUqpSTCLkwPlzScFIRzrTl2wxtC8Mp7FJqz8zgoReZ1ufXwEP1VddXR8wju
WVRNNVb25V3hHDlGdbdTxkbL+ZqWXtZZL8Ang1cUaHQL2ijU0J17sMIhH4C6UjKDlKemI4yU3SGE
CwjCggmTwZwN9BT6yZ4CAOZdoy5Hw+MZ9UrNSZyg16fzuyuP66u1veM0TQnipHcseUzgvzGYeyCE
AWoI3Mwn3JAUzndR8rvB/ljyLZwtRrZp8jtqz/cLSznqxJMaxPoPtIASqbRoAoboxDskAbFLqfYq
74rEsSyYO/DRC+7TdE1eyFQbNcHaQFPGEPJiWGZxxY/829078FghBi2W2TnMY8jfR3pSc+TnFbI7
41Rkx3jCsYZGvERyDUAtPsMR6VXOu6dxV6dcJfq32YAtTyzTPzeAFEels/g+hEbTnaPj+aIO+msY
B+izck3a29tRr0QGz+7BsEWQamzM5yuJrGb06Zio6lrtXkmNJUsdR9JOPdacJbXkyYAohr6NSqHr
x+UtoW9EF2F1VO3tvghCums25UBxQRXFSdF28uEzhEnBY43VHlqJzAPIXC+3D28Ezly8MDSAE29Q
fKFWotXdn4sDUcCIBSN06/wQ6as+1mxUJoQsznn6j0zHo6XcOTlKuI23SuwHCHmTKvrADbhARP1P
jG5tO+3cEvZ1L+DpwqJVcy0WWqMM7OIOtGe7YNwqow0gav+kl+xiDzPQmKMVo/0BdrvbF3t5N5/+
IDnhNIuLEOy4sVsCMfKcEBndz+LrkT1vaXlIgNJWMjpk4WZqPATa7jX2iUk5w655IuFsZ5GY+XgL
uBdprqY5j0hPuukiN54a/vsXIadKGjsfRp+wUgwGfHHdlK9PgdeTT8XeD7VMU7HebjLgiWB71AnV
UtUj1hEFJVqonedReCun6+YXKlISg610fsY65UlDGZ3DCkZqvawkBkqe40EYJvXzrvN6Zh8nvEQc
XjAMviJuQs3tg3DWDtqL0hFPf3wyi3alo0x5Gf+ldiiyfz+e9oPe/rKBxD9CENYV/vII4vuUnhRV
QKODukP1jOdKpQVq1846O8DSq8VVv/lX/8c0PbgVILhkti4SnYappHy2nsRAQZjrt6B9jp7P70gS
Db1o8Kmky8boo3hkSCMJO6FQe+NM7PQS6MzBZmxK1i1D168I5sYlrN5JUbxRn6h6OVRean6NLFxe
6UAMHhXdhcS5ulbIf+G6IyquLmMFS5Yn6K3o94SCXItudEcj0rNn/abQeyCNJFfDcJeonmq45LfP
VyJLP2O/ZmPBltrMTmysWP+eH7lqIhosqT4Nf2K/G/TOxuKT68Z+mHAbBJRWr9ibqXrGlfEgAolJ
TcTRDr9RyrnrWPyE9RB9pUb5o4t9cRdqme78pPB9atal7nZcm/ybhenLRrvjyfk0zrDfJgCdv1kA
ZFBDzj15E4Q15IYR1XAxd3gVKhwFxKJnRmlXIYGhwGLGI1S7I3dDOSuGrAzSNh5uUW1jLA9yW42l
8xOg++bJ4M5aVH/kTu2DBi1/IweyVVKWnzBXj2ttUfKp8mjqJHqP5kP5jb8VZWamVnKhfgNc8imw
zRR/Ve2iV+ivnAlyo2bNwjM+rnR9g5a3pFgXdRabklqE5GH49tzftexsfc2RG9y3nbDJgUJ1OPLl
iklm46/JfhFdkLpjkqKgDwDGqykkddrbDLwoyehUC2O7ZHHp7gARuiCC3j3iKlhStGWZh2ajeYiF
OApyueceI8l9T2lOQp6CfhbwOk9dD2aXecsN/fAg6Orkj4F94NFh17ALZhtsahYQcSM3QmMXkj/b
2HKKTzLjEADHM4XTZhcx66ycnpa7M7vXv8rK7bZkN50v/H5bamtiWPEK7/MnlcDK2xorWKVWPRio
nFuwSp96aNmmMD8XVl7lipmR5lXjD+HML22sAt2OQfcp6PsqGUGiVfwzC3X1Xgn1/BU39k0riF21
kDXrmORG/iLzbjzg8242CW9WqdwipdzWvnXSwmU87jsL5xOZXXk7Jk0oWT2a6ukrGFSVT7Sr1T9W
72d6BNfRM1kz7tkJnQRwAX9OxwwkMePbgRcr1qpdZEQ/RV0sp+t/GgnktR4IhwINJ2JuVxUnrCWi
ZnhaQQwFAepLwdhMeab+tjUZan4n/WGu712y7zKQdfTEGc5KwfE1s8itkHzafkDkj03bFePAwAHB
jA6jFBdIRARbcPA/o0BstWqtg/hJeEwStYJmYidc9IoIRpmR55jICJxasF2UatT9ZET553YmFdjk
rTGnm6Ca8q1MQthWyN30CH4iAGfPcz1joCf4NnVwDEaMi75RhVx4Un+yzbYF0lHicEaT5yKlJJep
paZK4AjNRqiddKci6Nnhc4mPL1BIXNXm5/uzFx4FbDImUy8zughC8XsDcEdz0XVrcgpmIRpUnJh/
wjsNaThQh7ug/evUTpIVwxEFbgbTFwFufDewbXdfTyzCqkSVaLJpf7vNN4mIHLX/1/xvztxAA13M
aohmzrSSHmuOkc0PYC64mq5wZAmKipd5ddQwuWmGWA7lVEUTtO2tnxNd0bxTWukKemCIgBQ+TD2l
8FeWSHc1izaop2XuMVwmE8uKhpSutDU/ETu18oCdoyTJTOndG853VCQ389yFOiRqX9ohjwVsbX9H
bwIXclXAaMYOcVehADGG7Tu2D0qq6eW/cFn73DIITsYD3xa6URho0Y8DV4x50bkFzdHV72WYvJi9
N5D7Lgz7A083GXrV0Wz3xxPS2yLk4cHFKykL9Uolhaw4lIEv93atj1AGABLPYo7T6kN4hfZGxhMj
ZCH3FFKzUCCA+sE99W3t5In4l3puLSCFwN8zhPASZhRkmhxkcAx0OCpydmm6OElEX3qGn86a0dF5
YV3IpfZkN2C0VaF1+xDlPw+ATcaL5PVVskH49BJ2gS48L4QtB5nXtIPrHi6VTm3lA5y50fjVw9Or
CYSI6GhmXaGvFb2VYKqvXdt7xwCby9nI1g10rQnJPfwBOKI5AkS9IJeTO8fphrP7r1muV0Fa4j/z
ZD9lwQzYQo+ZSEKwoFs4ijF+dMPC+JBnP9KKYbozny4VcX18fsrBSiujBJ2j4EweORaGzvrvpMFi
W6x61Lvs0Rdzws5WB/Ms7pyW9M0HzJkEsP+sWwBUBbt/fBzY0F43LJxtofbKzN3nDoxLFSwRKq2M
9fmLtSD3elr27Az6YLI83x16tsexBNXLQgQ7QoI146/V3eCBhpGOME1lJ1mFbs1jbD8MA6gSroVW
SVSgrLC0TkwHfnzY1FZW/EYV8J1ddpQZMJXJbY2MWr7tNrCaaVC5rsdiKX5ceatSLFMoBom2bDMp
t7bHPuwaCZO01nkPqvX1BVe4ZEGAH95kIeTPnfC7l85kGV0drLD9HrmX7xPuI/gqKfQtGLnfMeKC
aPlm5PzLPKmaGZboBLorgxWNsgPqGwKFWmiUMXLW61A1r0sQjZLezcIZb3tdU0f0F3iOZR/jMtnw
1c7CZTBxUQfgdOHlqpaJJVOvxjirSv+fW2Pkbz4sXepScNFaS8l23TLTIP1TX39BBkKFbU8QBRCs
ysW3vZ8UHQJVc0pHlk/h5fvQRPBm8hweqxrNsLqSWmjOCUc/VQKiLfZfvBujBx8a2K+q89xUkkxJ
RbcrYQ9WlEjxX/ISxjFH4VtUDWGJ6l32HvyRgq+WkN0ChxpykQLdS3ApB6J2KRXnozbarmxXW12N
ytBLUEieEdUAGL8Lsux/QGlN/kZoUrStHITlf22lW8pELaugQz/GS4r5X8M7tYIVtOa+plZcrtTm
YofU9UpLay99cTwDtqT9zUiWs199aZkku3//DYuQbMQF7xSDzPwNze6nAvJFolvyfyh7Px9ysD8x
dYKl8ypTtBit+042NaaxkNUMlXBov69JdC9zOfU/8cFhd6bXO7RkYwprXzQ9yCx+cEJgERr6j/RA
OKUxn3UPtPAm7APnUWt0z4bBc1cmEUsGX+c3t+ML12JB+kkEAyVhn4/ojzBJA6Dk8WhjjBvdkKWt
T8/n81eN9FJl1uW+TDKcfMXaFAeE19bOH0FE95JENDHu9VfBz27L+byL4d2xph7H/R7RaZXpfEsS
28XZr9NIRuDRBh9Lb5kVXbr5zYCSDxEFoVK1IOMpkY+fyv8dYgDj4H7wna1RvEaAIC153guqqSci
08jdJ17FvN8YrH18k8QikWaUR0S/zAhuuF4930Tx/2LwXcntbpQdD+Vb25gSFAW253Q5yOjPvRA8
+Od5G1YHA+rfQLykD9oOKEhWIofoXhwjwr9yvoUk0AxbOxKSTGN2wRAs6+kkcAs0aYz0Eg1lRWbX
oHJUnYZFrJiaQti6e9RN1p0iKs5DO12kv/PlmyXoTxuDIYJcRyK4/Srhgltd11l1LcYDq2c3ukUG
iO5GQLCy+hrtEN2Ii2UYB2uJtFpzWDBh1LbLjnueY9pWGVPFavmnEq1LpybBr0jS9GZrGkgtngdx
So9fpSByT+6fHj57INFmlRDRTGCvGcx6Qs3nRqWU9UDEXpn0BK0tdY5xiVISQbphxLlxrWIWNEfc
V0KC2Xfk8/D4JlngMjELhS4ujCTb0GQDs/3pySfzYoh3bjKkJFWVlsEvL0ZegOafI16KrDek2VV5
u/JGJAEAbc6JG6XPnEYlI4GNfFWpUMsswSk1tfV78ObhOaq4wAgrgr66KHrSEkqgdmXcaDpBhjJI
pCZRP7D8UY57RC+WNk4iwnVjNWYZsteEzzVCeWnxvp7ql6z3NXng7xjYh8vXjAIiV58xjtnf1ohj
UXGdQjX12Flgwh6Uz1KXqv/pnqmHZIn1oJEhXkogqK/OiTIrnqQxE/5UbpOSRL/uDjkTMtdXfgt4
X0roX6aojBBkU7n5s1Qfi1i21pt9jwUKPLONi3mCqN42eZD3ORZnvsn3P0B2EOzuUcZ/FxYd5LNT
fNVVUVFYVUFl6qnLZ9kp+UrJNSWqIYoRM6VdX/kTQa/7g8p4tuI8s9qJBM+wHbegDYrJwwJQLHeM
fIpDyYQVb57+QS6CaR7EnLG0f7zOxR4fMyPPkhwv6o6xGZkI+huZ+6Rhiw0OpE7BtfQ2/VTau83O
qH3F66u4MV6LrQakB4iytpd9nU/JBfq59DsdNBeOh3phrM3/QBMxnWx9umlWOL1p1axhdSIawsVj
9oTWJOqlqm9GZA/+YY1WE6rPURVRxLSaeNG4cl6X1OkZp1vfzjnXPjaZAjpGp7x+/oQu5Batgzsc
plBNqWKJ65s5HH/e6sbsihgLrDD7+aVKmcvYajgAZYdG95BX9LiCkupdOIwDW7G29HgZqPafBTUj
jJkDiLBIN2pkub5O0r5XXeWTDuF4eFfJ+yoQ20EoJDpF9AUlBdINWvdrrd/7gBkIXGUZgygDX6kl
KdvsKFAw3N48/4AuEm7xnJlH9TeTR7sv2+Psmy5//zfaFEMBvRHVTlT6z1/dgzCq6w1Zkm43UmJk
p2miK7Bp81XzxXb7AEZSRV6goPo+ofIh70xKtPkC3wln4i/N6mTOfXyfqn2TTQDZ9pxWsn0brXoq
YQAivuGxdppijWeRTc0sSKJqFs+j4GJanQh3p6HH9U2ZameCi9HiD0oHgy+gHLGcJ+8Evu1lwK2V
orXbGLOmZHVtrhhZijWHpZLAHEcDfiX7ftEKOBzAeWppHE3kM1/mrLvMgLST98WFsOl3PwX1qAHp
3Jrgs2cidniD634w/w2VsIgVaB7VDBiWANzCjgysTMmoqJXjF+v5AkWUL8dsPhTLRfuGP2F9Hat1
zUvsirOmDC4uBnTEk+UotCts0U6TywOh1DylYDLjFE9KGOK7ttE5BVBtINj5vOZxpjeGEBOkUyZQ
ttBVxfy5KpKUYpLzDDhR5cU3wTITN54UA/FpvLUdLO8yapWcUOY1ln8DsrYGvnU3xGBmtJxsKnlx
c6UPA3RR97MpZDoMcK55taTW92vPvhGcBk+InwVAyrDMmbwmFStCD/eF39ipCBybAoOTcYUAmTdr
wkyIImczAs5vBYu3Fu3g0sMDXfZUYPw94sPCzCEUU3NPpCBdhJ6UlQSJtgB99ALZvAEy4OjHLxZt
phI1g/pzSxdwVoec8yw4L/6qJNtZBaMUZAc8imvH3lOR+MT8EPQ7E5d5J+myPbfqPKfdbzV76sEx
UO6qPf2ZmFHS7nQ8h50uSb8cCMRpnMqdisInDad19jJlTviXc1+fh8FR1CHimey9/+cU6G2BcHyi
XdYjR+xHoMqLZf28fhZa4IOsMRY/X9o2e2Q3YAqdfIlb8d+ruwwIps7qQUjjURRI0DcGMmEkQOQx
0hoGr2jYh358uMIEaqXc0NOxxTvxU0j36CiA8wILc1sUdrgW0EHDQ2eNp/bsulJ7t+n5Uw7HNXqD
SAreT/HcH0av3hjgLGaH/r8Oz3WMtcpBE1mdLZ+bBn3KpJgKyWKhN7NR5bxIJYG0eySJv61C69nG
7RKDgEcYVxriQf5qpwBKcedyA/L89/tLyoXxpJqrx0zPWYMGVckPAWIuztWQuK3/LU76aMnSZobc
zzhZ4BXsmfihCpm0wDdNf2NWum0D/LHDcOH3BGvFh3LN91EvtI5UbUCDzKcGF7mXjA8kztyyFxrR
CRxgP8d+3Qhm/W+oeRDR0V1rb1rr0Vmpmm6kiZ6qHysiWM0H3K3B7VATotUPywvu2zRo76XnNDcb
C+xPxhgRam00zZstY8shka4k8bsnPn9c4wiFBuAqRpKUjMjzAKpmjRZRyQ4jgDOZpwHTBN/kY1+7
4po/KxIVQOF8PL09wjG+QrQkIw/bBBvjPLEnWPQppeO/hgeSRZX2Z3HqmNiAZ5k7VVDARsSkkFH6
kGXQy+tp7uKCtfyi1a2UmqMWxZISEHlSofy11P/151E+CPI0vS+Y6VAkF6EmVLLeSmNBgEeI50Ma
s9fF+cbaq88/SNBJUZSC8MijN/s9b5cHtMCJ2w7aZWavjoP7H8HRjE1onxcTKwAShLNQ3QpcycwW
aXxTEqNIYCvW8Xg//RpqhEmlu1vh0teuueBv3QkN5qKF6UHZVL4Crj5il+JwxL6Tkw5laWBy8Dk9
h9ABEBLJdgxA90DGInrG6WyMIrwk7Eq4XyvSd0EbLGB14nc2sv9SbelMcKLMKjnTKWFhhnLGhe1y
fbVGUFchjEZ73E1B2Jjuh+cRaynBz4fZEwVRiDdfrhLqV6E5frFNVnmmL8aH9Mj7k57I2SGvt+rN
fijNln24w+QxAeGOvtfFF5g/r5GDtJnSsSpXY1NORH3qQbZZB2S534ODqwacgXDA2y3jF2tqrbJk
MKTLXJXOO55J7FCJJfkSSfbvII7X5eUPoBu2OYVRWmnd1zRaO5gxeGT5QSXHXjC+yvVpUlizqB9Y
DPEAc4vhAtM1yPKG96puWvIiZ8rqYntNpwEKRvFehHxSX0ipdL1SHvQiWj3ErldYLVeBjYcRDUOI
nW0omJr8QxmzVcQnvfxynyOnVPaQF4/jV3kqYSxuHssmgCHfrfoPGkTktbYvzYLt97rYiR4ddlPL
UVpzk5ETj26d/WsxGzhvs9byAMimfLJyChI+Sv8rX6g4BJ1tfqYXN2OqG3AExVrYoNKD6TxymeLR
PIF+aEtpomD0QSnOROa17uQ4Jme7ekQGldVMgdjJG1Co8UT6Wb2nkuEK61lhCzB6uyepEBhE9j6t
BZT6ak++otAblBOm1UgUI2bcWTfKSTaSvweQoyQq/MLiuUwyx+4fIQbq/EQP08V557HJZ4BpcndX
YjEwsKJthJGf/PyPDX8BEygD+m7BECwVP31Kntq+EOX2zRgCL+qdgY8tqHw6nvETVvMb2hM2uDpx
t8AKCz63vk0XK6CdYyZc0N6tRLDVthVtJktNE6Qx3WAZEvvn+u8OKBA6kTG3oKBkyy8tSmBLoQxF
s0JuUH2wBRceTdfbILdLH3FpZp6182zbKIVzpAkfEc2RWoDYWXKpNX3Nx8qPQs1bjRpJtiflpGfh
wVpR6e/zz6qt2IQJqI68qefUGUEL95tLdLyjolx23ptsnSi9ndjqKRGZi9OBQxJtTR7KxrXPfKQ2
kdqkhap80yfWv+w3w2mdAygCQg0MVKTt0OamvOWprRqeB80xetcyj1ImYaM+pHJxDSDRe1khGTZf
DB0QoOV7MUpAqaDUDLyUqSyqQeYcclV0+19w20Kbl3/ToAcxOrcAhc3XNzcPhBGOIkuw8+xV6aMS
3L2Aa/V571KX3ztPFslJ55pd/V6C8w/Lu/4HXhidnAWoJnN/U09+DyXjTwWgmpT6bY5cAYGW6CRE
/Z97ssCOPRfdXQTbv0kq8618Fs1lnaFQPFX7sYSv2NlUXhCeVvAdn3owA80stIwb/yhcTbVTaA02
PBfMR0AG+JZzNCojse+jKOvBlwP356H3G6qOpbf6BdozmPdQX3kIy2rWhcgu/X2x3Ku2XimPesSu
VopKFLbvpfsVpnktTJ8SKTRZ1ZmsTgKkbI1qziMYU9VF3lPsyC/G7PxXK+99PmGU0+ejjrIYyPE7
Fv/z3CUhTSa5BfdpsbfNedbirBdjY2WMGpCvc2p10rm6HbYeWDv6dHQIW7toA8N4hAxIytbY63tf
pz/rjrCw/l3uCrMEv3KLIpcIOrfFhqSZfYhTOS1RWOJS7v+kp0AD+3ilCW944nxyfNPm9VvLOaKh
L/tyEbgl6p/F012uVzyFzVmhQP6zhp5VKaqdguQCSCW1+QmG9pISmjRAZVCD0fPszud81LIuKPmU
qtuCFEwp02BM6uOQJ6alORD1TSok+uxS/IGM3Tg/SN+XUqfr/yWo560NEFaXYayUNonR8L5YrrWc
RWAW1gup5SgmDksZo1SoSoCqVZk6bwLq+YmJkhbR9KNxDil2EQoglPdIKZNGD772tpf/+Tfl2i4H
iyw3azRHt+e/pK0/X+oQKyD/tT80ovjBXvWxwTElxPDRxpH2yFqSu3+lRaVur2qdzFD2eyDA2aEC
gtR7a/rqF7dXDe2+wungYgtCYe0U7ssvAVPZUMMRRX103bj+381BiKqmaXi9OGCDp4Oa28SYqn8K
kT8PBO8bHc4ciVdXjTNESJfx58nFclhnThP7GRfW4iXyD6SF2o5WZ9+2bo19FEg2Dc1E6tdhhL+T
sbOaljhcKss1IQBiMVvh2Wh4LbAPr22SMDPcchHRR2PD6Zad8PCBgrHQ2QNnhXCR0u2xhgADF6bG
9vBQurHumOD5PTJSwpPGzt+SGqfLf/TW4/Igltwz3kR8y/uB0/+7KwCCgxmii/agCwv4Ua1kwcq7
ayDkKgIc8nuFvvj3qVecETujIeYmph4RNol2VzQfiU3sLVzd+9RDF+rUSVyf56FQ/u0BCociC5pz
NzEOA63Rjdff1rdxaXvi/oJx+qkXbbfYngd6CP93Re12UIV6gHG96f/i8JNBIE7N9ErQpUr02R6G
kG8ZV8XFkByG9cCC+WaVTz2THzzQpptSQRzilvFOkFvuERshQZ3Et09k0pjwUa/QkyIxiJ1y1UTK
KFOZsAg73jigLGgCbvpcjiP2cs9KVfAjutjK4Ai/ijKXqUajCVhsX1Kno7Ta/bF4ywMIGKX8n/22
v+ciZQOdUDRCRtIW8vYWKsq1mCRDXRxaMCSwaDyEQ+Ie+dcXKeWa3bJjGEtNa2LO3aZpO0pm5E1a
5GzkvYxIDe8vN96ip+ytzNil1DLo2R1vaRNGKSag5WH8v0HV9Wu8b5itYGbzTFX86pjfNeiiovc6
vAmS6sgDqTZlUpgPpHwRwl9kGo54Mceu5v/4tjT/HxjlDFuemQgyDRT8MQKCFXgLZwBFyDy0ZPtX
IjM6SUSGv3QEKWiJd+Fbwz7b2JM1EZvlAW18tEosqk2WTMkC86OnccdQdGNFEAMgXKXHr+b7gGfc
jHskXoSOzx8tSDxROKrlWa1fY/SR8YGn/xN4RjPlozQDUlYpMapYgULCWPw+ztxtc7R4tM24yr75
jOeoQa39ovY1K3ky9qBxG9/8hkWE0yltD3k3cOy09eLd5A6e0cyTUDfKzJwK+UYJ/yzTaXM4Zt72
SH4CFzsdp4oyk7lw02H6l7AAc6kTAOoLNwUKwI9qwSykr9BIHCycGcFkNluuuyl9LeIPbJ+gq5Mg
ox1funoPAE4JWAPIn5x3HICVAZ0LoSmzaMSYYEy503rzHPfgeoTWgLUAPgoCKLbzb4m76SoiAiGK
lU5yXdpRdTzu3K1wXVdmE5QgRqaMBwRbiB3gDkQW489O2HB8ResKMwCLkunYfi6YNtIAm0+UY7UP
SDeGWPqJQttI5MpITT3CvBslvfVAIlCgsLt9EukPOAoCzmPXs7nx39v7eIXQmj03ySi7YFZw+jWg
5JWeg0szYFtl6fN6lhf89qpFG6osA5+cXUezsoQY0QrFp2RGvg1zALSEd370e1YXJSExf/lkPjH/
N3I6s3hrefiNZQXvuTVcseiDnCgodKg5Z+YpeA281noA3ihkNpGD26wnbGUZPYAV2JDwLeNUN23+
orTvgQsYjXwaKVYx+Z0983QhNDJHOii7pirH5DcMAWlX0GB/GwbFGb63uCfdjRXjSD36Zv9vzdkN
Z3nfEiRQwxbXdjBIVgHciLDwdho3hXfWs3vrAKj+fwDebXapTBJGn8zDaX1/MQFDSufkYxYqfKcS
PcyPq1G+Pcpe/Gwyzfi+7NsupvFtH0r3Otrkc6pBLKcYxpwkMrVhR3uC7hgBT6eY7LMFChwB6RNo
5X6VyAO6U3mDSJtKNJGmrRgqisJ3u0Oc8sCH1tnKa2jcAb77KLHWDVjRn3nGcXpiU2/G0GS4m42C
JBmE5Nip3oisk/GpzHUjFyr8tZOWy3KQe7xe2HIvLEegpaHNGxzsz36dL0G2tGJYB+cSxulEC4Yj
9FXiG2aBy96e6KuNYEpmg54CdHOlHXiVKoAAadrummZNRK3nlRaVmVu8F3gsarI3c8QUkDYXegf6
usmFIFKyZdFqeSCxfPglSCQLkDN7DkiABZK1CuQk3trfTME63Jchb5wHXCq2ATNNFTEwnO+kzdsD
a2LwUjMK2Vj9/W/FrfebPUj6g9mQLsUJUq5xFR6qwRReKuMIffarV0hnTs1RSRD9DjxE5eNpjMej
2O2oDvEC7TO307gLFVJwfPuQFcShUSvRDMxi41FLd5+hVz+6Psu5UxoO2lQK9xsalDDcBJVq9U47
pnY3kvaSYSQOYmNb0EaOzQwq55GvSylne1Eg8azp3DhgwfZbxbGDD5J6pg7M68T9haqjF8iKdy8/
vJ+BO9SeFTajpIzYYZs9s+hgxajjFBo1BTnB3F/InnhjASoRLpLoZWrfloTPN1hwIrhcJ4S+lPgA
XknUUIxevlf4mYrGQ8KSGuTXYWzYDhtdYRxBHKtW8ospMLNxsnANIDh3pRyedEDfrykcmIV+o9s4
+LMG8B5P9avG2Dya6gV/YDGwuvTVEDjoMyPG/jpTGUUYhh+HjoqkaPsXgCj75IRYJT44vTPbGvGQ
bWVizwIA8aeFSxjHF7IS851rUFenP0Q1VHu8ZIccHdNCb6wsUKa7NB5zboGNq5/FRXYD91Ner5FR
VF2WZNcmSjJ6JtTobkWs0BrJkVKJN5enlr+wimFfWf/zaacBtKG0o8SzbaYZVBy4nW6+K25kv4fE
GQuS9LKCXxCk7+/QpOwyDhPNe0XsrQ5LcbnySlQDl8OWln6AUNeuU8Gx2d043eLUrWZ7kirwLdO2
yf5WaxAarYZjiU29jBzx49ZutZf8gbKFrrPbFwaIGUt9d5x/F8ojIM5R/6UkZi79wRdJSlOe2FSW
BFl6Jso1SsbpwWEWVYBSvA66wqO3S08wDU8gfNJT29GK8jZwO3bmoMsIcnGoJ8hJcRL5V5B2/Gjf
F5s7M/v/kn5yqfvwFIrGopsNwia0nFbDEcYt+rFWWj8slHQ6vEGOLfRwpgK69F9z1vEgljyUie6s
kXgeKVllelVw9e+2NmRQvPVHRlXVsnH3XVUtnNqTzvTdFXuC+ssE7VoSVo1NBq0A9HP6Y4gXEnfO
5esiRPkUXxOR4W8T9iImfVIQ0T2hRj2ww+zxM03kVWKiH9sY4o/Mv5h9MOl4Fuc9diruqTfCNmOP
qwThDW28HNqCPCf6LkAAAlbEABP4kcwjTkrlUZs4uACc2xm6SpqEGbwjkDJ6T8CcEuX7kSSbOrNd
FoR/pA/78ZqdEkjFn6AMUQgSOdYB+2SHzFfsuTLEb95VmBVnWpO3wEb5Vv0MSaqRIoi87m770iQj
bwl0RjX9XsHjRkNrw93VebssNBQvnPUX9+VjrHSfXOeeYeFjMGLlqPtwDriP6gkbwl4xTytJ5W0y
zbSAS5VrlSVeAks9Qspgn2KqrSjWa1hBtQkFU1dhpaLi83XnQ0MJ+K2KqgpOfwso8Q2eNKpvQmuM
FEjwb44xNLo1fhdyHJpxW4Pd/Hmm1/9n9vy7BtPq0ItxqyBPnXfFcY9niXXaSMxpBLZvgQ7Wxmqm
bEgNnqjXepbIROZusIKM1hw4LTVqfhZkPDrw43bIMPrtbr1vY5v5HfSmeANwRwPHTqUxnbhugsup
yzkial0NEfpFoK7jCke4fFtlC+9svAphG66nBFH3YcJwC3wCIi9f3rI/BTQA3v1QixFK0XqDGDtW
2yKPOv0I8aZ6pHyhNQdDitaYTDQ81v7uj8mZUtDsRwaDjpkFVCWK4yWTjY1mGT98jXU2CjQFZZY+
+uys7Rjaf62wDSg4lkAMPPPmaJUD7ItvKZnRtTr9jddf50OVmjvxnoY64xHWqSJJkzJw6P3mRtC4
owUCn1W4UGB5mISx55Z2nzoWgKO7pbpR3nutLRKqP1h5rbHqTBpM1K04fPfDAUheG2pWbEj6VsLM
XndgdpO9KLC48TMGlwlmoNdJRmxUDh2Te9UoqKgJowz1LgITkTiNG9gpEBzK0wXtlW4TMds4OFoV
tRzwj/t7DdxkOEPI5uLRLmBL9Eus8Z64dr33e3WbGkPdB5Ga/mlOKfd1j0ZgG42KO01vggylNHfd
OFgUZiE8++HxLFpBvcHFRndCc9dDs9+JzzC3qVkttRuCltYU9fJmmgwBuqqvzjHsonSJ4/FSrRLK
Z1cjHgtXmTpDaddAZv/0KKyh0uMpgp4RE3buAWo4UKf0bdy1MPXIQk0phrcIheNJc1pKTbbpuRsG
/k/xlmCDHxjLIh/UpdKZRH0YWlQvOUtRxeF9xO/YXm7i4Y7CVwFcmUOv+qlCQrdqmmUtD7nauRVl
BoxIow3KWEk9OfZCZWq0CKt4II1qqk233WSkXDxqDW1ybbBYiGK2mEWKURk+CM0l/63u5i1PyuJY
uy3++HUJP7ErMvCOvg91g9ZK3YOZYZs1j1vqFAoa36kwJ2Hxlj1fIEcOSZX+Peea8o/kYcNqG2q8
CJZkkWiug4YNWtumQfoA3ZqXsk/lJQ+eZNNgWPy1C2kWRLZfzw51BRjmxu8YXEpvobmjluRu/b3G
NuXZ2lDsnkZWvCWqWueYZs8WPFT/qkKc0x8yIKhEhQXJ3kCDh5uxzZTjdSPAO5TS6hv56tqMFRVY
zT9l6g04gmH2BA+OoR7pa3cjElzG2vuU7BaZ8SbXLE93QSde5LHis6U8QHvo3SbYO6GPbsb5udtO
BIcGe5dh431phxmYxFwW5FCBxl6oXVbJalfPbVzPa11CDjD8byharc8sfXV+ypaBrBJ1KmdNgBCz
22tMZz4HS2ylsoAVSyjuPPEO2BVC1sLQtpyra/4Zoiimjmdq/BQOlDv85i3oMsFoKA5jsUyg61H5
GISECaP+McCn0M878+dhbX0X50U36GWtt9r1l7UlF/m0lCD2+81CjQl91J79nRYMSRrx/3rVdj7Q
H9oeMquu5b+BRPRhgV4FmjrISlryzw7cdLUvyE1H8dMaK0OW3wAJ++QuE/eCgfA1KnnRCqBadOKO
xDkc+GuvNlHbsUG7ky7gXUWUrUEocnP3XBMrZJJjapkrjCVutxE1j31UGLi5RKbH/Sg9+XqlEfvb
c/KX/2w+7CZy/cO6nFkcac72rRTQkjAnA/WhmnK9y+ctyTnAysDII3N32WwiUtNwds/4rgLIarvj
UuLq1LgCTFeJH5hTIJa4cyf7AMPhYF4HIn1/c3Ival/N5kaTx4KSCtgTj4OStX4tJfFav7Lz1qjF
e053bw29qxidBppR8+6tJ+sxE2wlZDR9/KZQE+LYF+qbFxmGM3pyWCtTLGDQt40nGcrfRf6a+X6k
vARWTQShZoKMWh/JQOachBuAR5PGU0gG2fIfGB8S0cDRsWAq4RcdMVBXD+Ppra3Y1MKY1XNwKJOZ
Vmo0eEqvXh2J0WOiUnJ6tGOVvUX12jKmJO9nqedrdYOfaT+a8YkRxp0FPFe3qeuGij6IAHE3bulV
BYuXxbBHVPgb6RhRw69LJFfyHe3dDOHnqfUN3uHLedTzvwSrIp1cL5igmsnS05WBTMpslDvF08zq
2SD7TPMvyiKvFYv6+0r2H+ua+IEUC5+ofl3jQ9iXLtrE+ANyVrZcrZ6OG1zrdXioeJI8hQnMQYh6
/gAANDKpG2RF3QitYbQT2zPjspHRtIh70PJjrk1aRdSLKxnv69o9t/8jaqF1tCfEM1td64hDrC36
iWNNasCfXgsJyTfcAQ2vDlPP6gA/IBaGPV21O0+2MJg/ytKOMQk5rm3pw/XVuIz2UuTU2IJLVhpZ
eIPCjakEczlxyGhwoF45n8tccYSikQWnkZIvXjlVhRvxAfmuakfoIMj0sLikIlfl6fj7ApUrANGT
nDtVv3FiCFgvnJ2eUvO++gw6nYrMqFS0NnH3C6GiFwtDDtuBdHhl0Rv5IogbwPE9D16U1vTpsIrB
meNC+/vWmmYZRl86g0U76jRpPAyYtmeAJuplZV/sLPXCJgDm4t3aD+P49GV2ui+kUt0OR1fGXJC2
Rz1NhzBV/BsVTk8FxcbQ32hP7ZUpnOlU2npFon9h9UB8LM7s2ihhkuXkGLC0y01u9PBMQWduAcyo
uNdTsSTVkeK3JPDDYy/0Vv7ryq3iS2ZRvqAkKYu3idqflhBe3McdPFstARAxfvFSbxxllwbowaFC
sP1dJ5AP59HVHp0RZ4V+JY9gVrC2QBGPi48i4rFclFoOoCj56BC1eblLH4mP4j+1Ti2mw5lh1wm4
OgQvoNnedkpRMV1pQ5Ge/+25lqNk/t8BPNy249xKuygu/LqQWqxTUjE+YBpb9vSbPBdu4/6CunQJ
1oNJdXWcQCFtdceJKBgvrhUC6DLfCQb9ISjOfo/LtJctgzcsS3OynRi6vKMAO/t/cmt++FMM7Kpc
nYQ/oYuWgni+ehohW+HFCM3VREB0zOM5OELdrvmLiwDWgxwnVzEDju8gpksHjRI/M1MdqJb4v6Vn
fnNRZfy++B1krxprUQATUhnRlDaWAsiSOfJzlRQnXf9dLv2la1iyU6iTyQc3D6Cw3eUihf2GJ4Zc
GgHV6wmPbPqi3fts8Xx2Yy4Y9c+p3CJ4lBIzB8z3zhlpfEDmhc/3p4Tfd6T9tiDdQYkTxexWj+dZ
i2CcktTa8c7RWk3TB9En27n00jVdhZqPh+hZO8g5t/daG0kTXmRRYoQ4h0DbMV1PrD0zAMRgNSu0
L8ovwUmP6tLIMgAr28QWhCkDGbj4tNgamSMT0rJrQAiw9VnFmcKp16KzM4Tx9ixln8sOf9YyrevS
tVbuGGDJaA0FN8I/ontjRCPQsoKX1mndQ5cJ/Fl7BbQwlLToSIOBnIBCmFs1RfHBVJhUKM3neKoY
NIkNWzrfAt5En6N8vnM8jEH3x9M2PeKbZ/dVbYCaEi05pUej37WekKxd5w8SpQcspschpHkO7K/a
49KyO1ytZM1inUSjL3aHYJZs3LoCpvU8WTQRfyyTb4em+zUxqlBxL4Q70/cD+P30I9uXGJCmw5BH
HnlMJOULI5m2o0rFJj7h8nPJwnc2AoujpKruqsL+nvX2TDN70ijR1rTdEgKa9KWkwShBSwi/ULG4
X6WyWplK0zGZ08LpsWE8Zu1hEm7U851WzOE/gg7DHrphfHE0dDh2gkmoe4zl3g9c3fasUKJ33t+d
1RjzbkdbjQhyK7sRdvRGKqJvIPmnI+NO56npuxf1g2s/N2Na9v9qsM0kcYX6BUqrxvRIsL0Iti/8
9qql1BXwAiECR5GQ9wNGspuHyL16G7rNfzivI8KbymssNLInRVb3ZhuS2gKx76gSgt52+kbwX9fw
YeUD/waqI96wBfSOaUiktc1ZhFkehWe+u3Np7eIC/yecZof3xIPNNYqj1jTMpa3NlZmQv5WlQohO
788LuL6iop+6PLPF9TT8Bp5PzA1lhmVlciieueA1KynCsllaIxIFjyl44GAuvzthR0zlkEaggD+T
C/2jwf1Vu4PNLoycMI8elRi0Mg85XZJnFo+/C0sNp0Nf28P/1jlnHXnLU2k93OyR3cd4Y3seTMOo
rA9IFRN5tqnRBHnEvl8PJuV5MP1ERcI5u2ZaUNhWlKOljaeWwFC9rIZ/T7KTaDl8yr8YWXej8fdn
esr53iYo1+HcrRKW0IpxIfeo9XAGgwEY4LqRIzeEWuFTnnLEWyqBRv64gvjh+f08fDpoBZMSu4LO
FeL+3b0Mt3CPTeQkqRRZPdkaOFXEwm4Ric3V2+Yy4DbTpFd/GAEn8wjqgbstuycMett22i1ZppIf
NH5ATHMQgtuPZTSDhdoU5aI3/ElQyAYJztxex/KmwRIROssrz3XAuEODY9XVzvURmpdFNCPlQOFm
dy5D4wzkGuKuDN8xyTA6obhH5m2x4wttIA9hFiVS5bs9BlXiXsutDMRSEHu0HqkG6R/TRc+C0h3c
7KJ0FfQ4pMhlycb/L+7H0GtGmm5WcGysefrMjS38ZLiTEEz6+UWQn617UY3qyZ793/y8Cd2ItPb2
HyGbNWi15fHdjQvz0QLB97AGcXXgWncu5QpNNxgM4Z4UYw78sD7z2pUZbvVvtrfnoBrQoYTChvFk
rXHByLrIYfEylDLwl5AIotsQv4JwjZ5zknW67lF8Sbk7ZHOZLdRzKfdN4ExkvUJtqTeerIVHIzZ9
0L3SD2xOVecOCz27z3uQqhU0fa/6KuUBfsph4ZJcyaeyo1LXasFLz1BNV8pt/uUsn8/PGU92EwgY
qTAUTEduiPRGVKMxmxc6PHB0HwIEYADLGIhO2fYm4sFfkKqi5HuKpV1/oxSuaa1vSLKQjLgQZ917
73mods3nGpp3kCZTy/Ocaw9cIwTGOa19ioyBsnUTrpM14YxaeOprsnij0yENxtFgVFjgaFeUQGd2
0Ruewv5Yqrph7omyc+jnpOEFb7B8Tvo+Ulc8eC/1R/PakzloSMTuBzuXqWqBaMCr1kR0OBVYMj8M
rPYiv9lzY67iFlBpOY56LiZDi7IBSmp393xpUr3KqZeUgDUTuQJ7Zv/W6riVhA9dpqHYnFI7kKTa
99SZREngYZqHh46/eWp5DjjMvCiZZwgJd/zwmLXWc9PEInenhRSR5qDndkGn2mDQ4OIfFRv0iKGo
xATGIyYm6lV+2K3UjeRSIPYjfwv9utB5xiOBn6Yl30rdQmgK204p+MuQvMZ+uy1ktKfy/o9sztPz
tBM+aJKqCgYs+JaR8DHraVsApaz6FCJK9eViDuKzd6ztHvT1EK1kLy44yDrXADajS74iusd12Gmk
HCwmmdH82VIoCkNAqTBevXuApYrlK63TitY76eYzkXhJAJoIQAzhHZrkjLZh3emssVH7Gh+paAIb
bYLTZDiO01MTL+CKMKAR4FJD0UTo8oNUJODZSRNj4UqPQmEEsiYjZtbgQ7ndfATCs3A5qW01KXv3
bID4FqRwKSNlsye6xzpC8j/xaabT89fZN6NKajAOjmNiTaUnm6wybHcBmll0TJaFBRddpEAIkOvN
ukftEWg3tKGIbbkuK8EnGRzq7Up5AxGz2CS54nbWi38y/xiU/SvyQOAr3uRGAkaCKEvS0nFnmbhq
TOrWGLE7cB40GzQ26CmDMyZPOaeUFIiSc4dtRXEcAavBJsPmpN4bvXt3tpIhtmMgGMMxswXGVJL3
ZWP9Tj1bhiY4v32RR0PdsGoVuPrS+ppHWvwHFnKRyE0fw7d2L3zykbDLXTsknoVejKgc1A6NP15g
p2KpZhnEojkFglbtaKEBJ5PfMXqHMT8bHMChVdF+vWX7w67KpgWuUgBbNNF+PkV8yiyq9xx9nfrb
vabbcip/1qmBnqBPkAcnR/IdFr6gjgMgQqRBuvGnuvAknMDtrRmh6ii2Zp1SHgu830TqVmSF5kyo
91KIRIvWQTIsayFNgHRrfYG3kNEEPcZmFTc4Q036ESICmrviH9K423G8C6tLNndBE/mLknAC2tDC
Nx/mgiCtPoS+jwmHLDKF+Txz30elFko/5sLx8c+xltVuBg8sW/8L+XJ5+qB6ldoB+qtoVatirw+0
gxqfUGiKoRjJHmI+O4UvmmAtPbuvcIop2B21lo1pVlTfL/IA0sOU1MIT4foTOqIJ00k0LvUqN9bQ
qqicjq325VWE8YpZl7R7BECzL5sPkNqLqWN7Jvt3eJjbwNibJYn/EgME1fWtsQgoRnbcHGmT3Kbp
Gde3R9NQ2EmYvY2pZj5cxA6qVUreeO0m3XUqcls1X13aPg2oW4kVcu4SESQHTGaLv9Bnv0Jxkqpk
DKhkd2PrhdoX5kM0gZVqfNRnmjOwUtjOW/UvyVt7F/OcLdUs7oWn+QFvoRH7aAf0O2g4k5jXctVg
c7a3qeJFwiEsTy8MSs3qpWcAa5QVVI6xut2HuHs5Vzm87HcsDVmlYcmCGGLFp5inB+8ZyvvTl7r6
qHwvJk/u+jkc9kzAWP0VOnQhHX8Kj7TlZTF5gWbAMtDBw1DBVPPvVS20sJTf1VZInSCeCBMWTL50
vEM/JgPKYSXDmwHgMj+BC2Vlgcl2uZqsU827Dki4FWWnePlXB2v5WEGfYkPhsCmTxavq/PokyHxg
xNaLfBHEwjKLrNaUTmnNMoH+33N9UGH5nKl7Gk7ioHzutDwJP3dyTjofxXOxkc8i+4j+mfgIjhd5
qF1MqkSwzm8AjfcI04LhTN50cH7JjepQc64MBTY2cKFGTzvhhf/oNrTirqc4AiYj9RW3YnMTV/24
xxRgpGCX/tXDyG+oSytlWUGWxYhJI1viRJtcYyyTqwfzdetOyJkqQS3FeJ+lFgAZMjJJKVWxrcBE
2NL8jsZZ/jKyMUBJ0WqEkRsLi+lrtmKdFl6dP2bNVPDz/BohRv5GpNtSnJxRRVgX6ZN3fKx+yxoP
x46KI+Jpa3x4R8eSCRCsWh2i5IFf389sC0/Pve51jFPnLJIFRC/yVtDqCYL0UdX6eQk4E1MMMWeW
mmNhllSLQ0DHU0B3vj+Yni0LmIWSYyfuLXhs73qR5QRBBkOvfQb34iT4afr6IBYlv0HIuKAl4+PO
xLkPWsET2F6ZShmcoth0z9JFVygm4PcJt69hMPtGb0XWkdaCs3Gs/7S/PLtClh2skj9YxQpqSKzF
p+CRF05tcJcc6zPD7+nuXi35C1r6BLZofxY0WEf9Xw+yitjirrxwN1/DtaSeKqZ6qUQZYlICqSCH
V6bQJtKkJ0RpNHNEXZ7H8/YUyxwIQb0r5noL+513GmGmf+bqRlj9lCoFNggH8B+XNIlzbFT3FSin
MY2Bmrpk+adziIJ8GoAVqFt+nYfrXZAbXap2mnXQOCntJV4680DC9kBOPYQ/GT1WWCH2+sifGTQ1
EgG2Iwjq/Ra6/vCJGvS1EZetY19LuV8AixGBkMGDNpcN4bn/VJoCAA4ukii+17eJX6SZZBfIBJyA
TJrV998uMkUQ46FJciryNGYQdmPZhtJycJY69LNlWtAdCNJ9PFkEEKNXZZJyScG9TmpK5aZptNTI
Boy2T7O3QnlIn+wuUn627FLJXa3xlyDcCcQyYcIAY+4DD+TxwjRu+7NSgLjAInjXsysIqZDud6Pk
06OV0ghpgE6sbXFiVFMw/7X8azeJUeKJMPWSlMGcN0PfQdyqjUXEaCYn/GJa/QHalvvwm6g2rrug
YExuISQlHP5xukhxzJdxCoPm7LX/rYAgBdWATRkcG50puiPkXrF4d//JhspEswA04qqVEm7lxLo+
SKJCPYbDN5zP7Dw7f0/ksltlwLYd+IUPcDpRO5grWlVIerNnvfPgrj+8ZLjWXTzTRFNubwcMLOow
TC+7BMxok4l3Ea/1Xt2WtFh8u+2KLYw+hmBVXVGTanDfFN9pS5NtteofgoELX1HXl72ybicl0DlZ
XNAnwNezdMV2tpoNKpaiEAqSbJWZZyYN9I7sZnfDadclcc+HrP3bKK+1DFgliIp3zfdYPT8q04KK
V7pLgb66rq/vTNUGp7ib9aNJY+2LsHKjIht9dH2nFwTOPKT77VubnzGlv8bkHx/t4S2eGiq684Q2
GAm0ndHj2n6SH/vC0XCnrrRwQ1gNDMy+f3n2zRRXre84iugU8YQERlg6tbw7TIeuk0Bk7FpeSLbT
ZnGKUUqIaX3/ULAoxFbFYIyKd/wzNHzuC5xXTEdiUfegKTkqzo3jTwYG6BTrcTrfUN4XdTqnMY7H
QfJORLb1o9c2TcpBPUgTRy/rTp8i5Na0bSTvv5NE9zbND1wGjHeUEAx7y7keSGK4W9XvL54pHeVu
GH4coeCA1u86geiOwjhcqhzFoY0oBCdt65OwOhv+BV51spW8KP/HDjPAQjvw63HFcayKtQ3L6QQl
xEXeAp3LY7Fadn24Y8R2TJRVrc5q6Ats4uy5GemZzm3IK65ww+SiFPzzZLkzz/LNgggv4v4DNrGE
KichN+av4GYq9FVR2hPdNKxigG5Ol3kmS6FE4TVFaiEVUIVjWDrxPMvofnWPwUiPbHWGIApsRKYo
U5NBCENNxfffpGVzCYkkxInWZbwyKG1pJuSbTtZipLi90z9mMbVBuN3dg58lgO1yaRN8qYlo1OYW
CQARdodb41nEvoURT6EqJfjCH/91Ez7uidVdKiY1NMJLLTRmqg058r8KyTlUq0HSE4QWlmJIE13S
BKDknT7ufMtBVTy1cHpfX4oKJ2+g1e5TmpcNiA81zsjdD6bsNomZwu4qlLAGsY7BqH3ubVPIbo/W
u3Y42f2rAmVJfGs1b3AZB+whlSMRT174JOFsdwpIoVfqFE3kqCxlemrrn1PweJb31fk/rd/zzt9A
pUSCx27vEW7THfGCYmEmW7Sg7jz7V5kiicFQqb/4EYRXOA3JRE19VSj7l0A8Z4xg6PaTWREAF9o1
m2a3Wsoaj+vSIIfy0VZAhgQR9Tnc0kkIV54JX39ov3BgWfg0fTAd4hr267l1ydUELepPvloeeent
vkwws7Y9T+Sxy6q9/3kjJiskEHUFgpeAk22+MjAJYkFBd2UtgxHQx3JDSrpftD/MGZPM5Qjb+DDP
7CTMrSoP+2qIdKGM1pw8CDQ+y90saRgfsKF0ujQAmJYSyJ2SQvQHFOMmoeC/vXAjaFlV91qSyCYe
Unq9zBGc193prOAD6x5r95QUhp1p7ynqx6BYK9bRtyt2WUkBspRiWci2GxskQBTvHj6kQ84BRXVM
2g6vW4Wz2E5Hht70sJPOtxr4F73CNqcSIq6s2RqTbxr5H2lPK/goaTwU3nJJzAK8JT2c7ypTdlMU
1oUmBL8KoK8F9164VJhBXW9J+sySWciqosFZ7YoEsvzZfpzI1cIAge0+TNDyMGtDbo2wCXQJc3w+
AW2u31vU75G0BX63HfVqpwhncGIrkcS6WKlyiwiIg39QgN5LRGvj2g6dMGcixJT+kTdlhjOeNVWC
o4aFZEtlRNYxGPFIbFSGUzw6WoFvhrLNTVtySRFukCKDu1gKkH2SNqSn2/ZfuBLRMnVU3TA/jhe+
b78nD/P/2Wjw+oPXqcqLK4muxx86BGWH5j5MIUyRy+OspC6DGgFzFf4JlIdL+weZjLZZN0dvs4S0
+kv8C1d8mUSYByzjwgyGQTIyYkO6qy5xufkFezJyzngM42HSpE7uMIghXqzY2YCOSLn644YLm+Dz
U/gUxFHxlZSEgDJTSxSoAPBF7rkT/OyAbtG4nNPRomHKy22YjBOJXWonYsGH302JkPfVgYNFZ/Rd
Cge1+acXtD+LwW5ZD64FSKmLxQjITzozFWO1grI2GJMHuDEVC/jwLbsFx2xdffOmseNDG66TCn8h
a1kA0Lc98SfMLghuqPLZ9+Ph3fHMAa+bktKf16grGxosNb+/n5Uls6ZJHvrOfhmqtAqmjU7JuvTK
RmscG7vCEWNRnWhzXPOhv6+8lHU0PJzvq8fumJO2aLfmg/FhQBMXcYCfTIagHI5YD2Dz5kJBcFrj
MyoJfXuLM7cCewdsmVtRf0lh3OYeTnkMPZCKhCPkjYckY0GN3gfs9ooE9Tmni5Nn3XAzczYzEY4Z
X7hONOpbFlBV2Tx0wCM5ASSvz4pQ4fz/VkXP6gUEJF8ApPueXE+ipITxrJhnh1uPtzB1qHIQ+Fig
mEE6QS+5CzcbZ5XrbWltbjNEqec9PGHzCcnHWIZS2pt8lumq7pkWpbwnfX/rzv7l1A9wVEXRCMkb
oaw/SQOqz7yKEFZ6iJZyeEBhIBGgvJYrJ73VQFdTXBeB0cN5ERQgEsR2pYbJvGXXXiQsXh0+N8bd
5mcv03qoSxBU30yfN57M53YytkvZZ1/HDAbA6ngsAxCot6nGB7yV/KIIO4u5XZuB2Z+hQ6IlPbRe
qkC9V3eKdTk8NRrgxXTGFUeUKFYWv506tVLyPQyugku8hXwuFrB1+G4H4vNDaWu7N7OsfQkXgFe8
H7yxNIMQKbjrGwfav9yR9vtLqcqsR8kmi679pr4n6QTJP3WlhK2w4aMyIfAFscV36qz4RPsSUy+O
vBKX6A90wyP/cxwJJ8WK6GjeOa0LgKQX5L8cFr3ys/s6kNO26xxVwKUg4HTTswXCGQWza5kXhNNk
BO7AyhNifJ93BsmtdnfFUvWa5uDfEcOguobb/17ypy2XN4itIeJoMPLRAz7dueX5YqP8qp9QmoEX
3i2b69cs5KRUDz1AB19hPQNkjYOb33kpOwdE4Tlre4xyMLzq8xc33bHavKpAzsMSO0MSSU3HCkjv
tay3utsyKdH5nrNGEh5oHXsrL4aTGjro/aNcjj3o//GuEfRuaU5sz1HR0zGTIQblehTQzz8jBjj+
kE1GcjbF3bCZbab4Z0fgQNT51YZ7Qow59MwwQtZrjQ2ENj89iIRCRe+QLB6YjS/uL8BRDl+8y9AS
iLIE3BUOGqFHmZ6zh56L8hWzacKiz/SZf6fL+tg0ugo46tvDpDvWY1rqH6o5bsh9HPTOd+DA9g/1
rNw+Uc13HlKPxHDTsSjDjwkcICQ+9sMNvGu8T0+2SQohVQzqELuCaP1Zq5pGKfLjfXiwxkJBg4MU
VUP2ZQSrIXhXyqWcQEs/f+8nb05gusbNscG/9hDeYTqTRGBFb6V6wvqczJuwVSUpk9EFol/EdkC6
l4VopDNwjAME8Pb8XiO9zFL8SAZQeGzMn2FEdAEch14DMKVlSIZUOgOHKPj1pgJhe4nQOFybNVpv
Z2NURsUAMzoECVkEZRYHgzCaSth4TzIlGg10qN0tmqvX+nOk/O2rcGI0xbuo3DK5D09jUQ6TdbGQ
zQjow6fM76sUqJGvf75BQ5sKAJjX5z69UKDE2YIQD9rU95Zu36Y6NV/mmoUGLqlI5T28EPiD9qho
gEId8Max0bTZqbST0PHjvmjG6ZUm7C11bFJigbB6CY0N0+5bDoGHEfsLszXxr/RBPi8f+QeKx1Dx
n36QVra8z/nft15vMAm3aTxlE3/HWsqaRsbnDnSUzXFyCxGJrs47bfv4VlqXJ5ArriYvWaPv1OBh
+pdZ2JHVPjWU3sMcQeVYnVVz6aplR6zUNS3OH5kXQbkFiW6wdbf3et6O9sEo/hPcGeh1+krfWckE
kDM48X83kN7vn7TkrJjZWeaNG6e1XpnAWQpby1Y0B51QR0/BEiir5vB/kEo+X9w5By+WPaKYmnCX
UxrWEbA3w8agheE1XsjGZOuQOnkn2uADx4dN2cAhJCPtTUPvtyc9miDqUve9chAHVgaH6jVXptt/
qy6Zht6OdrSPy/k+t/FsFCYy6rUCCGy8giYhVXBvbp9KbCLPMKyn7Nua9HpQ+EpZIya1HnkgoR7a
DWyCw2RzzBJFMCR1nCh2Llar7o+FFPA8oJJKNuh26WqHYqO1U/03NSP2TGCDCa6SUSWuB6DErU9r
yyT2XQg/WWCokLgsrnc97WDTymAVUijIikOb8ZXu6wkgcWA5bloV22F6zxKO/8X6tT/QE0rda1G+
CAWh2U0ee6MKv7J3PpzEFQJ3nlckhla/mFfulAAkOW7keiLN+XyVyKEmcePD6OoKW9NuAokettR2
h39IdhfKit5YWfXGFqNqUHwKIXsWtHWCqK7V5wIAT4PQLIVn2yVGUVshZOSqH3Hz8p2bG5kEgmgG
3CNFDz4mrs5v9xrueeS+7scWwXTTatKAMYvLbgA3PDcBlMKl96rFcc2e8E4kWDDn2qnUF6B8IQ6r
07PVqN7xdjMeLB+D8oSnUYT2e9lfOKYORQ0axbCRnSQPsdTnO+ZShlq5QZB65No5Eg2qv7GyAB9q
CXtQ3QkdUdDk+W0r5NqLYbIVYJNXluGziwbUhyMynnq6TvPfHwlvoq54pRvugyQU++nqtcJMTSdu
mmRb/Sx8NZXFTHjX/CVQZvSLAALHQI8P3oESWpin1qoR6e2naDflOXZf0dHAwVNAT4Nn84xgp9t4
mP2vDm5RRtflVucsI3kU3wwxfiykDFMtsFJr5X4jElaZz51Z0b+504CRo+lD+l7qZBtdVvVb5bgd
b20i3JriW3cd8liH5L3WVtb22KRVbhTsNjhS3gwhuCsWL2OobL/uUJ5ljSWFScZUeArHuY7dxk/W
S9KjSobO86p/mxJ9ACCwg4W4pwnbsGzHI9LQzLlVqd5Teu8v44rvH+761Um6LGQarCRBcC7xbTWS
4sJPT2HHm8zvrFvhdhIaySCWS1N9XMYx+LNNFJEpR/TXooDunk9jqTNzvfFs2Zdw/8MrhPWXnaZ/
XYN2wQzfZ73xk5uq7neowjjV4Fgq4lNdeGGAMv8WewBUU5OqardTPqY7kE721+32ws6fofWrzzir
+Xfprqb7MVLT5HWXcbB6pdDI7I92U2HbKTpxQ0885Cnj4Q/k3cgwtwGmuF9e4XIVhO1bgoQ9yZ5z
7sG8CcVO+j+UkYho++DHDtvKZIo/jj3RFVCiy9L2gWvpySaroemDKQQGNBzmFGw9rkhGOeTT9Ql3
lzxML+G5+lQp63mKjnpRtKwMCG1xfg55dtgAlMtvzhP5I9ZuhPnjRI3kFyKbFM45dTOnGY1BDDf3
MJdyXOyZP4ZokdaHQdkV6ebqWtHZIIPU1KZG/6Au7igBs91QvL7nXneAyMPjbQQYB7wMHHdhCL0k
ZzaWQUee53rOxoJfflM6A3sv0cNgKVzUDAUmQi6hbZ9RI4nYYLdLhRR4+PyPhqKQ6jWmgjIKymo/
HnX23ULMc0UUw3Lh4xFgblzK/sXtFn4U9xrKBEEt6L/XVkuomFq0tpITOTGjsHCLFrixywh3CTNv
vpzqJZ9QgvDzv49PxLaKVWtHvDvXHBLA4uMyDI/LFJDGPlAKert9o1MZLQ3Kf7R44kZaqhGRNbao
W5bOzJg2o7zO4wnOqkQU/fYVFYJdSF8clB/Zf1+kTmfTWqkdMLbT5E0o4oMimIDN6TLNsIo6qmBi
xXjR4Cz/mLqCCy18RpiPTrGkYHxEz2NSAQ8p4td5SO/zexHOWYOdDPrly7/3dI26eqmePhmC3VuI
5nQUL5uVM2gZ7y+oiX2szgIGUEzcFn0vPmjhuewoLWadmzRr56xBCkfwVOmjK/DjwHMwuuEPMt5R
zArZzY5mF292oj00JxWH+1woRnKE+R08so1qnfE3E0XnlcZZFiCBv1i+2HZphfaMsEPK7dRuzS7x
nwA/DHeG3i1XMPFNUzUsuyBh4rchpq4ftW5fOAaVLsyMOi6mSGTSv7n+uJr9Shrcowo9E/ylwGse
5oKzgvj1fdnqwIr9ALdGZoXWvQd4pFiY+ryvkF39mm3q6NhB+R/mu0sR/R3Uga0kfCUpkHEn6XxK
IVpx41KNc0tKThxhoLpmw4hvc6UJDcBxalatyyL5R+kSHDOoUasoCltwEOntn5OKPPg0t4ry94UQ
KInDgQkJfs3eXsxdxCJ5XNhQH/U98fRxUaiYGkejeCAUyiLvW/yUbuXdYFrl0metha8/8EqeJLhL
CDAz5k/tJG6I8I7PP9RGmXlLnDLt28qbWN3L/9XY44eKmLSGb3rSPoxUiZH/q5RgRGAebbCqicUg
9Jo/ZOjsFmRO/7iun4zgFEA/JIHh2GxCGpyg8CxfA6TBHSC+QIQ3SMnFSzTp4PG0Ah5guwH7thiE
Sn70oRboTV1V/UKD2dgwPA9eQ3OO03LMn5YClLwUHWTYAYjubIRTtn3Hz+Ydjqc41QjdWYJGGqnA
+ZNvej8ZrlOpIpUbgqEDpVR1gjcXf3A4S2tNPXKXeR2GSjkD2TJyx/CHFzBSTzaB6ac0RQpHe8ML
r0byCav3a+u64CoSLWX5ZUokIdEYkFX6uB0kIXDxLXOy/r47ebuRs0+2vAd2kNPGWw+maM6Vrf5C
zCpR+eaW0zMFZrVtn0Iqw4IkZK8qXD7VVmCDck/nTbZW0kFJxxftqD+AsTgTcjkJMyuIw36MAy9v
1OcicMsOpFt/HQY9kr60TzWSBkqYS9JkNjFH2qKDLTFrCUYwIbe4ZUN+D9oUPGl/YUdPERlF0o5M
hapTT7lv0UoY7H3Bh3ZIca9Pqwkre/PbntNTTVz7msb/9QVH8RVBHwtZxOimIBGR5QqE49+Q3Xv2
7JLsKG5DRFKTsAv4p7yA3E7vYO7FoXYGlYc0E9JM5kZ/V6zMNq0wlxO5fKJnUG5pevBes0c/M6Bs
2Xj56nQBjfKQEdPEN/+vKMx8OdmV6NYAHUfQh5LHuTOFbkuwAbyLHFiYxYh0sHbF0iNFdOLz3P5D
FoUEyV5QZNVULfL/VKBM03Cbh1OTPFH0vd+FPCpr5TJu+jxBVcPZdpLqwNa2kTmN3bP/++b0bfJF
hfNSHiURaIPGmGc0wTniHjmlWG6ljcXPOU6XVwYtKl0oFkeAGdt4QA/t4bYJLPqD4VPBzuWTYlls
q7wjRs/FM3I5yWPrE+8YXYxvRJFM5kufCYvtslkXuboMkStRuwTlow9pBdLfgr1zGvqR0RN9e1BG
UqM02MK0PaZvUxqSEKE6C1Wj9P6CIkOvRcO+hQNtNUuYVVkNzNQ1qBlDAk28nuZO78MbxWKxfVkr
fm6xE/qaNm/FeDvwftqItjJlPjERqWM+dgagvP5WqpkJe4MYby7lMoeiU4myP5FUsnUuTm8i6lZ1
dOdHRCnZrxF4LNszW/Jq2NuhX5aAbw4TObws/XuRYOxQCUs02njf62zrdBcBroPBjka+E4qyQ5uw
II3oY/kMJwos6yglR1HvN7QJzn35Xa4YIFd2OkbLFyniFWTHf4zgsaqsveL/vNqQZwbpjmG52KMT
XC5NE9VK37Ft7EkRme/kFAHi7mtw4slOAnT0VbQMl0P7mFUkJgmExiBw0lArHpeRSftENMhbmEvB
PgEYh7XrvtMQwuwpBZddS7Rf3UWwkJdvFvhu2pimqYMQgwJLPOJdR5G5wp4uNjWR35VM8QkJPNVA
WFLbdb3n6CxfPBDfsa9XWJGKP3F49ZRFQN2MV2C4JS/C2YjZqn4Nn0XitZ9tqQscSCsIf3g66UJf
BPrKjayz2HT9CBRWi95ZXYqOkXADLatJR3tcKWqu0U1rynXsltmrtd7y/xiZO8OLMEEKbcZxCnij
pmNk19OArvcAER8pJ9wGPM2oeqxZO10MM7Zgl+yzfpLgKiHjkFWJ+J08QjyqyRlzRV6tu11+Wu73
VFyOXkyhN12B1wJV8hQ9ppB7aDVHyL4PyCAutldGfhKrSlTKoj/6DWNtRPUtUzgwn2nNi+QDUYaf
XEKl/wHKFphxk2UfzfGekndYp7gym1+k+rP9uMjhNCj6aSk7Pb+ojDqahTQ/qwVZDn3HTFfSJqKJ
bd6+XRwcgte92utaFsDow7oENlZmSM6gGXtYU8DW+Q19r9bbsiDHA/g/ZSIqORFZg4WaDPMimr+H
t5WdmGxtGEoKxWR0esGm+jriFLnDHtfrh7GnjakuiqBnxBf22/b1g53vgQpVN04g8pcrp4K0qxSY
xtuaM1vL9/3gqrhR85KhPa7LKr0yJS2vWaKr59ZbjWAe49aPFvYeedI+cbkXhSayRaSdXcpc/WGn
BxU14upBfMvwzZIxASZlH8ajM3LOEpS4pcv/dxgzVhA7Qo5YOvSaef9Wz/lyQfE0sHwmxjlVZ3m1
qM1tfE8JYtEtjP+bxwX/OvaNc9qjNSPUPsv6WRlTC0kcdEDlKW7D1+imIZa+7pI1rXoZrP1PZhZF
sXiSYG/xDEJ0r3fAM4AXGMp+PaguUwrX+hPfsKWE4k7nJ99fwYEj1mnMp3wrx3ctSyUQnpHkO06+
ldBOPp8+mzifusvgYmb5UmQphkxSBn23pZg5zgA/DQ6pDGaBBLpsI0ml+JgwXACXXdB0cKsj27bu
ML4kULr1UZVm5HLsTRWicyczRPSVBwX0qzKTsis7QGB72CGT6B2omW8UqphkO0hnFSQZhjmOmGli
F+qmUMETXyqzOf4C8hVa/XWRU23bxXpgRNHsVmdoa+He5hRco7fCi2rc42dYFkfnoQxDNzSipEB4
WsFfvmj8RjF9gSTEcQeHRf5W6Uq83zNzBBlWFgW6hNWbf2pyZzY8cJSC0erLu4zD6zPzTg83AkQZ
qs3btIhCNA0L9pdwVG7iPhn0NzhbtBfUb9DqvKiPxb/NcFPMggosJSEk4s1p9EGR15bbgLHkoSPf
I3h6Z3TRWaAa8tZq9JFcA9KgpBqodr3u71+xhVav0Rz/BiMHuJH7x8voAYqARZSxOWyqt1FYuvgq
2MCDJcvT3B2iXUe888ui2fn7nWjYONfKB68LDM2QhNMeZYANQN496lAp9fSF3yARrCwD222mBqtn
7ezgYoT30I3eUocD7CFihDO8iq7Rolqs/S1eAVvCb4DYrbjw0yU1VPLAYYfaaS4I4fH81A0e82Uj
ja1MXQkLxMEXVZWKE/ZME3LVp2FvNxJaXskzKg33VjRhOWiOv4KLMcuqhPCl2FKZAqQDeZ/eua1k
NBk8HetgiA3nJt5DVmRy/KKBzKprvSxHNX4+eQdGkD4dTsn1ZrWaFBqp6ioPpZsTBC7AneYXC2Of
+txroOzyg/RDxru8aiQWi0dfXR4bz9X+2ZENlcWnC7Vk8L2fGcEX5wdmRpwQ/szKgjt1sXBwPIE3
5L/2IwdmmwTq4GiHVLneypNLbJviMGV11/JwLmL5uwajo1mNIkxgnq+iezAfc+3bO5RQcaa0FEhG
mEF6z53GldEZyPD3InZww+qWwOGUwd2Uez38QppE5P9zEwtT3VO+3uyH1EVz4/cF9X/cb++mkH1v
CJrPg07mGk1FVTzEpPTN2iDl3wKhgNNHdjOK0lDycGFUtfIm9ItB6DSXhbxyR+6kl9MLZltF3RQq
9mr5bdfZpMvU+wj/zszYtRgONqQhEQP1u4Idd1aEWq8JhZkxxoqACInSyaX/30OcYGLVO2nn+sWy
RTONbKvxDpEyA8mp5HIsN5j5Wz+eImSRx0qQMyrGn9fKjeciQIcPN3wE5IBeMKwdqPj6G5lhk/FF
JVy58++byOf2l2BRDwNlxULobZyEpkHayqSNXPWjxvVEybpVqSs8LvdAIydzdZWG/yKeb2wBbbGF
hb4GSxbENfKDIXIoI7I+55Tgc0OWbWZIasQB3geMP0tdF4OCU4gVKbaG8xmWupAPY8dUYuwqVEFH
fL+CRcSaja6rYJEZ3L/0IxSRQYplkZK9IP1m3pgqK0tupkVAaUTGiP8ZB0I+xiYUNVKViLkyszEa
Op/LKbbE6O/0exA/BkegT8ntY8YSyOqEPKe6ZQxQJLy3YI7XAzykbbF3de7nqshRc9mKEkhkcKVo
ySB9ktW45ZW+B9Pc+bRTrCcxOh4r7LJ3jQnlOUGMUJOne4tycUdvEsEBpTw0/4aQ70O2ww1fbXqc
zt3obyrQu6SB3kMtphC4kxzczXQSNGDCHZU5IE0g649sKyQby1bnDXNyESWwp+zYMz+PCnFWxURa
0vu/oG+UCeyBh+6vqDeG2q2oK//1/24AzM/G8SsKJbmNCJXt1JPr1ZW8L+SBYdCWNwKlhxZTolgr
De7BHAezEMns135K7P73/lCNzGgFSBhMi+wPLDXvmN31MxHZJnvwx4rbMCztE1nZSmpTJNihC7pU
rwCVQUhVPsg4hNEwxW+/PVoIm0/ljoDbxE+UhVejZiTowHREzdbDPL5a/7KWZ/f6raVdFsttqy1X
EQRcauVu4wGrek9AGudEHS1Azmh7BZBg91EYSBbv2R7eSWGjzmp9CqrPWkT72bOLtqEdtHNa2ERD
kdFrtIrdabKlBkmIy6TTIH64a4WIgS/yImkuwPVX88R7H16MlQSaV0vFB1xOs4eHt4o5L2YKdiQy
PpRK++XG00U8JzLTBygxFcZWeuLGGpb5u2bzAF1GmAsus+Go4Rt7EcCwgGPqXO5mKVnPPT4nUwuO
cM7vsieLt/lVLrIaaEgpXKhIQCV+xIj5owIUIkDzfpH2KOesCKRqdxkU9QbgMgbyAhSD9P/ex774
EPVYZpWzBFTzngqtE8zieHo6vI7vmgcCLgher8WLe3NsnQnlVqaNgdcpt+4lgY7gjO7eFQxUMdiW
kJ9TtWIujS27vUesV4CT4oPK+BT19b3MJ1VTMbkADqVuS52oy5Sgbk/hMyIj9lgw6dfe2yhUfTxL
vOtOVCnyBaVxgdBYKKpxeEsLFdlxPzUsN1ciqFM17PPuqFt/0WEkziPuLNyhQJGXoDYx73d8Nl4C
4qNZzH5CXGWzN9Al5iMx5lYa9GrmFRek+SgjxzjsNEaKvNG3zAP39emhjkBEljJIkigkl+4aZXv2
S743Qi5nJWUEgmTtOPMB5b62Vyi/BGuS9fVCZA55E1D2Di04SLc6WblPFSH3VBZ/+LaFhLaY8mxN
H1czTNCo/lSxUQo4PDpL8X3qUtZmwtLAkL8cQes/kVtdsFBIdhll5G7yKzEM01xn6uhYRQDJ8+n8
LYISWCbquPRd9NkmSnbX6zwsDJUYRR6kbE5N1C1umvt1nppoGBo8rr0iHN489Hv61kboAW8zlqxi
PQ5iRYPsffmzD9VcBHWgiFwTHKG8/VkXCCg3OCkXhdF9IOMD/OcpVkhZxS53+4LSCWYBM0YiTZwW
DzRnNYFMrWtoUl9tlka8QqzItWFYeC7ZDjum7PMas+OYE7gsSFPFqkO25RcRoYpkqhAcujQZU7Nb
cqqtsu2F5IGx+Hvoc7MaAtXlJ3z72gmLXioy7KFUMdSiOsF+h93QhNRX8sYjk6zadjQq4Lr6CxEX
Dk1NJbXdew+i/gI00/DjIV7szdO0suxz9JV+iJJ3qlZZu4Ko0GzKyiIeLzQvrmCN0p24ZGgiPS84
Sha4vE6hsmk3eNjpc19NB6dCtbilc8ZmXvQg1pokHTv+SSS3olrD13h0n8Lc8El3JzlUdSUd5qmg
qI9NPhFb9muWnqx/j0UQ/xLchHaT4uxXIUrT7b5LMvPHgxQMZXT5GnK82NlheS6vQf9kIfyu/U1G
cUlTTigCt3Jj/tWxD5jNThRRulmO+gN+SSWQRjee3++eVwpZX+mqxBqWSSRZeSgFmRqCEhGoBZ6o
MhRDdUAxH3MZagjCJoK9ex/JYta6YO7PiBfXvYd1IYjnaQw1VuCl+Ryirjohx6QamGYAwfyjOFjJ
hYHoF3LTL2sUB2/Sibq6zGqcPVWpYX+xYVejU3wO/pENOx6/IOyy33ghLVQHnwnv1ZzYx2IEv1sH
AwlGjwS5VXjLTuqQkEyfjUHiHQvLDAGgj3IoeRSCYKarwTNEgNPKe5qiLfao8xznUuaj3gKqQQfN
YfMUeGQqVX47fQTM92Y193HdHMXnBPxnufUno1qHb/R5LLWu+iS0S5qLuGVUfZON5kEZvDjuHAoW
FpjFZOsOv/Ff+C4XjirD4YGQJB7tZmJDQo2vn+fRcreasciNcBM9/4RPVBgKNf7otQ7Jdo1BYsU3
yz01vFHydsEydVZKhRzoHayQJ7k5qEg7UyZ1eOIFBPrPnnMU1+BQ8FjNvXIP1fPDyqNr6LVT4bog
kbXC3CK/ZqrwHR4uADCIsehaq7kCizJtSc8pKxNngGbcXs7wZiMtwGzS+dtSuRAyk3fYrODlMzJl
WMfno3miP2f5W3sDQT4Mw1SsjvCb+xKltRzrE01FvoyuT0nubRCk5uETTSTVHqBBiYghNXtXVDEq
bXE74vIRX/EFDscnrA1h/UwxvIlVBRd1WjehdLHtJrKu5sHLjB7k/3QNOQCipm+MUoV7UrsKywe0
0GFgtku4sAKmK/AhbI+2v8LpRNpGqoY5VG3PAw6OnPbCHQRVVU9rvSb39Udmrfsbnz7rWsmKNqgs
F63vYf+/cGuYkVqA51HFPg5+yWaVXLFAJbLPGljl2EBpcKOhj75gmWuixPCzK0cnRrEVDInCGTvz
3kOYAL6hvGjw+Kwxzq28nMrAqHz79X9EHl3iyxmLg1FppZZkcAj5TvJg0Yh7z2nwQcGSGaf5Tzek
z7OuLEwQRsTFdEL8/c8FOnkrBhdtXQEtzK9CI5G78bpPBFeLJKnrTYvYXj3zwdEWx8yW9lYBJYkz
QUvZF//9vj9RmbvNQ/QClXCMZCKaDpWnff+qfiLZiwfawiFrLlQmmoeQsw8jItxd+IX+AUjDL2fE
ZCvODxawen4G1bIozKiSDSN22efv1nf/2JKnjS8wf2Pcb6QW9pYT9eSaprlQIfnBRbrLivtOyOyN
WRTLp36J76LGbSVd3+MfFsP//MtTzIqFXnmss57oMsmk0EroScHwfvsiorw4yff1VoRSyndPTiBG
i8lJ501LPSrpkc1paXNivaoxD3pWx0lofre064/OlmxnzUfZuO7yVeBzc2+E0d6+ZxuM93X/WUOB
fsOU48xf6/7IT/C26Z2kGAKuc1POU9Efav8FucFuxQup4XutkW2V9fRlrSvRw8/SKjeAXgn5AAEA
gUc4x90oMQ5ov7QVRd5s2J/zvIMYLMHrEJoKqdQAAdVoXx/+qISG0h9qtW9D6zV7m12eXQh8xc5C
F571lu5h0WeiLlOm+YfO1pBRt0EVEuAJ0Cqm+kac0BRnqq3ipDZXpCC/tk2a94pY2lkBQNOn9PS3
1qXCZIZVvNU/dc5oS+A/nLA/So6TPphzCzkkA7dpTeNpmROFjbllIBWbLkengWk1/qZKa0if+VjM
m9rb/SD6cgAJqRJ5EDTr+I+J9ISdE31Xx7YhUrMWU9Vqu0pfsy60AzlLJRmvU6hYEdBFwQ4cEyzB
aXY5lC1LKwUfRAkfaS0i7oPka65rtOaZEPg4PgzHLi+eIjtE2vNhpEisK3yDxYA0ilKojENR1x1A
5Qt0uoEHwkPwvsEEARBLZ7lan4JP/WXJC97pIMRXVso5ou4y1OpiSpo0G3fR2/Ni3XgKdeWrZdgp
Muc5N/LYDEP97jGFHXK/gFRuwBcFEVnrzaqOmVPjjrpHc+Dav8hIk2A64EmeqPQrrIfmbgdt2rUu
je8eoLteCyUcDZAtvh5r/7+lnjsdYJfKTZURJDa7+jiSFVyEfw88BoSHzzOqK7pbNCS7ICQBwKYj
PWUIaeSMUc9NHENz92ucmMtSGTbFeb5vs/0MrPgG6AeVVFz7miNPgDgo/3NljgTrdzAnkkgTKcx7
BXJQoLrzyolf1keYpnF9rAjG3Ge3hI+70rujPsxcQ7Z1ekhx1w+qDlUiOSebjjvWyrfuMWNhhfyO
EucEHYYEkGY5dFh8JMag+7Le6127w41WotBg5l4Do330Qg0SNl8C1dRPW1bBw8qfgiSu1yCKYf+P
foV9uyww2NBKXEs1+7LAOaZ8j5E4sEjuv0lxgv/VTHBb9jW5XAZUQnBhfLiCxfpPYJZFYQRSZnI5
HJPMEKbkcNl8Cj7Q4PWcHfTj9rmcSjzdrYcC/1zhtJoamyTVTbPSWfjOamDUPp4EKD/LlqBeCwrC
WMpzVwlrSGo8icNk39miZF4Ws4C0UPK9391jotTqO2bSynCkZdkWdT7TwXXT2pXqPLHz8YGbby6h
rh9baoYXOX0+sknwh+jWnnXmlvFZYtr0zHvuaF+8MjGh8I1k8H1vBlTaRx0Wiy13rF0FxdzNj2sV
mZO5rWQGXkKqCGzOhhtjaNA+yR+1nhmfp7zJ8M5xAsFXWjYHo6ujzIweVKLzIfok8r5WcuUTw3NN
Hw/CznVqUfwbKgxgGO+ISLUiKvstmjXKjIaKNdn7bQLjGY6N+r/ffhauB4dnnqgDTo4twNw+HN5s
NjWHSGvaw7qtH1ThnoqK+KlCEVMydiHxEXyoD0FuksnfUZSmdpH5cGFCTyDbNNByivpOfIYBubBL
1Em5/TP3rjXcb+Te4CQVc9gpuiXVhEWKLJQIl1mrlWYvWv2zO/qVfgfZi5bqt6xEYXgz5E2d1m7V
qVDPIWCCHXhS6kuLKGOJTMSHSZwYspWvWMMHacOuJd4sl5wh/T0MU/0G9RA8Rpc2l5EVIlS5Kddv
pV2Dn4a+1U6pSbaRdGpBOSXa7RWwMCczk9fuhP6IUcwnnZ8tAwoGvFzyWHwXZsDsxYTqEsjcgHA0
/wl3e8BbyYnUzJ6lO8P0/lT179g7dUS3Vk09s+BgeZ22aHcoi2/uwNi+SArLB+ei8tMr30C1Ub5r
XF9dEh4ZnKg9FXSeM1RBtJ4uWgBdNy+mZc0CG0bbkuC8dpvEbXuBcGgKi12UBFOKJ5JC1knVl/S3
upc0ag6W7QxXptZBcTinNiyNYuv2DPVkj66AuQIs5A31ofH22J3hjqe7ohBP+xAjhnVQgL9oYt/1
Vpj7FQXcGB0TndTMFolfHUksy5ELcsYHFsn172QzV4lWA29P5J16WuVM+l+aTJykd78wz7aFDb8Y
WgQhVL/NGiM8bRjQ1OK0ODn5UeZPm0WpRBBj1XPGYUyWqDYQKmP5nWJ8yvOuH/pdQ9eHvknjJthb
JzxWt9N+SIK69IYgdvBFcLfvh2Zg630DfLPhbJCIzttUR3dJMFjG/9tpga206F+cECeErcZn0qhD
V6wSsxXzRNuR/yfxnbzW5akMJEXFs9u20iqCqLszBWhdy8NslntWrdCtqUmDdTBqI+DTUoJeOQGp
yND5yZMF1st5s+lCUa/fF2erMBno4yLxNnRjM4PvKHqetk648zjld733Cdg+l/gtmJJYjgScc6oH
GTz9gh/UIG1Q6TN5En7VNDO23dv2qojUgVy7ERkk/P4C05yjIlwMyc89qFhvXiRumvgf+bMioanJ
892mtAORb81rIKIThBm2mJzoyOMKVoYQhPsxnGRTuJpip0A/cVUi9BXZWaNaglBxas4VN6tk1WMk
DiO+dJyS6bKiCS5V+HikjUsB9Kk6SD09L7BBxmm6G1QiVH9sEt+X6BPAV7XPEp103d0QoMMud/V9
lPknyPCq85ppqRuPhFHouNllhqgA3wA6UUtL+6a13jsdl8FucMNbO3cOqB1GeWpoja2MlWzNsM7i
rpM4baBnqPTJrR6RBaCNjIiSYC1MxhU8cFEcMnKDBrYsKW3p/beXXir61a8VmHGm2Whkz86NKzcG
ne7dIDDgRL3SbRYrL/pAIQL1kwZVZwN5Jys8K5BhIDKnChJfUdJvgYz0FBorthQbt4Elbtw8pTyi
AXdHUdrQo//4sbYYkCNPtAqpVHak6C5+h96giNql9EtD/GS4DV6s9kuh4FaMwByDWaAuzzEnjABx
2s/GtD5Z+Qp+Tn/4/KOFUBHnDD47yzagkqmYj0jRYEcqJ6vjhgFdJe8VdK26hYf+cjo2EHVz6PDn
TO7o4pm3v9zef2HIoGDWTZfxaBcuGvutBodkr5SznL2bHbCUqDs95pY/1v1pa2MK89UrCEasPl2p
1V+stg9bbQIyp83Q15tvq6r5uSCpLR1IgV/ZLahfeQiAvT27TQPywmKPC5pt8x3GfM/lkeaVVLu/
jYgOeO32b2/rUwkPqIqmrJ1NmWcLzQvsZKps0+ie1qfwch0OvQBspGIh1CzjslXK3kdi4CsQZlFN
YpaujXR41ce/hGoatQpiIpLlQpP2ujDZk0ApJfuCsWyunIs+4YCffql7AMde+sNGgL0lQ80nLHft
+VBU7ZxmT3Yaj2PywvFcfHvnvxLrqVywh50DIwh0wJImVZxz4blwcEA+iaWv4HMhIoQbcJuFGwTQ
Fo+GEJ8AQEdvdypSSn/DdjLeBrKb6xYrzc2T/LS6icZAPiuMlI6oCRuWdDKUKSTHk2RY4dRi2x64
KXm0JhUBSl282RyaGqEW5CQTVJAB+//FfJrWJvfRryIciQ6RekxQsfmtSxbB22Q4Hbl7Zl8ydmTX
Dj8823/Tpn/Edm3JGbPZ4F3yjfOBIHEVf8Iy/mMd97cb5klIxQPgP4J7gaMN6py6J4gly2P+2Xkt
A0oVEj7nFpJxalfazrsj+KX5jUSKiwzBeuGwWt2ampy/Ay/ffc0aBlpTTvYXJtedqxfHTBX8aNhY
CtyQ2f3fCCM+UG6j9pxcswKEBNkSZmnoc90zbGSeJVgByZqUWLS+YeL7wR5KXFKFyTBLo9K0I7+B
1QmRFxFvsAMfNod0ENL2WyeUiAmLuo7pZ/kQ9+9Wuv7Tf2xFtXTxOQq5hby8o4CzGk0PZHv9swmB
9n/xZZXvGe1zsu8Oy6fXQatFYtgbaHL//8/6Kaam2s26jf5+/sAgDj92fSPxoPTBIFJW6d23U5xZ
Am+xF5pAH8Loh4ttd7MCAaY0ItCDHenNBibcKC5gNFqFhZOrb3KZlbTQ4zBQ17BYlNl74BKX4hvh
UEHfCoyxn9RiHQNgJ4AHRQYrwuAcr+VNXRzHTSCc7TCKlHoUP9PImXXD+ccwJQRCy8E1bbljk5RQ
+wRoTvI5kCuwX5XGLuvk05RwVZsAeHVG4eaNTnpNVXU+8fhvg4oT35KEkQjizN0YFC0IigM/iY3r
vch/0eIe8nivs+3oBWFHl8TNh2qpazrAsj7Z0CRub/AhqCkMtAmYWZupYqoGgPqQc6HJlOK7rGZZ
AmKYc+YnQA6wAfLX2minWG8/KFOoZ4w59QOXVo+v4DtDC+171HZIh09AD/A+cJiRFOi8hayuS6Rw
CszjRg8G4RhFd2kMHAeuiyeTwvYhRIuQXq2PoSIUffEE1HuBiG6EQLpe3zlFgvkGTtMcDG8UMEwQ
OejfZuq6p1f5xb4gs17iAb+gG/I9yUYUfo9bvrkxZjxQymoCt1KaD0CM5qtxSTQKbQG4ruDKtgon
Wchb8+1cjaX3eRWXg/eiyUfzO7U1pKtZxq4ikUhZR+5qs1AD1xjj65BZGHzX7obR7BsrKfyY3pWv
H1hT52xqMXgpkqaJHwvdeb1n1Gdq7KRtQHhkwHq6E1XYdWRM9dStwlasCpF6rOoZC7YgXV6Csmsy
Pu+a66qXNPHef/O9O95CV0CGYuDhpJeVLVVOnt+JnwWfxD+sWqmCnRXrYjvUoTy66jvnBN7M3IBA
DXUhF1H4jlNlclguSLWHISHI7kJHlAEtLMs5nb2KCEcT5/fv5s5shicynwqVByRbF/Bn/riRtNQr
I1dP0KP/DEnoFU8PtHz0yBGGCrUe1gYEk1oY1dSxHKw3HOVl9KDUTzcbPMSprvr4Ym0kRrjskwWi
CxDBh+sPrDRU2Np9IMewFoJ6tGZz2UjkWglmGiSvpZF++KaxolNql3xfzghc68Y4bvq9tSTntBOF
U8aN1p+qRohRp+ucJknqaLdmVoXfYWEfBD4q8eBRPnm+6A1o6valavnrE/b7uYAyJpz8wEqeSkSR
WybpQs8voD7yVjQg9swcbbj8EBOPYExTZ97M/SCHuOSEVGoK5w3yo8gznoyA4zGe4vUH7C3yeovY
CHA4roiZwAefvlUrp5c9ztLqP47DGNyqjGyHudxdc+wLM7YnfROK7XUBoKJVZVyM2IhY2ImdfBaT
LhqfpvEjbFnsl0w7Ex3wX0fWT8Ak2D1EaSRbo8W47OdeUE2LW9ipJ82aBzIOd4HVtexhOF+p2Bfy
iYPGxQCa10Hm3kKfhShClf/pnGdMXpBaribSV2NDGFn9feKsOLW8ObKknrKhLepw5aNlKITw1Owd
3ZGRLfUR0ITPq5LKrA+YG0bm0K0KFkdgxPxu0ovYsrgGn+6xk6Yo8uq1a2Icb16R+kXH+yPRslMU
5HgNl2iNIBJTOQ8RQNBTu1K/z2XmzxEd0xf4jWMUR187ZAi74eLqsd3FRUOHZyFTC+A1d5LUThId
jdFFTQRYMybqELXeTbyU/j03CQSd36aQArJ69BFXgiWE+fE7r1hOR6eTJWxcnogSKAcIGsfUnXWo
RxYoqiDB2MTntous8ATdNuRS56gpObdOMtw8i/mmHHamOBFXt70RTGXRYdwSqqZQQDpWsaDBH3ol
E5jc2M6XcferPoj7ZnPU78B2xLPzOihoyGsRsluNME0u+CW7SrXAKbRPjxcPv4EW2lAgdKSgfFBK
Zal+apBez1dC8ADe4cM93BecB4GuR+yikGyuLB58NqANTPHAtJTyVEFNOPNChMvxfMwjJHZNobin
n3BhGXWKbYjBYeQKuaQchXDT6IKqyF7cwH17Ty6u+kCkTQgIY8rm8r3KbgZyQHcepk9TxWTP2nml
5batkG9+eUhu4p1o2NqnQzmMM6nAlT7LLLgssvfpybhWASagjqk3U33rH15vHa+DGwG5kffc2ulM
cZ21McZyoKmpVFY+sk+5VLOjqNlpR5ivVTHssBFTMJuq4/HljRtps9qBP7Thk79lmn9j5nSufPw/
3EvANqz6ST1VTqzkHG7BXoV+V7ksfwztREJZIHLQIbPmXrdpBeux417kzQPIees3+Q9EIzPL+beP
+tV5MkbDil6uP5DNW/hgXvtxWxfVg+nq+7wVkuQs0351ijvC6Nmb9AZtjVIiwVuaGxnRJ1Qx7ffF
QU44sYH95W/CB94evnBR1Ph1rbEJ3uCrkKHlI7s6YfbY0qu9HCVpsEw5Izqt+kqBP5pgROKmoUGb
T2DkD1FKnEcn6CMmyAv2EVxiuQdaFlqYqanNfyBt/PWuiWRz3H+FwNYcNclH2x+4LwAN2FlFlWtv
cQH2rbFIuQPfV+ibkaNCeSOT1PictoUzAkAbLTSuN6x7lmSn1aO+W+nR/L6eMvb6lfjuLKDtubHj
Dgvglsc+rVttcY3+zCQ4Y25hyFogPaLXZwT9AeaTQRwFNKacnw1Q4xGmbHq1NkThnk2IVSQFqLN/
5EPIQRdXWFDcR/CNq2m15XmfXrvXBHwwcXZm1CuZr9yAoesYpjOX49cutdLYRlMv3BxaFOdjTSVz
ihhmn/bWejmSVXaQfVqo5Xjc72V0FsoioJo5u+1NmxEXAPSgUOP5ZyGQq023lfAK2Z1qozOg7eeq
ZLdOTEbRGegQSacBVop0bCq6Licv86mc+MAOUqxnKP673NOkHubPMA+Ge1zjrEmkqX7SRbASKIlI
crBW+U+9utJI0BcA+u4Lfh9I4TLdErdzaEY5b0beqFYW1r0IMJUcgGArXHc8OP2jrqNbne8k3bN3
pipXugxTJ2hHuGBdfOY2Kn25s3Sxa7m+vbElGVqyUJSN0Sq/gI9nVY/LgAJtv78ezYR1a5HbZaqF
EZLFY4D9MylKy7ulpgDqnXpGwc3Uyg+AecdVzQmzjQAfFWz96o+bJJjT6IrNPlIFbalaCxT6j2wF
Q4802ROUORDBOqQypjnEVPUs78M8ocNJ0wbNUhXOpiLh4YYb8PB0tb+RrxMmWUFjCRUZSBD0OcbZ
vZ+UIxd6/3QQz6D6nQc5Ii39/iSwlfntlpGX2CaU8VJdnXqYs+BxRpufasbv+9/B8hCsR7o0Lq3W
uy7EuN4bo22yqAobjnIZa10vGEmwA3KM4Fu9xPl7/gezCiDQ/MjQa7J4x12QsB3OQT0oL5s82CYi
WongaSsSbPmtP6dBjNtXO6QZfXgUZKSeooXdKT73pG64wa3dPmXuUf4/BOiHN8+4yHrBSgeOyiwY
Qcb+9hgPmNSo36lVO9U5iesTwJEt+UsQKFIc+DNZAIfz1F05ZT9uPiZP+ms/an0lE5Wewl57G19P
wL1Zo5utGSk85F2J86FPV31I6DZ160OIGV5i4GXLt3rTVCc4WKwWmK4E9c/Gs7Rinc4uRBZclNBA
Nh8NOrCpA86fbOdJYb/J1sXbi5mzECOXoMjy2DpRfJLAsYYszghAEt41d0Sp2LJ1QP42sphRM7gV
h4Xx1NQRZs7TGgULfGaYysX3dyPHwNNkh6HXj4c25c23DVbh9+UFnosJR01EnWby20QrkP4E2xxo
d5dkpbI3dU9K9qqe63sd/CO7zKPX4QJJ8lnxW0VMaRcEkrrKJFRM4Tqp3WkXQapEtJaAMWWwH+Rc
5ptMPYk1zHimAAVo0loeS/e5c79pGHrARWrW+4I/OdVriRQaCyG6aDO77M1pzahiZjoEMKdQcbBM
YrejTt5aTR8ZKw67VjNVrWi4AYR9tVnBvvMvC62ZGvkRrlar12yn8UAxG9jANBHxHUN3cOhoC3wS
FYvB8iXZ2HL6RdbWX058UX1qE7/MDd/qEZcyBD/a3Xc5KZUqON8GSMxsWK84BRfp7AL7GjVk6Pt1
FjsZHod8bTM7AGYwaC9xRjhY54u8JYWd5rAmFxI+Y8sUT4ELvqFN4HgrL0ZvKrs/u1zF4ifPvehh
e/YfoggZ59sTpWuCIcn6lVLkEi0RtGvLQrP2hFHPjyqqcpcSR3duVNuvznh+x9G4bkk+XB5ASas+
J/apKRA6A8Ms2dnD+YxwKfa8qV55842uKQhl/Emwjf0NBpmjJO2Porf1INVu47zTlNqcfSiFFrp1
ASFVfv4BScf4X0230lvJxqlvm7gZkx5775rE1SN6GeMWi2vwfWpIi1D6xZQg1elSJ/JVfpK75rcM
6Rnq5qJRjIwnafuoc7meqWesmNvbVwaTksMzyx/0VDym1Z1gArvAPyMTFQrCvsqezvgWelWvg/sJ
NcYqyizqKelFZ7Ks1jULlRkAkyEcbMuBSA0Q3PfISfLPOkgSSPd/tSyQHEoPmP72OqjhneEdZPc7
1/HiKl5MCRfj8UMJll3VGxAujnFyW1/M/txE1dPeDz0ZF+2BeYksby+zWTNd9+TrodU/Jn+6u60R
ASBWF9Y3UDKXL10uq3XZ8X2pIbwbIApAaCER+rLJHPjh7VZSFCj/MJm/FnxIRaZhaGyFj4oO7EYP
ytrtdyLNUjz1Xr9rfyUOhTIypPGvig705nDSW2xqiWwdguy32pvopDcZiauNH2QsCmUAKKgyNaUf
cSpJ53lT34akrDiGNnbUudxUuCykP62YMU/G9is2zdK4l8cAvMD5n4cCw3j3LpXm2gPEu/wnB0Uu
hDFf1mvewOCgfim/GG4yPxoaAa+aD6T9f2eOZ7O5JniCUdzjGcdW7hhuOdUAf6NwdpUi+JtycexU
TUH4KsrqMKOzxD6z5Io7id50j7+shlq2PqiH9P/YWQ14OrrZgjoBgmVxyfaZTPjnb7yE0xw2QPZp
6EWqnzt+HHL+8jmlS+hYp7VCdQaLW14pYmj7IvKwnSiVHp3db/rZyD9J2eGdcuxfhJR9T9QlFbXU
JXi6MhcftLDZOMjGmIIXajS4XQ10LXxDGazeIAXPBInBFUymwNtRLSMe8/Td7XONtQv0pKSmQIbj
CYWDtYF3WDbxw8BwLfxamL/sDFHgLpxocpA8tgFjdiwdsG2GMrFeG+Zq+MK/AFNbbkVUAxSaokbG
PNpAlA04U97iDWSKY/qmm88Lt6F0h/ZFexCD9lPxy4Kr1VetwJzLr8ayZpUVnsrbIhon4gJWI3hN
I3s/VcnsNEpXAvamUC0Mxs0SkMLkbKPunoTbGaZpBJaLWBB37ScL43urlvul9cF32SxwXfgTBpfp
SglMAiEkX1oYer0Mtlah2HbdMeXTMBKu9/VJ/HZg6ux2FBHtQcgb8i/RGk2kdFiqASbVFYeb+6O+
Jojf7U4Lb4DOVwVgFXwPG5M09uJmu6s1VsOdG34ANTONv3rHBRtEva8hDmJcDDVfFsSWvYQ9NZdC
OGDY6cKorpYeLjt+QQ+nnmMtOawpOzbNHsfgAd9AmrKiKE6TrYZiUCMtEG/Bd5xcC+saePmaAJgx
b1f8+PkkoOnvpn9FqnwFZgUXQpzWTk6EXYyab4DI+UhGU/4YeTe+Hsl3SZJ6G4ah2rc3Q21CQyhC
0W1l21IXGDmMYvyGCjV5rOuxKWW1QSKmUQfDWm+SzdJOkmiXLHW5U/a+ceU7YzFcBWoLgCFglKlO
QWMtQdCTZARK+hK1wK8jqljhi9QFC0SskTvuOA08LpCrSfHPnjl5WiLSg5nX5dc2XcikH6R3xyc6
WyJiVlzLn+l03GJcnlF12GwpJhcOJbkcplv5tK4++poHrFaj+b6o7yD9DMrKwmQ2FzJ2vy5sC1Se
XpNN49jH22DnPN2s6v842wKoO2YmrIPIVhBoqj831Mq+6a9axTdZnpaEtbCar3dtCnr0nDk+w99D
1euAXMvYq4E16/Xa2u6wnOtjJD0l/9N62a2oYKqpREQwTYx1jehtx2guHCsXUKre5eFw+GuEnopY
f5bzaHeqYultNMrvYqTlwDfZMDZbL9nEdCzyXiDsETLdDzxPwEjfiom19S/pBRDggZs0oyaNqP8o
1ghkczbA6R+jN3Uwxd2NmeuzoeQkT9p86/ci5aF+DF6OsoGIISP8M+6RJk+yqzk8b5gTuonmNF9u
liBMnxap1qdzuS5TLGQnRq+B9XC428+vByB6copiPi5FNmP1ZOTcQL+kC7SDabaOiU7gixb6bfS+
8vCXf3C+DnOpjg1ZO54JiIq4QwJ0pbURYSoeUNXTylYi1zMx7OSA4J4z4zQT9tSqIwSNs645f0Zs
AyPE8th8LBsHt8hAzR2SEDps6u3MJ2ltD5YlEqtZLnhYj2DUbAO/yzNj3V66pp7iyhHxse/Idtca
7CiB/FJrQXP6roHEX3VNXCCfRg7RvhhEaA5RJ/6FVDxxvt4gf+ilMX2okhHzyofNCVKdp2z4xhkN
fDLBTvnjkNF5RKrWdaVcqhbmkzjccJDfE9/afvgctLMiIkVuzv+sZ1A9FrwLs66z9qRwF/0snnby
vXpQT9Q9sEbhL7gW5fjd92aXqeL5h7vWJvpqmEOSQt25E0qLupgRPKmXzVjUofEF3zJ19qSIVkKJ
eF8OkN+BlKhgOQvRN6Of3lbU6WOFJrExzOnrNYljwgVs/qa/jbpjtpYbZok8NbNCQb8QuciDx+OR
EkSgIjwagxHFwrC7Y5S5NWKZd9UHZQdI8NHNgcZPYF60mAHjiBoN2UbBR1/lf92QcAPJ9CCFWcHL
at5f9yYHuoFDYhWrUKWTZZ4RVofJFZA8+lrABdkCFb+59RhuiA0f25QdL7dPVtv7RKPfMMJZYfdp
4jshYwsnvw4BMGcghy22ZnDPUwq5IObxG3e3W1h6y15uTGVXuI/B6rgabWwsFR3rkPwQvFoFbpQF
yANqbO1m62XhnC0faoDg4TWlBzlZmUFRnknHAjkqEipdfOp7RvrPmeyni8iR4TUg4EHsAF8OHrPn
eeT/ul4jz2x06+yM4MTySk8/3fUEDKfPhwAfy4eY+JA5xz4YzVDAbRDMryr89IhDi9maLxDwXJ34
rgCUh2jie0zT/M0NkA2QPBduCRKfxpOykBbRm2dbcsVIei4p9mO0AedOsht59XqUQMjNeK1sEVQn
ViAL35JnxkzchKwtsaGQhFVJX42zhOtvjbYGu92jCCg4oYc51y0gUsqzWrVyPYJIAODS+4HsIIKv
1BiSOtWmJV24h9rG/tTNbv1iNn3XXodAncsykfGy/mPa25JGvNp2Ej3UDEwfqU/Ut6lWsuwkyqzk
820ffWd54T1gFkJos5xHfrAaDGNifO1KYXDSD4cs6odrFfqwSYttMfnn8DO3XDv6wKMdEKxjvsXi
CT+K78xkN6Y9bMeE8RnjQMSpVxL/mcF5BF588f3yg10VjmUpMbJX41hrNw+WEGwPpT4NXX06sVcP
jcia9UyLWIqm3rjpgBSrATyQafrURVS8ILhP4dt0Y8YxidyzuzCQIB7gxvT8Ri+EmEhe9hLoiqjl
f7rQVJrU/VhZiXU9FMog+bC3AJlrPUJVwK9/Wxu7b0mIQhGqz2r6qnKvs6+pycs/5CSljc2xV9E1
bF+Yv/N+RUdKnBEH1DjE0A69cXGCaPDkuZA80knioHODNnIBBH9aPeIyNgaSlndhKJffYR4ncnkd
79aE/hkTdE3/p3gZwMIcgS7cJCos6X2Nh/hP9sYQWLM7rljnTt4FBPwqx5vvnG9xkDvRFS1qoylQ
Oq3kRkQlmZo1bUUqOEVixDYHJisHSSCnU2b6dsO3FMsRm66NMqcCQHHa92VrvZRJBY4KpeI6LCEe
1g2HM1cPfAIFQaXUTyC3StzsPK/OBvsksRjbyW8X2qGWfZm1DuzLsQBFNogjxO5UvWUhtA4HaLYU
0aznv34HuehVGxcQ5jXpbpVceRtz4p5PmnWtM3K+T4hmBPM5JPavScuqz0TUu8BH6PV33a6bvsdZ
tPt3A6dcP/1imifTMLwbvcdTc5TZLlwDDKKnQ/cKEtjYIUWmLkz0PeD37lqMpplfyWsw0hIKiyAA
gzQZs9Na+QNxZy5/GFzRfz8q3bVj2R4nkagosmywPaW/spZodmnSIRf7NlRiTevI/qkguIucljKe
tGIrKBdoYkLomzBRiuNqz8auUZabhbVjFCnsZVCov+Sv0ES/Td1XBeiSUb8EhFjpIWOFsdFStMk1
7E5Prh/pC4QXPPII5eS4GbbhTSCrC6ZzU6boxK7U4V/4lPEqZNRfZOdKk3kJtTD0kN5egSqw4uJg
wnevkyHwECoiWvInt8X8sdx6AHodHiluoGrTLhy4hlU688h9B5US8/bY5GipjulswaNF23CE/V1B
bHVLQ+WC3hU+sNEcirnSg38+LEuMXp7En78pcJrdwc9KfK8YZYwksBWTOjmvdhEpVNwM5Jd1U7uW
vVST7uvrb4DU3De6pgbNTAjJRqT+9L6X5766+ymLUNZ1qYPPwTJVlTzB7g/4NaEcrXjOcJKq5A4N
eOyV1bSZQ8Ps87ZI4xcCQggVk3jMsjxrh28C3ll8+7Cad2pDgssLKb4RSGYg7fsWmUEn/jwl1rGA
kfct2cuYAGg8grIS+lI1/9jfRQuoXBaPd0pDlnNuobbo9D3brTKKE8XJqXa/dGm4WSHAYTKa3y4x
EaOlYxalDdUAADYCUUrlA11DTrKcEVSvL5+piDlL4obw5WOkhKHfnU6HwbjUgHLlYn4t3xBf9LkS
UWf+zdCA5ndmBTLCsXQn9TV79+IHHfpEC2QPNs76WH6Sev00G2nL/m80iV/0kGGynHr9W2xW7VPv
anC3aYfBPvv1Eb/GtCv+X9jZiWn8kI5y2F/vGW6C+plePoR2fsWDdsquKLb6aigy/DI0iZWS5Ze/
ggbIlT1t1PK7a65IZ+goj2J5IhZn1fjdTYhPG3cNMp924mMre8i0cyMJjsEEJC6MGbyw1ebAcOLx
f/POtbZimFvI+NO6eu3hrNfN3rqjCiVKDUPL6e7ayGJTWPHeqIufSR32zJtGrUWxonZ3zjmU2ckf
T6NXfzQqtDjt9B7H2oWuDY+WWdJp8KcHMvBWv2Fx05aCUzvliRbVoElkBm83n86R5mb4ogMHfL89
nqtTMeyjbawaXO++yPX7GHP7yWG28LHyX5vDFREPa4TUVP1bmeVEe4dM7cdnscsU9Hv5ecXFNecE
2AVBAdfNaidG4cU7R3RLOeHYJrEnkSqyFYAnJKU/kvIcSvlLnXI0b6xFJ4AEHVPnNRSBarjfqQm8
vY290iS3+Ov+vdGLNLD4GZTcriFiLKSYj8q2Eq/dJ1WnaVvY7J/sSo/1h+mE2e8xogcTIelbuVpG
bQetvRAL/7/W20u7yMHqJkAB4zerRzsQEiOy+2Ga988zsw0aKoglVr/HBLKox3xpdnmuDKxAQW1N
DMpVybG/V8bNqR7hrd9CtyCtdzHsDsZHgCf0AT6ZNAnngZhcTFQf9VKFYmtrEtH0Jp4MH3AWOJXf
h4mywSZY8G3a/J3rZN62+WC+SBUqbsJWQ0TdooBudGRaP9pF9VLh2Rg+fw+jsO7z7WYHHIK6gVys
T17efpo2qi6lLUY79zkCl3BqMmicX4gi7DPZgtrhlVlVY6aVlHz3hg9LG2Lb9BgTJC9i6Pus7sWC
Hd1s8KMBlauWh8jhsRN9l6OIut1StCQGyHkgrUeGVrLQAefJBM0KGvSfHZvf7Qj0hkxTNtfAcGto
rJ94Zh4cgntAxAkmt0aXPEWkgjqU7ZGXzfuRAlLx+2KZYzIHcVtRsjuk0dXn96h/fQAqgOfDyVpD
THPUg53vDDFKQxTYjtcOvxLWuxWpKoUimRgENljt6MK1h1luCcwbaEJRpamO2kke+/sH7KJ9Nr0d
6n85/sT8ObN1RT5KoBPfvKqvku1CjvJGGQ0CDU/Y788/XPNx68I6+xboLP8BUvce/huwr9vnAaQd
8hAtdWuqyktFx+QheedpN8HbcJdImErmzULuacNsS6TsJecR04K5aLqzWCvfXFRpV/kozOL4VLVy
wrfAXmFy5AyAgoXL7Osyl/Z+8npKQBPhR4as0PZpliQXTEhQcz0qTk04dtRWX9x2CbiLQrn7yuNA
vQfoC94Cg1Ag3S6xX1dh1FaX4/Tv8tLNd8OAaK6wErCuRiZZC4CXXNGRSThkk4W4N/l9/NtJj4mL
LCfMFJq85D2gz0+VYVYqGR9jc7VZJpmKwhbi+MfAq3QAKX+1ur3pZ9+XIxgn8VxuuYpr11K56taA
Gl1IlxYLOSLT6X4rTWrMxXuJQP6GKY1n9zmyQOo257x7KfhZWmaS89h3UVYayaMtjRmFDQbXlbsi
hl0bQFnD87w11+lnZurDRcpGMthBFyWWbYyS3GRnsLU2Cw0u5M5tTNi4i3Ig7BSrbFKbgRhurTZQ
4gMpOaoKSem+NPXGNDchFr7HVq9cUEPuAiR6YQCMl7rliFLvOs6igyxvJrc/dtsfWvmAV/E/gOiu
5GjosRuzMBbgO/88YxCXmh/T7r9O5IroXs3AzJ1inyRh+AN532c9hoj+/TrJoAX1yvx+FZKcrzX6
FHHtiPENvU7mVFhfIgjJhb43tJefTEVIoFE3wJySwt2MeO+lPvbPTb8uNj5gDkQxdeQuef4Y1hdN
TtDHEoS+jdEV1Hdc9kc40W5y1ZCRpe8jqsW09g7/5/tspaaeP/IKJxh1jZ1zIVsZlp9oMRfQX2iT
74vgcdYgnI/jj8lCvyhwE8MYUT00uAQdhjA712A6R32eIXxKc0EkIvcBcw+ilTsY5yDCmGPpjrtO
ybPUNfn/l/U2sKUrqNPfThTL5VYQhKo3mtaXj90XwQgFhbltPpQRPX4O9YZ1BUR2/gPekqtE4uQI
JeN/6atcf1FkT1a5SJPN2iI0EGb0C7IGmu33MeyqYD7yqLJM9pr4hsvqkkv5dTFm2QZuybyfEz74
669ebYKzeag+gNgY8DiO/3ShE8FRyuZlt7aBJ/rmsAv+HlvRqasLewJNmoVPd19Bc7jdVpuhXpUH
HOOCy26k0aoVWSTIluefYuiZdxz1VgQu1z7+QITRVBZ0VCCW+a/rCZaCQgTjBV/qv0TkGra6JXKZ
HKNyd8ZTxu6uc0ldMzVuXYFp2UUBL4r9Wab/yF4ZrAdtozPO4yApJEe9Z58wkETWR3pE0NKbeObd
W8ncFvnIN0uf5MKVRMjpJhR5yI/l2SzzRRwHdp6QeGPolPXOpZ2jILWny7onH2OK7cdD6roCi7I1
I/yaH084B0t/4iqFoX493gjUYRokdYXFvUcPYv2+8P+0rRa+repGlIZ0akwf6lwjpPzrTM4oxZVd
2uRwXIlzWyhu0Mb4TP0qHUynm2h3WQwzfpbcRiDZTA243c2kRC1CdcraizPUXudz0jgh8kA89puz
5/CXe9un+9CM9x2wwH1EtDipguDbYrf9cvtLGwWd1XL/Fw4SAW3yo4X1t7+QbVaGlACRawNewc+d
qb95xwHZWWEC4yolmxIJDbPwL9eca3yE3xjRzNsEl/HW7Q66iGgs4jLDn3mHKvMcHOmjZuCMwwMa
zQtnEPGtOmn0qjKYCYhD9zYeaV9GHglDnZDY79cI3+RevvMZlSP/Iwm2z+MiOwlTrszMspQ4a4W/
mY/2jdBSXhjdXb4u8ZNMcGqR93RkVrAbyQEtq4Cpb+YkHX1V4YiBtdwRw2Z3sSX60pWKUKNTia+i
yDdJjv+jxngJ5EkHn+d71r1TnyuZ8srKMkNJHyfzk9/Azp/3QYmZVGDDJqrYlXBB/frS3v35ha2W
U6Sz0cB0z4772J9cbF7DBqBueeo6/FdvIm/73r+eUMSgGMdy5qwKYe0D0WAiZ8/GYp2VJZgLYydD
5Dj4NoJIs8fk4dvoQjd44mQAjYN1bkQUbMtjcc4qxoPSQuTjvNPFshtccqFglY2FXENbxwpGqwnr
wfVmq30kUGJtqUY37YUQmxk3lVJoTUSydaXcBE7bGaayQG2zYqyFGx+OQac/wfeCxVjdOfWKRksY
YR3a0ecjyrLXGkSa+WmDWraIW5l92IP/MwHzsg5GexGxfsUp8xp/sCSwWSg1KJ4JAhnTZEa8PMFe
f/RPBt050Kc+OxSk5bW2dZpm9msSJwnCN0ncw6X7c+Fw6J6wImqZdqNt0XeTSzqJN7bTV8spPE1Q
BltEAmLrsAoUOGm8DDsqjfuqG6F2sGNtv1TPcM0jTsJA/qR2K9E3H3IkmPLfT5mouSvZkVvl3wiz
TTlmTt7CqXMT2WiyNSUvvg2RzyinPTQuF67RKS3p6vWA1753Oz3jAac+2AVLUUEiKqdR1Yl6/r+n
ojvMaXcEoi56asmJGV2IxSQoyqNhccxHksB2j6mLo2ycqkN82frHwJrtlaHTFwqj9+8RkO84EAKA
/gcuModwOvHrCCVpjiawv4nsmtXTPjwycGDVVRJMKvO0/Vn0X8hM579SKzYhXXLX19Y7dlwLjCdv
u8OGgbDSPgIb3R0rz+I+OoewUOCkDwBqwx5vHIuEXmjKxdPPJYU0MxcrYyYbf6krN9+FmhHHmQ9n
BDZg3w0qKrzKoytsKEXI3LWrBHg61BW1HswCj+3wGm6tq9Hszxq2qFUMVNf723iMjq9aW4FRAZwZ
kUG3UGwVFHM1JZfawDKJGAlBhHktB57lPWk67jwcOzsW2T1+jHK5JBw5S9SYBq0UsRmBeE9lbJRW
Py6zmcLtc/oQjmooyvFzTZM2+VZK5w+URgOOO7CKbxKM+bpum9RqL5wbVZGGV3+I2kvNYFYvJnOb
fmcIQ2Ss1es16tAaErAN1oud0oUkoqCQmJxyBGtSKRcu+iP1LVQK/ki16fEnMPkbjAGeEoI5YxOE
zgor0f/CMjumkcHsqVeW8AWth2U5t+nOrD7hmfrmWQI/5WQ56gXXiMbrSJgpst/ckQYYkIWkjXrs
HwnewqNrq0pAQdTIWZI78aVKBEXqRWQIdWxdgu/e1mXIzwXwG3yFjWYyzpdevbV5nqrmnQIY5ygS
NeOMIO1fEBOp/jA3ESeWfZzzkPRY1aDpS5AUKxCwN8MP1fjkN2j+pmPXelbioGLYwLchmgiEnxs/
E0kZ1uEzNJK0WoiEmdLH6MDXOi6eFBjDWlqM5er5A6gvURkf0UZjvDT5EyfM8Y2VNDnScjtQze2N
cKL8cB4HbRsXTYAsu7fvKq8etwfHrz2SeHQFOZHI6pKHgM/z+aGr3Sr0NTZDknkgf1o+VJ9pR4uv
/qktHmZkmdq+tMOVOaVsn8vVYv9gt9bFBTT8Xi0f1Ww/S9lPexABDxQ6QxiOtxGtZtnT3bK4xXpC
li75hHmqNZ2ioz0zHpdt7m8QJyqkDDvfxq7hD8bUKVGUFGB8ip0YB7cmuarb4z3UGpZJbF7UekYG
H/4efJ8+AAHTBCm0EYOck4PEYSewwbATgUQqrLk+aNKeVMj1cL8NUYzdKOO2Bms0YpiAmLVQTwiT
WN7L/0adnVlf7uZsZ4oFYpl7muYfEeFss4eqvBtgnbxJpgXHTJ07ufOJeba7+7gTrXv6tAAoiGT2
0QpSn1U1M/WVMV8US+n9tTlWgoXL9wjoQPFltRQ7Mk9FDroeWuMbSt1zFFi1tU3Guv1OgyLj1R+3
T7K7iivtGVceGo02vbxCGTwz9xTeMxoH0RG5iQe0sUq2/JG0AEs0LH4C1se4rgdPSMgaZ1d+wl5h
jdXjJXMMCadAuK8FZSuGxniOduzAyvYOKFtvGwFFuL6FF9GFGUIW2QcrxZqdgphWYfxfto1/jGCZ
jSJC+ssSScQLeccdeUcrXKJAFMPvTudMS9w1QDxmrMRcSljG8lF3JYgH/TAszvCHUIPz6s1ci2Pe
6fa2BBoD/SzflAquvFq+ISzk9yow96XSY5V7G5flFAEy3vjtjEkMc8Q7LVmaa+qacnkT5E9v6AGQ
1arDjJce5z7y6FOmcqKavJhAFuc4cSBKyODHkm6XQ4D1QG4/5rEW7yjN1oA8+s10tOnT5u3FGwIm
tC18qt7JznviGWxs+qctLBoKvVoxv2ntRlManhuUZh50awacRRi35BSGCEAF4+Ezl2kAVcDIgxg/
m2b3xvf4uZY+/LIio2rqohqyWDey3lsVQSyVWHu16vbNZAV+9ZY9RnSd7xrW9mpB4sNXPnk5rEyC
jvSETwmEOT0HOHgrkKX3/u1wLpplRFjeKgdiNs57OOMrW3jC2fheig+VGtC6dD4wthXQhu8UuS9M
XqMrso0TGXo6d/NC6NO1Tr4gdJGmjcLNgXjS+G2JFHty6xccvbJaNzPnQ/03U8SMjXS1zTGEpwjA
RolZlzbUZsc5Yh4tjLdkKf8aKoqWyjNHl7bNRIluxew7DuOPkSvjhQxv9hshOJ7wvZR6hMAY7cc4
JjZdBZ80RZov75hXBLHnWOsxh+O3Qx74optdl+aSOazvp4yovN0h3yfmhLmk5pe3TpMpTId4vXfG
8YH30i76ycIAAPWCXSEWfX6PuC9S6PDcDAbAiM9UITmpMuGHa0j/TDbaTzYud1CsS2lVUnxYoRtF
rFntfvX0brWZLl7seJ4pfRJ7RBfRXJm5qYMUkNRxtci17vtur7I+yOYjlVXNkXe7eEHg8NKtaxNW
Gcb6nzoIJZX+xf1XISn4tpbXmRJyh7/GrJn+LQBIzOBXXzFifM0gUXG4jzeK3CiLPr3PfuCwvAoI
nv15YrzNIratsufX4lO2fWznbg4sQSS9BlFNQ1QY2G/R5YzEgWm9QenSamHCoXEZWnXn4Q+eV6F0
HMybxXSkdCSmYHL28hwWfqXPoL7U5X9xjbiOecsv7MVKrk/Cey6p32RHTFpSh25n6EVZukW3anpP
62Aga99ZxK169STfS1qZXVC4roQZMmHmF/WR2oOUrcZO4ju9SsyLkAtiuhGI5uapyiEIUiEr67jt
wD1ErxBclamer96f037Yd1WXqcbVrIMy0r+lwUxr72Qeyw6TtV0XgBAgwJL8Xs0pSD5t4YcI1ZHw
CNHo+4yeJ6htcKY9EfAbDkqcQtLDKeJvxBoJt1Q16RwW4DIfAYB+3/Qfw/O52oQleWAmTU3jU2gs
IXN2jLMohgqHlug+OKQXRHmQJadg4gmst8IOUPCNhJ6Cff+BnS74FhtqKQf5o0CNsw3Vm3y49lx7
ia82Cg6qQ/+Wbuvs3S9VOi81lmPGiZbBOdFsz9SbR5VegWCTmcD4bEFiHRhNa8Iyu4HmmBPdOBnT
wcD+O8kt8+f8DnY1GJi9aOkVE+3bjoPDTyDdo2BU2OFvdVzI2yx2AwFRD4TANYlBuNeELiNWKLBJ
rxki909iIuuEC1OySeEnMwNajHKWL70e97MbcCcffUjKoClja6TR0DDs1p0e5xP3eSp2N0cte2Gk
Ym3obvomdu1iqS3e+BEK08HCZQQNAptNekt+3XPKxgWADB5R+C+rmC3It16/Pusrdh2TFRiitmRQ
vkPtrfbotWOveMGDlOFb58mcBTMpehQ6n214kQ++4mu0raMhvPph63FfNz8ts0+EljUpdDCZtt0E
nPxfPi/L+JCJp6uZo1k57b9Oq1krHbxDgj+hIK6/nEAUgF2nAzE1HQ/uqDKF74qF4PU4BNW193Pc
UUvhgu4n5L08kiT7iu3qs4J/RD+2WatQArdYrBHfhmaz1FeJMHqPZAiPSEGNkDg1a3dvzsueRBjt
I9dPlUy6tUEJueKZW6cq3WVnGwiPjj73sLvH8pte+045jca3gRUPYhNPzJlqJc3LoZR2HDl5c7i3
oyvEN9U1xgfBZEoY8tz5+Sjk9MFpI0sr8DccAiTQiLHUINC6nW1YD8ALOdA1fYjo7Qjv+R5GdsrR
bhyrqQuj+kvH1bJrOxvV5fHMBG1r18yYXhAqi1GAy5whNSPJvrRz9Pl9qkchaSF8lUweGkWYmBcO
E8q0uxjRJ9hBDEwPnPARWd3HrE3PlajPL/J5mUnFU0p2k+GUEAPT+GlqK/amhgtNu9ctQ5fG75k3
JnWeVEr0BVojxrji5A+HnJuxIumjvqAGMEbp/VHKvoLjEh1TRPco6lv1ptB1Mf7ln6d+BQHvTy0z
Q8Ortz2GkItxrrlKOMjctNpNBdWq9BiglLA5NIbrbtke/AszhimoyLXxVA0N2gN7ZMmR7kyQf/CN
iAFrlVqXaN4UN684eIg0MQMb3OSv+gZfK4oMSxEs/IHWaYTauAfjS8RtPfzxuQ1JB+VqnQ0IxDRa
z1eu1+ImtiQk3Asv1YUWoEVNDZP6CiAOtlvBvz8DkVFldAK7zuGaiO9xMzjgEvSzWsN2upXEUjWT
iIHknoJ2g2i+YkzfvZOz+lW8cMBpKQn7DWeZkhgQeDMfrQZNhIHRieweifsksXvBUZ6xgTp5mvdn
vMERlkVOUblwnp8M0rFNP4+WkVABEsUk9HltmS2yZqalVnbK0mE0B2Jx6oNaKgWg4wX5YkS1IEJu
psshW4FdFItQ08i2YYciBSLXCbUhaNFLQDSsj9lVvCRmtVLA9qZuitR37HLBwHubiw9NKxZoHxHl
Eqt+hBt9qrzQaN/+GJHc+knF7vJTZjMz4DN54/gQR/poCj30MMZZ8RuKs2Pv4yba73/17ZEezsl5
Vgp2RyoXhMgQjPprl6mDzsVBPt8vE4IyYSrE4swjT69iFmTJxtFiqAyrUvmfrE18Zysi6il/orNU
91Lyl/hbl/FAjbz4WWMEJIAWgphpOaj+9HEywk2qp7S1QDf3jjkTbY+3SrK41hOog+hjJXPrNd6g
9zDuVr4O2JFdX8Zl6f6SWqlMtA/ZuJ8yDQgaQ0BSwbq7JpiA97SeQLi/muDmO+6lXr76qEO68JSf
6kDK5KMLXFBlp/yohUjTf3zzyZ3DnzrP5Qg/A8eRpAUbFwFMmifbARjQYlwJQKLM808d52Z7n7wG
z99JwhZ2PrRT7XjkkUCu6xBKPQcsoOXfX0gkfBkHsZ9Cem2WeNcaHQXSz/zyQpSkRr4CWs4w8hVm
j0M6gxwPuTn7ID3FCfohpnZDLFqObGYQUH7MF9Bspoe2xf776Tb04lY8nOX8GMSz+UBgrWiGxU0X
Sn85DgOPOyEuAm1c2L29CoQdM3UpoLpcv+EVMqKW1tn+Cgp/RUtAGkBzBjEtDTUsrXlJRXRFdrV6
KnAVYrjwdCM82gyHqzpLG9NcfB7TGK/nFr9E6mvPTgnsGr9MVOC0iAVDPNqXKgpdb2w1iL5wR71o
cL5v2yqnMyy9BconGl4EpNUxdxSsH1X9EE6FFeM0Wry6hwptgpSglofxrDAQgBC7fCToYwBwb949
A40noR9G+7YbhrSAfv4lg/1s7M7iaSrHqOvPBApre8ixFxqzwr3zsju9RfAw9LuMy9DxYSU5GyGo
JErYOcjpRnR0wJg7jS9kJ/5gEVmLTflasinE/G6uFW5eppibEWetWY2fU74piFQr7mBZUxgNsLWk
2O0nPrUVDZ62fd92Pj5qgvNCpkwkJrATeXURm1ry26RVjvSJMlA03hLbFn6F1yAQyusRt57gsd4C
E+frzZmeeLv29AEACAHTqM8RHXfKd4fHUcZ4MKQhODPBCC59cTK/Nk8tn4ZCb2/GYu6Q06J2cdCM
raSFcusYDy6URpOuLcYfBmyUXAh///2C9EErj2YVp/5n4MKqzTzER874fdVixEAkILiiQKn3v92a
f6gvWY2WvXBjVNgHgm9USF5z71hpxrTMlOk7R9hZQLunyPJKM8GiB2wfLKbfOeViIhGb7Y+DIWc7
hvQxhhCiwvTv7xXocNK3n4Wlb211rpLnaNfPhdAk/57xdUP15HeEL7QN/D0FTvLnfwKmfUGtXF9h
ERMcHgjSPvWJnKr/o+atNfeZDrzi7x/QixMKKt7EgVFVvZeRhUrWS01UBiHobDHJpBUJg3GrmT1p
JqEjiZUn+l/lpiUIsnzCRUv7QG1gmff3Mj+5QI5MSjTKze+V5uAnLh4UTMXOCjbgN95jHSjb647l
65TaJsnHLvOzzabm7WpaNQiFOuN3/SaAHJ8eFKnK3j+C6Q0W5bdfb5x6YHcV0AXOvTWhWhGPctvm
TMZIFwDYyGyQ12EoDtafztspCUiJmwDwsVglqmCWKrJWQOgL0SkR42EpnQoJZ8nOn6T60gsHAqHu
RGXOwWjl7PYL537GdTr+6nkSoHRAeXrIaOoEnlPnxFiH8OMG6zH2L8ym87zxtJ3b1055OQR/xyoz
PP7SiH5QDRBLuj1AVpACYb7Dywijs2LrgVXN5CD6LNWBlWouGHGVwueBhj7vQp3g6Mw1Hcvr6W0Z
mpCR8hjfSK1PIbXqmTeKMJ3gzLXXIuudVwuk1D6pvUzWk0jaNlWrk6ALxs4yiTnx5vuFs18r12y3
kNvENzqGfCoB8dplv65p8XBttiU6fCaNXqFcFjYf+hw89XBuULnK1/xdg6isjZlR7w2wZSgd52ky
3rxguwx3TW8Lq/na7p8xI9z0s1ThuD5VIyD5xVrRR7M3M/wpljLtu/Lmec8NxT1p6RQMerHQ6xNn
ahq/CZQ5HsPBkipg5qjqQ4BJ/QX8XkC3jGLvgWmI/XFsDhHgv+9WRl088hhioR1rQJpBYWN5XCMA
6Wnd6ELPRRckuqZaAOXVFu/tGfAkdhZzBzLGO6i5yRokQg9c0DNMPhNZL/ncugED599MkXLUCj5/
ujcvnbzl/xraLMSW1q1stxM4tajq324fidPVG4nVUhNKhg0MEgLTAKyko1d9ec+Kb6VGmrcQes7J
8NixO9v8ohIVLL0KFMm4os/jcdk91Cdw9A8gb0D1AtOsRDYpEjP4YVWxZb3xXXjN38Ot6O1+dfKG
5jsB5XESO3OgJFOsYw3n/MI+oTLhi4mBjxaSsHS01bBtk0o3+ExPJlMyMIL3+PVX6LeIgIeurQl5
L57X9inpan8YGhCmLVrYzY8aFHbG/zxUBrVuPHNL4tqOcxA5YRtk8DZ5o+cQ3+f3rCHkmBIzooWd
sYBZyGZQl8eH43EH6YXZl01ofZou/sn87BEN1jvA/3i5/fKLjIF1Trcucs0m2uogGC1ox7N+58Qm
/I9sozqIYPi1pmFkc0ZJz917jZm9FmDE07iMp6CnMvkPpr4vVn4L4cN3lJy9DK46HK0DUss7zXQs
XMrpEqKufBRuxgik2kRiDZKVhMIBR5yRWrz7yHJ2gv5oYDJbpGC00ptZu8xay7E/36j4nhtomtHX
RYCj9D+3avKxxSdxwxYvdRVf8evudy+NpsK9pdr1Vrx9Ext6klPRRUJfMJedHbhpu8xPkDFtcqVZ
OucpZoJQsh3rIjWElIaGQ98paBqgaO6TPq3wf3FMS1G0YXw9CXMQIxq1VR/CGLG9MCP02/EuC8+O
rxw+NaYrByYv38sGGVVDRu8cJPgM4a1CcDQUmZkQXJsBv3biSEWVISihDr904bhB9FEHEvpeLrcp
KnnvPrjL7X3/jTrzQqJWVDS60gdDbostyUPTkYp50DZrB3eSu2NEiVlO7iH1+KyXgxWfh8i86g3A
VaMAEHCHwAzKxuKdVJXy7aQpfz3EaRetYXEyvu2WwgHxOdfSpJ//NGVZj99IHTPAejoRdm+U0efn
B4p3+oKop/8m7mwWGQn5CsRNtkuQt9T1DdTpPbO9lwX2gCgEYFKMIAQsnu1fXlB9b56kc0OX/pZ2
nl8akJzpDwHvYYtb4uqoRYirzDzikrW0iGBJKFnFXt7Yf0j8dIASMOCHJi4aVzgGwyd/kVxmcY9o
0bTt24NDURqMUrEE1O6xnRMJQ3OLV/1jHFZ33IzntXYqr3SX6LS0CWK4TLuCewB56K2NWW6EA+vZ
5Vvrnt7wNrMJBjH/rD4E8J17U6e6RJwAqqgpK6e7sS7VGFBBKLgVqvoMwZuAW3lQtkXaVbbcSi3T
abQJNoxmk1o24iYwDfnQDOmRfl3r4Nox6YwtVPN52reB/hQBjRYDgOnzqQnEurm3OJBb2nDY7CSh
fMHpDBwPW4uddq2X78vaS83Xf4MITQ4R9UB4CQxnCtcjgZQQfizReG2XuDGh0h6cgwP/sRQW7z3/
/Y4UYtYdeLTj9FqV7VFMjHlPkETtUbbCueFlUs3XTkwljjLM3P/+UACV64Zq5ock2f/3fOgS5oUr
ec+KMoP2QJWkxPJc5e7S7oSVU0JHEud/lr6yMwbczjRrDeq4NUoXIPmbIY/hQJjz9WDGla5ZLtLn
u01uxu1UipTw4NwUelu6I2Ee3+6QQebZ9GL9CeadXQec4nzsuumryFZLLLG9gfwQTK+vmtIqA471
wPSBTS17753y84o46ZWJaWhMKUsBCPMshPWhG1iLhHyRKs590ZLJCKWyW+NFAagc44/TD9SOp/zJ
ntOyGiDBvLTG2gL0LslzER0oAr/PP8mjAuGjHdpkMsmZLaCEL9FzATnGTsxRNNz9pSD/itmX1WuW
m9RbAxMu3GstRPHKeUi11phwMNqB2B3amSkAXH7PbxBlmB2wb4RlOjJdAeuDpHfbkAqI8VyNx4T7
0Y4slAdnkdOK+Kc07D5tWgHuFO8SOOAQUC4eIQ0oB7jAyXhB+tuVu3U0n0+bDR8hJTTMCKsDiUUd
az1XJJWCh4sIBfrhOGijMJpS7DILTIcVgoPGy3dSCJvHyHWQRkRF7U56ewM85W1DWk0/UQU3mcqo
MYOFJQQFsDzbLscbh4Kb0eXortmTpCQNOT034F8bGQy77doTM2gXgMDu/XKaytGjx3azxl6ew/Nt
aEvHK8uyIDsplH9ge9beGByGO9x1jbNoLqeqxUX4w+bB4plXZbzltQeakGf7y9eOrXyjALEZyRd7
/8l0dg0zSXK6hNgfKVSUmc+8hvodEI/54plyQQsylMTliLHcNuHxoGW+6qyupDKYJ7iP94co6ZjO
AWfrMIB49YPH+K3+TlB2yl4nXLoPmfhK802PyoApEwwuaJLhTDJyvtjhqxhVP+o8m6DbpAuuB+ZC
4Sfz8WtT40siKdIm/LkkkuhnC2cRIT6eJnKfy7w55/E89f5YZgNk8gWO5b7xal2a8rxnr7NssOjQ
aQldTkdOiNaZPrcfhSr3F/RE8m3RAKG225kSDSkl6HDEv4paF9GXbC5m3gmZqfg09IAZlHpzTU3v
TPLW2zoMmteMWNHy11vV0bGQ3s89O/7IEo+xC2Mnr875H4DY4rAzsTtKv30bIXkNmmrVTYSkYztA
eO3g6BjVUUjQcFB8EpVCBLhDGcssP0IPkonoBu/mSaSeRvzJM7+nUMt/Rk8LZ6Lus9+V1lXZVpac
dM1GPt6MJlVhLb/Q9GwhdWnxEeYW5Gp6VmfQCXT3GRLZynLy5v+AvxXgEeNyZjOdiG/lkGQa6TjF
BiBAH6brP6GB4OVPEf56BzLQ02yWWnqtOVP4V03n47zBWvaV72d1DxOIwYGQLFQ3/0NPkZcc3JPv
31zhr1X4nS5WGNFxe7pggLVGvhAgHItTIES/mO6oDU+yW5PgdJQU/pIc1By221bkhjqi1DFk3hJX
ZWR/PXuz9S7kjRWtWW5K+09ILKPE3ixcaXLOI1yzfZG6/XxwpW2u/ip9I3qo4YOBawMP73JGp5qP
5B9Bwqb9EpUGki9s8sa2f9abWjqtOFHqJP0VDVulhoe2/X7Rj11BC7kvR9JCEMXzaR0czUWa8qbt
UsJEu+J+3sMbthheNgRiqQXoVxM6O+jM2C90k5X5MteEmmCPMA9GCSjypiiihVQhrYEbpbCbiejs
fU8smvleyYLx76e0qolsY1y8cShFkR8qRNmJmsOsqHt2AQxvIy2Ko75uQsdudxFBO7hUl4P9TKEO
NHDLh3GJf0X/Eb+VRxDmM+BVjqtZxUGV/MFIdF70Hkr0IeI4gBhearC55pNX8tKdedCXd2hh/oaz
r27ORReJcAt//wOYrh4kVQn+h1SUySJH5bU5zvroEEp8zZQHRJLD9GtANg1OHP+o9mOpptdR4E3K
gGbUP5Kafml3xCnxhDEgvvYTcGmkWMRbjjaN+Z1id8f3D1o63PEGIX8SKgn4oBeT1AXGGG0k9+S8
uHzGIiPeVkJGvIjmSs4Y00CpwMwXt3GIYYebhLtNbuKkLofciYgFxDCb8O2fSBeTSCcA+2BdehnL
pU/JuL8aF1DRsKi9rcgtT9OKc7dM96Q24tZs3Cyedcxp5gtF2ZF1i8fd+oghpC4z/OWEnpsOsvb9
znsVFWbWB46iWNZip4nCreH5rynMe0tou8tzolQq1kWwU+Cvh7e+AXsjxqlGItVyp5g1aS4jketV
8ImdU3vpJt6bpeTWlM4J3xehn/k5QnMqRtpF+dCL1oZS3adx25SUpRaE15WyCBNVN3Q3F6d9Ss4l
5OGDBuVjJcrktFIWcFJ2zalNAaArXK+Vf6sq6ABHZqhlOPUSFVYwOm+eSGwlV41j83s69CfGLu2x
7FcL9m9AEXl80iV6KZNFWTzJN6AeC5CtXJusyyl3/LWvwRFebj3jEGlZKNlNoSRo/oimzVAxSEjL
g8eed16vF44U2FjS7uTApQyw1ZLEYiEsThud9ahOcQbscCoQ0t2OHpvsycEirrXunt6jmefzdGlf
PGPurfUbmjHn943c2o1Sm9iM+QozBcqmfIhRRzdfEf3nNQUScOQt438IpMy7w6Jx4rw4mGvlZx7e
m3eg7RqTp2/xeCqhoCRjcTIhoCVAfX7hegL82e3N4EA1SoFToOQLvUc6IOevfZ/xnDvBPK4HTG9b
mqJgvTbGfo814c6riW8+aSufvoWErOx97VBhfjkASrr1x8KKJOIPffbuEMUEADb74WgJ7JkCHsLR
WyJHitnS/Nobdcm1ZALzkh6wOzOG1QFkgjKR77F1bYPhabhQvHFoseiPaelSMJQcw6vQRD9BS1i9
mCbsdSxbUa5kID+OKjU4hZviqS++cmBWfy9jHGG1RXNpEg0jeehJVHJw8JiM8XjMuHlyUjP4bx2Z
M4q8aDE89azR6RegTpQp56wRCLfxW+l2jUh65ZvfUTEtTDY84+asIX/8rvFigesPDy1PL8g06orz
+TuIOhSNpYED8+q2imWsaBHkl87PtfGzT8qMNBRmNjqBMIhRBwZUUzIBrIzGXCY4rb3b4jlU6kdP
h4/fpEXUhmzacxRgxZjqlvA/sNRVIJkzQF9hcajDd5gP2NKvPmVVQo7lL7mJgwOc+nUEmtQy7wyn
mZzIY5K0oYHOTuyde3hCtL/fXmtVRuAAwTKOZ0b8TV0WExjJJff1JSjmT+QsGgZ6/v8aqm8ni82g
ldcxo39xusDK4Ob26XVewizrToDxdfq06lMOCmw0nuih082lY6GLgqAs0vz4UdHJZs1GnVyAPIZ4
BRAojoDJZ9WLPu+m+mSFLwPoIU0ydoK0flnygG2vLKvwhNzzV6/ZLYYKgn6hpdEOom7qWmFWRtie
3CMk0cVLhY1Tdrlez92m8quY6s3Ag2dPVZ0HJTItkQE/nD0UDR/KOFKj3X+StVNE4p/JJFkk2Rly
V9sbYEcQ2DpJLbRqURWIgs7NPy1ahBtNr9nCpxhHL3YGpYvd3MHy50E9fgKbeigCef6FT9zaxdFz
wSbDyZYNvlZ8CtOqfjUr6hwf284E7Mhn9rlqFT+kqIkfbNS3GW+eJsst55zMfbn7+zLHGa5t3K6f
z1IQNos+08mPfJfkerez8n+usmobs2+gUB3e0gI8g7EVgGCSbp//CnJBhJ/UsEdTdkFHKiX0Ew4l
ZDmL9qF2xSRdWbhYTjSGTcVO6sTUUaiosxNteSOAx/dqCrvd+7QKY19B7YyD4NmzmNqoUW8S3YXA
h8N4Hw/t4NL5ki2y+a34JtZhflXI9ODkCJzz0mTgIscvZCn2SG1FnrJ6O2SqMpj6NjALzuPo8HXI
b0nH2qZRpVboT/lGo/mCJKouK+/fD4Rh1upJfiKZumnDqXnvkKNaejGGX5zRmg1S2wWu0PzOq0Mg
Xlpe+XjNE+DlnRZTrkKkaeNW+/+lBflbHtK4jYNbWh+d1ouMRDxItKq0WO4XAO+3SWwLzy0brdU7
z1yq7bL5gqHH8Cj4tpbxhYVg7Go0jcsX1oIsvwKYrwGcSzeAt8Y0QttxL8cE0ZV7qaDAqvanQRTV
9i4o210VerHL9uyOF3lJsADOrhhibQ2NQU+ITaWzDK7/gMZBBT1DfFt6asWPYpfvi7CYxmKBsS3y
sMx3dwt1geaGWM7KowhfdVqEZzeVayPlUzqBg14ugKig5oE09hy7FWR43+x6gmqYkmoEc91630fO
XgkIB2x0DMKb3m+J3lDYxwXlg584M45iCi3dKUYdv9Rh0dr1vLJD9ssTkay5IBb7KVhawFJTCZx+
s70C8s/CzyQadM2hgGJTSzgjE7AJsoyN8z3FK5yqoEbVkUniPdpGfvGG2OZO9kIobUWUnVHu4JWN
zVcSl5hABOhcaSKodcKkhS162fgm4pItM4PnOqEcrqCnSTxDVL6mTgwzrLgu1Rx3PUYtk+BLzF1C
1whYhJXdAolWVgCRVqIBJMcEhQ1/0qFjn/feN/iD8vqxpHinzkibHsTl3TwCnsaDL9abRLqEoPUn
v+Thmgc3ZF1in4qoIcZpfpt1068qYe62FDsIzGIRPmnoM6gUagA/3aK5phwxTjmVeA7YQ7cU0EAj
xS5fHXFTnJgDR16lYqKxc6RDm3E15b663SYLBh4gFJMo1SZhq2Y0Wo0iVmw9XAwJtl+5nIyklG1T
zcG8Vw4B7Ds9/rjpmSu86F3EcaZg0WMzLWvStwkWRjVACercmM6Z6/Jn4cuWNklj0PVgeJp4DXvd
pyIwPiQW3xigcRAdk3GnzWQvrsBYfAe0XN5+MjW5cEPa/lXWmhQ/DurTO3TXhCx889xhCVxFFScR
n/z0xZ2NmGuodBa0jAanIMS9bQ5pV7/IoAf0A62tk4L+RpVZ1TR6oBuRRMhHVEEZu45fCVvRCXma
ibU+RNFHz/OZKRkC5zJnLQ4kzyENRqx5gl/riOFY8yAE6XDbD3nOSW/KXZvARJiKQTHm1SbUlexs
siBY/C/JUfqqzn04NsOKuiBfgqaKoBF/5k0iB8fngsujRsqsAyrcIcBJZBeKrKc3+AsB/Qf6QClZ
NyfnzDkJvDNaRx50yhCqHmmVl9JIpBeFEY8j9uEFh1iHyE4Lb5hT6tyZzMnP7cLM+i5gMzFrwCxU
N5PVEoLWoKGm21A2AbRI9LeC4QumtBBo7v7UdbLZcCmTvVH8B8GBMtCYj/A/vj3FxO4wI6JDLZtI
CUzcjEx5AcB7CCmqImEyWX7Jr3veFkeryJb7Xf5U5Q+DlRApb80BKBUM3zxMA9RyVAfTEwJPHwcz
49Rf856VAeq8dV2KzbJVre9k/N+KwVw2zC2fyYu/v7BXZyGHYx4GWpw1yGk41UjpVRDTd5j2Eu8l
EnO4jJXraKluqIJEbelBwTlywjEIuRQgTS6y9NPpTpQKcwhMQF/WkSOMk/1qV79sDXX4s/rS2/b+
nuXl9SSuLrTzcb8sNLi7WS/qF+7ufc/7oQ0VLDuTbNHa4YS9/jO+FdWzBjz/RvwT0pTmYysHWw5N
H3Dz1tDuIpSgAfn40TKfxCqyOPjNQASm12g12GmEgcvlqdaxjHxJ9u4Zte94SQ8Ajvt16YHscDaO
9h6rmiX9l65DSxhkhvRpYo6jqyZLeLDAX12xvg7me/cb24/j8NJwCDfZrda4UecU38ut4oEi5nW0
QjgnphCOEfw40te0JqcirJvQ5jJegtVgudJWrFaZiHF4zm9TmwHr/NrmkGcs7ax8c1oI5SJROGZM
EB+Zceb03Rt9Ly2lbz/b9/y5L0l9mNAK4wAWbqUHjGCpklcOPGHPhMPR+d66Ki9r0ruQpp+oVi74
B74RUSOi/9DA7XARgOXlzNm+yiPA/3RNSomRrYg78nibdHBvrzknflIClYYUwDray1gqiqqrjBsW
ewp67Fr4wEf6DEg2mLOogy5n0MqbKD6wTwrRMCMJzzG6YQAS3NK/i8m+0vLIzUTCY34ni80IezuQ
qd7QIZADUbAgFSjO2Zektzqhg+AcP0H8+AhGUhdyKfcw6TxowQtue4rklVfIye0rNzZ/zqRZ7T5v
7IobmASCkZALtigUgE8tBO52h5LIw4npKQKHkDgKoSusT1kPWjJFCLENWmejuI+zzkZX7jvPD/g0
32XKkVQBV90ArTNRd0ZG6bBISFIKcLJFybGgxSF0hrYmuciTrLhuQKi1FO+Jmb4Itku8fTMrmYv2
l1rUZi7cyBfOEd9JojCCDII0YjKxMuKsaikDoojDmZe0VjGJ/7lUJs1Cr3KzjonjX97ZkAMPwDfB
y1wf+aZWoQsu4bUneLPtZMHAF0DMQNKhPVtrwIHayH8oCX4GFE8wF7H9A3947qrXft0GSxCt+lfs
F/HtTtQhgXCswRhFRKnRvptjjyggr42Z2K6LxgbAXCjs7Cv1C3zILvMX2I1TKBXVh7qavKS2vQRX
PsMeY6rzaHRfwbgz4W0Jzzj2eEOu6pxZl+2GjTS08rXCnV8xnzebE6AS5gF6WFdZyw54u4Wcvct+
NiaNEowcXRUTc33lwc4Lwd8J0nxx8oXX8beDl7HBzOcEkD22rSzNNGJ31Oc0lsFSOFuxehEScSiv
CUKTlhZhd1FJR/QJu6NHVkV9CDdWdCnxP+QuCrLRm+uhqTVfc9Y+TS+ev/ZAoutRKuzMOkNTHZ/h
WmGxQmacFYT5FdqryE8xYFnU2BpEEj9ZCkXByOmU4HCP7FVneqjW8lHhm/OQAj/QlY2qXAGghWbY
aAAu1d+JpWHWqyUIhGyE5Alyb5/B9tvgF4D/mssY4CHQ90L4X/9Dmk9pDJmZMY4jLZPkDahDJtRL
RWaQv/D92sYNyFDheMhDMmzFr5SJkZEhFr5edFHLV391uWaSqr9Ior713a0bNkCqxdcx9n2YsqO8
mZzQb8sLkM2AkEHnZQKboNtDD6+Y7Sl9mYh0C8gnAnu0FeTN/kEOrSaLLxD5fhUaA8esCP44XSUJ
mspaoVME4XbjYe3lEnnD0EYdTV1GDGFcWwDaBox9KCXWaYUMyZThzE6tpmq7Gx2aUC/vkqlog+JU
0P0P4uGg+6TLAL2k4e4aj2QYQcFP3/zh0sXBBF8XtwCfMMNhv+7YSL2o9UUMmwUmr1laZRXlwDdo
6OvvmOj7BS0XKO9glP1qmkG0dj18T+9iYuiCwwB7HQZx/KYLmVEf7g+F58bu6gYGSJDnJDBzlADB
Zvd35HAqa0S0wAb9M/NevImCRjud4AirG23kyJi0XxJjLXJ/5qsLQKpWxCPdf/SEXKtg9z1jqiWK
/dleyMzg/+emUdAKbOaPiq9F/Pdixd5XpDlsD5jnateaDIkRZZ2dkQ9UvT8UaGE/dsoEWW1E4r3z
51uMrw6/g+G6L/jtmioKF+Scs5zxFcc9KOB3NIpz8gB8C4n/81AlEmxiKEh0tzUc78MWNBNzSU+A
bGFXu7r9zqItL1e4399RP9OZY47RfIXwj+HythxYM7uW5zliOlagPzf3fdetnBehj09eXRe5lF03
ooYQDlZpf1+B/ojW1GFEiwbSPLSAPshm720X3YJaXfp0FbhvOLRhI2L6l6LEOZXHFC/qZo/ccvmp
1BIRSiZtmq98NbIXms8d7vlm1dvAKftHsFef2Rw+t2nPTqpm1/Ukh8z28tdH/N9Jtt3hKKxLCChx
RDSm7XXWoKJAwo2qJfjYo5LtQkbUgat9T7XEsJo4FFwf+4NhcDwh9FrjHjwO2mvl04ct6De5rcfe
CJGW0A2OTkfNCEQ2ScCtY+BAxKHENeOEaO+U7EblMHlehZxKUoMS8ctGhKMEX/mSZJWnEK/N71xM
b1zSw/jX9Ll4VvGyyAXDugmreILGkD4ZEhHcscfEuN59r8eT0ZudgirJ286MB2MxNZewogwCKwWa
byD5Ms2bFeu7Kk9sd7S7Po4891BJMDZr/Oy/2qgWnRuqXga9Q12NTteaqv0e1HXtGYcDIN9idQeo
H+/mWyrpqfsonHZR8s6VJ7kfN1EsiepjTKpvRIrEUCAGsErwM3NezrJJrbF5UPGWP/aGYd8XLE4k
YUEerpdRVqLCqNg3qiywGpCGGpb0fpgPcbCYYTCvFua/KzR/gVGxpVkwco43Xt8+M5g0F2SBwgFE
C/H1x2eJFDikXZHbMLgAm1VB1Ws6WbF0yYcmVXeQn8/sGrUKZVyuXHV+FJ5aBTrBB5qPoNdcf65W
L/kyVxMOBqIvBOp3q4GqfUuvFEVs0CzhH1n2s8e/OHZnXJ7toDD5InTAJCGmVNCWV1Cj2j8jXhzw
EPc0mCOnIobu5tr+HguacA89B3QzKFLsG641enzBP/QeEt57mgdYRBB+brVrE2bhUQUZOdQyJe5O
XPGSfmn/7LRUKFBycxlLIB5wgcEQ+1tIaX9hUZBABfU8QHhphoZ6ujoFMIdpLRisRICNaNpaXXu/
Zi7fTxZRqBpKQa8tsRZ8xp0V594sFRcuseRJaN1+D4258mbfNIeOXQMtXokXkzV0aUA5m0Jp/I4o
1XoZHY2///Pj1Hcrp3+QjOBPy52DzhQp28L6dAr35UU2pMUatT1STQhmzxs0nTerqT373baiqRfC
PPRCbyXStztmTd1R+Y1FJrJeMl5mgIj0K7mqA/e1WZhPT7e+ljvWWP89MY0yS+juiAnzf4UlqtAJ
ea+KirvnjJbPXcGn4/eLGFvuQQeyCA+Q0O1KUU8s9E/nK2h4ZdY7djefL8Yx7RyYLUMDUVpXBpjU
cOS914AC0PI9Z+rBtM7yh8lolNeV/B8tGf9NFNRxV0bKmBwLu2VRbGwOhKJYoLw/9C+kEmS6imWx
JN+KJcw5RZCDgK6UdKpjR4q0VfWPLRHKKY4kiENyfITkXQTcSxdiAEwa5rDnB3RpcPYIFHB3S4NX
VBHTQxxU0PoaKlZvaQinoz1nkJqT/O882Q4ogrzTVprz2FNvdZUD84aupptMBB4YNEvU3cp1HtO4
DYDoQ7m/cQIs+S8ZhwTRL4FbMdIH7f6rvrJ7MXwa8YdUUhhDf2Z9sYm+gskNRyzdAx/XPF0hksOp
tLGdIf8DPGAIIgc7T2S14gxm9hT2CVUGNqXrFdT9HgR2aVBaF+SNtI2jA5XwFGl1p3Yp+O9wcrLg
8T3slBeWivnZyzdq+6dmS7LR2x1K0TdCxJEl94RAa6hCqD8JdNa/zq+DJH9DWyewq8Pj7NyVL9Xe
WDJ5ZYddkVFX9nq4qlShdbh2rhuQSRV+uPDv1vY4yC0qikC2qrGiBgj+oWXyYC1/joi7Z52hs/am
zmHBLAW/Fx4z7jZtR+fZniu4BBaiEJbkqNqUuMnm1qIj0rEHwSLAqnbE14ufdsDt1QXVwolrHZHU
gSD4P3xVMe679G+GQkdTDSVhognk2Eub+cSPtNpSawTtEK6Bzxz8358J7BjX4auBvPqVYVIUV8W1
ApgrYY00J4iOhP3RWRT+YqY856bmy1TGZqVQaGQZqQIk5+31SnLIVgXDk8H2b++9a9g7BJXNNccz
3oSnUsmXeqQ/wEGrqla8ZSWSpPeZH960YBU7M2ahU4nUrZzeIbdGn91AdQeVUMWUelAYdXe7M9Uw
1T+2H2DaKVicOaxLpiWRl2Qt56Rn7l+dMXURAnQPm6zrIJVlEzTK7U8RgvZ0fP+yGjqqiqD4QYIB
yegBddXcsJCngw2zrr/4OC/GeAeo1OALCul4z+wJwMC7Ewg3g+dJp4MKFZzZbedrfESzZ69m/tOS
kcMHGhLmrjCMiMM45Lk4VPIGKQX2d96zz53XqVJfSjK9fqQ34X9ChTFDNGmo3J54GQAj0yeANoVz
s/VR60yo+OESNKhnWIAdWNCHrpTuU3TmkWlsmfzAHKk2dsKBShfupejbFUIfqHJFLCXmzZ0MkhRL
HS5TVTBiKftQdivdr6LBnHLVA+8+jyb3ei/7zXFZvFUUpR2FjaqBt4GHmAzlZKgPDMPGNDgUxgSp
OGbuRE5Cjxf0XiSHKklDfR98hR9t53IxC9JPzVrrVBT/h6E4gEyk9cskkn3lp+n3pChEvL5TGQ4/
xRrJm704bAi2r18Is9s1ph0ua7jqxlu8qduXKpw2P1u4aRrSg5qdS9ezcL3MeMwdfOpXmAOUd5Sb
GrlA8qCCaxnaId7YETyd3+qs38gTbw+cGBEzc6VbWl7OJUhMae0m3b7/V5C6/K9zF+napOnii3WO
6hjk03Njm7LOqKEkX135mrroV44BCQUDDGRdWG05SATLMUBZ7odO2X7GRU6S1JHM+b7M3ehmKys0
eoQWTyWtHTKmni7lDhoy+75A8WkQK5sNKkTJSW8sGNvWxJ8SM7mdd71riLuIPqTqBOEby9Sw+iH8
c3jxPJdp0SQxQW6j6vY7lQIEh3Ff/EeNLTDiVOw2YK8wf2T7ZDl5Nk9bX08KH8RrjFmxbyQeWZmL
q6GwZ8tku/6bhUpVLxjVdOuPtdOkor2dxCgcxZbMGRMkSn41tGFZCNgJSPw3Lly5LU5msNIvXjkL
dQszL6gh27o9hK9qdzsmT3AATYUc3mZKJyc2sWQfK4c2wb09IvG7OSvVBpQduSw06HCX1GscWlNR
yx5YiifCOH2GOTezIS/0Nr6IAGPkRM7JAPXkaGSvc0yVqnOmafmJ4CLWwGN6v9wXQP4gCWTHwjyY
h7GjltU7/ycbbXt5yZHTSw9/0WxLC4ze7d7pXL4bsRBwd3V9AF+H9IudjXmFsD3fiiHUuIDMnkWN
i4/vGvhX5kT2Ls0Dapck+i/RWDEYWsUMomDgvOkQXmBM1mabHrymAU7bKW8rgUvClG+tiP+/Snxx
v9CXuZed0L9hozSmzu0KiTSLHheShzYY3IpCJO5yk5/XCkKLmlm5dtSeQa3GCQndt5Et71nO7+7t
UteqWHpRKPWMdcRdXFw46OjPMENuN4+JfN5j/U20sbprbbT3mlUFeTa0LZ4YrWURQqsF8yAxIbOg
Lb76t8JpEOKHLxEEStCw0N8LGk55owj4tCG+N92pyNz9tGYyIYt92XAxFfOA/OPAv9kf6RQbCdjj
YF+LNPA8Dlr+rEGKG1rzPUpBzQ276VHElP7Pz2Pip0k+pWxjexCl9UBLbzbZ5WlKyjKs2IkdRkqv
bvuE/+SiVir+DpfJD6HMuH4wfaDhYCcQXqgRrGB0yhK0cwcRog6bQLZmPDW5pn83++XqN3qxxYyX
jbECcijO4/3NII9m1vOSWwEGaPXgBXzKtvOFHPESYFXIVTK7kNKhDj/3qc/wCkdivbb1A+rTlwel
U68FyWWhxp//DZpk1jV+2Th5uHTM447TEi5lC2c+K1n8QMW5BCaLp8u1b7EXjxwhJlM3iZkIMmL0
uC4+9Fm4xGJl5eL3JyJTpp4CB3NQFmVTKYgNPWJM/dH5VCzxBNmcHkUXgYQNpOC2mTi1sLB1zBdO
Q0KRctts2P6Co7jqXKwap0yerEbCdziXGb1iF8EWKan0E5bOXlyLfKj6HbOceHH76eWWiGZOHu7L
UjXWs3yMePMr8H1z7Z0eDBQnD9FT9NxpwLIyRHIMdorAbgQWNp9LLMMMy6Ra0ixd+58J0qHrC1d6
IziUOtQ8i5SaMpQ7LMHgmagcqVxn4rE25frscSf2/iTE/4GEz6DeuNshXkEnSLPje339PtbwXJ6y
uw9UiJZ4DQth0uJpDy/dUzL+p+PzaZ68bwmxvI9NBBXfOsHz75GTNaGNLqxgAGYmB6uTb+52XTHA
gLQcwuSXoA2KDbKvbe8kzWcnMrzmtgBYj7hQcUu0fjnsdG6c0ZNuCyjHn+fUSo17jS09goLJOm2J
1cPmdJZHQoucjRmgKv1FAVAetNbMZ1IGi5IE2cedJqm3pENermww1qkV8cFzrb/F91ky57/hk5LJ
pcRlf/hQFNPLDdsCD+bgmFa5bweQMzH361BOLLfvYvgLVmBPMaNbWb+3e+k5b7tQdVi8kGPdSIfB
DGnIKxkAPpucApnBsP6CLNuL3ft4tmdA0Z0FX7qZWI+aXH0uYjpV1KWQ59rF/9lgSmHN6PBCa1u2
tr/2wdeEDNe9pt6Yl19jiJNnl/edJsO1Hq+mzTAB4n6RBT13ztFX4SL7kv2n58KNUvuBU+NuOryk
udkxg7aiCtwTZgwxw4p0xsDhKes6zMdJFKRX3I1Ruan1nAR0U4qw4O7dkTw4SWXYNH1zNmGiK6Vj
xHdFZxlr9lDSQC8wEREPQYaoZaigbJmIo4OghrSOuWdxwSSL8Ivb+UPLYR5/Q2NCINMo69Faww/1
mX3dJt/fsEOsIcK7dRUI4cKgpk/X7vMoR9xVHrYjh2JAONcqv/rSSRzyBkQOhy6BBmvsj/NDl1ed
tUJSxRc4TkiKpHsTqx75nZj0LgGZ7rnvITO7fivcGglv7CQcpx94ceqMjDCRCdrqe8RrmmM1kKtZ
XlwQRwX51J3PlzK2OLBnj6q6LV2L7epOEttLVrzt+dtrYlbhJFI1JsRxhXFox89G5uEJHoNGGjYR
nylgfyJML5M559lMCsQfBCv7vExxyO/TXJu1Rp1NMzCke+XOLtEFm26+l8XLh6QHIn0EpO/Lq0CQ
O7rfvtOuhDJIqEKkCcgrtyryzzzydlm4qgq3sPf56kIORMaFVJE4u9/dQQQ1S5zH6rQTwiei+l0d
OPo/qJD0J0OQDxiVmkMVCdQ4tTNTnumqXQMsbT607MXKSpEm0Wcu+3dp3JT4ypSrcZVHtWEmEnGM
Ie7W0EyUuNt6Gwrb8Z56u5dj/S2CZDEWIBkehUWlgWgreNzp0em9wVhut8X7UXkiucvg/qkaICSo
KlPet8hUzXHIZ1NctZtWL7KCxmG9j++DCrxVGgY6FgPeH4+qciTqN79vMXusr9OX3VIgAt59+foV
Jri+1GZvkmt3itv9TqrKpuaoc2RfjGVzSLOVAEC1JdkEx9DrPJd74OV/qISOJOA+6ALIacvE64l7
AmL7TbpMdaZj0pGdMXP4qB3shROWJz5G20yKJQgmoQDkoqUgBeflVFwz0lRLqXCxxfHfOqHI86tU
6mr7QvaMSXwpGeTa8uOdKPW0Fjb5ZDfOZyS1vpM/izSTMeqAN0jbLDpc5mzxQ4Xp4YEfKX5uSCin
wI7iWnkXMTxeHeDMEYWGX/9WlntQE830J+J6ue+Kz9KMDUTziQpDdrTJ6QJEs7yIcRcb2+fpRjcu
4d+NS/15oH9eNE2H4rIJD9aGLfKaFJYcHUkA7eVjfOZ603qhuKzBfBZVY48SbZ9J/AXoOyEoDfxR
F/Ps/fFAc09jeI2Ocb8vzYEnas2SzKOSvT88ZxvKyhVvLA7taV9CnR14LfAe9hWtx/G6yiEE/ux2
uiWkL5d3tH2uJ+EOpNEPqniDJagfTfx5LQfBIAXTdUnfuUO55Yd9Hv1CWh+N3wJZqbokAk38RMWE
BqqhHqp8Mtb4obdGJx8qs38bFyqSYpZisxCR7ct+Ai8qQ0JiC/pvcfA3EQc6qik1F9hcbF0tuVLp
3A/B5l5gAxP6L15IBV9/PCi/De9UCV5guKa47LTPjo5vSyv3aJT4UcFJgAE1z6hR1ZdtKzo2OCVm
7ous5R7jxopZ7D6H26HKDgbYbnCKxup52vuk8dElQLoRnOVenbXuwKjNdN9ilfZgwfZV8d7zLXxg
6XnOzsWr91DdCvV0qHMt4fX+i97trOHBaKPiwWADSsdmm1aBDg7ErGYBRf0FNUAmjhTz5qFxZYVU
gE2jiBwEXOJuLpnO0mMGY2HiI9RaZ2p42K4ot2jo+KDTqvlULB4r11vfGW9LP2uP+mFUPZSh7Iwa
AohpgSm9FbXlnJleiTtuYpwZh+iazxwQRnHxRBSXOALPA99anb3VSPZ3KIKlZL//g+DX3XoyPieC
jQf3LsPqamkXPCvIko7ySb702dEHs0z4xF3cRUXRlQG8tZcJxt3sUz7puBur+XAWFcKQKcTNKOVX
ukIbgsNOoP3DQILBSWihknLMhcLD1Y+X8o5Pb+hFFBMTEStIxhLhJkseNlTXC9Bwq1uk0iAxgSMr
18p+k1FAd7iZqq0bSkkPPu/TkH7CgNUa0B8RRt5l63njCzkkoboJSd4zizkHe3IVlngi251ptH6W
9GwmZftEEhf/EaP8xmgz6tSiKAmUI39eaG6EWYkXIczj5wR5ovQ5cX1sFdoQdNIZcVj8u1+rklhA
8l0H9IuozfYKJWZGq2k4/rPbd45YjSHKhcfN5jrE7ZyE4ElRVq523XLpU/Xp+gaBnXop3pSjeO9+
bJ334XX0cxxreWmXYvLvLaU6uuyzMTRez2y75idiovYZx33AW9QI/++bisrMTTwSo01v1PSDLVhy
Jn9zdtJdOIVReQRBJbH5MvPs/KtBKUWQNjn55xsyNwT/tQ5RvIWBPgaSEmnkfSxe0RblBRkMGhqW
Jbd0VtmhYeg38keqWAVOZWErtXR92qfhNdLcBhE0+zwmfVjGSkf/UMaI7A7S1U1Hwy84S9sLBk8c
JUwahjATU2TyvZqP0T/6zvcoFhIDPoOnCR3GDmadVeTths5d0wi8BIFlmqMMpru5yYm0peMB8HgV
kFM4luhBb2/kODmcR4MoTsRDV4jKfIUbESw2awkhl6suljru57U2yvx75NnlxV4LsRMjtTW6Ycun
tXCWaCBHW4VJ9zg4kk5FhTwhU3+y6RcZE75ljKngEJOJ2z8mwrPfLOGVfVEdyGTvoet4jxl51zSx
XHaIiaMJb7yEYHqyr5Hb4r+MzLckgZUAUVELxUR09r2W/SCw60SKHPyXpTDYOyZ0UkqJA4Fy/6yd
KeIutkBG8BUMmMSBYHfzv/Rs+ReYacOyxoBHrYLX0Xu776jsd583EpQsCIcibUGcYsiU8O4AXiQZ
bAiUG9P1S4+3+Kd/4oI9bueDa3KhhYVkc4pjNRcK1ybyrx7aAcmVZR4Z4RC6pWH0COAvkcTugujY
MH0Fa1n1+W9OOJNTAxAXAlbsa+Q66ITlWHejTJJMVG9sFQCVZer9FoSBq7HdYWuNQ9sTGbfp7PGz
niXVktTOPB/yz/7GmgfRCgBbimjJqKst9QDP1AZ1Ph9iJA0PANn3wdhNnPqYkKfbrd9aUBA5i5Ee
My7cn9TE4lW2OCEXbh7Hl49Z9SrIYdPJlSaH3YSjBdHTeWqyCO+QhCc7v12uOoj4EFoQ3uv6CTIM
iAaSTE8U0eoCPY9vPVnlll3kAsiRAesFZgB+I5dH7OByQXoIE259pgkog8sVhPObdhg8/4iFUhbK
8QF2nrmpjLhhS2OVNrG34tFBdj6u3l9JxbaSCDDLHSB5BLhwGOxZU/4/CEG4uT2MogVKwDydWUhE
zs1reqblT79+4s2U/rOFSoE47h9LmSdVvXQtV+vXz1e8626k/kSJaaD6Tq/+2MTSf/WiUPjq3t4i
vzH0VK13yG4+MWqu99rFceiNN0rB65NuZIdf8cqRikVck0h4hmrwvgFKrUYarMFl8Q2RcWFFTYdJ
NeuDL8MmjM5Akq8T3jZzml+x1EuhfsDi53LEBUJy8rAE1Ouu3cHZ8IgIfBqrPFF5g5Lr60W9bY47
IHvFK1DuFwV8yFtfpGZ8OFrYNWdpJ6qq6XZB2p4RoN9pxRr45u2s/55ViChk1Dus/HmbTdr0wXk0
mzK5zoabSAbn9zCgIJnfpGVqy0Ke+sfotmBCwA7R2g+7ohm6nVBPcK3H3Rz+A5FW/xnElPFXrEy4
lt57GWZdp/I3xKz+Hl0ka8uYLP0L7VYUTxSH1BUfpsd93J6XS6fbtBFnIomA1i6YlaHqi29KqZn+
jb6YvUiKPiRStdVkaJgQMSYFKsW4byDYJwX6ejQui+aEJ33elnvB8fgp9PrrnA6Uo7ZzmDV5bvMu
wOQ+XT0IjbUor9zSV7oEZpUSz5iW41qwiKw6OlAplW253FxVv1Ushc6wfSUd3hRdXp1htl/PGEDz
x8vJ5HOb9aknCCv8nc8wm09ZGrXh+OPAE1xLBDNSZ+IJAKPN09ID2ivurFYsK73AfiMlupSDnXgP
if0QaeII3QJRZfozjou4Tr1NA3mk8bTAwK9u5TPWyf2HhqfCz50xTFTk0wL5eXKpPsZDQuxYPalY
mK1zVN3RuFQkJrYvy7d9BqLdj8aMRNo9/oLNNAAluwWGcMva8zn2BJDfMIsWd7F9q0ZIUCLmsCLN
rH4mmvWoXkcWU0YX8kpc1dgyFG1I3A1ZP9JnccZoiZDfxgcvh4Zxnm08iAkiAxIRiLKQGFZWiExB
rCKBsL73TdsEL8VuKCuIc1EZit6poFlBiOh4eE1CQNM0gE5mytD7FoIOa4OGaGYbdqFXBf1ZErf2
7cwIVEy9Ti2ghh6PNObG6ub96eBj1o6zJTTjLjxbSe5mkOGdSGYcQyb09Kw2hwuwKcDqhBhLsfRU
jegLkf9bnMpO968rTW/ooHrfpNRmHj0PCp/f8s5k2j+4MK+iebP6GFgU3pQCmYe2zP9cuEzvVe3A
EXl4S67vL5P51BgEw0QPg+Lxz7IbekxXIVg5iNdLrxbjYtRc+hGnYwpaqiqZXkKRdxQfo7xRkP5Y
mv/9JcI+b6dffZUhSUM49gzGNH+vaf5W4QJqudqx5TwAPJA1NFrxx9SKT4bpeXEFY+FhR2h6lNO0
XFBQoIQfuBlVuwwfc9vF/e5YglvQX4dPJFTIlOONpSZT138/HeXcjMrgBhW+QtsztzlsG4vDSbjC
RpRCJaiAmG5F+CKL4pR86HIsHySqt6J7qId02Bjp+zXUs2yb1lZzPZoDW6jpMF74DFF3bcYGJiRQ
XxtV+O6VIC0H4X1SQhtP5UDVfLj7S4LUv+mMz71sI/+U3TBaj4FIBuXkS9cg/WxBTo4ySl+6PXHo
/Pa73jb1T3RTlVD8YYZlo8l0AZLInd+W2MtPUjZhxGKnb2YkC9y6zjl6g7mg0Dk9CYYjCnSGYzHx
FLQHzD2i30Oxz5AVVEse80zoYYloxZWiH0k4gGPIw78P8yjwewRfVDmxuDRDeACWQ2f170t7Ukry
uN6mP3WcN2sLmJ3ycTUacMZchFKD95ZFRWe39hjESYCzX4DLyfWnp0oqol3QIv7fRmvt6Y3SPBqk
pvBPbXVKzAdCCqKDMG72iS/IaXiG8GhcByIdG0iTAb3oFjjBoJOnrI05aA0+CLdEi6kmZ9PB3/tg
qfyIBaRT4RtdvRjc77/whlF2JwmA46ZBtMKW9dnsBH2QdB/fliRqzq0BDjysnPVIFBbZfWGy7Lpy
dYWv/hTwptzf1q4kSiIdnyLTSDhHhkFYkRugs23+5N5HGk+PmmICbQglzmmx1arVL9iIa6B1m0gq
3Rv2DmY7WvA5v7oSbduBdO7DlgHSDTv03mX1TNhYelrLi+Nh3kcQuopfywkLZ6D11r7jNIZUN2Yw
TNrR1JzJDaQZnNSveoyoas764t7d5gS2sSO66+gtI+HGdu8BYhU3KPUJ4UXsB3a24PHnWi2/UFVm
kwnC9tzaIMWZu0pVLFzIDnM5jG27V99ye54Pgbbz2kMDveh4M6uFhrZXXWoKfQpzyL2pBScWYj22
Bau7+aq8HvIEW76hAAk/4ckmfgy5SYDRysRPT7DJP77+H9FByJAxRPy9yChF0OIsYYI0K1m3I4LD
3Ts+XdxqJTNE6abxZ9dx1fCl85HRnP66PKEV1d+Zw3oMBlKqVQ07nxaPXiKnLvsekzA3LN22Mwtc
lU1KIXdYyXKaRfMepFKd6mZg0EqhKsM4yOXXikZixDA10GKMInUzzayN6hFglVLq6B6duIcWOhhs
nWEq/WNwlBnOz8qN4m4WnTMoqxfq/278KLPDtP/CrDCUqVJUspALUrpcv7IqB/vdObGenRIbK8AN
DXEjen2E0FH9qqbhpciovA70np96cIcur/taBYrxMylUA+RjJzdFLroB0CVjPcbekpWNCs4VHLkI
s7e3tJntj0oOKjKME2kky8m+/jr6wkshU9u15emm2aGdBbD1Ey4jC0ek+3tZuWqSE9YNMsB2/kpm
jcn+jQBQKmzfGq1pIoc2BcEdnIRZTZXZffKDD+JDeazVqgrzV4wWwwBX8d4iEWodFpF9fqcOfxDJ
wUxnYKFBneoTu8fg1lvnIDodJQM4PyxPW3ezCsgqrCFZuCDnTGUC9RHMeoK2RqyZ1egu3FPFcWes
5E0/jzuFdLGuq/vigIWqJvqSgNgVPNIDmRJt/f7Qhbg4HxhOgHoU/rOqMBtbxJQNvFQKldG8B/Hf
OitETRDZCo/Mudei3p6V+ibhqIdjPFkLIy8kJjabOj27Na/IbtkI54L9BSGdc2ewyr7G3O8eMc9k
vuT0L+Q78GzvJjXjSIn3u36S8YqfLfYXgo//vtVZjlTXzzMy8q3AL3L3b4EmbDFa+vPrItMF8HPF
I31/szHBmt/fXuicCsivOUO29N63/EeVDl4YgBGrr8978vsNIMJZI6wHtPm8KKsQQTk0P1S91o51
AAr/gcvFpfLSDP0O+/Lp8aKK0dZBa8oKou0zW4HVwPH5w8+5HQXmijpTsZ43u7a4/ZF/MY17gxRv
SlqbUxqpMzKHenyL2ckXfR95KcNbD4tI43gfPFs4YAsJhfGORi1NFeneZc1FpdUGLrwh/zbfuOAY
REb94t3tIMPIn+M92RjoNfAFi9qymAKWhmycL4gqWxtW2vZcf9L1XjjlcmxlOHAbSrFOSd0tvz1/
IP3MXoUaQLauibe5PgeGGtQf1IVaPlUVfz6uAmJ/8wmmNyc/oQq8dCHToeNULL2pQBFoOTccALlk
uqFvNsGFtlGP8lDUdjqFHu1eJb+ABU20hI6zPLqKH8k+9uiQRqN9HP/Mz2vOwGvv857rrUKFTJEQ
k+1vIro5kkeAwBFmI7w5D3gtIEKWEP18x4nc70J7wWe6M/bInV9ZTdVmTyNCG/y4CO4EjQTm8HY4
m+8vxADwkx9bcZ6qI8ZknKawFroaQqs9wE5p9FIKlcpbit/vHEFMoGKy5hvh8u1N8xkfBAAtdD5j
moQ9btkluBI2Lc8c9E14rSjgsk+ro0v7EAJnNvh8kRpHh9sdBxANglYSOIN5XOfw5FtuhhwdJvtH
VeVip15M5HF9SwrIbXK2RjJnMLOCivQD4SWO4c+syfnSVVOFJPo7rD+FBTugT+J/IqtvAMysLXFb
jxGMqyhR2dSEusvCpHEYYWkRtH8a1nx/uMYciap/usukdbYLNOyeTJybh6KkvLmFaaQJPHFn3KJ2
O1+ZCL+5ScnCXmRn/MTUbVGPni7+1N0Fik+am9+/oDu2IB5QPENWsY+IZTQ5ZvjtZD720xkD9jYX
qzLVXNNkdYERyUlV6mgiZZ+JY/igK3iXPy8heFNXiP3jLLpKj7bvHF1bpVV0vQPf7a54DGoD7fLK
mJbN7/jDrXNQYtfbsTyFqBrYLVntMa3ukVXOKO/dVwYO0LElyQ7VHCmnHXTeZ7qCGD+6Pk28vNw5
tm029HeY9xxQHjlZO79jpnAglakCjVqTa2wWEzGlkRbrbBBnDVqZnnaegmxLVzmgBJQMhRKIRqsF
Kq0XJ57jPg+fjNtD+2jnoJIPpkzO8QowI2dMVlIWlkex4Es10hW86oEwDKEARLknJKsybzgwTCsc
7UbHSQPY4pDgbXH7r8CmTXZIKeezhyuTGI+wiCcMmjpyCaNbaBRAVA4+GwB7aW5HQe242MjSaarZ
IuLjYCvbqRUSiG4hLdjSGURzR60IwdwRQoTXDWPNtDS7gsOkVkrGEXufeqIWe9ea0heiNxUjnO72
T4hi0Xz+5EdSWvxBxHow+tTRZgJFOWIuK1oVZzYo+oDHJY8qsX0cBU1FZw2wNZx3EOcBYvJeJiXK
U4VQ20ZSluZQMZxiCf6KWB1mKE5mvzzUTAjANFbuGR6mkEhmk55PoWs97TefxKf66NTE1GDssSRY
tM3usUA+UkFT+ORUMzD0nyZ6FPnS617VBk7LNJpCNZAha0zr7k1xNkjmJGooCCKBOJ2BVxzKqYQs
2DcCik1kBagRXIHS4wfH8eBspf5X1KQVvDm76lURMPvZUPk74fVQ6Gg6PEpcXlFX+zFuo3wr9Oss
0FghCKMZDm8XR+ckqazO4bUbVz9OCvVxtmW9mt8zS+BKyk3WODaeYycQIhAuTuScoGKpt1H2QoMR
x9f1p2UBa2CwYd+DBeXqWNIwMe/8Rzx5bqA0OZLCbtF6uanh2Bx+cxkV5cSr8Ru3iRdzPIC5cFt/
oTvDGP6Ts9RvKny7Sr127nfu0SBduUdK2N9+cKLBDRUFjiAIGdoyxeesbPMTq7MV2HR6tRGMSYFK
ld/5Crnw67uuvpAUzt0rzs6XLLzqHCj9cYY2P52MSvZjOKAmOzos40FlIZ8bfwO8nbbrlcp6etdI
plp68QLHlDGlWAZR3HOuTPA2xLzez8lSKPVMzW8JfWYmW/I9ovZIK9gvCoXIsdrrRC1FIEbLR3cq
5Vi4mqv0BprTsLJjSk4g2LBW2J12/zczlvmh0KOphIS5A7v4C6alZZgILVD659/Fs2qPwKG1r6Yl
CEGcVimTpJSVrG7kYE64vDDMpUxj1yuP+S3+0uKQxR5Zd+YAAofukMHzMk5iJjbniPU1cAUxaF6t
47+qxb4mtwgfhVIXtURp5LIDsiTEaPVgrlrKLzg7UwpkcUB31VQ1Y6+ULxaEdB10NiWvhH4sgj2x
/OBQQ83g7Vni9C7YYyoaanZODT6Tx4aNNc0Sq9DuwBPJ3bGDPqZ0+pnR+cy9vWw7JsNBiwYJBdlw
lCd8SFp6ivb2CNsbJWnOHXbDN4ZMfOyZC84Njf3+ztOZ7hdds+JeCbKCl9nqj3S38YSJ92gIFPy+
Tz7DKjnIn32wufmd49uVI48D38R3ei4YoAiYCXa/+lsr1gJyNaY8RDp5cjXC32shiR57vhOXgprb
pBAoPfSVlLKLjDmfC3fKgQg3qpDICZfj/EoVnmOIXOvpBpd51CT5xdpTI59KAxIdIsL7ljC7VeUZ
Sfimuc/9/QAlnyAMDTbF0JNuZTBLUVQrRAZwxHiJhXEdl/SQ35tlxxxb+G8pQd0xXHZuJ5CYHOfy
SAG/HyOVLWE0Bu2Y9heVzZZPwVtvFPPAZXiS+0NsImIFRRVFBLRfDDNCpTpL9N3MaD4x7cXYWPKJ
YnWeukkgA5TM+drMUvhOzGHFmch583wWcBtItnhO5ry39E4OxcTlNaDEDobb5iBWgAxHl0932ZND
licymNvN1nuG4a2YyhOFeBH3reKtEaVhwVo1XP+WOMYhL6g85Fw3fST1J2nLerlAE/QMOFhDK3jK
mQqKnbAcnZDPEGxm5EOicoVFZH5YzH4NULS9VHS4e82HTVNhf0i9Yxbzeg01YvYTW7WC4Z/vW2XY
hf/QAAzRAw1Y2R6rQF62hJ54t1TjaLZ71lGjnDQePnszywdz42qevnGTSdmqXii/WeGHCUxS4xLv
WXrQGGdcxu/N+DbCKp/hFh+94367JsRB1v+iKTt8c1263y3P/VvZZt6yxmOEydmhd3200j/krUR2
ZO6C9/lQTpVnYnSCDAbMlxUs323NRk99bIMhDrXE6QwY58oh2kqieEE15MSrHixJplUva9nMSRQI
AkBoYTk4Wpr6+fwHDCs0p4kPAFdFtIrr/9qcocUJf9O1WdUG7MsMbR865eaZYabWEVjZHSDNL8D+
1pUDAamtsh734A4SEy4DpPhRFTWeerY0xaPwHcTC9aed7rpHOg6U5cKnXn/IqRZWiBDZCUczp4Va
MGpQQTw0NIZpwsfOXPgEtBlSogNoe9jvjDP9xDd/vyDpOjy3+WGkKgjXfd5s8lY53NsKnzJXcuZY
8rUXVpj9ySJJSB3A1aTqe4H+/FI9ech0wLFqBbZZsE0tdn1QkDi5d8GKdAx1rmaL11XQkBz4Prtp
VR3zMkIdFpf5bPwJkbYCdi1ypz/lqNpFnPPWH3/qZfcR1agcB5+pVOFPYqyiHz4iD81o5gr5tLyo
0R7R960rSZHt6DsL8CLCHF0ukh+0t++CpL6pZ9N+LkiZX+hzhMltIY29DLeI3M8wSZPmactsI7A0
THZh39XQhZrUKWo/RCuQqdU5W1eKGHkytYC69F6Msu3ROgMonMY1qFkuXKqZnZvkzio+dhRMDBAe
aX9yvs4+dQ49WoUUtLPrkvFSfz0kcYRSDKv+nwcRz/k03Wsu2+l/56KS5ZFlVB7sGmiSNc0hBnEX
Lz5EDD/cqR7OkyRPDKyr88Jh5u56IQQG00J1SOuEALbz73YaCgru1JYDaGh8cy0BWE+mR9Q4xyQj
KMWSMV+xJZtRbYwZXyCWoFixMpAknxW61QOmTQU8rIduZdiG7Dc1cwcnLOMmely4H1SRbpspmgYQ
S14eZqjsrnTQvvnhhS2gB+7CcgrJzYm9Xz4lNcyASyaO4PBdzG2aZPuy1Ju3aUxIN3tw41svI2jR
PeOuf/RJAuAZeqYGcG/S9yAhrIeXxVVPkY04ORRWaX/rz5+oWLWecKbVUEPo++h9V8AO8k1eyrnT
abOoqNDfInzpVq8q+tAQR2LTSt71Y8AFMDQOOcNmF5K3eyQwk0pD5es3F5YVrrfiFmwfEnjuAUUx
BmpdjhGgwnDYNP9/VGlMW2mPum3FC2FXg218FelOFwIjah2kMpBovsIgcO8N6w5mwXfIWrL2Toxb
DbOzaB1Mo/84hWTKQY7mVlZbUTFM7DIwEs7WZJvk3bgeHfAHroFcD2cShLNdafEy5+p+mI4rNHzR
11UOCNO/nTyJQE4GNg44RofdGNoo1lecY4CMkSOKTIx5w8oMBnkYHbLP8vMZth9GfI5XYMiWGUxb
1+g7DH8RebDFq3X0LtPjtsOc1g2QYJqeessm4rhsTQ6hg1o9Tq2PYO5BlNeuUbiFzjau0pvxEno1
sEGODcaMz7zRjRYC4gGnhrHcwA6oqslpEDLCrNUAQvMIdw1vX6XQZFz6p7cF9Fea88jWsTnv0Inu
CZClQFLNpFmhJ+61oaIHrAT9VPm0QAjpsONsHWGHkLUOkJkU6Sz0mTttU1iz3BD67BzMk+CJS9tQ
mlMWdK7/7ie0wbPQgqNpKSr2Hsk6Cwj+nDvKdfJKd1ezgGgEsFnwLrmVoAGWs0bwuyN5b6NwBqfT
C55wcxUvKIP24L3YGnIDPN8dHRHRl4rCKV6ZcVw/e9ne6goR2FIbOLqtFbZxLSRO/6JWCxO95Zk3
GFTViPjdvwpstpwRdMqVy6pdMou6CoCb5xqvh6L9+r7jqlwSRs2ITL9RSFKHsvGnngsR39LuEb0N
LHEgx591MniPcApB4OJG7cLYxAYUZekniv9b5Kiky9yam4RRLpZG0SjIO4kt91CsKZ4FpYjqspPD
cuci38IDbCiGCpQdYdY7MLOaPifetTxIlaslfqB+U/SWGfbZIpcCpOfFWEqQn+TDp0NPg4tnpm62
tEhxITIBDFwbMkdfAWN8WLTn3b7WWgvVhAHTOZ5AszhocsAxnGMqH2yGtX6kVZ+TO8OytPULwcvc
pHCqvhMNM88BPVWNZHw3jwwkbab4aGNfPtZSMiMX0+/2SIECBleLCB/bfaM3NFV/htUjo7VQbdFU
0a4KLOXhTT1189qSigPHT7X1VwCZEbp6syl+v3GsZ1NJMMnt6xjN7MDSFAsgdUHcun97he5LGVNJ
lHQ4FJFoNhXWvnf4mP0Tmqid40EcB/8Ag+MhPMTuIHFebSM3DSOVswGeubRfd4+oelM8crR3W/HV
AnDw0xW6veTmytnmpSmfs5rDMbU5TuMlsUY3LgddsR9Tq/1JLqtv00mT7dsQFBH6b67NQ1b0ndoT
CHoISLMlO57/Tz9agVgkfx4ajkf6CQm3xx8eqNEK2jEbcXvg8VwnNGvCmVP0YpZJBZExLBeHkGPr
F6RZ0uVJywhk/iELfvpI20S8nGqs/4V226XC3KG37Yj3LBTtEBtNrgj4quG6wqYo4ordgPsmd+3z
rbvBi/29Y5x65YbSHKFqCMbNk/l6+pupRW3IIaiQT5j37p8bYCrkY0iQAOU6SQ6aJ6Vqhvdyw81S
3jDDRoDhZA0ALiKjXPxcn4twFia2hDJeW3pzMb9S3+wUdZRHRj2VGd75oHUxKAC1rrR9KtmIy/lZ
4nyhm8BZnU43JufclJiy2SsFu7KZj4rjhNO7a9HWWRo32YkKVge1oX9H+Do+k/iJffu5C2dyKN14
+oxutmBRD6lRRQzBlkl/MZDe/wRhig4bBdvunlX8wvd2jVw2SmPkBG9HNVNNH+eHR6GHJI+t9YV6
+h6ePMUxcB4nhjzIZAdgJ2kzLN7U5wXfc2XJPxBOYBcAAqtju8YZti9jFFjdxn4LRYBG5UpAfIbR
noHhMuQCikvcYQ0No7WzbKINlQu1NuvTzm7CUj6lsNnan+caVWxsdg4o/MIqJAep86myCpgmFGs9
0cU8mx90yxQckFNEzpZ9QIF0oHM7bJujwZGQgE5Dh16IUAW+W/HuWTLb0R/7WEfkhgs3ZHQdIKau
4VXY6W0DRDIFNSz613tlgiB9DMd4AnfPZt7YiZpGwzl6YPB3ybEtRVuetC1gU9RTdbzj/e6dRzCh
PHfOqHGuFuD43V7AoYTfPPunas/umHe44QIj5mKuuy3O2SbKGB6xtDmY0s1TgjEGT0RGiLINALmi
tCD2V+A0lv3trjVzbAyrELJUlCVxN2TD4iQ5TaYMPEyJzKgb/VwMf2AMplTTxNn2rqVBwNuQqPqp
EbJnU/K4iMV2mAGPwia4xThI9Oh6svHxl+Kxw/CdNXaNFh4qcllJjN9qwnylg/lP2BvSwJdPAOxf
dkiVGknj55nGIOVoH07GuqKUfQBvH0F7HbOAB6IrISuV8bHOpb9OC0vugpMB/+23deNM9vCz8TOw
0oL4fQVoTBDsV4zjqrup1uJi/wXrJcSAChriZGOjhGxh1mPjcdVfM0eLOw7wQN6KMUy8VBA7wT0X
y57XexhT6tPRnxDlY+8XeaEhq9Crd9DmIjcsZ8bB2PxjsondUAQYKfMBuxQ0AhOBwxRK/620zP7L
KrT0CluBy6jqlD14JiZjLNVvQ2yW5+bLQLctH9JCe2LMg8EzovCIuesPAbZUYp7bbjgWk6JGQUPR
k3GX0pe6AL5mkRJYipLSGQylpvmj32AOfkjGMqqOzbAy2kWslW0PaR+s5NO2C3o/aOWRY3O0YAlC
z5AyjV2Ko5vMFE298XRecAvRFd1Y1oS4P6DzyY7QDIL5dORrgPup45TdtWFm/nPtHHpAUHVRxKVb
NGhUbcpS1xmgq29t3pc7N+cQqMxlmL8QV+zXCWykFTBiVME+PozyNppDbXcoTIuz6Z1qPvDAA1j4
SbSdjTeNGwnzautR4yZKIFaG/IQHkQoiaUBxCfDkBPN3xU03+bEODYxRAB8oYL71ybs50/i88pYf
OkeFHA0Ack7bBtEUUBQL/8Lc9VSrLGHIZEiTQhwLSYHJGbN/BbtyTBh5yn2p/gsBwOzEPSvrUH1N
chcgpkY540aShxQandTtZQJbhxEJiOgVgSO2L3CyoluFVuolDwdV9KyABO2y07hTgc+18zEibnbz
6d2XaMegWeeR/lu4gXWAAbeaFkh5h0xyWNTK/qsN/de5v9UU2J21xEZIOBm5fGTgJDO2MW9z8YBF
spqLEd/QEktU58iLNAGuOVM2fnngD0kMiK9+eResT5UW04cB6LaLV/OX1NshwyjAk/rBeB1M9KRw
kZ3ZWjBxiNxZ4HMuZA/YwyN7RCiV8gEP7111eFXapZkr4WkEDSIuSK2Ya9HDAtTMlNm74EJno/h3
rcRs0mFLd6TiUGIVPtqffOYcePH/rB3zSCbTtiQasPEphwtcLJPC2Ng/woA14zvhjgkKdwFVigpH
+a8Y9WGwoC3vEd0eMOqS+t8hzPP8wCU0zW698YiK0dK/qAThKb7cO9/DJ1as2yjvYxDRRFIT/0XY
SmtXVky+0mZBySSS47eRBwtOCqvl3nVOsuLMQmxiqucbz3DhPR++GJtgGMvkgAaP5+xliZR2Fj4z
EARV4BnjZPZLQF+SZs7HK+mm707/rd7appGzD9F3sbbpL/P4Wy8XgUcHYw7FaamnujsXu2VDIXKk
meqIkN6eAibPEumYQ1Ivcu7m7arJffz+fSHspPdkqhyrGI7w/ZQbpDOUJrWXJt+YWupoY00KS8Fz
jPvB1CYZP7mVuTTO9wAsu6OaJ/cnB0zUgebcegvwUr6N2TpT1h7OPbTjtDdRiUYWxx7x0QFB41yq
Z15T5aTUobt/tcGTX+M9uX6FwVLr8+o+WgQi2qFotM37nxQYrIcj/gW4BmlZyWByEHZ4JDN+6/ST
MUWllOcKgxQuIB8cadhFcxKFCxd2fBlA77yDAi2e3DybsV8tvNYa9qcAZfWqgM1XHc4ilKLryvER
dlbGUxtgbuJ7af2Bk4JmJOpsk7IHqGYkjBnpKVp7/hcfFbBr5zzgKksPiEXrdigJZT6HcKxpucDd
86XvzIvxQ6EBGf/bd3ec+BXP4yY20HX0hMUdE7kI4LQPPFBfx1QAOgSYQSp5bRjG0fb8jwxbSdGi
eQwu0uDH1bh/RDzT6P2ivKtJrBMegIUVWzTgMe/JQFHu19xMJL30fpCnewD9/yd0m5sx8a5aanMw
nRo7/7aYsmnJvLvfjKxM16xAu3q8l+GshosM/Fm6QFWfLtLaxFfYoUFujLjPciqy2wxsYIlm0qwZ
lhHqmnHIoy/PXSjhM5MqTPqHvRNXFHfPm4De6pOFQ1xNyaUMCYmIgzNXs0JzRMnaCpUI8VkPEIG/
VRaatDtPM7rj41LOz23/XQa47bMo4G9YC131k2zvFVm3+fESvKGvvFwqoPC03v4O4w2CwPHDExG2
exfyUHs9j0t4rNfpBVkOGtI/fmdeFVKLQ/2uY8J7X7rnRLgjzCTesbKPIRlZkSxgrVEJUtHnWbGA
KUtHMYpHPWjUxy9yc/Vb+t4U3t09oi56QJSEDFwuPX0w5uqPtIBJd8MppEAgxvl6XY2GR6Srrv2I
S+QMmPNFjMXhM6BCj7OWiNkPUjkzdYZ3rwJUJTx2QJHQOClGUsc9yi2g14s+WkZQSCSbbiKBKvC2
5+vCe32XzArj1MWZTYwv1eU1/nTSsISpvmhUgWfswzQ7QNDbRo8xFd/bdByZufVMhn20J/zJwBzs
Q/vwrDDaUCUxe8GWSbIQ5VIp009OHYg6WGJ4e71o5nK16v16fXZfVdeZKujOeEFwpUzEc8e9zg/5
+/23bdF3mNYfbZBxWO1VKyOuV3zXkB4/KOzciQn2hqcmAT70mZgkpToKt7xbvvA1gLWioSHgPpsS
mUXbIAsfRd+T3urt0ARWS3hDA5PkUbrsR7CQuaF+ZhFET9Rqd6W/ECJcSHBF0g7h/pI22qexaTYX
UaCNiL6VRNv8SrvYjGGmHnCmmmkmvW3BbEqxg4fO4js1WdwRbIaq/sELuSV+lCDNS/R3c6a3W8C1
LCaPX56esiYEcg9auAy1X2XM6wvCk5hDEPaoLUKq/ipC23aqDMj44rqwc5nOtG3s8t4BeKMbIEu6
f0+sB8aFiIcs3aODjPP3R03AtIdzwc51IX4ryfecr/yFpTOzMOIaMK9b2BcpgEBSTlBHzCOnp9p9
EWi27g57VMaiIusOy9tXThqkbEfGuXtXAoPNJHokmJWa61+eQ73d6z7jSuCyjORkmxva5K4af/+b
SmV5/6wOrdfKHokpl5yWGshYVufpfr8dJbt0dHj8GmHrJ4onGo5kwDtb5/r+zNanrm3X4P1xrVMD
45fWyQio7sdXdGa5X84/+gnyaRFH61KpKtgUQoWMNJb6wZ3+kHi+nU+tbOS8T/BOwx2CaoTDR+3L
rFFRRdpyeTJBFnXLkelecdpCI+TqEAgzG+1uMM73dE/R+cnqNs/e1DDie4zL01zsCVUKYNbH3qe5
B8c0LJPv5H6Uw7Eqq2QcwuL+B37rmKEpmkte4tfashA/bzKTrnulbO3G0iB89eciQEkOBwH27tfr
4+QV0s1e6naRxtO2sbYLDdpGSTDNH9NbxEdh1zQNZ6YGKPG9ZgBSBeT55x305UDHd0TftSvLdRq7
KCyuxoY8wZt4z82wIQlgwRWvN0clMY38bzxLKrY6151yATMO/zRTDWXdCfbviE1yUhxxKWiHy8N+
Eh4uJ3WAC9CuAmRoi3vqBIaIdc8bVWoTXhsw+VtnD0/Bn21M8RKWDQJHU1OchXHcO+6k6CDdDtxg
mBqkN9VgZBTrxN+BW9pwdOLrg0mDpBrEWFodlNXwOMvTk9VcwJVhnX2IWcu90RNpvPJCC8aWRx+F
N4wd05+O9WMn7r5TiToU3j3bpKs6wQj5LvZKcuwAMYv/y8Vs+q+nAJqynnfHHbb2M90mjqONyh+A
NWpcie24PNmgqLiGxa05oeInlDmqZ974hEWWdR7nwiIVQcMfyMjozyJb7UYMGwVaZm/g+l3IIQer
4P24PHG23U5zQaDm6zaXyVlNC3NIwoAMtbLgqBkjNnMSyq16A77Kbut2MLOnPNTCLCrBlZ/4JlNS
z9Kgw3bn3GHrua/HusI/ZH+YIyBoMWRuuWkrCQgg0Irx2WMtRuytLBnHW1Ks6+GMP93JHrhc6oDx
42VOHUZDEqYeBPr4l/r3SbV2vkRCC4UxlFNYGyBxWQM6seJaeEW19cMS5MTeH+b2OeIrL1f1PxPJ
pl30pASKIjDCFZMSSDDY+kmVTfHAxO7w6deVR+NYsbsJDNbop2+8ks3fdPmIHpHH/IhCmG3Z1bNM
0YvOt5ReouZzQ1QwCLCwzH8v1JCqfXOXo8K6OWAgFapxNLcX23fq8XTQnhvnbYJXlGWjQ2sQtI6t
MVIwJC6/yZxxFHB/97dwhWxwrna17/h+7MMHTirGi6EojKsubgC8YzhuY5CHHCvtzPPzBO7TivHZ
ztBDzYmXOTKgu7VX8f5OXh+tQZwClf7+v/eFlC1iXpSjfEg2Fzx5Ud/7K+u+Q3feOeg5UzLhZ/fa
mMNolCP+IiqUkCwRwFQBKw5hwRetCnukpImm8k38Ui+EZ0Z7s1t+/4zrMUHI+dfFPA9o8dXb0bL6
TwTDENYTMesqCTe5UPYru71DXuBNtK9vvxq5DcWTON5kcu6AvfepWoIQFyzPZ3x0uVEJa5Ze00XM
ApFvNfnVqpe0KyT0ydkn51ig9eQk+YQxyK0ZMG1SfEEEYbaxYJqvbchJ4lrHYz93DQ3N/g6P1dPD
/ZcNJqW04hxIJmkKFlnKIIg/orz3V3OhoB4+ZT04nTkW7p1EL7rVSqbULrQgARATJBqWUgBbnxLb
JP/balGS5tnb880wqpv2cG1O2v6hSIbS2DRy+YGgWFePKI6HAgJsa3pHe4NAkNSSSI6KtgWwiOcv
5AnI+dotOyaqKfttqCWW6o3hzxaEMM+piJlY66GOs+Yt++iBl216IASPTyyUHgY2uL4RjF+t8VRW
6/t6TDJXYTOwp511oEtTLNoLan10bU4rme1HqLwgg4q5S45n+2/uTamsHK90k/Bt/DtzDGuIKqo/
kVRLvaTuUbQo4IpJrKRm4gdFGNc5rtUcVb7d00ebF2aU8Aj7gss3yX4CKx5OEVj9X9lMaCtQHAAX
q2NV3FpWGGt0fBVKqMgKWW03uzifsvScF+Xz8jmdNOkNCiw+WvPkeUbIl08+lwuoYVGHik2AmKRK
0OqAEZxtMTaa71tx4p1jjciYOV2+Bs+bzkIi3REeJHqbOdUt+6oaF8p0Py/5gc2DmRZbDy9Rbmit
QIBjxMQdxOOgyidIwQf1jaWfc9nItr+ND5Q8Zgz51qK3aP4yaPXqf6hO4uBC1lKUk8E6Tiy+Kjg1
v5nFpTqT/LiA3IcbFfdH2+3vQ3qkjrAhRNIlU2Gzg4t1FMZzy13Bk+mxlinQTGTdgIy6ZpC1cecy
w+WwWRosu/GBYNrPbD314jP4b4vJzuiBzyqpqY/jXpHgrMxl0fplkCg163dKAsQlxH9A+P/9VDOQ
+XVmcG6UUFiMLTW247vNRXyEyEWjRsyC7uPBlxjHV/slc46KiAC3nerW8MPWpA3xLBq/IKP2uxm7
xhgPx7Z8L2lHmL9uZHUrlnUkkp3RzS72nDmCPOEf51tBSamFQ/Xna+n3FHomapaQMmGKqK3SP4XW
3GoxFkdAQj2tC7gxAdwKWc3KoiCQqujb4nB3BfdDq2cnaatDXFlxkZ1+xhz4/Tr0wPoT/ohO7loO
K/89nkYRzBWwPzHsT6IzoeeOxTiqWwrwNq9bg+o+rFr4Ja0OiQDaasepM4SjEaCrqEbxPQMcxtlI
MHDj8eAUfANxvo870BQx3Oshd/aCSGUQoksFk2uSGvETk7VNXeya7JJ6LNE8X9LoIyqBaghwm8w3
3ylfGiNUUXFGCf6s4EnWxJxKRcv/DsOg6lmE9Py5j3OsIQuPyeztdkV+fxzuboMTCvqrcogc44ME
VZX52G0cRsN5lq+2UUR8uAszIE1EY3u+zEcaBlybBxFP+/8WqwoxeLOLSbY0uu9YD8FKloI2U9Rc
WHlbmBqzcT/PViS1GJWPfBr3sMwMmx95tj2HEXC35S5ohstaAbKmxQIzGadRVsLWKzhsbCbGLjiR
LBdHQqYdRMOKCW8NrTQN9dnY09/9PLwxh0+1Afpjm2X85PiWZfspEIwP1qYLcDX33enU33+5TMoJ
sMQcU1APm4AuZSEYgz11I4b/YD4XP2E2YfmvAHOkYf5GyWzSj4jGLtvU9+B/bi9g+6SkAkfr6K81
MCeI7DADpGmQ0+HvJ8dHbddolFIT1kZCdI6G7tHJn4YqBpFWu9FW7aB7XFBF2vI/z+zHF1oW6dIJ
z7D3nt8Famhbwa6lbKm5hPTgCwDnv+hg8hxWKQMwy95sgNwrBX4mD9S9ZLCyCWme35E8GMesI+xZ
hoAWQrXytAt7+dPiT7PBdZg6MBKFOdfMbVHY2pjWeuz9Cctln+yvUY4F+nfAASCF9zGWBswFdswM
Ok/RCoer+TlwOgBcILexHXeGT/V0w3tujv6w+ZAs0g4NVZjsNy4pU0noNtveCd5B4W0c+xtDejA8
XYGtsBkVaemDJCCZ4q1nwJG+XCA7EDS/dNUyg8TafdYDyHB+F2HoPbqge9+YqcMjUAmjO2HlNIQ3
Jpxa5hTiKkReoC6e6wGyKtbZPTppLAn+tM1oasAIXe90Wn8ijqErg/lNUE6ggJnpxHGc6+hL4+Vd
5awAwl8neOCvVmnnNzqwDgukuwXWzeA+PznBhZnOHrk1OJUCBRU4/AwusqmOkEXoVNn2bd+TctRe
/LCovDm5wISuzzJl+U9sEG+pmtHBRLVxmycWvpvJYJ8LuGFPPCYPeHtKw9kbyGVYsPOQCSpS7T19
wQfYDYUIS6E0ANAekBzEmn6MEj7DFVsp+9hs+Z9R+GCBneWt3qBLA25lQUGp5jBiTCB+u440lI6h
yyKu+dNtVQwnfaHjbsOLI/4QvW0MICw75jRqRWjE8zXPmwWP/axg0fT6GY6Gnv0rJ/m2HZ0wyDRU
lFEiA4xJxr8rEwQQxDXXuuPgaG0ZJ0FdQ01DDEHlKpI66oe1b2qvuh69du9J5DoxaUIAJuR0Rt4j
bHjgdW/D010SixCt5DjbJ0Ywb3AAJfIHoAXExLyrDNUs6YUpA14MnI48aXKRKpxMUcRCGXpqdeNf
w1Hge3rMaDo7ZDM5J35r8m0P55FHMuBt9MM802nx6eQRLuwnGJUwzkHgl9dNvNv2owY9lL40GoEZ
wBfsNGY+PWWD3RtJn7FTKXNJW4cupJnN9dltsOENVzSY6f5Xk0z1LDXXrfDulW1sLzyXxZm2TaKT
lt6uAV+6H+J2rOKUDGbg5c7thw/of4PDOx6GVX8AUnCWQPWnmrRTasYsFHKR5qTyFY9Zkhx2GPG4
HOky+vurye7ZnmMf/T9hG7xYvCTojzo+PISPJQcbRLFfL9gsctHDwcT4GapjZ4qRfe6lmIMBP+HH
hWO8Z/tf0ThcXwmNnzyx7RxymHwMfGCElMVUi9zLIv+IrqOr7WsWrp7FdflJ4ozVwGf7W5j6Orgc
IMid62JojlFQvVRMDO7UkuITlwj4/Iyhp6Vb0Mt5eUK0LnuHOsMaiWR3+T2ND9VEPDC3WAvdgUP2
pHeOucNJniw9mnHdXwMM6laU3Cw25aLuGAiUs79o15L75zF1TiBRvRrJFHSh7DCViFo+yFACWaCl
xssm8K1TI2WW+rcp58tNdQUBik3sDqV97kUoQWgqGRjq9ewe3Z6gf1s+RP+ZckUknhs0fAtOyjYw
WlQRFbWsDzIZyUy4UNg9Kp04FcQo2LLvn5JTN+rRyrVLLB2dJr6luoQoTDsMwfUtOUiUkjIb9dSP
sauxJtw5G1I5F6PgMzjh50Xa7ptgR4+srTk9LTSoC/p6YYqxTXIggQNwKpoxWPHD9/p9eSnrreg4
Y9SKA+iBE0JCIRCORwJqKvKqUpWIwXHB2D0T0qwHf5A40JjL9spK7dwlrswV2kfJRu/omVDVw7RC
dzEX9POXLIZmU9psI8XQnk7AGV0OCHh+b2e0yqQLlYbTvAj0Kb6wGLcJjJEo43XiIrTgoU5+jMS6
EF4fdB5r+sldmjXuk8A419aeV+N7SamQXEKoIYn+xO9IqNnZGNMWa+cRamMrQpfkMStw/p3WtF4u
MhBTr1pCudDNxpEegu7QXBs8Bxet5eVQ3Db9bK2mhEliJ9A3mZsFCPiiIuMqUsGzQB/oMxjh8pcw
dFG6YCzk9NyPt3sa0tonY0dXdpmsbUjxJn92lQGv24ObCJvpsuvHKn1p8icRoR3rcHh/hGUDaB4n
wVpoLfY662t1FJ+sahwjXBqfennWimR3fwLbPOuQ7cDN1evo5R3H/Y7Q5VtUXiquoX2GKZUs3CHT
PT9ir/7vrsmgAj+BKILkeUpD12r6qQX5gaxmFkfnEp7FLZacPkZAYqhSDZuj5fOcxqS2z52eZxFl
34nbKaSdCyaKGVV9lSvy7RmX69Vt/pygjXkbRfphqK8vIoCJATgiDlXY8AO+bIYG+Gaz3Ap9Ci2h
pSx9spBweypgfjtDluPwMVozfJxGIKooeXWzzU9WolAnzJ/jbMpjcT6WQ6KXwAZbh/hv0PKMKf+1
sjKyOZ5hvZi0QI59gEc3NGcr/jf9vWPykdMmBkIZH5RCG1j9cNyfS9Lc0we7bGiZ8H6+A7NEoiLp
UGyXuD+fFJ8Sn00q0XSZLKaKaRiBBgpVjeNeMkjeQ7j3yBzKEF818x1w6dJpVbgLRTyRBBw3FDft
T5Z9u0/haGS6uW5he5wKonbGpg503VLIqr/U+wP+oJz7UqpjtKWvt1PB+YPZUumYoGRKPADWMzym
wMibSlT191uAShHhHHZavhjKAV1yrvFc8k4GBrh0ipsrAgQrkCsG/p+A5NHvuSWEpiaWySBALlbw
dIYTWZySjIQq2bUuPnSp8cnfb8LVEN0l5mS9j/EviWBfePcFcpji4aPJX8XdRL/HseuamKGxBOsQ
pgak80dhw8S5jKYcUlPZM8BOBrj4PC+umxk8NgEAB3xVagMXW4NIQRy64xwWn6p3/n2WM3dP0KTM
C9BHZr341Jio+t9HmIuag6WUwBNM9eiE9MYpNC38NMJ/ijw4as/HV9JflRASb9SSNLgTXf9Mabvn
8ZdhDx9PFmxA4CrOPJM11n8aLvYIouvm2G1Lp+FaGcSO10nsM5wnc1UWMvsfp8UgeLGYUfD4dLxG
YagqLue+AWu7orG6JX+OpfuAHkG+059dBSqkak9rDR0unB2boHytrLGw+zA/zFi3pbWlaNQcp3ab
PiLB6u7DyET+a3GlRKZ73S8Ms6ydPdW4nfMyUro9EI0znl7+2oH7TLqXK2Xq9Zr3F56vY7SY5hDq
fHnYXTmDaExbUHD+vNlj811A3swMVp3cUtHiSDBVGNOsvj6SNvENtciyJKEdM1xqQKYabqe6a0qH
b5WZJRa6fPeLGkValS+AvZFnv8jgLSW+mDvfpY1T88BjpA1Dbcy4uxNfUX6RWP3iaIagSRDj4s34
MxoysIigb7UZksgIS2GSzDm82YkEmDmGA1VJB7S0X4F4Oh567nJIq4MDBlzsU1fTEoGkivyd6tFA
buuS7f/yfENwPoEh3en7+0q/nGV8i/aid8m/hzcX1Y5iZtmoRt73Qb9EsLRwOX9ynujfFJC3+lep
9gxMB5X6jRn0McIt1J3SCd610tdBUG9adIDbjsltkyFI5ddu4IUIIYMTaKJqFdMOfGBTUroaic/a
za71Xd8Ak0+TM6GHeA8pTDX99nKOz9Y1qMescThWAa8/Cwib3HCa8UbgWtYRONeNKWI3689MufU5
/G4HVeTsIumVusZUzJbLME89JjEBsNDmreTa6QfdAyJSiqJC9yS6rTJfinIZzQi+qLa5wi+WGPw/
stnHCRoASrDiWK/UjQV0M9f81SROSEmQKuibEi/PsDN2sGTgCAMlNqubomYEOJZbcZsNJA/Rbtf+
+NOZIwjWoFRRmGk5cR2GR0rFHJv0cTAcqDhdaUm6wB2DAvZoEADYNSIixyv+mBymMDIshwl38Ddt
MkuEhczt7/gDvjB5KEZNkh4ENPOl303aAqjnBWzF8inU2wfvGJCAFnrE1O0mZcx9VweiuUktLvE/
kbeYSwmGWOhg36NCNPOaHd/Qvi42wT+A3VMNBGLSZWoDsH4+mMyPVEYpquCWV4DYUjjKe2V1mlGd
qyO0OsqaqsXN15N3ZGssuuPwmVrF4Qbu6De7vykentzH/4yGnQykaWV8Mf6NhCHvClsmjd4NRtmR
r5TehWJdknBJO969IkIlj5HWK6tEveewFpVoXyRF4hk0DsSiU4XF8g6//GNYMRVQKIMWywXIPQRI
DITL7FslD8hEJJVcb60s2N73jV96/gaLovFTTGGOgB5l5xR4HRVI68crsk00etjK0MxPOc+k5yjO
DsUFg5XgDa0c0j1uZIVDnv4JT6aQn0FCtXR8VyZtNdozY8IBfH/u0BQ9ZQ7rUdj2XaASkCQG2MRD
g3cGYG2KfeRxNTYG0eaWuUtSq/e0XJPXsORGLL6F1LLmomXtOroyBtNKlSQjV5lIwZOuPPqbWRpb
uzyTGgBe33ESDhBRCf8veapt7U7PJKsd/Zu+NYpe4EgoyBW2ld2x9DfbnEVKLxW4iUV5k6KH9ASe
JoS6+pbfTjm70kiwCOL2o356MEFDRU0OcRvZusKwu1HFJHbYe9ooGiozr2sxbaS3eRNozBN9t+Wg
qKepG9o9cXMcEqMhfRu4w1rUGBoZZzOA2xK8rTlDernk5f6OuJZf8Nu33V5K2sTJ0Z7sVC0omWA6
SU/4aZZkBUHjtTv4y3M/qYJiiGMQkrmNKxV8Jnc0nnrtrTCgxBPWF1/K4SKGNQKTCMPVFb9YucbU
XDiX5ekfiMb1/Fx47xae2SBqSFEkIunqEVI43BXwFdtvoHbmyugZ6P/7L3CbXTZFx4/uTn5WNxzw
Y2e+oHAtDtAsA1Q+WEjt+CkFyVyT29tRv0ssjmzH/QKYHwt4iRL76u2Ve4dfKNTh2JmPhIQMnSNa
PkohRfKS3lWMM9lBmfbMCFdXSSAU4+GHQn3wsMM92uJad82ZFk1tCrpgAyU6Y/IQSvItT49BVQAL
qKHxg8pcaKOEoFLMBqkAnTOM3jC7vjXDvp4ZDy46GPpMRNNi0Z3jwzzE6tYQZ9zE594cu45tpjdd
D70wenNfZtD3pfk5MtMaVQ1YYSxSDPs6pTAiTtJCk6TgcEvM+h/S6j9bsJn6bQw4Y+GZoa8kGium
Zs1QCjg21iJcy3Cck6yXraR7RyQdfH/O+xO9GHTG/uSl6MwWK3t56M/gb6mIvvqMpdlpBZtHzc/T
5+UZqtvUD5ifzQGtMMc0EXO3vvgV8mc7eQ377oGI6e9MJvptDaU69rqfxK5tzZEAp6l0GQucmCs/
cu5VmdVeUwHnbeM8YeEJhArrA0QOg3LDCxtVhBrawBCq5Hbwl3GeEwusvLB2cujwOmI0CjtvYGgx
itR5LVXrDTBOl6k9Nf56BkUv0kHdY4ok80vbwONkVlJ1CaycZlffHeKsYwoD4VeExh5w3MfPLy3E
9URNVGyCiHpcCFKErCfo1R6sXWr7pgCQR6xzleXivtjWT/jVGlZWycIHn+j09OFmUE3mS3AB9Ba5
Ag/x+4W6I1q7zyeOWwhAeW+k1aGeP38s+5d9TnT78Dcr/xdUdsoUorpDrUvDsdq6/52IwoaW33H9
97M6WDnZynsqchw4rqDb5fa5lIaOqCvm60V/xtOLtbKu2y4bHY0rX7BDfKTpJOdhi49jCobc4SZK
7DelGLSR/3ShOP7bCr5Cckio2BJ/CS/ugfL6dVnZpnfCagBWNNWBpvdBnKM+cf4KF6OvJZzWdr5g
Y/MH3pMGM71wQqUKxydn1UdaoaemgTMZ7UrurPGGpaJDCNJerd1D6Av9wycD29JB5XubQkhlL8Os
g88koy8zYTTXIGW1bjxL1hW6Ysb3lb60rg/xmVWa9tNjiefIT+c9DbYWMsVElS5wguL4Ck9M9CTr
Ep3pj0mtd7s45V9AVVxGyCgwVDV2zezUMY41zzNIzAZHPEaTLwowBiwsOUToqSmHi3FjVOtulViY
sxkQBMQk0RTDhNQPW7GOziLLCZIfodxQj52jMWgXN3zBw7NH/uMHuVWFjOGjY7uChPfqvgF9PD7O
OaWvSdGZXqF1uhh9VhmLYVvHSkhTCnSUlKvEk1wjW9Q/InnSxcH4B7PEESSwpgT+iacPum7u9xL4
FRoJcuLHi8MVsbw+Esnqj6HWTDujgVfhIcZvwV3/eEwRQuz5706hCvH4gTygPD9fuA+r86Q2eFZc
dWZfJYDTrXTDfZ4ez9fc2SxKEtbM4+cZz4OvBhUWT0C5bWJthnGX2V4AmjmUD7IQ55ftfv6p8qxM
ecS36POJAJ3KcCxi1PvIxKBNjvxsLZiGH4mdtnt41xsFB/1ZyHJnR9Amw1RDz0cFkMalvtt4A1KY
BApyYwSVUR9dfqtDKvx1JiWsi5V676MOZjlr54qb6fd4JU1qwsulDqFcv33D4g9k3k/PRtxPNUgU
U1n4qpMEGgUCFbAICZRCw81CBmqrt51jh/80oSfmrXRERBY+IbeqS2w/o/aFDDk+94LNHB3FLW1X
YRQuN4e2onyfRoxm3XZpZgtJnVLIb3yjLQTeEpN4ErAXlfb/d/cVZaUfuPytUbnOk39wYJr88V+8
MBRuMZbM5PSxzDq5NWqFpzxoegZIwZE+nf4zxhNmkPmR8Lj8EGoqzx9fW5gjrKTUlLqo4JJXrKRg
ru+d4UWP+0iXfgEA7DEbaEWLQmuKsWG3LwosKfPldfdsfEt4t410pQMxdwjn1Yfd5F1DE96uTMf8
xEEflF6g/CPWsd1EWZxD97mYbYogE0wAQWEo8mpTquKPksEMGxo6YdEWf5AOwknRjNGI3pdU5Ikq
diLjYPKF/isFnM5qWN9J3blzPl3R31x7rbfUMJOzCwfzTAfW0G66wNNnjaecPy8U3i2u0nVZK/UK
dGMd/vflUw/bbVI7SEyFx2XNA/j1PEAZzZpr9rIQra07X3KrXFu/P01QIyWEq1BM17DYfrHk8oKs
q84FZDYfMGEo4k9VlRtfZxV4YXsomZuVTZIbV4xlVElFQzZUYfPfmupdJNw30lE/Enn1MloWEM/+
UO7dQwQi0GRNzF7ogR7y9YU7BpOe1m/47dMz2fZt8OQ1MNo1Rq4VknKSxfzocxGOxFIfRZMa33QD
DhlCXWT6WxJdBIKRd+gKWpA1HEwX4IbWYlsIrfgkS7Cj+jomHnbIVk5SHZc1GFotFQmt+Dekhns0
JuAib98u7bTHdcCapH/s1NvaXBypyFSAE7HURvv61SRBJv5w11U7BWSXwmg00mpzkQFoD4ngLClg
uiwUSO60eMDMhmO2Rs7BFyOJut13OaLvjp7HrBy2UIsEe/pnovVMqvX/iqBwe724viBfK0EE1RZh
ajSV232yk/87DRl2IEC/qqV0IEX9FZhJk1wKG2R8WJ6RJQM450alY4eRwAQY0gtnO2YjBxlPmSa+
aCWvj65220xM1AtYY6ntaDcpghh1DHe0wyVcr4fqO44MtBzP7a56fU6UvddHW71ik34TAtPRKeDA
vTli+UUceS/l9lBPaWXo9R+3nf7/ZzJZ4QHvWAUYfuietYh1UA99k5QSZPgwsAxFguzhZZ4dKPc6
6lLEwQKbqau++7B6FTwXnk//yW1OM9sKo7Pz9znu7FXaAv+vEniLfjRHUYfE8XlBwQgbc3t5mX77
BfSuJD2tSDG/Hpw3VPzYh+WDpg7W4zm4jN216wFxsM7aWrGd75ne0wk5BqjTu3hRSt3H6mMsLyeL
uAZKzxQHaTzOy2R1s9TsNcARX/Gv991tBTkzfq7iPHLec+Sl/LuZCLRjgfQKMH5oklqFLoFhBFZE
ikr7z/k1yqnLaqnAEFz4cDZ6xqWQcDpR/opwtcBEDxeWoV2umJ55zgounHb0uy6lIeL7GeZv9bO2
XVMAlft3y9CiEciqf61BX/QWQ+VgDivax6MgFkRQQ4DRqhkMjjlR+WlTiRZIcFwXqk0JbZF/KLYm
CGYGkPnURpuHEGXsGssTtsajyN+W4FYnxtljzmnxACuJZngqh95NeIoz6avTAZOa6g19/kP649lH
S6kXUYxDmh6fi530npMPkiGoYb6ds0vRqTH6qznEZF2VHhYA9lrVKnXyfMluHHOgvNU395LFAWkW
vEy6pYbO0aaVHf7/NUjsIVwm3EbE1PGjGGkjv7axZvJGheMfIH+WUN76xXHa9t+MSs6bO38Gumdo
UVS9FjfxcSCCMetYhMI04XhDJORtPKG8gDRmZ+szcNwI3o/1fDoHjNwjH9BrqDnp2EZHGkqbsWo4
jdLaNKWwCioxacm8zArVjEChJ+KI6Pypp/xEJ3mWPFcsv5fvYc2bq0VhnAkthTUbsqdBuUHMgoBD
UENE+cwI3yPlIwqb1Ran2krGHMyKsQP20BhYrZ/ZxcYqHBQwNglIS6SViu/AXCzw3arx07ZJ+/2Q
ZgVw/XFvj1Kp9YlMGnSSg0nrIB+wxJjGUB01L2lMEtm1SeqXS8YBM1ARPTKbh+Te1kxooP+rFjOk
pvE6oC3FRuBM7rms/RQDOucU5S4U1zpD/3xhx7mMyBvinych5fu5VdECu3HCT0oBMu/xJSah4CHA
sk6FHTfD+khOptDIN2TCqEOXjjVUSBSKVWp6Hn8YU5Zbqnp3vFEzeu0HDUHWSIrZxBkBRuFo/nOy
OwSHneeeF6FASYZA7ZMAdK3YRTV6aYtbytZTxWId1WPlcXAETlwTTXpVc8twZJWC1xhvEHIuObxH
oCB9pqhsIP+IpBU1tW4KbkOWHdc5UScbUA8Mh7xiNmwFbAV3LK9Tsg5QVmmhWs41CWelmAky1yiC
8aQ9JaEqiHNxX0K1t6TgXtyl/CmCVYXN4jrYrSOCamYtqaK3XGxPYCNYdOWy8fiEpDT4CvVnyzWR
GSws2LwwYlFeu8bUkkxNg5wQBFM1pfVqDUgz/whTGU6wWFUMB/eWgm3wKa1MxHwFLSDSJ2hmrDV6
842QeF2zW0ZALN8sJNUfQAw+I43R25YigDSgLL3VF5lID4aoltm1unTB/0sygjvrOscG9E8qkJ7l
xU/7wrEWsv131dYVfIXBIjpnXXF7zncQh6nHcNvncFbh8nr9yStSf2MjyK4uC2PvICOXr/n8wugR
UPBqinkULRFHEjbw1lTCcIlCUiiDuIccBAIx+PSzVlo/lwLX18PNmRmy8wUE1EwHEPQxOZ9Qs0JW
AUrNOQ0X5BOQhotHAi/x95jGzTzSPyBO0YhvjcpVV3mJ2hc/RCNdshoj78ix2mNBFnAciXtrbq7w
r7Agg9NePsYmi2IO7bbE81lhnwwY3nCgmgr26n1Ixzl6DMdEOideouXLkLZf4Occigc/KB+G4Pg8
NSxEmgUdtccr39mbhXOcjfD6fUVYkTP6y6vtgunQawvO0Ucbq6IxZ9JiEIqa5nynlhJ5UiCS6qRD
Lf7bNQYxRsDbNxda+RbbbUrcj0sTuFFKwKKlQ0jKT7Me0BPP/RPcGc/tjlQGOKNa/GQHHFkFaWwI
9pQShDRwZIZWYRNhX2Sejj5B2/QwL28X1R4SPjmK3eJVIgNceFVS6ZR6Tdkq9OoAfW+1IO09NhcR
VgIwpFR1KVV5o181vY92wB534Th06sRDpZsbMgIYgJm9dqb0Y/mVBTzFrsIoyOe/bPZpNFyO1RrD
VHT9adtjHvItnpmzyjfD/PUOCqLodmHr987isGHBns54xgALl+ZLRbUD960Ci397UbdTE0sQIyLb
uNo3bzWi3neRLLN+zqM6HUmMqqp1zFvAgQQb0OZdahY6Iz82i7Z3RRe0KlcN4c7elC7yrMq35F8E
Q3nmqB9fMsEv5xTcHzfhcKNXgGTmJNCq8jQGWi60uo4rar56wypsLSduNbEeGd/EDtsne77xfaJQ
oqyhdOAAlqqqV04LZj/ErWveB8IssRvsumLylwDJvTgM5nShFejnwoqrwzcJ73A/sA6JlXwuhZ/s
TF3zGJPDl4O9odAxFB02ZUKFFL3Hv1i7zAClGPeEZv8EHovzcC6pG0isCncvq2to0272AzFnwMwu
E5R06xvs3Ovq4w9GC0F5dft6ySCX5QA8t7dGug8yGP0rvN2oBdSg+d4wTomQTC4DF/WsBFyZcRdG
wzWh7W3FWCxtOhgA2uDn92JF8T6Un0wlvsi9eV1pPuVHrPyklRT4YPzgMOOBnxbgDYdA5+i59XdF
5DXU9igdVpKow6N0o85mU8ioWDuUMmsnvoBsT4nWdwwJ0ywaMwjjVLZDa0PmiYmhtXvnt+2lDUxC
HyAfa6I67pyVgVAKoaraRSskAqoQ0ibstwkBn5J8o7Wp4dJkDJXh8K3pDc1xSbIcnv8fQwEe/4Jb
Z1Pe5a074eQAheDZwcy0HQkAyGlB7MIQLBkDZZ404JyvuNL8ToPOpVYljYnqgMzE1R3IqCgJFO+p
7d6CjGv/CegzZ6t4700x2S0tKA/wo4+ijZ0VkVxk8d0CTceuximuuoKu+zW35EGdHKc+89ceyBAt
5A4BL0fPFXkzuVkIrwCvoR7VSf3v4dt+QoIe9nVAgMaZeovQlejm/Fu66/q976xeuG1tUDhCHYCf
Ir+Ijm0p+yRffc7RW/1d9cH9uRYsjWvUzbynGK8Kc71yyN9f7DqZi1NSlQd5DNMTRYsfDaG83erq
vkcUXDXGErNE5K6DxBwA9dvyOtHtvJ+Ykz3bDJqK0DPnFlz7Iw2Py3WXnBm2pwrSCsRa42302YzN
4RuLYGJC8YF6xtpJ51ACmNZ7eN3D14h5kf13M6q9VzNvBe9nvruD1XcrbN5jXvlI7yoGHGPbtzwc
tad3O3wp3xyYCpEzVxLOxlAdxTNLm0uMkHShTY/fEVwmRJlXvsTnwKB0v44oSkZWwaqpm4+7HyPY
U3ImSpuPlLImA6by1msx5i1tPBs8YbNVypsj+AGH0RP0W/PkjtQmLqD4eMp3X0cpceOb4ndiqnnF
sWo/eLtVyg+FWD24KNsxGndPkLbH+ep9OR2n1J1+3v8dmg6A9WWuB6k65zdCbc32yzR+TWzArZKZ
NL049UAkv2AllIBt6kSemuyNBXJv6QXkxibZFfLK0zTrh6LRIa4M4fuSMSjUW6DPt52wsWdFz+Gl
BfheyKpqm4aj0m4Z9Q/L29y6zRcj1jQjTkZbsq4W2Mzlu1PiSkAt9xoY7Il6/+u3yjAM+Ahj9WVX
i3ezEkfCO1HyI/HZ6W6iFn/DfXMtsUzqlueh0jogK+5SKUV+EFPQCRTedEgbWknzEi8aKm9xIHYA
j/7uss85pl8vO0mLCF9Tw54GN2CEW5MbPfVEpjSB7KRom2/hh6ltitxKqqM0oOfkf2ZmNpmEuShx
F5EpUJR2KLWh13gN7i9XIsGojjQrrOiZj1UJerAHNKyDR2Ekks29m/3yibgG8qxnSgrvm+zlvZVZ
4JpHYI+MSLmSrt52zWF6XaMqNuI66CyXcejfSsbeSslXfCdBxnDZfNdWMvGr3rlfgLPCGV43unxf
bdcZQmMf+T/unBRpnUbcrOmTMccdL6VrSGeRlvph03/4Vgpkiq2/KoNuQ1GZY+2vT25lmFftddPM
FW980vXaFAZmqDf4xpQs54V8dKvH1EsMWQyNgvnNK8dvFsiVNkuJ7GbE+EwHIZZmlLYCXq9EByWK
LE7vRedGzIvi8lVlSRTsDREiPt7qip2A5YDkqvdlSOS7eV7U3hp604P+kSAV+4/QI+zKhs+kdBrl
7Wo82OkcDLnlc0ndLKwxRCPHSX8PLy/HrNEcKgtajiWVqI+nTgyfK7Wo6g9/v0E9VHCg3wedOKnU
8Uwqzb034ejRcARZuJiKdd6N84GvHceFaShhb4g3OtaQKprFDwUtJuSCxOIsYFXGNASjT2cLfQll
QVkZKKzajagHXxO1HIyVSjkTMUwVOBnQWK1nsAytHqX7mLzx1HwD4JlsG8iEsZFwVp2R/8xz/muC
dVpeqhF60tOOL2ySQxL064mefekRmiBwc2XtYjh6TYMtHmf/Z1A6GZr7iz6EXN5GpYd0B3J7OMsG
20e6JVCOO3xTdKOBjsAyeZ271fB9zC6JA00p+FgpmPEh5a7R50Lxqwxs0aNPjjuCXWObHQDw/HlZ
XF/WOUdAlPdEeeznno8PpyCR988hLogFyCaZgYMg1EqiCJvO8kOm/QFLCy+FW+SHmlZ1/YT+4b1G
BRjYtYLYTBRahnyWkszqLF+WYj5x968bt0G8SvfEofjsj0Z2s6kusJ08kLNUY8k7Hde4DCWgCBdw
A8C9v2geVZNMVVB3VFBSWBA6LZFmg+fH3u4JtDJWTpwwEqgO2YpXOrMKAIy1dKDOfy1bsloQICry
/bYDH1vpZDlx3B2pYVRYCMQfQHY8nK9Omw8dH+6vMa0KILjOy7Gp6tVEFbuHyuK5A8WHDiYU2ac8
GFuquqzhr0mPALx0J6ZMfspMpjETZbo5zsOFZtyEP0ydSD+ilDuMLW8zCneSpkhgY3nGJ0PLuujZ
9dSsU0jV/LDhflholA/Kr45/sj21DCVE3rdc4lPdcCmzRZ7yRpRZxFZlbWJZVhEcrRParzJMkW/+
NLdvwDys+SjvMxhJbNt9RqaPHJ71+9wWYKhoiOX466zAy8rZGU55QFzLHLwpBzxTk49kqBCFwUDf
pdt8FDp4dOW6aH2i06DYy2kw5s2i91disyw5SAGPyTqxwPHzjPJ7ztQ3oTpkc00MGoiHOkcFhIub
SZRiWxMlpXjEo0X1AgH3gzAGcvKayOffPIC3ZdWMYQKi8jAHd1unoAfZCSpiZmTsOSRQzkr95tBO
RyT1XCHA14tvuHdtz6wHQI5d2vMhZmeoqaCYSLPHh+qc3lvG3oqzOfD7aHxWoiz9LFSh9buro3W9
JDfJKn0kTYpUSPBvx9NlUQarR00JckfmFgXjnXuCMdxHGr1YSK93pQ/WYlZ38qy+wN9DQylXs1X+
d33h6xdiVzhCzhdKyJOOxYsABWb8cJjCGZhv3eHkfzC31od8wS7ni6kI14JrwdE5sIoxK3tbZuja
VBIF+jFWrRQOuqXOJyidMwtV4eYD7P4LBxI7byrX3kRls2tQo9aTUHzgdW5rNpzKR1iQYYRj7lpg
LNcNOJS9NSvy7uEDl/y7b938dwbod5O6VHiKj9Hd+/u0PoEBEfW9twRpes3X3WiLwkqqR5//HcJs
AWlpmlB2xwZUJo9cjM6amfiSp2fyEKmTJuiFU8O5f+AKfEQX7Q7ItbeysLlH6UMPKT7PvsudzsXA
m3vVFp2MocLvf5TyoBWMPVbYo4A8B+7S8AU6sfiB/wd5O94ZYXDG+P1lo8U8+pQcpWkL8EcLY+Uz
6pfIZTgadYDVOMP4KueidSWBzLfQ4cczso8UQiYdiVn0zg4SLsKIeiUk3/GkHyXDrJT5LK0EmPWJ
wq/+WDQYy6/ysYViu/5f1JS0GpjlL0TOL7gHLyAq93YGSs49n00Ib0rnItvBzZHTj0oqrhiDbbV0
R/JaSdJPSnzeKs82RsGkmlZc8l0wuUV6mEA8bB1YqLTy9/XhmP3SrPyb/J6D9l0N04oVCU3pA3jK
iffzlQffZy6swAFNOn08MvyeT6iljGaDju6puvz8AUX9fKLRFYl0XMMbDuYo0Y72aa0ZYHle5PAY
xtp+V7Cud+ho2D8MTzDSvhdjbeMNO5ViFQfvvgVszGxhrunv8tUX0RMbz1gaA220VFTlPodQGtrh
Dc616kS8n0aoisqw3yuqmKqvJVlFJJlAyJ1Kse+zvpcOSiLznjK0c/8QGotZmWD1Og1ldjzQFNyH
RQC6oeA1NbDdk6itVurn1Cxjqfuy/0FEmqLzPaiWaRHRNBW0UU+na9A3hvlRgXlqMfbGYDu0+Gfn
LnLC7KzkX8v1wVYmkvylJR0cMODLVIs9BzV6L79uU2fWrr1QANinIUnUIwuO7q1Dw0yXsl8S9idP
XoaroJEfVz22ix/AYjKRvpEkdHEGvPRT/CF4vq+jR8pqJIMTI2Hth7dMRMTlajy/CdDMRE/xioBW
Ec5GwDNBy59jhrSbFPzde2tVeO1NGh+8k1yAmoDEb6kLR83fDdfZTAA92othkD/bOpZajEOiSOLv
3dBWgqs5Jb/WKAsGQVtZOyHOpPJ/ZoeT55HhYjsPB51g2khQEn1XAIK9hjF4WBCTjY4q4ALAot/c
hY6tOzOUct87+kF6UeiFJhlcOrlE4TDcpn0wd54C8NsFdS4JjY6uyfAidPs4s2hHn8vZIz3TVINp
JvUS3PUC0m05TgRDNoyU7s1oOAYoQIbmL+Cjcs38dljwAjrPB6jpl/n0ODSjudBu20Tj5dh5kpql
atUj2judZinH2rfXmsxJJNjLt0yI2FSmxM0/cxuYkS7kZ5ERn4ZTH4dWXbWoyjwIrynGSM1Ihoza
WCWQZSW+t/FPLafC6uWs1LAollUZ45ev2TAG7ZfCoki/rkYLt2qFDZZfinuhy6gXs8e70Hn/PHdK
eZLlEEr555scvzKrcB/bgSViXp1n1X3AmTiB2GAIWf4pzZ3jFF+KgDDDU4OQXmT0VS3EcJVR8yu+
NIDm7OHYTJz94J5YVvMaRwESfB22V1Px0IhHh9XTFMLUNYeonp8RSdLLllp1gVeanDefbvs+EL4V
2sSo9Fq/TGRVvVHpRJQMYSQyEXAxWbAawQB7Cq7OPNW4ZkD5HKwIw9dXxw+uOAbkPKi45a6QFdu+
1zvtDNHmMibh4tJzh4Cr/mPUOkE3mqsO9IZMlwbmDlrDuPkvzRFL4tWJszCs8cN+cA9RBZi9d6k/
0cf9jUKrSHFJqPf9P5/O85NyeY8h/eS5jZJJV7kfQq/OHoIRIcKsiBAqU3rCZIIVVk9iNYD+/L7O
yiSQKyapyBMEbDFdype2gYQU5Lxulbul7jmG9f91zKVg2U7s9vf8UVrOrJc+f38P9D3QlxZAISaF
hsAv7eetXAtRfcYs6ZYSqhG/LdwT1LDvdwKlLv4AQH7ZOABB6J6veTwd8mJkJ4+k0pAEBojfz7Lg
RzNUH+eiDNq7rmzjYq+tfe1i1Ni580gOr5/XVBxiqiBOQ5jhZSBA0dl0CsN7IvkGK17oBPalxdSF
owEqMh26j+Zzfi+5L59zovS6GXgpv+JY9YKXPuVW7yA4YNNcnOW409pB5H+Z3NqOzQl7t2VSprxA
h3U54F4cmBbEMowyEayXMUUGjuc2dJwb0heVgr6M4xdRbkcJ1WvH1zjtRZYpB4m2K2Ktw5hTuOQA
HGKAwRjHeMiHG3PsiZlrlMn2x/LOQ7/ZP43OZUUf/z4lxLgRGL7yj4/PeUZ4GYNdPY3bIhrcotU0
Z+xoNkGFlLjCbdjlZrI6ROqO2EYy4CgEpx9iDVlEPHzjOeHelGldF+qGfw5ao6SjMl4SFr/VigCn
whJFvK7vDKP9kP9dTwhvh13FUuu+Tya0vWOp/RBaHq5ah2ph7nMYJ7uixA0SYbZS8ocbkbN+WcpK
hbqgI8HsPlVpUNAChZ+nHTjP0DweGlfSbGROENUksk7BvD51Kv/RH9lw/7XhbDSBcOtJttHjCp9w
Wsos6dpZC7I4gwzjMmJNT/xUC9FI1/29jRbMPCgXjJFAPwBh3g+Dr2SgL/fzGuEy/AxzfjIY6D0p
/1bxNN5x+SOCLpro5mEKMFueGPHkewds+rmiDnbNzM9Jf0fg7r84JRFNlpvxhiTt7FKNy7lwoJX3
OVx9B74vgV7LcZPPtTFgXI+Xfre0KXW350CiOk0l9h25TdwQSoM8MER3yVyVIDmevOq2dJ10+4Xn
zfmXrcNF1AXp0om8VONGA5B40QGgv+3qSEk28hIHsjE1iQ+ZERvLq1bJB69xWRZp/SC/rN1TiJFI
rK24wg2OWrdhaWMP0Hxa14frnGXGBMUDSzdlcId6aqq9aiLvdCYGMQD7utNmIOkA1a3HrxJOtZH6
Xq7Bg3QgMpClHVeTyCcwjq6vmQDRm4X3BDAyFy7qWVdf5YlS0knDfuyOG05+YLkm8wdBYZBOezBC
f+orV690acJVRRoxlu70oAkhV3tRl9V9WQAfS96+dFNx6BuNFo6KS0RZhX0rZ3T/iAStZCr8mkoO
kO/c9aVrEcSNnHLr5ZyN7Q+2WjcUL3RRBs6Dq8/yQhmbWJnhDRRky4qFiCBHt0bziuQWmtYDPgLk
FbJKATTLk0DJnc3lvssylsBpBjggk7ls5Dqlp3o8sijMVi3WOAl6qvBZE/C29pLlV6gVC6LWRXqj
MUeFdLer6Vbq+aVZqkdMOPhsYzf/0vKZ48C1oGGMwhOkIPJdt8fjwrNJm/ex0cTZsZS11yGBes9E
qe7pYwmfzHfUnhhcAoX9dkDz4A3Trwbe8HN30FCyFOCvE8QhQa0sfa4I3RfnookE4X+78sQIpX8Y
wUJYadxm2ZTBDX28gLKc7hdWJ403JoEOs8AYP27gocZPhz2m23iGx6h/yfl3tfQ9pM3Xce2p3cyZ
z6ygETuZQmHzmTTMoBOI+NS5hrlZqkQ2U9UkXoZXsIbqPnepmtZDaPYeQ7mWSYnziFxWNhUy+JH6
3J5Vi+m1Eiyct3pvBaXxvcSVp4cLy9IWwrtFCtdGcJv5I5IPZ8Xp021ABhyKMlLKOQsTyd17X/p0
FcQwlazA4EDuAteF0q327CER96Twnkt0LRq5a14gaJEe+gwFFUwK1zQT9ADrh3OnPe75g+uyoxwv
LN6eYmucpKeKGHqILdmeNsJeP/dYnumU0GO4hHojNqv8x1laLVE70qukQ+NhR8YJxjQ9kINiRkwv
FNuM0aWaIP9elL0RgC8oFUQ2TX1i78uneyVXe4bK9YG64+CEywZ1IYfvCA10sQuNH7jqSlKE6orG
Ems5wywJ41HotaWeKl5j35zIasU4mciBPmONkFLymvLl5uVaM4K4r0wxhKlXMQeN+RfoJRH0C44c
lHAraPmrmkPb3kip8nrM+SW74JdnBWQYF1NNV7IVHrJ5onOIQ/sFspv35Qy61NqZt4XUPbdNGdeL
+Ff3hhY1LbUo/69AoiY6mlJFg0MDCncV8lEtA+3eRBA7wZalsGm17//pyKwacUe+v0Y+7tGH04Xf
vrDX8xUoJVokPgr1nWhSGwc5CcQyv0XbEmGp0qeUVak6BhXB1SHJrnC1T7h8m+PFi2vbFpe0/+be
1Jn0KgfpQTVwTBzlRCXG35G3gt62VeP8GXNHHSVjU3dS0XC5sPtGEvgAGHzPIOeiVW8BBXVTlDQG
VHLMH99JypEro8s/rW6bXppQ60U5gw6yGFA4gLMQX3vc/2bCAKX3sjB5PvQIGVoKhfImJhNyJ8qZ
DjTHJzZeJ0iVkQfntGc83tXptHDQ/wQnnoMkcjM+sFJY5QVKdJYem7VfOtZmrYJjXYmIEH0Q/ETm
DAQPJXnKke5AT11P872LXGBrO+DFmr/TpQ12dreZl3Z0LTFp3Ca4D7Vlz7AVtt70hw2RgFHLg7wC
fTShA1a4mMY0uCRECw4Hd99za5Xf+tSUv/n/Ni9ghqYItSX4+Kk6NNb7lk+GuJQ8vBIdW2eeJwfW
GKNv0XOp+I1SWxFHwbS4AMc/Ivjkrd4txxU39+CW2RBCNOJn+f51A6j/FMY5lUnHpRwVm4hFW8uT
NiP0HpNCv8Yf4ggQ9lQxz9+pC46keTtO82U20Obl6vARvdYrT/OPshw3iqHxzDO/OWDXFaqmUryd
sxYQOUm2zYtjU0NY+4e9Eidm1kp2HuQb+d0wR692jrNn/XIQ3+u9xJGjP3HRkCibQqJPe0L/tEpb
frM7AnFl7CtW1BNJf0NjolrzjYiiNdWDwfRRMR24zwseriNRqHFtIAF0yBHirA+PxrEt8rWtE0Qr
cJGbWrtKKvWNPqaEjjejM7jJtxWw3CS4Yk3ZpSyArVpkhohloRmW+GxRRtdUdWftyhMhcU/L99FG
r+Dgj4Qh8Mtt+7sDe8uRKbPGGfF2uJYf2PjZuFM8/1MzPLgzbJYUXCSylXjEIuBo2dT6XCN8hgsM
8yqkLEpdhwYlp3uyi629BXeKynSR5wCitQMe9S9FHsqo3exYMqmrhgr1sMSA1OZ02uVXdN4Sq04X
FML+9hC67Le24EHlvGXgQ8aVgWZ3PUIUKb2SGX2nQXMdoI6ep18j6sd5KEDWydnwM/jHR9heMNoj
UWirEir1NcWer0rgHEktyLBIg9Vz6jwvHf0w0gRj3oEjvgE5ezFB3B0JVlDMt1xL827O1NDXSfn2
XxwqiDMdQrRHEWihZWuGV/wsAqBwuPGKZl8lB6TNkgjSzQQEX2ukzdbRPwDQeI77FHgqjQSTAJsD
U/c3FtUSy9oK1vf3JnDxr0MxAzhsXM6Wczg5qyPdIZ6SHKDBdJyonLLrq8e8mJ0mxmYWdXxvmidQ
MykbnNbluc09/49mw2BrLBC74wFuP0TSFSize96+AXiAYQPMbWm7xNCD/TNNDVWlcmsqNxr2ukg9
fBSCmJLwX8uViR8mXK6Atea6LtVt8GxrIBfFQ3/cqZLstkOmG4P6BCUj/U2XgMEk7vcwyOeBv+l6
DWqB4r0bdingSwSWf+YfaI2wMuyXsGoIi2riAP2jShL2j7ABn2Y5JrJq90dSW1nN0e8La2cR7EGF
ItOSiL4SQdvBhudrjTeh3lhlsnNRaTR+I0XVH1G8OZQFfSyhXtxErGLfMcrwb1NOvKxDQI2WSTOL
KA4KjqHziNbmHMV4E/ZM6A/1ddocBAee+TqNePsibb7UmIiq8RMv5KSv6+FbAK1mj0KsMo5vgkyC
1iUnhr/Sz172dialAhmrPvIkwVKb+IOJKEGjU9koZd8fT5OEh/q0+6KmYtGsdHDp2R92hhpMAlrz
4MPZ8N/iCfp2X4cGUSLsDU6foshemFXVkKhSTalEWKhnbLNS7u/oGr6wi5zkiU2w7B7sKjtg7qsC
e+En1MdS14TMtv1UIUZ2njaCX5UIDmfLwLz267oCph7KEL29dgKeJTB8pzccjmQzzYMfZF7pv2CN
Jg1RV6h0j9PHTwwntr7zvyDrjiqY/D5Yv+JETCFjwqe09fVKt3Va1mPBB/ptqJvX6dDAlQgO6B6A
kzF0Zy1bdjD7q8zCrpNXvDNFII6Eh5bx1n/Xt09gTr7j941bZcaUg9F4pI9u8uNwItRIPm/bUA0S
MmIy9LBm5/VApnNVMQZpYHneAJN+Rh0RPmTt2E91NG0ZCzFLLFr6jNgTW85h9Uti9yqjTSjzPQSF
w12xvVPljd6DqTG19IEu4Pqv57c7z3E8JdUFhhI/wtZ8aWgJf+mqN2Cp058WniW4NkK4PHQzwBei
WfaNA6rW+UcZNtgNXav+g1pYKJGp7HUZEE0rj6JsBzQ4esagevokvxfOXoiAKP5bImXPHknrOJ9C
6pj/9N5Wok4+DP5VWGfYrjZaF4kT50QSouHIs8iMDR8YP6Lnm+fCXtiWGU0o+IyWse/XPFTAnMhC
1MLk61fTegWW+08p569ggr/k04v85U8Bq8f7x7YteFcL5nFnMD+hd/yMbsPbeLd6S20/tXmswdJL
h6pF5oX6oI0qt8Sin4xnhma+9a7HMPIgs0qu9g3pGP3eJxoo0BHLdgbCs9ETPYQa/3vikiC75WjL
L7nZK8iZ8VL9hegV/3nd8Vdi0ofI70Q5ifdU/KRvZ1Oie7nVecbGlODx5EBgW18J06efszzW/msk
RNXi46fya6uynfiiyNRgeMIs9+ZMP7N1oXLBKLzcxjgKKidMh/TXB8Yo+1XEyru32oByN6s/rzdl
LCid7hCqb4sSb/gsDcaR0Kl5UBgicZZQWRj5kfHXEKxExCjI8Sib0GT4efxUmzeKrdPY4wKXp+WK
J2Zp9+KTDVqCws1IZC5zCS7efw/O8t3rwDKNFu7I5F/poDqWCO3W7N48XDqzZB19fn0C3irNbONi
akvTYK5QEIyWOWEKgXDF5esh93evJNPbYpxR5quw6qOutNC/JF1SPovg0GgdJCuEbiE4aDrrqVs9
rrOevk5ADYI9U093oUagXkGOPPuj+1eON+XI+Eon0CHVtLzPEoXg2t/QyXkD8Nc8gWRlGmHVD84g
tPB9X90k41vk6m3dmpL0Jo0ZpLZqXzYFP0Bdp8BKZUYsbZm8nKKuFHPo6OMTodVscCwCaL4uHi2g
xrm2SB5ivKbbFBib6gcO0XRbayZ8UiGmXmWPnHLbnZnZNHqCEe9x8+AP56ByVJiItRIZaNwg4c3J
qUH+DWV9+gZRKw4iWfAJaK2iaw71yTD5U9aKPG0tGYsbWQg7CsHWJDS5egzsCulTfz4L2JtNGxbX
QSgmLJfrfgy4y1S0qeskPSlAPb2/wGO9xok0ZO1mHKDBXHqWYSDtxne9IGi7PEVULqEpC5QZL3Ji
Z2jEG7WcL5lqS/9zSQ5ioxTUGfk6DArrbzI6BLsZwtFDE0F1oFPuNF4R3YmA4kUDChOlhpU4q9J0
n76qv5r5YCHqAeQPTcyuVTU5O7q1ahDsa57rYHfivBKwnnzBMswRNzzB5fHbBfc986fnly3A+FHw
05TkN8ncWHmim2S6RHUPFQ5S6WzH5hNKn3Kv4nM8GlyYPyRgYq9kmeEwdOd/4xpMI07F8xEXQLUp
m9QhMuervzmlx+66zo0Wy/sYV8HOALVYE0xoYa1X/kUANRT/LMQTYo7KCKWb2cXjLi4ZUVejaQhP
ykwanVQ99KFbGRoCDclybLmo8Oe3ByrB30YWzeO5lYHvD3UezlUQlqA6lK3ByZGFsk8MzPHvYbfk
yOEWZLGie91XQq9vwwAqUOXOC5cCyH/3Ym2EfMKRzlbp9viJxopCVRr65xIlqOAE4c/iFKW0+GsP
VTYzJaruLjDHQRNeQcp6DWum4F3z26m0RCgR4wGV2GIRGQQjI5Tr/rzWgABiR0NmqbXwEcup1E0C
eeugRpijYZir9+khl+fvl+WudXn6yPKxO67GQiw2k3ZP4PuSqsCW4mp7VzupSouPa4ps0cw8jBeT
Ewj95wLkrAlqsbBVZmsNy7kVNvKYt6hf2PGbzyBFPsrLdnTtgGWk7YSeShs6/vs9WpuC0+2YcuIM
nNTRZUlZuSglzGgm/WEYGyNVeWhTl5GziUn/e/LEIeG7fdDRFLmRtUqXor5hhBYFojOYGUlrSMK6
b2Z9j0/1ydY/oDXovXaJiJlaaYV4TxlceOQzigfdhKE4F6HVdmTqBKNY0TMbf/TZl4RSnciFUW94
b5Qb6YtItvCns//IaH5ZEXabkmCm175lt7j9V+Ae+gxkxUGEiuElIWuRWPdUVkNHHTfVNzDOqLEL
8jcivSiOJPb8khRYHwMCXCtccZ92uEiW1nZOsWe1++4sYZ1mihymU3wQ6E0wLxqFmrOegg44zFaG
QDmEw/ZVmLk8hiCMMFnbmJr1OblNuyzdqNCQ1h0NBn5GkCddwsgYzNvBjgSkFvRiQWeoe3YGqlwu
sN/BwpEr636+Qj30++AkhyAAaVyzIa672lkKbL7cAVngbCGVA7pTgU3x4KAwqNpfQDpRWFbLMJZr
Qs3e+uWA7KekOUnHhqiQdjsthfQBmO8PftxzH+Ds/6pEnGOvgi6SUCDQ4Cr8nNeLhnnH5nF7X9BP
GrHk8FJlFPRboU9+c3MgFPkpx+yv0Wy3m8P1ndBLIVcRvUzu4F3LE3BsvdrSmOgYxHd17G/JmtbH
7KXriKpc56D8/vYpKUtO9TfzOjNYnoXP1WUAZkrqsDllS/TzWh5jIIeczfQeDj2mzXWsiEVT1FpL
tltu0fXf8D3HSCdmVkcegWtB/XW8ai0rk0Q0FUXGn5XbyK7Cipkdl+VrTCRftsR9Rz2zKa79XChv
dHAERP9bAp6mvipHDyHQiiASa06CSNYY8vqv+cxIV0EMiv57a4+7kR/M7Om55+fQrsYjjgPhkeIF
9nND4LHVFtj6y0NSq/r72xVeBn+t1gFr+p1VrUytrQMbo90vLZEGjB8EUGo7xVr7t7TAQXxCMmqo
DE7Kx7FsUG0MqgR1UZzfRAZ4V8uqNyNuz/6V4a0/LRLRQQ04y+3klvU17VdKWLk0qVHeZ240K09T
hWWawQTMo64YsdNpwC3nxpO705JcCCeRNicHgkrjTSQnr8xhM8VRKWFPrqiY8+IU9w2XCd/MYuTI
iOeQCCYpuew/pFWNxna4b7gco6PrW73P5cO4m9OCZ/3sD8d3dphR5nhkIKZFF0oxxbK5Na8xK/IW
fhkHbSbZquM6gguDqE4a1Vjx2CdHamm1sh40+LPTe1084JY1Wbf2WB6s0QoGmObqVd9TdQcmELSm
NIUREktaccsGLh66m5xT596uh6wZztdxePxNcWK7AfOeeUPlgDpYfsiP8CRQkWbYiKiIxaAybDpt
yo5XMnPN61PwJ/qHq56kAyRqWx6lvjnY3OKtL0sUUT2IEGh1RNvZ2N5F619XeOFAihEvark2NT9p
4szBe7hDyJNG5FDxlfRUd+o89+rgS72OSVaHs37wVLbqZhZvoh5S8VZGUbNwb5LFRV8hjd+CYzUD
XCRsDen2rVrAd16gaRfQTRciE613l5jwEuBx/y4CrJv0QoFnfogfSrY9rNcpjn+ySqL3nsvRSedg
iW+GMzQvfrp2dmLAXOtoNMDAWG8MWK1Bup6Nyq1WAKq0Jav9C7Tzl0zNWS3DLN5ueiaYeGtyctSy
5USXI6ukARL3+/ultK/4Jwvn37AI3NUXJFQZQaoWyYGPAHrVO1t1Mx20ctGrDNEhUr+BFIwST5Yz
rBsojYeh2N2jMllJVp4GyIF8W1qddby5/zGWY4hckt546hhc7fS6HaXsiYhD2gPUbIfz0vqh7dBL
Oy4E7B8+za/ZgoBKp/J3Yl3Ixkm94SW7dA4Wk5bw2NPrXqCXOWbwmLhz83l0i8YJP3cjgCAJy6Ul
dYbxKRV+vVipN3lDq+UaO+H+Sm0muRyqgg80963YY3XDch21a9KC1j347Ci1UQLQj0+GiTzrmhFe
jdRlcC6Pa7P8NlABE4p19Dz2HJq+O6vokT6FjpkTlMqVu18xpACWe6Ndzdb1SQbcfBiO+2ZCqlUG
YeYqhUL+SDIUapNdl//Ita6uQTmQ3CZIyP9a4pnpMWfN//6Iu6QWnvySGAuiwoV0SOYXzb0b78DQ
n19blt98XpRPpIMte7IhZcpqmYbqL8RnR51530V3MUwvvBHAwTFKB8R1/E1dHSOLBUDcABYVO5GW
K335/mZZcUPJPrpon6H9xairsQcfRsdEnsCxE/HJLQka8rIDkv9BA8/0QY2+Yg1CeJfW2KMi15p9
0rULZdljIBlxhubi9WawOW6y/KnZH+ZGv56IGfo3iIRIEF4sbZ3EuTlYmUxR6CjQJBgIE0VulVR3
4aSFOsAIEtRGUxQ9ticVqfFnqIYaV10sh9mdFkFVfOSUkIXihIP7iekkFZPUkcBoIQCbOAnt+147
sAzoyBFKvkVT2U7ITXhYIko8pRaqRkdAz3hws9i095uXZy62ftLUzgh/fivb3SVPkXCPSa+bu+iN
fflHk7KMdNwq0UewP6zo2Rxmd5mhJJgbmouKGtyN5LFEI2LrBo7dl8mJb2clvQNKtbo9WNcHz3ZX
sacs+nXspKyjbcbwMEIfwyUgTlc7g7yHeGD/G1EgDlOwXO77CWMDIYKrSoXO7kvmk2HEcD64IaI/
pMFL86S4zzUNShlM2VUBUNhnHf6kuMk2bLjTIqAFCWZfcVJSTA0AfDOeCf5CBOX2z/letgQZjElQ
s0lRSR85+HRJTStpcd7S82Ufg2K9p6ZhQ2wH5h+CmX9VR2Je7FiT+o2dy5kmEWztaRJLIEHQ9y2e
EJzjEHwgngI3JfNELHTQTAACAgUlDVJre7vjUQqqBFXvJReq7r8S3UKEsTqAKNNB4E3uDG3jljti
q5cg18lX4D6hYwnKZy2ywdBPlMyLRbaXSrkmm9aAYPXWSHT9ADsQz5VSrIOuROjVxGmF/WAwhkcj
gwQxiw3sLp9GFzxP/+lRzpjs+Ngsoj0BAiVMY/LcZF3dVIJRLtg+reu4kNLGi+qUpVEftm199Zmx
XJiBRKEY4STwGWKI7LJMMO7nVZGR5eOJ7L1wUvVmP2GQUy2ZWK5SE6FzGF7ZHovQ6TQWFF+JIO0j
1enOvRqUMq+oKDatTGvk+C7i3Sltmd3aR/jWEghkzP/Ez6rQZ8i1t2JV+bNBjnjB8d5pqNIl1/j4
+gcbiaJ4vKrMFzwwf8PVDGK2O/BkHH4JvgXgNEPSbimLPvnR73EIjbCxh9cBcg3vU7/jOyj9kxw7
bj/Exg06bTuyp0W6m8seZU1bRUSdWSHruW0twsMuDxC8eLfcKZUf8L9PcwfFyHTV9HFfGdI5i68g
JjjBZrxC5ZqRjwcd5BmtMGeYC8NW8ESONP2MkDIzMX+N21QvNMnZ/7bB+hIiuu4qOkF0M53e3bvR
i1P1fJLtx/iG1/ZuU2xFav0ywKIckwBRzyrJxDvFLbOGg350EYvw70ymHBOi6h7VaELDWfIPGglP
pkROrq2PHEyB3w2pDrAVQg0gZFeK1ZQ8afgSHvgJmeaCNOArgmR42a9eogLfl0v1qe5/1hO/05w2
ra4PU7j8jXUdGv7XNMp+FY5zV7zCf3lladUq0JLfLLKuVqww2NDbLmMtipr4O3h8B65rxpEYKA6i
s02hdnCFNO1qZjo1FWzgSSk11zeIKDT0JEYIwDfrPD74KyySTukKKvuU23H6lZ2EIZFEcR3xQJxN
mksMXhyDMLo8wOn7FcfaeOTXNVPjqp7q14G2bxYzZrqtqNHa4b/OGeMUxdE6JJjfkqx9M4Qx9q7X
V6M+mTh69Q8x8X+sZY5G19NLjS1SRl5nfE5EgQ4/yzEcEkk8PN741bSd+QKY4sOvL9Hd9rxPxa4F
xL9e/kHf2baqgWQOmBhdGVEBE4F9fJ4/amAMeSsgqFFUxPU5Wvba0Epsu29//ekebo3Him4vKXQt
uFwcRi9rOew5svaoiXapsGuspe4jNZLvgbZwNngkb19QzM8MwwqWbSBkhbCKgVJ5W3O1uXv1lR7S
5YhzYZ8ta9Q32Q63V+3rcHbf0WKvE6LeytmEIfpCZmjXc2yiMVGmsFXxrJyN65EsCveC9JV4+Xe9
et+Pig8x4oY3WYFz5S/scS/rfsAS8k8jnzFt8NXnhaZGqoYk8HKgiUs2WegQsDJ5i7CQ616r59Bq
7ZiHtuJ9NXSDDU70SPE4kvWxK3hN/wFpww6Thh+K2S7rrvUHvBD5YBC0AraDx0WZmzyG7nixvKl6
OlZffb8wXnOa91XAXPKDxctUmflcRIQ/yCJMBfS2vUczvSEaMuHIOBas+fDoDRhq+kiQGunfJT+c
g4kWe3t+BWkLXdG0U3XPtEYS+846gluV6kudV/gT0ivw9WfK7YvEvbMlI/YKIRKpf0LXcEqFKJoL
FSF+klHhFhidHgxO1HjUnkcqg4fNA/Cf8Do9g7ABX8OYhUDGG3EgF17IXY8Da4K9swcAp9+iR+ng
r074a+sjFqShsXP/sAdISvEqhz4TPuJJ3CRe1UTKphU8JEsk1FWkBS4bJY/m5U4gPaPMuY05PfOV
GMXEa+HPYx5Z2cYAm2KME/2hIqUhtajLVbmDNLPHoH4SfQdLgnWBogt/L5ZgkQafxPdCeKuMVkzy
zbhiyTipb987ErQtdCEqKgZAq4qNyYZo53IAVUjrYKsob+pjVoToFsICK5HqL7swlgoNT104KlSZ
fkQkzuWZkhzplTvMTyyLTKOS1f+HR20Kh6Uivw37JnVOPJquLa5rAXw0jXUGs9e7TBA7oUSsihDT
IP5kMXBjbPeRSoWRixIghKkXVdUlJfOKXYBUcCTSkiBzJrtyYz4cMwOvHQLw9xnendNzLnhJO1U3
hlBLlERoYNXJWtAvCsrYOfanbkdGiDeD1s3h4jl/wfw5MhJu8xr/VMOw3VRH1bYTb0NI9BFpMcmj
c0Y+47f4d/9p1sC73cgmxpG7EBVbwDnnqLLbIHr/iAc2M8qRDWKA0nVZc9a4OBucAcAZ7e1s0AxO
VJLGyZr8OtM78vj6ffvsUgJ1/wRLpGBCJnm1wiWxW8HUVPOYXnhzjxKiZCZYOq7ddeb3B8acugtZ
zqeihCNR5GOJ1PcfUeoykI3KZnD000h0TNEqRyB1icts9K65SlxfjztIuH7xtjpuD0o/jwIH04eK
x4b5Z6LESzgZbHutojtIpxvpBA8i4++L7up1V4cVAjLgHo32wovdluEg7Xes9clstI54iyX1KoLj
3abD2GpTYGvouJlzOzOnWrLchzO09c/o5mD3ismto5xRAkJUXKD0+PTZwki+U5ZRWNWKsoyzA0Ue
+n9v44HrIZOkzOMjYdbnU+njC53aGaSkRpD7odJcAT8cYgVX3/MsGCpWSIG1IWnP9FifPUt5s1jF
WkJQq5T1e1sZrT71lvXvICX51XoECs71Eto7c4vIKsmg9fBi3gCwvTujeLIo/T8J8d7hK4f1PrBC
Zt2svtaBQtd2h3bIFvyCq/mrM5TT4bxeW1yceMLhebl+lXxMxYLI2FuKvZ5xm6Vp44Tqx9+DsJgV
88kkSqGbA6YESZO1/Jy7kB3rXAV4IueIgWjCWqF6EtVAguyIz58JkRurbNI8c2SjeGey/LGlDgdk
uU9/iwG2qNPIsN8L+AqlMVMy0WJAOfBc2YLWP5+m//tez4DZ0ZzOmwDCcQo9h1hXz2NDiZPTi/kq
AD4k3S5kILh/LI8QBWQWG/cql88XngCorSagjdZaqwkdzH37o3u5GRkZx9okwaHUKQukhxcJaQlV
FIhWEmjsUTG+YlmGcDFdavtbpRn11JNh8QjuVGLq2/NwknXcz2kn368BcJaxp8HHKAaLzYJd0x4h
dpM2SSsebVj5kwkHgRJgJFPs0NFu9S9JmYviBeAdUMjXurzgVIV16hPV8SXorvgT+k96bPiUboft
qBaPeeoe3Wcpz4JbCkuB4oo/658JALs7ZGBwDZtOzryjJMigtQ1sqaZRThpgRb47TP8nrh9x1sRS
bcY8OOS/yljCwT9tUPmtSmprGx4ifsQ+ws79Mcf9P2rxHaJ8PkLjGTf7LZA2IeMyAUP3yx5XAl7/
gBUpwMKDP71+XTGwX5QJhYRqp3J2pqbcxPI5S20P6eJTInQd3SPtcz0aSMGBjCsYKdhwIeBWV1GR
k8dS/HlRbmxBNfnWomUByFdRs5U/5cknDbhAfOGjdV3SgXf34tSgipsCdbed/Jatj2NSzINnz1i3
hp12yShX8C/dN+qDCswwVBAfdYJUcb8/e58ZLp8GvmmcrRsdF6HvmrUCm66yCg6S66aa8SpBI56+
RKOfpHyZeigS8/qVQEcbkII/Ab4vOfxfLNiLTmR6v5DpoJeH/RBgVYCWYPkDc3kfgFxW6AZk/2Mt
aMW40s6O8DA78MaoPOKZanmsDB69ReYRh2PXj/+mRsAAmpspYkWh1Q3qIiRVhfh6O//FN5VsXQrO
iFyS+94jrRd0Ecqf7aOTTU0rQM3Mlju6yCXSfaBytABYaZ0tiZ4v+9BA/lwxzbWuWDN0tUODmL4b
ouv2Jdzcjep30V87Xi0DkEKr+6rF+pRes8JOiYwhkREqpA2a7JqjfSJoXhjS08uqCtQ1W4Yv5hfS
dB2YMyZOE+nsdGmON1pg54jYM7ATOZsjL2orWP+HNZ4CK7KJKxsgPoD+aA5bLYHonVmr3M+w3wBN
72nWPJjbMV9Gq4QY2cSJFkX+tf51/xFLxGPpweFujbZAWzDfmn7zlFwEn1VVLbLPRdsc5dmgeMFD
yB+bHruR0iba0h3Mbolb5ZbpoxLsw4MJFNQaFoHlZLy+B2XDlEqGyuXFunceRnP8cS2ZgfCVOKDp
S8ldAYs5sfHQHk9YM8pPMQNZPIu9e1zR7OE+7XlnNoFNUiRIPCmCVisbgNZHX7txMsT2OCCyNsMq
j1vY9hstAWY7NV2pLw70CqX3GXDOknEw5UkhzsSmlop1tNeok4AD5+0dk8DyRaSe52eTOHKZxz+G
gFd7aXOH1NH1Tx8jnrn/OiVVVhnvm3r5Nh8akG11K+1qjwVpv53IaBkaYT4d2iYjL0P423xhV2PK
ogsBf0eBhQeYqmpSKd9+s+BfIPYcYMUx7+kOW/QA0j2EGVP7LmhP2DU9s8i/iHjdkmqiuqGcBz4k
/KUhk2ntSGlEv8WJKMXzTkIyblPM6ZPgyTp1YvGVIQKCsxGFFZwINclBrmOOZdd9eTSDVk1v/sPg
M7W9vKZ8CIEmji1f4XFZ2ufkxyZ3SwqlD+wn5T/tpVNm/bbA++zRfdteHeTeDtwF9oem03MmgcYL
Mm18WoebCiDVMKcGs8e36Vzepu77UWv69h2VC+yejesZ5InAavuQvBX/hpS8MdvhFh+CfhQS1JAj
zcO6IPuxSRatzJqpxS/6NYlWKaJBdh7+JBDOTK6t7pZJt3gai/gKlagTWLbLyPUTbRvxUI4sBhCE
8SZlpHGuJW8QpVoP/s3HizJblyMdAyvW3uYy5TwRuZdQOqgQttrzgkzwBPSeO0ausCUnZ4gH2iAD
DxEASAQ7IQgK7IYvUaA9jy3ENS1tXhU7oKsHhckBYt+hjWJ8TPMvMd5OPAeiD6OEz2VPSbl+lL2V
OO0n7fcom9frTAMhjuB96BuTM810Yy9H5yTPqHW0zvo5KJsMVYZZFaqgUcDpbv1tLqZyPQP3GLYU
gJ6eftY+ZgYtAPg4VTyMEsxP/rtrhOSg2iJoK8qfRikT5A7ae9aGKDLKHlv3gnfWqCM1U2g9vqNC
FSmqGrUs5cfP0I/M1FSGPYbXYEPw6Xdru04Tr3JL8XdWPHyB+DnKev8rouctcUUnUdV1FI/KQLkR
jEhCB79KVOuhF9QzsoJoT1G0a6tYe7OCbXbbgCQgM/FIniOIEiSvQKM7TUSg0YNVMmvl+DWiorNz
AQM2fM1AWJLGPlYhSix/FMxXEh3n2rP/V3hTTYVCoAeT0cockHfdXuqDNfcVQIemMmWrzTmAEeHV
svk/OGHqbCsI3jwQc8g9vWkJYZaDRMHmPL3eNsVkZNp+U595XUJkYBJBPE0HQ0fJWmjLlY53jRCp
AlXzr6K2DIV7p+BHJHL0TeJ2F4GlxIcPFUttF2RvwkC78atbvS+fgRblulo8zwrsIq5yi9bjg08J
YVkEXTWuBnuF/67/vpzC6WXpj+lqPvFVKO+TRPvGnHr+icJbo7vNDmZLKaSfu4PLnlXIWC72Se8O
P6q/ayucSGuTFQ39U3qk9rcUHAIQ3mKtML7XpQlJ0pU4Aiw/E6pOyapDyjHMKAnY+tcO+lvdKF7X
f21TLmEtTGG91iCKb6YOqBrXITkGp+mZiB7BnLS14ifWriXZFzL35XWNEOZ6xsLbS+/FxavPjMmW
TXWvTeSnNugCrDLUPY+sMLylky1JEBwDDqI0bH2H/wtiI5rF058izClKryJzs6cK5sau7Lz3JGda
1YVodpMwlGI5ZjyTnIc2Gc1ScUz4+dARfEo4vM1Z3udOBwp/COhqlYW5G6Ot/LnHTaUNi7+QcIoW
B/ne4eD79RLGqopJbJk1a1qtiWKNUbyCzmDZh5BZbxllWkbO4Gghrjz/HfS9x3TSipDQT9TDJdN0
Iw7RXRwr72UpMnWJ8XD0qhQ89JLh3wEK5fAwuZwZ30M7ifQRXbMSGXtX4NGJQk65BikE3yjRiBcp
h90/zDprZTrhOvprksbXyTj5nVWR7Sn6ZxjOW35fB8h+BmyyaRBns82subTwExt712OGI/lftlNS
e62uirXDX5WcdopxZMWu6ZpSxm1ZGyq6iQftzbLbsI6Sw6YO5cHHzDvo5Ufy5qR7vA8a/Ewg4hdr
5uwWdqijUzVSqBgg8hVcxSNWw1afQVTnTnkdSCOrOrC94Ck4neZwIYSfp15kl6+WDBG8SyTdBelD
D08K8HwXzGAz5Q8dqfy/dPdKuIAXccerf6g99d8UVDtdlfgQCrrJWxyV5tEcGDFj0GSX5syVf0J/
A84QEjn9FRHV6tPx1BtT5TcE/Q5mBRdpCb+gCxHY0ErqyFChDiwlqxB4KeDhM+n5Wa4dKO7lWf1Y
Wax1FjYXNYr0/0q/CxXaCYoBouu7pyei1d4IwwD0UYvUx+flCG8Xf4GNlyT7CoeTmz3P59PesfSx
SHRp4I0NiAMTR7Jj+DVgH6euAy5M1Hp/4CiNCj/0CnHlPARvmRr4+GohZQnB2RbM0fAb2Qa4qnVE
fXV1afP2i0vAtgbNKy3befyoB8L4JYnb3e0WACZN07aEoStQyl2+87Cp1UoMPFmyrQqGM//X+pI4
uahqUSgkCQDeuC+idvHKylpsB7K7sIc+MrA3vH8PEs/twaDuZ/DScyxw/hYFjh1k+L4XylcJ/8L6
ASZOIp8wHt3GC7tsSFa4PClptbLQx62iNnh3idF61kG09mxO8LHI7wUopYydC0zWBWb04hHMzNn6
XCVvVX6EriIZFreaq+oqh80dy2UaWIptLakUsuxW0t/YRXBaZENfjunhwuzHCSvNRLAJdin1HeD7
ll6x0az8PTLcFZsTAqvdRBjnYcJE9VtL8p7R6uYnHVzt7IKpilmNPk/Bom8LyUWR3nXUQugETmIE
sbDi8BB4aQPl7fNsFoN/CpZXzhr5fcdkBhjhbApI14LyPtoN8bmr49ESrgPxLybujoqOicPhRpE/
CfCkysPCnBLUjN0GGz/Isf0vf6y/pkKJ0ZEG8Se82f8ku9vYOlJHVhBbmAhupEOIh3yDnXePHRBd
0Y9drMYQan0LGrkokvEawHUKsxgETEmIWKRHMihO9JdUVOdbVMeDLW4FU2YFMWqBicnu99LPvCiw
3Q/wYmpnf2BcvbMXqIB284GfZmVX6aqnnlFVKy4v5eGou0b7u109c+cfiRVKCq3t8/R/2onmW0rK
zj6M65MEzm8bNNJaQ6Iu42hwu+yEEz1qCjf8y+GD6kn/7LpkFZFFQ69O8sKS6Upd0rv9DGmdImgI
1+bOeOEcMX6XIrQe/zp+hNbOT7JIna8bnddthqZtHeoZbkbevkEl8AtsNlrvJIxucLlXRphF5819
qqJJHmgIRUCgaw7Hf0yiYTDCDfzxqHwKYxnMkkKNP5p2T+iVgcXhzS7N9oai2VgQQH9DIyy0NkrJ
LQuYVDHgQt+PN1iGWIAeEVC8UTnCgG2mM4s0sjSp1uY06Qcqdre22CHUDmHeOlsl24WQqVoMCU3L
9uWOWEvJoGTZsL6KXPd5MqkiBabeiYLAuI7gXNQc7ldTFBW9TGSU3WWH722ocQetKEJnBwG0awEq
PRkeAuvE4eQXc1nJjJUK1bwZ0K59SV9rxsc+Ags08JWDtiyEyp7D1xzI/IF6IaGdCUetNqsauiy6
L82R+43pZUGmJ3Gr645vExbPiKQv7jWccfx//0fR5cENLkW5vqm1os6+D0PdSdxOM2MpW/CtjtII
IsStauwKj5hcySYSJTz5T5c8BXXVbcMZaA+UAXvanjFqAbVoTY0sNVPx3OqtQ41OA4qNSn6G0hUv
UVbpIGZpdkfuBab53f+orhxz/HABZj9yTgWciOY7kWrcbG/pWv4fXOqidfYtn76Lhf6HU7Q5+qK6
fjD+p4STH4pMsCyqsffxH9ihNjgQYMiqcMMQ+B2D9pPjENwlmDvFj2e+zBwyerFBLtbnOUUkcjQv
C4rfMUxYWMVQvb+EHDFAG1bRQeGW9EUWLPOHGWp3raB6tyim6/7c1krSLmy/3DXRBEy87cg/AlY0
W+ZialoGdaZm0uTCMUQIl8yMV0YWs/tKTcaP7D4olj+PFl57FFZmQvEHFP+BGo7g0/ayLHF/P2cK
+PMrQ0P+hQmSknIylJxeRL/2Z44Xqh02NWyfkN+TAwTe6q+Gup7NuU+99UHUWz7E8fmVNcM02KBg
GsrSljEutrC3yCcuPcPMlyakmj30UICq2KIxfP/l+/0NNaRdjRu3d/Fo2A6kHfRY1nSgYsgc/5Z8
oUmn8ETIENoidhBytZPEbyAgemdW65as/YsmujQojVu56s6hKx1JMq2EO/P7Mxfgi1eq4+86SOXm
yS1kJwKI+ubkddy/iL3tkgsP/SXDWFJR08NMddCWnmX+olNVgzb41q645epoKquRaI5gTpSgExKt
Le8Im8C2sMZobvGZAtDZrIqDns0eWo17MkJHW+yVlTBk4Elcl1eLBVs/ImuUCeU6wVLaPbMxLo52
tW3gyQgF7+iahnDb8eJTFhum0ZSo3RkgrHuIsHM8wgwRCvKkhJ7wRSAiEYU8kCJmhz0jSk/2See3
Awit6NfvM3HVnt2I/rni5BW9WhYbouCJ8iV6mb20KZzjbG7PZdM5EkNcN7mQKMwSdOmy2YwiqRQm
iBQCOGDBxWVRJKRm0zgs+/N5x4Vt3F/kbuHyr3FAv99N3rDxtYtRfBsCjAVTuKA4FBWqtpglrUWz
W5jZ47eTB8LELnIgiABJSA6TPeNYzeYVbrI+ONlVLXXkkOcrLpG7qfh7Y4/BrAhpum0dY4+F3RRT
rAkTqa/4tvlM6yhnlV1vHk3GaGO0OkVLUxZXHnRFIM/NpoyKnTsFX/wGa2XLuHzmXXxOzUFi6Jph
9n4iT7viXMT3zb51gpyKkTE1Z2w+zgU/l/b6sKLZjPfS48IeWkC8ijbKZiSJCEYDek1gP7nLhHp6
0lOZog4fAXiE4VZNhSPH0El1vUiinUuuXoDJXLK1skpZlsLZCkhacBjMCAt5Px0L+Z36cypXH+oT
dhI4AjFi8NfmC6ez8VdiY3wmtwseGl9urJ+u83R3PdKYrNAZMykpFHzu3t/wlw57q8/oYO3rX2uU
1ES+9vlk2aLYxFdZq5l7KIEsrVm8TEmoRdxvfL1qlX6RWE9h6P9n9CPPW+hxhOUI8gr4F2nbvEYU
E9xwZ3T8QyUoE07R9jEAw1hTSh8Pigru/X317lKfD2K0pwRLgo9cPgzvv8tSJjpceQDLwzFraT2M
MEzrJkDiK7i+e2bZLBliKyJOLVHwKUimg+sa6E91YwDZdsv55WPa4boGEIuWYjKMx87MrMUq3X/t
bEFwHL/G9EkxRsgJ2Z/tNSt5jcMPKD5g9eaS+qGy4iiygAQJU2D2oJiRHnKqAu6a3I3t/c8j3XJM
BWXXSJ8NQ7S6vZqNZlBMS4dr/pJBtUIkw9JxrKsHRSxiDJOfa2ZzWp9BFp8mFC+QXG6Hi+9Lbl9Y
c318Ua/cOY2Xgyf+/onBBtDdXlzUS2SkRvmwglLwUVfYrgfzZfqG/ZhLiazwZ1oNdG6vcjkjsisp
qOves3DK3Dqh23Kt3WIBsoviXG9Q1nNwgslneGAzz0BTdSe+sl+QuSCtpHXdPYbwZs1JYwmKqFXF
5QZCioUQmLARXu2jTisrJKGN5AmdRZgKEpNhqMXks76sStQ5EcD8w66we25fHZVaSzgHagYmfSJQ
FURsKt1luR5abXYH/53UIbtRxjY0ZYFJCfkcgeelPJ3zczNcT9/cI9PCKfScsVFNh8Azmgcto3xM
aiu5WwreGaDhol+DRJ9ZdVxTSAx1RG1wnDNswSYPt1Mv2vX3y55VvBNDwGKc8bAnTpPqNgUEXcdn
NghyOYIy+rKG8yMs+XEa4fhJ9dMmBx25J0m0w9wZsqsf96OcbIjX7Nc4xXaOj5+y11+euNsHKmUS
cpjnmeIiRnq43thv7mfI4WJP400CNxoZscSSt8EH5nGIzt45Xd4PAruEZxjq5hQ33+V8atT6TC7G
1bprNto8Fh7/4hIbTZ6HSggk7CWjXwpK03o6TZJBSJtLL54fTvOZ3VgAO9arY+ZZyNzv1+gZcUO+
s5M9zAvXXaGQbMO3HEFgBRfYPFs19OjUpyJfYO9zWb0L+iAg364YKnr+0g0RLJyRoSZNqDfVcymZ
PrzpRnqaPKCDk+/m6z6UJ0vkFF5j3OKCnfDMN8HDKCyVsHUNPYqnbxKBqxVhP7PUgGt3XcghkBSn
pFb08SIhlqbqUUrW+u2qPc6o0dbUR4be1yfUgGcr9A3P9KFjAtYds6z+Cv0Xq98x2i7sUhVjW3XC
Mynadvy53d76pKuQ9d6LM8ztGslFGWyTJ4y/w0zP/0IHKng2vlMhlZBpYLqFQV3aHa6S+gFKggvf
yoDvEnuSDIfKF/CHg7/2llc3rxNOY+/4C5X9/FsTOlh9Isxvvlb5ekjz63UptyhE/Az5EfhHbRdv
Df/ik9TwvYoTAg/Lr4L5umPyNBEDrWy6ws1D+3+0QtwR4QTVj95U1eAo8eJy9EEnIfw3dawgvvOL
qOumZSVV5cC78co1ipkCLYkHl+SI87kWaTk68wnqs1w2J66+ftsJcZAtk4Ci4vmrKVt3RwcHODCo
1fECouF/udBvCR4W0XB0BhfE6aOZcfpsCR9inTPHvA8pX3nb8OKPpt/ZXjKx088gE8ysDTM1mHKb
CjKx9ffg0z39GYmWOFaWennQPilp0fW33+5SNXvahQXYMI+ybqEJfyqL6acTYyaGJTA5kpZdOJAJ
UbGFvLoihke7k1WypAeAe5KNd1rh89oKtk9MDF1XJ3zQhzI6YRPpNJJYpWwHer1e3fpaoWpfTk/t
HUOwgEw37jpX/GQWfidceVQSci523OArA4l5w7tH4Y2mR3Zts+oObHro70HT/4LlMhYwBrpr/nzW
kIEUT0sZjz3uQmbKrk7ivF+aEIIzIpyTvzKj4bKPH7o+FnrYbHZ4os9786capX/boJ+Ozjnjg3PO
cMow2xzpvQ4BEzsH9P8xGURpADWkEgpVMo+lY+WsPU2rRv2dbmj4fr+ZOvdA8jj1yZbSQ9h5JxPv
aLHuEjhe/HE8ddeoW94AJoS1x0TfQdMMSuwCHf1kk3s9nyRrfgD2R5Wqug6GfCQJy3Z7+uUdP34N
N2FTVK5e+lQiiXUgwoHen496jF51lJmztsG9hkJPBIwyoQT6DUEBM6LpI0ysJERadc5Yq9hjQ3AQ
m1O6SEasZ8jQrVqzL2xJNabRdYRc4EiGRf5tkOFIZa75MznhHBBte8enM7WiALl8+mhqIynmNiFg
EToulrI6qg82z0Wwl3dN8t+2xOBFs6Kcl+USsyA8eMqw3V1Qn9hf4j2wAv4k2lPj3sm4Us83Ee5r
sikQBwWetQ/MC2b+uEVhdJM5V/HRiM7L59zzi8b+jht8Tgfy61PLj8NhaEyGOfTBT1AFyFXXIcW1
5vr3hNlAkRiglKrbiV2SNepQJ/O2vjzJkoNOj0CJADHMHd+78mLDTGBuJPx9P30dAi+o9bkgsrHo
eb5oONRmG1UsLN/8pqNX14Iipqil5QYKsQxCDbfzFBYp572suXfUurMcXXIf3kfKcIoyhqve7ViC
Ax4JDZHKGsBmRLnLVhjA6igfloup3YSqziJiD1DV2m3tiNtoJUObT8vP2jbcvtMV3Yjc52lkjHf1
BweOFzkpdqtWPJVcyME7KrBY1C9w+TDZRVAJf3BSy3FBtLFJLRAUYxj2tJYvJPFBWWg7BI7MYD0F
ZQanumYCML7pYebocGgF/BPJpMYYlTi5CSLMfiiGLOlxf8IQgd2ADO0wpL5nGlSfThf5LVCdVE74
hM3CPC2Dl9qHbA8JL+1zpOI6Oh2PxlPlJsVn/Nm6eGqTUIlM20g1U0YywMiN4sego5jdzRw3jfIY
evV3wXn+6v5kcBD4P38yLyLdjzBosPzA/bPahY3/Dk65NK0ccy/5TTnp2lTGuq4DBq9GRuHnInBm
tazgf9yu+20LyhoVZ/z1CDzlivKWK/8n/+JOgL0aGSX1wQrbwtwkRmqzG4UgTfQBoxDb3TDJurni
HJM6+d3QRz8CUUHm2s/uC5ETgrmGP2X5eJKCoie9cRDxu47rODwO5gC8CZZRq3zlBHkie6Z3eMZs
YfkRsaFh4rKWbU95gQx+YK+Qo1IHpCtmIogomEihnqmFu3ONnrtKRsyAfF7JIAVK9f3rcWa1SjBb
Nj39kbDxBFemajB3NzjBm5JtY9/Ss6U6I560lxp5Dj6B15qJ5EYrlgbAH5wwjlHH1gEWGrjzYafC
mhFZLV2QvdfklGUaNBqFnijQ4qHHt0PPQ8pUf54ijZxv0aDnogDmJVdHtbq3xuGEZeA8voxAELLm
J5Pw8jYCqb1H5ETuosvX/w9OXZ7UcZO1/JiXX6esOoUmY3qMU1fxs/48s9kHnIoSI4Mrh4r1kFtC
ZvY4klCPyJyE4YC54OsihbJhRIIA8kJOmP0+O1DfkGSvX/shWph+bfULX4Edg2ILgaeoXU7mEZYr
/WheNGR0bhhLFL5G7SjeMicH+YQijh2aEw5dsy8By5gNv9UKKu26OH0uWjTh49fMoWMNs1eRQXiF
t8xqoEnSnTcbYn06fE5uu72oX4CV+0VQ9GKiNEBHn0XWnm1qe80eNy0ZHBP0PDJQYuCUcRWZxyok
ETZX45xMm8qQy/6e+0u/66rDWom9G/ZLpGrgP9L4OHoAFSmZpdtOH2Vi8RQeV1fX+DGp27fqgu8d
r70vx5a/IrlMHVWW4Hdq60WuT3NfqcGggj3nY2/5qhDDtEQ7m6QKn7GdwX3RdS9KT9/ItYZwSsGa
B7XjmXHt8KpYwmtuJKcacGcBOcELsc4mhMcvZXxstAak+HyKN7CwM7Q3KzSp+v4v79Q5ItUhgo6S
BQZW+5HYt6BimravMz9FQonnX1DKeMs5j805I3BAIUOgD2N5jyMKbx4L+5heQnmL+h6si4HNUoSt
Ope2h/NGJz6dmrXnAoh+oYvyzdxsE+m8kOqTsKWyW2kVoj0I/Fvwj7yGJQDR9mW1kzchsEc1+eSt
tqrdHUKxKbWxfxycV9ltN5n1yg/S/JtbSfp/I6yPkmvxnJAjZJUJjigISPMSCaNaoMea3ZbCZIbi
dgMPr6DhTQmP3DAS+NWvKNVE/UaBwpdRoSRtSDZ+l7j7vYxHk64a/MNNnD2aaPKqcVWAe19jWzbo
cvno6ep1wuKUR4eZ5RQ6Bz9GOB/T7TvkLAusH+Ii1NJCIP7dfgGFuliDlqRVgh8No5ym4SWneAYa
rAQKSTJAZEKZ5V+MFdQLHG0EPMFx+2/tiB0hfZGqww0SzTIUx1d/mxL2fpqNS3+v+nCJ/RY00XNh
Ud05k8WAIwOi5KJgh0IM/uuyi29qiua4HB6IBgGiUqZyROe2+56mmXn2MhCbtD4JQ2yQxO0lw6Qs
TD6yxeiFQGxemiknm1r7w69dL2h8A+t4rMNpdYjgOL1tIrVAVrm0GZYO/iI3Lhx/OxhqLoAmpQGo
XIHbvA6TOZIuN8QuowXMeckw1Sm+j12oXeRmaC8Y92TH/bUBkvw/yun3gYWpcnuAJpbndeA1Y3B0
Ihrrd+aRx5KtjehmQdEoolDDa1yKmd7wj+UGLqfX6l/coOuhdcwYVQpPbS8XDrZYnGd+eiQjNcGh
JyZpF7j9cfrM59HXAQzMFrS6aoigcYFsiFGAkjAHjKdqXL876YM7mA+4LDXYwipmkFyVRMFJ+iW1
Wwf1prGIwLI+Hj8vJs3XApgVHNDfpxJlgnbDn1fctiu7TrfCAKhnsIRg/qgRHCRpYoY5IDJ+9DO8
/Tyf2vT9BLUdOWCaNnu7lpOqNWu/hik9mGr9P+KLdpSzHC8gl/ckXtPybTqVrH0hGXMrLqLJ4VHn
aQBGH2lIaAM1B9T0BfZd6cbCswQLBzrN5RJITrjz1FjppLb7VdLwwZGc5U4aAYVq5D1XaMFmXEwF
0BH/YBr66cRgLFVKIV9aOW7utP8bOWxkUEMhNyKWFH7TwumZGPkVb5ksbg2LXSzHIqJ3Vhmd6jk+
nsMlBOdfP6Ga9Ve8jFm7CPHD6w8ijbZ1GXIR8XLnYBl6/ob1ALSeBEmjowweYq0OAroVidhpRtjP
M/QLC6t0yznmi4IcHTxJ2E4sj1yNPXrlEwmVRSfMrctgWYZMlRt8Cp9Z92juDUtcPMV+tiDfOATK
BYA/9ci3v2R+plT0q93xKiAo0Qt7FZKrttKtrDA+j0z/J0wrsj1dwlB1hA3m9ade+dcnicKYmom6
OJWMB++CSYTPtZDopn1pbgqSzv85KiFTDaEIN1k4Qv7OrC0vmxf8bS6Xvy/DK3HHWInqdEvWeZcY
IaFvwmYnllQMYunDqY04Vh9xKnlB/oIu5yb+6LnVyokKzC0ZP+vNMc2WszybUtNlykfmex9boZtz
Ns8/Ahag+Auenuyjp7IBoyDz3Fl0oEqRB0lDyRRJLMccqxiIxH588xwvUza6cEINWxlA0R0iO+zf
DL51gGE6w2qlSCktcGbShHGw5DeOUBGqXi8o0p5Z1ogvtVWtMUudLEK56hcRgp+CB3GdrJt/9uk+
NuzynenTwcD2WjVAniQGft/d+tRN2aGgYJn++NctwnwTR0GkZp4YPgdzGPU2V17tIG0OWUqWa4Nj
cREenUq8dMKnJqnAaXMx2ysWsbIZfCKA90UNek5u+b9CoXrqcPk+dJzg9BUMJQqzIjM+J6LSSiJV
U9/CaqkZ0y79R2DtQaVtKUosUypuMYeptZloRZSS01jERFF3nVr3vdmrajVkS/h5lK3HHrxKtAAF
0HhMxzDhxS+C8blVIfrc0f2eIGJaXqo2j6awmMtKW7UtKg2CIHL/dJ7LhrgDWoQP678loAy7PU2y
Li3Z7k90rXwmlN2mzvzMggQ06XCffBH0AdRYTYsVqEy6zrSxLkH0r2agBa7t4/W5qPZe9YPMyMB1
laDbLXiskQO2awO2XO/Nyv1dJnZEg+Br8NS44jeEFCWflgOTb+XUSZg27T34Z/fc375pDPt8sYbo
Mk/qAufJyUAt07nueYpojgtCnhh/CLiOI3bTBbLuBbCwXVbMIXrgryIlWilLYYHLGp9DVxLOW5pc
Q5rld2mXWPLDKUAb/ZZ8qCOqFIerRI9mb0OjKs0mWXUO5v9MGvRZ1ggUvt9aBi3aZFzNIfqJgj46
D1zvNjp8WikYOQZNpBfFkQddm8oe76OOOIlcEfMTumfYFzDIhPFngytBtmO0YjNvC6274h1A9Kte
ZX6fARn8B4FDojqXiiLaTwrjVtM0I68Soc7HKIwUskhnk2bu2EmBP1dtVnuQGow3Ybrr85kDo5ZH
9L6aDXCj8e5V0LPiZfVFfY0MmdzXckvG5tPxUhUt/Fih3wjuef8I9IV2M3UHjAjJaGByEKLJoJdZ
+m2u/fqqkBVhYcsX4sZsxIzgbdEbBNDz05Q8a605cOu3op3pH0UD7Jp6bmygZvQzn1yUmCgyTvYk
Qxyzp5KdxFfKVzoRuWc74q0UlPLZjpXUFdD7w7ctvJOm95YzAPcq247MBOpTW/rf3ypGi1wYS6jW
3HNDHqRGEhC2GVFveZhjVew5TsHBi/z/QnY88Z/GLqyXiiFFHWQv+E+7zpQ+tdwYe2ScKzTHGeVa
sX0xNHAOMwsG1TCLwQBi2WfYiQvgs14zkW8jY1cujyuzXogVbrEZ3eY04KXDTiJOQmjK6xQjMTTY
aPgYWYszZdtzDYjkCIEJ/BV4FOJt/rvOVHapNQglp6umIoqp+i86rwlXeBoMkDkKpyfYdncrEAD7
b2zCRfvWVEhd16sFaWMsq8MQoKtuBIuRLNtp2tn3U2KYbU/1Ca9J0hNTVGvQj8HL16YLLCKxyDsh
I4RkWDeL8Rf9LXeYKX59c5tTzTKkxQ2j1Gtgl1KcYNwSlKl60xjxSqNM/9rrc+dKHu3xDeNxrS+k
uj1hj6ndIUBgM5voNP5YiwCDmm1jhvXbC2UIYBa0cKfmzA+5fvt+1OGGitmNTvfPTYwd0ewuHhEb
4svLlXTCDN/mAw3tDFjHVroZo+y+6poRrf4kBR4fxFyUavrRWOYuc2IIUXqMZ5XzJG/qvq8yPHUN
/j1l6Y+Nmq+0sjpHsT1FRGdzRpsbYcY6KlhPwGZfhFLN0NckwFJusajoK3HGdFE5fHdwqSw0BUyr
CGCjOWh+kiMx97ZGSSApNxYK1W11u6YWsYd016Sw8DrX/ObKiOPt/ySnkvngI74BnotikXJxr9jS
tHrqx+9N6pXxBV29vl4K3m6whYJba4PvbtJNst7OJtpxw7sxcIvwX2f9MoeU0PJDMWStREvNxdHW
VG0/TObbgccvUvqfoO5rvmLyzrRIUW3B1LX1brOHOuUbPAFMCLR8qL3K74+utPSrkEhfRDrDKbvT
LT6W5nfErDSXqFj5QAz0tY73jwpIEPcapI3oH9v3k3eysIWWFFWVlqKncJM3uCngB5eU1X81ONSf
lRSMNqWjJK8BLkY1fX8tiInh9fk9hmxbkIXAgoKvX/ymSWUnHAZHSbJuepOBN3/EqqAZjuYIVwKg
LTwUmiDp0h70ilgxQQ7M8vigej+PMbGdjubWBfVFuxLaq++7ooeHEDz3uGYB7znygTbqx7lK37UQ
BNfJablBT8PkQRtBCCFdEsnvjFlBl3/ZlyyIVBQeX35Hu1gIlmB4Eb0/aEK0vfI5ZFsHgb9Z4dUB
+VUGbVejtjNG58ccSh+23nIEHoDv33H8v18glm/hq+3Tkbf6uTY4fFdh5lwCvuCINmC/kWhd6kXv
8HBhN1B5Z1XTIg3PjOtC1yg0O1sOZGZ8rT1P1PxkTEhC3UcZ4t1qrlTvfkvi/Gs5S0EKk9Irg01M
4smJ88iUh8PSniMjZSOQK4lYiPlRFe6gWEcH6fS8WLGLEx3tHmYW2sO4vowOerBFcTyMAAkUxil7
HbrQSPKTlmSa8+wow1cXTBqseiCJzDsegERAVT9vgh6mP7eSvfKSX1dziNV2zsp00JvJgpilBBGC
MfOZukD0e682GWo6iZDlPlJzVBc2Ui7+t9p6MYmW7vRgeCTqh0vI3rENz+Fy7jm0clIoyz1K7plH
1xMie1NT/cd2PD6P19bsexhonhG/By/m/d71CNrWd7hch2PXrNsIy4t7gfY8x2bFj9rM28efNBPe
Ua2QCKNs4s6krAUPPa9WGushdA/zF/M4ogsQ0tyRyADz7zW/D2m1qsiiN7RlYw+cMJWVkGbu2Pgm
lzzELwU651s+Wo+nOS3ecy8iFx1WEuSoutJ5/3lQU1cdGUmA6HRAM/KfgkWiCEaOh8RnD0fLy0r4
JVdRk0EOftCFqmuwkz0+AD20jGqwyHEjt4tF/Sy27FtplDBOV0FoZ59/IZoi/KicyqATkKZcE1yu
O+CMLQWDq6/cAxV2C9d28m5hyH0RfzRM8xH8SZfZv+H3puJ9RDUBg1JQTb1KipA+wkA8Cqfs0si1
BORVRb8Ec+3OargPGMvvim8QOE/GSY2efxnmXsqdkWcuyGnBmkdcvEiqHaChZ1eQMScihIag4P+F
PNvVYMQAsiD8VbU5OExSIY9OgZJ9048ytDRQRbnNJ3vCaKWGPFsE0NTXwH1IDTGMAU0JiOxXiDZb
EED3ACer7KvUFIL4JHkBHfjnWNBNqVRmc06PGsHfro+c8xcGSkpinATR06JDj7ag84fwWFG1tSRU
Ci0B6YwTMld8nyL4Mo0EwYi8JoHT58ERTgGRr7H6hHIpKekGdsD/NN23NZKhQnHLe4n3e9kEoToy
LzEU1Q81Dr5sxrXNkdpPbs5XJwzwqUT8ephhMWbnCt+f0EzKHgQlVC5Fd219qgCDukzSUv3ghWbH
gS2Y7V49SwPS6bIjOU/+yKkf5mYETTaNAX80qrCU9CviYXpj1a5pJQI5T6eBcHyCzr/bC3oSRviq
fVlIoATP2MfmYPpnFPZ+n4kOcUE/SAFpmwzuBY+vzd47SRBhRfk5/9zg9S8hJfx65BmIMrEY8H+4
+rxKsk4Cz2tPb1fpyMZoJzqAOjCxAlQ1BM5fc/dDDvbaddzOB945LHP1F46ffkR29xk+4qv/cpVK
o9Ylw+qZFproHxnz2LPUVeANfHclbPC/DerEmnmFP2EQh40MjIi7+D/Hj5RJu8VDFIg7Q+PoW7ox
9GLcuz5dl5+ITEfeYOOqTYl2OuVnUBw9GL8c9IqzzYzcSaX8+eoDpHqf5UXOvGaEU4gBzmIVBNWj
4xzODcBiAnT7hG+olEyHiOtYLLa8mYVuCGOHayO/3EGu7ygDp8Ws23SGgXz7fFjo6SV/aUdLuTXI
vLpGD20DsDneQIxDJUE0xSzgvVMSZiEFh/7EI84llz17/J2Bq98+YrXo9xvc0wsreME/nMxpVHQz
WayUbZQTUpPCqGzexEE0J4JBD9sd79lB1pqWeNnEqcwDcylsqQLi9dAA5F2hDV+HoVW85tLViQUj
321VuG0NObncwEUpXz0NhS8zUEtbUDRZ8bmi6Sg1BjTu2IXbCVrFgdpOgyH0dK8OXnsBnV1E4Pzv
V13DR7xpFfXkoFlSwsv3EABD1L6VoBB/uSYaTVCBOu/7Ze4Fdsg61Ugg3Jm069gqlUPo8CBPbMMu
yjd4t6qSRq1D8Mc2ECa7mi5jm3tXGq3Uhn9GpqDoDAmG3xWFbRLBFaiGT6JqPIBvh+lMvT9b3t2V
IZhMzSpzXnlcd3u6BJm2ejDQupLU6LA8KYowMCNexbIwz97gd/NxmOWMabx1ZfOwKFcfxSK+8HFA
Cwo9ha9zlzvLqh6ZDgA4Z5jjCbDXZ+aWzeK9hMEf2ur4dFLQ2/XG5pBVSey4+yS490mc7/WRZgih
Jh5auQua3Nt2ny9SsvfvIhMVopqRHm/T5q/eKhl8iA/+nKwpMkS2MirfI5spJCaROUPjasU0h3TM
EySARNGdJIMKQO7szSMdcyPcNlfdW97YpInsg7qBe28dueCpy4Ls55DhgLAhax2YJAJNqiBjspgA
RPBSxiBololCP8wnVvzc888bgoq6MxqoFkEdBCbqJOuSXjeq9Ka0BzHmzskbxm1kzvBpRXFOqSAp
kJru5RuEaMJ08Z//8nmlM4zjqV4WzHzWTkVk6vt0lg30xbY5czGdlkLg7gwRGCTrEQQJAjKOUmhH
eLVah+K+fd5ucCdvBbMtSufEC+pFjw7D10qQkjBau5CMIArK9kdn0DjvkMYVBMrclP8z6rWPflAw
eGY8MDsIeH+E8mnWAsbjB1Z+tjAz6iFRES4tHrmunip1NRo1xFnJ8wEv8Gd3bxW+es7qVfsS938s
tKjCMRii8vQZYGla0W2UVY7A7hwLws6fdVMP6ID/bg2zrmrXyk1au6SHXiraZ0zkW1fCj7eexa/S
ND2FM1xf/tpKl3Y3uEM7XaD410XoXnqZjDALeqjr0y2zfh/jVAH8SIgOHt04o5ShtdTZNCFB9aeR
4RNFzh3Cvf+KxH82QSehrKzmwXwMeOZBjaq9pNBS/hmxQyD/ZMP0KyFfnGGE1DGQX1/4ygiDU/An
VsiiUClQTn28XRx4cL9dlcwJV0fJdtuuXpDS7TwzE8z3KiYcuxT6U4tujfzMkwxHuwvdcL0K6xIl
rT3RvWW+JBS7F4xg3o7q3XSqjyYZ8+CAEZxlcgm+iu4Kp7XpGZVomc1py8e5np/NoOkyCMMacSdR
GqmECuq5LQYP2eZ0dEsX1QbciXHtqSzIzQwDXLG+OsAyQeEXOp8B8gKknD/q8xvOR6m/11Zn1QXJ
aD+LSJ9wSeLHquoc+Z+RtQ0q+LWNzJ1MlXIo+hB5HtS/hpFB9bAo9mChiQ6HDUSDSwMk3POfyX0Z
n70Isowl09ng+rAK0sMybrPZAz4W6ZGJHI8hJd7x5c4HxzxQP0UZ8OIO2RHtqSyCLlVkg0JNDEFo
4iHfrpSYbCGaTF4+x3lufCL1H5g4jgzSEM/qcviGO215FXd6q4ZOn+JrVsRskNQbywM/Askv49iL
14GpxaA4VD4syxd0N5dJ7RU3WKxq8C/LCKZCgXores//bsxYVdBihQvO9TBNXXFlIAs+t/gqYjQt
Frpr8c+itIauQKAVOHrz6+IOQaaLDnqFzppnhncPM+alTmpc0R8S6e598T5qGP4S/0ZIAmTenM9U
bJnXb8Nl6Bxwtu6zAqgYQk2HXfH28ibLaUsYblCFaNj4xPal99uB6k24TbTspbFVYDhgIUooJwe6
kFXcxe1yVO1RZgd+BRuaiyQP1bTr79mQoMRiwnNpZBA+GzbvRPxFggOKr0v22jbZYGhp4zSmo8K6
tRASHDQI131Ggr3K4R261m28SBDjKyeGLTtzhmfCL77BgFotnD9qTJv1gyf0f+5RGAwVlRt88vDo
HD38EylilJEp6joGv536NNp8bbHpJzWV/f4PN1zf7etFvl1TBc5WteNPkL5XtbwIGq/BZYav9XBN
A0GUCwIphFgcCauLNBYeUfqxyDugwXy6zJCoQ2szNwsfcT2X1Yn/j7B0rlEd/2V/Wtxmw3qr9W13
ogrNFlp+FAlw+FLRKiOCqJRCX1uUclzGaMhmTxSxHb6/pThlSP5eQdgAHtDOKGrzcvTlxh42340k
T5F+2pWZbp9ukxl8jl9237GXs41I/I+3Dx+TzL4k/bVLdZcThlTLDIkoxzklXoQNgW4fxi+dWdZ5
2HySAXp7aWkWZ2rfzsJcGeNzbgjIj1Xyfsg7CWmZJ7ZGMd8W2lGOGjwkxQ6csGzA1vq51ygVu1PL
1YndxnTE3eAVPAHjvquHB3sQnCQM++EejA4mdFBpRo75VXi3GQieSphj90ivFQE5jt5gCeQ3pwlL
LDfncj9mbKknliIj2JXS3kBHuLD3UnGG/+AhQu9NFW6SB3504ZqNsFRC1hzwfLFEmwqaaN18AVwL
+ixvW9XkDq6zL3b7tQyr24XB4x3PS8/6BY555cUtqFoeDwOK6HPx7U4Xt4hHCd5/tFC9awPVFfd5
5+HxPkMrKvj3aamZ6Fcv9t9KNLcOazu1qyVzxBvP+EIEgQdUvoyDUBCj0gsm9v1M0ECyl50hhvmi
MLFoR2CyhwZ++Oj5jfJ3yUBEc/QOn+3+cWAhrKqeJRgKcJtMjwe7homQ5gnk0Tii6ir6nI7Zyugl
X9fGPxK+WLou+FPsq7WK7b+1FjT0lOkLqJa5NV/e6owHuhQ+r5Xi8ZB/KHRHVBU2R/X0R65m9yBk
HLkXVwj5rh5uH1xAQcSDXufM/h0VBX988M5s6C2AW51xcbHxvlnKsBc+g3nwmEySS7yBiGM7t71g
/q0UkXxvFFko1mK1IXq+/4dSIqTVBkWBEhZi4GJxf2sCbD3rW1f6O3AohKMMNW2M0uEk4iLoUap0
VcTW+oPR8tppVvjIQf1DRDu6+w/XjtKDBwmhHbZQ5eN5lHzUvBDHVK28U1v20MhU+0y5A7+WJBdH
JWA65z9TRrim/EQUNjfbh0BvJL5KIxER8aUX5x7C95NZ2+vISzMO5RlTLeSOwwCBoaK5piRQfosW
m9/Z9y7kyYbYuaZ2Nn11YxdY+nwXD0AInysTyRknome0xIBOiTFE1ZavZ8nX2Hlj1akb/7lfPAEZ
YH1jrQzKPKvYWRmW6Px5HrwLaiFlkGue+gYWdUGh1vryBFXzschGS+t3hQFEyGrIeXB9VnQ5nmLR
KYfMaeiLCNVY9xTS9f5RHQuu+96GatM3sAJ0iSxddeagcdpYKrGdsvGd0EEjvhFfqEbFcvUK/yNl
WndvrAmFLxkryjOvmq/FOwjoTj621+44qdXad1cO/baj+m3EcoBzUNFEZeSvL0FErTrD+DAAAA9z
yaZnEQCl6K8zi6TV0LPh0hnTpVNS2bQEkQ3+MuOZwNLHyEY0yCN513TzVQnAifLoh20gpN6x/Jow
D6f+5rlhfzTQgeF+GqCx4gjISgCWGisz4tQlFPt71Eeu2g0Ma/MfmwyF5ZXB7ZgdIcKSoUt6+ygX
OeCT33lkKGpBWIyvJgrKza35dVNbWBPXzp3oEAqjdL01llJFLBwvJ4NlP33zfwxnrDuNjSTjYR2O
yESJRr56iCyd0iRP/mJhZAwiTrOdU44Ta5VCkwzOEKV+h5D6C6CKvRZbg0+/rANxw1pwf29xC9Ku
KvJthXnO8y2ekLehnkEIGH+CnuTWtNSfSYoRtWQH8i7CVo6e5qAGBJKhZMUGEBkY02eOIsxNfpGt
F/+YYu5M8p2c70qLoUldLiQAG0Frc8qm6xtaxCyDHp0GeVMYMVp09vh+thU6ioPHHRV0FCzMwBVB
Vj7aiFOWPL0nrBA9YotXxg1csQkRoZGSaX/3n59Jv/R3TFAiowo6qsUGIIQPUatMzz8nUpPu7wtQ
j3Ly8dKD9ocMcfmr8Ccid+o8wQ/z/cUuI+eatmF0WZ64G+A7ijQGGWYyKCqqtGGFzLqAP+Rx4I5z
HAF2L8R/Dxrt5lf48KuvMIltpwgzn/NHz7qs1VnqbgNxTCSsjhMXz/o0xhKdR/oPi9cCDu7RE8oY
mkCN4cvXCdH4hRdNLjOoK909heluF/zk07H2MtUiHZOIt/ek2I/AxNSCkUFyO450qAJsln0bv00Z
6+alYHORbglyUJwHaobm0FYnX9+1bTQYXit/99L4LDzF82qeDsaQeZ2Cbkven2qky0TVRkBNImLD
0l3fekX69afvDgA7iCcGz306IbdaZndCShLP8GqhasY9zRESDJFA1YFQSjvHXqQmwCInEy7oTzNp
9VRZU95clw1tvuS2KhqHsSABTHMtih4gDpv+vEk88U69C2MgwShjWFOWuf00u08s2kWf+8RKyft6
0drnqbOvVpxEejT7lvRr6KYwWdA7qm/IRiwCz/F4+bg4hez3JRb6EFYHe5hf9+IOAIIk3lwlkfUb
hccIp0sok9Lmlz2X3kt3uptLbjhref0R1Na5H52sxPVGk7CSrTE2LD9jerT/o8ELUHiRAWLeY+97
QZ6IeT2LTIg/4mJAj0kYhRBjQ+DfEbtH1UgGMEmgSrD4J7s/919YqimX4wLcj5Mv7Kl5hvjmXhF7
+t5RWf3c5Rx/ylWldYba26oWb94bUvV2wgiIcTx8WxI6SQ7E2aGU1e2jIH35TPySEkR9ibsZqQCj
RveEYm/ajM/2Xir91HixqhXC/W1nw0yaCW8D21c4F+lKcdmoKNxZoJ+XyssnfRInGgwGbmRoMt85
R8yEyrDZ/AqCQzhkdFLGGAw25hC6875d/KnIPSby15q/bQm2n51fjMGd9sZX4glT7kk7XeMmU6Fz
xvV4QLVwDmsJqH+0gT1j+JELjMECSMJU6fiOs49O0bgmn+ygM6MwfX/bqhW6kwchU2iihWmlTe0k
xOsbWdbxvlsKrmFuWDXf6KgJCXLwDCg1tij6ORbQGyw8uE9a0+5qVTXPZodWudCoDmJDiKaT3BQD
E21NAX3p1HHx1tw7EgSSWUZvEhdcC8cxDTenRsv+KFPgWphPEN2a/dr2oXpOGGC2jLERQVa93ld/
V+QiXk3x2dyGXir5SOBKostfbRE9TSk+LiBm0/C9YCeFhx9KNhvGBwFTWRTj+jpsN3mHcWs4n+76
eb1XLdj2d7wqUZQBzJUkd9QpukDab/6of+XUdEUsl8Ig4ksqMJnSlV0YqOJIiOMbPPjOSqEjNQrt
67urFu3WpPvd7okqjY1MUVRLfL8yr/a5dRYuEs4Lr7hcvGc5PFmc5JEejc8fkZhwLQDcTRKRx+ez
7KXb154VNGInadAl/qnRHxEbaReIVMrYVOK9phzLxnlZh/4OBWosl476gtcFNAv7Mmi9oUIWswSu
EiMIlIIfYGojYMzNUS+BnzfykFGIZkYuT6aKD8lsv31xm8+dSR4DE53iV3gUc4TIWmz5poWOQt8h
7IK/e/c8N4dx8srvcaHrHaVTHxj+vjfFd2bNH9+g9LQamxYQMQqA2iKAtl/HeyYl2ncUBNtX1Flo
NMbsob5LniRT5GK8vxfSUCYfYSZd7oemhk2RiCgt6lYhD/Y+aEWvGGRWb5j5OiXxFmJR/lTdYKsK
GvVaE5LpUY35ZSZqmkKIplolBoD2scdAKK+QLmlxd2vyKPFnOJpBsgPLonbSqmVX+ksXmgMNDl8c
dper6kqPOFvT/+akm6SP4Dn5GotiGLtsQdGD7vRQP0CYagTPAeTP+1O50feH/c8c+F3JngPxW+Gd
DuKe2mC0bn7FhW+diiKaI4PBmaJ3pHKQWGTi5UUmh1/ifCXKULwMG1FYMI3fPo6REf6sX8N0unT6
whfqkHWUAFqshqnOahbWWdxoBukbU1B57t1p8PIuqbCtJq0h71Avdt681t1lHWiEGYHlwjhcSDCQ
qa8iGKm5yog7S7xJj0Te1M6AerqFUOIgJvyxIW9J6L+zvgT2pbtg8tpu47MQJELom0zoVWGETpI2
tK/arDHtrTX8utK3Sed2GmDS1Z/RFClv5R5VtQfgZJ7pxqIRPsOsZHPiUyxnOHYr1TvqZEHpHKMK
+CiR9+2AsXrJUt1tXKK5BHsmM5S1zk9Ha0H3eIkyKaz49x7mdpk8bFUonafS6oDSKllCB4U7A/71
4KsVOIqO5WTUXvyzIX9lELxlUhRD+pJ4MpNx2+cNvxE3YgcK+sD/Al28tuJloX8RVI0Zwt/pVEmf
3jlSrVEryRISf+ibUrcoHXwbgtQR7xK2GYotE0qV5JyARVEWuiKg2QfuxmrFKVB1unxTvpHbrq3H
3o7v5IKdERtMhKGFu9g/DLLnJjaq0P7HFRa8IVts+Mb/kmOlax/sOzBb8RAmBD4JRXrjBRlcPWYM
akqiFc/G/obDG44PizGncbIdLbnNCJF4dttn8L/2NUkVzqiIODEnxkFB1OED/5ihMSSILycw7T99
n1J9D5W4Ur1tQx/unyD42KJ5aPODdZbFD2xVjbp7M1PeDQBrFiGIl3SpuYWJc5uTHDr+JLQ9q+nB
BeCkj73Jfx0JGqY4+BKkfv8mbXZjqcxjUUlJmjTKqv+CsgcLKqH/gNTUm3IoQ5oy6czh/DZ2K8vH
Y9UygfUZsMa1q4ok1gjBYBG8JNiuuupM/xE23wwiIlJq1T5w7JYaYtXrIwy1KSGbMuAC5IAaqCa+
nKFAWbzrEF8F0fVLe10eA7MZP/vEAclJWJh6W2RFbsnGIcOcN6zfUAf6ayw2aacmj6buPjw9Oy2d
S8SLbH28yp8f8qnx5XHaVJ1R1MIzPE96nh9CFaFa08RsZ3ByeK7uR7GhGo/JfNqvtuRvIMpKzC7v
AsrcMCZRYBhLPnQDEbTcUjYa9IaUQjcRA1K/ZZadPj151ar/lPKp9hoemNJ5evHJpvpNjnuz6c5S
4ENENP1GMvV72lz0z1/HiCYR8L1mmY1BdXkOHs7OJnEGc/bEROpywm6bqfHIQ60Zs8BW2OkuzvFw
nfdzNWlYsrl63SiepwowccQLcMdLLgHBoO0oMr69jExzoRZEcokTOn4t+zeffA7F5fTN894hHWvb
iAvYYymmoRwquOnfzHl0R68zFTaZSViZo6p7xKCK1xbXWGuP5rMI0dt6h/Y2fy48hobIKYjVkwjF
4HR9Ld9IEGIMgSD3EZirgNSxJb+qHO1PkLMrXfNCFfmf+IRYuNdcrfZp5z6Vp18uypSr34QFs3Nc
B5v4UCQjPHODGF+C2MGvpSIhdpOP4hIiSOxTuRfYbz+z782cCPJCAFDiFQZ3z2jRjKuzgkPLh9hz
JOG9h0IRqMLegfhrGFJGap2I1Ghl9ikmBmnO6vuV5yliu9nJ5CMRjkCbNWFOl4LNRAPxkyrqhFyK
chp1PUHRdmnWRt+dxDonDJuEydNusTH09Q93nhmJoe1BEBhKDcI6tAjx1tz7wuJL8qKKoIdwKei2
9W4v5oWrQ3vONaMouZriTM4afJzjoATIcYhKsX+x2Bus3EHLgDBapWf4ZH7kh7n6QK7NtrpwFFIM
1Mr0xhMsRYHmUu7wjxQ1yTTDbSad0iE6I6dOCJjsgUYJPm4KlBsMFWn4yCxR4VwDVXIpQJML7fUp
jMUIJezbulIx1OEZ4jbiEq0jSQLT+AVGEZ9jygQ07uru8pdf4uWaUVAmPEj3/NWI22wVXhkwCeLV
leWR2ZyfbuBZQGn4F9HkJRIr086GSQ4856JK6c4qwKsV35V+CXMdco8J0F/WCHK9TrZiAiQ+B8rl
hmRLj5sqbBgZ0ev9ATh1zuqhXLItDd4O+pcKMFSrAffFAXpNLu5nFsRYfQPy0H8E6YtDpLjdxQym
nacLTJImiRF4D/Z/2JnNHZtl2t8Gro0DuBjI/+C8PHCH0HIWkOYsz64PZPFUSrtpY8d2tGqOJXhF
AqtpUU8upUiZSbfsnNdayUuH1SoEiPtMLs2ebLT34cG5XMb5w4fV1IF+AAqPfvBpasMUC+RAKCZf
tCsIKky6k1E0cDOtVHy1/QxX+6OJlui3t45dXmGzlJy6/xoQ6XKgIu4lSaMwdV/uZ+8ceFjSnI0L
vVqO9K3QoCh+CWLAjgqQjhLjWi2xDz1ZHl5hIwAOA16i0qMhrorNqesaKdNYxs8pS6VIixDkVpJY
ajbe2oeachqgNI9Scgdy7Za6E8/g3RsYYfb78R+TprzptOSYyLWxLe5+KyAKSnuO3SOFVeYeAGVh
BOaqFSUPsIE2+4EL2454M41nJlVCeMaNWx1zjgHRe7luIXwhG+83/03EJhASli/ebsy60031gKeu
WchS1PWtzzd0UbsGe3IOXGhh+b+yBc2fVWUNmQ7pWzInC9fKFS7LwR0xtBjE3FUMpMAkYD2NnYxQ
OfMvUXRF9o51TKT2aLfoBNMbLUb9DTLv1s9I5WbPNmuXtBH2dlo4ZO8jkDmqXUP4xlbOfO3TpwK0
0txJ3vkjMK2wadAhK1wzbpw1W2AGrp3u0Vj3is7eBZJgCWSAFRFzZ8J0pIQxQi4ph8TGBBYkyBBS
si/xh2PswBdqTNWcJU/XxzxQj1iqM1TfkI1UWZwSO1Z2IxoQRYJJnE93MShsZBEqmZsdRTH5rjMw
wBLQ9oMfDimfFpXwcFuJFpjf2VvXvWA0KUXsWu1s8Ej6LllHf9TAFpM0qjVGetnRloQckMdSLeyB
BVHwGupEH1BxQ9xkQpeubA++daFh8ziPr9SqkYkz2ae7THGqv1vWbGGOZLtp84WsFX3a9irgyfmF
bbfBoKuVsh7I311wsHQuwJjxfLBTvYqaTOzaA8/v+bKYeqq2NELGCwLLW6pc+aW5FooFA54H6bH/
cvdiT6R69rkuMR01n9X1oJGNhSjab8ugxteSdvnj6qCNvmqCOuly9Tiw/nGqHt2aFVmJ4lrqd3Ah
28I4qoQtX9yXf0jGJUCNcdlzsIXiU6LDlk3WPXaEpzyJlg3/70IFHGiF2U/Z/xV9EaZXSAkNVx87
E2Q7Av0P93NEJI2mVYfEPFZt9KEg3CucVx2G946MCFcjX7wcCY03Ybdj4/Lxz8oLDcWmcVquFoFh
vNd13E1/9l2/e1SYO2Z7AQ1AMzEsC7DdWjYTxi07IxhEMRLy/TC+tJM2dEiTkymw0h0N/Cb9L25f
rsa3vjF1H+4ANcWOLTHINNeXYAROGaTD6/FuoPEEi2zJYjauQMYvBUC1vP67fyUdDXPftHp5j0Mb
OkN9tsmgvr+loXR8R4fQFZ9c0ynVYD1IO67bUuYGtKmE/02Q2BNFxRVb7fiZPUQXilEccKaMWAKi
TFhwL+Qd5nhn7Z3hJ7JKEqdIlBd1iO3sGDX5esonO4vvidOB8WymUGiDv87WA8FqR8/Zvg+bp38a
Oc40C/6lLwcQa8Dse7M3uRdZfHXULux7u9K8XZlar9jw2S2eA92ueIZwnjIC2GDjSzfb05AZKuDG
wel+d3SXFd7YEshx1frPHq9szBaplJ0jum1Lb3bMLjvo8DCk3H7e5M45MSvbuUPwMitR2RJQJ6of
HuFIij9eYjQrsKufmJluxNT0/GPnYSzCj0zo8lUckTixlKLe8roEALGqGZggeBbpmNrDs/O7ZxkE
fjFIBKBAfc0oUhmRkTk6k1SsO3w2UwPRofzXT7bVBjsAYg0iVLYIuH0sKmP7ONkhLhvU6unWC8Ch
gXwbbR64dCPo3FS45FsNx2mr5ER1wl8nq7TSchorH9x9HX0+0+sI7WKqAx6wxjOXjubvgND3oTgo
qf2e+6PUmGg8Ur6WUVnKqohp+mluijDizS40s4AqcHoROCqwVaD2xEByAFZFQHDK8HiKlgCcOxPX
j8Q+Rre7M4oxIg/1UXxodlL3QDeKjbTM9FBptQhD0GUAVubHLNG7Kk9nApWVOxggmcYIWzXCz4ht
SKLQO/xu9oKmjO9NFQDmINbe4c/7hbE+GBQ3PwJ26cE+N+DCNiJP64pWgDMQfRMi7v/p9/tdnB4f
6eqYxbQN0NJ30BozzvWoxXUU6ZtzMqMIomn3IKNbCRrdiihVAC+Skw4aEOy4L2pYPgpLMAg+Dp32
qLOdoyRMsaUBE7pHL2BDHEM1rNO9YtpIzIPp4wHaRHE8VETd45Uvs/U9/Kk+YHFKLxeoJxLKnx8r
daWQeLzMYctekZEgCgpLHHIX4aufaSBwi91yr1bb+fdfKnoavwOl0uq5gF422Nkn73/V/GpWESM1
hcpMTrlkyH+i6rW6iR/aHRRjdqcYBOGZri4QppTZewEajurL5qEo2nKB5jv8Qt+SKjaTkkw0OvAF
vMVwbRFgVKHAtpxRTFrWg+u41pzNqLBo/9O1pNM+Vp+YYMputWJc6lALtREWxYhjB3hw5GITI95m
lem8X33+IE6AUXzovJ+hPGrwoKfU86dREi9e6gqj5ZjkV7NA3DDHK8Vb0zqfQbnFrnOh6b5wXoAG
obxgHbizTgW8gVatFdOdOewDsFHC3IcC2m/ewqQEhvTNUeDmC6jx0GR51SnUKb/pylONG3p2T6VI
ZZWsHoCQnKiUIBUJiARJuTDOelT6dBx0wjpjz2td90F5wWYqv2iAL5XS/2l4Osb2T7BzSWJbIJQc
if78fkMkBKsWUfiyPikW2J3VoGMxACw4NN0sdiAlJmarXLmoW9/ZDNjc0PXhgGKaQOE/tXcE8hpH
fbNegVGeRRU2tweXwulkoZZcV19oJyUYIv3hQedyArrwEVPwDZC6iTzenrkPE4+Ce6N/B/sVPm2Y
VwAjT2+kEeFyhBB/gC0lhoobrmVZ7lyADp9VhG0k1+4g84YS3Jo4bdtl7zlZRklTNB9U9HKzL+w5
wf3D9Do4ZamJsI8J+or/2SDtu5EX4+uGznBTE7FWOrNF5pVDCp9X2CmdT5hJ17PU6OceGFRZlYST
zc6TP6CKE4qvE6rtEFh8juWsJfqGUvjHbC+5CAJ6yk6LEFrHKP3YQRpMTadsZUXqzjGz0kIRElQP
uFxeybz/q6WYol23jcmwiN346ABTitJFl8gUB/cG2MOwYxjotb6nzds4/hLV6wFDbP1cvcDQ2EK7
5qvpu++ZiByzzuoW9QgL8yv4J8arIB/4lGTlr1rg1hGhE5kgLtyIrdIMpJtwwJ7tx61T7cyRMeaT
d8kQkBXmAlvys5F0Jses22t5TDvSU2U3R6DD4yowU2mFyYPgo8PaQaMwRyFlyviglDWVWwC9HhKl
UtNuorhX/MszrtvtqNfvcxunPiAg4N7wADTZMLc+kpHO0MWThsSZt4rTZn8paLG5m1/+946o3ZqX
J0XKuJVe1kf33AXiRE9r5+ZrTvqiVV2CVC2XY8DU2qV9v0AQRAT3kh49JKSOGApcdZQJMEXuOyAf
w6jPUQ2vOp/oE6lT0TrATcchr4v2CsaNXE+T0IuCKnAP0Abk9T3spKCcykvv/2iRir9zfItrPhZV
cHAgZpQJCZ4OLqrxNAHEreEJHwRmV920CAXhcBl4GlRPh8jBo1AKLY2Kp+a4hfuiKbFlLJxlAWLm
dy6dXvQgRAcWjvxGjnk/viuVYeWNpTOe3OYXnCRIxx5bZlB5oC4GbBGfdKLT4S720KaYCjDjayb6
qEdtw+yIcsNYDIwWIFAgeR3uo2gUHU/9F/Sy6oLcaN5bq3jT87Kv5MBntR5BDJ63Z/6bhWs8rbos
B1Opb54340sqqiY+huwmpYracB6LPm0dxc5xK7G186gibU6iwtrqXXYPXNfZ7lBwoVSotZnjCNCZ
sbZWl/FaL6M2TAT5O0CsvAzHv4HPeesrG/qWyROk3n4zewplG5BGUkH4V6ELApUQNyZb65r22nur
rjkQoAXzadxWAQ9lXOOimpwJzLX5bb8INjbZVIZVU43JY9/zo9Tbik9PiJKlemx0EvYtTr65RaxT
6jE3/f4FyoCeTkdbUP1qXsuyqo/JAHfxt6T8uLT7YSSlmVyTMnPgD7ritnY/oY3ABk3rldq6XWV3
qpYNmIdWD1Hny+IbLyu8ujzLIBHDd/9xtY9RGQzMhrJ6lZ2S8nqOr9+E3XD3QA6YVvzbDqISU+LY
zkp8YeF5N9iFXesJsLnbW2Wo04s0flJRBxpBygv/1A7dz5RTBdRK6HyzHkvM3MAoV/UgUbSL40aO
TYB8eG/A4FS/H3f6Dg0nBPH5idV/JwEoms0nMw5N/81HyEJwSScrkVyrdxtM5qkgHpMNZmiMwtLG
VwujKBgLu1za2ipkLr3yLwV829y4A2DMbrVF1iTfiN+vLhDvjAJ2PhvPmJtNaTLIDW4ffL5qDTw9
NWqXPnX5illwFftIVIkH4MyF+rn9jPdW4VQIF5REChQBt2lKy0yN7XlULc5Zqo7m+fV+sQX6wVem
25rwZJghmGohbwokw9cu+8oR3TSRd6sm5g5rlZfeI/Ll7QTLNSnf2iVVxRaAhhttPdJCNfPIkzzw
2c3b05weYWSZGRDVvPdZHmN41hr1Om9Emc0jYSTB8Q/kaCHCBnJc+ckXsdTI9ueXKmeoulYxmsV4
EuysJCkvXAjrXZFwSD2IMulEgjVH7fJJ/6GU6FrT+z+t8FsVCo0Fhdx5e5IX9yquEtFD361WZAGW
8oWNu6XEwjOC0GsKlFLoLUXDIIe1XBLuznxZNELIy+dsaKO6UOFTxiQFDGX4LDvmsqBGTfiHZHTi
xNmgchi9f3H+DXIRJGL2w+hMD/iD+LxYH+p1nnuP+4Qiq2xNS5IsMAZV72HrzQzRQX7b2O/Dw5Fj
A3ZX1yN9bOuaKVeol9RK+8SzF2xhpP5StxRZhVKI1nMR2GCgfhhGtEbarfJTS4wJz1b4F/RU+rHz
FB5LD2OEhQTh9m+AG7jtMEHBKZ5mreb92PDTGOU6JuNWvZci6nNTkgpOIDUuVMC8qrVqDFBwpAQz
SEwa9nZKu8/aXjR+MOlODII3LYkJScNobZMTcGZh2QTUDp8wFVz+3DOadEdOGeBI50RMu1VZ87qo
DQ9etcmxOPQhPRrpfuXVDVoYzha/qwwJdNGBLwF51lVhjw83zACmbqixlACHNHC/vWVm/ex7OhbT
jXJHxhagCTZa5gLlqAeF1H0zvGA5Ocv9QQoCH0E50gDZCrEkh8Y9ETAc8aONqKHL5IRhGkaHMI3P
Qqf31qsNduN5LzY1vPuIfJtFU6zw9IIYW4eTKMElkbrgxMvY48qXAttFla6Tp2UPdzfXQA0QA3Wi
FAboQ/98rE/kCKQ5nk+Z3Od45TVBcirfm1GPbotmp3tgFdF2k3CK/2GqT7mC3HlgNThp6R0ulHjk
ouzIvu1RmMN2C8W9IkId+hWyDLsrQmaLUcu7VtWwyUdld3GRrs6CXlSHLdhHyKKavGSEZf93uhm/
q4HkF4AIv8JaNPvYQSD/BUKRZMDF6rFUMIp5rzcKWhfT5BmUgFUi+cf263dktFO/+pCU3F5Qit+c
yyDJTf7TuLDxH6PwaryelD7xitukf1xvmTZrXkvZWmI5viMN6v4AS12W+CgWJlDOtNrraYU7SOcj
cBskzgrpIr7plTfVC9jRFTCZpg9fvBRNwOHopgtucO29g0Tou2Hzr5rNYFvEfQ4BfUwA5g2m9e4s
ImCr5hCRGAMJ971eyBIu4T+F7CQRE4KCMx8T6w7JYVFO5oIINJRfeqqfVQ8YwVIzVnYnPQpmtFgP
8Gy9HdvqbqNn5e9BKIbHttWobSHcd+IisgB8nHpYTHUteOp1EweKkyqDLZbejzg6PTWX2fQ2zrl3
JbTOd92ksNgYUT8Hx81zXJmFY0W+i+gxx8tjLf0xFLyPt8hFO9+UsAiG1wkcH+vBr7PBwfVWae2I
w8D2GXcrSVoZkoLhlpM9VaDQ8u+svP3SRcSO8QUHUdOL9zV4CJgXE/yiB0A0uNtTvwhC/qlzL0fT
hegdf+/ZXyQoA0L4ONc2+YoGmrZ8x8lewVttcpL2OuiEqNnqLrxBArX/mp29e3EIrPlOn8hHDLSQ
ssWYZTIgprZm2zlb5C6xK6dN/bK3XbEB4clX49CFArOk+QEdPtiaqkmlzdWa5BOnKFWp0vwQ5Knf
qjKQVR0HjkWatUfHoPWcsylAhnvKDu8pg4QXZPjlQGeJa57q3n2NZ/pk2bI56jMNUMnFAwB97cAw
IoeQKxosGT0/edUeoo+EzikQ1OR7Up0J4DF5UPm+h9FhFkLv4p+ZJ/AuO+54Paw50vGNddB5tONH
7br9ps2csd4PjxdarvOkBPUBNvqSsL4VALxnFqQh7HxxfE9qL4ym8fxzK7j0Kbsk09vUlG1jEFwp
F/q1pUGUm9DgjfPi0BjE5ilqI5OjPHhekP97fqwieD6ei3LWUPg5EXmhC8jKkBE2ZQWwr+ze1euJ
nSohNaBbbpFSpiJGMwAXWVBP64xKwM1hArjxeWq/OS9pLTZ1KbWvL2b0dpSid9e26u+k6miwk1iR
IEl2DBtZdvJdgGDGjsofufvKn+s/9ET+T/ckytm4D6Qvq+vTqx8nkOXPfwCOXfdGnCfSa5ThwSKQ
YSeu41Hhx9R3/hTWKiiO8UGoHAMt+eQwtJTS7B44a6JDFLAi9kQB1JzvsVHZ4a7ddvPm4lZ1n9V8
S9wgurbEb9LZQjIUBKPvP7v/yN+n9xfVwueoWbO5/R4VmdfiK2e0k+wEoCwfCEPYXi9KKK2s4Miu
B78pgMWO+QYANSJCcSafYOTbgFOC1kgl+gOBnCTb3uM2QjJaDd2V7k9d4DsU6R/Rz/4JUdid0MZD
vTG9RGRnRCPitS3bIYHrHu4sN0uhgehk2FvyszLqX1Hs0UdlgWwjC3abAtteWwXP4iC98FOOrQwv
cQ2jcSK5U+4HqUN3av6lyO/qbF+G9SIBLIxnigNupvHv+kKEE/JpQrSK0jluKe2nkSgYk6ryTg85
XvlFlyvuw6ErXwjP4R9g5pGjRHHZdvBb+fwGuAeZRAiTDE/QvAeXuCeLQaZZNvV1tK9dCj2F7mec
cDNcHCV83hoeIAEUftZoiQzbA2oXjlOpuwv6JpP8ECjSC/olYFH759AOE1NzMpoKMGbJDutrQvXu
+YQ/Y7vMhzvx843pX3OTbkNmpiUr3hlaCnJT+UQ7J1vWLblZoRgWNeNTWONS8Be5EJVWSbjEBtlD
S97URjvJhtfc37yGPAhfcZ3yv5kI23mv1D+WnxQ7QHtXgnsr6jVp6QRDlYmZ9I4VVzUDd2yMyi+u
dWpVvOCQGEyvGpLn3D4m0JlkbVJUgiRNxnz8sSpae3+JD57x9cEaPwi/WIoFBukjB24B1NwfhYEW
4fkfD/EuBiUB4Tp5qEV/knsRYWzOjslbc+KlSikZqShS+U9BkVKl4/80P45HJEMFqJT/pOWEJ414
4Ipnm9tMRjDT2VvuEz8yV+tqeJRHpjSsU/mLxZe2gxznOhHCB/tDYJePyKyTA+90u7H2DNOr5MPl
4T+m0XEV1ew9kwyAmgzJeT3+Rr3V247MOxVlFFh5sSmAPSIQtUGMP8BpFfkKcZJ1+46+GDhYPkMe
xwSYogAcEK0csUho5f+9hr2IvLlIz1hCLp8QMGNTZHMzBDCLCsLROS2/wF72PEy2Slo/PuidFQYL
pD245avLBVhFiesBt/WZxWNUCNDBO5emznzJy55oUzDpLbIeDxc9IzuuPVFnwbWIwkxzkuSf6gbI
M7shCGBTZh2IGUMCfq4XH4PC8V0yU+DJskjD++/cfpQgRZ0gl//zfUTbRgxXB+zywXvk76UY6o1b
ROcfL2c+S1Cq+hEXtobWBBd1c8eWdwsddqLtD1zV4dUT9pcL0dc9pSDS5WEvLdagLrdPQhhwcSAn
a6WDkpjtglo4saeLqjszEC55aK12FnOFVmamOX2RA7L0KFzqCUM3Vmo6CV5C6RzXTvrmFmtpVJji
XKhA9c0kPFNvze2sYKAwveAVf04hlZtmsfWUrBtHUo0/I+ceum8VceuCTnntNVvkJhJ+UpNaizjk
GdMoRAwirOM6wgh+PMOK7VIAufyja/eZH89rEDRdxXAt5EXpFI/Ql/1+ggfrAioBBYgVcXXDLnTh
mPFrDNN2mG243TmI+OnL4qJyWG7BT1wyICRfkgI3Pi1nJQuIChYWPmboFdO0WrrvD9LexKhOMetO
+tnxNt6kHiOvn+HuYje5bZeOO0rXYOASxbRk15JdIR7AKGEzBjr0nVquPkrBuyQGrKgzKyx+oIMb
GG3CvNZ0sWxB19JCPiwmI+qyO+5M3ORlEEvoaBfsJNVnkhuOEO8Rmgz2Ofe41uOZP/PIA2EwQgxC
96Nx1teOt5GBg2EwGKXG/6VDekaMVPBnJyFHCp20q3cdSrmFtshuFcA0KL7g7oiRIwpNqzUW/ZG8
sBnuQ8pYqK5SxvE6p3ejSiBO8f9JQbLbiEau/R3qk6FzjaMqys2i/Yc3skFl2J1e0tMpVzemIFVo
qhCw1V0/2K34bEX2ItZdtqdEBWXqCWe8cbbWYt10CXV3R4CreC4IjAObT56bvWVXUYCf2zR6zNoT
Y8RvCebv973/FY+6VTeL1mS4Iooh7a7vUCKHv93AYsYk1zSnPVTPbzhM6Ia7dPeNw/7QYjaLEPcn
kWTy9v5cVpFjz52R8cZpXeB2qXgsD+bbIQV1RYdyoPB1FN79vWCBilMWYlQQVIj6zPTyL1ls5Mom
AKUu5f33linxiSFvhOrE+fnUJWw46Rgng05O35FF9z1+ud+R8HQp8PWvUc0lJAJoikfTzxDRw/Lx
jISk3ht2RGX0ZV/osNt157ajPREDJFQhUjtW1s5FrWBVBcd0Xudg7ZhXkqxXQHUA5j85toZC3ZDl
ehOgQLCfcuiiLPZx4WsBmIXA/2f6OkN9nppO9nS4K+VEoucnWp9OawaMpaUlWIeZwuRoypS8TmEP
zOUKf1bPm+b13FEoDStybNw2B97K4r3/7W5Oi1aZy/P7BQTPkhxC+/kk3O59fxi/tbggfsvpVY6/
INFaMuwgMmimCprDPXNJq5a5UfRzXreInfOXXWR4GpoUuPK4aHb/9a/WzxNatpsMk1h3OlMK44ar
MWiX5UlRdcq6I+vwQkvFwzaG77ztDEtb5DfWnTeFjkKC3E6CiRNF+4Dezwz1LCqCd49wkC3O8DVy
ut2jA7eLIBMunrcduFa6Q7N8Z4nYj2H40/eltQS3VxfABcLbmduu5qN/+dY6BQpRN3MmhwhtTkeT
JsYgOFFYfP8yRG2NLUmhQGAc38VwDoI2cHHAOX+Fyuc+EbxvWFg2cWxL3+J+GzbDNUzwe7BKKZsm
tJ4MqvRnpOEhQEWpSX7hZjlXYPV3pCYXBs5NWlcASLrgccv0SHf0J4XKJ8PppfgviUY3EaTEhs45
k55VJzYRriAB7muByf+adu/1Kn2e7hymZ8QNi4lHgniyULgEp4OaSu/t+fC+xDXHtohw7e7yovMM
bL5VWSlPZ4oQIHFuUw3MX3LpdEV5StBS648Iacbr1v7SYt7IxF66PZvAkPEosvhsLvMrtDgIRbbO
B76Xeir9mlw7InyOpBulgLGacYk2y3211yVAKOypOqjRxFZ0YcEUz7HLDSxJekgBLjeqgl2lzRfc
GuwWiq+CiKksxX29EfUJtvmCmjLTDiwMczZuhfhdmvuZEx38gDd9otSHTAMyj1Y+gKWIdBAoRdbz
Hn5XGTjjYD4tgOx5WETNcBnuzPXsDj0hVDOodXf+gdYmvNPaEd+PMTaC9I+751Uiw3frBw3vcmjm
mL/2BSHkEbbg4ZHtL/sG6oIlJL9gzK/WOJKsHyfSeo4tAbAOKsRpijxcBePzbkAhWQ4fJQ/aP/In
wDZ2ZJn1nT71fpj/uQbOoIHN84P8aVOakHg/4WLXQhzAmWbRz+UU2tydNYq2MvaTtGUHlsN0KbLA
BwGhSmuFfKEagvnguXHqlm07Lq+xEe3Gr5aZrS9VvrM75mwbLJ01AD/HPvEoYW5+Wo8lOx/HDKYV
aAZMzgCs0C7iCjC478SRpJWWCVv8Y2jGcmlcgiFKsHqPgGo6K3VAXzDQTf36SqLWy6gHkbZvyEgb
F3CF9E3u61LZu8SxsifcFmccvO6hZ8B5Uls0WlaCyvcqJcCLWkgwFfvjCeepb1H0G7dmWrI6v4Wg
DTA4/+zzK6CQAZoRr000T9lOGw7ZCAQjHeVvbGPZLVg4r/wvgXt9CHhmQ/X/4A3RQ6g30+fcUb5X
hJnhYqrqi7wXMzfrxTdCqbotOBue2+ovSG2ZEHYs+ilm085XHyGJ7osEfmAUkWulJbOSoBcDsoDw
J+SebcBQf3aA2pH1wX77SI+linJGruwSbsJYZ0+U+DbNT+8NwroN3FjZLEZDUajBXfyGsDMnGqfU
e3bkLQEhEMgPnHVMwy9w4Q9u9JPepj/JQlmrQJ+vZoVMn0mSMKnRgcQV6NOeHlVQJ6XCu8MrWjG5
S6O7/PscFpj4/dsFw0Y9kpMFSPeZwts+Jj5YuDMHL4bndSiGQCBSETVLnT93kRu5Qmx376/BZrfb
cTveD7DH6txUtaO65ohfL4avrv7XhaVvfdyGj+NzHxWkuRhuBIkC+hsYyYbEYnG8j8LObsMIC+Nt
uLhMHljzzGdcsufoiEya4g3NOZYdLYpsr2wVq2Ur6HQIwqKnppSo6q+F1md3FBBp9YLuH4UMxvdR
bwrToz/SroY3FyjhqeYbN1TtorltPWihKsJF6Fkr20BJGemkbF47QLedbm81ml7+TlFpjQ7hR/1A
seHf4/wAe+3c2PTDCXymEFPtDLbexP1UwhhsTYoolZUK77jDCSs5jneRQvW79fv3RSjk9Q7Fm7iy
mVZEkqeWhcqyi4cusVmLlo/6UNrVumxk4LZhG2wWZw8qNwTxSWJpCA3KdktnnPUWr88q9aC04hb7
qloUR1TxCQDlb1GIDpdqdn4OREnOMsULe5Vu1DGBn3jrPEZBf7ctXkGGAH2TcFCtpNnC9gj/fKZe
eMrZ3gPK5X8HfF+3idRaMV0Yyt7aaqGuLzx9Alkc+guWURrQf5NzwoHzUClUXpb1eDsKOxwqV4bD
UwLI2q8Md36k4+6CPCP42VAucYMhSpsAi29NAw5Ziu0NCQxhkIQlf1NDUUStdhGGJOMwNhImgMQL
yujsQsldChNC4YHpuIrSwHRzF9abiY2Svk9wFKEFwGtdZA+qE7YzABukpBNoRz64y8DN/r2XDzNc
Eazh9AuAO878q9r3/a+GoHaEk6OXI4xIObeYNMPyXV+LinotX906BthiS+yqFCBpGRYFqa03lVL4
JxhY+UEzWBy0O2kTI5k8/iVS7cAXNPpUadC8Kx9ai7xh0ZKiFHRAHs5RyYm1e6ZIZWXMBhYEEWyn
7AMGXbRm1ze9ReMukPcNoXtlJxtikiGh91lkD9WJ1B18ObIS93rEucOk215TB5EXpDYyvUDvPo/A
LMeF+sWfpXRb8HDwvlkovS6nsIpK+ly8hSNG0CmaSa94Ql22Egj66+0LuLOVsTzv00aIcExFsEp4
RH/NE794k45t08VnYudrJ3EJ/zaTLJX7XgXZq/DnVjV6ZTbGWNIObSVU3/5mSrLV46VNXRXeGT+N
nilHEq24CN0l2IMHku+DgZ+Pv5mwuotUhJcSVevAXQoNlaB0xbjR/UDxIdvUZOJynrg9KIar5/YF
F5WTFoNeHcmuUkGwZw0EsQn7Qp5QKUQopc2zKqzn/0R+6ggtl5Qqsv+Ecnk9SzbJ+QRnzjkW3+A/
+YcGqwdbgQxbd9vbJduQ1xkWxSJx1R2e2hZWmIGj3q18Q4MFcqOtzcZwXjS6qVkSicWPl0AyFrjr
1QfBjuNsCMZqmnvG2ob3tO9Iu75llO4Z2t//EJdzaGxU4NLH6WaARYYpBmDD1BAMZ6bxhzxbUaDv
79y8CRURIP7pFz5skhwajd61MwUMsmwvriF6LXgDLvdZ3xHZtdhXoeNFnP3v5UNQlnc4xFSuyIi3
pI6cbChU7iR1xfpTl+MFqO6Z8FUSp2nQ5HdcGtdIUqQi7S7r3Dp0N2Byvb1t7zeCwgGVRV3Vwh+d
2XXYBbJtj+CgZJ2uHxqUtql05T3bC2/nOSwQxGzAByp1ftJ1/nPVa1dT9KVhBAh0vTvsN0MTegOA
1PwdWtUqBn1dDV6WEY5v+kp2PYxX4EN46CCsgzcnUBCp0hlU/5/oqog92oD1LP8S3NfzU0uX/TxU
FSryh96xjoFoNTugYJ70vDtNUTksg1UM0tCcU+EEnGRjOiZBYjrSv5jlgaWZhjCeqfp6uOnSn57r
qIDQNmXHuSQ041I1gW/mol51/bz+9d0O6qafRiQclMxDjQXc+Co4JnOJuBojvD1DvxoCp2JG7Vhn
TJNHljUPGBCz8VWxn9l35zLRkcSbjaznof+qSkXj05YfEG3U76vzHhwOmyQvoMXUMwL8CfNXmlgK
XacjYT7Oe8aEm5ZlzD5cklGbTUO9rqYWyLXQxJ2+eoInYF3jJ2nwKKtAPid0EV94KdjkOx8qMGjX
uN33dVAfIvls1GYxtE2rRuQWWwTheP98pFHyxd2dC356K7gaiJEsglOlNOTu0aWkVWPibt0efC1e
eIgNu3F6sOgOE4Wj3qy4ipz3GtUdRhj0ayWVMnGb56VRHXoeekZPekJyBSDuvJz5+mlxqrQriV65
0nuZskN7WF5w8qQYtUJLLyzaIuaJYatOrf6PRfrX/SWkq0peUcak8h6I8jrIBNP1kwf9zsc9Zxwy
cWRaMQD+ayZBo1QKWJCRspJOT+OthceQxtkOJdCFpN7qHVyQX/3SzgpMF3W+PcABd5/wZMPQDqBJ
bEjFw+/pS2g4OoO0UBKCo8HQhiwu0uJpflKQMZuJY5n6oA1D0PsuL+7ENUfJgq+0yQScdcn0p6So
YdJwI4hyOVdnU9GsdBDJC75xAxUmjqLKU8+T0gUQSo0qCkPbWbRVC2T291ml3I1RnPmnaN9V9nyd
MWgL4+qofsgQU8S9qdK6MFivBOTC8GaarMg11YK2E+WLL5xtLK6AW2Q2jTgSxIEQD32paRm3OMn2
tD4BAgfFQXf6gvKeKu/i7+Bkowg8wDOmbm/zqbDxQVTjUnjUSlpLm335DTUpYZXW3tPnPsXdSRmo
iubHwHvo1MuPpW09O1jnHV5nt1piiUKVvvBT98z8Ws4hsJazakF1IIAmH1NnRfb1QcW3rDfDrbHy
nWxRID0UsGxsZKY32oBZtD73szB4n2Knt7KJlC5eRDEOjnQ5fprJu50Ztb2FRu3QicRnv7r6BrX7
so/sgA1mQZt3hM4G10RlDGlk7IfBBuItVProMOjVa5THsmPQoEWexnH4LVg26mfKEOxMI890koaQ
mpCBJnewmaaaea9xzJwCGbwiaAdZc+e9MMxnz1p65dkOO+hXlkmI2IIiI2xWVF71ezbfFUsO6VPQ
Bb3BfpXLchOfQ4+2xqlNanvy9Fg5v54pngIVYf8Khxr0kq116Mx4XrKWjUbb/noMw649SryD5uIz
kq38zwomL7Rxv7iSrVsqLspklzvXQly4Z/k69BlNm/hBQkwdDKdLw50mfylFUbYYaVjASweSMlil
2KzraWBaPiPyqZI7sKad0UAQCFVEgtrTLfajVX4WT8JDRBSlZqgVhLrhRwjpIvdVCgnrht5rsxMm
edCoadDuh5mHgOCWXE3cEtgegdTVrSdgqq/vXAheoxW+I8OeA4bzUV9bhfqt3ZjNtxYZBpjWpv4d
yzd4PLLlgKW2pOU+lT5i+Emfi1O7Ey8qcJhu+6VW4T1reUK7YRKjW82HkFO1tqV3sM/qAn5QG0OZ
QY7ej0DE8DmLCD4+4Tqbq2YLp5GxFBLsFVyuQ+G2pCNqrije+cNrclJ9L79fpFwmU727uwF43vDu
toSLkdp5RAAAie3EfO7wXHrfPdLK4FUH835yGwnZ/ASaR4yD5syrLYxLLmEJoBIaLrAy+fcKILb3
fex1SPAG0I44f3qAO1lsu4L7/lawmlbtibJcaQAE8fX2l+Zx6g2LcfQD3/Wc/x/PtKh6x3JOTqLv
CzBalEhTjVTg/FaqeDatRKFd5P/4qK7ORdeDU+KZn7IT35F7ojVZg+QQE31s+qw4xODQZRutZZKo
df4qbHA1BOZ2Hg4ofqszmZDUl3JgWqvwcydBVfgGJKJOR+ehRx+f6v/MCfSifLp19LVOVDemfRjO
/t4nz/ub0LwvnKnR0R26t6h3VfsiySj8K0+B68OrwykNuakbbTGYm/ekGUCXKSpF6t+H3yiNBeFi
U7c2w0apv2PztcQOnp78I8lzv1A+2XMxJu7iv2sMEu1fhI1uOWjV+DsJLasIz4hvecXx04kJZGRJ
YIRMueLY7yfCruUIYWoF2kDyCXm5JRT1AmaMVfQcX0QbpTKqNFu+YIDI1RwRtzCqHMXwgzvGPAnP
Z5Rr23/wCYDoLkA8w3kyez83PDqgff78VUm/YbCKMk1uI+SOxUz+P+TrfvyZi5DIqz9iX2gCoMTi
PMHe1U3L8bXLUB0Yzp4kQp/ZS1xLh+7YZZMKDCRui7om+UatKvF3OQCoyRmON1EyAx92H9LVRUTg
m3dMXtiZtCFII4mm4l0FyFhMLHVT4zQC9mVLJ+ZIsRuTsU3LlSiRb0JVLsft7dzs9k4sBYY+JMEa
GJP+FabQ7dbiHXHJ/q149u8Oep6+4qIw0RCkbjv6qBOjOObNaX4CWk62tDCOfB84J7WNJa1mvdvE
0D9oHJohgPJpCxEd8LV53u5r8JiMq1Eg5vk5aeh8E7bUm2FGMnGIZR0nxasAS0bmvaoPSXZ/oBJ3
MxGz7d3Co1obG5/MEI/Vg/eQSzWMtHzS+wvtO4js8dfx9bvil2u1Ao718CYwUEeKWJv5jHY6c3pe
rWTWt+FdHLtAAx2HP/643y7iU70wlZxKp5afKwbILtZCIvaBWfTVlvAd8MZpVJwR7pevzqzVEgBt
/Q3taDiD7EsUIGSSOc8LYNsaF3KgV/Sl8HkECcyf4Q1xZ3uOaI6+UfAFeNCrlXmN4Bzb/ZcEw5I8
sr4sgMjTMb92qPyYuU/hyjvBdsEqjF07Qg/xh+6YLFzGQ3JLD8EPkj6h7IDC1Ji5uMtyvxw4cqOq
8RJ2Vn1guR1twQR23RWLQfIt3EqHBV2gH04+sdT3fnOTF1eoHGYWBmPkkY0Pvy09HejoBQoWNUtI
khRw2VkAWLNO8EDR7bb3cviIlbGogmQvwXKlX4Pwwoi44vhDsEHMkmrfbvouEFuoRR+FHfwsePQp
R26Jjy4+/att1P48sHRMznfqoMEkZNVnK20xGyYHltB8Sl/9zofrxxCW3RNBO9ZMs+AzPt4e6hz5
VeKA8ep57fRT9rB96bQJ7vrsZNwS0OGh0ppBz2JxhraA6a4DEFfxR5jFQeI7LzNWvbjeLIi7nmpx
D0X+UbJ20rqi4hkp5nkP3EolIs/cvFcEC+6rjaLuvVsCsi5IA5R41w56nHumQpRyvaPkAHHskhgr
m6MJCBz8u3AWI3sMsyhUUsIHEHqvbgAP+yS/nGjzQGimoOwYVcg29vTxJN7krOIU4/3ANgJh/FgG
N8MPahFeRO9eoSXa5kDWq3xESuA3bnOBez+vHJvlK7RuPtLtnUv9sk+O4XSpuuShpYpTOhBzYHl1
SRfLE2KzC4MvXg1OVVsVgTIoPV80/Ut5HSvpy8j8hMCTZUws5LW+pceCjWYRX2VePl2V80rlV6NE
xeB3M3Tf/ireF+gQvJdw+sqvZrh/5GvJbAyvuz2oauz20rolP8EMOqQNKA2ucCnjx08hT+SNCY7o
UvJ9qEiwwdmV5C48NFHBYz8bK3GfOVYQrfsFlzkItKfscoA0BTeblNTJ+eo7Zk7vYD54PidtaJW2
Qdlt+u/0Ny0YSPDDr8TJZBerHZZ7ODOtbVMS7+6d55/1sy7WRwSV6HuhlPq0HwIx7Xyh9/xgtOsv
J3Rzbs15yd1PRAnQ844Ow82+yhRWUe6Sn1dNRCMJ0N0vMMCuPQeml75cELCZvEXvm7UZpA9IXSI5
tksUQ1J2hKIMGZJ/M22xfY8JXdxjGAGjlmPYRMz3UBDzmVj+AZH3tq3cSqd+I11PHtgKcckS3Yie
tSUjP+5jk2T8CfdKY0O0W30YOkH3dGbzk3vQY66dq49qSjQ2x3ALFpFRkucCWvUkkulF1eokZfgk
QGKgga92ejct8vO7F//Yu8KJKC3sk4YBcT7ozI9PXyVIvnnITK0Gc4hqoWjKBa5NiWDwjwBuqqWY
ja/ywcXAnpKsKQFj6eBnEX31aFMB6VBPjKqpXK7Yt7VqDSVH7XQTaVx3zSARUgi3GzbQ2D9UE4pQ
2SrVyeeIKsNMb/yM5mjYYELTVCs1wMwFyVMix0+iPngmmTQRsFlaNzBjbXYOVwnKPb+su4iwzriF
bq4JItt02skkjzil1QShv8TkimVsdNEBYNGCmBtUvjK5Ovz0bxF3Ubj0MC63D0mPDJkEcgmaQiAp
ItvQs6Osdik+YZ/EUmR8lpOcHv5yKccRKc1tVwsYZaisg+r3dO09aFgBl4gKwB+NsjiY5aMJhbag
TzCpHn/xasQTyUd93jGoctPY9n2qEoFoe3NTQHqD5CtaqH0JugfNzyRy+1fKoJ5fJ+cbohO94g5n
lij5NSW6x/JGgRUT9x04crxhcRb8f5Gg7scEqaC0BAoP3uwN5A7ME8Va+z8Ge0DVKxWZJ14tkV33
94EzbQgZRx3Ne16iWsfjqt4XPB3jw4UuRWmU6xziyHVgQsVnMl4JRrKSm5kE/VkavOjrPWweAhhW
pgBiguDH+6WLMa/BPvATcD8kk59AZtVM2G2yAcdi/0uCSu2oaPxB6S4gwBe91pDcJgy8EbK4s/AP
Imkv1q8xIp61gOZZcnBzz8QGJBfBw6eaGOYYaxIC+4/YNraDgYCPaZWG3Y24DfU05zTaQ/TklDp/
EMNKPQy+O7o1MBiN3i2mepJ4n1raXyalMrS//9VEAl9RNCsGREI54bRwGJDg11PwQhlqNrCxKaXb
LSuZ6xeJYMtDteIS41u5kmlBfHRgXnw26+TJK4gCFJrPLVWHq7+MuRWJbO4JCWbhRYj7kKrvVrbA
9hjjJaFdHfeEzeHR3/xgurD+nHtko4FsThT27nbx8X2+UtheXEhk1MfoyuPEe5EqOkws9rgxqK4L
GKiLG/6sJqxboS3a/MV4ZdEQTPI+8GsZQ14MV5VAscW0sZf9P2w/6CkUcaHgJPpzYxFIRhFAj2a/
dn75+WA9+vxF0EdVplvrMNt6Upz5LkXG69BCHJdBrspaOObz5ZTPHNVqltBNIzTSMFO8H7y0r6BN
CMcclCpqT7hsa6rg99AInAP71r2bx51GT/htVw6ualIivzVii2bffFMwQpqICcBd398N+tHfDw7c
gO74rasR18UOCl0DvuklJyqs8tpM6oP/uZvwvrwYcCP+UXh1wO3xaueyq5cER/y5fwj+Za17D5os
SbtkQWN/Bmmo/qSYJeAcvoUR4BYTEuZDltP9/81TrY4nby/q+3lLBH9emPw3wo63Cw+f0wexdnJw
IjfC/VQ38RWX5iO1ndA4K94brh4YzyRbhxfJBX37E37/HWdUDJximOpnEbCaLLyvJTCQcumJtYt6
PpuCeGRlGcmMueYzU86TT4Fna6FBM6MT+83sl++z2o+TMT0rZTY3zEfkUjSQ4eRsWetP2SEVRO1Y
sBZ4twYH699rfiwoPJLf6wTh3Nnft0oIk6qtmVMkbGZ8ZsQ7bzw/+4QzGdtq6yUr3YDLWxDNANXI
ldISggXsbwJYoerYaPktWRH5wHRurv5HweCsRgBuFm00GUgAwAFSm72lgjEfA5y4d1czliotLLX+
WiHAMubM0pUAHhnVv9flvpTRIeSw89ZsxowqnyubozhGx7c2tQivzSy64xSuJn0G+8arSt6NB+Oo
/M7E3ZBKSjYp+riYATz3Wm9kp4enuJYT9GAdyRCaA6Dm8xxx3UmVV04dTU9BbCWNjzXIgrn5b40T
q6ufihaTVt2GoXDHQqWO9Xdo/hrV3hOvCrxoMn8Ld4hIpV8iAjfiLRxaPCyNV1y4N9oe6wIKG6TZ
QTtAQ6I4OL3x47WsulSDA703IF3H3r40FeNGdGdg4MfQ1Dy6AU0UDXzVdlqczXA6w2ahcB0a5Wur
xkRQ1hFZLVJ5AzLCWPeQ5Eg94QcjJrX97FoNkfcP07sGIbBUHH5MgpwUIUXjiYl2vW3DSC/b2C37
Ex7/rP/XXGbxEs260pFgu++ZwyvbqW3epc4xDCWEhLkbunf9G03iOhhsh3G+lgPLwUKcKgtEEJUj
xdSm9tXIEyOwj5KPwf3vw3ru8gc12wt67GwNIjq8I/yjSFcXwWNCWVG/EqGr2BWVNIsd35AWbXCf
aWr3i0tUp2CCydX8ye2SdDMK8v5v4F6dgonJqIJpvNKJkgtUC+1pJsKOh+t4VQPD4tzzuNi7AaIK
neTGUaWK1WkarX3ErCV1NPXgTjCS7ptMcCdDk4hVQEvPVkpxtHAcVcx351EnEwxYA/QrSHDgnwVO
ylkcsraJKfEYZ3WPVW6tuWYi8G59c0ioL8/aCLgxXq3W9g/CDlOXJRjd+VCbjHOFaXUNVMaVXkrm
B9afd1y5Kl+9F013tgopRJKdPe++grH9o+zEBz5/DXfj5wkJsuuXBAZC7UPgG2jx3EXUAvhSxrHA
6OOKRJWjW/NlLW8yzpKCLxw1X8+GyN1ZTnvj02hmNo6/iLRJFvov/jwzG1akdNJrhaVYQvPwYLg+
uExkkMC19KYD4gszAiMzbm6PedCCuMwlVLt6U0dXCxasrx4uYIbN3wDyL6BX04Z5HXnFjWhDkLC7
eRLCSoQgcYUsKQcBo1MOKZtj/Q5gU4fyrBXaTUzasq3kBNTYGf976GXNBkETHrhDTBY7r8wwgwqD
BHC2euJisso3sVmsh5MGKoepsx8G4erzdpVGoxu+7bL2Goo7OcVom2kL/kv0OcLa69H89L1kQlqk
qCwTZBUs+5awJxpsBsU9YMgCSUud5A8hpdv9665yy/RGqYyLOMXLz+69mBIGu3als4Gcz57iuAiJ
AeGBgxr1EU6F+BQDmYt8dqgjw5nIvOpK+gQMdFI7Z53Z/bSaiD3GmMUyzx2gjiqY9Qw/SPUlvpcR
jEGtvmDZqeQwPJx3XJaMIl6bl+cZlk1jqp/emFaeUQtx1YHIW033KuEVkskEHP1he1MqSrsdGhsT
aNkOy8k0rrtKOe0BoQmb7oKD1Jbv72TdZIVs0sKroai9jKEVMLfoqp83FIsWLwuzTIUj5Y44hWZ7
JxlbebZkoGCCv6wNQsvT9KO/g5rv7cR8ffE6gWrES8jfZvKdQEPcS84BxNakAwYC1u1vaBvXCoEe
5eVoL0ehC3LXGZwoKVfG6/P/SH06PE7A7G/xEgFoo8TboviWGs7odxMzVbT7uqrOBjDYtzWrDu5s
TjTuNK4ly7TxQT0+2Pdzirt9RFcFPsq6PVR24An4S4PvIGCX6mwhIvYXEJqbGzJeSxTOA3PIQOEj
DK/aBm9/yKM44LmkgeKVW3XdL2pl34mjYf9Te3wfBSmT6TCPRWp9juP82tTvw9zfCN9alsr9V/6l
irXSTmX9g7tbYYAzvfvoQz/cjDxn32xvtpHcr+ttUWS+raypBxlRO/Lj7yJQ3npp3JEjEcdNKcws
VwcGW79G12hOJVLRUJQ/6vzO+uICC0L3tx2eK0J4H8I/vyDcHT33t4mls88cVlbcFUpPLr5T2B0m
4ZlWt7Q4GKeRJrDDGs5q+8Po7nd1IsJPEtKk4mBX1eSGC7P7oYt1NRXkjmEWlgjeZ2kJe+mqzcEt
89hqVwIa9B1N4XY8B/RoVRz3KCr8fb4KPTeA+QmnMB5iQ4AfN5UcCWM8s7JQYNzcVpA5DkZJj3nK
Vt0zcsqXm1WaTVRUeyJrnWFDPd8FBWl/i+k4CTC06cf8mxxzHq+wyTcPrV5nlup0c+WdK57j1R8P
UroxayuHRlNyotzEVNBvkogB7g76UFf8BStekyr3qvm3cQyIQueToytGwHwjbz3Dz1cZjKTJaflW
XJHVWCy1brtLczSDA3NRwryaNjm4bFSmMPoPrpzYWtRwbe6MVnLByh+KmWyIRsVgvhjQbMNx0F9d
4xXMWVUCtif7hB4QzQK5d77s6CI38/nkm4S7csGg3b/7Czh6c+xFS15m4yANzlLUo4lQ9CgLd1ZN
0P10v1olfswegICw5jq7T9wPoyClCorzWfYieXjXY9pSlk1iwZDMsSuPWpoIPut9+YoDR5jsQPsJ
FTNnrm6Xt3sqzr4tzkAenpAyYY2FhyHAwoi2PbL4FRVMiHjMs730qtBREhbOQ/75/m2yWssTzpBM
Yg76gqxoUYRrnsnFqNtOanZQ7jaL8eUazC4adsuztdMV8Z98tBCCx2HgFKdVHNaN907UVT0le2HV
irZO4SRA/yqtf3HisJeAunH3/MF2vmtBrO+N8w0kVWCsh7Wgg+kg/I1+UAMVbWgtz+jk5H8KPACp
yZ/7Ec9wKcebpEK/ffFNualWSaGDAYqDFHiti3aeT6POn6jgmpmPe6ZQ/z45dbW7uM7OrxiglhrZ
u7jy0b6YzlUcNU2it/JCKw1WanpAeGrJhR44gvki0ANjltsQYeT/4dFW/vl0yS38IocAzOkj0rGG
1X9L6DKiGRy1cEh5llKKWUYToDye1HiHpPeQzU3fV3nYYPRRknffdS+ECBs4b2TZYSGYKzQxJ1sr
aiC9t2ixqEQv0XatwK2rindJ4YuunoCL9ucH1xRnhLDrXsNBk3cUwSCIFR3xHAGa015KE0siNN6u
mcN+5TBSkc2899ygnrQtHJlk5o/KDEEx7nAh6q2isavWeNivmpAa5BclpX4ZisHk5BObWpWsx8AW
cARqZ83rP14MIqzosT6jwfewuz7tDuCvg17ZN+vkebdN4qSzOExKDIyvLt6CMfFoQc8U5h/AiBNO
cZDDpNyqqK8jWsb+YECOHt+t6BUZzHsFVIOozUmptQZy6nec4aXItLjMsVkcOn6xqMWuKlu6kQcQ
BQTr5gYMhjK7/wCAh3NiFbHuADJWso850KJjXicsHKdFEPGu3xmWN/Un2BUHpFKXvX1eiDGMl2We
uUTxn58idSsjljpukcJPLziVkE0XZ9CdNWa3uhELjlj6iCQZApaOhf9ljM7Ih0jIq6HgskDg8X/L
+Ivl89pM4XlnnSQw2z6+3d7/BqD2smAkE/7p5GyhHOXNcPHT/DEzs1RbOZpXSTX5FVBwL8PtKd7k
Xzw2KPiN9kG4kRFcl/DQ2j7+isOZcdOiEJrAD5FwA4JptkXxuKsVAGlLYJ9hHUCoJMI4R8e3+Cuc
K7CfgWYD+xyOBfeeTusbSmzeqLh+hrqoDjO2yjxJIfb4hNUC7eKP/xZP/p2RXaDJF4CZnWGVX+vt
VvxbtwYglHKxT6QbitJyCpUdwq8E9cLselc8JFG3rPN+oW6dSv8JRyltB6hJNElJ1DdtkyMrp8yy
4I+67xd7aNSMvXlLG9vAl4E/TMAZIR2YY6sLxfdxqJaqNI1QeBpX+P9wZ/rZPJXHPFr5No3dnQbk
KQviLa+vc6VWU+8ggOwe9/PoLh8s5yh5kX2HS47ZWMJ3MVsoAn4WZ3AX62bmZLykSgj7Ec9+Yar6
EFPa6Nw3Wv4h1hN239hFsXdzPmb95M85si3HHjmjQqdDlqdXPoXQ577vJde/JHx/tiSWasrXh4Zy
7gv576Qaw6PIaElL70qk3pc+/8gvgWWsvaAoaGaVHofw35L9kAFD0kyUjM+qZM7S6vp/Z9GQD55J
WKKTdB5KxzZ3yNo+GcUcv5WazxW+uAQW/HDjb8H00SiTuaov5TnD2R9btL/Rbx+yAdQoGq61+kzx
fLTaBKnCppItIcbWXVsXWe2ytRw+3itCRzbKArSssjOcbc99XZIJ0b+jXXn4uYEtj7uzC+wec1Jn
IeSWfYYXOwrOa2NXk1xjcbF7FUUxsHqmWCKBHqZGFHYIf1yDM7PbZad2FILd6jeyDvoFxTxAhg1U
ZW0JZXjnVuWwfjLNlT+pTpgJbGbNIdvZ12xyjwWvudhtzJS3l8VpwTee450VcnU6OZbI+GvEVEdW
Y9h7PO1ge4TvmgWzLQ9fIFuf4Xk/Itdzz6Wq3ULm7pAmssHiUiFQjzpeCRLm5fFnzQySW3Y+6In3
Fv4zYnSDxz4PHWluaumPUMivb5msftFkWt3nMdG6+BX7fIS5iwe/prqG8yDryQPrzi8gWBQRw5/9
zyNgyg53jpg+WfIAnJRxNTQwPc/FgCNnOPxJnfA6vZyC/nC1d/jkwJ3Ffr7UbsKrrifECJnSZgtG
xKEfKC6jtpwbnbOOE7gDNa6KfiNgKSPOsXwWwp+x1vLQmfGL3j8MMzJxZOzQJCFueC8u7xzYdktv
04u6uYv9eJGke/Q7B6VznFWyAZMfgfLQxGXnLeB+Pc/nxQT0e/+AYRsrHoakW2lSvOaya8A8o9P3
r/+cjIhD4nBWagNCU+j188YPz18f8qfn0ag/Cw6UCvIb1PUYbFnybwJwNNB4fdFdw89udQEFEkKQ
aR37pO76ax4tzUSR2UBc+3gb0KItTWUc95/zHOY3uIOVQBRGmMoHJ2Y3zqe6Qf1YVh8VYPAK82JG
tsMoWjkvXJ3lPHE/c84ybprd22K6shk7Y5E+kc4dTpH2hnhm7Sg5mhwgKvbDb10Dgngi6NhahcNU
XUJE/gxn8p+bBsop3TByFH79L5nB4kw/8MR77iiDTRCElzTEVqqZb6yMYsFAuwmgrcCZmJzqb8rP
80NwAwPmcqXmtmou/p9l27zWu7/ZQ6NSJSbu2xTnk1a5+03KYkYgTamfuGSgvl2XHP9LJZ4uujjS
CA42eDOT2uhoUWPRqQWtEdv8EDY/uBQHd60FSnLvknQUYosyDUYwpqDAAgPIyBaKxn+wS50Sc8sc
EqS6SUXJPhhx1i4jQcxwbnx3/fb+bQ1WUZYzaKOboIFFIordj6mkP5UvV+hKfZhuvfE8ib/8pXrg
/GpH7EOcT3OUOkDbrMcYs/PFVLhXs7Tn0JFthKhcgJMeV1BXB084Xyl3VGaiFsa515S2TN/9NuHq
9uu9lWyzukeKDSaTqWvVVSGrTvAvkPxib76qS+Q2T0xy15VJg2uOOuIh5rjPtVyuiAaiCVW6GYqj
yWfPVZZNMKdYM7j9svMhv8+MCPm9tXFejoHsfhKoIBvb+FV2CrAeqT31c4mqoWqAXqWy0uitWJu2
IZoGJqoN3ntDSK5YMHETFg9Oeb4T6mwsf6TAuOf74Kp5+GnV/C+3Zk4Y2MQbBERwkXlk0wWaue3q
d0nVgvD5W/V98Xyp6kp5sz7RLbFiynJmXIe7QE1Ex7D/z2HFMjU4AG0SeODljAftcn+Wrhlevrk2
1jNwlWY4qoZn0s4NTbdrJdTn9RNtMVGoFCKFUYvJNQ2xsbzISIXkoMLX1efW3QpDvkHb6Uk1CDEq
SgmurpsJoENiBmYoYETg99c+SVGojqaLPqYlVcFaThm2f8MJspVhrGwcI22LAaxOyf7d0JCuzfh+
1ITc3jXh6fE4FMovQdxGCv5ZcxXMcedcCf4D1mcqXEs/+Wv5c4/ns6PDQkDL/dWAhO6NonKmGTvY
Y1PDTRxrV4eETWbMFpmCnzYmwGogIGc/8AQh6sxkPAtDjbLR58eNccOrQoijTlUKUruzbHMfcrvc
imW/IzWdPwfz5Vd8Evypduy+m386u7Ev+LKd2LhEaMOWnHJBRtb78g7iO7nKTfWODF1UvDTMvxXE
Jj2XIEivdai9nJJoIncecxgk/rDp+Jixu1abxoX1eaJ38EWNawJqWeq60HenMg+HGKK+naQfCfEE
ra9LjkZ1CZbBTXyo/RkpkjMqYPcZmag/RM0EvYBndGTL0owE9a+tbXbQsuy5CRbyCAwSTnqr0aeI
ainRyzTcyRW4UlZaJaZIc8ctkMxA26tdvRWuPoug9+yENdckVOGUNRdMyf9dT/+185IgKE6SVtov
XVIpwXT5KvJfZUoKAeLmcXvnG8U1oqoPizLs0XIenDvRVjDHiN4fOniCarbm/jou5EFwncUuJpLN
GAzmXKPj3lBoRXl0YCUU8ISN8fxuq2Za92agJuBTU8TQqDKZnbRR+0XhMharHwBZV4oai5xoRXGU
6y25nn9ipCZa7b+U1uAfFlB3lmFUEUuYFyKi8+3ruJl7e56VMgJ+5vHG36Oel5bpVIzha/09s7TC
VN77rdUmS3iV1cFTFHeSUOvKMtXH14LKJx5ApHIZ6VEBhQkIY5E7rmQ7WKg11b1Z18wpXMOEvFhd
WZVcyQXTmwRBtBnTP59w9JrSeSY/Zjp2SlrTyNgHGKQ15gZmlWl4MjKHgvlT4pDXITbww9f90dod
6tKE9OrvlW2VgGqe9kSrY6lmbMCD6Vug5foc+j5E3CUaMuz3mZMd4Wh/+vKpef+G+MlZbYdSCflK
983v2xh/+huW1OsJa2+0i4sCs110ixBYok8g2oZWr12o7QqBXzX+t+hqtKbvuq96eb9eqKJ7GiCb
zvgRJLltFHTB39FTQQDkLZqmHtbUw/yW4MeRvCwcJGxm6N99kDOq8dbgxC2MXDrj/z56ZHbdIzqu
/oLfAApDz5pQtJeztN6wQe8LQPRIKrrbO17dswousuRDQWGnD6Xt3uZ+7N57sIP6Tvol9dvg99nF
PdNN940/bReabiEKE9Bheu3cQRaccHuQPiCuIpUr4mi/lYCZ+I+8AAJ05dXVL/R+6W6FQc6Vwrci
Ba7BrmX101xvBhIbmdWVMGJz/UDAnzjvLqWrBrbRWTwBkQ5VA4BDstOB9IAnPvNnYldG1YgDMgKU
IdHrnriuUxx3nrupsNPtrGkASvgYRBnwSh4eTsj6taPREIjjJQAo7LXcvZ1lAIhR0MOOWLSL8lgt
w/cAt+bs4RynLF9/MUee07QTb7utlkqq7adgYRG/Gzh7eJyIkPDan+BG97f/rX3QVGkuBIQMBuHN
PdFvHu18l0jlLKWydZH5Kvps0Lu7Dz+k4Tbh60lrJSZNda/SUqvQrbL7TbI6N0GroIfLIOPUT16K
oiLlyosB/Hpmv0wmcgA5GgeGffbG8EahQd2IpohpzjzAdXxSHGfX04qSjxyMsqlnGlhmPFKrbqJx
HZ9LBwhZ5O773hU+r4y4Aa6tws9j0rQViM+dqZ8jxBldErD+/kYtjwIT2pAvaaRTTF73oES5alg2
ekzrP9O+PhVpkNYcI8DlnVlhEPszMmCIoev5dWf9Loi7o2rYKaDxPMv8smRRZBaTz+OFL9osQl1U
JhfS6rUIunSmN6JObXTcSI75ZH3NMAjFUOY8J1stZ4hp6FZRuG9X7E81f9rCm7+Bhc/Cs5uklONp
3uSmX7HbBmL8WD/J7tSIs7E8SBGBLxW/VsWTM9Pgv1o8ThshbbmItwz64mbGDqlMASpBw8VQTHrn
z3F3yjpv+Ctsg8ywOqHhKAyLAboBpeYeK7BVbZ6qJ/STrjIrA+sCMqwp9YU9pHHUDMUlqc31WYzs
UuleJ5CxSGOjjJYgQ7OUqMlyoCvwbl+1Rl5QrLp4hPemwiAVnk7sRE599+tjz8Gxbz+NTKM9uG+n
Pw/8fDFfJDSuVU17NA30j7u7QKCoTz6FkNva50xRXHqttXf0Jj57KaMRDTSAFGqSmfiG24RA7gOO
rGmX/KDtchz7OE+cF6N1Co0c5Q8S9tQxSgJgSU4FkXO43HHAA1wUcCGbXTXl87pBfB9gLn7oAK4J
ay4QyeL62132p9Gu5rZFJS8Ptn7fieWj6d7Ui01nGFsAaatt7wBUZld5ZHvliL9M7rSbo79B3ZZS
sbzKTGW+6cNMSevp17ckYkLE0jWa+1MVcdd0jOZnTKjAUDgzO8lX4SHgMcb2sA/Fas8O9P8h9TqR
CwrMzYG5XfYffY97sazbVOQozOZelNv+C2Y3RyjZQdrQ9qNWP0eNF1wjdOZFsIXYO1GNUyJ6v+jc
9xbQXAdR+z5GIZZKqeQ8UxlLEn1WZmWS2BivCwYoLNEWO4LzJLP1/KUamXerDzMb0GSzXIEuNyXV
6n7nqMhAhV+0+1P9Gs9vo5jW/AnrPnmqeygaDrywDBmJpHWcwqCBThSzrdwaudjEQVmHtaTij2vG
Mb4lP6HBNwoVAR6RocfREkq7EaLslJ5Eac6QCOCvrTa5EXwUn8WyD2QOSAiNPEn76fiEcYbV9TU7
fuqG0U+mEg1i7KKuHq9Ko/pnU/33TShIU5SW6ry0qOM3gVWGXqTaNb8VqztXI4kT14TFvPto6fQX
UXCPwasq1+TVmo1e/uQEVpiA/Q5TYzeMK+UAtgQC9vpmH/euu3rdcdfvfxyMZofIWQRGz/oQW7x8
zK1zjU+B6HRrD4IBE2LrIZWTDZOYT7vmfp9IaosPHOeMZ2VDU+kVux3JIN/M2ZkQb+r+cOpSCocA
3iGJR7PpEJi16K0e7O6gkqpiNpKgE3K/0EAi065i+9fFqs0E+TrP0EgZfasFOU15wQu4+C5vLVvt
w2jOKErAQSXv7c3IauAepO18z0mff03y8H3YGXYyQXLT8r5UD8QNBrJkwog0XOAAllzAHuR3/BEu
Av+8XX6UrcjuILDmwNyhm0yedUcxOhlZqFCKdjxcWKDEBet0eEbjXLAhsN0QlxY9in6k2FPRPqp7
w/l52auIOIBJ67wK4NENZMtCbZYCJfHKL9rBCbX6Ew8R8zdbc8i+r+7Hwv7wSuwsD/1sbqu/AHK3
AV+eiIjq8MY5Fb7uebkh0cL2XV+tvDJvSFf3XoF/e1QpZrtCGs1uSgBwC6Tl0Z79WXDZY04BkD5W
dc/mlAl/sBt2fs8ga7hKIVtmScvkkFoqReZp3eUCdElRqKKo8+Knq6SsG5AmVf8jBg+ovR4s8R5J
eeeOgBFE+7f17D+3kbAjjerXuzR4qRKxwKwXjXc7Ql9MTtLFtx65DwUb+rmX70wS3zIq1FWigHXZ
rVZhKVfc5kg/pz9GTDbr2T/Xub2dytuorQ027I1FARerdsIwC+z7h/h3pbGgcjbqtHL/IGrwPMp6
BGau4deu4yEgzxlPNw0ILuz78Q6SeBAd3/Nohqg96GA8N97OUmhsZKM51nU84IYOSXRu3ckfKhrw
/OsSo1cvdkwWurADx5V7UfoKCVr34Y7uMCGJcfXGHZ7BBT7pjTeW5BXSPTQU0X7T+Q3/A9hTpAop
eF4p98+VzXZUThCSw28eCV26/3Jpy+0wq/sIVU31aAMgbTE7vhkZvfYentvb69GRPU+HHoMqVj4s
nz1dYGA6GiZ14NX9YhzkiEU9z5ZK8pehKcmDPvmEOybKFWGpKfh2l2EYLTZuay6firFlgkepPj51
YpNVSCEb2o6XxPTc9mHGrDvdzTED8RwekNg8Qv8Qf4MCB6122mqrRSE3zzI+87DXxDqoG601GG/i
qua85xyJAByDBW5tUun1jwJVjbh9C706q/RG94qKtWE/kIQnbM94h3HfwDnOt2EG3i+vjJSH9/9b
XofFfGFuZVeST5+Mae+jNZF1RUu9j8/C9drpgI92R5dAW391HQh5n/gvVJZ76ps+QSP7IWqKfifZ
NzW+RHZ55sXbD3gb0y2us+XeeHcAD8B83UqRKr5aRToYxC5ojYqbyx5CaTac1vs2R4dWDE2vbqbs
iAm+/PkA/v2jugiz5x5nhozw2DoKHMy0szuD+PkWpxKaopBcBXmh7wdaC/83MzqAsAKEeuZrzFXV
DNR4Kss9jcYhmbOKYaHEvzOuvdnJwW6QH6ACsph1hUKxzsF2lleqEedWa9igdjYRi6d24lvChEl4
Y3z3foXoJvjcMAMmLFiJFk+iic3cg7+MUiq5lD9UzahcNVSjVtyl3cfHr6WiLEiHy4+dxw6AyWz/
GLSJ5v/dTPypKj66LkL7LJ2ZYCi4uvULR14RdNWoL9ZJnyJlguuiavDdyABHa6S6E/mavhPWRiQN
LmujpMLZIuI+IIOIO81eZbvmGE01EaRrOM5xx+dQogLNRcMwWHIePOe6/UwneJatXXIempkqrHdi
iB1XUIG7fAnwZ4D5AEy0GUyCBpZU9SNdlQmI93YKz8uUCjoRyMRBEAD9mlUXIwhCUiljN7+afsIb
MzYoLbSu2QSE7in80O5oLJzSZNmLGPKnOjs83zAiMWGs2lCsDoktoh6n/mQx0YYkjJrf9jbCV4zG
GxVJswP7aVA3dcDZxOgTOkT9VeX+iAKEASgOejTvXy27ynKNXodRrUu2zrjt3XlPOe0EqQKJ9vMr
zUdkA7SJBZ5au7ynL2lsXUqxXe0+mCgZ2UTnGqKzplRJ0nNQ4btzKrul/QYRuseG9gZXIZjVGLNO
Ex12ibU/ytY8AigcQ3UxOlLbCpnVV+Av9NqdYKNkTyJPjdOBsjIDpr4F7gV4eVFGkDZVTEx/LQhu
8OVnngprABqKFHPumlvuZFNDkvdFMhunw4Iw547AQuz8BrkSPZWd1nHXSTwc/TFt1baqu4tRF0Ik
e8nQxlsFI//ShG8YSBUGUvb+PD1o33hFNs2xrdmXwKWyjGwTyc26OD8Rt9gPC8tGFgpWeYyJ0XyI
dmBLXJZlrYQdV/4+GN/kW70f30wxCFZBehE34WwD1gE7NDVas+mbSgcTT4eNQ43DFFGaIrV8UtWC
6E6NNBjb5+g+7kvIr+cbjoQO5fO+RmtS5l0pSAHnerp61HKR7cKC7a+UxWoyP7J1h2yhl8bQrvz1
fqTXqba4Vby5Xa5kh8ZajM1iicDC+hWqFBjFZexjfuwUCRf3ZiDlIWv910B6mZisAjA4+B9etYM2
GDiLBkGtL9uyZ2wXVF0G6Qljj5CWpCdqSD/qL8+OnfNxIWM1nHqE0rKo6A+dVwHXWP/+fyY5Nsoi
/yfvaeXZe0DbV1kdHdmF5/Gm7Vkug8zvbi/2wkYXfLojHSfCOXMjI0J0lkwij/3TrZfSlqJBeQen
c6Nlv4N+/w/gmui3Ddt2IgBGNnViCHntFh3ePpmZQtYUafvYIPRGM95OVqBli8QK0rNcn/Tbug8q
8ko/oLlz7xBAOQyxZ2taKX0dj5KwybleNGP9PKe7WJ4A1aV2heovzTzH9xK231wbGELdy5Wntg9K
CsdRmd1AIx2ErXH+s0rmL6dux5rgHtyBa2y/55OpNCAfJeo0OPCCwGJNF7uou2tSdyruF7S86E81
fO+qWdhvrd1MKoDd9UUGJi9fGV4DwD1GGQyZgO25YhBLlOdMBQAbov18R6nG+2yfKyd/RcCBY67F
R+Ey7B3mcZaNhL1Q6MDMVanGio8o93AzNkr6ehXHLXZYXBxZWtq8y1WnsmA1Bd0CY4Wz11gnzXsZ
bJoDRFusRz0BuDene2lsf/hrAVhmww30c0t2aW/3l8RQ02tH5W55fiz6gR1bcgDgKYdetFyHvog9
e+UZD+qw5JQUVgBWEcR+zmH4SxegpZYci6Dyasu72Uu8o/XiTUVz7Iv/sVdyAcqx68kVj07rIWjp
YzROjkEcWT9D9NVtTbap05cfsvCKTZ26y/Wwo9TsmZTfZc/aCxcIrE/EG6gEFz+llg25GF/GHATo
EQSY06z3gmmjI1/U8zb9JmSfoltVDAfSDgwPQKToED+1xaIXIsBbRyic7SbZKb9mNg/l7FTcHY2I
/gl6FSWvSAT0iFD8HlY21n/fY6yclzDmfF9+6LMgpz2vfbZUGbkFIvAWNvymxAiqOTPoHj5cIs6B
UFRgiR7iLBpCjUU3TKj2imqK8kOle/ROChxJpntaLxIOkG5620PYrYbAejHuNNLGPQuItax3xnvI
VP3LM109xCRRE07iIf1lic84Iduyej3OHc9F3jxsfomcE1z/EHWmVYUExkG5x6HtgRy2VjZpA20v
aTLMyQy6FOr8JxUDDfehCeWJte2URmV9bWti3kPHOC5piX3eNmC31Oxs/qcNe4bcpj81JCCXpwkj
geQbZHaKTPnkIYPZwhk/+xiMqOkLAqOTnlKPut+5pC0715JBpZQAxl9PRk8I5+wdebpJwYAwCFZL
BzGoJ3hhcW4JOjjxKXCjmD8CM9rdKsDTLW/9FN2lXPMIaMK4yO7xR5Ksy+gxqe+Zukjwn07Y1SUa
X0get1Oi7mxxMHnJXGEgPGly5TMgmhe1Jtf8jzBZVT+4/9wwy3q9JO90K9y5hTl1gmqvt5WRmS0U
kM19f+JVCNTVIElGJOmXQqKAulQAHWLyRqTMtS44qb3wMnK+cIyNH7E0mvlG5YT7Lg/OsG0iV99x
vJavZNk4Ewju0253Q4I2sAUiY0AGLodv4/cLeHc+dyj1Cp3HAO8dz1nDSOeWuLN+hWjPNAVGbq5k
rKC/ESfkInUHmURc+ijnv+0rqh62xIh9Kl/P955qRMDxZWAWAG32rIENzsc5WS4Ae7gBVVKvXSzF
94s+oDoZnbrcxThi5+01JM+KUKB2kMbFlMUNbvo0g6Mi5KwqKJnPc6stK+nn5b7AZfNJh+f1owcN
i2MkX+VesyPcgCqSAcflPsNMLZOYksskYJA6ateM+nz2IvNpz5UWKIfKyAferPyOFRh6Mm59MpJZ
km55sYHQR6FtJ7OtinBCg4dVPGNhqUOUB9s+QYUjXyvCtg0qHr6oG1DINkQmgzFu2KvsBT/zes9a
g8Eh8RLHxB12GEXZ98gpxGmKZuGkYmNsY7YNe1KP+bHenCWEZJJcLpIuWc9wVoSwJXjrkGsqEniv
/0RJ32NKJv1w4HoBR8teXEVMsAAf5Nwv3/SYaP6+znTRvh8AJx8BOZPtvgi6g57xyoFNb5L3yTRH
NyRGlDdd8C7tQXgFGNRiLFzp/nFONCHeC6KuPJzd4iDDPepVzFd5PKjNWoahmZIVHtUon28WDp+J
mqAJPNREO803f4j1Q1TzHHHuBlu2NkrenNIHpnU4zFfl2UP7Sc77A3wWdfnCPC4La6qTR1iDjw8b
HyupGmDMVkWwEbAxxgeb897mcCtrG5NJ7vfLvAJJg0YuCSW6HbOJAlfBW5zsz9dt4xCPdudU9fOZ
9KyuJaTXqNZy6mPZsTKTFlcvimb4Ma9Jw1HbTbT/FY5mSsjVkqc0Ihw8VZks5F4FSrN8cK5IQDsE
hpD/qQZGFA7aWIAeitECgza0oohYPceXuMVjEUL4U+zpXq2mpT9uERndoVoGsuaflY2qx1xL/qI5
PTfzgPEkj+IZuIbTID7Lc7as1wuyeuu9+f9/9PTv8zgJYVWPKtMao0PkcquBNlhtHZddGUvDKGf9
OkU9mEtjoF5burNaBdP3k4WI6ltfNOHQW/Hm5qZUTGq6GQpuZzPngtWGHbhAh/S6oAkafqwYugn4
QM9rjLU0fSfdnAA/IbXbYkHWXqwcRgOybICOp9mnZQUxuXZT96DGE61X3xoNvb6iJ96oT4TGuhTk
hatPFBEnAFBNXAsfIcxMRcyk2kRVJN6fevojReoutqzT5HUpP5IWmYKp+Hi+Ejbq0FYEY23seAE0
5D9t6Nc/7/zmz0Uh6HqAT2ICW7C1rFrs2hrsgr8fEdZ5lUotlxoKFMUuPa1O9Fmg7YMaWBlSDLX4
Qs/nfRguFKXCh3n/Ol8DdP7oDzT6JG+PxWioAah8sLhocmkK9xZLVB3n5KAkEZvYDOxCnA8UD5cQ
rYo6RWEwEHA43BYDIwN2O2OE5l4ruWkIoOSUZFffdcI9wil2Zg9ioTUzgiZmifETJnKyc/w7VYzm
eqVm6d7V+TUkTB878AefSVUMQxNCuO1bxvX997nBDKg/8nlTv24Oyz2l4NR3fb6pYQBE0B80/Ds2
L8Zh8F0XFJC5FLJnW2guccMRJAh5/5q6rbMZzIWbT4y42GkgQR+Rg76+12I9I3lm3YNkkKbtjkRo
COvUCbOJWKST0hrJ49sWtupG/dTMjFIi2C+RP4yQxC3V4QM9O4qCVq44aHDAU5/wDXXt4o2ysA3m
kbMhm8oiZ3RMYDc9gOLXAeqRZOdhchY5pn706K1O/DCn3Wv0KQC22pTw8+9agf/2mkIIyFDe+1q9
vviKM25nGX5FwaWyzgWEp7xqziPzOgvpdbrDd/6cuQftG9yAT4hU8LXirQMr40yTXsnANYkR5Dw+
R60/kQOu/QHnSPgaa/3/xqnlqnQimv2u1r7WV2KlbHVeQ4cZRT8RA0cKfO4t8bmtl8hU6TlDQIJq
pStnD4orehA3NlHevB/IksrpmSj5UiuIIOUpr4ss0xYHdwgIs2bpzO/kH3e5zvICyHZMcwospFSy
mto1O4ZzlebBAEYXYz1nbcxSze018bewYCJmLZ+VogweCWY+LFjDk6f00ZbpSaTJhvP/BxeSpgz/
QNMWIrKZxh/ssZSP+Tf0bModR/024lpBPVzxq5+RP4t2p9f3dk8C0hUq08x9G1UC69gQG6WCKQ/o
+c6NPQYFEaJE8Fs84tWJ748TGRn8blr1KzeLx37toBP0sKhc6JiF1il85+ZvlE6lWmSx+OML5dX6
Z7CCX30YtKxDjclo2OEbqzflvfhswGkqzzDSBAlmoI3+BA76UxDSukA0FqZ4MusUKaBN2ueZvyHd
dQj1JfMnuMejosigg6FYeO/AitppfMj/jBcICeGMrH+VbMphysK3/MN+9pfBovZMblKmc2Cl/f6X
ZhyjcGjO0LNyMwX4SQLDjD3xJ3ieQb8eGimZeCcZZEmp7DhlPAKyrGDUrYDTU86nGQ4h7M90Oins
nukH26gLy5+17aPp+Q7b8zkEKyKYQ6V1d51Ht8S4CcyM/3oN+Gt/r9Udn9lX8GQzxbJzUh5gCGev
SQe8VjvhjL+cH3mNKQ3q796H+hMvhDO+ropeAW8MZN35O0V+SvK4Oxhw8w+9rTpPY6J9ZSeP+WNz
FExhO/8snLLtbi5o39zXTs2F/+0jP1NQNwpsZpaum+FdYhw+vylohWq31JN1RbWSlRXCryKKJkB7
06fMBbY5f+JtzSklUX4gbIwRrDgQ9P9Z3VZjTLGZjb89RUfpkbuPqzHVyhtFbYEtJiSekwYJaT/V
FkpjO/L0LE3Js03R68qDLK/Rrm1QZXKCksxOtwV3/whYuAuHcEieoAOLpqqTuA5x5NzDbU2+KUhU
yDMp8jMT8TTnMSk7SQx3yQFZzi+Jbme9iaxNYSW9jkPQRuG6gSFxd+yKD8EBrBP8lakVI2nfY5mw
VPuv1t4utS9mq8LyRJM/HV+KpokSHNDn8iMF2465/8hTd+ly0DGy3/CphSUAPROqM51+KGi9BYtn
NBLc+Nlo7T+ZBcyp5QsgpYZ1SaUTUEMraI8y/SkJ1Cg6xQX9XvQFkgn6G8Tt1fMjdvCURxsXAwaP
ti0Ouis9stGfZ1qIK+nDWXb+xWV5HuYN7aS+ox+oGXKQ7IzEDlBbMeT7G6e4KoUd1cr0h8KYma8S
LYqqSxP6Z/9UfBJnTLJ4yTEAVGKb7+3bOjNw8gRKoJG9TmHpxf7oIVEiMYxKY6YvdFmYi6187mkr
gMmNPCCxhaZ9ASXkXkec+7cVnnY8H5jc60P6Oc9PbzUnYdPzXUwpe+5UKs9qSNSqs6dIPUl1dLXx
yF/dbHLrHPARB+Slc8v0UQKKnnB8hsUrthhnWMrcWo6J/qH8zWfB37LH5tkF0s++Oax6bkKskU16
g/v6lM6z2lp0ArFRwUYWetend2nReJ4Pp+5dZXywWxPsU0qgjczPfdULIdmkNrSTlPuQ7/2QuNon
2DIRmwEGpgqHpIIKUWDtDI7KO2ns+6VhAuwLONmmZjQdqpwnW7aFufCUvmH29a6brAg1y1ODMtF1
ZvOulQJ+xFdgeMDZs/RLbN4mPD8TTd1F4kkcz5rs54pHYLZJ9BRODSB2fI46ks1YGrjD1+zIFIev
9kU8uyqjqbw7ajQYOYba0Isvnf80IDcKuEbk5JAIHhzPZDc3SVGmVhe6lmiw200AmH7/G1MPhz8X
V5LoNmlit6dtpR+xV6ahQ+E7rl9MmLeOYJMrhiw5nnwfUoBZKD0f1XFO6ZpgdvV9zEhddT7mAUx/
PtBADlg2NE5S7qsI9vaJjjRASsw5SBJFvuYoHKo/DrslsTjuMvLaawnAFfkWgE8z2oUgwNKp6I+f
hquHuIyiGgXQaBE24ZPwgCdSo8SPQ8wGgoFKIeIOo0bITzHmsK4XZmTc5KiSmauVROWXuXs8rQCB
u6FYSQKgdOWfShH6bZPWj6LivEGzN32R2h35tkmUOyTiSY1vEn+T5AAeVu1Oac3ruYYt9Ka9VJj5
VqADBLAI6nO9WOJj0FaHOuyS+l30svannAYZJ7UMI7J3XqfKzfNm6tJR6BBiarKjnDD5cPHoDpIy
d1N7siR1xRkWj4K2OFmL3EunsQDi4RdQ5O9wZ+Vgo3xLIE6YjiRUAhxE72YilqYMvUBonfE0OU/c
FXvCzWVjpMxwGn330Gek3C43FE4+lme0srtjLL19BBmMNlabxl2vDAzAJ5BWD69Bh2CXlu7inwQE
rHWJOerC6XYgx0DcEmJhG2EA8wJMPM3DgIQCJRfBvExtR5xZKdSCNR2nefRqu3msKk/GysR3BY54
Ya/Osbd0Qvy2VPh1sOBKsDQf/AwqQfWgMAUgQfOnWOqZoIowfHDLWEKfttm6OtmOhVpGGosnnsVI
iPrdvWIBoJVfJRCXo8zffJ1rGqT00kQKjesbKxhgxYxwODO4hLNO13bq02YwrHnUlMbzOSueHjIF
5OnkrBZ8D2ZFD8EWCwXoWgaDTwOtd7dvimIyo5gDH3ekDPd7KGNgwh+XqhCGMPcu5TSe0KIUvtTZ
o8vNoaEE9BFPfnl7HnU4AnHzbcrqmi6UF0KVBRJiUFyFH5lxCv8NKymIIrYIxiGP+W6XxvWFjYOu
nL46UT/a+WJbozwTKeI2Rxa1ovwjOkstXBrlJdh2bcGtO4rw4PLJBJ7udYiE7f3nlQJ4n1kv10hd
MlciFV2IufA7O9D2vwn3hcpWveXciLJ9mwR//9priICBujHd2o2zHhlKCrsXEj6tFdTArTe4X0Kf
E9fvn3JkJbuIdy/OUNaHcUbw2PnOGkvNuCdv8cR2GVpHqJTOpwwN2+sgn7FTiFvFwEEk5zxBeHIV
Pauga0CaWB/wEaZ4lkoqt3ts5I5a1QZM+Q/eA1szRCCfb+Eu7eD/k3yED0S17QKO6rrUx1y5CAPT
lqGinCDxNBHpkTXvyVAOjHubiimsJthKiKIXL+baEpBTxOxc+x2Izp12hufM0iLxK+Mi8wkE2h2d
OZDsDIz7Evhen0m0YOrTrgm0XXXvykYc09xPNAb1KNPe0WwA0M76cYVnxn0CIMrdDoPc/6eno36r
IFYuce9VtF8CJ9IwKssFLkqZiX2tQjRJr3xywEG4TIhBunpfjb3Yt1LeBhtDNtbjwLSHRn4qAnNy
njIrXk3/ZpEzpBtivTapbb8AQxwolbrhzj0ioZ0rBgwNYVMjoTES+U/I1Owmc3NtG9lZSt8OTEcG
rNk5tIu2mj083w3mY97hGABEhXAsXdU9uNHCni5jd/T8MiMm9/YZO1HBxBo1I6uzapO+ZWWtZfDY
zjADEcuznAesbpSg1snw0Q/oz+KwMhL+fQ/Be+St7hoCYMfEL2mbXqaWTwxvBAt73aEIPv8nTx7w
ohETKnyf/cryCDMZKcQsWuzCqyeQhm8vj0usI9Aw5z09n7F+hyrS27ud9gr6Fb3EW1oSMddFWrE6
tB7mXW3iYThJi/WSa3QbkViZ/D8YDVZs6RSLrsfLvPQJz++GVgRboTVwX+/JJuBgAzxzUYwiah9r
4d/HK1lFQD9Hb7cQgRNPOMzkxxKT0tHY59TqmJ3RyiAhPmxNlUUY5tyX2zEPww5lphPPMGGywytq
CDt+7EVHG1so8smW8phY5oVJqSnUG8Jv5qTnWlaU56431K99D8zhPOJEFTBQ6sdFZXGepsnA5r1A
bI1tthXNYag58EoVIrVh0eu174dyqLs6GVGerpPX8AC9DS44+eXD+6I+kGOsLyJjpCZioV1LJCbh
EvznNV3OqKXl0e6TsBZnAG+p9BPvsyUK36h+thloNay1eAxqaMWtyiA+F0vQJVAnByO4ryCHfAGs
5Tmz79loHzsasbZh3/nsH06HWDHrg2rr3OhALIXLM1wnGAHXoAPoTqmMU3FpUCAPzD3MQROHQwM6
s/BQUoHmLXiX/VU32f5/2QpniJJtXzSjsYgox4vjgcIJa+rNE8U1OkIhKxUvSZrrnpTsSev/Ndhr
mB1ADvjhKLKg6+2Z2rcoHt6j1WECdAgzEl27d1cGCm57O+k3lDM0FOapxNK4qAUjFV3BfbodJ3US
EVz6D5JTyo7gW0Km3jGpsnQE2htsPlpMWG6VhhWUIJ5DbVShIY6LmnZ1MyCOaU9xU0Qqmou8xFwB
EJxI34gJmeN5nLHVaYWKS0kg07AN3g19ZOKWHQkrtkgdgO9DTbYjtb+SHS18O2yEvuzB0Yue54T7
65RYijRJM+tyZnv60wY1hmkut0nAhiWIcQwZwIP0nSnt1JiNkTdDkQMHgswP+UYzjIx67cio2Zzn
tfdVbHPzK6JSllm74eBTX9IK9Cz6I0BwjNeU5HYASOMtMhNUXWtlXKu0pABGiKu8UfWLHkhcoJUV
UzoFUwdtPgVwcl8VCxAKBZzWot9qkXYIh1Adp/oN6iv2hOVtkRtQxFYkL37QRhPV4JR8lh9xhz8W
G3tQxa1lAL+zk+gqDE0T/lCZ8la8ORUxIpyWG16zjUsJO9WyGSW/2rzetTMd/NBr0j+TGf7PaITP
xUvxU9WD+PIPhaJZeDFU7Y2mFD9HER/ZB0S/HdGJMqlvQZSOBSjkWHfrt3MB+ISECA76hBNSNm8V
SIPxKIyR97U1TWIwdvNeKgmYVGkzn7WdXN3JRgCnmD4u6hSOF+FL7s4djLbvdjDlN5pqdvrcPc36
q5XyAxDnkw9O6j9Iaznd3+2ZaqkS+6Gh0hF1L1Ln+5IeKNKHT7pvtShkz77gCcRS41co12PL53kc
NpDE3YkQ7dSGYgUuiSV8N0O/uiwbAZb3Q4yWyxneKJ6SHt3wHgJe/jNsKTmcq5YO9pkg6Vr/myuE
F47yt+6PtnVBQtwI/fsjjGGUViffu1vQMSLae239gVBNxnXDusRj+u8kgK2APoY/sIqCtTmJqE85
I/bQlmI+JEs1ZL3yAsZ72zlnuvEQ8I9fyB6dR2XUtqxJa7SjHpahnoeUU0wI2tsYEAemuD/ozu/A
CBRjG9obrQiD1Nu2Lq7JgjsMld+pL63SDR5uw6CMV5HFARnA3mjPKYwSK2gWbSNnN0UI4PcpUKJB
fDxV4iVPrArWtKyNP3yL9lVVy+L27ijFFuOzvT5QIvmefzQPjL8NrPVEgQ7S7dFkDGGfzbRPzQcY
KZXwqT4h0fOYDws7X0oyYryR0E/tTy/+50K6TJtzqXfqRjW9pi/lIhQ2YTvles+dXoHVINyGOyKv
vgB1lVkMz8NPjgwwggYzwdLkBPMFdxoaimyWV3NINq6SBR5wmbAD/NKo+xYpgn1jq3WDDQZqxT3M
yG6eRbbI/X7dmTNUwM9RUFSfQ6GmLXzyMj/N9qGIji15ivqe8RyNXwj7npaaEWXOL7inO+k/Eqp6
vJZjK1Nrq8EzMohXYbayRor72PaBPgwvQh+zRm+FUjk+oRl0DUEyma5VlSgP3+FxP+rVbX4b668w
csdYNnBgFgaFOs6YDwLGgkK+DMzu/IZWb8mp1iPFP+5gEPMAy+CHp4g0MYinFHF/d26bVuKzN4ky
dapBxtF5CI+4NIbe1+yeHlgFcVqdAYUFPvScFTkIUy7/dj/wNOO2ymfMoii6I+6V3dBWIM7GgMmU
W7lOCqyCuB8YbXVQ2xatOqvDW7iF8r4FLjqrxUKXshF5TtpQLR+2IeSrnzka7jgicV09UlslJjXV
MFeWtvSqmEBMr1YDqjibLMiFH+L27f8IAPJBWySXJCxnnWnPOHPpL11LB4WoArbpu49sm9DOxS5U
YhzjdueDYQrsmgbuYW/zsSWOFZLRlWr8Doo34wgIHzXLhrPJBzNQUKvV9QooO4Y/xOxwOJ+tOvpT
qqoW0f0C6BWxC2RdmKm399XgvP+s/f0gP9gQhRAGNtl/uFiu/XmBetaQdOj73bQP1TgdvGp0MJhE
tFwLA7bivj5Mjbnz/WETwLfO7+J7FUH5l/N787ExmfehnRjn8zKyMIlNBY/QMXZLJn0ILClU9gVc
982jT6upPQyKLuu9qgldtKufzm5/qOyg5TEr0NVh58M/NZYHL4/YwtZuUKJcPAPuD7M6zorBmv1G
wOD2bf4cuP5yFIm/6WApc9+2Fe4tl7eY86+oMdZ9xwtrWOMcfIip5pm9ubAjAMTY/vebOdyKcMlB
Z4NmQNBhmmRtoUcb9ekIASZKOdPWFuiCThPf6F5dOi9wQ7oFmFfz5bFMGy/IwCWnohgzC9f8iiV8
7rc50gvTiDjUeyaTw6PKlydCMdLv/49Lr7TgJMCAV/BlDAXctd0MDUJHCSXNhBpfn1K49bCvgQSw
4KveeWzZHSysThYjSbwsCyBEw5PZulKvkMau5WPPTyae/ixTsvJdOvufjB9gDwsuK7gBndvugcq9
JiN2r3xIbb69CofWonFl7wwGxv82vgFRSsiiMAwE18Jxo6T+3WZtM4ys2k+Daq0GwH7fcJstbOnO
3SbLTuBmc+/tby+5HqM2W1ez78uNUuJty333K/LbYEf6hE7U+DfXdfWEmsYFEpY7obGtaBRHykZi
P4Yos42LOJzTBr4gYuRbvfipDsdQfPKQUzJFLJioX9x+HT4vGRGMCj0qLePMrWQu6gj0muRk/Chv
ZEC2QJCoMgHCi+1mw4kUGhltW8oNZhWmpLnLwxXn7S5qojIq/kxnV00jvOsoMit+un1d49waXON2
bmLuUkfVqgLiWsmjhOfdE70sVUhfuKLTv+sUh/MM71Wv/zJCHFObw5ggS2zU2xBlSEPGjNVMwabR
KxbCC4ktorO4W/GTrmx2ECJnidF9UNmxqbTgT7rqwekYtWKpuRnSItOdfOAFXWMTHYiASQzvqmw3
LEkRlhSU3eZRwnI4cyF2hxdI2S4HCn6JMtKsusb6GKKxy+0lvtbQ6iPDIs6zCZDFLbU1j7fiDmcJ
AY0lAH8R/0mwuEKMIUgb7K0jqdjGZP3rBrW+KiYBldPQ4MHuNbptm5O1X4VsN8Y+BGT74mLO55Q/
VNiKIE/wznOLzlegxZUL2JAHP26ZLNbgHhAdziwBYBLRomjKOAPWEJSMsjAe09OIPHFyqXGQvhUS
KQhpcBXaL9zoeZU40ZFMKi4s9QEfk52gReriV0VGO8fx8BqePJF2TfU5NRO6PQs12M5LKdpzn/Zm
V9BHAZIU+KQWT1m3bi3HtY4TyuQKMnkoRrDnLDFeqApxXzGDN0ECcbCr9EuNKANQLDQqofz7y3te
Jy+XpENjpeFfYVCNDMjloRHfqxwfPKAHnplHNhDIvYtQhxaj/BaNfbY776k3esf5KYE7PZyFeOPt
pt75hSfov1b361ynDlcCN/0vQtnQ3ia6K3IAcEP0F2nNLGNCQR5c6wAvNB8Mgvjn0cRfwFvgchr1
d/746Mii4G5N1lfOWkqx2rkshWynvoAL144GEZF/JR+YeJ585doSTdaNTjeJIwAe/EKMM4mSRYj5
ouvqsjKhrf9JTyjK8qYSGimVOhN48FWTf33S/sfLgVcFX4Mes1SedFlZqWL3tBKUltmTZj+OheqR
lHgxv+N+uG/68WedbISFFaGiCbie06R1nxDg2dgMmTk+hPuJJEnpK3bZd/AiemSj9BD50OwDmKbi
anhF+gyXNGmVrcLOOP0YadDefi4gpotuwvE1Ng35qYExypAfE485RwI4/D7xO66WoRC43/BUb7+p
FiXnxKpsYtzOSHBjqhoWS24hJChSZ53inU7guUUgKTnRpnwAUGcY/rfNGyAuQew+EtIX2a7+POcA
dkDcgeI2SGH6A/Z6OaAEqUd1YneFTpvP+NLkCEyjwWgR2nTa1hyGPFQdlt/VFIEFkIy+AY0Ohqdp
2Ig5P4Sd/A6yR0kjLklTxcUtfZRVOtF+cf7GoZ0c95AkcVYrdMhpbOLS8Q4Y3EsJzHeRG9xZZJ84
kvMeMn/gHYFiLjhBvwYAlAwO//IiO2SKjx1/5EPFHH9ciskQYlkSx+2/1+NqDKYT87zYVSD9R+ZT
+XjRyWeKFs/aIDaRilUztiqDZ2exEH3SBbngNNY3jVHcsXoBsw6lrUfptgqAgNHVBzshFEKJWvxB
sSd+ow1P6Aaq9JV+APIJeQ3Rd1OKmK4ZBT4K/md1T7+p6jFIb0DWH5ePkzQDePfr0816MursU8iQ
LHJhY7ArUY/a1JrV4nLwFCgyD7yltgHEFbFvlAfVg53IYOyF53ZZowhxIAvicNBR2kjl7AJlFPpC
xonSpkRNOHkIU23Pws6Aso0+TCk7hUaIiTGK9vAqcqGkE3qM+TXNo+oAszOrNeB12w+amQVzMQuy
+DqFYbBOY+bOcq+KBJp72+1SOHjgv8Ty5ZrA6M2DqvDckGyDTd4TwPJWWWmgbkH2bSIhoWujWP4U
qINrhlovPoTm5geUV759jWyx1LTj0CN0Ll1LwFp++k3eEpzrvqsSaaWMeA6acFakNKubt2KmBse5
WUBIu7K47zvdxkHV56/mp3hxnKR+VWgoD3O9A40UwocDrzfEREhyL8OKZG3tcNSLFH+GtiHxqm/6
P9JauZDdziVZaTJZjwGljAHEpaLr+2jCDqenpwsiqDj0cuVzqTEMrhkgbDN8qRUAuHrsMhWdE+FW
/QTNdlP11PrQCPf3PITsEkc2vJfpRDDnPwicx7xY80M1eUNAeWb7i6EHNVHuuJfG0og095zQ/u+l
Nhjv+bLrQxgGxqaMiVYRvsDXXWRVDN7QKiOa2Lb4kuvUw1zxtNq4RpoZBZry6B/FphocxxXvcHVk
HCxxwy8xRR3CNupNFSnAzfX3DYpr5t7d1+pKzUvaaFPBroyuGsmNUuPYGFn0A3h/yfzJXW2MTS2d
YLK1KiC/Tvg3dWzP/26g/VTBOfNNiOyqeBDFUev/4BWyQKCeDCk4A/LcCOPBaZcP+s2GgPpuCiFC
KF6uPJJbBa9kDzm5Rt0Hf5wnhhJGcTKL8xrQM0c5HFKli+XsXRErPBwNFfkqkRjD4QAup5laSGgu
LkYKVip6MnBy4Ee54CeixF1l6go36wo5M9bdu8BPHiqqRUB0KtABL1K6F8E4T0KDi2Z0jlVug5R2
UfPFPA/0xDP/POlIz/fSdaGYQnICh6+6gRUvK1/PCjuux3zjRftkNg5yce3cvCYEMbL7RlPAs7/x
7DmCvSc5+rX00cG4Vc9uQv8F0892w9UYeRgg45oZ7zsqRh4PZCbolx+Zb3/26GFWrIirDzbliX0A
QQ5Xur6ubK0G169PdOhGku78TZStIbu8FXNQjI6L+mH8L1kZHdfIVHhhz9snRh/kUUSA0hJMfQhr
51XkNpwu+nX1EOgXEQyjDb6dN/LcseBeDQ/1BhZjv70MIRh1Kw6z4u4uiixGVmVsoaxEf1mUGg6x
v9j38btoXvr9AkHIOlrZhnlNGtmEG4/cCl7pi0UqYzX2kwukxc+mveZ8s6BNptjseSzTN8AibeDu
xGd6+bnDCkR3nGv5804ZhYaJ/pm30bn/ZN6APfSLhp3vc5WFc1dGQ17O/CqoFtoicO+PW6/WKzjJ
DJVgrMpQOMLtT/WoiKjrDSAFKXyw5LDxZ11V0wrUbwC1yLOojWtJJ7eFtQSc2jzR8quG731zvIlq
DtOeYNYY9qr6R/PEjQHA95Chuoghc+YxLUtI77iSjUcq2QIBvdeiLVufcQmWU5SeQcmlkWwPGJxI
10q1+eNZ+XOckugF6CkNzWBj+NFW3AiVfRwSl3Zy9ERZUd34s3uyFij1qv9/Wd79CmjFZqhINsFx
jCnOA8Iffl+rRmqBe7cTsbhEL6f+7zRkrYV9WiDKeL9ObAiWzBVxq5dc6UA5D8akp16F2PIU8zEc
vw+9BYpQwQFnTfbn6l8eUQe+pm5uXLWr10megBRnctdmV8OukIs86nG8VAcdrX09BiWR6oJxCWlq
dbPXX9u78hchoOM9go5OzVv8RyQdpvAFdFUC77pUK7M5uoiixQD1rFzBjWFJB/dom+uNgzDFMfv6
vpmT7KQoDLdHASnIAbMgSYORxrbh9jT6wi7E4KUSGRgYahC72IwZAGUfON1TDjdky5PI0HC+REmP
aD9Kv8p1xKYPbb9ax/NNOHHFGacIxQD+leFihTVVth9PaRjHHWTZSKwIOa7DbWKvBnFm7G2Ck8fq
a1JAYQn8K/aH6EsFHDH1YOLXiB7CDyGc/T1Wxkx4T9fcRQsa0/m+D3zu4v/C/pTVIyfGiUtKAszK
MjtczHCkVrINHuJPXhKTovGeO3el8xgCSlD80erJTjhs+nz6Ap9E0uzgniYU13OQNEj1j+asJoiw
kWE3ZrvAn5OWk33iRSnpb27+IupyB9mTMRySvt08ZF8P9H/JjyD+FdP71ZrHRMyJ2ShLqq4jdSXw
+36IVMeAsj0qEapOVtBzULol9Pfk6fzwjUMiyjl0Zb1qXbifhH9x59PbLr9mtebhBK55CDI4eFIm
h4gb/MsptFaOO05RjNU88ph6wvn+Q0A+CpxLLwn3Pqw5BjbdVRauoS5K/UqvkL/Il2LGtNUL68gE
WmX17Bmw1Hjc6A0gNVlCSjZsNAEjnzEQ3l6dZ901UkwE+mDrTTgeJkNDFc4q7Z0nEeIeAUcMI0L9
B5hKr3rGOa9xhZuFwFBsoIeMBoUbTXSHId2spHR9+q8QjcgUyv1iCLuQ87eOsx7zecdlFVSQs66c
Ygvt3rhDjbijh3nGojD4Io7C1xxBi+aje01GuA8ytbq8OY1yAPMbcUd4hzSBgQPeia4Q9F16Jtei
WuBc19z/f8nOcyI2/0CLSQvXaAdqz6X/AfB0SpliY1Nmi/iDmXPysz8RMvQM7Yi9bpzDBXJQEiLc
a0CcxDBFkUkDTQAY/FyRiJCQHlsoh9AZgMJ8GHpmxKMfajTTc/z0xJNGTjVESCQTW8hMmmuqhSxE
ZPNWAp8Ru+iWIYQvv2w5MgVVv4rpzRVCm8Nr/cph9reAtLnEMZK5IzsaLiHoCSDNdeY7eKNNklFa
aHz5FEQIuOyOEkW/IMB3xhaEgTeQKbX1aBiEcrDsOwg/SfzmrzHJ0icaoSYynnwC+/ZGkVTvFif5
Gi4NJ+fTcWBI5R7owDPQzU7hT0Eot0VmPFT1hSsGlXrKsS/aKam7HkRcwhSelNc5w9Rj18hzDKcj
qI03I9mieBy6y7Wbo0yp7Oug5iSpPJX9kLcuATPWQY9fEPixv2SCRRfct/WrEmtF/GJovf9mePX5
eUeS983skIAk/xKW7iOnrOOxnYVt+I+0uoSLozuFqCufkfk32Mnm17nRFKmz6cD2mRcic1MJiL7/
3kLJS45YZacCr2OQGIfAvPJ42Y9ntZ04nsj8+G1yIS3g26xsPaKxDktTGMH7WdLcXdHLNk7MMvTu
tmlA+xB5rPssf25sxfAZYYOfVSs8IvjJ9NtSeolYyZlyjIkiAapfslEqOVnkud+hR0DgL/G5dSsF
I0NbXRkaELUFjdWJg9C5Mdwz0mB4hJvNISFARz2Qv6SSoRpzDzZLiI/HiN0xABfvje6nOv3bIYpj
7lw7hXODsSWBhyBImRpH1PXVTV6KBZoxAYbJtf5GdiuOgG/ToYSxiJ/AfvBcj5cbjm0z/NUpZtP0
iCCWmcSc2dXNLO1TMZY382C2X3f52iYax5GdjWYSRI4WhnQBakvlPCXHC3k+71R7b9NiO84pDk+b
g5dVtAUtFzf9z4RIij08UFpwYGWDlkbQRqxaZTF+YbiAyTMaOxOPZ7Ea2zaTqP6MohOclkBm6+8E
zdPqyAtLPZlBwo1BZICioXYcjdDP5IzFQTpm7cqMVhj014Nk9MREFN03juzJQNGzIZZhSukTZ6tr
5VZl86nHg0Roziwjmeoq2wDkkM4Zcu7kX18VA724cmWAelXnJZZzMFbfpqGHc3zcWk6Acl2K/VVS
zplBSqlAh+MdCtpjZRIW/8zety4m9Qn7Hx1bIJlkz5hcORy4ZU8espKYgMlmRoyHTB8hOf2VKl3X
FWYYwUCL53q6K4rF3rBSXMTwAhnPs7bNry7QNKgMrOts7223l9jVwn0zj/3xUKgrDF+tRVKsAEkG
XSjThOeXGX0Gq98EQxl5KCRsmDFcqlVcUclq8BR9+nJnQw+Ui1rYd4FFRBvopgY+JktGzYdEJBRU
uj50BorK9mqHCtkon13t4/kdrfVPxx2z58dpXloLDk174PIBoUZvJ3JnJzLgFYJvS5GBD3xrVd4E
OYpo7cRlXV2mnkVZ77eRYoFJt8okpHracMqo4gPWrEp+BrlvlyAPuN18lS13cEVdGft6J2TJnk+g
I/+nsSO+6Zd/2fenLhF2/DGuFbA9uV4e8MyKBwbEcVt0KDKVSkzXS4xupUocOnp/hreyCcz0HMVA
BT73j7WaNPszQgapoGfeqXcVSjY4lp5jDAAoui3aAgs4QIp6Xa1hgAXPYR7YxFZaMAwbZB5SobvB
XRaYRV8+U2eeb8EmMhIZcMIHqDjQIAWQ8giHSh0WBqhekAdjU6WeqavYaXA5I98FC9siscJRKwit
mqQX/TvTVocBybon9mLn/6rQ3VYhyuzlDgxoAXCN4ilmbNLHajlIvf9xFq5PCW2B9ri1HdgPsTtO
qeZoBulsIv/o2eNQ/Uu94x8eLdGJz/3KxohiUaah0zXQ0bEeJnetWMziq/1yAOLv2RCAmxhrTMIU
cNzjxc8oHcpkYpX7ljbGjg5qOzvWBtlmCMUJDFFLHRrVLHIaKR48zyCtfDzrvXoEoRrXwNkhZB0N
red022F/1jM9KCucmR2O4k98icz2vQlvcEPzJEnbpZ88pbfq4RmJCy83m5wAdhTLTt1S11gRkOLq
WVP1zTzdBEPwzSF840OfIVS+BY1yZWCglzU+9Wuqm0bRhvCnJ0LJW1jm2RQupT0lRmatgJnDHxZo
l/lhzldMfAbVnv47OHnum/absEQBY25Vkc2apGFUCIMhFEGiBp5XgU2JSCLYCEwnU9IrTeBk/zhp
CZO1a73UV5iGi+9OFga7kBSnCxHqkccUjbNmdbc2oj3WH4co3D3OSxqXnGj+esZa7Bum2blnv/yF
iJzPNuIjltYaVwAZAnCozQGsSG/ihZPwNGV8/KasdYgo3p1SNxq6IXZucomze34rWFDSXNkA84ti
Wvho3xMD8HB1E0efgRxnsSc6A7KWRgS5hYnC/3L48FBKnvS5WfMMo2vdEqnfCe4t/76yavc7oAyM
J6pT3Hy0QiFaXx+uyR6XUnk3Cgu3iuLJ+InPtShxgv1Ml40/YZgqkN547qqLZvL/OS91yd8pRc3h
raKCmc3SA2tIggMbzROLX/0BnZPSOnuA+Ydklj30JnuQ+vvoN3RJaIPeCll9ivsebx36bHp03LSM
NZwvsN2I/R0+BzogHxPzvIxtYvMHM9Or5paKljkWZ3ywIGXaPQUIqciiOjM1u9uLbmNLB43eiSSG
jt3TCnwMSJi3IKRNJhJ9KKEONlQfBJk3yFEODK4pcB85jJeNv0bwLwkLKZYyFgXJPXPhNsmrtYwn
FAW6sFrW0hycQDLHWbjw2+Q6oJ4CUB//Kr0gW8BAvVw0tER0QY/XagTUonKL+lQBFznIdNCeqkwA
eSCIWcmc8pcK+6dpnZQGHxyivTZO69lPcNVBNZ+P2DegPzTWvWutMIqIWg2cZ+sj6XkR7qcycje4
dkZckQEqxrihrmRHPviZJcs8mdh8Tr1ULDgLWWwto5BBrmfRiPVui4BplhzXxMwadW96vmIVZzjO
NmkRn8mpK7M7eExJU7Q1l6vKuq6PAtdyeOUWN0W3xaAegiOfaJGd8vrxgq7+ofMvLybP6Xv5DFz5
tBYHbdqOjNz8HlaUunWApTNf2sMNw6gmWCu3uxdisyFdDHix/zm63EeC7zBiGGWRFazIIxwvdq41
ew+qjNX1K/Ds9hjSWu3Bg22NqL91IgBdcFZFsePVz5CbWeFAEXWMfniNJL44DucrZun7LXtvSmPK
5vMo19UFD96QD2JiXBDLUKVhTEOWyiu0ItSWTkZreV/qdHM4TSSYcmeGpSMq8+i0WytkfJRLGe3b
d9HcaDe1VEvuNAZS9eEzFAKXQPqJvhkH55VrHF9ptnLuuYNV/uFYAoyPalbQU2vmIz0UC6imfhFn
Yj/pgZKsaqbxBWQO93km8yt+6dKF0WgGgw6P6CEWHLa3ilW8H4y9YbvpelsRUzQslb4l8CMv/jut
CVI++hk6xt/cf73RchVbXT1ef2PL6WOi6ycQ5OLMDpcE3E5SEW4L0HnOZANwRUbnfZke4Ke/iz8b
7XjV9S408r8iNmYlGFfPYOOIGGOm0vFrXBl3HHy9q/1uv4aUqVd7AwZsfQv4kqE1n85yNxzhcn/u
KngMD0vsnpYeYzIpX9sccXh0XTbUKQHI6BK+FAqvRvyizSiRByQjZ809FRnWr4IXk/+floNHsskL
sRzgqepNIbeQNNUNT3wveszxPS0huuB7u1equTMLf2jlLP5i/JClaVtpxc/btINaSMMbdz44d+q/
AHi3f+Wc0HztIm54gBhsDI+BtSd9mVpC0MfwD79FD08hOgq8MA1rKRywy/YnlegZgQo7spFIlB7X
n3Whog1YBgldfx9oFfCAHNu7NmP57w5S2nLSHBSUu8eHI9D9FMpDpm9Lhse+LZyTTJY2IBEO2Rcw
52Tg1Ro8fiAMaJ+nQp/BRGCqPMThN/cLvRyqSWfkXATye2tyIdbGjpvrLhqiAdwk8Kj39gttSemj
WbjTD0v8ndpGWTEphMMGNrJdqJQkBe49LJ/MTQhh0Rh5Poz2qPf2itTcnKObkBHTDoxqpiR4we/0
Mvm3py0ZOBj1fmeSOYUHqSTEtRgOLIGx4w9TTr0EvM9n+y/6zcICu77pUBUwK5bLnleIgcGW0ym8
Bk1i76miHqKLzu1V3xkUzBpOB0j5Rd+BkQGX0nFSoAMoujM59qHVA38KKmrqE1AbXeQIfmI3O+mX
D2zfkWubahUmplJsaB/hcLBVnm9ZsvQfPm9r2uuzzmjFpqq3Hpo6xXBhM0xT5kZZtOUr4jByj1TH
XTM1W863nYMVOXGYd0tvChFO6TSDzqrfwIvkaXoy6xBbrpGuYLiH8vdbJfEjrAl5f9Hu4O192G8w
ATchKOk+23qiQYyoEmmzNM30I5IXtBw8U5Q6m00xuaSjsHQrvPhGXZ4jQ3QJ7CteKHP+GcZGVN9M
MEwWJxIB1eGa+tqQatSXH7yNRekwWKFSkCsOcVAfWUmZyEoOBm2jNy9anau/igDaMajQZycbh3/0
z5LGlEM2+HeHjYnbZ8KCu+R8eHRvd3YhRoIceV0R9GKUJeYaNQh4B37Yn7eYNCYWtmb+B0Z+LEqT
RevuB28Oyc4gM0VcNEH6A+YhkypRI3YH4ItTq4rkXxtNDq1E746OQUqp29ImXB2U+QV+7l75HON1
BjiazudAx0u/BejmWl3CtlR6Se+WElCn55lPDV5384exmMSiwfdhj7qIxjyjaQabHaJYqkzxGIM8
CKJ7n6YLRBtMCm/te4HhpwAncYy+6EfNTrCXqsjBRrDb4zWzHmMFzyLEm53QKCJz31S1N7kh62+V
pV7l8Hr/m3dHhsfANlfRL5b04nRFpvtzH/XoIgM9qZGh9ql5UXtAD4DRSNMsrkLYNks/GToVinJP
OBlJh+6iXmEv+x2V28xd8T6stuhDba5/ZMiIamGm/Hq5gPYXaTH3Yi1ZPMq5P9NSTTnSLlkCHFGQ
BVwxV7pw9mSgAJGNPWEytfp/r6GTybqOGNPXr10vldLVwhwALFI0IW1pNKgHE7qDeQH2nfz9temQ
lPR5hoXBUSasmD/kdz+90nW2l7sdlJKJVX32qXzeg1xflNFocImMOiii4T9f/qMeo0iEMPoOL7S8
eO/zgB5tu28OTamhrzJgKdrYJsXRP2EaeD5lXPxBVl3KReC9uEYmaaJLNzjVw6lygboprwu6Q1w6
02lzJAJfOkMKRqcfZBAgDPAg1UPqxTKkyEl55t/l4G1umeZNC8wL3VMv8oPv9AjUjyBi4098ol+l
Q7cZJScw/PemaJ6F4CveLWnGg16rlaMUCLtqCY3gKSRPrUNAvN8FKLEReMIySjlapEaFlHDScWo0
LJiZ/1kT+dVCdLezEUcEW6QZ6el8OGbS/98F0GiXQTwShRMyEs+/+LgLin2Z+yixv4jTMsFjDD3W
6xFLgqdfqSmQzbvas7QTG5k9qB6cLKPF6GZemTd+i9kgsnCy+jpC/mDrogO2kyCQg9h4R6Szx4QE
CChDMyvEN84fqJvuC9HTUvrHibxY4nKS8/7+lrrWrQHqQLcdwT4EKUmmmjy87oAkH/JumvAlhe7k
Xf0FVMco433TWT6BcTH3fbR0gPcF+JFG4Em2Dqav8/Dkh9z9XQ/oGdyQ3giKC6USZc9vmD/yKa5p
b5MTr14O/mfH+7P8jrWjfV3yTbAKSnKdDgA8ZMvBSIK+vDYcCMIyig2HKhcHkahPv3AoNwLGMlZh
Z/jQ/PvKo/9VDK6KLrCddWJ5WL599yNc5UPQtZSkGfyXdY0jqh3Y7rwyx/I7FrGzDT8g80su2OQV
k01hJNhiM3Ml3lMrszzn7HBmMMs4N5vyhiDVO6T2I9jhkpV/f62jlM7wJBQ8HzRU2gJR7wbCWgUE
ZPkpyPUzqIkecE8+B7UTAQ6EaRmFwiUurHAHhaa0OsElkWdCro72U5ACOnFm6RJ0zIuoXyR885tH
+qRzFewhHyDdhjfpA7ZFLs5+gHFuDGLlw3L/mBzSjtedC5J5WvFd9/oSj5mzHDqNmW4IRIDO3nTQ
KGdQ/wjAF3txcW9J500EzLjZDV4Kkid1lhGsM/Kx0I+4+rSCJpXC3VsjKMQHsbgHqo1jV5Nij/ep
FBXtnEiMcSWP5BRLCdy162g/sAl9z0IntkNPoM4iyjrl60MyTuMzm3BFLbLmR7EoCSxiFHyMCiqq
+hNbQ6rnAssApiCRgUvudB8+RzFTj4tEdYJU6VzZ62M4TWvjmc/i9rL6TPDri6/up6veq27+Lhn7
9W9b2Sg92CjiIrzVSX7N+QVlLNqVC2d3a2PMWv7qg2YqzKXwM27ykmChCnV4lYiGLWpOvts/3v3e
ZfGLDHIVmiDTg+p/tGFQDtaYKR/0yB5/l81yV/uGkJLXwfuSL7QKi6PbieeoQDMo1kvE+f0JMWdh
B7eQkYSSeAhk6KnKmCek/ZidH4aktPgWzRXXL/4JVPgo6yBwO/fh8V1Y2qvleIW2K91Os7nAzTLP
F5EjkykaJd7LNYj34Rb5KVzDFQ9sFgDzWXQUBOR/emGo2EditqeOmXL5vXUFrixHzrCvH0ysCu/9
t8O2KV52WuincyRmk/8cvZmOcwaNQNBhp1XnKa3eIcXPL+73BhA0nS6WfPDcrlinf/QnLwoIEeLK
U7sudVU8ipEHsLf5wozLmKAH2c0AQ0V7XK+oDkYOdkT1nqz6oZRqYB/1dbcenx1jUR1lTo+08Bk7
Lh/I1X4Ik2EaKblVlzR71L9HY48AO8d4rTZKNGlsvZvyrpfqkRAOFO4v1qFu4iTCHfVAUk0j39Iq
RHSK0wtQqKQhKx+456F5OZfQ3Fbfcp1ggzaAxQ5z7eN81UVqVUrTJdPRGTIJ0DVa0Fy2Ke/Lh7FJ
GiUyDZwVjdq9MuNrfGrNHeo3Bw8N2Q+OmM0jTd+mR9f8b1SE0rtYXp4rADz63UeSFEzf33s8St3K
7c2X2whgj11+faC5Ji7frRhT37MJhrrW3qLBVT2mZs27M43+FZbiaqbmXueEc7XyvVCxM3thPOEM
7EFOSXH/Raq1d8UNJkKvfrod0Cms+aLbnMt2ffKcoCx+bNbRFYV6OA82XMBA3Gy5W0sD2ZyumZoF
rLi/Vb38HxQTKpsyCtFFYEJ4YkB/Evc0NNjsRlqg+AqjBQ5bItqBWHjRfTCxsN7hFHgOm64xJfPX
PLUsqGtSQrg7+BTaTC0FpK29AfdO1lRYvf7Ye/LPlaWFrKH/JDMBqx9fJVStx8jX041rOhMNhkBk
+IuIjL+sZrotLscw+xk8iZE3m9+dIJ1axnHQs2oYrS0UjD+ONnHRMIzCRpH/yd9cJ8RPNzpfEJOb
TKattIMapC+fz/8GHSAb9a0xqbkOOIdPxWHt/A5TLllbJHG5jrjp7MA2ilxmp3s9rcUiQMqOXNWe
pLlUGHZJaVql6OqIs4cRTCL5lcE4fAJvYZUpVXKBfHDWCmHHqR95JsojFqJUmeQLo5pAgIIl+NRm
FTOKBccFh6T8pO7yYKyzNPu6/2izyPWPE58N9Gwn5606PBUpWNEpBpVZv39AH3tUSSgrbGw7frng
MHx/KTsxQuzrB4UyAwPfL9RrY4r8lwpKAR17z3nI016icftjvqpKq+z/NhmbLanKNnAV7F5qMGW0
bVGHFsO0AjcdPcu0MdX7MfMdh7b03FrqF/069RgE2k55tyMK2icRSFOvpMV2fodIn6eNx2IDYQmA
GKbbP8JaH9G3hZUME4pyfCiKAws7j4xmcg45NNpJRDfDrRU+VDOo2cwlYu2gktERVdwPz+0M9Sn8
kCrbHqDTFlBiohrRuaieVJxbYv+pMa3uJs0wOu8WVE09hrM3oWsXtAfkAOPNZJIgUEhjsSDAqvRK
2sQvfhcrpGeTnhlnGfeGOlMD/As4qXozM5ngIF27Bslwn9xZaSqcZSqM6dGy2ieDRwm+q7QpDpNB
dtcVSYTbCvFJcwZr9B85wHlWjFuglWDdzSoSrMLeIle+N6M66+MtkFv5l+CzhdZIVZtQePE7rU2Z
oIPPgYi7PkdQQT9f9TWg9h1FYT3hjW58hNL17VLyd+hcQ70RwAfnHY+0NsUgaUTM2xVUEurzOLI+
ixt6wj4/G9SwKKIMWYMiqLpBgF8C6lor2zKLXk0fyTmQncBkS18jT00UfTDNpArvNfnZ+yW2uDBy
GAckvtKnjoavD+eo+bRQTwoQtOLUWHyLR07avxRkq4EzWORxdHJxP1CXuDwY7xXq9i5Or4obXOnr
i+e8cmO5qI8FNZXmsWePjBcjRAIAjjUAs68QcweeTlE4/ZXksomAgKqY1JUcqe////uqjBtVcM69
uNwunqffes/FQgoFOUUVw9GKeOdRjD9PpHAGbXy95Lkzzv0vKb06ZEdj+7v1lkjOt5nlgGiR7eLi
rokzfuRI3iUqm+AKhrrJ7AiH8u9xaEIg/+UoJukeWU9xA7fnckZxsk4caFKUGrX0wTkh8iwGWdMT
Ku5wwcYpEtyGTl4+Tfijc5GFPjE4tssMWkYQxHMcHlQXWNQDdEWoSyTh5F2pY/N6EjDxVA0AxE3j
xvx3IX8lEUGCkrjDqlHv+CERjvUYio19LMGjGZF8j8xi46HzMhhveb+mvu09evo5NFjr/wAWDhmh
txsZ+sknQOspb6u6fLjWX6ZS/9GJzOymyI6cYyIux3S6DzGHxIxuu00ONsR3uVAQVKpN9xdb9KvR
SkRqhdha5jpLORzzb6YtTqX/sIdGPHRUqv22q5t50W3cQ62sjrMQGmr8Ssz1UnMI9shDh80YM4Nj
nyECbJ/YzpVDYHvfKCeWs2oURD3I+tmqheVRAaHDomHWwWzGxEW5AKVEUUezvqHD5f+ON94OISXl
tJbBU5fjPUDbaj+/fm4q1ykJKvKfdklLux96djy4IGTLAzUUJb5mhdLjtlIjUqSGj78Ckvp+gVto
agqyXv79bXTUq5XxFUG+UrXr8bsDhP/TgqEtpmV4wLV+qwbcokZrknpDJvREGKvUSnBjMCg6Ys8E
sB1eS7U2fWRBKC2c2T9QViXdnT1FVzVMSqANQ0W9nZhtGSyPt4KhUDALhlBZAv+KbPaXf18y5LdI
NQ3i2Q4rLQWb3DSuTXowrgX/vqDwTCFT78E7W1KGpHYK0lkidaMrsf+0b9tF2NwhYyaBuImiZHTo
FO4M1TfVnr5AUOQUhtyO8q1g9FdAyy+wLsNJRnTiqjYGp7U7aCqpMzj6KgNQfoK8ddaKq6DJtZn+
w1quap7Ouvek92nZMt7v30TJTi9JLwGX0YkiIxt4g9baY3CN6gxDIQXKuzitWkURD2gxJ3WpfOp9
YNzUrQBNomtsCtv6Xp4MwNKthiEF4iIXaYl3RdG96zahXI1DPpjQsl94sdiey6T1OuhVV/kkPyAt
RH37DOw8yaWNP4TaJGNYH+yV4gY6YD8Am03NqNvHeHvYFxFPkL0jb0ZzCOtZd+RaFVPtsY2S3lzn
j3DMV3p41g2O1f3a0quLO7nGkWdirj0mzsb629nKvlSOLQtHxIUSOWMCxQSh/z8KZXSah7ScISGS
oIW3qjgNNhufg4Shy61dFKVF+g1PW1vhB1vx1/vsp/qOuJoEOBmfaNtAMjbTj2oajcAaWjpu9Vuk
zvOLojqVIG6ekIqf8Ev9t7vdh+eqejdV9i45pf0dXdoKe9v96+cuwDDpFf7mOdHljuUzTEk4020m
JbampR+VEmJDdOPUEtJezwSf8uBlWTSlVelV112HYf8Ae3y9obdNRge/QVnc0vvUA1DeNnIwhxzl
q/44iHOqX8aefy/vWyLWz+G5YMpJBiYhMZeRmRS3nDj8I2se2r63/0eY1aD0jwRp6uep78K2WL2E
4QpoyM0fQdrg+hYR7rz3HpLZOGCJtznN0ewsxBpxbJIot9FVQbGH5MYWwBBVXIcPsS3LOMAaul9h
iGZBveszxx5j/5zuNqK7Cjoi231awePd5qs+m9skDBLQfhoa8AEqdVeySZxcrcXFJz3SprnS+nko
2CzbDWtEAmKTy4a/bY6vNMnkvbTSckNdDCfoO01YEZg/MEuqpdIHv9OwcfMA2XOROSaj6yeQjJ4B
vUBPw2AbOuNx21F+8pTpDu6um7QNvY+ZFyk9kyA9Mv1SNnXYmkNsTmRAYZW5E2+pdT1dyra+39j5
18MxB+gCi/0A0Bor+AV3MBBkMwaVGWJDZeiCEEXKAhBn16bBvHIBNRKlU2jxvEtiPd/NqFcPMtfg
Xc005gRpQwY4hA8oRRoV2KJa0uai7SekfKrkh2pWwF263ZMksG7q5GXVTIWpJ9XHVwFy2vWu+0BX
w8LSJbShyZ5l+o/itbS61bX+jDjRK6w99QwlNDe73yzZOe6AEHbBGvWM5iHmBpY6P7MpjEvnrrlr
+Fo7vnvd4Hqw1KmFxQJN/RN8EdRlPE8L8ekYcR+nFhOca2OH3hGv7I95sEKb9GxemLh7crj2K9TU
SJc6+4MDPde/ezDHIy1mRmtMDnhfCznTBPxk9p8VsicbkmO3iQg2UI+xkxbjVLtDlZV0UUvKejve
IgeyTAADTbP5YL3jDB+UoCA8TjgZYllRhFXWuIRgxoVFOTRZWB5EgBNoPzsO006U07UyrI+/L7tm
c4b1ca7PqaZerWhWXFgGkv2rJXcOPUeoX3XvamzJz3sjXWKWbkvSuAV5yx1Q4H5NQdqASjoDKRNk
wuYeJHfEHy43b4FkrErEx3883TA0hxnQX8b4hEr57hBtoyVXHXPMF0v41IucG4GA+/3LNDgw1NhI
pTQhfvyTCaGdt6tbATWd2zDD3DmpRqtyW5tG+aPNTBnqCsnAQLuF2zMfZkSWKm4P+fU26LwOFB4n
V4Gewa54y98kJ53Vlk5GZyWAg5FcUog0MeaJ9dMDeK1eVVsXKFA/P5EomxEe8jCITMDayzqw0+dp
LfCS1meEc4532X7YnUydWwlZZe0ETvgSMUBMjpj8iVdXVN6D9+Dl64t6yZJa8h+aG6wuDpu7Y01C
xzbKbtXN6VmViSLikjF8myQKkzb+4/XlfjpYMgbvI9MPrVSFkN2Huk06/dqrOM24YweYUfCYI8CL
i072QNBwo+/84cDuCxOlcp5pkwU22/6otFkaJwwq/JSKYAYB38iBv2JXb5yAR1IaDs8h0mB+ncBT
FfQ4mrFsY5NAui+gOQRLAac0FHKqUsMH2MwT4j1K9isYSEeqYb78mh0ikPvV0cLFlhM+UUjkfdKM
OTst7RHjx55N1Rv0LGCo2W4Z2Tocpovrm6FJp+IT4+eyd9M9rH+BCTAexCiEHmu3X9jM5Y2V64CV
bshOvfXDU4eEJobmepDW4GmxIg7qPiPYrt4WkYn+L22v4HQyOclgataF/iPDspSHyXbgoccxue5+
3oeVLJJGp+5UzfDiG7VPx9zjRveE3tH7lrkrj4Pn2Bac6TcH2fqi8bMqbp563mGNlmDtux7hvMv8
vHAT3FWJRSk7iQoErEL8NLAijf+BWbDPTAdNMa/aFfvdv22q3wHp6ZOKuKRkeapJsdx6UfeQntTM
Xyioqdjd+fppgoA67mvO+2Sstf4V/GGavbSG8f6zKjGuhj9t4tXtAWL2KEI3OnYxCMLlurFnZlz+
YwbC1qdErorxGnUAX19sXOq1jqFpull8703gKJyAQMYKNmMfwRZViLDR2dlgx62C4Tq46ictE1N/
LCkK+WjlqaYM7XM/eZsuef9rymZPaCjnJ0LEJvgFVI1C2jKS5PcY4nLg3IDUWgP5BKrkEBpSdgbh
q+jEJSthcglQKlMVt0cg734Jvu0U1Gv6H+4bkzpCP+RURfxGNgvHkh42vfFbXaFe1xtpF/Jo2bn0
7NnsYBWyhK+/kE1mrdMXIXPDi1qUiN0R1ZeFfeXyRny4PQKPHHxlK02QcQU4hDgRtCBfKJnHqzYY
R4C8A9oWg6CKyuyeKiznym7No1Pi7rO5EivNTL7Ixw3eF/L1+cDEHZEQ0zxAhrcwGuJ0zQwVP7kS
ETkeTkLy+pTc3YGM0+7LGk9kg/sNFoPm+iO+l1ZloUwHm+yXh9h2XKgoGNLPW6pe82BLb1xTHwlC
CA89ODCfYh97A1VHiHwc0+iXGLRzVC0XIFFNbYAvFLohOUp4ds+kwKarJKQfsGru5oOLn5db2IYJ
wQgVl+iIcgfXk4tCbTgBZ55V59gM/pEgfSDLUbsMa+++rl8wimmwBDsa/D58dv0OvTlkQFgdF3J5
IK+NTHiBOCCuWuGH1KOqqF1lpVGHv0KohN5ptdqX2fZoWLQNN3fzTUk9My0Z8QzsEco7aoHdd3Cm
fauvOZym4dntjte2iX58yH7S4ORV/WXHH0dVzKZXyFkI8b/5ICFpwK9n9mIFMhXxJtGqe7yZY3+I
NXelM/DNVj/w4BW2HvIYKX/KrtG0+wokCB/DPlDr1ho9lhoO4Mf6KFUG3eo0for3yeMjOrac/q4L
GUnNrqfwxGX0Ub3xNU9JZRnAV2L3CrSvxBLKGyZMRA4LbGPVX0OJpYk1z8SGPxQD28aZ0+XaPIXT
nYYq+jmI7f7Ysb3Wxxm1pmeaImBr3/aAgRwP7TX7SaATx6f9mHAFxES2xUPKG9aWcfAoEbTmtxQl
64ZyCcoNRDjZhezavv8swJpwP/8Oj/SPmjgN/t31BsEEfZX2Tkh4tWum2JBLMNe3OnsZA/btDddp
qom4/oYpqcKAxbiVbr9z5m5wczv6N/+3S+0V7r88ggRBLVCPlZhhJFoxvGiitiwOhKPhHvehytpQ
9obQfFN6YN4DC0v573FhFZWODrWyeYEJkABEpUJ+d+BXSWiEmr4Cz22sAdMQcLgZmuiP+53MR0J5
V33f6lbJjKEC8voZWRoE/XNSLWU0UOeaiZwXtThuXv4aWI40/nTYHAmgYdgk+IXQwcitLs4Np27O
bqlk/8wAl3zKSmWW+PHba6IHjKnDKej1sKWd9cRRaOVjsUmXZoXA+Lg91gqh+8QK3SXVPKDPuhxi
6/PlzI7LD5z2P+EXisfXgNK+IXjnNky84tMOzUYPa/pa0PmsuZoINyFnDTxTutn1BvCpGPVrLxcx
4uikNgaC6bYLaCPMn/E+vQXX74Nhe1fYLUnWLldCsnZrNlFugxGcboU0QcXWAOTbnWNql5X7xD9f
CJdHvPuUQy02Q41/bKygmKeAWYwgMTYYe7FPJMsON1anPgJXuYb7PB5UOVysLTEDHResoX5Fk0h+
BCKjcuMu3NqSoipMWNPBXaCY4WS+97iOBOzrdNJ32qgRh0OfW9rcvj85BoHOZebY5aJn34SH+Yqs
JMRo6dkQbJcy1/2ebpqZbN7XAbphBeRdnj1bHUYcXWrAFQ8IW2s3POt2D7n7F3k/EF2nnv7D4hDt
X5U6BTLnB11n6YJvpi7ZTs+K6+fXz3J8Gag+tPQdORoQwfEJepG5XFaQqaJo6aw6066Dbwmk/xci
96+xFe4CM0WUQ5VGUikok4sHBa5DD9ziuPjn5AvITcrEv0T3j67JpTHvd0LApGAiDJBBoMY4N1H8
gzxJxP9UJJUggYI0jRtT2rIv2ZobXHyiMJRfsDJhPeMxfOkjZMw6iF561maVM9/JiNT6dUOZtE9a
fdGSP5/z6rOBFWbpyocpUrYg9IDVnocVwm+EseWZB7IKYOwLUIKODPhiDbuVFTbYSsZW+mXyJMpg
/xMX7VfOxMkc4eR2tqjhg+f7srE3VHfgfXMBKQqNM6yv24Qp9I6cT98M+puP8l1ZJc3j0c0L9clz
RqK/QXjvMhKK4rFoKOkwd0HM6AO9wHv03gR42BLNJJFJfL9Sj3r+P2dab4Z1HjM7OqRG5olu11MU
UpVQcyN8AYVvvnjkhYuKtY1jgazfPT306WnSccxOYo8RwfdND/eT7xIzOpbbvpCoPk7U3NhELZE5
pKnk6a43Uiqlffw7vvAMipeJoaFOSe3HMWEpEtooPP3Q8ovx5nvBpTFAElzMq/N5mRZQHDMECHjX
o5kH93SBez0sxm4sjOhDkJ4lhBL728Jgc0HNddXolYfH5pyQaWu5vBCCFGaIQUU8P1mj7xiyXLT/
wjZEyHrUv/9RqH4ozyWwkurwhMMpJYKfAeQYx1LCrnvUvPoss7UBb1ummnb/TgHvyo5QE+b8LZly
sQoB+xGMDzWFScakY/dPHZsUvdEYIqbMT+JLDKAthxdUgGqN10cujQ8lCDD7Nmr7n6d4IYfdUdg1
VzuT9kA2VOTQ2eeZHAev5PUAYz1rclNi86mrUVHQ5nggNt/wXXDDGb2OWbFtdPWLAeLuMpPNfMKU
5wsRe1TvY4rKltcjyEhFiBddbuz7dwu6+n/WsQrR+HgJirzSUGr5RqOLyYIj1Tpt6mo7ZcbBFsu4
f+IILx2Fak9OLz1qqCzAPAGOCgwznS5X3t3yI6X8Af1EOc/HQ3ujtdywmFuPaLurKIroCrbN/xVR
ay1TdSOxF4U0mMUntZgxZl+32wR/bMZbrcqEMobNvmKqbhsOwEN80QGQQuAxhne7ypRQAoSFWQoR
Y4hEbOX1DuIGmG9PM2YFgPAkJCE3IpbTQlwMQppAhBEdefe+CbwBD9b3psa0dHLRcZqRocnsuQUi
RUehpuu172nCOOPQLQDVgG2Wqzin5z8IU42yrLTgSaUj7gROZK/TCXwDyzqcZXBC4zqO+ip80NPJ
6dU0L374jMvz3AwQOdARgCpnOmwAOLuCov3gAx+YGuCzd1LUOTzt3FykjBp2SLASemchT0jlzDBH
miCwvFBE+lbxJ382ixJG/mHTqs5AtpgkSJqmzx5i3pp/Hi4LjZ5izR1Q4Ai/GEFG7NB759PgwGJ3
RnWpXcaseJSnkcbdhqAfCDThT2lPouTb/WLyLKK326URxAEV+ccL7HDzT6B/5Hisn9qWGgLXE6vo
PBtCR0YRe+ikFkArXLU76GEnYXUmzLdfrfmndVlzEQPBbWPgpysV7mSI2wUZgFBp5HFV7UJCr6iT
hYAwoatp+pF+oHapYTJKerwc6zZLufIAG+KO1ibZNk9kp8ESExGLd6sgQMDrbklIdmKJ0KApJ7Ai
EM/tSxMUR2VmWVCHqpe1POGvFc48MzfOhjMN4Z/JiMwt7CfU1FmDpH25t+0saJmUzD43XAT5VMv7
c94ImIQnivQt+hZjQlSRW7V4xZNQ52jzQKBscCoURpbXtpAEozreIZYe+9Rs/XIi5zm3xkoU7o2d
gTYjWnzubvb9uzYYc3vYbIg9Zluz4Z2AqwUxgf2HqL/9a5qiq5Ifsgoci6u6ZtdVyXzoK5Zd1Uil
6mR/rqOXKqaD6pqFeR/czlnr5XTv8H1oan6ZKAbASAUZuF8nPgxxMtk7m9UzIb8JmmjrFVH3eC54
kdzLOw9jPNI2RbyRV9G6crJAVd1/k3ChRfGIwOHSYr7pVOOBFeVmn8NOcJH2I7A/db7H9+UhfRBA
xKahF0TnnTudmz9qzl+kYNN6eNLdInWdqt2afLeQ0Q0YoIyyVGa4Ux7PvHSOWEvMDvV4642x5ZZa
6ps8vNrKa7P0PoXA2j/cca7sWzjMKAEtk46eMx5cjT8zN4+BV6As5vqBfY6pKEvdY+vsNUwEz+nh
5lyZSzuvTG2kd1y+I3awFjWQU21xiSI8FiC+Mx8Mo5gukI7cXGAddjb1FWBP2xUXOhLx6Y7KceCL
vLidHzzGlr+674FU8v70WG0gXzXe5TixH3x4v/EAD+Xg8i7YCeHn1pELKpFAxZsdO1tdGgLicOB+
NLH9HpI+g0+LFAQ4+hAk1WC8X+Kl0pgMZodNZZ8l0bP8TcxNYmlCk4cvkI855vy+4kbX61voyov8
MjZrUtC1R4u0xVI4F5eTJoFHrZfpbYPEd75N5n5g/zCk919lObb/s4ijsp3uPXVXkJI4M541uRmy
SbuAHakyJIGVUyZlWUWGQ8pzRUrVwtyw4Xj1vEJ4Dd+FktuI1oxNlyd+ctmQ2ES2JhuI9P5hbazv
hcr/u3/jTpVgYLJsptdzNxgvj5tuCRFlht2fSyODUVFg4ifTUMYAnSZUZUlOcKecvTi0qmnbeLi/
/KJkxtOfksGJjvAjynaRvMc2wiq+nrA2mW6pNS30ouakkku87afKznqvRYC+8yJp3fugLJ03X6nF
TtUgDXNN1D/C7ErH+1myh8cde7CDZShedTVKEe76UlAktozOoJNkNwxvS2sdJnSZ7R70spYu7liW
Qu8WHiWWUIhGtqefdMHpMhTlN9zq+kELfM3KyCyGZr+NgE+0UzaR3tX6bl9Gt+PBLDEcg4RxFa/O
QPSU46BkzkJ0MnogiOMzkHD28fVrsG+rNERblfojJ3uwSr/MfQLr2mlEXG1muYGCDkrE6EuxGoYw
23zcCvFFyNZc7WjgE7f8CLJgEk5Du+bOfS/UKughgDWgUhkc56kQvIl78wOtzZBpQvPA52BtW11+
UST9Krc/qKd1mSlGQO24stHVP+e4PQ5N4GwANSDckSP8TU1uhJUlboyj8fyA5h5bbEK2Dobd27Lw
7TdC/y8yfMWBVkn/vnnMjqz3/xWyeqj5OK6V0/J6YagKaEs4GusOeaA90B64OhmGAJAziG5z8M1W
uWYH7JjTO4oREEDzs3wSK2U5Oy5qhdXgQsNHr9YSVeMU5zRBPmYuih2GewdUqAEJFckWzYCMtLFA
o3fXZ4Wvv34/6cLZ6j9KoWeU8jI66hldqOp58wqLXTK95c6uGf+WdpDHVgOzFRKz2hOR2wEqvUno
ury/Vk0rykb5C+i+/9s4Nvc0A7c1kUKTNBKPsJ1NYDzA2uyJ+9td2gF3Vc/DNxzPt5trd3bwfj7Y
ZZ4DanNDhvEYIrjzN0WXmLVyzAUGnlBef+k7ZkiC35DnDr5H/FFFHfAJHYcrdU97UUazUiHNWt2X
n2hXHVoBLASRLWcBex8A3d0Nfzv14tKv37gMvb3vKb/IVAXoqg/h5TT7cAul7ohOHtVd3C1GFCbg
kNrNIM8cXcsuVmmwH8u8YFe0y58rzWB6P4n9glZcVYBnveNkPlEFd2uOkNfcfgOy5omsi7zwLMVP
yi3o+Y6pO1Uii48YOgKbOp7mVhjtq7Cw5+mwq0WBnyySrlybDMVzKlnyMZb9ukhUQPinJ1/DQzHo
1FmEKnjxTN6iCEXpJm+byaM65NFfu14KlZ5VTNYAm5w9wFjm7kJytVVNCKvqwb7zwywBSJNWJGVN
YfLBzMFpF4yTc945c8s1cDrBN8WUYCss+a6yAAzPTHZtqaE882557HXY21NXO1T2A+9G9l/wLG/t
ucKUvB46AdnPqutYw031PnNpmoKKGMNcV3XIcBFexP6VQ+djudJqUwx4tSjgAlvwGTJXI1mnTnxB
dK9Nmi0boZ09Qe9ccj8qS38lP5NA1wRU2yo4hFssZX0I6UccKuRJjXMTF3wZo+1B7MsnTiA3fi4G
LDw01tOIbbK6jnAdJphv/EeRTf0xBXlQh6tXdB8D+Jixn4Kb4loFFQG3peORMjbjGuU6TWu7Qhvn
uGABpasBfgoSbzpquvKYIsxPzIXOsz2fR4CO4N+31LYmDrNFG7Ai+RkMcXaR+Ot417q79FvkMV/J
K1LuSGKDQb+yN2xgetod37cEikGtYgSFVrvRiw9CtO8CJVlzxARvEIjFRwQAxYzwEyTdRIwDh0Vg
uacasPmDyUZXU7IcBUokJJ6A2/pLNc/N5ZT84UNtjZrj+TkN/YzQJ3QE/Uza2D5OJH+F8orbMuRT
Mnqz5DCWAKEF/naveiGo0QJyQCM0/nRsArzHLWP3/we3Ldliu55jIiB+tclKKVOTeV6tBJT2Grfx
Gse5qRkN/pZaA03t+5H/n720mp+TPey9jZElr5jCa9u93HlCf3CmYwxD7tL9SI6yQc2gzY7WkEul
PwgEchHSkb5HWUqOti/EXcIx6pJ+I6uI0kVMVTOsVHhmvrK1tcIecsUwktIh0sxYPKZyJUa4si6M
cGV11dU0/uRbwPSt3b5edXf4ymlCCSKL0pSQYOZLeYtT0DaWdMgQn3gHW4ojDsC2YcrpIanos4Vt
Q7WIlHGfShySkjigzXxDpIdAADjlkCdlTsDJZPwJ5Xv/96CGFFCPO2n5ubEJL1mj6m8m4uLQW8G2
dto7uP5VITTZkGPm9qRYyK1lo/aMxSMaJt/GN3dAiWzY92GXo+wjw9GSSOJKa1V/i88DR6MZ9YY7
BG6aWZplsRcLb7/X4ZbDK0IOjNJs00TTE/nUvvYt/15Y0gCgAOLnRmUT2vF7mLvYGn61GsXpZJNc
qUU/1L0gloUfopy/sUU38/1WyaG0A9UhyocSlnxsHu1WOfolY+k2ZvPCP6a1Wtd4UkZa+x2Y7pAT
51gNsrgsFrJUV7tnUzrETfGNib0MKwwVDf2XNoJLhsVbqPl+KH8x4siReI0SgoSs7HOrl8nHKR34
KP8C6hxUdfytOxslDR5Om0SwnEz1jH6DxjmnXDhKTf7Qn1ygWRU8Fp/Qz5BVUWfJOqnPI+ZGJYE9
i+HJszLBlB04f5Efyr4YamSrWhBl/VOD28ZFzANBPqp9FxYTATcwj1O8/Cw8WdFcp17/y+NylLIM
7RuQ07zh263bWD7V088SdVk6tSD16KbDeMzksA2Znd4UNh985F/i4EmkceT4XQpsISIQ9DYmG+AD
8ZXowvGIq7wF4MMgKZGXkkKmFZRuzblXiXThx48wRXPNpF6gFawRLZDZxEh8UV08/Tg/34q30s5n
so3BTaDrcna6Fa4AW/maim1YmPGuyYjfyR8s0b/gbCGIEEzQ1K09sG5yj1VmOc9fqcdbtfMMBVHp
Jj+oyw2dWtIkKk9hrC0/wdGYJkG6DleJp1eUNKm6iE0SNJET4ZdJfj+728k9ry1EdzW7g8FlYkLA
uCE5PYeeYlFlnrjJnFPCLnIUYmMNuDpr7b7AdGl2ciwqnhfst5gPTZacyRNeYHa/Me97KLKEO6Pq
OtMJtYy7VG+0GSX9a0S2Y77wgqZdCJAiH3r4FW9urN4jrE9df/LE2dXkuAlWV2kgSwyD0t+yRSB1
FU+saZdtb6Ad3sXj+kkz/G2SS/4D+pXyd+Ty9CizJJvmqQIp0uTqYYG8AujjQhFX++haHNNDWr/8
7pamYD7/c1u/8qRK9lWtrxd3gA18ga6O7HDg/EQl5t3rzTHRE5nwVNNJmapdPOBkA+Rt7j2O8ltF
0Z4lQrq6Sl3rYRiuF6lybbuAIEi2qIn9klwsY6ZhnlCV9ASgSsHo5cIP6cX+2oMHnlBSN0NayzUZ
ExwnXyQVinwNTNB0J+itLmZk7cJxEqF8DS6eiIWXNlGdc7xwStT2UhUSnIEZHm8baLK80YNP/1im
Tgu7hKYwW/NMMV4qhH+PKEH/EOXyZlas+tYHwdnT9Hf55ct43CdD4JUuKqNRvHWZ45qLoPdBsMEW
q8+h+JmZxpoS4RTVrzxBuvkrn3EWgxtGQa4zPpgs9MKsCnExs59xcMTs8HF3e4TkvoVkdQEKbu0R
STxn8ClBnk53Aaei/w9C/Eyw1ARZsW1Vsc0KlV922ejP4chmKImve7zB/RaYCJAYKI6dFBiQXiR/
LuEelMZ2DKm/rovRxzQnwPMoq4NuEY+Kodes0zCm/4gOoRdbOMnWWSrrdxVa/e/d/EJRrboJSLQf
1DFqevSjq9O2CszARYvAY0FCLZ4dANxppAtxXMdjZF9Czq8BPYoX7isiEUhgcfF207TOAXliWBVm
Db5Sr3mpArS1mKZDgD9AfK1Zu7gTwlfgPDMs2yjLTLDaSfmOFnbnsIcrideNVB77iQgDd91UyS40
+vRK1RNcr+Qh21cfFJhx1XBOdLKbqS+ECp/ykIgxDBKqXlD43AWGnMksGIi8BMSs6cMYj4GCK6ZR
kPUBqNodhOzBqdrCmV0FNkBWoQWHg/OMbBCsAGiutqFyDarX3erLR6tcc/YB/XXTnmfj301gFzkn
yPoXwucb09vCn6VopEDsFzZdqX32jLsnycOAOa+HgL70qo+Kgqaz2inNgdE8qNIDiOTiZz0TPBfh
afALqEHDIiCS8VRliCWINYk9jyUVvcphAub483dzWqE/131a6ogl0DjRLLwGW9USbwKt2ARZRWK7
giSWai8x2qg5bqe6bhYJ8JA2/6kGWzQsQx3MerKWI33yd2QkUVQ1CBlFktDRk92pECRc4mbBc9Jp
aPCAprOjo1ZL21QsKoIOsSnVrWDq6ukCKBOV9XAC3+Q6Sb3OvtCjjzBNqOp7kkXCFOa0LsFKnfzw
9lzT5SgknW8tWvD9D6oefncr8Bs60jNRkfnaffwAGzNX3RUS6CW4GCsdN0JQ8iq/hGVzAVij+nNW
sgzzw4LqRxCLtEiL0xOgOEJhgB0QtYGdSRFpsVfORbva6T4q9w77+wDLC67Ok5s0phJn7U1h4Z6e
HwlVMuJxp/BnED0H26D+TguSD0I1uukN1O8DawLKCbyDHyrmxbskMXoSwf7UtSqFBp3owHkfxFot
hu1BJ3BHLDKrVFq1poR0NhriKXBxzhnVZdix5AARZdyV1rGUiGRrZudFlA/r8nZinPFj64XUdnHm
jIQqq82NaXOndT3tuSzKic0TOdzQmrMIAvcGy6TTdSG8iMHoX46tJLSgagvpP0ORSj4bT82QjhSA
ElP5sPn5f5leZ/w52alqd/sBwUWBr6QIloSYd4o1p05srsDBfqqzaARFqbrQllWHu7TOq2uAKqXO
s6YaXz2rfo/q2SMxfx//qDW1I8TIDyUrfQTWR59Y+gN8cDWTy8Q6JbMJontWzWQjnKRuQ3dRudeV
Q4jsH6R94pWEbRVjwKt59Z3fFPmiVcDm06EjC75solrYm61T8B2SISuxyZt7v5ZM3hBmDxhqwSCt
QclrUSsaWsKQ5LxcYw+CIXoX4pPjupBE6Yv5BxHsz9e1MK28hbyKcFclbdfc5Jfwoi5IGrFIfnoX
IecdqhT+9lC87RCkdvPQAoW2AIx5imRdLWoWOg4LbhnI69Kp+w2ulItSxxcNzin+qHzc7fpiAfAR
PMNLEtpA+T1ag6WLb/dc1EYz2mdRUalIWSM9qJIQJNNErO8wY9+e6VOURDe6sa8uXMZKPl4ypGZF
MkAckUr0ocsS5SuwI+MX7RUusJS0iUV4Us2gvakjG0t0PuZBUXwsy3wdHpMUP1Ur7d2ucfSWxvMc
Zpj5arWBYaYjTyntnELEBGvWWmH41tRNp9LWzVtIvop0EPUj8aPykvnHpkLmCij5lgWBYkww5Fez
K29CbAT05wWhkImeKmokJ1ypAYB0ocEQvMEAiYiAyAMKRRtIXh8yhumhG8wKuQw9OlXreCwXYY6c
g941QqPObOIyA6L5XCKcA5lc/RfP6ubJAZzA6yn1dKJhhpeXnt2R490uVwQDqNxgliens8D8Dqi9
F8EG+J6g8E3+2hYutDXzptA4F+++OOpdLWN32k9gWWJdjGl6hsVN2/aAm8eDGrpv0US1d13GcyHu
VqBJvt6/v1Md9TKDvX07Wojrm5eOYkN/01e0WqYhJSakO6NEbfXKpxywHYTP+xyhzwwbxST43rYP
7DAoxoBaQcQXQL6m62in53t2fJPlvv9t1zkMSY80/VCRfNfNq+OGRmKZKKMXJ/aY8h5Ox3tIV8w8
KJvbO1AlCRR/HZPch8Zdx002BS1Dxf3kxXOXciaLfan1bOS30pkjC+S0TgtMU92H1LkvYiDMjnU7
1zu15c0GyhAUbgUw/Pw6nid7HKEvLYC2PThJi7Z1Alkpe8PCddSqcUvI4JvYzm2Y4C+BSoAjyoHQ
Xp3Nlq6vxZnL3pJISfC6RdUd9SKeH3BI1QeeO2a0RgkMlDPWEfZ0zjt31odtWlP4nEAHjE7Ugxpk
xPUwvBF99WvhpqhSHLY7FdEXmZSRwPdh/g0DC93TOSSRhg8oCS820MPRPJOhztqTjim1mNNzhSjc
9EiYfrtTMwNrsz/XbG4uN2aFy9taFXSeXgh/J2X5bINqPNwbqsbs9oIG+MSbvPS+hfz/CS3T6ozu
aPgCpchCJJZnFDWr/xbODs5VN0LNPdpH+FlOQj/TBTCsErkp/E/GvtyDeAeT51XKBG4RMpeO1AT/
5t1YQ+e14Vsk4GgB/GRJJAjGNk2Gx/FESRQQ19wTbcFbeL+KUYA9xuJInApKki25jo8gX8/dvrh/
Ck1pkFTfNeVcsjzAn7hpa6fwb2OSsN4ap1yMmGxHzMvwYh9G9d2P7ARyjHF3iVbo5Apg3/zxHWv3
QC5wwQnu+GEem1CsheA12J2awzNfWq6dO1T37F0jlot9BeuO+B21MdIolz9x2QqaMJ+yOOXtTCvb
F1GVin3vtFYKXzOlUixCQI7IrLXjFDSI7/NAtWBLKq6kDbqrbu+17BTn8cXkVO4zwUkquQYCxi7Z
TW4QUL20LUxiitpVi3WNqvxNHeoNAR6vtc2KYW6lHK5AKWYW93V31vee9zJaWuKsKrDKZOpGEkds
GfiX6hhgMJxDSOclehtda7naQJOG/ne5S06uQzGJs07526zr1m0l3GQwHhI3ZmTGd5T5/ZTCsSps
A1ynd/kk/v9qyoA58+lT7jtSzHcGyuLwh1GTtxq1hWSvRibRzIHULagCUlhHdzk+wk+NY0BcYVbw
ExaYebicxFHBzB7JfnkBrOtKbYYlSC+zFQZoUaSniDV5xP7u1DuiFbbuIAAQ36tUVRAWPqVlhzRy
qWPns9MnOEfQN3fBF04jYPL222F6MO9HSX/3GBkGFhu/XjaqutWpq6QJu1brinUnoqIyICcy8DBP
Y/lxB8arPb6XteIqQ5pB42qL+EIBYSUlr/rPXEtl5bzCt7q/yoH9gewvuKJjBPYHipoUHlrmtXDp
sOOrsYFEBRx8f05JNey7m/v3XLUjv6qnPtSi/LE8touduW5dKfN/1kZBeS0d1B0+MxlmwHmxgslf
F3BJX430sbUIaxj0VNQu6AtmWQnhBQdp83U8jsGui/H1SV+Fi4WCVZ4czu0pLRaB12MZpofxPxxb
TO8ep3ZdDshjkA7ICDhCP3x4R9h/ZZ5NXcd2TxQVf/DMo6Ju0Dh8QWcyUgyu/n+MIleK+fYQ6Stx
aPwulJXMS7yNZczQobadkD/iUvI9Yj0R21kZ2MZuBopoRUOd+XVMsuzajxsBHejd3ceNEkCLziuy
12F195Iv/RaWYnd7ooB0Yrb5xsp/rKoAZdEnT+UWdz2ps4A0fb8xuXRxVdtRtthxip6lkIVeCEno
zLhlA6TMscyTfQqTeQLAslGC9yFwjyyWqBBE1FIKcL3Anj2DNNUWs/1wyed2P5kC5N3cwhArQLl7
vguJLK1sa1QZXOz4nstbTTaPieaa9IknN/vAGpw/rHn7YMk2z7Rsju1d2qJZq6tw5zYyfsTsIX5d
ySzsDjJ7P13aVTGeluRPcEdUwHRX2LvbVTCzcMDs9MeQ+CnUrKJ6m2YFWq+qIBMnLWsc7rMl/LLr
oKg04k2PBCNKv4Eklobpf/m5XV9AAvng6KF6bq0njs55ejM1x7R7RIMy+5/G0ySoP+tWw7iH49Sl
Dd3IbAJ2udB1LvT9OlhGknvWsiZPlqBmXuDFLqQwx97BtShwK8Hros7LRGrpi3NQh2JC/91Fq2Eo
L3Yv1GbJZ/YGmR2IFnb6hrERJq8QVtVhCIPlBm1gsXXnRTm0vI2zk72rQJ+NrgCcNL8MwFgwHJAU
wfHLLYdXypnzlUyojmUAIDl8r4Fr84Cj29BQc7RpNHOw9NpJ3PRNHaxPMeJ2M2JqaLBDlcZRPhfC
SWY/hmCnqWnTvC0lIa1JGGryfANdEGFiweIYmC4zFGDpj4EQB+u+asCzKvWKrVj4aOzpG244TI2I
AACylFgQZcr7m//uOCSAle7sPh+d6vwAr/6Xo1AXmRn7iWhSoazQGDNY3nLewlAg3uRjqjtiWI0f
0On+qkF/+2abAP6OHnLDkxaSf8k91NPjhdyyeMGyuEyRFeIm9McyDHhNJ6Eccsjnb38Cpx5p1vK9
PIBQMz2JAgfACMqkf/3rePZaeFjVZjwbdAUDudstrf8R4IIm7wFdPTTAICRsAtTEp25ESe5Dg9Da
t77NI76N6NaGqxRGEhpZqicS2BS3+pQFrXsdRG3MYlSHsDNEObVgAbLkwJBJFmDYTptQfjXmwMet
5MKe2mLrMwSZhyEKSNxg8SLdV/PMd6rnfwSmZ1C68WGwTJkRAA9m0tmcIl3OaBczEBmgUHKn2GQn
JeVVRI+aTtznjRF2gJL94X9niYhZUzcgp23yhA3gtgq1yy2Lrbe5DlF5VhIMh8yyBi/yG8j7WXYR
WiO30FQa2kTUQbz/IhQTPV14Qcq3dW4OSHTClgWvRy/8nFaMf5m0daX62diLDMZ6UbyjssvTKhfO
/AQFhgE6y3Gh7FnHDiPjgPvvXciI4NC4GiqgMhHKOgo1BmYDmLkr5FAK5HAmGcggBxKiT/s/EPOx
cYUJ4v/OyklVakWxFcPnDez5vWyfVEFjSFd9V95U4mQuADn2+aPD3Uk0qmyVkjeK/1LRjlpNaTJJ
xmJW1MkrGnPgR0Tr/3u9b10uhAOzFeX0Bjp31CR5eqH7ixg/6HUzuNedHfD4xQLMan02YWYjWv+G
wh1U/GNXPpTgnfhdRE9e3tlemEF6NvujJ0URTLHhnEy1nIU3OkI3kGNPiMr8lY9gxhPn9U+rQGDN
/t0xo8niXb+EGRjc4xSdnbWdIelsJbKJ59ppy/XLGrPfglIrn9BYq/HnTm+43zO07CfokoTiqG0T
fwcykYRHtuCJRh9AL0RIEhavfJ7fBtgV2ShJMV0yzMzNuNMyOJR5qAfl28NlV5rnw/ohhTWDZWgZ
uavbKQBlL0O8SrV/9XYajPRQifIyQoNtBRHPn5F20xfZvmYDsz/LA8pSN9BnTTsKLpzSuFkINetz
n3oEtjtFlPv4Hn8qGrd4GoG8NjrMhDdAu1BRmF1oPr3tSKcCJyeUCIRGpg1EfpIqW5+yMZ0peQLl
oGA6tKBzmsLBDbxVI3vyu1F5JFWgZnNYw7eGfpKiIb0FPWQUoyHEl1Qwq2l6SyUbGPPTTtatF66R
C946GOiT6NokYm4gUbY3XHd4nkWfU5pyKnFN9dW0Px55q4x7Tht/mkdnoofISdWpu4if1kZWvueR
okEmBSyy00DwqaCTRfZ87zOWyqklpc53AChXzjDkSOz8oDwKgTV9Byr6SDjlZSxcnXB068O37Ddo
N8X3pNz1+GKdwQ1Yo6xsOwfM3pQYhxBKEBVaV3DLMTeSbKhW/Ubp5WdLotL9R2KZyEKBteIUk4E4
qIFa9c/kZCwPzoRhmJpWed1wAtNiz+dr4w+nm51/AxXJhENaaWVhfGze71uMkiOsKNeiQxXtoyWY
8La4Mfmw9kbkJ81TTfzpbOwwYTSaa0qxr86Kzc9ajLPZZhb6PvyBgT09UAy7bcR2sfycVsBnYaN8
mVBFUUaXUIQdH4Ljj2CU2gl2JvHCxFNluQWCwblxvPfbUHESoalTt6u5Djfgg4Bg5yAt2fT1S4dh
U/wQKK0kFe6q75HV10xcXhvVNxnmz39uQNDQ9+Gs0RyEs9N1YT4P73UwC3DHXRP1IranKcE8x5GC
U+MMK5TxSBYkju9JVlnMQrXa6E3gpA0pgP0SFVnS68pm6eKq9ZhiRb82aTtG9oudfLRJ+9yRZSnD
SEyOW2GIvTL9JZKUGV9yZrqjlCOj6zIw2QxUhTn568sykS3PgOPWSSoJlgJ27cGOpRGS8dEtZEGu
E1fu5RsR/v6mQ63WvKyJOFTwVYCTT0fyWzVgBYt/YoCWW0PRCUwYkHFTj1xx2AbzWio3G2n7jsEQ
CK4F1NOjTA7AqzXjwmCuqkZ/PPZXbJ9jJ6aS4tX692SB/uuvDLf8IWQx39f4uc/Nz//jr3rIvyKl
4N6ZAV6VQLk7/4v7q3zGBJSLDkSrtssmG0dJrweKxBmEAXtB9s/pYCmEYE9rOGG7/nMoAgwmH783
1d3uUmmvnTtVEkwH/zuf4J5Kbb0OicS+7lYQ4zQhVLtFkzcgEvnMQ6GFgkEr9Mxq2jDJEqfJzcuV
lxMmtie1LQct4NSs+TU5CJc4w4to1vLAB0xXtP3HnyYdPKdjmBeN74cMAJ0itmvs8HhCXN9RNWVZ
wwf19x/EGgMifOQ4jC700CGZYDWDeuCIYLvRGL0mz1mbK4Mr7vwRvVpEmP2N0l0w0azDTLyNFVie
jNUHeqINRUZ2JJeBXN7RQyzTc3HibLV90okLp41tDi0bfAc/fm3H/KQwaFcvBtbvH64HhUeaSQfo
COAGn8894qTi7YXNFW6K169Mwc4Zqu51z9cSkQAftPIGMXjy1T5B3thp25igw+ym7t8LN74dKt4s
FDnhwobJZaYIrrwRa9IzGlD85eCTCNhGx4vExRfLGYsKqSuHH6ygsD5g46o2ArI4EMIIgQIt072l
sAhUKf+wzcMJpgPcFmvM3d/2rdlSw4cAt28sQXfCR/c+adhfqa3JLTbsvJSvXHH3Q5NaphM1zqhy
SO0lE1K7Gu/8V5G7hIZmdU2ApU3ILjqoIC+vZNK53v8f8Gq6XiwiXUDS3I1FxIw8p14IaBFcu78p
0O0Csc98+FIgTDqNVqsyO448UNa9vIIuyh1vaZm4iwyy2xvYt7M7xY8zxzrBoq8HIth5q2uLdFmz
yvFF/gscYvwObfkoIFrUy9CFhG+4zLFbfMh+2R8N2+ZmzG/CZ4MrhucA9iBdD3TqPb5XtRadX6Qb
JXY4KT9exQj8dJmm5Ae/JPjKHmx27vKCLRziMkhq+HFJnBWrMzF+ShqI8s0vNruSiEnhNR78pmQl
oouAgUm8W5/4U5zar0osacUbSYqKv3pItqICTgwLNhvPPu+TXvchaHUwsLFRcGUNOvTj0lkXVrLL
iuIWu7JTcV4woWOSfRRSU6sbYJTujKaKkfxLouD1eABlJqh0y5ZjBys5GCRJjQqLDKFVyFAtjBm/
YXnmM8ZPxLfVPepLkRPMHQ+p7jb6LZIGHljSatb6tONrM0y6KVcp2koOW0u3eIparzyPrroV5IM+
XzGQpnw+5kyR2s1i8KJ7/wsz/Skc70GNgMB5WdQTJz8vyuwyao4xbmI2ek5kmWfusoVmXcGYJ9Ot
PFPd8dxkESponIFymJ0JQggQnfSylWraTluwGrlVr+kdtfI5BRqZz/SiRQnivO+TRB//E/SZeDLN
Zsu+wnBm5fDGag3xYtqxTuqUYhLWxUrW6L88sDJJO0IBqnsHUX20JAdkc4kGgEoy6XOActMCKDhP
jj9MZeXI8zMoD4mB1Le5yXyT2JfaZeFsK4A6pF7AMzMaAuuLmYizV7+FnIYqSnhDeDW1Uf/DaWuB
HiqOPJJMXvSYGngamSk2QtAjlPS1FMRk/ryXGFZKjUnQZBict/F1YpXHTlrLks4DtgcnBaTDBUgg
3N+WBRDsOXKHo/hqIcmFpkP4adsGlmrg5FaEPMpIBU2kWpphlZir8GAnUP2YPeC0YiRTMcl2kF/6
ve1d+/5KM2+/uqQ9686UrKgtVTlUWbEe+BR/eqLjwng0Pgl4xHp2N+0cPe+wefN6KIpPnyRqXPpx
DxjpDYqLPeaA4WaiKOLOilUFiESlfx623GW/gelD6hhWTYMCmo3eoMCvtdE7mxnQZN5dF9WyLwWI
PhVdRUKVGDaDv0+ENBWiSxoUuASfqQYnyBvNPohAQEdCLygKlllorxANJGzU3J8hKAT5itExSvGU
xItN3FMu6HrkOx9SE+cyBIzSj6nvGiBsBHQTo25hHhesoJsS5tnnk9VCydzbdjY3rHLsq6nKFyi2
mFKFgKdqidLCvVrM9UeVEktsEzCakAoQFsmfWVKVTswing0zfsCVkPUOd0NyWQHpNYg4V1pKkJYM
NKY/b8Cutv2x7BtWgROguczcZTGSpnT87Q5MBJOzZd9/xmO83yJ5p7dJb4OoymVZSUe+aokA3pRS
fyaGoHlZUA+uSN7iofvgYhbAAIoglKDNuuARyy0CwpC1P2wNOxsS5TvLLUyJk/qMozy0EDqgPIPV
8577u27eTQvxwLm/gs5FEUMGdBXent2v+WY9jWDd7udP7Y96yctNPrUQWqfgPTE43s01uWsjM4fx
QBywzeKbz9bcyPeoCfQUNBSlcpIjcSrugfCdSe2/MYgWGyrfh6hnNvZ/8F6FHbJhmj9dUYKRMOTb
OpsDuvYbJK+Z0L0HEJVGAVCKGCZW4SiJL8hOv765Eu8q3uhhmTal1FzCsz2s+KvQoYQak3XvT0WQ
TCj39HMNfyR569ID9bUg8pCO/9d0yjy+DQ/ReftKnZbb8x/P3N+vlP+fMpBQzJYN+01SwLaGNERx
HBmIQdqr7fD0IWsMqnLCB5Tpo9QbEH6Ric5R7RPcjhaimTIDdiHaNRMaCuq7GdgBCj56LHnl0Z8o
4v7rS22bGaP1kJn5Oybjy/zY4Q0NbGuwhmiwkCcbqvoDAbQVLC+PWv0dblN9Fl/ETr0Ckkgi5TIu
mcwnUcUIehv1K1bFpw96CVQQErUAuucEivGlXxADqVJyaHIsg96SiVWFj4RFfm55xTEko/P3vkWP
PAPS5Zo6H/or8DG/QL62aiAUnBMA4N8/oAi6wgjSQKvHWMWj1hIMXEoGg8cz6RdDl1fTRSq97UVn
pUE0XyjGXbZx7aOz9Z3joMFd8k+3Du+/EfGxYVuWZYnEfU5h2ApPvBxuxKYkGVFoLmaAXvrmAmLK
BM+89/jtuw/w9eW0Apy0veSU6/uv+CB/HdgWz5OZl0IQNPDqhAjKfC4TgxErC2M7XWWVLl9WYjQP
EsoXneRlNxtdMdrPJ6cgpNYUQT2eOoDLol7omiFBE81ICHtkXA4kvCqzo+YmQpMvKH2mJKB3QvJf
g92GAuCbbT7xyijZVZaAJU4dKkxLZxDdzlxNp7iczyES/UE2CSSDQKLXf9u6qoZWk4qGU6jFLs05
Cz8dc7QHQ6KxbSOoLqnCJVai84KEM3RHjfBpd18VXof7VzlxxI07IBAV+27cZogziMaAChmWnjVu
QcseFY7jjzsMrzO9vt4apQ8vUX2lqwE2JIs8y/FYVKwJ97zox+eXhwVRhGgWC9lR+A08VPP2OROH
Hdfqjn6yGLg0hMvNg5NxuUtOlsJr3cC1GGB8H2tsGZ0A2i49d2MZTeil3tgnelFvSartMAdrlkmG
Ewsph8OXDggc43ny9MZWLtkva6yHJAdKCvMugM6kvgZIsXfLn/+q7WoTQzZOvV3MADDjsV19BJQL
nA8idcGcDRg96nAiaTpa4AImUTVNbBlEp0J/Ban1ht7h1Hz+a0O4pzFNKGuXvW/jWWYDYESkZru9
7r83U7OUZBWo3AYPJWMnK/3E8s7GrYXmJtiDWajJ91tfuVgQO5HkfqFDj0fRfv2ZI8KUjKlxCI69
+3f9Rh6VkkWiGf28J9IQbB0TFFRv8VEA517h9SGhAxTUXfV2O/HFE2AwVqmrdG2LXbsQPTEV9koL
jS1BsJkNv2RlLVK4+kunKQoe2QuK+y2uuE9ZB56mt7JGjnKnqVN7AJHIgXkuCDqnFt4Q5dI7yvY5
RcK8NYAP+PCY1RQbhIKaykmf5bSl92f9PJPNNZPrVSeB0r9SiScrr2vJzcgGDZpGCRdliUGL4xea
VavSRE8zOJWyzbdx4DAwpaxIkXGDfs2Uy0oiIdX/BT4Nrwb9e4x6AbY56/hfaqZquxXEZEaBY1In
AjHZjCXpko3KbTS6GQ4YrdWbJnRnrj/GnyhmrAFSzCM1IwGIf2/Dn9ruIXwrT0shFijXMBAvKvYo
ZQATBSsJPTeXEsOOf5ToXdeFFYaRMp/5EwswW3MQy+JgaG0TsEJ136cEDkt5aJsIBM7KN2/apJfd
mAUYG7tBmIkDmdQPXmrShI3LzIE6KJ8vhB/bTTAbU2d/Z/8GSKKt2qP/EycQ5U0A1bz7txAbfaK4
609TpKJPOzBj59wKbkqBxYaq1MLU2pcvXjgx1zkM6hh+s/EkyGwpGhDKDxGbmmJKkYjexpexnoQb
cre5271RO9lay5HpzdC/Q4bBEcPlm3shzAHC7JQYdfMKe5621lwyF9GbkULV2i8kzGkHChg+es6c
laCYPSux7sqV4zWOLwnhvyfhcJPfgXdoArka3KdJFcutKyt5kUn40nBUKF0TZi5PcoJonUsOd5xC
uMVxl+HgcqYMDvl5J8byLabpI2+rKiQknTHtxbyr5bSn9uoKckeF6zD1RJP2IReJh4RWJNMxkWDO
pXO7DZRQAZzT5e+Fp+4kZ/VQ/sAcjCi1KA0nzA+spuqFAgjBSqdCLZvz+RSCay+848h3/AETPiwM
Lx4w7YAoTraxHazH/42VTIEG7IBuqsjB4Daxd6lfNAphU17LDgxlJfHkwivqVlinHROmIGmgqSog
d3OnN7e00oYUnEKxIONmWtY1EBRkJe/bhINRitlm1ED39BVUrvbwvJo2Z32jQlXfM42SiO51Itq1
nuWo3qfseWGwQf5g9TpVbjKBTE7MqySVjsq1Gi55IFsXzmcY1lUNeBNQywsxUOlRMmp25H21PtSS
reNqcLHsoy2FVekqVurV27mj80q8VQNrOeP29OiGIC9JapuJOx9cBnp9QLadvALAUdOS3a5xcZIq
QpyXVT3kXOXlbMoDUi73NJ9U6AFG+oOUcQDwpcb+VVDbOvGDlfAbrT88JLI+4zMFFmgcw34Y3Jkt
d0/lFJxij3mvpc6zMSUa9VwTZBTE+9enStA2ICCQ9tljeiWpkM4LF4XUZV12xM2Bi4BTLZemFzfT
HZ53NOjk1y+VNirIpousdtrvkYQOiFfVsbTLFeRlq5N8XC4mTj85dVvmYnd1IsI/E2iyCVTF61+U
oETjNhrZYr7SJL4TgRWANxZplwK2KP3MmeYdDPyjV2cWuPxgCUomYwojeOb8ueLngquk9MvavZ4x
vJ3PBK45A6fv9EZD7fJWcb7OuWvoyHuJ2gmOvB9s81dlHXWB1prisycZFZJJbTHXm8mbd4090r/l
YqGvrFPA2e+lyBE5rMTUmHGWM2WUi4lZ6Yybx6wzQczrCyydrmvnr+my9ODHkyazLmxryf9beDk1
Y44i+MOKAzJmkMu1IKIuuaY4vySSx22AimLcg1ihIeMIgstp7ckjNU1SdTpj4FTbXLDUm+AKwglP
5ibKRiv2wtADMI9qOuhwNDhTU9Ov6baL2l+4f+DGL/MFlipD6nFBJzrfPJYyPjWKSZLCgTo9rrW8
bWY1xfDPKeAHWAabJkTbvRhI/e0ZW7WDo5iUd9v/n8AGlu1e81BgLQAe1uBK//J1T6r47oHBNegF
vdr2VaGB4UxlV0webOy0X9SrdKr8ua49CAU4NxEon6mlFcpd4v4gMALDJbbftuCxAgLZsqxVEoa/
Pz61pwAbLjDWN3rpPenAlcTYkfPNZ/qEbr4GsobSgWLSqbVtU8HDtY0EbA0lAo2xcQZJ8Eb9AaVd
L78pHZpCCZBncUdIMTHLqdG4EYSvpYLAzWbKCBjEbNUPVOdvZjCZnnJCwlnitRMLjzD+bx88haoG
KovD0V9gqkwoSG5kDI2d21kvRH8IH3zG2yH39Oq4RrAZmLt4jDr9/MKtWNN877Tl3RBPNUrBqmws
ENeuQe6YlaxIpDELrsvJsi1BSGTrqykIdImanJlFBF3Fla34XE0gAU2psaYdiux4aJJctEvMqc5/
fEF6nsTgQQ+IwWc+id+l/LTT7w5sep78NNKghllicm6EmUU06fzRxz9+zIz+ewzRjsXO66+dkBCb
j/ZQYFY0j6TriaZfXRODZmHqK+Xz6Orr+Y/TddmiFiakZeawhD6r0QwQi1RBkeZg8wswGzskfd6g
aIanfEfbskr9YoXYlVBs7n7qujRApLK0waZUzZZw1kM5UJbfS7rztdbLPz3mTmjNYGm8P9PQf0/d
82VDv8Roqn71FaqtZPwICcWHYa5WLvpcHwpVJhMJb0phn8UAF7n6TviU7vve8W5/Wg9b2HLKfTVv
48iSYLiLhLVXd5pDRb4djTYxozUNpJHqpz+oCB3413xRzXz0hCAyYwab600ZZPSukqNriyOWaejG
d8atTjqSMA+uUrT1Iey6QlkrQgVli/7ne4GFjGuiuQCztp8qSX+cmUkKsHxL6QFs29103Kzc1zl8
uMGFxLQeYdbburtyFt5ufRusOMZ8BE1XG010NOz8BmTP+zpCwtWoA8pfwM6Ec6lUfAzUQUO55oGl
/IXtBkjME7cfaDy4akUmVLN2mtS3BgAeLDcdHLVeiQ82R5vdUvl5u6BfPkF9i41P+aC5ULP/ze7o
740EXBk/aOpI+eVyHeHASUXaiZC0whR/Y6bnki9/TxZqt+Bfl/70f7yVjWqh721haMmI+AXj1YO/
ZQ9BsvHhF3XUjC4HAYccymmcOtk0SceYqGUa9LjaF4gNUK3E9BU72eBU40JLa3DE+P8Ot3Tbb8iW
tQJf+IiHDfqwansTPftL7Y6bB5xatgbPMVJPnmmJaDzHM3DI+KjwHBH2D9ryVKacKgxRr220AhQF
7ylThbLMDJ1vWnksxpnpS9o5KxCKMAam9gU0eotmwcvH5Zh3UpJD6G/8EdB7IkdmDd+jQGlpBS6Z
NvhD6P5L11AOsTHu2g6FNAiwESXfDdseo28TE6VYtL9y0w1OTqD0Zx6xVHsDUckxDM0bOLD/9GLU
jA/CTvoBF533AKBR7Hn/qiySlWjZSkIdu/Td3CSPEGjG7tlbyq/QiHziGVK+5DBYv7rBkdlC6DMF
eE3X6IJGqZVQAasOF5/tjwwXsZ71o269FVd8pBGI9MRVhglsEGIchlaPExDZSEJ8aAmi3+kPbl7m
iLbAlLyhJitJ/8pYgbazyLmD/gdSWur0D6ng84sfLS7/2mZ1FmnAISp8GUCV/wq5JnKs84zJFdy8
ETVvqxctJfaNWjh6XSl8nDslFx08tNt4csG1ayAFgqXKkvUAq+oeYATpOTS7RCZHS7jXiJUU6lxV
XKaN6Qivl8xs8PMVgdeCfzjazONa/0adiCxvtd5w/1bPubX4q8SSsYDTtmkMAaKdUEEUKkspeE6c
sKOIoE3Aqq4qBhBCBGCh0hD9YRiplaX1RBWScUbIufXlWh5MG4dTaqhKQFpUF6mADxywyjL9n2o0
VaCJuRSfY0nlFDRRxSH1CPj0yj4dTzdEdUg2D4ee6A/rZr5JipOdFm+i1Vn9ioKX46pLxjYz9Ih7
mvlaQWQRTl7/cCLjdChM8DJUnOQaPay+eXRH2SHNAKvOZYY4b/7U+KLe5II5YFGa9LISgRf0LZ0D
1fG8qiTw20ExRfUBQUAN1BBQ2Pd1/jC54WFKTuRsTAARcSLomlFPW/blrEOmun2wKDadW/oveFAR
8PQSXYWsr0wvIQJXnasWAvCay6zbJ2WpFV+ZHeVJXndeWNemJ5df6NitJWfI/J8qGeW/7MldTDr3
xxwyOfmIp/zmmttwgBn0JsQ7LluMYK3TtEA4CKLTGz4LaYV12M9Yysfkaodb5Ae5xdxGWccz79zK
dRoF5D50pKYBMM5lny4XdqG9O2Gpq/viJxUAS2hXRGkiyKBfkS4IOASOAZxykKDuxkooqjJkKlhH
ix87u0xFtLrRRmleoxuQkvjfYgHd+V3T7vNqEI09PrbuTEcEc7z6jt3IOP7Hmue4gUh4ZOi/0dsE
R4fM5A8/nzyQtJY+anTKAuPIwSOtwE4TFuidPWEN8DQhqYqWrXMsfDgCN7mrBSsp5ErgI43GBvNC
fNea+nsFihFKnY5gsVXMfeFcfACv7IyQ/9E0jKKth78wG88+xJo8WiyDUijZKX4UcncCoFnYdA/2
zXAHlLtlvE8WF4Gx6+cYI0rZqpsLyhEXxAQfp0rQrlhV8r1A1827gegyyG6FTDgKrIyN957tNS7r
H9nGvGZ7DdzaDkh28EElt5Otj21emECtjC6r4jndLGkfndURPy6uJ990SqTHeGOO+UKpxkHDsmFy
wI0uY5pIlr7qRCCjSyV52fX82RG1ByPx21Tc64KdKQ6kKWT8O0yTWTy2wJNv4lAkaKDM1VoUhhXo
TurPjpxHsls8CTJ6u9DVGXdshMZjFsmvDzIVqjUhUw5gX12Op72iJjE/AYIXzrRkYKBbjv4YKOjt
lQEQVGAz4anoVy2aBjRDwLLIFWhzxjuDVxji1cU+vpRp7sBcHXsfaHz+64adNZGceTi0flfJnJIr
AgCWy2Ym3k9emnDRNfEp+paryxepawUXPwy4mbogHwoeXAhd0V/7H2bbcD8KkUzn0SOJ0v7624H5
sD36qpPReBb0H91YNMvZGCBUV7Sm4zbtW5sq8+8RpdeRkCLZaYawsP2LfttOC/uQuQ4JyDNP3ous
j+gxjMHkS584EBz2ArCg1dFCDHo2nh9KRNoWxnFmUqzeaPIFx2UOt67eqcbRYU+SCuvSAHHeUAmo
+hna4JYz3R/AjlqmZeez3V6DrqI7dw/kt9Y7Mpw6qu/XlkwAwclQorQ3+r9ql4HYfF6VwGnzrC2N
lHZqaLuOSM9DpyMDqtvJuemH7n+rCG2fCLvFzjLloGH8/75ZuhgLN6KFjD3xeU/dF5S1ICSo3jK3
H9tT9AMuL/g/0RTHniE688JK8l5YU1KKh+O/QPbRlzkXvKalGzGsxsP0t+mz9XiIDhUww5FjdAI4
A4l4kgm7DCtTvPVLL0JpLZopspG8bkMqwP4FzNJUvsfvkFw4O5Ico7S5ZM1kebqAVTDE0KqU5t4I
LX+BuGoDB2Gh9bbc2uCMTX24eDtVjyh6/UFe7dklHT0SNfIyo4HWkwXNUMUmfmC2KKmxITIzxK5g
Fo/BDHWeEQLOhtjhpdIj/ip9bU5JQYcXyBuR+RrbrAJabvSMvNkW/3OakcKjxxitYOomgjeRuXGI
nZSASVK/Xjoxd/81lgjefDHLcjV6rEHiubLY3WjUYWZDndcCGFp0PlnSLfnvJfETZcNHL8oGGGl4
ccCPEW7OWPp5Klfcsuw03hQfUyqZ2nV/pL0BjZuT+ftTwr37Vwq5nQxjgpkpHrG6vR3uINaP3wRd
c2+NgEiiLUfuTxkL1jkg6vQgaJQucZre6vDrSR2k6vmyxNNiZJRQul762P6VjAvwGQghL6JLjv0c
qU73JxGqWFhr4djH8lzfnRktuyT//YOvEo9FOXFlZLHPwvyv7yARaOB2WTtWOxYklzOQyi+XipaK
fAvKdf6cfrHogEKwCP8nqOhvcZhLAYDqXZ+88MQ5TBOQLINkwgtYNsyU0UhqgQa5DuiSPFZo3VRB
9NK4ejY2tKLNB41bmeMOaM7AT7VpbyzM0LO/rAZOt9OYJyvviQziBpE1Eaj5aKFvMAbiejwh7iFW
phJj2JWa8j9zfh5ccvKrW2e76UGaIokOrfoU8he1A8Vj/sKKbPluvrbVb1QUH7Z4RAM/AiL2QJvs
/QBEr5e2OG4tcNfwUuOEMQO13MATRDLu9ugs6eBEiTstwvveKwj8JoFMXqXgayMPIH3QKB6UVq56
Esm4ygb7wDucqOA8b0yPmcqSEThynKJJrnO7xzx00zoqN+Q3E7c2tcX68pUI2YhKo34vb+Dz8AgV
X2ZrocE6CB79auvPEy4OisqgX5K7taC+fuOlAmYACLBtuVWSSdGqt3uLksxjSnt1sJzBu7voh3z3
ODCK5MyABFuZc04zkcImBFElaWB1yIiDxVb9VBtzCyd3Atx8v9Q4H52DjAKjmA+JOay4Aa53Mzdo
aVBx09yX36xkdbdpOgem7+vb7q/AWj4Epx1xgVSkK1h+2+XKcWb1md6N603itB7TZc7ofO2Gq0to
ggWrTCsjMgsLtq1dwlaga/LFBvDlO1l5fECx5jG1HcO9pkeMkZ6DIWVNPXMxHj1QoSx0N5PXUcZO
XVeN4Mv60CVf1fgwFLmyT4us7I5Kb9EiFgeWkJdN2Z75dZSqD+jvIJdYSGBkaMktgtTOElePLU+Y
0W9c3WzCclCet4cKs/QBInzGl0PrexfuhXp2K5DBN7AUQrBZYoGB1r/vESHtluvYtLvwqSwZ9yeM
a+zod/KQmnDlECUVyxodVcHe3z1mZS2jxQN4EeY/6PeAjcKvBn/ZyopwC2Y5qCG9yNYqtfv7LvKg
7BQGHVOc6eZk671yG3Xr24CQb4+Jwp5DfBaNk/mvXSugzf3CsDrXfvdjAQBO/faQeeoGxIq0G4Ly
yhNKkSbIO3JLhm9fZybxvjh191mnkWdjqKB+GBh0SKzh8XuyGcyF1qzA3ZIzJ8e0Li/9dMJ4Czro
/+eKnIUJRdLkZoTZNgyuXT8pozLYv4rb60BoY0SvnDLxFbAseEwB1gsS4OmG8rnLe45NCJWc1fdQ
SpZA6zbZlkhWO7op4Aup/U2SJf+JWkx7r7822Yk5kkrbmo1F2MYBcchBTPhXJQsO4El1efYeyuSK
srFxevzOLpbB2+AEIE5Mic3sYRe7lkKjGbD87EAI5LSjcWoibqsXytAGkhTi2HPaT8SDNVUR6z/8
+xG03Krs3RJliNdDRjsSIN9sw/MAEwx18MY7Ly8mc8Z0nUWXOZRWAqmKM6P4GuRkZ/yOc88/Txuz
y9F/9QXD0gyy6ek86TwQ0cbe1TixUo35b5rlTWH9SUd1j6LYHqrAShquawBBZbk/rgLGE92eUNBZ
xNSQOhaSCg493qliPYIjHdguD632SsH1i2E4JZ5uEmghXRlGHLOSobxDUNGCHAPapponNC2V2gAg
Ycn7Bmz89E9Ct2dWhfM6cpaLx5WSrWVc0XRfMXiKzxUF1QlBQEP5TY6UywdmXZxVkd5Hj2TyZLRz
/GRyEwgIu3zlrILzRCV05OrFQycgIWHoPExZzhI6XUAWO2abRo1iZTi7TRtHp5ffyE4HLSa70KsJ
KtRyIr/Q/uCqcrFBqKekOfXD6JmEumatwAmh2c8DFPVBmgLj4lpjedxydYQsAsk+4zKY1KCsypoU
5lAfOtThKa5vrP6A0L4SdQSHLhqE9QgROAj5twe0caDHAhw/hW97TqiCS17Ci2ZYtDyE4O0ML4sl
tTicEJaKO5SW+rEcTuyldJdKIPJ66fW67weRaMIKbOrYImVW8PQtiRQhhTOFkls7JKxPZwCoNXv7
wP/c5QLDANpe9lVeBdhkAWf8tkk144a7Mvxrmayih1sNFWSg21YPskfbbX/ZAeBMcxufYSc+09fn
mQ9Y515uQYIXlrI5a/OQgHefHAF8pR8fuNie2hK2P7kfxIWKBccBSdnVrmHo4VHzUBCLOMKIHF9x
tsUH4jruSuPrdOD5rd6Yk07WiL/quORH/l5RQf03i27uPHs62mdSStmkt9BoUr74KhAXtPs7Hmlp
8vsfA2AX7EqwGB7AJ4Ydg4YdM9+sNusIBPhMt+O3Z8AcI4ds5M2ZoUSfFHpFFiad/cHqXhafd2z1
3WyM5ZhXVpcgbrmVczAtjyXHafln6WJIv0ahXduk4VTzKW13wG1Kb8Cb8P0gBtpjXu2cZ5NO6NEa
kRs5GstPvPRsNllK45+h2sWXd7vAxGMAnWgEfXX/rVci1NCUB/y+CyFYxGnY7fF1hZQnfaLaTPrE
1kh0eExjO+N35VLtxPtLBHMnKQfuqqxV7V9jFr/72TDVOmizGk4oz/FYvoAISj5rdocz7cKGFt6O
KIGyi+gwfj83KqyC911c4643XFjH7e/Z2ueMJLPdOxSl16y/tbJJeAgQAMOMqlEI0lu1hfUprf8z
JR+5D0DFJG5ckLPXHyezkhnb6UE1s5t2Lv2EgW+66H923SCbWJ/3IbsOKtLYN32R7T1PasSjSzV0
qh9xz3BPofk8463scVSmgHJAQs0BTJrYm/HRIx6fNvwGxglSvo3RRv53ODLrxZECrHwq628UK64H
s2ApNvIkqTxaA6i/+hRhCs3pV7Y11KL90+XX2naKzWMbnHDT7HDt3yY05g321Md3JYfwLIkCYH/P
finM6eNYZIh+JXnwdZ7LuRXruOXDlaCpPO7oKLNM9pUC4Wr207i/moQ4eawu0BEotWo3tX1SXDgX
cLhMPAPiJWaDRWyomx0fzV3ciHvGHYNSamsIgBBey8BvvWWhacdjbfhdOST6AzXtU48Ot5K6teH6
6Bru/8tqfSiJe93zNaxaJsUFhTZK20RWkzopphv1xdTumg4jCNLFof4YrTZESLENs9Nsf+DkY5IO
Ph+LnxDSZoEKDoQl52fmTBQab9J3xbHsgHE3EAI96czfVoOFgWa0ReuC734LXbxIWL2flrzrzP88
kLLtacDhNuBABpeuoI/Ehtb30AsrrxfxY+PmW+9oNrVEsYueNgj0iPHy1hrpT8hHC1M8jxuSYjUy
u5pJE2KIxCb2nDlZshY9hHiZPu2I8sglCsiBI/hsT8Kk+gsMxjgjpp/A+kwuso9RZEHs81sHqGiq
iw+RVanCx0c2SgxssqvNtOpNP/1+PDyP7AUohTmO1uGW/XW+80bWXwM6FcEBNz2379pbqfEQIKuu
F2qHgYkeJ+67b9xHWqma7+1ZL1tur52rrS06H4r5cH99nFFCoYNrUSwS0VUhehPo2LzOM7FfxMRz
9avqrF26V8CvKyai0j7B4M23SZjOG2p7I80yZNX/nWu6mHB1yG/vJLSEVjG9TXS60lmsBCVnMDQj
iFbeG9LNTr0GBMHCE5+NVy+jTdRYC88vjYwGhka/wc166IndaSssTmxqSNSmmEkpcDq15f6uwPkb
GPKnxie4eoArZrXjqAn/NSjTlZt2vuJDjOtoW8+hwjIQbPzNr1fgNksh0/SFJwvoS5PFyNOKkjhB
lhj/roJvSF/ibUPuTgJ0V7GMZbYQRlTG9A3d2TOhGxmnhQVc4oODflkqvgvNj1Pr38f5N3NDXuRR
wbG9HL3BJTkIUL6fjwt8FYbiSbSovQFAKM+P+WTm/GrSkxEICYmvmHFnCPfRqI2XPe9+y0Hljk0u
07W1vZPqWmmKznKL55REQLWXTimWPTgxhBgCN+2KbYdfIfino2SCBj3zvV1GfTND3bJumng6Kzmy
ASSWyfMDZDyLBmHJ3/KoeC6/3DmZwQwYsWPhfYaSKxfz7YJBqquTsvdrUB0Vbic/f2N4euOhVmSq
GyFYJIjoLp6b7f5C3JGVhpEyL+XWCgqYI1boHSwShfxIx7WJHrX7Fokw6KfACAGszoGGC6VvR2dk
XCH+O4dZ3u0WYWBDkV0VPgNEJRIMiaTv88F+VYfd9RTFkMxPaqnmvnH1Qb6QUJKP/882BejmXGAN
cCixzkw7tgh6ETSH9lKMhwMLsfAmQ1Wf/vFbYpWGfYrrPjIGRJtaN30zrh8nFIvRA7O73NS79atA
WgTbqzfksjh3b40hUNud1HR638Be/DXsGd9VwbENHin5ib6DTtK415zIYR+0QqXZixu6+FaBdByp
YFLpy+i73uFqxSEn2XD1JVuT8rINU0leh1dvxXiMMm/nJKZXKYgF8IPZpF3tlBIMMvA4cxrvo+Qq
Vo9Vgi6ELSElF4/y6ojKhIrpxjjF/jBpHeL7CWDD6yn4hRfBPGBtie375jjbRdhcwDrMc0qXT7wL
2sNHtOkQgaZ/4b77eicdgheQLEpvhHWrMZumpsiIiaDlM0Z50sLdgfKlWDCHiSyNm6/RnANqHBM3
8f97MZymupWjHof6ult5T998MKwE97ywqztJW91LDXO0rZRiVWEsBTsgvgf6/Il/2fNS0JjRhABW
x33MvbmnSnQ6IUTLajNxbivn9LQWPnV4XE3NxHqZVKY6afj7I5Gjx6xcOTHKYvOf5wIpjTTVDpc7
PYI1E2CtMQkzLdeuSvVmVFh9T4BMj2kl9VnP6tqAHDCM4txPvjV+9eKG1FJtsq1/Ut0ZTbbICqhM
xqg8G/6CXO70pUgRGzJ/9FP9bBe5F+aDgpxQa4eWKq4Kg2NU2ZIVhTx2bLyitCDSX4B1zOBni4Sr
3fVZc0nqHVmihjOoS0VtgyFbSHZxnCLR59+lz3XeE1xr9WMxbhrzy7Iipfn/UMqaURMmKmzTRikS
iM5RGzrh15BPYRdrvnujUckANOcv2TMKx1cJqI5uR2+Qv5NNKzaO8+GqVyfSv231K+TmtWmkAwdq
ZwGvi/4YNQp1xfg+sRJ8DarNGaNxuaec/tuuGl/KN8xpUt+vMUBj6MRU4xP58fhHRbPdAmOgInJX
gVjUkw3y6hpadPB0+TtIinmsA+KSxjJe6HEAXKqlUAr61ttE4EI0lDl6TpV9mMgmhVUalumWadmU
GDeDuCNMLMv7cS5MypyvYdqYOjhTz+23YcXUBrC5h/11is9upPPiUMc96ACShcbVqKSPYR4ksLTe
AXsUPWRo7RPvLYANvdtvmw1nRWjh5THAl3zjyZfW5FzfUOdcAH1Qif5kpq0zltV1N4ycGaHGwY7k
avdrQDy3nndleMVl1n/wKF7zmDX69FVtTYISyXVHSAUWlS2coBn+TvZagcN/QGMGpzZYjgr9lYpL
kyrzg+2V+LWaOXh7dXacfVYPXcMlqEoHgny+ncQy5pIo/6fk2yLGLq5yDDyDXCABzDTuhusOkjz8
NxBa6HCRXPVoiABQ6LbrpKzkqMVrsOeECegVngZQvZWyjntCKGt8+/a15CyaJIfPakkMNGQPZQX/
Lx413EK4ULepwJ8lVx8BvcKBcE/5wUaf9AFLpspxSXndHUoZ4sFXpwjrMxBC9EAZgb5Ni0mhCOy9
4UPgPLtfTORxtm17yRmV2utTaH3gCH9dqmXRw7N0l3h5e+QMylmy5ibwbA7kyXtcAPHuLb3CZnrr
0vyJtSjY5GsV0z7GfGnbeyudRmPIfqHYo3JUEt8tRcZljaZZ/MbD/TnAFJWkMJTpv7eSzzROoJNE
xAnHLdLOS2DR0Bhc5uME0A3gCez30GYIn+ArMJ5quqzY4Ga6p8YqqQmX4LIxzaV9vNh0jOW3fy9+
LQZhjoVqYGzzonHxaCpNWQNjU/X79IC2lxFiQs3yT7pWRjV7k1rv5iz73YKqXFNKQvkJy2tQlhE/
xcWZQxsGUElNnyyokR5L+BcO+MZ+QcD+79fCkF9Js+kdFaLI474L45zzx4dQ4GaJp8e0yFGTH2SR
iQbKyUAxMbZO2G+NJG3XecZRE/VID2/Hx+ARNMMhRDbN52jMDXoFJEf4Dxkhy4NGliVS89HhKo8B
+TE143z/W4UbEFs6vMkkOUv0OZ3s5nQ3sUPNmeTn2tCK6Sbx0BQsvD5HdNPTx+rHttaNKnWSsztm
zQIYyGVnLc6HkzQNcLKM1HVjXH9decKKxZHFWobuiT/Fl2u+g/3PIUb01JepS9CdsAKagE7c3Rze
b3TU9jAOBWgMtkNjI4uwKSEkpuqU8ijBlcJjoGIedQtLnEy0qA77Kozjlehmx+fyesslvjQDnEiq
Yo15De7TOqzb02GY9PvIjuw/NqEQcTMovBrg7PUaJQpZAfrTJx/mdNpr7Y471oFyqbyiAyt/QWVO
fWoDI80vq7Pjc/jg+xqsRn28nDs3XwALJT9NHkiI9Bjy7/3vRzGxkly/c6x1r0AXwfOgTlyzxRMm
0Wrv4mwPgiCRiJN/iIAExo4fXX/AXz19/p/w7XhC7iey0hADKDYTYbWb02/ebcMq5dKn9wUTzFI7
WDL1fxYfuDrK98XhjD9O9GL4xDgs/025qZIUlwLzISGi206DpP3NtdnxI/k0FvlZPIxiUJ5ssvAN
n+79zVWInJpuD8y4Z0s3Kzf4ejAguYaMRc9ccFlD7HfdU8fuaVlu6omxZ41p/kToCG0wXjCoZDYh
Va18h1uZjYqpeTL9OpS9t2a944k50X+WMiZ1jYJgEjjkmz1SEciGqAj3ZCPa+dSR0AF66Y03Ni31
ju9N1SoZEt3N13rKcXb17a8xJHtLbdFr3VT6xiI6LM0kc9XGDkO5SgdBt+3XDqZ2bfXaUT8f4ixB
+GxG1HY2eVssn0SBht1urRkkqRsqqeGupI3HQuzhXpTWvokWyFoTlFNa8gyAngjIXfrwpdG+l/0U
CO90rfReyeT0TM+SyXpfLLYtOFyfhVe/dUkcvwBoB68N7DbJMbsahwcyN3KviYpsM5yI4EkqSFWO
Vn0vacE+8PczqjFk1SggxTXQiiSo/ujGa4UctP1lnM+ykQu/J8t5r+BsncnGNgDIvAGzxYPPy0ND
vxFg8eVf7v04xj/xmGEYBVn7mgU8AFLKEcMLf51K+Znckyw+1kFX4H3NflmtWp8/z5qm6o69gAEW
ebrKKbodcduQU8+5J0eNR2bc4zObZqY2p0YFSqDlexSUf717VLdlU3zMBHGzCWacRQuXRiJsxwJQ
xeObtx/uXCeNukgsbeqg+wlmjA1EJGWURXhOHLk3g3dDKvOeFEBg61Yh2tpcuCupNZs+EuDxgu1E
Yl6E+69Qc3X76bwa/NJE+TFzmUBEqEhwGUBaOHBL7oOPLZrD2eY2wkmrtRVPO0N4dbHQN5IJIbHS
H7n2a3fvmO4FDUwOhiFpJe+fChe1ivQUmtG41YVPKaBNkNcDfOmJbARA55fdkcIJq7HLJ6M/VFzH
7H4EZW880m3UtHkhXkjBo1WxKFyEqPSYBuGyeFIMdb6hf39wAqAGUZCPtEuCwk/l8UBWczBDb/a0
OIELef2wdIou0YGcVWuog9m43vudEvJAuknmydJYCOVf3PD4M0Ov9L15qOZzjLU0b/roDRi2nchY
d+0XFSN0XeY+mSFYYOOdMGLlu2RvsiWpJvQYIKpC14Dcpsw1fQmtzCHWZD0PwjNou2s7+WCEQlOr
tVD63MX+96n2CA/NOQgFVPCTinjqb5UQZs3hGMIuC01/QKNiKjD+JkCB4u7QD5eMNK9BFfYgAHS/
fXFjxbyGwbbfBcg4gPn0Qp9cz0X2jET2Dfz2UgrCxa0l9rSy2eZCRTVhmjkSMUYJm/8l09ru33A6
UKpYKyyRKo17rDmwEE1mZUXT9FmZS/g17D55DXAE25Jr/bHAMbVzk54Jnrecz6RssnqeoMdz1LeV
N8HBjX+2lI+Unnmq55w6DSBl9LVJ61uLt6DrHCkpyfXCQTK4cZtnPObVSxZZ1PRJ/QRdY4ZTfKeO
3r8xb+0sY0OjhXPub3xSniYsvyN6VatXP5x+D0kek3rUddjpO3FB+D6w8orGT/TuGvyDNPpHtERZ
RAkb6bHwIi9T1kE8FcdARFx272le1XI8gfOErNam+sdF61a4j6U/65CYlhGnfL9QnOImEezZMcJe
rkRRprD0OI7Y0s6hv4z40V/6MJxwpfvK4NJ3IetIspZuHsx5uyqgIjiDM5IHHfBJB9+6esF+AWlz
HF9KEa3KXRaLoVEF+4OXlKkwqiifjJvCd3myGb08hVnU7PGioQl2cK1tTBp/uUwuuJeJH1Ggyiso
eL1u8x63/OVk9eovZ1YgkCzS382PrO5lP5ofebDkmxFTE1NhSw6XckBHd2/gDoTtnzsm3JJAyTo9
K+92vLCNs+BjNJC841M1SM8GtASLuZ9PqRYlQ8/pFuz3gBCNDWCh+qAhj9yQt1u7lD4J6Foqr9cy
vuXgl1y9zxc8JPABTMchKJsDY7N00M34mEri4q571RONg+fK1B/LYwzrCIzdAXgbsK9KL80FPoYh
lD6V6BbpAn66jpQny5eGEWzN0IQ5hJDBaNOdgjGlZ/ppDxnGjsktk2PdYJBdLncYQm4B37Ufp44m
LvE5mxl5syyjPxSz976EVgb8pJPtxselC3fRTULVgRpvUoFKcWhA5Ahn2jqxyWCs5P3qYbcRXcin
InLHdzUkHSWqrHY8fUrDK6mggqyXGuE2il6tB0iyHHkCuKbat7LGNtRgWPWeAn6n+pq/bamFCXaM
St3IEDHuhpbKTvxmxiEX33HE96Gs6gIc7rvs9MhdpSmID1QPDPyILWH5u6CFRQtBOf9muyZ0++1Y
nvYIccuwsjGReAI0dB5tE2X94+SpEiJA/W1f4MqkfhW7PcR4wtOCbVv5XmSgcHtvybsUXx9Q7m7r
juOmaBsB2xvRA4ZG64jI35pjjZ94SyX/S7eGZbUOeix0D1u9Abgmqrjj9upl1PI9Fa3okmMWynQC
si9DRMtX74NAjwuXQ6DzUr1a6584DDcpwZfyg/1EZuVmldcQqmd9Hjr5795+aBG/cse2BoO3bNnu
kqh1SRFtw/AbBIPIlX/1eXo/QdezSpODiM3mRYQGuThwKBKvgP1Me0ciCzCyUdZkNaj2UJYPzqzh
1utwCG0tFj8mJr6aa7GqRfAPNbInhsDisqs0V/3coCrw5Yb13UELUlcGJ9jxnhBnCx0R5tKUwkf6
onsXbozowXLMwMQydAStqKWVsVP7eQ/Z/fa8or8gdrCf0shlcX5tgHrvgMKUN2S5daCTj89Lb/vJ
MgU45q7Px7FsZMVWEpDzA3FWUWI4F27SEkxW7AEoX8bf1zew0CgI9AD49P0INpMGnsMBybPrBkUI
QVdrfgm2waDeahShL+fQHMkWtP5NrHfRTrsmXO7Gu8Frm56uFL85Tnn/RAeLJ74YHk1GX3Yt/I6A
OPPexGBaT/SZmoq34C1F033QAxrsBg9fOtA2ATz4lYIvyy3hYYiEX64KkewWoP8+j19zpqWwXd3E
FarGjl++4k26H9wrYDBKBTG+hmZFDNvyQzu/rFg5On3O5aPELGnD42ROwzAGRKJVdDBVcwZNf4bW
wek8w/FpyPfGiWPy6MekS7zDJGmUvPBj3ZbB8AIoV4vxvLYI/l4vn3C6sqIbgETGxivuTiCS9D4W
etTOV/Xgm4N2Nxj/6Gd1uLjeRCK1hN7EMoDCj0BM+P7EUmrl52qw4PeLF6hGidJIPCJF2X99Radb
bskAKriHqtVin2ORfotbyFPl9HbXlePS4wp1SL0MOqel31CRCFg+TG7fo6w58R4s9QoL0j8G7/ho
lfoTQ4rWD7FmhJlOtipeZ2jFuregConiI2AN+psOHklDKQS7LevPLeG7DpBLO+fA4hDe8F4DIZ1b
UXjIXXZaOPS8TdyhHc7nKPUCx4KRhevWHPKV7zBJ7zQk2oIdO+IsuwgVXs/0YLm34VdvmV252qxu
Qj/DeaK0ziOPzZl/dkxWE51Pv2TBcg3apL+MXBV9hGGAr9SA/Pxl3kJDO6pqQSTeBdTb4cUx6+k0
7JjB4pMAy4SHotdYoCRpd8M/DQzwVZ46V8znJVa9n3+0qn75wskQIXelVW4ZDMAOEuGNpuiYSi6H
5ZLipwJ4gt1yI+QQxFwHOGabhOIMxhYfXmSCiektQuH8WLeRxDBBnQdzEk44H7pRVt2NXBcQ/BQi
P/WJLYFBbGJIhSFXifbn9c5NnxN2bdhJXa1kEM5oRhN6sDZ3BRHjOkBYdtFsLcNawceJX82V9Ogu
VziuxT7fASeBvFmj4A6kBI8phpg3RpwTrfK9NF/8y/1G9MfKPUr579WrDNtt7n8FM1dknaYzVoTt
WGYcB+9kxqPW+ho8PWr87NR5XarOX40Ct/Obm/Fg7fwW3PxINdP0tqEGLsyhFMFq05R+OvoBQcDS
S341EQHdnRzWri8e4FP1+hlIVn4hEO1iIRE4pmU1VAtOuD0Kfp4LHY576mrNUIFUwj8zFFcyJUiS
v5ZAM283m7PPr0BR5UB6oQulsyI12jA9nFTfUErsWXCA5b6hb3RKx2fnqD3ERCu279fDDxncbM/z
4OUfQhtLmGi+vif5WoUB0xDfqKEVCFZFLelzIuIx2Nbzqv7kTR9ISAkLaBIHnto9vNBxor96/Cf/
jzx4MzMKSmHG3RmId2uEs3kRS1n2VRy7GGAXCb1Jqh2cnUuUbSJHlk8Mdy5tin4FzkPS7ll8wYJF
In1WUETj+H/OLguoMBBbh8E6Up1AvREqYGuMwtMsuZEsnNLT45GyayLv0bVkGi5HAZysdraR3BVW
tZbH+d4IbxjNYa8ti1sP7kvHlyh9hsphVi+p9sqTpWqAJPKF5Lc2tOBIwHGOtYtsYuTRfvWUsT7S
cXgwpb1dOktK94K41HNQk8YJO2b2nqv7qz84rQcaavMpK7UjyLRj5E+TslCIPhIEYKS1q5kX8i1R
4WmHluwR4BVtwgb6uONYBLROdlVvQVLIlJ51xf3IIIdCmpSJ5jGzva20MENmfhmdA+xIGVfvDwrJ
/XC5nReUHbRADSboRY9EaYQzdPM4P2sAVBxvFfORb+5OgcMYbOi6JhcqcESgBoX0JogDOSlL+TIu
4DQjVOYU9CMCsp7WFpUz2CN6QfkkwXDS+VxtmoJzIhU2oQULIYOyCIInFnA4SkUliXBfKRRodoUf
UuU+eZYHeiiQ5R8jlLJR0HmLXhANYpCHIgNhLHhwHapLU3tk+yDe421aBxN1XCQOT+X8nppv7Bvz
dNgnMoPvvVv+W2YiGx+iMGgsDpON9vGsTNNrmpbUVGOtKrWp07prUzohxB4pr3I4/g2J7/yis6T1
YxySUMHYi9q/v07Nyw0Vb1Ngm7ZSi/ys0epz1KCz0vDKUUc7ylXssTVvooIjmrctiAUJTJLajWau
ghC4RwVuHPpSDkT5toaRcV9iUPg6FTVObrgMXi+I1XXKh1B0fectFrEspyzbhNDCOeNqnmdzYYke
bFxMh2U/NLGqa5ptpj+kJAFPV+Gk8XpA+1GkTL8zsTuvRnUpKPPR9Jnt+U3sW0ToT9KEZ2Fqv2xg
e1IQF5M3i5VoL0xgdm1Y10W0FPnsWMkL08XJVzeKDLYZaxX02d+Rui9uqWRDDUpjETYy3xreQlGU
nAeKbRRuIskiDrHttaQvTwNh3FdZ0wXcwUcPxdsanq69ABrspGSgYweZm8Z4GZ4J+tZtkzvtrws7
E4ELIYSKI2wVNZHF5JyYFVkVQxarIQjFddiYlC1rXy0hpNZeUszHIsHyXi8oF1gVNgtzDuF+qoZc
fv2c7Ex001sNZBzKAFeMC32uXNTF+ec/j1x+JWrztPnEunHpLH+tgtoRk11gyzJxkiV8o6ER7u3e
0AQr0etKXZh8M4661er6BBORRmTIHsJw1Pc608Q3dC5Hu2u7ixS9ahaKSU9dhLDeaoazq3npYTui
VZeXLGVs5f0+t1KG5n+sSlkZ83XcXUu08BJ+fBntLHtzAh3ybJDwH8KhipLVLlKCjjzE1YXhijlM
jygB77Vt8FiOn42rlczY18OyWyb7ZmZDHpFeZRNWKabDblGJgAy9huGLkbNPjVL8VDCEb6L+J6V+
mYuLmAIWAcQIEbRFgcBVaoaAbCJmSq2vwur9qFlIbLko+D5tYY3rImMppSYrjuJtO3bsZehoyg08
xHfL81EZOeHPpfPCcvb+JwvE/K7hMOhxh6QUy92+W2RcJiwNYnU98Lui+DIHq66orM6pbE9I2hiV
W6fpVAOApN5sBpgtBA5dMmwDasjEMdUC7cj7j4+Tv9gYXWH969YaWsMq2f07OZLdvlMSTFtI32gQ
k35YSMqcSta9DFe2x5dOKtoPTiGgOwjOqVKtFRTJTToK1TC3d4k/Zn2/49eBTldN2EzOlBP6V4N4
m8mhHc3X5GxuEwjAWo5CrUvc0PMQnQUZfAQ1P7xDnRVRbBCfxCFpER8ZjhShhx6mFL3nh+Nvy58b
ZJtDBAd6T9+gq+IbSXIfFyDBU0nBMbv7azQubbmZoH5c11nb4kM7SkxuRKQDtOPd0BujgdvrZIoo
N5XBlQvbw+SSUfBDHCSqAeYEERo0lZko2DSl5ihlu/CVVkEv2fCkLOXAhGDDs+bKKiTugCIVfTLx
Rqddd5aB2apuM0NDejf+Zb44QQ23hxBkmCEVfYW2ffzknINrU4bb6gPXEwPCBJY756dayXA/3T94
JhUZr0Pi+kDDWhwWdd025hZGlyXw7+G4dedoejNmYa/DBpgXfq1RFvAl0h9/RXRCuE6jNEHAo1if
JqsPzEYP9eKJHNvsAEUVJQvLXFw2Kx3Vu9JHMZJoV2Ec2GkQNwl0hCi6P7kQx5IU9R3VNS/+AnYh
9SqES7pTAYvdbd7abYvOQR+HO79XcS+yv+CXGX8fFzTAT6qicjXIeMpAuPfosJdrJn5u1Fp++Y2v
c8zHynyD5CuZ/QA+TxTzrSB7U2HdwiTdNpZprJDRzX29zMgQYSZ/Z2+YKnhezo0NJaY3fbdJViOL
3g11aaL41ih8Uo8X8Oq9Wr9uQY2mbIrmhiULJwxt5gLQgWWlFVll8v2k5zvBcEDoWtRymhFP/1Ee
1J6R/QHyaXI2/Aq/6VeaKwAlD60aj2Awv0VDfoOPSk4+1kZd0puN4l/bbeKQRydZP4dyp9HWuFEX
2R+OGp4joXOtKnAjaIDgMazc2MF+K5cTtAR8yghU5UNlA0C8/N1Izkuss1jcATdnh0c30iibjsG4
3JtOYXgl+/tjryZfhAHOwVkkd86ETqGlVUlP50pbsejXr0uw3MjH93EZDAoDme89OjA+35ICopJJ
GrNFM5odM2q6cRsZH6Q7nKD1A2YiE2oaoEmKtlQrKM0AFQHS/CG+tue5cFttDa0/eCtVG8xmO6nO
XYE2zqm/Z455W44zwBJK1ZDfgLgWg1nxNDGIn1mlEwLOxBKItCPPNUNpJ5B+TKRcaSUNLjmtv/oK
0bzuvTcI87yp3cNtKo+RebUgAFfMshD33v/YHbfRcBrMl4yKKVJqDJ6tleEkgE7pygbJMBZLNzvt
3Z/4plEEjObF3f1+xjozCPfOGng0nbIqcDTNrlZ0IhNK/cFuXrDLpi9vLUo0JWTjeAt/6+qneQIm
XQEXxyf1sML++hp+dDkG5ZfJuPkctpduu76Jpb20MaVDcLOD4DjOFirPfAVRp0G3V1luvNmWiTw0
g4dUWCEDLyRbJM6HhUSrFkmYjYVJdyrT7Y2L75ra84QslG1s0qNxQPY//LWJ0Xfoc+JJjf8E5WBu
FT7wHuECcFhirm+y6nwOayfgd/xNxCgEGzPAm3LHukPXCMo7XjpTXYlqHf3fawgzvk7E02EdDpvM
HPoPJiLJDfPTWRl6M1KAGJLb5sSakLjaK53iVwBTOjS1/ct7lJjVgKbcmNlOwsmMyURiIFj20JKR
Q4gVmaxmw2GEIRuT2v3pck1QtrQYbuTsmhUUICY6OKw4WW3PeCHbzSeBzNC/a65ELlgcy6cITfkG
EsMrHaq+i2ffF8NftSOalaNdg7/i2EIb4ojwJj/jX6+JbRE17qmJP8fv2+Eb5FQxjHcneTuHQ8W0
vGrKAtL9OhdRjzg79ndOXSOdqpNAIitTNQS9aoWGFyA2bz8iLoL6RUKVSewsBPzSviuZfIfPTuhN
wn38Ts+AC76SzBi7sgcxETZGezPh6ji7o2ut6bTXw0XDuOfQGCiIUsOYtzh6Fb0xRjJ1EIVYv+Vn
03BN0vRXip0RDQOaaRhVVjwcsTrHITMp1zWI++IQ3WX4rTOHCAsPpSfKyE4xv5/OVkiIQrgYwWxw
wxWipzunp4CO1rLgt6h9IqYaLfAEU/Zqcoqmaxg+HWOopERX1v/vgn45qlUiA8kPwNnGKdtlwlKy
8SswcvImoaW0rF8eRZwTDNqRm7PlPT1fw1Sj5z4UZRyZLUXZsb3reE5hEIOdOTpRt1yvVVSJ6ZCU
THvyOK7ziX3pAJsfcgsttiwwAIxba2ORbKWyTHRs6LvOWTx3TxjNK6i2/gR1gP8LH7zC65qkxTBl
Zl98oT01Szn1Mbga1IqOnOEZfZSCeNsLSw738HfK4UdTSWkVZGrT1j5aqr3B+5A9mfu1EdWdqAiZ
wf1iu5Ww2sQz7frsA+QRko7X42mMyfIiw7Qx82uzAsbArDRH97Om1P4hFlc0yVxR/QZzE3AESAb+
Falw95Yre+2xbotwNEGKFhh4T2kH8F4RYdD5rtqPAKeUVz8K1FU/ULSDCLnbk1il/gIWk6jhzGJJ
HqDI/LuqpGcb+pOnjRzzKg/pRBpyzBSp8zVcGVioYxXoWKlqq2g6zXtsVn+KdAXp6ukjhr5e9ssl
LA1WCMq3LVyQYteMPya2MWlfoSBIVpC44kI6ASVJlJCZ7ikR1I3W8oSJMDjltirx1ZA/bc289eaG
RyT3G1kSHX5n6bxbjx8zBHtctLbILit/zxKiTPHPd++5JdeMCzeNAabxzxLfbwsn8nIDjkP/hQa4
WqyaOGBtgM9EzdUSOWiafHpU5ry40WFGGaFP8ptigJSfN7j6NnzPz+Fgf+Kiobvgl0giILHsOaWq
j8zqd8p5EWdVrHHWL1IGuNXubrcsMxkFvLb4Wb1zfIr1Hl/khqH7moR5lQ3fne6bJ4Z5HpdYbh65
SI8JS64bfEg6/eyoUHFHFsQmTn6itcBG2cyD8pRIDFAkW/xly5wa/TGP9bmxHn+5KpSM95CXy59I
jUxPqXbAZzGBtyTK1BCCCQzZOrDlmiBlvyGdy9ZKEeHeMm2oBDOAXoh22h+wlsLB7T/LXfYdGuOX
LAWrr4M2ZAnt2nu08nEYEIQV93im32GjGwh7J/vv1yqkYvT4NKoWehaOe0fH/D2lrbhp9a+wuOhl
WvWqvuFumUzplW4sz0P2uACbGn/SixDlrXcVwk+hscJB5xFml3x3Y4fQg/Q4d/IEQJdGFCvoF5No
3TCZ6l37gmjupv9RTX4m0pQjF37nd/mNnY8pYy9NBynv6B1+j8b0HBYEb7kRf7KirxB6EhzzR5kj
a6S8B/ZKET6H2HTFq72uqfk2Tj3Kt7X5rP6JxTUzziows48NOWB5oXf9MDU4/6O1x0bBEMMDKYRe
w0/NrAyQfeXr91AbJKkACAj98PzYIHHeGnTReZX4V5Yx5+EVrkkXFcMeM110QOjzxgXgqkaEyqsN
M+Lkvu2lEtO1GAjQ3yhAE7S+q9RFX3a8w4rVJ9ENNOvmELem+akckRfA2cvLZuU2Rb3kFZK8u178
teYTwQsAchHnp32J85K1ntAIyFtbq42lDKN6lc0F3BUsizD9Nu551noyZgQAQ03AW1e1oKBNck/M
F9oEOCHw9aODVvS12Rp/MSpDciuzmJ5lmnG5FWkubVZU4O9nuJED+QYxNwZDek1Z6yBYHPPqjmXU
QZ0UjJon+M9tTo3GNprA5YhCr9SMLUIEy9WrEaLZRD6AqAbgmUj5P/xIeWUeAEfm9meecyfApmOD
gbHSG/SOefs1bW8MDtSnSIsA0AguUoAzwRTl50EBp5v5UEfH1hHsvU/eNEKteFc7mFnPIJ5tvLWJ
D1VLNJGKwFAqnZs77+CHV+t50DIxHbvA6giUmlwSvACZ3Ha1LDcTz9L6ZeqVMJPdXZWNwIWlfFQV
rNti07+oi6/GHYW/bdjpVnPSsNlU/euMZ66qEzMxfQA5h0/XGO4neoXMbXgDqNpYFIk8SD6rBEVz
Iq0B7z6/xaXXAImxIbLFWM1DV2s3LeJDmSsNFbnk2bm7EuJibVEvjO5bQs39PmhoqO/o6wPxSevS
MU6/nBs/97vNnSEB/G64pCJsUnNi60Sg+vpEqY08v/sdpxVLKMnDXOt6anz/NzoHIZmuO//roIXZ
QeLvEGLclLhDKOa+eLzwhKgq6YvX/xz3egN2X35ViRV0F6iOsVbCv2wL622UNdc/saFMTu9cvNVS
W35tsv5RAMfLcX7nhHyEgAAy5PROWGtoVcr5jyTujXo+JkqBtvJytd75Bbw6xvCKcavwnjPhyWhZ
S0dlFqZVJ06lItfJjmCVA0PcYjxzKiM07DXI6DAVe4it3aG4gvNiohyT/GXSsAnkD9We+kIcSd1a
+SaRiZKa2doX8kheZo6wncM0g7E6VREA1sscJDkaScmnoPbUxe59Fi78a6ZNnX9iDbCxVOBQnnRP
DTjZt2uhoU1beiTAQoAFwW+gyHmywoZiyETfgcXjU818wavkCJdrMCzlCgshPyeDVGhjCoTKWpPO
tYMuyNKJ+KYgsPAXMXn3aP0OWoPtpGAxWpxQgEGyVSR0UY7tz+IrettT1sp1Tio4NqW/eTAdUxz+
pDC5y8SxtNrfm5K2x3iLcnOfI76rpUWFR8wGJ0Y/WI5NrRw/VZ9kzPoOUbFgm2wH/6VU7yYJofdP
la9l3rsf6e0e41GsAPvk5EeEQBItnkz3MPAhBXtTg5JogEWDmv2EuaHyWwxGsDapzLljIpdIKs1S
8l+Vcpbpcvp8Oy2BWmBCCvAwA9l6QSGQecVGeK8wuAAoo9dlhyJxYunYhN6Y00YmGVpWWL1eZBZK
ZN/1SzaNhdqTJQVzNa307kJfIOKuVovQGK6XYzuUmUCxgZExi22W7JnSCDjL1HwJLyXG52PANIdk
ypgsnSaPRovEq5peUeUJRYjOaIWC+e/W6gSuBlRoN4C8TCJkXJtCLQvXson1dzU1rX22eNmSAbzM
424uqMrufx/aMFYsrw7ZG458cJx8zFL1MwzWT/bbMQkjXJd44gDZcgq/pcnNBKYA3x8++UoTwd1x
qNFe70K6ZME97sDc9L271ZYCdSnc6cMBmRLYKeoLi39M2A3jWo7d6xa4uVyRoyZx3Ir27g6Ll+pB
/jJtS0aF6dUrZcFa+31BpPQ4MYMscDvW5M+046oHwBgqD8bDdX9Bl4CX3MnnguxHu5z3gUXx3fkK
3b4fc5QPGcoUUqrCJMRXJwmwlhBlFqRnqHaB6LWQew7KaRmF2k9p6KzRben9WYZAQxc2PQLKJIfj
yO+avSuhFrRj+w7XppvzOOKdmxj07IQrWX1CTsJofsdtdWbntEJ7bhlvoEa2Q06jKlccybm95X1S
Zx7LgAm/Jdgd1T5qEjYwjx7OBkWTOLzJckX6hiSRR8RGaWOwBtJoU0P68d8a7CgwzbEictjbNZ5L
BNMJLaewQl3Ns+7MV/7PzIITqEOVmW/S8RXwzDkcMah1YdiKFOVq1d+HRjN1GEsoQqLjuSxoZPrS
ylooiVa8ExOfxSMOlEUD+Iv0eAA10szAd3girfmUmpP/Ox/DoZdvxtGqrYkJpBzvBKcfO57bNbCa
Wg9JVmT3p+nFUAL/p+dNt0MamsA17RUWpo4/fMukWjERfhYCGvcAJr/2+IiLEnuliNExbOgIMOvR
xGQDFuSTYtPkmt02u+9DEI0qVzrG4xnvy4fKLCDlAQi6hdKhAvYx1DCArWthMccM4MH29QXl8M4E
gnoa7co40VRtV/7I/8wwKGcIEHRdKDLC8rczipyA5b/krWDujaouYiZTPcTXZxE1bq58M5t2SbZf
JxYJgkz0Tro92D9FSgpu2lJHhwy3X8NinC3lM1gPnaaMvKvjjEmZwQonNBFoI9ItOagyixrVFWCp
lLgD/WGV4W1IQtw/Sv/M2YdnIGXeW8H7v3XrF9fPTC5E8mOj/sIDvO/ltai18/Y7Ltz3MCI26iXw
Gk4opZlNhLxP0AQ0VpcmpxSpmmgBk0NzQCdqY97S3UXBj52FnHBgCz3GPYPmzTiThfxWDVIHJECF
j0AmBLB7Pbd1xx0toFFTw5yDBHImkc5wAG2Tq5L9rBkBg7cNP5poNZSA91Cby+XVrLPEFdkzZMTn
jApVimkG7GGahi2TuE3Lgb5R5m/P6ucojBPJnvGZgeOTjndN1oDZa8b/eMHsA3w0MrsvgNQPIlyi
QFfxwtGuQmP97/fmZGLxQoJj8oO/ybFU8t3c9ae2HuT8HfxUbescCCQePhboYk2qmuuojdm1IGCy
T4keMcqpRo/n2SnOwFAdVGkIkuIAdbL0ChRnOT/gjnPIIa3foJg/jpkajWkiQo03a7NO1CaIjy0j
jnWpzLyGbFWB2qfhGJcSqfDMjaVYg6Ra03qxlidv7ANqeZ1E1YNrNwriVqDu+MkXhDJZtN+HWpW5
wp8soL7IDFJ5EgJQRryYAKkZJJsdchUoniUA7XFFdAzTu9DAhkjZjdJlRVkrbppvBoJC1ZeyefWz
AI127J4eO2EEXDxeqwTyQaFNdUk1V2rLLDF64ZkTF2ZTl4PFtzfWYziD/BdBvasmfwLaQ9wpgCYH
7Za8RNr4wujf1D8hZqLVEB6zzH3jbi3m2wrz9uwGwtxOjFqx5NkDm04NFaadIPC4KptvXjgN+ajw
NlQIEaea1pvMZwohfMv19+bUmziVXrLC0FoaNbKzgFj8NhyullxL60vuI2mV56UQ8xdaQGnuzeeL
9o3SHW0ocIcnlt0ElhT1FVaJVBHkEFo8Lw8bZ7vsTTvl3yN17l8uRCRa5ZHldOV6rZ+o+AcOYclV
ykbf0WmavpRzeoHwa1LpYuphbgC8dahzKFJhMkhnuewwhQD0J7pOZZxhhOkaPBKftXWq/zDBgobo
NjSfbdx6oZAoQabSod605vLjLpJ3wYKcL63WvW/RAmqJlLcJs1q/SReWFZ84YFIDNUHxiYKXoafq
d0LAA4RhI2yck1e94f88uro6pqangv2yrvkMU2G+1HHzsHhuc4j9DdCxQhMMi9OQM+i2+FzyTnls
zbyNB8UZvD2ubZWo5mcS62CfmoQtgRR0q9cd5F/YiTTohEpIlcb+OYrQh65xmcsEdjAB4LFKsghP
BEF6GsLHUsZS8olxsVdeJm7BY9hxwL25H0kZQoLdqZulbBym22joWMen/k76cIWAleyZ3fTGeEm/
+nvT3aWXRxB5GCrsp4X0UC3khUTD8TUW1HE2LTxab6cQI3+LkiXtrmgxGZAHOz/kHrUT+5tYDW/S
jLGWJBx75t+pv0cDiSRDlGx87S50lCsgo1o00KWTCmbry8pdnImHZrwmw/5yhuGuqmWM1NGH7pZb
fkCTQKTTiB0W++AzaE6sNwV1e3DDoCNHPjJnmW8AVX3X7PFI1MgjugYN1cFIrniYhpG2FEcUcuP1
hFCayMy3SMBu3ICVFzMDOGz8j0OIVU+LW9YI2SrCyWyuDscDdxyc7ATldlxGsu+rzLNSrBlah7WO
TCHgN04MpWJjjsYHSrTUyKc3wfBv8qHlF9jPym9LEREgQd4eK7TdA7lCqmEWtJF79xNZvn+HRF6N
rqLpVV2hD7zYSqodOHe4vZpjsfGQgBfvSA6qMZ8OHRgjKEmzxKXSUGKI7PvPL57qUaGNQW04ztXW
yzV7wrlDvTfH9jmW8Y8F1Fyz7HD96dxhxrTf9XC2rAFf421Ao3cLsTlWFn7ejFRx1iywD4BWHbhT
U3vCTlmGuF934aoBgBS/0Oukc2O6jdv9YbFecXOlDKCDPXZxpyjiEptHm+KhQGxxARy8QC+/aZyx
tJP/B8NAyc0gGr+Ilh+Ev4Li+TGiUGmSD3+TBVyR2a8CfaZsWqzqH828bfDLpnR/34I4SV2FDOqZ
wwcp+PgDMVtM6OfI2omQmUzS2zZqJykL5pJ6CMsUB35eNyaFer6VXiPrvla6+uH3o7YiH0JSUmnU
L/zZgdmsvm/Ec5ZN1EMq4ukTtgxlsodCYPXLsR7K+3qktqbYK5Ue7lhY1t5G6m1KayK1D57RVeut
6lYDz8pqJ6r2FjBSS5OAPMSAg7ZUSmvvruMp3OEl9k03iXNQI4fQ7wMvCXnwlBlEwdU6BLNNWel4
cqxE3kK6xz6gIHRJUp4bjrHwviWuZkqkuCVLLxJCGPve0kXjUY5xibbRU7BMDu4shcZALD38PFA8
Q3JcdAcF43HJjZdk9m1xSK5XEXTgWi5n4+XOe87solsuD8le3v1zpy922B50tPgvO9ckmm4ezevZ
rkCjfqv1fDBMcotmqu+Gs2IT9hGzXSMOlZ8oknWulZoL9rYkJXLG/zB2XKP3q8NDAB2FVQ9DKMnu
zqWczDinykgJEsRtN9mYIFaa8L/1cdO/Ei1JJA1mmDmO2NKozwPJ1d2hdn96RYfWQF77h1noDmPZ
/4dQj+hoicwOQm8CR5bQYv7bo2OI5jurEfigQyKVY8GCDmXLwyJ64qnyorgxFVnZeIsRjqK0SAsl
gOXgT7Jra5kFcA8qwtvGD2Q21P2VdYF22PdI2UKK9rjHxhe6MvRGtZuwBK9y3QX/rBsJCizT0+Df
Sfr/TWAis9w57xc7IaVB6wRfuaG3a0PLREbLCE1ADrHSG8DAInXOfqSdK+ZcGtgfH4DcShCzES7x
4X3ErMIEWVJGIeH+8RGUglVWPo1v5ih8vRPFY6i7NQsCIoVomKeHjLdZIfGIuSwsIUKQpbBpbZVD
RtMKuz87+58lBBwIuKbkjnXjRSudWY7lvnnXz7WPKkfewUHfYBSlWdLTN98IGCNSV7tc4taQ6Gj4
BBcqslQFAM+9SwySWA5et50YU7Itp9tE9yiPQZGFT05ZYL+8jnF/Kph4eQph1HcCQ0t6xQhkuHKX
IZHc1RCh8hEcx80jmRdNyO/QJpdHI/0FmU0Ne4GUSl2ralw+buKgIWDBqs9OBxdjuvkzovqQsuiH
VCDulbz17VkkY7mr4n+MvhVRT0Ud3RiKV971W8PMxO0L6/p8Ni2dWNeyZ5XWWC3DAB+MaJSp/wky
Y+r3LzWa2duSoVPLvsfcx21O7/dDTO8csjcqm+tJv6B9qfOvGjNC79DHWsxHCMhOqmUKamhGlt7D
KsXCFfdKiYp8c56s4J1RF6GetQrSmB9O7lgRuB+t7cUWi8zGJBzWTGyYzwJn5dlzut9Sgtaamdel
pz6hzHjAclhlxXdC1M/x8R3/yLzU/BRILNJXgpKoNKhs4h2r14oCQTiEExKO6tqQ6joCNXXXYfMv
03mRJKAsJEMOmTMUMpzSZCRnLjAmlb+m9o9I2SPtLhOp3JoneQBJSTXhynAf3TzIzcLI9VIRtbU7
dUU4A8FDjOZcBwcoiCXhrtgzD3uO7mMdeuSLNHtdhC+TnI78dT2atJMCnHWEZ7EGRfRM1JXxnB5W
apivhJDRd3tbz7dOb6qinpbo6N/Hqi/SX3nGBVaJTel26Ha/D1hJpT1k21vuZBaUYdmBYQ7xF6UW
/MZmcVe0CZF7S9CiZzUq3fNpHEQXEeNNCz7CxoHP9vVcCDwGJdKI0y+EZvTuqYsMUjslNzhsOXL9
FOm/CXx/quqfrBuRl3SuvTU3BanYmzua0j/wITYygh/JtfP6CYtrw6Y7SgWJlFoq5sX3Y/YTrjIP
FEUhdUwqrSG4GqTKj1H1MPyJ7NkgIvesPvxc3aRhwwyRK68c0EDcN7m71DAxw4avPmocreojCP92
bc3QOBVe7/ncGc3dNTYqZAinx8zfD20lykz9c64ysJ3QB4aREn+g2+lQeVagrO5UCx2KTvkq7fv9
5VTn/ZvANPemb13LBucDQBouSP6G8bDExoFOJ83K9DuDYVEoA9fZZbJaVBTKfCTDZI2TRIYhtq1h
Ja/VTJVwh1vLbB/91mW71p9+a50DPFuz8glLYUrZ3tIeQRLggwDV1ZPnmD3bvVhYj9T/uwm9M2iq
YZADgnaySYkyQnf/pZsyjmCiF8EB4Mv9z4zsT1mllnAcH0Gj5PUFDgMsvmt6f2hqj0lqMjhg4sm0
un5C30iwzrqE0zqXlK8y+/KMkUmDc3sclDu5loAWl0x+H0hcuz+NmWPQanGyk0bPaRIur21QAVR5
orRLuxucbtBfPqGtN55VSg0RWpSpa3pBKilj5KjLNA72v8EUuDSDX9yytuozXyy6EZ92Ju2tqefY
0Nv3pGAAOq+mg4GVzI37GVaZ6++3p9JX8uCEjyaXLUpmf50TJx8b/msmgPmOHqLIkgeK9QyyB5km
KaKD4lcXw23Hhd4hnrsSKsFGXl4L+gUaFxUQ+Igd7uKR8+2PBE3zh3L5q4Oa303GdfkBf+l6sJE7
6P//HlwkBr1pzNyO8APjyt6EcfbK7maIhXUlU0EphO+dQpQw3ECeHpRLoL77MdAqc6S7Al65+qrh
dKgqNY9dzhHaAZ4eKTDcZQsKh9ObBbGvmT2zGqGhk6iBvR8xqK/1amvGTY3fTs1AmcdniecAilHX
Bsny8S6GOL5jhdfGbYLBS+qJlrI9clz7i+vdFIR2sg170SxLVCSNg/HhsNagTCwL4H6nRdIlWyj5
EHxfe87ndFWOP63uC4Wol7JFOMRUDNr1BgFy/m/1fpX977X6U8340CWvG/aQlpNw90/ublDlAowo
Fr0dIlKejJKpjS4Y1OuuEBcCUOHJW8xABSEMt+PxGgxjIUIkoAy1504Hz3rXY7erM7f7R8/QENgK
2Lgg4eD/3xI5lQIw/vIxsAgY7sjb6bC3OxqHm0Fb6DedOJL2RJuHRNRyy0hjDYg6UT3KMnBL7M/z
ACsc/yPOHX7IeMIen54Gc5rPLlU6hj6gnxfeKJwSsMjO2Hquk+uuKeiUxWXttvpQMkI2AQgI3C4l
9ErtK16XkbdA+/zcJE0wl/4c+0Q9CReaMjXk4iBMhBmQr9czUIQ3VgLSrxNJyI5QJApAXiggZtHK
3gHApb5/2UKzqvqy0wX82fd4aiSUrhIjuhCu6ZOGwl2yX4BsTDS2gg8RDZUhTeUtbucptNxGhZTl
UNZq+IDa+x0Kxn9be+fnxX0DAiLsVpVROCRoknN9E94jTBNen3oet2Alhu2pfqhBPp3A08LpFT/+
4QbfWrFDTAWOXpIRycXu2yL3jbBltgvHkZtsdKbJxq0KloC0UIzrIrQIswm14iWrqdo3VS6i9EVH
+iqSiQAgd3KKVjj21nQFq61hblJVSj0wstxPl+TatmCCk0TiH/+uk24tDnHGiR0s0ZUADsp9WhKg
O16KjosS7VpCpv0apJqtC56oRm7kjDOJZK7evmoNVzEFyO3318WUd18gCsoGTHWLSCgTR2iPzxjN
lHLa/A7d9BTQxLcfULo4Tbz+xjRJxY3DV762ksWlRZVT83QSeTEgBY30IxF3mlUJxDaYcD+W7twp
dfttSP4wQ1wdASWYM5cvjeI6063w+7vGg5I7UEH0YzCpvf8pBdLgGjN08Q3wSfFD7C9TlOsPUBtp
yAVYvJPiN/QDc5LGvLxCnb8azKyBKj4BbY7TOVDewUxHuXRp+EbO7VvJIY9lBxD+zwuvvKOv33fj
9E2ou7fTXeJBmDNQeCqQoqB/g4T7qImgnR7Wmk3i8+p5+qz4q1egVooOk+FuOHByJ40cZhv1bTrt
Yb7K7KignSdxFCKq5no41BbX/BXjTfAUVfyso5BhdgdOcB6YlYEC/IJ6ZkkoER8qvR+4WXDS2VxV
mrzyk16BNDWc/Mc48enPCl3OaataprB++5GDI8NAOQ47j4ypBcyD9nIFvExfPC/fUWSS2EQo0oQZ
tEnqv9K3kJFMqYDFPtatmVwD/aUQv/eUnl7rZjrj3HoB6oO4c/oAhDDQk9zy4RwtDESa3K5js8Fy
D4B2+4LY1IsUY1wOAFz2X/C1FEAaFGYS6pf+mvSit6JqMEXY2NWudpkOtbuS+2qpLFpw5kkimxy8
+jQHfy83J8rNcjZWVxYp5euPT2ejlg2Y29i58EaCnHD3VBiYByqhuT+b9Cf37zo1WeZ0q6h9o5m+
5VGekPDSy3/rppRjaC8ItSRoDMuWBXxU9Qigx60EYEagEWGa/83UFgtm3g7SJRtoUaAUhk2TQygL
xC19cOO0+P8otxWbol9+k0lSBCwmspkvr2itRl2eBETAg2ZMkYPJZ/6nApBtV201/du+nzUegBNg
cOY2cWqoq3WtghtwMpxJ7JW4eplqQ2u6G6i3bXUT9uqAJxMgaIfu5eh/xK8hZfXI8r7vXHv65fqm
hXvyc5CT1R7zTZkf6clC3w9keGV/wv7FsfyhTgZjeFaXgJNctwagvN5Fz66hvM2OEvURgfWUoOWb
qP1jhSBI/7OO5BYHuJ8RCkKh8JdJy/j57jof+m6g/2SJsC2kAbeQ5jqbMAKzUK9rQ/IyGwM+G+0Y
xIkAsbSHkD/M7radlTannhjq51bElUzphNMMBbRKtUWclcfMlBuY0Ur+onqMtwBVsydy73OM7XLu
XUsG1k0k72v1BaCwsqdwL6G9eSpccwIGbNP6BjaXIosWgHh9JslkoKzY1QSwTLlh2E/1/6ustTp8
WmeJXOdsUS2r/qi6vus+X0qPSSgPaOFmgHuoZIY1F24zJVDPaP4qZAENNw46sZxSauY5KoDFPEPA
8VXPJK0UZOO0pXzE08bL6K/eh3KDNV1doPIP2MvRnq4zkEDEughMF7g/5nfP6eeGP6MkNf0p11L4
TZGieBWRS2ME8nsVqbTTDLktzad5DeKy3lrPEMjBuUf2yOjfTkBR7LsOZVn4OpYi1c0gBNFMcAvM
Zk8tD9+33iARmu9QZlwLtaP5KLP+0XIsIlddwfe7Fy5ZTBcc4JkpBNSJq271NWp/Mtl4f7vWD59d
dXcOa3lvS6UxEt3PytPzDA6QleX67pDkvB2u/veEajIIuPJcDdtUJt0he0GnTbxlNq5YhrB8ewk5
T78R8a0LgrNcHK+VMggN5o+57NbG6Kan2eZDIMSTgLn8lToPaYZaQhtnHWxi1LyXPUmgLhAQcn3m
G4stFfxHMqGaGEza2qscxrAXRj5QEefcuc4aJ5hhu8nR6yppzeQdQf7ryeTUG4gHHvhmz/P6/Uy6
azDBq6Cdl2emji/W2DCelRbVu7b2euRTK9iEb2fpYaK1VExf8Io5n36fkq6se1qI98JsQT09sx1H
rCpRfLpow9VNDy6+gN1SMGwJb6DwgpxPloW7W2AkNelTypcUW643ncL9GO+q0NfjvRNGxMQbzExY
WO91bCO0a7xDRvdfGzu6JhPe9xiU2MOgnT1J/NlanYWPkOGz8m8G+5WmKKQbL6fk4sMcI6JEQJqt
Q1iAijENkJAow5jE2KXlq30msTgHBEAyRJfeCCtm3c0GKZVB7GGd8AhsTbz5ED+gW3C6XpRcNLT2
xOW6Mb6pEuZ/zuMPVfRGNLVpEBIJrI/Ymj/Y+fWGpcO1GPwL46Q6gPcSRL8yjhpAN8qCvvKt19R6
EPACneZ0Lmwn2lt9vUf/K8V/7BLDEkXj16gF5DtdYpS1mCBDu8jY53RSHqx4sFvZQdgNDUlykmUP
wKkjn3HtfyoAjNmtHTKlnKpXe7fGFW5kp8LP72epfXO9nnIrlMltxskKHXifCiRPHUC3N0JZAoYx
GsziJ1iOgOCHafnPp/j5VwMnxhtISyN4AV0FCxTBTM1CFOVeprlVUdjFktWqZreORSOc/0O4l2Gu
0ve+KXlSEQ1mAipIoGlA5YntgA2vHShr9f2t4eLWKlCgjEhsA+jA+tZe2wupytMahBTYLvkxJL0p
UMjgmpd/H2ikOHO+JPZVjP1+v0C5M72bHhOtzt+0FFiY60ifRureRfVBD2WfUP9Y2SWkFuorS92p
QyvwLxFmjU8SMbm7cb79zWbby/mlDR7FyKeJ9Q3DdxFG7DRbAhC6fpIjlGXfHGTEkBm4tYcl3mAV
rUnPmh3NWp9HW8fOAo8MgMQ39Q9MpmaVJXoLkDokKd64qjnFkWTwGNt46/Q9yzqWHUhZqaHjGeXc
tnxJ2MkVeG+2miTyMz5wRn61cC6qMoig8EKZUb1dRfQaQIEINZXP0SbJ6lLtyH2SadEGKnGBxS7p
PokQsWNHeP9ruPbg5+DiS+tlFkmCNITTW23mt08f2uUYh/K0BsPk8lXXMCXFCWFOhjuPz3F+OhAL
yraMYIT1rjX3I9FthdP3jaNv09bljZoYxg8W0e6M5ncmnefc77HO8C2ezgHf19io/x+78rfkKBXE
Zy8f4XTV7vIjqwYZgA6HcFC+iA7o18s0OOL+eHHX8maUXmydV3kgpMB+b47sWxxIsDt/mXbjk1P7
ZKpVIf/H+0CFIiN+ySLrJOOCrUT+aMD857QY4JlP5AkjQkflIcY9mRlSfLOvFynzMLjl6VA737EE
WxnocOkJ1S0/OSLl8ktAIbvSkjqFxNCs4iXdhJIlNX7fG9O5gnoEag7MgFQ0Dee6G3bTwoB7CcM9
ZfZD2bodsNt+YkJWq8YxBJgMH8lyltMwdY9DU9NoooYhX9xPCz0F/+aBasdeP619FQQYehAMnzoa
EWkWKQGaKHdsiubTsmodoIz7chAi6joHDpmo7+60GY/h47Fdm5YbHyC30D3Ly9mI+8rBskVOzfgZ
pd1TqOiQjoiINWQd6nYeCN2hUsL5591ohX/sCkCNxWdl5J2Ri8QYdvcich2AsRSa3vN6shhT8r/2
zgqrqqsmQDXYS6WB5YoboVUtmWmJss6YxFoPXoWQYgJNCzpgzKcLFrVmVSdzwKbGv0S5XDYTDyU1
tcucGDJ///cmeVIC1Zo/EtuGpejuf4unMOECS6sfFqrrj9CAJJdsIm1jg/7KtkQsgEWUx41G/Khl
TtWQ2Mg0f9aXcsiGlaouZfzuvh0Z+UI9lgeCCNP/mgo+zfaJZ3v5BseVgefFXVjgvs8l9FG+UqOR
qdUW4C0OtIFXF1OQ/72bxkIejd01Nhd1flqtuyzX0bOi/8aSUplx14iKglZHB5/vM9fDHrKr9sGn
oUrlgJYc3PvmFuwNd2ElEP7biBrupWmp+6O30BPaDfxXk18/GK89kji1kRwO4GDzkOaI5lZXEaSr
1rB4m01zlp0H0STnDrq9CfMOrbioeNw9sVkxtmjoVQA+SLHMKzywSvyk9o48dUPt1BZIfi0s4YMh
Dvi2VYawiwSvCHmtf650xpWzKbMBeJBf5QhAr4rrB5mj4ZmdG0utN3KQMzEcqrIf3Iyi3nC4I5m3
BLUwkhfuWE4zRKiTgfHP2/eOEILsr/ifvfyqTJAIu7I4UJvNowvETPojkKAfOPIdPxU4HmLeLWs/
3OJO89kDl1vcJqUTcTa8PtSXjW+1diU1e0BPXXh91vW6SxIse81JWfUvS/m9nsyVpj0xG9BVRgMH
o8FdjhTqX1GIF8Ljn0oMeRGMsZYoGKtHMB1C+17rOhdXkBzMOxFHczC5z6UPvL+lPq+5oIWXzWKK
5Xn9D6vUmeilwHdEecjQ71sYIsrXBjQW0xjbZwGgQGyEiYxBiSycn41fsAeXCj5FWJhDfVLEt4c3
cr9a7GTydamf2ds1Y51CxUKrSpWj73/EYfhEcUHurqucWh91nabNqcLkGKXn/O1kyEX8gf97Y9R4
loTK4pWmld/Sb5/ZkKRHxTkm2r28e12YqKRucYavG+CGRI8VkEsWduwhF2Et1Uu9SfdwdoM9rNPb
OSSYnCIL+cz6LhgbdcrZVuItp3fcDPVAuvsib53Is/ne+Rfh+1b98101HsYFahZE8R+CrHVynEmt
IVT5amnAJhrplVjiPWPzFZEcvKC6hLh06l0ydUmgb4aohfi3qs/+l6VqSCrqEatIOv7ZR7YixT08
5Orzad2wH+2ktesRcpniGO1FssfYGlfnfaWS6QzDibX/iXS7KTGdR6TjrVkihr6pUDRjgTw30kiD
6Mq+9BGWBZn6VA43ogCpqz0U3G1FjM1qarQtFnxR2J/rauknVSze/rNu6fkIZWbv1zHUXyw4i4Wu
dHf2cVWQuBhDZVTyEA5OqfeCmCeSkZhUjsv1N/ZlEPxQDzqFdYmw8bcIAIFH4pe+beIF60t3dxyx
Zkv0PWhw3u/S2hxzKvFijoXExhmFuYjybR7GcOByD6Gy0SuszE8VreqCV6ecxOig4ezkkO8bWzoJ
XMXDQ9O2BY8sfpBEaE/+1bSOCUnc0CFKUHIa3k9UfI2JVTQn0NvdgOHJFJru4CIb9gdxrIlW8kU7
qIsqjAP5v8dtugJ/WCkNoyE5+Ah1GdkAwlhQ2J25ZStcPo8aWwlfIcWNe5Wf8saJ/3/oU5SNF54l
viDfyk9iyDU2SgvdR/7zy/PxR8aVYx5t83869Xk5GsczxJrCfdZD+DwzHW81SXXzoxyZ/T3ESz52
n8LjUfl0MYuqAU7jT4fr4EeukUzbvt18o7gFK2cZnMP8NqVoUroFsYIy2asVKKhOt1U6RtAenEr4
wFqKY0/OE47Y2WmWiPICzuGaa1MJF/9M8i0SuxPn7wCFJp6M5qrNGq7uOtWdA/XiTG/v+lVVx6Ul
yrrcwgdkxg3VFenZo75e1Xb0HAqA8LPTYgWq/wgwz1l6mqx7+1SEGJUYt7Qb2uPdNYlJFS3TFNFY
yVdhZhdFIdZxR9FV7nRJYLbPmCVuX7HfU4kIpK9FhZ9sOkpyFoyFxrLE/Yf5OAXei1FQRhsuC2yj
cEGCzA5MA2C4HJEY/dnUp3V+SbEoc2TiioTEl2CRXRuc3XWIhRGOcaA9sZY/+mUgmiNROPIOr7hJ
Who+FXzcqtIsIrmlPqdmtvSqtUGzzQIsXaop31KmP8Z6IIRjiAFGb45EfDR6J3isKSsgkTnzsLOv
W0Hbi5Rg2qWNrXNNaHMDwIlcUwINtH4M7KKoJaSYMhtDyJ0yN7bQVynS27p8yrGHW4sMx/vhwF11
nrXdc7nvNG9lWYFGsZH+BJr2mb99CdweZcxTZPZ9vVkuR/szw3dkSPZ/Kee+s08V5IeddXmtixIw
FfDEPYh5+E8DK9jz3aVXtmcC+N92i1/5kfXW/Jy+ozJDz6iaBEBT/vjuMSoKY3cCVQTuRhFUNJUV
Kj0TcyFGLwHE+7ZHaUvCL0LuJgjaOJsZqOSlwj9Herff0zXBB5oPHc6iSHB10op42Bl89KQeu3rh
KCULRnZY8IQfIm9TAAP4yB+ND+3EgEQn8O8EDs6oUPK32YQ8jJ1cOdQ7VcXN6ewU5IQE86/4hj42
cRX9TrFm1Td9qShI0tbwCwGfmXTEg/9EfDYTJvObJL84ITkFKKWreKCUFOW3lc0fJRWZUGwPh8E0
GDlFmiTz2C+7uxNRLVFMAI/lLYjDIl+UybzUuN2h48sR7faueveJJk+01020UKFTCQBGQR+lTeAE
6zvhkBBWJEqFFALrqD6iiQuYxWeqECwHjvPCff7X4nRE5IghJ395aOwHIvNC4QG8hADPEIb/Ugig
tBrkdxVc/9Snbqbflo0Gv+wGOAM4PH20gqFHtBEs6kWbpeVWYU352zzcfIScjm0ZHoPO4K3iu64o
V/x5fSWeaslKdVjxOQpPbidNew1kg6j63lKiWUTAYBDimJc+G82o3rb4n8AUnhlEx0vFDe7xBLsB
J+jb1Nkjbxl1pOpIqmMcC/DWv2FBWu/mJBJmTWkKbJqiTfKekEFSIiDcq3TUVL1Whl9/9JlfdGbZ
2jQ/uR0fYHkfNlV/z6Tavb32q0zzGcIE5ceJeMifLU2opxmOhbpOF+D772c3kYV7QGbIziCyWnjO
0+i6bTnisoxNTFXUBMKn79YivkX2dDxIfZPx+LKADwkRXQ06aHzYAR78G61gHH9u5fwZuxNOx8xG
9eGfZ7KaIWdNE1LlHSNXcQeWYxkcOK7c3QBczwSV4pyvijCiDoap6ig4TaIsd7v0Tj5fGXUV06Fv
jCGUBw81oXAAFGTxAqPVE42mqG+Z/mbOkn0KeJ7k2XNXocytRcNnXuJUWNaUU4bqGFBm0Zprud6N
wLYBqDj1FEwVUGjfLJtZNUZnu94g1eKp/YNrW7IedsS6qBS4Zp3OsQQcdRhCHD8XtJzWlrVtKDNJ
avTCsWIZZ7eVKpw7fROEIIo1Wvx/HPYgHMndAi7olbeD/ZtB7NDfdD4Ntd1l7gDk+Wn47IBVdV/N
McCHpq3R+V5ppkx7dMImIUH9QOYc6H7/6CXyZVW4rsHHpgG8Ug59oJXhYPQaHbgtWrEt3N/gnRUG
CmxRccJWt9kn1wGzklfhoiSjqd2wCEArFSYxG0yJmVaDKDwYmYJXQkfpYL0aUt+6XH5Zbc4EFHRB
LJISDG6BWMB71yHLmZb09mLLnzu0cl8oW0VgZa4byk+V+Y9lEOi7U/HSlWtqnG5LszR0VR/R1fxb
X/xIWYboOdpCs9nbFUuK1jJg0tN8LySP8f12LeGN7wwX4NOkEZgTaOhZaoYB00U5ES0Rj2KqAB4c
yuRHidbzgaItSxkXWnWZ77dSXgA+WGQk+moOKroBq52HixBOitLbE/THBcm07CXf+NYniKSgAnq+
1wdJzf6/sHztMtPIdhQBvoMRMrIY45yvsfsOWvoCtvIM7gbEuLRvjK1jZKfyB3mxF2YWRMwByJ97
Oeu7lrJvzNQkyBmahNtDZqA6WHhZe0072Ys31ElQrm376Sm+synyr8ryXghreQ/Sv6lQ9JKMvAC6
+lU2GlJNfIa8kIw/WnrWAhCM6mkVCUnKoTx+r2OdDP561wwrx8GZAHqTcVnmibgPjAkRPvBHKnKK
W+1VxsAJZvEwnWFwzN4zKjRV3a1ueI9L820kqAsP3biTBslRw5Fi5W6heo3D6zlwSZVZb4av0hXE
PUpBG1Yl38zoPDP//mLdP0f7zEFYiKmf96bBkMe7gknBRvvzLH2ZwNc7LiRD3UUMZhID57GhXd14
DkB6g0R1LnzrH9hVP/cEmn+PWBAgp8OCznr28UHAAXqvRQyojTYIyP8L4oUppm6jmcgTOfa8Xc2x
kJnicN6R3uYYdb6SXxhdfdOuj6oUGkqZL1kLyHC9mTt7jFqpif0zP6xvLza+NbWxACS7fZo49QKR
wtk4ZjX2ccMONdIglDKaYB5x+uc0j+/uul8VYzc8gBra0ke0p0ZzI9lWrmFlv2Wua4S4HWVz5rcv
CtmuDNECoLu+WUEWP8iweVEFmdifrjOKyPGhINO2TNWIPMpxPFK3ybaP7CE+McCDE37xvNzc4AQ8
zpWdojrL73i4gohOCsprrXKtzj65MdKYVg7jOtjYlecL9RVKqDYwJRp2W1ZoRgLwC0frZs/YT8fy
VLOah979ofzfDjjAJDNp2rHdyi3SYx+hIEkXN5dgLaxqC/5D0toCRL4NGQLMlIkrFJj0InCjlQf+
nhL4Li0Odru/bvmqvcAJl55f9nOSJtFywDdqLBmF3IBRYJvL7l4Z/sOzijdXF251UkuaUH+U9dTm
ikmrcqdcBUQbfLNwGkvNw2IRvu2rZJfnruCMwsMJfdxn0Kz42S/maNFe+TC3ESZdyO7DUgEOVpLF
B9ZYaOaei5d+atJ35Yei47vv2nEhLMPegwpG9VJyvl2/eggJ5GzTi24QrMmfcntodrPYfYyLpAEC
7wUJuPSC99Mw32fG1kYFyN4zfROYqqIUdaa8Tv8MCI62XNvcGP1nBriiuTaVinnilwtIrqcJQQKK
bOKHJJelj+tPw8f/qhCZoDCiEueou0I1S2Q37JO5zlKaow7Z/KzCxMvZhcr+7zFILrEGxq3j42DT
TtMwODzgMGJfj9lEyiQ/E1NgnuPsN6bjTcbKDoF4Ms66xDhCQP3tjJGUR7+Nggw8FuLMd/Ui2WBb
WmyfHMiz7p9vBLw1Ub7kWDbVVAx/6mnRg7Fl3KgZ2LdW4b5GJW17fWX6aZIQX0TFzl24t4XzR4Am
du33G3y/5CJjZw2tHezHiAf7n1bzzgCurCV8t5XSMams4jA3y6Oit+QOTTO6BE7EWYZlwZpTWYY1
ecw79dkztBSWpBp2bouSkuc98CLpOGgxz6SHxKKcaeDT+/t/oZvYHtZxxvNHEF50/rAqBa/SJing
XpF8mSdMbXrK6dcuwM6/8yIhbNEUBx/8BvXFPUKHmPio4gMzSBtQnUFEQ0P/UHIDdmvyEHlpJenM
L9+xt+l3OMN3PTMWblqsFPJk1bOzpvyeZaW5uNX9pUpvLo0OR5B1EnpjpqVCwozWzX4Xs1i0N3Hf
RGi0BUBAb+n2h7Jg+vQSKBnHx4EiuXdZXHDf2xCxlD4fAiaOfF3J5QbGciKLqG9Nzsr/dTgLtDPQ
o21Nzr6DtUsw/Ps9xMcv38K4mD7a5aEsH+CzxOvVTUNYPpSwWY24Uoh5Uk5Vd5rAjhPOWbaFYfRB
fLpcncUtzkbZlrgKSDopsmmbxioR/lry5gfxbFb+Lzvj/DcN2DwQDUA/77EVVYXs1sRLjcLNUoXQ
q5nfZNaQvPq/ECnJEOcU9pLxz5uCFnhJpYPbfZzEz2h34aNGA9NVwBlY5bCTvT8HIAxtIC5goqRQ
dWAdEYqVKe6X+YUoKF8AfXzfKZcwPrWXOSpDMw2CYGr4Hl/HF5vwrFR0/6wMua5wu0jncmzVUFmu
eMU2ViszTLRCF4Lx2tUjj/+Svx3I6T6SP/p4EyqcTeCvFJ7INoJyK1dftQMfKtngoqpbQlw//0ad
jwOvqIjFWQx5DOe21G3FoP8CHcKtkAUsirU0+Rb8eVnKXs1rAsypT/FbdoLsbFzZaHMdKhjOfDCd
fucmo3cmx029AOOtSKNOnTe8/AbZbkE7SsyTF9n4K9yk31a88OV3ex7axa0Dmtj0lEdS1xq4sw0V
EutbVGY2rXKq0MKLCKkXvDXtxpxeQqr4YayOAc18CRvfjKS7XIiW7QVnMozOecahIafIHDNU56Pi
nhIXFTXJOt4Ujq8snIjhltfZ3PrSGyS7xnBXRGKTI8V2XKWp7Xx50GQY84qiq5cWQEK4pNX+296P
vF/ulsI3JHKNUiBwu53V0Bhxora6lUqqAM3uezDZvkQrDwIr1qUk3XMO1TiJcIC813xH8upk3vG8
TAdC74zxstMjiH5M6MYc8jd5YbUuWjfciYg7nGU/t33H0YAEld6TDgz7jFU8naWH8B/NgpV8vc5F
+kTO0svS0R4a8/6l0K8HAySKtcGr9KFxncRnHo3EYmyWqoegK4g8JIr4RtEaSJhmr0UmojDQY462
5XmQjwr8OHzzalhrY7GAjLxgLWtFLOm5F43uJhY1i09YtCpdcfbbuuGinEo8sEzsfpYtH9pKmGNS
3D4NTNAJjuBZ6GL2E+qgQD0gKIpCeh752JO9e8XBbgk/LCrimX5iEznKoxil8KVHDFXvBYBB5M5O
0eiVjaJMZqV/dHZPXuoqMwFK75c0zGfheoIS2s2NeRY9BssSMYoZhDGLmnmv043eRD2cP9ISdj4f
mKq7GwNNJj62tyl87n5EMHT2I2pX1c0x5l+OOUry6llEfWsich/3Q4Z1PiDUD2fTmbP4DeGB2cki
euaVVgnpRY6dwL6+AK0vlTmZnZAm3s/pw15u2nb+gh1q0GbUaqSShzLjUsNqK87UW4peB3yDtXlz
tqofHmB6fVfHwEXmtEln85iLH0Mj7iRoFikZdOLVZIIam4pCcvmaL7BJ/QSFYm21ULoYduzXw0Yc
NDersLf9EDQD67UAA+DJul1ccXknHG07YRg0x9s5WGM9ZLu1o0HANqn+aFKnS3KDTCQrLeZixZfn
KLN0Z19KKwvmAof5OHVxCuIA3QQvdJsKZL3dNYTUdT704evqKcj/7Tpw7cF4nTUI2ZcJKLNfEtzL
P01CvSRXCLvgB3M6Scwxcx8HCU57N1vaqwCfywXbPSb+l/0nm/o/av8B+tn4N/DBKlxPJgRFIYjE
7n6WDEk1oMn/ZqR1uVYT4RYh8WXxylzHn1EM3sZoHAWTj9bvkqv3j1xxG0UhyVXIhpXKtkDqXc+d
3WSc2XisiLmdwS41rOpcIxJVDyrJgLeIA+ByaPZGIjQTB0hk30Zm8im9guPrUXrC/MQ69xoBC85d
jQs3aHWxl0Ss1a36vRhfceKgQd8jgjBUFISHGmjX8NYPcZ4XptzmQRp1ncpEyMQ++sth0g/f3ugn
qF2jipJLQRadpDFq+EIQxd66zhXWnUtI1kkwguoBik7PJZpg9uy2qGBspwFoiooS2LxSJTQWsDHr
BFedtOhB37RmY2xD1nvEMAq1mPviyBmstfsQLXcIrt0Ty32ZSE4wUP+Q0Wpd2ODHrqV9GS9Aggel
Z3gNiK3ASmyuIw8twKW1dV5RpuSOoKWL8IKxeEIV+W6gJFhSd0TcKIWi5nKRPyFTpI9o8Hrvw9zE
+k6nBav8qzCnHGvOxeiikMedsVqVqPkZ8I5kavwELDNAU5dJuO4utPid9Y1WQHHzh6PrBKa+nwib
rglaGYWsx/il/ivSjRMMJ1b8zEQlc4pQIRMh176xnayyl7bF+fxOun0ddgOzEHnF2KYHHFS/ONle
5XegE++WcW4Ybhjpp2HmcKD8e9cuS5MJn0CIaNOhsfkWcU+zIfwHx0HSErjcR/jV1XtcBHlWsWP9
ft2e09XTQd0Y/l2HTCjMl1fuBnRRVDyOTUAcX+NPEl3Td8EFhpZ+vzvo7H1oUArxDRJByrADOkvl
5O7ZqsCRQAhLQQqQ0ohKOLsGzMVtLMEYsPUucDDnBIZfTXWVfYrYr3sM9oerr7Wt/Sumk8AmznHS
6F+HcfRbHQO+wtBwBVbKMJMSixgqKjS6kEqC8u4l+gz6Ciih4pKfUdpz5z6kOurznCRhC604Ns00
bTDorUWZicZRSv6Y3Hee2gkm3MRuhU4pSKrsrm0CNeXII3L0k/HVjfDe3cnQCS+e6xaZka2pAkp+
sFlj+m/lJdl5v8m0d7MFg1dODMPXTT1cQ7mMKnI7PAAJ2I4Dpx3ZhDCIt+51FNY8YuNExiACLdXl
DdoaCWBRGZAzqpe5CHPcce5CP7dsX/XVuaLzB9wB4h1riQw0eIJ6+fsd1kA4mz7Ezsq1WWDR41Sx
gBXXZYzsgZYRk4OUz1xopqGHFCBMCbpzj2DCxdO6G8waNByS2AuwatV+bTkZ1ttN4k5+ne7APZbi
P3OfWCnHrn7yRD60OWtBrZXE8CLFixC7SYoiqZ+2qdVn6ywPFyphxQxu5lss4KTfx1ZFWsNaDFg5
caW2+bh0TwMwJ9NJe/X2uUlzRxuuMWig2IOe3mBoaWmUzQMiocWhMcS4k/zzge9qcAaKh+6ZY1EH
jQWUnXOYuNlLXADE5090HjASRRUG9+Yj/k3AhiKEpHYurnk1jw6oGQ3geaQSbOKDJrGiX4a3iGe8
ambrtZ0ivo4J6yhnrLbmvr8mkkTTn+fIG9hZ9j11sq9DdV4wjHFVMvS+mB1g31/3DUrH0w65UV6V
hfK6QGBHjEIxalFyA81wxppybTyE2XIUdU7Ue9yWkX4uUT+BmfshRXmiqAAdyLJTdy18rDkTp/U3
lX/3VQ2rCf7aV1eLnNX3fIxqdKVzka/aDR99n0tVppFzWc+I/Pft9nN9i1IHcOOKNjEwiQNqBYcF
Y+cjSGtrhNpykSYMgTx2mwgmStXhyQ3keDoHdBWQvSkm2HPxgtFmF4S6nTkNSZqYmlm+UQEFB7zf
cTmzBD7daj8HXvskV+9kzPLO3dPR1uQPMqUqmsYkpn3PvHpxb0mi/W51ukUwONxgOF5XXcian6e3
/2IJm7Ycqqv8G2Z1oEy+S4eiEmMl48FASMvP4UVG6xoVEfVLzOUrLpa7u/Hpapd/ZMssi5EOZ96q
VPjq7FrC1AlWYcRhd30XDCDAPrcFItJ0kx+goXjP7tGiaHuXVS/+vz32pZHC+QMlL7vSwBhEgXqz
IMna4fe67KEEHRqELln3svZCaukUWUXjjrGw3Cu1fQLK18NCQICHABBqxwCFiKmU7OCG8C+APodm
fzj0gpBLhM3rdIacf5kksKPcJGwBxmo33O2fs3UuOQBXyOageQ60MRAEs92zVwRaee2z4qjjj3Rd
6XJtOTuze2eIjIEZIftutpbUbOTXZ8eEekyqoWaJZuUKDu3kcimvIzD7ueItZmzvg0c91rVrxrXl
5cak05EodaBq5DqYrCONK9OwxXEzDD9OxlndwAuBnOsWE9aYDkCbxm7gtshLIOjFaH1LWfMoGc3X
2iwEYqOBIpTO7RGIrIFUCWE9OzMnmOzkMCbd7L+7ck/OYVpzOQFhrlUQyxZytfHSCgCLogAEKlvD
yTq/n9Qslx8sx6K84Wt9epKTEyDeQlYWijbR/vSOwC5AGh4U5f7HnARrLkinkq+Zal8gw7T8vJro
NN3YtqoCaz8pZyQFx9N5uKJYpkU/bSJVmf4wS4J1z9yQZ1RYjnlLt/PLTlKoLQT7IZxEn7syBKWs
Eo41EUv67jPJ1X+TiIztjclkNCrbD3CJB/vJA2PZ72BuHfsYYgJTMaaR/cRtUmNvIUBR9yNuGBau
5R+aowiB097ioJgMQX2d54vSNK5FEEB+c1PGA7+l28/ovCq89okNIp0FtbTCwhhP4Ve8BZD+3t7p
01Og299KdmAbIvdz/rLlUs4TJ43YWZFphm0Q6e3XsjX/Rnp5LSIR+96hdBOeEwip5BqU/G03wT1z
5VHp/pVkYRq5pX6s1BshKZStzgU/gDXR+UQedKiH+Bpg1Te8fY3GSFVMwxSMLU10QHfu47qnP7tK
132AJpMB6EiEnvTJ+DVAFEcpKuCI8YV1n6YTFViuATOHpzLR7gwjxhRKu+5FzoPvILITZfruOGkc
75C0KbOmJ8sFtsVMJjfYKbNxSrvWvvF4qfIvjkOMbc6kZPBZo1VTYzo37VmzqIWlzNc8XfuYASpc
LT5DthlEeXYd2xqkyurFvHxHN+TcEDI4WE1CILt3WyarUjc+plSdJoKZW3aWkHrRQq6Q81Lg5jhc
yJnfhc2xVriqXnBQdb1AUCr2xzfg82F0gYjfJZNldfN4IH3RimLUKpjxs2eRf62kU7/EQVwIoudm
MEaHa8bhqQ/8Oxi8Vk30BGc6l6TwdqNUbg6eJeWPRyUA/uJso1o/4Q9Ot5kbw5HSaxi3LR9VLbJ7
QUgR6H41Wt5xQVhQjbDxymJMPQ9Ahv+h0ONFQTQM+pLYQ0EfTuMdpJ/zrVtu94Je7szT0ZEXUZUb
t4apidByzbsGelIF51Z8Of0etBQROjXVDD2ynk6Tsl2fHy69tRE9KNGqGJXJ69GTD6ih97OdbWoo
vJ3ToFujK/U4RFaebKhlcepplw3TjHwOpQ3tJu8BOlagabavinQBa6V0eBPGACTJb3WOu1MOIgRa
8H3nsADo8It5nZhW0zMrnnK/MqYVDO6CZsfZ71OcVWYEJE8TkqozC5JSIPArVgYHgT7Knwfao9sJ
ObKUC9HWVysOyrt+OS+LyL8dDbPUqU2xuKeWG15DuPEijWR5AhbbH11j3iZ+koP08TluLBVBb+ds
pAQ9zcQX1M20EcH11xLLYH2vPBQJStedIKfefaXNt8RVg6YfShGNYh+g5+JFFHAmRbd92qMtMtxR
dqaZx7Vn+mwAp2dRlAkIi5JUOYrbYCqiiKQowiJTsgiMElqnO0ohb+cxB+6IpFyPpcq5AV+2TX2V
ra6Q+Z3IL52fldKrD9greNKzmJ5LpSBAyhyMkbE6rF+3x2PuN/LraMm9gpKiyqyAwktvYl29qx4N
y3YBQYj5GeYC/nqyRKP3czUgzxcS0VHJQNESi8J0saimpMNVWlH8IOaRgpI+Jd2wnfkzw/mfnO29
nYhep2Nfs9t2OKiwTkAHclnOD9DfT6tTRuwgDTnbqU1gCcdu6YG/EogJmpW1qp/4FIx4cu1ShkzP
+MQ9APGZEeTAcHKcdNqhbI8oT//lX0/VWuPhyuCsYbqvgYN6IedTio1G2DFHeZWyvdfxc8KiZwnn
8I5AcBPB70GpsaV4x29cqUM3mRZK4oupdz5FDlnFGBTmzaJks7qTK5e69hlBe7cIW42Lt6Vp/rbV
lcxwjE1ijqXLjqN7sqOgi9fQ2fMDLM/YCYQxjqVm06027jKSUCaP81A5aXdoTO7ySMqorNrj2eSa
VOQKFMOpRumt4HipeCClM9o9nISXjFZL8ODr0JwhfCpudy/MN+z0FYxMvWC9a9TkPiL+01QABL8q
rx2Tk1uVVgPKfZm+G0KrGii/ks+DeSoPB6Q+FY8NIpY6qnrBq7ACYFY84eSHFn/MN8dTx8Sw63ta
k1QQTGyYXMCvPd+mLxifeEOoTutBhGbC25vELfba4OQQpHzq2Nx9VkvWy37b9sw/KwK5Vz2Vj7Ev
1VuKtgxg4l929RWiRxJx/tc4DNa6OhY5Xn4aX/EfqYNI9lk6b1ZDagFM+roGhQhnal8cEyTRX5ww
1wVQYvKlifNQ63dqOi3qnIZvRsMDfryw2n5TbA4Ysjjt4Ve4IwM212ZvS5gP70FBWf35y5mAfyOp
Sna/f7MozEahL6q+vupGcoRNPs/Lpki7vymc5l1c/Z8tKJHCJaEeAj7SWfEh1z2rRFutZgUy/Z+L
0tjZTTkmbqYtSktFIpwLosDSsQ2Iw6eIPlnj4knrYNMneDV0ldNJ0oXKHgKk2HckSAF2iVa4PiGY
7KzDXPnZ162sSL+yjtjvxZ3uAMDwjAfmfqMDDR95Ri0zuf0z529/MW1Nb69H/pkcr/UhEyfi5I5H
EXMo1OeC3n4gDNAqHxGtapHCUN/5zMKZiw9HXI2R144yA6qXpDP+sflWkDyJdeeD+9CifPl+Uei5
0UW3sR943zmuUHhi51reFx8XbGI3pyKDrHQPlsvwDSwSwK0HimnogHn89yx1UjTBTH/mJ35bGANY
sPxdsbrpPK38Cv0vMP0yDpzkseU9+SRsBwmfK9kC3vDh1E7YcC9DEdVigDPz6Ku1q88j1bpM9w6K
SD4g4tyRzUW4iIrR1I5udt8TWAM2Y9thlXVPDN98A3cj+ccv9I+5fNRIN358YQ1mWBJ55kCEzTAX
jNEMILx0ClhOCDCAtSBS7onQItTEX/9ZQqTrxNFKhH2UdH3qK7bfkkluActU6gpssAZA/rQgYyns
U5j8AyNl5sCdgXf3PK3a+4K4PocnAYkaNMZTiNfIAFed3KAJo2RSgONc0jFdfVAYvKBy8RXowqwt
/aJ5Kfx7cXc2K5Jce8k46tGLyctZxmRggwvQstU1ARf38oMQgJAFQtAQoca9CLz+lhtcS6er8+mN
f4Q0kqJlU7hPyUIefescpbeDM9JCnK4HthweC6+eJ2g8QjdFvQIVBhepLTaey+Q4guuYdVCc+V0d
YlbsjFRR8f5VRziimDzHHtUj/lR1fjcqXAzjQr/plfGjRMcpXMwy9iArxBflLH51MUeWl2p6r4l8
cmtpSaN3qKxdxjsJHWpT96cYR8NEmU1MhdfX2p8Lka9VIXQOvvTi3GwshxGgD/Ez/RN21BMN0UYp
hrPYsze6mywpbKGhoZrCKkBHdMDJa/TiV4Gll0ZVFZNwPXILXBbzk6DLRG+04vM73McG11jnd/AV
DXx5QTMkRBjgx1kKp3GpBuGwoEAJPaPws6PyKmopowtOYYTCOzhxx95NpI8mUKbV+PdgXCOWmbqi
YC1mSL1KJWplh2gUAGO+H3gscq7Mjmsf0M08HYwXt+T0+dhspJasVV+fIZZrYhCYbVuCP5tyJVWV
kdTLIGffHwFio57v2pdha3dp+KDGk+oqMDkILIqASpAjpw6cA2HaRaO9lQGHTwgOh79mfLASfySc
7Y9MnvHMsqP7bdg+taXWNwWgmeVOaiE0KpGuh4PvTWgZBOyqD8j/yEH+OA+91QnyK8XhTmnJ5wpS
AublRcaw8nwqU62Bakpds04Kx3PjqNHnTNWQ5MQSXJgDAdLAobHHlro7hc22yWke1bA4/WCOa7o1
5oJgZntatFW+YsiUvgh/pOLsYwpv7jrj+xAmez8TuryZLrp2cfYmk7pxL9bIRVo3RfOx8+syacMV
EHRnShE0kZXmvY+imfa+rHkcwSQeGL65MzHsZKsLEfK/fpw+y3FHJl1Fhk5e+hsajikXPse0nYI0
YmK0Yj1k/jxcwJPuoC9PhKZ9UcTfsDicBRAgtn2Ae22XVMCJ7WyJDnPuyqmx1EaZkeAO8oMYHOVc
c4lz6uKFj9d9d4onSJSRztqWPX/Ypcejy8qbdfoI98kvPTVPZ2as0kMf558eOGrYAhtOU2E+oi4h
jeuakD7lF4tSoHIaHm5MFXEg9BXmQcXQvudO2uT86JWemdV1mxWEViJPBHwbmUYiZ+dzKoDBQR+n
/bVKoaymnvBwhXT4eXtu+aJxRhD6j9sAq7cQJvh4w7iuLy4wwnkIiJdZTsah4K2zRb4mgqR4UH0Y
rcAslGqJeAGEG6yXfyVoClacK1fFhPKFogV4/QF/yCg+JiqJRYB4M3jNePDSY+/N5YHhgxdIUeSX
AEXx763mr4bMQwylp47ikyR4zovD4u5J/36f+YvfmMyD/MA/64562RXnN51DpDiQhSLcTw2smn1s
tJ25uZeTsrH76qzE9GcO/+jz7oturjF/1cAeQP3jXJrnr19T+T4C3uzfWTTrXNi5bPnZ+HdvttWn
9Skxj4ZF9t/NjCOh+Pi+YlVGfioi0ji/m4PNZoB7AbjkBOTz0KkcPI1xnsGJiVZiC5pKqT4sZTgn
UlaDK2Gobrlbvwr8nEfLBSTEF3unfJm6H1JUdxVlkoDQdB9XH7uuN2/4AFL5ZA+TbHRBO6KAZIs7
CJ34X9BEnLCnuNGYembDHJuVZueMiCVHzCGtTU+6oBgOOtPEYF+Um1dTk0wm63rVW5SPE470oWWu
fSbUggjFX5ZCtlvUGwpZJe+yqgsXSkAzapv/3VW0IyWW7GK6r0ISZqw2gxq5tVth1Y3mPMwjxgXW
zpqMGLxWcWRmliCizfVhsoeyq60KfYWLgqmxX7S7KDLu1Gair1YYm8SZnFBHuTUyooZLNOsBbRI+
jA7tS5XA248t+vkw7vIzVdShBrDnBe/RWJIk+AjLJY2BaUhiDzI3jqzfoFrAGLo5UPtY9ziTFZg+
OL2Tel9LcV/YiUoK773VUhnPEpjbYkUGUL9dZCF8EFhcF9o8ezT7ztLX7YwhbHoSR/2InKrMfida
HHdFB9C16eFWiV0ZrwR36ijbY9UlGRfPA4ASuDvR6Jk8L4ZlfF/zKRUfTpxiP8a/HsTTt3S+Bj7b
P9mcvelXgPABvdNeY6W7BAqUdbZdcqV3h5uEKRmP7v6PHUvB+OhevpOb2OCfDqlYxPDT7hjC5tjC
vaj8trcYVqUQmdquFGgb2BiTRmnzZeBwwP/eQ5d2PnWkGxcrPP+H2+Mo0SGsE1vcz2uvplxHJDWT
1QJGp7/tjF+srG9oU6PxoSjMvWOxuXFPP6NZlk1ysOmO7TL5Ac3Vx0mRmgp7id4JSIryZ74WdHF6
leUtHGT9sLxiKdBCCWf/01V5Hr1lVcPzOCw3I+DfrhN7Hir0az2FM8RP26DqtHMtOJdeFUsBVPgd
9VPNvnatKhyDcE74msK3KZDfbjhhvDca2Upeb1oB9Hf997OBdRd/KtVA57i5gYLME2LdhCl91fyW
VI3url+acyrhVw8LMY00cTY5bOlmZ0OcZRnnMaS3rft9zAVaun6IFvxsioOFLqdSMd+RTkzgvvRM
XC1fkeu6sJILOGplgmvgxIERTY9q4Shi0MZ2IJ9mKMcC1uW2LIo1aoMxkpOlxGdHWuMHAWOJ2sma
U7KCi/pCfCzjKGovnzCugsyqukj/OTjwGlHLhdYJJpOJwR+0kz5N371+i3ylmkezNb1pmbO0foI3
Ypcba4C82NRGIogVQl+C0NJ93rMlAtbO4CbIex9o2pQNZV51qjtIdGaPdeC0zFNhbWCdarfxTIJJ
PIkpkYexNOGca1GbyWfozDwn+fQ/bttbBVpMlpWiJCL5PIg+v4lch7rINthvujyYAQKpbXPIFJR+
oHqAVjCz8DrEsmazILR5QHt8fMxlcjWUcwN1KhztVEI5M+F1EHdq961Us6EDbySU7uRr7ogwsX8U
V60aoMhjb0CQc1XQA5iqkhYrNNMROPG9SST18zVnslkws/4f3uTEaV1hrwejY2RgRKKr63O8DW1K
61E1LWX+cg3Ay+6W+VbTy3eZyZBe31+nJeengm4oQa1/Gfiud8QBcvO+CEb/sbMCIPYXE8IbZcvj
41U8WjT+pUDy2UMUx5wqG8QsjHIv+CDRlD1ICDlmgv5neFTRzXMy+B31DaxbuMJR449ibKmeMyET
GDyp2TeQ9L/37BXgmNnXdkbH6lOtocl+y1MMPqB1+OR7FTT2rNNN2j7106QU2DyM7BkCf7ruPQC3
yF5j6lxm1HSCF+KcOoEKGa+CSLGu5H5KV9FtRaCa1Ls4Qlq3BaXZIz17e/HB9OfRVMrfSPsEokrV
gwnUd2YrHmZCuT7pOB+Z9vIdDgYqR7Ty2jqcKF4OUlBX+Dipq+hiTdp4YjF1pkM0KXGSQQ75EDVK
YwtAuHUp5yf+6mVpT3NyZKC6hSw6dvrfI1ePDl6S/jqKF0uwcOBraBC/a632X6Okpp/ftnS3+fFE
F0Rf6t+DXD0LbZMmGvF3jZXRuPkrBxlhQ4z6zubUGFvnV03ysSq377DUiMoPPtcI/VWJuWrDWNag
4LzPW5poWm5o+dk9c7b98k6vj2Utxg1qErL9NDoBe0sPi414X5udFmR+xQGgpfdY/k5lrS6Y27x7
tsfQHEhOXkXp/ecZB/4emkob1+Da2PYsERDANlhd2CAzGohZw3SbyLh6bTcR6vVktziotbKP/eCV
Bc0I9J6PgHhy7tETlsJegApTtvi1UcF1IPEYyVuLHRqYOjrw/8UL3LmAcHkiF6Ysu/gg7Gy0isX4
YqsKrPicef0SoY1m92nE48mLeoQl+zF1W9xVo4oLq7aME1onToOOo+s3JTaDcbIi5iKI+DikaX7u
iuVpTyF+6JHWR2wjtvijw8IX4juHRmmLzBs++q0d6v0HWLIpGYBWFPz0gbxxwslnUSYV1oEQ7jCC
XVI51ht+1h6l7Xb5YVAhOX4OcOWJV92zxqcQ+Cw6NzB+oHIfJPXSoOmg+gMCLaJUecPHOJht826i
VcV+inKhBSk0hpDM1nLksNgi+4yrQdIhC7qM07rHujJO2ICcMXZBRfXuRInJjixw31GO2Fb/6/fA
KOY9UQvvBxlOvyx0yEWghs4FJvk8e1Om1rBK/Grv4unNFkWWjN29RavmDJgXZNHznRCfk7H8+Qbh
nM4gzHDfQAU4HX5jwKD0fC3TPjK9Fhz0D5WbWTMf8n/3zW/tbOg/IcQLBE4t7GDmyFqV7z5VYsDz
jJ2wyM+d0xcj+803oi1SoyA2FXKy9qFi9xM7YeJacm1YmzGgsbXpgM6msv/q1rZEUAcy1yIx7sjv
xY8XaZP34v2w0ya5yj4uZAVIYwN9XmOa76Y2hw9Aejz3MMeqWpd25QCw+vpQU7zqj0h5EYx57B7+
u+VEg1Op/H1tRoHybYZTRu8oyvUBXvJ66sDii/XHG0LFUD9Gh+w/CloWVBEdGlJsw7gKz8hpA58X
17e4T7jS5dz6ACgPS1zKAh2JadPtVfDkoULcY/4U+WY5lEUj+lYfwmDWYVsDyG6LrxdZbLifzXZn
sIg257XzzokoE4jncOI78GpwYHSO4MDBhR0V7xK3sMzRZWO316xYu6hF6L3t3ft1/X3yAO3tC2Xv
Zkn/5/h8iZjAAXg3WPEka8nIP1GCXiG9b4f0PTQo+zVkq7c3/ph26MXK7io1WRSN5bJ9YGZv/B1l
WPkGVdFCrh2ZecWlx4BvUIvh0ulj+fCzYWIXG1j6F/EYNO7S5Wit2rfEgwgoJQl9EyObIr8kLjL/
lRK8NY7Jiw+7dmRUtKqEXkcHccjRVOco/Nk36emYm+BpbpyhWJVBLGAWj1mEu8rvNYpNrvIWDZvy
fNOrrWfvTXJJzELIxHDgsY4A1gPg/sOhNC5+GBjM7h1lfhrxCCL0mvLt4btFpE2xJO9FF3GK4Nrc
zXXEy16+3hZDk1m/MoD1tW5uo1f6m/oMV1zf0jeztXb1v+yUBNVTGmr34fsnmu+IE8UY65EngKY6
2UaPmxiVkEMsNQabjA+kKTxxA265WHMJV4BrSJpRpKwKdgjQVOqntQuqvBNls51DSIhOAjp2/4+A
R4f97BBn07SA/A5WCXIlJY6fG/IN0NkPD5T9UBSCqPDCAb2JMxFr65KsDdr3BCfJwUvlubJfAVJV
HeGtAOtE9gtkSwdKjv0eh1CpkERjNUdGG+WWDqGYt/x2d0n09Xx5nTkMn+wP3H4Fj94SOVxbRAhJ
yrFDu+AXYgT3LSSGpopyzi5//KBbGsuth8GohMcL6+4uYDG1WQvAbOvjcx++/cx9EcSLfjVhkvPI
CKRmBYvfDlOI+SpQvm5xhkLilG8orKRXCnGd151LPyJWxacQZ/VZgWYbq4f32/vQ7N/pvMABvUMt
1JICZhcvZgkE3r8/2cuGBfmh219MZK1YvscRhkAnoASSunF1zwfXjE7mzk1iipKD4PdZ9EBtUtOZ
jTqTlbScbIiEwYPtFrmiUugO5AUsjICvT7e8kKdNl4sXnrchbrszMtTkT1odHmzlSsZtw2C3MsNE
y4C88dtN9OvgZRl7iyLkuvQV0zr8PVu9V++HZFMNkoLz8h9Gh5L+WTmoLj0B7UpTNw9QfJ/m/uLw
oV6UtWarQvQolmAJ5INmZYwxaVG9SwdyRqKYYtBl30AqNGL3tsAyQEq+DwiXPnEd0WRK/DwuiBuu
Ej4eIdU+8vKi11uaaPfdFROq7H/nf6zsmKqDCdADOgYoBY+QcuQTmPJP5Onan3vPhWF7j/IUtCQH
RfCUdbvwD04MOsTW7Druegn7XB71PgkGSmar1+JfFHfb0twvHTZBIBszmMzVCzVPf3Zar9I4Vgg0
mrSiL4U1gxXDLQFOSG9D83ZpEVj+yw2T3Qj91Zi688PPofR3Ujz6Bhxr/Hz82obwSZB72DIito5j
47I3c/d4P3qpMUglJaoHEXAi9qmsjXhMwZJ8MxRl7/i9w64xGgXy053tMhUxB2+1syI2VKir0TtL
5fz9ZEwYY7eXCSMvDHZjWagHD5njJ3oeCY+0wKfVzN69q3gk15f7F3xuupT2bfRBhX0/edgH9SaE
SMtgl73zCABBj1XPbY8LAcKKGOFhrqRq46llcg2eZdnQ+k3jSTrsg8RvIn+zzH+y4R59SrYmAVoX
OVcdTDlYhQpM0+4PH67OGirXatY75sSscKMNmKzNPVFbfCUCoIsZZodAJWe8E5i1Q8ZRFbng61re
wrFPDSjetBP4poscTpbQo3MbGu7i9I06dWfrHTM/oX2T8hAKJnqZZzoU6CcTBH2M/L7E7d/0K6kA
JRGi+myUyC5/HJFSoU3rv43hsdYvqwOidQkDYVr9EZJ+4E6aTBvjRirzCTD4HCS/fsLR5pfZeayo
j0Uxu2sURQR5nnD6uSkktrJivBJpVr7FsBpCVSt0K7xmsc20qG+y/TefwDOboCLnoRCQH+BrrWTj
XgUHgM3zULhdCX6FvFQFvz9qvOaGEr0PwR38K+UKFPmYrNs+V/wPT5JEPlu0tpqRoe/2n09n+WMC
1ztrQX2rOJC5krur/DrBY0gya2MMQjygaPgx2EatE3GsVK14gWbBRYtP3QgNxVMLl6LD5crBy2+M
HDr5x87G3vKVYxoixaW04tOMUg7p+G0EfmZavP16ftVjQqzof/Ij/XfrjqS8eXQuA8ZGho1sU+2+
T1iIjUP84SmlKx5u1HQFh8iSflIjSQ80uzZ3I38uh7NMEZe12u6bIatD8BK1/gK8Stzoah+nGeHi
Y9x74poII3nOaxryWmAnjny4grkN4h3s4w0S/rxqVN+0GBEoU9RWGgdaFixFdacvwwWrGjFMNwfE
3jHoSTX8iAWrUlaTzij9AGNgLBSpm4iT/R7fJQ+EDab+dcL4DUAOYk6LEGn/7w9AOQjkoxsUPjiE
BDi6j/RZlWY7DngpXFeQ1qh/xrndwdjqCGhjlI9+8kugQok4cgKNIL0CuepTIpZYMmIq2VDyGgRh
OHFX5bdbIWkspRAv5a4LjmlG0oTozFY+mMGq5bLrCmXjMA2W/pYZfg71+dMo50PtDX3Nf9QA08zy
1SnFraW6ZXYNMAdw1mlnwZnhII5RZTsuFI8yBCofRfmvP9juxafVtgUendSPGIIMAqu+H0JyXAsw
ueUeMDYMk4v6Rky0XkrBRAxLVX81VGOOcu7bbf6+lbPVDZUFhL5Gf7euRmlVn2ZGqlhRwt5RukvE
poQKeo7KR3wupCLej30jdCIHULXSIus3HDhpz1sE27FD6/Ww5eHm4fp2A4EHEbmCltMXSzNMVh/O
9fIpsjb0/8i2ohWpziOBJOZtNfw1lPy+b5c3midI01IH3hQxKWfdBNLCrQuaHnR2w7vm34Z+cs+K
FSNiaemZepzCbL618PqnIxth8IlBuNCONzPUIF9xmRFEI5SKB8tbEyJCvQudGHkObdyodGaTkI7r
fUqjDHgaJt7aLMoiHy2kIO6EF6qiJNxcOBgyYeo9TvnFwBQds4w9T9P2QRzZhO5l4C4zTCnsV8xT
+/BRT8q6vHi0ZTExxRKY2Zf/6FtTUNnYSTWN9/AB7oKc47ALymAsP0zuk4rnRrWjyQc/AYHMZjHU
LVJlEGeBnw4eR+FkPpiEhyi8ooN0/FcTcpYtKcEnQptzl1RyC8Dl39L7ltIX3F8bvb7VU3Axrmfu
lovJniHMpon42kBt6Ndtx+7hX7XQgxYsUBm1WeMjZTpg0vz9GjzWQ21Bw5m7YnJQdtmxoJH8keQb
XCdLNUn3iJise9I19atiIuIn6X8OPyaelfbLDBuyZPM6ZI3nLDAJnDntxm896nzKC557rsjW6bNe
eiY7GAxSPO2dwQbvdsGo96CHSXdw5j4+/N0cOIh+YiaPmJDgYgFtuN4qYh/hZlYZ+3hnOUxSA6fG
+b76O5uQAMp1hOxxip3JEDDsH4Vh9KZOgYMsG/K0mQhOYTvRFCzurTgy6f0tDiFtIJV5abmmgBuW
4Mo1eFyh0+kPIl7RTVVw4qE4jIJG8T7bxnp6UfiOTi8JvtiOODy64ka+tzJO4fD3FaHE+uaeHfD7
SChHqROq2ZnqHtGpYAAfs0XD7If/PZE227pALzUeZx1byQ3jupmwyYu2/wtFGyKHExjkADVO8BNS
OBALW/gNE+EK7SE7fYi+8gkG/Q9+Q1V2uPLczcJGlhKm3qS5uZ8X9R2XSiuVepCpyDOV6ddQftt3
FmeDTTQsOfmXX+V/AkoctgvBiuoJPsmclARPSAZbGWHsL8+nIKa9NhBF7kauCBw0q3yRLg61ztsG
tT/K74C+6W8oeiOlpzFEUAQ/03thYbRG9L6oYIMRLGPXBdj/auCuYOxUgSAcRjj5l9pXGHOna+IM
+w1YJtUJqoE/6Zm68p+C+BSYSGzlA3kx1J4Dblqlrw1ORlLUNuULR+vpH1GJw8KB9WGKiePNkehL
TVAbdDiHoxaPfHvtmjYvbQH4B/s09qNxn3JHu+Tfo9x2hN2OR4D2Vw5eoDgF6Ct1p6euGj+4TjC/
CNqk16+P/uXnDlEgleKNdkzq3iqNU7ABIDJGpGBMdE5waiyzSLF6aNkOuJT20hMZ7FSuQIn7o+ey
QcxSs4H3GA+vdzsm9OGiTP/ciEeg1n9H5h0Ex5ofOt5Cwj8xeV7AajP9ewDs5yq9WBPUulEVXTUF
ArhcHdq0p1zcKAa6bAWlZ1+iZ3x38JzFFtH8q7HqhHUVfSOPLDaV9E62InOtU+s+ivVsOzhA+cCl
QjMbkRzYYu8he9NUOXrh4zomQT1PKXIr6a7103ZbTwsbn6H84GIgm+WxCrYdP0BVU6kxa3+SmkE9
ZFD6Oy0evJ0goDgBasWtmleeWD4FmeI9O67zQDSczv/Gy8QH+okCsyooGWrKMe8JWRV0WRI83+6b
qM7X9ajJUx0o2IRa8luuzvRIkMss14B7rmVH2MHrDOw5UXTYlpbGbJlJiqmwm29u65iNULPTs8jH
SDask5gBwCuAC/Y1nJogK+sV2+lkjuoY+FZkqwvvwkdh3kHdliK2XxQb3XMAwcP+NCnVlEfFkgQf
zQUpupDaOeTO9GsSWJiPHIxXhLSMyxQ+led12MVbRyujMNxx2hKAnUG8hBU1cfeNdttxOWG792oT
QakhNb596Y5JYhg5vF+R/CWGYBjVV6b+gczt3kaayoJtVNNDGrc35pbH482UR4M8VJdDr/X8YWkJ
+QRBSmL3eerYrMuHHXWK4Jrw4d/zYZVcIvXxgzy7X8V6chRdl8Jl77sHudM+U1NOqdnB2RYHHFKP
74kYJ7W3+KjXEY31P8+2Our/siLP9FdGEQZ8EVE3aqJEWySOA1UxTC99lIJ7GpdoMjnDc6zaBsD9
9LbgdPcCGKSoMOTxq6pxoyQmJZqAvmyovs6Sg2ixyHOLQATlcbn/KQFjH/pHsAXV2uPqNByxAWDj
FumeleKDSUFgf1DscQe7JFXe2tP2lcOdoKkyzuereLdwtCB3Epm6U/ALa1SoUhvoLkdJqvA2sK7i
JE+qZxeaKPXNQ+zx2ejDb7ms4GNkJQAdEul8e5Cg2JblyuOUvATwfUHOfXLdtMpGrgnsNcPGooqP
kn4VtUcqOlTCVwWrM17LYf0XHBRO9mEOQ6XgdnC1/2scmI2pCUBR/MCT6PvUf0Cg5jO1j8S9Divt
J+eg8yA3zhs87vtJYqUXLJ7oYJcf6qjO78NSRjhIdYmOjBhowjHoOMvl35eB9D0OdcgNDq5KPrFO
QSLXgfu1hZASPkEQpp+0lXlhIfE9mMAuBV0sCElsPo2iq44WF+cqifAsujWGg5oWX3EzrWeGca1U
HW8ETMAvbsdZtQwu0MVhSLkNrT1Qau+I8JxM8sJo1a0LGvEhb+3Hz3JPBj9V55GNowPZ/ol2wAK/
t+HfMTK7Oa16p+U0MSlHZQ2POxbxLvXBaV3t9hmEXigmBaYORtLn0RNjdcFWWEy3pYj4+HxdXbcx
1wl+DB3f3ZLWO88KytKR7pf8iZotPc9P3DaYx12uKEzazXm7k4KIvOYNbyUErKysxTXutsUGGIGP
x3UzlnLXA4ERFEPs5TBt8a5keBeaFsDUbsV6bcGP6DnmAgIDnO2gw20tVneK56YExQsSTJWCV6U5
NojSnXoljqwcVRIGn6kUIVUK0/wX8DN3Vvc/NxOJvb2RlfETWPsjQtE9xK/ezHuWfEgN5+DwvpGL
v+9DWN8yyf537TiZBU6htvZ0nxWov1kLweEGaPNYaAigPcjSLOF8XUzhE3pPufepB7R/3NkrgnLx
M+ZTFf34NG57rcWgz8AARCVzFFqnVxVL0S5W5rC68ddw/EVhEOY63Ka/qkyQ2h/ZCi+kB/zYTbjo
mGtLrQmajapYp+gkB66pQdSNdm6om/ImEnc8uIf8Jdrcv5s2b/e85I7syMPZkvs+gi6Fe3WpLxMl
eehu6tSYFNE7iiTWnBKp78OAnz8tcmY/hh/mfmM+De+WRfhGj4U5Y2R3bKP10gyF/LUhjg6+VF33
WNdEJM0CEVIuEGT1FmmqNkFvWhHftGF1v5Mqzloh3tCLl1u5Bgryh6AKnSbYLMI4Qxrvn33DDNdz
5R3yfkbGs5NQiLjlrEcO7RXmggbxjUPrZBolCFd4APHKQhVm6ojTQIcnuKYILyqt427JquX/RNy7
Q+NjKbWrOUnT2cOQsdRCs0p3EEOm7QAk5exQaTtVO4IwXqhn6V1GcJz2zW+7QpM6wnVHiu8VKcuA
bxYrihe2xbthz8ID1qDeHI4QqdB2A05l3TrkvAWsGUR0K/5nlsw+s/wKLUfHQkc3EFgsRB32xCbb
BAfm5SYBkR57U80b7PlXQaCArTEfE+DNy6D0Ww3cM2oNl3ufDkHILDMb4l7Gt4JXHvjGV20cdFHE
rJfOHylZWxIQljGvNUbgKwUy7VMJJsZLTIzAlhkrQuE+BeC5IsuGHQQgzWhQivazxVILSQB/rLwV
mNFrPJHeCB/jRcwa682LVdZTHBsRWGKR9QCv7cHiMlWyZajmAdQXrrmvCJazoJPQZ6NUt9+YjXm6
YfsBmfNqG+6J6cl32hF9Mh/HEqKK92Zp9o5NyeDcTM8psZYP/vXKkCOKW1WMijq6mkAfuk7GZb1G
rz9aUma7w/42IP+k3dQc7uy5mXvOpWzhoYE85CNo0YaDnqqw/1RrgAK+WTxlFb6EtZDNcj0FY6jo
+oa+bFXJM6rZre30SGlv72ewmskEEyqLqNgdeSmol77DDPcQc+OHveTxnFPJyuEtGtmHfZKz5e3z
AcomRCHG+fuIZzx3j0inENFlfxjWKR/33J4YzBjbR6S5xC4vfefEqMdXp17Y1UDRZ6hhNm3cMGL9
cmc83tmgwUKgbd35pYJ6586FhDr9FfRZT5xA0UPSTsbYudQfZtGl8WdmvpZNJGWap6+Uo4kb+SJj
XfcTBjNRmyQE7TxnglQPZrCiKPIVYnGhBmu5UgcjsM2LifzB6DdMxsWPujrbyJ83qXOK7mQQ+ZF5
E5oXXPxWnWeTV5OR5bh0KydfjSwU4kC/+21nSPcvQ9qW4AzKsm1KYfDM6KATeWNkiVPSVMI1YaIb
TfYVR+rhl+MojzJ7A+sQA8DvHt570uO3v8KkXGfNBMtLcMyj8pO2SjfqtbbHZGm8gEFBBHWMOj7V
trN9T+nPfAQqSQo+P4CBZ4hvKaH719ixG94sx0yk8H3HBIwWBj9T9MqpU0F9BHOd7u5KC6PEUF3q
1LKi7QHdQTCV5aARG3vxYw2imOoRdYprTjVPFXwJuX/yLuxOdylbNN9B2UN/WX0LBeqYS+1x9KWK
Q1jiIbJ2UE0g2ZYHL/Nbj9PCNtC7U6a6p8mbKppAK8LZYMgLu33T39aYqjxu9apBtkgWkmXuW+P7
wzh64OAnToSYUyIM/rl7AvwdeZsmaBGlFNDW7yFET9PBCywCfHxkbNV3uPYbl9UxPibJ+TiAyRPk
FbMWLjhZdkjRdcU9SSi3xuc8UbLP5Ab87F0s7e2cxZwDP0gY4q3tB6kGbKlkBiwGs8gBXsHSx1IN
owgyYojc+KxgmKcsVLLhTZ1x2lYjnQC/6Z79KO/sNpkUlLEd7omipkvLSBMR1Cu+neD5D3hkkCSH
aTIUpSuIRA6Tyimp9XzsidR+rQ5U0s6O7Bvgp0NLlp2r4TCVsShoAhXr5NygUKe/GmV1lFoImiIn
V/dC9k7KswmKQgvvBZmJ4aUl0FUfVnZaRn6wxdl/UbCdhJlhKXcS+qTnHjj9ALM3zunBZbKsh6ka
TBg8/h9k9eD+fVtsJsoQoEROk2r1pWXWf5jr858auUWrbr5aq28P4TL4lqf2SACCB/j1M3lnjrqa
UT5j6ZL9nIJWuTrkO5N7+XVBiSIRwhNpwn6NJx7RkJsl16VlotL/sc8RBoe7MjKCUCESteiY9s3t
7iuFdPk1Zfs6ddvGLGSwmRne1wqDyKh2ibdnO8QqElo0MvAKRJ/tsToZLcgGWDOerja1upwkHnpc
6foUuPBSFKPahstGfeTiw0yCEPNyfVyLKrXXcfamJ+ug5kwDFxe9gPJWI3yv+xh8ZN7gTJYG4gUY
/zaCrP8z/vwrqLqN7Y768ToUT6EdJYFCPhfzxOORLfhOLd3bMO3M/lqVbGPbf4cHtJ7sfwyw82JD
WGnpwyO8xf9Vxn7ZtS/hrghn955sG3cHRd+BkjV9w8qhXu7O7zVn4IOh8xG2e32WYIZCJp5cpySQ
1eZUMAZqWV7Qn5gDly9eegb4jI/y1QN/cBwwnGFrumAZ0qFW8Yobp3cUXa8i2YBAZxjzQsM+xcJt
x1TCqakpBvghrO+a7J59arriHwkRkSNQlU9ue4+/a4oOF+Jf2Rv/Db9kvmlvOpeie3VoyxYSvn29
3QSuvu1UffW4SbqGChH2A9V9m21piypUo3VIou0rG2B7ZW9fjQJSB8ZtDcpZwBUBlOKrbdOIOk3J
wutCRv6vb0j5R5gz/XDwn2/e0UVCgdk4XlfEpWrFVQpoCGEq4tkOiZ0MiXc5cV3K4azUjm+PhnAO
ZppRU3uUnJLbuikpr0wZ6JVMRUEYYcj/+DTMI0luuUZC0I9wPt52qj9KsD1vq/nhTazRvbiRaOm7
+Ps7KnmHfMbU+3VPwv97dCSRpHBLKaH6pGUD6OM40oh1IIkaLsmUCOhmnolmZQF1zYXtjctn0cY8
GqRYZBbv2YV3uFCFBScTxU9aRf0uvvHPsD9MFOohL3NLjBQgU66dXMCf1Oy7uMNDMl7+Pe93riTY
XnRf6Ea4MQUsktKz7Xwziq6G5KmvsERQAY/9/IaIJN1Q5Pskvpb5M0XzqCwxgblkgqIE2MmZEDa8
+Bid39nr6oxUHlCzanZc76R8WI7CMlJd1LhUGelao0Yt9UZSW1jqFWnkA3EitIDPQaSWJUc3o0x9
nO/D/3iBkjS+wUwWsP2Jwpo1wxP8mLMDMsjWOLTvq2Eo2TbZ0NemYhnZLEZKBsL3ID1tA03MA7Pm
KD2EMYtXPBmW2t3Hx4QfCiM8/irzPkCgBipZoT7VmUAdOdd3/YfICK+J3dC+ertRkgwL97T8EnAX
l4JwAb2yREsI81OnuZTlP+mU7VvADW1ZhcTOA2Z/Pnlje0eXpi54ilywiruj3fgPg1+hikUjlmyE
9BixDdMlcK6NFjqO9schdytfYfClidXN9BODjgJfrQqPodSvaCqGxlO/1IfKLsEDdHTV45I8bVUq
d0XMa8QxrDAY61mE3pCMoBDa+A3CtyJSS9p2uCP9Yor2kR8TYRXTktICihXk4b1ZavUIJR4imfKo
0OdHKmLlosf3a2+rsOIYS4Hv3M3WdO65pByE+11ZfFIBK0+yKSJ+a7M9TKqG06C26BNZFK7zn0jq
r0jLCWlyPV52u0ucbGFvc4VytgA+66CB+HzdgNLN/D1l1vEvppUWJugsImI4lusOR8HHCWpnBhSV
umVAJRFpKpIANnzvneKXT+UKrtLithar5HvuA2WM2Vl9R8VaIPIY2DWtjYGQPjsrjuG0h46ZuUHt
zu/gcpq79qD+k6gmcGMJS43ppE3n9LnOUP2p8Vjsu2oQtR05N3Vj1wQCqWk7P6bcvj9SRJJFGViB
DJDx7sbUGtsc04ipX+ry3aHPBNwY/qLqJ0iDRZQ/tQj+bYsXoza1kqZJkjsBs58HnVjEjCeNJAfi
IB5E/XE1qlei58VeR2uWBSRYHjSL8ZGI002X7zqJAmYmYgc5x6oiz69SdDKWLro9YhUYZ0b9lEsc
GiCeRPl4eLkgNErY/DA4dUIvxU1YYpLAr1vteudEuOCQZuB9D8y/3y2Au7Yh0rmfmZOePhK/LYIN
JP8p0GnnC8xMglJGNjK/LMYKzp+qYbwQ/bOjGBKgfu9R0BERQ+dLAuYEjagZT9gO/Cf8INpWJmgU
goqyk70bxH7TMNTfcLBrpzjg+YCo4Dd6xnBl7ty8NTGWqOLA7r191ooRXkQT3Z4bp3ExFfkz8EKu
XBEsexm7kU3yS0/mfKAV45zz07HPvGW6CZfbUnWxfqOqM3gS/v4IrP8ojGTeFLbVF/xNlo3BH+GN
NRxwuClWLNAcXZkS3gEjGbsPpKa7O4VMiTxU2xV0zv29C0DMcAQ5DKs8IeGpGdLiD+6b7UwDVrOL
toV0tsQI3f/JGkVbEtDCKNtG/WTcx7NtoE7NnzJvzdv9b4IiaMRyvxmF/RukH2HsYeX9B/SUgOqp
RJRMuXDBcgEfRIyFH3DKYbmkB2vj4YE5ZQ4uogH8uwaO1J53cJoIkX9fkb8XPajXxuHD6SURhICd
7OhLNDKpu0uWHWwaUb9qMQYdDEJtdJSgrnd42uwUZNKLQWQFeRp/BVas8pVcrVDCeBKMNSQbqOaO
VuvAs1N2ZUbs/LmAvfEoDYYysA3VxTh9x502cvSCsItmkMByQFKde7Q0SzmIH1uu686L5KX5rm8t
BJT59KravV6orDUtQWdBlnjnfdgh6IuJ5UyJdcmPZ6vX5k60Vwqbk20y67o0Lrz8wcQnj6IL0uuI
e0js+PGlFKzVkLbsuv2sbT+FlJO8Yw6qSGl2hpyN1aQny1hRAEX3Zy5jLIymFhEwvZ0X60MbmWCA
yewBbVpgETx//cA9Sqf7doA3Js9MGzLGQ3mGPTNpOyNyZPqHFEmcra2aAlYYst0vCmUf4RPTCq98
SEethwgO966JwQ9Fdbuxda5ESZjl1pZzxV5I3Y7JuFRCCPKfzT9WHsd+0oHFAB4vgLdmC8fepKTF
u+CMV9qjcAAswq/oLCgJ64fzV0v4jTECCbk3+MGHc84BwAJjOSjD+a0Pp39CiI0MoGtR10NOoGbW
zKfY5NLLfhOn6S1wkESy6jXaywuJNt8GqCxgAGbSWy6ZYTbHGhT2ZxDEs7VRbRhrToey8eZOWQDH
yPVwXOPGwJuXSG/pQjptS4oGJz57mGxVAdSAn3YE0I5h6qlY+QryxDLLb3Ra4iwZaUIWxN7Gjqta
+rMyuZVLDPieYnJ0J0qYuH9CqpQNcKqnxsy/mgE5PgsQitQKWJ5ui0wJrRb1DXcyrlZrjb51i5xQ
N+CUvUFJFbqOFPCPRddI/CFfgWU08HNNKrXFfuyRbXGhFo+pu6OnFccPGg97F3pNxaVOnkSAPYLy
L1aKdC/dpbUwD7VpuiJF9hXUF8y6bP2OAYp3G/2+PhiqBpwHn1HzBe/aFNqyTqJh2yk52iFNuejo
v4g3dhOyUq4XdYPD85Cd6bgCAxDB1Jdt2cz8TJnrUjh6JCDumN7reDBXWvBduFvyFdKjeO4X6xQW
zkFvep48GI9EEIAZGv0joQOwdji2rBvSgmuYh0YyOk0yyAMK9wQAGWFvqCVxFepeukbjxlOomwEB
sj0NAaKJisds+SfBfZ8V9FsK9r6PZoX4VrzRxHNfBwqtWXw0lLsW1CfB+7JrCJ67D+lnx5CAbKfR
2IekcAlB9pHvp/jR1kJoFIudr7r0FYI7tnM3AgtCMXYnP5//GNw35iSshF0IX3vGBtNL7486otts
Id6MvaHTK2fUCTCQiKpQSEDHdIsajDiN1Ft8Nf3n8j0t3iT/b+a4JaN+JIGUvzFYiAYdNMsi2691
xeHsLpe0pbUCwgC/Iephp3+PABDDyKzXBiRq1fmRcVThvnk7gymwp+28HPF5/hyUGLZWV3U+hFHc
2RKu3ZdBOtw+p+ZYfCsRadMWf65VmGAbbZ/SjbqM99zKJXyLY8yoCLR+CzyRDgvlLqd8dhyWpGqj
RuNu9Wsow0xBXW6C41o0+YOySS3pZ4wv9bYY4Ch+UAW+hwjoKPlPJeYsCoWjo0/+ew5lSr8bcrvV
1/Xl/Unc/KEo2Z62DvgnzcpI7cQrL3LmbgcncOIUYiB8UInbY87a28UY4jyTp4Nc4x1R4I9BmLpq
OTThE2Zs2nm3yTnr+UWsXF0QgtE7tIia1inNC5vYCW/OjB2fc1Y+HjhrC6YkL6UmHl+xtRPJqXUZ
Wb3J29hNeFGip+DXo3RfBiLix2vHNc31TBw3ZNobFoM88klgPk1pVwEMIhpMyhTb2zFVpkpoCgJG
xBhiwQUBftw+EWMgjRktZVRGQPaZXdV+/fckIeRwDh/Axg9egxk1bi4Fg5KVB7R0tw7PA5tyizsA
UYN6UXTqcq2H/LI1UUCGPlzuwEVz2MFzotnUJ/U8sf4WGnEH4oTRSqfc3wYHXqWdIJ76SLFCJ4I5
CJAu2LLzKykCZfxvTOdXgpJcXx+iP6p8XTrf1qkUhb+OFRulmgnQBwEi8rK4wj0YAXcY4648Z0B0
KunBeoIQ+ZkC9J7zl14MZvNHN2R2Uth1wvT5DNcVPs3GgCL4IB3x4uc3bzYsowD3fqSbnFLGA+Vg
ziaAvv3JUd8EMJHq1CVMwli/uKBV4P2PplAfmvNLWXlfTQGY9nRotsI+JL9xTwPOItO2Y64vf31s
aSoi6zTUQJRrDzoc59NJOQqD8p6xFMWCsRSTpzm24dcQnOkdfzMAuijLmBNGh1hUwPD7Z4IH5H/y
FlbtBf1HQHfwvYaeT6q/o6Unw6TD9yEhOBUPxgdAZBevxyTU94XyvRz/j+5OYCghqtxIXBvRT+j6
Y2PUytHaSEVai0eddZ4SWNjTK7jhRVD8r2VV89PHMSGT7GmCiYiN88aXMXJwLrawa8HWBa0abTJO
db75RPCj3lgOtFmY6sHFy5xYK1lcr39wU0hfyL+usDrIZYY7iuLvS56hkCKZeaPC+h7xWpMvWoCK
dd4sU+kN0q970xlhYsCYTHwjV0fYJWOKw5pyxUcvezLpqDYYH3nCsrruaVZy3Pd7zGBKipJoh+nT
c15G/9XLql5wBPu275zNjqA87MqAlHnAR2MhhpyJ2tZE+OrEAO0y6D5eulympswVYxeuFgfNP+z3
vtNr/9whvNXq0zqCVsQ/7pTzdURW/LCqJajVRbrUjXTroXsu8s3UYphNR0wMFpqwCUbTiXfocuIn
fHCjd1M2Uh4lb+WF6rzy2LOIOgMtHd0AYph4J+83xFjJ1xqaG/M7wenoz3g67i660MmSP8BORcva
xh/G9GkhJjsrlbA+RjnVgQSJLsmakGbIW8RtjRZSxolGw8LYPlhKe3cUZ3l8FRvnXXbH3TY7WxXS
fzFeMIF4IHUkDK9TMUiVVcKRoH3IhNDgffMV/0Gjh6RBAi1A5igqJiWZtrTTx6MI5irphqdGknzN
SAske6BgssbDBTRXAjhmlJidSAIfd7H5ro7LQWsiOAL0KmGcvj+G4kHbLyXH+IT5ywKopX3OwQqu
G1cb4Oyq5G48xChRmt+U8wbIIRpCv3EbAfTzmKPF/OLvRL6iZ/dxzhOdAppJTWlDntqTGtMGT6LI
PKafruc4Qjd4GooieQlZ7kPt4yXXsAOUww0A5S/eHiRTliJiqQ0/IspchTOxHG9OAXt5Bu8g+n1U
6Pc+inloAaMNn9iizzZLxV2ooTelN0svV2chvrmDO3yu2YTv1iv7Fm0g35eG+mI38/7VucCAhGQV
WhlUR1enTZDVPzqlT+6iJyANujFqOFAgXNnNhRg5lIKKVa9PMuwPcJgTWO/w++1PtNDwDR+REXid
Ub2VL0nihu3MC0YeDabH3ff/NeWgSV12WFotx2xWIHJKa8LX+e/TODBtrMZtoOBGDZ6ScB+8YupZ
s4Zf69b9kX380PMJ+1eh3AX8+GAkUk+TKMKA+xixWEiASUPY+u18WSAuiwaJQCSXXQGXAy6g+9Rp
1urKX5P0k1bGxc4UKYNlHffDRuwtsdR9K7j3LANwZZHZLnbKkFK1tQzfbcjkNOUUrNDein/n0Avz
zP4pdaDTTP1K0NRqTRWpM7UjraxeTYGnVUlteXdqseUQN0yDtawc3ohwntDUXB9XSjlI49KxqaGA
v0tPUPHfy890KqCsxCjsbma+s0AMAHCeFxFPJFefs7ZJ3A0ATaOKh6+wva/a9QjCjFM1Mkvg9lNC
s7JWTqOMhbzdo68DqJH01zR0HXqYyIMUiKGdL6M/FROL2BTjGfIjreSley4Gt3cj0W19sicLWCLT
5WV1G3DHmafesxCzshgHfn5RlsZqmnjDaJh+NYOa6p4bSTp0Z54TUWgY0WlH2/1JdDsYKL1nLbrW
brqBK6YonOxmTB0FKo1QEBN8Ey0hJDzc3uWK8Ex4pXM82v3Rzu61Im8hMVC4cEq91MsbCAUaRamI
N/eHlLnKNlQTHfgV8dt3uM+V2OxbpNe0tLD9VITK7zRjpjHgBdt723t80/cOgbtEHvkdyw1Ii7m7
EkStHCahv10H6PfYxbC4WohG6V95+pRD7t1MHsE3Kr6TJbEyAWqmaE+OAuh0gXOWBTknkT2biYK0
G9eTSF39ACX8mACNnh+8PYGaB+n479wcrLKDY2rzEMP5iz7DUJBo0szgXNBb4JLa+NF1nduVpqMi
hutAfrLsMINvNPlacU4mhcxM5Rzw23yPhohB8NwTXICd2JwgC/PLP3SNj+VJyvsTyDyNjZju/UpM
Jp5Xz7/wpl7CFltqxnrQR0aSSPOon5hj/TpPNjU6U3j+QpXPTj8MqXYe21WwzcJW7JrctTcXYIcm
ly8OxEKaNcAft5ItvzZ9kCukb2CD/Px0ZfIstKY4XTwE1CXH51KuLlEzxwZXh602clmxl2s1QxJG
h8Lli0vnSf4DIyqRcOQrcbLW6S7qwpH7hLq4hWz3QptY5yp/tuF5EerR1I/QffbbnozWRPMdvTmq
w+nW8bdg1seA38nG43WOBdcxrsxE/2NLY7oUhU8gFzqBzet+eRj3OWs7mJemx0BfneKT850v0AKR
Dvki0gphC5ib+LX+MpixkqGbAStxblnwrx9tRaOS/ZHBLiKfh7vQkriSwp/cnoF40gVuL1usk9nw
2IIb9OLEQfn2iGIchYVtdNOUz3GHaV/uccrbwc/Hx91ye+89OaNPvCnQE8knelM6zuiTX8PekLiA
ZPUbeczIVfxcYtpuX1RFF0v/oZ3gQwMw+Qnh4ecOt4p/M2qgkIHGbu7FFaE3GC82I+PwBzlgbdLG
Cztm5rLBIQAlg77zFCCOlQUTkAATlw59fewU5y+vt3+RoJU8ZbHlrgU5jMn4fESJcWr5SXVF/lDh
dwuqtyfCqOOk8G3ialO3r7v14zMJfTqDQt+PEdPajFlv4kL8OaU2xJfmF3LVvFAe5BTPiJnOCQRV
nB24L/KwjH1ViN1tLZp4BsWFYeZ/aftKmom94PjMK1MJMQyLgMY01BwpkretVDTaCLNtEsgH7Zy6
yy4T9xn3Tb8b4Pxl5uj40qXAtmaNJW+XyyFngUjKiryERvyW2+HpYOzRUAElujPkWiwDH6J1sSB6
SUGTt++ARskPDwwVmQuza+VevfuPYloq31W9pAUBNVQlMgc4S4pavSeD4Gs4f4NnAVBGFeW09mPu
ncxOQIRf5/mI35nMBtPfKuuW7d6pfm8vyg0s2jjyFqu1PxSJpdkfuThJmb1N1cFTlsfhuKRYn/ra
fhNWY3Jh/qx8F43Trg5qKnZDqcsR3pwAjwdMRwWrm3dvZzXeNWeQty2SEjg9t1uJjwmvS5Jd/mnW
tzagGK+AqAHC/eL9WQtsr5xH3O999/XOU+rtCzEJvwWftIXoZN/L2Mhx59KlN09wx3DSEfcCOWZi
UBSdTnmuOumIWgboENJI5pgfhL0e8QFi4no5mtTrHpyLetDW3bJSIZfH9pb6igo9mX+D7JXHMAEG
qkHRBa8tR3TylFwk1G4ksGwssoPV5+ofdeTQ7ivtlZoUol+A25lrTO/RUaXMW6yzzq+V9wXGOvvm
sdCLJrZ9/kZbwiTemcKTw/LskM9KG6c9qitDII/W9PPo2l3xdPh21nDAizM5/zfzRE8rX5v6ewUe
3bfhtI6fvrTKhRmfVqbQH9BPSEIDpXoby5ZTx2ems8gxiaCDk3NzfF9FhWhaHtyEPEU2wqBek3uK
C8aj5WuGa1Q9MBUL/BBhxVkUOQxEGczFHS5RcgjP1KfcNHmXChSWOjhRFGrsv6VdANprs8tH5/Dy
rI9Y2lucvbp1tNRZ6kOtDpwNisfOH7xyBCOUjtlzvYQKQOC/8SmodX9vBtwwDewkhz2pXrTmwGxf
BpFehxk888b8Ngj6bDb2+bAsc+E1DXIqDkrJ7PX3EpLCpPNgQT8Et5wSKSCtXrKMSOonrIext6gs
QkgsKa1J7zGpHY7+4fTrW+rDl5ZHK0rLJKMkx8ljxqVHj1L1cHb9vzUw+rXalkcj03sD2Xz4aOwl
uMqpJjZgBlOsTX67lziTLBN6GZadh2O23dzREYEH1Owq4ysWoLHQ/KpRJaRDP8ThpFdxKoiYE0xp
kGBrHR1iPW1RNysVdfvGEun293GWu1CtZhzYfH3FWfjdCTcV/ApCKRUL3aI+yWjaNvjFF3l0qPPW
ZmwoJpY6XE2mNHkRSjFvmgV1t/2cYQXF3wMPUo7qhkRARmf22quIMOuViSeYOiv3cVF1bQmnOcOr
gi0pUbhYyEd2ZhZjQFQchlycVj5LZkpQxKmmn9UV39zMb7GMxoUlLSjsQZjtqksJs1x5kZQjcaYN
xx1ehd68SilM6MCJR7veUFlhPW+jFlZGq+X5X/upZtePfW0sRSBpImKLtyNK5iwIG9yQgY1xx4JL
BRmf3NMV9nyFjQYgznA1qeUdcEJ+OcapQ0F0epD+6gu9iKZ5p5IVUUmTFI8PcVt2WcdJXvpj9iVA
VoqTkE8y8w3mepIofpzzfehaokJW++pmdOBfDEupXCjyIBC9onUZo2RQZINaupizgi7VKZ26Qsv9
uGs4sRIuNoMxSf0yBK4lVDDMe1gINlcpCSuADHM3A7nPuIBonNOJnv4ahoHJIOwkiUR43BahJ1ai
6h7zTjLAZadWsjAeCGW5rJ+aejmjw9MbOw7lE9pdG7t2mAyq4VMIk3ZWhYruEGguYgXAAyUhgfzx
evYfyePXs6thttPRtdB2R8d/4U9cig+AS6y0b1VZ/xkOFz9Y5GONfm3KU3kUcDz7r8Py6cSiSZCG
6t6M2QBG1ZWA+qQHTosu4XdldhFVG2Cyk659aTqQdTP9SsD5BrhNeO6BcC0ZT1Bw5mIabI4RiS94
gBqe8c70mavwwaM8v1ZwbrWHWLwdPqLErZUU8Hc1QHNdDNlY/0T/2+8VyAI3TKB1RhT3+fnZL1gD
E0JvoHlcLc/A5V7MwXPM+vWartFPbh34U70/KCd6ibNrCZE7xI08NBllacoeV5jyGdTDj1mRZL52
LKIuYDxw2EYSUqTUTxkQcBxdvJlTQTsNnysDS4+WvQK84POwaO97r88DTzgE1XYsX1guiSf4LD3e
yNDKqJj+VT6zvN3AVVG7lPUdMauFmQxzJ/iI/geWp3FoWdzla9Sx15r2bycDxbv0/3L2O5jlWble
QR/1E8iNZmwUUHhzICNpvr5QXp9RWbmJRV/JzJ9zAUU40o7XoXWjdSXSWr6sHWKkZFOUhP/3zXPw
yJZk49sGI8h8YJrWSYeEzrM3+33KyREoqsXUShk7S8RRf5AKZo2IqizZ7T040iE3elRqmuy8a8ip
FiMNiAatKYhYeWZlmJUkhDfnb8VDFzXA/DtM+R+99x7pGL9Klk+JxHyLmNWfosyIjnb3hd9h4Pkv
JtEnVVNR7IAPKGQI+Qy5RrhQGJMe3Sd5IJ9ATEwcbU19WlGcVeF52rxmmZ6sSL86C+PEYNcIi8OV
MzDsunkqkB15iW4G4hgxEALha0V/gPYWDQaujC7hRnBzD0r8bpQ7dCvp74URWF6XY0sY5cPcAUKR
kyRDXggrgiGV3z2mQHj+gdF9iqqBEjyCiprgs8EIojZr5egL6Or+Q2LfLphCX/FoSGTiCRZHkHtW
yAPQYToQOjohqtMGYH9XgfctEk+QroGIxqhsEVIuw0DFDUS1Xe2B+BcFBg5s6aC8C+ECeg8p9nLN
z+0kaRsBdoJJeJnMmfoGe8XSPWZ/f9H2vWQQQnlapeiFKzlhIOvrVcZ1xe0+7xk63dqmR9zYqUzF
MXTFWWpx/XmTnw17Tu2ikc4XMkqGyX6lGAEPoj7FvWyyzahyuBEG92fkyK8/CjIxZ9bOTK5aWzaV
FKh9/QGZqUj5ijiiQ6je6eZ+L2SWVWgepNk/IcmD0x3cr1Qi187LPSIdLsezWC420UfBuBf5AIlR
+iCITuhp8TVXr+uHVcqG4lwmapfIMFpXnSXCaQ5kPmtyI6AbtT/qA7wUbMxUvydhZh6R4I28SwBT
/WIrDNq/LX2uDU5KY6oFRK0iigycAHt4zpgGt/CJwOEqbnO9TPoloF9PXNBsoP5DVsjBwjlVE4aE
3zGyryscN0CwHELZRh9WVlW79h9ezL6JBJIZruTRcMWNP7B+NDYCj+xeqzw5UpPtZvrMeCJZNSTn
A8e4dyz6hGmdEei97gDzGvNZ3AIIMKrGRYdCajasSUYJOvIIhWVjc6+lES/TP1maKGzWIhSnD/ZQ
gwijYl2shRSvnyWMCW5lV3IjQ1LmW2y4rpLiNvByrSXwyzHLseJm7Om5ciBA20Ms7zk+WGQ2N2HL
+q5NtR21iI73yKCecfIk8Z89myATTgzSrlXydowfiF8t0HE/A0HUInh1SShy97nt8iFD7nmZxlur
yy9bjzXPZIt0WwHfItignUAeRCiNVja1NdbP9w0gjC08XI/HQ2+FjiKB8sNy+XIxb74qRwXWp9wO
j035jsamZdRfe4kEcMLv6zVUQf1kwbNoKmQPc5470NVz8HMmbJm+N2Mw6KdS5/BxNNrOw5zLfMTm
EcctCvnghhfA2JVMbNfn1DMGFr6+kWdJIDGk2026h0pednJvXmI5sM4Xv/m0lmXh0ZHp+kHGR/FX
HhAyST4Xe84R5hhS6/+50mnS8Dmy+PCmcS3WMqrNEdKkgl7gev4UfPp3vDgN9vvDbW6FFTzGlmWJ
NM23LO349ELnuvK43vB/Qp7NQTh06tIiNoNh3oLMzSuVxtWz1iS6TFaaluYN5jszGajsjn7t7I0c
BxA57w/UUdhxvDTmCeIr6iZcz4jWgLF5DtfVCCWdI9Csw95Ou7WVgw5j5Gc+IvvAEotrQeMdlQFm
5UpgKBCmTwTwxe19lg3aoSDG11X/kkPa0gpZulf5OdWUccC2cD3fkpA5GHXg3ga+aCsBluqeJBQt
ltUH7/uYbc6kRPxxQX8E6jTD6HWqhZ3AqriuLfGPLVr+75SI25DZ9pAU6mnu5AaB/N6oyayAONdO
heBjYMXKZNw7Dv52genlvQxL8+MArCPRwqFlI4AWKny93DuuMgDQAOiEe23D6JUYlXVGYqHD3yrP
QIsU9rndVOyHN3Kp2nmmRrptyPF2yxASKLPq6JCFbDk/5/TWUCAFmBETTPZl3DSnA9sVWgwT3xfR
gIJZjnQYbUnNhpDLYVNCXr/U7jj45Yl9DbAjbetvzRh8MDYjgM2mepqBkV0zKitddR3CFVfi4z86
pE8Fy9QkEq4pDDoCzY3D755DaAnzy2J4cxPrgPjoFY/2I/+13cJS9FAr673CNTyCvcUl5kifmsKi
O7/PQls+zOa6Qcr74AwjuBUnGj2ydO8OFwKsz6vOSMFW1demuZAo7FzwNeUfp49c1X92fy9YT0wo
TVkB2f/oNMoXu9YS9ZaxMI5frAIoKixMXtWTU3kw//7HyRpYYAP13AJMPz+3IZuVjDdoh1rkqA0+
TuhJMowIiXlF1jvkqaY2YXczdYYCImQucVofV+Xon4T+m897MCTKtNxoZnSHb55StXbDpSQmFrp1
fD1d8zf4Lun+8GMe8n3V/3z/9hJD7uMh89Dz3kXEChD3IItZZkAqaOLetyHWdQAhhRmk9bAxs4a+
7kQzy+ViiP5NwxDjQ5MQBt57u2eTcdCQH+oO7/cK/BXRI1knfZpAkS5YBk//aXJvssEI+G8d25Oi
8nGFn7r0Xa+dSjlGnbc6KUQFfcVYhHZfSjsMzN6d+Yw3jQ/cBr4kpDpfajxVXajxCpkFsK0p/Q6q
mToG20ouFEnKnKlsw/QK3cT77ZF3iPFu8CrfO7LcvTVPQg7E2YjcY19lE1tDOrVxKMISFD7QChdv
gnCcAgkiKbWToeXBJYn629j/GDMB/WFXfCUmOivERoougeRPqDKppqiIZbNGxVPqReOmNKjKkOCf
8/DIcqf0Jbe+651dSWXz01dKrVMEtbmFSQwZt5qukgnpYGPpO0iVBMO0Ww94XlORPi5j7ULg151t
bSWkwomE/FSiBRvXu/N/22bZ1wkyjgYA/he/RVtFoMy4esYZzmgOAmAEtOuQCypupZ9nMb2pWDWT
kmNVoEue03q1Z59ccnZPuJXr9N4lGH1FXa3BSA3IIAS1uW9wrNNmqY5+NwMvCOopTLN6wQzBSJZm
RWURPRbMn3CMMr5LUQSR7nnQ1G3RZQ+7DVf3r7NMQ5eKoq9zOMaKvhN3AbxhtTZg6tIbXs55RXmy
H47FxPuDG22UVo5wY3pxYbX2MQKorF1cL2ZBlkkxfXBQ+lQgL95UarLk+GE5IoU1kzpq3UIW8FM0
2fZWatzA6RmHi+9k2c4KfWH5m+e5qhmt7L8LR1vVAMC8CvZTHAX0bEQPj0gKDzbmXOVpCMEbVyQc
dnFPaCyyCo16LFYlo8VVx5M2atYPtKnu59Ot/u3bOBAfEdTnsEt0gRPxmI8+amcyMZi3038hYN8/
L0pTkQ9nEs2E+mJu1PQy48WaWjF5BHbovL4NrDWJupelqNDqCcWeW+TyBZ9LDDA/UmeWNJ8FAHuP
5izqlFZ4uptIsn4HO4k4eXVOQ46cIYCeO5OV93AA1trPD7jLfHsgOCBO3oGeRn+zA4hyXPN6CnhQ
yjbQdNb9k5K6XFRePp1Y4u1p5mrCT6PaPlO2AgG+lfS3a6rCTPzymKyaQVNM29ZFKQTITRZ7GMdC
kbC56PkLTkXj4kQGNrlUAK+UDyZ2n0UgkPTwPZ0GBlQirrZPz39iIuudlcilbWOzcCiULL2XSewC
eSjmZKa3pg8GbsOzriY9Mk4OJAM5pl8WvjZkfPnfhcweCW1XxHMaYH284ZHPzuPpVHiCTgLEdthK
v8jP64gRDrHBewEiJv0tFlcXOj1J/D7pVr9iOUpyZeWMCASMbIxmHcREK+B3ggH39t+UGEfgEL0x
vCjn1N0lKXeudPdFVQZ84npwNU8enHnCMNRMo55nueMHq32GF1zy5YRP0W1LmU37uYF6/u9P3+76
9PHq3IVDbHPXvbWBWxeZBydaEedhIeUdZeFX/QBXSiuNpYcmZS6xbOVl4s595VTL5SshLyI7apwn
ehvcgPYMW8rbdCwNBJuyLQ7lu5Yy7nHnyMgfz9F6Yp5iBr1weA1edpt809g64krW5kuroFyJvXv6
NAlulYOqh00xwMTBuTURdbi0MjA/RgGrauJTeLctTwVFvn3pUTVkQfAkOmOAu6tm5s4QGLQhNMs3
/OhPqES0B9mGOKcIQimmDmNCMXMixaW+7vBBU0vhdVUpnB7MyoYBw+WEPb9WI4N5tId2mrPTRwIE
iUlSFjnPw7E/qhXRJ3ZIkZMBvAWCKPnzoTV/VLEWHMmqDR44ouh0jd9lSCQK3+PvAyDh49bmxH52
asb6S395XtNv9hsbFNcnqNqww0QNKik7npKeSREoDdYzhQXM9E1w769Mv1w4ptXKULSrvKbOUGcq
OHexmZRtRmHpOeu2XPEH6EpfK+qjmVcoU+fGAQa3Q0e2IVB7Xz3Ih7TpjMHRNSZk0C0mzPK2Mwoc
TvSgB8f0qRFMBcs7iqchRVBI+/sVmL+7j60yYovjr/PH7J8OLi8AHybMpaD58o3avE4oNa2DO98B
4iLaOExDhnVG9/T08jqj2RsQxIptiWor6c52eDgMRP3YxLIhfQ3DOPNCFRE7B+TsW313Ocfwt6YF
Gdq6csbKQ80OAQvGJtHBvoqTt9EvGaOPHcb72CxVC0QO00Q6CvGdxlbumrXZKbfPTD7P/yKHApMw
NMVmmqYtMi8D5ynaj+EkhjArye/cgFYdJTt1Vn4dttmYNjta5ufW7Tj2NfL+qczmd/KT4flyt87v
Uar3TkqVwgxgiwoJi3fXbslTlcF2eGdyq/ZtHIXIiuz7jnpP0sHoKZ4MTxyJTJKh8U36lCpgPWTe
NFRaVEEW5vYrXz/hx0buRr3XxUr+Br9bp9402JWVJ9kriJnEptNV0TfAavfmlNrKfExfVmS3aMvS
7T0zQkhvV4guaaAvTSIgRxGV4PTOidDXOXrzJ6g1G0gfK7m2wtTSVunN7viXbhnOchFePZR01cgW
HAj3dwx/G9uACXQ7yL3iBNYpCxDIUpmKxF3AFzOXofWqhwckzIRAJN2UpqCinXLCm26sB3wfZcc1
UoU9J+aYQY5p3vvxy7vCalQ9WTsZpPCHd9Re6m/Gq7lEj6UgmTuY6FlkiIfuL+g4/ui/h91ZWLF+
4O7gF8tdRFMgmrxf2x7ZnksUmuKjSRqSlPofc9fb5RI29s/1tNJWfwPBCqDKEyG+0+AZQsV1U+3R
vvmVWSxvMjxf3/GSoI4HLKq0D2Uh5OnJj9dPkUogeTDQoFVS7pRhwkDRwQCTXmwwcG7NaO57LbUj
wqc52KQxWMyPsDiPWEF0xZWuJlGRszDF76XOJaNtKwEoI18CxAIHwJOYvORYSPV1GBKdWp1iKmLP
FEvS85mjVAkAOG1myKhJ82Dzy3r7PgbtJsgeJT065yhvWxpuiE73fs1bobTenwIxa8WLdEAQv26z
dD81F4EmPBS5/g4dzRg+1b9RmrmfkC/7+nI5mH3uabDgf3Uo+aImHNndZzbp590p9Abxpi3zLYdm
y0Lojc2lYWpvZ2Y7CSSlSwmY2rGQzTvwUlagVCYE9m3RqtIBib6CukhvYvRwk4R7sOu3hLJzdDyB
nEA6GHHcJIuS3XSYfTY29L6TQdYu1AvgqtQ/6Imxvi0iPCq08owxp50rYXo92tGCseEKLl41cIg3
tnBL62neAogE5XPKGKRlFLrcIK+1TeUi+kqW2Fsk3jmndl6tmKgNvmTixyevkWH41AcGGBB/6dhD
3K69NQuEyYLxBsbN1YmS0qh67SnlW0kkj8hOhMK2eqX6ha/5pomVxqPvFSlTbmV6mf+tgdzaoos3
1fpzZFYaQPqwbPHiP2O/3ZklYFtFZ9ER9d3Y3+JYF/G5G4NVPaxd1oZw+hIxbQDO8mxAN6DRXjz5
VdHsL5J8LJbB3ittScjFra1+KULZS8/iU0FoNRmAE46+Dkii9nuFgvTKRbvYymmaJBR4Rkr3WdFW
UQ3sTTK+8Oy4lC9udUeGC95ovLF4aSZxOOiZ+feGBLis7VrK1gQ19IGhz/UBhEhPf9j1NZp/b5XP
ojtw+Cq2lbeZEICXXZizWR8adSy4Jyas66AcVo9GXHaFwB0DQAAdPbJ8j61Zypj2MzlIoj129dQN
mbnR7HeN2E6/D8vgv8M8UkkS52QBQS+N/y+e0zYOosTjRpMMafdd2oVZ7iwcNNABkglT3SyXj1xj
EQHMbfUDk2SwDJx+f3DsC9aH5Yhqw8TTU27L0HEbP9oM+sJm/0dF5yMiJ1ZvoPeagru3U9Ooy5J8
p7C+G8I7VnuF7MJL6gXm5Lr4rVp11i/83h28CqL1y03V0UwWcBli1sdmmg/LUnLb3ROIgE6WQt5w
vUATPHUwj9/soz53YYTnZ+0BwTtzwvbnBwTjwbOR40VfKuTvhk2/JeYwlT1BdA6Iw/IISw1il5Kl
OPesJEKfII+LMLJu5xbacDEoiqzXGM/2wU5hl+SDXXHXy3u3Ni9smbHJSgGD0iYvTo2RxlxXHmM8
5tIYdbtvfp2p9BV3Vr2GnpDo7PwMwlRG9Ks4nvx89xRb2pBfXiq5qB1iG6W4TGPDzEy99BqUwwy7
shjfZz59qa+b1/4EqsepoFlhqlIAXI5WCqNz2o4yTmGwxdbcZBjQkomS/sFVmwo7muCZypwFtQsy
ZcncQRvRvbhGdVar9TxesKLRaN6Qoazcgw+JPgE5dze8zrxajpX1fYmh5YQk+3l+7NvydVfLDj6/
WnyA+vc7PhNX/OVBqNPo8IaJDsjcCR9OABoMKrxG6cE5IN/rjUKsi5zkoLCSaJA8zMEqTz1CmvJR
MNenKjBY0VGpfN/moD1+2YIu9c29RGjnVzKOzB8UHStHKKf5k8Nk4lLfv9Ksr9ELDZrLa+qecsIL
oipCf9lfWUXn1X3bKIIU0SiTyYyMMskKfWRZxXf7DzjsIlOoVL9YPa+0g9WlX9B0fu11lvZklE1W
uumJ1YYMpk6PDbSteAhW+azg+PeA4i8xzb+yeafc2vysG2gBrPJKQ2cSgKW2ThFunY6ipdHOkkzL
QxLnrqUorFNUCeI32U9F6GrhPrB31E1DOVsiy1X1LqpwJCqS7qMwFPt1zFKMsoU4ezz2838A+4ut
af7Ttn0qV8+d6CkYYfXU5921JPkKP9TEXNv4w6rF4GlaMQ7u1VHi+NzRy9t/B92jWmT8aRg9PDcs
hnrehqpNEDAwM4WmKHxy/op4GBasb1FGiX64fCVCPA84UFXBvh1WFZOMf/cB8kPZfUnbSsAplN4A
zOp3/zvovVxGlQG2KxJpvutqdGdG/4gFLMBLaRAAN8e6yntSELvVkqzWafTbtPMMObAK7tjtBNbr
g5XyXqbqSOjKsv6d1CWR4wL25SHktYrnYTIOlFPVYE0H1+AkXmyt71ppUx9uQuqgzImZCAo7jaBI
/idXqfyUzPazXJqXepXctSoTKsO0uTJrVBD3p5guZBxu5KaO75RIQvI44/rKOy9LukS10PZ3AAbB
aKuHA/06dITSuV9DK5LnDi+YVbvKGfWwlZXZSqvkgy9Xjh8y9jVpB/HQ//8PzYE+o5WiRiTJXuB8
VoAfpzSjzG5YUb5dmFl/KhcSoACd9UbyldMMplLERx6BJTGj+oSujXBCcp0GzhgCXH5aoFCGkqkx
EMZib94Se3OW3yN76ZZrzFq9ViU9QoIJxyz1CRxh9+gtaAM4Olckk+j5Wp4jYEVnTBSZUSudA0T9
ldluhKBjB7bJfDzA7wiNTYjdUk82nIoqMCTnrKGvNFLspTOBt7fzE9sj/wHtUITJW9Z9saWyp007
JHHJIN5Kb+1F7z4jLp8AurJK+qCJt3LXzP7wXwvBQWlO8Ut9EI7782Ontlr6hIt2oDKUwRMhNJNk
gmbwRjYdO4Ca+nok3BYZ8HQQn9bZP9raKMnD7UcfPrtDGywE2qemRwHJIs+6ejXfP0pgv0ScM/eX
hwQLjcxJ3MKfIHtCROV5mQ9GwLovFC10CkfQI2TRza07IQSR1IdlodZZVop7RqNLJlq9hnWzbRJw
anZ/LrfbMBpMe+qAWvKSS9vXhLhg/EK0/A7GEam9HITdfsQ87+syneDnC1jUZDMKageoDhyiuSLj
GVJn/91BgRu4UuH/O9eRDl8KtLHwzwEE0rttEOolcwzYANWFXgei5mcgN4JdOKw/AfTw/HiE+8il
rDnNbgMa21st6X0wBQZZyz1ggdS283DcoEAvx4sAtpFdndClaKuQVRv7fPX5ynd3X3rqqQDsZ/R6
OprcYs0zEZPlqbMfwrfsAi510lEV6ZE3fvyqKsjyvHKh6g28wK7Yi2EfjSPXKvN1A9NQQpmCcwJ8
OeK2Xi9K3gipbl/SdCTBmiGIQ3kUYJrOKsg4VCrPnYhierODXgdHnZsQwBtw/EX6ztdqus6Q3hLf
laeKGshfpnWGDpOHaWsbTgWWgxp0xJgfsRXus61MR2duGw/TGqfSjJG8Pn/EPP/CHjMCKXNL7B7U
AzM3Hi2GV8QT8Cx/pQ6OepDrMH5Yd62w9r60BBEbPSBkST5LUsPQQM3ThmaLFp7RWP03g94fP+w/
trKaFPHfsaLUYe+EFhgDUm0NNxDy0hJKQQTUF5xw7duBaEmId0VdNAOEAQsJu/96uoih/V9cTtTL
1RSOdDYLT5JkeTaDdKOjY9OjPnfrHVzSC8bXGAB1atIL8Be+KmPkKlqBWKwt7SVP1QY4RXLNsQMO
NNi7TAzMuX7cBba491ozeNftTQp8VhzuuDByHlq5huwh3920HkVjY+E4M0DHdF4n4dfqP3qUSGo6
qU92C1jMNELj4UorKrGQe2GdW3Ol109F8MfpNcMfGIqWKaF0UEt/7pJN9HzAxhv33o+gqmfYLRF8
HwMvHD5MPgT0HFWp4FnXAycBTpYFxipTw/YR1C+y1QxJiimZ2Q5FeQx6RFq61mcds3SDTX2uCT6l
PCovY9Uk936qSCkbghiiWo2Ar0MBdtQBOpQAvIuwBwClw1kwcaJzbP4y82QIRm1CjYHA9SNn1cbp
nV2CTdP5BrUYW539m6VLglaMIuQnR8TtYECkfFBikD5mwxI7VUOzu/EeUoi/15GwEkLVfMyij5Gg
G4jwuYyzO69iFbbg4mgMak18mTdz+CWwh7//QG5U38AUTr5Pg4X+ax6qeJr8Irrna/mHQWa9WRZu
I//TIOAq/HUtXh8l4NHNsU8zmhkXbu+ksQYRVdFVcdIbstACA4mFXoWt+7s3IbojyTJYMwOsFAXQ
aXYuZCX9icjdCl9VwmE7jpV9/DxNFKjqIDadgYr6AZh9CHEXwx/bpciwo39gSB6spNayPro6iInf
c+p8Z1NY1NsR01U9k6jacgqPgrNugYsR4FFF1ctpFCutd0HIfD7ZlX3byYyq8vviKEcQcNtjLH/o
GyIQ/ClyliCiQwPfqx2/bKCyi+ozWiz0rIW6mzdyPUWX+d8zpmuErIhtZV0+r8Bb4fCgrwAQ/mKy
3Gh4TuGc8qMZCexHKZZ77LVvXbjSjWP3EPAVuNdNpkO8Q8XBQ+I58ui+Zmj6KeeFBU5867yjH+iE
FvcdL+U+kLekgnzLeS8Ryfju3w2ae6WvWKXPm2eL2TjH7Sfn2c5z1Yuy87QL7FHY/uNy2bc39vs4
AbG6XIGSVtbyk4ujtlvDOBZCfkD1n3NeWSMPmBVnck2sZiC+MI3e6NaTswQT/ULbx9n4LOuT4TUZ
kV/M8jY8GXrt9uARUq6ls9ROmHix7TuoKfwnpnAWmW1Ahkhc5px/Nt95wkuR4nyWCFwE4tXDqcK4
5LfgSi40jupbgcAw9uckEl6gHfFVnqtjpUnEsGQ1s955/QBNMk4QD6vbjB7MQUgclnxekXxXTgfG
07JBbYDAoCgvAM7G3xJxv8I6pkwsxUrGzgiHv4b71f6D3rMydbVDD0AIIXgbGMW609BidtVsqILi
iAWpFWgBM0f1+HtGbKBAXCIV5tihw+e5QxPl765a8hzI9XAA4+4RSJOsXORZ0X227jBagijLRcic
k658vKy2abKckRt9OcAtKyy2XOYEl9HH1UygFj7HnY/i7hxDhtQYShuw19+mvnFdwb1mZdfZjcRY
Ge6xZ3YXTpRfOsl60Vz2WJGkg6NIL36ksOtl8ivFsj0z8bUR8GwGiTKVWPGMvqxXwGaxWoVGdg8S
eRPtZCLLIxJKazVSaXPPsXUUTvsO220vXs5+IAt1kcA2A7dfmEVS3+stY3xDqh7DHkCJB84SVpLr
M/KrVZ3xCeWdu8iWghaC4QbyvJsfMKvSwWQUUlhCaSqkpSM2TBwMqmPdMy9RFT0L+IyO+J1C2JXB
SxlIwkAXdJHN2pESl8PKSRcQy69oFr6fgSL0nfY49UIC1QgbOQ/Xq34+rDzSPfXy5yNLKZAmR/KU
lwWHUpV4oL9bdIc3IvtMM6wSin/KMAJDiZ2vyCuGVYvQvwhG3MsUqwyyTo6QxC3KF85wu0aSd4tL
D0RKeJFGvEjz3LeErjy+Q7N6mH7ST+s6YYpQkq4iXLKI7yOdjdCzXGeydO6lTfr9qcyby0mIZyjA
AG0vj46+zZiWcXXZBI57TxJjReqwXks8E4CVrTHZ7bL/1Wq7VnF45GLXU6WPVN8eFa+XZn5L34gM
bD0C020ZtIItVsAtSi2mgHzNzp3A7J7OcqKLqNZwkXqPXBRkE1M75n6/W+AwmqZVR9jc9VDg3iuE
h/o7kJwJWeQiT4wlDhUqkdqGHk1GZ8QYWCyRnqqQgHqCe+wuJ57gbRCgDioFEzmwnES7/UwaF/zy
Y59mIqdxjragHqvoMkEX1sx8yMN5H1VFHcMvYMbd8TZ0OXx27D+IQq/fESRw30o9bsB42RRQbbAj
mVkWk2uyfUhqMu4J7dUqjaUgS32umg5dOPEAvjlM1H8JxqfBh4w8YvqOJZgWvMGT99X6WpEdcR6j
lGlEba4zzMNnZ40bC+vV3Fwb0f+4RHPD9Jw3OYj7b52GJxpQkyqEpD7GuyydaVw4vG4ZHs4qOrV5
Sk13BJGiQjoqZx6hL4ksJUPHnb/w/BdsW9Q5JSm7tj+r6CqvfdRoTwEz7mmlAqEZinQ5sNjgSXuk
I/vPw5gZcSy+cEeUkSe0awrqpQlXKRA4VZeQbNk3ONzXvQRxaCRt2QAIukUVLMLzxop/DFtzwwZf
CVKpcsbLTq6BEpyto5EeSK6TF6FOc01MKSYJ2nDTdBHG5MM6gt7ARkG705IPDGZ7vmRFS85y7VeV
dtBnyFqBlAWnP9Tw47dZOZRV6CCcalWRpMk0GZYb3vU9po2MjUMweLGQSvsmlCjZhDeYgTlCTNzM
wtd/qS7edx/q/p0PthQVk8j/ggwdAuwUvYBKlUaq1AwG0rBY8965u1oUpsyfSUhCOK6klEyoW9KJ
fmQDk9dmWEJojNxUmPqfTr2mqetS/DmjC1UzrgI4wIJjX+f+kLOCqwoa+lVb0qumGrNpfU8Z84aA
ikX/kddrbqMjMjvd7YMASvf866mKgAyX2JOPNsczWg1Nx5bOe5rP9Wbw/J62ng3fbw5dWpOCUgrq
oNDIFnNbJCccp2nWvyB/yyNS5gPeBWXzxvl7RbgSgmPoyj1MOSgJ5xXwuXEDgqSzodBEygzZCbTw
jVInFri0fpNCoqPWQTvvYHqzd/1jv8PSNxZZvhf9aCvgVwKhHfcP/DCNRUWCetkULGTbUwd5eZSE
MqgYZcqGC6PogvnplCrWDImLKSJBKmIVqf82FEQw+1mZEjxxjqKrlh+LWDABw4dWIV/ALBJmjbjP
d0ECKTwgQmOEhkb+JAMolZ7407AedhDpJKvN7XdZ1FdYzYzPJ7/y/dONQd1XigBHXHJs5iTnYxUX
dt9yOhhENvmDwwnP455bBiKcCfnxTuk7tauuwp4d4+7RzvEq1XhebKfk+lLhX0RcOb7O8NQggJV4
QKF8xbAUW00MU694ZBPFezBBQ6caLxea1RzCKTAaMyWHCBne380jfXl3VSYMt0ZCuWxo8unkWet6
HfawMaKop0rUgjlOiy1FrfStquIhHWYGJcl5/O8AdlYNphe6qm7agywGruajQiDbHMEC4bi2yM0J
/bUhRbm5/64jJjzPvoLnrKdG3/HY34BivGKtAAg0zFYxdKi0P4nYqAaNvIy1Xvg9Q4ROSinpHxeK
zU+8102BIjRgC9avKuVB7CsbawwLrs4XASKOm+DHftrmkWZFWYEIfP8EjqLDQDGPl8VP2IFaPbJp
s0PjHwhKzgNhr0u8r5TkOfG2v37jKkYHKKO8BiBIE6vYTEyqsF2rlDYgotDX2DJjyD1AKasHsweP
Ha+dd69q0cnSJ4pZsSHRqQKRwq9iuRcBA/GgX/0wsKLqkLVImwSRFqnQ6YcXRhC8sm11Il6eyTa9
xiysKuiSJk7ulN6NqIsGWlCCDgsRqu2bi42jYOAnFINBcL8kFXUdkgpSkmwAsvj1CjdYwBCZzetE
ybXRG9bE8NiOjX/IUpx/ll62+dsm954PWwTPrQPo7cVQ2Vef/B06it/JUL0fQer1GkU7yV/qI29a
537y+qzQZ1t8mFzbpwq/71QZHh+TJcjboJiDIfDUhc+7RENjMatUOS1Tp6TDuP3zTNd0PL1BmrpP
+3Rk9EfycmvMzwGjTPR404Xz+CM+DqrnRBuftbIXmi4KBXvSiLqnP4Gc01H//jnBHCjGBSGetPc4
RQ9h3hyAblR5+ea/VY565Z24Yn9HERb10eFe1cs90Pw9x0rXtzjPRp9MDokUuejyZnkFtn2gSm6U
h5gs8AooSUdSuGY0GNoRbMWd8O82bGQeuUlzrjtNsitOdVeWUkaxhka6mtOeTn1kwQxNVTSC367X
FZ/tADKlkLCxH78go2u1daj1Ymd6kXgocHe6dEjOhW1bA62O8J3UeogPArQ3jS6ZpKIdn7Qg1PNV
w9AqGnCm4OqJ73LX8Yc6K2zZtkAuZ9hbxfNVYTJ70A+ncZJWqdC4cJZsIbotMCmdjd5R8vI61vVa
mLIe0zRoM2wNBNZ7BP4qOD6zreoajkD0Au9pOSAmTlVkZkZ9ki4l5JOeBD4/rq4AQRjXHc5Pj1YP
q82zWYnOQsCJ3UrlfSGul0lhVbJ/FqbtNKuuN75R6xIoAew++hD25JV2stWhV1aHWMBNl0sGnbtO
wRnYeTEjvt4JvFtC2mFe+r1spfbjwLavg/zF3Kex7RAqQYsHhRxD34e9Pm7l2t/s3L0Pz5oQeq/H
5noDIdmXM6eQ0gbq2YyvBQiRCG2SwnmpBbqUB/ZqrD0qgv8LDqCLk2cIacDsSOgdc13qwMuz+eOt
KOX4xWoG678wLB0S1O6tPxuwVMsYO5huj4GqROq2qh3Da1Gq+fYtgdqrPdRNBf39Dv0GFeMIyaU0
FYuPYh22eaTjzLQwDI80pq26G9YuzjfyxW99NjDMfQ+GJvRhEGLJLrq3IbrZCH2OMHHRqNliU1zQ
G9y170017295Op15hYCg+HX3kzu33qBc/sstHoe8xRxhEV6JH4j8NGRG9h61v0EbuoYpCn6W5VBp
UO1cP71gjF/1/U8pb4jz7CXHEkrXpqUMy6E2sP04m+L3oLUnmN45f2fX/3nwKFTHUOrCkr1QQIuG
Y/wGWLxU3+Pd3X1XMyoqwJyXJgos0RqB9FV1yprWNNpBEzRJ/weB/HlTRL8OHptC0VIYNXk0luA8
hSiU1uk69cX8aa1qK5DGyUpbOfXn6lTGKpM0qaAO39MhHHVXc8ZCW5FMXEHm87wo9T5ptUeByVTr
lluoWpKZIsnuMYZcjoHSfqsJZ097tcVKEVfjNRqsgWz53TkRSL0/d/xB2M5o4qlB9UNzo3QFUOXT
kRCtFjMcau0BUBRhPx4wZ33GVd+Si7RFkbbc22n/cELtz0Q6aghBbLlbL/F1TzhikpPjBojB2ipG
kqO7cswta3pdU4DB3M+nhkBtOXTu8mIQUsRrnp++AZFcRuVjX2r973y3/dMfRZ0m5ZsB2xYdgOqY
CIxC4rpgm1oWLlUvWUlayWaOr9GjDv/9lsyXEufhmNg/EWzUqzwyB/f1yC/rkNPaIkQcSigh1m7W
o4QtqA9tBesP4O4+C3D8rEfP3EM0T0VzdYw6DU7fjK7VSOp2xQ6pKtBbVcUujBoB44f83pcbqHle
gjsW8pQi4HovisNDPU0tkOudf/T1HB5vyolK3mPGvC8idNJCSe5iFkbFQrst8e38sobLRa5rwt0w
z0juPdyIFN++9LrG9dEW+DYPVUx5xh9h2o2alcwWPTF6etHDkAdnVet8yDk3viwfjA7vSSClrkHD
rGOF6+1Lb6CEBpXNyHOL9FTPOQa+9/S2nCoMd28GLAqr3aB0M8r4oV5Eg3TM8IYu3re+shnSC8VV
GYB/grdokdcReIm3Wi9KAuFJs1cQSWZbuYMoRcFWLDBEoINtnmma7/FfuOEXx+u4K4qtoyoECX9J
4FOoT7hWfCqBS8uKXiH5Pw9i7bNeQqEqvNl1HhY/i1tj1ndBkQqEHipsvTfha+rPa3GTPCjc7AzN
gWjr6srBr+dftW/bQtAysMCEFyDmfjXvCI6ftvWvpRUb1EHqYjJvbKoXbZekKrSMiA4DFdBwUjdb
WwrrB9kZGmrhnw2O785Kp4QpMA3cmvwdvR5Bv7HahVimPmm7gzO9UDJNy8gq6wbNfcvrxSqKDlmJ
MPMVkPbIl8inau+JMQcKP9XJb1GKaemz0JcJNVuGDxktJvcaFhAVaboZoJhB78SPeYt8IMKlgw5N
RbBWF6sPjnutJV6BX1Z1nWesqR5uaK1laHZg8agNYNYl01ZaSG4Zy6322tYef6zTlD23jd0lzkBD
Rl3TawY93NoE8JpdcdtUStegX2RTiRBlAZZv2ISrucBVYu9yHyCzPZZc80L41UQEGaL+6UuzLKEg
AIQdjrs4h4nZaKoXH59pEy+ke2Bt8FyIjZugI2PQvf7G3XdAgm+wSZcaCDfZHmnjn4/2QpijnSjB
kTOFLAE6yfx/Od/S5LLph6wsSpbYmNltHsyOsjjALsPE3QcCudktAzLx4JdYkF+ODBqn4Em3YwhW
ikjcKpjD63bL9reeo9XalNKkIpgEsQVt0TWaeG9UMLErBhvvr6F6fsAwCfacZiGg05MV0tvmzlHm
YEofUndWaEgMAH1UXBrMMKPqyWRULLabU+pSwdF919gymkEuSCb5rYmRFJDhBCiT1NHjMUE1vRrm
fu5THLz65AwlIWfoOD4EnbdeQFN/WAFMhwDN2yIiPsv+SuN/1FxoDWdcv8OtjzN1RBpO79dh4Q6I
iLt62CmHwz4p0oPt89bEU70VKrg0trZTuOsggRCh2zmVmJGDOSjDBrzpE8XvGxJlMSb4W4DtSnmI
HvUZJCAfZfAz0tBIznBQzYXXiHLt6c82uXaCWnTuDAZMBKkMZbYeigpgWxjSytEC4dpeyzntmghN
V7O9Y3d7cuy7iYwKQ3cl3MAg5I/uALzr788blM4gVMe+sPt7VArJa+bSK1R6dxHMr9RQ99IGkE/1
XaNV6o2RYU3aIh0g51H72tCVHC+0Jao9HQSHkuN18mMurFZVH0xtmFN5+x+3HKb1gRSGOljqfjuk
TFP+okSKCC1gJigZX8/XxLcv8Rm5iGNcOw9he9Y0tbhOEF4atxXduRXCmiQXVT/mK5J46hIvK1Q4
a7UDGUQLTc4tv9BwwkxZqTiUXj96ae15hQ4tlvyCrcsnOn/bhF+BMS3epucUIWmOrATvKYf3KoUb
Ks2eHnPCn0uWoC/Y1WlQL/AVg5pONfdEPETFKp0lUkCoIoArTznAPAdFu45ilQxuc6UbQSOIpt0C
FsUbb0rto2JPBkDGFWMOPqjr+DTpAcLL023nh4Myxf9zGYSKzlz2LSRITzJKPcZLADjroqG+T0hY
p9A3LKxhy01bEz75ueQ7GK1PQoLotqCcs/U3yT7pWKefpDstIxcDUK8+5+P5Y/5Co+146D5WpHO4
AdwCkA3j57s7mhIt42iBbv9yeb0jwjCRhdquwq5GA7hofA6iPkHDmk2/teEQxzJphU/a6J6uYGoY
1lZTTFil+BTugL/rP0+eumLp7BFoF3JjiRW+k6NxkxlobBRTP7kmX92lTJ3CDdCwqJ9sw07GxdkY
JTUmWJZ3krEciYL3PJlk4XfU6RLvHu/9pMak12r1b5yeXWIeRjVKA9tp9orrstJ8dTMlg0kXaZOU
yMxmDJvtJTL6Lj25c05vEJcRkpyVtjPrKYzPl165G3OWiHO8MUlnAKkZIPCM4NzqOJnJW0lNKO12
eyecEs54tN/WjVNFN1tVQtjxIn/s5FT3QrcIU1MUxLjJ73VMiRKUS2D6pvLykznZTfE5GSfOdrAb
Do0ONt+VyTiRS0UoSZODbQykQ8eY7VPce1Zr/HP7xb2U5ylRrmIVp07tYoOYcVuA4RJPobgFye8D
6LxxAtDuBYd23qWpE33XHpgIr+42M5P0/S47OTx2IWvzHhUxkaa4dBqVtYcYYuPDbomkAqZ5M+4Z
8iZfz+mkUFJi34Wdd6TwD3yluyI+WymPegJX8vsEbQ0s9t4ObH9N5w6lyNCXmUorybqMjwfWnlHh
SgepOX7dTUA8Ewy0bR7GRbysd//RkXFcDazH35vDogNbHhA5eF7+GraCZBw1WzG8Aeb0sxW+r2hB
BzlK1OUpe3W3sujcPAGEu+zE7TrKQTaSOOO1WrAQhyQlkphuWqTjuVU5c5QPMChltOPurS80dJan
S52/CEyjDPgkkdM2RC6m8BQx/sr5GbWyH4fv+VNIgD7si6rwNbNCgpJLWL+xVk8FOhiKrzj7RTC1
98OcgDXvhjkS9XoFDSP3liTasUDONdBOmv7zqDmqEQXgBPWE0pkd2UrQsaaEI2QxIc6tgR2hGXgZ
AAm0Ac4MpV9lrd1kT4XQiVtzn1TBaxOQsjnZYF7+IWrLnKEEjhzqecPPFEIuMjr6m2ap8ajcIfXE
Zrl2QTE0mmDN5t3ILa6pEgH/+WChywR+eKuzCwyz8rkfNYQkcTxr6P5ZvfXF1jBUZdBSUGqolJNH
L+W3+jhrJUMd/04YaswGG+4fimw2V8/RchyUuIcrRnaOpp2kBFsowvF/iHQTCHR/xV6GX33yoBlu
iT6BdXZr3Hb5PRhPDdyliap+ntOWPUMmzcR8cP6YdLoqxGmt6XEiAN3cECSIhhSMx0ha51D5A4VO
c/knbubKsvZtnDGCEclJheE+Iiijjexok0hg6vZJsNQ1GGvT4JGb5XUBG4IAIPM8QLYF622G8dVs
sabSCvN1b/TAfTAKS4tsYzZv8pNxn/PhkKuXo4TlTETqMukg4R20u2pI3pbrElAJumGHSNcevprT
0OzXTyu6KyyQB4UIJEn7dPaEprLfBAJfUrGq7Bx1BsGXUaQoTc4LC84pJeycvGJ1T4O9uJeZN1v3
WFmHTb5arHNJpD8RPpAsQ7qpSNLFEvfHO2jaIiqN0vlIJEQz2qWXnmybO0T0MG9xciuUWC1lCuve
KSuGyADZ9tY6zI06jCQi5tUecH+vX9iv8M7b0YPX/I+o9chbapKly5EBCtt2244hdbg+NB3BNVXB
2ZmPS26KRrhRMHV12HO5fn7hvxmuMHG4ZuLvWTiMnmleLYNH2BFbXzb+8PnA4ZD5xrqE6BtTExXw
9Qi/M/sjzIWBvk918DU0gKv9BWstGPEqo4Z199r9vChLRkrVHv29kvnwwWZLnTzNWj/rp+wJtoHX
NRhRZEjF0WsR4y3jhJZ/FKH+UzBvT5euPOBwpvYfl7TwmtUNCB0kjETwDjvrpUnDrxYg2V8dmYOQ
wiuOif5nCp4RNX9nZ9+l/9dmynaowQN2YDdOrozyrs4ztniIHg4pT0vb5/CVLU5tictiLTvAVXww
z5x9SZda9fimNwQuZAuQ1sBVcOBTu3WW0jAI5EQYhIDFXx2eWketOabiAEhSflhdcdAotuUz2RWS
QTkiLhcZkyCqUbqBFTbCvtmD8DczWmhbhP17b/AC1E+tuZZEb7zim8M5rKY9XvVUxVHF65UUKOBJ
G4lzu6deYXOky3z6PaB3srU8fWstuz/L+B/AbjETTQmeaCTTIpT6VWw1ORpoRw71SobTLofG8h9o
wXQX46/1UR3PlYXqdJFkG4d5+90cN9OaOM9GiFd91aDimHev7Ap6n6+lL8MQzYCJYnHHeeD+X/Iz
AJX2yssBzE98Zf7J/LnEFoqKylB3Jq+d74hc89tYzHJGPBmDl66u6QBVTBBsz6SRD/7VnCnXxSHm
elUr3WfS/FNtuA25E/eJIKDyE5pFXPP3rv7X1C79oHU44KWTTEVpcmJmGS/3pgp3Hn+nFejz6IyZ
mOEXuUYGwkGpqoffRrbe2uoSXsR727gHGXEHcODobvoRR/BrrbRLd4pMWrEKrVhHatwEna+HuMVc
Lesr5QnWxCd17zIUzRzuDCJzNgrP9tFwA8NlLQneY4Y97XMLP5eGQRLexb8lKAXm1IofAiFrg+SR
zuaR7afuOF6wGqopHGtnTh5Nay8YJ8xiq3x/+N4yDFtaPNOe2skZahSTgytu3/0dx19+PZkSCoqb
avFyDkp9UtBvADWD08790vLmtq1qQfPrZOddkofgr8zBdFXBgSLbRSqzzGY8gFimtxGnn+aJo0vv
RYLqW0aSKXPAWNFv6WsPubkQ6gQ0NqD3NvvTE3HyAngLQDivsvEqDTpVp84Ppg2XOocIa3baGt8i
3aU8uT7dGuIfZjR1aYBeWX6vKs8e5joGQmlbgevvkQYlD5grg/H7bPs1oMxA3rVEpOjiIMDOnr+i
xMI/qiVpzuHyZGAA2qK8xp7PMuDf8SBTx8UYchi6wJyz9+MC84mDkYY7kmtPiE7Z3FR3pTxr9Dq3
kZgUMU+RZOK99aZaOh2JH12AOFykxMRPiHnFXCs18LJjH91DIhjgAkWgT60nJJpR77eF284gVWjW
7GrsDctTT6BLU5AXsAOpRUQegHSHO99J/ZZVETVx113/iqg6Qd5CAbh/+StSPnLFZD+8nkn+JXWE
wVoNffvugxVYc8YCWB/kcabimp99+T4EPBVxKIX54HQ4TLWMsMIZsTCiMn1Q/ehbn1mH+UKAxfMk
fbXkwewQJYyQmiqcn9G9w5xuXPMEZWTU4vr3BZ+QCTcYk2V/m4zft8alHiF19pkTxNABGwCQdqFG
3jj/YAtKrlsz0FgdHtHzCgyzYAMf2Hx7lhUAY3O8ciXkQuuCJR+9cGHX5eJ7O4Hi0SOCj+5/vDNJ
+rDozH7NAO2QuZJGkTgBKowhyh+Uz0QgQXfXwN7O1pIi9NRRl35btuSsBvv8ADqEj6Yeol1hHzmG
gWxzjSjriyOdNeRTPh3E7LS/fLsjmZyWsQe3yal9kXy2lFE3kd4MGpWxAgCV8L+1llpRF3kUpWQW
pZKjnkjz3kCfEZ6ca+SXn1a6mQkS457hoj6DgALye+bDTI1aj4K0Du6r8RHugsNV9dw3EPXHNSDh
NdDkXYIjRtQ0+ZPZUfOI7YKTdBr0sCLxRXNAcOh4wWsMruLUanu7MPOIMIAal4alEbOV8ahc3A80
1++Ncy90fqUyzvshwaSh3sEKCPXa1HT1LIZlA4HZc4j2ep9+IWzR8vlh2xqoG3CIsyv8vYF3nvoL
AI8RpLL5iojJqyZEBGwZFRZgFnGkr5Oitn1peT72BaJjn0xiuo2Fhgnz2Ccq8EpNq76uj5hMy402
XoBPaoWZq1FuiVsdE0Vm8UXdPMMveq/Wmznt9GGWURkhJd4C7J+cKyvIQ6bDMqjbAhioVDpYyiHN
dd1b4SypIuYf7GrKSxU/ih/rxMwNUPjdDpAwz4N1tAg8tTMuEOT6mxboKE551z1sbjKH9oA5VHUD
u/RWCBiiHiimXoNMjabNoc4KJ6iM//P3x79SvuYFuK2xAFGUveRPF8gTK1jv01OxwVsg+xhYpMRV
2IB32dt+XOy6tcVQ3fp6xXyb8r1EmPU05799IqUxq/CovKGwDsTUcga5uRy8uYpD4tl3ooVHfsH2
SHJf4X/t6uxNsUxhD7c+T4iL71DvdVXy3RpeNV4eV3J+nosIWi3esDLRJrIt8nTU7sXb5xsxNoED
SpjNJuvwTGa1Lktq3KEaS3r6AQiKcgjDkMMT7o+g2Xi0zrDyB52+1q9W+f0DxszTHEDfoURlXLWe
Vb1jxl6matfN46ievftJ2Y7paaqAMtr+IAc85PpKeI27qyaNdL04+qPWWA/t9NxRe9D3clxndEnU
5AYXvRyxgEowJbsSJVgQtesW24InbViw1LxqpxEi7bWeQybayUzt12/eKa2PhEfkCblpZw6wDDX9
iVmcNl6vzO2P+0+U81s/YiUWIn8uBdHw0Vd9NDRCy0MfCmkNRSoKFvZdifIbIP2/ZU8tF6JaZvEg
iSTv4KT8BPOM3rSS4jM7Ndr7jROnIdBiz/dNiWIMP8ivLV86FiAJfkHLpy38+lIpDMO+K8mZMM6U
ATVPhvD5FfoB5YmIJJao7U+r8Vd3DvNr55gAp7GoH3faNRTZgmeR9yyTlnI0L2VZC918HHId3kpL
BoG93u9+ib+wcdUn5WiWNKX7HbK3TW1AvakeSHvchNkAfh1dTzJ1qz2LOem29v7iwnfrIPV6z1ve
h+qBc/r3vqN4X4N0hIqHTigeDhAGnmHJhh8cydIvQDB+gggruM7YmN0lEwxScdgLrXPZPL8lt8fs
Sd2eJ9olH3SsguYfFxNmQtdZCAU5Ucf1hqFRuCwx5T7B+kEwL1UjQBUcbAwua+3JRAlllAN9FEuG
F2RR6k8YeK/2vTolU6zP0xsF8VXxfi6Eia5MljHbYivBRFk8mGPrsPQObHExU2VSmlJdBwkqpI3m
ReIhjbdcbaMTjBu0dKOpQ+1IGcr5aMU9CSjCaBoI5DIgAi3L/poIHrB7bY8+EjCPrBbeQU+AaO06
mDahUnz6J2YgKMl6ze3FrTomFnvRQtG0XhjdqNzbj1W8ph6ArxMoR6cUtjY68aRjMvjbsNY3TNyS
TaBv/hwCPrOgYpt9U3QgR4rZh/FMcGk3lYkoJyP7p0yzd0RF/L4Iv5R4PM8eZ2UwFD+l6VUTbKkZ
rRKKs+944+jBeP52q1cS0u9F1QxZiunDqiXF3rMDrbmGePynDfSGkDvjA7wYHQq9BCC56jjwcnYX
x+rkSc4AKQgsJZ753DlPQMdPydHBNlAuR+bH0dvJTZZhuLhdnlIgvJfsEbHRhsd/vZ9XVA5+YjXz
iewalGdDd5wIpoWWTq1f8M2uQobHnssyYeh+ITfZqfwUI7Gy8BJ3/ppKQbf8SNXwV2yURWuhRY3J
O9SkPwTH5c2dOxxco+t+yjuea975OAbxL9rJZYHNlWL57Wum+gt6ILbywfWNueZID3DICa2MaMwZ
3G29WRWT4rZ4b57j4WvB2pcemOC4qkc1BegU9ajdWDap4wMTEfeUDEVCNnCwWtVPpD0R7dg385xK
z8CSwZoBpfQgDhGjzGKceyW2X9tKN3+5DwD7OcFIkxWKtkKE9bBg7SKXzkLR9IQFy0L0M9cXq8sJ
o9HWr/cdJdhNx/TJu16IZcfuGJyhNkRucdVxUJABc8w7OO8iLingTk7woLvE9MyolCdyRVNbgvhZ
QmR9JQG4Qk8IWiBuMYj4603Ca3al2OPyd2RcOC4e7v8ETufT6hpnJXNbBWNJC2BQldMlfmXsl7bc
C+9GxA8dSqp80dW760HBVBWYMEh6wO916DdLgZJh5+j8raZUEA/9SiZ2UT/UTV1zBGXHwzVq+/xm
J4PlNZdBD0ahIIa/kjwu30KyQh/+Cu0WDBQnw51CEyfAhqb1CI43wM5IN29zd5lvHFthThmmJZVr
TNXYi/4zb7QkVi7Dc6+86yC2/ZMU9EhJ+GChE/gkyiAhCtPnItvwX/q0kCvK0d438UcuMr1hx395
Ai8jKP7W7ba8EkqluVehQTQCe/WM2GTfpdL5SA6F2fIEaOnGsQ5BDSe0z/L9b+unf5evQGKQGLFc
QH/vWuplMnhQrg8TzCbmgpVFmfofWstrgsb3mYcFrCbxaLYMRBozKBN6NF98kqz6/dKJ6sG7YR4h
9oPYuPOXCcxvmTHSVkkZdKC0oAlUr5Mcr56FZVR7mgZdX06MHdhEGHJHB2miysykUg6IkXGjhYBX
ID5yKeq7mtqRl4d5LEBrVvlFkRnviDPgZ4iaoEiUGi9CISF0+novyurgUpm9y8SCXovJHqN7FMeW
1/T8nHKO+QLb4CTfpNiDzfh74P59GOkIGgyQtiuPjfVwBuCkFeHMNOjvfKSg0/WklUEei8dv9W4z
C5GwTAeFUGmTDuPSQI3bY1UdpgsJu/BVKjyOmH487DFsLGdQdCZ218qY7lSNeXC+W5muLAc+FE20
J5gPPefDc4sQSPGd+h/2iQ9vMsYr3xVY0jWvRqbkteZPgDFlsd/zx9R5CMtlNAkh8shCCzKx3tnk
Z54RTV74/GaAZ3fMWCAaSQl6nZpF4Fbpp2dwguAsxJ7Q+CKcoP1Oi1cWKFX6Pumoot5HwH71Pe1/
RGMCbKfNhkDd/7l02hfYLpsa7r1S33QfQisaia+IOxe3iBOnBOhuuuy/blRcWfqweieAze6uwsSK
Smtihbsptt/5x9sBcqnG13idqEnnPO7YNxM3fLtjocQKPi1l+wEK/LM+UgWzT/i1z6ZvLMPLFPxd
JgM/oUxkDneP6Tf/YzxVI9AXhzLAhVYH07FpsgED0zcnDfzBjYK9nb6QjvE5zVGpvagG71frzMSJ
Tq+ho39TqgGFv9nM5DSZugwuo+IM1zts/YIWbhwmrqjZdpF9AFBnBGkLLOTX1qUYO21ifZ6R88jo
/Vag0+Az5XAfyNyGnFF/coZ8tpL7tj2D0GbAEDyPDQCJGeuRDnDavc2NgVrNrqV4+hdNnKTNMhb4
MzaUMd7n/DR3b1aFYugQbQxtvBGUeg1vHEnxdPKrD0/al8x9Oz9eUlZrm6YnWm2IXdeZDZcKFVu/
tb1Kp0tZd3EG8OSIHdKEl/zp0GhR7/8RehC4F2gKPVwnIaTy66rXh7YC9OrgqFIzI8bjvNfEyJa9
/0Eyh5zqAgQHDB54M8fK+1RLhyYO8DgATTbuyB3JzfFDuZ/TJY9Y+WPGUt9xIXiWW8YWr0PxPQGR
1usewmBn+b7cVooFWDMx8NnRmM6HeJmWy9H2/PJsAD83afOwg7qRcyDhu94SwSumQHhHwJ2araqy
n+CkiEcYW8F61SvrGGSNCqm8cM0vFpTpVKM42gS0jd4GGQ63oul6GkmFuf7Qg2UXQyhtu9FNhpg6
rBWqJkrFEj7CvGHYb8pLvRerwnJeivqW2A+IBUuCO32Bc349tTzk75Pibb6QniST9hpc/W+ZcHz5
CTdlNSpfRq1sj4U/Pg8eqr2zLUdaYZ9imqArlqvX+EFvNUpeObKHQLycmkzL3lXrfAvQdmrWHMYH
niHvBdkITdV2tSQ6IsAR5afKwpljWilq3JVcmIEYEsb6jptVGK6TMNsyVa5o7YJIsXmv1ut9zYY6
n5ic6HEiMTCsIX+Hud1Yk6kRidVItO83SxilFruBHsIsOuwJsssHceccSXrul1vMYD0qsBIhOQov
2YkO1YH48vJ5l1xjFBn3Y1X2cwhHtDfl4s7/WSFvQS/5a+fhejcSAghOBc0/wNOkWdEKsPDqXWxm
90kaq2eYAKGePrSc1VS5NlWf0cp6ReqZ81Gkw7LqROrlxHRNLRT8rrrHMpA+irpWLyavxh4mTlJl
NVPflZgGohS0Uy+VQVF43KczNYHbFgIi9WewUitJxtUalIfiyyBou6RsWhegYCE/Scuo84ugrrR/
FW6NkDLjIkecbAUFEwDCb3K7+Z9l/LRxeytC9yhuH7XBC3bu5dFmEhhUhFMBUNIBsoDrDwwIxK8x
JWmUA22BfE6JjGQbYnOafa91JWO8H7paB6H9VRsLFV3dNTc3TavZ3mxQ/yk/XWxqCCL6mLMO2Zhg
L/HkVWgIt57zHtI2pgaI48QgJ4B/v8Lo5+EDhi6Vr5NhHzUqQ6Qoab+/0TTHFKUPzQAHf27XLyEo
C8LCT09MzlRHG3AKlS4g1GqW/2sqHVCRvlVP3n6yeGQIh8Zr8HB78SvC26ux7SSM1BlHAsfcyRmH
OpvmPVdKSZm7V2aL/KfadbrTqaOc5KhYNg0XZzGG7+FLjVHGGtu8na6AhyBtDW9Q086T+0WjNXil
46sivaq7Eysv5wK7kKvHnc+lhncrG2sxQP790i4F11K4afURqd81KIg/Pp83Q2FOFEvWL2LYwrq6
UUr4wJUVAI8tYkZxIKqtsDY8kRPx6VbwkINqgTuHfSsA11tXGXMnVsRM1B2NhrV3NBtLLoOT6kpr
Q6aGwXvxgEZ+zKLIoRy2S8FOyko8zv4EoHsPKcthEgoxiC3j6O6zEXBY1/jIMOtJGpaQZ9DU1BJD
OUHW0Hm9U6wYMQUkAyi0S5wHtEqqa5F5ptKR3z8XrCKK3yNesrWzdHdAqcRXcqOK2VTZOcj/1Y78
+l97TUWUyj9tlEoxJC3IYe5xbQ7y/5+zh4LSeEJzYrtWQ1mDSuQBn+JyFOAOWkYYbBGiOlfD+k2h
VI3fCu9+OcoXbngbYOnBzxP0Onl/nLvQFuZTxY8XC9vWu/K6JOL6B++78NMZzAZMsyoLtW6UyR9g
XGbRS+wDSE39+GGRqWsDj/a8lIEFThlbuvKeqng1A+yg7Hyn0RN9sKQffS2ftpSwJ9YXtBnidWgQ
BJrEo7HPqJTpvzWUqgXhOhwYRjHPoAgQmlbTgv60prFdV1UapNhChI1YlzUdN7fv/Ns7DrXYdPz3
hy4LQmXjGe46bRBQ+hD5/iRP/L2qFFcb/sX4YvezZzsOMnaSg+jUvmMKP51WlIoArrQycuCI2xJp
E7tmalEUYCvH99b8Psw5Ta9zrOJZgqZspuLnb479EDIUDHY+Jy6rgU350Z5arkTK6kCNafGQxolC
bRrdXl+z+AamC8d49jUouARO1ONt4jvtuxqg5vIqZPDqtmHMCEINYOZeDnAfZlNWxVsska9HV8Yd
7wx/L0DI+Bp0X1QTHQDuuINL/4rWPtisyivnhw8gQbBsEIFmHZNVXUssTZurdzItE/L86+3ar146
NBc7R7zMhI9giQUwbfT60UA8XvAuJbS6fZSGQhP8tyO5TeV2n3vfYzAFKp78i9s2qZpZ0qHdwa8p
FTCWKlKlfOBwus7+ZbqLYCFJ0hiC732UfbhbTXQuQlRH31T4OLL7UxJNrINOXDVHZue1mKMKn19V
scW+QNCkxa1zO1f1cFYMeHpdobodTgepajKkhK8og755n8hv4/eBZj4mmyi4s2SEn3xysO1Qv4iy
0Cf3uksuq+tZF3syBYi1N+lW7O33fgrje5+NRrPb6tnTdKNxWINx0RsnmxS9nPtdJ24Blhktt2UE
WfFCHxlE6qgy5LTmnhicl8II4JSHOiVrGqhZ6zwaLuqPms8zxfdYHDXxGqYhrea65BJdthbEgXTy
mpaL2EhH2prWW5zr0eNM8AyeI+ds5239jwW/ygesJ8GzuO3QDUI7fdO5lUFCYLQv8twG9ThrtyJQ
MPeBBVV+CZFJFI7EbLqfvisoYFMw35E5zFC75uu1e5U+Nb2XnBw8gXhgZ6Y+u3gFQRXZiu1LGLGo
W17ZASAjxyZ6cKpIxoGk7vxSY1Z0uKvEVfTrGQJ2e/IG0OmGAIlX1F9ejW+JpyXfcd/MKjI+/aWG
oyA4M+kTqWkXuUos3n6AxtQKumsTM9iIhLSFtrW/YNuPu6VCpR1WJ7CK/PYmZ/L2mYSqy3QrF3fH
IStbbt18aR5DvfEq8qLT1KpNVIVHfFZd0eCY9t8VrTcHRLt7RdOpuuXqeE1jnpMoaJpA0TkQ46mi
RksgbQC0jI+K4eWJFCQTn87CUe2GXrDeo7//BisA53vLAjC5zkhJYjIaGJoJGLpcAAx37Qm3m9D9
Kibq7aR5G5cKJcaUmBs5i0e+x3zktP+CIpTEmjxHOWwIMXbPrZ0RgyflOYdJap3q0zo9c4F9WEcV
Jy0O4mIfFiEz+nLx4GIRdLvX8xlAD0Yo1niv6Ure2cSz5BJ9ed0VME5sOmbuD+2Uz15um/2D89r9
fr0wkDwIAPE3UcvRoBj04UK7/pDbJH/GA4XAuDZOEOJ9kYyTnBN+QG5i9fKZjS5DMlWBHRPwsbFb
IoXv6Jtv70YQcPV3YA7oVvYnt0enCalWccybThm3oQOkZkA5ecHGQpaa5K5LWS8flKzz11XLY4eQ
SY3OPhu1ecnNa/UsfHeaDftJsMKGJ+H9u5jwDc9vz+eXeEZDACrKiNhotHPkNtspiJt5Zp4laBvj
GRH5opBGOCPlJIvthLbNoo4OSOJmNAksn2rbcqcmAs19kaNrSjWljdgLlyPlVOqfZYnrB7xWW34C
HB8IWI5jfvX9giX+XfjOzgblMhNvCKjtpMpHg4UAo6Lr6ocI63CO1O+uxfrV2A7wHvMPF4XkCyMf
PPEEC6Q6vM6RHYv91QvUxak+sv7/RS5SHLubFcY3CIUQpjyzrDcCBT/+he8nENo8Rq6Ru8h6sv3c
TRsUdJXaMEcewh5KIEhChSH64GlHFG1ogzXl8csgSFaIkWFXjH3Gd2batDi7r4wrrT28Vv6ZYG02
t72rcGk5684ZZNiLgrjwyPhLTDFN6NuNjc7fJIlCXNCA2w2PjMPJ60TO/LEpQsDXKrVKfkv0a/Mh
WHzIyn3+1AWMNJgviQ5P3jWxJXOITipWJ8q6jw1M41wYPIkyrHXbLBI8KVqGFnho6EDh03OrbxSE
xnIjgWmgn3wIPatBMxk8L2bucMVrX+8mI+FhJGOv1t8c8C+fx9QwON1QbQ7zA+8J2eDjqwckS7ai
Y2I3qB++rwKUKiKCOGyltWRDHp06lwjmoxGL/O4tpNXhYXYKvBB1bUaU3AiX5CVudXkwYAS7/kmu
HHcYpK7enPKkz4Q8zyB7MhichO6w7o3r79eH0noGVTTmZmoKV9uVXmz1ibVaA58MG3/sLWPWcTQ3
mmQMfHVJ12deSF8J6cvXbJrG2m2EZEhY/yOqX2bbbvwW5oTNxPhpFg4NRaMKGgJbHdpWRSVxCFqm
VUyMQlzoNrjszkaxTPfTTUaYeUZdenqZVOO1+/OAvEK/HXdizVDdGf9u8UF2P0tJR5aPRWOONXwx
RN07dt3mO7Mj12sNC3xCJ9iBGG7PGhT8PSHN1CHfnkDI0plP4xpPU4yNW41JlohlPvNrgCS8YEk6
REqzffcEnwIIC0B6H9pjtHmbLWLwRF7lnk2cT6Fx3vmH2DIE2Ig5Y5UZm1Y+J/PRBH09j8YQnXxA
KtXUwjos0Xt00KBbhG81jiwdBMkgJnghKy53oC+W9uGmJ5boFp9BbccrkTBidnkxM4G6CKeJkcos
UagSFpRN4RUV2QlHrmuMz/C1hWDtrCn4G6J0Q5LvaK8oyy7I3TfL9PEcfSRQl4qfm/LsrBQ4xQp9
vUyuwIITg5j6VT1yLeWn+amTiNhkR6pAUhjHBJ4YLwTUZa2h+POz1oA2xnwbQ+rak72KpGuLJ2jd
5JwlkoAm0+ADv6+TOlfHlWIiw7G+J+LeXs+f5Mte3paHrZX4j1lbQPS2qrZJxwoNp67/Z7zwqV8/
Q09qlMxgoU9l+OImbagfrcUBlt/tv2qH0atBQiALg35PZp8AW0OBmjfKnxKF+tYJcgln0Yn78e/X
hDfJWS5Qm0GTjmDxl4wwU2ivi5m5ZJK1NopaoLt4Dknm2BTMheJglfNeBeq0bFg8nPnXQobzNqum
Z+sLNZPowrVEGjMsT1pNSopEoanBYS2QF8Q+mA2K0S8cZl0ZgrSd49Gqh5NjlgMfkgp3+BZd4ews
KSS+FIz+3ly9yWRWSkLKTfvlfYzPYDoZvPZdHpHuH/Ts8dfZrtw0lxIaEbIb446c025RiLRRff0g
lA7/H5Q2q7GiI4YNq4EUAzTh1czqSA8m9ZNT4u81UqqnUu/9jmZMujK1v8BrnGBRt2KZs4WG8DMM
yRVL7hUe5x/sbTIcpRDO6UfFRpl0Xqyd8V+uMjvh4dEjyijIn3dEDwuEvWOS0tgU//UJU6IaW9RV
+3shIgNLPRrfCXUb7gkOcXk7tO2Ygu681AbCA6z8+vwq+qeLV7kQSZbqUmtsBAeN4BfgBp1TlqEI
NAQTI8Fc3sFOM/ztDVH2g/ASSn4cVtqqRWbWKH4XocsxtkufAawDRizmHfTiwQykHsLScaSO1j2V
6MbEvY9SnvGVViRSo3K+kub28gGcBXNEqqIzjT92anX4DvjMG7E1jqHVvZO17wqASTrT+z2x6576
0gLKLFTDuWJGaUDGSZl9WxToqB+F5wBL/WmUM/DvhKxuHxLq+7pIm6u2m3mdfZEJ3O0iBnTstN0r
l8oFL+0HEBgNSlH1uOu5F9fa+HyMApLVXtJYCenSnC5TegLyNwBxxg5Qv4zvOaEqvCQCnaRQ8yi6
1XXPkZLGyUUdHQqXkpSHj0uLRa7JI5CepRTeBK2lpj8h8CorZg8gOobWWuHV0MfBGJDMs33Mkltm
aXnWtcWGvA6EFea5JjYV0SQqDnVHsrDIWmBCATYwpqR0pDW0ZeQP2NiA9m5Qj7Z2KJBmISwHHlQ3
LsFFQ6J8MhPFPRBnNVo3vcBzBVy58sM2kR25DDaAKxYP8Uy8RIclXRpSKl6qGU4mTy/8QGUy1DD7
iFzVPdY59TnhRyQsMSVj6uDat+fo/pqSaAtbyqYTK6C98H8TIhZ2iNgcQhZy3Pq8s1zxQdF8g3pq
yNwsff9ca16aLLevScoii5amnbe2PKo4weDEOWtBZziYbfRDFfx1PyOknKt0w8i4Rid6o+Q3wKYB
zK+NgxhoxeDuuNmWViw6dhMD63/juCCi6G/SpjCGw21eRaPIxSHsyGk2vLGsrrqSSK9vtiu66Cbt
3sx5Y92bSy5ZRcGM5qHUq1WPgx0EtBnMzsosaoJfDZs8H7tnzHEPQCn+N0sDcUhfIzVIxhxuePk8
ur9Q24chkUbUeek0JsCzMB1YWwmHpP3T/q9umnUdgIWYJxFV8W/xAggF7AECxdPycNY0++j7CnmV
JTsxvLWY9apZivrHWuZ3wYKuMxPekVD4nwMK6PomOoXgOQ3s8nBvyINzNGNiSHE7OxboQgFHJMGC
a4zRY1IySQPa9JBbx8MX/sUPad+jedMdDaWNXDw/i8dwEHSlFJd/oxlbLn/PW2FsSlb+3vwkKlOn
YpNHoD8MeCNm/UetgGi+/9zRv541A/eFqOZsdtO0WvBMOoAIZNzNDZpIsHwH7iFApJhHAgfrtEzF
Xbmv80MlTRPxVAmox3fa6xSENjBOksDjfIzaKXNshWd0kP05CtDfv3h3MhTlQP4ha+Jiu3PF5iGC
0Fn7nJDk1q+8xA2prv4BKUK/4LOmS/unp2jtGicJYI05RUd+5nPHFMnljUO/+JQmTZ76/ebbni3K
CKDktFGSVWAmgCOzGYrfDBb0G+kqru2O61DdC4rnJPUlfKt1Ii7M+bqxvlnf/v4Ssn2T3y+aFsne
LghPcl2wz3O9gEsr0b56W3sRpyGa/YuyNaOQ8ii8fik16OyiWTGCw/++Gp2qKYiGXRYdDT1JanOR
gtOuHplI6vJ4YkGwUv6m8jmmdgEAfcYaAcPpvFVKNcE/sGjyyYeqkbwaGHiIkbfqYHg4l9SOFiRO
KrOiyH0pzbtNkKoFoUDwuvueUSkf36SDrH+y21noha+g6KyDBum6QqH5gKD7JbH3WaUx7okR7Dqt
Rba3fjevvqewM8Y/BH1+Uik2Ojvs5p3cjbR4XCrKmaxBTrWmTg+liQ0HwCNh2QmEyO6dWxLStmOm
hFtMclNaRrqCR79spiP6ypRVTuflrOhr58IwO7QWC192byzwAN34ShL78nJwq7dYPz0QSNM+dCBg
ENjV5/eQfEvflzIcFIKOFFTyO8dU48qOMjzrRodlCgO8l1VU1QT1iQWl7A1x+KTF+TITiGyF7C4G
M2HMWk3ghT5hpgUfxCY1j4iLOdszzwohNrZrBDK8YktVMb6OnHACQh+f0BeSY/ttkDVYaa7Ihc5d
Ep8T+T970YE7iD2iXqabT8gAMw5w8GygYwbT4v8q1wnbeJ60BJS7l6FmZ8o37zEE4UQ3iiP+ckxB
jhmxCBjaFisgZnT0QuyzcMXwzQnmisH3YLMgs1lgDYClQjFZ3ouc2Fmy2w9HFIaAXfsECHq4jZNx
vYGHw6dMNjB7wp183NPqRuAqnKuw/MD4HkN+xnSyDl/rsO+XswZ1/rLhpvxGqPbo3pbiMspmNfwv
LGhY7w8D/6db8JiYtaS/fBBnSTKueYnrelrW9s41BbSBHvZk66VWELQkOIKvBPBk2A//rep/OTka
1mNKk4G/WIV6H62EtfUwk8rcpuCSeDVd/WIMaHThaYRt3Vwjeawlc4j4/8I32gzvhwyNJJ4Yr3R+
GeXpHPPpuAFf3yLQXk/UMN7MrdnTWWIlro9XrAGC8QJUd/LrzWIzP26bi1eLyevjYoWSFBR3WUDs
TiTOyYua3A3UIlLrYbJ34lLf5nbbgmi71pVJ+RpMcJ4yYOlqe+Axs7+ByNms4fgxJQVVPlwCl1a+
xl4kiLOzjFK7Nr41wsPj3KgoPykOWjAVwQ0FlTn0waFY5HKYeqG6x6eBRETgPUl+y4nVbH+7SN0n
NilzO5Vi2cNu1fNcBeDB9uEQtt6N+HtaWd7kThsycnWRWny9Jaji4NWImaXUslsG4zHBnN0zQGmC
JuRLZbF5d/IN0o8MbzlWPWpsTPeJwv6WtkhWwAZJpp1gvaq3QvlIjueQF3/XG0mKlNhuQ0E32nOo
2reW0kpm9Zg3QiskK1L3MgwDLIQVN+r0Xcczd4IFrLDEtVMNslYUcZYV8pL9L/USLe8Z5oauZO0+
rFextyS5rmGNwp4wm0goAzm3NmLKApunCnvE32Gwjz/ZTrpYOMUMOJTpXRX2QCqFG01eoH3Ur5o1
OiKK/DJvPLFDkl8Wmyjih1nFTRtv5KBxd8X1TuD8l1kqOOgCtV6+tQhA3nBnBzLkccIWAz/W+sBy
Y3D554QtZBodv7Bh7d7Oqstb1qv4nfVMUDomy79DXDHEjRRC+Z3g18oSUl6sa8gJr4xSeSOfcHHK
lB3df3QiEbbpwxucYtmwzMVYH4VOLu0ZATAwm1Sxx2DFi4OH0/e/sfZHPQxCNHNfi60QlKIUrHla
OurbxC8ShiyjkIq9xrQ0RO44RvrCMiP7Ak/p55LvbtJIFPWFPB/WGX1Yi9DrQ1v5inaafG8naXKe
29BMN5Jb/LjtsNcAuDrepytJZD0bx1XvpmCD+OlIvxxT8KujughOp44JYtO2lB349bOclvPJAYmV
2+nMTo3eKWXqpziOI4pMv8V5WhxC4dBzapO8DjRKs5ISbVqV27+AQKpjBpUj0Fp3lsSWa1PhF1Gb
pAZfi4Lk4VOTBAzOCdx7urGVBmAIER9RGozkVvhsbOzn9v1B4LkSSfey366eC3U4o0dS5KU7loSK
1LP0nIQ+lxryBixsFdcWICaGg94kPAga7nmj2hbtwXWgOmdTRSSrsw8vU92oCiRqQTRViqKZfs8i
k2ViDFHQU/9ayrvsmNn5nxuIjgOce/IWqHmgNc4F/46/1aSI0XSnRBBv4kWkMM0R3xrALzeUQ1ho
Wm/1LbdE29CMzQO4LjdHLYM4rtHxfp5aiZcJFtdXnOIakLXitD5gSiv8LKC6aFVS2sdz+ASeldk1
rkgZOl5ZdkCz8oH2rZhU1N3QVUH+kwq7GstihHWXn1WNRfhQZvoLs7MXrmwWS8MYGgOyS6zY9vn1
7XR+QjmP/EPMxxnArMD3ady7phAz4dm3NXDHiHwSb9OySuAagAkXVjmuysDHm104gD5SdKvM2D2Q
sk/xn+iBe2lNe9UlzH/Y9LxGqGhxdCZ4ymGZ5VdLG9RR37bwO6Q0PjycEZGUy8fVf1G/nR4mvkI2
5/90PIkz2Ynt5soEt1KDVmQQHgS946no+gw8PUT8E2sO24rDqQq/jYEFr1Gddi/kRHirxf9bbCRm
kZjMn/nYbURgnx1K/IoGHC5uWLTU5liNSXzu0a3ecAdhN4mXgKwnLS/A+UK2CQhbGCfCvFBo2CTF
KMVq51m6pP/XdHidNA+TvpQHmVHG7ZIQDF5RdvjUoxQPe7cd3RxtoIhLmZIpXFR9abvv2+BF9s4V
7X/arE6TgoFT6Vtp0WOPXjJ/KdSu3u3xEFvomFrGtT6xz5oHxgWg5bpiXF6UqQCUUvRcjxpRGJ5v
nqKF7WuxEZ/XVpegc5TSCB0VHULvKvkfvMyw44dvLb7E6INHea9Bgxl/HyHnBAYlL+TLf13pN+Vq
nAn/lZZDGNZ4pXpzZaLVdwNYzeATPJoLTvl1go7pE43ahzjqeZXEBr9Qq8osIFO1QW8kyq61ag3W
NtnQIXMs/ycktep6bKjiy4w7MfdESDQRJErY7xrWFPr7F7OafUllLvDkiIuouA4isy3RtwCZvaJ/
fo38VzBhJnkIn7HGJUpOPIOaCltx9IGz/qpUqqw8SKSF9z2KYYNnRxPV0M7etBwpXgkFzicGOR3e
3uQoiSr8QlgfoS/v7b3d4LZGlnKbtc0bMbv1Aw2u1cCTJ3eB0DQXpNsl5js0U1tEhE+5q4wUD+xQ
lBrGbzuyiHS719xHpKsLYjDviy4gchYVYQ7eVL6FnXq5m2Kpr7m7+sz4bIst3tJ+EtuGVIAmxiiq
k/boelh2PRrnbP2pHR3roEMuHeRHTSiA+FLXdzxrr7w+6/AbtXX9TXmFxOwclHikh3yAA7GFas8e
Zolse/yBb1vnAsoAA8BUuaCniJsK40ZBf90W+utTulntvyU1cJl1y7V/lPbHKQR+orxj+5/sO8Sc
Yd5PfWbPmQDTcWNDkSqvs4xYOwDClyeKL68sDqIYGDkp7AM4Y/txIj/m84wa22u5IJbE1vlET0lG
Jd/iximiSSi4dU9tDZZK5j9eRx9heuJZZZb+8azG/LP+YucPNrdjFIKULEhOPsvQGCQhtMeVTIfx
r8affHXbrQRq295imeggU3YqWTyoPiF7DcM706NC3wf96CSzDAaaaBm/9tBPRpO231uvT7lBOx+Y
QhwAfT63XlndRTOL/KBwZj2zEhzb70Zy4+HqNb11dFuiG/vSRD/wpVdV6MaHK/hz2khHg4/VWhHt
qH4RUjxkBoUryiRt8UG4qvrkjBDQgti7fG9SRBjbWlIqDMOchk/YVg5DwTztuxq/kjfc7Utl2T3g
Fq3JUkACpCVNbe/oK2jj18F1gML2ZoryTqh6iDYJgIpc03en5ss+8KzkZ0ygwrPnSMntOEpBuSyQ
SjR80BKrgZ9JFv0srVxkwbZSR7DfqcXdEuqK9paJU7jRVdI4A1XkcFmocOVEvfXHH5olkvj8Xtet
lnQff2Qh7IHtmbTUHh5sTkyvB+LtkKCTaYcZYf9gEo0JD87Fl+VnImafY/rZqEW01PvsoeDhlvVI
qeLydmNoeph5A2q4KidoILmnfQ2VHeMWgRAHO7r7WilEnbS4kWWS9tuY+PAg2xa5pDZ2tkh//eyh
Vd8/aUPMxAGzN6rIPMVx7CdmphTQoSI49WozSJtwiolEMPswdo2ykF3yRESwDo/+x5EdFJFy1IMg
RiGdoF3WSGeujconMcJk4xzMmDtl9D2edXU7V2qbQgAZF1oMm1mbKjY/YIBbi+dPfuYcrk3ERrCp
39L5khvRUypU8LwMrh5JymJUIUKZ+nVdTMrNlaL21tuMPI7BwZ6OTO+tfz8EUG6Tn9V+0T1u+aPI
/nvgQkLE5LdycCUNoKL7ZDvWkR/ZIskwLdKgxSNCrV3otU62VHXdNUgY23qQCWaicXUHm0EklOya
ctuE/MT62ZUM6dDPc/Y0wpPHuG4kjo75PCGe0MO9qsQuVJM73RDpIELqnMlWNoY0EzQAjpz3p/Di
JVZ8o/0du60h7hh7YzbNILOkBunEofD4vuy/Og3TGOv2lba963ef+cU0pjFkD9nKCwnMWJvbXsic
SefkO10XOcL6vXe1gh9dWXkCzt2YYJvcE/KfdZRhZw6gAM5A2JdsVpc586ECb9uYNKi4zXKJWYm4
LPYejI7yeLDmLVkpvugNl8MJhkKXR2hgNphxpTr/84IsC5T71YQDYpVhF6JVCJJW3B7AWy4/eP2S
fc8ZKSQgsG+nvbrQLkEwVLq//2uuhT5CjGv3MaQPMuSAF8vjg3VZGJqe6Df6G4wfjLaeu6LV6CAS
0brDM0hjGJI7DW3yDdyomvp8OCHjUnCeen1jnNOUmPloU8WYrdYyMBmRbhEg6FDJC+dad4LSMvE/
j8xt2UYHWeGw/a0At8JLa0wFtmVqcdeHv/UGU/jt6BpmT3X7OyrCwaOXIyaifsUWXARXaYww2ZLu
gBJ6hAbf8qTQh7AjiuMAZ6cxsrnjQijsVTOD8f+YYXf9vrBkc20on0aE/FeZsK10kziXsRgBaHZ4
vTf2tWHxm7t8E2QFT2HP5RNsQqHYkmiTZien0mBMacm29f7N/YbfJukuX7EtmKrgVADBeWJXry3W
dz5cY4oo9UU0kyr2m/8M9pkqiU6EVEE1kIF8MKQbtsy3MgvKH3sPs1U+WRx9m/mR6J1lQb1CY6L3
XUSyICqkC96tWtLloq+0NJrUmCc+dpD946iMcGERkcA/p72GAvOzoRk8BTiZYFsAw3LihhcBWwC1
EHboT7K8fidJbrLXTNPhDxPiwVJInQgVOJfw29liF5UyLuG33L9hhWtKvdnwnEZsi6gQ2YDxBYta
/kvdN2snrdkGgg4caBnQEmeMPaBkPPlHQyL8XkKHfs2Nv/2pXPG6PsYrz+NwYfjHXjBKa/1Wgy06
K9ErG6TifB8OWvmFAVZazEfmaMDhSrCrSQVHEtVLEDQpa2/qeKFuXRXcdfPaJUAh2f3CkiPJzFz2
/NjsMg9GfBtXdsOL79VdsSA1wPmmfMUVjA6FJ/Iz137eiu9VU/z+nzsAIV96A5QQWPwZgqjEf+YK
sdwEY27f5pzeh7hL84pVUrBre10ZIbTi5aDuceiCLrB+bFacgYPXE5bw4M6oJMMhpQM7RDF3WC34
p0yans7iGNC0oxtniveIWJb4SKrdHCxdpQDk9rHjqDKVZ0qWmh8txz93udIv6rUmODe0730xEzFa
WqoL3GBbtJs6vgW5GjqkILkAuXHubuXeIRs4nEAGCJocWMrq8w5VMVP1bFtKOx52yh1CdWoltRxe
xGni5uiYsSHbB3zAakaU9L510O6FOgkR9KpcZwvaI7hu1lsUBiw8CWkekzw9g8oThK0f30VZHEzV
2WBbgC9p9STCSxYAbqhPrIW+LgeRhRp1oD1pzY0zudWKfqLAhaOpklhooK2g7HY2hlH5jayAygLV
2lz7+OU06soUYoegpMa8W8j8+P5tNmb4Ivt5HtGxoPMY7pRezw9I3+RAlhtCqPB5pVm3Np51OTym
/ewGbScVbKD0Bi1FNm3OBB+8moC/NtWz+TfTOswrdiTUc4g3JTLlrnYnthrw8YzLN5Knzreg4ROI
lcCRpNT5lXQzdYCMl88QyRmsUllfYevSCOsDJjFoWiQIyoAGz6+H30EBwF4T8SjSoPVyYUA2wqw5
T0WTnc6SNKynPsE6JeoalTQzx51cev+vt/50pI1Ph/86xI/TWS3okHKVYCIyWwAkDo8BvKySHBpb
7p6GfDvcsGKm/lKUzSaDc9RgA0lSS/L8HElBY8FtfvsbAcLs6oMP78AJEIQiZB4kzzgVBvmsjNs7
nZQ11thqXo+HBwsWXlqf35uX5PpA6FgeOZYiaoO5CXKNZyLNtZjE52hkD9CGYxo1mW8fG2QKWnft
7U+cc+Qc7jt6g4tbN+imfhEfCJMhf4DmS4HbiTZV692XrKzue57Oja4OEIe5KEXZVq/Rfoiqi6wG
QSnz0obdMZlcgpOp96nFSAvXMqYgrLJO71uBd+LE/nuh8sgfE6jcjrg2Z6aRUlWqAgxcTLGFvwQh
Bs8399gG3WI8+SBk+ngbIrBFLFfbfmoqtyu8c8eCtBesqdylMibOo167mqGHUEHZ7dGSnAB16at5
udrNacX/LwRW8HO44/WVNTs8xGrKrD1Tr4hkojIXFZHNRDMNB+8TliLGaop+ClXVSh8gm+hntt3e
iTMvu2Ye2sBFGeV+qtBqQVE2pt2d38XScLz2KJ8NG+uAlWRKCb+bc7x6RwUKOiL4wOtntV5hcfid
JwqSpWvJS3PIkHIBT2sJXURqXVCBy3g4RWKovIDY7lGl8ZWZ5IiIpsQswOO9bcWEarpYaV77tM1A
MbZgyhYcWDi94GOpBXgGQPZVKdscT2FKPFrT6sTEc/tJt245iBw5Is2dpSTfZDYZih7Anm89LZm/
BHLKdakPeKnEtXmpF5mtbvyj2Ov+FK3hDq3zT+bs6wIP2cBf8lnxR1cyy8VvsJIsanPjbbuCDn3Z
J69kbQnJlQBUBQUW7/Qsaqhi7wArLADqtHCKv/JYHgFAdPrzdb1LJdDx7VWbkSwWhVliwEXXNhpZ
ri/K4eqMo1tJ0nP96YMYVyno5A8xhGf98YCsYElglZvLHx4N4OecJp/0Pk+kIcpxvymxe29e1hv+
Is9APwwQ+xpZ1LnEAvasi3/IZDGcjZw0jBvJGvwGS9glwCXyyADowIo3d+1UfWARVJprxgUtcvzG
QUVuNFveHbRIVQEwexBP8deuD9lDmT2xe3geWXFS26f+P/anad1c0DuGpj9hWnCG0Q2F7ACX7MKf
08vQhvPMSgbFSKMjSTo+XmU4UQRxkKRVMFPBKR4Pv+vvCCNZo6E3WoCgFeCcsvhXY7gUp3inpdy1
KN9WbtGmqaORvq5BL31X64nAERrDydqA24Hh7kTWBVjkisE0qZlFlXs82N4iGvrODdQG6WScKW0k
Eo5Zm2IHcMW28Gxcvee9S9RXiVV4o7fDSQOccF2Ky24g+SYUkeX56PeIUxgxeZxUwVO3cNOAI1rn
xEzYv9nKtuZ0DwNTUdANINY8YcVpbIl+NQKhGPoShx/2nlV7OOqXibxybWnSHr4d8aozuwoBNvtt
cXEyJidDSfRsdgHHAL1gvk+bt52PcnpbK2KfSDwn1yIGxT5pp4nCOeCFShiNZg9KFWpt/jtzseg8
UGs3l1Y2xqmprCb1RC6jHfCRJ/G/rixRSWFo+SzmVCUNBQNkDIqq77gemWgZpGVeWHK3UeJmwLtu
LInImV+ok/jTAFbqkXycztEOZNgpG9CQCmlqeOf7syQ9oYVQapsBG4xKm3/z/uYxlUxIUw7wgvnt
4et7V2G9SeugFa/TD8By/96K6MTC0kiYfMleBciXyFygU1jYoDCVWsZY/6zOkUni96eSm8oxR/tA
chT/IyGEyQ9nS7g4uoUrjPdHwqT2yrGWdI8s+cIDQqCmAObKmYHKjnwRBSdkvHNuEMifjvSAhbx+
CB9Ql/OaMcip0/ogtEZBaOS4RJhrans+ppSPIhqaJY74fOzLHPd1aM7tKottnMEbu314nV4CNrxY
eA0soJwbDcOKdemOLFp3ejnWUpI24pDnPb48ZBZFGpGGGJN6xJ5/UOiv9jtWLvcA3anJMIpMytAF
XpQJ15Qu39Xcs1Jqbp+qhkhfp866naiO8xz2efYLBS9R24ql0ZLEaB2dQbxgdQm2q6jQ5KnA8/nJ
ip0b50QnCkMKosou0RmUax62mwYkulPkFV9ZqyTn1TWSChOr3iPead3/mToPz5U03ZiCgkGy8I+Y
szkM9sU+2nxrFhHlDfHXb/skTVOYgHMGy/cRoQValLjGLErzRwcU4HoUCk2Sh43zYx9/3q3u5vDj
galoAmUlsvilWPJQbZMkrzp28joJFHJm6UVSeTgQmftIpaMd4XIpKRXb1MpnhcXXookeZCjg1KFm
POMULnNlqrtdN7FuswNRONZRs2YShBLrjw07LnW+O1panly+KW4/je3gph/dtfcPQ85bD6i9AiAT
1CR/FPjvSObMGlXnYrasgTQaJCfV7pwn+qYtTlwgYjqzkTTUlG/YoptbrgoOiuF293IFMlfZSRzL
BgDKGmNF/aIbPfJRb3WBjD5faLo4c/r7C6h6ZjbvdqPnPLJHd4iFTljGgdxdqZPfmNJdqbXoBx89
HHDED7K6X9AC/0vhrb2gYCbpVgF+fgncSbEpKKqCtV31fveWWtYpXK5QTkUDZaIU7ESK3UqSM+Bp
FrJDp5fmOL7W3aSv7PamzslCSkYcGzSoL/1aQo3CRFzKH0SKFPmvUIlyoR0NJyE9P2LmwrepIsaZ
kgGK2vfuVyLg0YmCeDWgTvLIyRMLhkBXgBtyrW5qUId8H1otFci65mBAYXQW2hsfM7rBbR6SNWSo
52LnTP7237iyd56qNxAKHZ0bsloHIHYpU/1qz/OeC1sWIMRwocfsOgV0Ls3nvUpByZQEvVx1nRWc
c9t/J8fXrKYEa8flMSCTXntH1jH2XZcWLqVwrr9mZpxkucu47Gwg7cVn8eL/PbbaCl9ZRCYvMCw8
C0Ds5CEkhBQf/YAtmgLjxkvu+iio6rS2yOTmnw8O+Z1kbGQZ8tACCAuRRBG4Rsy7NLnK1MHoVLVn
M5I0vyPvOYOQRmk1NMupW6BDniy0B0XZbpnN50Sj4R3jShRo1SLYNh+p+/0jFD1m39EZj8CMa+Hn
IcGhF2HbtUxq8ih+KCgItOYtEZc7Y8WlsJge5c6UZVgtwZjWhfMf1jqlJRQnE+wt+JIJphfQUNIX
euktrzA+oYtrTXf/JreFLFisJIrF3erbDnwnMlqiRbfcgbC90OF1u6z1oMs2BkPSPth2d4W8YRRX
GL8O7zW1JfpagColDCTavSgBp4petINuqYJ5zCFt42XmeaEZAv1hFsVsYwnGtY7cDZkbzIrrjuOe
BerJgdRheeIw0IZDXUCcrtMLY+Kog1I68N17RZ7Ue/N6A4cQgEu/pP5FtYacytgCDFWfsjZt42ya
JU+FaoB3q7SQ/JJb1wjrgt8V7AHHa0/1aXEfaJbrp9KJYJaUMgvS+3U2icQuqeT5ZlZsFR0wJIj5
D4J2V0sRJcUGcLUdoeqVHYHFRdqtPQUV7rQa3Jat8L9WnH7UrjZakaNJUL4+Ptg+K/B22mFP3Tqi
UiS0+O9J6Qkosxuk3lxSG2+Ykj6L9GvnR5WTG6P74wf3VxqomQsoHUeW7O+frTJ9QkEHSU+E7oVx
zvabswdeHYXDSzYqXd61rOpDgtuNgrO3cNT+TyzKqpjMPv4RpVNOu0fCO+oSjW9qadcOuwCGi94B
MREUm6G2XpnK++m5Ku3VdMgGFIduUI4YaGTAYQgnKTuD3hWHiLaucF9152oSyFu8aWCaMCixl0PX
+1BDCuUVpJUMK0lppWsgU8C0NbYbuQk/CB85AItrqtNPQIeKiT+QxalmAv86OwmGzf4oAbfDkxNZ
JX0QezFolcsTbnmYwk2GP971XRjjRMwJ4VKdm5NCvfw/qdqdIBvGE/D4z7bWajvRu7IViMXLKgvl
UoMMB3MYNqmYVrJdBoIOIq+D9IePiFSRUKbGZj6rIEhLB74SntN0F8ZEsfjmr4r7gHxcZQ29MwVS
drXECEUhXaq27goXGFL3vaMDym+mcHFrVc1TT88RXyhotCD8CaDwmwmsdfXRF+KquclSUxulor5R
A99gYjkBM6HGs7ggd+XR/3y/Sf6FFdt/ucvzmVE2Sxa12YiyOaP4aEqwOi7P4p1CDWG/V0OHFrAW
JMXp3UAradljMK//NNB+PO+hXbRyoy0wBTIsCQ+8gxAO8OUVxn9F+GZMWUZYgl3vEzBqxZyFSPFJ
hoiQaiW5tRCZICNU4riW5NPh6ok293p9VIdHEXICxh+LHFubpC3cQth9JKhj5voZ1U3AlZUd4vbw
d176aKUDzdWNlziGEHXcbbyLoFvMU5mHIwLBN5bRfIYn+g9O6KJBIjGDGxOu+hxb+Xt+XK4ie0g8
mg/z9zaSK1soxLRsjScGZqIRNRJNQxyhW5b2Wx+FFKAoXtF1e7Gu2Nq6bLi/2tozG7DSUv+sXIIV
wVGvTzWUwmCSFh+Zae9WQ9puhqLbewCkHQCmKV4Zr7Nk700OdXGLsKqIx2zdcpmNPO9cA7Euf18z
2XtKONGd6ywTWtIZ+CSVSDcYElJAMuHsv1kJBTEuSx0P12j7hIPayjXiTxQCoYF2+pwvi28Ur6Pv
fFPS6jggtkiKydnslxfvD8JXuA5bCQipqUemkwoc1LzrsHWZqVKwL819sV7Dem8sfTY8JQRFjgp0
i7dOxD6Suy4II0RRFAiCZyFoMkfOYpx/JA03assJdsG5RhWx2skvzO5JhIBmzCpqb3M45upA643h
ySDT/yZ9UXkees1buMj7LU5MbEEPtrhv7b6++yc2IWjYdmEBxSqxGpcA/UAM8ABf0+n8eyCjoNSh
W3lynM/JzWfeswFv/DbNP0HZM0Kn8c14nJG7MWNfQm3cHfS7D2ELCBvAzcBwpQhgyKLyatrcIulZ
HxLGwA0Xr7yEpQVTdsirqlVn9siPuApr8Xdov02ZRS6S06AaF+rYKogEVmxw6ClACuCGWP7TKMEB
lGIqdkZOIoUQuvhVPfBilq4yqrBb2ZfL4MulJf5pSjK3asQ/UwbGCcS7dZ+/VPzc4baZaIOqOv72
aUMT6y7gAlV/0MTnG221GTk9mNnDXr038d+TllmyyNbJ7TObVGdboQISFjAVrhBB+cLjivXUejio
DWsobjUtHL3Cj5znBrfsmLOfCwP2LA2cTkG+7ssvIXnz3MGy3jn2dFcne1saFuBla9zBlrB/rdzG
jdkH5O6C1IkvnrHyGP97JYp3wpQAY2FdQfP9bmEqIk1YOlOYxz30IJm0ZIBwQT5B3YQ27fkCRhw9
Kpzjb+et4JjHU9738+Xt+OVpnnbfmDwOd9HZyvM+k8g1urb5gZ0JFIeaAspF/hsn95VhUFkVejyH
iDVpuQGRP2fCDklxTx1ToUL+3pujCZC85gw7o30V0vAYgA9KQzzsbcP1l385CYi7Vo/V1Ag0saex
he4aobyCqQ5YIliDPpG3N9MpqL5rgSvp2H9rjY4G0X79j26f0pwjMNJuMYmIBQCZmJnd7Y/jF7z7
xUteW6Lws68w5jJWDNENSMtn9k6nVofcsbgR5KyFa4TGg8KNxaM4Kpsqz9kYmj/s8qkA2+gOoNZn
89whIjE7NmIdCtN3080H+1fa/eAHvbIwfPCjK8AFN1X3LFwyMfGG11Tc6wG1Ajap1mbvbtQr/8cv
hgJ5dBO3oRvHkkIAEJGt8XzEgk12d95ZBhsZ2uDvisbJ0+mJT+jFbfDJSR07CAozc6r3oTwjjzGH
C3W4THAeyEiAeRmlFK3RoFjrDMEoq/rmPgp3bki+rb8AqDXw6n8Ce4ZTKtkEkYcE+cKiAOQ1f+eb
GA96UKQE0VpZjeeXQs4OTK/Xjuq+Ct+KPifAGAFIlTuEvOusKor3iGvRg8RZF/etePWXRUQ187QZ
+0udrMYP8nD06P8T6rEH9is020TG4ja+Fe14rn7KUNOsPmgazxCD6ld5KFrv4jXBOoSZgE2gMo4t
Qln1CGuvQCiS1g0ElLXmFtG+sYSjZhFifH+T6qgo7C/0FHB0U5SDE5nNaH/N0henJ2gY2TLWCRYY
ECvO+oFeeBWOOJPuM1wyWTrwCIJmMcChWwaww1xQS3nJTa//sthWc+JF/wTF4K4ThTbZQ2veARuX
KM8cQ4aCSN+i21JIK4q7L1cxEqUZwYPkLPAmTENNrobsru3jh+1e51R1g2CsTjrkROdU/DdayfS3
47whF1EoOXuP2Iji+zG1WHMa8+12rsGm5+kfNHpQJZkgXf5lOKwVlF1tAYSvVsAizcgAmiO+o81d
h8zBUdSxMUCkYJQnen6sw6HLvcxbp5ZqfM9l0o2pFyihPUtbx6kG9ISEI5vSyHSI3qcgYD4mBSaq
62/dzMDdw4L4Gb4aeb8eEa3jORVV+hAY1955O/Fu/Z2gN5uftR0pkSe1LnuVL/5kPsUXRY+9ENMy
zMneqS+dAaSfQCofRcZ+sI53HtoFl7cA5GC7Ndta7PpxGT37SswzIynNqqihNh8YzvNnushKZHSu
Khvn4m+BAO+UD2hVy6xdQJGZ7wkTOcTQKrD9IktPQcbcqLIfY6B8jtxWlVD2GBCMUI0JIPe6sPpO
DDjPhuX7gbI3VrOasluZZCv+m3GBZ3OGxXUcOMK+QvKRQdNpTKNwliec0UZWmKATvk/T+nMbXP8z
+9dhi3TLaxHu4R/Ns3fxJQQ7ST8piGN8prtIIs2qkWiWdmGFNqcOyvkZCjbBM9NtLVZA2KnL/Jjd
uJMDdoTY46EP1aqO2XZigGo2XMLtia9hPlLBtcOJnXvXj76G6plPw+Fk3xZBIAI0ldFS4lO6Hu4C
bSOgKP+8js+mVmqb+TriMh/RuJKQs8tVccP1Q+9B5SVawZBtHiHHHRz7FaZXY6Nl56Ua6+7YoDdW
9F5QxM66A/eRcEB5VXdJ84SGXp4nUkv/zlj/Cvq5X5dxN359xWakam+xHezaypv04GZgiat+tiAh
3RrYSLsrcurhmDSku0miMn4Ek0f+w1WT7+67JS2Q+XcpY2w/I4Sx1QtSX10dhAwye8awrGCukR7j
wA8xS/qq2cdjii7Q2F/93pDXtiblZ13soH+udY9RPenxj3cfVHSTOeSWX8as1Gqs093HSFeam9SH
ArKlJVV+PPfbJuRt8shNCVtqmqnjkM1GdCeq58LX5+y0IRNN70wxHUPKhZCPqaRPOk7PXPl0gqqs
SZkuWmx/DbmHJl0Kj62thKlVVF+khITf8LjmD1ez3LLNomZ6ApIvXV7iy+ViE2wjREboItK1F6Nh
oR77vHEii2zS3taVFgXRmMqWzYdtTYnnYFNDdJjV9xjnHR7EgJVNAix7kbm38JCt4xkcqZl5dw44
xfAwEhHUlGAanl+zEg7kKIZoeUx5v1ZwlqKc8UlrJrjZtnEEEbMmCpGJg55xtBU1ZPD3VdIaexkZ
NMpM1T0ve1YrYFhV9JQOSqRoqmwVnB5CshLuV0vkPJOcHzrY0CAYOQVueNyHJFYDhE058OAJHk7F
kDE79+oE9dEzbcMKRz9u4NC8jNYLzB6EOZdM+erVwqUZm5jEHE43MrhqI2PS4ENICZypkxiq0x1c
pxyqGDNtwYQjAjum27QL/dkom5dqKrHngkahkuYvVXseE5Qk6IOn+uo1HTFj4zhbjrMT5VNjsMDZ
dXTgam3ljGy7RWZtgu0UPT9ZOzzIqQGuCSYNVoqCUSYHYlRR8kAgSB0LblYjagSpoJZC9IcsD4Zi
jXXKir3bgIZYAsDKYVueJwXqxH4+souymQDub8zVz4C2wg9BR3BGyQ+jQlZ3Wj7E80MhrmudQCir
mYqct6io/zV9WGqW4MkVq3CKE995frQZ48KvtTS2t3FMk79dj4hTrHJ9CAc8HKs1K2SmwriwY2qv
LWPOQ7eEVWNEBiiW/icwhPKIRLw4zA13n/R1+WcXlU9K4JPfZ8tWJ5naHuPdgPiP3adZKGyMeB/w
GBPu3U6jcQSdHE91bWNK2tEM2qY3GWJwtmDnuAKalqcsI4Y5rLi6+VVbqB59djraoFSmRbJA87nV
s4CLE8UNVTZXLN0XnJ2tbpbJ6DWM415LCI+Q9SeaMpkLgCsXTCjNIZlqH7NcYn7DQ/5rgoZG/hJK
IN+zb/Jd33EcYKf3qzAXFLGlgA8O9iEKVhsWOPrTh2utGsNYiHidDRAHbEHotb3HJ2nIvZd/cVeh
JD48gBwmGYEI7kjlFHn9UuTSxeZLtUBL2YESHrP+HtGIzDlQpl6P+0JQj6RyGMea6hPhbxItv5G5
vJSAQpFLn7zHgywSEnt8fmG6HXrc3p/YyjzrQuARoxOPXtirARJ+vkQconjmGiUODCcd57Xb28kv
7cFGWTH6muj5dMGRpKGsBW59Rz2zaUj2YVA5g5LIi/H30yENW65SqKsetwCmMDIDNUZBqfobD4gw
kfnqL50EKh5W90NBcLMR3t4ZC7WWW+Ciup0WHLWTDNoo0WmM5zn1APD882NVz95UXhzmX9tN7fWt
eu/QlchdSjP3qPOiYnWC6qzuTbBi5jo+8MSyjc/A0vAejXtIXSXLspunGHwsAlrHQMXyVxhY5wk4
nZ4Sk0a4Wxk+vemjI5HGM4M7pltU+611X6JH4Oma5563DVn0FG6xfWh2EF7NKsdjaz4jEXFVHCUb
eCp/E7ydNWFbc+0MlE2uKY3yRmiYOvim5hJONpbZ0SQ0ubAuNwo9yyBE8LvAZNa0oqMWFdDzfphV
HW17EXo2j4+Gv/MF0SJnKs6vTRGlNuMhDFTVpzOArZoc1XO7M08RbRuhafbiUEepUjJi9mwj/Ppa
R7TDuBhgqlv0vviqbpm7lBmBb+kf1q9RVQj/H4A547xFeFc1IofzA3/zEUFOuYsiELrR+yWSSDpb
Mrkjdx9pdQwspko5CiRB/04QlPH30xahk+Z0iBLo+tgezHJI33p4inmdy/kAUZlyQNSRqnL1NiWB
J2LCexdRXPrs9685hKLShrSVA+0ssxPyU8QDIzQ4aB+ib3iwCeno2LZKgg44rx7d8h+YdfZy8H+0
lp/6SHvaLQtQzI5mr7AZrNPNEqswnTlXo+n2AklzWnQHXn6RYeu6pe9dRPIIkIsdSc8/IGi+4CiT
KfFEy2BHf3os9tRhQCm/Yfh3YymDTw1F9WI6RfxPAqIxw5o4Aj17/Z3kybl0FxpMmtte4Pi0iRd6
zBMCHlKVBjMUnmNVGxBqkLjclTo1mWxhhRin6fa09qMEi9fs0yqDVwR0Zm5jaNOJq5AMUR/JWJUR
hB5W912CgI7i/MVeqLEdW5ojtzqucEOMe704Y+mc9wM7pE9/49U/dxQ30bC2XnaWoYns9TzD2hMp
VIJds4F12NVX5pReDLPlBAxS4uGliJ68Rit6153WtL+vFeGvNJNAuPSrMeN9gPKN7c61k1JxSna/
FTT2mT1ulAJKUySR753pT4hxfP81ZO1smQ6ZrtNf6xPUxuBrj0r3IMwhTYUV530n0uGNPHsJCx7S
amMLlm22RPwnQH0b0GC+UTAEcw3m+VsUxyOWzDUwmSKUnO+V3xbKdaLJjLLvGcVqwHUvNr2nv8aP
atg+7rJeGCVRV1C2fjyNhRqTQhKDSgtVZkQr8gjlvUvn0l1gg8GO9P7o0uyAc6f/8CX0Bvsmzalq
yeMRXGzDp8fR8Y90DBiV8+Vt+9kgF+JPH/vloBI/8xspbvb+6Xg2atYKfrl8hQe+a5sNNXIbQEFM
ZCPc2nwrOfAZXMvDzBlapsSgShoI08hMo8/HgmyXlFokyDEmqdFc3T+dn2sszz1hfblN7zskpmgz
OzKdsLzweKGkwvP27Fep8QuYoMdPCHx+K6OQD/mJcvLH0+hB7OEkb9llWdiIE5Kqo7arPg1b4LJD
WjsvtLW8WprdX/xA7rdAIXS+xo34lnC8cz/4h1JkvQ1N6Ahrjmnx35Zt+6Cf0SavhjEpwpB5M6PC
uiHGnXY+byGnz4M3HdHc/QjNmWx/KuvUeFWh+5va1vvWlBfgmv5DlEgba4RPM+lyXTeTMRRTcCS5
2rg5q6owpzQVnsH9n9c7VuMJQ5qDK15QPMgypeJfPOe+dxF0jlbq/ym3Qv8ZO/zv00PeB+5fxuTl
vJXmmmYlvyCmqgxE3Wc/QLXrbOR6WGBtpGGDnAKzWipycY9Ns6fWprv9F09GbpWA0brfl+yLeB7y
paMpSNYKmDnyPxzL1+9InJ/gGRRxW2JiOMkjYQ71lUbF3EBO2am5Ms+Iu/IzjMIt2VqOAJS1d5tf
HpYZxBNOAffccLq/7BaRotCL5V9KCt0aq6FbuXXr9lgK2N7m1DjsAnYpCxHUROYyDgiLxmTgtO9Q
sn0Ove/Hjoreesn4YQTLy2cQrOpNsCDinTYq1F713xDYyLWeCbk+8tdDAMwaLmoUaQtBftKlX6jk
ke6yCRIePAi23yY/vTLtAnlzciGErRiKEB4N/MnbXOCflwoO/CyH1ZOTIFINw6UXvXlUsya3Tt3H
f9xyQYOZm8/qSnFIu/p4ce5t7UVDvVW58eVLy0vpAjYFdYYozRdHYEqDK4X3E6vS1S5cN1H2PnyC
yIl13R2clWTEPn0Cnm3LK6u5LwCneF6UBVk253AZ8x35rtYOk0i6GcLFG8fWUhidmUgPvMj7bMaP
g55Zm3rcdG3xGr1CSSXYsq6qk45oBw5xG/wnv20WZEhuBBV4NscR114aJFGv6NBcF5s1XGD11Jm0
0/HY4WnaQdY3ug4WXxeo9MnDQ5YADXFZQDhjCS+aHR/8xl7jVim+3FGcwhMhhKF5hB2iq0HxPXbN
PqeuaYclyQapucNRk2nZIEi2BGTyccs2cV9VOz4/oPI8s6322Qx+gwrEUEVatow+HJ2UZ89xELQZ
HBx13WzNrMZryWn0bjE30hl+fPJcIfTJJSHY0NWbxjJCFvPyvswkvHaq9NIgCJfW760Aai/Asdby
oA7uPZgvABU3yVgLrrOS1Qkpt8QzXQVGecoi5/cQYBMg1zMz2Qic5UB6bJfLMzqRID9xeW15aSJO
NXDqTLZz0ASHgfFs4WY1wWnlA6a/JhucO7nfloWp00Kh74t1IvUGcHXfKp1dQRhb4GDtyL2QSdFa
CqucOcxjJBVwiZ6Fmwi0+0Ip7OZquxaQsVWtLo0+XptBU+8bOb1qk9HttSWre7xKXXdfl8mhzuLO
IdNCSfRq9wmWIrG6INBaE/l4i9q+u2SiVkv+adrakcxXcfJr7v537nIbQmkYbBWM3JUUPI/m8u5P
hhdOeOXdnEhqnWYNxU3oN7kBywKPPckOmLkRYYTGHXMvJSHFjGaKnzeHSIGJx2/M9H9xM9jNUuiQ
G+5EVffAKYLZXoPh6z1vbGmBcJcoWisUTkVtDH2Z/Zq8tY56Tpn2K3TehQjskWoPGzJ7tngGGC6U
s+GvvJiTVRKGcmfC3zpMuuOeSZxFGtPMnAcAnrnqsm2lEmbHloGRTk325uKAptIKWi9Q9XXuWRrr
/rhtQSXyWUscpdq+vdRKZNB5b1cEUQWqlOxD1Oz6GkVLztrGRKTDZKzrXYI5m69yZP9jxnbwq5rv
EkaAI7ciQEZM3/8GhRMuQvhx3v9h2RMyYb6q4MsRQy1zlNVM2xpkk48F1RI2UIITjqIs/nerA3Co
XvA9BaQL2rj4HKZAUpwZUEyQiQH1EgyRoWnO5npKrSGePURGSYJe1SZ2t0374bsc6IYhVJXOSs8J
jSP1E++OX0wNRo6PDSuZu9tcEW/4vQ72l5mafhQOkKZOe5Pq/BS2Y7dzCnryBq9wd+GC4sBMF3l1
YK2d+QP2yvd6dONmiqtOwYOlnjw/apEl53Ow71E/nMXA2x35uW21Zq6CvYhbqIcz/5He0/hA/STn
9fq8YmfLA2Nu9TJKAhIlzkUAJB+IgWZJ1xQWJCEuqo3Xo5mGRl6DMsOIvPqQbnwQLKuLbSSB1Mc9
3RuoYCpVj4urnJVJI3RUdNl7wboJk6tLYk9RJDByeISogYSpfKouQdB75+EbuRRSzmIvhQukVIb/
kz/FIeAH19QPHlAGxzXeC2pPDMJ41HDBWTy93qqPNnhUOzPioLQnthBcEk85T9yCHOoE3bnC1XDN
zhZ5W7rl1/oy9r+nXx0BTckHElNj/zAg5ne2t51YxWdd4gK3O1OX2cSqfMnWqnie+ZR3ZdqDHCC3
bLebNeACuaBcuoEIy9blWC6OSSPP+QPIKitMvahEoXbxUpEuz5XbljotNZsjYa9k+F1jKL2KctJK
7oXQpAqP7LzZQjUnGjC5qoNiTqoQV8xEddMudYFJqwNUM7UWQF6WOgoc3/2p+bcXXFVHYpiORkL1
KiSZWib9L2eyikW5QYKH/YgL9OlgndD/uQBbr0qSr7iWPx+SzUIHuJkXB0UVDtsCixPynt8yk9bR
JKq11x1zpwMqCv1fWa/Z18u8XmuEsUoY1/1YSZjVqLQbrlRU/h0eysfZL5XsP9KRKGZ8MnACzBU+
rx0VkpRsbuSBotftU++ra0AXCWzp6SElsPByVirVLONXU9ePXhSz+iHDsbOIt0RTinQbQofF0g5d
XWgg1eDv3fFUFmUIBrADL1WjziMgkhDkVADsov+JP52xeiKcWeP3+qcQnVAORfMwHl6hkIxvG3yr
Nnd8/pK4aIPAqhJFFAO6Vjmn98OgMcpfQ0kjToE/1TWx6gPO2jf0BcB2EDKKAC5Cr2+hOkDxj1yn
fJO+ghmahb9urFThB6lq1BQOF6s71/NM28R/vIWyUAk9IJD+bHgwrQ6tTHk9qbTEs0GRhMaWXd8B
kMojvf814XKOAxs/VNLT3n64WAU+p5WEuZbVxB3aHXYqPQE8xUyljUvim+1C4aIE4mRs0h2jTaIi
YNuJ2w8+4UM5ISxRj/DuPxzZUWvnyIY4nTYF94IVCN+q4h3iRfdti4AUWtJfPD5iiUiO9KAbygse
voEaA2SR60dnypwEXZ6i8f2XyGvEwvZLyg8oOh+qxXnaW9RHedFDTjiS6/Tu5ci4Z4nyw6rN4Jw8
JXB2eTaQGyEpkyZ1629JE4u/hTuwHd6hk2okSMXtoMjyKHrr42d6XwuimrV+iHuXKVWwOGwrn5o7
tiy7z+I76CgerUMXzpv9vRuW2NP2YTdAUcuE8MhBlhQEUSui477pSstJ9+rUPzfiwsC9fwkuRa9f
ZDbr1PB8UXbF7oT0xj7VN1fGJMTC6HNU5gI3em8xwpnmYVwdErKQ8VXsZ5L+2ZywjJOXQYVL9E+q
9CIp0Xj5oVr6A1AbXBISOXRQ49K0x26cWAhM5WotFNawFw0TAFr2MSca3meULNveRfzvK3AVwrjC
PUe8v6MamDPaqg0hMc22TwNOc5HpQAN64SlaOdB2EmfNFcghKIE4sSgd3w5wjODLjpvRD2137al7
cX8tMc2ZWqMOJF6c25Ar/wV+Xit9r1ZBTn2KzDhWqHaM0DERKuc+Rq3x9D41bYcxvcPgAhhrYmiR
ANcUSUUWAGqckGGq02DiUhKoOus+5fvqkGGbb/3IlWYFxCnaW2sX9r+aIHI0q7H/ludhe7SMvhYR
HTKppSLiZ3qCwRMup5qV53Nr+5LlOZiUZQBdnUCt4q2e8BSQluI+xg+a/v/DRYBjASoTnDtJLwVI
f1I7bj07QJt1SC2FU2w6yCT3HOOp0LwKwwmDiTBO5tQY3uwYiVW55tvfScq3a6zLVkbZmPa9LIAF
wlzOyvXv1Z8xft1yZg5GeHAUImTYCPFQk4hXYTd5u69NQZX39qLx1YbRHFUNsq4Nr9U4MHMnnu/m
6qAMk6esHs66QgXHzcPJ28WC6P9/qhBe5ODOHMnsXFnw5aqnkjjOr1WS78Hj6oWEcL1KtJyf/bZ2
PNSmmXtNLP76cmZtWrAid7hTGi46ocBfbcPr4DRQPa+g86g21Llr5B68v7WYOIfH3HbVvAbZy+HN
Rmu+lEK0am+jhh0nd3h0lgJaNSNPonn3fSPU+uqY2kvxgUUj9tE9H793hVUPJdpYNShWGEtpKrKZ
ilnlS5z5PN7bY8g9ywHU3oMaPIh5Nt1bK5J9qfQH2Gxx691jarwR4KgxSHcTHfWy3RFN0NsPu06J
zSiqmA2+nn0zgfyZMOj49cuEZd3adX77cgOFxI219JbVzCxpR0GsuOZ1ZYORGD5k4Q+B5gNG4ISQ
aPPmZRXOhrqGIZJFhL8L6N5P4CoW1ISvekMEuOAFCtHkJi0EIYQVqOObpeeSOsjKrMoe9DGJAC2y
mZLmpCF6l8bF8AjH85oBeFLp8ajIGLcF3SLNMmntlu9t/7dGTHFNzG6hOG1RPf6x2FbRNC6j1suF
RNXMNos1cxoxOc1actzayxavd/m+UcF1/XP8iHzk3lruxAOOnG9Ia3iHYVGriut5cj1euGRIvgvW
rwCXlBUA8x2R9sbOZT8MXypEQMJpz8vC/6vEXRf6Oh88WFTKW9cYAAx+ZxOwpayWeKNWfB7nRq9Y
Xt5cdNQhefwjAOFRsi9h5izlR9CLOIhXPVCN4egbZv3V+Leh+rc/50MbpgLanSalUuqrxjoswYwk
eavmBPNWOKt7S2Nc7X9FUjb06Sw0ABbbWTCR5B8DoEDzDF8+4/03haJHrL0qotRwKRErxFOK+daV
lD5tqVSpvssPuCZa+8+1AQ6gzdaT2vjo2d922QD6V4iqTCQzpbKZYblRLtWbZOIfe/t2BXom0Htw
NzoVPyREElXBaq3zXWXF+tnHPnrhLAaDb/t2K0c2T6m8QsQs9en4aeCtdy/+5rI/VXer9ghttloL
yvynUfETd9ZNBi1AZQBQ58EZDzqKubN7P5IHDiGHs12axQnypwuZpg5aUqVXcvAvXTDHTuA8EyLK
cFN6Fz/V2/9hYzo9ieH+n1VYit8Za9n4Gqe+wRncJq2uMg/3HoJaCPjqn2TiLpFcAD1vaSUWCquF
N5wKNnX2pa9CoHTnRmwu3Syj6GyCvnMCQq+4bFlQKVL9dlH+Kd+5whpDStGe1jtRLz1lmQAewfht
sC2JKhGOxLIiLd8MkjMT2PiJifpqe9Jt9oVR0ZVXwJlj2kJOb2EzZWjhZBgU2cojeJeHXL+hsuu/
KrpcA8Yhfn8IhRzFI7B4QS4jJ3MEjn6FrsyE6OfxhuoWckP0ijy+xlBoc0r2wAhtOuIZ1OiPbjap
03lYP2xu8N2YH0KstieW3FDqgabc7agNRcVlgi3cK0ePtx+WoG6C+zbBcnR3SN8kr5Uo92hv/I5j
fcIj5KI8sux6l8ZqZgs2PsRnnnIk3YS5HiYxOnLirwh5lbL+6gCGhNtJKgPUnKG1mZ2f267xJhlK
76CBoiuHFzmI0ai3J2ivaOp5u8EM/HK9+w7qBc9YB5JBoKcd2anKhwz74V2BzuhKyPITaKU+QQBL
+1pzivp+isjKYdJTDb6hVU/t24u5A79dCNz3ASETg5NuSRbXf6it3ziYrBYA+VlHDOnx2EGcfF7f
u6GR7Lb/cGKysNTn10v7fN478RQXekgGLjxNhXJco+WN+IUofeFFUdpsYRkQC7UNuZ8dfMezkHZ2
EXljaVphhZOwb9k7GgXpqFYNHlf4Ttty8m7YlThD39Vki7RTkxET7QScbimiIvLicVjzpCJ0x7e8
ptxeQmr/nh5hPjTODl69plGz8TfQLEuAnKd3NupjjSXG2XXl/S3hYqIyWXIbktLLEAJwsOuW2Yf/
iCwyxDIDXlHGE2CaJnPpmgX1cYpTqTMyN2iCDyIUb/Fl48nXXtu+oACgbU5noR96hyIVqZyU55o+
eDrbvDyBkxfjR1TLVHNi3aYigeJR9Aslv+kiSpBEoNnigGmSjaDl2VK2xbH3yW4qhS3X3Km07mJS
bo6NgRsoHirnM5Sj3SEOXkwwg1BISk+htQFGBNt3n916fef7NQLqipLGgD9DHng5jMAblj/B2Qbz
zaYCvYwxt+sb78lke4AbW+PP2BCzfGmDnQzZXwyg/XRSArsIBQgfN6sq18WEZvHx40C0qtFWYVOc
bt5EGlnIjXV1rSUk1bPaaQvePTrP9kAhfhrZaMoJjjPHOZ/hlvyhxKgTIng4qM3neqQaj7sXMPpT
7pVKiFuP/jdc6mnzM1AW8EHHTL4A0eCD7fOL6qH6fkId9jqLYVpAIZEhYJdeK2q1iaUPDaRTY7y2
rP4FP8xj4DnoyqcKJghzbD6bAOdE5bmuyQycG3QpTa/brzGsMK177WcvbQvvTZAcDIzZpsYYWCPX
4bFQ+BWWMbacqIszsXxHnrpRlq9tJxA2ksKiuRACBn3cbOMEt3Y7Re4KNi7ida+Pl3dMuNR/dv9A
p+QDgJwYLPS8N8pHB7Wv1i+WKJ6N5Be+0TrEykO3vWWWDsv1M6giKxVRqnS6GLgquzKkb066c/30
lHf3aLG0gW1yDUrsvD55eEyExAVN7Q9mGqf8KmGrcpEOEMYhprZlSHCmIfyx+JG80JeJGiIZ7G2n
O37htykrEAFyiYCcyt1QRl3/6A4uM0ksakEp1NHKe/iLHMoGmmZr+hBlJrd98ellb249T2IqYcGQ
vKOs6ncLXYx8YI5EfYhzIIc3gJO+mCHRt1VmlNNWo0VVRgge4F9Rr2axPaWsMUpICcxcnhBgbo/t
fHIMN/RjaK9v9efVTYCjMdGgDJW1HjOJNnXbwWXTHoMtHFetCYmpYp332D5K7P6txSASdqN12nFv
GQPQbpcHRzgVLTO7Z5iNRUacfFVEilmYe2fvEXDC5/NzKFz+cvrCZ2qX5yCekWliRFPmTORX/gr3
Ky6jUPuMqGccaSsb5Ogx0vQecFpfXV3TCcFb5OfYGJ7U6/9ZzjN9t1GZoqnyE0Lavgx+2DYLhor+
i4Wb1Vc+iyTsSGLNL9R59xrU9MvfkGK7/yIle+NEptY43erd25M7gKAkZiJ1X8lRbgOIxODqMaSb
6h7tc7Aol5DvhgPKTFB/+ywz2Yr/uGRaM4N33avzQjfGm3iyaUujCHbm6slQb8zKhBGWJEESBVKZ
G8ONkbWDkzWsNhSOGRtgohpw6k8MTU/6z2XhGy/VHFAzGfGog5Vzzw94nQjGGqOatw1bAUOjMaKW
PwC9s8/0Uca0WVr3URaoyTh60b68GHoAtz6OJPIj5j+tuv6vKmcEW9ETvap0tWelqRtg/qK5ozmA
04JBh8yYlasm3RpAx9URzlQrbBS10tiIT3fVW+IbIx+OMFkKOYalD/SUGhq8PzLOkhBG/AyflxJ1
hqQRk3tHx2yAVhkx7vEIFHmjdq0+fBPiakLaLjhfjFcUB6STQyBO0S9W1A+dIDLsG1D1NtH84WH8
FQtPaRwww4q50xB7FRnmqFxyoC0s61HiHHt5RwpKD3D8lK6cTsZm0VTdcY6IcFubLCaCuCcL0mdi
8yIAOnVpjS8JK94e9iIzhXr3TYYbdjBasFr7F1Y5MXLp6bTOSTrInvZ9VHCpvk5LF41efBUMVqs2
+LXsdhV9/YTabq7iN9dkvITrMyk7Ka6MPO8WMeyaXMNCfhVJWeYJpZc6jv1U7pJz9dmlCVIyV50j
B0VowbpMItMD0vxQcaCRO+MV9xOdgj9/Wb7rDtUR8b/2iUIyji+/0g+vAfet/7gsMV7DySFP0ogE
TL7mlodgcCqOwcWnfl3IY3iZNSIukqaXPvFQ0+J/HNlj+2kdU6jYj3xUhT/CvzlRLuNJYZhB9KY7
fTrqLJG8LjkvKobdcZY9sBqJPPfSm8wQJ07WqxHcgsjVPMlPDXgwuI03lLcIfjbcQWHwgEjJN/yX
8CUPbOobjZ2p1uzdjd5vzeGrEuuLGsSbqPF1kOJalPQwv4B9st3iriAwEoqYjwsfPM6haM0i+QJm
smKbgNRtIbAs2rl57uhW25bwwXXCRALNgTSvKL04TBepSd93D2Ir00e0MyT9f/QJr6e0YTgRAmg3
OXbKqDQDQk+38eKNrLti98AjjOUVdRs34iy1cbrWKS5iBVqFRhvKUT/N0NQhjimTD/VLMuQPVpLN
ejkgbEzHwfjyrPW0Or4e0RenUE0PIE0PNmm6+3C0cgMnu09snz4mKo6oBdEcRkaL62VneqIXBYZd
x9DBNsj49ht/x4R94cYMoGPJollbQoMA8KQqH0iIW677J/Zd/27ZcvdMQaBho+rD21LrJqAOgfI+
8B4DE/oO3/nxVbzZsDi46iy5epX0tXMdDwcxrIecR5nKeFxQ7+yxpX2oFv3jRgGWlf/AZKe0LNAy
LrnRsHeIcikypmPiUOEGSS1Lycw/jvvv+v8ToPwEUW51c0So/6pk9d10lLybfsM4XkLHF0Hb+D3G
tthtqL+mDQXdvnxQ/Ri48T1CmzdXijai3/yEjSk+h7C2gTemvIcoQhfD7LloomBXv+2RGAP65Q4/
lLQBWhES08r/nV1t5bHvq1UD7tWktcGjSkhVMLxUFmnLJK6COhUvTceMzhNl7BUjjVfVClgvtydL
1MG3X1gPmbnvtdUlp3W/XA1RAilyPLRBI12aiTroO6JXEn6OAAtnZ8Ap+vZDe0Cb6dg00HkBW5ru
6MZE6tVKWrpcDVWzJJhjxChrRWbxZ+2Oy7Cf8/+M2iZ4Pwu4MSH5JmzV2nC0wusSl5Q6vOs9hoLL
2HquxO6FBxiQZGDWeowPCaO9FtXGBZ/pq6Yxjf7COy5FK0xYmdDr2A4ZtY+F0TD9yGDJd2Po5Xeg
vqXzA1qHduexfZE9uWaupsLZ7ZLd8vBn0bSAkjPaEpUrUuY43ViGXb3QBd0y5yYRD0hiTMlVzCvL
q0pJMbq3+Xh6hvKzJLCBRLnqg0g+F1TXOWuwB4p05m+k72dbEiWSrGd8wzpkbuYi150tSjtkWbro
M3Gg/W9/fwlCF/WUC5C0HtfGqySW+N3qcvn4DRzvZrBEaoncv70q54BkbkKSj8V21TyI+M0+HFXd
R4ucjudpvH6EijlJzKJ++5jQaoEkFVNhfUY0Q6zez5+jBn+LGY8bmnXS8jUYeLuYuproxneZQDLW
yRdHsNPcfh3Jt26Lg4IFpAsdsKn2UPSoqR4essqDWpqx5ZQXrkciuyW1TX5gtiDEYw9WD0/4XNJX
iRjOGLYbh9cHgIb7oUt/Si9WUp8QJ7QzThW61nZh0DfKplxTq364/cawj7GoX4FvGe4FoqGncOUX
ILkVeOAFldfv5q/v/GxAS+qvegrzPK4rogXW9G82SUD32PGHlt1ill/IA+2E0pEiBWkT4QWgIHSA
3rcRzRCG92bztUEYYMy+kErjcyWfehwpYZmGlbYDsN8mnU7miWEXEtjg4VYegwi7M3gr6ntp3Odb
cYb5MMUAP6vM78Ya4IFE03hmNg+gAtOkj9NVmj5IqP2PutVbnacAhTM8MCKSsumZuKHuU9UEwOq3
Z8ZDvdw78IeQP5Z0Z7srLlgN8n8fRVzhJKMKC6Kn45ob0BhZ1ws6ex81thGZJRlTNIl+UAKcEUgA
6jLJuRobOi/goUp7I2TuW/j4xUAU7HuNCKcX7iy/C3oGV56K8EuEhdq0nQuFl4DOwMO3UepuevqS
mT0uCxEgPa2zrsavZgo5brFJxiU/24QWe1ZKxvKup7PI45TNxz8F5IbH2DtVQ4gis3NDSTrz0s2F
ntz1Bm0Zx2STPguPPGjA/9Xomf0ZhkdLNNFHYKlavYUEznUrvzeOs+a2Q4/JTJVxlHj91Z+PydVx
cZSmsoZUIFsL3bkfCs2M0GTX1N3wnMxvT1mzWrkokmWEOEiJyjEmYHNOvd5Q8VMzesynJnlYEoDX
wtEBsA77jBUTr3FHrSJiVx4bCffj3ruueSDSozStQSN+GM5SbKy4OO+3hQfUYb38kTMSpKAusaNl
jLsbKziJ5j/bk36hqTVC/iejBXmCCb7+cxVhKjbu7oDPXCOWYVtXMYmhzGN1VdcCzT1gBVr7SJS0
N7EHJZEcdaQC69DiCUl6oWfhL2jT1VHSfcMDkiQRzNkYjKTGvjdMIXTQdrIiscf2nBsFb/2cqY5G
9jdxCpAWxtGxmGxKu/Z7dAl5tEoOmwNahyRdMUbyxPNNG3mYT8fs9/cLo/OIDWGeyiQ9gnYmaEmE
J490p6FVF/2IifHcvUMOF4Of92pVzWfD+i6hsLkk2aYEzA/5/O6zFdAc3C7Kj1GEC6l5ob3a/DGq
qUSwgaYlRRP3PRYw7ELoUz0sR3rTCDK6MXW6L5LwDefWPAZ+SLEnqDmIrMUUMeUKFtkskH8mt0/L
x46SPrHvBB+IuhyZtxt3c3ivzyMdu8IVAVWvaNYTrYLhfE+8F2/cFwOmCkdUQSJo3ww0o8LnaqEi
AuIm8h6FtisdOQ8XxxIZZqroNwws0wpcqG1BMYDsPMHjSd2n+qO1uhjx3HooxGnGdtaUxTexo+KX
FMLaoqYJMLlFPTAt7p3niYqrXcwiVOwLS7djUZwNvCjKp4ynwKLj0y3j0YJfWZgjI780h8R8hpF8
nsK1Yy6Q3XR3bC+UGbjcHJWCLHC+0s09k63ITJvx1BSdxHsfPEAd0DiBu9HGNvJomEvaHJUpA4Ra
FhxmaIW61pRmjohR15OxFZNUwq7PsSFfr1b1BHZ3maE/bobDJ7zq6YhcIueaM2+2ZP3F3g3m3LXR
gGQGFv0h3A1jBn9SXhZLVLS9r1r7hzzmjLol3iYnt+bT2CPwQ3iYPxW+QUXJQbAaxTZqnMMx9nab
GK8FYSvNwpGr9nazn/AerrF06Cwx10v5SKsrrsrK4+OUm38jhKp5ngq4VJc8K+N2Sf9ni2D7kIv8
JGZcGBM+yfZFKGobb3lMvSoXWZ4dYIKCpfzeLkOopGCf6XjMMBbwEYVMGj5hTT2u9XcN8+agquRT
iOaZHZ46dUR6SPBqCcP8ad520pMxhh25KL7BKYd5mcjYMQudH+WK4dKXFL/gS78OfIsX5NTApOkK
FqcOircLfN6KtL3WpVLIr4yVLFl2vLZ0utOvUs1Xggq1Cn3QZQhdcS2gd5/45koCEgFgeYIQ285I
9GJa4yM1wAOKt7Xcf6aVTEW53meGoIumtnWCjXnt7QzfkglZ4aW3ryjgUFAwROiPEyFqgVJx4WKV
UAbjXG+DosZUK2rFFZ5ZtXKg4NG2jB4jw9g4G/9F1aHt8M3VMLIZeEUyi1T0/fFzMPaeeUVaRg73
8x+olM0sVa86jttbq+J5PR3CzxLb8MJi8VF3rkCdB2yK5bthNsv8/btpRjulOl5z4rDaDccqh2rH
QHPaLc3z/vFl5txB7V17FWbmFYhJbnJnZhtb6FeBlUF/vUhES1UEhSOC073pePsxR6KVFO0TBkSf
FriypZd8Kthh6kCq4PJ53ftnZ/aBnJ71to+FHiFHxgrbnhT8KYY7UfwaIDq25iiyx/lTductM1vp
Zqdc1YouNj9u2ubhkh+dBsiyPgqkEKjZw6yS0iL8koIMoBEvaVf1hXQJkddTyIxJa6HpAVEK8bM4
VGY7uC/8RHQ1WVc4Ey/Z/uixM2m8M+puV0TMe62DWpcO6HT9jRDHy07GT0051zOm4xtIKQd+Fal3
Ev/IQTzme3oDv5/teIzYZTqzQ6VINtrCnjboM3ruFKC4qq+dGPotCcoKa+EyeDSz4yUgHzUZudE3
hK3BNQYhvqd1T9bqQTzimY+MUiil+CAJznsWmB8uJhDEJcjK6nW0Q4by1O+cSfxvVqyWIFVPXI1Y
JU08+zqseGrJ+mo8JLriomT1h2fXCJt6zMISFK+Z5tGlqzM66FljDuZA+kLwfP16UnP2p6H+/96x
XGUWrC8AMClqxVLijchUCbCE4gCqW7hxtyfemCscOwRH55OxAJ5YeGBUJMngCughTGEVRUTgipLR
ZGR3daNnDVnSgLOmxKCuxAu6zRttmEAShG6VvrUikO/bneU9TAnRec1EkToqdnPKyekkUYIzKRh1
g8ays5YxwGHvPKzYmBdlQSgVQP55ZbrLEWMjZLKuymp9jybRFVo3oKZVhbMW8Mx4ii45nbucgxn3
b80Nm8jjHnPNWjBa2gZ7KGqa6Lxkohba4iU1AeQTeZjcSx6dkiS3DYhwrs90fXnf1W7ST9Ki5Ytl
biaJbzRzOoIER+hbBOXWUklPMC0etMxGoWEjWfvVNM0PIGD2O1PuO5KGlN06nNbjDiL+W3qTtiSb
Nfl/rsE8PuQVJdHA+RcTP/uhPl4Sf71i6UtXXCOKkp05cOvGPPp73/4wiTF7TReZtDrRfbILcPmZ
eWKoXHOl5rw2HFVURRg93SJCxhOYPnYQju1itcWApo8V3qEm8OlUKp4oeKOcK4dyhpiAz+2KqLQO
iaAPYSOfLGjVTRfPo+Xb39pXC5/CkZPFDG+vLqFX106ZE20vUsHfNAweukdofGgTF/+5rDuMZlZP
JBLbvLQGeOX4IV33z+G3x0+QIAAzlRq7628Dp4ZFXeLbelQyMbQWCizIO/w12SAAcw0e1isLecUZ
EpjyFe+Wo+pR8nQz5d8ktx3/3eBkOsXtvSKYtWOTtjN3zg2MnPhtOD4FCrMQY7RBURm1vR7HlvuK
ZeJwq7AyEiY1063Kzj+OlN0OnYA6Om+Lb5PwbrCSQOiuLxNc15jM/prMu8jFzy0uVJ8NNx94hM5y
lUv9aD6dt5PlBSI/hdiVGqEsv2/GsoiQmy01/1hJ9HXxb1mz3qPerBTd12n2ztftWamRod5IEtn3
0MGA6zzcMIApzW8vTWNQqFGakJjTEcSaCyuT8yOk/NIAQAE5tiVdCHRrbtdOeQZJKWehaDz5vxN1
SUKqp/YEVq+ITGluEl+PSQLg5Ws9CttkuNZM9EtTe9xCSlhi9H4DbKWcQLD8hGFbcPk5sVtAcXrw
SWQlRG8e6cfU5IHCRwth9gtPIKUYBMN61uyP5BhbaJxf+cfVrvxofODar/3h/Z/FhgVOI6Nn16Lq
Qi5R/h4fw0Lqi4pCJBql17nw/UlwZoRe4NpUPS0D0zsm6ssmkEX7s3dshFXRrvMHNvfglv3Ljxct
kkkU8AeMVWgwHngOXR5mhGC2OsAiryEX0Qc3TN0YnvMILAUqvp9wqHFya6hYAW0QpyhgC51FXxzZ
OFls/ovmvfLkTk+l/tLA4AReHum6Bfd4wLlv5C+LccxgC+JOElotsjImtJO/BuZxWuvB3Ebq4BB9
8z8BQ3PY1PxFjOTdwwQbezZOGr2h3/z3RkiLzINttaCNIcVPVo9rDB+2/OiE6AG9f3eYLrgHJWQs
k3/xu/z1VCjtLb+oQzfioOs5SpDZ+4w/bXHhstt5n+5V9sxDukvSD+7cWOJFaoi+hPj0zu2l/Pjs
WYBCSMq0QT/tjyq6LaRuDfqaAkbzsjfzvHcfb2bG0Qm7ng8RGN7ZSVtHyk1WdsfqSE/Gha8HhJAS
VwSUiIav/CIdYKCFt10GabWtRFI5NHLwFkcgugdfN20GOIQ3RYKPbbroUMJRBKCXX/8hfncUfNVt
5a0Gm7RL1CXmMjUKNaxaoZvp2WUKHxMm9t107681Jzaz3WJagQURLX2V09pDvegerGThHAw5hdSg
hf0ed5xDV8u5sue+lNVsqw8pZxS/ocUQKdnBJtFO9i4lOgjlZDBmZlhpb50QHJXPwrw9rFqN+Voy
mxChitb7d+UcRyPNl1x7uQfgKL5bPh8RJJpx1fMOqhd6iuSB0Zqn8gDnkSV+G9DRbUZWUWWLdhvw
EeYmEQZU63KrvgX8Le+KAMU2buA90h/JnkbBpp2e+0D1YAbjXszkCSRRDIlgQSdDqeERNAj2UPrM
bV2K1nS4UKNe6Nc0+0Lxrmbm1TlEezGolmmNMgbN3BP4WLTaGTkmFpTL8r7h0l3oXYDjti3w0cZK
LDUllSw4xwU+qFZXTVVvVWBuydbGDPa1OAmLMOSoU3OEn4RxCPKbq5YazaCFWtHA9+wgOSBoBjEw
4sndnhbxX5MuWxMSdYJzqOLXQKDro0FB6BGmU7gHjU85cqbalGpQLHVZ/mEI4pK9FrQTsDHZQeBZ
/u7GCObqGZ5f62FuniRe5/V5ontLF/9k+S4AigyZYgtAo/fFu9SLHB+D5vAg1Dbcoijnm6Y5yDIE
1r9cbkmn/5FTzPB7Z86tmicrZIc4A0kEwfbVGLGx1FkOqaIKPO0Zlv5kkhmNRiVS/K0cs5nkELbm
0yNvHz4wRizBnvfPu/n/fR9YgulXeSIwLdX8kjGACX2ifN6PaXBJuOR/P3ZBA9ezpfpt13uK83GC
4uH5Rk48fbTmoTF24qk0BKJ58GChUpy+psK6VqS1fHHrxhKthx9pvoVUduab2UtMRS5nIiKWLOkp
XvzzENhjgLGIgpLxDoeZxn5MBfnEUmmEgfW55DrwID49pjyfu9yqLeYRKtXCnUXUbh2aGnaQ3QyB
G1HkLQYglEaDLW15LN2Oj1pX/Q31b2k4amKuuxLOszXPTMQLIB2M9HokWvaEKck5FaWI2wIheGlM
n0F5HCT0KDFXSnpDUuvGp6oHkJz6fm9T+/If4bturL+ARI35EjHuuZqieh425Z8+4ZRWkVM5YAoj
PL/er/Vt1wJufyi9GmtodlpeR7HtuPTR6pQXh1GJn7VwKVpxQNF/ARTMZVdLTOQ300nwSE4UwBar
xtMUeBSKwnX57C7NiU1ix6zp/nt8txkVOOdBTCE5TCj+cofkpcCW7vVduPxBR2ykbI4y6QdlZowX
lh3vrKUPmB8pxlYBRY61nDWvry1TsKpl8CjFRfRmOtiEKJYVv9fKP1egK6wKmXbaUjJiiq1F/Uir
snx84CxGTecPrPmLM+nR+f1EGgszE2JlM+ttU/IwtqvvUg5oDEsCcJn02oRhbun3whFM5RQq/Qrs
Rl0+dynq+6W3/QbcfxToXFrq5bhIY7Pkslxb2m54u/oVd1as2NmdtlBHYL541IMnJiz/qcDi4FFT
i4qUcKoa4q3/c9ZFWNoSH6K89RAX7+UtNj+V5nYVLrvTro5E9OUOPOb0d8kP73nKJGwHIV165bhO
gW7xIitI6LepybQu0Zn5yrSqgB66ulg0NVdE7hGDeIxYnjyr7hEx+ia4H80jbdpLhm+iKCko3Jvx
BBKo+Gg0kX5JWowpzxsdBGYaZyRDNz2k3yiU5VtuHbUw5PohhyEUTJpyoZYlAJhBB/L/EOWt0iEj
EZwy8m/h1XeuAbJeMSHSZr12JuhhXYYZtFnVwaBij7B/I/iOqzNqGzwwAhkoG7yCojETHhXM/Pik
JVgFN22E8/rDr4aq3HfNDIqUgw0Uker7576RPeDhZX230l6Hb4jf9AvQnU9tH93MQuYUVao2uHdd
WnlFfJdMjAVtaHsSwuE3II6l7ePGmss9BfwYpTOc4BvHY3YaYFGWmeeKaLbhfTBlmtU+VSa353G8
RtDSVQZfaZHWyptpPIw/obQn7fS4EZne2MCKP1Hkz59Z5vy3gkJpRm1FcC3HfLsM7faBTBpMhTpz
eH6vEb07XN3Puh5JUlEHQ9QfsxlgYwYRMJhI5WMwK4grQTD/iTuH8VQMhPJuTMAS5Ip8Fklli5x7
4Q2s2RshpjdJIN/nZKQrcV8DP2CS8EuXj3J/sW1GLbCTqCrE4emPslPYCpY7IHFLnYnBz8KT4mf2
u2RcPTRHBPptf49Da5hzf3JocF8hJ7K+mzLV+XEA5CGLkQEb47ktJtja9H8ecR+g1Z0ome7rgKfe
4GNnRDm/ZldwSP1hh3cPcUK38MH85RJtCqlPfCv4feZQUc8c/jNj+JRZjbuQOc4xA6kxpNHpMLhY
0KAFxKaHo9KBOj+7RFMA8GEL7jllpW+A+HpatT5RnNeWdX4iFWVcVHnrxghJwFTFTjDiFgBUg6yZ
0BvQ2L1+QbJR51ykWqKNVIcHF1Tg54vrGZPmNjDxQOejSu6SWsS2VWP8hNEMdInWk0ARyFl8/S4E
/NV795+IZIZy/hUe0gCak0XMV04EmeIAI8ONPNOHp9jtI7hqzAnB9PK2OXaC0Pg0dRalo0EGmRQ+
zLXug6lWxDnZJHU/KTOl0vSZvG0hNe8Qp9mHa8ga5QXBqjdmwpMRvYe0UU/kFrDNpQx5TFHXkKBT
tDS4vsYVjh1y/iAmCMQr+C7jMQYnoWV+X1TRdqAqmQzxyxDFhldgWmxTQfjW9id8pyipIefKuD56
LlBfTGfD8h4b75HfwGAcuWre7SRKAd4aZzkNeGi0rJbCwQLapN17Y/SNRKH9pSMIeUmDaAyA+dj4
m02icVY/soKA0KzbHM6WWk7GfOhjmLcsgsnQ4Y5vkFCv42J+Mu1czYN1AVpZDdcTL5hN5T2qjp+7
wAXlxnFop6vcDa8AaRQzGiNwGDdWVI3Uzu55fYDhieYTVNMcsQqEhiqK6yvREhPy81sQwnuWO7GS
iFc6LN4wP7tqMPAZ4jrJKd2MEDALnSIE8xMqycodvFLagrmLlsxdB4Y0Zxosic5PgSbkc0fvFwqy
HXQNiPkMrxXRBPsOkxDBgCX6H0XorXuYNfOQ3kd8gySgVmyQ9cjaBnHDRiPuC7fSachTO9iLE+lm
D35b7o9pca7HlpTg7gflkRAH6xdcqUrqw0ZtfBRifSWUQa1ATQ0wKolFierfRl5CjVJVbuqmzXzu
zoqrMw0FcN+QfQ76BK8RFdLxzjoSdLpLEzOJyAUcw/+FR585dVO5W26Jc5yXxu01F+GUjd4hlpd0
jCtizoVkhT2brerCUoa2ikW5fF+QFhiD+M7SqNjTNd7P3JYsBt7zLGxvWGlejBKYSGGA35iZHYI4
v/p6Q6rKI7phliCg2tQ7umpXgeSp4NH6HE4odyKj6Y3Vla7bJxYffruzs1nsiARooQsJDQxVrwkS
5Mw9VjNHSWeNtZ7Kj8gQeoFc7miKwOpEBWHHuRqf08rGNE6IpZMUtCcfdxwSY2arwrULyn7jWOMA
inmSgH9YUABrLTYEpLih70eZmOBlCRoRrLqPmk4qT6Mltta7d/b16uf1hSTv+GfkKC789NVicJL4
hFmvuoxMGhd17DkEdvpIErA/+1BVNdleRsKY9ZEFt9INK7PVcDda8EpOEbmyNJnbwCwboXvVuJ6+
WKfgYkwr2BOM/TrPVh6yAhz+vdVU+nCYpx1AmwUHW1/k3Zuf0gTk1DRZJD6jJn4xVUxliZO1Zs6M
c35rzssysec+/lE9y1988p3IG5h8+89BbMl/Zv7dKne1xzVSdIpoGMgeq5q5ZvXxwp+d6LBaxcqE
rQS2f8Pl59n4YpYWOqxxSdk1dT2MJjZUsO/nAblDUzl8gcjdq1wpdfA0VV9YOF3kRafVxT6fSuYt
jNN84IZR1gUhGxvcWXbsi/1tbJmHrIqTcNCjqy2kWni5MaRw8fEi6LM/GqIdXtTBJ5/4okFurPoh
yI82YqwPR+pm1yYpnwz67TnpQ/YVBsOGT5BEibwC7Hl1fFR5W6psZyoFA8kGCfobZxJF24KoMQGy
2qPvy3TmxCWDL5mDJ9yfOLp1WJLrlOgy3WYrS9koJS/abtIqol1WMCKlbdwYqyM4iPIbVjbf2M9L
ZuBll+CZb2a67/sh42Xv53uMFwh7IwqLWtKWDxWgFt2mbcz3qDBRabdk1F8TmF0nuDcrHJz+4l8a
vPGWHdzA8Y1LQuvWHBaGLc7dpJNKudgaZCLlPm2lqAdkcxZmDetlGDkYRtCDibr/+d3qEXjklfO4
5T9eNyD8/LiaF+C0OPNzM7CDrGlXGaxcr5zok9C4Fh3dh4Tsku4EdQwFKA/UNEi3q7VA5IyIbhFM
DmoCHQ+MMJy6cLTaxlRpeQaHIk1aB1yAiN+6VYUgo800Q087i5kPyJzfu505xohdCvSczxEwlab4
fnsawSh1ifRmVFC8SCOpdDHADJ5Mv8ISD0idWAmQsggL6mk23NWWQpRO+LQ1vKOz76MLTc7PTwpz
+C6cGrxBRjhXaud3lPX7U+/DMKf+PtTZmBChjXYpzhMiGabl0sWqCj90X7LO2g1dFFpp2InQ9ssc
xSpviZmYQ+Ahaqh0SHSUvIuV9AG4rYQBJYe6tQDKEbxWt8c+jU/rA6276/rlU8QervJO3UgA10J5
DfXxXdGZNNz0jvFEYPAZjwCnQ33DvvN97ETDs+0gUy7NbqYlMdmtmmrFAIXmYQGmaYTR7RHpxJYD
drofJByLWYfwKW1+rdPJMw24BM238r01ErDHNyJQyur/AhsP18GNqxIETmgiS2uyF2LaRhIOCU1C
X/XtfOIik1aPdwnUBEc9h2etUHUPyHBMSsFfG3wENklHaa/ESjvIgD/zJWPISCmkZheo+e3uRvnf
kjHCpzp5a4oikT8NrZZYpZHEA9n5e5n/7eV9ZpGaXMIu4DAN+Qgzj9NiZywdEWAfnLFUErLlt3sJ
O8mWmw8ZVmunvlHAercc08SYWo+JjIQOnx2eo2yR2zo4ME7u6VlW3aoNiys8KKDRfFCgAaCJxYb/
FRnUe/kWmiL2GjWjlcl+JC7k6mbe5eB2AbVI8N+ahei1p/dLps0JKmN8TDSiSYrKiL4PGaVcQFpK
756hwuKaIPciunJHuZulvfH/v26ZubxvsluA3XUi3cRX/NZNCe15lq4QROJCxqwevB2Aglt/fw+W
xXzwwRHyDOxOA5gKulUpX7ibW7Cq+/j06C0kgPhF57wuOO7Nt53mgDear9eiQclqIj77f5vkpy2R
bDj1gwYixwoVENA0dNhPioll55cEz1jD1ibwNEEAKPW+2/toZDASaaUA5DQrkA5+9Nh07meFJXRz
r2620DgUlXmicib1muJYmOQtaGObLzWSoNFvI2OzOVw3xdLs4SX1/IXh/M+pqepDJzHPunO/0ieT
HyWByjlR0u3xWN+TV7RQ6dQzbVDKdAvGAvtVJQkuP7Vn4Po91bh2jlaD/i5oMbKn74PMgczlWtFz
7SZFD5NzygqTD6ZkhjOi/UESbyT0hjDsCdy/BVLXHn7aFb8kfISwUbLfl0weM3jMwshzYmVkd8Bj
q0JLSgRlY+2xdcfY9zlsoJpTGRsxceqp9n86ptGPttDoCz5vLUtN50vWgtHmHAsL9WljI7Biwnfa
vQ9VYtpBlpkpjJuN7d4BhIn3KB4qgiitifjTDYwSxDx9d1u3Kvh+Nbg6to2rJ/oF4l0h5yzeH5px
SoVpWy7gZI8od6VPG53trmln6fNpF6ucKHC2hAl/YryGxC8jfdwQxgo1uWeuMk5vzXMwDhfrudtb
okVLyNZo5zTrUQcA5xx2bqvKoijhRU8G2WLlH6akQ9jCoiOEaFAAV2XA7KhVTXLr0+NArgz5uHt0
53AWjcyCv9zBOTvtdhUFeLG58xIIEELviZo6CcfTusDEsM8v/jBW+K8CR9Bg1Q+JwsxmpAfeHU1l
Xo11ARvc4tT86cyAhCm0AwB+nsKpTwVoIX/w0SOKL7Eut/8yPScz4+h2x2GylWQnbbLV8FxwMQvq
8LE6vKOp6MUrWMKIOMqArYhFN1hlluSbCn2uSYxwv8Zu5qySk63BZRLgCSeomfigp8kZOoBshJ/b
hlejGCoNa6DpJFErEfomz8XvsmoVlLbEibu6LaUsTDvIwDsTK/Pm4ihGKHo8SmAGpZER7cCu895y
L5ylMl6vZrN+EY55C4Agkh/4Y/9vBCSIjvN6PkMrU+KuXtk54zRODhA39H4BqHmy8VmzRhhB/nyl
M6mIFLm0hMUXLRTBFMrjGBPzni7tWh1KyYYj/AsxBrP6oys6nIVCLUssewQ6fL/GHD6RWcCJ3wDx
BSNRuFddxmsrYvBvpiMfBXFnfzez4mabbiwxacmeVs+FjSM8wwGF1VOHwqSJaL0AgwMUfHcMaHKW
qpfKFn8Jq/YLPKyis4VJ/bPmpGS5/yRIAnFZmagnrhsB7UoZ1EfynnE248YK91M206gUvSJ/HgLH
Gg42WyjLRMfSsHwuFc4LOn894v6lJ0zKQrYOtXbYPnDQSLJzyjFpZRDSPbzXmcZw3ePFBYDIUPmP
hCJQI2/TGwEO9lSrTo3WT2ZDFCGzwRxjJ+UWgA3ROPZmTaGNt1DDKEOzqHfTel849KB4mnIu11Tb
Zw+D+4cTCCWySIRA+lW8wijKGsOpIag/pU5FHJ6XGvEZsPiJyoviPm9anrB5awl6kw0YM5URvGyV
8ZYl9cYZo+Qa2f6+qwZKUFPBH7Fc/XZKF4NXljSSx0w8eQKNz4qxGVk32zSAkUKiWzGLBMdxNuWq
2kArFpPqQTkBlyQXThims7oCMKHJPq2iv+E5heRTNUUG9KoHMd99j8KZHq4vlIbaI6tPatuuF+uQ
6F8JR5bnVK3vQoEpAJi6V4iyndgJ9zHI+0fe9vhh5db5WSy54a1TLseMtgRedhFp/H0S4A7Noc7N
PbvGVq4i7NCwu8Vm46K6dYFFb2umW8gQGdqK1ryBCOJ8Om/OeQidz1EDCbDs8ce7BVn4JxOlycfw
+i02t4hl2mnjh/VJsesjBt5af/TmluAH2jifLVEXj7ry80PNYlikFw/jgKib0IymTPEuLGY5V5xC
Xba3lwOecNP0QtgspEL5HLXpmQc0BR2onM4kCTeccxmVwgAr+7gmrpnU5Kma3Cv/PNv4RsCcMIwu
ZzDzBv7uYDN/e75Sg3625WuRMkjt2aNva1lqw+IodnD4siFuNmHMFsCwr+hYXoGugIU6QygHJ6uR
Xz0B+qkblWxmvUAKdLyFHxRWgYGG6Q2d2VtTPF0HHKBZcpjXb4DUjsXp5vDIiAZpVPVRr0gKLsAF
VcKJRteFOjAiv5WRcmQXcoi8V0wOg4DzsIt7Ma8veggroth5bzzsMh+ppgVSoPVlmeFzQV7jO9h6
ztHEyWVt/QNsrsUpAgwFtjyaQv3ez+ElIRxMKqdgpOslGzDqa9M47BR4O0FUXPSn7ILE/muFWhos
vGJkCgy77oHbhoMlH41tnkMegAAmmf8kNQZdxjbKI4qq0hoJ4JR5NUpJywJywu8QPDi+Z4u297xo
xhf3+1kAyfwMDxmBeFTVjEdAsBz8TzHkongCD/dwy2TnRrbvpwijOxxhKIXZRapnqF5Y8SjTW3K9
hB3A4ivtBqhpfL4zlgDSwdk4shtxUcfkegZkHCFHlpTR5xH6EUPdqhMGba02A/QjHBtbF2813M1z
dER/8iZsbN7Ah04cA5GbSjpfRa8OQCdEPaiwypNo2uS0JIG+FIoJJ5ttbbE2NwGxKwYwZNcR7R1q
2JJ/P2Ruz8OoroRxRHsd3ifpQl0SEVB/2wCDThsHk2389pklXAOwwvDkvD6Gbx0KXwuFlu0NlTFL
wS5ZX8XcBXzgfdxub01aIdipwwLkURHBG3p6e2jNKO23FAjET4TzXfCYctyBbcjp8hJm/Yd9U7qX
7pT2NAmMMCjxgiz/cjGucSZc3wDb1ppPMdX+kIA8j5axXUl1Zprt0U6DjDlPmO6SklrA3JXCovZ2
TP0YwWsU2zbYwasfZ2oT87FEVn8p96uB0ZADtx755CA5P5GccMan8+hrQhGeBztHTgvP6FWm5IhA
M1X1xhc4RToliCy6frSLcFC19xSMvOFtO7LTvok/YOgkWhUNcR2674GaOCsq42NMiwBNVjyPowq2
5+sODn0q36ZG2/bKXG386IzhQN2srFWbypVMRZOrsclTfN7cssu80MznE4yWyNs5DAEZ4fqAvWPI
xwpBZFXMjaciXg9x6SruJNZrO9Lk4tccklJvpFQv6QI52QfT292f6mJvlKthS4vEqMWm/0xKpTlq
yNxtIW9TD/XYts7kRcTZFDOdlohzHQA1jdG7KjJyC74nab8YfrMMK9pWfDSQaWECReWGyV7qHUdI
aRmY0ZJGRaTUEqL7yEZF9B7UOPolBtmqFSKKHzRTJ0LW4PE7u0tWSyJ8hmXcz39DVyWh/rt7EmdH
HHl232sf4PtgzbQ1bIcirROoCxrPOAaaM6MWye0ECrvssXVgWydQvm9UY1gSzKuy/KIjVjirDgR5
d/hjNBm4hpPgo5nt55ft5pn+tN/TFt+N6+fSCrMv7ztwiLatu3UxUhjkQ1581QQzqR79a5I0wkBn
0IZzybk6+d2XlGZj9WsIk7HCnlZFSaRVWt65DKwJhw50oO/22OnLriRgDLU+4JalT/ntNGVZp1fi
SbjqdN3DnWv8vOOgqFuLIVE6/S8TsaSafMCBLWGsa8eT/rUPHdU15QAEWXZwXo0GECq7960kJjv6
QMp9KXEo/GAdrGvmn/KQ5LiTTrfBjsfIwjKYk6J9CCQ3QmkYjY0O0SqO+QgpJeK3sGcvRbhsJtMv
qB/BcOG+z8u6CynpoposmNYpgBz3k/QEgI69Wdr/WCcgvv9YoH+nL1opShOwazE9lFtb8AKjb4WD
0aprqcIzIMwVe4k4ilu3qam5j9pcpAL5xQt910oqKahaEaME8C3EcEs2V/zeO18GB74b09ppBRE8
m+5ZTMRKgu9ehaeemgPxuxaQPxsqhsLzaulaRiERGquvx73+vvbbRvfj13SvUDPpZFMDSHl0fdvC
e4Tz8ZUnjxI122r8FwaR6fH7nSWBmajPSbiydD8JUhEyfm6XPgf7fbZJ3xR1F4ee3LpMxLdFFlw5
2Ywz4qp4AyLdo2ctnUVkrYvjd9MazbfSfXzjWBmpxZHp2jzO2jSUj0Lb9JKmQL15KtJ2IPvXW4LQ
wkxlhBENjYv033c9y0P2JZg3v1w2+pmWTLLgtTUOzBj01HHkSp/O9FSadDUocFap3oNafyFxVAho
M6eYw+rxzdq9b1jwfmM8MhuSd+3mHbwkXBWqsF5Wt6wx14LraH4TnQTlsbaG3hNYp8OXCMPjfXmW
0pC81PIfdiWMaKmRtDppbDo61QscCMDHnZsVwATTwOJxVZBZn1Q+9M6gkSUOWIKH0/3UUP5D9m86
D8FEn37nWwD9jqaMtVHUNz8JnUyLaajnm8rjNUr9u+NfWGN6UF/Rx5IQV1VlAV82/4oisMDWoVVd
gbTWIzaa4np9ywsUHaTOpHNbQsEEKhTjUP6kl5NlZti2nlTC74Z59CUKrlxqcJdv49WkLF92yVcP
vye4QEsgwboc+jMZkufLD+xfGbfGVoK0eysXmjbv6vnOfZ5tiG3XNiExStel2z2MjNx1sunqPMxq
Fkut9jYiq2Ih0EshZSYYzspaNdhnRTuhoOaeZ0Uc9ka6l2DnRzMLEiqBFLzOeuX6R5rrmgk4zAwJ
YuQxbOvf87Pipyq1laNDbQW0tnG1u0WdTrg/jyUrL81WZXeGP0VjK7Bxp6+Ogw+sfojRpJe0XNP3
KkumEJdAtjJsonGeXkuwfmIjxtXgeomzkAJBB/77bIhRy5Nf7wWfR9074pRxi9zneZES3U7MCOv6
ayCCWDhqspam0g8wEryESwgijxIabt4/w8eUa3Hz37Z7uUSf0+oMRt5GwEwzpGhN5W5IBEaQBlnP
clxrfFBtQAmS+bM5fo4sjgSlsaMULKc53hgNiuh/FrOUq/tGCRuHJJ5jp7RbqJGg2IbIgZ4qEj7k
ov+xvvTIFoqp8T4QHGjKpixSmd4Rluu2gY85VGBwtEQLiK0MTtuvNXzCsyMUL+ROwcHQ4Ntap3Wu
I2Jix8o+QOoteeXqmTnoMt32WSPirhwzufru8V/8cAg/BLZlFxbyxd7aev+GjxhKnl3V1ZCy5ytz
fMz4sldzERO9slw+4tjf0PtDLJL9lyzp3l3Lf8xGby9n1FGFwqvAct3FfRTiH/vKpEfaUDPUtIp7
kT7qF4aR8kG/8xvOonF2avdXiQS0jyviUTMGSJEXbHXkcfAS1IbRHoxqz3+me47yJ18tauQpEyji
AD3wbypSk0iKLv41SvEaPdnWT5qXf2IH903fzDWo0B1124LrmhRsKy3Dpyujb2HJGOMqmoElfvNJ
vZBq9NCyAHKTXp6LlC13dQ74Dre7XkNJx4NevI+UXUT160OAZC0MeXWwt4NAnmxIXAOWIVwHeWXu
Io9rh7I8s78yGu3VzZhrujtkIvjyYuTr7egwX8rRmd35/AXJIgvDH5ixrI0Uc+gBFXMUY2WpKNvC
lohApXbjUXotCEf6oZ1DDZK/7Z+5lWbzWmOLtbYwg01Z1XiNA6BroiRv3qu7WtOzqG+RwsRfX+uR
LQLt8ZluRkSnwkbownq8L8YFltXD8EgS/MZZ/aAqPnRC4C5TM+cKYRjMbxRG8BPT+KdpSrHj20I9
p/UzwPh0Wf6GUp3UrEcGKbXbrdtdGb82XM6BG/WIiLGn/wZN19x1YSZ9k0wjbQoIf970eh0jJvts
GuxJIaZW5Z1bSP/Fu5YmOBIa6+jS6wFkLtEZODU8ufhmFVlIKm5+ddQ9LS4jOUfuPKTixQqqS+77
qx8JN0jhCiqmiySTWQlsDQpCxEKurdoojmtQEXBWTSlGrQdl2g1J5Dv6qVrd/At/g24eLhV9hjch
UT/u/sxbjPwuGo4L1XMpFfimMxzdMfSY82s08BShc1BwmJ10DkYucPKImjxHrGCvqjcJQ4viHwtF
RDQldpZwaXT1v0TTNogUA+FNl+7PZ1SMc08yPiPWdGL5t0M+/h2W3hbk8viG8fwE42tuyl3uTjr5
Y9j638ncxMgq7bUyoLTQc3eYavcCGFzufFV12EQHAiGtiz+NLmXUF3DM0xeGtBDKHQJYsy7VgLto
6nSoe+pVGTL99eemzXt/8oi9rGjtNU0d+EXurRxVdbMvul13n/iE8b7oWJ7wwAFXNsYu48ctIh3V
p8XU7kb9YyZ5uOWVi8dxmeGK/my+oyVsYrIh3UcY8dhNC2HOl3F7SWKYg847lEKjD5DS5mdCmBM/
WcG/KfNWcue/KVMgxLv9cgDTcEnYVwlJq1U6dRaBP6HlpXB1mc0yOmbtgBL1OB5VzJYATo6g94BW
gIMrWc7tc2kLI7xRHQMRNEBztnaJNRe00uWmy+K86eeZLKMcZft6bo0KYXjq92gOOJD1NBGXr0cK
/QS3iOw/7HmxPTYgmJB/Ly5OLzxnJWjt2BQ6SC0Koso6zo+t6NkRajKCAjtzO09BT0rci4zjrzUG
/LWDGa2D03IVb3Qo7Cz9qnJy0ZtQ5zQ63e+twOtGCjJwiSMFBRwi17abNd87miw9OXbDSWCK6nuW
N/UINSdvyOr0SlVXTWm+oSFqmcnaxIgJbAEdzcB+4S+tKCSbHW0ZAhTOEUaFTdcT1kYrlc7MMK1M
gwXTG5j4C2sfO/97GP8UVUFK//JnU5Zk3lIWBo0oCBrJZL8yH2IomAUkzQ1i+CDWvqZq0UPGP+Pp
xejnksUKXU3PnJF9SaJ3nMBQf4uq3RbNQbglM0EiYNB6Je4S0VRRybtDVGNMhecy45P8qvqE3wIW
TrGBKjutV5hK/nr2AEJZoBlD4tef+WAztQtyiZif5lPTM+VmQVFbQWqui4XKhH4ipcppIgYWs8kx
thB8onpnvc2qddnay+hU2RXcvmqwFIAuiT4zGo1CnNweVdbwjxI3ycHxaS71V9DpBwpVFhmh7OPV
q6bQMX1hh/qhm9iEgsJ1pxkYzXxFaBFVctXsXrUiz2Jk8j9Z/MV8uwWtyGa9p0F90vAWLWJnIF7/
zdBfl5EDtQ9SKomAyZaSA9JBbq7ijML7oUesh9GDqtlvH9PldABY6hZ5zmAI/z9b4LRNojAvI1PS
M0TQO3+NBBBo26g6Bg/3EKdUAxcAO3LvxvZMKaBQy9AvhO2RXupi3UXwHoM+8glp7nDwg1ysX+dW
qD9sJ46GmFQBxKc5Xa/OhgRGlib6Fs/zCtTwfzwZ7PBj5JWvH/ILMRmLSm7wcCR1ppygGcW11Lcd
+erSGqeznODM7X0EmishsbW09zuJ+81VrXPL9UKGcZ6yO4ADdzXVazS4X+DVgcAfWl4fPYYS1IrT
tYVedWzIKzFpbeOo4aoVkUc3txMNikeyruGAzFd1tAuYo1KELjg8wbwnpU3aiX8+j0DjI4ftJU3h
uFGUfsb5IMAP9yPsPjugL77Lv8lXBA1rxXnPD9VDYA/9C0GcCsHMOurteHGwEKl9pa6pGm8cirJq
TCTdL+ZG03Hqe4h64bt3wTCFk7DM0xJRFbKLL010+BR+KEle+TA7EeViLaOXTyeiovbiA4sg9kcL
2z90hOZjCIu8L1SC1T3WFZ+SYlo5PT5CSpJsL+6gbuC9mqVEclOdmadGbAsfSj8JuEkLgTKZCD6c
vN+YWRm4J2a59OAleBuG1xYT2APNznW3k7f+EHZyUtCdBDF/xlOixnoNFVU6vs7Hdeh8wJuJwVXj
U8CC74m2uOd3IvBoA1scSz5bHa22WOH3CHHSmTdQmFzSVbZn0xt+ao8u71sHaD7CgTdTSgq7HQC+
7gGC4Zr6HC/GvckqRpfPneasE3Tozkqy8pZ1EMSbVSzbF5lrCTmaVtgmoraG5CEULMHDOiSLWHdv
iFU1gFekfmf75w+rm6SqIdzo3v3B29O209MheYrpGej+rK6xmnludaFs7jMFpets2oaTgGI3zKhf
jLZ7k4bdEdznXui84wjemtYo/AbEeN1myo0dJPD9Pj6yrFMmSsTubTnzO/79svzSpmE+hRImhqbk
Vo47hactiWCJ7LYHoC+6e40amUjFxdGXPoQ6yiNv8nlLViwr7XzbDkjkcxrK1Nj7K6YFb4XFoHiW
bXKAuHJNn+d671j1EEANZUYOIROxbPsmJGPY2eyrEGQbiPAczhAkk84DCbNy1i/CpKMHs8KdOqOT
aao7/qJuytzobGvIKLDCq0URt+9Q95acnAnyPCihzvL/SUUSbc6xzCHQAqEWQehHC87pFFY407CX
EGdMEy07gheyYBOMINgOW3JdYRmxFjrpjd0v1SlCV4JHl4K/6O0aHNXsUHsTWsHAMjPcsBsCr2rq
gtg+FzMBlzPwogOu/yBZl3i0FFSnJaKTsS9fnIPCMh6BFItjJ0rShgNMvpFpcmvw8ANeV8r3LdJx
lBHY09aZDhBARndChFc//ba86bTxqdAVi0eSEoILH++uCUeq627c0pqYpUM+B8iT3IgajT4sF3ef
S8lDnUYV/8K6vcfwYO/m3bL4TXT78odKU30OhQ1I2kJK6rPAqRsTWrOfqUD0m5DEAb06+XTu2/u6
0hyqjQqB2iZhUVwYI9utfHGpmRp7gWQZU9c+jfh/drvbHAEXKEueEVy3ligimr6OphqVXuf+V/kQ
NqWAZuImSFZtFzI6983n2B0py17TzFtKP2tWM08DDg7ZVeDheiTVkVBSK3dKDcwfoeDsgLdqB1hQ
RJ1TmbLG0wPuKXPWevdfFuIalM6l5l7/CpakW+LQv6/Ce9U77W9O1zikEi0PhCnjZEztRxfq8t5L
y4Sxtrcc6KO6Alhjy373Ic2MoA1VYRf9gpwqwBJmBjMDsRi0aD5lDCdTaDJrizXbQ26rM8nDvgjK
Pyyc+t5E9sHt0rVko8sSDJn1alHyCkWEUWe0n8kx/hMzX+tJnEtqaTfzXxDKgbvVxjReIRC39GXr
E6fH4WUigwx0SCswANIB3aztycNYLpvdnTT6/f+MjQQv06wHnsmxU77pW+DAB8QT8PkyCnRVNA07
krUUuBoVNWVKPnlMImkqTWm7BwwFHyQs4Rp7IdDJwfOVC7DHnVpVL/bx4zvbXqQdbpTcRpZ4gY90
K6X24FTIYOWZmW5O1h7rFesAgzFvRxH8WlFWnGoVcIt5SMsStJjmdvW2Ff8w1ZxGw2/5zBKACua/
x1KsFgqg0hKgMJtH6hxjW/zGAtM9OM8/yOwiZWSZUncLXt2sHk/TVgdaNIsVlWGn86tFaeslOTep
rI8VFvvBNWdh/C/KvE+TE0IB9qyuPA24TlGCduQmFoPEUkL2waKfW2WuVLtshNQp7997HxiFsrD2
oxmR15tuUssgZ1QIC5vXN7E5S3iZz2MIgMAO1/mytqt1xwgfQ5zvu2cMrFtrQRcG7MDuY2BoD9ov
0vDZG6y6Z68W0ZoifTMoQQDy3Z8GHc3brudDd/aumnhR0qMC9IPtr8/tsIELHV9VcuF2Cu5zl5Y6
6fOOkVFQdDbNf+KVVv+la7GKlIodOAKX3kN1bZ17IPXs5DOCj9ctrEw2UU5wMazW2KRAY3GEFi5Q
4qZ7/LzAwpNNQJUfdRzcss5MoM5c0xKPBO+GCSOixq4oMHsZgP+undT9Z76ZVihQl3MgbJxMOZkY
nEPF6sUxhu4refEbVGBb0llD3Tz2f3ZHuGK6bf/PT2tRRLbr+HD/5URpgWeofTZbyydCJYecRK5+
3qq5rjk3gcSS0ypj9kj9O15YIh8oZDkn64E+2OevQKDjokUApmDIyZsIBaChpqZ6vMTYpwVNHr37
EbiYDa8j/8conaDGhS3aBU49WOExmCwNplS58LJQ9WNlbMPcPLxr642h2rYkgKyKaHJS7OVj9uwv
EYa538wKxSJyd7ZfIv1HXRltSQ9B+vbLuW8vI5985Zn/74OlFk2fYGvv+rj0/iNF439Dzrhl6X/R
zts+MyP9PImfcpGAQ3vfV8sB0BUuZzGRYFh2/qbpDlmBNzsaBg8hX1Wr5R+TfTFNPkgDxQLQBnhC
UofKlR2E7DUAbFbeaUN1A6GHXY744PjRvsPv/PW9elcP97tFk50pdODSxuGAfoCCPAKwal6b0zAP
z/BThCX5uKUtzmOKMjFn1QKCMzKxPYGTf2zlU2jRcqSE9tWPtiVNekqxs7deTMyk4pO6kObET9DY
1niXHx69uIRXgEm8qqr7iIor1lNfu96xZgnqkvCcK1vKYaEzLbGpClgmvykDMgsMCgCni8r6Nzrd
z5HUsM+ZA5PP1v/xCyTaRpe/9zc2f1JFuH5kDJpeohuq2Uh+EACKHFXSqGQQlUFW1XqHamc+n6jE
QI79qiHI/9Pj/KzomjVUK1x8eOEP38GZ3wV5LXCzd8d46HX0O8pDJL+URT0HpmdMkmGLSXjyqSjX
otZy2xluj9zvJaCena+QMOoe4+dV2kGPejCjawBE+3+yW2wwcD5cppO7xIF8gTVVBD9ItO6uthBQ
q9ix9w5dSZFWHziQJ5vZpTcy6XLZPqNmNeEmT7BJrHBgJqi7Bm2Y3hUqTj1lyI0WRR+njw4Prps+
iWtDUfeu9ewgnB5GXe3l27c73oDm4jciWaIexUHJ2wSZEL/kn2O6ANBDTw9oEXz9XPevKVT55pNr
7tgsNvg02JVeXVUytQnt8XLiP/qpp5fhVR9G+L/J883zj0wzWFpIQ0S0CYwxYPAK7y4+tvzuY1o4
RXHsOKp8SYyokvFpeh8kmGImTP/Q2CqP8R578ovL+oJpTw4J9PQoAVQToPUuIOa5t+VCPpxLkdvl
dRe1fyYvqF23Y/sxRUMlGw37w2139wOQtn02j9k1AAtTcsejFhe7MFyYtKEUoEIhWC/DpU7LC5sb
tudP1cf6+uyGbZSSE/Q26k//bmCWcj7jUthJd4pWqSLXcpQ0okZjBcvjkUDHMVuYApM+VJL4slMs
iLDYK5FFg5wgZw2juhaanJ1G/2tGf/9mtVuSuXA6EdwB3M//J1RBRM3878ztOKEix2+614UU5x3b
xiD7ijDdqX9gJ/r82S+BynXtU2bxvYWzMMguGThc0THUbaKhvnTtF3vGILYRd1eFXkPFvKVyI+bm
UvbBjHWL9jQBD/FoJaW2eOQGzXMTAr3YoMLTpxngVLWiiHvbqEDfg+Jk2BUz9igK2FDJFRzMs8cU
DyhaksHuGN6YyH7dZv9pWDasZNR+RN5CvM1EKf4aNDsJ6DxxLiU7RLJA8ybDR1gaeeHZzVhvNXOJ
59CTrZ9HLJtsN0kQb5HwgRTNef09gvQLF9V3s9yhEOLydJFNgLmRd1mKoHFaeGbW7HlklDhdd/e6
hokKuPnX6NzZhnIVookZ687CQw3pMQJg3JzBMGeYA4k5W1lPOgVLf53DxvYgk4vEoCQkQZiKHA3m
4/og/fHckadfpxuvzzz0CSTcnfXCONxiLY4NFrW29uDNLI0ep8EG2PRbHqg2Lan4HGetExrDaqnK
qT+wKkMRHet8kwLINm3yLweugO0Xz2BQBctC0T40HP3vkkw6Yi5UTG3rJX21hPzVZXuzfBPL3G3G
Ojhs/3rhkf+uKZxZW5nGU7qYQIfi78LtgTc1KmMn67fkhuLIYFSUm2ZslVX7Gown2Ob0vunGskOu
pJUMKXWjpU7mYdgWFPqT9W79Sti6U/K0moCRcz38Maab+8A9vU/wI6tRDSKt5/m2cavQInn2lKyi
hLTzAwc+lnQZBstRMI6x23U3j/ZtrHGtk0YgNCe0/H03Xo90GqRdfcgySwdFnjxnyD0eZdNq4JhB
xKofANsDMODjcQ1rB40dK3RWl0FV+Ie946YU6iaclFzq+QeN3kUZRRQBgmx2SoFMryEktJufKr98
3k4fcgUFWlMkipYSFz2tZAKOmUhQP/1m0TyU6bz4epPWCagECubXGMOGSL0JgJvP7VxypKzTNxL6
q9V9DN35XckFlrjXKT8OmbaKwg9XPvZkxFMQQ4foVt4nVjjPqXRxI6fo576cQ4eWC7WKlqjyEdfl
V/FXpBNljVqympSPqst2VnGvrP7ligkpXtxThojvOOMqN8ijvWMoQDsKRbygs/6Nx+Xv2UFvHwwT
pEVfScPgxrfGsgSMLhukW+ERJV/XOZUc9W7VlJSynp9CfA+3hIwWQgV0+4nIAsOoUzsZUIO57Rzv
vZzH3A6vcODChesP5n1heaDbXXCazY2bpHjYg2/S7Ac6ceveg5sSfTLl94cIpG0F8bcWcQiq6lvs
1u6jKJVsIR8azoS3iYPVdJjmyUadIjILIDkWOhqi0BGJxA/jxpKdqZfoR3gcIMu7tMdBygikL6+6
m8Nn9N/NBw7vCcGfF2+oS/W+ZreLcHuq2a+Wyh2/BJlO0VLThvrjqHx/k877kdX0uHczfcmzwVbb
5sxl3ua3PwWZikXGkJGkIDwnwgKnscxtSWnWS00jxvqJOqHaTfBhFhxXJJqLjiqX/CiPy3hqWA/d
Zg6trU/SRL/O6JqjqbCQclCMyxyxpdz9TsOISsoCZFuOftm6pR8snh9uXXXXTl/VrXMBUm0VisTp
vcYYOLadDPkQtyYqpprXSb5nJ2E+KHUquhsTWDm9IGPSUJa3gs6Nm6TKeG/vl2TeWUigyUZ9iTGs
luO9vTN0WyBBupDW5tL24J0ceeb9S8imiEWRgQ3FNdZ9quGE1uSKyYhsexRuP+PS7j/qK44Q+vKy
rfyWGsWFqPtCdEkOCL9cENjeEFNKMEkvklDw94pTyT2wEcS68juPo4aD/eRAQw5kv4x9/jY6DNLD
n1G24Tw3IP5RnltiqkKnhUm0Mu5IMICpXZYqNR9ZnwbS+neYOOS0dyNFWvZh5LAJ0kmJFzTwJFBw
Wm9eKg5zLu90C6J2d7GcxZcTx2XZ1Piu4RLYZzDlMXnrr0ttrbg7t4T1+Q6cd3OQioq8wW65eGbO
zgUHI8RAMw1ZIiCX/gAhP12RDK56UAqQO9FOjVm5W4/4jLTuAMv7XCx0WKejfAst/CKqz1aTgqBT
ngHJ7QyRDky8Y89MPRlyYsb/4PbL/Nv21DQ1/PLUIbjukRDDSWA1zgwuU2lnB63RQyNq1+gYq2/w
0cj9vDntJtH9ax0azpCiV5ZNW0k9RATgL2KA5ozb8vHh1Cloa+DZIsBPmCzOJG2pc3Rhpxy9Ukw+
RKFwnyPAXjvqN84rqlaqBKMFPHZWhUjPRbspsuC5F+7MNk0kIQiDMX6FoawigAI1Y0tBIh3A4lOe
8R07JM8WLPAOG8MYEyH04haNKFiN4r9RuUmbqD7gZR1FJM3WU7/bEl4JLSGfpJ6sH3zDzZEslH4F
UnYXCksJSl9vbkd5VpoACS8DMUzmzpbLdPgXPW3C3N8Q7jMtuTlAhpp5dN0zZKeJ/VElrInZCNqG
JZCFq0wx0rIQ2eZxyZYnSAQL5+rClbATvS9dDtJf5S9Y2eSex1N3upe8/vw/nTm3YekxPE4K0shg
vLIUNSkYFklYC/CDkJQ7QO5VZV2Bpo3UYiN04tnQuVhr9u96CTwtLztl1OO+6dfmSvLoqoLujHm9
9eOcuQyTIljob3LGynN5G6wNKk/luiPFb236I7v6Tzke3SscMMidunYgfF0YospRg0Zi6CjEsyx/
mk439qwp8/L3+nKkpzeZ6cUfUapP8v/W0brG/L7uoLdPHKpsB621vsYiDR1uYebmrTYyPBzBkuDb
rJX69ioKWMroq3bJt5Gprrp/qIPt7Hygag4wuAVdWGU9YOFrupe4e2uG+XH+wmkyYzuf4v1cpzsE
r9FDj8RVJNegeJn0VqVAMFx0SizDnn/MLOq08irI4ri6CUQYtLGk0qp2iaJ94AKx3BD8Mz13z0Xx
Wj/QHaXU7sQweaOlsoVLtnkvjjZdz8FsJvnsta05iJdL0dHbnkYXOPUCbkdYdQD6Hu45jzP0pncR
KDVBBsi6n1FVd6opKCVkJ11Ovf3MXyAZxfbUTO9j8R8bIin15MCLrzbSKNLe0xuOvXwuIyddNTdY
UscaTBTpARD9A2PaPk+Yb4UXn8Ii26XXUPaXaJ8ASTc4Xfw9/E6ElpNMcBsNo7HN8WUOkRZpwscO
jpwF44ZnwYSpdRtTYwaSnV6XYCkAf2gaWhij13LmpAr1EF7u9s5mL91rfxd+KYW0CLJr4Wh3g7om
vbdK4l9oHJ4KbDhgsMVJ6P/DpVneLadUDp4+P0aMtsi/k52hmHWLcIDDmAa735vLZ0Bphc8CEv1K
Wbec3PuXXLR73/ohsJN3Y76CtHevOtylXXlBD74+7B4jK4/Cos73YV1MpVp+FWDVyajd4gkLSBgG
3Dm2CuPpNcu13nH8KFPshkUyuP+oIoYEjJXCrX7r3DgBw13OSIUzoA+7d/sVzmAhaGK9h94HHStU
b+O1N0MepydT0HtzjclH+mSDcujrNPu7ABlzQT44F9xu9rahqiCHVFTwc0jBay3WwvpNpYKrnMHn
M2nligNuZ+qE3zdsWP++wqX4/pcpdXkS/O6fZ56UP6jQfo9zxqxv55UTRcsyUuHWQADkUWg/Ag4y
wJIsdKE61p464B4ccZ82k2t63ABWw9IjRM2xlXlb/alzmBerio0c42SPjCr0Qr2ePdHCreGmn5oh
KoD8BbMPma05XEKrWpT1icMPn0gAOorFWoon03hz0HgPxFSpG0ujKvbabhupid2JNNMT/M1pGFXN
H0ekh/EWpKSMUM1s+L0kA13QqklAyzzhEN2nhjeLSI39DfxITXq38UPOzV/Wo21D7QQ9tDgPwa0n
MGdoEY5riPLGgA1b9U2Wb6I1D7MGGONZ6po8ojDkS0KVmxgzUL33lXN8j1ITDFCq3yVuzFrsoLZE
PrUmI2YiHrfvsVvvJ0dGBOjj8q5ZBinxd3fng9uj2rPKmAVeHh9VfDIapqPhuUONf1vfspVtByYi
i9yZXtX8HfZdDu8z0SrSsFs0NDxbzKqBN06NDbtrdzmwfD5p8XcrIATTz8Z55OS4EdIzRLIyKTqq
0R0Pfz1vKHKdJD/718dfRlp+jUjNPHpOAJKrsyYUc6f7YPwEVPSmzRttOJwWEW0/KqP0S65GKG/S
+pmppcMzbbCSGGfWz+RKkSoKU51mM3qODjzIAW5C8W/1dvim/2Vk2+hqC7GbYm9OrQZIxBsiqb9Y
qCGwyIyHphXwx/BOtWLAvuI0n+iRxOYiTKrLsjFXkKQgYDQsL+lA32voD4gyrt45rRL0eo+qcRug
44/SOHrb+xeu1Vtba6atavk/DhuzY2vq8b7TCXvHLPZaTTF66PLDS+A0Csx5UqEmDkmWSZHRQqIa
uuttxZXkLAtEH+QvYCb3bX0LPIWK8xSe/P32SoOI+gVFTehM7+UHLB6Fv8pNUzn5Y21+RxwkOjPB
OHCFETSMfwq2AHZQk8EGzA8zh45TeS/HZ1lp7Nw0fhw0KaFGxvSLAVpI3uRdVBpEdMMSdH66z5PS
vQQJgEcTpxls4dem7FwUkcCH9md46MH1LXv+X/0LJ9PyjGQtYTHhaNE5dfFL1HE+aQbSr9rXGRMw
udnOMwhInawjwBXuc6UknSqxTV152RkqDRdO1BDMc4kvksD1UMj8i/tp3bBA63zMCltIbLf2CtET
3lhJtVW3Xd3aHvMIBw+Q9QAFWFk9oNkLPuqC/Lv4/+gN7yVxCTcj29ITgFBsq7WuOKACQaJy6K7h
m4zWZkfcDKpp17qolyPRsHOzqVAllnAYuRaZwr34nvwB1E3h6lv2cCCi9bPLFVuu871BbsZ1qiiq
1JwCPujjNugoCo36m8yi88TdsnOanCZGApaZgx6MvIxr6ot4+2YdRAOnFKtCk/x2TLKgIcQiGiq5
whizcIr8KKsUiNLshyqjxfctl4uSPAZeCvNR0md2bujAjlYpKUZrAbTcQquoOrIEzMKVHU+4Ojk0
FsfRbXYIl+1JN0lqbpMXOUPUZnKGdcYoncEvbIWpFuRA7xwAU391ModHpBRS469E+z2oJH22o1j/
ReqYrzc5NX/VE2Hxruf4NlPJXQPHTwZnwD+eE9/z2ypjiQh71GsygN6bq/Wx2ocXv/wAUafqeqPY
WXb7ICGZOJCMCTOGW/MviootR3sjyJnw5FWikmEm7U/KfuACYCJK9HKF42J2JHI8AGK7KQIs4ui4
kHHKfwSP3f/EJnkVyWmdWEjn3CP8w3qUe2TcGedAgwBRQPWuwtBg0KLi7JiqNf2sJv1NVu1qsgOZ
SUliXDfQV0v10poVPf8uV+IIs1pymFLa0yedB90pIHi9xUUQN2ISxomH/Q1kpCT+oOYyAYsRy3FX
HZMtVOVvmKKDVy2fgFujDPDvlXplyNeM1Q9qisq2dYxIhEL9PQbJq5+BtSsYnq6B6dhvVCtgn4yj
jBxN+l/PdfZzLEGvpTYFCzaya91r/dIX8Pj/DTLuGM2oZPoPivU1yyrF2Ab0L4FUad1is3sasRRi
Iq9OEJGfeRZqC7HHpe2b8HAXQtDDDGQiF76F+FYDUqa8t3R6cKI6Ruu9R44Zzd7klH03fcKr8VLk
IUKxFor0HDchwuSQl7v6sPo5+UruAID7u3PZ4Pl7THH9Xr/qH9IZ9SttMNVx5HuccEc8iE2hZ1Ei
SbLkP14Fku51lwCwJ4G23PXdhD9jxIAgkR+XdCQaSVUrArqenc89SBUxwfUiE7I2dvLSPZ5xPfsA
oRcZbIPJ+2Zw+GTl0dWZpLq+SeBimc5srnkjEa23mI4GBPGXf0dAPivKprFsbDzwSc452HmN29/G
R3a86n8evKRvK/kH8AjrobFKbCm4LuJzHIkgo/IMTmcUIwhY0KI/q7RKN/SgwoBKnQ/zOLmr/Kg1
v2rEhdUNPFDn0IfUZbytL4vnaCc5WpEQXriO1Nf7kRDJKAgqBu9QVrd4Yi1jwDmULhn/ecXDXlWZ
wCXVOL90Ff+kgg8uEEV9MvRd/amLOYtBvI0EyW/zY9Ujt3FS8Q1o4KJZWrhKFwRyG62s5JRASZd2
1z9O6HX29zHJnoOD0qr13PcIyXU6f7zacjFVur1eUchxAct2AZz4Q52qjwnzepExG4u/Srqi15PD
1Usw06ZymINQmgFsUXwPUhBpQgcPyepwu3sp//Rx1zGRyI6ke2FGuiirK0gkLDGPEazvkwDCI30P
BSE50d6vNl0ItjcG2mMZYScNBAod80VA9Rr0V6r4sGNWOMOf3f74Sk3ufdQvwpDyODS4/woFJABl
/DbSviw4CluQghR8G/yNv3nMo/QM1p4qAuG+XI4MGpLa09jX5gnMaspCEF7V3iTwCSzoZDnejP7j
T3lJQEsGswOQM9m+Vydq7hvTRUVQVmPu+doKZG+hFrIkRo/mvlpvWcrRHlgaN3Jr6DIJxEUwsLdM
G6nospGCSbfBCMwSkDnES7dtd5m3JZL40wK7IBgycGSo7LmlBXNTZDhb7LV8AvzWT460ujsnjRMN
2u733nghAuQ9n9pYRQsyvh5/jmXYQvbhjJZO9wXvzCpHjOuUIQ34d4hE7udMLwGxxobhtWEzjZel
0kDTnT6rrD8ARmxU5Yw4J6FJwB2twhXb+WnfREJhqeHl4j7ZlyC8aA9XPA6vdY6t6vIjnDDJcO0k
G1uBL312aa2ksVmxk1I4KkfLK/I8HV7FTbpFXRLBHRK7GUpbCyQa5Gfg0cbbEDFNHu9IkNV06a63
epgnVrGGMQ+784MwjkJmSXdeA6FBUOHx9hMCiEATxym90rLYACKDdhnDgbFFpAhhxeR+JK3Drpds
6xfXi/huPd6QQZ4ymmESLDaOT5sG3xdlOEM4AhQ3T3ajb+TbAK8BxERmC6lzPqkv9qQWgBdifwKe
k9OkagZF+ovYnpiNYzexow9OdppYa8twg+qNABx337bLL94U3tDytnpeZ/brUqPmaenLoztaUl7A
0ZhVynHgmzqOxOnGjKU8qUJR1YQHQXTvzRdNB6m6urI+S7Qw3F7E9/gdVrNaiW38e86YUwJOVJ2i
DOLfbmb8LNnsJjkwhjOnhym9i1kX0ES84m2/QadFqGF0sDo7p4ZAd0PF4VeTI4U2vLuJo7N/trAN
Y0YcnvSI+x4bVFx7+YpFj3fJEDcWLJkaXW27hghOK4Co0HDrO3fyuD+Lg1Vppr5I/hBNralWcoIj
fxXw16jXSBlFA3s1GjZ19HNW2ihxIvKr9D6RvMUryg1j3PHktuPfkt5aQaaAziAGXUd6ekS7s4y3
iTdmGtFLWrTFLN4HIAgSa3xvfM5uqMUFED/YHIABqZGPVjO/rOHFAPmfSP5JqTrsNobHcKxqUe6O
1lU167/gaTcg5tdTKEGsLNNj2oiE4mlXLF8KlnbGaFPhuLefsKdrtBxjC2tW5bRZY0rtrBhXxb3A
2+ZcE39P+JAQDbPqM1P4Sr8wCJ2rH9HwPs3VkO8D/VyjFBoPZ+7yBJSzWuEeA4zNP3rDYTmUnhcp
uyVoXamNBkeDS/6JulHR/z++KhsiBmqbwKgCaVQrtPrLJtSmZxf+HgPzZ+YmHsJr9TRJ/WpSQUR0
og6w4UXO9I8YLuaCkc108MyQCTGP8LyY2XSvJsJ0AnbZ1iiE3n/471d7gaCPXos668cVblEg9XhV
CW1OJ1R1OSccYbYaYvEmnAsC+a+oA3pknyGjzamv8jSuO1GmF8gZZCIzxf/1eLhDH9QugrfTwpTI
kbbppbhEPySLzbvR5mfxVyjE9vxxUnmxbjpMcMyU8aJGBtzknx1EZTTq1HtD68c320s3QYVPCFjy
rVNt+fa3A1c8iRRaQv70/xqe+mL6x0VJh62ehjJg5Lc4pg9qm1FdMrRVyzP1v0cQumW8Di0gzsG8
HG75iI8Hjcs+j4Ilj31apsbPSrarIXAuFiGsUB+JqdYYrn+TsO2hclSxqR0qwD99iLo1IaMqEAM5
DHO1Bbj+HMM+OiF+Ip5bSDL4fHuAUx8KhPTMyD67fQ8aCMV/IyPwmwCpI9xNfn/ingyfJ+qsp0og
drX4u9u0elokUFe4MPIdxUwSnK0vHSCm3nRi6n3CDFlHwfm705Utcq0XhUc4UfNEAm89rWA/Bw0J
TGT6bPCQsjCGm5KCi5JppopcuYHDTNuqbehn9s4ub4OVfjUXl/BizYAr/RPpim4+MJHMDO92brLL
hGCu1oQ1YCRC7p/W1DHyTT7TzD+JFy59Kl3Dv+uvcC2GRzy0nwsglUIEjaMa5Za3d6xR1imsuXaE
TxDxUhhuqEitySDk0tRKNfKhlVj4xV9Oa3phP1OTPrly4mZp06/oPFd1X6TUwUCop6feMQlSRiTg
YJ3OBH/hJVhAegnk8qAauYpmfcxa+QwH0d3a+95MhSVfEuF5gEACm30Z2f+S4aU9N8fgT0BplCg8
GL8y6b/8oXobwePjhQWtch/7fk/QapWbhfS+DHvmvk0fGQkazyN63DBKMjITKfJndV56xLo/q4o9
Nug29tmLyKaidKmFD9sZa7nBb1kdJL9JY26p6TPNmw/KnzWzoqI1SlgxajTqwzlTHsE2bC5MnTfo
wS7ZRmMwAZQ607hj4Auf3kqeQsOgO2C4IyidzJitV2kokOCly2UMwM0U9ZA03HMJC7FHfvjZv0XV
l0caXjXpfqK0bGJRZnFvs4bujyH57iYgNDR5y67ImG0ZGvFpMx7JYiX30Jpm9bu3Mq02ihq+D6rH
SgGz7JkkxVRIpnKHzHxyFxq+UeYk3FcDysLMshVOpNxDWDE5Wf6l9n3yvijhqfLc5yqOuzoD+dZ8
dVbW9SnKlEvMAFZfjyx70tNd7mNIgqCvVR/57FWoGTfTDadzfGjZolNLoeU4euFwS31Ud8IpiyKi
IZOzQb5uj0SR6CGYWYTTp0rUExffjfxhBnQOUw3vHsNmFiehrifvXd1/QyX8HEcgzmBqvX7KIJ8X
eHOfwJL2IF5u1yO+A/iZpgc+IYg7GFION2VVmdmRmNYUMIlFTt+ok/w+BIMnQVGPqUdNJNiSjmmE
dtnUw0fqepCDyWUAdvOowSWA69m+J4rI1NKNlVV5PNpFxoCf+DtvhRu3A0d4S5Hts0Qsto9iTJkX
iSXsvxlbQeRB2hwbSemzj2htJ2D3i4Igl+eXcG1YAesnlcoHnPm+GUkZU4EwjVUmnvHMKdxrHNqq
+znt6egTLD0x//7JIbYaLOiynOCTwIMEN9gZ7Rdoem/C1pD3XKvU+j8r5MVnLcmkVbvzpSL12wgE
v3C6FCbN/y8vxos5+D8J3lluWJHaCcOI6iVaWNMWGuxsTA/HvEfQ3EwwK/DcyhuDsIglG654tNKI
lYqREC2rnlcs7Vfpe/mP007gqcvtdwZjaKGL9GAYPHCBixulEzI8CxiNg5XqvGkE64fx+w7QF3+k
Uf7H+/bTj7MullLfcrUHnw2detsFBM8C27U4K/+I4JVPfHGsb7anQNDDzECnj9tslRqjUJTReyLc
s+rxE0naMWWh9uWUewLxRj06YGejprQRYCcNBDOhPr2Av04Q3jfOIR00SwDI8Em1OWuRDoTupHhI
FhRC4LI5UGfhnotkMoIEkQv9RvQy+tofMMJsE3A6C6nB3UVPH8q9dg5HzwalbWcDO1H48jPyP4Fn
zZgw5CZDTngdpDc8IYLCVxaF1T/eBhmxlUflrZZKJs7f+KAPQJbLCMTFaI/+G+aUGnjW85Y4fpTO
tMMDcURBxz02H3P6fnP9prnbK6W4SUTEZv47sHthSdLw7ZIydwaOASXJipg5GmnqIk8zu4jJ/SCm
jy3+sAQjxKUM1hRFUPfcev2J/9NoEMIzU2bX7HBPLg7hFEQRVdxDMLihHCm7vBnemfCA9EOjrpZy
KThLGkudrAGCm6bxlsipnXMMB4XvXOpfEH7RY5mp7yU7yfU5GQKFo4D9eatzPMUtr/5sQJlwPDzd
lteQUmbheDkCHg/lBHOdhoOIU88miks3QBlPeGV900bYY0avdIvyeLyl3tBtngcNCjMgSakhWmlc
z/smIj6ipPKOPAPlaE9CtVjZEkrLvvs6s1Sat1GjeuX7nNiO0HdLqiOheZNlCLSJdsBmb0oG/baa
RgUBE2IAcs7U/J13ens3BrPIlUAh2hu0epn1mnQys1yVcY82qqP0PwFreW6C6ynmd8BR2uMA3jpV
O5yFAx/tOk+13PMUWmJdW3E362JLUqiDm2J7SBcG+1aBUguGNdA1jeynQ7W7NRRf7I3GpR56zB4O
9Sk8bHDltLXyAJCi9r1LHXFBBWcRhoITTNUqCyg5oetpQdrfczhIGFMUk5bfFfA1lpEgEJ2x2XG4
e4ZZ/7vapHMhuq2UTHjJ+Q6KUxvqBvnx7GI5+OkGlInRNjyLbB4wP72tuwZVGRxh/nnlqHJligdA
W/V9QWDVxJDiapbPP/EIjDP+gmFu9HkK0lGjecmVF8RY3Ln0kZuGc48BHOI9A87FTJiCFMkr7kxJ
46gOT8jmYSIF6mnwiVYyYjXg/TE8z38XEO9+THLQivq1PwlgeZIiMDK7PBpKgCBQwq2NUD/QhVAb
DqJcfL/5wfqRjztQQregVqCXUD37BZ3Uz6vIdqKHt/d6wi7FZbDB5wV/msoKeQ1bzLLNKIujnht4
ZDZy462OmLd3Tg/BvMvcxL36FgnX4fwv15DpWrVfKg8ADbOc95hKHDp1VABb0bZqJphtNnwvGGX+
IjTPx8aKAM6I+YQFqYjRzzPcy/F/9TDKAmAY4JHtBBkjBolUKVDBzDErlhgrePK+4KXdF4d/Y7vZ
dmQQBkoPIIRcNpnHLTlSMABpHJSPNKXGyUevkbI/1N5kHS/+ngLD5bsSVyvz1Xf+MK7HGPkWzqUU
T80ZAIIzEH44wsOxNBkoefNKsLNp2QgiZZO2pdc/raYcN0oIeocvH5ID2cJFTPorkk7OePRXwzyx
TxaqCH4+ZC1SYcBnCFd3dh/gJZRU+AWY6eHyD4FwLnaJrgLaHBxArrYICmEmMRLKF1NJm2an7QpK
oK3VYgOIVEkL6XIl5CfsuhfwOngJkd6F7JOH81mfcDhtkdayNlh2YBuE3e00DhyazWwT8iWoVI8t
XnMxgO0/othZAkPSzhdnPAw4Qgf2862garHSyUKmDcAdegRWRRq6RME9E5tPsWdbnSwQrmXVAktJ
cYIiTlhcH2xuxirs2kHTTxZ0lvV4eexUnx+22GoeZzaTljs1dcSPwWZMrNLL9ZJ/J7BGrU0W8qP+
T5s31hjWi9OfXKzxieCab0jmzsApp1a9Nv6yF032X44jErEHjO7iIwH0ipnBAiqfctJxwaViYXB2
JNNwv5fwCxXi+lIPo/yNJ0b1KNMkNUo2Fc9z5sNm1Z/1o405D3lmuBKdPpn5W+ae/1s8VccMJSBG
gibzHyUrDBzycbJneR0uTZLNjn1XlFKSVH/e/jGG7+uOW/fjchntQemYrrhulNqmJ1TzVdqAVCc2
V5wZoBeybONofYz2PKL7Fq2plVVGN8eJH8rEsaaqZAFqSW8lCjJH96KTKRlI5W66JtIUR7wv1JWb
72SKX/GZm5O22S81zS5I1UaLJeIlv8TtWAxlpvIe8yZEG9t6mzaOXzQTgxI7TJUrGJlse/K3RsGq
+ieBoV7a+JZNotEcU7rtr3haYASjEUm8pB0N6DleWc2pp4kWxoykgTuSqgEACLcz304I3GcIg15s
bTdWDuZ4tPMZQs3hGuEmUHvyk4uhAiV2XAluXinsJxDTg/vH3UIECoOInVBBStx4G/yYwjMQEB4a
NaQIFaQ2HUip6SxjR35D2AWQTxWRfdjMlm31q0uPnxa0kq4+pFPBZsd3CIswfu7XS36LXnxnvf7q
VLxluuf8MC1WnMV+UZv7j97j+V8zR4xbQcv/274cyY8BYz9ICZFH6313rHSEaPEcXlUq1WNYZlfz
j9x7O2kxJ2aI3lhiQDTvlL1XJrnHGW4LdXiUSHhx1fthD7utobn8+w7rO9xgiGGoO1N0hhVekaU2
OyOcBnKmqHgBAQwjd2+9pOvy6yVH1Op0JvmkGluvZrWWhJIzdVisJiFfZwN8hLwtldhF6HCzgnT9
usiN+pSqEQCSIoi0JfV2vN5s9JeiifSBG7PM5uyLMXSnwi024oxtKdwGml//mEoMCXKN9oVcpqTa
qKEbYpXKF9BxIN1ETdGB0IZDxbkzunVt0R8/joBQ3kvr6BmpfU1D2f48CVIIx0dpRKqFQu96SHPL
1uQInFwnmezb7h26+AIFYgNEldKI3rcSV0XL/zDykBkXN0rriFfvWtoCRcXeI2f+B6UiV6iLdcSs
oBU0KF2Ty2QVwElBwiPp6V2Y9dOd5M4Zc19wsXSDrMUIb2T4+rH/MEOxQc0GmzwRBw8YZElP7trp
rOmjP06O+T0YGiDldX1gfvk3CPfRQ60pOvD4fYpccEEvdpswTv+9jymdtN+dQXiUGKR7/Kzz6Rsn
e3nE83E8zJKJvZ8KXPPegQZidSVSW+2BxM+KAHweNuVLODtOMTKYB4Z9O0X1hFapE6tmNZ9lpsa8
RjRXv5f1hadAFcKXKD3yBcwUHyxb9A+kRK0zmLZk1S37tqoFc8hn6d6F1Ux86o1y3JHmqxhLCddj
6foafz44KL5Z+WPsGEinhuRNmGMsU6Bs5iYTTPYTFZ4Ei33DUcTCaa5/3JKOJgI8/GqOe/IoO15R
G2je1JboD0YT+0UhFA1egbrN9tVRf6CavP+UZ75adzjqqSqn62lZ4yjC5EYU+aINrmozJfo6kpdL
gYhqOQuBAzx/P2vVZpFzRoC0k7+/RRJBSwPV+55MwpAwJoToPI6Ph4E9pnyTGL47H1atHMiUoDHl
F121Usnm8BAc8uy1Azyd+obM+ORZpMSM+haTLFbqFvwhDNx0qqnqSdcijLYzVWBQ6dvGslAmSsFV
RUZKZGqP1fAsGBJxecuhbFD8MYWjDIW0yGREubz3aqLep/Oy6y7DNCMSf3o7WO0K/38aNkcIvtBV
oexwKhKxHMEStxQvcN6esI4JLdp1DGNA35IpaIa2DXL0z89NS2hS94NkqE/naHIEsuwOZAR57iJN
WNBKumzqWuvclS9Krk8XQjH8BbLDUTq760/sEEKMdfm28+V8HIC8EDxzNg3ZM6XEQpnGqapzE5JM
neks4O9bk9wQGvI9BrvdjfhLf5yxX4hTkhzRsoYf55uZkgTgmC6gRakt2wvLQUMMTqrgT+NuBy+S
hSb2cn9ky0uNmP+DtTKadGyCFW+zxmfVuBasKBMiz/zEa6rnRbD7aOfvVOEcgIgOCnndLBEB8dAM
6PAHUTBVMeWtea7KHT78QclOm9IA+FBLZAe5mObwXI13EhAjDfPMrG/5CJd/M3cUQm41adyl/2Nk
Akq3EetapYgSOtMtossKKDOiolljQYJoDj2v/DzhIv1HazV8kHPi30g0tT7vX6/FV3Sh4ZuZyTJI
79UBfOIijktjLqboDpccimPMAtRx4IabHmVKuoLzGyebV/CqUlujN9tvULSavtBex0jHiUQSJCYp
zFZ/4ETGCzPjjk58NPqBCY9996rLdgZUf6RgfKE3vRuseC03VDhwN9yz7JAN5iLp6ikgkrg2jlN2
23+uxzRiM2NDyDvKqpf+BZWog0uFz0Bp2u75jN/BmqOVkcr8f9YoiSbYUiF1mYweGZ9LqoEPun7Z
vO+gCq83sLOVR0K2XwWGYQt5hb3e2cvY9tNekLcNYCcN0PyAhXOBoB38M8rRRDb2SjENmphjMnCs
0046Ar3r35WXCXAtncvWecez4/lg6tog3MsA3+GOxV6aqzaaAzmjx0iX5egZdY7D+cojj05AdZ9D
DqYwD6q6v6TmkUMNGSBAtC9gQtppFsQl4QggMjl9pwopigFnHXnym1XsB3Fl4TQhVLylREsgaf2R
/zHGs8HDYI5k7GNdWLyrBQ6rPtTZF7YOQcHGCC6anwlehSoSyBij3g/i7QOVyTsgDU/X/39qXsa6
UqKGOgJmfBKVddVSF5QVw6ADCkbuymz06+h/r9INVmaNKD7iNUM9PEXV4SpgmbSAL1t+mxnKgyqu
ukKMz0NNYYz7rzawiXD5uHOL8E4GvR0BCYaf8K6FLGYD+brb1zZsLMfYkQPqoneM3nRuqQrCA1g8
Odh0b4/BbTg5j7t1tyZ0Fk579zD/N9qXz9qnXeZCuLtnxYdn+m0KR2aYYefSN7KhJkrMf5LO7XbK
8S0jFoFSqtiibSFelHzHwcFCGHoS2zOw0d434AYy7/Gxsi41RiYDCCTp6BzFf7mRZF+3lwwNxN3x
rjKyUVXkkiVdovWpAgCSuv2qbtWw2FjwneI8K/9xX9sQF5mB/xomWrIgh1VeKryFRA/80z8+Wpu8
n8ZuX9sk7Bb44QpKKBaEI4g7QJOc2vzCB38tCMd+iIUKbbnlr4Z5HonWcLD3W3x7tMPRG+Vpk45s
rJd+QiZXzOziuzixpiQNHwlADjphzjFlgK6cfBWTAcPDOBEHZwui7eq4C89asIStykiaVovIf8yJ
wOxVZtoOKkg36VLD07PuLjBCpUxAHsF17AEkTtOZUbKP7FLr/YN++8m5/8AtAWe7ixWUg1xwahGc
rVlKVTp51/0cjTDjrYpG/FBawLE2i3xnd0mX1WofnLybUpz0dPlWfbkdLgWyfneAtlht77LcHRXD
Uai2bwV6EY9Zt99+qdZ//iFeLZdsbQZ0SWw+xzE2+LOTj4EaOjSr9uFwO0kd9vG/Nu/wz86Sazl2
BpnXXbNH9wVdi0Pxth1Tj49ZOxEJoPzMEY0Z/pEuLYnIem81ZUYhT8YmkZr/2YmGDD49DEtPaMqu
qSaUstOH2L+ofMTWW46qZYOw9armR3BkMxEibBlwOuCDzrYQFITkLCA2FRplnaV705e+pc4dQNs1
GoC+98vr7sLYJpAjYF5TVu+TkyntbbKlO0LY8eM+Sj7yd+7vS62TDALVzeJfbMryZzvgY2fIMZpl
H20JkNxo2obwvpmDqV56Z0yCUUD60Y9MN+BB20QvZFp6ymvvKrbxTf6852m0+FE8VCDaefZCjNtb
xdf+Oy4Z7P1juYFTGz3GCPrKug8B2uoUsYhuewpDptY3dF4A+5U9PWvpgKhRX2vHnyWbMBI8fHVG
6cD1aDs3+jBX8TIMjozy11ffnE5u4QBToxJDn1hrjCN3nYtHYvD/+cKmudktwU7RMZGZH0Uoswnk
54rhTnRq5tN1Siu2O5/oth2LZXD3kFhuKZp6cd3422YeamhY8dyeMNEtuID/eYjVZ7SsLnLrvoM+
tofGzZEiUtiSlBON+RdBHcU74ZoK/U9xg+/FeZBxdhYHewQZL2stPdH4gVi2OkHWRxcKoyqjafgW
qz6vwdOiDLJX+rnO1ClrVYbGio0PnlYkilmsqXTeaK52iJGf3T7+noC/dxf4qAOrwFVVWoBWjBOO
SV3hSwTLdG5ntikSvQB2wRnTJGAVPDkzlOtgGZvt+0UboyyB8TQzHAdYSlr2FnHw6LPYk6rAlBGZ
WUaQdT3EQ/osFb7ySxRUCiu2ZwMGNbNepec2OILnnbKOaHUHBhaLCGMpZ97lyJD9+VTRI7sfOlJS
ASfY5QlUtAzJjREADtKr4c1CE7IFLZWmN9huQcEv5Kd2FggolsDvFNKl0/XXKsl2m1V4uMmboJhF
n2ncntoSYCua06MHZsJMYD7uLFUQRfrzW4Db5+F+CFNgCtiO1CTzbdljR+eulxicuIgoBNilerkR
CtIqUpbg9jzMRSKK4TjhwqpwVQVxdMI19VnXr/y/o41uqGiVqc1W31SMJsBVLBp0RdpIzpO9Bz/Q
Kok3gT7NT8RkxAqD7/JA7f7AZCe3sbCi2Rp1BesrqHPt/lYWbK2h9Z46Ku6IRHMh/odeL09m9A+0
NnejWTcDgai2BUvAtIhVLHGFnEOxUL/sMIh7UlEECkkc3mhBnzi6YSriDw2OkjJC/zh7wc+4IRA1
1nqswOBX/ty9kMzNHYbBBUjnqzGt4UIIYJkzK/4UIfZqIqAJqjwq0gkb6U/kxHM9rUr9bcxNT0ox
7pNF5X6dIVA5qD4LeeMcrPTA/knx7a6I+a1vM3zLovOio4YVtiAA2yFSrGJ3mNJdPlPQ3kprnCcp
Mpb/JHZ3VPvWSJL+GMEiBbmHj3mGp5N5auP2bL+q2Kng3nbu7bsaX73ywr/NfVIbfiLR1Y1Mzb6x
G/7KWBsT4GsrDN9QXzin6qNUaWD7OOx7LcC0fnr0LpuvxkObAMO3ADHnFrycCqnesSy5uL2yqAGu
lZod/bW6NcrLJ3vBdgqkuNfHVdX5umUhFdbcrM/wCGcKjuIqqy9jwk0uZaLWhdwrcRvsgNgkJ0sN
oGWaw7aGvmUSqA3g90Gu3uJMBOGgFvkJSMXvPoZVzDssNErs/wt2cMIfTdwitHzNSF71YmuqHjje
7/lUn2hpz/dOR1RJwsdORBmgo1d8vVrXqzIyZ6+p9NMlHqwSPaJ0Tt711bujZQnuX7QFvc/Sk+LB
I4P4MJdhiUoOU1Be3VdNHnpA7RnsMMv4j49BQOw/M1mBr2whfcN+WeikleDACBkwUtpAh8lZT6C9
3Qz5FWOL580X2Nyh6koQvqipRJu07yqMoxtC3sBz9udxecZBN4CKpo1xg8Qu+4EuDS6rMnCWntyM
Eq+2bsnve03qD238ru4/h8YBWxu/kwXlFfDQHNiS5x6FD5H2FWlfXw73Zakh816/dakF6sTtV/4p
lQZ1iQj7vKJNHY/+7gMBVturjW4QCZCJqv/KTTFursvXVx1GsfKuYcXV3zdbdyapYHvGFxjKjJeP
X+90LkbMWpdMSB7nSypjNxiFwWVtYSgCbMlUKcxBL9xe8qTI7il9IjAYfSqStPCRF8V6ZAw1IAoY
7bvQzLhV1nefDZXmrbtKjbBUuC1+2fMbM59Zv/p+vl/oa1M8fm0I27p5QWkoAi8CwSBwQjBgKUPp
vVZNVXx0SpSDGAVrMlDRrZhuIJSuOLWQJo+JUgTLWgErH7FB3xpIWtv7IciD06ZBGs/J+re24mxB
A95KNz0j96SZPNPQ1nkLWSqnAOUQIszUkvvAs4ZJhh2mmpgUodBkZPsjnH2JD/ITqXljPf/YlSeQ
Oa07rQRNQ1DRFDfrCLVlF2uNTpjX46fOQCdhJ4pqpbp/3cggYlrJJgUXmI73NxG4ZR46vQQOvos9
1Om7m7/VesPQl1XcSIxWJZtp8F/gYEGYvJ3z3d7pmMKct+QOwjbXy5N3CVP/+L1XIV+uVr8H4P9R
5xw4zyET7cbnv23QsgDdQ4bY6bsKtN2iV9qTzkAnJdVHe5Q6Irfs1+VxrJBY7L8NYwsMCwoilw+M
4S5KxLNU9Tb4nerAHlKxFvz2+bKfKQOQZpE21PxjIGJ/7/AJVRyYE27W8bdyLzLgQW8dDsERzjye
NeqDKraYGOy2uWBQdSHytcNUnPSmOQgzvMKOYcvwwqXPwnodSDkPTn9g/8bkbGSz+hGT/l+rzUYg
2kYWgwJ0wno9+Zb87Vkhjdn585Y1qBxlAZsfx9rD8lt5Zw34w+3d9/7r+1lWIxH4S4Loloj7tsNy
sPzbDGTx1wlzxatg4SUCIALFj1/x0zYAYTvTeyddxw5lsfgtlNDlhS2gCx4sOg3KIMrFPxctRCtk
AVWXiqSpJ23+TzZMGnXHVrJZHIkSM7v2SUr4X+AHwxMAY4rEusT3K8T0X5gcUeLX9bDdsKOUeLcH
yb7z+upH6N/dOi2Zn6epZBHGQ2vTdmVWcXUGkpCJTCFlHgCuv2gEzIsJOiIXHQeIgnggNqvu15JE
vMnxzYRWuwz/oR+pqWcZaRvf/aIdk0K9n/asYJtaDqXzw1zwYiDqhaP2dt/L/dhdF3m/PNpEajkz
b5MsymIjdQkX6ARMuQHu28VAQ9owffAwO/aelH0v3vY+7MPpp6Sr1x/es3XaqUnhbU/Y8Cc5G+yX
Oo68FVt8fkZgUQFI8MOXQpIcmUkxVigpUm7DyQbkxuPnsKOiaJXaFImCFwyCQbWH9EdyMWaMqbkE
f2gjMkLgWAymW4VrKX1JpKa6IngjCk9y7I64UG18IDj9yy2vsCailLq+bwo2YcC3CGc1Xs4mTBSu
PKKUpJLfYYumv0LKanIHltFwDQIOwf51RxB/8mkre0TQgRU8eAdwnlRlo9W7xEx6Xt4UUUU3V83z
aZsT33x+eXZs7f7w+zJ1Zq14Fa0kUUha9gbf04Mmd0J3GlHzzZxfFNLa1yuRhYxTHL2B3SPVzMGO
NQgYdh7rCfMPASFL/Xp/h2bjhsMfUU3vRdRX1FPba7WGT3kKKQxFjiyr9HBOo9WT8fDdWOTA9tEt
Q0rsj14pGqlsVhNwTbsSXeoO/VpiRRpbrRDfWvOMe5VpQFytG2H7icG1m/eE9MSR8LWs6M05+MaX
RCGfAvXycr5EfuwHXW5h9fQLj7f3dlIhuF6xNgqOX9pvpTpXRoVxYv5u8zJY8mySdSzAz24U06eF
3F3wM/K16aee8bapf4y9hnGXh8u4kaXzQowXbKBukZBh3L+cIoYOWs5lytLM+J4a+rps2lmFIOUS
9lPVY+s6LadDm67iznJDyT44xjxe1h7TLdfYW/J05zMEvOgaCXf5xRuWfqhZn8jKP6iuLDp8QjW0
PWJjyX9tJklsk1X83A9AnuZLBc8D0+zzUu6Oht91MdXSSFqMot4zyYG6iXl/tkQ+WNpmj0S6t4R8
aWjiFGxdPBqBEGe4OGK8YJVsglOFMc63nx/rU9fpZIAEWUrbqrBnZod4VguX3CNoexOUjr5FbfDY
yhLuuFoWu9PzLyJZw7+CHSh79qBge9KpwAHp8+M8IWhizNDP4K7kMh12E6sFIj7WkuXF6PRRMV1z
e9UF8z5Gt9lSeatY75DKLRzQRVhqFtftrWpD51WVvKURUGeyGobyNK8RYYjJQP0/yLGrI3wjqa1L
b4W2vmtg6ljgVGh50PLyVlcoKmOpJJBErtDynsZNxYzZGAn6elCFRT/gpphefAahtheUv61ixO3D
He3/8c1/yYKWsuPnAjLKqayF8s2XGGSdiRDx0ZBxT2XVqUFTvJricwzN+UPffz5S2BaYxchYxQbI
5ELLaQl9+EFl7r+/K2kcF0kam9eeJIfeTtb7W69T+un0t5NGDLE16P12+/KNm9qtwqNkhYlHUwHw
ziyR05TxMgROozqAqtC+uPwz1Fb4kCIDmwclQNvBrRMlX0CwipG6tyZ6qV0yKjbaVEKXThMwoiMu
ED0e7nFeP/ksCFhEn/vVVpa5v9KnPjWGJcgrMDpwLCP4+54kesHD4lO3HfT3jaz45MPyt49ptbgx
LsfpwBFq2G9jo3tnjDhNbGMGNooiu0wiW+Po8gGKmvfhsmT78TCoCkQaTvzWe+tUAFCXhA8rR6+A
nI/UjmuVqPo8tgSraxU8rZ9/38b+N2PR+Em4Xm+AFHMRExv5HRvAhWydAIj0PKUGYsj/Lgs1E5Rn
OxjvxXRyC3PvJ6jFBI/zs0LO/THnXSnFEadZwEAqlE3lzWhztQnGBlmST6XGfuuOWJFVeUKrKjht
bCFNX9KUTJ/IfI+KXQZ8g23tTpfrARD+dZNPvucYycGNEdfXjrcx5GsdV3opNmGLOZheLYpboCiW
up0TFmK1ZosxK6gchdsg0n5metMBFJUGXV/AMVvmfaWNL5trB9jS25aN824RF1KuAyNdaLaUyLye
Xrb4KVibAumfrRV3tPVm2GoleXC/DnLFKYeOPrBRwXApIX+cW19RhCsluAE/PGjO6lJ+8Akxujwy
gmdBQNzje/GCCL1P5YJsaBxEA9a5y6ip7EKZ/IevxuOSJMjOd9OoyC31jda1GH1xUTdUTxwEnwbm
mTJ/xb89UkzqlV2/1FGo3Ud2xgg1ybJy9SeMiGQKojN9SLRUGJRQG6TIcTLy7eHh+cUrRzFkMBUU
jG1cX9uLJ9n9YO9yWCWuGhY3Jlw3VApksIw5KN1XqXrMLaSkT7CpCyWAw756N790UOYWyNlhXoT8
X2qwFD/UqUU34hqx/4Ydir/3qxDA1xnLZLzQz8GkpBSpkVkqyeQJtngMImrexgqSvhaytR86PWYI
6JJQyf0bJ6kHMgxswx6c3F4Pwpj8kQiY81yQttjPyufO7/ikew0A/caZDq8i0rnVnCbsz9EtKh71
AnkupXWH6tULch5snvu4dibSk/OCicZWgB19DFLBvaDlMV+ahSul9h9wDoEzZSuoQ3XeE1lbMalU
I9KV4+CqtLJkGZHXmRIM3Uf8xVBb4/KcoS+k55wrxZILhDZ97tvSPwJM7IO02aUfN6rlWfbnrD5l
vrA4mAHTc1tESgOIrYdswcIayh0yOhjYFSABn+hCfLtj0HUW73gaJQbVEf2hx5RAItXbPuwCRzZr
JmVJ8mrGbnwvMnWjNpB85L95p7oZHI7lg/WG4f/3fVNNKd6B6VfEXgMu29UjfwGGmrm6ltuPesja
poSBxmfsPAVAX3TKSA2mkeCa9oYHhpVGmJwb3+uls+Jx0idISCvBnApTzFKN3SmgP7oj7XgJgn2d
8sG56fhYTZj9OBHI/9ulfH8xopmp+wvJXsZ7bltZMMI4nJw9jHZn++n/RanWvgdBRZ9yr29O9r3S
4eFQ2Rxa2L8wle+84a8jkl0UMXx+akACfNl6vi5KKklVFZnyvPhDJsnGixeHXtWQfywFaXSJRPrV
mVlz5QFtihny86AEbGnNNCekpTpNO2biAwPrU2Tc3k6NjIAhhm9aep2Vi3EecxKeDEOoDMb+BBDO
yiUDEyZ8x4bpNog56f+e/RLzwbhif0IKFjlfiJp1fC7dlnC6LWQM04J9dm6KO9JcUC3p3C5iofya
HgLfoF5YVdYB1wYFqiyEyTeeHuoo8PWL/AHpYa3RImd2WItuAIeal+6m90wW3tKUZmEsmNsu20qO
iGv/rfgl6WGXxavrZk2i4gwTRl45s44cdp2dFa87YhwTvauMiU5NnJFwij225hSJG57vkyF6eshU
3kNh0wbfci+Qg4jea2t0BadzpnmDZGad1eCOlKamRqlrpPfPIzCVrLImrUJlJHT7BALhGvhClBIU
CyEvEeIohNfBpKtGEFnSfJT5pXerrsAEyoKI2hQls1ANbiK0bEkChvb9vebI8eBEt1p+CqQ38kS/
gXzJRbJ4yTUf+wVRgJpeeMsHxoHbvl7KQnDqMneUYGp6Swl9rlWGG6AxBREXjYaYLwWKPIn8Y2w3
CO5xuGi3y2RPpb6Pl/IvtvTqeKXojSrVEjdyM33UY9E4vcYZBzj5hMAPRZ7UkyFoIOcXH2lR7js9
YLSvYeDlYWt54XGuG3twffzuI6th1zg7z32F3VNiR0/gzIm4sH31f7F0ZDLZOei6KKbS/n06I8a2
qrF3MVcLORnlYqqlpt9Zjzc0hx2lo5ShyBPq8qr40AAhOeYYdzBpq6bxruvMbhKKT7/dTp70CIiV
9IGDXcVADQ/0jRw4Fmr+v56QU6TKmLG2fMzkpcz2H3mbfAUfpvZU/Bp0x7HLdpCWzETMrjKrfAGG
M8MuSPOIl7qD6ORXYN4XFoTTi1U4Cn14r0+Ok0WtnAmIRdgY8Q8xeI6q1rFDF85U4SyHCvEzuGn9
iqAIJJ9CHM09ztz+s93ULvsnTX2hMTkC1281m8bq/zF2w9P3/N+CZ9q3G5x4Fh+DYwO/vXnezwUs
pPy9SgJCTpM5Fl4sTPiNOnMn5ltotpP0CLXSFNVpzAulQdVgiGI+PIdg3aN8iDdxXPpNyilsiwtj
h+PG8GhqLproGiE6CU00AkQoUHzjWNgi5Sry/RSOiuMtv+AdyGPdhpnm/ttzd3r0cdasaNePWSTu
oNdDEVwvSPfEhS31Ix6ifF/ACDbQgzQ8e992CWlVREBG/RIv8/NAj6N2dkVXuDkur/4YT705ig3b
fURoZ3G7l+G93MNpJHnT1GfuxFQzR1WCSpVQQle6UKYe5aamxvFpGCqcR9qtaWNJw4p9B26w4DhG
mFVzc6QqKxxQ6m/u5o6dpts8G5xSgMYasUabG4ahWl3LBEiN4QHSzc7Kpj73XA4k+ei/pl3yd/6W
xu5XfFL30LTJi9XMFBNZkzBqnIVK7hccTxMXqbRsQnR0V8dMB5pj7NTiSaGOCpHeuRRRdKDTW+JQ
bQbS/tPNAs5IqPHNRaDHu2GRDKpnGaTN+y0ntAKVYcpfl25YYvBiqfeRGhQal5OS6JyN9xKtxBSB
/ijwiF3iLdNmAm++7NUh5AMHYsDwHEDsmx50MHS12/AtaKDW7wvkp4WAQjkfVsgLqWAgTILW9FOJ
JBz8xf03q/MW3vehXwd7zqrto4Aa6twdenhf4HQez13XxAk89JQwhzPIjRMzc4Et8I5tpiuZvGqQ
UmZkes8wj6JNBDZfzbPPfw9aq0ordo5qiFivOc1OgNKd8emzlIYwpDxtLS0WLLNMowTqNNmI3fxW
l6DenTGQsX8eXwMfHgoSXcnyLUqV3tv+q5+lB5H9SArqkwsOwWNmv6PeFVUq4ji8l6J+QD2Ld5tj
Knb0EyURzbbquMgh3QZ5z/qllAg+VurJLPSrC44lbF6xPYX5M/y11O7+UW77PtWUJO7yrIG6WzMH
UYQ1aDM2uIZ2lPfqXtztjgrzds/n8xeUZHmS3AcN6kWGMspBcFPVfwThRxv4RK6kXcjGxdSheqCz
2mDqzmRguOtByK6p3xBI/TZ7hyPX6sOvPpF0U4w+UDG/QTsnsfCh+IkZWOfJ//wPZ/xYZGMCQ2SD
XJSH4foMDKNPYxazt1B7hiUe16uDS+QF7A9c1iL+GMmmbs1NZ30VNMuvP0M0IG2RF7qKgBRo3g8v
b86RRQuw1M+3d5LJFmEIsX1cRPHac9OsbdFPK+8eX2KwwlH2XbolqhAVopijK9btxFQfsBsd4GNf
u2Fncjz24EQnoaBPemrBqsHGCYhC/rPY+b0CCiIw4XAuOEKIKgpzzCZQgj+vena/V6Wwo1FKgqV/
1I5xZv9uoziw2oVzldCW7NCGv1B9ekFQQ6EwLV3hhZ33Ei+7kKLxl7ON1sBL1e99LfrsEZLU4VSe
oNP3/z1MyyW+1CtOOhIxzNKNmsZ/2EkpesWlZhq8PHlHb8mWjuI1IYUmloxfMTDhqE8w0wrVGRQe
WS43tsh3JsutGOVBXF5uAtIuGtdMWcDzViqP33sexJEb8BFiQBwVLboTWCGlvBuIWGeEE8qR6uzj
dex2xaOXKIa5amqxB5TogGxa9ZnTytUaWWZT7cS+xwLcjkQ/cUanhw6gr+cbeRcbdZptSx7KPkZ9
CWKcv4FMe6SRdvjl+ANzOaM6Y/sHtWpy0MU5WMDthHkqfz+jiAJFo+bRzDMtq50oIt+uw8v5byl9
d5girC+12H8GqEtaa+X0b9kuLUfyoiq0jpvdUBKOk1+rD4R9ZqJ/EhFLy9ThbDgCdeJQ7uQwbbOp
22ngoNda+vThhPJ08hhRbKJFanRe8XA+jrreV+gkmRAVXkKsVTnnNVtlj2dJuB9J3HyDs9LzixIp
ow2yv+HJh/AzeYYt3JKMfUVvr0W7Yql6gmRMbeRaDusPkd/pWXsF28kTBFrzL2ZTdltoI3jDYrAa
4aVAasW4/FfoyrOIJ0g9x4+xErAv4HQIQ/z0UWdGjCJ/MujZPMWxh84kxNVobJbQIkZMce4g/OJB
pASQ6kWNIyB6yKFqFAw5iay7SJBpx9G1+m1Nmn6phNlvsRi8ID0q3HBZE9X+vo7v1w/s4xTYg5Dg
bM06ClENusYJcU8SJQF2b9DcYguxEvo0aGunDXqLC1++FnpbuzK9EfWNuEIQcCgYf3vpEfnvbT4E
V/golWCAwinEPSe31FHiNwW6RxjVK8Gab8vZP22+3ACLJ8iS/3m9gS33nMk4W2aVwD43kiqon7e2
KVZBLmkhjkpFW6iH7/hINiMOmZ3eqLMvr8o5jOvxRkaIH+R7VQCiZ5mhOuNKJYrrMddAsQuIphxf
4GAkmcWJuOl0UxrhAUoE6ncob2wCuqxi9CKoHaGSRBBwHr588d3VdWuZt+1CJNEym5v/noIPzxtN
iFGKipYFo7luOYVFSgLys/afp0c/jTGK+Je/jN5AMzKoRN8WXwCnBYkqryO1mItpGUitWEJi+Xpw
7B2PpXRTtLoRaxFb2whx2v0aKnPI6wRZ+uFxAhowxn56mPXn0gAI4ou4M0mkksFiKfnn0+l1fm4Y
+rb+do1L0Wn+S4LmltE9tEP/42GfsLF3kzyRdOEL/6/76lCLacDU9cruolt3rlI4G5OmfDX48F7L
B9L724NOrC0C3LZ4zi+c1pvUoVftUGUmOuKtBuMxKPB613z7F0S18oeFqBNtgE6RsfiPUBOzuJLp
AMHNKFRrnkHmW9oI+aRtP9GPng1ynsO1UWhLHqfo/CaeX2d2qWL9HMA2Xq3O5Nm3g81jX3aO8lCd
hjz6VxSKymTHk40ccm4qJV6b2W9vZWY3yff/tng9LsMULHOWdcZCWHZ5QZ1HYjdQN1njgmVsejD3
jxzIqHDKZkCitxlMEEOGvP6Z9Hd33KynH4dKW5MACeaJnwzaf091+e5FFnnmNFKeaStjG857djXu
Hx0Qmgvp7SSfONf8MoYEf7oyIvLpFle+dx8d2FnRK+i6pfHzMtzmiMHJqWuu5f81up+VzFo+jni+
iCXD9t86oyCRIBnNun4jdK/9fZ2twry+mKrtL4jKX11B5u/AyVCcfp6zPVrbKDyUQtM9M3UEqquE
qSNgAeJIM9STpCIkAyDx2dPqCd8OG1rat4DHHZTR3BMyA1vRJ3nsAwsareCcbrYjdeOZVslIuBd3
5yDTM6ZSy1A7GgAuKFNWe6owwsoz9Z/T/77NHW3JvM4Jzyhf7qvmCD7DYkDrl1usoTmWijeN91Sq
mxZsKOLZTYc3kCukEWyS+RnNm/emZEbzj44OF6hljNzI+SBW6T2T3rVLfvAFJRobuW8SAw5eY74R
uC/1voF3qyFFNB0fx92SqyKg9ITdJxlyUC5iz16EW+kPL3tEl3+YJY6fo747WVRostHQpIom0E6G
2k6STj+eAfTxjYqRCeCYSt17pmisui2EmRq7uPIASgytNYytj9QUX7Va+72UfNfncHprdUXGEHsc
cZSE05FnWfTb7mxttnJwaMOGJOWI7xH1+dhkT08ffVoqbljC53owiAQH9rhIZlPaqekDtgfoO89k
0YTppeOIHg29ShHVrg0Oo5gH7MZu1i0Mc2ZwDHU2x8/WuiQ4lLjiMhbmzG7knSknPJMjK+IEgnWt
DBXWR2muxY2F0BTX79olKEm7STG/dypmHBGPmgJtDrsah8z91chUP9YNw7lc4/QYHki8AzRZ8G8V
cQiCY3yGQwjQzEAt03l0CKBcKH40IoPj0D/lWSb42oTsWRSAja25OnxmMJM2nxpFkg6rEN+MiCnp
Z8Q6s0lWue4ml2eaTddo7CHujXp0OPRnWUfsfQGnDIde+I6TjhARQXbXY/Ao1+XoSyuBSGJbhnWY
iCYUXHQPDSFvo/wC8bJfcbkPAFv7HgcZnjsZpxUf9ImsMrtFr7UkjZr1ayAeiX4BpP4ofLJMUYrR
n18dCqOY37hQ9NS9P/rRTwmgNsT4Joo5IAkEbUOwFPB2nOwis1fg9JkEBMd2+K3tU3cq+Btv5a68
nKnSDn6yuzcAjrNSLIn4qaNG67uLKJ8mkmeIlobpsY8C7PFN5R7wngXvg9ATJ7liplOK9bS0O/pj
E4KWIQ66Q2VcSNtH01B+w2GRVWFmZUeb48l+N997r5dMPOHQ3/ZvY1c1o06ORUEhyWlBfECuS1Ar
ac6nCfyrdeCQ1Zk9zBiVliA+5c//ZIJzQPXdOoa6std65k4Z9x6bSEJcriB4pFFlMuEBAn/0fJb3
zQm6RZ4NGAg1eSRhSt6YQbgEYj5sSOB8VWz1i0eZmIRt8juSZXRHsXGyJArYoHEETCLZa1iZdEqX
ty3r7tpsDtvtNtrmV5YCeSA8MdyJQ+yBNr5NRqwIJmJ7qHxZqFo8R9xW7JOFEBfPwPxUV9Zz+nXo
4zFZGbkmDaqkh+sAtX9vfRwrvsgvxEwvXhpD+IU+mE4hNiDKEtjto85W0SP+jzFTcoXDeDmERhbC
+rRpYetgqDZLhuwKIjRb7mQIXlohDOvToWnWb13cnp34Kibh7oBmAO1OMZKgPH9PLrqMLvP/cyvN
2ErNjKljqFjAXdXevrBzNSlgHchxCgH9wErLW9ymLp37uAXgkPaBjuti/S9tGOgy7hHgoo3HEkkl
QtN6r96r8JsXyoVCISYKnCqiwafDCYWLAcC8SOxZc75UAts+A/MI2cINe5mu0jmsKtmuKpF51fkt
mDsNG7MJfubfdjmULcTItWOsij4GHxLHPAlXq5yRoXXKjVHO5hP+J06fMWCbrJt3kF0OJRewkTTW
qyOfqAkVsO/M8ZSRg35Ept7/ouWQetA+xYt2AcsG1yqvcq17Tjj8H3Hka4YDdM3WIXfkpzBUC2lB
zThdsMNPDorPJ3f1GSo5ej/ixiFUlVmkJVPOixpGhS2aFWjEuU7TZZbLUaIE6dJe2Z7/9N3XnshS
Nh603McI3DpVZosK0rK48Uw0RI4uPRhb4wHJo0u6YjQ+1P6AbcRFY3rFNrWf7RfsTXHM0lPRJIJl
RwMn66NAbKlC2xKCkxBENSL0Z+7AxZ85oOOMMYVPXXPIjt+9xegwDT4z2bes+pzPelsyUq+p60Bt
cgj5aywxtgddEOZHCtFwSlbJhpLiAGI1VM328EpMJG+AksZ32kVhm2SPdAJ0y8NLHMOU8ZJ5wlxE
NDlAOSSn1/GUBDeT66pS2nPdarYkojIQXU8ADXkH/L5BtPZaXELBh/Ewawll0NgoDRWnqGPR7LVs
MvRIuiTDcnyvG90flIZsAsndUJ2xn8UzbZjiS6sddDqlN26GjHh7a0EsXDHwVjmLKt0DwCnlw6+c
uYEa8WtGaDpfJLIgKzVVA4H4kxtkxtqUUHMrmnEC3x3EYkNtc7MrbsObGOYiUOcXA8L7xHLurJ1d
SyW3gOAgnbMtqG65lR0exVxgB3CEWZvfg+3AhB5qQAjCSWpLwErkhfRd2sJSWMRIzpyZy65rnB3K
8VL1qVDGHfXF8U8dl6EBcjDVpeZhPDfXOXSSe/ttPZEYLnkSo1OiNYFgoCkGmNEkzHD8mO+U8HOz
m12Utrm3PMTZZM2xUFtgMjc0adTjzR8p82pVUx/yFRhx2yFvy/9U6Cb9vCtPXQ3L1c+y+JoGoIa1
Bj4zvJLAh8ZJFgpzR5NQXingS2uG9OhrbPMRP9NKPNDeJqdIYOBJaraUWcpbtddGHztXrjmUnsgj
8EcsfTUF4lr8GvxeGfw/bssSYYWn5yix4q5GG6QCk+t64nPCZHNFSaQS4q/Ic9akjWPLinOpyM+3
7terpkzUCiiyMfLowOcfqEujDWqDOg18YXrB1kNNZgth1Wea03/nYukP8z6jgiNcV4leZVfC5epf
eHe+/YA++nMnTwOib+NFSKgkbcjcnKyYg5V9yjkSzjNSPFNv9YyF8gHecE8FUuXRQc65PfpDq21c
047xfg4zxQo7j/lhoktgU9DQVXUoddUYLK6FYARVEJBnfRfdwREVYua0A7siIud+aOBZIWItGg8G
UWAQAoW5ukNwBCis5pwTYY11uh4WXjkqzGFiqolNA4A3G4jGp/slGTUECIcsUNiAAeB2hjIl+fC5
m8QNRPqWZuEHO8Y4Lb2FS3q3dStPJUXfpV0wHHRMMuKmM5yIBnQ8eRc2KGMwy3Bnhs5gOvNFwKNv
sOrHBureBtJePjzTir15S3HwDxUpD18vx9Eo8QoVHxmkOGRdcq/GZuca3wQ53j1hFj892TXfGjdj
L3xWF3BHZXUKoz4AWzLqCzjNKZex/TRbNLiH8dqwVYVG4s0GmxYTzSEBLMTzNUrvBaEgxlNW2Vjn
/pdgrVDo6JJ6z7UjiwIAWkBUEd8V3hgvbRqXfOQc86D6uMKdbj09nkv/EOWO8H7VVxadLlJg/lxI
GbIKpNdNvjdFbpHjczkAKkQ9SO9uXv7xOZfgmFwMU+m49H5U6cpOmtS1FuPYWuaDAxwSXCW8RDpi
nkynqPcgFQTktwx7S63mVQi/fHt4xPzLyGJGEy6FsPgt1EpE108Q9hTDVdeRtuRGp8BqLOQptAFh
T/++iRgRQ9Z8BZva8fti3MBN8T7TI7YoeA4MzVvYLnPvolZxwIzVivJtjDsODpPunXtAqBCiREeO
z07h3sPc3sExTybH+D6TIdUdZ+ViJI/u1AS4IkPsWMdOqg0JKTzGG2LZCslsM99N2HII24iARAld
Dh/mP1Tih9+FgYn0GACGtNUXsfuLVCCkvlvqTCy1wmDfbGobTHfyvh8g858YnEta4O3MI4EBCb2E
NcwKaa0ekn9vamnAWxvXKiMQlMuagBE3VAePmEUIrIzWQNyIqmA1zMe46+RWjO9ex6FKuiT4bnY9
siXDEFQ20MVNDtVBd2nZHmls7FNe3sGTnkI2GguJ4lgxNmT39bSed2qlJSi+SqTMZMAfvOhAOH7Z
j0ONBsP3y1JxeAFo7T9xZL6ftffs6XTN8dsR/rgP877SSW8HADj1rPvErspNqRytt1h37YGVN8KL
ODC0igMwLAFOHLtOoGcomHX2DngRDTFc4f3btixtfOTE2kmGJuPmvdwf9w85fJChB+8+Ekvdq41t
zJBvw1V8HQN5RV9pgaML3yJm3WZdd29hh7XbJ2K+Y3AjDGh16oyXnZWAwL7PGlnzeHycZ8l/qwVv
M+7QXAzq5TVJqwHeOt8Rkj6uatoo5mQPUy6r9d7WC2LFFC0N1iV0pagj8irnmgyAt3yElYwLVzbM
7Z83CpbN0/iNDxqVTKl+DSvVi3a3P2LTCuzbT48Fegu4ksQ/uxgy8uhAbwjiH3dhB5sJV39s9w5m
HXGI5m0nbR9ZQ2u/N075fROqNcylgc+VtTiLOAKSGXfbJxXoK32X17pALe4EYIsywlZE+Ndwr6w5
d91wZymyudRsZu5GyzjuA8hfYusuFxVV7WmVaYbSez87uA3GkPS8krm9fNmyn4K+s9KEIYNzrRIC
Jpf/GqtiHJpIbEnBvVrT1eyPtI9vXSGLDKZN36RQ/6mConP0ZGptd6ybenRk5Sp68CIwim2NYxBs
lEo748bk6RdqSRaHYH7sRnLIwOyh96dRaeXnr2phfAEWp0Pq43yASJMVqeqDY+rVlh4qHeDv4Rfx
I0AA4PMpVnYOD/XZeKxr2B7H/2gKkSj3gSMTWQA9zxhGHY4MxA6jx01zae3tg08xSZ5MnB+he1Ez
GzDUuxt0jS8XXTsDvxdlB5uK0LvkexXudsCXgzfECM+uDkI1+vaXXxVNcSi4LbNsD3jHm2RDMc75
yom2MPu8Va0q9BPNw7Tg+sywOTA7PVVIOuCrgBJIF6YICNka3eHSj70CBSLxrOpX2Ls3nhyLatgG
75BpRVUS7+R4ms2cGj4gAmwn/MbpNJNyGYO9HI+F2m0+xV5DpsZV6wrRNegv4xsEi2r8zY+79naK
OmU2kJtiU1xZCzw7d6VbvgsKGmIE6C94mY2YdDH6vJu55dDDYKTwE0kkw56dkGjeV9yMzoFUBGLG
Wn5LaqSzsJAM73Eppe8mjvW3K+9a4qd0N1X3AESG+Hq60yj++56EFf01qNkD2NflQ6mVYWGtMcrt
S0M018SxB2NLlKR3JOe/fIhbUsdXAn/rycVb+Wsh7eF6W3rUUmUwqd7QmCJIUn/R3gEzVLT3tSFQ
hlicebngHPbe2RAlm+n4DOpNFfycbj+XJVeesz9IpUHufgfoXiVct5Bt0edeFPTK9ARYyQkKv2ti
GaoX2Xv9liZCXt930wndTEZ/yppRPqz1W8wObYa/PR3S6FU3fkUEBg5kDCrWxo5LhuhBhFuK8Dvx
B/obbRW/wjeX65lXPkYfL7wAOmxy1bgbonz76angswFIXB0xD5YEUe4wK07iC7IPG6q6Q4m2Kjw8
i86teW4Lb2cpWgj5tnwwN/hxbkCE9S2MJ1aC2QXevMFjXli8stSVu0kne8LrLWk/pgmCoIunI3sW
QYWvi8MbZcQfTvMhyNAEUzTLM30vciz2OCr3IaEemNyuSLiBeVFS3gaRWTMxBaTRt4VhAxFu+NW8
uMMFS0iOWUg2bXRgRQnaHFSoEBXglId9TpYc9d4L5vIAznHuvkAL8P6CtviKbv455mBd6yOax6Zl
LFXSC/AvrWONobRFqHGhUcEvEnFQaYkF18Zu9XSuk1oqzFoYGN/EmdR+lhYBw0UBKtxr7Pnp+3Q0
BxK8DJucgrsQLK0FTUyswWkoUZ4YAejxrJvcqtF5vTfjZsGBzW05BuB5iwSydYD1nQkMMm8E9mtq
Rg6nE1hr5xYNSuwGq9xl8xgRKYFFIzxfQRXn4Wrn6QM/H/mP0NA+7o48wbee93BDkatAUtijftIp
Vb08iAxvAN4f/SYlMjg+tLyVQM8wGEL+fWZdJL0pdlnKGn+hMT3oLpdAbnbLRazVEbUDWe8Rfmqn
GmUWEHkp7IWky8EEpBkrwXyhBUtC3Fz74ZotJfRAaSyyarvYktWPfmFeNH+g5x/82UPjiRX9NG/+
cHItQG7i3Zt2kj9k3rMLlWafyfOBdTB76R/phrjrZfsNa9k42V/9lEmXpLY/FYeKNeB/mBWbsCjY
cXwin1nJY3Z0fKVWqGM+6kvEl0zIzyRCDfSCX3DcZivT7AVUjbHahiPPBZv4LGNlBltCrR1i+3vh
ZQOtl0Dn8EwfGIdzxPXaJmU/GQATmRUHEkEk83KhvvjOnCQMdTh6otFEblRFmsQNVOo2JwHfHMP0
jt6cqaUdq3INuccJRyVflzS4xw5O+aMi3F1VGrigccrnlI1khVbfwU0fKkv0UOEq7GOtTDe+uGzv
wxysd0fEjtmNgTaqelgfBsJbqmpGzc3TXjnVMUDlE7DtNBvkI/7Ig0liPzfUNP7Sm3lsh8TogA0T
lndTfsJP0PkfTV+WJRESwQPxLekJjw86ZqBCiOCFDc7499w/wb/kW98ES3DIOyjcTrIu2QJqiXSO
ueinBtHBai2vcaekhxmgGu/fg857qKrDtF8uxTThkA/E41DuadLqKNfPlyGwDoSw8tHAZWnTd36G
DCz/E7fi0OpQbD97WlSosolf/pKxieV5rIsj3FeDY0QFBRDecMU0hdAsG6ry48+jCq7QHDgbzfKJ
IBjyg3kOhgS0Kh6RXN5mzKWWDueuFIiOVVR2epMop9ChEgzX7Okl0HehLvSnXS+rpJ6RnB4BBHEX
bwktey1klFpVAzmh6n3tgmhWpgRoJ0Zurz/SPvgA/1oK/elTCyYRLiOZAKt4lAoz9Nw/nwxSsJ/Q
wuSivewFM9Sinp9p0Cn0DtlXnqvJ7AgQdB1bX+Y018D3Bisb2CiAsZyc8Ar7e02UlyWJPulmpnrb
eLXpxsQ0SYRABeU+Uk0EAZisqFBrfR6l5mMS4X3gdZs85KJoCK85xPxNCelZEfepCbhT+gZm18kD
e2epD7I9Bi+4//taY2x6Fqn0JMH0JzH8fwIy7g6pZfV0zdosk0LYqz/ucgskR/jrKEzEkENw9LlY
XxcZIrRh4NsgqnWqdjBzI/8iOP+R3WBC9IA1iOw3/tJYLeiIIXIl1iL+2PEcNfZw8ChA+5HNYcPi
37CdQFAsZq9hAwyC6/z8KLUjC2+LBOto8tyNTFzUycKV6V8c4NRlMiwfarqvi0vanZsV/KNqe9s4
+WJMWJ17Tq3ZSN75aYtuaN27C4r307UpeCIIxVBzc1e8cm64GyNgNAZ3cbmHNVjLEzGhHnK1XYDO
7oP32XT1KHCCpIKBC9kqrvdPsKP3xFebmy3h09vtItcB99bkTRL7RPmBPwPpWgzjJ5VFfbVNkoxt
vaouUQEAaYbmc8XcIVabgKCd5jZGMvwP3FNUGlpZd1ibrONqIUgJ2wQdKfZ7UBlv4O2gZy/0Rpxe
3KXd9xF/At9rOuTBAeDxof9yNXM750Id1/hYGHzeZIYHlX50kkMQuZ1Ck4wR8E1GPTEHHxAyUbYK
JAh3aAQihDmwGMaQBCvWPyU+vcAa9ftTpwfWV7C+rPv5lS0DVoB6njbXIWSB0UvfiLS3dwFHzeDg
trkpieWKPXAoeobDRwINayGh1rsLJ7OPR1EpgzVic4Utf/4+rz3CQSCc8/nTDGu2baiiZR+teIZE
qiTbOIsy3U5zJ+3bmQvk/8+Pf0ySVFF0fJYjLyOe+pHGnYu/kBRI+oXHdlSCpzA+c1D6So7x0aqN
F1HpiXe7JU8zUj0ikId13Q6vuaL4Po5XU6ratSeyZk6oMY95OmuSYctYO+H8LsjeFAAM5xojl1wY
ROFh7KO0aB2BtjCnX5u+nIwJM4ywPA2J1T0/rmiKdtfaECvLWEgt/GFK2/hNsKSRcbtXlgJlruA1
8BoFNTUof+ambeI/UBToGAbDa0HRIqoNUQp58U2mRBnFF+tqPBmLBArcHGzw729Gh3MqyFcZnmwl
9u8k91O4oIHF39E1vxsddQzJhCvHmOhgzomkfHA624QI46cKWQUO0JoZ5e+Qqdag6soxqEYJj5mG
VxQYxbDfqDJ0QmS/mLiKGrIqaAr6UgGqOIHht4bM8FEHZMC5OGDvS+y2yucn7DboUNVNWZs3gWNI
RJlLJ64b1Qlr0U4W0tUkK4NBlfmcl1ApP1AenKInbX+tS+3M/eNG4Vjqrp7H0ScNdxYyHI4ik/Ms
Yngf168Ri+TO7zftkvmxBLXu4Z+tCGIzg2fmsdfEX/frfjzjG6GBgYCCcgWm6n4u1B1iX/u80Ae7
F+Vy/mQpA2LPxWQPUvpEgNHVYuQGK44zoxqvK6Z7ksf/J5YL3nOCkIyjKXu7Lq8+DEXMU6tqnQdz
PKgSZtSistju/1/mNyMuGqY98oKmyXUay5FXb2yYF7PAhB4U9WbYyc8b1qYKuPFce5+7lZgP1I9P
8ZGSwZsagjAXVAQ9uDFogwydXvNgH3hKozYF9w66K7dGVq1vQJyzBE4MR8+yOJfc9qdyIuonkBrr
SRBWKJNFZdi3fnSwQsoxPUFfKdkWZ0CFLfNi4Qo1oZ8/4qu9YgycQwH2e3W7kg1ggP6Pe+fcYMEW
YhM8X+l7KGjPhdhRlVNQE41zrxmcu+37VEGibsyNkL9E1qMyJhZtwNDEacRH6ttPhfpICaoFvD6Q
7lcpY0r96lH+PLOMY/7nPNt0/ZKjQk+uZOTT+q1rFpqiKxMmkbSfP7jlETWkNrjzj3eoMVWiZXcq
2EhvmxRwmzI3KfbjkO8+pVOUgosc8OA50yNtXuh+y6pVEHa4KvhV0nNiiKAz/k3+VsuQfyP280ZQ
RZ/ZTyqeTh9qBy+w8D/FmJc7YyO9M85qMJGJcqkp+e/yZbnmY1VSCNWNG7JPCNQEDXn5RhIAKiBb
8O+Vly/9L6MNDA6WLjDfYqNkLrkRegNP8k3tMNo86pGJLCCRFrMTD3O7aOnm9LlhSiSWcXTq119K
0Q7/MV/lQ/vgLvJFB8KqQW8NX4rGoVB4rjG5EsUWjrzmMv8qFhuDrQIde6NzgKnnYhJu0ib2ciNv
LVVQTBOXX/WDuGhWAFSq1XZOyrKwAOTl4mdzfJnkqSoUwnTsR6Gmpi5J2559LWLd4ZVFlQyGIg2+
HgmAWIvsCVtIKd8JMxTX/L1QdS2f82fMOEK/N2y4vGWqqcI2G6T+UV23bLyxlciHjmNmc95GoQ0V
E1o4jOFAR9ZsnIJ2Xf6d8WZBGQ7j+b5dHZovRzFrVZbZ3IfMOs94AStH/lhtXk+PDwfa5+tDF2JQ
3+RruvLsKKjbl4IHmMHF1q0rbM1h1DfedsiHeVOfETcVM5oGhzEGS7GgkMQpNjoWw+oSgFEPvZyj
OLQgA26V5+TwMjg9TlGt0VZKsTrPhGF+IyxrPHcHIE+W9Uj9X0IknY86r16MyVt8lwAssUrT3/KP
73D9Wk9XM9QcnSeFpA/V40dxUvvW2z0oYnGvPnVfaCuDoOTIUAtrZveLfXn3IOcv92ZbbTAOcmrq
8HBWbGw/saYcUfV5brsNBq/y/Zb9x7BOnJH9ypNQPNM92sgPswn/ZrtpxNHgZU1wC5gmYHqYZZhd
jJ9LAkKv/e1dCLRgmwq7Dn3JVSJtLcM+r205W5yCzjd4gyio9Qd0PePBHU4QTO/3aGADquyrqIWF
CcCc9yZvKFNAS0lD+0CVSIpYrYVbB1ZrZ5LaAFpSuCytjOyGth3vTYHxf2dnwDrgYESn9RoeKOv7
5jSOZGYDIGxFvtGEFboghG8tH7Ex5JBZVEaqpOJ0XVmEqMo+LAdomvescHfsHbRR2DqBsLS+R0tK
PEM2hixo5nFaF2EydDtYdtvWctFr0SX6Y3LdTIGrCKu0O6CNfR68N9eUbMTajag2ZJ85nRS2qU/J
f/gQsk4iUfk3cbQZ2aF4zRT74A7cJyCbiBLGo2roF7Z4zG0eVWIo01ph2fMgHbY5oip6Eoj8lyKO
rASHkwx6IdSkRts13RvD0X4F+34dDij4wJ2KhtnsUy0eq+eS0bETu5FL4sFZVBXWFv8s2TKlnMCq
9wbetfISas1cEoQvwpHrxIB/kRAaR3FX3AN2W5lHk7IL0VWkbwdz0ccv+lA3YHxAH3RNOSiJQ49t
M+CVHjMJFtEW8iG3h8ez84dH5SNAZfbXqVFI3Jl91z4W7HSgywuk7LTinzhytLiW28pnrqJ+EJYs
Sbwro3TH5H4DEWQWPztZS2kNtlbSS+2elWEy56TG7EKhvS6TXsTj1WNFZtj/EQRgLSvnPtv6du0M
Y+9MMSfLhX4mHQ2QoxLp8T7G2P4pQp4Sm7ho5cANVmTosZAD+XyjYkSYrQkbUO8d0FDw694dmxKP
Ze1cUZIxq8XDp0wtBCTY7P92CTp4s1CNjQuB1tZbt2LwCOEmD6HAEsmxbJokrfMEn0zQ3JZNfB95
oufl4mtHawGHj9gZQcC1y3MrH4s1SWp3nuQmGbyvmsWVG0bQ38MgsSNo4GXrnzy6o2wWGOa3rajK
gsXEDiKQabrJORFrI7Nai8GMwZRICitWBWd7uhb40XqXMIu5Ak6NqpNbbEljNp17Lw4IHLqVDJD2
Cgn8GG/D+gopBs4+Y4l+xG2snYzeN50ZRJ+ZenByXaJ9XsTtoC+mvbwCRhzeJuqPJj2RU1t9XTcg
rcVIq3Jh/LcOUE6Z/quAefGGXAojbXU95qILDK/U/8CDuGVPF3nC8fzFFaM7ztPm3AOfkxA+r7rI
8DIVOlCav2Tiqxq1tIpZLrrg99f17cZyQktRKKSuuuW0F21QANQqxm/S/Pj26vnpeL72C2ihjXL/
gDLvT3fuKbhKAQY5Ipb2fn6LTl7Tm/v0TM0tAFAz/4LzuC4Vj3MAXodxYlCS2UCyNubOqSs1iiin
j471lJsODuDoLotOp6d7qraTxNIvRpYYg4omroCkUfGRArN+koaKL+4/D6n/kNuDMK4C6ZhH47Bv
i7R2e6o2ICPc4wK6UdUOOdNFzonVwAWWWJtjkWG+tyekZBFlpdkFAi0ef0KWeS7jVPKd6FJ3nxR8
MJpnRrRHbgKIGxQR4z0IG0EY9s7aOD0LsC8N7C045x5WptwKnWx42Vw1S/Uq+mwQ+s+e2JXPNToI
PrzsFzeRmuUGXqCIJM03j6Qv2HMiFlBZnJ5VsSo/F6TTlSl92v3OqKG6vuiYE6TDQi0fqonIt7uv
f+efqYl+/LoYBCJMB65n5M2Z7icXhf5zCmbcqyPbIBDyaFMew70mWYV/GeyD5ix7/F6IoSJ4gz24
ULLz8PaONFPwtstfOykNwvm1lrD20gO7Pb1iYiyiWLeDy/JXmmUbAiR/RyEWLZB/UATHNtZ9Okyf
0WaBlfU+fLxHoGVfmLBEpDrbYd/q19q26awn3J0SIp9klqmdJqY8p7TJcd4RdMlWiAxHXZwnmXP+
9FxWCC3rG9TqF8XycImc7Kl929UzVyf/XjgCE/8XGtStRnQ6fd41+kFFPl6GBHCftIniBE2Yerr1
3ZRDTUHw89Jh8eTviTE5lzEazNSy9TrqecAm/I/Om0h0i+xsZJt3PGjOx+AM6ZTGdJAbRYHj6Iyr
oSvjle6pOCbmdREXhOQ6/SK0/V/ZHm10CC7tVfe0CbzKuc5qP1q88CZG5iZNoFycqb6S12PaBwb9
SFu3P22nuvfrgRvVfVLKree1SDUbSxVyXPwKEf5KxSWNxpCxFfF6v5EaMAS7X6BqAxg0OY/lm+DI
CgiF8IjVQBvMNeofTKJLbCt6VuuV/QA4K0w96ohYRHXSAV9RLGkGsTlnhPmOHK7XJ56bsGR+RNYt
pmKLeczTvKd/f6ePqMbzJ8uIC1otFfUSHGDGA1+/hENORug2iHMkpbYcQjKC/H7m+8+UiCC2wAwI
K68VvdsEsa2Ba4eStKeFOCr2QI8ctEVJ1VhS3F0/M1PESUdNlCEaOGi4R9nalfb8Cgw+/weUogMM
eoWCnJJiEmuCJVRRGPO5RQatdPuZuTuI4OlgMQjyK8F7SX/IRYKKO6oBtORQNh7U+HL+9yMKzkke
cJdNH9Ga4ww4dVwmY6kOqOQnt5Bl51AI5XiP8O/Hz2FQs5ya9uTkt1j6hPiZvD9e90oThpb46OpS
2HCVBLajMLidQ6rzi2EYlvciHmhoIYgNjfvp5DzWzCemGbWFybxsGF2/0+0shqdGRg+fWP4SkytO
OGJWdmC/rcfSPMvK1PME637ghHGlhEuwdCuKkeMmkndtCmidM6jwLmg+SgdfMufgcJk8/Ubxl3Vz
Fi39bpHJcpnzZn6tqC+rIxVgWrPyy5WblYaJnw56FM2sAUqFKmtOG6U7JVRNKMTGLQK00dVVujiK
9GCU+wJ4bzsdKyZwUXEbNTGwNTwuwR49GBUuaYa4nboSVcDao99vJAtFn2/yOcDyMDy7t3LVh6rp
ztC5U32OgQpCqgBJ2wHw6NzilX6ignVcHGAb6E5JNefmi+sLrEPfCxZgVQg5zMWzcC+jmvNHwx7m
Y0Rlb3Zh8Xa174f2mXG8IZe8l3LEhU4nxM18A8DOo4oPLGRSwytZoobBm7HU0yafragau9lqLFUC
Ng98CikCVdWDpYzpQSloXsrUeKKM3RJhU/mU8sWo5e/vLyFMPl2URXlUf1w+wQld8XwA6XmirdFu
26/tnCsOqq52Rq+AvpLoOeBuAK38qBKJ1+s5uwxhpXmqAeRzhgxXdP7b84j0ryL/3IZ71RXWISDr
+f5tDuiTPxNqewElb+s1cJJpcU2+834KH9LQy4HCXMh9k6eJN2CTTzdkimBoJyCoot2+8nwqvxWQ
eDNf+L1qL7W76Mok5wabOn7yMxy+1qdyslDXkk7omO53tH1HmjLv31msbkgxeWbJzuBe2COySgay
1+uwx3Q1NDJwiztYOgde45yAnHSqFhP37tQ8/IW9wKRdtgL6zXBqpSASz8o4LoYSkFz+nWZGySz2
GbqEPKVdA6v3we/ti4eeG//Tyjo3Aj1CBbKTyUB0aYdxrwJy57WGW0CpnWgGVfyun/E/iUM6lG4D
EkSFfNaZ1+2+7kD6pwoIQQQMSUDzhOZd1TdOOjJj9nJv+eVepgQko7oCrECY4ivSqpAc4JuzioVT
7zVkL+p5xZAaobQpbqdAreDz3o5W28GwnsEQfi6yxVMRbneBlcvUSi/jhJyV1UfAhSy5JEIy3TCY
Z8WbAUQaY4SGA+dKIydBg85RwqP0SC4t5Y0rCVpE7z8opjNzh+3kQmwm074VzN/NrkCS0NFHn1Xc
SbONjTbjIq0/Q9AH7RLOAu2osjhQB0CGqhCpu6kQn3CvK0nMMtPUaiuotaxv569Fo8RUMZivoUzH
WC4rnVYUwikolMIOQUhkOz4ppdyz4Xh6qLl6/tyOGbuot6DZz0DbEZnTDyoq6fVo75EJ9ApGHcqf
lBDf7lRsGW8WwcucV20vq2olz9zYmysyTGGpLkYy6iqdUWqwFwiqAyuE3nodi88so/6a3tHWjaiC
VaGn7cUHrQTZILFvaupujd4baDtlRIYRHY6GBUaOdZoLgwvFecZnzmNXzO8Dcg6JfQHitim76/UN
Zv8zm8V5a+Rk+lCC3Yp0xvWjbDEPum/o3l8zWuRbTGVgqNh2EJqj+h97rE5ESsDRrgh/2Bz1PSvf
TNy7VINZLymRKMp0Q1k1Eq46NFfK7N8fvS7NfX7sEypQQgcwqKAGXAafCrWpc9GxFS3WAvtjI31r
pn7OF+x0FDIG9gZ+WfWJLuCLZweDCfBGbUzyUFt5oUj9mgYjC8AdNxyYHoct/OI2oMs4s4kby3GJ
0GL5jHym/N52AI0aCjaP5Pa1OFCRbu5U4xsgc13DQQpUW2/2cXMCTcHoKa0ZrxqmmtE9zTaGYyHG
ASqrRw4DvboXJ4v+nSpAmv1h9E9NIvPgPBAMs7JlN6LiXF7wm7JBkIM+GrfyBExU+iZ6r0nReHf1
/S127vaT6LOCN1tqeVWXptw+TQA/IEIa27rAk6WHHyjkbVlMGUBY0VxSHg9rOzSsa1ZQRRR1ROk8
zL4cvFiZBkq3coyA/ItBOSVkLYfpvDg/+CW4AIin3G+J0C/p/c0JQQ1hIveiBbXwrImvQk7OCPb3
qvpHUP75LfOo5DXkji6WEUcntxe1QDveJaRmuX9/soggg+ACHeJ0Psg1lCCgmBfXIerPG97w1szC
QFzKqDsKqp4sQrHbJ5Tr8oecNmFjeSID5JZ6LU/o7FrsFVnFbjurL29ojPh4e5vC8SHLK9zbQ0IB
1O1/36MfJRanE2L+CuC3TKYCJF0ZV/IjleBMn8OrEFW+wR+2zlm17AIAQ/6CmBNnOaBKahIBnKBO
2fQaVIVakp1ost2nsmjP8FdjzrvVV///0LY4dsmCgn2B6/lpR8PdH6u+nyLcngq6scrD/BPUx87W
uJU6uHbfYaMvWFDsWtdoeKXAf3nzEdu+3HLigETBlwnVkEe8cwInEbPfNDGn7xXHOihYK72qd4Ko
IKWK+HxADxDElUi6Xus2/bFCjF6EPhOvVsQUNR42cqQ4IS4O5e0ltbrTzBTet+MEmr/boBMWgyPp
HUuKwIiE7VofS0Tn7NavEiPobbkavVE792CLEUgvOH3UNKWR5XfE1bfVmR/dtob0aD+ertisD2O7
QgPpMnddXD+5f1WM5yaxgQbQAyFWQYOqo7XWUzI4PX0Fnc2EtC25Q899wswRkjv01BQ97saYjKOi
ubvgBZCf/rQyPLyX3LVsiu+Cd6+/3IEJN3FM6+vSQE2Ho5J6neZ2dUnRx2JyhdLQ6jMMSOgqW4U9
beI7/f3OuCr3SZLQqZilibu3KvjwhhBP0Kb+lqTVUgfdKZzJQwX4lCzGWwdIdYHtxkiIBQ668NO+
P071G8azfm2ytx13PtfgzkqJJTyavye+uWCgJPGUZQ1gYwy3SirptWVfHOUxuxrFMvKZ2PpFMSV6
yQvxJ56NLGtwpwsujWtBKy4MXJANxamwxpiRTBmG06GPORMBVfwksT9JwufIpNdc3njp5Up8d0hE
NqvcfF6NtR3ziDsnd56XgfwIJm3KYH1ciM+JyuAJfV5oAG3F/Q18OXl7bDQdVEJV10K/J78OHFgj
oBPoIIggndBI9KUNfAfk+KnFLkpVvDQYgo6YlVh77knmaPOYh0VFzPN6sxbWAHCxlYBLswi3kBNK
rLuVBRIi99PhAhBxCVT1225zHYg4d5IxAJdW6k4+mYX1Zpp/SoxSVefU8XcZhG8kSDXpvwmNaqYJ
w+qPD2SaiunBDgdwR0xn82+4ofJXRhPlrDDSYnFTvf5lW9Ctw1spLcJY25+e3jseUvO8dZN9nKYS
lNLq8njQyAht9yd5ghSxKFoJLipXXY41hlTtQGYaB51L1gj7Tfdt5pImGUtHoNKtPRPkqtTABWT7
4bn+OFyWmVSMYWrNu3LfeOi+YtrJ/BjngGefAH4DTBKpWgfiZ/G7tuWlt4fvJoY/SieYpA5WtZoo
fCplecunhRWjFdqlbVXvCM35S5wjnhsvZKvAfidaZc7UVTDKnF084ESRWHnTzfp8tnBbRia2U3Jj
7nWzYfJT/Cvc/x10sF4USW5P+nZkG+oYh2yz6IBk2e3AXqUVKfntJjNQp11bn8smvdZJ0i5CNsM4
iI3eJYe+xSDXDlSL8dZ/2KkHRmjAm+FHRdMwSU7kpQ7eZQ21VSEjb1uhLDpqZTJDnlydhzMhgtWj
08ZvDdQDmxOWbyEdUnb559oFgIMwWQdE7+eH75aomfrZOAyoY3G9g6mn2+rxHVfktBAhpxYzYYpc
KdaMfK4KipQzuzyL6+reDEfG1BI606Rj0MNY4t5SXNwiCDRZAMSTc3znW3vWUNA8bGZN0g6VBL8D
RVtFmgH52/WPpgswBK20JtRMdO7NBvONtrUuwk5D2pLM4qZrhuiW0a4yEE78dNQmzoovNAFyonXI
piaFh/qFdncjvBc5jagN+VHrIE0PGOmGkqXcSdFqlGLAnLg1CiJuhYZR/Ghrd5n4k8kw3Qd54SG6
KsC+18+I3ZHNqfwbj2vL34Cvyi1fGMt0Wfnj0kq/SNzpG6rfyULBU76R5Z0pS0LMc53TZMqTAsRc
+pCgsUqgWS5AwgXsLhjVb+fal91DFX/UlF6l8RSM3bBpthUGSk/z3sPZv+30EorMzSrcrlyiWnZX
qXSikbLQxZSS8JwmT4gxfRtLq8r2irAMH0nok+yrrW91FS1lBgzrGbFcl4VrFNGn+/UFyOAMBiuT
eYFntu+f/bM46hnQqv+J91dgUHmu7QUzHEfu5SZXuBiWeE0gqYO6mEciWVmTQibnXrPuw1lxTabc
XbKhjsOcPmkAI8gblvqFYvCMOr2ej9t8oxo76d6hPaYilZSxOZ3RmfyMFeGZY0cRev6z7mMw7VSk
szQRe3TLD7leEZXp2lf3bPRe9wmKn6arPdFqhDzYN1tZWru8SKoG78sMyA+dYwOO5ZzLm9IHxjuE
D/ohzkZuDwuClOFiGsC+6G9NmP4U5kCc/vPObXOfipee93ZE9A8pnFiXi6UXmR0Ffu1tCqPzkGaF
Vu0PWKkb4BbBI+Cf5o1yg+wsSP3vnlahv6ddGYfWZCLebqSwaufVSgS5OXwZ3YbkwDrlM+NAMXsN
TRXyuX2izLJCnIu6EqRcE7R+P5AbxZIp4wBv16FcWUKPD04a91au3je/AK+JZeR+LHi46glEqKs2
VQasgD/yitxmWMn8AowmaN30O58ayS+lk2iqMGAUZVbQ/JgB3bewREZzmIvVCjgamxyFQHtROjLT
YtiSH25LBiYF98zAApXF9PCq9Y+wWlAeBtZGOnNnXMPFrKSsAI3Lc5jyj63nRbJIQ/NhsuXkEgNf
LNE3w5yHqq/TlAkhPLD268oxoFicQTZ6C4+/ysuHblHAWulrzyAvIiYphqkE5LTLdi6F8KIcylK5
3gx9e+HVALznTvy166vDAK5VLE8K0zZworfG7Ky89ikv909wwpwuge7i4NWlsrhbt8DU7y/HFa2I
ps4Bb5XfC85U7+1CvamRlB5eqCtM1O4h7lz1y4mSJCwg4268uZKPKIEgy9DWaDkJEE7u0/vJqhtY
dUsR4rsjyxCV034RclS1cunUCdiuKb/Tdj3R5GPco024E+xEBVf4thROC8OPM9D6ZHpLPApXwwhu
Jsm/iOO5o4hZLpJCgr6FHaYYWAWYhlpXaVFRGz+nAMmpbZEauWDKUdPx24zjei6n2q30m0WgzM9y
5F3U9JzRrUS26H/qwMIZof34HCfmvZNrNCYE/0CR0evrjE8tUWtYWX1CZy+ZtsgMF5f6Wdb7e6D3
i1TeO+65rvu0BB7olYKW2m9ZKB/i1T2R+7AHCPuuQ1/1iv7dxVoVyr7qnyjRWiC5W6X7Mk9b5EDb
aDkC7z91NQlW7ER2gtr1PxCauEIA+V2sTYYeJrden1lNMPjlxm5XilwDQhpJjsoq4hub9IusmV9s
K8g+bRq1CBC38UkLOMgByoRvE3VLtZWjUuJkaOIOTBydSx50RZpWwLiEX+MXmtte8xkIU7Ve+fQf
JxGMl1+gWqFNAa1g7Ue+DE6FoFXVC5txuo+GeB9ruAEK03mFGBhGzDQl0WVbfAufTQuFXxhEA1Bm
p28ZxrtBLFIAHuweSrybJnqzP7r3DLdTLxk2p7lL1nCPG/xtH0uPaDdqr/qT26d4qLPnIJQs4s4n
A8pF55+LE2qeqo9uy6Het2s4RFV/gZFZu40N95kRZ/0Dm6eF6RCpz6uDkYqCblwI1Rrq1bNcn4n2
v/kcJ80wQeNdOlgTVtnOTFB5C+U1vcdPZaU8hTQVCVIV4QVRdNsE/AuHcpo8ycR9UXSisf4ZIUoD
QzIq97Czo1TLsWAiStYhxAoYDWXYz48B4XBvwDQI4+0Q9Ymi1fiKVmo0aTOfGESeSMLwwpopcuJ8
jksP9PvSzwxFh/yzpcs777xyRC0yg2k5h8ujyHv2645eM52fVpQggn9y4H9Sm19cKFdAcAYuL8zp
6aJ0S/j3xVtoqAlFiwrVCz2Da/Ij9pG4BPWXBbMAirZLaREATAKI9mkE3c6tb+9g77MbBHE/kCjv
mvFfTuMhsGXLaTIdGQMZZxDLstOa1ziE0ZSH7QMinQm/Y5r9C6MDmLwVYQpiIq4DjDVjYCnCSOp3
2YiXAQr1DVZS2t3mxcnHPQFBka64ugL4FfWXckC+atZ7p3AeBOL8QE0oEsNbi5yF8yDwwZZ+VP6p
cDrjKNm7uWk/FlrYQSPXpnGSoKlEkLjQX9RSYYR5SOjZkXNLf7p+fD1prj0LX1D9HtuaV/NDBKna
UITCzroPchvBjEl5yYRnd0pz12dleqOfSOKJiTonVe7wwV8WbqO/rtcUg48+Mie+we/1XfzZishm
9Kwew1LHcbiSmE45M/SkwcewDSmI6o8a25xo+jGXjiTMpVXjdgwOSQ7n9hNA/oFrzyYi9f6SJo02
kxEiL8etFwyZfOmoXoCDea8b1iww3d7IHyoRGAA091cfsPCbtK/W0glNn+WpJIKrfyC+clW6lW2+
L95kPm7pgDN8UcOxpBva45uC2LNrBGLkRYrZL+lxG56nDYNVKLWZrt3jvbUSDawuUc5oQm/Nrqe1
hNPi5pu2t/DfrEqv4VNG0LWYoSSqeY+VqZ1WwB3e0Xd3ESRK9zoMGg6nVTyYwXNyCx/gNWXPeMyc
DRtpNOINQ3Hxe9kJ6FNutkSvBtAqL7mVo8iARt7d5vKKLDFXunypqCb7RBaIyH/MFaOzY2rJU9J1
9TBcpbgh0Wxot0UiUKhWWy3Z5O8t3kccM3UPFqCKp4t0kX/fhevOVV5ccP3ObPehSc23Kv7sQApq
LpD01KMaDEiKzfncWnWxxNBLdoThBkjHsw1sL9hd36QDXG+3ivLcQ0VxkHXSUbPyUVi3kqe/pRw7
Rz7WVtVGnQVb2fP8L2IbojywJ/lEgO0We/4YkFSkN2eXo7BQiolxKxOATsHveBlEfuSCPMAiNTaQ
5/oEUQv79i1s8HIIz9O3oXqU1UZ9Ong56y9g19cHlL51i/o5thuccr2EPo8BG26GUOmcC1Wkge35
4VFfxfXcLTbFNw7tRwLjdgNmhSculdcR7sWPGFDqs6CtTl6tSUMukH40CYChpDHWIMhjgqCuNrXe
ZrOlUf6Kv0WFG2FtJlUK2NAKwWHkWJ+pmVqKG1BHWimoauMhf+eaTSKKfTlQsOrPcfXI3jNwT6Ft
2bdhGWoG/QRScIAnDt9ySTHtFRkUMFCV5zqT5JhECAL33XwfIlMK4OmTvsVSnuaTIZxn5X/hiiTM
qre1dxy1KTh2Hj50VMhewXH8ezvXR3jHbymO2m9/ElUz4MA3USXFTOK1LopP3WkdC6SWMdsOdInd
Sdfs6HsBrNG373yeZiZnD5Y6cH/19qgorGTYKHRFygmdth9iqyu16/Zcq9jDYDCjtxIJtgh5XAva
QXIBdlrEqobTQWZJ+938C2am+3q14gW+6ZpaGjvGFrCBT4XABFC+AZvhwhaNwKp/xc9zGUedS85X
MItO+6E5N1wvsMhAashOj835dKWJjPnuUdml4p/hscnoArncRb9CQhZcIPuhej/bQi4uR0X8955L
d+oTLf/VCdFcM+chtrR4zdoI1biCTfG0RstJfxU55nfzbf8yuEoV/segfCMjqBeAqBT94wv+PT+Z
dnJdh8DhOzGSlGhCIRI1aJPg+twR9pUurIiG6iWtxbVJmpk60Pc4xOVU1XexiqYnEZg9C8a6bwu4
AETISIu0AWMw+qv3hh6ism2M4wwcNAlh0s9nprv1euWgNpzJYv7bWJyNn4MJ+pKRCfU0HYZkDwPE
JscRDkZKS1ly60BJCMiU/5cJYHRii0CudxqiMiabYkWB7hvunJrjoR+ulPfYR2s9N6lcCs+M2NP1
89yrwxHsjCHoKNS/jzzlprErCCGz4NH2VGzwBm1mLME8qHyqxLQ4WMs3r2QUDLIgQkxiVTa0cTKL
7VnEjxOVFLw8kAlQ2nG8KP1wKd8Qt+vaaooKtQ0iLZo3+WLvBT31FvmMW6OjWD+5+MBwRWDvVb9w
RoshiQfC07UHx90e04wpi08eKNutAl3eHZOtJG84GQJtXfWF1Cspl0E7X4sbGR63R71IjAW05UnP
SvYRbXHXosgyvjxby3k9+vJQvrbFtonqoaN4F492gNWOwZ52/OgdwnMvvVkaWkSeaPvCnyy81ynX
HObdHgOC8EgazXjGRVjqqIPx95XoTot4nVzrPEmzGrErAarQhqPhOjCkF4a4/MbAeFDM57rY+NWS
QkgvCKVIAAtQQFEpNuJNNmY29N74N+41ZqLUwI4lhSG08gew2LxkBNRMWeAXLUYkrFUCd87m1hGt
kSqfL4ZF9GanxuKu6kfob9D1PYomB8Zv/PEhxTQ8BipqkUXGzRQ7fKUcHU+eY5rjLFZQ2m8xIgR0
6eoJeuIpB/r9znh38mN7p20ni5dHlAyyxZ2os9TcZ5u2/AEm6wdo9fipmlBMH+9JrreS/uxOnKDt
JiJD3hN2dxBUE8HC25hK92a5LL7qjeGBPd4UUKehkSDcFCHDkQPSMjnsiQoxlT2+UvKjHva/09uC
WIgRiZxD7KuTNIsz5Pxx4KUdxerX7M28j0YgaZ8yh6iTzwBXZ8M15v3//FUQkeRUPHprM8KlKNaS
DVh3YtVCMMVAXWm4qqhymEeNsTee8JXBKRIfBRCXbnh+MxwiV2scEnN9qVjnVlsfTi6XkbbjXW8z
wtX/Fe5g594er8H/40aHulndHqbAPin03r9s/OCTnZ3w790hJjJAtqavzv4RKKwNO2iUVFXNDy+7
RlvJvKTdUyoOkNDFqaSjUapP50N0IUOIeUGWfpbccVNkAmFBWg2/zMu+twGA4pDhBl8n3Rr4CHrR
xEzNwN58yWTcbf4TLMplmpMPJCtymWBRvIIkS4DdAG0ANxO+qLiHODZidZ8nv7iEvXmCW3TLHmUf
qovzA60okDt/pXb/L7CL1sE8mKqIolkLpJjZXoqq0aWeK+qYJGMMzHxRLFwVGCWL9ktzP5UuyLq7
RfXuu6PrBA5v6+IgGFERy5efNz8Ws37z5V6k/nDcRmsjqYKa0K6JlHE8aYPk36qhySm0V8MHBrJO
uWE3IHZxgSWA7MH77mPAyUXWI8zbF6TNgGk0Vbu4LeY8rEabYAS9Wf5x7oX3At7Ljd5lG+1vBKFs
K5Q0z+KU8M/UExllJxRWa8aGLTqCLSR9C0fGFLaQcQ1ref/vufbGjoGB6zmFib09evBDfjTYUppi
Ag5yJlcyLUxlL10MHHaPCeNGnunXs1H03X8fLTUBWqHCa8ku2a6nrLGXSb2oAz0EKNf3w3kjDwne
wQUCVhAnE60RV3akhnjX0gz4RSK55oJWUyNcEtzLjsXhs3wpqlNjbgBcjnGTZ/kXC7E2qb0h5hQn
XQy2svV7+7TEiBi4k1/ORitgTY1BTm7M06gOYzFiZWq1Qd5UlyYDiUI6/lNpunD8sjnOyCSD2IcA
1QDM3sNY5locHXiisNiBbm1O/HMhXQ5iyvZDH5MgbJV86xoG2sczRY0S+FhCzbK5tLAzl/M7aZBF
gS50yopSR7DCpYyLejsKvz8oRa8d9Tu4BXag6tmMzxhnllofLn37R2bkGnQTYCqFrETCBsWZMknl
szAQZYnPb3LRqj8L93W1nRb43ckiYIX/PcI/2sefgPOmVc32c6I482z4g6uo1FV+YIrvufqkTWPv
YzOw8/KrflHL8A/vmbkSoskP0i7+DC6H5ZeHiXMjh8/Gu6e8fN4mDgzjYD8d5GXd7pPZKIY2AvJG
dPPjnh3ph5zWMsdovCax8TtXhNwz8cJOU8fgsTHz4QcSU4nGurqaK56ulfAayKOJ/sHh9/WT4iq5
XS+8CIxvFRkc/ScGnPdZg8e+A9WNcHkb1nSKrV5OPdR7GRWmdO6qkSex8JoWpq/TnO25eOp5TjLd
/nKB8acS7jCy68MtC+T4ri1KKdg4+h0McfSDtjC+mTyXJDDn2+obvVqXhqprI09u7P+FxpNh6a7F
r4vFCozovfYOapUaY3ccGakpUneqJw6lTtF6ZfOhnqns+XyfQCxxKLkXo7C++wKeqXvxpFCXX7Oz
Y/CskvZnSP+1rDABZqUIXf5w/QBQXH5gxzlmizk8N6dIw5ENkn3zkHLDavaMvFBwmi8Nfb2U2bAU
Lh38hfe9n+BcBzkQXm/TOlAjKwThmUBO28yzK4Ef2yxtHMDckTmdHVOWZQBW3TmXiR1fWV7q9v6S
UV8m6d6cw434u2Ao6ij6PAoS8F6o4tZR3nDWx8sg8afQreIb5/XC6umloEMKI/yzc/hHkxg7vpmo
xKS7gJaZIqsL7mzfbDUgYMEiJIoJ0cz3SeQu26c6OBYATbiqOLqpKARwYg420ttbV/32eZWazP0/
igyU9ovLmlvlcffFNi2MvXKJNQ2jm2G3QE26Zr2KBU+C7tYMeI2gUAbT70W5xv4WMtScuJFNUcj4
Vzn0BVUdPvRln/NsMx3lcVwpupGLDvb4wjhgfqymNliQwfFj3ZoSqLrg+S4prIhbfK/VyPXce1Rp
IP/m/zW7tzaNeOHVYLRMbSQJ+papcWaYweU3Oum/gY3jtepRSQ9IntLnea2rXJ3AGmN3L8wPykdO
B8AYvtSS8lnpjQ7QoOmxf2ad1KfkMnWp9sybXdwZs60U2IrHlzCLDw6RRUnFx/+5cC8UEBl3KrEa
ltkioE72YjErDSuUMzJALLm08Bs6QR6El3wCI9dQxsw6TAHYsN9EQlHx9/E9w+vq40mPcjgMS3bm
9XCtlddDCcwlF4Ud/0t/spk44Y/bheDcPU1cobzbRvfa4Qhw087YkPvYcHq0UFz+UNXuQWD3cEOA
RjQd5lrq3R0R1FZ3FJFarbBf5aQpR1Yc21tIvxNm4XmWjdljy82MbiaqhGzv5vjmkPOv+7UIkkjC
Bh8mShrMUdY20kEJb+o5XVGNnytUqt/GJcnpZFgmwO2RjBRVPxyBc5v531FMCjKWqp8G2Us5JajX
yNjIvg9QHhj6fgEWW4zfLuO7L4GfccVwuzoHvmCL96dR6f+nrcc+EkL/OKtfd7cTEPvUC0P7UdQL
84+vHYvGfJLWNPaDKZiuIgFJjpcuryB/cHqh9HpfSGzX7WRsZqNe9m9Gnviita871guJKj3XrCtb
2e2gsYelMwPqKBBeZKZ5y2YP/kCTA4wJzkUm/dt6izgld8e9Oej8O9V6zGjNfXPD4Vk9SDrPqI9I
/4Yt/03dPTlVAeFHye6paLAm7uMvigMlcCXlnqtQN7MUxwehH/rV7gHX+KA/52HILc6kq/C7/SbO
fpo/6NsEGWMtX2CkVGmPZPGCQBDydDrQJBlfxtLdXu+WtgyosoO8/70GgZP7WySD+afm9aJYiwJD
QUf4hBiXxVTrogBNgPnamR95QP+nDwlxmdhsi8antZi92zOXQdxjfzZMSF2qRcFa/zbhGh7uODKD
pELOovbJaG/jWVXlbxkbcqIZ7qSUjKYC6tJqGB785qQTqlDDxPv0pe/aL4RKtyND75SCjRZGbcEv
I7UkJzlBtcd8w3PGAW+B6YGBezFs1ugMbDGQYdSTE2ZDTLosA8gA9V17QO7CfK5u+4ZSldHZoWuJ
i3CbxkKSuGu6ZOjpAdsnq4IgtfpvCsf7E8Hzz8TaQ89DE07SiWTD0p9jhJCAVjuXy/mVcNsY304E
RRlnCyMFzB4Arf2sHL4tFEhkPBbxaIP+c2mu4v7HxWkKyrZ+LXOMIt+imiE23KV1Urmtab4r9gC9
t+USWv0KSQwI+AiWwBxIrtzojc4p4NOaNHechtiZVBcvRB3W7KsKD8MzttHdrzhpMtZ2SH80EvVx
s5ps6A6dO44GiqjfMuvvNggcHMbbcfkiGBHszXqU2H8LnHrte/CWp3bwwqjnuYzWuoHlP9xX2yle
FKJn91Oqng7V1pvRxCQpCzWzzUIj171m4i3fTvgUdor9BsZOMBXqtqqRfAOnnTCq0PxEg8kE6Q2k
dntvEmNQLEh7ZS9nNfWfVumCv8holCft4htDyBVraKR8ixsKp50+IgT1goSD+o7kOjKB4b8nBXmJ
AK/4cGKJC/3QRtzEdpLPBnv2fOqvxdI4yBX+e9o5l0HymEagaiKa04ApeGCEcBGDFSYIbF9f1lgf
mGph0jlh8B5guzA+X0KYLkT/b4RlifRVs4eyY+b5262UP48MTw1yA7ehIk/1kBiHVNTPnkpOd2Tp
nt4Xlp+n6rwCnAujkALjbYYbYCLMbVGmJUW8pgx6hCTXsT35ArObC1BRT9vBu9IXgzRJx/g6QwVK
kVoDXaUcO7iz0KINlPB4Ld7AJOesCSl5OU9OTGXqn0ax5/aoVScOAfCPJvYlz4OOLQkH349iewG5
45UCNsE+1eawzO1smltLp/4kOreogUEl/Nfq6wvbdV5x7lmc6w+EqUM4sm/Wgnha4uxgRPXQOZ6Z
Ay7EGdiWrO3Klz6N4vwt8lvyipT8ZatvR3+4TNoEe5BM8jpn18SzT4Y42iezFrEl1c/7n+cUu74j
FTpzYbbO5FyOlw4oe9Cmt99DSNbZtG9eCbLsZAUPzCZYnirtWwv34E0rD+RMD5w0cxEVKyiLKSja
Friq01ENCFIHBn0YFME67hxQfvphYSACHDmGi46phoyzUdTg7da0hpE4wr7JiEFtDYnqsRoQ4XwY
EvtJHjYqMju/FUMxgoQQ3U88axXjZPqSe7JO++1AlZeyiKqo/aozsMd8gGDDuFF1vVLb0J2hrW4n
zFAgMRZWsmN+UO8pLHE041dMe9mAgUrj9/2EI7X2BYXRZ2tHjBVHi3fZriABr/zYvfIGw8/W/7Wj
ZzcY0V7EhH9slLpcny4mCGDBwg7o0rjcgLyX/fc+h6tjgaTUicviHowgO4YAbGyuiG/KSo/LhFqB
sRACbRZ7LItWnOUJC25uDGZOLZl5Dpj283L3PFCLUXDC9JzSoAbHxQowGiIokWAr4sQhjKyWGSQL
8bHqD/lzHLAY9GUx2eoWPEhHcVupcE6DV0SXklbswXCnKhrRfW31qeLNmJQXwoS+lsd2mpHQzOwy
Xxz1/83aPWO6jIRiC+f9R5FrL85EqYpMOerF0YFIFF8z5TOcyGxuR6c57cHGJrNyT/jI2L7EsTEn
wPZu22nfjKQ7o4olxDaIUws84Xb4Dm0wUCmMV/PBrvrJNtBtT7FxSrNHLtp73jggd+oGeJ756hlr
cVN+yB8AfttrjAHeBHoXk+Y1Ad/3OGA33pqNWrqMh94joCZjgyZa+V+TctWYQkLZ+mxxg4jXbLy8
khEil3UxbQHi+2oRHwkPEmFPV5DcZEHR0R0wLi1H3nsjYeRcbszpKRDESKjBDT5dcRfiu+DYaCRE
nCGsdxUYSi3Pw/+/5R6HFj3O3QY8PCjwn/lpXS02mgo4us3YKpUu/SAEyjcK8XCkH5bZtM9NJV0E
igGCddeqZV6Hb1ZhED4rjEgno4JOiAdtAUw4hhHp3zX3Q88gq1daJQROXJ6pAMjNCePSgRy6NDSk
cVHKdNNRDWOSGLzHW3m5mqr81vMyFuxQAackZ58MLfME17NU+Ji+NPHYtUWC7jc2bsIPlzCL2DKw
O28g/7zS7hhgSmgguWEfWvM1gtQFHDMEwVrF62+9eTvIXBA5pNrlA68ICPANVmUhkbpIHfoof3Ea
fDUF5Hi9zxBHoDwf+/v+d1bPlWMEfV+ciAqQW5GpFqlYDCn1n/qmL0y0zJBs44ZJtloENZuGCRVZ
BZupt7501lGOrw9iaiFyQaEKOqzobNoXlRTpu64GX+G+GNuj14tYr68yB2cYJN5+FzCKJcbLmBGS
CtLlcZ1wsqHwxaLH/ze1jV5yop8hEzpYlF+2FKEgV8KDRxZW8BFUVrbut8U1r5EjJf+PKrdzsFtJ
NspsnxWhS3HW5Ew/TbBDRWX2Sh/70JvFLBpgN53qU+a0wZ0TVIMC711YmdUh2MY3qwgO23pK4YuJ
4jaL9uD/HzBfKyZ1tjwjtEYPA7BcSPH05r22GLACkFqAwkHRBb13vGKufKasYxwkaGrBuQfGELbT
iSvEYFv/1dT3H+fZk8I56h+oEyaVe8mNkX99SZNHpAnL7IbQLQB3nrQn6FYKVfzf1QhyVAXnY506
DhxSG7VQWE6vkYWkoAX2FUxveVOuoR3QOYwSG5x31l6g1A5pwSFKPRV9b0rTXSMVz6Kok3TD47K2
5HCMBYOV2JdG8PJWv1mB/pXW1G0UU1FjoTrqtG6Vqw34JkMWNanV/gizg61RqcLwdFtOjZ0868Sh
aDEaAEBSgC7vfCNKx6WVnVJE5fifbRZ9fy9jTqum3Y2l5lkJc5uTe1r+VrQzgOkwyahE8yRAG9Qc
cvX1vba7HXAyPWna2Df2ZNDXWYOa0zHJCwVv+czRjb1aS4NIZrEA/0Q3j8NVBP5QrxKKVYW12f5M
TipqhG7qudyhqEplVAJs/reRT1aN/BhW+WEfSKZ9gnERpJ6Ukd5Baq43uOJ1Iu7EO9sbwTtHp3Cs
z8XFA78pJg5+vR17oMbBtKMlv00B9DFg/53869ixe6yWMtiIyUIWY30zw1rbi7XMbbYtANSXmMTs
TcFOkNxkGRHKL7JCCMVmyl1q2xslWoM3TlL/PiV7ciVhKHkVBFjqyp6MLI3cF56QgCbuQ0u3rlnZ
OHTDTXJY0BBa3ReZUrYEtT+NXB0tW4+CvbDl/M5Vn/Iy5Xe+A1nm2JtQNGqNewJCgshJMpMq5SEp
GEem6SXW9aG1+QYvq8yd2xuFJyJKvniyUBWT9g76dGeO371QWUX8L+SYVDTAud0b9KRSPVPMY5Qc
cg2FX0zo8uUCXdVKXjxb7pQ5LdDgSImaFmppH2iS0rhLrsqqqxyMK8WsbdsWKCuqzgFA0vHvNLjn
dDL9sLnO/GB6kK+GXNbBo7C9cOh5BL/rsmMVQviEg66XDyuWduWxqZB3uNpNaQPtifzj/1miQ2/b
VRDB9piDTDLKue4iO9FpLuBCsbceqk027dvKTI31hIp1QjMYdViOsBk8PiKkJlvwPxrTFKNKUbnS
hjbCE0fAaK9DIlyBiaAP6ACqJkLqzRPeWk834DThozSUGAgvAvuZBxvgFYMM2O0DlZeTlNrfUk4D
MCboe8BDppfIJzq0GceAg/M6Y/TAzcx33qlZuce4AuFjwgXAMrYbIbIgItTFRAs4MAQi7CZ7VrbG
cBKuZ5G7jBrUMWBzej08/hkT2ptxPLala4yCnBJ89Zg0aFVjNFFHZ5Lfcxf47eCupDrkPYvKN6qn
VfvXHGY76Svc2Fy8hPO9R/YBX1CKgaFizSaWY1JSR0qy9BZF1QwGESlvvm30Jq9l6I9blJsKS2lB
KCxH2DEwULf3HS2Ruu2Sa6QfVP5lDgZsFyfasPMAJadmhD4F4l40DsJ3uEkSrZAHD5TjLzVJw60r
2vManz915cMSJOZIE+x0swHgMJmqb7IEJyU804VqjTWHunqS7zOP5BGKOZQVulnbgqvfzYF+MbTs
LHr1xKuy1hjw5C6atl4aAr84nh/wHw8QP+26WbXQ0D+etlJEZmeFHdGJkZpxexjl8dGoTFrzbxGZ
f5V9URJjvW8Nz/jOsqMfw9S6UNeTfdEzNOkW5IPxaw8Njn9mIBBAi9yJsqnOIAMgUOAjvcJR90c9
sT8bwmKVwLCQHSjygwG5f3PVfKjN8EVQgYfVka8iPmodVWvKv7tx/T06OUElaVxmJS37vKu/2bKA
3En/bs9gZ3JTfs90WZ2mm8riFePqHrn8Wt6xEqVfx5nxal2UQyyJrdCa24AJBEkAguBrL9ylbuXo
GxgCfmwbiwI9XcEw/KuSab3BqWa0DzXrBSqJ819XtsJZdDNURBED2/XZDP3PY74VpsIGlLsl8uM7
xP1jBUe60RWDkooAFhFMjO63QFro0WoVYIavBd2VOMDXxq88SFud7sue7cVgQrExI0+2oWNwRrYc
uGNRzxcf5do9eFEMuofR377fIwWwLaigCm0mcRvQB2/1URCu3nw9RyslzMnudLORLMHYqA4gquGh
RcKirE8gmRWiEJFTo/Vp/7Kj9vLlFPLDK6/4wHg7V+orXUc364OYZ+txH4MVgTQ+ZEqABnjwFgWM
UlSzJcXoe9DbsXmkvN1YYv3Ku0Artv4bhtGaTKLxQAwBlJtaptjRqL65kBk4ioC1ePTrGtguXX/2
2FJlN0pgeeEy1A0z+1RnQxr+gBxWsWny1AZyjULTfsEcHJ8eUVbruKQtg8w0xz1jsY1Qf0xq8rIx
WBfCKAgiC4EtzdDjTKPiq184R+rmnOAPZ/WyrIhF/cWEwlZcanCz1zAd2N8LXFexCbyGXJXfMAVR
Tz0NnH1C/9plANeU6WXS8Is8D47KYrh5Pbi87szGbr5e3MbTL3sh09ifb/RDc7iXkpzCjOTS5ECs
FTx4a59gLNpVdENOeR4kvyo7qeDbFnhTL5RUDjU4+1EhD9r8bOo/+z4RLnsTBA+bKZ5Q0WA7MHm6
l+m8OW7WWO2BFKRhqgsntqZgCYvcuM5vUAYGQBXhqbRr3/Im4t+rbrL5eO9yQ68KR6pgGHLYnZgg
PZos1RPteVgkp0GpoBS7Wn5ywF4v/4DMnqE0rr9cP730n7QuYHc19B39Ky09nrlLGJ7xbft0lg8w
y5CNVl5CKg4mXZHkTmDv6zkoJrErZEJI+Clu6ix+wI2Q7u9oSuu/CzzSuPG4wp7aexAw7ryzt9X4
3KVdjc0y9iLHLY5HypZ+MlSK4UN+vh0MiuL0qVABk5eTgFVkvpDoQZdYM+0TVIJRoB2WeZxnJOj2
LPNaYiTE7zMHYxaAkBVsOXbx+/5wR4WuuRK3SkZtSgr87ybB7Kq8/jxEF14A0jxcI6903IAR6NTE
XxEhJNqxNn9vpe2m/RHuOKe/ODEuofDfQtgaxwz6cp6mUsm2hYxNAgYKQB5bWeLQjsoEKHpcwqBE
H5ojw6qmoqZjieQaaKgW5IVg0PJX79Nz+6PZHzjlchh+vfrABfZaiGfFMX5zkuFZHTKETmHuKb8L
yTIfZ8w94XgroX/oVmqkZElzJd1F5PKJio7CZliQDaTHsDRYQhTOTLUJP0muXwf+i0+cPwIDZ9GM
lVsnKDu5vFpX6HfSnvABjiw55gNnbJNSmd4CRPMBYStB0qc04spd4nWZnVUfnYOgrr6INUwJFH4O
rlXZU70vtAQkyDy3N2F1Tm5QAubPWfpIQSpKwy6d+X/rTEVByXCAHB9Rob/Gt927Un4rnaPXE39I
ZdMOuAd3ABDhH0F40AcJafanGt9O+sk/aTtkHayDsWMxHjxZD/WMKx2ZFVHC7s3JFL8KOLVG6T6s
UKlxAwD9VKj/huwwJCTyvPihk5oLE+zsuXqxfCEQrTCbQOH3Ysr97x4ICf062Tc9aMxuieEQIC0f
X3rV+RsOyGGetU8l2kqPDmfedLwAD6+04VwpitKJFCgW9duupWa8ppIxFMcTkARjrtoOGdHp/ftZ
KOIRdn1OjfS/N6PNPk49WkfUObYPWO1WdGD/V/MJqD/x+ueFSV1l+aqkHMQEf7xHbHy8hCFWsKyP
0Fb5/U3uRWXx/Nmspa846yslqz9g9csKo9zC0UY4t/6XzHgEUsyGYdtkLUkEpstshnTbf3+m6X3k
ih+JDjHhb/40jSL8XBquuLX1C3rhNjwstEOQrnMMWXTQnjKlY22sqtGzLhr3Q6+bB0Q2us7GgAkT
+8ihEerBHUoE/6aAPTtWpPrfPYOs4Xbbxsh9IilN3KGg8suVlA6bDVy91gAmp2hPMi8XXmzekpUh
6cgsE2s7WowU90rqtBqkHXJ0pgY4AuDLLy4I3xhe4X/zsdnB56T2fm/IJiHeyZF3zrSyJniJex0n
ZS62ZVIJeLdosRBdN5t3GkEvLrSQiTDKVK6hQe1pGlSxyZNEaZ3L2VN0Cf50TqDUMSKCm5W0DHPf
Vq3qAI1mWLZV9voeswe+osm/d6uKoiPqMfim+kgi8pwk7SG9U6UMTw83tosT7YENTq8f4qkor1w0
TmnK7Wzft8hu18pxYVv1QmSXiuFFseS9kjVVLwes5ZZL0dIA2UCDqSXMTcv9mEJJa40LjGaeimWn
r3Wg5WgFA9bpqfbaK4JviEAf1HNzFzeAhpBwZ1cD9e+KD7a5NJFWdIeH32X8HBgHkVG8RiQUa1VO
Jdhckm/kDJJPf+SKfGt17m8PG0Ptm5sBxyYmWWXJ2YsyDV18/0PERAbrKZb3VQ0H6dnnpgKzJQxf
SwkOPLD3L0Mn48EB3+IgAMgs+sij3LZssVvB/h66TMaXg1RpM6YsarhJ/urusvoLSglumbBsHLON
3G0Nlii/xbZw2ze//7MNK6MG8ka1f3tp7gapYG1OgzZmYmAmSpUaJZKqb5oGk4Heq21kTJw4aRhg
AeeOr6pdVTJ4szM2QHmuopl4/22aPguM5/To1EqySVjBdOcXnWGDIEkKQKY8rWlw9yAUjRhPgMcl
1p715dDV4airdnVg7dsEhhD1GG+qjMYI5Fbf7mlbIXCU4j9v1iWo6Qo9TSb/EQpvHjTxhaaTOkqc
VFoZiXq98kSkCUaMg2PiGSErAf6YVqLTCQFVqeuCKyrpMcojOBHfsw52kmRbIQdqBOf2c+P8nIxb
vOY1KyZQ18+zLUrlL5D/OcpKKElxDHnJ1944ppRDWqU0ninuDiMeSDQgC6VK+KoZDg0xgvTW4OXF
1O0r8jAsfKqWPH+c/aWs0X/8ueRiGzyWgpG7EzBlEI+4/OCGhy1a3l+J9piNCJda+A8Ozv0svouE
J6Snh3hEs914DwXOniTGHZcsW0YGiAm2qeVhYPPPilyCqpOHUEGFTe17HK0J5aJFFrsJNhCP1/Pw
WWKCKg/ryjUwVSwbe2feIAMOHb/+kFiYn6kmBDIKZ8RXT+zN+Cc6PUi/Jrw0Nkzblz7qBwuKrj2T
Ofn5J2M7LEF4C6DVFXq71M+RCCv0jzw49S2qofmC6i6f4J4yADohrQtRrdykF9ebojAiE/IS935A
bBvXl0KVEQeUyC+9nhUxSiFnJiTg0DhM4dgThvfBLcQYH5j4dy/+pLwV0jqFU0cUWkNHsqo377Pn
LRONOQ4WK/Pt4tADz03dK8mJLXxm+4qfMwx4C35x85fB98fGoY/oM119y4/v68y+vpFiUESOHtd2
X73Lkg2e/w628SwaL4j+8U59hFrNBtUISDW29M23VVX6UCOA3I3rALQKjduuAY3OKNMOEWbAK231
fiZtsCud2/9XLO+yWpk+EyNcDgkDyQ6CSutZS7o8lO+PEdR2rogmx0bANl3pSz24uUZlh712M0hx
4tLrbR+xa83O+pIqJKJeUXoA/bxtQopyz0p4POzY7sSd7wjiFnLRMeCSPW2oGRLYHGJZwMKf3gDN
eSQUvq0OT8kmw3EXWzYSM82r9oiOKKZ62rYMlQJjELUL2TuvJcVgrS+mRs/EEzvpR5itYyMdSYB2
g0d7hsbI55mrFCcX8Wj1BWwSpaJYSPLFaY1IEpqsjbyX38eNOjhhtBksDvwch4TQPalpOsKQa7SR
JS+Pr9BFJl2mkzJayb5mYbxtdtg27VcvRwC05Z53Z8fKBtuguOREiU2YpFTQPNmlCJLPnK4eHeGj
2oqJSnCBpgt2hzlV4BfJ3BKwIYe+p26g8Q5kVKSVObKggwDG/OvbZasehVsw+E3QFhYV/5RKMLV2
BdtMih8GcSdcQ86FUQDFi3ejlD5WJNl9koX6Da4PZ9Y6/T2zKgIaAfU9o66YAcZHuR0Ph9x03Rr4
x+V0Jfc24h4OFWjM5mtMla7m7QgtraH5Lx2Yjd06u0axOb38jhDWBROGvEE2WDVPyzdESoPHTwAX
RYhBTV7F6VaSmoGwAIgLQp7do87M8E6vzZQsazo3aWnQx203xpqqDOCipfxRSGndhhPIdNDZRz1o
pAG0LqvmPELM392pOgP0p/j3VrD0wMws1bEVYqVp1l0qXT2ECySuKalBnK8h4IoSM0Tkm/vhaDNU
A4FygOEUI/Wc5xuXQ4F8EzjTfLCveP3TemkJwn4jEX4e5tOb6R9uhe1hbqbBEs23mf4DeQWpfiPA
E64RCXXggsNc64fAb0hKEHlbCJhKGzhDF4yaN4Pk1986+A6w/KbFl7T4HNI7ehO9av9zVsINIvg+
1+bWO2uu2GvK6hJJh6JbZfVD2HDKWWYzyLsed3bQW0KGqiqymoNjs6Y2xwLAN07d1moz14CIA3XR
iR1APGKpRsUQu8e15OWomc/6XuQL4i6eDvsFJowYk7EOQzA6IszIQZbl5inGNfJQnMR6ExJ9n+OP
yhM7NF08MlSviBmz5rUs+Fm1w2CvGX6QmB8veaGDtG+l9ICSZJmasnoHmm9XG5nx9ub5266Z3d7o
RBlAjvUusYxGATi3DH+yHWInIaWZE5GmgL6ywReRwzXkIqU6C74qW0P21qRoL6DHA5DiQ+WxNIvv
lsXDiDPHRtWNL9t0NFhdg3FBpRukUlzaNlKf5gpw3+OtURs/GTE46G2bnTb7MY7oDHUl2LseJuAz
JoYFbrnKmLgKxY4ZhAQeDqGyWFcT804fFDKcqD0NZhrxNf77B/egDgB9c347Uf8ASWiTgzNoCByk
1UtpQ/LB1yzD05iO4o0rWztpOkwqhGpxBjmSFntDYR/9zw3Y+H/o/ZRFzdJXgzp3is+ame99ZcpB
/YuHlSfsX/SKFtMOatWjwc2cAjvfBNf5CBn2mCKGrcwwnBGTMuxdwv6OMf7tZ3iAFb6r9uVk60N2
IeBBVEp/Hfq4AfFefwH++MLgoKhQip4qrr0nVjgjPnV+Ayx/efrtWcY9I5ZvhJMmP1CxxVJb8TZO
6GHplvPD5qt94MfjTZjSLa/OLPQu+E3eIl8wzFd6+g1CKAYzvreMSFdCtciQAvgm/3ER1HisjsOk
g1vVotNrsPLfigODpFTakMjnNSkGNaBPSV5yBiAjZCVSaQoeWHdfMtO34l0EfsU8k9fBToRn1Vic
GMvxh0DSs3Ed3BYHJbXxBlIJFzYfhG+G7MTnJ5q3ROjhCJD7IB2LGbEdDVyGDM402Rj9E2sq7O6q
2kf8PYapY/s9lz2MGKK5YiyP3Mo7rNFw84o0HfFJ9id7516v53BciBNsPnqSke+SmnlXdHYlLqt5
B9C/BMMBsa/yiN9q9zowSYDUm7Mtg23zfcfKhX0M4nHqab0GwqL9chVNRXapN3G6BIvo8YFZ3jbs
cKh2vUJ/9ZWcQ+xmm5owrT1mFEEqE1gAygn//58c2cMexXgxuwas1DcWjHkrAFDCmhu9yJ+9/5MC
a9vMiM0hIZ5qYQP+IoyBYdWYOKDGSTUt0a9jLWw5tMnDgPKzrR6XLNPZfPFsydv2Jhn1gTr1+kS9
bUjrmzD0tYePsbJDuY9EcIKx9sozF+nVYSMfq0iQ/uyoZIouS5kuNI0k9QpS/rNF4X1QUYYh9lWl
E/tzxQaCv/M8ZvI+rDnSq0qjOlzs3x+0fXbHdrbuPAcHrNynpece4CCtRte5PNMIywCdRTN7bEOo
Zc1/PhTcqIgbf3e2b8ixGpp6eAHQoCmyHRrWxToQOpenhxTNN6nugTGqxqiGWOFNqwAaG2Z4VmFO
2BHCj+t5oHPnTJqeiYfKKcnbrC/zN7OWGW258skOKzSrNBfB/PoHaaSGP7mPOUnnaWRdk+9SPK/4
o9bbcKsxIfq4p2FTtck6WJjj0XHfboeesdZJYXpwI/Rb5zZ5OZLBOorXSYWFpkshfDiDter42mqU
st3XW9rPHrZRlK8B/jEct/8e2SgdGTMKe3v2F+8mdDug61LsEsotKXDM90ScbGRbehoU5i4H7RWN
KZpdfBGI65pjFZOwYBylXRLn6B5RRDLKhoGaAjSNPA3i9GeiZkycg7XIKUzvqXkvpTaCfjMAgwtp
OwYOjD+sXarWgT+XIX5yGAIi1MU1KzmBhju7fnC7O5f2ZjzZcqH84w/Rzta956BXxbv8Qh8Kwm1O
H8Kg1FeSrs2MGRsjasKNGzSQvCKiDOOyS2x4bxfOhDp7NwXTSkS01ffa0YFKBvKulcwLkST7E1Ei
VHnl91Yko/e4dBm9WvJ+TZg/qHnLG13+tfKwPrVQs82WEc6FceXj1sYbLIBEGcLmMYHvE9viB8tS
uTHVRJMl8j9u2Q/JMf8Z6/svRT0Xd1ayk7Xse7rC8FtOHaLP2V6xM/abQvt2LnUOPLBitE0DxHAn
T3kGGc/sfJUmZP38WAXWifiK4YTpzoN4d3JAig8nEqD6Tig5eGaeUnj1k7OzHtsCJ/A039wpcyVW
ji3DdMMhP87itOfQrwhriVrFn5v1nPe2fjuRrss/ohFOCzYAv95PVO4gKG2QV38ODDQZp6IFM7Xy
2YvOJIHWqJebueHVz8frd6b/C9iZ09Wz/6Br2MEIw+pyDzW8078n6xLYrUgDM6la7tc4xhNX6lqf
KRqPmpxgApQdOW+7rrVc4nV8qmORn5YZXiXO7EFhJj592KM0Oor8BJciTksAAZzDJ7ycJXVwjwGI
D/jy20Zvf7cbTNRG4Qxs07a/quZyCrco1fH7b2jOmb94qj7sZNxAwYrOSyFYloBe1ESuEY8u5cjt
QOjxBE91uw/ysM31ynHQcUSDXQUZGcUJGncO1TWVnr1SNrwbw1z4HqOy9PeDfXEw0Ws/jqtGHFay
Spahq4AxobYpS/nInhdL8mSSc38PczbPpixr+8DiWQyIeLKTbqcaoYXZTHRO2T+Jk7U/eNE6m+7k
djZoThAaomlbB702M/9YKWCkvYL/bYeT1Uml+lhr10SZfDTnnPufa/y0v2+Ecafhg5kDt6jpdTIT
mDY6fnGaSTFevtVwYJvtNeyMLC23+t20ilOFgAEPR2dllNejDtG8aUSrEa0UNFbn9v8gZAU1Xf2v
3BziA1XvEfEU6E16W1qj6ZijmBEtu+zTTlPiYV61k/PW8O7EqyHhUfdnmflw9dbqQcC0AnFMB7JG
LPlKNFymggQObhUzvT1PQ/fiDVMluoQDIpz/e36lBHXxgmn+67SMK8o6Zo4PFlg0ur58998dnxgy
P/jIiKv/CwJm+v9URa70HLAIneaKU4Uv32mpdpr1TR+mwlonhjviC+uwHiupstnCmRmzxhKe+TGO
8gULapQixz+As1hJGtpr2tRVWC0D4LN1MOzegeCIOBj6Wl0d7ZxHZLSLknCM+jw624xNi3F8Arn/
QcP6knfJMs2Yx/A6XjrcrODdUZllieKb/tNT6yNjcGdqnqNnSuVmcZKnj/5w7tyA/0VEDsFclC6Y
2s9vFpA9xXM1GodH0ayFbo/B4Bx7sbehVGvNeLO8xmYMv93PsUAbHfkgeBdvOtlaJSVA2asATfZ4
bdBQz2B/k6KJmK0K1IzQ6FovHQdpyezSec9CeMH+zIKETi07/EuenMr+XMw70BTwuxnnUMLUUJya
ofKIjfY39l5yDbrjgk+1bDVg2UOBsCtx6oqoBkLi0spe2NfA4xoFq72fL7gJLdDmc/09bYaJ6aP6
EC+AhNVfTsNnV0tmaaTitnFMGFy511GVnw6H9dUmwL0PT1AlPe5gcaqaoWfHUdi6gwUvFSmmiBIk
dp/DegvEv5ELc+3FRfAVo5HZafjEhDXMO8bbCZibUSMslLl9ua7jMafZU8UlfIMTNgi/uo/5zhnV
+DbApKDUSvYI5Sp0w2m79y8QbwFVLmFVxaphBQcvL48nOL6HO4fKoKe4rw9zmNB3AgA59BMir8nS
jKBsQ6OtnF2QidmIhgiOVnLTJ71/I7DEduRxkH9xw/dg6fGSwvost5EpPOzwdrt4+hJA+VH1iZbz
gLSmKm7/khNhCO8e4pvxjYRMpUmYfzJu0oX+dWCSQGdZh58zomYXjE3bwGDk0tvQL54UjDZfIy1z
TyYdR8WMMwoe+w64MFQTt9PmGEN5KIuNWawxnsREGzi+KvFiYdv/s8OXLDs4pxCQuzYtchybgBxK
Z21J2VHqOARUoBj7irWbph4lhYNBZer9BZb54xgO8sDFF1cfvI03bOnZfdJdcfepW72E6BnSc3/T
iw6gBMTyhAIGH/ZnJtcwjVghRoxKsppYcdS8vEc1o0Zscn1Y/qlwc/DFpyd4XpqmF0+nFE7ki9KA
uY5R57gRlpkho6OJ1tj/VDXGMyMFuMQezhCH/cr0+ClQnSiYDfH+cE/IkPIaI/9/AS+dKxVHn9oc
QQVcMTI2LbFIZoN7kAHF5/ZbFa7OtlEv74kiOh54loVKn0fK58ciQCHh+v6WWwalhTLYv4WL9UKy
c4mEwoIYnbQiru0iDYD2qbX7oPbxAcqx/V7+wR078dQcgMIoc3QtTfsDUA6LAWFpOiV8adnMi/ei
6mkFZbPIVVtX+oZrPw5XaPIkBx/cH3cOTwYGAICnXQe9tG9sA3+0MQ5RoHSyqEIqD6RtW7eVfoJl
O9XvifI33QY+b0kuCjjh/N+7CYTmkAVL3LqoX2+XBp+36EpyRTQk24m068nMGkvI6EcN1lKPFbYO
UlcbEozjghZSk9RkND/8BcyeAZL4WdFkvDdU6Qxrlwz5ZXIHFxLHrQmQhYgIPWbUMClUW4FwDili
lxaY76QvZUcxgM2xPNnP0J7ObJ8CMGgk0nKluShoo3eKb0If42NlJ88nrO7BLjIlCDLYxTz+8+rh
eUWEmaklm2WYgrFI3iQWrBwRgolka8GPzBEVGlK3eXYWFUzTJRMGL9lFWcWzSMJva0epew+MkoLY
PLHn3cu1ghV6U/ciS+cQAp6jMJjH2Sy9C2GcNgsYMhxLa4o8e84hpsncYCyY151tpCX3rHNWeJzo
aAAxH6VzUpElfjPdR8uCJn9Iq/jKujQ7POHle44v64TfXNcTPf90bW7pEo8TrL5maEYuhBn5t0Aj
Pm8SSMZoTJsahFvx5hE71k9m8KyU8wrbIJx3kyz/NLZ+rgJkpzyI0s79N3LfbQOvdKW5rTE8/7eF
UZ+KrTToWfxgNTMt6PCKqieJ0ngZL0YOYdRUAUvKplUVFvF9q/xxNJ0Zz7aywg4zBRD2wkm3HrP0
NgG17b9753oUXyjhXlZ8g9P76bxQNUj1UZpINYOykLVZi0u1Yv2/bIkI/w4S2xCWopbzxyqLX4Pn
Uy98S+yii6GNd8etyTRkG7RrhQbE/BJ1UhT62WpGXg0phvS+VmxDIbzwFfLI6qgx/ZLJX3fTNfM2
FjP0m1AbzMkZYBDvAxKA4FzuJdA80/I3vDSc+xwpUHS4QqiDU6G2KjFJPmyM1tdorC9BmaxYd80f
Q2uHXq6daF94zjhcGHnHrm1SQOuyfx8TMwoJUXEv0RzGwohwjQ6RNwPsIhcQ3ItKvCLkkW+rFcIz
XKMP6z8578cG8Dgm5MTtsJoT6qc8My78FchuK3F+j677N37xa0y27ZFVI/8KrRDLIFVuzZ20g1/J
tLjc11MTzDEYTxF9tV4bhDBzu7lquND/Zxa2CwzdGeYXkusK4ZgDB7ebhE5FUkw+oInwOO48vRM6
Ruu5QB9Z7BuvvZyNaPbJOFuwysVtcroe0H/rdA9TQbY7F4dMKXPjjrRA4OGQ5rPX0oFvts1N9QN0
uPOFmwTyJkWTjqeODfHMJEAlje05UYGz1i77uXdngaZRvQABTZ58jUzsTO8w3OsV5FqvP05EQqpc
2PelBstwmwmzq4uNBBRzQxN7tSmbg17HInAeEhDhlgLaQtxXc4YwIVa14s3PIoZTpGM5QkGwM+JN
s4DKgNC6O1QDjG6+suiVAOhdu9gIBC+9WjfkKrNhL83r/F/VOT23nMYB+5AykAL4DB0B+i9k6Qnz
fP89Ci7gKvZ8AILBG9GwHxfdK3oKu+fc+JGCRcix9e7yC1diLvZIwUvD9AhqjXOP4My9w2J9RMhq
91b3ss3/rKk2Q4pfDyDLZWHg97SV7LwSiAwEIerDcCRFlkM5I5a25lxTr7LWeGAVtZG/sPxyZMS9
o52LoRoyvp/7I3QDVDmgGnspjg6huXPb2FFy8+qwFt/uWs+n+TyB07D3dNil8DbvqCACWQ0EgqXW
m0/GBRL1X6rUAGRtPKRt1AeoCwGooqyZNlk1sak4foRLrEQu5UVC/lK4SDLYiAS91VSQ7Ovx1t6x
ulUzOG4KHh5NYndCth7EZWQKWNtiLsM3KtqnFm6FuPyS2F4N9GqcryX8uNVgeBLiyC/JHsuYnS2Q
i2oxO7CDbLJMbMmAlCUvoxEpDgWDrjmyTUNyMd/QgnDYnflaB1wNvAMIbhvwMBXHLQfqBNKrN2q8
L2gkND8RTv78f5MEizpKxx0v6CiAHfQnspa7kx3D5xqmrlObXYT0ELANpB/r4aI7RWjEPS6T6TKe
XQD8mw2AiigdpmlYb8AhQONFnVgsbPinF2FrB7KoIYnoPbQl1mgqavgMeehQY99DsLxSDv5zRXAp
RHWFK8u6NNmsBNPE18HO+ip7Ufk9cdZd/Ks9FQxdiznzHYqZXDxhorhaAE/jIEnz4CJz8co1PgMF
TFApOoQ2HrTSHRpSRTLf4v/BZVk+jMUmYqxSCKMfnmQ8gl+n9bTF6I6++VU76t46LhMOBRJ+YamU
gCV47VUcOR1xLqb4h0VI83yuS7oF21Z9+TkVc/F5YSSdydf2nwUjuQqQusWAUuBEPvyzAMttxpO7
KE/JkX7NVTpDu36r3Ka2KJSpHBdW2DzYDfrB7j7qgNyJP+sHVJVY5wAdZGqY8A7wFOeZRn9XChbV
b3EugqT5MYdNWYFLoDYtJiMfx5Spvel+NSn8F5XAISCbbK78bRJ8kbOaQf3ccAqls0hdqrF02w5z
gi/TdziJNpuHo0K/5Nvtl4vktu+U1oC8M7lrmcsWDg/allZix5EYV2ZfEpl9Um2uOA0nzUO1qZHr
x86QWnC43vPP8PhFL2nCI+T3vTPg9nbeIqh6eo9ZOzv5rDFU2lbnppp4xol8/3CESgPJUdVSbDb2
ZBjbL+IJUHIhG6fa72gII5xJg7n8RkkUQkMRyu7Vie0PIJ3GI6t8Npa55kKBea0Mm+aysrpzOnHi
Uq7v4WSFevd63IDyEaCmWwHJ6ZFn+zpzZbijzVUVhZkH7x5lmpFPTXVZaD3sG1KMI5ElsNFFShwH
e7U5+jScuwWnJ5yDh6ZcQwlC0Jr3nqYNZPw5eySlyTRX9KCbQX5lBidCOlbgtTaHuxCmAe8SPlIA
0XxQ1JYpcJJ7e9roTBYRAdMpjMcr2JWBa1ZUqgHgSHs5HQrgrORHM1C9UVH25oHM4X4J7xYu1NUL
tGyOweYYLKzRe/g2szYPWPfn1iEaNmSjuwteDUPenVePN0RtA0KJJnBcIg1bhkovq9IYNwLy3YR3
SuW1lCNMUdmtAmk8a0rPetDMTIkMUOe25aaqFmsJAu0KWloRQqu7SCEmQLmCN0V6lGkmYgOr1ahl
PKBSoxQQbbYve68oLDB+8GGvayxE4D/ICG+Xv75NIvMkNgrOPxj6HS3iGGAeAQWPDsEtB0o5y6Xy
9XNIoFdPRhZEUJaRiUiZFd17DoGNq5ZpKXuHEuPz8BGO1kja/pb4fk0jYZzIJRixTm4+f+R6V0C5
YouJVUx4hsgl90oO98ZPeAbZn4+TLsA3oXdn+nTez8WzqKmxkvXp2bz3rqXpemkY958SRSpfyO4i
ckOuyLTNc2fuJIxCzUszqIwdkVZYlIkrDDJM0XYnkkPu9pci80G0dIk/QQlyDKml4JIWFKCGEonU
b5XiHmWvOzjjIbzMINOY/ZpFFOGBDPv8NC4Edbj0T5P1SGAV+r85LavD3cSy9Q0uwDBYug3tLkFO
3X+LKdZDZNOyMWwkwlcpqMtCbHNFmYpiS2kf7mfKUrs9MezNcRzBLZxwNDdXTRNsRb2za+5+Ad3k
oDRdvqd9UC1PFYcakyg026v8ewKaAVG4JbIS8tm+gCgVCi4aBvQIJCCtYzK5tnvSblJkrpCw0ofp
dtbeNw1t1/fmUTfSLaOOiqqeCmmtnZJnRlEQ8O9O8v8u2TM8po2vkXXF9vnNsVBCR9QdbCNVR8cx
9hKqefKfdf4+ORbc/ytRymgvstt7ebuBtCPsxoW3Doxfv6gThXwbKSWxmEmUtsQkGlO4HpxF6d7e
nNJ52VBYHovS7QUS8HBJFTsNaul1oNSC6hbuXl3nyW6BVTAoOEbs4Bnrm66+4tbj5RmUtGoGh7oq
RpFhe5MT4xTuTOvYf5uoxb2mnJtSDj7iF7k+PgEKViCAXgdUPBgUk3V3x6GhMQsDkiSlrnMmiwfW
XuocG3bPb+Ye/GN+nBbkgzYn95xFy8BDeJ44oUhrRcW3zfmaFpAHcEazir5midvCw2uqxGaizqU/
ADsDtkhI3ZYVDNZxNqgWfMP3SA9FRqWnFluSIqPRx1N//3tP04ZOC2fLqm1eBKvuWEx0RICY8wfj
2A7Et+EE6/8lDk9VRMR+GOcAbfK0ptFQxEYv5iONeQ9+rpTfms9H0owUAAMQ0NHZNbhmYVUOVw0y
XB5slhzO2qyBbSYWhg1T4BTQaqxIOxkChfjhbcKM1BSNysqS4Iu3aT2nle1+tjYQdTZ53ZqDCIal
rBzT4Wc3NbZyB+AVRS4a/iq2iEbcKozVu0ZybvAbqtK/xQioperP0wqvnDoBE5UQHAxEt8q72Zdy
WNqHoSqtjUoic+Wwkg7Mw3DJ1X8/eChPpAX1EVwf/6gZQQmFS21Te4dbeKm2T52nnBJxMipVJMNk
QaOywpCduKOmJY+QW/A95RsjT7ieUhW+1ICOtvEk1e+3ZwooYdC2dLNrdZRl5WaWEx6BNeVgRDv/
a5fauipQQqwT47KXP7O4MhLDxXuzZFe51xuyPwgKBrR4utko9lJk3i69pTpKGxUncoJa8FRJI9IF
bRCVZ3QalPK4gYsMaa80UnIKrod3aw4pZZWz5fTocYbvBdwsod8y2VS2X+fdKJjcPGL/YWMs3v61
e+H3DxPC1yJc1NTyyoIUNNtUB0A2uIUtOeKDnQ52Ys9zs+mi/+RPC8Bpc8rz8n8Zq2Lry9MIAFCg
P6mVlTqEil3vduB/v0DVhmSnnvFSBjBpiv4Tfox8T3OOvWA0zC1VWEldU3REbcbCKjBk59x56z+I
isERRqw64Y8yib8tSCI9MuqBTkmT6w9/2uEtD93DLZVQfXDYbvsMu383ld5N3L73xJKlj1jUhKAo
8FVlGOUM63iyjoADYOmac00H8XPwtQdwS1rumXzKWGxw8D3jdl5dQS/jZwFhRde6fejC+AevUAED
W0YTBUySPIXXZLcdETRqtQ9MEeXpTloiuGiIGsRWV1Dr9GJeN2nIN14yr2e65rSuwbyWgdkz+6Tw
N0SfEKIqubqZegx6TQ8GQw0MkEhwntI11cnbaV6pP2RHqpPXBZMVHLJDUSfRngiLDKy3tdWd6eJp
UUISZayvHWhTiI7GKTt0yEKUMxGjs7rTwijQZZKYP/gwsECUIzkAXryw7Jtlb2bMCX4aZ8Tq4PJ6
brLm1GDnMqfwCcJMIOUg8VVmR1Mr401J40s5KCF2nvIxXwZZ0VsdUbN38IUl9tKuRDQshwo3N7hb
GbvzGjY/0Knklw2Y9hqtbmehdBoHJQog/PCLk5DQncirRzO7awb59fkNVmzmBvj260kR6i+J2mo0
/mySUzp66nUsKG7PNcl1EtTDIh5vipshipMALXgRMTsaKkUndJMGsO3D2Z6Bn7A1Cu3wLIllfkin
QpY3HNglNcXQ3Fh8a4HcrZ2VUMFarTtSL0SY+ge4WH5A4Xk9tCHrryxV7jZaZleM3vnhKWvJtYQ8
fORiLhYVNINy+uenq8qJW/bNW5mIRlgHCzxDKekEd7RhNreElMpd47hAs0U4R9x4yT3BmcvsQKhn
FrQWovRZDbptwoWvhel5dCbhNjxKlNUrJG9RuNSAJF/ojwiG80WR6P6ujRJ4t6MVmma/DmZTg2PW
5Fteab1mmiVw9Sxg8Bs5+7GrT9If5Yc40mRo7kOvgJGM8O1FIBz/wpL1ZsJa4/ab7eGnQzuNh/p1
xPxBgD+KsFknCwQpgyfn+lz4pRgyBNLaIVOIX2vUwvsFgP996UhdahJxQeaBVl+41NVTTnlOpMCe
a+t1/QReQtY6yuXPrlcRyKtEd60HhrudapWW1Zva8V9wIKkKc0P0OQcISLHinh2LtfVS5NFFr/Th
1pxkH052k+HquSMFk5NrQPrKMBlea0JeAQ+d78jGJ/nbOHZbWOeZwovkBb+FDm9dH6nWbuhqxnnZ
zqoPojGBh+TE7Csu51bRiIRGlcyBPv9q9bckDKfTaX8dacMb0SS46GUUXXxm9KdJhlAovSU633Vi
BLQm4f9PdOSxiCKN7c829H+joOdC2NXrs0DhVBzpxOQkiFZDeDJzFncsAwgCAkOwBLuPUbqPFU/4
h01dEujF+5K1wlzG4QwdULaBcuRyTdzhpHLRltP1vmTYFYkVUJc62zOxmOo8CqQJ7+0soyrjoOPH
s3E+wqr/YVJWDXmhvj5gwNv2HNqo2yIemeJmQhLScbWKaqZ/yGhwhI5RdWL603PQe7HYf+1YgyPg
1isZ1iWasOcGNWHz+iI9qeMoI23jmwcfk5jYTnCSeZLIzjDCI30hW+0PxoVu17lB7gn6qIX3Z9Vm
2gKLTUkhF/vqsdypiFe262Lkp0gDXmgzNfN2jzVDnMZkjwwSTZh5XKU1T5lcrNJKEQJrkKO6yR9A
Q6id1aO8Y68O4VJUsE+0jvQ7C2ZqkvP52ASklpYLUQZGOegkQmdXWfRd4yO6BtCT/rEiLjx2FY4b
lIXBAXrRxdx1jdJbxMjWiekmXY3luHU5IccbCDnUh+eU+gps66tqmWMbT7q+yVG1rNqzSSjXPq9K
2L5O1qDEwhkccDLj2VwBqmk/jhh5WsrI49iGT3aR8C0fdtFLGgzSqpFRuAzkhmuv1k+GQchnOxNE
6kOFG4ZtBs7ELA7q8hv5qd4/xEzUq4e1QyDdmJFrxy+0o5OWO1WpBxzsHAkRQZZBPc7A/PT5C3GJ
izJUXFNPFNCxJQXE9q55LLmm5dzcCoU0KU+3k+KceaHImNwa9VS9a+KFTVVwi+b3RGfAtHifUC4h
uDQU7petSrYf3y1q9mGlweWExnwVldEF+SqPStl/gmZW2a96RYWdA0qdAuF/VgAyiAWbevhllHKL
Nag8gZhSPUsHygVmF+5RBwSVjf1BeOPSHGF3WySH7OHz6VmUOYrev0k2hLqeFX4n+RbaYJPZeDKx
vAfFNtB2mdT6Mq1JrFrbsx53jcpemHHp7jNHXpNd5LvijeLOBqjYFfVa3up9NbFMeABHgv1KogXU
ykL4OdSMxpsSqMq/kAY0gMv1tSYtV3dlvK06fy6qH8MlVrXVbJxguA0c3uX1AZ7ZRaOEDtZqfY1H
sxWc/ffGL5Jlm5BcuEgFhAkv0Dht9FSz1eL7+uwY6OO9g7cbrQAyDyS57iX29w4KqkoVlRVIdSvO
QFlxjLVNJAtf7ZYi7q5WOY/71B5Urc4bQjvQ/ojtF4LSFqF96hLg3DvKj7RDMjOTUMnCN7cE/Llp
Vtq9oYSOhPn351pFeHfNnouYgkcSjxjtCJvC0G7Fu9K2bRVE2FAAXurlTobfXPDCiP0gks24My6u
MAq5lbCv8Ne0WelKy7j5SxHtvvMWsFUbBREYqYPQlWt9vOAamEsAtaNxPkRcARtvUpi28n7yHWS9
f6lhzIb72l1yi2uRtiVJiqiPOWz1M0o2Xcx7I2+6iNo1zwfLDU5VNLCqwzx6N9ninT0N0HAfeWvN
FJHTeo50xmymJqeA+Jj3ceH5xOBAXilPQno6/PxOMxYWb6tZr3uo0ZAYrgy66+wPnkBbvUSGR335
DA8s0NyTQLQGwcxf/O5sAd0Qo5GZ7OANe4rh2seXLTgvR3xx7IIHXIZi5RP/3fMny2ut8pdPbLDw
VeI/7juZ+tdW7IPNdVWv54MMY5WazdAX8+xCs1u+nLY26t9wfFsDpqj7En+kErUNTf7FdCp9yM+0
vBA0JVu2Cqb/UmFJjGzcI2pzkM6CHQGwKoZDaaRe6GrQstsgpZ7ORbTXAGyFWkie+25urhBjhWHu
OposfjGwq6oSMzIJQEahlcBXU0ItNoqslyo3JrMMs2qsGdet90m4cd+5IAINz286r0U5HhITK0uL
9QsSN0VGK/AjA1DHQwZ2/qYGN6337s80bJQAIhvwn0Kjn7H+x3kskbtTzhyXB/5EUBn2i4LcDHpp
LzRfDJnhJwuQD2wbGvVxHc8rFe1QU4YTMOEEfxUxVOdqcQwGxz5nKgJ1VBTnlpQcovE3onomVpqO
KsRfR1cxQnxran6yMADRPcfdtFGfzb1w8eHRoh13IOHJFSyHcSdyCeVzug3lBdpIULRBc9G8d6Lf
t+NgdYalLT44kxpBBF2+IgPHOzRWCqXtCkpUc3csdPcG/B1J7vzMdi+vLGzKzsQGSdp0E1Bv/KdP
KHO4tywzt17GjyU7rtorc1dl9SE++z7eBcmv2fuuHq4NfWS7Dn3nREcLKSfd/cNSvo6qCHbJk3Mm
laaMg6wvCbQTL3vplWk3rO/02jGWpd2LKrNdxLUytr80bzqbX5a+sDhJ0UMgZj5iPI95xsR+153x
TDVEJQ4Kn4mIaL+zWn4eM0DEoZMRJpF70h2Yf0iPtbI2N3m0//M1bFsJ+jt8BWImmlxgomXPgPHy
/7vWfXGvNPt7pAc+0Ic+uErP4isKyljkrXP4Bc1Vi67abx13duzitUMujCidasyA0H7mzX8u3AUD
h0QeiYzL8QK0PdZEKZqGMWsR8xbATrGxICkLRg9TcWdBZzVOXhGb3MZoz5VIdaMfp7BMXPYmIbse
eaUkNnqlX6XVuIJgd6KdofUrsn+UJCixjU9s/Ocei+krdWjoFCLMBtFxJ/Qk33DG2pgNwwY6yq65
QmAxuxpMlxjUJgEH/eA7kHvnmUjJI8q7EtwBjktiTVbuEnq2iPoKS1Bif83uSdh4nIgOpZBvL5qg
cBa39TNDLIRhI3KSzL1lgFVUu72CeAtUE9NlUGhtZewttbfWGKscv0XJiCvWIZOn7YlSV3NFdUUa
DacJndaiSz+IiHTUalEqCOtUz4W1XYo6iWzUKw72t9BEYMUNc8e+f4os/01gMjvUs7o1XZolxqUB
mw7n7d/7LJEADtQo+bHBYdQDVNAVeFbCXbimmhiWVFkOz5plqjRwmN6oTKy3FeOghhBJ608k7r48
Hqn8WRY8hay0pPDkAnGcT+zblSl87r1pu/I4elnFbpJ/Ahmwo1fayAMDz78dMISuRvozKc9UYVG1
oH3Qssh8uKvILBq+GmKuOCdMWD9JRI6UwTKzAJ034ZV3FcuQXoj8q51qGmlNsC/i96KJ41Ywm+0t
ZB9K/aAH//nzUE5AbCHxOyzeT5Rh1DIUlOtIninpqxod355CpVCkG7fC+krFuCTno/b3flYK095l
RtNWmBLheQ+8uvKtwLH68uhZvBLDz5eYTrdHuvGMN3j719nweCAOX4yE40f8SZuKJ3q34tVpTa5f
WMHPkuz6q5bF18SvLhIBAB8EkjzUOFc9VJeVuLX+omMt0Qhdp6FhOoOuY60aueBaTW7mpDRQXqTc
cR86rlfanDdhjPG+3bqGUeidzRMaHVy5hSRa1dR26giLc9/mrzVYGZ+2GW78OhQpkQcrHUGTAd+M
5k0gwHsBEUnZLA+dlaFsxg7+souJo+WBQdzJv1aEWrm1155d811TsfRPc+mKMQQGbFaOGqwK7ZZJ
EChr9j+EG5tln+BzIS8tlTUnpuzEO1PzTk+kdH9JOTexOdn+ZPwGkDNmE/atXEpOiFofb8U5cX2w
bhk962vQx3TJ1X2ui57TgmWv7worfAchx9ygyLCLL6boUN9ifEjkp5C6bQ7AXrIic9LHPdZIHsUi
pkws3fgUEwpeFiKh8ddxxQCa+dRH0n/Pxz+HJVJtUhoHS5Hv5hzMTD6Ew9ACGSp0Fy+BQ/h+nIgJ
iRlGbQe8+oZXYagmcFXlrFD2Q+0S4eDneZRIOeKmbN4G0oRwRdOW9AbTy7bSaUvTrrlRe8ZwvCcx
sFGABGRkFtvi4G5tGeHc/jvk68SIlN219SoVT5EG/Y/QqX48XSG4G41MLcxD2DQdwvDOmFypHFXP
pdq+W0ta0NdKfkqK6n2pC6ootI81mwjGpvv+0sD5PDg4OAHrtcop4HelVlPjQ+oAKQ0TEnNaHvdW
qkw6mw80tKeSpnvL9aZ9nhd4YpT71PUCackMFr9+5PYbVhIMLnqT/hksAAnSt+7IFKBWHANKnRSg
CtPKBNpQ9G/Dzl96YsoQ17e6jConCrLMPZOQpAiivlCrQjaOX3D/t94JQvPTchkZIeUycXtsoKW8
enbBS0p+RW/hbtEq4/rYTO6uOyeb2Ey+zx2XRVrlx8B32tJ8E/ZhP40EgAko6Vz1qGk9ag8ko49F
wS/qoTX2xw5Qpp0nyZuLe2/aD69ZSwYq+W8a3tENHIjhMouHWQmm99dFk9ismlf8hKQyE7Dety0j
VneG1V0wrvUDgB52ynrpohgJ0pBNGhRrMN+4mV7FAOG6o4D4wxIZYJwHUbgakMx+lDtge+x1bv8t
7t4t/AjJ3x70RwkmyH60A7dvuV52iiUsXvz9uvW8eZ8b3hlByAthYyfo1o2owqw+0FNOINQtvqZT
0LNtXP4KcL44JyJ0Ob6BQ036g7PCMm1g3xldaVjC+94ghTtputxKQ9i/ScqpNAdkNydUif24TK7G
WoH7DksfBHNoAUbsqdsx+k1CKcitCH4bOibdSwDHOtLhMwu7i275I0u+i367c7FarGm7Yct3HyaH
OlLjRD0VVn/MOfnY0k0tP0AACV8IsxtK3wSWIrf6HgenimwN3Gqxq0TnE+Aq/kz8YhxzbvBTGGlx
roycdDpZRQUkAhwchozGTeKuKzeKdEvPLo8/eh28+iZYsmzOefa/vpqqTOez99oXWVkvxOMst8FY
vzoMc5+BOhd/wTtKq4XULH4F54zp+ZIVLQyj1InZtvTnw9Wcw18hfeYDMRvYz67wavVKo/3Q2/iQ
MtrY7GDycq+a1oIZaHYS1LQz7wxsLC1gRniTFhiKR2d/74GZsY1GCq6g+jGBFcgL9tj4Is6yGyf1
qjaYHaGMbwYmV/J98GgJTHKCJ6qIPNVATsr0cZ03x0AIfa7+qizoExoJaMBJ6RGnGFhdZ5PlcDkb
wdCpq+JzjuuCGU2ka0ayL/dj5hHPEtSWpb8UuCFY/tGuJ55V9BHnazgdkBdTBPb9N2S9G+CWua2D
X0xC6dSrENBuyGpFqYx4+Z6QWlCzKbEGU6XytjBeTv3sYP51SdnJ8PZQaPlxSoNv1G7bnyBTrSOf
sma1goXf3m74mtzuSRSyYLtUT38MF3PYeWEfXctyyQQuZMmPKBxVMDy7nKGM2v7K3rkrCVoGagoN
/+pIJfh21KNsKA42GTeKxhyP5GQRYp5vURXkfMgW/vTFpbkYZzeb+YbRgK52HtdxmkNSUQp0xRCi
1B/NNw7IrWw18riOv96ltkwIZfWuQJw4QZIK/XI/iRvz3cAIlHJd7oe9qYo/b9hp2CU0QrAz+qcE
Bmc1vxgoIqH7HcMujUJNdUok82NGiT0M4HA6TZ12ZWVX01gJsxa1CaXy0j5yiii0DSAGXomv7JyY
LD30XdQaOah2IHtKYsj8Yuw+KNkgUum0lENqwnfTh5ZGpAezwocl57+pGR+m36EOLSiIzi7O3mrA
Hbn+pXZqI9xj6jKQW6I4tLJyfEoKa6JqNV0rYO8Jhl8l2wZ7C9HFD6eTsPiPD+B8YbH7YsQqe7q6
VkQpKy5s4SDgtmXcIfVz9KwXctDM0vJdJHPh+D7o4APcI4zW6LKa3IV0idwxWMwPdGWnYScC63qu
upl18t0zDzJy6+oVXtABz7s8V8KLU5YipK5GdZmOA6L/3t7weDkm5vNV7sTHgyIM5wCCK5TmPLuQ
cb3OIe1Tez5QxL10VCNCF5VCB5q6Pui94ALUF6am1RRvGJj7SrZS0K+h058Frh7KcWgBrblCGDo6
VkG6f6IH4k2RLamymd+JIkx2zfXcnlEhwGUeFpfg/zn/k50wgQL1h1tqbhsZM+OTZjZ+xDOoPP8s
MmAAbnYUyrjvk6zyfOnnXcX5Bjr8fFi3UfSaSph5qXs/TP4Ed7LVbh46GfQ/l+/yDT9Kt+Idhy5D
IWaPMWmeB/zjmKGzSafeVBGi5msyHC+sTlMgOuo5/Tcxtr6PwUMcI29Il/cAzkvSV9iIP9bAMeRJ
BkGYTASmRDAZS6BRm6/3yPli+VVgLRKsyVYVGoEmdT5MIKlXomMsIstSGdh6EOfBpzcxFARrsIXr
Z5OJ5TcFhtFlVLX71po056N1zVnuSyPZOy0eIXiiATlLfCI6eeN2XJAE2aQfUR6ffMbE5Ec1gCQN
/go7C/WDAHCc68yiNs/v2x4WFjlPV30OHrALtprs++VOn/NgrEVeA1yIgcBd8V5uE4PcbJz8F+/K
PBqIh1lEgiKYDe/PFpm9dyXX+MdOo/yfYOxOkQHSvagooh4PCkqpzdW3WQN5U4QU5HMVZ9RpfR0r
FZ/Z8a/8lOh+By6f082Wv/wSOROL16QJYDH5V7PDheMfjkCMfNC8BkDQk/Ipn7EgR1r1fAxc7q4c
qsz1ypYygL+FaxYHgMTaXbph3YJFfK/ccHxRfhSX+XPa9+IrQ3cWyEsvL05moCE9ZPXkmY8unRMX
1CGKd9K8uZQ5riwt/Q3qQ7EfWmWzILJiKyLJLyIC8PlBa5Dz5zOsz6mDefj9Rsqa4udyYdO7kV0T
aYmfOhKBEdnV8gYbFOEcWAVxXXEmLjC+T4fV2ioKIlx7aGxSehV8OZfM6ebQF3xIMHjVL7cOJQlE
7dNjcp+QVj4df84ZwNQFi4/ggZ/yylKx9ry006hj4mPxYAmP42Q8uYjPHsSj4lEtapWl+UUObnZ6
jIzfvKcLUmGQNRharpdEHIQjB113pstWWblD+5RcM/EnryHAGzvrSfyCxyjZP2kjx3/oBCSK4V8Y
HekJ+sWoKrOiEoaePb4P+7fjdcpSAcYLiz8HPxvi3ymPwqYm/Hmbfr4GUyH+EBCjqcjEHPEh3bse
IRMFo0zECNw1X9cGJQwTiAMo9+MtixElEWwrMQjzfgxX06QRZg6lWkKOEhu4XV8kUt6Tc52mQJdw
HE/gB/Qq8lqVnqIPUyRpJKnQ2o79dXY6gJhCqETxM+wreCFNIPQdbURM2wKiWuxCqUGc3KYRCa4t
WjjD1kXXz5nz1/nBPhpxmXFsUA73EAqL2vujhLR8vlUgs74r2qUcdjrdv4w1s5AV+wu0jYrXPRX5
la0Rj/264hpYEKGORxmItQTQr1QtQfqJbMjXad06WOmvh0TmnqT9Z7Q6MckqfTB+pwp5FJuHT2Q0
J+XvarJI3wcwvAYfBFJDvuWjEgNZUEYgC81e9ROOcGQ47LyUTLZGk2Jbhz2VgPmunzyqXfNeXirI
DucSjtuBsuiOavRwte9zhkYlnfS2g6Fr9v475ypuuBil74ckMqxhO7O09IripDc9/lIQWD76u12r
HsE4/tOhGl/XXBFzduSAqn5YZpFbWyFgWhLWgxASgfodFPYARDXVviE5Qnhyhj3m+BYOX0Vy1CF5
7g63GiIiGOry+HXqRVCNVdma1kY6GYtYThXXsXMyzMckJvjJ6HuMX5H+y/wFFFNGJ85wJc1T6jV0
su+e/U1/rA8j4u5JKqxQTdmGJsfzsNKM27M0viZXwA8q3/EU2xnM1Z03axtBKr+zZrSqMcbK1OnD
0Hv+uyYz16z1drgyUW0LXeEtaQk35K7Mo/WNZTz2VA89dApv3BaRGOxKDmc7dOMl/ouQMMWlz3Zt
cOxFfcQsNArQPc6/qnKHCsaIxBSg43CLjMjObJZZfjOZCTRj2zkc/e8qjZmmaDW0u9AvO+HgyTqD
auS2tispFE7x1NEcrAnPrR2kOFTvza0KtT+05NssHbiF8LCxJ4eBDtxC1rjY6ozVITxZj9luhk5+
h1s+sc2KcG1PE4ShFP3QlTkRi1RrH3BfuqNWN+ImHXBFl3pKO1kMHHKY6NpAT2hk3X2KRNPgLJkS
P75AEGxkir9QprMxdv5Hcke4Oc/DZu65GQqtzo+YijRogCyrOoEg233w9wzTjRW+Q5+SE2PpfqJS
QhBuzWZDa6nKHdB71vMYJwvQtDbrNrrhNiMTamROqXfl7DVidmqUHcOQcAHpWz9J+9LcTicsP2Sb
S+lWoRndMatiIWwA7xBzv1USyQYF2RpInNCDyC7EZezKXjcSA5HT1PacyFiRlbPJ/DNE4E0EIX+2
1yrw3LLPl0VTRhjkEeDNpkD3zFHTyL0VLnC28GeV2scrt4AdaIsxCXMO74FCeeQovfGtxkn0T4YA
aMXxzFQHIhbXzF4kKlL7iE3CL96yj0irY9iY+blu67Mil/K3HDty60jrV34cvbM1T8mx/hHuqHWJ
mdp78A4LCRqKoE02k36U0+qQ2YWvIFbBdVEbu7JWVWVTXlwn2sSlnw1qWiq/EgylL0PvsYFpZhEb
BEFfuvYYB4tp4h31enHtsVGuSVJtSBNkaO8q9i4TYvyu+pVY+ANsSXz4BPW6e/5qF6/mLCkRuRI5
l8WFw/mobEPtN32l+PsR1VIQp7S0DbhAS7fCqdb6T8iKTYi3FlXuEI218GOX87fF0/j3vqCav3Ta
d7K5yk/NttY/58oGtXpDUbejS5c36QiHVpSgIHPrnENcv8Uxyn3nICviSakRsv97hcOqTjRc6RrJ
fAxl2qi0dOMaZb7Vrg9eVWZdakCshhV/oKiNnkHor+Jc+z8bELdpGu8hUg3OyBE+YZAgE0Rrr7qa
SEtG0ONL6Arb08Li2JhsPQG7jXZtCDODLQUfIC6T6+N3LVbsX0uwMTWC6shmDSSQu6NzfBGd68lZ
gj1zCG8MP34tuT+xzOXAXofRV95OeHs1Hlh4sHzHmJs3OL9Y8ptNBxfRffnDgEIkTYDkRMeUFAJP
JRX5G4sjqks10iJ9tAvWrwWgjxHhuOZw2oVp+O4uZ3bujQyMEw9e7JpNwQPJUBSmttuuJ6mjEOSv
M+Xd5rqtJngj0el5fMkN881481M3AcV09GtY49ON9FahKDoMNRN4xInnyF68YY4SShhMW0w3/kNW
2aXV6gUA7A9c+Fdi7lRtPaX2RKrzD+MEhX2vWgTT0/8/CY1bR/3/81OhTU80S3LfpleFWdpPZvdt
sFIfYBlm/mnaTHbW+n5oEK8JKaca8bO8BB3KIVLjC8ELT4/NgukH4WTJLD37feU7RL3H6BhcsOJf
ieft1gtAoCsALUT3uJVfEx6ZwBVAHgC/cFcFd6PeoF0NMpJ3R4Y2Ot0+SyyPNrrynpFntvrryVXk
1lS7mBIaghMOtI9scFg1QLyzScNWli7JIoK/UnOs4hdZuDXhcWjDj0ky1LM0PhG4ZustyJAzb7nv
Q5PK3cH8qEx14HqOfo+wjBN3m1F143T0WgObqAar2i7XWw2+XZf5e4mOIk1muN9TzLtxsVt6fYOd
YDW17BXF5ZehdvxdWp8W3U9K4YL8FtgfsosGV91h7kU+F6XIPaoK10Rj03hMS5qkO9Pj1FDkN6vv
y9hARquG5z6+bYgnFnGUwHxJicCkE+Lnd36JYSIgQ3AmRoU4ttsXGrp3bqOk3XpLUPiE+7gJfjMQ
0BlzcUo9+TH69sYAAE1LqWqzM3G9OqCXU9PVBZVovg/TztP45eIb6yf4MIiCOAziR6h7DWulJWM3
AjnOAnPyDM/p3GpSmhtAYIrINFZm417dpAuRQIgi4ehz/v12qSekNuTDsSe+XXOT15QhAtCTDDzk
FyAcCdLYSHV1+s1vw6Q+VtxRABHIZptKBVh7fk+BmO7QOoZPSYLMb9+ANnBZ/6AALGyqQijSiGKy
jICYjOFw9m6LIMV0+2GsS+C9ABtPX/d82gbXIdMFBcJNwpCVao6rlRpMLn4w3LYvT+JsbWmBRNYs
2rCRpHTGvhESCahyBlpfHSRY7kUrXTYUxnmHNPikyciu6WSAy//emZd4GYpGdLbCDvhK95kONwjo
I3gLFzvSscuKwbhfnQeOTV6NMd9q3Q6RAqOTcQw9EivgV5lNLvHjvwg21/oiqg0otwSwWjyHt1HZ
1dl4xbKdKUiUlx0ahWTZTJu+h1re8tvsPkVAKdnBoup7ofh20N6hw/rx/ynN73XaaLLCAxpot+An
M2tZWDUUeueTkRPv8Iz0Mk349HQtfx06JoP2ZtniomerXxUQK2E4T/+KtGtZjhKnaq6rNLQeVBS8
i724sqXfOcSkK3Ipxxg6EaN3hzrcRyMQkn4jM7dNjnZSay0THI3y30ZbpTHlrgZzXERDKyQizLbw
zgswp0LorQ/0ACXgbO0KXiVPIqRA9glPPSRoBoBGclE1qSmTUWelk1pOh4tntmMiKIwuNToXyg9D
/ICQ4Qpm9nGeoUvrqAIwIqcCzG3UmH4zc5LZHS3KpshpX2SkdXVvUCHUnwZAeNsB0uvOp9HQP/k8
TmGSBGvA/1bOJg1xvPrGGWoi4+AztgDhbjmwFJwp1jA48iKXDrHXHtfIMyBLb8vPZniaMZsPB1LF
1AQnfvzvFW4rSkX4c/IXb+FcYxfo7jq3UGl+SbtEoXEUQGER4mvCY/1B5bgHeDqEp2uCbsxslyuz
hC9HtlN/deG18cvqAhrCcr9bHJKLxb1r4xRXX9IWShVlHtMdWr0t1IsFjqYlSrbzoYPMxYE6ljOV
Ik4vjz6/oj8ecDOaKinApYNxzkN3evw/Hv+wVy5ICnlr1svkxP4m1Mite0397ijSxJzR9xQU8BtE
xyICapXEu7+ianoQQMYej9aDw8XDpEY0PbFAA4mwpWIzZC3zV0pjvWU3xUfKvJgX+1K4Cy6iym/z
LZ8rdaUevwshaGSN4ZFr1bC/d1qL6bIJ29xGLEddRJQfsP86NtMCpm60gmFC4uiQKmM+IPtw0KoB
5jkfwxIGscA0E+6BY/UR+M7wcCkjl2f2vKYcrXS62Smioso++K5prOlA77o/WoHbLWJP64YOHVJF
mZy0oRvUE8KeH6ygU3Oq3sqYY+OIWNbRCAcfwMgfsrkTIRtse9L4aObPaqWYyi56YxnZWNuYT4xE
43AbUkuK+Mk6cU1hRk3KNkqQiAOtymafW9Ck45+JfOj5+MsVSoPXzuYWSgrkT7xtGqV0PL8WjHaR
E+2stlX9QPTh6J2Vf0TcT0WJrXlBxhekZgDmvw9EKFBQHJ5LxqPEfR3FFCLO2tmfzbwP1EXyRkxM
HsZy37HpGec1aBkGtq71JkobyCH2Hb7FAlXRS5k2JoQjZjgXfOCJXGL5ZizzsnI4zS+po5POwrBN
WHyisrNOx/uw0Rk/6SEARtMtfMnn3e+2uQJoh1WAsu9uIM13uDQCNUkZ2nJTD+Ar6KTZx4sruOGF
Bnv0xPKEBE4nU55BVag7/Wou4nA5xKiI1MywTKNFOKWWkYO7/Q0/QX9PegA0k5aAAgkb0AveDgxS
ZQBzcGycdIpEgNG9C8hmgWwIA+f2+7WU12J30LmkuroVuG6IXPP+Lq5uINsGBtPKGJwQCShlzrnI
zNq4FAMJ0GEarb9GAfsOpBKehicuF7dtrYaOURBgy/rebN2DhB8kao7AvaXHlULWng/lLp7Oy5eP
u2Ve5DDFaxPo3P9HRBj6FUoHqSyenU0b5AYV37m2UlYjhpYr5cmWtLJjBmVanmzrlLV0J8ncoMg1
EZ0nRs3xdG3Qa7FPjy45i8dRw4GLYAhxduduEMrbMIVliDiYX8pxaqYL7fLGV7hho8+Ol8FJ0bKq
IJ2WRdaNhA2XJ7JJsmxcKbw88nsWRaYwWv4zhFeqkqwQ7qgpSaPfIrvhr/wr4rSRK80lxI7Vv2kW
aHxYfv7TqO1cNntMXKQLEl6PPB2qp1hLf5k3Ii3QdZw23kzeGoFPsM1wSRXKPH08yqsVgNXfmAhc
sdLt2y86bvqE5Ss35TmZPwP81dcpHpTPySi1+Uu18fDGfMlwVFIOdgcYj679f15DlwHiCpiAgr5K
VK5TQ7T2VMu7qUoAgcZlxQ6Dmyqi5+50tPeOaXWfLNr0axcZ6HAqUNNMX+VnrDpMXXbjkrjMaKjp
oCEYqqoM3yt6BhQSvMHb0AdIuvMuJ9E0SaicZ6ftgtlUVwLaEWp9kKb0OM20jW9NOTCmlrDzWOLr
QGeMS7ZuP5B+qfHXK1Mf3Rpzjdp9WvMssL81Yv80RtInIOQo2AEocIrqCJqkjrI2yGy2Kl+kWU/r
o7nD/PIKZuOPD9Q+z7kut2Jgh527Z6GOYFPGku9Ugb5jMVGQU3tdToMYMEg8fgM1rm+spFCV379u
VexmPAE+8p6366UACwyQl8KfHQkdJND+kNISgxClXlUJ05Yvv+6oNgcTv7IG4hmrCIWji1ozpZsD
dk1qbQ1MZ1No/78FkEoDaBxeb6SoKYsWXUPYr0cDAuLUetE5ai3kQJyJWpyaefwec4D5Q5OS3mct
TdkBClK9q3rQ3Z/LKROBlqB5F7wy770ZBLYA62+GFztb3FOgqXYsL7axDYBTcJSEtFW6+tIouo4h
D0mCtd3BLjoVUcYBJXaud1WTRlswnAo7YCMX/dUrsMZSofIHQ5KdjtKasMG199YZ4bPacUUHN1Ex
G+RYTT1LsmMeNGWI0/RIOw1hyyHA+6+YKlzDzMp8Vl+Zw28c/nqxXpw/gdtNqxdXnn4msounifn8
S7fQLnMwRmQaz3QWM1h65s+sYSgGNwUhVT2NUqEaxV/3a2Q+1/mh2OsiTAHV25eq8tZYhnQjWN3U
h/XPQIBPCLNrGgxTE7C4aoI02yJ3GjFgMFE1zR8UGzU9HMzgZzD88MTqTdEC/mfC/hpnzl5SXbsc
dkQLSdCkf8ZYhEU2dUF/lpJdvxmh7BT2n7TtGStKv5ANjupzwSi6mNt2WVu3/rFicEW9k8UfwO+M
SfuRpTuv45MJdgLjrq80soaNIWDL0REgo11XR7C7cqFBlMFxfvPDg9TG31LqDNRilT+0Bc63d1WH
IxCJx8ew7fa9Pktdz463L80CTza11KvQLQzSFjPq6iBFLNwX+wzsaum4JO0odNwmoSB0i2X9xk3t
0bdg8KMCajUvyFAhsi5F92/q/qqC8P6Q9Wt8WkA1BfD/pXs4k8nMPLUe3/LAi/nCeLtKnxN/M/xz
X+jeb7qS5S2dC5QSrZ8IqEbkKjh/9bdaDtGtPQIj8XSOInXlSguyknNRMZ3GNF+VBzFWwwuIsSUf
yWhJuXEpCGEj9TTqxc8DWy8r9rwgqag8Hr/0yr/nTvTgDLgARCSBZupdKQCa98r3k7+R8j0nFZe9
+rynhP0lyc5WJrgiYJvbMdJT6aACyjKYv6vtkH/2aMnnRIsope+cVMQUEqUJISZVbnixORJbeNn0
fGaqm5zWOVm8oP19wm1omh+V6snKkS6rPkmxEiv3bU4L2AxioACgNvRf/hMssM9Lk90iHVgDXoZP
YcMQ4I06ZuUaQh2QDk/vGIAgZwZQQn6f0L7equiHWo9gGsLmKo7u1aKibFApDYBHfg6/Lt5qrG4N
vlEgPvtgn9bc1by+Tkg0rWTR6AQGTz2bBlpZhp+7x8B3zvX1JkbSxrqxJv5F0lDbByXN8fubQ96g
hWMt3WCgd9sfJSD/eG+vvizXUNAOCWTz4djRdsZAwgJIaZK3ks433y79muCCPkUTF5ebKoi7zYe2
Jq6VIQuMRNibPwjGfxeGXolq9PW622FRLae8TvE5N4e0AJKl4mjhoWhGZ3kYCb5OkcVNHUcm5ijs
O/q8iKlD1W9XEX7Q8hboIpLuNWUD0mFcUAQqN9iiCWHmF4Zp4NhaTNbjO1KJ8BjCpUfKbsM2wLlL
X2VblpyU0rNsUXBfkshbHuM7mqRFKgvSqtk9rfrPgESlyP3SsPrwI4yQWPqUJoSIoFcdBxN7I9HE
LNr7mnN9WT3GbdY7ZkUjtAwvQieeyCO4gw8ApyjZHG+C0nEwQdyz9yE+77FXckYQSjKWORek6V16
/8gAGqiRszD16zi2RIjLk2KqVKGf5y9UgN5uHKc4fD1l7cOTrmz5EqaZCFn1Xzx4fvWxO4+rt9Np
/Q8Bemy46VlAhwAJV3f5ugIOvjQdRAIfia4AiUyJQ+Ub/rt+aDTj4+OMsxw/TULtj+S++7wV2G0D
2rxdCe3kV46p0EBb0EWiv/3WtiUk4MzuDPAoDFdymogVv48LB4no68fm3rboz1h5ZTnM8M2v8KmX
6qliSEvQ4atyPFzZZ5KD5m6ZuA0wZDz1pQnc2efpieDDHrpVdiz2nMTIhC+u3C+iHwLi1EBwN/P0
bO3QfjF2X+BohjkCkMlI1a8irsYqaf+tNwdivKywYbp784E3CFHCYhQ3ZJ3wlzjcRIEDdMZr0vvQ
no8oMrazXk95zUWIdcR7ZeB0koySQVn2nfn7vNTiZXB6Nn8Nnq5tU78LhvuAaSGTa/aPoXgHko7l
Qw+Hdk6IbFumlB+KrXkKkfWmp0FYhTQjz5khPd6pt9lE1tm7wv7xMALhvFZgZhF2hWEwn4s71dBn
EWLb0vxO6gqT8t7vjTmtUgs4Rdcwy9C/D0qQEoh19/l1o7ZACnjAarnaiWdNKrFWGqqi+yN/YWyF
CTak5TSHWTbX11rEfI4r7CL1xyntaesp+iz/kkSqOtBuBtf1+jacnD8u8Qkp/WhQyV/tDh6V6kJm
rBFEMtbO3kQPQ0yOC9eiNZRazl7oai928r5cPhT3ANzhryTTE4eYPE2Emq1lL0U+RAes6chCFnjB
3j59n/l0z0j4CtD5T1Ht3EGzcHmQGudiEfdF/HYwUwEXlDLV/2z1f6ETfryUkVkdyAVo1dOM1ihi
PdyfAEiRQM4AE7c8wiwdSkOof7M1g3U4zlkLp49npHKbBxdtsrcRpRHXfEEAMzMgRiGJVWz4gFYw
Y6x7r1eIB2ZBM5IgQGEF91K/j7Hx1uFfgzTgaha+omKqw2wEY4F6EPTGXXrn2WsetJsdByofqTCE
vEZ+vjuPP26opEDRQ0UIoCFCOeUY1LCpzhamkBmq2YbJ2fUf4iD5QVLyaJjmAxX8DMMjDvZwc7mQ
cgTuMmTNrXoZYp0qe1m7O8lNyKPwTTEU2P1WycCQuHcnJ1Kcir18h0MrtTjxute8lnImGII41i/B
n7h25NOUkN32crLiKx19r4f2k6iFAhl4u9yb7VEWHaPoLj9CtuZBKPuBKXw6nyY7rY2NZID+ji0k
IiyIxJqVBvzVZncLLXK2tfoH/EyiXZN8mn+Q5xvgKvDP17i5VAk6zU4A4EacnUX8gXI873W0nCdY
5XDD8h9p4Tn+/KwGHQ4G3MP4+Dy5TDfx0/q/oCUt5AZhik2kr9qi8of4DJwsUY3f9MXp/GjWPsyg
m/qsW4a3W3hPPsYMwKvwhi2594OszUykRTPdBoxL/h7pemD3xthD6Po91F5DazW1bKtCx4R/C3XC
K0gCVDyLgvsRsuX5+b8BmemeQZCD5Erl0fvg0qydoRMA0rKjHL0bhoT2nmncuiV+1BNVHNM8RdkN
DXjnTBgPW0QBpTFMJk4OJDZTpSDdtYI8l72QWxtFNXlH5FxpaB9m4SFf8AxH4yl6JQOT8+c92ubz
WsBimUNv0hLz19IHBFVgO5XzxS3DR1YjWA49XfOO5jHhI/ru/RN0QedL5Eiwu0PecijYZFVIGwxK
qDI50xTPpJEhKZ8Xdj1nN+lCM8Vt6wSoYGhDOen+rPMqNJ1h5Xav7YPrkJT+/NZoEF4Pr7Qmd59k
IJVkZhkCrKMBjggWKvTUbO+EAKZ8KlFJvVaCgtVzu+SGHS/vIy6shZUDzdaTs4L7LujWF/llDt2c
5K8roYFH5ZnnTklE2LJGyAF4a51Fstr/g4ButOGma0EAhb4KPMFMyoHF4Q9lpQX3jqRt9gO+c9jT
ItgmoYsga0LcKZ/OYorg6W4kukaJEUeL63uBG+NV2OzXlqi5WVxcGg7RfVsWBS2GU4kPRlhi+YyN
JrMd49p+Vb6nyxLe25MP53br+VZQJnI9lR7mURY4GF+6w9T3j8vgiKX+gR5XuLDXHoRvB4M2f1Jq
XpS48dW076GjCJLFjzeJCNVjYExAvCh7aC9Xd7cPJwoMC5mVlh/roUHaYHBaKibe+hktHWXxyAn1
jNGpYQFX/ta8zGMvCyLm/t4j3u2g6WH80ytr/v5BjERnEidRUfSkx6VkP1+PVXLxZjomyeLYaT2I
3kEd/9Ci/4D0ehSBkhImbTHrdxURmbK+4x2NFIMtEYsKkxyMztSTKDdNCAJ+su/mSfI/IzgZxqRM
1lIBX9GGMiogLk4EaebEYEWmTMNYPyKjT3zFy2auqCxDe4Ke8WyabKZx/Qy8WfAd4HdZwnvHC0qV
OieuKvXyerwAEfeXrW0DAUSKSv+jlhaECBXezDFjDN0Ny+UxNW/aDH+UXYP9kPitB77VOE0ODRQa
AJq/uqk1w9QlKd8Gh1IENvhMVnNV08cf0Ujm/QW3SeHqWnV73Qmaszrr4ADguWOiHEWWQ/bFVzI+
klRwFpKXn/KM8FE2jyqYNoVKN/2ps1ssDQ+HIPSLe4ZSsy015+2jJPO8j4lZ5xq4Fyzkts7vtte1
CXNO93pSYYr7aGeFCPIn2d5aH0hJvqlx1KWK1k9pxsK5hdgSsekShjaSYK9/S1duCZA86aUO/Qh6
PwSWleFg8hNT6kHAl8UkfR4HR5GJUFhNR6F+zn1ZBU27tQ3GsD+EGsdrwCaqMzyhkhRoifQekDdb
YbOxFiIQDf8RAv1DLRytwt1YGGw+v70mx6D3N/zl6QfKd3jFul8BDQS6hzEz9DFwUYtQvKc/obqM
W4Pf/xd32X+4DsyzMxtoBzd6AdWn54D+5kWgsYBBC2izTn/JZZxwBwDhuZak1XdGzCimRS2OuDtJ
3QvceZNR8b+yIzA+W+Vma4ntf32IUuHTlgT9O+T291FlNJBtGEQif5XRnkeQ/lukfzmQ2h5VyFYg
ioPFJ8kpm5Un95qfqseUygc6FxGu/gSamq9t1kvqkpJKLk7wUrLCVoelovGUhX4hXBhVex4nnoM7
6JFdudJcC3tJ7tDpCuiRDoVMPavtcw/CEZbKuzb0d7hQxfOy1/d8+c+XwCSUJ952uWNlVajMEyEE
EQ1EYQHdQ0xUt22X43SGMQh+TNged9liR+SPCtCCT8eMO7FVnzk6BH+pxmNt3RsdXPj3qWhZdSBa
eGJUE3TjxSfng2JG93dhIqkM6/UIp/5mcNYiJiLNEFjCAV58tmq5hA8y3+T/lurhTO98/BrbWASJ
9axF0lHY/bKgBi4afA3kx2kFWWfLNq/HYiEWYbbWVvHqqfj4jOk38/SdZVvDIOZWywz1paGEgrdq
r4SmqWntwUXr9iw4Wo2wbxBCZ9jYzUs4r6I0NlXGWVNtzhJssASD5+W1UgirdqFIPYBszQH4txIn
DQ8U8Ly7O6j8IulDybQwcBL8nprlnIf4D5rrPjKSnZj2+YnFq9UqihxwWhp9lW2SQsVQRLq2IlM6
2Pq3tG4pVUD77dtBnLNBotJVPMdRfO4DuspMRakwPVgB4AowPXKW+EeLTVbjfWr5nq+hnFGsNdvE
ocdWdihMJbJsFSn/74KnhQuodfjiripxOJyFqHY5YCZEJ8oF6T8HeppsHBHA/y+iQDrA7+Xomk4A
TcGpe4+9E3Wt7RDvK47s3zWvqaGTB92ikkb9hWFour522ViXpGo4CEux0sWZ3UoJNsyKWFxzKjS+
QvVYBwpUgC5DUP1ag2uztuWKJ6RAsmg2f9fnFs7tVDoGyeDhyiVH1gp45R3otwVDMp7O5VRMVxY8
GaBcpG4OWuplRkkcv/HaxMr2hZ1p8GYzb0fd3VSuT5MDyvKMZM0GnQ+sKIE3Awe1FBAXFo6H9YoW
Kig7uJ59MX6tOZy76XHe9pO9X+iEwQuFUkLbAeEwWfrN9NEIxh/qTsFBMc4d89bs2Qi8qQsR207K
PStNnKrm7OEe1a7BQWxB+l2LB4PVr1LcvOFC1+JgHki70A817CMJ/HAAbg+/KCea7ywSykv0oPFo
0zF9sjH5x7CYO0m+85Mjv/U6CfSPamLVLTOnmU3xrjQ+FtGqh6JD/yPHPPvLUpWCPRrPE6521yMX
fiVG3Yv83RR1xsLubS/6JWl+Pvc09+K8guIV7l1kW28CAUfigynz3lo5On30+0c8GUI3c1dh6mBO
IDcLaZF6eCfc4o1S0ObExMq98a7nsyw7ahEdWaVBUu4r78YJ8l6g5R0Bt9CUErG0Au0v5IchEcEF
WJwgh7mp4h4JgLp0yx5Y4RA84Fbg0Ly6Dbua23ZYo63xV4h3M6tXvb1wmvkKs5xKiB7se2ZqEmDX
mX9NV04zgAaGMJYCxTlxzufJwf5+XXW4qRArz9NowI0rHTNhXkCvK1mAVBRQuxytLhUbfsEUSizP
B2bI+l7SzD6gy74vXmpPJ4ggnI9fqvSnllbY/7l2ZIUhCbTBQ5E1W8eR0SX92j1jMGrbvaUUppkz
a6oqRm3E3GYQ44HASHuRHP8vn9BuiV7ync19d5ZrJWTWy7vPyzRxtATPoGgXsGE8yv1AMtYg90yf
Sbts7R0UxLhquG/mzrmOGrczWoTE+8cgPdtGKLEPQegbFpKs4UWsId4mxmEt6pYTvblCJ9t1ddyK
Z8vTDBk96iPyFseXzNAzCt0LmKOv1H2Lj+fMXdmwFSZ06xu22z/nKRWT1OSikLoM7/9M/cwynvD6
9+ZVRz+zYozjMuFVqs2Eu8iA7531fBuCDPDJP1xJhJ8W9ZHzeDXedsUGMjOFXyiOeF6Fs+cBoCYm
MlgwK23S7NfBNr7f1LaeWKE9asrvHqmXIwjlBAaQ1uLDVMIDEHRdUQymkFwpp2THFoKGnbJMMn4s
5aC74H9X7qjI4RuVkkrlLFl13m7Pq45U9a3YvS9XAuXHTPLkrfgt7yiDXWvUZiLbQofZZXQIQ7LC
zwuqBZXcIjxb3fifie8l5WFUey+9J19ZK8WFtSdTtbJUVap/nh1wwxp+WUNIcmeUVhE+1mZt3m5K
lBy9FvAOYF5wbCJf92c7rdFPqm9aG+LJrVVw2aU9mxirnJK/rzN0SC57N5qZIoPJCz3/BJ3bv2YI
fuFm5lS/PfIFjrqJaXmPPUnEK+TMmYiTpwzmwzYBFEGHP+FbtMCG2ysE1kiHLgvHZiOLyOrmeo5V
TYjeVFSIHN4z4iESqpQZh4HppMsUUvQKgHyeiGcG3jrwjhPERqYQ18hFxCKs2cWbJ3lGT1IO21Ro
96K4Th5OFSHrteAsucj/PdxG6sj0v3bEgqz/005j5be4RYBeI4EHbHjI0Vrb275jwxjvUthc7mVD
AxjlH9du3vz7FX/U2Z04UofVciP6F8zKmcHgkiEw7wqhSbDdncmeQGAhl2WlwBDfUCe93F5Sbz6K
hhxsNfqbouF/PlyLJ1lTiHrkO4CXHQobyxpS9L/h6PI0UjIWyas4a79GClL+UF99tzpprfWYXzso
d5aLHTbYr32gZ8zGriGiRlkHcE3R/S2dg5A78Y9+ysIIOr7hrwS259Q7M7qTn7bSlINQDLNaqZmU
U8zyy/CtIRCBxqbNd3epQNkPyZtqeJ4d0Q7afuK4QHSt2CSCV/Pe7FQ9w3YxvupTpkonYl0kE/uj
lePXJjuD5AQk6uhekqBFSXQpqGkJwGPwpHfXHsrIQqG8IPIve5IS/w0n8QwsQEQXt/P+R7he1+5r
IWwDmnD0IxswDp4jzetsHlE/iQ8OLyVPrxsE9qi9Ee6wkQGxB6ZIFD14/Y6tEs9032runhotX3Hh
aXozZ5Jx4y3BR256sgT7BMymWoFQLyfCKdup8pG6tL1gMbM6j6QY5rJTiR45eoose6gUqWj79zp6
QuPA+7ZSln3WhsRQPz/hdpkV2smX8xccTqXsztek8Dbsz6o8N7/6z94jIIgWJ7W6zG7n1jDeLa6d
tJ/sI61x5KKwDpIqlHlrwTmhe4VRGL1yX09bABqCfldUT0AHSYJqwzv5OQ1vy28c+Rnbnt3k2aBa
XXkBYqV+lTIshW3A4Q2vocxOYOruMa/Kdr+OZVCwKmmvB1xgmrKCjmuwaU+dsvNEwGvP0Ni+fbsg
tyVfY6zg31Wppb0PqpqmIB/IghrWFMLqDZYKjFl9GFgw3js1hUdSKTktJfDpLHx2tbaEgPOYZm67
ili6xlwkU+3agl2cRpMOe7C5i/R7Jusu5SRX08WM5/UwctqN7BsVppyGFB4US8nK5X2FEirduENx
pbqh6FZmI2PRXajTytO6j5BKsUK0gbJPY6JKdN0ry+wd5HUygSVrdhjnmpIEzvG1A+0d/Q1z+08y
1S/5vAcxPdCd+CQYF49S3cEsSNNKednV5ZFjA/O9/01BNd+Dw69IQRozy6OZxbhkhTFjrx5Gce2Y
VyUniORYGAXQ/4vIvZ6CkjrHAmxEX/rb9pjgt+4eDbVeapIrFT2M1+aoeEeKCY7rASIB7uTuMuVr
gyx/7GbenzLvcxv/AVnyWERGrbB5+G4VRagTG9ZExXODGnqZ5raF2xD3TGvD+BdZI7BBO3LmlkLH
9noH2bHz9iskF8nDkO6mXGAsDvhwT/3+SfbmfgON2zvHQKzdltwi+/wruwAbnx8Hg/uXaY4zU7xs
YeqCktyQ9X9umSSpKuhvFm0YfqLLqXhUM8Lu7Zvyh6cUwiHbMdZ43zJXVayUQcGVP0FW44NOKSO5
63Vbn5UC3JwvtlshoxdL9qWG896W/KtBKlMHbo0OZ3KWGOf7dabF0Hc8P1h8VACRt1rpuNydIDRA
5wsOcFgT+ljfuPsFbFvp0eWMWMaGoB98SjlnCWlAh9SKoxE6xDEVt4iabRTOD/52U/D/5tyJ/lf+
ISYogLQuC3LKh6IuKp+GDkh54T4mpwl2rOVCBhubqWuS1HV5PCvcQljUa19C0rmqRrCYd/G44+b0
aK3NQ2XdR+5Pdmvzt+piSQOwp6bofWyLHEtq9mRJBmjHrpbbJXEuKfp/zZzylnfNR3bqj73QbQxu
v0CdYa2b8DuRtUZca+mB8dvQMvn+RRyPTCD6BcOu6RSok1HkX5UAb/Ki29vFcarXefKN8UmahGLn
3t1/iszsmscJ43nOHJAHD7F11wPwF9C40xkBoicGyktIA40OuKY44C2b4jfflUtb1c2IOO9FTeMc
ekgHEPMpuzXO8E22twe2nN6YDBwGdXz7vCZeZQoUdDzD30X/1u69+y7dODjkUs71OQbPZbSIXjsS
lE0SWC/pQ/IjP5hTdPHBut/7QkwGFWBmGzB/Qb+qS5S66RQ6D5ESSe9PRfpQbHsM3DYkl8KohIAB
d53ksxzFyjjO2bBBdTRcMoH1P+hUde9vrFwULeBK8bwlPOEXrR86oOjrm0LczEO9ELh9Bw9TPIHI
SYj9E1nWwirvdaIjxZqKy9dUEZii49IrJ6LM3LMsKS59btPJivOggMb5zsKpLzcxKPBSNBULhiRy
JnsXKWdqq/B+sWhKAhRYgOYcrFc1Rnp2ep7d9K4b62449nYWJ5C3MxU1SotWHP/UsQYGzskEBsXq
SLlmSMiXNfWruRtSGqxQiIJhBQfpQEbQSSpYTDgRXy6jK+ecEHGpiQWwb9PxW31T0FTXqDOH00S4
OYT1ysjPcRo0hofOVpWEwFfJwEkZpmsmex+7GK1D/e1b4QlwH4dZl69w6Atc26CUqA3c4LtyNROb
U+b59Wgmg4c71UzqiYvZ8B4kC24SIigKM4vPf4qHQdPCHTWZFHK8riAjYt9CIG/NjiQ+zcPPyVDa
qvho9pzERkVBYekQwRm4mmB70v9xZMjXKWa70olfpLdwiSvPbal4TXE25EJSmIe++xccyl8J5udq
CwGtoTjQs+pP0+wFMRia1DUPQ6DVFvo14JXMYmMMSBWOk5Oc+1ICDYrmiMwfOcSNEIDeSa/sOT67
5OS6cYqJ+uQjtQ6A/6hKHVHs8V5hnLhmrHTYRk0R59rhMko2syrEUxto10n88onlLspElYx+4Q7D
sdOQyHtvYrKywNSgH6iSLeCAjrraDNa8aPqq6482S5ecKxVMzhfAr9sM2BpdcUSEXP4QWImlExDo
/SWFLNWIltT+GpU3DtVqRwn9fIx5We7tgkU7o56zXDdU4w6FRY1RQPlTe30hlsKVR5yAx8YwJ31h
UUJZ7oN1Q6Iy10aV7vDcFFoOU2ZcQjhRPDLCyGk6poJR55rcg4mpMpFmRcGmK6/jFXDl5af6rXmO
KBx4+OatzlUhelY0n52E8Tcxv8vV3kLzpc9aXjZFrBnvofHQg5Mys6ERYWzs1AxTCFCQ4XqyxHgX
7Icn5rS/wS3BXaHF6pXSdqWQqLhe76of7c51/dGPi4z9bDMPLt4N/MnKL06aBr509E/Uwq4MZWye
g1ncfORM6+tsEUUwSsn2vvw2pEBCSbYuQPTQAz1hOw1o3Zye2Rz/CDM2gDkgiwMHnz+0pe1amMmz
FWJDeCspuzf2+zYH191+1rm+eH4o5GFLJF9WkDYYD8p3BCzvnnlGE5PAQ0MH6l9ppfOWNcIefgUc
lmOrP26zSqVB0+kN5vIu0kpzCw98+rtaq6l0Z3fGKscrlryTGKo/qhcdUq0Si5HX95K+/nBKAKMO
G7eYh7BqVwgM2YgDFGeOQXTVxMBVT2XiDLss3YsXoue+70Whh95iPSMxgRave7jiBZmPxOEK+w3o
bv9wuOlnUK+BgzQ5zpONDUcf+TN0J/tEWUSG1cBmAsA3mOk+8OHFSb6KD7Mc2EfErIZnRQXb6KS9
GJ7CtDG0bJeaEtJjSEbS4nigEvGib/67agYbpGQ3gCXDmQowbLTNy5APYoF74TcmJH9jQpDkjIur
t/khht10KQf2EZKjkzskrAA4TZJTGgXOh1oJhIM8hFfAdT1LE3F3s2Y0mSp7cRH7aLaYQ1y6lGu7
cAJ1x4/hW8zFLTJzzHFG2mlrj/b8kCXAyZBx8KBNHFCcYqq5HPjWPWuA3bJxLnCbWNFJ/cIk0mmm
rOBN4nvKGvnrUgc2yTAVHNGyIXFsyjB87CYzXTsDAo7sBBZzAwN1VODNs6xm8PMem2d7abshuXTb
lckohpH+OeDrF1KN8PDyXj9T8xRv04abA047C6hw/ZUy4gCnsTh90jYgLebNp/H9ewzJAGDbaZJT
yqteUyTDYLxL7nk6lNqQSpRqFvb++iudDKjoLSibKXAwgtVFbbVImpKF+oj0jgMXBEB6m0o0XrSh
0RzeRq7zbjdoYAbUZO2ErJSE2L0a+OKONAq2bwG/kb8ZEd7B/VUkjKhJ7s4xjE8gZPgySmDz3rOk
xY+eCvQrbXB+Rj7xeVg8Hy37ufkJKcZ27HNp9uoTtStCP6DAaxmyLqHAHLU563+sSqYeg1K8Trzm
aunaGdzhhRpqk36Pvmwe5I0oEOraqzCNSXB4+tYv3F1ZO9zOq8jpFkkTpuBjWZgypgAeriRFV4SD
BLYzZ/l7xDcOKvqnCur5KgcMSmE+dEOqVx9nUp9wpz/PN61SsMUX8yqiC6MoePfCwLiAHuQJ2GDN
thsmd6EKMk1UeaVCx4KYAgDfcJu65QXmUkeHUyMVFSUrkaDYVgn2q1hskG6NjXePW+hSNuv5ddX9
7rTfX6mWWvI08MUOQdI21SDsIGvjHQ1Itrps8OfNk2t/cvyc0FMhW47Rd1ubFXfkNg5v0HquKk9t
YoywfoWctIDX+ImiLf4+ayaalYESmQCuYIYeeN7LgYDDbENfcszFvs1Bqg7GsGISohdaO6UYAh6N
z40TvYb2LOrStGQRN7EiRhhxH+1DN6m2VUW8xqtsR7ADCVe8Bzlv0/zpuIpIYKp9xIXwiqqiDgQB
HMIN2CLPED3I5st9x6SNQkwDQGIWu2EdoR8QaL+DhxDTZbctjGP/7lomG312QCz4tEYgy/+NT3Vj
f0ncvZFByc+q8qMILNxsWgmKOxgPFhKSSTs8yEhAGYz1983KM1v/g+j1Yjg/AtUvXNG8M3+vpkSu
13z0UMWA3uQuZGZy9ylsXpPsdwfBebXUBhHbF8a/y/aM5DsXBA9rhEQzXQgXxX3zR7IC4pWWw3ID
Ox4hOSpng4gJhJv22OO2fgjzVCtgfSKgSqdrDvsQbvr5wqPsTylc6/I29sQflQBdD3G0AbfF8aCq
cCa9LmT35e5GiJRAp5MdGhqz1qbCTAIbF/ZWexTZSKm9r/wwkLvnwQfA/RvCfzMcd9RxGz9a9WdI
nyI9+1qxAnPtVEAv7MNliT/3o2G7t3CTPJwbBk4XWxrvxRW1PTe0G0yKtkrfd9yxC0bD8pnQH5Wo
RT6d6VOmLxCRGOo4aiQGlv12izvuTmPm/GcNBfIPGpAvTOdvS5k4/6NZYWj25lax1PsvOlgFg6FX
fC9+/yGpOVDjRQIsN3AOEAIX0SKuTTJV//oSXV6Osr3UE1pWoAEC1E31zClC401QsbU7vESKVv7H
nDblA97SCA8vnFMLVuRbOvK8uk9aulHuj1WMHA3F2KsDJVZ8bXfSG7KbIbqrlrWPSMBiERr/LcSL
CQL2d6Uh8dAZeiWlq/vwAKkQ8qpnXS0KGe6yWoiw1Ihkjm8nJn+MRiU14Z3o6n8OLpr3yw70QWAq
R0TNkeCydY9QTgc78QuOuQqsgqdHi82ds2730A0nV+HZzgIPiUyqy1yR3yJMqIfTdBfe0Byh9xjN
zGY+Ky4ZF+373hBBbrJlugRdRRGtMuYy+iy2HGSj9wY1o7iWN0BJcx8xJ4a5FisyYJ8/m7zIbRr8
95e7j6ktcfS/ZKkLpniXyeFxOJM7NsNzmg8P7E++BeBzd53MX/dYgvBBHL1ICEqoEhDjqwaeSATk
j/OTH9pPv1GrdlKZYOpWkhnw9ki6xfM3OuEyxStxLcOXJM8md3L/gJYZHvlytLEx7CpXHCf6rLIn
v4JOs3Aj7WGNN34eB6NrWwvItZ5Jg2x+n1TtL/imyXLhSmiVWq6Y9WHQ27LyCrO9LpCR/Gwcbijx
7In8hwRCeYhMdlOG5w3VldqIaqvnTYe8jcTJec+nKAu6LAw69dTFJq5OoTHVJA687WLU/Yhoe0BV
LPU7/ZzzJA5ZcM4LS8LKRwSKZuy/7ysuMnfi1ZDtGELQyXM6AuaRjNqhML/axKliTXlI2edbBrT8
EG6tSH3rKggyoLayh/q6+H07jgFV4U19Vqhs2qEkYQgCLBrImGdRLGJPch786S9kC3IsvF4WMKHw
Pyo5Mcr4xAfSLEg+B6SdzdXCTMBpA5DFxGhDMSXcsiU7fLy4LDth29ZLaz4rHWm0t2CmswIcsPCf
M5eoocIC8kjiAdRTICauUDwEA5BPGyzlZEVRfl0/7BydKDZss/UIYo3BdNOQsQ3mHVi+fhUQI/if
q108BXWThpt2+JtM2mgXnPN9phAuuF5T33XLJ2yyr1k4J9qg5sIrC8hnMBe3WQhJu8FXBrmWoe0X
OwZnRPrtOgH3j7SsP82S+BeqdWpz8Tjw6icpRC0go2GrQHi6mz7r7d067a1el0ONa0emAN6Lhs4X
yT7Cl1aNyS/IVWXsFomej2ed4bl0iPIKWuNMvqrN87nY+k1bqv/W2aNfjKXjMql47P0SF0m1q/zp
Az032onWtIm+BMVNQwY4zuaFZkpLMpDMJ6/pM7oFzhHC01FhMDJaeSSamJRPeyLskr2RdOfFLRdx
4rY2A2gxgmTuirF0a9DWYQGef5CjyJskfcbr0Ld3JnGykJluk5ZNOenPtSPOH7vc/Lh7n6lDQPkT
ZzbggdPf5hCbExuhhvoPRdnmN2pLoaY6HBWKz8l+VjsZvHGauj2uJLdGyLg/lmQRrcx1i7atrSdP
4lJHEZ5KtnmSRHSYtxz2vKqr0wk6hcuNfECzIJUOtahw+T4lsOLveEam5mWez6T85C0YiOCWe3Ru
8myNDfmNsfjg2+vyVaxQMjspg7FrWhQ6yFOzQLEmzyL43VGv+rAlUHFuw/liP2J2WZQY9q0xoh5d
PpllWSzFcnGpB0LE/eA7zqj5Tvfqxh+z2D7jKwQ+rCGPyn2O+m1hJe3W2M3vs1hQp3qE3KZKNWXz
7BNIjxmhQ1gA2mAJquzmWo1JUHH85Wht9rW1Ny/bD3fbS1BaoMmmKpUUvjYPQQUQQ6jc7rESzBqm
/QHZGTiYsQ1LTRwrhtwAK6xagIQYSAMqOzI0C6TIJaBXqM2QOyNjBAOEgE+iSsYZU++rTYgtgID6
zAqiLDNpTrAslelGIaTi0XxpPYPuUbIWxA/fo4ZX+nAypGOk3nnrhxytEUZHzKgRragEL6RFp/2I
Y80pd5Ps/Do5GCdy05E+eXpsajfPpTd2dXH3+YQEWgCltQT35AfZ50qPntc5VnFd92yOiINku/tY
G1/vOeu2mt6KN+qaSBaX3t0s0LekCA6je01GGX4rDnyvU0dMNVhhjouTcBJaPmZMPDbOG2uEIDcu
QiPg3KmgH7IxBAYmI2OQ2+oPtMVxwSw03qZwyMT2RefltMEXwrFtTnJUCtQCbWzBxCB9OSLA/YCC
lDpmXnIaHBZ5l12JfaEyqbVmWMK0Xr5Ukvw6YJ4Rv/L892VTlbPfrgT/tbX5MFSsTuuIHVRBPIM/
QPnOfcuHVCwtS6la0oL7CA5jC1YZ5HGvdsmMtSzDW0osb+XzWmsTyGIXY2pc+cQuzEXeqoZGOw/X
d9fs5bVNQCQ5ge8v+7Di4cEiKX3CHTaI5MGiAin0TRVvDnJJGkdF9CyTlc2UaG0E8cGki5AAW1KO
5koVxt9MUvto1AWbetpOmUbPD5PrOjq6qycDAJtDi+M9hGzQN8YTEd5uR0660KTSbqVH+NDRJ3iG
sV4LGH+TTJX6ruiv9ioCy/36Ry4cjLHROc2tIqAOJ1bDCHdVa8HS4D/82zGjdVIjsl8y6zZPNVXA
WKJKfdJIiLuXkdPNwPI40HcNB/aQnreqYPkP2ee7L9lHu/MOFo4sE4eu6SvhSq1xEGuyBl+qZa0u
Awy7AijQ4CKviSdKYbDT9nuoCJ3EA0foAO679iZfBhm53BpB2hRhqfofWIfYdCDyP0lJn5ufhSwt
auKiR5WuDDgngrMPQF16KG8WcjCc1bBwrxg1Vw92SqgFA701OxrIz61n1RqHKn9wynQsrvtv/Vxv
dSBPZNTkUkdVCUj9leDLY6G7vKuBtXFqL6Zb9bDzImBUOOvFEXxgFbV/Aq+LylmyMPvy4z+4PKbE
Lgtk8vYAjLKF27xOqnuAUdYkWFY0BNRWaj0sEPyYTaR8BVPzq2Zmuss+rd3N8gZAF83w1ZtU8bdL
3580j3dJrNIEncO2Hadu0dnSBINboeBXh/DA0+ac9Z2+iUf5DOqoZ8SBQapdo4DKlNwRcLSlHxUv
GQC4DiKrd2Oem6KUTWPXR0iiAHfjlgJcrxjjN2ei0igIGAdjXDRS8sKFKcRhBYCKjxTQMfdOfcfr
gk6law3OtDdAByfzdELJ0yT3Sm+cZyc7vBAze/H1MbnhgsarmVap5KADDY4PPxwQM/IdVLPXVBOC
qFGQp4rQtYkmx/0QP+NGKaSPl9CjtWS9vRQIA/1tnP7tTTAVi3zos6nqRgkxN7uL93ow/VmvsChY
LFMtuWAC5P5wodBpE35T9NJ29VNsNhN0mFB/RulQ7Aux4R0Hm+WdivDb8a+A+j9zuLliXzflixdT
0/gIKlntvS8UluQbG8bZrayegxJjBACpXhEqXyH/46lTv+aYVgb9qJ0HLggnSJqb2BWJsg/79llo
eqE0H/8+kgAt2lVInBFxAISDjfw/bpoiWC2EcPahgpksX3cyTDyR/ixBkPFc5X6C+d68XiGSIya+
E3B4q+1CnyeYz+XIU7qZ0K5lxiyLU9SF7//B/04XbZ6jp9bn0AwluEgJEnOnPvXzoScxcJPKDAni
v2jIWOWTEOsD8ar4UWqcmD0CypMIuZl8etpjtpnKVYa6eIz29oLKkkqxmZVYJVJEZ47pNop108Nf
yDEyUcyCDfbUXCaCYFD5rBOoj1Q7YcScZ0QbDc+l2XOVqBHRa9IEFS6K4VpU8QygcX5KzJ0/vQ4a
rZCg3+qssLeEGQhYlxVRe+TON6f0YxMRXmAtFlLpkHnsgnFAbJNP9+IX+7p7+lE9SmVhlpoSH0BA
6KD2ypGecCf89PjO9YdEI1/sj5c2uyto1B0rBR4sNKjZsLvW9Zb13IA33ieFBLFzcaN4T26cGBPt
/UnIJUEXpmUKCgXBV88SaUGVfzJgogYo+Oq+4oV2LqHvTOO59KRtS/HRQAEWf0SWR0dSuhRgvi76
gWQo5ARa4BIZCS0dB4btFT8gO8qkLAeOpWPQEJPLBhf1aJfaOk2ayiQUgvw2CWwrZ+pKIm2MhT+P
2RmjGhJWkNV9z3Jn9C3lOwxbKXpG9iPEtBvb5Xy0CQa2WBAQE3h08DTldOLM0eOigW7QNibmjYrM
RCaqa2Tzenr8JMKyaOzmeRSX3eymaQNGJuyYUwYsYfRAQiIY6sEAfKT7FgdSo7ovCR4WEXdG68jK
9iUkYCzJ6353cOChgjeIMfMcEVB6vTBUEnsUhQMIt1tPWsrRcma/ChVhmHy9Nr7lqo/srI8ExNP0
GxSyE9fcK88cLa7rsloFoZ87YmItsV/Fb1J8lXa1rC4it4oIR85PnV3QL0l9ggItRrQNDZexDMIW
+KHXWieAe9W1yiTBH3y33UKM0KzoRLhSZj1toY50rEcTb095a0uIJH0y878Uhp/rWolA2GmqLgcm
2GZF6zCIA0h8649WtU2N22i4HKAH+DhyTC7MY7XUVRxamsKoF2SNX3LWqhQor8RK/GjbiKM7BTda
N25DDTXmvRuvuiuSv6GAtebegPXmQjoaxdnxW8oAnNUpiwYfD4U2G0JEGLF2KqeBTPlnfj9EAgG6
XnJSshd965PvB2jAYbwQZ3nwqsZx8QA1Ekwxumv03by28TDWF1LmFh/A8p1UG6f4LvKIVHHumaI4
fonbQEpf8BfxrctFRSN9MexfU9XBpcieWc85Rg+GmySgvrxV2Uxpb7lCnQJSYsg6rdu5+1eJuZVL
CDpM5cZdWYDIit9aKdiwagKzsaQtovndtq09oZfXZY20z0769B/YGpu9VB8DB/Laptn6AZp2LZTs
DhOQTV+dN/uNcHP+fUJXXnMnqwy/fIMiSR0VlwurNDqulT9UYd66r7O7w5OPsrOxpNBARx+m1fPX
pjK+kGCSUuBPnSLd01elwmOL/gEMQhWDb3+V5GczLafGp2HYgwKkbcmfOw+JVEl9C1O/SBL/mjpu
Ifs+twfWa21k4OpOk1C8mlRQ+pxJ4i6XzK0IF1kNIYv7rJsfkdCzivTf/VR+rPZ3X9dsb4/GFVHA
gYZmWgyOU7j8vANPToOlVVRoFH/qXxi1wcMDifpp7Dy4uj4JvG9/TayKMs+0qfCNHRDmZ8CQLtjN
jyV6mZZXE0rXJUBlPD6dnmMp6tal5pPSDf6Bf70Pb6UafB2DEQx/YRW46iLaIrVD0ywrFD3vv2Pb
kgGEUP5WzxOTcZrfypO1jEeeSyR2atthmeFN3hPoNqRw+k1fzi2nDyt+0GYtNhWUna//LMLfx1d8
1tKh4cmXJ4somZHwJcEI/sa0QShh+viavPy8MOM0gzgMm7PQ4djsFRnA3o1sHT/XnArd9+mcRfiK
jM53WkpXC7HNlYxy1CHgOiZavLNivwiAb7NE5H3X4UN2xAwk5Yfdr6NRBthS4ghTUJzj8TGo8mA+
GVck3VObUSP6OqgInXH/QlhDr+TlKVyoyGwQt7hk7DIkpLI/KLpjBCXKPTDq9ymb4PYUVHuSDzQG
1zz/UBEX0qqX6UcBdq1CQ9I964dUR36BYdY5qpItit0uzwv6/xaf3uyWhPCK795MGqhgC/UC+i/E
taXO5TQ3za5HtlnipSn7ZrcOpnLpi22v11n1PUTAkSdtq2gowrXQ5iM8vkO27harmx54ZNtPzmdP
uIKWK4AzkFHSw29Tx6JjC3g8VtzbkdI2W/FLjc2FTrNYWlsX6cACmTzM++zVyJd4T6D5R7nQnn4r
FNr1TdI5uj+KKzegQtICpaNy46GotZYkfm55vs72AXadr1NCALNYHW9QjKpHrWoB2xYPsDqDFhnj
OP9EgXv9qa8QjFOjZT4kxAKJb2R3JC4WyxfnGkP+3X1eDfLhvJEEPyFrVA4T/DR7xSdOva2cS+S+
PEAxaMwGtD0vjLNYihLQlEmc4emW0aKCw55Ia/ZWC/IJoPH6Pa9m5im/tU9OhT1fz1p+iqHw/tF5
I9rXdTVG+xQJeVauVY7tGqDwz7YdvkzPSwRFzGpQ+PCxTqNZzuAenwhAoQDIS02igQXFRisxBVGR
IuHKKhU4aIM5RJ0sJx03HPeH97pDCxjCRWe4HIyXn5bjDU1KbGY9WPR3I45aifCQJa57HcjOpNBq
b45I/FTSUu4uSYnYiw7jIVKQRNm2L0RNvShL94N+wqK/DvH2umBwhyAiPqRROsPAhUTzcgB9h0GW
jhXb6mvewURjqzvsfRvhPEzM5gVebRtyrsHKdgpzQkv/1wBZRsaZtN+/uirI5K0XMXMafOGZega7
JU6sSE0IXQxW28Tjk0RvtKmW0IeWp+ZLLCBzkvMx/XS43GTzjQJcVNqd8iPpM4cKJu9qUkjIBg9q
BS5YhDm7STh5j6nuWcvACA+QoOBMs7jKbgf8hgNgXuTEvLOf+RuCqGsd8isxcvBt4pEASUxzs29A
kQ72Wb5PqnWw9nJxkgpMixclTVd7bhjw6+GFGHeG4miqcI3UCiGa7Ai+YQeu85uCLx/SR6xK102u
ERDotrmnPF3NhULukrf3W/Imt7HL0jMwPYGjTzYRGyoH7fWsbc0T8Z9Q6MZ5Gku61S4JOT89HI0z
Na41Wh6AhsDypO5BPjjDEq5GKtvYnUnFV/TmWIGd1Dsu8YwLVP+aNEWfaQ/0L/nSNC9VAkHIwXxe
ygkB0R5KlV9smaZOqDhKVN2gDaxNDZzmuC1lqiq1fcV38QaYHwKHsNgJPMSZQbFYXrBfUdabtldj
LBiApwLw+ly8jSrbukiSrIXYPHivJg2ZWx9qGZgqviWIFelK6DSzLrh9DyHhN8jtErsjTkEHRbLe
e9taxf92yH567XWGXYsaGLT2WlrAyWZQb40aYN1nt6hsypjrHfBfPqElHmasRRdWqFYeY5zkS9V0
eNI+QlVhwFf7NeUXZYJT6jV/vkvYItJa8FgrbFrgc+IuOsJBp3zbyzoF2JgMQdaIU5KBu3VLsj75
iVGtSl6aMdtvqg+1zWLnjYDtbGBvgEOEjpwx0zzChEEUuDjQRV/ZLTVK0DdLtxlkbefL8iWXeVYM
LveMqPV+J5EBP77rwEzzOZ/68RrHi0w7scqj/Q01CYzkX51i3BAVFsKKb6lngaLZ0sN+QoH6zT/t
32v2WDNWdesq5uVU3fWs8+KTuOQ4V+uW+L798pOnJvYj0UipWgFdHrsKZwb6eeMD4UCrrwKWagIr
ky4oWPUT8AiEKmeomL7NeK74dvrbEGY2Mq/62x+oPNhPbUfZpJPB6VD26kO8TjNd8rnSQdxR5/w7
EOA+7NxzF9y3x19PpvmCArQP2fbPN3SSZn9fIv3zbCfaDnlSw0wvOZPV/cCXDA0bZQP7Uuc6FWJu
cCU/JXm60js6vFp50lwXIru88GGqXHxHspN9isPHE4pnZSiBIP4pdopI0ef9Hemgk/kJUkvNbwlc
9ZQNkSENl2KPb4/XdLwo6E/bidFAspHLQeAIwuA/hg2kSjwLoSBKCcXER0zY8DRjobHY8ji1khQW
J0x89QHC0NDunPa+eOyh2rzqne+ccDWbIzOgA+V4/2LoTt2KVId2bQAwVJCicLTdARIhcDlTMuGJ
xcxBa+UYxrgJzvQu68mKKGfkzSG954OirlA0u7EcvO+hjll6x2CcHXMskb5KPxkSVveV+ng4UO0r
N3SJsrkq7BVU+vp3DtisaVUipbvNbsmUgU8tiETHsNoQY751rHhdWCQmp+5DB7NiAqMY7LlHMiKL
UxKw/PWWjuln12hnSXEL9CVP08lhgoJY8urhNVHhRKVdBYKXJD43/JyUvHD8nV8eSrthHsdpDvPF
kKgGE42SI8QizhilgySTn9u+WfWUa7x9OzZDQL/kShHStCu5v2dNj+SHyU8LthE0k+uksMme69bA
xZLVnX8qGaKDxDS4WOoLqj1USgAGVtaqByqRgTi+IeLoGJFbuVLcO2WxNFqMAzdOjObfGPLgTCor
PUbl2QX0Jb3LmkG6dXrRK7BtMqn9i33zZeIhmvwHSBP86/4RZyKXL30COYVCAMVpdRZbFyi0Acw6
eOovyEt3/7AtBmAu4cV49UqmfbZwEyaxjb63Ta8xwWptbQAfWYd5Mdn7czAZNA6Mnjk1XfwWDg9u
8X/+uO8aO1mk4OwnY9CYdXpSIuDmG5FieRTf5QSTiRpBp8KsgV3MWnXMyPgKQqGL9EbPf6VRYiEF
GoRqwVLLFSHalCsCEcoGAuxUKtbQtPdXgWVIODnVgZDUvr4I6rcYW+/4U1UtArAuU5A7NyBiz81G
9SU07YT27ZX0J2v2G6g+jYzSgnLy/uPIsTm6ftyIC5PIz2yxI/hHtTxUt0S/501s71zyEHRSpKfm
K77HrMSxc7XOqaixQnJzMOToCLOJdsZs3XA6VhL3NCs6Pp8tc559TReJAtDRFYRSzDukX/GX/s7h
0cklX+sW3e2ifzu2FokBktepKpqNDjgADAXL4HBsYj6gh2tAh7Bm6EY6X3TdMLUYyfyDe8aqH8Hi
h8U4gFum7Jd9J60oRRDFejF5G1tBF3AUYih9EyrBgCW7FAvXEnEIvLg7CdjvkKT4DX4HCd7Mp/tv
Djgzix7UFi5Zczc5fE3FDt6M+4JTllE9OkoxuNw4y4Lr26/24lrHVcOB4PIZ2mv4KgnKE0ZSQ4M0
dLQ4DPbwc0K0apv7YLI5KOXQf/4zg5GYQsN/iYaoBb0RQOwrbhJKINC/bPgmMiJ1PEjxcvhwuMbw
wWPEmy06BCvqXUEt4EDXVB+1e/R77SkXaU8YzfTr7XiNfNW8t+ejZVhMdtZcoT4qV9gk9gMbxruk
H5sBNCOoAbhIh3Ep7yLSbLdS7bp3m5JM5lUD+RRsWJkB0kZnrwHVpB+ecZSQ2ai7tl8x2CAi90k+
H+Y/YVXBFH1Pm7rhE1A8UVkksx4HWJ0h/qrfdaTkljCP1ZutBqprycAKIA1q44rMDPN9NyLTEyOW
yKtKU29V8D3Bb75BnBtuQUl6oxMjtK+efEGUufx2Ca6+YO+XFrOrEayIWo21H1iJaLPdDR6RduVq
VsvtbOWzVlKErqeo4WGqlt1xUacJNSV10bxv/VClpPa+SESCJ3LiqfRWFq3iQFJ7tvoN3qWRQNlw
HcI38yLTqlJYQTyeJpuTjyB3S32bC8G+re/zApVZDx01TrvRibHLiVAZZBRkb0Ess4hnkr35m9dP
9zQWCsHL15AhzyAU/e/LxHEL6UTpRNfbf4WD15wIJfMx4HmLyZ3J5CjDSOLlu33Z7a2TJBDY0YLX
upaGrDNj9c6IIwXNq0Xmi/gbYo0THxf+kVu7OD5BngfzG7wPrlXd7uYJPGcCbpuSVQoaDGDUK8HQ
WWJrq+j5HN0ETmv6EM1ASWDd/ofmE2SmmRQLQ3vwqQTrgrWfp47kedo7t1X1m6JOEVF6I+SUAB47
njjOEHDnV3Sds9Ft8flyW/NvnCaAwEtQE9n6Xxawc1yGq4cYphWTBFi/GmgXYJiXkVdCx0RRzlFI
k/PPFw8e2bbJAPxKknSzOKuyfJnHicEGgWr43WHjVngNo5bVryM5zxFKqVOwbGVCssoiPjcGkvQV
bT88kyl0Jtpzua6zCgZJhwVk5CqZF/0EnTCZaC3kVwu/Lzqpu15nLpLLLKdoGJuyRaL502rwRuHt
xMOcuqxvgkjP2Jb1AkGtNiXa4AhQI5W+ma66BJLJpFxDZ0EnGtiQkNoxaW3I3auO4aXVv7wENYoo
pa6WujrvsvtfKPSF0BDERfd7X1uSnvT2G3FVSC1Q9yuI/g0qcCRfD2Bx7UKM0dQLiHT1dboqK3xX
SkoECXJB2Fg+4oIx0bATIsjgK/4pDN6K2QL3VVfuoie6wNj+OuEZ8SR+/NkCIWYq//g6KoBJggLf
wCKxlhR/SghPsSvPsej9YrcAS54ncHgF2VpIRNMcPU6+bZEHsGJJQXwKQeq31rDNJzzXM+pMRltT
0h9i4YIXiBtL2vyvvuvJqSOiRlKdLhb1V1acPXiYnwL6wLSWDS+ZOhd98cM59AJsVNQx6UooqERI
nG2XC58mm1YmLFzhorOGyfMgreQ7lex74bCRlgj6mbLgqhANEzmEzV2EUAlPiWkt3WtlmbAqll/B
iQP9FxZKPncySNLv4WbVCZEQn1CsXRgyswy3IC1mjayFYcShFZEV593t7AIGTYn39ChED14aC/BU
R1FlflZQDNgfq4SkttAEu++3prQ2ZrKA4Bk4pM5mb9+0RhFbnxmFwonM8KyboRcHPJPakuglL3Xj
iCLJfY0eZNSoy6EslHfAyyNEEnTDvg2/tln8IdUso7njhrC2Nk8on8uhG1mSEI83LYwnbAF4RsHD
/KWFLGIhB+VeTE7L2GySPR1RxqfN3rFPYu5UMfDFxFr4cP1bFKIU3dCjuN8h5flvOv/95kG8UmZw
13CVxaasNcmIl3odO9/NQFw2zZjHtDgQUlA6hXvqIzYXVQwjcAmqZPAslKn+A2/Iae8sG3Z1qogY
o4P1D4Kzfhpq0kBfypEoIDfEoR1nFsUh30iiQZrMjBderK/dgDlcA5Tvp8WYN8z7mR+bUO0RXaqU
VmDuJMXjoMVPtbBsSZYSoO42IEGHVEazH3fdQSvGFPS7FU4C755slcRPOfHvehWp2DOtl2ox/2Pm
zOFehVvJ4Z/uBDg4904PYWJuXUZ37EIqSU0Cum5Xop8F3WI8apIt3glMPHOGNBSzaZ0jDNdj+u5c
n0RSxR7pgItAQXNs+AHej6MRPMJ7nxr3zV6bQJoy/n/8l8k/RdaIZKCrD/1f0yEW0h+6xvB2Vlaj
24hioHXHxXl5SQCQG1QeDxqbb/6Y8zg0gpjVT/zAvmAZ3/v0slENt8pDehBVwrd545JXORavaaRI
AOWFkz2dTttRJADZaNXhRVkFGe+6Xo4G1S+dU+tNxIxT1DMvyrkBJpqb7fdWvHpmD/ii9fIBm+Fu
07WT3sd4ZDdXR/DsM3CCj02TRr3L3SttOmP8a2Mykjrz5UxRM7iqmMdaZ+OdUxBALVRhgQjXftKm
Y87DdxKDrnsw/wiAZDr/WNy/Fkd47mY/zVonY6vUBmA4oyCSPtb59oo3cIlvxxqonB0xcpE2jCVw
VSEwXHrgFCf/GkP4GhI8AJMMK4XHTgnkHWa9JPy0hS+TU5xDw3hw2eCqpHZ8nzbqN0yJZUyxOHaI
s2Z9OF4Xql1yWhHFaTYOgsdGQtle+gUAuEjQ9Xq632mOiJWPNopEH+LQAnIO108uJzq4/Lh0c6y1
yaW/AKbKWf65omQ3O6x2VblHe8oD08sykTm0MsMzlHWpceA3jwhq36WZgj1awoYvJCC+3zDpFTAS
x/3i/gfP4spYomz0rzbLnhJMih0tZHYKzIyIdaZGb1g2DwNNlWNPrk7N5H/FIsV3BfGTHG6tgQc8
Pr+sTbndMK//wjvfaBl+TX+UXQMfrCyc6AJiFmwRMV4Jlq71s0UnSASRfutHaAF1igxMfovYuV9A
PL92Ev9cSBD3F/j6MWvmXuLHsBmslVUsvS1r7iigyQY/vEa/7iIZYKw1pKmceD8tyimQGwyl6w4V
ect1eZSeBpuVBFdQTm+sIAU6AItAByxKJ8Xix+k5MucOl4oYGIm9Psg1K1oCW4ZAoo4a8Bvhnf1e
ciqG5iZRmXC0VX8CYaagQ7XxEQNNSMeebkx+Enyhbh37AWSXAMVGXqRL9Vy9+A1RSbXH56aFIgSK
3DlWjY0Wuc5H2OCcYQ/z5X9GvYevgqV3AJC9HIRY88nnAeLSKGyyiyxyD8lXBdeskl0B8j+uebf3
cG9WjmPnbcUtAtqLOHLuAp6OYbv1tfVfa652kcE5Zy54wrjt6JerqXYyc6NrPcho0AChcwEcsqDx
4MclNoZvT9qSM0V8q2XL7Lrp1/XhVpXI2+eWWL7oTE60ZM7HvoKEcwACg73t8U0NdGIoqm0mrPSj
KeA/oM5lD6Dptc5gRc0iG5seLbkq4T8ci3f+Sl/K3jv/ZJvHqzDR6cWBgAGghNjzfzKilvJnZKmN
6FIOP5PVevWcHnBQktz6S9vFe6E7BWPmTu5/P7BkiSNO/GWD8wP2kRoVjzvRjY5Jrq3Fl9C12A5K
d5UGUtjA4a0WCGnRZIP+ucBys4DNGSVjYn5kbA5bjAiNze7a/pquj2bmQ6YW8hAFebGpEeNpEU9b
l+gtDnNS7UBct84LVaFY3LwRHSR1hfLYgtLn1kcRm6BEvtiEhxcXQF5ulBm2H0D8zNkpUft2DMqE
uDTqINvjtjEYoeYhZs7aGUbb2IiqOK8zUaITKIzUZCLL9+vNfS+DwEceY6isVKuzgyOZWAah1uc4
3fbWW6/l/ruKDTpy6FTUlVWIwc6wxsCmS5s3zNArd674T9tiaxRw+I5Z3t1pDitYysIeDyvP9BDd
4BDgmfIx+AfNBOHKX4hxgSHDVswK1VPwHLds8wRMGIIcnMgRp3jEHdxHLEFfNoWMNKKTMyl/zviD
YN6P14K+Pu1vtrLnOVHmEQ0zosuZcOi4sPzIl0Yg56ieWWsC+eK6EixLWxtbZxKnrwd+lHSffIe/
7SpCGfjmPVbs3g+uBoFZJEEV+w8UtaaObWdFVoTHvbxuM5rhpOdHCpEnDzixcW3JGgrkWkLXqrbQ
SV7ZRI1uUf0Hb7RI7AyVdfc4/3T9CZXvrNpOzrgBgg7d2PDmfRuKGjj2STuyBJgtW5TiIYWVfwkY
Fpn/wrTrXUBU/RFN/wvRjl2S6fxra8cn8m5IIh/+jJltcyN431vUPDSUAULDy2nEm+21LqFwAV6T
tvoKx9ppOUXddFvTJzSIIdWut/p8hash3iTCy6yo16KcmstTuWR307ajWErxNz3meJR6b6ki9IHV
ex7ZoZ+ad7KxHQtNnlz9sHOXosrncjV7MHvKIlFYaACXXcmhJCbyyb8J+XXQDFr/w+Ym5ruwApF+
eoWZeI0ypNLX+cJ4FinlXyWcIHDX6ghG2OP8iDYMJ63lo8wb/irV9Jzphl7g4PMn2mCSLqPECx76
33jOgcg6Ob5/NwRdVR+uLQrGh8WRQFGl/YC2i11cijLeQafCk6nEJ36tbSiUDt2SfvZnyPNTizHT
bkO9NE/MPETLDYQW9eDAzhsTZAuOa/fzWjgQJ4e0rc7vaE1TYaUM8pmmeyTG1Uy153rM0ircQ51m
mpB4tW+pEJ9P1q0J8TzN0U2anAG2FM6u1bFMLLY+TU+zN17Tz5sziCp3gJ63/Nb+BmydlBFUVBJJ
od3ocUs8OFP/CFLiFGtfiqitjijv/rSl0EBtzuHavQ0KNRM1OVq3ilw8dHuj4WUsz6IzXjq99OjS
KBjOVF5vQGJ29UmfrmXysu8Yja/B/h6MZtmKuJDmN4hyY57ItuJmhVy5HcCZrhZb7/yJO67cgXYX
bzFSTosWui+iiWq3y5Qjb7aRHjr+KsNY6eXgudD9TdRP0X28MUy3gDRlYsOTd8/a/IOpryDJMAmd
jbchveiIL9R90EDIhRWnsFqoQhJziWhuxhHYAdmlMvYON2Us0TLa0h3k2IcsyoKupIjllLaRXLgS
gK8KAAgipc5Az+NzSEetPr70ce6VCYGfktte3F1Y0V0aAwLF8/sN0NSftMY0h9aTMMQs15jdOnlt
YX4coE2QNwojpm5ZG6+z/yMnxASUdHnsSBiqWVAii1LwmI/st05tyEAsErBm5njb4wCxTFb7Mnjk
QnZIPz9u9ttPJapvLOhBntFiAPgrYMHMJOk0RTQvnv6W/EYlegGv57xgM52v/Z9fe7nIbzbHiHVV
ffoYikeQdBk3jYxiUy2xoQtRD7kuQA9ocaWMQfn1cIKyW88+fAGPtM02YYL4H0qXcOJ6k/ZS2u7B
3UDsnZ+eFkofuVcin1+gNZ7Meph6cQzRpjWWJxdKbwfVgp9xntTBk6qnGKOullBBWKpoI5u2AEt3
5nIf63dgNhOYY8CkKaRTQ1gxU4+AO9hc/vl8B1ReoqvroIgSEC2idpVL2nWOtjPWzC1VrZ/COsfz
qtuZyET+lPlAhWfh9SggMXKjFu8wQk3+UQKfkm3Vhm6nm0MffMJgLlszo0jMm89Bh0zMt8qB9Z9G
BpisW6dnRjRAkUl+gsbnWUKXHt6yd4XLyaKNmszBCji7bu4oyDRC5VW/Pnv62qFoeUzh2IqZ8oxW
9etzp616NXRZue881XQ0qJrkEMwGAKm9e5Nlyq5IFXfj3VGay09SUMqUg0QQN6C5BDSJDh3hO2v8
j8Tw0xywUj6NueGUOZhqaYc05YKCEmyqCPaxSm9CEfqydA9TqV1H7z+sYdHsOHpCGAeqoMCcNMmu
nU4tGIdeC96MVikfo6o30pQEeOg/6l46XgfZESw7msmSBaGGuQl8nlSDMIoMyN2RRX3UdJxqUry8
Q1m6MEU7GgWIraXHJReVaB/XnsAx/reh/PTMpHwPSBd5wdoqLNSxYCtH0XC8h4YvI6JhvnWNEboc
941l8U/cTx3dMQAd8roPW/+gXe0gLLLa4WCIbAF8/kpJnHhvTRssThJ1wf8mFvJ9edUMjc5PCJVs
JPmiInQ3hjGaWnzoNvkClgsBHWFWl42Xl63KEaK575Hw7JuLrb6KPTUowNMsNGUKDj/NvofvwCvc
1Tn4GbXbkCfKEebtcM3Sh6zTVhxo6p/ZTHt/ihNCpkqMOoY8pDRVDku9zyv63toXyh5Scp/0Zm3e
ywmp4LwjT77HUb+TAD9LyJ4dw7OuU/wg9iX+GmKAZ54AUKRJWmI7onhNYP2bVEFvqPwSc+UdJNQt
a+kZU6Pap0qx1R5diGEOTDHG7iOfxCQBUgYZsTrJEnvdKFBXzUSgWxLmJXNofWAP+eDoZmA586tb
hGNmHbKb9iBm94G+Y8XbVha1vYqk8JSPHrUX/xfutHToAAfOSu3wgrrl0ifo7mtQCq8upu4TOZgE
wzoME1HRJ8yi6GPFUM3XNVEZyD/MT/BVNbGvqUvetElIFooh1MauOv3LWV7L3jXTRRK6iJRh1+NI
yQp42JyyOCzp/raa7iBYnTb0FbGib4CI6KWsZmMR757e0/1P8ZV2dg4M+mkx7TTfH9rEVe0q9ppp
UAUSuN06ETv3u8LdgKhI18i36YFbHwqilDGshprd8OSlqZnr8hceNIDj0fOvSx2qDzU+487xrrCK
GO6gRrE7CmitcR+N+E2geSiCY5AcLVPNvUkaIGIiHmr9a7VcueWdEbHBoW8DWLMrkVJPbk7vPnxv
ynASUh0w2r9Im3eUmHQ+iXN2M+gIfq1hvZikrH+P9bQLix8lBAozjaHp8xnDUTHByrCWX7SZdKSF
jLXHWh/hhpcZnFemLLsWEngmOSPDZm5Q8oufkn/mxzd02tznRMFOLY09z5grhjU7N6T/mcMiMov/
xQqoVyYmdesSPJi5Ah+pkQyisc9p2RLeIUOx6gQNExsUTvvb+fakQWMOBTQP05/4m9evR4KNafmT
qQN6PV3ztli1wXYhgbbPiWUc/A9I48RDdw0Q6l1tV+/6LvLBwUPr7SyLiVpRv7V8xYAyh1T3gs5X
ZvKmKX/kJ85/zQONTlWU35hl5TjUfznePNUOMaCezuJoP7iFk7C3o08iNQ4WJn7sWji+/YzzYA+q
Am+zEPXzMt/MMWWG2rnF/pulWvKujHVesB0geMYjGZ9HbZgpxhpeUDUkct2qsB+/pmRbxduSbLuC
S01yP370A+FfuXQByyoWDfCdgroLhShMHn2i69kDaIQ/l2x4yO1fRCF5++yAhXbhrffB4qKWdKQz
YXZDSR9uruYvrdQpo7P8xaA1HXIt9jd8FT1KAKDY+zgp9riFknnAUB83ehC97oSEbaPCYKWNTeXC
D4E/S0kAP7T+mXV2Vv+R0ICqctmK184x3GwfIk8B+YMAm1QnKEul4TlXeE+pCx5HbE4SG+UHmDr9
xg2GjBUsnE67s7Xe9an7O3/rFJNlby108YU5qW1R8eAda+ir8wqEe94PZmyz1633Ao9GnWbMa/EV
GC9q8BIQU8KkzxMM/ZAJ+jdpYD1fPc+5eFxJw95ghL1H/U036C2g8PGfCTsGsiqJaERSuVLb8IhC
3RNUdi0pmERSrypVaRHKSX83X6/dWLCReITnlXVG3F2JsdMeL+qZ8RqK/48V8NE4Ro/Vq2MZrDxC
uVWhQ7B2u0Jx+En+9mjCuxkE1XOywjhukWZj/g+oKHWw34muFNxG8VwhuXo9EpXCgEYBK6vQGA1I
4ZHMPXn+CV7r5o0gNTqdTV07zN99Q7wQLy/iSYsodRS1NfCKPCb7lY9Z8DSQy/MCww13TAvNMZrY
fiXt4abDIUVn6ltFGm9c1LaDN8m5VSiPl/Ynuczl0FYir/wlxPJ9GsjtZHa/KsVdxgOjoNH9UF2k
AZWQ1DPAhhoFpO4zboZhDOmsYBmK+SWxtGgVMmZrHuzjmDRsKPgaPn4nWa3KdsH9v3KksgCsCh10
xIlToOyWQvAWosGAArjRGbSOvqjssLJn0ABt22glVrwcUCJGhxV1VOSECbYakqkj6qlIopY2K/YH
BAGNpQAGp09sUhRrdcuunQSpV/DiwrPEdm23rC2D599WeNt4jqHjVL0+k8sT8x2M+bcbwq3fh7Ry
AZ+YJNBrFA+d43APIZ4y6AAEFhMMfqoJR28rBqHsqia5S5L4wSUuNc8ZhgG5bpht4RcyKGHedR2a
hpxLP9BW/8DXsKOZ2j4aWWkn1g9Q/c5Rl9f3uHko2ZO6ScTTAbyk9D/vU1OfNNibPXxzseiV0iiz
FOjvrdpZ2onLNxxW8iKnatyUy2ITKRa07+Hmw1RsApmxzSzE5PeNcfY/ojULL8beN1z+JS2t1zhB
8DjYPH4mvhHpcO39KJXcOsKY7eE+N8JXEVF7ZzFMVLQl8F4EEUPnOqZVEEdGPIJknup6f1hJFiww
Y72nHjcGE4uw0M6IwO/I5xvUCFnMVXgKSJOrJbU3G3BMWolIzFWNlYdZ/jraudmUYQ9XwiVrvRcP
Qvo3yEhGlSsvIu966I3UC+7G14Jr7N9besOMX9yY0kdSQy+5YYgbczHUCHyas4zTLFUja5JeDxkM
rwdsfA8NSilI85Pox8pOOuyPSFoayzQI1O+I7NUlxKOHcdhF8cV2t4JEShLr9d3t8jhYp5xIESdX
SyIoE6+zUkJDzNCyEiLgWY8kEDR0mQy9QPv4tuceLdSpGqs9waimS5V/AGKZ2jyoJJTzBDtzX7MK
hVSgskBtjLlKPYEiQZCYG7h+72FL/lvjGL7W8oAuE61WkXAa4CYZQS3i107tHpnBt8R1jpHe/Oyw
3n0V9ixr3zd4UyFepMarbHZm8nOrVzf6q8Ruw9at3W+wT/nbO4F6aaxksJ4gL2q43i7krRa2aDwd
j4Kn07H4zaIGvJUckqV7sB9mUQdcYlEk3MkS7OEGtRX4Fc/n2c5r5ArcFeJ+nc/0SrpqtGqMCNng
pSM+APvcaPhe71kKx79AHn4aWJWmjnIwppo8jcSg5mIJ7s2knLy6LaCN3MaY9UMHAcWZem0wU5dZ
z+m+eK3TUleNu5RTb+JR00eBO4XBdCF4JnbVP5pjcrqZ46UCdQ6r3KeyorUPjttRRq1AWLfQcSfi
/WKPZHdAHVm86NOFVKfRJW8oQjPY+sFzCTyNCHASCy5duahEYCY5jJK5DNKkAZUQKdtg51gp5Ts6
C9yO7Uxj73wriJXMzXoIB5T1sUxn41XB17frvEc2qfmzUNNbbpDkH9FmB9YCRh4WqNe+uRzAMD6/
feRjoeE3Z+qVYQai7we8MSXnFptwzP4WXtEshX0Hgvk7vYysxuOlXJKkj47nXAS3T4HcWS/mToFA
0P5FC8V0TCCnusWkqw9Zq1A6YugHR8QOhi83aA+NFBcwzUIMefP+zER6sXWHoilgVtOPFo6eEd/E
Di1QbkxnpsAd/aFGg5G6j1dh9hwoqa6tn8V4TkdeEUSwm7l+3QwYSeOZETGPxYe9/bYII/p1MkJA
VhvrNCxqIbpRKzT3Xd/DMaNsWAPnd+TjLZWZZdj6RVSHGbc4OPeFKMGSFEd/UbYPl7BipsoAxdzT
bwxeZQYoN8oUp2oApzjT4hkKF6BseU66HjZkZnspDIQgHD9GPVD0gZ6qfkZeVuCQnj2gizYF8i1T
SEohqLpVtkWJznihS8VhGOjjTYdLCDPQxD/hvwd2rBlHMKZZ7ve6hlCYeBCHxTGuRpt+ZXF/nPBU
DtqybIUl7/eFW+ecrCa7BfPItWXl9/3ZQC4+NyqlNIStbjf2gi5Q5a0wlkYdTFjwAgttZFJ5waTq
NlYIFWdqC3qiwFHLt5AelLIgApkipc/lzrqgVif11cxUTpKc0fIJ+guC+JuzXfwDK2pSDrRRDuKX
fRIxCGq6KB0eg8wNaOSqW7CYDVStnK8kvmfV+FVyef7nBE1bwsF+EgVGes/gTtaS8TlUHYO88voZ
Aq9MdIznLHfyEH3yp512PwedwY7E4O8dFGFaWu8NXO4N6QwR81kQyb4LnXMT3ug81+uoQ+2xT7op
CbJs2+FLanbfdYWUSnEdIGkj7yKkRNT3Q1j7Tqv642sTiThr4OhTGjl+g0ywjghesKa7f0nU2N9X
xBn552lj8iXMj6jsFJ1MVaD4bsxIHGY0f/sZ9t55GIJyk52PiIP/eNFrVSu+FXC5ZGL/1o6mTd1y
9YPE6L3h1F+7H8lPo0pGBubpf6VOF35KQSpmY1MgfQ2ALhtmm/NU4sVKANUrhBcK64xX6K3NuOoF
Kq9Gm+ij/ycsRQ+P57uE7EjCZjsOuOSahepGdNVb76KuD70WciEU4w/BlBLvsN8IsYr8OSeRLGc3
4GUFGNjNPwwQTqpwWVCZJmEK9M4PDjC/pKSXW28wyjM9hG+4e87sbA2WWxBmUXu1hTOZIvxla+n2
N+ibhbomepVCaMTj6z7hIGXVm6tiwemNuf55xUgC4cXour4GqBbiSA6gZWyXix25r/KlDakp3LHc
EbLUHmNWnynj15iWSoSqmCvxlI/EyLGct37q/QKbLTjF0lMnES5yLci9E1aCsbrdmgoeip6Sk7W8
WoQzhBjVpIbMNg8t+XBakQ+9PZZp59BpryEN/yjrZU1W6vuB/7vzsAlq1tQOrDlW1tH8/I9kDZ/u
JAmcco+mx6+hV/b25UwhOzMBul9Npw3nfXT9d0Cz3cAMGExlW0gVwZsdgwsZjDt7A8PFoWYL2rwO
9ITCQTBrAtYhCQcEszQvlM0dU1Y5ealj22WOG0u07kABlgtSfqxYz92Lp+iU3GUX5uSZ67N28FRk
14+lPy0mvGa7L5KxfaZYtg1SZLGc8epI+Vy9alSqhgTn6j11GgMxW9Le5wLHRM2xrPJPYnlmRDpI
zeCfxn5cjSC3R1sTl6cIzeHGPW8jHnY2Qn4tZ4kbEVe79u/oGCmAAtUrGU1PQ7IxHQHbIzbXsS6A
GlWoUhVK6zDViKSXJRxpuKQ1CLIPpfB+8j3iDAC0a/fiveJVGBL8jKChutaZ4HSeGy4xMmul12uK
bdpaTDW7sZ6jrakz+OUv9qfHUR4jYNdUnME8Rj38nEYqEJmjbdz6IQ9ztt1cl5Misn9vkaiiKtYF
DylfiQFBOaTetyf8CDT9DfLNXqHGLEH5lg7aim+MHdP0OUehreZHjt9RW+rzltzbMhlMVc4ST8tC
mpuM7mYpsfQkM3kh4PtDnXdrFUN8wlrfdsa57/KdNXR+4oqeF39IPveb6ix5V/AuFI+pCyEyybM6
DM1CEV0GSk83SX8q7ZWOH/rDCo0f5lDaCzDW/mzZlWk/CS+Bpf5aqdpjJSxDPhNLibwB6SwXlbj2
idOmvfzmD8+vOAE2C/zV9zZQg03265EqzyBu2PeqYwE8kF7cRS3PsS0Wv4WHbAKsGEpdQ0qTgSkI
OfNEIjJI0lu/oH0PAWjRSKBe9bRW3ve9BGSKoK3fAEqSfykMSnFsfN3NuIEtVIuaCVa8u/MVbQIH
HfG3Ym5JpU48maNvlyBmAZH36Abs3l6KhCAF5Wnjnjhm3Tdp77grfLr05zcHTsfjlHyDW8vbvpix
IQlKiDUCXAVWSgyLeOrvSQHpF4XCOzyYQU+jLAfOQau0gB8IbypbFT5QSR5NbDMJk9h4GDJifof+
X+3igYiqxbjZrpxzE2eMNVEOqOP+/dIiQZta9keTD4v0eEFRvqnM2h2Yidl/bKxIt9+HtERJwi6I
223I+3aXeA7k/8cFJEyYs0ni+93TNkx/2xALFYjT06DY22BvVfs8Mr4PFljlNZQxTuXZb9OvVbqO
Qo5hdNypcK2dWZxIBWvXUXlfgH3OKykj3z8lSRLLUeKQxvxgNwSYxRU3aPoO/rGIP8N+c8Z1pGZw
pHL/Z8FuZa3RfF2w7Yy1x8MUui8X/fVniiua4+DjhhQ6FPeVX2mB280ckMqpHDeO5Gy6EkXK8W4m
XLfUPIckdheFmMY2nkxfurOTTj041FCVxTuet1AxIfhMlv86hCekc5nq1aPCV0TLe5ML2c3lrxAH
cUr5TLcxFtUGs5rZgVczCAOF1bZQRWmvER/nhIwvpfltIhH62h/+aL4/XDL5g4ZAHSVgmrYATkVV
7PxdLvSox3wXprte1InoIRKOYBJPGxPkncpr932Ax6/obZ7QCBMiJiptBQ/ypQVvYhn2cxJLhah7
esJ+VLTPcOEKO1OmE9hD6YzF6UXr/YAQUlMU8hrVZQeBJC4yfSDJYVDmUF00NDyjX+4uOH5ftFyc
zVaAmKwpdWPWPan1EzqV17L1Adjab3IA0pq/Z7i0KTGDvvl2uuP5VLAzYprO/TZPlCrAIxZqXGxJ
yDpseAixErI4V7cXJJsqH2I8PuoANQj6c7ab2QEbPLcJVsvw+6geadVHiJ2Q5B6bJtB5TwuKBewF
w8mmE4fpcmq++Eao+KAUUGYrQP46vRbJ6o+B07/FZKy9fBDNqGHlpF9J2+2xbAX+0zg0dfy6gm4q
48ryI9biy7N3NMD5o8w/rkp9WtZu6G6bitXezw/PPggr05C3ET9d0ffB89WzSUYI5eakpR6lUupu
mWg8JWH7pYv+XxtkpiPQGiVEsAA1yCHq08QoMQXtyrcjnjHjhBuhK/MwMGWSReds5WJh8oWAaiBy
/TY04ZNm4c/DWCni+lArwWrTkrFOi+bhTbsztUCnWWD/KeMi+wzfmBmFtkWY00Dg+d5/LkDFrTHc
ppqM5uK3xV1CyfPyqHZ0ijIp0DGW+hO6zFC9FQAimh+qNFy1dykMFYR7I6L4wZvNmIBONgvUHRL7
YyFtCSa2B8DBwi21mmOjh9RJCesC5yoZLGsm/lA6cZhPSreMYRHddliHPFKrfnxlL3ilJ5YH/buk
jxomvLdbpYAjdTyhFc0ta+B1mqfzgpHR0w8R8n2Kmu0e8OnwZabY9U6/qjiUGc4XYzuFzsVGesd1
S52J+8VP0eIJH+QnXXsNbsr6VkZqvh25xx5KBGeo1dgwk4DVj85Mt39gZSkImkZqf1g6M9biPn9m
r5QHcP5Kha8TAuh6xfG7TqiCgs57I1UClyzMf/27Q/yAfqbN1AuHzk/ydaQSljadFX9ckvKAiT1l
M+u3Ld74U2k5UVBuy0oEiXM0NETQlVsqWKB0M4D8Yb1Zxmaks49KMCrdNPvrZQ/u4DvvXuF9gdOY
+rYmxlDysMlKv4HC+A/fETMbGHRZ7VaLfT9b67MnhdEGCfPRKd1zRhGnFfQ7fcO8n5hXMgKH/Pyr
EkD3Zr76lE6S4Vznl15N0u1QP3EABriWicZoT3Os2dN4Q4Dr4GFTeCZmkKYZoOOB3TpIpsR2q7jQ
PLiMCS6R9MDTIVLdoK52q6g0sUg2ZV8rUAeMgm4UkZ/6UBe8zUm+CCs5eCYzBB0AV9r9zk6IN5f+
tR7FL4JSH9CmRvR+otXYd0e2+bf4vd86v+SVDDUFUO7gdk24+5f60NSW8wFiu9Ttoao9LtxGQa9v
ak7G8Ne9kTSv2sl0WN4xz0+KjIqYo9G1eZB8B1IOzzQLEvZi9koTU0g+5Dt/Zah/DromjlVOgBnu
WGT6AD4a8SBGiPtwoctsi2Cp414XBvTEn+I4oC621EZbzy4A+AGHSyrADtsO3R3Gum3vT7IxuMq+
r/5DLK/RgzQ7v/Da1o85iU2u1OgsZqa6i7DC252gE1tShWyOz68ZdOtZmhTzDVGuTebWNGaezcRZ
gC6EDOcp1drRmCi/wJk4SYp37q2u27CaLcFGNsuECKklKQY1Z5WrTznWOn+G5d5jwp+NwqyqGPMy
wezKfffD9/R67BDhFdwH9UqezZyBJsXBToLfrH/ZMuvxUP2UYurWSrlTHH0ek7Zwzfmev4kPfjvn
8XMofdB+Orc16oqWOAq9OPsutW12oAdZIBKpJ7uQaIeArjf9CrSntLINoaHYs0cYTS6cGEmf/3e8
iRZhfNkJjhQMM+ZR56q3txiHhpIJZhi+TtiHBGujb0JOPEf6NldpB7RAVIewk2u7nKRPE4Hp/PKP
at0QxxfTXUd8KTg8SK00d/AVqLs3CebAOSbDnLkQYZdeB5yRB3juR2PSuIS/xzC4V7ieN1Rv4C0i
K1r/wtCWdN+qktvoQXi9BnutFS+IJM/+8qwHChpMG7LUanng9O/9rg5bTxx0jwu06BQteRiGVtDF
ygM7LzoekKdVVNYiaxIi4sbgeLo8SPpROE4BZ4KfEVBWILbTPVfnsU0lKift9Xk0ZXWge2RIphFF
3J3cWDQtYWsBzputDHJPQbUgkhMb0QJju1moYplykaTyh00DyeTiPqBj2MWplmsYuB1qCFXYi0ZW
W2euH5Y4aPd73397WULpCBeAALLMMLCsoiUN61DjJ/X0UHM/jHyHFWLJPxl3SuWOI23o1UlQbY7c
OmVn74XR3L3L0JmRb/GyQy6G5he0qA5LXK6YawZxgD4bBqB6PyphYwhH3cs1HBnBQmBJyc+swsgz
Oz4tVNc2l23dddlht+wy6hANRQMsT1GE2lTQJnox1xQUkhXEkcBPgvNboQnPxtxCf7LvzKmX40Om
Cnl7THvvvhnAzwKtt4DZ7W3sewC9hLKhk9U1m8F4PZk3v7qRIn3xZqQzX5M86gPyJAnjKEhFns3A
CpCEarmaeusUY9IgmuviQIsUFolLZFyi483GKHZ9HhBr6TlpuFGMP53bmLT0ytXZ8F4PHqDsNgh5
fOPA1QBYn5WDJTnsMVGagiDYAqYTuf8wYfDTfKvJd76hdDi0CZ5wLAQgDVdna8ywVC0XNJKdPAzO
qORBe2IGil4vyYz731BpaAx7S9GaBAWHg5J9WRNSIUQofboZzocXXTtSma1BDlDfo5k0B8p1vZ3Q
2SpV+TSRi8+AzslLc34EZk5PDRy5ldkWT0i80BsCbD/57JunmLenH+3GVzg9pXuugp2KJR3N9K8g
hdPgVj+t8/O4iFryRP+hM3Bhev86usPr9vog19UeQaZdDkOwO8Jf+x+C3ymgITuXVqwgNSD9qboT
y2/zpzG8Dpw2fuv+jJxk0E4TizGfBnKDjuUuZljZ3ni0Q7z/eJhCSoMZNrmD+Y5vYB80EWxY3lhX
4j5DRIg7u+eFGV52oCTacUY+0X4/W8OkyrKgByKv3H348XhtZVcGJ/VO9t74KwRyzCauMfS1//sO
KiefyLrkQZ5Aqvib3nARHiOfmoPmlVQtFpPyVfIlTSZeZYVaaZzgudGmXQ/++iRnsJYyfwCeAFgh
Ke0O9OP3NJ/IRPOUxdRP5NIr6wBhA8aovLx9hUzz7tzO5xS6P8Abq3Y1pYm08vO+b2QjjdBN34C8
csQzcgIsJN1b0T7tQBztTvjI8gU6r+7gVeZ6BLVSjCFCjV/pmEA4CVioRUpLMbo6Q2Rp8QDsGk2g
fqpWWxJ/OwK4P4U6kJNX936x8pyYtuzliAC3PUIC6OnR1GaVBEFEgM98Nkube0UAK1nwZHi94wzr
gtCegLu3AmFBqKAA82cEqEOV3/RDXVoASQ7IUzG0IDzychd/4zxRJBM0jRBcrU//0gvVNWb0nDMc
ZeTahPKYxMwyYoEw9mFzXY55Tt/zKgaAkHvL00LOH8bgMb9KaOSO1BdPFBoii56M4cPOrF8y5u10
1xYTrHOtSz7cEFw+K++/n87RkmxlFgQw6XEQLt5gkSUCKjj9RFl0uimsooeAWX3BG99++fz6O2V4
/QQt3lxYvH12thc77xbWZwuadsDvL6GCkfFlybm8uZuQpaHPiAw3kAILr0xfY7MoSC3gEDZKsyyf
JJdH9xdhJxKO2SBd2hOYR+UkYa93QWADA3Q/2Up6vs6ilRfYVps60H62qFfMNa/xy4ira3fsUH+E
SEZchEWxOG+WXhx1kp0u2eVi+ksQm4n/M6Wy6iPQ6gDg28aQD4udAAF6ulnnsWzDfe2l0p5AoExO
SmmMGWBKeJFlBtQd/sHYQgzeQG54/WisVAgrv/HI04Lp5AYqIklT8KZcO3ZEEMWq8+NNX5tdL8Nz
Hl8QCG8J//AkWzHkqMxjJKWXtnJi8gAwEuFVhVwj4m+M6FGrD9aXkfa79kbvte/30LQYGK3PUS+6
5fck8lf4JCGTDfgDo/cFWUeOQhLW+VdAeEMmsP3I6ys8Tste7/EOZOovBd7q5tqVvmcN+Yp3L0cU
JMoNWizdHw7Hfd2oIuswruvxVyIGnqngZ+7YNxpRQQePmYXhMZHYHh/APJIrhxQiBZ7H76Tuo6Lt
RmqCWkUIZ4UfX3HKoSkh9Z0e6c+FhIaIvEq1NGExFPLM/pBZyGBgzl3I7XXA5gDCSbYyfXt0pz7P
gAAyaUZJJwXY26VBNYrrqU3pcZWKCUUxh1fdMmsXW5OXmgxN6UJP86D4FHx1LrSxjO+SbfOKU+HE
lEV4AlL+Drsi3G6RLFakoPCh7LFczRld2qtThdodBDFiuGn63ppMTIlCvjuTb6DPFmlJlH01unkl
S5avYurcH76sj0XkrqKVgB8fILyouEa2KOza0UGzjcUsADgjgTBKUMgMq2iYq4ok+nA7Ss0M+ruc
EIWLy9HN/iCj1Kps5P8crivVNAhuQMJXL9OQEE0t83/9znvisyJmrApIeF+9TwDlr3ZYKoRQyq3Q
f3GgLZE8dsVDZZBx9XVDPwTm4E8Ip+6v3ItK6UbSjgZdw6hcQKNQDKxc75Oxxk1s7/YVeL8X2Put
VPYNQDqqjXV4CmhVZjYSRMSEnz28685Tz0Fxi/tl5ooACjdIgkSipyePPxIlUvRsiispIGM+QFp4
pmmKNWS8stcfx0LuxQUwR1SMriNl+47al+B9FR3uZe2LOyXQRWZiKi62GrLifKI+6kK0naCrYyOJ
+vBOJi4T+tdXwJjUbKshIGjkSIF9Qxu82d+QZiQuqE+sVftw7/z/VoUq6RylRCogr0u/9jfkOSb3
zKkE5m0sChFYNwgdkpgaJwrDYEDnAr5MBVJM09WX6DczieQUgBy6KHNza+msNgqhWqOhVUQLDUgY
V6PwSc0Uqn4ZkdE2M/wq1q9+K4QTSuJa25FHNq+9UFWmDCRCbCfkHc3YpveKY5t5prcGe4+oedNp
iKzi302WS59TCqgI0PDSr8Svu3OoE+l54pVj3rw+xTdXQTwGDOHnrICOONFK2rDG5XqtoTe5vEje
3QOnuFmAV5aD7QGrm/fvMRaSHKGTshpDnqHB+NHbBMLdCgkjIFOcPAWegNWSh5bFrmbCo+o+nvyt
29lRQL9IxCbz6evZhtFYqPbMNX8RrkRa8Y0mRj9ptashihHzl/s1mdvX63Am4aULW0vb1hgq8rdS
5bKiWTcPQYzXWtUnortAAd3ILYO1dNoSvrWqhQSu7HDc4neA/rptRts1fpY2fg0P44Tw+zVKZR8g
KecOtL7GFWLkKm+ssb6BtaosR/DDOLgjxDCkzy4mBMFca3nl13gqKQYXc+z7I9613CZhB23/0mYI
q7Hcm7macwndcWoiC+9U5KpKMwv4Dps66ACQaex9qjB6/KnR2Ro8l8J+3FUh3zRcgbdos1cyG48b
DF5X1Xw56CwQhvwPDAkj2hbeAVcZtAMiZgu0dZDiJd0tu5c/74gGCXxeBO8CHB7UBpc2dXXUhh4x
6XoAerj+2SGb+1+h4L72zv5VmF50zNNz1dqeHZd9MFB2nSdebLdETjCz8cxYzS5KL1nHEQQXsVbG
fMd34ZWO8CrITjCqW0W3W2qbqydJ8AZWN16OG/YForDG0sIeDTcJqURvjotzYtFZXBRea3Sv/DA2
+JJ2GO8PK9KoGLsdGfzc3+873Y/x/wB9WlMcPMNx6B1Mgl9C0FS756cLES8HhOLiwlyXzBa8G79e
5p7tmhSI1jhN9vicggRwDnCZA6L5C8nzImVEMeLi5/mXarsh3k7h2FUU/pnKsjehFnQzPo+l4/lz
i9G/dT21god/L1qvYTT1KseejLN3/SidvW+YZ25GTZCofHkrNB7msCncjm0eN6bhVp924u3nyYfP
RP+mZWLLPYliOE9Ymaun1hBNZz7/2WSa9evt3OOg5XsFuuTKxIMUqxr23iFCB/vgMyzjZKDwONI/
yX2LKG809/mb8GvOMt3v8NA7z9ZIBY7BM9lFCIu9Zz0YgQMiXUNEhI7cnAWXMM3QlC0otNFq+uLp
krArOz62Xks0V5Nlu0MU+pjXLz39xkDXkqE+LME3RNJbgGVi3pODKMQAopYjRa9hoFDKumqSXxJZ
xZxx0gl/jmrypIWZuIKDeCWJafVbf430aSOxggqtXkVYe2/iDF5G044VjPd3Vfm0yiRO2WB8DWy0
w28a1C4F2RkPXu0joOamlcHMlpuVUXFa9BxMhbVBQ2KZOE4fIVRuoa94PH51KiOHVPdT6z74leJr
6dvxA+gZpmbrsbck+DJLtOI8hyRLIUfFO1DYvlX/jQRGgjqhuE/iPs6Ij9573UVOgVhL7FMojiWP
GPM2/kOa1pNP4Vhh+ZnPYMzGfDFJTm5cFiC/VfLdnaDCg9mU0RYm+O0tGb+k/V6brNezJpNYmPfl
ZAqT6/yuC+JE2LABCZu6CwQIZWDBDdBEOGHDG1ZQuZdihe7cUqlTcLvoBLpTkHK//kifytOlYgaS
d/WON9ixQQcA45jzayFKoPzCYyEEB/rf5ASQr8Kkr64wuHdVJBEmc/Pbv4n6HdWX35eiKgcpc511
zs6p47jw95oDhcOsWI9x6CT4HQ35aBO2CvOB1269U1CWUwuIno/FmvZj9EjXqQB8GoerQjy39FOw
TKxU7NCVLzih/c7GXA0TBIR2QZ3keDSJLGa9RcZKTolJH0uGT5gRtTmtTWEW5dg1208VMIFZUNou
uFh5Vu8XkBuCQCvge46+uRYDFlDfRyleZA4gal/l0+nef4XUmhbU0maC5qz6vnWWFvcnc47JwMYk
p2odfSdL5eqKRkTor6eklLi1qzj9m0VaYOpeahDNUyblRDfD/njP7T1VmroxWWlE61zR1lwPxvAl
iKUq+5PiRLAHRm0WEtlDowvyYkhxZ+fak7eDkwyIe3BfS+uQXR1GKi7WE0xZDLLWPbJMTQVd6KmI
3lB++/9WPnAeK2LlTIWC14/8Mgyau0QLXAXzypT8PGbdYXcSgU9Y9qa4cYrfXyDNgI+tGnobf5Su
RVbt2fkkqM7bkc+t1rtXqpZD1Ywng6TAQjTFN6xkheR94i99mbBgSpTd8qy9SMqVcUxPfnNjyTDd
FZRXj79+AnDw+95JJeDucT+pJuEmscLTeNd1g6RC+XeTcmNLIFgd7fT35ZvcnS+dzH5Hk56gIuwd
xYV9Sv9MDwbhzQ6u9IC7cDf+xOmFfp86b4C2YNCBuZMmzV9JqGOkb67lt39CBBbFGsu/iYDm8KNX
pXDO3mgj23fkHkB4EoIudY8QizkuJ0j2vZsTjzrrslCqzhrYP78KXtkyZko/od8awQ/ASE0p+0FG
FZt5wbfuOSdJGpXLhwYvHLpmYblIy/hGelxn3722ClAuiN+HPY6//1WfkpoEbX8iba6g0zox1yVY
5Q9KeL3Wl0GxNW9u4uTHK5pO/YAAfDD2K/mzWqNdtOtfDNRxhTOUY/EB5RfTBZ9dafGhiT46YUKC
veW2vVBrHTyhUnHu++qLzbVkR2Tqp0hT7HNSID0yqxZ16Jw234myvrq1/S+QfAPFvCKxyty34A4e
bpIUeI3FPR4X8qNRp3MMRgsQXrKOOVIS8T2VNgwmYU6KlWW5kc7h7NSCMpxe05w160CQkj3kZjDf
MIY+pYOBfJUU0E0JgvNXc/Pi45WBTj9d79Y8e8kdg2cxMSzr2B51tz/Io5JLLEWV3XOTdUuq4K2W
79Q0px1V5/gZ2BxjuRiMCrMvDC+dCNBb3LPMUO/kvGrNMBpl9yNVEQ0aQa5RXnjrK5EHUoRKVMYn
5nweKrhX87JBuItDhCEjm2EOxYrvxWLnK6qkwGNqAT627XMEDJUcO/usSi2ozuT/xLIA2GB3hZZ8
GQ5TtydxKNfBuD5A62bLa1xVasvR2XAS3P4g1mdb5u896pK0eP20AdImLGui2vSqpf7t6PoRfzAR
dMRiNr57kj41TK1vYzssiOrf5t93ZFjl98KUx7UajzHlprWsErDkcb/EDo5FAnVbZ9/5Mr+aXDVD
FMTWwruHSiWeW4B+o8OOpF6vEtil4PJrTeiwhsY1D8qtClE276eBLIkP0P7Vue87ir21l8u/lnan
1yW+7SS6ga4y43IIqKkZy5ubbAGug7skKw8B4Ue5j1atbOouxJr+jw6E5HIOwry4zoYvuurp08NT
tAzOctNQubfoPAuo5/XM5B2ik5zVwv0yOQSikeF2ldG1gUix1lsHn2qCfVQ27hNeNONmJDO51Nkm
K9eqK5no+6LD6GPKkdkXAfdMpDdvXFWr291vYP2Ga+tAYV1g0rdeG79FWuM4lsRVgtOp0JQOcnU6
yjEKtpG5MCTVst7mowBMnO7u7SDVCCMftlcPRXuo8hwnEa2/8WGBv4N1f/vX9M10D4UHObfqwP6f
lx8Z+bvkwdePeJRCUU6WlcfZzomleI/ZTudc6ACukOIb2iFZFyY97qtn8IZbZg2lWW25ugCSQ28/
ur9JjY8YqmcDNJQE21H1xIKJQYStLRmN3vGU1QJqefbTQ9AeQsp5TKZDLy5CWsv9+Bm+4VUj2Fnd
v+eRCXDNyYOY39G4X+kDFtmU2GShHKE4cJ19ai+Kud9cx9J7Mstiq0ZXOIZdLTYEOiM9mnzA1y+1
up8jJRDDy8ZqYdSPex9rvzhRKV6m8qCOeVYB7GLVfZAjmcifKKrnN8xMdTbaHGayBUD2vSJmPwuG
tu59x8VPGMZ8PWm4ESVPUqILwm+aLci+j8KFf7spYoN2G8r70t+zZX7XhepwjSaG1xH1NFjx4KcW
jbBv2dYGeGc16hglROC97QSlT22fXsH1jXnv2PXOD9+Du1i+N7Oai/ev7Jf0ILdBp/so65iLqMXn
BWkuVdlKmxiLCWsE8pWRvXYwiQ5SjSWjeSmXLQwHoOgrrPnhvuk7mW+MLGSlJXJRqBRZ41xrL3z2
0V+J/zOOIGmUvzjJ5CdF2za+ZUzuhOOzsNWroQ1qppDgKoMkWTdsLhiUDg2nehVFZIgv9Ptuo030
1qe4Y/j5R6g40Fk61JjwHKwELsIvgx3e7m6zxB5SEmlVOY9WQRndU8gFGYpJJk763FefrGA3tge0
ZgYCV7N6ps4BJLJdVrF7tNW3coS2MULTuF6ZhAKc4tc7vLxlUyZ6yIfAGDtMRa56dKNjkHCsfzcf
kdfJFqqEb48Fmf30+Demz28idECT7/N4sXrrfOa0V9Fr1OJRvOZM0qFoG0O1kxiwwdM1q+BlNXlZ
fqeYleju54wmEohme3kyVkBhjplZ6VXX/ywzGhA2yQy3mKtMMeaHuwnIeR/nOUXeq60cs6jOBOYy
28gw+FHAvrwPAJLCpIumLelFMydyyfK/lHiKLOC3+qLDDJWJBD4sLu2LmjlUVeibCRcS6TXMpjUb
H5VZ5P0s4AmmN0tDJTFrXtAW5b9q70cbL8OAylsEJLtVgFcbCROQ2GwMYASdWFe9/GvxKQyjbEfp
vrZiR/aTaF43iBx1Q8903q6fFUHVqPeSsTyLLn2kbKpgp43EGl/KFQmrNT+3P0qffKuAz22APdl6
6+Jb7WM2slomIABgYtH3ks113y9JAugWo1AyIMxjAA8uys8jXfVr8oD97Sc7UcBdJovbFy/lq9g3
TO0+T9n9JLwS+GwI6YOzOwolZmDyL8CWsRScVjUlpdzVBFlJweWoZCW4QIGVng8l9vomnlsUl/is
CbJvCfJZTZXg7nx4zjDyUtiOKK4VxAH0Fr/O+7vi1nZY/kIOAK/BbExuSiwr4SKsyExBab/OIKNn
WaVrK2ZAiXqv5TSBWL3dte9OjLtpI/2qYs501xyoI01mzGwUIMJAkhgQjDYfvm9G+4aYxdlH53Ez
j9wxpyqfRacin0WUJr1CjSGGrn4/b3lGX3NiQm6WSac1SqgIYndSve/K5xgkIqUz3GMktfnzNoog
Fn+MJTtirg22r1p/+36bSWlsVG0fUuoTlkJyyjr0LK6/y/IgtHSmx2rv6kuX8SQ1Q4gAp0fUF3Zf
ff5moolq8BZEqCk+e7vjyMhlwrgZ/9m6LWZKumZYh0+lsRqyv7UQp5kOZyFaIZ3PCqBKVOWmCm/m
4aMiABD5aXFw8j/NfShv34rGHLsKzMhz3lbucYcEZus4hBO8HRL/+gs92geM95IKbh0PmbQ1R+yG
euj9F4/7SjADvV3mCgWl/fSCGApMBLF0R1dD1e1JILpWxL0oQi8WjZrp5roCPOYA6E0oK+LxtGi+
qVuvgBfzRA/8hwwg/KtkNeV/UsOa6zs0I6D/jA/EGvgnifWMGqQ+Ue5B7z31XlKcwt0upc9v+ouN
jY0sTTjpbmyXdqC+GDjfyvBtfg4uAsPknZGQkzIxjV2yKCKsxTzbIBOqa39cgERZ9viSSqLB5Nnv
uxsd3cXfMhyqQ3ufpPbyGl5cOn1x6YPitnLoWYIqkG1O1oIvZvmNiPS7IQVVLkqzcARHHrTThZBo
bTgnqQsJh0c/mS8dVjcirGvChJ880vbrcZBFiH4pOH9T0n/MNYC0l1scmYAYSA+9q4cu5KYQOdXI
37OkWKwXPQOXgBYBH0iwkGY1HoJ+iKNFl8Ppi9vZ10IIk/Mc4hdmk9tu45G7YGZPWw4Io2HZmc3I
FTkTIk4TtZnW+Fuu1w3tJdWIQy1IuLi8yTR1t8w68R1408HZOEaCJXhaF4eJ+O0elDx/IUibUekq
NXEhyQqQx3sD9kSggtHb0Mmrhn0lst+eE+/NHZXYQNUXESr/lbb0CIfzVt/FjtsBKDKSgPOJ4xtE
bFzqVXhF1IL1EjkTYEYkSHiIFbzzK7M8uK4x0HqH8iH4+sq8cAtTHEbak9A0JECKasxPiqhv0M22
PJZ6yODW59OmakYpmirp1d77dnxlmrr66SzLikDy0/VP/wyXrTQPTKJWHJ38elvw/bcImQjxlPkK
5WtzrjNbM2LZEwF48DJkuETaXvIomJypAEMtJ2ZOR91Ce4ZDNopTTy2ggMElVDrMjs8aRM7EGL96
/CbewZEgy5KDGJNj7chpJ19gBeKBt6c1LwlXUEYiO3GAptsVe+1k3UIyB3RRTwg4X4w74XOMFWZj
Pnso4cs5DI00t67G7qweG4vkYpj6UjIM0/BtSymVKB9YnLmCAL4peNieE5HyC21Hs9JB5U7H3F8U
577uep8ksNNyEYXdHOFtJLQJ8Y3y48ZLX2+yMHyYljqzyVO0KQIBkWOUqkJHWDw+hJOCL4+xzRpr
ggptojN2I3cOczWP5T9P8pC1bG6xhhQeJXQVOjZlbjE+C5uhS7nQ7aNWqkO32vN6317y+3CpDtIJ
mXTOoDPi67dxmrBNgkmw3pdQHxj09FocpawMzKnM89b1tUFzM+UwAwguW3ZoTouT/Nss36dgIO9s
20Z80EcRpdtPTmerBBDBSO1IFEeWzC2OjIfPtn33LIB7gmFP5D+czf/wPlPWwZGSlvvOc4UdQbja
ohWCGCH4P1ml2VP9Lf900wUkH1Xx8CQUbifHfsAWOPtMmZe5/hZvTwvjhvT1RN6YcFt8XA2iXiHj
Pzj93pTymqWdMBIt9VRaELmdxISf5Ek9JSVx7WiJtTzAO6g4/RTRfKNb41+1vX8CP7ZiEH+fVZmC
9wt7htJhByvQMA9atMRqv/7b2049NrTxtATs5dQPZWXD8D00dYBhZtIxUZUs0BmMYoCURrWFsYzd
I3yMJXAgtoNmy2N1jPGsXuWZ3F8oRYyw2SEdpTYS4Ukwu+ZvKsfxNW2cAqoA/Td2afE9LJp1I5DO
ONbySN/+IuuRyzKBUrlABiCcFPWCQk0vIP7+gu607Jz8cBhmCfD/MZGOjMS4hahLFHcu8fFBU9Xc
oOegWvFdHMeW3WBm8xwoGf9Sxs8us8Bht3Oz98VGFnC8vSeVQZ+JZJpiXMGtcF6mSaFJe/oQQhPt
+VnaFyMrLPrOvIZpzRjaGb1y/RkgpHPZ5qBkYqHY5SEWqREtb6j1FW064A/FAcQh60KJJFHtiVGU
VdyduM4b9fJ8lUN4hP0KpmU9/nYGl4IVsb9dJwIKIugfwYgWL27ffWSD6ti+Sk4nj9ZaGpvzbmwp
r1tYA9y2pyf1D5CExFTM5yrVmw2dJuU0UltdjkDrQrBDYFFuLxvYk+G5bW4/vOxH4g/wgrhhlkw5
JCj0ejoTxjtCw/X7LS+Y57FC6NZ/o+hF6frq/cj/wC6H9/Q3XVyZnIviXcc5Ge75KsQ4adPBdDn4
UlsEddl2ZnhmDO/6gTVDas531I9Yl2ZpA+Zn1G4CSQP8Mclvd3ueVKMHnbKBZX/uXQJ8gplOJ+60
jwXMr9pg6Pgl1ja4zUxFlJdFz7liA5C3e6SKbWqMCp3Z5Dy7xe6zpc/9i7WuJIvEhNA9m3kOQYVb
DEBUJv7cEGrHGz/56okEJZ7lHFpQQaGjB0wOJ582el7SrhWXlC14vqzOOvR3httlkuWecfQXi9A9
4cy9+DUpC9aq08+vZgWpQyaFIj2gIn2guebE3iJfJVG5uh8eE+e6wJLtoxnJR1io/vKdKQ2Eo1Ko
drrsKWk/+TVhVmoZarAeoFW1c0VGxj8zTyhG5Zn2WiQU0RpsXK536LJ5R6aO7vcuvRDaDZr4YOnd
4b8Vc+b7gYepGNeT4qCPwiAYZX0tPQg0noT2X1x7fU8i1dJe01hkPOdOpzCmkV5b3PjBIx6uYBuv
XKj3BHuENLbrcdC73n70PiV86ax/GetDPDpGe/6LssVHW3rmULpmaviutyi99Ci5g66SPRLbhlgG
fCKUuhtRfksC/r1A9Q96Pv1eL5MRFfDnbo1bn1F+O3EP9PEw+/VTdwwqMt2rU0Ov+91UXDzPthdg
ihTOCNgfFxjS1rtXm5k86NHw+aFYgZ6znde7YzYje3r5PZNXVaBuqLMAa6HLiAjjc44Y5Iz9vkce
CVqAj4S0c9JZ8iwygUmKHinATIJ/7NCQAsMbVD12u/Gq3BZ0EjT6InQ1q1FdqjD/DLo+wWdC3YUJ
8BCjE7Z3BiVRRjwfd8Tv6nhgC8WlDfBhzfut2/Y3Zhzjeuu5Ak/KypZoZwH5dF6HWqMkzyqOOLA4
9r426LJeZt1uT8fNPcSKP/kgoyN0c6lMjpKcuuAPPwZj0f+uIB7mxcP1RdWKM5pLaQ0kMTlsJ2Wc
X3lraurP0YKbLA5q86usk2Y5AErx9O6/b3v6BLQHJAtZygIlMwFp1J4ECI9LuDH3cOmFGEyb6agv
wKR+jkz00DkhfU4lg7HpvsTR5NGGR/NeuvtuYu+xEL0VdmlRDuolHgJKbBz3EKBWJLECPEd4U7pU
i9gv7WAWn5+C5jAW1VYeIMuqAcpbuJGn28Zmm0WseMBoROzc5LEhpRB/mwATmHZRPMU9UOwrPknR
n5c3ZVpqCgK8weF1+dyT7IPz4ByWisVFh0wzEYHeBvjS82WsHfOhYaWBBHfTQictM1ZWY/QARzKW
eRx3FmfIXD93OBgu2/baUKYSmQaFpA1mbygdQk5oX9T2xpo5me9P+YGLgojWIfrW/2xwYaEdGLpk
nIk39Sqqb60cCP2+xHZJHW7X8+dkq9TzOVlr8Tqdww52HN2P9nCiJoq6tZg5zBEEw3kWsj5blNhH
r60wwhRx/P4PKD1feGzFaOwr9GYhG6D5XiDdEAunLHvo50cxEbTtjCZAwz5uSCGoxCgPJQBrHqcY
cDDfizlD9rXlVYjO6RFd6fPWYXWv38/GTCD1RQ83leleWh/EU/GE60OYEaIc7ym1y/US7s0x/9cS
qL3dxKcc3woOmkctmLoBHg/s29OCAbqjPslD0/I2vC2Z65Xv335w7/ss6OLUiqw+vAlcOXQisDb9
kdX2phBC740FZ7X2Hdvr/B8NN+N9CAgAGxYpdaRDP7iSHO9X1F1nmStsw3nCHsmWUaRsKPu0MBxv
K7N4XbDCs2tGdelWBuHKfeUMpWHkn1WzuQvKwstf6OU6ufbnu5FK1XAI4KHTDepzPfwVVtFl+I51
dQ+w2HSEDBuHEHultK7IX6Ot5f6Qsb/1+jbYSETttMxuCuP8/rRdBh1suv2Inx04M6MZQa0XEfeD
GpMKiVRkH1+HqHeqhEBKrmywqH7XThQItooL5L7xa9GBRJVozpnuvD+KTEoibbIJVx6s32Z1b7s/
7nE21wIuxg1+72p5CpGoGXig3CYT1oJ2N8fyKiGQfPFscPDHnH0RHQGbeDjWlPzVLFIRR0i2Aubs
1drYf1lRrCrG62PB0E+Kcw+YVkfaUVqQBGtOnCr2DSuZjB5WVpjkVtJ9FpzA/Af7exqaF9yb6/RX
KmHu+db05VgZquxHmy9cgL2Frzcp7RAwN0vuJjbO/lacMtVDsyZbNh1E95EkzhVnnXxXYI/73Usb
wF2UTWSN1H6ne+tU7lfHtQD8So/0KJR+POHKIlIXiANIKm2eX+UUg4HSOkNzN3oLkaOs93lydgBZ
zgl+F9G2YVzbX7nHNnDkhWIgOP1l9Zgu1F+dTHxSVtc6e2mBe8oFnhwSdtEii0HVSgb3E+L0ioQ1
XYuLWS079RFHjXYGAISIYD4OAKIRx1kcuTweymticj5Si1jApg2saVzQ1cC+fleiaLHbMzTYf5gu
dGUe2B07lV+qHJ8J1NKjZfHxqSTfKgiqHYvvyoR09XvwOuxfLH2b6vHgIKYHmsLueEW4L1nUk8Pc
VefMFmw2apffj154GrGDhPMjzcDwArTjy4u2RZXzT/kqsHthvhnZumyF4/Z7CKZgLXhY9/zaEDTx
OEPf1lWu8Y1BdhPkyjvkDH9ELvrS6Hv8TEWNWPFgQG6qroM/mfpdFOQxmpT/eYxgnTt4+FyxvgtV
jd4DnC0W4lpyDbk0fdNhpLjt+Pz8/n4hacbH2sqVoLCgMnXGsPb3t96byPLqowe26t3QHQ7p6y+g
6wJdqB/E+CIShSLrBJ4e2zgYIow+6Cw/5B5b6YwdbX5DtjM2YCbeCMhuM0qsH6Rtb3XSUK757INV
lEdl3yTwdgYV08NP/gBN2AlpaAgWzeCDpixnBaRNSwUDgHIRuCqC+bzg0LUI1Zo8hnqjpcvM8k6u
xBoBeikXyBJkN7Dkjgdr+FFIimnNOIA5LbG55jq8xeb9XmjdU52s2NVx68vA6X4RvMtENAfX3OQp
eGHcQxfLdb//V/E1gTxpVJNub5TkoJewlXquTy8JSgIFemgRwEPnW/kMdzIgARFS+azHXTZHUq+8
4gXvH7e8t2dSbbQ0g7UG6ekQhlSbWLxhCW8Mifo4GjxQBKGYMQCmV9jbLPoV0voBnby/d7Q1lNjd
L8CcBlVEQE9EdCpzfD/kEi7T7j4tExT+peP08uw/1xvpjx7PZhSjSXeBdvhGGXWCuDxuz63dVJBP
8UOiePSZE+gpvR6WCYV6Bof3nTQjNJro8P6JldM9eSNuv6V6keju4DJmi6R3cjXXB2gWDh8nqW2m
+WNrxKoTfFl4tmkVB2jfoADa6mTIv8pChPHUEHS+fj5Y6cZq40a6K/G9wb5dnbZr7EoRY5Nkzc2e
XX/5b63RVQCBxqB1ZHZ6PeZAHb8Ru8geFaZ9nkpNq1z+/J0NnPWOQ/a1wQ2hsBxnvrxR3a/qT0D4
EkbGzKa5obxCnvvsKfJVmkQ0aikJyzgQIM3sSW27o5F6pigjb9p+ycyVpcz5KHohUaDtyIvV4ehx
Rix7Nxf0wUhn0prP2YVqqHADDqXopbv2Urw2rN1Afi5ZdewwtNmp/8mUufF1CP4J7YyTMAp1J1e4
GeL4JagrONiqpaWM/ckEQca8oYqRdRAakbxPIFBNXSGrRcJ/OiRBfo6OzT0h72y5KZXx9HPV+5F4
HAjzk13A9NSpCyR/llQvmgoxXN/hZXwLR8l0km0Rh55eGzV8sphFhDJ6aMgAEp2e2DC5znaLva47
nDXva0juVhyvXrsE2S8B/Ok9iSyUwaO8ScRf7zI9G25k64ohpIXTmjv9SDW3FG7MB+qd+gFINT/3
Xsk9GQLZNPjL1S2RZ6GJw/LnLtQphQok8K/ajmF7awsmyUmAWRi55JmH4A7GW4JOPsxxp+twAvJ+
73UR40h7YLTgp9rDyRGMXfyXwD/DbGOFipvuf4d3wYpSFx3s+P0oeaSfezfPjgnUreafxSBCi0fT
s+8XXxn2+hoNXDqrar0bO/oDvTLQPLnSXmr8qwYMkVSVNHXerewZyEP8LG9/pH4Sh3WcBFEAKNJy
f8ugvNbsWyhDR5Z3m9DmaoY9D1Vkc4DgovDqSNggK9qWbIX5FIohGtnzLYbANh80HwP/Uypk8D8x
XYHG2NhWuC/dlHuMZVAnu9xYNnKHL+TjQ9JkmDvm2fV50XgyP+PsIcJS+ZMzxTz3lL/tOHL1nT84
YGAPUorAqaiVbMirgzW/AoPBwmmY7SV5ILiFkR2TtGxiB17Z8CwSXh8qx0/PD0GjDc9fswHOi76u
qvKXc7cbGHUZZTJTXsiwiAIAdTVBwPg/tRWIDa1ehI13JVialbG+v9nQp7KFhOf66MAbLTBT3ME9
iOfqEHygkAZBzp7119jpB4GmVQ3FaoGnxoIOeS/YfqfiS5cYxc2Vn561+tQ4F1VzIBGQsznNFyb8
5z3bz4o+D6RPP3UkoNTWrtOxQgcQKnbr3z1P/EmlrVHMq9Mn6zfqmCN1raoWEUDNKtuGXy7pgf3g
NBnaQSfXjLZc0nblFLuFTbOybnw6a29jXKOhQ4JaMLCQ2lYvk4ALORlXJVFMJvikdMkiOWAM6qVC
kV0+TtLOTWHtRP5M/cSpTNC45mL7TGCzJNiP1w9xrAqXpc0C4AdG61DdEjstQfJGHMq/1qlzOd7u
UQYmzb6aOILNg12TFVxelbwnzJqlTy+ldNKQcITrtJIkQjTLZ0bIfgSrVe1s4zfPqgOLs/t6uBTS
F9sfrARZT8jG+YJSxIO0Tepgo5gzaBvMOJIMAUNJnbwT9CVVn0H59g4SW55oBeMm/papmv3PaEZ1
coxHv8QgieXYeihzbeV6vWG7E3PmTpfJLab4VLqVBe9yZnixlmIYPZ+fZZ0iZXOWkuv6lq4T/hHs
dXCBmMzI3sZs9oCY94+1YeSeEeyPQ7vMiGKC1DQlCtn1plfarYbYuhiIunILi77cpN7ucg0/YkfJ
Kclw9NXQ62E+TwHdsJDa7HxDVqcz5/nUCUl5vE6eIhYQEOW8bMn8SvQE+ynk6Tb8/VoSwFZYHOvw
vpHY60G+2VYyGftI+Exda+RXhdkxQvL90kFHTS9ZfTfmHuC126EleA82jhIE2BVXutO2RNPClfOe
6Li3JTwJuNrQbgabUgLToHxHEKgAw0XXxhso7mBicbybWA2l03ln2uanGZJX38c/AwS5r8YCcqig
qcTbiwXQ9w6lRrx/pdlNjJneURNllZsrAB0hMb/JXgFt+M1IuhOfel5MwRLeB7PB+F/2fexRfmdz
tFRzzZzHfuXVTWh0PLhcEIkapAfT07mm4Qb5sljNGvIpCtasSZ5xes/CVKBM3EBNx3frW1T6GAzl
RvOwOziISyhcawXo23irYhnQ1ZQ2nnJY/AMybeNhvEjWV/5vLxkwgLBnQkh8jiLD1HP1LRhyt1u5
9mO9wITs6WAaQ5E49wOFcFiGvQaL0Qj/XRUSPyNGzM0RK5lky4KAk0FDI8SMi0AaGWPDa0j9AvLv
Fyp3gdLpHTU7iAWNPGC0Vic5Iq/L7iTbhuxr8P8YM3vq0CCh52ZsMnHOhpHstfAYMlJp84thzhXc
RXexqW+eMQ7FoTMUjaR3AFiE74TPARpp6uUe1/m3N4ZW3jLqBJZrV9JkWptqVbOO1Ms3nGuj59GM
7kj1FeqWYRgDwsFQ8I7yWitglH9I/eK2f1IBW+CRgMA+99yz9CtUI847WaXCru0pDpE+Os+2Wyxk
S5DMkoQ7SY2gS2eSfJ/KJNJUN3mEj25Cmf6N0RXL89SJwm0weo2tKuoczBg/M9ZBtZzMu/rj8HJU
Qj3PDcwvNpZo+YdqRgLrEUyvfga4JpzBXCTpCRByKu1SpeO9PfBR+SPfBKCsCCfoIEResLxBb4tZ
TgX49ObFHsCh/n2IAv1v+EpibGh0DanaHIeV2W8SD+2yWKmT3UKd0HctIur5kcsUZxIdV5qYBP8/
3eUKMBSVs3IehNhwDKroY6kRDQGffYY3L1Ebp7wFXiaTQCHv6bZl8/gDvJgGbAimrDlRZ/A+N2vg
aEW5JGgMtyG1CPNfSdC+dZqPozTeUpqkMvRuvv3oYAk3BBVxd68SOB66b7BmEhppBKSBQw5TydiM
G9XvpSG2j/9DwvZLBm8/sjMEIHGxAruUIVfgez9gc5WfHFC95Y/uih8o2C4FOi8MOuWLcZEgdZD/
VIFb1KsRhl2YTafwbpfjKNf1EKa1gTbyeFDSi/RtCw7skr1MhWWzsgzFV6nZuGzbm9wuLuZw268K
K9jtWNpsehmA7vMIqcbNRfFHOhxd7GG2ml9eNQ2uMTJPH68vWYrYMRgguTs4LtarxL5iTVUb7UOL
hrAP1fbRLGnjgCMdH3n+f3r1Kn3Gsfw88fLLf+rVAbGhQFaDUOYzJl63BUIblNAP+RbpkkLaiLRq
msJN/Mv5Iqr+/HnIeQsiPxgiyzDzO9Nhw6F+cOftDIBTxJslQkf+Kj5kp621s9OZg318bKL/9Hbo
MKKvhCZcKRcbUad/TX7eNY0+Rky9wV2FuhEMY5uTzLWXmx8Lo0kY0ly9pJDIB2svOeGbVwUGhPvw
XKn8ME9AYAWEKe+uE7jrSy4snsEAJJsRzFVz0evtAzWlVN18BYzgs7G/BcuEmFkJPd2Eqy098RWt
JLJyZ/vkt2NmAf8NdmeJCQvXMhrHCdR8OAUlGMa6vV6BDmMGHDxKUxqR2wIJhANUO33XVz865c4v
GXsvYTd8nCwuEcfT3t6XWSNgR5nS+kYtVIZYLdrkyL0q24oUHKCm1OH1/o/ToiqnYXFdvl0Ui0OP
130uNZkHFzg6zj9GuQdewfJ/wnVIA0Hc6N8D99Usi+l+U1kVP0JvpzE0yKhL0zvYdySfeGx2Qcul
5j9rAHm7RfFIYcX1jjb0ZFyMQLQAapMXr4XrzMCUTjMfOpngkOSiZ3TUrMRE8biAeLR3GzBL2toT
rzBRbMTTvwgqdYOl503EqXQVb9LM6ca9YoMZop2D/iZgn+uHWsQ+j58XjnIy4xEvX4Q/zbMqks90
/5Mpl43+go3lIailwWsiI/wneg4RdQoFYG2FAb5wa93BCO5LZJYdhUUiJq/4zJZStVcpyd4IrdTH
GMKqRBOc7ftXCjvLHPVtgFhkT+ckY2PwmEa0+KQDIlFcEhn213ZTS2LOrFXe/LwTjS5kaqEiB+Gi
VHp18QKjsrEGt3fpx2bR1GyYObnv9OuRx6znUX3ZdX96GRRmoxXPltvCAHVn9N/FZOV5QRpGXtHK
/05Ba2a/Nz9qY50vgvT4bL4NgOxsSBAhKVy9gEFxCxE7JKU7WRum5nWlv49ePwShtId6rkMcP6dK
/KSjY8VZQYOBP+uTSyRApeRAODOVN8sRZed8xsTtD/c88F6FKpZjsSSTheagPm9wz0r59/hRs9Nd
fWHdLCKoI9BArtAK2oqehdqSZXqhNBNKjN9IyxMG4qWwF9nubCmkaQ+IUoSfhMNbibPJZNBzqB8+
JTc3iyU9wsXsAlTKKerea9VuEqzj5ulTrMH86k+KzTmJZuFrUDvGIUeuZV3bbxLQSmTGARcBpsPp
MfJfXfg0K7vLedS0C73j20f/xGKgjRjhDTpUNS8OhL5GGFqdA57O/I+D1/X6ih0fyqQBCZE/Gu72
wZfz+8kENrC5B1odzk45cRzOWyEo9egxb4FDy/lZH/v9D337HkiLfI9z1anE6MrwlczB30BhyVLe
AP6tg0gXCihpzvWAVUde28WXgPs87lhE4H6yi82mJZV8Oq8Ro4pOJuJN8Aw6PHEEj22u2BEUid3b
THe9o1/xVUQxpsw0aPc4YIMHfeE4oDPtq3sjb/H5q0yg9c0GECsXRXiXztZ6BwSwuWcLh0tbEiXM
ZkoURRXjUAZUKwPviweH8eslVAiuMtSUjTp5Sry97yFjuM953BeaKqJWbUEYhBHBU365vDmlYfn/
57Sn0Lj2Vd/Fef2Afy2VOk/lSlLOdV69SZTCneQJld/LYLqA72b2WzvwQwW8GXvHCTzRqEsLZXk9
jSLKV95ev36PRU1ye7+OLYymTQrc8ysG39Au6JszCU3FXJF4QfC3jVzWJZIZaCBlDy+FHcZeyM/3
qDipb122CmYXLBG/boxUds0AftXk2iHPTaxhRdKMETxDspm24ah/3d2hOwIb3ahsW1Su150DK2EC
ww4YS3/Qpwpi8gQ9kvWcSrf7N92r2vYYHsM3F/HNEVe2w7d9rcKIJRCJbQS2AJZb5Gp95X7WKL7d
irs1Yya3lFzUpX2FHK3P/TVcNW0QtctzH864S8LRRVo3mWeD3hgRF94jtAagJc8lr7qbKzYAxHvE
W/FVR0La/RclJ2EyAQgAdmX7ntyq1V7QIYWVbrVQRB5/1uIrjbOC80u0jRwy7uxM9xS+RBWWGlsU
T5pcB2ME+KMkG26RFWxSTLgykUcnnS0rF68NqenQoKzAYYd/zPjCjmfD4/5A3WTaoErRBhq4/5Fa
o63e+WyxhN1SE/g5bOE/UWyjcijM9bXZJ1i9kE8jyNf5wLkIynbBJaGZ8DUPQnrVVfbkyDyc1ikj
5a2UZr6DYeEE41qlnQz94OHUidNLl1s/m8Tny/EDJSKxlFvsz2PnkSnC97Tk78arG6NA7Z2sByAT
Nisqo92ui1VHeUQotkGyvYgk/ceVJOkkX749B83bQBFYfmVYZXFUFnp2wFvyNMJ74gkatmgq9S5z
hSuHSbCeHkT7ndUan1un1/ktZs/5KAnAcTcjjOoZ8sTid4rLoyAtzF+q547TI3gwD/CjiR0XKjyq
ZB0etlG8e9x7lz+1IEh72pWAMKwS2MHA/hPGwMX67kJ+KNShLmnU2EFT/DsbO9j4/WDj4zwa6pnX
L2YwrWwlSV4s/x4HsswQdJ1nV7OG/koYWuJpE9mTaR6IpF66NhifqZIwx55tbqeordHS+el7cKR2
xgsTxQQkIqxRPYrpdkKUwGZmOkL+2H9ePuN+rV85HBljtwzQcVrCJYcG7CKdyvhvepXktb2wdKzB
gC21B78oJ/PS5nZlNVnLuymj74jIMj6cMbJVrYzigtRjUxBYCaJPhpb1qzOh6rb3dotyO9PxBwQF
3bXDv8gCaEmNjlTUwM5M0vAN1lH7P439xo20mWoa/2jHkghiO0k14O6bMXLynnb/YPUTzhnmmTo1
Rvdm2VvfPoQjNevcagE+B9/dv6OU2YJjIwQ4o8TzvHwZekkI0A0fakVQRZbhffNRrzsMp5pJEB6w
m5/FXllh50/M5dOLfUaGcX8mlbmPUzAGC0gwQOeAA+CTxHemj1W4+Qb2Q7q4UsdATIdcxuu8MDZJ
77Q6+y83eY9igooSaImmxzYkuHV8546jF7cJMSXw9w6qpAiuMCPJQBIByRhw9yeesxARCyj8r6vp
ArliMdJWLKfSf1Q0F1YI0UaiyImaHpmzetnPh7nM0Dtxna0GcdzY2crtHitu65s8neSaUNPyh0ja
jBIy63LMJQkMM92WAT4NN5Sy0vAPh092ceg+lo6AKpjhKexVssYLDjkLC/Q52TZT0mHQwgb73a/q
KdVgo7J4xPCbmYEGL3FYlllAx3adsa0UXrrUGHQZZUpRWOCRME/+L92nfAOZwI0DwZ2RUeKkU67m
mCTqGMvSK388C4ZIy1VCj6LXEEDWQcWeS+B5408kIrRfoBBpVBt6KCx/LQJ29CFciQnHgVfVcgSh
BxxZWQ4/1OEBy2DgUVB8OdS1nKBM7zh3cmoJYoya3aFweyWf95xTIgLG1vPt3lQqc7W7SbndhWPg
obnpKpBbvUqaPN33xrIva7wYVzt7+s3Z4iM6zwEVtr8GZIUL22Eqhr0OipVvSisSsDdD3emj+0Eg
YEjHQfPRyVJVss/F0faxYkN3cjtcq42WlToul+SigQrVeE2RMLX6LElQa0XVctR3wZ7ag//3FxF+
V5EtoWNJ18BKXvwWh6QViK0zZbL8MFowrH5yJ9ikLCyjCwaaFcaGkzNTpRnicwqqS9FAR/HDwK4K
yR5KDnjAvqe++ZpjyqnwFoSP7ilPz4eS/A7igI+bcDhLEnAWtQ9Kpmcf8cSY8rY3/Bckgf7ocyL6
3lwBceGqHpt67cm5vqbmKnMmIeQPk4QCcusD/lIKpV95XeoD+AsbrmkP8ZiWX12/13PJjRQZ0E4A
cEdXKzkCAhvEYAS/5yo73cxxFaSf5UnYFnWTDUlRxdXEkufILbsKLgDY8Y38FeGgysFXwcUlhlS2
a1SczBmWHmkKYTQjuRYHGhaaAeFoOgCQUKc540ytTgzH/BQPk3cNLchVOltul0lnCbNxabD/44FH
DfLptkbg+EG9J7YjQWrWN8zUOcr3e86AuQr9Elv/cCV96itFVBzvQcXHrXpg9BxF7zUF1A6wIaV8
vFFrRLO5/96ClYwwPWMOTglPolkEXm63WlpJXfiyaD72zsWlcH9kN/vDv3sIBGwgi+LKjuTE9zA0
E9LsFtoE+FKC0K+aAxtjfjb0GiblU/F7cAl+QjvsN/bqVUCBMI9UrcYMdgk2wQGoGLb1dA3dXtSS
YpYycVCl270+24B3JvWov+/f+7muPBLbZy19/JdDYzPOvT+8RB+hAFr25L4gN8syqAN18pY4XPhd
YYjx/LHtdQ8E2N4o5KMmlRXjXv3EcRsSrLWtAjSVAuNx2JyscwVxqQz89tjE+jhxmvKLsO6W/3YE
7LrnddMN9gt4sK2aAeAqCN6ORbWft3AAbmhOViAGfpejue58kd32lmevi1GwNJ/kM11KsqU8Zhh4
g0IZ9efgRMjJqgB221GOiYK4FGtkidcgdWFzqfW4cCRGWqgKsdkRbuMuKbRJESfl7ycQNpbrsasj
kmBZM6sqgBYA60Z1f30jTptRfQOuoRYiUD6dGCJl8O97ZepFjKzh408xW5QNVAOgYAznoY0/q8Ss
XM9gHsw7apVHWwp6Bm6J8XljxYZvTX7J9Sj+EcIFsHRyQH8qpV1Be5eHGLEr23OXd75c+5LbQe+p
fQpPsTL4X23f5NtYcBORtMmDCAdX3aEGN2QvhC1CHVYF+FGLRTBdV2KXN4aHa1KBE4Y8pAOJZtya
DhMLfK6N8UoazEcm0ZN5i/zongXA1Gz+almJSUIotDnzdX0fxDmyeCk1OeSpvJOMOv4N71vIVA7E
4y5j/PW8nFuyiLP7jyt/chJaYjjB7sMXjb/jMi16oGkfdiVXrlT580hTTt4k+kG+6LpywVsTzc57
XV4ERETfK6k48JFSI7c/0cozHuC/2c94Os0sDJ2kI4Za+0P45J8vGTwxSnrnqIDRMcnVAm2evoZF
kQu6Ejmi09awr+xj4C7LDXv6WgMm5SVk5RBQMbDRThg+XqMaCg7vkml2qs65PsOyYx1vIGPHDUKI
MYsMQoTs5rlGDNt2U6dsNAtFzAh/bH/nvWX6hMTij3UXFMl/0a7i8WEMWa7u0Pj6KwKMMAgUeZGq
ZO2R6V8GH16iBTeaD/zm2wLD4HC4cyxOHaKhiZzeYz2XR1B6nfXiRFXDE2c35VJiyC1pwD5rAyrZ
s0Uc6KnmzFt9sl6ph29Nxt0uvmIywLHkZwmZ9gKpwhiWIMi4XUIEOZQvXY8noyg0ObandiGhJVb4
sY8RGSFTFc9D0sGsN5p8psELk92hc6TtER7cBlbDNjR0kBAKzkB+gcNiyUEbXF0PJ6qMCJYsbv6P
cJlhLHvTNtnlroYFBFIvlZG2uDASa4fWJ9lrduaDQy/thZ06gy0k5qRojz5+kfxRXmlxzNzg7nsC
8UkNuCE9wr0GVfKT5fwS2DDzZIFExQFlAsM26dQSbZKFzPBlcVowyfxP7Tkmn7mXrcMKaMRNlPqn
BMF7m8/d/YGA6/M5EyCOr8Iig7k/7bJ33ds7oSFZ656Ph8/ZJmnD2fJxbBhaX1k0k9IXHo5hHJ0u
LfcdNXLQBkzjtKaC7ijMCeMsin1vrmJkBvQ1d0xFihgDfw2yoWEo0nR7ajJwP8nNzBcd5DUpqowo
cHMXOcFj2oWl97E+XTTwwT8vZhpYSCkO2pP/xsiglzGPGWAXbe2r5x3rXceGxPrEtonQJ6JOWXKS
vuu6juDZp/1fNAbyB0h8fYJFjbcdnYggeEClmsTErZ1JABRGWWyOGn1OZu6l2DqRndX0YFHqwMYq
ADEj3OKlo2qjiE6S7/md7zi5ARAnu5dd1VNh2imVzHo7XWNhsGRAW/a1Bmk92EFfdzcjYxV6ytXh
K8AcykX+J0ltQG3BYWZJu32boiwRYdWdM1gvIwa+Dgt3X+cIY2YkqiQG4viDciUWvR5Oe5sRhR+Y
q6BeIgwPZ/y1IcbpUP2a84KXBSgDKhT4Obew4mAiGc8YDbaFEkOwiFzX3Sb5puUlZ2FN3+Qp/W1j
JDH66BuKjchJMjZvvcPuomHvH7SHzXam0o0bo0ONqRMtJb3jTuNNgnenUyPAPbNndoIuLhfFSrYD
E59Cv3xbIGM7iFsSqEz7425U3q9sJ5zRiu+h6mUM1IWTLZavwd/lYXFSoX6zVbhhY+G9r3uvyb7M
yvZba5nqHPGwJtm2YjOJ48f7Ais/bJjvfiww4hE4AI//71rTy3TzUNL6Vz90GE4zlcdP4Ia2IuBM
o6ftHdwBn6HM/08mFcUEAHX2PtkoITnZDBej/k6cqqCDYFVzNSI5k95CckJADHBzyXp2h/5AhNsf
NR75ansOV5aJ1uLlA+nVLuAyZHjkJ3GTlBcEBv5XTZls+6tT7c/1Zb9wAzdirYXY/JzDFPKZeVCc
x1DLwFiLcEHzm4HoIi7B3iS9MJ8itnaC3fsQZbMOg2QPgeawobTq/N/+CUUyKeYfmW4cUWhThlyN
/qg3L/eizkUxqEbRgG6Lz613/6GbMCPdo1UJl1VgHJ25OXoe7uwULkCQAT2C01ZHJFklkoUJyUB+
/WDLTbQbzc747dXtIovLIEjHsVtmr3ksJXP0JTb7xwB8dIki4+UabPfvsUq5bRyPFOu+ta0qRXPc
dEpzsZlzmU+iSMcFRmf0qOvh6l/olIU53IpYumvVJwwi5Anmdp7qY95JiPGMGcZJEB6n+dPLM8xO
bpveV1I+fb1vrA0S1QMIrCEAB1V1nAgjDOWlpxYbJEKbqmJPA6AH1JUqubk9Ql7zkDXofKQOBRJD
K5uaSudUd5U5zadWJ6z5Ntpn+279Wl4JtpL+xiAxdwe4S6y/YYF5hZwolONOXOMMPP4EWf5WAuMA
0C1q8SHOt/Nfd+QfCz8nuPStq+sY5GYCLOfo802YWZZF+g6NwmE2HX+QznUmY2eWgfYv9k8KfVkE
o7fqrydixcYvtFAbAxKVoAcr0mXTDQS72q4Dna+UczpV0uV+xUZiP+RxWwgfxPIs4ETbRs5njRcu
ey2iku+caBAbxi+Y44dsfBzlVMz6XtQOWHWJibpk3T/fph1w/JLZSL11B8mDFRXNO0eH44U+/j12
qf7OqbOTigBGTIOO+KBO8288BTv1d8Knlio/+6bcu+q1NA+swcUXaU3UkVl7GO9zovA9j0PIZSw7
ezlOzhcWWFM5Cq0j46N32Px0h0Uxt2uKzPa8WqGoxSGZTUgUOz8pmF8d1hw4n2nHvDI5pDbsSogu
QbkCwTTnwY3SlGuwmev6MKV1Lok+rD7bYnzZlA3G74OqlEK+x0QyvfA56m3mKtSd+yHHG9BKzUXE
Gr4MdNRLxAzuUOF8qN5SRyciI7y5EYTBfBq57OTWpo+EbizSF9xn+QjfRosTu+yFpFmabdcApA0u
xfEoSQA5CkHyXhZfvqXXFLIscIddPMzzPT//0dnmaLSQzPIGUWAsVMcFtUh+gAggG56Hffmb/yrr
SSrH0ll76ZAJOg2r1llUL23jSXe/YsO3eP5Wc5j0qi5IRQAAn71G53GWSNSBR+vSpJ7TU1U3HoWW
Gvq/pA+ltbGRG9qwWUfwIuCUP3dUor0S5yKDqr2gCwTveK4NxSp5snSFUsbswXU6BZuL418lS72N
XEY7F5SopgDIGI5VuNhPlIqXHhKK8yW0U3LMyhFRCrEtVrOUgZ8hnhXuPmtpxFfxaNhLepVH3Bqc
QOiobOkFbL84VOhZ6tEl9CyXwCcF5JG3Z02UW/DV0wnzN0u3o6iSdpIuqd2hSJRpEzUlk6jBSbLc
Ybc+ee9xBJ1xHLA5K6IGVf5SZSLtl6WoQnOE0R5M5+qrU3cApQM/VIlR+LNLqOKLF/tLCPdU+7Mg
TmIlaE1AGx9LglAfp5K39VEQBmc0Ulk3YsgUifqqwM9skIEd01Y06rxp13VzBukA48mdI+VsRPQo
PZi0SGMIDhEw7Arn/l9DU6X9nXf1xTd6HlrTyZ8R/n1dYpNAURi+TcWRz6XWhEAqSF8Qq2JADgBZ
u2lHB7AZQ3Anl8aAtBgMT45m4WDNlxivwd29jY8PVfmv2WU6vVSVVJKaG++rNWExwiyANjHWEskp
onGDKRmTBfvBxosfKKYIbRAjm8UnRNCaJ3DnkVFa7n0dSyACqSvnGqTX33YPvGcOxRaNa403FM9u
lSOElxP0gMqa0Ds4ltqU2awtQg8hjAq2c6/FvSmyjBAQ9NOAShvlZel/N4nn7kH5gwAc7Skj4Fa9
MPRsFVKVdhZI0u+kkAUOvB+PYm+pefWpu/TK8ieLkfCXzl8MJRUKMd77D2T2HIe97kZOvT6EiRFr
VqZvWXP1YavB2YEogk1BYLQo+e79puB+jsLXyDUvKbG9EFGjacJaFHU9H49o+ug3MAUjUyI19BMs
2TCqrWmTt5K15BT8UTpWRlGiAU9ID+WQUo5+okgeV4vW6CS/0A59sRc1h4XYGXnP8l50GbIFd8pc
8E04/ikuIucwHGGtCLr/2UhCnH10moWga1z/rLGZ+oX/mtIYws3bUI1V0EoTJwlYIYFNrf0ocT7S
jyFwuziovnU3ElT91jaQSjzJV2cOEFzgGiOZE60Se7TV2lUQIekxgzXzgVPdJ2gacBdZNMQM7lCj
rUFUxzmChvXW9jPv2xYyPcWluzC5Arlcb2R0PzaHbx45hWgahYc+JOytK5AAV9b3gyOCYE8u7+aO
y09gjahwbac9NhOe+SuEuPiJJbGZjoPB3mKEuW1Yii7YL7rfHoXlVMtff0ZcDNv8hjlxleGJ5m3C
lVhWEt0RjGAox+Qqi4gBT5q349KpghzIUyF/CEbFhC0Sz6cZCry97RR2V4Q+CmlKHkTlJaFCGB0V
QDGSyF2tGv5SFcca04NfsGFoCZFqrm62Cb1EpXJz9G2oUnKb70dT/+Y3H9U5qbyoR1Z5glxDtO2Y
5Qw2bWE6rqVqoYCPFPsb08zaxUsLy5NvqyNUY1+go6sR9CzEPFvBrYg91Ym3921Kg+i5jIHDY3Jl
kGq0KL8gSLnu+jrbdw8MygnTLhbIylkjKMl/9tx+ZeUXAdNURc1b13Y+bZY+XDpkMphErb7F2TNB
OZ3o5rQrTS6WKQdqraisfXVXQWco6zHMQ5M+djGdG0nnwfuYoTseal7aoYl9iJZrkrg/aNltMYaO
DzLgKpZBya2jKRbxi4Z6cJDDCaYHZKj2BPmmRrYqUrAQirdT8NfS1AKBsuS2x8yQWrVu7aAkisPY
XkYXIpAJD85NizoqljuOMZDStCn2lq9uEvzcsgQm5pURI4t1hjqXIDCTYkyUHPMFSql06X05S+iA
D5ukQlpqT+yIwM6WHZUBSyZAwYgLrhpZBKduhrGsmleJL4Wdnxj0pHgidTXHijaK2rSglQMO8E0W
34skMhII4Je5rRV6AmGr0ve9m5no7tSEjFekmy//k7Q//7lC2ycF+QZcGWHF7KSL+JKN3a5p5Pn2
9dCYIwu0XPeHBS/jw9XXR3egihp0pxGKFXKeW6ww02PkyB4jHlSfDR9uurQuug0qokStDKFMDFGT
qkSi56FXkablhizy9BOHUGiM/b3PYfCyEKYG69BQbLManR6twttcomoixc0ODy6iwuM7FgFIe45n
dlWdWiPDBjf1ahquzoypMTqggnaszhlT9Sn75GJxQw3DOni90tEDk0jNlW/2colzKVu1BLbDEyC2
OnNKnj6/TR1LteFxnnOy+psI1xzc2ECIJi6KrqmJz3HdGSHbmuuY+mte5nXA2pC7a3l0agu+cUzH
Ki1o8hSplSEBx7fjMEROK99/EL/SpXGi/qDR6VkdaDhAZzePMMBz1jxSmplyHHZniBS961zEXgPT
FweSvsna6GfyDUNCPz3KEhdkX/wusf9kkr7a4TVOSNkZwar6+bHaxzTlWbS8S3Eqt85F+1qnmFgD
CQhvyPz6MDvmVANmr4USNR4AEs8hM0vLNxY0Yhug8f5gJ5Gbl/Pn8tzB4kEhlMCoaDb95ohjDmmE
uE2KoOpZzMKBahzm6JMR+1unXycdtGiNDab75vQJJb+UwHv5AHaN8vTcIB3nZB+hBQxcNwJTaE5N
HjRyzR1sqX4bG2HB8CUY50fYNX/yWcuJZrUpZEVFiihO4tL5xeX9VZHzRFLXYGjrZJsmycc/IPq0
sN/E1BzA1kqqsS3u3HI6AnDKTcR83G79flX5mAzqbT0+6BZXpsyhn1g2gKi0Koxw6SdFTcZaN/6+
wzypmLaKqRDcB4X5e0sZAU3JH3CCyzUKesJcehyl+gb/0e1OuQ/6w/pSs0lPR55kSIgnoATTGn/i
8gCMds1wdIiq1NESM0y/S1H4wMISSmqYLjLRYeUqfycd7w54FOXCf5UExJScgsBZp31xtnRJcJeG
tH1UgIytLdo+If5ZeCJ5kYVoAo6oGW63RckMEGsW94Q0A2MDaiSJsFpfzNFy/DZqQ4uqTMIbc0MX
y88Y+fFgO98qXCzLlHHE16LX+ZjoLkMW0Wi1Ix0N58mgYiujdKOMZN4b3fJjMdyd1+8xNV5hlZ4h
luvF6wiRmiqyZ7cNmCbr200JIwctdgXynkIAMz6aCycL7qUu0MREs4kMCqQnHUjTbQxwY7ZcJUNj
3mK84aSsbC4kH/xn9KjxZKsMCcCqCr8c250J+DAUAn17Tdt99xgFq/eWeaX1H9nmP8SzPtv0Mr8q
o2aevGXQcOipKRZ2nMvFY1UC77geNRxYdiCG95cAKfdXA//Um5TP6EGAL9Gvuf+wV5h1ARwkxXPM
FxAlb2Oo3CyHkEadrrOzweLFY6n56qGthP/sW7Zozqsnf54O9OpIKkrYIoFlaz04Pk6PEe/QF3EF
N30KHZuUozlmAOB79IW8gHWOB4Gwam3BesxnO8KC+FPjRzs1bgPaMV7ClD6tFDTJKE0DscBT30o/
OIvS9gua9NEAz2t+SW8O48VDGnFfFZDCbOOLq8ROuaCcUMuONr95TVkgjsyxzoCij14VgEc/PlT2
WB+idvqreOJcLBF1n7Z7x1DhS2o/UuJ9vbSUrHko3NuXvTpPsZLqD2gv3vdM2jrlMKmxcS8nn5HC
slAlaa9H3D9OsgHlEuYYqCx8bgh++U9F0Lz5fq95KPqtqP4DQ93FAbIohE4bS59Hvo+Zm3fp1T7v
+gYbo2hGbF3buMsbzWKb3ldWFZvQTikBBPN94m6gZLt+xoiwZ67QhSUyU+Kx25IVLLPUVehg82w7
hoiJt3mWDwt0rnIJk2AEH5yo3k6yPRPHDCiL9kCoLHgt6HuYh9B14oDjDMoMODD+VMaKjSw8mg3v
hlMDXKQnLSWRe8GkqJxVOArV+Xv14PLMPQJgCoOu/WIAV3G/w+abF3RVtG+28RenRBaNf2kDhDFv
vcjsf2Ll8Hooq4tF4AONxKwJ8vPEleH7zGwrZdm73TCVQpXvXW60i3KW6YWUFafh4USU2oQZ6pz1
70txlSBO8Oxtbu22Ze+usULiWTBvxyyRPDencglbKAfeWFh0ID6MTDVhMkx2U76ZFbnBJozk6MXp
mZKmFFEO5f6EwPuO/UEjCFSinVZuK1zrQCqe49ULNmkVX142jtGltzo+KyvrQK8ZFVv+NMw2ZRhM
6iz8Vk1LmRfwclFkUhJBid4idFM81elnyfw1Vx4INSbBflCaxFDxfx6WE9xIrtqlFfcQUEtntgbj
P96PxrcEAf6utgrM6VtA43Fzf8yzCxydCz0Czo9cdw3d5qqlSZnYieMhPXNSd45vCdQOdK2Ysmyd
84vgeSObByHLaOnlB8vjEBhg9PXzBZa3qgtEAlTGJUX/Rtw/vFyT4IFwqSADfSaaOQEPRkuf6nLH
vyuaXr4UHVEdx/N5qvu6Hm+itKLQSpBfoQ/bW/XdjDgrVgHAz+GTLHA+5Xp00CW9FEoYbPkOe903
KNxLSgFrpNBEQW0iQ+HnOLomw1Kq3gwBFR99pVHZnqiSy13Lwvk23tMJrp4qhx7iPBCDm8FS6HO3
5uql0MpuSPMPbrlHITUFLgHRqMEIKhjJP+UuVgGBBZeJATf4YhtMqqB/CvTCblLyYEHZOPd06j8N
Hu7rJs3tqXklLrZGUGqUySm6CeJRrCOxKo25TJesyHd3H1j+vAxzxSfjaQCmvx8Yvmk3Et5/UMiL
qIV9maSZRroR2gdzdtoz/Ip6r35mHkNo19ou0ZGRHH+JSQh4IQV0b7q9K8Es0RvInuajuH+3Unnm
Jk5j0wnqksPuCQwLnQzt+LdZflsbbTSTqoWwhYFRdYHffpNTLkiP0s6y43YPjklo7WdsIhTElSr9
WqmntzvdFdhvso5sAL3kaX/ETY4pWzK9VIM9bFYR1HLMLTwzQJUyDcLrZCkrfGXp8ia62Rj7BP5M
OpUWUg2oWjkJwk6sg1vlhAAcNe8bu+EiDgO+pLXzyJIQyeW+vH8Np8W0NQBXF6AP4RhhJEoGgzXZ
5MMQR1FCtHxJss+lKhpXbzXDhSkx01w0+gPIRbnP4s9wTKP0F8N58PCqC96QxPY66tsN7AAMgzQz
gdegveLFMBWsMZyDlhQwbaDGoMiQ+2Af295Y0P7p1bHKQIOrMIxXkVJSmgCsB6jzwtM5n3aHHzOR
ILr/yYG2bEPGjoSHiC4pGc7aDZziTXzp2V6NonEbMODUK0BO0rlyPxwY3VAJm/++nH/Vx0/QKjH6
AT2MVxLAnCUGA1xmW5biMkk2fMtRlTcUoHFPuopezYkdEpN6YeKbgUx/h9eIphzoRdebiEquZsRC
w+LyY3bdCr1+2MnHui/M+cUb8x9mvDWCbHk67HB0Ex/wcPMuBS8Arskrp2IaPU4oMR5g8F+Y6e6w
Q7GMylunJ9LxUNLa4ziiIDuyp8tqovl64S4jsdR9XCrZrzMEqfQ1g3Y8Z7e6aRnVF3j7R7gJIwXD
j/mdMYD6WORx4WqHX9h6IBzPwF72UeM91AwZuOaB+eLchUPhl6Lz+xLd6/gnwk8BgPk89SGQD6ES
rTJO4VVpLOd7O3s1ND+iu6hi7CZ9rTePrlWN9AJ8VgxTmhvrglGKdoUjX/gGqlPocx4vKO6wbmrw
4aLmtkj1O+4Td/vF2LVzNv3hJEFY0UpzQobh7KQX0XtN5NOIciP2OhUBx2sQxQysN0gDBxK+zX5u
bp5xjkOG9dOubXFH4ZrU1F0hjucrTlG5EOrW3ty50rACLydRd/jYcH/T8ZhyI87P5kbCQJgY6NXK
R/XMwCAZ8o8AYp1JiIsvi0ZnOxewmRrcmwTRFmiwXNA1BvAxHcF9XQ/isgCF4KHLyqBqGnclf/vP
HfbueMXzW8oglFFQQdvB6bP0660y/Ey9IQ5Xd5d5hTIHtP4EyrN/Ynwwc3bfUHHiHYJm4MNDcRTO
Zhxy2sjXBd5I9re9xkHOR5GuuLkscUIWUvxyk1QzEjsX3PplUW/bj08ie943daU0/ZdIvgx/4uhq
h4UfSJYyERTI5jP1JdtGkfT5/x5UdWcBiYe8GvKoawCJGq7L7V90UrE1n+4AzJPN68GX1kVRt2ns
x7M/kiOOaoQYF5HQBT9N3+p4Bj7QJPhGQvPWCa+8Az7wnkQgXN3XpcLdIJ5fMYLiMF/NDEtw8HJC
FyJV5AIIIJM2jdEV32HCcs9b7/vH5LF3oFbu/frmBg7dx8edf/Jt1g0bJREA8wDceXwqg67hd9Dh
Hy0MCawq053MQ8Q8h+4+GcxAmhl30qekOKKfb//MyrFEIs5KO2Kfo/qRj17slc8T4JRjlBDl+Mqn
kf5vy2SCO/4TgZFgoU23FkZ69F+0HlgaKgE2X43L5Yc/3DSRAnglfwdbR8CXLKkS7bMNln9PIWRD
NYsGOzfbVasjVq9UD4Al2aluLwppkn/HeeHpqzYKdOiKe0Khy45sCParILX6mnl7fYFEMA6xIjYT
Rz0QL2s1dsSRp0IN+PYaueEptVI/9467PJIPvgx1z3wMoitzWKp3bKXiWXkrcLEMtNMzkTHdEc14
6js+5izditFyhcuGDvtcuurj/AqYci8wZx2UToBXoO3ke2w/r1klvTTSSS9LDAd3gtTgXCSsfsx1
u5fjxIgHYz8vCsbvYYt/ThaKZJrsTNu9FsnlDz+ZuOtjq8NM/yET3+gBghY1gfDCtgaUWdXIoWlH
cO6lvzEzsti+74fAfb6JRFEIBkhkLGHBqO3mOab+3siIXfG4xcQeIEbHB8sPYNIkxVKUHaQ/nP5R
tGFAdCeQw+k/lvBSibB33jSJL3E/yzRbwi/o3x2LGFLLKsa8pLfnrqjPPy516IwZYetzMIz0pa0w
rJaEKSMCxqovbmxC8a4kJZQdyXJvslNVAlJZ0qo8KquikceGnbE1344SsvGY8jegGM22vc/h6A1V
EFEsIkVVJN8hzz1n/HVgnfjyxOO0wwtqjj8T/ovRhcdIbrp7JieueVaTg6vg6PFZTB4CqyltVL1N
ROqF0HOiNLSI5ToberB7uEYk3cg+CKwTi/JG486DDqlQtZFQm3cByMp8uqrckOWncZSwkPdlGXZK
dAxSjm/AxLlAPVQpZ4FZaCSAVlr9gsoLndu2v/EcyyO2O4dOG0d0CGYJO8G0VEIsoZ38E+HhlSTR
iHcvgDBo0V84CfIKiqiY/BLoVNkoHIdIMbop2ksi+DUd5eCLnhDbDGXmyEcRAGTiqcYp3zEvG/YT
zHkZfu59su5Cudd6aDnGyrBMm8S47Q3s2oJ1Z0ANEy1thTFWT594s60F/cpuGU9IMfzYAQiUJYXH
PGB0yBAa2Hl6ESHTW/a+FVN4KKJ5ptyt427Fm4ECrk2UezpoZNMuSTpHJMpT4IqZokreQ3fOOPM2
nWPMuthFxqR23z5AbpEUlqIfcEB9RjBmEbEm7+EOhB3N0mvTUwJojHmvkB+doFa6IcaCvcDrcceU
suNDW9HX9ohknFo76jUGPpzvFZ0jFJnSi/pL/G46jL3iHnTz8Z2kMpTqCSJQyuQNrcsiCGdom01D
siO/YU2kKByqzXiR+2kN0mprgqqX4NyLlj71XBBu+LUvveUxk1+olhvss97pB6lxbTEuFDhbY7DR
OF9IlKvzyAGyleQosh7fTgNOUKTbzvFFKT/a+5khCMAJHv5mUClz42yFpJxNLVLihvt1a2sKEDzj
z/okB9wVcI1XfzDxneEfPnsVZxfl0UtKs+r+qb5SfsGWZ/ORY3+YViW/LQZkHUZeXex7b2UhXj0J
P2/WGAlcZhPrzjSgtgxof4mkrM0KQi0Qt4KvimSpzrqTLCQHWBlYDjAM8FccsmNwMP/Z4LBgwD/1
dNbHNyFNE6CJqOGzynqKnoVTt7vXgvcIadbUmZ48Pjo4p23A+Nv8VENmdlya7JoFhWcGidVaga/a
5oyVxJVqjlZkIjSX6AuVFLLOkFfEOqZ2VT5C9B0FPuTkMZ/eel7i+I9iIi/CBiXfoN7npz/2l1E7
KvxmQi7rJVwNfo8jNL5YbAxUm1sMGQqzMMEoKz3s0D8cTWCdpUygJLbXzU8Dv08Th5im1dcN8mbT
en1BU2l01HkbNxwEMOvmLt6GD067VmhdGujLwNT1BsDstEPBEcLKArAaclQddjh0TORw5s/7JxWf
9av2Qf1CHDmOK/74gdOWKTC0nuxycIKuKw1Y5Jo7NK4dU3/AgJkVKEdF6nLETw0XmLpJ8gpX5NAm
jSXxWQ3PDbGDJ7SDJjyIZG5G46LWHX6tWGPUgXroSanG6tg+Bbht6AZ8zk8TQg2H8wjKY88JAOHH
06QQCf07gl9xMobdwNrPfeZrNatLzGmAOcrzSuwKa0nEeEpgTIwHShhSDmRlQQHaEalleiXnVNZh
NBY4LxRpd/mP6FNve58Y11gM1Gvs7EmRi8rktdGyT/UjdWjoLFEEIQdy6tu62yPIl6tzm4+7OsDV
MYLGadQu6CGbqCSoXKXY/ZW/e3q4j6xBMKyrATbT1FTfkzRh/3I18bElVFLXoB79a09iP7MiIYBj
oAGBsmoPf4BOJPJwAtkXHnEn0mc96pTxSvhMnj6I3P3juQLZ21ldbdmuz1WIetuQjLCugMKQcdMm
l1uD4jDMHARy5pnJEzVI1yQR6Ex0X2oUPtNZ9qqdaU3VkBLKgg5BXQe4hiAgbAG/Yr8YBbOUYuyP
Q91kUQu/OwUM63oXWcdyjcTST0hMqp2q6r3sA5q2LLj3TsXqOWjw/iLnWYD1o2wwV9ilOTVu2XGM
2jZ8krLzBXF3WnzeI6S8egFuK/bv322BwgjWCNEO1Rfg+MQ73e/yfnTO+J3V2qKlGsEcqqmbRkX9
b+r88fQgLtm81VPuw24EAnXzSC2cpi+6uwo+44OE2uJxGia15NedIfF9Sd7mMk2/4y/gTaWYiIe9
2BWqFFHZD4Y9OoSafqMf8GpmYMQM9FjnDHzQu/NbLBH0S4IGJPJCnOoc5U/nYZOLDweNys1zM8B9
5GpPKssatf1pozUOIuo1a0Y0B1jHtKyM7UlY+mSkN88/rQt/2+JvZpBqU42ySWlne2OKrJ7sqniG
HjVlDqjggKlBKWoAKaCStSRIXnuD7hgzYAXPC0G64ehlcjoVb3DlibCHAvEr2udC/BQRzGh8sFQb
4oqvGUedWr8Il4H7wJWXoRJKzpDfVIrEK5g+96u3XUWEwGJpPD4y8/fN+HvUStVzDJmp23gru68k
0+TJaufOyEPX4z26tMXv1N0AtUOo6Krf9IutNBdgGjXO3MTx2vOYMtEFe91YxOKHqgCgnVqdbtmv
o1Io/nDmjEXZ3EhOLuNFgypK5s1npJ319On9ipYBo8TKaqKS2Wu9kNIIaHN+RCGRTTnijLJ9rCrA
lRKOzGqNN1D6YAv4gUgOAJJ1dwUo4jmqRgbo+n+r2kiFOGndyL7vszirbvPHpxGcaBifYHe5UK0i
ZCU3dFuxbfNTHWHMYcaz+jRfIrM+WSk/gndfWcLauc4rHGbp9ZHcNB4wMZXBpEp3QALtZjQCu+CR
RKkALIuvZOB65ks2EzWuORUU6CMgDWXVEamFDWqmTDgQpQjEZCC7UaOgDFJFgry9So35wWzk7Wui
Uzp0PsFai7uWx8Ycgs6xymwnAVMr44PoSVMN2bVY0jW03ZITumCYFXPuxSOlMePKgdEYxtJn612D
wlQrtclVmfpJ3+dzw7xryK5+lhfGCGnBcuEO5AfNuPsBvnroKhAuB3Zjb4GvzeVMjNHWolziHExB
5JTaR57w5UrcUeRI9rP/YC/uk4RWdiFIBZWZVz0mMZHtJyxVVDmRJT8s9uueWfEofNUuCFUWEKKl
rKy3M8ulUGm8i4WqDcICwIwtgNzshi8dn4hIb+U5nBM6ERC4klRR1AhNboRggR6bgZulgft64tRR
xi6r5HEc3ZfOyeF6o40Jt8nMW0pvbjR58joYcUbFxqY9GtYa+E+/2jCJWFCYi8pah8zSdFNJsSt/
xc3dnWkVDmB6LR76CdMvJ+faHRbZXPEHF9SiGcQ0ewlQKjqaMA4myDxI01pDXpWmgxk933QEiHsO
kiOVR8+zk8MJ9adAXhRs1KtUX6c915cmeJ6v8ivi5bDp9gH3L+iMhtuoERbjg9zYuinymhxtGNM0
3icV9RatkE75PSKUjUwG3TcqiF/PSomteq6vWaV4G0wJFsgxDLo3MN28o1V08aARD66uRT3EsHgI
fVCpFLijElT0SAG0x8jXYvxEtlxjSvyOnD9XLc6WMmQIPDrFGXYQI9YfkIPlLNwYI1qhiIrQNTfH
dHyBvQmCyMu5zmftvtg4o/DF8T49qrmy+9nijelTlOkMS18CsoE0tfMZ6QB48VOyKirP+WJ/6bhM
bm4/R8Ej3+EAi1x65dpFX+WTPTTdHjttwtaMkVBv2qbt62JxzKaxNw+ih6IPxET/+B1UBldzO1C/
Ac+ksjxt/PvfYZxfh1bfBFPkbPyEXf+YaRdi8lWVSZOlwHgtocPZ27wBbKIMqvCOK7UbRgmUQxR5
n5irOJvT6e2GqALilJlAfj7CFyrmbpoweTd9m+FZ9qEOeDgrHe6WGiymJ4vibxZFOn5dQdb6ZVMZ
D3hSMpLGMX6N/VMKkhzkZQaLgmLHNFm3SBms8Yhjyke0pDXkY+rdTJAKrMTsMeLqHa1Fh7wwt/ff
XWtyfSqqcK+/q7AWCSHjimwTTnCljZuKzxZjwLq5dj798caO8iaMfyl2tVYrsJyjuDcKcJ9/ugRn
T/LbsSJw7lvr/a87YLsIssLKZsktnJ8GtRg3MN9F/RZa5R7vnYS9V7XNAeCNEmm6OsuG0IxDjg/Q
WYMl66zeFTls/z7efT7//HnU0wC/Ou5sZ6tyFEIwusrwnnP6TBTteKyWsv1JC29UJM/RUmvPM4mE
KLe3dMuvS/frApT0SGzLhC7XTlXZ4mvGHgMtGHDMFMfUN8coKbWzkKRYlZzRVWfoVUYuSsTl1m0b
h2e9Ib9wF3pQnxt/HRXkYsVPtatqtj43WVudD104B7zPWPiFplGMc6RWvWDZNqz7gOjOZvJlH1Al
vPtG8M++bW1rFlzQEDUkh2W1d+7xswx2sZw4CNfz6rfAJ5JUz402wLQlHdttV+NGXSfmXqFVTk2q
0rgvXhX9Qh6pV1tb3Vvwwv5htyzZedx+Ho4akWS+WykQaDZ4BpW/tknDUmzRkVogcYa1kRdL2Hcp
pc53+DgZ3pTDKRo0DzSrTaEzn/YobqpHOHCAURtBdUYN/M9XVyLeSsX5zAsJ8e+Arf8b2Pg+4AS/
Jmow/SWp+473CN1W2UGtncuelprxeIbunwRfNFI1oUcN6p2CaHp23Sg2Up6Vsr5INLVcXuOBCXqC
rnHD5ckqGf1A/GyjomVv7MUDWOpY/ktDuaDmJiw+Oyo/pi6pYHAfzxpp5830denHZiBMuIQx+Xwd
K/Yrsuo7SwHQFtzw/VOt7W4P6GkWugEbiSGFRmHMztHoEYhnIOysIvYq2KMLyD4rhD/4+x+eYCy6
MA9U9xdeyiz6BGEETmVWmPsG2yBuwzUWIJ5ERl2scjQ5pwwzkCOoDP8SKw1ZduFKFxTdsuMe6l8W
6XDvorXUP6ZhjbBql79LTQo5Ulmtv2YDvk2qvKXhjpd70idNpOHerDnv1yb+7B4/BoMEpyriy5tt
wCyOqk8Zr1gGPuW7GVY51f9uIVpL4CNTMK70LE8Vaa0S1RR8NTpuLs3OMStdm5P5sckWJfoVwnxF
rzMiwwpJp2PHDCrxhgr5oWEOzpLr04zDCxQ/pUjpXo0/kwe4EUCsgCurTL3/+2mDtaI8uCm00rJK
5ynr15bwS1ibQ8lOMjS7VaKuIGGDixY6689ZjvQCfEAfy1ohz4wy8Kzc7kpW0A+wp+YVxDcj2o7y
tY09tPaHSNGLAK7IbUlC6nXmSimnQp5FyGDuSRX9auHKdkmqoXQKnPLcPvloShy6nlaN6z/32K60
qI+me0JtrsheTyk4EhQRX49MATAqTV79jLO/Jk4B4pXceRLa5jzxLJw4/VJCDEigoCzpCdMS18lp
9otF11pimpOIfO9xFPCMCaoBYJ904atwVt4yaf9KSGzVFhZ48dTas4RIwL7EgmYvnGzS4SY6uvA1
y53aNPZLhb+CyMw2DEG3pCUEYtD1oTfJEyPcsItesJDg8geC7c5ocTT5OMst4Rbbbh/LmH6BLGqo
vBY/L9khbwxH+mfKzhjtdnGVMMNjDja+El4W1mOQwxxwBMGMIX4fQv3XA4fHQc2xMQNbJ82s8eFs
YFYt9H2EBZ19Skq8bk0cmsI9dSrcjjaucrLGrUkOto31n3lFBUrhvSuStP31yVP4jUgCIn2Fteb9
iGaBh7iPDjxZq5BKj1K60yg+lK/fYZEwpQT20Kl60JcDc9JW1Ap+hFr76YHikh7p1hO3It8s8pgK
2qnknf6VBqayb64zUXyGAWRyrFQtk2w5Q3Dsz3XDhHDZdCf9XobjQjcVuiNMfYQfs6uC1NvttnyD
T4LCfpWYcSYr9Pg9tizJO6DVAJr13TclfCD+8l2Io3YikqfE+Sl8h2XQycEFftLjxWAPK0XmqIPz
OTMfnP4FQz7/U3Y0uZmQQqWlbCXzouEAW4DkfEakB+F2jHUuEQJOQjfrs6FkOtIHDcAsuNkHhQGg
NV1ERTfq0t1fHCgz7QmtPIwYN1kWXEF9rwYNMBs3jbkeqjLgE4LCChNm75Ibj3Ddjo+164K7Ns1k
3wso8kAGoWFq63JpngKdiU0NSIgt9iC784Jl/Uvclu/Le5omVYJnsxYwvK1I+luLdS7RILpiWA0Y
2Q0TMNAlmugyADzWdmx0scXrgV1PgFHGFRHrVZW2yngmpYlr7Xl1nqWCz62SdRei/u3xOP3/VO8c
eRV9moccY8KZni+0Jqo5A3qPSwlE+gCod652O+VAwAqo72gIDOs2d+ydFXibddXOAZ0pQYVoKIrP
KmzRH0HlTGMNrE3Gp6LBwtvf0DC0akiWupEqjttIT5Ggnf2MqiKCGSSjksqCW7oJQmHE7j7fOKxT
SfQveFUgDh0M84jEXUMfVWsSVD/K2Xtuji1srnjxMyNYk67XzeffctuV/26C+LM48i2NpjxgX7j4
nwCrgFOBNPu3hwumzXlQgVigON4IpJs74JQbx+i4iMDQlHdwTczUbY5GsaxunCNOFIMfj1uznm7M
sBkje/NRAuKnC5JGTJOeYydpIJ4odnTBArjH47Ja1tCxEd31P4AdUq0/Sl1YaE4kzNgMi/7XvOjG
2CTOyqrmXPV/hRZVPwJoh1kPOxzP1oZdsM0Y5iQgMCUWzpF9XcbhoZLaq4SP93xdBnHwa6XDSU/e
UHuBXQXZr3zbbReHXXjhIzPYknDD/0FC9sCzQ5P/iFRzrcKfCGni/rAIvniJNQNNzI2W853VUcmA
HckovuLjfLRgOWvd2Ai9SSwh+SDpAyPwRKAH4R6FaXrd87u2Iith6lcwg7lBWYFFBhD70vcHPrmj
4h6Md7UUGVOWcDtxGIexQRhg9uECrjsbHUwaTc11XHh4PoiQm16lygoysdkfNJ3/CA/wPjBYfHMm
fghJ7pvWETYa/+SfsPMaRgqKqCuq0Ku1aEfY+hTK7adQXD4VQkz3vAaRtlvt4avN4nMfCQkSYaX1
uUgJJ8qm6KwxxDi39fMwZiFzJBjqcHCpgHXzZjshW/OPCq3lu4m7nyyhuqWlKyufj+I0K7BBfgDg
C035V7PjHXNwH/UAoo/26Kq1EFKFCW5/2re5wOjTrD06LUGnEvg0wULTR7cgwiACMJ0hn5jZvxjj
amXPLa40SpK74a+v/E3sgqXEWVtUuiemVLhpmCT8b3L2X7kucALkqXZxkI0zD8ObbkQXCuzBbzpq
H0Q1ulGK2TYfMqkl9teu/B/sgtZbb5w3QBU4UtDuTiFgID73Zntj4wbC97aBkqeQqslCuh+YMYHp
yowaI6/Eo6SdrjE+mSyaK30M4GVJOWSH64ZHnhgg53EF1MNLzI60+1L/xemG0+0Ve2SlDfuHO/m3
a4QhqFAYc0Q/0o68FKtZ2QWavYbFGIX0UavKc8llBS3Ch4FzNeu67mrKHgFT41j1yqTFqMXuOMoW
JSXibxHOYEIadDZolPHLY8JGGYzj3fbdJKOX3HeilxiE0U+YcQuW2yp8ceL9SjmMFD0y0onC6l1f
BrEElYT0vd8H1gEIStu42aLgic3SxKS4qTSMbH+in9fhxMuXKixXpwqFLjRDnXsk3svshW5mJavo
1W4f15r5iOgwMd/Kz5vQWFAGGgm86pYSKC37O4loYiICXGpge2u15KRwRBLWrmhSpNBnZ7uk8Z0c
EODKyILo0OxYsRZm6rxXsO8C2mtA0qwQrLzW6gS7y968DyDOR7gffj3orc1bGqyLWmC6I/S1o1WF
FbMIv5p+NEgd3q9sbko1C+t6pSJhnGDf+KeMqDZdov3jbViqBplXgemAsyO3tNmDlL1+lNpOMaGI
+JTmLmNLROpAJ26V1MpSPw3YS+93Dt5BmgC7KzHTEr0iSs5o7sE1NSXijtCQlnCaTjkxOo/I6l3A
8ObTf4zHf3ni/sUcId2dosb6tnzM+AAddidXaDwRyZuc3Efey9sqM/FV7ZygcQ4T8nTYKrdVrxwP
+tRZ3LxVkJriLg8CCjDpOW9L6nZea9m5ZT+JGigfdQQVzq8+d6fp5XiPZ6XRqQj8337tXBc55ZGN
PNtzeOa5KWqZlsCxBXzKQCakeJzMnW58czt9MdoVr0RrU7pvl8aS3+lgZwemdwQ1UDgbNaPtR+pU
Ef3+Q9Z5DFRYFez2fuKxjivh+c+QFJslMTqtZ3z0hYzprK3svZY/58WfRDuLMx4Sf4Qh33ibALAQ
jRIu/XnbmkJ9cR8pcXo0z1FM7yLevIBzuVpVT/n9wooDIdExqJX2SfjqAs2SCk2VdGSzfczmOUJR
2xmfeGQ53CStO2rSNuPVcn5xQX551/Aw6Ex01kjbo6/3A5hs66zRtFhyXIw7SygmBvrysxE6l0Lm
XA4Bz7nSkpYLbTu8C87XIlpxMJbKsYVEUCvGbw58JY63RJKGStHyW72uR6MZvOUouaKaUBcwUdDq
xHOrJ2DGycgbyl4lDlkWXSUe5EJgZhk0d6ISHxQJsekZfLJ6yTvwFN5cN/dqg0bZzn2+GBHilj4I
1QCyDWiep8sPdPYhRHrLXJhNGxRc/JRFaFZ40nVKzHtgPABV++y9HKcz39bvvD4cpFd4jeSCYi+K
F2UtuzWHxDmF5vR0U5JUc2dPmiOad1//oeNEGw0JBDnADI/J8vqVmZIwA27Opv5jplcIwZPYjggC
7YYC0S4JHriVVd7FMGnuQ5hUCDyLbwKFQQfahQN0V5gCgryYvL0PFBJ/6f9H+lBVB8PXUZQ2/uby
UPI8MPTYKH2SfvaHH/fveATZr6WwaY7WIuBwm8Rzouch7oZ2uD/pWx4GQ3yPCN98tZoSDzPXEJwO
YWnkE6jBymRGEnfvL5SnU7ci5B7hJ5pd51ncTWbCZY72DQBYTSJcATa0T0Y7iOtM6lZSmyXiLEqz
dNpoI0XAh0ScliYz0Iy8uaJFYMIydvAN2QoKJRn+FIxhBwHQT5fohMsAsPoOsucWCpx8cFBgpPnl
YaOBkxwpvMeR/G51vOkG6c6yk4R/GsPGarfSN4O297C38Wq/XALYWahGqq3VlYaKvUhYg6OrQvcu
GT2GikRgDI3OWRksz5/1VBl7DMtUoLp7+/HI/TbgH0cRcIoupEINxqk8f/VI7+hSvtNKQaLBwLEY
SxMcHIRYIT4ppyGXtnSfVMLvjCRS8NjzYKCyRPkPFWwUNPGroMtQYBnQMcglYpeeQ+ZFQ+u+inW5
KR49SIynZnxzlIuC2cJHQKJHuGHHpsoktjERHpXeAIGHhnmQwv8e7+WHe6BnRdNZAxEXQyndn+US
yhtAjIz577csjIIWBIqQIbRs+PzpUjgFES8iS2KYzAzQlA2psCdoEp6p3Wm9qqk+JT8MxUUX8RcW
EQNluwzq7ydVZ0Uj0S/8QKD+h9w3gJ0PDXryhxUvt0i6ZZdoIJBZmasidPL/FwFm7Al8MDtnnCp+
xkOdeQWCXYPNmwBS1WoZGlhkY/HVVfDxGrFf/wUP/9dNrC8z4nXnzope/dbkObdOCLjxikponthj
MgscX14SojQMKn2cLzcfSpFfuWplX79jJlaHUvC7Z69qrOzcpypWgeLOxo2xDZ7oKbCmwPNgdQEX
VMN0k5L9Zgs5pZXf6lXtxrnto4cBUXxsk16s7F9LuDSR+e5JAIQeYzugVjVfjCeELYDUq1sp02Bz
AyMv3686YDYn57VQxdBs9MxrZVVtv3J4Sdq1kK+R+v32X6cB6k0S0XJqd8UAT2CUc+Y7P6UbO2JY
Cu3uoRp7MEX2okcM7QuvLFW8St5d7YlwKSW3Na1GV4jjqRX8s7Oc77NFNmRjFqveVKSwRPsBPyoi
OGWEBnf0S9hBimLoUaXGyGVtNX78XS4qciwKnj7sFj2SBE4WMexZTJVyvlckxtAf4gqpg6gjSP7/
4OhMeWZiugBB3pppjt4IhjRFkfBv5U3EVfqzrpcF36i3zc6OqjLuVwXwqkGezxWvr3TwXAbhNb0x
LPHkc1nRIw580QtrcaeF+diXf14sLQ0p9H5TsGczsEWkuk5nIuYy61QczqYTskhUB+DQ0AfjDBfP
ylJkzFu+95WyMORlIqbvfRYwF8SwM4r9MSwC1d90kdWmBBiu3oYDL4+AD8yd7khtM9SVXYjiplWF
S8QiVT5a4N1MCJbJYTQMtPxkGKJO+NcWCeu/2glTx9DCspdIHlyfsfE1zBdKazhPIjQId4X8E1jL
J1O/91iuu8nR3cPoBaQasZWRzUoiiKpoAb1gJfgczfclYWehiB2Ctw9LLqfBSQCH/Zd7zMTPNqPC
VSyeHrHYCTpkUGHSFQLxo4STwox3P/PS9Rpy15q6iG1V1E/Qc6Tv0Hcw55Fc+Q8cmoz+6IMWAmDk
leE7iQhaW0ufp+Se9PRYYHtQ5mhZiSa1YnFmLql+dO9gu++OU1E9VxQ6DXFYLCXl9+Zu7jShHhw8
qO5u4RgfvHjvcwxQfq7cUnOk0t60/M+dbLehNEkpBQ+QsFB2Hi1q/uD0xNr7GJGCD5ZlPe3FvBE3
9uyKfVOQYELI6NMiuGghrB99wKVU0hRvqdTiBNDn4I4pAkoL+Y8ND7g+7qgnQMeYTj0TCZ4fRoT4
VShvnVq3lENey3DP6X8ptm5itV12f/pcSmlhwdSs01FE23Y09M05y1iKvN0b3CojQR5vcMdU/4Pj
N98EOzyY20toO1Urfd83+JNs2vmj78kPJqBivGXRt1jSvjcEMvfItqd915kZdBfyqXjEB6qMRR1w
s2AUDLg6qRZ/jWcclUX1CntIms8WJ8tnIZOoc0b+3rvXPe3J0rRiLE0cn6/Hv+Tij9M9k9WPfUaX
cI9vbxPi3o8O21aHj7L/+fu5vgGTy0ZRv4E6ZzVhMwBISmZTkOMIipQIUDjli1rOfUJRIM2cAPvw
JHiQlgJypEvSTEJub+ctwgCSXWCr4IhvVVBdjGNtwy+uwH0y6We6N40p8JQSudOoZBUbGKuV7Okk
YyEv/GLALb3AngzYHBkPV/XZAQrvY6Vfx1b29VgizSZDv2NHtvuycHpCm3KABnlghjbnEXk1pIBR
2imyCtFJ9PSY9y9i6fI77jLuC7LVRv4ldEvlUYoCexJe5HHub2zajdQxhUnD+wr3rwrlN5tegCBc
pkFesba11G40vA5tzPKtOnSTnFMYEz/r24Qo5/dW5zjiK3OGtmiKIguxTRcpOFgz1FPCNu0mghQt
trTwSczq1KV6xB0rNgz21gWjUX0skG/8F6m0oLeo60l5p1wO6GxlwvHFnF9WM60fHqYQUpeN65cY
Ioxzu+Ut5Yv/3ynM9Ow+m5J39+va+/qlJuIO08JeVY0ilh6O2hSwgmAKGPotIxQp9+3ndBSTZyB0
wvayp/hjSxbsO66W6863RUhiy2bM0y4srlXOyCHVg7pt0xgTEn/Yaoh6lvs7r414HhTOdVq6e3G2
XF0gei+oeKca+47kdD7P+5HKOUH4YCgOJdq6RrgzC19k1TU5YAQt6CM4lHwhCkcyMZuXFxXJd/gr
J+oLN9PDNplh7rd8VVMB0jqaVXOlGl9i1+raP0up04CT6fY7ZRUmkVyYbmiPlcnPbWZ7TNuTtq+C
crMR9x40OizG7wBDGV0v9zxuB5Houl1wlUHOacC//mUx+nTRSAh5kGvHIVb3VhTFCqymBmWbK0xD
Pf6omHd39GcBSGXts9FqQrGRnF9WPFbG4nQ4e2Cjm9ir2tLRgyYLmZ9RfrkGPRg/GgDC3rkQXMFA
7VDuIOk/OKLHJv/M6g8YDWrS2HIE6M38ZeniFQ19y4hkf3Ln70O8fsFFEzVTn8BykUE0JeTSHwKk
IGrXd+ycn7svP2nI+gLQ9QfJBvETymJGJh4jliV/vljHjAjEEBtyZuBCMFYOfWFwUze/ZgCQKyS2
prT6o6KMI2znoLg4oNY09sm884l/jDb7VxzgopJc3/2+Z2e9QO302UywzYSMgEvR9CuiqMVgC46h
F0+rMclGdgd5wWnnPTIY5zqYttV8kXKYgrhdHZ0XzasClZurNo7d8FgwoWoFxyLPN0YGa82ialpV
oBJw4nzBObNF+RbBSJ18EsolxJH/jpprdUNMS+0d0cKVEO7QwRq4A3foWvTzx4aNg/Vh8zp0zIeR
6tIMgUw/k3wA2BxzCvWDZLWHJ/zfIP/fMRpKDJBzRiyqzCBsPc+c0F8Jo35B4maIsnY8VxD8Z8nH
sNM0tf38DC3L4vgMUsLCmiaM879INplY5i0IJj2IvMTnEHRwQ4eauncOuM1uFtJwhDyXDAZwHLp2
0zMlLErznR6W4tBmiFXXKKIZf3mwQjaBJwRj1kN3ZrqdhB+2CjX62SuXQJcDRAdTgyVo7WJgqQbY
UFiLnpbbToEIlMB1T8KMhDzE4AMOqTi5L/jRElj/VgA6UcFfGwVV+5I4A8rnGCVQ1QmiL2tn0ZKs
1WuFzcN7eonhIK0LniTZSHQM30OxtNOTRhCLpqLUGSsBvriiRc+qzfKaKueKpP/IVIbtwrkGs+1J
jqSz5v8j2T7nL0MDLlAcukWofXid+gSuVvNap4u68nY9DvTwR3iwkktmHdk4cMI1AFWvJ/U1V7uV
45yyP/hz56iu4dLri5o+uG8XJZGK3tbicS2ROVRRDdo/inEmx5Km0vKr5dPLJ0jfED2nGMnxsmsx
BgJal2eweYFl53+xko4/h3GywVtGKPW+Uk1n3oHv7MxeRwcZfomnLEXtoUhWMBGD6uaqUF6Mw0Tk
1LSerDg0HsY5IDU55fWvwGTU2S8p6hNBrGsfajLTG+Od0ogJZbIHOLoBswlXldkMneZsqjm0lUH3
JaICMocUSmRtEEtnQpDmNbzm/GmGZ6g3bjRtoclmZGrb21mGLhkD5d8xuOVLt+Q0I60FAeY9aaRq
HwZx1vRpLC9WIOJS51IKbdrO0Qtl+ZnFuNivOTGZohiECXMANLLfPAApxjG3Ww9LcWs2xK+zwBHe
igVbSm6RiRZ7o3HVZGQVpEm9VJc2fZwlNkqCkTDiAQfimFGHiKMlpVtNbrnyd6z+baZPlAcKWzcC
wd5j8iEkXXxx8zTZRVm2UVTBp7qvtaav8CJJNM8F0TZPk7ZZ+yw/AdmGYq0jp+L3xLLGm8Z7eegU
yC2X2W2mCHexH6uAB92mkPIugs4MxFMRPcjXLNEl1732pGwplnXHjzhXUYyRzusAcPe5Uty4r5FE
u2aNO4u1+h58zrkVnWk1GEjYd40DvgUjyoq55uu91m+e8KggkrNjm+OU8KBpJFfIrqc9XtJ811jA
xdsDHq3HzUuMYKY9ouhbMoG7jW/h4uYyw2eSLo7ZnQOb18cufYmzgJYSI4sM0v+oO+svd9nwzl+6
hzCTu32K9SgZ71wd/9S3tn04o4gzl6iOecQbXr0i+4M3OZZTSWHoWsQO/tTxLbIe7vIxxmUqOihu
yMhCdCqNpzafKHqb6arx2/FPGCDeknFcqsKIX6vJFuEiEsOa4bEnAx/SMkP5hssKD0rRYQ47yjb1
7bGWWqj+/D6OZgtY3EwNwzRNKz7QyDtd9kp5kbGzier+sO9i2GCmX7wIIx+03xWwPBBU+UJdTQgq
OO17xzH/c80BXLDU0nbHuBBkF9gg1U0FYF8kcpfXNkOKIURezGGXoWGAqCAbnOI3vpSIM5a3zWNs
NZoiSCNIWXCJan/c485/MKkfQcwo33ujcJKT/7NHZtJgCR0qVLDVQsOHRWMQnuz3WootVNjoGpgj
pMI0z+yCWNRPSPBUBA27H5jAyvEMAgXD2bOtV6pxRtu18cYDy2v6U92wDgdzc4Dcl6xN54rzsHUo
4sbfTFvobJg5lLorNOJQLv4Oa771qvr+fVEyzind6I0H2L/tU201qCWaOBOqOvt980ewlU5z0uOW
69I5uge/dUK1Mp7S+i1why76Ptxj7HyX3ZRtWV7zG/wZDBaTitEBh4dGxDHE+PCz25OmzVi2mqVG
k4GWnW4ULbrcXAFr4r5KEsGKMoHoidwl/4/n9uZTtQb2Ni2slEcnKOhkVuHOLDNFUmRi/JXEuXdG
vHb21l04WNKDw/QAgVjtyspGcH3+cm0ejLWE4s2G1MvuHy3BZ0z5bo53EuvfcRnH9ciyX+Wd97HK
WNU7MDdOMeeF3tjCNSmp/r+ZZvF1bdLYvldxL4xjkmnNFUBNuPf+GFA/lArOZQPowBffxhYTZ/KY
jMTs/ekUzyGqdUDxfV8t9m2mNPWdLSxgPlE3B5R4Qy5iGzrN4sSuwaeJSoQvsoiJIqHO5uLjZLwO
XVEGItznno5rC5zzgQfPocQ14GLXLF4c3Toqr+Fyn6cyTyNxdUafWv2I9b/rsjA3bo/WOw75IW5l
l3hKfnR1KxhWQw50ypB/ngbVUtt3LziLPRQVJNNn37nKR7pHta2S//kROeItKy1RXvZsK7dReZ+4
+mKDdOcLPtRkrcsHJ243MBrms72F+VAh6Iu+1do92WI4xS44QdzK3yucOufJGR4oiwJjSTSq0TZP
5xDfUQVhCfayMxfWQot44EEZ8nAEhCxKVk8dcKrxp/JzyCTfiQR9/8K+GJk7yzm/zB4Y7ULjRqvX
uYaj//5OwOdbglkLHq0po1WX7UYnwzLxhkr+jX/hKHrKqewDUJIX79m4A3v/HBMuRX8S3ZaFtv8V
vm1lcZpSo1Aq2HjtoLNMbuTOOkrpUzga8UEiRNr1wkERay7MsiO4YJGIwJw6tRUcVKcOZ5MgdLnp
4gB5flbIqi5kxxBeCz0JtBcXkMA2WWCbRqVtkOag6mmmJhlO2f7A0xVrksbaADsLVjKTSN8TCH15
MmZ9RKYLrN0y4y1AsktHNe5gRYvWrAdoAqnFaXmDZUkOPveA/Q9mZjFkfGzLEggR/Dyz8X1lgkTw
QDaan4sVGBLbInP6CaO3I7ohA+A5dENg0NzWz5mM6hq5zZdDsqXLZIiEi2vXX0/1+YncOZwgmozZ
Ovuw9d1D+pYC+07yEIJ6wp28/IJCgZmfAhrQwNnVMJIIrlG9SaK5quXbJWK5zyqcF12Vu9JysApK
xcak48elPd9PKHSSqVSy1qaukhMMNWPZ3AEdcTHsSnxSx1GUhiF33ZnHCvg/xqqz6VHbRdd0QbA3
J5UV6ZTgQ/eiQFUbkYTtC5o99wJBDsVj7hq9IYRRO/HnDDhmsbjKad6SF4qRVVut1YgR5Rio0Lnl
ComWGJgEiNDnqvffrg+ntMpq9rVsDnDy+RooIc6fz1O/kjT/T5/lKBs6ydOeSPXHvOp+rmyZtvT0
CxoiSo0/3uRv3DBoA2zgXHlytN8K6IHeJp+NVufXhIKPxGc8qMrtRCNyoJ55IZUgc9+EwQRsjN+p
3cZM4eEwRLn+/0KLIAbyxVYMXyOyLAxbSGnzlQHkmC4GWDJZRHZxzrVqwJtw2jRHkjLSHVFAMPnt
U8f2rPlLe5C6JsEqokNjsCGn3xkuD+Wh8bCNIG/CFAvBXS3aM5TYRbcFM/Q3z2hb1fIXC6F3lWmh
RsmRSMD74u0U4rb/fHIOOh/wHJ8k23O32kI6BQy0leTrNArUdJMtpj46KKuGSA7jTcx4wcwmCxt/
l0LVY1afKAWiypaM1BR5iLQNiLE5+nOOc2lIn/Q1stb0MI2XQ9i0wE+DhV507IFzRgr7q9VJE0ob
2BgeA3fiPA7jNK5J6eLwyQnKBlLMU0HhQg+0GG9uXdtEIFct289ora567sIqy0cXRD9fSZFGgxdc
KbxzScURhSVMUhINiUSlJJo/1r4vFp3WLVxwbMIvf57xsbiwKdkxxAdlu8m88reJahMaltRDIzKb
XICyPyAMN2pnGH/yQmXmY2y9PHNQLu0lJMb+0KWxIsYcwZcFwGc3P9RCEFGBxe0osu60QcNB1pfP
D1j78iNT1hpMtJEublsmmzfaVLvxcqOUx+LTduYuIWWD+hS1begvV2hFRp2e2zkZQE/Pbrg8y1MM
goW4vMQGplZLR7Ror9SgFFZ6PV7JCaUEAHuXBjsMFB8D7uap7EwMNoJueo/0JjkAn054odjMM9jv
p7bKNZjyfI3hZUvr2ma9kmAfGvrgHrVIsroz2Ue/ozFhmK13yU/JO6GMlBkfoqUFIm9wToTck606
xkrl5gVpD51gXK6NE1W73Zh6IbL4uvuIDGXskRzAJawCm/2KbXYpPapXozOz0btnGMAqkj/rwuzb
y7d42t+bSZ8EpsVxoah2whKcW3PENuKGjmhQp6iWP+Gs5zkq9WtV8e6YrKiWP/4MWRsLEQt2zCET
AxQD0NwKpymYXWnSM2YUUW2tZ6coNtHO3XHyCfxixn0/+8ASkDneuLF9A8bNthGqLfUWhlAjiOBe
VQ+fRWBDjOCA9Ts5JpxpVF3mvsjJgsguoBDpWodWyhPS/GVXLj9ndieuF670mVI7nxqB3Clv9721
2Z0BJXiC15d8rMvwgFz3vIMVpYZH4siTDYpuzWwfvKUl/G6YzNai7PacHILUe4UMz4anPQcIKwvH
XZQ6teLu9rq2ILqNUDPnI5Hm9OhTLwza9gCWxNSQIzWPhXF7dUb7OOoxFi6O+peHt7LcEgbKepmy
etmahtCyR8s/QK4OOIeAwRG3cgLm0uYUAgSPB2Erj5YSQaWhqow6ehp/nCmWckVkdzjqvF5sxz1Y
1VedjSp3hStwmeSDcK3Czi6ltSWu+dLjO0BQqHnD/tamMd4YEnAB+C0C/nZzAhtky35sB1Qii4M6
LaoYFCT4cBZ/YyczplKk8RIZimWkgi3s/p0aTMfQsgUvZqujwejsnfwRCsAgDXzS+jp3V0UH6unJ
gj0NCkhSFH5a7HDYv2FiKY31GjiLtVlc/3KVdsAkphJvqnygDaYmJRgw7/m5Yibt1uyNgjQ4EFXl
Rgh5bVBjJXMv4c1q2BZmn+kwaXONb72s11unrFJ1ZP/Hhxn7DnKeYSR+ApLGdlxyfCwfeEpt4b5Q
IUoZftVsm6eeXWCPJMbz/rOf7De+SVDXDPyIhL7BZ2CYtGteXpdLicGVywBGEe2Q3bWVGfxsPXBg
vD8xzqLlbDbqSyK8t3wmdm+VtzXDc54EIY2Y2rLQwEabFQZkT4ID61ofKyXZp2GIfJsbwOgszHl0
biS+qEHWkJbWEx3QjUyTRx80ryfKtUN8PHvxyWF+NeG1pS1fJhoM0rCF64BOp8pTsEGqr4WfGJd0
4M5zjgLiMwpoGuNbfquLQj71RzSIvwR1I2qTup2Uqk6kfeYkiljygQ0/a+r4iTqESCXqKCZjbgpq
dKIU1XzK27w7ByL1xo2cLG7apVED76pg5GmrZJbg/C0/9Vbz0IDPBXq/2uqBL9tCb80OewkjjZec
YZjKQ8WjgRKSCPzBHRF8ibS01wc53FIXVCoG1u42Ialy6+C90KT4zO6yQkiv3+FXgV7s+KfkFFUI
54BiUiYa1LxLOIxnjgq5A9wzOqMu4/Bt3P5IqTG2StfUeNdNilZfaoQZB1yYe2d83WEzWntlcsuu
88J1CBul8BNmencR084riw9ZoYIzaqDZv1JugDQy9ihtMP8UYjusfsdXJpz7Baa6BZc4Ealk/xps
9IuRsRji4dQ7Q1HGFINH39gNIxwodTfsBQenMXKpfCQ5B7T57kkW+rsSwIRc1Jb8HQkjKIWPZz3V
sQdU4XS/20aFyVqSviLZvBtpjra5T9DOusbcZ+CDVr44U9XGaCC7mZRYK4eb01tRPwYsL353eGLo
KnoQc59lcfjd0dQ/r2IlSpgQFZmCIL5eMENNI+MA7TrO+pwZMRs7Xu3tjEVgCjn10k2/Sj6HO7qa
zgoZNpbNJ5lQMZWD92Oc7sHUxKobIeN2ziBP3t2dC0dEcwJXPzvMw0LIiqCPJYcsWe5pNdRg2E07
fqceHAxzfbnNexjwM8Ygnr7BEfkutX4fRgoAsC6ezNO82gKr8zVqzyXAIc5keA15UhidD+D20cL3
1AYoe7XIG3+t+O+ztF4v+5G3BJuMPH+47Kdnj30Wfpf5c42dyYFB1bf39MlF0cXx4MhBWNOrNUk6
8HQ8HTY5XS43OPOpGMxBlBdeN4Dj8yhm55YWDGzG3IRKXyW8qSn5m8iBoK2lNidStXyrY5Gr7kw4
9QU/KVhG1ULSOjtTDtZrXLRxMKJgrPn8xiys+piMPzOXGX22ZpR79uUl4dhlmxXssOdVsb1e6Nel
OeqmPWHyNeNyjvN5V6AgFG/I413VhXyYR1DZ6utTRyVZSev9rI3Np7T5Qet8XabOlwgWmnkkJe42
7uJcSZQqVDo6i3YESRtZN52/GRZfzOKUdz/q0vOv4xFnCPhDzfnnNW7h9WwY5lmYp1INXI3JEeKT
C4/TF9p0StGcNklr362wfhfhE0iLAXHRcxwQhQ9yp6nTNzbWMWh3jjm59jlQ0xI8vkc5h4Ik3Ag+
4mTYpecRyD0lCEbgO9fR5m48yq1VeDOhs7SWPH71OHl1oPFaqwXfXreAehVdNswPZEEmcLg7l7Yj
iZthHj7+RyHo6rQeahmg1fldRdTgkwOHaRmPG4dx/tNTdm8IjkagaM1nD9gKLYD13MBYsTwqewa/
OpnMNHcm2z+8PyZXCt1eix5nDjB56WWCjWl3f6KvZ9by6BzjCwjas7+83tFvtMNFPhA7g7yJiFeb
aSusu2I3KLOptgJFAFZnEBvRT0COkTy7C2/HEYhOkDQUjlLZyiVC4U0yCOzI6LAbIELbnJLjUFhO
iZW2ve3olHsYM3V6EMEOJfhXSzwa2aTWmg4Viiopl2ssZRiqr8aO1TitBgbkURArx21vIGKC+nB5
nRhau4g6YpezOi/xTbSVjgoNhozafcnjKDHWi0o4ujSQIJ5TFMSiQITwv3GN6B3SRSjfH2L8JBgM
3PFdH8xtYtVirZEfwnnFRVs43h32M4N0/+yCiP0rrGs+0Su7CkGmuJ0Xvy2ZHWc+szY2LIMtH9MO
0dcQukJE3oh+/OtoFYYX8E62MlN2HTjSYPOYnDBrSiUN1a6zMK15vfXeODSstrrMOBo18A5xwTFR
MKVNBfksTapgFeL6RT+jrz4ntyUzLLBeWYpC2k8oCPAxmeq9B3iingH0Dpt8LMnrNoxXIk7GZ9A6
tvANONSd2K7yiSXgLhGd0CiijfSlpa1kwHoFjl8jrMVyhiYM8fRxmpZbDn6pYHfc6Y2kJ4yRh/l8
B4gvKOkmlMcBUh/b2FxTa9NJuvLuDtoe0o+xXyS47RXsAYckhahXG3tP8jV9FYwEhgWelZY4X3PN
92PxDSvnoIZtSNu7QlaEISQw+cCwo4BtNTz4P16fNRKMUHSIv0n6XjLbE659o8WhaIaFB6sL6FLy
fhPI+VVD6ZJ8lb+WWwYV/lVKuOcIM4/rSwj6D+QEFvC5Gn9KXOHBxOiWGJbjFyEqGmAp2yLGKJ5h
FNjq28KAldzpscLcpW01XMqXoZYYN99HZv9IT0G1yTsnTpmNxCaj5O0u+fHGS6hxl6wvEcQo4ptV
0Y0InTm9EZ8R9QVbnkE31RYDAOGi3ZtVpxAN5dqlI9Kl9hS0CGgzkXrXRkTDuH2pjWqqDCyKRyBu
52raa93yKGPDVaB0WhAoeqF1Lupllt+HNYBJ7pLFgNZ3lIJPRM/WmIZo28Fci5ysG0EKJY4W+d+7
atlxhz5VbumrahP8VHeplK7eL9O6ALBCXV23A0VvVTfR9mf9GILwl15r6YE+fQaQuJb9y4VMwrpE
u3dS3EpQqO/sv1cDFIrN6YghL4CnzWWgCzCutMXTPamGGhyFiyYoCkO7uP+gVIbevQtIwg7rhabh
wGLeI5lAz8UyOfwgKKdJ12X0VRAj1b63uISYu5Wp6u/k0kV+bx3WdEbBcUfj3LnT0HcpfYMNvgVg
Z4y6RkzakhYToFyUDsOYuJ6EmcLqGqP5UcbsKqm0hlR4L48veuxEf/aqUYGsUy7lXDrfI3eceg5y
EwtlKWZBGE5kUKr/juyyCmcDmurwrA0DL4TGXoXg2Kxqa6u0uATiWh+K9jeEwIKGLorQ72sKY/Lw
l49aSzcEoWMn7Y7C6hch9VRPtIR+mTKZ8qx8eBVjPWiGRhyw78i1B8ZfebxCrsXdjUkpqz7PoQJt
eg5Y0DAV1bbwL9tx1SC5il6zKneHeBGuRy6lyjn2atiDh9EV1HdA47NCFbtFNAlbzRNVFNYCzMlf
/66HF7n979uI/kC3U2+FhWqfnenYqwP7boQUmLFzXtzboA5wygy4gHHDL/ndiWFOAu9FjPHkGmTU
dBm5vcYJR6ZWjr44x3YykxD0l/q0N27OPhtYTbSQZrgASGt5ZCfW7z7U7evTqOJA1nqe/4+/DNaO
UIR3CO9DXrgz4nvo5EDdrxWEOG2nhg1yO63Jl2LPGH0gS845EmoLS+oY8xbwmeUFCMs0zyDXaDcm
b88E3UaMy7E71uYx84GT/adi6Ca7qPkUTaN1FouTDLLtK0MNgwOe9nxf6T3bsz3FrEqJ8QufgUET
E2UdZ3e4bWR31++rsj6bTmQnVvUaLCRGAnaMRcSBl8rAtT7Bb3R0GdyVG3voDi6bHnS5uX6MEc8d
pGhC2QBH6YpWLqQtUy1JG7rXzf9Okakggsmpbbvnot/AkdTwppWEntNx3jog94lew+ud1SO8p04L
VpyBZwviD4S8Q92dKyU1ztZ/Jpnv9o5ZOR0FjQ6OE9npe0cnh7RwyVSRklQtvLir/Ij0kiaiF0Ce
UMDFfxeS55aBQRc0w3EPhQ3NaEkXquWk5EOWr5+6lEvUYFnaAgdHAeN0WSACpcDVpfCM2feWNbe2
vqO4UeZM9WEjJsyUyXhje+BvXA4B3WSOlXgQ+OsS5MZIxPCzs8LbC+xP9l2/wCwP8nYPF7vzL85v
cTIMy5UzSq4cEvYQX/rW/dHijrM2eNJCSc5P0NF2UyujaNEmVg3nu7Cvgpb/sNjnanSId9BExQBe
M+U+XjRzvn1Q4lt97xmmx7d1AXrjKVmfIzz0Nx9CYzAxvv/K3OzeZmu7bNfeU5tlpEXUhp4BaWLC
xmOzjzfVtCryX6Ktp5ViDaHQTlTr7Tp+PWJ0YGJgEUKurqpFqO7+j5j23Q4B0m1PuZg/kUEUmB6W
iasQ38kmV8jz3dJwrnWoFO2jn+8IuPHh0LkxpTT77qtsPzhYDLbC26tTB5P2HbjO2C7txMlcim0z
l8+8NlUSXVdnqnGhmA2JFJfrfMntOVF63zALfG6s+Hz8HGahjlxXYvPLmlRsHQhHHfNj6+4uyWB5
ZKOkhrKer73tWeHkaZ3pQaOmvRXNfI0K9WTsDWAZgDUBewGnTwV71Kyy0chSBvJL0BgL8MoK+NGu
O5PGZlJgeSk/O9X2KfwbO+xlBYwoEgtiduW6J+3RpbETVPDytjm7hWsNTfljtPTwALjYh9eUtcbA
UIyJSXuzptia70UINbFuZp0KB5DC4wlC6tg0nLXgz2I9f7r3OLk4tYXNJSRGSt7bmWJCzEzG7yXf
sQkieT4mXbflFij3jSylL/O4KRHoGS9ZgcklBThJmnNOXxKUH2QKK+m3svNH5yM9DZS5byGuVAKu
u+beicOZ7WfR1VTTeuuD5YynnH9Z4mDrY+hVye089VmSIUPN0AKTXQyijYS2ELGSZ+7mVIDP1Stg
c/8mRuZ9ACmzZCD3tuyI4qAFLbjPp7y3f/8NjfCBki45cyblbdEiIzIz5l4ekewly3/HmvTZ3PR5
0O+gcKabmZ5yAiht78mrKlFpToU2ZcWRmw65RlCPwq8IPlKq/KqWucUBIgHNSl79tkvJg5UZI3QE
IdKMPIY3VbtU+sVYaO6PAI3w2C2J/6GTS/v+SBcb86TrhCh3wgOoiooc5L4uWw8V7qOPOFxJZAKH
ab9929PKZjWFgXwg08gUC/ZBCG5B1SoO6FLfAhcQwy1fctiOe+oXa+vW7CjB6Laim/B6yjvuEbvD
wUxI49c/A4JqS0uZ6ARv0pE9MGNrg/o5JP8Jq6D52mOkkSD9gg5ZhVZHCi0meeyNAwvs+ffRv+38
YKJC4eR0BSqdH1ykmvesqQRnb1bLbhLpfhW8pSVB74tZq9bCb+IK44K4BxGomi3OqJJslacGHu0U
IY+0gH2ORQigZ8c5HGHpjPoshum0PuxlobcamwuAGMisY6mQIwt2tFTKsipF9V79FdWBdd/MdkPm
cE4ITosQASZq4CVT6pxC5IWZtQmnZ90vdwRi/mxXEeBn6czRTkl+dmJlYTVb6AuGVe2Y6SCYtL9Y
D0n2wsNYycAw2brLcKnFCI4IV3Eo0M64s61LcrCV9r36lIbgcxyDHvbBGn+3YYmBRScw7Q+5TNgc
Tbsx/Sr5H5RvjxNk9NTUQbQ3BQfAFsnL9H7o2vVxDzOuRcAlf5W/9FCajHfYhrk0tz3i8PVPvzSs
rYbrgIc4sahqlvWU7o3E5vvpuOe5oiyDyHPjpp3NDLixP+jVyOtu1nLwoFIdJdm1qXz0LTbbgK4r
Q5i7WZD+G/xj0A3ZSYZM8JjWTM4g3V4ih3tVp1N5ytGIfe2qLXxEieBoR93fCc7PJWQDLNU4+PL3
cdoYvgYKqx8xyFtQZvC+HEWWYxKd0bPRKf6thnABHM9+XoOwjXOjoiPrvi0fOECT6segqTrmWLDF
0Z41FY6GucFD6j7eDf4+PV7VhV3PWZOwjZObcZjC/GyMPNXvmbduQOwKX8SRlw8LovBhk1peX+hJ
PHGtnizIv+RKg0K3AsW9P3w1E0ZG+9HSzMlGLy3ZJc96IkXizGZ7Rz27Va2V4mA+3pSEZqtRKOLp
pZ5v+mfhaHeQwjI4Fj51mYzOlDQwnsIuBRU5nVadHhczsoFvGoLY0HluEb/6G50PGacMiXoENJaq
GPqjWdmMoJ60+OtceNyc8wJn83pVv7yARKaHKNvPwJvvOLO/FVHMbpJxJidxC+d4agKRX0zkvCln
xCf/D9GG0vBCJKBhFggXh+RPBWvlC6kRdDHwQ9r3bTC6BVi1a8cQbnDDN8jJBDBze1OmkC9v48tP
vVHd4M/cadk17ZGAsIEgXVitRGwTZPDT/HKErZJ7JZJFU0kGWEm+EFgibS2SLt/QG96W2JFEvLrX
6UTsNnZI8zVHJI7HdGPEcLP8AEOw3nyJkVZ1MuXb5IK9DqV2EGfdX+nJIpS0V9rZrtna5Ex9QgBw
Ch2ctYgiYFOgBMPNCJwUFQtL285gU5Riy4ZeEQF1bO7p0JjzvMccsrSTVg0/e4wXQVwWbroND9cZ
C/PcUaKs1ioIQfTDML0QCUX4fQd+t0yUr76A4oua4dvVhcR0cE3G1m2TPM5m1UrdR6KEODEGcgJq
mBIeWIr4m7OGukg3810FFf0sZbCTpV1k/yji48rpzp58o0LuZAS0n2ruv0xjPpTS2ty5yTIJ8wIf
EKxf69Qah5ViOafQ5zLlH7Cp0Ji9D2c/vyrnogOOQudU0DSZ+Ti++L6H8s8hAl0nSB+M8hxaq2iR
9+8CbvWGLqRNh/vYPDSyxe3+cofxPGg6Gg/WeDlYUd35N4iGsHSxw8yaJfA68W8cyp8njldJ9jjL
AemnGziPAAL4Fnmc1qvevS8CvvdqtzBY37HfXK1ro4V7AAAfxtBYkNDCvf3WBDHcEPJYvvLY1FCk
wTlGIgwqYCdxy3kgjzpAibh/AqJ+uJEGW2MbexR3HYnynH7IT9EU3W457poCkKSgjvjCWRfj68xk
A4lM6uHjGteaZJtnsbZtQH5ZxfxYR+EUsgJCPfuuofsRHjvixxzeSJFxpMKbgle6T/b9Z4dMOzbv
tQ0GF7TnSQKw3wU9H4sDlT9st5IGnoCoBvkxywSx0PZ4dVTGQBL2GdvoRt3DgMyCiBgg+VaZu+iw
CLKMoQ8lmZH+wIjyIHEaLdFAvFacF0yad4rX8KK+Cxt/DSEmEt0FIaZITokl1F/JTZZFR6PR9Clk
2OBbIOzy8wITNwTwmvDZ+CIfS/AMxedmrbXFm2EG1yKHPeBs5/vBuhuyfOHwdQRJfHUjYDl10CWC
c3XSg182pPb/4qcsxSVoqkjOmJTnu4A+kfpgjTDb5ZZHa9hJp2AfCIxa+OmvAERvjVHjrSLIUxSM
++maei8Ju2AdZfxGtoccwMF6UH00afspVhWR43Y3a30FJFu4Pf+B/3KYJDl0w9GTjAQQcvpst2mn
N73yVjHFODpYauA5TLkI0LpCiZhsM3op20mSopMz7sBQZkH2RrfXBlLfU5XjCS3NFHFVOGMQ9FPu
zIrKw9N1rNZPHwGa/DKHR62wWH/PJzi0kukFzfB+phmwLS/rwexWNTA+dy0NcKVfMZYp39wigrdu
g+mPsl2JLo5nexgelJArz09ip6ztCXtuM4TewQ2vsb9jfeHZsrgBn7efmuItYlplZbAztIgpPRLI
nsSHN2R8/KRoAaPNxEa0H/o6SGpCjxDHXVZyL3q6Ixg8+dg3t5/UzLa8almw/fPMsNiq/iHWBBVG
kNw5cQOMXDBTSIFJ79f+eKMYURsUK7lDvnQtKrsS6OHHKpPLotnEID6GfaD5B1b7f05hXoBtB/gL
LKQXTN3Pvk9IShwSegtIikmnsjcKS+1p0Cga//u8c41zL5zkOup2NDdVOTElB++1tj4tVGvfGL9u
9SebCKUNeeKA/HIwFj/ROAKv6BERb4lF9JtAJC0rj7ZZOQ25zTvtPvBxsY4BNemM16DJhGF8qGij
8HG7Zvq9pK2OmcaIqyvB/1XMjo3rXEkv7Tckpku3Nwmk1ugY6EsK2Yhp98SYZerPNjmlzB/lef7n
GdYTXSjmIrlQBIH5Hdm7XgcxCs2tIbBFOPyWwuARt8EYsQdNr6tk3dmNcYwlR9ZNuNFt+X+8p550
ieUZi8uH6E009jynYfQwE/l+piceMly3pzNkmMfbWPKgeVZWCJuIJo7UwbVgSaRHzLva/NCknS2K
WvPRVdhbOFkjeeit2vDecuoL/t7PPuuUNBQOnbthgJdfAcjJUGMbXeNXiM+JIXR3NrdqzguV2ZNS
wff+Bb2mqZUKxrFGBe+d4T65/mH3EZdSiKirKNihDODnMMtS8ds62AQ2QH8zsvsLlw3sW8Xs1vbx
7N+K/UpGITP+XKJ1f0d9HpLPvlJiRjVaE7j8eAyZd1oyhob4r+/JxE5p+KTWTxVbdKI2ASy/CI4K
sRFlC5UTun/9dRPYK6tD+h8Ocy3/p7VuLXbENrRiwnzqR1RTTUptfEGAd8+vOTOOhgdZRVF3oQ77
WGOzvgBr6QH6r8jKkMt1MkLnyqMa8WGkHe+DHFMpUeMUm/DN9l3sR7hr3CVAUFQUmyt0GneKR+wl
UmYLmkc6euWWAA17+Gfd5adBqMbDVv0PyN0fRk4LsCfLMIRmjbp34uAL0jke0ZwAyFvm3BMd4sm5
ddPEhwPXcHkpFIavhXMXIrqpJKlefA+FZcrC0XGe9uL3bqDeydJemDWesKpMs0QFy2x7SCe1PuRP
CJ8MVSqeynN0WzEmgwvlJGpVD4KYfiyAWa0gVaLwR/ALvzTElYLwhDri+Pp7/5RxoIRcbyJ8gohP
r8fgHcEgQ8+iTxMErc9K5xmEzfqd0N+uaI7Bdk50PUcm+XTzaM9w+C5U08zM/NzmyuhiF2Tg33gy
lEctkrx28ovhbErR5QXrBaRRp0IVQUJTSkEnRz3WmxJg56vPD+F/zHvi/68oBlpBvA3M3tSYIpLO
5AEb4KZ1ViTg4sXuwutnvqr39a4ZKVBzROcWuuDOTPiSJKNi/hHQs/Q20Y2DNqdVTs15Bg1wYAdU
aH9xJ52Z70caYN1a9lzXs/0yaSESnxAcdzILnjNO1WCBe5yULPfBkIk4+DylBkPcL8AWdgrIe7tX
VYkcaJ2CvU5keS6hhamrjTylE23i50YTR6H3nnv6prw6/Pmw2d3Eg4YzAlVhYCRFR16o4o2OzQFF
GMVrfFHcJV8TK0Bv2kGD64Fm4Hn0y4daie5wwm9cD9OqxadeOgsaww8DBeSyxsUqe/Qh1PwcwIbT
DvcoXYFpMWFmxl8dkOTCMudXA/Oyk+nhZT2vcYOxXWCBiAtioAHGPlnW8/E24/VdjXiyPbRHvbbs
icZ/0q8HBlt7hUcwcFnccY7IMAyKeCMVOzlxIiu8jD5P3HAMDmbUvNlSlynO62BJxa82D0MdpfNY
SSsaaeXH9bhuFWkgrhzrQ7m88Cj+B6QukQX9uTtishydwyITTvOLgkmDV6ZadQtSs7wK2z+tzShF
z4zjYcp6PpRrhnaZAfTzUqo3uvXUdJuY6O1MeH/hVjdUQxgea+Pw7yP9CPCSP5ieiqoG6GEAjTtI
odJOSteloGxG4QQxSVhp7UpsTPgriie+P1CL3vRrGtMF7M2lZD0JWB0xau36YRkdRQ0fmSH8o76n
qrMSjWoXI/MceHHOEOCwJ6Uu1SMEs8Emc96jGMBBq8isVPxHP8Rm4iJSVEId0PIU/GFEugll8P9T
o+q2l+38k6tTLbRoczFr+c7O36tkDc4E/lwKtfs7yS4anj9KWLolMEJ6I8TacqgIKgm0zrYWUK2K
DJiwep7UKOiOryhYSabwa5cwHb8DhkVJRQQLTUxuH/UWec7UwqUFCf9twnQvo5zXXtEals01CHxa
tvRlrhLGvuHEvancPxxMBG+j2tIIRMMcQQ1fPwA8sETq1IasmmgQilpszk/+AhaWJiVBSgHpTCHz
CC9KaG1Y6Ss2pLGvcycJS/yr72M+j5rzrzc9wK0FGk3cyz+l2M5BpSrIa64CZbW1dJV7X9H0MKv5
68/bkl0Q4i71WFJAJM3xVmqah7/19U0gCKG4fak+REC1Os5A+tUhwyXSjcretoOiFoaHxT6ZxPqn
DIqlqP9wSnFY5lxSoSxhx4kXNwYeZuL6lKB6rU22vfh5mfuf+EXaBO/gM7HWo9khROTmVrWiEo5P
I5t8PAyw6hezwuTFHr6tqqfRibzbtXGzEj08Lm2l1U3i3ZGr0Vpr9zOj1dHp9wpw4ceE1FrA2lWf
VIqkdeLcuoFs9W5R0kdqcgEFm+iOQto6FAVwP6agDxf2Mcx9FoAsxPJeuanQC8h4uLY4KwWvlte0
pto71Nr6N9Bij7vsnQosirovbNhq1cN++I4U7vOW2U5ktxdWwKjLK6d9kBGeGFrvMegaVriNdBDf
ICqezzO4p5Dgl8N+1N60AAk5xu3nqHestU5UdnSufgjyGdP3Jth7hszklPf+AjcckcFmFO3arJfq
m9K9cDkdNJQuDSeXfO5UgpbJYCzKCt2hxyG6yoodEu+73KnjHVv6Cl1MqaIIzpbK81BIjQ3jnRBZ
o/+hnEKBQAPDzYR0w0xG6fKH1wqntwURSJE+X7R0J48PcA0Qg8uIATdYYeXP5X2U36otvJjqeJWr
rDWvm0GuRowD7BH/uRr9zuMAAaEBsChNqVbauJvGwbuhffGzBaKTeB1InOrwcZEcHxFSukAf//Jn
K5Td0ELdv9NWvFwPySqAJSGZf6dIYk0e4w+MODzV0J9eo8O6EErN/loZ7FcaHxgOwMGo0xP5y/Cw
UScttrhJGgiKmXlk7CmFms/aNjQnZzAyYlvZGXl53XSKKhCkgaD0bp36zFTVubzT06SQTS+0U9Y4
BWT/IObASDWb26UGO/lB0DIC2/A5daLU7mYAnv3s5gjmMej5VfEoEqROiCr1iOA1jd1kgjnGa7TT
MCbtHZq7nYSzMdvCsCH7w1MFDqUSylXN4bn/5cs6EX/XNCDF4+ETKYNVLa7axLfWQBE8V2r1my/V
1EODWyrvLKGK4CJfFuwk4nFBws0gyeBKXI9nvAEn/ezuYeToKrt497LtmCGUYARoFht6oaD9aInQ
7JI96vsETa7qfMT4EqEnq6pASAbQcETnu/gZ0Ffv0ck2pMcztw6O/2NHNlXybsG/4RCk8qTZ5Y1z
tf/n83dQKRvZ+k+QkunqIDmm5AwCX1CE5ZvXmNze/+ZIfTPYYWQTYPqelsJKJhqSyFE7uMtKV46d
Hyt9Jje2K0WL2aX1bIanY+auwba3ejejQzugz+Ff0BcH3rRzJHuFSMDJOC6mRhwQGzUyDYr/Qxw6
bNJzcj2rt5TVA92aK53zZqFqUtLclM6xnuqgBL+M9P4lGY0jq6QnW2n0oy1jwFwPguwk924oRYNg
XHPVF3hL5yKzc8es4dUh5hlCR5UqoGTjGbbBNKjlp+qHDKyTMn0wE5JPXN3pwxj5c+P2Jl3upiQN
UQKHKUPl5YbyYfGmQnc4nI425jJE/l7iNouB3P1pRsTtVl2rOtKqmop9s1iJVHdV5CY0YQFdoLJH
DOhUlUIzr7fMAtNcD9gqtfvlgNFQk9BfTkb39TlylR0Fo5Riz4LiWYy3/cK+k3EDBUIBVDg8oUXM
HqhTKM+y5GM+kV7s6dTm4x0vd3ZN6MtzL4FH09q5L/j1EtalzqXqId32FAUH5v53gy7qM/TPQihU
YBtC8e3IWu1ssWPTxEzjXbTS/xNGrUKpTTnkZIg+c0Z6qBUNq6JszaGGfD0K97ke+6USb11dF+nQ
uYsNKYIEAd0RRjUELO3b29wzOOT90BesmZtcLAr6Dqk+0ajcdVXdUcgjzyxyzkFJD/lCEBnze6A9
q8GTziTWEyjpFE2vkzYtavpU3XywXU3IYPUn5izwt3W0lBrCU3CU3xgfepbiKw2l3PrpMQxqwdVy
g7wKS+Kozvq5R5zudtVgDP6aU3mH/lZhZ3TR7hLMeG016qmD1SS/ZPgskzisnOgPntIvxKv43RWu
hpVWK5fXxLZP3MOyV0O2DAfStVnuB2ZtvANwb+0ZwUiqCEnppHLvMfUQchp9uavzKSYq1irmvtUC
cvzcGFCSvhnu5uroGYS4LY5KVL4QQnuWzb2StLJfWhavBNdIGONgpXibDuy5yNSUNyyjN00ypJq+
P7rAdCXxOFLCb1VpGap2rqSTWAKGGSe7ZGvv8d0QA7NYGAJ/NK1uECQKAfJl6AvYonQ3/PXi0a0Y
I5vQQYTTqlvCnZl7OmekKZJ57jMU5+SE2HrIK8vbJoOVeoJCGjl0JMu1wzLKsPDFwq5j1TNhzu5T
DD/6FvrCvogi3Hd4KrUYxKSq6Hrgz9wFclmHxRQbgc0PbTPveBN8PDtaE1Ab31j01VZ9NRiF+Rsg
h8UDDwMeAsl8i/58K43iSWMa+W4eVkq+atPFREv4zs70Ur1aWeeRsmLroVUmkei6ZhsE41K9mqci
xq5rQ3jvvW5L9CtNNoZhwcu6wuuwPPmADNp2TD+XCcUcsvjwrjyG7DfKgKXKrNG5USl1GVQ/QRgj
eFQ0fas8oB0QlisphCYKr4g34peissrKzYKaJoGQOazR7EcXnJowijiN2XKduzCcCNHgNEtXsGVE
vWMFbN2bSdpAxDjGqi5Z1V1wNs6o1dGRj4lHbklpbArLuFIjVGHNSFclqVlgOUg373nU34Tkk082
yStUBIpvGIhLmauMOOhzm2SQuGb+5sVJCR8VWBAiryJCy/XAkqA1pQOFjb+hY0QW38aD1Ayu/A/w
TDNamLJVI2gXIwuLaViSEcC0ZthDZJS2ZqRcTKzxClgan+86teOuRko1d21RgXUnSf7SDis98exy
PjXVUztyeZSRcdh2BQXAbYmSUMGK1hIcAIUBXJzlGItip2ScuNdov3/XTcYDmLeijbcrQoIS8R56
nK8E++4MALYAAOrQCTK3v1vmQLQwNSuKrPVHvurOC+LE2/TeFbG0RsyjlS+UnQ9SDlrze7RKzxKY
uMRV+NA1tNkaVy7SDKbHfoS0Zqkw3LK5ACWCM0aMRJ6XBSRD6KJfXcu8SdpsEoESHELyPgRfuun/
GkeN3X9R6fJ1+93CE9s67aHYo/AKuFZw0g5/LeHsXS/yiRM1TQ7MXAJs9/VSr75NOGZGH/vZ3NRz
byaWkxJ4rShtXiTHIIMqcF+MuTVq12VYjiF5BIWCXoEUUO2/UQLyIpjk9P+KAYow34RJctqfQKR3
dnp7odkHhmnF66zAbZ4Y1+5tw6A4lQ3AUQ27AQQlNyvsBlFkOpmvxn34LR4TT9ORckgXHUKXRGwZ
X5HBEoZOZ96/kUYOs+joHb5usw8r/YP0CEh9wrSRMcqsCs/uNJ8myRXevXzf6879PIynr3s25q7p
BPZCg5TLx73zVhhSkacuzUBk9tGonq9ax5z2v4UtbNAnHEjGh06JY7i61bMTNTv5arbHC04VTH0x
Z5AA4AJu/oX8cYkyfQgboPF8INdMRL6ZMhnJ6nJLURRSWB0lm9P3AbSgMJ5x5sxwVPTBke3DqCKm
LB/x4T65WWGjJqKoOHfiyd7C4L42Wlc+DXTdsShr+S8bCGw1T827a4hOSQQnPwHCZBUfC9CcsE0l
61SwhhIGo+Nt0MQdMewPos1yGPiX46COc5Llxc32HPxAmactu3DwU8wPoq+Z38MK/nuI36k9Lo5s
eteOfiCJeFeEhrDFbFVUEjW/tgRrPQ4PaTOj7lMdh6eM85x2//B4NOc+MgBOiIp5ZVk/isAjhOMG
SAL+XsvqIyLAR3vQAvUumPjlZS6lQ94IL1UEuauWFIl7tf5zqjpqcnYxsAVcYRYSQ6fc6CcWyJNY
nQ2GBW2BYxCyzoD4LwQxtwNdh6M88mizQuE/a8zgvcmZV17UIBmQhVoY1tgjigrUwZbQDL9gTba6
N2+PY0pKktAFI4yGwy6y3UR5PKailJpzqG+PpT/kvpmKdlBma75AAbJY3or4c7jiloKdvGkedY3t
bgSCkOmDWGUURCT4lDhaOJnrVTPCEezPAexpBEEkQp0mCOKDfY0WmRgw3+KFv1+K9uu7DpfPemCo
RsynVAsmZDr8eoGpKSCs31oISa+X+rCNv+vJmC7gbsRoHml2cTkAzzYV7ZB0boZJGUMdrl26DQ/B
2vtSZfWng+tHAiY9X9CXYBSyTpc2BEYaoczVItDwcF/hdBwKUOlaPuwOaaVypoQqVwdkMcQQ1mn/
nOXiSimfRqVqUEj/qO5WRPFtdMnfm3qTw6oIV5dcwmbxHMICFTFE2ymLqGiDerjtSmBH0MOkzDXH
3rwi0OGmwoVrEkY/nKFdUlBit4nVoMZsV6XPPTcLYoALkv1zuG3KrMQoJcdGRCljVzgz2AS7MT/R
a3FiMUXfDXjhFEhgg/Hy+Ug0YnLAgbj7jVEfpTTxNwQVpboPfYz41MRFsM9iCetJGFRmWLvGd3Qt
q+g2xw7kE5QHS2NyOzBl9oIJeAPaBzxIhWW5F4/ONUMdpvTsBhkYRRDDq/XtK9BaM8sVzT1robAS
0xfAm3e5wT5uHGHH/UmOxYAilD9M4Yure+u9f2v1XpmCgGbGkElmtWfRN2gVrrBUE9m/fwLrjxId
I/y7QnGy93Odi8V3EC5gP5J61+57DH5OeVZqb81qtCVigQo5V8d0iuY3s+geQRjoKS1z8aizC5nk
YgKZAwOMQcokXd1f8DrmNsOUve53GFrMno+bqWRCFFazM+JJYKyqEnEZqyNzOHQaUjv51tpCdRGL
PnQNIA2beDCchCdzYW0+1fzVqQZdrLVG3KLU1RuDor26H+8LNaLC+EpZriU1SRQSaOJu4RdTPr5x
bYnL25VwKpxQEyRaHS24YSVDBOkjDYJjCpolYI5G7MGDFEKh03LSgWoTOuJB2FHPrYJnjjAcwEZk
Ay0BI43UL6W+fmmAEYK1grTu//n18pWsilhRCrdZKAuEh+gt0V/R5TPE8quMyQBwulyRZhF8UEcE
BV7VONmMfvCg+ZACvf5csxwahEj5RR0hcqWGchEvkZKVy2GDlT2OazoYhvE59lQUMhFyT9qVB2IE
9INZNEwfFr/z4Tu9DofH1J5xRnofIwITcNEGBcs4ANemnR2yirifY+QAwudcw6QK492Mw4mQRns4
gZOC3rzYRuSw5RIyyJsAQ6mfRw2e7tE6jx2E19BuzjU9j3exZcWoeMpS5Rv6soQiDLxxtdBDEdKi
YzU4v8O3c54SPUXnZ1rTsYJIAFoVb08xfIvN08HxSwxzZWQbkg5EZSQRcXvti5ChxNnWqz88TnRs
iKt2OWZ3BNi2/XI5BzoxDqJmNaNXDehv+L/+R2NCcQAJ+ls2lki/csQ2767ARBNKMMHYoHY6ov4M
1Tp/rKWaPD5gX28akuqsBOXAXyUo4v9SgiBjjLRABm/qNePEs9zT48Wt71Wi6BbAYilhG4XbxscL
+rgBh8gfBm7d5nMszWADX9mA2wJ5JfDeyLsYQkudojXtQGGPUkvazS2pNHg0WYizW8wTHULwBk4G
Eizf4oEwbzn92KbCdgkILRSmi4T9XXWMFL3IbaMY/sXgIbAYSlwTFXxwSpGi602+JgOz+3b8HL5V
D/UCpAVKb9lyQq5Xw+S8CPwk56jh07UA+o9YTHIieJ3b/+gJxXkBOm9rrmUYGPwT5Jr1euj8v9MI
OpdzbsMjNBR5xSAN+/l0rhFaQ9r/CfDfqyRESLsEHo6eMW6Aj92R930uUC91PlKWcuHwxKxrFV6I
OsmVHUIzw2KtejGFI6BpTqVQWmAY+ajK3i6wVjH2KteF+G7hESGEf3LFC/+GvCnK8hcTSZuAtDSB
eR2udE2FQyDurelMMc/AFL+b5jgq2TUzqBcum3NtPXiEfrktRnhZJF3zgH9+tFuLL9USRzAiVyYz
57xy7fJO08lhn3dnTfJKq+kKXDyVzNkqGAP6Rx7Mcum3/DCBsf/Xv2kC9Px9OabhqGMY83vfTHik
w9Ad6GJOsVSzpMq2ZvxB0zvosP/bWrzz36uVWiDC7f+69ieX0TIXpk7lkaHbFh9fgjMBkifiRpHq
/diIjJ4uDTESVfhON4kuURgg93RJH4+LqGwh+1C3Ax9nkd4U5tWwpEq2MtiugYJVwwvQN1092+Ge
NJvFVZxh9MJ+yW+EFNrGtxv5xDYgPzLDXqGuSRPWETi7+K9zm3hwjfK9k69pUnQ9GAauR4UW5e7Y
xh+WcMBSmTGinH3DjIMR9ASHniYlVYyiwkbGh+AJnhdWtInHna8ogn0QdlW+6uwu8iHQHo3tJWDW
glZQSMHDBceQoSowz5p9gdh1xGXs9cHAvPulmPr9oATfl5O6WoDVA6jTy0MJQ9l50fsaRpNuQOVz
39lZofIM4nxk+57ujDkG+2H9MoWq32SxLtCnFwkD74VkDoxotLrhjfPKKorL2XtuGzul0pAUKLuj
KcS9XqY/jUHKf1XF6WLKaSidJzulRUYd0gf+r+I55hEyPMLscktskgUoDsLiyDjlwpXYG8RrprJA
S+uLvhMkfjTcUzw2DflnOhtVP1o8Jbv4lJRKdb1ftDqF4wBzPZWortn9hxKqkZEVsiI+tsRn7XwC
HN5QKWmkf2juMcbGkk90MWDq6eH2hp1VeFe+TnjbrEiXzcnxHBqLPPspRhcjiY1wJ7XdI6m8xGyw
TiwNXDWoZ1yjUWNZ9Rosfsk8k7mq0dHh1LeIoEdLMvsefIpiVT2tgPas8T6GX1AuURinvBtg8zLK
Vn2BSEjxPQZBECYuWwaBDl1ODLpJIeufe3Y8k6dfrG0rrZYADAXcs0KCL5KNXlYOO5R+ikxol9xW
ZvH9eAyFJxizz/CwqakAqbWCu5/jqazuo418n5e6BRD9o1IVH+N/BXGWZEBkEYnQTRNcIUU0PGn0
Sg5GwfgxslhqlT/VoLLVSIp9iZrfs5etz4DQZArizKIWyxLf0r6uifpGSCTbgtrUiFvA7+0tImFj
ycPCLFdbqazTnpCmJC/bYx9QXOXuktdbzN6ueFFtudea9fqcaj4mAp45vokB4TZov9SbkChZZMpY
lZysUspnmUPptmDnVi5ShDeLXDMB21kHhsnBso2HwxObrGtqQmsqJ2Pf0JdRThoMkH4S4b3b4ukg
AFUVS5hJiui0dNEHDkYiIdznmF8AkWKA3MbGHlZjoLOZci0lPvraAQ2knZMCXwKuCpgj6P+W7/wW
y2IHKcs5Kw87WgDmkZy1YqJCHeIjn3qVhEe/Qn5tXkg5Gl2zsj2kkhzXI0eQvZTuezQtKNPZ0gID
z8BcAQnI8onRujpxmyRsLy7IhNZbIYlQhqOnFaW1R0ezWdigF+JZcdfEUH8pKvOUyZb+fhFG6QP/
OdLHWkfymjvHLB4NODQc4vjDyCNAKiTbqR5XRYeCPAPxKxoVEtz3wPISV0D8LOiUPa73bCpMYPI2
JTuVAFAW5PLseT/lqfcI9wC3UU+K5xUK9ci+DzjZwJDQoBw26WLkpmgNNHuRg0vpE68ZfPywdDc3
bwWynKqci8Lc080eHIN2s+sXMPUOLnjfeXTSsR38xMPnvwWrY5VfXkGoqLUwBXGLjBvhc5WQEPIp
ddU6qiqZn2Z+QHAVLMK6dzjG6CbhSQoJBu1pdDPKAisSRbRQpZqNDR37rbFudwKlIySj8HuV8lrH
RAVHrsJg4yiM5JKMmoG3gxzvA6KixrhEaXoVJpaVRiQXyEcjmIsF083twDnEBCLZGM+3nghsAeTK
zMrgX7X/d7qN8MXm7A1y1PYqSXt3qKdXwTvOvdp/l/XFkNa7y52xaefeahj/E4ghA63fbA3hWo9m
5jOQKuVEfNRX8mAYDjhuD+t2nOv7wn7hGrct0QkZff9Y7WPd0gy4/BKI/L+oaquXd4hxVjdxaGZ+
sAOI63jFmheRUAF3Vr3AvYM6NLTUbNmJJEW8AY/jLL2OmOyO0bb3LRF50QxsE+Oychb/UaqNPVI+
J7kc74YczBc7zfSrJrRyXofbB8bTO9u8fCUci0vYvdE/7jc1vV4sIXPOhXFtY7FS1KVwed7WM9b+
qYXlr3njV9jql9NxMII5fwNlrmyGsX1B7fuTP2VO5TUNr5AyEORk9ALFgB8CSpAkjNPSqSfyH5gM
JI7KOl9cf9uYAvR9QlHGjrKb6UKtmOYqOp7P7AlGBeZ7C1D0NfJH9CMILWqbDJPXdhhnBRxCc653
WNPnmYsYlUT0eWQRT024Z0AcKPNTDCAOcWZ+A/FqwvWwXD3w1ah0sZTjS0X9eDV79RUKRBtAaKEQ
JPmHdiHZxw/SqHz/jDhL5/PzEk3V9NcK/EUrLuAr0bbaXEe8AktjbidncN81HVNYZnOn6rCkOSDu
gtgGSuSBYa8k/hRZ5ESsSavzra1nIBNlGiUemWYcPFeAFPRjT3N8W/4Ty1C87cJ7XM21poD0aWxg
wEogf9A8Frldze6Aj4oaI+RAVuA0wrjsE/L4i41caAE646RepjtZcyaMlTuALnAAt7IZfzmRpobQ
/1f574gUhm4BULNlUfq+hvUXk0kEM8hoGgYQo9FoBGFcYHnSFwqNwI4NR1eCDrcQPXz5c3D/3527
Oc0URSubQL5sjjnowo630EXmx0dBER49ZrGgRvFesFYPvY7pObR6KAkPK0dFhdL3faxJx4tCMebu
RsHBMTi7ojPuzypLx4vP0ScioOGnHTIthNuSbAo6I9gHdefBQwCRVsFtYYOc3Pyl7GhskFqftHdc
6UnOc9X4xVHdJQYKFFX7m2hZmR0M22y+24GhlamrLAMMD4TyFc/2DAI7o6EfhSZ/EWjGLGCUlv7w
Aiji3t/Y3uZb7AH0dfhn9ncsYKTmcskwwldDuafSwnmFH8nlQwAEDfK5GlG5GXSLL6OFLMRyMoeb
fgznyQMsuSv6iVlsk7R6VCAxBp0iCEJRkH4bCddCA3q25s0CA49XQcqrQbmtWFjPgM8C6Gy2YkBb
vpqmmR+9SCb8Uo05IWo0ZgPoO/qfmyYi1Z6Yt1aQpptyZ9+Q+zjDQP+RedXhNANw/GYCV8ZuX//Q
1Xb7xZvYL1cZlrC+6CKcedAHIkh+lcUDCSDR91CxiGIwsetPlLdCfBx+aVMsqakgMC/hw1J+Ue7p
XOZguDsiUw3HDr6QsdaMACNHur/Oo3ip/EuoQvBkexRLvPAtabbWpDHZkibYePFMMNaePEcIrSkY
vFCiieaohBO0W/qz0zJCqh/RikGevRwABkbmOAED2zetJaHSHFVQuG6HNZ7x+0VyihKRRxBpL1mb
lA68tvm8vkK2T8DqiNTs0XRAQX2G+Xe6LvCwgL398IY5JdikSzCzE1y1mTLLmOw5XjLs82WyCTHf
W9se52DAmriurAvWFX4h10pNVNTMUEdaL4fiP6KDfwTtDOePNoYDP03QSZcBMh/Z1ngTDP07HNhb
a+LZUhBaKmT5U4vUme93TovhVN4c7mBXz/FdSbNHZeys0/SntjZ8sHcVgECK/6ozg8AcKZmF1e8t
gC2LfsBwifUVtymNe5DNVRlRMm9UqWy3vvIby3cTaUaQXnfTp6IFV27IK//K7XuVxsfkCRiACoPs
QsUyy2PQdbFz+MEOs3VQRcXiFuQ9FkKoVnOO7shxC8setr0XpyzvjO1TB2Ref57yxEh8ybQmn+6C
b0FocZrmBoPfkuc/8szkZ81bjSe3f+dLqoRDaIcOEMHv2iW4ob+OS9g61ITle5OzM3LgZKYgCeZm
qfEaLSzwKVkJaNX8GA1r0WCGoGJEVPfx1zjqeUA6Ff+axSfzDjLr7qZInSkNL09v8SLOnz94FDMT
Nvz90GkppdlILOzeQIlZXs00D456JusCQPx59il7ZtFceRVkFBZlOSMKLpWnLvIQwO7YhEhuJhrY
uFDQ+h/dhrfcmXRcI50yK2n66+EEJy+lSn7snpKCXXruMElQLaPU47VhMqDqqVi7pdcfvRYbIeTK
VgIatZ1+z9Vr6XhscYczkIiZ8S6yhQZq4yDeYAFW44KyQuhqUfMYcgSdsJibIrkMn9OCzmvSjBs0
lqUmuDoxSdU8fpHfsJ3Y90zgZ0CDhKzR6o7onkW+kQYlj9EsHC5aFHTbgAaEnDWo/jNnvriGXELh
bh2pHPW8eCFWpm6EcmnCBNSL+sYcoJsHIa62VZWPGLN+xa/YGf9NfYqAO8OHw7FJ44DOjytYtHE+
eAqSUtAew4mfpM/0etOF73J81qUm48eJfAmE6YiitvGecKcejbpQDJDSstTEnxL+fj/ccp0ct0PH
qOYXBViIOXBBoI7G0MO0jhBW+OtXijvcqFx58H3LWNmmEtE13bDvAlsUtk4n03LxLbKypqWhf759
JTjr8d7jUINpOAs+4P0gtQnH/FW2opv7oGhSRskSMI0HXOiqFBc+vbpATcNMOLEjWvWvrGRClRL8
0bpz7XZssRJV/tHIThm0n23rCeNUYSH5Tm/eQY75jgG6vG2IWVG4X0r7Q+JHE/pIBSLS1GtYXSJC
gH9yDSrOZkot307aGPcPUXwGB5L9F3C1ez434sYp1NJv2H96+W/a+kP0uuE+/mFWWbNZzXoKR851
Q8ie0dejq173Fb+qnz0lFMQ2pbq+aBIxPaWhDCF5RG/4tF2fo+PlcS3CfVVng05PayN4F4KYWT0A
GavS3iqGwB5rlZCobrPYtiP6DjAqdOPFGwdKW67qYbgHdObI5ozNS+y1G6Q+K5uPhVIMpdf1LYSk
DYzIB2BuogckaeyWg2cbnTcFVf4Mujjz4T9HVHbbKC5bADvOfJYowlNgHDkc9uBnCGMA017lLnrL
mw7DKa4sdoyxkFXKkrEnOwwyGib5CU396Ib7Bk/147QaFa9Nr1AtlJlHgxyebbGMKYf0J57EXR+h
bt8hagWH+t0b2bfBN6N4O9kgaU/735wlZKVuO9dFphMT7LPlv5miYI+Eo6MjML+olvAc1qWdidsv
gnVmf3nVE8+zBAQK9rRZtPDhekqVYkGru6+U7t5Q6LQ6HhZophxv7SEfikhPFIxE2gvQdmAwi0pq
YgqxlVqIH57kPTpT2WZly08wAX5t+kgEKWsh4KLBwnr2n4BdIPtT8ycO8JZeSjBjGWUazPecvhhM
s/T+aDZilwZJbX2Jv35HSNEB0nTPJzCKTIa7CdnCNRt5CfVqrEGaa265mN6kpGXc3ZyYTMY1yzjN
hmhlKONcNs4+wY+9MYNyA1R4h818zEW3PXHvGxNbr0mxwDxwYF9UOnHpMkpOBy4lniYhZTlqxV6t
jiv4SsmeHD8hNWsNWvsVr3rLAtxmRkQ5JH9ZaOOJBj6Bf9vbdgSMeIeB9drGAk7DolZV5IYRMh0G
Lyz6H/I8tIaYGWpx+vMGarE8v/AJDBOhJVDtU12U8GYmaWKueaIxqw/LkTpzzWpbqsLs4V1KXzSi
af4VPzpMG1TOn2tcDv6dAaIMQoTthSmg1FLMgSZUYMH24s7rpZNCc1+mT/waA54SrrDrExR8jYNw
7Jzn1h9+VavMB36CL+TWe0dDcm91nTuXnvkJPYOWwQuN/AaIBKbnEtnbOUs9k1GFuOvkmSZnhFBJ
t4aZFsJ5+cjH851V1N8CtaQVNyL4mMBJsfp990ak256i7/N1KrQfWRtuevdxChyA7zGOzcE1QGiU
hrzbphQWmw3KJIfce8+wyYxz0JodPZsCxaNs+jFURms2UcGB7diLm4wYOhAmqsMUyieevYUKmuJa
dyl5HZ2yWXtiFqIhoRQcnGD+yF5zs12f5NqYmObo0rzaWcAMDNnYuqBdokluw8UgXuJQQZOyVDDR
sLblPGvq79FYzeknh3uQPQXN9dmqxfjjXuAXU82zfzedI/PeQ3K38Y0C1nmkM5H95mdwwiK19DXS
KIvEhkKiHLMC8EiRf2Zw9kuOe1rsLsGb0zRXsC++Q9KUsRSzQlI6QGQlYM2EZ1PrxdWx+QxpEiLA
CW1dpxCbFIg/hZIZwOs+Hjx5woMtrMZCI4Pfxp3onOZPLmKl6leQwB6Ojh2HMLhE15qNHdrtpczG
3DE8EDmkXv/pjHPgSFxZ67O2y9Ew5qgt8UMe9l6+4rSYZ6NpVSBY+SBqdaHCj5YBvJlsf8oZtqbd
ckH/5DcGIrraMB9x0juK9iSf6xUTi1HdA8eLdjp5IWmhun2IgpXX4+GxM6JfzVmg9BtTltSH8K/R
N5aPDY3KC3038AlNydGoPACVrr1clntf/EIY/l0bt6bfdv8TseKBaSu/Yji0WcDgsvMsIZexanX6
/Hj1H8E0/D0b2zwADElrcj96FjxY1k1fweFS/SQOtB6hs11vWOzuaCPyW1YL/RNZ8miKA3Iywx5g
JfpPLmIwUH6+lhF5gWr/+TUoP67OF75iqL5i0Or0q6okjnw687AVCxzXmAg/pZwUgz0WZZ0tH87U
eUamTt+ZrkjyRvpAsvd/0CVT8Gvr9M1ZHUKp4aJH5MWvr8gvc/MOeQUPpTzoP5iH8Y/6ONgk4jIt
T7IN+7RxAKdF6nXn82LK8uF5HXMekxZ+hooJLLT5KZL5Uct5o7yLrWXhXrCAkX9kxLQSvpbQxmRN
0yoiJHTPfosiZcRCM1IxE+HO0sJeDRnTl7chl+toR1HDpO+9VSD7jzZNysi9NdwhRfuZNGJgmBFg
fOzHyKo4EB0vsaI6cr3uGWr5PCP2hd57CEh0wMvpLXVa3M6Gx79nGbioVkHXhVVbiZx8I74biI96
l8VgBCahwjibXr6aP4Gh9vdDUI/9HpV42kNISMVUQW425v/S/Ux0jC0W4uUwY2PjEIi4i2q4sLUP
OGpLh+OfEi2yH3FbegQFFXC8GmVx1METUwuKCTGNab6E5GyITXnDNSh8XDWBZ+2rI2CxAejRs7ck
H5uUX8kqWsnlAauBY4Aq8YLaDsNlFtUn70tALCV/DNRoT59yffNoq3BblZIYl9icWVMQA867I7+I
Tqw9QJ4upCGgKwcdYC4g6A2mJTDzIeTQorpzi+ONvHtHf6hLKUYxhSKxBKFOG6+WlooNXau2lSMX
YzVdmYwe/tDe90VjnU9v2F23DnSnRcKTRt2jPzfOuONRY8zFxwITZgSgkpMit75fKt6lW5kXnFlD
GQkCKLxrVIzz64kUGvTCzDloaRLmeQ00oz3BDP0zsGy7cuA5Hv/PXJN+eef0e1dUu5hPkVSF0h15
EN+yVdAFvi9nxDkggLU65QMw2lAVBKls3xnBFygcBIryDW3ulAtIKdH1dOtTFpkmTo5hNsQ+8x5d
TJJs9VKKfX9/lbSRWb/LVSDVpNOY5wxofVVA1i4qC+lu0MtK78HRh6xobz9AnqydGQ0Wg5PpcPS+
PilsVgTQ5+8pBHl2DDX1YbArGbcLAiqJMJ0mUX6oK0HKnYHMbgDJYQi9eUUQuPSUrpW1jZ1y2hIc
TDKd5anZhG/xZACtEBpvt/b+UgWSaHoNlpm8/EsUxysyDxslsfkGmfcYZLEiGiUNeNjzGPMhGum8
n6Ng6/HtHrfL700Wk813I8sgEE34EJxih/GdiDGRmI4fiEpYDjbiHyLLsJ/H309KNWGdnVfrrx0M
78+g4e/tno1TRNoKbEIzW7g/HRlEzA3c7+NB65faaJRnYLjirQ/ZM3vWEfTVEh+tyhd367hwafVV
8VKo8OXJplsXtYJJijjHrXlw1w+Bd2qwPbLzT6FChYUeiK6+jM5KILagguuSQk0flJ3A9ozmvtUG
UpjXDi6Y2b/i6w69SaF47JjI2Uj+CA9yXlfTdB2s0JxGOA02iOSNIhqrc36CyoB4iDSqHIhjj0AP
z/22Sw/XBw+YWMKL0B5m68jOfak0LBUmCt+F8BQmCLI3pdSVZ0CD8hEGZ2IwNqU/3LnrTW7dQrVe
uCBHH/mg1P+CnOE4FYND58Fkeu4uA0RTxoKeWibb8ogwWfV8RfJR3FxrjexAegaSjmu2KIv4uMIT
pVgPyD6gbaqPZW/8iY7WiZ5TQfkpjUt9zqs6IHHUmn3k5e6E9jGEN2hoZUy1rbzrvYnzSwfPGhsp
+/FXY2/wFGmbgGgbUx/O+v4Zqipw2NfegbjrxtQjAGACRu7pWKa+fmoYb6Ua8Lf+iFzg1/nUjMPQ
uQ+e6/sz0q5KGhgdttkcIf+UFWEQvSE+oTiRnLXDh/Gin5euVXBCt7mfustv+ADp3Gzi5h0ND452
dTRG0ehFiqz94J/LVc2QAHijc7qWaae95seDbqVslMtV3JyY5NsJd/68WGKjtrsmQi6apoPVfrOR
2AUIvNF7zg4O+WJXj7SaOJ21U0fmPwZdnAvdkE6s8r8Kfq03AjhLzv66hMbE9xdKeZhwdxxMY2D3
J82DQfIJah+cC0AgDh2a/JSFUjvYAW0U2v9kG/atOtmfetfMgwc4EZ621yOZ3aad26qdiGf7Qwqc
FePX0XEv/c2GeuO3BGl5o8ZNv2nrTh7X7qFkpZWAbVCyTbGPb3NCLlTYdPc6kVXx7tsS271xlZy7
BFsE9WiSpB8ZvIZglH2uGH3bvCd3MrYq/dBoQrqcH4C+4Y6XnUcQqwKhs2RHVrUr4pfTIVt0xTWg
GIracXUUZS50FFe0xueceCQKw5OpDEccJcKcR+IQeLEQubhqao6aLYOp4abbhhGs24syNIxyyDgN
Kc+3PNEmQLBMXQhfaN+e0DxEZn9RBHHPPefvZx/mhqQeXGJEB1DIynWADKG2SttbEFTgRqkB1njM
RSrmMirKdqG5s1pCC0Fn51d8gNCnu5ZF12kqUHA7Q4Mo2A4+pD9u4MRWtO/rbnWjhHJxKuWpl1rV
ciNgN/7fsGhE9jghTBsB0gvYOzfEhsB+vIAk1rLNibhQ4+tcPmQTKo+FApR99sTCahqT71usMYeR
g9koMsR6EVM6usdVfVoa0sIY3vy/rUvKXAz5nsZUR94auhyI1QxMw+QfiOmQKja7DYA4EbE2zhW7
gazab/XAjiAEx1HX+oU6ReUpQQ/imgVWu7Nb25opu4PsgjpqRh2+SGGfoHT4ducwiqT6SpqQtV/3
A7SeEbu9hHlBnGtWTBLCibAlomgd6IAtCSPkYBqythGQCXkti+4VlqtvbxqyicDVT87hvarY+d/F
JUUb9HMaszuEybkwcF1JjFj7tJ4zb7s8cp8Z723Z6C8khX1xsWT8hn+eIp+jcVHCvx85v9P6mSCM
arZi3NZj0+xIeuShfiUA/kisl4+O6+9xLr5E3uGEqUrtdfSBlIq3U4s8bEYhq4JVzwueQwLWssYL
s6WzKfrhyMOI4KSzbD8RagR7u0kLObeQPgwp3YwGLUfVfpwsWP/1Q+lyN/yfL1jNmofVxY4hFC9/
dgKN67fBAuO2dyncC3fCHKdM3QKKnvgOdi/b2y7V3BxtJi63bU3HX8FyY3NrnsVa+C0WJC3512rE
A7G8WUKWfa7IhF7AQfL3FZHeJzLDaVWg4dz0c3HFXxmmGyTQ13/WHhFKVPdegOOtVXG8V0YontAW
cStWdS0WyfjHF0Tf6OwAQLg3FXFDfq/U5ZOYfRuJBIz2wqUWFd9dbbGmPM3pk8+XvwJ1eILxcJ4V
nyS9L4dUb13BHlZowE+ixnYOn9Vl1HB/pjwgB2FgYUDXd0ct/z/yPwhQrgf73Zd8/zHq8vqmOKxt
c+XYt11PdzU+xt7GWgT6oxnrpXW+VB6nKDZSQcCDvFTmXybgI+RPAsV8r8vnrbnUox7rXxgEKKT1
2vRjcCs/6bulggzP+/UFa5g/o6V8KF3iLzQXrctNr9a3C9koFDZEUI8idx+oea5GfaKQ/G6Lb+nj
xtZy/oN93a7KGvjiyPt8CqSnqO+ieNO3gisO4ra/Pjl3iKAjE9q353FKgrRd9GkTHEuAMT7JmwT4
/tjvZ5Qkxcpu+JQ56ccLrQ6/LZMwLSsCEUTUUqkYIfbGpxCG2gcYJ8mleXeWjK5bERTlhpfh3zI9
weh3p5eujjU4RtRsw/tqOcmBvxXS7wY1ahQP4iGEr2YXCk/aE/L3BRP3HkRfh6t/eY06IDhanAFR
dXrw8gsGhyWp9W6ZJsd1phjeRxGME+a7v7NTI4QrXcuOJGQ5I6cTiQee/o2Nn03QqcfR15JqKUKr
tQQuX1GLrg0NUCiJSejyIpYRpSzO3gRPyERk/vuHgH4yLxKylxiIlJl31YBVle7qahoJLSq7WZCp
o1j0Lk68DwSHwyUc57sBvGsggtl8IS+n6uCNVPdSmI6FPW3na0b4TlP5ej5k2yvpJ6pk0b0uDBBZ
5mD0iYbjmcGZvKj74SwXvLuLR77n9E6l6BZ77kbAwZmGpeT1Epya0mZJB4NPz34t1M1gyLZ6VnFr
p/RMSt2iMXOYm3g2desxsu1B5ysfYfEgBORHtbOQl6kfjyi0fCIY6cY58dpz+vCJcm2XdasKKp4b
vSEc9gt117bV9Pwm1LeOmU1RWDx3PZAUys1o9cU9WkP7OcYAt4AtEqFfRco7r6okp5qjmAczmpMF
4v0hLKFnXYrmo+4FwPkJFEfUTfgGnA5YOUP+0vXTo/nBAvRIhm/t+jM0jN9SjTnKgA7DsZY5jn+6
i6tYkfTNGjifwljCmyw6sGLAO3DiM3jF1TyaJEEMfBXFY65M/sYp6WTsdFvkbLfMiZY9G8KMrA1s
skT70QIFecSfKbzgbhdfldolfuICUNoFSO95s6xzZr72y7QxBblcigxjpoYNyTjzsQHKBvBtvZM4
Qd+XaKiQJSX9yiGxwBXGbWy2hF6VQDinb6hiB5IxfCaENiGZUdniNifeHMY7ifWNsj7poeM5f1Jv
3hxQSWgAZZ5pJQutvzWoo8SpPZX3mKkgj6ve8dl/ZXzxYhXH6xal5mcrCBVYiDpytTBAyEKjqvH7
EXdaLatvY1F9q4GKu8Rkw3aifztuw65HzaNopaDywtzIjdpLCr+H2SKGgK638jT7ZKxFB5+d+pEp
bMXzHHfa49TcbK1tNQYcm7sUzng7CfwI5gzrVsf0XeOsIUJyCCypVH3MyOZbth3K4WSDMWa09ASS
h5hq3SSldGhYw+45D+gkuhCyk9+Qn6yNof/fJrDZ/8iStL1AzRenuG7bbuODrGX2n4LxDsHuSrqL
UB0f0UKCYnc0QLTXKV05sbT6hoemfA64iEQ0ZI8Di2bNQl+4T/kANeMoWrZRRv2mCK8n81z2HuO/
l4ZHt7MG37mnc/R1AQW2MS5yPUKPD5U3aYGcZE/QtE4KkwQHPVNhFSPxMvb7zuCHn/EkgE5l+FCy
xHaopjnuidmpUhQXwLPIZnqsxec35OJsCUYfguhyQShirENXXA7mINw6ns3RyF5RmEljqrzzD/zQ
3TTeVOybDzNPadnNFO1RFNZdwaSIAE332Pj06wFYecp7mWRgH72r9VL4/i8wuyvc+I4fa5Z3x1k0
zonz1uEislVRsFDA59+q0lImnfaqTA4zEsDqM5yVGwWrI6QDaGLFzi5hGqTnPOqzrEYhIJyya52o
PsPl1njMSDczYSb1rZY/2nju8N+9jMhCxqAtN9LZVSFpgfte5RN85s0cBnn5vjGYCoYsp6j3NHdr
gy/UDR+9pjHQhse86wBamNjcjWlHfTY91Az/uaCUViJ8Y7JaHR6wt+0on46hu/pT68JY5vZqmlgr
X80YzABQujCoSZ5YndJxzVoS/CS6Nk9WW833K037kOWEwj3+SheE6BE7yM0QatJ9BU42eUkmG5Tu
pmdZ56k9UzVqDRnJgcpPPCz7yKxGm0vJLKbrmW/9/wrNWAroZsQotKINt2ZC4zvZ9L0BAkvyhGCO
Pz2t9vMS6FCzpkpaSJcZWm11VZqUK1OmwTu05HEEbDmTd7J5rUCWZWBu1Ncp0xF4YbFqWDPQpS3z
GSCaGrRQ0zt63wxN2QCK5fkuduJL5Vx4QUh/r9Og9A0C9urFGdTMJHxrAEsnwpc+13fWyQy7MdjO
RK+qY6n/RJY+xutb2NkitZNyBNTvLkalElFVeTxrInhVU7jSH/JLklAM/4QkwP6IT/9+GbvvZi1t
5LyOHfejLMzYEdQHVTw+Y7ZtBLYh29KUA7lHWAbh1nxGDBsVU0cXyISFAF6m1fvyzJKTjzF+m4HJ
sqq0/yVeKLgtxQhQGGzoKm3uWxOpKtXlpK8zxrO0UCcWy/jwZ50BAF0KhDQmoGKn7eI9RTP60P8j
M5chHrJLIpiXOrj5DU2WMGpvIxD0OPmOmtOJvYAUUT7A7V5HWbU/Jpp0n4ebySS74h1R0x/x07hp
RfFBhTMNZbcjO31rQYVJeTlHSW4fSEdA2fbIsTbS7Gm4/TlTCVsTlfcijRnIcwPbqe5HuszHPpcz
5GyEUGQsID4nlFf/Sy0dBfW2jA7UXSg64fuSYOctzc4JYovhFjsF3W09q+kXEX568VunDM8v1bD2
pSlAP6B+8CyNNnHJLWXVg6Y9Z9mga3a2HaF20DQZ9XR29jP9vV7xHoSls8rcyannCalOatKnWhA3
SgYQdcT//L1rBenP8FgjKmR8qT4VCmt8wfOUxDTjP7JpSoajaYoHn00boeRJawm++axqOAFbK/N8
iAQ6OIA4MltGpmS5yO2DywdGHQH4IWVvX+16zADO2/V+XuYGWjcuWROuNs4LRSJjx0uH7Esh+5Pw
pkAQG0Drvg7M+vRYhml2JVt1DuKX9c/EH2a07ruO56LBsFy9ffzqYvfACgcmDmX2yn5jYXAx5qad
Tosq1iVCo5AZE9nvBs3AEmxq7bncZVK0WgD91+/Z3kLc0dahf8groPtfDXrVGvEYxRr3lKDryZJF
l6BTUhIj++2LxpLu/yIrF0kPzg1H+yVZV9gFDq49cmdFxxQKY3lfUXPnruCDySHMXG3NAq7/tnUm
kixX4Evz1soGG0MwuNgfxZbr1ucFDCdFNtKUxhkVOGxkTlj1WXho1p00Bewi9zRZXV2gk+ozQ0Z3
ucZb9ho7qohnUtu/pKrIj9QXtFQK2YiCkZIDwHptH7UbmTtTHSRBOdnl/rUZpWQ/PZnablDyZ9kc
2KS7ekZ1xEH+l7w4vj2TAUBt0ukKxxDxj8QfVZULD8mfSUZWwfQTrcMxb5nA2NKFc0PGT47YNmJ4
6/IYlTjiAdyYxyi5biNQnLSYv/52d54e7rfh1q42B0vWlEt93Ck+J9h2SUiiAkaI7MscUgboQqMi
LpfBU+BD1WFplEeVmoJvCv6gPi2SsBRf2Gsb2h+T6MmkWioUzpAnRmkxqb4FeT+4r+EBEKcI6Q+E
AAE9WIYrTFyTCCXIm0SdFJRA/fCiSj1HXqdCcbsEleAt829JSEMmWJI2zqmK5nELlEYzRDEjugUG
OBaTOrROK/SuqnV3UdjxLW5oo5nr23qTv7dmLreavfqs8TaWGgkpQW9WJXZZJj17lsFg3yTJPfuu
pGy2On7gwyZl1wFoX6nXSDxAOqsmFgxEVxnnExtkk25COgx7NDjLthP7FdzCiHlvWMATKRH1Jwcw
Ok0IkqnTujaoHHHBKbHpsG5NnaH3hgggGkq34dLAkw+KMsY5O0gfO0+e7qx/PR9nQ+ZQXL77csNx
+lVyrSp2xwWXP4ywUswDIxkb8N8wm5rvzb4RvwgRuPXwtIpfa4qguYzMeytjcPm8zozgZ2GWuV6u
jf7kP2W9XMrVGi+fccf74+n6CWG0P0obqfFG2wr7yYc8FvM7ZjbUHn9dgT7m4tcO1T1lb8/t43eL
G8YW9fJXGr4BJ9Xet/ElfoPc312a+g7PTHOLxwRb8JCfaIZnDqCZ0gsYu8qhL0tv+SWcX0ggxpf7
+XTC2QOl4NggtTN0xIy7Yg8p0tY+SCtVMMaahq07+m+5alZ5snFjd/3qTluhP2iadVqUFRrwWE7D
xASPHbDYFLEuK+bwkTpxS5PT3L99vrPdkTDV+cbbk3jbid1hHPJkRszT9wVm4EWRZO2G52iZUwcD
+Jk4G5S+9D97/9yhmGEsRcdpLWW2kkXHEbH/sEl1bdislBThDr8nwjvFQF4wfU1/xDRGZ92CzBwj
MduUKHxC0P1N0qS09nef2oQ38XYUfLIb3qZia1ie6O7ucx4sIh7P+ZmiI6wjMBt3pazq5pZB93+9
kbtcGJCmDdMLCYJomscQx1U+4FTFyRtRR5mMGVxhBhpbSWGuwd+0IwZ44kSzBgmRE25arEMBE1D2
upAKs1MYlLyn5wKrq+XlD/V1bDjWfKo96mcmAISVHlLu8xQ0kHqMMcCBqjrb1jApTy9bFz24BIVk
QJyb4qjrauJ9ayR6J2RrDpIgvAjZaKVIg7XfzTSfs912U/6Hk3GSrZUYi32Ek41uEogrLAxR3yP1
ASIh0g9+qR71V+vRyeCV8tkJe3hL5d+iKIjLOuvDTnahXLhllXuQDit7gCNMEok63Yet0fsrAjoJ
fayspJCv++rpKi3r6MkqEqIMF3qozuJzPBtYrB9O1LBnTjfPykh5f7el/O4UeJE0SRGE7n6yfDta
6ZsvQQLOyMyKCygFTJeqcGKzVX/sK7GJIwb8dd9G6ZxHjMyd4wkYzWTERbHcw7kevMW+mn41Wo29
uGJHvFH0efvRem7Rk7EYXXAQkh2p1oSKiq0+uGHLwZ00w3g9iudcF1c/t4z60jDlO6q0VZTUJ35e
z3DP7ihRnPMnALmqyGnJ450lUrKhcoNKOcI6fRsr5L43XqXR+iN7hPA3Vbs2F08QaeJjrjfie7+j
yT1kh7UKU2s/IV9FJv0w/t8yZ/apoA9X2zn14xztiwv+KO+zFys/+dia6za5HPjLc0PCtHf17pYT
uW+oJPKkNuxR57AQsN8rEB9bHVFHegO1v4Zd1uchSKcnmj31cFzz5zs74IzkXdCFd9IH5a6kInXq
yUttqZ8RdM8PMSrUXhzF6FHnfy3JZobNABZ1H+b7C8gh8+zJGFFW+KZ8E3a28/ptk82bdrfDYAV+
pvHEssGi9w2YgFJqiyVK9LSAxf2XBCgLdOhpTCdfQRk2GcC/uQVhLCOvaKUVrOAbQJinx0ZH109c
5rwnlHKPDKg4UaYT240wOPLxu2Qg5RYHKdBSqER+/cnAgRuuxSfkmRwCxzkbJvJGpHwhqxOP41g3
x/Gr2mktvBScULE9T0Ts5BWtf7sytnBrOm/wYZP8ZLIWtDOcRpALZuVYkOn4w+2ax1UelkwevWVz
5e2E2mUkNl40T4DZNMTHUJd1FdSVSTOfOXrxLiOP6sMravjcbWXEl/P0CmVsonsK9yrKHB0aeWqF
zfWcLdYJBCZu+x6vYmuTNBg8uxRRmUf+hHsHP50aX94WbpRwunRaiyIQ1iJrWV4IQd0dCAmCmkAV
wcTYlTH18eBRo6hqytsoAErRs88H+l+5BK2qR1dZJYkdNRFh5swB2FrULHGaWjLwViq4i2M7rINV
NhlBomgREeWhBi2hJYfTOwmp0y0hX8r3tK6YaVqCrD+sM0BMYbBmuUUZDvt3YZ4aa82ZGr4NxhTi
St4FpUPRbsl8428xQypSYyzmU6T7WKGvEU5dRd2gZBHEdHZDHCY4jtNuo6PEoEnHaqdm/8UAXTGx
JPNgtOHV9N4YqqcG33axpPMsXMvDy/+flQzZ4SJVCtVekof7mpOO7b9FDH7M5lu9+NEpiwKOKm1Z
WFQJyUPoNL3HVYDKa7Q2c0Yl0/LMIFj6yz98KHLA+m5ArYzZZtWKC+C92rVLsQ1Dm6CEjNTWKXhF
SzDZZ1xEMtCawqDXESufuJ/UgnSIi5e8L+SvpLyaN2cA9SG8WjShdcDFVamgmkqXy2/ZxhTaUQNG
1GBeHNhvbp19ap3rXIPbUSNNzoGIXO+UeT4hbB/odt3s9EgRif+kzFJlAhkhoffqcPweVvOqOPra
cyj1Wa3fBiOrg8fTOtifg2U+tR/mtXLFKx/Qx7Tb58l6MyANZntseBulOEGy/C21a0LDML+NymdU
YqiXINCLrvrKBCDsDSt4BPAosYMZP8Qvq31mwcc37m3ir1IiO3VpcfcAlHmR8QzmTVVyCgaLBTEB
Wk38kIRZr1YrSo741RKGSopoAgG1CCx1rTPmQLWJPQ+uNzZ8ZRxQaofpcWhvdAfNfcsQnS9jRLEH
NZs/sCWnJ935+32A3VVsHXlEBvSLpgPhooVhfHCdDRvVeInY2+llpy7gib8RqlMWgtWJY5McXK6K
/QkvyKHvBtSoM913AJv6vXehoBZJRSFCMgARl+CFLP7zLjvreTR3dZgj3iwblWbVZvWDTfrtqxur
gPWN/CedZvC2or5pVbNyS9Tl+xTUO+e4xlZovw78mhftLPTjx8LAXJl8BC46eax+Vazd0zPWDiJH
/mZTrdgPUg5arpzAjQ5TWMgFPAtsBJ/5uUijvy/4o2hZlcF1juP4Qx5yjZZTYTsvtvQOsKj51ljh
z2zNttm71m/kRb+z5ncvQRa8QMmYf679H8Q4ANq94QXQSYmdzQLpSvI/ixItjojVIs5NdQi1y6Dj
UsAOpfyotjJzrsZ3o95cuIIXoKgei5GzxjMxivsc/KjMwrtNlFtXWanAs5wyusomkXHQ4Zu9RCyQ
5KDQloODdm5SvYRZa2Zz5Ee1xNKaeqQZh+M8tfxPfn5ugw3jv/CbIPL+q9gcY5VqMAjoxj43ixM+
JptXDHV+ShpzxhylvoDd4hnVyDdAofixLkJxWYkXGWOA22YdtMPjsbHLc4Inm8rHzn6MeEZNZC0X
j5YGlt/rrDkgv/yznVK4IRjlVeiYeWVrhHkLabGUE1//PBFYBMJBDP5J1p+V9d8fWQglMWDFquEC
VQfEx/+FIBzeVXhdEIvfam4OTSY9LBhKrvjW147uBREL/NKwhiy1kirOAk//xKMSlFJDJy8o8/7W
WTLyQPncpG50onH1kpeVMxdkWknrO6m6teaqqyBJnoZKWECVcT38Iu0LkUnypephNfb6TFI1hO9m
8OdTDfocKLrjZCjq7DSXLh8uvPn+dpv67Dojllg11FybJFV4sVMvntByZFxd5A+1JQl68SMnlZ/o
QuGAkgumd5Jhz4U90X6AoaT0WPGafTUd6uA7+efiBx/hQ5ARYu+8hBXAbTTn5BgDhpwnpH3coFI+
Xiw1p9zj+14fbJGtcPLXPRo9MagzUmF8Gp046xhArvIJRH9BP9ilATIshX4zhOcHETu9FBQ8S8Gd
EXKZsbqYHKoYqtAfK6l2mmdiy7IZ28bqqjLoNOvO4nbRtnrH7qZFNZl2Gm4chMBS6s+/Fd0jfmI4
EALKFPPZqK8rSyyDrHU70QR/8MxX21P8z26SoWJx6nUGJsv9k0tZ/0G9RW/IMQi9oJV0S+Kdz8Dh
bI4/gUmorbtOT+WwF9pZRfEBsyjitaeaGGIfnl6m9pe+x5UQPMB6wathuc69IN0KARFdjf7DXMkl
7Uu/VXRh/eQvpdE16F9PYyS13FImtrK5hjcsz/L/ifh3/y5rkyOJlviO4FALCEk1DCTT4moVwa8V
N9RtnCfi5/avwc3DuZK3vKR/O42YUvlT5T/zKDrf9rHtWe1VtM4CyLjXmffewYOcYJaTqH+FvFse
k4zpskHJUGlxtx3h76R0rNFn66sGY1Omf/SHX4F44lN8M6Aa4Pt4KhYLNAu2bElbm4xWYXtwJyq8
bnTHQlQZHV+HFMG6vCinWLx2lSceYD/odI8B9xp5uz1JWo3AhUBsRHPWAX39HL1zJbcNsMDGQ6p5
YCtGDhL6bXzhclyV0sTldNBAl9WVcRQO1FhAII9zjbedVdtKxDZkTY06kYs3A8Mnex1Gg8JE0GVK
wUakG+pFebROKAKhpO8UhLIF3xhvHWAEuFBsBBlLapnW6YzTrvQEFVV9kUS60Sl11Rs0JkKoZdel
Nq+lXBSe9o0kAg63fWFbCn2KVGe70fJ533toBn2sxx8wlPeCnR1qqH0vQ3bJUYeo/xdLHQ65YQnv
mI0SnAByUuPu2pBCAOiPTASKU8SlkUBro2IruPtmQSwjdGxXJwUHZfmTo6GI7bTMRInxXRnIJezP
92TLo8fEKpMyZu+8iO17MHESAy7D9lWvbzIThJabnM0Cey3ozAupl8hqRg04HXqaqEw8HiL34RKK
hfUIBE6e4QUYXeP26xYq5+eRhCrqe3C9sJ32Kfx1KxIzXcMtY8Lz8BhgbhX2veQmhbpd3R7WrhNZ
Z6MnNxeXGmFyEi00VLhnLdR34O1p4AvvtHTOiSBCPgp4N5dm2Yt8Bj3bY6ytBsfEB9aireNVzVbk
752t5SJVEgg/CvLj+tFwnkJkzHofgR0X0lyPzpdjUoT1DKKovt/qkfLNdgxx+aML2p7qr0PD8E3+
xlJOKRidTysdynd35jV0Z0aP+zFbW3hIMayaVhrs2keKYPm7CXUL1nCXeDrvl1dB1/zGI65Ct82O
dbZU9R5m3EAStTn29+FwXOTUBiQ3JA62PpCaBZ+Q1nMQ31YbIW9AtrmO+a90emVQAPKMV2lBV3PN
e9TrTFMliOlUdMOehhEredWgsk3HckdyTWvFPgvjMJGfoBcB2kjwcFmsn/6KxDQ7eHzY0ZW2GdsP
cUGj/l2k8s6VU5KMEwGzD9JEwu3Z8/W9t45lzkmSSKPjPYj6PdHQ+UGjXJyPyT0pcjhEtyFVQKOO
ynD61PbgqpvLXzEbiOf5WVq0yYYvK8Qip6OLefFWX+Lz7BhaTLzI+zk5sRpBwF1QI+aB04suizhg
vaAJeLW1yQhogirJLi4x24n5Tm2+8xbKnPUkWqPuk2lK7icKas8169vWTmTO0CTcB7pW4PXpPc4s
yvSJ3btKKs9riXc6jeBxtyIDd0Tmp2KfSSfniNyYGVhVXlMOXtjRR6cYBW1adTyhFX3PvOwUDIJ9
xHa102i3jobCmY7LtWpd90S2vyesnS56xxamYkhOG9nyuzIGZmArTVhv5QmK7L6heO0eoaUo5vVk
Ir7WmTSgREyCo1MVbmZMks4x0q5sCkLgBpjRvbPkjNVhqJWkyyNUiskWK8egWns5RL1Otq9lGrbZ
B7qKNC2xHiLsSoEI85GCJ0iTpqikJXQt26it0wsXag5JuEDf3AXihzlO8+Vc1OPWiZC5SiDYHXLn
3WpqPkhxyxkl4pPFoO+enc90L2moiD3UKtROQGkNm2ykCXrxlK9Hb2hjK5n7/ugKFioZUIuxqSDn
p2D56mQ+tyH9NTI614CSJ4VteIDhsJvGJCpyZ4PeOmRmlClyqTEJEXTAedazI1QewdwCnBgymW3w
jGFFRC3lsLejIoCTWfDLEotwFjbUtNFAvA/EJ89Xk7MghfajP/SQX6JmHzJ4X7A/3pfVCJ+1TxHC
jCPYGOkGg6r4nnQnZynuY1e1jXHxY87vtLh4PoNOb4UcuMftmYrdtY55olJGQODRYfTMU78C3Amy
Uy5xfvPF4H30RwW5hzHmdQb6Z4NEVirOs42YByVbbOB4gn6cxuiDmUwDC1nVRSDk0elybqwvE3+s
jLsSf+DaYNiuMK512Ea4miTVaUjI6oxya9IukBz3z9z5cCSB4Ok77LanDsJsXLArLT7ppaF6b2ia
ZMJvFpwKeHF2Q0Hm9dWymqhr6HNYou1S1tXxok3ai2JP4VCdWcRkfb6LG+ObIj6kuUlgh2e81Rog
99WYKrHz+lSOcq4tMaMamjbrSiYI9FyZCpw1aslNLcFwfVkxI+7XM2ttfIfsip38//P0+MAG2UWa
Imjirsg5a1/cILSW2QyOH25QzxDwWAhqt1kC3keEUI4OxrE0qezIM/O/rcnfp6jZSp488tXnEt4u
Ib5stgdjoRCAJdpsSUyhJZEYRLqWBIzVButUkPBtJLNKYv3ciHUMZJzvqaPABk7J1VGAXBoHdVYc
FSKxZfakXXvVaSAN6BXeO+Z2afyJ7SKIZuxO+VI9y07QxfQLAcNNpFpdbx+fsaaALTEhEC+DDSwa
s1cPuMqSzWOvFvrQla+bmcMyxLIRsAqWMqmqfSblkN+VMrLXjKsmo09quOuA9SiwT1cmkd4V+SUi
TDqGgaMpLvxRR6Cb+z8HxG2vY0W6eddgD6LVRZwA6nMrwWV0ivDZAl9xjMaSTv6nKLikmvc1YNku
ell5RoFR821KOT3A5Yzt1GaKWO1YCyXnimnfe1CT260nCbeoW4JsCnDj/yRuJ/NsNY/C6uz4ittw
nK/XG9n3I/69oQfDVUAvN4u+1rp4j0brtJACDFiUHgFViO7o0Jvv3W/xn3GPz+v4998FKWsVKZV0
Db/d+phH5z84Az8gP7Tz7hoiFKaK9gWYOmlqOb4oAqE2e09blMlSv0oJaTYVHw9GrsllgM3LYoJE
dqctSz3qaQ+LJms1ZDk5VCQsRw2AHcpxg0aXlGYZJIfbyRnsSTzGmy0EvOUfKxeG8sw5nRNUSvSv
/uMrvBKjofecUGxA7q9+P+xCVtO+kV3Helda4Zis7WkE6MiVe7mKKPX0OYR1hw4V2rj10mnENO69
iESoqBbmSxFIA/3BTOKaBpIeNWsBJqbLOGLG5ftFyAIv3Sv92guqs6+xkOa9lLBzWCF+84IeJ5kh
KSPAnThQ2CBGoYHGKBKpdP6Hs27RfJvoXrHwtqBcx2m3DwGWitqUaAJenoIZy/obuJhoECXnHzLZ
fvlz+Co4OYB9kAAxK9LnA4+RzG8Y/MqCRJvmVYsdtEiOtORQxIOur7SnbES7dK9OpVTFCWUN+qIe
jW6JKVAKZXO7PHQov3xrG0RDtbHu8zpzp34R6WGwYsGxUf0tQF+NcFDPnRqdrl6Qb5pdDs6pjRwc
nhr5RuqyGQXERmRSPUt6eUL7gkPIWQXxn8BM9uuiSkVDmWLFSEg2da4DnfC/+RhSdwCsrLFZfT5v
HyalruCOngOrRPtKYpYYcr/ay3+Er4fMzBM9EHv/X/0rc3YF6qrojOR4ktPPRxg0oY1b0SfG/Bli
skRfVwMPKcQygPei2714Xz0BaSpXN/WH5jH5WzS1JVlOYD5KVRO+0BlTszy57NxS0mOBSfu+JyQe
j+tI0WU9tlSrLAa81LKHHYnzUiY4PKtK8UpK8UXN2kdUJsBeSA+R6FFo1jwS1v8IjFWO53fgNr9N
TbXNhnIxq9bP1El9liw38QwBHdm29YK4SJU5rzqOpFegb6nn5GtH7FxXHCueC77X1E/X1ulZZIGr
vPAeAncKze1LUMKUAT6dO2wvihKHHsAAdY3u9urgZvwmIM2dNp4/JZBIILKnLLsf0cpaIw6xvE2p
WTlXuT6HwkldQOEhRTcqHtk9QXsFGS5FQB3Q/mUafStwKzYfEbsoXfD5J+KlkfMFgjjUZS4OeGrL
R8CxIO9so5A2x50hvYDecCoKa+W6lpFeLnI2Mfl6/DjiyaE07ziUVGI/Um6MQiyOx9uOrfachHsR
tSTQBFLnwz5LWso04BsikjPiTW5IUWi3bUoDP2eUffR95kZ7rlPc35r5qLFrxO57tFXQqV77eWB4
1KPotTeNS9q+N88QHKm6GSe1ZJnVxZeed+RCvEdeXNcV1pVt9ouXeKDmKuxIkqHsvN3WTVhBowAx
cf8e+f4AXJlZHLahk7gwPZpmFonqBt6Tk/mXeBg57mcSbZfsEZkLKMIkZaX8+x35g1/nuhJ8H7if
5POCoLcNzz4w6aNza9E2UVHt4UsO5EFCW3IqtBkjXO38v9BWiPDomlGmH1h/IwhenKlXGcHujfqY
1YKnH7oNy+5cKw3v97ndVN0z6ARuqP+pDjfWg7s7hzvHN1AVUS8cyXCELfmJ1gkp64/pxHCdbhKS
8vDzKlyz/cUa7I8Sdn73rdIqg5xbrIE28d7wDdbLMMVxBsv4Wo04Hdl12HOuRIdTvaU6kx+aqAhR
l8fYiKy3//x9xQXy5ZCpDoXC9zJ+b5SFnx9TY6HPDqes+VxWXAHmBB34KDX72SepvfMxRRF536Vz
K68EZx38IpwcMWusbdKuoZZ6VKo2sR59ksBCeeMZzHM+McIn7tApjGjkH64T2jbxhCBR0RA9B+vW
W6ehCgOVq4bk4vFzW+JZqLfbkI56TBUBGzXMHbHqY8IGEe/tpF7WeA3NdyfukebM4Az0NPKKCL+m
bQmGcRCTqpDHeAvlf7U03bWu3psNFOB9cAm8dhinHWR27N2ZKD9lut49QjFF7O3P0GkQX/Cobr2j
1ubaM7xtgEO87O8aZPFYTWsdAnX70CYFSg1CEi5Ny5qdeRNdRn2e8uCRBmFktEXA0Ce4X6my3s/w
YGtD2Un/ydv/o/d7QlbAWhf1cXgCJT/FcqGPnYrQwNAaD/MiFuM8sliN9+5AiZKBWJaubRlNEg+T
A2uuckc3MP5gyPtKcrrvL1b5QiQo7qlRlBhVaLW/EYVQ2h2GHagshcsJFmfMV3j6j5itGInRigAq
D7GYXcUdYIuA0DX2BIo7xZYO0Ni85O3Wk2qUzW0yKuT6brLFW1lDNyXT+C1XUpEIHrTaO3DCOLei
p0/gs/sTY0TjmP3sPHvTr4s7I7wwNXaXY+tWzJ6cKeIgwhWuIPFJXlk0n8biy/64AGhPXKeKzkdn
cuj5KbfW+NuvVjmXOeBwcwvaKgdWCkigUWLbE0cUTeINmZDcMVJBCIWNwLpZz1xtl0/TIUhvEpqz
BOAWfhFTlDB8/33LIcTEeKKTrFg+f2Wpr3W8dZW9/5KN8x5Q1TNSSXsPrvPXWjlMGwYPvOOJ8+sR
mAsuEBh24xucnPTH/CxYNOeiv2Gkk02Htg9df5we4NAU4pyb0aoN9lFaxr1r24vXHNEJvIsBVF1Z
izMgTU2sc2p7+XdiDNrwlyFnNteWXKqtgqmYcj2hlPKZ6oxDI9mt1ycIsS8JNbAHClOZidIZxi4j
vossM4FbHjNwhqCmW1nwkm/guKgyK5YoSGGatZS7/VhmxyV1s7P4YfhDuVy07b6gwjg+isBfP9+w
qpdSZR9zLzVaPUXtII9fVu8Zk8HHVFYNlzq2XKLLKc4aJypGZlcdaO4rrJDK39KWowkQ+35o6CHj
oqzj6WphGLA31yAqFE1ZCkrAndE6Sw1hicxt3pO9oJAlY+O9A4oPGlg4J7ShQogGOr/9b/k39KyX
B2vFW/V8kZLx1qa0YTcDH25wbs2uwLdNodIvdPiIMwBpJJzNKASwDVb+HittuqVwsowtEQn0OYtS
MO0/s0Rh1B8qbhQNonmR89xOT4q5hWHZasiwE99/32Axis2Nx7sI+hC0ULfeWJBeo2UYcpflUuCp
8VabWq0yoZkP2D7/y4ybV2pURv7amvfgNEAs8W/LI7QlUHGk6YO5e5Ya8vr4RCMryiV/lYdwK0Eo
Fx019RE2eruP1kRzIrhCU511Qz48B8i21IDIDLlbShdDjgDTigoLRolyvHz5350cJjfJvoCehmML
0c7iF4mDdzWxROKX1/IzwfWjxRB7PoMPTenjE4nifrjNxwiML3NU6ws3/sJxiUNSasItJSXYAoMf
Gfd8aMyZOAWokIXN6vm9K67v85ppBZPxAteZDftPx/TDt7bqdDByDx9hSHD5xQ0bWU7P+YbZPr0/
rht5BTTX4XTlXoQLT1R1ATGZWJEiz93bzu8BDZ9uKclssBQDRAN9zYaWT+oODOXer/ftaXEv4Um4
+qleiZnJMilQdlJTON3E1JLuLnqeTsIs/GxW9bY6qgA9AmcywWnIkF4tSSj3mQTn7GkoPPcE63dj
Q/S7GRAHqXQ4IcVkJ+/vxKYY5nPWPJGZQoZaLKmYnDWFwewYPduo1Ri4A4M5uLzZDnXwDOof/m3r
xuCaxOQ6d2TfnSI9t8/5Xlo03hcQFqbl6gtVx8AXgg2/xpzrA/RNr5CX0EriD+f+OpRaBR7V7amK
D47YKFsisgbhOs3DvdCr0DkVw+odwlTkQQIAdZwa9W3J6ZZ8ccTrHzLMrODHYeCP6OV6cHPgunyy
3xJ2MI/z6lykP2Sh6lPc6CzaWIsBwY7GYJxsVCq0FcQCIeoVYX6muam5Z0/Cflt+DlhOFFxPKT9s
3Xp8no8pvU0c04JMMvh5gJYBsOfPpvWgAR8zzEBGDbYtOecp5FXjRIBLqkSZXvFhb+bcIMO6c6Z5
82h4YoDj0pNwaYzrfhrGRks2U24/WKoS/hmAIFrDmUniyRxKV7UFpmb6bM9fVjLbb4QZqAgRGexd
Sj0qo5F3lKMFSaQDUw3orKl8pdgJIYiTRlROmP8TiQ09HxJYrfOeaCs0wmJmPjZ1P9PbWHviEVkH
hXpQDXYeFbnPTiMi4LjP7ReShw3B4tT6p81u2jRi+gyFOraUI0nl1bd5ido8O6jCLFWrQty4MTPT
QMLFGIIqyN4lEUF4S7/HtVAIOLHnF86tp6J97biwgSpDuTY1qSz3MoxCAczozERaN/0AVdQThwiR
cjtMedt5DLEDCoxYyp/Ah0MFZZcVNqv7xJIkuwEZJXVtubScj0pqI7mbnxpfw8rhnYhPRoNqauJ7
emM2+af5utuJVXlyAZDuDny/PpcTdGoWKSQgdv+gLBwOYMe4egnWE344RoN82DCvNgQcv8OxtjXD
7DLpREziDCaSUT35DK2ryP9yDsuIvx++3WZv1sWeYEVn3+ZQwG09foPiBYNXcmE9CzI0EZs5v2Of
5uK49jZdKV19Zy5dC2vsN8vMAk1uUXbz+BDiCaRH4T8JXX5o17s2wy6wVfLiBb2e0ctQ3KMbe5fg
MOkc87T29W+2lsciw8fUQfC8aljXzxL1mMrR3+DtBY3S9lKYzq+srUGWz+m6zPyXjplKeqegj1G2
xSINCpOtrgKqSP86LP2pZo6E1iUye9FuAcqygIg0vPeYCypuvVzGQgUarsUn4pFoOCVJfp2HW04x
fVA+SRvPGe9N277BnHmCdWpnZD72OBvKOhTiniRxqCdZmwuw4YiErtFAMwm2PN0Nku5xPRXaxyFc
OPwdTL65FIjwRxAdwxCMCw7mEwLQee6BwvCc3ll4a6kugYA93AnRKGyr831xjiLgjjKfUtrsQEJ5
1ywSktLhPdIZPN9NQilfc94dB7SmhOl4wAcpoOmYge1QfoFAuilex0SQpznNkIifznIeSPuDfgqb
KwmiYuFRwfRdR8TAM/F6XfjW54z8ismcHr0m/J+cLzOey2L1xtCOuDjDTMoTV0LuuUlreVMMZdgH
DbSDld4gafpnMEQ66IW4M7otprNVpP/2l3wfAjkmIrbrM2smIqZ0DZWotTVQlonWWFmJYodRHFC5
oGGRGub2pksVmdGJnCBD97kQs+0Rf5yGwC4/rCs7O+PuwaXAz1BQCHv4pQQYRUVB4faffqbRn9wE
hYw0J/QOsFyE2W2vZef4831IuPGSN2LT06h67wRB9IzROGSuq3XA9drt61T6NQYzH4rjTonir3Jo
g9me8ofjCXwcDIUOBOunbjNglwi4Kau9y1lx0C14lzV5Wk2DhFNUANsr5zRKi3vFzGLCUBoXXg7n
+qECQHZ+XTYbr1GbAiTbVUxCH5hVzwf3Yz40tdfExzVRNboiF1JWzO0AbFxlPWndifZvr560tH5W
Cj7ZByoZjmKwI/Q2Ku6kz6YWHAPlTZVTGTKS7NTwYHOZwrw1oQ4VkkZDYhKkMvMn4OTvHhx49Xze
/ji0xF0Dcvj926SPeG+paHZVH88YFUovV9nM/1Ba6E1+QXP4ywC31wozZapyrM09vqN195vFygDk
F7689KWvSf5uQmi6hvE7ePSsvUNu+QBctBln580pdErXCyc7ZCy2d43v0d4wMjFgtrlTscEp2quE
tMrWCK9xdQW7g45UJB4L7/Z8j8ifACDEIl/6tF3HvXGXDXN3dPsD2hgXTTD6FMXVrtOvtOANeNK6
M8Aj87P7/cKkRyCCAJLG8Mc/WUlYmMKBss8O3HvnjsvCryjv7IlvwMRmWvUP47sbGtSxzeK8vqPo
95c8PulWSEpWnE7ciVCPQFlU6pXABjFBnwcF8ODN7TcJ5cAMR9zr27KuLAeA4jtS4ZwodXN/aZh/
vbX72riRiurshR3KvA6SNkyjcvvqHddTxweR2rxC6ZXruSzr43JsBdUAIlHnT9jemRIRs7WEVCrz
72zjWQWsxjQy2syz1f8WPmCov4eDgX1stxAZIPCPBAeOyqzz1zTUvK0qYcVz8SSvzQVrnE9aIPvz
JxdbXEeRL/XbLzaFNSFxlxFmI4WZUH2soB6xfMW5c6bQxLPwJDIyma9KKLrp0/La28JUmd1djRuj
A6Nw+GhYSmMnJgnKoop2cXuYL6AldufOXPMGT/zrpwPaNBdyncwJXVW0z/LONMCZr+WLPoaEERGL
s7Tjvf/4e9RUPhAoRuvurX54d+aotPNwaHiHeFuc0sqXjPyTlgFSj/A4djlGFGIzHSJV2yM27dCt
LQdnWSHUzGn1GAu4tvSgmVLmDZlMc4zaCut7y2eupWSY0g0kRdyTt1lw4mUdk8jKRLYoAfInIwQ0
a19Nap9JpzOP6n5sU2TPp/irUXyDRvsKhHvBRWvxA/1dpaleuuO2phuekxWnwRKqzXnI1fyx3Uk5
dKGywZp7BwLM7MLTUvIucEFDBj43ZjeHijlkzM9M+ST1HTUr+CEzb2LvINAD1qnx7C5InL1cyfGI
AtP+O+j4aLXXiACmZ6TmYVeLP/h/Gyag9T+xfk0eWKnQUlUqynAVnjh6F8sGAHjnYyZULexILC7S
fVdwVoM08ncflQR2r1XqtjjP2nu64Cj6Z6X7RLLQ2rxpS6STpLlwyy0GgOz1ZTFW1Ga1I5ceroDs
IP30c5tDqgGp86onweuvGeb2HsARzk9GzLvIafCyn7tCoqCa5LXqWxXlXwX5mUnp12P16ESM3A7r
ojcgFjPnefc6bLDjw0sM3pSIzeh5astJ5vYmpJOABu9Rh57mQxl4VYc2ygtWHVlpi1tvPv1fdUal
vhSCfhtSb32v0AwRx+EeDvMD/cT4C2ejR9xM/M5/wEAh2CHgTjsodIyFH3TXVQVF9BKR2DCnikzl
BdoxriotzHlMRi6pfHJ3AKhLpe4qHVJb1t151FMAKQs/u/mWvazYmtOC0QKhJKk8wwuzEw8qL/Uq
1b14MMiIr4ZD2KNqQTjNQQ2jpqgsG/At3J9V4g3gM6l8D5YtlyMNdJpEDYc4azbkl1TDG26nkw8u
zPR8fZwYHE7fbNKs3MQ5MBG2fQlPS0cjeho9q2WwTM6QYC196NIJdfzbtuk/SCuMDJnJ04C1mBYS
E4Z85iNoMnFLRcFdRy+8OaRcl1PvutxxLq60T2GScKQPt9KH5amnLKHPtw1yShfvP3Jz/hQDh47w
J/HO4djr3io19HVc5bPvDFkhCRq0QXcAYhoP0uG1rIri9tSpB/1ssf7WfkEWgwbM5792Ln3FLoHe
GqfWSqG8Sc2OFdTK5Y8AW84LhOmfBjpM+chtgmSCrVrJ+7yMJbvqMk80UvB3kPI/MEmL8YX7dZ8+
ChXYYgqXmIRPHxxPbC0jK7NPp7lxOyh0xnu/SQRipz4ZS1QjNzRp/nJ3S8y8oai2H2yofcDv++Fm
bTtdVZf8ShMgIGRjJ2irRBnrkNO5AAf97dqi2KEc0zKJ/gLHfHwGaXgga7W25JSZOmmdh9T+McnX
F69RZZOUhRzd6xkrnvV0OKOTPp5q3SPY8euuCV9aytILbzICguc2Z3NNDxtJ0yd0QsLkdMJV11nK
uiGnct9dZ2ZvW0diaB3JCSLDliWOiFSgwr+2nepTtDWdMKylC3sruNbJk++E8c5zhWUFjbErmJRe
wIEFOqm039pETdjTMS0MKmVCqbD0KEZxVWa+zoWPolV4WiykHMH9/9bZS53UxgrpyXl6Va2d2WYD
ZwmOgWXBtNf4ushnZZlBGY/0q6+Tjc8ygMn3UbGajrj3IyWXDC6MDIprE+2dsR81v5s++DP6wQkZ
Cr4RE+VAaIEeIoTMS0LRerk64I7b6tgOYTfoR5oasPtkOYV/pWSeXv66205fqQIk7HNvd+3LIuPZ
p5T9lpiI43M8ALanHyq7izuS284xw2YHkrWvmQXg0FcAIdrDGTYE9klkWKVK/mEnPjIRqCWdvOJS
hClk286kknKFv8nTcE4zkmckpBuGsOC32crIGKv/p7Rp9sKS8hlOZJNC/VI9sUtH/Car7qsPBVNq
MFbj4osvtMR1ad+oH6ns1NTAMKQB+stNYLJY8DNsz6n/h2WQ8kJL4FQVu7i6Mx3EyeAXnKklv956
7QHwQjL5IksZ4lrIWrtlTBXEEHtqje/lqdNITsnumrpoVVDDdhb2Wg1GA8ZTvITGS/dvtbI/lo0G
1mcA4o58figcp0kkYJ03dLmOIkqkuQoBqoWsWHQjSj1BDYYbIRKF7RAvMPgvJ6kO6v8LkUD3mTBR
BeEMUjEr0+iN6IlKScvKEzRNIBP/20XpDP0nhnvy0LAYqkj+XZ5+dLIyNmUjFR2W8+WbcRHSEQjA
3MujKfDoO8+OcnKEHgBbqU05EOFXsH5tkAEn+fMeAPULvLtu+VgTkSoyVFUJuc/B6vjP94Lmt//B
6IhO2DTPXOAXgNoqWlZUo7QkDaxHU6ogHlAb8JpHuEfoZNC85Phe0lwDx+0sbUg+/4lfIFkeRBYb
Og1AqyM7QiRJoEXO2tvk+j4e4iZk8NcZQpu11oA5oKx/+f6p12x1aHfZEBUD9ODo41RXmP00w0OQ
QCeNcvIcV41fR2hNaMq9e6R59X5XtuntIEGd7V9+zLtXsxkL2ZKj8fV1DA/t3qrwCc9NXjwbbfuj
3+GZawzFjROV2dDkgAU7JE+UXvFUhEuv/BQYr80qtbKRhuydMjMaEYVas8M+u5AqMMJlvLYyiVr/
zyQrbzpT2OkqHh4G93V8l9WTOefHClEILkq/eeScEj5AP6whcuHfd/8oUhK34NYNsb8/3OptX+RW
XaAJSMtvvMWamr4SUi4o+EvRVnRJCcLY/2WrZifNZwxKxzHu6dUeNXjPRcHVnV2ybgA1WmKQcAOv
Okyx2L3If6R9GXkWEkymaPus05EBjbBdMnlWliDdNiwafXPzHQb+pbcZXX2mnpi+J0pTaVQ8Yl9y
9Zpb4SmTC+Cug7N+OPWdlYNBlFJFnm2WjqisHY/rWgYVC5Mb1dg5JHMh/InQ5jK2v7cHR0tzfMM1
sH2JH7vNeZ4cFQ9pWfoPquzXZd8ZdVBiWKcq/w6qQ73n0XiAcn/3Ti+H4kKQFDV5C0Uh0oUnq1Pm
FzbVIBy9Z1ZMG8qoWEsCVFDkh9l9m4eq63uBX3znHRBZa6iqLgMM24YLjov5+dz0bnjZRHFVZ8pF
/UCZdY30y80IiC7N0yISQmrGpIsSMpvTcoZrviFNopLCl0/ZNnTw/oN9U4LReB0fz1ExJYMvHhMN
vEizlHFbyxVN72vQ0MnsFQ0/CiIkCgkrgBUoNa4qnUHUCiMrs2ydgYMEEwXAF7MUj2WHev5JUjpF
aDG77bHyqikRRXWbTvYLYKzp9oEhXIna3IuywUiojkAKFnJDxSqFCtgIeApnTGaSE8wM4y4H47uZ
+IIiQsmmyh7pvh4hzDElwtQQDtT9R+OOrfAvLceq0EpsSXy9He2jmx6pwGINwUK2HfJnDFB1NEoN
vBSXVGks+GIEDQufa3IFamPC9iYswtYkItJzPBHZ3UP/EZwb1d0iFW6BTsP+qPs54jpfqC4V/9cq
FruHZDXv4tD3BzlI9IfiUDd5GaToCcSwDhynuqrsxVhp91ieScTT+fqlMj9A17K5xFIzCU4K57Ys
QYESsui0bPDfJzzPwtfCOtzZ2H/f59rr7CDhPakcOqbaabgxp9ZFNU2kfrYxF/VZZ6jc5SQxMTpn
7U6Qk8OWRIBk55Sx/5MP4t3BMmJueDIgRG0G2YfzoXVv96T8kX9JluisEt6Q5TspsJQIzVVHuj8e
ca6ECeezX/L+7DULvv/rvG7hwB3gwJMiX6JkWPNHoLgEKB+k8emxpOtNRvoFw9NsiahM/B6Hooae
kvcLxl8BOeTvWhmgHy/yHbmGY2OI89aVMuckn3EzURKgwKUdYNH57C2d40FHx9s9mLNmtYTp6VPM
VtqMV3vSYCLtTolCsrODWOTQ/xHEZm14gffAbYB0cfXCBn1ZvrYJCCBD0k2DnwUDfZ2kNOBrUG8U
TgaH72p/CYPwo+xQHpvGeoMg6b+m3RtlfWnjlv8T+TDNzwIb+oUVLMc7tv84hPdV/grwM9o6TcDQ
vNcbPp3Tgofg7t/t96lnbnnCsxEx1X+aoSFre0BvcSyf68PhWHwNxAdqwxmJ8fb9jCteg+h7/tn8
hkj+gL/J1t2FqhdliDvTe3AuESVMIjtKO5Vbt1WdWYryd4vF+jR5K0G8jRSawfHkAic9zNuH2VZ+
9MEUI5WvzmSpaVmnVb1DV3s0voLdI555Aw4gENOfunR4/x75wYMSlkkHr7FFq6kmUtWVOQ8ZcEJh
lP/YvdTHHBuVcrUZVHQEYHx+R70Ic8b+zE4Y3iZNfyuFPMtGRT0Pb/REPQNFGmsZpnai5suBn6yd
i8QT1yVshfo3iScSj3B8bDc6D5FiUh5i1a5RAxr/8EZBiM6+kjQTTmPvwsCda0kiUXZQdCzgSDwQ
3lC+X3c6KJXW6Qh2RrURMb+nJQ0o3JZ+7zBiOcheeApTkLFsc1/yzo0s3VfH8m/UDgqS7tqUsUUC
hO8HgFzsCzqkjJoPsxBR0+QL0KY44ZfruydDS5XkV8TwxmlxqdCAtD18eBzmOAnea5v4BJylWudc
9zMN/AjKGqg5WPufUqT8GBxTqKHU1/yoWVMuMZU4CfynleSo73rY7znFrNxC7HSUjmNoVg5B4i+S
tQUO5oqjs5xA9GhIUxUMJlquRouMgMyV5GpXDljTEllieV71DagkBM1Ev+VRyC/CNX66UcHPZ1VM
9BbXySj93eNJma4fYjC5heMCqVi8BChy/goMQw4Nmuqg0HrG7pAlqqXCoK3i/5cIvxp2AhGo6/Wz
a7ksV3qCZ1IkSf/pjW+a6m3C5ArmQa1eqrB4SNpYA1q6OsyC2A8l972LTstWqHCaIn9xPcOF6+JL
N825Ob/xJxLgybhUQCWsoVrkDu2cknTBvHwYoGUWDSSQWHZ8ZD2Z41pRXkyGTQaOPYKJM7YZthzm
EWNPOwbEqhGGSLrp33EMYF7Dx2UP0xLRD6fAqHoMpjhVbDWeA0tRcKhkAoh4vkBzlMxw5ZCJ9yT7
ODVtWWN0oF67Or7Q0p/6Y/aUU2FcTOSG4LCYe+11MV6VbRwUKd9NzApFjwUmrELlSFn0p2+we6EJ
JO9/7hr1xulasXrDHQq63Ae0SIdIJ5RN476J5skRybVSS1Ap5HuouS+SZjaCaNQaYIicABgoWXDf
9GzsN7ovC0UeC7BIyyuWh31Zp1iIaYrAkp8RrKq6FbdnZMLKzPSCWIzXUOdo4Ou7S8eYOqN5F5N6
s6IAl179JWN8jspk6YI0x0sXmJ4Ca04RUO74dtmOV4Lar2XnLMQHaDJyB02bCMc5Vifr5OVZ7jdQ
chYAAefM+Td3Ysk+jRmk8LpVRY18r49LpHJBAA2VJB4m30sraFfgTTZZsO+hN+8J0SQEu0Wpv7rj
neK9yaZKjXJriF2jq/QvJzwivz6uzs8G2HXqV47UTYd+T/Fdqian0JT/jc2IRllrNRotYGTcsyTC
hH7iVMoucugwg0sZusBdV1Rkipj0qEpBRM+Ibxgkn1sUD6r9cfQK9OG/E83O5WjUoXGX15dIu3xn
eVmgEKcyxPi4L6U99IAiQjHF722XNlui4PU6/sII5QrNb2xmcVyaIGXYNNu3JdF6qZWMWFtENbGE
uG5qGUDorlirzUJv1PhOlpEG1tKpYqS6107a8ZwedAsrNx2sMcfL95EEYlji0QxVZi25WSRrs7GE
bV1UM07FjpbabKP/lHvUeGIZCqXeQ7dNFrMOr0rH0QR6Lmk7hsVygz1ui3Vta4M0ew13Q8HNrzy7
iLx1UvzUDto4migNmwBKwsJM/Zfclqet9hSJ5ZQIO61tSr6XImAnhr69/x6+glTbv0hV0MfjYArB
OzRs3EQby3DgZWFOApmc6/r2RUBIY+8XDULM0IqFNJ5WZ9L4ipm8YS17pOi50or9AuqahGgJ+tHh
X0wbtpL6V0S3/veHsaQI6b4/gRRZ0gfXv1Y/9AdQ2rTcRZpliOwO4PkrrMbYVSD4R8+DGPUNBASm
v1uOUiaur9pm46mZ/tEk8iucNkGd5tkBflYajzlPk+DvFx56JuZiWPbwceCLn1REp/HIh2ILr8fs
Ims+S7zQ9rMJBQ2l7xUrTCeS3JlmfHfZIvHxpTMD8ON/YfGCifGbUm/OOcxRr2CMP6ZEYmKBa2n7
LAcnPpG+DrIzhNwlgRmkhrUC9m79HBiFMk1eUHtXuboJkdXP7DpJ8VtOrhVHFejL0Iym8kKBs9QO
LvKBquLNda8FOfwfF/hmc20qH26jDSdGMte6qJZKDNqYem9nkYM992gForWjcG7Dm3QOB3gXRdb8
rlmL8tmNAlf4rwIPg0U1TOQRbe8bcl9gvBksH4B8R0W7fwM85wNfWJCHRECqXLaAQhmgwzwIV4rV
6nn+k2DM6yhtZ6P+r2cQsb769F5O/po7ET1r35kxD2jJcoyYlohZ4HwsCPxrq1XQuOUabNMALpqK
5vrVSlmjQM66yVPfRhW2TeWlEQoZ7kg8OdDefQApj5ZPGbPRFUTMzbKzr/icj0kostDUnVhQ9RBa
4wF6x0klXrGsWo3r8X3Cfd8hmoHgk5RLnhjt3N9JcU0hOYPtMWEihKpiFFC/7c++XlAs5sq3vxG/
YBfdplr/iN5Ljxu7ac+25W6lHwGj64Q3f6EuyeegsX/kx3Z9qFO4R/CPffKYihw5RAyDokkrv57R
cTCwkIDl7X1pKaTlZryuez09RoWH8oQrslevH1NJmyHu4cx7ny7lAJu2kEWPUDPORnISXPLWxKe5
P8X+BwrNaa67x7pYEEcKZz3nh83Ra8ea5JSQ94pDmuT6BR5hAmn6E43abEOhdEyl2UHqY+LBgXr0
n/5Jz/HGeGBhKCXteZaWjWlu3OySqDtkfeeGNzjH2aZa/8BUCA0aejQlP0FMwAcnRInmFZMBc4Np
cvlG41kYyMZ0m2CFOIxlRF5EX8RMYB7tYC6AFUjd2xz4u+SUy0x16xeEh2WbS4ow4PpHif5WeUHm
hHevm2CdbH3GTe2I/04aBbiBaFqMVcTFjlAFeJxdjkt7a4pqe+Bat9LRgbMo46C8wX4uVM91QRDD
nE84M6m4T3gbdS00v1xIu7LAdMJ3/h0/DPGBL5PyPuTfgJKL29nqRzxvCbSjXM/+2gBxlFDlvYAS
ItQgftTESRTOl74fzfsDHsCTOF6ciHcvC0Wn4PL2F6PdSwDDT7yF7YOKqhZKlhsSU/rkZL7aDJrf
/uFMgzjYMtIrzDlng30eVv6Ln4I8k2swOSRrcs3M0orALh98ajL6SgGS23Ix2pj0+DLS0tw6S5vg
pjZrP3lXRmyhGrkLaGKTckMtykV7VvkkGCnSftsvTpcjeFvwCJ5P0IgzuXJomIxejUPZiyi/jf8J
VfXNjl/+wpUnZXGsuS3Gb/prg5kuLZL+0wNsemBhf4Y0e5VNnOAKmuBFlHdNia2TFPXTsUnDfoUV
O+Z/M/X8qKslGg8Ja59cLDxphMh1ZFLy2OT3Z0JUc5hyD7YKY6Ib2c74Cu+iUnmmErHXmrARO5HG
Dyx1hpdI10elhpu8Nvt2tM41E2n+fJjwFB9MPHoRCsO6UxaMAMmctN63Om616gy/5uBiQIf1EyUU
OcFg1CBS3u0zHrn5k3pjJeZdmeQmKDIFlInGBd0b9Mv8L9WuvTJWI8ddi+A8pbdXwFes3kqY/vL5
E6dXCDEWHnIR8muCDZijMnqajyOCiPPsO+I9fR7oCHiGaYbOGCJAHmF3LhgsDTeUc695b7S3yaCf
dT87Vqw/TKiQe1rTW+W/XiTo5e86QFOAQ3EXfUcdyrruqTkNqdRmkaD/poNNBvKS5JLkFQc7a6AP
XKj/w9SoX5uNR4hrTHEX5zBcDO30QmjHee+autQfGe1Ra79tUZzfidFoCv10UR69MpUzcCsLCQxj
TsbtU1vNesMA6D4gCF5QnfNv0oLWS2vzGGG/EeuelMoewOwsR+thQaswxAfITFkUM938SHcQJyqL
JDyfbJmJZQzm2bV/RMZgpxLkbsGa9XVxtz0MtBj+IKCj+aW1l3DYjwblvKB1aavGDAoFP0w1R6by
9MT4pWABUwBz3fGYJFDEhKu23/k7YXD6JpLdIeZgEaieylV9V1uS4WVO2pSHMe8DtlmXsHDG7S9B
DSJbv2nBGwBw1qQD3zfNJzT3d01GeyTS9usyYA90CQGwsMySvPT53xxXut1tCugfBrTl3ShuB8Om
umODDCdnwvueW6mPqykFnVE0AX0pRfwm1aXzL/kwPennSHNURdsGOw9rX95Gk76ouJQxnqsSmzU0
ozVTdkFmV7n5S6B2C8v5efQMA1p1P3oaxly8J4wCvHOCIGMYpNgwFDJv9O7DE2SAEwo9u0Nt7Z31
Py/MDCQPUcRB5gV7TVYiNUhig4z5xRKsxkRh7sE0gmEKp2QIhOwLOllXo/vCRKioF4qmrT1FsnCT
r2KFRru8znHt2Y5iTY+jWoIOyMOPuBVVnrmQQOwei6EYDqcchn2NKcZBbqV1SMzraX6G9rU3zzNo
zhrNy7xyofw08KXaUthntVyOzHUU17TM6Bv2eyfUXhUTM836/dabJW4kaXh+IOQ1Lq0A7dNIPgn+
D+8For7YiLrCoXuF7+bDE2HGv5OU+tvKBOy4WxyaohAih87OyVvavPsIPEDk1rjvmMcQ8y9MlORp
t7+3t1O0KdE6gbWSrV7IB+co7OwisfDcxcoMBQzSzinqYtgGjg3VEcbOKGJdAg3wTXRjD9A4VdLC
Gba6+h/4IDCjW0nFSxKi6icZQ5AF1xY0QwQvuGLp/H9MvT1tyMVCFx5cGDG7SNjZFft5EdY9hKVJ
AjKrf7nWnxKu6fx2NSUoaVZ3kkxLl/qLYV47T3AhWW1Pa/hJX22b4rD11vhuRPysuOzVSKBBFQKt
AahBi6q3vWgaPH6W23mOhKQ6W3QuFtRZF5N8n51sjvTuIlp1lgKE5fe4ijrmoI+BeWKw+lWeRlap
Lvhd+SMu9Cv3T6TbWOyDtxQwIln//HSKPCecT0u8uXrG9sKVBdb/Q1TQ8k6c5Dx/1PFUB3vmFbIx
BUjwUW85TMVbRHvu4IjXKKlL/AYSFf3ouA1sAGpwJDRDABgsUQiND0Lr7iu1GimvA+L7M2AZBAxw
2MTacWJbYnTdEm7y4TNdXOAkIkNpp5g35VZsdBocOJCJo6t6TvtUGN0vTXBNMeHaOcqc3Q8GwcAy
GIix9wWB4I7/gCl6TjXsL0DGbjpQwM3obEnXRHfZxesUvsNNv5SNHjyGPf4o37u535C5SHteVL3F
82wMlfMmcLNXQ7my2UaTa0++smI6jv4mb7CUcRZ+4u5s7wT9GvQHyuiuKRPUE/PJIvJOWlIeFwLQ
D/w1LOO78DRMMQ7ERFWDjWpiBKYzDnBOU8Uqlb+rINEx2ElEWREgkSx0qCR9t0mESLnE0okEpch2
3BJCM27gFA3QGpJZQDi873iZN6zXlZHoFVnnS0s1SvO4sL46OOPAjGqCtssKSHYjb9CEej5ec99x
IRoytZd/6wAOz2RHYBKYbJPAl2LXoBzMeVmPiiyX7JMoZp0r8Y5kRwkFJqVfdtIk2Bvgf9yd5NIM
hPBsnMOpMky6hD5ygy9ajJF/sthYnU/RHRbqsKpRZjLdHvOb1RnsuiG/ps39B6awfvBbd5eWKq7I
2o4bH5a1pm4pjSbcKulwP99blo8mIFqst2TdSwOXHebN6q6TMZl0apODK3yGrWYWu44DUKSGvNAO
Ps0EcqRL/+T16H+T25WEuEWbeQmhrcItQR9XoSkgO+o8JEn4CmWZCqdWrxXs5KI2kwTsuZgpeBFh
y+b7ohfQX3bhjh1Sqon7P4yQrjrC9wmwOkHHwXanbZ8B9JpdI6RV39OZ73w3MVyrfuieiJ6ummUF
9adpLps4FNVQ9tQxWxp1RHo+AfiLh9sM5GmmIsgSILaneNw5ogQvEGpWjtvkcaWGYPBBiCFMxF0h
5RfqAqtrHTwJ51lBZXQTIqJnJOR8/watgYBVmGUYiBXAWorWkF1r7lWmZM5a2GZXlzUoRjerkq57
V+MlERm1zWdHvC/44eTmHLBO1d6+v4J2M93gF7w9WpkowtQE2VLa4P/S1J7bz74uFjAtQwxwMlPv
nm+CEW4XKM7S6J+PHFxCBkzvNTfSmeFPnMKTUa3MUKSV5BroZscps48CuKVj2CIJztRVHXN03OLB
FZ9+DmxbYV5X5dwVNeqOxuZdjy4n2YcqJrLFsccu9Jf1If7q5HBJ4I4nJP6w2wZeFcQ/YDzMBLtn
JtrkJiMZbxlB05Wq17FuQH1IdU8iQ/Hm7ylM05LqTIUFdUy4vCvnjEsglMKqlI2g/p9q73NP/rEY
KB7IahqacYcITLZ90XQcYg7KWquT740wMrh9QBHDB8iz4uv/1+CglQgtIE0e11eGxXbuztr3AopK
rgibigaAN/oh6U9N5S8E3WzuYi3JH+L94rwuI7FliTcpGOTWULsV68/iBjQAosHuTlNhHULv3DGg
GVM4VKlonTiG9xGNZt3pkt3/P54Rvyu/qM3kpTFqDTGTkUOEadd4qh2grGKgz4MqcSUqRfQsiGxi
JIDm7KGMnyljalnbRFXqWenO5cq31w1nZJ69K6ZwxTW3fCS272mqspGEj8wdlOpHMvAd23rTIu0H
1DEubZzyYUG0YXDcCpUCpyXmgLXtxGiLA0nTrIoyZiLcK1g3Ta34LwajRD8kZr0ssQ6UmmyD4Uxf
NQQxy6IKhk/Yz67roZYZQwxJ1OIyxMYfFvrgGlWVYZpA/t8Nu118ThKrVcOPxwJWbPmFD2G7C8Sr
anCQnboCh2XvEpdJeh05JMKYWpg/d2WevOSue1CZQNY8GmTZG2gp0yp/egURtug3cM426CRJiKYN
uK8TiIai61+DeNxO+0qND42FUo5OLc+5K6gU7/3KTJOwWMBmh1O1EgKDrrsdAIs9tXc34RpA1+rJ
rIeK6R6hR0EDRvJScrRDChewYy7dx8UFLDv1WYE63c5jVzU2S4LyYDRfJpWA6/G3z+uhz9jNY+5X
YPp/HPgXFjc/PbiUrHu0V31/qKtfk1m19+5XsMfOHa59XHo+bOwU0877VEjvPkax+NT+BfNXi+M7
GMU8rGyyr+4uRamURBl55MQJDcyaMbjZA64rVwq5PiUFjfSp7PwovItAZXx3OxNKaUgzvEanqmmU
y5rsXWDcOWlLmEr4q1mNcdtb+UJLAsnLXOok5QxRc8LMlHdNDk/6sQVNobb0/QAjXHRQxF8PWCmD
8Adtle6KoHRNV31crbyrmkDK9sMQTb/ZjoCytZTdjBL4xtd4G2sUfsewDyDHIJTkH6bE/+nZns3M
tJhd+OcyPzgAimY5FmJ6UU9jUSvbpG0RxnZ3snPAbhDd3zuuweL+u92AuNgnxxehObTLvUHG/h8j
i2NR29olIHosicTQ4Gtvcl8pQm6jB/kdNuOIFb4uxXFy3hp1dVijJJM/GVTaqCmHOD0fLO2cCzdA
KKIn1v+oue3kDHdxEy6fdJs6P1gFFrIPW2PKhwg3nqDOrLb0Ne8f7LfrGxrfLD2hE23j/SnMmYyf
7RDSbKbSz2hfX/WkoEy7NyaiueOyhnSmNIBz4CtwVkGcsL86WUvx8lbCjl1CkDTY9eGPeP0Vp4MO
BpgzVXXT1IVT8eLtOgZI1Os2NcOIN+CwNAkL7rx2HdLak/IRnRJOcntALplzHiEH0gxcd1Fb7UHC
fYairwgEAywq8bFPDkgNnmBUAYFF6z76ETPviJlUqSmuiqRA8AfQkUs6w0W0HK/W+3vojcdGBiYc
h2T4Kwr7OWPxl47JqlMkUYun/h7TFBO1BGFyqn3Oy+X9HBQhPmCF0IwK5tP+8FJRBEBtpLrJtoQo
qqam1UUtr4Y5fYcuB1xjgF7dBI0IvPEVbcqVwog8e/R/W3mpLRlO5e2sTylT7qttQLR803QAcsWS
G+j/hl10DZJd2usxHerDMVdlvrLOpAoqRg2jNY/xWNPebGhxbktxKnB4wtmHtaFbkm7HCUdcPJuZ
0PaOAM24BW+APSHgA4GMxi63dp7RC3JhaUCLaXrCYqEwW9lDs6ffPX7dOkNS4EbpBHpG/1HF3DAy
nmfrqdxmiYV1K9q76NXIpzy9+5G9XrNbhQoKh2Izo723gkrzjyRnJa9/oB3tgMl9o69P8HVUmYck
7ycupzNYrIvx5AdS9kfnXgcyND9RuMp64MPwLRmfra5Fox6/UQCQADMooHV+p4Dw4V/IPRBvHiZ0
MpRWqnMHMf+roMA18E0z2UIk2CSlMTiVB/vSMYbKaq0r4cNMwrL/8JrTZ6/OSzNeAAlcXOsNSQGa
FNQKavv5/9pL4nRgD6dYERb5pcvOeOoSUwoHmktPs3VJyhQFTSVLsLMpSpzDoqMAx/zX90s9VCcL
sx1Cyy2IJlrI8kcjlFZb43T4Lsp4YvEfLqjKl6onCdgKmnDp/e2UayXcUDKsdal/z46HCqEc0oDM
rZClwqG6Q3k039kLuO0UTWqOST9h/7dJ20ldbzmFMHhnI23BZFzv5i4jE3a02ARVrI31uDu/xM6F
LGdbHHC5XfbEOhqafp1z1x8Wi1aP19Lob4zEHPs8XdaV0m0J+jl4sQv2AyuDZKU/lL/XBtOKxjcw
f8uYAxPZUwfvmwqVfGlNcWDhyE/SUy5sdiyn+gAUnr7ITe7sR+KGYLvzpZvpqJQLKNMfXWY1f/ed
smXh94X6ZcxiBB9i5PmmVWjIQ4Fa/tbOmjfUhpisJDiHCP/bp6V1tRHKqY8ABp6wXRqS3D7xIbwu
qRUbjyUeFu2i8lNCSUAffBU39QoGjbr1MjCu2LbxjqxEi64tBReIOB/EIgvKIiS3hnDpO6JsFBUb
VeyBciKc8JS6U5d6OAVrD2FRZv5iIdH3Pzn5zb1KA+QZo81cv3xLCMfEPcHMZ/XZ7rpsdpN+O73o
3aR/mjs33x/Zt95/TrfmB7biT9QIvG8Hr0pXof1mATEZRdCetDtazyOf1yekuX01OFGeR8g+HgHF
BsZZnU3J8bzORITxZw9JJ+hwFUcmPK+5iF5UFVhMFSpNunSwRTvVvusAnQiSxAEMLk03OhgxjM07
SXRj4bGWhPrCQBu/VbvKFYnLCjlxDTQ07l7zeSDMdeLRUfo1ww9XWLgxzV6lNth/wp8xg4S4N0Cz
L5ZX4hQ/oGG/68L8inB7teVjM7MGNxqoiotd6PI2jeq8OUjju4NM4uchbXsGJm9VWtNX1P7gxjyt
3F5ljG2SYMAYouH9AnudDeJ29PUZfsuRpnYSmP+IkuFjSGVZvp77dK9Jwk20xj6uKwYrcfWccW90
513Id1QcR/Sxja2iPYPmMpJA+1n+jb11HavXZcI2usnUFTrr5zwnZYvkCN4QrugBmQoWFvMON5xj
2qE9XIhF9HX7Z3o0iF3cs2mB0foTSJVh/9RYrLfvVVEFZAgnR7+68jlI5VnnLMe6O7voQbHhvYXk
6ryVkkNLY1SHGo9zoP1uq0WZdimT02UcQuEN3PFgzzprjwzOkD6pNasnb/K8fUhJqC2Lon2hCD7y
GxKsTC1ge4ApTFQdlbVPiqhS1SNXb4MJcytf4s2rJx9VKO1KpSd4Oc5IyM118bOgqPhFX81L2rSc
eS+Hu4POBjj5Eo0POOxhdM/gW+LcjRHd8Oi5arzVb0CCnTEmAGw3F5202uAq5WQiaIk9lH2PHAAJ
PA0yeXa/4iJ3jbPhI4vEfGEwBvlBGfe6GQdaHDkeGPjF/xJQF9WJhZAwyThgNEt9A0M8UPhIk237
ltW+mijXjBvlzHsPeHR00eJR1wpg53ug4lKtCCyXucYTtKfwqEptHgTvjRAgFWgFExZcnC2SC9qz
xZx/gMzgFzVUjgokT2tWIRpKm0vyohkciUFO705dUl/uUWu2j3OksUAmO4UICWQLEjJQZVE+aQjZ
XOEngql/xhczUfcA0/E+xdWctghzoQW9hUNdzAqV6xD49+J8GjXW2xBz+hyf9yVwUwKu2eydWDo6
BEKdlg8ZnNTtamdVELJ4FVJtFRVFdmNmashkccYtuahizEqYQokDyct4pQkixduDsR4b0Oh2dTdC
EPGbc7cjK/nig87yZlTeUlfUq7qpBi3EBgohxFxmVQZbh0EvYUWdAjl2dvmpPGH1rn2uVx+ntURY
MT9IlazPaXimCOnKLZpeYQHKZdH4hTGr1U2WvcXlYOkWAcGvYb8R1aYenLJ5T4m5tjk0rOp8CX1o
vrAbnJbvIAb6C9ozH3MVBId3j05SdwWGSQSQE0OcQAj8MYDgbVSNTPzwYgWdx33wT3aWJR0ra2Hp
0O1c2PmG7TP+QK7Fds6HfnC4jIier1yAxwm28iSs2A9jZdmH0gFRaKR5fJSC/cHlgKfojm0gmL76
2A4BrY6UNk3T4r3NQLIhrVRhwjA8chj4xqZHA8IkBKdo6lfXGpsE7okyf2JMZOh0UbIm249RHBDH
QfmKBmq+ty+/E5+UxIKSQWS7L4yQiQaNcoZAtYSU3Zq5ZHjxjYZJd8Gs99Bv2zyu9ZE1T/4zkBiQ
BB5KFiCXz7gdwr4jxq2ksC0J20yAoXrmrFsNtF4UQhZx44QTlhka9XMZAxGEkRvC7ZY40G21ijXG
MND6rr2espmnl4sfmk3zBICde5u4d/eOnDnmZ2sQ35KisZGkv5qiTX9bR71WNqfJBiTroNuKgsDP
eTBaoSKCemaYFZ3fNchypLH2wBxMEmyIUMseDjl1EgScjL4pLHisQfr/e1H3jhv9UodLVbDQ0oq2
o924yTLzs/Wf3QvlqvM+giMQ3vbqtW92rGr4tbGzHHcSFmZ9p+u+9Vb8PVk1tWcqac3yP7rG9vEd
dQlIdSzkW0eEBYy+ap2PW6DGPrVTedx/nYYA+05euLSIkycZS7ZZ8Qh292c7i6XX1vE8iJDHpwdM
U+Pt7ITY86JOdRsLcT8xVCrffx0wGFuyXNb4i5ltFXcUvAgGd0/w3sigE4wVFuSXnBbL9/v4bbO6
2ze0P1MB9VhnCXRCUYcBb3Vw2N1rkjQfCWoXl/cyCJU+i5LVqK/A4Ugi8uj4+7R25WwVVvFYuTjl
h+HQKfptJ+7EXeiva5Wdkes2IQaIVE19TKUb0XOwwjE+zrVAZ6x+9jzQqM3aU45Qz0wQxDuePN6R
B0ce4xh5mYG1a3fPalSTJ4VuWnNY6XHD3JZGSYOSMbjQkY5GO+vNEZQoKqNIyQaqIz+O+BEslJqm
G5ykt3gGZSdrePLgVPmWCDcyi7fGwJHQ9UJqHbIp1pYSfOfO+6/cYyuRLQ+LJeluNXGHBUV1/QdF
jsT23QSrLk1xw7c1dJVlrudppGMKh3c/NwuUyHZgys+V9c+FaHMaPT+P1MBED1XAxKDg5INuwKU/
+/IsWU8X5oUcMaAeT7SAor/nSqhhB+jIPK22cay5DV9YgZioAGDTSUGOl35r9JPgN8+jTiW8ySlj
EU+DAslavBkL45KzLxKvqUlSwXqcdYUAvIeNu0Rsn7CxdVKfpXEcpviV8nzcq3SFWaY6NEeS04ID
G85ikIakhTPKS+aHq+o2MJBY787KbMSZg7E8ZVaSP4nbKol0q7xPBVxGSesfLF3g9kYF74lBvFPH
PmjuEz5hL12yLTYrFGRvlc8DdiLORpgCmHayaVXNa3qnDIpjXYH6ZkVsWstDmHkZ2ZTEwIMFpH3D
k85HhT2OhTuwK2JYmlDBHVvwQBOsHUvMmhBvOGkX2qT0QE/+hu10eco77imVTXDBTgOMA9cGMsnq
Ts11cJ5ZX44akxAQ3wc+ZykyzFAdf1BZ9NSVkKXRNLJsDO62XxhtrdVU/XTQIfFx11v99/M/bZlq
VSniQwnefgCuRPKWg+/BDOuMhSEA5WIWKy73ZU1xucFTCW/UBj3KBshIVz1xW4PMhPRAUFV5h58L
C4zgCM6EzhFuM4ozzaO/SSwqirNljXsurZMML/YupTQJmnhiyJcQXAsgNMCJuYqZtKwRYHmIW8wU
7OXd1Z0pPiNjwuM0cxSuDudz8BNhEhlcF06rQpDCFB7zdGK3QCcWy1EW2pSHMdZ4IfFjgHKaIze/
KaQli2JPacQH1AQ3zzEZITvaY+plcCUOp/JthyQxLzHR808fEXG7PnxJHaYpAmcJch2kk1S1Rqhb
p6We+XhQ03ooIECvcniZy8s3FeQEunoOL/H9VZLJfp9vWA4d3hpEA2GSmzeeSNih7XLTXPSlq2tg
63D0yjLPIAqzNaQ1+Ibbj8o5d2WMaFJjqzpAknFGHdPiCO0tMY50McsE/uU3JpFnzMfgrC4ypznC
e+pO5aKRWWRZOEMEtyF/Re45u0mBpQs/0U7V2Oy1T7HkrhFXJSDH1XumBlOwpMiu1Svw41+PgasD
Rsr+7RNo5jXi177vf672Qqk3anNBjJEPYhjqXch7M9+AKGtd/+y8fZLsAXDXdjOE2Fm1tDmyKe7N
Rqu0nA+IaK7KHXXrB/BrOwKx8tBgDFhLAd8j+4UlhrFwu/nK78vDLy0+mdxUEyGweURGvDbPqffe
1P0S1MaVCO0vr1tiipNTfhRmucrXMepph0E4S0XVWuqvLkmlwrjOQwC2FR0BWX4tyBN6ZiMQBmI4
kFSbYadQKqZ5Q6itTujQgMXHjxJVV8Ln43aDnEa/aN5VmoHZINYuTKvNpq2Yng6xYqn2W5E5Mthv
1RcJ9kWU9jEpRkBx/ZYxSFR/2x4iYucPVSVW+U1hFNfn6LwVqnIc4OXsR44Vn3vptA3Cpc3vZB7h
EcuO9I6gZSyw8398/IaAuL9h3lUeCN+GQpb9YLNjZ7WHH/6Oy79LXrxqd7TDw2xx/lDSIJ85pQis
nrET/znGEG8tYqEMAiZm99V0aJpot1qcTGSCqvuDJ2vcfMjBbcWtPx2X03zLKYrhc55HiqVr9XoY
n2SF6E9W1CwoSIYAVVewCekfMLF10eP7Ul0Sprnr/+1a6vOFcl+Y/OevTyvzn926FmOqdTm4eI6n
sjTpGxaLeij2cVB/Ewk2a40KzL7XVLKZPtv9U4Nk90/WEUlilLsOkq9rb/0beZyb8ckmEBWohLc9
pIt6/uujoIA4qICxIq3GoSy6OEA+DTT3iB2lH5HtymU3N22zoAMKUGwfCCqWQQHX3+kzQiwvts74
3hWVppsrFwHZp/OVr4YKgdwaI9bjcDGq0cicuxhbSugUaE5KGtqIgoPuaDCmWmjgl0DjCKHvA2Ng
gPD9Gvkq/U/f+WLr1hETmNnO7SDcYdHj7XvdbWQBXeEBHj1YlM3ImIL+U5i1pYubLaoQnjY0JLnh
kxhF1jrSsWOCHQtKRCOXpOChodT/UBZ5dmjoEegcF1HKZPR1D7jfpVQJmw3cjdYh0sV5AoHs83Jy
xkFd4AhWtH2+C7R9np8nBnhpyyuclC9/e2lIfa3iwChII34nYOvB9Tz4trUH5GIJaQkMAglOAQ8V
FzdBMnJfkZDJhI+VYQMRRRtHizxGo+EBo+yeRbrK4FIISgySy/AiNw3vQ1LZrtBFEjD5+rDRC4Sv
7BqkAvg+dRxNjbYd0XlCyC/x5tpMXPV/kSyWbYO2VT9s8NaQytF0Az/0Z6whAi+qxyhgrT5KpF+H
R1xtkyctiX8qdBUmDVJr5+UbY/Nqb/NqLh1aXk3GLGzO7R57+SRjHx+FcH7/CYldwE646kdk/0bN
kCiL1wrL41FSY0UOLUg/W50k++tgSH59yIaeFsCw4kPDeqhd5NOJxLJ5Q9LCuh3hpNVJ+SdhS/+7
owYqIHQIpJ2IfsmQkROQCyLV7l+y9dk8S6yfvDHLGguTpjdxOdFl3HG5YeoMuGnqTJE0yMjtLgYO
MtIBj3WonYuOJxMsu9tOL4WLb1rAD0QBrSfmgBsaQHA1POgYeuUbU5qTIlMXrPDTxLskT12r5Z/y
aJhGOVEpME2g6GuXhQSRNfQldM5cYB0n8HHagpTwW1/MkBuVdFgR6/pMeyPgwCt29AXK6NBQhErs
+Rj8Ix25gBA3e0qJyU8KilXKcXJqaeQ3q3vTieGRN4JtJ07T8/EH84jo/XU7O3NjG1DJLgEemhqT
3VMBg598/Jys1DPEYJF+MFhY0bDUjMa/qCwtFhF7c9+Y5IP5Zqa3hJuG4ww0Lk/0w+5iFkHZLf21
awP34jBl4jUt+KwwWMe5OpTZJ6vrI7/ohAoT2oUO2/Mj3yKYSZuEH+UHrYBZzIAPsTad/CLZI+Lv
8uu9FyJoq0Wb54CWSYxY7W9oxiHY2X+rd7D90MIMBzbvf+9mQb6eDfd2MANjucv0/cqY9W1DJZ1u
/QJj7xC6PWdxGFdH5qx4SCR7BrQ83caRez+1kkw4fysayxZgLf5q0xuzjHxGO1WUw0mxYQcLdP+1
nZVFiNFDvxDfIKU7xTuSLEx7j3QfGiiIbvkNV7kpKYiXSgByB1UstLoothsKREg6twcYNC4vQVtd
h3WlecjHBrZonc/0a/cNG8ypYGbY7dMCRgv3MoRKkMteAkUNoDVpkLX1SgH4ZqTnJxXbroR4gkGw
8d7xBVSkWFFx4vSNXYZa0jqHT0kSlNHA8fSiqmQHIwhek10Ro8MRJBm6j23MZ02EUTjXz4IPuLp8
mWqAVSG3OvI+Tc48TnNKy1yhDkrJarC9OqbnGnGLYhMNBu3zyMq8/zTrRXLq+fVt46NcU8+dnhmm
HhyB8zfAXqKOAB+nBUt3XNT/dnrEHT6Yv20sXz307UknsYEWSQ3x7+1QMQtmd9+srPjdz+ZBwE7A
9KDyl1HEDdZQ/WeYXHf89oJtbvgoZT8IsVuA7JOYDbDBsi7yqI6YRfQoBS6ToOvzPyKk0VbtKDQQ
ypBaTfHeGHiyqT7XLabTgsh3XKdpxwBFDgiivl1jjUO7jp3GV652KVy3Aqld/xMTZXdmj8clfttz
wnQpbOtvfj73vgZxkApcb/oYj9uFYmFZkeZ/wen2D5VhzkAASlFfx4r8PddZbBILZCYN6zTWGnFl
hzx5AZfKAn9TuGKIVF7e0slZjJIeNeYhIW7O/FKIFCkmkzEJPqohpb09ivnCCh9bUFgL5O2w0Jb7
UU5F/LzFfNpvSItOwYFqjcAnlvQ3F7FRZyiuuTMvQmMOWRfeNetMWJ/GDT/EzVilj9HsVLvxaW+H
v284jro444UYD3af9llBA0QzBPU1NJQNceh7iI23+mhmAaBAXqj6gH26yrDGrWYLeAj0LVXJFyPM
gMnHAuqqMMgyDw9lM/knUMV/4bBwpu10eY41sSsqrzv61edvvPxthfEJnQ05uJn15uZUvUNmAIat
mI5jVG2Q89qiiHJrUuSnyu+tmgNGIzKfh4hreT7tb+TU+jiEQPDmOqb3+LnkkV6Q1OTfHfZ/a00c
fgjqS2PO/nrPWHEINAY8C4WK/tivf2gDX5V+5CioKrMqZFC5bukkFCmYCIPRSTa0GjW1ffeoofP+
kY6pRIRLFjYprvOFw6ooA/gRXTCE+fRySevW8/w0ukNFXfXdnZpanD2LqfYisXTDactXM/rUL2Q0
/ZToL/PeK0o6IbbER4VM0PDrIIVQeW3pwsT0oksfUMdXAAZEVoxnbrQ87XwGH4+ZLc6LWST3bhbr
pjRfb48EuYUci4SRddjUJxzLp2Lt2iDEGzUGoKAlSlpC1Ws+r1uQJHdY6UA524WQjD4ppcNDawvk
yclK5LqfnfoStkB5Q9xFbNyXE04dLUKF6RRhAtKQtdW/i7Dk+g8+7NEJEvtixWeWiA6hrGYWJuzi
d87dAFbJe3BHAbhb44+ysI5VOQWmI+kVdNiB/bpuXu38ruQ5uG+QBJ4FAvir1A23MaaQ8O2Vc+to
eCXF2jtD1N7hTjZzyK3N4IBgDfN4dFKBQA+L83xKta18Mi0hDbgHYDAC6eXTr7XHmvWvENgCft08
w46MfEejnxPidblOimCvn15ttvsxLINJshz4UGxocTksYjKz5TpzeLia3oLeGWXjJ+nUEG/0SXH2
89EQGe1NLmZ7HcKunA61MdLFgJe6py40SBI2sKOoRd6vJvaaCPjGy+dtTlMf4Zql0tTgxeenu7pX
0YcgxXCX1vC2hgOtFpdX4t5tVCF3yB16kFLSaYVWGNk1zLdqkOMJNaV/DuuCdHJxrPzuySPDl0/0
u+OY32M4qIitN7k27uMLBSbUCz9Anc4CMj/PoxjZJ3RbBCnViIozFw7aNAOQUBMZfUVSEFrU+0gr
kWolpE1eC/VP0BG/GbHe1+DkNlWa1AMgNSTXYunEnY+OEGPJtxOIAXzpOY4YiNpEq1DkYIgaA3Hv
4ehu+GuPmUnJ2xXvibBy1HvfviEov3mHuCdixj2I02RJ/qOiDC9Ju63DlmSuZ73T41Zf2ujdHkD5
C+xuRHbrB4t7hXkMLjg81UhY88ri4GLjpfSthVJSH3lUWj0xHpPBQ0noZ1C9SD1/Kk7cf5Bhidcn
615kU0HsfIwBtMg7JJg6fhChDWYVUwBAvW+zS9w4dQf4/vH36bx72vWR8arCu9iGlgU9VeYwc9+a
1M6nn3EAbUeDjQlLLt4EPEib1LNqbfzh/mjPb4LCF10XpKoyZ9mMCaNh0vI2ld+HsfA3oaZKJ9ep
gI2lRfvYB8275RwQoHTzJEOIpaTIryuVuhZ2ygDdvTdYWHn7vc49gEzSsVmoHxnlQZ0MhG+ecEQ/
VW9dJuKehv1YfwwUzJOhR9kQT9/k7WATvTX0ff3QaIHxPmm1CRpMo58FfM1nAh1R7NRXgGJzbdIV
7z213WKgyNuVmlykMJhIsxhmvqFQt9ID2qoBlX7HTwT1Jxcp9LEGJMRne22P1CIoD4pncqYXBiMp
rKn25pYybY12FAwMKFdFwc5m/7Huss7cp+vyxRikl99mk7ZhuI0UowSNZNjd2gznLa7i9v8hmKPb
QmT5vUz2s/E2eT7eY1ndlcmnztbUgs6TlyRaLpjnURNLH6UYsN8wx3/HgzyAAQJNA4wqsnxxiHaU
xBaEJ0VZ+ioWJ/WLThjo6RImAy8LP6f8kpxqEMlbsqWySx8y9pcgzBrIDrwKkUkeyDZUr5NSToW+
s4yjZ71qCSbHhfy1VhLxaFRi+Dh4TwWe3PD4uR1bU7jBABgqTax91hSHUxg/g5f2dd9uSj8LizNz
d85ytDiJPD0RcIOmrY4l+LQ1fj/zVUaEbdT9pb+Des85KGhd5m9I26Eu9pkXiYdU7K8RqJwRlf/7
ROunoAOun7sFeEoSohDGoD3E/2lrX+Jl5dRncpZ2RetIabaonJlu017MT0Nx71XgfGdLbM6vjSQ5
Y7QD+HG9O9oV96D3e0HI1fGDAy/lMoT9uwa6LLOOrVVvdDHxmm1+rDsJEorzj9TN8NPIqVZoHPpK
OI/VI5ivINkYMfcIq0yGIzEhPZpWBWHxbI4Gc6DVfg5cPlHwKMt/OenGkKyKRvAykzxY+q7ggPy1
10dHFbc/ZrlrBMqXqj8i+d/1rWfzWxl8m/06H5/nqqYFaCpObrW4GTxTIcVrLoDazzYKr7O0JSEl
edSe0x6rdFsw1Vdqh5Qs6UQ5v7oK0zUFdzn7RMtcCC3H+knUZpaqN8LOmIf8JWjRCu1aA20vJtBA
Xk42z1qp43eZgvprbr3X+6bNHbhWjma18DGrstSloi4ZfWy/0H41FP2C/sSWRg8EjN/DKF8oLUb8
aVUzaM09ruhUyi0dD4V8rXqFJMvIBVbvVcIh7QhYpZETyzBBC2pcQzOnAlxpjhDw/rpjZ225fZD/
L5ii7dzk+x24KC62QWih+Iapvms4OEvJYbUM+fNnk+6US/g/so9HK7BC8+2cCvzdctumlapx2b5F
O6ixD7j++44rtumiy5IcTTJDSi+B4fHJ/Hxodwnzjjq54djT1FHkvXGzzXmSIH8LLRN3dXYP1SfY
dk23REs1aTER6I4v6iljOk2wUBpOeWqu/TJOQAxjLbFLwyjBet5AxqGTLuPTEqJ0gdRyVFr1dDpM
a+dFl2Ik/iq4LjEWupmZA5wlQpzQEeqZKCWdUAqRnwhInxZkJW8toCIXHyut6qsNZqx0hkb5KlTa
B7cyOgfFXrthhOrGm5tmg14iVadBDG4uhBcnqiETRfx42RXWVEY1QoVFg2ndsAX2HYEG3oS5vjDh
ogiR/+oW2YpOdMd+CAR/ZnH8nGqWEHHzdL2WpAJ/TPZhQgSvQpIJVmpVZGKWop4ScHVvDbVYMvVT
9vzIH2+rqQkWW1B3lU5lu7V7loJXfYKTpjJtjc3b34wApqPQKVeSHim3kC4A9D9i3Kd8wlaCELA4
mrCo8nptVEVKFkV1CJK5CbOsukE5jHfhIRn6wsusIvZik2n7FlU1nGmLR/l3+1mTznlerrccyF7L
k+lbKJDUBViN72W2BqkiqNhQNxQEENhnZ/JR7GKs66ahDcjsWE69hZAsq+tClIcCOwlpohsPk3Wg
tjr6CqgBWLlEdzN/qv8cQidRQcULJaXQ55f1r6JH2rMG124YTZvnASyMPWYwFs05n3j/EpZpU7Uo
cFJEeVVX4K91cDJlkz70OYJFB3aHDOHK/7LK3+4iAmkvulfAuTtxymSTAv94DsOsa4YoDVMyURyU
aY7wWrPgN++7DO/XAzuZkSW1hteQAb/1LJPxnagAmEOvhFGSIPuOshHJBiqOTJcCnt2JKtwifLNu
q8BGy4n4jMRJ1txF9s3q2vTPB3nUWdG+JMBYXKnqI53wVgejh7szl/9wHtdtgeqvQRnteYAk/6Fg
zXZFvQmRmzePWuRTLwnkrjf+p/xOqKK5Ws5wIRiCCXZaZXg7WKHiW/6Eg/Zt/hPV/3n9ZbTmgx59
gF95IcAKNiPsTmqfPZhyBgs4sm/x6hP87way5x9CnuHUbBMPe2SR2xrfxxqkoxZ3O+PlLyiq9H+i
P7I1r+VM5X0bJBi+yiekP3PUK6yM+PMuYeO3zLMHvPkKj10GThFpvzdf40wPsLEAB6MePlUejQKv
gkkqpWCDJGggV9UZtSFLIdvecDCJH7UqjC01pzM1Z7ppWxr2kx65brTfAK01988bN2a4a4BWs8Qy
+Ht8QaqZaUwGP7t5QVg26MN6bQBUxTVPhpjs+Iuznay94SAzuZbcjVq1tVHJISfO0qwu2jxe9kzD
9uTgW2TdG7c6Hvg2KgI6CsWyrYGSut80ayUG6aV7g6WB/ZI8SGhQmTAC+ZIBSGjEThlRm/u1sD+m
Rh92WEAX9Nf8DnfD60mcqxwPXgw1yFMWyIq4bqFcc9NuyaeCo9aJhSZDOtNfQYRdxXQ81lxa8O7c
ktIauWKTexTaLZYLm5oivwmCySpXI5V6zPeCa/0jlmwVwRzBaJYrV+mM6t3rJrEn+iXCkCsKYa6Z
PiB7vZmGGoELlpp9W9MPRR8Yaak+XnCPNRqoxTFVhcX+8olqECVhW+23XlpfEdIyAQdEjsNV6zo/
eg03FzlV4sJ9VyyEum6OIv5IBG+47iL+K/X3onWWpJKYQtjNEr/dplifzZvnYB7kxfU3KQzkKiuu
4pXn8ZncYWnekoNc4p+MHr29vVptCAKQSk0IhRhTlZrYX3is9GiIgIv3inFnCxDIvWc8ixa6rtFV
zMnMoICOiR4QiTYxDP0k2PTMfI+lwwrhelZnqMClexyfXThdrHaGw/+DH+UOB21//2DvPHe+LO3T
rTHpwGdfFWPbywIx35fjxOk/SruQQMEDPNbRVMc3v6QVdzwxxc5c5BfYxPc0cVR/gTvXLV5AR25D
Q072Pbg9O59SYMyJUDoNAnxLlvIe9+kmNkRKjZCF+ydGBeNbxf5G9GQgMZwXbJ4aGpe6F/1SLtqX
H7Vz6y0JoFgDIF4KShzMOpMBDGlfmDUHYEtgERyp24mbxNqQDBI4EglCvc97UCezyxpepyUme6tX
h+Bb2f1L+xXAFjO8/yay8LI0fFsIJFW2dcJ289q/kEh0JKCpwdBBZFDFoL39FDX5yjQ3cYsPF7Ts
37mPDEHcJe3ZC2Y1dCfaLJ3yWUmLz61FrxMqdzEn5xCvcNK29HMCly61TcjK/5u7yUGsKEUYaS0a
rLe+FT358bxySIvG7MS6FdUdV0rfHyaZ7OWTLGzKlMnLBe15iJzqStd9eAKKWk33TatoD/CVpDWV
uLCNofbwO7+0zqfJT4ckm/4SQ8OCJ5puyfYCcjOXiXHR2uN5Yg/26UMZ6S6eeKLlhsl8h3kKYHXf
qhu5gaJrIIXtSuJ8g6lM/gggqlSZDHUhQPBgFc7VElFsYjEadORkGmTFhgnPjCXOJaRN74bH7/pE
csJbJQ4FmwO5vtBzB48wpeNlH8jSrv/F8EGQaa01DGmUBqgkc55x1z1QtsieqT+Q7bBmyn6fxwWW
WP8Bl1fCN+hAblx8tKdzEZItR3VLrLnY7YHTuZsUBMIPGxrSFR4vtsIZT4BEjy46FZ1V6U2YIAAb
SfSayT/rB2cHn5p1p/wc4Y+Vshy0c75PofBGbkGMFXC77TLebXTYZtCvjtz2GJAiXja9khnnsWHr
HSw8Ql9KxyPCdLr+759ZZsHmphDgKHEf9ZDW5AJf00kddD7iDaS2GTVKuvHN2wgZhvLpMl/s34Wk
4wXWNzB7AXalkKO0x1rQxdq4/5ISb+TjMbNzdMXDP+t5qnbQYjKkvdU/Ss234eAWubwYVHYbSfLg
N2aHqL3g3aAc2TAFd80KwhpsiBWeZ3a6XcdM0ae3UxIkUacBzAoeiIl8zNUccWvOG3jpXCQ75e8O
ViEcQuMDloQZsJAK3cZ9A8Q1fdu+B+jqNoDDyvzQBTMshsfqIurrhm7H0IJr0taITyjr1jNqXxib
ff7Q8gzOAWrWdjtJNt3gepx661lEa163MQE4gaXFriffURncER8B7YAju0E2mauE+zmauxGlbbV6
xDEj8B1qJHfS4Cy87PtrRF7mmN42anlFcJpX5j/9QgrfxWP5AXZEgqAXx80Nb3duyvJMgwT6ZAtB
rG1oHbtimFZsL5UGHDzExhkT82y+X1PO13YyCUVKiXZP/sXDfpZEA9EdYlg/kgmcwdlAkcHXw08C
ce1kFKL8HfQY/Rl88XNYtkpe9Pw0s9p6Xh/F34Vpl7mJJe8408KuogWrFbu6XtV7KnTw+zBGad07
fkcQjpbLChunhEjc1+LxYJ0Bao9ksEouftzsD7wo2qE0Xlj2/VdHEhvSN7qMYWAbeDW8cpvhSmxH
wdK0KEzDLxdBfnYbmwYJZJYiHYuhljyuNQOOszcBz9J0hzKQHX27D+NyezmiLH2SQD2rQpa2SkMt
txyqIbtDuLfzkL7/MIfrWse4zd4wFXI6ZUmywHgSdyuZ6kq83CxlA7D3ZBE4UFtnyHmf/ewIo4uC
HI/ylJfV6pXIYKfKUOpthfl5005XJOwSXt1BvQvn9C7q5276O4ezuAEVA2L19eBLtxdqJ4lwhtS6
czy5yTt+mLkECfHCh7UmLEynQUFxkVGt1k5Ss+bEGyDCfxHePnsJSu66DRuKjVKocDhxAUNl3dl1
9hg3uh2+BONshj31y9MXgMWKZXrDyrUQqS+MB/aUzDzt05z1apWz5YifvuZRei4BBStSM/4Qvfzw
c5ejRcOjqRmNA2qY85oFOoROHwTg49pThWlmnuNBxNoRMPuH8A5h+6dYoupZwuAvBwaW3KlT2SVG
fqUVMvyEndymdDDnSOhdCxfY0I0on5YuABJIf/9OBhgDhtLiqk2nKPglXxLaqWonlQCF/t8o3q2J
BlWg8a0IMp59WopzAd0CenSxWFqXZqhLUbmCg9eSbSsL3KKbcQm+AXBDI70XaX0ElUIUep0dFCr3
xY+McnfNsZYM/SHnxhTs+7fPcc6MlOcw0w7CbxzyU8ijFwyacn7vAYIXmITWTfiK0xEkU4cTC8OE
vem1j3+c/LJE95YjW8ogvQqf6ySotEH8Op1dc22+VzGGvYglEWH253x37CQXREi9/SkXE47dF8pY
MZYXKAvEMwSGbQmMLu2dq5kc61xzNQNs4i6ok7gBAcyhVNSCG7KFZQHw6k9vaKo1NchSLQHdTlOI
Z95E7QACasuxT4CVxJC7jitgR8q7vGRiCo7HlUp5d0widEDiwQApW8epCjTv7U7plUeCkV+8KK67
71126sf7rLFwQm+ezIvaH4/aZXkN1qyKC2VFs0nqER1n5NQ8sn2wTkPItcSigyDAh8N71oDWHs8K
nO7Hn9jmvZX5Mgbz+G3VRvwj9zMD6YE6Oi+wNDMuDQyYtnFE1gWQkbAq7lXOzr5JTVuv2aI5SIni
9Ua28tCEnhXC+XYyxHFeYxtY5M0PCu7G5rZWYJejTXMoBbvXMcfN1FVjbavi4pORSCYQwd7j0NdU
d6TVKsnqGJzMqssxiDCpWcECHTVvA6J+B2e1l+O0DOXj3IZ3KLhRQ/XendfNUHX1rsTiEI7W37FA
BoCQYrITcPzK3TIPdnBCJj6J1Tg3HUFDIBWsAn4AkPy9u6QRodYFk2bT4PS5Jt5fXoq2PT7ZfXLV
lrA/ocSZY96t6K5x6CTyAWtIJ43I/se5l50H6vdnTPzSOP5H7spZnMcGfB0RI96f8z69IEmMZy0r
6OGD8a1Xy3TOVPfZTKGrRbcfaq2FP8QECL1zyXf/1E0amU7QXaKoFlGf6xDo1tEnE0rDrfC0n8SJ
8Qq8kn4gqTlImJnGVNqcPkFIo/+RSuny45E2klmPFOYA8B5biRm+lIbSc+FRmkJGBG3cc1yNSD34
MpdQHEIS0CBPBgSoyP8yqPoOSJFQ/s8smkNg3ExzaUGMoRCah398MC/Pg7EiwXGRlCwUroQEoo4U
J7/8cYd/zQZ6qiEWyFlqRcVThA/gk+GA62aPzTy4+b2Dg0eLWdgsWRyuuc7ArhlUsUVDMIf8Js00
A975aP7C/dWcwiWCIJAoNHsFVrZB8ECKNg57sCYhV0HMTsMZ+BtDdPBwF6n23qvJo2t9ZN3DHmsQ
UCRQbMOYNt0UWZZ41eJuHSEZniJu1N3wJIOkmoQL0keDsg8Yby4N+ZFiSawZQijhRRISjf/BFbPU
xiZABKcgihAZ5lCnpqzbcZev2aOdS6nMfTL4imA7+/uBy3Ovs/eBwisuODB2P0VGriNO/3M9vMHi
++ZKet3H5AJ6auP7k7sPThqS3Jprek5qhsU+RhMkvXHjKWCgbNV9TU2IsYe56WfGeUi+k/ZpIaCp
WYEGX7l2ov4W6Lt+W26TRhj9IeyCN/f6ydad0mRCIivwnf2afn2EzDurDcMHqsNFmSQYrC8vaL5T
31EJ5ojwTdoHL8lbCLbI+Naa17LxgXbGK5lT/NA15Cper9ZaBwbCZqBZdWGh+Ht7ZtsQH2ue/in3
RUn7b02YjrNF1SU25pNpij7KlCnjPZqjfL6ZmIdaltj4X5rFVEOKf9RuKLEc+NHtIm9mdxg+Tecb
ispkPqqqLQ30djIWjpVgy31eTpt8m5ElnEF5kB0LMgScwl1tCEvnpJSeK3dk9mvmuhG8VXZ/y5gc
0uTe2iYNkKmw3kCYnZVTb6xtiBaWdccuvNtHoH4T1Fcr8ZD+1YDDf83RWHF+pGt0xjWo2LVl10Cm
PXK1hWtLZcVFPQrT4VKImyiJDQbnDUD+zk25zPingLRncpz/S+j9P2TP5zgCiLsGsu0XFOQl98zV
XEoPm88y6LMWSFI4Q0X90M/27led2ERs/KgPcckdv1bn0B8yZZiAIWS7wb+J08SIAs+AaFE1z270
SP5lSr0lr0u1CbLECv3mvI1oJcRKeB6nebC1uKpncxW8qIF0ufxzaWOTd3SuykeFbZG9eT+Rtnob
ILVfXlOhqV9a8gng/mujElVZukgoONFsiMilvf1YqpWpEH20w/PHdVA6GviPXXkYSvozJQmALxzh
hUyL84Gmxc1H6LxqFteAhBhVSQ8bloYTinwp1V7RCjPHF7DWhN8O6Yaw2cWNvKJ3Xy9CZkdKtGyn
I2J3WUiIHVi09rCAIlOs6TYAMK482mFWWZP3In/M3kOJQC63XbaAdXFXdZDmrkmX74M+5+ZHf8bY
I4hv4IZvjhAjsNsF/FqdFlTOmloTJ5DeKH1ju8T6hq5hKT2KOAoej/hF+ZFWNmaFsK9Z7XmBOs0x
j8NAo7cj9REHbk17BnfVR+aPpiP0w8OvcakLfJ0jlSKfgPXNPFRb/IArMLXBM+0SV2ha5wtGL1wf
c5tsfd2WgGc20Jl3TKJYTqavrSYVKWKJ3uurvuJ/vgahT37vx2OqIitWWJfTlGFIDwXJhK8/y3eF
Z6o+i9+4ubTLC4ddp6R1diYpNcXU8+R1e31WaWW2DEast1CWA1fgq2dZOK0tqEbcO/qoTVgXr5Vv
68yCpxXZx4HyGkX2D51HE9kx+KrJW47iB14icHWq/iVjX9bi/QfE+r2eQQbHn+svVb+TNBRXZ4i5
MSaJRF+PopKcc0MGYZiFN8KTl9fb0HZw6HhkqDt5iGCD4qxtv19csl0s0Omjjkn1SSxRokDj9B2O
6+QtXlHOlU77wyh6F6yL5loRdLJgAZFCB841WWDPITMKGtWqQATaQ91XuHYwYDoFUDN91E520zxy
hJYcDXE0tac03Y89rDP1Q+lmdSuyjIqomSUlwdM0ZlvLGYL7nXFQ0ZcTnVA4z9/qClMJ91jaKl1L
hDRzyfDikQelxdO/TFI6mReeFlJZ2K3/aA3NgzK7SQMGkXK19AHuCXK3cLSSrKTTH9EyfeNGCnpJ
OXsQFMJiqhTM3KbFDnwtd0h2zxizAq/F5Vhj8n9aNCYMsuBb4/vDvcfzmuWaTCzUSKlUnQk5Z3vp
Ee4WBRoMY41mWb+9qcmD07D7myFT1oKTjEFsORpYLUmC9z+UiAlEqKW8CMjVPAADdiz2v4mlHPWw
cmY6Z9ZkyRurm7NJtbax8im+6MLbOsputcra6IAmhAsGyk13SQ73H3UMek17IEFmdB6PPUW6ev5M
oLVPlICNRPOkhSZNjCIOhc9kbeqKr+GXauBctwF3wurprS1+NME+pkThuKeaxXyUgCoU+V9yDbnS
uQoK24XUxfbx7xRDUMk+R6GdlLPMzscw7vc2CkST9/HwxoiDgdUhl/KX4+M5sWZCWLt4h4m3qBKK
AAR973xYTzjhYhxwStxJr5Q9UMEmBmf97R9Izi3FRzpHUVrYoacHB2LxK0rzNRMmkIWXhrfK+d0Y
10qVU/eysUZv6/KjrSl84OmtUNNe6zlzt1tjgKPvlbqswp0v/JoOgkQJtJQKBlAhpCToUybaVKst
CaoPg2gyCPvh2yvFI2xdriZDPD6ShI3YerOo2ILTL7MW3VArG1geg5UKLapQZMJLEszwwaoSvjz+
o9mHAZjhgxg5u7MW4U1HErKM3vGSMFm/Ud5+cCba0uBiORnJ/0iDAbr2IENBKvjAUumgJyaU8C71
bOUWqIIizbB2qPfL6YPJ4+dGhiQdMbAWxqfMs3Tv8/ovB5H7nGEOIFzkcG3GHko0ZnS8o4+Ll3XN
sceSjmxzOwjzfDRAQqVvbsMF5Wn46bYasaVUC3xRNaf8O7YJJMtMcBauHvUQwdHcntv+DYB03Xkv
TheuLJBLU03qlvAPC/7QDIq5KyexnjUWPhSp8kqaUS5T0aDQPzzQRwKGEIbsWbu8mcCK41XZzmKV
Q0R9AeL/39/sHYBcwu78GweGiYUDCnyx82Ry7qehTYliTg4W6Sh/R0coG9MN76GGSCEVkqYUQ4a5
9tkGtqc2W5vpfqWV6QjlxlQGBJIBI/8PjkxoF3VNyzaYGKl3YOY97Na99LlX7tnh+Rz8jQFEFLh4
Ig/ocyM9AWJtbGnaot4zuqXCbIESuXQAI3RkqQdfTtqOKXdWhYI1KJB3i9zngkvaniaS2Uh595gk
mExR73r5GZo14Gok27UB4TnewJ4HaK59RDbincjWEEKIQX5xDCpZu47qoyR3KO7NQGd6RluQmFVj
RJ0rYZu6Y58JSbJu53+o9pD/cfmEdiGgcxOtRJLp0wW4DoSrDZsmakBbYvA8bptKdOtq5gD5H9/s
yK3xZ67MTzHA7MwgKmdc6s60bDpoQJKLft/8V78bCedDH8sFI6qIPHSXEbKHB80yN934Qye3GEzl
1qyMK5BVmEgISMUHWeatGnfvWc0qzYrQlrOHPZ+4pCSvkH1QKzBaEnFKDnQrCGwawvX9efjvYBC/
Z7OEovBiqxjP3+yeOYWoORsIZKsK1rFvkwHeuvU9xk5fAHvnQk1GwWceaESDrAUYiMEDKhVt1kI7
o6zYGT3ShZ9xyl7tAzLxQdg3SRiuzPi4ZxebdX8ryJlVGUO/GZJHBljbUZEozvKdUpFRN89uwgFn
Gjlvu66WjaK+KADjbLgvArzlkdNqdmgWwo1Uppe/TBv15F/o+UPg7xXOPajT7d3PqXxPuIjCm1oH
FQfVWFQFZrUj7AMOb/6yZNgtmqQwQR9YnSG/QWaIbtwu4Y5ZWrw92OZo0bix8+NBQcgjknrnPegP
GOv937t6tzS9PRBRQ7iQQ6AXB4PmoU/y4FTHbdtRVynx9gT7OfIB1ixZ9kW3DApWRjs3AbHMsV5X
KoLHxeF+dW4KtW1Qp14FsRB92EuzYns5738iNRPassPBnZ9007QFWeinNLiVwujVhnOnVLIRWd4N
fLFELdb91lhoVIeotdNFDwiBJTggTYTllfVFLyHshkyLXe3biFgTrqdguVFtAwnDxi7YS7fbKBTS
MplHz+FOtrOSiz0duspQLFas1pwEbuQObvguod1EPDq4JHR2bd4XIMjLCne3xwy9cx/S+Es9S8WM
DmSJDe7fPO97pj50kVFyd7CcX7dv7qx8YSQtnLA9gvUf+eLW81wMiMznZCeIEu7qd0TK/I1h5S/6
EEbSQUiKdKCw1MroIR6XRRLszvEbXbhg6H3jxBAAB1zEu1DH8DnykSqsuWdBBpe8o0PxZTDghwBo
8vJXdtOBDsEP8nbMgqsfcUG6qkEwo5TlWHnrgMRLNv9Y64l1NeeaerEEt9Y0tUEshL5Yvo/ojyep
0WYzDmzJ6aJyVz3xgWWvdrl0GYpAUfVMZFclXwTw08C+9nf+S5wP3Yjh62TRuDo8FOB8wIC1g4Nz
MYwEUMItNEsJeSJXPPApr34/geX4sZSnkC5lOQaiPgVqQ9T7+0IURPAbVtGGkDhqp/Fto5WKpN1e
3dV8e4lIOPqbDUaXgrcNYUEWmyjEZ9f69P4otuFmgVfjny5a1s1YeqlafW6XVDNX5soZIYskUdnQ
IDclrcwS09DajeY3LVzyyfDHi4uqT5YNH4qy1OIi0wBzVGxYo5fgQ5U44pJOkFAwyqT0EkqoR6Aa
RuSFhz1ZPUuj3J5Ge+y5BRJ42puWBbxNnV4VhK6taxYlvGNTD2rVj+9srRjx6Wf0AIfCAc6P/eTM
DfT3dNoxDGYIhb8hl3mISExbOiEZ2QNd0AbUaMcNgUANBGSaGPiff5JjTvyjS1xcLER3RVT2ETHB
eZPi5n76m1tpJxMG7+sEA3M5Af9EonseN3fmfrf/N8hYS2Ef1gCUCa5xZ1gXYXxc3RIqjLaEQsej
Eds1XZ7oHjDOXflFItPxVq9D5pe5Gd5sVZpTm8u2lqGlo1D07Nw0hVkEFDfkBj/T5XviiCcILkNn
OUbXutb7Y87bS2s8R4zjc8H5MuIZ8JkO8E+S0kRyh2+OpRwuDznVJXn6dkisZ1qLm6MDl4u2CO+X
rSnDQFg8LSCanoUwYs2RS49M30AgoqBgQ9gEWDznMc+qsBmAxa+a7aSfnYXsGNDl6iCNm9R/NL6R
18BMnKg0JChmiyTcpQm5V0ggDcUpppL5bEMI4C6ume0IS0Iu2lxjYhiQiuxZs7M9anylFqusIy5h
C9uihZWaqIxU3MIX13nnImeu3ePUAPZqERztsM9FmMt14n3lFtRqlkS3ul/B73Dj0cIVR6Zy7gGP
dtuZ0kiOnbCMFcQYvPXDbfxKyKxeQnBGjLSUBm/R03eZ9ysn5wbyK7ZYezod0JK+JuOhWWop4Mii
vzncVJ1wgdR6tpzpOL4/tfxLYj8uygRT/cwOspy3jCAplIAy7wdyFYGsVcRsq+528RaiEA1XDtao
KbxCpdwmE7U5LYj7pePZzn0dxeuGodKu26vN66zUfmLs7NCRZ3XVIIqJYqV+xcGd5oaQFc0C1vL4
rNlfxaMZByJIwQkJg0qy0fgWtqX+gncUqK07SXuLd15RYpAHfQUKxwQPsVlfp3hWx8FgvwO4h7Vo
B6SlZqyyPzVN+f7Tb1+XnwppYEEJoXxsMBYYyZqxN8+5GwEmnCY12hw0if065Q7/YzIoKxk8rzCy
/BFR4iZUOlajPsTnOl5IlHm0BRQB66UHXPwpnTZcM+XTY9kYWBqjz65eFSdGVk190exq4tVa3LWb
NTSjJW1T286lB0dw4CsKWM5MGQLU/1lipDq6Zj+2XZcDC2g1licoZzzsiiYJjKZNlmgr1VGo3kR+
Ms5ICJ9KA2D0e2mckhIUIWe5nouN2EiveXBgfpfdmI9R8G1vTRv9IYuhzbuIV8+Y5JFwL37nKZVH
Guq05d0PkpFw1dnekl9H6JIX0cYbomK07/AL+9bRTtzq6VVZnd/fXImGc5XGE5cUlMLY1SlkOfN/
fsJR32isZ9dxN7Sd0fyLrMbEtsLKv/ZESEvsf891IWlNM0TTWRfav4y85M75InYsFDBR29ezdC+z
btl+hlPcoqUATd1jl5ERACje1Tu6o97lXmTU92kFftDclq6XbfSl4538dVakk1NkzLbwm81ryRGS
UmmsQ5HcWenapbF9VpuAPrKvpQa4GnMpEEjSNWeeN8qUUEkW8xPsakKbeoaslZSTCHoN0DXCQpBb
OUIxN+bQTCr7YdAZ+19RiJl+mL1yp37rZO5QKv+DwSvcftkK1Fi9Xv9IatrOyAvEbbW1ZJTc83ok
s7+LfgJ39cdGam5CCHTcrXoZApgMGfFlWErGYHK4MaZXdiNuSCCAu3fTbncvgxuH5Yuydx2faFDw
646clAMaFfgpy2Uy/UhEV0IjMf1g0/juQDmIeP8Rqu/JGFGR9GNsFJTxkZQnZuHfrRR3DvM/2j41
KTpiPjD4l663qbR5FV5U+nk+6Y4sCPf5BpO+gmpkdH/4dCklXIrcIvrABMeBQ9VFqXu6IodvNdlW
cql0HROpxDvXqV/cfY3k+NbnqHYAQNRK7Y5F263ksHedBO5ZX62Jn4C2lzGVHGYXEOITNkaJ/nyI
5Yh5lnYFgdGgtQ0cmErYWngyUvPWbTPJv6mNeC9pSka5LSIevxraUVhAJLq98H/+s2RgpsEKch83
Ix2mPeTCpnp+duv79G9v6FBtgB/52ypg978fBGq1aDniJg/0Nn0iJrDu4d4hraRhmkSGbkfL/4cg
JfiG8Y0LKX6y3SqDHoOKltThcPrQAwUE2BXVLSdFkozI47oMW2+zfVp3gkxMvLmz4KcwOYgyAsj3
Xj2O8T48VC5DWTvIzHLtcMFHzxRCc9HkbbesfBIR7Uvb2PIb9fZaAGy1LTKQHi+etVEl2vjJPquG
iUd1iewFpyDKIfGYn73OdDuIeIMdgnZpEexPmr8WyXVVz537w8QueRFVuRNZ1VmPN24Iz77nuFMf
J+f9Xs1m517L6gKM7SAM2NJyYXT2+Bz6gIReIEQUaXSEg3v9h6hlCaZq/20w0T8NgaS5pTA6VhO1
KVXXM3fgGJ6O7O8by61Qce01lOlzmtPfUGYmcIMX4pD1mvAH79io1pjC/lXu2l7l3WUT7HB1FXYe
gpSqjqFf/moXV4UuZ6sJ1aah4S+YGBxeSlYQo2eauwE5d4GTFE4p/iNpDFdnexhvT7d2PXbviz51
a77pDvCWQZAvCzbOptXRdCO++4NI2gyOrGUSV0MADApvOim6TBr+Ze95az1IhtK4y/dWVkoRkx2w
JWf4QBnk/0xTXKO2yen/8IeQNOgy1hbnbRgmCkOjFggh1ud4gAMTYa6oTM/qGuqHmT5pME+Cf0P6
ZccML7mmfwXdzqCRCpDj30NiLw+5WBUiQcuumEX6rW45bzPMzsIsd1VKuiTWqQjcrpSaURSg2Bh9
x/5PYftW6xxDho+Bam9hR6LIiW/8GCvwxUB0e4ghPyRbUTIo6Is3bxU0XrX6ogNoRSdYvxxAM271
SUr4dNPhCJPM+dyjyOJAwO2U6Z1+C84W9Lbrgwyn/iialTD+lVWcfORUWBM75SlqUA849Sd/22d5
DFWcgU2gIm1UH8yk3zIL3jWSSMkR7MtIWgkdJ1Bf1Gjnlb+aQjTiNHWvbUh3mxd862lk28H2sXHX
4COdDTAVQG+rY6Ki4OX8yRYM1EI+eaaOojTaetAFbTSId83rj/9kbDvb0qaB3aSdeuGgKED517cw
JEsPs6R2XI5TpuZ1FUHFhFkrGFdSqcm0D8rz1U+t16W6/zcqdtk/hVXvL1RAlTaErE9N02S8gV8H
cmUnxGRhyzO4igbz5GePk7KNXloy8Pq+TA2RluOmp3B10M7tISKPHpjMKpwObTxByYnCcwFNcZJs
TyX1NO72BKB5UZ5QRjrYsJu5lJlrfB5EowZm8IF7kc3m6v9zZuEWt6RjnmBUVxddQmeqAbRchen2
l9uwzZMB6McgfNZKF0P3Z1/tyIa+4iwvdyK/NotLMpIArqvo8QCX1A+qvNLvozU0yD2ApT387lBl
9+NUMGyvAfPY5QJY9sPZcJhZe1AV2/zq3emXe3MRoxNBgmgzaOTtRvObR4cOluj7eTy46+hPATYZ
baZ2VNIA7CE8OOpiVW5bRhoKU9fWVyxhtqQSzoWhs6ZPyZfMxaIk5uDQlMPKMqcITVhLIfl+gkHs
56142C3gszUn7rm14z4OHLWuBKwjeXzOneXZkiJGVtxpQaxDy+3jhLpYFIanIoqA0uCIyX5yptFc
7dO65c2DL+IBDNcipDsLada+nDa88sn/gjXywNw+NyDGmAs62qDpVj7LqoTJ4x/DN7DM3jquLL9i
eTiEGnVhCB5XMNS+S4R4gwLw3H74WapnzDICxkykLn/Rb0n3KcJ4/PGlTGSAKluz3iKFvOv5sTOq
wTxQC0/JyC29LgJPSgXzW/HKatiZ34bVzpQj6CbHuvMD6JN8rD1R0jTYRUf2/c9LDbpxBBb7e++j
Wb/t+oI+AsgxqYUQQ+45WXPgHKAzY0+jY/ewXiPiixvIxAFs89sl9uDPnk2Qz0wBoNpPxPIlMfoK
Yy1PzaSuffsb1NUjMG6fo+FwVX+fpsX03mvJrxp05jmqto2L7AlX6IFmwL3WgAcmrTe4sppnZfHp
4kMvnqYuoFRZNrLYpvw5a6IGq/bWzA3I6xED97iYzM9UQFQAOYNID+pIb7KhE1z3BGQzG4Cxephq
atR90uKcP6Bb7V+haGb044bZqK7mf31BlA8WMst+vlhH8HgZSJUVOqk70HUbdMjKWkfCN8ksKafL
05DNrABx3bOHctst8uVzqbooafesAa6fw2nCVKUHLSj9yy574khSfWN8/nPfxZTavJkqp31GEPWL
U+OChtmMu6/uTv2mVkRIu6yL1lWERgScpfbJ7kQpwlLAFq5s/umS8wDqr3DYDwNF9BC62Hah+/nc
MBobUgJpScfQESNthFM/oenceR10n70X1u6VuGCLU+rK0T1YTjiZCBjQDSz0v2M9Od1BUmGw9LBo
yIG4+4hQrGImiXHZkMh4/6n1yMb1yIvs35YBYVhITJ6Kt0spkjgp9DnQEStG1IfwlNHdOaX1IziU
YMyxINXhgG0se3s/zM6sxQGS1dSc5zjRwFordh9evpxw66yhp2qc2q3ZjTsDYnGjBdGqV6xYMg6G
BQ98Bpg5KOmD34911u4FfXZKF/CEM6EoOOzegWGYWrdIB3I71I7IpQ/gTFfm7AEGm8DyJe0Dtg3I
mjqMM1KzfjTF72NaXZZeBdq+uASgXwYQO4qTx64NZXTbzSnA+1EozqqjlkoWaMaDhOUt8dZVNSmX
etudMNIWoBABbTwBA34Z2A4JzJZqek88iSThKLE7MSLaGkh54eqSacTaAVUkj9mzx3/dN2s51mWa
oYkwyhDkQaZou2bczo96/exNNYYzfBdJ+E6K301Dor2PPUQ8L3qXAeu96K4TTHhTVRmnz5dJcY+Y
nT11wB0xAo5Uc5gtnkvRWa0prptHbWWk/yFjDYYvdRW83NysHm4KQth93E5I9IKbUSjl0Mo8a7WD
0Wd0skz6Zwmc0J1pLG7F66JgRgLxHXRNqP++Jira1+7E2Yk3CkRs0kbLojAHhhtzKrk6u9BKdk++
KzWsaqyl4oq8VgR5KiAcGIdqqZIvGA049KTXlneMHS0kbQylm/skgjPBJY2desDIeS7dC/2g7sW/
Gwex/C6yKiyrD54bsfhQMzNGBQ2vMWQ5yUV9E+3iW0YnbTeEoiVz+MmW1AMcpezozIGMLQkOs6fI
MxMIMSBuTeZz5gX83jWTY+l8Q2L4lAajZhuU1gRQVHF2lN5D/1fu6BMWNp/X4RQPBRmLi+yWZJgK
HfjXnBhMg7K0eaU/vF0fgxuC9ECU+azUWFypr4Vfzj6BlwKnXfVvGPGW5ltZIbrVa/G7kMmJlg5g
IHOhoPUR204+rMXqeierSS438HJnztKolalAqWpbB3S2faNIncMXlP+L3Y+kQYt/aqes8v+LVoy9
y0up5sSf4jUVernDlWYfAFsH+LdDz8vXzFrxCoI8J+yb75nd3v7Kp4SeWo6HSXERqA0ddYmBOMLs
FGmdWGU76Ncndp/o99a3jVUZypru6yL2KAgOmeGDAXvKt571LBbJQq2WvYl2bj6ZnNOTrBua+nPy
3GPCpdFMpIcX6xGVP9cGvQ/zDi2/wqEBwa1SabywW1v0TTiIIEP3xzpUIkK+GG4rncX8MA5ZywW2
9GxX1p06SDVSc5wsFPHlivR2aqcCgCu2JzNf+Ll1ZOVqbYDNW34LGGHyeCgSsnzXURvi9sVItwfX
gX7PJEAJfADK3BpkORtI+UEYI30JB4QNKy0/xkS6L3AQpPbBejbgNFvpfVftGysQ3/OSGIXIx6rF
w7qwSdZ/JOAPUX6PwVEpE/sf0e4iq9Wrm/nsu5RKKgRav/TWR3bi3mSH86h+s26BE6vanhfd4tnT
4FXKtKMypvaaeeG+yW2iFaEj+Ssj2GA3GRWZInfOi/h9758wtpldH1b+3D6ADBHDW/NIKeTwSkZg
ZNm+hdg8okaRZOjvC8JScebkD2jdUeiv1GViG6BrhsMB+jCpJc8SOlHzoJi/LwUzNkeZ3YxyUmdm
Zh6YutyvyLt4H2UIH4tMgbisMHQjEEZIaqdrAOuE7N1NsV2iPxZm+A/dZB4D66oZBC3ZgF1QSW5b
ICbUOVtjl2ykXeNxW1C0l/IB2KEQxfU1psz8NUyYFhaC7uR7obIv089lXB1vA6MhM/XB83YsIWPE
eYSQRj3BAiZN7KEIkRazieCYj1/GVmc9fWH3goQJHxqTRlKQdSbSRcUSH1x6l+FTiZHZfUdUCFlw
WRcVi6WCjfuc1JjLkcPjmA55crHZmBl69dnEcBVzYFC+Xbxd93yWTC4uJvSmC+TBc4gvlrFpI/pf
TsInikjk/1vDvC0Ub4yU3NvyAkiPuUUVU+tBMJBRZOEcTKIRAzP98WQfxUuXP8voxKwnmsoK79ub
cyFnae2mmTg6XT63PYrdxMlr22IVD8a+EWMHaaie2P6fnarb4URY0Kzzoiawcs1TT3rji/X1Vjqg
UQJL9qaz13PSdc4squxnPJrsi0BDcrIz8J/Vbi9xRalJej6juydymw5ES99R9KKWf5riI+gylOIg
MqoWCtQ8pvz9iF03mh+BBx74Z6tNiVRMqktFie2bgGXyARZjlWCeGQFn1BwsG3qfipYemTQBcWnX
GNCIke81iqv04sQDyzgOxwvSv7+HRpKzH58Lrw0rgvljHMkbn6GP9UrAnN8TlsLVLdUvliW+Wqvd
vNZEBUM0KEOl9El/1kORoVWdzFnj28ciYupROvOZMomO0x3VG/TbNMzUZjKNraRK3CS0/lpZsrdk
hFCEw2qksjjp54gLAUvKWQm+CK0utnT+w2Fjh1KpfmhIwuyNxbBV22eUKYrII11U052OrmtFssdG
Y94cCKJkS5EMlfiYwdU86RETnpUrnAn+lKCAiMi2+nnTDbHbsG2dBAH0p1jYHjrcL2u2vQX7dl97
AHFXDE3iQHegS2cI6Trv1YE67da9u9hiQTdMD3LrqVU1dbdE+PhtvvXpgaCopG37FdebyKhVntBN
sRdtDvj/mbnUIRUsH6Qua6ZFSgngRrm78X1mhF1XLuS2Lsp5ejH1f/81rDu8fc57fx2CGfljoi1g
+mXKDBjuRKrSQ9FhZkGUIdj/dEVwbkJ982MFcKeTid6/LQuq2bdsgRJXwRCpSEBhehlHyZ5PLTo2
l/FBHfFOZ25vIl3txm27rhi6SDIaOxiYGuHrVmhP6mwgZis2+LxKFSS9HmUsv48tnMZgSBOs5SF9
jHgKTU39LlFuifJNSqgv1QWyyJ7enkBJFhjMLEu921WEExsYn1jQ92T3rsPUUT3UgDbtuv0qTgh9
shCUW9IBn1pHCqCeH4TyLHQLE4JA93QKnIHPM7Y4VkmlJfS6p/XSD2u+fFwRs1WJPIzDBUGct4hz
VwbXmrh2P8eKpIneRbuTpTFv8jTcjPgxgF+zvfLns0TG+ayR9ofOhtUa7NiTPm7PjT4Srp4KwvCm
+WuqCTkEeqIzHq35pesEBZHgL1HvQPskyHogQhv3Hnp2SkmQARBkazNNUNmeu/nwAoiF20vDeLPv
swEhnDnPidLkwk/XaaSxUmkppjbwDpLzCQGnNKyQkWhgyrE2Vifydlc6XpjxqTUcYNfnWgxv2VSg
cxnIeWxBqKT8GdeV7ko9BzUJWPDWdnquOesTHdH7v4IXfd7IJNaIzJehqD40JliZbRYbkEZa67kN
yapxoPcAOW/MVnUjae0IqfL5Z6zLcZcxwGIGqTp/VKSus3z7p4sP3hGmvsAGMpkP/+1SQe+l44yq
W5+R+NAvpJp/xGNrJ+KHEa8q0pG+Y6jpxfN489TPq218hXD/IZ7GUMBjeswk10R0I9G/idtIz8EI
bU3+GoW37nk2Ey16aPKD+iVxWS0pcT15zJ2Vl4Eyny4k5JbMAbRfsqPn3aU7dPfifEctHEbh8fz3
kfio1ibkyUe5sYnQyI0djF1MbYHVr/9qO78jfLi/j0SjGgNzoGRYJM6ULzod5oL6fosoxFFZYfBG
VQbG2AbtYtA397U4BzvXEyry+Pi1wz00Mob4j0dCG515QYLajYMpeKFNQbdL4ZwqDUwon1lubB7w
fKY5vdgNUnD7c1N17EDIA0MY7JRtyvYJk/yOIJHaKYPqG/1BNWw8Y5V623cnyPYLVyretq2HBk9Y
vDgcEFyrTyrmdDYho2QOwde+4WmDlX1ErniyDVe1+8JDfVwbxU/YsvHpz9o4SWbC2I5wgoo3itN1
n4pH8chgleni04jCZrQ1oLwX7DEI3iHocMrUaL1nmYVZ+0DWmsC/e5E/c9sQyfngJZ/C7l/kgYjU
ghZo3wEtIeJ9Hg0Ni54cKb3AlGVFm2iS2/obFbVwhbGD6LQ3El7PwiridO7UGGoCy88ccF7zJe9F
4VFtWVUm1+Fm38cqNy2zgE7Vh+SVkdwDw6GVX4T67f9I7ojiQfToSLp+14F+UoYNko5GMKp1f9dT
Wp4S0pjFCYJlGzzLhTEzVSClXj/+iPYlW5kyRg4UnjFog9RSA9n7rcwkdz6UyZqVrYo4nOERgf+F
bSxGogeXaa0Bcz2tlfkY7od+uEBuwsLhFwyAVny7ygIMEi41tbKrLRNeBPi3MlqqiusFxussdlUf
aKMFvRSi/xqFRUZQwbXipJOdXlEuNjDLP565UIlqgJ1r/Us5/iKO682YTI1n1whPumFUh/2VLB7s
n/gzjW/XX0bfwWjGrqQgDgZVW6qSTW7DhEZ7hPIl3AzePNRfF+htmTprbUwqa2arvUaAFRhSflZ8
2ytlaWgjZ6OuW//3KX9eOvNnqiGDI8K2BmcVn3ll+lY6mhsRyDs7JpWlSEArVIKzBpnlfGOKOovX
oM5OjpOLMcObJlqlVbR8AzrY5BcjqE4a2dtwmwElB7bnwp093Q97YCS2Gm+lx1MUmnhg//Voj8WK
ds6CEU5nQgx846mevESW6RN2eDyVoDaCEkbaIwz5ta4XwIqQGGc67HpC5paOpGvO33923Ptoeur7
lJNYt8oQPfLiaNeAFpCYwi7cR2bGmLnvh/3B7+IqzXSV4TrPsdtDSbJm74UVYjYfTREMvU2WcY2O
14YYjwr7Iz3a4kDvF/3NU9hlWCwY+Y5xuA+1Pmd+EKHAeLV+4VG7ozB3qhNJdNJauL3ZeY5dmDFD
Q8tWbNPw6omtf4OwlkY7V8A/oecSSaXqwJPf0nXAMVZVoZW1178FGs6IOeZ2lsq7gb5ra26njfFW
yYZiYt64AlfcbimPtQAOVD4oxU1y7g2tjqHyET3DyRWn2y0Tpl6UMQsWbuC7IGIzMHr4LtKV/d7v
1R87z0fdIShLg8cfhdta6MRaIScGLnVdms6o0X1l4n832UYasmJjM8sHujI/mTRBzKSdoggfSmU0
Ft2JcGlXNQOSdATbK8vLL+D1AzOxo50rYL+nWX4mLR6xirY6WcWjvfMlcETda/U6+poX7Jb6n0cL
Q6zKg3EBN14zcftBZPJRrHux+3j+YwO14CUGugfiArlZZQLPFXJxcIpKcfw5+JiNwUJo30jIgJAr
kwn+49+gBByaiw8d+FV8SiH1rrP5XQ7DlUvtzp3YVzbbBfSPsM8gBDrrnBBBD2cLZ2QGOc1FRKxM
cwdXxdB0SeeKMdYJ1GV+1MRllrwUdb5R8z00VEJEv3RUvIQY7dw2htOXtAQFdKTKwW5U66eYwuMV
6x5JzyHLbkm5Vv65gnUPEPH/kkop3A3uQKk0x7VOZEM4QU2PWodq4A/MzvTAnPL+Z94FH2nCS8dZ
JQvjSzQS5kSTIgCehq48Vc2Eyba47osF1olYuDaGnNrkcX0ZNSiX3K+dlU4iqkcwGSIBUm4GnjJ2
EP55l+ORQ3j8BZA8nzHZvRqZE4qEEy4M9Q6DdmuX8N+HpFsgEp/y0aKJ+ELRU67d2D+LVVdXpbp9
HxD7urPptRw+SKi69Vvbp7mrR7dsltrOYsXehLPin/X0lpWsIkMOoY7Oj7LoXxaew8vicLacMMSi
1IlitBmPZZoDkgU7Zx7AILcVTXLZ8p7rvNNxEpfALC9IsHK9HsP5gHh83G4K2v0h2QlMhIU5dI6p
BNEJcHJ2JbLaawUBFtjfSpvlviQ703oX1HlYnEfA4VkAtZ4f01cCyUiCqo6aLHzC+v29CF23n4tj
MB1Qk5vPs8U66n7BmwajSJiY/eY7YXRiGou1ulgysZnlZ9nhFcWZ8wlnVKrNq0L+wbE7jAJJu5dI
tsyecDEkPxV4aVCVjL8J+ci1mgTvgRv4wdIDL6iKdKmCK6uDHODSZE/yRbEMKWUqhwBeULQq0GwO
UOMy1Gz91ytbXaYQ6Ni5JNdY2SNbtfsYS7VvriBXhkCccaam8m7aLo2DOzAXbt/gbR9czIndJMI4
TjK+WdfgvioyAm5voSpnrxlA4A9ROetq+EPVVHDzxR9ZYdtoettsBLekC59sxvL3ww5GxsNbjbkK
tFZWM+398e2Edy1AZb0DYj8Srh5ZbIL51WCRIV4Bo06QGDQDvQ5pSxJGwyX2+VmG2s3a1RI2skDZ
8xIExU9/Ev7XxPDqcrKEQ4zE6uMol+tTVtEx5AbUE2n+u98SIG/Mn+ivxDLEfzrutCz6vkJ18WLM
cf3/3FgZYLddody7ECQwjqyBsZQS7HeUwOpAqzxbc+GgVgrYbvj4jskixXFRR2oDC+Yxes6hqr0J
jIIXRVOqly5YgeX5cyzKTD1hmQOMnV+oMfTRJOdvl9SU/cX006GS1Hk6a4aWFFuvn4HYV/Jzn7dU
f6CscLALSvaUQnZujfr7CEj0uZsAKcUI1MYjSoazKEAcD1N7l5W5rGWiUrF2yqWUYqDQqxgXERlf
QaTL+IZM5cgXSWLORHTGM6Hqa6v1ZAqQeSmiBlL68u5uhx1IvBcxIgd8W30cHL9//xrnLrVToNFv
ZdaL9B6+6Fhy6hCYfg41kUwx+DissrlmZwAhccU3sDR/mLzALkyz91UoPYlRq9fxs1sconB/GV/1
/JmuzwzNyJHyeDMjkoxs/fA8/eR5a7atR/cEHfwK69iKiHxVFUJvAh7iOjA9Qh/mJSO5XQxlr56H
T4h544S8SFqU/tnE+ch07aV9hqS5RN1ljvQC9eOO9E/Mur/zsLZJvKKPHh/c6FRixH4+R61fr56g
XUSDJoK6R7nZjbBOIfzwPPz1c5sxW7GQutwqjNAEamEOAPX+25yq2ceL/KX3SiK5mD2yqfpBAX72
zIlsKln8UeLp6iOv0IjhltuuIsVOCt6+bd7OPhkNUTbpVxSxNuvzhUDhs8Ib1bY2ky/ZfJOlhKMl
+l4uX1XVZZCRRdO+4+EFMJbrT9bkWY56Mt0hj3HcnjAR7tvKO1TzLttQN8WJrYSyO4LgMSEUmzri
Fo4vGiUTfRVbzpaWwyaaCrCXyf6r+QV3adeTcWk+uofNVjIsGntQpe10TQWDGlZLxcE9xGQFblLV
BzPdiG0g4iI3Bq/VCJdBq7roJ21tFYYJREXJRoCt4R+Jcqyh/IYix0CLwVQjdCUyiKCTc/BVHNO6
wX83e0I6DElasoMS1lhRA75Z7nLC/Diz6C7X1j8nWSCamnB8zJZlxhNbr0HsnZ9HHidZ0fUw2boY
jp4PjDvlXSr9P1R1S5V8dcaezhJLbzEfAF/uJVtcNxagYn/y/JG1hQ0JWR45ZWvbn2V5M41H7/5l
EE1jCpyHtB6FQsT6YCZ05h3Cd/Cu2MwM5M2rrhqXeZN1EGuNamFenesPD5hQFVJLAFjB19QQkgIL
zmeto0d3D5UT6P2qytDBSExnVoozW3ZHUttxiGXzUI30ENnYqAJBtTjh4Ef2HtQNsOndlmr39Kxt
rxA552Wyj1WK7kmXQiSr+7VmhNbsx4alDWnh2awRz4U4HbMF6pkHGWvPPF5Wbr5wdKX1oRtw02SO
6tUGA/1pg3j4JTQ16OhaeEcuT5UW28j7MzoWu/JZ2K9EB0d//QrFh5yzaSswE2CGUP8sffKfe5iz
vRuST6+nXSMX1EI2UOrWTNqlwTRvS7Ez1+e/GAL5FLBHQLjwhR4EzeYlNKeuyJsZIUgIe+lICe9P
55ljtWWqtLwmAvFh36vqlK8pJhzH8ocbCNl0uuMDfAZCi9yTt4nfq53ivo/8EgnDfyh+2oq7DtVA
2bAaQd2V3HBYiK/hLhw8J2ERqszfYSEvLwvd5z+lzUDAVYkB4NU1L6wzDJyz+i9OFeiR01vOtZMk
wWH+6fcRyjyedivUMSHxBqmUSeUEusPgzcCxoxlX0i2rPuQafgKJd1kz1QN8u0hg3tcJ4NA7aWc+
0S2JDraHOW4pYvVdQ1ZzGeRYE/PG3zUkqX1Dc7CMoThDf87rPejccylzpMVENNAJlVJ4lJWnlmas
dGAaUD/g+6U6Ia00RStx9scpG0NcRSQBVDN/Xwh8OvcIy3Y2NFRw9uEJG3VLlv+Zh3mpgbSVDaKH
vsH3hF7K1CQJHHS9cgbFeALzoKlaMDxrxTAzR8j4pCe4DcsGuTngw9WcDItvSir2Hd3hZ5q8SMgo
FUGY18UWSOjGkVD8d3IR//diJeFLUWuKTJzRKdDBiA9C1h4d/iH9JoGjD59jHmEevg3hMN/maD2V
NMEgOljLDSjBVe7uHE+mZ9duoiuMuQ7DzfO0Aa6hX7X5pMIk5+M+wntknALq96DBBMXdIjfDXGHf
ttI7LAOJxNhLcDEQTeIqU+VSIBPYfCV71SXv6vjMvQ8NoIk/j+KaW4ebx4IM0TjTP0ogyRsDlWWp
N/MMSyaJF4FiIcJhwNc5tzFwPcjPCVbHlL4KyKGlcdDOktKllksOgczvwxCIr1UJbZioswULsXkE
fbWXCCoOI3DcVmu8PKG4kpBBUFI8XJjGRavpgXuKoyaB3PQp42bMnZq/nuVtPtc5GkmMN3T+76zM
2JuCx7iz3TC0gnGvs6u7p5+S1kfmUdwKBUr2OtUpUvlIeF7l1Kom2R3LRS0rn2AJ/fSFdnDOahlN
fGT9eSok5TDR3fK7gw4hIEXZTz0UQMaViQWEQOPhSnlg1ltbI7YyTfLp6Xyr5FpCZ2NesbuViNun
MVnHixJimX7a4eE9tv1dC3XuFxQAPNfmFjmO8xa1bP1+roYsrpLAYAfm7pHX6pWLTUBvwJg/ct64
tdVh6rlo0gkodn66fwncTISn5tTeMDyieojMTofpMkl+dcOFCN22zQePlV/4u3x0h+xG0CM/rWZc
QGitEII2hshssnTc0s0FKKrFq64U0gQyHu/ZGxf4qLvrtcgXYUDLkiXrcHf0Lj0c5DbqJuCayUAm
GgiqV8vuj1gJqCw/HAgqY1sQKMSoQbCS5lWrlBwWJbMJPlfYAghZ9sfJIWDSimBucSpuXvcgDlhX
DilUZ8euKqgBFZpihjwaCUo3PPSetPZUQmH2VQ54m1J2hdhHuQdwzUNhFLnOgE/v7cHLwtDM+CQ8
aSSRCM+DW5eG6wHVoaf9vqjT/Qv87Rahma7jMXycezXMaUwZJ3JiHsqMajc4YRHoZRuFHyGn9fa2
PQyX8G5EaYbpxIALIbcxb08d+HU3eZdrkrJaBNb2hIe+sXlHxgc6iJhm6YsINsVCSfaH/QKAlf1s
aVZpP/dwrLunsU9XynmhA5ZMKax0IP9dVkQcsuJA7P6o1gvmsmJJkupvzJndQLtg097iBiJX5SSu
hjIiUI0dJVWofrdeE06XCelP5+7YPvR4V/V2nlD/kxr2epH4AgNVZ+68qDzAmYobk0DNViSISpkF
of5e+wCjo+4lZQOH8Yn6yHhEISrp2MYuaQxVouNAOOwBUTq2vzdYJ9C3pGrxrvHHKm+briVEaQR6
cKf08wa9J739K/1d0bUIsDFVGppJ7KduxXqiUwN5c0nkDxf/So7JYBx+x2rfziZG59oQ7Gx6uSLk
MrMJ6PVA1MKokvgc+PV8sxXg10duFUBhNDIbNYv0PvIgZpELtoV0taOIzLgUiL7PkDthjpdMiLsZ
sCe69oi6OJPZ6JC64fhTdXpTvHZIQfEfsBZpMxE+F8NNh6ydqrGYKZH7FY8Y4L7Ex/cA1+Ct3AKQ
wY8Kz58bVKSMgEAHozFsE+3AvsECxP+hBp5RmQEdiPsMnHwQpp4vPtIsvtHpCoLMDjC2Cpu/oyuX
FHvHXM1oIci8StE4TFuCDRupNNdtQRCR2DVkKrtClLcGie+SR9G46Cnpo13DsWryflsJ3FUFvb/a
0q97LIhuPWQyGbVYw678bAbZilY/K4aB/2tlL3FOLCRMKrTzim9kn2GtFyOF22vS71gdHSybeHk7
WKVE9I6JTjeBvVP/DAZnQ5BK+l6OIBRZLYyhIIqE6pO9XC4qQUoo5ir0dnoedUNtTiZ6i8R0KGzM
jDu1rq3IVt+564Q0BVSz4Wsf89seWzAO55Rra9r0gBGXHrBJjS2AW307BzvjlZmWE1GOxfJZr68Y
h9NrBo8DlN4Lghd3lhRwxE+de9Zmhs4MIDdk+EpC3tLhaYA6A7ix9owrFQVqiuVK8UNGvAd8V1/+
LdREh63eyymc9p+WoHRgjnT1BgaVX2pmEYMIEnn5Uzmu6wGtKLUWqMEyrIp7ph1VNjdkPQR9mryp
EWcEJSu9cbjuFiYMY5LjQeaQLRwNcaYZx0Hq8nfNW1ya6VEOTsf3cx63jihW2YLqplq8wNf8m1ZM
4v4Lf/qEPwC1JLjFnVyqEnwquMtHuwoJufREfKNMFvZT7oLXxMq7Y7Ja8YYkCb/cYroT10mXWzzY
Wmnuc7NqOOYt+gz0HQbR2zsvA+5johXI+Y7QL9WxlhmUvMEa6GK94Kj2v+iVHN8Q4iQ6LP0i24Mw
uanIG4Ol1tLC2KzyR9QyG4EsDCAxKzY1R9Mkeu2ngaXtik+MB/Obj3YSaXd8kvKZwJc2KTLLwvee
/SLEtMYYV0wezlWRgYY1XvlxPsVrBCx54V2Ta1SEFOtI7JaiMC+9JFegX+OO4xUNPZsyeYIrMMcR
n6o5EZTsIgXeOkpfN0CdLYzpJ7QcDjuCcaz4Q6g9dcc9nO+p7VZl07aBEn0MIaMdfZ3Bf4dIjatC
cDXxO3cukuvrnvgUv81GRMBm6ZKnF4BgtqpRxNBiuwaArQJ2HVWB1432hcDL1Q0idhd54ZWbKQuo
lRzTIYknk0uDK7pgZ/8JHAc1B0eiUC+wijg77guyrVy5wtXQI2FwYBol7ySEK/+Y7yvcwNdRnpjP
NzCQwMCqhOfWrchOIdgWCBgEW4KY/H77PmMp8TVn8LF1A3eg0JK6L2wG9E8GfbyC9JgMu4Ksu9NU
j1GV1rqPF9vOH9ggNFAQGJeXZLhoBuvZYNy1zh+2N6KkcW/AjuMDGsj6WAFiCtogYFVRVBk50ZAQ
sDgYrwMCVo9eaJdOur82i20Br2uRyq8mfMt/yyHIb8lX3hjI/EUBNsjTiHsVVhS+j9y4s6DEazGf
UOgcMehsDgvuQJEgqeE4dA+zoGIMp1q96ezXnbyAkod/h2Kyk8afq4DAvgMZyFM2THTTJ1zFUr3x
RzAjFGEp9c2OrCGOvEvT5cfvxlyuJZXVR+dTv2KqsSMNPKynmfbCdbEqZS2cMXQ5dcsIxscHhy+6
FEUAHY+9HxXQVmX/cyHKI3APGUt0VJNR5MTlW+pXwk2U27vIHGE5aqrDQBZeoiXHeIGnkT9SadfD
piUjsT6k1A8aebsU7tozEdS2aQF3WfQVu+0PWCZDjq9ZiZ7x/ame/f4hV5efb0Q+ektjV/JX3zcz
0zCmpiGXJbn3eUiKZvGWxgtAaksPuNJ1uIEG9O7iFJ+vuwPS9k5OBANNDKjgF8amSZCKW9DHU5Ca
ju8TMxGSZuxi7iUzD8ReV3FZzevWpnpqj5yoE4uR0XceVZETUdGeL8GuUkVGVGKoJfa9aW0S4jdh
hFp9LhmzeVFsA5LgY9aNEnzhbv/ZQrzXNs/32UW0Q2tI/o3/T3uenVkWhY+xqeBHqvsPoLxomrwD
JNTxzWC4Wk4trdkYhlooFJDN/8aDLXgCAxivgLDoG1yBEHKh03VlrjB0Ysr6XNffh6O7tEu/ONac
wI6M4QXbx9jtCV6PgRLP0OrwNb7H9rrjqjd4i7dddMZJshgclDG/38W/ruMOMaMI0nK9/u0TIW5r
MtpqUNL2hZJqj5KagDt+hhlSEQxknaMPI9ReZGWxoW4f+a/g3oJDf76srVVnfrKJDfuE9EJ+rihe
aSHjd/9nQ9IjGdz0ZwZeceL56ZZmZfGgrGd8w5gWWwTL3sIOY7iW8Ll0QCkEvhefVATKh141WPkv
4KyCdNWZWN8e8sxB5vPEOgF4mB6u26NHcVxXUTNj2QgNSFYCqgjD6v2bfdROU6ZOK1gHOts6SvIs
Qo508C0WtfmVuLcVIDydPohnGZqJ/eUTOeA5dbvsYXtbq7FkBRketrNhjxPXQZEn4ojNPhDn5Qda
+gWt8wpc5wBqcxo0fsgVraqRvIW2YRj0kyEQSUN/ZgjHM4L4QKtxCpbk46/fUgoquiYPe1joVuRQ
VL2wJElr4ie2fHTuhN3EGtpw8WE4HcJXk1eoe+Z5TNtdgSt5MBFEQztBnbi7lln7QsMAJZEx/omp
uWBn/swUqIVngoVCeHRUo3eqylVhl+heu8LNzsglw9pR/+103eFROqrVSlnaf+QhH7uM5LpmWne9
gQSRnI6F6AmcZ9zCImikjM+WHovSH2xd/AQLEyCvFT5nCePwiyEQ+GryTMVmaabXmuHp3SP+Tvxa
cPs0ETn1eBA1KvpqDVNFvVxSb+iE0y94LE2fInC/TEehFD3BOJgLC9dxCxREEwo7YlAwWbUDe6XJ
Cm5xMyE06bWumEF2gnjwl0XWjWqnspZNJBU2i3tccxiz0Iq+4dCyToTVpI+lDzXllWIDSgTskZ0j
APBzvT0d/LO/83fJTvQTrReHHRF264IBhqH6d+RSrxMSwwXQdlAPr7vxsF4ug3iJH8SvGJQd6fmJ
e7nVRrrga7aI6fcYnaEn1v4OwvsET+RgoAfNEJoDMfxrL5rFsGRW+e6RcMB1gKJhPRIrFIiepnBn
1jjD+cwIM6jF5YkEr4P/mDADgHZvOinZIWotJ3lVUuqHEeF5W3nQUfuY4TeEay/Bo39/EKDpO0A1
Yk7MTT5qHMSMS8xKYnOkhN1n5wRonlSdFkRG20ExgKCrQf83rsnx3sHmqr3yV6aXZoUUXhnS0v40
QvhPJ6di2CkQYRB8HfOtTqEbyQ8+HS0QMMz4mhIX41TR9Gf/MO9lC2f0P3CAe/ZbIpm1Bmy3PwTB
ZBI/+K4ppkCZgwnWsUSJ3Xcdg0ujE7W0sPTtWhIyUCT7Zu9VDgUx5HDrU23BpWqHvRGxJRyeZCyD
GyC0aR2Jy7BwIaNAHEFM1A5yBs5kSKSZW+L9Af13FJFnEg5XjeBJ1j4nft1jYsodqzdYRDReoJ+5
GylwC9fTZvjV7woQavh0FMGmuqoaR0acUn7t4TOm6OeuAxaAs5B6pjyg7E1o1cawv+yEnyRAOzjz
3Sdsipm4xbWukmzPbsr9tCp4vw0zwJzY/zxipt/pCV4bJjDiz3pENFLz1tqcMphd6A2XhM77/4rm
+us1JtS9Eapru9ch5cFkfBcx3Y39ugZm2Xh5XjgddZ3l68hQKmRJ2hfVZ+UCBQISzx5enbX2dSsn
qelBFsCXCYOu4IPyOqn6gR+I4/bose59Dtm+EFnSxJnBZ7ilCWf3KReUc+hOOnOvdT+eqPTEi93D
CF6SUEiDE6Lj0dGgb+cF/cPuplQ1jkKZEWFqxIg+mKneIxfiG+OmxoHqcpLzz8PjmMej1XcjiTup
rqabT4dSTNwctvwfvgemUfaoZdV/lN6tKebMvZlbHqRw/AJnmpyA6jSk/SuPvfMFjoCpxx6iQabz
GF2AtmrnIUH9v3jHZItjc03PSe4YCj6VN5/0vKMywmpSEMrjNS1AE8XU3DK96z6YBHweNTyW5o0J
tu8qn4w7N2pPuTkN+Ubc0O2sQxjmigPwfeQrqqzHj9tMs87JJMi9L8R5G15cS3o6S3jstuj2S3JD
sDBcI8BqRvF7hzAsODL/tiK51m57C4HpQjMoe9Dspsb4H+XfBpW112zQgThGdQx8/udqTFIQtM8K
DYH8cnUw0Q4HV3Xc1qINV+4r67d5d1/jB+jldVM4PIWJDuEPliObA/t5b8qqEApaiuMgRWHEm45B
fP5nS5bem0gKjze8XVlcatI/HQ2NlBcdYZQMzGLT2yj5zwOqAWqSCwJ2LRmLIM58seh1Jvx0uX1d
89YSSsgJ3r/wAItf7T4L9JBcE7wg79HF7NNcH9AR3a1nH8PGtpVLV0PYpJF7L19wPd5vsRqOHMpt
cUha09MD5ga8HzIisRyGWVItsLsJw7mK6NDMHUnUZAFD6SEQ7wxt0zb6xVd03zR9hWAYcSmMRjwA
W6sqA/E1aYQ3giOhUef5Osr6hGiodU16Ox8GN0++ycrc90d7GwTDpkZpqw/i3fujCe/nF8kxF/er
D87bmHEsKXDA0JawWcFFCUrW6evlL8LC29mTExbPH/lEptLBJPGLRFzhqo+gSemn5/Wo0QfKTMKr
44FjERBHcsVO85NMSARyb01mwQrRtf1b+XNAhpFsJfw2k7b2oH1QDGbeihObDxNgocmD7iGSfi0E
qNeUp49J+mve18HezibGo3SrUu4xyc42HR1tIHPYZql8blIQeadT8LyzIUUsk7H3DWi2f3kPl41g
g4sbVHvpvGhJK7Q+N14+XInczhu8kipobE2d9EqGWWNhSq7mPaAz3+fW89Hs8Jo23TubEY42t/Nx
7nV0qHscUNCEG+Hni3nwUeRJ3Roc0YGRmNQQzpKc8zRgaETMQtkGniRCJ6ymtNE2T9xJBiq2a4ur
V124AtXlI9osJP1Pgedc1vnBP5A4pc62sIfuaiu3QYuaJi+kg93sNKpzWbJh0xpZCrPu2TKqK+jv
zMuBHqmHx0S9sx8LZct59tWkg1G7ojuMXXMxbdPo9l6dZN6ahxvjmR0Ec8g6SgH3cQrHQ8JeTdIa
xTrqzHzkQl1u+ZM23xfOB7K/YFRMadroaDt34TgtliAfDPmafQ2zHa5JTK4/4AaC1sF4VXPMKL+5
qcGQGRxqi9Dwy9VlM7qL9QtFpK4y7b977zO89gL2ZGSWFu6tZX3sIMcxsKiQ7oWfCuMoavG8T2JI
kHTIxrQnBYQpb2ojofLV8CtBQ1G0BZkA9cMvHatE9Gg5UwQGsvq+UUg1dLrcIrjVxYgOI3qPLhYe
tbaaCZPysvky6/SutI7es2fGxD/udwlXrXs0I6GFe9qGtdrA9z4lpaCQdiBtFrl2N48QVvucaAH/
sJAuLMWiM7ZiDlWuZ0Sj1Kko21y1V5G5muIOIrd89Y86gC/RZB4iUZcNLnq9F43iJlo4PNoGCL+q
BiDkSvn7bk7n1X+x173TQg7ECDliMOvZPlFpQqxZupWgY+weQnYAanb4n8+t3S6ZCRjteTvNtT/s
yGH1m1v/nOoEGyVnUulRulNsp3wbHRACbSkzopRbifilYgBS13gKtECunrGW/sptHWO7YZiTKfvr
1ADg/9hGZGPQkJE4pg7PENj0PIr7tSDrRZoTw17ydiXIf/EdviDtlBrXZWJu4AefwOG4WIiksZI/
ouj2I3VvGqTJZJdw1Qbg7W3idHgmt/XsCfZfLDKG9sGCs+4RwE0mIM5sTSyRg51TjxAApL0m1IyG
NbG1GGy7gVUrJd/Kd00sMaGwdNw1DrYMXwmMVlJTpFy08pefX/tjedwEFlN/cV+jCwGQHQBTA3I6
QP8vZdcmNPDvP5UVUs50/XAOhHShNAqWHm6wjpxZ6HVqFA4W6Y7Uv2IOEJD25mVnfdzJZW3laCL9
ADF6Ar6NvuueJrToqEjDBKtUyrOF2Ze+w92J9YMHWiyzr8XJpzb9e4Zjnxl5fPAyJIj6VDHfD3Hr
Ry+SmlK+1PPCZXmVCoAuW5/VR2MUc1QIHTjG3KE5wH2IGxGpHRpSaHRQl0MsQKdNGi8xmPA6QfzD
wb1zzFCZGVGMmJVR97ss+LtpBLO1JhAvCutsnL1tukaFxaSYFlmbW4p0Xc68QLn6Yd1R9/8ZElxG
4hwBa2w7/e9SDCUh/ivjJGgZqgg7KhUP3KpLF0VIe4cY2gcrK9UNt1gg5f4CiQFQPONpeRRUjs/B
cuWnEhFO+zG5Mu1y23vIJuDF/jqhQh3q6SvOlNjETV0+oPySiAu4KL8F/oF8Mhm6VcAW8h2Dfv5W
kJaOK0DqxFxHjCIfCtEmI8FeWuN3+/iyYEfzUBmPzyNpzwbBfcV2IqqUfDvM4QBpW2EE00pVQhbh
v2xWcdNaIaCSQiJRvanxfIKm5XYEEXNf784jMH7LD6gtPrXtdX3MiebMWi2dtVD4f99whb7206Ea
Ni8+skasWnb7rujBfhxY5UQH0g868v2K78MvJIPQUVwpCjnOgeLrneAo3hcqFzeTx/7Rh8UnAvnX
QwHeY0y98tMPLa78np75jE5/dmZKrHQMiOgyAHpFfQ928RY1WEecF1k35rpUmqtNrmHbe58k7YlE
g5CEa3okLnEJg7feaxBK3/sSHpzMV/6e2yBGutg/Xb5ZPIDLTu3UOnABFZ4Lr4kvrX0aGASDDN/n
PjItU6t7/4O0ZX4HnuAyktYWuxObZBaEVHsMm1dxyBcElsRfK/iBSHtY6/qao/rMRW3JVmvSq6j8
jutdBoeSIeKjkNXkHeTfkwx28dCiPY18/c/2bVl+53ZFh5T/NXz9oF8CojQ3CFCEHTGwelPxRjna
Fj1oQKbxS+foHGQE4s3lDyzeFF40S58UlszpbROBwcT6mErQVAIG0FZcto/s8bYMOGowbEfHabGm
x0ZbFbYgh5rSvddYGgxJta6dIVsBfd5DR2xWKtcEf5HPlZ4FfcDIePrNXmMUPuB9+Xp1yTZPGaEU
wDLASSC/ezYOGKe0tr3X9rPh8SJmfvjlhi0m6GshhuEnyMTSgRWSIcgG7QRJKXIlXqk9T1OHgAJK
mhmbmmrVMNETBvnUXPlNQQmI0ImkXCVn2YH9v/Xzl13iC9H01fUhy1PXOvTwPpCbwTr0608+pOj5
XgRRvE2z/Jo8mmXnv+YllwC9InhN6E7Fd3utTX/JGaHc5AYNTAOlmxIl4kaEc3wdniQw3hotQ1Ow
ts0WKb9Ju6JaFYidYvH/plkRUBpyL167KqFddrCGK9yQoBjy4bMlhhRdlBIloRoyc3IN7a/o3/25
GWYOumcKMbB9Kax804SQoP+AdJ3gs96adian0mEMMTbhMNsf9+mFwA7J8T8rJ7+ahqKfvoqTdMAn
5W9idZfKF8MFSo9SBs2elyTYBpeqoDw5v8BE6fj0z9pNda+NmCpd69mVvPd/41P+1DwEqGSfFQFm
AwC0kKvXgCAEpjE5r+rVcv7lVaBKiPJcLuwidIuo1afwfzcUVGZ4MeX0AnxCCtURuXT0wkHHYSXW
AwZmNZ/9rm+qUI+QCwpItfGfutA92HinN+P09reTdZB2S/fO20ggCrqnSRNuuDA+XFE+0P+1fDXv
JI00etDWqF6xhzBB50IDP/iYFr3SwO1pJ/NoTl7MH9jTxL6emyNlUktTPdHcslePFx7H0q4cfhT7
As0S2z5Zo1OAVa8UCPV63CrWBFRTuuYZ3Zow1o+W5HLEh6JxCVWGiLYxkMn9GTMpBow9+Hhx5kQq
bONK99W7cbrqJKZivR11okOoL+Fp3aNyuD2/lj+gwuhtkuUh9Jm1t9u5RpMf/bdkTPCwpRFqTlCY
UngGQdM4u+1ThFC+8xHNAoc6T0RKG4FqVzDHayazUtRmlFh0Ly7gO0wgUWYp+IgIMyZIB8pbTjtn
Cdcd8TmAk7y18aszMdvKIV13cWErrpy7+ciqaA2vBp3J7YL6fYRyjo+X2isbPvHZHPYqPiCscLuH
TAbE77cT+0vEXgOhsjDQzVF9ie+/LmjfgmgX1Iek52Mxq2XrZdG+FNS4M3d8WmmUGQlYvSPKV6Yy
HNSiOYJJuaAunxgyKEmneowqWH/FycM12wUQk6vgBMpFpmT/iGJ+pir47mthydYZ+OXpUqKFgCAA
0feTzCHdngttw5a38xESRVs60HAvpfNW+VWZAz/mwOFd89m7wGO6fV2dsYunkuMx1ZtNArjJwwIB
AfjmgZvmD6n4JtANYGtZNeTZ/n/4EAxTfSRtSeePZ4+I53PoR6nZtn35TeLS3xICmxyTXzMTmU3K
BwI/sIECMrQ5Q1ejoMFOB1iXHbPOql/a5zJnNyZ649lSMRzC3w8tY+RYMiZcPzDJgTofq+HGoqec
PPlZPMcRB0IaVhGwjWqgVy74UrS0Unnhqiv5lWn8ALWVmdhcPPmwDQgxyS8E4NPrC8wylEf0RLxB
+Y4E5fMPqKf2AN8AI4BG6K0FYrZMmY0h69kwJPZaJOJs0CVSxD3xx4gDB2eqOFwTjkE9wtoLXJ6e
FRJYpG4E8rpl8eEWbwRfjmc7jCGCTfhiK3baQ7mp5RlXEUwv6TQzD6aTSZBQ/JhzeopnOm4ukv1j
1KILUUvSBWh1PmKo7LguFMJOMkE+5FmScbdFmqNmmy5YQ/4e09bB+e21wlU1WzUz6iY36OnOJXuy
PTpVqyrEggJnUMOnCqB1LDw99BEa2XLLMNoPwFMKUVLOtbW2jXIGSwr2hj9Dcdcuh29tTYHo1eKG
8oaNyIsR1bRKYJQcIrXA4jfcr2ueb4WAAt1TLZGg1mT2RfGJPpYIx03hDzvmgk0LQGG4BNvm9HDD
7xGI5eXEVKX8YMR8JPPL/iT3LGYMklJPIfOOhq5XKkhQPByv5VnUKvI0Elq6RZHsbo+YCOjJfdx7
E9cqxcGWEdkDSpAPG9LMn3Uc7i2yT5U+UWzANHmGEXczy4P8+MpC55NBdXg0b8OlnkolU30Za6ZA
gninRDkl7THq/qXSseKQkAXBJr2EQRFO4tGfRbpemyO7Z4kgmR065CgG7g2oDyCqbMAwVygjk+Zk
j+OyqfPAVRxfMTKFLl7s2460WYqrNu8KfbmWPWUD8sk5i1vrP5vYY8omEtGIScbqOkncoRmk4wN+
yghwnm8xP2TGl7HQ5UW13+CfqNZ7NtsqNyM0HkK09dK77WNOGSUHDe9N9LyacXJq5114qWvn5n/R
hvVC09c74Hn2vH/OU4FvqNsUfNSKCLyX1qJIEDcv8MFM7XEV8/IErolJ2GRB4WTHEYKRZhYXOz+S
/4vV62y02sJhG90Nn3fd1vYFr51ThBjQopUwQ4VN+G5uzVBySw5c9QzMVJVr2W2LMVNq6hfVNqke
eIw72yOc7BwFayHAjTyZkWkUKI+L+681Svyku7XLAAicwDmX2/LgrBZ7AAPMpKkzp3Uq0bzc1/Wy
6udwXnfkcmr3JmMu6eCoZdkJC+t0eAda5grBQhNkf3LrhiSGIEJyWws5QBYage3QCqezIwzwudnt
k1XpsVx2OptHzwVvjv96fb+sYR+bEqC7/qgmZ2fRdg8KSB5BdTdK/j3yaMiL1IymGu2QxWc6ecyC
abMTn19bhXPNNOBuGzWXf8bLOSZg3XbnCdQ+VLdDjhgMx+H52uIpxBGj8t1DjCHt+O/666QaW29J
WKYVJ9P/wOF2uRw/gDtcoWb7qSdtedBaERnP2tHVtAcrRNn0FbD7O9i3FnbPNAsyeanBpYbFwu45
5zTQoGDL4POrL4AKvPq1OcQg6sD4X6MzJ5ZQ9uk57ZPZpbmUaZxZ+pLeoWgcT8RIythRmIbRP2gt
X906d/aSpWAKCdtkAPa7Qpem1E/lW1wfzXaBKtNP2zt9RCcH8FbCcZu6+tqSbRKqRGsH6eUhpOcV
dV9VyDi9qyDaJnrzeK6KW724QqVMqErtS/JN/mokH8BPtlGryCXBZhG8iTuK/D/yMdWg8A8zjPFN
5wizePZ4nFlgGmzowyAA8GUD6m3PaOCx8duBIuAOUiNd7TtXKi89grLlAs317XkbIiNSucKp4wSG
HE9oUZ7cUWn0rFvnBEklJABU9V4rsyC5ojPeASoN7DqWGFWueiGOP0O5eiTOnen7Yfzw6823QWww
pHEb0lLLd2snM9nYin6homfyBQ1PaunDrUJSLkn9I9P6pqgYKpUKp7TfPj9r8IFWpl5flbqUvhuQ
v4OBn84JRL3wBFM6kSo5jtTcr338LJSVbr4pSPgVREiK5w/JwBwg1yC2w7r0GwXflS28xAEtZ8IT
QGCjcz2UnawO3sEUR0esnfuxSABEnpp6qfQucws00sXtiRcfI06iRfVSW8MTUT/mIuBnI7oG3++H
XYpM9yTrBdFY8g35qc2g6aMmMGPnjpOFH1B5EWmyzQhK8A4VNOk2FBegh6yy739X9TXz19VX1zjA
IqnrJnlgozC9oFMlSExIO7Z7YZPix9HbjtzGSydZiJF0na56oMjAiK3HGU7KmtBQhxdLXT2JgmgB
JZjeUd/e/mS1RkBz0ftWu6AOgkkvf/l87dBfJ+gd9B3hnIgeJEA/iML9sc1pxn3uyoVeY7RBeKqA
RLfRDC+iqa5vQWY5Q1pRvjVGlOAYb25+Y8xaqo8GEY5+huyHMpSMBc8o1NYdDHGCWuwngnWNVOAa
CyfyQfVPb90QPDtAe+MN2lZ9xD+kIPGXqBk974BgEHX3DjcHcwRkND6ltn08wPoWRWPkFfjCToTK
oYZBCiqofIca1tcFXh0jEnaKvA1mrRA6cRMhXEIeHYNDP5Cv1gT5l/GkN4dYyrKeKb/P/8HmLHja
lMDQs4SYWhQ4N/yR39qK8L7XhFJkjlVBWf68aPFZV6y82Yzg+BS1my5IPOL/EnuFncqle3rcilDL
YzmAsvBj0XyJ+z1oR076m44UdgMXz02HSO1feRE/kXURq14iDZmZlJPgS4XiITQTKSDZXwy9nOAy
n1SrfsaYAI9zZZqmnzJL6Mk/aDyrQFu6UK2DVVGGZOOvYCuyxpvJEJn5MbOv2KT0Drnzf3aEGVex
yuTOKZijD+mO6YOXAA9LC56lbrK09yWNrvfsGx085lKSbArUEHF7ToZSaUJM4hMtnpbt4I/Ie736
KthobVk1jKG4w21bur3+CDGiVLai6a+I13ByID5ijW8uQCabHbAywJVAAINecTfCAIKWr7VXm0IH
xbqsn6zxfMgSrEwLZqsu2hp4/f1CtQaU+RF8sV/eCJBQSOgnjAdksfG9syGMGk8vInD5qgGZTJRv
SDdBqmOP9R/GFsDvDobGvSRX//jt0YnlPrNrYIdeL7v6wQi62GPEgSnpxm9XxvSM0K3NpHI9tslF
Iccagdkmm8m+XTTcIdxb2IqwXkq65ZMnyJzHNK8PZM8qp72g/nZYwsY2l+AqQeWoldypBlpXpMqT
eh3990oCSRjTGyS/9JDfpHHQHqfQ4mfL+QSuX24h3REQ9mYHRuUln9P27wic6czdQ+3sRsOHvyCa
6zOCKcstHneUDVHo5zONYCgB+L8vTnEb91lc99tJvo4sakL2IZmaDrZPPn+eiS2BouG7JaYMk6oE
a2U8paT2NYO/1WTBHPFXQ6F8gVdiFhnEAVBp5iuuaJSa2hb1EeooNqyrTRfgqLWR3advlrFUYUmY
5lJAXBAxUcgTg5TWkXdxJGOq5WE1CfegqjWR20THXf2h4dXr+MJF4tHTRSY9G33nEGK3Le1GkUna
/P70Gzc6LsEyn7R7QNAp62yWhnTGUln1YmdBF4iPJe5gnhyTr/AyMDjZftYMUgKVVIWLYjp6jvx/
1EUMt42VxF/BDikztjXq0eIlayKU2M7PZBaV8jNt2B992TkyJv4uZczGj88vrN0RLbGOu+DWlZqF
CPC2h8qBsehTOM9G9BX/a6XJtqS8obwZgAqqKVZvaKKiEmISgPgVPLXRt7y+d2WO1RW3vZ6vSYbF
yBdkk4v42Z6XNjSMX/kddPm3RVHuype2H9rKaTPmlTFVUIsF6ub+GRoa3e/9rup2JOwNAciC+uV0
H23u9ieACQLJ69ZPRuJvOm1NxW6ulnZy9lZ9OTZDS/vPuivxSLG5+Ka03CcdtDT1KRPEKCU8eZoX
PgSVrlAyFFQ0zyLzETfB18lsTTBafOz2WQuGJhgBSX+f475r37EUOquryD3hbFd/R1pugm8YVhwt
cAZj82FXqOAQfLm2BfVIPbUpGj24Vv67yOSR83tTox2yDTIuqVF6Pj9K5YA7sd0ZpnbgxmwkJIAb
mu57k4bWIf4PoZ703yftyBEo55JHiW+bqVsUkwxNm4vqNVezOORqrWIepS0YuwZ3Z0qTEUyrcqO7
6tatsxz6PFWNWUOPpqEt6X22DquQ2cq7J7WRVw5KCbuZqTn6zcF//LxJ02+RL8U44udpKrWuP+wl
VJqZEEC3GBwS0BYaD8VNwL0P9TsSpiiL1U1SUAqjvFr6wifmrDprqzGix+4ipwOyJ45LkrJfHUl+
sgiQkyLBq5A5hvHOM2jfSH7NfMKpIKDmhGJiZgPfCCTcvMzHah5njDh/hj2gerYcsiTkkCXM6E75
TBezxBCDhjFyh6RUtrc9RLYU/9UrJzZbf8bgFNLVisUdLdELvfH6Hu7CCui4dk2Zo/HT6ZMkmEqi
IBw9l6ZK1YY60sXgKZyXCuGynpSd8d0wWGN5DFqyWd75L0jJ4Uq8rtqOmlyOhoJJrXkk65qSLkx8
wzPqDpA8VZeoj3zy2pdjqrBIcbjxa34hxJvxGBpAfWjxY865fbIbuClwJQCj/c6wzJqeLubmZ3+L
oGX8Hcu7hY/wi47rZl5cDYvEVK+hcB29q+LftbiT1/GCKbi7Zyo7UEk+C4A969x1zBqIrIJwa0mg
upwmKfcmT/l9dPj2giLJ1nWcZmVS2OiBdftIQ/4yS5X7qvGjCzulzaHFwoydCvTrkxna45I0BUoO
mc5f7WP+8gL5oohNw4zkNlpc9xoAMmgqc531GzelR0Z7TOe3wD+g8TD7rcD79Luvtja7fGHuCk8L
1NCozsYYJBbEl3jc+X+I/SBb/Kt973V+qnmHkWQi+zicwtv8UTS7+TxYeZS6YpXm8B87InroGH4c
y4OCHUyTSSOQQJPiA0m5jcOyIac8E8hMbi/ymV5A1hm1Qwqv0THu2i8ulUqYn5iI2ti/M+NXM/JZ
lF6V0UN3Nr0r2EmpnvYAQJZ72vIiYClVpF6weq6WLEJsOpVks78yiU6wpwp2Pvw1NnrSGPrWGnaV
kmrfDyJnFznwF0NTvraCex2sbgCNcYpu6I1lYR7hszUX40NGQG527NVhhuB/3wIXfAQyBx64TcPZ
+SuEd/5wF+R6ogkPWFr/RV0iCiRqX+XfuEYdplsKltPuKMkRPabMMHSdWK9+gy5oaEKPWPT619ss
wfCM/rYGr6W1m/fSlZOJlFCSHvTlSoX9QedHuKaXPP0UhhVEyo4+YTFuPzwyzhEFRqM61fsdh3/f
v7QZ1kC3L605aULiA+5MBW0fph6ec2Uz/69G6fW0S5Sdwy3917IKNGrG/48/4Vlhb4lsiiJJ6kR/
RKhqCzFuZLwR295mJba6E1X9QAB4lWds0pkc1ElGD88JlaybsSh4ATZYGC2sl2jqKkxVe3MYX6jX
uRA9ZTZMkh2RXJXx59eTW+lBrslmxgqnBXiglnHHhB0r5vhYYQnjuYpzE5STyFN+yBEzryWsBPUA
SvR74Xh12oAheb+FN7y+zp1uzaMhdUxQQ9Mx5tiwircSU4CjjD0KAi5U5Kiu76pDdjNxf/bcKRIx
7kiVZxcgsyOOIUYdBBihX4qCa3q2B9vLR80S8+5SenJVIf5mGastC8QC4qHWFE6HdLu4/bnwffK+
gRQjYxKEh/b+duVPW5dYlFbJVSGTw83U3EQIjvwYaaEGTf6u0VFEQ1uPKp2rxXa71cSEsXQPaKN6
rv1EQULbZ4AQH+w0j2w1wzMWLe3EdAg1ECUyIAvXSzgoxx8Yv6w/KwzfcOgWtrx3LIAWmcMCSpln
POM90ypeo5g5gqAWqgDb/hQBq+xfb+yYntvF40vRhZrGxa/lrsmEPXLDHpVlMavP6+kjqeSa18LO
OoxsTrsu/pfMvetGdzd7rrCCaEBFr1gLdS54vht5NA1L76U8YXV32GGeaR2kzCrPbRYdl/2LTQQu
3cMVpNMdyAs0nFxg2ndFL5HB7iMbQ8Xwet23xQxCrAFsMz4zYCsn7+dHXjJaacB8twzpDFOhmrAN
bl5t2waszkBcKxLXv78I3rWdVum4KAZj8/mck1FsuOW4lYivYb93ikvDy8ZCxKSbOvOR25aeOPLK
tF6nzHQCPw8MJX9z9w2xs88GwfOqje21oZ9/Xj8qhCdPaOkn2UghpywsLYwO25JSGUxRajna1dHX
Jnrpdn2EcgAzO3HLnYnqC7qOhTEbYf42ZJ00CjdMXi5+ownbBbJk9e/5Sij0ouYGOJxyEJgI39a5
sbTBXVQtnEGyAMAqqISLgKnV5BAB6vFioyTODN5locijmxPTgR4xxvhP3qSt9HzK4/MHLCmRQVNx
/l/u8aj6lxcVDWU51j4Q32txodtmG71Qg/8w7WqzFM+6X1kfiy4xE5793WmnX8llAwLDAlhKrft8
mjjuZgn3gIdSgW69W+UpHoQGzuik8ZkNo8meSR8odUB7K4Ta7MUHFbx5zj8DKSY9Ublimdmi1q76
talFu1PcgvJBFTVJtp5ZNmsOKBoWZziwGbrWD41M8oz4Z8VjEDyVAUMJAzeK93rFlRRMSb+adjPB
Pv2KuIfA6EyyFYVNAJ2sx1SReFhzZP8EvbGp+bV+tXcDfzdcfQ5jkJ5Trv6U0Bf1zu7mBNPVugBc
UKXJHgo6tPJYf8zNnQnHFPPCrWkkM5nK3VoSXEPyGFELPUuk11e4i5HkBV3b6rrYmFLeTRWaZTpZ
ZhnxqwlshUbG3q8qmjOs04FthZVeUj99MhTcTgqK0Aa3ggmDFFD8sipQhYZLP+cWj6Ap6V45VvYM
FSBNY6OCcomafnziXo9dna/TpZrEflACgqIQOV1ifoDDoGpwXwhIm+fC190xf5cniR0N7BXQJaWd
U+axqpMAgiEWvJugl/MfvSIHIsZPJR/BuA5omc/QwvyLKtQBibrg7dFiCGYYzPLjODNkpmO8W61n
vG6G8wGqCEXclB61myjcsP784VU3lxdmxwfyww2Vp4zbDxkwZvkpchbrn3ca7j1NucJgz74fgU9w
CdhvNzVxQEBY8pmENYY/kxql9/DDE6QHm9IJYOnTq6bOcVlmicp7Vcet4qMjwVhe1ki7Sd8DPr2K
sMBKCAYIEKcp9LcIFtZrAjYbI57eTzASBUYPxUvCv+A0z4zj8Tmhl44hnBRXlJV1wUu4AHuZeYgs
gN3Si2ISz3i3dCoVyi/XqrX1ipfOLbaLIKIBubdFJANB3LFuQr+42P2H5srTFPeAUe/v8pQpXyCX
6kHeOmWoc0/JM2SqvsWUZwZVdHHMrVzpOlkrNehc6acrVzUg7iJ4PjJAO3ThId/5cRXT8pmdojHx
3Zx9IA+EiG9X4ZHgZPArYbDR97bbM62xd79d0SILXXYGMzLhKwUBxrXrFHoJB8cGjbl3Gq+ae2aE
/n9geYcYE/2CK225VJVlQmaMl0E93lJUDgUg2mvFnll5jw6Tqw2KZz3sO6y+otSatBFwwcRJhjuB
VobrKdWdDKVhXGRGDEKH3/ff/IJSiCbOAmfS1ViWpJfiG6LbqLJLLgW5GJllG6XWcr2Ba16y/Foe
z0chGUqgy+N/zUcix8MyN58oNLgwumqUattaftBm4UUmEyW7hLmmLRomn6Omb7rMJXlCNvh1WmVz
bkLbw3c3DFAKh2b7USQnZXH6XaQDVcXST95nOMRfa2FF1JNXb61c7BVr4Aex0+OfopepyHxnYB3n
icVQs5cIscDH1mlvVd2IBvxuxpzGzyxYhCDUmSzaJvhuT9WA4hbkxQCsFas+bgPFw9jlhduQoubg
XOzW7mg7lnwHzFQPdfJgriix2CmCvALjgojPR4JbvPmSO3HpuPF/e/Rap+ACWBXlxsAnL+/7zeBk
o7V034qsZ5tOa5bbvFWlSIY84ElrhOV5ij+xdFWwXLs5dVXcaDGe594zND+si+Vde2XYX4xM7NFh
E4LpzZ8dCU7YaW/Jm0/gTMrIt51c38Y4KQtYSQcrsgooXpbbxdeGfQPlKs8KFKqXZFjzw3EIP8Ku
M085Yv1w3HnDRDF2JPEpepWbMELeKHUDKP7vI5lS8AhH3p7/snEJNfqRaavXX1Vn5OoK3L02Kf6t
slnXKDM6hIVY5/izofps6YSV1+6HBOnbv6x6g+0Z017zPc+oxpggzIh/EDNXSWzKhd+ScY0re99U
inJxTWu0KMM0MmgE8T0dUH6wKrPijcUhcuGSEYeOkIyKiUNP1MI2bgs/Be5m/1LDZPBGsbg/gdI1
pdda+gk3N7oz8rr9N2qt9+fAfXc5rFuC5Hgybnp3jHaNetaVwJCgaLGe7GXuNgVNxygmAXct8VnE
aSEVOR2nDkP13/NlimLTN0W+9J7jY7zxLF8VN0+OgiTRl1BCj5Nic/b7eISDNiYTSRcO0/LzBOmR
ZqViDPNeDBR928POAokqgX8lrhfLLMC19Hyobz49FjQOmiamqMRBek83T33wUMj8W4+HNnfEW5OW
EPLqKo3rJIi73JeL+bLetlwxiwE8KMMRuY0i2Smbxfp6OwzxWkVv8OUyO/01mnAQ19zSFxb9+Oj5
Z9SRPAeHExsjE3TfEYs8gM32Nqbuyf+8k0+luBo+d3+A1bDJBlbhhoDobtQwOxpdOmnO5DXr/U4o
cKYcFAi00uE1lL5+SyjSpF+J3D4KqDKH+vPHdopqlKnq0N51E0Ul2INW15RK8YTBfXuJ8tRS/QcD
YHoSSuNetQslmxNWeUyYvIZfSvHXNLrlA9DKGCupKSlalJmTfK3C6O74SCTnh03/9Oenil33ksFz
ROzgPSIUWVhTMdmCu8xY2OMSEjoy+pvKBTF8PiI+jU2BstGfzAHpNHVdRseVHAKCMlT077G81cc4
dYXJ4BXWv45v/QHaUcFeN5kJwIqNqaVt0Xbjpz4N8u2fGs11vweN4KCYP/+MLBp10pNZKkeUWNGT
nbrrpLBVnzT/YOocWcUbceXadTS6xSmY1ye99PuEvuoID2S672hVcSfhVHUhXTgWCQZkSKpHS9wz
BMX6DOL1571Aef8ItVMkG9KV2gDMDEu3ZasKwkZYw2MdKwHSphz8EDxRISUNg8gupl08vcktshfI
xmWLzl0KMBFXBc0tcVSF4hikg9CyxOiGytveKWFXKRf45IWyfLj4fpKX2+yTiykBXjTO5hLMN5+T
aOJqVYFRwjwZuRiwqrh/a7iH5aPD3jBNdjxZhH2Ss+uJt8zARjBgwCJG1pzhFD0azLipo0GZ4h+L
i9FB7mO4JJ/TL0Apfgpifqs1OXEaT9q4wIx8PEESgONXQRDJ19ddxZGeOZZjp03FkMbcbdoeoQcX
13U/zj6xlqUYJfsv9xlZ1LML/66/wx2eTu2ehGeANeJxpWync8WXoOJcePp9QuRNvyYY9U1mTTXd
b7ND0b9xr+AkPWLjUE8ll1b22sdJJXZM0jk0MZm81dpY25AYWlXGMx4jhLP/lkHjnFDNGCAgEhee
NyeBafJeg1FQYhFO+nU4x51XyX022NEphhcq+m0G/yao7aMlksz4dCkzTEQP6hnbuJFWOB4LNZsw
1M097YrplryYEnx6FRdsnps6+X7G5lBQU2s04byQKzzJ0I05E2evSAe6gQ8/Kp/OxLQMHG/T08az
jIAbJrufL7UIPxi+nkhvka/6fXkhQQuysg+KZ3mGq0NEs36squdZ5veNNEBwKNYpsPc9ec9sFPSd
R6s9fxzN2DMXvNSo9lACamu0jxxbfx6peziKfbQ7zAZh1T9vFnZ6AymL36xfdXbEGEBled7SoXsS
lDCpeC/+dZHkNIW3KUlhDNE42ubMXYK22B3lz5fU0qp2m4e8mnuhjV2I3arPYYgRIZjzrmf98Mz5
5Sg9eTAAJepm07VuNomfkPaWf+yxwJAUYuYXqgu7SyM0kjgQw2Pqs5QtAmk9x/vWVC9Vw/YNBzTZ
BQtKZIHnsfxhT3VUawOvZ72GZaH1p/kiT/0CNxX7GKd3nPGLDOuNCs6S3ipMCOVliETT2EL+ULFt
DSr+eAhvvESRDcehGZxRa2bKulq97vYK6Un7ic3EgKwuXNw7WwKzuPdWmRiJutaLZ8SCWJLXGKvw
qp522wTOlX4ZTAVk02e5fsnZomoH5XLRW6pjzbE8N8eR3gb6PfaIJjJ2t80Gsk6q/Qqvj++I+eF8
g3VErqvsym0XnfVa196KpdX1KB8hhY0EHz0rwO3ixAjNDzmzF0l+NLoFvKPDq5P3GEf3VO+R+WNA
y2YwzP6/20iR6Tjr/97J0ZHOTYDhkXLam7Zqw4wq3HImGosa20bioPHJPNX2aZVaTK3TbkRGosO8
MfUbUZZzT9EaPpd3lZpzThDLsqkOyq4/u7Qa04D3K0z6ZGoG3pbtxmH58KhVvk1H+aEJFYmz4IUV
UcpFatfeZUz/ScrM0cHgynQoHmpT6uH9ltmBcQZfA/svf9z1zgIk0H2ynu22tr+ScCn5sp1HkzCD
vfSaEA7aiJ0DgwW+J7ivEP/bFFiPWQ3LngxCh69tsorD6ndcvl91rCCVRkiUGhOAgFEmDBmKxtxT
Kkkoc7fqJmNIFAD13dXn7mOjLtnGQRxjy7BVDZeWw+vNizJXSlKe+OgCbogUcOIb4dKqdwBex1et
IrCQztZTWN1JVZajAvx6bWM9sEPMpq/1dNpmgjoSYLYM/WuZitoXFoypAej9iH65Nql+JQ5IL+n+
Rho+cYzub+iwQH7+t2ln8wpuRyLwzt0ubB2d2oPNrXhC7Q149Qazd+MX/WU9BYbCoCY89EbG9ruP
NW+FzDCvo/Q3+WhP45A6ErX/fLp6EmIrGZuQxTYSp3NhmIRBnYVx1rx1SZ72IQ1IZ03EkF0Gc7OB
sBw7eu6t6kk5c/sf0s5NCwpZ4yuA+wWabtmUFeCX7Ih/cHybwwNFlFa50bbpp93QIx5LbdpIJBZh
IygwroD4ehY+RA6RhwQp5w7dUr0DAw3TbOoqsLmYos7STwkJusqxk7GNrAxsWanhPnITgjskh44V
nXhzRJUsNACZE/BAYQPYvWXnweaHNJr4kERtNUWYHENqD8M07/wmig5hfuKYbS0EhOhIsL16oEc0
kugy68M8fYcfjCo0wLp4p4oZQwdhXVWS+4p9DR3/55IbtEacLMc98PSy3JVxu8oosaw7xBteUcVF
W9XYS3HK0mrp8aa2o8lZUG7u44W7qB/ZciBZV1C6Szx9o7g70m0p0b+vZRHjFJ0nzQLC1VUnpAa/
iIBMSwe++wB08NKXVUgQKo01RJZEvCK2vRZYkRsk4F7La7iwHZlufYH4wU+BD7LX0qM6vIPX+TsB
l3PRtEVzwXrvZAvqkks8QL9ronh6q/1ZCsIpP7GYUrv7J/YZUKqK6cc/iv26xRxkh1YPTrQkKqI2
GhEqD+Ka1bk2Kx131xueuImpeEaB00G27vk91n5MN8DtHGGNQsKhfAu6VCOrUuXGQe19GKd1Fsm6
YcC4HGRSZHp7aTtfGBNMucDY5JLpC8qxnLCM1qy4Ll6iznTMFuFw7uBgyQxU18c8sjomrs117oBf
z4ND+IitC5PKX78Lmsh9p0OM+lngbna+3rLWjMjuRrKUn0N/Rh6yA3f/TC1fUeWKfLVts7IU6LsC
+vOvut28k2uH73+O1jQ1KH2lI5xX7zCOIf5qno3zhhI+ClYVI71pCYW8PzbZ568h/fYGDh4kNgts
/shORiCHvkdt9jEskIg6kU2kOjSixft1kleO3SM2zawIr9GzL7IUfrHqQvyZBMPfpusCeIoYP67r
rshPFT2/barf68W/bEvPwf69SuB0J2WcRWV8Vl+pDgkfJTae1leuxa/UnxHXPk7PFpmg+fvjipqs
kz9o2rBkATIw4S2c08zgSgoLVE5S88ccEqtMdmIytFZZOibZJADb6wEExVYmjFq1jijutFS4qR7c
3RLeqFsEpdkuuWmqHc/E7HDFDMZ/v6jijJeZkKWOnvjb0HzQhYWGxq7f7vYi6r/ZTwyb51f60ckD
KcOOoG4Jod4JTsyK22q9hyAO3Bk7WQ6C+c68Pa3m2K7jWfDdBUxj3lg3RzyQ3DxWXx5NSrWAUMqf
0yMUIkNkgXc/8wMwxZqlENZ6LCNNlHtoFCH5unQ6mWQ5RvABMXXp6/2OvXtWtoxekFjUG2jZ+U7N
faH3sbeRa/jh1Wn2fTqhfevd52B2SqXIzBDaRkjBH1sx9wh1ltxL9FQHLNdP/+ZYMUxVei4zg+Yz
1aKRBvD0gDomY3Yibnp7n4ESlrB2T+9qsRm9lQyvG+btJmMHfYEqU9UCOx4CEMw2bFvPAwN3ay5P
4HJHUIORYzeePF7eHsbatutab2XFTXydMmxUjdrPNNi+2u+JZEqgWG6mLY4xC/djfcU8Fw55Rp3z
7E/5o5KcKf0ocMLdA2C0m7d6jzaWhcwd75nVG+ad830zb5Othrjc9b0DnPP5ziyBh3WkuSQJr8td
8dGAcxKSrGTJpONauMHILNhnoCaQLCh0a7Tx7N17jHUqdFUgYkV/tPi8IaYm1Zi8DNxf1oIKv6I+
J9vxJrFyhokej7tFUrPUsLeOs4FVnu2O3iO+odfpuIPCsIiZeB4bqFVl1XCA0RGkyOqOqBkpX1sC
ZF/MlQgFcU27AzY8S3KiC1SRNKgNum7Lyfw1zWhM0nge05/RIqSF6ywqKOT6AvQMS222UkB8y128
MIs6MtN26BWziixf42vqzx4cFPgsfndCesMUdz++6jEVbPHhqLwt2Fk1oXt0jsf7m2gcgXUw8bjv
E9NIKSBeDZOyiva+aUaPaTWdk4KlJ0vhsslowuo3LXwE9jeVJgTG4pZ8r9gN2SCbuRmzVEsm3Jyr
nYhbp1ZWJ3nde2lM7P45kbXfZEstQDgGA2oFGlV4pzubjDgrkMyQ4nUV6S7olt4MRYYtzWN4CWYr
clslcZqtX4tbCofiW2uaLFEOJg3NHtlMgZoBNLNf6BRlR0X7ZJZn+AyUwgkVNKSAZQztWz05M2d5
vgM0SwpoUZ2Sjd6SxEYiyJmVRZlpdjZPybF8cx3V1ZAufpz4MjOmsCWDTkRuOLgivcDStWOZBxjp
7RAM8ZpaMfjIFGTfjND3Vi1YRd8gmeQr4hI1be9uK83xLQ4FaIbIDaYDFj521xULK76uccVJKafP
7ZaxD7hqtQispckwpWlVvWIS/yd1kwrA+TwzRRUWnhXFC1CZQ5HUxUAFRk9jXQYPeEg40NI6NRDb
dwyQxKqa0SI6SY1xQlgsOgI9B/ESieKWec8HsyxG4bmjRqpEjRBujPjD2/1OxrhjT4oicCro0cjr
UsXfAAYiFL1pO8l0aZy2lPxh6UtR5IJA1p1kS5ko2WizJdyrlCt/s1FvHw+gsiuYgg5s+ZwFlpbG
WSedOetuPYj+WcMsluh92pYUrf186f18xoYS4bgaAlyYPF1zcPcPEHJdo+VQNXTBbrg+mSh64Q3Q
8P0caVVbv/IXrw+yiQZQ94QY3ltEYFPRNktQGj0d2kCX4CgvR0dNfQAso37oRXKirMo70dfnGbQ2
N6yRajzo9tX7bktBn0Jkf9RA2g7WLCW5k5qY+DLtDw4Bbel9cjAW1fHENZQPbD5hFKPet0EVqhdq
KNrK6O4EQQaVoTrZFROmQRObDVXU5a4eUW3MLiUTn1tqQL7NzVR4YynObkKZ30gcBQ4aWbyb2kxV
6R2T2b3THH0IlI26Wi1kXz7GfdU+uUQhXpTPDxzLuVZ2vYBo6tfKj97sbQ17RHQ3aLPoEeTjk8S2
nXiObxdzHQyfnjqJ5Ecx0kWo2+9fM2bQ8lLYqg+nOqbpjvGzHdA/69irTmDGUrP+3poq+sP9ag3a
nOmjGtDi105+8tEZYB0vYVLnTHV9XRMirVv+vr+U0l9Rkm2CB7cTE7ngG7EADr4Z8w/3ZoWfYjSt
TQl9a7eAzWUTpf3RAhwfv4fUoBdytMeSIzkUxme48pofHRij7pycKts8JMHy7lYp9k06BvsiFC/8
7pmh9Lc8rDl+pNI/y4fJnTZR+XmNALDvvaDp5A5pv12yGzaJwVAkpfhuo3W0WEpmCRQlZ5gp4WLy
1ZNWQidCKryhCdGPlFCpXaq+07LMNOdxTskxG0Dw6zhc0LcrYfRqNA8B2hWztUETS0dZdNeYALeC
UU60cDgdCOUFvTllTjiSEiwF4eIBxv6Np8a9DWSDZPQs8U1ErEgCMtuR2o8iPgq1lzmCFNSpXpit
v+HxcTfFrMs9UL55Hb3viT6teFDgyCknhdYCumTZhpsl6WU6Ho4mX/bhDoHrydW/2Xp0JBa6REP+
/34/faFNHhmzOWjg3Wor3OgQzyiH4Yn2jWQhm2Ern2i/KGjRoPRvVe9iMUY/jXG9tKvRl5pOPRiq
lWgo4NsebOgqUsGDNMavuf8uJvMZGQe8YaEEEEn4YkTVMxO0fWdiS61I9OETYDK/uTHK2nsgIUOJ
4C7giH0e9w3krXx+1d0O52uwXfvRhTCs1DmLBLE59yMqyA4PvvrDJ5YJjhsFkm7Bdj9hu01juFta
gCsm2Z5g8Fb4+OTJZBmdopj2uh4hu9nb5XOldxQ5MkWfz01H7TYfn9xj9Ta/UAYEGNyS+fgMv5QH
94TrzBr5tJaRt23kmRsKeirgGSuJk+YL9YUs/npqw0dbGpCoi3He5+aKqwcXiy1DhGYXSr+dtWJ1
k6UxzuzKGkMVVqH1/p0pDyYFvWe17RqKft6BtF56NBNgYkOhnKtrDtxQMX8eVkwJIV9JgbLyxnit
h9cwIX3vstF+46XoNHFPxTgaOUOVH0D3CidP5SIvmGvbU668NON2hxSOWcxKI4kqFo7CLy7UIJCz
pdwa4GlmX/fYxVlySWoWo0LFr2GkLZAogZu9oAj+nzHeM5uIxmsZYKwqgM00A8L68sFfDvpYiRhm
3LiupE/aNujH3n91FUNw4YZr3TfKnhsEsw+zKMoK3Zi8FefGavRRVhGv32g0OwiRHclLSCfyr0pM
V0ZB4Np1hzlxcM7XIev/AgbL32BcvP83hILMIILYV7RGBtkIUYbgTS3fjEQlGZoQVuoFjQfN2kGo
ifKjiFtU2FyOxUP5hYY90+IdIiD0A65H2G899yeFdEU5Vo1Sk8aNOlr0ymtP2zfjXLmi9qfLPWVw
FGcGyMWb+3cd86hBWr2RIYKgm9gK72hTeDqt4xydo7yoW+Ck/TN5693inwZ4olQYg27+B5QM9/wV
7+csds5UAkdehrdF3LKlX1fa5+fygRJvnGrQmxa+hH017KYQhkIYn36yKErVrRNcr0mnMNKGuLDl
YYrqTW+zeoOf/iL9yCCgg2iYebhATzLKiSz25F/1mHuZZOuyD4OgfZBV7gU9feOIZt+i4C7uD9tV
9Pwplmhoqp3ODlYKZh2A7fQMlJnEeXL8fB1mhZk7Aqzh+mVbjGy5W/+LVFDpP8Ka4NfQssRNikuB
mg/uy27OfL/MmLwJq6V5yCEr3rt/Dnva5HD3CbZqTFqv69KL0ilxTnWwfaisGwekZfmuAFeDRlf5
iSB2QNe63z298qvpv94VxT+65MFq4r3g9/DeQVY4SIe7BMjP+klHB4ZtKwetGl3Ahs2/XFqK2hEm
mS8epMq6SFn/QYD3DEnKlYKuCLKtDfpFsGFBMSVGJLqtzQIXrKdqFL3UQoCLW/sODPiWSGGdJ0J1
5DsgBU31HGQ4eE9pGLob4A498pQTfUMKBu5uTTubC5TE1zV1Qbnq3LVMNC8Xdtz2DiEbG2HVOuZR
0c+/Yp1hGA8tC8TraDZkeOGV/PL13fMnraUmAoB3sv3pYPqIXiquyf5mFmWXRWs47Xhe7ZIkJnQs
DyrWBRDREGPli+6I2nXisfpYsD5bW1B3dC0PBxWsL/xamX4gtH+zZzTO3yi+FeDsk3W96zVVk4eD
JTMmdjOUSh5ABQc7aAoFPuHFNQrg0OUfAmGA/Lp5fJJHnDfrX8Iy+YBbuf70SmfCwRZrYkMGu4IO
gLqRiyIKIGo+ePbMLflpSxIb9OA1OD3p/ymFVfTc2d9ib6xHF492KJ/xDUpPNrqNq+G22Dwt98qo
jMKah/eUia7oeuOklg9ZDMMljvPXU1KZa9luf4I1dL/X23ADKrLVw3+BbiDdmXWCEcMj1csTEL9L
tLSmHPpXxiukNUiwBijgbahOjXcFbfcNow+IUBZ8gwxO6cxAYg93IQaN/2l0jMFBbMkDw8oc+AKp
Y4T7e612WW4nmkoOHvv398Pboyzai+XpWv1fudGBZtdStFO2zIucu6MJ1lo5DilJcZvlyzjMAQWc
5DBRxZAG/gEo1uRs7mIhy6bBgAsWh1Bic4p0a8u56CAbBJaZhPj+EoSkYQswAkti0OWgriWV09AD
2leT8KecPDZrmezbgYpRzrPa1eYn3bvE0COyCIoHDvKQJcLJb7K4bv7bTCNzhFzidWlsxvd8hNZq
yMZwqc24gwdbCriA8QOOj7H+nxGahPUcYyxv0VInZ1/pacPrUhX5QLMbi0/mhsOyii9hoT+sD5yA
kYgits+5Kr6YP2o3vtx2oovuKHwEjxYIlJwqz/xcfJDd5Mj8v4r+58fVoa9hqhHFv8z3QjuUxqvb
hgvoacYv8D0Y2WctAeSNW5eExADlfDI+55d4D7xx9cQn+Q8qyeF2alS4+d1FrD6kFYlPchC7bvuZ
+5+LTDQAr96pJwJ9L3aofVET/TTWa582+Mn+VrvSbzrcEE6MxQYDbshCaOWca6eDpbtsS8b6jnzY
vVbOF4hqt4jqQ5fF3xInjR6BbUz8oMzdzyuI1/iNjTJtx32UrKulbmfgAC6jf4OBJ5pl446oXpwx
IYC3/EgGpT4Egg4+4itvp3i+pMEdRf4GgcboJxQcreuYBf0nTSzjl5+yHLAxoQLDrZXMTIaEUexG
8gyQG/JDfkGKOfFYMpfY/G25FGZnePADJysYDCy82s3aR77b6r5gWDkfSMv9iw+BHMgrFb9lxdxe
9aQJxTmClkr0FE6v+LQYz4uIPlKyUiWGrDuJaFDsdEFf79+4SGWQ2dID+wGf4e4kpIhTfMlieWU6
BusWgLLDIYMw5r/i3paOohBsK6HMLPsCoGd3k2pyYSGcyewvwYmRq3Piy0wh4NTny6T/iulOcukb
3EVSMQVN/rFciKFXyJqvNGCS+sXpJkYhqvh0iAefLArqTY98gfvRQfgiUlp4P2McZDlaNPa71wWo
JEsf74luQ/yyn2sVIiqx9NCm++6lGA+hy89GF2BlQP0JkiLSYUe4taGgW9w7R8iY/snxUrB2cBrh
RU6MbTQFG297R79DrfgnJ0/Md6FdFLd5SxP9C45Z8WCeYI3K2XEJNk46vH3Rvmyd5NiaE67ef0HB
n8M6xleQo4gi6Wjpfr4HkLrh0TH2yt+6mP9Dit+M2wiFxsh08qC3mvHVfysCRiKz6MSQ6BLWDWdS
onxKqEV+uW4VeuvOhKIEgXyXxq6dntuYW3C+xY8pPUxdEx3ZPT0Qgm7pt1wBBzS9lraM3auPUDIH
cm3bY7NejitnCZqrpk5VYhoDza7L5Ei83lQsOzb7nyzh6Y7VzY2MnZICwKHf4yrH/pYkrvwYDc++
mYTKJe4NQXEo2YqOjs36oSVWWEsekMDnHB8uzBFGUV9S5XfN9/BAlkHjwBIoYlFUBpG/kCTGpPlH
Qubxvw9UXCuIy0cvqAiqOviEowaLnSkYMEG/wltHmmxVlqmCZH37Mg7y1TDwj23TXyiRy7uDMBmr
l6wUS/mXxqlbRU/qj0Bk6++wE9S58lhX0vB8NAM+YphLSAT2wR9pgoTGLx0H2wt39BpsP2KniiG4
WPKF6thHn1oNgjftWQBYF0A+JkZ5+0BO0lK9jyjoA0S9qxXc52I2kwPyL6EozhInDPbJ4VlzMGUZ
GrO9ypitLnXzqeAAXSr63cK7KmyQ+uhhReKD1uETGJEwmFbL+bIuToLbi8n1sv5NfWc3CFzbZsEr
SKTLdgWbtKyBIQx30h/HvptmvoEZGri65tziQi+KNZHegEucVrrN8dhD+D2Vq1nt7noupwmR23ee
EaEf2qNmKwOo3GezbWTWSFn+APVAoBy+IuPVTzQ7zyIwSgY+Q3rglilPXTDZoPYROpVXEiuSII9s
nMGQC4b0z4WmXWdt1DMuveufpDB49f7prEz6lC38aVGvAGKACHv53ALo9MOfyy116ml/aSQGJ1du
+6EdxdeFWeFmbK93kKcqRhA2DKFjohcHBin8KUwcp/sLO77aQB3q7Fi1Rw8TJqP67tUyanMkynff
ZFgkjQKdq9PHa1w93E+hySl5cm7ATiyQDQXUVvWqF7MpjKw5qjiUY2PfmDfCavXKCnxAzVspHM6t
tTf6O8O/kHrkvgjP2YBIfn4dOFgNKRhE0Hy3KJZP9HcG2/n6JgL0WulT5hYioqOxG066Qr65bIAp
OsmwZ2CC/GY6Z2FxnzmZ+4vwXhWOsGPkEqZEFBENi35fOrQl01VxwnK+EYZ2lOI0lxTcbEbSn+x6
sO13Z5j2hHDsheul7iNmgc94eGv50EGxpQ8W3oGo2pDqMu76Ov0xaNdEQKWCfooqrNdf1hQFInw2
UY1gtOxVHcOe+npJ4ZcYQbVDBg11sUTYgDP1cyan8B+Bewq0kjmngXVVP8v19EcE6KkjR4GtPL1w
dD3Re2FMRdTeKYKv/8IFLGBfjIvchSp2dqdvTL2VcBOfuB+Zy4us+jRTSxi5lT1o2aG0+nKbj0QG
yqcGUDHQclrjK+vMXF/uCU3+MghULsxUw4wKqiigzQscYko6/IvK0zbm2mgh4GUKQ29CWKuEOoPJ
7ELQM5ndIHJWKExnDUgHlb0GIdJZA+JUAOpedfT+eqjEgWgMcPZee3dbMnUbMU360e201znfzpHG
mQfLBk5q0NV1tqNbRigEVDBptr234gxBhNiXf+/SvDW2I5MvrtVgHnsF5lkwdUI8eFR3Niu94YG/
54Mda3OzoXeAJ3r8vhufl8aax36jUf8w2XOOPFG8rN+4tw7t517xn5x0i9htcaJygQ4cqoppE1Ak
IOTFowBKEmX82S5rivJKGEv0pE7tUyvnp+IUX6jWXoA9BKQRBv/++2jJ2rBDyjQ2H6iBEAZjWEfr
c1k/2SLnQ2IWi1q2C6mNdqIm+8xrx/wPGU2nWibiisfzagyBEEKxLj2yyg6nhh30EyTffRXT11fS
ivbuimxJWJ89bqjbIA8obV4bAJ2Hh+WCR0N5Y92wd30DZKerPcJsNaaLLOieQypOykupLRIIpsiR
O68N+OaSWgo1outcfKXE/o+O1yaY3b9nvQiokqqhw4ruMVOsJr8qwbOOgBn9Y9scVhdwVibyRgkR
SsDnsgrNSdTpbYZqBqFWilNS+qCkAUIfOFTqUw+vKdgvdfshnCGUWOt0KQc0OQYycbBPXa2z+fx9
DgfVlpy7LTMKtiwkIfVo63gxHU2slhVEp8k7teKpa06hG58cpAXAFYBDU9zn3cxZ+dTHJ2BMbZoT
zVFbqank7FLNg8eBTUVcpn5S/Ej5hLCs/w9uyriHlLSVHm/iyC6Lybz+3PrSMAU4QyjukXi59nlu
PgIjW73LGRNFk8TTctkTord56q0ET8dKbGJ4XnGghlQV8E45IrKaRz2p8lkioUnX0HSrHyTv6m/T
Ty4Y4Yf++p5qdXqMNYcIy+CbSvKMb7tl7TvFuwKjoO+iLsBumJEfOX91Sj40kd2ZwZb9GhpOnhQZ
XutXo4BPmmu+s3mwdsM4T11l3JxBxDdbfUvo5owmCW7sS0i0YRGxfrDL95Rnhz68kxE+3WJDngKQ
nJ1tXea3zSWWukbncyxIGbylngiJwUjn40oufyJs1I5y6A57RFSxSTAdPNmRACsGItf1p7tIPeky
HA6veV+7r9kVuur8LXt+QHnmvF9ocqdoaIm84C/4XV9tl+E3OSf7NQhhR0ZYdIiwTrvyyw4LwFdQ
+B1xvXdP6D030I6JQ6UgFmB5AOkUtaa8/PNDb6J7vEdbtwDTU3AnJjTOcR2OUdiS0FCUyHyiV92g
4S7YuTxq0eFcGOi2nj2CRmJxoEyZ2ARCvxxRk3CycctRIBcG9uYa1wXsxMEEUIz6ihXHAA02i4Fr
OQNsDntWC6W5RiTVGDvo6v0ogVRmqsY2krXIau51PDhcKGaGpEa/2TBQ3a0zj47xbHdAVKMNrKgC
lg7q1G1l6XLdQZEe+fzDHNFpCL3hjOS/vbB9gjEOmsqrz6gvDH7qztkwcOwDDGne6s961idjoY7b
S9ayIa7U47xzUskENxh4hNGwY9/zuKuKoAPOEfeD6/GpNKdKm0Y7CyYAbQYm0tu5fDH/Qi5kstJ/
LDaGB6YCXEKRIlfXZf902SY3U/C6RK07Mxs16yysqbZyG/9NjFpu6/MaPGWSbRR9NHrezLTxJJsz
oxkm0sN3kW9kRUUqYeqzBzrsXuo7EnHAxDTnKepZel+YguNqPtBaiaAdSj9eA1roeT2Nqx7bVVdd
Q8FtTlZHk0E4NcK4I557e0BDKWzjUCiawhEdUcjj7GwqsfiQzcMm6T3QuNStXl+u2nk6mEqWfbDR
r4FbpT+e2N9oYH2pFt2EFplgSwB9kgs2zoaZ7U72j3VRBv4tQw87e4pi+PsI0rPa3oCR8Ay1FjUT
V2t24HDXHkUCvgxFXq/kfaYvqzz9VClhQxWTD/ibo78F9M+tBrRmqBOf+XctaLy7JJ/rgS8Fy59Y
Ua6r4eHCa1uZt3yG84GvTNyLmzcWI5bTdxCdY7nRZ4q4z2xYWdNyVTvsQNDPGSbH1IB3CNHOrnR6
r0vOZgYF7Mt1aLaoAoNUAsYgIxryrBfapuZQjdU6dronugASwWD6L7yF5ARSt5Lvoptof6p4pi5D
4e0H4c/8xpQ7xmKZPzB7kzb/vRgAtyc+FKAyOcZ/P0ARP8lCQW/Dd1zDGIZajSi+IGq6TAhT0+4G
FbWANCsJnTm7FGTjvQ4o9SBsB1z2/P8PQ8uDVfHbcosSFdNUlfQjz6WmxMDRZ84wkK51wAf4xv14
8428vSf7vu9V6UyFy7uWwKNT64geTe3fZdiRfJpaGApDZ4qNOb89+EfDV+zwME7GpoKYjL/cbwcq
XcaXXW74cD8Jx532HUas660qMNr37eyYS/UflfzOh0OOZ9iAIbJZsNENPPg7ZhFv3tfJXam593O9
DiKPdI6nL9rXOl1TQ8dUuUTdhYymZ4b1hwkX8jnlpiEyf9HHEgU7XPULn5rjgWBIMGC6uT+MuHAZ
REpGSsgnuZOunlmySE3NBUXWEitU/r1Kc62u+gGyxyLwZ4/5v4ZOEPzrrqdYwMOP7QyK4MrKa6dD
0EE7NcxioaHA3+WDI/GNcBzHrsjeWGOvW+EKqhwNNRFjR8Spe7jpiakVowyB/jGpKPk5egCphAgr
u6NHzIwnRMNH1NgTFGu9JxDvnhSngYa4NYpIzSaKj6Q0jhsbnU0MD0wOw2ZCQwk+boKAMoccu/nz
E/uIEVwuNVrBFH74qPmWo9/+pCdKVJ4REYAp2m+QVljB5HbvSRwJmSDi4iDiX+BVMhDoBS1JsrBk
5LOB9TKyXuId6pS2dNCE8TT+JhjCyIsVit06BZmWWoYm3qn35dRHrH/vDqq34Meatb2ZqYQ9c8UE
37UmS3Z5nAqPp+Vo13GLPExVS6W68AV0sDkvVnrnEcDVrnwOba4aPemzCHQPltMpVZ7HjPX3aKKq
L0Jur1wj/LNPB71TJGZI6yBkDJYaQfr+QRt83I60vIFu9t6OOFrA97mZUxaPHAJAZrBVGEIeqJop
ZP1RzE43IrhIOOF1jFGJwboEquq9m5mq1MIXyhICGvMStQ3VFGXCkRNs/nlamhlsj06g0JwYqN0p
D+E2DJLYVQDOG69L6gicwxEGlHLw1jK79W+VbV88D74082A871YnYi007sU1qGIzE5yub8lBmOn3
nSj6C6eLKbT71IJW+HnB6bgcIXWqTknS01qXMaX3C66/MXeUiqjbG9BEys5KFCahLdTpBqVHw/28
UfeOt+D3lpH9v/s13ltJXkKUyFkRmZRUKNZnLwUBNWwQGcF9nCVP0+/L97mem2zEestgN+cQtuKX
17KyaG2H4fkOOL0Hw5sRuiFNi5PVClbd1oixMNQDbJuDi1JXcs42FAgQxuPGI/S9prOYIUzqUMbZ
j6mRNqDSoi9yAs+47QDCPVpewk092pBJcq6BWMnFRW/I6B5RpsvSd/TRJWN1zOb7bH9zO/JNejO6
ASzlwm5dNfpP97JONLGruOF6RVp6lRFh8o2J2F2rnE2F2PYW+bbEFZMkwZoIZbEZjGVUWSX1fwvq
+XLGHGxQdsP8FMDynz9+bhtbAJvo/p6qlIPILGQGmYyu3A0xb/w7wedcRXqOld/G0f4Q0SvEzIJq
LQnDD34MLZuOqd3xfqoLjZSJ3+L/gm6YN6n0+7E5B3B82krOlWkLzJs1vA9rseFvy3rfnIDemAT3
xkvIkj3XzP1jYZ3l4nw4q1skgC+UYwRTflLwCogrWGH96kDcBMHKF9qZxsB9wOuXZx2YpWj/eWad
lfH5gI7PhPwwEFt9JdcJW1MmghqkbCz9ePtvAzbf1jVqlBcSWYDoTSRTJGObaR8+IDgAqcITPsQ2
+T5s7hBkMiHD0oF1NYCH7j3oztozcgS6NauteG1XFUotcxhMqPoPBNSREK9F82hu9K4/CSRJxOSm
b9qXvzMN6IKN8Dx2rlxH05a9yD2ich++s3thk/FYTrerr9/GwVyUR5FW5LO9QGHhvQ4WrZvvQI65
pLsaxfVD+4Btjru2WMV5QN1+6VE8GpX8YO+XErt+B6r5HGXA7Y6lLy3WosvzbaL8Y4F+0rRyV+9a
7RM8KwVdOPCrR5nSefOzDiGtLPt/jNKPvC+xQ4vgDmcbnLYgPoQfqY/Me0nh8ZYp/0SJSz5WMxWz
ePBbYOmwEEjVhUtLKsa4r3CNNXXQSu5ZdhnfmQDDxi99Ygk/NECdhfQse9jkvR2pq06yDAQMysOV
KYGkqV7wvxvDHX8a2HjSPKEvQDUPZp5V6kcJUzuBWdxjCcbF4d86CUFpyTtzSM9sZrz7enPjKWIP
qvhseSx6K97p8vlXLTPxMvSGmp/p4gZCi9IdOSgblGHpKJR899It+Ct7AGIwc7x7cta1OZO1S52g
6D0whkEXnOfB7QNwm15JefyV9sFEmFW4iragJdP7+W3yIMal5ktyUsMSuGjvnmqWDiisk1bAuVSH
3232GBJUjxHn3R5rR6B3JCJ9lx7ORuNtugpNb7Qj8VmHP9sCxhIsUOrpSNk9nvm41wGF4f/p8vwO
/q9ZBbFEMMk8QPRz5Kr3T7ClYBO0pdav2GTbvN42DCKXHcm92hfCHeJX3B7PjFKXiCnv/NK1kDQu
hOtvON5p3/1wI7b38CMCHlJzrcGyMlh1QgUH0QMY6iMWoUM883nHm6JnD7HeA1VVUwhSdi0S6tqz
mCnd7MYNjSfILOPFJlew8pwnlU92VxJY/aWqfCqVm9B3ev6nFR7z69ktKMQyHNXrUmRCrOPp/1cf
dsvN0Ln/Y8Lz5rvL3j1VqvqYci0K5syu4GDdNO+U2r3tWTf4vZzw+PVnY+td81JFPLwwuf6cTgXm
mDHgBpGc6dEttl12bzwZDQWw8lV2xt8CNXUxOdh2nYGEF4ZUDVWOGgmnTqMg7PaaUikkcrGjWVKa
UO0pYsMzGRByc2oMvm8yliMQN8SnKhyVu2ysUUa440iuknMADQT3BdQYguGfPNvrcFCZJg7NSfL8
dHh03+ZxbQYAreQPDGKVi0py9e8lOruqjRDM5bNk+Qlj9CQVAQ3tSZHm/AcX0xlwnw6bFMqXnHFp
0RzQyi7suE6/rs/w+K6+17l0MUS35GpkyeRjsH7trl6J4kBSMIIqitBozOZNu9gnMRZ14vpwlZul
NmcE+te8HM94TrqFX4J3gdjxfJzrCkLmxjbJdQyPpWKJ49y+mJZds4oXTscBuisp3JZEfx4/K7a0
wJoSp6DBmRrqycr6c7jG7+8VUujCb9anJ9Lk2tnc8ati8JwVGLJEW6l5vB2iUb1rKmn95TpBdO+I
FHy/OzbFP2v7SB+HW30SMpV9v95DNtRiOSmreUP0u79oGAEEXegWshfltDm19W6F9cyC0N/5ihXZ
uAYFutbSlSOrMFnD/D8u+TtuDEPu6zKyP8qH7hKKVmKeb1gQipjHWLQai4Q3ipIVnyQ4cf11H+Bk
j0GxpAVAjyDTDerPAZ0bCM8swXpRyPLr8ZAIp2gum0pgDFXLm1EGe3InFh+VIfKNNQxzRTizBtmg
tF5oZjAhWiMpVcvAwme0JUD0tFA0WO8FssLfqJ3YW63A5uV/ISCGzx3itUAn+mZ9PzFj4db9a2gH
wwLzsZmYN3keJw8+JN9b5uy+4HXmaL8penOCeSf72CAM+Zxx9yDDfzJmsxjAiHRcFR0ah/6f+aps
VuiZPTAbk+XOu2csRvlbUP5gM71voq91cDdyG72KduCjBMHtXauakWFuQr6e5L/8gz7hcPGExd6i
NY/GtQg2K0Dut196Ev3Hz+UfV0sLZBOBAzYX/Xl+I3qLIWMEHmC3PzG+rh0LJ0A8dlBMb+9P9ozC
NDswmlzrw3fep198zzeAUNXQ6t1brfF7TVOeOB4mbb10Vkoik5SeacBQk2ECZRzaPBDCq/+XkG4V
cVsGIbXQk0x1pH6uPnf3ohY6Az3UjZ9/H24J6aFab/jlUVJYryCqv3ka0anetsY9+5Ycj3SEtvxS
/8HFfmjLOA4VEiO1MhMbJ73iOOHSX7POlY9rJO/DvEhqdUasvgoBBbx0g0nBgO0V/kzdUk+G9rxa
5Jyq0PfC+vcqao1IFZ/dqacvg1IowyRMJLnBmP8XbZuAH5H4iJERcIaOZQkT4aVmmsWEcY74mKX+
psT0XXIwPppri4HQ22IWZEw3IN9qluWQacTDYztpNpYItEGM/KhHPHZRXw2HoJ8cZgqODIOm7NFq
10v6b8af2/pZet/zIzbir+BEVnlFI/DEWo68PMEAhycIJxAtGGhAyUWwhSmVoirtSTAxuUmNTom2
C4GKKvLAG54acXcNFJ6k4nGBUNuGtryt8Oc1U+nVZcG0HZlhwBOQuUZbNM+sT7HGoQLoiJ2OUn0h
BMDNaPfdXKj+d1Mj0EM7gS6N0qgx0FE4ObBDjvQr9Le4te8y/FrfjAaJHxqOWTOe36pKNNGCUD4a
wLZnMqSCxyCQPrXvQwERH7vUpU30iwDc8D0vTmZMBt2JqkSezeFlRhXpJLCtzVs1WSo2asRb4iXl
mstRxXyCFoF+QLaYioBSCuC/WBicnL0+dexu1wPurnCA6/KbM+tiXXNQr+xCbg3CnEc8LYxN+ext
oc24UNmSYibxns/CgJkeFjrD3NXOu7t1HKdh11GDVXiiolwlcrsS4kahSLMoIhViFBACqsr8g4uk
rv7seu6/noKaxOpUcJUXFIuLDMILWbW4yxy/jY2G9UM39m+V5LVBD2AgJrzOV1x+yVsQZF9IrLQu
gOd8YJNQEMtUFN0FFK2fxMB2UqKZP/TXxgQa1D7po/CLB07VAUGqAPDclHhIlqK4b0y+CPpzdI/j
3Fzr5T5qJzIOPFHiVkUafeEURiuS9+11uEMm+q+rnZWdxq9aolq0bNnqgpUZuuIOU31MLv9jw8M0
hhMz6Dr3ll41Icz75lgeAgQOiwJJkc2Qo0d85rcJtq7W8bqXQ68ee4YeiB3ghHj+cgDuRpgrTbqk
XpXA9iMIH4cfanDCDjjUnxDvOSF3PV+4ktDSlmc1jSNcBO1raSr6rcWgKXTYfLGcnHESuX8K8fxK
z8DXYv7ED1FQQm+zg509pecsgr/r5lGlC1gPyT+d4nT+dLka5oPvS7QMZSLrGU8e1OhG+9Rxg3He
xFQw21/d6j/dYAb7KLi5TgNR31eDHa5lPJjjZ6XD7cDKjls4EZcaxng70KVOmoR9v46N64HhFkn4
r9lRVhU+v2Nsj5BBdBmq4xg9TpsSsqJ/xfs2JiImrT4QP+pSIO8PdDY1cn7Fx8BKb9b4ihf9whKu
YiCG6/y8NhPQkzvG7Mqe85YBE/ClUF8CYZfD6+7Vu6i/AJEj7lTMsgAAhpC1OmXnGuz0FH6Z1kPj
9m3794InvrBpFcbY8wsY/Ho+Z9zFE+UTf8Z/r42OZxHBLVJAkwzpQ6G/z/NxfJb9y55zgm2Cs23l
pzB/sMAA9s2O+04UMQPnm+FAP+yeyJ2kognS01e3u7voCEQnicU6QdMpNw5zIZVC2Ov6oDqKvkBp
ak6hC6eTHIoPmvgzC1Bkb0riE5Eu4GO86+09qscjM+ZZ46TGbdkNbDagaeDdHAv8julwuez7s9tC
Y1joW5AjO72pw0AcyT0ZaXFIkXtNqVn90OO/QcVE/fcv28c1+8OxDtBkso2L0iZ0jaVY9j69Oox3
ELunU5Z02UvJIXAW7GbWf1yHXeX/cHmFWYuV3VXzw/kSt9kCp012t5Z4rQmPTHrUwkSpMFmUYU2l
yCGYDx7+EaVg/ItQXc5dB6RdxRsQZ/wfSEoNTpC5UEdgSOfL6usDKBqz7yYBU/KctlYrEccMF9Hl
/aq21Tpnu+ZCMIB/6qKOSsSwvXGIhQgbAVoKD74s7LGZuGuQTcb22EvJLKanleVH52sZeNlikpg4
T1UqVDutgC+tvOCr7jkv99UGJaehwsOlgaPny7xWH4anT5CIcKalpNpgGOtUYBnKL6WGB91/DTb8
koqGnjqSoqSIOlk/3umGda7HygsHXLD+Jea6tRv7XLdeX9V0088vGCwoYcRVhuzF2n4KlbMXX63S
jBQ/zGTXmwSgNoyYTaaDFtAKGO0KsnhjpsxDDrEsByIq7Ltk6Wf1LB029oIsRpCp94f9cKmfhmJS
xuaEeYuE7qTXWfoHP+symoz+gtd3Ax+xtj68LFVaE8ui/n/siyXRBN3+WPPfqLvkQKXselVRCo5u
gOmn/R6Edn5TQD0eaS7b6z4q8tu9PLbvDM+hIGuFLTevzW7Ed1FZ2uqaR6B59nXVZWa5X6NNkEPc
6iKAiB4lB1LBr54WSq39C1uU+h16JVEhGFr2pHa6CuvcYRGsGrizqA43RLhgAB3DXx0/i3DX5Ag8
xP2Wh8CuD8q7KqrBr979FhNE3n62T2QdutTnUTva+3icGmBqZdx8fBjZNhf0Io5GvTloVKYTguit
srlI4zT3EQVPY5WkbVHVLeXNpuZ76GsCS0YaKLjPmfhq5rSkNROrOh7J3qnfXEXbMGdhej4Irdi7
gDccDu0Ei20Ngjn4k1Pej/ILL8C3hXPNTxhuT8kWayPbInSYAhACSgjpu0bwVvjIhjIKwFi4KyQl
NkbvpV6CQH9+gSHZqPH//tVwazlvLVqlmB3e/vWy4qeMXAZev8ZLhsNp0w1/Pfbe1VWub6Y1b6C5
tfrUxyRbF1ThqMnWOYzRWIsqhJEb0oeQRwdam8XJOGuFTFqUhm15XU0a28UJxqnN3HZRpXmWZtfZ
J944JXWUBsuOljfpoVELMA1DN+VCS63AnH5oHKRJw7CqSkBFa+lbF2T8xcutZVZwP0l2Py7QUi8C
duSkYq84A/An/83Jua8F0+VAnZ/DIVavBvZ/HXevjXHBgk14PKylt74BbG/Cm2BOI2LMjvbYg/Wj
Ua1FxmkIy3n6I59As9E5HMSkuMiLHWTcpinw47kDpqCZUoKOWqSIB1ixJYfZLlC72H0sPHAN+qOd
+fe/tSCGJZmo+u6ntOvqpqFhp+jr1QEN00kCtwfLf62JtXqmVSI+epUpe1Z//BZ0QqMrB2HJaL07
gGp5Qd3bz1v26/gwqKvlwzhoENCh0LYloxKfHIij9urD7q8pTU8htEar4KYdXNRgpQk1O0TaF/El
u2QrreOeelMUsXG9hdY1CySkipus5BKUywROJG8y6Hv5GOzaoa6y5nseVj5sOzqqp7k1z8WGFdmJ
LvQcQCCFEFMm+DzeVbkgi7cv7vXmJA265Fauq+0TtOCHA7OEsJbKZxOLKed/p9xmgijW5aFYsOMM
u+QfJcp7yntPe+Av1ewkdUzZbiC03Baegh+qqtuDERlh1sn9zmYdCvJcaSYv6Nr71tRYZmwXLSt6
xDEmm/avnF+JfttBrORqMImv9bn4+6Bh9NiBJWpO2qq8f1cgou8On4rwe/0dEg4jQUimRd84oJoi
wf9yPUX08jNxQSvQ8QDoP6QGtLFWr2bMBxPVLNo4IgQaL/eJ+OvowJpPq9WZQTELJcBHD49U8S5i
kpkjJm+VNHwyeM06ZOI5XqYxKggxAFEL38WGzKkuq3kFO1iVwaUP8YkxxBabPJqbGZ5ALvjEukTf
AXWlF8dzHsI9GRKoP+VYtv6tOf/5DquP4znTYki4uI9UIAXRjuxxze882vc/BoC46Z1qPa6Lc1el
cpCKWx4UPIM8o9hl83BYrJUYcynqKO9Fgldpq6Xr3yZB3gTQDcZV8x0bPlswbn4AjPbC1i+rJLRC
F91Me9aeINXW7DRBF2UrG8ijWJ8E7DQV3g6WQZLOdStzO1SUD9R0bGLblJ7d/Ls0rZRzXmwMveKe
7DIz92oknfCfIWzz5oiSI+OO1mOpZUienvzRQijorbycTSNz5+/AIe/F2E9tBdpi4ZjWg80bC4nE
0gjWZMG61XVNAZXBXmmTEzKijpgDBiqd9hZCUyBaJuNUDxWfa3OYL382UJsy90qYveVSF9oBNOAJ
tzxj1TT1A6aUdXXO6VDhaOK1pRS1F6TJAoIhBSD94FvSbLnoUiphIkfK7rfLRZzNy1WTxo3wBRsF
fxeHwJx/BjLtFv7zCTVgkHAjfFel8FU4ON1/lNAnFG45WLLXwxyiIZg6OJ1K1f1ezvdjyTzq8Mc5
u9VV6V/uQJrnj1sIaG4sM49oQf0vj9a9sEn6yhm+HK3uC27opnlFuHNsVC33eMr86CkTO5JoJvj/
HeirTmL67djYaY3dJQvAPogRhhbBwLhrhYVR2ta2Rxuv8ntu6RY83xXptGyaZt62+zWucgUFA+c7
BAtoNE3y8sBZXEbFOayVl2QEtzZzvcEVFCBNxEQKQ1/BgKl608cq6vNNClSoCivFV53ucmrmMYHD
SYcIzpWd/G7yCld8qHGgFBXS7QYnGjKOnS5iSDK/cL0pIfmjk3Jc5yw9mMte4oWU4R3Ekcj8wnfy
NaYMP/dsKmpP7BnrVqEIahn7soWJckruT9dsCw1biFsPxQ7ESWs6nFc1zN05ggYUyB2Btxw70Iev
sTMLQ/te15UeuYoYmV+jdgagiHcpuc/NLEorDmAkGjq5hH9DKIJF1HUMn1hHHarNTTfuyJlfuNZx
FZPqBASXZ8RMSSUZ71gz4DEYYa2G7PPuY08P8SSJlOJ3NcIDXUK29Ts+hEc1VPn2lUW4FpMVrvzc
5layAdMO5wLRPWHJxf6vsB/2kH0GEWfaJpwjJWg8dlTltUKPVV/v8Qnt4Q7jvVbYMgULM0wlxz/h
R+wzZgJnjv0WhNoBf3EVOCzR1kT4qJqAyN1gC8uCaTGvMDrSPo+GdcN4DHwg0UmFX0kznNCMBm5n
dO1zSGYCQGloaSMY4pd3GcjeAlCPMa/VX1d2nLGFfpYE4/l5cifkOglCx9k9X8DK4TDuJ9+x1tQl
aNmaTr0YWeAaTuKamVrAM/B+SIBXGcomFly69qVVTa43Rda6imFCz4CvOJsMLkX+8zGtdGY2uMWY
L35Q9dkkfy96lEd/wIYt3aQi1FKou0SWXYUHo8P8MW2KSAjNDPyCIEtjON05ZnslZAkeuo8aMf7Q
86xT7dYzKtKBbfpaAz7vcYks1ytXqyF4JpeaHCs9IxFuIL303PvjBrToOjLRAHT9lKWrrMHEJJLA
z0NL6DaSRCkvU7tOtkzm8Wif8nRBUfjetB3eaqOdWfr23JDJnxxcpbD8n16w9/jxcgEQZ7PixPsH
zq4uLPuBLFOZXdwbmBHUuVhUmb61XDtwMdjehAfZ7o4f5Km3Ijwtm2cNjiNLFSgdmhZZxwHv29jR
uqsL6BAlSJ/L9oN/xlBPvxP/19YXEbfuWAVyQOnw0WIi9WBmkNC6/Xd/QUwt1c/Y/iWaf2lKDX/q
/7f9N8oNT606elI0L2oVD/1piojgvMJZJgERu3Q8l0uLgk+6iEWzaDYwER7kwWg8ZAL1veBzhErC
LHfTEI8/BtBPU3D5uacBCeN4TINwErwsKnpcxozwzNubzEdCB/gKxgn1mSJ3eu76cnhrug1cLE1g
wlxGsfqQpCULq4nI09Dx1Y/WNRKLnmz4RuR2In7U5cKl1lWMOZ/PHyDELfCFXa+EXqt0QR0Fa2Ll
kOzB8NUypEuwQZmmiEQPpMM81hF/R1g+uy4PiusoA0E5sLqU4+UuK6ClY0qUCYsV0nAnFFQOp2aX
BeKonyjG/UF4tPZVpcLKc6Q/OlPpQdFHIyJHpWaIEq9KMdPuVtAqc6G06IQNOp1v6i24K11BM02E
Jsp7lUxW3tJPvNq27otnl1GNKzrYYqxeLoCuEdGqTpK6M2mBmUxC1VSX8u48SocjnezFf6Y536dw
7clx0xS1YkmIgDMVeLpBtc/nDx66O2QTThM+dsIFm6aAW4dBQhSDGfSoW8rxgvDJFhy+lFUDMmn6
o0xXHk0Qy9E8/j/cxABRjVPisUOofp5tTj6GUz2x6IRoAYghesYjhvbfe4LD3brHb958rGrHMcqT
CJseIHierAwfM59KLsEFpGFLlzSMyUR08P8SJ6xok8VGgO4nBhyYf+Gs7MRXqI3jsdjBWLFaxU9A
S+xRc2hnWRaMhM3CEXX3fZ3BPt9I8a9XxPSGq71e4Zsry9f4lPSNaJd+sbkvd3uRQYCb2JfCMes2
dBD/NaRVwue1my8d1rs6/sLSq8EziBMsZxgtyrUo/LOAS6wCDHi+2AQnCWYowBXk9YwRF+VCkCZi
7N1tZVMRyRn/nzJ2Erk2WW+z8lficNxMkfVdruSZLwI1ZhmCtJkSNr63bkGKdPR5Q57moDWipuXN
drUZQ3DEjrr9kpaltwQk9vM6ytWTZxBV05ds3mD/2oswydVDFPpZr33MEl3G0kDqNMqyJCFYAzpo
Vimpy9UZIa4evxWfMZ0gR5lJCCuDXbhKC8qatJZLk+emAaDqOqyO2E2Oz1fcmV1yS1K3C6MosG9F
yixi+ELwKzI05sOE2Ygtwy4+rHl8uAA92nVTgsaC75qR45oA0A3BQATonljaszXudKTOq/O14Axn
JVzUXM8gZW/tZKVSVZu51mpw9ajVz0rlpQ4rQdH7kmvIXSwkuY/aEfj+fFjeSE64bAt6wkEeQuhc
i/5wUnchZYxbI742q9Wp768U/0KznZWDYPpjfZr7dn5fC6LwjGe2jNSXlAbsa24o6hYEXuwRkVpy
XS/kfBWFtB5uyauSmY6YdTDADpH+XbapnQNWs5LeBD9oRhGU6t1wGXAP+xAG7r/25fb7R+iOyBN2
7oXaypBqHnCL9bTLt/lyKNvp/fNRJAxR0QtPDOLMgS2fnKYo+Sq1YdSNfwwUahN3Uf0qTc0Y+/nc
d3qnqH7TPwSHI896kT4cFAAt3h8xR0TfMJnoMNJB/8omKmhunMAER1s/GdoZiOOk0FGyTTt6FDx1
B4rqrIoBvE+JcsewBpBLRdJHgSwGERjR284n70MRW281isGrxswC4JuUs+b8au2FWH3uNo6JAdeB
tF6bYkizKwlraMbWVMPuFO3NunklkhiYz5X39xKbVIsCjNIHuwOkQrSbUMxuDvB7LWAfU7OGB5zF
wb/b1ghV6oQ+hyKCOCgr+kBi7UkOyKocA1bPXYYj4N3MTcGf9iaw2gEMae0sJw4FHHrPomW+KkzQ
S2/l8SuPnqJ081IIQZjOGXeax0OOa9ATB2AKFd8Vp2RgP/ZsW1Po3CNFuPNOYbBNXbwFenETR/QJ
ekiHTgwyuoDI0zqHxAsDjEfPUQ+xWGqgBCBxu/4vUoCnnLi3H7jUfTiGGzIr1mEl5OqGHRTClOHl
TNdYzi/sO5yCjhMJKD6Sd3P3ir/Z6ATePIlAqcxi0ZO0c/1EPWxRIfAM7TinmjRXzfqUkF/Ro5n4
+2Sv4d5ncO/R2HeW0nErGXdqLBa5AB4321k6FnRJ4OxDuP+/2q4iYpcOXzVVdDEnhXUd1/vz83Fy
pOn+8uqH7ZeOB0QKHXtS+WpkDrMxvuMsbWCpWoL1L1j7bbDbebeP7WhcyAZL2JO4qNWIy4bfqrIz
GVwq1BxCxTXs9KrOhD14dJjdmxe9HUchRo3kR5xNQ2TdxnjoaHWwz12ZDj0XjkS1sQIQhly0xIy3
20iSZKzYo1rP59NEYNf0vu0GFd2A1PVqk/Y3FAzFdWgM6gx4f4b4MN1pDvPdNJKYGlhsuDHtoqmA
+aSkMg8Czx2BpjH+M5YSC4t3y2UIs39ffKpwg1r6MB3wvxSPh6Bw0Uu/3ZOnOR3uQT29XG8oivlN
g0P8KBPL9rhs/kynSP5xUhT6Fb62RbzL6vfuJHupnUnheL7i7EIvrenxawfwylfs1+LwwbWKfuXA
tJVYV3b1qyQq5Vru+XLU8O7TJLsCL+MyPJUbtBjYnSPUG47M5c7vyMAiwEnb9XLTrrVQPb5WN+iK
ghvPhQt04CyKYNA2mbg/xvHI0seXl+ErstjGQg8ntL4ILItdQRWN1fjeZeGwn6t+IRrZWUrCDdVG
508sdxR240Z/X1fNza0xmQ7teGnJIAVAHetJ27W2g9X38tiouZJv1qIBpiqmw/gmdEMj8ByOdvAY
tX3tbM/aZA4NIhzZweTpg4oGv2SxUvYL2MUGn1IyDvYC2zvHu1pFRsukyTSpMorRuu98dbhz307o
NlUWXmTcnLx1G0eQ4g+Sn04M4VqHftUzSGbORgx8lmRxSdMVk4OUQSc8Eb2QNfoOcSu6j6kksnkI
KlIUofAoDkPbMI4nDfYLluOFgiy863yTex8i2iH/hCsg1rae2m9oaS3IBa97AfA6pF9sNVE37nIr
HeTtUVrip0/s5F+LdHDbWuKlvsnd1Ql+n6jNE2gPZMkV2LmTKiTQglj0ZPAydvMFBHVH6EBohqK4
/9+j4XW/BzUQhufqGMEqNwWb+OPIBrRsvkvUNP9UtFDyc7m4izWnhLz7Q80c5pGyT1aFDTnGP+2G
dV3GK0m7EvCC4LWjgvH0PHmn9dTgwOxk/1se2DAugzyhL3Xj/Dhl+nxQF77uBJ185ejiB6uun95d
I+r+k0MzNth7NM6DyzssLqLFn0BbzZEDhbqbmiqvgKo9CMS7FQLGcOeXKavbI5v+hcSiyG25yMKO
53V1tTp4PG6+PY6PW0XFQ45p2fTNQeyrGT3tDFF4yq7OhAuehPWzMy5Prd9hSCfYRCy7JprsWUYm
u4uiRNXrzPegjsi5zw9x9xGM09x0MiBSpXdjqqx8KyBqEESw7WJwjIZMqhHxb/DyF5KCQa2Co2Ej
wLWMPb1jkOihjnYGnbrVkn8IaTTEeSMm8Tx0Rv7QOhlno+e+cFkgbVaOrnmsb4KpBHELzev7t9Rh
PYTnOvCaMydiA43w9r9rxs6JsN4ImqI4mc3j7qQGCfE4viGLxcFzRPWggQRyn/Ko1gxYT/vV8AuN
GbgA6EJhWVSbz2kCMO/sPQjiCLoC1N3mxLZX9MHUm5Cq+Y3c8aqlpNjOfU96n1HH/5WI+KOO5rdd
BhHDA0VLNSHQqKaxV2FKujnjuPf05avVljxUI83Oswjuzz28jHTmh5tch4DpFvVfrzVUNBlWiBD4
cRb2ODB4QdP25JK1oieJJx30w8giuXnkTztFgAFCvpfkpMJrhkoFIr7/xWqa/5+Ck7Oz+b+sOi3U
wkYi6nBD3yElS5UTGemue7wUblh5silLtxq0KQ163zpbqVACWMfjLPuwCMVF9xGPOUO8LA5PtjUd
5pBV1lPjttpSsiEV7a2hzLBDMLcmcqe8aUmCDy/UgTvUYqyESwm07FCEo89gfyajARn6oq3Z2g2C
ej+eFBkPALJscJBHIGJ9lRDonLIbAcDhVEH4B4G6TNfw65pUC9PODQKPn1PKhjZg+pUeoF1K5SXa
qQhLK6gZBvuKabr6alJLX2LWCQshBIqHNSsvlyOt9xj8eKu6OIO5Ni150hTuOJmyhkjhkDHgV+uy
/RCSmO6mSX5fAvOwiT7vDwpxjBNFA3wXAWwSCScCEHdx+mEehKkBd/auLTn+zH6LeBGbfFPIVAsM
TLJQTChqMtjMV5u9kcuWJNfwFTEbisViKWXzqsELvmUwkCWr1FyvoTkpTlmwUegAucuy42FJ3Qi8
gmIMh14laag7HUAp6haG8tpDvmMLUC6FnQZxoPYdDMkCWrYX8FzmjKjuGlOPJTgx1msWhBAIIGcK
f0aT8lXKUafgS6L8ih8kFrEqVIiy2ix0ZsCL7CCGiYwDWsaiNUD5KjSQ2F5cvnMmPjnq10cFaKva
v2hS1ZPscdlWx3UPvCjTW8AWpqc5jznkVJeOpABLvrcwag2+eu1oIWThkIPQeGgpX0rIniMEBVxE
CO6SCaz4SHheEJHuL6Y2OAdilt14RB9K8cI4ecDB8c1vEfHaSgiM1/p1r3LU1IZl++Qw3q4gVHRR
HBnQwPYJSpZmZSHrpbQgHiU4Te32W+aGBjmzpk0+NJRlAdVBWqMcG/uZGRcJAcXcT6owBLy9ceyq
dcHbK1BjUMlx891YhffLZWQC9LW2dBvtcJRkypKWWrJVwdYzU8A9IfCur3NgTwci9rvY6n7XR7RW
tEN4N1ZHgNsctZKO1Bs/+ILHliJ7jcUDFAUKdtkeODkxDgI+8KCUfiDBViuPpD31ThZpliOtc9wc
EaC+eRrebsYRAQs0cabqsYPgVBoSk1vNBX6NVDCcSgddaawF0mRljLxGuM5eLclICWX8fFQKLD/D
GZ6bM3oj3uiDMECs/tAYvrY6rDd9/H8A+b9h+/r6g3s6EVr6D3EAI3B0okFlTBO4r8+haw2/X+Ji
/7ns/1VEJ42mN/U6Yd8ebbxPsK9xvqWFBGDS8/2+robpYlz21/mKwNqYti/DjQ0PSHk0cpbmPF1b
ygx6OEPmpSzRtfUf5t1nwXUn6BD+twFtbku6D40mjeG8VLg0Utnu6XSop6RkVNjmWJCROt2Z1/gb
3fVWA5FQozvt88TDnrXt9E/n273HLJAtWGw2s7d8lgsPKNhtrjl9tCEJl/eZPV2j++1x5DqfA9hP
E4IFwWyad3X3d7GP1hZ5g2QKV5zLeGx2ZEAFl7GHKOrJR9sZmy60CmHBd7QPwve2MaQGKz+y4J+/
k+hGbNayglF4x/snD4dYVWTX86lbRyQb7aCnq3JKpPWe8oLeBeCuJ/H+Z7qCWnLMCPfP8faVw6qU
Fljbq17CZ8XoXw+6VEmsQFzPl3+8s6TP6xjEuULkmLT6vYqJLV04miMaPVQ21ir0OGJRLu/yj/oj
wFytLUgfbHoz9Cms4U8191VN8og7SPf+vHMmJKwYHzxVSFRHl8bj2LGEAXRNCJQVmWJ4VtZkfcRx
5ho2wQ51W0F8Xrl+cXyx1rXHnVXIUUEfVQtccICJnBGUUnx9+yiZoL5SDap0HOdr2wICTiwz8niP
TV6qKD63ZjFLADunKqfjFyyNogfj26jugcJ7FFrH8rIMlYjmwHDCBN3jgNHZ7OntbtWfeW80x5qC
NQoXGoXfAVOjkox1PzyK4rPATh4Rka2yCyGQHmCU+Yb91jbvOCgyYji6K9hKKkaKwyUQEQcTguUl
/1aYwm1u02TBTfeAzfaepcTDNwsszSsQFxZ6diDF2X4huXAKK+vD8jiDEbvVw7tBAzeexULjEkY1
CZ/VlyX9PYVQjvr/H5m1oEyQmTNUT0dcJFamrmPb0EIxyRJ3OBpUctuchNumYAIINXTk4nR6WHk+
P5kDMThJDmzHzNIIWzhKRtygWWH2ukdZ2XDOmjHuUJuLJCSTOYM/aif9epfHqJzZSLddlx4A+16c
ClkTziapzysAKhk7n+Cfaewqw/umum9kweqDd8tmaZfTVdQniv6iUGGtv2m7meCC25rFvOm7dCYX
+jwR+u48HHUa22Ln8ULKB8ePyFYMbTqXSubeR9cmpM1q3F6UwyA7NcGAjCB8x/k0Dd9DdrI/5mzg
WANvGguGHZKSK7bCMV28zn9RF2eQ1PE3uvPDvWIH/Cybrok6WnDuGSTEcklVKO0tbue6ehu/BbUp
Km0fiJ8RsLASFQCIE/h7oKxEjG6H08LjEqc4bPZm9AvohF27JXgivQ8fTbFSW807LsZxlLuwPziO
lnp+Qcogb6lBzIP2Wf0mVAmmq86Oxqhnegm3ZFyJbQHAIkRPOMr9yUiwEgeEd9rlQlkfx1kC43Ib
356LRDWl/UmwmQ3ceyy4HGRSLfUWNWJkj8Vyds/7RTssBsfPTkLxJLXz+h2VWFCAywiQ6NAfqrcB
1Bx1piNfT6YRanAY6Z0jdWcN4dIMS3gYpRipQOFTPDmHUhUw965OHXZyTos3lK6UpTCtjIjKRh3P
NXh782Yz5vdZP9GdTrMfB3Z8x1x3x2tNifIuO2Hy9GMU62npds0S7ccqMgw9zUqGk38n7TyJxTg2
v3w5ABcJhbH6DMARI7Tts84EQkFm+zskpMYuwWbOvVq5Oi4BvLRYI/54bgQiHjepsCIjQUgb49XR
hXSh6vWVfXNitwwwi7wo2MLEKuf9uyzjrpxzKfkKCnRBuYX0ljm1K1uUiEw1mvbyGU2WLKq4lKhs
BlKbeD5h3KQ2OPDRQwM5LN01nc6TqQe53wneMXU5IFl8XEFddg53oe6Aje0Lj7pV7BBs7kNyiDxo
7pC3jkZcBt36KUoUA1SBgjWv/ftctRMdtaLJuy66LxO7tWOsCv7cV+gTE1Ao78lIzLnlm5OWdGkE
5Eu9KEhPKKvVdzQuoHYazZCsxmgm3OYYpgiDKQG265sJ14jzraPMhqBm+M05RMS8v9UNYm0KZ4QP
Bs+XqiNEaVjaJezvw3lL3Y1eUiTSqzZXLR+rPSPqoBpacJl8G4Ef2DBkueQNRfM9aRbH1ie7pBOP
VQg7kgq0d+Wj4o1BT+5sBCvpdS425IM4j4w7zktd3xyMvfe1Ts0DdPVaIXPiuCJCvh4/wBisGvG1
n91gDaK3/OjV/1PsNts0fJsqc9Spn3Q71HtDkMH0mLvhmqwMg7T6f40e2gQhyp/Dbq9nC5qHRfF5
HpLUA6TAmhtig8kFSv+senR6om11Ylsy3TtAKmkIMBP99PA8ny6shyU9Au+fS5wFijT+XtSjtDzY
pQTqlVqZJCkXfHxoHvKRFSmnEjy2THfThLeHNTP+kGA+yvzK0K6n8C00AED9GLYYCHjSnTs8UC7O
2PFW2IN5YJ5seqM1Es/D7KJdQvwavIrGgiIYAE5g9assyOye4dn31IOwycG42h54EdffcC1UDBtK
sf1BELXuamOORAPlu39G2D3c/qfkOFo782SXzPIH0vjQEn2FyWXH08GiF8n/61yBsT8CfwcM776N
bCYBVEuzeQXtmvKGZLbmNZubS8dUmAmhNV+mxLyHi+cQYLRTq8NnnC2N/k3fPku/tkwGnBThlE5+
W2Ro+1rBD9CbpB1KhAYaff6qjTLp4GLGSZUkdBtWHw34q5ghLeLh+dRsCaxqwt42tAbhsuJwlNC4
jtG8f1zaPCD9JrVBqcbDsEXfFBLLZM3uhGKjpNwneIRYLsGkYt6leKITQq+vUmptQh2tLPvBWsNx
bg23TqcK/7M6y4AzdFLJUj8VtUaufcnq78/6bFkVkxm+NNaFgjbJiGKQHxdNP5S3SfmmXinOZ10Y
nKLiz7kA2MQXNppI84EQn5LO7SeRzrJuSMhskvV7AQTv3ktELbP2jkIIzZ1rumJI+WPdbZngo3im
3mZi2fT3qDskzPFfKEYAs43dts0S/8FbLiUiwnF5Q3HqTtmvVFgKhoRtLjkHfgRc6ROn7RbuKFUx
Jmz9cUheQ+KHj4yHmx3MA3USQ0uLFziAX1IVXenyFaRKBWgIgYV8g2gzKOe8kwxpN8NMwnK9cgV8
rJ9BwhedxAvL/c3jghYNT7va4AyPXQo0OXLuzUwPyO/eh8fTT8n1aFl6EHbzz3DGTPciaqwzEpfz
UwI7hgk34eiC47RloRQIBsw6fEDwHXx//nfpWhVEzi7NovRWpSWTVqA5w7hWdOWOQHroBsZKg1He
pe098Mueni7Fu4TlOCuUsHVOaagDD4stYBf7P/DSzrSYwd5ZL309XWDdp4SqOZ22JiCesSIvO8qA
Gm471d8HXv0ZGCJ65vhfvrNgWc5kse2qyh1q5s8jAekxequMqE6pUF6hcXqwb82hTRRZ3ucxZgmN
9A05WWLjc1lDqXO/Kt152NvK+a32GEkEf9zZF/F2MZ0do9b3TeCaihnw60FU0P/ufyjqM8Hu6WDz
BNa2w/CPuv2lAmHwa1TajBNjWBeB4fR+7CEMQ+P4NzllH/wa4Kse8HvhV9vm0cPmlUsXu8sLVNkY
/l9Uehomn8B9KVxp/Wj6JZNE+buNBC1QdFbJLFS2vogpL7GszQ8mJeAx5U4RAh4+2uk0VzUEfNUL
F6ylXYVyAidalRQi26JU4FFyuO5qFPv80aQUdXjGMNtp64ETJ3XKFrGWjuV644SqEReL+tPAtiAW
eaEpVUPhtKNGKz5qA14J0QfAHX6Cl+pRnyoPMsIAfVT0x2xnTpb9vOJZo2Mh6jz5ZoOSgwGqF+RY
JF55haX6CspeLna8a+PtOAjcZnc3ABRwoaPvQ/Sh1cqHN+P7tS8CXO0MxoxNUg4DDloLg2sKRt/d
mQo4OtjOzyUX2RXCSbQ0pZCHBOP04QCOrx74BdPMVHjVAHaBlgTgHqwLiI3DIpsN+y7mZOqVvSjp
hhBx4KfLlMZ/5rVmi3X0OiP/QIDrSY0eUCPciaHY+HkTyCIij0ZyD4EB9OC2Muqi5ma8EO3i9f4I
EyJ6lTwKALIMNZzwGCuHwHmR0/ZJE0pcssRfNsYcwxjc1jC+aX0gKnkXaewjmFWUhi9+H49YP9x6
R42oHpx0tb0EfkbzJ+kxBpxtvt6tMYsgsqzAb87vDnqxeFxDx6dRqF7SQfucpdcBneYiO9UYjbo9
jZdbzk6tDaJ2p71xC0UnQO/hOhwGU77RZY8zOh/kpwfS5cldRPp1bg26ZNlpFWQpMQMuuQHeR9uV
Zy8VlPaFRT7Jc44AfaTd5u59tM63Z93ffq+NikI/f5wpRvgjmYdyDselF2CqZdYiYeATmYTWORBR
zzfQ/z4NQVRfj3vk9CmwN4pdBmmpB5WTMvpr/PKQKeMCTI5duUYLQFpa7Jir4vPWhh0lmZ7UNQHh
FV+GCUd19ggS2zDFXoqjfVytyJUiPrYsiT9E+3S0yn/S2SYBeUYI22VxywpbSi0y/A4gQVXumPWe
cS8LqQksOXNs41RGgsxQUgM4DKlifNRRv34XrWlOdwSxd5cwmHJDi9X2bqi3FKX26JdSuLm4gTcz
1VR6/nvdVKPfHZ7aV7jKwsSHJ96tTQhaRrzlGMGBrFQbdWgei//nsI88CGbxNy9DFZ3nHN78yP1r
sD3UrqFfJNfsipXaMZM3VTO6wgYezCUNn7T9IYl+gq/lyKc+CznjOdwShj5hc+GUE4S9biFW8I6l
3mOTN5XQL+AbYqna1sx9LvLA5gq0BG5/e7UQdAIOveGk7FPF2lQU/VMAW62PfrPx4VMwNd+tHlWz
rPL7obKU2YW7q08dtsujgSJxGXrQJKmXaJ5hhByc1dv8HNGzVJ89z94IcrEyl47QldWJ4eTuiD2/
w+rKoLX0jjQlHyedb3iwgt9cTzslbMdxSsKw7ib25hdV60DkZjypSJsvO2+JGOdbclLSsG+o1yo3
vD7+NBY1qVzmfwHrpTysyzIuh3OTFGSTxMtd6JjQ4A1PANoWCvWELPBcF32q4QDSB/eXw5K6s7Ny
/TsncnfJdzbkWA7ZeDYrd0TOl8f2KRWc/AYGrkccnRsXfpoepMCE6yrE3ul++JNjwUcxGKJDc1LJ
Kh26H+mpFA+npGLPpJCtiAKnugamVrdUS9UJB0crkpb7qTyo8xz6CKoFYQvstut1EW+oaaQezUfq
UFVsxs3cHjM+z3i5Hn0dcWyLHpeFrCbRDXalnHWXHyPyVGU6w+n3IZYK208OGbLx6RE9MQt3oq7G
wo2Pehy9RfT5Ig7kP95l1ThQijTgRH1GoZxwZ6A11gPTiCqWwkCbif8yYOFNlqnfvY0BmfabwgmX
TRIfvu9FOVieLNfFiBkMg44TINfw5wC/zjocVPqzf2s8P1HePPw1HBceDEcJRNJc/2fkSJFQn6oE
2+JU0NDl09LqN2V+j6XjDq8hzi+6Y+xMbdz0UQ4VI4lWRWJn4u0OFlbrN9HYxF/nfd1LRStiImDN
du05bz19uIw/MXzZKRfwaGBPqNkwXonYyRs0vcajoWB8D8GHfEDA3uY1lIgm/6j8G64BUeRFDfza
kbW4lrCvrppvi+KGylmQgqISMZtgidqPBuPaCZeOs8UkfBXLaaNZ1NLenVoRHOusJRxvTP45jY/e
yth8+eERPfWikEXPfm2V+1RjCAtMPo3ZtYbrx89E58aZGduOifRapczqzTebkj1nVnTdeH5D1yr8
RQML5nbVqNS8lWNdF7OgVuxzF5UacXXeETJxRxizotnr0xTqOIavPMTv9cHCzRl4E9wZIKbPBJ17
emF+PwaymDd/b1v6KjmpqBlCRLjvL6IuCnhmjS1af+jiJEljn3xtlYFHxCmXt7V9FrH/xGXnYsYR
xBp7n8egQc2GIQk5pAm/ibUQwrMXPDdPioapQTV3o7A1nB9vHn3Z26Cq7WjNWAkUk3k+PrEWi37e
9glUfFgp8n3kW5sLkD175X/FDrzMUqiMAaFxHAn2NTdzfxjD6P1aXHZ91FbYEOskr/hw/iyR7M4L
ZImQkxX3662dogF9oq2XHR/B23S+ElKj/FvSlXcOtAgZxwIq7h7LpjMrMjpmbSuVdupS2vzknIzt
6RLcvos5wn2/9moLyugUBl7CejpA8LQjvnDUNGJcZmwbjP1ixJsMGNFpAdJlXibNSczKsBAOGuLy
NyHE3QGU3y1FoFolGepeAKtn5hXFWPYOYxP1u1I7R1+KhmylDUTmeHs2HM4udOaTYQ1FXXkyEXnE
AM4BLRK1m6eizrhizCmu+ZS3M5J0CEdc3HmhKMANeP7te4XJvNSMV/o/mxm6dMZuK8EX3yPYyhk3
cY+MCmTanj29Ws2Hu0FeDxySat67q2HLuX5eJ5gyJdvN6xNr/Dp2WZ1/zoRuf8vfMS+xVaCHiRMQ
ol0bJaMXvI9bXvPPyO7EN2Ye1Ei6ZPymm8iGeWERIFwclhu5hoZMJxnDhj+vLkUFUZNbJ6wU3QG3
F5ha8YH9y2i62QFQH16WwgCtS24IKa8oDfLR1xAXmTvPoUBNorf8dFRgXjSly834PGipGZr5NF8J
VNtmKWYuTrqlMDb87BpIHt6X3O2O/LYMSqncQErohIHC1rGt5jUEEjv1HXj9bO/BnE7TcEfyiRXZ
m32c7LWwFbjjCvL4p8xymcYTgQvtB2LXhPXKX+72W0IBcTpCiekiHCqMzu2M9ty8UsKgN7fFnn5v
EMqq0q1Fw4EOHpemdRTpDWDJ49APoRMH6J5NH/l3330ezWSi/QL6wG8ETjvquWe+sKnb21hTxnZH
WquUU+RRdV9n8NyMdd81Tl25GU7mnwIkIGSVmnv5iRyMSd9ulA2U3YgsjMNDSSaiN6jq6GCvkQU9
YSvQbOGJNEzuVgg80XC9bRiBI8fggAHCUNVibzd4Wf2FpMHqs60Sm/Ig396Bznm4jkR8mwtzoW20
9C9R+VNuFQ2jKq/hTkRcUVg7vFWyPB7sxQPHUrJg9FdS2gQjo7dh3QcDLS71jzRhBBOl70gSkwgP
OdeRdN9lJovtpoFmnFMCvjPVPVnziJYIy8dkgGuLvbN1iKn2YzW+lPFm3YIH/GYbF7ETK6gCeKBT
9Pl9p0Yq79g1misvbvA2mPs7fFkJ0JjAUmmloaIzrSEAIvuFDlpa9nZDLXCzphm91Pa8keGtjDs8
It0zel2PWEKth15HpiSVIfAmXCVAGi4cvWM+XQxRobf7kN1NXR+SHaAmQDdDDtlx/B5kz83h5g/u
7/c3pNvakG+4qiAFicJ1GtVdQ1isRM9J6s967M1TZmU91xcjqnVMOqLqv+lE5mhUk+wn5nOT1GkP
kixCDBQs++BhG3w+c9y/Fg36Ox1XVk7TvUbRa+v7pQ/Z8001M+J+59DTaOHG5+Et5Lg6PiRDpIq3
uBSsb2TB6sKVlfTe3xL7zZQ4Z6nxeVllc8ZbQjny4fdsfhKR3nrKrfYSXuJ0iDz2RlbIMC3z89+M
KVIxJj2D6VjTzF+kiD0rYByYyE8M9Vw/HaJ+zR+At6z0upekk6cidF8MwsyVYOOH/kAupIJEH338
oGic6bm33h6ziuFaLqKf2BLtcJVKNAJPVf0pqcFiFZS1H8MAeDw0beTZ5EDwVYDYpIv8lLr20tXE
JFY/7Q+cqJE3IijJgcH0NX0dB9Okqlck1E8+bysTP/g9Al7YW9MpPRaHma0DOt4QVIGdvHXRyP/t
jGl3TF8o22QFzlXO+slFwFIOQU7kyRD/3UV0TROhYn9qE53bQEDDxgqfGvz3jwPNk1ZYJe8/Sfqv
NMGRKmy5fcHoCs3fpJJtoxBSWV+gbP+u+Hu7Si0GKbaLMZnwwZxlHdfq1drHsHgyCuMPsUxlHSsJ
Z/51651mqpav1nK+DFcH921p+qp7HILgi9SO/2BzYZPmdDrx/TaudcwYYxon5pdHteAIpyFibZVg
2K4fx8qUCYQ+W6XGofuHmW2GcuC0vgDQnpzKJwE3SecHOED3s5FpvSKoamNRxJEZXSyDyWz74eCS
VH+zUPyINVGdyeDNsPWzzaEdNfkj18JauNyyPj8HowTChMbt6E4LmcwB0svpCl9oL/cApgOHGUoz
EZbVsmO1S9ELiWrDjnsyDbEbInlirR/tRMNUof2NZpRRull60eEp6LwOek/4iCyFj58bLRa7HWb5
d5G/os9RmS0V7Rt1CdMh0eTfuynk00Lneu3uqdJ8Qmlm5pHLIiOoGtCny3aP6pxSPXu5wcw51L/s
eGEKh9O+Idcb9Pe2JSfAkX8fLLduEhUWNchEpGL1GvGpOyqZ435xHl82SRpOVnWm06QZAh1o1OR+
fd0MOc7EAe6/X4OUb/Rhx/yksECNt8zyUxUIV6bej7l0GqobbCQCQn8gGEBZEJKqgg2scM0oL19M
FEsbAYCxw4THKiy07jOj/7ZFVCJ8dgOMw8R3pk+LTfzUvFiDjALJ4sngajHDuSyX42EHOnb1Eg3L
odXA738O6/oi/JDo8/HLN6pfM5CwvnIJ9wJWVuChl8uvdK3xe3VFUqEo6my22jb/8y3pMo5O51xL
c5HrcBHtt6Swx4yOsnd0oU8kTruFQPUr9OzMG7WxhCfDBsVsTH0Qif6V3CeRpCcrCtWXXX7MxTtR
NBvEmzCWs4dGBfMUCNBZf+DAkt2EogoCgnut6ggMN8b/yl4omkKttzX/bl2R5KbExZHh3kImNhJI
U0QUD4i7AQhnSwtdPHmmVUSyr8D0kraqUVkkjQaP3hvIx/PzV4dOO+L54DEqNiJoby4AvCjXJzUY
yfnWN8ZXN236ZSM7MXIEVzvZJFCvaKwm1yIwbscbxOZX8i5TlnWkyqHLwqxY9Nc4HtDzoBuIeovE
NCfUPVUA41YZP3L/VLV58fAcB58r5jXZo7LhS2CkDvA0NSduK2KAZnpV5LQURkEF3QctNvYUTEfl
bSFfxdRgE/bJRsyNMKPhCDEYnv76PkbJOatF1xol5Yyw26tHWumxNrMBy2D3WCwbCK9Rh3XZo8nb
Wa1sb6htDZWIwEEBHSX3+v79wWVuZH4wp2/MFCISCLkWyv5TmyCNX4jzxSPB4SXzmF3pGdLbU8Jl
2QbVfFz/ZWsP83yaKpz1jR4Jnm6Jm5ndXEEHAk4byF4Cw3NSACy+dmNAAwPfa3uoCx8nZuLZMVFY
pe9HMvCw+wRfnB2l5mJwxspmpL0uOV6OtWqSTPdgoEe2hqnoCk8zccqdkPxJpsuUsqOgRLGuILRc
GO+e37JtdH86uFxY/gH0f5YHMSjLYUDKdwqM9c7HJ1YPiEkV9BUqJcRvCvu2mZ9vVnqqx5AbY2Na
8+UvXSKU3wSGYdrpQSUo8Z8f/mgX6GoXIKvQivkP6lGge390vFNX/SX+KtlxdIULMSeGL1ApcByZ
Mi9hov6jBv5pNXp3Uv+08Y9amWhqOM293OHgVp985Tmh1ZXYXytw8Z4nHf4LfFbGxd2FiQGys17B
W2EgKGJ6lH5u0sa2rAh4ca/hww+FVcwI9qUNlCbVQNtfbWX0eAlg2Y6NyyY1sqJxUPA9OuA9rN3e
m6ssvZE8wrrpPe80WO8WlHunY98j0MXKSvvj+3T0ulCiZWNU7Xd2FYOCuNv7ViwBKoeXmxSngfX/
4JTvFv65VpAL/FvNxZIN3rzg5HReTjwm3BDkH1kbUWMjRZ0Za4Yed3Zqgxz+0nA8x6I0KsOvQQCW
Z5RjfVv6nz1gxlpuB9Azx+fwQ0bDOZqj1oGtGF/Ya77s1KbO8nCt50oszAXGlxdDqEb7QnwwK6v/
d0Fyj9hyafYxex0PMkptAEKNyumB1WjELQAvuw/96X4nf/djm7H0KQibEIxgn1rBfJ1NFJ+xMUYk
mkEvmY3Q7O1q9A/sRt08w4ncCSqtAnUc+VpRq9b3kB5/JwZzEkcsrxpd8q6R+/OxOPxpInRxkQG+
C7LxyjSro3fL13HUef3XnYg9V/vlUYmTf8GcDDNRRHBRwOTVwUAsRHI1Mct4yYNLUrYYZ1pd7UY4
ut1RF9nxz+fqizlNf0LYrwpYNtp49DMBVUnGI9rMrHPbwxpynGkgVjkvdppuOcnFNFcHMG9tI5yY
iQtCSNcwZE5s4iER1wzFfcREKciH0nyOvcXpXWZmQhDwlMRD8E5zOpEt2W9OKKv9y8cm85EDBEDe
AL7WgOogW9Vhu8cel2X0PbW7wwKnr7HZRS3ckdTnY+4elAoTgfKgbtJaL76zUrSjPrpNgsq4zVOu
lNVaMdw55f03F88C1Nzq17073VL6m+JtdjpJUZEBsuz6Eo4x9mcIl1s9IuCFZZ7QCRcVSkrtYRI2
7VQpGe2Sk8cskcnV5Z3CJgZn+VzyTbG2qtVzXROUzceO0p5bs+dhCMC0IgC4p7CqGKuSCR1mSY8s
VGJb/vuwXojjcn50pzcAyn2DqrW1L+SppxdySliippameVZcke+AOGnT/zcDP1b28AWfI/QHSKAc
OZ13dmJaIYj/Q23XnILEKiarkqiMsTfhxOJBSV4/lXmZYc8DqtHbTVuInKds14CCYFF5EzH6k+oI
Ofy8K7NRE74URMfvHYZbCw8yVWm2VW04n7M/gw7fyo+cVI8BiaeyurQe3otTxoemD6Mf6g1qvdl2
F9nllsNJsyWMjKtxUDkgt/nrC56bpWnRGHE4tGbPIQq2LCI26BF0lRCWIOoDYhTGic5eog7D06uL
1BRETDr909lk7RFPffPxPM4gKLImxZfWu8pnTkY4SdFBuVQZYM39jQbJ26Jy1326qUWqpz/WSDDY
tylNN1Mki/v1vrC72LaDqdZt1g2sJEqdj6lHEf4nkL2sr5hRznXvmlXlbvm0KVLU/wZxjauywBE4
hmBapJOVtApDgarTPp3Zn8rhchbWyxR0rd6p+HKkF6nc1ZMdDXJM+LTVuergyD5+57z4MtYufXnM
y6pQVDIsqYc1OTv2yXoYGp5Dq45qN9NwxdSGPWnImFjYNOhwICsQCy4W4R1iimsrC65dHW5td7/Q
HoPncHuSU+ezLWxBiIzswlWDiLkWZ20rLpbnG2Otv+hSecOJZmG6iM8dWJWWb0KAjimBwAce+GXz
JHhHmWjRQbAb3RmkvtRKLhvo3y6+F0bw+L2BfHqiWohkZlcHqe531CI60IvMnv03CE4OGimd1ETI
I+S3JCot+W1q72AqIDieFfqXd5DpBBQUtEeGiZ2V5OWYNuivr9U7o61n30VcFQbDXn6W4ZcSCJLw
ZI3uNFoM1BGxAKyzDo7wAuYh0dSVHZmmkkIYk2p96U+vPyc3ckH1HUDNTdjb2L4phQmc6WTo/iIs
awHh2zd8nTFlEcEQ5sKIvZcEDdPWnYn4TAC+TTbNZ/oGhoi87Sc8UsIU9B4g9WoHO7SJ4w2FK+Pa
t3/cHwus+kSQZRsc+EyTej/bpbMi22X3blMAatsR9qHOVEHbmUwHrrnB8nyXT64Mm6DTP9gH06XQ
E0PqNS9dTyK3h4fOg81Dvl1rn+Og9s63xHezg40IWe2Ylcw9LYS1i0z1cGBw2YJOR5R4qCvOHbKA
vbSelsciYqsXwQRgGmTP7700BdTw3GYlpV8y6P+XYe+YDzfYTOeCqDA5MwQ1KxeCKcejZrwpsTue
QEy3AYD2wg1AJe19KBh9iUXERB+QG31bt91y6SwhF+MB/gGPX7sFK9hn5oRZeoEnAnNDMVYeQmKq
+2fN5hTm8FoDDJTen6RqZzndTQ6lf26ZSBgeqnmNT5vXy0Gb5e31rP/tIdELpfYe++xJVXjO0pmG
QDd9HQPCyhhpaYhmtmvHe/2OHvv8xLB2xb3SYId8TUDYcieuDb0DXQ2xaTqqIriljqvI2U/VuN/r
7xjTrFzFd7I+erHJp3No9XyOUytdTnoLU/7crxI6yT+mhkO7bT7Yv6h738DnywvPnr2MMGJtV2FD
PDiRuDPVlwSHOFg6WRm33N5qkrhcpxrvqVYR3iLRyuF7H4QtK+Fom4MXpEufoLOnwQYvDp18wD21
9g2vcttMSHWnpR4D4xh9ptbGX/8o4ph2T2w7JXCZ9FizTi0cwRfYzfAtZXQpClFHdA4yKFdDNjFB
VZE4Ie0cQL3KZP3CC46Vg+OU/kSNesJH2hs9Uf1znOeTVFAJixc7JWKcCI6oALCcPoMKGq/C61z3
C9FhLLUt81P7hVHXQ8kj2G9LyENa5Rp59ocYTOKdL23AtjDRHT5Xyajte+RTaPE2Bp/ZDAQM0tqM
xU/d0bwded0eNsbDwFFga4p02B5MnbQR+N4cKH2MgMpITGdin6iXhq8FLG0BoEhyxiCPWUilrxD0
EWa3KPkDVLaait2CzaVlj99WY775WcOJthljU7ZFb3iHcXLQp1aPV9M+Gu3kIgLYHZkk432dCWQs
HMC92v6ZODGgqt5Fp4W0s9JQaPmV05zhdhioAxJVGfGU1lO6THW4baTp3T6jho/BV/mVagJL7RPN
qo2JQddIX+IDFeZvPnXzlKi8WBzmDIaeh83Ns6wmFW4EAiUpYLmcZ4C797iCXsHdhqsIaHdiXGZp
DTRh9OMBQhb8BlRaCHJ6K9G+1GI58o6GGyKahc1H1NICG7ux7ZQh7h2NsTZD/qf+q0GGTzTEKdrr
hGpmKBSmoaxnsk2L2WptIR//xInnhVlZ7f9PpARfOz+uhoKMcYQATHWz02Cm4NPN1I8/+QAjwneY
gZ1U7oSBYeThXE3K7Tl0nbGmIb3zTrfApYijziMXHI2e7j4bpwO7fhglACU4aN0y1MTUKGWm1AfZ
P2k3ghm/UZijqiwX60oKOtlpjr/kopOYRH5na5Bki6jvs88CQoMhPP8v7H8KT03OvzK2seXudNyd
cPTMckk06V1fy3SuC+oEZOs5XQxFgWFTBSe0+W3MDumErOoUM3U2IcG560blABlCYCRQ5P6ebJPI
jtW7dm17q4o4EX4udw15oxfu4vLD7mocIXUtnCtOI7KuB1ggwhChNoepvKZsGGeVzaFIqIWnMK4R
6EdkELhFmQsUShLZfziNlR/1cGqWdmVKVpIPa0ko/Udn6C4tQdcWr8Q9kTAj+TVW1B5pUl35zb/N
Gj8TlBMcUMmElv8qNNZ9321RuzzeHzDBtMqaaTdK66Xmzf8AHpMY4LvfSkouFF5JtnZ4166usBVG
/b0emlhAnClR3Lck690LIfluTcDo8qPrFzFjP+nvhHC/OkhWf5/mA859f6d3kSPIV404VhpHDiXi
PMQq22n6iQFibwbDPuCWYIlhR29rIrh95zeXBEg2L2yKAGi8cog9GQqMGqT+8DfBLCXDkbOxbp1i
Jhh6b6BPn9qpEWaH3/fN1RyEs5Dv4e+ggnhJaPGGBfcSO3MAoNjgOQo9L7K+78p517DyvqGKLu60
18mrU2mtWV9Jjrj/ySzAlAJ1ZrmsarkbOvekJZHJiqvyLcTMXUQO0j6BfDrThy+4N4ES5huNKvQA
7bxSLyFbo8Pq0QfRYJ2F1HhZ/4HUBtVnM918HNNreSf+pukPrROXIFzn8QcsJjkWPejTYPep+STH
1qGnXfFVlBEsCo6I6YpeSpGIWZu/D1rr3lJfKETAuHNhotaKBYN7NIqnlG10GZ3QVQNSt/2Udl0o
JL1pZ5L6rYNN8LuGqYjnB42GxIv1yMnwUay/8GhzTVOrS3tYtrBJ6wEn7UAU+GlXd0ljO0o7bkCY
zCsfh9uEYbpJzLehwH0xZqCyLCiU25t2S1a3Lic5cSoKTUF9b5Py60j6x6LCnOt0a0W82cfI1x2X
Fx/C77ha9NSQYS7kcDcnNrs5rLnKAt9D4HEoB8XCulHjwPqri0qJdDSd6l5qfxQBFkOX+71i4m25
xi5+FfX7Vpfr4soZRfVzTgHgOk7kD/u01YvE7tWNgCL1hsm6Ai/edXsQm2mXNCj5gJbjhi9iCpsp
dx09D7LTeBbu87MdRqPFgTJH/NWdfFLg5bPZZgjJXDxZTOKe5T7Lq7Esg7EsEC/7mGjm76EQyVkF
mAQNqpZoPVeji+Npl5glC/XYazFmvZ5nalebt1hdJRC2YrD9RkxJmQRHpzX8itQyvFN126x9QS/w
0PsELEaMpaI8N+yqNCOhPwwoEpy7Dxo51ngEKud5oYZwlGeAxXd08YqSbIGD0YhViqucWiwWcGZk
6cboYt4/rl7B+aGhZ6EiY0L2N9lLNITBY//VC7m4H4lZkl+7zYokTW+a7jzBOO0lKGSnILrE6aoN
9HnbTaylce/iwiWuvD50xeHvjs4AYNHqavFEcvvyZc9Dc/5ETCnkvxkY0DOcFqVXmqwG8oMdXzcD
G2+4uwATvBixNG+XXGIKZ0r4mH9ArQjhrkq6a6lQXACq95yTrOhVhF7J9P/CCBzdaRudm3yUkD6v
Th16ot4PBcpPSouQpFZ36EhNtUYNfCXz7NZuzxPDL+5Wrbdc/2FQfdZr6m21DXrD9c6+igcq3FUf
2FVhLYq0tB6sxW3w8uP3rFnljE2Mc1WGIi36cLlOGcYP3NgnfXMIRPqFJ6M80T5HVMTbnoqvTMxo
V93DVxtqE+PtncG/sqJubqjBePAOemTsmd1IwaR4zLg8vuPf2x/16vGZmbKquoa0rG3PTI7/jOMQ
F9Fw4hgJz/nF9H1J8kGU0pdDr0LTXUmjNvHFYIUXOljNXiNZGrT6xszRWCXfKiFru4Xr/HlVt2/o
duaE3gkZlnTQmwhFBoKsM1EA12QZzz0iEnMOCb2wDXDf5gCiO1lPfNltJToqq67HqqelMSszxxcK
Wd3cU2VqQKrmEitUuItLWNOjVy9VxcDvrPCtpCrfWdnIWYQ3CmhFdctuXNdTB6w8ch6/xJbGdVVS
gYDC/kRYdJLMrjk1JIMlT5Zzd93R1/54FcXP6gsYh5yRcOqlMI0fCR7zoH0wOol7j66+zaFtd9ir
owYHyqNlDOAoKi11Zs/2DQi8fRZfAP7YPNFwHfy8xYlsP/bpmYpzgzh2vaIS/Ome+vIJiMe7AhYp
wSNqFbtUcZkmti7Sn1lGrv7HkIoXTB8iu8xxyisolWhjfR0R0JQ2o3Tmbi7BcIPJMcwF72y3w4Dt
yVpSKg9SkmgNOyyxGcXNhU+T2KDtfHD/C9GojaOv4TLgIoYpseACxezO+Qqy5jRScyVDqulDXf2c
ajtwkduQ/GtWw6AsdwZ0JIYoQvNGFVurdCtDTUtGNrsYQHMDMCfouZ0oKWC8/VVdDhjwm7qW0ZFw
896WO2iV9mlGyi9YXnmXDKMaZ/AQ1POiOWyN1+ABlsa8o8ynmiIaOTMxotbUuNdcz3lHNKZFvoQI
PMpfKgFsq1fjY8ByQJxnR76VAbRireCcqFrk6dgGpQb6V7BTrzXBfh/Wwwww90yK7AwayqXa6+VO
8R9DuQ+yWAv2/ngAJx1WR7K0PXRIaI66XP3wPWoNkEuOv3BTHNixH55RZQaDllf9MSFdTiCZ8o0C
wMRs6lkmeQ08XR9wlj3pk/jyM/zvnkxmhgLcdxoSir+oK21KqEu0dGAwKkUaGaL2MM1oNKyjO65r
IZw4t7FdJyMnl2jhcYd1QNRfylYETYNByyb0rATYE4lXaFOV74vYbsAxg7LL5dJAvG4pEShK6rNo
Mm/1zpamD+D71dhtyGF8r2W6JY5OAz27EZJkpQAmI3fZXC5If9ZF3r30k5e7/zQu8l/Tm/JCnyWb
JYDTX8vTLpTR6WN8DCVVLaQ3OzncSGNUvpzA3zmf3naOLwNKUXwYB293TG2OKmVdZbmw7QqVWNhx
P3/Lhe4bnde6sNY40yacyTjvPE2Evwifn5yY4ApVlKMNnrz+rBLroQ3I7tgwKD/bARJBpxj+nHzg
yEvo8ULGuhbUoJ6zIPY+vlWEBGkFH9shfwkJ0vrcl4MjuTc8QUl4OE2+LkHIsNsUWZ3ScRYxX15f
i1YgKZkvtYWgMKPw2GxRi/10iNkWFaijP+/hovZnipqIL+5sYkgWgnANljfaNaF46FXBPitu8HAd
slj4AS2QVNonkolzxW/bQ7wbxaG1MlaQ3bPPNiVKDRqXzEi+XLUWYJtcPEjelXzPp55LoM1rT6+w
MhA5YsEXyIb1jq7mdttXwchzsqrv9LfL72aZwLQ5mHGLdFNQxGYA6JMB2leOyYSFsFU9ocCGV1bL
PC8PWQZbYfNvqFb1xPcU3tJbZ7fS9rY9Q73Cf9lFqfLCg5e5g0wA4sXY0RBfMlv6d5ntoBEhFXKj
KEMcYs28fidYLp2krl52QA+GGO7ZrCYWE59Z1WRB9ByzoMSOLAGd/7w0Ims9jL8hlBrVZpCJzolp
fckoGxVPs3ppg9BwToT4bU2d/5rmjypeZ2R2aiBMFekliAXpQ+NnN1XoGZN71SMI57Vqq+dvrzJp
iJjkj9DSHE67b5aNWzG7Tev0wXuZCwrtqYLEvoL2ydQzRvd29dGXiH9nklbMhsAGmNi82qUpqx4h
U4O7P+Ir6i6b3E3KuMa8IZYt0ou6tMky/7dBfys70t/1rwq2EMMmNElsV/rAr1BeOi9ZV3H1SCX5
xTukg1iE+ybmJTqalNyrfN0Idfb7hrpQhf2ph3aL38wIzOOVF63tILEwuP97NQ5qH7/5vh1irpFf
Xis7S/ax7Bk078ULZmWUN7vHQi74Gbfx/4H8X2U17chCgAx1fRDQtWgamFLGts3rN5uFIGiyOXuD
fdLCh0bSGXyMhId30RTb1UF12oo8VYqO3aVmiDjmt7V7we8jDHgYYvPPYD4vafc5FPDlMyxR1wTu
7tz7Y8aaM0ErgOpIi6FqHxi1krpMc7/5oqK5pZ3ycArEVuW3ITNtRS3IPkxAFLujnyhSAB9RTg7r
yvYvfSPhgcVNolbp5e5OYmVrIp0axPD+bTcSmvSeshJax889xkZyEbrJxgabhawlh4b/WB7AIqTK
C1qeCjAisNXwf0YXGYqKvWGChqBLNWk0yTMsVQmh6i2bHuRtmCwpIx6nsDBckZo0qrxDd0eBTOZ9
EdpeqaXUh7Iu97Gl4f3Z+ZwnV5HdNjZCe8UzhTBg+XZmTUGcGE7f17KFF21++3WMYFFjwK46wKlt
4x3/9LS7UyWJ6LEvST+Mgoi6U//17I7xuPjCrcCjmiE8gXSNjnpg405a+JPtE8LbGZkaiIU2B47e
55Cx/4yiMamYuaY+U1Aarzbj5ct/u4O3jgefEY8ulNxqbIF1Hobgj00u9QStApZUBY8JT8JVsfpk
kqddM0245euR3+qce2qJoM086+zGqpOCHGhtXzful5Shk3gO5WkMUwFGpNmMYf6b+2zJ4dAsPNd8
UWdcHFhtuHgfCvcjt0hfA6gqVa20L3BalfeSnKlYHeWmgcMJF4YyBuS+MFn+CQYk0Bp++6El5czK
2RmNfZxaOQKA/2fVpLjnMbUqM+/EZOKkNGw8TVzZii8h4bqVel0rMh/TKpGDMUwFRuwarkjxalrn
ttZlCTciCy4OBudSJQzMQ5T1wOOFglv/HmU9mk913RwLjX6v31TGlUUBFJHi1q0z9Zp6cyu9aM7D
rpdrFPR41b4YaHEguoBWbHAFi+xWm0li7C8cVI+qtcygDfEY02ZxPx/8PvjIeOzTnnMXU8BnCvPi
sGXxOWa+zW8jgAXB0zJhgO6lT0f0LfiVrRRdNHhDA0d0mlvizxK68HVsmz8C+pR55n8WujoxZenY
5WOXSUaqtVBK/eIQBoEKalssgbhaWggPWzPP476vh1hXuiS8YXMC7B5JFKlKDPWySDYqmliRJKyp
uSq6ku9Epunis7d9zwOf4ue3qnjfhvWW7/edzLAjnWwHX8HhD5pQXl6Uen3xQiU13CZKv+mVLbPY
tjqU0JMlIA+rkUHucLF9rs75VMwCLqvDPraH1lDtF4zsXmTOoBqq6AqozNIrBkiP6up7snpJox+S
A1IkDoKVe5ihKbdSLApr87PAPPHmXylqj/idrWr6TTqk9lpxy9WgRgATPUdmcZAh9J3Dqur2DfYg
Chs30dMfhE6eAT5jqF82bmiRN8Vz4KYwMSc1FZQWDQHj4LhMBe5iNpOZ8egtTm1SUHD0cRBswhGR
X+LPO8Ewi1s+7HZHQqhXnggEfT0+zS7Xz0/fVlZhXw2L1megRF5h6LpN5m70FQCsUb64agtNzRk4
hREMM4QJHrLKKV4Xpub8bCsQcVGB0XA0yTYEnpTmdaGyIqfvs1BLvDXZH70LsbNzCkmkdwcz26V1
f/HBNbKVx6TFLohjSN4kx+UNTa06tfUuKn/ToqWk1RcsfyIawavv48OyzsDmcfyf+EseawCCCus3
GvCMh3nSmQ+vavhuKwyGc6xHJqTFiZW3Z9xu+yyDhql2DloGAP5OpOO5klSV0DM4bdaxCjO0GZ/l
q1HVqGCEef0XlOQhIBF4bp/hc7Qz4t4UR5e1hzNaE3BJimAQWyX5xpQ/R5Xj4YQx2dTLpcPzvt5n
oBeC3HWKeTAV9xlt09ZRqimGvi4O2g2wFIvy0uaC74RK9wLlPETEnxcd5ctKl7wyd4CjsClY+jna
RtNecor37+1Lag7JT8qKq2tr1cx9Fusn8UN9nR4KcmnppxsVFrFFzlOZMCzOmxHE2mpeZ0TyspYl
IWWVsKT6oN0XNhWcldrMOsvKKoWtYnVzjNLd9fR1ezHt+0ARPG+9j3dAQGNCVz+3abIrkYg3JrpP
G4WbQuTN7lCX+dmiZCe3jx1vUTn0xpx9e+R9fwBs5Vtcjzv+jAYBL8w1cVsM/NtDuKBBk05R3tMV
KTvcLL5Ss9r9k67cht1aiRVzqZR6NaGNSGB1+akl0SxQ+z1JX6ql1JwPHTsYcIvBb8QRcFrxR4OB
uFRXBC27B2iwfEK4VvUx/1RFuF3xW6RVmTNQFpZbu5FFyBGyl6MTIpUnAxbvDP5MgM1fa/LrY1DW
FQ3mEelhnAywkZnlq2cyTK3rb9Vt2qVzhSTGplM1qQYc3lblgqBrWEL1OS1pZNGW/NOhDDh2Y+i/
fpEjtL4kq8H2g+w1MSFwJmOIfDogm0nDAGYMCNGTnM6Zi9fOYvzxO5jK7qc2Q2zwoRm0p2z7ScpS
ilAxL/IVFrYS6cBXypg4jveyI/NEWHmF1Wy+1M7BWfS29Zit3rwp81L7fbPloZy1tHBvlMw2Srx3
PekWRhTMaRBW+ygLPsxFv3j80AHyd4W8q7qoOTn+oe+dzKkb3+T4BzbPBkd+P5SGAhq4XrJM8rrR
tE7b15MZN5VAZbgBCx6RnsHjfXh15WrYbW1aldVROG7Qx4M21LwLoAmPEsNngVF1Icxqx8UZvmZ7
AVRQDzxQDrpwpVvhR+OiwXWPpOqq3OwrifGAlRwh9v+DS5N0wNlilMx5BcDTMLCEW8tTm7IcpKVZ
uI+BVgI11aqWO2ZkKVh9JJzBdTiPHQnyb1CF1lnK+LaqJpU2MvwFNhxwUaIRejBVu+WEVKo91PAJ
WwBMSIPPPvPFIRxDMGwLXEg4MQkL1p3Ua0k8KKssE5e7UE49SwhzGHCR7zJ4JrWFSqRyc0tnt31x
LFKmhJFnCHDM4WIYlRzY959ETFUMk3xBizp88Daw+7dbEfUxfYHmhustqxsYjvUR/yO/YaQlcGgC
BG8jXolsEG9ibhhRPaYhoPtRJppmA8cph8/CqqCLxDiJASuybSVks55tNPFgWs2KvEfbzMWLvFtc
QkWJEM7DDs6NOHLPLq3fw3cB7vzrKDZY01e+DKLzObx7t9XYfZE5jgWaWTq1vXIOnkKCtb+Kbnmu
OJ0DTfxkGh7W6POOqk0NIS/I74fR08zcS5FMMcoXXKKZTN3IQoTOZLlKGNiolV8rdkeMEcDUJsbO
0vkizuybQGXKG5nmOJ9IpLrsxMKJS7Tv8a2tSoPbVDIdrf7ziHPQKWsi8CDHN2pSBLyCKP+TnhIU
IlVjtcmWe5FmKPvl00nqDgRsf6GIvArrP/KZLr5AY5/C3IIy3oOxTDy+nJJaWklqd7oKiiw07L8t
gxxRQfdmbDjkJBV+jjYYoGW9O6Ry5oVk7lImPDV3VCBCAqaYK7PXsz+tfBCNcE31pRAuErq/lD/I
4yfmjYKHciqeXF2hQU2XGtaiqyCRhA4LU0rtsjDTeblJFZDqz5QzZGsOblvkE9xawy4uG9uSk2PF
AYGNgz5KwezgccXtGLyPPaHhJAIMjNme3dvw2aq/6rIEahAOKw1sot2qCKSNshqiPDQjcil71gLS
+1CbL8gK29WCogjcRrMEvXwkkD/+IdZYXmrt3gTZ9Q5h93yc3CxI/w7GzZaoN6pzo/4gTjcHna5v
uLr+k0UM+ezwfahNt0kNqGoN7WklZ9kxVpzazztFjBDURtAZPwFF+4biJo7boDcFTE69E9EN5y2a
ynapdRJVtuVWLm8fy3I8ggSk85m3QGg2slHRCSPv4ih5W3xUIrC7kN7F2c+7cbkUvdcwhxqnapkV
lmawRTc6vXIejTepxPr6GtWsPyw8lAN7fcKXgvD0L6hjrbdab7jm+jIIjE6C+7k9KxZsU5qVaTy/
bQBlZ5UW3PC8roQIlLHV6JKZMWG0K303vkQKlnii52N+xQVyB+xij0gR2bceJVpZ8/ilLcIky2lI
uZWpUjzTDEfD+Qmrr7B4utZO9HeuTKBWOwiYTSO7BffrcxJh19ho47nWpIj451Qh14bxhmoXTTRo
v6c32XJxEqJ99AYlEz7NYp916dogsTTocgT5GeHs1vk6aD0K39yqoYVUIr4+XhksGAfd3cPPKZRH
IiqxaVEVgHYKIJfAKTHNQQKsBKBqH4p7DjW+c9krObHN2vHyLnOvmV0fFy1sMxIV+kw7YB6TxlhR
x4lZhGeLokSuuGkdIg4+UR4Db3NCUIdGYOghUFG4W9OnltmdBqI7P4eGMq8RgtVhhvfnbUcGtMMw
hRex4VayH3zWNGZds5MEb/HimnQO5lNuUqOyX1hLS0Fkuw0dlftByuWbCcdqmmUWSPECI91hWRaL
XnXVQnQ/PxfCrTj+xKoR20n1llYVEKdedo1+yja6XqHgSeattLZb08MW/GluYFIf7Ku0V+1FHIou
Bip0OO6rLosycnuxEqy7w7gaN+SbvMZzQJvUnCHAtTmSVNb0KLCMYH+LZha8oIb6mCJg38McdVQT
30Sw2Nwqe5ksfzKu2Qj8RLZYWXr18CXJ47+FoMm9znuOoTMqq+YpKDs/rzhb70+6xRZhtfki1DFQ
IOlxF4zRc5DeboxH1kKcK9vXQHD9Rpp3YMJ6PQvFeGOM92o44G3+GF+jXc7/beWLuwDa80BMTJZc
YlXrk6BCFyQr2WOTldZvUCZC04cYe/iz9g08oqq5qMidOhuExnzMPTVtrAcfPVQOZ2AdgDI0Pj+U
aTXLxDCA9QIOtnV+kwF5Zmn1H+Cqbnc8jpPv4O30ag51aaAfLgazcRgr1O+9l5kYbsVQ6HI3LTqx
vEiDVOO1WKYSbfuW/pXGmvwSBgIc+/SR2IaH9d4IR5umO2ZGJPQcbfvrZJZTR531x0BAY/U/38zA
C3bSiRTkIi6HGg7zrU7BmxxI7DII/ItjXZWwDzQWyjHWHa8BIHGYJ8fVYpHJCAYL+sAIGJXvwRME
qqslg8os1fcOvMzPc6JVNoFyFt/HwnapvRG3XMvdAVG6qu3wy8nee41O+mupAinG4DOpPafZATB7
ENl/0JKJz4c/XrNq2ZlN3iSpwvSYtXO/ib5RVUAyYOIJuAVE5OjAuxqaLkLyq3zvvNuFTG0xNIQZ
JzMMGsVrbh2KiEfhPpvZ68oGTbWmiP6HuBxe6PmSVSu5QyHEn5+B82M8re/oONOMr7scUTMLPhVP
UuFKw4ehT6KrWK4puh1u3mKR96Ki4ETOW83B98UmbITMu5/+uk8fmPRKBrVgPdZNlCcRQ0XE2CXQ
j+QRVW560OlOXt1WwzIVKBK2Kp1Q9PDICKgIBwc39bsAH1tYDeWDnOgJU8iB1xQlsov55RiVOLI+
QPlsPNZQ6NSEXwCF3S4ICMM3F0v0MFFqRNnBeqO5BvwRXqW102I+ern3eo6kNsA4jrJ/3LRHfZta
U9g6H4fUjvtiFiGe4j8K9cvyAihWlNyzb+nkPTZftSIQEsDSHL/1ib7sP6JJnrmvmdQkTZUTci/U
kf/un8TE4wIWQRxnD+M0TKsEsbqJWk0qgLe1iPrQaoX0bhZAZmEBUqsuUkQYmaDDA/rFOqr6vUP/
jXceP45nySrIBnqUdK5Oj6ex6x4s9IMh3VWxq1acJLxT2fO1ybBufgnwKLr9vVKLenxodpbDA8pD
b3o7RFkkUYWRl+uu5ZjGbPHX0o+lmkuhlx5mkG+Difz1GkovQ/akLS5Q4ydMcPwJRjH1X9pKJQTw
uUXLO7hh3Zo3fOg9Kh3srMbkNjRvBveCvSyBDUTuVgzwn++izzvtmXvd+9K7zdULo1bTwxmcXe2D
FinEbg4DaxzRwbKsCtmcQ1vflZeDpbaE7Sc6z3L0QOwjpS4r2QaX5ySBg7UtK0fAIomB6GUbp1Wc
LLavtkNWTrgNQ1WgUk70X4fcOyXPItJ8gEx9Sy/t/OKTdPltEYDHkkzxHfl7DzSaXZbVZmEuO2Dk
/L2PDQ5tgRWdikfi01Q0W/gpcFzFjIc28BahjFQtNmrgvmFc4cqhJtIrTHm6GOmAikjwZrvnRnXp
TlX1K+3lXFcDytwPLblWWZj0GDmetUlPsQbGbyErRlGVCPnGOzu7xeGSkNwvucB+E+EBX6NsvnZk
EvQThOeD3V0xivEUFKt0aqj+AW2iQKfgRaYO+qsam23ty2f8oVauHLndlRw3WYXz/TH73AQYMbzM
u+UmmqMo15ty/VI3uQmQOtIuSeCMAB6XoEvoC7U0DnMxvycMQK2ZYuZ9/zyOZ3SudjtYWXX7XKxA
GRMij9z9WaAA8TLqcqbfO2UGe9NZJGVTIBt8Ff+e3PysQcjZhHi4cgzcAF3PlZWrJFBb7cz88HlW
z0RxTDs1PZQ1f60XkD1eK3tsbWsfULBOHgkfU3nfcGHFknEuOMS43mKB9HU1TOB/XyIAevGxzFft
rJC/ayFj83/XOb0wGvpQv5szOBuiRP1v7XSVofc4jpw4pMC4E22/yb+X3KRJeErL6WnP+KBQWZLv
rfM3Wa0qjva1P8/p3k0nFpt9988HyVfE0fU1buOuk42qLokEh5d3KRFDOfsUZwUYFJ8aIqxGgAs4
p/sV4PP7TkPeU+GNODWS0FbKgJter8zcSs35FXhxm57GgTvWe9Vly+5m2j5cOIwJrCYMY0+PrI9J
4oqmKw5RRKEMUOxYl1IqXk3NuN9SUXaCWzv6cOzbd/U/oEsMWW+tJm82svqV3w9HHLb6CHNi40Q6
WkfIrrKNWhr29xgBSUcRt0dCvJkYSpM4EOhkpbS5tFMA6I/ZqnMDaTXgBLhv8EcBDSkWn/65sgdt
XX/ijcUqCfpyO8FGR0AlS+UGwGvsMNZ+h3pUmhXSqITSQE6uzW/dDUVCHnr4t3PLM7xAGOkW0P3c
hSkZ5FBXR5Z0BQ+2oxwLhL1UDFhvdwaQbCjOavmu8q2RMKCRCA1Frm9KjmW5tcXaKFqp2PVkqaRP
oSqL5CRNPVrRyBG+OgCinQAAc5W89HnZJJ/6mP6L9YBJZUcevrFSKWkVG3MZeXL5DSAXf8BGvOif
uKgF9l2AgeSol2YsW4Znpvt57aigPDLMo6B0B7xx+ocd3w2AhdN4OCbpZfkCJJe3021FyJoLfmvQ
0A3WCUppfcgraSL2MTkxyEEgTaO8OiGO+lop1c2SipI/iIi1QP2HQ5fqFP/Sj12vbbIU/mOgL4NY
YaYMiqS5WDk1NuAWcnCxLCXNtzyKGJM3txMDCEQ3oT15SrWXlcd+gjB7RqGMZudQAisOJJQiqBda
nFaMm0nDX/bJZXIfa6Kdtk6jQNpJ3hjzohpIAkc683m+JJaQIaQs0tcj+7YxI9oUVEsU91x8FrDi
UnsA168pAlJ3n1YaSL5FYEz0tWPQpJcZ+RxqSbbMUaeiUUriDsZnCJqAqMwd5XswBV16aQXqSW+W
Z8H+wEwtTH9ZtpQFFx3YpBA2HZ9f3tOuUm1eLjTavJYJKQo5gwdbry2E9A89MTqIQzoRxV1G3tYm
YbXPMy1CXm3XBAkLl0G93tqEU+Po36u7AzJjf7BsD6Njwzss1y+JNuSs7zr2v8NbDqZ6/LI7RsGV
A2QMjh0UVhUfKSZkl3m3j2lqcgLSE8eJAV4PY2n2WftUiPDxehOjlvLV1QKOTMPQMWMYVXLTzTUA
h3nhARA/olewTILz26jzBstKOwH5iEn98fe5ETyWnZ+et0U/UluvImo6hWIKjVuc+Auil69y/EeV
eaEgavR8ol8aMz+wSeVg0YDtkqf2itrM0xicOCaP3OOq0ZsUcvjsGNLeSOk0qgQGd3JcPZ+Ppk1d
UpKpCQmdq265DTFVZHdfM3JBb3T+Q4EvVXnzDtrlXciGuxcq2N+vWMSAZURYNRNHhYXjnNi2NYlc
6axK2ARM6YmYa322rkI3L/yZnQt7FiKEYFUVewhet/0a/cGR/3GrGZ4Nbtdck1v42uf5n3t/qepg
cZlQWWuDSF1Dwx9Is4q2uWsG9aUe74dqENIJ/QI+pt4WtWFTGWsKxvkPZw/mya18TEqUnJF47ItX
89jUXMrn1j08HbIS9pQPyWPYGjQHAQhXrNM42j90RQ6PXj4I5T0BFdWA3uDDNCtvDbaKUNoEShzo
mknXBZHAPbiZzgHFkpziw4iwBrhYYbMvKoWE2By2p/NeiY4NwO9JBOozunVoyClXHYBIjVZxZku9
yvoAzwys0o4HrPLySpAlNUahX1vTv1MpUwf2V5Xc36ZZPyHq/pWqQdw/F32mZatnGvJG6W1VFSq1
qnjA5FAiT23JTcgZnjOwvus2iEoa1lF32hvME+kOoeSQqmJ66+KvssTJc0xzqLphxRujxuBki7eE
64Mxy427RfKJxONT5daM5KlXwKY5j4f/nPEIiIdCg4XIwK6/jSr8dXgISQzfhx2iHQCYlXTENjDG
/uMbRk2wCsbX23b9ObZcI/yj8ZpTAYD8Z9mUCGtGRzgNGHafxLKi7U1ysw9AhCEc/QXSuXY8FynF
O+1yml7mYsOkxpzKe8KmuTPU6RA0mM9VNek+5ysu3nJ0aN+gE+9TIj/6qRto6+whMak0YHlpvqHw
ei2HZH2C8AAtnalsJRsWy/pVHVQDWFlPXMTiZ/AjGZKN0d91zp6TYYqDb+IPsKQ4H6q3tP3huXk8
SqJjbnWgVJHuS4Nn1P+LP3VdwUcw9UrUTODpVnLKY/NRGEEgcypE8QqHzSpv/GuwZcNd0Vdv8WeB
xV9Fs4wq951qJULzV6TOFAYCMpsxkp3eMQnbb8xGL46ACJEUdVq6N5IswDgYLgXdnD2fp8cppHCE
zNo0SDx5k4ONb/9T/LB5RCtESLVU3rggyA21tTz5A5zx77LyP7TlIS1J+Vz7dPHD9oxU9tz2pCqK
ab8eTLayTSCrjaClfnF0kDZOTPmCOIDkpKu+Js+QsxpWhpIAGLGfhDoAQFGU4+Kka2qJByFH+pDF
X6RDH8BXgcEeHfUlyf+8QfWciLI26c+rCBWUZsd24DX8teDSOaf1aaPoMlGh6uOt+qWd7L/DrQsj
omO+x3DsTsC0R3LdG4DADYZa/5HtQ4F7jOeNjOFw3KuYAW360dQSpJwPy/Dp5oUVMRvmljgFkeCB
d9o0AdSx7RHUjCqpN/ps+742Y3uxWx9lm0EHWZjD/BqidxIiSZ5NMC2ZERzPE06Eh7yK8xn9h/4v
zKHvzlZBc00++bODvbDoOcE6XIG0B53+LX38NsqX4LpoBfX0C7rfpHZeyA7Y6q9We3yykOAOP95R
2MBNlC0a3TFOpxsa9bA5A+tweeNwuJrFo8ykJidSsGH8rriAOokGFrVr+tlkcEfFPw+Oupp6UKNr
DvcEpQFlQ259Z7wfj13MRK5FSZT29RQOlNSqwUsStc2kXD6Ae/NL+Ldz/gbjN0C3EZwRsT7fv6t3
gZltJ9seVvkyMz13ZdFkmcidawpfnb98eQXJNdFtP72fxbP/jXO0TFxi7qBA0YELINclflO3U9XR
p+yNlgee5HeVzE9W+T/HeAvMT4Q0fwJtfPW8N2mPyVDwgb9DTEu7xf26DJnjyg9RsNsEET0pBB4x
JBgFlcDdUBXyw6Zh0kJJTOLZ9j8sNMuVykCeWpJKN8K4uUGdkffL1QdCzOmSERPTuDXkGA0IK/zC
J28tQEqaQs+DSl2E/fC2/2bNO99bfdPMk7M2D+3FkObEGb7r5ULWcwjhSavcyJVe+aKO+aoMV1m+
Quj1c8iFOA+HoeA1WiOUTeVDDAwQ3XWcZSUuh9ydSazk/Sn1jC96vmgTqyNqJewePP2gMLLucJNe
4ajVuY5JcWeeYA1iwVXaTzDofNoXn51UB+9VAnyJz/2Iqhq6q1pyI36CZGnuV0Inn/KkDrcTr362
d1J0A+/kcUR9MZcpFRQqsWLSk6pQ7quQO3J+/vIgKnFuZ6gGEXXMlgBAZ++U/edzEShtVuHYIATD
f80N0CNpAof1rdyfxRvkZEvAvPMdVwSfC1u87vnLQ3wzASSnYgxp0TrguE3X2HiJUkrdIaXBwfIj
9jP3B4lDZssXOq16q+DtDx/YfMpCmSkGk8HFxIAfgLPNh1DQsdvEVmKLaubW6XyX9ndKDsKCsvj2
lB1vhE+RtgW0xi8tq5Xx86sQMAZXdzk7IstdukV63LKadNVi1puTPBpBBrCu57jpLNC2wfveG/53
N4ghwiyH7qCWTh4eABWAXtpufdX9++Zx97iqDK2pIdn2VFvJgGcLaL16lrNqQIeybrOExvwuNDw1
kDzOa/I9Fqv1NJEgs6C/icV9wh8Q9W/NnvcAoy5aSvpeIEge42M9g5f6RF8UZs2x2LbIPp/yFWC6
TX0Sytgs+4bVtlmE2SH5HDuerXPvMYSP9RYZHViRkmbGgJKZSpQ1lT9pWnOMs94ymOQmdQ7xTUcc
S8Y/0KqnSwy+ls7EiyGd4efaI4y1NbFFABf8BBFiJDl+JtHz00jYku7qL9wndLMzfnUuZ/if5MpT
pHkcj9NAMYl1/BGUOMWj+PIXwu2uZPGq2gj0D1F2cdmLB3iXFZ1bZv6DFNlzEpigWDgp44utIL1n
PUyLbnyUyq11HGe0t4YgptB7GhPIH+N8tsEqArUhm2OW519Ajv6lw+edNnfFkI20xlZhFfLegmrQ
K8OIeCEXU8xezUNe38lZ/URY4f/KgJprOjK+Uw82sPF4okOT9o1EKGH2G5TbTT6tnB/yBghdwb2O
GrlZXNTTeZTdtQejJGsbiVT9Hijjb023zYoIGnRBWMZg49ZTqxrqekH2XqA1pMARzhGVj7AP2Tab
i3t0w+2Xwy9JYLhrtaAk3156cxOCzDwLOG7eHmR/nenQdiTNa2nEJ9HcR6NK6ryG4V/yHfSG4t3P
1kTjbkiUI3SLLkc44FNsAd3/xieKwa/28R7TiEGYh4F97CQ7GSdTa8a7sGp3x3bFoJ3D6xtD4eht
xmg8Pa5sVGy0unDlu6ZVTZBUzgF4bVcTQz/2RQmOQNlrWITPQJHD0pZXcDqvGsUZCpe44gKTguu2
lJtL5IydfcPBDzA+b39E9YUb7W4L9ErFbWps/eQpq0Tv2PKLHr1ezBTUA9b0f6DHwpItwMWr/zWL
KcW9aUn/6a9gaEFo4piPzRigs8q3dRz0+BgtTq4qAFs7jJ07+nYndAEfmyQGsn2AoKu6avyL3trs
Jhes+E2sewbUlrebCzepU7vyG8o7xrSOKlRKeG2IGuTar6T8a5o3i5FXVMQR1lSztVK4/GKx0oYg
wF4dxkBbIn3CbeQj5ZQ8R1keYFekmJcMowk/7o8a1/cCmc6YpEnoRPu3ke7siFIKVwxY+HWIXHb0
mw5CJak9TnDU2dTaFiOqv64jSeVAUZkX+vvziJj4DzokdGD/q9Uyc49CAJF42MiY65wwEEd2lc82
vEBjzlUSghaYkYGNm5LhArEh2xCUxl/Ru58tZCFx+m8/g0Oo9Q6AUknyQ/dln4tX+ieoS0VvNTlG
INe62aXX2WdMEaSDd8BrHRih7Oq4oJFTmkFzXF/DdJO4v8NPTCo1urBfYLkY6Xy1jJnNCdIeirMo
jz7B41R20yYr6qIYDRGQRPzVLydHqGIJqPEjl+pc+3rg+Qwag6sPI4FLYBpjbYx+OhbhLL+ZzuAW
HqTX0GvL0eAbc0d4coXf5pBvKsg9dJop8M3CAdRuaxVLoHwGgwCPCYLI51XgxQ4scoA0xO+lQhEW
rzFytc+NVNbdzc8tpSQdF2VlwJyv6hYmzFfJBl1nDQuxiSG2rKtjh3vyVhQEA98p2qQDB+/51y9G
X+tFPYMrZIne+9VhX/P6SLzFdG/ds0+GIAUZmwJA1yvR5wMk5zfJoHzD5wXZdWFo0Bf6wP4DDHLR
bCYqilBf4xkp9guX1OqzNfN/O2urCI2jIpBVk1uxfpmAZzgCek3Wmav+kDDPZhvb9D8ATd4Sq/EE
UAGQwcNG/JQbCCkEPtxSzIsfcqc/MOgqzmYf6F2Jcsk/UclGr64vmHrqNoSidjNUpxUjw+46vEB4
6aK4WNkxbuixBuR/l320ro+03FBeK9ZMI29yLkBPeZCgnQHTIWq4HQIzZl/oAPRPHxXmECkgopLo
bwpmYkIP9dvBLt4HPGYCN0tdIMkxcJZoZCyJ6ITw5I7JT/xUD/C8h9HpeqxPiKD0MrkkfmlzTTFP
YcWx8RQseHRdi9qYZperzCa/8SquqxV3rwUbk7rNm1OSqrdPWc7e4z8qjZnZtyDr120N+iRcMj0q
JGK8vdZimCrdNlcrRjIFIPuv8N9ehe/wspoAl2lzs/JtdOoqC4AUnHeRcZO4XzTrIdkNg3EVA7Iz
RSo2dD2O5ALDTNZvr146oW7L68YCrBHm9Uea7MYdnd8tTwzMELpjmL+Ltr5inibL6GMSUOpvlv62
55mmzjsFYLWw2CjZePKqdDIoQVA45ntKWSx0f20ac4Hat00HG0AFKtxKCLQyBgVZZeCk/sXFHxd0
cQC4CFmRknYjU2VyTRPhArrmVnrJQfktdXXQ6zNZkkLUixIZ1HVr4QaqJ9MfIwamM6gFv5M/0qjc
xu0pWlUccpXKxSG+B3SavqfmSlMsM7ngO6vO0Nj7IEJSxkbegePNRgpnz/LkOtQbNLUIISr7dXsb
WeokKtA4XflX+eqcRfnTs7ydtn6/beQF3LlVQIz0Lty+Fj52367EAS+VFla5U+9ygPGO08sH4xqo
Kx/bUmwi6+dDY3z5dgiJxo0/KzUE2gIE1HE2J/XK+zJbJOmvxRuPZ5PrpajfHggPv7SUFIvB6p7K
C5jVgYWf2stO7cJC+3I+M+79Li5EfiB8xig45aS/J/aAiWapeJUasOy/O8oGk9WfEw5DttgZOuNc
FEDevIkeFSzIElaLvQ3qSNJ5gpjsEKurkN482T4cBD3LkZ4uHoqsihBfheAeyhkcrLug3yyk2D7k
mY50pBaBG1fShqRVKBr587smv1SMlVgL1fisB37K1vQqGT1kqY2v5RfGq0UnOswCayVqoZCcYduL
yRROA8jzkBJqLf4ANQlp7Oi9i2b1oGvK4PrR03jhvnOclQdzzvD00Zo5LD78P38Ou7CaG70eXbtx
QYX5bLTHgoarhE5pQ5k07EZmYpwEi48FPrK8FoA+C7UocFju+WXcVlVlUohrEDA6N0e5cGayfcYh
nYQu4mdmSwgIgsqOwhiIjbzqA1lCTDf7fdmx3/fsT0yrMoCiG6FozumjW6Mg9HiLOJ+da18KShcJ
XZ3MmIZ+JbDaYw+TwJwrsroi/Ykzq9q1uE1x7doDPc3xDeFKaQfHTFIgSpGLqtMOxFLBOYtbuK20
kgKWOa07Z2uNmGdhaBN+b5q+SjLdSGePCy5688nuUOxXVQ1zUnvPs/lvsla49z/SrgXPinzgEuO5
5zHuksF0j8/noKqNtz4bLaZwtPwa8r8z+fQgVoP+dKI0FF6Sng3UQxZ989eE7SSyyUnxt9ShUgvm
gRSCcW7/L6UIyx45aVXhJk/cmbV9bcCPdHjcRiGW6UwGk+ng5kxjEwKLGcufA8JcwiGdmkUSdi+d
XuYDAK7P98AHB9o4l0VIZomxqEly87In2LfncL927t6ituLKwj3GuZeE1SjN3eIJUHnqJJVv2leQ
SZFdT+altjLL8NliH8Hw9vMfh3/pnHlw1y+SxjfSLzE+w4V35dxLJn5FiEuclnxMZRax1lmTyy3o
Za8uJZtpdy7F6SsKYvm30QbCz4U8Wb1Ke2jNJ7toSxajQBCZkOKJK/OGMUjHxyGP4Q5gtHaKmyq0
cO7j+425YGf2/rP6oRQVIqIiJURR0ee49WkqhCMxC3YEOh2rHxs3gSGv2IVH1zaeMry/aYYPdjoH
r+bmgBdjl90Agv+dn3rOR7qTZMVVYlAKIgI78lJ30Vnx+MFpYItbhpB1H8QwASJUMny+DqZu0liN
HvzVBDhSfqq+f4pm5nPT3wNZl4rHbWKYhBJ/N0JlqV1EHrdGfQT1G+uYBkmuUh6lX9UAwWGuXa4N
jqynl9e4eBvKIEzECtB+qvmAL91PdkUJDQ5+3v2g7pCYamOgYmLN9fWrGyNBnuZqASGi3yLtLROa
axT3sXZi+EBhgVptZ5u1tO0yurTMOncRVDZBjq7KS1MZgZEP/yRVFqEvou1ARO5VdDkeatqpt6jG
Pgdza4sQz1kTMPRBEtj4OLWNkdBRI1Bxr1jNaXtmm/3gJUezz7e5O0z38rvnkkWiC9m72V9Db6w0
cew5OogxTQDgkJcHFCOmL65KbwFnqr3iRpo6Y4Z4k29LqY4//Htb+kLwLr85IxtIUutgJLW7btZO
wbZHH5cnRltjbqsmdXUaEtRaAEQgZWdy0+KtSXzPDt+mpMOuYeIFWz+CHbgvA/KwKB2n8JCfLM72
vfg/W8TSDPveWpI4hFW6HV5xaEYPdrh8FxEsLBTI7cBMdnLtYS5nHT5k34GmSMpz1o8w9hz2zJ//
qaFjIu8uvcSBuHt8+R2dwhS1SJeNhqSOHt2oaHdtPxCxhvbEj/4QvDfipHWpsIClnABoxccc0Hvf
ChaKVOA7G4BL1umnzQnjypC6veSR90IdN8p0JvwE4pqv1H8u/cbD0CALJFzabDyAR5zS7O2h6wZh
A3XC0blphZUqDnH2MCriVXprO/jo+U/ZgthBk1eJnZVQiyPhbdKD5e0SSEZgOOA9olDtr+n/pzKQ
u6SjKDEzukH0N0EFGs+SwHrLlwZH+jWECyG7QxSLZVBPzOg3a+4F2B3CqSpUzZSlTg7bIzqWphHh
ix2vsIBpPnEajSGcMECQ7d2OvnECMszMn+MqGd+CnG0MY0sbJiRLrxYYgfCqpas3lx52tg6ozv86
DuATjrr2LH0xbEOvjfljWdqGtsOiWajnJoP2H5JVJgUMrZgLtFCwMorJr1edZl7miuxN2Tkk8Jn/
n8OW91+4Ie4avLsh3qA/J3kU6+ALEamjq0qJoVS5sqmnycicIkNdtDIGp2QjWyMh2UW3/HmfG7Fn
zpZo9ja42oH3iozferyh28PFmD/i2tRaWlPYvddxxg+cspWKtjIOXAFsU6UFpHJOi9h1U0dSIT0u
gJYbgFomDu6MJTXKCGufrhtJk+EYD/M5/Yx79613MiBJ+sCMJp4aCQ8jnESxP8sU1CfWXGRVd/ex
+HcnSbGAhcv3Rku/pBPJP9jEHmJa0caHymR+TJi6HSy9Voe2TwbW4gQM5aCoJ7YBd++DR0Jloc3k
HunKYFjUgBaIcVxL4HbYsCujizAbB7WhFnc/sfp19C7FnJTkp2rhbxQH5l9Xd48pwvJnbuQjop8k
1/G6KgTsxmIFmurLQYdFLsrif5RfR8Ey0p7ghLP+QlNbtX+J9quwTCn/lCVWfqRTDF+kvyYEGEmL
aDxpMkf78545mRpxQINW9S3cTSzovwSjNVpSEG7bEBIIdWQijxtqeiRpKd1T/vKTg0h5qWdTykSm
FycKOyNaFqoO1+UJWDqFq2fpL8SNQ9FsSppjUmNp7aI0KRg0+FtR+RdqGvJGjKGJczPZHjIisWcV
5BEJaoEk9NI++i9Zc7YeJueXdVk+HM1CTrArRJUS1YCRRX2BJFsZdJ0qdFPYUPLv1kEl+2K26S+g
2k0a3vdJ2oZq0ZP0BDMAIDYI3mNGhuqfmBqqz1EAKg1ToEN93z2/5XDAF7qeAqb+CCwDAgdDPgHW
5csbDJzPF5pZibUYi1PgFxBX2T3yM6YswGqlceT4cSSFpIlRilaNr1Tjl/DFmXMX6nMSbUOmPpt7
msWGDXHCC3kN6piwK9QXmhSN99QXFOBl7YLF0uc4fXxttAC/0UXPWk60K3ErtX/0FaiMh2NBxL/2
grq1BbwluCc6WSS6N8nmvmDotdZhzcghuI/+yCaN56Cl8zaywPzZ3igWzemEZ2f6g1YJ5OJCetgS
0AogcBiw5YK/tW9q3ZRfMi9eEj18orkDrBG5i31C1VMCqGWnXLIGMbuZCRQe5XSVgOIFiBird+ge
/Q3cP2GjLtNC4YHzXwnxs+dnQ25Y0ryH4xhQefxlUhjsaCJZPR7dtbPL03gcwiwPGPo9PgWzkMPa
E+v3TsDnwEW4FC4IvDIFpuuDjV1FslY+FkS9x5h7FV4GNEQxoJIyWiM5ENtbOx10vp9ikDjXm45P
4lXoEgb6BGrSU6ROQzOVEGaGycxbVNg894zh8gvhG75qlv/tuL1Tvmeos/RhRTxGqTLb58i+1Nah
iK/QvPbkp+8tlg81ZZppaVSQfj/r38NhR/RzRTVAVkYI6GZNG6B//eVWyoK6KdCnFnAZKh+SVSft
yDKRKVZdOrC/NHVpvt6WHHxyjntdUBwH/161B1Vbr7vfiLGyxcU+YnN8/0LzOsx7Uj4tIZ1O7JFV
LiBHVxrWPT4up4Fe3V3JDN+zj3l307fs3jEPyvknnEhBiO2kGCtrI9P3krlJga8twOGmFhOfJgeA
NMCnNeq7l+6qpL9U1+Ga4XrZyXEuCZbu7smxPAo+Wmto+IA9OxfgPE74eKBBwDWXJrf+er/2v51W
CZ2h1TJSktMxvHwcQylTwmInEtdEA2iYSduz5wgcGrVtckMApSHoe9hMDuBo2FDGcKbny/i7rkOP
OGRcl0IKkwukOYezi/eiYH5KrPLZIJ3DJNWM1Nnnd3MCHioCfkGeUBKWG3Z227ujX1ZMP6Nia4Q2
4SBR5gDvJSaAEvdbQa4fvRCLA4954ATsGzjc3ZSAOASjtuO5SHYbkDJQLlP5WX+hhBv5rj1icmDk
uWx7Pt4DT88Mq1fBp9VzFLp3Nj26BMA7ojZXwQr/F6uEaDwbOXrX9z2IvvjuMB9GpfkYdHuN+Exo
FKawZ+c4sxuqnaOPkK0Jyv4kgIfKbK8W5iwoSD/rBjBE6af+ZtFlj5fWZtSrfIg1n24d8WmoMNCJ
cT9G5mogCR/rc+tR+PfrwfmksvD99qh4NJI84PmNDUHrBqPYeN2iWJysFAw5IaDjnYzfQQGMEMj5
IHXQMrSPUMT8vbYOXlAm+skBkeofUaR6a/PeuPP8LB8vWhrIpl2IvVrBGSfEgAXsKDbwNWBjbS7G
Njl6nhzkTmWmzBqP30uR+SMHj/W9APrZjRuabUnpqW5IevcvU6PyRhsxWDcBxQPHUw3y2BmNxS8K
3PyxFnmgFetfFgSVaBOfI5aYdvAiq5eWiWJrHzFaEhHrqmcb96z3w/zUqoDO/30+pJTvUnv1Gz2s
njvdpImQwZgpYvgJmu3z5HC2UFQcM4vp2TsHWbn1yzIsAYVG31CmBXVwTn6JNXp9b9HnHxjL+gr4
8dW3aoUc64r0Uw5OuFNdz7zdI9IbBuZtUW+SHEJY3/flg9psVuQQSjeZo2QQdOc52ADfSeSOxS+0
8bbDjgXbtI5AmaDf7ss5No+qUkSekVxjjEnB4jtbgrdMmz5v0rU/fFS+KFNzG/KUXbkfvMTh7uZM
BWtr3XaxF0QN1cqOVG8ALorJfEqAmXg6c7AYOOKWXJ+A/x7+tNaVwc9RxxsYVBYSioqNfX9GiJu4
epJ45VN0zAvUDoyyZCQTE1F+UDA8bwDRMZUF4qSd5OGEbai1TO2JYOUcZocQQepN3Ggs3kmzzEcr
OqJanMHija3paNI5yxW5rRKDCUSvV+Ym50ycS9UIN5+rGA8GlIermBj3UBp4k93kNJ57tyWdWrF/
a1nsx0FAgKU/OJ/rNmodFKem7Q1rK97wze3n1jl+/cMVuXwcgyn/l1MW+nG1Jp+oOw9yz7rO+5KK
WW4WdzuvFFYZBnfQMALsJRK0j8gQYbpGTPrFcCLmSb4C2CJFG+8VT572GFxPw4bfmCopWMaOgVb7
WAc8Mqugtk1RkneCtFxRf29HWjPQsP0+LdyaKQvMHp/oKhIASFwi9A59DYqXGJf7qxoZDasqUCX/
HC8E3LIdccdRTOIUtcD6bJGtYHJ/A4+oO3moAu25MJGzTOYSbCEAErnDR7nOeCtvYeRTytSrugHL
ZD5QZBsTCdoZ6q4tg8pzNPUSiwFljkAYTGfoEETOzXGTaBRomd73o3wleOG/caPPys6vdZoNFkqV
KdmKIKIRN43YqXWKdt+xhltrnlNjDMQMQ0QtgyBBrAnx5X0g5des4PkQ7Y4XIEZuyCb+MI5Vp7Yh
C6edQca21CF8jNxk6k2HiQFUrzHFGc9VUbhV4bB1502zjkl5xXpddvX7J5IYZCMF3SYJSXK95wHz
TuQWCYWMQfiotmJQQpdie3uBmNP0Ea2Az/eXNTcpVYMqCHL7mhm6qf0Qm58Qrr7YlPCowijhChHx
G8Cg5ddO5XwlnaM+uAbejvtTYP7TBAKtXn8JdfR2QX9XyIV08v2KlmM75YCZPIAUEsmsVch2Bd76
tpHsH20C1TBmofoxeVpGmhVzzlPQfcQYtfKCaBnHL+XU1EMRt+NJmQwSnQGZCwfR06MrkXGYwpy/
yhBEZDRwrgiGCMwgh61g9eiv3Pq2BvorAjsmbes0+WaFTad+idj6K3E/e4DwTqAc5sDj0j6AKME6
/9rdeRqR0pmfalHQJ+PfmQu8lAkQi5G5aMsHhnyCwrkxo8cp6MFLMniCHCcOSsft6Z9ew+MEW1lR
Po5wbcGjvVFzBBf3pbvy+tzcRcEvpFu6T+1Ed/El/cOH7oOQIeFWJ3xGZZ6AcE011c2de0xUQrFV
yeg7EioVDlJ7KDdpci7GWN1roqFUJu9rgwyF1AIJEy8FynDiEwrLd0ewlGMU1dfeduLiOzom4qyX
I+MUU4LXW9KgYe0Vppw7Hj4scZE4xzqlAoBtcScQ0fR7K247JUy8QxoQImMaRAvJ3E6l2+qU0F/h
2dUyGyYmyxbMklr494mGYjGmoADzd3n+OWuyYtQA0mEdkPaxuhCQsFeAmwSMaRG5M9DL8y4Zsx6F
cSP8s71btxdFal6D6Sk2X6kZn3TiilR3vZu5pELI3R/7DgBbteJ3oKYQq4mcv/T3CiwN93WbK+6+
aQU5r0pxhIdKMo8LuP4lqFB9JwQXyZwm6ke6+bJKNajO6jsXF9Q81KbZR94DWcxX3kkxmdZLUnbg
cVjwHKImIc9rH7F0PPws15Yp94w+eOaIV/b4wQuqTFO0mL80d23YcEk2zZSphcqufffGZn+oTRtE
nHe1PWZeI/gMmITXIMGstP2/N7HTgOFQtKl20WYRGqxCA9Lmt1d0Isq0aehLxdwpe9k/Lnyh2VFZ
44fLYyMnFIeqq/WgvX9ZCAZID4qPsKtNbytSnCR9iBeAmcdLbam/yAkrUYSlEaWmqiaFWPpNzePx
9HUkxHDtPbr5J+TODk84qnCdsue7iqJo64sOszWNTVXsmf3x/0xaWRsfyJGGHDSPeGRkbRmnhO7e
HcMf1HMxLq0c83aF3iq1sjFvufDJi1oX5qBTz1MkxPyz0/mcMW6cNWeo4zL125KHpd+damr2RXy1
AJVNVnHV0nhXuNngdcpSMkWrpkVMjOygztw0dQyjb4vjDVhxpg+oNBlNQ0Q4YeQPHaq9wVPnpHlh
pSkbnkuPxZ1G44U4KAo0QTHhI7TR0w3n3E5KRVimXz9mysbc9ek2fRSYXarh7m3uYGI8/vqk3RVt
nCwc7aU6fy+LdG2LZ4Mq5g9QY5HhTHB48JOCGM/g/Fx/v46RYc3YSBcE50jejkihQjqbJJazY/+S
pfyj3YrrAL8qd7lEAUz8hIzZFmfKrW9GSbrPw1jLErPy1qhNbJZ3JxXZ9hmdxOhK71phfp3XwmE/
bVf8nXjpG6G8pUfXrYSbcsjuV0eo6vucaIHzFTUWZvgSJbupuBUSMdN1GMGLMVBgcFBtjhLGJfPh
5pZTRm5kToUMV1scUREX+PLH3TQo4uyDs96pRBUNKPsZJAq32IIxARSxD2+VirKyaicXflhIGPbb
D1GEg93AkgLNWX/zOcUiWgFc0VEX0ih85V6rseHIJaAjWTyl49cujcqCG/TVCqq+TLXVkdo9NGu4
wShf12mXkiKEHykkcgAcg3k0z26ZLpv7eyqyV2LPDg/Q5O8jeKklTMxEQxOmQtIAhy2ijbFGXorE
4m6laJq/hY2VV2AcmdMu5E+kQ5O3JRjeBqWxaHjiHDRLADBV89hAS3wXR7Uvor/4bfyCnaC62zbb
CIQEDvEB80KIBZx/pUA1OQB4q/c2mdkXwnXq5rtGJIwkhefIix8Yx1ZfB9Vj17SI0Iof94wU3ENX
y0CQrQH0wq7/Giq0zbrIv8HQdW68Kd4NqLuiel8K7K60+D0vjTi7sT4FKPfwvLVg87ya1XlJ3Cy7
IxZWI5DFB4U+G2x4aADDdIjOxboBGLdx/LikiqtQl4EztbTrN8W0IrLAna/wNNRReHrjoumtO5/H
fT0hCy4FHvO/rDl/uGQNzZvwDBJSOWOYYEpU4KBRpGVlRxvs7g4u8ajSlzvy5vr1Mr/ZLhQNecOW
prgIozw2bJMJ0WZmP050FyH4+v0djgckZS1o/uuyxVlOlx4peFFhc2oNGaNP0bSdHYAXVChz0S1Z
aMI++/Lus4SQhZvqIwg4UatO5QmxvviQKOOYYwXimMXOF+QnPWA+FpnFmZcxvovGTpIi+lepvQYH
oIqsDEEx+Il1V5TPacvLKKZDfpJqV1zWHeejUg8a0EkIRsmlk7InTx9c3X0EAMUHMlvIItftUCSH
6R05Hf4txyIbb9zP46miALguOBrmnEFgaO4IgS1BQtKqbfTRruEyrkoAZC0GqlNV3YcRrbd/uSZm
sNqsHEWb++r1nleYlc0v+GI2487eS1m3dr92rQ5erBGwG/nrc6rYF8nMN4DARx1eNf73kj1B7xIe
lyb96M3AFzGr3uyI7ZB8MWczUNT3jNSydcXAviUnMeRtKf9C0U0C+c8S3NbUqOgIPmaCn7C/q+CW
+3AZj4WA9OuuycpvEE0y6pnjuVGgXKHPowYHSjlzJr438J0SocuY7VVqBc34D8jpotgeRqt0K5X6
1aFfv2GYzxGnXx0JCPCJhQDwwtqwvMd1dIi4iUDZgi5ZdpZPxGHrPSnxCJRYChoWEDQ+nHnxC+SG
LM5WDxeqeE7pgH3gi8WbMRPrEpXcfXcKT4WqwjcJJ0t1H5/ZeYpqYj4rxvTYDdGUaKOaNjdejOFf
ZUYipPvfdlku4oY/NGSxLpLGQUgxA3hBJC3rmikbr4cOfrgUti+NaNqU2R2PM89yGcclsMLoSzfr
HuxTHiUfkKK2cL/A2XgIsb2cRR42P28V123+NYf58JxvrgiYPMgy7sdaqCYx/u1CEcVTZM6VOL8n
PxkJP5ojxJbZb1PXSBTarOFw6JWdGp5SgbnjbdbjBvWkRZ5LZnRWhmoWrFooyyqgYx+BOeX14Zcr
Xkx5aISojDJBb4mrXbyG0ziIrc/F98lwHyRVT/SyPkRftQ7sjrnGcXVFLbJgNgX5EExPLnmEdTGD
4BdQ2qXN7BmtOAiz9Ct60Kcqh/PqPXFyKeMtUP7a0kj5KlEIwckz7gGhm+SdF/QiQdljOWLi8gNG
cgrwWLUyIK8Jx8sALD0eUD/sC0R6hNsDfXFiUaaXNOMeyILLY7MNZCjafvgPhjuEi/1I/DLHz2+V
MEqyl71SBPXt/HfgQQYblAjfPH2OZAX59L/tkh/invjRqSODRQY8qz7sYgNtmpJWmbKIgKoFafMN
PHZihrN5wXcplKayVYy1a1n/1jPw9T48P43wv14yhMSUBfvqBDSHysVM9Ot1Nbr621eoDVcyGbYk
XoiTHewGgFOfb2v36ATg7go4RY8jjrdAQglYV38MReUDL+2/8tungqXC+mr+QEQ0D67SLwEZYblT
KlqKG0R3u2EX2cHJq/SYSTZFLHZw5H4dmrryGm8uIR11D9tiz5HPfkdff2PxYrk9c4xWkauMXG6T
MkXYkk+x6vPbjhdpR++U2cs4R1HyGDclrufhtXt6+cigARogPOfT2TgU5NTqakffVv5JsGxRC/7E
hFmivR6VHWtzeCtw77cC7Ar83EsAUvdy2H7fQdNnVDZeOtB8HrpZQIR08Kr0dUNyUB6tJ5tew440
j0RkMMr3eVaaL8N54Y2Jw+mSWxV4x0Qe/Kz9gKlBRsM0pPLiNgZ+ziea72PHey4iV8khJuCiEOLe
JlQ5eMwe2t3ONFEgaMaXI+UeLBxvaF5HO7ZPNYFAdFTZsZb5NXS32tc+QCBn9lSAW+Ngn1H+B99L
FfZ8NoBqIgGoqJnZdtR4bP8TziVNKEMqSnsjCGHC/m1n4RNUONeKaVQLYe6j5zlFVGqZdnZAVqLh
AfHksPkVxB8CWynwPupov81cGQysqWmJ/wooHVWcIMNTfjMLurZhQ+OCt+ZprbOZQcqA2NOqI2vY
isw/nTbcoBUpUPSQDFpbHJYozXYdXpwFy/lkyJZ2O0a5g3ufL/WLX0E3/wGeFYBwMuccc2y/nzrm
mzYsDkJ+bYrruEBRwE+j+dghCqV4t0hAdANtA1YsEcnpsAqPSniTXO8LfkLt5LhI6zZuQRPyQP67
8ogGYLIW9SsAzbk2/sISp9o6AZvUibgY4OnYZ3BusDYIkcpVdyBeQEsYbqaGvFYeIhUgt1KSJskA
Zju5b/r7hiPv6ERTXCHcQ7pJkww5SapF6ytV22WVE2hJ0Xm9dBMn5H2Lc3puh0legHBKljba1kgW
2S1JSC0UTCx1QiGhgWRV7/Yl5PWdzfwGFzDbnVr58tEl0KTSv1c+4SkwI9Krsr+OwKa7g1QK2S6U
HLbgeCAYIZ6kkIBExcmsAVZooyWhoqlsAcd0KN6jwQxGBJLkNiztSygrr8KNu2Jt/3olH8wSNxjE
P7pqg8A6R3niiK1nG8M1/NCEfGNN4+Fw0dWxORuPiE2X+sS6ZHBJxbyBFTTjNGwL/3KYMXk0SS6i
mmKCICl00KLGiTDrPPTNzU9581YF662BuDEoQVyPasb78ayaLllppFPo0oUWPePKgjOOfqtCskaS
2tjVM0eqcTFgoEl2ZFb9FuFLsG3ieDafkPzGrPrnCCQdMZgyyisY3P7jLWHWzyNDU7h3KHxcFXMB
Oi/FyxR6W8kvnY7pAfR8O0MwAMpWfCGfnf7rsbdUvsNnUoD6LidIT/BvAI9Gap9f7ezLFRXrMDj2
vC7JuxtDAn+l12nxl+pLcqsTQLGLiAvYdRb16FLTtQ0Aa01DL6BGeeucd4JVTKXNZSg63K3hjcSi
KP7/1TSqdUQ8CMpC12n+64Wule2x5BIFeGBgQ8OcExMm7vskvy5JVwpzqR7BlvP3HsemGm7adIy3
zCNe4tqphyj8uXDkuGClfBZQxRtbeE5R259xqRgyGMsDj4Bf92NxT0pF/IPQco8K4GYPFNgio+tO
nWrePO7ShxOjCUW/Bs/lxElQxpQMrSZPpPgG4Hf/ae0F0ZVfjhAJ1nH9EMYwexHg1zi1FCFXmA5f
Q21uQe10necNM4Joe9eQtR9u73gwy0UDDskl3v48ajRsmc81m/sHm32t3ZdMUlfQmczfPk/kbGqr
RsYUw/RDeew7o7Cl3BXLRqJFMDyAxGfBxHCKM2FZ/OhfD5Ixm33BKUqHl5O1wH6h8YbkqtHNanIf
UoPaEQiFp1MsV6xQ+53OZ9eRFpWxkbDZe0O1qov6NTGcTOLX04Mynsw3WyHZ6ns+MTn4AwPV7HDS
a1Q7nKj0PDoEsBUvhqx0w0fy4xa3gpo/FrMM40A2vI23ef+Wy+pMeXIs1iBAGalGUcDwI2z9KyZq
zUK0WXWh2Yw1p6MopTFD/0X82eSv1OcDb4BVzEr80/Pz5dfTrvkjXdbeTPPaecOIFWWreAmXXWtm
oN6CrHQxaOwWhNgtsD3UUIyKrGlXBlq2Gn0O8v3U0tJ6IkI6Dm52MxS1x49txzPUGBGt0Xb54jGn
1MEOb3UKqW5rRLF7hbp813jU4t61GZgfRzVoRIJSneiqd6LA3DepQHqYlTet5qdXpD9jxUsNE/tY
vsJCwgzspLigE/pUvPOC8066hb5Ix5f+N4HYrzVMmJs4W2JS6FieXiLagTDGAhk2Uh2tW8wqyv7A
/uTrZYr/MFMaQXpZVe0f8o8sJN1J42qPVsRdLKS0H9LlvxNSqeMPmEP9CblAk4RKxdvnLvjtmyul
yyHqtro8NPYuSRVtcHoZ5rQu/6PKQilBffphDhauwJuSJd2MyRiJI4FE5BRn4yb35DfovIiGE9LI
mpNBqvsI//mu9h0GsvX8Z9J2SaYQQaj/HfK4+q6Jpn+Gi0t/WKUsa71MRjBFZXQVQsV3XDmxDo5I
T+JhOULQRzYbR9trWghVDwC/OHFQUN5QucOLNm27s3pThjCapSLquoaqaUHGFhqv3qOW6cHsivvm
QwcdazfpkJkbkHSUok95wm5y3ikOr//8DfLsb16mCJFFUtUVMwK5PPNTB+y5PrBtbtUYpLOCZq73
RlEiJGdp7hb1OBd9BniwKMY2olhQduU2RqyKzPBfoIGQO7A5M5wAlMcza65QOkwdBZuQpILmSrkH
lNRgMMlWORRrm6Foof1+6qI5n42vP8PDrUPyCxmE86idTQl9PecgWD+ZDXtUJxhjWgf/3v+mMG8e
XwYudhkue/UOBGsKc6tPW5XU2FT7PUWPJN6CfaA3ZxYhVodQLdWcE4bH2IvIGAWPRWkKAK9Ve4JD
+eoenTSGmXV3rahEmwqs8K3ESpzTg4XOgJCuOv/2FuETUZiqWj6RjC5eHE9icKuHjk1Zu89MEvQa
BdEGp4AAsH7MmWDynnQqOZmBIE7u9NAtqf4OcCTbswYis2geCjP6Ze7Nonr7eblumDfJGHfbJpPa
ZwnHs2MnrTv/OW8kMwm994N5n8w3vm4Jq7xFEqZ9YS+w6lLWh9kQrbJYbK87IH+UMcoihsvoWiJR
Kj0O1Ggj5EUwVLWuRE4yGZsJfGDgd4Gu3SHHz8jrdrrfLiqooQcN+hKBv3vqLH3JyRld445Hdw7a
v175oe5fZPzWomKARNEJ6aqF4/5HohWFaUiZjNneL8j9L/fiZuXDQt3ase0uHbVf3Ssyi51RlMqU
o9IUWpBm/osGqzuMbLq4MIZWUM/IMA+N7Q982/OAl/QlwoecpzJcIcZvUGwNNCfZBbVwhbk0wyx7
15Au0aJHUB7tI3NhopkdwrjHpYXZXGz3JIpTSV2bSoeR17TO+VkVvXjCD+dDT2NYjM9q4vG/IwK9
tTbDdtqm2Panuw41Vl5J58kg2h7W2FWUOUF1TVMA98F4ZSWm4/WV0JZ+B3wvaCKnSf1V+NxAwO2A
zo42z9707j9ED90QMOonw23qYmsVX5guf61pzkFfv1CPZYpae1lPzbv6Vdl7utAIitMupBfzOVIC
EO1FXawCLJBY0532H70NTHSiY+tbCRusxPVsA2/dKYgAT05a7niypYVhiizJqKCrMTYZZotG/u+8
DwTWE0xHdpgweEDe+lpUL5cOXqEtjURYC4qfNHNP5GZNegDfT/W+0aRS44zGMS7qGS3+wQK8gQ6e
S0Ot/YE6Re2ZevVseJUH8u/xBXdHwgQE2NFNuCNrScSj4zkthDNxl/28nw59iYezjKK/GjLccWze
9egW3RG9azV2c6tTuq2ZZYjxpmbxgBLwIcGp6demhUpyEn3fa1G7+lBfZ+oQxlsXkMymIs4vqAXy
cqGxAnSfN9uRSASklZI9mhTgDEuEcCVTnb1EthuT93QxZ/GhzzJmq029uzRc64uDayLc54q/D7gk
3vByzYJU+pn5347i3IASyjV/C05i7HO9dthzgtd9fhBcp09xXhCp7Qm0SOl+A5rXiI8ZESVlti5G
braDUdTuTynYtN3uj7U3Y257pK3OUaxwjJ1zPWsU066lLgsO3oV5ptq2yn7npzAYwBcGqhjWctSN
1sXznAkbV4V3DaRKk/OkGZrJ8UgiuY8hmB1l1jSterDwwlHqM1LAmbt+B6EapTT5/8SXqNBh2wiC
t0qq3doNJ7yXUBESQaS+E4RkYbjZdy/An6+zkL5nIEXBmSBc4ManaU8xWNK5dTmPR2Fqwhla4m3H
nng79PshBLHBcLpwB7sth2XqArBopOFVv5RgtQIZm7vkkR27aWb9RMJgPcXjTtJh1wONhbHcPu+s
9TibfJ4z3jsJazbgO4/vzCI8d23NbRZzghNBPP1TDhYmv9LUtN9+2C34Bgt7irI7Wh2FYehrqth4
mReqNqkMmmbsnRCfkxVL+cjYzbkTpsTjok3KsSgCSGj7vnT02uhBsnYr7Ugaw/yiAsK02FSUlYtQ
Sgv2U2icqpkbkuYlJPgVFnDcvcbIo3FddaIZS94F8Nj8pSGNuRMsesRecSwFPwVCQrhGzMxHECFj
IMgNxuwqAEphYQOL/SAs/zfTdjJ9T1xPdnqiFUuFyM9BcHLHOOf+rvrUlox+swDmvBLhkkxAzL6x
yrxclPjN0y4PTAQmMmOTCj8y02pd4kWii3kfAS9CdaIQLdqz7gwODOsUb8LnpJ//iJRnPNgGrvaT
G7cy0KDYtxakWvutjGReciUFM9pidFTXs9XUK35njWT/bBeOSnlXNP+UQBmqxFtAa4qzG8vqbNdT
4w4ZqEsECMhlSE4cYiiJTj/pmTYrUbzFOl4M16Vli+ndBDnfIvp3tM36eZ7ZnCUpfbIHWYVZhSqh
Encp8jeWojY84bZcAzMIyWRwyiNOwtgIXA+ex3sTOnOIp6QmN/7pRiByRcHce/W52K7N8MKMcTnE
UAK7dXBnWaBCmL/4rPf48ejU1fokftLvbsIp0aNYhMJkLBF6KgAKBM0RchXpTyIAVMvrwm1ZpmvX
p6u/OkAzw1Wk9IVnK7eAwMLpgCGO20hqaQ8/1xIlZidXXVGZIOn7g9MVBDIscFpmv/K7rrXZha92
boNE/orvVYZND798MjDkBrBDckH1EVd5iWzhoFFHHU1JpoYxLd4ihu09IGqZ8Nn38UYHwHk+g24U
vYRtWJeM/LASXvX1Hy+i9qCP3jElh2d0QSOxakkxjqWZUMeVF0JA/R4lW98oZ6P3UQ34XAsAm6/B
O2FFCX1Gr3PNGM5a7V6zYOVxkOX/rl0TdqjrqCfum16roM7iJpIH2Dgo5zsX3G4o3x1ufHw8hhNz
w+OQ3L7hqEbpp5pL+nCaqGmAwKNTfnpzjNSnnnX0WOuS/fDX3gPPcobBM75caiED0MtdBMB9GTz/
WExUUOxapUN4QveVByK9zYQwTQaOfChmMkv25L2qOePNPaswadzzpW16INJBurM4c7WFRxakl0iu
E785DofkWRD4eQtroHzDCvu0ri61pRg5GQ8Ngu08MOmJqUMlUKwjXm8hvyQ8jc4oWjTYp1/la5gH
ingWL2yP17Lz4lt6VzaIzbV7yU3zmpBnWNKXEEEE8beb93bKYPtebQqhFRtlhJHXvFEEWd1DTUpS
CEQ0xU10cY46FMs/J1LdaoRSeUPbg/KfcAthkF6cphPnxbas74ahZn94Wl8OQ38s4aWMd2htPO6X
vE+4lYLdEIBR92WPxVLDAFrb+OERDW/fA+K9PpQ7reFNytruDX/i2OtZTTf9ynKBn+lxS4RCIY4q
6Ecap+ecfRhxF0la6JRKw0cXjmYIf1rSMvkgdTDYp2GwYSb/yioWr03hAlOyVA9OWTP5ORgd2uwI
42MQ5VBPdOX69p0Qi0FxlT011lK0lJX0vRvSr2I80q6osK00AQsxstUczyJ7EgIOF2iV/SLvKS82
u6K2mQu09FqfpkYh9nqK8YVfR8msEKuhgzK1EQDF/JneoQYWK+ouoPDjcWTW4PZs/91fxokrJadx
jFP59lbkY7hXbJHB4hgr9ZWSFJboSSTGkuIZgNuPjzCC2pR2Btd2ropYE/NZY8KL+NQR6dMHzmjk
z29QBR/+wmpQBJSwU9h8jJKmJIZzF51o/R4TwVPc33mrq70ngExM6t0Ok8w1sbqKqUUlZ+lk+lNH
Tr6/1ugIx1qUtarL7dLZaqW1SrgeTUC7DCbxUuFsozXFmW5F2MUlImB2wD7N+4UDtshiAg/4y4aU
b8unfXXwYYaSdODf+DELQHpIJpHghOxDNzkx9OxH92OrynKQamQy/epDwbGp2sh4/mUV7sIjwJXM
1yQpqPLBhe+xYbIr5FKp47mJ9k4yQ/7it4euYvdbjBYsLw0ub3p3vdS1AJ3VE4mILacnRVeadryR
EuSPWdP+Tc9sdzWM9K+8nFqC+/j0h0eqBj2urxoUixjzAX/2+OI1wyJEf6PaXv1WjBl0/KkFnAeq
CWcz2bqc9frNMf2wN0RI73gY4LJmjQZ3AQrBJJYFR5wQ8jbgln4enDJqNXJvMh1guQO34i0+FASi
nkmGz4QkroRlsBQhTXNQXEIkb7333fmxHBUl/zNf5UYWEyVN32mIboU470Ckj339rAUh5ye6aJac
huzeAEn0vSMwYHmBAa0LMpXvHkKsdf9eWfrrqFQjwZCroJE+S9N6ffSc26+dLp+LDnxSt0xV7SY+
jNKET4ELsMnh9BnsJwc4x5BmL2xRV2IWN95aVZ20z/aoiBIezlirjm6zG2lOqAihR4YBBgC+Bqqf
xG57A4EdbRrsygSN/t3wCIjUnnW9slAb08n9zQoYBB1xuEA8e29ud+Y3K4KDdEQI7zF0yNL+3yLp
VVSWQzOVyIKB7MqNM1Aut3G0r1HsvGU8+0rCZuI2n81r/XRnGjYyiwQmOIDXDLHfrsiwkWQLuFiV
TICObNBXnIW7H96NWTTlugRIGZZ6Bmant3H4eFo9cH5ZflWmLpTKg3etUnxEuPoEOfckWv+u2Iww
pKOgOKc/78VUo31KUl621pohJyBQ7He5ynrymIfM1WceYbTXHO52GyjNH5bOADkoeDnHA09ExBjA
n0mC8yz+ao7bsXQNbN8WLyo7+FzPMfPtSOOmNEkL/nFSbFBtlgJtT/cbjcxJcG9AktYviMuR6R9i
/behCp5wYOo+M0p96ek5H4gAnuNr278uUNtqHchLcZGorKUJEkrBH/VcQXJxg+bi1VOrqA95aCWS
uHWnXmU3VuiUJULSj2Wy41jNOhwPP3DaqqJCdTJjYAvx4xqD6HEv8BcW3HamCQbgoKCInWubQ879
h5kJdcr0pjjvaueZTcrzK50XiF8xfzengP7ul3Wk41F7t5cQS1euneCbEL730R17JesL18QDQjxu
p+qEQ4J4IldiAHi3UaJMMdK5PJw0Qvso5Re+AGCfs6amXwkWUiqR1PcHxnKyoyNCYLiFQP6ejgRH
FTedH1R8rWzIKAgRo0bTwtYZsO+JC7JUKCu2GspkFutEpPQ5zRVPpFe0OIjSPbLx8C4Edh65rI8o
B+nPS4PolRCkZxjL86ifgTfb4b5eOrn/adWtqDIqGuVBaZRfWHf4zVgJYR3ZVH80ob5Q4qIu0mY2
oWN3SGAz3X+TGQl09JiVqeJWUuQ9q2jgz/D7ujTBOE3Ebz85Aws93t3kdR0pkxxXgtdLM8V94Vcs
JPCV5AjcZPGBU9/nSIR67AR+E7F6Kqk59T9DlSER3lVJsNKPHG5AetZ65j7knReUTSp2xjsJptXX
UQzpayXfTlTOyhkGksDJGY76avZz5UAdWooBohHRuFnQXT5b5Fm4IrU+69DXQk4PuTi0jx8VxjIZ
9ySztyTYY2f2wg3fFYcGtmHG+uavOwrtTB9xRGwEwsyo+AX+hdkitsrdvvD5OG7d3KYOut8xPyxV
qSieFzFjikqGn30Otd6ABlcPQMz2llDR97/cgU8nRxx8OyltTJMb3WUfjFZpCdeetf0uU/qb8f+0
QaRXtnFHJk1FJx8gjLHefoQSzkY3yFs2XrFbnFBnAzD/X8XbNvIJJBgSvHOCmQiBrubPbw8FqEbH
1yoDgdvxt8JflzxDPhw8u4GrcF7dp1geSY35IqjicPP32MsLUGNlkgKGjnJnIMPv0O43htgswdDW
4q0LHuTxCfVcVPhOAsYjizi5tk88k87scfWINJ9Mz7sVZNbBCRZzlE3XPRj45kh9z5sfmt3xQkRf
99sgcATM2wU3A6YUGPfnb6mz21d7xMtfAD+LQAVs9Gbz7lLBugcLEW+JiV6AhBlDnFtZInjPFr7Q
n8nI4k3rst38EfhJew9hLo2r4kUKP9p5XoiNoNRUx1ayAi7uKr+jHQI7J8lknYZ4V5DlID7r9UUy
9vgZR18xpAZUwUaF1jmmaLifZdqJhhPbOsv4n/7HgSb9K/zVKA2y6Ak9/YH3GjUpG3yOHN8DxTle
wewOUY0q4wpcZYYyC0EF0Z9lJ7D95zw/zT4DoEsJV64B+OGBV6JJ/WQ7/Jo3rNPC6ittFwIxYDcp
9W3AADiBT4h5+M/DA787MaB+ChGhxV7pIRMPjlS3gtBeuLyRDdlnjDgj0GiFzC88jOWHYBWnAmDw
lNc9fjb2XtxuVBvjYuesjFhJo2zGUlrci+9H+9eG/rA1P+U/IWDHeHq3/NiuPMp9v1u0HDQ59hoJ
jgmeCT8xDdqU7ks4PpvPiD3yyKtXo71B7sH0o80Qg+yNE3Fnr4Upb7P+P3fkpQnAyRQJ+U3RvVKl
aVsxzidqoTmQA6TMJrwW3ExeOVCLDYEPultPCS94LVBU7w1mxnLLyW0vCyeFFy6T1ZC9KqwDGSSj
w96LHKOfspIXYAn84Pu5C4R8WyaVXcNikV2L86tMWaJCmEvG1mXdttmVypq5GfaIhYei9/hDl59Z
eL1ecpY879HqWZD5U35aLCOSmb0R1v7BbNo30IaKvLb3MnxhYgKUTFCspuD4UiQekht40HknOhdJ
4uS+6eWwlwjzRJP/K9/SkA+7db5fD1QGzZTyr1XkY/iDXCbJew3mT0Ps2/lNM87TI05AaZ216n1B
surFQD5Od5+J+w6G2EBRkrGYYTIyAyMIfpmv3WG+402HqO0KGHrQd1EC9NN7TXCiwH7cdIBHLNun
p/5Sd1cUfVjg7Ov2fjJYiM1JlOEcJPGm1bE7EHv3jEkQKCn1AM/1y+cI/gskGZ6zuB5I9hehYYB7
C3Cl5FqOZyCU8v/ujGGYUeAV4m8VhJlSMYo5ojJ1FkRfUineVQluzOZuuOP16t7FLuYRB0LkOB30
TFqZO/5htbL1Us/239UHO/y2kBWaGIElG5x2gBffhyi4O9QY6KLf6zIfODxok2Zlr9/FSG9dEpC9
DGH1m/Tzy5qmPqVgJ4BV+ZSgnpwwmye8NFo+RgEICNtXAhlq7/0RuJhetnJuMESrKKEmBTsfvE9Z
lS8ILxP2iXFlRfuiYCzQmm3I/d9iX0Ciptl+tk4lF6M0aZ6QiOpe0Y6mKxpGMo1WiTBjMUGww35h
wPNDFp99RZ4jDRnK/9VPBwBdsJX6EhagK2Gl/svtqcdDTkDo6PtGE5iCiIs1mArAUkvn+Hzd8no1
95MAup3WvI+bkYqr5t8pUcd4wwTgOPYOfyqTj0YrDL8KCT3jm3pDmd2ur5Ywc4rWtAkc4B4O5w4H
9q+4szajwAi14mxxnc/BHi3ZphuleGgYp2bvTRkqE1EEWpcyTwvnK9OjaL2HXtSkMplhE5xH4Wrq
cwgFpiAIALQh5l1+tusa++MtB5FQNdmJR09sbWTxHcaMxTf+YPJVklccJnLp4OwaT1WL7z8K9rAL
fifbIX0HDBh3+74JP5osAoK/7A1m3yGDBCDGTXjjHgb00BXwDcbf2J7eNwre4hPF7k6X4fxsoXfc
ZW8kz2l7iZwAYK+K3NMv55IGs8GCULIE4h4hVVK4WGSgRjLyv0EQHBQ+4KciG5DEXHa2N/AnJx1v
fl9iAtSaZdD0uPL3FhNOUUd2tIreVbRASXm9ay1tv9i0x2EbgeiIViPVjEIbQ02jm4VAsWZ+/ZL1
w1azXAWAxumbK85Zl13sd4gQxMq7FCJDwNBuTF/FwxUdP7+PCFmciCWV4DjsFArNZKXnsqViBTZj
TC2uZlon+ma4qH99oXLyh7a0lUzrTB4041UcbhqbKg8qsPHOoJIgUV4kJ1mlU4C6a64LpmBZtmQs
0SSzstMDf/7UUnJbBT6wfbB0foWroC9V3eDsSalb+0aNeGtZDWwmD4wU8EIo95nQA7uZ3ZjrY++U
/STfBOKGq9CU4X2dyNE3fQiRVpShhzpuP1FRCk8pMQJsMt+oiedtMHzBkzSo74dLJ9yQaogVY8vA
JbiPxyIRcKV9ecrSCjuHayh8DxKtt0B2xJcRz9i3gpVcZfTiuUWmkK1y2Xm9nYLtixUkGavdgwSd
LapSK+eul25e2tP4wFf4Qr7/S9I7Ri1u2O6kBQmbHVmseCjSCmbh0nxHlXEMkev5pmvLLfhKFE4l
Wv/oZV19ck7314gorYnnPH18SgbqX3ZB6HXCmT1eWbZoqYSJu1WcZJwnsnkOkqRvs0cYfI+SMzgw
aJcyirzbasApeVdxueH797R3I072nxn7jmAdG8HriO6tgmaXYfgarStwvRxUFKMo/SawxU4faKC5
TBql5c6A7kdlqrZtgNPYzQxskzZTeG3mH+m/NRw0TpIsgQFfslpECmoGdmkUzeVLdq9eeFMWRB9q
RYzap5M6cFByWu1QEAgX2mHSqlZw3iyBhpsNCoPHTmrIgRQFPP5y2oG76NUKqnLO7uhMTaRO55U+
XDjIxGJ1mA+caxQ9P8m15s6gjEr+azNkz0kTue42LaI5YWk66AVwXHajvqjmioFvE+t8DwPWXAcA
dQpBuQXahBb4RV0vbLTv2iaE/Fw4DyHIWDTYdwH/jB/bim6jvA35do2vix6vSWu/zFjS/OLeUmq1
f7R56XSTOijay6jDHUEHKybNhbWbvHCB0W3XFQKN7fDZGTxJ/sI1+3umES78ZczMtGFFDkj92w7h
aUXV1q3HtIk5jWcqKOyJ+bju2C4QxWUC1pxc1JHu6Yj5h+mfRByonStnvIHL4sXqEfj0fN1KCs2u
dotaw3+g2rjCl2r/CUY+IVCw1/0benn/Kw4OEXmy22fcEByjfY/7vSY+8bUodzBSSMTLD1gVT8Oa
AQETVMm2S+XP1z5VfYOiMvTGYoNO9eouVEYu3cq2ymEEVgfmMjmz6bhQR+8RgN9Qh4eBCS3/KA4w
Vg99S8e27gnEo/LW/cSys08VoHxPKzhnrmz4898Hc6qunbDiKvaw8Cu9+iOrUwcg3IuJ6X9Ho2xI
X2WNCvSmRn/JExc3pHzSyIfLsk9AAKtBn4SXs+P2KWRiD5OpnUtuLCGU+RakmwBrfDpGFCNotsC+
zCN8bsoGDTJo2IVxhf4kszz5moq9i3gYdd+aw8I6bOYDADPa1/81c8z4vOBUCBvSATwxh+GYZQ1j
mO2yW4L9WMyxbNPbt9nWirNa/GcCzebIfSdi+ynTGXlAdsQN/EIf6OdnhBVdKtUZFGDQaOQBWspK
U2TlMI5tjs2txuVzclHpxibDa3+1vYI/1D4X1qLh2xUU+bsvLa8WZHkgBS6UgedQXYQtnTiU8NC6
sGqCdEAC3SBXwbEqsjI+isb6MpJ/fUf9ctTIaisCMmB3hbe5sx135X+ESjfMWclCrBYljJQZBGej
m8PxMwf65z8g8axVUcf+8ds716MGr48U0fZMEKdwlWiq9uwY4s+GdMBoAdBhQ2fVOssKBn36S8sJ
1zGvPZlzZWdaXWxFPeSl33c7Ai4VhDuA4rdez6djWWLjybKHQ4WPfa3qmbM6cDdUqDaM/HKyaXP7
iCZcq/q3MAkqewQTitCHJEJVPGjNRwSFXywrhe4ru2+3mApU4SobxfbkYrCH0s+svnmAL5B4nU4V
CbBWTp+7BJtqU2kD3ewG7O8KN1VLbfFFCeBBJWTQL1Wm12x3trmuCTAHXyYSYHjLqi8dkcIktpyZ
euhQKlGPJjCzmpK/0Ijw+6GBNKpyUpIVMsVv2yzQjP/ATMy2GrxXo9Yv6/bd5mE5AiDcfR4UJaFQ
6yB8k5+f1lSkMZSyXaquYhrLS15nkeoxYKJZvzfBqjoZrD4fDy00wEWrBGyGqylFejlsaBdjQHQA
gOCIaW0Fcd1TUEkMsWwipRLFyvMNgOQg+XObfHD3MmjmGxGj8cxlU0zPZEjwYJ0xQVi5LoARmA75
b/tOUTw9JpH0egvavS17fgKphjwC3yCP9tpYMFCAQSjooQuS35bkuJBgqwDffXr5x//mf/XcvK9Z
xHjspBPkMMlKkSH3287eBWWsqh+VCI65eOPUeS8zC5LIzs8yw6MiWShO/bG01yiMwpgMXMm/aHH1
tPPad3jN12qUdvUV+FO5aA+imL8Ut6ZzAdnmcgfxpu2Ap1tQAnj6tB5Hd5OTlyKQw/L7uAj2pCpc
GmZQbkTh6J82mqGedWyj0Y6HZlelY7SAYcyVrpU0Ct4E35xFcAIxcxD3h8/OGrPYC3B5xAUosOD5
Je9u/Yv8ItLdSMSPXSr9ITQe/l0HZUO2WdkR+7sK4R/M51PP3C/4DFi2NjsFQoDGd5jc/3Xekc3k
PtAGd2CQI6tg+MssnkigjDQVvQJrCJd6XBJNM2lRrk1sn/uQo4mnarvEDywy+tvDLbJYWsi/uWmi
3j0jDUUS2bSE0zS+PyTYXr0ZcPodAEA7xT7rQp0crW5sWmS5RVNS6fWN9DkthxWx3oS8wTKUcthD
oCUY9ndlfyCfxED2zLtczqXfvucEDSn3U3G4BapfvGKWyGDtawOq+JF0riRxBzdvVpAlNgG7V53r
N7ozlOccBG7JFiTlJXlvvhN1cIWFEzWKpw4TdW0jqMigxA3Tmh+R2IzSKFXuURNFOL1pO93SEoOZ
Ldef6Z4iI6n/mpvUSEY44OfUbZvYA06FkNBdNWlwa4iHsVZQP1CD0bNb+RO5dWmPI9Qjf2f8X26w
6QiLwyJr/VVF0w/WnDqYLnQ5+PkF0/9C7a8AUNRf0u/DqwOwKGau9nh97Uq29qLxyD5iqN/M4wgx
6bHPMhG1pR//AFptJ+fOi1djG4bpeGbRSXMqPYcTotSvD4Zj4Qzl3QoeaHuCvU9SoLLjsJ203WnT
nycDOu74p1mD4PXFf1xwUQaQx1LnA/8c6bUP8kn/EO6u+fxLKoihPcdfh6z8US2X/qoqFzj/p5Zs
p1toFfCFoa7bsRHxDAZ7I2YE1gbECRFLAX6kXCTTzE4krcH95pU+PuMeFNqNFzDpBcMWChNew9aJ
FA4FUjQnSPTVKemdRccUts6WKx50W3H8Nhidlt6YQ26ESIcaPkJVPtA4BlLa+VaCaCt8FGwuGkOS
hxoVWGqlqkZShSkJeIIwPnwmuiJZsPiJFRVtFjyqnjhAtYiMex4F1gtFzlM9Dmq/66CQJzEgCqVs
9bOSRHHxoES3KMTusHdWeLo4Ol9Q6jbu9B+v1QiPJsBjk9JnMh80fVb5Y1NU0YPgGx7FeHOFnHu2
b5bl9Nwr9i6mNwUUbOdqJxqs35Fj9a7CQOgL0MIArN3me40ZRJX5VAqNo1x0p0eFFg1+WXBOJpAL
RBdblxfirZJ1CcCD2OHCpIVdpxUhdcZxtht43OSzNo0Ax/cZnXxiLFLFFHRwPhY2jyZQmYC2o4eY
fJ5jYPGgeOh4/Xq3Un5vfyoX6GwnR5vHaV0oMFSYqsk2TxHFD2IhvbsCyGSbkw+bvmLvZ81g2DvN
dgGHxyoIgWBaTCR0MlBmfrZ4HQznJqPv3A2CL0RQ685Q+vI4VD0MFg3MK+pqHfGdkSbRcf88NQNC
yjM2abSKyqezEFlyPL7mQa1UCYP3IRJzrWg341Nbfw9FFriR2Zg23ShAf4t1LAGc+xqfpzm0aY1u
XqqVHV0lDb1vfnJ6KlijbpwUv1gJiO9sQg0wmSRQeItaJgNyOiu1pcWK+U89uVZvkf1ThBQyDIWD
PFEJCQ5s8qI6+6f2W+HP/av4OY0n5dGfa4lNTD2um6csfysYwal4cCYURK7oHBp927PBkcdMtS5K
1av2MGrg7p8lNK0dINPRSXOoiquptIFIz7Q6pKn77k4Bmg70+cdBCxPEC2/IXCST57BAIxq7FGgp
43sUGbjA/LRaXRCOpAWZQ7NY9imZWU4+O/DISGhAL4VL6bwnCgr+PupItiPqpg894uam9UKU3+26
SWKuNCtauaPZmvM2jPDmG8aOKMliGkqW0xhS3K58SZIsRQy9qOuoumVSQjA4MS4R4CKivNElobzK
HAwscyOrn1WWhiKlpURms3anT+TZd8Hl2xx5Sdb6QiJIOkD4PdIZCdN1h53Cl+y0xsM9552qxj9E
fuYRh+crl1JE+ppGi56s4HlO1AtGTJVXs11sfQ3J9TzKMW+Z4p+ZFa0EQbge209oyBRLGKr5H81T
9S0eEZ9ivziUx9RR4QmwVZSr/mG7nJ0P6hBOSvPKVnSSnCnrD6rY2ot5nmxQ58GvXIXEJLtidk/8
aMqsTjKQHox6SdBz5loAqoJfqnttxGUKz5i+C8zwtGxeU/lIoTRm7+UiXWVvrQYpQ6nK6vQQNrb3
+OWz4maIIcJy0jZAkf0DZ75JRbZUx7cOMx1Co/HsW8bTKD9euKCNp/cxHmfhcqlXPlWcVo5LkmA4
RxcC1jvzYl3uRul1QG3ym6+4eo9y6L0ubFHv+lEL3nBLSWL6DYkpLT7fnvJX7qvD/GwoV+7lE3at
sDDgUyGK8p4P+JKuF/dCcuH0vOwM59kOs2iw19oSPUlDBX41a/hM7GANlVB35N8kxlJtrgd/Tj7P
urb7DWSLylF2FSIbii/a1mttil/PwNjwKq125owJkMaOuz0V0qJ98LW9GYtCAaqWUKzzL0IBP5OI
cXVItGBFDUdfRVhkso5lAm/74Yp5Ad8PS+CWCvYHFVM8q/nCicAiiORJwuHQGVwI8o12arnPVIMH
Q2WbqQbLb6//G2JZSHMlQ+iya2qtJv7F5F2r3DszwLYA9OSzCzflJq7DDn615EZaV+DtCxSj/41f
qPDu7dbGL5MrBGoJQpmcHQA8ZKd1qJepJiCfnV2Ypx1xc5Pajn81PypUdlFn1mgJ3vXo7gosiWoD
0MXO8ETkOCXpMPWWcM38uWeuqVFqLD+kR1tzdtE2EnZ6l/ZD8nG/pw5LsKJEep7luemlNnW/4ffn
rTcSO7AOnNPoo7VF8m9heMZIYA/b7zNCqhHeXKWgHNthGSocZVJL3gWiA8sA/wewPvQhB7aLpk6t
OJuFgH8Eec6jDpM6eajnZC9BRaSMEfVBAy4w4pCvu4s4ekvvPmKYaK6UZFhBxZ22VmcLQsXkpCTK
sF2K6RjND96AzW9TPSxkq9g0r5MA2eySAHIq69phMKm/JMmSd11suqjS9SdHJEIXhHMBiH7+9TU9
xBhNMOzUybwhsDx6LyIfLyG6t6wQC3aEegB4WCu05FAR8qO42J68ii3mak1Tam2cralEfH4ujFVY
0GZRmJKDLFlIvo2gyOiHzaeX5Hqe21ZtUT0y9BtqHhLWoNBwVWXU6pPH3Y2le7279F98P2SuPv69
6rJ0oNwhg6dLn10VjdI/+81KAsd/3SvJfabfvE/5S8z7qO1igdPk2Q7YSz2xlewHmcni1OiKLOcI
cCAWwpMah2IU1n7Y110QuIXCgW0R1rjSkPTi9uaw98tMEZ5aQoaHK8azJgxPJg9e2PEi8p0P0luB
oArLa1CqVmbucvd6dFxBbjDiofzoocd2kFfLIDzsJqGIDXuYIYXN1iZJJvMBujs4SJFonjax01Dv
uk1VQbGjeO+IwaxnqJRDZSdqaTWA+ZMFYlmvN7xtQrDARTKYncPmqJybtZxsZhKAoXxbbfgCQHrL
pWaAxBSHFRBUT6hbvRIx5gFS6xS4ECjJTNd0eR/t54L/ZckqoZpWsrVSgu3B/eriWCkp7+EgBesQ
m21wVz4VWbatP/D6rg1Bef3WenH+H/tjNiQquSAKXMoaKpqytLtG+/a8z9uD7lm6oPv6FjtbLP53
NDbb9Iy4VmH/6vJs2ADi99cwxVAftqyJ3H3dWbUbyM8nLkJKGBH1ZNt/I1r2xW1eF42CQX89PLBy
jJ0+z1xZjait2BqosgPWOPgtniZ278n7/tdxCfw1Ns8mdJ6sn6lWOJW8nA+AZvGtuiU5QYLSBlH4
hfrly8rGWQmmc82aoIbtU2DT3LTQh0hcAboQdcIv+Cf5sb76WTwwdavBfLxG5PXN+WJyDOL7QrCW
I6vjUIC1095jam6/MlO6X/cNbea3kOnSNozldusg57RtbLIA4y4IrKEsiUosVESYhZnqGZifE4Cu
7oPvFRL8wARuVdIoux3+xE6F6VCSKDXnIZMH6u363wvW+1O0odHdg/K7WcI5ich/Lra2a1asR1MB
CvLZ5UhSzzPq74gFyywPHakwQlAg4IwkeNvMNdVwwrhsMbWur592R8Wob+bLlfyuIUH0BA2XgI9h
G/9QtCOWDd75Es8xYOo+Q86/Jc9V9HYexPSZtZfssFA0peQlzxs4KxYNxK8R72SySCzelf/ubdU9
PiJ6Fh4IRAzGfbIUi8aFMQHH7Qp/J+moBNjXoOgDgnJIetcmtVzFuzrojajXOYYOcpzOR3cgwJkg
e7vUmjoGO3N9SdKwp1zlbmymrMv0DXbolGQCBzLS08YKevX0VWbPK5Xwu5dKE6L6T4dtwaFm894C
/KFRK+6k2Pc33a1d7n47sORI9OQWidN1SouwqFNwdmqWHm8fEPJ5PXBbYaR8r5CdMRqWcQ8WRT6i
cCzCFynkF/cXzScrE6asmXKkfl4OpzxzEm9QV/ZPfQac+iuG8HY9l3KjDJnTGboqu40cJiezEqad
K6IhSHxojxSOS0neikCTvo7PpEa3GHhAozVv7FUfdzR+bB3HZ1OIK4yHja9Sknab04tlEA0Tzwc0
t8OKAWznMiKyZPTwzekglBGhrB2yBzF5JwQDr/PwBDFOy3jE9Y+6g0rRrgiNmiUs+/sbVbxvpbVx
+AOuSwoBGkC/+hhEEyIAskP7Gi/eJJHKL/1a28t2B1RNdW1joF2KqQNIHtrWE4onXnFHxbfTE+HF
5r5jYqT84wPa8JiWdlPs/g6wY8VJ3l/jc39JR4mHREZ0tSqRT7DSixuu9G2LCsyjY7s2EQB/8nIS
kO0EKMizGDvo9p/To9qQ8PvgddssnGcoAWwNjqvERgsrPxtZHumchT5vOziRBJtInfAgCCATHTX/
DYmwpHqR2wMMhD1JPvVjRmJQvY6UfmDdKwrd4zT+nbfZulZWX72aM6y+Hb8BFZ35cDQtBq42cODp
UfTPvnQVu91T5rGbTcuk2WMjAc2Si9lUni8r0V/WdhXMI5jUWRi/6/oG4+045zVNYz5hfMoKDlvb
Y93d7yN0/1x9KNrhP96sUIA7wMBFXhHLaF5IuSo3oKfTUWeOq8LxZgQNkKPDHBbxJefPDNfqPW1l
xV6kC15JzQty9Ow4BurJwKNtplFRQdl41yn8CtfZLn7k07tD18BuvfqOeeNbHvXU7Y12gXBiP2d8
TCaHwd6ReEni6ribKUuMQr+wI3J3uEJJQTonAB+1rSsz3He7OfIHkpZbkE62ZNKlGxoJ6sdP+q8/
AipuGy352sNVBErkWC4I4ChcocOabpd6Wpu6d0amoikNIgq7+jyHJSToz31dcCIIk3+6EbUdcCXl
S8gYmMRtuMpEoSahASQcjBGnUk4kkQhtiE2m0rb+WsWXDraJ0jhEc/RzJV+HrowagsaVV5faYn24
yTV5IA1JIv5kykuSsGXyQbG6ClU0tmVy1w6wHNlkY0oHNuqz75uMX5lUQWuCCUo96uwxFbkXEiw6
dcY/jwdYca8sC7WH1MsHCFhgpnYOuveRA+MixbL7SIChvAeiC4bQIILHnp2+oWB1R52T8q4jGHWX
gtJRT43oBepxxJwihpfqoM89ktrOBcwJYsfTM97VdT7HN56C/HXDwXpzzLuSirg35/7uJlqXPmp0
h7o8woOxrvWrbw3IxHrZcv4gsx0Vb9PlmR2MP+TibMtz73aYUYNSVUijdSCcZTstukETbEzVNreq
nGa9ZoOWiOAWT5HtsKbPe0TBg65TzTNITD1k51nFkp1Vf27RYdcuWaajryyqqDLfk2SBakXlN0rW
PanI8B/Zna7/3UvqOoAlyf+A/9EYhOsHWVIsQBrLgvSD7zybsy55/aKOKcLOPgYnjFwSHVaWqlGW
enE3/pbfWbLiuYmgBG6BAM9VNvedgXE0+Yb95dUmHQpDILQnXuT98aUcf67OY30ZAbMv3/AsIVbP
q+K3wEISjGJSAdx8oBvjl5ATHNUKjVUOojaIKtIgi7uoGMfuQdfZpvonNp2KJUawC4S8Rni30HzO
gzJ8doTMPlWdmLdu6exgjwiTRv4CImgv8eF6reL4/x1scS8s7y/8+2Cb+9qsR9l9UWBeKp4Urcf3
9S74HdqUT9HidR/Gey3yeXn3uQku0julma5LOOf9b8A9TID/B3ai5Ek6ZoPcX8OCpo4OiqYReDij
gF6bYKre0XRAy7oWDx4GPP7J2KFelG4jdRHBOB/sqfWPfgdmElC1SEfzNAibaSLHx20Aj98b02lb
bRSViqGNTb0mf61Bt0oarBDfu8+Cy7KOcQnU2j0YN6661R8QSRjpy4w7hakDKkLEa8jDXe9j8ctx
XiNAfrpdWmQw6oeh+sblP5EYpqPR2HZJ33LV7GURCU69EDCp/LNi2LY77FL8+fU6COYRP7OFCXnC
tcmT5drNkEOUSaWFDmHbzu2WmnQaBkO2oSoxNu2ukgIrHcNlFzrtuV2hoBUw0mL/n0PDdxn8zWE5
ZQZzIRJUftDYJt/AHFdlVMFRtwQT7TPK8VTjcvf0cnVITtv1Ds19KlBZdzOe2BR6G7dWjitIZMKA
aaC9wGvEcw16WOvT2bWWTAZRO8xEoipNyM6shZpl/5gTM2btgABg6y7S/B6O4MVtjIRpOsG12Smp
qQG4fFpunS8Otfz/uAlJ58ndKJfT+vjU6zXnNrnt41xYqORHOJ3cN5sr6HHABPUibiOmLYC2xY+G
utPZV5glFBvWgi8YuX/ba2O7kpg//HHWj4m/u1TWmepXlO+Oo34fyay7EduZxFH5dksCMKT4u6XT
FnKWRX9xUKmT5h/z4H4rOtOE+dqTCMxSJA4stgzhwp2I46LbpBpv9PaDjkfhYP7R7yc9t/tlu/P8
zbVBoXJXFhIUAhovd8oIqEHpai3bSBebZM06EYD4nstvw2BQhDIP2G+PTi+6D7kxFPSPtvjVYSow
vmFlZv7Megb1cWFk26b5i8n1b3AgyipuDUqmd0xEygS/T1Z18+IGUNvWy6wwqmFor0va10nDr6xM
RxrcAN5zG0AHlNRpCWPVpOXm0vRqICcjJ/8gXJOcZOwkY/PthVJ2n22SE9r5pNFwKeJussZVgFya
rhZI6xfW6L7HeznojvO2bRv0P4Wb7oQp1z2dr+SUtWSUadU00zS0tM4Dm1zbZZMCbM5B7eTwuvhK
gFxmXEFar01m+tYvQiVfUHD2jrtXkE485Z/IPJYNQvOOqXVrlXKSFlrYjMFiUG2nos6BRkARRwnw
WQhR2+s0e71cOdIn7Q5CWx1UHHNBK+QBd+IaWgSvTH6AtThwMKywgV5Ki9BykoExRh6hsb3BwoeD
UjBdG5w0pkIPbitu2pYBTgzKMBlqvH3GSzAfQg1TZNOVXHNTRgw5QaQ1AnLfm1WBNJgzwY+tYXCE
k1QRE73Pffn+mHkWaIpocW1RYvh+4PjfZUsNB82GvPNs6Kjk3NIGBKRVx8GbQyLcZZNQDnczqff2
NytuJMz1nzdvv9Ui2tMw9dSGPsV10EKVjJ0drjvzqNCp2nxKDJpNW5z/RltbNOwV/Cmh2qGY5UoE
7XhlU9wzeRZBGVq8twMbS4y/FjD645Fn7fbAsffuTHoDFOyfSuLPUZjGky3+HJUIgSU0I7H0RBtp
FD49uELJJr3PlOWaHK3ennd47mNRdf3t0LYybw826rJWvlUmKlaxL9XijnEZjQnl9w55uziubEUt
+hJmehGcbPJHkJZdqBqpLua9txknYnkuvNOsYBEK1aR3M7wL0LYXB++1F/kjhJWr7GTd26fkyjyM
j7TT5AytLMmccaBSGDuMTrB2hkh8csEMNjSfZQZ75qgcdg7BN0ffA4VO7Unl70ItOXbvdJBeUyl8
cIaPbdmx9Q1ljCLD1N6L1ezgzozHX77va6lx3S4sdv55vxmtC43oHkwHu4RldsGLiW+Wkel1qS10
224gflD030Ri7zcwQimsDNpSreVcd5aP+OObuBt8FuSZMosqH7o+Rk8QARB1/5imf89KtwrfaS6b
yOQ/eQnxKpGg0H4iOUU1s6SkYrk3sjTHGCZX6hmQsL8uOFS/sJwIXbu9aR/MSNYA3hbA4XwZ+EQg
B+t21ZbNIeIRjnPuhFOI8wVZXQ7MP+iFYOiDoB7lXOieJI4mudgTkyXazbF8tUTyg2o/k4GxbSP8
Fv8CvAmNYEXlGaG2thLjidrPSNSFvlIxmSvWzkTTOZBxw5movN53BoaWG7vrvrVITqi2tGWPAv8O
YMaojEsamwtgmNRRZSsDlXjR6YlUAj60qsc0eSyCce+SgH8Qzbi99eTiax2LdmvBDvDrfYPyCgk0
Es5omqBPb/y3YCFaYNEwgu/JUPhM7A9cPfD05XrJxPTW/+3aW4qhJYmX2ng/VHHq+IXXA6d+Of9d
JeW6D6GFzvj/NDV0ji/4Tg1X5ATJkDcp6ATc6OA8lSlW3bjPgHiu3tmQ0gANTu0FGFnGsP1ZjeOs
qOJ/jAnmDhQgjLMpmElNPT/WPHM99Rr9R7blBQAL4zagnIlcxqCHNvRiZr+DEX03bwMWh88OOHzw
8NTdXu+saE/fu03dZboygnsXxIbL9HnlRJ9nBmU6rlChYsRdb1dGO+w+zI0xtHHDRdwMfqbdDbll
r3vh+fn6JwLPsvYE/Ayp902CFN5jCmKznjbL/x71/LYhxsZ/PYbEM2AhYmQ+Oyt9s7bEn0zggW1J
b2z8o3EoLh4XXHk+24tD6JBe0J8xvYsWwhI2POXJonrED1lh3anDN+9tPYhAwqHGW7q3uc4yG3zw
eLGe4L+pzUPIXrqbJS85UYujTz34SPdxFLRFUCSGkjypTG5TJ8w6IFdSUjE4AjBBWPD9/d4tlN+o
+XEWP9ckMzs16lftv3sM/8UQD5rCZOvQMBl0SF5Tc0az+wZln3/By9tHxjisNx2bJ3muXmfLE5Bo
cq0XoKOjqUE2CtVT13+FVKRH21ScyNQDgKIJ8+Rqxaw48X068F4kOtPdxZqf2/QThrO6NkyEfrd9
oiks1Ho1uQzGrb1/vG3d4BXRxvSuURybM/glUDroVO5hnaxKSNjdYSeYpvjPE1Ak1L1K6zNStaLs
W09/wbeDObgpYcAeC7SY1nLaySlJDPHKekAUqEZrQDw5dLCQEWddMHCN6UEiBr0q+yjBlfWU8XsV
/BUW/Smy5fVrbBcnHLbqOIZPA1yAwuJSznidmjVesYx7wsG8pD8AlO3leIVjb4TUBOvrjvQIHQoy
iblJjyPV3jjvcTviJHmlmotorW4PIucMiwoWPsLvJ7CPD9kLxygTPJ4dymxwTlf1qHebuS4yZyOq
BE1jOSIGWjZTxCoG1sLZlC8u+U/COBDNqqVX60ln/ibQMDkuuR7xOgH3H7289+RA39Z3U5t/UlLJ
EroZZyDlY0nUkJ/d9/KyfasiyZvvdK6XWacTZD77kEHcYrMgjQTj3gp5zIqRzQBb/Z7Kh53fA8zN
BGWQZC3+G5jioHRVM42hiZUVqbbfEI03AI4iUmWL7dmSVSwJ0WLMkBL1LrkC+0C4DUZYfsTga5mD
P9F0gG+U08JJmPCO1Eauje3rpedpQKGf8VesTJ0kebqgaU/s61KxtE5dIZv5Ja3VQyDovUFao1AE
T2zYiYwWB0YGcDWxq3jJOl/sbyRTQvFXTzN18p9gQ5EC5OFyUwfpNbMMojYa939NOBWMkOoLHX9x
aNsPHqDguWf/jE4pgy599Wu6ZDW7f+B7uk5SVG3rSustEYNSsg5eW5AFiZUYlWodRQkFehUi5N90
7miqAHORAWKGHDPPzSSPjtdwPsnGBcawILTlIUkqQv5hYw4wBi86++K2Ow7eBn06FxYWIPNJlpWd
+n0mPQmq/hEOnVdcBvDAhweGgMIfjkoE2JNcvZxc+uk2TJVIBx4Na9xJXrr+HTLpsD8cmAU3w97J
yk+vhn4AiOseo7KYRJ139foxU4CBXIliz1nCz85HXfgIVLu3xCWtY67FECRr1mfh8og6hgAN5MNG
MLhBzbop+Zl8gca0/C0UGK3ekf9Pu7GsYWT+4zoLSbk8t9Y5gp31MQv1U4bVMlGBuzaQSIGvtmEJ
ON5bf4z84HXa3JA/joD8blqBQNZFb7/p2BIhb5v55dC02tuLpbQdqJO5uoyJyHLLNTqicprOw2tT
GZZ+IOJrH+cKMPN+AU2PZN5nidLcEBsJCohGdaXA5VNerfhJjawk/EdygBh12DJgBW1mJfwtwedi
bHvNdoz4ykgSaFYYbz27PpptXNIkd/zjC3tm3A3JXpvkgKGRy5j4bEUzeoNOkj10Tzzhup05HoEt
wsSQrYKKmZByMy80M+Nx2Iyqg7+cAmDdRa85UhBdXNELVwTKbqP0J+zZD1OSEQL4RyMPFgD78x+O
EvS4u/Tdw6BJqUWJmVWxtYffiZdoTl/PvIBKWpl7p0IgESaA7ms5bbEKqvCGQGXZxodn87+mUrNZ
QcU7xGyMjhBSAcczl2ZWQ+CECb036GeHFS3AUNK0Gc+4A9aI5t3/rqjaiRnZgSoq5lIlfgmp9guu
2e4egIxcLqt8AbeDM/f4S7+OH+onmEaijpPp0BUPk/8CUNTsnh9F9Zu4M3ko5gjxnd/Njip1SQMn
v8WmkFebyMFiq1/TASGlZlrVFic3e6FzdACZt8gnpgEvWU/n6L7Uuf8/oLhPhMj5JQ3IY+ctHn5T
rf+DAvQ5bvvDejyTWqEhEiiMMXOXUlhamKeH+6m6cSqEMGnZE7H553Mqwm3WRkrA2mVLfSTyEcQc
vrZD0p4jXqlZ5FKbOItvu5he7uzWUYcOH/iLLj7HcM8dNeuIAWanIlgnYY50+YY2kBWRB03pWyHl
NRP2je/cBifGTmkKM1zm/aoZwRabpyOuYdfyNL/T7IvSUGr87tBaA2Zr3j634gLdlFJS+mJoj2yc
vg0bDSlntGBamQNgWm65e12cIl4Y+oWD5k4xmHAJJt1pse9+YwgunWCxIv8vaViovua3+a929+lY
wNqATc+tSwED4F+KRLeSUs/RSpASCEkMuCCC+e0io+GMMF+AoVVLN+euLvKhdcKBEEzF1xT/7nit
YuzBHziCfJ/pG7e+K6E14l2Yx36tThHLh1XvlVwu1yswehNuStdrcNMzuofUaq76RUooLaRIo4vo
82NrlnFJGEjZiRDytB+e+AHUSGDT96HEBhzR9YNz5BdBwgzn777kHiqAvLFgTpIuMpwv9o8JItHd
fMvBw2VC1F+zClSVr4AcSAcgE94EJ/2SUk4n6Dt44MI0u9FcsdqJvO95yXTXK8dcCxLjA+NEtUN5
PYwc9keV8bIJNrwovQxU1pr37Ez/RyWHIKeaKSqdjo4uoj9PvrMwEP6Ri4xHXAUrZJuoUv8onX0d
ntbXOvbIlPNrE6vTeJ3ZLBUMqGYzLd0TW9gLTir6YA05vpb6pv1yFDIXcn1A52TuNVY4Y9v3XVpq
gx7gE6q+jPmQtnlqWUgE6dLQrcswip0YpQUoOy4yUcMN4ctihoWH8lYsOqvzU2d7dn+soFTbHGIm
zgWSNieEol480j4qCFbbT1Wvw9Yyp7rARRdcB8YhBbJ/KaPLaKMpgccmx6wGWfacQxTgkYCBn3k+
R6oJm1OMDQyWc1w37hVhkiIuX0IvRvMau8Le94G1rLYahN92aIxLSLgen2Nq6yKY9xWumAlaYbma
JkduNtUhmUQutl0UMaDK5/mwrOQgP1JM/qLm6c0IaPHyBiChC0tvR/vULUXkUM5G9pog3HZGpGxt
rHicbPm9qj5es1xDTrWdKpOLxxQ5fFIcfuYIc6cOv64YRqyFx+TjG/n0Oo009zq2w0s/oamYEJGi
L8F3QPDum8tail+gtyzECYMYI86NP96gr7TUg8Ze6pEbDQJ1sBaeKQK6++6LEXTLGOHfGA3hban0
QrK5199uGKl44JD7/xumiMZRTKzrA0qMFzfRaP7aigloiBzUiUhLOSj+jTuUJN72P1H8E8UTG5t+
xKXLif3iLCAHx0zSEX2eQUlqr9WdUvKVJGVxfAQzknYI8uVtBWcZ4qqG9ozNiaWypZgrh08G9Heo
jPUrvU2BFv6sCXWSMkKOul0rgHm9P3VjC8AFoT0wEQp1SCefDuN6NhFZHQ2NkjgGYIF7XKHf9MmT
0+qTZIAdd+uYQmk/du19/kSWbPfWiOhctrCVuRBYKgZy2G+969y6a3D4khaAX/TgJQHcZzgHS8q9
hgdqAyTUe3Ya3K5Y0ZA91buElEDgidEcsrNPjUUwHYo1UmOgfK9NT0JEcEYOpMrmFh/8B/FPsSuj
Nz+iqHL2OOW6qf6+eYnlR30gDCx8uezE9CkmPEcgJaNwAkjBHBOIbqRisgPP6D+QwjhPgpDpdndL
H5YU9TSgniVC7Ycn9ertmpji6FUMcWHPbEgO8cVJGnvzqle2jBa+Vv1uABC0f33uLgAftsjHaPub
60KyjQpZqQlwokB7JneewHZBIxd4Ni32QXzbBBDkpbwOG1SN4+gkTJHZx53UCG44FGn3jGKNr67x
mr4grR1ZNiR/m/9zExJ56haUaBsc4//NlUIBR6qjjfbmPSu5p5zFf2ZxAOz/sGlGISzoe5kmhb2a
+5bYrsNoZ49fBDFcqm6DhqI3zZ2xtqGEV/VstSahvlHwv0SmiyeCGqqHiufkVbZsNFf/iOiW39kY
TBbRxt55lJ3PDLQLXL2NcmWcYnDDNek7Bj4OzdGCuFEeEgxmEzc9GmX2o1BgWP6+se3SX5c/A730
FXF7430oNRR+ABi8D0o2IFKJ4HLrCLW8MVkZxZ5SdRXaJGWX5yllIVmK5QDYGN1zxeZvEg8eMA2l
0UkwQsD5GeQYxxaeNj4Mv/wtaTIlCRefsBd1Q/tmUgSv57Vi07GVi753z1XGfs4LPYgYYXmujw2U
oUpvlEszCLpbWuSvY34OTLWCbo6s++e7wUBp1YSxTUPu6k+IQp2E1Sverx7/yHy8NEoU5SfjJJXm
64jLQ5plVUzEJeolWSw+d0iqkA7NrhYHz2bVktLapEtx4ZcI852Kw0yn23KoFia0Ug33O2TcqOAL
dN/P6IZUdiz49Qdmyb4GPuS2N1iid9h6Va+/WI3Gr6EBk9t/KBzWCGyiFDh49ENhQXRC2ANiDk5m
ZyEchJags0Ow95s6XxtOxn9RUpUvEbBhwuzH2/ENy2jzGPJogIzbZg6PIcNKyFgBc9YvtmFHDJWR
yec5a/2YoKscsH2D+vnr/g51K6/6+wGdPsDxTFJe3rk+rpEmPFCUJ+C5Z4742gKCIT6n6UWGzWC5
o/jyUpHLxl5tLexNiIAGivUv0L+Aj9iiQtZKxXOQkNemzGqxteOUr86c2Ykh1bePO2A8bvha0saN
d69F75S3Kw/IFkLu6sym4rGdV9dDSPHR+ki/HuqMrv8zdeQ0/7g2HIC3NY+XU9BskKG+k05HZpJv
iRlRXMVf1lNWc7+w5HaN+CGQqtTn2vQg+36KmUgxJUO00o6cj7wN4ukeyIRzNgb4RHxHfRCiwy3m
t/cFdeIBg5ZaaUblHIGGiCBubQHx4uZAkZ8I8yHRX7a4laI62/yraJ9I+6gNhApJmOoK3aS0dELG
IOp4R5eomwQGD0gEuEmGIYx6RtEH0GbX1gtDZn/eiwPXQLMDSVQEHfw672G880G2/qZ4n9jTg3DQ
llbro55gsyxAqJja5iY4a8N5lHh8iRh16mXxvr9Xbmht7FsRej1m7bgFU+eGyBRwFfMjlfZrKl1A
irOPoIKOSSlAEH37So99ku9eBfRqZO8jJlBNqMANbdjjiWnS3IJJ45KXYiSolXrgyyjWQgDX/Mzt
Gs0uF/h1kjXwIMZgJP0urZX/bm4+UWWX2Q5Bh1YuI2qtR/RQACGO+OhnfxOaDPVysQ6xO3cElZgX
ERH6xqY6riKVEF3LxVIk57WJQFlR80AJX2C5bJKNX6jLB91N3mfv1t6SdSJv4Us5xo80jmTBsLR3
fiaKcbYXHb3hB7wtrO38vsd4eayiqcaHrcaijYHMFp7QWZ1rDk1R2hdFUItR8m9gptzjX4Tf3und
ZexTm4z+v84wGZz4eqUbGKl8Ct+REBOdM1XbKGcYjb/1gxavErL3FyQ+5MPKTO83yF0hRckKvSDx
BBhZqffUH3B5Ji6HJ7IlyjGT5Xm/Lgx2ANbExf52V5v/0p+sszHIh/GwgQzeb0mofs5r8kdU7IHZ
tlail73Y4eeBYkxprtzjJtiIL0gqosCEwShYHqxpbbbTujbBnJA+aO9oPSDqdVkNDAwPlqHBvHqe
kNDdFubUQWncIzYSyecbhjIOs0/HZLGosBpsgygr5Zlkow9F2B2Kbby2eJ+1XdBam9ni2MxtrkDg
r6LNq9usIV4On5J5ZHCCWc3yp2GB3At9Qpi4meHU8DvKa23/bUiwOJTGL+empwbuUN6m4VtAmlWD
6z/jkF4Fb+MFGrjLcQ2jdm+6nnGKrQ7UzX22oHds91Vb/soJmr6dEjOmfjZq8/WiXVql6ePhymeh
2KZ4DFGceKbTotzCZnuNlnP5aZSaz9qKSECO3Tp2CCU9rdaJQi55S8CnJoW2hX0Ij5E7y1y1XLKE
AUs9CnLbS7cC9Gq3fP76TNa7uXVxgQa5DS5VylSCEFHRogyVSLL5sLfnZ3Jka5Z6kkDxLORzWSYv
3iD3BtASSOUQ8PqINMir6sGC6fQuA/0UFD/EndME84syVJWdeCKImbTQhRyzBFC6iJkBnYJ8CKUb
1gI38FFMvnu73e2vO9eWNQWh6uTT3OekSaIEurTeCvJgzEH6WJWTRS6oDLJV3/eWduCs3xlP+5ip
briKanPT5JGtIfH/Z47B+bpI7e3CxetSbwb5RntwlvVBTbyvz99YMqw8Qo6bfyrV8oj9TC9xXFpO
YgiTDNZI4HtfYZ0b5k8isHpPIsVHBx0evW5uxlFqnIEGCQijQLivf5cdqQutmCwqWOUdFRfv6lU0
wprjK7of1yl87EUR3T//wvYCncP3D3WcJxFxtGbTZBgikQuoF3tF1oSmogtYfGEDXZvFSqmJCuzM
4rcR46B9iisE4D5iGCa/PPKPNKeRQ5Fdy8GNUttUN68RQK0VYw2rWR2je+PrB8u0yuSTbvo7f9Vb
YuE+G0ucwYjdyLPdj8/zvgREVa/g4pnZdz8OqXWtmPanUBIjuzW5sLiA5+HwWGO0Z5DRD7Yjiixf
Po3BwzZVvHl1VRQbjPU0NwiNx1ixPZFqUQxgbIJGvCiKCCzrIYX/C5prHjwBOiR8syUjZa7yqpK7
Ver3sP1JVbP3CTxCkJ1r52vYofR2iUswpQrG6cspMaxBBwYMzdu505uX9sMiIiF6sHAY6GVuNdQp
utcqzYg0vhke5p/g8WcfWtkZghN+55uBfE8wBNZX7EKhM7epYJDzggBpr2LgkBXcvnaAabnlIm5h
1DRDjCssgqUDoiwD8roYi42+4OR03izbWT/xN4n8cqjo0ss5bqO6mo+PKHGyJagpUWnY6ahBIhxs
MtJS5AlB3hby35QeqDlYikgHlPSCAdqW0oAodYOYDLyScDmD3BZtw6TUsqePxDdiirvDKC5sGtLE
IkXzjl6RnvhTsFuqi82g3YslDApYbAbRUxenWc4rJ7GOHYTptPuQY8ujLJHhakUJZpc/aMvkT7rA
hvxaV7R9nlflmxvMyj0WtZp5sZm9U+3hI/z47z3rnKAJPQo8mkYC9pHG28bEyXTV2AkEoDuO675x
r+iswTw0ycH8gIYOwSwCc5N2VccrXv3RjnyvcWN3HtVyfuuAXYr6TPREhxJgLu2w/rSq8oTdvAQ5
cgVdWmJpW3cGgYZygNMZt2DmIGbMVivbGoMTWQBESvaFqmG9MsNCB9JGnqOHUxo97JHQbRjkTeYi
Z5/p0kphOewqXwN6vEakyWRrBQb/j79ukC1ZRbLCQr721tRVcK2Cwk9txy/WVY6k7TPDrlJiTMpk
BFPR8qIF0JUm7kgCtf80cf7VuUG25+htI3oKCzf5NBsfCrxqkrYpfnD9EvALCSsbgNxVqKOV38I8
pq38lfW+W+B7HzaqEvKcsmZa1tKkoam9N6nXBXNtSvI9cfCCLswerKR3n1vYw+3C787X+XLsYqph
S/WpCEzjLWGGgLs4L0XvMg0fTkD15acXgTVT4FNiapnNMlhH5DdkFA5TykFoisLpGO7c2RaYtKBe
ag5j/APrcQ1pX66oWb+pUnuIlizC7UVGdipECnmHFBFmuczCio7e6CdylQz/85VXU/yqbvz62TbH
PUUCf7maDdgbZJ3pBR2V5QRG3LqMYBB9LNqIJareeVU1nqXPOLXJZV0c1sAArFceOyc+F1HK2p3V
BlbGvzvVwnURZFli6TKKm6fJA+0OTwSSBeLDoIRCVYOa8bJCCZGqLpP0T40QwiZL05kpman/ilhs
fai5ckdLueekXMJzWu/e2DZ3g90WDe6qpDELgTbdUXzUA5o5iORoT5+AG/DuP+kKwIs5NMGdbm+2
BC1VB4QZEwYJHAq0UoZEIaKku59SXzYTA0MnV2iGI0Z+PwKM7FsMGphjy/nzsA2ACI+qoa4EkuTR
ye5F8daEXxp4TVGeTSyvbeipaMzl1Xij8tR+y/8Zhjs+ohao8YHmX28t9duDSYMQCXom9qFQ77JA
N4lNPMNcKvcvxauChUBMOaHyiVq0OMFCcMBKgbtfukNhxS1uOaykgS+ozPb6yJvQwv9EEgWbD5Cr
Zk4ay79KLPmWo2ksV8MT/uk3OWvArCzkjpMUg1PrT8Nuq71Mn6Pj1TZ3baV6yt0JQWQY4hRYsN4y
EXzBBRX5+QG0MfkoZsl9uEYPAj5JKHXlN1lCH/ZuK3jSEvwlgY2+OOYn0P/5TrmTz9upfvTWE9xw
d0jSLCD6nb8HSb4obYwSHiDbc4VuEKM8JjMaaxRpeq0ngUcOI8ObyYHlGoENfLaTvdNM55djUSzC
ADcXwRho2BKmsbr4ys+mLM0npjLKkoB/qPk9fbJJp4+EQuKmmGyv15zAgprmNEug6/qIjJiwRPh+
JF09WSjmEcjr8raln85IO9FFL4XF7zSSRIt4htarrNehpFHX8Mu3c2zCX+LGCUeJ7UCXh38fv/9u
CQvJaOhVEfbUBprSF92lolnXmH4vNsr+lUZdwv/BSNJTuU+xtIEMRCqAF/5irtdhgP3uS1fMEhdU
QMaoxcg4Or6MFSaKMf0jXL/8ZpY3J+KLzQTNy76in4wCUmTCo7MfzXHIiESwEFk+tbNJLfZBTzPF
O0TcKZwjl4TBD3I6sRy3hayml9N/REO0RwMevJ1d/lMr6I2vNzeneh/7wcz9fShZAMwSizNTttHJ
bauLPJDDo5NI+TfkanKqQb/vJDVomTvUQ3F7eRBeCN+QXuqzl9PvHQYvpn0zq6D8Gjj1+6sU2FiA
Rl0rMl2ZOCoMKXeU8t6vWL0BCteMEV8rw7tgvT5DVlDigU20O/4BjwLtJSqr6jzL62ul8h3p3EuT
NpmYefftDzCcO4D9g0alYuWsne6iBTCo+U+x/Kgr2gnPlPrWZhWN/qs/ScZ7qGWe/3i5ago+PC4S
6EkdPpgqN3Vt1bEtsyIEruHfqFGrOHoUyhRA9KQ3kea3EIOylXGOV6foZvpVvHDtzAW1vmA3F1EH
juv9tlGPsJG9RDTZVbD69DtwP4a+oKPlA5rTBnXyd1bDSodz94Z1eeesxvhVg0cn5UFeuS+/7OIK
H6wfxSqIHup3sh/0QzzzzmucM/i6ErFJr1hCFharmQXxw5dTfsP7q7Uy9mloiHeBCVdpVQeY0Rez
sIDAmjeapPXtruuHNadai4RpKUwEOKRel56MDlJdpk9oeA+k0qbu24iAh3rOr+Gm1WeATRS8dDVs
i+G9zvOaXGoXgLimnu5S506VBsQwc0XtC0izlAKtQQ4liu3oY88Udv58etzU4JPqUqaoqvNZQfa8
EGUp8au6AE08vnAc4fFn9kxml6uHTIRMivbCnv5VyAsODnb4xokoBGOvM4Ob4EKyZXY9dO107r17
HD5OEaF9VG0HOzm/h80lYNa/GuhrbSZe6asJurTuyw35DuRBDrQ6fRU2f8p+82mhe8bJkZxw4+6t
VUh+hns0hMZu8IjXxTUq1aQb5AzPruBaii3W8xpT8sU4TRXoSIA30nlVm9rHU7Zh5tQzSfK0N7E0
Bh2gGM3EuTjutFLci4QzyAWLWwx4ZZr5fEmBB+0c9oyFaomh1RSU4J46xEV+0GFNm7TbaqcJAWMc
3OW/piZ/+0Dm2MJujz4POeqVv2oHCZNOVl86J75Q9rAGrTVhp9hVaHYKOQ4YHyK7rjks0+RXzfWz
svNRJbhSOgpqfDvF7MkFp4GcqRFs9dJVkJiD2xCrub8TXCdCprQcrtnS4W2gAjjxEoDvPOe/bWr5
AgtojrlKfoCqBge3CaVXfjCUbcpe5cQIZgFFnTGcVqyPf2lLsIa5UZVpUU/6QgENSQT/8oMgjEzs
sWggvlbGC72AQeiRnFyia19JA4fgCK+UZG9u0jwHlWV22k8DfIFToTyQs4kVsYi+L+UUpcRyB51M
a2U1ER6Jd3Na3e7YdFbgBlb6wJ5e+ZkhKcrKDfufZjFP6iGt74VFc0jp5RKGhJDxRs0gHfGiNDwW
Sw1gANQ3vyXfY/ua0IhBgIi/hpR2hrpmkDDpZ7DxTGPIyWsNJpDWQsKQ+xkboZ58ZLPbKSxB4jp2
EKZfI+i78dElYYqODhcQHaMaLmQRSDOgdfKL+hOHx7R0/CZ6qS+C01VysUIs81nIQ7oa3mqKfA/q
BS3kgRbKVGUfVT2LSO/cFKbvaR9J01oEaeTBR/MPBMLJOeNaWAm99Fa/havxdNHrQ9GGDwE4T9iB
iJ3Gf0EB6B0ytMDdK03NXfbUNNFTCM+qfnVljCvlR0bIFO2sQoQf7xJ82zE812ZCoNGTSzKBnP2j
x59cLlDxwv5PQABkeeXdcT+wc7Pq4gen6PdJsVIYk+ge6lcTm7pnoX4vIF99KI5vFUYvt+5DRAwA
/6J6YAsFYjG3roLVCtWbQgco62/gndu+a1RXTNSNez5ny3BQfNLZAo1xzYQOUoRh2SkbgIa7VYvD
BPkH2dqpjWIb6ifsEHBAKiD/R99zGc+8AiKOAkPezTfTpKHNCi3M8vK0tiDDaaOftReI25mwo5eo
em1s0rW6tkgMHGin3fRzuJgQMtvLGaBlc02JO9Lvi/QE/wWW0SSaeDJhVVFeujvA86U9zsqE5HQO
LvYVOAKkU1uncM4/TwRA/emu+NfLc0f0S4eq730smxyrIKUaXVD+4K0LfGi/FXTDSSRaRYpJzH+j
zwsmv4KR58H4R5APzTil3C7mHYiDu+RctDIsPBZ849k7sE5mUvqsA/9S48hhEtU3Qb+OnZ+3JkZ6
eM3pl67+qSLEo+PhK38a81cxm3AvTi2vJCoTt7xWh+wG3FEqZgMrgavxoI2Siv2l3bykjGTwrxnD
8DUbR6nCcSDtIDbZICu7lx4vcaXeus0yRKIv7T7DOU1kRjiHGwGAsaDRs/MtAd+sebAvxJpcoyYG
80HOpTNh+7BFqxAF7EmSfYc7PY/rEMVK8NAOryN37k7PILP7S97XoRqVGYmpgRHV2EULRxkOXPed
dgaeOJB+AQQNysf8TzYoiiq7fTxWUfw0zDTlx/3r0WqcynoJK6a1SItJdtFwKDev3Vy3HUcQOA9L
eFJ7JHfGtit2eDCr8pG2bPF9hDORSxoTRPATuHKJBAehUUEZAL8lKV0GjxEeYl2tkPqSd3HBmuP3
G+Y39AOy6YITfDDGEH6GKh+M2kbBWggZ6w8fDon+kgEb9Kc8fU27s+1Ow1I45YW3UnHwIYRPYyJN
rMC2IY547s9KbnX33/9Tqrh0GMjXAjBsBYKlWoNFlf0EWIiizAHJTuiVRqckmnQoC0+w8JlpeCMk
C2PljvZcJfW+KVZOkfff2u9aF4EqY9kSIg/xcDkxlBO3dfsS9Blyw/GtXiFFFx9KU0g5vla+n7rw
e5VTAneg3DowlEarkf+0R51JFDA/OVGvU17UTscIJEOobdz8IBjQG1YSR0RroI/GX0a5Px0naO1g
ljUkbsAcRRdC1QgmHuj6LvwqvEx1zpKjagIqoEsEkN2gyHBNJTo8gVUuP5CnxNYVZIe2JBWxIOg6
Iwco8o36PlLd251IyU9IkRoyJyJpv1ftheN1r94oX8Dux/NXSbpShB3DYt3G3gMcDMPfungBamwp
YXKXmCznLSqVXjU+0CnJSOMLZtxMdw8ccAvuo8FCtaaP8aH4ZQ0LtavydlxdfY0CayGuh6b5sVIK
gRF7a17lD6LZnuTj/uWbPCTMXliNQSJXa1c/gdaETk9JdQujmYUs2AsVtobMT0+Yv7m+i4HLpRd8
GhRNrlgjCB16o5cUGH7NhvC2rznCG8qvVFC+mUgQjmSR7x3zYmOqb5twfviYyV9ApdL7g+FGuFE3
mDcFVhctg4laPtdYceA4xBynVHZgkZM6VzL+sxT0+w9xGweiVmhUocqB2EQEvtzofv0e4Kfx23WG
YO1++l8tLHAtPwGuIJlSjvaxryTS+POALyXz0Ap3VjtD4a4OWoMzUUxN7grzKQp9k37/eByaNqs/
v6xdUVk5fDHOgjncerbOzSJqVmYx2qoJfQFuQ0CSm8PkPCjDumuIde1K6YcSx6gIg1d+EbFm07gw
P4K4D/UoeD2aSkk2udHkwXMo5ZIk7fKdPvwDqgXI9BVAgYeXqptjHI2tlnONPByAIChlAsKOMdKV
EHdmhUrvHmYy6I9wsKcRRUJxElxabG1qOs9FAkwu7B8iIgbKWQJnfRgfbmqXSkRYr0ipBJiIpZNk
yFCMAys+8QL2Tgd9hiIgX0FjRaXVLS87KXTn68aR+emggd8VH3JkQ3RvGm/5IJZA/I8rakcI1slL
fKPbvGK16cZrYuY+/+ETNfguFJfTOSLCoGPhmXWlzg8KX0OYMCXRtbh6K3j0lnsZiv3tjlSj7n+6
3nVPtU871yW5VSCv4o4OavvRb1LA9Nr9BFmvX1ZVoLEd5xfQxIIdBvhxeunwOhkwkWGPJHiFgZ0J
uZ/3YpzqdGjrGeG9y7eUE3mUr8xjA72PbRchByzFJdOv+HhEGd7EflgzTmdNTlRr1y7+81/+XREa
oL8AO9BBm9xRVhQR02CyPeMAAjDBDocEKzwAnI14ty25XoC+6oo3i+ryBCF67VOSuoXauRYnS2er
RrNOB5gNMK/lQx17EI1ojmY9p2MxEf/yiCCeJPvlCBVPj2+xCVcOlm2cp6YpyjX5vQcJ7uJToNcr
4qOBilT2uZ5PNIapb3iqVOdwF32Myl++2miwkJfrYJKrpyLFuo4CouT3gM0C+8gVWUs1FVYDGSy8
Q+f1NkGdYgV/oa0kmSWovhdrM0Ou0dmLxNZ9IE4PAnOgsOiYy72brhFeSQDYwn4tNkHq69wBsnpb
dJtnwLnZRN2pTLIF/57zlS2osmNtB5RCenPeW2GvhGHryrEClT3vhyRwTcYiEzKd4vUju5Yr7MLb
koOF4c59ZrlKbD2TKlnmhmIh1HpkSYotzr/o5NydOjZy4C6M/J3tMUOJRXrnb5DLmKlLY00IYHkG
9Y4vBkGtQipgnuPmgAB1NMsvTGzKFvHCnmrMkrsie2VOnzPMXtwJyUpisFGv+QXelfEeZQq1FPXJ
ILW3Kp9f7ucC5sGN6uDRnNxcFbncbhy6pU3pK4JrSHJN9kLKCUUUPIiOerPmmjLqrdOI+B8yCRPG
raJBGL85exFlM++l2VZBk/fMTet5NYaw/AhZZVEEN9MnO9u5iWrMXMm+smTbSAWlKYaA4As2ROAR
qPFMlNZgyVDOgs3AqaKdlo3OA2QfYpO38xPQ6yJ4CJLPno26BelHp4fWqJaG41lL7OyWo8oC+j1E
c9oKOsbxaq1aR69qB9pMMGZUwNsBNbHPVUTKnvq/rCypPi0pyLYEkC2cn2QObrRFYG+oAHPWi3RT
blWqu2WLHZnya3WGytYdzKrKPVi+VGqQfFFIsckXgMbRhGWOX4YdSnd/CCCyTfBS8p9TNXyXcd5D
AMgBmpWvtykl/9AkqMaX12HKr93kenzdKrLzB52sh6XIettAXRd/ZyB16UjWcBhQUF7v7wU4ZPt+
fia7xwVnKTvPof9xIyI7JlGoJ9gKvdNXObJUu4bT8Se6yq8mCTjpr4N64FR5+OO0Amd2nw23dW2g
xlav0jFtAZaTOegPZWF5hO3NHrxP7RoJ0RRF6GQm0WTHfJZGJyoDCKSUQOYCjZyAe5IiIUMCiCPu
0JZZVHCQXA0ym0bNKENUgYMCZcpsucLNXL9I82+5W/ff+ZvfezGK+9BvC5OtaNuT32Zxf6963ljX
c7NuW3PIPZdJh8muonD6X33LeOB6V/u4J92OpduormSTPZDCaCoiEY1rUdeGBI1E6CBvJE3i6Qd/
jYYfETTrDI5Jcd+Wfoh5T7VB9LDw3PkW+eealgHrfSrjPx36E4ljUmnHzjJjyHRG5ZriaElcp/WQ
gnnosRdOT5UuP0nahywZ5VGF8g/j7alxWUI7CEpURT5yNN/Tok38nVgibziFasynv1eODz7miwjg
xowt/1QsMpRL2Idt8WcrQ9zsd1zKFZNiDJ6J8F6UWqGqZCgQIUq5ENzvVC4CXo/6XHuNC/trGFL/
2h4P/dFpHjnBoEmaZ1Xmf/lYV8j8c8HbzeUYJyj/K/+wfAqQnUAHE58O6mfkrGkcnmVK/NLWV0Ps
QmJZhBxjIj2M8Jyz4oe37pHi8eET5heCJdgfIzI7N9nHvB9nSRIXCwFu2mef36AU9z1iA9Jj/VhL
Cu4Wt9LUwqmi7k3RGAFJv6wzyGzBZd6CvyD4yTxMnzbVvpuz2dai0/U9tQF4G5NfUqppk/3To7v1
TAW4srs1NdwNzGJXY5acpOS8I7VUjRFaxfEXOre8mNlmeb7nQ5KkxFPrUQYzD/1Qrk7mUVVojDPU
LWDZCsiW7JIfW4C5WB5CG8hqLWEzsSMlmrJ+HNkAfGVnrqn1s5qKLYm0vbniNlVTaTYDnSgpPheo
+0F3GI9bRJa8KsENUFvhhU/9sp0eaBKrbqqVDuvMoXGqx8RXPycK3QPp/7kyZtLbxo9aXHUyzSZC
F+spn3sJkOdmVQbU2KYjZ80naMfi2s0F6I90e9K1uBIG3H3e4Uv7+jje3nqviPPXm6cH2TXZK8W1
vJrWiY/3DsB32u9Ivwjdpo4HA4TklT/Fj8XtYyRo9FqBbXpO7axewcmIg5k4fzRXVwRHivTtGk+O
Vzf5Sx31fTNAXVkOf9mSZy0HCz4r34VP3z+23VVZLU0yq782ADbNvYcY/fNmWIMoRfEN2WLCMLIy
rSYPDegM5Mxw4ssZ/SvuzhEkFaGcboGgnAPmU3peE3rudUtmMTTMhNWWMuZAjKGQq1jJwjnHYzS+
xjJj23NjgYsgXY5f8t6XOxMVPFRgpQjLYDef+CfFgHscj0D+6Sx1Cj4K7n6/5nwNaxCMuM6yZbAj
HzpfYhQssAhsrllwouvtdghg2hzEzZHXLRLi3BIIqdkQd8pFqffzU07kDs2F2CBmFA1/PP76zEwQ
JlWwUyF7NUKa7WrQubs3F2rf7MishpEp65Pf08fDp7frVEFHugWH33moBy+yawa36ZIh/bXdjPvZ
BxY0e3eNwkvdrjKyFmG6U778IOF2QZhdWvZGpAfYiUVKnfgNj89Ghmdk4iw+QB+zyiBkx1is1LCm
Q3BS6iEDdmVAeNjom4+o4W2zEBmFDt7pMH3uwyHr0u3xTYvThJhv7SNU1EoFofLTGk1vWW5/Rv7V
QaC+go8kST2Jwad52oNeflzlxuUgFh99kdza8ZqITwJLZ00RBZMgdf2ynuh+NsKngzFlTvcBlZyZ
vzSrMMYW3QXPSisYrwP6kmekWJQPosfWDj0WjtBbWd/6z3PHMyFVJccyduXvb4xlelfkVZ7KH4yA
KK6bAMUz+IWmY/+UPAaJSVf/RBfs6miWj8IfPJ/jTqdI/WZ7aUzniVxQH3tfwuhoLCok/M3dQ7de
cCoRP3FwPex5Xge5R5SBeSzeB22tdtgNg4UsmsBFhfOx27ziX4BU0DmcjxNtYMGiX0DOyJD6KqU8
LVNBVisruypbbxIzlyJ/SZGJMV+3OQMcmSFAs48c7yGOYNJ6BLDFSVFXLa0kSyCydYKb511jJD+T
OjSx2zvhgBUguZ68vg4Sv2EiGf8gQ0isksky1a/myI0eNaC7QeftvcCTVz2ZB0rkJBY6vzbqsDf6
lFovxNSq+13HwUl288MCeSXcGw9ad8oCj6Y1unad0Q8P0j4If3KW/wmFl8j1+SZkgYiXgiwRJd51
cimdsIDwHz76bcvrd3buyDvpT0ARiQtAAkgT27CADZ6lLW7HjqTnmcuk3uPcsUOguG7SMepw3r6R
FMpxJ/YGgUKJA7YfPlUuigaJjgcBoVFrAxyyAjuc6G2Ety7unL2HRSGFJLn/rVfLZxalVkJ/eNP2
RbRuN263ZyQ8nAFLcmXFxQjI6IKNmSV5tNR1osQwxjzHL+Tdcs/4NZlJJgRczJrZ/IbXTUeVSj26
WWyNcl/q030QlQuorYzn9PielGx/G08hwgx0zWGntKaZ92eeFEJ4oujN0PcAKTTPg/dcmR16KJJ8
ULJQZNFgqfKCehrX0Tkxr2ntdRrfsjYyM/pwD8UNoWFsdVEgNagb7uB0/gvMUvgW3xL8PKsEnsnW
fCb4l3BuMFx6+dRDC66ff/9ipL50fctH7lyMFEY8gF9fMtGTfnNqmk3gWY05Y0cymP3c9+gJd6xW
sZadBhuaW0ZalP8qOWQ0QAljZsm53z7/AuOsPgm4UqmDURH7p1CrViwRD/zkC65/zuCZrt2DLhFS
kJ+HGeCemXuXDrLjYMA5ImG6V+dx9odOr9tx9Y9NqLyhmLJoWaZ/klYPX3fhnC5xAQ7j1uO/S0vb
00pGmJ5VA7RhDTJxgA282u+TqmpgDvCahFyt1tY7inxk3HgEvzeqiNvJKWiaLx9rweJS/hJNnkUT
/hp16srBQbZR6TdGjAA6VNeC8P2JzbC0Rmpbw8xvTDM49/mPtBkBzWI4rzt6/PP0p6Xgr5CHmtke
KbeToKv1qHH0vPM166ZOw2UIvZIS45n3Kvy/n/R6KKlHeRq37bW2BUR0SUve8fmUGCaEaSeG1KOn
1x+LvJXvyyI0Uj8NGmE1WuMXdj2R7e/RrH/9sLKYI8G62S2ywMcoTIfCF5AZvRufh7Hyno6j1Saw
XJ1QGwg9Q0zWptkUoi8g5u+HTFmj1XIVD8nz+BrRiaKoMOLdkn3ZClq8en9YuJX5Xv6pakBOwlTA
3k29D4OS77iX+TpFqee0x3+BQ6mx2SJaNcy+okixKcVWU6oEcizehKWU2fydKSPJIzNkvGalfC+M
g2Ou5s1Uc+uiL+G6roenAzgD7G8Wk9gXFCbz9Ef8ohB0Jc4+sfQoMZZsIVt1QOJkSBX8NV5ASyP3
FQ1vbLLJmVkyH3kgaAl5h4/4A9ivifBP2SASQQ8LOEsU846TEZt6pr/WJSxpf//yzIj5usH/y5EF
WGtOE5eWnmeneyXQtT5fTpErRxdxM7OXaK0YFKehdcbHjrDhGtD2r/c6heUEcM3MA98Pe7t88vTJ
6jpoOB72bua1BbrpJyJZdlLmaRKzcHlDZZkP8xEmKzjoCWNk6aaRRLEiz19G3D0O9BEQfJPXyc32
lrQ53KkpQBiBmZHTxW9AfEFJUwpBP0Z3oxOjjUWWnWJcL75bN7FbtsX2Dk4MvQeBDLDri5xMEuBF
XchlTD3TgjqgEdxITPGhgKdxh9lZEKzfSiFd78AJL64bg+rOhJmk2xC+2buwAJJshqdgnOcaeWSk
6n0E4N/eA3241rqzGowh9uldJh01Ei9Ldqqz7eUfpKq/zWD6NX/o3i5sAJbTZPr3DVg8md1TqzRb
PIB350/1s/lQ8dVDMtmYV5x/xrVKHAa01dKjJ5ElQIYvD1mav6E+2vP7yIQFo6i8ipeNiaLVIPMD
5kc58dBOfspFHXyWU8lzk907nvZc0DAS+pG7gVPbODuBGac41iicyl9wRCO2YayABeUbPjuaLXT8
WpvHdfDbm1tVaM7SWyynktrzWilT5L5oOKU7E200OmnY5ueco26Ul0hBXereuho9ef2+fc4ljcpK
xLvYBohoE312/AZQqNsCr03hn1ERVCjzyQYh92paewlsTSlFj9EOKdilB/jPterXSERVOr/bszBm
VqFEDQuANNVh4W6IFqKuhBn3adnfbjaALNnDlrjJhfM6lVx1QVW5LYPO9UKgLM11en5hoFmrBF3a
SE1Lofk9IjwIJUzVK1U30FhXrSaarJYY9TObSrCZxU+EminSyIld3ypwPZa/tXIGcWYOP6cN8Zld
7T6dv1dnCXoIatsurjnbxS+p1x2QGOKJ3ISmqHiMQsGjobu9EosflrL+jebie60GPSka3NF8QWRf
JXSdMPG4ArnpSGQxDDxvk9XP91Fxn/fPOni13z7tzpKAJJwS4YeH+ONnBbrywamVcvAfHxlvAOCp
1rRRXmW5Sq0KBYECRAtgO54tCvM512bFZoInJ1P9amomRWKHc2jsjqgVRwBeo0QTZI3GqPo+L8HP
5VR8Owong08vO+qvvFMwk9vh4ioKicDMjAE+fLX95sqK6oeKsnTr3mfIhCrHA7LoSPvtjMfsYys8
8b55KrnGXHHCKMWsG8uOuHKto6KmkB410hE92J46pFWnufCW7SXOl9Ujxy6sIq9CIeqAQdzDdhT2
qJb+o/k20IURCAzCphNSfr5IqPa/0zvMY1ZHGMqDeFZG+lt0Dy7nWwXNKdKsB1VU1/qcbGL65iJz
7S3pKLRN5mYDMc4oPQojgTRYaYtbdz9+6bF8D9hbrI9mQNsrjgTKUgEsYDMndz2zq7LJ1Rp5t7x9
m+ISrnnH9a9oMVVl8o0kI9Bo1lSgoYoiTwvG5G78e9lXcjB0UpnJgu2pAObmbr/qD97IjruYsazl
eDIt4j3uUjl1Ir7CqlITg5TwSQieq+geKZYna/fIiXkHWs8mN2kPeFRMQYezhzFV/w04Vvu9IdBY
ACDc3gCDX9J8NC3x49/Om1+z1CQupFyY4Z9oHmTKQtsfBEsYq0NfNWpGtPWvhd++seUh7VxLS/tZ
8PMYi8NLUVIqSJaBjZz6zkdg4mzA1FY6Bd4QA60jnpzXlRCzhG/2z0ry+hlWQo62NSVNS5vTWEYI
2iv7PZa0J+q9zKZ9uLKDxtEYp0obIhjQc9I4yA0oCeZQn+g20cL76hjhx3R2a1RlyQyQy6ZGD71F
pJzfsyAWLZXIIS3wngYnfhYi5RK3MUyXovafYvWBQesWYyR4O5fHjQVgCBUx3K+uIMxWlLb7JEg1
sk/fiti5he9r+rpoEYXJYNOAAS9jllaWwLVFm60Pgz1Jhn8cPnBsdz9yK0z8EffNDk0eo2g0Vx54
jCGZZy5+oC81XER5xfv0sSB7H+iysLeN9lNsx2nErB3Kpmsgqt+XIx+iqpZ6/NxDOxwsi3KEXY7c
A8wo4s9c1jz+2NaAcD8NDFi6aUbdRa9tTWTRyd25UrWDThxzWBplJs0pTM673zwLqzLcZvdE0nYh
ufS21zeXl0YSkMqEPJFluCBRG+ER5C6B33jmSojIxYzARqKJ8CZBwlRsonWOWSqFbuovPprCXuHa
bcIGqAKyhlQmTGslUeZS9WvCjSQNyUNGjnganHZpw3+YmuDTgCUGJQgjNAJYzX4fP+WVN98AB9MI
OHVCIVWkNVvz7+r1js6HNwjtJaH1x4ehpg0t+5If232YApFyzVXNSi6bogwzkqeeNVteWfoCV9r9
JIozojL+x0RNUOGh16StLnIJIMQz4i6VZjNHlKH3atgq4xrDmdluV6IW81no9FG5nfNgARxSJ6sU
UoZyrDOmSxz3oN7QYMfrTc4WrlWeuHk+u24Do5cJZKS+MOKA0HcdMxfUAz7ZTUUUC9+hHJrZh1PH
cuGyeMehb6nrY3isrQzrNW8XQ+cVBcmt2cx67MEFUMLj03ESntmM84lvI+zsD2cW8nNKlR17GXzY
/sUTUUx5lCXLBVPDXw8YlNsOAnIeZYZhPXlw5u5vBw6DPkboFBqLcfDxahuQ2hGGcCF2SAkn01eb
JtG7g2byg5Qblee5Aw/2ujOI7Akc/VEBfvB/UAdZTyZ46xxNG2AXyVfU6PeZfRx/Zf2k9DLfMb4f
bVCu1iEau44atC+Xq0Sle3FbN5Iorb0Z1D5js4N1DBnQtl8yiVxB8+7cPO5DARpdNxSECPKnRHBe
wx1ymwENO23L9gF/6zJHxBoZu3zTetbzN/lcYaf9RBFV2aZuwmtMQiCypIp+SQJxKJKNnLUYzszM
QrmbFFO0GRVDcnaTt/+VCSP5LHfE9xGkeeiXBy50pDT9sDVrZnVs81iIe0CmvWvPf9YRohAobSmr
NAOthBWVCN9J0cpqlgFkws0ufpUwctgYFUndbRkRKcMvq6wSuCYEL4xKYmB8rkQcLr6zNMOYC5sO
+oV7XCDufMdUb8fGiTaIQ9zKYtbUjLd8IWD9yCcJi0uzczwv9hIeh8bBzfWX+zeUfeXCQ61zk5Br
usLsO50bQ9yws+n9r5Kof3u1yT0u3+qIHF6Pt6y2Kw+Xeg1Pmii5l1b+BdixQH2o+L9E0Sg1UJJD
HMiZez9VhNEalMH6JmV1nahPMfbHGe55hM5/6CQBMEtDA4vdXtHH01gYZnThw+Ty3XAiP8WNOjkL
X2oj8gTAO0XDdu7UUpFcZ6xQqyBF6f8SYXFJtuCOfFFNw5m3x+LXjJUuBSY8x7RP7tICXJLCxvP7
8SF+W9ggjH32wnMwgfJP0UIuEjN1PFgws8YoyIAqt+wLJ88T2xI31RtbMEjQNupFBdcAwBh0dwF0
ndJM/3hnWJdm4sF+yM/3KoO6OXYZn3Ht2+3W0RvkVbFi2IxHFDCOlSQfuncKndVbOsN13fzDf9g8
XFwaM4iPYwVzAMTyfHB4Q/f6u3jn3poVjWDyXm7ifQSeWtd9rmWJPqVzvCJ6lNa7ewXnYf/QYGRI
yuGAyP1ebXAfE99WR4R3o1nY7riyZxuA5fuEwWzrX4xs+jCeHUIOYIsrC5d+OS+2t+GLJQZfnkaW
VOX8h+/ZBNRCYaYYaPQG1Kt8ngtprjnFXb/L85M4KVP6CYVrhGBZfgSdfMUxDfhxGykRJGQPKkDq
0mpn1H+Y4Q790On4u0w+IfJcx3c/OtEqhD9OIMJJFiKCOjSaPI2ZMiu6BMZfsX/rm8H8Qd1gDAKR
BBv4f+9I5y09sh9hftUexfgfbsz9MAL+llm9qZA1SFpNWrtz4aIr1FbrFQkxUZ2CDLHdflX9yYuU
ycy1HBo1+GyENhEJoPMEDO2nZ0DmF4nhCtZPUfvOzKWg/M9dlDJ2vx7BPTasQrnsQus/Wy2ckk+q
SoBF0YEuR8Vqdx3qNDVP1Wl+tDKJnJuJ2/PA4tQd3Rutln90KMcrHZffCvQ52KvA7eYXe4Gy+jaI
w1maAKUCL/DHBIi+BVxeoWdzeI1zSGCgWyYC+VMdl0Z8gsZpv+xxVZM/D6O8kBHBIpA6MqiSPq5n
2nlnBFiwhPpgNbhrbxJFO1pHeLy2sv5SqVywjuk+tJ6yee1VNCnYsuc39lpv0incwOO4c2kNQOqx
kUAIeGFXAQ0gB06btk7jmAgUYR+uJSBIC9DnaCFQTb3t2uofHy5a/s/46Gxw2PA8eCw0BNAHTdt8
bh56QJyMU/1T18+ax8qCxadWGd3t82syuRsYcGJFaU1SB/A/7C06MfrV7ZC6WXwzAGLuSWu5v98s
x0ggsCPFHiJfYOJc28ll98mwB+mveDjwOydT2NhbBqymAww0S//v671tGpxfqiF4yYVLVt6cgx8J
qLm+sHQ2w7JA5p0WQoEQr/JZSj/ljqAh6RYxRzsXYvUhm2cXSHFl8iqK3O9Ed+X7M/Y41JqPaskE
yXnMq4GjTVOsj5S0+vQTnzvzNCXuIR5OfsboeVqNlA5HEqCiDU6nO37egbcZ8Nio83rwmmsli75L
93S9m9SZhtCF+pLylwf3J8EjV/T9L3z5rbHx6ivBsmnS8GU02kbNksb8wAKmMuDGMXA53pT//ai/
J4iOBRAHmU37X3GY2hJEx8OU0mJO9yFPBXZLVX2d2OeU4NDwr+O8Ht2Cpmn7ZuFR1VV5NuYtHLIF
xwU6wjSA9EdJ6G2Q/lWgCyT/HbhWSB4g2aWWZVNIudJ3jr8jN4qQg2ULdYjg8spuH8ZPVp3f9F1a
YVaBmC5ROs+dL+U5ZZmr0FmqWv1T4tOKl86Nas3UzTOLQChGarJo9Z7axWUa/9O0pAz4B4vcU8/k
i1faVJxvYJI4pjosUN01liYS3K1AUPWnhcnjCYUCIKn4AS2R/GvzfM0raXZ0x/AzxJeynma5Z5Pa
uH4YVZWnY+zzSQcstij763XSgph3kzjePlu7VE290/33zdMtcafGejNYIDsv1wRCG5ccIJlQuGgR
3ka/mOl4/rGXWxs8R0PgSsEjuKJHmcReuJRqOp1/NXfZF8oYT+mLorACyXkybWKI6xauo1AGfu/y
2bi6fSHFhsNB72iQlj2aswYuTgjLHllAO5uZE4EIvztfq9DVeYJDGJMe0b38M9OKMhjvd9G+RGFi
ildK8SUsgjl8jtipfVCVLXBRr77kyPusXDaennujw5LOxOKwuqzkUl4hQfQrA1LOvrocuy4b0+7e
cuigD1GYeV0OsE50N9sLEyYzCO+PfhpyIfEENgBTpqy2EGudSVUR3LRHQwCSnH/gmRx5GPRC0qQz
iutOXOQaFQydDOoIWAuQunH3NGdvrDPYqhsc+Hm7Lb7ts3VxE+LGJnr6Hqn6AeCGwPFnWBXMLT66
V0mtDSxxB9X8otgDgR6QNOIwhT+EP/XMFRpo8kAFlC0M/nolzmNPxa+tP2HB8MUgytey5N44PEBz
hYEnBsO4bPONuDjh4FatRt0w4kuA/jDHYfw90BhL2kdGrAqPSXPe1OpIvghKD2VVi6HAMHGWnSj2
7HjWpiQ2fjBUL+1/63gxjbwGIOBYIJn63K6fNeXpE3xij0DHYZ6X2XdsYkUJ9WHZqtjK4+JhDi4F
4103nCtU/147g1o4IXVezyP3BW3MCXdcH1U0/mWbHO3NU5M2xlJXC0y9W2ZqjHSHpMT1gDPvT1jI
hsJNuZrx/YFNZmjVrliEoVkfvwTWzuxc4ekQWX7Whyk8csDbpfBi8gZY+ME6CM78/25ZLuqxrcjB
8TmwMHrcVs/Z4NUljVEjhu0ETQtmgs8dUWa+09+uAhLYQP5mSRIZg94EAjpqN+MvXDUyZwMw3R7x
KFGDU2OcXrLnjgjuuPRix6itQxNpP8pDIHsNouCeEU2z05Iez30BN8ZpScG/6Q98rSOcbgDIf+Fi
VuzDNA0H1hh7iTbFYhHszNHNPrGGyrmPwVsNkuu/lur3FxyPQfm0/FBZzplyFSOn+Hx5gTYBS5o0
jKVHCAC+vB7GfOj78n3XYmZ28Jf2zEZLxBsTV4PFx0+jMAbIcVGy9qJ16LQYH9/mVIpkcwjbtrWG
KsZGYZWIb2VCm5d60s+GqW5HITaRPvv0OgPExSWTD2FVtLXbF/Tjq6JgfajOngPHzAVWCARoD9wu
yTYEPCuOpXZtwiNCL8F4Ga+9q0fmdVA2rVlG88ffuZqYBhK1ejUv3CokozN1u5QVoqNXx4rwz5I4
bermru/CFK9ccSu3qoYbxqHF5IjMkRxJtGbDuXT6BQda1QKyUJ+UQH09pK4DN9c6QjhjV/y0YzVG
8Nqw2y8C+x71IBhmEbq65q5+k59taLfAtRpmNy0OFslwmCxENmU2xHaTV9W1btMNLOtgnVy2eiI+
xYpbnS4bY/OF002bS4q+P/UhBunROYIyFn53XppFhK8y1IjBJ5ET2ES0n/SiT74op8sroL/0FzJW
LPyy0XmXIMRcI4E+i8F2uWdVxR987zoKGxAzqHibWWB+VyIXtOfDQbu+Ztfo88U4z9YPT7KRmXx1
FhBw0VpW9F+HFqCzjPMwB1y1vvIaPE5yVNDNL+lW5ofDKGSlzYuV/pkp7IoswJVDQpVt2Fu6WLqd
nhYTo3r28HyDk7qc7ln/U1n2eIgqOQFTNtDxWV3m3Ee84NrR8Pc2LpOkGqite+oz2ugmC6trMYUi
qtTt11w2cKEIFiONZ+RuKH6molGDoc40HD6EQvabatmMIkHgob7IMclwL7tUInC0Hyc4aJhO2Re1
AjvJ3QGGV0KF+WmdmyvJvwdAb82cvVztdBNpn9aklY6nK99CVHfLBFLPhYKMAnTQ+GWSafcFFp2y
7MuOdFTbE62TtQD6bz4xTW/loq3EuhyFPJCdAc0l6ZgfnIYg4c/3IaDZo46t8xnGaJto6LnX0bUh
WbFmX3Ec60RjJm/b0iC9xSp+Ze+cw3Y4IKwEk5qtrOSCkEObIjCduxXaYVdPXiMhwN6zDQCvXy40
1x8CHjKpzX7qy4QJbonfwZzIrbySYauBjXo5hn8bVlkIL/YyWhxXQ6kenG7PKpw639vF8QfCor+D
QUKrDQ6zjTd0rg/QvErdB8op2J1Gt2h51eiRRY91XieDYHe51Sz2Dm0PHt3kGTtMVJ01U0/pdXUn
b3dPkPy+fz2ETLUTNgLJfXc8KKQ6RroPiSyjDG22vlck+S8VJ3dKqqZjdPaXHAdEC3zQc3lFS+y4
k4C4Pb4dAvCeL2J9T9DeBs0XDRWLPi7+6JXkpu3KoREIRTu+g1Yu/4uwbmopBIKZJc7bSHuHQpr7
u7Vh8sRgskazBu98ccaWqztUHlluTtawn25SLNda64NEURdh04aLNodPD+uiUjl7YDi/gXqnTzxY
IzdzdieAEprHz8xLj9KPsFBOKNISl01XQNSa9DkM2wii48kLhVhwKe1uORQUtpL9KneIDfxs/mbA
S3+u+u0CdTg1QkdbjZE+X3XjVfkuH7Rp7DimOslCh849a4MD98FkZkh9UKL5xictFVKZOt8V69JI
rfcVtvotE53T9NpdNsuONyPztzAYMIJrJME2bFaQ+IPopuGnudcPDYSYZMo3X6JkaPPzMNFWjp5H
O8kfecWR1UAJHTAnGsEHyiipbYXHHMRvzSzpTmJwQ+CR+E/+bp0s4t2HPFUbqahYfXhNm+eUjoKq
n/xXQ9s9aJ/ASG67XTltZ5yI3MKQLPwC2oPWjGwGFH+esYNk/DrKowLuocuwwidolYGrSf+5TgvQ
hfi/hIKwD+lobhZFwnKY5CqEw0KvK3BUrv/XzzsiJtJHZ2yXJsCsg66VnIPzm2TSS5B1uuNXyQxO
xPJBptvlU3ZeEt3NvSf4r2TmjIuGUCjx8FmFYdB6EmRYhs6vXlfl3r76i4lEXQyKW3ISUPMNVe8x
owPn0h13IoHghDgNVsdrhwO+p2LSNU7qZzjRxRI+eTfNTpCY7xDHvtcg60F8vEBr1QUIJBpPLapb
sTZRZ9xueZvEMba4l0QV6cW6LH2wBUXoxrQgCSRO0mnMbgKF6hVvUM7TkHXwTtcKXKC/8wtRxNqT
rPDhyN60Gb/rPTYU2N6LNA5fId3tPcAL3vfh2/HrgUzuYefUAbcLmFQP+bba6U6o4Npe7yBaGrvG
qTTQZRbKHXx35y+iKHS1srWg6ZORIN0pycggb3Cqu9+ZpuFxTvYySSCbbl4sH40EtI3EHEclFRzn
SClf1g6S00jSSX0rb1vnnu4dftnSpfwceXFJphtsw/hqiOJFg99mmy+AEQ9Df6XpGyssJKB4uBfb
2/OtRE7E5vpGQLwJ02eJqrmSHUkoUmctqX27yGk/t1Zza6BuCvXZLb6JsRqRyCdHPRhlSORs9k7a
DatBshG5Yydzfka/0UZnvdd/sQt9IZr218Eqh/nMrWHLpnKb9tQDTQnCx81ABV99qAzp+f2KTEr5
zJIkedmSPjQZyb1QpGJ+WXyt2LVwxZ9wKr78uVztXAacx+obB/RLp6QqbxxSQs5qwW8AoxB+bxRT
iKhlFKGItKDpf048P4030dnU0RkOZJ08dYAq3IesIjiqvYgo55LBFI69v1WYz35XtqsnCRQAHuOw
f5VLkxZV2ZrZblAro5MGuc+h/KU5y3RN5cscEp3a0YF3qJRbi0/abA3KZU0+uClgH0XovddSWkU5
NOJYbzkcjGHYsIdwf0+ObG//qr72CbtvayqQFa5sDBu1vmEC2swfYYi3qlDc8hCtKHmvl9v0I9yd
vUhD0g1rRQI4DQwSaTYu3bAI1yE2fLZ/qEGttTSFF4hH22p4BAPlNkl1fw2TyMB77TvKojkdsgcJ
jttSfTUooDwSe9VRhKlHk6vEf0rbJLQVGX0C1adiaRcM1IBVQtBFIOHjBfFyIu/cKdrOr25ioiEU
UKy+6XGgg8LmzQszU4vFstqqGvhF7bGCgpj+OPxprY5LP83OPskpwqMapi3OiEy9eYmQnlCPY/wF
nVZ6pf+a4OhUmpXt/n1VVVNm4E1nPVu3aUS+XzoihITNXghYMCRSAycYcYl6Pb56KLdKPeOLBfLH
x7XVJDbNDMuLB2kL2Q229m1rF8e8Jj6sb8+bdvWkAToxHuB6vqUSdrtIrys+vfUT1E1Pi3JDgIH9
DqRW+ANuZnQkTKAfvZg/5Dso7us4n93KirHjD6W5mVOF0Zd3ReqC/1ea+V67q8zQo+hFg97eGBes
DK/aZmqx5ry3JZbxribKI3RNY4Wx3TXFWZWBd7VbNLzfLA/bOm/ibqvcV3tYezCe+91k2ov5/nMN
oDfJ6fwoIhuSYjvzkPTL2519+a2CTamIbHnr+zX8EJQMRPszg9nEMEhyOe22GU9NoEKuSX5UQauN
5ClH87xYAP9akMRa77JElb4FboBQfL/wzC6sf6vhZnSbaZiWtYMjSXfx+vE1Ly//BcRt6pQWGKTj
Rn/5Lx6KoYJw3mgpsn/ksaO0iwIJZGedDZXWsGUychFmkVLwKatkk9jQkpgMdszwWz+rGDFN81y2
/e9ANkXbuqnbPQtviHu1sAvFzedY1VoZG+Nt7KSxUTfw4u2v3CZ44AkFaNUZyATDIgeVy5IJQDKT
036QvW4fr5gMiVZw450Sfkq+WBhz4LmlW1V7yP2rsQtPbFVnNXnlec53563O9x/g+FSd4Ul4B/uj
f8LkJA/vupa+BJD0QpoaLBY/2ss2L47Xz4PEd5i/oBx+Wd6yHVJztU0/v32UovsFQcpFGnW87ePU
JyHGngLWS9cpWoqcvNg7HIWjR8ixBnI9lRcRHy0szj/5jNgGVN+wguG9iKB5PK6dVogLAPhEl3o0
h4g/djWiBlJYKBgNRh1WRcjk36Cxvy7RqHrJw+q3sFlhal4vIGIrjy6byi+ss2q5ouDsvmFtKYaD
PzFCmAUbPSyHGQg9136XN5hQ55vnIbBFy1bUAS44Penjqwk+bdMVkwGKrqqK5KrmlRu5cvMhjggh
76FA/clgdQA3mrUqirroWVDNLR8/Bfbl8Ggxs/1eIC6zFawFAEBMTtFqKp+lXpu6NvT5o6mcjG4x
AH9/Q11FoeNMXhEiF9KOuGsaWFd2GxmFR1fb2skAnIfXtCswuXYukU/jXOqfP0fuQSFdY4C0eij6
OZtzwE5w7g40uNpP8WJdhJdCrGAs1EzOqkypyjp0r5Dr7u2mEVKcbTirvk0fI/7GFeq81yhzsQuT
CRPGHQGSmCHhENJRiyFvKmLyRWr10xPju73iRh72oDEaGYYzWjXjOOHZhH4TrmN9xVSbQCYPK07b
krQKYICYmjzbcjJ2hOs0dL1nak1Sv0xPOP9myVSzZK3WFsk/bBmy1D1bKQY95/kL5n3r9UeH13rG
clT4DFk69ZDaRXmOWtuACg4J1hXvtRi2Byq0u+IkxyaRsBVEs+8jBTnGcNUpOwrgAtHfWkXm0+/n
ZGNzzXCFnDiaPzUwKE4dvroJG/BTHLMGhp+YlKo6GbfgDL/7pEtGSEqisRgsWBrYycR0NGVnIxY0
YXYrnR8XGB7TD5EOJbp5JuCffxk3OPBAlas7PLliButoYDZgKwuNlgf6/59NxaXQKrXkwAEgMUJw
LXgX+VTfdu0nQbpW6zKH/3DaXT9Crqh5qTFsFm+cMw6Pn8e2Kyp+YYjukUdw/eWV9gGyVqgJkYcR
JqROGlBl4AzzOs8NZUk2D0vTiwZeA05MSfm7AE45JEHmY78+ekDDnuSnDqp6Cb8pC+pGzZT2ptnK
7NsYsY7fJttywWDFonfFYHCOTSbfS2VeZBW964mUkN+DOp2RX1dQk+AO0qGoVoMnzGFzcmK6cUKe
e7aJnkjSzMFsLbHe4FDuDJCm3zKN46SQsGwUyDxwWly61Vn8mqcmfBz3i0+WRg7C+LgOSvUydFfb
IX55i0BNM/fewClgSo+W04PH2mas1ExaMmhGW6qeVcHQooYWsh1de+EO8zzuEPmuEczL8yxOy/uc
VktxJ32nj+oHBn8iVug1spDSRGmwoI1jLDYfaBu1ZkSk72l19Kl7Oi2DuFnS20iS2DleZa9vT1Km
iq1h88lt2Ttg5drJmUShp5FxhlxKS+UoTT6SPC/FSoSYAUsAhUgujsOF6sNlwlZEYmtwJ192rfK3
eZYpAH12fNXdc+yOsUka2rY3pscTT3INhnHyDmd8BDt1cK/gydU1/ALgBzpFVbTYtUBQqJha/Oqo
8QLzQBPKfKWVerGaDd0UCdp+Zr+J4yeq1JwpS3wre0hQapZxFeVXvYE0WcWPoIwfAce0g/WzCfQU
ZYQ5dXFf9O+cWnwbffJkdC4KMHasAagMx5CjMa1FTDnwQovNdOFpKVNigSw9xJpqg7gcBSv/aKF6
9DV87UYpSg5Ns+C26oKmC73NzeJi6IbrzLGNLsPI2iTgCuyKo6pldWCd3z9B5VoaqQ9G2Kwm7ttp
0zmjFKP1p37UqrTbhcl83QRWIQ9I5o/Wc+n1tdabDWtaIJZvMA8NsfQo/0nTLcX3Cq+clsmsCnmm
RKbVOVXJphKKaAEnvTyTq8DOLm9TKZ1Fbb2DkdSQg/4qKlGB3gEVq2Sqvx8HlkK259LpRs0st3pm
RAS+rIvW4gu6bCh1PnH2QpcurAebTjkCKI6btKMFnmI7lByrfaUx6UYTh0mXSj8qYvcV+20lQy1s
gjF7FdfIFfq8x9ICalZdIVcKdBTYZStaenLoFnwqU3lKWNazju4kDGlqRW2M/kfaJeU3BN0OD8o5
UMkoWaxUNG6qqTYbN2hIaiPBS6DcD67lsW1//r2+90kDifMsVlELb80xnkyY/UewDM/w82cua1jS
xxHg1uM1/38G53CtQXMYmVYuooKQFEJm9rT2G/LlSyGoGQ81+W2xbzOITqfGKEeoVvaSZuwxMN6/
K+OCq411J2ZHq6DwdkH8Ufz9tZtQrgtJeOuaDw165564S152qVqR+edSJCJ8e+D4xhublPEoUZRD
/jiZO1A3J+Ebd8/XpKcA3gEQeXPGbdrlJQqhJANxHK/KHYkCbMuR+VYx0IaugSsSEfmCp6w1lmIa
6q19m6oVsghXGRF2ceRG//5DSCv3STIDheTQAhRVC1HT8wdtMcS7/kAdHOiFnoUx7EJ+92vePZot
KuSyCIk03ZXDef9Z0l9LnapbxoVGV6t60nljAV/hgdpPpI9DukNzyDCk1Vc2vpt6GlSMK6WNY8zg
Hp+xX3O4WZQdGvQqs5AW9tKTlFIZAvynL50ZKqt+3UOl/sKi+HGeOkb6V+fjEuW2Ym/15pmNpDBm
xxfcyp50HQlfhR9ct0jjnI/aK9F2xEXl5jWbxgUIzIbZcjz/XV6TPD1dsVEDsVXP8WmHFo4EWaOR
iZem5C8+12Fh3XevrX0Zy0s6rzRph4o/+ACVThS4418WF3jKt8p0+6RNaSeDUm73OgAnNzqso4BT
j0CKRZPLPT3TkUsjYR3DqB+YUNfBtTU3493K/p9ypMQidO00c687bQF4tKRPi2SwiQLT9SRkRJJJ
PwMlokGJcUkCLgTYb6+uq/1hFo3h8X5gWPmqyDvU7M0njpptNYFgsCJtaxW4S8iwypH9vY88toil
Q6W0s1jkKavuw0aB/IgqgIUaMonCucFJKnFTZ4h40d+ItpQJzSX7QJZl3RHDcFtCn77veu+usmnM
cE0YPugXWomZVLpTehwOecKJWJA0h116Om2atjphHwfftyuUmIVK8Navumu1/nbtv33z3/zWU08/
YweZjkLLL3cbkTYJfX1K5EtaaLXpyc/dm7mXAlqu3t5zWAOcmKERHg7WBLAGXbUCDGygDS4Y8hKE
hyTeJitzkqMNy7yDQni0T2TWstXFLZCQxlxQBNnDtOV02BMWt8H+LKZGwZ9mpYFFsNgVbUdSTrXD
VFPdrohg/Pg1U381E94oiIcjH+wCtHjgCDkm7c5WDVBl2iTaPR1E/nXiBw86hLnJY95SrMXInHMl
9qUUyQfvlooXnTwcwOGkfYO3StvimvwtkxBjIhdtl5KZSjyHnVKEWukBOms41ZHcF40dR4pT641F
ygMS/F1QXn8lNByHD6+SsVikT7ZQZpu+yF0bT8tW9XtdxDAtJ5D7WUD6h7xrJj1eVlo8TEw5Opr9
6AmSJpsGbuPfA8AtVIkfpG0sWVghfKUpptAKCRhFYtvFm3GPdY4zGRfzetPfupjsntOnhSOI0wj6
M5OFMxsx69KfZDTIXSU9Gk9XAZPiD0VQjjGi2Eyqmlk0xsVgYZabeQmb2bQSxhUoIQ6q9y05OTAq
LPaTfRe92vsot1BN/ZxxKQUtDf4TOyNZRp2sQyHXo5RJSfj97jIO7REmJJBGUG+DfaS2pbmB7fvn
mDfNKBZxJpxbveqRcKuTCRKDVUirGa7wv/NsGAORxLBPBD4/LhftwMn39hIC7FwYxX45G+0twhC9
JxiOt1wNveTBzKMFfBUYrtpl7ymTDXfQpNusRkhfFtrQb06OngGSasXqdHpQrrDZu3bdCVx/LbFC
zOWqLuNFXhjYOhRZhIX5Bk4t1W0A1N+4QJ/dOTf3t9HaOKFDhLS9eFuN8ok35A5Tmhmo4H13GFVL
Jj4V7/hu45k2Y5ytee0u38O0eY8JA3sIN4/AYfPYeaTPA9Vh9XQHpwHufCXF21CkVXrYNheXTJHG
8+pWAVyaAHywBdvsbtOKMepp1QC/uwLh8/HKlb2Rw5BfyLQIKTX9itf6gjnGTcHCbdFNI/xMoIBY
K2GOMzBy8aLqzTkFyTUF+Sc5MOihlhSFTbJHIQx/XorRk1XaSKQ1wnvjvR8Riat2JVjzuKXHODxn
utU0jGh59JAWanVJfQhkEEe/onwV3Xxn8jdivCE8hKvLll+lis+DDSDP3t0LF78c2McnUtnZZtNL
kk9+w7w347TGx4Mbtzpm85qI/vSdecC1lY5spE4XAm5OzJcTsbJHelJ0WSAarn3dQWMJL/27ckpq
unCyy5jZhK+Thv+NVtaDCgdbwX0CrwqLbNtzndVTwndOjGlZzSd7g1rPYGflZaCJ+Q2iuETauDP+
1ZZcA/05NaOlVbBQwMXNIk9VRrAxR+yWiApuJ+5t0oXu+r6gztvFEh8SbFzUvYSuLhzFQKH2vZHj
7o2/Nh1eUJR7mH3a8ZemguW9x/fIeY86svqppCkjI5XBhqCYw0RmOGqxVbMaOWavCi6qyVFPZqMY
xvvzRQcwXMoh/y1GX8TIS/wRQPHVXcM1I04IBtwQEhjJ2egxhJ2X8oRCMVY+KBmMtpi99M/GwQ/V
z71XwwObjGWEa09zsf7Z+7H8LhjSSeJ3EPe1v9xyNw/CfaLCFUVIVGXybTkMPfvmSGuszufwcjYa
ev+BcvJjz7/ZjLm3BXDLA2xbGB9dTp3j/5IVSE37BX5BkHMbn8M0oCDOz6O/PqsTISqEr0G967H4
c3/RYbmTeB2YXWkES2vHPI58kiw3tjpr1CdqrIKlm+uQueXatcSGGP79ELCYNz4YQMhhx3Kw1y8T
LV6vSGPP9hGj8T9/oJ87WZ5wFAoqlz/gR1i0epmeK/pORd8ljHIdQZVICP/uDsfI2vgeCX1Ua275
PGSWiqk/S05DYWsFkAA4sNJ0xJ2WVp5G5BHo1mP2EILXoJH0hHpRt8iMDdH9K2KIeqz9FxCUJqTI
fFJtHj0MSbvh3KdAIflMgkB/jvrfRuSAygbphcxoy1WzBlbhhGvWO3JXDLxrG7Ky5VmLmkuSIdiV
8cWpU705rPNNRWdjlHv20jGnQD5+mxbDPb7t/3J8u+AZFahRORvedSCcW0iyEsAiax/A0irD0gyl
e+vRqwvbyfGl386sTbk0RTTX0HX7k56ECwRtxGLfn1bEbLioTnYrwMfC0wnVUnflIu3unIn21zI9
rIAACJzyLV4ddXtVvJB4GHkgT/pfWkHBNT3w4scaxHe3W3ize9MHyNjpbOT2bClt9Z9nOfgZz/Fw
XkQccbhYWKBMywAiURJwYl59AdXmaM1f6a5tz1ynIouhdeTkpd8BAtoo40onV/uqVbwR5DVwUF1w
EJUS3WkLbpNwpsO5OMmeMTCrv2coelMMLFptmVG5wNaMTJH6XF9t+o0wrw0mfvsB0xDa7qjAmRSR
s/d7Bt+MxyZ06yRNjEuB2/nuDxj9AIkVrAEEDIgruoVq+K979xEtifO+zkw+K32Sp87hgGmINEFo
4+3hhj0eH/wCKms0mrhu3kiGX5hVKTN0OkcSz4VidosbcfzM4u0VGQwTssb8E+vq6buJFP7k4kin
bPO5DfDELEoVztzjDnrsxdZ6Mw4XHxh6QguMHkv30EuMBTEsqM7IJwP06zSYIr6F4KyUex9nWVkn
oIOiyX1qWXdiUwdAy/wlXjHHUs8o3ZSDgfi0UEg5ubAKbL/DAgGo0jGlj+13NhfywOOmkCicbrqh
A2IxdvQd4ZDvBuBBFy+M6XWJYPIaAXLTRKiWQ2MK/gIP+FHobhSKj3QRdbps9yEgoXx0qaFieB6C
y1SvaM4xBgPNBIa+fgQX0uL5RLBtzrU51lyEil1WdCAuTON/IoPgJAzhAt+plRKhfV/lcNfKXTQy
mX9HHpxs/QNz2MfsXE3jiRnZ9op+bNdq0D0IVHc09YR58PF9bMFmxSJWNb4QHouU7Ouw7LRCS13N
CKgcPoUDp1yB6CIzSTrnhsc15elXUNxQNwwkCEt32G24zZvHBMZF9QTz1xBTly375gUOyBDpDnoB
bosQgM4JAt6uLm017GBGDX99NKOwtV74Ed29EVpcwz0sW1LKlSi4G+p3AjuAG5u+haZPwftrQare
wGbug5qyDFFd9WdpdHXPoD2YJUfVKwXSlodZsD+RQgX9iuLjZ5UWN3tIL6CV97D5T0hDfRtoBZ+G
xmmQ3G2BVWJ6VG/km0TdISnolCG89JwMYz+VKP3G3Vusg/fN0ytYLSHSFB4QodBJxAEVW347NZpS
UL371fabwG+fL8ivbopwGAC3kWZNUMy7jWkvbZVZqXVDQXAD+kaWWa508+u55RPb4dgvDJGr4YE4
W39A/MrR876UDfKBuT9xFdjvZc0GX8BRJ4Bur/WyXZgEUXkXbpXhNQWwF4/2njkns9EuxodLDQ0X
uAwPNzqU0A1qLhCU9vBibv0tX2wu7wySKDlOp916ji95BP1kS3leSbZh63hCaDFUAawwXQQWU3e7
nOOP5KdPCYtt6YwTuKuFgqsB0hyOdoxomN16fjdnRR8avUvdAHA83TQSjmiUHWWu+oENIqmeS7WQ
EPfLTO+fvGo19rFWTswUY6Vt1XKvVxULzP8mXF7tYz1B4YgxhDrE2AXkZhMZKtGHN9vX6puCj1VG
ewP2iWPboM2qCrCTSsPzOU40qt69wN1KRa3UBb4C9CSHuAFI3c8wOCS7AsTuU3A9/mhZEE85eFhn
uOn5Tao71meQiz39j/5dohmFExhK999uofqADStFKgSaG2xCr/es9fQTVmPv6aZ1UJneexdKIUBH
FNyoyTOAYLZ7D9PSyeLCrGtEpEZupFa4WBCZt/AVkF8pDotaJmFTR96LbcnblaLgSHstvXh6SKsW
zomYD3vr0IEGxRYy/WnWJ/rr5GSUK9tOli/U9NZxnwiVstCF6czRW6xp9TvIiS93MjKIIkPddZQi
H5aPq30VZNAmMVIqTtWIfPlgH2V9dblwV0dvxWUA8sjuIEFCATIOqKS0qIgxlt83SZwIOZZk20dR
Qo58XEhN574NR2cd5hXrGcyp4468xwDvDfq2zi17+LZZuTohgaF3jwLNLoWqzz4C+NWf0TzpdJVQ
RLLEU9hAwIRZDIdjQO9mssrntXBIxNE1zKuNUfS6MoFKU6Xwq11B0/NVV4M0zGGfTc68BaaKW3Su
wwHXM4OAq8EKrf6GWyG5pRf4KTMQfho7A70Q+vJdY19VVHiHM2/Wn0hexG80Io4nCLqby/U76KU1
eGZyZOpL7RQcVmC82Efl7yAtIQetx1PrasPMt5xEEIUFS05EWLQl1TUGVS0RB+gRY1ZpsQtLxHCD
WzOtsLD5HZ+5WmCeJBSX71AYIPnMCCFaDPmOaNZrxYR4HeO35LLLCnuEOYETLyHuFiWDVq1R4y+/
5Gl5apIbVXOlvhKYs9Idw6c5DvWB0qi9Xlzfhu457fZ7YmFK0+1RwJQtCLMjGt5U/YjaCOjAqHbN
v+zB6+u8rgeVwePBibnWA9jWh9eWn+ZfV7uLpaz+Pybui66JluskJbXXH8kzvC3kANN8LP+oJUau
65f+42HKQtge8EEeiyIaA51mZ18MT9hEyM5NzCCuqqVQpcVM/uJLNdWw4Q9djEiB2syhfL6FtjII
tlIlG8ZCWZNiZKnQzrFJVsLemRnhyNnoH+wBgtfYWkshJxfYNBtGKBM0dX62CuJKOOQH1Yh3CoM3
Vu08X630ob3mVqA0ko0+baPR8f5gJoqXlXvlQokWm7B8oZExF9EVOU9jM/yPfnPxSCIckBnHEolr
kxt3zvYbGnA1/cUG+fw4g/Q50VeJ337peWaZturrIWGl5DrnVr6v/NFVZhO4g+sfv16hhj0GxIf9
fp/8RIqZTiO5zaEsP045ASaJrNd7N8jnsKekI7Iz2gXYsGFWUVEqrdzlFZPQkI6BeEAcWeKu4hX7
no9JqPqQmWiY7l24TnzZwoox8ReA/uvytZwmzqtufhoWeWwfyLN4S8owUbogyw/GVAGj7X+UkO5v
SoMfW4+++k5TIWjxk9xODe92ML9TvrwbmPvd1yV45SVEqkDwB4JhbnC1OHq8n7pME9Z+w6V1CU8Y
tE0G2rIv+qjFH2dVjUbomqbOVdL9360HM8rsyUVJOKn2VecqHNRsxM01gypg7fO3gf0Ro7NRySZ7
FudQ+hNY1SLwOaX21+WeXvjoOxVTePDGxZY/GIhKPIM9AtTz5dyK8gM/iTk76P5PSqiV1XerDtOL
9QOOyFg6wjUZpguZKlZJphgqOGBWAPeODAcK/7aJ3QZ4PPskf+mUnyprt/+W/UIjNR6Vr3/Hmdo6
Zcd05hNx0iPcHlGu01SXOAzI2HZVBSW7Uyw1lCvAFdOwCQ21zHJKY9hTKyS7ExLlFmIqVpqUNC0m
lkjj/CVKhCOkptAAnU+NzfspAruZZZpqXk+P+Ym/Hp6Geijx1HWSoOlRwOOH22WAhzYlmmH6RjW1
pUonmdmGNWtQuhXhj/+StSbynZVqvvxdaMcS0DLTfDppz05aNPSx5j+Xnr8HFudGKm/0bzWJaFFk
om5fNkjt27Z4q9LPZK2SGBFs0uu3fYhyI0Uqqgk2P/WTo47VKk3udzrmvEo3qp+8Vdal19lewtx5
kx+8ErD9qbLFU0p39ZH2VDzIfAL2SvgTxHxlbW2nxdMk6BtGERZ6GNcmVx5kCw9MwxcaJH05fSbF
Ylog4nsvYVyeJSjJKDSBIfLWaG4juh+nSq2bV6L9JLsJPqowf2wMG3EuCMcMup1QRf9FID0+vyKs
pd/9OCKZQOLuRXKQEtDEi+CAhWnjswUn5jBy7OE1ZN9DhJdxVWTFj3YdmGp2nFQIjDPVflssMWHG
pX8ZgtOLvC7Fl9Hglo8akKzCb8xaVOYVxQdqlMDHFj+x22ZDRwJseyr6h26QVf98UbymVfmRnzy2
eyQtW+R8nhCVm9Leh8ZQN2z7lvts91pIfyC7pvTDVis+Z6EjRFYjIASlFwfJh3PYQWZW+bxtdUQB
ixrFaxHgnMj783sNQ1jbolEld8tKsw/q8z+rbiqh9jOv9E94LB7fgmGfwhEAfWkYXOa6qGgavax5
SuXRvR2XS0cEaQs2N884JdZpF33DDSJxWCwyfOSycGBDiu6IueSzB4ttmjrslOv4nqIscGCGuY/x
O96/sacsoHwFJFBMcqj78yUD+FdcTrsZZflUAq7WTN2UaOiVTFV5OmBC3o2vR1aemBet7LkSd/ns
CZjBHLRZb/ZAPD4tc4CF6W0d+eeCoRW5k5P6lBw8JEF2admMhZRdTwekYaa7zKALW/YUippi7zs6
CgyHd8G4Vzm98OPUaiQXjlkzaX8I8xL89Z6gBOzynEGd07gJQYw2KvlvydkcubS4yQe+9RzRhdte
vXHxO8m+VekhFLkUrNE1dvvN4r+Soqy4DLxCYP8aJJOuMQOSXNwT0JY5PYuINMj4ppYKc9T0gjCH
jDqq2Zg1v7T3x5QKmZYMAeuylUctO0LKv2hsk9K3bjV3gPaYyfMAjRUO2Qot7kiJ/Yp/Pmk0PPMo
XFDh/hBGKOJxlho4y0t2LTSC3r3l2liDOvs9R9ckB8Hs77w76Xeep4h2ogbRstDCjE6WMYhKr0d9
nMqrlDb6Kmnr85iwrrMSk3qCUTZ9JPCa3kCmqiPQw8NSFreK/7KzxwyxxDyfJkvH76egUQD7ZD2b
hCY+xOLVVZR6uLwMgTWi4cpiL8fua2fniTOLjJGmgR/tIs6AAAJYw8MJF+aJ6V64xAdz6Wy6nwH6
2vU9BRpa1HhI6VSjG8Ub2LwF9q6hfddAt0GVDbJ0aiQdyjInXBDKQbs70oKT5eHlk/F3vj10ykKk
spIKu4Os6REQot/FCypUCSK2icRTXyLe9fJfwGtn/uJppS55hhYgwKKIRTgvAj0BN68PZ4bl1gxJ
tpGbyGtHndezi8m/JLk42I+fYQEKtwpLnP24LqO7wH9PD44uCLsTjJLnZcBh9aAl2IMIyINdC318
ZwHymhKn86pGL8ive6/DcyLEcqJPZXDjS4zY3LJW3iQO3UMvzZFW/QN1hn2XmHTjtaEW9FYPtuId
gxAIQHxni+32mrrGCtCSoHngzFrn4Fi8+bIeA7XE7rjNFpQojvqHf9XC+W4vOcrBViScS8kR0fTD
jrp8V42HyoIGwU509O1vvd0RUTTmX81BmsoEY5+cGLZrAyo7gUgt7nULDXGYrUaVehjWT6Sd8fv/
DIksmOvNOEnU2ixlifdV2aW8/NHivL6hlvGJHw8S2PcJ5OoSKHGlc+6NVCeO70xbPck6YLUf3pbt
JRBPyJWe51bwVzOE6E4hMPsow8hrS2D4LW1nIaP85qsr3D5mFI70LH89tShDwo7RMAPyyfgt8ZTD
gl1MHI/GDTeVIpEeYp6golgjRmccGLTAGSvSbVZBzcVFjwZNrXlPxl3HCK+qDPUifB4wSwNl0Fz1
eLApFoCdj5rkXVWakZ7W6sYIvV+O0nd61ptGHvqmhq8GfMoNfYgKyMYvwgd6WVhwEMmKIdOoymFx
AO0RL8AXoNrIQAU9IC6KI+X0ExYDi40ae4oIJOh6qGaqSn6C+qS7c0YVOPRyWC80NdtOfWed3ILz
I1qM1G+h1yhAjQyOU3c5uuA/SG21ZQ0MIqJNbqPUuqBnbC0Vr5U+3yqM67bNxrIXSeW8oDdZj8t2
RH78HfpMKHcTp/aJc7yoB1q1asOjgD0IG29KYHvMqewawPdLSVYfCUlogVEdk4wMoscmbXRere+K
oX9pB7m2w7NnnQmgnqOacSlF7WLWqc+iJf3moqKrABgZqhVjuOr3I/Opc9MW61YH46yv5n9KxAm0
xdwfwmWaiUJGqfc2Q0aN3xtKXkIo//Q+P5AqxDpWREOzXHJenu7mJAa0bBHodEqXU6wgIlXCWciP
Kjbvlla+t0To8bbSMehSofBWMUxFJAX3I0bcTrpXzDAU6HzdkGVttVM0Ii8mxmse/IcRwB0iiHwM
borh9uV1Om+IICsgpNJfIQ6LeEqwEHr4uDCvXS8hymD9OhJ+bkWbPPbnlW5aEl8fOT0+MngKtF+A
K36oE/4TlajgTtyBC6ByHn4zy79RsJ0SrFyKUlS80sUuWxyHdYwRLp2RMFmvoIsE5Kr5KJTSWP5M
oysJ1d8oS1+rwtCyEvI/ssVpfbWd9PLBlVQQEFEL5LijOotsqIAcqe5eEXYSwb967wNJooZzwOch
h2eIMLNnTp+YuUdV2l73O7kFhLzRZJW+qV8WuJMXKYm5Azn1l6D+I2o4/LM9j8eXlhHIwuXFxsGQ
3LCNMa3lT61SukOm/l2+Xxr0KeJfaW8aJgQDxDLGtcKWTufRBBlPNqDljbGTsYzRBviaqpQMTB6S
vup+rAlj4U1QXnoV8GuyKpQ648YQSDIKpHm5M85D9qawBQDzNwwWE6WuPMfaSh2BSH5o1eeKh1qG
s66yLrNv3AvSnZ8DdYG6nPeVYJkBufDoaTRIt6ORRoozKTg7EOmMSfHxnh/44cFP/7LR1zBs8N15
/70WkMjIJ4j5m4Zhyk3PTY8suC/69HiF5O9aNurW3rc6O3QCsO/QTnwjCYtsHCMo83cwsdAA1l6e
c/diloKiGzQAbWqbuK7apqabI7/YmB7DxD6hcXltPRrAeX78IRdKromvyP3TiajWbNH7y7Wk9U90
zhdV18h81wx9ibKBiIiMbT8zPcUBo0FZOj8jKW86L0WRak63Dx1X91J+jkzCPfNVMpgOAPDeJrO5
W7o+pEF8nJj4ymngiWk1ZIm89WV4CYcTx5oNxJHzbGuh8ndf7+ZD0WuiUb+VQ5lREJc4h6P86fhP
+8nlKzC/5XVu17d2i2drZYHSNQQ9tNAe5J4fSfLHNP8m6vMWnBk/gVkJ/nQxeg9wOkpw119IvjV4
3gs61LyMl3ZhilBQYJ+VZLgAER9u4tP2jgqCc9nTJy1a5hBvbNdQ/PfNJNecBy915SSdQ6b/U6JC
ponMMyrpxTOUmDwlJqDL5LelsQ6yfM+jzuUkRjJIJWOtmkbRENVXOr01n2OfqlGRhW2bASBMw2lI
t2Fr4+ClCJkotBgCDn0TVSxQ5Y+6vqnJqAT8/Sw7aGGZZB6CMsIiC53i5jEiewAe3ApxRCXmGbmu
ss0LLbYZhJnlPEknMPsE/0FFbgibYiZfJQPuT0XUdyDT7wDkDqNT3KbNC7vSa9K3sS1vnHn7CKiQ
0y/AkpUgM0P2ZpBAqn6RXrpxERJnxIoVA8llVwq/OauQNWN4g6sogckJlUO8R9j5vQGH/q4h/OAv
/Onaayx0ecG4KEjFXlfqhyIxxbRvZIYeb/Oexrg7cVqCGwS6g+TETjcwHrG+UfirpqQB0VA6JTr+
a0E0GJiTMMT1Ia5RCTDDsDQVtToc6MwY4+KgHvMPwc0dF0c6ZaEGwW+nc3Ajz0cUD1jce0LTa0qP
0SnE42aT4cxPWovaJlDTaEgPuCsQrz1icK7w0j4eyFa6BP/RE8KDN7wWhPtKy9fFLB1PdPboLWGO
x2F3+iWWPxDA5gFaRJExa+7kvrVazaUzJg7OpUmGWaPdKJuLfU528LmHqAF+UOM8mIm2bs6MTe8y
Y7UNnFoWunDGPL/auKM+OoSJrDzNnVM3zVSBV4oegHYoN8xTmz75aFZuJHvanzaYeLHdgwOPRIS+
PtSaroePer+OC7E0zF9bgEhWJ7rK7Sy7bNm7c71H5qlgQvoM62j+KYNovdGFaOnKL46sCnqhB6it
PWZKWcyAFVNggZcohVI1/2TEs1sSyAPtNU7C2MsEaLmVzNH87aGn2jRgeI6F9hDMs3kpNt7RNT9N
AwBCR7MjJY2EQw3zt7ISp9TZBPU/c2RW65PmFUkZAIJm7wk88k9qOK6aDo6TbE4P0DNNgRt7ZknJ
9KsrUO6yePoORshJDziKy0LF/R1Bx00p/LGAd6OToRW1UHWUEtoqAkOZd11V2MM2keSNjotqFOC7
swJ4q5TsNJHdRXu7kMKgGgU18xEz0mxgFk6/non0sMCkQV54VBQnPLVLRoTM5U1Stg7GsZ1xwRrb
VvTSyTTLL3TGafXgU8R3xHMzTQkbaKt9gVZUgTqdlLUzz7e6ecoW0ACibT4DTkdLW8RmkT+QeZc+
O+SMxkyk7nNsPQwVat4obbnuggs9RuPh5aYpbuyrzQd0j4tKnNt0y8Ew0s9HEM1peBpewNHop9T0
0b7JRx48M/rlT+ciZ8TDcaTrwgEo/g7iAwPetLaD6Zk3B5Bz5BoHLVCkTe/2b56Ye9bbUyhRs5E3
k0rCjOZMkAuJCoRJOteG0I0S5IKNDoni6t+JTq8oPlgRDuhfn/V9hqX4uiGjlF6ppMmleWz1odc7
uKyf9aqskyB/OIhdFwS6362wUGiJDBR8nhZXyliVE1y9IkvS8ajHzJtI63MGA0Lp0I9Tr6BQFVGz
ZUIHp+MbBKXAdwvrCgT9Kb1w/HKDFITriwFC37zSED/hmDY53XAs/5gWwSwAJZ3DN84ZWr24bFW2
wC5cVhSfy/KwEqwpo4/z81cse/zZ9Ij/MTdgZ1hr8xt5jZWfEisFAKebX7BVu2yDnSCVOPq8LZtO
nhCf5IRONogfblpf030iIZ11KX+H/Z1d3hCVxtv/bD/frzqms0wdJvhM8+Mk+H8XfzJMSaOtzNUW
/xIdQdy7CAG+pIO/frBJf4nGDRvueXZehaR5uJQdHBxd+S1HKUXsg9yb2CBFgHdXzTGeaug3jKa9
v2/EE4dxf0mlYhvTFklsWQRnJCr4BdVNPmbFvb2ymLed1JyO/WJVBg27HUBBWFmD7iRW67X1gEYb
VuRdqBcPFgpkGSQHVSEzKplF9VCf12Kg2QAIRaFR+wP1xuY6mX1hZkJHvxfbdj4yw9buKbzsaNKH
vJh+Tk6PQ+6H0GQWndnSpyxM8PWn2scKoWa1y9A3+J9O7yS1RKjYSiPprja/Vjel9UTiQw8YcwIE
pCGthbWddb7Z13MYu5QLwZviAC3CifYy+k2eEZmlw/+xFIVcv5Rv3MHyeZ5J6NDcBixD11XiG8A3
pbcXoH3ULOFaIy3XY/XOsxnqumZRbSAnBM8UjxD6CA/ADvdFs8FL3FKbLOvA4DfvU+Y/pFHutRwQ
CUdwsSKh+A5pnfxOQfjNzXie/dXnxLlZ4k+uGDHRMj6FFNt1FvHGcfvnojR1Tm9CEKo5Z4BjjXfD
VLEIBZV62dA6nlBMbv5v+PctqqORt9f01Vc1I08iEXUmiquKwqCH5kxO1NDfUCv7gEINhwAA4zIE
UtoOLh8oNb39HOmHAs1leDXXYsxEZN++jh5f8DYE0pRC8cIO79b0c6IZeKq307HyD1Eiip1FHRoL
rlEuv2vZi6cizsxWO5nWzy8WfWS4Bu8Lt8oROTILM5BzvUY8hz6wQau2iWnhUI98ylVSa9JtaRfT
fiyz+9waBuFSgnvK8BNZwdI92hz3g398Uf96JIgnnpA6H74UHJJqr618uOApvNuLpxS4t486IGL4
SzWRVO+gYrFZ7MN8LG+fqN9Ia9kizOD8sePncJNnQBHVLMiF7pnqEhiSoMRxPrlVedPxPgLA2sZQ
4O3bg8iU5H7gEJ01WgtKuvZX5hslcplOBjNkOPENm4gVnVDj3tVgaP3NbsxEL9wALPnjs0b9HEP3
YDBWfd4vOYlpOzWdkz99/ITZzCohPFtxF/t3sey51hMU/axPlvL8sj79i2pi3q9ZYRJBJsJJNL1x
CY6CYLsdqnGMCKWqymwzWsmmlyOLYNAMgzrGQs2acno+bYeW4nS/Tg7gRG7agqWVZItSl70CJQ13
2pQvO1pYITAag/Hvdu54m+BeLbRaMMFdBoR9TKU1dykmt2Ow9sAm/yhlw7/QL1erMkpABbjb2Ooq
dZIrtAKLwm9Y2creO1uvMtUz6/XKlTH6P9Or682SR5kJKESc1UNtDqpQ0SdUG8YTXW8fpsiwTfb9
4Z1sQvaSzrpvcx5VqMHIL2yGkV+Wbtx0EYl1qXsOSkIuyTUq0wiztphhtsN+0pw12OBhXjyFCdCx
ycMkNdNpnxwPkaqTbmvR5UetYNZt52zUWnLudbZNRc8S6aSf3INRcqFh3fHBOy+ZqaNvxr0z3tZb
bQHf42Tz42cxLqudU2xoyEiUvMv1b20slO1V7a1ngh2czV4hZRyqQ7ucZ/RbTw14/7A/EHknHkyC
8iSnKKMiZJLP589nOCWztCZABgkX7bzB3WuuVsPG0QJRrdiPaq3fTXQavE/nwZweq1/xInEXhpfX
qrlJ6ulEF2FX19hiVFw0Gb8tzk9g1vybYsuAuIZ8fuKYxkau5GKpj9cI4vqfbzQtVA3+Mo7P95DJ
GAh+9ZTEvsTaaQ6Gyffdqqdyl+JUja2uwRUzCVAQIzMHuBHo9pNX5aBIiZOtJWQkczW9yEcasnaM
kOz88tNoNlRC78jbBhbyJsMgOWcv/XOVEIUBt7rVdo0j3rId0woRF7X++Dmg7DTbBy0cjMdiG8Xr
kC1oOO72/PWnW7Zxb2HaJEY3CS2NzEEEhAgFu+U91S7SYzDo3OZ6TogQBMLMSKVgQ0b3shr2Zutv
gCxDRNOuXmuzQIGcLrwfmJYEAIyU/2dx+aTJ16M2B2w/FvlYg1EdwvOAAlewvZRoJ2/YWU7HLA6h
O2nnMfNqKKbLcirzO7rFYLxNFC+MLBUtzWn0fvKR3tQ1jmdNGDL7FxnYyfBzSTXkhZVZFEAA3QUg
DX7E2fTqdu1SjKmx4e9LhD2VFmzAEs7gjl8+r90ak+oZfdrYwAhve6OujC6Mf5AjbQiWj0T+vhN3
o1BR+gs6oJXOF1vX4sAWrQbDuWWfQCQRZ8qMHaXoLK0p/+KkMQGLwOG2nzTmRW2EnZSFCswNioDC
Blrsv6RW3vHskLXHFsNWVcCOdUC4XJipbz+eDKZ1txsKlTexx/Lqm6UFMP87xMM5Gy/+8ZbM+bH+
ezHgGY2K4Z2IJqdOSOjdQSwhBrIE6KUSujuUIjsxF9NNwju7PayjAp/7v2ABACop7W8NTckzjMbU
58oZPR6tQAhGWb/5JWq4UvaJv4ncgDrMBMDqCO+DQ1w6Wx5ZBFIGCwfjGkKAmoQEn0vhYmeGcTaS
qtCyuv81P3cJclo4vwegfK09FxFEefTFv/h6wh3ZF6HP57ROWlg/np3SPQNyMeUiwPy+1Y0GBbsE
+2yjFzrsCkj27myDeOY9P7d7BiYyDK3/w+3JoJWlV5ozd83BRpBXJ0lsEEzsWSsaF3FUHo2OX3+Q
lYnil3vsFnlzqkFeBycywYD9VjK0FBW4KjXkYqOcBxjxTC9jveYomGgizx/A1gS+cIO0F6pXxqj3
/UvYICFuwJl/K1RAemMi7seHo7H48jp5LHYivMQzK58p7K9A4U5DrSGJEs2nnnfgx0bn1azp8dup
fKPhHBPB7ijoGKs7PZY0WQ/d438aYq8UIjU71qPQY3YjqT6d0tWcnxHE74tbGCcPyoRXA5asY3AU
dBnaqw6m/6WCq7TtIDHdbLwGZxep7/JvwZSCUXRKAvG0YLAhU44zDCpw9tmzIN1OI8s9SvSaCT5s
YbYIR/2S1YwvjDnRbYT92UMOw7uoJCeSzLiAhWiBts0A9EOY7m+ioKqxo2I+CAkh1LsN2n6NRNZK
9n/5crmiPK0tr+pMPm4ASvJ6UoacLC75qUDidnV9MpsoLvGTLJmK6GI8DwoHf+MjFuGKfgKCCCzx
DsTeMsmS4u3KTYKCO07ON5OI1FGWq9q1NdI0QaGycSPsNaeZJdIQwnOhiIhpH11zdBGc0fA2z8xM
X/fiQce81GzF/80h1Rb3BBoRTh2fTQF6H18AqEIQvibMsqElNLiByGzXsfAjiQLfd7vJQzgt/gsm
OCNh0IqYmryyVDN1+QznoD7lTNqEn0xAdlNNcwyPpgGjU0rpbUacu1/Y2LDAW3p4SbqHdakNoPqV
xe9SrZwzdLALhp43oeuFyk8EoaA0R3/CXYoiX3T8B0mee1LS01ZB9+V5zHo68GtHod5Bxn+bB3mx
y9Wx/vFcHJ2x/bjY2U7HPcsuymyV5SvOYx0nc1zd9Bvyba0TDP2wSk4hwd+nCajell7XZDSyMhOw
3LA0uaLXjglVBMw6/Hl/rRjekr/sZD25sQewnMZbAwBOlnEr/dbf93pEwqWQrEncd/xCT/rski5u
AJiLPNxSCDJjBoX7al95kGTibZce4PFhXGRhWBe2CU1JnnWRJ9TuOX2N1bsab/iedjqzzwiS2VD4
+O/gVoExuIqmdR3QNwVVBr5J0ADk/eSIZpRprO9GncrATQiHevyVRUeVM3N8XmTy0a9EPqEVfArr
Tek6TspaOO0SO8bfhIEgSg78/rltF95J38x5Y868m7uU9gcUrRZS0D78bkxvM6w4mn0D0/MJmB8K
I8+KYHVG7bV9SzLo8kOYNlp0rANwV2ZHZUAYLTDEM2CIg2eMHFvQmlLoPU2wq07DxB86KwLgI0Z4
EAbuJqaIJBF7XOhuec8Pu/M9jbloRE3toMWDt7tBpwI4XBeayy7gzJiVxMuqViTILVk+799q25p3
ZSE5pbNUeZzz6btFLqbRTt5tfDraXa1mHLWn1TTrz3vJuAUiDdKqUjxk6ANga2a43n2eSO+Cd2vD
5SP9wPjMtf598HMLpopf3WMvrRHblfIUxOqYmyEubTqYiJBXTSZLy7tylHg6DyZnqwfZDb9u59oV
2Ue2tnjrenBDPcXIPFHXgwvKWl/MvNiquiB2rw7omee0ND5CLzUqQRiL2AOYRHWAfyAUtoHzozDZ
Z2RsQ07+30AaWVfwYhh3XP35BzliiobZ4DXOSN79Q9XKjOjQcYHQ97djhXSGi6SpypoJth1n2Dvl
3TdJYAuFiKplMtij3evLxPtO+eyQViDWHhqVXZ46ccxjR/MFSGkcd4uyP79jV/+eKfvJU1JrivQl
NcOwzdY1dlettT+12zzgvI5JLgtgTM1Anh5IF1zjg99rGYhTe11YimgsDVixgxtqwtXoQNf1XoQ5
7BThEa12sjA95kD4+tHlkLHqZW6/eFtGedlSwpAj7MrjoPgcKUrWPTWQd3g9tCsSRwRbVENZ/x2u
9SLjlKOwCpT1bVYMCXnupEQU4ypcTvfSqZIaEHvH/aCpFtk5aJQbNdmMcnBM5Z1Y3/HzKeyT7AAJ
wsjD9sIcpZqiFPvdC1lX/M984/8UEv4lZ2XdtXeKxEWu+wt3cfGhzJABAGmnsSBj6xX+a9GisT+/
UnTLf+MuUxc4p+6Kd9dGobaf+snQNAixJdFo9XxmuHdFWFJEgpmeIyip19E0fT5eh10Hl8zx6/Ji
ntolQJsNOPHoZ7W/jC0C1EZTwrAatggyzo+sun+6Iqb8P3yYWTuCFz76F0AVuiZqZgT0ot3851av
Z8Ia8Bsthy7ZHdioJrodXm9PlWCvAUh404quWQSr4cI8CUjhnvibRvF14/axUc+aT9DolXGrSpjx
DCzff6zE7hhEsssvzL60bhRGYswDIi4FvHXzVgeH/SCrCoEmzpVVoYp3K8TSeacojV1AhhzS9KjG
iqOG+ppeIeQ6C0nxwgIOwhFtVmTdE7aLhMMl1Mz+ShGCXgW0TdhDSEk0SbEeFYhUBVLyKqnyrxwv
jdQZQd7xKiSMEq18kn54pK6Wi5mj4Q2EJoDw51YJJ6UrtyydyXj7cWV2OaeGWccNwn6t2Y2tuplo
Mzc08NPXSlnwlrAnjIbbG6vLINOxDXQZFuSNHLhdxtD1cshRS/dsSGHAeCvey4OHkDC7E5e02/cd
iOzJoJMMQWHTfyUxl0TnRDhPl7S3foAXMmvDtevAsJAqhhUNJ+b6QJbP6M0z3PJlsFj4dkSb2YSJ
xZ7LvbZ9td6EIj3zXEJSZF4fx7nuyjhpZn5UzfRDceDaGexc5+MFMmYAZ4xFZdCIB1sGy6iHOT86
q6MDMjU4raWo7qoEU3+OyolvzKtfXVW709MbloBXR8Db1uXQIjwdbnTRgIdrJdsD/3F8Nq9+cBnR
3bbmwsx4CsseH8M2QhdoNUf7ahnVwCA02Eib8CHdTgFYbZUv8UPCekW0islIMHmt5uVw6452xzJc
iOK2U60V/6I8VPIYDrXp3WTljO2+c5qXY+SF0/SS/1FDgvsBcY/++07VDWggl9bGb1ci9qsKzzzm
V83TO5xYPwPXwHQmMd3dKPor/9AHoufgsCVzT5xBVYHFg5caoxr9fWVNk70RGfG9Q0zlkSkmS4ud
A9YlkAUQ9ocaDi9Xub6rUBWy3mPTEAR+G4c9ijhMcs1PyRMKRxLuUrUnnVBCvlVPlzvW1C7QI0dB
oKkJLsJDA6o0nfTJzpcZ+LiKH1RULZpuv5unrT3hIkVeWZa56tlIgrFbOFfEivj7u+eYzIgfM20L
ULRTekB8Z724eMFYjdTsyGvxy2alaV8rg7ZnqZc3gkNOovw7cTrfVRT0ccq2JD6sMTOwnELoahfZ
BbKLKP0wNAszTb5vyGUY1CV5t/mupDWc1cwhoA4rOAPw1oXEau7oVVIwkNAKv3jufQwTcjFQVjQs
Fkrw/WeXUQXyADDUrO4+Hc7nf1myBl+qUrk/0xdUoOWWNYY2DSxkVjDz792OGkQRF844lTK4hCPk
n4CwLPpfW1Xd0Iu+gLvYzHhbqwkr+y+VSTsafrp8/J7E3xXRLi+fKyWBrTxSRDq1wRxazqhCpa9t
1Xdpel0ShqjdY3yRGUMhnvGeiPAvrTRAbPDht/5z1XKMiWFSzxi4P0BsmRjmfa4UETetLI3xZil1
Odzzd/jYIpBJmSMdEV1uVMVA1aPH3z1NijZd2qheu6SF8ZlnTvCYF4Zm7jZtw5vydd8NE9pMshNx
lv8sUibsY7i3786cRIb3TIBc8ItAOInnRgiy3I78MCiJTSf7aVym4Qi72c0aOjS60qqbeTVbqwiA
LCaBO4T0hWb9k8GGdjtTp3BhXDS66m2ovWhi9uz5REOcyxZuklBM8yNbd5QwzX7Aec7r4eUwe0HP
xiV+4zay9LL1x5gvo7fudl/86F74k2hqDWS4Gwk42aqqbyDCa99kjxfdmCs2gKPiHH1vNorNztzE
LcKJ2Ng1sOE8DJXQi+hdXypbvjFpCopX8Z6QOcyS4gZWAO/jFcEMLV5MLBqObSySURHN8lGeYl+c
nd8XKvRaPOZXJnBwgeDBc8LUNE30VFvIF7VL7pz+LGOBmjtNQlwAOjowGKCcbXu3BptYZ49R78Zo
TpmtnzcX0+AzmYtNmOpY3Vuu2mur4oD78H/yXxQqWQcpthXVaWUfszOw80Ny3a1NtSIcVRI7QdjK
nlPBiJE3vcUA/wP0zcDUrwMroE3rh0PJz52LhGKag0dAuFY7DlZBAS7g03yf14TvzffZVw7QbeqI
gvl9hkirUYXS7J0DxgW18zWCC/xP/fzZ0CcqFTipCfnfcC5gDjJb43IUjBYhDMn2gTgHvH5jS8E6
fsdBdb+DlqRMcBtcvVvOiJhVoYHVNlep89+yB5QkRyTW182RW3RHfGC9UIlgQq9QH3KaZAl7K9oO
d/fEwU6vcz0VCGUfOtZKZff2vJYaaxF8P6bYLgTkN2vonmdWr6OAOXm0alYjD00Wmg26o1aMWYpI
ra2WmbtxE4U8vB6CguMSscNMRXlfEQ4Dp4af56Z7a2LsXK/kZY8BxuJievnyk5ApTvMpMhKeN4SM
LEwa5EDnf5fJIpmC7LbdsJ/FOaXA1ZKcMPbptJyo0gt0rCBZm2sp3wus4+yW23JApbSIz5T4Q4iW
9dg0mArctDSqRP7nvse8zluvbO2LmNazzGHahFdp/c9042kfUjjSvFtfvNMP5usTcTOW7A4Rg0Yn
w8jmfV7xt3NbYsuvctIFgJY08ctRuqWAB7T0aTC8j1vqBYAWgIaW3Wyz2IDQTVTn5Gi6cmg9HdcR
jbbL2Rh4FYaAPcxQZKa83Chot0p7kNe9z0VHG342YLWLD23fxkdIuX4YjxbrDdBLz9vgBJMKS0PW
xLCta9AhBsSpPGiGFzRj1OGy6bnfbJYVZbKmMY/oU4XwTkQEcf/A0BYUB7TTo6CfiEdAHlvIm+Fb
+JGVyrNwLxKuK0EjEAmPoNCOUXDjDXhl5btcYRf4Fl0FSfQJkBJNirWXqAfifBuUiRTuMjWBZxCh
6bl2RiqnHARAsby8pfqNlFSXTz7NuoYoPXVhrppQZTT7GADbvYq3fTzl1g13RXHqpPPvtsfrMPP1
2ngM2NHIycfuGjbMkGu6kyMwGRl89Xxu8KDeCWHlwOxG2lHH5cq39ReN1lWAAzUslsKFBlraxp0I
Mx8WFI4PXlHDl9MYLdzQZKTfMNsvDVjc1j5LphrK0HbWckGNyCKF0k4opiz9Ge7EhShrIT5KSx0Q
Hn8tzuU1W/2RRzc1RkJbVyUc3EU+aYqGHRR1ceA+78sAUvjcdoWHvF4V2rAaZkqguvOJgaAr0stP
URuvzrBt5T8kv41hQdyKXfvZku3mMKu8RauuVqNXm8vx86llotk4noup8jTfYri6zjWGN09Mfcwm
0pOnoh3aiVUw5JzLrGMtqgqI7uwnbaBlXAUv4r2pCe6RUkjRfcmTmtjpC7jC6RSlmKG1Sm0jkxuV
gDa7w1wOKbsC7d1Hw4aqwnAJD/AowoVjtMXrsDc2tXe5fP8dwlZqPjO5s7o12n6kbvsnrKQQkegD
vqGWyF4wIgxvWTcOWNdkdTS909Cj0IBrd8UAI7v1/388eDrItRsGwLPqsUrrA9pWXo0YYY8We0zX
T5aE9AXrWK4hO3pFihxtdh3uMeKqvDQeWhUmETcqwLrlqywm3a9Rm4lnkSvnThvTBOY/szsOevKO
tVbAP7sS/Ed4tyKmyKuKL66GdGBj8GJs2a29ycVQj3tpyCmioytg2S7tSlzyB1lSDBIsQQhNASiK
dgUi40iQzYpP+bPhGQZ46JFtEsQhmzQRQusEitoctvCaaU6O+zbRoemJMfqh+wpIwOdUMaFgxNsB
ybFJ/6iq1rEgrr5Pbxj6E626ol+rsiwe7MwzPmgpKCzE5iUBqNeXomv/H+1/L6DY4x/ney6wa2eg
BpNuEg2epNRwl4thq+GAHOL6UjVr/ZUoxdAF7TfReJW+V9RiVBl5okeAE/Fa/4Tx8ENzszJRLDSr
lfsDBgyU2kcOCp8/QD+FbnG+etgHj1A5Yy66QABJiytUcTSW0f1MahaSD74TjyLStqwt6zuJcPpO
a2CenvTvN+BXgAU3lv1pNqrOvicKHbBZ7h8SmKF4dtqOB2V6iZfcUirNri5ZOiS6ukTICoeXtotT
rpt+Ns1hrt7u3FzFMegS1Vp4btN4ci9dIJIF8vydOB+sIViKbpLx+d2fRNz145x6gNOjinICrBii
EqShsutcoWRtDmEAwFDpmsUBdp2Rn71RmmSf33VncsnlGkla91TjdIBAW0YW1WqsDY1TH6vfG8se
KLfendSApBdDTtGwSTvchNPDcJp500AwTLXgtEL372UG7tPaiFymKHjSPsWmDybpgTnJfBeQpgee
V5rWKjLw5iqcxnrzmEGstX+0Z7NSeDlFrZpzErtu3FBdiJzq21y669GfgeZR3qFI61IG4xC42Mfd
jKsZq7thcyyK2kDBd9KGRfiirX0r8MnM1hc5VJj4W1+H2/0heWmaRxVzdJHEtDsWEWWDMj/eRugW
hiQql4FnQgIPJdAYm2doAJztKvbAvF5503tQat9iU0q32xv4vucn6el7W9zUkbbwaly+R4ZYStLY
uJyOv0tBSMBglALZhXlBcdrVzlfqT0d5KNFEpU2leS8hLYJyOL/eRqCobkYDjCgl0sNN4U1e6su/
JjuMX8Hs9GXFBILZ600YW5+W/zEaIupjIbU07QJDyH3BZzG7zXN3XlfvmvDHXE7BHWAVdg0PZNqq
xSijt1nKQ7NHZhjQ38dMXVCzyY/Tmf5004qPe2fgCtO6Yf479vhmdvLwVHREv0981VY86YtBkXD/
qPGY6sDP2zCgWMG9rr1O/ih9u4zrizF7XtlqKaDNqjIiP/NJpBswG5/JfFhHIknCDKKAh62A8ERK
07rnrym3HAAzBg6RVzKBgMnr3HW5GH+3Q1ekmBXj00QzNhJfEkiY/ybj1OtwRtphCobSw/E0t+MN
tpzLhKGw9aExXMuwh40RFGu/tE9NfahGRFFwAKzjlsRJJTGd3yUUvYU6V8Ny/pWw2hATdgp3Bgxp
2K4J3xvoxQpGo/P9ctNDjlgWKqbHvtA+CYimE7e6LhXOOR1xpa5Ma9j1IGuCmOZ5TfLm2TqkuABp
qqGOkZ8ayckbY8KQ1LCxajcc1Jasq3Wr+zG1TXbUAO0WxgxAloXlFCzChR3vQwinXcLuoO+ENual
6qw4pzbgtIBNK9H2c8ck7L88j/h3nnuDutIHtwwigITwgA+XRpyxvQ0KeSdkQ+9xCfdO6s/G0Wg4
QK1SpSbIBM2rP+98QgbmWK0WEK9LcZfUdc91VkMsVN1IMaKXULc5jgf318uemX+6WJLpKLfya5k9
gnLx41AxAUP0pyHWn0G+7PeESAAYjaSX9hQJcbnYNLACIKHY5XD3qPDyD5JPnF6l0Nt/ejKYY/QE
6qGY9vkaMY6VdoF2PmV8cJLsG/fEom45wFRLMCtc/htKQ5WeOAy+6OHZb07PlT8+O24fMxVSFs2m
eQaoyOBLcemVSFeMyYRaKb/rptgKmx2G+ha2g9nVZPHhKJ+3SMVYFc91KcBnUsF55nnNwvJGg0YS
eJ+adajrfMaqy47NJNitom5nwQ+mftH8FfuKz7MmIxDqSsh6wb6wRzF5lPAyA+ldUMJ90iPKuTNr
dAxs9MnUn+EhdzAZHdoQJ1wrhDEfyyMxQ8Oo6yZMErxtgLvSfOJWWOfDSJBjau/FS+bmDXxTrWXB
UeYhXXDAW+b/fHY63gskcPpzPGjnyz1X1xa3embAMkfmVCi1GluvPkWd14dna+EL21RQSN8vlRj3
OvvGRVzoSMNvDTOZArW30hnW7Sn9OXr91961daZvz8bzHU77oIzGNep0aVSaGp2wffU7Zo0PfsCj
wT1ewEefltdo6VVefKWHuGfLdDnEpRR3NIs564JXsN3yxO6y/hdqrhG9uP4ApWVYaKVEWSq5XDH4
MWvhIbqMRN84jelBXc8Sl8CY6/13TGD71zRP35dxSjt7jgnaI/GzOXmGS/Uo3SOyYz+SyRQj7voT
x1/k7anu0tzAurPBNojPfhFNpSvmkogr4RfsSpuvHzZobb0xt7ZWDlMq0TRrmdJZ/Rk8VYKM+hwk
I3t3OcQgjuwCEaV41v9cj8LvfE+x4pUu9reWeXlfC1FRQrBfJosD3BVGcHQQUk5JyyibGb2TBMCZ
LWuvQ2KUcGR3v4YFyAGNyJJIw7k1VUTX+QmetwZoRpz/2/hRCpYF5aXCB2uyQQn41BK3WMuMe9iL
fqACGqpuYkYQyfXFoWrqKZi2l7NnyBGEW6kY+nbb94XdYFo7lPU9H/p9H4kxT2eg250rRd6gyWFE
FJBrQtg8UuK9uKbpRUrAo73G65csH239g47ps1pn01oZkeBBns+z+GxoddGPXWPf2Qzbh8n9AjYN
S0xtU/32MeO79tI9l7ZO3sZCkVkK13NFjnxYp6CUtVF8G3vRc1PUeMIsJfJvmk6V6XWIfhgmMg2K
NE61yHikVj9jAVDuyvkanNrB8rE2g82zedxOtKs9Ps8sNadGfVKj02pADAFDj2i+CdaBPdHUnDIl
RpYFkbK9G9dBe1tYbbCravR21Cy0LK1wWD4Cw86zmkADRMcOgAMUGBfDTEgXQf9X3hYCiZ1Y4Hjo
lneeYxxTH6R7Kg681fYlq0roTn+zwb0A2F6xMUjE+PQxWLWiK8rog0K88CBOmccDuxdmY4a1Zv6d
IbV405tQu5pMS+NRr0rhWmuIhjqj815hIzBisRnvIWHUXIpracj6Mz51v2mNvYwqvvdzc6Z2E/Q/
n3h4x8yPis9eV3fVlnxqnsu4Sd85/Y/Ft9Z0ksY1M5B3lnZMpL1rYSJKpspKgiu/0g2nDlryfIIN
IGd5y7aGoL0S0A32xXb1Qh7gjvT6dp3bCOSLVr4P2K9dxQ+q/xSPXx+6x47JCgZa+jF34J7Tw9sB
aU9YoCuUtqAvM+zDp57GHE5OOf3++fsXR0WQw0OJiYE2/TzgionTmPeTiIFCOxz8sj+Xc972nyE9
sxsaVRbd0UG4k3sG+woHp7HsFhPk1q9BDfVdBvjJCwBj1nTjwNxckXOkDu8Dk9ZuH/abc3UxnjH5
B2X9cWqvRx6rpC4IknlaeHhfAgtT1P5LcJFOm9cK66Y5ctsyHCG26ynG00sFyl4+3wsfuIh/dyKa
MVq3pJDZF6z5iiyDcrQ/dBc6uIpWZv00ozAp4EeazaTd4eAjSban96wFVL6kTWNEs/iTRQPxIcSp
u6FPaxxllyOeawZF+QL6FrD1YCCz2f03zSg5Ysa/RIZAqXlF3wpLwLPK00Og3t3YAG9fFIVy3bdd
Y0bgqxWrpNLsp+NNfF15+B2GRC5u3fCQ/ESkwjag+GLp4xy10F0nHzeIC1UpDbW3NysEhhpG+tgb
XwQbf/bQ3xBvuqaU2mJ4wp5gdTO4ZFDcORgfgS/y9nQdeaFtxEMHufAV9jIZAsC07oUYuqWK3UlR
I/OUPVpNT3FShjzb2UEThFufIlMu63pfhU9UDCiCwAHx6UP9K0StZTq5cYyOIep0wcNKluvt8mPR
Zg6FosMRCf4zghPnZ/ISuiQGbxg1C9Q9lqycofd2gh8zqySUykc9PWqb3CO3nWdJVE3X3XPO64+C
wAmcjzU6LuR8QboHPob07V8E12qryuRf9jMOFG7/e3r7ZCbo+RCme+tUu/g4GCUpv7I4ObvBGE9i
Ia03CRHLV3CiEPy5H2QGD7fHHI4mM31QDW3/0u+OLHAOJe9DSi9Vp6buH7cDEtn4facNO2Rlds3q
3q8qPauoH3BdPq0mbbDeOzy9uRw9ZFGMPMqEAtFES7QLcI8hKnw7p8mXBYr25EOHtYub8bZr0Cu2
xc2ITCFgdf6Z81oH57ZfClFF0JzgWGyIaZyco6c75X3PcszlGsqHgzfl73SP5X6jk0uQm1AZi8Os
6pbziw+oaCLE+vKt++L/sM88oNLXJW4PZumyTeV9DkBU5GX0FeVdpVna3YZUnofp9f4tYv0tWE22
OWcUZZS64lpo3QitZjUiAY6xmjWT8sr5oNueC8h7CVtEswfq1ANk3NA7/WgY6g3UAzgRSUS1Uo9V
/k8T6/uc2GxhZ8NS6Gc1JsYLAECKi31CIJ/sjl2A1cLbTByzg72wuPI+0tmBlGmDzIavATJRLWOC
bKKB3IQOqp7cQpB3qhSHORPygKZnFXc+Ccgv4xx5JxHgb0VWNGiRoN3djM9U9b4+RgP6uZsOsRmn
Ao+rCbxdz+affwGdfl4hjbGmVqopZE9irrxiJsR1SHKtDuUJuXhqYtYFV4KuSuJo1hgt+ElnNh/C
6IGKYMjWz+qtmWCk/pgaQpLkVGRZUnFcFBgRfopJLyoInKGLlKcFRVNJ1e2Q5Z3MsoQUKsvt/vQ7
f6W8iC6gdI4jfOBoNifwhLjQUdUKa0tuC06Vi78wMqeIDJhj562gaQ/VFqc/NTepZrgneeyjAAmz
QAjxSZwGsoafA4rH3Up1ph2YtZkRuhDdfN1OvSYxeUdBTgu9eq00aKemA4jHVNe0d1ycAob6bIRQ
XOa5/rJbD79juXBsQmY35pUZHdhWJLv3q28TyQt00Ag70EEC4mllhEnsbpmCh+aeYYnwB/9CUNdt
NBm9AqHrEuwr4gaFfFxs7izkwMz3bLEU63k1MvIeoASlFl7+BWv6vkMWhO8FF8EoNOjvSFFs1HP8
1dNTPntkxn5aBtW1QcpF0buffYsge0/WOnKCRjl6F8xJAhj2V08KDJJAJfe0VtkE79fuaM0HBywC
7lSVfRmwo/uFages0h3ldy9eC1jvVSBsxyC7n/TcgJW6MeqVuAql8DwSwVIYRtWr3nGLULnHKTZv
tmmXYDeQEKo2Sz0gWl/+EZHJXSOx0NqxfTAzpOTtCK8oCz2N5lDiEA9N+B0DtX/Hq2AwMs/4iXQT
Zkithh8x7gtTOnNt7PE4Fws62tGTgi9OaAvzR+jVcoonwQeI9BLQ3xGWZQ4G4IbPnFJQOAtNxZPr
0tn8tPsHs7lmxU5tHtvHh+VuH+xjneOF9V5kDlZSclrrkGHKY1FK96A/sDy0+BTTG5ngt7IdW9HD
Rq3lMF04//OaE9pXYlzjR+JBdtmUfJA3RQ7Aly02yOpLBkGttDnlTx/5zRQ579XS/vkMvcDMgD5c
h54PysVVthVEPaYOYfLfwombc2LZ/LaLXqPBP7vtA0LptbYbTlED9J+3vI1+b2Dqt/wsj/Hxb2vV
lmluPjQyVzvBM2d05OrbQ7ok0zWZljDrfahWU34KlNx5Qx2dsNNfd6YK0TFxH7fCvCM9oLQxn67i
4/U517OyNUL6Y0XZ7UlQWoJ6BACrbJMpT/RVz0DhLRJ5fGHkkLJp7ZmXboQlYJNXCNLAPj+seij4
NA05ePNjPa1Zzxe6zkY5kIQE4yXoNo6opjZCz1NWB9wBe5KM6u3CYyFG0dt5Zs39HH+RzvnmNkda
srxATM90FuvcjjKoZo+9YQW8h2OVX4VLQKGuZxOV9rU/9tD7hWSiikxXK/P3LLD+BTTiUFfS1hNk
ww8RV07+EUTFjtg5toqHQ7RAY9yxA4XnceAcPe5UPtz+FStLRLqDY0/HQyS8WYtYncoPV5CwQA0B
bVaDiHEwHqL6Pu0/xrUbHwXoGjswF2TSmVeBogOzZI0OAF5bCohu7TiHkjoB8hVlClb4v0N6Y3kF
YFIgdAGv8NdOeLjWThAKkO06PD//Z0e1QfccqpLaT62NCWEgoUsxXHLpKLaVU6hGo/NdsYN6zYjx
MdLOlbYlUekQbV3ML3g2GObRiL2oMCLnul52ShlPlGbRprepxujojoa7pG1XfA4TTyQacJFdvoEp
oDaEy5kQpGF3rK/sottbcxnLr2tgg0U/YDwi++lU5gKE+PsuHlCMVhVNGAl1cxCGeKVTAynk1tit
7nS7k4OCoRGeJCuS/as51TanOCg5QCxZ4eguX4kqXTcLOwL8y4PrKFN3qn8RVyv4p7tbzrc4NI6J
9YiC2vyOkWszKjTY8bgr5LPUeplehOJrS4KjPDTrqR+00JuTWgvMLcCH4dN+pfoTQuZAbJbsYyv+
ljdTFwXLzSlAmzHwuRHLqQPfvtAf/N008853SgJgBvSwpaxmqDeDUMfn5WVjkRcouUACgre0g+f/
LS8aukqe/OE2VdYKmQW+6QGHtJNp51Xc5NMnUs7aQeScK7AdspHwv4vsnmBC8ewEiqSc21abml8d
pUnlM0yCN13XebMgAQTH29AC1BcZY/uFlX8dRIrVnAMHnEMnXyyeYQtG7w5BdVNVamzF1x/M1gwY
dSe1Z2BbCGFXHGBBnviv5ZnlSn/DN7lrjTO4Pc6r9YZIkEes9kI6/6ppnkB7OLC4yeuaWeWVM4TC
mQiNnYzkCUiZYPblWCBDEMm5+x/e8goYEm48THtM1iCOMr4ZaPTAXmrSfw5m069uy59X8TxO+TYH
6ajZfvFtp4eh3I6JVLyxhM+JwkNDjcl51LiisA4LOoaWJTSMFAAtPKEhw9VYsdQ8b211Ud3VEVnQ
ZIiHnK3WswdES0Ut1bd7l8sRbqt1nluLfBe/n0renJSdu6FacflwRkrlTtujFf2fAHcx2a0nPuDm
YiC8P3klSdHNInLkZEK6np2gbILnruD7NS8PuvplOauXrTNOfUFayssMqFg1aIIP4a0lfi6ME3yA
Z5apw627GSgiJjDXEm36csvoInJwYrFMhP48mZrrvNV5OGmGJxEQWmCAb9mCTOpqDMmOS8uGeZXq
b7DiKyzWAx7b/CIZp4tQVbJr8d+DSzVtERpHPLHiueoDmVVYcYiLKJsxFKsZmru4YI7jBNfE+qVL
XkS5LskMPYpwy510Ph1xwIu/bhsVjPbu1SSrNLIOjCfmLK7gs4BEmT1xVN7d9Kdt+zOuItGkUFos
Fap9POreWU2EbI+lkAjArJzbuUKVQpzi4y3XD694qmNXDTYsnXXG+18s70b97P4+IXVPp47qwB1l
tpfOn3rx+OfDWjrgT0f3NClH4tEZzSa59R1+TPtktuJF4muEXpRSJb13zA/wXy9JaDDFgE5EN8lF
gMNPqi1tGvsfT2M6ePWYzcxuYSjd5fx09Xb5QZ2Z4LERZV3aS3EMYzh8V2QB/fRmhc7eif52K/cC
ITZtBskw4isA0kuTbpseNdC2ah5vDr92CRbDTd2qA7BVNcNxFcFA+YU2OSy5+sGejeCuuULYh9sI
J3zmduKxwkGuj2F/nkTayo3gBiwc9kyk+uLRyaHYDqlX2W5Vju4+3EZEza43zVvHepbmSpmCIrAL
BARx4daRo/0GomkCa3D/F2WuF3KqvpxyapmmZ3W1+5RCPSVW8w1JbOJhQm6pUZJu5yXQYmMZSnQ0
0lHxvdQMTfL4rapAg3SFYMUGJxkn9DdLfTfhiAUlLf0K0Fmkwojh6bOTgFBF/tx4UrefObRfmICP
MdSKgv64bb1Jr8gIjg2eSFsyDU70DPvrkF4BaoViadFU65R1Eh+uztxqv5sx1S98s8DKNlbvfATW
FJvK4x2hU0uYWBKKQWPKwAZyIbVl7tlvcv1ZQauYIJOWEX7t2wW9M+XryqNsx12QVwep4MAWKM8b
PoyABtrLoxznUoutXaXcpaYTvZ3YwToLfHmluQgoT/2cziyjkfuHNWnlF+6fQsdUL5Mk8k/HI/ze
sUvqvuqzEVNeFTkoLWYBeF9Cx1zH1Sm3vlHe15iHK6VHobueNMyQbQeweA0uvumexFFYSNvOg7rD
tUYdVRi4HPGothrSjEeMk/e8KQxB60Qi/19yCmhF+Aunz0cuLLOkLweEBgKxD5mNG64dDOCNesZO
qai+0J2vEfzYC0HXEwXZ169XWl9NW+xQZ3GvrOet99o+qLKxWKonRP5zOVFHD8hcltaSw1kPVWlU
HrGrVS9k5uPpix2Fbf+zi5ri3YKMzD+MObn3CirrZ1A8Ntv+tawma/mCzcGsMgv+0ArObOTpLFsB
RfebHeVcib3pceMirgIotPRPYnAK8G0njqsjVn1dWVvixrtyGcsvfKDixe/4IY64TGQ70N5i7ibr
jP2rdWL4zTlY9IrsI+T8PrYxrd9BXjQ6N3Xd8AlqvKQp0xxx2NngJ20ZmOk7i2Z5hdojnVsOIY/U
YZ8zcWRt434S9ml1UIO90KW3WVrHubAoFqhk8lFrDIFYZJJy8FnJa4z8XFEvGBFfUrHbMqijExRG
wJYpjRgj11r4fm4wbCipDYlsrZ5Jb/TkN6ZwVeQY4baw4m7UAt5VoMbKyu12L3ojAEyS7uB6sL74
s6QDFXxYTrC8YNKuWERx3gi7h+dVc7cOwbPXZ8b/rzEki0G1PlYCfnrnZJbUvjn6uzLbdy9fbmaV
154Gpe9wb1tMyhH1QZRIDxApmJLVhIzYWE02vvDJtcV+mdnE2FKkNFoGyUHeTc+uSffL+dMqDqiq
/k8M6k8yX3cnKco48LoYS2kgGr5rlZOoufpcaavHJeYue2htHXPCQ79CEg7NvNw7ashw2qw7oz1M
J1oAVJ8oLNQDOzF0yG75MuqKTIPklW8678QxiH5S0xog3kigMhuJ1XQdcaE7+GG3Y1k1YMw11USF
ojgDHn7RwMpd4E23ZZpTdRzI1Uo631KafG1elTRPWMytwNE4r2tMhwk6fMGeELjM05+ki/HmEb1U
RH9Du2CVilSMRLw6+2wkkPSwKTB2aDVaZfyA4Zqg49oEzP7rIqf1Uchb2Xd/GkdR626Clw1bwX1B
vTP+ASMBSSfMde0tLOeKtEU4fwgM/Jn7fS/brLLQv31tRVs6xl8jM50CjBqSXjbwkA3dd+SLNBdS
REjCpzNzPODOZlphbogko1x3YYEHOFLQGLUQN/j3D60G2VJ3lbeMQc2nKCU5WhPuGk3tnbnw5pWp
lM7cKwPlUhZ/B7VTXiCKQ4ca+dRweyHsB4YddF+zHvAATzBN8o/XOfOg8c3pB7hIpAoBE6FTiMrc
cBtbA1wJ6L4KeGduTLyr9t3zVjTgSzYR21Qdn2jIS69X+2Ru6LYj/m1qPHcmW/iapYgnX1paSANV
FEC3vrWqH7hOFAfDShE988a+GxkZp0m9MaG5kSGPubxw51pv7/1IwENEznEyc+HD5XlwI+rghLPJ
gpCxB0gpE2+YtYZr6cIsHmMQRlFydV0sNvKZzYBPpcUKIb5rC1AbcwDnLL3kd6MfJGb83rOK6pOo
IQs4BJKAnPpz2IwJP7ZfJjpDCA6S0hGntM+Vzh9xsAgLpJT2ZKH55whlc2J077JS0FpBXX+7d883
YToedt39877S0Nmy9FkwYmytMSmAG/aCH4e4wO8cDKRmZWSeOkreKbkVxs47tQJhpA2AAMKIU2/8
B/jKgwpu0OfVArdV5XvGS5hdtK1kkE3kvF5SiZHPaM0fiwyrvoaI2mKylfnYbLtz4GjgTIw0wW2t
77Q+NFbwApnBqWE8768cfRIGCaH9JHweR/cIYFdU1l03hwa9hrNv6w5Ri49QNUaGX2dt/MslSqm3
x+/c8Ko4dw+8mdK0IuEKuf+/hpWunSsVBt/9c3t3ydBKeDCC+GIMucrdGpdUM1cp5YIde/M4truY
P9P+IaUiPwiFscxukIGssOpbYb78Uqe/yf1yyudWRkANCaNj4dKHekYJv8AazZrtbWvw8GQH1lXy
+cphBJ10ZmTRAHJpMq//v0KnKgSLBtBCY1+Lnon/Or+Avq84o8QTr2lkGQJ8AS/moSDreMIxZJuo
lyxmMQdUJWqotVvfgwDTC+pEvBZFHqgvsQ0MEcNA/SZ2q1GyOzZSWH7tR7B/Hu/1LaKqIoIzg4s9
9m9Bma0fT70xM4D3Jtrzw3jK42Hs4Jy2KXFdP6sT3F0vFIfYC9rVf9ySmVeelRUqIuOwTfKVc7Sz
HhVdDE+0fCARscDShoI5rJJChjyppHicABA01gWirk+lDv1i9iz0+pnr4DXLlUbCPzMVgEN5lMjv
3/ZdYCcL1th+V1V65AJeCr/tk+w6TIqgYg2A4be6RAdDkxxCnQicq3Avylws0YPoMJSusixqXmwy
tWbxKz5V2mM/JbUNM5ZPgN/ESyXHcvsWgkP3VNK7eN47hImCYKllUOr4SjYoyosqn8u6DfdPJ0x8
Ea7yJYqUy3C4xB+pqBUSLgbDd+O8BwPtVfV2ieJzrCRNK7+EmcP0gdScUYjSu3eUKn7esz4gEdEX
r388Bg9NQu//pI15z/Ss65E5MWlJTqc7PGI94RDK7gZqeD/GnQOW9w/1DMDvEgojcl+3AQrSTroo
TWSDZhMVDrv4xD210LomIRHpah0EeUK77sM9cnWGaWfj7VDJX2J5Cy++sM0iZpEXNpIWsfv3T3do
P0bpkRfZhXQLN+lEUpRkQ7Mhk8yauCfp+MERPFl+LLrhaffDepwxia5yvBuVD/FX4L0MloXmzppy
+g8E84Vq9KI/2o0TR/rmDeGvRDeuRNPhEVgRd+pKUXxBeLqCkdG/TACuGg/1letKU/pVDVvGEUo+
TftnqnreNeaTt95fLXdrCI/bkOZxryK5JGVNSpjuQIz/L/1JqZr4Irp0CX8D3BoAalW4Z4zQZMkb
r52j8gD0xpaBBI9+3vJ3ojMdYaOV4D56SeqW6vY86mgB4AZrg+MQyfVLtj47721/LmgLz3gkLfOP
kJjJ1RmS0R1zFmX+BdnKPmQFAwItXCuAVaUmL2f8NJ/AUD6alCycHydGpSjtx5j3bAOLaZ4JJBDY
ToB3QYTlqcZTAEn1irVg37TtMAZHJTbYJCt/IJkvQxnSWgkUtvg9CeNlFZk+gJ8o7OmnUCcZYfTI
tJkFMTuKjN/M1R6DjAFok5ITTE5zAYXE8PsAlBVmNc4HbgOg1jgE20OJIPe8PfCJDgqy5PrDvi04
ByicG2v/F+nEpcXzqi8JdmcyIyNsU49ry/8Ev/+BOv9s6I9ClBl9h72ajaPjQuV2qIvYMSnihEWC
B8h2x+vQBI6ANi0x6zH5BL4RLqe2z0iMg2jnibhVkJ78GXBG90cvKRHnNku8uAmTsXYGtSOLmZEY
wt0eg+BMtoIJu2yunr3UNrL8F7IA75gfdn6Em5//qXIS3HeBZxWatYENTkMYsOXDSRACt4w6Xxmw
wCWulBWjNNz57FazNvZ4fkLuNzbUKvkPGUQUzCAEOhN70W5qu5zrBnNazlc2UqAa2/SNRWRSV4HK
jQUgXDkmyJzNFn6cyaxEq3GMCCLJt1bbGQDKUXM8DbJ/wy1bECRzfk+xFYP6G5EaDujU6nEcOxA9
gHkxjHwxdIVd5+AxPQ6cI8L3uqiXokEV8R2sZl+OPv8c7IFevL/0VQMlrS424zQQvNfPJ2KgUXCg
axnREPrTUxqNiPvygZ5/3eCZIHHOKBKEICK8DapzTv584Hcl0Cf3TRpxpxwgOuLc9ObBm+5kwU68
6gleTEkZVG/reQZDlJPS7i0RGXUSH572smpfqUqDMLjGGJTm5sbSRsfuekw2vgxiKYgfgogtwBgj
yz8O30vecdvMMaojGybhI8YL4UajwDFqfoR3LLLgb6O5573FbwuUiRx8KWA2hgTijYW1nl9JNtKk
FbbmM7cDphfMW1x9nl0tMIcOVsVQVvW9iR+MNCqPc8+xPjwwqegpQGZaFFgxSuhnlQiW50zOkjjX
ge97RqqgMTlX3o3wbBL7vLoq2LJR77eOxP+fzCVE6BqUAFJOl1K85JeKNGufAoFbZMdlYdZHG+X2
id0shViFidXBcK5tcYXdJHSVfKhyMEFxl/PFKN/dXgo4111tvpM5+btW9VHUcn2mJ8CJPY6P3sn5
aV9dC9G2rYGlksqbazDzE3HyEtghZ9+TpH/z0aJuh1NwbMbV9kwumyb+iGljWpENtkxHKQtHMTGq
h2tcY+4fjKGPdWkqIzSmpuShfoC03tSYbQJ0INkSZLolv2Ry01CU5WKw6yenzqefnK5Ha/Srvz8v
zAscns/o1ciZcVTHqOw1vbWJbUz/KU2CWw6URE7ip2GS/KX0VBy2GtDF6PM46BUytWFXntPva9ml
TWGQvIBl8GFgUveMo0ubDvAbENU4zCBtb6IYyEfawBB9YzaTDW/15Gb44ApHeDl8xjgyrFvi/Bko
NrTYCdsFqddNh7HDXJUEdFetwkUufCSD0yEz0B0B6iRLOPyDQ8NiHPPY7ar1mHChY6o5bdOmvk7G
9MWe6uPNiQg84VC1rdcfznKfzIizoNrWpV9/y8x5TyhHKVh/HY1l8qqNeYHPuiRuaC/h1mnnvgeH
npbiSfVwOiWEs1aJzJ5iWCeXEvFqdWC6oHNqCtDUq1xdxqY+l+ABhbx8TFDYups77CfKZfvv/8hY
B+XzsIj+RKYOkQPE4+Zz4OAGUBtnhCuwyMs3dJsWokKBGQ+qQaPGmyRACL/5jH1BR7cm4bYTghFR
nbLllEWYNwJQ3bPOiDUdl28m0YaPfeYr/llPVmDXb56iamdhPyNEANISbqyJkw313t1OR41KxYvF
o1zJYbarkOF9LqFyzHIaTu9DLlbHKL5xHjYNFhMiU2UoU85ZwS6IUb1F5/ilxUYO4WSBUw8ReZFs
fCkqo+n4LtoBOJkjz0PlIZuOFdUPV1yomYaeIGOiYo5t1WJ176OC3WVj5WqXCyn4+I5sLknW/xyj
CoqYctNf5zhTw+RkW8jg+S68nFfRZkaUpjuBt0ukT0FR4DMjQukeKoafmsfzNHDuZx+Nlxgj5dak
XReDacKkxdCvkoJzDAyBFhKLETBIIsoL/yQr7dmufqa+ebcce35sg+27gl1lJXTfdjBZQQFjE2oh
lUjVicdC2lpPlKgLwcMtFrUmTwrKJd4ETvPgYoUNRJANjX+972N9lt8SvjzKUW4ddFaLPw/riRiJ
uhBurht+K/+uSySU6SH53roAZ88V3m27G7NPVNXvVbfiIulF9kfMI62wzvq/tXpyMz1IN29HxacH
tiYLv/p5TuN8tNBCBgC5vslaETtCuD+di8/xRr+qRtITgPUUjdAOOzkUKAoI3KX6QE9Eup5Pf0Ww
m/XAKvW2mFvPMccBYYtVl3HPM9gBLgAFvfzwAMTAO54codnJlENPaAHrvNg5NwzQd3fupStuVskh
mIeHhMl4plKuELW71xhUqh+kbBfgjZ+dA4Q/y+LXjNgJHiXN5g7dVzk98ERSn0nSZom4iybUHYxP
FkWK+Z6mV0+rXNcr/LQH9BhWZWNwrfBXxehOL34CQ+j90TYfRa1sDbgjwQ2WBXinnNmJgJpyOtXD
PK8lRDyOApIbUgBTE1jgPIzM2BrT3GuyQJBM7xlhb5fGRA4omk01X7FybvT3OiLGPAHSaZvvlf7E
SbiQ75iFwlfdS7h1xfU8if6oYA7jm7QCrxrjRvxFBEcxLJE3PY88aSNcO+qCQaqNztVCEPtKU521
dreI18NApeI3HS5Be8Qw7q11+m9/vJVAOM5O+5xR33Ob/ZBT+GkP1OrEq19kdbh+nEfiBCSfwnp5
YBjmrKNiR9b2AkMgs5W+bdlU0+NXvYD1BLuAPMAZQtvDnxn0FOUXvK/BPsLZHUSNcFPbZGrPXoTL
B5zLNmhmYUjYmV4XTrQIcqSbiHRS7t3I6z3p5Wrl7SzcL5bjqycGiaTEp2YCaQnciVOOVWrE1IXs
oIdiKCaYBg6Cu7yxNtHd4LJrvHuvzaR2RZmjONyD3MW8U39e9ZssYbXmF+q3QnqbQi8v+FRPjZ4k
HZiO0yy3c2KcpSXZixX3A2BzVPOkOanIynQdqhTJDoLRqHC7ez4Mwxedfiy8VVV+7FF5Mi86LT5v
l751f6su/KdK0tVSwdE5Gp2byQOzbsKWt/k2XWDgff0YBXIHMVh+A/jqMX+2f+o/KVgRKdWBvu19
vg2JAqE/FBzlXn0xKug5E+tqnpsGJDzaV3fqLBCFYDRId97MrIi/Mx6XP6QbO5JsUvcwOx1FvDrH
aiFPuyRLqauuZ7xC3M8QNK94Z5GFszOrStT48d9URv7CWB27J4irzH0H7fudKM6w+aq95r++05H7
4j90vxP/+nV/BG9FvJ5+i9KCPGjPJ+Ac4doO1+D06ZUoHB2Dy8fj1i0PubZBshrT9HhAACP5G0T+
/JirflVKH7C2l3LQPCKx7Jd30BBjzyN2ZemtLdcckzqy6Y/5TA6ESnqe/Rbv8QTKOyn/adzI6S8G
n/z0xjaPPVgXxBx+zWjo/mx8YAVuElgT+BsnRCA4n6a/TeE0qcoumDhKOHxUCIfOKXcC5LzZ83Zj
Epp3X6TrGrw+JTKyrzaNMK4trTBvj59KzBgtx9g572ZEfoo5zEz9i1onSTxiIfotbGa/K5KsHaFm
c1/oXwbbdG2midBdUpj+tkKUb10TCy6yHL/vAUC0Wo9nUgnRyV9lvJ28qct1ivL7w9lG3cMAtvzY
zjYS3LMmdBZSJ+8v6j0lIfmItrmN5P93sx6HdFhvl9deocuL+KC/OA3mrlFQP+4fogLA2FMqqF9l
s6YPiT5Ef4+Gdr+znnqDWmP9NWFowLHMhek97IoXAHtwSopRPPfF63T21fXOV+WxvQ8g+NUPZyvd
V91YFfop56h7mZCsz5SynD7lAVQoJCWr1xeeLe7Tnr2GTmnA7zCOjzR9AF6Zz3uji2mjBjPr/9vF
av4D75bUTcJ6HNkg4MS/qKv7k/uB/DUueiIrzu3hP70JbHEQAV6tMnuQW0yZSUHakxzg2wMso+Yq
AinTYM9QExW0IiQ9cD9oYjNaH6ong5PxNNFQuWzFybXGdQzP6MfrdHfFg9MwI1pYQTNLECIdlia5
01uEQDhLdc6FKXqdtdRIP+XC/+JLJRA6100eWagb71tjSzpe5WLsCxpCYHUw0ZX6s3SObTRQG6s+
/Y89qwiIRAzxgusPvAWa5phCfb4hTky20HP2CQBZd05ecHBfs7K3dESAH2iopc5rdUUfFunVaSH0
3McfMtY+wzQVVZ1PM1hA2JI7G+YnKSEIrZLMqUUAF3ThDcPfJRJXSczgPqYYkPadTNlmjZ7iYHIA
Cgq5SEX/rSQ+qJyQWRbgbTmRS+Pwja9wMAfAwtFYXDtnP0AWMvVX3+Lk1tlfnyLJWOBznLSACHJA
w5AE0aysv78+1OyN8IGDLQCrkWATOy1jbQZ6lQfG4VGfDDu+a8ow4LVIdZARJtIFQpZ/bsA0GphS
kCbWm/sEOX1X1YmqRO3rFkzjECSmeMDRYwp/gUTjZp4ihqr7erguAxyJl2sBEDEVcVq2J8HMbLfH
93SQC9RLlro6kfNZMeY0CmHofyBnyboNg4ThBX1vmgSAQIknWnKTEX5yHGnhk50IB4H//jhKzP8T
GI2mnMGcF0WogdvBmP49jBe+4/Q4jjZUPw9Z4TB5qOnU7xeRZaB8r6/gzp6lMN9Ra3a8z/eBmepg
Tv6scumSmGTLC376cc/eFsMGy8CjccWskN0gg/WFIOx/GwpOMxUDUn31D6qa/xXzqt3m9dwENbEV
EwJpr3KJjt0vDN8sWi4EpyO2qYu9a3uCnzUzAQ2/cSPjpKRnwz9SCaIaqewaKMJETQXznZ6f/qiC
jOaL/qtmFYjFEVU9nf+0qjcRBjKPsWgh9CIXSUTGX9fKcvIBfydvXtGqmdkm0rbSNbtcgvRK8u/3
06Z9jWSYJbH/0pXgCnjMmKKg/XmOVX8PkcY3vrVMPmsRAxBy32jCvM7NKeDRd3l2lUjW1HL4LZMj
LnbtT2XOYhrYHsGJv6u62Ngt9E3aY15acPwU94t4awmV/ZzEFxVf/owj/ILebt/fu47sRr/ZpwQE
41ldGSW+gVtGTEioI9tIExtMENmuiryoyDlxW3zF+NMgDrheSf07gtYH7Ccj3Yu8ukC+MrxR5yPb
ckVi9ywF0n3l/ygJclGHTCnxDSW0yptUo0BkarQ8r5jgo2hfkMgQfi9kOBnA21P1U23s+4VCUSOs
BMDsJ0IhymRoSCzpwU1Ybnqwnq81nLR2loezNj5e4JcXz2WpBRGFw6+QOgj7pil9zoKqth8jhq8b
fN4D9d7ZXUa0eA9wA7Zf7xWRTef9YENHRCUne/UjOYY5nBDLxfh+3SlK1EWAoGpsLC1NzjDTtOws
IbhUA8o7okbVGmxm64I74+T/Bt5HZFAf/LOaiwlhgnDwoON/P4j1VA5ovz9go1X3PcZcQ6BCuu0R
vmCLvQ6lHazDODWqq+s0TRoVMf97W1KToWzCvx0JcguKjypuSEag/VT3aEkRn89++TsmVLlPpzo3
FJM6brXgMsMuKXUG5UQju0r6fHbO/ag5lQZaTIAohDo3lWtpECiiefuwjyS9Kakd3nlsnNCW/MMQ
qlPjq4RWBlYwsILuo1svV0LLfDtivUuegHTLhBXwCp4RnzKBytM2a2EXhlLLf7etgjoD1V6Qkvpc
h02wITEU+qzhfayakzdVWMxWBdgymivt85qCCgWkucFYiyYnyZnn6L3wiJoWykpJHmTTpFowyy1T
kdXJWNcBeuK6zJhKEmVZeYf0+TkXXixyovBFIvqi2TfkuBGOzz6sv3aCQsjSHNOY0FbrKgsDmsYs
Z5rTip6cRH0TnYiZZTvTEoXOlJ8PGOpw2/vz7MQj9l0gGCutIEWr/EnEPdRh9hxXD+4AiJ7N2tO8
16Rdhsqc7HHtCGP3hJbxAXX0DdnLXPrbXoiFq4GfrJ67KDce65zBFOzPYsr5FK2pNhs7/NGAd3Mg
eyXJlbwS5ryXzDKOEOT53VnEJPuTTRheZjIxGavSb49G965wjvBphBVeSoiSiO8CAVV1UW0iYhLI
aWJAaVPbc95+Q/gKtJIwwWQAasDB9xYb2pzNegHCqMHXFOaXtyjEmc2xNlxhdNlZ/0wMjnXAfElK
zf08DeS/n91BbSTbIBI2mFoqx6GplaIgeSSS1ItE2A/Pdt9mE0lqPF9YjE5R3ku7I7egq9ehLaej
cc3fYjyH1S4bS56RBwsfFFQj2D4PMXr4TtGF/IaEUsO7omEZDqL3HDwwTnO4WX/O13WL3QGgz7ol
QA0JKxllnaCbRA9x18krjxI0nH2fBSrOQWRBzgH7oGToDZFdzG+PCQvllJzxTfLshJ3UC5k6OsTc
txNccApgFH6ztYI1fMAYNPAxueFRVEDJ0jYqQAjsTPQ9ZWldZdmYGyFzq+1XBj1TYvwu+6CjMsUt
ZJuIsu4GYY5nwVeB0RhdL0dYz1ceCc/iSOG1SIsU2RpQ6nAtCwGl4PvJKUxAmFT/roTxApR0GAi/
5C9bGSAa/H1NhhsL7p40MmtesUSCkEULmwuRuKAmugwJboCJ5In4GmQqXe9sSbYIfMB2oDNHSgWU
57V6ADa4okuBUA9NBURCblv79oM7e/Np9lDbAW7Fu8PFWcCORE923Lhn6k2veuEpPE4Scg+yKXfb
XLNuHJxL9aBBulSuUvVD/2rffMmr3DJDpBkTaDUBp+g9IEwxsNGfKs91W8WrNbV6Opur2n5it4tK
IZIXVm62K8M6+NHUyWlYu+pSg9xsd+MEqOtKisGt+GDXk5DaQyJGhU0rN+LgzhF5/vdNtxM2kdnS
K154kAmpBw3C469YgFxl/M1sv9OKHT2eCytLXRSvJdOhRMvIaS2/aQql6nzXusV3+FZHVNakRXGw
WYfHY4JEOEye8bnhYpMTQPNP0HPSeCNFgxS+Mtj/XSpqH4WUUHoIdIICI6G8s4LMznppRfJTEeJH
qHF7MjcSQJtFJ4V+7lmSWxPnqFQolsQR0tB2aIlJsgtrqbo6JD/zqRyZx6nUty7g9uU5hpVIE2uB
cb/BC7Ly+G8259Z0N7+6pVqbiN1ZpUcW+2o/iSM5EX/7f8PWmyuDNEpzE2rwtmR6ch596VS3kxlA
1OFjysajQ0VJES6LmhpghGhgca/Pa0CsmTtcEfzWOPJ0IdA0iWFK8fGorEXHNcVBJntqbkVF3/Fy
ffBN86ge49X6E91p7QBlhkZ8kNJrCDSCFJsMZEXPfbikvt2FQeSdra9bwbg8h0IeprJrJju11hkS
uutVMyYLw1MJz15IKFoAmNKGeWDH6I+MnLm6QwnFLz5upo+YXDEG62BQvH38iRL5ZngJTPmOMkmH
3AqpTJ7+PmTtdcba+P4f8UbXUCjsWKn4K4zEXMQ13o3nQkI/OA1SFeccLEYWKwMELqD8ncb24h7v
mN0ceumBysiIYayRMxNYcjAtTsUX3cyjBJLWxBSsfoRj/GIF8U4QZlM6Bt0WYPl7W2AvD1YRNtdP
34eLewihBrNWWYiAhfKeLIUUTK3XtKykoR+sFX6cvrMZlDA6tElLgbw0bpNtJQ5hrXekdNHk7d98
iJuFCRbJO2hJpJKEbSgCcVsz+6x8G+kD0cnUEP9rQGpBaD/JY2k6g0QdUnRMunv46B0my3KdGbQz
J+U1qBKndLvsPUZAsEHn+/6LnEChTUOzch+ferdaByOCcX0rhwU49/yCmgnTH/ftCJepeHabQXJt
KCJskcabnwQYJCOLqqtwUlXH/pWX59OGLzMzj/Xq1amysXQ0kDBGEGeG2MV6oNN9eVGqDtKRehKz
9OZs6mQn9l4RTPv+p4QRMI9bXVZjqlQYeUYR37O3uKQ6KNU+CpXGLvFifo0huHlYfEJorNmLBDbs
31RohqEpThKOxQxYKNJOaOKY9aruRKay0afSBADPfbq8g77v0OEXZejNyxlZrT9jeT/cijZlVnMT
HFtY/R3Ci1B2zqUkdyh0/rk+j3ri7IbbyObWimeLoCw0Iuo5gi8hRCaFLGYPgLWCgopHUu1E2Saj
oHsvrDinJB4+lZBFo7S06CUE7eREiXX8Amh6uZP4VbXjkOP2V7ViIT8SHElcm7FmQASXtKgDuDrD
Ph4c9KWLcENS4u/9v1V7Iydfr/m8/i+7ssFK4NCHfws1BZD+n9PMHipLW8KWTlIuzj4rocJZOGn9
i0ubIwBW2Df35GStPo9Bl2Xuh5EtoEHOEUbIO99RpNtZ21V7fuu99NOK0EAGm3kpJhPwxm4qN0FA
HQ9o3Di3D05exKcvXjRilkbfEN0n8QhRL1ZW1Ugp7ue9cu0DKhq7TixjFKz6plkqvhsfmbTHFZNy
yiihi7BBCZUgRAzOKk4WVomzNMzV7kYGKhsQu/doiud2fWEkm1EQNl5HkVDA6fLdFYV2U72S7Gbx
wjY7vfBDqfhXoGQIPxvL+qQoj/NjoO6Awx8yXFiQ8Z4uvT+xwUqfY4F1CwaZxku/p03TpaIAJ3Bk
0PDbVboga9xqsVF4BP8IP+ev8WUaZ1RAPOwkHwfFF4mMAfWLx/rQciV3z0zoSuKDJKWQfxSwUl5f
gFcpFZHGGUavGpCa6kbE8abVv/0Kv7NKoCVr3ROZNrJx6tAhPFniKFYt65qGP3bD/UQ3Qt03aT5S
W/Bxp5lBXttkBl6KpaAC41tE4WqbrxG6y/CclwGNIq9RplNb2NR7ZnC0ghkB5J9J/iOTVGuVt9Hw
heoejq146JNW702UzUj6r9YFjjn8sRPe2jlMd+Mn9Dy+2rm0Bo+R5JLHDpwM5DwB3fJyHKu9X2Zf
D1LBY9A/Ys6ORq2pOJJoRAJ7kk/kOYI8mnce02hwdtmhNVWJQwmOOVRa2G3vi0ABsgRYbXf+JUxU
AsCz70pxuJWGf8MxdMksuH5q1cyn6Y9cBPGIF37XapouROwWuk9mf7c1ZjaU8BmJguTaYzcuaSNC
oNchouZQLQvQ39y6eetyYMgcBNJ5dswyV+PNmoyW2yZ3tEEv5MduBx+jWmqZNq0iiEueTjS8CTLv
+9MVAxqYtTSi6+QMYIplzeXezfjREtfO7EYykUSVDdyzmY9Pn/ukutwkGEidTOPVMPXFgsUMoJZs
mG86mJYPiHUDRcJD+meZlRyNcRt7zDO+daHHmtjDl5k3XxSQ0WaPijFjKLHYlES+rmMHhpl5u3eA
aWBH8971EcP8yh3FxY/sa9/erYrVv+0TyVzFLj6IBkODCzZBLZvyTq9zzMT6YSsHhTSkGYirV1CB
dGoqoKoZATpU5F/ebnPp5dKd8S2wigzM6uLfrfAPgMdHV5uugrAJnEQxt1CUpH6lrtVAPiSillDE
jwAgkowzARaTQnqfJGmMiDxHENg0Bj1f6CycYrktFTNALGbEEFVh9Pp/mS6obAlftcw4iKJX6QIz
9k3TFDPy2nnitAEgx62EwChcYhHQHBLwMrjQZF1I4DyGXqI6NusvbevHXCN8w9Ue7jMQEXcopyAC
+PSyDxZ5V/0MuBYVcNrzR88AIJAzQFXYll/UogP0F2xsT31aXzUm7G5hvUa929H7tXCJp0Z1ym5t
4Mxnu8Ecg30BQzVCkB7IZbVsGUVx0KUtLKITq/TMWMUJ2DcOH5zUtbxvGg5CmBLcj7VwA6xVD9JO
Y/n7ONBkzFfQYU+pL3QMH1+tGMoo4agIfak0gb+D/lpZwPp7/ZtkODZGEmZK+jD3itdjt66Y82RJ
GiD6NIKhYiBjAKgN4NVBwkZ1BqjIevcaUV9A4oc6M3ILCtzdSKdWWojyr7t/0xuwMQzb3xPMRx8p
ZJGsNsHvU/ACrhHXno8h5xAa5lpbRkqNoSBipgy4cWwROwEkX59KcSLXsqN8lbclxX3GSUH4l5ae
u71ZNSf0DMns+gluqGJtydo4AleWcaHPbtOsHHRXp9tJuvpB1rY9EQeWFfECtNrknAnu9eAOn2Sd
l+x+Wx9vkAm2+xOQnQB/CLLHT5XFr6u4WG1g5gVwyQNJGPpWuc+53ztIYBvR7rETbZB2ViPoLkgX
hh0C+Y/Mqffar+HnFW6WJJs4AWuhaOZy0DsjLO5W0SfcMjV9HwUcQgiQT3jqQwFvz7qI4hCOvvDW
K9S+8J+lnZBAvmw3PvZtYzZNNzz8eE7XJtg/MRmX9BaYK9pJpO1w7NzsLxs6V6+FvrVPehUPiHxA
fzOcRjYMqaZJ/HAdEfL8vBqvXyRGdNE5kx+PEddGE678Xodb7Bsh+KfgFYhL7uGyPJTXEvC5AgVt
eTFQO52z9Lc2byetwmyCSQXKN9XqvlnFFi8oc8QfzWc/EJ5/A2C4/X5zZnbcScH/hL5MXuZusrHp
F0torXPMdbUMj96z1zdlmgTWWwhjcj/YBKOCel8OacEFHGGGHjmClihBhET0XaRllPDn+dv4tt0p
W07CmOMxhfC4N0YOXdDg806J2FM7PBt5P1OiNuwOTMwMRv5IJHnH/vGtIvqdwvx6JsKvEJLXOUnm
F1NwQ9w6sTo4irU+38GSEJM0tW8qFNYz0yPZaWciuvcaPkt91GW4Jmam2NqgZxkzJ6rrbmDpTubo
Udv+ZOucTWxpRS0YkNreKZMbd3VaylR9d9ZOCR0Azu3aTbNxpdop3LvQynRRwpnnGtE6AK12vk3Z
FNrWpz/5Q3u8IwmmcqFKkemkXjfoOWRzBljUUANoBK6uefjWQloov0AC5HZUcbEalSwpCC/c29hX
1OLAz/q0YTTUaqJ+kTmPCkG+Rg/3bS79TXiHgduv7gO8glI41Rqkb4tBDgHDv3Nk9p5eBTc1ATsd
eP4pypISZf4SWULoQAeC00BzLqEhl9Uu8HvfvzXLfF10mU7ACY0a5FG1HZNIKggd3VPbagVNheIC
I8ZJkwH7/8wfKtP6A4wbm4vXcTwN/2itmcweU3gnuPAUktxIxhD/SsBVS2KeseLDrr4AteVJOUr5
KZVpEcwuEMRvwBPD03z6N1G067ymja4sDUZGkbMHEQsi0QZP06FUd7+8rTxyrBd2ge6Loh2BjgJ2
e65pXa309NcCL7hwc8rSW46eIQ8IMySaAicOg4Nw2f+XqHCfViEbccsRV6wElEZOmbRdtNg3bza+
/Eg3LmPVYGdJKDmh5q6CYqO9xIVHawJioti9mTbSgk985G1Xpdkz+yU5xK516Az0nAUK4+YFqwmM
qrKGqTNNPgTEmOjCqzVKuDdKsqwSE9mJfECY83f1bRN+7I68YDZUdry6RF1KSHteZbStufp5fy3x
GK2vShTKR2XuHRvJu7oIGBMZTiu+mMBa26cv7eVN/kWi1Hu2d9OGArN+AWTFlIqwLNxwwoNTmH8O
fN+9XGA13fT2iwoGvnPZQa4SgNYnq8TpSd+ZVuRpxKjFAQEoURCmoPY3pbMTUf3+8NS+8UEUhu45
HsesAohSiuHKggd8IWpWfuijWPc3EkpZNlgJv/WhcpOzsH2+XLZufiE1qt2sCALTz8x0wsbsoNQq
I/gq28gAV9VghmFfAC+DnSoKT2YITK78z65wFYy7knmPcwpgRkVXLFDoI7zeZuu35x1lIQEv84o+
i03zLPSCaikmQn/ix+75Z8QFzkreZp06phy/ZuASQA5GlaKl/njfqlemA8IJRxpAVPRxxgsYMYax
m5YpuwotAOZ0qVeaP9NKCt7x28o3yvswpyrfCLnO03kjRYhLGeA8Cj07hT/X/WMDRcahF+Vt96gG
fX7LHeKkgXBtoGzWb86hgMbpcQ3UuzPrfdHRPTt9tgx6DOCKcWUJKRjihJ+32tu+/YeiFG6EtMu2
j6mUx8k9GpWASHwSd5fuIKG2pKGOLJHu0g1gSib+Iv5cEvSbqVLfMiOISSyJvmvqK63ord5YR1B4
fk3vs1rsNxf2JUbeRSPUFpqDf+sIl6DCqOAV9bHWtgjVxudE7eN878wgmiI/miYPz+ehcq8dC6hp
0y/FpAOlOuPiyrs9RBzGxdhz8SCXGkL46XqkGbYWcTaheKAIReIeCa/7e20nRzODEBs7GPR/ru1w
Yvkn0wGUkXu3iE3ANBMViXeg7QJxdZ7kYuhco7BftKG6aKGmdXHJE9/IUM2t7Vhv6fW2+LVE7x/R
gog1LBgn1Ghc8oqgYen2ZUHTnGIPexrkb2IVWc2O5UWPtqeR2HyYeBtrpGRGzov7/e/r2AoaZ+Ei
G5ZwQcs+OqOEKv/hlHNIMr6xXczcnguJy0USec2HRNqQ3XDq0Azv0e1I4Xze8oHS8I0wfAea/9y7
6AkOZ6xZpAs+oyH5sMOhjjWszhfGPJQY5akdPat1gpPCDF5nh5Sb1Eec9Wd1K/6TJX2P9aG+zZpd
hsmDteMmRcrB4hfxahHgyWL0VvYwEJ2BjoL+c2xGDVkn40934IkpfTLN30H5lcKvniv7GL9+zcd6
zNQfq3x5oS5ZsE/v60LBb9qRBbkSX2wWgfrS2bP9xDQp+2caJX8ScdxLJcs2YbBQG0CO8sLm7fFv
qLo2/5Q1VqlZUe/iF6HBPjBDmDAydEvap8m/W4oPW8ioyO23u+h2y1INkGdomya7ox7r2MzWChYX
2PBdqeQRQwUwgzLijUZRfZbUHIrtRCbs6r1+ziMNdfAsaz0ITplZ4WL8Tw3xP75wlozvr+KTaE2K
XDlSPMmfvJFH2aJuMZ+xHq/bOBxTYbP5+D1RyXNPxrz05nPQO3p9HwmrxzN9aT35Y1jl5Ppz3M+g
r2X72jx+9yoyXLZOdvZa5bXKdww3DK3Lt6KlXoQ0BW59RQkmuyEp7oIQ91JCkkLS3yCV6zRQJHTY
UMaCezDQko5/C4vUoZj+KVqXmHrWoWkQraBGKkKejW26FgUzSclliE34ubnBJkBMN7HRElglKRMf
5uq4OFSfMRbfQsFhHwUFA5X+6OpyjIqSaZrvmJPf/OGM2LLkKvUxJgvGH923qu5cp10TRimBtZpq
wRTDLFBSydS9QtiPJyYewrbYGtBM8fD9WjCclokWv2w9wcvuAddnTxDDxCzYKPVMxBuCOcgzTfmb
XZDmENaN4zDTMH5y49OUa9rbcNG1OtGVpJNOa3FaKhl5v31LEXs8XMniZKRWI/MuMJnED7IOLCBZ
3qPOZaw8Om4FSJ/ZQ1OmBhEMlW8bO66afLxkQIoUuPRIaYVsSzs5IwgEpGqaBeqmLimMXulsRE9C
49noWayKOGn0aUOF8ilB/KpY7zCLeQJ/8dRZcwuALlGOexhlc1gpeJLmHKaiveBh5ln524Y5986J
Fs9K8IB8Q2/Gtcn021e521Rc4qO/dFCFUYamfdbckqux/aRjGXLexkI36lgx9KaHYr33n5kEcW7z
Ppe3qBpkf44hcUrQ98skidwmYsl+kqX9Gi9YKrHqL0txRCNCqs5PpEd2URMBVdradH//aAdjM2Gu
vzyFz2uWInAJzl2+Q3FGcFvJTUR3SC+caw5t9eHEOl77wHN/V6sp5MM8V0Cy8MaRn9vCQup7mz1g
wzdWyxAZUFZE1L/NQozeEHhYSvWZjQPrOj0DtlgFxRI52zAtly4yEMmLFGAJESG3ekwaB/xFa5kZ
4TPTWke4nvNZN1zJbsuIs1le7OzvBnGN9UYSWBr4HGWQfJ+aHHDvTk6kpclp4wUhk80bngxMSZPN
2LYegCBu1RDBVo7zWPd8AwGSGVDO3pZHHRjkfN0C6xQOu6PTUcl4XXUGSk/eKTO7CNmNLbIoK+n0
cNDU9iwOoWNzeSm1CSXGHOyt8drVl9TYundf/Bl4YTcad9TasnH8xZbHZykBVmXHgCrNyYJmnYow
zcT3wxKScTgg3vVx0XwgSvQ7I28UJ80KMutYJqHNx7h8CY+OVoeKJLJEEtx6Is10QAPeF6jap1Mq
+Y9lA0nq2AS6NSQdOOPnO1cD0em8q4OCWk7z6adCcd+7fPtbqm8Tv+pOXRsahhoJob8V5LzSI68g
Q3eyado79yYNnnWeiT7qdHuWDr7HE2FpJZFh9kjjw3RlPOzA5148EUqZcfTQqSG/wyUgodmh3sRH
rJckGzlKc6+9/97P2lt6Z2gTjblIIp+HQqsXv6TIJ0W2/9YU1ENG6KMhsD065y9RixcddYl7uvsH
VlzZQgRZxLRo8h/qy5Tt++uPCmyxRNr9IK3VOhS3zeotEGfg15JgJwdGlChkuecfZUH6urlKQB7r
g5sLuHCmZRrmHiWfl63JYuLskA3TNOW4uCcJBgtX2/FEc67CHrJWS8j4QZkcWal2jQyzK3oDhhm3
D/IdYuvvltpQV9IokP6DKD6Pd9jpAOQNJrik7pvMvvJVCphq56niVP4FT4kLKbvoW2qgvUrdlz3t
OFsyi7zScFVTO1mgFtM3MzgPiAIkNBZeapcpNe2OPYQGddURiXZSYKS/b4m8vFmnRHF7Fv9msONF
WPaEkeZhMH7z3ZtyKEfqUqM/ippAnMzxyG+NOhSqjR41ZbTn4RnbQAQlr21sqQPyx3bnBt9Je5Ol
fe15Ttbg4FgwrTba6Xh5cwvi90UR0QS6/GevwSiah33wPV55aTgmRaPzJ+bl6TrtcITkrzNMqWI7
+NJdflcWECoQE/yeUGPHhtr+CxdN2eU6mHL2BfMaRO1OgUePFSzf12maOJDfOVBLG7xNQqrk9nob
wMBSCQgLZ5JAQDGNL4auEHq59M871hX1ziou48FoR3N11ZqFAypvxRq3usvotpCk3z58Crlbzafx
SBRnE/j09ULz/Hc3mKA7bqW9hp4xu8M1fQUaxw6MhmIKEkyxn5f0ilLJzMtTmv8yLbkhda+kHyZf
uCzp+/sTjXY4LFoZKvTpFFbk4c5yKWakpSFQonzHkf4lmKB7uHqHCq/IGrATChy8KNg0/8As91hQ
3jijK3G7MtwKTR53UnIA0zFVoH9/RGdXMy+5PLj/G4aRDlMVvxNOGQEEuS2nxkE1/oTusSEg+w5/
L3V3NZRm0LQDQ16wLdvSBu6GtvnMHskwEKTWhtbInfUliA99otnlW15GfyhpgbyTnhFCyKlOQl4K
krUsf4TlqAupujq/PYyrEfO8JpUZejyfD6IKFbzjL/kM5QaLSX25YLRCMO/rS1y7cFDmmEBpmIxx
XQ1cPhd2GR+UDkewNtKhziomZmzEnIqa9dC7rLvJXqvMRr5y5ATRtNj0piITIQqDYjbLLZO7h4mK
Bxwt4q6op8NlPJE1e15nPpNYakNrDVAP34FnjDICdkHMG1JedAOGtfYoxuYSJIZ6uhsGkjwEcMnN
HvrKcRFjwbhiFZdBXaBOEohs68iibpZvExlOpsuaQ/bpC8NUJZpqeNG5rIMtk1Fb9DMnZN6xpLiG
dbtt7blrJT4+9T4hVBgCSunQBpwe7p0j3McxlGy2ySg5Dvlc8K1DWNCZ+6Dw/vsWDKmsrWSaKG7z
4ScnQYA+lT+Y1aJpylS3wdyctb7Q6aADNR7JPia8iYW//xOvXl/LIxS6WOOh8wV2a39X3X3UIGXs
IaoMl4r008oV+MYa15QpVP2sSj31qhN49LRJV9OZl/VhARwussM0Rl7aevVSF6AWphR6rCPy5JXK
EriG2pCAofpKh/RTsfUCD8a/AqE4fyUcpV80cH8I2YCw/ILwLmTeMiZ9mCaVP/6tvAwg6azmgyFH
tGehgtawpPjnvcGd+99s23oc7fXSOOQEnxiqDXbZ7bzmCahyZUWU3cwkYZYPZTlGOwLeOSbm80n1
xBnrzhzF0DZ12nYuov52/xthJwHxgsghMrb+b0oTvrfzzqo9SWogyFx8mQEEQpVN8mDO+dvMzm45
Ma7OaCc6fjQGCc18tm184mifZHTb4OExkYli7/Kn+DHEaoI9rZWLZg/R7wsOPgXY/fHss7/o8z/e
TFpcR1HGkiTBe9bGf7JSxcif6bs1l+AQK0jk8hNdHKQmzxVTQph1yFY88ToOnKX42XrCib+4nG7s
6r2mVjPPk1QZWCSa1eqqDjIlu48OeptMdmm2d2GDrBJ+s9+TZwiusfCHBM7HKEGphGa63sqgGHdN
nHkIPbnskqZHGeEvjk3cTybVH+PM9XOnb+NfNgJSjX0hfsPrjtbqwrn2Zy7KTbIG6QD96NyPNVbR
5Qg+CDmXvMnZgMQxeXcaYGblNq7RuwEMX5laFKTmSy7iS+GKrvLlaNdwp0Kk+nn/6yjn+w9L1qfy
VxjuLI+2OLbF3NM7i4bX2uJ23d8FbITUg6qVADSLRCYZWROOF27qZjx7u884QEHccsnxG12wFyUX
Sf2NxsjmPC3RCHoj6JDtKCad4dSWN638Pu8ZL9Assyx2hmZ2zWYzsrB5TBR+GwrR1o6H2xZ7KaJc
WJeOHM9Z9lJp5+m2++T3MlzW4xo5XJ0UJFcyDgBHVzNkxllbL8W8YPgIRGm2YcWVW1yNLZsX4mOa
566deL39CI5N+TOBVkFv8j5h6NIw6D2F81UyX/mrsvlEKnxYq0J3rEr/fiqoFmJRtqK3z3RyJ7Un
xOUfQrEphr/nEXbYQD7i1+BPqvGrnCX5VYgilBjCOEQnG3uO9v19xL9GJg9k4NCVM6IYpEk4Kyrv
4uvJ3goJoULlNtof2FNsI1j/jv7u52WC50BN4wV5GCemQKCwCHB8HUarw+S76NCZVAdWIlYaqSoH
9w+1sdhy061kLIglhLcS+zeWHSfz1K7IZhBAH0tmiMG3EaCgfWOKHxHSs6em5tRuq1CqTjHpBgvl
o0o1ds0YRJQKAUbyVnz0rxXsM8vX6qQGKv3jWdPBmZT3YNPEKjjrXdRSNOTVxETHy+8X2Vh8CfE1
jq4dhX9oqtwxBX1lydt8FTbiKqROn1UWTPuR4fuh0g7WuD3CQlcHyQssXYUqQ53F582Zj1w2NLL/
qBh5hozWuKVx82x5ClmX1zUjpG3HxMd74fPuAEZgl9POhdNXq5JKkxeIUG61jBJSVdHugXV1v4rR
xoYonU45nrrjY5YTwO3ql7piX98hXL+Y8gOarlUIdeH0DIPwwWLIKyOQL5cfGZcGhwlV02DZuyCu
sldj5DvQ3DMIxXlzB3qs3kZ5zyMNsQiZyZw8DvQ+TEfP2z7mDgJ1KaHDTr6CgB86z6hQLOfhERQ2
sThGLIwda1cQRWFSqqg/OPaMotxQ+mVteNY8oGbp6L45SmmcOXjQIzXi6SINDEmeZFDyNXbYV3AD
Rz1ju+ekJPBVf6DlJ5FwlqKpJAM47lYheIAQf4b3pItXnHgvW9x3NQmQQi8nbR1o0/y12w8PlH50
AjeX3b3kqaArWUL1eA6lFuEylePwbao1QXeuCY50jPuuBhyrqwuwkCcFsKOBm0H7720zrY61C5ts
2rA5qllaA1EQiptKkzdJ16BwA6e0rcAkwAvU5J/2ViZmLmCkemESYD2ws1CZnDFr3Lq7JIw+Qwig
ncWiieXBe9nuiBk7S2ekrxGe8e2pj9qFLHGz7l01MzLQdGpQ0ynDXJaq8zjvq4aJw5R+lbh0gAnx
Va5Xoap00Ma/mFV5JBjnl7WtYdWEVocaCvgORR4wqrZcfTTGnjiWa5L/dKf7ZB7HsjVEC49AbDRB
bZgp8C8FlQ4nStbuRWKZdH6gIuyncgE0JI7RYqExmMPSepoUEkZkJPuE5C+qPEx+T/YMe5hOQS+N
5acVgr1bLW4BlDsaFilRWCFbUQ3xq4ovqq3ml0PnyZ7IEV6/q8LKLcbMWLs0XXS3bsHmSyzi4v+K
qfogDVqEcbOj1uiUPBlCLB+cjZAFnp6PMftWX3LKXS+F2vY8JnZHhejUvbZcDBDgXIvawmGFgT3D
UF89QurhXymWFv1kaOiIeYFf0P9gVwDnyIMAI4u+inkImY9xHOn0qxP6B2+kDcIq+Og2GX1OrFKI
eyasR6EK0xCKsrSNuVDoIAIOyK1u0DDh8g+rbCs3hBVwKl4JpfQvJ2S/i8ni1P0agKSrNb0vbWDU
XfcIBeJfOAyUanGzd+MOwJN8sGQD/aF+h4j2fEpn/vpwFtbgjwDBYfZLK5nTyBBiyyvYGj+Xj6Dq
1BFqNKZNWpTPlCjUJ/k/Vakx2tDZCx7TLSaHUM0hNp5yZGLPNwS0bxIS0qZ0A3tzp8p3k7xw9OWm
ZwFLS+iymmK/WBXQyClpq8AQFBYQJg5Mgnog7A6Udlm0z3By5SVrxQnth97TkG1e8sl63h6NFI6R
voM4YjA55kVTJXyEh2VPlFJ4mB2PvtH2zOE6nUzW2LQnnReUUa/sZX9UhuT91LRt0IUYuyrvw7Ew
97bgZvYugEQfExYI6UDBTd7TQ8u/0vjnxHCWN4s6kPWDP/jc3hTjze3m0/3phODkJMt45oeqpKt+
lVQ0zh0cEgL59IrZ8mMsyLkfI8nI66WxtYgIvJ+th9OZdk3WXZILC8rfj17I1nVncBynznxOX7m1
ABEsUgyDWUf9+eYw+KEIeBYvO5X3qi0VHH6nAdbFKZvcLiwFZjOqizugUi2ZscYMxIRWFTf0QhRH
MbIZ4huHns+lGvx/zFHto9K59jvXttc1kPRmsHT9ZPF9Ob6sUgBwO2XsWw+bhnHjJkTgSLCYn8+D
1aNRHT43wqdC8x0GfP5tGD1mEvfSqwN+ed+2tNsiLSqI4FZkqS7wVRoOHKqUaM+sy9zVKE1832V+
DbZC3BjSvInVW5ShnCEounocq3W8lV/LPilfOVzFw8XvmRl70Viz1IRh0eocP42rL8MLD7UNeDt8
Mt+H4Ol7OVs2nFxz27ucVg2IxAccZWLLCu6LEbaj8B6sueKQbKqUrHeUE8C9jVBov6Sgtx/fZ8Ki
q5tpGwZad+cCiwM1SbP25irykzGAYhyb+ORPuq5yzudUSyIrJ3xt1+aVanhK+u5uIJ4Wb73vC6aK
h06rqHGJouTLZDf50YYNISMwsAcDXGyoGA2A/8CRq+Q39MK03fTrlcHCu9bRn0aMvtMVv6oWL2vj
VPAjQ4PDkEhCCKmWNR6SkYT78Jb7gtZRLnhHOoSv7R4HzfTthcZX3j9Np/ESzGW5oJxraUMarww3
JTKLbLuda2QkLdBZsE8gjDMKbyJvbZ0GLSeUEooyNjL0TIYRFbx/KjEv4ycZ5Z7zCMur0Pu9hAin
pfnuKKrf4G+QpLO5whFKqmt1/oPoMT5JibVHdcPS6UfKf+t+dRGl65LvZanKqIv3F78eRQltMYnE
W6JtoRP5G75U6Y7coYpcEOI+Jn03GqZ6Q0AMWwGIEu+T/HlOkKZzWQqWsM3vC+xhEF9kM+OgKK58
WPa1A4OJ+p1MkGpXACfFp06s4wy11yHYIrUeiTn3kCoG6YAgmGS/Hdrk4Z4mA3U1tXUq/JWVb1Tj
X4GU1FB0C3KlJgBGSnrIM0/myrJTtI/eyf8/L2yiKC8u6z508sjbVYVg/Av8q6zOwmil+fMrD3MP
KITnE9hv4WDrro72ZAoDkOLXy4d5AA8K2hbxThG+oH9BAQnmaYycsXFPQlD/zdEFbNr6745bdHhi
GoMmXv6Ply+0kidRovZ1wJzqgJIsLr0ic1WolPh1weLVVnkOUveo1wPxMT6Ge6Wg2X3Yce7lmM78
7SVPf3UexaKPECDup2+GkmnaDzq11T+dFtw9I1QmeRHvyJLD2WuswIgW7cdUN7QowjaHwmrrd4Y5
bgcmZcLdpvAX1c19RrcnJqsXsrYgs9dxAKhQAtKYKDBzbAx44gnKmHV/4KKCZnARHt74vgsHelqU
MWBGrehMht/VP+4KbhPR8js/ViI2+QzRfuKgbkXEq0k3Qck+YYNai7HMWHcSb8WUje071n+OIhIB
De/rafO9ZVUa9yxt+r36VlnZpcIS0BWKsSetnisW2vcx0w+Mac2cFV92WfAZiA8p76yFwRE6Ux3S
5DIVp2VtHyxwT5BfYlRlrNmCnsiJoyH3RBz4BShd6OOQnAhyD3HLV/iwyRP4llwbApGxvInFtSOw
QT/mYRiGHDZ2YXDDtWjMY0OXxQd+nKDhCyXl+mAopjJOtgLXuzFCqRwwTcKLS3S8TbJqD2CnNLXu
M4Yj2dbYBqcD0yyHEjBFgjNajyGQPiYQck2H99MP+ytzAvECne9+Fa2JvVFZaQ+ROE6VeNOgXxFi
cDavOOdQ8HcDhhvlQ0AYxFwNNrrYpAj62a2bLq4MknWEjxSzBzNISsp7wAGQNuj/0E/wIMT2jKsu
Nre2AZL6HKF1xxnK3yYOUfR6dkZK9+LSSOeaKNbcMZUMGH0S58DbpF9Ihq7fqIdy5njeCuK03BhQ
ad9sdsQ/NjF6OT8PN4ULyYc8kY1EHJ6Jp0aQq1NOMBwVE+ywkNnMMlKp8h3nNtn653Ifpuvjw96R
v8LP042vM3igpI+HvBRDjBN2Jqt/h894QFIKgSHPim/plD8fsWD9logvildGZ9M2OhpErHQYtiTK
tL75yCzqiQBQ80DfFJsauZVbnoqok5jQ2Nlc/gi9xLGcy0RHY8ISXZh6EBDrV10LOsbvjfkMtt1N
GtQU1Snc927TsqJKpnpCIHiyvWCbixfmn4w6weFO3uP5/Syggl+SmQx4hhf82uYuN98GWnS04P00
6TjAQOKTdfopjfOxd69V1Mp97upM6tWTdqjiyTEf6HEvetibqbu5JySeNYhFd9NzyDnN5S9Eh1Pb
aTlrFMad9cd44cXKsoi6WaIynR5MfJqYpxw/uKhj5Gwk9XZ9J47Q0fXGIQSf/CKrc8iyHrekkfFU
DCQfDUcKHNZOlSEEx639GxNa5YwWpfk1AW9ZPQuUjNqXAGx/0tuvlFIplPC0lULVqPb2nul+AA6c
PWcg+3nePi1LUuWsO84OujmPFM40v31aTMra74YsNfE5hoflK5heNZtCs4NHvX94fvhX98XCdR7B
QgvtakwcZ01II/cyCy/mOiRHvKqlPU22M3+yH8cyAmfbpekyd5QDO7vpczDYCZRfzcC2Oxm047mP
mMRfTGTrh8Po1Jtym3NVYK0vy3GEJMnBTUY4uipjjxjv+l96Tuh48ebqUSKZx22y0k2byxUn6loO
u+8IwAi7QoUtPF5tlssufL2vPeIqydqrdcbGAZmO0F5zgX0jglSlSEPRKbwRKTv6NqGc5fpmE5sB
eDa5ajWoYKadtmqnX0kArWGCthhIfuAl4iqo5WfZvS5kKk4y1+X8ri/xcT/zW55vhGtLeIKBD/B2
EgjPp2a8rFgrgNHF5Mg9F4nAeNIxMLarHslUrPgftwlR76C7/Blt2H3cj8NN5eHi6CdGKIflTVXu
14Tq5BZEamVjyjdNI2MnuOCiaoQf0xQf8i812WgQlBTWZ5b8eiixUAoTE+6yI/dc3y1V3+aNKB3G
OwB3NhkEEQc8hVUxUszRm36S2+vpEd/vO0HBSF7ENE1ZXB7Mru7GGSKhUbzOVxMQLE956iQJqN1E
qXDAHl+bX/iC72DDHMCWyVltXnXPZEjgJjpdL6sUp5jiHTv94qQfaubFPSuDRUt740WCBITwBu0G
DuttILadaLFac29yEM1Bf2QtJsaA2leUm57dsmqU57wyKxF/8LxAQkcRpa0rv85guYfDb8utN3Ay
FBzEbskbynKTPPHYhBgunBOsO83So41/AnjsbEPwxAjXKIs1bS/OT7xHjgOYOWqSDAC2NN/rrC9j
2whnDpfdCS+IoAcI4wUxZAZQyWsGWvR/r8HrjxjRDzIKdu1s1DO9l5LUdWn9lzBqz+TFz86PGY+k
x1QOJBkpmp42x5Tme/yhGxLNTZH5sdKqRB7I5hRdnQyK2IquntlySXjHqd75s+4FPMimL3aOwSpO
Pv1gkylVwXRxmNB0w3f8mpsiqNpoXuNIhYveuP6VP647uA3dPqefZ8ZFYRLAUztHmLyvDGcZT7UK
UGQxMCSFrdfybrmRPbkl+O8KYYvPeAIr1HYQFTelu8n8jp0PJIU3ZDIj4l6AP7YPyQ5C4XTUMVyP
JYBDhHshNaFkZoxjf5q1jk58+J6yazqIIMG+cXrB3WjThzuHxVtTXL9BwDmvNETcq3c/gNN5iuRC
PSFv1S4KZhsHLoPV2wggD6eksfHcj6QYemhLG7N+qNvf6p7TtiO0w+Bq7zY7tNzxAflT7SNq/JMO
DUIcvtQhcFoJElqD4YB7JOlI4NkpxsK6w3bya/zN78IdEwA5yAXV+2cDmRVhm3E9CvyVwr7Wfsdk
Kx8Onf09sSubH2b2lLRnPm3TPjJiH+NSgM5fgsILpQCUy5TlB1Gl4tjdf+uUKzeceRpRusSz4FkU
K+QmbDsI2U4fGpry7c3BxOA+cvAubdKPB1/zDq3MifSTe7u7YaP1gBIxnU3nsPxYMKy1IpL/B1YH
qnENkc1dg+LdqkKZ3CdzuKP/QeXvxPuQfsfJc1LtjIysBKaOsc32AXMgTBdD/2yUkp7Ap/KiFCMg
ywyCPgHyWgN283Kelgn7wWEqFJT18WqwBTrddsXpZcGpWDP2qb+hqagXd6E7AHPnZrM35Ato3qoz
uG9TOIMBvNspMkJA2lK8VSNVUjF5lZt7lESqcPIT06PxOCT/5LD1G0Y0LoBaNT8jlF2L12l2nH4F
8+iPohBISZ/nEVpYtds2Dwmkhh7SR45tTiJ5HfvOcSfhfucTDoUrlVMHMGeMjfQzT1HEvjUlzWpX
nC1MHJxY2Wmimxp9vNQRR/6AfcO5lKJLv7QKUu95bNobbfbnDpGGnxre4zJwl+r0bYxRhmTqnFKg
YzDI1IY0yf8pnLUb1YTNnZ0QsZBeoI6itVCd8sPM29hT5E4kxXoX2PXhHW3sLdZ75pQnABsvQknr
Ja0sSDVy+ppM6k1bKaRuogxeEFOhCtsA53OE6mXIolpKxETpzmiGi6IYRebycpPP+20x33DsGNtn
9WvI9cG7thjGyHj3F+8HzMW26TpXTCGmVsEFDGgfUb2xPoPceO0u1iGav1/fOnSdO+y+Bk3o5mRo
HvLGaprBDmwj/9V7s2dy1+n10CXzEmxkVyqg/wsMqD6RxDNvemgpaiZgPe3MtcyItkjawVQjBlWn
0bCQ88usW/BqmRVV47MFVQ5f6ugtyMhgpRGyzi7u6jTLc/s8Sdzuo+fJmeuHZbC6JE6FcYYI+HPp
E2uFZN5JzPWh2H5YmgL6/eRWoJsj1a85ZF73ST0OmTeF9459uaIr/BEaeAy2zpmrwItQqUT553ou
DjKI6jo33IpOkgCll/ruxViShK1gmMFPLKVMxJ+nsAPkVPquQnn+I4JHy/0tnoewb+sQrorXJzmG
eNhxWNYo/l5aRVSeb0B34SXNlGtw0yOUU+zyBAjyEJ4rzgobJRzSOYVqMkSfeSxWUZHBFWJmFr7J
Eod3md3ikxx1K7t9xDrZQgg0TAQ5JSFMXZkf28LnauFJ2o67A7HXFNald+MpAyD+0SYhnNauSa45
Gk6G0TWj+64xphuyJ/l/hEXQi7/wpiCXcI95UHifF8VFyhqtqAwzBjAnB2JuChQszqHG7s33Uhmx
rzHOTlymEX0gSw1L6Z5p8QGZmU4J9RfTOOh8uCVqgmDzeN8mpCjLoKBTnvUQKjdzjU5aXYgBJF6O
43wpBv2AdW6w3b7nmWK8QoHY0ldvFWKQYSkaC9Pp1GbsbK3+TiYj69M/UrOX+uLOVaX5WEsKmyf5
o6XNtCCB+q7AJSrHQI7vt0n+vV6cThalXlcwZleU7JnfB5DdaYRm60dpqTR8vCJ5Q8Z/jHnvaSaF
cjM1sEpaZdH/tirUsoha72xYfZDVFLanxh+BRi+Yhx0RxrRm7SG6kSMTCj5dTsGeGFyvbV9rE65X
BUNgm6cu3FAIp6ilcdcq1XXCVykwA+D4JhDSM57y6Pbri6Qu3QiunYLGHhSdu+m/9vIoHjt2VoA4
2mkEBEvgUY2EmAracd6MoS/NiN2s4yD0orTlgpjHnuRqZsTSmzZ14TwWQ8mhaQj6e+j/byv4/89c
LXBPUA/jydLyJkZM1VOokZJ3g0xwAc+dIJ28QGjOHr8o7c8Q/1A+5SEwnNKu5Qf6Xni7JIvFekXl
ejaV9kas+s7TK8QYXH54nWBvNiVFj7xPvFStNQi0g634FyElHLBPPDMcPg3W/AvHp1BYjVHLQDD6
LTDuYN/wmDhESCEW8/ej7/bDR060AlsdNk7aVvJEbV5qu8Gdp3w1OP+eeIW0mWgTiVDAoHPuLn3p
qiz/mGWrdkuVX0szCYn+uJxjg2kPigFeLC4kAhO/+sU0hx5J+7315bJ5QKzz74di1ART+BNvknjq
IsaBjxwmOVw4h1oXZ6Ocs7dqoRgRyU/hTdCALGHMJjspSG2zrAbyFbnEBS4b4pqCB1yqqLwJJmur
2AWArrGRzCHptCXmE+xjUIycpRUfHUrtxdhcCLPNmOOaT13FN7Omar80du4CNyGmm7xONEVv4Ys0
0a4w4DHoP7ALJJ2eweiPHI+/8vJQuRWbHH+mwwVAYAe5mHzXdL/BnDU4mBVLe6M6Pk8wrRu845Ij
Er0WqhJWoN4JFSxPAZEUFctXDc9a3mnH8u1MtYUoIoMFfmjDqEptn4OQJ1ALRrCSE6qjY937yu8R
yF+KSNiMXyoOkdMcaCtTb8E6IFjBln7gyIGz4lgJYKQnc5Ol1Y4g4mPEm4CjhAWLQUkJhj7C+oQk
xaUi4yLUTsAUf6ucqdnM/MPSqcScpWjI2IysGJQ+iPihF9WMQjzBUz8H3HyhLpqral+Zms/bdlZw
StZAwfrQ107VxHzm+MTWObNLxFHYRC9nkCSfm60zIi60+9RRY5bhoaRQECv3pP2tFYKCw8tivzY+
QoAhdLQ7o8tvMLYidlsh0cHQDsGmCRap1XBE23FBU26ccIQmJNHJXZ402TjsoM9byUbjr8gmzdcF
iayppXL08NVPfcMdp/6zOSZYPB1ra+n0rCsrjv3T/nGhdU9TFwt9hSsKP9WEEYvKbyqtQAcL0szC
qzvQWtXlCK/CAIxP7cT5J39iy3PXHkT4uENCF6/ceoVI+vhm4e8M5QVQ01kXiQKMUaTVMn2JXUiZ
U3JPaDjwJhMqIiaOok6RFtNHLSv3EBoA8rPe0SqWPdvwFLWJq6xIau94gDEOSD1GOt1FlKmB+Xk8
De86e1eg+o5BeoCaZYDV0DR1OUSjNQ2pGoGKhze+5fjeM/ais4n6rsyMFyg+50J6AasUH9ehx0ve
cLVtISGQtuFVQQJnzul9c2kDGVkJbSrUR0jD3bgTsIDT/BX2UHEKddp7E5zN+62bW9Tya5Vulbt3
Ithukja3K6Zx1MZ0TKePbHQ2Xzp8k8VK7VX9UQ30VB87SYCalPzv/BoNpc4zOiB2zvhAs+c4kBYZ
h3no+yaDxR/YsbdIyRag93GfZ4S3bW4rmbMRRluLVOk7CltxTxq1MhKYCibtJDVny/179xPPYIYu
Kdaod5XOwwq0iTZZ/plJvQKwt99mELIFjdDgfgC/ywl5CaFqVlMurcqSJbgzEhim4EzkC2U91X5p
8Fh8H5MfJa/W0vIT3eqR1wCQZzUCGxEVNUHo447Xg/3uOAP42tiiUPX/raWEdAznR7LxM3RysK7D
jWMgQPriiskkDby2TJgfOikFZ/5ksnY0Uhv3OFHAKjCKHTSrcYJU1DyS8jsxuuqJt1ORdz6IVjZc
8Pz33hVy2pEyJSJz28Va69JweBQEWqMyZ76fZQUYf/eKy55SfEIlQVY3EmD5YU0qQtMiNlIeuOEv
YAf+1gk+ZwxATEmlpZHGID2KASIlcA1B7FOyen8LiX9BamNJiOATFLI0bi7rVZpTGSIxD0ecPzZu
klwSkTZLx0v9xJgUiaV6YT4gYRpO2qh+V0c6vMwzBMJytWaTQ2IOtgDxSFdGpRGs4YBME4mLJGQf
d0+weVqOCeUFSpxxl6C18Wot8qDj7Gl5FYehTDzdpqFg3Zuw6R9oB3I+K0uAPmHSvT7akFxQELYf
BTSW+nPT6PcPP6DI/EojisX3JBsjyAkXxuUyzx6lVnCklMabAoBj5kVvwNfMX4sMkKWyU55lYwJ7
vz+pxHKvu7XKHO50H5buiHO8VI4JvIFpqr3PaO58X4CL0rmlkrgtYWXTLepk+GTCb7UzBtQUQTVb
a7AtVzeijjmqpTp9e0B6h0enOkXbYn+aYPRlDcYc1hPzgWRcuds38mbzvqjCNyNY5EQjDhARfRhQ
R04SboaNchGGs6STludblhHuQz2syiaY14hBnxoAqgQmnjAxgbDC+ifSRFuUxics+59PfU/m+W2M
gil7aKFOpnq+nmCbu3ixgeFvGnst4VfdHoTOIbAGzQ/MQCFyw/jllrWUfSahIwr7/VfnEjc+sS/Y
A8G+YeYiA8sGcpgJKibDrn3s9OaYUyRSWRthCu7FsWLvMvgmEi0tzrlbYWGfkkox8+XpoFighKG8
yh/mcqZRqd+JuyxNa5Ipu7DuGvkgBuEv/cdEKeEzol8JpkQLPq0iCkGMWuL6YsLso/o6Hy9n0uKF
JHolKV+xni3DayGKY2/E4DUc0aWetMgCmojGPeghkqRaeCOeW7St9spoEGfK2c90iKFBa8cs/1tB
9GthqueJ+dQUBKwE5ttbAK79xtzdDHr/o/2x97hEx6aUnLaCd61ALJZayLz9WHIEnQS5OxjpoEh3
w2fpAwuhGZkjJS4cOQ9Mq1l2TLu9Sa2w4xli3DtzpnuXDeeFZdoaXCZifQW0FFeczAboP1qHhzc6
+BL2sNFhWEcPBPXAsmm+pkH0bCZxd6VFbf6d188TJg6G9z7Ws5uWOJ660udoLsAOY3p8gXMz9Yqq
yx0MbEXFKpokRURFsFs4KaAFHCYy6NHTut2KQ4y8ueDBFH5SDB/JFOh4QTckCPrLIOETPZiePnxK
m03pQhv1+Wako9lNZUT2xIuaLEl15qe55NUKLNU1pYfjTMgzZQzEmVI8Nii2w+M9dq/De3iO9YSP
208zztPHGZyXeeTS4yb1DZRiYRlTnGkHudqjcdd9qkCw0vbPIxz8F1Ddk+VMzY8mfUMeUdnoAAC6
8tKEOSCfEaYwaJQN0IYOqF+Ta1lUSA6c04mS3s6x1jSZrRWe3uRf71HjJleaQnKmkhmCRSc+3LmP
tumH4O9Xe+A8vPHpjipeV0FtXZRcax0TeoCZ06HjRmKVSnAHr/3eXyagQ3l4nKmK5rBD3UNTJOQ0
pxCelbCqbQSA7eQlHe4qu7PZsim5oSujgDP4nSuixUSKqa+BaWMqg+V2/uhhqd2RCRuqIRZT64RE
lS4EothxdBEgabDcBug8a6IDz6lPOxJnAUrraeNJo4ErNuXCQuWPQOCxixiRKUYHKpDHOVbBHgAt
rko/qaw6DO/Jl8xZAUV0Wej5SfBRhA/jajq/FB3d8AoRxKLZ0OF0eCX2VDNKUIudQjFAwnuTbprK
8fVGKxZYzURavDDKGO72amXXnqBU7w1K4TkfGufubDLYtoKwaGZgidhNP/vzjQOG9WlX2X4UHeq+
UDj0zw1D3zAn/jRHiMUb3pM9Ewe/OCEhLFIVXrYGx8/lYZHziHs9RqQOtPkg+9TPDekRDoGJs5QQ
KhdzB9Mj8tVKhm7qboD7b3028oV+dxByaFBQepkssV9ntqUVBmM8TpfHSqsYASKNv3GQvId/bhyO
xojbPI9VNV+e9fuRVOqw+3V+GEEx/+ekQKKesVyQOUyDdlWPTkKcgaK0ytz4GrcTsHitlaVf5gto
G0WHaLy7LTQkoraQ9wHHXsvyLv72z2LtAiHEuIMhdAxFKyUcCsFgemfSWS4ZtrOO7qKtf83hZhCr
R/DaRGvXP6kptH68qtfCo4dQIeIS0RxDyoco59Wff8fi+zxFq5tLWTAy435ONML+S9NyWHa48j+G
tpGVtzVqNVPoPsBRmc66tJUTvzbMNtSe73s0WiF73FpyrvnRgARFpqc3p1TM6k7YCsmHZnJ+xlLa
2KC7WwbenJrmyFdcu7xz6JFkFPQF2d+WF/2zgFnCMuQrdNPz8OMw+U0mdRpf4hk0I+SS/7QV4S5M
SxvNKLzmn74ClhX5muBI4cJfLOgNJrV6qyeT73+EFxaXOcEEWI3Zb0skv786y9rvI2Isl/nftKoy
1SnOlYKGEpvF5mdisf0k9nJBOVnQuKkKXukaTafeXTpe1lGjNtfsqWYurG+2z6csoYamaHUxGVHZ
X00U7q05qnWYd6zlaYFPIaA5DDUSxkRp3PMrK00AHyGtbPTcVip1QZGnIrYwAZNnhV4sFn/5mQRz
WP+vo9ABFT7UgeDT4sghzbKLleAbGdYyUpwBxEBvi+gioCG9G4CNf6YCRCuYRuDjQW0vM2Zafn2M
jmjfQAaVvYkJ0PVB5cWKNiBNxUuq4mQVA/wDeA5Qe6rK8LduCZ1B7fpufmsnJzMjZ9oF5NHoK84H
SxuD+iG07rZk1pyFb9BD1BkPeJO+FXgNzRqG4mquV05hzEi7z6EY4tD0KK379jl0cC2m67c/BOOt
TLa730dumgA4GAHbc3ewEKh09bOmthjQpvgOZtSlIoyd4yY2S15y6khe63H2kgKaH/T3eEJChaAg
UjhCx2CL0G+EMgMILBZKjt9u1Ted3zUFeuyYLdKGlS/Y1wmTuqTwFDE3qxnaUThCv5IF3d0BQeol
cO+bvesFwEV2mFct7Mzia0LanCZ1J1URIfxJ5zp3DeM/8g7vr7+oTfcQxmiP0WjeUDABIKS4JQG8
lNUdMNRUuDjHvsipjMeyyAuP4TMXXRkzk2CiyT1d8+H6iuHRgrDALTI52kaCaZtCPd820LJxoyD3
87fjRHLNci779pUqLtCuAKl5lwOg/ux4QmsQEPsNtSFbdqg4JJ7jMPDPAR9M8eTCKmU75M7SCdO3
40FOEIlVdDJGzqIvdrJPN3U8NreHnMydnt0lCM2bKM4LoR12Mu6mu2KAcNe125I2zzXlpZMVWpXd
KqjpscP8ZNXRaHNakYcsvwSjDs+OF7XImegrYbECJuClVq+j8kLrLsdh86/fDq71OT8ToscFa9R9
g+Hld17P7wUSQh4PcEeilO5/ihbLODRg7miUjL7MZvsYySqcGtkQVYwfVvJpREpN3i2oRqeBXvoU
+PRPd74RKJ6h1bkG36PzbOm3Ji/dBN6zjI/gz4eN3valltbRCgPuRWwx5GbwvKSin6zk5i9G5xVw
iHLUcc2HtHvmKJEac8GrKyCvBdmMq70y/NNHfpabiGtz6WdXo2GzebE0Db7AJ97lwYAG4lYZgs5+
ZE1U3F9NX3v8JLko33Ykq/66QVFDkg3Cozl5xiUjaRjTAkvRYGNQUqPj9tGnezN3fLISMh/v+LFm
ia9GN47knPQW4rcia17+UD2R0ozk75p/0cxHPTJTlVTclFp2g3LNEyzIB2tsu0Dqv77Gh6mOIJ0R
0HSJL64D8m1KcHQDJnUqDGRbi3FJLlfiZLmyYke3iJSIbp4a+LhR574PlfFOvUzAjmqlqZWSTVZK
x87KTboW7JXMbRw1YcVL/48ypfdlZ5NmhS+KfIiU+LC8u3iZlzYZCxbdUtBi34/6TqtrKNSFW3BC
xu+kgg/NKWUOiCaNClS98DE8LAyvnKVmamzAEx0ObGH5qXBC0yYVZ8iDhlQMhpuzgpbOaWPYxYJK
kxWHKhMbUg8SOsuycfYVvUGQyoPitXEbqxy6ryT2AswYlDKOgdD8Nn/V6tMRmucQdQJ0IbH/tIj7
EvItURIgEKhNGLLCYuR354X/IA0aBEz1oFyyBAh53Mao+fGhZ+N06waqishJ3dPtbK4OlhjmeTI5
j/u3mfXG6m3jpGotxs42MpW+k/cHQDkJKc71gduTkE4+4OYngIorCsQe0KrbCqq/1D2XozcNqSof
9Y7EFkFozJoxnrtY2cHN8skUIFjaKB/kqa9C9AdXn4/tRKbP9WqVm9FcZhTNvff+CkBvzxUU/l5L
G+xpL/upurES3VQnhVwwoutecn2Ta84r93FvFwGy+nBpxoaMgaH273osTee9JnQmE2WlKeO3X13w
KKac9ia08VjyhstfBZdjJIiEkkvNO83mDZlJF6jPmHMIWwFScq0C03CHSk1QdE+BeB6wjEGlO8e5
1yd5g9o74NpTz6IFIt8lOWnbpSNuKDjXLM7rrdf8x9Wm/y16anOwFuIPwz7UgP2xgqEA8rLXy4i4
cYpASOWKhA1JvzN3/qQ/xVJyf4jN6MQPguU+lRAxbJxqmGXWbvD/PKdF+/84HfiLkFkTe+1L29BQ
Gv0JgMj3QJU5iMDUFVtpmNs/0sBIDGB/I/dAPfcUmVy3Wae2DbMW3scW0Xf1EuOs7Qpfez1Uedat
TNiCmBe3PnMVttu6If0tq6FvSMX+PPsAAx8VMZ5MmtI76YmGP4b0YZ8woBCycfACcBPT2RoYXnxI
dw1rXNMcGwvt7YNFC3Sv8rU9/ELt6ymwpk/w0vVdTjosRtQ7FvT16mMPsSoI1PwgSFdecf8EKIzk
Zki9jeWk7lgPvu0wjHxdpSq2gttNj8dEWwm+rUVVZuF5M3A/FnaISghavIIS2MRfXraPMaMNfJZg
dwBRQfTrfMp2oQ72iSBXFTjf1jvspI68RKsBG5yITMjVa9dwa1r1UdzsImuNr1ojjo1UvEs1E4p+
MZrymCHYfO2rwbXLShsP5fSmUJbVwsqVaqQ4vXtH28rGltHfNRFro8bXiZAaM15vgNiYozz0taXj
/FZDq8qlHvBVJ0xmhaztwUjg+DGWFCVuaO0DN0f8N3/XVww8LW8r+veoyT2+5t1ruO/rEq1LvUXs
bCV6J2uFa0GHHXfyvtVGtPnzDM8L8h/UsfnYe3n5GjIQUTavPaXJ8IWBFndIwlrS9M+K+iJnQU9P
tjBKt5SAZPnM5PG7cQvc6YXcttE4e/uqpe3OAEuIErOI87xmfI8QanEVGEGEp6Ph8LEgQ6fdg7rv
R9FHNakiDDc5m6pllFgLKnP9W0e3gXY/3W+yk2uTNjX4CYjoHz8Sc+ZhZ01wLTrTjMS4WRFAOEYb
p9XvoU9UV6k8zcu0QS8dzqLZ33eXe069JhbbjamkAQiOpdkIIH3RFP6NpQAgTbyFHFMlJEhM2V32
kVx8mvq17Ed51IcegnBqoqQzLH5DhB+0N9aQ/rkusVxjFM/hjBY1T7A3Er2FV6+GIzSkOPMQZQLE
76UmSQprKZxS08XwwHPWiqR1FOVLcaN9sy8UaG+rwb+NdvArBgSNoOxNAdllOIYbwOgmkc4/GdmZ
iV05cf9TQjU9jXBmAYoPV/rEZqYjTqiaXhrvZvDkkJaLSo1PQcer2H0bM+hH5peJ/ma1hkw0IvIY
jdVPALRmfJVLiKwZVq9E6GdGr6KgCs3kutSuEf2XC49Wcrz7U7HVzYAo/7ncqmeyCo268YOTYsYp
8coz018GnHw4QZBVKpc72PZiHn9plOCHbVooPVc2TAz9GK6or0kzd40GSWs9rBFNNHRAgoa+Wwi+
hCGPcLCffjgDBWLl5bzpqNbhKW/4/nKGULTJUTLH7NnmcYSxni3XYjXHx0mZYl7Od/okQBJPkLeG
nQkZ8VbbVz14Ycww6VItMCUAGTo8a7NeqNCnd2d7IhERAqEYSzKbZVqRjuHHfe8kA8oY2z/CmCSx
jR5Z/8J7J3aqxjRaSAXdJdGPGDZEAFge44dbw+0gWEnNtofusmT50zVLQYOhaJPT7qDyvjr6r/Ln
Vt1hd4hzJdVIjl98NGAevD9Mm7wAwgKmvbfFyzb6OHAHv5MrtpD4egQYS031gAKRj84HTzksE6JV
aG+3pbL3L2tRMBCZr5tNTUVPGoLCM32s6H3kaPsmbKuLc2DPh2rSADVWOxCj26ym8agRc1WCTeA2
jzCC6loVLKpB6Ni7VRT1chup8vvekVfqLbGP4W5IEz/jsXRZ+FthdOJ6zRpBfjAYXrPrPQdpbyZ+
eBd8msvGWas/LW5tlEqEZ8v1EULdMqDf3qOTWqdIpQpvzF3zLhD3K4o72tzbz/DozU+dxzQMNDYj
118iswVHYuvcPcaRT+4RzgxP5yLKbaODRCXrp7TFM4x6s/w2u0voZ6u0rg+Jxe/E2Mqj3CG/QX6n
ru0AtpYzSy0MQjeZPXLd5YUKSUgGNdCUiEIPCzNaiqzHzU4pdbP9SPv0LKZIi8jIKxteW3bLolQv
dopICq/SbQ78fAS79tswCdACR88Wu0DmTT+JxFZ/yzj2oTraAXtYTMO7hVCZ/5UswkBYxBypknHm
p1cd8mFUiiVRU7n/2Ix3tQk8hLWWHWJZ1wV6omKkI7/b22LOzS4O0AGeir5em0tNhsGtTjLNkg6j
Jju6P7spqEsvgM0UeuPFXKjHTbQ0PAcNH9LdzOH4P3q/jIb73PEiNiJtDN6T+vbP7saBOOPtQhxQ
Y2VqrWIrdNyKXAPSz5TyIpOB3tEFUJzjiyzKQn1JzI/jyBGY2uzVrUIkQZ4ef1Za1AwG2KZdKaJ/
Il/t/B/6Qv2SiGUUTMGX6z79ZG2PvndK25+LhYeG1wBOiloxqieEXR8B4kwFdSvWpBHczKTnaafP
I06ZHW007Y6JA5dWXSyvbdJp/DcjM7AQZYBnR8fSGE4g4TfPa/0x+WuoSYVwphJxl5uKGHBMb9db
zU4bXWL8qV4d0yi7Y2TmNKnUcAZXKMiBuBoW0nreXpA3bZrKvDQd5TL4YJbxyjBWRTjOY6Bikrkm
imUsQtmdY/BIkq8BHKSaCO9WfXejDs1WKswKhD6AKz9irlJNN33oOyZLIt1x8TTmdxRGMsslnz1U
tXE51izvMyiP3DvwCQ1UwgzmGqAcWKnlzpzTIW1Ji4m5A4PvOMTvO/ImHgb3tbMY0VhWOgdZbuD/
6tv9INrc1rLeFp0eDr5UcCXCmIw5kdUtpfQjhWSqkbz7NnsPSjZauIoXUVblYwNUC+ckA8Jvgyc9
YK4RLbkytJ6y/ZJV6bZ2LBAcsnplnFCw3N2MSR9eD+gwCcuVHCpPalkqQ+T4gygcqWWk3UYFjzjy
yTYGWdSJhtBciEkQSsWSGoTgDoriwS5Dvhn769zaJEMQfcz9yjANQDFf3Ryiv7pJ/MzUMJH4wHsH
mgLET8zsYtfYLJ7EFYbsrEHzqUHh+OWDz+tF4AXSFbequs8QKq6ES923VOzbNiGICa+Y4FcfwmsR
Q7Er2V+s619PEM1i1+uPdu6EQNH5E6M7d1f2WNdnOj5WuNOck4AfWoOgCTbefVFZcpJfW4kj2VId
UE459qs6CjPVTEYGg7qdA8XQp10J+JwVFwy+Vdki0JH8KhSwluQ+HjHltuJ+oxR8tB8zXYyo4PM+
arsZbuoHvliAXqFkxYFVDHn615IO3j0oco2JnRCaSBiJ6J/w+3rFtPjI5gYbxea7v/QBXLVLPkcE
2wuXBRiPy/22KcyTfHRU8sai5jyaVIl7RSuzgU6MIs8hRAFbE38rKHu/kSpipskF9zZpGWgTSdck
VVBqTr15C6sU5Oxs3vZnQHylPCjtTBY6R/j/4hhlTxe/ZQGIX9CTPGTOMT+dIIgOLwg1Qc+3LxtT
1ViDgiF1sey4HfBJG1+4MuUtfhoH4zB1Wd4W4ViEkVrouNhWn6HtJyHfRBPFOFsb/8527buaDERa
1qpzsH/sX+92ge9iMhw60zCWVWndWkDMvY1rQFQSaYxmHqSva2HBn0sC4CeGYBU/r376Vhq3LzVO
8l/M+wlGS7IxljmL8nP9R0OYolgzm7YwdQlO3qXi+BJrkTzynXLfHhph/nFomalyVOq3ieXxB1NF
/qcd1axU6tk0LhAA8cyic9vSVDZjC0V8pIDcRfqm5txcxETUbrBDt6q0XqmiCUSVGFtKED8E+wKK
5a3ZTIW4K+1cZPfiHBcy+z7NhtVmJD/Ky728hYNoyVhDcuyAx13l/glQ44bBhp6WS0Mjp540uFBu
IWdalI4bwke8P0IMYBv8yq2jYt7gdgjuWrvKvwZDzuQgnIdtrTRQE6mzwuSfnWfkR2XvLgcdosua
nPhOaL8v035p4tTR1p5J86BupPOfBACscichJ19P43lFHvDXkyM0PvEOmBYUx2V15FjCB6nO8rV7
OTofyIbL3qaZ9bcI5jdisSt5l/wybLUl1ocBitE8kBDJJUkqayp27OWg+vt9Vk4R57JXbgsJJ50/
UVNy5BIDlzWZX/NGqbzC62x/q07aDEvZARB/dRZb9+f8qyB/pk/j1uUTm3sx3bgCDEX5HWvr5Ald
wEz0Fr/APXupgfgGx10dH5rlbS+xRHvYzSha6GYJGPVeE/cl4F8IpJ8o7dAz1CuVWANhRHx9kAGG
EtSlMNIQmTh7h6LeSNOZOESHFt62694Y3xpHo/cUCdwKdSl/DrLHGMS8zQUJ2ksDx8shqwP6GGRr
fRzEc/iQcTjQBHNhojkwxUyx/DZtIezS79IJ/NEOcmjujx3WZMHC1IYNbDjsudkoz/cTpQfUwBYf
tDN02GxwsDBRVY3Aq510JHR5pCbq0c2gR1SOiCccDk2b9kYK6kvEvdB9izdL8doapnkgApOYAMs3
BONewVl7LvR3YXfu31lqAOlk3/rkW34ex9VfpGFO74WbgrNLrKTqt9X2n0Hj4DImpcsHijzUsXU/
m5LzVjnFTK2pjH8QdjO33It3dH865rYU3AmTrk1JqOtya0R4369Ck4Qf8jSCbACHLMRQmgo9rRf2
I5bLUUrjzZgMHlckqv/s9bBaFsAuG//jyfe8U9axxWxIUbJir84WrqNc+QgfPB/Zr/DxDN+3Rvur
xiJV5Ij6jeZ+TXrlG8H3ZgcbAcAmMlYRizuP2ysCt6X9DReUKk3y4Gr2kO11drvU8OS5OoGwfyPt
AMIeKRLHavwTtdbIH4+k9cAswd+xCaaXPKL2P/LAaJnalPMr08E5K+0vHY8KMBwxLCrAhIRv14i7
qejGiKDkE4cwOMucOsD9j8tnSFzUbQm800FYUh89Ky4dnw0jl0V+QrQY4sLEhM87Kom84zCchvfJ
1jzQKXexc1cG3lTQdp/vsKWqDuwuLXjtiEqFBAHYoiljfUAKBojOh0Whv21QE7jkhgjTbjJ6sjjp
xC3iFNp6ngLXhnqa2LYPY9VxaqAEJFTPfjVbUP73faXZwhHqu/opanFfb8UaCnc9548hyFK2Whvf
vFy621fxyJAlWZqwgbEo3gYAvNYzTGrur407MIcK7FV0HEYklo6t6ilrxJOxK7NW1I6vcbv1BmsV
jlVlTQPJRVtSk+Be+1uivFP4+mo++WM0GxE8BLGrY46QtxNigmPu8orE8Mlx4rCAu7FXQaQryA9m
cl5n4iTXb/TySO8sw7UJCqEccIqulMGc0f0qt8zGOl7uiXFt3snhRIzYKKCoq5/0Eu5gkB951XxE
fnQlUqcLkoDtdFE2lK3SYbHwkzn6k+0Kb0/7s41gYbAC/RRRG2O2xCwb7mIxBNpB1NhXutIUu024
7bmLrShqJ0h1tArztnM+y5UiBJcWDXUoFmNbdZAG+rY7QzR1oDadf18PT7Pbri6kqIXcBLwCW+vX
6YBJl+y5R145QWq08/1SwylyOXPXBA+HfkURDBlLh+K9ToiXeKTg50pCWYszZcQwcCVZKm3hTQXt
4EPCW3d103KTRIYWHVettrpFqR+jNsHb03bM9XVJQtOv8lUZqdqkXX8cBzmYBUsg6Fixpe5dpHux
Xdq37a0iRhdbpiRSmDMNHAgi1XiNKs4YXRdxcQuI7bo4jMqdv31neeIzq1/0/UXgDKLlAAkONJVr
VV+HjtZn1SUMu7u4+70S+3V8bw0hcELm421HeozPfsG9x0RSo3ZsIc/fNnpsItj+cWDpN0CKYPep
/TAvrLIOBouNgYO7JjHKdFkjAutAWuPFaN67tj2PjqxPx6O+Qoqk/hOE9fy+fGslUUGCqOls0shY
d897aEZ1RqicJ30Dq32uyaQNCt/dV4MqrypkyzFSUtqzjgthR10xS7ywOGXV4N56wC5LCELBLAJr
m88ZJcFn6z9iV0fGmi5GBjKffeGaAkblqkzvapY8FDSk6JrPTBCBNoOhDsubeUB5pNqE59fE+7k6
LW/qZtpGM4gtA44a6Nm58m2QVUemYew6i30E1+/TaE3DyGi/qTqgYUStxOVaBoxORJb9vKVZkkuh
kdJyxtlEZfgsTCLvJ23Cprghq8sLV9OEhacx4GrQcuhBlGtC/A4Ogrql03A3PBPIsqtDcwyyHRVC
JesLbOzkMOF9JFcOAzqyYX01Mk7SuxjRd4BUPtIvCggGD4MxxbV+YYYsJUUMPLK00gkMz/ZPTxJ3
h1tHvieybmUpFkAh+zaUj2ayAOuxZobwe36wGAM2FdBsDRWrLzDILejz1u1QE/dfRLodnIMO6D4Z
AFHsKpdJWGhc1VxKbvLoL3DdXvMukQkoTw2phMUBUpdJRY+bhTP//pSzlKlaDoY5nrfqwqbZqsLu
Ms7dDPM0pPyiMQ4/Wlo36x5PzKKMJ7x6gWR/bPsUkAFIogFsP6x7DEuV4DDoBK3Tw1NC5c/0nFwr
IaLEkW2vTqlP6P53xzCIqcD7O+KZGbj+yGHsfyR5UQXPsvTttx78uNnHLWwAtYxmNUpELUPifVne
cA4EyhiZd7UpfMSfG95dNXSd8/E4343eGnRzdi4odkRpoD2zXNLxAoSxK/m7RXxTSnRVv34P4XnY
Y+xb4ZA9/8JUN1g8DITxy2cPxUWAJTsxRKrDnv70PDfWVGMtGW0iquZHRuRiEDhn6U9aoAmIsINS
MujCd6z2dhhUSrwysxQfx+uVzQnTNRW9XNeRP/YQmbgf/hZvo1Z6XMLWoV0CxOR5NNuatdEea+e3
hxxvzu8FqT0tsxZS7hyK8yEWmpGD17ZCHOgFKv02QLQYtPoEvdddBqtcR84o05UzXM5/IWA6M7HQ
xj9I2WcLay5Tg8KAN/vdni8ZxkZAOaRvyuO2vxjbn9QJoC4AIMupGzEtL4wP/SMb50/oKS9QiJbz
qehT/FaoGo1SAmISALC1HeHgpiOJhB0plX57eVa4c7eKhFSmKtWl/50f4pc3YHZoOnmw/Dphcd9t
kjgA2BYolSLYNheV3er3cf0kRdXggZombjuMVhC5vNrMvtWdXnamFPkiR0/icHTpeZd0vTF/v66C
+ETTApj34EcHXVC0STnC5b7tNrEUEaHd6sOwZRCTe+fE+pnx4icVhoyPwOAvmBXNYsn3cGt04wrt
zB9kYANgv1S3PhWEFXzvNwOfBJ1vIpuEzeEj6opcqWh0+qxYBAWdCf/cDUESVnmiZZRboFgg+bSN
UKS89hxyQ06CiWY/kCm0xS1M7dFx5f1a8rtA9YJCX0HTgD9xKpAr1lJxy87xSRDkg9OJV4p2jnNy
aGBp4LbLMw5vBMt5kwyS8e35trrp1aU7rliIkCqS+fB/dZgVegIKPcFYB8V71m7wSGf0MA5ssZ/z
yuJHT53Zxkx/4v3NraxHpSmxWWhkNCe3n2mQMgSs6hOaptP+gO5frZL6bEjjXkpXAqYVNDXsyNSj
maiRlKXUr60tyneNmYClH2oX5OT7BlhoZr6jfQIztc8FgZBpHQM6/uaujCKls1hRAmAMfilghQKx
MQVgzH0NoVDRpQQSECEUy/L/5G89YIMU0e5wB6cVdTBEjcEet81oXXIxpc1lg198pQyzyLQ/YSUz
7mdAh6ewriZOTMInmGCVgk3t+Q3E14Iexbm0UY28i4grcahhamWAEaDlubJdnt4Box4I4Kr4CbEn
C0l9weck2yRAdhmhGs2IPWoTeweeqcMohBAJvCRl98PvcIRzlBJhfoiTHy1Ab61+ZTJFoAg/j0m0
1N4WYyhNydP5Pz0L4nCQQIsKJ3yQvgxZ9HeuCC9SkKEGgzMvgSRN2B6/ixXF21dXW+5L0RhCHyNw
QHJXrotC6AL6y1mljfFudYD52gq7DblbwV2hpHfwCTyYGBe/huHr4qioAjrZCwSHoxzQN/8btUNb
jYTSnvc7/E69KBr+s3x7nz10ifiwbqGD0vlDSNK6hEiiXDIPc21i8ggDAsIW3C1Ms2hzy3/t5HwT
rVNwrGUGfOn6wuPXnkrzko7ZKx7um2OLusgP1MA02xoJwjFXaXPbUNiz7Qn0vc8laNjGaCT0Hdn6
5bihe5GCp9+hFP8X7ywtF2HUTOLY5hI512TwvyOX/if65w3CXFm7y/i/e1TRJd5rI9omlxLiX/rr
utL8UxzDC7MA519ip4na2SJEtnKg7QfMpvPbmRgAXGLOrHruo03WZyb7iuWWkBu3UCf5QQbKEZFq
w48A5ydEWHFuIBM8SOpzZlFLR5jb+69YQFOQCJtweGgHcGUW0qISDQP0zVsirhHJ6lCl4uihhuuu
OyzHBfbrnswO4Ha7rydNC8OmX35MLHCwX2BqtVyybD2f/LvWxLLWSQ1Vu6XLllIUD48t2P9LjYJE
pOsKJH5tIk6L4KBSX44cLV4fAtRUw55/+zgfasoPAvE5JakehW1o8BtZ0zFRyccZLRTIaFcOMLAd
oDdKrN/UNiZP4sdRnb0oQX0tkmkxaUqgHUpN9VIquPMC54GGoSdHLA9JsHLvThMQ4GWg2zMuZlCN
vkSToxJTw0KCfjjakVAzndxvDyOG0bvHDQfpthbDPsnKSXhyUmI4S4q2Q4XdoxLq77D6KVbpez5b
mQl9B6QcO8ndgfV9L863isnLdxMOpLLVQ1craV1oYhzTFH14tPRzq3ed1MVOP54551en35g7GGLk
oTmOLYvHdoKCFeF4RWVHNxy10cbcYhzIvK/PFE5DcKErhVrkhvoAwElRPFCUW15wPaKDUOBJTIqd
3kPGzK0609AqzT+2R1Zu5QpFQPv48xJ7xlFzL9C4k6GErkk4mSY2ol+pgQO/0A6RU45w4SoX/4c/
6tqd238UNWNBH5BpZ0rRrGymmJFyKtzPKVm7ybT7Tj7nB3bU1ojIN2aJsG4JInMIkxPqmDchFs4i
LVGRx2R72jAbPCIZti/dtl9NELr3OziDRpTLV1Akm8wFh2C4PZRLGa9UuLKmJXnzgl8VGD1Dmp2d
xm4kDluUg+wM+udNuao8Nat2FFBlNpGUo2CKpq90zDsBa/mHQwRwD08B9X2QgEKoa34Kbs3lqc8u
eptyfS07qTGWxKxTnrwTP66i9mXukUXFaHJvxactoB8J/YauyW7oak6D8dQDMASSnuy3uFRrptcr
CDNRv+9OVNstn5/Gb9iF/MWtKHe/SQpAEL5i1Nn1SHdrHibaCOc9QiDoNNj5DhenUvPiv40t8oOw
GVed8z/LDI3CmKckRUIYfMMo5DY/iQaAeuPjY6HbQyxoaDyHmECibBbIyx7RjrimhMkBc2w2nVOo
g+1s/ZHYYMt04RSufbqnDHAiTLcelsitKMmrEleXg5G2D4vNLJM+1xpKLKTy/OSgT3LRvRAmaXpE
8dQstm6dbqVhRrOrMMDcyBdTYl3JovzDBxAwcaE/PvhpnRAm1FaT8R8KVUtOO2QjYLXaEgBvLnXv
sLzqNp1xVHntIAzgFzk0zCdrPXQFmqZcXvntLbPyAcw8/2VIhyMintQDLHRNz0RwQSUZUBmcywSB
QN596cudcTkz54UvxqxzbR9u1UpPfJrCCrQg2WNhAj+OIyeMihe0wkzn//85xT8lDVL/m0/jlO6T
1a/m1+pacavfIx+7FEtRfZBRawrgnnj6ICsmg/aAc/MFNIm+q0OxuhNTnqTnpVhpBUdEH5AiMIxg
31WJufHTpsFYH1dhsxPtngI9NIZdb3Xue5GufxMW0QoTLE+5ltMddp7aBfmcTSONf/8ERDK46mM3
k/uTJegtD5AtbCmSfkN9034tFhEomtujsixSTXrobAtK/yYJxlptlxXUPj663G0BT5cKLUZBv0jQ
0WCZcWdA8iBN/ish4DefndOfYxW/J0jHS1BiO39Jfl4rYJDZBEHXhQiV72/z01Ue278yiAAcpLNG
mye4bFn0TEHOez1xqCctzcTn7W8+O+A8DUIFL6SFpFUO+7QXIyrBTHH2KuCDhI9ftnLtUXu/Lfcu
PjFVcv7xUfRf0lCgKnca/jc6AIszv6hkkdgvb1/miOVV4tbj0dCzXPjKk3NrfSrXXpgGqjb6gq4B
TAghDOeUfMMQufzpz/JgOonCoJAhIRAI8hh9ONVjNMvJiMgDQELRncEGzO0TRG0Ez+jbtQzVtznn
ziZiGYIywRVUeiSf+ejC/C7NsNiCxjdOPHwZT7RmLO9yEALXT1bbuJIp3Z0qE5ADN17KMFq3rpMN
YAcrUpDvegZt2Pi/v8d0pRxZujBqGolmk+u5e+JnZTZHpUTMb+WlSKPvH2T4RpHALIHnINbXsz7Z
5/wQ7fWGWly3AShrb9PhMutJ8eDjcy0loK6qXIckxynjZffUPbXmyBrUg69nhgv1wwDODYvrIJ84
Fc8Y3dmBSfoytfnyYOIrdR06DlNJ7IK3igoADP90kSE012H5G8+46Sf8HAinlm4OJRKOcfg7l3Hw
medZZKCCIWOt8MKXDngZ+BkT91tsNBJNjVS7mAXmBCfipLj/fK+u8rvmyMGKtQnSpt/06e9Y7Lj6
anQTKIgUNKaOHj7tpOUXO3i/Zf1oIVFrhVLEEF26bGlKiDUZ44fBcg6TzVxNhZ4WSZbD4xvySF64
AOO01UR2+mSGVvrsSVGqdYlKB4xUrxX9C7+Dl5qS8dllvVOOx1qEmq+uNUaYgbXF6Y9mqB19UZMp
cWEK/eRFqqbjPz4G1KkYf6MoNcvoZgIEkrqWiJzGIcPdHEqFaoezu9OQz2p67ceKFieD5SispSu6
hsuxJadJ4v9evXZtwr/4UNQgJKWF0mg/UIhu0PcYy9USfCpSXJunkfzD42Mqcfkn7jm5G8Uw7/09
H62GgeALTXJFm6dObjpYK9XtxYrU8YbQeMxknpiIDj5oFgzazTFUcolyLTBQzuGwCK2vgMJ7T4PQ
IL8LT/k75GLfk4oNBJOD+R3LM7dnhytCwVXNkxcDk40CUqbik6jxMOSTPUMLbGHcgo/jXGgWaiMb
zUxIm9+nWlAcyP4Exab0Djae1rjRjST75orm5akPT3DQ8lUqdtg7SkThzUBPRXPXpw4ETXRHyX+3
ToFXMPrI6Gt2PcIyKJ7nOsitbNoB9yhLemZgv0DgcId9EZUMUm/jSEQBCdx3hT4QGMCmzivDKmoU
JlvFWsAxKcDGaDf6r2o1sSzprC3dB6xtw71rWCmH9rZll6HmgpurbvBUird3VnTfJx4AO10gSri8
e7u/JxE/RBulkX5y6Ix4zP2juVoFGth8oww1Jky0XXzhiTaCdVDGnYL3QT9Rsw0R8k6sjGmDukIQ
Jb40r+3z1IDWr0Aze/DvlobA6ttnJIGK0JWKRKhEzSGD7mqoDyi0rUjiBLInTnynMuRFpeEBNEyW
7Os7peaa4mITfWVWxnZg8v0IgBf+Rr1rpVcmmWoMleYudAW5NS0sMb1ndrtDJQAvov3fJrg/DmYX
wz2M+InD2gPWYw3cCXjTFP+7DushiYFyan5XP+kt2nGSMcajdQLxJma6YErE56SIKx20iS4n7SHn
bzH1fTYlYXbN3Q46O/UCr9fi4NGBe9USUYiXwtwTUm2kfcGIYJIpPUdU8Eha/S46w0rbpjto4B+m
eUVy2U7CZG2GSrBs71jsTxMlSW9Y3cUzpKlIZsUJF9lDPwblv/5g5gFeFq3nycKg+Zz8kGRm/Xsi
0ufQrozWaktA7lVW45krp+ydgwMQtAYp0iwvvbZcVxSBR84vaAvQYR93/C1LhDA31gE7misxTEq4
xZU5X6Qii/wPaswqG/ycbvMQAeSXz6EBXaq7COQJeLU0mc29EsDrljhhorCd/N4kwsRTTKsF/lSO
IzNG+oVNpQ+NuhL6XOmP/0Oq4cR1omJcOJR5ceJW0S0piv0iW96Vu7GRC/o3Bc1I0A5wepNgHEfd
Agn8mkHI6uAcOIQ1lwXqW7sA5vVBGz3Uh9qpLY6RoH8MzAOu1M7yTGFHFkEzX/R3aLLxM/vRboVd
fA4Jjqin7kdf8uOeV/sGbQy/DqTeOOsEhYNUnkMwtNUV1yQGofnxOQwrvFKPFwWx2jrZBiMW7512
pyuczOU8R73pUtQEftux/2mqum0sC8mopW3ghtZQsfi65AlUwiOc67guZ9O7Fi48zk4EL+3K3uR6
TCcXdUjrcjHo7vWC+z4vNl7xexJbVuL4c4FsgrGvlz/SPfSK9PLoQy+XtJQi8Zl/0EZD5x1Nwmsy
JG9N2VzKrcZWspv/mvgiJDj3h6ZQWssqZmhPz2+uoxxNVCwMHK9NNBmyZSDo5vANSZwe/yC4Yk/J
VBte0X7pZRO4Ad3DVAxacdVYCbKzVYdJF6ZXGE049xXS0UerrscQ+hjEXm3ixDqaBChyB7n/qIEM
Vx9bVS/4m8QxUz5pX4EXOuyjc2gg8aii34rAfk3+/CIEIlyZid/gtCyfn3S57OiZvIs4qfn9bu1R
tzfSfOqw8Q7spcWzEYe1QB2np+B/ZZVSqpvhQXhwTRLWgSkQvmhIoMRN3YriapQzNnTEwgKUAIMO
AXp/zjFrowIEWPZcNdPATcNIxTLknuX1VtHsXWpKSwiWqikMfpSw+GUf/8q2ggygXwN+kaVYNd/g
24DXMga/uZzIAzNLWLiBqk+lMMrHrcbVTDWrxkB/JE0oMA3+rSdUQhsh5/wIEbxoP3YfqUT4M9M9
HaxTfCqumfREeBRgGBY7CzDa9qce+fMAHrfZe5CkIN5KLQ6n/qdGJkH7fI6qMVT4hGFziCBMleOn
/nOMBhn3JYbF0Q64N2U/xGvJfsIeUyvx6v02U3GJu20wp/To9zHWe1Dwp6YMr+2GVN9NRTCSdXfh
UICjuTUeves/dvMm/QyQc8iCP3M9jE5zY3Mla+nHZpHDzIxHLFuexmgVozjG97OHDVb6+ISWmL+I
ISNmWlC9BFl0en26gZM9OWHFDCNKNCg7urw6OBI6yNCDq1hDL0lwb5ln+nvOp36ERx+OWpHElUbH
ODiSyCb2ECpWlwasmgZHgcJWY3p6JmsxFLaOuM9940Gp+ny5zsrFoV+2PpOSGexW1ltOcisZm9PL
m3h+GxdxhgLN4wWjmX2Oo4aOOUS7GJxlGzuSIKn8J67og+pFhGy0m4EZ4lrdWQzDgfLP6rTJRZXe
fJ5lOcn85+1XOkwU777fnA+TOGmbzk0hunJc5TuRnSoqqRZCj0YUvfg5Sn1yllLl95jFoypjhlYW
RunfpML8JDgUwwzjBMQeb9JmFfwDobyMQyUglE2L8iE71rYiW4b4gZ6ZGjSeQ/BrNFXmF4HNRJ+v
v+wPibHK1vfezPNdxmQigjzzp0bYC3CCL/9XVtEMADBOWBAsvYQb8d5mcqsk8aqK9V5AbwOTapLW
dXGf9iDCwcC20gsM8ZfZ5q7wKysLJSXOBbeV9tuyY5M91GErxYtcRIVKFq66Qnbn/J5GgNWoM6h1
tHmQVSlE2IF8wMQ8RehBI0tQWOGy8rcProvnS0VbCb5rsyxzVmPIOpejuqStE2yZwy4aqnSjMG47
sri8SkJQ9ED+W11T8EAC7dye6i98OR2/ZOJgKLJlHxQTXJ4qETUmr2T3uDSMAaCopn+8DM4SXmHg
d8TFapHyI+w29HG6UMFxVJfUpMB/V3TL4O7g2WlQ9CQcUidHlwvYha8Go9QM8IeTQZtHv/vz5cdW
W8h/eQppUxE8yCXTpbVmul6uUuj0HGcjmkllHkB6/Koq2jYQod6KbDoiuDDxVXpjrX+ypdhApq9g
Kot+ao6heak6dsPToN7a3Hja2gtbqXWP9hxi7HSBbVLSr68uKwfF39Vun+WcyGBrv46G4kFMcqoV
cP2ZQwraVaBSI0UTLa+S57gX4EgEqdgokVLJsHh8kjqusIRanzIUWZUSdkfIbuxng9gLD9YVvOy2
3AQChybe30o/lecaYTZetwkjgdPpN2VsCLsYmhHL92851ADUELhwgOGglVGHp9qRalVMmrn5oss0
XGcVhsdvgqUzimdLbDzbs6iAEZV2PRIThYznpVWYDrEGEAvJVTpM7CHxgZjC8+U5+m946+67HZh7
nmpWyeB/1RWDjGdPE418hSYiVSXXq9YVU+el4O4Yco5e7ZUHfZiiTXR9rOrmLKQVyJ4SZs0ZZrDp
RjQRgKK7WCHz4dhPOKykloGKO2IPtSJJmytvBsefP2H064ZsncvRR5rkVsP8buGxK1JU3mJj/NiO
mEs4uzQNOdvrPtPlAeVSMlVOXtNHkZUTwq1RRDqnVQvHds4lcz7sJftur8/FYVd6ymL/DrHZ0GPu
AkQJG4OsKixNgRqH2bVOf43avPwfVTOPnDCaqudQTGGX2cTA7ARIl5s2l8oDSG7DAhj/JQEqF2bL
5u22nZSnr/Sac9RrHtkW/RzwFCh//9YXKNqifxt/ngFNFRlKwWUMebTu6asloCFpruqZIVLQM8ct
r+ZbVRdI8qD6UH8wd+Kh018KKOWyi2CURgCPpQv1CLS1wPp4UbOKWMRY73fCwIFPBEtH8KK+5KBE
VkFqyArLIb5yrRFADPBXOWqs5fY89V7PQ7rF+TOLIgSnW5opFVkJEHjd+z0fiuwlP47fPTznXZV4
aCNeNWtg5y4PW9PlVWQSlEnQ8l9Zz+IJ8f2MO1DRUuqPkqTTbU/F9Es1HRnnG7hmXTiULD4zGdQU
U0XA7J9o/NELAhPqyGXENu6eJviIZsDkUrasmrBATRcmjAFfMgTU1BfY07aZZuwNr4q8YiNus6rL
KO8v2Fztu3J3ZqIrmvhID0u85B64nGoWMOvmjJY0VaREyBLBrWNGweQUl06ealD70irmIjkj9IMk
mH6rVnWdO54Rjy4fzFe4N8jUI0QPKj0wR7QKPrq/YA98fUk5okFeGF+iD4p0k1Op89J22Y5kjJCr
VLX/maQOgfvWUlu2J48TVDeq9USqZ6FkLuoNrfQMaIlz8AqMzu2CtkXtrvcSxOmblYSzuo3yVtmn
WULuOHTLBv9DWNNDFNtqE9J0jkUz1u0odP/wmfaWFGcdOkWFXD0Tl7vC0Mu/B0rtO/6wHfcfYibZ
po4LzErpOz9Blxl7jSaynL41F7HppBQ4d7l/Sh9BKbtHoi7TDFBXxsFU27Vf/VSDcsvWYrbetbPl
C+SEp/Tay5ynicgzm30BhD7DlQewqJgRR3+mlfxNAM4z639nn799rQiZDzKSpd6HawFc/lMTJUmt
2/TRRT9IXDBEFKHSS1Y7gCHrVumYligdAmu7WHkP4MjYQPQNTlFnmdkRUlJjroBxVuUzu7TnVsDI
TC8gD8hmM0hB8+6QSJQ+svA6kyyca3YMUG/oRR6rKQZsU+xDNpOCiPWTrgYvBTVkZ8/+tgGAQ6jE
LdZVp6rewZfkTEcj2BCS5RfGm+881vSCigljnvsZ5dMIe5H6zNA7GgTISKh8StfTxb+aupmQnwsY
qxVk6t6uwlFagaML0QorhQQXOQmE4yJ3E2VPbagx2MBCdfN3ElTkVSsQQT+Sx5h5wvOYG/SdN5tF
eFpHRzai5RWb4ClkzlQnKoYZ8T+iQ/6CVAyAVaiYocmpmSOdME//d6sYmGwuuMWLZVR14aRq+WPz
RTD1SuH4zcL+Xew/aYSLTy7joYDD2i/rtvBYb430PkYWOfNxyNZCCiMxBalsLfAU0iiw8paBYPAP
O89DN+PEibGJCIU19c28QSQQ+u4hCb7jWPzAOSW/iPFWLB9FLJ1HoZdCNvcSONdSahhTHKYnYGZd
1ShDIEhla+x7anja77QcN8Pt+J4ydSMtOyNrH9YZ92AXtuqtCA0IWLuNzfrRw5Iy5t8b/6ACp7AV
VmjcNtEtj4lQtk98mwiHyfecYpdB5os5gBugXokPhJF8SZEIbH/1BZyR86bg/Mx9PxnIew3OW3iE
i3k+EEXfIUfjWx6CtLPgT9qa0l6y73SAsmSFuKxpVBvP6y01V+P37nBxBDpKhDjlAah4sj/53xH+
P1bTWfzw3Z0ULZ5p9w09NBV0xNsckbSc4bb+V/lS5lwOR3oQPrCF6OJyhU2jRL3cN2vqi3FcofUa
2RR9URUprmdfXC40OfV1ExCQErVk7h6l9YM7ME2LRPtYEF588h0lBjdv/HKUmEh5JVp/IwH4FPpb
eQwpMYaAraF9kHt/FHhO7OgFi33hT5fPhcZ0YgAt8x/aF3zmwpg/sUpq6cd+7OfkhemMkRu49xTx
GFJ6c475UES3xnU3r1oVb2JFkisjIZVf032j6tqBoW1yLuJ9duNpN/qzdOQbEVgZXr1X8aq1L0Dt
qKX4Y6gDti0QDYABb4qYjlIvZSNfmCf9LFVyghKpBnXisBoqxKkSW1QwNlkP3oyYGZGs5cTGQIQL
oNruBk3U6CySezzLb3LaIUSwq5gZ1bsPulG7oVdAbnnrEQMJeD30M8ON64xfdPCNuOHPFZhC2wsx
hjjkYwko3x9boSr70K/tQFWFMgVF16Ubizl6lWTM58lh9NbEvIqEVWgcPMl913qWK6rAk2mIvutO
BI6tjCgX0xgWR3Nhmj7f0LWWxJV6y473KOUBMRqJhAtC9bY8xYr42qz2+ZxbPEhPMv+ElDS2uUSl
5kvXEdTT0unCyeQkhCtsv0ZFKKb4ol6/9Kxy399mUu96J7PLl3EVxYLgE3V9uz3MJklZ3VZeXH53
BfQM9tIjmstcLqSYmWwBpgqxx/wo63wwvchyfKlyJ4TaB6wLi8fsPgszU82YH52AnOFzV9MMpTSi
Q6fOG/Ork1laUBpitq8kq3wen6V8VXp6QMzFSNOwPTx3TgsxBipCXYGo2ss0rvnyo3eL2IPef08K
wUVp2IoSEakrZsY5mPOvD5w9qe8dxAqZAMz1LECnUhjTqSTk0JGTF8RGuPF+4gd4cO+ku7uc5LRy
XkPekpA7zJkb08BKkwUQpsm1kzry1OxqD8ygUV8pBmBrAEmC5NQoXrOmHy1F/xpvGjHdp/SgwChj
Gt2gRuS+Cd06pP6YQrNfVdOXIwpnAa1KWZwDsjyrRjujsxAKB6I+yq2pOm0TG2HAv/ZQxkPJF203
pQJzujfayMEpH4ko7B+ryXSLTRzeN68Q2gUowbIt+aOw0rVYP7Qdc4JsjmgEa4k75himg+YbA/6n
MdN5tx2dmmL9acJ2DaTGLvpm4I95STZfr8u8TCTumUBPVLuJS583io0J2aIj98u4aAfI7vXskL/Y
5eUlVPD/+hH6vc/zSI6qI0RitkILSCIAEwQ7POOEDa0eCAASOIgdLlsl6KHujL3X9FZboWa+LYmH
1UcduotxGLGiazYlhTdvnLTRy4O/fIxMZT3nROViJZHlIjIuMZfipPJFLDlup0YmGpHQj7+jDV+5
2y0wA6vOXPniQ+4trzrHcyHLsIfaOERK93/QqdmBiqxYYZ/83QottR8qmu5eRHMp4DI6/V4w8TYm
6+j6RdXSAihuLW3AYjm5pCWxGiN6QxZiStOFORcRaYE0Cv8GDR6umFk5mkpWPcDX/uolQtgNBoB6
NwdiVZzZebLIp0hhDZBs08EezQCIsGI/sHgYEMpmju0RDiWf0u75izc5u9nybs958prFJe362LfU
xQthjFlofOj/WOWUkWa+tmYKQiy4Ap3DfZ6Fh6CvMkpdWZXvSxMKEuoaIuDzkZhEN9mbqCF/D6mU
cEXX5mACSGe8eacAfUq3VVOnwt0hAxEA7Q7GbuCh8Hk0/BWQKMWQ7N1Y0pbyJIQmOfCqWgVkYORH
Ft9twxZZK3bcH0aPNoJwXDTNVr1GI10GHw4n33GfQYkcQ1xR2nsXdMO0nAmFN97YN8aIwQPWuvIe
4i3b1Pv6/3/S3/i/hicMlzEN0m+DMqv6T7g3Wcq8Fx3NV+b4asoFXMabpygwehg1nW0klCl8s2iW
tUechdScSStNZT9pV7ZtKJlz/+TQQ0MsOkXGUvhLNV6SB4NZgW5rfLgOPPSKjkcnt9katcG5xyVr
HaKNYynxCUUynguQdZ/ae29klh5fy4OY+NAFDW3TQtKL3/bPoBeVCwwBHFu03CRNlHYLeRdcORBc
uQ//p1L3P0d87sMhVi7xh0uRhCyf6PM/9mZzAuPYLu+Ffe3hlEoDxVdNN8qIJof7LYa6Ij+34QMK
GG5F//F0zBPO7sQ9Kawv2X1e2K1txAd9X29pTPFhY6Q52bo00zQHn5xI14b8uNikwl+2aGh5n9PU
5bzZU8kDbxTr9yQN4VA5GUNOY4V2ku9J8ylQ8d3S12nR4zaKAJx6VmLfFavaSL9/LnFrZrZ2/CFV
4WR7WoGxc7VBdLimycujVbqYOXND4uJzAVuuWRjqr2SxdD7PUQvN6p5ETasOP2IGoBMsY6RGHy1m
4Mcm+Iler/wmwA18abWpFbwNeYsqef2sFW20Ru7PZc9p36k4r+yh0OdMRBPhpBNekMMmoCFE80Ah
yjt/PGvdvCANnANsb1FVDIXako/qAbpMnXlBLSMzSvsbqn4dCY6eoHi52RxhSotm7BMeCUgSn8Aj
hs5i68QouZJNDwiSr6tQL/Rg0xnRmeUEto01/CLIaPn0frIcjgsLdTjCtDmeaZA0jpFLMoXSc6gQ
3V/JBiNkcbg4zYI7cBfsUvhAg8UEk7o4+/zlGXpFxBScEW9k+bLadeJRXTuIwMrh/TvEWrx9j8yf
M1WqED4wNJXTROh5CzMnRAJr1YNMnbGOPGrlU6Kj9p/NCSw8UHRZMr+ryxbE3Oet9ZcOC4tfYHi8
S/AegItA/bQP1EC8wlOa4XREYcvimJrGJobvLhBOF4y32ynISsy1pipT+TszI+K37ubN94pbOprk
oUaeAmvPNK7EfHDYp0dXkzeniXPvw4naqM2dgkrLOLPh1MFcxF7zFhu3/ERk8UWWRGsxjqWrzS4w
VLasX6EtIYe0pJvszsgK5QlQiqwWpQzq+ySrFlci2jvdLQBbYR3p5Z8J/p9aX/2lHD8X3p3TSB0H
6C/ggRE0TdrYIxIMxVIM2KAU3Bp7fkD74W/Riw94/sIpuUc4ckWsASPvNY0b5awqyIQs24zAvVuj
oW0BzNJPO4iQLsQsUtG5ecaBL1XAn9rX5HgLQ8VX2U797ySdHgduY7N5D9lx8ge07VKpx0Xn4UdW
hUz20v5Pe9ayg0d463owALTgXX81XVY6v2rAcn3CRZbkO/Dp2mxgVbhWLrbrvW8Idsf0neIC4I12
qGF/GRh9hje9Svrn1Oeg8T8BBUAJTtQ2Br2K+QYqZ1TNtq14bqy8dOPt55Ok6KGZs87G4Hx7FCvy
vz+ISkWti9gPYbnn1mEZP1kFOjD0F/jZVwHE9fTEApMzyBy++aZlSG+ifJ8jdbvyw1MtmTwTZY+2
dehV1HTkq6Rv4as4qe24tGph9oL1+umaV8an7LR5U1jStseThcMFvFo2KxB0EePr+oPkw6EOohG4
76tnO26Tc9AN64xZIaGWBqgXTmGJ6T6TfYP1P7zUcWFuyyOpTCaRBKKu16gx2Vnd0omC9XcBzYmb
ReB7nX00hNuZZMr2d18TAi8oYyM7IaloFLigjgUyC5WM8mHhytVsnLeXP5OgC1nC1Dvn8wOn7naY
0tbr7AkI/EYISml7qVfr4g5pSkt0To+yBHGK0TbAOOE2PrR5/9RD2PFe7XnYnkTMoI36Kn9b7wbM
I2pJOAzxnbnZ1WP2HQudrVpcVW/yXjP5WTeId9rW7CyJsT79rNYlbKoUjXQMHe8Dbo4wUxK5Na2T
6lxtrVenVKcpIDy2Qi+pAGyaa7wxWOJhbFDqwRhzK7iawlmMbu8eekqAJWkbKaEme6yUooCusY/q
H2sQ/UiiC3RWouVVtFf24jqjkIiPmBT/h810QhgH8v+OiMLIUpfEi2eEjY4rDffrmcPVoYgddkXJ
UtYFnEmIcx/g0RJp0HZeNkkhGWCd7m7CZzQJEt1CFEk74rxKWxLCsYMCo1mTbUocY08aJZudgG9h
ARnndKsXBi7YC6EnSZPrg91fWK6ZcuoUEosl6iCAnGUAbJWBjT+NikiiAisDNLdHtRT+WsZnNO07
12OaI1xodhziVa0d3lihlHxc+g9SnVIDGvxX47u6KHamJI8ZVLZfqUzjnkg0mJLkH/6dR84gGbus
3e4Igy7ltpn+EsDeWQAUBcdF2XS4zq0slriVl8w3vws5Uem86PaElkAgQ6WNfEIZo4KW1iSFIDC0
Qul9qTYfhAvs/gEvDW278Qu3vjJMygnH9xh5yzcNWW95AmDBLB7zZw6WrZEbyeRkL9p5GhKdYd0A
K+d8zfoZ9rcOIuvXinxW0M+eFSKLv9iVto6m0Junt+bkXJ/XX0KXoKJOyA9hv1d1c1ke5esZmZSy
a5RspJdt10YRuIVGUgyu2zrZQhorRTAV/a88x3eG9kaT/cntgHtWT2h+fqFl/j0fdUkPHSw8/4W+
/I/bfGCE34d7GMtiqZnEg2RvGdqjq5fDUalz0XVdOCN9t2RiiNaRpGch4cKcwOTQcGT3JihIhG+t
TWh/rRNdw4jHkSeMEAT9tz6DUPE9IQnkG62KAY8Dh9UdqSPvQLhkFYPw5ENkuKq6JjGmtBIRMw2x
/r7CfrScNNrHjg9Z3ZKfH89jFkXvqEFZTeDpeuhLj/8YXq1cfgcKhszr5bQTjjVekv51lngEU81u
l/6BMwsgQJcLR5cKSpzGT8dpoNxpd211RL4s7ngvoLM8SrprRdym42jIO1aKRfy5QeL1hAs03VNn
BZYQge+zvAgx1ojMdGKZUhTm9DySuGYSVBswplrImw4i47DQEOGU1Pr2JAyQjYZb8h3jXje0tqft
QTEHSacmbCwPGOMf12iyeplT5beeQ1N+Yvr7o31Uim6KZ/9XKqfluVy2AzzxNYL60c5g8TnxGQUG
uOHyCcNOZ/UAQHcQD8a23Ko0pKzjzRXWR6pRsSht35L/Bg2WES+RNVvIssWm+FqbMjZQURz9iHSY
82jtAIfhSEMqbKSxARnft0wWHVEZvNJK13n8konpXAdXtcekljoicCN8jZ4vjg6n23RJZeag67X5
oCeAtoJfduC4AMx5IVp7lHUxN3Ble0UyBIMFt02nfFDQ03asHbxgNhkrw+u28We00dK+LQYUAXJe
zCdfR0wAdlEf0bkh0CKzJOtlX/5NqjnlZNgwB6FdZQwE26HvQEAAUCgxzPegqFsGpd9CLO9AVkNp
6Hthm0XCZ2lLiD9RNewEFONb1pLQySpvkNVzW+5S9t5wBwracvj8aZGpWRaa94TlxNuLSlmiHJwK
vM+yslPTHdq9iE93rGd77iDkOMLM8FjT0MIM2cVhEJON1W/NswuMoqGLlPFHUf5GcOW0Ltnr58Fg
RAWF2vQMfI0fjSKI9qB1I+yAuMNLQJ6Mu4JJjrKHm8XypUse7A57/UlXX3kYubjWTi7rE6YvfMAd
dIQT8lzbg1oHT60LCNG9ge0Y1Y4YOsBBjgh/xEB8hGThfBI1VpYYFBF0b1HuiY0VS8ZCzT4Ff5RU
Nfmc7VyUBV3kcUn5g1DMBdYbV6VlO50FfP54lxjFMDZdrgiR+BhmZSe03lGM3QuvX5RiBHECTicf
kXoapPVhqO6qHejpuWGxXJDIGlYOaYAbmMMIgwlVpZi81P4YLEGw9qxHtpp+wLLHNCz5AgImPyAC
eviYTgEQ7mXudNi3Z85vH5MbduKQpHtV/V9R2w1vqVQp0YYAYrbDa30wez0AakF5ys4MSzhlyX93
861Xf/NW42J9L6BgNCsIs5RPOtnyIaH5Y8faulAzXUhjAOeRr57rF1Y5N7QNeUUCTrCxlllIRkTA
14qajb26/jLBcYQt2+RD2im2r7JRN+kKJJtXq3j0m+8oInpU9FNWqm7v6ghVIfED4n+QI/32is3G
FV86Br4JenFhzkVglr3SSvW/ej9K5kZkTGSgQ9zOFem9X6sMlXuIFdq11vE4XRO6GNACiGZiqwvU
0zWBjGzwPJgQ5hR+o8vnSULsxS2y+7uAPjEL5vGbjACHkZ/aysw3P2B/5XwbN8ssbgX0CHwF7Nds
alEdFw8LCu1fX4EvZUVqgyk7EvxIRe77JqHCDuwUTaKNURILzqQteRy/VSNzEwsKBWJ6W0laLVz6
0qblLZ39FCmFagfl/8T26cS8P2/Ucvy01lAweh61Y1TonKnxHL7I0nFC/7zDB5sNIV2hGyMAKbw/
JMFSFaWIdackd7h0VXVrf2O8cvu9+sXiHWcerdx+tZVc2O58j8Knb0kYVy06/Y0YHddxr7T7uiC9
3h8yagsf194MEUsT2tTX+8s1MlEaKO+uQd/O7jeLW7G1nUV84fRKeWlLbwWsK8R9DKkeBEJ/G1en
P5bhDbHtM/QEpjn+F1MBdvzYFcDUlZDz5o4MHVx0e17i/+W0Wbxs8t6OkwFXEiPuR1UsDn1WugA8
K9Y9ZITjmjrqNeCxm2WleQITdbp/l2pDHFfwBnbBqloid79xrm5C5WPaIeuSGCloFm8XamTynROD
S2X0zGpjIq0J/euKH4qOsPBlcJBBbfswcREzFlSf7nfFX+4/ZsvmFOLQqbNdH/MEI1xfeSEkvuZY
mUM8lpreUIOJI6x/Mx1gdXkKbR/bsINIxY2R6PhY588FuP99Fx5Ea2rYCFdTLbUvqrx72XSdtG5A
vUROF5btOah7FVZ16MR7TqRxHj6/TM6LgCHXguJezPWIClW8TWEg+1uczXSbOOBh3eyp4nxgnGdp
Z6Xzmha+4XGonmQo7U1Iv/SRRo8bXJd2oGuid3cOAhMckX3akkbUG8z/UEanyvN7aweuN990HQyc
1MMHyRdElCE4i9TstTwSQmxr+TvOpagnRyFrI3SnwabiZbOvVClFEn+9hZbptd4rzPN4XVwfWR7r
mRUZtGmHyNbpOByQ0aBzUZKr9qxW9x6B6E2pwzVuE+o/1JJHfgLxozgmnqPYYxcQdVciji2G5o0Q
AYWXbmsKBIb5NHviC/QvzzeaqI9aHvr29bIISaLpojgwVbsjTxlqRJkWiJmwMKCrHLVAtU6byqeG
7LMS9hv48fv4SSoqs9GJBYPXC+PRlFScytUpMAlBjIAnNeecaL+Kr89yXPeS8FMP7wxVXFKjlfpX
Xow1Ed0H8wvaVnwZJZzq2DEsuPvocSKSaxq7PP+V5N7oZEPu2qSa2kJSnC70vQ3HzIEfWMxJRteJ
c2l99zt9mQQ3/+zk0cNwHPq0HdAnYZBJ8Q1+gwjX9lx2MQVVQf6OkXGlLXTVUb0iyY5fL4vIC9Pz
H8ao2D3CN0cALlK56ask6sMtHYdeaZJ5Tk+VEGV7TsPW85iNiH08XQCJ6Cm01Gma3LIuuiW3Q3KG
HS4B+ll6hVaITpmISJdQEOKclg59JXBQ4vN7FtZwE1rLoIJbgnnrKUtjhHnVY8rpapZtIBdQ55np
yq7XMot7gLYUeUeUEFQJdtBhxPIsi5sXbYWDhe4Ti+J6cixwLQtCbnuQ+ChibeLwka+n5SuiWvji
qUl3faWVzoPR9yZvx7SHZnfg9o7SOploOnCBLLbV5rt3J6saCkMyO1dG8EbHVJyPaiPw2OV7sTXJ
7rg/jgZJaxsQAOaFLO2dEaWx7g783geZmJeXJoGrvJmWQLxrqVszFLlW1fEqG5ELzFB6wBBY0Ien
IuGYZZAbtBwd3z1zL6Xo/5r7fixTyCVYdH1kzVs7vJggXsITD3T42wu80XSvj2Cjiu0SBLmUBXTr
oI9x2kumEEXAUgj238uEBZ55tOwk21vLK5Ja96Us83Z8DplLBcdbq+A2Mzp5naWVsrc9WquApj2x
dF4mlVG3c+TJYPxmx4G6lEj7qjcL+7/ZLHfcqFKZUqO+S0QOcHfU7IAcgeay2kAcSvI8mfJsYqd5
N3HdXaCARx+MPfO2mXe+nP2RRgWeaLW0MJvFYvpwSwx5ZPBsAvy/HybbdsOPhYjD6YJR/8TP43Kt
pTyEg57sdHuh/4gViBIpb7tubGoBEgH5caPm8r2BaGws0eBne6NaPO0lhUyaAXbVCgdM2kKIHsDc
pjAL8QLgjZAlD7wO/JHedvnUKtnkWWvBxnW3fERo91sHFT/VqJUzdWOWAioiPvSu5FzKwi6ZCDA+
x5G97RqmhAuSgKT25QUXGf4ZqnWOsFmH3fj9FS+K0/WIDx6VhJWcHTquu38D62l8TCb2ZlS+RM4c
iLd17Gz6lwK8LCwTpHt621bQ8byO+w1/+OPqAnRsHLUfJ4VVEA10K0hgS+TsZcvowp2OQdKJjGlu
zqrQIStmyLrPEmYQesuCmMy5kzxdpT/E5a5zP3WtZxdDTj1IenoPwy29i9lKdT4n8jC+oX+YtSa5
0TRW3gCFZ8LRZcHlbP+4DGgg1R+PMNwdzM1Br4VVrUgDc64rBEgKxV65LXxXQDYguBGoveJs2m7f
Md5q0L05X+ONpGCcH1aVBuZ6OCLiIXzo2bg/qmEHipimPsInrpXdW8yTsXaI2od0sxmS6JcYi6O7
59OSrchBvPsqSSntiuOCRy1H/phn6gtchyT+aVxDhZO1EAHdtd/J7yLTHC788BCu97h1c9owOh9B
DK3ujmmwchWTq4K6LUVu6rhoiSYL7pJmNCYcxr7dABRwN30qHdd+l1hQQ5CPUtmxkZ1SppndT0Wy
VG7V+Vxn9FQrQUmQMEd5NYxg9/yaMcrfHbhHR7MKZaGjeWbo7q8RxcSQYtG73No+oD4+KrzVbce9
kh/JVSK/ztSJPvVL+jKDUCDrkV30XHuFhrtE59FQviob8zVA3aRMpb7gNnxAqmiieDRk6SW2fET4
9Km7AG8+Clpr9lPqEdSsEJukQqFnx1LmqPa+A7B1r9/HQAw3j//lvr1P4u+CS6VoLlTl7Hi/wbiy
nl+CyR+EjuIZmG+VvTtACPixjSVZC5MQMpcER9zu9y+pRbrZ8+DCiHh1h+gzQeYXXwYcS92N52o/
Tf37SN9HL1dHaQYbbGGlb42lGHUu66cJ/Vz3p0S6QM9Q1kXUFyPWMtzAlj8D90PwTthkNdwmk7xP
+P417cGot5FN2uZyM78utioQIR2Mc4TziRb3pNxtDBsvMH/SgULsYV4yFkOi0EmvrZenrMl9rw2b
gyydcHO5OhJT4YE0t55/i/ecxa1Bfs5xBaw75wXUYYOz7wmcFEnjOa3j55a3RGCohxgLG+RHDO3h
hN2cJcuWi5uv/Qjw8yFU+E5NTWvO1Ue3sulH5JKAKZwpEKm2muji/uh02rzWfqEFtPFhxlWEim0y
bjOGzI1FuzpeAlSZw5yAQqbWv+aErgFa65rnLz6lgtp8nFGVzUiBXpKb180BWwfXV6k9tl88H25M
r1w8hk0cybnIGdqpex04MQ0QqNvLEqbrFwEldUreQXyAjE5V2Bbysbh+NrWU4XXpZ2IztMe8KzCb
WfEHnFSIF0wHJ3FDad82g8IBj3Xtl1rL3/7KWFr1NCrcDJG8IcfiI1Pf5M7CzMyHOWPH0xpAsqeY
fJiMIdK7Vr6RQLcyqz/qSq2cH5fwyj4t5UKyQh7r8YkbNdo8tYYQjfStFpGoKDS1Kmlg4UlHlBsM
zYUr7EEUg6a3Vqtq/D8sKOdZcV6h4iJ86BXNGvgef15MgDEH3vKGEHOOcIWkb806T9ezzyF1AhsS
cyH3VWTZRhL73tFlFwCaARJn+gHy0EH0jX7T+1QfhBffAxswXTCd6S5tffNmSLAFiaEoHy5nfioJ
Oa712C6vmYuG3AoQCD7PPcVNeeqEglPIrvmGK8nE9ncmNYi+BG0Wq7xnfyfKtSpT5Ab18ngZ6ilc
EYohlgUCRYoOTzzNBy5qZtEJQrE7Jep6WvsTSJ+2tVToX3qNBbMEqz11Tl7myRBcTLQHc97xbRxH
gZ3ETwZLtylSTaZqd0A3436NmQ/yx/6ggdIXN5q15fyd515+B36iYLs2exrMWeBQdtNyFsutfCgK
NMY+VSiz1aC/ioNT+a90Xz2ZboMcla76xjFTLqeAii3frHFokP2m2okaDp/bNBP7VuBp/WIKJDda
Vl/lhYEjx+o4ajPKPNZ9QW/UmImTOhPb/jd8jV1QXRyaH26fdwWER3k+PXQn8Z+aNL3AIdHJIFRk
5VeelfU9wjevpvg0vGZHYfWgGYMwOEK8A5FfefxBB8IlYE7CjrMCmHh9HkJ7nYMO6HeSoejA7RIC
gzigyzadwMWUP/6mfZP6RNUatkU4SoQg0K5iZn/KPjS8Jv0aWlmvya2kCVGjGgDsU3uv+CQHaPUF
+0uP4c63uiBDHl3e+vfL1wPZVqgGz2+EQzXIaaWgI5B7Y+SJdkz0DRx545bBl1Frsoxpek+begub
lDWoZ4to3DMu9cs+ChRMSU3REwXa8xw1NtGBVYfUGZA2nQ7/Vn3xAlOdlzph453FY7gkfxKVtTX5
fOLbPGIKgUjMUbjo/1+/vWbjLeLjNMfQSI3/VSnVi0m7q8yez0ytrI7nW3ta1g5OnjZc2X67iBjW
eA9TGqu7FvQ0ha/9dtT30zBeXbGNxRki3HJk1ctR369STKVLRTHSpW5ovM6PfvqCHHRsSdNfXDnl
iIKH1ucxSeyb//5RRgVyG5suk26cdulxQSbESYcy//y9S26N8zxlWpUD97orRxkGMdr4piob/2Hv
W6dxZW3bPVOvknQHNQOfCvnHRLMGjurrgMmzSb3uqe8Uc8et5vHrLanLm5hyfgFrwCR9pGaBUrt5
GedqElgvd33oJECZJb7vF3sIrTfuJLyH8NRiEtUdEZzcBXKGJN0uNhxxCuUZFgnrjwEFZ2qDN5OW
yZud3vauv1PK4WQ9gsvF6f+8qXhRJwm3zABOklww+d+qLTOWraHe0C1Z0ZKa9aGhyobqSbgIqfGd
bBTv67jb55t6uZ/Dj3Iz+N1XB6n9gRoEMO1NqMXoGI4mzPQTtKQLJHwA8//xN8lZ9wtOSQ0IIcvw
7AN4Vsgcnj7AYNbnNFEi094/9cSw74jHZTK4wV0Za722WNT0Q1maeCFTAwIaX9hWDqcfVNmAdwLO
In4boEpgsr+cHTMvO6n2nzaVKxDRtiMrW6Cyq2EW5Zr+rKdIK+b7w2B07Cu+h4aipDC+7+Sc/Kk9
yCpx9ZtQ5137syjyiLvR7K4LMN3OHFIqGY1r6Y/WOAAvS++fzor7DrK9vgzmeYvNxCvasVxH+51h
EDw5+DDvy386besMnLVKekJH13IFa/RymDQm9I0ESYUc+t6Y1HZ7UyjmWMqSHFfWVH1oPNFekM8V
DT7d6BosRtblv9xe5WkI+gJWSp2pL2AQ0Ro6ZSx7nn3l2P+YYmDxDtgtqclPIY/vLRerWIW+OCG/
OxaHf8WuHsQxtSoYlPJmOEQaFes+fu0CijY9z/+UH8W6GruYvwnARalOb5hXhVXdhL5xciNTBLlt
1Mykix3qcuTiLUeKmjLwEKTgtym/67g7htcDbtbUQPdKqWqV/48YVhuiWdZj0NNnEIBrV8Bf0whs
D8AtzFUS4nYdP/rgp7GSBSOrGJwdLbtc7FR7SUGj0TIljbGNsHBKkEP5XJswXu0Dd1dSCBIt4XON
4IYSbDm4GI1EJf+qnfjQTmVe89i3hEL4dldXFUSdGoW0fzTU4jhVsFxgXgv2UW+y4IbLC+uf6PYp
ca8r5ffXX5owUDu+9SmTCgAOK0Fm5AT0a5TOgE1e/tBSv+TWqiZ0Vn03c5QVuFelzP6GIXxTzAbW
GZZlWatKQR+pV5MbrSUNXBDomk0wiZ96K1nRvZPL7hB2smFe51JaaY8GaqZ5ckIrZiorfilCV/Wb
gkmWimg0ip9iTqJBSo+/5TASj1xITzmwJ6fQgYm+bNPjHB1EUT8mI59NvfdcSrLl6gAiR+rTd72n
lA9XzZ49Pdf7wSjIhsZTT8/8TFXo+A0cCyS/NDh3ols6cLN0tLV+Nx5rrrfo/etc2P9lr2+4Lbdk
FGd6LTEqTizIfvASr4P2UJ/3BYXKanasJ+Y1S+0+nz3wklztHDNS3MKfe3dN3ckuyAkq/3TkrsVr
eK9GKCt/ZOh3SYFsszwaePVg54p8U8O3recZJ2kO9mfzRcWOL1f5AtPI7u1FCUQmaxA7seJ33ZtN
1iiPr2pyd8uawflfmvEbyq9sDyVZpZJgfXE09ui+qTwyJ3bCXkSqJ0kWNbyXXvqMvbOfQibXXgDr
5O1qZSCzl7KHqq6MULPb/x7qy/qDfrjdZO3K5V+ljdmnx6jtBIAhKYcjyD6W+NONoGhP7luyi277
lhgEgcMY09oIOBdZFKlr9aYyjdkS7PIhg6lgFE+E1GmzulPzcwKZlpQbL9mipPHnNn/3ErZPlMDK
2qHZJtVlAXl+Uk5BZOOmxHX4byFoPsmYE8/03QARKGy1+DsDtGIf43DCwhFDpYefclKgifR2NHgO
aDJfx+YTFMfgm+jrbpoYgIx0/+Szmh1b8OIPWaw+peiYnXRCi2/4XXq1cdcEkikMFrwoJLLdP2Ih
mbf/du5OBAGfQVWYsh5rB75U0Lubra66dCmqOfF223ptpSkX842ErbuVgu2KVyTR2BkiNyAlTrtR
/h7h22p1us5OR2fzLd0mj134ZUJPtyuBNJSL+RcUjiEDPGg+LzjPRtnIP6R9sGXLsn3U2yKODttZ
dP8VdsyUS/MlqpCv2u5sTCSRcH8O8vZqn6w47tmUkMYoHP+8TnL8AXpPPMmwC2uc0fzmVjNODk1g
NufP3N0Ode5X8c9yj8nRaKamMsgccoM//cnF1Hp5WkDd79Ezl1u6qubtbV02DokAXR8UkLn+rzYO
jqV4Qr3ZhC2Wgp2kFm5stEVXb19pm7HzNqR02OIupnDrmxk6pCrsj/AWk/5qeR1aS60JbyERRpQJ
Q6Uut/KkmmKHvCbfLy5oViJLQm+SgusjFfsFJ3vGIjQicn77S6bZxEcl5CazrArjHBJA47+qmvQN
1jTJs8lMBPex8FKW0WkKcPVUDB7VU21xVVCk2wtdchOvwtXwADgeu4HP+Zj4upeXbrJliyElg3h8
w0JTjemQwKbZrQenD4I3SY/8+lIgviHGSh4j9/jPftW5D0E6OHBjXVD/MTgkw6nTIZXMo5RBvGOh
H7uAgHKkHN/PtVqSE13bbKsgnm6UFddRRA46UG9omjuYyyjC2CrKN3LbFA9tb74rSMn3vlTMAHy/
QMmUJk35i1qgUzFvHe1Q8InsOyQJ02skJIGBRoOudDqJ2sSXYKISv3n/v2+3oeRcrDqHWj8+2PWe
0A71Wyo8s8dUGxDRT3l0LQVqrpqNNO16zosn/bl9k9xht5Al+RLm1fqMN1nTDOrpxP9xJMrPYjLS
7vcoMkuSXirHuALvE7CG7igVJExt2bwkH/n/7Xm5ljbjkgr4hLYzvuIhqCf7ZY9XoQre5zTWAsMu
q0hp2NTHg7z9w1jyHF6i8Caz2yinlNgNfmd47dVcgTP6DyyG4lapl6e/qAwF1R3ZqiiOlHGMVlSQ
tSI5ZhA6yFQ1shn7ctrYfAUWlz2cHfIvNw8j0xN/lyUYRz1vN8v01sSIaWdY9X1pvA1ba+aYESzk
e6cE1NJXpxasYZzfg6q2vbTIYHC3o8ZevG0tdmrYx2k+gJKkKZBIBZk5x1Q1kp63IpMR1NkOJCHV
7uOyiSX85quGkyzSIBPPKUdpXOWsUOiDevahoB05muSH8GBorIe9JhotYPVz65o0iTGoWcICG55n
XdSIahH1NV9rJmlFr6tVpGvzVtq6e+xAnM/KKpO0uj+8YaIWrrCuHZAW+RwH4fSg5Hg2q0X03uNQ
OfWnLQ7s4lD2dSsMfn3mcdFPnU3eUgZ2ACHxPcUilvPdsG8DxY0GkXlXPL8aI6rwPE8AxL/ySEDy
QXJhlpYb3FohVRCg506OcKrnUAs3UjDGDFnNTpUXFUVhNt/x0vkOExBe/NPbMjeni6zfPxtxF/0V
aBv1wcO1VWL3eofFWbjB7DHZ+6IuP6R5LLY80cFRz3M8zd4zMOH8lJUq/syIlNF4JpC5FCBw2OkM
S2YORsweFESQFAJMdoxfqIjuOOIc7oxU2kGxzR0KS4Y9aXNymSNGV16Enaj5M1MHJXLdndVxiJVM
XNUOeOhsftPc4reqzrQTX/7Z9zwmmeTSzDkqohxnboY2cNq+vHB0CA1+M/J6i/Phu+B43430MZq6
Hsauow4pyCFQd+P2qfMO5+C95KL3fuPHH6vHgNMVhIt2gV0VQxHGsoxsn+0EDjst527+hAT7uO2U
EpXcWiwRDPEvqeq1MdDSaAKc3GJhHvKGJ3E+ekbqikECcvUs7+Jdq4/JJkDhzgPa+hnUB5n1UPb+
xX3JIvoFHFqLIbjB5E6ht9/j7XDK71KD+0iwBVg1vLnaAlirRJ9QFyjG7q4vCYSecmKYh7UFH+vj
ueP2ESqFEHmmaQswRhc+FaBnZpA4gPPPKU8iiQqgAsyrii2ux8SBO6zqMpS6V/QXqmWFl2bLGLDl
KQfrYv76ykUUbo3NFkJYWCKlwkrMxSbQZlTJ/jR0y8a4tqV32DYmSgJr9G1Hdv8AfRpq6xvyLBcH
dWZP03RTZ3e8O17UZQxLZsh12iYxvACPh+6hM8JkSUdGzyCSk3Ohc6WCTXdjOGZEPiSbPNbhKGpz
5Em6oIZbZbwKemiH/oPpr6BVjsbxrjPnkCJNAVE3F87qYEkdwcSmE5A1BDV2uChZkjOC7UurExxx
pbeyfHptlEP2keDy/PtG7s1W473MPT7lMa7pk3UWZW5AewHOZk4BATOivEuU0F8Yj0YZbgssuNFk
lUSkmZdL/NBRAjaqedOWbvaGdC30r3/5VHoL/08o1nPGqw0Rl9HbKpyuyHK1LeaQxyVeLNaiWOuW
CWagPWaLtuU2HTqlnoUtRxFkjTEs2HE6kQJBKyvEheqLJq9hFaiLpbIlTfK37SGKi5EBMXbIgXNW
eytJBY7gBlsMJ3qblH0GPLggAkSPsnnFeRyjKykVPYOYYzi6uwSbubVReXXxsgFsZCTnZqy7rJz8
blykfeV9IVMNpyroxBnhPMR18aEWD5qgrLDXx9cqmI/FArhJvQjN7RHtx+fXzKSXm0piye73n1Jl
ey5JOysSF72Nv6QWy6uldxDjEDUehtxiC8LSZDMbqgHAOT7gQApdoNoekJWSip6CpB3jru7zYBct
5hytmH4AkNqJV06t9qE1zmwF8o3V96ashB+SflQRSoS+s0pep/1QVFk1PtjzuGaeC7iRjZgBmea1
j6YYldb6H7gZpbXa664bbDNK5Rnqhiz3MeKxj8I//ZD4KXmKE4wE0I/xFpN2JgQ9Z7i/xQTO7Sgo
htMqDNYDt/RUIxA/MdkJrDQLR68h85u1w4Gl3CVJY13LHX+leL/H7GNculgIZjM4rNVszI42X4KT
PaOR0VzFgDalhPGKk0bDCKrm4yVEFkmsYlCBIukCnY60QcUz8cfLif5gZGL4HduhzabSCNVZzZed
SPO3lAI8q8AGmhfS6p2qgDBgm+xBPCueT+llfCDoD5KWo+xQ+2zUpgbIdApgT2tEV7EoJ2dOMMX6
AQqyZfHgxXLwHFehNKaKcXlq6Kp3j2/0YjCZ2D59ZFbCyNE0Eap/rWmMMtQ2Dt9T4hRk3EHv4XKF
ruptlVqBZtXWrQgFza1dIqUdRVg68LKQCSESYLzFO6hOjjB/7BW6968TK1MyZ/4UpPaLBkIZF5qp
vlkUdiokDGGBay3W92BNXXIOpFX9YLsdMlsOGKf4YyU661fi0pHW10u80wR0MqHTQ05ETgJQ7+dh
FwiWZ2uRSXM9vZBZAQ+J8njSSgKHfJ4I7PjfgtkFvTYVNKBBbsLbN3gan5H4rsIs3CvQNxdYO0AS
NqXOyVfFwGUmKH5GkB5QePhbKVWkZrrPFBu0plC9cwPOBTfPtTvIQMAzh6Hh4JR5geEAxcdXz3bj
TPG+ddueGAa7uAnghjjA/Wu18rAKnnr1qCPbt4ZaewetowyzGBCddaLuF8zKcrBt0HxGCGimv5/s
3OpW/C6AoFk1czNQVVkXXDB7yW04NBm5Nw97/Q9WP6G7i6IWfUXLranxOx2S9C6g6p524eA+eUNw
KRLLLq+oxlSGQTm13O8JcoOCY0FGXKeq0chgRVLx35a/Bqy8EW+7MTH0moHUKuEtv8BXz2stpXze
NLQefbh2iIy9a03ecTUNVS/w4CHLIX4tPl9fmdZxS6Sg+p41i41JuWIouBwP8PKq/ZnD5Gy0enpI
S/T/EM4WcSni/iGGgm9nw8xtNJx3RBW8f8owtE8CiDxO4Pb7btl+ftOufZxvZP22/ebFeXBeOyDg
K6+11O3xZVYVzM/GOH/jEpq74Xg3NQwzYXgLJD4CC7T73X9bDKm4kT6vx53feOEze6ZX/n777yqo
JRmsRIPtPbB1h4HCyVZvtPrkul8VP/Bk2Wsw/3kCVSmKUdVU7oyd+WYMqFrFG2zuuE3e0OSWDjcI
SbG/vooxW+jcJtjBZyVutQbrkrlaByMq6Q/1fu/kOQDW28pLP3LegWReSfjQtMnGHjZPZrPrfpXO
evXEA5A7S/+TxhwRlSHqEnziS9y8WM8X1Am6oLbT+lI2saG+Hq5etOVN0kahX1V9wbUjg5M1ZIGc
XC5EzCFLkrLW3IF2T6BeGuA+ZdZaQ5TY34mPoYHhZSQypFOfrRqk8ACqgMgVzFJMbvVJ6v9Emo2q
BeHPKfAiak1wuYM3S1QIcpql/D/WXBIo4cTmh0Y5isnBXPj5QQwRX1PFmI09pU6qNlW7hvNgV+ji
A45BvU7cluO+k6oJ8I3pfIjZxYop5GB0f5B+r+AqW5JDXiu5vSTctPysGmRf6erKE8z/FfJjE5yh
M1PG7E4iDv1BD0zQaC8kpZw1TYZ3+QA29+bW99nOtvf9i0RhzPjLk7KH7/M1C+cmyzVX+tgs05do
xab6VGa1bfwxa1fGKTdhRNnV9P5BIEPEHQvcARwHymdfQBqSD0gkZKqO6US5KgR95JTqRY6PlU5l
xZCg6UxWu52TmJlQ1cI9TypfUMDjcBWGO95mpL7WZtF21hXaLDhxlQxJXKzgxZtYeOzHMTsMmNRp
kl4gc3jPxQK78tHF4bj9wbIITozDBcCP2KJ64ldqRG73rVorGsVo2EuLIWez+qjGyzQaDOvFzQ6t
jQzLhRPd7Hgn96uXtL0xszZC1ebI2avXt54jRNFBPUa1xEZUonKxtkMJOMeNZcjvEZ9FrLCbGlz9
QxIg7MgecsJurL/B/cejTXIoEwDLZ/YdIpQGiJXT6hLsw/ztaYGKJTTgmV/x2uXDA7l2m8abwW5t
8fxZ8iLwJ2uZnrMYJmLAC7UzPI/x0OOAa9TjrLytXsK+IEHbHYAGTAcGPpwWmocBiFZh+bMokKp/
uB6XoEIIFM2EpTkjEMDPghKxCk1ze1IhRDx1JGcC7+XvdTy8mgiPdQdKEoKB1zsVLpPB1lCniyIr
YuKKLgXBrWm0C7wa7TqikXs4QlZUewjZZrRbvMpyFdkEOH/CfvANwm8pDvE3Z5hVQNvE1UFuHEch
HS4A/9qneimb74iXzkICPaaa+BxSaiH4siMMNEsOEEzr6Kg+MelQptr7yjU3YcP4uVnTRDrbnzBp
WcKzC5tj8QmFccCmSOzlQd9RXsoMpSk7HgIXJIx+1dnteAUgvPh5lo7XJB68eNrsaPeFJGIY+o5F
V6sp7eNuAG8a7k1GO7Y97Xmo+19YTZn3BdCda45d+9ficbQ1dhPxMyfhuevw0vTjdfesy2mt+hYE
Lri7Ra7Ig7DSLw8+P2wOVGanj8tvJ/NoQPpbHKgb1nUaUPaz0Ufrk+8NasQohVsxEMMXOKbXaNbt
msy4bOhno5DJcnWzmEDcmT8cIR8ZhMWQgYtwfblRBE1C7g6pWrbWDaTpItTJBIemh6Xd2PUcF/Iq
goYoEo4i00Dctyriy0QeR/WHFHZPaflZKiAuMlUzkLpnrxYM3deaPe0qrXRnyO5wmatDdPuGmCVj
nelB734bJyHepOVZfdHTxehTs3/UQnPTtcuO7lSEBre8YN36nrfgGHMAN/ygeTc9OKdfocH3QLTE
w/abZERDLQ7fgLjfYMFgvglNDdYCe/ialoSZtYs+hKSSvbcOQx7hov94sjVRsuer/fKOl6GNQwPA
bn9XIotMEhvbNl8iBVD/zgOFZXhbWE9qU8X9SaK0xGVseX3GZnHNO37tZzTzdQLzwy0MdzSPcaT8
Ae8FjooxArzEiApiUGwk4qW4noLcE9lXYDtm2g+AX0/RVpvebjQC8nT0FU0jV97BhwWejaejfOpq
/FGl6IYOdcEJeosi/yfL6rh72T6n0hxR+kp9yBYd0ZBsXU2D8gbS5D/X4Yi5dlLBLrd1P2srGeu0
gys/JVEe9FwccNDovrCZDv4bWvFrQOyP1jkURovE8J3N8u6p+HX2B93gf+mLTCAS9bTfpg7oM9R4
X1X/+CEuZOEFRppdKkG2M6e4uMW4yEvudHFKTHGDimiEBxwSqgdzKaTx7sfaLrqSEClSE6aZVfz0
RqLK2WsqR+fgEf1gia+SLjx4YydovvOVD9XIx0UrfJw63IcGcaM9OnqxlQAxZaMmi/7iz0OwxCmt
4/buYrK0CXqVCsAhGgh8qQVmqF6yhmfbH0q6M6NOyBGVvp/lf+b6WbFTG0XonhELaHWRXSoFF330
ylBmmJfk8mE/yayw8uikTIdjffXKgXBQP2JK58yqBYMdnWkhi768GgqzP+vM8bvZKQvJrm9A16Un
5GRYSx32gMSkzZhwP8dZPrTzz7Ok78t0FRK1D4NILYYsQDm2vsOzZrnoUEE0Xp5ydzkJG3hz3eZV
hCryKbqB2LWG6jOFOaSrjU56zXGzpOsJ0wwChQ38KhjhCHUZxpGp3K5eC8YwRwHiPmUZFdZ+QWx6
HfiA5nO3tyfBw5TRYHAl7+D4zwfbmsJPguBXUA4xz6tmKShGe/7A72+IvMBy0RZKrzw8uYoeyOyV
n0lCW89fBQ2VSrhuTZU0vHgtThJ5TxQZD918h62+VPd6GNgHnnJ6bx0iI7n6YdB8/FAB47lkWEC5
jBxVDCWbkv/qedgVH0/Mk3sAHPL2czN4tV9z80iFhUattOnYXnmQxqCWrRnSh7oXARpnBimIdaZE
I44XExmVoyM79qFXNfycFl80F6mjKIjbfLTOyM+qkamN0jGZhd0x+q8eCp5Rp0Mu8z4BN5YuGHoU
4m5p4bb9oxz69DR2IhTo+6SrR/T+0L3mmyVegLsfo6fqU/FfIOqwkmmhW/5j3bDg5AMJiuBurK19
v+w8TMTwke7Uw3GRu4ZmRlxKJSqF9KQIfZzHHUbwImRDCasktimiTZE2YQ7cnB4SAWSnMKiB0NDB
bKpiFi00wx+ySVYeA/mbY2vFAKDQU82fLNJe2MeEyy/poJ0RDqnxX2Rienb2UavuOY7FZT6/X+4b
dLJ0yUr1D1U/vf4mBk3BxcjhVJu18l4GaZBXawCGQSPDwQZjF8HmgAGAibA1rGwkOC5wnmTNewlq
LFQBkq+cfspdQEoNehHxYWnX52l/Zwkui16w+5WqROP6qQlBW071AR03DZWdcMsZCW9hThZRUVri
L2461eMyCuV1oDl+/5egONspYzt2pwBvlUDHM13v+Cq2Mp9K52zTQmRzvqAlB0JDS1+54I+/WSww
KgR3jLaF1RSlRGCQvr0333Ih6Tv5uOiDmO0qUtOislk4N/UZUHFpXhiIK+Oao7pPTXRpZ6ACS0W5
PuQwRx6IpuCt9IemEmBjhcwn0SfTCSK5V6LBXIz4BQWPlFFv2ghMBeXFOho2QWxHyULnO/jvNZdg
Jg2Rrt58ryzhoo7vTK1+Z8zQ8O+VZ/5AVYYPJsKXe0+bHD1MmVBagojavdNxgYW21BgdSJtlch3L
VdacbgHjZIHdvhr1N144K5fRL5L8yHK5zmctuUUyyeNTW7FLo3HezZNuJ/EvlS7O/vnr4PkF7xhY
wlNcr3PVI9BE9TaaqmcEpjaUFy2B4S8d9oi56SWwFlq3OaEYO7dUDHz+bIz5UKDPIIYfGR7KDNdr
mRt+zfz4a2DuSyMuJ8Sro+Z3d1gXf5Oq6cYJ/e19oDwDa173RauYAo0FoCHJaOzxmwr3N4/FDLRD
Ll0zyZaV5JRyI+lPVewzDkGJiAQ5g7kQsFbs+3E2F4/wwmoibIErVVdNW4IBgbBsJJBep66M+ptU
XKBTsq6qean0EXh6H8BJ/82LVwirNxt036QajJpgxYBio+ZW+UXeInGYHoS/PHqkWHN1o8bSwUmq
j/Nmg111svHvePxhqT9kvlBOUJLOFDokNW+uNjC2zQljcuGXMt0g718E6nlXxxKEoCpNOEdqS+Ia
nuRp9nfuxov5Nok37MNTePg2VxtWXu/gqcPj2c8gkMFqngwOiY0e4+ZtpUWCAuFRn2dwyzByfLyr
MCZtB7bfFRLxvJDF/BoHtCwW9bwbB11G0u+7ort7rX5pvxG+qfCU0ytWm+qMXscNZtPbsk2jkb/E
k84RuuHbU7Xy+qgBJwxGxZSqEaqtJxIWpv/FwOJ82eqW0b/eMw9kMGOiaqtuk87pfLbIHmPlNC22
Ofio4pIANQ2ZGGXJk74XROzi5B31ggEeRGwGS+7TROw20oBpxJnNtkCwuupq9MAZ6/Rq4m3pFktP
2q9hdxRe3bE49OWm1z33QjgzTb6Doks3yBIWI5vVEXvKnW3eSYdwPVNFJbRlI25AQ128kvf4A0B8
txQ7FLkpK3vrpJglU9zFnBRHC7qs/0RAr1wPXNL2DjCTKYbiSwvPWwx68bL86I5CczHqo4S9cxpj
ygYM0RgqshqTOUirEUmQJq4Js+3uipQHrPxwm+uHoi17JgaA5C9Qqto5l7/jd8L63XAQxzboL4jh
oajcNmqOoye960tdTY7KiNMXuD9fzYmVNKw2sNg7hL1WO/CoH6XQG8YxTYw9+XF/cIVgsOWtj7i6
0XYYgM+LIZRegBX5jBEtleimzD9hbbD+wxgb4n9NOExFVUA5NbmbsQMUZOAl4OOubWwn3ZWe+jmz
aM5ULtkfcftcJNkOAtkqEIXDoV2c8j6Tx6rNH4fI+kUIlkRjFJGHXj68Da49aXSCA1Bp28gJtWDC
2Zuw4sGdgY1d72eJlH65ZSatXdt8WD7U6E4I3rZhx39cTtl024CzWbc/4HoSQWxTjsLVRGtQcF8h
2KEJKsWtiUa6V/csW20wAjXuUs9F7rTRUBI6NzS+Racdu0p6Ldt7iqAyBmSW3CNR2v1Ji4uVwMvH
9Pdy6lz2Msc5iEk5ENe1MMIGm7SlWPdpotTouQWvljzRSrnnM+txHJCPGIYcbpmzbuT94EnQ55rM
zgrjRNGUF/TXqUiEQ5+DcGSRzGj6VFbzBHWMqbCOmN8Laby3iR1BCmQKBfn8BlyaurYVVbIMdScg
Y0OjtAPH8K9CHj3e9+26EVbY5pZ06AZCE329OfI7d96ZqVnAnN8ET3zVzkkML08LWp1rP/ku30Pk
s9xJLI4ivFXnO1Rgd/N3GKxUbSAxq1Nze/g8zQnUiXDew3/UBgM3n9pzbBEz/dj+vWBKeQHjPa3d
Y2El8CHkCYdZGER8Y0JLBtZI6xbdRZWOFPaFryRViBAaASOaRTCr0eXUsE8e5FaELz3Gkivw5MEf
YH1ligeZ5ANFKiVDI+1JK1MQdxc9eFenMS6NJdr9Zdmy8UFBsEpbXRx5lpNhcuxNVyNVkdKbMKR+
dDUjnpwxaouBleT4MFXzJGfE3YAv6Ct9nSLoNk45t1rdQirDXM6WtNOGFrkgcDGXEKZUB29zSliv
vgX1FzMzZU002n8a0yUszvN8PWyxnD4zfsM8xWgVu0xrg86yn6fopY8/P5xQJPijwq5R2visy2o9
bxIu+LKazv5V4TLGkVgGwT4fkN4aEfqj3vp5ym01TKqUKzH3WSeR1HMR/GJrsZ8VL7+R2WEc336d
MvOw5AzW676N7Ei1myRIiQaueMTpZsFBbqbPppOEnmuZnKqTmR33ym2rmpEqwi3FVzX+yDBC8VNT
BFLVB067AbOqRxsp5dF0UmG5Dne8hRN2g8V9GFQQtsLT1F7It/mT6d5XdhUZZX45t/t9wdUwilBE
vs1CbkXnVYgTC4fk+nqkaokWGftD4ICG45RnViWaCx5mDErOpHBFMFfSw7M9dPDnS04ICMNvnkIY
luNL2mn5zWIApndGbJYBZE+AuzpkeNQm/YzweAkl7tOywb23YhYR8IBO+VpNYhZm9vFs9rwz66Tr
vU/ggEdiOiR7g18Fxiq6SGx4GNPEH080QxbkO5f/2wpoRvfs5HJ4Tb6RAXZZkVLlAqO90W5uab+D
KzhMGUbOIonxHkPffP/RyQMon0+szHHD8H5iWaqSB4s+Nt/t+DUEKwLj5JWCV984jWa/BZIqScP/
kS69RWFXlZynJYe+cNill32hO3ejml+zZ2gnfsX+BNeI9GfV+rN7N2YCePh0m907tl3Sxarq3csc
vPlMWbX7ApZAQ+aDiLe9bCWyXQAUc7cevqZtGoCpb5CmAQrlPOzRCtgFl7clDncIABGunUwLUyXA
FAHh4BZmqcB1RjgSmroZdBlnq2mE1hYeGh8doqCJDNgNLoTt6aSn8o/ndTaJjsB7B2DEY0Z7yxkD
kbd8jVOZaRaUn7z0dVg4VTwj/Hx2VUGknQsvtU+WX3UxF+ntjt1vbiEm22e/u90RTqNpxhDnRSnz
nBsUA9bOHiPYqupsRGVmVFG4sOBQhpw0Ho2IIVE3kTnetIoqGK1S5+DxFroH46fI8SZjRwXaqFLy
+rInJ6/CF3oZ/8bo0heibgk1G0+8U2MaqIPQtDE7rw5n/FJSiP+5bZ6jiBoPo4WMVzjVIscNBy2a
Wdmh0ElU1p8X4x+wSAMY/gwzVne3p2X1tnjO2r3GFRsCfXFpkumDajY5arSwgacH6wH5vSNmsEP3
jW/56ggBtQOSeFt9QmwFsVevGJz9rbEY/JEhCC65mFndY1gDBP/SbzRD14nfZfvsGpdTteXvb/yD
Tm+wde2+VqBBlZSuIyOqHpIh0bNKJMlmq0yKtzcYsrmUlxLltlkEmRPNBuSH6dhMD/PzRIQuWzgt
/K8y9nv4fk4AqD69U5/ft+Fy2Xnfl50R5FmRkXUla1hdtGyVEHpHpm2LxDIzvDIUJFNndyy5g1DQ
tDFbpWOD0RJV/hsigLHLh0w+rVnkIk0vPFNbtpEswgh/k13md5iqECUhcrcL7gcoZ3C4YSV2Uurq
8v0bjMN5eq+1ueEPIGn2+faIhvc+Aw8QBUmSYy1ZwlPkceYoMsrylBD+cYIxsptxVojPcPYalHLz
nzw6kQrufzjDVYqAcU1ARI2cZV6vnopzcXR+LVzo8ztp7Agbkcg5NMcauN4Royv4ZH/Bqj9BI/JU
lRCa64p9VS4SQiS7T73bincu0BgnhSRKsS3vdJqfSeSDEGLRdLMUCucFzllwNr5BgnIXty5/Z32T
CV2wAAroRwpkllZlN+NJ0tF+BKAGHQohsDKY3pRlc8fVsZw0QsUwY73cMWqZZ39iWAuLQeLYdDfm
mTzA4FcHdxt9oT5a48/oxJ2v8JxJYkPI8A9w0q1uOJwvemTvMFLG/2l82Q01zmGr9YqnQ6h4eQMf
SZzjsfrBaDpAXzMPCR9B93pBofD9kS4qtwuHW0bifA+UWELzoO1d+A868R3JZz+oXqbYfNKavHpX
9j5dN/cjRjNwmVR/JRYS4ud4v31ZYmvLnblqCYO4Dvy0nxAOBkfDfxk9ksn1NpkNF+p7D6eYswiq
njyvc2mRoMK2vdRPtqbU1LsDdHsbn07+AiiriJKzogOx0ZhK66EYD0KFeGvKmqRvTet9H8/iLXFa
gkr7y7YTS/MhEKvO7LHoD4bBqoAgjXDryGflX8AbwncKE9X7d4ZWb6sla0uWk8To6c0DbFQaYcyD
aF8QogI5wTZYGXIqFDWBUUu2+mcja54kM5ZpfTT5Ku8NTPJdsfEHVoYesLARgVITdCKPANXm5Zki
7Q2HYKrsz3i0tdIiRLdSemDRiTGTxPm3AYITDvYYYOvurSinbUgteHuD1dAInYX2hehGE1l3++Tp
jEeK2dR+j2z15KX8uLDBCfaYTQKbJft/9D9VhXodIekQ6SbUzMJYuHMjaal2LcXBI8QP5aleYFKw
tG8Ncdn3bJcg+lu4Ly7/h3CJ2903DH1yJg0UpLzGuzZp5AeUtyrg9i2EN+JJdGzjwNynCfoBoGK7
bOCdnRggYJwUXDwu+/TcTr9DdBgs2l6le1oA24p8ti5DDFwsRO5vd4YNJjEd588WM4pInuIdpxTd
SREPJtwkfeHQUcVFJpgKLtQzPqvulX5KDJZT9D3MKu391Z37v3gs3WEuMbt488UiCnuL+9jKc3QB
ZEb86Tdc5/OPe3z90COr/XDKFcK0Y0Kof2Lf7n8tMJ+M8WHtWH6S6e4z1FYCjm645GZ/hhmwKn7C
IJY0+gozbbiJxAWjKGsoemxoTbrmHkRLcgrK/saL6t9K8fManrXq1vgBIpdWGeLjkpPfB8JWRb2y
omwOWZd7+ovp8UMs58p3aVCXW7cPpfdH8VqXl3IfWHW/y89aP8l4f0cpvBT07AOdgWG8OlgsUEfj
e9osnw9RVZl606D5RvZ9tcCh3R6kx8HnaY5IjXdpoFeS/1t7qSp4xmx0a22iLbEWCDFhCsKhZ5yT
eQqNNXmXvUeuEk8CmBU9pUaokQO14brb/LNJjeNbeCoSJo6T2wospbGoFn7uHqeUF42KWUA9/BNt
cvEGlqFMBMrxgHfnVFB0jTruPBY+aulYcA3b/bZHXs1mV7zvJ/PKQPOP6T0Zhe/ZIuO4ndqWtyiR
w8jsnwi1kJ8dYuRGPsO8soctpAUdRucxSmAc4jrK+eeyp1iVePHD9BnW+pldqtPk63XLub/x3q2Z
fA4XOHz0cZQo+xtFq/bsrHZ5xuAAvLP9zG2WVtzoOJbaHWWox4+BPwHKzx9SJjoDNmo19Zs6FbfB
faqCOmyv3CIrZsRT53Sm1ZZ662ojAKWI5Avh7uMLECivWmJ9KKOMxQ+K3Pd7rAbQYV7EBFpkLYDZ
Tt1tixCaudbM4WelUUXABSyLpDaXbNAzktxT6/ddHhyxyAlJub9u1Z/TPrppIqYrKAedZGvk+wKW
sOoclOXa2Kl7av79eV2SahFZ9BxFXBnOJjmWBkqsLraMuZeqKPFWRWnZ7Ypwwe4Hfo7ATLghXvY4
4Z3C8dH935gvyUDxPRiyXKn5kB02xYc7zm6rjP/GXfNqcDEJGy4PyxplZgIEKXYo73QIIBySnexA
ldsp50cJgfsl9SeSXZOa3Y0TEKn2stb+mJM99njrTEeh7ZtY2Tyq4ZGUD+hAWLdBeHAAcpSMGCv4
EA+2olutOOzDLKXeeYddI/9MxHEpOBcQxvGthY6tR8kFK2T6TB5g2xOMFPLBbHwmK8MLoAEEMM9O
+xLh8ONRTkPsLciivsYTS5nxMn3mmCy0dh6qsnF5jUUS2bfcOmkyvppso6hOsCz9Kmp2TfanltTs
x7GQL9BsnBA0+Xf0NxVLhPeFh+/RahOuHrCg3WtzCpHDG3zwFy+ATC3TJC/Z/guGsz1LYm6buo3q
uqh6qsNDvU4Ziav1CCxtciM+FH73E+tie6aFrqLnOgMlD3uxUkbNvaFywCio34xOP7H12iSbWpXi
V0JLmc3HPriHT0bCFo2ThlrHG14YdifcMQJ86268qF6T3IbCU1DokzpzmLZMW5ZLzh3tDSeW4y6P
JvT5ud4Ynj0VOLkCKlSxLdHoT2jj0CL+ZYRlmHSL3Bkf/wmR8nMcprAZkOXLibj0uHr5wuBX3/ce
5rFgbpu7Q2Ah3qAzGXXaNpzEvfGKeBonLIVo57Ebv/OhTjrivMx6lSATYe29YIyOUfCnqz1WtXRo
2PCtlTrQZUa74JWviaSOj1hr84UfgBAOzF/yS3ribxmwW4NjI7Y01+Z7wSrNwKjTcaznUjkLOwRQ
A8URB9Nt0EVb6NMmogd7U3q2zjcDpWrweQS7UwdIikh+5IbPVxL9eIWM881PGsDjyzLyHTVJL14T
BXlgowpgYkzJzIP6e+7XUNmI5eaqMCJlKo9mYFNjsPju59Xz6t1fGfrmsCNRTRtL14OR/F92aOKo
Nriw/wuQ9ypjx6Kwcy/hGSM4xC7ViAasqNIukKUfr2Zbf9Jnc4KNWU0NZAlgH/+V882Df+TOXBV2
5J5H82hTOQoVe5tNnvbg5Rxb/GvTq57ozA2lg7BfPil1FGgwIbuQ1kn5/RsRrsYUOShlds4KnzlH
fc5DkT+xArstdG7uqefRrEQi8AwL+sI1xNUvYExtLbnuM2lUlqcQ1A03GoTrBKCOVovBc01QFXn/
xvQ7hl8l9YXlLY82qMXruykMYhpONcVTJMTvR6l4jTSnnMfUc1Xdw7ckQCwFkyrrC6USrdqzxJzs
fSU/4eWNE5+41GXoOhq3wqL4hZ2wlM1Dnz8h8KHyuCaK9Psb5OajA7JmKhiyYLxnaNotE4y/5BKY
ky8ZXST23vBcpnDX89kMPT1QNjIPRmd5BWn3eXOKRhhGNdBpOf8iRbxapVJGab5mzvET1NX+lw58
5KIwFZR0zEtIv9hcttduJ6ltyLprY62wkyiHHzhklmMws8PLzq5KvvpxXe2sGxqpkANJEigY5A4I
eDHz9kv9QdyK7i3zifG3poORW3BmLpCUqYY0dXlkHU5SIglaz1xCYNzA/tLlvnvS/2sVFX2nQbcT
NehAIAswzSJCfGPoo11N1HzbZ+FxB8469cUQ30uLowZy/JqopRBJEtmWX01g8cRVgOTHISeTSo9u
f2b6JIl/Q9BO2FQd47z6rpqjwjsHAOH7uV2uy88xWxXdL13V5k+q69azm2T2+fBpQmTuihuTFUmQ
FLzAG4fKACNTz/+SefIlHk21eyL2FJHIJ1cRoLkVCmvr+1pG9+9eyjlhyD3r0mcGQRw0OqdzMN3T
pJlOV1H9bLz1v5dbVySs/BnZOiscB8F912xzLybI0sOKBh4oWdZKYu7e6blmb8CpcQVdlEnUfpYk
nf73QG6TzhwBbA3/j8Hps0wj4nnoDwAArKdOEtxHl32MMPSKyYpO/TSug35kpUPwRr79ddrvDFQD
+igBLbgdS2aYNDohgMB0W7GDidLxI1fCeVIo4htLpsgVM2sciMZxUDLVeNNA2Qsm9xZGyR+nN6M4
5EunNY71vQ2kZXlA+8z+1XuDfhjf2f5LpC/wnBL/SCfUJ18ny+OpR3bF5rYjiuT39V7YXANUzlZW
YveJNu1hgLkT4Y0+IvTIAkhNRpEMEpk33JTHYC71CIKNRICPXULbEJmmJ0asbmDT55OMB9OvBrfB
6NZGtL3TO7XQ2dfM/vWkJ45I3ewKFn+iVcFCDNQkeVZF43F0C/ASPwasgmPncCa+TMOr1rIkebSk
pEAwarsMfRIH/ZD3j5EENnaIGJn6lDAKhaGTi3sjnKhTDjB2Gr26pxJkOYwplQudlFV5i+brjL5/
mZHCXVt2W2g5dEAxjQTrxCa8md9N6JVpYXiHDitO3klaVPeiaE8UUa2FIOKqS52T3wi4qiTYj1nN
S29jaLgMsfGIh2v9BqIbwErYFhll8GXxO1zEqpL5XYQ7QD7lyzeMLBL4EmVxNK5849CeHpn1qFfI
1wXAi0+Ker8yPZhFdjLQTaMhOrxD9LJ7l0YWMyFdXjTiQnDAk4gv1fvH/zr5DITEHjy+eAq+qBBv
vGT9CDFdG7dVeZ8wROpOObyS+CW0SZHY4RdHeVGhBNZUtxX142IA5UPgj6TFiUfxuWpM9XcWKm0w
ig2eiZF/W3btoO46jv4+SsSE1H+mBAWm3nrCAQzRtJ1eVjO9XXGiR6lCVMCTQTdQJMfOUuxXPiek
HW+CZtVUmxrA3fYKEQuxt+MAOV7sinF90y/5AeATLHybThjcqmsRcIpIKQVFI5T1P863ZpOQ6YcJ
t5NE52Yo2GKneq5i/KNQonvPycqJx08KCUVKhS4HOAkb4eyMKxb+rBrwnjdvHdtRhZuWuqIeq0Xf
DR4mFrdv+Vm9eT1LJsOqUODeWkCSuRjxiyclFNus0gjNIoyqLI4drHEiap2iKCoerM5pG6ozZhiv
h+MfHk9KS144es0uZmuMdBNTuHZvW2tP1XwXf669KWmN8laYtB3gt+1t3KIlTIx+pNL7Gaih5W8q
jfArydp9Hf3DMK8ghG5TEnf2RJtIiH3Cv3mLV0hmjadKEu98AAHxbCk5jtQBGOVWLYYss8cOXD7L
YSt56PUerU+1GlmnSXuaJjmkbdWFcumVTvAZMJYAezdLC7N0USzCcBTxD/+s0r3RftSbJjWTOCTp
VTRPcakOXJ90sREtTObGu2vBYMQADxcBjcjSStqf923NxNfLulQc+64HBt4wntgmiOFGIZZX2Axc
gtEv+nnJ6jYd2nFrjQ7A0rKPW7lmgVYS/4exBhc1VtU8Xpj7jb1+WgvqYHZyEjUw7bX4eGUm6CoW
LEFZTyXrb67V7MsUREdGE2EO0tF7rVIKYxu3Kr78t31/1ci1u85nRDAsEwPYRK1ay0yEJ4bUwizU
AXYErZNTevSZirWb9Cw6MuJ4n0QEGYUrNoK5fRxwvaHYbYHOmUy4BITgEC0CSYUf0xP+vZwa0H2U
lFKv3oWb53PZsaKibqqvEFh4W8O4TGCaGEE77fM/nyZLlLrwsUgaVzsjCt8wXGSgpI0JFqxzzzly
rh8eDf5nqkkDdfkGA/QVlCuMd/1B46Bpq2q32EF/m10EYjMxbZU8JPVWdAKP1BE5pmifnhzr8sSV
MMr/71ib0UWU0EFOSEuTPW3G2b5/HM8rbgZsMcQh544NNCsQKx+McsftJu5V/qwiucxnPgLT5XTo
72tUnH/OGavJh8bkU/+oPG7TmwcxEVwccG1mH6O3Vwqb4Wf7+Y16GJtm5uo5kTbmUFGBETYQnI0s
/cKST8oZqn05IP6Y/PY3AuKFibcgaYOzaQ3QfHU5IqNP6X9Gp9ZnSUO0Xggs8vE5utqOvsIpLuk4
qKnHxSol5JFGGKWdQReCC9ZGSDKXJe5tlIcf0F6p8M32sYmaZ1oiFhnONNLba8bS29Vx6r9o1Jbd
RPnvvorQNtoZWflPkJXZ6ATDBC1cO5w0Vprpy5iq5GrYNHRYLpUqTBs2l01Y5NWNYkktQZwh4ZXP
3HvrTwJP2qeRcxzFBi706zC6nppdhjju24i9Crt/2SYohICWve7FjRMQlWxaXc09BlE8Q+bduniY
drOaMb8xvETXYP5SK9WoN0eAPFPdmsKwqXjy/vgYGgpJT5zMfCvKgfO06UM4ASa2nwbspV+P3XZm
FXj+/mzwdaSG5fij9fhQzD/xDSfq/GHgw6ia9dUws0bWszwmVR07J5yJWp8UQO+cmqHoGYU3Woha
CSSlF58iCiziTJzCTi3dkzzkZwBkpc1hePyHXbngo1Kyd6P51natHhGvoiA6HyK44KBKJmfyAevQ
SvxrIwgUrDvqu0cuUs+9fpfE/ctDeJJWrurGVQwnYA+he2nwRaeI/hQBwR7LdHQv7kSiUI5K1pT0
7UDuXSK2V79kORSfxdtlYtpsA7CE76ZkiT8a3HKpjrU0wuweX5ZeFJHYW3TNoBQeuRfFl2D74y1m
mCfkUM2k/dEdF9J8uxpJS8yWUq7CfmU8AtGm8iv3J79yEpJ0kOY/VyDe69Z9XUJbcQNv8afx7i5N
Bib2jcoBhkyHnVBJaRML7Lz4Is/8elK5Od6TaTNREYVu2kU8/ATEU1Az8YnSxU66gjiOI3/0XD/p
J5pN8b+cTxZZlyr1Y699UmAmveCeeIKcbyjhyc51GJSaxp6ydB+vwtvouPJ+JG9mBvtB8R33KvNy
XAGOzEfjyG3M2lGVCnlmaiPZQg9wUtOJheDU4Pjbuv7z1bPVagWQYRfgmUzziHrvjffBGnfvCrtR
5nu18O2nIvXSnDRESxxgOY7Ns98YzYeUpclPM0iLSOdVLkGsj3Iy5bbBZZinrrzCCVpzE5o53e2I
034ZBBZuqTySRpREsx0PtoWLLsEvhxV85X6elaM3AlvwlvfP1/fWFqyB9KFFcFfUbVMyHKlPWgYX
d769b+5ajEFwSOeLG9AoFB4iyYa1UC5zpsMg+TqyTJO5kAoXXK0+AnTsdR2k21poVXjk6pcWOyDi
vXdsRYYw6X67XNYPz0UIe0lEDRejMRbLobLrIAGIIsGR0b4m/DOW2Cd+payyFqy7JteFKnjRZd6d
kCTSoCOiifskSzRBgI4qOCfhHdvUlunnFQgyzrRtXZBGFbbtgidS00w0pWl6dEMp46mJoG1QQIZa
0BUvecmBkgDFHAh37IUS2CalVZ3vtHdIzY0u7mPgHvw4z/kgz3q5PotBm8nA3kZriGUfbSQoo68z
XK0KRkNEiF5ZUVFUnTB1EWdDHe5UmPRyuaY3f5s7djlJaBOUAL0qkoTioVaivm3oviGqwPhiYyGj
3dM8lfvgvaJ5M6PnE+gIcS0TVqW6zSTpmeAF2EGumQ1rkkkQ9cabOUFVp7CJSsketCQ7/A4ZOUcX
wF3rKPXfOts4oJe7GeIWHGpzxs9IwP0mvIcDnN64vuM63ojN1fzV0qYEandDm+f1aEsvOAOIwfki
4KEJM9mXLfnNO7rRhvSKtYGNzJNRnpfmaQ4CZ0IOhSCOMyAwo9Z+/g4yllJNyDE9M16EO+TRQpuC
HmrvVzdEFgnBaS3MUz/EvtYvOd4XarjwEjtwXfuCI/a0RQ1sxenln5v6mXi4G9tEFwI3dR5uxkHk
NIBMfRRrahD3iKxDwUwiG96+6Qp37d+dU7U4MkG7TaeUCxIXEcPTxcy0Y+54rWNIqrITt4U2Ijg7
ShMpsbNEysToNxP/XGxq5OEJ8UKtBnoFnweCSfgsX0jxbLC3d78n5LklQB3eG8LpApiLzDC6IAmM
Y4TX8orz8n+9haygTyfbkIe1hvAeeYChUm/lXCBCyyi2rHqYKdc0DZ81rQjwbuprr3ee1w/uWh2p
PmtBBnujl4I3l9LpqpkZY9/m4n4bIu5ZW+V+DXQYkcjQ+73Ibg6F+ArUn3tmw5GUGBiSC/z5lJm7
lOLX0zVWx/VOFYUnSuvmQ/N0yAlGU1xkkA2q6JCYXaMv5Kb0I0dEpr2KACOKQy0gNjrrNcuHUYfq
f3ENoh/z8nq+ebGJ5QrbEqBVFb88TW+0kSnQkFXNjS/zDs3HIRoFyiprPTMOhOZn1j3Pu/ZBpXzW
JXj/+t72qv2zhcXlyAmxSwysielWavO0gflGUEhOeGSml3WTPJWLaPArkECO/cmU2PRNilzJHDsA
QJZpYx+LafayA5cRQGmERlbteS6r9PLUowp7jmHvGBGwFvccGa/LDuXfbRQhJ5aIUzUXvMPFn4RW
HZWslxnnztwPjPFLLe9huLVUh4bpmLmA+X14RUQND+W6ixDmr8DgKVmUWFneHICb/q80HdGH7zBG
Gd3d86/eiE7/RsrMi1q0oS7NbdpiSlpnsAlpYX6FylP8axYLACtkdBzqn2XX+n79CY8O3IEqi6ta
OPeRvNunxO4Pe50vJB6qN/T852rP9B8h691g2cEWnMXnLJfpoCezxzthdLJR52+2rmmDnLlrNlXR
55Kkx6XnFSxNLWXHTHQDAd7NbO4St0hXsra4+LlHM0B9dBhHxIt9KUjvANGN1hAJCNdRCj45zkYR
zKEeOw7/ySiSyHpS8JFhlFa/oUK2Fmj6BUFkAv5gzrRlf4oVcxF192hpwXjfVSEmvoprOE0HK/X0
Mo4btAovPQ3XXOouylflyna2RacBHNmSmcGXz8SZt2PaEtGY5B6WW7EG+HK8XWtx/AgXLxljpOtV
e2ho+7IS/3aJszsSSPc1jX/QZe+9ZligF5u3Z3g6G/XdWSjia6StIfJV22ibbKVYEdmPN5tCUxEu
yCj604wpMCCrGugsFpa3S8UWSbJAG0AqaZLlQQlDoCa8MD9tFce4Q0t+3JOGFsdE7CqcHm4ov9mw
WW6eZAMN24FrvmOWVqchkyusdzJpHNYqkvNOUrXDci/fOZg3HSTobcIYtMf8QkxfWrdEHKLa4oRs
EjINpiywU/+RdrqdjlUKcW9ngZJTvPj1aBRkNLivgtNihw+oY2muyTbpzBORZx2JuQVt300R2A41
5PqfM4VZDd7AXYPxQG6RCsCjPFvb7sF1B1CwDoONdE3T1fo5v9DJiIGjr9hcMGT36ce34M9E8twF
KKNulESS+aD+ogfy7EBdwAbGq4lyShsd/m+fqJmbxFlpEuSeCWC6zzaOvLj0NbYcgfOV/iaTP0ms
njHfJZFevHMSrYx2iLzwKzGozq3WwXif4vw9vxizxxvt1PrYE47VbFyIszQR5ps2fPZA5fEbrK7Y
hqgaGasxF9QZOINoAtVW2vyqbFizk2KuF+L5RNsiknJBdbmlkKJucR8o0I9dRJth3tuzGDyR2Rme
FGGbHg1SaTHPRciw1jI+yFu6vB8DyCGVNSEh9QKaq9Ut6Ta2cAdIz+quP5MsWDEtGHHT4Sn99DgT
gYjMGMa6TMxGjk8QxH2zds8CX+I6FOpS6+KIn9gJQlr8rk90ZSOVE1mIwj7PEGSqnLBffYFloYLR
E0FvSrBSJ2wo3fzFLnJgAL/VjrGjqsMHYpdrNM5GwYoUFZ5J+AnH6ep1MTJ1N7mJVkuHjYTE+R3G
0EpOultmQ6beirKRtet1jk3z16KJ+EJy7YBfIvqvXDZGUECdkgR/zZ9TWiQT/ZLgZ2FOYG2lxFDn
crUI8ZvW5OXEb+Hd6/f5iyDivuYcFUZ3v70FeML/wspgpmzx5nsYHKJq4TSdUxFYE5wmXHaqutOA
pEDF4Gu4s/Y3+14lq0Rxa6h2EEug0e+iOq2Ioft7+cloPJ1+vmW6aE4u2eW972xy7U6IHTx5aSiv
1XZWp0vdAseHcE+sJ3+k2lb4AcKb2PTJayeQpOSe5YIXwX+75QH0jDbUyt+NDqij6/Zeb3XW/GU1
rrGbTI81ZpkvlrscthQkjdbO+AYbduNfIq2gyWJwEA4g+yxBhsXJyB2i4uhKVO4LU7nglVz3Rviw
IierNwHiqIY0enZaFqV7PzEr/H02xNoPN8EqCwbilzTrd+GgQKHCZX6HLKO+DRPj0z3nQJnwnoUb
Fj8zbIfYKZVsyTXsi+A+M+gZv4GF53mHPa5KJ7QWW35G+nxwFM4dxFn1DKjMGUej5Gkjy0V5jLrp
lgQQeCfTN8/AaAxf6j9gUrkx0/64maNlEjNWaJaSinMk5p77E/Zi6kcpKaOO7W8FO6yxcBxPRV9Z
lpC71K1IOIjCsKlLhZoAtyZwsoqvnlrfop6xMr0Lvok6M0n6eDLet6Z+wE7YEVJDIuXvZDzfofpL
j+Z0jjpK5G7vmab0M8O8C70YPPgOf9wEONiYHFsmUCzT6rwVqPRM43Mps6qfe9y0aZAWhEOlqFLK
lSXtGHs1/Fl5crOj7dU3LncB5/Jhi2UURY14HURfcYM/wgXBvwKA7kXhrO30xZ59dwhyd/aRZ2Q8
yWccmB3viwUQ/9FzIyBVWDmPB9XE3ArUMi3pB4r04DZHy+2WOvLGez0Uk11JLyBMfqvMHORQFgbF
1AKpfJ8iOLU88KRxxcdHmCvJ8ZHFD6m5Mv+9pkKTLsfcG7I0eIfGHhgSppe17LwHOgC1f60kMNnD
xs42KaBgUWJq20Gwvll9eYqeXsl++PTSHF+zDW+l5EF7vbY6oQJRNI564Co0WCFIWsToa/Mh2EdC
f8iCAD2wV64HZAdNHqdD2g8R2QmokfMRJ+0s+JJCSENCOaBcSd0NZ5ka7gVFR+9gNOrE33OpEOnK
D06zdK6VhV5nNjmmZGb5b3Dd3UZq5cNvESKHnkMdKLc7udmasOPykgRAzGu6pFKjcFDpc0yrw25R
0DNXMegnDoWXHVLvHnjDtUE8XBHFWRlhYQGagwGhYJyzfKLWboUKmiG6YjibckWKmEn7a8dsRHl3
um8iE7eB3vkqtquXMUCwiUQ/htw6cHnXrBN4EsWijut6tDdwrHU1JB39i4h2/iqpG4hwITOcsAkV
lrOJiM04EZeMdCgIueNVR+oA6C3QEfmlJlfihw9LgMgodi6FUG/T/sx2iqvx7FyPa3Qip8SmpwiO
TkjWS2LOde05ZWyXDaUEZKjr/FYA5al5Ujk7b76MSmsu9JhVjAB18MPXOlXyTqFaP8xTJxGQyok3
rlUugIjmy+DlXMwC+iKDSM9jx++Navlyg6rJ7gDIA5rEn/JNG21PolDnjk78Zw4Mclp/blsHHvaI
wkLoGwx1vxRtTAQkLa9cgZX0p4CyJotl4rRLhJCD/8OIZFZHchGl32vXQSY4A9PVewzLjZca99mD
pN0JN7znZZssZNbqohoIzEGiQs7l6+KLU7qlTk1EAWh1asRN0dAH9pT/NQsmZI0UAiv+TQsSzGtl
xQmSCLqRN49af7d8XCFJAdwYRKYVbrZbreSmmI1A1TY+tgWrWpT/+8pA93O8F9sO751THs8H9jql
oP1tmP2qjavszu0/bfuphFC2p+M5690W1XQP5bmWYVdo/Z+qwSxkQcksoKXL1n1wMmVbXIUMFDPC
X0vNhw5hIsfe13TfZAl+CK9At1hH4PAMdPdpYOdIypXaU/cLMDCEbvnFvGeLZNcTClaVLhH04cPv
6eE5qBBv4axaQijv3jwk+INDjOZwTurPLtboyYleIj0Nbj9bxILPt06Xkx0jrMyzPNUBHQN3rZrS
Jk7zNyRlWLA2dIGmmlZaHZJfOKZOaU1II75UPQoEllCXNommCsCD/hI+45E5NVTW1MzX5ta3w/1Y
1v+4KwEOdQPcBgPWxDNp4evLSU07eSeXCGvTo9hd0IFKu3JUBewzu8n4uXnjLQTe4VWpz21cJ9rz
+SY1d1TSmgavlSR2OQqzAweYxq3yVHVlqi6nm2Bw0MPf+kg6udeBw+iJtSkGUJVLeovgSKvxCfyI
RmHIIkr4g037spcb4+avF99ax47Hs2akRZBWegeOpvFqfFp2mm3MvbFqNelzDJy6zfSqfFjMU5f1
1MtC9XxplIqDvQdot/ZSJStY6PCn1JRlbcQwjLlzP2g2fqdR+jzt988s2twYAMhnlCrUA4Jwklu7
nCDMlsCEE+U/EEpira+tDHHDNTFc1nfDP5dCYoNPOCLqVHxs8l7jaayXBa3uHeJg7Onkx1RrSclM
n4sGvnf8sf/u1q+ohpUd3PU/Op5p+USOW1wUk+7p2RCCxWEHFfwtXU5Ol1+N5TwLPfx7zFeYhMHV
dfjNbaF1StBOQ+sx3VxyucLdrDh79CM/FdW31bdmS9/w0ztOZAT2pT/xBV5YH8Yyb6eQRaTI3GuK
whzfxWDGursqMXa2psg8HRA/ONZXgUgWNnhqhEWnOT/g2wffn1aJ+G6zmGFu6qQJL5ABkPw+1t6d
rQ4ZZta4c5LwwhJET7OqEfTAjtTDxI3pDSwyNmueItWxonewI6NNnyZ831Elqnm++l0gOq8QzZg3
YbB/GCnsZ5yFkcruzITtXIIFe0hXK+9EMUjkb8MCCVa6Ygok8hGOYf/Cq/brswPvGLZt2PUqJWla
bex03c0aiAMnLegy2C+Pcbk2hHGkeK5gOJA+PUobPrSw4xFQj2RoksUSmS6eTlCNL3/gLM6BM9Y/
dPGL4OBgcQk7pZNjuZeAuGiKnUqCHa1hpW6dorhGl3pxUuyQx0+vGmb1X4GZgCVdG5EZxO8qPqH0
b12cvdzakgfFgsZZa7Fl7c3+bf8CUFmgZdkUtV7ogV3qOAAihGGIRB+GIJGGvYhsgqGOBhJDK+dF
Xi9LjzWfgw8JJ01IbB5C5EOIIzaoxMzuOERSY4+axv1bQSpkb653/9DCDpi8Hr9SAm1hi6fGihGH
Fl2WqxTaUND/nYE3FoKaMhXIigapS4Wt9qb6bejV1AVNppKutNNAtLuDnKmWE5uncSRXFIKY2vL5
FFiDYeg08WrpvSXA8mgZzOZ1jzi1GQI5lLaBW8iqSobaEDv07QKIjR0kz8FTkR1rowgMsNIPHEqW
/qVOOZhwKzPQZJKB3y6THrq5zv5t8vf2LIB3ugdGLkDg7LNRKntVEuEhzoM0CiyuyGF9snHXHzmt
/qyb+Kt+XGLMrWax3IwJUSDsVVKXgJ3YRseUAG+b60leOGT1whmUBJ7BMud+rA75yPs9esycW7zv
VsoaM61U8jSji58ISYKiN3VwwAVJKy+dS1Y82kAHXmCW+Ui3MOTCzKuCC9rJHJAzfEhULDk6moUS
Je4xJY0/Acs2RYKh9lhimPlSTprarsF6vBnHh2XyrYpDYks1tp1N2p8n7xQk71gJa9uwMnLFb04A
59kssPTIaoec6FeCoMkHTNPsob0tWuOVOqXXrft2QD9olJPlTZFObIo/+XJUilaae0qzIvQ0sCro
z+iuAzzc3+Ncv2Ybrk9nWKog75kEqzT7+zmAtUbPg/067/qM1K9kqe8s/umLsvwYW9DOGdGIbay0
1XP/8ppYRPBW5Y3ot2R8TamJI9yBoxjVlpohwfFMh18diqC2mUiYKceqGtfYVdlAcGTRv0rKZmIM
2Mzo/CpTlP150tEDHcrqlHcLPjONOO5VXu2KNm6rx0blTVLOu+Hg4PzfssDlxYSbrp8AZTkudtm7
ir2hbWISR9y4TEVjfIx4yiaN5/hB9+8IjU2REjlmeoz9VQdrXOASJkuOW3n9/Fm3+PJABulASNNv
r2y3WwK/9mOX5NwM0pus1WK8COsH6tALhvMYatNpYx4iEE3G+/is25lNjfJvzpQk34CYnCMn1SVN
LQ/+fwaDuUGyL6yTNRpSu3josjkXYLWLU3hr3D2kjJQeACgWbzLwYIqK0OKt60wrKB9Jo+tHBHwM
wMJ/6dQdzB0zj8XYGPsPhXu2QR89u1Nsi17m9nNQPKp4/qSiS30y4EnFcET8U3l3Lmr6FhVbzb3j
0tZ2C7IJQJNMBaXk/c0enlb1KCoBY+d6diZmiSIsAvuEqrKH2ncvxHm/89AL+AfqQM7OIIGpiK4L
JtYJ5C/pwBNL8N3eXFq5ujuUEOhNyKq5pDS9SdhiriSiCZD4wifAWEnuRvpuPzctTgYHAEew1iuA
jLMoniK07SoLFHArS+QvghRxBvCIXkkj2ePLmQj12no2pXisU+7oBvjqFFDFzbfe4zOVPjfgPIVM
AoneVZslHyrrpQ2m+LK1JdvUAlRQWZD98c7oxqtimUXM6xGb+1CYYLss9TR59JSFcsn/U/u5XI/5
ga3IbT/7drl1r2Ws3ChTs0bYigx/MNii6/YCUONgpXPf9HEC8bNSX4cBGVn3khtyMaW8Dwh+UfDh
7BxEM/hbhwP+kYmPmxnCKv+eFnEJU1yUwWshdKhUSfC29uUWifzOZOb3tyMsVvSFbSVqHNtIfZHZ
MH+Y98AgHdQ86QQQ4CPnoZg45+2Z4lyVPHpvJDRiQZVmh4vOGOcG8t2YtPYsyKtlyiX2+WGfuxY/
9Vy2CkxlMIFLO46bebJ6pfTU8OA4kfaqp1JTEeLwLGe0RVOOsialU80/rZyiwwjhJRUX0rFy+ak/
rRpukxjPW4RujblWJc1zhjS8AqZ8APnlDbkSO02SUTSZ7TsmRzp597C/jHsWTPDkBRJDdQyvePoY
VEWzzFC+85fWAMI9ekbFZUk/0vrDLkQsbehEjIJVVqCbk1Oq1N0DIXjWBViasVhr5qbiDM8rRv3e
Nzrzz53MMbFR3vegY4GPvbJgI8kORaR/DvrkbnN2EaqA3qAlmQiePUtgkgQeBqAYObATiMcdvPys
rOuPe5h3C52EP58714+x8oyfNpxjchVccZRASKApcUGm5LakTvEsueoe45CCxlqbm4XGA82q04Mh
D9yevBHDigHKxjebbpeZ58TAYF2jlJvbkSl8aDHr/WzzkW3V5kZxx+BSArK26b1h0DxhYXDMFGyC
iI31hex7uDrDXh63xGM10Faw3891G9/BbJKslNQI3gBENpkJB7t4e5R0hmO0MGTSKv+R6kGpZMuT
hfraJokdb9HA4001k1ySkd7wUArYiDunUvofWu27z5jEflaNXIWgQr9pSIRDGcuf12C5FN7pmb4T
o5dtlNovk7F2I5dtAC8JrkSe0JIcCZxzwYHX18ZxGeWXFV0RPGVOKM+XW/1cla/IDdFk0ST/pYKK
C3fx2rQTP+0uYxvDVzP11/B/c9Nrd37voiBoo1rptFHdpZxvh6bjLHAtb2LlQcbayk/7hlaRjTia
Nf/9oKpy8mq3WIh/97g8iz5CfdskcFjBDBXg/qiYmm9JPxMNesXw/u2E1JP7Y9+dE1fFokYONz/I
E4cn3zdquiGSU3/p2yTEQywv07FXmaFoz8hePv1Bul+T7f2YWotTQekAPaVhIlU4XuX+bYB4Sp5G
LFYar+q6q5imTVWJNjWTgd/EOT7T1m9/TSiiAjQtB5xsJO8FocuBR8ELoj+CZ6Eft7UhEFFJRhrs
l/VLOkC0pzGm6DKRnY7TBU9ggsxWgPSeJmHO0HeJLpw0rgOaPzBGHhyKr81UToSZ7ZRF6yZrGf86
r3bgqxby17WJNHtE4dEwtq3d95U2NywwK59iKFszmh9IbVlMgPW0Hv4sz61umnHZrZQY/ZiyxG47
lnANgifjAO5mVFBQypxTUPJRqjVfBp2x6UdSu53UG7ufvPXVa3qY/sDVOJtMdU7Bk7pXPD8iYdCM
XAmRegK8BaZtOT9oE0B4Y9fUfk0DYdXKT5Mzgz70qNrDdnHaPgVKl18QYHhOy+swNU/2JrCJAR5u
3q/D0a8Ve8oObWPdyLWfsF5aEd4ncDO/qc9F8EQsoUv2z5F9R99jlE8BTRMmWoPy+PHLvJoXt817
kHcVZU9njpmat85W7p+DycbcbWo267A3RPJgGFotfq4/L7kE3heHCjoC3WKcPc01qX/G03FAhN0m
GGrl9mGk018uI4xF3NwUBFB9jxs1mHmCeXj7J23XQw2+ge9J9LDwfDgYNBf3hwOiGQ+RgE3iNx1K
fosuB4FDQb7YPBwSHq6R5bDzyzbBVwE78vXkLMW6ROAewYiaHXa+p0lTp1a+DgtXlsbt/n6RBzni
vupsQtjYfslqnm9OZrptV6T9oEHod7PO8E5DzBEOu+Ax1d9abGqZ97vtmL8MK1NrovVYXK3Qh6vS
h62/Xh9Ohc40tZu9si9Q7/1gHDxecsJe0Itgt49sHDRI9r0EWmN913sT6oLjNGDxHZi5Ry0Zx0WF
4XfM15nhrtfIkoBfoiuQsFjJfo6i12oFOwcxVAumYPGEz0CO4tIoptm3XlfLlUbgezjeLbVodUQk
yccWUplkN2EVcuAOivHWZaQQ3r+S2I4FGXitlkUbkvvd5kajuVaI7YRsneHyI7F76tD30JJwC7fR
hW4SMu2Qq/5Cq1R5xt5Gi3lDNC8sBZXeGtqEmTwLdmBUbjTTRP4LHS8Dw5gVJTBMsbE0kFHNfAru
PypaIhQwhgvW8c1LKGBupcM2zJ8mmTqEVRtiEttQLHGEXmPtqr5tXpLBvf1Xjra58HmX1TT2iaoD
tSJdZ0wHojIhlUiCJsLRy3flKD1IMqWWhTdXdvwseWkGHGxS9sn67+kijbPmgumF6i6AJu6uE+v6
QB4TmO5Pcj8zfVQk5yNEQYUuunah5xWUVHfy3DGdWL+Q+SsW+qrqQhbsVb/i0n2uCxExejSXJgmB
gHLx/4RMNiUQm74bx59RCeZI7CGZkk7J70ZpnOWp+YTj9Vagxl3FJFNRDcJ/tB0ZHkvxPSbHDeDU
SepodKsX+Lg20EScBn/GWwFaa7KIJNLQ8pQu8rCBQ09SZ+Uw6rhtcLjz6TDU8BcYuPzuNnLKWQnH
RRDbabKCOYyiNR+7n+soVVebtCc+gYUz1vi7K5FJd7ipMh9iAg9kwjhZdXcHhvcEmEgMfdS3IW2B
kOf+8cEmznLggfD0+JbQ+fdBDEoYHXgk0UIAhXQVhhPuzZ+1H8gxPJeNd6jZxZLZNniEXCSyEVsA
nSJQjt5ZlVXovJYPghdUHUyprePB+pOJ3m4fxztv+mxA5KA9YuTTeG3zArGnqW1gpZsmtHtz5il6
9aBpHPDFFa34VItkf0OWOgL7DFITl90p2RM5F5QxwSFceqG724JqCzZ0pf29deMTbpU485qFDsCZ
U3D5lh41OPdm1lik/teczp0rP2GRQQwE8kCCSRVWgRvszvonzIW5Cuypwe+7hSvL8/Ty6jWX5Zi2
Dc+R6COybrNI3dsh1q04xgWm8GgKCQsHwy0/Fwrly7Fvdk5riBp8+DeTt765GbpblS6zjraykXm6
ic+4F2YUpKRloI249WcdM7Po+YzdauIwJqhRdUDh6dyTVFj/ERtCNAtpWsFRx06dmdbRk3kCf/mW
FuxEPI+4t5OEj1RjwVVdnimkNpJ0LlUBMuwizhP2nlYmRs6EJyQ371dtp5ocwfL115Utw3j45O+R
xg9+5NNWCRGhwSN35wWV0mLLz5nDMrGQWwQG96+DjqmGHafXA6IXyCo7e4RUornFGeMd0H6+NqGy
yCRo0Ecw1+NrredDwPTF6r26Vkwi1ig2Z1NK9IRfQnH39HdThQ/ABed2g5vbxXHlbtXnVrxeZT1t
DiVaPaPnE91da8HzQoEWGUywBnENY2aykOU87onnQitcqNAHYkiL2ZStMWVBJKJWXnw9ZLUwLOA9
0RZciauLhsOWM+fI0REs1qeOYBGHIGoSpl8fhxXBpWqJE+BMadLEWaogosE0jhMEl4o/ANjI3gAg
mt6r5oAYGwTEx2EzeFwJTMIIGgcjv0vJUgSGbN3bFEDKYk6DyzGKDwbHxHtDnV8B1z9GXrmkbXcF
ufb6iEY3/s0Gkp6KSgsPzm7xMD2DMdCZKiJZ21U1s73qlmV2Mg6l/EQaWlrsh9FvDn4BLNbnj/Ha
s1i2OD6hv0Zk9rWl5YzQd1to/geKAC8KvklHXZIoWJBupD+X0i+FZuQxJv61ZGCfeLUDepujcQeu
KT/A1iKApRH6YjjzSgk6DCuryYajOADisQjsYYu5eMOaxlQmvU1s5zDsYk8+gnfAT35YdoK3Iebp
9I7HSZAlxXOoiv6Jh3EKjrcwRuhqxWj+5gP6NMSvqFIQe7+IojZYRfdlooAfZkR0OFDQ5Ga9V7Ux
6XfyHLdT6WVhC17YIlsTUfHbEIs+3grmOrRHmKclJnY94uMs2nkNQSQlPqAuABf+HjkwYEqFIkF6
kyMn+ZxwGOwumnkQvoG1jZkvJzWcaqHPju0p6mNhROYszwPsxo6GWTeQFw/hkNWRt62WE7eoQyWq
48g7S709Wf2G7qROYQInUGBjQpod+hHwSWyUp2XKnkUO97k60Tpk03gam6nrucdvUy6r6Y3QVby0
BZhBDJoUy5uYZ1W7befhjr/zuKvLfXsQjvr4BMKznrPaTCGZfiTSRDdX0n2UcjnFHVt+xwvaJsYB
gWLGpUMjET2JqXqdoYRloW/EY/QF116W2KVl+7Ne2yLgQOgYuoDqzgHkFR92Gx1cu72wX5UTAIfe
rBPWD6zwaPDrb49f3ZpzxRqrqg6wA8rrE9henid1P70C1y81sSjMuSwdqr/6bI+P3eVTxwYRhaNm
V7L0QxSW3zT+2ni3WquzVAREQvCH4yzHhWRquhFaKS0mzwomGN47PPoodlshPyYVfPuIO+SCY29s
6nsUGxPxvjJs9F/kp9FKxdjkQgUN4z6XxLJHxgRz45JGoA2u1yhSIIEhdcgj3CAGpZYQm1jiVqCq
3bAzxSfTi5wi5QLhgE4WMGoro9ZqvgifC+34l8qifckWzaCFu0TJifZYFXeznPXDdO5Vx9cA9hFZ
sJhyIrwTAiZoCSTyaDs/FaZAn8mR7kWoBKOLeWBzYtSGhSjctmHfmf7mL68kwKCtf/dUcoKj7QfH
jIQyiOi6NrtuhUiIbJKzR37zI726mE277QMrQEHk6wU7tWLEvDczWo7DuwmpPmbZTu93wvJBx49U
+pveh2jdkMxqRLrFWEgQLAmQoEkadupmuIQtbSbQtg8KnAvliaCd6h9fCzFwXJQ0wgBSE48ZYqnV
t7beWovdiU177Qj7LpkhCWOrFkiJGAmzpeXQjtnoAR6Ho1XAFk1mQ2BvApMO9fHgWLMKAdA47WtW
zLZm8PC++UdvHMd0tVCdzwIjlOefLnlpxNtLLCB3a0vxyV8b795mAoxjf6UQEhNgq2djAB8Vdh4O
9VCYh3h0CHODsyyWBlql/+YttriJzFafbY8Tf0b8qWjnTlU0dUkrDvl6+5YiXUcd9nU/yVijjcD3
6RfyKlEdEHeXqEQyPhrGCGXnQKBMeRiQ/uyxV5oaqUQG9ci585NKRNb94biBqt2jQVxVRe6XG9bq
89KDrFuLsm/ZuVhJ4PQbq80wkp7DOGhgRlwymB5g2z34eyG9HZBCDbMe1S7LuX+9ysb53CskkesS
J05H8hn8bl/T7o8f9Ipl3U+E2ELghGlzVl+f+F3jcfjQX8/yc/0kJMQyRrMhYbxEhT2b1KpFSL1A
+tmhVtK2a/m90gzynbz6XgiXFEjHgnWJhjHGCPC8fEKp1TJTMCCjvp3fZzbbN6z7/nW+r6m8PwNB
Ab6tHoXnk2WzCZnjexfKPj1FHCOEBFH6La5r9Bhz6NcM6tPuOOtNTUKemIqqKQxtRSYmaYmII1v2
pdF3vIUxtECpooutpnP1VzRHjtmXLZ0NEnY72Lk3TwCAEaGqCfNh5LZTRCuW10A86c/rGIURDioW
UlZWXdpCkHY8O/l4cvaO9G8u7EFHcz50uBejyyjH/8NsDgI48PAxvpAo8ozVjSz4xDmqkbbzHJcW
X/T3SFyHUG7YUvwKn/uDdBQNvgZ6rjks70+aejgY2vjDK0xSYFS3HMkjRUpnkWK682X1B34a30YC
/GZdLn81T5IIBDjDW5fTdZFc0esdwb8ZNhO6nnz1L5FtjOpbfAKXB0zwc8EQrseJnawAxIrnmj7j
IaQ95FLKzN0+z1CSKRTzLgi8UBfKz8XKQ1hUyDsSrBX6AsHo0NBY5Q7B3vl/rh5YSVEhCIkyUR7j
HzzOn6f5+ctD23CYsWMPJ0FWYji6N5H2euy26wlbNUnj595sPJvTzxi9OaRUBWwGmNsyeHzotQjN
lIBtKOhTKDojAaTAq2+uXZxLpzppFNNIY1T8lG6WT74p6AukNlKSUIAcGDxB3KDfUyIXZGNbdlc0
yN9TOUFqY6rWlqusDSYmZsRoToqhjWN4Y8PuS17YIhi+X7InsQPWMG+OVoa9JI+BfPc/8HhUYmnm
lCcwvTTs+Z6chdpM5f2CPYWn+pXBPDC6OG2EKhWiYcbLMzEjZhyAU99vs2/YHF/mU4u3EMPDnLmI
6L6R/ZC/eeqGscB59jnlAnKy/IaIBv+XEfLuCXn16ci8kKOtAjugEqB3sM4wPxoLBQHwHJDrUZm/
u5bO3tPBg812l6CpGMVA4eyTyan0fD64l7j6lhwWmrxlASb3Mx37t4TI53XnbdHHWL9SGnaGP+41
v8zhysyw55Bs8RX/DG2BpPvTowbmgex40I+uSZBnrl+G1VJMWyctiXLdLHSPkq6u2+FBu+jVIEeV
1dMsqIfDMDZLQr7lwfo6AHGGpNOnxNxIJKDAjaIhN4GDzxZ9jicykG1Td/fa9ADylHdvAlyb1vVF
k86JDIPcwadjPLTdBT0wB7ycA/iN13onriYahHZqrMmIbj3wtzOK5rYA075soJizfztRdRADZk8k
m8AoffC3yKkUTReO6BmWZaQGYBxVxbiaqAhGAgyKCo2k2Bt2Ac+1+b9ap1D2eu9hGF+7oY8NfBr8
Kzrbm18M83IxOYb31ScpPd4c2LHIoDPcQqO2Os1Q8PkyBarP6f5g0i0D/7zdsLIGhsClMT6JHOuB
ubb22oiD7rZLT4xhb4f+41ysucL4h0YDZvPKAshuRpltfNXZyKdQD23HKIB6IK4z4GOO0CQoLJ9I
Un3QKEi2iFB9ofpJqTiQsSUjbN9rpyO7eeJdmPNK24LKtC+UQKeur5caoUYAoGnbvtKj5QTdPlEU
JGOTZhgVnW9DZ70Bje/G+Vmc/iVy3ISKTuCntEcApYJ3VpWnGvTt6VWsJyn0j1CorQ0YNYA0JsGM
VksEvRzZ6daqPqFRdWlJBQQ06TZObeU8hgvwzXbBVV1IwaTz2RE+rxAREop9L8CF+GHPAgwcvJRO
1nggy3ckI639w/yV+OYeniHbHQgV4JyRmhnKNNaSrDziOsvPqFg7pKLgYjw/LBwPghEgaFFJSRY2
t/OXPkV4G8q7rdvsFLNwlmTvjYKqMpK9FeznkrtEvYMCjWF9/j/0ys9tzZMKv7SkeyepcovYrVGl
2NhRyPjwklERcUx6nRPrwfQ+7UP2rv0Hh76NnyBPa09H5fh8D0DI7EUW26b+nQplFvHTUYDQ0rVN
EIDFcUMsokeCxjs1mhwJDuAUNLgTFaSFJaBzyTkY1v5EoKnVxp1E4oMP2Ycam3E0vaeEKVy8Nm6F
qD3R33Q/DpzdztMoQQcrkNpiUvinLwexqRTlBeCUq7pPmq6UM91+/CDmUJ2f74Dil4Roc96Sc2Ji
I854QoA/xz8fC72MiRhNIpMuRaYB9ZtmI4PtJn5cwbkt84wyWYBatnyHktnH0n0KJn9p7frdYnh9
Kk9tRC+zUXegpP0ZFNSwIW060xVX3tnTbmVn744ZBNvVTy1/lRCcLJDPVSLt6oekCc6bVG3+MT1r
lGSOk3Vmm4N5AqDlQ6R6MtBYsyoxSMmY3N2UQDFL2Sqz8hKWYvSZ4Ud6fvGSdy6hUKAV0ezk3VHZ
16OTu7zbF7WIdJxkznEfoMlPun6UwKVCNgNv380V2EUKJSTeiOnvXN79NMglnXbCzJ1WLyM34HPY
jKcD1rsCql7OdDF61ILBDMGRS1q37B38g6PpofIMMtqQeC08dEGGAAK2J+LJXPvzexsQWZjejmNC
nvSbxsb6X7t+HjIDTANVxUxuW1HiiMe3fIiqp1j4mSLeGEoFUHcl8LtrAXYGugWbRhP0d/26St/j
CFdJ3VDmjXa/jcWDQF4ya1bkycaTukKkcfwpwZ9mk/wtv0YokgqPr/fGca4Bv0+gXBv/+1TTeyec
5ipOzBw2CbrdbgGVzJczYGROg7zGXbHmukTk4fqWCAgBWXqi5rcDaDTf35b8p/LKdEo63iH345l9
KrPRfVwnxXZe0MBeQL7McXW+qdmjsm5XoIW/jCPTUtUFxUpczZeu1gdVWxK6WJ3WL6mlIvlovigq
WjV36oo/YgqIU4CZSQtaTarGybs1sjQZmnpelDkHif6fD8++I4C9Ta2V+BhPPPaf9tFcp2B+Q75r
pDFnx0yuIFoZ+LeDEUqFo/M+IPHRQT8aLawrcCVB1OvLnZKucfM7p3hZrnWnozPDV4ph9BsiHz5r
QMd4gOoL3IxDwSZAFeJtCA9XmolEyV4YTlvloxwiZjUT550fTqgI5y7/LXu3SqHaE491LOrZTWp1
Gy76nsOX/kOsB4q7BhdOsWmjdqww54BStg+uI7d40C3+N/6mgDu9sOeHwlIELak1/7Qx/f/wqdCi
s1kdFtkJS4Cczf58weXKci8W9m4WDfPeAaI0zlJ7asvN42Myaif56JIc1yQGgX2BYRIdSqPdLIvY
38wVpnW41NthJzEI9DMAKn9xWItRvnunwsn6UNoGFnxdX19MUBQpZ1dVJjaoJ2pB6RCpqCJpqAA9
8TZeYnGnihW7hxrg16RZvdYIWw7ywzBBY+RhSvdfLl2vqOlePElwxDQb/w1zbUgbjo81nt1y7mS1
1EptQfSse5EkNdc4nAjebT6t2zij4/WO5Ug0sKwZnnqiacXDpGK3ojy67N1QoNR0crybmUM3Uks5
9MdSSAHoUz3OFOOnkrj6NHJCjo4Jiap7VV9g33JX9l/CYpzq3F1xsGupyv+IiU4KidR02GXPMep5
hJIZVOWooZQGIj0yhNT9wcxHoj8ccoHffDXgT2xiJLkSDVJwwAXNNJVvRGMTrgYGd12GRHlG6Fpk
vSYSouA0tAjp0+jbpCpoiuRFWaWuuHkaTVlBixHf5VO9j9JnNZPk6I3kxBZWHurxomtdfRgRFHf8
Zyj+mTubXz5G8wou6npZ7DkBUsnNXxDM7ZimfjJnsHfDhkQZv70kFpB1P3pABg9BZIagXdCIZGcI
AI4xGrKrLxIHyacYgsE7reIYBY1Qq4IkdzNsWE78IrNLL2Gb6KUXAEAvd79wWvDUDCPJLBLDMIg9
VG4+EpHP/+hGz7BaNhHwi+sQ2rSO+XGmh7hiTITe8/NHCH2cz0Nti8ynGJwFF6kYe2doGbYUQ/on
mK3Ab+X8IibfpFVMI6gPFnRcswtutL4nTYEORkXi4skwJ8AlA2jf79XekO/+H8pkwHvt0Ryo1QMp
n4opBSL4S0RzO6QA1EurnvAjUIcOzlRmQomjWcTwk59dq9gjGPUgEx0SyxH0nJOlOWYrzQca0tz+
dimgUR3is5lSGaZggVJurGkk3HBvM28S1N7dJalXsUsHaRzdc7HlSyGvvt0VYS6rFa1gaKA6s/Fd
QRR0GmHdPHxpAVA1oEU5OmhYARmDdHMEli0TnlAfzKOJqNfWWtarmSKC6/Q+2PHzwK8C6HM3i8/k
ZfStBMO3nRu8IrxM+rkO2XfMvwrgpVMr3RIDAD/kAKsE4ug7ECvpbsk3zf6/2MAc4yS/enN2xWg2
cQxs5bINlkyTpP4d7KAU7qY5Bnoo97aVbEQs8B0e4xzG5RmtRp/aEBkG5UTOO86Z+95NBSp6bAmh
Wqk/j3R41AWp1EfyDW9sDuQ7Dq8QBKMSPFNhEVaz68U6/1zc43WVV9Vwp+0mGCSH3CzfnhJkFKT4
mklGc5MKe+VB0DJiq06WQnGX/OJbbukf8Mz341NiGOH/3pfB3XQOfYdzG0KO0UWASQivOCWcqnun
RP0mXrqXWr/5XBoFqq1VKONFP5/ZQO3SKzh8LE26GluQbaPXsxUkE91TWQ7Ptl/xQCvtDd1eL3Fb
cxcEuY8pdwf/wY8bs/BBhtsTD5YKHVpf5zsUsC/xJbhtqX7v+kTZO79WbF565b+y2PM9c4b2AW1/
NBA6A9hV5eglc6GbDGAwCY/3l+YDbe0lOjFpILK6v7H2Llzh4Ki0ivZCrSkn7JeR8V875bEJrbyy
A4NUz+taQcsCUzYAeSkXnID1MlYxQKu/lHuifWqRGQYM8BOyNz3nfiyMuHsNRpsoEODYQMCUYkYP
4X215rIG4MrObD0P/a/7BF8Zv3lzuWzNB9Lj1sWuE6nxSS0yQkP2c5O82MNcMcN/mBKZLleIPxS3
mwqKi/YI/FoA/0rbkwMEj1PzceIuvzaJjh18+jwjugeYNmWNL8KPUT/myylJzqFi2ysVryUVfBVW
Iev9R67+zjOelBqy2guWIEhfwxhIwADS/5tdZhEAmr56i6vKvPpOMmGnlCmmCmdGKjQ/jDBHk6C1
6tapT6eqsEscP7qo6NsdgeQr4Hlg7mY7S15vA5GRjDt31bfreqBurqlCmEf4oreYPvt5BtUjAHDS
wRyNDsIUYJcaCdG9p/+fVz2AbxraabfhUfVqEq5qLtbSGQ6Kunf771rk2oKb0mfCwsE6BNO8Zb8r
QqZoHPIgu0PRE4N/hk/HWMLPcJ5fDGB32tQkEb0cNVvSOs4ELqGl8vdwYqM8NDimBnNqZ/o4/ZGh
cPfAdqFVfsdJDevaicNX2AeztYFQqb/JAaIeSCVakvkGvY+Fs0IqLc6ZLrEmxhITvh3jhTz7ngkh
jqWTrVJ8bMfj+vw4V5NeGSuOznGZ3otbjQwfYhKolBxBA8RiDoPr6HcgoG9w1okfSVrdWDbng+xg
R1Owb0oLJiQU+K6vnDtfC+aJe/6EqQJS+ghV1V4ezBDQrFnEW01W3UxbufDO7m3NfdmM6pTeRBCe
2rV6QedV4k+zYY/PAY1UwieBe6QhaQ+tZOgMgkxXMsJ7UTJjQ+E9+tuAWxTAhuu1la2IesA65BgG
ZckjZ9DARd+QlxNO1TcqLsELc63XTyxzwr5QSq2GRcwA/wf0iWD41lDFs06wOK67voTJde+n9u6h
vm4Py301n0wyOUGZEcbqIkDBwSrvof0F0itC5CLKrezbisye4kGyX+YBEnZbIfcn5LZ2qBD2ITaC
OMOwKXSVjiUtJrUHCOm6qld/WOKW4kSns9nB/PksB5O4b+qn73XBRkyeTTxsePo8mYW0Z0fHvwZw
fmltyyesK0glSLl6P2gr58y9yOc8DvY6I4iJmajZDzfKeYyQ19tvPHJ8Dw+apvYz6uflsQi2JJzz
PLRCtvEyfdV2Tr9SA7gEWhyIe5lEKu88/tT3xKX0eeIyD+0Ow0WAuCj6poTGXHCPrMQgRa+rC9Wn
3fLUaXS0J46LQTMAoutmDKb2tpcbH2S8WYChJLRwIM3Scqk/HI4q+PI7vKaSvzeQCf85Bf9/ittj
zJuYlBs0BvZmWd77mC2BJBpgHBZw1JJYPcSL1Rb6WCGhuYmFeESz5wrcq/hL4qkr9Z/99lLECbxr
K7hvZi3flyV/YWSZ6JUVAPtX9JK2pqhgrYnjTDSRzcU8HN/3XiazsrpZIHeCtv35lNgkAPF3+ZXy
5kovf/6ifgdMzAiRtIqe2i7TJNlD3lMGbkd/Jrr5YIsmIa4G9Itys8qcrMJ6oKhWpCpfu/IJWMCN
mz7HETd8kBMNeEpWnXkj8drrOTWEqFxuitw44Mxhi+zQBt4TkMZoluu2mdyLs8N5E60zueUIJtAH
haZdLJIuY1MP6+IEakav6zBcNjuMnuO6JEFeIVhTuHuX35w2zEmguud0dUT0MYXHop4iAYBo+XL3
OhgsKa0LtvG34RHz1KaBnOhdjAYgNwxAQJ544PJm6PfJAW7Jw/5/DzYNUvv3O5Uh9W3y2ax6D+OE
CwrExg6WOQxIwyl0nrIsmu1JET3Jl5LljFHOQbn/rhGiTc+wa0VhAYHyGAe6TjneLpYj4TYJz6x6
FCUWx4dkUGFzJ1ulDhVJvlW8RvRVX86s+LfBcQx9j2/7srF+om/FRvET/MgnkPS4mjs92Xsxg/Vx
rpnB+JCHUJwEs0zmcVqKPKgeIiHOVUdANaJe4aODHgvVu6fTHgGAKy78L3hRoOWLq5s7nIL4cZ0I
JJKpTSi3F4hW36VPXlgn+8nMy2qt5Rooy9c8jV8vZ/o0NZHnzpP+e1ty3PyYq9KEzdvMz+ikuS5Y
55NQMNE9zh8fzmImkXg+WCvrlfJHFQPlkJQA6T2HPkl1Pl8tlLuOJS3maO/udfoqztERey2NV1/3
s0mL157kHWhgOG6ZNhUjposQvaKbOHQjms3E9S0TAi3oUKAbN+FdHJQDPOwzdxemh+OrroPMcmqt
69LAakM2yHMrhhvEDXzIKbmgI8mVvBJXH8JxYVEiAH9UXjF0zXeQEUI0aQZmf0a6pm4zw3Zo4z7U
HO3w1zdJ4njYcmt7TC3zte/rilXtDiMUZJu3Hm0CzrpGJ9s0T3+7fyLOvtNivISIGOybH+sDdXBC
yV0jqmJuly55R3x6KeC1Ha33J0SyITEuuz7HicIhG+SzgUCEaLy+Z2/puJmjFbL6fVu1TFdRbjyi
nkMVEwXwkXSYW44V6b6f72nyY/MGOj6hqWcfGBtNNwmmwGhuSWxUFD+FLdgAs7gDq8um6JU9OypH
JNtMLuHdJZ3nINuoWJ/CAxqD3DiL5eTk9S0fPHN3xzyE4FuD4R3Y5ClX+OciXwMPKf7oJYAux2jr
7Phao4v4HfEhauBqZzsrFLKWsA5GVu97HU6qAW1rA6NUh0S1LFLDxuiEmYb4n1sXR3JWQgofEP5Q
vA/Ab/2nFlozmA2XZ07qeLewPF00dda/Ih5S7UWAtbtI8QxkcODN1s9D6+1cAJGDtibECX0SpXE1
IrfNWmx2COpUtjbrbM4iMbdtZTeQfdbIqG9VXE8YsUSGz14Vi1aDUMA7ts5X/DTgyeetFzECHA4I
CCUsv+RnMIJwBLzrYyD62VPkdt6YUOUoynmuneOyxpcEDXStIyQ7my/Rj+oyJ2yfP5DtS9RAUW0Y
lYQUa5PcfQbylki6RmUSPj4mZtioH9tq20uBWWBmBAe7dGqnFjXOzvYJZMYSlRF0lgmIHqSqnsNa
NYEyQU2KUKXxdp+7ObwXpSUa0zD5g9XMEKilEJRvD8SX6IjOUkEQToeLPeOCpOXhj9qRx75jw322
v69mgueokd9FA3skB630nOe5UWvBZ9f6glrTSLQf1HnihO0uxnaMtyIDXOibHToUkvAjVrQmxmzC
wUg0J5obBK9N+GhT9y3cXF+kIIZv4JTjNk5K3eXNeBGm7gNN5Kt1ZA6xzXN5v0cXy8EbDyOkurjS
km2gfOdi7gd+Q6WzaAfOqAlxH9ffHNJnnLaClfkzDPnTOxJt2UmW9pAdYHC4CNacfXhYC7p4T7T1
6cEK1xNs9ELPVoVgGjNAG27ef1R1bEUfl3YqWSNTUWKu//iSQ2m+h2vtK6JlaAumtySA4TndedaL
HLw2u/qQY3pLNqsmPf1Edl/fRsFuVYu6scDMj6mgU2eXjyeWrxVA3crTpBeixFXmdQHD4ZbgW/7y
jDlvKp85qvN00hr9SJsdirRB9uBIeTkRPXFF9+KVEYRjzyT703Klxz81nhUbbhpoQvTfQ28RTHb1
FAzc3N1X9QyT4m0TuXWS/vvd5CpVINPk+aDLu12k76Ep78hIwuBEovxVVfSdvCtqeW9TY7Jm2IfX
uYV3O4C83AYXgfHKKlMZivIp1PN8wejmhFD0U9OnzeaZBp4HP+pbS8NucAUbfvVsE/VjxxSrVdE8
odSkLwB8v/bxYvdRHxi9bbDXyvu4EeF1v6GCNWtvhy7Bba5kgVXOHGNf4VuwXeRjkhHA+OdG1u9w
ZwenXcPkAqH4ODaRn6exMooWbLgCnkVbLC+bmk+/rKNsrLddLNoW/5AvbzoNinYTIcWDICtC+nXv
uKEmTHdsECBIUTUxm9+tMM0CCLQg2BYDPFUQX2IZxMyz/GbY7RZS1+5DPgMve33qRG7Idcu49jQU
vDKE2bjKjlCkU6oSH7VS35p4xcWtI8ejdjxEL5p1N9gJvBImrObaKLp9bNND1IX2zA2haqfz1NQ8
YpfmtfsjamkAGLdE163/+X9cIjkQPWzWJmHqqmoORMMXzHJazGXPDbAxzfKGP00ztMRK/CIcF/K3
Nb2NE3u5v1TlhYtz/DMVOLJ2j942JpIBYvOUt7BHKfzVGM71xZgvhsABGBwRRmm0kicTAeOmmmTH
lDVtd1vdP0Fl4WHZjXANsOtwbavms6UTx+IOh3JEYO6JAHkqbtCoO91Ftrc2PELON7j33p5Y2M3N
iv6nC2UdsxCRjZLkzPsFEuZp0mDpWxdwwKtUWNvnAY23mx0i972DQq1ks1FG7YDRfRgyQQhXAh42
nyVYeO727NqcwdyodFApIfZesX3peUtdTQIMsGPu6+VzzO7Uto12JjyoyGv0Ry6io5vF4OHt81XP
aXOLWpbmnUZ+e4lGNcsgd6SXHMoNUm0ZsHWVGCeqccS++95nv0JsCdpaZVBfRakoprH+qHe2SMnG
aJ+rC9dU44wbtMYt7wrkaSLur5vCEWvfh8G4XHF//FSdo/sEDCAbSqKHPdMzjt7OCz1031Gz72yD
GtTRxWhqbVeqMAmmCMVwmdtsqjVeyYnTNL3t8hH/GVwrijoD+f0LFUgFL8zN48/H+eqnP87hNiq4
PzsIXIH2+2HyIIX33b8TnkMU9RQuLG4pZTjokT6hMIXHIndvn8/9wu6pOIipSls+OVjCRe+4LLH3
r94EpNEahvVz+P5tsx/rvENWUakJ7shygG2sYsIYi8qtIi6RZ8NeExLZDUhx5f1rxS7xilOkQI9R
ZpvnbcasEr+CV6L66Mf8GvMd+xCc3VcXnRQcjSfNTjzNHyvgEx2R5gWorI4qTFPfx6xQaootEL9x
1sH4rJw3VzXIb87f3mA3ftmLyVT8NktYRpJ4DPOahvJlfHTUWHapDMiO3q0g8RmLu8ICNGkINhut
lDEkX8N/T1KMNcrsr/7Fcyu5nmoHBeEs5gdeSAtqjwNEKbS7lCx1NY7tJJ8UM3FW7Jj8X9LKtCnB
IBza9qTzm3/kyNTpi4pFMFYCQcrdRgFYyfkZHK6ivDJpVFtx3nHL6TKDnm6oi7cWc1rFBWrBkM7D
aWRvqkLfZklssUjVueMVwRA+ccI6OV21rqvpCnqGcVDgMLUFaP+2ToYvZsjUP+v2yZdJ6ubncEI+
H1ariu3OY93gOwb7sDevmckxXN3V2wl6JMjnutr7ibUP8S7Bloo7fJs/R9UWgcZISYb5txEXzx47
sdjnYzd6JMoRXOb3voZzXXDWzZYrOp6F2snGAnT0hw8xqDWrEmCsvvi+JYV1/dNBPhPs95rD6PcX
qKSJzdYnXeXozlsYQBFIebLYl5dOZum7RosT1PW6zKV6nnR2US5T14byoMNyT6nl+SYAnDWEDW9p
Hi72dtw3CzpX0ROVufcOlWl4QYfIyQqMO5akRXlGtzRbHFBxBw96Urfnw9p5T/Ppwni50U/oNxeY
Ou4I94p29U/YZstMEmUZMP/39w5XmnFC1t+WOqhGJY4OgBl0UKEQVduu5j5xh+IaXBLKgspQSGB+
KOnBPbFV0a8zjK6IlQx6qmatzHLanDpeiaSVAjdV7R477HdaQkIG1/LrWoEk3MUqjA8mbhXa81or
xsGbXI4W2OdC+3xbbXMh7VD1hQ12VWNjeI8vt26C9eg+cVZvQjYRY043Q6LCPI35hO5/ZsbBndD0
ixKXIVCFb+y8otxQWdTEgvUYSD7TbYJmiVakbxc+wA6wsreDApxXFoGKsHRXNFZswnwwfSEsw1Gf
WyqLcyzOMOgdct0SBFrvQwM2YsPJmmRhP6gWxSNwdOmIjyQs17ydgCpRP4uMykRYXX5S6976PitZ
TMCXnY5kfPnlRdjmeP/g/pKTS99BhCZNbydDYdG+dgymLHk10+EnDng+Fta2teVXXz2YQvQ5FO1o
kzgZbOKGCHThABgaiCp/dUwQBN6vXAAdK1O0RqoJm92/9HtptHA4FDW5WcvXhYEw+FfJED4/Khs1
CureyjdQGj4nsWTmB11W9xuWlRGZpDAn3rLd39mllN3t6lSqlL8G22Vatp0AcpAVopYR4B8jA3+K
f+Ev6CuaO9jqlFhjlVpA26fU5Qg/PJZSSmYti+7OXQ6PCky9dqefJ7yaSabdNLCC6ClA3tq2acQc
A7JeZATOixl6dqPEoAkgCTUuqM/ITXr1YN6opb6b1XTIMo8Vp6VbSiLaBh6SBwP3W/iAKae9f3YN
uC9Ti0/9mpVjPdueW+bByN9yYWSHKjjWp/rBY88Gy20PwlB8mTTSZ4uujDtNz7Z5VHudN0T+CcyD
+/cOQJW6waJplkM9R3c4GxN9v7ujYddwx5526p6vKcpoU2ft5D1ySVSeCOzvT+0WplHQaKUSoh70
CAeuK2ct4R3Xku4u87E2RftrH9oWH0RDSPyBr4eXzuUrT1z9UHdM1PcnQ/QhN8Fnm/kRhpx7Bars
rsxLWEJwCOjIo/81adBLu446BPAOuoqBwN4RKR0KJ++PFLijnxuTozToxrkLGX/ZW3yOU89tzgOf
y1rLn6PC1W83YA7Xm+SjMJ63REOj54tgGxw5sAcPEwRevsD3EHC46Q+GI+YCXer4n+RdcZa9JWgS
H1fZ+4Cg3P25rgdtOZrGsAVyTURBK1dKbLOD7ysAmTldYJsn4AYl9q2MDi2Q2POAO7YTKQTXS5VV
vB3XWO3gk70V+6PLaQBv+H70d54BZMpfN8XK0q8rAGcxOHmi2ii9TVAuzKE0yFbkGAbGATBNxfHI
hOxyTYhaSYHygRSzVUgh7N/q6Yj6pcridt7YEse7GmBEgChQRKDNcZHaLn8sBstJABaKPFlHjA81
Y85NoWlXOk7YzPyK/WIuh8lmOM6jQowzrJDsG2GzZ2aUwXbtXnVHqVcLuE+xgthFIrYD2tdFXxv0
bcxg0lMfJ+bH90/q9ysq479GbaHZ663WwRvfEWPhlDs4MZwGPj1sK1QLBQDOrfg8US/MAI0VH/Py
7m3qVt7fSnW/2+Px6Ypf3jmlRQbISipuIXpn6RcXDFTGXHW07pGQGXZrlTohu/Ge5z6eSsrM+Epf
/m82CYv2CF/aMPT84kxBp177bFCxolBwNCa5eZLuGXEc7mGSPHZPZZvc+z8I+o80stYx+t/KpZsh
+iScO3seMSCcyFyzoY6xghKscFi1yazpZ9rk/ZOQjN3I0Y4fwfL35/qzvjMrtK6i5Tb5v7mBpbYZ
6LXK1aL9ZusFuB+R30nvp+2E8cNxOihXhhZi33p5sKkVJj1YgokHGre7Wr1rVTfQokBT94IZJQit
5ZTOvQg7zE1FUjt04nL057a58JIpKUeDZoUn+LGekSE1RyJZT/VokKlrKr8BKrfXoj3TsSm2O/w9
f3JfnUpbdsp8bJKRAbqSahK1bOIMN8eDdxQlgWvXKonlWaxRXPDOfK/xonhdPfJCwb5rJ9aQJ+q+
tOUhPbrzINbWVLvkLH+zKiRisccxdyEPasTUPqxpBUQFmXraOvQURn4kwOoUTnscRpYQgWsTrVE4
+Zy+qYvse84iYg7B3uMCpRy1YefaOSPqZbOmk8UNDYxi4NSzVxEnKCteF6kwcVdaEQMNl2J+2fSi
qxNxB/xx5UuSilV6bPgtYE/GXsJkO1+UQ7EmwWL6C22cdqECDeK/Qox+NuXd4DOu0imQuQ6iAZuR
2Ekh6AdzHw4IaruYQEjHJfHVwhoiDeJMMLd8lfuxa3Y2tTPcYXckrSfFrDvO6gIexUsgy95e/Mvg
egKEKSyM3S1mp3mkVJv4wkZyhjeckkS26qZrHiZCPMbuq3Qs1kYUOV2wVD7UewNzYEnXfiLaJOTo
b+5lWLExj0ojpUr68VLQOp24rArdAEzPJxTcLAbP4TSh1zSJntYG1mBblX/vdwpcxrYHIZD8E1lW
6IPWuKI6Kv1dNGiO5wqpYEcbw3dFBkmUCKX5ALOQywWjOKK1DbN3AiSnpVoe7Ximk2d6zDaWAuVc
32Tix1J7Nhyy1RqAnQ1OzjEScbDJoQ25coLy0QFSb/yw+L8EwNcWmE5E9cD1n1diqWtQRf4cvHuL
TH+kI7G6l5JnTZHt0Knvpk7Z63ZEUvPJGwlvcbWTWdnzAsB+8DNKSicZmgQSu3why9oyabqCW4HS
2Bi8oqXM2gQUe/Jl1OBWP5TQ1hH//44of/iNijhtypeZDGIsCAV7tMYAy10+t28U/UZJoP8D0URN
73qSRCP6QaLTQVdra/0GPbYK67JK6Ucak7fVkmwgWcgqksDJKqostXine+2NknnL5PKsBVo4RhJa
Q7PfUo9WF1iHBWz1Bl12fFpgXT44Yz5CiS6mzhMyfSYJL+EZrs/tM15d7PXdoMdTgUXvuk/+EejP
vkCZbWdIMcJk2H/S+4fPDqrhaQXQCR/xw/szUfug5FhH9QqQEcKDiGPgTWYyVhYbhkoT/SEdi96K
Hg9JEZYWjk6k8zl2EI89dtO9vdEEdCLMsOIMi4LsP2E/dvXVjbdOez8nDol7AXgKppDhJTgE5U0M
xY76QRm4wLw4BbqPgcEk4bEKzvuUqJ2jL4G4NiY8Sa+yu1IXB56H5sgwi5aQHHKF2o0z4XOtrruk
Np49vvTH2hxTBCDDi26UZZRLlzOa3nywmn/Z26mI54jmrC0Ejs31ftA6vVMrORhoq4/DdJxjDfBI
ZwxkvoAt/Xp0p7rLYIlTgCjjKcjFrBPEMnEsFQ058FWDUUcWY/zgD+goAeqNArt7z3JcZMZ1uLN0
+Gf1mgVHJlUDepErAAhyl6nl0GJwiEWD8f+wrSLeh0MFdAWmf5ynnTQqkTAAMJ6o+8t6c/l+WBb2
z9YVTNYKNogb1C+9gOfOQDivWS1T3agnfp2DkWaat999Lb5fYSf9RcY6ek3peA/aya+uCFVHXryf
mufzIOoy/2GAzSbWdc8MfU27chpjPihWEcG7iVFAgqKw8WzyyRURcQ5Xv/6QtXSDt0umkBKot/Of
abnwXps2LcpHBCWTCOCuLMJGnWpza/gsbBDrHjy0XlUe8ocuWaRtYdmwcklP3aZ7KQsroM+ECUmP
htKPOYjUiLnxpGSlF2/zgE2WucqSh7IkfOzgrUbJrU40m20ykxdbMuExyHC1giubcbyIf6O3jBIr
+TCOtXqd7qZEW8exa2IhHwK6kIpJpfkXqvj7qVB6CYyya6sbtdmWXhxApjm2279Ls9POArqefR/f
FST2IAkj4GUX/VDE6xWAMnzQnRw2GbhnL+80KqLGqcWNDChHpxjUU71daE1YTJq0zT+Kb8s1tiBa
DoUmXo+iYt8N9ip9DiomU1hBeOHIrjv2lTnXqwl47igkn0gjRsPY02L+iHcp8U6bxRqp3cEWSdGl
3ottJc9d2Rk23NuQ4Ma3XE1537DOImnLt0cnSWEh6LdbA3u5LJNT6D/MaV9zgnLWu9RDehRLZ//2
zZwcqdEbwCb8x85K+Tv/wkuVyNQ44hMUjQhqOusH87+cMlFbpjvnbgL6AC3JW0iE8jpqJLDTuiwu
NavJ9r7n3fr3BJlEF8X52yl+9QWwqw98p9IahBgqfhzyFWdrT6I5Al7d0Uxi0bq+Flkp/xiAs9RH
e6XvpjrgiqJFHAZFwIrjvs+NPcsHvepodSSYNp4TahhSxiY2Y40lkW5jSicKHLPFSinjstc0dE2L
ZVNN6AJlE6aPG9rBl2SOyy33Jx5MfwVON5PEz4xsu0hGrPS+si6n8+DsQIqglulS2BBupOmP9pdX
LzuMU0WkgY4xGab53EntPgv1nU+WBvAxLCoXKQx52WGQ12zdn+HuFuUMnwsf7ZuAiiehz+J2G4Xq
BL/OsGMDTXQtJnLYL702FsiXWAMo6l8zHIvN3zxUbwJ2oNGtpNkcvOi9iEYD0iApzzLpcZetSZn9
224SREoOyYIpEvTDNq3JQQKsmz8BHEf9U2n2w7CvPIydQ7Hn0KbD47Qcv+qZJsQQcykiXAOjfY1c
hgLkWrha60mCDic0CaJrBNrus+nq+hgURY4MwSHpjii5eZI16o/OebX8oT3jk/Q19z+xarWEUBO3
ywxxsrCm0lhT4jNRu18PsBT89y62C6tlFvlp00V7ozn8ZhHb3m1vIgNmPHVf5eV6kq7wth1K3X9E
G9KE7pkrW9BL483StqBkdJ4Nfh5tEjarJLKAPnO544D+N/sYz4y0gX+JrW7czucF9JK6x/DncxUg
6DinwbwH/4WD/xeN5Zmau72A1dv6MRgw92jm1+4v2j5LSdt63OH48sq+8j5bj7CNA0WC6nR5Btvb
Yf+Fi4xNpfuh7XUCJ9jqUhcWkuxhOh4kypDfHqvodSLF21kwOV9MkLaVaYPACILx5cG/JQqNN1td
DDGDQJ0bLIV3U866MIBmk6mykroA5f9kkl0qMv/apo0VwZdr1MSIIyxbHOnOb5oNANofwAirnXxO
4qC3jExHsl+apwfEOyg+1HdZsKV5FfQGxgMNZeg8jHr8kvZ95M4OpvQyAnHk9K4eJ6Cv8EMb3vaG
S54UCRYR2oexwKQbZS/wU0PGgNUI7IMhFWk3EYaWFjUmcXU4dCjSzqKPP3OH+Gk3q77FqQfGeTGo
2yKILpeTZeR42ZHMRhpZnrKVHZo8f5ZPng+MYDQ2DkKKTENqPf4C7YCwDPxO7H1R07g6EV1e6lY/
7JZCK5/9IG0crqfYGc3Rl5w6UC1tUjjJtKTCX1fUxf5Rt0tsKReeXrHUTRT+qcU4xUM1VSfliYYq
x3b/PIA46+8gmgfaJhsvN+SvbWZybT6Nd+4vg4bJHxn441qmbrobH5dfK/pRlj54uU00uz7z017W
MrlqwDk9azyFb6+jsPLxRUPUkhDI8sBqZlWsDl3KXB+sNmEUHWnIPyb82Tx4XOm7/kf28q4GQy9B
z3Cb/Frvjw2UY/rJIj0NMmAxwChGbTG4OhK+z7APYXkU/QRprU4fIUaiDDOYfquBEgOPowIOp091
SVLKOSU9HCRSzntxO1o1Lz5x3Qu7tVA9545IdrCysCpYq0afKA5BkKHT3wl9r8qH/Gc49Yl7SFDe
ERBzPzPfobwcUFyi/cbdJTi1RkhuquBV4GLstvwvwdGgD5XUXkHZhouw7VvKHOnnr9RriDJPkj0L
hm+m5GIniR8JGLas8ebXoK4F+ahLTIZ2STTN1ZGAt+8UkUy6ympgOevz5IuQPsRPs5od73BetBrQ
DRzy6sl9uIxrMc+0slEhncJOZZ+GS2mO7kQ8b2QVrUof2J3OQJRkNzMcS/f5/XQSoJUmJ6f0821f
WXicfZZwB1P81azbzVOVmfN1itnvXUWkC9gc4Q624QfSmVOdCMfIDgnhWCP6qxE/XyTacI7Fai2L
B2NlP80QeOrhPMWmGwzgVmA4QcQxZoligsdvM3iG+Pxtn0O1iuIctx1CYwLg9zquT75KbbUOWTNv
KZwXyWTJxzRSrlXjBaW/tHHlEdgXRKgeE9Re4WUKjNNcxMYuiwUO4V3jB8Ba7yOhS1o2IuKNTn5C
ZKAnCKwgd6iDDpHVBUWyqZt5DHq6dabazHCGrQoqyZ0XuSHemzJvBON75Dh5n3YT2KdfvZs+C6O1
y9tfNAmf755Oezz/oR41eNPPH7V8rC9YbwJ7qiF0V9gkY7x5eem2rSPcs4qO7xlCl0oQgLj3W8ga
Mo0q8grq8yezTbx3SQPtJruJ/7Mkv2H88eywz+txWezWZht6yd0kq0Y/F6sXm1K1i2mTaYBt7jeh
tBzcAqdMT2drsV/+tuv7EfvpWl+Lr2rc+Nj6Ghp2MzQiFcc/nvvQsEwraO1NlvrDIzZ7QUvb7F8+
wkuoNVPyQy94ulCmm9242osPE7zDNXxG5bDTYzb2Jo+NISldN7t07YcxB16osnFGv/T2RSS9D1P+
SRzoB6dr9oQb9IhMvmeNpyjfKRUlso0vHCv0Mvh8XhyozIq5vddB4Arhc8nH8yC80DfJRoYb+QqU
y/qg7xNmBZ2Majd0eYRnQASdHUN0B6devSbFcl6+8hQT9PmGEKP5f+Gh7wo5R8c8kr1ZlGw1V+k0
dG0vWdnU+MhHIZV4o73DiOvHIkwAMbLFDXtZ3QytN2qaCzI9vDnIOtqgnlgUmMo/4NK5u+25AsiD
kD6aLuwL6I0UU4F7cCFXq+PXiYrduB2PBGxjSeSW/HBGMJ820K08M4f56bwndC8K0YiOAec6DLWR
t/v2uqlqcIdVzQQxsBXl8SMljXBBNfma4ICKO8TdsAoiHUcojxXEnT9vCa9dOfIsH6XAijMz8/BG
grfrtC7q3xOshg0zEu/7nlEdwZPwgNLOA9Lt3cAv3O4+Ns7aFS7U9ZtIq2terYyuhPcxosADRdvI
h9Fj+hcEq9ylzCo+J0ZEYGu8dJjwRiSqOrOSgoTxv8oy7HO0O94BP/nlhtlnTM2AtTDox1fX6IaS
CpgVQMwbFZlEMvnj7J6Y8bh3zMVLe//3gCzMH/yUmV4/V9HqMiH4lVEZCNXYZ77sgbYGdJc2d7mK
0ZRUk/foNX9gp1bV9RDqS3UsP3t5LbJjbnFUpf8IeCs37NkrnKjtDP+ESm9G4IuMgbn8b3E8llmI
VZt/UGowZJono2JrunPdIRFObkCAltXTt7hcpqdZO+akSJouWpMvb21u4nSwkKhR8LVvlBEgRSlg
sroYC0cuERXZ4l0QmjFvl8OcTq4vgFb+U+FCF9GCrCJtPoslRyDoUISbt/dLJ8Mwq6mQ5kKdoye8
v3WXIB7DgHABtZzmvme7otcl+NCITORhn+QnECklAjx2lfjBg10+oSpyYAnBOnLeUWluT1C83gOF
w1x6wUgnLmC9V46924mHrTEhR69TbF+9yNF+tv5nkgoGqJCSOwtmD3PO25zcuDNcNlDAvEcPYrpK
VTI1FgjcSA8uXdceiUOirWw5AtPa5Ko5q02aSAvHlfCWwU3MZ7zQ+HFDWci1KC2LHeyU/jsU8lc9
qGR0X+iptu3Ld1X9PVjg6hAvcBs7FHnaylemg5fK5TfHTIPBAn6Nq+X6WiPHz2IVd1vkrPKnuxx/
d52WWatBNmRGhjsOW9zwtSBozKKbEDEdAqFeM1MJad9zkjLOPZ5qFsQgDoem1IiClRAbn6pME3D0
vk3W77MdtaYXs1LlZ+uDsuLok/QcdvdAnYUr9ktIqry0xtm3u780KGI4O2H84vZGkXJHQJD9EPIO
yrawzzsUfhQ8Cuditw4t3N/mHrt8V/dnMrgJdetiTM5AJrwzYCgLvx2uiBUDi4r7ZkxYXEgv58vh
nwBk+NpP7fsYjLZ61mGY5EGjBnm8oG5qP4P3sHMr6st+D8HgClwjfzUcZJAI6rRKt4ylcFx1HGFe
u1K0RaDU+dcqXrE2yK+3Lcib4eTpCfxc7ixgRktlCDcN1zAxNLbgiMfD3AbYEgEsakKKAK5HrcWN
urt6bvxqBA0+9QFRr4EOflJAz7U4Ivrxpzrgz6qCXbzDplQkydcWQxn/8IXB4YncsP3RrRHUZmO3
hMRiOjck0KJna6geAQbE5jDyxUyPM33stbcC/YyZdHnoXMiQHH1He08v7cb6CSoBHfhWVYK3/rSe
T9QdB7zcefpxyKvc+hLMokm1zFZLNb+mEOyovzZtLR31Kkj4ijU+MupbMqB/m6/Tshh0x/VTIJzW
fIKI17UHRYnIP3fQhxzNlHWKWUxaflZ/2+oZSsvY95g3Ysf1GoOMHwJTieMBSXwjcljaBwG7Vipb
4Pk5Rmlu3oDbt0wROMsEmgKEOGDyb4FW8yABdOQAhbPN5F1B9k6m1rXAQ1ncWVePwcyWSKRSYg2R
YxUNHhxfKRlEuIKbU/yFKn0ij1tK8oKJRBaeWYiRKebbxFB2G+9oADZVmwsmuG2P7f/fRLDwHvhs
ztO9SZJKiI9yCiQr+HZ7xux6WWeEl04U0OP2HBkGlsEerIzva3E4yGQfOa0V3vjTdZoJevlVchSG
smG9hGTENkQnLIBhSw+ZbF9kML1TMZ+xOdxL/uhEgREDxc+kRGlozoPVSYTUKrL7lLAVz7h3yU/z
rI3fWJKpCD8eldf84od/CKp26JS/CQixNr3aJyI9VUZHYBJkTE90+lYEDTnu66MfgFpgM3JaRQRj
ba89A1BhDtDHA67bap1bK5LAKMPN56h0XpWb8FJ8JrEOBuI5q/iOxeaRueSDv1m/fK4JVNGUzh5x
2SQ6ptSoohv8A/dGBS2jHm3IdA2JR7tKeFqRe7myYGG2UOQmWBun0wdBvG7vOYz6itgrSgaIuKfj
d9dbI1n/T+ivbpI9eckU5tzyvglMaBrfPOyqkdlPDrJe5tvEz4idppfUMoGkMPMzOlPhkOGWaxUT
yNL1eJH4I5C9EJLtFV+qIlDtFcTKIJ3Yjnjuy2mcKv6E2Zcq1r1mcDQGWghp/wEBsX0BKbbom9pu
3bgTDZpO/R5nAlhu1R00wJQBDHHIpFict4O0KL3o+owtaQ0w5KfhmW3B9mW/mCHh3hewekWwvua8
k4WGqLnYs9RUnf0uZTd0q0JkvAvHC/29zAom3t1oTQN8kH5ctvAnKY9WTUVtjoeg82aq8Apdnpdm
H2l+bXS4U7krf+cgLutFh3U/zFyVcg4aBKtxjn9jRJZha0G9dSeWEC6aK001H7C6ZdfmBGW/F1nK
3fInVVJIEuBKECJYZzvsMvCZWVO1k1o3oaEF2y36YBV+VQBdHjx8z3qBY36PbbZloXdIyWJX4i/E
JPriauSo46fSK4epz/H3GXosXtucxwD28pTg/Za9Dj4vy4hrMGH/R392toeIfvkOXv9jIjzkxmBz
RK52fn5PMFtu9ZvrPmNamQRiPz3GNaAkxydKgSL647nUsIALFiZkBBuXm4nxAixnv/t/3dYwB+H3
Cmx/NQL470TDGSDARRUutYANan7+Zw0EugMMT2DrDk+WXsb0XXIWyNb23jX/2+SkzsV8d6TCahuS
ysWDqOwpwd55hPPHW4xP5NCHDsoqorI6Rw2USoX5DD8kB+UYtznXhscBSKeLjNRvXDxt67J8R55e
m519Wx/WvGhS1+4A9xPSpGYh3uwQ/2NgGr919K8jnYpkEB3EB37fib6K97PDdpa3oa+cayinXpOH
OjYnAgB5n0LOk6w241CLXqZJaLu/jTzy36dov0mqbVZc5+Dc1TUfQXxs+w4SbXIA4W76fylln/dP
fZ+arEkk00aeI2KQleMipbxB4bvywG/wSVopZJYKi7xh0/VC65o05b+ps8bVdPaN/8QnedFAe/je
fYtVlpj7r6miRRtLO1mDF7uDwJesKqrNBYQXok7kcyuHmg8nOFqkoJdcdBaxmqAiE8c54OUq8Phs
/oXIThhtJxjqGSIpkyTFLnZhgPWTWxPZMyhQNMgO1UKkb45UvhKm3InfTha0nxRtMoY+55emp+ZO
4DHeye1Z/xnAK3j1FffsZdAZr7SUv3qBsUO/oz43WmoVmAKrPbrkdABhxVKawHy/glCwy3EczorW
wrZp+i4D5ehu+4HRpnARWvTejjcANX1BQ5w49yLdPEbT6r0h91QPhwSWrabudkWZlrlCQf+3l8Ya
G7vsbGO4yypYN6wgOr8AgfF/uzAQoMciaSftFBwuiYFzgq1zsX/WHZ+sz81zYn6mKSVks1xq/UtM
dP4kX3RWqI39NNiqlNB/CQkRd6cSN1sspUC+5ifIYdis1aQPvL38EKU0stNunDK/AzXqVyiJ7I86
Z+0ShuHANov5waU6uaNdg66Q5DK5lq+zNI0gbgGcgKBlmsuPCjrSnTG7rS2K9KyaLx01O9qEoY4u
GeMoYOoKCCebwcGwg2uJJmSeaHiINlTJfhmNSRwgt2C+iJe20QvaUo4vW2rIIVwWkJ5JHx1gEq2/
iVGTX8E4A83WXgxFXOxGt1rgtw4cY31+OFRm0uDG9Ggnnq9gyWNyKE8g/Gc7JZhJ2nBWrhreT3uF
cXZevrDjxd+1auxYh3OZJzguE8YmVA8+QLGRmgsEsofmRvbyBZxlSnzKkiRG1EUhOJkl+rmdOXzF
nwfH1f5bLnQV6FGj9/rbVAs5oyyagxx1B4n5zOjQFO5ZMkOcne+jXJw3UMK8yrdSDIz5tbT5uakq
UYDP89U9bI5oauNXROoMuuDOC3qyakiu5GHc5ks0BViqk27Zh7bjEDSqBFR1FJEydsF7x3/oe6jv
Zoa3/LWrjog0RRVhfelYIZ7o7eKBipvYsc1XRSyGifzGirRe49yuAMHQTp0OMDcrK31Lc545lESm
RYf2lEHiujaQR+LH8ubT86sk0AcnO/ckFRWEG+oxwhAe/qfZiuSFUAzsRssysnu8g6ftmJ5Q1QHQ
B0XQouXNOIA1SfTSSuROdF4FwJgCbsIh0q1MtHSKK9m+Fp5j5gsD0f9rpAwTBGFSAFMjPnw+TuhD
DP2QY497bbHpCljCqdUQm1eNnPxN1LoKd8bPf7+nS0OKyLm7hF599PXC4YkYPGLf7GIUOVXpw+8h
KC0hbeLI9NTdA/pCq/kKgn7FpWV8IAyGEXbCM2ZY4HrjQC3V9i6sZMLZ6WQQqs1B4CciZQjvHUzO
264sPHSqMWwaq9cGnrYzIhPrk2fgJ89zjqrx2mTVLFxIJr+LYTTWGtabaW8lm5r3DkIMoOpZIUly
We0rOMtCCZOqe2vEq+Ead+J704UzKFGga1i/3DAFdLyOQa1FlhaTeLdwxMGrtbBwWyqNlyGw1mVm
nBfFcDILntQaI+GPSGwiKkntpXoSMVwI043AET2sSmZFbRDxAaiedhet4Kkb7eTEXFWAzj66mBgH
StcOlO9+ynL2zzxGnZIjGHsDaeNNyq8g2ww7OsPUpwxbYHLfp8wUkrhyeX2Vnn0ZhcCaJBBsQFJg
+C/mSeAAnc5Fq34ayou0fz5pqInO0OmRH4bbi9x1qqYc8ajr6PXttjXqD8s6Bwa/xFqsb5Awx6rN
uui1F2xVL9Cf5AlkW6po9ytYnkUY3C5tBu8KwMi6j1kjLo6avvUvy1sK+eDh++HemnrWbl/LS2HH
05AwcSTuOoAjl58pYWk/GG6Lib5xZCAB0PcHlBXA7pSn+0xTy1m+TkminxNPL4Nz9y4Yz8SwZyi2
DC/F/shbhbeoPvH3rLWOxeX34YNkwymbGViLARZOiMzD8eOmYJYi9t9p5/bFg6xrIIGYx8maUli2
3SqCfT4p8NcMaItHPFRHeH/JKFLUzF8c2KEUlKOBLtr3A2HbkrHLn6RmCDuKOBV+wSCOBTXHVDuH
OJ2SpkGno4kgwIJ63SEkjd7X/lukPKUhhWNgtd49pFwVKGgAJS2FkfCMcXRfViEWJIJV2Uo/hOYD
9xpcwZNEpe/L5s/wHKElA6q03d43KRMXoV8KZL036xfpOUl6O4TgAhbRwQ/52DeIXR7ljhnoqxz0
MIjEpCnPTjJCoEy9jebDfhM/1chtqNUaGnVj7chXmbDfxONjPCJ/zOEEcZ0lDeShpJ10MF5XjOV1
08weWX5p9RtmFpDHGTTzcFR+zjv9qxGileOwmrNpIMfDNHleTQVz+V/8/OU2HnsQcpKkLc6aPHqQ
lrc93d6zXFO/vKIx7RnSazs4fXLCCYclX0ILLdGur2LVddLASatLHMd+sMoM4SGTqEPYJibNn1K2
zp9re9W8WS3s4SPBvLkPzACU2JKQwKFrwFT5zlDuzpg6K15XKmqO2CrMkJ57e3+t2Lo2jLMvKP6a
mAbx3So6JkxEjrOf3t7sfLeGoo94EZNzyKZzyrs+hryKOZHfJncCSM45e8e005M1bLwcIbSXJ1Gg
OgFQ3AW1o7D7PfXq4yRn0RgEoXT26+XKTsH0KOYjHmQXC4XnWvzNWr63kPeW1hW39lHbJMvVQYTT
KeypVquSCfTAZd5HE/H2Vw1vCVh52e4+/65kQmNKae3xAGbKqLxKdBn9kwjZRJZb15PGHpb1fwlc
1YR18BL6XKBrDdLkArSOFJ+dxEW8+pcNV5/NAkj6hHFleKUt3PRYUFgDcTSWWzNIUNJzJKTGwBPj
RU8Eb4G9W11E74lJN91A/B0HFKhrvEv/NGpYM77d+QEYCDN4OqqiKl+GorNmt8dEGx9WJJUQaNlS
G3hfEFVELtmK0ABAU8YxgqX1Q5PbLClTXwaFnEE6B7ORi2SJIIe1EXTaIBgPzh/sbZcqqoRAeogT
8kk631ZQ0IrPVpqNRFld3ZqNNXzpu4jxyvcGrK34SpXRPwbM29eIIk+iBb8Xt51B1Jms9jKJZS6H
BlNx7G4TKt2+iDz/Fo+2NWO6WZz441VSwLV1iAmLZxw1FV9/NG2COr8Jx7is+yfhc1ARXLdSDaUw
urSft9JLd84HfXHGmJr3SNbndHRgSouwBBx5NGUTOz14ZGc0VCy1kq4cJ1SexW3i3G+9W3mC0TSJ
cfEimKNEkLSyGop4U4sXp1A/8Tbs1P3wJRXeFw+a3WQlF5Y4PashLmJFKk5OGOMUKgJlb3uKVSb7
m6vO3nUuOeK8V9gYknFisVZIcOqcgPOa958v1L+pW1XLn6g2SF8g5hzLJ6kaVIZMuaZ2o8dyHVOV
HocO5X2Ci+yG4jpJukUZrO3gK6E8kNrbvpAQWVe9Nt1Ckmv2lj40/8GUqr7fyEDg8CyeNQRLRUcn
7QBX/b68ufuo4fwZU0jJ3YU9v99IJ3TQd9RwfzH9VKEo2c6ixnCYQCraejKFDElqKxOojEeI5chV
P0XuoE90sMghHEt5Mehv+2W5r0vrTrBihHidZxsfaiDU7axJM/pgFSudV6xdgGVZBUfA0euSq4md
JYxJq+7BuHtUWyNsDIc4gWi9Fj29KU0HYwPfhDeyn0MjOTRGFLj9hmtuh/eFslPGmvpK9qdTN/DO
FJh6WvLeLarSqwbnjc2KAF7rfzsIY04WTXnbT2Gd8tWoixTWgu4tVebOwxZES4AHFPyKfKdGtIzk
N2QBCc0aqX5NlRy0O6EEG4nnPUA8u7J0xGnTqUVe1xcHwiqi3kbsquvs4QRyZI6XWto2XD+Djbf3
+X8ImygxrQK0wNazlpMRRfmSr5fvZoMPh3dX1zJe++hpekUZRYEQtCl0HU6NdXwtK7rBY3LZq/PA
cbLSJV8kGAgNVefz8zKaY1Mpyu29NptiBZL04GuG6ADkww6C4eNvoOLtxsfQXGKiILzcMhcjWf7w
mOlwYFYH49qnHF97LTn+zZkkUOp/acdmlDvjyB97s6scnxGN+BHZPmThO+nxBn8+fahVCvVcNGA0
Wh20Wp9Y+0jweE6xmAcV3NxIaLGEWIUKq0Iut2n/acLKj8CyuWFYFGp+X//Vyr0c64dIWPUXrk3T
5Lrkte2ljdIoDKwrh2W83XfzdTN6bbsgoSZCcpQOBkcNkO86nd2qFMGl24rpysfYDevfDtxXckNP
dWWzeYHHNSqbyq4D3cf+YIEV8jFpYXFOCeKVYyC7wd7MKzikCfkqD4dRIjcwlSv/nDY7hxyJT3jn
EtqHHuuCybTM0pyybbl2HQQf2zLBISuRP5GZynNRj3JxH5yp4255bAlZmSpTQ0F2TDKyqrjNAbIe
ufJUEwTkJwe55yl+OY1vA2181NJuS1r6OJrP3vBUPqGurI/aMUd5UQfNRON5pzsVwcXyVASiBI86
QOhGdGGqV3daamMCRyJ0y3HOOz2RO/upzXuZJnCqubawJCh3d9pqh6qIv/VTjcbQR+81twRau5FL
AmwzTmHvC3mkWtJ0UUrtjDnSm0fpPMaxekrTof3ZYDIMkvEAtYPjectvWX6yG+28Dj9CDgXhgkKr
lVxAlivoQR6FPG7mU3e6fGl6Cg1Yx2hpC0snUfQICmPi1LnJFxrIF00y8YopmXYGKvQLh52suHD8
pxSk85sAJ6jotesHy/TPOamKg8e3+M72NNr1cGIB/2fEbrxRFmHXw9HIZ/Pul1SW0FYLSa5hm49R
9w1aSnRzcF6jd8AtNsoMtc1U8dx4y1tEDP0cYSmBkCIR9QCY08zoqQwCD7hoT8vdEUxQ6tMSNVm9
x/G3NP+ZJNUEgetAcFNbf9p1vR8xpkofcI9+y/dUqKNeGF+N54dLHxPvfDs/Hupg4mc70MJupr4H
8wsqIygeJcOgIKhw/zJlnvSf2GQGEAUk7knE6upUnc/1l+fiIraSusrhvvh2zxiom3Q9p6ApTmI5
YuxOca1fs6SuFEPqEwZHFo9vl2HP4DFW3hak2ZHHZYbkVT6hl0kKWcvpgzbmXLF3IsjBx4ZWhSk2
NXMxRc2qS8+6aM3mR3CdICp4EogB39E7nBH0SvejUuduiF3k4PW/n2G/kPxmw34Jz2W6ryBdM4Rr
NgyxfIi+b66purniMcEsPZxON9U9MEIynxajZzjJdUcwo8d/C1Enpt4orsnnytvTvmkhgadP14LX
gCtlfvtIEx8xDYykxWV87OzawPqXx68zg2bqIN/RYPeZ14lP3N8yGSLswUndjzSRY1eCFvj9EIPL
1RWJFVPhOuNlaHQnNzVlbY8z0Ht1kopw7cAMFIoQnWv8r4oN8a44ARA2OhBbFCcB+6k/h3zI1T4b
3+S3GJ3XemTWz3vTUv7PdLkrDgJUJdHMSTDF2XQV/h71GjiA1n/44FC5GabVlDuapecKWWOVzpUg
vTRC6pwW2YfRG46rHjSmMLT6zRswQABMNKuTVTZdB6zjeRfhTaiZ2N0SF+9P2Njmfyt45QZnBLfE
480IhMwliDG65Evesde72naf8D4CXOr75Qa3HYujtGv9hXvMFWi0hecubxuiwdO+/pGRLPJqZGtY
hJk3MJiSIw85PjoguBdgSMTOdAwRSoEdYy1gyiBnwjqN6M/J7yYoxHXxQU9ZcrqOujG0O/ePNLQ/
K7lIi7WWZvxkacGzUE/BAU/qImbgjjs3KYub6uI1r9UJEp7nGIFkx8KXwkhlbaEAT47zjOqi7djE
2++Kc/M+p5qYpaaWgBnFycuvfUEpEMMcdq/hHk5Uu9xEzhbashSC521Wj0ZbhaPANnk9PKWRE20r
b0VI80T/KgM/MSrCvQNqI6RpQr6bKUMyR/MjPXenJFDMMAHhYPcdHK81B4H/VvMcjCl1C6iuL0lj
TZNjhht5shF+ZBktujbbzYgEsYGZF36PLIZsf67Mr9Ri3VeghoYeNPMbMjFCNLGB0QIglFJMZkVE
8DekGkPJDLsL1Eft9HS2pIkrBjOOR4GHUINhI/32JaM+WetGBH7Wr8Vc2w6a0lbvJ8Z0vg2w/8XB
B7X7GBiuWyYijAnx+cBJ5Z2JZNFhIgSNsn/CXaJqT59YWV+yiG8tS5MkjEY9saMae1doethIPjc3
WECj/QSR60TvHlerFF70FbSVGVOSj6qSdF4NrKBYqYo8kaGs+HHjgOUZl3I0ThbKCoNEgewxgY9y
yIz06kMejx5v4BnuoM/nYTdC/YEmW6SulkVPWgG9wy7/WYP0s9VmVwfzjVcsAE+ouDIeRATFy7HJ
SUeGHMdpftTaQyK4BBC9e1EQ7OZdatrgcCsHkSn1t3y+Fb5sd9FEWVTCLwW4iLE31DX7LjA3DF7s
OAr64kZ7v2NvTmD3NdYyHjpqBDj2F+lIt8fEl8vIrsFNp8hxTEIkG4XGn+fVa8Z5AY0rnoSLmrQl
i1GfG1ts7SECrLMdmBcTBqRGXqCe2A/nrf0Uvvf9SPYWOm5QTv9U8u78LPsY9j9C/Y0tpGZeJ+nV
q2seQDDuTTsd98lxLZDpbctuTZj3137aW1v6pQGy0dkwJ9lF+gzHLGeuszMJ3FMKsTTN4kiGWdut
/IG6x8G6dFgPO8gyDzHBpHrVlTVdUU2P0Mi0gjSeNShD9Gc7Z9eSipcnbSc1w20Zw3fkX7/2JOuX
2VcmrqEgxVYyJKoZwWLFy7x2HlZey9MbuMFZkAvLhkDNbimctQAMQLb5zkAWQmpEXdvkI5FUaU41
LhxYh0P/JSLzn1wulVY4ob0fQxaPirxkCwxd1dJ3l2RUpfaQow9Ef+PurOFXQjexk0stbzbzOmfB
A8uSas66fD5IDYQKtdZVl5b5l0w5WYF26xCHab76HLM7PXbSbQkuM5cV18RNrJD0YQJG6Kh2/EsV
+/yRUW+KUZWfQQnKqvpEwLue4yG3PAo/BINhJZxMH2T+aneiSLjL0g4NyZP68bUpSo641ksJVLfX
tqAyR1txDgXQjT7erTn4IJ9Kl03Kwi9n1GPJv2hLEgP6k2ezJspgUK5YmOe0MWghDnF3Y+CicrX9
lyJ3c+Jd6CZeXfILK4xw/bO312mqJbnmFfSuW4Cp9fricg5aj/2k2T77P+gSXL/j9mBOfa8x55wZ
nFQ9V3G2tPk1GrZQ7P9xXQMZ6JJ3fTTxvajsua+i5vlnfycaYflT1moU4PMDvWrZ7SSd7G6oXzqI
2Hlk4BFUDTRF5bcL4R3CcBLYpLxY/2E3oFY5ceNbNw630661g+5neF9zBPeASRZ5LipUbA9heBGr
UMjxRaQTPm/OJC4paC5gXwcvmnPgrAytkYkhCbdXg2PEAlUJg8yCe67rKQezYnikSAyD/Xyjurcq
teYv3MWtH2AqcOdZNcuYl6klDJ7dAvPAcO2Dy6t0Yjd6WoDNir0fBPt4Mq1c9+UKijDa9JDJH/QY
0ORz+JDEtm7INOqD3HH2NFjNLChPlQugYINvq9Ea2KKAujMkjDJVBxboxhJFjRt85LUMQhUBCA9T
JWXM8XS23vUMKA8MoYYbBqKDTCMUOOjwSYXJ6F6pg9kbvnH6cNjldQV2lI7HUCgHXMdV4hHdbLmA
5I0LeFsX4GWOGnirz9Fs8YEz/I3fQ332+3OwwwX5cvF5leRtAKiecSuBZXjm9YrifwUwlZndtBjQ
44X0tjSCC8XVX7yY9nfQKxTx0IQs1ALU8s7J9Vu3r+fe5Bqjapg1vYU4Cp8n7e9kgpBEkCZTZahu
bu+WsdxTobeY2qphWeLUmnxPlj00SqMkOXZC+J6MxnmP9FltwhYnQ/tf023/Og5FhVw09zda++NE
21PhSCTu0MPWE3a3ORJrFL2/Ynidj32N+9YmQ/BnlJiGlBiEsOh/Z2FlDRyku6Knrank1PIJodih
AFzs05LqomlcqEVsPuf1VlHwE0osSC566fy3U7+3JhNPzlAHs9bjh+XrP7ONCW7aZxtuEB1ZrWiy
PcOUDg17kaitfJKLt4IJQxWDY3aRKWc9x7mrbLdej5f4YxkA137eGo4paUiF7fdPEuu9+LWpsRj+
j0beIAxZ8cyWkGyEJhDNlr8PV/OWUJq5nSpjkUsMb9U7GKzHzL/TSmuJBdxTTZM9cYQ/jXGgrae0
i7JpCZBbxbxAAR1wDEJpaVwJSzkIzIe/7RQYER+j60hkwx4F5wZT2fbRf2SFeKPdtn5kGr8MdVEi
0XYr1ASrVWyYJNUEfgWE3dKcqWoEHLYutblzzTGpDp4QimuxqZCZWO8p4umb+ABC1NBhr3CLXHPo
VF3XLy86rzRG0w8bhtXDpZnPYkh+CAvSuLfpUaNl27XIV+BhCYpVIFHa9GO6OXv6DP89lsmI/aGS
IqdlYxwIMgPS78Z03irqR5UU/urkRZy67GG0xpAF1WOA0Z8s4wlg9848Un0BThSGI6J6c+g2cmx2
4AscG2gPlKWcjPMYSSD8mvqARMh4/Zi9VbEAnAU56jwVUyQlkCchdg0rwqh8aEqAl5MzBgXbfl9c
JbWJhyWl01RsBDO11NMp/xQglqujPxkQPCaTbNKVkHG1kwpX1o7BtL4CI6fds6kF7TVQ3co2iumd
5MwOyqKHzGJIqG6PKRl8hadagd9xCXhGjLWugo/jBIe+ik6AiQDxTmSeNhH/oI/m902YRCPpApOJ
xV9fjcV6layzgSxjrBrzUOzHxbYpwA75noIKCuET0BLCvEArQtaN2Ww+rv3hbjzTOyhPgtvyTuzV
IZXGJoC4vjKt8JPxGz2jgrPR67d2irW/QHKUdq3Fnf1yR3Gb+nQbndezQyv7KGEet5iv1xOpmueC
sfPZiEraDA/zB6ljpa3acZk6H6gmwVTWlteToLCCvo1ITFMUiz6MgHW7IXiRFYJ56bHfV85irbTo
lzQqmtgeFy92qsFQKecykbt+Baa5zMGrG8yIPxK6YF43XpfuSUw11AekBHAb2XyH1oc0Di2jILZQ
FvBYmX5T2TnpNFGq9tjvrXfjse9q33eAO/eUr3lh2Yraj5dM61101UKYA4xvuli5KQffr2Wuq0Tl
57vUV0qmI1mKXVS3lz/WfMTwGRW0zE89q16O9QrxHLNA8QuQKmjZRMtfL/yvgPKf3wMsXneChbUm
0gGkuhj8bU/RjAs3prCR+VxBmjutyH77v/xZpy3b/EmDa3VbB5Dbb7KwAGpXkZnAOoNGk4R5nMvW
/3+f79SztLsXgnXpeD9trIfT7zSJwk38VgtpM4LpoI9B4y4FjQTd6QhBC0cFonFINE7pwoPsPxeH
Ozoz0M3zYfpqeh99SGzFZOvww1W6E3Pq3IGgNJp0mKnbeJRm+23ZmFMyLk8X1PBsbDNrFlqqh5zT
al1hh+0oyyoXkrYOeGH+UczTmWw1UTDboWGzmsXBEzyybeYR1ZbpXOWBifdu3QHTSTFFPBBe+wae
nGrr4Mxpttp9dYPVa7Vfa9Ajor1UBzYoHDMqVHpS9i+Cclg1ZdVTegG72fuuPdfPENpGqcLlDPRJ
73g0EEVUW+48+zvWSrWAqwiweszPcMfkoBFV/ddWVWP7icpDyevjdORjZq2SW12hWx5TIHfLYkzM
tQnLAjqzpZteagi9l26jTIb+355oTlafkUxOWuoKpZQLtN9nD0mfrX9zeumIjXwa5xTldWiaKUUA
zUNBcf7FI3bj2VRea8EL/N23mfe/pye+BbwtAzRayx77ULVhonRX9tYarMWT9CKHrcY/xf27IYHc
xliqwxGqal68LS3oe4aErDh26EiFGwdfPvtUyTtoJpCaPV+5FcbgnaggjkQsv05YyDvTrm5XSlbD
hcN3g6P7RSklQTt0/WilHE4dPk4kocB6VKtdKU9jLdfki66M8e+8bwVxj9tuB75e2E7Lhgu8waT/
hmqWL3feUMa5S0u34b4R7oVVJZiZlSGGFIRNA0PKg9H9q9HqWW/PAUo4WJDDdmwGZZSUqjuB0e98
nHUdJKS3UouJc/OZ0m2ARS5I5qW3y1IJot4aOBXJ/5kkNXlptyw6K1G2gCoMIU/YieT9ZKwP0qbu
yKITZgKVdEtMelbNyMYEYxVkA5bfWlHSbF6oZBzfoicQHel3zGS717T45rFzwucChASGDBC3AAkb
TXHWh/61EfbgRCQq2Qdz/kuLtcleubxCrPRZMCyHeJQRXMMyMfkXkifBqgIZBVL9Vrp3VHIBP6Ya
p+XZKw5t3oreFhfMLxWQ2frHVB02mHuNoSInAuV1+N37jP91v5zD8Nu8d3FZtIa/rHetqJs7dJYZ
cDlQyGkpo6osgssZXAPjc+yD+tcBLM4xwJZXZGIWoyBYcMtvgZPA17H9ECeNCqHJALeNs5MbifNB
M37EUlShHwl5RmK5GYbmwGvHquaFSGZKwrfGOIiA8jUj7WAY77KZTtGo4WESGQ0Pds2ovcf8u0BB
iOa+3+mKLCJP7hSjITp5gE0rhHHMINpyGrL2nP0pRbrvy40G9qsHaG2G9IfmwU+DJBBAw19PuKf7
IhB2oxmyz3FzaYg9jknCz3IU+6T8w7QnGtSilnt14y2H3Vv+q+hPiylt6fjKQCTLF14JGIAJC2Ag
aeBbelNKn5iROh/Znbp1bAuQ41liaPAo67Ny+dqP8ORHcI9uP/vzUsxcqIP2SHZY9g6RvQi8TUqQ
3urROcsoIwny+4FCcSHWfJCJLvWo39FGj3DxEV31f8rDjgxveqSs7fl8TTQXazFHGwbHAgyu52UT
xqXf3Mtqfo7nHKqaIx5JUCZ94Xl1S6L0kD9Zd4NOpsxn63TQlib7cHSklnhOwNAb/DAvwS4xxQiP
00R8DRvpAnKfBZVGOQ+HX/nR/zz6NMvLmV3JKSnIoo1hDLHXgwJUTLh+DpD4xoNxq0a/AzBLzu2I
tZNMV+4N6FCPAkfM8fcmV95FU4PmOtSA0O97GtVXMDxD7cAssuXZ/JC9gguOtnfXPHWkdDwC1pnv
zzjU5ud8979IsS22j9iOwKFCXobQTHgtKO+ATQbbzJleRk5BRlAWbi4QNfIwqv19tb3D0TIHw1+C
+SZwCbIqEY52qcQUfJYmKe+epcI7pyENV5EoYPsxiPWBcNMIlf4q6nVcvLeJGATCEGCPFN4QuEC5
mr/F07COw4HQmM7IHqH0L2sDCHnx1QgWbHbvSPA4AoEZ6v73+mFeiqSKDBMXUvkVg1G3n7lAda4P
qdGEhMi3kLmw7B0bsiJlGKk4LkItZWtX5ibhy3gTvjJoCznk5ktt1kUfn5+eY/qL3fM1bBwBgwzB
TeWD+2P7GlICnrsbvpOaTI2QNVP95DaBoxndJu/iZZznasfFMexDejQZPyRHoBVUca7nWC2iHUXe
WH0Sd3Csyk7oxubYghJI5hDgWTvTf1e1Fo+UTiSajiSgbX3hygTTK5TtW4x8fXEMFQ/imtdjdpXI
tevb6QssDtHOcSvFRMoWf098FpoYzAP2TqklRuwB/2NpeNbdmf386R34wfdGQC3Ifua8xAw1tsFs
lBJturmqlmYE0HqkSICGv4uPZhnr9FgCeMQNBhRycgyF5csA35yc1tL/8hLUwZIo2KirwSv0TMWG
5848zD0D+f1kEGq+OlNR4Zzg8k/tInSL8yYTNGbvdQcfnLpasKpQS9s2H7k+wMSCFVxaVpECxiNF
JuD2UmO1J3GrGvgSQTsQCJo25fpLT6yMRnpNBDW1aJwSv8F8p4dlbxejXSCDhU61gCudrcV58tdW
sMOCha1j3+hmLqfiWbxPgwdW+Grr1FtpRhcQSJyhddvSBpSs/4iPcR+Quzq1TLL7MutpmZh0vS18
OY56tIYOtnDKn2rOUE/BtQcDBXAq2aaJyMuBlEyO3K9Br/dTbBdK7tzjM9rdOhytOlFq55mec/iZ
xMjSxk09SDXhFEq/MSe8vzOI6ch7e/IPhMGQFWiKHRFeqwor7jggI9EYedHoLOqKRsnPuO/zozqp
Z/LMLi5FotN162RvKIhjanpUL1WN3Z05hdEWx88H5OxFe4cqlabzXk9rS4qa10AWXGYOOP9B3y3V
vVUAJcif9w+8EWRj0amqLGNlvZ5YVXmy1vhE7OV+PRXIa7bXbqMcVPmJhAtiEPTCKAM4PCmGKbi9
pEKDB8nriRRCG0x1sc+nG/c0YkvocOCbN157jW8t+sFnAi2+37iyViH+5yriWeVQBiqk92rXrMWR
4uMJjt5gsSsmwPCXwq12sYRXTY/B8DR7D3dpAPyw+nh6yc4WX9PRR/b3Cqcey93TeEj0McyFGemR
r2snlSLTZpkkvTa0CK0F42X3qvPU3bxbGXpOmvjbo6NAWPYYaVbpSbpIlPqz1J6C2nKVNVO2Xp+J
0UY6gsWbQKckBJZhUFh4WJqyjv6ok/wJszLUDu5N86yZN6u3diIeFeN7bA9z5BQ2uPhVTLEjVYA3
pCGO92NzbQQ4ZNC8Q6rh9bbFf7Ep45CRGoDpmUABmfwoI/sv9p/LUb3Ln+xjK3sjAtX2ziEhvZtl
847KD5+aMsvKSecw9sadZTiqG8OIV/QkAfq07fJNEeD1BuO1/hf9K7VIZm59e+KOHeFGGc44ZdAf
c/dSgQ7bN3q/NCeoOIrOmfiZTp33Rya6wwmc3OVeBcbMY2HxQtPDcptZlVgmMLbjiEOeoBH10m8b
IyDm0mCzyxZr9YscKc2xSdceF3FypYFuVKrRusEsBZbgjbzvX8+mhMX6gMeprtCMj7zyDdWSkyBV
IfbJTRKB021rjWvbsVJ49yOcWCiFTwCkbwfjsUPBwctZK6mZhDf4L3YqoSOz8SdjvzhMbNy7mOzm
XFxZHiOeAA1sVimDNFbq/G+v0uf/ZCG4xyZWZQvEOqLzWUFBxOl0X59QvjaLi0IWOa2ufgXtOGLb
uGtnytRDNBqwpftFkJSYJwswHZlF7yHr7zofjZhaoijNrE43/jSpbi8QMUpsk5Q8tEp7QUnlDFt0
hF8X3RbSn9lmcNoZzB/5gAh0a5CK9qrJaFuWVTDAa22S9U+JfrT0iBgyW0AcVk7JxFL3Y1X1bqvY
CtzU1ZvC4ByiiYqksoScVHU1b/bDFYrV+iNxRC3mFIqmOPXo3mWZvRhasObdPnBLCN//moS6coiV
rzzDi72waqaLH8SCR8zXzYMhpYb/hnZCMqP4V/PRzvVQ3KYtBMBIP2MLL/o1MsmeTvpbhRkoAneh
AtXp9+zclhpjAmeJdiXhfv9Xzf63bJFdfnlYyl5I27RP6sF8bLZyFs3imdXFROpUrGNjUMaigYsE
WXvFk9ofOD/BqfWWFlg3c9QY6QxZMJkhq+AfbZR4DUq8zV1qlLjtKSYgQDHJCL86DbxJOz4tBRCQ
iSwOQ1JJkgWo6cp6bwtLnyUqf72yGHxRo/uUVYWjNce/1jzsalkoM5YA/+5ET6EKLf56eqxNLL1l
uuAVmcrdzyOXuUKFXQOmDUsB+C0mRgsebOBpDJvCuc4RyNvB5ck60d3unM6J40tKLp1MHt39X2mU
PygEXmg+Kx0x280LBZsr/QnoZTGHwhfLXNkXNIScSTFiNuQSSXnrgzl0PxIKsIzr/iYuADqOcl8X
stOe87C53GZUfCiRBYzm34zp1+Hgm3lnFun84dGEOutiA0k+Hai3GB8ll7XTgL/TeIk6wfPB5Cj3
TW+xVEkTo997Hn9afl31L6K5PZdq1dWU3xkrst6EaoPpLNbXzFLqtEOIreWB/O8Vy2CpTgvqHzVC
ENYmhrb5/qF5L4D2KIqCkwgZ68oPtrp1ASxpPy8FY10s6h+nzGts0WiGAdKufFTmMVuY1VEjsStO
hqIptizkm9Yd6/OVkWRmAlSeyRFzFXX/fnwtLkSN0A0k2ezdSVJIPfLBv42uBFMsGuM+5IGxOhkL
8UkZrVyvasq5JqPf8MPZoliIgchsDxr2opn74xyIPmHxZ/PbizUytk69BuzmKGQIiKGYKpRZQl4R
vJe6JQUNOrOhcGL6sLXUXdSmqx1O2VXOz+WIrHIr3ZhZ4aVxqbRJp+YCD1DLW8DGbqiNjgpQSGIv
deCmpvQ+Q0ooz32UGRdQqog4PaGJm5DzowvVt8ggRU0L80dmc04u1SA8SVF0g12u2ctnCOkf8GoN
O4eLZWzVQTDbsdbnWrP/dv+FUdhtNSLW4Vvas8P+7jVbJgONDhvSzNujc+cgvvg+dcjvFtgk6kzM
5V/nlmxvYxvWiGM1OIV5MQK9F3oWXGrC8YNBusuRS4eDcDB7mecfpRwH04ErEb9KGr2C0PP8naZ5
Mqf68E5d5wGb1fYY2OAnynYjtO8awPwkPWWsXI22UHS/gdEOj3Gwf7RMVCvRkD3Q47HqQhQyW2DG
7Nyu35fAmvJalhsOzo45yse7v6QkScVTxquN4yuFogQKB4awi63Y2+Oj35sfOoSnoyHJjjjtoFXe
VzlSnYHvVB3QhZuSMwZV8zbgMr2N1ZNyZ++8pJST6xRTZRoie/UKBzc9t2LYrem9W8n9wwen+qDb
1AxKkjnIPIZqcmQGxAs5CGR0KmeP75uIoYU9jSHNdPtSrXzTAzJyraqrxKDpHRdEBzgK4zE1kUuA
FPWgvG1OSBeEvqBVi6CB0U1BzWQfO1R5ViE/bKiLzYPM/9yMfoAduBtN4NqreMudmj1DxUhIZgeR
hC7nY/ZzHBU9LryYpScYt98YnYta+ZT6SEGfvRcs/V3p+KKiXPyMA/gXfH3v6n2XmWoh9pfH7Rzp
KnzfwP6mHw1gpTd0ENpLepoQwNXoFeuPuk+3KHuuONifbRdKGwviQ9TqkWrdOu81lIDpcjc9qFWV
jEgSQWdylmPCZhqSrfXGcwK3lKNPEfYZVA4v+0xwYalkbPLFq2M8spNQ9GWCOLVGy2WEuG99OKZZ
aU6OORb3DriUe84SGlds6ppc/WzCF57IvNkATyNDWXGyoAf9lFL3E2FZuDy9SBxFuAd0sFi5QBYl
acHoxYC0Sgpuy3dZ6DPyfAYtLnPhbqTWnUEDwu2tmnKZFupIUdYrLY6cmyAwlB2EqGkXJ7mLPBNJ
frzUApHa7WFcyYTQcWVVRIB3yhdWm8ENMbgXA5BgIfCpIN2+egZPyuY9cCkBdX7HPUHBXuQZcBPe
BkjMWTfYqqrkaatPc/q4H4pdhF4bGIHVgMTFITcG5AS7LpxHYRtJzeSlMv44YK9d+h/k/2YH68JS
6mHD7VduXWFlO88rP/6betQw2aZDg8Ng6NNzhEYQzNX5UK0G47cotjMM5RJb5Naozed3elORTI00
H0Wc2f/0ZdRC5vw1wtn9iGJ/qp1glHQIQRF0GE8Gygx5SOjkMub60NBPhfNCyn76eFmnAZk8bu0a
gGAiUfSycMrzx7NEA6w5T7+8NdEMiOVOD/ltXWiHT6OmvkMmCxXSEK/L2hqozpyjmrLYy1T6uZzW
TF0KDlO/T/47Q4IxqtsI5+rdaugpO10K7bn7XoJXSV3BCbJWmjKyjxENwe92VJfyO0B8y3lmbO+o
YqQskU0C8b2BWa8fTFCLa7a1H0cKzZe2KkYNJRtexTnSsylLlP5Ep61e60ccbf6UORQlZU0zUYRG
5JVb5HmckmigW0vuCGCncQB7av5rinOqRxjEijyLZqKV6LRWNrXsI9tcsL6bwtLsFVfPxy2apN/b
kHes3LLABRr9cxOL/D8RbVTX4K1/NtxrmT6WoBjloDFBU//XQQdlAMaj/PTwPAPtyQpp5P2AZMWh
hOtOe2XE7JqyKdx/8bNVS8FsE3Q8yC6gRZYfci8nDNoqjQHlpd8SbJcgHKJmZ5c8jC1Ee4PvuhGW
LxIXxjY2V4mP3hp/a7wKqaFYy7t9xGL/FxURpe2jMtTJg52mSSoB6OHPgRTH8db+xejCrhQXRdmZ
H4H6GfcgY+PmTi5uV9YE24ubBhsHg4IvztcZnTgUzkUIXldIVy7I8cGgpWxMDtZLvDDpGYhFKHTE
guW5dO+TDfEV5gOxUUAaK15RJ5y2pEQTlFI4vhddV+hGbA7rhYUnwRLPMGeL6w34mnmtajs8TinK
dHcgMTxTlcbgm6UzLosA6dvq02912O0xI8adA+qSYAmn/UhiHhHbFOmnA2v8Wfudzj3F4BbywcKV
IRVQiMbuLz5hNfdW71vwcrH6Lr/eKQ7ib/NBy4KQPlGDEeAzTsUslAJpDjiaBmEHRjiPxYyLjiF5
5HCmPASXFS4NwI1y/bLljfMsM2L9r94KBYoXZEStdhKq+QT5E0p55PDtPBnkMYHuiNwWp6hi3UUv
tTad6iC6+Hu4I0A8yCmXIliouwmBM8afcYxYtVzw6WM3SYeWuvdMu4oQrztCuSUzIcblreNNNtxk
6M5YfeI5G97Dxde/3sa/AjfdG2ItKKWwvh5JkjNNptnnybIXxvhz+89PxglMJXnorlfH2gUc56Wr
IriSEf07i5TX9kZX91e5giR/FjOB8rqCRKK7P/pGdAxUrvDf423QsSkh8CDQb2lH0pxvMFzdnIXh
HQ1yjuUHEMSQ783CzUVQi5e14LBBm52MqSTKL4XatnJ05qCMFAMxTLFhXHs6QA0gHJuzaNYsJjTF
wuzpRpZmvhwszCN5GwybQwKnxbQpH5lSnsKpyJ+QCCYmFP/CYoYuBHd1xZHsDyYwzHt0e8FtoByq
OuMPu92ZO9MLUWwINoO5eBwh6/b/9fDFMjYrqwvw8RrJn+HWXZ1ZvNQDCC2WVC1ql6ZzCnDHaBqU
qYimv5cbwB7kf+ClgV9UJ0diVGMC7S2YoCf/J2z8gyM4Y+KFgdmtd4cMA0We0tQD49JOUt9CR9dw
RWc00vhUqGYkdGSkspJ2oxwaX7TJJ4luxedWDvO2OtOvlLBk/Pep22PU53O3AiyHJc3OdDE90C0B
dTBkA8IfswT/CheDvEvd3NnxZTEkCkD7OfNPQidmw9l+Xzfbq/sZuZ2y4jz8MHaqQFRQdgcXdlvU
OPFKlSOqBW7ylhldVE5WtvcMcqHo+fbssuRJ0Wjc/1mO7kZyePJoKd/BGMMK3kWxmaPGMUOMG76+
ShnH0LpbOtGCXbSDFGptqpBPfLGY9J50Aur6yDZHevAfx54jmBlf+8WnYgiZDjFuyYyahmAStbA0
LL14+n6sW6DbYdFmnEDPdNW9rjce1WqC8FP4huWZLD6y4UJkGsg9USRP3ZRQoSchwvx9y7kiw5TL
KkiZBsxoYFSrH73HcB3s6yiYvno+ntCpdOLEQZ3qCbKu49mmeq8g/jussa9eJtgtTpVBRKu+Lnc7
ZS0IJD0iJLKybc9bCEHjAAs8KxgkbFI4Le1Yf1FMjf1R2nfWVkZJ27ZztVbwETpLQBFKhF2nbsLi
jhKiKGgZsWIA2/b52AMrk917Yj43/nawtOTOJi1639xzB7j2SyU3n6p+jieRcP2Olah1Ep858kKH
cv+RFHN1VbR0KAD2wbjDjW17wUYFOT2EMjhmIihrj30mkp2tT9k+eXmvvrI9nk/8IeU6BwLP2eGK
HeOiylMZZBteVNytAjNFrUIdGl3YRCyhvx9j2nXGVYVpMASM92p1AlrIquJ2CG0s3N2AIoi0Yf8y
S7hGTm5FQmslegCXp8Z9pZMXKWZ371rCjudyfyIENWh/9hyDopwmb5rc1H0HCYwcZ5MoV3Asst+d
I4OMOCKnp2lbXqipWlgvEWoVoRkIlT3GQ3C23qoOOFDw6CnL3jJinIPE2eYD2UFnxnKa38qMJc2A
fVEn+LvQeG/q66fLsRDnJFbMgjsN9pzT9wUxSSqmGPPkPTEpbc0hL8Yuig6COfPsz33MJkNnKOUu
IF00VUglyDhoqlUSKuuOPOvPMuKD48gg946RLiDCLF2ng/KKIjVhJOcS69jN68BvsW9QMZ3kbm0Y
PnejpoGMXiMvlQj3/bqso9+z+OV/Bokizq467Xb+eKcqufHZLYcgYz/SD1L8reZzvorWmNFriAxS
7V9L5NwT1SSMb2bbVfmxITmStBGW9bABMO1jHV4CRp5gKs/Vv8Sr77zO9c6307l7Coc2DKCP6bV1
vUflGdpttcefVFhNXUrw+cvH9tZpruzItZcSA0L82XkDQCCWKVtgLKgI13kJKoIXj//KL4lneBCp
R9S7mnyifHtQsp6+tmfRSvcoMes+w4WhjUsygfqIpvY3KZt38rx+8irbH1PwSJkBntbzXHKVSdfN
IK0HXrpZflkygygUBjFq7LuJW5/fpTp8VtEq5t/xpuHV7/WbffyMQYgEoLUSRx3q2ymbvCh0MXrQ
WhsdyI7xSZafgcm7afsyEiGKd+MHAgop4jQuNZrLVGpRCfVl4HtIhW5Ode1OZx1xynXCstxI9cSw
cAHz7LHSyRunMsAl798BcDUgHZL7TAm5w448RePOFuOlSlFwC9MGZ4UB8XugSwTYoh1lbgq46153
E1QbDLbL3FZiEC1t0BKNzCusVYZ2C5Gvzckv2L1WPm1zxTgpuwdwmYQtpKfQkyCFLtnIj7+H4v33
Onb0T57jxm1jeoV+YBejpo/360f3nji6LqOjvEOs4jAexTVnXiw0/nGvcaFCuCHCx8DIe1gPQWiL
r/1XmFSI7IpvShY5hGmGU2040YrzLfm2FwuCd6OWGj0fpkVLpvj10TDbyzUVcULQSZ5Wea5+hCWf
8boFxkuWkmpBgK18NhX7fqu2J9Cf3k9SGFyhX3fmFMRH93h7ni/97c3XzidZHTO1sx0GkM8q4XtT
6DWtnpJijCR0B90q0VDeR5IGCFWlpWrnsu6Keulgoh0KECUYRNQin32plHBH9JJbR5mTbsT3HdSq
gzVD8hcqn121ykf5AgS9KZN/+bCbnynLE0BbQApcPpypcCBTOhVUcESnriwQps2YlMGZOnO4NEgS
nATPQV8fACmOTHCxoIwXqtjpLSwjxKWCXyUVR28NMD6eoe1ZOKym3vVkyaC6zQSns0JR1SXlH84m
95IBrIrtWpyFHvxeaJESrZsrPhP7+6TxVe6/iSbQIoPpl732SVYT1YS55QImCWX3NbuTtyWdmUe8
YtIVQ+yhFeAHvUncDHVoXj7DK9G3wlxn2KB1ea38OTMynIupIMQzDZdf/1nYNKgNO5YcJMRqtXcq
a9bdkaVVMhQY9YcjoViW1M0q2tp07c9aCZ/u6mmmBDyXcTwoKlcHlwLu2ghuUJTaSU3rbugxQdIo
K651QimaQu1AyGLJayqOFTaISKDFu2t/lgooKqxRIU1K8claHPGx0ApiVTEvX8RQ+4JE4VkqZ7nq
M+LSQjUZLF8IigeTzu4bbUeXgqN1syKiSsbbE8BQblmebRclcZhYjbEAsPE0oL8oC7BcfhnbePt9
v/i9qv1v0rt7k4lOyLymGNJIn+fdN5lsnWVScKUtXUHgyZLM0KrpDndTRfDk7X5fwj122ma38psw
v1NPLmla1FovygFTj7JZssB6z8GFUgZ71yM9CaF4NdOl8jZDfhI3tZ02bsp7a4+nQHsWjG13VUJP
SfA5Qy9Xq7bWy55HwHewIgpkC+7kDtKFXuaVmMe8F9dkk18i3r3KI5noPhkEfAXH1pbZ5KVY3hrK
vAqFzbeiD7stwkTUMq1RdBeIHvQkH+8ncL2tdHvT5W5EBM+WF66PpBD3julQpo/C0LMK1gfwhpog
/tXSh18x+PZxRv57Ev49kaIUK1VU1NNldmMV85bFWZdyyjWUxQ7wbd/Pr1okgkvG6nbvXjQMz8ZC
bL+u1GVrCX2IFpUsgPdzM8Q2ydW9JWFsbAGSdlqOCf3ngAzEEPIYzrlF9IhT8QsxXVzmYlHHGm/i
i7BR08ukZtNhdAaztQWQq/8G6FcwwSMbNdvXMWWWvgRK7uGfR7+EvrAg36SrDD7RXaglDHJ1/S9j
ulCujShDOsFMxi/q3ePy3O3XBBIiEz/0ongRudop65BH1gQgDuokXCfGMyFswcMDUSt8PlWpBEey
mAnhd4bCZg6+I0s8dLji8TMe/8etzgN2hr+Q0iwzokDZNbykbh8IRbxpTwbrjVWqMO/84mw0xM2+
HJuRd0T4Hp1widuC6QSaQtQAc9xXvTQ/broYDjeWxKW9Dp5i1LbgrJE1jA3hh4nRwtxJEXY+ZzV+
nwPgorl/rUYJkEbOJGTATz/5lm6y3ODw5BWr9CzTejnkow+BsWUNasM55FiLBO+b5Xsjra056trT
WDiq6DIUU9bnKCZuePncskYci8qZhDGakqJyghf4zQQUdtv9Zpa0g4JqKs82VZqbJnqQMu77+0lk
y2jUf29TQMd/UUjrov+gbd4t8fmhujHwwmr70ykGuhppnPcHQY1HrDQi5Oj+Geo3nFg50t+YPKQK
i6mfapVZomIHNWVP4P/PsaqfNAE1wxD7IE5YTbhjGxSePmXJ2+yVKjQrC3fBYwtv9G+zNApSsWN7
FJYnJ76KczegYXoeJhO9WCXzEVnbBPL7cFm9Gk21hipcMAwmZfnxGQgbxlX+aQDUi42N46KPPjbb
SdEjAsuSmWTMqI6eBnEOEUZQ7DLb/6ZeP+ek9NgQ7xDV/QhLDfy8jBRXwWrM7Hx0fUnl1OP/ora8
/atsQo0cU5QmSweZSlxUDTGcS97/f13VL/+b49y88meOA7iVASx0zSCplfaN2tBRD9Kw9ZorRe4i
gNXD80T7IkaOP3BgIoOtxqrSkRouTSmmsBbPgvnHc583nQVaofrWs3M/SIJ7eugKDTDZ1yjkZ5aL
/8gsYspyFghCAeIsc3mJsq63wz5Eau7dk8ToiaHpBrUMmLQq6chKlW0orNuSMYn7Lh4ad7/MHyw5
iRKRw0FK+lBfOBhQwoIpjztLj3ZPxYWw6efT9y0mSkdQnc2UiqXrjLAqzAk9G69WI6y9+uN1CnOb
1Agl7sgmhXRtpf9rdiOP0GuZPJl4gUxxn9dFyVzbUKGyiXBeVz16Ds5Cv7ujWaRzHd9aeqd9laUh
Y9wA5eOkIW1bPqhiC/kFGBrO7w3kn/Yb2MdjFk74wxBI1m+OTxcSlOSTDk/sInx9x9s0jawWwcT4
QLsVFuc08uHrZbVq97a/BqnqaLd7wO120M7hcEo2pkA2mk6e5UFF6Zq0hx5MuLU9HFv2peP5jdEV
/qovVkute3xbdclRQqCOngYO08CGPXn0V5QFd/WxBrVfZd++9IWzGG9pWbq5Xrcloy4JYVxWsNuG
VVC6b6s9DduP5hdV3qfy5PUOWTcqFtDj15Nh1v8wU782z6dXlSbdYYl0IGgNcL5jfIP8NUW54dC9
s37ns38J8M8/0HEDBO7Q+CCnY3cMRRwyeRGX117GZWmS/r5yrwa4Ia0gkaACefGByg5+CEI+E4ZC
tten9gI8Ps9q+Ry+VCZiGNzLjRTndNt1U/Ub+OpwfTX72JQPwJv8daRkt/QE2pkC8cshgpc4uWbS
BFAI5ZBuszPJEYdcKr47Z5ixD50LcFwcVV5xdsHUyKbLgTntG129riAFFR3r2LuJMMtsfbPXjqLU
rsMErhFzwFx+QCTIZTYRCRMn48+5k2pZM69CYgmWZ0tJo/FtD6bfC07FBU2VQkSNIk9IpnyNktLb
8k5198CfL/WPvgre/W2XbH7NmDgPr635hWoS+RFcIN5jsHDCPBM+IdeUz9v34xE8veBH3ZayEarj
+6aNRJUGM4kON/QCZ8Jh/NlE/8b7SnNnehaL6yEHCHPLO3YMQzN0cz3J0MlueiNaQbV0HEf6FwME
lRioOIG1vw3ZWRfuQzCEUPU0dhxgPLNKaPqSjCAxUQNYxYwWOD9wjY7qhFRmrE5otjHsZsYcVHpY
QBHkxwy/lSMDL2IrVuZmjyXkPqLDk1N7Rh6Aj6FIu/vNETUPMeGrLleE/eTwxsCG+Nh3BXWrF0DD
fS6/M9eZbzV5r0slow/Udw/b1P0hCNy8nZv23sb1z8QYeXvyOgBRxOjRUoC5iMHZDwzBXLykkTqO
xJ+7MjrzrwNygQ8x/Y2W4osWL69nAK5D7VOSoAVkRgpfy4MT2itEhAVCnnnmaCUwRHVTrmN9lkCz
T9kizLk0O/jZ2tJR7gQ7S7vkV+nILyk6AQJavUrLpEE9zls53UMDneuV1wsn6zJxycGoJJyeuBEY
NYug0d1jIuwsnu8bPk8YD1kMdUAF/8Gm7ZO1cohbAi6b5buMNOuRNWMC9GIxTDAuRLeM2JUvovud
Bji1ibpFxGz2EXIU1lCk2tm4PJWW3u1y1lemAZB/ffuCqQ8sI2nrqf8MdYVIX0EQ2fNQ2CPwCLAw
JLa+YaaIh9HXrJdO1ChqDFQE5S3PC6Vbh+15cdD6GxRRQi+fDoPCoPM/+gSQzDhG4sPDci2yImZL
KWYn6TYiUmS1wjuEEE+9rmZQzbo6BKOO9iNOBGvX1YYDH16/xayFR49fLDAB2IBZBvjIlapV5BtX
vQ0P0rBOI15iUui7lYClaM9CcH+vR2Gzw6lpVMt+g8wEw8XDgHtb4U9LtPPFmAl6Isjt3pXYUDq/
C7uph21/MoDU5V8/2eRUeiOyVXtwAambdXfN5F7FWhDyI5jA7vPPh3gbeEjdhh5oyM00zowp3EkM
vVvT1rd1k5dtEBoA7CCpztzQyC+nX2Grl52pTEfT69sDK1wu5gIzEh02Xen3YjWU9701VCpO9Ewz
ZNArP3WEmDAMQSqsMpSAFCy5ak4EmcU95QCslNZ/5HWroIrBcVMrGNVknQIgkM4SIKiqkDckyeGf
f/wzftyBHHb6TM1X2YHysehUO/Qm/yMpXbmUINPGfFxxaRneHrwniniCj4S+AZxIGvkjIwkR0EAD
+aZs7/ZLStGm341HNuQH9zvJijQIw5VejYpz1d9l3IW2A6VM6HJLNZaGnXOc37y7TXm6gHEJ8G80
jDqRIhsGvVgKP9sbeQAyAhtI9n5eeMcF2kynq5Ds4A8yaxReNUikgtzm4LXSU91Io3qTyO/5TSq1
WsL96sZAJD0i6HFabyxuRLiMfLV88k8sVyFsfew3cQio3SWUOkmuDNBjcI2e3ITAT12DHbuPMOQx
2dv3t1FlC7Avu5Wvo94oHwaC9w1umsojzYF/Ry6ctkrztEjqGeST2L9ZpjwmqX+C8ZM9PwAb0+f+
fdH2fR+2iEetjES4fbMt8Casx53DPMP8ajF7FRE+9yPvXLaE9U80Lew9NWViidLi55llDVHWDhdk
yszNYYZTArtAjLf4n0pOgXV06292EvBpK5vB44FlvK6bxVYhkZilEVmf6RqOa92cEu3VO1VOS2YE
3AV7vRBG8jQCHdXkxiQtIZl/4uRvf8xG6uNDIfnst1yByGNI85Ds52MqY2r5RrwzJDpfY1HSt2Wi
CASQMDGzyeBQ3/iWrA2uOWde1vbIjnyQ7u5Q3XRTuE3chomIpkyO8BJCwroJhMXOOp04vW0MqD3v
p9Hd7SdrpVWY7/9NYbPOaT4St5GKjCiDDRJsLiBsZ5WdINxTvqFz3UavM15IveNpN3dlzIcV9teL
WLmMbhR4+TapeW/Xjh0c39FuUF+1zdfDb4FU5h4fBSWdv7drXaZ3l+5ugRPge9iv4AU7PeLUm8Se
FssWqADovFB6KvtsWv4HA3NFUkv5s6gdMdwgQpZzCoKWvFLGEjpaN+W3w7uKm2gecV9R+PTncsoZ
TT5CEOfzddfp97pYKyduhgerWZGS6f9MkrHlGf47zXU5KGLVE0mkH8PIINdUgv35vyOMwMDbqUxa
wm/gxxAMwY5GUWePhgI6Q3uYkGpQ+6Lk+m6vgcxsDSL1cZFCusPa0WCJv7ExAu47jImHW0s6xRMI
ZtPgoErVldbPLYDMhd6M4WrPU/04R1TZEWkuwkhD3UUPjA6M3+VvjyCCVKd5//usAsbBhU2gyg2y
f33MRWZC188T/r4LZAdduMemgt+Z0nhRResKy/hE5T4eqx19XaXw9UJDXdxHOyX2pepHosJE6Ty8
LDHsHJygg/OQB2kO1par2MfgPVj/P9U+EWu+ba94ch7ZAYoWS7RPOZ6G5K/wOZJehweQfFsHlYMA
PpV+LRW9z0I429DsqVbZPZrAs7LDKPFc6xnsN1FCKQSRqMviSTpXr5Ma/rFREuQ9iEtpoCAGvGxp
LTZGFALYgPorZSortc/zX5Uq/ehfzaIbYpxiP3L1igfcHTHPMPvLNxL2KFXaRRoKb1VZbrqROWrr
nWQXYTJH9CAyoaiu177a9s5VlOAWhItbGHcFOqUo3SkHpxjh0ksYcPtUF5VRZwW38qCi9nhBRWx9
u6Af2OqXrlqLIn8c6lCXdXrZCOh/9NBZ6R+jHntIhNjNqYR0NzklC/CXRO8nI9a22GHP4BR+KhzL
eP34KZR6QslBpBeZBs3w6g9iHIGMnsObd5WMCWQRkhrZxvyBKDzT5V/IaqWb2HVNWtaa/x9gYUZC
I+izKi1aVbg6Ah8flaoAeejQSRalRNs8cjgX2UOiH4baNx+eaDHexFRmUuC3e0pGd7pS4EDaDEsc
qot1TuPg6Ijs4vmqsLgRQ2z3LmMYwuOkLXWzwt46cxDZjAzTPIW7QNmOC5vPwg8aXP7TsCUdIkpl
ViIRfVmAv2Xn9l1kUAMy7VexNVTbiDmXngP8k/Gn6qsnofOiE5H1KA/ZsZoq2P1kdHHGXNYRLJPq
3odeNth8N5cc8CGfTd+TjOit/TBPhvm/oiuC4dSm63OMVBtppefor93TDv1XB8rcsOOlthAkkKoy
XPSDEsi+vpmjsOnC+yKdSEfv0DlDfUNot6m5PvVQHacVSNPYhKuw8M5HXhGOqoC6MY0arXggs1f+
xa1Y/tPCauGowx1WVEehgGAadHsY9EgpGXfX+ogVAi9mbAgyHAStJ8eazltYO70EwKx7v4MY8vH1
CN6wMK8oNBfPhYzoGTWOJrrPht8Hfuea9g00/TmPXA6wMB7KOQJ/nCVedaE7DXltAEQmdRBrhjzh
+qbuTPVEqWVWV91Cu1xFbmFldPpBoN7RshLfqvFo2N1yAeC+9f/h+UjCyJTC9QYwAUnnVf/wQ8LV
XZMlV/O8fdgOk8D6smVuooFFN2DFl1URPDRuG3nYgvC8Ubt4B8Gn/XUsEwZQjZtGjPDSjgkN5e3T
ZMHrfm0ETs5EcMtM913X09cHym3qbeGkuplaqozvZeKE9jLJhoROrHqnz4FuCsrIT3YeXPhGpLJF
1nZ5JouEgI7tOitBV2B5564v7PmjYNaWIZ3CVt5QlsWSoVN9MZk3Ogo6milmqyUMguQVaJYuxvbR
Zl7f1Zf1KhFFafLWr0MKwx3SF98fGmt8R4UdFsaodFJiINRqSw1cupf/qTFxggt6sdPF7wKxKPf4
lwhgzHnl5vja5FH79h3gE8ojGvNboutTfM9UXOXbCwDn8g+kGCGVjAvWOc6F+jiCFL8Bm4EgbE6w
Gtemqs5SmFvUBuSGPafDretfR6QO0K5KBoo13HgA01xyP83Ls1DHv4GKL/BGA8Kkmy+WfgQ8hTtw
M36N0uQV99UWRDRk0/QKjnrzjd9tFInjQVZVvQVyexYpMpK0C+AQI06olgQdCn7OxJDP0GK0lXyL
UpsdWfqMPgAbI3iWlm/wOTsW5QQiNThQtjEGiE9+Fiby/20YIk/bUEaye/+YwTNQFxfUroTKrzs3
0orzMkst7zzF99UENO9dgEGg8yualyR+em0wvgfmpgwt1NsQ6bMotPKskW3KQiyG2j85dP1xl3b2
jwi0RbbJIAcuByCPVKhmShIjzArRNAmcJfnXOG4Y3FVk0JWQmk69ZO/strvpCJwru3tMt297CKkq
dNu1/9s5avFcKWjaeUFs/DEciLOWW3fHmCaNlxJcmLarpQTZTyO9c893esIk4aJU/wQ25JIDxtM1
RqIt2n9DRs+gVaNgq5wN5tjfaeF2GIOt6BLzboh9QdyyufypCzaQSPMvIbuu3jIB2WYGfQY6x3KY
EklEtuzAi4pSXGti5CYoC/ogDNitIZAh6SpNXM7czMJugMwfkZepXc58KUTNJx1veNuZ2bTDCueS
tm9DrFwjWvJW9xcBIstAp5VsANo43xg2T2Yz9VIIUe5cBgNc5C5WO8AeShjz3W9Rv81izieR8dJZ
uzGPv0dpxrnoJtsk0PrBxl6ZEZoTTTY8gzhzwPL5ob7X6I0hAjN+E6rhLJpAFrLOhoEIAFGVzh5a
0GatMtW3ocvnrXwvuhMijFYbRU9+xy/stKl5EhFUaC0JlLItd9osyzMcwO/fr6CSl5rN0Bwc8e51
gsGeWxVRyKdo3x5rpnAaT//NKQpF3XgSrgiC3cHwgX4ENX3TWuwolyPsJbDwdw522Mh7OnwXPGpy
IyoU4wRp/k5DBW41v3Zy1KNWMkk0s0mQLOKR5Xo8LRdzsmRVnbrdjJALxdtmiCFWME7CGs0XbbT7
ZLx+QA/2XtDKMM3qmbIOnwuEpuUJrU91yWDbX3ER532sBn08T/z88mRfEVm6ds5uqXEXOu4pXHyZ
UBTi993miPEPwSa6XR2JwNbnWhIlU4gZyWfneDBXRFDzzZCY3IzLfjGRF1TQnfrTtyGMYl31B8aM
WgjPeGOfnFACNHKF2iFlXjcdwf0zMLxMqTSOJMJFBIAzYBgRNMUlBa8A87TM5gEVzu0vMg1AfEht
kedCvkmLVKhbkIp3n4VXOKrA4MsYoP0Z/A/AZ64mjqm2bfSKKOEsyuhbLtpAcDqcrwevtNPqVD3q
kIFf4R/VlNIcQybUSEgzaUsZFSecpAK/+RnPat0Ao7nr3Rp+KRfT1JNP3IbAr8dWC61gWX5sc02X
AqeftHWMC1Ix4/ORhgqoMUr/zj0e5oQd03PYUkd1J+EbUaxVdiX/ud4oCKtCeV2ojrDz7HxBd7X1
i8uOlEHKuM20KeUETZNWs8QS+4fkJYHszcc4KyHeM5AWslWQloAaKMxLx4Fp9sqjW0myyzGpwq7d
RG3tfhceBfhC7vw5Fv4jcKDkXw2KwsqbUmfhMHNheai+iS8WOmLrAoqLWs8ExOCvY4oSa9O5CMh1
RJcTHM9ItpQTyW1FH4Aaqit9SCI8O+RosDHTD8bZAFrjkLs3jxcWeHSjEX6FwSs2wLd6XJbXbbMW
3C7qOyb8H9V0+OZD5u6muph4WJtrag79OFEFEpAht93j9qXsi5spqaAR0ESJuujJ5jRhTjqOPM3n
jSGu2HEF/lfRvft8R+b92843PknJ8nIKOmwIsm+Ge6vZrBeYC4NTEgHmCpTg3Uz+ehZ6ZLn/jACP
ATv43Q9qS7ZV4BHHt4Nu2X+d8ECZqUbShV5ygFldCThauycRJ4vsY/OcKe+8nq/2LFSiHETe0rsC
dtF29QX1ZcYwsElewsjFavNZ/dlqKd9wLHwerMcihgYYfTB/Xr2XNhHHp8gmu4iXSf1X5l0WnN3C
LePiWpOpMfJ2I9nfuTx+PR1XhuRebqw+UjSAfZw+ilfHcL9DdAP+IgAvcFH/tQ6Z8Dju0QePHRm/
zD0mXcoKH8QVORXKyV6zPpnScXOj3mbjo+3A98GFYqZ6M32Tyn3vURPZ9fWL00Znt92svfMFgSec
eAC/ASDphKKkM29/EOb+MCsi+A8GzfalBKXfScmGOYqvCfvDLrtiR66Ijz3tIxnYE8mAqbh2eQI0
EU/jgYZJcEmdRcvkIsWNOmHmirdhZifdCP9L2BFYgIkjeadRLNrDaJMiWm1lcLfIoMAA18lhLhxN
lG/lZPiZRLdGKY/xwAbtm54SDWAL8y/T7D5hMtwbVrIOG9jbZ80zbETxof7Kd1JsnLwAY8geKSzY
4WRY6QErirTMc1pGq7D/rfF/7EYo3TiYES7wkGuhgKUCr86r3JHL+HK6ZfoBY81dbwDJLrxStM8k
lWljfFa93mXw6Wr+wQ15ku01KbsLDYE3vvQIiUXrx1cjEWJSRAuIJDC7YNxDqVJA5eTK69dBWVtx
fEjdIBqleP7q4/sTIjiN0lvo8elNPW2vJ8jSfRbTND2KEBCmHeRhqLTZyFRqLKLvidQCjSvu62cV
zcwgTJgMhqyktseoUyYwwt8Obz5YtISdpLtw2ze0Vlp6Z8RdujjhNx/cEkarn/AWYkcu9vNeBGEe
xtLmwplfOX9m5L/iJzOpYG/YWNm/iZjvJn3NTPGrTdok3WZm34mO0LIRpqvzNY4HfalVyQKLIKj/
MnOBU2d07CYDIo2UbZsr0LkkQ5G6uj6pgvUU35cszqshlg5Gpu/vfu5dCALYWo2vQaqEtBUW00uY
yvB0qfHAkbmxq1X6lgxy+jbFH/9phhbedvwfJKqeRFZWv3wgV6hYait2PXJZnaCsmyeCo3OvUX42
2i49LOp3kQJIj+ns3c4tvO7gOdrHNryAqwkE9sr27MILoH2Qcy6AmSq/48+vw2PUlz1YfKmTYM1m
5n16zVYLYDw5ln5c+tBgkS0p+k10IyS4baa79zlpiiIhptXEq2AB/Z310y3fqs/IZUbTBHdkop1W
0R1QgHam+J5MG0zVFbklRuQey3bb4m4dH3SEgT5LjQAg1rLbVBqnc+p4jfR9mTRQ8TEZ7tHGpy4H
Oeswlv/PihGc7LYiZE82VZdRVh1leN3YOsTsu4m88fwn0KZD66dXSeF//OmjLHfnjtA8R3OS5Kb9
2rqRumrkjpyBNCRLM8xLfvRi9YKXbA8PFSgPIzivNjBNzBa88YUmT453XIgTsAqL/4tLSJQU5QkT
oDAUGXUn/bcV7i8k4jTxvyQkl7BYDZulrv9CfehxaRUhph0q+kc4WdWfKfzA1oYK1wxzgbFEFi+G
W/yrs2R7R2spthaX+aJxcfOT6hHELifOeEa4quymdIRq57XKKklSHRq4jwe5SSboutvnQF9YPg4b
nz47GsCHrYsfFJvdMyfO7UAeT9Hqy1m1EIYbbadmZSBOY6MryDvVNsQCdO67EjnLhIiya775BPyG
Vl76kRvsXa66GdjPD6RAufKE0zPOQyKee0bgNdeSgGhm7a+j5aeudhYOaPSqifvj+xSWVP5GFQBj
QI0KHUaLbeCvWZ1ClgOfiDjHfcyfNjLv5BSfR84R+WWzeUsjsZ0pGsFyJZ+Sn4HFcX/Cybar+M7L
MYu502UysYlVJ68vo8I+KF8hthpGYL29NMKXPXojZKHXNv+YVECQl5cohqFPCGJz3jN4/tVIu9IX
cv14FH7FBHVjEPhoMmsklEccuHRrOKfn78ywaNGGDajnrtmQVUMREKMDFNhAvPR2Bp4Wcz5iLomz
Fz+J4yt8OOakMCgAnBVsI5fd2JXBcIkv1jyUwi5MxU4nCUtYfIsZ0d34BjpLuF/ltzYiHQdLLy3n
8UyttjPS8XsvnBoAOqe+JS8rHPG6umqvnA73gjbTpqXpFfZaUH3YD8nr1HSZJtWiiFHsdY+dQKt2
Fv796zl7GNJy1kG4aa0F3SEPm0kTZGVSeGf3TA94rpHDjhzTj6XryTo7CuVCo1Sy6086kSCfzDmU
ESbMZKWaeErqeLATiMoguTWUUWDpmwgXJcI/E0pnharolpU60zGZLezBWSaeDkuAr7+eQTgjDNVU
hymxSgwsUumIyr5eMLznE6czQYyry676PuoHTFPKlaX1MFFTRDnTeykEcu0A25U/vF6fyRB+VaG/
zKYSsqf2vwOhF7dEJivaWSn4pyypTBkT6KAxurdXqsDzC3Hx3dfNUW1rnlSG6+ZGZy5Ob99dBfK/
TtjN4O8ylkyXFoylgZs8KtpPF9Tvfv/2X2gJPyNqF8/0D5xLzy4yInpEfVLTVxttHcFcn3kn9e5d
O1ig+cFaLE5Y/J3PhfpvesA9GOHmacOvZAal0hhvCSN/zy865RXQ/01w1EF8/VExCBFhXdxhITva
SBP1hXgX5TDcxuWEQJ2m/hmUWOxw1M3Iw5jWlHAl58dTOpF4hPeR+P+YhvYozjjtlpHpHP83COnc
v4vvCT2PTVKzKdb33ZQ6qFpyBUmM6O2XIEPKKX2m6dT+K9H8TFCovrvR52eTh5m4Ps4Uqz8veimF
5R9BiFviPUPRtZH6f1ooVHUrw3mijhP3YweLZ3VbIoUgtC+rJrEtRDsXVtWKY9I2+vFR6gkTeHdx
enoyq8cTn/A32x5R6yrLirVVdRjAuM2eaF0bkOs28Ons/Gbq7yTjQSm1iJ+fRY37Z9bnIELelc1u
J28bGA2zCVU4nB44DOKTx0BGRvMXKLcpS1aep7eWgRBpnmzR5Nw4syWX+qs9K7hTzZCdqiXHq28o
BF69jLdDKI2+/anW+JYvqBUS4rKjx/Y+TvYULaelCAc/rUR0t/pi/nQJE/gxG8o9kbwy4/DBg3XG
4cfZl4g5zHlir1lIlXWWfu5VAQjR0pxv8UPIwet5cQA5vSzIPZJuBSfziAsd80pKNCJ4JZh7dZNr
S71C3p1AP9JZXE1NullbqMQUj7ddVHbw+0wxMe5zzvf6g3wMcKlkCQF57mzSa4NjCeKeAtST3biE
ToNd0tgXbgJXL75yXhutgO3FiyqOdf/4l6DVbehSYwNutc2efEIoK7p0J01hKqkYe5r1+Aqb0uVg
/L3JT3V6qNt1BN/3Woq7VEZbcww5gvwxV7qcZKQpnV4jrBMHcfmgvnn+44260eH6NVkFcbJkpFE+
z6wl+8PCWrsEN9onxV0ialWQdyxIQSwOT3mPqOzUhVZdW0UYzWIlCpQ/WOdGcCUKnDYpVEUG1Xde
39mm6T56xkoyb0q+dU1dll1Gk27L/8nIkEgJixyk3Du1vw8E4pvuvvCElU5StmitsQeimk3y1STt
c2XrglGX1a7VaT6n8dPDHr/fJEGmHCaiK2ERJlx0XPRk5AOgQBsMsip1Zs7ClUL9iTVHVBXsBHs4
vErc3k4OxKGZb3qkC/4WzCVH10ljMkFgpsrYP6lr/a1YtVofPlHxuOTmMR4yO2gEgUrI/c4NeMwB
y2Oeorrg+Ls47CG1GxXpPzQEzdNEyUIdM7vcd39bSKo+pWT0UpxdWnkLfth6VlCYukaKHn8m64Fw
TLncAtqD1tZUOHs6TfURiEG5/hxfKaCcc6rH9bLZ4pwsXcrr3gFJBR66/3GA8Apm6XegTxr72lpW
zOXXX7IJfHE6A+wRXCQQTH6RoMN/WpsViLSsY7dUSDcdFQXINrr1nQgLBAtXDYfRiySjV/ZV5aqX
hv5RNhIgeen0bLTBjDp/roj7JKMGYHMGneVxmJYXqmLMmc423LbFaD1Szdgc4N/ry2EZ3GcPewVA
j3nZmrnPZmzjn28zME2DYoy4BmRCuRcZTJ84xfvaBe3ArkXvFyZP1w67GGqHyml7ql9ZKapgMKH8
mzMy4bhngWdrsVs+E9UU0MUbuWYhJVttgEuh3uD/zN3vjBpV4JDwl5Rlw/lZ87IccBuHcuk/MWxM
KR/cw4L+FfEXkhbewWvr0BobgGCwRGdD894pdSqAfg4zFgtrx87CwthCD/JeNDdtxBHPt2zLSjKM
z4cOiFzC/CceWvMNf/vwRF7XBk2U7i0Uwc/Qn9FJSha7nQALd9MWVqQZkez8DHejb6h+hjyIBPjL
NGhOmnAwKJscln+Og10FVTao6i0kRvy9ZwaykUCC/CzdL6l/1JYltUuGg1ZmUpGB6LVPzdCLlf3Y
MeOVdCI4jht0Qe/xi3gP03WBaqEOD3MtZEpOm0ygPUUyg+CIxDHZAPp+CH6hoKh/uARj4ZZBCGaE
Dbw9TkMWF+B4UGFNPDt2r1aNOsFsXS6gRQ9m49eooOpAiGVDGZMWzVPdAY6Xog/Qv8l3OIzlnMLn
h1PtGhVHj1p78g9OZuJWFKSc9wp7J78Dw90dO3bFmNbBBVO3iqmdR5jEhVN2JkduxVQ2FmgRLw+O
SId117cn3zdskWJuFZcfmjHf5lHOfSQl15D2k8bXOsVYCvwf9QRmC3CWpZrbDkmNvw5PClMf/XV8
8znU3grnAiCi1ICxiQ+ZdhxugDFCkRzGKFl+jIrFZO9lkuN6fwLKHt/ooa9wZ1qZxBW5+Ze8nZKX
wwu/WH0u7pr4E6MZbCnNtnnjWC+jcZPjGT2QDiqAIRJ+/et3M4caMjrz6CWcRuqbII+5yL2RU1cb
3zvakzd8wWgwditv8K9Bq8DNz4KX6zWuHxNH6WYNCVBr7JhzAHDX6yBZ7f0JW1YZMpNM+kUMlV15
KFIvZT4YIhRMvHvBn1+wYmO3wHs/bU4GJQgxwTiAWyyO7toZltdzcQuCoWtdYhOJhIjZ/PIogHfs
Jq05c8q64nOvxlGmKBxC5jwb4uPH9xKnTforkjWddar6HekZKRYUphfzVm/OOWPFjQEvja+Wt37d
K6+X40WmyICafaa3QvU02oY2oiQbnPvOMynvWxf+aXGue9tvPOtgfljYfHa0FcPNR8XtUz9JFfYW
/vsCABRuqs1IH7tY87v3F8yg+gEo/3UN1KC6G8pBJweC6hY8PD5ejWsS1Ap8iKl09xGOZlDwKrnI
o9cqYdOKBI5rwj339+JoQryXbYr8/cdc0PnQXBQClPPDOxMAuYwYwbVqavWCDDR3lgXDdoaTVc9U
D2n2sVFIFDY9vUpkkc66iJNFVAfjVXiiMpeF73MJLgEGC1xrs6VSAWlTcW1J2/mVo2nz/Hkh7650
uVfSvS5deLYjVGTNrvtgM4f6S7wL4lmP/JBPKI4l9k/NtvXsksJmwFcWBoSKIdu+nfcaoNlPE+nH
+uzlLkasCyFQ0Zbug9aJxXZF0n9KUqiEi/q0ULNdG577rF3+NdrcWyiaoVFRltN0bJxc6u+LM0WN
Bm2YVu7203vkCFTSm9HIxMezjkhEGNLCrK4CDNhcAZcjH0D6MIy9gJ6LbYGt11yBmytnVXu4MsW3
UkGIjfLOXVOzdBBXWeQTVzF4uJkn2McbdWCLSwOHOpx9bgwN04us4nDP2c9QMOQCSClxljdhqf+q
RrskTex6V25ZYilB7TGOgCVGcXJ2M/i7h0r67/3dpvIEtODunMWJ3bZM/8VoC4LOEkW05qJ7joNZ
cIkTmzNC4b+rj82AmmyPCyHZhxaVIiwW2Pn21fCg1THLrulH2YN5mFMV2R9V6Vhha/YnANblszkE
YT3KcYUQpZrYLpObv0zWaql1niGT0lZvrfsEqXeZE+hzPMFQYgT0PcfPGyJ3mXmt2Mpdg+D5GrjD
XGk8nBoom8nbT6DmbPNk7CA9/EluGpgCXyEOc5oBT455ppWlf0HL4MqzBoqdJXgL55pWqoHXKFfW
RdUW5u7MXTwyFGFPrf2VWKSSSRJT+aj5jF+aYL8c6CYLpmjGwzQ51HLTzTKaJUqQ3DQRAP1dAVzJ
ziFmr4hftuJJIaC0j8kUVYaGiqfJHPuJwfd8rr7BHxS3/5FY6ppLJ66novH9uAz88VQyqOAaKFgr
XRiocQ4CuHCXxiYmzw+Wxazu6BQizXb1z4rQ6/8pAtd2a59hiFrO66AGHRecwCQn76k0eHNPEDSK
XZzaCNSwfcSWCq8xVzYdBOGNh9pug61PmiOZ3TU7xt8qjGNaNK8rGUFFMCEHcRUlNEm+eRtRuCQm
TDVQxMGN565Gx0470bRRjh7PxxfvNZBkdlqI2d/w6I4ckp56lQFNwB5vvilxDoKevj4Tk6Y3XFBI
7d56JQOv2mfK5oo+vgrTYamGTtkvV5ZmczmFNZZLNKRIzJ7G3Dwn1LOizJKKEjaY3kTsOKTVaau7
7jHhi5uKyyC4nGo8W9P0ETkF0M8R5rPzxiv8PpyLrymSMx5HDlC8AAjIk1dIrVJiZqV67LEs1i81
f3oT3YXFF0rZkERo4/ZjqroymtUDUcLGWFqjImjD0gJkpHjDY+4HPelLXd10E1SP4fKDMnf/V1/u
DJGsp9pTJri9W39wffsyNSCAnY5/7LQcrNRt9ptOSX/SZI6JaE/qabsCWQWtv6sd0091yUkbzyGe
4447MQjfqX0372MuCXaIU57P0JTrxgx1BLFN7Zs8Wus4bOrgkMi7fICtW5XkxhZBSJ6QRP+irIAe
zVgi1ZrbZKwaP2bprC3Q4XBng8ozFZMYS+CAdWiinMeA0+xauYpDjWj1t/fzpX51D4GNY7Fe/AQ5
qPfNzyoNTKMoeqM/Legn8JFwwxmlP7wqfBL6f+07qlI4S0rm2VBXYyr9Zvh+gp5pGcuklu6KKwzo
qfaK6dFW25daFEzFZ56WmrdRyeGC/zi1kViYcQOJPBQrva96ECaJVvri9NBqQWjvavmdNZcm02KS
CVNWdOvLsjGdb5GKEt2Z3/gKm9qszOLnD296ghaDFV3AeRVmd+2qHc872WYFBklpfz42kSYsUCI/
DBNGsFnHHAU/UAKd2+FiHPYYSurGzCOLIeHxC8KFwEYKWjGkgz77ZaNo6OUTdB3Bu8LSkcenqea4
RRfNmUMBtbQozaK3aYptBtK3kOloywf0KDe26owCddfXgouJTec6prJlXVSA7sQbUwr0CD+ulT7C
zRcZh++yDReS4G8L9M5Qq8PvI7aF2fDv/2oezq+TmuOeG7JrgRhDtyFa/CGLCOJHL4vj+EzwO8ea
7ngNowG1dTjZt/spKpttQLEQuX0H1uditllH4ut1T5z1COBbxPbO5PBYBkeg3fsbhAWml00uQhTi
ytK5ifUb8WmCowMXj09uvOBxwi43xQVNEWSFKbYjF3meG4zQBkZ9LUFurKYKu7A3vEovPM8vLE43
dCfSLypYq5T6ZQhIsSo77aSbkofy3RTZUSn7IgxQdUCYz85pfXKJ0SSJbTI48o1ixZcJC6EQG7u1
TT67M0DcMIw2zYkqgP+SqDjjbxonz1Gsvn5TQQxg5peQuYq4tj7OKqegiYMltqQxJc9rLabIiqTD
AJhpmcCis+rg4HYT4TyPqXjfpUXw/5NUtCd0BaagIDuCazXMJJAdsYuJiay14VqWC/q64pPYti8A
4CQxnI2qyO9LyMtb9diQyxeoZiOJ2ArZeMNq3rzK/nEj20r3Z8t5XpFuq+1oTDN6EjEqmCQXbm1W
ShO4rT5aQr6PKqdfrW0jnBzYYkZ841NRxTm2rGQr62pXIPvls1327ApGd4j0ktnU2G8S+HED0qG8
dUDbreneXAVxLxG8/LnFS8/SQ31ZgzIfF1FiGig5W3eas6r1tTidA0VE+RyFn31YVByMzBXazFd2
/yIItiKdUyY9iDWRY9hoordvFfXrmug6GKN8ZrtzBLZ5Eb46SENpTkC+oxq9UVptxhfS5HTmxnK+
wA5DIanfk/2Fzzl2W4xddFYNtn08EIJBcipioWwljAx2OVCd6CKNNy7m/v3R9F/yFew7lHy1uKr/
SVAF5ANqOVR219Hd6z08a0bA5n8MEzm/J0Lp7YFXBcPqFj3Ohdm3G11cugwz2QpeZdjZiN3+BQFM
iuYcZHxRF2WtS6AwPAHABhJ3Xt1avZj541c/Y8gYXZ32W2zl/cU7tV/TAEtPNDvzKbiomm0Uoy40
9pWcOjK5PC+CdYMKicfsraJ2OEsWvQpRjWK0LbEGCxoGCHFMtGRYYivimRAsteUnGJfIc32LBbGT
ImRQHttYSCv2E14uW1bkD+9vPaoXSDQlUkpvuzYHhmxzq6321EaVSSEJyofk2sqCVDx6eD+TKjzJ
EIeS55l7YCbCLDA4875oAinwdWCUM6Xb6iYtodjxrbGIVFJVaEcNLCpAnBSdF6esxKrkUBRNybu8
SjHznpgpqghNm6itL4wRab2M8UKIbLGlf3rca+LVE0rZt8NMSFTT/yK/jUnH1uqCNhtrIhlbU10Z
CiEcvW+gi4573Cno23m40Up2wFoR3Iqk7zJXRH52umfwFkln9l5UOjTtM7pL/DYJmJnciuvilhsH
J3W+7nOWzQG7OWsYtuZbj7gvEPN+eF/lXI728ys3E2UJla0ZtUytX/42EIT+IFHJvtzD6yB4bJa4
azkYAFkNoDfF6T8LCyJKcR2W52rJluivSfgUL6vXPer1iAty6jPuTYW1CGXgSimSSkVZiH9n4xSP
a22mKAy/YVK+9M6YOHMJqNt+JjQVB0pmBPY5Uag7oXZU/jgErrxeaLfAajJieS5slnPOfFtyQVVV
12g+IjvrvhjVm4gnm26Id+ZmukDd5YsS9X0l0oSZl8jcK5tyTJSuiyquQrJqBVe8PeHJU5V0T4cj
rR6imrx/EwbXo6dtReiZOQWCh3MPDWBKMTUklnkS7Ult32botem0O47Cf8K6VA1ONWxkIAQb5N4A
/pVTN2AEgwHPD8uPm0U2uJSvAUOZ55T5kGobCp2M6tS6uFjMQ1ujLwzvuUDDiFMC3MRTJyK7XKUu
GW+sCmywioc1NQnsBg0RPkhEDhDLpOtjSPI5odIyAoqUemf/YsCIabEpazmwJVZPu/nAWv0+o1xo
7ZenicbZUuXSoi+To2TmKu2VeEMCYH5vsOVrZW8uIKsd+m5VbQTtCSMZ+jtDvu2eWoz41/vGfQ4X
U5p7q279jYd742FrFy17yf4jVH2BC2IVhaY0cAH99GVvQ8tAZJKQt/xOvpH9229Ue5l4/PqZWyJ5
4+l01V84rMSuN5HLpbFBvM/KCM5+OdGRPfmXATFlWuwahoOFZjb/s39Ws1Pc1NU/+x05rka0CcMt
XghDE9M31iL3g85Y+bVvSHXrYJ0MiSSvcaBk9HlOUaXTzJaIJROSjH2DgxjB6wheOt7jiLeGCvXN
EvQiNhT7cH2/8QugdMb0t6sQJYKValhU3aseE0vwI+3KmYXo3ifKWLLakUCxpJW/miHQz2d3LNDX
A/0SeVsN77vrXa4gJDnCnnPoiwGLzY4cgEhteNach9Tf4786rYgP6OX5daDkpvyNBsprVEl2upag
owkrJG3+MOexNpK8k/1dX3c5jRQt0H7NDvG9gMb7R8SYQa5CtTovaAXSWjqtCBTURiwWKh+QErzv
6YNjdN6Jsgy/3hBwyxdiZRC3DCKorPIrZEgwJVIkHCmVNTwv+8lvR+ZaPHpketlU+wjaug3r3nUv
wHXiJSv5RcPDQ9UBoMyzmtsv1Wc5LksCsKhaFaQBVPnS1LRAzhhAmGJ3loT9VhdBp0KjEnBca0s2
TqW8hADFDkshkyFF0mseFOnoYNtWLoJtgctkDd6qGyrwZmzz6S/Kr0GDr0a3sN/IQUTOLnJ5pNZ1
2rxrhl1G/sH4yJ6kDb+eh3qoNpydkBzTaE7GOjLYUwMgZ6K83GKlDRPOePiH2+a8D5huPKKLSG8F
vsDjVDBBsT+MHDKgScN2wagz3gQ2e1MIE0l/XktyTSoDQ3PdDHbC/SReaeqMP1VAwoQhMRMCJ7Oe
DmI6EfTMN9OewwDFaH5qnVPk8Rjglr+eTVIcXXAlw+53g5AD0rDmrtVtZLyf+vCil34bot9KlQUZ
jvK02PZkxK5AKoRtvzyaGlTB15/2RY8nz890KRNS+QjuXfewG6Bd+OHk9ROqbGpSu6nzw+d01lLI
sCa3R/Xlq8SDONpEqjhbKq81Km7M2QvWGR8swekuyMcxMPDMtdmclVZbLL0AwLJFiq9F+05Xm57N
6/Qpxb3+CDk28t3tH/xzzLkuwueBsy1orU+Cc4c7PuK8wX6mXRhDATDp3BNxe/zl/s2nAAFvTmjw
alaXdqMh/j5u+LYQC7dXz9vnXKD0sx+mHJVemKWlkGad1/50cM3BrwH/OcLJq0052afr5RGZKM5I
/08ZOWkVpIGgQMygfbxS/fFUpSo2duPdJMmrRcKTvDLTsrdLvwx8Umvzm/Q5n8jbTazYwzshjny4
Sx9JuDvMtCyLSPNi9BYEjG7gCoY2Ne157rVTi2YOH2c+bCq73a4ejRwSFR4gnOzOqpBzDTf6t9Fk
AP6Wkm7/Y/C/+3mezcK32Jv2PBQS0gP3ArcUK0Kcyc2Kwrm9CFTXn5hZoGyeXuZ9Rc1JCAV+kqaW
HGk7MIkEAytGDC9F2fWpwZh058hhQKwSLGppvR8WCoOimGVKPz0D3PFeAWfhXvIkjPUrV8iuGb3v
PZWMRegb9D9U8LPM2awV9ltA6ezf7MBSeTHMrdwfNF1i2U41rEzw/F6nyev9d9DHMKSplyeP0EJw
kXh7i/wiUc/E4PkOIi3pOx+WTCtfKSZniRtfZ41t27w+UgwYumCK77n+gSZQjx286WBdjTYTuSNH
uZmGXj0cCrcLedP2082F9qhXh7+JPxsFR5LVJ664ghHNwF9AqYY7VWJB5dSsCBnNFjt4+NbUrb7H
10fZtP79bzFho+0ARX8MkUuYEKEwG3PhdOD0fIsB3pQMTRDkeaJAH8sAfVNe91KXlE55bzls5u+m
ZDbMSMGHbU8liVXMmjCTw1r1UCm3dvdrpPlgY0X1NT9hDWn7tn1wGHX4WCvGe8Oq55cd8YWC1aUZ
rfjihY5C3w7X9eEuy12tjB3VjRGnZ2E+gVVZGkSrFhtRwiFnlxHQbRAfIvxp8oPCaLH6FUoZjo9d
ikzdtpePHCeRy0fRDrVB4JSgNUdP7TB6iGzXvUcudfTm3EnhtLlgLGhg5rvIIBE80dul7jmDfkml
h5ap81Q1LmpF+wS1V/YkQMabfGLXiFJq42l+1CtqukY2Z/ytOIL15ZHTi7S/dwTsuVQgnJpClIuJ
dvSzN9LchyNFVL8x7uFUBrU309gXcU1KV5nmvrRc+f7U7PtZ7kQuoNYIQLkSGWDYJFrgcptGs7Fq
RZkWe+SPHv1xr5c77AQcyCQ9pVnaHHz1jSXetd66+rK8GGb0YfqnX3c9yDpI5nokx8OmCjPUGaBN
w+ECv+AgW45puI0rQigL5IxDXtfRIYrmHnjW/tA4zQpIAP4NzT4xsUvuBX4R/l5fK9Yu1fP9jtP3
TumXxgylSOsyS7wPtPQjAfiWGaQGUaU9YVq5LuV7ms0lr7iRxJ+vy4fcVd0MZpt2wM+OJUcJm075
egNXqFut2ClYFevhu035w1L5rdN0QzkBw610lV8IdqY3Vj7m2T+KY553iYTToDpEZBEpJiwTh2Dc
G7HS98dTMrYIwgetuMulG3vUSKBM6xexz1LWBj4zozE6lKSddixlTM9caCWe5YnL/3SsOP5FV67d
3LnJXN35rqVgOZqDnece5UPbV7ay0KhUD+U1nxTgib835F3tJx+ZQKOUBlJwDuQk5uFGopGSaZEQ
vb0LDVstP2uj6d4ZpnMLS10jxVQT3HW5js2voyL4In7ZpGmoZQ8qXk37c3GLO5XD+tRgPbBXq3f1
0HLbZcJqLTYWUmldgxsRYERqzZwFinoG8epgqnqFwqjBWRtR1SDWRu11ZrZun7f4NS51vLasiz70
jjRWxVLP2PiwZ8mrEbRVciC3mOGFjkPiNz75jwUwd25gm3jQLxlDSDxk/sozkC1rrII5b+Xp611x
orc0qhx95pxQfJNjavYEKIKcN/j0PsNuPgZRplYG0zpK/q4SOq5ATsqSCOPobHZlT7oB+UA4X2gZ
1TFMPVi4N4NzaU4t1vh2R7Zpe1/OHrM4FnVDandyyn2sjB1+802ebncrvzqb8yuvejGSAQyZ10dK
dtpxNuuqzYQwrUUw6F2hL7LBgcFHdqxFPH6Ieg+bCv5jCFWEnOC2PcwYzAJXdPHDDM7GhnXeqTz0
lovFinUxWdPY5XRVAXwm459hAWZ5oDM6cYhC6y2yMqE80Ib+MAVPfhPmslQi+A0zEKJ69j6NRt93
4d+Hbk6Vl7tVYujFLJt7fmyiTB9VmIdoBQX/BSwp2/uHqrXQCpD7mEKzVbYOt+swaxeYs2zyoOF8
kOjXSdsILqP6QFfAS4el7NuB2OSnPjO6Un8adfhtC4mmmzjisDKe8PdzX9CPkQXqsrc2VsMFRM6P
cKD/LMxwOlG35scH3vcX1blJdn8Bkduws17LUeX2GD8yipMlsK9KG1kZkqc0j8BK/Emby02Bx7rj
IkoKjal/VRqwNjhr3uza0uf/l7E33WhJOCyoFQoIdPKq4/4RzTg6PwSUE985O1TvCqxKzHFFpQPW
XskcWfE9fzmXcBX5OgPXFH26lXGpjR8fCaAScCuDIn4HvJNKns/m07yFNanxYjlL2EjlzKLDeUAC
RlSNYLa2xmg2ieo1tDosdOomZBZ5MIz1Kz5zLmNRd/5fO244CeNceO8MoeY1bGaBxZP0qcSXrE/m
Dv1vNI/fhLjYvaq57CXZzJ9cMJ+45sKbNz+esZ4UJpQqeZrREkhncuXmy0tiNVZvRs7H+1XFaa8N
mPqhmpzzL/zTWcsYbi5BjqDaAkJOvIHMviCAjYLjIGdjwwr+m57I3V8jCO1JLyuhe+MWyoL3Djiy
jyFR6CZkl4XFme404j9dwqYGphqNOYy5us24Ab3nomxyuFiuK403uLpjV5rGPY3ksp5H5Olc74G+
0swjZcuwD4mQfXW9XDHVEjZbVTULV0jzlBoOnzTDJzLo/xIqX2Cu/qGmCBhh4uXDzD5JotcgiINH
bk31j06CzewnkNCEoadsNG0TzxuJrl7AVYNEkOMV0dXpvVR/SNW561y5XEbFBjJEWz9wsbgYW/RU
NPX2e0WYsszk67PkoKeYImONkftJ9T082dQ4BNBQ68KOjtLvHuJTPeNxFNyYIna47QUSvC9rntic
OU63AKvTRHVQ1QLKhujsEeSqSRzWmgYdQ91A1b1lzllDs+LKozbs6TbrKgMyxbt85hLrUa22M5Us
KG1qCKhQ4ZnabvVj2VbRyzrEXKx36EC8080B2VNjkwxu9JUExZpUe2NIKF1rYzFb5r/h86OaXZgn
mkfN5O/NfuXCgBpIZ2Uc0O1CtBd6HC+tCF0rL887SPTWJNmpI4a6o9J3SCFhVMQYfGaowDtAO1Vq
ZXE1vwpfLwo6ahupEUR5jLZwnreD+9Tk8HQDhWIle3HVWcHNGgRgiFxPnL3digsbBLR/4ajUIFdG
M1kPdJSG27E2+aMLdG/5jq4N2qSyiA8w93FHO56sLLP1NLGr7/7JOjjim+Ih/wan28VEoJKmYVDc
y3CnKp3s26Q2nhlnFWzWy1ZV3BVwpoyudYkKhEJ6uk9qU9VED52/FqyHIRrp0gxQRhasYkkGFj9O
Gzsnp7rtuHOFTboU9gb2vyySBGzPkMQ/LF87CeYVYhUyu85Ls7V7/JiC8ehxMu/m2aJwDqwTsU2F
fR/iGQog845lVVVxMkdNuqhQC3wuVdkh9LkLjv5g+OuCXQaH95Eh/SfFqSLiwpTzjGdSMV1VV7Z2
zNthhtyvr11XqU14JNsY4AviJ+YcCzt/3RDEE84Qq1WVUlEZgr5epkVz+f5GqENvoUcfCTeGUZvQ
oJGiuCozYxOEZkXHE98ACEezc3RUQjsl5Jq+QnKfET75v1ixZ202QwV+SR9qXqFXpUd4r0PSlIPs
X/qE1fqUPLtoGOunazMV3pFgvuu95YTLgmH1+Tx0G+KF6kVUzLXh8+sW/FTYmNZ0TOBTRgY3RDnQ
UMdZMbi7g1tUg4o76/v82rTkjmonQHzIJl7rJ8d1YNNdm5nSGb52WFPod47GG5qtJ/b7IlDW/tvN
zZuuM16ZeXiQ1VLmsmPAiehRpeoXdG6qKQvpPhZVgFqgJtgldDA7BVfQwJwpGSnIl6U5aYoKYXGM
+/+38ksmNgDSLBpZf4q9M/Pk3tl1OgFzqfu/YgCRXS5ZUa0yafzVL5wEEHwn5xBQHh8gIoa1+72K
SdC5eHmUnIKfULDCQpd7GQnC8miJqfYEuMbOap1xKiKvbxr6zoeSYDBC1fj8KGORAsAHtr9Jx07C
CNSLVvTvr8lnnm2piL33m9Iue+0pZrwMVnaeCt/z6SuHpCeY0bO2G2DvWefgeHNcgi5JzjF+pAgW
b/l7EC99hYb0UOaEWQ92C1ukHtmAvy+nWyYSg3Kk5XSH4HTSJXvgCgQpyXEXbngoUwhzfXOPDgiH
bcxaSjhAhaHgTrc2b5DyTy7P+x7UV4CH6IqfJcEIexqyOiadWyJ8yjz0j+ec8X34tKbi69mScvGj
Gy8MYG3eNTsJJfSYM2mepdLmi91w57jZFLFEZ0hy7dLveoq+lU5uKN9ZBABRHexldN7EeDIBGLXi
pTQn2QSkMHGyFqgAdSygo5+TWT+7utH0Ke2Vqc3uS2nRuIGJ3Jn3yCZ2LeCQR5i+mxCj3NxNTJlb
NuRGYBZSWK6s4U4NAqYo+S10IDHLqZH/l78r+/Auw3LHJrXOVqiNAEuVHrLhRCLGeWoX4zxzDIzo
W9rDAiPgX5s9i5O7j03NomACJ/uUeBcewgYYNepYoxUfm2F2BiWoZ07aB0H5Q8QQc1wWCzwFoZpV
cH7iI8FNreEeJmiTwc2/3S/6n+byAZl6Wy1y6PTMxUYxs4RmmbMkul2HKCG3R76VKTJbxG0dLGAO
Ore2VA+f1sFQ6B3uqCAC8U1vU5v2ZcblbP/bead1xGW9ORmX9jfp3+95uONybbDBweqWJcbeP+4c
FKUqoTin6kkXWr+Mw8i0hwJbbNH159JG7lbpkflGpgITIfh+mCWOhnQj7HdahfTF5Q39+Mrr/61a
U5BxiDfV97FzGs2IzY+KDcRI7Q+VRqWbqUkhfdajcMXPds2i1QnV/ACTS0ybPB9RoshTtsFww2fV
5JHey7Lyy3Da2WzRzM1xfQJBTYtHGhPZPnMiHxkj3ojGfjMERVL7F4I8LJSPSCZAsx7A59jWNYzZ
Z7UqVIr3y/sX57C7rJptbgUOfk9TaJUfkBQXfvUAYwZj6a519bm2SUuL4GUOTmb6LlzkXdKs7lGt
VMZz31mjJD8k7b9MrJxehJiEWRj5U+jVKPRFoZGGdZk2xcQqUyFt9vr1W+0SHxSDQpL1DBoZEjGx
wCfZnwNRG1YLpLtmFr3smQdmbWP7w8GP1lhAHV8a3x5eXWSt5Mmai0XnykNdMsAOvDIefcLHwwdu
BbEM/7CWwtFAktz2rfc3s/yUYgEx1af4bxBjYrXJU6H9AHuSClMR99yf310+yuF6XHsCr66UxRsW
8CscnIosUh08sYROYckyAdo5VmgQHDvt6q0wo0u5QsuphFlKMtqReBtEJfjYBo56PxW30uJJBkA8
LZQOR3Zv4zuzBBRSJnoxosihqt538DXsvJ9YsCgGhOv6HNuqG7JKv66sFtVTelU7XP8xSn4gW5Um
NPPwEqospwKGQvNn5nXm7TB7jMGUhvPm+xilIWfSXisYcFosXiiHEVGTR4wrsaPeEeoYW9yx4i38
cujAHdsnUfJgSv/i1DHaY4uWiviDW7dMnsDtBhBNADOYSUoz2jPUqs0PO6Lypmr6awyfuaPMZWui
NMG/6XaTMW+w9rPIs7Vc6+fhdzN1UWzH3GhQ0p+kK/vqZWzxITbeP8x9gQ0J7s5u16vYvjmIuJHy
ZbyHM/72Vr64yWax0jK4lqEb1e70JrRLtTrut9uixPgKsqZJLFQ7olhrVUe/tWzHYUWVromSPjl5
IEi4QOCJjTLlOdNm4xXBuzcOg2zzh+6C+Gj5cslhD15IPvw3EhK49Wua1XXleZjF/6ry24z6BEjq
nl0sVLA9Fzhh0ITM5+5qkO3G6DcjVvTYkjv6wfYTv0zYNi8GOtOEHt0u0znNZM2dnmi9x1OWFmJG
cT8nwy9xCETTK5m+XfxXuOypGZhPwZZMjyoYuBMmHD5897b5Mkb79IV9dxL4YEthgZoqjx813vZI
ikao7IMbzjB0o9PTR1/t5QusG/wgoy5SrF8Sho7ZWq07Ql60jluScZJkg04WzJ96QAB8Y+gk8IuA
3W3xKBdn1OqP50lu7UgwJLj2kbUBpBjE7rGCxTjUhedWurF/0tU647nrj23n7qmRSRd6ClhOx8Ef
DGCL9A4PDF46RREbvhr2TiMz8VbDIcgn6oamQECQIUkHr1xZun4LJo9LblRwuk/dKka6JoDqrxQV
I0uMf30vf5OcWSbZIHO2h84pKrm6VOjYEiLxKmtJPgqSZLaTjdrCRfjhrv11U7Mi709MG/u2Fe4j
J+U2ZMc3SS5xf/LbjA/bXxaaBRZyOhD+BJePb+tdRhqFYeSNV3rc4sh5qR7vuuXe+WJN5+Ww2w4w
jGdJd0S1ay/x/MKuZSKb5+xvfg5DDtBHrxCtU2noul1nnuBX3v2T1HfPVTp2yPhkAWNpH1z8j9vS
lPzsOwBF2T36t5k79DOC3QJx1h2Am9j1ahzUzhcWEmVVi4gpHRgpFqpsc8hMXKbQljqcLRzjDjQ8
ZYql1sdY1VmLlVlZoBdfOFDWI0tbysI47BqU/beFdBsnAUVuTqoTfSRYmFEX2YRXka0fV0kklQfo
Cqz+5KY8wmcvONggBrCLOsIV7+sfYMWRBQA9MJR/PS9JFQi7O85sPWJzRZrUtkuAdvkt4seM9SLa
zXWic+4/ZXKUugSVyn6MxpJ25sJvAIfQiWno5HkK1bSHGr0uDJczHV85+Y0TYIDf2uWpfesarEP9
+ApvIEBM/RvEmK/Y3YLoSdHhwZrV0dmDoh4rzrBw9OEB1dAxxYW+f9mDfN5/mxdtIEo5vo/HQ0zw
+jzlqOlO48u5kpWFgH1HbwX7QjhIsT9Yjwc9Q5Q61nznypEAXYjTVsTslwrTjaxQ4V95Drft0Dik
l9QBDoh7X9C7SlJfG4lWohSkQgECqMrNOA94qBRsAsZe3LidbNF27oQR/XSII+yF4nHZNxlBScRi
zUqIflevNpTs8mNWBFVusqanoCJ4vUjs9yfoM8kpOuJaIo5J3HGAkZLveNZhuMIZw0jTbKiyimzp
O41UGYIlX4rgZfRts4fFE+a88xqVNlbJFD5vu3lsp1hNqOPsZ7+y0yLkmfoKW4OmVxOsHj6Pmif9
5zBg/q3hdi6htyPV/96eyeoENCeAEhhL0M0bzWlvX8HXqwQseHQ+zSfnP7c0Kyqxkog130Rsx/UF
/BT0uHM71h8pTZ4IAHSH2YlRpaiOizvXnXQcSaWmROap/X0naA4FK+Y4wb7C9OYZv6X1N4Q762J7
wwOdN+0dysxoDsr2dUpZ5ws3lW4vAqy6gxecCOd8ffcrqwyyv7td6LxptzdADXXYB16HJsWduyQ1
TTNAjeGdGKKFEAALcsgVvYSJavxT/fYN0CLxInofm2h9xx+BhuUia3XWNP8Bhhlsv1dEbt7qlgyb
jT0RlUtlUaH7LZLjW8INy3ikWM1+mk5u4o3R90v3pVz0uVRkOwCm5z/aXv8s7CNrufvk3nH7FZqg
D37ixYRdIre7cyX2rh2ck+jEkv5Zoc+2JpU+ibqdoaQBxn86anbvaNzRCEnVvkrvdebsD7XQ//ZU
mG1dgPa3WeHivBAp5gKFe1uyt7yIEg4Ay6/xj03JCQJORZmRno9YY0Cw53i5U1/gx9GLoKe/NVTb
vyBqIOLwO0yWq8X+bDZdsbpshXXJtsodWhtzjLKzIaBS5btkAtNg+7zMWYLONVOrHKr65jZ28dkB
rm7YvMV4NEjsQgqQn2dR9/FFzzAyKGdBtMAica1UvfPJoLzj7KxsvVgTvrC3tipRI5WI7Q1QgNpz
753wgkLKznhjyvZoOSprEjoLlOGfxbVbIppzp23c+kxSR8nQL3qtQKYFHUwTq+JSv3gWX0RqqK+o
o7IdgfVO/N6h3c8tKuSYtdPoiQj5rSmZfzqzHYy/nsK/O2AmPngdYkhnPZoyab3T1uN9zFaaKN/v
lkPZQCe61QG0a/dUh0RU9LB0ZrPl9LEebtVpWv0/SPJS6Y/1bOLrBfWKM6Kq/ZV6KDwZ9lSeiKrI
5pz5EleVqa5q6KIF5FMczGgxEc7x+5ZoQcDgTsfglbOv4ea2qUbMpWqfdwIThWRVAaioc+RbhD4u
cTwr31Dgq2PQVxjfu9oOgm+X0fvbVcP/xfIDFbeHGBZlVAPeR11muYFF2eIj2eMCnK4uDADENePl
X9a8nTbq5uxuI2IKboTpe0IF/mE4qh460ZkLaYyHsVcRmdXZaPccA2eo1x4vsWwZ1f0VGtnQmXRn
NH8zFKgNWQLXJolL5mdP87SB5Y4lv6dWUheFU9lqLOv/J6dwswOoF7qAWPHhzwH9eIi7C8Ni9W9h
dy1lGvkcBadbvQmRU7n+U8e6IfUQg/Sjni9cdvUDVSbVd+FOQjwYoyX3XEqGNZCMb9gA0vLb/XFg
H3IOfU98WtgMNvKuuQOIEwbozKG1L1qHEETi5EGJKJpbiUQj5ZlQImws37MTeIp2mBM7L8Ow3+bx
MO43PAn1D4D03d1+nGB0YavoF8AtA1rZSRALM6vyhtdF5BqIHdE90Yv/DWNELVcwVKfU/cNHTLX0
cGt/o2LOG88BES7ohsq9IBGQWxeojWfulVORhRkSHkaX/GVojVeao8usLoe6kAYstp9yREPmR0so
HYDEA1JISKumbUedJ9eaEEvT7pNDr5rjsX/xYSCjhZHvPFb84XI46JD7Bz9XpreceDoXpIkF7f4W
UR+3mmS49cpvoLv0cqxtRscVBZn1QPn0KHz2IOwHE1PnTM5/qtAQ5J6ez5s0cWOo9Ea12EULKQQh
aXyXd6z4pNgN+kW+ep1AnXicElP8kgDpkclA55O816l+cFZND7VIJNqg68zkEF+A+vuQw/971zTH
nzBiP2gdaZwkigTq4bAyHl4ojKQqciqCCzK6regYc1HgToq0o7vqv8g6WXu4axljL7GGe1O4eXdt
4beUflyUDiSyT5zdFb5MIURYXqHcFCP1Ot2aXSrCzKT18zy9lmpwuld2HQ1gg+ChtBl6XfurLMYh
Ym+u2pAhCsJYQH9sizeEh2nSkS71bzFdFpS686JDXD4+OLzrTCX3KI2UTwHpnq7HLK7vcVn9GIgU
Q3zEU1JPQvLaHoi4NzBVAjYxKDeCk8+4YldpImlp+rfm1+T8wH2vsTD9PkOyhtsOSysUrGJ++q52
/eBKGvGuUORgOFmF3Ok9v05uQTX+LD550up1dDLN7CKC1u/YZxeMMJvLBwf1zrO/H6AYoNrUbY0g
b6E3In5wQhJba2wkZuklf18cGTeTJpxGsXzLYQiLbO2GLhSr3aqaeOnrVbjSnqFY70u/pOzxUh57
4ux45vjQ7LAOcjnGh/hJoblgHHSLemAqq3+BpOxMMa/QvLqBpJajpMz8BaHlLk6KrmTgnrO8Ka5R
dpepHPqneNhHaMJhLPHfPAMnFCVaVo4Luu26T1z2UXssU0q8Isj7JeuBU2WmwKIPJUgaxbYAnyoR
xZuzwhkkBRNJDuraAIoSqSmWPc9vzq/7wT582p/W4kMyo0D3yEJ1lBhFyFgkP9LDzpPCAgzw7ymk
3iFdZTCSJyz7Z0bP5JTGJn1ThMsNOfRXpgOlweiSo172ndheNF3Uv+ZrY58UXT8TSJVhkn6xUD0R
kFsKHi6ECsRWliVRO6aJJA3gfLt1aeKBZ6RJLSxhX3UH6f7TwF4nSDh19Rkp6DqvZYcUnFq1gO7J
FJzkkAdYhMlEvymQ31+Br/0aaqMjVXKkaXCTdfeVS7kuFgMnilavsutcUAVWm6JjerYpJRyL5hem
pR5fu9nFQyRiI7gKub1gdJWLbQVijw+nk540LfHwjTRlo4/3m9vmqs+C80RnhUs5XfDkBh/NgmBm
LAMjpvlJ2u4LbhNz/5T+HR1Ren1ZmGJoF4d25a3bxnsIr0X4zyo/IFCkxDzaz7wm8Y10gfqNU9vc
NcG4q1wkKHmOfplOQC9ZjB57pDZ7o8NFf34WasNEYHigONjmbg1Vwa1q9kjUm6Uu1F+zjmgM14hx
SgrrtzYUscEXyYO+Lfyw6+qd9fR8nBNhhob4/cM9cO7vIUqDfsCWTJ6uStDsY0D6/TEMoJ1rHvnY
D9zF+NeW+Ly6WoDX+XeTuk6B2+OjNXtUJ1IFWzwrRjkq6JFOwQo4K85azWQTS/KAvCT19P/t4Hip
FvHDglaL+vm8FRnO66fNZ1dOeO3s9syGdlzLZW+ucJqeBD7SINs7fZdKMJW3BbFQ6GwDsAfjdNKg
WEKQ6qG67B6SlDCfu75UGaOo5TmTslrAgNFVh9HHq6aKdcwOOsb+VAJHgt6H+KeiHLbuc5NeUroM
XM4Cv+nK4OdxAgJf3h/+ZMMSVlf/lqOtsg4zGorfV7heJBvjsDkgTa1YpDDt39HFDE0j1RISQ5dC
B3B361p7/DrMO8dFH9kQS29vAuw8s5GXdXBcXyTgYR43BAJ4ywEcRlsEb2rXqaM8TkM0TeqU7P6O
E69r7cHiyOppooNVl1Br49aT7ULKDtHbBoD7+ZnvfDoFxkS5CKJ3Yy+Zzdk34SMf5OhqrlepIenB
rpqP/5K4kcFr/iFXnQ7YpM9uNi03dOI2F5yuRMtD/Cfr1/W+0U+4AUamU/rfoBmVavidlnjGF0XP
PdaXNnBOS9Ipg3cuKnYe2+HuUDbOseLtrQjOAIXYY7GAskb2ccYJ146oyPQieNpBZhtjgcX+Sjup
99uV40wu+ytq2FUkFfm+xYe0cOmbutIaZzev4FDhnnlDD2QJ6tPHRAlHPaCiIFwnjtpTxTxZswRD
s6nUnTrXIw4bw420+v5giafO7zAb9e+Cqkdqk0601A707GtFdRRPWdYPewB7w7meRNRBuwM1iFqf
e5nWlN1FbmF76LvvxjDtmtwQkL/JKFLtvpraLW9vxs7K6D2DBO+VFpmqyZ8RuIsZicxP+kXLWiUx
j8kE11ijE7J5ZIJc4EPYdpDlKHlBMmfjB13rLm/Z+o9PxDRwcSJMFQMQ+YlvoNy0/XIkCIPLx6z+
dFpBZO1u7vFsB2UxNYC664sUY4cBrC2LOi0OS8yMngIJm+P2Y0cdZS3XOGrCOBY89nbU9iIoFjsy
p88szkrhoPz7ZtPuavHzNQKvZoE4hUPm2t+t0gE2dogMzeHLrfYuaGRAHOlS4I8wOynQWlZLWfKx
HXCybALoX68L7Oro/NbABeDLIAnW0lIgHQtGf73ipNEM+bZzSKDNnicFrzkdXWh64KJ+fDuniAa0
CEKGuUlXbLf4xo3Vh6qqFttbA7/sh2ejPfgqd38v9dQ6L3Pfxf6MsVpSkrBSL00iBIGvXv+nPsrZ
g/q7HbPKcEfcnS9KJM+SJnVF1YiSmwobn+yIvu4mwbCiHVMIaOzLKbifnZnKYAODvjB+4kZQavqY
uK89uGctIImrlXpa73J1h1rFDjiCsPnpBpYw8wOJPM2DTfkQ+2k/xyV2HT+T9mtGGg5Tb/6HxWU1
Cmhapa/aJ+jD2JjIq3kAHBRgDdfXTHr2Ccb4olHJK2ikF96iuZAyWZmN5Je6MFk/baTV8i9fHx8R
RNf1oIaeLbZ5l4xSLAEr7xae/2G9DedL8GZq3Mp3B+UhNmx3bo7zqshV84GHJ64tm0Ulja1GgnNW
pMBFwIyKCfu0PisWyuDdL1X7vki3dhzImvmUQCmCwbLHrVk3p0Kj+T98rBUHEaeQBYzqF4cxtfZ/
BwvEEbgB456u3zd7Tz1Zyn/skIorjasEG8YVQkm0sk0FB3BwPYF6GtaIkqTsoklzteQiJIWQpn5C
DWB6Xp44bVKhdbUi48npJZbzqInSF22r7yd+V/msF1zUuo2kGJYRVinq5p3y2vkWMsefi3JbObWy
tOaNucxwliBOZ4x0u6BNxRLOxqS9H4CbJctJr5ay1o0s8K02JPudjj/0F75WOK/zzJuS24AxgzZe
8UAFodCBkJjBiJCCDtxfWEmZSCKvQYR2mwdhCOc+z1oL+zxCA17g+TXu8OIRpjabszaablujK0AX
U6CBHkx7YJERKNph1LikDxrGKv1mm4eQAsMuzgpfkXvZswyRHjgxqSazBsn4FOUwQXjlXxFFf904
iXqM/hJkscM7yul6QFlUXIVBt69No82VNXoVAOKcL96GjOegESyzchdhuatgR/VZDxRm2Ko+1sS3
Vx+H7ac2aUdGRHzN33NBPXK94jK8CYk+c+J5eHYRH7vLeqlhv9/y0tYJ7jQ6J/BNv3KSLBfJ5oAi
y8yYM7EEV9CO43ivj3J/uWfPqax+KGGJzWwQ8BzlRPWgd3oSYv0tfcwPaKP3r8fmAdZh93ZT/7aj
D9HHpY83UBAYmXTwAJBeiP4QAHmOVSI0yOuIWZPAxpyItlH08weDQxyBy/QFEGXU2re5MiC3AZ9e
QuUUzJVtYHYNUCCrn3Tt8b9mzwT4hCGBPv+fUC5z58oW8+pfwFxG4h8imRG33PH53xhxyswwOX4m
5yDiqU1ztIPOXNrjSs0KCfT3x999Dsan3NfIc5IYi9HNRFSNMoVtxPjEcbNcuuSjeph2B2TovK+h
Gn9ek13nmSaSjShQzlIC86KvmmPYTuwOSTJX8B83/GFW4P4RO7CF5XXNfa46yjJ1r8+Lmq0np7hS
X6LDGOgYzNFi7Mrg9WaYfIJydFQGtVSU3T64zETbdhP35QtkPLnQ1FR5jx9dWJGoA2VTgPyYQZnc
aHgkIykpNn4T/49wi3Ti4b+X6QP6JCRbuQO11Liq+gRGzkOg8liG7bY1pNiK0q8xrKLec6WrlemU
ow2Gw4BGq4/FTWLlbFBD45EeuyuzqPbopD3sPhUdxlzsmZSeT5I5h17CFdosZHtPmgdpNfwwhcTX
g+S4ZMWAAre+3wwOInI+Bc576AGeT9VL1QLXexy3Vm2hz4F8vQoEKuqSIku8qKuuN/mfIOmNuyt3
Mr0NkpoVudO3EeKH1xuAHht4k7aY25BQFMHV08IztpxUFaedAg8GYEmRPsiKhByKBXzCZgnYc7v9
PBhhDVkkXJ7zWRqYYHjjW8a4GyK++mAtG6wcDf+c3BNVLpk1sfYhHE2fucXAfyi1QBF9Hop6X2wH
9wr8t/J3mJphxXvvK6nLcw2BNDuzB8DiX7zmoyiqQTLqiFIoSimo3feSg86qxe4O/lc9u8HJqcP8
Y48ZWKyYgXW7Kjgh+ErP72GiFc5IsCpwc+6HTBqZTFSr/LfE8w6Hiz9clBK0uXk0ms9Yy9PUbi+P
HKDAcFsN1KbKR7AcnwjfLKqKrqsaXe2EbQichqX55kenZfVoOTP8r2XwayR76DhlCkDIw9XmdS4Z
Vnq97gtY5KBCxK8eiuC5O3tsNRYrcRqv8CmFUspbMI4l//7XQerDXooWnWCXdUGMPgv+q0pymYyz
lIB/iaAQDEa8aAU8FImyRge0shKPJbxHCP29L25lbqppADO8GH4BF0ius4AYKbAo/o/yZtbE9Wca
AysgNj/3uuIkbkMroP32S73AQz+zdVrCqJjbE9162dunTfL3NKlGDjmpbAfkURA/g9u06275nmnG
Zj+l4Xna6axkWlICD32obiANV9zF/3ZfepR1IlRuC95WgtQkUZDWzQz9BuhHE/+3ovDP7uRWBEi3
49zVZ82cf5zoTXKep/fBvu2QuhrJ2fq9XcvJTzOSZ3ixCGMs64Gz8JXKc7HDdK2bHqKjNj7MG4a6
FE3PwZkAB7iHPLJlVKeG9O2Kh5G1MAELaLiCv+dIT4E+NBmY8bRM/ry1R/CAljGacKtTG/i2obw4
p6Qof2l6ul80FC4bjNgZrYuOTmkjeysHZRR2rcrS4+9T9u8mYXzV9yLYlTYbm8pd+urhQ7nikwUx
aj01aOMgnT43XCLhFYcVEjBfKrk/40pV0izwmPxoCqagTWCojFcMNPnH7xT1347ghFi/M5pET2vQ
W4nAgl1MA3wGZy4LLgc9DjiSTygg5oMyQT8U6ivBmfYRvIKehYGJ/ZSsRStsF5etslzhMabmNtpv
xN05z+7C/btcBb+C5Lbr+zxDZbcDpCi78WOy82tp4XsEXjStdg6vf/PEqqDxjj1nUM5X9QidMnvg
U9sF3x8qqSMY4oKmU6EXZrl0r7RBsKPtbjbftTqk6OVQ4yKD+j40TqpingDxjobtSoxisNupVNKT
83NGMkX1RozXFziPP6O0s7jy6XqEczUPVYNlEQ8CtZAzaAMegaM9O1KV+TvNVeMaNs7khSvC2GaG
JIwW1stx8xT2t/w4+/T7hCeUIUP82belvPx0cDAv9pzUNxKyzjRzyvEfe5cBIZBr9I5G/PB6kAx5
MuomhfoPlaAeJ/c/Q+DAqkYfKCIpiQXsAs7XgT4/kTWU71k70mdN7rFyLRKGEPgGKNalBvCMmOtg
xyGToPZnTFzJ1w1R/YzdWNhP/o6euWgL9zk0pkruuB4zUoYVO+0foZo4KI94NDuF38Rysu55Ufk1
YmUP/rPqVdeWh3i/0YB2we40sp4kyCH1sXMguJKlwabdkwJgKHusTDw3bF5smq0di6NJqgZKbdWD
fduj7aDiqosr1T7tZ7JuTNLFNZD+hIHqNMo8Hh303Bbr1ytOKBVc6Sic6LLjnpe7r90VVE8nJkhb
z1+crSNBXPOpL2Fj6m4WKa1PzEsD749LIZDXYUFUu2ACgbZjypO9uiAYjWteudJC+SwX2DlJgDJJ
weiqGvx0OmYFX6YDQOTQnondJbjRVh/cFkMICQC2TWi+rwzCThNS/MzSwahXEVBeBQ/I0V7Dpcru
bv4iCh3HxzE+oLyja7Eo7BfU4WtdPgnrI2xHd1jSMSBm14MH5Ip7Myrp++HAScxQTDpNxGlIkqlF
gDufd7P39yOrWS6OaAQSMp60YH9GPZsj3odw8ZHfeojc6aCmGsQZpL6Wb0CopEy3UAuMQr2d570T
Ts3cTjYZWHJcHqP7SAraGQCJC5ZAyZsnLaBdTEt4Fa/SIjg3FFSTQChQc0aQ0MuOSv5xc6oNemoR
oA4tSMP5eTdsjAAzYNGHhvHfVuiV9CXMrtgkXsnRgzx4elHe4sSziX1h5YjixUXfaHzImC4Ec1ql
u4mKflhFDzwaH8iwQIb/1qLuvBEhzRFI5+tUBS7ZO45g7ySPMlqsVeLBU9Iz+B5NOsMVE7XSwhNX
K8c207g08i/KZB6ZJVzLPUvjYdebK2YL+7lL4yKvZxKSPaVbOtQ6A+ioAn/WgDGOohNDWv3n5mZj
t0yu7MivFTD2mHmKv+JgHl/guZRVF7sRUglv6jWZ/DVtmBNDwEf5GNekNHppwOoYIACI/VWO4YBa
0NZIKAVG9Llj68s4SJ/YEhStdBkczk+1H/AZ9Dw3/V/AAWMu7sk5lTKKknihcGxMBSPhP9akqFxI
h9ySPlrfHnKKOPsOSGxgMhNIT5GlANr4yTTerN8TYulUrbqCx/1ZSTu5VUfarjId9N31Fbn5MNWj
MAlu6wUyODRFQ/EMcAUbETXagcFsB5szmsTUOdIGipPA/PzXm9W5KjXqmKJMUJQa8zL3x5yPPfga
dGcQC8DZLW53D5mJ4E4queFnxG+ExsupleVG4FChn/uMm9nVOplIOAcM8fHlAhi0Rb6nBV6pJCwR
NgIeGnY59fGejFNHXTx6N4MjI3ukWw8dRO+1kbEmUPhVQDDRNY/zwFKOFwbjD4goCu/LHtfC8sR/
0NKfMyIq5TIcKo2t6/qLZO9b0UKapp7+4mahxVP1bdfdOILo5iCBuabs3hB2sFWwVfJ9X5ylnSaC
Frq+fKKObmcga82/Hs9yiDG/aZr9DG5tEcsaN2vP6+pQPUtvE7ME9AOxh3FSx3ErJ6BOXshdJHb3
rAm5jmVDhTtETErPZIUMnp1sfO8n6tYTlzh6st4WAyMuMQr0sZRTR8rMJyYiF/45CKaZ5BAG3naH
0/HG36qXYb42bPfLdDynEACw145OzhVjhhnL6Fhk8Z/m+KAm0PqCqy4nTtNMCmm13aV2MX2Yxxq/
5/t5GO0oWPRHl/3ttB3z230pGF77KrKzR/Ukhw9dnZDeCHVrqJSzvT0dbmUD2xtpsQZgLWhJKpC+
1bXRDggo5kaNO/AjsqaHG7/XMb83nZL52stqKsyoABVaZuJvMMCqSIBd958/jJumzUAKjDhi1LWe
LPC3r4x/GqN29M4FPDKa6f9oLFpM8lmESsHhuNKis/CpELxmV6LEDKopnp7quGUJRTb2Rt84bfpx
wTvxacy17TC37B0BDchtyEjlj7hvwaokyGFXa+Bwo8BMCUp8NNa4w563R0PkLx70+BZhWSM/Bw7j
6bH01sM6S9JCTy87ILHV+9rWtR7tmCljK35z/+htXXM2ZX9jjWUxJ5i8K50blmokRGd/jZu99dx/
Zz2z7hVF3+E1bRRSGhjuczIuriABkARvVif9ucQnQDizEEvJA9zpfd84XNkP5Rmr9Hk4fHBX0/0d
nERkO/aLXb0y9KTO1MANI3ibPpb94hGuFGpDtrGh+EEULrlF3STSwQfawYQHfos0eOhvPKQUPE3n
OEBuYAO+JIsPOA00y8bZZUzXN0vY+QUSO5x+V3DPSrINf38+71lntcGWuQvS/pvcedRDIM6xD/EI
xfmcmXb+u7YiZgIxZ6qTJ27C0X0woTncfC+Zt5FMj2WJI3WyN/uPEm9g8VapX2BSslYwIknZwd8M
smXXJyzqD9YyPkMDJdTxCkqSvbAZJuPaFfLQVxlUAvYfsEH9x/Kc0seVuht7OuHcH3SN6BjbGkC7
c5oKj/MZCo39jt1QJOdKvKCqWbJMpI+g8PpSJUSy8qS7aFeAO6FV0rGBiZVrgKRcha65FOlUQWpW
hqqAOMqYzeXvv8Px3lrbOm0LxxrtLspkzUQnS7PuQ+wzzMp/jJ0AgwX8KkfYjeIZkg+qN/Da/WH0
+oh4g3hhcu31sg0jcae11FmScnb9V6B1LFR7TzPF8p+LALUQ35W2Xk9sUiwOlohfHCcjED9LRTmn
tBuY/D2E8TmAzXBoZOkqup1+hmZf+FV0jxeKzXYjQAGHWB7NuRAEya2PZ7jS9Ci8PtNo6aCh8r+0
AgPdBDgEFgaaN6ovYDtibWP4vQjD1jW2NUrB67IcuVaEkF2z4+fbPU7TA2w2fiVImvG3+r+iRZkQ
wX7c9Stk1JlGI/UfvWo4/PcWbcE8RM5RDzSIzmBV6cMs2M09srrTTlj41qHWu0Xhj647ZbOFHJKn
t45ZDDMBulWuTr0PXAH2vuRWE2Y0BfCP870VbhN1bI5ARht0ppRApSk54+ngwsrAgTKTOrvbP6oI
tH+T7l1CefKLiDJiHCUol/Nv5qTVyDLNk0EpymFSiWmYO2Ic5miS1WsVc/vlKcf5Q/cLfA1jdvTH
Md8F8TZEUVBTDVTTXt/Te3Zig2GQyOVzA77K6zM5wylSXaNqUXFgYgh19duQEP4idevHSCN7Nhrm
yV/SRT2ngwqhGE4AQUz0H0++rZfTcQ1CIZW6jtlOvdlYGqaiajyH3x9hZ95EET9JiILgRcJfrSMb
hH410tGojVNkG+D4QdnSxZT6nwSnHFFpiV6ThRGrlBD4T1+iLYCrOsMgsYCFL00+8+Yjfo0i+wTs
QPik2wGOXfQGPhnY7Ue/Qs4GSies7JIyloXc0gWj+NEGpYcQRCmwabpW5//fTgah6GVq3lXs5a2V
OXMBAmcaEfovfjX4KBVPqNFAAm1StN12RM3aa+Sf38neBJ62+7ry2ziiXjCfd8mgsSFqmicH6nIo
A423tuUbWaJvKP5v8rMREQJDLSqByO4dcq9n3msxIkzp2aL4kugRDsN0tHZHQaYQtgprVVLdze0k
QGdgb9vxxhG4aggN091/wf49mnAsNt5EUACMLnNXxxzJSBnXIJXCCT8lr05bBhPKdEHvryahfPI0
x2lJRvVZfjm8LviUkivvZXHPjrsuM6FK3aISZNXkqi6LuTmPvk/u4NQtxK4UWb0VsY8vZBkBMvxs
RtiBOfo5CbJeqFbDCqxk5tB6PKOOEbh6Kh1YsNzQKlaOrnR85F7VqOEA5dG5l8P2xaqlmaZwOFUM
DIZqzrnXuoWDA6Z6lvqRpR6oKdrSNy+o+4RnjQUwmFJT1SrxjKnVFrwv93FCaFcSWPBsVBmq1eIL
Li7gVh4lZ/GTbJ5V7tOG9lzpLjxP2Umowdm/gAXHzwlq38ikY6TqOh5+5P41AX6tWBnPKYuV363Q
L9zX/ZhHn4DH19bPdloTKFQA2GkZSQ1nTptyfgNQTSTx9M7n+QPDFzL3mdWHqs/ikKfOHYalCWSV
2AHd6abDEv9bAmM/dLxqmSzAAbtlJqXKyXn2GEbc+Pub4RbhxsAfflcm1QBOJJnPMbczqv0FmHol
hnujPDtxmgFxM37PAw44m95MAGziqmpbfYAhuB2Jn3P0VobO9iy+8i3clGWdwxvDO8w+grcvca5A
PGuQ7SHMSaYbM0Uf8tlfEvB4U/ZreJlUtLKQCpw2s/R9f1oWO5kuRQDwtRyjR0gY04cRUozcIV/i
qGGg8BIW1jOIupVhbjinACMMG0vtc01/Ni28cKrygL4/loIgNUkJej2LOZ5aeeeT3LtkIyJ98QKB
D0XeqKNH4HF5YFgBsmTts3pAq0AzxaJPDTXlCR4fz3pOiLNy8ccdsIWQwn/b4RXVQ3gi+L3+ocAH
DlHlPRggKAKWwkPppiIgM6Jgf2bWd/jv/VM6gDGAQEsPIbWgjXSbh3af6qJFuBrE6TUHtAZpSvL2
JMCFNavfLro8JKzQgUJ0IVRZEFFb5gvqDxmfHYSNUUySp1VjPgrk8n3v9nAp9f/95CQ6kC0Sv1F5
Wgw0HsK2y8obi1lhsNRO4AZmEN0fiPzUL+3ZVZCE0HrP4iNbthcjJGDQA0eI9Mty3HVcHJQB1bro
SNlzWL8bqs34sEgj1e1cHyyjsCCDMDcLiByii2i6Ly5JUGJ7+GIMaMOIAYAZ90tjjqbwgqQYxAiA
UzO4VxJKEeBzYmCdkHoOmR6zsmlb4d7QuV39kMgNxNOXCjUubfP9RpXZ/bupHSoy0IaPCQTzJbbb
YBBnh/AaCCDkWC2Gamu3fZj+/gwgPeRGVd1IBXEhhnm7/9P9MViLp/az5DAVt15efeDmF3//6DIu
T02tBBndYJaVk1wJWJBXmbl04quhmuM0vZujc31gpmBSm286XaDX0PiZedoovr67DhoihF4oiFK6
XlObNuWfTOcFrk+afIrduG1fMcrofKddNBD2wxtCxDTNcXFbhRqPcDMqQsFwBXejPe74xTD2m19o
9FA7gCy1k1/+L82GuGyeMjEQInhSlcCwoaVO0xyT6Id1XiEU8kLNnoBQEGDt3tNrKmOYO/UktiSP
zeyukNZc4jVGz+i34UtvnsAC3eotKw+In/FjS+sgZnJvrpwmZwufBYZzAxNpAI67F3UVPpboIPmz
dggfw2zPiJVBm8gNqXRj/vEwFaXt1ngWJuEkL9KqM8rxfdhpg4q0ufAY/5/L7WfhWM8IBd3P4dYX
62Dqc+0P4T4mps6Q5Sty8SSHWCVqyZtJGFUD6ya3xIZas0L8Fmd22XSfsax5iAliBPN0Iu/uSfOe
MGgAr6jTrNwuxtQBB/FsJiWEn+QmVpri1ZHM0xt/hbLkxtwp84qAlsghRmJHBESK9pPHETKdcJ90
OyTvWqvBhRv8XaMQN5yRzaNZyWhwWbb3NING7SwjPFAi3EbUNKrN8SgGbyMJu7vzk+AI8+SDBiFr
Oqn2+DdEMdItsJ7qboNm7dNh/q5rrthltcPHGdCO8E5PcueiS6H/wLNSC6Zh5NaWYvxIhrpeDCid
+XQkuOt895zrbVBZUOlY6utT3WtW0ZklRhaF6yPSo+CxJiGz6AeJRHOp/vYDeuQXfiAjlBCo3sbK
bthhlZv/iN4EDhDmn4o+Uhys2Q/uiKv59A6lURvxLU8/4WZXED/Obr+f2KMB0eXBfzAeZjXXqfpA
OYxSwmtY1XN6ZR5HfjjdX7KoETmGPktrYGmIVNhvc5yWqftyjGzgvIt+hSax4mwAwGT8Bw2p4LMy
zMUI3Hk5Mk9+HKJJbsG+Ajl4E9Bs7ZF8cUSBl28g9EEIlzSeYfIwW1okXR+3syXIBS4hJNZYJDgW
ehXaZmI0c6Aq2vbqUh4adRMAux41d9bMhu/+o+5qvRlg7agK3Q/JO1F+WCqMSYiyb1bcUosPJ0Sn
W8cawxywASW5Fgz8G/Cd1Ee7J6yVjaO9KAJX4AhUkzxWuZ1XxGo7dKSn/2FZ0JYAUWDyuUvSDmo4
bGqSvsMSQboOgk+bQUIw9Xc7gAkPs8/lcyFz+G6DJyuZiAhGThg3lN1g+gL1uEekaoiYtggvItFH
PRBRxpQs0rFu2AZBCuc6I8AloEs1vnCu/exse/iSpdETvVWrO1rCSrd/LPhtttWxQv/PgfOXcQF4
8/qNsYV3YkdJkXp2v3HCS+mI6UyBWASSGZQ+J2wVdLhkP7PUKqIHczbc/AX0MUg7XqVTSdBvlg5m
d6rZ6Nz85/vIMRCAJVwxHhvS+0PkYEvcOB6QzmjLVMahfvgia2LYMzNPbyyAhr/Uh7Ppsyb1D4WM
ur3QFZV8YHDbcgOzkgGlnKP8Yp9klGO8gqQilb8ugbF1cf+z3yGFnbMg+VdPdx5kCOICiNAuY9Hq
Nx43IE1KrSsNI38QLneeFd82Eye+kqIY36Ep55NVlWuhfflEHC4/0YdJgP5gOpWjxvF3KJIlVrPi
o2RBjgXJp19vvCa7DeZw+cLp9h1DiaOrk7n5dQEOlEY7VQWc0xd+XQjBJt3sq9rYwIiyvtdF5xMb
iPbaL69ea7YsUm6y6C83JCjcWiEbHp/hSBFo2E42VmSAPgZX5hHCUJE2czhEG9AqRsVEUNyy6z5G
ywp0At1jRHiz87dUSoRIrliZGnSPoecFHFKi2L5Pw6uDMp7tHYLYvx7paRUIL9XYYzapJf5YKSE+
R4R0LIKFyRjI7V4hP3KoJntGIvYVSjsUz7fE+YFb4tjroZq/BYs1eSHedCQ7BWrluP0KmyMID4zp
PREiuvh9EW2380BIw3L9xJ0wLVzVqySTGBKTmhfdVXaEmOkFyge6AXZSm7LrI4qOBgTY+AyBvrUN
Ffri8PIGlcwH3USHafhpqnZG8HRjPR0xXySscs1WQUZSmWAAcmUmqyn2zbXBgQ9YwOr8m+7O4849
r8iKX8E+wAsibRjDMBTEmiRQ7wCMK+swLrhJwn2wxS+9RWddY7/nyxW2uiqSz1TSlzFyZ5/hilTV
+5XZzJH25NsbPk7MpaXW+pNZWM+Yjj8pf+XNayCYQYwPpU/3JTKahN1IwaSNpV7sRwvVSZWmP1zh
kcboaGfypy4ZLNgaadx7s+HXw5aGjCHyRqsVF6BeN1JLz4VOzhQOQGVI3+buAEmV/aEZBewzYfC0
wWY18QOdJrFcC2ulRdNbUbX4tIic/95DQHObW4N1Ga8+S8bWgOJDWT7vc7I+lvPwmX71m2GE3hMX
JlUCBe/E48psFZc1IgZ3wgjEg6uw+gDRXuw0k4pJQSAj8+tw5p9fWQQ4oLgK2MekNu3fGUEDSsb3
PnM3i6iVYF9qsQZKKffSUrogmBoST0Gl0pLmXL4SudCpzo6tipFb52pl/RUICwd0MZasBU7fiX9F
nz8p42KfTfzklOZolopW9eelBFOO4rtwsXvrMEGboAhJjrL3FgbbTLhoIYSPdSeavU+ii4p0qEmF
TuFJc4+Z3p4Fp2CG7ooxzm3w3cYiVSQK0iy+MzA27kYbSAGcS6/HWPgC40A5t0HPWle3tB9MT/Oi
UCug1HxSbWxO/v28b5sWsSgXFlyOdrNvvSAFYlPiOjVsOd7sxCb5hQ7S637Tte4DoINO7H8g3pxe
jda5a+P9oM3wt17F9ffLkzBPh6ePj9B9SZJE2qj6RpOga/3uSufuk4rIW6yMpAwsMcoDWfqbrcwx
hVFU6aTJAj/lPq3Gh7azI7WgvcQUVAYe9SZKuR02jH6x5bPLw6aHSPCx2zxc6nRMY8EVFOfQhRla
e2WEBuxjmvFtjuA3KI+e56THPn6KWZDIXhl9JS/l0bQEA/JVAPVB73sJvhGOMjsS4lD1dfjEwfY5
jI04TjAChwIb7h7NguGPBGjNy8ZdUWk17YqQRZUrdFHOlmda8s8/NOqy5ZEEMQ2gHsMy5MC9IZ10
kOZvuUZZewB0Mqf5NcDpl/N3sT6bnmBymPQhXM6YwYdUJICjwtdIZw3iWkiMW7Lu9iEStlXUOwOJ
BIUGYAhhGbave4D3FOA+qRDPnJKU/azgAIEQkPHQNMUjdo13lLqzdPQuU6of7qUZoAYxXUI9nnfn
jKvZdBWiXU4OMgjpX8xNFVk8EqvEwtmiW5vuuDCXyTmlGewZNj+OmOinhDTSjSKzM6h9QLVJclBK
i9hZJwIqdQyhDmieY3abn3gupceAX+Jcu1KJ9htTR5aRFZsVydAHjjCfamAbvMS4A7I8EUc921hL
KxsjoclNIvxQXZ1WF1OnWCdWS/pZr7snyI3ZX1wn496xniHnKR09ZH8BjC7TKhAaC2tAbL45Hzuk
u05aZQmLXjbyZPPn4x1tvoEnuBUVvyjxqnUIEWBcitku97yL1O6s3xIV0uBFRxDZp3x3WQbDq5ca
G3hCxKbckTOPBnULBX5NRUy+SiWKA7PRqJ8548uFQlPA2CUMs7mqQOPp/oWprdmreEsky8s7z3UG
FsuLyH9li4uPBg74IxV7tHw3KiKe1K/uTLarK4vzgOy16sKXK6D9+kTMxFi7qnJCdEEOPrhAZMzR
diY0BXNKHMcBLYqq4F5TkuGsP+1cq3T8TlbXFoJbinpeu/JUlTR/HlqvPGSqcc+INbJPb1A7enzU
yYAMObVJS+NkWph1xLU9GvFeY+1yVKMQYQtdqlUo/GHeeMLDOfhHGr5eb7qHRB3T7pSAw7Dqhnrc
YW9TpqHBrcPf3aKnHOhzq1nEX17xZZCqknx3L+6yNiekEbWowukof/2NFA6kCmJ3hibo4GdLRq+D
AlzUEcB3mGFSIMTvk/tvdpOs5VVkQ/r89uaLifrP59yKJTC7CcNTY7y9g3z0mL4jJWDSca7RVCaj
B4bmcOO7GbXNnu9DpHiVUaOce24aNH6nESYsiXraTUL16QNwehQjoKYbuUdYlWGGy+B9qt4JXtgj
8hxGbT7gsGtDP4SI/H5Lbk+EVdHZeOqSUL4F4S+dj1xGOs1sIFW4mZfu6gzMzBeS0xWKAScUqwfX
pGrwo1GVvkXtogWKVCazWgDJrVqUvySQUQ4X1D90NTzdV67GFJgKH7cmREXNL1BJl5D0FxO44+mx
jfOhJb8MZAyO/wEcK6TMKDcMvCFTuK0iAYyfSdqh2q5yHHWBgEU1K7aqCbOeCOnmM48i0MC4CiJk
39TvdTszc0Xw3IK4wjBzEqEcphG6ZHUP2B9Lq1JEoF7F3RdvsREyr0G7sVi+hVE6ycctLuoLJFjj
wvNfX0S4X1/udZStbAEhM0Qm1ev+ZZivpCWNSPFKaqZwoiHaUKqdSACFU+lb5+iHUopoDuplnNPj
nL++2FokdeF3/HwiwwWQnSklI8EDVeEKcf8fOhYAVafGoetFEmy2elGD/72wo/U+HklFeN6+Sffa
VeGSKsHhXT7Nic8xGQdgwdN2UG496cGR3u1gY6lyOJDCK0LJHtdp0raCBobTqqNj/Y2a2BFRXZ7N
kOTfZsxYCqgfFHkjgs8ykzeZbYjp8OqGkLF+hMC6nZ81HSKNDT7V8tr34Gfr5jYPC6lSoR/YpIJK
CY+uzvnvuKna64EcfAYEKLAt7ioHzyBZFG/raNh8Id6ON2EGsSZ0zxFt0UEW9JyrblXNg5IqaYJ/
XTGizAVy1RnK5cM5Z8TZWJU1bwKybfN9m79xVAJWnYGdI7V85CZr+hvLG7X/4DzvY2FNZd00wiP1
bWQfHtp5qo6BhdH2KnyRc68sATbIs/cRKeEop18J5oUmCXUAyFgwrH6mEJvM4o5PnVYSgtvMJZH3
fu1lVh2g7FfhTSpeVkbKcPSuKTCsIZWAEMMMktCpgklDVeU9zq4r/MkH7QppU6HRqtRfEhBLHr83
tuveSON+8YhJ5UOmx9Lwtns3ICVunhIbsxSmRoLbjOTWKe++Fm9yNyuGGPZzcb6a1PDT8Q59XS96
U1e4MWlSjV43dyBHDa7JIzV5LEFSo+UyBETQS8uJV8+7yGTPJCGBegiPR+eQAy64pv5zCLbSp755
QDjdpI16S1kuIIryApXnGgjOhza9cewiwU46sBswK6WCcshoOl00u77944e+DAO59ER3omk+ltXk
YjzmOOOjbXGtQObYbGXmfyLgrd5OF3WWT7U2lmr47npnUN0en8wWcveiMGl4350+gJOK6ooypaPv
ZdlKBDaqYyxL5QdJR7oEellPsC0Fq3OiFbg7KJeIEeBOlpdu1+cfraOH/0mbElqFuOkO+uIIlngc
GjNV1+X1npy97rcSpWO0EUTIR7SZdg0iAQCrcSODS+p8EDjRA1Sf9Xk1j/FGweb+1GDUd8gawaGS
53qMILi96iekdZ9ANxgRlgEoCwKTS2pL9ZEvBr9YejRtyl0HN2ahiJSySh4ngmEYraNQsHhkOc+O
YEN67FyTjNaRk6EtdG1AdIHL0icU0MjCWaD3mFSDwjE51RQlGALFmouf6xDwKH+1ZizUy5TytYpX
J7d0zJV9XHTSAPLu2+8fnqz1wDr6wNIdRUWzoBM72GNlIkoDBNuYdOR03iXqBInxkn+JHYVvrhhD
Fh1+fJnirc7jJE6XZYbj9to8XYktZAL7i779wCDtL71xZsLEvMuO/MU5Zk4syT6FZnezVFKC1Sum
IsvPxDiOEd8ZJPTCTDtNrbF3/IBfYmw5MBp3Clfmk86rI3pVW6JxUucvcWbzOpwY8X5/PWwfxzjz
qo1st+dZT2zSPM0vq1ATajVfNydXd9/6Ewp4K5Z8ut7FFozlXFTptMHVISyiXP5CM6KWvqkCtvSj
pTxXsOseVz1xrifoHFU7qa8ezY5fLo1WBmiHhJmMGDec/A+cBzjFZZ6zXy9A12Jxd1Sk2sGa7SUB
wGxc0CRxaClBPzgiFyf9ZKBj4+L9ZCcmXk680y9yoqY5hBIxI+a38nhPgfuxCcQKwxuuOdHa+y9m
u9m+PHoPOtw28v8Ll4ZRrNTBT7/o3nqxvByjj/FyK9wG0Xfq3MHs7vKuy92/owjnl664GRG8S0xj
Yu80GJzZRM7V2Dgq1FEqNOJrkVGCAxlq6dDx+54vpPnfvFcFrhfCha5B3dO6Rh4hJLU4B3YpwDvA
E39NMXHRpa+qqmBy+n6wJXSGzymL7QPbFNe5Pz64FNpLdmpbq71XSVcEFzEIB+mBZ1wkKSVG8/X4
If7bEy/QoRBFLYPARj9juMOdy+ALig/hrfiz0DcbaGZ7r4qCxfksRkeAL7I8RsjIvEaztJAyXhoe
3M+hXURO7iq4X9WUzZ9/lnOyGiABUeNLGuqQnIQbrPR970YS4P6zjLnz1Ze2CTvc9Gr/1BWFvzcI
AUmIi6kseyghfOOerfo7Pjs7UK8FkSCvwSE9MOPS1wtSJqX85VWFWgWDA3VMKobVS/WK982YmufK
ifb2OVFEfATMThIRqiBTATvyEPnDRIpEfgZw2slAS2rIYyTwB6Q3wBpNSvWW12VndZrBKWDRukfK
UnZhbduB/Bz+v9Dh8aPr75Y9AxpPe3CzmGLM6iLUHZ26iiSoCfoBdVRCtMvzRFN33FXBhQH3lqs5
Xb8s49zHF8mzbmjOpGSN3usuonuK7rJd+6nuPLTZmeCC4ARk+8BjjGSO1vLeVS1tI2is9CYZTLe1
pEohhtEfy982QZkftwXQFmtlMSiYrhM8r5UkC/Jsv9wlWtkohHcE7hBNL24ZhZ1M7S0cHY7QTv1i
/jxQq/mEQR9Cooszst/g3IgG0hmTddhGIDhnNSvsrI6DtTx792qS6z034S1m3nhy0qXNu2jVvXnt
zfz3KrscB3ndFQCWdIWksZ97h4GNdEOtbgMgKBd/0YLlmUgz0TBQ9Y7G73F1UVy8n/JIpwTrksK8
AXrHzXio5zxAA0OsyX39G++xd53kx1Ly/2FjHpWqMk9qHShDei/RU5b7h0pV6rh7zFdJV5ejmemR
6Zg42JQp7OD6DbB/+O32gcN7IV1JbT+4oCwPbN3jg4zrgmJCDSEI82EPBoCheADZNyREpUvS25V7
nnwIShx3BYXBr+FV8FZZQJMwdZfLp4qajhGaoUfuO1DZpgxeq+k4R5FTGPtDnZOuN62ri4PwDSSp
lkCPwDXoNdsYZGp4HR+2JdP3juk2pdo2Z1ciiLNHugbAtITG36rsZt+Ck2CyF73RGmR+LJ+Fcckl
YeT+kPEzme98euB/9IR/3xzyLM4MvSHu6kR3Scs806Zs+jkhHh/pMfuX49OljX4m4YDCbHftC8L0
7D0oGF6GwKyLW6c1iZeC1JqF6WR80Sk8wZ2ybqJNVfjTVWxcgI2Z1O+riVgzTV4oOqPH7rZdSktO
ukIPUqW2CiD/+73jfZaKHDihYtzA0jrRpLJO8F+5lLXgIZ9qcasjeTiToSTUdvcQWSf8JuqJxonD
grDZo95ueWbyXnbl3SimNDw+3vIS7tYPTA5WJGyQZLsB021+1Rg1SUN1daX/JX4KuGxCrq9APsxq
8lJ6cYeL62RornMxsnyixbFXHrA+BahiLskwJrBhNTiODJ6VjWrz+WDBwzHo65yV12Ams4YJ9guO
7+WWqM4oEKp0R3LxWvUxTKkoRw6r5U9UF2qn3/oyz7QoLJYB2qGsDEcG2IBkbozO3zD09w2TvBO/
JpDNvYhazOOlxB/W5uzSpOLW7U10tvnMbZTDZWp9HR++9DmheuRLUFs5HPvIRYQTswe6iRxDyFtA
fYl+ydOFXUo/7/ZTC5uI9YqPszulgzzz9wJO6TqYQLPJ/T/ng4iaPD0Vp0JeCwvyblMuEgdisJ0o
AwRMOeKqyQKzYiVE074O94/Tv+by1Ne2IpiDQjM33j1ImI0fq35wx2hYXCqgeWcBFWH61aMxNlaM
cAfWpGGr6cdRMNDyPGWA7R2T4v2uBAkw5kWOFLQ3zhM4nLjJlN4WWAL54U2OfLxZ7wxFN8qtk1CI
4O38cfQ1y+TyH+zaCXeTLckrDDGJUnNtDY0xAuGZGi2SALk+pJfJhTa4dnfmlkKwS5SrLOhlBzdP
6KdSau9Ikz2xcHlVsgMiJdnFcZYhUXJSaglv0OoCs3FLbyaj/HWC7hVawZpUkZGSyrXkFy3CBgdX
+DobQFHev7WCqqX2IUTIKz/CFgu3OsfGrTfRI3ONmDkWKavSU0xX1FfVThwzTYu5FUi2vbLFZrZY
7cEEeF6hEmGGSsZ2ssaJpqipPJbDAbB2Hhf+16v80gEgYC0JrNvKwk4bhxXRIp7QVBL6pYykxALy
hTYnAVqkbMq5j31Xgxp4wv54Sxmsv9gGW0P30tmq6FAHmhTyjnDUc7mdw3ItgR2DENEwC/vFJtDs
zUZ1TVx/bekcG53eIYNCpwRVavwRsiBamhFsMDdYlfEp618V8ODKiVaCwN0PUzz/thpO7hm9s2TV
I3i4NZF4wFJ9zb2Vaa3Ur4U/RVJi9BWrMANqPxAor1FiqtnK53yAbsGUrzCGkmSPbMggBA2SwYZL
7BFQjtimZJi4BwKAikeITVA729e1GSmi1XQbxjkwgYnApiyUYFuWb7NAabRmk7KunxGBGtmtCokz
KZvxlOx4GI1oXY/uJ1bzqA/ih5QPdKlauAfrwhAzJLXHPvGO5v5hpKm9cWhUwe1r1xmn3OTadGt+
F6irav2C80mcxfPlVFZUOA0VJ/JklCbYE2DCIlT1dlL2/NQEfT5f2ly4YswtbhZDupqc3XrDH7pu
6AmMwqb1iJdMsF58VyHBucjyMeqPyOc063N3ZsYSoRKS/rE3iyafAws6Ksw3wHZ7E47ikNZl/ASy
AO61dQeFCz+u/SKkrvt4TmDySQMYyTuJGvW04jGurb1bKaXGy1hpDVBSruhV/Wja0I5wEKw4Ar6G
2o7wU2xBcBC8Bp4xZsR4S3SVqcu8ck939QBvvrl5O78NJYzZdNRXqEGSWqf5eUPBTJTnUPNdV2Lo
0PlRj6zTubhUjl3JgQ8h+khX9RCyAkHYP5KcTRUfD74VYYa2CmxXLOgmgIGCVWtHKqMQJojfdaF6
echSNaYxPUcp6qrdWt1ISbcWssgzGewRMbweHLuP1HZeTJv7uCq4viol9x1PlTzsUNkAPCUx9nbT
KC9X4jLOu3+NLzd1UDlAB9A/cq/2mINE/+L6bcFvqB+WJd6/MI0I/BrplrZObrM7NScV26hg6i71
pXUHiCWHeQGCcy2t1UZTqMu7bv7NJZZHHFdowLrRBoRwU+ILOxwF05yNPTm4/E0u8qfHXWKt9Yyk
GwbOO2AZlawWwO8ufPDFDdDowaiJ9MWg8aU9aR4Ub08gROpnQdhX3854kqz385RDFwP6AbnRPN01
S2xmNywBoi8bfy9AkphHNyq5kFlfI8UeuXfjxjQfh+jEI0WR937gxmihHf0r0KpFuQ4KRCin0ojA
5D1P86b70vKSGOMKocBymgMtQeabq65eycLlZnZ7Z1csTWoVEzF6rtZ4oXqJh5ew+QsBH+Y1deM2
7OV9/p3m8ZoxeTBpEAqOlKU8HbnpU5stqPs09/6OZMPN8gieq8I8rloIzKaGBvCppRVTTqld/5TS
OFA8HlBlVzg2EOwpjiNXnmr+MloLnIWb5CZIfu+zdzzT3IX1dtvAJSYk16KpnynBZe440IFPrWFk
PjtOYW7kVtqPQbrDdt6Ud2zB3jJlWC0yAArXWphimeo73P5VVjcC1iQxb6LbB2cuGM+uFL6nsxv3
y1/O7/RCsNJMmM0PFGGXF62j0Tl0BC95UA4HGenH8hPEzl+nK8lgZ8dSqDogXY6CWWLjK4KXsRfJ
V+9QWS8blKlZKFgeLDHg7MRHapec2ntnc723GgmY7AAAK4UgeQO+phhB5cyX04eXPPGYJ9kCyFiO
skBgKh43qwYKPhrlpfwkpB8IAupHlBPTm72x75Oi5FVepM7hvHGXCG8+97ltjXM8xnDDzYKfysTw
tez8aJ+ulvdD79/ts4gxI0WgycTXt3VWQs6jlVOpKLrnC1+L1/2yLnqupkJNvpY/r2CGeKPpyV5x
bNi3Xo4kvp8HPBwa5gfXRpA63yd/XxXcM9u1YH3GkzYU9pBMrec43M6kWm0BgHfHmEftuGYQ5JgG
5djaOAellWNYGd65dI4eIBbxa5QgcZnuqevuRwgb94El4Kcb4zqjwTvjwTSWF+vqEo1QFRPqZSrg
W8eRUw7vzgMgMgHzq+GGvpPcaRa8r0zBcOATmhn175nB4BqScjj3Ug73+x44IssY47b3Yr2Ey6Ea
ZYlmoU3z/x4Rsp7OE7H9CKyCPXgMzsm+tRLDxLSocxwChAm4Bisy4vs03Oe0iBbfUn0tTTgsZOth
HiOFc4wfBb4mn57rMbsuujKKihDps2S6M1j8Akl43TMWxzIbU1M8Cire3kmggV4C2phy4Pwx1HXs
rsQz8mQCH3g1cKPbg6ePV4mb3lxR+lzmRdZs44DTbUeqCutmG2JS236CGXL0LYXHlnRa6Wk3GmjP
TsOVrZvu+fvL7iQyYJVPQiyBJMMTm9cnRR0omdsFRixnohp2AXvv90uNt3bu9ehH4BiS8+gV2Z3e
r1zxtn0hIUvmS9hUv0nJsWBtWwf5hUWho84OVqfUtIHfDeqb47pkRg9sB3ou5Rt9eA5XB2f1EzqS
sE8Z3gWKjBfaXIjFjYXQJFQBU76KcEgIibR/gAKrtmtEJA/kISE991BqHQClNGumTA4nfHLMq/DK
moo/YG6DTNGt5K2aelFOOLnusIzOroQwDnUakaFJbecw7L37bb9O46zKVqe9a3nT+un4VbXd7lSw
PmKqDNfxmvSy/yvHG+j5ZWm/3GtZCBcylNkIrhHUbYUX3bTYpob3MUxp80j0yb+pYSDPxDjHn8/E
lwUTa70Uk1/k2W/uYzF0eqq6wgKE4RZ2KZxfUg4XmEpNS7AYVl0at/cnW+R0c0sr17WG4vyQwesX
MPzgQNtuU3gT9HtfmhNOS/Cg81ipF1f46y8NVSm7zfZs0rBTeMYaDra/c8R/LV4K0TsswFNRtpZm
HWzAbmXSupJGLsHw5si6h4VTZn9XTyPkFQh9JzXals5b+NukcyjYl3EsVeT3MN6bxAOxhlXfB3dc
fjc7hSnLzGc8He8LnP5nOUl0VtY0nmpUQh9ZTRhl3PDbnfXAY6WSw47Af7mIzRDkt+N+rYWGW5BU
X/VjmSPr0HKRl9pl0GEAO6NGshTnSr2sM6fbJPi68au8mVmbcRlp+tSHsIXudhzLCXlEUKPXvZ8H
HAH069hfeenxL6HoK5Vr38IsaS+lJVhj3A9wVu9fD2JzSyZ9OsGAhutj8XCO/cp04Ki4+Ba00h0o
X5jW9K9/fIwf6kg7aeM2wZVzQ6nVQY5Co9BDiEUwSM5lBNXSde8YrGLMnj4SM3QNrTZRaKs5DMmp
dwfil80fP0J+b0h9J/slkwq5CFs6aWydqUEs1AdVUdxw5LoxG0CkTU9lvfB+yQ1RTyaeq5Bg8bli
sK+b9nngSKXGj9uUghT41AIrCbUKWiVm7W4RH/zudc1DNWbqPtQs2g6F6fOQ7MQD9fV2xXW2NHgd
QVGN6ZliX5fACmWhgbQxM02qOlksJrY/vTWAI2rG7os3+TmtJCJfLgPPkzpy4r04jOnkO0OUdbe2
3v93k+L5P9kclZqHBnaXkkqTmDwQpbPCYb4+ah4bRWo7nzLK0B0Yai1yehBZCzRvlvP9vsLOkzB1
QIgJ65jwzERDxSPKwjnomyqs9VmpOe3hUDILXN0CQV8YXDPMbv3WvDXTFwGLaBlxmrhnv9C15N1c
hawg+Kr9Vu8u3Gjly44chF81zY8k5u3mynMYFqVq2KmTphY2JCwGuF8bqQTfDh6vDZ6VgiWwOm9v
gfVgt5m4B8dEcvA9alYutB7OvTLRGwMEaCvytSex9uzsvQaH5lwDBQTyrq6PaX8uR/1QOZtkEd+g
VFOcAOjfoRuLCBPX2v+YFCCaU0AJOLLH+sdCZJWv8fn3RfHzBXzd76Ed9/lLHYOcIpiHoEzVdAGy
yFjDhTG7KsPOcYhS6UkB7r53f8nfBaF6KhfOLR6K+m2e50iof+6t1skYdTtQXLh2dTkqrqqD2oIM
zcO9D0dBouashKvtRp0q+32oMlqZHt1x7DGrwBECHGJ6mYec8lloX0mfduhFyDiwctotqYaWuvQd
mTtPjPuzPbS+0sHl7Ojr+TNwhvd3f3EZZIEbHBRfSPFaw7814dxCofgkH5V5Je8YiyLDKpy4j4GN
ruPKjcWTKo7X3bHfJ+FW9N59YDmBZqjNGrNJ36DS+uc/k12vy6sNEdZO7gVV2NMyKl9XkMZeJfvz
eZv4PjVpq/s8l1erytITo00FkVur77tDf5qkwawSFuEHg6LKSexbsQz7KYsfDcJJzPGr1r9R/ZjA
zSHZD297Lx+qH4172Trz2mxqOnyUi7FOxMqloCELOQOh/zPcJjB+Xr2FgjAuNVQ6ruE/n5YjxYeL
vw+L2bqIC8uYnJpC3kqVNUxiWqUTINorCi2AQiNEjzM/cQt7wdYS+BFrJ69rL4lFpdr5fjfEtjZc
mlUA9HfplCa6UWuPy8hNBIvXFPhzyDgL6HfWcV8WelfX+n6oOtAjW840T7zwkVpQU53ajWKTw7oF
mS9kmqZS3zdA+idzvaMS88L5PDxUlbJcQpN0RKNRuDhcouH+DhMiE+eXCzvOKh53bDr4iEgoEALs
kbqpzt84vY4r27jVbDfe4LFlLIggX2LS/LrGhMA/r4DMKkAxKnVOHTLsYvNnwxWa9f4cZlDHAu48
KcPBJL3orWIO+XY4bAfFs2eiNtgVOPgSQmSogTW4EPVnzEpmIX4dv5BkSGcmBL6HYC6GVZk5FZ6N
g8Vsia2Vae5HrJel+TsoZ/+qKwTeTtlu7UBJ1CBOORfio3hn1MSEFmv88wBIT0bp8yBl5WvdLdYI
7pXitM5ZluKSirWpbEHBIpok0yut7xM/FMO7Zi8i4xkTluTA+QaPBL6wl9wWMnQFuw4V07WfjjVI
n39trG+a9q+E0NW+fiofLVM9pFLdL1v4dVIeORtBQYwzIdBtHixnqo7hR7eEcbFIwdw3d8vKXHe+
b7siTL6fgvKUr8A3bFVWusC+drY4Qys/2QJDPYJZDlsRfeP/3K8pa7PPTHEpgfxU9h/DMNdiX3Vb
TmbqII3hqbD+fapHPAVnX8lrauvZzJyM2lhQ/gbvsOp44Ng8IbLCLk6RLoV0dzbbr20T/VZQZubW
rKXlIocYTQSlXhsRJdhvAsYNBqx6zKjlfg5M5PHvr5SOMv3iscSBd26naCmio/FuLoHbZwNyupzu
ixBJaxCcZXaOuKcDz/Sxu0wzax1jaUhjWoqcqcy/jc3jJv0BievaLFbq+lOuY/bn7LVP15ltnDlN
rSlcfQ2npJsPcMyK6QRBHdnAQjJxVJFvdFTNih0KMen5STTHnyDSfyzi6eBTROlbpLEyzWKFRfZd
v+0ivMXLWjP5oWCVkYwJgr7ARdlkTpYqdWl6sIjy1lY/azJItd9DtN1fdRRJ/WrIS2t0N8DfR/9e
V7x+JKPTnFf5pr6tGTG4I7XACGrXRJMKDU0omF3GwDJOdMCI+988YW+TSULbJMXHZ3mLIq4AUZLZ
9vW1Z4rLayqH/TFMzlqEQAbU1wxFncj99yPYk4fiyTbnRX3zVL0ZcFweLciyBOv9ZTBCjV5o+Ww0
NyyZ29EfUvb9KvXYnS3ddzMjJWGKFcWz0G+M3JPSaPlMecNa9IRkSTqdC4V2uVdqpEJ6iMA8eeUt
HPqJu7DyHI9xF3gMCgYXBknjSnbpS205UDzUgPxpqePe7INNKz7bXns0aMSSqNdvdWTCQt+ZLPIl
rGgToJ4n3Z4OG3ZOC8O1/VsjTqBCHFnASMf9D5G1vi8c2SWA28/gVhiZ/l4LDbVNlZ83ywiTg2iA
004kmObixZ5H4U5NLEkC8lBfJ450fMOm0Q1fgiFg+f2V3RF7FVz6y36ULHuFCVBzU/UKLbd9wsyD
1e8k4wFtUpOyEEcfm6JLAIYdlbvCqU10um7ePc6FMDdfyBrdF06IS2wLnFk4EdUiDbEf7xCab7nK
CYk0JJ5omcosGzZknx6KpPz03yjJjF9wuaJAqPGbVXSH8hC2CN7Ym1LjNbGRT8XzalL6F06aLG8j
YtIGcQ+6hEwJv7JTybdeTt2Y0KICGCWO6EAu9RQGNjAzDUhPGoESbXeViA+QFAfQvpwVXvsgu8JT
7qgmGl67UYSzhykVXmB2vXZt+5eH9sIlTd9j2tIn6Z9EflpX0ErWbh5aSUKB4t7pGUUiNxsafi5Q
Vn/0zZPFIvtbXSFOGyIz2aoJTDKwkIHFj8+rkGCGimv49DSmfuJJr8W9/bXrMijsgWq3F1mOdngB
xE7bhGiFzHeUHz+Jdv19JnnU32dcTtXmGvvs00+XfNU01wTCz3uMeHXT6IYJ1Nqjg+gTSrrhHZFn
/25LACBFerT2NsV2TN2NzmQn2a7WG1JMxWbRXSq1Iq2wT0iI1qaJZXEJsUW9AvKhBOdCdu/mp2gD
/oa0TMmURbUoGwoMkmCCXvzJTE/kDrLtrgKhD/WvptYI1H0jra6Bqp6Gl0qQ/SyYW3JcUF7Qr78E
iICgarjbMIEl3FwPQ7qvG2nJaEapfevsHXHKrCQHmKksk/iA9VovlVfYcfcl6GGBP6Zdwx1obXvu
w7HUayJhQYtT4ktjgUBV7AHMPOJCcC/iqBzW49WePm7UE4Ovtalf6Rm0O8sit89M1BsacgTJpBVg
bcdFgn+lGzGcXnzRhzoyP8/2ftG8pO0mM3XY8FgEaD6rp1pvQrm0+F7LZPvKim8Sbk91JBhNc5Sl
RwPBvP14MW7xOuEfRvTc8tOMsnPWWVAXdIgAIhvpjtQR3kRsnseVTVKKdf+PX7dCbQqxX1TGflrn
z9grf594rsizEBtRnWAAv3lckoYQ6n2cLYXlouDjV/H38go/KkwImtdc+7kezKZY9tbMdUd8lQPd
fcW9+Erc0C/ix/y83sWu+Of23mSka8s7XMphZFkc03i2g3yeJi32LPEAS+9b9Wmp97ULyHzzBYtJ
ku6GbzMIdm+GxBRicjRkzTd65f07xy0j8RQF80CJ2MXCXt5EqFx2OFNOhtMS0qaTNaI2iDvnse9S
PHktPfLRrJIfLylFjb3JOul+JPpJF3seJqetKYP2nOYKRGzy0vreld5Duu7z6sIzg6BEgiRmEYTB
2KKRlyyATtq1p5QiHbLDPvv8j+2PG+n/SD/I3vlVcifXLvrQvI23fkWzZGJ6wzuk9pbvrzq63Dr4
Jowq4YKZcUH22qLyhPNxBQkTZ6U7+XUI7TH+ezgeBv3xekeH4MNkY/oAnWyq8XGSpXHBf2LiXA1t
zv34y8n88mSudM0b13+AbQ4brfMT+AqP98BYL1cyntXJXQlzKr7H/2guoTEUtd/eQSQ0qi9Q18UX
tqq1BoAGKkPWOX+bMzJUp/odfP+wGBAgLGJgiIy4N94BcUndau8xoYc+OMLu+0zvPdeVXiijPEIx
VWKvWvW43iyDAeBjBqnGrpMENa7TUNEusyPBEXGLQZBYzJx+aTKJNhTkJKGnj+WQajKe6oQYx/7I
Gwx6sEy2lJk3nhPTL/TBW4NhWVLyGRd931wWzgrtLF0tFOO6fzje5jOZMrLQ+uKMPP8nB1nbunga
3cPfqDdZdjD8iPJvockUVRiEbre2RDaCkZIjSIDPa2ABAWtCNiu/nH0O0+AbsOGg75abyO3mkhHI
QVNPtQWxmJwXlV5IElnRnbwYQ0mn2E2i5P/ir2iqs6efUkJ24bfivN9G66KWSL+ZBaTqptkB5cV8
JOrk+0UlGuOS9bX73MVj+btWXpUpxVEtyOoQVpvt4+T9LpFMsvrqD/VeWjzN/Iq+7U8zaIS3FxJe
wCyhMfFti5+CCILqiMGdxe7BalMIs/m1Ph7vMAkMFHl8QkGRINEjVT7NthKIHTMen/ur85+UwTRz
Gx2NGE+OV9c7bv4kutDL7TccRI5sg7jl8UldMLqZPSgCE5qVjcTj26sidzQP7YKH+Y13nPkCeCje
27mBT8VhgQTH34XedXVsJ8holDoTuUTIQX5W/OwCmbLnUzm6d/4rGsGmDicLRHY+KesJhr/ejTW3
g6xtXD/Vnds20KbYT9Dr5TcexFaImGJHh5ATh2QfJvYnPEjiwlgUHkHUNQyIVDl7BNnCp9k9R5QP
cd7L58gvyqANmO08Yu01aOJe+i6CDA8sHn+0Cuye5Ty/yBQoiuIYV8ylk9hASJSVN2gr5FFxUtjz
sRDadbiDSJkTyDfoXzdSUL2oD14lbD6QQoqNNIb5Ez1JE66ttzJNVWE7bAJZxPLBO4IY2uiyEz6T
AtrOXhcOEAXzmWA97mFfg4Gu+LqjIUODwC7sJiBWWaLalT4w0So87DHrwrgQNSk+nq9Gf9x/QfD3
U7v7xaEVk6HD7VO4EIDdD0yJHEuWmhT7q7FxP78FptjfdbXNyxaIuhccS7pP1TluCyVvMQTzKnuD
Gdy8u6q8f+90u9ITAScD4y4M5pWdLCJO3QFzBYIfWehK1DztGCspyibEkrv4vIhqX7asCu0fY30h
QQ7Vs5uU6TyiRmTmffbK0+htcPtBZlBAXfXAt0bl8V1glKtTEuAKJ2AipgeoKHGvovG5YJgArkoq
+8yEDzeRqA4XMUnTZ815LmTa7pfq3lFTBiBx4Qd9EoJRrTz3d3X+iHnJ6StJHGigwS/9oMzGYk78
0qBDflfnRKgsO0AG029lvh/0nvNm7mvo9DzVKHRMtFneW2jFkkGVJezWHWKDxFiLxux2ny9bbTqV
I0ZbMENq0PEou1pGCNibb/ZvA1IoNN9vsJdtSiVLf99X585kvucEnclW1QejojLWTyNBAlWh6KJw
fJJpChBoEPhnfizNoV0AocGPG9heVjDv2ACaTRKX/DHwll9L1y0d7GW+gq+/cjFLnuhXvF9JZesQ
n8/rWpZBdxHHQH79fr9JsGkS6IT6Z15qDMaiUmJO8vI5YujER3OBkVvXzGkcM3AeM9hO8QQPdqwt
3+4DAMnTwoovCjD4XVuK4/GNz/peCIXxzcCescflQ61P0lm/OR1MtOv/0GWq1nyIcEPDoZXYpxpS
dHBIoL5YNocPFemG1zXFCnPvCScrga3FuqwRkDeG6vF3AhMSrwtpf7ckIcEIzZ+OpHtobo15DGxl
ffzycLHGcxMoFDYs3UxjE21ZpU+aoVKolMDhF+538+92U/ANvpJXP5oEAppCLQBmwJ94EtO+zGBC
1oA4hIHl0VVvbb+WZM+YwBZXn82IdJQCVH714HWovOsF2B6WfsWcDpfykobbukwMsVWyeNgCKJAn
nsJ9iiQB+Q+s34KiQm5XA5tb/0D3VJL1ldL8uJBEk54+Cv3SkwdeOmJBusfIOubNo8oyUN/EOcyW
Re9fqRTo0jyZG79tzGGweI/d2RfjxQuoKtMFhwMqm+bDcjkeUwq6m6dPTkdmTFTecE9i0EUuFKn9
77Mto1Rpayode7+F625ynSxA4q7qsousGqX2BdxyzclQodbMbl53zbwC97/mHvrFJ+zFU060f7MQ
8D2R2lHotzyK827kDcT8c/4J1beKu4sXouuUcyVlg3g/VLhcNHY9qEO1g0jDspqOJSlEzCGsMl8G
UkBitQTWtrigFHYADALsPTesLyTPFnVTMzM+gWxcKxX38aDauS8fZymyB+mVS5SUa4MLkgnsohsR
FpKJ870GalT5OV7wWPZ08kLVygvUWm5s7xs+RU4RgBi6KL45dGK/72RsV5TvO1Jv4BuzUbS+h7t8
8cSM52p3E7AllZuxc/+gmlXbdXUSQ1qhb/af3607dYOzj9kH7+SK7JQ4LxGnUBCQSiw+Ql2t+iv6
eqxl26sfWLVWG6Vai/dbOXGXHQhvOOeQL2FZcFwfX9YCbruueGtmSP1vKRD3sVj7XDmcPE900Tgv
p1YL/pRhQs/kjclnGqKHj8BZkiaY887cUGPNyP1Az8kWVtVVKIagwpyMQhuVwUoZJmd+UWN65Hlp
1da7/iVLnTlpbIE3XWG4qzQlVz+CMK8X+8/IOcRzO+ncaSCGU/o4ABoncVPV1S92xCqBfoLc8FoR
T8832tA6nQkB80UFs+UoN9nlRpj60GyQfKJdII+XKmLYIgQv7orOD4LoEYHPmmNTjXJm7pS+YT5q
vx70/23A36cP6uOrIrqh09zuroQMuX20Us86EwbN5q62ZuK2eX7wHJs2WaDdZQfNDIj4JlXUFeLv
/R2t9CtbtIV21OFeiiW0W9mmIuzOgaRX1J3OV2FxhT/Th85cKFoSsEI8UBhDlGZ5OPIq2EOCol1/
vTcY9OCiR/M9N8N1+SPVPHmU6alOooKGUf08jSbxpn0di5vzlnsLIRd6crEMnM/ugaGGgNt2iUwR
SyLwEpBfDHsNvOmYn73knemO0q5YJ/+jXgj4lYtMh7lTaZUabmM9YjpJMl8qfx69mqGR2CCHNjM2
MUtXgbQp8OPbCrqt43FxF1w61i+2w+0/j1aLw9FdFRAob8+PPy6OjF8wIMeEVEMXdqtWQX3VNjxV
Q5K3TkAXwe1S3BSBO/iRiduC3cYxScZVZsdKNlor+JkGDx7rg+6CGWffa/agxBlCE/9yKb6NprE6
AksVE8Em1ofBs3E8HvJQQLfysPmLeXTnppeg6rNsPgw8H/wK72b5A6h387g+Fl5XWV1kJ80rr2iz
SUo6FRfKudPFOTVfnT2y18o5Ux/n3RdqkMqxI3WEciZ4GTqb5sKb5W2mQFuxIbnFWtFun1h78JVY
KFpV5i62Wx5qOfESqD0mjQ4Z1PAkycV1DENlYuriDSC2NBfgNA4ztzCneFxaPuv+HSG12mb0Im28
OkIBxL+EveZwPtCNUE+xd9/5j42b56qvNFWS6SxVQNNmRllR2JM0ngd+QRw3PpYvwWkA7IwRvLFD
G2Zko5q0WIMBLfUEP3qxWejWirCxoHh7rXFoVPB1N38u/veF3JZKdH58CoF3FH1RJ0dDMrEHYNO3
kHSG7TBC71Rufa0dzkq8HIF58SXqHBBdiTYOzaRWyimph8nYJxuC+vKpNsFSIxs6S9+eojB0SO5T
qTyyvDtsMB3/v+fwnOZ156Qc27MVXyxPNJtmCNX7VdctMCX/Ey8gDo9r7/tW2iPfHE4yWGkML6aI
rcAvXIEB5buBjNlgYH0yt/oG1DTUrplRsQHvtsLR0iQLHjJCysWP+hYcmYEVp9THqaNOOHWTB4Jb
h0EOSnOT6y1uUFgmT8wLQomTsRzucvBOWTrEug0DvDg40FzZiUhpfF3ZpdW+0S1ktpQbDVKCdPUO
qCg+plvBRVKFHZLXlRplNetA5Rwhqngh5jdC33/d/feePfCWBLhxMJ+SqwB95WEU/joNcluTnSFe
YahdUhOmAGgXYprNoknYoeG+dpnMGVCEFwQX/oove0A/rRA1TbPL/L4WVww100RklYp8snvN94uW
DXO1NpyrTV6YSESpbyJQNHfYyNbTyPoll55UjYYykiC7A7tN0HzVdXGP9l09KMK9XN/YRPCkvB3I
q0HUbmQBxe3AlgwHKzSx1TrnayQYIXCy8lN1Ee0jnBRd16Kipozs23VeyrGp7YvW+SQsf0citrzD
lg7ABCfzcNgxOtFK7pKkhHgQ80hlrQrX9bx4Zk4poxzZzOSphRwaBoexEfbZeZV6PPIiB+awU+gM
J2R6wwkDuX/iD36S1x0BLBxuRghBwnIEN0Dzoa/sGupapcTA+/oqY8jIrZIFFf5vfc1qtgKgHCxC
B7M1TtsAIzNAHRjMnCQTsUPvE5VUjLqV43JxseT0ueIco8HzPcM4eoLd9NBoMQ5nCiVGJOobyNYv
tz5FnvlaiXpQCA4Zt5eEVlsbcWY9oJY4K8Uo7/kr3HL8AS0AQeO9uQBxAQNebPZJon5Y2MWmGlkg
iKhNQ07Exw+i/+Q37Qlq/P8YTYqT6CuKUPKVJZ4av1o7lFOgnjGbWnv9DjerM1fgma48qU8baldx
IJXDp31h7qQR/xlrncZsBI4uGjXkR8p4CbJtjgLyM9+vjMh+7zRlOjYU9cSs4CJXo5nmyBeG/QHp
6vZB3KByjtg3mKtSXjreRSWgsD3+mqAqigS8AviszHbZ1Ppd9bAMgzf7iIzmf9uwLLt8J65n9RTi
INneGdDbjYUeRrsZPaCLYHqjNEqepzDQ4eRaVMOdlW33q4qEC97RrOEVPoQguVX/kGP1Do93Dfmz
wA/pYDsqTWYY2n2nrBbNydEpmqDYyNI+dad3mXnyGItrHNZrp9fQjeX4Lgt53L2oL3Qale/p8tX9
vM/xJqhwTwzexE1GmmN7elWsmYIbTwumcwjliP3iUQkYDl1EaXk83UuGZMJ32WF45dxnHTXkaSV1
Zx4XvgAbhw/Fsy4WyKTx4B/VpXAq1Wh3RLrK+uO0dge4zSqee/fTY1ftvp4eYYOzisSX5D7M+lNg
3s6NWgnsmeP+KY17SZAfuFMmDcg2gAsHJKAHLAvHD/yIDp90AmkZHWt/2cz2noIAtkSd8h05DegB
1yuqUkUpnYGjzmnsPySbNUlWJ+7q6UxAVrDTqPDiITfkNlGW1cFjU16P0W+bgk7S6Mlx32bJ9n9d
6iqCC21bsj1esJqUsraijHD4lqn+flLgmFGJscTNTZZt/qHQQV9Hu+p3sm37VfxE6489K/uzP+vy
11NAF0K1LLHmiTpuFbAOqeQ/0cHmOejtLhP+S945qBNaiJrGVknC+eTBAranDKqK5Rr/vrAAylva
YIPj+UvfMnLbJGcpKW4YH5Wz6GzBl1HzHjXX2PEp4SrhgVjvcmEspfkViG3tIgu6XT+gWs3VohtP
Iwb2er84OGdVIoYQAEnEDWtzl0hoPeV16ZUt5U/uWEucyMpHQdcAAD6fK2AyPKuZJ6Ar+GoWR6d/
/StBGFEwXz1PcKB8llv8aXKXiG+WTecoHNY1OWTgAlM3wIqNhCiME+bz5um3n6F/yZ1vAx5PMlIn
00cPadDEmpblu9tbV+QDeclbOG1rdFszYiR1Wn+mj10di11gKskhPtj5Faez4lVDGQy36vLHJWwm
NYWL8P6kiTwmLDsiUW4s/RiEPeVNEtPMWluyQrKiXBqlOEr0G+XfjJ4IhrDKD5nDIsZlrd5nYszB
wbkvOiM5MH/XKtkvJfhJ3MG8ONVb3sAqk+cvWuwBflLGBRYaqskn2O85277q5r1aB5J74iZ9FsTa
I9Ri/6Bk257wdLerXDcW1AfOudACtSUPPhAWWF2g6dT2RYYqaOTUq/tL33oBQ6E1eRjETy6Woyxu
NHBO/PUKbl4MtJMfH4M1Fid/0smAg5WWYXnlTmtzAtaQlaOfoTQmlhNKI1k7m5KM1PPNInlAXzTI
ReHHSeMbw4OWrD8jZN2uEFQKlwmaM/OyfZRJMGaK4Oupep28yIGyOxz8HswwOTHCIfZNdZyaUP8B
kMraGNtE8uyMc63xTCrdRBzNm6bACWlMrge4alYRJUhg9yZ4TyvrCBu+zLa39HoOCt57Dtvfz2ZD
MuZd3nafcf2oy/iXgTpbTeTisSHb3oxXi72Wm3xgpZQKMz0iX0Y1N/9JGcxh9mvEuDLn+OqRpAXB
WXQYsBrySYrF46n9nZnkgJh9gzmqd9x4QX0tGdGAsD972J8hF5Ba2eoVstIUSKBg94/9RepzLrLs
y1nO9ivRJp63D5B0Is9ZD62fbHMoShjnbf6+eSgpId+Yeq+N6l64p5SkbwDjMTHUMpql//4UVhTN
1VhpBY33CBBqRCcRIYwsj9tj2n7TnySzAH610DLZ5fPXL/2tfiQc87aA+7+F1ZQ+4jVZmSh+aOE3
HguxvqrGkn//yGf5AXgzRSW5p3lPilZXq6U1MKRaJJJoE2ET6Z+EIyVzKHSbpHCAYY9ZfdyPTs0D
nHFWm4iGZGmfh9nbKvMGjQggODJ/xg6QQdqaJYc4qVac4pDt9yRMLHIru82Dy/ZOmH5BWCUop7lC
ABAuhjdzZ9xC1EV5tQCSReWEc2rFHz4PKTRely//fYJ+isMzrVOOnWfXU30neH1pFr7iXWVvSWx6
2t1mOJDv61j+ToR5zkjbIyU32kH2925sJNloG1JAU6Hp5B0ohRcAbJzvcpq0ROSqwS3fchLdDAE7
JoxtK7smc6fUPOxpr8rpWT00gbwYZ9Mxu9yEB/627KPRmAFkl6vNB7YiyTYF+iHlPdHMQWFo79WY
UFLq/OPsP5PRddbyTJzG99/CSFfhfO9VJYhaiYm2yGC/lDbm6Y8wBJUKHQH9SJw8dbC6UjfRUgln
2Isx8RLoAYO/ywZScEr0k4j1+kgdXUm8kncdwbn3xGe+LBAW1yvYg04eFg5N8iDp9iSzOeQTmj1V
iW5II1G97gjNOlUq9ukm+G3lG9NfwxvoCDNVMCVgDdKewf5k7gbNVE3RbJARX7iBdaZPnMMXOgT9
1iSdQsZzAUbPXzmwnXqJi0/FXdq8Rbu9dyjm+yC8qdluIVKKVaduBFHof8CyffsXDdcC6xdNO08L
0WfjKcoD64VURu6PzkXtZuhN8RDHq1AO2079ZoII8+v72d/15Ik/DHLfaqhM+bGhVV/dmAwjDHdG
1lqT8p6uRtTxbR0SC166wMRMmwFYRjdlRvVO7rJTTZB3yekzE4FaoaSjvE5ddzO1NOhNkJzbl8jh
Emx2L1Ow+CBGpO0FlFhrPslbdIDSeTSSVCowOfFNuf6Po9SOCbn7hySr/BtmARffYDLGkdKudsPl
cY2Icw/weufSv0oTuZuIpr5eSfxy7jMIbdOXZ0c/zE9BBXWVnMKwcqyOvZ3vxqrGZquDOL8Q2pcn
jhE/iokPF4KpKpx6SL9QtRfc0f6yoTPCAUHhb6DDKD0A9GE+h09cLDM43t8CBVJTQ+0q9ZFkufap
p5JXOp/+X7FskcOv/JjHNJgM5pi9JTF1Wm6QS/z5wLfXbvkLhOh0v5VdeRsh2YTwUv3GMSgrJEG8
OfUKtW1zfz+l1Ku+Jg/hu69TFxoacC8fvRkD2qrDnS6gkOwhMGOLYOLCOiXJqs4tyyajPX1+bbBn
TLesn/bT0W2zrogW8oDIz2TmpGlBFoETKueEpIpu1kTJ7ggkuBGMPbC50X75DDcg0rM9Mog7Br6J
4OH/YAJcRcTuH2mzHSp4onqJEupa2HKBNrsvBPwu7GsjXOt9jp3VsIt+jYoVs7W7F7WxYNMKTwp8
zN3H2iIj2EO/S1XiPyW57LyrIc3AxXHd+nFH2uDsq2MPn5UHFauLwJ8JzI71ZgHhmU7nDKAyCD1d
hXqpfTxhW1WpqCsp4y/9vOX9Ht6GvqrINQvwHtrvp3cfhQ9PR4TTANtFezz016A+jKMq1o3d3Dkk
oABQ6YwWASvQh49EmX2Ehi9acBRVJjw0ff2iM7265BJoyWAtfWX5SYCXIqPbUCBnX6K2wEyxdNQ1
o3vWI7u7FNcp5GGYkNg1Ds7TCKaTJDAqa9lKotwcBURMmwlF/Z92RGkq8X5uxJkYkKhn8V1clk4N
NdtXt/YQeF2GCK2c2dmJ4IMuiLQmqMQNjh1s1vnCCrEZmTlkWwqLbCFEjCYVrnk9cM4vuZfjl4d/
i/Ky1iA+T7Xu1jf12qisHvrS2Vbj4nnb8xCrva4ll4D5e/ZX41FvOgwdSZVVCBTBlOuDdRtuXH2K
zvmd6qpsfIMwY3bNLo2S+rRcP0UF0Fu8AYhRdim9PhR72U++Gd94ot85l8jySMpI0PoXXyvtNMml
wQZrfJok+TY+adUs/JCIHhleLUdo8KKUeutX78of1viyja/lgGpQbVt2b1/+9sbxtHXVxRKzWHjd
vZQLV2yCq5XyiTMHcxBWyKq6xyIc+ON2pCmockCRuA5usw8VgHjNrOfMhzaU+QOrU8Ru9EZ3/BLW
4B+lia0Gk5CTXy3KNlQpFOOjMuZY1fRyjVGFYShwcGX/NBNA6vQL2zSumgQxyjpjmGLfkbCzKS8i
2Rb6pXhqYY8CbqwR3WODIyDoNs6PtYBZgKCxrQ6QANhZ1A+gQZX0tDTRolGS964JlIkhSvJ99e4M
zAybuHSpK+eoeiy2qX2ghERyJgodpZXxkXycV8u/uUfzL2lqXl0rxrbsi4BAjKsCnGikpOD/dMBP
cenrNzz5ZfXvX/HeyQG/qHEq6/zOGxU/CoCZ0vsZsGkNyJU0EVi3KzwXpNvzS1AwlXKEaFgRJ7IT
i2k+a5C/5oUwNXiq4YD8FWTfjCpSPymyU25i/ow867ESr0gtlug85s9D5wNaOo5HUgIv88FednTC
5VltuV0CfqpoJWzWa2OhJf8ybtHegwdLDwFEg9YkV9tfdZIBt0Xb6refGHz1X2HnQs5rz7fWjFAI
s7vUk7stQacKg5RS1Cn25LR/+VX1watdglyXENAXYVGhMLMTMxOaG6tsr+1nAAvRntiny7iA9lJ/
9fw/UR2w64ooW3fEuF7hqj1GzeofFxFnJzlbHfc8l24g/QNaSqzj2Q48zojlTvGZdhJ1LGa50dMK
A2aH6voOzquC7PNfKV+pJLS1n24igEgk8m3/fexOQC9h73tsI8AujLbTBs+Op3HtSlf8V/OHlXnu
CUIvTJOw6H+Tcg5DIONHJGIYRezuque2XHYSOBUg6RHiUMnfDf62Xr76GMXXkC0vfdY0GK2eExoU
tvtesVMBpaBEnIhEkgWQLE+MQknA5IeonQVy05JTaBuXjpFPXqik77vUlPnlpXvdXCQG0XN/Sn3Y
H5Xz6pHWlsw64li4HV2EP+b9NfE2ImfwPZsv2hrLMKfOb2KW/K8F6S7yTphB2qCV1DJKzME11ZPw
NOhB66EpHzveMEijyYlhjzyNJTaURpipNQ2Z9yFVyONVR1lPQLT/xuIXXTcnpfcLw9EjRP5JGow7
XiVahs25zn3PeGcnd/0nnpXCF4K+lzTnWul7aZCbSTYc146XP9HijsM4BXlKc/Eqqe0X4LNZcc6+
H1twy3IRUxWKDhc5x9DggrLjisUsfVF9iDzBjMU7ZE8z6vUxz4REL+O1QNeWRaE/NGkqz921VOO7
OuhA/JgbKXWRR7YJj2yafFEft6TDAEglxHOM+pljNemsmJjTGcsnoKVCU47HAxZWOJ4P40LgmVbl
DI5mHBgZdaIi9vRYGo2EQQJAvgZZY5JhOjzkYHqqsub586HJN6HFf34PTTJsvMcC7ZiVx9Ex7gXs
2t9YT+XI8uMVQd13ULXkpRhcBG4j/uEYoH0cT9FgHurjr6yfvLzK8YqQ5scqX3IZZ1VqTmy2R5AD
6HllOoilD0TclT/LErivf32I+Y4JRtWJbC9V7zSlO3OEG2nSUjJhwNyMnMOHlQoPrNglxCgXtfC4
htHUpjj6JaG7iwLE/aKSJuIKLyhTwkMnsLMXDvz21YY9o8qomNX530U5v8WudhJkZpPYRKs5SbMp
g62UzSF03DGJ2dFPAuBih41CLg2lAYGUuMc1D076s/qPGlkGadOsqZCW6l0KowuT3mOQc5PAxRkE
AeVw8sWO4rsXIwQHfYnBrQTGa+p/rNcddcVqQezjXuAweAiE6VSRs897z9c4G4O1LAIZY/zXsnny
1vSKbf2mBsxs41gqE3R72chL4gJJmmZjPrcVAM8IJX4zNBWHfRESn2dI89n6IdjpUH6gYBaufaI6
wRikghSd0cQr+zL82UcgfVTBh+Za4FENcd3QtDzzpyv7kppGhToIG4tYd9QXmj8+LT+CiDeVkBiz
ssE8M1aL8iZu/9ed+SOP+Mk4ilo7CELsxKhcr6hS+RlldgNqjVKuVtPJ3or71RbMmXNpW1vEd6CV
3s57Q3Zi3a5HkDEp5LkoRPVcjPhmuJ6oSs1mxt3R/uhwuINuKE31vw+MRRGt9AXaVbJwqtwpusrz
sBamSdp58rx3AtH7SelVDmWE/NiFd/WLSl+0k4u4QdsNRMEnKtzP/MAd+Netu6H4USEMgz7HNdt3
xYb2DZjqOKxmwZpqj0InnSGPeOzILrkrmLG/8D19ZN+HyO4agmAvebMdJPxPUswR4I8XUQF2RlLG
gZRouzBaZLcXjMdzJ1Ha43fOvtenvInPL5sJiEA40WA/HGIl3A7cWHY97aN6b6V3m1BzeP1gXsaP
7StaxAy6pAAGl30g6pz63pfOPfjTdJV5JS/jwklVm0K2Sxivey8xvhAXPUpoyqO7eOR1RKLtJfAF
CmUyJci/DzesIfLcKxD+3Q9xoQMavFYTLXy8h8tBflUy+214DLBk84cSapEh5iN8H4VaYQHbRPt0
LcK3fssSRVHmtPTXIxxzq1r7n0b9bzaJQUvoZSbksoKudfY4ZJplc0J1tPSInHhJX+qPlsHH6yKV
AMXQa+Geusp9ykJ6HpHW8cIFP1rFZdEuVphjMr9MfzY9xgukgyAw/HmrIZqxGIde2b/i7y0KjGwO
Sezs1pdu/h2h98Dlwi29HwyLLV0tFltdxYTqc6fqsW7SyDJ6bsA7l3nbqqLu7mvoSWyFFgi2os/6
duiriMdRK0aYq9mgq9Jw1vR8qnbr3jHdTIC+OHbDninAUYSLsvrpy5IwzH3LvZz1GdmcG9ApNZyK
3DCq+pOqTSaHUjieeZ3X1epdT3FStjqNe8U2mqkGRxt8CBRodtecwm2EzW3DF99nlR0YMPco1wZf
0J4zmIiObuJaE9Gte+gpbYB0NPFExruRbA9nl0n5YaGbgCNY1pFSdk6bwqfGoNiyzJpwhYM/KDxp
HLMh1vn42Qmo5lJEgTe9HTUCEUxce0Mqhd1sRR9Z8lDtkQJmsvFNENVb+ou5kBJmGZDIjn7nRRp2
A/eMaivvi+5ec3ebGg/YHBupLdFB3OxyoRUiKNRYG/REBZ2fIjGNN6HY+ZkGkc582Pt60vfryTcS
uHd0DdXV6Of8zm/KpCFQoARBaRyuMk13//qxd+0q3ffrL2apO0XL8u2fZ5EvNf6s9sIDbZUusyWC
hioG60iXX1hVm6/L+SQ4n8AcYkCgIfiNpGeNJDNrro/vDFPs65dyOjoUC+Wvn1atJSF2NbV+YmUa
oHoJyATezbM9g5ghhjtU1rx0rJbVICjeN9D+4CIQK+idn2E49MZbCD2pfjidCU4AYBhjrrC5JOTs
L5GLh0Tkteb/QBSQMMMMronN3phoubyuDQnEvAcyMAERhpQN5f6M5TVwyRRwTUJjKjNAvaspMgFe
nTGBQTH1VVaw1B1tYZKuHaB/svEGflLX2PFHXFpB/ntlfbo8FcDSi8ZiKtKQDF+t6yBxSMqb3PmI
eiROwT2ab2udljx3TXxNu+UPyUBF9F6lRd8lAGNVRqD/cdd4V4B1VkmXja+1qFL9zlVqCWe8DZ2j
x/xjNYhCB9w4f0mwfB6QRVsGYDcgbifFhZ+b+ijKNRCUcm7/Wf2yE5gXQ8LWL296jEC0sV/Ug1Cz
etTk6sCoR59Y+7gTzhebYME5MXoeTwZX4s7FE3XDQv4AfYHtVIczUq/AqZMfHGuxIzLRUUHAy4hY
h8elXrF3T9TFBzG93f+YZj9cPVHSWAkWyFlzKjGE8/Z/KDJlL4rJpGoXz0+V2R1T/ejk2BNp3i7y
8xBVy9GX5r2spCuq99FMC+JE4CHxowbAT7lcwI0yBgKL44L2jdZYQGpKFVz3xR5og24Lss389yMG
fIsGjg6bumwRYAahlf0XVJjdusHwQqLPgk/a6ZU4MXGFS0sL4+a1XNub7ZJyh7SNfMkjsMY9daVB
uWTMuFz89TPr6HcMNNjYtJbqoyvlNWYeK3t2fU3FMP6+FY+34hmHK9mHAQ+CEZxGFs5ijvtbD5R8
rODTB2QttzUO8wTxMmdMqfUIG6/OQ82zfH5wSLN0sQ/ArKf9p2E+DwITSjtxvyYjZUZH9cmGgRjy
XUth1T99PWaeObt1M+k6LRlJ+F2AdlrS7fbm+2jfc7Zg5K02dxam+7LuJ0yqa985nl+mkcXzz4Nr
UiMV1qDUH9YsADgp4xLTu6RGRVsXRKxgSx9E1mA7nymMHRzbPma+/zeBzo2YNPEbwsSm98RCH6oc
ESJSQAsQGnwT2g8Q4jEKRWQRd8e4LcmHtlsjrCCilGp03VitQDgY/qKSrocpbTL29ynkJl6HAEZR
gOgixaIJn78/awwCH51vDHBEiiVJ0JXtURQiLfRcRSBoSaD5EVD+KwnLAFK2uj1YW8xpq0yvvZus
vAu9B5O9sZBqeAz5JgsjyLv3p1Pqzuwyd99ignbyxkAhXVOeZLhgTJbwmZ8NChYtBdx9iKs7WLr6
S9XBrXs0rNo27oelx4U9VA4sa2lEjWLaBkTeDd/jO6PasoPVuglYCYx93v8ioxawEDQw0nKT+cYs
1XTCSX4J5UQ6PlGVVPW4sgiXpUMaGPU2JTGlgJSLlKkLZKxeJCrTuRCWr1CcmgR1GcFuTWcE2Xgq
nReEiy7dPf10CjV4C9ebkdRESb77Zlwgd+TvgPTHwB8fbAk8MZQPXZbRIS7TgmmLYS3+Z8ZMeoXI
gCoFqDY3cRSBhxBJ+mP+7OqS7wGV4UynGM+6WE83COMmg54/kYRrkugtr5p7qUE5m3Pq4uhUicLc
8HIq1S/1hd/AE5T5PTpwpGmB0ZMUJB42oYUNrCHzbUq5RQlbWHtrmejtfejX2XpJQgI40ypcZ+nG
Ze9jo1ao5ta29fVU8WZx9ILg5XSkrMuZyk2QnGBGi7JQ8L0Uql9m69Y+JPLE+USqG5r3iFNIzUh/
Cx4wI+Y8was0uHOwRIF9IcIQKDLNz17WadtHsMcQtbjRWluuKJiRjgfzz2T6tIE4aAECb5MrKXKN
kk5lbLTGFquxA+Qbd62LgILUqWCNrdJn5HEt88LnNUNj7KzoQpKQerPrT4kafOIsKaekVEScXw3S
1aiP98+zdp1dfjf8lQeDBlRVHKxTW/EUe96rwYerr3m/4ccBKJYRDlrqg2hwVbyqr0kukAT4Nb4f
7tOF139BPnWO1xF8VMDSzg2ttrJHB3xKlnmJ9VIJir4msxivS4QNxdo8VOr767wN6gF+sAOQTz9W
ZCysFDj0RZWJeCUXUpjaIkQLPUdSbB5tSpIXdLXciEUs6qLXknMotg/R0wJQYPC3noMR+p61HWa1
TqshTlRPRMvbnx/tXH9o842RLKSiO0UcANbYlm7j3ta0pegQlflAsQWhcyWXJtMp3/RFA5kZXcg2
coqliQiSilqiNgBO9BgVTtsc9ycdT+BCqnOTs0nlLGuGuJxEIlXIur0WvJdJC2ljZLu0Ze7T2ExP
zXmScwmfLT9x6D5xIT4/Iu//cDovcDW/cnWXpxodesi+6Z83QPWW9Gj+MEbe731HAcqTFkEYyd88
q/sZuo+ErDUdujaiaW7tBGRoLtlW4U85MFUXCHt4WMCFSwvAA5gJOlrDdS2XRlpA8Iw9ALYwtIWe
aBfogv4WMP+sT/o+3nPMvsCJXK11SVOgcmargfxSNnVwNDmwvmk2T1+42jT5n/ZKgHVpcoNKwBJK
QOScfOj3j/PeKMTQRj4u72pUBHx0Ngl0xadTId4bx8DPLDf8AOB1gT8kDxU2OTikEZm1HHHzKOo1
ar0em6sLZ6rtbjmOloAsczqhPN7+GGtZhNOYahWRzjrBrbMOR+CwUAUCORhVWAPLZ9w2fVsxMUzp
vPPiJxeuWzisUiltV64IuNFFee9LbSjkGADy2zXiOlUOinhb3D8RBLK7jlX/RL2JQ8DzFsOZ4kaa
3G9KUItzE+F2G3VAUpY+EddQrAf0ju1CTneY3MBP7hj039wABoCLpQNd9gHkR2crcRlIRDLsxuRP
HfXmnwpTcR9Yf6Qk0bCHftlF15yRfAu5MsOkUIfMaC1D+b56j+2XAaBoFJFl2TkmPnJZZ5bVcl2S
AH4A2kxbctJ/42ksCWH50CJ1hYQuJKQ0VQmcKP5k4VnJTGIa2PZJ6nmCJwNOGfy4SD7bKSfy8Zq6
TZbF0qFOLEFmSXMggbykgMNiNos/45xN2MyfQ30ju4o+Ym91t1R2VAit46J9wThNQ4nqvm4ssErV
uWzB0kEIdGGkdJOjWf0M0bzhEO72q4G7lSgkVorkxEUgT/YVUI3LOYXVvkSx7lVuc7KPiArQjgtl
2lWwjv1eyHXOb23gIu9EnBIhTuMjGhODw1CmKioSvYAH0xcPnOYF4mH4aQgU0ODukPvoHoR/tawU
5qLqUblL8RNu+pkeLFPFuBVpYKoIrVKs7IH7BPQCrPH1WOQQtCMfaIe0ZySuaQu8lMBffP/jEpYW
4hMOP0EARfbua2pfJWZs8ctq/x9rsnuziPrcn2eX81MGLPI3x0WuPd4/xzvFAIEldqfK3QlQBUi0
J8pJ0PVn8a+961zSgTKZiDJKHPoTzHQNUWqjhbg/KnOMced4MsMew1/A4dch85+mfIigaLvjzXO5
x0iNKcpTcbV5k9ey1mzAk1WRlKqmCCPENtIw5CNrKDxtfs467rPpf2uLsrmIMNY30KAAGaEulxxy
kA5fX46XkQVIP0gxEWE6f0GMa4NmthBu3v5kKSlOg3rnvU1zovG15dGUCU5nyjSOLO+1N8x1lOiu
7Ex67UzbOqN7bAErD5czwkeHVHf6gKWW8y3Daz0yJd/MoEn8zn8Vo2l/BrWGoH6CmgGmGRMQ2e+n
yiW+08NuJGUL+weOxIdE/z4swHQuqOvQLrJ1cFw63PFspXVBvz1GKaI5/XgqRGC9jFytmLM8KRG8
iDPJTUiw9B6ivaimSt3rx63whYVxHgDHWZnRVinDmXyGdcLjTAvV2zhYyi+104iSLDr+A50mS3e3
IUa/yxWrXXeYVpTuoUSKMytiu2Nya5UXWLuwRAxgHZf6N/E7Gj0V5XB+3zb483mURqi2OZPcXrIW
WHnE2UQ+zTvbtnLWSMoP1ogEHsXcl9C6UgZ5TGjIrVkfFP6kgohmcp54ueoU0n6bDRfHFeMibBU1
TFns8ZXf/2rGk2aOlvpaHb+WUDwNfQaDoeS5ZA2A1jM9/+f2DGRSE2A4NTg+0qMnPjjlNQ0+4FPd
TYSCsli9RispBZsKnqULmOl3/+nqucBH+lYIwihxPDUdm67ezNppKDDGpODSeqotqJGBfTxOxaOu
Q2Fe4iMe7HO+2lw/ttx1tYbg5NMDzQemEJStNW/iEyZrpLeUBICS02mFEYpJbotuAp3/Q+c3OspN
Tp2zU6e+ZOHNHojjp1GHIBz8hX+0ZUD/yDhKO2cIjl7HwRU1wNxYX/2aFRQY2jgS6gtIUDiq3Jnp
QXA1XhEATh9k8k7EOgbJ9avBW8SAH60Rn6Yrgd5G4qOaLoF7fP9rSujGmxNkIAIZ38sJySoA5Ni+
aaTMTQTloFJKXnzRsXy5lui2z72ncG4/ynZ8LwsLEK8j1jHolvAXIWQvnJwohS/HonAUSI0ReR7+
mTQaFtPSor92xM7THX1vSWAiLTgYQcg3gqE5IJmWO1dEigYka6qmo6AaA76Id6R9+uSQ0hQbrkPL
lLTgDHnJmtdkVqEuVfFW3LaLzjliB+yuaOFc5zVdZqtMad2zi2AGdb6fV7UwykTq3UaDz+1SKmxq
WxVZyKVYxJqqrRT2UfKiYChUccUpADHsJF884eRyImGK+79IC3th3IPTUtI1Yb+NwHKYegK0SJxH
0jQ3jHr7fh+XfPur3kNWFkoozp3rKxmGBbbTDPWqvDnLUGcZzzfrWy1rQrM3Ra/udlMWmFmg3aaw
o9+xE94LelpQ2x+tDcBqShZfaitkPoyVt3+XPAU5DF7EvcQhfhuEVKp7FyUuzAlzxshC7NmxYjcT
Te2XTzKhTpLfotLHx6bhy5zCMGudE8C0Q7GvXJ8KRWGzR3I6InET25q9t9CCS4dFeV6HxZZl7jGb
vUegZ5keAeo+x4Ei6/j/Oodaii2Mi2Q9JnwkGQeoC4/1I9ML4Zs3Be9UigBaOgQbuwnbbZGjEFg6
VljsN87F5QtR5h2uhhf5UR+0GppQSxrXeuOAoNWRlaqaPQM9G8AlPOkTOAJzOr2TJikAAm6NwOh/
/gGr/ou6f7q4JC5MA/Iv4I0mh7wMyd9Ot8WAUxBvEsowgV/8Fp3y8xRr+8og1Zs1Hixbs0zsvPR2
L9QziIjFxjokSTlBZVCs4eckBAvsflNnwILQ2P1ZnGC3Mv2bM3n/CKFSoYgOlg2J49HpPlHgcZar
66z93BqDAyzK4s38kiFh4oU9EkD4aieWguQ1tuDwkzxwJNu9dpKa2+YqNXNRaqXDhnY8Kvd5+hiB
LPKkmjDXYqqIb1WHJesvqodKRBqvpG3xD9DNIPX5l4sHZwucZi6EuuMGfDQBFmWTpqqkMxadaDzf
ps0WytBHb7HJI0O8gMFzqgLUwskaMODFLAYQDip1UANxMCDoYEp9Ll7cXidvIu3dRz5liGlXBLUi
kHAXQRIV4PcQIkf8WfOvtI7qeLng0V7QGTfj29XWN+kCzjuLYH7nu/offa9UWfdxnbXKTgMx7n2K
oE07Ox/ngF84XLIHLY13kGQcm2JrtNKIE6f46YwKjI26BxCgXm6ajlC/8SYSR1dO6tqsSgtPM37m
G5hxITc5c3t9gWIl5OJ51YgafF6wSkvFvCxl+0kORLK9487UwZG32OYBtMtgY7XYkXbTZNqoxpao
2f4XtY5pDz4rKH/4jTp1u3SRWx0M2jpfJHhVjJBb3Q82686+CJZ3BxazQRV4XpLxDuGK2tXh2wAD
Bru/KljYhez7BGUK7R0wXo+rPBVvCo4Wop4ZkrdpVqQlk7jUt/9Dy0QjOe2/tYSi2yxU09gU1CIA
IxlsAvcAPE4sLmJluaSCpIN32c6GCgeYSS3vTPSgsaWBBajK1gCm9bJ9TqESPgMFCLnSuxfxYtTq
c5GWOQOX0ULfEJtD1fLmI110AcED4XtNGyAXWkSfAyR3t0MkhI75ODXqmrvHjYIUcIVMch9+QHDA
vunYHtNxeSshgsbLLFVuy+GVkuEgIGDkm2mRKqtujOHcWPE1iL6bXAbSYQa+jR3Iz3PUj+9zyoct
GJDzHEUMSQTmO767XLQA2wG/XpAZTBOxicX3EaMNG63pIgRojrv+741HR2uUeEJJwnLx5C/VNDlR
WPJDuQBC1Q6DhXpU7gBz0sL78awunpkZLf94DIuu+o6yf8cu6xPS8zsM3cyLE6lco5EOeY9UfiMm
WzZRxjhyGtO698+gypcXTCzWaAuX564A1kPAC0SehmekACgJykkKsLE0oFo8OKoZGKfP1dvQ7n3r
jcE/ZQ3S+T3X0JzTFU+fnWyF7eSC/+KECJcCKFOhyNs7forD8C3LDiivjMsi8Sss+S+wIdkFtoGw
c9ZeICTjfrsVTrAzijCkDqqvuCIJ4lMmBRQ/RbMv+tg9h3/g1CDn15gLfMN6j1UXNAvhQsKL0xf3
SeAa2/5yi7TlvoJQqXvs0TUmFd4aLasLTJkmbhrhQG4yZnJ9uMgH7/kIRT2VufpT8YZNWpv4ejNX
yAZTyGH1FbHCFqPvGDMcyPKGsIuo1IM9Qivxw/M0HNta7d2SvINNNshDPamHg4SM0Kxo9BiYEjeE
81+7Z+O4ZCGHsgvUgooA4bopQP5GJmcxc+GjjG9tBu+MkVYziSAJkIyHODfs7pmYGluBt90tAnM0
9wwoKBJxZDtbhralUXU9KFcczHKhxFK7BSTFfmDXya9CfnmMce6pbs1kz7tPho0l+YpfZSEOs264
+/r+tR5RKAelG2lUCB1wY7LWnl263cHLfXNzKe/Rr87NpGs1h7nJVeR8kz+4FJVrNg8snaFVgLl1
fMoWr6K9ij7FtCSxZGOL+S29x0DVCeLv72SxG8exQgtSOpxsNKvwo+CbMap4YBV8/GCF361eKc/X
70iVlBH9fLMNVYUU5LV5CQ0MztwwkoeLjDo7Xxw+rCWHBwKl+J0UwDI1qXpO1TL9NpUVajaHAu6G
CszC5eU9WPwsDVsIE9C0ts0PJlVne9/883WUP6S0Zi1Une9zYHQL4SYtQTQBiBFVXemgXeiPQyGs
N1Nx6Li6nGMGAWH8BflQoM750kJmbJ/SJ4mKsPYNKnf5n3HWj5kQ6+vkmE3Cz42F1oBlkn7glIGG
QQzh4TUsLsB4sanmkjs2vEw2Fi4SnsmtIeG+NyoF5W6PS19kFk1BZOB3HOvuDHW9Ay4qPdQG5vNX
REmIQ5DRxYsWJ2oSMyPWw0lkewpYPVHsIUCApTxmP9XEd/aUhOHZz++wdXuCQxk/VH9YdgLbx+4K
muzO154uEaJKioWCfQtCao0Av/gLSmmS3D9nqoEsPOBL3Vut/vb0YiBFVHK26zQWJshTrxWGwYMl
vPNlQzWJAbfkQ4wJ1uD0j/0FZod8vI1Xn5U8FpIyB0Dcwu+gWRSZx4AEVROc9KdfndfM2dRlCPwu
tmWS9YlaJ3kS14Vnca7uFCXuk1oF2jv1sM7b5UAbSZPht0BIf0CV1xZJbZ5tbaokNLLC78rmLDE/
qBjY6NW6C4s7a/apVY7RTeWABo6Ok29ULnq8XHKoUT6lxCWM/ffw0CksBAuxWjLs/rZLDYMb/oDT
lSytmGx6t8RLeLKHElGk0HJCljv8iUj6/M8ue6rCzgZplyk7RSrXu/2Z6rXSBUvDaOddsshF1sTO
fGN1F3I3kgGiM3PNLUWBBUJSGTF5BjBs9CKgGMjdf97aMp/Bh0IVkUeU+F1UPR6U06OBKnVUu8Cv
gNRi2eDj3e6HKxPJKdRb5dq8vFmxsnjFpawh4EplGLJfYv22bIhEy+mawGMiHIh3GTzmPrxwlrYB
gtVUjd4720HNWsgszZt1rTHhpphiLjsOC6+qfNTDgYivgXckSCc9st8uodZ1as7sPFLwjV7/TpqO
NJPD7bCnu8FT5BeXENohtnjTvP/xSM+AMG1XsLhXDS0A+xeu8bZpIsd73RaIZeTxgBOgk3CvyEid
UPAs2Ajv373P20NUBvgXJLOzYrKNdgVBkvgWZFosq3/eGxKg+7HdpJNl6WGEabk8xqA5jh47Vgum
9lFx2Z2jOgTyqegzvUaFYewn0auFD08uL/2svLo4ncctwwFued1gEoAcSYUw60VLjRYyjKHdnVos
pWh9x+N7lOxX9novuMoDeDiCfj7f/wP0guJbeoEkAhg5ZwMzrB+Pxm4fO9gN3mweZUbpRexTfbmh
lCwyMRWoEImoe3TkWy0t0pCrjIgZBqURMV1f8VgXddk0bqa29j7epuzwY0ZUY3q/K9z8IBH6gwGB
wnlAhK9JMEx3WxyKlol8g3YEN0KuWVgDIjSDiKmcosLH/lF04QTRE6ZBinLlYuhnIQ2ZUUexhkKD
gDF3+jIjH/+zljQJHC+b/N+ei60tz1G5U00xIfKGYx5c0YMRNeASfDsdI7WcxAmxMEO6CoN9rp3c
VNJYigk3DqrsGnGYzQ5GGXMGn88RLQRbJeXkC6L+bZh90SJEXye+qGl1BTFsxQvQklRnX/GfoJSU
f9LcyfEyYA+c3/bFJSImvjYkza6Cs+xQcpzIMK8gh76/n0Zarn+WPys01pdc1y1ecctBDYstpSqe
nU4+hNA0D9X8Jt3/fYgQomj6vxUfoW3lJkyyT9O3fgWSZoRpOq+skGiDlISW63Y28niVjwqmCf60
x/qPc9Haul4ad6KbUtSX7rKpGqvMPP9RldIr9GbCDR2ZI8O35rgqzHBq3AfTJrY9yfcZRdcwYnxv
jQkSigVw0JnU/Zm2fNOzagebmJ7xog1jNO3woHE2eC/GEJtsAUD3YnsU+hJiNR7HFXW/VxibqLPz
2IqEI93gesKsPiO9zksBjszPiyhJ7VrGjKpbo1sOhDNUnlkNfM/bpaKbn3QweyIimgvU/ALtknib
UKqtIdS0K6uawpF3/YduX91By5lQef1h81yUqRW7YSozDyvlQLp3nsroAW3erSEd1oii8nw6+Rhy
7kBtLWMkSCg32WLuF35B8Axs7+i9njka9lTe5eZMF3FzoUE7Bw480dQEeBYnLmPhJNPZ4w3II8kl
XxWwea3DEUIhhvryeaXNZVSEDw1fvdQ9ZhVA8Wu3wH6b6HUxy/3SsWcnkGlbOXte1j1q7dsP9k2h
n0Zpqnp55zRVnZmouj8MuqixUQKNTlzb6GWoeftfCftFsEgT6WjZ3jBCFYB54fm6aPbHpbw/74/y
onMXZfdt8W04vasYc6kH6CGUKGtkvyO7K3jSVb+aKEI3XK5l3t6GYYIUrIvfdWYp8n8exSM4z6U3
DSF0jDC5Kv9kCTdE3aDzrK6h5s/Sbw3cvfa0yXi6E4I2a7zRRXSwunO79if61un26depJgSrV8D/
FPc95KEkdLdrY1B6WRSVKFmaMaRUUgv5ZzgIJMVrTx1JcN4cttYdCuEzeuPLpOmjwzCswzV9tJfA
JbQREWqJ8xE9E7p6TEeBAyWuebtoe4+QZQayoT/xtaWUVWfrBCpLverSKa9MhywtwEiwL5WvDWzo
ZvzcUfcxLYyrj47ujrrmxjVOQAeu5PUvnlfG+iWw7aSt1dD6+YSMs6ZbIsVYbjDul/6dnmfPZHT2
3JgkC2dcToCtUqvzVZMZaIO4Cgaa7UBrulEK6YfaThUTmC32ZhicgYxPkv/xh9NAvPYsYfruEDQw
HwmQqDgAvNemRJWDLGTOWXPcojL7oCROeIye10GPbPbw0vCrMg2EkqEa4hDrICIumyvqZEDQ47nn
2zm9lrg7tr/c4wlKVc+TE1QW4VWRAf9n0T3zRxJDwR2GUCiMhO5xUIqzKemodgj29FSdCkfgqt3W
Avap6gKf667uFqncw1hKo4SDk45YueW55YJ9PX14cvIn6PlyBSRu3OjaUPUa2X1Tinng8aqGs6fH
PrCgfApLsFOJaODCIfgHxJK31YTWAFj3erho32q8IU+OP5FJqAzK0lbTYz/osYEAJQmlHJWmN3JX
oWZzOmNibyPFDZLdwlZlS0EiA/EPzBZs0RVzCkQqEEgySDhnh/WT6tpSS/IkIbvSi17ArWRzHtkx
OUT+HI787rWMUaUis5aRZakwGIUOGN67ja8f33P/y7smpeQ0zHAluy2a3U4d2xGZoEcgdOKh/eS+
Ia/3SJYCP1a/eQoPnJCo26+WrjZsWe5h4opENUYx1X8BoKlP1tuXRA3194ztegsuGh+H+OAY7/Cb
BA0xRwDhvPuev+G/z8CA62TM1FSEdv0wglMpGm3Gp3eLN0SFczWwgpvbW1nWMiNHb5ZYuBnLlzZW
BPjcPupyCwWgXfovWElH38+C4G/qFilbo+ignKF9v6UL8IzX+0W7P2iLckVtHnjSLoq5p1qNQita
b3GcKB9jNAuggK8ticypCqGz90dM20OXIy+y2hZbemV3Rx7ggfo1U2n419YhXLWc/sppzn1Ohzy3
DAgiiaBbFyH/9+oXVOhVBSEZi/zleZV/y/kWuBt6hKg1T/ZTCjydCzlgfNcoB3Pzkty6oj98u7m0
hrJMDrwXcCh012l2383M1ltISyAFzSjVJXBg+VnwkK+mY8IlHz822Mt8IIzS3ibpcmQpizRLWfRf
KyyB6Li4pxW+TLPA0FLwpKFvMRtDUSYECVhjop04rb6BfH22sb0fjoHI4JgXLDKE/YHdClSx0t3X
Lr8CxeRdm4kktVbL8KkMgNGC3L/V3DYT7rNt6iero+oe74ZfWHSLl1dmry4dg4xfsY3E7kx1aFIJ
Ad1kzglP/Y0h71sTvh8Fh4G65RRAULzi7xVPbQIft3ThZpxIQdwGKusd2kjX3+aCn+AIXT4lw/8S
JaoBewno1IVwV+nC5Zw1n8847U1CKjEuXCfNZvHTi/AS5S65t6MUuv/gVeTIFdTC8mOWl8szXDg2
Ork1Z9MzveC42EmCb2NvMeqbQNT5yJv4CEGNxL/3PmRFLCpgCr7pw7js2f0PX6mcAO+1DFLh+Vbd
OwK+uubFBtuOyP53+fawmaQJc8Wl4nR9mtG6AqrgoD+iai8tmMo/Qe3QIfyJH2avswWejp9jEV+w
PZ9D7jJ4XIHjigSgrTQol84zfB6J+XnllD5Ze9Lg8iWUECMs14pYdVhdXTo6doKdCYMf7HZSN7Yr
gPkTiSZRaxSVc30u3J4P0SQnqcNOeoiB+sTKjYXaex06Ge/4LNODpcL83lnDbKQnZP1lDZhj8B0F
orHsfIiSzN6FF9JCwali6/HkMcyDpmc8CFMzWIJmLgUMe6U0kslhaVBsnApGzlW37pcq0Ra5Sqt/
HX72S4uNPRrMH3dhZThR7pPqjJTdt5IvEt/KRTCWqhbTkLawgw6kFV1mtMD94Pdsibph2hhzY75p
sS7DsfQdH+TXeo3xQPN3m8k7MosQh3iaRBGo2elsalJRnAYBqUU6QuWa4+XVIodtkHWpg3xo4aFb
zpzewJS6+yFrdNqObdhQX/LsUbpZ2OQmHRFQIVNIEoCyua7U+6L9k3TxpWXvrES2gxuFBr03zLHg
44wjG5nj9aBFW1w5wmTIqmrpDk40ScrkPcSHfe9yqyhgqyV4aLqdUQqygD4L6y7BMaLCdoc4Dokb
Lh9QhWoNtaYKQdEdXwd0u+IAKgtOD+7epFiXfKguAxpRs7LBFQao8B83VW866uIiRywAsahTQBB4
IsutGDqgQQPerEi+zW+4BSZ3jJHiXKd1K62EK6/z7eUY9YV2o8TuoI5VeZQdMALzy6SJ2ib1h7N5
0gzDzL7Xw0LRUPCuxbdVaqCyQwE+KyqEPYBq/pkRaoLuIVveE0p99bXMdFB+obSOMcrFGcm3zLCW
TBkC5X7K5Qffs5dlsaTIZFivdAxS/ObOdJQTJQlkwQ4wDjVJgO53kVIk0xN5mrcYFWe4KzLQEx60
U618aMv19/jVJW2i0+pWNimhqU1Tpxud3luvSb69KkzRuQRtW5v/lByeX/NuKDVxks5ij/mxQC0S
CSU98ZNYy9D7F9Hjk3jAMi60ctW1oboqnnmer7PheE02AFHCiFAYpeU4HeZQJvKuaM/oEIzBv9J2
fLzQyCyvtYejNRSsjAqiF1uFkOTGNCw8mUgI7SnHeMurU94PjmHxpjrYV5nsHkVxPaQPuC0heHQE
tGN+1KH06D2cVjOOgBL4d2U1YOkljnlkgLw9PoDWEMo8+19AsAV0UFC21NvDN2o3CIeraZfoaENz
LF0bTNzAWN80Hw2Z8miV3IzaqdOaLS3rjlHMfk7FxoAPu3W9MWQZ20ML7MRXk6XGZ0K39FxMfROt
lvJYzKhocRusb2hxD34PN8f1beG02doMibjiqBGKd5CpP5ULE6HYfRnQxGA0+k76BEKdAXuds3mN
B9IdaBgSbQS2MfyCNqyaC8rVuHlLxlJyKhGo3dEajgaKUXheHRfm6oueFjlg6ylhyCjkaFTf27cr
6MbpJ5zDkyiyJuLPlFG5IFbUGdf0JjIQtrAeahgeUj81Nhk2wGqmWKquLvubBYKDAzK9oaU4oTzs
/gRDNPZHEkcYOxhxXNg0XD/p5yXvFsPMSypSCAzVmthNb1yH+Q5HIoyQz48W3qMu425Iui3EXWXP
Ye8nJ1syaF1Vk5Ag9PJsq5dOwYDCJGuO4or4Dh95PutdU+IMO9JMz8nj0FXImStiw8C5DA5lBstu
XD/trhxVt753C/hYxIvZ5EVoIvLfOv6F8TPcG+6Iy9JPH0V2+1EY7CeJjWAhekB5QHizbEGNF7do
cumPveLweD+8my1+nmq4d/YBojGTfPBJP9DppCO1Q4tRTuMs1c1onbKPr4Lq00mNIHfqzWl04McD
YQYag29CJtM+b+QqyGUYiyGM8cuRR9dEwkrrs336PZeg3vxFUzTAgLeGxM/bS6MKfnS/+Zaw0ApE
2Zg0E3pvmOsh26GhZQx1fxMkNPUWB3dnr/33oODiF8dN7zbC3iwB/k/9sT0osLcINUMDFezSgZzT
jMJ8GTxu8mwB1B/LaeaG1fCRZeydhZ2N1IH1i8IW41Tqj3QlvCSsTI/RKAPp3JgLEc8V3jfUityA
//A8w3hnO6OA8M+2Yvv1sBfWH3q7X0t/vA1SKCCPc1yGihB/wNLfTmoxkVB8NJZQ894G1Lp4zLk+
vWcsxFbCzB28GtI9vPRP3f5Kt+80KtB/YJY0ZReSrYIfaF1UicP7nBiKp7C6QEoFyONUsXM1hOvk
YKrn0icxvdeAYEcsirR95cilDqF1vAmZir9GwPuMCOzxhScE3MBSridYP2GqdD4rT3UXj70+8uUo
ThzrSgTvhdIs0FPABgJxpdoPf2xb3uQgq/8vCEc8zdRqOh6K998l6Y0WmOuf9vZo/pHUwdk7/WV9
gtZRXQXf4slUWzNOi64xjfMd9WYNUbjlkX3mu6PYIxpyhyY8pOkxUT7DSZHZNdr3cNlS3pfGRXBP
rHGX9x91EyNlp3dpLnVckNkeOWgud+YEA2x1uIl4K0LLiLZtVCieeR7LiKQ0olU0MX6JgRNezRjb
FA8bJdRoIV5Mt+Sq9JSqSkQRchIKxZfWK594eOogqOem6eENd8PKu1piaIWSkPJXXccPtH03qE9x
2BhPuhkGy0aWF4gf5ncHDUOisLkHFw7BKa1/MIcs80MtHUgGN9rS6wkQAG+ethN01Ey+LsiF7B0N
GUWfmEEvlbLevNs/7VF4n/O3PP8lZ6NBq1h2pgvnCLaP8yBmuki6REwMg/AbrscSKwxgrJ17A2Je
SZERhyHaIhsC124f8AHpRmXsjJbxujr9MuwhAdRWvSK0jaCazbNUHEWscZAerqnT+Y+0U8xqrqZ5
SXmI/aGrGDCb09PAi1Eu3lSHnU5vBFw8aZJIuMpyfGHdcRa6D39w3Y2QiXdScfJyy8uj2zrqTSRZ
HPT4gRboQtBphFeVAi7yBPLsaCOT6yK8jOOhubab6E/TGxg3tU+BNLMofjgTBzJ9mQ6JqNfxcy8y
wTTaEdhCCgX+MGb4DojG+siaShdzPHH4mHMX39bFiOCJUWOhO3AeBPi+uBperV2vaNApZLBgKtv3
rzuSlHpqewFsWbVLfsDWDENudvYKS1SwUgOdUe0mZSyGmzx7wUx+PPttSOFCwd5AXUSCr5VoxSoA
cqIQfML6uk2BAQ0cZZugqDabiDjQJCz8GyX9xfDQmA180uoWgQ+Cr/ezg24LiSlbLup7jaMfnqxz
u8NW3ggEGLThGbsdMMv56pEBLrde4hQ71Lff4JPmeovouhvesDjtdjgHucGPf/IBsXTx9vqFhXe8
PkK5atbTvEHfMzDabwul5WS7ASWRj4jbVuL8TvdLa6UwS+OJIhFbt+i6kWcATqE95qfyn47tVqui
cy1e5Ir+XrieVR86r5yOKlOedUjDvp+99e8isV5zw+5LDmvvIeOczuCsDgWOVEbcYN94Gnw6Ut1i
rJ3dyjmYzMP+lNW3thVyZ+Oj3SPTtLWkt1X3+JWjSJREfrBtAO87jQW4jzbNZ9bDYYtJC1iWE3Vg
uZJdbQnzmBAeWof7A1sk8fl1kOn2tCd6OZG4sNkIy+xoNKcpLKVuN6spapVadH876JDl/e/sf5s/
6DbuScbmQu+IMN+tcP4/XQlPZfvTRsDaYlV40Ye4W2i/NceLYmUamVo3Od6VoQxqauBIvkfoxRFq
4mWVy1g4po6gWHofW8GU6qRFEMLF0T/47UpLBSEK5Jew3eXh5nZGbmecmDF2GsBItN7Qpmix6Ebq
0YVLkW9M2cC5a3Exo7Mav+R6pWESvjqnu/NiLAlm1VFTHLNdAt/OxZjuiK287k2TNDuo+bDmd1rt
RGSQMQFZMfXKEOvL2LCUKpKUyCBEZ7mttPgBTo4F8q/lqvvEVxk+175nLUmxBcr1m4+1kHlNmI2C
uwoX86W47PqI+UEcK35o2WYYXN3Zc0lXAmnf3FMk2S/yjlixhUaC9ZCasJBLpcAbOWhOgva3BfHF
6BJ4qZTUKXKdONlkUk5NoP//1G45aLI0qexY0INzNgk5EfkOY5/k5Mypg87ZWI4BDRrGa5kX0og2
SjW2ol9xegXPaeo26vL9WGlSFee3mxEyWEbcqQR7heN9PTbbLvNvdIgJ+ebrkg/ESRVqv4CqfdRr
qPFNeT+fRP5/aVLIJ3UqSExV3Du43myOF8i0wSOT9a7EaJFYQh7xirQpIvQaVjwizmJBJ4g8Curl
KOiaZr9lNWpP5hAWVT1pX6PyiOCZCDnYOMB5KQu6iQ+pClS6b/TbZn2k1fkeXfo/vCzuR4olUOGR
d+0gCA+u/XqU+8QTdgFjzo6OqqJNaytQKbapzFOipd3fvp5AloS0qGOsZ0k6mIiCfT07HYgk0u19
ukSpjVxx8sU5buyRzkLp8ICheAclKVGCyLd53ZcIk8n7ds92vHIcTCBeColcxa9h4PD/p+If/5kG
NDxxgPOz5PiVojtggtWoRA+tPx1OOvgckVA7yuqjJ+p7/7septZWmoZg6aM03zu/Z41YmAegpu5m
DrUWgYn0gxN/ZoHlq4GRUlCWZSDiL44go3zJ2K6jsAlqEgJuwgAra4uk35tqYgY1qFHGxEV6c/mM
DGsgtONcMaU9rOK24sAJYVShJs5y5UbaCMWQtSycxCy86Bt8ZHwOU1yMxbwSTKE20UCJIrQqkYDI
durgR0JLYtj85ZixkUnQdxaukMymOBYnHtzbq5eaw/PedTGbOEb9Amxr90rAySno8CM/DGrrYJZu
2IhA3tI/XsL5JkEZacFz+N4hnJUXZdUNQBqRi0c3AnDZKuXKwVnUJaBnz935a5NUpwqRKYxin/uK
3Ad3j2/ioryvU0eso3dzasiSKYSaSKX2lhgSn9SuF/Q12LCC2ptGSWW67Ed1bebnm4W2DeiONCnd
csQogszCm/Z6GOaq/0hgrhQwhAWqJYgpau6xlrom+hofH/1Df1dhVO3SvOFVF5EUR6kFwk6hhmRw
M4lGW0nSvYH6P8AxSgU8EJSN9VDiGMLQSW0iQIk+Hc9yDQlIDs/YFH+iMdpedTop570niGEy2CYR
Mo5fvf7T7nRHUX716RCG29OwNHJXxle9KRIR0QrzeJMw61ZYU+8/TNtwil9D90U5I1PhvOTffkx1
Jh4bCkgxWT3JfroF3N8BUKSvY6V9YHz2SyeZRzmIwkBfO7KViAACZzg6Uy36ZezfxbZRxkPvHbRk
0G8ByBe11RlrFbkb11K/Bv5ulHZbhlOAGyMslabeid/iLtqvBciaDAje13D7Atl2UBNfFIGpI+rt
fcxggX+x/iQy1uO/LcrajWOWaGk0WbR0xtM1VdyT6LBPlYbZkzuz09EsVGrNcbUXJT9C/dyiEDMu
EehSkhgiSBtcuWXU0vjWcnehS/OXCS5JkFGizLZBJODVxngzaUSBfBuZ/7CsM1Sm8q8SxmMNfmrZ
LQWGlR8poTaIhTLZKfKQOjVX66na6D2Cb+efRcAeFOaurYxVdQGOw0dDkiQLBDZNJDGSWHos40zn
my0MWkB8A2thT6cMg/ESfrZmQkVyoyG3EGyZU0YOwBQ8xsu4lAWBFudDi3MANaAchj80aoJ8Esvu
HYsOWjMMHwLA6rT937pFxmbkhmxGp66vW2kx8tJRSqpyvJKnecf+ZwZU1ZmnmhrkOFbzUpNduvKD
hqyecONSjUr6DfstrdhMxNr+QKBooQ6WNdCLDb9AQpl11casSshcfNLQADHDhN1pZk0RoAQnJPrZ
jm3fmuCdlsQ0AFwPTisQEi/lVgB8jkdDzkIyMO0zCV0+6K/2AMFSRvZpxsaEFoOZiohXPo08OtYf
VudaIdT1lVLNjfwxoLxwB7VPA+aTv5Knh06Clo6CkX/TVSJwx3DPQUdYM67CK/4557zHivFab6lH
HBQsgeyNqA63/Iq6EjJLY1bTI9IMGz6sOdlnz4gPaOyWtPvg9Cl1Zhg4ahq7bi2BC7iwj5TbeLQn
ofg0jE2X8M12piBJGJgf1sStoiQkT3CtQzBPK1YR72EKicLUMWMONptIdwuqhPbvm7YffgvD8D5P
T7NrnsifIzddCr/BtWm9CY7zWDQdvfHfMJRa6aypxq2p12Nu4Y82vG0InS3UJUPcgfuLGIbsicXG
+HiFBqaV/Kmloa5GcabA4h+z527tSQ0unZ8uV3ys6mRu2rmqa+c1P4x1z9Fe966dmQv+x85q7yw/
xpKpTF6Hov8/zHqI+FIKRfrleeNwBY/ocNS1yfvMrFAU5tIiUMCM/n9m+gJ3I4AhiJhKLJKaTDz8
p6NQzr785GMc9+lUB8gsIvGuAj5BsPPtpHfL+Fivl6ZfALzIF8sxFYIWSL7GkM0Qb+7F7N5A6Z1n
d/SxjDMPrLI3nDN+nnoPD9T9vNI7RfHujMeY8XdD6Bugrv21BU11oPmgy2Z7O9Rs/IDm0GFBclYc
ZHfMV/vjmj26YleCWL1P8/wgH/KEDzjMot9TukUFQZuDTpyQ0MZ3wpPyWoRigN4nbgb5URMirGhS
5zUM6n4Dcq1Y8dse7anqG8qw0dxxk+8RF5GxXJWBuCNiu6dX0C4HVldbMQMzPSqlCGrofPd83WL2
oPBAdA0qRdBmjMKZKK/jyh3JjFscvRZUG5/T/46biO9ieKeYY2rO+zzfkA76v1/q7lLKTP1etatw
6mTuJ0vKZFz4XbEg/M0NskP2fe5GoiwIP22vu1Y6OxKtIr4tYM2gMkxnap+EB8fFcvb5jBQnvhbZ
SrRV7FCG5Zf4gIJogcP7wMmgua3mS58GsYORxJr1oEWyXyE7syI5A7sfStb70Vut5WdR0fPh5QKD
AuMR0ycGjGPNn1++NRmnhGglQpldfinxaswjsDtt8qTun5ebzQkeOb94Pdr1uIiKMBwq4GyLoGcH
RqbqunbQKk7F8UGHTa51tV42EdpOLFMJ+/TsNOV6pPXFs3ZuJqu3ZOtHd49hYHd5ATVpPdm2fxNL
asYcZJy5qsuan7uW7jWBxXaOQz3hi5t8gJ6hwci+b16lraUsPWx3lW426yszFxxtfItg+/+ljwbi
8RKw7J0hl2y0CnVfPQ+ZDJ4NUedN/w3H2MxImpXZ94aSPQvryEwUNAlUPWFdpBgLIoXuCURszI7i
knBGnqJxY0a8IwDmmA8oNGFnujVQ8Aa1E7EOK304sIeNvTRGpEOzCYCuDQPP80f5H9xRQUTZrw+/
5Slow0YWztXZCTUni0tf7ELj0067uPXhLP4Ty7gaop0qQOYUm0wRrfj4j02/mGaXtk2zoFszEE2m
VbB8suDZMSlxgXmhAj3bkpauwNc1zqQixcHGUHTPO6m4WdzBMTxAxmxK7TnIhO865YSqeoNFveDL
5nm0LvBx943XMAmIaO5RkgXqVOcXy5orA47NCVRWcfXNw1Orhk0jHY3Ytz8EtMd43mne7OuPyKt1
O3Y/zJtAaNPobyoxIdAx0lJQ9neIJqCCg85BeNozHSQNPaeja52HpUuKx4fk494U8fF0P7zOn+WB
24CmeL1xZT+gvkTNn2BFZsSQW1qKvloYD9/labMwus9b8I0hQpyG/0ydx9BpJtN3G4GxOGkVk1+s
R1YvqexeJU1dVNcRs/BiafzxuzFxPElbMn6oxVfMpn8/wgOIffO53+kSziYQapgAoJYe2QEopZtE
BOR/jTqLB7wuzfjRKe/TlEduAeQQj6v2yVWSDQ1KPW9zH+irqMlTXJcRi+7ckxrSK/+G+hF7H/iw
p4xcPWTTFI/n9YnDiZrZrtjC2yUdsHCL/fFLlJSxnIMFSbIU4JSOBVCwfFaQ5jRRqa1efzljnzu0
esZTiuISEYMIAC0yUEtFehBbIweB2zmp3E6PejNoU8q6wYXGB1i7SzRUJwEy0HYNewTUj+nWM987
GX02UreD+Jy7hJh6cnOrSTA0YQLQ92zPojS4ftHBSNkd7CwQF/XaRKOFG5HH48YVxxUgYzWcIgoa
6MCjZdaOOMSJfvruw7066QyyWgpsHStPn21rB4zVKSkxrHf+uh5+x+IXu8b/PX4tHX8ZVeV9d5oM
tDy7Y628y1ReCB1pzerVQXRBEG+Bafi6OJf/dig2BHU8Z88MKjm4ReJk/caCt/VOaT3k1mNaQiGN
P75//vJ7adJRY9FSUTtiJat49yV88735axKxLFf5mYK7/6quIlcyXonXATfCBPrwJ9dhBTI54ChE
QoPM7Mke4tBCbr3VGPGa92JijIlMnrMDfvh41Y6M65Q3pPQjRbuM/YkKck47II+L3Hen2cZEcJQc
pwmB0BMVL/RMcphtuNx1fI+SbFPfOLp84K8KDrupIKeTKaPqBN5bZ5WQF/UOlGCZxBDlYSQVafoO
HYrTX+OvJHGOAS5+pSqm+dIBZyHgaX8/z6ssObNFYFRyS9s2MIzU+i0pHub8BH1aTR+DzzKfss9R
W9AhlexFg/mTm5ZMzZnNeyMkKqG/5Vv3MGmtdibICDWIijq+XVxewXaL1oJJJCooAWLqtyteWw94
jKu7E3gOvIdK5pHSpEw2ahGolI13a0YB2a+VTo+S+mjoK73RDCBdGbnAYQOXO8lK9f5v00ARKXv6
vdUudOChitTKu/Hm4IOY16i2X8VxZBaEJZwkinJZWreaS960oTXquq3/D7ePpB1wIChp7sET2qDf
uOP9AU0ZzgeRXExQFu2v/XNq1WRaRhEWWK4M8z7EteSWMuVwAMbiv4zS2nPD5Eipm45LEUfvx817
5AIiEpjDdjCRVFGn/isLPKspfKK9ZPZMI6a1gc5RMQ4wkBtXAaLQcL5v/s63PYHU4TdgMgDJNcCF
4yRwodWNF36EzYadkcM463wK4E4hFurG1F3p/cCUyA+11V3nL+SPBluxhET7o9UB671TXefmO6uI
hmZn2Oqr/Orp3ksLLo3qq0AxBM78DqMH46S4gx3boVeRYRA4mZoH2yb5Y6/WZzBX1wmIESFPdgAb
Anbaz148QUp1tBHsqY8HmSGGXu8d5IjN2Tbla/spa3vQnVtc6yTEKq9cHL0OLu4BHrWoJI3o8zDT
g9QE+O1DpyjuB6uprbSQGeFzmwIyT7+fsVEslI4IWWW3SfIRDsWk67hrTZB4dnOuC8jokFBTajFS
av7hvM8s5YgxM0aHxgKwGb29qrYwUqvNgX7ah1n7qT8uxxJ5fzjio9JcTU8YrYgRSpCQdZEjzpHm
Og2DwIw+g+2bl8zXfR5n9N6p/97J+iAHyHXn0LWaUD0gI2T61zoodkGr2NzuBAd/OfsHfkoUq3Bk
qn0fYTgphE02hKEUhRCse9ovTz1WBQFjNzbfjT5Z8KK2xC79f13c/hbSPq4AjLPUc8+vILEMWBpE
E/28uzG6mIeIsf9asNEM96pc1ljKjUI6GnmnvcfJsZDAwmwI7xVHGb4+c+jtrg9JVXYAihpM6xvO
kKFlXxTuXPa2B8eDOcqmbsDLj79SFkZPJzguMBFWXjacmLU2qwH6z+F60jnZDMGwC2iCOMNacTK+
c4vhYeOOP8j/GgOf8BNtqCVEaySbnKn7bxv7dV6vCeCsKsSfXeaw3xeOZcTkn/aDWL/dvNRHEAtE
brqaruDlteF2boHkzwPxi8ildNQDQ2r7dWeaPDb5/CaHmMr0fGPdXejaYDNaAhthaLFzbpPBDtCU
KjM8U3gq1ivaIA2kbdw8D1qEJKaMrR4LHhJ6ZmgJjJX+KztzVO5gyllYiC4fkjwDEoVjxehZhYJw
r9D/muHY4WJvbXCegZ6jwdhEMR89vCOSwJ9HU4JAimkE2GErKi5AE54Dqvv7H6wjx/oOtJ/5MR+R
FHYdMi4gPy1V4bx8eZkhRVtUjAhMNZPrGA7xEdHWJmO0P+3e5o4lmxzyYWBawHYiF1eFwxZXJG0w
+gEGFvMg14/v0zns/JSSLs66NuyBZIw+lsCl5pFbtZh1vsXjLwJ8ZbAtgHIu+9npNDAC6JXATiQN
7EfCzwRBY32D1r9+bW9l8yHL7XH+ycNjZhN/lMtyFUVVjXt6LAOCVEh9M45Wyw3lv2j+j0pQGyuM
mkkD3cnk8NdTh1VuNXTuxasKOKqpVOWzbZzYTXln4f1pkyqawGUEeZwLAC8aERbn7BrIjGWTNTro
qBYtrL7BA0wRSx7YuCs3oHIh9rV68wJWyM+Ig9/VSyMqRmenfVGuxCZXjtiNQunjApWZSNefZM5u
QYh8Mi1UsQcUVI2t8ZVVwo+qyIbYvweQBCxPXRTgSWVAAUwuOMRunUkCRfNE2Bp59CaaLL0NE0o3
mcfcXVg/522bKRe4/5zmrs9MKODvED8/mV3OtXJWRN8xgb6Q+CMZNIUfInTfK4u3sWMrIGadJG58
wUh9oT32u7pFQLdGtDSygJWXrO5pOpSRMN06SYGOv5aCUkyomWNHa1zECaz0PDDmHbg09kzfDFp/
lb60Iq0WVXKVi4SSRrbBatv5imWIniWLKHbbd0soFnautp4nDdA0vP9jvZQxJy75QLHunR8hhz2G
8ephk9UWs9hC1ByMZV3kFO9B/1lbQzJf6/kDFve5AshTosSBNceROtPbliKebabd1BgnLN2ewDN0
jyzn7IXVmxF3sdbHzLL8FuNeuL0GAIBOhBWP4nC9ojcU3DjzaU5swMdJpS2n405mB+rAmBXUWDux
0MZ/cWnIErPD7MGyPMzb46r8K4RCV0fZtFxVI+2yJ5w7L87EW8WQZXAXehBsj17gz3pUs1ZsF3Ov
5W+IzizBMmBVPDsiW9qruPyFxs//OKmd+MwQHc6u6ye4n2vGmlnvo6a4LBfu7mn6FNjYIAho1/T4
kFK8r7Rf3fi9ljkapqa2y7CcXeuikcsCfIq1awOMsHp6EcP2jJjZlpRppnZ1r2MEA4CyWpvJQSX/
xY5sMOJrBXVXBPGRvRo8pRU3nVyy3prMZdL14/uF4+DQOB6YJNxuCmGJUajW6Z7ki0jDXMt+eetY
/lT/efWO86je4RnKw8tAxurzmmOtuzulrDk1JKiXvENF081MxqpAKQ6nUXP8i5DMw9SHb8Kv1+zG
sdEFc2puDb+V1Ijg7eDW9xdWUIHWbpsf62Uu+rc/1ZZhmYmOdm6zQeBMougRDf16diX7vvzqoFkQ
nCvorO3+wGvm3AYzb1F88oVzUcnzbHAgpEtECz8hnGwIXsZFcp/9lOymEhBRiOO+AR2f1zhjELTU
TEnG+48RW5qQMODn5b3KMj0DCjC4H5ntCk9ztZ79QeUbVd+qVmbKOwzWlAy2xLv9qIjk7rBItMzM
iH8MHhmQ1rs97Sw71BVoNt8AVhseniznxlj+gOcdAaqe9FbbjjR16Ol++0iJiT27LcdQ8mrw832f
sE0UbtzoNBvbioCZPrpguwnX2GW1CnlDU2RqgsB2pCw+Re4szM4/3Wp6+o4fbEmDrDBUg9xR0UUs
IILneRbzVroXk0Mv86y7DLMcTVXID3XOBZtKtjuooAsRFsbsq3aayJ+JelLqnsHJnAjDErrX8rZ1
nOI4zybolbLTRX7J5vHcI5A6cDviBxpXUq8I04/Q7hH+oM6ZsI/18+HLZkXIJgN65zhNOnvGz+zR
BR263KISHWoyTu9VMSQOT5GVoAlkeartl9MnP8UNzXaQpFu462bUav26jSFfVNaftT2iK6i4bvCy
4PMlWcjAwaPL1y7WT+G4nEL9VrqTkKtZtMfP6M4aVDU78YqtFn/rUJBcCClwbiEAoxk2sQ+In1zO
YHeMGqWYYE2EJBvvdBHabS6Lixe5S0BWAORiDJEnGSICGmXS3Z26YD1yec/n7VRQMYtAUKnr5YoQ
sVMhaTFKUKPRlbtc1ARfHmCsS4BaLM61FHh4T/mPd9DJFFavJNqJwk6v71MBxi7Av6WRRqUl/dmL
frZe8UH6LeeGJRH4pIDZdxs4iBtNriFADMjDXAyOmmqS3L1b8+69qXnlQJYp9qEd5KwPVIvZJt9U
eh/q6eXQC/EKqSYM0woc3BQMPtHytKK0W0u7DNGeYn52yza0zZGt+kQk+P3xLoXndZYMyUN0EZXR
IjLuCmaBrwQk6S0zFJWFP5lRPfVgoEpqarowLxTFISWGHbLr1X2exlwAGIveftWqj7rHFftcIeVy
QCtul8Yc6n3yJhqVJTq3Hpl9rhnfcRDDg3Xyw133sVPjQCNFeB0SV40l2uDT1T/zDR69re2tqbhw
eGIaygF1FnAPXXUW5C88aMCoJhOjsqyG4h5y1cdXOJ83FdhYtGSSFn7LZKAXIzUcRijCfKvLZOq2
QLyw41/T3UVMXJvMMAs+5Chy86GsQscLYND+aPSFjDMmO0o23sO8sxuJUH7URsM2SiUAG66ThtL+
Md/RdYKJ6RiX6gpt+m0JN8lgtYc5NKzeBYl4SE0xlcF5C9uifid+XZ4qfZRwG2S5RVEuwsTTtrMq
wgoZe9gDB+JxHhBjzIPsO1QJl8ZlAVUUuOmnfOxC0u0h4g9/eET6pvni/KBSPPWwmlvQBjKJ6ehn
rzOuW+wAhCXOvIXPF3/e5fuj0Hx1NcbdBNkcVIWaXZwo9kkdeHQy195w11wHLBXmfgW/N6tahusQ
x2H2x5MVgrMiKF/T/BbCYVuj0iwW0EPyFwNsO74auzM357yzaUllSTP4CsKhOqcQzAa2fPy7xoce
ecdrxYE+umFQwlbVgQSgeG9CY+G1gzzi/i0NI139MXiyDqChRz36AuWbx9+xZfMMpbMa79sseDWP
ao2eef3q31FJYG8LtLhiw4Biyme5nni8hCQSU6xJbePPTGLPpqwsWR1tKODgi0W+oAZhLO8tTUk/
irr4XgeGMc3DAY1BFax9vgra1yuH735fVvvhBOfqgrM5Ccwap3FP5jro+l02QXFxvYot85xhDBSl
ca5Zw3wSH6xfiClt5+j7b0w9RtJPSts83kA/UWPjKyPuQvIfUOygnlI/07OkC9rQrRkxxUFnG/QI
43frQ7DtGOWTWigislW8OX8/IujYGip8gatGBPgxy0hX9FnGQIi7PLAcjeCIizSgLjRUXHJ/3hAM
DHxHO8FV4MUaCQad3oz7fwdIXpAwr3InUIdyWwX4LTqgvw2DxSYzDILCnG6DdmhgOjECadTSMEzG
0tVVlsH//edV/hYfIYUT3mKBuaeV5peVlJS6De7jNAg+qQoJnzhLAj9Crnykrf6IloodN23e8uZ0
uXaHP/Dc3MhinXgk5TX1MMub+EvGkPeLIp+3qjH0jc1kMObhpoWa/v2xiqmI8BWCQ+LNnl8lC/JC
D3KZgmFRAAkU38wDvAkWYtoG1XdgM9OWdbUKHyNlK9Dt8MTC3rF0p9ecc5IX1OAXii0KbUNngSLU
F54vX03tR7nyjFoWaUKeOQ9B5s5LqEG99hyx1cy5RUFuTWzKe/uy+PoTiyRPDwubK3V2Ralhgc8L
UjZ4DSkYXJlkFVDZeBzXX1pKlADCYCkwljJq+ASqQzfLInIYGQuV/rEtW94hUnGLs7C3yhQ5TsGl
RhlAESnGPUWxym7AKHxmdRe7wqHQlKs6zPwfiWODF4KT4N3J3ZUGYkLtjlZINjg5tPG+5dfaRre7
/hTXUJ7GHjhS/ddZw+Z0b1pl9kXRDV8Ua90EEyOPNcixBEW2aetU1TIz/YhcSMn/sEsBDKqTyC5u
iUBvfB114xmdVGQcR+Lqhj6Ey1XzKJB0/jSVZlpdEBVGOgM0+uXNAxu3WFAjvweMGV+HP7Io/DxO
8W/vJFAPo7cyQIgt3efHtFpI6a4NJIXruLuaml70WzUUnp/dQd+g2Hi9OHP7BQjBUiqo1jhLKYO1
UYEkkXjYR8OkbBQGSuAUgP6GV5Ttio4LHPPoxNwshkBAXB3RlGmGhyGo7hr88N91blSqJ8xAnJfq
ZyU+xrO64NwhMTGSD443atMfaAR1AlVdSTswUTWYz/g0SgR1qbwrHgYYTGGpDWlZ29MLCSChmqpp
ajRvhCPSybOWk7A2wRLiWhuf7ptuBHr7n3gJcX2MUurxCsWDw76dhzNGsce+Gi4RGZlPlZ+r0acc
yjlZ/wkEvcBf87VcS6wcu1eh9S7maDBBSkt6MBzG9/2mR1o0qRYKGfVSZeSh97VgI0pn6CWex44S
PeHx8r+PZb1g2W9lmYj4xO0rcHpBih5A18A9ln5cyYFC5FLUKYIIIkoC+kWpT9sOp9linuOq+FT/
q4SavnIRfQF/9L05cdLvjfBsq+FzJfSBbWDyEpFfyxH86Spp7RWZ1gW5t6hNn/Gu75wzylaPmQaz
wN9Lq7VKv1XzrqizzlwBFs+fYBgJNVKkqS2maYSLk6hDdesziBHvwnq5SBf8xIuPsHSkqgvJXaJq
mKHVI/jssanWgf1IPeVqQkNbG0nux9JXkTwr8W6mwfTrUdaG1gGjCul05THNTSOo4bUy+hyx2gv5
IWAYNTLJEbx1DrT8pweifxFWTgaUc3kgrftKtFzASyLWuRQ3kuit9vlynsjm5rDqslsmpuaH8iyq
Utcj5AInlhcXPidFuj9HMV7lVBuQF19rs+VZyPWOg7VZ19Wgk+zyGPS8ugKiCVAkFd5uZymniqpg
dSKXZA8Pqa34BCeoyOqEZTwWQ0w/FfUcj2H7+FGX9YWAzq7M0ObVg7OU4+e4ZMUlkZttLJ3tvmLR
JR/RXWJ+q4Gju9tPY53lcEJ2LySNuo8VlhRcWqeAhuyFxfZPw4sFLHbijGK44yNWq2Yt0TpuHeji
SIl8CX3Cu8LKic9OPI5dUoemFJxSukTRzRc2HcxExhkA1N+UWAuMOAXnF1on2VEKwFGr7GgKsiRx
HXh0tAgoSP+rVPwGOz/O8EgwgdQ0P2IOJvxWrgc8SRM4Kt/Eg13D3oqcaD6jyMzyvsaJf4hPk/wm
6vtFUtiPy+nknu3wbYfXNdR7V5rN75l/T5zRB+Zsb4mqT7BFg96Zobrte64kurlCrfPXwEHLJgim
Bu3rGOo+L0tMOc7BxE6I7Mohd9UuXNezwyqEz8j+cqCaDytK21tOtkKUWk5asfJvlH8o/wrHpfzu
B6SeHwkNiz4HseERsEMPTYn1TXlnTE0k+60xXXnB8h4Hb6/eAGcILz0ZCqSQ0Ix5g+SpXbq/nkcT
3vPbeakg51HDDWKklBR4twJFA9Wv7hqDmS9wea3Nf/Qc2zlkM1DVhjZsv8q5XkzRbjaUlHgr2D/p
eFAVzTVXzwKNRB6twQfZGzNQoDYHmGZvhi7rXyCmu2CItxj8Wgfzi8RqW/n2AUJAzgO9YMcRjNLd
Ipq2UxUxhgNf/DvddUo6MlXfKgO+ZIId7tzuArKMBcIcehJ8zJbbhkflmX0e4KVr+SX8u2OAYCtb
hTKtbOZca9iYjud1C0jTCWxa52zVjHQGPczkeIkhYYFBJHBcEPZK8gSrHfVtiLFHy83CgO0T//en
nneo+3f1ZjlOPLYqPmMjWsHNY2wZoKyr0WBYpHMw+lbrJRkjY0AhhXrrdJusRmvinGbNaVncdKhG
9fYN+DAoza9ZeB0VRfmoQC+FBEpcUK/lJG2/OHPQiMAstcwPIxNHqhm/K1F4hLsTHVfakp/uTNxA
suJ33tv2h9APR8aConCVn4zclQVgtlOkiT2dm3+fdzLOq2nDJuwHPgkxOhKJ+F8PwZ/iPab0Iom2
kBvAPs5Grvp3AXFXYs/3aoMtwv2ij5uKhQIW6wMyLtt4aoVeqcOERNkydhK1zh1eMyW9Rr2lQFx/
ZLxJUyLCcpBawx8C0kuac3AcYfbwZakMfrP0wnIXxfcdsR1SNK5b7gH7YSQX0dxlrAI4pKFUXVMU
zKQBIRngzj30YamYLiWmvteKknr9vhOvP6B/jAt6V7rfVNuEaHBkCAbGeyEW95dvknQ986sP+0Rj
8zuolrc7MLATPJvwjc3N7puIiLYyEGvy8YNUOeNCbi+A5Lt8FybdmILAcAjzwy1N+xtzfCDK/8Rd
mRIoam+9rD1rypAt7tu7/4XstdOmfuprxs0ozPUkba/KMPQ4zWouBZZ4iTYRSSAI0RSF5y+nDgQN
MONleIEFsQRFIilq8Yr28qe7A5IjW/sdudD742oe8Qu1KU0urRt/hfljFlV0/ZQ2Qjo1v1KCsPrD
APsLUmTOTObCyWfkMgtatuWnz6eM2CooLwz8KQdsOoCx2gSzSeFO8h/IVKcSk9MHt8f+4i9PA9q6
M55/ubFnwb8F2rvNY8VP2kA8o9LS4aH3DnjklJdCk/RZAVjiHiCYiTlH8F09usWpw6CQS4SDpAnM
aii8YXSVdDDI1dWmglUJZ7uoI0/oEWrF0hHSqOYG96niYaNHtIQynqURdfMd0xlowDmi+juafsq7
TTxRDNUpB851rx6Cv3bgnUD/gL29qJXDJrwaijsIvi7vo8GyHCtS/XVWm90+7WeaOfntb3pSoc4K
Diiho51CGfLI9Gf25LdxUF34uSv4IEhRv6D1+LTiOj53GvcMPZ+f78KDLIcGk/K1SdQEicsBShXM
li2N+VUzU9f1d4lv8ukHns1uOC4utzWCYIFAuDx/T7jEj6j+3nImi901UXOgwg7UPDAsDU5HViDd
B5EZa6plJBqG8vOsqX3e8IV/YO3ZMrNTEMgAjoZf4X2Gh1X0jr6ewZN3HP1ALnscXaZ1RdoeK1O+
WC7WXXG0qAvEuTO9eFME0N+RSjmiwdnn5rJOyKZPkGPAdiUUfSsRaEkkNLkQdTszihCbq2yy3Oet
P2sCHnZOK2vcalkrszQtP54JQRe82dtnSgy1BsLu3VPs8vwCtCDwowE493bTyRxyLbsyEDKan9Tl
V+FLpo5q5WLC9oz4t3Hkf0PM8v6d2bunR2fLm1d70nHdL7so/edmhqyy5ROQJXMsXSPbijkSiXqg
AyUdew9TrQL7lML2xBNMzeW3ujWeUeywnSaQW8iIzhjwdf/n0ZBXE5QXmY3ADumTxkonSsjatvCG
M+9w/OA3d6g8ZutkH5TZ7Pu2IT2hGd67VYsVVz91zHhgDDxKhJ/INZq9xupqY3xn183sEgmGKToJ
rj3fuZ6PgSTipNgvE8p/g+xs33IDE+JWWpYPNzFLojqejEI2rtHEI5LQeqyft7LK1J7qOn3FXdrI
ur2t9Kxf7xJrPCEmnPkT+xI8uwwT9rYbDp7m9zYeTuCm9ExXNl3QKiaq/NEkq8kgHKPOrS9KyeAM
yIJatA59fYtu0CqOIKar7Y2+hT/yofq0LvvD5ntZZ3FhEEJmuUHrHAftjR+OWB48E6f16GCYRtTy
/mofNefa5OhGbmXj+8DvnWluhvGd8RajVxWQD0yX5cjDk3ib2T4MylTucitcs8mURyissknuYtp2
MUdvbaMxQF8aF61RK37D8xQMQ0qX9yB3BZJo5aPKqMnSp+wh/Ghywk0R+/PtNpdJLVCPS5+FXinG
wwXdiz4L8OE2OWiHsC9f1mOeor+UnCPOl2QPh8BxTZfWcp5sxbq8j+njkkYuQiPV2tnJNpnuhcJb
1+fsvxTt6emfcaiW89nq+XXw62JwknCZ4TRbl3crrVxaQkKHVF9xFhnpQQpRvePc5h4+tOjnMuKZ
QKwV9ZAN4Zv0FqMcOVxhVtA5/tOL/M2QIlRd5vj/0EL35wGrKysOWCRK49aAdxSXu1ktKOeEliLF
lg1sizMZqQr5TQpLOmY+7jY7dqtmo59JCB+OhqZdxeJ6BMlzjWJaLPInNDGVThptw02eKA0bOLbp
+72qCbInvTst29BSn+sIWU3wW34ngdyrWB5EA40yI3t14CTLcB5On90Wpc6KQCzyJ3Xo/whE2p/f
mRTc4t8K6sREAalgF9VbfEyEAS3xW+we+SpeVRiExXEegfjkye37nHL9eNma2mtjZ5qL7DGud944
TjMWBOrel3xp2SG9WKWeZV6P1Xa1DzstN7hXb8txykhPcDvHF5s1ObZwXCMsJrHeFCXhgla/TUej
XYvWxgg01yhxv9OO7Mudni4rHtyZtnBxLGt/y7ZWRdBMkes1KXYKu0ThFXB1Nj94+Dlgbs9/QEpW
uRPeGPrB8OPv9HcdBQqP56exiEMuXpScGga4ZBVebO62smUPT33TpvOHvvmerDKuybYT/41WxnSK
iWT2+asfZ6ZubUdxUGqkMrhvv7xJJV8zTy64dFnvv91oljtBcMIL3yiz8IjnLFYojM4ZLN+D/Tuc
PiAvbgtfuJWnPb/9XxivVqlFifiWspIDyOF8GUSm5LzWc8hCoaPWxUjHD74rV0tA7s/JQkPanAie
hxX9EzM8SXHOL6Tqy6Dwv2KCV895TUhw31uyEXQSlPvndd9A/jiDFhRV2GvhcTbtG1YWbwHdcKpr
ImlhyZUJ5i2cp5csRWZAi5A1HGD9kUfijSFq8JKFDipCVJBG1mYp9Qbw6jEyudrHsyfD2ZLOm9d3
FTNF2PzNvYvJfxu7/ORVY6Mqlgy7Emn6wd4/njZAtb1N8uACsiae928yNEUmf/rNo7yHDUlvzz4V
+t9b1ZcBcjDgu/uz/b6bi81dO5of+wtnbbXa19yUvyy1ocH+hst0MnYBdy1BCbriYAwOXDoCzX2b
23kyqPy9yhIfQFeRBerMUqkMqnou1nPjxtDk6FHKtDzlI2MIN3O03IcMrWJQZ4ZxZxEcJIeGhxzx
g6Ec1vXLN4K0V2S65sLmzfacnoyCX+A3yfS0yXgyQWV8CHC+MtWmrj3az2wkDgzTPMT1EMYjVKgl
qrCIfLPJhQLCEVN+UwKxBgc2jtc2m2oK7Ez74qAUqDQXY+TTKxIrFyRZT69+feJzv89avbB3SNuY
PaDD8XKNLhP3IAKlYjxwt/Z+ardKDBotGc1gKUtFBtCxDyZKi3fHAWOcl/PsUjGRQoGFDpws414+
+gaC8VhypHVOtWU6nzIhPJ7xiDdXgGYn0fN5R2u0gzmYg7uaQsx494GePPxMdggy70t62EHdk3r+
A+scOWL9DsPQLCsrYnMggxMNmh+uvX1+RofI6MS6Vmw3bo1kEd3EVCJujGi8EkR3B925f468EuN/
4wyo9ltBz8/Kpjwd+Hx+4PonKEBwgEry36JtziavC47+ZZL7726hp0+AoGGwmedZut3OttpvZVfF
uQdoTANRVdvRy8pV4dpw6bpsUASAtIEULtnNBP13RgaxMMltbTA3/FHSfQ2W/BNmT8OMC1yYvPEa
lKadM51qypMRkNhuzl7C5wH4KUy7hAcsCRipUMrTVp0uZ08bGJLvVfO4ufD6aTWLFeCvx+dLfYKW
ULQrE6eDcKR8E1xcR9R5zL+6sLU6HBIBKvZgIf3r9YPXKIJu8Pqw/rrib50QgnD2GbEHii2Oq+RH
32D1KPoQZSA8gRRukHfpc4LwCzTJYfIhG/3cc+WJpgVXRKi8+rIau8WbUknMRWFwq4cEiK/cSw38
CIcViCCoi2p3pSg9pRvkFqb5qn7M6GgfjFTlv2FDNlr50jq9URrQ2rIzbCiK7vFPPyyUjNPtO4j8
qdPZ9O6M3ZrNy/l4kGgGQfRYO6fMfea+TcY8U+Y4EhAQJEYOwAQ/1yJRqVP++MfWcvtctAnnt6Ys
loatqb3RX5HiD7BPs4ZZ7uCU5y+cEpgIicVsdT5hilPgzWb7QpIHV9FrzzF+QAJN2MxkrdzSRWjV
BdgNBGvj440JzYtlK7DfdKSn+Pq6JDLTeXy8zMBZK0gBH2ljLcCTHx6ZRX/63C6thhRxoVmdmCBu
jeVrmAo0cp+1B2ztIIDpLpZOLu5QzEoykPpTwYWFL5PlGR8mrZ+AKlgKZT2RFdBVPJA34SZxUY+I
cTKs2lbRYWcs52tpL0nVcT0TjIvaN1FVmT4yDjth1+NKUrVUhR90b7dkYC+M/KQsqIO/r9OSH7Q2
GRT7mgQu60EJr/XKqLFV4Qoe074clAFU6qHP3OhLqBEn4F98RFMXmg8SoRWCtO1XBd5qrF1GXP9f
HqcYOPo0BflYxtltga56/E3ceTF/LEr2AcoKnLJ56fOk00zOZbosnrpb13FDAdjtiSdPtspO7StF
53N51ekEH2Er4RCWLe+c+Fjnki2s/uu5noYBQceGsx+0EojtNNFzaenejdYjPaqj+oyzqhXYxAyy
mF0fHF6m7rCcRd0E3y9Lh9pFxtGwrI4WUushnf0Ht06FwKi3Z5zzygz83eWvE25c1qWyLgxKQb+X
N3kpJdOGNxh49j0KTEkLeSA9UJGQX8hXoJFS+alrm65q/E6UxUWTcL3ValG/BidiZj8SKj74yEgb
qkDVAPCr81jd4BjGLXAyB+O3IimekcNwOf9Gh6bI2p91rwWp8PCIzhfPnK5sSSXWg//CVi8tNque
sbm6brsk69JEzKHdHQXd6jBTFZwkVkLNef7ekhSxFpWY2O0XDpT/U72d0IwO+ij802ruPJo8MKJ9
azBzf5Z+/Q15ysAKUyjsQZDYNJH1/PT7eXrWm/EDsdTUq8dQG+MYh08jxx2GTnBA/sYGv9P9aPNO
oZOO6bMcUqHu7ZhQ53CdIPscCy8Syrq4lo6TRCT+a9eQcc+5Aj0EiRXlxrJdMtq4k6lE0JUh1Ckp
q3BbXAh8eMoB2uT+4re1jZ7cNLfJs47acfLFoDVcGGkrJ4/awCk1zymDZJ6zy0Eh8CgKMXqDnQ19
mYFRXzgjkyocXl1IFqHfFyOEPyS8gz1Oy/NzgwLOWqsMJqXaqQMFO+8s8jrGqIWe6F0DrizOexvo
CnJAX/FYVxGTGrX35O/uuWaaxYuFpPf3iFvq8EXOnEE9MnFyDjqSlz8I53TBu8615mw87iqLDqDA
uim05ld3GexzW4N14AUnN9KhRGlk1HpJDMpCHVPgDOuRp/Ol/+m14MGg7pPX0wMk2a4noIhRXxhI
c6Gc0C5CCrJyxVC2n7QcQCeKsAYME7lk820UCI/H4hMW9+zkKkbcNNUyeePFhjF1iDi7B1j21vZ/
sW67pjFrnWJxt1Uca/maMefly2Uxq1loWZN6C1zgawqXxYCKGolYjYHhZsU7U1LXH4TwXjua+6IS
y9s9auoGWpbN5M3LCBBx6LtSL5gDRWhbDRGmhuYuyxY68XihesFG1M6fnrvKayIhJcSz/BLNWW38
BWPBTTcoscLUBb4rKAqi5eqXgWaGSGQxa2F6OfgCTxt2fD5kaR06FKWxpmmpKpbBsWGJO9J4nDfW
96GA+zUTMUZ+6WfRnjHHldm64KojBqhAD5tryUoNK3zDyk/KcTTocUkgBebnxHxw8ZyRSKcWh+y4
KMIyPz4Mmw8INUaIt5mz+XcOWK867CJarPxqHmw67Ht3O3vgqx+nxDudsfkuMKnUnNSU7if0VGME
4bzJyGpKxkJMr8+B+434MNodfD1KXAO0XeHFTVN0aGDtiGk75FOy0CEq4vgBorFApakhhC5udjeP
cOdz+QBCWV0AoexQIJYfYXf7nMTAgYSj1ogSMNw1Y8i/5qlcUlGUnBa3+SXlm/Ow2m1kWZC0YoOT
N0UqQSwuXwNRA3TwvEnzNVpJdo4PZQIHnb1W9VEWp1q23U6RZYm7QjQk052U3SjE6vwKo7FGz8F8
QOLzO5fQRXoR4gclhh+o5Fx2TPUUBjv48BudZxgoQ3th1kdsAEyEeXKdpKMxeKnCuEFdxThezoQ+
Zf2rwV1rQyg3KELRwZeRLavlCpeTrBvV+DbSXicKBRUpIQk/2OCQt85AlFZi7mTRbQh/fwtHu3VT
vl8Yu16dQKraJHSvtAsWxsGr39nw/oWJBHdoDYDSoyXOW54UayFsMB0/jMzf10f+pJIiW6mp3iRx
edJZqOmtw+I/SyCdtOlrcl7Y3jfJBIlHlrPtCsNyVWmfXtOaHZgc/NQNNfr7/lYEGLYsK+aBzR1W
bK86OLOEwvqP6oXcOYuKsjYvu6kRrWHchux5/SyqS4XkVIQC2DoH90LOBsxr3ADHsUyoN63LpGuF
MCYNJ6QmKgZ7p8yDm7h3VjsltV0kCCdE7TdLit74mJ9hd6OgFTMeSxqLBnr3Fhwu6EU7dcI2OujD
gyp6g3xv+ydjZZ+RSbOYZ9Dkus59cJDGWJOkvDzoLnEecvGEMQwZKuwiiCbe8zgdLrg1LZcIXpm5
zQA2Jju0LWh8EJizP/LNikQuiVnbBSx3mYP7/s6ZWZ7CpNkY4Vwj++I51C0bj2w2X0BCnYvgxnGS
vXtOnxWoILbOJrbcHatREVWG351jhEI0g6JoZZb1ig5uWjDrQVKl5+J+Ogc8UnKh8Yrov0CYFCam
dT291vACp7TXxjGN3usoBUAVzta6bFkAWA/iBTxMiCvdq6kBR8JYcHmwz7BZ9EBqK8RFkizQZujq
9ypBCA7fidrF1izEpPRFTPF9W7Yzzc7Vgl6JX3LW/mVFMmoA9iqlC6YGSTXN6+PJ0m7azLF3QqWA
U3ZIzbuXWxRnfA+NAt9sBoq6S9asi38oPkCGFmbk3Xix6wfQ9rbx7vFHapWOcxSr5/idh9b+4QDt
QwRqRScU0b/SxLNdvy3YYVCRlsKWpctajssTZ7JZ/WTLzP1RH4FIqJ7HGBjH0Rk1YgDtfWfBCV4U
diIhq2RPrSzK7vFIu5BkXByhjsc2wEBvhokt0PHIsAHnMQLgnQifSgSmraV9+X8+umfaUpSFHMnZ
dEdj9Fn+jFvJGcjBBXUrjV1Q7G8eGjP3R5XKewCnluaDbhrJwgERX0Vm4ciUnu+veqt9IGYW0QHn
9ADbkD5ypwpRJlnlsHb6beArNkAdvyYlG2a978qbQQ6zhvDzkfrLn+Emi3CNcMk5Mz1uyAcBKWhz
X06zT/jsCDpNGuAop97ca1vfOVBd2CfL3yFlybwHTOXB+v9dicBvV/UMYlqQuWSzSinniuZEb2JC
F0steJ8Ie5Hmx7/TJJp/7wlfGwemFSjctpVvpgNz9txyv5fayee28dy1EI796ro/b6RJfGP9rw7t
lrRbFcqx1IlVNrQcYrTHVaK0T2TQGu9Fy42OR9q7fhwHuHWEaiW3U4zHf2FJqrqjGHm/jUm6f9pd
55Onj8aeRdBj7vyc96RhKZ7arFkjj+SmTXvLd8Nbx9EotiHeWFabjA6tEdfprttvKYcJfLgZHw8f
jhRN4aYvCTTgrZ/cmedT6DoNB/kODSKBg3cr+ADu3BwoZ45nzSllGRfLz1kO2CuGByppHkfHTfkb
mEzKjWYA8yEtm3oicbEtIowuqc754zqJ+lPRRXVx99Bk+t5e34idTPAV3lDp9k5Uvz2l/O9Av5Lq
6BLX2kK9nnDtKMTkke4pcxL0uvGaIi5qRXV3vS8BAny1L24AHTroANt7bqPriZXqbKhaz5PVnbNA
0dk36wX8Zgt9zjoJDIiqWZa3xJm5NaUybcGcLkRSE58hAEsFfVma0nLLtuFIoJeTELLA60trqIvD
eFHHNVdVBInZAI+SvJ1eFJaDTtxTeMlFk7RkZl7hsP3TrSGgY/ffEQk/sXdLJtqNajsn1WVDyb+z
Ihfhe5RfFz20vgwaMAT2g1YpyTb/Wy6PYpduEMNBzHIvoRj7+j/Vz4gU4vpykDN41eNH3p4EhZOy
4lptWllhzWLO0uWHfY1Q4ibcZg+g+YK2jpSUs/mab5TAKSEIx2uZGs805FXQ+NXobalTvZWd3WDp
iwI9zcI+ukSxEhYnJiB1JQThL3PdjpPirnee7jLn/T+i5VsaUESNfClthTI9SMfgesTYMWmTzRDt
HnZREOcjN754uCNHcZ5ZYuYLOMD1gM+TEx0u/4VE/Lv9gw5xDdaRQfbMCELtEmj1ENjf+MKQUin1
p69jVaYATfzY9Df8NO6JAZ6HwqWV47qG7OELDze8hUz3nysNgFqQT1H6JBhym0KuGMDKHJR9pI85
hET6d6ycgZCQAM6pb9jGuXjs3Xj7X0MUMdYEDGpe+/5TktHpFH+3AQqTSiQh/TauoP7lzRXmabhk
Qd+oqfmh4QXpOq0QlPWg9eVqw7yGXBqbqgNp6iwZC/Z1RRZ57qqtxWSmTIONFjItSIYHI82gWYMz
6kfoqfziNbAN7OYvSuOe93xAJNi67nbMeXUEKhw5199tNcv+pqGNJ+YIXxn+tuTOpsUSdlrA5jH8
WiqDXxg5dWweVDvWvZbS1gudMjfSLKPTq5xc8KPMjY6F6Vv8I7Ve3FL+d/a1QnImtkJ3hd9JsY2D
SQPFftPCBVqUI5FAh/1m9fT+OzWiMN+F+q4+ymNcdjdqyMzs/O+20Pb0M001y9NwKN+u/28n+FRe
+oEOSVvWyTIAdCJFntRn7yaxeQ10vVJhLcajgeGO6If1S/amly1YkZO/iPnWMpoqFJbeLYBv8OD4
YkNAfbPzKwECJZt3UiOYrnHaSXT1ShlabZ5LO351JfBqXD97A0mB63U9dzfXPB9ZWGtSQ+HW6G9d
jecP0oBgucCozDl7Us0Hc2W/ICDPcm5F/XPQc9kVQOinbRfbTvh0BlDJRDfCbo3sa5FqgBH3ituq
NQEyn45zdt3A+ArERo+wT6x/B+06qpo4ohAGFoP79QIMhX98uq9OKcwD8OEbwieQVw0fYslKt7dM
QJKNTxe4sYcR4D66wiqC0hv9NopK+Wjl55uNImIULuCBs38vmTCzUt19i6h4Lp1Uw3Xnc6VvN0im
UiPtA75W22109udh2LhceZZXec4uK0Y7EktgrwjCWztM8LxrbZWXN5u5Nukpo8hdgLxQhi91rEN1
6StnxlElU8DxkO5TtJqLJUCzvioq0DiHGbI86KAwQOnFC9B61gh4E5jQf75H+xMfvbd4Rz1EXHH2
mcPAR0/6uadZJe/fOiAqfQa4bWMZhYeyktNRY6bIYOPX3ktWelXSs8m+pxe92SFEAiEoZeZr9BJl
JtX15omh1nX9hn2N6RZHf/ClG16TCxUSibYVMqeRUR7/Q+TZpOiC3wWntP8luwk5w+pFIZMz55tr
YQEm0GFxocX4VLG5e/r8Hd4kQvKSlAjbiS6rq+MF5XkkQskM1C0jEBa2mZ05OByCvo5a8we/mcUD
GABqVsWAJZnKZ9jB8ac0WiwSdzKsdrOpykMQLL9uz3Bp6xR/81Iao4N440KV17hAnwdRLuNqaTXX
2uW2usKiU2AedznhvMCYh8UbwtVVKrefSigqDlHfR6Ot8hm5rxV+0TWbJ/T1VCbS4OJn497R/RPs
cdm9ErmDJwwVavGQWPjvZ9RhUJn/liT8VyS1orHVdZFXrHSRajnPF76wGhLQXjmlfx2q7+9LWQ/n
pjF2F2FcdU2T+yNpQortqAOeW+LrSCw25xtbAzKCBrFYaTVDXuS2i4eh64j34DtN5j4EKStwy0Fy
r3+K9BRLrnw2C/yf7YX3zk1exF1e2MF+xfUSptpaGFQMvBr0pOQX5srZHXvXzQ4w4NdrZ16bXGzd
pQXJxDydrUspuX4PaS4UWaaGfiim2//0oW3fLi/bHrR7W07NRNUeen/nxXsZ7DGPCObTnVTppqTW
QJPOG7Un+OAPJ3TmR8I6YtMV1IMy+MEBDJLl7x01bK+EQ79X2bzDiX8IJ9NCQSIvOdneRZ5AOI5z
YHYSFodSAopVrd2zEHklkntQNaka3Er8sorye9fByRoRtykk+C29gt0LC0FFXvQnTar/IgWZd4EZ
Dw8QqLGTpS4PsgGAouJ4JdAdKAsqFuSwPW8+LI9znDcwEMWC+HgnlhOSKIyvyAsp5ZaDyrfTrFhM
3c8OPglzA0j7+qoJRGzGXcyTZUduFhTetzggLFpOaszY0G83KOAN7VGJuSl2gDAqDpahiffYMqZu
g6XCYtiTQu0hNHI94JnIP6StBXuHYgIK0QIUPKTXUgQw9xiOPzsjBlwOJCXriSZiKZ8xv0DmWpGu
Oa2SmLRdnlAdYyrFgpiUXzjK8l06PEoz72TeZtdwg58UFOvceVR5DsL1+rgbJwN7719MMSvmIxCF
UrBiyL/fdGfUeBgnJzJKmdFBxH6dYWveNB74IPlNiwQ/h8luQbsr1YuwgyxVLLx3Fd7CVd+V2N/H
9NxAK4qES7dXRPyFxFFOJDfBDyh/IFymWysZ9fz30agIBRhRgVHSSyLb4czOc+yqx6qO4ol5RgjS
aOxY/Q679K3vGQxtlc2FdRxx3eBlbodgmkY8DFAbN0jTcsTQmXexqcOUHDEqAHCFr7cwKlpnDI/0
XoHFqkG/DBXE3waApcDKenMKmi6NuI88+6FZROFmzahNrZRAGshuvYOpXONvSTp/UMHmgXatDrHg
ptcW7BNfm7IPySqAgBwIKYcX4xL2XP5ArxnpmEvIjCprEC4ww29UqFKv/qt5dqVjGhQQLe9Sw4+9
8pV5p+1GhUf4I0mBywtkmfNEZQ+tkjdR0qPIkB2pU7Bi52wvaCHJw0kSo5WLgm3SH1ATPqYEgmyC
pAwCJN41rxqnp6PiV0hpQ3YJdrZHXhT6T5FeYJiqFwEx1IQnFf/nr71HYFl6D3B3bORunRHNK9Qh
L9Wd0MxmFd5LBPGxmsk73+5FHR4zn0/CiK0i2Wtsf6h14xTR19lUFWDvZJbSz+hQPBwuzEFy9zpV
Ztv3fEXtv3dd14xYM+KWn0SNxUMGGq1B+D0TOGms+VPGHLgIv6WUEDk3zOlYuTVO9eFy+TTQbgYV
wxbL0jvxTRYEQM+6dTvvBKnTJQwhN8jZXZV9bawGxGb7HdpZMsJF+uopIZJPP81Ik7CBvZiKxspR
hFdle9pdS3+Usi2NHN86neoCOdsI/Tt3EOwkN0oj/f29hxVGZqWkmhTsHQU18mHvTANE90f33u5i
o51ayAtbDNGaUXd8vCLy7WR1Cfs5AONxU0D0e1+jbDfIOAab7deK0yZXqgWZmsO58soYvSa4oaiZ
gp55JvMau8zhFgG781pWnMaJkSPT8eRp1MOmK93MoC6wOP3JemV8PK8Z5PDYeYtytTUcYGXYmHIo
uwPIXS5hs0FUrr6uNp97dhPVFKoMayvh/MQGgxQdtWK3EwRfbd5s0azOTjLHcEIc2oXj8qhHLq/w
n7ERLHz9JcUbPhO2EL+cZ4IfubPcgDcMn07xja4vUjlDcj+aXl+XqVh/6AUOlkNfmoLyafAJDhkD
cU6OKd9s6McS8cA11/zdgtlvot1U6hrZA9l8u7dqsR/yJNVmDD400MbM5sBa7/4vDlu4mbx4umFQ
q3eaxKXfFDZytYIIG8w0kmMM/SsZhwgsXw8DpdUMtZd8pRNPmZJ5+EUHvc5WOds3lkWgPgMxRz3T
O6Dqt6sK/UdH0XR9EjzIAWOjp1bWw6l1vkLOxG7JthPm3qoEJwyKjaT6eB4Sx9mWPJB8Ac8+rjTz
Khj0n7R41S4/0JvMcr15rox4PwIRli46OLfS4W1LGovbJB1RoPMNx/SjR1Puzwccd5NnFEXRWHMu
t4E+XhY/ASYbRt+G7B4pwFSz1Q+PlKAfOhtB1n+8meLv5/+HPZbJs88/V3b3dGm21NJRgpD83qa3
o5by7xzwKCOlZ1HD0dm0ksTO+8ZAIhfnwtwsJh4XXXGP9pTc6z4ukXV+Dbnv8UxFM2Rlb5F1E5z4
YGlmIbSsjsXuFeVwb2kPKwxAfw7lbS4k2giDk1xOQ4sy9aApBf/8rrtnmixBCX/UN4z9JYCA5GSQ
0BIuKFLPxdC5BIqCU6tT96JRNTkRm8MDi4n6da66pAEma4kA96zXO+/Ikh4wxvtR+kkn02CE4NLI
tKzWfnxwphvq8yvKXbIeK/BPp4AV7aZnjkSNruGk59qgrDyTBhL5IrgVj33bGrOlljO94+wyAHq9
AuLuJZ6nJHXuN5BSE7eD0MlHIhg6O6PjpwIRWPu1KbLD8F53Inv0f5n3GdGI/PUziplsUMIv7OIs
3b/YNWBobjg8XZ8iTTCdNGFwFvR2nIixpmBmlpMCdHQMO/3QDFuYpv7CW9MukJsOifBkbriOdY+t
vjsg50S7NpagdXJjtSatrzIeeUDrfV9lBvGnby8jZXxVds6EBwoKPquZvJ4FkeaR9w05DgkwMYOc
wbZL2PfvZpLpkH4NICwyTq+51gsCHJYXGMxqFpGGEZRgp6+rJGl91SZSVBIqv14X+DKmwcJf2Lk9
E2SLvVsXl9CO9IB3pUIAL+Wx5/FJY8IvCXGO9mrpCyvz4d2K3jZgGFr6M8HFuKktGfhfXldiTVMa
MVO4+8tF81GMBh51RKG5qz2jtuRdOBtKs5W/IeyK2GZZKocqcofdr9SNDBKaL3JnDOsol3h8aiks
n/R94MuuXIaJd6zgrjrVqLGdv/HIfjp3LIALnDThbHEkuDzAqlbiGdBYnte1TGDUIYyrxrD+1z+m
xLJ8BCXVbGY674gCCRFy1Z2NiU/q/xzDseOJQ+fA7cMpo96aFM3cP6j4wMXgtAgT6/GHNwnXcCmB
so30E2HpU6gSDfx7JEsd5Zq+YJcoFNuW0ls8VuUME9v6UqbjsXbPEhwb82PnRHfZLJUia5bMF7Lo
uiC/7q+mq3KlugfkApb5mxYlK2tEbR0p/XLKK4d4rvogKZ0BLyNr/OK8lw7YmPIh/cgRLg/lk31U
XCOmTgfbUhhHfjByjE/+NwiF6NXtzEKywRdttNgL44TgczEuvpUZvbfnWBpbUKN30PyPJTtBghIC
zMYd844HBBvGD8zhAy5Wz9WejNySbyIdTXtIpLozMZSCXWOQlCJMGqVYUWFn5EaBUj4m7/7lhrSY
fah+fwfV05Mz9ZCunca3uaUH/T/RXdEs9+fq8WsqyjXVyqfT3+AyDESlB2Y9VwU0ySPAWT/iWHkW
GHOjkC9OmjLEKxesnrklGlwWRSOr2PRCyn3kKEw+Vne+iM6VrX0T75xeZko5RsSvxJKVfHccQVxf
ReCYPFz1meSXfle3/LCcpGPugQA8mdECG7tRaD1vNXzdTVaSNcQJMuk7dSHwycbW1Y/ZxaOqNz/W
x/O+njTQxhGHJoQsXARWYzDt5s2SDHRKCYBm1iHkyAexOX2THxrvJN0Co7ePDfq141xS/uc6YoFg
64oSd/OkDeXLjARHxzZeEV8a80siOVg53rg1BlJ5t8mYIHtTZzGczm7EcYL+qXeJyYFKu9fTeP5I
7udHB8uqqMsY+rOqLO5uu5Jvb+2vcj5y2glYKXAQGDVZs0w4f30Y33NjeI3bAZohQgbgnDVXX+3d
Cj1i9VJTM4jr4Y2iNWky7lJ752hZyIT6FJcK6IHiMCpfum9mG/ZKYop6zHEekoSZMeIocokGquyk
/Ob5MaHm1juxU4cEtZG9bLbtofEUtbHUcoenAaFs+8AQEZenMM4C6qma5bhgv2SqrhcY2YlFKCCE
dRm11wVM55g4Nr3/yYtzrJEGJ0woZdiw1ukEfo+o6/1xhGMAuXNxW7U+Y0nrvK4F26STRPzaR8cy
nQ80VG1sLZ6ZqMoRExJoG2DmJgVfHEQKk05331iF2GG4wGtuNJQbOqEHCisYtlwjljDLr0RVs+SX
z23zreHl1tVXgYpDcmJNAUhGLupU40KysXSMUXjTCmT2od2+ACy0dKjS8mBF0PKZoMUamhhOpxGr
3h/GBkPbUARdMY41+xxxgacuV5ZtGwRIQFA1QI7TSSetekjANAw2OuYwzqlBhiHJwdFQmNg+Jr4S
Wa5ScekMdmJWM/HSXeqN+auu7hJd0Srh4aCLfzhBAnvFzoNsWqt999Eev5lhEAqKlDlU17vhIZnC
WGYZxJwizE5oN+Cpc4Z8TjenZoOl63cx2+xhxICdNcWbT0a9X6lj5zZiQo5lD3HVyuXe1Ax05aBl
2d9G0a3PcnO6K+4jo3zyRV6Y3vpe2liCYIeHhU7ZxnS17orx9a0NXUdArSm3ZGMHt1WKcztcj6ZD
PaJfStXu3YG6GsQEJzwqGwo2cx9Idsn7qz2q4ozdkloBJoO8Q+mXJn8vFoRBjTftPbIRtDq5D2VN
HfJRLRM8yzIzDtO8LP0V57UpN/tzBU/LMvLHRjEdXf56MDq7sjmC2h8STMVoKHl7xMAw/UK+JbiW
xpVnTLlvFHJHi9/90xe+dTxrU1N3lheMkF0JcG56hHTCKCoRoPK/IDuAa9CCJIbeP2bzAUAQMAG1
OgEKNgrzbAvSqWbk4Kek3Q7gCOQb2bf2zn7pQrPEnwr3b7gewvfpi+dtyOOwfV+m4j5+nqNGXOL6
BnpAZNl73c6gL7hpXxQtifB8x/oOyRAFVlli7u76YXZ4NggB7oPrroNckip4POvJQYXvlzX8JvmT
oW+SWtL5HMqpVrKzuUHLgwzdUPvD9dY3c9139xFP6xDSBa1y5lj+cs4Zafgno8TbmD3j7T4VdAdV
DenVXshBHiM7WXhxByAd3NAQB+kg+gtIyaJNX/e0YyX42iU3LwKBdJjpmislVTdnribQHUZ3lvFG
U9PAaRdZxJGVUGQJGTNRRmQCBGq5nfEJ38o4qDIaB87pGvtnzM4RbnAKKuC1tq9JX/u7eV94vGs7
X55ZTNTYVnuHGak+jW0zXoUdrYziB6aRhv2xgR5tjhz4tMp5kuDFFvayoCOqNWDmFHruD1Clh38e
vjmmHYdg66pNMGsZlc9T1Nr+dAuhNhI1cI/fWbI7eZCNIB7tYn4pkMeClMNXkJ+gL4lgC/gwFeOr
Zd6opTR1ZuBu/rs84//nnJ5fgay5Aj9nFDhHgiEB85HNV4gOnyHDjPTGwCR+bTx6/94+uEQBDS1V
2ZbBDthXC7fxfKNcLa0JR3EiUruU6YnsyTbt80N4zVWeaasjzlJbdtE/pFZ9Q86YmDYD3YKlsIfX
GNFqPXVjVo9WYnaK5iunxYyq87qqW9iX0QtTi7kk2xfee88Nc5748XRJtx8E/9Wa3Ap+6jgLbevu
XDlTEDd60bZXt7CNKAi7ACgTWD6L6yAdOiyDs+AeX+6NYJUlSKAWxk/tWxMaalR1MgvdWSdg88QO
jRBEe4NR3Y0K3KyuBcJEgahqPWawDs8byByZMuv/K6KD53ikR8ad1bT7bHQgW46KfnC1a3aR6ukl
XPcfIux43Xzr9gzQ3NzRXv9dWIOfKTIEo31vYCkJKzjMqUfqSjqRV9ioyJHvu/eVLQQIgOKW7egf
pRKHWXXHWD2Sb78uiT1B9QvZIXb6ZjyxCxpHeW7FV3iP/s9oRQ5vjq0fdXYXMaoseLVWnsBF5Jzw
pC+Ra3YEFb2lobsrLVOENuu9eQnF8YmjibNFnJTdMxF5hX6pOxv34Psj/wpo9/EWQ7bfFf3NOgJ5
0y7BCG3eR3U+KA0GvqYLmKLw0s9aKR35VrF8ixcijQ4YB/vqZLK1FU5rXPhKLRlpqFGPynFwIh8j
08mI1fRgYohcqubLwdL4SY7q/Xh4eypZAtaHL6jcCkwUQek9LKzA7u3vdIjSiGEMZiWiOwRv5pfw
7S95b3Xa+CpPjsgJGLbWCtDCXUm8a1WBKSZbJ4hH+Hhq4h1As0WiONU7YFog+lQEPIQZwaAcB1oY
BYD9PTTNGRERXJDUb76wz82rIP1obEWAib/1EwFZduvF5+cZiG/cRaTuba7pm0oWvO5RHDWidNSM
//jWR99y2FwTyeGFKNGVyjv1GgNN4Crwb9ELW+PFdwiJ3evqn32i9+sgXakt6+nt22kxtlywLvO9
2dNkKeGbkk5uiFliOn6BSX/avMEjawCkcq790eFTjR3OmFieWq5MkxLypgB0HXE8MzzSvbzYjYzY
M9nig8QkEVdSPF79KFNRUjYeVn8NiCfsy3NEbO9WqKPN7YknGhts2rMVe7LtMTziHqojL5Z5H4XJ
SvLg90a2itOgOp1aVAFlElDk5azEF79KB1xiLeltXXPbrlSs+Lc2Xv9ZtbOGgJSpi1e6OQ7ij2Ze
N8od2deXIDRqEt8lYzIHdyttqK0mqR660azOx9UoVddVJFKLSFQy/4aUtAAhH70OBP3Qvj0NUh9r
jOuGw0rpXfu1nmjblEGgRrQm9z9h8i81iNIKX7OdGVhW1k+2wfmGwHsBynbDNte00dmB29enAq5q
N3P3h01WHAqAhYH85x68RcI6Ql6YcmMzuKHupAZz6BwsTiYTnHO502SuK7DPu4ZCZ9++GcOEaK9H
7DNnDGOcWZ9KjO4MM/CpRnx+lbGc375iA8iJ3VMtcfsM6QkmAu/WeTlLh+nPNLtLMKYIWiIGl2aB
p101+ii5D8XfCvzbVPAeeay4gvPNoa4jX5/qQ9XGuRRw3S6PLAG53IV9UlDYTX9qlOyFWdNSbS9G
/cqvtMFjPQeVntaqTgJr5k7kepJLXM1jVrxf2Tm6sbihy7WJ5MZlQB4mMShgGRfudYBFzOgTo1pM
zok6EvObjPUBwa3QlRVpveHExdNQAFcb6hrOqHt2oy19SuVr+C4Q97S4E3QS2RGmzeP4hPoEvQ9w
I3RM3fi09gBfz6pWPTOxU5XWYKmQg8APfcu0KTli6bTLwI6PoJz/1q0dljhtwHnKY40Htu9wJ5yQ
BpfCj5zvbQew1Kd6Fns7gpQN5ME83PuAk6FbU0zG3xPdBqkiGK/XRIKS8FRPNqp04PHNGMPPWydG
AJuFzoAJL9fRfQvdz9s7eedKiB/ATEFmFGDXpNZsubQjzLTv7i22i/TrxZpjmWDxPv/VvjvpWsjJ
Lesiz2YdrWerah+wPVK+JEjQja5zi8pjw+K634B6qqvDReaIyfWzRu/vcHtyXK5ndvc59a18FQ2c
MsJ7iA2ocLhPeTd9tG9ZPGqNyBWjFLDVFPyBcmmjUGKMPQA6Yfle2/8vemgVq9p4IH0v12Rg1Dt0
bQ1VV3goC8zNTNUVClnfujDyhd6Mb5DroSPnYMIVr0c1gbr+QHaAzLh6+zKH9MAl2kJz6j/yi4Dr
TrGI3FzARUCWBtd7CtndS3mKXkvixISN/YeFYeiGrjFGfm4P+XVKZ5k21dHFTkN3sAAe/ihvhwtf
Bv3+9eJdjgGJwHFod0ePS4Sq0fT0C+WhDgO6ZVU0AqN3MHjNG2lL9mhLMBKTdeSqZez2EIiLOb/Z
F5zTBGTfra2FFB+YCqbvnBPMEWrCW5jruJaYdBJTkrtqbMb7ttH9ARyF2Y8kczqS0oy4FZ2ZKRHz
D06vXyHIgP8Qvvez55eBxiqaaAc9muq9RDtU5jaAXo+Yx+A3UH2W9ion1vzFs6pq+ieiFILzgyRD
ExaCVwLXpiBJqeBmrbKHjz24Jvwnv501ENFVmPpEiIzxMcw4ZJ9kIWQAdw0EZfR7P4rjEh1+ecNo
BSbIYFLtUJ//yGvXlmhw4vsM27bBQ2H8+Q5Ck1tt/sK1xuR+dIb9vkpov0S7MLDplezepVaF+epn
g2VKD+EYJy/GYEKgms3nl1TfhUZeum7m94cCgNzvNljoo9aGTIF6VhoU04gtoWXLBomWETtzqctw
fz6/fzDKt/g9ZqAkT8b1/PkMUcSavALgbZe1/pzQ1ecspfjmLB8JpHid+zKEf9V5bKSmZ1TxMMMJ
gt1+YmOmOVzaX+LPOdET3J9KmXI77YVU+Vi19A1ev1dA+gZUrr6D5DUhitVlBf260DpU6Cxf0PQR
thSsZT/N3ug5A/+0m4LRG3n1IdMvk8So2NDLCE8XKuL+EeEoPFn4OQclc0lD57tqQ8t6ZA2iCRGO
lQrpnSEOtOV/w9KO6GanYdBs0fLHiIR6qYUD+VgIkw+nkHVilmk9J9V+2VMvgd1vL0TZJS3jJvN8
hURB4gyCD8Vhkybdzcdl/dvJ1O4RzyQsn7yKHLXbSN8JCUFa06s2Dx1xyIuCoS9KwJ5uy0yJ2wJT
6qcZFwGMjb3auaveJwxiRJe1xMiHMrQqOh0dvcH/uI5vE0zziD58GdS4stInWLRk6wxw4neaK31E
XIYsdZO3l4d9RPjAdMPY5b6MIVp7P6JrVf7TMgCpwL+1h3o+I8fg/TukVUW/HyJWMuWaGoRxbg/p
qfucqcandBtgmVDWYzfnZLAsTyz4mKrh0HUJxY3nhCENh2Jj6gkbfvZIQAIStbd71XOEm+hNZk5D
zQYVj9nGCRCyfXA6Zu9ID8AphwT7MPwZU1NkIFGWsjhHEcr4SvhofAHtkVghCtB28GYaOaOx9jSW
VL5J3w7Kl7RNFE4uI3yj0VDK3eAmP6oP/m6scwh2EJ9oomjl7Uo6s0Bbq1S5Q789nIW2woiIjtU/
0vurlwFzujhvHnN3dilSM8JcMxPWvJRMZvV+DZ0rHCmd47DweGTT0oSJAN6fbSBiyjx20b1pD/ia
E0HTHEfHilIvMSj8cbsohAzoEsY7fBKBVUiHcFzLk5NGVvT5CSL6SZKGVmUFVG7uU7vZfMu0Jhkx
AYvbgey7KAEMYifbNNNVjPW2Sc+Fl51lHGJvk5k7u5LP2cNfGZJ/+n9AZo3ht7EDS0U6D0lFcYWn
UISKHYxRebPFLHRHysOpOhaZDmbP5hmFEFudRsJ+XC4qWXCvtdGsnZL2jm2l4uL7VhhdPkgQncWX
z+ZMTg6COFhbsg9RP9DgbHwr51VCnmmYF8AvBjub1RdaKDZaYDDRdAaKSb79sZiyIQnyLGQdvxex
4SRVkYUcElcKXohjsfdVonUZRMZ6HlgZ6gIFe46yWvvyHc5NRAow/+igGhUKVVEBy7JvB5gc1LRp
5m0q07GQXtkVkJLg6Fx0KLEQphnbG1wlH0N0ZkYPqNSRlw4lXhTHFEDDLK++EcSRLe7OrZlpsyUF
QwV8XMsGMXkq06CFt6NwA8NNnG0zwmZBugI8gxZr9mXMA7mD7SYFFcug8cy9GNH3PmCfHxtiXUUX
uSP/N7TsMDZzu9Ijr0mQ+NhBL4SS6tAbkGq/xmkNu32tKVHByN19ZpGM4H1O96cC/hJmrMbEgrEh
gXWR52UfpeY7d75wWf2oydri+gWpM744+eK5OlpWaoCtoNmP34Ly2W3tag5tdmKGKR6BPY9e6TaF
IE4EH88+hQ8mUaqKXlgw/AWAOb2Bgm/xVjRXYqYzzgJa3N7K5usHsl5jpudVCMI4rLhiH3faKT0q
F9CzIo0WdTBaNQOHqSSran6AnXwAbUFv/9bA9WuXihnvpcvG8E8zwLHkdcvy7WXitW53d4cyWzOA
G3xV4BHVFdMbe2w54ZVN0+xTSEtMsc+Zblg9Py0E0oALEbS/uf0p3vd4dlTb6GSzo/ZFG2L1y2sZ
qEbuOOPy6lzSf4fYKvsyhfSg5y2q1bugGXG0ykRsoX0u7kB4agLsi3+xUydMNTmOZLPz/IP0VtOo
MdUWtUMSNYvcT8FfkztSmjmMMuFhM/NAuP9HnH4pGVT8vjuug5P7akqWS7zTkz8SXdpbzUTe6Hxl
wCoiQcsMab8NknU3Bs5qb9bj0RrWXp8b62n5LZblcovyNxTnbzLANYXrfsgf6OyPGsved3zHEmRu
0XSaCUHDn5BN7YbM/VToy/q26dtkEakcyM+4gY58QNkzNzF5rG+Q4HE8vG3Tuguvsf/hSm/EW5DA
aQ4QB+IFkKVKDibw7pEGesWrnDBfIpx8w0mBYOQRKhzVZUeQFgANj/T097SdfjsebM2Z9ZBUy1AC
/o0lANFRJDzaSornebRQlCp92DMvxAoNiEdmNnLeJeOWbq23FdsUPGx3Jst9wRC+yTLlhhqp9HfV
wTMKDWfUJafCUrZIBYrlc7jc+Xd0aLVumNjRKscoEoEGzkwcSSGhwOxFTtZ1xz+tB8CiZRsURxGF
YqrhK1KHtojufNgoWBel9mXQGC/BpIW+y2TI/O7NRWw4Y8gJ1stChFdwojbulQ3V8PRmr9/46nxM
bmFP+lawBu5/6Onfel5OfDDw5UYTk4tzEPp9lcK6RbcIrq3CwrDKrarLPq4VUKtzs8HYZdkFjlH5
/D628oHvUng8udGPQ0fEzTmafpbgKBKmLvHB7q+8NsvCbQ3qw557XaOBUBvrKfRbHOPR/y5Xcnjs
yWvHtxnyPD0zgXF6GxiX0TBknZ2riI4/E0dpPlbD4XBVuZcynSSwrkzjwSzvDCgGfUOFObrjM7F3
9pzrr1uTUPGa9Fz8440L5ynpkP87u+Jhlt4ExZNZy51w+YFb09um0XKddUCaSsk2niKOby8uLygX
Y21/ZVajdatDBwN1a9kR902kUhRaN/6sn/LN/CzZhc47IFNc6eUoKAcUbboMKBoHrgUVP3IBe0aj
lAGSQTWjNxkE9Djz4LSBN4f16dKsddOvN6E6Y6qjmJ5Br6bmNOOY/H+8lp0h1rE9A/XBDkMkC0mO
+KDbaHlHzdzpMghR6Tir0pUIphSXhLhn2Atsa7bcln199PbNrd1xxSNsd78d4HnSDlFegQWk3FCl
zsP8i6v60xPv/QmMtPgsvSvahoT9U2ONy8B5Am3+JiMNDzcQ1FqbucnTWQC/nOSElOhj6yAC8hGV
hmFr787VGTrzbkKM88raAC5wgkDT/SwoPFT0AsYpwP3/BmIKNmAjoiVzinELXlgs2utz/3gNVV/r
k1X6lt27TAEyZC7yrnrJHyG0SI1QvQQ0935w9Hkx0oPGzLRJHbveEFG+5dTTxR80IaN9r088jR3C
wXe8P/Qgo/k68FYjfwI5N2jfGj/kYnBuqIf5Q+U52RYH+c+WzpK1pALPG9gTqPiwGRZ2YvpP2zKW
aXF1J31EtrDVnSQPuHlH9hbqV/0pWFtoasWjMCcrUd+9RXGjUuAMnmJYbXvd98dGeCMbYBezsH7/
QdT05x7YVw/nwY//99JZivbNiNHJQ/6J1o3yzDxSnkGfFNFDjIyVMQmqelNNGDQmvX9FUWgnglaC
xrYidD6pZ2So9gTgWzC4fXKkhczF7WZT7hryJwgG9keLw05CABMCyRS7LA0L4sfDc33ebJNuRRbH
2yRmUvUenHMFaG8pS5BQ/TRcPb3fukN3BFjX10N1Ung8YRbcONA3WfDpCwZqqIXcCxjdEEYq6hy2
D8TSKJlAPW+BlkXj4JRNWdKjRH6jwc1ph3Em7jyF+m26K9zb0/j9Lc45pdL3eKR42lHI76astSZM
1hV3n6+n/mraTV/4YJKGLNLAOj6qYjD4bmZpRF6F+WJdhPu69pwhEJGGTZyGgWovm1Uv0RRfdoPF
8A5exGUbakIlgA1FPY+dKvC48DpZ26qElwzl2HbdWZnspmlGkERgLo8sn/Ean0kR6flL5j6PkDb3
y2yyrXs8fLzd/RkFRxm0NS0a4OLHqv7g1mTj/AGIQk47BdC6fZ4LyBgryLlkBztnOVTHWSfJQU5w
t8d54uft56RoU+mKMhZeOFgonbkfmaEzRNTjqAHjLnoQBe0owcbZfdIGRmT+YHU1UKFq+ZVz6zME
A11KgaZzCPUzXuwQto4EdY8thxQy3qvPhpd5KapkzVVm1i47EC+El5zwcbcGoX8FDDZIP4U713b+
4xlcLXEkAghVHE82AR/Fs9vKSNe71NaJPfroZl5aBGdL3+5PxPmBIdCialc0o2cASW7Od3x7AnpR
iVeIwNK2O9AgajQg01YKCXYKscnvGFTVEZvsMfqDNe1LPIGv332MumWomPM0ykYKAmsIOu+HuePe
D9/AqM3+VKkiF1fSJKbDPqPGdJGyj4DH4JhAA/e9Dozs8E3qFaA0NyP/qbttWUldMaeAep4GCGe9
zLlxUyUrUc5SEaEO5qrrjsapBXKgH6lOp5zskMJf82Vtog3tCKnw1kBNwSPu4jdPs/w056T5vORv
Ov42euCUB47w8kXf1Qq4k9iI9uPdUwQfmPBpNEJHQje6Hq1O47Hi6sGkkXYHfhILmZCL+N+GNDrY
w3vEki/TPIgRwRKeHMn0RSBlHfFFhUEL4OUNvr4kilkvBG3hrBEenEfCK7Lu/i8PswvoeMaG1JGE
k+afWDvC2XCdmwYamtCAryvUSARhKZlZeugdtjzxdu/TId0fohj/B10V3sQ/PXlciD3CalcTTkL8
Jj1RC1phfon0xNKsjEwhUWN1jgHMEGJ5gIVInw8kwYoCEqT2KqxxnQJhZGyggh0cUQaOYgAHeIOJ
l2CymMtz/CqKiLxXuWRi/FBnjTPmmNKejn+DagOcTpzIG3CbqY7gfO8SPalmHYQx945i8CBJP6K3
57hVNPEfAb6zLKMYp+8Mi1ds3owoQGVztbnYVYIlRGJyKSsvAP6Z1Na9P2umxz8PX6yBq6ziEwEU
4HWMSZPNFhCwYm+lMIXsflEkLp6+vsIIaWYtapk0x4g9YkwdhnCrKVvJFn/KPKPVWTVzhycRKX0T
AnvM794HHt7mzmV+pBhd2Q6tANOwoyRBe1VYlBVjb7acqZZhoXdDXcDl0u9JGujqwwuNKLY0d2kn
x0ngxjByRKniG6zFV0B3xeWYZhJmcLfTQMj8onxnoavFGpydLeDp9TkS3pmAHiBZGzjT9Tb57zQC
xryfA3AVKkYCF9E6wHNHJa/D2RUwukP/471NrS4umRl9yFLuA4YjpctGb8q3zy5Bvg0l5QpQLjMn
MC1AnlJ2vYMrFHas7uFV7E0vDFSxiA4ac8FHDDfJ610CJiQa9anuCyqzaA3j02ENoAmq5s3R9iQ9
1472Z+QNvaWLwH3pb1YPe6hIl78bF+yXx6fmr7OV0XgwStDtdIrJVN9OXQS9n+yrkPUGUb4w6jHM
DYNnjFNhHW9Ypr9gbYBQ0YTQJ8US2BIqSQ6PlsLEPfWx0cSXji6V0lRXFXpWN1f+FnnY+jbcdWvW
IdwrnM/6UVCJDxzH5VvNIIjbuamsr85M8ihj/kntxkeq75Car7pnvJYS+cnKDWPisL1/Okdjg9YD
vjeXWC9iUWGruy+tdzGfpeuyWlVpbUQx6m7GvjIuK+znm5rxN0EulCtRQ1pzCswZop85gQ07rlxl
jRRmeak6pWD7TR9PqtVmowSv1fZl75zQ37uMNVMolE8Ly/y9zcjzYagSZonzPxcXY61TVZT2xAJO
Zjo7uG7ljRlhwt9MdscVb2zuL1PDBMMnihb4XnE9P/90jqckdNZ1kKIyUs7xt+CJLiuLL0vPxrl6
kH68KtNf0EUAjBdCICB19KAtckGeUU9eg4ZgAW6idJIX8ChQksKAhd4e4AjBrHPVSqMbf+mg6328
vvTxAElm6NboK5n6XQ+PWByN+W+8Y3f8XI4xjzE6/7he3bZdKhPgQ7CHaBdVDZEJ15lhHG/capn/
7FattYAshNFcMBC0GmRcYjPQg8ZkIdayILHiH/pihn1A5aclXv4/oi4sVtMeeDleCb0zpvn9Q1xz
uQmzy7vDWM3/gJR1esp5ubu63UAbv4Gh64u738MhT0rU/6dfj0z1Vtbb9Eyi9CbB+zUyClEdqjag
MGsuK8BiOLZhNS0ZTaoPEyi7BfG0WV6YZaIuYoYKbHowIpt+9GYDUKbqQ0Pitdofw90M6pj6F1Ij
FI9pjq86V1d0fDb7EHheNlsjJHycOO7RtwO+f+rgLLThCL9zxR+z70ZRKSznBraicQmNV2lXpiW+
yC1iy16tGm/iY5SoKJmvb3FcRCjxlmt/l5y+L9e5pY9XZJqupxiHA2QjBqayfZkQLLwThoiW7aG5
PsKcxRYRAAgzPbHx8OXbEPhY+adm3wTJS58ogeIqyxXeuzmugHwcel4Yc2M2t6/9n3dVK4Eg+LkM
g78CL61ZerNmFjKIQ7+NzFdwqA17i3Go5qKUraon1ZKGEpOQw81r8tQB28ijKxGNS4aW82doajvT
WTFqteTmGHJl5J2hkyy2Dlyqrqjmh4GMtIOz1M07rYejpztdUHgF7YDwqr7q+NGSi8UE+7Kz0aVX
c1OFMg2o+G7Zr90CglPkIG9mG1ZceiOBb9Obaoy2IWJg5GMZI8HvnxVv83zbFinDr8HE8cuCtmQm
L7VdYiqmuGEdBWcXSElsIpuvMJ8v/dlj+/Jei7qBI786ACoZIjJggfyh36m1tOn7jBp5C7i64n96
Nv9VlwXtW2sE8qnktB9o7PV0MOdAjpcu265R3lIp1i1fkJFlE9F7+cOZNnf8jnRPPA583ovfOgiJ
HEvZsNvPwh88ZvaxfKGsz8DN/h6Id0FOb+Zs51e1EllnZfC6nGIG/CN9iUjCLA4/SCQKe5WDKd5T
jqcY5kQBqppUhK0jPLFrr3DmEimOPLyHs1GFy+lkT0KN5XfmDJ9TJ8ckLwCDizRZ+gY1e6a6gZPx
J8b2mCVLyUqM5HvVHhO+SLGiFr6xUu6tQa1z5UuQj/OtfP13fWEFweUE920RX7n9+IJvIOkmmiD4
t9VgjlELvsOHyIpgi8LCidywTnibU4vqquW4Xb4bAEEHpP/EigQ9O7KfeO+XF52jldkV38Jybrbm
MK19WzwseBrUE1z9CQpAfzm8KMiIgeMTHFDc6FYzcLq3q5j4SpGZZm5iLUgoeKmszytSbo8LZ5Xu
49jvUv9n8ZGs7eoA374+E5yFo1So/NjsD9C9uMwrBrQFFCew4rIugwCiRbFhvC/SlnD9zj5NpbsA
7lorCa+RuEcvVchh47Gmrq4HqG8AQHQE8KR3f8Z08Gflc4QsHPNrB1xyA7p9LocJhP3RM9Ms9PO5
mFev8QvDeEnzVWkiqc7WoW3/ukzQIoOTMiMZ7jIAw0qWM9jWePt1DykvrWMAqa8ptmoPlay/8FP4
EK1wixyrXc2oIyytLQB5nlw/50r2xvC9qrOd0M7JiD6LLWGyRT72PxCe+vM5aFHgVZheX1pda4cn
SvAjSnRAy0npoHJM6m/TrChI+1B2jqm4P1nAPCMCcl6Xcw5nkLroU68Sh7s5XwKS7JYyLxcc/GM9
vyZUGti2Cm2txU3CuyN1uDBNZFUw5uqBfcGvCJD+cEahM52IASuas0l/fWgAXGa8AUil6qSWiXF1
QoeELUgqzK1bM/ZPbS2yB9PVmM4xGdH/IoMkNp+wRQ6jN6PfdSaTkVDUQAb4NmzGbRTgQYDDltuz
tVfBWwXL6sX0g+4oJqeH0hT8rK24A5cwayp94/jPV5lKOFFuFezzUtqKQHxTLyDb8BfHKduHHDqX
I6vqMCJzQ1eZY+oZ7AhC6h8VzWPobhgwrAN1iHYJ4qisAZl9Ho+XlXqgcFPJBBUXjamVYrPvDzG+
5JnqPcXcHkmOZrdc70Q2PFKeC4W6N6tiR/6A3q5lsAOWODpNbu3p6Z3txhKoAE1GN0gSiw4wI+rw
C59VGNaUtPUgRiY3daFxT4mTerMZA0At7SaCj5npv4HokRM2Pae+OvJjmQdso61RxInygk0d2ZGW
XRRurUXCF4Nau4vHq8AncwdAcefGRRqboAAqEPQfHQ7wZN83HyoiStkjqkSJjlgn8hLml0YWjiGZ
1S7RBylsJev+8kwpJ+DCV3EFXhMjgPKENtXvVaj7H80AH0SNpYy7fYD9PE8XSKVHn4mbWw+dlrk1
W+nsc6Y4lrFDEpJDJQQY258gU4WtYN3nyXlG8llEoUUTsEDbjxQCJy8cFUGoLiY61D7CIXtA7Qal
lO6E4mC07kYEReZ8kHEvSguNxYo/AjA3mbRevg9rYOp1fVmenbaZl1jSfSAhQ3p1F9Q55mxxzu7s
ezVbWMLhwNKvoEax7xpbiT9r9nstGmeIXrthCYyHyXrpNXC6i4C9cr+iZwCKdurCs2qPIz0uf4m/
f5eVcxvQz8+UxXKXDrl2o5iVIExmgbt22IHMlB6lm+8rFyR0RS7+1xeDvYz9Z6sZAIwiqHx0OaDW
qdC4F2AmILK8O1rB+y3mV8rWD2tWlDf99bt2oh6W5+hwnJEubnmliCcj4vHx6dZ/Z6nq7npkdiUA
F7nuIEnzbsvogJsjIycuHg364IZO48dYf7Jp957FRMZPNje1aQD+V5Funs/nlyEiaiav6ZaA7PLu
Lzvo/6/5BRWuBvNo/z4wIWyCPajZcN/162i7m4H4z2ID674xfUKrEeJ+pxMEBrhVu1cdtSXekGTn
1QUk44LEaYGDzq1YAA5KuusGhpta5YYVSHvNmkAa9F75Os/9rlKt/b+PqDLntkghWQg/eA1FRqfs
y16eYjSiXqom5gOTeY6PXWOf5AiMgwdIfSq+/rwRkfXjbq9HwQKv7YIfom9h4TRIPBWN+eX615yz
swVJVYWRrmzvq5BWKgNS78gDYjhr/RBK0mFv6+F7pm7Y/Fg/dEuiFShacKqOLkfY4rkpIjKz2H+U
C02H2qZW6EnzVQoiQqBNqHbAcEu+PAVPT5rX01KLm7p8CzRHais/J3xFYT1GHRmX+XR/Q10M6t9G
i/ZhF2EEuPQSf88Z49BvWjiQnCpDb+zULdf8EKN+yExsQTkxrqi8UuIfxiN2iJ0s+Cl1Q1lpE4Ts
ywvO6cZiQv/oExQf3vcrAjiaicqpa2vdDZ4KIRLNdpX5Q7mxu4SEavGWc8MootQ2afjNBikVTLTP
tNMYBKVdHNQCGbPPFIAogb/UoEqHOWX0NqcjfciNYptHpNVmEceM6p9d+4Mmn785wuJ3mkxmiQxO
5lXODYUltwVJ1HQYComTjewBn7X2DnOkT+DBwTujhtiR6CZ/HpN80aWRoafRDgjgC6s+t5eQ26gd
WsdSk0kyInDYE/WIPb81bQZApLHOCbTN4rdwwsWcdwtU5sqMeyXNUj2vYYYmpXx8edkKhVd0qMmq
bd4Yp5Sz0hmRlo85pZCM2aipA0vWzOXmRawwsFwa6iz+O+9oeWILzZMHfmC4q6zz8SsJz1TslaSV
+oXydP5D33mwxa/vuuSjlQs9ZEUN73506hB2d2vnCyD3x5G2PhvwDT5KQtrNqlbeKHHYq/I7BlsC
2KKsy4lxfdkDu3t/G+Yymi2w6NyOQiCSNuK5uweW/YKlIl4jLaNOB5dzZHEXSRQKsvDn4/X3iBX6
suNljWyTerRE7V6y9PRn6WfpsrLuY9wDPLyp580O9Nh3MOo4ajCw3VzzsTD9OMamCzaQYfxtSUiy
FSTkKI1EzLyI1N1f0tdc67PLca8noSNqdQkAm3LFnpXBvWEehv4emZ1HpqzlCPrNkbxSlbh25od5
Ma1ES1XKBMBFneOEs+R5yDsP32ZZtSDClGdCtYp0xW6iZT8xze5LBGITh7smNio2estGkE0NGVLl
bbfCGi19KiPW62pKbpvGBLqyMY7o4KGUQeFdEWhD8B0B4NUS+ddrCiRlzAwznkvLX4r8uvCkqEGa
S/uZ5XCUFlahbDEaG8pPyRZJfLAMKcLmHJqXQGbQBmrCtm8s5q/b3+Ee3PElZ8+vKXsw7dNC3L3i
PkS9qM9PQmQfEyHL/+xajvbMPBhICgDXsf/I38JqdUO8wo2SopkrRvMBaiaUFiUoKeBS2u1RLGyE
CKFVpvEDWIsEXMxB0SRdJemu8uS8/SH85fvr1DbbDekLbB8i/7G8ObUpeRDPMI9RUIuCeoDOTVin
NcoLARkmqBbbpTdXGa7aVHjGnHpDuX0xkuLXRL+KYKRHlZSDlz8sXYk9vW5d3KA3deSmGegaxKi3
U9Gyw3B+7tb0cKuOa9RLGSzlEolYVqQOiAFdf5KmxTXTLGKJGnBvGZWqazs1/cF69mOnYE62/QLv
+1AJwxNCKGS8AHxYefhTFhfbFAcposbIq7r0HXRF2eK+HrVY7f8Y+R0sTKxSjjw4fMr/lk8d8jDJ
B209GmMGBsykGoADXcc5tggT8sj0ZGmd5zW97A7w7NcsFeP0C+42o7PuR886IW/WOugcFTA8v/zT
ExzmwOvnu2mDQ99Clqvf9CCxSvTYe3U13SqhQTKzOdiLytc/uhNmHSZuapG2D/03cAvZDbSwXVhS
7bw7LcIXo15p4L9TBXcDHUaOtEU36v4ZCzkCrE6QJrbKv+HwWic7iD5PT+LFS3gjxfuCNaBCP6yS
QYeudAQKqhKwS5rdPxk5VBYGiPyqT0lsbRyD9s794HwM1/f0IGaCyJk+x9O/uKEa/kfNk97UPTMB
UVQM+Ow3ifZeZARq/85lhVesPHW2sCidQNjav3muTCC0Tt97TA9a+GRGLu8R20l5QU0DVAzNzJbZ
G00TtwkKNwifksfKov18M9gfUoWklFQXLr6OrGDMgxmoYphl6WRSUUSfb5T1NW0Gv8aKQdE7hJqq
Zz79qwQxce/doSSxUH4jyKgR+YJ/TD5dSfd24uPqh2KycyDc50hS5KPni8rUogZSnvAwhCk2h+bq
XqeoFUN6kaQ86yrOtDNfFcpLl6hBUq8Y3c9qUw1aNs30S60vTSmp/hEHIzK64b2ry8h+RvCA00FX
hC9+Lz8WAnVxvE6NCkX0dCJB8emVJwYLUvo2+jw58OuhergsZtSrThkg3KjYUFybNc3n4d5ILiO+
0HWUgCFYqi1lDakkJgw6H0EhLRBgBalJx7TJ6+blYPtC4hVv9XAqe4oMJrJq4ED9YvqA/2yZ1/+P
q0ZnQ3hxU2ZARZJr8LsnIBxTpIwKM9wM1f/M4eIfGbIzyDAzeKFfpaYpRP7ba0eYF7Qe33SGTird
sLEDYKwB/E+AgZBpbrC8lqAwVuS5s95zcmNVgc+G2m0X24XMHRteea9rOgkp3Hyjp2YlKVgOErop
yNq5l1SujkjMOSRA4EFwE7u7oT9Up+pSTT5o4yxwLJwFrqmsmNp2PS0N7kyTEAocDJs79sUF6LxS
JhsuPTE6xUieQFVnh+TX9G08xunQDb8pJNryyVhxhnz5CDHNsGsR/+MM8rJsU+3StFo4Tj8enyrw
4rISQjmfRpFMYAVIsI3cNG+iWjamHZwetvHfWIK421gKKS0wwqKJTLsjgL5wa+H0cTD89M00wVrB
2xtjtiz/eZK1jSaauzaw4kF0X0aRQXT+Tif9cZ6+NrWM+laHhdihFokt5Vvd80bPlcZ+KTh3t/yF
qw5J4Ufl5Z2I70Ll3pSPx5ljqf9xqUTbu+5NQ0Xt+sQkd1o4VVANhaBp4pUR6r159FJfO0biV9QS
XRAAZpMuSTG+jcFk+VpAlqCRgBUkIBfMUX9+FLuUi4wLo8OLcJCWfIfY7vlj7NfvXbNeUPCcSMQy
lAma6DwHV/JoJuiFmRqzkTgEBIj+Yo4P0OiRS5SNVvmKomMiLl1CuoFoANKYptRFCWQqVVDS+Z8d
h5N60FBu3nN0CYn7bdXSxsaSMZY2XnT7CSol6yfhtojGbMY3DnumpLeu04u15ZJNbI/GheSIZ9Ya
6UAG5xW3wfSQ/E4TVwmQPR1/tZaI8YR0U6zkwidV3/56yVvm1LedYRUHc/ADdNIvDEs+owgXVJVv
zgU24vzNpttx7QYN40vrevQOr4LtwbrRzIfy/L40LqZ/9sm4VgAv0R91lCHbddSlXHb501XZWOjk
HuAwSwW+TSX2OqAQ3qnJhDdQDb65lD0hSL84A5g5BdFTBhpxww48cdmWGnLXlLXoEF5+BhIi0Ejw
7KoeXuhd7voMDxdawfpQwPYroPT1/zvwD0bxD+7jIhO3Adw80RcvWK6xB0od3KWyk18zTxDmFsp/
3E+4HxlgxxwvrM25onLSkt02O5HzHl1uXE4hVWt/k2RucrvozHmOXH+mV8wV/UChJgg6h4t7hzHd
YI9nHLFr++c58aMHtDqMRtMMVJMT5L1Er6V7a0QtXQZjcaxkSeILwNP5HdwY0LbhN2FXQ9peIFej
NVZAMtaIOCns4gQz40/oru5vyMW+WFGpdrq9sdZQ7f07mOCBdyOg3VHvomsvF/9oIVlrITO7whn7
3EqBGGRjB/OafbL82HtOmPNNnDI2z3/E+GkM+kAIZ5sDjdkvlMw8oJSGKhN1v8vN1YH/b7byX+pY
AHcEcQYjEXO4Q/kOe8fkWqkIc09BZZJ1hYUb4ffsBNC6JFEWi9IKV8/3LmbQTIdMJVyCZaGUPLio
62ZabRRtPmq+ziAYXpCvZbvxTQXoMPgJYnXp7ASF4E5YM7oG9e7hi8S6JyjqcOCJZLOeVarD2Nmb
nImMX2J79ef2JGFypvJzt8KLNs6r1ovZWkWlHk9IH6poAYzaVXeAzBO5wTEq+m27CvhtZ3J4jiDK
efjpmsfO9e5VofP6otcPGaOoy02cejrC56MsOBFedqtPBWuX1v730CNDT8+Y7N2zgoW8T69FnqxN
8EsL64axiJuHflaCwq5sSd/FeCXaZmaRPDXkrjoawnqZ0qLofycx7tzHraB3fvEkUhd2RNFWNEya
I6UWhWOBClLY0/v1tG0zBUXdqaTSiYZcYxoEP6YbltSitm4j9yoqHeiSGWpbexdsYAc0JMikioky
3KhWc0Z2I6IL8/bRtSuwfbuuquZP6HR8/ENiy4UDI1jMStNPOnkDZXzC9Y+W9aMiDoA9kjJTJuxE
FWFvlnmBiiqBkApdh6VS3iPClBrY7E91EZLPyegon4hO7aoDOF/e6WfWfx/Rr5bRvgY0d6k9kMQp
I4oGZ9WjWBStZKykKGNt8W8wupaRIMieYTuqhLys3q2ecg7HtlPuZuHloWZvVPecwQguJgiQVbOV
d7GcycQ6RwsuzyF09v3oF3ELgD8W7jJ6qWwdmscYRNZX9Wzn4i5G9RMJPLYQBSASUNQnuU1KChPo
x2eQ24DWrDBtBoANR6rNdMxR0tAtz/Q/LlsNaiiY+lDZz34nrWfO77FnT6z+cqqozdyX+4aozoxL
Fi5UJdFpju8ugOz+oKBXTs4RiZSeEAfHR9B/ucTmyNV8w2+5LyFBqoePqqBloZzsCGnfkMJn/T0d
7UtGsO6eIC8RirWokWXTq6MS7hnsM5Q7haimG6atZT84NugbK1fBpC+fpy4t3eJa/uSSEBXBdEid
IcmTCP1Zv+by+ZzqDWSJWjgofT42Ka5ilGnXYGDkwFxPgc8bJOTBZgf4sJWIBJrfgsLP6G7EDOVp
rPkmIlUA+O7G8tzRNjCdzmvwmxUtp+RoSuybXUodkgIcVaLU6y9BaUpcUloTmdN1Ge9CX6bSvPOK
/ZWEj7N41CI9+sGWjozMBtTaqPdlB86WhZTTlI3xOX4Log/0H6SE0kBzg2uNV9JH/F+FftsAD0ok
RWlxy92+Jprb3HqX+cKYbwaFttOGGo0EXPKqSG+1sswVDzqT6/2UPt3LM0uYZnC/znVNdtmTf+Yz
xtAJX8F7Pl6yDJGVshQw616HSSrGHLjrjS7gdFKZQMiT5D2pSbxdjY192IeliO8nLa9cl/4ldaSv
b7KW1CCMaOFyeAMiURJ3s4jukTB766LubLYbPb3Be6plNGv+aEktApRV9c78i0QgswJG7ZHUjhco
HGAnvbsaR6IJqaSkbY0VlkoEqLNLtrhcwB0jBUM1dcfIcqjsklVQYBWZvPP3PzSRBi3Pw6dDUe7M
/ZNqHwmfDb1J9g3LPsqp68UXGxU20s6r1iAFcHFk02/U521NcKoz5fOKB8kM+W5FWDIUELqjv0jZ
ic8gdFIjXTi66Ivomb3xdU63OeC1DQxNUhpCUdszZ0ld4tb/ir7+glhibiJrz1YU8URfHSD6xsoR
vQk2MVxAIlVY1VD2+14gxNuYGiPL3V0dEd4DQdz0oNYmoIR0DJEuskit+X9WtBX2hFU3G9dDTNJw
EicgdjC4W/Bxiv4+11bxn8ECcn1uAcvUrLRE5f4TooANn/wSofNh33gu/jcSRs3tFsJnOS71QmGp
yUAZmZoJK7JDLUV25scA0kPuBlGEEG7SrcRXw44/5Kb+J3Hnl0xks/5rO2NfNTsNDetBHyimfk3B
3vYzUntpWwb/tPCByNWYw3zUe22Xyh2K5H+YJjqvn5tld8DIhrb6EoLkT9XBfWIY8vffuKHJ1BoJ
gY3gVAmUHZAspGhq/1B6P6H0NYrXFrK8eia7iTZPQHELKaoV7aPtxWMCAH4mLlTFoqtNuiCdU1/K
w3v9qTFD758gjIqk5IoL49x2xUWwBi91Eu02uLw4H8d7C1Vmvp3uivVI2vOUTVme9RH9wpUFRE2D
f1to4NU8KAJldBlKE25V5CkpmaHBo0AP2z7k7Dbm3H/FswYae9jXfzpsnhBux7GG8j88V+rKH35j
1JEw95EM2/lMO66fUaf9PYm+g9SzXj6Boj0wyb1Z8DMXgUvBuez3iO2Hac6qDtiYCya3BnewpXvG
/0Eo2z+U3zF/5cFhUE5aDnCeIpCFGdGKdMiK877VdIHjsEGU3UCdIrAttg0e1+T74gcI1qdaYX0Y
ZLZ1avpTSKw6A8AB1cvatTD/vtndQ6Ae3PjamGhOSZIuBBXZzsdYbb2OUsTiIQWhYPmLBOLUnEeZ
j4GE1aN9uC38pIVzzlju2TajrF5IYFF4xeBAfc0q2xWdgW2wr+ysR6ps9BPRlpImpejsa1xZnbd+
xSQaQseQ9/2dUZq4m5e8YeWYqzY6u7kXYHSmRP8P+ZQnNhhiHZ3IPqvR9CSVj7rvfCU6/qBRKm8C
CWi7kbfDeakdSW+JT9yVYAVsN7ZWRG5hHQMqC/Z6VigR7UcNIgvgCE+9ZX25cOHhecFkpQxr6cCh
Oz0krkbcBf4VOPDH6SndLaq2+MzJtIaGL6DtkyzJ7pv/vWRzELrH08XPgClk/sT0TDz17TiCqWIU
NVjrOEN+xq7Cw0uUQarscbkfZ8oYnUVhpq/rC6zSmMZPSrvY9/NsWQGuPEljrqd4s2ELncwmN5ao
llQYgHw40c5d456OMBddG1ARxYJkkGIbRJVUz0NDaO9exzWh4L8uUyJdSEXdLf4GZljUvOKxkwNH
NwWiD2WlqDJbf1rn3CqSejzV5/Qxamnm9g+QmjMc0CijZ9XybT6p2NNyntp45S6XCgE+BFmL/+Aa
w1CZTlMEQxHQzhKRfFLx5FeesTchb2EC9YosZWIG0s5aNLf6d50Hk550OPjzI+vxwP6EwnhfwYiJ
agd+hjgaZWswGRkub8gsT+K4O/urxbhVhqBx0ccQ6SJHv462vHOWJcU/1W5JxneRDeBsw52j8UId
O5Td7ECrNazmCCGqmdRDhXFiGhV3LmoCOB8KPIt9kWUqkrW8FRTtNEHV7cDEpjng6DBhaJpOG9JQ
1xdQsFzIg3IlHFBvrvYwSEyZq7LK9q1U++umpBoca2Nig7leGEep2pO0vrznIxatEAorc7bd6jYu
1VviYzLx3xibVgC6HIKY5e8Uw+MoY5juWUHE2qSf+gVV28fuK07TlmgAlKLg3VSNeT0aWiH/liZS
Cnx+0eex0YDZumiVEtKm6pj3zHo0DV+8X3KuE0/DfmX0wsvEUhBamC2dOPZcYbPoXmXGrsoVWwAL
xzN3kZtbA0IrcDvl5Uk/1XW957XYZtpXjp4/KxlFpPDEugLgOExf030J01PJRpGdxa3dW2EUzAQe
+GHmfj0e8UceUWNt1fhD0rShi2iiHCg1oSSeCeZNf0BDezYYeGeaoXAMynTusKTh1oDtqq40Vtxu
BA5xMzb9Mcl4HrD1MviUS8HJzX2CMUASQbM6QSolYuwt2i0mAOG68t3cV4iuPslbtIkXgRXskqwf
Wq3CxLi+5Tv/y/CPjwjgBkfwnqDkKUCcMaT710fJC9iPrZYp5uTXkRRtDaUsQayPAC9gzr6X/hXB
o6uvrwwyd/1BzN5UdKqnXJ8lK/bWwy7FR3GMXwRHA506L7pN4Bh0qJxbcWnhCVAM1C/Z7SvL9LQN
SxV+ZGcPA5Tf7e+i3nqss8K4Tdz4Is/wCPqn5qqrOhUAoZwaWZlr8b/pGvpEkG7Efl+CXSR/+MQH
4svRI5b+DGU/esCiaPD94HrlwKL1XMvNRV3Rp+l+vdx8WOJut4wQwVg7uZEHM+rU81Sw6WFgzDBx
W7QVWdKI9n9JHa3pZYIa5YIBYLAdEnlTYKgTDM/xwBKUOGz5lWX3mknGGIACpmN7NQZXbTJgBRs2
6gPPa4I2NpIyG1TmOOgUk+8KYSDgkWEVQFl+MAt3jNv5sHw078WBW2ZI/Au4UijYP+B6z4LoOU86
N6ytV3ku8vbhzdRU9aesgKYI1Qp4L4w6gjUdy1HOPG6+pWtIIlgQ0tTv59G/JpAhyNnzqPQc5frz
4SbX6RUG2j3T9cuHw/FtUBaM/xSvsiTGt5fw6cAhkzMk+xrhcRPrKdBVtN8OJdmVtmz5Blyziwwk
2nln9eaIoacxPiGImAjKymueSQf/ufrV6XIGLdlQ+W6Vs6rgEgv5le8IJFAGW8I8u1fSF/Rt+maP
uL9EAvvMMXB5Xejy1ii1C7xxF6fG0ao6etv895t6qLJpiKcWWk++Hfs9MpFRdEOT98IozLs6dcZ9
dbcVuTd1+nY+arkZMFezJ13gjwCaWRD6f034u+6QdYfjUxtAkwOt/AhIsKvjxdAJY4V428fHLOW3
ReQIIgHTSvVv+svYTzgEfUHTZfvddYZxh6qmuafKmQHr0iWY0eyECymf2BqidVVznwXl0uzekbt5
FxICzN8911bL2qs4/s8Ug/WkepDW9YSYk11aUB3sIc0pgk9UNEAQtQLUu9l3levefu1A9JxYAGW5
ldU+rlpEKZZc+ZcPcqYGnujS6Nc6xzHnJLqEXRXclHCR41r1N4j6kglUYyhYcX+QZ0iFX3EDNqSZ
I7ynGyjmvjvdzb8Wnx6KSR1rkAHH9p7uUCBKfS2bFtflqr6mvDwCawv4QFwnHG2g+nLYIehYrUtB
5jNv6Vm8Si7isMmcmUgpqMeFm2RtZJy4Zth0CY9PQxfHRdnS/s0AdJFvwtVbV8XxYhgjAIopvoJe
qRcmm/tM3hXAtQoaCviKLlbuu9LQ2cAqlpKuRePGPhTyXv0AXyHNJ+i6qhKJ+hbqu+9utyZg/KfZ
6e8xTLqjoDL53Lq3eV60cGQkMvTE/XU0XG6UwwqrChatf1fI4ugjMukpKGUu0gSPewWHegaba7B0
RZBvd3wvd3eG7h+VTEvDlSVvRLWfMG4e+k2LsrRdA5Y1+HqTmZpEB/+110vYVNrvabsDZjqQb+Tq
ty757zq4Uc38sr68Wdpxk8kD7bgP/a+Std2iN/n6UDwlmSrjINI0rm5SCuhkYczO6O2b4Ww28EOd
+BMFTpFlOJTyCN+EdCsGVIWcNDi4WMiVVr9JGLXAVkoBuPR881YV6+LxzjbRSXYeQ3zt9zSPW0RZ
I7XFQpisnZwvF4jXYFa7AU3fLbbj8B+F9jjccSOwBhuw2FX+ZtDeMX6pjHi5sjHOn2qSry2wytFw
KzemDH+LFAEJpXZk+fV6VtByAVkWVGBNyB54qhn4vvmkbkvuXMrRlR4UPZRoi+7WI+Gwr0D4neQE
Rmi55Ni5dEAyLNyhne2S7WgLBzfQ9+MLni5e+IP/kI0JM1PSxAVjN8y57eC7HggCE6N4MVNeNvkV
qoJCKX4j3lUx+M5vWlP3yyJoWeo6vm8jTcLbiXCidc3G9ed688HMYlUQV5TExPdHa+UQ5B0UgFYO
ioujcRhjptmaeRFgrivwP3k57auRddFDxVUVqeQ2tcHP0j+62W1QmGRqwVjud+3haH90xfkt8D/Q
mjFqcvfXJeg2vhoqlmPcWneC6svKxxO37ZOqglK3LTfDj7t85uS6/6dU3vx0K9hVlboTDRyBeRrk
Y/5sR58IHJS18ScF6DIitMpKuvm/8PSi/mDJ2QHaKqsREyNjSah6iWfeVly3qLC2aZMaLWN9hAAO
CrbxCcnUaXytAyXqqo0jOxCZXLIjG44FvACPFxuw1WMSUadMB5VtmYb+E8CKru60Pmw/bh7iavar
Drfi7+++YDC3YCaBITfRYKKEut+UWS7cphBXUO6ZTPyKEbJ+uWnn4iWwb1Cz5+4w29zQpOp1TJ24
ZRk7NLC2wzzmcMCJrP9uhDwLRZ3QgmXBxJJ/iWCFwIDv32WM3m3izlBbqZgiWCdC5Fqtl6bvs6M6
GNcdrcvS5r46wLqdRPc2C05+cQY63nj3G5xy58l08APgGC82T14F9zbydU+loOGskQg7srFAlrhD
TC7kkfz3p32KwncOQWpLW9n1f9iLW/swHe7Qlqr7O5KoyLegM5MpU9iVF8iMW/NY1Jvcr6XpbTTl
n255aB56ZvHBMmi7opIIAfpptE8PccPrY6Dyr+sLtYlUBQHApYIwtkEtQoac21k1mZObQM2ERkXI
PBINURDt6i4t+cW4x14b3jcetTehO7zdm58Y5BPXyLe3LOSchHSFbqDAmQc5V1LNHGGy1KhCBZ4p
zymxOoL5QI+7lYkp6qfvKOBIqBKR/Sz9YaK0v5x5kOMvPFAHlJAQ0r3fsHGB24A1M7+amF0SW+T0
lqCXMoaS8e+50CNVAnsXeJ3/rNkcWL/74B1wQJdDsYDbWlhpQqpYR/LL1RHHRmz8yv3PJwukFM80
IJ8u6r62ZwkOJZgUAd7CcPhOZsxRLSycnd4ZbNBBiyQZ+sSGRsJrL1azbiN4ajVPQV9Z+FXJZezO
ZIyvKYntRx7ti7BUJO3zA1WAo47r7717QTPPut1NHQhdzY9AULJ+zfpU7DPbOD8gx/GpD28tMIFO
sA255AP3gn1Cd2rzLPH6DvqM4r4JzKaOukEnDQwW6V/nthWhfbihbIDJTFvu+UQqG4HjWusWaokS
BbYouEUTKn7LTk0K3K+daiOijCiSC5jB4Oc0w+1EtkYScjh1balWQtTZlslcdgzQoOuXx6vSwyeB
mPnxGSYvRr7vTGzmtmGPNv2pvRIMAPxkfWxV0MtjgEuiyv86QQZ283j5TptyuxzraZAoncQXhVRc
/cv1VgoMHTY5VOBsWC/HCOex+4Vxma47Pd4F+U379LK4w70zEDNlxXTPvfk0Y4H9wotvWwf6/92K
BWZkJI2RXNi2j6yIxb+d6lszT2QDecVwLHfWdKR6ZPl+IEWYz78/tAMiAOq3ZwpCBHgr6tb8HatE
D/XdYFh9SX/siRiKZxIsQ4S65+pjIi0aqYvlPYntl15K3WWP+197an1JgwgAw+n+qJvFnVwbbHfb
+YgpRZe+gZy2v7USEb4oCS/vKbaqNKKs8Oe6r2Y65O8AUnutQE8z1bJyCRa+Ph2C2KJn0HkZ2O91
W7XWCPRDpq656tVFiNS/eAMCfXoY1cE0tkjbs0YUNMzHqX/5tidySgwVBXLwKig05Y0bZfSOWHSg
d3Z3sodF6LAtgiUEKzRLetSxkURs1NXjhVZzNSu8/UUkPX/42dXk8L0uACykyjV7T8bEVdmkNlLm
HexO326BnemvbLgtByzF4AABIPTsPKrhl4LFOiFWySFTfyCf27ND+QRsjt36XawKY8XQDYMBa//9
XuelYIbI6243V8XqpH7XAe2vBPbR7CihxiMB9BD4aOtCj/q7FK+Mk/8tCKtWdMJZX9U0VygQNW5g
0ev9hkJOwvJBamQR9TZI1usSoQxyxFBzI1j8WZZ9p1WJYF8WxGmepbKQES4ixmiJ1FvpDc0XQgRg
hyyL88KrlXd/WbV8D42uLtT9BgZtVXBqZ5i+H/l3y8dyOn03xNJRYqvK0QCHI0v/npdTNwqvBymj
Yb0vURLIN/UyzFu817mTNW++M4zgiOIjlpSxOgwFONhlW6INpMz9dgE1H1wgd/+lsLNtkobqZ7e5
nTNRiS1f73xFq+0qKlzjrCS4DJrklRfXCh81T3kJKeqCjJa5+yj162IR2MfvNFig8iJLkgRr84OS
wJAAAGEB3sPagvL46CPYTTBuvGTbQIl25XSqhpHxvOQ9FpCAJIgWPqK1IKwAtBP0WDJKs7IEJGTv
YInuadbIRrYl4sjxyFqc90/xSbuc9eUjfeJJeNsZfxsvci+dtkm8gruFaUuMoKDEkiFJooh/lsy8
HrMJ0h0cRyDJeLe8EU5SgTThz7n3cEYHmCuaDXwuQqL/RtlulO45X/ueMVgHMfMGBY5FTW7N0Ens
5fZd80OrddvD3PFJ4uC8IVQTv2rSefgopYzXy4hCJy4XhodMr0hFtl/HJEYZgtPB2gj4tGsqgSpl
wUe8ZqCAVKKnYM7p5bzrZSTiTFwHjvK29IuvBFKYKVf7Pm1yBUY0PYVVgCfBZA1tJN7Y8MV4pifW
Fbipt92a7btGAHTTm8+p8mb1ybN1H5CV0QlkJvN/6eb+Wg6xhvqtkI0yLFRmh84QOKEcxP3OJUwk
Yjk5tHPOS5IdXTrVhdbG7JGePOwG2l5flvztrB9Eg5NPBRwOhp9JHSwcK4KD/EnII36sfFYzMkc1
HK98xk04oXB+e2nByAATW85L2dVCL889Q8O+JIYsWtY/b1iDEB4XSyefXxKrgUxl5eYtqxUtDe+K
lo0w1iT+hQ8cfFaYm4mg8n6zrEM+d0eNOfBqksdtXkevOiYruxMIWbz3INOvJ7MoC3BQs1hOQMCZ
2IBqA4tVJkbduiD38uiKHQua/GhCEZ52Eh4hnOQVUgZLM1kCsWbaKHKG+3++Tz0p32XikhraUf4z
Tc9D402Shf3eOw+BIMXUDXt3Cz4oM6vQE89nx+5flWCbO1ZYnfjJWRIjsbW3NNqNAm4T4OjbeP5e
mBBQLePBHlUVv9PLSkg4eLUsW/YCk/9U8PVqxPjoUL9fYX/pERJg08pfaBaGZ3qDQXoCJ55S4eia
a5eg9vI6BpWnFbWQV40IzwSw9YYe7qGZmVV2+n+bHagBSMnY+HJND07ffog5OLmYv1MFTipBhtwp
OD+E/6P+/y1uzyRWf3LlsGwuW+u0F0+M3EDG+OSIpZ9kxE6KQG9xevIPduDZh+cEAiukvauUqUTJ
thqhMdSoMA+vykT61pA2K7QDmtXFd6IWdIeKRYARaolYTSOufaBoIv+gUbz9kZf10VZNSHMywHCE
RsP0dXLyjxWLI3lF7rOnwTpQ7xr9B2GxXANnLJkAbiJZgONHrtMwVsIHlMS8pNCl4a3LTo4tP1Wp
02gODO1wwYoC61F7vI4KdJByf+4CmZsVUYXOtH9md1pC5323JaOmbs1Qbc3euS5miT3jQqJU4qbI
MrlqmLuJdns/jAV0KG0RQkla6IrhA/yTLTsLvTt0JX5GstT146nB3Qgm+uo+uwq9RuYUz8d4ot2b
v1SLUXLplo55gwaZ3lHp8vU6QqUl0/YwkfXJnYSFteufuI1d17y0LJqdYnJHiyXkea2+PW0gmnb7
omGpkcmY0/ck7gakv1LUWbUY+VMccMztbPOKasef87atKzJgyp9IYMfmK9J5rot8nua3GJ0ToeqL
YNy5xxVBOHHPHiuJK7lYX33YpCkLcPWD2kyjqPHY/KByvDE8DD8w1i1OWXo62TzCyCVxQ2MVRZzP
nTz8S/uJIDAV6kXNJ9fbLU7pmC4zMVT0WI7P8FVzpjFGOibt9b8FXYluPLk/9Qj1CujdqnKbvbRE
QAZTT8+ZBXWDfgc798zEooH8L5YRJdJh/nu9TrXixkIkoswXyhG7qgH7nbwTnjxeUyMyAif4z8o2
EbFjX+8v2gb6P8CeHcPpgo21SaFZg5Um80BxPPNYIwoiOTC7cMNzYeNnY15PeJPxHHRBV4k7zVj6
8VZ4iTDwNmekJ0OqQzjlLlo7bFd61yEcHrYR/RWKgBR5KAayxfM8n24OXFkCgMQp/j9OWH1VnQHU
dEveWA5j/2mYnnrqd9s7qeeDLJR6jphmoCG+k10delI4bCjvlZjW1Hks4hiaCM6nArPWq9I3GDRM
tyJ+80O48oMl7xNbFYGn0J278ENkpOGIumoOdAYsnf2VckV2m0bsAW2kemcuLRMDz3GVglE+FVMc
umc0UJ8kg1fInVGAoPg218DPJBdfr+q/IgmjOBkyMnEqJeL0VCOagHQAp24cBuQGJY2+EHK+2r5R
f61CN0NekTAf7uo0Tqkr8kHmctwS/XGsWq7RbLmtb/nKI8jrDIKwUNUnDU/wLekCHnplZ0W1rgye
x/3h4T2VQ3CzxtLaUcLeiYAdxma4baPOmFKeeSjeSVHn92hZ4wOx1JyA6AtVJPyoeNlzFKf67+4j
czPxHUsEK5TGSVC7rv39oPlA0LEtsQa+v81DMMger0kWJnQ6xUPaAlc7395/9Ki93e3qEFmIMzG8
krnOCypMNr/mJFg/FakdOvs+jLmTbnETernO47hn9euMllLbKUPGX3dVQeuAyI2OFQnX5JzPun1a
82OBtv20TarVAvBw8ZunO1KaAo5FNcTkmOqP+1+kfUrWUKSPHgUmb8CxFy1Zl4uV1FEOlcTWI7Cp
jQLXjv22/PuU+lyjyTA5uN7YGxU5BHyoYBby1PzooIThw4xdpSPhfSDz4F2TbEpEn41uZxsos+qg
WMDhzqjYJr3GJVE4tdUiFhk3ryCnr17iygofB4l9uGAJafFHSGGEJVMCaRP2U8lWoznIYQ/I184S
DbxSPnGF4cge9GPjHcsx/p1qhgH1Iu2kZ/Jjt7pQM7nzh+porezvrpZ1JjTRl5dXySrhvN0ErWr6
mjw9Pm+CGJApNOKZNcJi4zJ/c3NXmKlZIbhl2xsq4K4BeTAemQMMY7BcXQ/Srcq3FurMJwPv/QX6
V0qGTTo7Bx8dlHWwlRgfkQZbvoZNQecSCJikfwS6VkGMzQoXBnLehNe6HNSZN7mAsj7WtQ/S45/Q
OFEuK11HditUPOnsx5gMEvMVK06nWqvbeNUZOU1D79Ahj8Kb7cZP/Nxw0Sue+GHyKuyEhT1KY5lx
IKeZdRI3WUQUxswJcSMgs0+UHgpviG/iXmbiZdbS+zc6kxbv4ZGdwen0/bXXS3WLs6GdjfRKy2Jl
jmS+Ss9szGN/EIDnvKXWWqMIvdqt9Qe7G0SjQjbdxagX0SBJ+Z1ndAiwO8FOVnfwJOSBjY+Xib0x
+bmJIio6L/bD+oj7vGnvYWnTT+WgXQ6EQ84KJAmD7pSCp/CUqzmcrlWKuL1hjjgce+2oEvEXSey/
Aj2aq6y0M/MfNzMV/MfSZVo23XVZ2HACUMHkJ/7Bj4qkubjd2p1oVod6ohZL3d3TYE/FS6XiF6rF
/7IkPlE0gCCsLw4EhIYuePToCyixvTzPqwqCzfLKq1cwu8TtZLQc4RfsUkV2fTWiGPywPgTPIiPk
1C9mcrklGmVF/AeE0WAGdIYyof2gqDx6SDF49GPiaCD2rt/fcPL54MsuGrf8gfZK9XdyJd00/S26
VRQjHufcxul4PjKbmmaSihTuhKSby1b4XgPOoTTm93dDwIfAqjdO1LRjT8HWM1LhpMZ1OlujK5j7
4yUopfOMC3PSaWGH1zIdxZJqWYQfn5Mw9fPVA21e6OTY5qpdWHe4lVYtggb9AVmcocSnSg0LRlIx
BJbSbmy7UQEA2SCcCqVxfCoAZ7mU4cWi7XIuDSyycgteu3YqrRpV3m9QER1wDVsgPSvkFowNo7j8
rovL/lMFa/GxpD1q3KfuRFP/CMIEYfQEFhevykMKB0JvAj8GEVxEXUVuouAmVb+z8AhULho6iGJO
2gebhImFx3wlchKl74G7GU7UYNyVfAi+QWj9U3rvbQb6tEbqJss+VSvYCrViSincP93t5oruWh8o
/f0Uu2nVSsFHcrpLsaQv4YrtnkT/+VBssuOZtm5NaV11+dzBnTP3tc7/z8SZgNWyp4rcVqztsk4D
dSpZJ9WKg6uOzNXaIwMXUqNlWb8m6Rc6OYwyS4Q5GEA5ZtowKsvMNb1cPEOe/1vHKiDjsnVOTwgc
iIMzlheiTWTh6st4vKT4MFGjkeNLYpcuS2PaV1yWS7+++2lvbI4XqOYtpzeJq8lKU6qLIidg1H+q
3Doau3jnysk1CoFza31lLNXNBXRIwTiYLK2fNBCUGm8PGECV5pqiV3ko8/qUUT32Nbz7eRrMG2uz
wAejqT4BoPVc2BIWi2fZLWFlP7PLC0ZI+fVrCY5+16JEPKTh3ugM5e47OtTYrCt+qkjZBp82ukqa
3bCtmjLpPoMobjAfQEUWaHKQ7Rx+7EfaCtJzjok8g9zgOxZPJvHdydx1xzvoU/kMiroiOA5YHIDo
iPbkMMzk+KGmy98a0qGcQd/CNwpX0rp2VaqnN2kXVnxDaFL12W+qUdvjpvWQeA1pGVCoxQVk7a0k
oOqLTNKJMhV31JO5Wfp/cMMEXIiUblGN0Ha8wUwUqLkPXeox4+Vcdszlfh3u3enYsqDzbrQEtipD
Lg2ZaOV9+GoIkAibZlXb8niiJngN1lHr4rSGIVI1xmddqFeVFptsiNG0Zs1AN8k6mpuCbnbJF6dB
Il7XTZUTn2XLmt6RyJMU4txjV1AW+/t0jLfpwyCK5Jg2OC/U7ASGJqJ7mGSvUGF6Jf/LOHQnPto7
xKdtXLSwQHR8RthmpJF7dDJ6YHk6hpNV0fQ514zmzkhULV2Yu4m+hX/yGZ8w+ZySCnm3IKyELpc6
+/rAbc9baaEexPd0/PkJe50MK3QaZZ2iAyV0tf5JePKnfpY/mIbTQTcaSrv4SvOa4pTTnzWz+CUo
uFb7u+K9ARYsfOjWQJS4T6OgkB9IxrJ0Z1SWPO7L5UoyD/bdQH5gl+/3Y8SiHFemNGCJZpuiKfIa
l9PApCMM8Q+OMYEcfOQQdXMumhNZxc5aEJ2dNZtWMX8j0KUSZ8XqeMReHPm28Eepa3m58C42qLjn
eokQSaQWs3OqoC1z2cZa0yQ63V1uzgJuJAPCUN0P3mrTEWEJHdoGJJE6uLXOpzj3B9DEh12Z5P9O
m83GCCXgCjNSMB0qM38RX1pvNy29v4/2JgvWfbeqCKRifBEc3wdUiPB09VxJb4muFrjFqLZnxuZu
VJdmwEWACNCYxkZhOBDYru08CDHruUbuOSlJ7QhpEMfWBZpV0BmSpZRvzn+9YsZe5g7uYe77Y6eO
m2OcPd9ALKm1OMINp3AtxvsPra4dQ8/dhbs4RsV1yvNQ8wqvMo2UiswGjGYA4f54a9TIAYRD0Ncz
FgUS0e5q1stMNC6eisa6u3DJ+lbLYLhNctwjvhOSj3xA9sw/k3Z35tzOUiOVKwjrn1Gn1roh18ET
jTfdiakKkC4z2hZsf2nBEx3r4KCxfLQOQmavFBfARF0EeM8jRv62CaYVnVN5il+7E9Zl2cg4MAna
vIhu6VEaAmACgofE/EO6kQhXL2y7Hn5g5V4op7t4bLc24hyUtMJZNh/J9tBOai7l1a03vtRj0LNm
7VlVGRKJAHOX0TMkHcK39o2lxeHW8+PKuoEncV6oXDj75rpZsD2QGgqEZIA3cwZ80S0ypgFhS9D4
OYf7QexUv9Ui26/d2i49S2iG4QUZybuMBt49iEV7HvoDw6AEzQsuaImJYuwDJLIOBShgWN/VIQX3
f9+Wk+fqksGtF5iBNhea6dBIn0Ilg+OHXOLCc7zqTDND+O121DSyr0epX9Ud5dQCpG65FCJDKVuS
L8BH3/pA3KJeykoh1zR15JNfa/fd0DnvfNKX8SRoff8fw/YNDZCPWmFzd2U4GG4a8XUE7D7CfHrH
C5eewyDS5RV9QgRY6wH4wZY/bFIzVnpAUAsOkj4gj9I3CqTsvDBhItYnkvOHH2kZtPooi2sdjZFt
F4DcGgz52xv/Cxeexia+0NXEoG2oETFPFwfawE29+n7ECGoZobSF2UZTSOyuva/VAd+yysvTREj1
ppfuIYlLm/GY72b3ZouFnUhHiICyITpF0QzGbg3HF1s/zTYB6LpuUUeQIYEndAacQKbxAtv08JmF
COXTapaVzkxgV8xfxSbfelvM2Hg5TIs1HQcNafsRfPRKUQ8eX6CbEnc/786Xhj3TqDcNRPHo5r8h
oNq7x6gXrL8R5kdmzfmg9THI7UTES9vCMDquRm9qtrocPMpULR7kuEq+o++Dh7u+rM+1l+F7ig1X
fE4nYa33wZl9uxoQ2PYCcXnlshGOukYhyMCl6VJHAaq7UswLLCYphvTbRt6/giS817m9Lavz3lac
EUfLLmkilOu4bUV2shLPxy7M7709KNMOf5H+VC/RGqcr2vRTmF25iKqG5xVgIXcjQnCUX/o1FQ/z
v/nTkY+wqYTyh2iZ94Mj3GIJnNhHhd/Ikmw0bQ1I+ouv/7EfLEWhApo5/4qI0s0jTVRaEF5+iNi/
NdBPVQrsjk51lUSWh5sDXaAicAdJfvjRh2mhS9l+mUOFxBjvCp1l2MxrfRWA330pMS7Z2pXQobN2
BWKqfxxqVrQu7KN9svGDNtGfxIgiw5EGRPdKKbebF16kP4AgJKxvUO15Pg8yu0GdcCKe/MrQfjhB
njp9zZSy5EhWGDnolhU/H+Icnt5trsYt5bOAePeaEVBCMoPwyeq1HgqMjghcT4GxNnjpaKzqrEzH
EI+hfoouATQXUDO4pontbBLJOnE2qq7pBt4FP9e/54csnInm7O52y2o7PtEEM7gcoNlVgYcsagyI
sHVFt4DdYrLPy/vciRZKadvXZDIZgS4wVl2obz4vsmYXMNaD2PUvLOdgZXdyWG0MJRctyn6WKmqh
gd0iSjLJ29/H+yn1k7G3MaTMZ1cL7CxQzHtoCGqzehaqcdjYw+vt/0wlPhQCHyS4c1LUu4OW4kjg
X3tVm9Wb7f5a+AaRpfHLKx7RehgRXnneCOzUg5K5m8lX+/lxHecPbkeLkN1E9iW3aTTCTNThxuy4
ZUW9OcXXDP2moscdYg++Z9kzNW8+/NGa/PdPiWEIn99HJ96hXHGzQBnGg42vuGpHNjBXEzWGH9ec
D7yR7VICceLgdHwE8NT3cq+4+SxEYI07Cc+YviCkAxZ7BEQGsxwk/6UhZjGtmGwgZH3oJzJ39EOk
JjdeK/5HAjdBSO0sCjZQ7AD8tc2eHzMet4ef3bkenmIQhSeucN/GWaHPunGd7ysfUE7Msxmq3XhK
I7lobVGemJ1Tq1a+TCRF2OTGRukoqxrJzFi3yFliXM/Mav2wbsfdLQ/4qQZr4Zq0KJAAE4kTtv9r
P2bhJ6a496b1E77ihEE0k2rgo+EL9L7uRbnBWo81HMdY+5uI9KR29WdqQoRnaJy7OlhoLhmp9hDc
G2zkAHEki4dk6c98MWAS8g0D3rsPi78CpuMWAieSwknjf/6gaExO8sPxWzbyu/idNCC6IQf6idvV
0v85a2LEFEAyNLdmFvhfQr7TzyL8DSvpUhuHzLA+EbwflxzvjA6Y930cg4GdhnSedYkpya17K4ME
M2ZhqND+vBsPldvU3w+/pPEitoGaoVY9WTjSkib4YuCVWzIJjO9Rw7UAIqnoZFjK8zqQSiie4fNp
8thiKZQYw5NJiXxX/C70KjgbiftaykxhBJs9dezyc8dFSaixe1k90r33MAGyqlVjrl2lFUL5fB34
3bxOcLp2lpar41Sn+OQOafVi2gW9s1yji9O+tu7BYqBl5k9bcnOdLZ9W+zVIfVI0serzhn6nk8V6
KO+z6a1MCbyiN05cCJr66Birlt1deFSXkCCJG+i8dn2UcDjZiDAUsWA2tI7u1sZWmAEsRJhwov4Y
ePAcjlG2odvOZqDKPpBbAyoHjh9hhlOLx+svF3K93opAKrgmT9PGP9SmmZmu1Vxhh4fdlR9Q/Sgl
X5Sp6M77hDc+pZPWrgGJzuRk9dvG04I8iHFiJOeLBprQAajJ2q0/PWxtnTwzG8b6Xw1SgMqSJVdF
agRcZHArwMnNEVPN8G4RB9MMwRB0OYlaMVuU6JfRz3wX3ZYvoCJPOGgwnPAzLLroFR3Hf0EVsqPW
R81AEbpr3oMwY6j9rjwUmmx03NjeL1XwjanM8Y+h+ps5NEdPeENCvkue0jSerf6tU76/So0KkdH/
mCEjWffJ0435hJb9wToEkuXx4s6YsfQN2Ikf+XbGeZ5XDJa4zzt0yR+biC45E5z0GVPcMougXf44
qcEx9nXdgVGGNWnRupC3iLeF694zlL9NWPml32Q/K+SD9pUOI7GwqC6EMV2SG7f9i32eD5rLPfK0
E/0p8Tpmf+Utm8AoR1Xkzvsc7QB2W6xeWI7IcW7C3qO3YrDyc2dmmXSFSJIgidF196yBHrHE1Rp4
elCPqkhjx+VOk8w4jH9oyFAtypFrgmN8381z7DcK/b9/N1BINWQefh4zSrIbOD/UFRL3XBh36bkb
yredX/LLJK+KyDFhX8+HttOcbI8O58DxNsKCAMsBJpvoyU8dpjzpcUQjsgh0Csm4EVALu0NVPnV3
to62mbwOGpUx0vPjwQNBNvNcwxHJD1eI6A94Aama2oDoz0DGbB6cjqzvqrYPb9RIWSoEPhCJMT8x
cLLA/suMF6Pd96sYizmTOoKXFlfi2AWabOIxwOV9OQTfBFbBRRZ2HjUmPIUwHe3fUUnxDTATLzF5
gCUlnPMlyESANjyWU2jgmz1eSNG41dvaQhnlhkRF+pGxIJs18cTYTN0kabE9o8RgdfLVGnpWTQXD
Xs5pYaexJLY4pHcVw4CSaH2eSSYMAQBsi8n3R3uH1IezkEcKapQvLa/+1K3sj6ur/BFBRfVkwasY
ASg5IbemYbnrhJKHhZOJvBvPX0msO42SJUADGgNVeftGBhPC8vVGUaHetsiIURm9W0A/Lg4T0jil
sdWpABEmEm3oPjCNYcGe90eqAOOs5gvRL4FwfdFSUskENfhfnwXhSZMqaeWsicFSKyqIj3BPieZH
ICXLVNmRpHa13MM57eMOe4IRj0onY86ArIK0SbYBsI1bUajuLmkYFsLZ6hH2bg78bxiCRb7mvJ7q
bMEb92J+jwqlcgxFGK9L23pKTDg4B3nKwkBmUlPrntPYL207CkJfjQUi0eqkjMuE5VJuoXYtLwmd
tHmITXVKH1t87iFwaPemhg5o2fpupJKZzJb6Zuf7SOMJzNxiCTmU00mvu1AMFsW2gXTtYtPixfSu
d9C33CbAw7p5noMcXRemLIEQEGJBJ8NdMfZsfiDM9rL9BTb1WVbk2VYk5b5InOfyrM5TT3RF5Vu+
wHBt2BPzbXFsAKjqYTgU/kOUgAmGaU4ZNXMo6PC982fzVvKofupnCKI0NfuKcVmhVnfcYuDYyH8k
PjnBtiKA2QDXVX/4NFKo9lcAQdflRSCnpV9ZLR0GqQCJ7lxgRy7lNGhSRH40++DUQMjQvhMQUiLB
Is4VRIstUm2W+FQIXXzvHveEjlpubg/KKGUIjPLUX0uAqz+nj1O6ddyog1WkdtDITd5PdrRYeI9C
H7iVJMCtSH4xJUmMjL3oLK5br7v59qcx5Rpk7KlkPHIewz4mHYr4uwPJ/7DREvkGN/aTi9m4g9r6
mCb6ErRfAa3WEEcLeGF5vvaTNkkUtpNpz1EVTTBz10YIUJ6f8SMQYiYrqWDZLOn7Y3QssMdWaNOV
06B8QlBHFu9ognXA/doib895gGdDiU0YsCkSSnTKb4pFQ2o91OFLXjxhj5SOq884gd3H/4q8vOnA
hLry/EWNuA9d6pESvmlTrzXvVTE/sbWAeX/HY4NmagyYm5HluuYCJjANTEkboGXkwuzow2Qotlgk
uGpr/ACY0xiJTMdmW+WzWT79ujRkqnV83ZpkMbAMu5zdDibKnzihDuxLSqnA6Q6eLafD/f23zInG
+zc0zaOBkvqR7LJj8t4yra+HHlZGlEDwghbj3HkePDZ0WCrV9q+c9txITyHn6okaRFNDClXL/X/k
MxnMxg1UQkQCx3WdrUUMg2GAk8j6V8aPfw4M2xlp6Ae3KFfaIgK4TWZvBcGRDXDnunQDj/+URYoi
DYnfqG7yhI4T0UNBwLO9i/K8wGSyHepFQJwLRFbE4sqtyDV0UphJp1IszVBjyH6J6TVo+yddHUfr
bu1U2x5Pf2E7jb/VMTBtnL33KSQ9Q2QbtMiwJ3OWG86ECl7HvRN6yPMGGYo59PmO4jjCBguE7Fa/
pE2iPLwa11rXU+rAGs7O2sCePLjRib20umkNuo2cgx+yGTzX0smnogR6JYd/mTxe3iwlmxsyQ2Rg
ekrkL7nW9BEujscL/scLbEtSbj3q04Gvhcg6FzYdwXc2xbbjgIMnI0X4XXFmhfjdhdw8DXXcMMv1
FI3jwTeCfso9puAeyQEciVAf1Rt+pV85V30XrPKE6lXdYbyNpzvjSYv7jTComVIi4vJ5+PxDJc2j
2C3UaQESov4K0UWym/F0UdLnTM7O9aU/VI4GY2iHmSuzdp44flH1JsGLLEk18VxFqcpYWoMep3Bk
psGchhbUJ27z0nXok4B7iVM0J1wqPoCq4nVZaMrJaSUs1j8B1Eyu+qLu5AJu7gYRd3lbYhZUWYMr
8c41TqK66zru0tby0e9FNiOnpuqWwpnjpno4Zb931OOc35JN81saqnwJL3JouAs1aADsS5D8l+WU
Mxq0PmbyvdqTtjwJkqqdn4wwTccIPnnrFbxmZoY6zo9uYI+zMLT+cZl9AJTSv5yuEwgjELbT+Kvg
5l0Gc9B4bUNBWVuBy4SxUE4ad3c/sw2FQxyC8rZCS9A1sJnFadXiyY4zVMSUeCjKrJx8HGtYBBgH
gdBeet4hvL8ShaV1LBVDdTD8TY9JV1WCrr3scqsfdNZ2ZKseDYrDFSP/Cb+7sbNVTUb+LaIYBifT
VJ92mgAzc26lSzaefYP35Jg3feruBluNi5BAb/Y7sySAE/x2Y7WdRrM6pWurdOq9+Eia5eUv1Wbc
EwdYThFA6RcKi2RJcSLhjGBZPw59cjvFLDYTTGxGFFPwqXfszlmQE9jTggYdzTEcdKPvk1410CFl
jCJuXWe2FVLD5GSlAb+kyhC4yUmy1zACvkCBvjH2SsDgVndHNOo/oo9WMrCN4ZT9fVS/W5Polbr3
sgex6xVlSkj9I40uGgInV9gLf7v0re319/pTEidDkfrFMNQQdyg4lFyUv3oR3GGZRhFVVADkFCI/
VwBWgOxQLDV86rkZXHCcgfP7PLkctLp96Ma6nb9kvrN6B9jXCZj2KM3IemzCN/BJWzqF39p/QVJs
qS07rtWxUPTyw2zA/SlFKJhmp6NQpceBeDOyxv8mYq7+O0juR98x9T8Geeozs1k5HkuKmL06JfFI
b/4nPQw8g2y3Hr+Gc3M+YwZ08cEIauFK95zvQwGbXyfdEdcVhHm8hm/IYpjqhoNoofycEwN5EH5e
hXfMEqb3VGDr13yRh4tCBbUO1d8itQwLScR3YEg9v2ztBEiFZnUZJwdWNVDJ1eQFUUkdgvlw6GB8
YHRL7LMeNWQmwgjic75yMiD6U27ImM6Fd07aBUe4dt+bzzOH4L+qgZjQxeaKu5LR2t78ll4Xr31/
T5rm6UyRtWp+DKj/plCnKdjny7UWbds+OAA/P1sLUcOmokHUlHW1GwG3r+u4skipDkhTADHvTPHQ
YfgLX9zY5nPA2p02PcYn7O6qZLi99trvaqYjsT+ETGM6YSGzJ79UKwCGW6b7LPhfFEGhsBMCkOsw
1HjXl/xaYGd6HsHgEJMAfQPq86VDe6pgBtXE3oUz7/UzwTTzJS9wtcBpJNqMbnVsUTKhnjbVqo4i
dh6ahRHla6lWTnt8AZz0a/PlyjQVvigmnXSSuLKZq2puJWKBXFl6CKzLJeAJ2ol+tAGio0MPIs1E
JmLSBUMGnY3RCMf0ysJdABFNKsIt5rCbsig1JSo6UEqr2HKOsFbM/ZP/zOcHkbQjJmqmLDS/Pcdn
tjn+DbUn8cwA/KFGXyeOAd4iUNLdszo+s+c633MMluFZOcDN/MlbIAL7RrDFmJVtMra7oTC5bEsb
ZaB+NT+vFMw6I+WIU4Qqge8jBDh8zxVMhNKkBKY5uPeh4l3bZYlbjwnTg7J84A96Cv94pj+oSnHA
sEYpLjhFKff+MGZrWVlx9nBkm0YwAEKo0WmIWH3qLucSLPMc1bXL/NZoBLSa3UVI76vEbinPHshB
2M/tDsv24VPYadek1dKV9ILRoKN7zBWxKhLiGoW1fMg/izpVfgdRjzYSA1w9buwdVCy9EPu9UZ9G
cj8YzFukxRHG8gBlPS2ZCZx5rbn1SbBKw01ej29dAk8N31EjPRIAso+mh2mVCXztWcDN5UWWuBMW
inebLyu5nilZwGHba4fXltQq8kQxKOzRw3QbnVxdIY4Q7Bb55lcftabp8dyA8bpruEq4PZ1LcJiL
cdq+Z/ahNs+fXXzUIlAAXasHqgAPBXgUHXnOlisimRwhb1gHXcEY9miwqSHNn7oX4enxhMNzdlcG
XEavf2OFl2MGbl+HaKV/XEIa1hql1oepFyhOsp+sk6XAsHJG3KqZXDkmaTZXNy0klOxuKdJDlWw3
NajvwHXyqlwehPAmotjIVWeQAnJxDFXqVITOjORgBQKMZvL8WGqwCKrcZtmizzXphFHifmUz0g8Q
EVnNEhXDv4aF9eWtgfx6raxWv5RI4YPPps08ke62sVDpm+mRzaUIvgl0+IJKZjS4HvTfl1QyXYpp
RAkS4QCTZkwS6zOTL62LMm3RvXh+l+elMuP2yrBBTClPuuvSPoAGFmxjg78Y3SliLwr6GxjYPpds
pVyfhs1ShlzOhzNexA0VsHOXMB+46ODUe2VASQ4gNQ6lIAoSLQSZqHZR11/KvQBHsk2i3ePxxohq
j/HQy5S+KdOyo6C4NPj8AX/SPBlzoewj8v0qxlulzT4wm9VCjmY13iXVuE+4WMeO6b+t39HG3xT6
Yt9Kj5fsid6r7oI4CDn4/dBOddbNScHge0xI0yJba73rJffUBTV9RtUEjrs8pcVL+QnLKf+cnMoJ
VmD74UhyuS+k2McM+/jjDMw+v1DDqbyufSoYAemVFBXD+DhCUEFLB42r+CV5bCSaf9Oa0F5wKvDk
sBreGmVPH3ggC+6e2gge7XYVYHZXxKHMwiii4oA9XyaYrriHXM1B7LVbCORqLirYhwJp3zRGHDgW
1kN6rxoJSpjtq/D6Fos4Mlc3SNev++eLzIOV/OAM3VUs2uLZEqmcuMD+V4p37aLd+AzeibqDw4vQ
ZKOMV6rosD07lKzHGprGza1MwsIcXx6W3gnMNXEbvgdWcyP/FUHGZrTwvlT2PnR+fbrzHJ0rfcfd
N21eeC5chk3bo7QCilrV8N2W38YzuPidmhR5BUmvjs4lSzN4hu1NvaQjiApeKn1unpPkNC22gyWW
9xX/AXeGwnZEz4FuPG2Gt4LbIKg1hnztGlbm1NcnP5oPK5WBNrOMRQ7nn1HthtV5q5N94i/P9m1n
clhHEwoZpD/qwipnhT6wNo1xnknTARGNKsUbgx0P8Rk/uMxhwQcKFIQST91wTs2PBUxUquK4SRoW
S7YSHxG6XuRTogB7q55xb61Ecp3v1XWiUI1NlPB3seXvaeCiZoQIagqfDCMIGbBlQwXSOwbyeoU0
qlqlNGlgTHbwC9WCigTuAPdgs35E1cVGNwaWMRfhkN45Il2/Y2aXdgOaCYVLH6CCIFt1Fy0GXvd+
UWnazNB16Jf+SeI1622GN3pdRY7PSmmL+Bd92cmEPP9ki0KZgkvjpQ2jiAisB/ovu6IZJKukQ+kE
cAzQEjkBf38+KgVY+E4c6KbLFFoDdcGAV2duwITAV5lDT6qUSXC1G7F+IWhPuY/Tr9iG2pqTxuo7
jg/V5nQffzMmo/dRb3zxa+XwOD/iGmZGkrTIo8KhtC0uMMvgFcDACxrZ3Fc7pfmyn6lqlKMEy6CB
Di1SqDQq4N9xHSeqU/D6SxIW+PVhepfM00xsEfSzc470rnCulAiBT83Nhr6YU0GMi5Td3t3Uomfx
iDGWd10YjPTIbjsS6h8GwnaNB7FZ0xlO6KFyOwFa4nxfQNRj4BymHfW6sqaCC1+PR5PlGlXX58Tn
8sVVUm2Rlmw2mJ+fJzuwhw2piF5PpPBxlkIv77DJEWuf5WXRIBS4nFIZVIsp7r3DKv7Czjmq7S5u
u3WqRgfyRdUCkBD8J6o/3mntFVBBCuHthwsCW0CThQ644YgN9DuRSbVRV8bC1ssPu1GanFYvjUC8
Ekwpy7Jah6h4wcUDPGEc2WBB5jvWcyHNlblTjyXWlEfQj6NLTOXVmoGRWMMJodhICMapTfwm/m2A
I6lHk6yWsuzTGSATICqnSBnbi1Fw71hDqSMDMnDXQLowvxOZQvToDc1djP29UC508CxZh1IHzLC2
/Y7YFFiXc66rFAG+tnidCHBA3fgq0tCf4zQA7VHg7SE6GiR5drmdKn7dg9vokBixeMUHhOlLxecZ
W1SVkbK/0nkXIJ+glMlxLfVMetDaEJMUbBnJ5SE9EwvdnS8ONXZ52cuppSupkIqq747T15XDeAW6
HkA9luMSY1l3iiN5hCrsT6MmLA5AzmzoVfFvDgbnpHJLjWIopxnV1DHngPuPaUGlyfoHq/bZHOYT
YsICfBZF9gWYyjvhitZnk0ep0xQsrF7s1xyV7AqjnXxGGQUnaMhpoFlZalwMeK5m4URIeQFa+OG7
lW9LLL4qW+N9q2n0b2VQdHaItARFiw0uqO0w4ULCQbSrbmvqlfV56KDHTpq64c3pVOuyNgvJwY3Y
tWoa/MrlbcI8UoJBXYJORMSFCfJEiBUWKK1haIi2Ap/fFR0Uq4nL0JXxPnxd8Xx35i3Ocbd6twHD
BWVZQ/qQ/NVPhjpyYmW6j6/sVl8TtM6ZSKU5uAOz4VlBcqrZh/lrQwgRISBxW6TGRte1SPqUJ8De
B2tKYprdYCCUWenfj3zrS2wmRXy+xx03gqF96Agb79mRlY9U3kzriu6cKxVyD+b+5ZO2RXLY5DNl
uYZKJ/xMWF+6coI/x1oUTfzPlnKxC7I9Xhqr1X3r1/kJfsoMO3YU/0PzVoIopeNQWgg7NVOm8qVR
ndH1V2nYPDwNI57c58DZ4kJL5iptbH4PppV8PolJGDVZc4gJks9WepFZvlRg09yl/Wctn6T2CDvc
a+J0+g4bP5k9vNqzhWTAAhEVfA4GwfTDTP3rN+ii9kWSoj9CvqhZ2wsqo6LLrUOClZoQx8fYviUs
0fzY3tIMkTjeCLFb0cHP4i8cP9HYita3d7yVE+En3tiWGsr1Qf1v7jCOUIn7xa9hoIQFOB4wd+Wh
MIGSznUh8Q79GuYJK5AW5LQ74r0zkeoJ30KRTYoM42myJYyxpO66CpWLHARKqzMoOrNeJGsQpmTj
GP+k3ttbVk/vBGY5eSMaKLHO+ScqbeRlz0oA6jRYCoXwFHSLC5hnRaAenYC/3PnHFxAQPCIgmb5B
BsRS0kDY9bur4qvjdwE8TwxkUS0MCHT2YiNNpJGpvqU8kmjZ41D3DH3Hk8RLj54aHwTQPQVKsvvo
vEO3XSh1D3QtV97cu1abgVStLpBu0HglwjwO0sT6JIQ/NbNBzVAFl+kNrkl3M5JNR3lP8VGe4FW1
WV4DzqVrxNr1Nje/fbTYA16DWHF6pkZBwjZ73R7yrHpXTWoU1R6sk1C+sMPk5NgD7v0HnUWM2Bwb
h1jjQZmwRs2MDAysICe7MeZMmkFOI1HujEM70eVLkNOnsI8CD5IN06fNTRdLYJ62xtgvmstls4Hh
0QxIKF83NnhZPbkSrC1Acl6FI6PO1iGY+jmP5rfWaKrmyDn2ofd76qi5x/ZlMtCf0GnJF78rTPd/
P/eqb2VwSTUrW5azicLvJKl/v/AaZyYf2b1dOsG+WzPGqCIPP39u+YuwdhptMSSNocKdW/29w94y
kLEBDaAvY0ncAV9+ClAjta8f44Q/rHRdDHODTkj9MB8QyIX2FOcvhuOlOCntTEbzFlhg8QpRa9yH
JNT+wetWZJnEkfvWgSy52Y2tHicAMAyK9CU+ctdcRjiisSQ7TSEXZxOS/HIZY8+5Umnk60wZBVWv
q3vltQh0vVMupYYlXWtVph2eO5sY10rlCDkxeBNm/nt+xEVf7PTYhZm8XPdlvgJn5zec9Jae6w8r
xj8VfOgRQciaQBrhUEwFVbAsBofMMZ023GHzF625vJIdwtW+fZUHxl4gA/FVbln8+uV/Lj64URPU
m/qlkvnZqXVsJIbQouyuCrLezJfOD3dSoEWqeWs+dE6/PSPubAvaUGZgU6ouEuuMFrgE+t00XoJC
V1UHNCPWaNA6/b2iq3OrY/4CJxr0qvfsI3oWyuGqbw9ce2q/rlhLdwj9yvhDXppBDbae8dU6ATio
auJYmdBYf8Kh7ReJlR73MI5dp451+C1JwdW0wtfPjIHc0tfj02HJg99h1xe2yWIk5r8c4rD6DAkI
KvljXNNdx4XWCYJ2OmWApwj2x8I8Y5M1NIHBRXIAEcC8kVDKN8O5IdEtPG6RjWiZb26Z/YRj0gQ8
lLLaqbueGcl+Lh9DqREV8W0Vur6LVoIKJzI2eiTUhsRTnksh6vQj5aAMUCGPcMr6tf2p4hWOASyQ
MhKv0FERl0+D6wnrPR8ObEnhoDLsIMPi/n7CUCm6cCAagucK1yLaFVrjoRvagiM4+Ce6ibPz3+Ul
eVoXu9566OGT9Gd8toNZD02poS671yg8IxIys3EXHKO6/5mr7JK3G3J/JfYEAGs5zQO8CvRSEUs8
kTqW7wwm7TSdZd5M+ZG/l1XmX6/jLDwvnkWU/rGAtXJreT1B/ajZNjjQsDfeFFqMAq6Chx9eQScs
Mw1Qne7Vh9Fh4HoTWz0vJMQCvuBq3h2FQV/y7QMuLFTqXwgPpFNYwybpr9i1Xogz6DRAvGppIRUE
+drMTvdUSeh50CGlq8L0lLgHvoE7I9LTmuWtJmqe4MLF47+hn3Qjryi/qmWiX5bJXy9KRtNMdq2d
OUY9gdZvYS7fvRR2VLNdwq1+frNnJrJMtcTgOrX/Kqs0GRb+ZFbO791lnOcmp92EZOrwFB/iHXRP
RUZ66CPCwQBWuXgvnIQLRTll9T14yuNBFhqfv1rwf8ZXF73ajAr0PiMDLCB0R3mNVm1dpcmwvBb2
g4Yw4Z+6mGan5wMiCvF4O5Bs5uNU8Fz+d3RZ7MdXF2CWo+JSuqkVs0cmCA9lsY1cb1X2KHeKH8ii
yh9wQv18yzVao7Zx0NS9UEMezKZmJay7ARj6JJUdFVCmNglXDs37DzmU4bsvmBvJK7hWM0xNsGeW
DOXiDkvvzyH2eMuhieYYjeC16DJChqHHMdlpXFROAgheoikSllcCb2Tp8PBCAlPy0huJ/BeoB9Az
QGzQVx5jbg2MV76G6sg+UDpApSGm+5vLqQPj6l5XjAd+PQiFKk1bTjgvGNIbnhuX5F7lZa0eUvpM
RYtyO62UUumCHP2Vq4j44oNoy1ZUdpdBlNhQ5wApVsTb6Bo2nMuZ+xcW6PX04931mufBEAlnd6MN
6L5qv8qY3++OYFmPByAe7m4t5rA/kpyTcf+AM0343BPyEhkom4LXeOPrGfkZYm06hL6cFZ04pnzv
5H1JaG7mte+28vS980wNBZxk/wM1BUoZII1+hN+MZwG0Zh33bgm83rHDr9qpX2fP/qzHD6ZOMvwq
8eF0/CmZAGby3NtTo1ry4X16Q1uue91t/Yc99OdwvgGLKFhoGJtED1wZow8ID0b5sHXsev+V0YGc
GrqmNeXqkjxyYhf8/t+PP8GTYeBUfw55QwrDwE3YMRnZ/X+kmc8E7grqzk05yJMK+kujMgJ6c0uf
fAgqS24Lngi8oTmT0DWD+K/4KsjmHmLOhZyDIVOqSlNA4GZLVSU1H2K7aEvgmQF9W4SdKTPztPAy
mxOjUJn+sKc1WdP5JNWRW+/UQn/c9VPEoJknjQeVJjkbOvOzCsRby9N0Gc6NHXVc+/gvBLzVMmPX
1xxCEc7oW/0xjeOhCcA1BQ1VUrd62lxhaqCwkU14gbMnMEO4jMdBgPZFCsYZ9gVUD6qFe262NLFf
aYvRywtcIA+lY+/auSP4XNHBd5dp1M3fr8DBRky5H+kHk1SkZgkqsvMSIP2CRBIK2ePqCGngQNTI
Tal73UszQurqDOvBZIGhr+OSIMzNJu+CHZYrsyOHazUssnPleTmWZwioTQHbAP8f7NDyqt1KA63V
J+Q/STgIsY3dI7krSOXYwtv+fbjdfEY/qn0cYmfz2KSifsqu2zNvGozYWCX76opDkfc4gNAMkDEO
Wv2TSIFHeJPAFX/g8AQivApwzhFp2vj3XewzW6fgGfZ3/wMZY7CdZN+m1EDl/sVpTMG1atnvqun+
mdCvuZKhwtAcNXGNwraaYKr7v9KZODA3jP0BZZR1xPJ5NHUKNnbIzI0Ng9+iu9XR31MeOUkjebeV
e1AnV7F4Yfz1MxSAcrVowPsrbv1acIi3KxTRfRhmxlBiZZkWSFsSkNNyqTdM1aH0izb3Z+ipjEdF
/el2hy2uwrVQm2y1m7JQB60D684+eOfyRrlN1FTEGlYy7zPlHO4lz2EW2Hqbv/BaX1+ENuCjv85b
MJtfi1JJTdjPPkbYSEknMr5k9OSy+ipV/gQZ7aFEKnaMWbRoxza4RRaa0EqljhXW/ovQKQ1xsiso
uuRVX233D9AfgF0ml2CW7EZlNLn5CNz+34/jH1gBACdPgAFFGbSyhZqMvLxROxoYjkFOiKMPicPL
Uuq5yH0rB63N3pMjnS2m4Oi7ezE0RGCgkyRnon/w6FN/hL2ljb8+3wwJgL7OhBxToh51W+lnG66d
ZAapKVs2xlzoDkFeuonpRdlU1fXH1VXdHFYfEklolT1bP8vwoLkivZWZqb2gr9HuXa+wumrb1Zma
mEeaw8bPXa+BK+Xxhv8Tj4yNTab4O60uAHlVaMwqishwj812VHVH0PmQdWbI8NjtgK9ru9zAuyV1
Hn1Gw1iKEXlgJUm7xXyjtGfAcxcGEFRNtkB9RCKqEJ9jEsLeBZ8BYAEXtaWOMcN4/nBkmUb9mP93
0LjcZb8HHf1GcQzuamTnY5hPSz0iCnfIfRh9XY/zCOOe4M4UW2Q5O0H6YiBoFZkvbTnIgV0dqcrx
Kjpn4OXMzlOrNU5v4Mr8XnpqWJlW0P7u4FXXRHS883HP6weqm3ZJD3PMv+dAvMQh9jzeIMW+DAxG
9ZlHzggqTIR34U91l5sN0TQt1h2zO5I5thrNLTRzNLbQt4hsfAqgy3d71Pm4EfQx/AHX+OJzaFKw
gbCxrm7qnLLDDaIs+akaE5Ux6suqiFouVSYWp602LPy9e7I+MKCUN4Up5I0njAah8wPv+2CDjMHO
upgTIbTw5ls26BGPP9kYxRQPUJeLA9YoxD7lQihybzPEXpeKWqxzazYDKi7nyyjMel2GgznpcQA2
5XquSWr5dylAyL6FklZOn1OIpvz6XiLcS/RfsEq91t6U8jMZNOF3F7o5tSvMm3NckW2wj7g1QkMi
6AylGzULR4JNKHrgMcH+uRMupDCafNmY2fFA7uwUzBbGtiRcLKFzkbF3psl9xEpLsPpTFg/BUSC6
n/MSWdvdMXYCPu9jFv+tQS6lE46vRg9fLC0VzIkdOhBibJabyWQBaBPjsNl6uKdNfM1LEnMsubf6
Va8QV6PhRx86Jpv4dbtys2YS8rabwMlru3D0jEXpJMe8GqBcTNU7DmE8mi7kOMgbS6UdzLU7maEA
RB7P7SdbqfSAaTtDtQYRnQxI3jov9iutdByZ8C4vQfmijxiyBCAtMflC1mnJJZi2vCqyspzdbZsd
JpK3N6B/qJ7mlcPvHKj3m8Dd8NetppMr6pVEMdOU6WLSzqAc4E3YhzBThdXxqitNT/PMBbl4zIpq
3FizKIXD2jcmVsPcxv1qWoo5C4Z+L5RWUE4BkfbisxdZEZhY2K/e0RAsPQ2JLlLnFzYYUDUd/rAc
6y3FTpVs701eBdkcinmDbEE1ubBFWzx0I866lVxQ56QRCVi0aiT7gvo5JOocIC9ARK/99dZT+jdi
tizzZyJLYS/lRs6E2PzPgrLChtMFqsEP8Qynq/qaoAcIicaSAntjkVF0qdTjEg452AF0GhwOW6+U
oHE1geqVeddhsx1sN8sEgzalb/zZVR2RoV6UskImAwekMqfCsM393M6aiq5TTSKz0JLSq6fwDe4m
jHlbEG57IBF+x9m0nv167ql7MqIzIiYMfwyp0uGW+Af5T/1eI4/MFKdMoZ9hZDh/AM9ZhTyBijYB
mvG+of/d06lpgic/Nb3rmIIQWS2VclyHUGltvtL+fD5YKGC8ycExr/Sn3TmDxUUZsNvndULPoV30
avUtduqrYMs7fdhPq/Hyre3Fs7tFsyJKz/IN/kU0+eGxz50y+l2OjiyxG19N2p+UQPuU+sewlFxo
1/Q+zMgLFwWTdYTPpn9gLazMbQLwab+scKL5jBqexbaIOw9aGhHO2yH8ROKIRV4ehNJ3hzPG36Sm
i5mYeBkq5OROFiOc5w660oFjrSKbzNz3h6QPFc/jSJqygIZzOqGhHmr3pxE3Q0939oo8ZSjvOwiq
Zt/d/RKmOIsQ+ybHu2bEUQYCkUk5FNYXMaObCOqlM48+nzznXQ+jpPfTFoi+Sn4O95tvbuIPaf+B
gLGHlqVTdPSwsiIV3XVlEZNwXV56k7Fe/M6IDtg/JhLHUad3qtHiWnmEUH4ZDI523BIR55xP6XoZ
7Oyx0cS30y8A3esIGvZHPGctaTS1W26Gad1vxZblL1EzxHCWhlKxtBQ3yKNzrlO9HISKn/8zf1CJ
CWBigoa/+b1+y/5jbmgaCOtq+h6yetwOQa9a5nMZ9PWgzU3BQ6R8s5cdcJvtwyOyP/Akuan13jyi
q5AlGCFXD2ovKK2V6H+XaUsnANWX9O9KoFI9u3vzV3QQNyHq/FIVVfBZ/nNC7MPN+hrt2uvmyjci
j2unmn9GAK3D+cjJQgPkGJY70lQtN0rgskuyZ+M8HDpT9FYQJ+dOLgdDaSqQ27NMXjDL76dUYmgO
F4SsX/Dl4nLiD0/MNekXnTyFO372nXZC1YJH/4dsnN/naBq6AoIUJASOTLEYXsV3xQv5HAHfIboD
CCL0Ie0yd24DQDT8G+KfodfTQSL9WnZVOLc7f8kzofu4xKir20R+kPs8Bh85z45Mw8V28Crz9clm
3H7SMOVz5fFP92lka7f/JhFw8c+4QpItka2WVvR6JP0Hj7h85MXzmOkA6idhDO0m8UCHNwConwaE
PFpRToqAmwq9nYtqZSE5tWa8uAwKdO2namQjOP15sILvbLiiwHLAfjv3POV3d241/9TIMXnk+e86
fVl27wNb8F0yxjmZmv2UxwPugqt5yT15Han1y1OzCBhuX//3VXDe+/NE0iqnK8Xoc/+KQ1LHbwkq
KgGyThelXlSpetXcNqY6hlmVlzvLnOxAmeDxh9uoHcDJ3L8W6068ECd/YBUVeQJmszQDjSuybGPw
ND8v7IXUyZs8geeO+NB2dfGCRUmtQF8t7KiOzcV1Y3AwfyaQQurWluSbHF6XF+ORWSxcOHhuSBKC
efbP0wbatX9Y+KhP0oYgBQ0ZKppDb2NIYfwqI+NkmlHvvqdeFgUecEaGU+hUNhDEqQtKeuATSf3o
6cBCYxL+HJVLXY2Fp/k7tGhOtCBDGemk4jwGND0rtEwTFRHBDXXHv+mnpP2PUYqEIBE0LgpCObRj
ATi3j7KeMxYgcTWdwFRXlIUdUSwuV1z14BDnhKe5jPWarlyIGnY3UNJEvZP+HzdDhk8UEOy5bPC6
M7wbw3FQhQImEPYGJ6kS35tN6TD6CvgAya9Cyo+5mAmVkanjSlXul9HBAngMk3XDUpzFfi86cWiK
17ECyYDtvgOpgBLWo3CPmhfq0MdkgVg/PKBXt6bxsOAkIYWjskTWeB0uXE9T7JqGjwAQlGkRtwcx
8M7Nq0Lt6xCfvkuSGs5uxk5Xx7cltaDnu+Rxt9qFpo08POwan8FnvismP2AJyiadLChpK9lo8urt
OZAl1TJpbnje+cQ5mjfi/aCU2pYGnbnd6naUEDgx0hc5E79kI/c4F9FJ9/+oA/oDz+Oprou4ql3w
PL2GzbGCPaZSXiKhLX/9HHXKPeadqOpX+JTJZMcDmgUxoxX+4UiNbaIOvZbg0jk/XtvQAyPm0bV3
SnKfaLJjxR+WnwbJIWJbk7IGHNMhk4nH402qkZyVg88NE0QSmCJ5JjEWIn0gyhH+lPtcyEcmDteJ
EGwE85MMb0jJGFnuL4CIK84wnwKO9F8xyNKZix+go0NK+xnvK8FJgr4e5FmipnqS+K5LpMAlojDr
sklydz8kqR3w/xsNKIuFHLl6qb2KM45Hp/uxJL1RLFwI0QQl0iIXjpFODCXUVzxq4Ib5pl8BD7rt
y/I+mOXvXiTkHA2TDgg7xfEYa2auVp0wpYJVtzSlVy598uH6aFRSY+MA81uAIDItrmyOsjVMc4Br
w6+JL/X/wJWqQnMIfbvf4K72l4nltKGmY6xW02xi+wbHtzEQCI7TlsY6vCLwZMCn/9PsqK7DXjj0
7i+qqCLZGPQiU6uyhZtrELe4XZvc+96wnAuoIZcDwQ8BIpkbQ166kSbwF/yNGoM/6mBE/R6WTZLf
ewxLMoYT8pVpAT1Ix25hshpl4fXqYfM7SlbOzRcJ/mSI2+KnmRtkCQQobvBkSeJXF7kOAJxRVKLa
QIQmi10LLmjeAc3pWgittpWKWd72Dn6XMqn91REJFLoK52XtW4PtqjxN1lWldCIZJtD4BXC7sTE0
RxIBAPtB4VSnRxIk5LljKoIvFQRqPfqxFF1KZkp89bSV/vKxwtraJnan05TDfdE/1XPcwleVE+Bb
bzCx7Le19/Ell/u87KHS67BSIkgm/PFhzi3E/ksgrx68Fq8L4ijech/jbZNl1D24QSqqaHiWJWbc
l3QXEtbR/hu37a3NBjC/koxRL1yXvzfp/jAJEytGuh3EOsBZBtXaBfP/c/6TeJd74XgTsg/vEbOn
vTVDuWMun1cfd9fWS0b7kzZwQMzRtIKYQz0yS/m3cj2jBGcgwdbUAwtC95P+mCr0GjYfRJPW94T4
Sy/b+0KtcXLhJyYkxY+lBC7WZ12CNdlTDUN2llBQdkjFbJa7xOg9ero2qO7rX/zzgQxTGtdTrj0J
WBrVKlyciDH7WFCypEGULl6LuN2vyp5SLyFsxzJgWn6pW7/580MeRkjVRz6I7tbOrD2jfoH4ldyt
cwVKHoJ+XllvYV3YDrgst4HMFcgYGFunwp9F5e++fiBjaxjZLZuwgFa43ndR0fI5RhNMLXnM7v5u
sz6VVIeaXgJ77SEvZZ3XX4ScZ60jJNeFbcbQmIXSit+IEPQkO9wbsCJk4Zs1aL6QSiCcjG/M+MmE
9j0rSwvDabSP9jHRWWIa9x9xXbbcPCasXXV3sHxcmhf9GuKgvqFkB1chq3EnFhmsbOsGRTK7FKEG
sDKjb7YMj2XZmBOjqK6J+leGQvZz39x5AVItaRVt2vc8T5eDoG4aSKwyw8/nvpDTB92nZsAYcRIB
SFiyak4/H6YkzAHvQOQ+CEu11m791JvvlRggypbrOmKCJ65JeF3nSGA366E2f1y9Z45cTZClj4sh
876FCUnrgUDwDHBmQT2oPUbskzltSNYbSHsYu3Vk5KHVTgR1EgDal7kps6xQYxBTznGbhPVK8s4C
iczCLl6hwT50rSHtcsFyU3qqqjlPPkCfy3cNuq1jzSc68Q2fV9rc9HzjN5uFzT3F36E+pS+UALAE
7/kiixyrj2+RP2q8QfOzmHfzxhggyZvOv3gd3G0tGN2TFNGRIsSou2qJXnuAvHmBrDryy0ztRyaH
PKzAENayShjAICr/Iy89n1i1GTFavcBE35XVxh8qYasHFrP1wolRLjdy+SoA3TfkBbv+Lfu5L1gA
qTrcmNfvqQrqgUTgNWrG6AcIjVwlJjRPTD5deWRkvL3Xrq/XOphOiBDFCUkxyzZ3TCXcRbHPxH4N
Ou+4us4i+J9YYlANM9iPJI0AyDIaN/L8UarJ4/g7Yh5+b0QxKTReh4JSBWQZUK6gyQXQjhJGuEXc
hASuvm1lWWSAV1NyeBsMVeQFMZerqt6qcFZTrP6wV+eDWMx09cgSwO88A5WWCeHBVrA9AsPPdreU
gDesM8JHHasrBuJouS9devGtpEDTG7f5qr6NKTgWRFTE9FENEvUbxAWQ71EK5eDuYr3MnZn9d5tV
B/DwQGbvLAM+SCS4OQ0d/ZJA99N0p1QRY+qVsDbpO4xIz/qi2Rixx5LTiT/P2GCs99qMJ8qQNYjE
P6AxfgmENZUcPvZQq6ItcI3gVBJRoQwoE7eRDrsbiB+iPCzicCi5oXdI3+WQ7cGIDBd4WvaEI/xP
+MecuEwNpYRLynu1ueHSRmgkrBVbPXmg7vC7Ax5fBPGrESw4IQUhhRRdcM3iMjnfFcbo4X7LXeE/
enHlT30TM5ofvahW7mzzDpcg5wegayGlBs9Fpxv7Xi0MiXclsqKjJLoVZiB944dx6YtHvKONkd3T
g/ECyjoBTDZt/nW7aVJEOR3ezb02Dq2RrtlFFzXoJvPji2u/fJkp1PnaJOkqhHl/dVU1mQ5N3o6U
6WA/WmSG2mQCXJjFD6c5BtA15I9/ULEbindKbhyuEdPX3GgqqO2LGy5lCYaca/rjDdSXe+ri5kYc
VbmNYpbjLMW6aRhQPd76w2KDfiwaWd82mi0MH25eTzAKexiL5w7vyH1pY5FG+40L6K4yguSfqnUO
vfMgNUjzuFgm3d04GJkX05czxSL43BK5h8yOBN1pLSJRNmHfiH2+4vo/61x8teFNKK7wDXDJSa8A
4Vzsd5p97RvmsefNnHAi0b5g6EbJ7WiQzsy8gowItgY+d42D+/2Un5uK77bTpQWehv1N0pKDDyTW
jS+RfOgA58shNjqkakz0AwyyZEmmbCAelOdmOmgv0AlwsaLQmjVdbrNPS3hruG7rltvRuAC70ipI
7mSxpRXGbVF96cKlKXfw3Gb6pdgfPIK/tqUpZ8RpgtO/cN2bBqaJmlD0xbJDBonVCOEpDhW/kimN
+QT2vdIYLqHv29oM1p1msGDN/2XBIuvK+qpboGn/9cHKijld2VqHgbfD6Bigcmi3QOIhlvkytA+S
y8cjnrj5rn37yzp0QuGxhlu6UHaRdAQLyYbsaghMsK7NxOXAeU3xW32g0+pqqh1CJkjp7QqYe1yk
GshrmSZQBG0U1VcNgILQiHU2kLfWNhmi1mS1nogDNw50XzhRO0o8FZ4O/lyv2144bg4v1CEiAEPJ
izRff+8mM+ezbMtr2ANaBWoCDV0gikzh0BaaAfG6R6BrYmRRi/IABqx3OtMqzEp+dQUJBpJq0OBJ
SRjLRrqi5hEYl3c+bJvLYUAafNkPhXx4/wGwTlZNJU4rdItfuwjFRDtThJBmAWy3lMfR010oOmE2
FG1t9lnBGBXHs5FpjMznl7tfGlMj+ncqgVgSFqFVfa2Lhk4GkIUqhV58scYBKgh/gdd7+kibOhiE
kdj7MwPJvovY9f6rByqhbcSyu5OlsakD/y/sslD5vY7nnx3OBz9a8ezr9QEG2nHksAVFvLw1/+Fu
yK+5qVknkU4SAKGke7RoJEajrOGS+g8QuAniPWg+ozCysagK3KTwwTMTusatzwCXtKoURYweoBch
c7tBkVRRK6PKZ0UK3koDO/XFUSlfBtB074FgWAFSM6jxDJ0I84GA7YElMCYCG8lOHJCU1xDbECl0
ne/1mXqonirYYgqsJ6i0Xn/iwhqNE+Lk8lBZkMQAnNg1a0sDMUjBU+2Sabt5CbaBW3ibENSkDGFW
zESUtO/MeLwEWliyodbFXO+ipjHvcz5EeaCAQOVB2pxFP3B+yTn0oq6g9YVCc1EMrXqUZKciMgo/
ka7KAFdvmVICM4WadIcbyN0iqPLrlBzxiPlWC6BvscidofefiS6REG/QpFolOyPPyEPu+y4wHKpY
DzhgpQ+Uirxa52+aDuIMcuqcGajdGJifWWDh1LwOKOajl6uVqEMW6QDZw+r8Pgo3v7h8fj25k/wU
Dkh/SqlCysVGAOXgaYr6QG/AiC38XHhNXKgR9Tfk7GT89ZF+n3Gj8nsRXQmPeNpdAWKCrxDNeH1d
aQiqhwNy17UhRPBadfmUS2dFjnufUsJZoNxod0GldrAex5Wpmyv6Wn4IkKOjKVktDPwWe1koIZ1M
KSDl22qJjbThLtNkPJzDLRRxryw9bkgnZznoO4lS6nXGptb8sFMZMGSQ0cPlUUy0OXONb9ViHzcF
kzkZKGkyn1l4weQZciMuTZQ3OV/CCbRUZtNUEZlrxx3tG4UPIkX0/TbQpry4xiZiOEa/A2BsTBaE
pCExPIZjXPUL56Huqyes5qkXJzsZgoA+j/JOm5W0z+3qVTbKKqOY1uLD33gJgxM95G0B9SbuJDuw
zAUHQXFa/bPrxuAMQ0A32zLOdUOmXiKEAYaVmIATdsE9HApi5mnQsPEE3kdPUHHaSuWD+hLXKGva
W1TLidN/GTAjskggr3zqbSH28+XjYFin7C6Mn5+iCYv3td9pGNi4EWn7EI5Ob1plbXNLFNAXQH4u
EhkT4pE2OwXkfSdmPXrOLNpnUwhfqMBktoOAm9qMUKxlK2fLYx5npWJ9HSB6G4miWHn9Xn0m6fPr
EQV5HIrO0Olo7+MABQHhwes7+zUXquIedfZ8yPKvL64M9C5RjKMdWdKMbu9Qi5DW6OfsHLIUvOGj
XzjsZ2Cy9gh50vA3H/5DdkV5yZ2z3gPC9MeBlLqTHnRmxG5XuSx4/aX4Qp3t234BgewZNAmbwWSp
Mbqqj2mjzG4LVaHXns2o+bC/Wx3lLCvlVEPUgscG2kyzgIFXxQdHi+LB5fM+E+b3TWjD8IFqwwTt
NUw/reT38d8aHtBtFkVKkepk76KHv5GQQn4tqy3FAjGBJjSvUXbLFT5eH1LEJkcrG3WkR9yEGmZM
RWc1eBV8DUsXDsUUplW82YoJZ88VrQxd5cU53sl64rg3sEkLIw3P+PYqFOx2RSXqf2LoNZbtKIAA
q9jQ6/GJUYMax9v6nds4Qt+7bDFMkn4J5q52hou4cwZ+SOIF1aEJdNefAcGhUAh/aVFu78aP0RO8
lZxgL46PWz2S0ApIQ/CKniTS7X79xW+XsvNH/f6V++BdVipwhLmDwyFDLkzdmmBKE3eFaYZe9yUh
wlTkgJONq1ID9kJ4m9BYknRb9a/MQ/xipW4uWqNo7XlPRrpDPXzuquoDBXaTsdMWF7yD2tLQ6brs
l41Hahrwo0sOk4MCFIVIwD4SPTaErc5NjXRtsqAafmaQ6VM8zrcdfeH4t7F8+Z9Scsb0HtW4p904
CNxhmcOwLXS6o7YxPZGEfvqrdHJxnNr5hd5SLpAb8opW/4g5CwpTHR+26XpZZD3iLH0UjxgHn6Ua
cRfXtypx42WudD4oVEi7dMwh84+X/HygW7GscheE1SLBYy9Kd3TUygQylKuurFryH1zasdFMQTyC
BI7Ozg0W3OTryJy95r5Nf2/jfs7QUAePWB8lxUOYxzikLb2hRZ+WeRvu51tFiYYBDrHqAUOXNUpS
Ka37Hiz7x9Tq9k6z4BslKCXiNQubgRofY8BGDAF4Y78iG7zNZuWfggsJaHZrdZ9etRxVosxY92wu
Cz8v8UBmFmOPxj9xvRmD0D7+x+ukjuQkyeBnmK7RA0+pcJ/BBRUb5qWpMRlyntU1NhMJ9sh4t49n
x9oZIIfmNL/3PdiQ3xXxSi8g6OoWcoyK6yHrNFqN1B4m3/RYoJAPOE5Wkers5Y/Mt7F+8B57s8ay
KcCYLbIivHqoQAMEF0jL92rY/uAyfJEZtqaWZn/s6jSVxh79RIrsKzMrUHfCZXaJN7BoLTdVlML8
jzk0qkg/X0jd3V6qIfQV3xmBnEXkpmMX7//5NgLE4I2eMG2YeoJLEfmbV+rSCNxPZ8ADuR9vtt7W
TeGUjIX2ib6xyztlQ0fquF4Txi4J1KdNcY7+66T2qWIDXFb/nYQKsCJ7s5ziqrShxozmeZZbKsh7
MHO/NRouEFhSt+jZlD289tsKpd2ol5RR8HhXBx+rIGNRWEa0+eJQZh5Tw1Osf+eGwsXAs68DUUpe
uycIHDKNxyHlqDY61zUYlQAA5GLTIH1a8fBIRe5XKGyD9Gp17jVjS30pHehEUVyZxRXqBAFLYHil
aglzpJJX1qWvVtUhAI18lYBU8qiSoeFoxfpPSbi7UwbBNrE/dM7xIJX1oJWY1IqyGmE0vTJUnzG0
9jqm0qxwwhxhwEYkDhUDc1ZydY37yVPUivUr/9q6FtV2hyf9mox6hxVkgTtpVFYBMW/s2P8cxOn0
nT8YXhz2Sx5nfJ04SnDwONLRkP3tDPK9uHeaslpFmBfOTh/ATRa/gGjyp7HR0r6PoYfRqpfGRnf7
4WHQ078sUQ19jHmydugs9o4xaF4xM2PfMBPxSv9voJcVM4zhEpagLd1GVmz4Dv+gG67nLz9WgHWi
v4dO/4GrS/drPMN+Qw+JwQikycClOhPQCUQOIlzO3vPqZlEqX4khqSfUJ33s3RHhCd15V3Z/bn0F
wJuIxf/s4FB/XRBfmlG0FFzBAfDAAK4Ca5Z5sUOCqg+Wi7UMOSDSYM00c/HVzNFS0y5ZEdP+7p4h
Oz4loRy8kUTR1nZ16ptuWEUSDG3LaWp849tIgkwANZ3z0zQzPylhhpUmJQkHFGQ/DyQTM6zF6xHU
fDEtpUsFJ15ktEdCl/s3IghVyA+DrXWAWcNwhlvGJJDfRSQGOtGJA1A7oyB/+8RsEH/hzcjhmpA2
kb7R89YPmAYLJ3US2dNE0YUqchFsLXeqUNsD+c6qtGFMBNqC4rfXfIUQcmyAvNNZqmJGNM7NDXCr
9KtAaTVXkpI7MqjuepU3UYaUyZIV5+DDrmQd7UGr7pRr5Y2pDzGPFkWQB2G9Bth/UTqVLF7O+8CA
VXFkdkv1IFoPCUCNweGANEcPrBFaNT5dXDFpOQp14/S7dvZgs43Lv1wLq02687oUjGPK+35ZEUmY
5YxBYuHIIaYO7BHcFA5Mo+0Onr3wwsQy7WZ1Csk/RuwEDP77zLJMKeGmoOxFx8FypDrbOso7cAn+
iQIR5vvY3MBcFpcGWmX3XcrX2lpdZm88FOXiFkyXm22gqsAZAGh8NdedEcRnw4cAajT1jkx6DH/g
7A6boysphviGEJlv1CFlxlzrAhJ6fcaN18NErxOhl2cPs16nYy4veu/XvJPNfRRS6/VFylgPTugs
dWpUoUesoOsVyvyToyto8/GTUshqsBabK8jm9GI5n3xOeLNmvSAX8ltBEGHHD/isJAopPOT6d7JL
luQrYs5AfWE8M0FdY+RVqDL66FhKdnBc4P8FuwAsk7bWu3NfqukdKlQ7+FT984GUemEivsWcxN/6
7WeNocp2Vdy2qp0c7FEHIwy8DDcfXejoWHve/EBkAXSOL4ALQEwlOimi9xXWtZWfGSBfvk6/cTxB
KpaujYjwuVsc2hV106+pNmUOgic6oQRYpuxdIOOe9FN6zDXvBNn3UMNz23y3zR77uQvRfn/sUP0A
ZflZ+ICRajfXTtJCBobaKhExaxIMF/NGDp/85PRy3bZKKiPwIU5p2HaOENyMLJu67YIwO9rgaocE
RphNbuMOyZWQ8SFGCPvhkN/jq18uvPEfDVP+NvcaBpu4ULL2kGxLzql0gtFgPaTHkNnvnktIvWXC
CgkJ0K778Xp1yrhgD8dLmoqSqaGLJE3PymfTaF+jb0XN7nw/CT5e7ssM041gbux2OiZl8oka74j2
iOkZ+dZHXu5ft6PnIaheFytTWD4detwjuLsx84myU67Im9QgmxLJVu7GashuT4XFvgWp0o1eYU4O
oMlWy/BWWbHaSk+GXsQT+olsPxN4BowYQQmH0Lt+T8sP4E2S87uJ/XTetn1kznx1yxNwD1zCHhgn
WQFUd8sgfxF7+yTaHNjOlRccqfMRnguiAbEa20Q/Y5Vpmgqyg/9O3vJRFn495MQVMdj7fMHJJF3H
RjbBev8vBEadLyjbY7yUU2c+flX01XjMBn6IvnnCWJ45SiAw6qfbUH6u5ZnUr3bSlKtanIvj7W/8
L8ytDpX/O1jN9tIO2qrRoJqrpFq7QDo5smhMdgKpl8g2hXoEV9PvQQ5OoOWgN7I27QEPHH4nsaTx
22Edqh96VvaiV4FIGeZlhQNDA+sddIVWBK6nSpBQYIrElkGapsSgiM+4ZfqVVxtwKtymRdeS/Z/5
dx1rQcCpnSijuRotYhjTIZKLLrJrbvk9Iu59c62uAhH3TqKtX+OUbYgkaMTK1pmL8rwYjq+PQlmG
Ix0DW4+HR41VDDI0mGRPvgS+y7ky7uKN60nYfXBNY7xfVYaJ0lDEwYBM+SgYSD2uOL5M7lbLuSYs
7nKi52++z71g0qKCGlDxBjRIKKF26I3GMmUP9JkHlIQBU+AflWLoaQHI7Vxw8CF3M0H0Qc31AuHN
T4vE+/e0epDlWoaJpSUnhLO4lkCLbwjOWdHvSumx5yq+KjrK2+P577EB6g8hYPuPzqthqnfkVe1w
09cWGY7Iqt5Ap7+IDNSSAGSg+dB15pjCTAFvLMnUEsvPfuW1ckKV9e/VUipxL1itj47oeCSXuobo
UJyFLGgbZ6Xcot3FmBLJoq6CXucySJkqPwQiRDB1qxTzW7vKh8WmzB2VPnBLfcV9emZpUlZ/907U
BggN0yUr0unf4dvfLm/9Ma4ckkE3Kv73Sc+XvQAH9BGZRhxzB03mYYy1HXbQzAW56RU4RyE4D4KC
EXHN80XtdHyhcs97pCQdGykDGIaLn/9wsCPjBXgO452FnIElTMrgxsxxGo3vz/28D+Op/R8h3zga
BvhdbiPVyOF8SfrS2RWCdY13nfTCZI/crH03g/bwsibaRhjZ7A8HmkCXTh5+Fb+onIP4bzFFQ/Vp
dk3ovqrYlmfFPhy6qkvftO3TlB9jZILdqn5YQO3/9Ze9bf+0MoG5TL+wTOhjfl0EmOImxXmD6Uat
7qRb47epMy53sx2REkgUTlrUhHoXiPEU5q+hp7TB1WWqbp0sG7Oe190Q4KbbEcsHIIj7R2WipRfO
2mN9XwEateNUuCxbr4wVYGMVmXNZFZATP5gppLxZREwJH4MtMvbWwmVntXkKmktlYlklnqbzZayK
Zidrxxoe3aOxu0+8mjrexKXFh9nzqkr8W4aaw8w2qnjCSMJdW+Fe41lgi1JBpYe+1rq9ZUQ0m9eX
EGe+d1QKUE3U9Saj8cTHdrWUtaM1bTBrJx01jd6d+BepghNkptImfADi+eSlTs85HzHYDy7JqQs2
PZpYtXD2DNDXimq/8by0+xgOk20GX2p62eYhsC+JyOvQCGwibD7i5c1IUa+ubpeKKREtedJcQYm6
m2XM+7DGzDBpCsAojXEq+S7luzVueSBqrnJoc5IqDylw/nJitHqLJynD0qcGLXoWCahU8IEAdrQ/
OuvwPMRBHvaW7qPDWoQNCp+W81aj74EM5YJOaS0Y+/XXhwfJTf2IF47Dsk4pamOwxomBheDGAp1p
URBjtJqwD+4qX8T/ed41LBxfby6rSqgzxbDxp7WCHsNAth5SBJZCcuKUCzLstzQSKrRdvPkcN/wE
AXbz+evjf8eY06/PoY2up7tZiR6m8ri1frOafo0epK808biMJftH3ZeLYZB4ycrJlgLy0+LZd6Va
VflVMdZmrUKqc2GwyR5XXsA2jeRvaDRcVAf8zz8JD6ryRWzN2ESUOly+p2RZN21S9/4DB2cyUu4I
+idkKUrGK6/hDXn6j3ZtYmRgvrR54fs4i3PHmC4jB3O5JTBAi4d9HDlwgOnX+QsYP1bq+c1xjbS2
0lfD2vRzTcZSbvIWde4N8Fv0yziZQUp65J9tNWrLC3bM15/ETT7L0aU2/aGzuCRajPa2SFWixNpV
ijeuceLWMWudJluSwo+tm1HO0/59yt0bgXb3j9pd6UdeT4Ii5zOf5XtSOSmiqK7qQ3x1HKPGAbgL
3Jo34zrVJWGPKXwF+x+8Z7nRXr9mpg9euMP7uj2wsjPvsOxjf2p92Z4qrow5sZ/vIdtQx1u0bp03
i8joj4UNYmddkhQtmEOgyLQwdN93LDq5DDSZEhZHBXSvN8UVErIfwsEnQuZPT2VL8qOByE+GqyO1
KjpUFefGEXmCYS9gZsRAqhktPx9oTzdrgmdfz0kuzY0dNUhjjwGx/U0ne1KPGTceei59yiwH2/Uh
EO6TSdm06bEhrPZj0ekkVcGS5H7qrGsIsimCuaQddBHcafiiS8iD6G9aSUtecg1yvR08uI40tSOz
XwZrL4vluLbg0YdEKB/397opsVC55oYLAd3J33xr33saTRwQBfD8YobKoDfVyr3YdNO7ubKXYBLe
VMAfTfe0QeijUpAafpMYgp7lkfA3840s5JLDvTLvglX/Z4DXmGnfNtI/J0IL6Xx40z+wqWqtZIuI
sJw6BkTq1aIKFPT162usm3sWlDFkZlL6et9nruedgfpadfLNT8T0UKTjpTF421mwe/iTj0LcJkhD
zVz+9yH4ehIiuez+jUpnjPj6rBZnRos0JthyJyU6wQ5Y3lbM5nCmsWoLVNApnEaLSKdmnmjlyDs5
JJEishw91ajBZte3k6f7GKrg0xN8iRcwtRtp0qg26A93Q0+Tr9ikZJoO9BMPsnVSz6tzYDsYUc1x
LN6Ga0E5uk0ZcA6WMHvJb1FmVHI7cpmYNH4QLOet/6E1TVJ/l70lcoKokEhhP4QEYQRzkj8etTzW
pElCp8YoGsJOBYPT2CcdO1D1xzb/kxO/9UHp0t+8tzdS2flJYccS7PaZWwHNOlcm+3xVdBt/Dzoo
Cn1NYZCkAPfEd8GHSVbYPKR7NXoo9GVwZyQsPoGvAJH/mOcHgeS2i3sLtiNmxsy9Ke+cDVHRI7U8
YMrJrmWrGQ4hTK6UjKFjezoMUhkk9NIng4LIZ+M0j1O7P3opbGArp0pTxzUAi+zQL/AT5jgW15s0
MQwaL+E4sQOdEDv5nvABbygkbQ4mu+46JHYoQ2R6KVau6i1jvOnb1itbTRiruRafl21BVFvNk4C2
1ZYwBiXiyoU43zrQdZZMAraENY6nN/+fnF7OemmThfQySTmyAKD948sAJRDtNh3/WIGzV+my2xLR
DhoSUZHPjVT2GnfM7/c66VHwGRwYRLn0vnvwmL8qHxY/P/8MiNoLaTo9Xdnrs+dnwCWpGwVIcGM4
gp+wEl1nbu5UooazbO8kNSj8ELPHzBPOcwucKNEG55Iu10Ka9m6cgaUMD3B1T2IiTS3KOufeinBN
/D7y8rmGCH5BxHeJdgW6oAnlYb1KWlbmgfZ9xny2r5/+YrQfw0/WGJQvcS7SKxNqIysi7ylZwT6Q
020C70KX4quAPOtv9m7+JnWsgt/okdQk3uUig/ocoNAWMZ8ANr4DlnpNg4cGRAXz35e7LStl2n4+
kZy1moK2ODr0JK/vzoHmWuB/LHr2G6qGGLI6ryZbP07R09LbcVC355736RgUt+JgWgWLLf4/LQko
y8yaYBPgVmpBTXUQPWP4WJBGQNRTMcxcShkYDWFzUnGhXidNgJvQaa+l4Nsj/6zGf6IZP/c5XXzw
2Q+Qb+0CnFHtwvyhieIjjtGScpkF8OlnxnAboFjyEOigx4CL7tsul7g24l1C2QNGL70SAWz3Ruev
2a2Pubeijoxw4Y3uaKETGLHFFSoKnx6Wi9RjEe9Pkt9+tn6yRHQvgqhM396WVGFYePFtfu4hzlfo
07oC7POXCK3xxttjdF39vV/cX8Bw3YPwcrLlrHqGpHliyCLa5U9TvWwCoZqS954Nqh6695dgCR7c
9d/YJ0VvVqa+uWgLZ8uOxoTkGBhzD+jLEzthtfC6jUWrSGPj4begq61hi3OPY033m1nkuPkZjs6U
CMGdLj0bcUWg5wxlM8lXNw/ubFIEuIqYtKWMfivpYL/7MgZiDiaJcm7LTCq6RYCs0IncZ3fOw/Bq
DvCovbhBhqevc7q+DNDMDs7EOqrPTpXjdB9zWg0S+oIlje4vurp2ZHVDv5zGyA8/9lx0gq2B0CfF
vvFSewHZ6FQ20e56htkd5fdnI9jSUKygpYqL8esfkPvurI8L0DwjNgOo6iNukAhXVQ/78vwewOeV
16iEyjx32/RT6GQfWxujZVazlcBzUrb5FosEtLxQK/Asn7uWF7Pu2uF2rb1FusTN96+sy+attSrh
WmpbkKNQA9DZo9VBxMCIzhQf8VYdhwUGKdDf/syWdmtM/pdDkxW2VR8YJ205zJbqvBB7E4amPcM3
UmVJENLQcyDzV5exl4zjZ2r+CsHM2TUEONcAV83AlVfhTw+z9U2lpH24y2QFHV1kcxyKjTGNF0ew
mtYYLOmdrxY05qdqx4bNop2RKdKUrMwmrmcdBSNTE+51yTV4kujaf9WLs07bDpSNDNT4UGMy/MoG
MdI2ox6aLaOtKDvWJKAIdSIjX2vMiY0UntSw4wtlVJkZPMkF+kBqqiQnv8yI+pdRBvRZw209/JqH
M9Uk/q3g/sn0odYgX8h+7ykNk6zGeG+bzsKBJ7Si66R3hjRYqI8a+v3PH6lonrXk81YHFZMJ7XwI
14GAW++iIBdLqt6qupQQc+KaTIdeKGJ5nDLrEJfzPWCI2Vw0S0lonclgVDGppfjk5AC8dhx/1qgl
5kbWrKIVhNK2oJFzNEKoVSJYP6OnL/R9jWerUMc7gj/Zacj3uqoe/MP0s0VVMITIjUW1BQt+9+rc
Ge4OlaKgpUCxkwvbvXhC1QBhCfiEw7uQvL3SSbGbfJY5YmNqJ9MDsFDMF6tGGnN0+HOMesP/C3OL
wW4PX99y4FYdKklhI92zxCubxuxMi/ZKRDSHWV3DytXwRZSAFFBbiFKR5B8u/PcjWcZJhSrCcibF
ONfFcoFdXPW/Y6kR6uzGgPV7AvUTsvL8DMyJWQ+fb83WIRiw1pWLV5UW/Doi0hRyBIZLt1ex2+22
BDZ49A9ACEvhf46wA6TypyNzLgVdNrzEZkWNmtr0utFtMwa/AMO81oSXbFiaJ/FxUnU8Z6APu/8v
JGf3SRTF5g7vGn3iog65SjXTfKg4mZNw5NZEMtqSMPE1idObA+p06PSxCVU8bj283YrC8j1Fkdo3
5sJXtt8X0j3N2Ie1Ax41ZQCvqeRnsU8flCHldWD3/G2jPn2XPF1NZWCkzcZiWCYiJ3rml8vJbMAN
1ulyW6zzHDNmufMttSRf+Iicq7YLviw3t0Mp+L16dqyhVTanPxC4fuT+Izqd+ww04qM7X/j8Dlof
GzuHyRyykowv6YPrHxEYhiavpJkb92aXodANEUXvqf/DeTleSXDt7NlX9XkIhtghqVHM6k4TiNoJ
XnmC4vvr8zfEersROP/vdW2W8W9ypDtLfYb0Ekpnw1d/eXDbYfKjjEqKbM6WRLfXeow7ga80tK6X
B2qKZZs41OAiDXstdiU8RgYkF7yeFA+Y++PHBRw8zpx/mRH7enggiZnNGBENp+yDRAT4PJzk+std
j5dCU0WuzVR4unMznwl2frJfkItC2LQyeIFLRsaxlLvwnBcKhLvRmKb5eVdJ6wlzye+uqQU6yFeK
zEvb0wnG6ti5e6PtjKYjT6RF8Z15Ujy7xidLj4D3ZtlLQcMrHNtqxZdDZVQ//a3b+5BvfKFBVMLI
QG6soYy5ol7/kRiggmkXD1rowqQ/jNEnM1fp83Np59fmEMpI+7hM3GVOVdS73JeDazQsaopND9Es
F8yg8z5JeUbIwMSwRFqyLJj+kIb3e8SARbZrocw6XQPyzPqFqouviHAWRyej6BBHuURmrz30rzN8
HGYIqtCJmX9enm4TQrctD/x+3G948zykAPTpTusEyah7kRV3HCodQLeXwFfxtvwt+G5HneuvOF/E
aEtBa+rUXA7aOf8W8PXBw+SmP1YYfdVB5AbQYsOyZtNxOKEJ1TEC4kn4f2SzEoga2xYSUWNoncJT
NSIAQzs5tjItZeeqqKwM49zXfk1oZPmkcVq7XLA55+p+Hx/xzn3a51jh3WdYGcgXXgs9TrBorT/Z
hv/GU+Di88aIfwKzmAWsIf2DkW40ktow0c0Xpf5f/UBUJmUxmlyT73rA8NTQ6G4cbpU+nq5SxZ30
KgkN5nHD8u38wT4pGXZFLB7RazwsuxkIugEl/LRbgcQtuSJZUAiInqo9DDWVdgXXCrNko/NMmAkm
qc16jy47IBwEYy5PhDPSn/DTuNVx5fuNIlaVloih4x32XYOFWAORhUIF2BjCIjwMQODEqZu9feMm
+ewelsPHSw5HEtxoI5nD3oCimnnkjzPjFDYklckS6i2nSVBRMEWWfkj8z8tfmuNRbBrbvA+Cfhqh
zYhtpaxJkZdNE9Ah/iWIpNwacaKFjxE7TW31OexXwpcLL8zKBsSIMzhdYsYWQdKe8R7P2th1keRc
UnIPxwmTNlJzze0cYVSRuDHJKlXxNrdpQB3esNsIjo62kf+VX8fJAcH5ji2NrlQOeJOU31krM9j2
SxR7RFJKwdxThhUlfr4z57BDfwoE6pz7uzNSLLGuCP4fadNA49yILkQD8qjNrKhc0v4fNSYheezH
qT6l85lblswTofjdQd7LRM55uGXF2so1munoI0QT/w6YwxBSVCl+ehlNgjZKW2pkPFalcg7jroJV
anVl1jH1yW4W9fQv3QbvQxqVYXz5E3S33cijy3xUgn8d//xFXl40JaU1oDv0MNTbDYMHButeiu9b
1lYyeOkoKBF92Uhwo2+1dsJuV4IJ2yUi+h2IHu1cOXFXvbvDAZOqR+pALRd3RN9JRCMcINV41W23
sfTp/J4E0vZcQOAIVpKOunjiKxYO1oaxUPLdtGckZmOiq0RpC2ckRjiLgef2uwmnk7TFQlGeQIN9
5YodjOG+gjrps/7uuSxBxJnr50rUwnbn0XZUKZYF8ZMVr006sMraH9ZmpsY259RNBc1XObFqUD6f
t1a3Gw0kWc7fjAuWhpy66GjfvdcHqQ8SgW878Olsn2pjaT6wXGRHYTJNEe9Tln0KH+m/mAzhp6uK
5hJvz9CuGz+BOgMGx2C3VV9hYgTyB/VCy0Yjvu0kO5SiJbLo+XOLneCNc1wQ3YL9lJ8qFRFH8Swa
F9h4OUK5rw3sIWm3SuYR+6RwOkkbW7pod1Ryf78z0Mkmup/TH2fGa9VLatPTGSriwLTpWq0WrMkf
O7OH83IPTtFjnhb9cDe47eBaG8pvoKYbY8pTG8rvJ5PGazIQ29rfmkGSkUC5UOJ71kYbwOYaxlcE
QYAXZUvViuMPMcnWvUlm99VYmKYqCatY1eXU40IrQVKM0QI6LhVlOJnWGNhh8/qZ7hyoPJGG4KC1
CZgC37oGPo3FKu5vqBSzZUGKPYziYlQMU0n2a1dPrypRZNrZUUBPS9ZYGAEK8qPrCpATFXrT0E/j
/cjZUkeigh+wZ6qwW9WHNIrvpqu3QxNVO2cz07A60IaaiLd0Q6SCV/bHgcWN3gWYqhDycXfPhVis
22M0s0FtPm6HFhAeBfPwV5to8Q/bEzS9LHQjR1m0LKKGfhygib8vZoB5OzFlVkzpqczkcMeipBSY
W50vc2mGv2Obm7+xMX2+ZNsw43OGCFMtXQ8kiWlN3nYQKVmxaX6BynBiY343Sm/ti/T5RO/1OUdF
ECtybAAOD+3+c8ZEW89/I5IgQWwf2Y2eTb3KHPn42cn3PB7tW3xYR3Ou8iwOQI+SrIzqIXwVLWbt
zN8BuEzpw8r1Xp9bACmgPe7o2T+NzvZFcIZn0Wt3NXyKC+KoZ63xFwUfl4qQph75YD7PLPWjPp9n
DG5Etlcy8Udw4MPc+QT8RRKsRyqhzKBpBe3ppI8gk4gBj5jm/5VeTPz2cPG71hU6puhUbUsXDnoQ
pHkV5xRHnD6XGkBRWgmTpHfticQaW4fIXWZCAKxdCQoVNzyI0IkO8nDxglHB3C/g4zm8JHzi6ugc
v+tLxV3WYWVmvta3zuphRZ2nWzCzf8csA9TMHoc/Vu40YZyuAg6bKaNjZ0aZT1v97rkiQDFDd+Ug
z5sBsspWvaBtfWgbnwhTYdjZP0ovn7DFsTwspdxXEBGIWy3REwSubhCWbjoTlPfx2Otcp+j2BsNA
ek39rb3i+QN8G/OvKFSL1psraQvEgX92f/+Qw3yd9ZW9Pr3k38WvNAIpfoAbRoif/w8m0KgLWTwp
FNXlQmNrEkcFHyRnK/75UlggJd6cxQf1IpbecFUVURfJczmKK3y1htntZHDnd79YGjavIiToTwji
Xl1foqZIYKbT3sE+24QGVabTQQrFFk8foaQ7AJRXmiVDlEFubOig7qqkALFpPlF6S7fgbye1OUpO
2fz+x6qhjYPgSn0Wk8YP6mWKBSmn4j87Eq4cnfBZ1AwWUEmUF3lCERDX0A9PAejYsdqTwNQjEy3n
w+yBrVIF0xxqc43KoVFtUMUHiQJdRbhKfiExto8xGBrIg3NqDo9Oakzf5tss2XQpSpMfrOWp45Mf
/eiLWIsPW10+gFiyXGC73GSiN7C2HlTBK0QVSFy268JRcu1Q+v3v+wJryhcMdTNpH0gTTxj2Cpjm
jVG84PL90ZyLywKF3/95yqYrB016FLE3lcZiCdKKQ2iMiZ1kYEj1FBRiM+Ev1M1fILcuiBKQbK1g
yA+AFryoSxa49A3lkajhasl5X0uC2lF1PnOJ6Iz2Zc051QiYu+Z/wzdVwwRv4afSzipo+zmIgTip
RGGAfTkIo40S8CfzvxHvMxejE41odVBgXpJu+NrXsTmKUp2SrtutNOseHFME37WGwy8AR8fAcToO
VFZa7F8Dt/0IqzzEnalgdX7p8iw+CiTq4g8xdpRfmlwYgJPgFHJ6CCb6LmtdMdPwAQgJ5ke9dw8p
SGTCyiMZnggKfSZ09BLONwiqhpKupUt21vp8UVJQOMGXbiHsmsjzp1noQxLCbTcTYkR1VNG7Yj1k
m2ztBjdt+sKKDrooKrTp5MvbkAinbDm+NqMps9vwldOkV+80PWlL/AfwU4hJpcOlYifC/BLPBp0m
gTyMyTuzUON3mw0Rh+wvxLGR8e/lKSJXIxphIV3dIUnv/4xO0N7Vy2NVsvEiAhZ6MKkKmZgmiX6R
ttsQDmrwICwlKdic9W+2ReQH8n8I8yS/DhZfBbHYb+SFcCmd86CZMg2YNd5kC2TyvqReNpAa9go0
Fg5icx8izzNNMsM/SotH4eVl92gFs3PJBxNJe+72qWHnczcSw3Uz3VOW/NQlsMfK/4WUiOZVXzqZ
xWhJl17xj31d6YSniTDzl90onidpwwXFpEQYY5Po61W9qjVHIsH4Y3GYO9zt84T2Dp1fzNLBZhSQ
LWaNp7f6+r2v00kpMhSrdg6BUYub9nkaofNKDWpe7pPHwFxRQEcCP/LIeueMLepQjATB4tPL2Mu0
PZmnbKTKVa7TXpz3f6f2SOs6y74R3kB8Y9Gx0gjPz4VgcHOXE+3kbj7wUsZ+91+EbMwsu67IKWCi
cUBENe4P2RtP6F0MvSCPIIBNaxr0l1BZDlkSnQPhAVcoD89JXTIzHPHr5M+TT6o6XYNUQbMWgpLi
JRu6RddOXgqlmvxrCX1yVHyGYXaiU4wHPHTNdctVyf4KfTHEmLh5qjnEaTaHyrkiteRo6sM7LFJG
UK77v5Bae6GImejvC3iASLhb2MH0uXTnKcQlfpsJxeLtARJvXrHWlKuzRnpxE9sIcAKQNEEX8gPm
kw0J2pUdp7WmUiPi7XsocC2qkJlYFucTo6wY3/NSF6KpaOfS5xm9eWOWXDRryEQh4wK9KrTpcbVj
SAU9mJGw/fw6s0MRZln3PkndUEtPqpB8vK8tSSHnZ68IEsDnEmxvNec8IB4gqG4K06AiSBm0v/3O
Trs7CbS58jgygShD+47oS1cBPsrekQ5wff0h/4XBz+osJPCO7CwLIqEHgNv4m6WxoyIQ7aNU3Txr
fz+lHdJr5Bi9chpPLb9cmO3FFSEtwoxPj3N0VVmaUZmMuPVc69NGRsV/J4r1SzEFSGGWKY7ExoYG
ASpbH4OtspQydGTZ4UVWo/mpBoh8o8KU/o2GmLzGv+FXOTNKC26Um1+49KuLEB3HDtAPCnQW232f
t2j/qCz+OJ2Yexp4pcDQRoVVGltka3GqAAzQg/xTEez5acuW2ckqbNRrwc75RPGfEER86s3bHSns
M8J6C+T4ogg5MYKuEkckIyd6+IDB4Q1UkfqAoaEfRWFGxJ0yJ3DPO71Li7lN8ZDIcIPFPYIW8u2A
DUeVAmgPLoDySc1PDY2KkFKgwvcCUMOhnXmYNluEN/sC/SvEFmlHwv7/0oNuJl2/wGbK6Yuezp0t
yz2PiM/iTThwWdX+p9l4SaSAlFhkurJR/Tvjc2nYM/2PqH7jTX+XQTNhnQshQ8MEao6uGvbHU8P6
OmLk1eBXZdtbIQgOFlWkPYGlL/+pX1ExAO66tIcwP06P3yoQXmx21HKKLqdYTGxJKTZxqKaJ1gnT
FBOcu/EP/1wgdFC/LZ5IuvkrfOTnj+IhxNIMK/yjtLd87KbdsKDAoXD88jmbn1GSl5dw3fniHmVX
cgMBuptZPOj9lmB40NelM0dgXwS0EjaSLcX1FCkah+YPN1VQVOAKpMgCbK26tgX/gvo1nCidOPbO
44gFL0B9oot8uzjRH8t9I84H/FMfvhdczeQwymrzKE8eqxdsKHP08hcohQG884zSD7Wd61GR0B4A
M/ofZQy2xgbp13WMSRJh1h/izrRArRokRAlim71Z8lnK/6su7Ws7TiC+wBApd5z6yweq+hliaMMw
l/oyu++5oPmKPRgdpsAA5M0q0IRk3RHAZ4OPec6CLW4eJTxc5UCOthlv5/W80/s8maALHY+2XCT9
/qivERbl+zM/RQxBaQQWl58aGNB/5toGogHSfFEL5J0ae8tO0dFHDVfN0izcLhO/j6MUGURmVWv7
mb5ENnf1/SWKGp8/T5N9s4Yn8JuK2KBLqqzx/lQKZyeeDOx4RPG8VIPv6tALd09XZdh2X4eezse4
rUjqQ3LmMzxqc7O6N2h28T0+rwcp6NczRqWGu9G6GjUVmXPXhqGzozgl2cCK1r+afVLqE8GmPU0v
fcRCuutD1hCceN77tOJtUNZOGmW2AnfvNzT3otavSDPV9nX4+mbrc2oMnoTo4R+acK3KkzXVyjtG
+rKAXYcPUhBV6RfPcc3LHlB2H4f8FnqSpnO2PgF+rZFWkVozBk6p00wl7KGz/+lQ677rS8O94UD1
Z1fBe+ECA6/kCdJwJa2IyFPhyv8HHD6pauYg8NAf8VqCWOFz7G2dkUlIh1maaGu9Bmcay+a4P66/
Stt1KmSZbwGB53EIovpl5sGdqvpCiF+OocMGmXlSFKOV4g66FBiTivoJasFujO6p99mdE+EA7aEY
EH1qcFqHzXnz9NxyqeOjmGwuauq7l+XtFlCmFayeYJSY2nxM6i6d0bhPdw9pTExxGsDsWAfOH8US
BZTH7l6/kmgWGFuZSQC51nRZ5iduqGYYK5o4pRN2BMoV2PRJVCLHpech2Xg2NvBYRc2MKAmAlRF1
gtSb6pFksyulSVz5z9n+UphbU8uhYCEXP63Mwktca4YAsEJiUPQw7hIaJxkny2lxF5XL3X9DGMqR
NVfAvkXfSRHuFmM3ndv3zGDngj6LuSZBc8gOCmUVcHwP5E1rzztqh7O5BTomCD621PpKnRahdvoP
KHWsxGZ+lutJjaFgDynuwmHRp0Us81kI0UMNXUV99SPO3ANmd+OxPH5cUBXh57qBXuCcEMFwlCFj
G7g1bhCGpeGJyOHMA1K3hAjQNAI/t+jgSd3F9j1lhSIgCBedBv4C5cgvAq8JpYqHZGbB3zRCmwjF
UkGWC13XcGp/6Hc73zvbrW4djmJ8+4xjSH/yAg8T9MErLbPjbKDHxtFRcQI56f1p6mWooZvXH8ke
LEwQmM1RHFVEuSQ26gXAdxGXFFIq9fHQb8p/LdXtcCGjOX38fXXAwoMOqejcJkynGERsOyKVM6Ud
PQvR34tbmzLLf9O4yV0r2I6BnMgkaTwA6aCsVHRxr3vrVuWj0fvB2Ycz6UWlZoHIZFZZFD2YTlvC
PxVPZ8gUzGb8200PMnddUK4NTe1dOC/5SUqvsFwr1/Z8cg73ugwt8aCchrnkPYtNajl9YQCt21YW
ZYE6OGuQ7QBeQBSfrmeq4GxzPTHB3FoJB1RYxH2PMu6bbNYVKm6DixKievu8mHMSThFhr8mnR+qK
U/uW/XQoxgPLcaJVS/SvE0CoDCGVn+Icp+U1VHVY93TGnuzEOOaFbeI2cLV1/yGrwEM0cVSApocK
XBqiqETi7a0YUl+fySSuVPG+EkRignoAAWrJ1QhnDHQUg7eJeYUIMRAsZryj9ULKn3eJMYnfig+s
1qFq7ckZB08mJkK2hHEYcvTxa2PSfTb0lUE9Q7nd45POG7izbtfRBh3m/RChScUsqcCcdWFuj72m
VvhEoXbFl1l33fTHRJaHgw/XvODKIQdTbv5v6TJlnhLAOJ1g3QEKV8xFaM4Ygi4UQrjmHHHJ8MA9
v+4oI/yeI5h9NsifhcWX6A41ORkCzs9zEvumAL5Eh7zMdANxIYps6f+41nYrcS2GHtfCyPmm3A4T
tisKlyOE0OzbzOSS6W8vh0wODMh6+o48uzNZ3gMah7xTTUD/KA1y1IK0amTQLMmit3EoaO6Z5d+k
drDolejm73ujcyfqnFGv+X/LlNEffar7IKXUZoVdDsRLNN7em8iij2iNZGYKAigfyFbCNzpJ/j71
THaGABvoipUbpqmpEjNkoB1944HgthrCZ8x6RByIR0atVEctNaadXHecmLIbKJslygwDJ/xs0svr
PlUPDyCikq80/shExhxEkjdHtBi7KvyF/YyHrK34xDmT0CDf3kqp5hYDM/zu6CVOKCS2N+/cO/L/
UVuAZCuvNuUdOIDDAERIXsY07Y38zOcqAdkMu3OTGIDJa1wZ7sS5t/POD/QFXxCn8ZjdeeZ+TqNg
Il/CjC5YA7mTZZXk8+RDfccwN/TzuezKSPMc09yqNYhD7aHluZvxY2ZdlNZ5fUJVAYtvVT+buiwh
zebISmQi7i7tb9h1xezSod25dls/BFdz9GGqCpHnBkfBKcFwjUf5zTmf0gLaUotaW4GsYrm4e+pB
WC3UnPjpQqF+PG/liPSLpa7cJab5xVm2nYeyotSdzFPxaGigsDViOv7ll7gdlbR/TQR3STLMKXJI
OT5b1G8A9PtyXXHW+RZzoXm7u1k3Up+RnH5v3oZxTcn0WZN6uZPjM/xXewHG3ZaYQC5oVzB8hAEJ
Z2+UqwDAqK6/fvBqe7b+la/1BNBC4yrrnYZz+snn7mT8Vw2ixTf1MiTE8To6bCW0bZHwhYLoL7f0
ea7uXIMMreTkX98HVizE/iP8xD8vVzkBFt26fAdVParSne+l77I1xU4QK5tuz1zk+XbmgqFLYZAR
5XqkeQUYsOohVS8rkvzWzFQH6MEvy6DTfLTZjk0miuhSihlrEiTGsG7BoUamd4crY8LkF4+u1H0l
HTYNOZDrTkfy/1as6cKuk1WVZmRx4DLcWPOn88Qw790LBNTWt2kothEl6eJ5NHWEvuonHLBJUHex
U65p7lk8YwaXqgwN6nIf3V4FLBvIufIlVBq79O0cxFma3KTOp3aVg8Dxz9lcWKyZd6NMTreoFDGO
B3GNMlsOT313sOkgXRlZLlMbaGxcZCyf476szY3wXFmS4rfwJukyrZ/tVNfO3O9wEYS+6yHgVsDb
/zT1fCnIR9AHV10VqOPvjZX/vKtK0nGWEPa6iLUoqTu3+Aaem1Z1Bm+buIHY9tNpN7116MvA4xV0
P60Npbxk7moVrR1Qs6LfqkXujEjf772OPaE9WSRdPYN0RwGpgLyHWXPBYG4yHjqPxF1Oo33Vonmh
DfH8RvblycyvLEOJaXgVc6BvbkJUBvbEudMF4bZcpUCZlvY8/5n3g4Owr214WILkW2AN29UVPUgu
QJRXzovuT20HJ3+9TkI2rGtg1ELZSpYwCHvPyuGvHZGJTB9rYjrJ9QrBmRDjfIlUPdg11bJ6hIS1
yu0GAzBt7CStCyiUHriDO9D+6r5Evnx6sfsyZsz52yO5G9jFM/Jy3buxe3BaGjyjoUfeoeIfsrTh
ARLCQeRxqW3+T1i6Dsdw6tcie9KrhtxJ3WFmsnPc+WheohZ8du5pdCF3eApztrK37yTQSMTPTVZD
7KcDyWt9uhj86mF9hSuNjJWJSmMCTmgbTjhltGPjnpphyM/Gf/8YUma5d42qdbrzaFg5PO25PWSJ
aJLfmVmtrRwM9FuCw0cXnDrXY9Ov4/gWWamCm8cwUT+7Fb1FxBbqGGOmJfFMV3pWFGR02Qk3tcf5
q1aHRU3J3QzslSbusozh1h9r1XwbFJ+rYnUfgUQ5c5G+AtrqgjUySRgRoy3ABfa7pzatM63FeOUZ
3YmdUjar7feglAgTNFyxMriVOKDShXYbcBcxj83WJjuw+Ff3hDt2gx0hztofzdyuyvPKXC5Wnkma
1RGLiqWe9m17MARGb5DEfJr7XZZg6xCxclMnxc5QObd+/p/Ai0Quv38xHRZnF9V6Pa6OeSKXZhzd
j8Y4ZmhUX4rDcRbmpm/13ukFn/Z+ewVbHRz0mWKw3RuwkBYoqCcPiV+hN7K0w1eUElpt+hKH4OgH
TIFItZhMguU/1y1zQNvtITKPRHCN6mSTpP9+zXH8LC4jMN+WlgL4Qhf5OCn4CFyDW73Gs7QOzMje
B3JCheM3hJiuLP9Yr1eqbOZOniXBpyHxXTfknXOj6fFMOys7j/5Le6Cl6ftolmOb2AkPuO+1r5VL
2A+Dw7fnMZ1U9+npUtpJh0mwMVc4fa4Pp18Vo6f+0EC3EjiYMgI19ZhQZ/SdyK71WkpbqZJyUT5R
sp1pj/1YyLWw6NSzeOakbnFn1kLw4JtYtXMilKVd3gE/sz29E3uwjoaeGiagwnfyjyjaKwUBTSlP
vgCNY2/g18+pCvo9rmNXbBtdBzspTpXlygwpnMADYmctZ1+g7Vr5Yod8y1MzyjFwkfq8yCxsL3Rk
qf/G4DAAccFFDJSFHFN1gKLMTLsY5zadhGb4VUOWukkKF0Z1NUPmReg6ydBoftU5GOKEfslygvzv
9lDIHXzxc4hOIKg0hl1cNZzW6bhHlDzwOe8zGaK/vM0d/fysQLW2EVpwcuuHGDW7IKXZ7uxEJUfD
YKrzb4dc/ESYnZutOGezb+EpAxa0XeY3sO4wAHfN4aT5Qe5cFdhpQWUogoFGNH3Ie6NHUpBfPrwB
1KlciMA5ns1Sz2xRf4eZgCnfwL+8P0KoYTRNuJfmNsgg+zt86SuthMEVxFh1YMdw4ug3TXZuInkq
LTKmshpNkgjun/kKmK8Pjxg8rfEqzQjgDoVTc67S3Ee9P7EwuMRRak7ARPzKWwXtc6EX+aEMyWfq
JwZo5/9zZ871lEvQr407PnbJl25pdtFBWnJjOvfKuPDpH3qIzxCIPdfGrpf13tAmIYB0dGZDbV4d
gjeYdCYqZzKQ0Y1r5s6a5wO6NpqU1mRk4mvJAp7ZMAGzfFsB02Rk9zoL7Wyt7jUQBisYMNEJUe1D
QNrU0ieEHwRfCEZimJiP4R+QoQCvZPqao1VQsNtqEqm7hNGy/rUZDmLK32KXDMCwrgIDkfJchKXs
/bFSrP/lQutO4GHCNlH5MMQGJOQIU6DuASELu0ePYcqYVSmhz1FTE9fzSIS5eyMQ3jXixL9qtsWX
dzdjlATY40jkblj/USurWApCuNJS8nl+LvzB4UWXnhP+DATpj+AMRBnOmtj7MEROwdVPI2ClenaD
i1t+Zjjqpu7Xxhzj1hNijoEiDiXal4rNCO4MaM/OspDnLkCn+Ac+3v3q+H3mXD2fKOsayqO11yLc
cXjbT4YdZ/Bnn30fdGjgqJz7x3JrcL51qvnUO8498w2f6ZybE7ptoCivWsHjG4nmc9gT2L7UVK3j
ny9QhzBQ2hCklGO0PFj4NwYkt0zor/jYoM3/SwUHkpSlkojX94qJZc17CwlHJiJS9xU9mIpsjeF6
3Gp/9UlxuNlBJ+c0evz0HEueaKeBqxuEuTMXlNCJOOItXaojRRoDQEDTn38YeHa2708T/ELRoSBp
tWPEvtDt3IkiurMlNLpHL+mfJde4mdNPg9r7w1u4wqjmL8z/KgoTL3ujZXVc85VxSVCc6+8ElqZU
qiLt1LYjmfpLC6hN5Gs7zj5CXN2i8dSgrEwC56lEXGb2vwQF8Gn6cX8cTXC11RYMedX4J3qAWEFt
nrokDPa15eZ1MAIx41bDL7jQY6uz/tiq7VwOB7mQS/pFRk05AMFbgFBQlMq3K1W+Nj7P7MZJ//fp
7o5DG2qaeSFj/KDa19/ZVs9sMWt8uuI1/Hx44BATl5DmCbAvvuAO+LMWZ1XCWvupkZiBp+Yjnwc5
V8467g05lEy9v1q9n6wkimS6qdwBsm+jzG9VYxmNQRkrMB9VIgbg5VqJXDF6kWYXZL9tSE2wWe+M
mnOk63darDTOOk22IWrYghhJIQBEEDWxgRZTmQyaeYHg3vFG487tdYJgh9J/935SGyB+aAQu0H5B
ObecPWAjhrgM/xgfUuuibZ61f8VWRvHk4iMHM/vlnM9ZCvOJ6Jzv5pKS69BmxSS0BXug10Cpylj/
YeEKj9o2G+FR6+WDx/ZIB9qk8YXtbly1f3A3aPKTxe3h88ywkn7DFTz0Rq0ej6XSX8/4WYtXr+2R
5r9leL65sQEffPY8LCP9V0kvPOHznH05+fk/yG3Qmc7ns2DKOx+g8+DCOuWIihBrTwrra7RBCGVe
1Cy3RHEQl6aW0+AKobKMIEhdcm1S7oq/5ABD3W9B6GMs0MeaJtQeKnxq1fovq39n7mlqDRUyxfLA
nHn88IKJZs8mXL0Oyiw+Cb1H9RSrR1fWo3Xp/BLEoObpAvzQMb0O4YvMhA4vIesoECZ75OqI3Uw/
nhVha9dwQprkLTXfKH7YdCbC5DJG8/N5MuI1LOYXL0ZI9Fp0GgHOUgOYg52pfjAnC6QdRFC+lboC
baxCJ2BEd89njLDnOlxQulj9R42Ns1HENKWfnb006xZ6xwljUDEUDNLTiDFuhwmMB2TyRe5RBicb
R16xOg1gKMZPELXCIATqbNEd9NZVt6EP0XIGQA9AYEl91D8OZgR4yzL4WdQJB1xzNft74b2i5HoM
4L1aEw7nZHGTxYWgoAW8VqDZpI05V5Q8lOe2BcToHaXana/Ve9DyWBEWDDUM9j+fCmLKRUghz4Mc
DyQHI1MmJXYa8LwfIYh2db/dwEZLjlLaSvkWdq2N+Zh8FTKVe9inj8NmGUOUFDgVmCush7lSB/du
x/T4+x39PGc1c+m/2MWyEXOkmN/bAj7LVTttsiLZSk3Uwnlpm/s1B3KFmIP8zg1J5edDFbWFzJHp
tcrjfBYI7JG5BifJcy5f3UdK2ieyy7zTTSArVsuwEx4yb0Zn1EtWHQvcgPeG5t1djOTvdJmSVp9q
4wYc+skBh73aAuZZyTtuZn+/+xqV+O6iC6xYRyGWPZVA1yDoYjQBMNgaL3U08IA250V//3aMO16Z
wb0F7JEYqXN3OLEcOwboup/ZJudY7yg1/JnLS90SOejRYEA+kGmuRQYdU7A3dvnqGXgRBQIa42G3
X5zuioPkuZMVghLQuvOD+citrwtjovbSDLScOkZcmJxNOSZYM1VVdzyhV5bn0Mkleu9LVKiPvrp1
ekEYON7zw+RR4K1FyOlNc6EUSlivhhMnLyGS4GMLlauPbSFchI/+UcsSwvEhB+gRSqy5Vw0Vwn1y
iIH0GFjOi8fgD8YrBf2njJ4/hIHzYGLeYEJtnvD93fqfagCNBvyD6RD182WWQhyNtew8PTL5rwuD
0jVgwKM0qIS7Smwy2XO/9XaoS8sVY+x9dU++2CvzihsQbQoL2dnJZCCyuX3/o1OKuF5JGx3DMsZx
ClI/XIvG4VgDSEnQttMh2+4pgnrkjtdMzSNRyQKWA8FzR/j911X5Kjw8Yggakh8uuAGdza/t3Gmu
38sA6NdOtRsQPnn0KRDVUsPIeJBjaYK5vVj7Zq8dhlpaI3M8qvTWnRRvQqe7iOIc3bxqaPfH9ooh
zgcQSToVQ+oIc9UFo9Ljq4O28X8f3iY/xi+Z8PEF8OBo8Z3d/Wj1uyC0cgaswvsrlufn5o8UCvxl
iMqLdQbORfMhV1NbtSHNlNo/wjklIqyWpIuuUq/5+0nCpbpbF8zrvZwfxbqDNRoQp0FPWGWVTAfA
EJjmuM8wUTEa+fdtZEe0G06uRLssg+YaikloTgCpudgWJw1+xNqx2NY82YurVYyoQr08bwfXLFty
dSNkLRVKrLdqRhNDJ+3nfRehtlE2TmB3znnXMAh4aw+7vXCy00+rDEH6AVnQdHL3HU0M3RIDypLx
NxLxvVTiWYP4fSdxobaM/dpgUzWp/sa3s8Pz/JDnOCEAH76ynEdr9ue9ESLKRfBs/+6pTBZ50R3O
WGT0y6HlRQQWLvmARCaAGADG9GTYwGQ/rh+0glBwMaQmwV+NBiKENUiEAaYwE1i/5D6JQHOqH5a+
dhA/SDUzrfdksTb3w5ZCEdy4LYYBiXVsAsX/Opr4wRa3x1itLw8/0N1EctG7dNd7sQ+NRhOdFMuf
fDm7P7QLWm2CGSvjkY7wDREmq1h2BawDhSkGx5Rsyz9rfADMoTAcdp7mMdKbd1DAjdJl2FrEYuBT
DE3oBZgnT65GbLYrhRjtjibh0uEvD5yrIr9bobgxpKrsKbfwa3Qe1qJ4pMa/R6LcEYMcbEONMtZ5
fm6ot6vw8oONQ6ONgZI/B2njPhLdZ4DCbDKNcwnHhYS+db+PTfZ/ZzSP99BKCXv8MdCGHiuKue+N
uiU4WrFasgknUt20cC6pYKyXZgudawrWFfWqrZxAtvlvvjnjFN4VWTdH9A1iuh9KcvOu1ycc/InP
O2D7weXzL3LY75kEfDHAeKPiAmaxU9EwoHyWtxeKb2T9tu9m53/yK5FK1NjBtOARg3PteTF1kkIS
01InLhq7H59rxf/vo5CepBqTsaqJtezVV1wXaCPC4zmx/pif6xp0j+XV89oJzlLsiF9fhxrpTGBB
bl9OqJaTW46JnAolPAcNOfafSdGgw5VKLVttzI0csn7Hxsb8CgKHGkBXXC7yaiqjnv6DOCf/z5Xb
jDG5GZVKYloSSnboBH1SaMhzZZOsBfuAQNJ3YE6NWaKcsWnVtynek+hQ2evUy9i7Xjpq730oQ2eu
nhwe624H+PDWQurprxIS0cn70LW6MWXXZ1o7c67KpYvFkbRV13sjcdHXCrPoHDEbCcq/gCodxMGo
64OHZT8qODeY1Hm8I12cw2oKDakpMGAsSeo5RarTnON8o2ZCEA/Q5vH4nzonBs+s5GdXgO2GPWNM
haoxS8oPaVuv6uw31ClGmj2mMm8cj2SU+qa3/dvCkW/viZkSrnJNybeoZcAt7DNUzAtctYDG2+46
Bz+ackaaIT6iYtiMHq6jsSgycA3WUI0sb2yHlPT8b2QLM1L8RgSpnp05cJH4qGRV+XZzN4vDU31t
8umgrF7MS7aW9DLgLkQmv7aW6CAxX9rNoiG4x3L35OUOwB/5j+WxQlnUnKWxr4MD2lATrwqnQG0+
c7sRW/Kroq467NVYWfi3c+9U46GnayjAgTwn8nCDeQPm0OpneJT46JFHqS3+VJIk3KCji8jN8u5Y
8z6JHqfERJDnX/N7Bk7ta7h0jPURMlKV2fGtQDNo+9KqVMPDSckWuExl0cI2XUbF9nOmH7fg7Fi4
axZtmi6mhlt73jaT3bib9mH4zM3jPh/caiN27uxD3xkPMhaWP3jR93s3dVAhyDpJb2BN14dd2Q9B
ctTw5TYXt7CWtENvVQmdTMuPEAK3iG2QzpdruqX9u02AQqzyXzvWHgHNsMxEA9C4GF2zsp/2I/uC
rZndWTIetlOMgXys1QhMq22NAHGpehkLmexx8J6CV2Kfcwy8dzhm+7kS+/Yg6U2McxWmmaSOvI0e
hoXrvu1DlaEZicJo4pV2lH1Zdp71otLL7g8LvAIcyXhecE1SZIR+67reMdPk0NaGM/ohgmAQmS0A
BWaCliLBZJ8wtIotJQlelYXq5BODa5KavyUMuZvt0SXEYDrvvLDuX/g5DuuLHgMJqpEjOxOcBMvX
5ZLP2VJ3PeGlX3vDFDViM4iFHsWa8RNoi7J8pg48lYveQ+39jmlqLQo6Pml6sx7m6vRlXqbs209P
5/acmcJSgk+9pbtp+HpiGyNcmu/J/8ietGxyAZfd81YNNMbwL9hZWAtOEkzSNBhfTqAa/b1CCxWL
vIluCkbyouH9hXroCj8igikThiluJr+uDSmUs0JFjIq0OBAzFIyy0+a16MJmTnV1CMmiYlsiN/yG
jneOToM4bbaguQevaIT5InU3NwuztKO2vd6UEWLBAkGCMc5eB6KE/DB/Nzx/vzBCuxhY4OTpIzQ4
Jf9q0LuI4A0gj8PvjnMrGRZBWVgPPtHH+4ytA+l6+r9F36ufoMqUn/qSBpe+ezLAbNPhYrVKkkJp
fDXjnTIl82sZGliRLAVsWmU29oRnbzsERzJFFTpxSr1vajP5MeSMVk3f+aZ5jnvMppoATDl0Svew
5stbvNbFtylht0SraT4wYrKzUIul6TqLI4AcfL3pNZh56IkxJgbo4c7bzUpszpL28AdXKchaiNCP
KxrvKM0OKP+ShBc/jtyPUfy1oef8leTRj3e2xv7+LXxmKagFnIVNFupnZMMlutJDKAMh5Hw00dhY
gLgqX1QXeo/4P4nsJZW/z9XGxEyFtw9fz/Ex4snDb81QJp09fG9JklZy88BOFRgDxB6UB3yyiB2S
CT5YyfEE/Hct7F8pOMCak0Po3cAw4kzrFPZ8tbinouJ1qtc0KSvKMl+dgykyf01I9/Nlb6uuvxtH
C7TwoV7vVeMbJKZWrzGGia9ocn++jm1m60D5K90SImxHjswTm/GiKfa7hzPoDsqJD7OccvAcMmmH
i/XW7YD0i5eBHYgoXwstw+T0D6oqGiIT+3aQ7HMziidngf3fmQqLeuzRJ9C9IYM+SgRryUtKJDtV
aqgtHMzmYxFPtTm0PD0n/UW+h/cy7SDUzAwEs3Qx2hyS9PgtHYOqaYwbjO7Ez+1hKc+x/bQVyjef
NuTf/OImaGGAesaOwUYmWbPFvMn+FVNpnO3X56iZcVHg17Hvk3syvRg4tt47xgSsytl5rh0nsMNx
Q1sk+iNQPNZB5Y130sflmDWK0X25n7Oznl/VB3on6xxVVB7vB4PXT+pUZ8O5jKZqo1Ri4u4eVs/x
wo0DkcNrdm+cakQatBOUydRVaChB9bV/Jceb8zTR5f56pV00gb21F5o0qWDVuzRCh9cVLaNwgKyC
1vKwhfQHYGtbhLEyGRBkgTHIdSN0x3Mv1QCZQIJIG65E0PwJINPOUWH22LxnTGmERkZ9dd2VN1x5
a7ppwjYDxtskS41rnC8iGLHwHXcewhHoSyD/ktE3ihpqJ/VbsDYQxNZsPt+QiXz4VIBWskMwjVg6
oDOL1t43zTgsSsCI9jQXJd/UhT5Dm3r2HjwGC0sjX+mCcyiYY4nRbNjFE3fxmOATy6p4spgY6TLn
yh4iDAgBT+2/w6z0HmkkAEXtglJeOqFTQeVvzzEcbybJiJnp8DkeVabsco5J0z8je+lU0xaTaegS
ONnSqGE6bwh3dEWmM35M3Y+ucyabVjSRoep/cBkFD4aFkAk813uoot2m4rwZ7w8NRzAiPK3glqg5
zG5sjCCPkPYEqowIraMMSFsPc4hL7TPBGy7n4m46aLg/SzdqT4MnTfqwkaz2EOE3QbBbyQOZYp+a
2UxvcjZo+gbsvR4V4HUjnftixFvHCg+8E2cWNlYY0YfevaCMhMtmbeBSZ0k3jK3igtAFkKBSSj5A
LK7MdHXHHWlY6I7FEaYnHGVofJfSNB3NFaDSP1KF7pkJZebaA7vs78RFy3N+D0Q/FHdzsN0m6R7q
E7y9q4eMmU9pBwd+Sd/6/TSt/qHLikYvzVsPA2y9uFzxE/wJglxSHjs/AFeo/FyxplRJaHiTjojq
WmSEZZvRXiZmHBSfmN58VPrD9LPs3LcUhV7GRUsMilVKtSwL+aK5lt4EHjRelp0KNUqXUPRRr0eD
Xsjcyg4MfwZdblXuuEqtapnBu+2bmUyu6BlWd4Wsgrp0dcZBRvUB66Cxmi7IdPNPj3R6kumiqybY
Z1/yuFEfiUMyxoga2FtC/IJvdsa1b1kP2VK93IEB5INdgDgXd9ynn5WxXXGfCcC19Dkdq60rI62X
RBpEMcSzzMMoDWSf2A/IOC42kWSPJT3h85K311a4EsKi9uus1AR9VT7bSMugdWzPXHWMslM/03wZ
HqRJIoLokaeJNg6DQTO61Ep2BemBOjkGc8mo1Iv76ravLSX6feC7VqnY48UxNuIHsTZPkZRDDi2l
WEdKsUd0t61yiqcpcRmXTwSgUSnb14dzhFm7zokNIjw5UWyhHY8XZ9B5ehA7U8pO3ELNPBDSMYsP
rEAnPpQ/CoHoQhHgbo5ddBOhSb/s7bIo6ZK6PGqf/n4Ar6dan13W9zsgzaEdOD5yTsRr9mnksOFD
KxfEz1QrYf+aO0L+ozWkpNes6daD21RH66p93TOwqW5Chb7oISeq8QD4Ayy/2sghe672i4lJMhR+
k6XkiW8+si3wQ375/lfZ5H6ijmyNbqiWy5kNlgagm5mSHA0gUjlEmvSKO8kkDDZjVqoCZAwX/0GS
z2QH8PvKveS3jUic7ce4UzS7yYHwEBGPVVwz+8URJY4uphY3gxGUmXTOCWdi53iqwH+/zTCh+dsX
S4JLJFYHh8tXFFT/I8xUqCdLLbgnItmX/ai6THeCcixXwNrVTZKaAvfUuTgMQ1P5S5dp/1vZxm67
4aemgDCjZ0cg9hFZMdSg+7ItqyNNGOZ/s4+3I4OX+Km8kWy2aoWrpKGibnm3QNONZuwR00FouTBI
CteYo1Q3zkXh9Zq5Vkpk92cJd8tDdu+m3wdUsVDYqcM/1QnX7k3nvC/+uviDj6vIgb32qzlBbC4X
6XTyw8i//cUrLPrx1iZw6eOV6ZBAuK95YaXrc/GK6h3A2FysNQENhAsWTWGxl68GkBMDhzraf279
9031Q0b+dCgbgxAA/5P5t6RQbp+1p3k6xYdH/l/Mm66NTTQh5w6urS1zSbKUw33PaB3BRX9kzvJv
CMdKv4nCRYRM7n807pxLUY8ri/Ka4lMThPw5cL8HesERIUWPpuyAVtphOgEmFoq2hMvMhFof4S8Z
WaII08CA6OFhuPn3DIJb6OUBBpcMnyGsV3raciOip1krW/c4l/ch3pyCxocHCeiqvvpUjkGlOGG3
iFeF4O02GemNgLGx+bvzzIAv/5dHK+bw7yXQ4iXsm0Cu9eSymvbtSylY2+8zLU+Qo8mM4u6+qlgK
tyqbVALZSzsKhXue8m8kUFF5DXOfXnZXwcGO1aeSwVyOxk3HMWDoQ8JeVSfZaXsolXgPvwxzlrDC
2cPRg8B/dsIuD3lBZvgRloxzlI2gDjxX9nDY5B4mPW57HjsNffXeIu+GEECwAZtyB0wM5UOej+OC
yZzdQ2E3Nctv8gEIAzqlkQ8cTbUj6sfkOGBxvsKZNjBKBWchYPQBg5pFuJeu9fkikbhSKWKe/vef
wo0KWE4ht0Z1+E9i+IZjR4JgRBqlv6IOzzqeC4n6oQXjoinmuHdShlIFGHvawd2LbGr0j2Dui7kA
dxQVjSRLLx/EPiCaE0jtouCMaKpuldO7R4VJGecmXnr7deUL3Jz7Jx3d+2pav4aiK7VrhOOLdgLc
KB2vNwqj1DJ3Fs4jLxswV9KyXpII8/dsoxuz9oteQJjeOLRT7TIDf27sLG/Df7+J5LL6DeylZSaO
DSuak1DuLMu67wZgRaYs5ouiu9ncRDyTX8sMJNZbmTPtcYHfyfRy48StqwIZANOf6SucAGe2JAQo
4EI8TVtPpuT3zlx+JwfXj0dHkXyiAzCYpaCgFXKHLXDbegmuBdcnOSUz5cGN1uLxnr3rZWoKVaqV
0Wp5ulEs1tSfUGIFgGcwPLAIwRchbooImhjDT0cRDM7CmIt0ArN7Mi4LViZf6DtjhCBe/LQe5qWU
MjNUiLMhqx0Hp5cOFwDhZ3yGpO/PM0SDCLHClhfqKn5733/cUw4gdUD1sr5XEb2LM8LAqDs9WD7r
4B8WBWXaWYg8d0zf7Kvn0cOhykuSbP2l4zV2dKgGwTJaPI51SNsh4FSCeQdcmhZ6zXVV+G7OvejO
uio3Thy2L7U1FzoyJZ75PDNl5i4Q98WpNAKmjxsB7uy10Nzyj3bTpEkGGX7+nxCl40Cx+81+k6Dy
2zxfN8XXXSp/3cZ4rL49Dp2DazLzPWM/h4lVLEUrXHsKMOM4+DvXhTwg+mMJTbmuWjffFJjOz+D6
TuRhS7UVaX4rhExsVmM/YeteLN6JjrzQqugXPBQWzcM+BERSHuZM/dwcQL+0YwTQKOE45Bt3eZBY
XU6PcVRnypUa5G5FVrZzKhjeoKW4qRQ0XMft11TArYe4m8yYiYphybYvdh3P9Zdiw8vMPxr1EqkO
XlVvGwHUvAPpkzkr9eu8UhuMqBCOPDihutJ91LJMEQmdCvetj77XHv9sttQ6MOq4GdxFxHmm90eB
0sWEKT2jXLfTp0dL45zbdTtj0XTAnaYuJLOAc7/EFTsrgXGFk2l95gj2lO9sjoM0Ek+pJqLPhEP/
bLY9hv/7BA4pR6BN/h5rQe16O/snBaoo01ZBu/vl92QTphgmeC+8hSazm1ibM2bo2X11ud3VtLZu
gTao5gugFRK7bhTxvTL64sVjgZcA0CZEwhp3M85Xk4bOug//acSjLrAuq/CJcSWm3HJ7RmsB1Tpj
J+X+pI5UQcc0CKCV+t53Oipl7HLvq05msUsgYFNdEGP8es3MLvrWU6WCR1KgHKEGEpdp9lt/0JsW
KchZL2ZvzPCB+PkUZTJSk+lfDTFk0IUEPbLHGyPz/Uwo5pQ8Gl1Dptatxr4AaHi9dv+RnTp/H4JH
IU5dAGqVrzo1cCGc/aXKw4T7CbCC8Oooo/I0odTZiw1uOyIEqM+hVjHYWV1jD06QRNCzS3bMEs4N
vlTJ8LcUZR/5QGQs50v822fApySfGljz25txzQKV1a5NAg/so9UP9r7HqQxflNc4H2B4pCK93/uT
TqEEAMxMG8JaGu0IoIUc4knrX2ARzFx6eQ2CXXYX2ibPNAJGz53b4f2FVm/s83t8f3uVfN64Pz6x
A8u8gatYMqEQymycsO0Q/HDEc/ELuxfSA8cO6e9+q6t9rGpibsiJiwMW7PUSKL3WjoU61LGZCqt9
9XAaw9MihiJkSxOsVpqTDgAW/it8wtBoxwSVDjQBCm79hkal6NsOb6VwR+Ga8B5CCE8ZdI7jse3B
WsJueuXf4OKjLm6tyZmbNz7OxBLUQhJ2/UV7TOgcKwxxBvZ+AsPqPRg2u48b3Dh/JDQ4I2hOzSa+
FLfqRJO7tfU5cJwgXx66NLqJ3vjo8pILMoUrGrbzHlq90r3qNYeqVJnsW+QxBAjo2TIjlgmbbEty
hDOtRf8eUzveKxnFNVkhTQNamCiBm6flyxxCQ12sKAae1qdh9xR8KB3jEh1QkaFa3bQZWxCWa2It
8mGAcVVutKUh6bt/I5fsHobCVHlN9BEaTtCAed/P1twq3j7bqRNY1udYJ6XV6Z5slqf5ymqkOnJa
7nuWAJ2o0CSRyPQksOAA/ROT5XB2oI+sWywqxxrWwRJViqgd09l/HxQn3O/enN5WTF10beIPMvxg
p+uWoxfb7gVb734C9WEuJr6Tz/LCtzV8aRnvJ5QtCnprALEW8bV/5JPlrA1TJPXCrIUywyZ0JZt+
3FsC/0YboQ7wyxL/uJGvSkk7NhlbMOiEqZzcvBPy42pJiwTzYg64prmPvSoCOw5yOtLyg6DG6FSB
UgQm/DHYfULLp5/TRzZZHUjY2RVJDOIvAGvjCoRHAy7UNyrq1JE3p2IIxam1fGFmfeYTVzsVbLca
k8TPwFq31rG5XFtOzWEhQRSxaxBW4rFX79H9rqCGRMCranhhysMpIDvTB3coH14Yk/CHAT+rGvwB
FF9XSx9G24NCLK4aLLW7jgN7xhYdOahPWUZLICwJFlmBuhToqNmuPqwfCUBS3F3yOa22PzqeuURt
fK2Zr4rM0J4bXAenVOxdZNrcRQmCdsYJ8ZJrlH9SuBbnkndXG0Lyi6ZlNoAzpFKjDgdHo/RKeO7N
/ra8A5yBVCf3Bm9jEiOligwqMcfhU3J6PGF7YkV9uALES+GYg4QeoqRoPg7gwWO978meFjlBoLsQ
B9nBvA/UbWrh4TVfvaRqnFpgSaqDVshPobIMsDX0uQcRIjIQXQtJx/dTgPtqTElJIYLJ9vZg1Jq4
PacFK2Bcb7wo1ye8clP0FOxJSTBhevHBPqAy1AXAO4naG/TJPw9EeSrqvFzz+ejz8GNN6pAA2nRp
zr1rV6txcQtFUVgkc/ociS/IztnTHw/1ZoMMYLlRJMG3awqht1fN9brRyQzQgMzBhXY790E85c7q
1af8DJ2eXO8/vWCp9XnTjMppzFmnZ7CqK0IEHqzRdWvJDse8OowNVgLRbpEOswiHkYZ9ekN7VnFe
1RKP8EIU9U6uNFkxpEGhfhdp7hR7BT+dCLK9Brtj4OZJJQQxdkA8Wz4SO6Y/TqnZMDBrMK+eIGHK
7ciyXzDjq0iSjtSCqHKMu5HBeqvy5mO1Os+qkFFph11jfRnM4csamGw/eiWIcVVJZ8LuY84rjgYE
c6HEeuh6KJbihc0zHQKvNnR+bpK8+YjJCv9noozSM0RhbXKktCm9PLrq9Y1S2JmSIXjcAA0TPzVC
sDojimkiuKDygTsZ4rRfK+QIS4s8n8wfwtkPIf/7Pq2onAK4hTQuU7Vgtt9lVCSWc5BBH9LhpelG
3C2o2AYG8GsBKClGEBZNMAmFRd5/s83QciZR0kUTKYe+2OOPJ8DzlfR3AF3ZGKwIIzJTJ+FdfuOH
EIXnN1+CN1WfQLY5QDrXeBZjmnV3p0v6SJ3BxQP0gyafhR9AsqZqhJ+nqmur2H/WMziGSalgAC4C
vGHhL3t2dFdgwRmVlmQukmQfn5IJU/BN9+DLgVL0lZLFszDWX2JVmP1SR4CXW4XhqkKAGoxm5l2k
++6qi1iBwSfX/2VOgAe/cueuCOkCmddkt9AbUncAhYszIMj9jT/77zoq2uMbAYy5+KGuPojjbEDD
h9CgjJTtd6WQRu0FllwDwNhUULtxGyO7V5pA9z7mC3ywwEkzxYTi75Qa/tpWlPyxcisbkKa6Dogu
2aTEfeK9Rt/acPw0GilqoSjuLuQkjj1V3bspISD+RYcX/If9yFj7WjSU8BMgccyu91r/woz8eQfq
d7StPenwInFky9AVbr382JT8WCusTx2NlIf+jxb4fc4PANyrnHkHoVkLlH8wBNw3U10eEdXylb7+
1K7p2ElLZY7upASbC7gVt6YR4YhEzDUaW33I9q/2aWT6YJ6YoHZBe0TCRkFn/jp9gnhV1YLo79TG
EJO4Zsp+gzEDKatPc4hbviGgduKZUEfS++Kp0AW10UUXDboTCa10nNqhsailF+ExlrRfSRgCT5EY
0VSbNB86GNppaQjwil9CGRSlsp3BvREAjeaorpQT4s8YWq9gyu/ScxTPVRejBen8qr3aaiDhiVvN
N6t11jMyuFLPrcwaVNQnEnCAnABWBEFwEN/9BJbNjCcrRhe9gXfZVVUZswUnwE8sIeBmw4Ab9Vaf
JA4vUjbSBUCYMmD6QPpQLn2LJpaOjZxjcij1tgHdxtcys8YW83C7fR2FopqTRwGi0ZHJFK6hctzU
eNeGS1U5Vx7xxEBK0BKCLe+9FCZwM5jTmA9wLW7JwxSJD/sbfQOi7oiSLzeg+P0L467RNnOAlPuU
Hm4+zLJSKBNxcFpPyU6Q9ZWh46JoWWy3M2/vI62dw34sGD1N0CgcIXgY9rzkYjmOokq+FP2NH6Ph
eC3ubNQEfS6IMO2y5D/h1TKD0tpO4Fc8SfIlBy7HgkgzPkCJ3ol2Cbdcz03YY/DRLF2Y5PToDvw+
UnE8zDYVFgwuKk39YCRT9rNgSkLccJB4iQ4oW+giXVJ/lhQyz+qRXhnRjCXaEZ8gzNPB1KyBlqMt
ml0H/chAXhI8cgjRSduY5cC/ub14KesK6ehS1IvFcF0aZ+sORIfLDscq6N0Bj+uB+lGI/MRWU3xB
nwldIn/0KYTEZzxn/LM1T731AOntXw8prZ+Sleh5KkgWymtjUbxA37vx34QFJzis7IakHYwHZ9lp
AXaGQ4MJDIJKkq3XuSeTw4CUqFyCLEgynwMyIHmCf4WuN2Mq5QbILvW3SgxExTrERfzI4H3CjMyq
ahfBaFONgabkG9PrM/DmHghuHSz4HV/lBRpTKVM+54ErmZr/wHr2jn/duuHjZ+P7Ty7e/U/jDexu
PjGNQq0auKWzFNFQC745sa6RffHlFwAB0zIosBAjvx7cELCZj5h3g4LlDdRMCyO+U+1R9azxkcg2
dMnj9JDsNw8Vx8KXmMnY43J4+EwNYUyjYfMmAGsmZIBvtWMIDzIR+p3G8u1wAS8FN4mRht0OgDdj
15bnnW+CH2j3h3c8ziBIGkiLXJTH3qPVtaZHkxbWV6Zg48045ZrcSF2XKB1k1/FSsUCDKk/luPNE
yItTLHPcHAT/I1gksGFsAStog5FjhCwlXpAjmb7FbhFxy2c1b19TRP0D0fLt2j7gJ71RaQTYT526
2481G8BaQhUHnQcIx9vcs6dNmKQ3i3/drWif4ubryQia+xFrL/AT1YSu8UNaoAh+2KzxgVBKPssG
M+jA7dGk38FbL+SD1JbxOfeNbT74cKcPgZwefchzSk5bzn7L9lE+qO5FARoPvg1Ebje+/kfWPzUV
jzFErqlrXeY8sZe7qkdVK0/BIfg4ZdHsgfbc6yFLsTOd9x9mKX4LshEMTl0I6HUc2N4abF0e8FER
sztS4QmBl/nG2+dfczI+sBKcYf7SwA9jB47jPx35j77lWQM+uT91VXwmL2l9Q7vVna98RCcFg25L
uFTkTPrjcss7XfJerARcVThmK83JJOQWYwlJ0zO2e9fxbDqihI/M9L/X6dEpX8dD+k2OeK12QeSl
LIs/LBxwuLZPrF6yzW+D6tRP6cby6JEB2yJzZqoeL8z+uSMUyNo4yK68nRwLNCuefZ6t1wHTAjlD
HdVO7hsPZ9KKlVD/Kwa/z1rYWIBii9P5MBBCoqS9wfK8AC0/CYf+/by9MoUrVUcQ6J4mdjKyNCj8
4a8BRlTU7Encc+znwrJAgGdzGsgkYwiyYaNU7ZZLe03jYkHsLgJ5ztwt8XvBX3aUIYZN504qoQ7Q
Wj4BI2/3bpmVNMveS8p0Y9wyQ4qSSCiOZskwD6RYdqUy9pfqc0qUIDGEyYQVzA0mviGZO8ugsahY
cuV7evdwIbABH521Be7zyphbFwTYX0NThL8WRfJSv1W+eu7MpEMhNh3wPGC9ls3nxGMQ4Mrk9LBp
PbuIt40WgMTv7l5/7300CiQngNO2HeNfoB9ihO6a0o2xFy/55oYZLH3iQvCfBi6GdoCkXUv3da1c
YEaJnhy33CFzTfrjlyKIcqp117pkxb1VdSPKYlEIK6jQUfXWyfbXK1ooXj6Lq0fv3iik7xd9Z4kd
0zTuhhz8fs4Tnt9HCAga3EA5RPAfFjAIdriA2Np78RKCNH9r1x1f2lak8Eq/4LkhKt1jN2ks7iqk
3I0eNSYqMSi+3+3mif5dEUMREc++UiaiBOnoDLqCRAGQhFH2pdMpPa02WfZwGDWEWGGkqzr2+mu4
zq6Q6r3c2hqhsMygqCQsn7CYa9Oi702sUVxittaJW112ThAIlbWHRCXwz0b2UYhdD7Z8sr1BdBy5
ovxC6oPBwmAhIMHTYtfKFIPsfDwMg9XUdxElNhfSfHdsp3f8p1Nwrkk9/M+8q9epMbLqYYjPjdtc
A5uSkvPOYllf2/QnR86hcgl2OXnHiwBe0clIDse9dl9Imwbx04mAUfXqIfk9nhq/8LjwYnSj/MDt
cKDnEYlixJ/P40P59Vz83VQx/rWfuUfamfA8Z2QiCRkHckyzTTxo2D0Q1iM+6cqrqSuRE5n8xGXo
Y9U378VkpzRYMlZuNJkHxXkjUaqy3OJEA8HO+bd1dV3VAVw3y0h1kZetTv9hLkxof8T5/i0zVq9D
uVnfwyKOn655O7Spv4HPBPCBVrQMCoj3sE1/mX0A7LZ/WUcwH5q3USzPdbLqjc7S8qZVfVT5r52J
bhTrbiBvK1lHx9DnpL/XtsQDG9Hff1sbTsLH5UplRIV5xNvi9UhWnYNJIm6kbPX329yGQHWR/SfI
RjSnHL043OxzUm8Po0ipvfg4cDgtTgD5Bq3Qj8FE0/aUVE2e3+VwDM0U82NIZiFK03IEAtJTqZS3
6SKJQ1WG9ukq6vyY/IdP22UXYv0i7o45xXXlicwym41WzEinS3NeFEBMfsmTlMLbWwgYKK01r2AM
SpatO/NvT5SFhQ9GYadnHmoFbNjFFch4xXn/ePU0WYtlwmn+NQp1WDq/IQ+qSYWGz5Gc6FBMWGy6
rtUlC9jFP+V9jMBt8LEXx/7PXR6y2m/Hd7OrmaxRxWuDhK0c1/hbuRi82S4QmQsXesTpOdO6Z1Jf
/lOu0MoYFSLnwD+P1+g4jk47tkAbH8EeKVEG0x+aVeLVHQEFkNZPa8TnDPsIFhOC5/UKstgsOFUh
b7XpZlsSrHVwQ0N3HNbHGeNUfsacgf98yFM0mtl2W5846KlIC97w4HnVpmktLAtte/TD3RHetnyz
/zNuQWNn6B2EvFQs2by1CbSOtvmJKskwc0HW+RBJhrD4TgPxLi5/XZPNGSItUdfEjVkV9jqybqaF
SbxkWn+sIpnjOwQSOBkJY7RtfQK2fbQw51A5aHYs5Dm68+9Dlzh/cOrcYpcLPetCbJsHOtxPsTZl
NOugVMrXopuqQXFE2ymFW4TBS69hnNcomKgRaBdF2PmJmyXGSBcj2zSDB9EcpphhvGC74DRK+UA9
9PZNaClDZ9hrLOK6O359ki9mdhpqKc/+TjVZIkbuwr7mmfjhvfeR1J8UPeOatguxfufV2vfS/bOF
kJdQPsckQ1hXtmHHdyEp9wa7tWhJ0oKbUu0qChGiRmfDGGwhfdhNUSLSEBKD95sdda45UtVF+VOR
p5QgI2/JYukVlHWbkFNhzCVy1rl4Z4a8ndhAgNhP9YKnPQPRtURqc8Qd69hKcwk88yf8CTHtKzWF
lS6wpsf5LifunDv8/rmMcsnz4h+FnyQ7/K8tHY5HawkKtufoMO0/zmtSVoiGuLbOqUwECNhXVMgp
W5FB8vr8zer+JpuDmih7l9hHCImszOrvfkNOTpJNvtD/hwfG8/7ETOB+bvbAr+d7Nfb1Y8bv3Wz3
gSzQsGkdanOg6uBBzlkZFOY/E2f9ryEjtqyXatz1v/v5RgjHxeeTeDgWHkwa8MGkb8R+5gE5ow2T
gRsMCcggHz1Prt/poF3j/CcoMaKrW2CLBKyOjmlYCTDYROGbeuj04Dxo7xaETg9HuBnrn8bLGbRW
FnxBn158ulyKJu7MFKLcPvzXOnivCIrYjgNZSsyVZAyq7btoCrYSy7m/o8Tk8av4WIFjJCFg869o
gDpy8MiInTOUTnh6CKuIqBf5Gw3od9qwguFoqS9MgtbslW5yNt1pZRjTSP/rC0/rlqErShDLalyF
/ztJPLlFg/QivWSpTAPKvmY1eV2RD0AS6kBRPAumwKBhzOTI7fYjOE0Mk1lX+myKhSBnLWfihz6J
oEHtYUX06rqjWzL4Zt8qX9RdtgxJFwK/JhP6dh0RhVKqM2nFLR7/kgStCSKKqgc2DTzy5G7nw2yE
QZCaqkOkIYtGX347h+xmWhYZ+6AsCkLdzQMXQNNGgT7kGu5otI/gdfSVazntWo5L/sNmQDomNYG3
MKLNCCjRLnpbnfg3yFJwhl77tl4VLUnFh6HgewiFEW8uOgGFg11ytpsvPCN7ozuBzaffEg+s3Mxu
XNN14b3pPSF1zSxVs3OoTEbm7FmeivqO/Jrn9SuBEOtKLQiJVHnrzgMAmoY7WlNDcY6n2ud2NxWF
G2qig6Bmw5us1gqJXz3tonsl+0L/QsRpcbIGh1Ngz+2Uh1Oq4e4C0q2HaemfIiGDHA99xFV4I1TX
51irgo407Jx0dRJ4ILBQENX6ulPVRl240/PhIfMCK1cxP/MTVIPftIYcKoa6h5qLEDfxO/0sK8Vv
UzP2nXv4/2Z/g6uObQtyJ4UYWkTt0DzF8JBiYwahSQ5UH9MP+VtmyDI6l5l0C4ylOgJ1yjIASkPf
GDNy3EsxJwF7Jrvbb1yjOFCBLPHpINykDnjyM24qsx1KJkrwrMDq5MgwRxaxpcQ5ZQ+OBp+6DSuY
yillXmJMKZg1bfkl1/KKMwpCS8zA49yBSzpmUiA8cP3bWjJ+KcEIBqugJzUeGbdnDEH3fRCyD6Bx
XuISt4zC/zSYKZ+ugWnI2z0eF400GIlM1gA1BmYZEgso3eBRASc3IgjstvrpAaz2JWcRweHZ4OW0
JSwb9UEszkLUhOeq+875UnHYk9MXYPlCZULQoUHTCwbIeTM83suhq6MZj3tlwzD1w+4uZzoqXs9D
eWSISYay47y7GDq20dQVrMYOhUBRmQLrByEVzbHHQpdeKO4JQcHnoPrmHhYm3tGKBEpOWMLAgc34
e7vPIVHMZSyKxFgAlJy/RNmNUYP7UmwghgX7y1m/WxNMK7axXIhn7yJY2nRPndSJrQ4JqxBgtzE7
PZ8BDVmgb4IeQVuhu0Xo+3RAsX9WTWPNBPYDz9PJmrsflRcOOLqwlFa7y2ywKPRGMDSx3FRpMECd
+ciGhmD9zERRtYCewKHMFytDpzFJFsFbnP1wK29eVZ2bhez76QsFzID+zAkdOnKfrQWwW9SPNdtz
98uyjk0+0zH5Hb0XvFUkKNd2CHBeaGnSeEH89Y70vJ4fUezbvlOj7WemUXyRGRXnjnnTToh92+4G
C2M8NlyEqiy4n1U42B/zY1N55Ux0aHb2VTV2UcFWTQM6C+zGpFXeDcOUpc3ETQju8Jsx+KVQkhqH
MDYBTpjbd/n2QY2SDYs209hPqXif872IZaZVbCR9WbifZK81v0h/hnrG1XKhuoi07e46XUmyZ8OV
46MoL/vAJthAWq8l7FW1elv/2jCNums8GOEfEjk5aSw4kKVSKh5cFwCsgNVwoE/B+9oEI+QkqUn7
e3JD7yk2No2a+dUq0Mv3XhLgi9/RqfOF0JgXAGg+r8quyBhtPJdMLfiuHmNWrZ8APy44RRxkHgRW
SBHsd86gjem3viaEudo+NAexToTZ7ZybXBMccz1eflhxwmQA+6+OaFTVSfWBtsKzOjFas3p63G8j
aG1aIdDhmQZmgFGJpeIwYiK5Lib9pZeAsaiQo85ha6YfLZybVl9c7QBwT0Z0vcbZZ4Gfh2ntNf0r
POkgxoCQrCnVQclQFph4G9EDTwnnPL98oV2VPFcccLHlCxyIKqwuwHosAm6+KwzIehLrIdWV6aSt
2fDbJ1B8ALXZJkvSnbNRmdFi3Ilu0U2Rry2TwGGUIeOfEKEI7VtiUmlNQfBZEGeMewCVsixAlyie
NTVSu2Xlyb6rGM3z9VDJ/gjtqxrkWmEjQJf5pyBAIJBlWjOw1cjT6zbhbTenDMOeZrPX94t5q+qE
6y/NcZEg3lcrPRAFGk1hlSDLJMoVFqv5Rq81eFvL8W0Jd4phWaN5wgNTZEhZuqtb6ENFNhE6X93c
nEpZ8yi4VB/kSSzIGXDinSAqRmq/JsCvBUZ9o3wFRqT/dywGUb0iPbFkMFxppuQ5ZVcbq3yqpYTG
HxnNQ2o7ZLQPCIHO3mMsUqwlIlvFsGPP0X8UBJmpkX+WRE24FneLqu+V63jXGFM37re36361LmaC
21Yw9/csPwTpQjdVrOJCHb8XAjSPXX9fVX4ccRtaksNAvfMja5c90h0/HwsmeWIasWKre6DVrXyc
6C64Z+RSFVxh7GUU7R4MNVBN2Z6W5wfLd/QIEr1naltf8T97nVXqKrFZyy4sW9DJrCo42o6ZQfei
WlRFspAhtvq7ue1I9votiHOVz5cDq05p7Fi7baFXq2FqvRD0qVdBBhYScd1F5Y3lU31fEmR6vjH1
GynDyXQKMT7Jrq95TBU7dTxOd84qxnr8paZqmFMyn2eG/f6T4MOIeoahJp3HTUgMCib3xArwkGlV
YVprvzGbEjnrmorAhNVV+6ugqRDa7edldjm2IPs0rvY/K7iBd5+7Cm0kPcWjnCHoR2k9Dopwg2yZ
ePERb7GkKVs5RhQLV3Dera62Xb4aK4uVdvpTtIz9xMm8MyPfTpTQyRou7r6WjxAIFHYqG/Xj+rNU
EIKmzIQOxHfsnB/gMg8cDG2og/EVxDa86wlOWtWwDhg3pp6FL5POsa3MS/YvwSwNllEkRZy2vr4N
PI7ux/waIHkYlDSy0R3+yKvg3EeXLO1mKxbfMC5W7hOAZb0HOoAQzVcWtOnVBrcasZiPzCT3x1bf
Qck4LCmufyQ5S5JYBumfROcO5CBF9qIvEovTVTWyEOmzf3cn0d7vWN6MzWur3RNd1TefajSEMNV/
VC3J8lzqYhzn9XDwjp4tmQVvMGwGU7aIHBNvrA+3l9IPGH/vnT7gi4j2sumM+aJew6wBe/xDH2Ow
B0lNkKPPnIo4tk5h/Q2oJcOHq6hbwY0ILfmJktbSuxWk9xKE33yuXEr3T46r2/sVRyUaEz+Z1B/i
qt4mkpw+IWz2zM1+zUwibGWea9EnesoMp+ltfOHQrXhZs4UwCfyyfJSsw2O7VBI7j46OYTOGSNsV
pMBW39ST9oudiier0bL1R4tTTNlSKNt0FyfTe8cIllN5zISeKqKjjG7RJIhK0cu6Uw1dVeDUcRRJ
8RePNhhbpuZ2hkMf7Sazpp2PCF4Qp08GmEbCH+uPv9UwQPVpr4N2letx8nSdH2YsZwc5XIfn2r0W
cWG7mSREcazXWCN/bxMdWkW6RSK7oYsRCn+X3lKGDX3A/0QkAaNTAqy3I6TTMSi5Hkrs/IRQYfpd
0ouDT9BU3iViKQa64yw/2w6m4008opJRsh3MjsEM6Jp0b+Ioz6+bSyEKMKN24ek1STAKcSu3Fj6h
VgsxQkUqSUwmmtFZWBPpaXnogrpHGEdBLpAF3eZ2qKT6GOyy7ywLc6hD8PIleBTkA44tnn6if2tt
HNPjOmjtnmdPP30ScQQBsHQAl7mpxV0O+cRJWmcUCc/+VemTQltnFI6DcwL9leT5rQaRaGxRAs8G
0Pb6rWqojvOCWuM3bbV5yG4J/AtN2CtkmstzoZfPeYDajxdv9e9i/9CBLiZJjH78THPstcfDcyZS
/Ac8HtEftsp72mUaVJ5tCnoU1Yi+Sh0G6zXIXfF2fNeHcyLsA89fdbiVcHPv2qfua0QM33s18wfv
8SReShzdrRa57zaDUcT59Y+JVoebIUOsBRIBcyI0tIFxfgfoh8dB32Ph0E8lBGMJVzTyi+Bl4Vhz
gIwUC4eqRR/dC/h15vrd7NY+e1sLoaEqFS7ay8SnNEWUF9DLJvqjB7HZj+FcKbya3g5+nLXnkTRn
jiC8OikDJBtEjKLC5o4g7x9dZ0ph4dT4DnJ0gd9qNAMmkHVrcwW7pRqnVZQcwePla90c/tz/RDWL
+IsmvEl/TD8gd1rXnBQOdEVb4DmRaS26eWZJOuOq+zjsXmkDyH6fCSa/q4Ld8btUlSdiESR1Lyeg
xmAoS+7u9aUGqu/2Wd7K6upPfhM5auBdMLsIhL8aVy+6oYZwwg7W9j5fU+rLnG1zZJd4bcbXTnfE
FtEPj2KuXoXxociqaWLytsd3pj5YsF1Z5lPhJiwoMHNTl4GDgrLJIXdxQwRl0V4Vy88rWbABkfVa
t+WUTP+Gt7QisH8HOjl5FkyJRoHeqgYKMk721Fc3vbeNzUtiRGVRVLEE/JVcvQw/A0T1jQXeIvpZ
itV7vJcMxH0QoT2Nw9tMKem6MHwcCYZM8cY7x8RJKh88pAJDLA6gxTxm/cciEldD14dTgpDsUCM0
OH+pbU669eIQLve/Rjoa5rIvbV4gTQz2MBzIyvhc4bZziPenVgE5osy7OCk/MmE2EX42/XReAx3G
5G9e6THexlyBAWGzf9XSCco+/HG/IdH6EBR1PogFr0StP96PsTfVnmVCnQ6aTpUgLnBdGr3lK8Ai
qsZD8oWB0GF9Vyb/LFVWy198mtUF265aqhSIEPrhBxgJddDXRBd5ArjwoNNOEhoUnHf8IRsL/beR
JJXxPLAhfKk/guquIn62g+xfbuuMQCJSCSHKs9bouGOzDZP60IHpqmrSB3T0/JlxDSsT8ass82wR
NcryAr8Jpj9vtyCuFV6QD6Bg0MMikXBVVtdHEoGOzXNf6Q1Q4/reaZuczA6xsMSTVqfXdVi24MNk
Fo3V9rjuT3F7O2bFLMbdBcZuxryDxU26ZGrvhbrqLCgolFySVHUma8MmI+k5rK5RC5Ysz93a7Rzv
jMpirC/GavllsZ0HqCoLzdfxHFpVIt1QI9DjsArJyWubMPpC1BLIYAYlGP5fnfzBDvDd5HiL1g5x
d4V1L1ZojzHtQSUeTNKOGr9E0Rl4MMJMk9jeDWU4021wJuWFv/KgZP24BIjrVQwxrSrJ7Nw9Sqqy
aeYfDml5XisT78rzIxRR0nBMCiyeNIFW3kYFTFfGP5VOePYlOfvuMNJqnyZDydgQyY6fWxuu/6HB
lY9ek0uqhIJCH4s63WLKd1jzrlVr8lqEGSSpfk/mEKCImQTCMpgOSts/Ny2+/55zbLQgxvFdjvYG
Z3ksEM3pDsNUW13TD10PmTGmPw5EKqqS2vg/hODg5r2TqScJAL7k3RHmgYUZpyuC5CuNRWejEANb
BmzR7WL3+rVuLiIFF5rUbT/Fpa25ITc8MxAmfAyPUd7Qedw3GggNb8UVucRf0+uQGz1te9JbpkoF
gkyiAIlzN97VtiOSNAE+irKQ/5w7jovnBZjBLSDpUpFto51w6dlOBx4EwjC+TGD4I4/rgWm3YTz0
r7eqEDxia+Yk55dIqR3H8KoAFzb1v2mIwtuZAY+VsVhyRjDw+VoavsEJoIDGaMUnuMZCYdbum72t
CMRBBn8qER85nrO7h/pyFuNWgJTHYDo3G/J2JsBgrSJNFHX+9zny6l/WQgHDR5AcEugm10tukOB7
Y6XLjcijx4gGXeY6r/QUDy9dzZ/fnY/FQQNJVry46/kQ/Pcqii0COmptmqbbsLWdNtfhrtm+8fnN
/bjIRaMsF+I7El+wIpUdeititntmLGZXukEjjLsVAx6Sl+yNM5nzYeyRt9wPPZPjaleqY4gr+nMe
LPGkGNcyYf5RI+jEBrXk1c79efd5a9c/wpQsLT2KqWhPfubRU900rvcF1WDgMlGfEfxT65aMD12/
HdARdtt69MqzAlhQU2t4Gr2NJhCHjLUwivm4arCgXpnfcKExwhDjsCneceZAS6ktCNEegqnbRGN4
oFB5BLeAuZFb0VAdVFGjEX3OQN/snJA5Fr4SSZ0S6qM8TDWeCU2V6HCBNBXa49MimQ9Yks9pHujK
lyGQx05l+Wj8ch79sqdxfLX5TlfwEAAQLsZk2h/zWoUAfqDSEFONnURbJP6hlNwNXXSsHPnyO8uh
gdPtZZwPM16BcgGntDssSlS454Hun/n09zgXjsRMQs6BsOA9Z0KUTzENib9ETQEENskX1wZCK5qz
ZLw5wTVcAG3+ZyZxcMz5BvobQGPJKJ2DiepbpkO9rbZ+xiHxcfLg+zTdmowjt2+xB49K9aFr4j2X
0tsO7DPfvQd/kas8Nr8uBr9esZq4kGj89EUju4LMiN5GTYBkR85Z4elU+wQ56qiOWBmjer8b6IIj
WcSrtZCR2YB6i04yGZWn7+YvQN9L28u0+KrkA9qiZcb4D8mbsjG0zD2LEsHg+evIMQV081POh4ey
gY4OgdxdD05bowRLUTk2rtgqIDUs0mOT9x94JQH8tj/WcIDMGU31HzqzCEyFzhIR0y+X+oo9/VZ+
QlNPImQhcha+Vt7cf0a6qZW7m70eJWlCDqnx9Ka3FgDvbzavBCxQl/ZOGd7oKjLIVLTzoCcEIHdF
8CnqlpXLOg5kYpWkJkve28LbxNYRUzD1Vt/gl+tp7bdQ1VQPpp5p5M17gAczsRqi6kdvoH8ji9Q3
5+RDWqHBCRMIAyZOu65t9LcIfHW/pUNwkzjL3M6WWqzsq0DM3KeC0+yf+ikS0tIn8Tg9BxPzz9kY
GSYkKPvZsLmt1JJzAWtT1sXAVc3Ct+FrAHdzybMGisswZkhA1sxOOvCPV4zQzG40hCT33ccccy19
7nLWluZxbeQAuYEWZD9wjwTY4YXfBgStxRgUFKJWI83yaNsqcMeGNtKpViT1BbIeVeS81863+XMq
GLHzaOvu+0wiciNRvNTdQAnl9O04vWzCOLNYanN1+zDijqB3zEoXAKAPnXhF2mri9xx0ndXfjhRZ
3jsWI2EdMnuufBtzhLZ9/iHYcEHv5z/VziBjJqzuasaonfbcUvwTHwKqN/PLBJMFZx1/eF/IhjNi
y7KHu2Q3O9f+I2tgtL1Uwi98CggWANtxsWx1/HjujR1aGtQfh3HoQ3vX8K7Rx/9LCROS/sNiDcGt
DLiWoHkU2Ei3mQs8gUQ2pNq4CslziFfrBhfTUO7mpO4hCDnokaft2K3zqSqnPshnwMZBIf8R2a5r
Mg1U3f47jpcSTVBynPjDpwAeLnnLcEZbhU4FFK5pydhO/00KXip5XZJPpypKJXtl7dobA588Tudv
IuvoozzMYXwbiZWe0Vb9wcYPD02z9+6kMJWOWRhp7ZAly+coyuBYeFkRmwjFPRs9H/S46pHS3z6+
AO2ojvORnIx36R3kaDhEiSfFaG09fCc1b2jNgLJJL8MrzQOmA5D3tAVtMjonb5TMaDdFore/Gn/2
ZU0rvw3piahkkPIHhruVt+ur/KjmDrvGRBmklBejnfscOeQyk9/WMABy2KZB0QSh32cgNqU/1A1R
AmgL97X8+491zsi92TDJaP874AVacRFkv8dEKVWKEvKkNXucUeIwGAj5xvEJpDiIFSyP2F9EZOBJ
Jt6lvE8QFXKwKpkfPKMDnKO3OZy3XOSynKSivjf+BYpCpimSFHcqoOZ+jXzdj1VN+die4QMWfcRJ
JVhSpgiwM7w6AVObXHEZEgd1+bItNSK4DfkD7t8C5xtdKEe48meXu7k9nlo/YZwsfZSCDBqiiv63
YFESMNk6Oqr6leUoOZk9TL5SENdtCe0FfCGQw1lo87pbbhynKNDSfW/fNm3s10M/u69HXI8tjJd5
uApx86gJS5F+3l+A8mGvzf+ZcYHL6x6PtBepibjEYZMpgVLaE5lbaK9ZR4Attd+xNKa8avaG5M/k
3Z+oDSI/g+5lZ6xm3C1+axD/WGxI7poUiwKb57paSWvni32aLrdXAcvtT6LK4gv0Dmel91kBpMeo
AWA4gEJTXyCu5ZPheVudcj4SUlQodmlB77HGoDgL+7fHLKhuSUT2BYaDuAa3d64zl0yi1eaVQrAE
rQyPIYqH1tnryWgKkF8pjShVVoQY8XPcGZUie7EOsxBlkYIsgDlaAkKQNlvINCO+7BCigXk/cqib
Hgx/GrdEKU7PFMqmIyoCLcOs8RU2b2U1Zj3r61AAcbw+s2Aj7npgslSeCtH7EjWFVD8oBJpkuwsj
l1FXh/bsyDfpgByUhswx2UkHtFNTFT030BhtmIW0CdWaaaZ2ErkzBlRidr0RWBVfrtGXyze52jDS
eC0ZedJYhQZ3GGwnyrH+C6BaTPfgRZjegaQ3JLluFZOp1pQPrvFSHrOC1bcJ8XuOy2J/a+jxIiw3
96VUknFRPNo2NB9S5P7krsT5CXPuBy4/dwFnVdfBFx5FB7ZlzCLZ0rOVWWzGLrNeQAN7MOt0mNW+
cnI3H9kxj8Nhh3izjWc15UF6cB5aLpEQUejBUCCCAMmeB03dIBZb00gJYEo/ywklm7XfwYLMw+wf
reRJZ7JdRJJVQPwDwsadXvonBE4/D0GgApXK/Fe1V0vLPcmIwMkAFxzmnrfGkOonKIJQs7ajHvQK
TYwY3YUmdbtjkRgLmehePHTyh5087oPziWnrPydW8OF1V5hcSEJRUWhfLWWS1VbWpndi+oZtZwhN
J702KRWC6GSAz2OLcKD1bgIs4e/n/L/uT6qTycz5rdrStyk5hDLGJ92tO36JDonwC6ZK/8zUsZF/
4PfHwYuHYYk8R0IKpj+zSKakdmjWh3cCiQWctwQE4YiFb70rausJ/xfLEJqJ2G6j9si82sngO3I/
zN8plO+LlC4/VNJR0pc917yuYPb5rh8DDSvYDBrTZg9Gtktg4MteAthdUbEtCiom5WrtRCUJsE7q
9q5DiBaCz0561+ySwQ8crYWFuG24JdvU8mdyQqgmy7fP2symYtSupeMGiZuCvH11f2Y08tjDflB5
DwerKcosEe2cOg5Ui842zxgetj9oF+ZTBoNZGvP55OwB90Sc7u+O61EOxxX443/dIhIuzX3Fhi46
lCLE2Q/AxD15L5w7v+ic4GEXF9LhTh415g3Nn7Gb/ExdwpxLmI0U5eQM4Z8dLgoskkBBp576lqmq
z2bqQP/rUYmVGCrEFxjfEQ+amGsRBXYTUtMUFKVlFcyICMsowRUTzs3JN30xbcJMOn2/lo10jQm4
207kMfoTdXKAotkBGoGrHrfjQxtKrlHZYFBwt6BAXDG8lPqqks0rUiFkMC0Sm6WaFLCS8aIPryar
5B6NbFrQwp6wDbFp5tChP0y+16q2C3uiah5TwX19p0aqknoPK9oGZGga/4kWbHftO7bFJqV4nqRC
MGHyBoA2wXghF3MtoNisulI6y5Zm68lHmy7dkIlISDl+xrFsoD3Q782R3EZwcYoyAhHJxk5n3b1/
SMfqiUR92y8akssDKZ2lm8qtm0aPncZKhL9raNk2WwD5XaSOGhZeOYm80JkTfhO8+ou28Fj8G6DD
K0G/8DZEvZoF9xBIgDHBiPgn3CfvzDjlQSoAzf6Xyvi6Gkbd/o1pV869x1oX0U8O78PwQrkegOLZ
ifZh+MGYL73IVRbKqXawD/aSKzgJNM8Dt+CYFLlMM3xdpzW5VfNKppcdzOMBQn0UNK1GAHC3dbOo
zFwMFvc6tFBnP35Y1wpTCuaI1Wn4B7AxusrLT2PDyh6EGaw/6fHhwZpRuwOVq0QYwmP/QtdTQxTL
NK3ru+HenvOe1FcJsS+R/cqXu2XW4GfI88+9CaTDPfR8Tbz4rTD9BV/nA2/r3mu0Yb5mZixscz6I
QjkzmAvCUyMD42TOS3Wjnss6xW27QntHga8ay7YsNDq0IkrwmczpkkCKWlbfmi9M2Zn0qOt7Ijqm
r+jq1Rv5V04yUBLq0iqo9XG0Vdd21YgYi5AP8mv15KJGNKSRnK9K4knJLhsdQ6UruiHGjQ+Cwp/P
hVoIN1S13oJdE7E+XI7ntRwc2bNkWTeAmEl7ODvf3RnC1OqKUu0s59NqgEc9lN0ab5DlNVfw95bw
7YWpVxAsWHUegtIwHusiaMRrsYsmMLGOTIci0gEOK9FkLjHvUMVCrOJRBmitcE2CEZWT+j94Khhv
q5L4NHIvsmaQsPB7NrxbPlV1WHZ+RtWqaM0M6tLkegwgtYZ4I4Zhfox/HHP6zFOiEjLhYfSkk/JF
0DigFQraBbOBtgtK2q60EHz8SsLcNuovUrMphgKVlQOS6uiJAUaHGozC0gepQhaIgCoaKHRMboMr
fs2jLCZE2lyvQTjfHnN5Br3K8cWn588KABkluVmOFA4BWM56BVmEZogzBLhvhSSOCdOXuOb19NlP
0dKWD71b3ArTGwUFLwIFeGExGFNWf/PhIYvloWwPbY+/t9JMvJQtJT4W880JE3iL9lgTM1AEpI09
BFwUVvHifmyUcUbBOvYo71zwTJMeh3d0Fn63TwHofM6heImwtovUy0ZUT/MqQiP0TZnT0Hn8SBNb
Trj9SI7Y1DNI7F/2wgr0yB+z4IGaUvCN0hmtUpfnAeKp5tCruaJ2nAgeIR3LVeUv1pCKxy80R4Oo
ZRDAQzSY7q0AwbVFWLwrPnrQBSUu9uGtU1ThYSL+S9QHbUka2YwA6IZmLMNjU+2X70ygIy1CPN70
9R+f62eGa/zAEdr6iZHBYm+590k9UMNR3CQhPOj40+C7nZnETrUjg7NE4U8wuHAnpckCH7EV+eeL
Dd1kRyM3Z88IEIfKKj9r9lE3GQj21D8R1+YAAWVbHDr1S3IVn0l/pMzyHelwFNV8eR5Bt1U0w3Ft
CUQSELx+bwQtUlTHXf6o5L0tURjIV6On4CZHtQzrb9JlJkiZmPkskqqIB68EXvmPCzA6AQrruu4a
3AglC8eiwhsz/cIOBOmhkc1In1hVwRbchy8ZeNk6YPCj9IaYlMY5dJGId1YB6MSFLJjePZViX0FB
C1URM8LzYDvAMrskwqrUgr9qK9pcMgs2mmlKzUtQrkLEdbb2bhkrhpzNA0O/t5J4U6FSwtqsvxqb
rPeKbiZgEwmwPQDPj5+w266FlCMfxuqNSZc+lOYVvOgGsRXEPvFp9kql/tOiV+ni1xLy8Wpka+ax
0DXmdMXndGLpFj7unpY5DB5bCi1pWTP6DyX1056aav2NIdvgiWySO47K9WOZaTTppuVWic10oXtT
xookmOK92O15VUKZ0RY7C/aYuQbOUFCONjqeXc6kItS4tXXpND/rprr69KuEun3ppHtOjpTv4Arb
cG7i8RXfgbEllOAhs6D/VxHCS3Vz3dt7D3v0hgEvNyBFCNL506YZaXr0CJx2g3yxh9rAFNYMpmgQ
+70HSYw+v7GCLzj0yPMT7liefNUb5OquLzYKYvYNYHiflhR8qfeuGx9VOOzRSVo46PxIZzzGPlfe
mj2V5PruKHTJOae5i87Gn3eFzrSMZOz14YkYlWVv3FFGCcg8cKb2MUurCVsO5TBWwKPqn2TFz92C
yLin2cjQyLHmx6lu1bGz6nXWRI8fafaK5jyLKHBCYczTyFowlkLAoQafltWaBeFxVXcXQ+lxej+Y
mPQlwudxy04DcizLsZ7RFKvr5auZzzSD3/widIF8Qifq2pjAMvFkBuYWBfY+vxGabBuqbFh2EEjV
D41g2g7BeGjb3uCGy3fYAC1qTYE1ufB8z9CjDDkifoS4yJEq06t8ykmLXTCx6jBmemZUZZw0+9cJ
NKcv1X37FVLMCPgtznDmsh+srbh0R/8l9gxdV/Jwa7d9jM2NaCBjNGQVlcqZ1bfMDWYzPCKgr/UL
UqnwcbIUauBf4MHsSF8HcJYlBluri4ZuSr6FuWKowFnMRCyWVpwnxouIMAr3xE0AdoMSQjivmqFo
lZN0b8cFVk+IKxzCet34ZEEUIiiMSHKINN1qvrD3/BayvaK5DC9fZFXV1ozMc2MxIws7K51w0RHW
p7tCIlfbiE6X2VZoOAkpKe8bhpdbmFsxNDdk2W5ejxlXUZ5cCB8jW6k31h/Zq97f1DURzTzPxXta
DRKT0mkDPQmBEmvTkl3XM17TfyhRG9xhnNy4mdqH2UdhRz2E/iTGkEsLv++1RQoxONlm85e/v0Un
2ckquiOqx/spx1/mbzumAto2sHncitZEOl1iC3Gd4BXg0B5OaWDM237bm3rwcdrCbRoXQ0LCsDcm
XncA+CMuvic1GA9moh2hRWGt3IH1hsCLpTQ1T48qiN2aHTPBEBNfnXNc5YyyHuVRGWmNIfGDGGbJ
saW+87w52k6EpHWQueSNt3Nk5KqYLU9uZVvfIMG3kzhm38A2svluWoptIhoVDckt59FGq3ioHwdG
x08ePw3rlSRpjtU0Lvt9hliQnKHwyh06rUb/qWvMy3WtCPVj+l95lIYcPJwSVfcv9sL9z5XIjY7v
YdVareT7lAT7DqCYeZP8UGN1C2+23Bmh37UMUkhpwpN4SVlW0Sv6Ii11gD9/OeuDZttfL11b0z57
oPX7Eml+FUyJkE3QNi8bgn4jHI0t8t46CYsHpeejAgLzyOoUZf91CSL94PSOOTtXLKePrYrUnR1s
AL1Yce+XLhq9zx82CoYlwrvN3wJKL8zdMcYcWUCPYUsAE6Gn89S/+aWnn0NtK5B2FAitaok1/6B6
kPcpVU4M+H+xaUQ+0W1Y4XxIrnUQbfrtbRFi5J1KN32IA752+lI64lj+7+SUosoHXI5ajXnE9e6j
el2OcHNeeekIqfhAMS6TDhFz8IXQYIun+CoOir4RodReGYGSfDGA5RaJrAM6Kb90ZLKgW+6eR9Pj
si1wSqQnkaynJyQsU+natkgqWa1mf5sd2efZ4eehWVL8QlT3qtohLJi0xQfMp0yOqtgK/E4ialqO
MnymgKGPPZeNQKL9rLTTBTKL1t4aDZllOtcLYL8lWssbC5JUGyy/Ysm0Yzxm6upn8heldNBHKuvC
/EzX7VDU0Yle5kdeDmCjh7R6DJOdUagJVbsujQrGT9orHAF4V8ePvtOoUDkPgoP3CopxPKW1aIt5
QllCFjq5CCA2QNBsYeuUe2NJMXVf6I34M43UR4L/icP91VU2D/bTUiY8nqz2ptdNIVghbaVbLllE
D6iCb2uExPHfNv8jwcJEgJ0itj+3rvN6GeInZn0dBpFIru4DRQbpfQNSumststmpKziwz9lvgkn2
rgrzui5M7Go4RSZe7WoFevHcnIx3KCmxfS5LCNw3ngsR/Qy3vJ4y0m6JK5DTEO7xL+xK6psp1rEF
CP3rGCAcIN++RKaN8QzKf/4lx27OGJlCoLgpcEA6RgZ23CUSn5rEmI2GjSjebAhAS9OS4yD93yKJ
274MySMTf6FlGUWe3o+saCRQiZJpPDjxHmE8vNLUWPUYxfZyZi4ZLzkVifZZEisKfHOTjCOq30ZX
kblDKVHbA9PAh3CiVQQpdljD35NnLHtAwbs7FAfGvNs3I7vF1CP7M+L+v6PI6L9ymuBLZ+7Qxdc6
naqRGYaX0zIF9uu9oij582lBksuaVKCSMj+RQiF62FlBSteb9neOKYaiLqjUom054ST0yUZ9w3Ks
VCkHqZ8SQDR9nYes9Bo3rT8CoDwoTzSe5o+2Re1jT5W+fxC3/bMkrNdE8Fu4DblhgeCpnKwRhgzC
gOP3KKcz4B9fOlIGjCmuhzHnDsA6kd2QemvVpsVXSC45+Nn/XR0EExt4onsuTqI1//7EoJz4Tl1n
1S40XB71LtELlrOupAQcEi2IB7vgGtg8XzPQIJY9qbl57iHuSGJhDtXd21uuPZbEBUmigZSoHEjP
+PSXj0tBJ8hgMrouBJEVa5r9yBu1m/7uYKlvcos4DF1Yx65E3W5tZAaMIWv06wmJl9f5i2CHghWe
fdq5Wsbo5Uxk8n7qX9XUzYOAyV9RD+cTfnucZhqXELHW/7g9DbqJ20+QXMpHgaZIvLzUDKAkKbzp
6e5KTEI+Il7Rf/2LLz2LxIlnenVhA6b65L3dlqCLFyl44qU4LabkVPrhZ9xpS0HJMibIMV7fmAsH
RCwIlNce1mJpkfJbGUE1IQl4cxYto1d0VnvcnpM0dbClhXRkQfeztsYD54ke4opWjARE0ueV7KYy
7hAlxLJtfTmk+Rq6gk1Rz1yQOIXCdntOWuXS9CZJXKS/OaPOMsdNd9L4uTW1l+Wm5XkM7/TY8RL0
rHYsBi/Z66uDaCTXsLTFh3SMfBCTNdTUJ0cFMRqXmMSE7alABXgd1f3MfBAGH+qiajU0jh5ybRj1
nlxUUUo6hovakr9Vl96iNXRltKi4XNll8WLMUpW8sToXDjoK+dAGB7NVM/IQMpqFU7wqEeaWkl2m
gG3OYtaxlrBZDlb2QBDEBacmSont+WS0jSerjTDlIdO6AtJdGpnYNTY+CMi5cBDzBK2yIW5z/hRH
Ad0GNU/8mqftfiX7//Rk+0JvUAxNUEpivYVpCvf6WfihjIHpg8npb5pxak899DCg6UxOrO1q29Zd
sRGb3BHac510Yp8u27iOt2LEgNhX/LtM6jKVFEYoy8318BI/1Eqdd5UxlpA1HzaB7/C12Zn6o22X
PrEU2Az0kzYgyB9+MOB17SE/z45dN7f9IWSPwuXdhHR5BGbMvx43SnPYQgaEGVSspEoVOgbLJHay
ypGdr//cJWRQztHggRdaE4g6oTerTC7jEIeNrRTOseL6MVRyFsKix1aMvuXeHBfvMgbalOojN1Yx
1Feodu02nzqDEvYqtCk4/XXvnWqBeqPYadlbhW/EI9rWRjJTp2RRh1HAeF06M3r3H/la4G0q5/2h
hdbrhJHtcIMsOrQi97G4tJMqqlQ/otb2Y3Sp+y8MV6W80HtKMyGWV9V7wes0TbEeF4AZaQDdg15T
AcgS5JMID6pkdJSOOsBHBoBKuIznd25R078TdNBEn/esB6MTptRx135zrZt6FLSOcz/bavFpeS/j
5r9UPb7WZH8qrWF5TcTYyWpgOIRRncivwEvvSNTKg/pfbmF9hfI095XxKTOX7rf05pE1T5GnaPSl
7j+K3k2M2uGrn/4FG6hdHY7qh6ea4fHK1TsYi1l0OYhU0VjE2fOi7Mb34qmtVa9IgWMdV/P1JMaM
bigqL5F7oCYO4TFnGNd3yY2FiaH18W8NhVKKlHtjFfkmzrwwN83X9tt8YTt32VQRbcpxmEMAZuEs
oiuHDuxzGh5F6zzXty/NyZwHEvBiNURxmBd/RC4udSqwxjI1hNs0zanQbR0KunK1VfGLD6Y1xfos
AukS4nHcsIle2fR3iWdeTTFdeRtsHxp9Ex4YGbKdO09GE8SbCrg/zae6APU+A+FwCQI+/rz9nEia
0NNihtOjU8dRExp8Puv9lYJAHDqpicJzg5Yy1ek/m2dpVGNwJ8tDEzbLubrriLN/QlJKDKuUMXxi
i2yDlD5IeAXCcT6n42fyvttLeoU0iIfq8kg5fUAEES8vKOsVbaOeAYe64luyR5AfBfTH+IFOS8SR
mY3lLMIMdQbyyOqW7i/qxYyHswqesAx9bZzRol7+oaBPtNPZ1KFMOPVlOUFqcdtgiEIAyG2qwTXZ
gNt9a+92IVyDElBEP1qNXlt8UfCc5vO5zWlXs28i0Jpy+4r10w9gzmUvhBMPYcu2wTHY5Bcwdlmq
+1Z58zXcFWd4Up41LZ7Z//B84K9QrujVFEqy+I/+LFNmNpK3dyhbcDoxr2pvFJN8F9YeSbSw3Mgx
wDxpB2FKmqV718CoET02awikxeByT5PLD1um1AtGYk0ZWRaUQ+pUQvR6hGdvCVqvb0EzJFk+1dBP
IsZUgOv0ahxrgMm9ayGU2omVy6vFiQ6bWPBzwGHY4SKS3SQT8KVwm/M/hJZdENgszbnqDN9Bqd+w
1tjuRbSnq8RPEGuVIuPJkAj3GxpZn/xWURI+q4rKuErVjLLLQ4pcsWKdtm+wO0dNYkvkV1MBdqH6
jeNMR6GBOqHk5XR1pxLiwLOUYr/pPLYx5J68pFs8jmZyy/XZCcbMWqU2VFGQdgC+SZxTLYmMDjR4
G5K9LxHgNYZMb/LUneyQgZsGnVMLtiYCmdEmlvkbaPnbkL6bg4E/mfYmX36Fto/l7Pa3px9Q3z6f
Mdia/CflsnZ2HJb/5+TJ+n11rqw0muS+pfRp8cYCOq5Yp8kyKBWEENGO+WD+VE5Vt/Y3FYtq/eWy
8idNAKSOtRdFTgQNXY6ne3l8l7qOxmWYzHyw0dfexHpZxcwcgTADE/x9teaMBjwCU5KevN6hn4f/
no+abn9DJhKceuUXjOaKatEc82YZBFZAPnHLKbDzixadK6k1PynD/ShWF+g2R+ud3sp/v5v0Jd6S
AyYL1b39kEhnBWyk9K0eBQ5Mt584i6Y4g62V1ZnCaUXQa7chwHxLgA2ur3SKU/K9LBU4TJZ06F6b
/EK0UtXvyfAekhxqewmKcd/6uzWZlz0t9utymXWQAVnRXxIJrM30qIJkNexI8Gq8m8gUNKK9d9/e
VjO6DIP1u9JQMoYYvhh6Oip4nPALGNpFmZpXln1t24cuG8y5u5/U3LR7cQqTfTxIoY/W5gbFVy6C
phHvEDUVfmsO/H453eefMQvQNBRtCKIX4NQzeZaKETsbDngYD4TKiKuuhjVggPN44CDGRAhZUdOS
NZ+ET/FIQIlE98tIx5uW476kiIupi/ybdnbXT+JvQ/YpjWfzxeRTCL+v2cT8c1CZOxwEJpLoX7zq
54TtJtlEcEPIaTUm5r3UCaCPNINx7bOXBk5Sc9U67d/YvO7R8UgZ36t46jBgBa9z4bryyPi5FjbA
YtWB9JHuwpZd+eryptTs0ReIp60Qgb25jMbWZQ0hJX2oJReBFQPiNwvW/kPZFt634h6qNxHYJKAz
hPU5hKNT8TTjj/7iReNZuOkZR1thAI4e/xmmYQAztviWRXICMzpFpoIis7n0J8UEYstpwVHyECxS
6dbY5a0PFJU3+tk0tIt2dPvaXhIlHD1fB1ymjKD2n9CP65PDVGdIeIAXY7kFR/qfzcUCe7KQNEe1
PwYjQ1kuduDZYVjYBRrAh8XW8c2Kwt1mUvaQPlqnI0FC8jaVC3elUnhCM2pxxLyDurjeDeoK/aT0
7mdoGlDeBksbKgaOSQB1NDALXY4vNVfgEAg4gSsMD8aHKewCv7R4WjBgS4U7XW+lkhWzvDl7tw2X
V16b7x3ekuVoHsyJOQ9by2OZVMmsdy9ydDaUV46QEpxC/JEkuf4DvLKvfThMEWDxqyskHRo70E+R
kMF2d+ccWfQJWTDPeftrgWy5kOGEPELqWyd+osB/xGWRF/EoehI+je1kTIWrxETE1ci77MQl7Vjb
OpgxfsU6WQd1jiGdT0ZipCPoAlVOfeFkJEe1Ww3wmLsFWf6zTFF3ecYY3zImSFXRL8XU9kTht2nf
Ap4SPtL57yTLe4IGbqGyUZ0WGh05EoQHvCb8edc0jN3KNTdfFfImOTUIJGVx5JAW5GHFkduIgGnX
CxY+P4gbUQZCSd+0hL1LEMISLHEDJGqo8/Kln9GLcPAd2Yey51tbrJA4T6SXcTYnb55kKAjjz4tS
BxfVODCr35aTHgbXnCSRj9yrP2tK/r7pWsWjCoMkAxgxhw6foJJImzi9qBNeTLLpBhGI4KN2sHBV
lQH/Go42eW8BPshHP1lN7+oEvppWgdoGpYFjYYbWPGJixPlx2KnueFeg0zM/wo/nU4rVZH6navoQ
0DyGsOEN3RiEHcNRbvE5beKg4zD7uWH8gxQ+iGPVWklfbW6Il2tOAaizL2+2YRWqnyg7nuUV/0hm
75T6udMpl5XseLIoodOOTNPQoX+ZVC/e98iqqPaH8+UO7D5G4BYB/4QYdgn3p1z0zaSmxdK3DUvU
/iYa2GMrw3Kq1asRHunn4RUeJ8T67xu87J/LLj1TI16WXNBhzmoWdbMXq/drvPGx37dYx3gA1kpB
Z2of5henhT57+q7Dju+Wj3XJ/pnl1dVPE5ehypUT3sgw5SichUm6pJGfI/XeQT6nH3tCgtpjtkJK
KobORZ5hoCr8Zu1r8Ovik43zlndZxwPPfOGxTql+vlH7MJ4d1tK0lCyDPFww5s1NcO5Pn3Sl8/XP
Sy/YmoGhIv32+4NWKl1ZvUqJW+CuH4cXe+sMLa6lVY8sZGiDd/mC4Ys8X6mA+xCi4+j7f9RWlUIh
huyF8EGoI7Itsqyo8q+udk9dBZr6Mxn5NdZ/7HRFs5JjSmdWoqErim9nxAMfaJXvwtPUBCMp/g6D
EO2Qm3l9Nx2s0dgrtFMyChURbis15BFjQ/wSTsPfYHBHRR3LUrxMkGCAW+61JMw2QidOCD/2De7V
Bz9dC/eQEKl1P6+NXwS/DJleIQZ7o6Yc/W2yuIQaZ9E9xD48grYIXVavvg0x2I50ABJNjLmJCblU
kEnO/eV2008MqvWSSBaoNoTmgpvnmM2NyQs0j3LGsTNQV/BcigPFK9gk1ezvslQmxCesP0dfvABA
AaMIREQW6Qlty2IMdzDmcrr38IUs4yESXJq7DnNQ+JHNT6jS5c5vbgAMC1bmnQ8rWNuYsPCTxhno
TufFH7KSGXKgAFHrTJx7ZEYwEyNoLSj2JeLT0lRUTeM3Z58qj7WcxstStXElz40aUoXaSnxRxtul
NTkkh5Y5ggVcSQmveczGczexo9SMSr1isxULX5IMtCqTLJiPG4aNwos7JeG/dzu2Xy3bZBYHdYVU
QHqNZ2zcP3Vt+/fPHdRj+eYAI/3Ci+uSna+7S1jo1jS2vtLAwRiRb8oHoUpfTWqgQGH+u9tksluy
ieGWNy+bzKgoLxsrdX29uUwqshzMC7rTOmb0CYbvlQe8BdkeiKvR/EIGWMaTVu+sc71S71Q3dx0Q
l3LJDRzmorzh/i7NXWBXVkU7b6YhCkpIyRRATOeQjR+LC4X4ihQ+ppqXr28wixGd2MYUssuZl60U
IiSgrH+4ttyo9UFBzY4oh/JBmI0l5kcA4z4yCwXTv4XSzqfZHLLjKP/ZzUyaEZwCCGLR0wCb6EXY
TiRId1kfPxxF/LTCm73KGNoG0zpcOt2R8M+su3+Q8huJXIUandlM5Jn4GHFcR7ejT6b4PKzWIhKU
DDEv7r0d303vDdaTAIwSRsXddeqLbcJf3fHL5GKrpe0UYJuegXPz7WPXaOJvDBgYXv/TM26oiP+f
51eY+8BK5gwcRt9fSDD5MFcUcZ+a2SgErFReSq36RZ01kN8f0kAUJcwH+S/Yopl+RVl/PJVk0e77
JjIYnSQvFdMRaDN4wb6nMw+AFye86WDmLGknGJRvWl+ZM7R1thTNOzfT7OUCfwExwWKc6EZJ8G2I
pqNTtcTJT1uPn5QJNmFsRAdaHWuYT97Hs2WbREgC1af2cld7Sx+iElLBmXIE7uKHnswku0/6nAOg
W0FnMojhj3plcoZsvEjGtpPGR0FubT7kgQafzya0XBlt0qnJsv1RtCqGrK2+G9Zoq0C2WiydYvGW
uL6pOeeiRALANnMbrxZfjqVWkxzX6eWD+j85Y8K04bk4GcmQkj3Vo4gsDcQ0tYAEzg1Hs69FmdGv
HdvK1S5+xJB3SqxllPvLx6Vg8UbsKwm2/SC6O7+6sMpqQzcn47gObjWNU9ukzymf/mH7GI8jbEwk
x73UiWbqB9bKrTWqJ8YuFYo2MSlRugBmgd+U6S5NWSMu/cesPFoMmhT/FD76/znIwzM3j/Y3q883
huwc3UaC7vUYzQrGPPMIeUk2astF+nAIfVEMwk4u4tRxtbCIXjngbgJssnENFlwYeVbzyj018lbb
Ij7pVj6y2JKco15UwtXNcm9M8mazu2Ma/z1uEEbAi2k+m7GMbHPOT4dhj35Mm5EaKl3X+Scdxo5q
GTlxsOviabZ6GasEMBWbdOgf7tRHT82QBbhEsAHD8Wt2EcXmGR6YO5tHJ/TWVR2Yqf1TrHJjIIXD
pWzgOwhCIVGermOGJs4FK2btUn3qVBQTAwVIkUtI57RFkueYktB7+gk4GyIgiKmNKeJMF6YMEeDA
U/93gFtvHD31FpAMXWcqXGism4wA7EZ6X2NQwD40tivtSbq2teQj+n6V74n/5g/J/IkYEhuDxN3q
80E9G2Bl/4yF+HUg+FTYRJkQxsf6tbAVxm0Qx88B1xGyNVqZRlH3rbfQiK2U2P9zE38HrYEzcK0L
gysJ4X3oMcTVGmlkrilF4Drop1hDficoJC3CWnPj3NM0X6+/Tw4jvXgRH+0bO3+NIn/ogLNAF5iX
iF6unaukUHqFWG7SB3u+MbGFJiuaHSHQ0aWuvG2xYz5bpBbe9EoFaoSB6UWzTC2AYL4xdUInmj9o
PFXOFZHjOHSh70Ea2cQIzSs4o8pR4+VB5h0rDKVR2mtr1urqDluthTY8iLV9HTcgeZnTQbLGRnEv
Sc1Euzxb0Wqyll1K7terfR/75ePa6JBUUOpuQ2k1zngECJWSoERkM849G9TFoinIzMJbl78XBp+c
nxBX/8V+S9nyFFaYJATVR9lzi59Avkupt3U36IGS3UbQnCI5fb3hQe/2SW99fslvCLxTCBrMi0KV
x7YUUPSEAz9J/rtMlzRTCUK8t0/+DO4qgePhspNY4RqJotjd00ow+GIwfQPJSKic3+KQpm3c3T4u
x7iAxJUaSSOZDg3rpsA1Jn7Vy2l/N5dgsL8bCV1H4dQSRLdU7c82h+OcabKXct0exAxRlT/3u/Fu
4BzNXCMXFpzJA33cEr0bggY19qmfuWn+Azh6pdmowNIfe7CIUqn0OzIkwD92MO6S6Y6ux258lBQT
GSzd3DRh7KOgwCb1FQuGsUnyZ5qqvg8gfeCazhhVlIJ0Fgn4sRb0Y6KXfV6j44IwVpsTD2N/C30Y
WtgMEaPE8joo+mgWIcA1T4hD1Ie12/z2xvleuLTM+VDNMpt6zMa4cPYoEyZyXWNNn8Bw10+o4p4Q
Fz0oES9XhHnE8+NE5yUfUzVjhppkdNT2mSFsMRUlmxv/v2tfTonK66tiHwHeRfWWjCnvlS8AvHme
vTWfANceCiIr0OTYf70gsdUJtnCsIaz78qzYXmT2HmJh1PYN13ny+MwboZVPpqKJ7Z9AQ8m7YJ4L
IlcBCvkG4VmtY48tuFn0mNYsX7nyfil/kFDMCasQKcosh76bnshLSNcOSX5tKEEgG57Dm6l1vUor
HCoFgbFkM/o+/4Kr3VqUeVjOqpkz+J4R//fYIlbKGHhSv14HgDaWgO4uQhneYVkl8CVbvY6rAgMy
RciedpLOOVXOWMB90yHsHUCHK5AAur26sQ/TQ8YN9V9ZV62vPMI3DPYBgbQHAiuHJfWD2EJTJcSR
E2P9WE2VOyafdRzCenxbyhaPVLUxV4SlArdJeBzsHrH7isZkRcAqLKsMgxliRisk1HZPvqkSAdYM
lgYVxBm3GG4EG/Zqm0PuR3DwcVJsiblkqyEOJrMJ//R/aDPDPpsZpsVffUFpdLLFJkgQ6AGu0gHP
jYQQUP+6m5V0WL28htxF/pEWQA+m22+waRxgjIv04kQMx51FdgaClQkUbEHjNfwd0M1qqA5cB/Mg
Q5+k7To6dvdi0u0CKlD/UO60dRU2Uqp3eKVSYAGzTcAnqv2gO4roqGseg+n5lC11Am8XLPyF9YNg
brGIKSe3F2ei8Bd1ezoLLZ3ocZ3zH2feAhPLbHS0R20i4LgCXiqfrI6G5aQmWxpetjyAiwwV+HII
CT9AcKjoCxXbmXUUpBmHjt63TVnx05XGEfjkqVlNZwB7UcskAzrV489mfMt5mjtSgKMoWiCKV4+5
7j1IQHxwK98lYnyFtDVBwISzWFtNbhVSowjS6cz5WYFeE7Ws8Y+xAkCiQeQpuPiRRFaD3+mW/z7K
w/UoyKvALCjxY7V7u5dPDBuvUJaoufi16B2GR7R2qigw+lYwQmiedfbxMf8AXbkw2GqzGrvLmSmp
vGwfoQO5b13CgG0Fh2OYNLQ39mDqq+Fz/s0Rhkp4PalieDJ447cn4UR7shev0VgjuSNrXnBbiNMN
5BXDUm0bGdz8ZZWvZsgfAzpaswU7Aye5DmQhd4uqdsRDdYOhSoyHBY5ZBcRE9DSRnpaNdJSKtbIn
k3U98XKeen0OG0wgmyfT5lkx/DpzdeGH0xRN4hlfJRe5HZXKUSvodFydxQ6UlOmuLl3MTCvELcUN
f6VL91wNB8NEX/Qy60YEdWwWNP9xAyxXAFqcix6lPZjWzlQO7DOXR7bC7ADOJ6O/O1Fx2t6egeOo
jH3qfXjkc93b+RCRkyPNb42c5SSQLHShRTsRGi8RBdlBCa5sipVUZVtXJOM7CMNEUBjo/CC4WqVL
OzmoGkO6jwBGhdp355HA8kQVQube3ejlBtR9GPZFn3+W3Q2h2Nqn/6EUM9Ixyday9xX+zz9PUtMe
dp3xY2nOvrUVW8K4vBzMjU4L8BkF6X+FMsKdk6Rmh+xMsgq7R1tnpWB5PAbjgmgAg2EhR0sFOuJd
I+RnITgmzKqnNXM0haf6vNLQiatGaO/1/5vq1uY9l2AN0kxltKct1vsAuXawd03sKu6PZMu7KMS5
6BDUWECJO9+4cIplXiGIhcArg/SQOf8tT3SFFW7xG13HyhEcJQzc3zugKjei/Y5cv0/bpJTo2Fe7
3zUr9+I5PGB5cmKKSVfp9TSSpLfQYG4L9RlgmkyM5fQnzJE2WV68q9tMgyH4N6t4v8k01CqMUwW/
fu4x+j3KsPbPfioqva1IppM+6uBDNv2VCHNRopTGml68DzdlQRhNGVsUmgKr1ZkhkSqIV0KY8yl+
a/s4CSmmbp2KaEVnQ2EqxC+WlkgeV993a0gykiKnTU9GBjt9WCiTMMfC1EzaM/dQkHPrb2Q5GsNR
Qqxes8oQSyq+wnecI2dCEGCPeV9c3VSsk1y4nNZGznP8FEjydAV8uKc7s895dZkAMW79tQZte+hH
jIrxQbHNjmE8iqj/dxXuKvlpuTx6s/CvV8orp1a8q+TgowAjaKBvnxv1vZcAGt5kDM0MpeJ8oj8s
bN36fHVVg8S9q4bqjKlrErPULsGPgq8Y5M32oPSvfRrAvYyitzQZxoXuzqJ8/3fFgDGxlZLbkUQY
NWS9z4maS1nV6pJl2a/xEuylVMX3nUQ7y2qro/0sWLGH3lqqCz/Ize6fs+kKSRXkD5xhTKnz3SCd
djwsF10Zf84hxS/OOiFz0v8VMz1cLe0gXjHG5yqgo1bXV9760rvZfVa3JYNAfrUc9iE4nvA7ekes
ZY1WTlkMBvyq3CoZSPF+2TeDnd6mOknkQcYtpLVVQ9mj0NNNylFtA9NLOxj2U346cSZL/HF1nQPu
6QdMtQQbAWcM19FM6oLARBDzE2Msp4L7rtxL4bmMS2Of6lBhLrSIfkesj2ziSzmTRWt13LtuEtMJ
TXp88fJxGQN8zcrra+XXfS+MWJj9o2ESSNycttiZG9pz7EbOK9TXkhf5P8UGW7+m6uWVHuUvSCuD
t40tXZ/ywfaRa8fSTr9qN/lWYYn7Jj0gUfHfJlBPBm1WZiXX87MkD5xA8/hYP6W161sirh09rfI+
2/nBipN5idVhMZbqhRcUC5gGBEJygFXrQo2atDAXQM8IDre9ZQeecnk/+85Fiyf/a2JGbIspmTLO
toZL0prtf3XoJSZ57u8fIpq6DEdFnY+l/3WvL+yQr2CxrmMllBRzD+V4Fk5VuPoC8xscX6ktj4gE
W2cr/a2ofUBk6AWQvYCcU/ArN8v/c2iMHUGsqq1GgBwrrGnOj+bE5VDID0tuTLFTf7o1RJ88nmh4
IS5uv6Er4SNkG/T6YZW6cuE+TpglnSvaTFHc8Z4fWlMk7isGM6gUB++aYq11T8hPmUj/aERBKG6N
BwUw8gyEihLO3iRBUBOI9c6jFY5jES26riILC7Ey8zZwEnVZi3ASgb2UNyswKceYKsXaNV2IU2jc
z2Ga2yM6KqLePThGPktyoQfBb47Ap+V4/OdcvYMYLSxks+hDDE5x8V7MxRCmqfTKAPaJzbkqofik
+0KjAXf8Cbm05RKIXGhIFUOn9TZf+nDFoYKDb7OY+b58AnQ1D3uUvqwXCBNjolgBIQWRN0Re5aiK
/g8osERmhspuqA+6pgFEvGhMkpcNUZI3IJ23bQOb4OIX6kwKSDTDVxWZ+2LRtO4pQhHN1Zxgm+5f
xRuAGRGcJqMu+csaqwCjQgVCCaxR+2CHK1LRF4kNV5iLjQZ3RJKHsAdBAP+JN9QiMTGq+BrW49UB
XF+ID92+RVzSd9W4GGhdjYfYTQPbi+Nkd3Dp+5kuCGbEWQkr6ZR7QghPKLWq+zCM/5dt3OosQhXJ
rTo5tjyhPWpKA1MeNwsy++dMt7gCkSP7mTpya/kAoKwC9HFn1mnTs4JfQ77/QA05YOV8hIMLgf2o
67NzE2gZ+DHm4hJDRiQd07VnQm91h4Odfkc7TWheSrQT0Uwli11Ditg5uPKUtsI62JSDAh07YqNq
0N1HyGQ3n2NxXnHLlIz0g+ImNbhudMEMq59Cg5J0QaPg9ATU49mQ3mksiju8qWfjOg0PbWYZpsLj
rot8mFXgDefVBbxwdMCIrlX6bQY++gqIko0TzFIjvUaEu8LOErkArNVJG83xmeWNCLcJvEdIL7nL
aMcwAdrtrcMJtcgGhf34V+PMakUx51y0crboEkAZ6JYP8NpSXK4GtisyjI+xxCeqM+AcnH4Axphz
wP48SCXN58sUzuu2p5rPQmpAUlUnyAcSLRLULr0duTgJyIOhJz5YzIg5tN1FHnMiKU7heyZD5EiW
NaTcCS1sLTQaYzdgehEFnrGcm+6p0LQ3d5CZ7fqP4ZuU3OK1jp3l0IbtTlUZfBfYkvEXDxUGmm1c
XjccqciIkTI7/yISBG06VvDrR1aLPlCIm53jpeXIC1KNw3VCD+dU7zVDFE9S8Lc5IABhUy5CWo4o
0W7yCe7ptzKvbkGzGwPwkwnzKihE/ZMeWTfBzp6fWxDf8kIb1OBzD6QoXyxDTvJ8lgnWI84e+OvT
R9jOsoV6su0t654xaMXMqcb1yuWikT2azUgi50x+qjgbInZ9c4osv841mKXW7K94p2BOh5OjWLHc
2Lwn9886YehqW58uf/NGTRA/Mg5XAaRZUjSotabzm1J3CY3Sx8fj61jpUIeLZGWfi0Qbl3BLxuag
3TH3Ic8m4AxJk5mlJdWUsW3YkDuukNW58W/2CptcJjgyL+dd+Tk4W8DfI+M5gscI77G+fbu6iD5+
znbq05vXSooK4hDo3MnuHNv72bioXqWsmjkNmplq6ihISDgwncYCnQfoEavS/FfuGS6Q/r3EwKfP
FOqw9d5asBSrcCBeZyC6W1tJmWIwcmoCzFHJAHEOGRghbrKJNTMSPnhZh+U2hOClyXGTxoPS6uM6
jXAdCF2WuRMeH9Vm+RDQVDAwSpKxZXwEtVSrNEiSmP/LaCrGVAgzTB5U7dQA23K6spJMuol1YrSN
6lyVidWjREDH6lZA3t5ScidLem06iLmVki+Z+LPXEw/tVvm8OnvPbIdlVLTOaq7GZARtuolxXZm2
/ssbkrRlNiM4jpPGIYHxqvYoxQmtetbr6Eg70KoIVryyF8Q6laUM4QFStZamY1oxZwdKVxS2G16E
S4Pl+Jhm55QottiblOaO/kotLgbJDHa8EA1XqXJUKgXkTb7VWLuRhxT7nUnFO8uaIbGqHwiEKKIJ
DVphAbbfpIL+YNp3t132aZ7JWeghrXAEaS+VKRoF5nLIBcmgUS8O2iTqaW+jSMpdqv0TnqLuaOaZ
DbvPyik61/eYLJ+cuihPNEnMRpOKj6j2xTA0Ii7j6hKVm4VUUnbY0i+ta4atoIVeViqMfJkwCgzo
4c7Y4b7n4un4mWkOCxFb2pHaAqRdaZ6ohcplqqmss0/aj4qBWMJzhms9mQ6g4wRZA15Nlqc2bcD4
G5lQHbpQIKNCoqdj7Yd3Y0n8JGMSLw0qOe10IU84vhipVD2IRjYmQSxW5MQ3Mfll2uXndlBXAdIH
97v2AZsHMkKdTpq6TyVOa8uW9SVUyOQ+cVRK3xvUTK1hIgNCBqJbQZD4fi5SwBdp5QSen/jYE+qj
WQ9tzh/WYCszpOHuLgswRP0Wi5bd+IulRaoA7W8X41GNICuMjZ69CtAmTkqbEtWbSjMRTgRbmP0J
z10OUqYlU0LwJ22PXOUMSAJxQwfq4xgo7skcJn2VW3xwQesm0YlQQg6ui5w9V51+997pqd18dsra
XoqCKPt6dMn4+gPBfBm1/gI//EeDVoMw0B5CYSmzvElXdnK6n/qFN3yIEiA9bx/s0vRwU/C6rzzk
rslZzoJzLiszyA7YmJlwxc3ejuOJe6C479ZF6WnRcliwpi+ZDMlGrLUAqLBmxLKNrYvvXJb4hsPc
cShXpKK5hX9Zk3q2nBfCHaCznnxeHYI3+7VTkkdYcLXdRAqL377FwrJrqb4v2EkeKzGxyW0XH42u
I19C0cz9XLI2S4szdqDYr8Gv4BHVH3XwmB9GcJXmHM5vngFrZDSii/hLOs6QFQBfiewcFI/+HynF
G9oTg3kKVZQB7FEBSCwqaHAl4I6eecRWvkFX5Iy9iNeRcaEJVxvw2pt8zrii5IPb76YxTDX6FqaJ
53JHAoaGNQbqQlSKokcXFnpnR3ZxhPS8WYf62X8cUihk0k8FtzVVdT7FaS0+Q2dQbGRnhOVRtxUZ
VJ8ytjZspQx2EluOtyuRjqzImyXiqSrFcjDKAZ+jgtQuQr4kh9N4kbkf55ts3wLDTWFAzfon194Q
YXUG7n7S6m6zdxwzFDrCYW8WgqaSXBffbBcPaGluuuhlxAiR0bT24IUgbFJ8FJhuSl/uGDiqzzYM
Pko9wzp+JOWbkbzRGiscCvFtIpHZOBz9vtTmVDqut9KTvbc7xmpDYuwaiDWZFwc0RWxQR51r1CUx
hrHe/KY0WmF5xjqL2xHjrubUTmDqJJ9EtRisguEiHoTieKIc0ZbzZPFPcrXY3RAvStnXRFxVJVhW
l80AGYbtviN8jNNoRTaoFNBoeoLRj2Sgy/eJ3vJx+414d66BzQiV6R5ioN7jRmcMHR3GHeajFAN6
IZpKr/N0F92145hHNre36FaLytd6M+XkqBxOHQI+qQhMJuWTuU5XJJ4q/D4e8ZmFOgEhLnXClqxF
MIPlAcLO7dLumAJhgMawQTFUHhMDfnFf79d27WSOSW6Xziy6XaqsbTyo8mPQzHlA6gZ59TwYfUQW
Ei8as7wqn6WB6767eSRaOVPB0D7INjxqngya9jiKnWHeRQZE37WCpsVMj0fykSShTSZYsr0zbXaA
doZ5uGQgp/C6HPxDZQotS+p01mYKpPSmjsDFtP0HwmPo7zZW11pUiFiOwbQ8/GIr9Qsnwd0eYVgG
ElFZWch8cpQge6nQBGxhagbXmriKcQClhDKYfFLmTo2gOwYgp3fXJHgWU2iIjrT46cUSqmAB5Zy6
WCrkwTPoNjgDj8Oma8cQZgwKQSGnZqLlEn1FUcPHyPxzeVzmud4vql2XiwXjbXGypxINqFZzKvgr
9zD0MoMUGATZzOyIUmsfW914FkRRXnU73Lv0NfNv+yFjzUcpAs9hke7v/0aJ+pSFQkSFHDkWXjUM
47nw8aKQSLrK9hX90T9I7fbBekZvGRrJehzpJDswcBCEecwAC0ymzlLV3qNDTV1SWH//MVi6SbMM
qjpL4oODwRvjKDAUavyKapZkzSP9gVqOyeaPpaMIlDXP2llKI9MFZyVCQJm9q5L1IObeBrCyVQMk
2jUpxJBm7b68xUdqnh7a7LvnFmRYDiZbH2TPJR0KnnEXWRtw5ax3iFwc/jwx4bzlQ5ND5kPc5w+P
4eOrvcltMV6lPwC0UMZgU6pTj21N4Qs055OrPnVphBklB91dEXjk78I/I5JXNhUnzbnV/oIziEdt
1utB/S00BnoQ28y8jAiMYlEa7v6ZagAycg7pyBg12vPxDPSvAoifaf6yn+POMyjTfg1Q/CXMaUvr
lrIqk4lkyBcHA5jcmXS/5gGiGZzepNNI/zEolImfk1SE1bMeYu9ZKHpSJq7kjWpt8xKEpHZ9Yh1o
LTKNwhqdsomskqq6MMuY1gj8qOTji+v1NbuLI+nDWcuDzltISHSlpkzqwvh00Wmw/ChBxAN1949O
ArbN5kTj+SRYGJhbI83SdG1eQaHLPMq6rDQc6UCNxIA6KJnexKdg5E7aUSCeTl/cToQVLawDeqMr
k43AWHfFIS9JN0FG9/7NY5ARisr8+3PH5bbyQ5TSeDeSHnL51i0mfVYAaxuHT1AhyA34Q5I03Myr
G+5MnStuARVcc3nEIN021PuGLCOqNUF7ey2L+g9/K6eSfx5vxNgAe1wqWl+7IAvPQ8EDd43FLJ8n
bZTA4uvuuM0gvosVo1UBuGJKHRlq5CIG14JKIRgWKDAdd+NSE4PNmZnGsG0Dd5P55wE5MclXS2m9
8gs4FsUgADJuV9JfAsy/ayQIEd9RmrFhJ0yR3Q9sG78spYQSubG5nrBWtohsBZ48/FYV1T4hjvNW
Tc3wkRA4XzGWnghSxXWYLBntRjwrw99KhuOcRCpgFwzyf2agkbzFeCv2YdoUqpQQsyTkSmc3h/w2
HLvwu2M+xL0E0IO9kXxdAVBDhwNoHTyUvhvl2Zc1K+miDefYkKh2jM4jaGyKxs1ELn5fvqtLR0sK
zrrtZRgIW5MdXZiJQ5ivvq5YvyMcANE0MyqQ1ZRIV5FIw/U0eKdMCHx5rgMgtc7dl9ZhMCB4+m4H
PqGPEKmMtUBJSzLajcxoh78rMegyaramUTlWzeNVjm5SuTeXCUeTbRxdB3UDudusiqNgWP++VMXG
Md9o4VZHpavSbS7vOsNvqqY3OEqbB589G8MZk1Xks1vd7OeRsLFrZeuBhwVAnANrRc3wW7e+cKoF
CWlbUFA7I/KohoGCAvImO/sYv12/ZcFZr4jvWXRdAtiA/Gsr4CY3eDQEUE+yvI9XGWuoZ4cmp6QU
/Pq1EKWUCMM/qoTG/R4vvAGdMOquotgn+IzT6NRLeTWLyH0F7S/yfqI9IPB2wjUjy1gb3zRb4HI4
zyGUFxidzWYNX8QIsKVx6dltMYrCwtpFUa5eJoLLmoa//1asau81Zf1qG6IlTOLXWOeSNXJvurv8
eEdOCVfLJKC89VnOZh3YOipo46QLBNzopjSoQ2wuxxJZqDmw90tO3+/exQCpq2FbTxrkDA8g1Ss6
2p9wtFT9iUZdaL6LHTZl5rV8PLv6eAzNiUT0tij1OKQKruYryeWryMqZwjkIzETdJrSUJuWY6ne0
bQ4RXVV9dFi9YStsvy/j126///MiWoKPvOFG2Nfkm3042M8EpVJqDfe9voqRVvQzT9oRUD5/tQGC
wV9dDMfcE3iSByzQlveZ9YZFp62RdNfWY2QWFQeyP2LMKCroX3Y55O5jbi5piOwefIlVeaT+K4aM
qV/CRu2L2qy0l3Hh5oFmj7Zx3B1jlx0Uw8nTbAHY1b8cBlK5CTXB/2qDs0ND9jqdmmyUGiHU0twk
xb6teYYseBeMCKWvgFURBVWvB+IM4u03eYj2q3uN2Fa3Mg0H9FZaadcdPlgsu4Kai70gFlpepKBp
h2Q7BmQcaTjEo0B5kXBNA1FD6nbQMT/viEtIKspz3rvM/Sy2xQ0JDjrrhlLwyYtebtlJ/pKzDdZ/
9NcbRKtrsKEx2ayPLWvmOMdDEUobJG+GnYZGjX+hw/Rh95k5mWkiT9hy8jBRHMZUXh05qio699z/
7ekSKM+py9eBfd8bkotsY9ocHwO+jV3onoWwnvkqCm2ikyo2dxmpd6qu46tx8+3qAXeS29y6/46b
kwA1fnabaXwim4U2IsYkxDZU6f4xzGaU0dha6uZFwojz+lIQ9+AhnAf+gk+/MqDkHaVS9XKG/IVv
5Xhky6rveVwrhSKAg8ZnyEaU/2/6y/V9rMedPHubeaOdYbBozNwnMlX5WW8qjUz4sHyhI/CpN6r9
CvxWoNE9iMKq0b0N99MiqG0auyu9Df5r9iIc/3NpUHY2lRc+O6IzWsLy1m9QYMW76B3qZ4KpZCw1
cvU3PYd/E1oir55jMMAqeKvNOcWSR9DchZ22u+n9QhtZ+IBtcRdyS0x3S+Y6L/kEuZx07SpZz3XB
wRAF6b9yuwl8cUrI7FPz5jXtnsaHlHPFBc2LKIcBFKOoGIsnph8jIB+wiPpZkW/PE7Dkuk8xv6gn
AN7+bImhPYk8nO0MpxfEfzjWMBYKDoUR9lJAjJ7e20t4p/CZuz+IVx1xbmJAG+7PW8DHM4abRpof
ACLEBAzcb4Y/Xpixp8hCmkp4EAc3MLLovCElHydjxLLKw9aQ36G+VoFG7k3Lv9hPqZsFw7tDNsV9
GEvfhN/+tmNnT1yJ4uwPw1anl2TgRFh6z1tWvI3KPg1KkfpliXFEfll2UJzXOGlZIGdCaDtqLN35
f80NIdgFIRPZBDrtRyUbxpJrCdwSnkvPUlpluJUf0c6qRCuyXQRQCCUv33a7CCXUausSiB6cn/3b
bZ4cswABmrKlyCZi8x66FXDJNOATd6O0PvICvHm+qQ0oZr8uYiyC/xGLGE9e79xrKWaczMm5+ScY
Yo3FdLlcmOy/hMavMhR4IAHFIPrPl6wjLQBAsJ9c8V10o2sJXlPDrX/sNsk5eNkjK+V8QBkNyC8J
zeEVwm4ACpFJZhx0atetvaNHPT+nQPQByjtuoztJRNaifgQntkDjxR/zpp0hjpfydnRiCVCNOfuw
QTKYbYZ7QXpNXMcJNlSz+X3pgDqwiK6Ge7sWWq5OblX11oCqXi1BW8XQyfEYMgUAHDIarT5Obhcz
pmshLPkGbV/U5AbMPG74QFesc0sXcPkMwJuQLr6ijIEAG1S/i8Df1LK3dmH56zMBmyjcz3INpBmN
x15jcmUx80i8b71f7KJ1H1uiRIaqWAv77fDUYTNzKsaY3uRizFany9+7W0tjlgS5mIBexgenERn3
RsWV9oP5w+/2N0PlNjGKr+/jAhyaN7n41xl+4yol/RvjHWYn0OgHYZgs87lyyk+AmCjtYoRhmK2O
sgoDpFclu7s2IjaD5Mr49/R0MTofNsGiVdD1GofmmD32bheSTDu3IA+5M6ZcOueoefGIMERr3Cq+
i1LHJGOcdofcyAe1DbWkrQOm1KvpHpq1Q7ifKlcQarCGCusjD0wlUgydky67IpZd0A6ldaV7bNTv
MX/anuVTa0s8+4u9wWvKzewUenUQDNNqbGXUeFSA/MjJ1p7lVitN1/EDiDs47kH45Q7Hp5N9UZoL
LxRouY2lEnY1vpU2SxGVMEKH0ykzQ4tbAKKm3F+fGJXJAf+agISYpOsMeTSmXuW4HSQQ0jROMPHY
LkqFqb1mNwZ+Ku2wlCmvD3GpbOIYYOEmV+Sp6PgaHR7zHNNEjzC1fnuPj4SAT8XZhy619WT/tJO+
pXcJGyLZtG4WYWjkECRGfV/98AXxcFrppJ2Dclfo8okGWjLla+/Bv72h05y+KUtV7kNRdjLCb9hB
xjXKip6JgOWaXUSPxx/YyNPlav2bIA4wJXHHbw/On52QMdXAk99Tq+pWwFnSHDVFjEpwN3AromsK
+lIIzbapSVleQpM2HLdCynYl0W8igcXJV1itkueQnA01knJdi0y0WD/uNf755Snbtnjcnmp+n8JW
cB+4WEdNNVgFM+KeQQCwDY9TZmydC8YU59/thiKFzudgR0rZYhPgv5eOm9o8CIvBm5n09i2m5PI0
Mrho6QArFiqgzecZrq8jAuHy+UyJC07w3F2vStk5ythGTd1cd0M0ffFB14+x0jGJNe9Q7SGat5RO
bCsZe0SovF9isFt90X5X4PuUFkbnZ9sDk75UL3wg0e/GStHrndjCZhNMalZ187zFM6t52tTVzmJL
dA7rcUSVD/pC0YM3Eor60QhAu5id4ZRo6gybXkxCGjQPF3QUxibYXZy3grLQNYuJH7D16Q3NzZOp
OeWAMnsBxi4PpZjFcQotNHE7mp/UtWF+fDFpstq89CqSY8yb7D/37Qh8+jIWajfoF/zT+JgXVFnV
QIfQERBhaT7xM2V6x1Qq2LPm8dM1rm18+w0J8o/Xg55YB1dvsp+mGpPE0f/XagAfXXnweegx/5Pu
Sd7D7UtroKAQcJIVeFnYwnDDokhc6aWBqtNqYJqTtDxMPpuUoz7LlcgGyPrvMAayc/ZTB+6FTma8
4E9zmYhZpRFz2Xa08Ig877tDlvEGTO7YYz9K/M1VcMQR/LkEZz9GUGvfp1DbGRUDcVzyL3h7ZCjd
Ewd1ir+NIl5V6yf20LzK0sW4+WGBZQH33l0aDtM6LHv2SvUWZbExsLOnCGFjBNCM4EQM/hDIGxXr
RzJnw5jreW3tJleuAG0xRmmy5rQqsy6Iw5jpk1f7ugJjj81fyC3wWF1vV1YqJQy59yaV/2ScTlEK
BDSCHOrtu9ChjyVrc8PAFUmYcozbWdstTdANsxU/scDIm2t/lJfX4gW8DDcxNL4JVDr6Ph05CPRu
SpjfJcjE91AEjLIkhPk5QHE+/XNWqXE0yyJ48IM7DE/Xn2vfnc4ISlOu+kAX6pbIR1QeppVvpQp9
WbPxcMwCfey989VKk1nmCp4ZoixpZyG7SrTpj1S8XpINnXeVTXmq44D7p5zzi7Z2aEZEDHunTY/O
j4cKqzlpT0XpsQW9Suf4Od2zbL1M1qoYQhLlKxR8nJNOXx0wllPvPckFzep2TQhATdQ/tTnk5tZh
eEUxohTW+3qgowoH735iKUi0A7jZPHee3tncCMwxxNmpJCxS5evMIO3m2lP579grMhYm9VQs3v1x
Gw789zlbsFGsQyDPFmN5CKzyllPxfDLLYTyZvNykBTga0/zncRpHqA3CcgN5mfGlNwZ/J3q6AEc5
qSQm+j0HGfBmjN9c3omi1x+q7XbTyCmyDFjdk1aI+IljC73V2okv/Kdw3/9lM3X/rR/uqA5JYu+S
OkISdLqyhzTL1ZZy+gJpmQFl78nrg6GB/d5KYvmUV9izdwP6zJLUqo0J5aOrtXZIGiNswWL1p9na
hrkITtI8vztktpZZOpNS8zaCMi5F5lZcO6HODZU2yBImuYEJYFQDki+rkj6mHfMf7DtKRB3Thepc
twO3LQgtM0fHhSddSzGqCK5AOVBtcG0uadY9tiT2No0DddYT86K8RTRjeCjO+NG84rl+l9IYInZM
tensy06ZPA4f0MgQCaALNr6hmeLUaXbol3tgCThtcFlnzKszkkUB07Hd+86MKWKShT/rgC5ThR9j
6I9JrIOBL2nk1czCFZwYyU/r7xv/b6dhMVEAULKCGUvttck9zMswX+I49JZuB7ghuIsI89A3EN6m
0XcaHZQtvzC9d1itqVKaTW/Q9ZsfVaY6o5xI+1GdQq9kOF5AVsH8ppF3GDKrPWQSP7iAVo+BxCUn
yoIkkwolD2BbMnoYxTsOyXaJa1oLsfrp4NkA/tSu8CKd8s25MDrtQRFQaA/6oFXGJW73KC/4TU3N
+VF6xdY54qQG42K9tQEE/QYm6SU8c+yfkxSNXsMu9A8b4/m/8wM5KZ5hKPe8X9Y5UGHvKLljYFwk
iScGZwAMJ+17qx4uwyiL+VlJvpZpzaSDvDIw3LVOoUMWhtTmZnTXqaedClekr9Cs2TqQoqlvcGBm
+2TByaxaTRKJVIgzcpfsOcivdVwTFdLhA729BRbU+WRgUmhG0LayHvo/uCmhB0iL6/VthPBVqZi5
ogQsloSXjSRQ4GQDOnzVfqJpZzv8h2Iw/A0ou4zYZzncAUc3lipmGbMAmplTmEtK8A+gg/mYM86E
5mMe0mOe2sErlKF2S3xRDS/5NmQIVlfyYlw+OMu7xh0sJaJeCE/UwLYcQhlmpE0TTRER3owk7Z+O
jff74W6dthg51EPALJJvcG4ZUTz3g6oOVbtr9AhaUsDK9VaW8+vvskIvSr3yz/jSVXqgbJAjqc2V
WO0kPnVMJdOurdgcQ4VVz7CxA3xYzz7iiDoVJvG+tBJghl1C1HpqB6YGLY1Y+LyVtEYegwCr5vJp
W1dJAi0snhB1KU/TGkr/ooRNWbJGTLcYFIyanUbu27oOrKB693d/1XOnrreAfirCauLedEcGEsTH
DgUOBaZv7HMVIwm9joGyT7rgmGCGrnNYsxx3u9opnMBW8Raa03K25tBmrMd/59Ehwctw0nbsy+n5
27tRv5omWJESHWInty8NAtGAakDyt2D954leP38My3njdANZdffzN026OUuYs5mzD1YxXeylbNu3
dhcRDlsLxJCVTul0vdkWl7KHT0zx5eBQwV1RF2+rSWa/80pioKzCih+Z4vT0oriwKUTPWX02E4IR
ZxSsEqSNju4ZIA+bd6OFMJKfsZPrPRzsZPdXUdRMWO3qxYS5PXHYJ13e5OMbnRfYme3/qN+4DwPx
vDi+pXpeosoDDCb5Ta2Pyl9uYWfHju3bx0DJ8xB6izjGbvtqWPILKrTCALIVK0uwPdoqAmZuBjYu
cu03LxDtrUX1DzTKfso/cgUY9xnrQMB6VzXIU7Fp2vepXdrAQKnVNVNWhfJDTMspMmMo0K4k+slR
nxYbyz1IwINKcXefiJPSdk4MQFFIWW4GFNBcadsTDWl9mH4sYlvQYZQI39Kp34JuKRrCUVBSG/+B
LkjpI6FY36OSNVRUl5apzbeSeEuMhTqpXr5SvFuBAyMg8sz9ebU+O/5njEzK29BorbL2JpLFZEsC
IYNP/5oTSvCACdVAV8mnnsMm7RXgYUZozNS/8M+ofP2kBbk8ChVKGp99iOcs8hZf5tc8b1+insYp
4fg2knyKtGQGs/Cns0/E7MYzXHbxmjjWpRmomsbeLFnCveS/O1bOu8hyXHxQT5KOi3boeQP0ZzrK
5MhPoqMdA+Dg9aHIbNZexlzOVFQ3D2F/56etqkYB+a9BGVc2n2aocJ3eq1YMgL4yTaXkl5XhgmB5
D3ZzZlfmQgzuf8bIk/oOD6DnbM3fRlJMSp/O12L8Zzaxq+SGly2tpWLo3bv80k3760enFH9AadJv
ScOSxHx13bbByZ+qDEW4D/gFtZe9kGSbt9ZD1wiwR3ew6W8lrAn6ISHXN4s2/Qi0OwZg5vdSMVyD
/HehCBAZzb9hJxKlIUX+XwPOL538OnyrL9H5gNXN87dv2Y40Ape45y1nxc2uQPOhLDg05Qhm8Pji
+SP1537vr3tmQBZFBB20NbJSu6mSAdgv7Z/k7IKoiFU71b3Coyi/Q722tGNOKVbRUbGK6YTscZZR
LsIcCROV5unk59ojlhqNQNC4HT7FYmppC+OxS8t1bThNCJLGWtkL75j9YxNrW5eMHrCLrLghimnB
dNSwFLkb1lfeZ/u4qM0rIXoWx6dtTgeSO5S/t5mH5Kfd6xOLvKbeFQBZ2bnAAe0xg+xH3YOxYYYa
HIdBMckS33kJF5N5Ssa/bEQh42pQJYiYniUt7wQ00MEakYTL4Hj9CE/yXdw0JwBsIZLjYXFhBAYi
hmHfW/SwrC4cWVnLPLlBIklr1Mf0ge591Xg54/1QYJclvS2kCiSiHvg4iQ+IlmJr+B55Tb5mf2Ca
5E6wDyZcIj6GqeNJRhVc9dBHmAeUGj5oFfht9vhIYu3gWYgkuZt2IOOWhtTjcLQYBu75PzylroYQ
ikR+27ACAN+mlD5HVSkZ8UFG6skkDjMZGIrUK59k/deS8BZy0xFmQIwQDZCVSKMwu89Z42+IOSP+
HGU69XQn/vsmKd6MklXsdy2apdFVUSCs9P4pk0DmHlqhpQashOPARW6/rzNS893xoFta9wCxTJhK
6rc6cF1H85Hw0Pgy5bpdEwLMcXsyrvGLWOiBt6e0X5NqVGpshrf1DVuBDnh/m8EpEhPOu8/goZAH
6Ama86tE4nyHpTYgqJu7XAlRnJKvT8a6XLzudiS4hrqMriwtB/g28+6/n4ZyYHR+t0I0RlqC+Ni/
Epe5ysUffaNbst1Tkz2YzaePxvULocrepFHOZDVU0EOEauQ2bISLcXd86mMyMkbEy2rthY5gHbrh
cqO46HsHffrSugBG2YSKpJlZ6uINqfdiFAXYEqf/DK7nCB+iNb55/BGG3D1yUjcH6VNeFf685lFu
u19MAhTmHJ1g/3V94f9z0qoSh+sNseiAliiqGrwZPmf3bbUBI7RYtaO7Q8aAEjw+P8Z+JYyjjWUZ
rxA663Fyvyvsn7ShZi+L/hYIJWUaOPdegox5t3maBmeBsRnX+vOJfoqibiX1J3JcfYNxuOfWEwq6
xUalrdBo5Wj+eu/g43kVQLumvpvKapZsb28a9L3ZZkCOiZjZmTLac/SwKbQmzg6iAyhbER0nz2Nw
ew9KdJLfl2MI2K+JZ8Uz7xcJM7Cirvouq4BxG6qe2yaR/H8h46tfTJd2CgUz8QOZ7zUvyfw+1I9C
mjVVaWQZUC0PQNPyfiYJ6jPB2rR6Lfsr1I7++jB/OWu4IAf4bCu85jZxPs6NtzL1bUhT+MSnZ1B3
WfSIY8a39fUkpIYfLXeM2KNSlHWh8gMx9G+SSGdqJpE8JymXOhOEtAhjTuBT49k57a1G0cdlIWgw
0f49z/w3LkGVrjdN1j40jKmvrEmjvmFbGvfcwwyVVA3R+Uu3XW7goAlr3yq0q1USKZsU45R7jUEy
JJ9AD3x+561qqhxCNUi0rEL5eIclhIJnLNGaUsA74c9O1LFIW7m2WgTqT6k2NPyrY7W2/L/IaECz
EAPwU8fdaIztoBbbF9WyBMwqMVVJwaXsaBEou7vgixXaIwAIwwRKS007QaLjDIS9FYTxSXC1Scwi
ztxIQppAs/035NHdysr4f2QxmlJ2hMoqcb8keKTQjx4q96YNUvHrhnLlajR+3dbomA7i/yo7fPp+
OtURKGsL3RCinEW1b05JdgyWIYe6pXMNPyZ90emkTOB6WHkaKJIzo8A5X2i7RrRNy1IiGFWgkoaU
xJglonwlgXWarx77C6Q3dYusDjGQk0KP19mwLqrDV3t5V1WMN2UB5uTCQ7PGIXkXu02HncGszu2N
fWQPa+KRb+YyfXvwAPR2MgQK+1cUCffhy8dtINcfjeYV2ty3gEYdW+kD3shol5Eil5QeyyTIRK2G
iqiLMDuKaq5p61S2Fnxz/XKkAcLGP9IRzciwQYk73M3lE0NkImgNtqk1GMJHJP8jYy6wL1MjRFtW
a+SC5shAgBD7JIjoX9VTOihwqQG/b1SieaeMRl9vfRUv0VvpZQMnTIHFw60RIQLMKR7PkuH5Cx3V
UC0uJa4uGjxbUCrpekkeeFEFE637xYavr46fXmRPyg8ACWSXonTrz/e8IHnil8FKnim5JybMnG0q
Jf9l2IWvBdmjGt5CXkd40XaBqzWL2/E0loeXtlO/wppElP4Mzsgvoi8/fhu1EGBwvzcWTFzAloRa
7AFDKsYs/++ZRez+14EEp481nDL8hMX1wPzgSH5LvZUs89MfIZXwbIYSA5UNDaAkFyX5xufTRQdF
yDKAtTaywSedGleSuevqdnBPaFvQDiGz4xxC8bGrN96UHlUjy4J1HMXJ3aaRivJ57KjM78ChYjRU
we7rHsY1CWFYyf83UGAdYID5Fh0uwQ/dyM9KkLtdVGtRBHrYyqpd04/PpLMbMZmF9jTRkgAc/JHh
+AY5SnLDrgvix4zPGQ630TBVCoQtsLT+1CK3SBWh0LcL39C3ENeyRTyijHU+XEGFWNoLNe3c09z7
Ii2hPvhB1WzAuLhRE+30L0CHh32XxTi7s69qJpWt5RGFtWWcruZ/q3JzKs6wLQxJZMemBlb/WASJ
NMSRiYmLk4LMIQ+nxJW2IVoK6qfE2NqhGExbqcoeVfgTwdPpg4qHtogoy5N8sZQ2AuXHhiseF8WE
+CruGEADtx0vCsTEm+wNXpnbjN1l5Bg3hFMrcmFv5F8nSFaNfdrbmRDZhGZ0jHkXUPVyMaAMo9I0
qQPcbVN418HZN2Y54EunlRtKgqo2iQZD0uzJfyAmXiMXrx2Umy4B9hpW2Wt6Pg9KQzOzkQS/+KRj
AJTSJJdREVBHVbzRV/ZDiCKrUZkctOQOfgMkY0kXoXN4TbRFHQaP4eCUkDbPnKpoY+Niew8VFXdh
URU7Qq7W8Fil0f00J5GLuKawfdKZ2w2vrBqvj1O17MA9hudpOn61PbqdgsyouWqYo+lwubw65j3i
wlRt1gUE/SmnNo0aE7eHt6lxw2mbB4GS5ak+TKroMAIo+Uw7y/UTa3hiWYPPmPZAHQOPRIUib6eS
coi2sq28rMRp41eZkE7zaaXwKDVMSdkomTzKnb3ilsj36h5KD6LB/69vGG0RiX3vDGjiH4JAXA6t
1fZqjkMIIsXBsnm0iCPXzcW10PHZ1YMN1Ttb3hxNcSyJlLSsXDi/reZwmZgTajFENPnw+VGRfb5a
S2NYGWzfWm47aoQpt3BshM4L09pHNlsjwsZ73xezqVjrg7p6WAJYL68d+1WrwebrH+TzflZu7ajs
PnMrXSLEmvX7CwhLNPs/vUgas8gqGp+6Z8nsxZkP3JHswcQ5c+CL68KWPVbjflxkqJqpE3CJeQg8
bSe9NVyBVtMOj5c6RdBErkJNeTnNHqiDzP+QLS74B5KgFFox89s4PYLVMduRJvakcGA+tDKfUplM
elhH0ad/+2WbEkBKIrB4JagXnMofJRTKLJ5CLD8B8YPNbLWIqKCSvJd7IWQToGXO4tNRoh7nOMDO
rLkPQVtdV/IyT1c4/VvpKWcHeYx5K6snFGBxmrYERIIv+OAyM1mHoyq8Irb10F8aXGBq6ysv8Tsk
kJYm//I/io9bzKoQDGn4ap8ho8ZVmBFOkQNELAmNEzV86ztQ6fKbh30xB3ad3Dj0nkykfirm6//Q
X3E6/S/eRpBADkSKzIvoCyQZ/NcrKQyInMMKpkHzRr9sar+bUsJbarYYoBdZKfhASHZWct90x6pL
M3vRGIug7h07THcRyaxmN9PtymxXy7iPlWXf5Zx6xh6OQRjCu5XUlCly/x4E0QSZ2NsdKIs3e9mb
189AWMRkQwittXYnW5eJwSS7fmTUdkZuiteJoO5DJDfJdo85Wb9nsO4GvDWHGHV/FK5P3glgI7s4
9/CHZL+kCHcgDirCrzXJr99JFXs48MwDBODxtad7C6PYCN96ufJFvHV1OCahDLSNVC52Omz5Gc6b
zAbN7YV/tXKBvODqXX427TV+pfD/7mM8aP8f6Rgj5UTFHMs7sL+A4R3KSM+REVGGajQMo8gHY8Pg
A0ksBktC/2cchRGbikYQ6IRaJFXGWm9c9Sb4ebngbCV1K1bU9GSwQ0G0dIEA5P0tip8rUvh1IHn5
/tS4HRN4pr/8bBBJzi/LCKy2lcyYIxlR75I6NYYxgzFKR1g2TPO/McH1SsX6dyRdFNdxywNpOA4C
HdZ1tc32u04esaZL4QAg+/n3BXMIe/vEfy2dD5rPb1LXYE7M3Dn1eD2DCGfeKoKTE5Uj8lwb0KsV
szTXdGbISjxZVdApS6w4rRg8n0DZBksaKiEI5vqTx+DzO6SGzvEIIDGU/9l+GR4bU+iYRA29R6Ti
F8yL3cIvwYPlcxFIWDmxEyoma41DKi/Owam50Dzshy4F6HVrE/bWr/CS3OtWyR5n4f+fD1SX2Ojo
dmBcrYOX/yRKaxkR2RaQMKSsR2x3LCs1cLpq1goiYaJqIeQixHjtgNVEaHr+EAfs5sOKmMmLkyO5
0XCezvybvt96zdQa4OYfOnPI7BL/y/mmqoczGM0NjXqoF8md3nDFK5HIQefqzv13ovklAY5gFMlY
1uEXgxRqrsVwX9A6ek8HtmBmFBRJ5vh7nfhgkw0i5EtY0v5G8OzdiqQHdvCp/9BPKnZwDTNFHrjk
TsBaWE8QZmUW/4HO8Yw/eWK/jY8LHEI1DJQvxISQOyV/ZkUJaWypT4kwh1pI+dzRRV6EeQzSTQwo
ciVzlA8m9K9hEK5lBu1wW73Va00FgbcMiClxFQgKA0ZayMDL7fS9xkYD/qPUj/jKDL/bwdPz724Z
tNsXDU25GmO9SfuHMnQGA0YDZTiOqFkzoK12/u+2r66FF1WiDd72hSOJRFm3p8mznpfb1D/Ixh56
o+2W7eyRLCcCVhk7wHj6wcW3VvOh4BrfsFBApByOIiKaTWpDIWvUVaxzy8mOqUlTNtvsRHDDSSPE
5+prQIPSjEJtyJrIR4iXNG1IqYluzB81Soajl9FzUCc52Qu3O3KlEoEqTWzYWp3Kcq+YZQvSrJzK
DDPPkxy0+ezpQGPwQKGF6p64X4mNtjb4xzzUOlB4hAhcQlN2pecln6oOqUGd3i+cdTwOoDesgKxF
jRBvsY/47WrUVo4/Zn++qYhVmXpmDh2uq/qGK+IZBYptvH+XrajjmK7VrEcTK4KP2b5gytNxGvvR
MDNIg41X5tVER8XccOcY6HA5xYcnr/VFJTmQrbSp8FKzjOL8+hROhXA9Iadgm57dyTtge5BO6NVn
m9e/k3M9cNKJAl4ue04ekgk6GR8Sn/FtXFvFKmaJHCKShgGL++5UeisCqIaQc75xeGqvJ5okhlwz
OgPz5jzw/TNq8GCJ9AA7M2NugHxpybPtZM2/CWnpRiXrwbFZM/lFwPNFEee9s5+7kiZLYiacP/At
GAonkmptqn5cx6bva5NsjXjYABYRbJ2v5PaBtvKCAzO8YW77wZUUhwXWPaKYW6eboJxt5CUDMUOV
2W50RjyvCkkbxL56B5GDcG1AI3o+s8MT64bjok/9SkORJh89JsZRH2hxiqewpGaNs/b13jodtrIN
XW+vgVlXEI94LYFPwCO5VO0PYlcDTCXw8SdjLIBGceV/rTJXJlvlCCC+CWS+eMLGgjrKj2AdH+8d
63Kr0WoQytP1jfv+W9AhxFCo3aKlfo2eK5EwZSFf82xKkwmRy0Ml8Z2TlVQAuG9uW801Iyt2nZRa
fwlwqCOQnQ77kkGxhHQU9AtFsjpY5VXzs2FnJX/A+DMQeqKJI3tx7MaJsKr9CeIxwIbAxy2Zvly8
Y1ikitGWJexMZWomWZhBq4aqPmuUrimtpHASAoRkU+wbSVfZwSkE82OHGTlH33dEwDOpnte6mho9
bFiKDJYDUIgCTsnuMyu/DV1cykk3pfP4xE1cHOWydAK0RwGz/VPWWjLZDw3s4H8rIxWd593/lszF
LVgK39ZaCq8g0XGAIgLABPcNcDAHyi7i9wupjhUKhUleGV+uYWU+QvBmgFsWHF7KLKV9x5G6KDpP
B07mFKu6Zs+vNSoawNl/6iFzB7x/jjIbJxIJ4kSmsfnaOrGdKMdEjAx8dOmwhHkwwa51jasp2slg
aP3ZFxaoOV5IwA4XJf0s2Ziw3B3BBgRJX3y53C+gFBgkMN7odTlCWaZkHRjMJB315OBce2gQ7Sau
JTBd3yHz088I3gcgNB5s1mz57oKYL9UxlZTVC7p/v+7bJRVzOpQju3BQMK2lUZySClFkpDVtiEvP
hmMJZ+M5Qfd5dlGxEe4Sp2wv1i8LqvvWQjC7HS0yrwAKj2QxpvTtxlVmAOjUTF7c3DrCSsctNM8F
yn0tbSgIwRIMu15XWfXXoPn9/riYpElqp30GY4faPPWtXdxcqAFmTRsROs2C+9h09HYeDXy1SBeg
8DAx5SeNQBz8GG5TgwtfjT6zpixSF07Huu97Iwa/gzbm6FK0sHiwBsLgeEHVx+RkUOX2S+raM1AT
+WVKCeJEG/Ao4WtYiF6b3m+3a4meJSwiE45vPhsox0HAg0cegQa4VBc1Uws2EuPjjUrCxu966/nl
V2A5SLsRaUxB7STKaRBxqd7iLjx839bosEWI4chIgZvpKI1w7tA7TvBfYaknZmjh1ZgC4D2C+ihv
XxckNeGOKeQ9TRHRTkEGZFrNyS4HAIv9Cx7hnlUio3Y+r/1HIDXghB/rHd0e2HKfnSdsOARo3NZG
jq1j6QgmM68JmpV++jtg4blvsuQ4UAJotV/FdqzmVR1FggHNoEbBVZEN5xvAa9sRzHXEeRRxWc07
ZFuYeuq0ja5OWff23St0DqEiOt12SFfkjobF/0q442KU2SF73gQquGpdsTa6Pf9MAA+6h3SMShCD
0grtrTxweGU+HZiKY+C34b9j83pyuiDJmPcZ1EIntMBnhrgGrIliaOVVREKZlP5Tl11cCE2WbiPn
1+cVP9i7lHBezVDTRhV9DaguZZ5CfHa2aNOcYGaNqMf0kl2K4KVOr0GY8SgOvYHJuwGmtf/28Smi
7wnrLGNHoTl22u0GLisFw/Ufeljm84pNgM6bJELsfbkAzycJPRNhMTDN5j8MCATtUlgLosBJTpDT
1ZC9vMJAIwgjJvZcf1Lo3zevsFOy4lWCLO8Fo9hMx995Uvg7DB2VFM3uFc+uPg5mogMSe5f+xvxM
Rzi9Mg9FY6taVMkn+9/nl7ASIpzrfk2Hqswg3pl8nQhNnyXyGTX+j5h1f9HxBwWaQKpFumx2IsX6
mRY/NT99LpD72LJUaur2gRiPfBZgzv0pUSY42Fy/s2XjhJP6VtsUPxE/Ok/XRLP/4wqX0uzHzMfu
b+4zXEMbdrXj91riosg3/6LYbHhNVISO6x5tJYlrASfID9SinyZ+ehsNeCvUFUlUNNGREt4r5Epu
hdlEXiHvvxnPTcskILDsoiyO5KmOX37+VWPAUwrhmMr8G905bxzkVpOLEyXaLFn9NeD+8tfyZtDl
CsblBF6CKUjZPWOgwQUGIO0MQZaio04secZhTuHul6Rs0S5OhxPMB0Xx65hr+5Ceo11v6OnZO+M+
EJZBsV6PKifZtKHPrWqFL0t1t1H8Xir/nDrJbg4tNGE/+jJkSqJrkPkUPYNjUP84VjDh7mnU84wk
h87pfAaLTpg1pUcp45tLhr+AnQD7GET5v/onbK4SdOLXk3068kk5XXs05kRKza8YO6bCb1hxECZq
yyvULT2CNY5a/HbH8plPYv8tp0Jo9xuNBKnx7Sul1uT3F7Ih89KF7anYoR7tXMvMWpaDhYWVqQ7g
u+5XUy4IHR4D0oQrC45HfJV0+9/pWXRVm/TWOvgG75pIMP3tOw6vQphRm16An4hgrBY11ylrlFa8
IzXKHHbOqwMW6KW+WmUUzm0RLavS/g2XHPURqTTrNjgz+FMIoO0cxTjLyRI1SzsLVPlCvuYVbJx+
oA6tVu4G3Ipi+6zsXxpb+IF9EE1z7v6HdDsGMT/p+ynhG1XsZaAtiv/xAvXu2HRqTnRd1IAzKQ82
+qIB6ZekIfmAnaazF1K156z/mqmaaZ7DMnL1JbItlWvVdg5HRx2ISDSiEYgrQnjokGTd20nMeLUa
y7EPoJhUSy/ADXZL5xboKfouUIEL9JzepK4XH/W29dkYiadnHeTp0AcXcywTyp8fBUmD9RuUp09w
J0KKhfou3SHP/6DWBugD0nqrd+/CxiBjxt0o3MlCjrl/T0wvSihCzmUwIliYr0+br8sCzrpEWlhv
yqJGu/Flrx2q73Nx9ZFgk0/b6by9uBy5kNeULIH75nQVFaBeRuBfT94VSA/PySGkCzEP9iIBaKXa
b9GYtHD36JWL7HGzlsnj7/TXS4sp0V5rojfN+bBHy3NjnLv/J99EnI4HEAuZ8NWnjEK023Eq9iO2
fiOKme2XD6inuPWL9rwi/U5yD4fpuEPxVMXuv+G4c0lhKFZK2TCuJJhCiF/h6LTG0YkQqBqESIst
DLL/pU2qGWIwvHO/e7l8N/Pu/DyesagdyCS1G9hty6M5UjKcxqVoEC7KtxP9oMhsCX5TUpNIdkYi
t13vgJY1FRiui9gzLlyaIHBOF3z26Q5ivO5s56QX7OzlrnIpJ7TDF8K2p0eY+YxOEasS73bYduMz
3Guf/w8FV4/IYzaScyPw3Fy8i4cCfPwLYleU9En3a3jKGLYuykvGDEUC6pkQy6L5D3iEiv9HrVSM
OTPYMUhxUa68ZAb2tmtOiu1ccaFlU4CrGlBIPCQdgzn/678uaNtvl0sg3QTf+ekEyfAoeHZ4Vy+A
0E2ttGUHABXZbtVej91qvlJ0Tw02LGKNJcyuNypwaknIOZ/xvDVRHZUSXUf7KVwW2J5iw+kXVMf7
DGrt4R9gh4swbu2txXs37CsDmH6b3bbrb0t5CGL+V/TM/zU6mwT84Yc5b/eVV+S7q6MQ+lF2xltB
swn5onLkvKTX6yS9cBlUDvs++DxXI1bREbLMO84UH02AIba/EmUw+0hiS4T1oxBrsZZsjuHQYvnO
BkRPZyaZbzZ3Wk+ErSjqUNE2ljG4mQdJ07VfLSUC+eGe3XDgD+FlUpf1Lvl655ab9eIowu4V4BzU
UrD8FE07L2suxa2KDacpjLkIbgSAsx6YvfTryfBEzUteRaAh1uu/l8F5HtesR1BsMPZkrsWc6ekh
eqPYqlqCT4BmY3GZPGPLDLw/b1QLYYNh/pb9IxHXoKzfjpv/rswfrpKAtoYApo/TvpDQtjC/cUp2
n+XV/iCq9EYKHELRxkKoDFeXjlnOFH0oeGCApyFtqfY6YFNql12Utrs2ihC5My3YqrzwfZmw00x4
TgDGvjNsPQWaQ0GQNyqjXktYKkPD+3Me1LX1nZlGQmrdhoctCIXPxvJUj6+YaFB9Eb4ODfQkcfS3
OINJjtXRKfTGUp3GoqhRhFFHfMfrdGwhbTGIOtahKP0sjEC4XvOt4tF+vH1GU0twN7IZRRjmDHjp
52BVkJkWWYc48J4Tdl729LkmvsUCyOIWSWIV0H5pmQK6nkZWDMkSBUeEBwFcBwf+C6oBxnPPYAdb
qX/aN9Xq9cgCXirnNio9e6ruXyz0d7Q6qrwCKCCIoHh5rebJVfNWCFHfTx7j3tKukL/dh1Q3qLKz
Dgh7fb9Uoe+RZ2rpVrq2yZXOOwbey/9FSyzFbStWWZZKVTR0ii8KNtAEO18x8eR1Ba2pxfWjyjv8
wY7agP8sZB4DxNIHQ+oDl4g0W0bAnB9BRvomECBuFLD/Ny11ljm0rIRqs1+EW7A2LCEukzdN9XaY
hxgKfQPdEQdAuVJJhbHebYGT/s+hluLeoh3O/7ReoDij+YDMPDN9qiUPu+x/Dl6CCQWOgMyrpsSz
7juwSTmNXI0D1EPOxy9M269yW4vsxT4G/dKo4r6DlzblfZ8rcJiV+1ihhJP4XCozt1fErXqKVqOQ
J07RRzwkYEIlvtWfQUnlNsB48HWK8kMd4+lb6ZvHZONqFoqo2WQTxmZwkgQXZGUA+8cZgBdFq4Fn
aNlhKa86P9OzXW1CARfGpKua5RDO6sbI5xzwfoASBc5iwy5v4/JYrN+ZKJoWB4Aic+8kDaZbuzww
ha8MaAu6gN8edQxxCLOFdOZOP4JMNVBZiYQbbtYBYjjlRubhMP8kaKZeVRz3VetKvLMWYk/dQx7k
59RBrOMtGdzUfZ+O2N2ZS2edqgoSrgKjElLbZP1KeVCW+97NRbMLEy84CzAQwKBgK29Qln5p9dDN
HPb4Bgh7RRqQZS1FpbeOVLsXcy2JBygfH9iLlY8RtUogE7v5d+aAJq8iughfoSfZ3Q+pc4V5jkVW
dfNvacEBfqjjOrSxVm4FMDdqluxS0P1U3HIAFWSR+gLZnOn95UmIZC65M5PlenW5KtCX9Bh3fwYN
war52CQmU0QkGxRZ//W9z8H6VAjRZ8zG2lK9IhNqFRI7FUebua4Ut8PSFP0+J3qRYaS99nIZU3qM
YPfzHh3+wSAh9BFxKhGgY/n3LIBd1OeK4BkuUxtj+PLyPlD8s4MjhGtPFsd+MKMywUufKpkr9TyE
j0oOSU216ixUYXNSsBl2Y/sZ81T9N0TUUFGcj6Ymuip966WR9bN7+VS8moMc4wVJ/YL+nPNH0kX+
du+nfD32fIpL/hE3eEAUvgun96BGPwErWA0CCti9NdFtI2/DlADN1WXFbN0id95wQhnMgz3q8EM0
o//E3wNuw+6ClP29j5P/zwfzvt4jwkCCZaf+8hFKmfWBzyMpzqCHcwgFxH8MuyFeax0VADU3zSYm
zR2rw5y20vG8JIFq/nE5Q/cKawxzYgwD5B0bkG3DXv1jvrW8mK4l+IJZfYwschB4rI1RsBnFHAyn
N7YVs2S0o+bH+8vlcjsgerHfHgnGzJg/QGPM5iWyRRFk4bztrhV4Z6lCioLOzClqSfcvmq3bqNAG
GDT08Xxe0ABzVZjTcljvJkOHb3m9izWJg/RBin4Ee6v3Ki45wBmLTr/KH1bkyjliwV3rJNHxxhrS
/MIqFZheycH2Uhgy4fpQGFjgkfKjen3PfCVr+/rnSjQs1tvJ7KaBMSONhjF5c04aKcd+cU40gyrv
0Hxr/7rUVn1OwEE1iLihYp9ae7hNVzA1OvHSVZtnskOpo1wtGZVbeQjQa31uwTlrnnJJUmSK8qHq
Z7TdosDv6fsqKMPJQswBhNOiE7HYdoypJEp/Z+wNvNLyaD/HxLsYpOIiPcNcGAM4ASeyNWJdhufI
M6suKDoqBAaEV/PQl4yFTtozTiWoxFDws3cJvxiAoxaCF34aH3JjlOS3dXFW6t9npwWH6Zui+rwp
n7KmLCBLt+QyXp4j2tv5oOKnwOqF1ChiKOXrBO9mi2WoOeBuVr4NoxtCd55goWif4a1tDwjIom75
6g/+XLPlVuh19au5zluIfWac8FOqAtyppmWjbQnB55bRjqPC67C3aahi5RC8dpaS0y3+KcFvSNtz
73jkVIa/snkpFibb6h1kbQHQNXOxyGqMnexzWZIum0pF6MB48iTEwvtmqlEP2f/7sVEzUVa6EH0U
53mvG3KUTf7eJ03sMnj/lcmdifdp48oxGZFZR2liACBJvn2pYytGdGCSGT9tknRGzM10nhQfCbOi
5Ce4BpmFu/5MlW0JXrpt5oQU8jJ/syNneXcMm2fG8yS5JyIU8YS9izOUaijtA+/4uFUmM2Kx8PlN
JFBXqoadTJFhT2/UoRaed7YDCLtim1axMOqyx9l5d0IB6ZKIzytJzvpYvql2W1jNlAvz+NaV9dk0
AmZPUOGk2uFsNH4tD0oSUxcETE9HGzhIW+gRqYDgLZG5yogUNHS50Blwte1fB/CU+A4ySyzHA0rJ
gCYqDp3g+J89Fje34KubhqS+Omql+gVB8eTjyeSi0DbSwVwgaLMTqzGcYubve32nMEn6k0VJfh3+
4Nnd8/dJa1svUrX6+3tuZvDsw76BYY4G6WCOQS1lt+LcXhyql0sG+fzOP0Hh9d1MldBNgkpYuFWr
FS7OtM0KvLcdHRQCmJLKdSlvMZ5Q5bZnD+tBWG9RnyTUVmqwOnhl/RHyo+hqEu+Fv5/TPd/aYwrI
lHkmrWSIS8O/wqzeTnjxR4UT07WWqZhPxJZTgMWZIIeU+JsfizrCTFcztWqEk+rBlfwCboYI/Wue
EhA/XFprOz5eLfEfy+AUZHIdN3SZT+LU3/Lgtn46MynqAJCTpfr5RqTPJLWWgbXVbtQ57vrzqgcn
jSeugTttgFA82r6edeJOg7cE5X4oFwmXjzz0d5uYlSdMt85fFHmTLV4ujlZZ3x15fEKw3+ANQ7PU
UL+9cuKgitag+QhltMmesdwtJK4n1hpubF4jHboRrVtc+ejQ4vKK1VH/M5Z94KvUiq52J1pYal4a
fQQu4k6pTp8TqcmcNdNiG7xdc8kMhm0oMJN5fefAQmSdDQ3pJxc2pnNxzldht4jCv/J1ZwjbiwOH
SN2EEVC0eVZvW7zU0C4Wi3WAImuoQJvzas26LanZ0tR7Y+vblbnZjYuTNwAgu56mHL0Dsfqbr6eC
UfrOxuS/xTZRqcO75yXDL9mJ0UYLh5T/lwjOS+cFpNq+P20pWtmvL2fo+FlbpEeS1o1aWbbTuOLJ
omNck3m48HWydV7pjNx7uTUc80WA8osB3WHrsvt5LMeDmvPY0tl26Ul8oSTNztI2WBcsC41jl6Of
SVyjJUJvRuOLNNQ3b2w6NFOnMS0nw96GnODPBnV2h/3UDuUC6TjQHlbVJKA6/MOv0YW9MxDAlpIg
U5ajImwXvKQetN68bJCErFZst19M7QN/SkqwCoulHFD595wghLSKrXeQoP80JzsJctPaYPQUkQ6o
v7rQ7xbf5wcGcIgrO+jVXMBQYkmFwP3+LNXGLVH+f9usTKUPxIWa0+BbKPaONG98nuWzk0CYHRrd
+Tw8AAmpyVdDeGCzAUiD1lmCpXPBbZ1EHK4wO0HPjfy1BYFHbML0m1YFJef5SnICWmNLeqmk4Xjx
FmEVW0Hi82RhOkursX7UlP36YlxVybdcsMFuR3m+Aipvc7fLcEbnOnjfLv3+zX4h24UmpopVzIIs
OsgqTVy4U2URqmpQGCyPI7sfJ+/agDIhaO6Ma+Lb8C0rLj2Fgd+ZXd5MgzcMYIipiiVYOx1Foq2b
1MSvJEIfjwyYWP3aJ7Lmf7UTslXccjKJdZWCvfnlqXprdoOpgGcRfnN1s7vS+KR1Ph9+kZhlq89y
6uMNc9x2BJZjPmAZd7xAvIGFYwTTzeTpN3JBKjgY6R+tkylus2OmxjzrIdCu6MhsCONkbt5U7DWC
tl4R5T/ZKG0dwPhKrv+GsU30CshvdUaru31taTuvAiOr9gjQZSJKP5sGj2P+UTpMO1mpLePRH/9O
r5v7yGSzj4eCOjg8d4lfxB2Asp9fJ/Q6pFkjRBafyShXYLgTqDmoxU6CvCypEll7AkaT9YgZYEoI
xkucXXAJrbpUEwQlqBCpcZIMusck/oRq7iagOn0KohXWAEBRjtiBu9PpvesFRsfhgTmzxkGJ0kuQ
TYQUQQZ+CT0LGBt9R4mFzrm+krLo+0hcT8NNYSA4BSjmszhbarPf7/8avLDlXBKKKIaGmcTQVA4E
UIFHLMVdC9CEX2KEMW5xKNKW6+bil70FY+Tglp/O3pPp2RJRzb8tC2n7b8lyR8tSwMSXbVP+YjiK
BqHHUqz2GbNR8TCsCMahyl7IhBbhY1DhrO91DDn8rBqtKYuHSICR0x+JQ2+c6rakCvwd0rNcuPL/
Ay5b8vZLCSk8SZNys8WiaUO4Crm2G/5hLMSgZ3XPfgzhO33shlj10Qv59DJf19baarv1n58i6RFM
jt1pXL5OIqPrm7wO5yeiITFWrEkZQrTjBHPr9c7O7vyYcJMD5unUbDot/eNQGeV7cGt1M5TirJAr
hQVtfhCtWtzAeH1vWJQ8SDF8bFfgnl85N9BIq4YFJywBQ37IAgarwAQ2qtySQSF2Fw7SsY3zMuDZ
Wtq6SexhnkXllk+4Vok1KfEs/4ATH9eU07Af+rd/WT4BwYF1Elxa96akUh3RvpLOxfir2qcULUg2
E+bNax6JaEwTxRBOvV1Q3p+YB9p8JY4AuQKdVthx7EQlmCFXVGwn05OlJ3KkxZb/XV7yrbwXp9G+
y2N71qS+Le7YZ2igHeYNq6jTn3P98nKRblcuFhU8Y5rjVjoWQlfmSQXSqdow0DzpC0oDUZxtFu47
8GsRw97cjqczLe2Ojtq1U8KMoOX670lJ+dARddTxNwTG442flU5HE6IzkBmMBZHG3ucqx6LNrfyh
OOS1wmhetnWMUI3HS5Nl75n7tVQu8DtG2KTyL3RhbcB9VXZ1gOWFuaih/KTnWd4jExhpKnTYa58c
Yy8hVeT7WYa2rjGq6XRWQiySO/G7A0HIY+Ci0ltRk0Sp0bTss3EZgFx9Qi7cfbaagSdCSY6bi2rt
nAsmasgPTi++wM+zpMjVVVnSIlkyKPBBGRw7/WHMuGZQkg+KIj3c+or5Xw4ZI1QOEDQpxpA0urPD
/SAXpfyAHwiJLfnMn5z1z/diQQfoDi1JWi4G8WmhMga1DBhvuw9UqqAMbk2uZ4QKm1nFTJslF+5Z
VS216vaTT2NQ/tRb9thkpp4YismJE/KDELnUxjZ18xZgofl7Vw/0TjfBgY2nwWh1zjaBtYZfV+gq
658x+OA/gpjy52LR/1VPCsWJfSTgxA2pcLw57QYNAApt1vjdT6TBhA4Hl+vN9mZJxslzwv2ngri0
En1JjilVESM/n38RMmkfokiGUEMohjqelWGB+rhBxt80HmyR1svbqMlTH4pzyeFPWLVoCX3OUiGh
OVH1Jbf1T4ErDWupa4bTU+C62nvKvSRRKs3rTa1KiKplt0JVLHuo5bTxN8qF0fkvhDU4u9QzaysW
WTs4720s0IadZd4HQv31xsnGv0kxVEKclOcdfSrzchobmtNxAWbEP57ZGeibc01oeu+XUpAJyHTw
FDXwQrQUW++mhfcFXX11QXzptmkLZbjGsaWfTy0zgkleZdhBkcSFFXkeC9MAVBm6BMA+ctqfFIQz
vCC01ugFNGP1q3i0q39s5f7dFkcKqWliI2SQOeVjjILDhVItvilthIKb1kUF8/tMMhfo7jL7+Q5S
wXgOTunLLSJojrkl62qQ0s5cWaP2B3s+pyl27MA3oZBm9wCuRLumxJOrWba8Ur2cStOdxVhjXYjo
reRVFtyoyo4Xgjlx2lnPKELCSzxrUEhyVFmx73zUPtGj53N2IDe5k8m9Vetp0Jxp7qTxUkipB+BU
QA93k1aZsK/gPw9k4dMqmZgS1Rq9K7SE1N1bU5HcqzutKmhfpGQz5Zt0qMN3jorDXFjcIjXrXYWc
6FW6e9yHn30huJ7Rwh9eM6lIAUAJYeSmuo4I0ds9k4YrZGzKKssep4GdPeSytmZFfbaQfZOXBfR0
dTvZGVr2zKHQ8HcrXZQvZ0v4LIvub3V10rW2AipGY6Ir6RcmXDOCDoN+E94ItIWvnaYE80SBxeog
7O/KLm4EG5JLXyqnTSiYYhHQKLaZq57PoThaVmtRJ8PBEo1p89oBeMOh6hkdG3JadOOHxOhsWxix
4dHTlNXwyQivXq1eygjt2MkmGaIcka3dBdhGXHTz63nawIbAQVnn+fjMjdwYUzQ7zuWTnWzyuMP0
kzxBjOb0sYiB6S3UDLjjt8mM9znsOZvPewDLaNvjaXQ2sJDYntCcLyWak6XVw1P6Ln/hJrPD0Lxh
tPdINVpvmzfl+g2B41MySWqO+obZz7/SeSl94g4uX6EIZiOCz2/1vCcp2JhLrWbW+1H2DjXiCbyl
6/GIc/AZFBDkx5ASZ+yyjJ5oRg7KVsHeRdMyHlrhrPLkcmwjpKS0btDQvnnvi92E5Zvnq6H4XYmw
BRcGu4zj/Vg5UrE14uTWBoACh79Y00laWbiDGkCAoABR0KFmNBiJlCs2De1jhVjWx+HPokunP4W3
3LfpbU4aaW3MuArs1tI3Rnn5Je8bb7ywsWKqUtAuWCskU162H32Eett3WPfgjrdJmHKkn0jlN4XZ
+wLp0I/NSDBC9A9XO+WLDFTTNfHOr44G1U3TX3n9PfPkc3+OxNw+CvjbwC3fAOAaQdxLAwxF2ZqA
56BcRnqKZrjAAvgds52jmNTxd4cOVdwkipVfy3pf+1Odz09oERXca776L3UnUz3Y93Hhi1eC+0q6
NBfOiLbiQEDrwyt1g1oGds9GBjpGeLCmWXWHUmrygFJDyAQ6hIQxZHTvq7ULy94KM+TPFfR+GmcP
AizdIETJ7+CkwYN6hNd5nCYvDpw+Pd91ZHC7zBBfk2RxTXxSb7Dlow04sDrWEptP3qKKT7PkfIsm
cSnJwNHS1iLdMmRcrAZcxxuAf2g87W99yecG3+4sC3CinOyeYivUnypfOURg6iyPfVFKDZSI/QUF
TUZRkNY2AlSxkpyfo5XXFKb0swpe/0DfRhjWv7A4EIsyw/4ZVszxc7NG7QeewIe38PHV26RBUooI
XexO/feUB3g7sgQyQ7+BK8/5PFw6V5LHxfEtaXg3vQcBq0c0wIOYw7zaLIu9sddM/nrExSv2EUsE
tnZsZ4Hgakz5tB6DbjlthKItrabN40GgC1WM4aJqmKerscE2xWL8Lozzo7Zk6mrhMnqQRQ/Ctwun
r0dNEM5d5jGsZ+O3ouv4yBzkD0rHMTF9jg66D6mlMN3KyKfHQDqP9nUlI9CFcdHlL+Mkg/NEwEL4
1iEWyqORiyCteHBufZ+0CYcqdY6dONL9f/Inw35w3T56zKDg7rv8wzhKz2A7ppE4yFg9HJsuJtcv
RK28GZzSK3/c6Ihm83Y1vT+bPGOsp6FtiE/zq2yR8p+/MY2ae/U7RrpFkOCFWdVVmlIANnuU9n1v
2cafSYabrRDlZMKv8tO5nTaZh7aKSuoEGc82dulOzFHtI3YeCdIJWofKkA/FdcxYJibG7h93prLX
qe2uxHQPXQIP67qYK5IQtCoEybYG7FXdvvLjI6ZpXiJa7IOg649ZcMyKVnZdI2IUt9Ma+MTZgwAM
+YuVq7FBjWQjixkWNfISttS1ITO2FJrVHxSVjA4QDBktGpf6wGtFeEyig3t1JRPoMi80DyOFJjKF
YMY4Zz6NroI/IuyHLws3s8vSMljdYmG7tApBgsaC+mM0QH/d5eM+0JIozcaiTSnS2wWL6h8xsgtT
Rx30sEVz9VxHAZl4VlHCvdYnoiRJ1klL09o51rT5RgBuTC/wDjKznTljDEWONAy1YQKscdUpxfM3
UxTmwXjcgk+BGlXTqmyxzSR/4S1rSzKRGcL53kgefU/a7ivHQ4f+1d24ZRwvdwiI5S6tUKqt7xLH
pB9cOlu1a3CEVt0UOrw2y0icMBPgeC+kq4ir+HVvUHNmPSbQHIj9QC0S1tw+yqmXF0p+98DfPkHM
1v53fMJM18uag9F1X7p97EVZ8IUVaRuYAymcIO4ipiveIpFAmX43piqMgSg4lkrzFWdBveCMI39X
ZaKyOZTzxMXhn/nThm/aHchlAR0XeAFM+d+u+WPE22pkRDRsbTyuVWcN5Ag7i6apu/ARfnYX8z0B
dmZMvFQQuwiBQwNWidIz0WgCWYGAtyTWAvL3jr+tTqz5GEXDeCy2anS8KZ8sQEgYwmkvAqslThrf
9Fn5hbJ1BopC72k/jeYB2CmthJx+DjSf4JwpbR844u9aJ2q5lHXobI+8KgWbYciyPNi3FoDZhgw0
cd7K+mhWDkJPblze+DVxqpfVgz1WYTEDcirH2UduDdqtrzqkSf2w9xEtyjRYlXTFqm2d3as+QYni
ZFkkCciD0+E2JJl+frpb/E49QWQov3Kk36uZvjjcr9d+BBBoJcs/HRvQyr5yRxnWSw54XxqXG54m
QBkBhF0vavEBWkmmeAS2UvaPYCvZ9iMWBeVyecKqYb/WtmPcadqBj0gGXEEvcC7hpQto6s/QGz9X
GNoWFRqiqHQJKsmRtkibsoZ0WKJfYASPjZYYfzA0V8y/1CxTqIgx5jYz108n08W4qW0dckTUHNgH
TcdX7H7HuCxtrSOvMObtcxPasABvIQuWdNdqenH3XXNuMElq/dEyNx0bqRcVN83G2h3Rnht+7kgA
3WepgvXXCI/W8O3nBwclxB4fidcj5y5s/MbFN5QY3a1hesDGXThgtQbicV5fbEGTmOf6txFJHaFd
LxXlu4lxzJRpOrsr0fpsVNUCI64/esn7l09q+ZEIBDrbICe8gBwSeYwh3ZSdY3ZoByve63n4dLY5
baTmkxcstPryKrBA6I8AYOPjo9TyUy50Gvs82X+BwtikPWQzMc6VD+InBT3IGj5xgEqXxJeXlt6G
TeDdL8IyXiz+CUCJxB5LNFB7apGGKGdobi1nK20NcFjBOJuMnNgy+RPbBOWbS4QnnSYZ3XIMb90q
2u04K5Q7aiAe9GEJkZK1RPHo9WpM+ZVLLhiW3DSPlqKFSu9nGR0uR9Rq4kyInF7XU5a5CPc+lmsn
3+yOakWnxv7ei4zKe/ARsvBHcVHefEA4/MyPf8+axlaYx583OqIXHATJ4/PJksSiZSGDyaikc5Qn
GP2C+Q4YPw3viYo8NXYXt25GomaM2MUAJmCxDLF/kNCmh/NiTGk8la+Zox7a2SpM3m7M1mgXaGJm
p+stf4q3iGZ2sBsMTmmwjR8SURJpf4zUvBipAPblD/z09uktth/OXYB2Hc6ZUrPDealblkAxJcvC
tdHnNLTTQ685Fkf2yNuau5Qi60kL1al0NrM77mgkyYcpgG0XBcmYQ32d7GkkQb+L5Fdp2pvlLoVm
BtjOrR5H78Yi8oOAHX8Se4FwnDnOYmt430OwNdauY4xeMHkqYXf7OYcH9VsUp3Wkz4CKC62A/PS7
AalW9DWzuIrCIy9+A22emvWZyI7Zx76kzZ/YTmT38jykQYIWotepMkkztGeUmelpJHtXxngB3kQ6
7CWyrzWr7tPoKiPK9fQNeU2pp28uWGVApv/hXB8WJ6+lgDCrqPhGnuy8ecuAJ97CA9PGbXmQsEMB
2UGLWu4FuFDQAfH+DjhjrJmNr+SOMf6fxGr5RFE1NXEylgs74P3N5LlURKl7tJiCAuqjIrXMOkg8
sl5GKQFDOF808org2Gc0TOMKx00lC1L3UuTvkVm+8J/zhmNMlt+MUP5zWe+wlwzb2sniu4rFq4U+
HsJVPZHOFmfplYLV/kWChU9vwI+uKe684LR9KHCnb+o3BqSsyQWmmSuuKH1n9k+oa/pZ82Lqm/Fb
CdULUhx3eEyA8dtQsyH4B8+XDUGo6FCUoT1ddEsyo5igTnInXvnmcHiX7DNC9v27nO5gSm5VBIva
TH+/8vzW+EAXx0+B8sBXNMNIAAIBJBXO3XLLiFLpHERSJiycOr341sip6fy09erCdzMS8YGiMRo9
FuwgyNN0bR0Z7Kx1sTQx9JUvOfPyBNXA1lLGUMny0E65/hn0stu06hD4epziTjsT6TsG6yxNWZvV
lAtTaNLHArNT8fL0s3k0/UpPSCJhtXvG1BN5q1YpaUt77geJkKBQhdGamsIuUJdw9tScqnLR9GVe
xRI/x9zjU4Ji0MYLAXaC+hBr6aXqiERBQKXOU8qSmB9CWTtKiqPTlUyNYv76RdyvuKkrRz/Obqi9
VHNc+Q4TuUP1Osc2dt7T2pP78uadNn5vaLd7l704EmSUGk0ZyVLkKNDUweK4CIbQW6VRGcdCxwBP
Tqbpo+9q8AokFPx/fj0L2MmHFhEM/CKhjUDw860DqkhriNGmmqArgw3q1HsDRP9oZb+6hiPPmvMl
4ooXwAo3qINm7sQOA8hCH+eFdTHh3Z0Rh6VbPS6vbxH4Uf6bXvH8xmBDm2qBlABH4EmyZmJpIZcm
BvwPQI3zpgY7UgJ/KRfUWh0+epGvPChTJ8bxfGyk6ji+tn+giNwHt4HLD9mH04omrBet2KmpWn07
7fDN5kuENAEP0ZXQchluMnjRHhv+I75xnnqFprdNHh/dmh1k/twIG88yn+Kn0WbRopUd6Paka4F7
88fjv9FKJT64Rxe1EAtY7lsC8U7Hk7y4hF6veGtLLhku39MmxaS2Qhc6fwb7yRd/Zor/k/LNt5Sc
3vLBU7F1vWao0z5mSbJrAsanxRoA91EfgyV4GqwXzH6AGtmaeyE9kReiDCvAlKlPmYa0QomhxKze
UsEN229x7josnCkJ2bmbOG2AGGm6vvBmlXtLqofM9CrPmajFiIyuASNfu+i5h9J01hq6kxw0/zMU
6zYqBnQx+6BHgJxzvHjOk7liWoj1lBKs6iqkxqsqMdMXNu4IC5Jle5eW7pRrrdXjIClGa3xd+epX
7xBEt6exuiZkYShGVfaH43WY/jRc+5cQ4JYd1YiD6Kk+n2WUg4YSUISfNt0lV2z82fcZK/6XV3hX
n+Xw/uLL7MYVTQVmS/7bP6DsqqZX1oS+b+20BEa12zZ0WGl7nb1A3y1AfsRkYxyPsgqDB8GhMHnd
ec/JtHNKQrajBxxVXtT1Ekg9WEdOgT319gO/pezXY1ISnvvd974EoUXlZv3J3U6OCIhDxqMAY2jF
hSW8IX1i+vv2b32XE5rXjKxNPXb1hO+wMWdeAndbkHOvJ0DHGSMp8xp1vd8bfpzrBPPfbJphh7p9
2o1jo+zKTX1gVdZocmK1IHu90sjj/rH2iWHFomIvLrl5eNKNc3pbEtKJtZUhMan94vNVKDDCQWix
wFsaldWkgrPl2BPHINDnBibLIg83o7ROoyiX/6Jeo703l4eYYedVrl//zee6Pg7wzcMhK0pWXfFg
woLkcFTS0Ece78eaVDG1y6aLOZI0vjGxOVZ3nN1+KWbyZVcsqiXbLjTsswEK5jbTDan/QgGKWI7s
5gulUHF6Tq+UwPlbC9JJVv9fBT6F61pqRSPSgeg1TFs2DdWRiT8ib+Zmos3FZ07tIbFsYzOQhbg3
Iix/6JzbhOUeAmAppgNTsObpHJgenXR6V8PI0CE908OwaZlnFBxpjg7vLp7KrVGJAQfT2gG7gBRB
VdmN5CllP5RQXG68AtSjaO33Go0J8Ze7fpi8rwvw06G3SGB8b0lrmVENtUf83dBwd0wETAyqz0gi
kg3sHDLfW+3fOzM6+xGeH8kQMgk55CSVGqUbN80rqGmh86ABgos7swdu1wv2jy4pQx/k+/NhJvxY
2khmsGsoWyGRBl91i1HjrzIqppJ6Gh93JkVNukEowdQdMf5lWKM/Xu/FRmwSp/Wb3SIHwcmDUL6U
AzTT4KuZZEZci0W+C4TVe9PJO4ACmI1AXMjMGWkwdwrEnPxmsVcvksqDzGUBvUAlQ9i4MfrQli5N
LeZBnbLcxGJnsTS7Xk/XwlA/N/d9NvhNQUVhXj7HvZ1Bg2zp5bchG52uXuzXplUqaiSSpmcsWFn3
Pn3VCjRNVfe16SzUwx3+n5e54gSB5fEIDLs+K0JEKUxdf+FyKGepuX/QymoH1cohI9ntdndryCnN
PhoUq3WaKa3L+Ce+ynQCwPGsK/QS9B8xluX0N9ciddHPzeIPndTxL8ruWFUgsFk5FPAXD82rXD0t
rovLjZqTFvThftWmi9+b54nmUm0Q5bEcNoapDnsgKSbEzbSlspTudJP9hLM1XgwjCoy+cyD551Vl
h5kqNPEzZe0UNXlJ6bcBrM8NICj6upuM9oLQfY2VHYyt2VrcaApU4W9dYRcayuPU0Fr6nWBHkplS
9dupfAHZikp/8dEE2l5N2HK5TiCqTfrkzeVSNXNxihRVgxkILYasPRIMF+PqfnLpFUYDtayBxIzs
7E/5PJ3QQhUTtABH3PkcK5zeCFLLrH9fQ4P/MofqL6MowX0eB3dMICvl/ZOvoBXIQlh660QTD587
Uf6oeFHagVakKUOq+0xLK8TvqMakOqyzHASdGjCDAUFDmEORxf6irEz8o7E323yjh+MVP+Nbqzcq
9pGbC2RcUBJyiPFPjINh9QmPOUFUC3SFKWTsK5FoNXNGiSCftTMDBwOrda8JVRdQveJ7FcqYBrvA
p1CLHX8c2PmmFLxzE0lidTOxzrfvustjLZeH/4hbkXqpHkaJ3+BrX2+UWdhPg4YrJyz0WsgVDGcp
arb6NQl4D0OiTUX8vI+QnWYgQ+28TlBB4mEnriP6FarM2hbR+iMI0PCtr8pIS9H3A3B/hqi4rYMn
lWrM/ZMh/6NIVtp/9pbwg6U1v/XEb0iXTbB0sxildFWJwKzUg3cggtaJth8UaD9VZTEOpluEXJms
UqruL+g0/XnGGJshp1LriJvub9VXyfVaYPKIbFNse+ZqFtm2c7rrLkTMR4DVQ42nVJAeOw8RmkyE
Jvp8eb3Qjnao2rq2NhZHT9P7O94xgZdr9jHXaM3j6R8sxNhfRc54TeTG+PvGZWRNGi03hDVzg6Bw
tmpzfFYU0vstyGRWAQAlPxiHjIS1XyDlvFWYLaZQ2e/9t87y537527QjuUJxNtcrzKIXsXy7jYyV
a6KkXgrT649cvVaJRLfMhLNEe6D6f2fTXrO1UI/RR+2YRZeL/K52vBBCYw60GN6djzrgTxdmS926
s0aRn2NA2lVc0dK0VdPVMnqFDTRxOUmVerKx38D+nCky12s5fwzsoo/s85qCMvIt8siZoAe7OUjM
ewb+LY7SG0s0HmnxavrIEzStKvIiHPsQLqGSMXBfD0ej0NZuVKFsshQCao62sTuBC5r+R1m9N35l
434e/6dknxjBZwX5TyEb58so9VfrnR17eMou2nbfAyqsaXsqezfyVP6a3kJ+JBmP1xiRw+Xdynqz
JZX8zErd02le+hdt3C1UVHnp75ZH6HsRd/ud0+x02KxqWMZg10+An8d/rWmFpq1nAtadvqH5OEKo
9nt9zkmx/ZcaxTnSrqLhEaoyIfyalcHol4+i7z52c88b3M9/7hZrmlTosxNwJ/uhOUngk5lITmyf
lCyKbnfWB8UCh5KeNrUnbQe7jkpoJqugRB5LCQBwnvj6ksRpWWPAbygUMaWO7+sNnLBurBr1b2Co
3kiJa1TiSo8HdrfnVeK+QuWo7A89KHvlsRk1j0/Wqifsvu29g0eRTKFuMAmho6XfOzLMEFd76oG0
fqLQb6f8gjxfH3TdSqCCtBE4/2ZgrzOlevvTUBg3K6XEYP0bR1sKPLeIGaS77usUbpB+l/uFtl72
iUivpltC1TgH7P6jcKN6sjqzBlM7+CAeGkIQPxUG9w8ngHTds2aJXi+YJoe+bWCFX5Jyej3FK/9T
u02EJurZ+iBBNn/4bALtsZ6E6/qQSqiE1+UyH5WCtfb3/MuVa0VNO9P0AUQex8m4+HSEHVvPmcED
S2DJQhxU0HSW3/vlwh0Bq3OW/iDKXymaeHakDPNivqWmG+yBEDpEh802slerKvQp3nURC47m6YVm
oZ/jAa+SDq2ibfI2TklSJiKctaC9JfBouZhiT7qyg5GmlGXRoiElETTvK4M7wFTFBd/njTIib04r
Hh/ZcDi8QpNgOY7YtjMZCv8H2KI4fybP6K4rv0nYuh1E8XxK5xJONquLxwXjHdg8lv69qA3CdWm9
rfzlQrY3Nctm3f/9jn29b9rfWHWtCSOINR3wqT9+uazfFTNdudXtDu5cTCPIgEsw0XweGfP0YhiQ
Q3pOjlPtVjdL37IASFSnqAISlQb0hcI5el+hYqcLkq9mGJztFEbly7tDWEUfrgIWOK66B6NUkQSp
lbw/Fyi1DN4RFBJHx58qEUgyKVp7olyRlbPbOWt+LISRg1iXeagCxY10qCqJqzrJJ+CsgrBg7Exj
NCloZlcgbtDtDlsORTHEKgFZAQb6FzkMgiMrV8F4tkeT98y5oCLR+dTdsD4stcUshWk7muIGYkKo
VY/QpvRH+jMFsQnWXDMik21y62vWNeEzFibdGjvjwZiUuYE3zQwaU0k6MAGHPs1o6Y/ML5tdaAeP
GyoakdxRnMK2bCgbjLnPcnbJNHjmLd6xndgO1+p5OBGwExDwgkaSEwkxBR+iQF3mlv5oSru4sEYh
tQvmR4+crkmYJFsI3vaTbzoVvY3rVbYRexPwM4sjfcROrHy/XJOngTT44ElXI3ksFpuguglrMKXD
Je1cqsLz4hvUwc3y4WrRwMcIrLkY/QawaFYL6nh2R4SVUeEKOSYO5RD5b7pZG5OFsAZd4bc23lf1
v8YpYTFEOns8e6AwDyDH6TNojmZ6/z5e7XJWv8cWGN7+TMV1vhXFMj0FCj4EJ+k3CjvJJ1WyeMds
gl40+0h1XsM8kL3sKBPCtsErgyjL0ANfqDdAoZS7j0WYGVJKFajUWu875dosKPqL4GGxxoXuYjRa
wBusjw3XJ9gIiynx0BzQLLQwm+LW0UKyjU6o0m86LcHUjYRQd0bHNcnHCobzt/DSUBRhjrsJx1N6
zYeXfmhd6Nv0cowGxOok5ym0tD00Kw/Hewj/xk4R3NX0pqW29iq+nlIrw6lpkOsmnt4r/+FGDu3i
qtuc3YkhMzSLFLNv/pun7LZ/q1kxqJ68DJ6j2Pe+wwrbVKrdD5Eqx4g77ahNRGVWFWpkjMRDLGY0
4EVwQ3Onur7sveOz9kd6HON/a4xanHM7Rs5t/vax1+TIB6DIvzpjtu7vQYjBW8V7wnqphulLQp5C
tG+auGgju/v7Q0t3K7ZYd2NHTceD9R8pxEKaFKQp9C68nu8FC9eFPEtK1DXcYfWp9ONamp4EeJ0y
emndPNAIjWinwr8wX373C9z3dke2gM4VBcgQLe3cYmhq2pVYPnJV5QPKnf/BW5I9peXCPSOgvUIq
92VETFNoi0Hu0sAwrgIp42875R9owj4g6D5Rt9me7Gt+PIzoAsCgon8SJih9sDUtyCpGL8kh3cHW
atG+HzD4XOLQcHYNKOXycUPNvQJ2SPBpL3dS39n8BD6xLZA9Fus3gEeprJ3dPwQxg7J5VVQUWuKf
5RtpnGxgWIK4FuebcRAWG+PaKcczqLlsZMVXBkoZBd2SOkCXhy6wXqKrMXGSPY5Y58PfWJyvAxXm
qCKGJRU2WNKDnvsgE5l7ZRCwNa4NwRVGqY9u7Amwg3nODU9UCBy5KLVqtMfq/d7j7Xrl/NY4f1+y
+vJpImanFK711OxQZx58+h1ToLKIKGMJGy9sGWaiTFpdTHYsad2JDFu/B03R4tqPvtXroGeN8KWF
d3FjUc2Yk0lQ2z/aWbTKGn+geUOcjkYo6+JXFZZhS8MvdajxGNIN2faHYfDTJGXoKYBHYhOY7d+3
t9Jv/B+w99J+dt/9CCjL5D+gaOT+K0gNv6jH2fSA13R943fRdCR+nPfESDyNeoOpH+VYcmArfVLo
8AHNWfdSwADFPzH4/Gd+aJKLbELCdX0aDwUcrv+S+UbGJoeIxcPcdSNm/PTE7QoFfHQV3cgmPDpz
ysls/wHFtou8B41xNV3oj1pegVDgCDvzZVVjUtueTvpv2OIP543qy8I2k6Eytc6XlWgQCnhV/3hA
XSjXInR8+LopleWR9+xxPnrWl78GJOTMyjAcPfbxNupT96jeoc8oThX3ki2thWTiKg9bSixECLOR
aNXvEiEYe6INdPUARNOOqt6lt8VLvRy+LJoJAqrE7Ls1cSyKMS+rEIrQxiTTdBKAwGsCx8TjMuw5
noFpAictWbAYMB57c7DRykK1/qkXBxKDrM3lkfIBZpBg76AteEtV2ak+SMTR0rdcIlYFTnLZ6A2h
kSV+scxo19ccz+IkYePxn34W41dizPbAc73Bh5ghGNty/q1GHpIQaQFj6YuydRUn8Bp2QlBMYzT1
2uF6AFhs/4P1sPJCUM6EwDbzvxujClUA36bMjbmZZVf40ERT7/8Txl0V5UWj4BHU3S8OurNloJUJ
dtWz6l4yLBiOmmkzWfdCeeb9pU13masdMxXo9Nvgbp/n5DcWisIKtpWxr/8L1fF2GQxMMpMub3J7
bCygJJZydG1H9fVfzA0LwodTVhGbtTEcHthlc5HCgmgsBrEFbrkwJxTX8mLjN3wgD/xpEaY3f0AT
5+FsezC57aV+KBqTC31vtiwTQKEBGCCJgjt0o3tmzVpf8jIyyBQ51Zk/42vvC3BbXdzjCEtqDXwS
UMm2iRkhdPoMh7MjCgy5R69gr2hzlUcnmo6m9H94M0/qJAqJgxoWBv89iOaFH+iyiUX5kbB0wwCp
2PioScHYBodTRbXuY7Qj5vxHGTyVMoi2WQPJCJ+wm+NZbiM6Qvg4/fdqNLb0udhpM2EeOD7WyT5U
DV4TcwGzfn0bE8Qlin7TwJJpPqBwnomwXw8DyPCK7OvndDc7VlOu3TyZMfoIK+wkWfsj1RifzTu6
7k3S75+e+RffGmgD5Zfy4yv8VoN6H1EgI/WdgOgDbsP0l/XQqeV8FbIs9dfscdZ7D1rOd2kKhWVB
iF6h1c6YOz5Elhfcflnb8EMfCtGrkygUeaoeR/JDwdrVUrvFcR4u8Uq8ukfPD11fnDb8+FHhMDDl
DhK2EUb0GT/3eFF0kjDQevIIT1R3dII0jQRrJ+phA6uEqrmo5a0xGz7LQJUPao4jQHCnCIC36vIt
kUlYOInHQcguI/R6Zu5HNu6tJTMhCf6JQ96k0c7KUtcNO8+kJxF97W8fEq1YJr3HvqKBxU2Hl5EW
MmxCBjuo9x0uSg+1MerzFWpq+4uLk4WuWcuszYsY18sisdICQFMuAyocDgskA9p7aJaUF532zHrJ
MbsVXf4MdEM2A8NyaLT7yt7flWVFvydYyqrh5R9iwYn2FmKVJMVZB/Z4VCdJj5e2J4BcLe/hl1Te
dFZnMJyV2Pr+xJrxbzSekNQzLaFm7Vg7WlZaD6cNVzQttYSDK8gPLhZm8ofi19h3fTJTdloZ68+C
94uK82Hy+GM3UmR4bDydVNDKH1PKktwnQvl4jPoUrGzyC56Rx++u8uR9p88pKNPvUNkt0+1fIxBG
eV/ukigDZiR3lUQzQJ2ABUNSvMCyMfRxqEPl1RFKuwwDB+sKgzmQruD5adS0wpqtLNbv3L4IJU/x
1nSBtopRtmnzBvta+RQKSFy+X/1blWjNYiQXIdBAq/Fcg1F+91G/wYx8nv0Qnc4k5+hxFCCWKAES
Hum4beQv0BMyk06UOw4YtJiL81Uo8jeKGdrsfIzEE7IQNCt4rXJQVfZIN946cRxuqxMvDapcHHuL
I5zSYdXd+OLjzgiWgARKSNKFoNqf8Nwi1cs+sBYGakp/Rx6NUc563GdeXTTxfNWxBxBD2plKD8rW
L5YzVlwc2XNsaO7Ww+CEG2B+7m3vNfUDusCBP7ObW5E1x+6dmffTF1yp9feTE11bg3HN+aVlAufM
rvBZrC1fG5h4nYJNAV5RR/CLGZCWdE+3WvIpD31ezhSPJPqwJa33vb7nR2sYM7JKfNjEi3692BZL
lRcXhut1CVcA0URc58amCSzg2NTjPRx13VVms9D0m29GoBllR5N+mKYYE4Df0Sh+hTcqaom3ioAA
EK8jNUQhcaOGa9OoiiV4N8bbaGfwHlQqUEByKrs+9xZqlLeVKAd9Onh0jNwvluHgNk+1jffG3A5e
X1I5Y8AZgykyVuiZxQ56XLjsyC/5QwwsODySmbMRn9UkQZARDIxUAK4rxMirra/GPFBX4Q7vp32r
DYieuLqRf8C0cCUahzsuBx+r1aoFYg71D4Oqf4BV+nLtBvL7+OhwI6QlzIJcsjGCwTUulVSAxX1Q
lvHha0GyasHYekdx2+TkUkU8W3RgJL/L2H5rYFZM505A1aBfbZLmwdvaC6Pf2HGjz8qpXAsdLdkZ
elOjzHINlo6Sn02piwO5iOA3x4Okj6JLqLb6Cw2wN5MfuKVS7pu06QnHG6yHBS5k22WN4IDvDOea
HqdHV5Gnh5MtIXglLSmjEuj5xN16DIS9c6UaZ2uSVhtn+TnJKcSpAnsHtdF5BCfJGjqwZ62Qazpl
5Q4asBpIHrKzshoStO9kNwikKR3YnR4J2G3s5+NNAsYlaXAfnCXYnk3ygId5NSkivfxePr7cBJLn
Ubjmu+iPlWPk+oxWjCEFpncpiO1j/MbQ1qiea5VnYKjwao19gMbro6kWpLUeKT+hplbU7rLtJpT5
k2f/69VML4h4i5Ya1m/ljjQKIACT4gKLtMcxfs8RbeOx0fE8Iw42S1Ao4IJuVIjV7b+KwfGJ3dBW
pOKzq6+DYxZ0t1+c0l7yXVm2EhqCyP+7kxZ+5y/wJgF8dvwXxqmrL5V0R5761Pj+sBh6/k8WBsQ7
fynG329q1Ds4cTxqagAMITqxk8KmlGFGLkDECjH4C5L1jKZXKPTczSiNNUUmHSsGoQOyZCQP8GOY
d3A7+LKl+gRGoYbc27Yxu+C0BJGgFjoYHYSwyKLLjk6bk0SKYNuD/3qqNeyuO2cImaefgeFO0AJn
LMfmNNLMYPwwTfsvbs7ZbR/gxJnevEnvrzp39Q076nu78MQXGmnTKcRMc5VCuZ7Zykz1qKpQoi8T
egywRuA1hZnJn8rVDCopR8jzKQIpOWE9C5nsCmtPZz7qSiVdxi617cdRNe4cuGAJ5AJSiDiDIhtg
kMKAsZ30eHUaFw/SJs9hLCOnHWCphZxZ8COHY2HxtEtHDEbQgeJgRJ4vgRZcY8jah6nZt0ee3rQi
lWeGPTcnurFFKhLDKFflP+fyEIBkpCpyzxrEBYChd6qoXESL4B0QGFMT7IGkRG065loKTSRiTBxj
/NBzeFsnp6ZWuwNx991P5Szhvu/Lesu5GyaVrIzMFI7f7cZoPVEu+49I0yQMO1gmA9ALhIRjYtr7
deQBziySVCbT+t8zKc9Wz1cQrPFliAB4HRheDYxVqy1AAORdHXdiePOX0HI6/Exsv01Kybe2bXRK
QuxkJURw0t/ozwasNC8U9U4iY0hg1gS07AtL3wQVL4u50cyDv4Ose9SKlF2gPCH0FE6EaLLJT9+f
bqcTPqWnGkyzAcRX7pjkR+jNqb3gYtBX+3FWVJyDe5L1B+U1+VMRqdsR0W9wLGtzuaU0YDlgmt5t
P0vfGSNpPUKV9URaid8eZCyhjcPS1FoND7zYmqbkJnirBdJjLnRZfEe1CqrQIRS0p8P2IeDHIgB/
FDpTQ5mDMsw121hTEskQl5EkSafWhsiiBz/6ujeJp8OaX3dTa2Hzm/I0vM9TKZyB4GEsfDefefEl
GsdyQnSj578A6y7Jak3YufOts8nDr7e6JZ24VoP1MWhZl4tvvGiEb6F3gqNDX4WEZmqUOHd+3chU
C7FEH4A5v1qqkHQ/OUK3Np4SGyNgYwLmT90dlGkgOhFWhcsksl79SW90kECiZzwfEB3jnc+qJlXQ
7KFeF/nJO8HpNDro5Rqzor/btQJtBx7t1X5H+iOIduFllWG2SK+t1Q2nWRMnS2K7yxhS+MoAkbOr
Jo5cK7frgHQgQrO9WMO2xNgx6UJCQOS6yq7yZ766mzNgDXafnEAObIzvkKFah5ZKnyDGKAVC5CJp
wsu7fIFl7gZ1+UmGM8IpZXbG7Ri8xYC5iC8F11w0eIpc/xreYyEKeyyc3zuujszLWdl5c823XY2S
rXs5ovsk/Wxcl0MmwSLusWUBRKDa7/Wg5HI9g1cSHcj05TtAklQCosTDHyJK2K0K2QiBWQblIPqj
4ubMddqKX25AO0M9vwDlZ7ZdX/8E8aUz83TWxRr+uhFCBt9LS1B5CrMKVtrTmu+fg4sdbxF/f/iA
/BcpxMBs4CKGr/6sAIjwR+MLgMfv2vIzjojvgHTNjCe8PTK0+C0H7KwHCdcDFAixQYP8TxHURagz
2YF9C2euXiubsKn67uVnKu3KNVUXvAagoSed6GIQA9lcfznDVOVvdDGt9ZCXrMNtL0wwq8h3VOgs
pfEGxNrOo66z6W3vhFGEpX57fRjMyg1lU6pVZQbvcIysT8UiWKRjOwctYM+EuJOV/BBC1RhukWIh
zzhmt11kL4usiQX+eQIMKY38+veHt6QqAYUH7N5dx/0jg5FMb8fw+Y3Q2uXDUsKZQZg2byHsvwkX
xeRD6WD8B/HcpgT52ZY42PwmREJroHE38pUo9Y7iHT1qdRlOjmKVNbZr2X3eu2hr99FKylPAVHKZ
NmIVLQ2rfoOF0FWKgRQippnTp5jeU2Y4Gfe/rrkSZ5hLIxb4f4BH6cp3+NyBydAGvmF+rnQCm/yt
pBVPu9W9g9c+99pTSYADVzpLQf6gotTs3pF0F66ISRW3loPdzBgD4zZlxJd2gnZekm+/iGWULTtO
uzc4ONC2pyDYIKEjqCmouiBKprKWN8v197mrDDVCvDOYAIjAgtMnGbSS8ML5Gxsu7wdXsrh7ZaDk
MbIUfpUiQ3f6XiqchIVH6krciIz02CCj6xrAbQVFEbE3P1IGfv6ffZprqF+P7HX59hkyb+oxmJaE
pTTLLAhaA9zJNA+EWqJ24iPF/j7NTZQgWWqE2nVCJuHWMdVAxlja02DtPdLMlUVV32HiHNvB5Ym4
cRAOA0LLhnX6mMggSvMZgNnMXL4aiaN65GUn6DFm95B1hWq0+dSdq0hqEAYx2F+VLpe/XLqlMAKj
SOGehi0uUhsaBi2MGDuMe6S5xFoEkRWU9xH7NBSQRQqmNp+FrA2XMNSBpm4Ca/+brd0I1V7f1ed3
g2T/s9lui1brQwvaO2OLqwVmnfwplijldaYJAfkiD1jNEPhvMS2DhQ+NDANBooMdZbTA1+rKVWMP
xn2ufzTYu+0Ud/pW3XOKsRObVblIlR2NTwH/yLiF07kw8F3w0emBYtRD887Nb/I0NkLdJ9xPJ7fv
wddVihclOokyx7YnLB1UZPbaUchFzatkneFqhaDxKEux5+gGA2lPD7EP64WICNZtI7ucK+B1Pt7K
yvWsLHtEBMi5kQ82rcCxVCCogJk7EdZ3dpZJsHpU7ywh+gqC8bNLmjG7Sjy6JXFjuaewxmrL61mY
rIZZ/LI9Y3v+dBcP8orlc2mOE1m5kPTA9LhVXbJcrKk1aNiEkhns2lhek2s28LKGH2Il0dL7ZYt0
U2bp2Wlp1XAaFILjN5nYIZwLMBlshvUTGWmkj94bwwsziotBytGZx8LkdW2bmFZe5fZ7DVcSjk7r
TpC7trAgv3P7DBZmJszI8Zut5u7zZFnhi7haStQ7U60yBcD2qtIVOrK6ltWP7Wf/1/SriYPF7Hc+
Ex6ACkb85+VMiS7QolICyE1vlaRaWxU+3Ei2n/cTixTdVKaXEhRNkzj6D+yCwO+s0PmFEnZTffaz
WO6aNpnS6Z/bFzOc9zgQqhvsemeenQP6WItmnwd3EdpXcYTXdZNb7yevQrmovpxCYoHn3PJtrzx+
rlgC+nl9y9NqvY780rGIXIiOPSklu0UMJp3wTFdcbfRSlV/HZuRXJ3cdw3ymf7laTDvbWKUJ11FB
nJ0PInzU1IsqN3b6JdUQP2ZEcV7Wft0ePoAazjJbLYpC5zxtGhfcpm0BbF4BM8wHvvF9VBrFnKrJ
gcy3P5coo2EvxJbwLmVHT3qYWGI7uXYVmKzd/K1NazlQe4+2gVzDmoeERS+jFjfcl4oULtky41+2
I2vbXlneAfGxdtk10TMs/2FECU4CZQk95U/SLNYdWIVUicqA9x5n+useJ9T1/Z50NFF+OiPyksIA
SaZvJcd5i3qyoKJ6J4XuY5sQT2yCzSyQKPZnlqGsX5nbV/gVQeDCkdh4HClpNft4MJZ/cUZLR1st
BFOKNxlrkybiYfgr900Jm+B6DVaepfv/KsEms8+XSVUIfyMby5AhYBCjYFTy0M6w1sUADZqCJxtF
hrcsymMBUmx5nUUqBLc7GPo2IGHHENfOYpjUfC7uzCAhN6AEH3eSDfafpBuAtV0+WWNHTlY6i7Bx
UDQNFPjfS5bHn+yCPRKDOGmmVcuuPpYDTVXyKfVBsIhcMgEPhrnxTlt17qJvyTFIusBKJnSPqePp
r+eNoLtgo3ZbM8MPedCWOE/acnU8+p18RvR61O3dQE18jEJklpzjSkZni/m107t3Ej2ZoPPeWNJ+
jGGXeO29iX/aUFlETy+XPt965jvImGkdKBwZ3wWFwq+FPbe89oESNUEJeXqLBJ+AseyHcWqYtAk1
/LGbvd3RTnWhJasAEUHxTaNaY4keQRbnMWKxOt6lVyvSZz3WyxY+Y0AaM0RjDyj0lhZrMcf/2L1i
GOjsdYEMrwlUKqhU13obivYDBHmTUFUdBKtGhZ5Gh2xKDoCNCtyjmCZYcOR52c1WUNLTS9tqnhLf
rs848FcbmvAtWyJwVLEkgaMMCJH5j8ahF3Ll29SEbmxSXMHQ5FWNYmnWgyHwy0i/BEEwRz8SaSeY
GMiKFZispxZhpUSOwvi9jURVjbSrCev6MPC1lEJuGtdYPNUVPtVjAaHvJXc3sPrE83OFWyyTBL1t
ERONJY3ZipN0LkuQ+H8lYUTG7D4JuEQTcCDR76kMTj/azvhXqIsM+GVsPW5VGzdL81IpHMBkqPZe
v4Uq9JsY4O4aWG0RNIkp5yaGr4O2IEF2luC8x70FOZhCmz4xKu/7+GoD7laEUraaickyxoVdnfK5
adfCiqGC2ldgSzMqVrUU5DEqwHytCrKPsLbxWV8cwwMUK1czjC74OE1KswiOLLZZG4wsDsAICdza
rPocyUuVbg3Zznft9OOCqiMx4TwuevjwT9CDlPkrzWnNgHo9cYxvIYriw/engZHoV4Rz1ZK6Ce59
pMb2p7RYhFCU8Km74xdOYMPDmQ+oiL8wd0mYqqLKnXiXQD2SmK/o6Ed2oRqWo5dZTBRdFmBlpQux
yFuYF9nLmTT8BlgHAVr071V4a3hRyP2gWrHwMG8POBJ7CpXyu8jkfCH7kbwYYh8l95h1vwIRrdaC
UODfQT0nXasrUwWKIRc21fJrrAl3hn+XpdJFwYT2Jvy/7ahIJZ8NsrbM6KBypQ/EYQWteoXTe9zw
e9S0u+0dH0W/22CWeju+PvuEfsTmL/z8l63ypOzoqzRvZEWZ3vk/9wy4e5MDgxdiXp/g9POmpOxZ
8B5Et3xPJkF2V8W3ajOc6HLxgCO7FeWAofdqmx3GIOsRnn4mEcXeGSS65BxudQ8cm8fY7txOpNkL
NYOUYuDR9YjM54UV1PiaqhBpIMsSS8B89sUYpeqgO+K9tUGbAFwX4t/G2sSfrShQldh4CT/NAtK3
PYz7Aa9TF8C+oit3TgF64goGE2W+wdn9EvjRQHm9xoJPBnDFCEj+2GBlJaTI7/dA2wuitzuGzOIB
QH1KyNw7JSLv4qimkCcxpcZC/C4KUtX5pkIHoN3PGNVa+rms48HGXGTWOw7jRgzJnx2Le62Ps0By
9M1lJWIzUADTVT9+0WoZ35jHDBIjeUXzzpkhxSgy6Od70tAs99noTbrKpTpD4IYUobbnjk1Ow62y
QTOS9D866Ol/SP3Y572411gligY0ut2QKl4RKBuwh28G08aPmfupeGZefZuSJbihSc57Nxkf7Mm1
ho0VVJmR/6AON5I7e8WCFsAmyzmGkrSnj0HKLwHGBn11WjEAm4pZviTu9yyMY5vm81RlFrK+jD11
dk0jJhEUcY6NNS+YI6cJGEJXXUSp6b+nLVCl4yNb5sE7jIq9ikh19DPTxZ440XI/4nu6vrkxnQPC
LfWsMqLh7zwD6/Ww+L1fTMsas2FWskWwvbwRJ5m8DOcfJQHdps1FpiEkXJVsp+Jg6XCgY+L6zH8I
pYXyyPjuk/tAQGiwW/Q8DqI85GsKulLEt/beHDllD5YpFCGWPmSSd4f8/keVz6Z9mHwmzhJLqdYr
lyXeuq5ay4i5X3lGr+2H+QNTkmK86wOrA9GvpywXEg6cO+j69tZ/RWeDmrPYjYOh0NUOrlCYhFDJ
AUQi1ucsHUvaDEwRJ2EEVle3FryvEE7v6P0PLfSzmd0jQu988bZfTgogDOdQmJx5BqjCtJ6Kq4Vb
xSejx8KI4jZGENOdDV24Bys11begGA982b91inkpeOFwKcnUKlZi0CKHA/MCcuJIpsLevl4JC0fo
4gbjWGtaF/V0M68949EULn1bSCdmtPO50cYO3iXGzUJApKPArj3MjMLuH4AYJtX/bFlnExlLAGAo
xKfd/hH9B562t5M72tw4K+21ncDTKkIjk8yyeOqdtmGw5FuLWd28VCL2o5LrrvtUJafervHzSLtP
Ky4ixc2iHcvFNE0lHYmXSmofwBDdiMKuMzGb5gnLSYrMeGcivKWN27vPLlMAe/MhqtspVULCW7bd
Z1kjerNHowzRWvGhXkky6yd6yBihIc8ddRIaMIUILTbn3KQBLS/V68ZOOZIdd0tHmkNZXeTjE+0t
SrS+MdXvVE+zhM6D7yOmUnLBzXWPi90ys76CJY3BebGRDXuz20tVU3Wtz7NRPGqYlzlu/EHY/uLI
8Z5TizOJnSaxabhKcoVXmGw8LfOfHwPnbVINhGQo5SLChPcbKCfZs15hZG9t+ZVjsUIxtZYhfe4m
SfU3IxAoa/T8LimqDZ3WOMNz4a02jF9dl5O9uwhUnPAanalqajij7mkbrzBTdtTJAOA/6hdJeobx
8EMKiRuHUpMkWavxJyPvT5kQsS8byO4L+n+uehM2PDMaXHJ7UIutnHbFIZTg5ADTQZzILde9JcjV
zovUtMcWOnmI8v6mBYwuBRQc/mcAVutgAZ+Eknnhs7ys0CdikohQTEQBMqylGBxMQvrOtKlphLPM
xoL6IraML/z6fU1rJJO76KxUZvfHAYUzgiCtWfyctu/6pFe9M9whUWDYNyTX9ctvg2CuhW5qlPF6
IevOzfCkHNEPRn8PoXTiA37pgVJyzldqij9nNB4VwZQsZBt154dKlbyKklRPfNG3fX6pFSZHS6jS
S1lsAJUw2+JuiGnn2DC4vAHG4EvuXsSb8tC0b2hxy10yx7HJgC01VRMVzkIG1XFWgL28L/tPE8yU
JyWDxWUrM9J4jH/SY2HKdiD4Ej+EMncwqoJII5ZM5O+YLaBRHcGQqm7ZlgNC1xmKOyd4qDGhd2vN
CSGqmZXzTYS3etJ0xE+QPuO4eY9MCn0jRbou0cJTiLt4hg06GUpgyCH+raZUQsRX8q1131RP2P65
eAdHLXqXlFuFsGwCrrR1UfP/0bkp/FUyocpLc5rz9N74zo1rbR6dAN6SoW8pdlgHDrFKE/RT7z85
pOgM0xg3CMljl/X9M/wN/japd89MLy1/SBMeoa83qnMSH+aODVxtLd56odct2s7UT62w7LQuvyJb
Xe38+4+zfO9Xfd6C2jxPbgAcH78F7gVWLhpbxm5eRgcFQrSzJ3ZOs9iVUoRWg4TxkWK4ubBdK99F
0EtLT0QqA7v0AjXny+fxjzLdXo7Sb3UB9fqR31JsFO78TqulGM1n0Nafth6n8H2W1W5MZkAMUahP
K5GYRxx70cNw7hD0RyOd52hyEpTtt4Dn1P9gRcPuXEIC5CTzEIQ91KwYN6T+yjlsV/4ycvL62o2V
AW/MZH77fOD9QoQ+UbZKKTkwckRAtpz+U58ioKTHKxKcieMEE4zZww8q9sjwbZw5c6JJtM5Sy8GQ
VeVp8psxGCK2UjlU4G220QWXxa26XmA6sxr1f0SxzIrZxtxyXDHTKpJ+oqe1JRQ+ukGme1wmWFnC
7BcoUPrlHjfpAbs86XumMb7huXTAUwMg3Ffv2a9xyjLNzcSA4uxoUzNbZrXT5RYZ/F7XKB7ygEmX
7FbTwoSz2+JLUatXHlzhPN8DFv7nyySrbb9gFAomjle7LTF5ziq1Ov8Au2AySYaUJ7EMHdBOb97m
SpIMrxaYPc+Ad8hLyUrwYjmT/68UN+ou/LO2q1wwrrIFPM7yoAycJ/OXBCGyNCizlrQgcVhGKe8T
wlxJmEQ/Cy2fcYN8XMXDkyJi1A43/DFVjptON366UBh/q1fC52ZbpJZnAj0Dj0q/Au0M87TP/qjk
k9OL6IwM30QEUm8RIWnvzdfsMX3c8h3kdumNnCFU9kLm2+Xh7IiCjbgz4he0C4QV9tiHnm8QjXOO
yl/NiYbP6TaVo3uzoHYSXKVYrs0gKr+3zvpZtYK3tRiTHYM5DgwzEN9HL0MVCq7DFIPJpMcmf4Ju
HIoHcnwIF3mFQ22Fx0u3m15ZCPhxHuidavI3znZhNRTKEr90G+ifsvhvuv2LRqNRTBOFgEWSprtd
BbnajPuInAaCGTm8buYD7igGv55PZ2hO4/ijl2jV4dQ7vzv8OSGbSQR2G2ATHfGZ0smP8v5ZBnwD
2jDTIcYO5LrfFSYLSXsGTnwfelX9+u5cUeohGLJyZ92lNz9hCPTbYMq77XUoe4Uo3XsMkG0rq1I+
ZZP4JssIpTFm/q4PoFR+UkU2En1Y51PbHMFA9R0WNKw8xGdbrEFraK45++yNXsKeP0reVEH42/tR
zmyCp9TwJSpSEKTWIoQ+mnSrh1SZf8V9nWLv1e7kk97z8N+uVYQUexgwtp/Q9XEvc+9e/xp0slSN
88laGPtCixRbecZxTl8e+dpJa8u/LPkVRWPYmMPsuxbvr2KiPscpgKMw9O8PBQrvX23+dbOYGPxn
YK+sG/sA6I8o3ozEga5da8EYJ7IlkGNreJbhull68u5ocOWRRkb5BbcgGws60Xc8jDsk/RmEZ51I
S1UI7tXXTF6HTL7omeQcD81Gw8Z8qwMF9/IhPsA4LNvogq+UnlwZXaGspqy6jsrjIA39dSJOd6G9
t9M+OCwfT94B89LGuATGxi0tp/iJs0C+i56sYAyh1vY0VgP9Bjwpn6+HpcaONK/a1Mwvn+IFK3nu
82uEl/k+GTkjZ4DfKaTyST/gzWBAJezibHQScOIjfviyqA83tbKTa1VnspbQkLqRHNh3awyyrz0f
wuZJ9ZQh6V0s7D6m4Ao6o5WeXqDEaUg/V/HKeTthzL5ywB5DQhSD8evzuPb7QRe8UfDMaYN/GHJi
kyBTkQKswFhCeVtMVdItsrF6WmAod7b6HQhvpUuefEIjsnFAeJ781mNgkp5Tqodk9KoqGdB1hgdz
e73VE93hESyRcadqHuy8C0pebYQ9ds7/SOwLOwMlb8jG6lODkV5s37pt4EOGit+A/rABZ9FWprtp
FstKbw49Q9p3TOVHWhe5S27AFYrgxJ1Y30n1/NIGOhah1QpdYNT2xEb+gD4k4jasXilt58nEYbTH
Ls+Qfw1csmSJltiER937hFWVw1rI9PyUeeMWc2eRP08ekIKvw4vWNoIVObAe1tXr6buJ7mgURHw6
UgGK+68XCIB0HYOMroFo9lqjpt/KAh0g74lzqIz9SYxtCLbgMTUt2nakNuqqWSk4PJrKnBjvWcA0
5P9Wc2aMtpdWXjK1ArU/ueeJtHdGFSvnRDdEmY8X2JnlIXhENngehQnegADSnKAABPttTllGdXUZ
eDZoxbln0cyB03eFHM9/ujcPuj43Xb2ZH03VKz3eQpNTOz/FJiNegzspaWakY9G138mVhG4hL1P+
ZSgZpJp7Crk2PtLxMvi/+5n6maN062pXAZm/LOBv3GO+YR/IMJFMNYdKGxTrdmmUyoZS7a8Qlc0f
bU9LV2nBC8QYO3JgpYMFlDbr7Y9L2gt/JQj7isIwqt2LIqsk07YzjrxpchyEB3ENcBhU7G5OZD0P
GTxdz1Rx3huvjAqzr3W2nt917yBUwFBH34bHZ9gEyU3tYbSX94batq27dsCNQ6mn7sDhfwRVbxOM
QO/Rkk4RlvjRWMvHAXlVdmvKKIO/qZvrD0Rtk0et9MSoa2elAvYL6t70jB1C38VP0zjobtyGyS6T
91BKHu3pnJFz7rSaR1AiumEJNQZIn4hVtUkqUn15bYNEO1SbKhRxQDKwWEsApTgpBd2k/bDPTyxY
W26p/PG9PozUhp09MzfYLjC3x0STPcHP6najomWuWsfGh1/vOlyk/LAp9qnneuN9EGWB2DY4v497
O7bOml+TuRM+bYCWaEcmlE24LYZC7tYGBNpK8pJOs/Or9ZRKm2xaKtThr5Ro0OR+YrxXPa5Znp7G
UfRP08ggr7gMtzaJSODJxkdKKp6LpXnB5d55DSdU03FO0jQNkSSXx0SydfU96ikctlnpir47dKQc
NQ+2kCeCXYA0zBFMroA2/pEOdbRWb7r8Zyqk8MFXJv1Out3ZGyh7vrn/1rzjTVXdkKhxZYetN62y
FyRD1yZV9tvKtZ4qhRCf1gTMBC43k71imhf/U6dq2gxFP5wmep5HutjhzVpT7MHUuUfei6byNDFQ
kbZ2+8YlsoLAJQlmtsguG1yRpalh309LWk4b3mUz2k+YmWtjWK0zxgwAJweyKcZ195vkhOQAr0wn
fE6PQB904dD+JjeAEVjBaHqvQDNZ1mcqg8hVY/d4rXpnbbarMR+zcJnPoYCP+EuCl862mLLGFHbC
73EcVGeyIDvi9bPeRzOHl72+Vn8dUOKOF9zqD2UGCq7uhjZ+OLxsi4vU4Sdac299P3J5OiVeVwt2
ScoEgfFg3T/N51YDo2nSirG8eiBGcBE+aDRqz7Q1DxJ8lEXUA77Nh0a4CqZWZTIoGAOX2EvlIdAI
nZTdcWOSm5d5DzYlOqRuoHhfB9wl/mGq0a6I5PmCHVoqnr7NaD013YZgIHxGVTwETj0LUByQqOAz
98Sr+J8XZLLRxoY3Z0MFSzrKKDpfc3Hknhc6IP4DWK4xHIyM0mmT4fHNMigaavYQR1YaLE3J0UDx
f6CAGRiJcFwHm7hJU4jn5FLRoicwat+MITv21vTDanH3YRfmqYsjeiInMdmUqW1D2ecG3gAGLCHx
MDLuM8rUH8FI3/03zS7dCvJlU8qEff7YAzc77DoVFRyOrFwW5fWOfP9zt9mCpjqEtaIrY2y3Cyrl
9Fe2UDr4t1RlTBZmxX94C/lwZyH5vQUhBvlzv2QEFdpRwFVfwlGxM8yIAtfCSHkN/8tXRep0sbY0
+EwQmMDlRk1xqf9bhO29NesFMUPrAuih6YzfhVoJqVtqSQs7GzgPQqgfbMCdMoDZtx+E9TgUDz9N
iytJZoKTsxs/Qf57Y5tfjO0wTpkdpXe/c/A6c3e+shR4cVtc37fe7ZxK1S1O5R0ew7tUv2n8NkbO
XYjSIJPq9Sj3suBULipsNeuQAMwsfVgj+160VZiE4rRqTYIiloyy/IwyaTWAFJKD6zI8DLclVtfX
4y6uuMj2sL3U+FLI9rB65AfiC5Hfe3QQw1RrsShUfncHqVZydoV1gUtuJR2k0KN6ER9Sainq2vJQ
qrfObEHeg2Di5zXs3i3nMPxTrqUFLbA2ftIDbO0QGoplABHw/8g0f4Xi/p4qfXkoxPrvgOxiHm/P
DRsSWKiqxydYPenBGruqikbWImh60DtBxt38SqHbDRKH+vcMeddZrO7RCIGyEs2pe/QMox08Lqak
oClzkT3lslDfPTniLHxKsRAeLrqJAikL8sY++a2nrHo/SBYeNLZ4b7SrJ8qod/TrElT0LqtYSFKn
3Xuhm3VrqFZSGP8K3YTVmT7d07uUn9h+iJbXw2ZNFaXUZ0GY4D7wWjSOsxdZ21coZ/AmNngLuTzE
1sN8cEnHKgNDspXxEAn6AiJh8EyhFw5RMLnZTHwBBmNypJkTJAZLXW6PA7rP9NIxWVKlwkcElCTy
sL4gXi0Nhs+omiOYl6j/aiaf+zCTQFPDAhUJxcpp30WRSZxFjDZVnUKZgEp7f4b8MaYCd3ipWi9x
Pyk2G4Rjpa3q4Tdz4K9Y+RJBFseKH1UlBR2vW0zQveCQP7VCe0N5hARSWkPf7lMFPubJWGu6dUhM
x2qVc5Fo8GCBh5Yp+467ZJd9E5unbyTdL2aEhLurmeX47XNz4qF77IbiAgBUFqCcFMFq2hD/TIan
Ht8GcDbbvYcsHK01bl+JynPHaiO9+j/LB/VPDOMvsvUbvSZ3azYnRmoctAIrxEt1kQfwRg08CHxz
a2nrbVfxW/3uIUn+SZa4n43uNxMlVLID6rYB2p09EkBJ3LuWQkdpmslGEWw/Y24I58ES87Y2D8m8
PwIBZqajQIIWV+LBEU7dBVjCBsQRKBHxwZxt7DQvhxUNRbCSdkg937ykZRrNFtr+YplEO2zix0kd
WDxPWbKiFh00Uo/aWyMn8sxnSkNw5+pkNsq8aPQ55RrpCNMfovZq4yzNnZ93Blo5qK5Qy8UzlpmZ
7VszMUIeeNiU4h3nh72rCcA8xdm82t0H3idIFH8RU1WE1qDhnrqXkmiDLPdqdUemB/v2boCZpU8X
IkqdWIfUT6FKierfEh6YBc5BUATFGYMmjdm5XdnvQUcxZnUvWVlBjF43COKgcecOr+AoueHNBO/N
jL6Ee1T66O24RX0TVDZax7DL7FnkaKhs5oizbocch5mv9vQvVxveIj52bZ8wYhbbp1W40EGPqwUn
dBhNTM/Pjyc6PBZPzR8rKMtqLEvFq8tuBdv98EvJzIUwP+7oCQJFCDKDO29tv3k68TAVV8KU0v7H
ejq3rybXtMbwr2mBYmXZRoCHW0X82XmYqVxpCnoSpvXoUK8/L9peTYbdm2lsStLM6VGc/GTRfvN3
xN4WudEslqvyGvtHXSioPH6H9evdKCOcNoHJY80wbhjxS5KSIfBxnjPMZTndaT9Ch3jbLC3sNBeA
QIWvZn1J81xXN5qmYdhV4Y3Tvyjd6TmTUUgZZAwxBbrVkKKEAwMKb3wBjzABraNL46+zs0LnkOBw
uZ0nFReEv85/a7Ms1vTbqd2NI0vXSE0sAIaYV0mFWo6e/mCoaLfkWicxRrGnjt/bIhoaAsVQzR2D
9euKSCMH9736t/6o7SLRzNY+siwP9lbzd3zhbsQkVjAvzY2Ubk0NhtwGBM2q2y71p82UtjCmps2G
XkoQ9GwIBbiCjqhvz7f16tK+Yv0081IwjZufWYHtI5mxgItEiQxjQnhHlgpmvni9zu7TYtiXvQo3
ButGTw5Z24kPDUV6o9N7sITfxAX/MiTrqi2f/MrQK/oxs6btdhRfUfODv1ZwoYaRiMlwWB9WWmD7
r+7r4tEzOrgH9YuDIgLIDDQUuz36ytETc1I1P+YZzfnNp8U+9/vFa7fusSt8/I4opcuhvrwKIhT0
GB7NeWsPwANYYrT2VJfiifFPpGJs5HV5uvaFT8TwQ+ttXBQgzK1D+AbRzvB7IJTG1jOlnzwt1/hS
PML8mHwubK4iWb1QQPumv0o82nEd+t4WdijA/RmrcfTzTKUaC9T8B5YnPENpVvb/ZqywmFdxrGPm
+1XPpWDhdl3S69qgqibl2Cp71UItd3EoycrdcMwQyCJ9XO4H/b7leSw602TawVoBTaRQ2uLRKbUG
nk9WMG3EgII0qmTs0bzMcg8wsue3RDerSGsw8x7WtLMU19dzfK5WP5jyr2SLyTemiM76FnUH9OHn
q2MzzRfn210oqDmtdN8oCeNz7wrGZGDq72lB79vTNt5pL3RxahNG/T08BdkTuqTm+dKl8abBaIHB
rwwbOTkGUbsfnZcK5v8uZWNXLqmXOx+xnEe6cNau6rGnpQE6h9mow8shOf6W4NVrCcbxhrIwzOt2
BIVfgpTwpdh0cgJxH0v51Ca1PvYHizoaxM5IE7Ofvk0S626BlgFvLjrl4TAHQrUX0vs1MEbBVCFb
0ymzfhjgyNEb8nybEAigvy4h1U9A+atCK+0HD4TV6EP3iAS/7nD2tHB1TTVuTRLpq2PwYbzL43lB
slP55NDmAdguuttWrMPGH/ziZgtlbu3IVv4ks/ZRnaSsqGaF46juB8LNy9HrjwsOnV4VY0dWW2Tg
cnh7ZDIiSHyQpCn53YTPW179dKNS6Gy6+mB995Vc2UxGA+TLqEejPl9PmeXzjFEG/kQ+H+p7bUcO
m0636vebyV7od9L/6zgBOHR7GZ60WcjWAkCSYJeofaIm0hBriGROal6oEaA5uFyg1r50KCytdL5O
tmILrkT2neTixCDQp/AUZ8EPvPgumZphO7rEJiPQAUd1sdgNsyebyn9/ZHCVMZOxPRPwzGh/6l47
2ATmhPeUTB1aD07iNcDma0SJXDI0ndBtuSABG4igEw19i1e22DrMosrReCjbeCEfF5aTpFCFAlPb
/gWG1mIDpPQ73nYze7HZGGUY57acyIuvQSgGE1vq4rvtBftLaVe3ZS793SYuAM95rqgxcK4WL1Jz
mx/2fQzSQI+2StwcOL5SE64641/kN39pEGEJ3dgWTmZAS81PLI7FJnjjOjpPmBRcDillDwI8RrVE
C3v1OUmRPld0zaXgLzP/KEOLgV5Sqz6ilQTFCDmKwhiWpGuEjbWBgM7PlxiSGxaBkTSTdi9FRRwO
rbyBhQbO0IGe4j4Q1bEl+GvQJH1TDRZjbN8YQHOQ2yk1+aleDl18rmDtynOwg+ZLwEgDJhXhQ1Z+
6Mgn8J24UliB3HBpRX0Xb752bRUDhgS68q74UHP2rXF9NlzBOeQAL6IecDHnG2CRJxHx1K6N3COZ
AKR4zpbR7cNRFtpXEYSE/QhVfVXyGUGzo9GQqpVh8U3Fls+yFcpITFHJt1Kizbitil6RSxauMTkF
KDN2Y8cZGrHyaZmBrCMbgUsO8UjgSzFoB6AJS3ONufomvwrideVNyPG560Udc2LOa0Vp9dcwuv+y
01vISOBbwu9lHillDCt//sHJZRS5oA714NzJvfQTDShIk7tToURe6PhdpCK931xBCePu0gtq3GnU
8VW0kn0igpnRwxPy/+bAYqgv+gmB/SaxZ+KNzBtPpIdTeiFXkOfrsBqK4Pkg9W1l5zEVqnCb/Jsk
L1ixo+MOeokZfK/rU24502wIfszvXCcp1sjlpRCFGY0dUcrGfyL9Xqng7d6cUFkSINWeTFEhThop
QxBP9Wew2U2qV5FTG+Jill3oc45AS/+wEq7Z+GNUr/FZCkRnFNVg4TYqQ2RUaJQlapIui/BSzJAd
XERLkjbxGOlrJ9smkhFdNZG5pf7tIlJ1lfHNI+GiCEbmzE9J1kji8goQByg5KUYd78EtAqiYUgsO
oABtpLBpZYKecuczYnAKHBIh2z3HypaIPMBEzowoubP5i5NWwf5iA9oaBwMEaRWsf9x/zv5cliZC
hHk6eJStLO5TrzBHZcaA61QzHuvQt9/MzeAQGTAHOGrhoTruz8wGjDqJkAFL9POm3ruQs2q5CpuF
sn9L+Ahv79nm/foUqerykY5cYAT4lGlAXlfGhfg01QD59nS3MtZyx/d7W/WBfBPNaYq6qD7dxmrp
2std3LFjKD8W0GRcsXq0vPEhdagVKnV41uDFaIz0vCzQXywX0Jdi6XzXf6ChSPTo4tEqZsn/DPsm
x4U5IZXi3SmWFY9b56yzCWMrMXvQ9CGuB0bIWcEpxp+z3NU808B8lxAZDdnOK0Pz3PYTTRU/Blqp
IU6TCmBes/sV3LRkdo9zDTBhW03lvb0XlhPbOVq4rfMy4CaGF8h0pScl4T4jfT6byMB8ciRYG5nx
V3yNK2MBBOVHpnh1/DVAk3MN3m1A0XPSCASJwuB5ynnoCRYcAqvK6XXm6o1wp9DJfWFBUmWAkKkD
2OaVJ/NZes0y56Tpplpg7H/jRXNTLJBZ59zn5nEY00OEq5kEo+kkK4anrSWYLg3fo8X7X4c56G1x
jlt6MJuDwOjU0BhB54TxYMDR+HoFKePECsmBptPHr7JSDYswv/kXJMuL5P8T83J2kfOaq0brqxaJ
2zFb5gy4HM73jPJ1loUJx8N0ceEg+okMvM8GZj+zacAFU0WpH4OzFFc9BQpQGJIEYFv0t3oDVnGy
YRTxtqvdgofzVGjrAeThKlha66u4Wt57EB6tmXAWAx3oOn3HhqpYfXA56FyVD00UmEV5PHAP5Usv
08D8GFq5elqz5TrrCKH5gEwrbyIhKWdOtVYXqOtLsHbr6bndrRLrnSfcZh+MB1A1SmazoQxz2B//
o1RJqGJGIuxJFkev8dCv2UA+5QWK6z0ot95EKbHntxZDeuYw5ETf4KSRsxdPi0+TxBbBHL6njyrg
bmDkRmdN+9VQDDLopfAy/j9ffvn/Kwntej5d3MECW85NOo/VqFeE6AllG9tf1xfN0FPNKWj+0Iux
ICO646tLIEfMpS8br2yVE3GnURt3H30iyS/2Avc+4NKc+mmMPkCjef8wyfN6mBxytbyQKlOzbvcE
3CVjLtq0HoBT9M4gsu4QVYxqQ3PiZfGxpExrLbGV3+8MuKxVa4yyYuIprPJ0nD7AcQRPGHS62yJw
dtxO0XaOgDiy8JwQug9oyHCQwQZegvuctuI0CU4hPlIxpemvosC6X1x3Ha7jcb9pGfjlE14iff/2
f2iGkqHTPgY+T2/QYVhp3IgbIjUfW7p06WFlY/ctJoTg/8GRGQ2KXLN57eZGoG3WEAxaN73uQqDH
aelba3MziO31i3mgM6JfBsU6JwWt4ffCDfeLOdj4Hd43gaJkYrsvN4/N6xwCVuT/iv/s9jPtoCvs
CVhbtXEnjgL1dOOHFrg13MdmjXe0p8WLtTqJWqPsjntUmUadnl0maddsi9CzEz+8qAszbcREkRvT
FbIVKHLW1WsD4YdNlkjTDFth9N26ASNJZknfQbgjNkmOY2vwgpXf6mko6rhVMyGyvPFFLVbRD1qb
XnEsWxAdYNGepitpnqANtXtrIRO2e02mePbAmLRMjANZ9H2Ok40HfSMCyXjvinJpVbonN5wst4rB
YD71I9blzUjAuxXbkI2LtXKj6/tPNAUSMg62Pii/8ZLoos/s68ASAb1kgwt7Y8DTvHk7nC9+fQAO
C3Y4HZAXxNP+9T+tLrMEz67uhtX2FpomlK3Mj6DvEYoxsR23E+p8MOHRG8fnC9Kn6pTS4hsLjpEW
xuFJ35wRSwp18iR41JCF/SBJbeakqxHuWe+aDVnE02SrLtRJwuQbptLudNWnV2mgvY6XesVsDaM/
xdAiWlH3ATIdiXPAFKviiFHabUlzBA2zHXEI9gMv+BOQWsg1iT0aBi/lE5w9uOGhSqL7a4WDwOao
W7xRORtS+9HUWZqqiDKQUrqWZAUMG7AmgWaOJMcEIBxgku3EtsAmjSrGcBH7qfFyv1Z8zqc3E+FI
97cCtK/5VuWVsMnID0nBLgtduDYGVvuPMSmzHWJK40+LvyJlE2xj55Q2jrIzeONmAGjKIdPXWXfo
9ziEUIp/BHVMaQVv+UlSiAE5p6IEQZeY+tY6/LIBuj+aqy73uugYIWr6+TCUovxgZa+jgYrRMWWx
C3hlJDwqQqahvyy/FXkOceRzNJAs4kIj9vhbCUOT2N/guXDkNrEHYv9Uj+HGyz0JMe1prVKrJZx7
T2TuryY/0OlZMLXelVpvdCh52oMltAXH4h+QI5vPdS+Y1RF20r/4Z6F93wm40BHvPxlHq9j9iUzE
GNteGmmkF5QpWTq4b9HNIdMVnRkYizjRaXKtxQFl3tVrsio1PlGwfVI+l9UGjyRAXWAglab9RWrZ
OYH8/RqChiahowQPua15HI4pwaOQ58HkVweyFzpexFI0MP+7757iKdUrvR5k+k62qoR+c+UWKVPO
x++GQf4HdbAdq/jCzsZtRChQ0rca5GcSvXcz43GItDKgMjwzK2lQRlK1zq0X3s2TZGGXHcuXZw1y
IAOdO2M91lwXELDczKQq/ziDtuLMMRuZ1IDtz3wBbk51a6Ka2rL3XuTUyduXl3uXbbkmR19TGk13
umAODk+1dyqiPVHgPcrFjptEwDa0tRQziIYJuSQsRMz5PWiXAQsqfYHx9JI7n4G95aB3R354Ngr3
863mrtpAtXCnjoF1qIY6SgCWJuo3I8M7QE5sAqs+zN+3WwDygYHT6gjJN3xFCAAo8CnKptj6JwJJ
zDQRcHU+hpTOr7h7rORU7EOoSTBmk789ZBguIRps7cDFtGApvvqVkdwNpCcC963nelBNcTCgUgUA
/krwWwEWEguE0FKDtOpbK/Hbhu8NJ5vikkx22Abs05n7eoYl3Rqx1Ym1tVxtCdnsxPpDKmEVvqGF
8YCGFkwcZaq7XvTFdr4tSGrq2Vg4gRSi9h1MY3HEbGsxa/0IlngTkqRzy8rFByJocWpcDXdqeq2G
CeAyDyvP48upou3tnM+Oiap4R7EGyQHzDnF36o9YTwlcDuuUrqFXtw5D6xGVu1U60WKGqr2K+X8j
hi0Y7WgafpWgwrTIpsrEyIM7eEQH1giZVbxtHzzMoAcJl2LmhoGzoh/itiqdzcLRe/uOboJWLUtO
Ps3z3WLsF4LwfFVUypsOR0zDiXwA/R1Iu48IDeGrzkFOf2rnObnehRFpSHD3vR21EAa/yQ3w7mSC
tTkbRy8Cn7zogdvqDPxXL2sgWYI0dieEXWVUvyyfx0Iu83gI6WzMtixv5snwCxSdVgqS6Z6er5Fl
43IRSxZmNQ1lgzhW5ubRG6jWvpQ42q5gOng7blMDeYDxWIONSyFe37Slk1msY8aZoyTpTgRVSZUX
EjbgfcAHbcA67dEa+BJthenw4PSO1fGCQfTbI/zMrOo1FDd4q5/o+VE1fLBFUeUOS6iZFjSpF5cZ
gBEaAvAWraot72A66J3y15sPjwPU9k1BLUA8j3WP2vLLPOdcENR0QE899sx7UPFPloOH4Gqtpe3g
1PWL61Tgapk9HMjBt9lADcQ1n6v3e1hmxkLUVi+uI3MRi770A/jav4Q2kph9iSysd4s60HKG7ey0
800B0thk/g7FpT07vszF+bQjarp7GLGgWXTacA2AqK1j6tU/OHys1wwLkBJHuNAH3dH1eQHq6Ciq
VrkH5TIO9rpTr8EVUpYj/yKbqBSH0SuNvDmQAZJbTC4JTQSL19gR8ZEz7fjRk7yX5kdXn+N2fgWk
F20ZqmNcwd3viOoqLYFp4qKTB7E0IDSbPHmUdMNlxZN2cK6wTVsZqTKdwn8rR3VAxsgRQQ5qKEbb
tmzlch/PnPEgYm2cd/px5+4HUqaPj/p+kgjo10rlup7FP3NNZALAO8ea3GFMd7nTKv511EyA46Uu
vP1CMlh+phZsG1eadIsci4g6xhDWcBZcKZHK2loleELz9fme+R0kiKa93ogdcvQEcN2KAldAMf1i
Kvcs7NSVH0xZNGGCdpGRYQ9AhqfjvCFMG9fhSl4VqFgOjiQiDU3rsX6/675hi5wKVxSzpm9Ty0sE
HEX8idEIjH93l9EN/ZUe5iM8i93jVUvb2+MCHet+XWk2mAFqQdS07XK9JpRLV0vtStmC/oUtJieZ
H47+TzngLTx26sKgiVjBw7qWov+oCULVJ1dj3TrD8HXzRwPCR2oxLnQEMpO704tKgSkNSn9kveeI
bJlNOFLFiUnO2iKH7Hluu/Vgct7HRsrf+bok937/yJZ5vxxf7Z+CIdSkTyPiP1A6cRHyrLf086+m
dVyljqGwawSXPuApfJHq5lhF18S9LIJX5vgbgtePxQMec96XkgT8v2q+DRJBrrdUlLjKq8MFm4RK
Bighr3jm5kHlcEyy76qXDkwPiSMZ3CscWW9h0BDA8+/BOIswWqpZT1SS5wBMt6VUTp58vAZZoJz8
RAOYWqAh+xwoLJHHEHWJNpzDCDeajbeM8il07zcJFWhikc+lcR583qfgbK3tRpq9i9zENMXch2CO
YYFPbqeKvzhuTgOtSTfZXyp4Q8XWCt7lL8aRIV7cPcd8CNVZIiqAbs4UunVfFybi022hctEQZ4BN
7ETqG2FltqYsYvNnjV8d0fHJnhkF6cLlJeHPzQPDL+afKsQkhSr2SqkO3Ov4itK+rgg/kcz1KRad
NJA9kSrIYAO/exo/gVylB1VSHd1WV5g9tYzDu3B3ZhhXjzIeIhVXwtzNejuBNp1UFe78jRLOl6a/
f8rtXek1xS3od0kjT6e/+VKKhya0/WziMQyN92j+r/hULU/3eAYtyDfgdQOMKLsq91AvMH8CjOpG
fKCSYn8KX/YlOZVk2I9W97hOKNIcjmSFCJm/Rg8HpBQB02jgSyqMa2yfr5dqu9p6zHoqFmF5Wifx
fqaF6HOJJDcoTeLy4j/1NnxV91939AzayuiEMf4wXbInsgdlZqwB9+VTOzlAd5Xq/7ryzxmhanQn
vJXzCyX5/J+jLA0KvQtlt09nscZHHlrsTvEN2KkjN+GrxnJbHpn1eZkKIosF3QTjNEwmg1d4rJaq
hQ23QjguyPny2CXHGDjaGwmQg9e4XL86am+dGLE5YMnB/iak8Ez1I3SLkiBK6XAOWcaexZUb0VL4
E2R0sVMmY95z9XEflQshTfV6IZh2DG10lqfKj0lYpObu0NozrkzLYkzTSoNzVRaNrRtxH+grRm0v
iX3frtubu7jKSkkrfD5D9W7qdTVWkk85I5pV05LPhBIkEVtoLWoURQnp8reFdWP6/aKhAVhTcoXC
AyUV3EoZyvuFtB1kZeIQzxxx8E06yh2u5euhWi5j79KfCxbIM2oE2ZmCJDJKSKTvVWb92BHqVaIC
mLt5tFIrq9WFtnErfqP6IaMuPkh7HPmR2pIQlpg++lT9Cbq5y8c2zd8WRKzv/3o48sjZ3Y/I42ub
SzR/j+OtGa1C4eMVZss33hGvsW/30ON/Za9M3WokqvxI72PUnM+Wfr4/YqQIRAVhYD6VEDm177FZ
I4E5/pZ65ZhSufHejw4GgOsm3YZEBaNwFfjQfYURIwZrn0RpcrfSqh+rYT+/JhIcF9yERh1SSAEk
48ZN1v/hIuHk6raJVAPf4KUCfpNtLBCGEYWI4G1Etu+t12lLLPGdvadUX+yPnQMPtJnIv+vJZoQq
zZ4j0kZdi1DXTilW4mWZU2hgEwlNc2hM+A56Q2FIAxmvTT+K2moEGWoTp2ZdZkAVtwCXhqzjXO+f
GQWQN1a82F5bYiNiuaDNsKN0dw5w2mOsXcIjWiIo/vo9GK/rSDBlnsmDx4T1rCruSyB6d55KKi9K
JrEh9GWr65J7BISwNWMyoM3lVisk6Nag25H6250jWgzSK7Qyvxxe1zWvV4HGLfMeAqBSQ0INK206
1tLtuzDYR0c6U8HXMdn9Kfsdk/V278QI2sKFTTugPoPn/TypUzCs7ZvyPKssFycKAF95Ipd5Hs3f
ZF1E7RJvEy0vAUv5ZSEJNHZ0AoIC+qCmydEpEN1BTB3G/XtfJ1/+XS6kFbBz7DQ+g6zxmKbPUA2s
/LsshN03whQtbRrPMgnaIeHYYDPzOwSAMdG8QWTgHNqdIye120CjaIZF4vSlEallFutux5l08u4r
/XImTBM4y90FV9oGjRQyFcwEeCHq5oiYpt6Czu9h0/0zCbAD/Dxq6XL7BGCKB8jaBTS0x14uWKbM
aBIpj3NZk9ag9JyX2CQCOVjpRomGVAp75ygfCvfQf3DdukXAnip9cZ5PclCFHPE4uDus/2SUqGNz
vWCtQXsaEIYiVomTJoYA3YEJIUiKAomdV6+qL8AlsCFF37Qix1E6KJx0g6mUVVkFuqFmsyN1+SPH
5vThMOivgXwse0A5mZdc7D1LfqtzLMNIPm91CQkqgUt0MbrEu3VYHfNWyetAkeqW4QjM16iPPu4z
h15BVSGw7X0Ww+oDxXbf5v6RdzeF+jC88TLWbxb8okjJdtNlhqoKTITfJyKsYuVE2k5PuyDS8fSN
CmmAQCRLSEtd5m998Y2PLosX2+mZRTM/fGbKkJ374D0PaClmlnuyR/jCIHZqjvMPrU6fP20GEkM8
7hA/cs3fAdRgjo1CIAl6iHYgOE3V66zG9kLycyEImj3/sQlV7sBLMIA1hfDhWwVqaxtyhElBQ/pg
6XwSCbE+ML4GVJNZNB6L2/E7rNdEOXaJok4gQHczm/h1MKUr1O9uKSxNK15J8NvB/0LFoStvVhGa
XBvSlqTZ2qbqJbGoL6v+9waJYVAtHGlmqMCbvxtdUxzcTQOnV4ZslRo2nBxK0/KFjy6x3fhbkIgk
wtaOHKOhAhgxNsuP8fealoEtrn3BJH68iVeuwdXfUTrXH+DYmjhYzZqoTrFV/72+8cQ7sPdBlpgx
9Mq46Lib0HPk89J2JBaI1a7oE5g/7Rv2mAAiRBHTab7nVVrUMjvVZtHqOR5JaD0NI7hSw6fKs2C7
UjJjO5oqfaXuVeApWVEXDjXqpMRYox69CP3MhSaM4yJtdGr2VOjl/kd8yGeIWdyYf1FOKKp2Kr88
JFj5r5zX/siQub6pMjp5xKmhP4WalEFGsctN3VOvID2AgudmDRErXWBIUX5kxcg/MFPrIvZNCpRh
rt11LuzUPZIhsP7JABLTaXtbTAl/0elRYJnQftZ7kmV5SkcnfwUo5ikFukL5O08YE4oCJaDd1Onm
IROd052UA+X1AxJdPj42ferf8L9tNssGPcYpyudEJYHCjTfGQPwKavflvih3Na63l4wjxxZ7lCmr
MfmFSXcqlkSRy1jIVKrWPQpFzY2P2HTvXjceh0cvX8XmWSUrq2FRy6LKls1CnUf+Gml0PGMUF2wy
W9Fnk49779DrMtytHAOWImS4MQayYbMjrnrV+XLFz2beFyHphxZ7AjK6+7pw325hzA2goFsLmB4h
Kd2Daq4nyc9mvRwJDVom6eR0BIDPXfC2EL1pStdVgSeS1FvH9vEfX/rbYNaE6N4pXhfaQc3BDdw6
MBjEPX+EMlLbGWtOzG+kcRwQ1oQfiQ7D0/wDooeNCxLRtIbMT3uWtlQv3kaB8hmKAaZS0zoCouEL
VJ+dA6JXI4Z7fThOXQw/g0gYmz9rEj+G6fggz1EPlGklkWi3v+qSHI4HRNC7okeKq3yqtxL6ffpz
WW8+xaEEWKckuzQOye7wPZMLXUjKy/9JqHLc6cFqYKmLVrhzBU/HNfVm7UKBnG1T/YH33uVC097o
RZnmdubZop+XVd8xPXmJNscRtdXznpoSb2xOdZtdiC+SzlLsz6wJUO3yfiNBnRiVGnrxVNkLJmGz
APadbkN4DAtKk5LYhQXFaGno+hGU18a7DqYv7H7YReecb8RDCRzXT/SSTG+lyEvbHno5lgjmE8hX
eFLOSkmNVBVq4ll8aXJU9iPro4h1FrDp2TET/+NT2PeBv9+ujpfgHa6OSTO6YQjTkc1MGOTiYsMG
TM9HbVIoqHlc2/XUtTYodyj45ondHlyYxgiQvKIrBDtzte1mBqlSD39/gaGnCvQGAk3YNzOy/rtC
e/m9yFU9WQgPhF5DoXU1wxE8haTGKRhLkrY7CI8wOHPivOdiGTEIJn85uS3rZ0it50EqxKYzYN+5
4KMEqz5j8txhL//lDmLJAOaA8/bxoj4z0x7CIBXPdlRh1kGsbsLanCUtrBuv1rO2VdXIHJW92WH2
OQXHxgEuRpajCM1XFTv8WrknjmjgJmfdrWqz155Pe9RRZYVqLR9J3ziR+XYMfWbBg2TJQJEtGWFN
7OX+axRxiYlRg5AUE/tXE3Rz6KZQFO5ORXN9+WbQL6gUedNb+5/jDX+sxvubkncLZZ5ByGcZBh0o
EOqtwMH2Dp5znzFZT6ziaIzxVtQbs9OyaO3sIGwPCtrTa8pKgQWTH9fcQ10J2woHErhvom1N1f3j
VCsSdiwkEM43vcNxRx9qznA13/Lfe7hlmbNF7k2B2crbngHKYOlmVxoDBkI9NHsTJenQcFqlRzx0
Xk9+TJScWtmrSt1FzN8G/nSO4RSRRN0BwPvC1FMTZCLcnrCjJnqB0/zJotTKLXMwy1WbkpefProc
G4kvzr0RUsQXvlCQ1LA0lzU7/uGMNQBHzTvuXGr6XAyDboiXQyPlFt53HtJwK/bc7hyLPvw9IMCK
Z2olOXKvGbYZgTxqSyArVlVmrOu4v1hW1fFX7S7/FjhHk5gfsOzxKahWIgd68s/rtKx9Umwz5zig
uRAh6enN/w20m6fmV9o3SGMc1RFGKAUdMqxNGcCpPRgZf+NYrogO3jrnMetxzqenL/7QvOcwWmw8
ylCc8TMbD/GHpQnS1TlXg52v0qfsuZCHo0obXRIR8IyQhtdzMpV39J7+ouCNFUrpG51ucpza6aTI
eE2IIDEw9vs+ixas8kyd9WMTpeAWaa3saX435CRkPIrGABmrdra7XrWnYjbXN881XInZ72RX0/D/
Hc2MYiSwArQyVFMEKJq+3F1ll0jeuL4vDD5BpZR62faFJeXzhvCFQ1+u3thpcoJpcKwShLeyJ6/D
TEvYbaLBZd4ipZDeHh83uUAtIW8bbGgNUX0Rt1amvDcgxJz8d3vACChCEkVaLwT1v+ArPUD84TaA
dQTGxu2V0CB69M9Y6cu2ayXpDNfzeakKjV2PinmPiONCMesEwH2jJCH6hzvSO+L2+Zsw8vb11Rwb
yuTvmeDFJvZrFTarGmjq+s2wOxodX+7AxELiO7Qs26BaQ8m0a2WEDrpKr3BThxY33iROiG6elRJZ
0fyX2lPVA/nj3SGGrTxg8IXF0gF2MuedUyPzFMel9DNwh/ksx21AVi/4+jExh24HZHiR6Iyx0yBq
Wz61BvpEmssTblAXqrD4zGytOdniua+MMaiEPY8Hnz6ASjbYI+9YzLlAXJ9T8c1cwZF7cgsem5KS
1HZwsX63S/VyRmol0zAKDQZ9E880ijQy8fbQ5EYkzUvmxAkto6ULQzUUSfTpvc89vcejw0R42tKG
Y0fQeutIDIw8kyf4FIhnO0V6K/SJyTFz/skokpNppfLgFHSIXWenA8YyGqpI8Ovj9POk/8nFUir/
T40HLJHYEXPdM8bvmLmNyclFS2+gyHGpbPi62q0SfWXPToB9c9h2VGSiAi8sNQVF6/wEZs3Wwqc8
7s05TSOUC35wqqhTRlvstWSIhXJgNbv7WU3w1WAYOdd2sdkRrBs+EhyAxWOEqDFbGO/hv6q/eHrT
pjdzySwH7F4lLZS1Mb/NHRKHKB/mzbOL9yFbxnq/bZiQUKA+gEC/0eUQ3zYkW4M6389PGWwLMkTH
J9Mxj9pkggQ0xUc1pQiVgVMOvvyT8k2wT1OXts8w1VCgyoJ3FOtB6Err1YUXCD4xaBccUcGNSy/i
QSapSTlN2EqZU24VPcjFBL+6mMy/+HxEkE+xXgMUWP2/bO7PkAc73I8nzEi5hz8tCmuvdYTIT3v4
AR6kH9x/1dKV+uBedIDqy4ZvPw+GbcvkiC2zFHiuoj5yTkGAGFoyrgZBJT1acr+9bFp7l5Z6E8Du
iqBBYvwoabXuz1rL7di3ZdvnOFYnVj+iHRp2zskRA53xXR+A2cVLa4ot/hnsAsalcedFHIfep7lV
MtZOcTJDLtBb+uoWvS9qVK4lR7FNHgsyGA+6+XfmKOxLM63187lSTcYW+1STMm6qGP81GEa1EICo
RX3DaJdxcSupqM/r/EBole1o9CZnU3OpDYZ4O3Xa7xbIVbvzlT6hcbEece+3IyMhlCopvWt7PsjP
wNuOC7QUSynK+DhNf6ILlwahNuI4f8ZdWAGFlx2mZQLRgvwRJGlXgynhHuniP1ltxQS49EQx6N9N
UTvEZeVnt5H/XGuFxBJ036j/EC6JY4iD7h8coBoxAuDFhDvblXDfczgjjkgdHiCFuXxY4cSXVh+l
bFXTgARd0MWJ53CKePjoVDJgk6LWMiz0kAN5dXtAgB+XEtv3Q+2vo+z8ZicaRlMvAn7diBlPD7Ce
bXamhZyMw/jGgRGuox14DF9nYQEawMTeqK20FAIdg1p1w6Img7DGneLbOc0w8kIIJagSlcMKBmjI
Iu4pTif+UcESJd+ZMZbAu+ZGBdoW2HBX/8KvhA9M4ACAJK1JVJfVKrRopfDTFbE95LEk9RZGY8Tg
lTYY15u+JxLtw8GzJpveibnxl2BZVSDfrVl8o7g3CJhQZ3H3yUOz7mK92xyUNhyBhAFcGf3gO11W
pAmZhIpZIDR37Zpkv30ZWKSu/Lm9Km0UXlMH6pp0PMSrcUZh0g4EFzGCATaDf5japuzDEPefshie
YtBomYqvy47XRqVlQ7xs6QFkZ+Wl354ISsIa5hfFFBhpq0FaFDqEnL4nKWPQqSUy0uBWwjzz7BLC
H8lyK3gFMAw9zLvT2+xY/FJow7f3KnVAVoJ6GqpryQh0rijuEuTBKsRPwN1cJqcClwOhLG7WaPD0
vqYMYBa/RL9/m9/6zPrcVZ4FdJjygpFlQVvkA/Roi1hAXyMAK1PTsFLjDV1TOIxAj2TfB6RarrLZ
Hln4TzTMJRm42ec/9MokzIoNqwIwLSzb9xXkxwY5Wej+AnCrsYexEM1yEdMr7EqcR+ITCdoXNW6f
lfU/SLSBFrm9CJkGy0d/CwsXa5qeKuhQPD+tj92OOPzS5MLnPmMw2ObDKjYrpWt+zF7e/JkoRNi1
AgOe6Xr+6GVXUrfHJTFRBVSQdfrahy3SGGZOvtiwnbJos8LyMqdKvHJDRi+K6jdAntHCPrhKMzXc
I2HoxCTCG9/p1wTTUufy4SzRXNEfoPaZXm7kTQVHBQcjm0RNTy6MaKQOUD3wZxN/f0hAsAhYqaPi
k2fvYxl6jbsE5Eoe2mbBnBdE4mPDTqqCyPrdYAwXny2mLji8Phx7elWON5xfJUCbwBgZAgKunJ96
/qV2blq/ufzg949mDf+W61+pOptWz9TrxKAP7bT9y2czgxdHwi1RRUUROZ7Rem1k2dYizsHeiVw+
aVG6fZPzBfqTHQHsXhpW1iiHKQk1L1lObe2UJp2ZfAYSkem/Qsdcjb3aOE7iYiyK8bJc+v8jSEu0
0Wj8A703vj9izoB/WpVtvGZLA2ZKtM/TSS8TiuM4bfNs9UH9BJ6D4ZBDYvMKcKhkoZ95+b3SawUF
TO/c9KueyNo+2PQUs64t1ib3ZzGkgwO3/JK1GCKocNa9iqqnnymKYi/ASbRnxOUIFcq7ZzBN5yW7
v+y0l4swNxqBeSCWa/bxAFoLBTSqF6QytITC4g2Nm1MvuxGMOiOzICt7SjQrvuUfw9JAb0E7FVlc
M84CK5z5D5ZmYKMjrwAjbZqCIfcxqtF+Mtpj/JPH7AOxtPvMjJakuTRehzErJde1Z8f6S1cT/XHj
/wFIezrLa1hjZoW22lKu32y3TrJpgP53O/ElBS+50AbPTmkR3KvlmUw9eXmLEGJexxi5Ln2U9o1L
a/nhm04wHiubUxjkuzCb5+rOTWL7aFZKt4f2o8SRA6s0D6rsNHCM5lY9RWSMTw3UDi/HLvJJZHrY
PUjQd1SOcIOR+umesMjo8z+EPJ1Ur0QIN/qf1uzyy2Vp22rG2z+fj+bPe4aJzvIR2ptcQ3LAj1bO
Mum55tKQHKb5cvm8NxYGDiI4jFT1gpZpT1/NLW6UoJZDQ5FMOCk+2dNUSf9HXP2A9SzJOKlHfYWG
W2dVdStQuKDMF2jIEqmeUjdLK6qHitlOQ2con74i+NK8xQrv6Z34TI9WaJy5p6ax6fDzyUlwnBxZ
Xwt9Xb8ZrDDw8WbIdviuCgFRYQUhxaZAfQcFo4UH5gz1+YeorliOk0mjiVVWc9+wpm6+bsbfsnad
bKiTgBeYg/7QoEHeROqRcWpHYmlMJ3vv0Xhc6DEEL7/AybI8ucSVm/6GNKMTG3FCAaaCuuVHOjOm
RnhPfADXgzMV0FUZD+Sf6WEgqH8ht0jcYdbNNHuMVp0Qc3QKroyLDMTbxDuR6fHj4wo3YxQ7nA5r
rm5aSqM1icTYbM8qw0yTSqGggvYePUQxZsoppWbHeFacxi2NZ7Xz9lc+HCi3eIOAzPvgNUdG7aQl
9jVs/S54DZ6BvHaNJF3mkqwVITlxDhbuoFm85TaxAt4cuUL7WJc39ilURurVg1FxWmC0O+YLP0o+
+aHxfVCQCKCBlgfom5WwwX89xGIQ6hUFMmwnllLdyYY1yss2D1fBC5iI5BQzkBi2LkMVvqWvMJaE
AvVwGIriJGKq5/dwsLfAMtLRN1Bu8nPuv0lXSCimdQTnWvR1OaEt/b4t66JgjOURDTjlcC6d7vWv
wV8qoACy/uDRP0K24YAs1TTmz4JJDeaMEvcVv0wMRIwkYU+8BUcEOGyzwLnt1GGCvsfU4fgfNjmT
gF1gB43xOAQK+aDrHJUNSKVUBdUOPzNC5bMoPJLKJVff6eKzDLjyqrV1xBIPLnYTFbankC4mdVCb
JpT2JMK0oZjDmzREVePM6D7klQ6K8XOudyI83hiY8eA/XFS4wqdEpLCRhD/Ysg+AwJ7AnewPeTzj
cxI8S1xQQReDgxg2vQ7L9ekN53xb+4b6iaeOQf81afhEbukZ8Y/ULyO7nkfTakFdiceXvFR4twN7
pq+Q/1K5aXr5uJ1gGso3A733CFqyr96biAdWsLoW9jfnYi/ULIGOtDleiD9Z6HnHdUnO38i5e6WH
fbOHabRrmmSlwD2r2BdUx0gSbUrmu+LjI4iUVE0A2v0bRNXWDtPJ2kCeaOG6bMK12Eh/+PtnzN7V
bKz8ixaier1y+A4ArkdqLdzyHCVXVNw61WnhJ4kOweqixvSr4CS45BYKxI31gWNccwPm11H9IIdJ
NuFq8K7v7e1+QqDN4mDgH9ZKqgdTGmUFoJ8JKgJi4rw7ydROULvOB/loa2VE+kSKCrQIHao6IDPR
88vUUdJQFgr70p4Lozhz/WrycR4IOQsxf9+jWQWtEE96YG6yx4F4xih+7ofU9I08U8U0wpO+zCeH
OPXgeouKBxRIMIV+f6spPSong1Hj0a5lfwE7+AU0GxWd7vqj5wpj2OO77/HxZdkgFLlG+LNdzw9r
4LYtkWWAmzuqzDMIGdZCfmvrM6iW406hzsqj6MISj5EzZIPHD35ZpNhL91KybUsuWesB7DmKtktn
IxT6bmaioQJIYsFADE4wmLoQVjFXNyP8R9/0vhmKRpH0SfAI0tJHfLs+ByZFHsbPLaOMstahmU4g
/TkJpKyNML5X83ei721p3LxEdJPOW7W1RxrYfEM6i+75+MNUs6zXU/9JbiWhA4RKRmBMwSg0NReQ
/JoH8u8/8h8+ZcpnhZ8N35/R12Xea0UhUZ1Yiqi8NrPobowjDUv6rupoN+SBuY3phoLsYGCe/5NR
cIpxHauvYubRU3XgjNXy5xn96v+rZrRhz4JrFYgbRKQjtChB62QMKeZfIF+wN6EEHicGlmyPOElK
dfpSGXU+z0nUFCuOu074VjSh9ptaLve4+92Vkp0RfaKas4pD4X81tHzxMYJ2ehb6MAvoKo4sIRwM
kn172aQT8fdXrcZR6sfFWf4RyPWMtoE4Hj/1EaU7f4p70rZyPPakJQrsbADc0HUD5wiXvz7V7wPD
Es4dOoxqs0ZWOKMXU8cFcuiIQUPQgWDVqhS8DTt3rAIeVUJyNEQ7HfQ3KuzDldq6GXqKxgmDc9zI
ZXJYMnQJg5TwtcECDHbU1nzrzoPP2JoiL2UgFrcW4BmW5OK7pNbRwVKuQJaT5vpx38Lf9zCEytsh
z+DVrwIKH+kK0Jjjhbi2F1sZqrOalN14gqxmMS3E6vnQEaIwo5q8DYWFKG8oX7gAZ9eeE/Zk1jaO
IcSlBR/H2vLpP+4prPaHExtjLci6GN1SDmUlGDn/GFzIE2TCr+3vtocpoUQfxXoWHtNfpAT2hwdL
iYtuthQkxZRcM9yBeVBRG4Hk2fR3UrHgLTUfg5HEARNL0FdDk5pEKApeTBlceOFBpQJbAdYZlNsd
m163LhYP8BN9fSat2Ixz6JNphH37+mQ7hGdTeup343qAUpNYS/6HPhlWE7sDREGTde2P61NGzNlh
Lu7FlmjhqxOD6rXbyiXrgpoj2idEVgibz8v66iHcdfGp6mDzjpqbJTfXuXfqVSL36luN3lBYM7pT
xgtz48t7zrKOswB6obCNPS/NnqW967EGFPYc5UOEn78o22j3bWLKhlllTL2beE4mN9LPRkh6OpXn
qFBds3UbB3MfWwpwnQ6hx0Cao4xV1tm8rtQvHPgnGG/cg9bA9tfeu7Yoy7B/IyotwocJUcq8Qg5q
bvXEQ9DoJjCn3IV+FEzUIlbH8TN3+oqBhXfIhp5wTP7lNkaPZBkFKV7mGTzsMcKMOWS4loSTs56H
p7yc4hyeNlEuIgckiS2KwkmypO9VjH1BgjNTQkAI30Ku8TiqYmNHsyoKdDZbsrOnBDnp4kp8KQZb
9pfRElDGhsbAkimudQYz82CmATHm3RtT9triF1tmak+brIpisXb7ja+ojJHGjQAuzTvSY5q1g6K0
SlKWpI5l+/WaVfgIY7VLjuJN1X8HyqfdNVLf3Sqvn51b9xhJ+NEpejVQOCUPWwA6SIdEQ6Sf3Q++
+JdfzYXIuH8iUUZ6m8l1brShJTSFJh7kNg56UWj02vKpLBcYx/iCIwYPXnxYloVGGiYsoSMSBXqJ
PnMPcXwfdJNYT/tQNUtP9FF4OW6iqIERtzpm9ismRIHeMXffq9X7VutjbQISGfoQxKmyvLX+pprm
Tb/AUAxXVt9dSf5iLMpmr1SuLGz4eVDSSlEXEdIOdTP4GRWUx8+W2nmwT6esVLdc6ZrdOTal95e+
hJMvkat3a4mCYWmKuZdNUjZn6A9gyN9BKz8jHPj6rPhMMF1gjOwC2L9bUKHsCztCUSjC3cRE0N76
UxyZ1n33gouHa1zxYBkPqQZfaKKkYn5mD1SyU9HBQudvjk2tYDa0C1QGHNPRoYiMqQF5TzM8wlzY
c965D2Y6Qr9cgpemRDXJEjkpDfzPGrFP48uuqVaET+dKhu6KC/1dC5tNjsAHWCRSLRfSscNqC724
r+TlEg8u3arj5cuK1ranBmI3TOA9WmZoyxLlnBYzod5KtEy/KMcZRi533olL7+Sd+88KjOx4p3li
WZD+ZQNdMam7nrE/z/hIC0s/MiSzGdJdOB4i1MwlCcaFOGHdUpelkA/G9Ik3kuzWHkl6a4SZM5QF
bkHcH+VprglHHhn5quuzS8ryhic6veyDDdqCvd+66lzNo7/bN7kP6Pkw6veSYh8MWko9U3t+iVj7
rgK4szNLdaekO2CMJKHunLS/KL6AchQTxeD5lnzrxOw09ngAxPVeyV1XqnGIz42++CD1pwNlAASF
eZCUNosLqkBJ8n3RE0ZyIQqJQML3Hep2o9qXDse9IOBAUojtM/gcytGRok/B9wkEgj8+WE97uLWY
I99bJ9zTJRg+fiRT7tCKvFol89acAZKelkD6aZzFqYtUpwDxHFvU63ct8gUJ/SthxvVNSvIEGnS0
Q4Uivy3rMDfNXgrTvLAle8blf5rtBljwv6cjTiIbn5RM+7TQI4DzoAEwICsHLtsfG8sKpFvFTsJz
WMHM/BqrSEvJrSaImekYIfvMGjAvUNcZHgRbWgMAillRXMYcHKfxE5572aD/ZL3okIsAXZWOA1kN
Opc5W64KSenl2G8RSGpGX4qeB5iNWRmTtjd17sCFbT8Mu3u5RBxuYt1Ujh8RoGuy8QgBgZo+mrH8
Yz2rKm3CRmmTYpAzCO9iFTwjiDoQqfCQaoNLRsKDC8wXeyBqhPwsKieai4DtOj17Bx/c3dffW1Fo
+TF3247JiHSj7ajDxE792I8k2KzsHqc+eaOhc4DHNP3TXFUElD0saTTujG9i4DUohgty5RL1ESnQ
zibuIZl4dQrFmuPNR8o0uCu7Bbvkg/brzkdIPtY+Ti75y5E8AmYrHgRR1I9Y60z7COkJX3Frkm78
x577DDIYuSujkpqnbj6xhmQpIXKl26yUe3owKlXIEoWqQRpmXvmhWEhUrWeKPUWrluRv/LNcPjPh
iKT53JMjnOJ+5Hm1rYclvL7R6QWGvjwFFQUiiUNfhVie4JsyFXKorupeiN/t5eyyiMUtDWai834I
g9/OKvO9XeFEpEVC5eIi1Tpt0jnTCZT+3+7+9tWTEmwdcJW1cYaFzqHLA8uamdmXctnxSzer0Fdj
F3z1IjpAOsQQaK7HZtmxpq/vmKv+wab5H1MXB/omt+WgXiFWX8Wv6WqlvLHK48hHVa9NEKd89CnF
5YtMrnO30sbC5aJc5PrPzneHmizAMe9E6WNtOtHDwEiBQGoX25OlU29S4iZtuUKhmGnQssBcUZjq
FUiSL0Uw5oD37POFR4HAoXEO1OJYBLI5VZSBQyM1IyBTJoQPzb5x4KM36+uRtbUPykIz3n6OO2W+
9Q+O3FD33N2lki/DaySwroN/kI/IbezKD4mZXHStdcxkS3n4O8+c8kTDsPl0zMZAfx9oFi+wVK0Y
BdWk8w7Eo161cUVACplzyoybtlAaMZsUxWdlEZNLq7jJk5trY/HF6MJFbA3sTzSD0frRkVvO2QTN
qO3qPtN90BuTB1zjd0ZokCLOvI+GpZPN/XLTl8KxnwLt+SY6NvaNM9UQ1G4CF/+4s4hqH1yjmzXl
6ImE5p8heyODTk5kVyEAfWF5M01UK8Dd9EjSSYIQdg1DECVBkqXokSfw3ZRW6cZqSPfM0MnMVDkl
oNU41nqOp/tze58cyk1I5VuY+XtCJoig9u/rKf0v2Hvv3yErbJQvimHvEd4BZfSJRe0LfCAizZvZ
mA74wyyQGfhMLCpTAmy4IFUhR6kR0Y7SiiLFqUsJzFk5d6RkfWMSh2dUAWGIF+ZPctOZNJxLTAXU
LjBnt9wh02QgFarg/JVYxzUHIkEGEfPoc4S+2zuXQeEXqQhykj6E3hseZSyxsLFyn1LZzZFlfc+U
uxJFiU9quZo/IBE+/quyOyXL62zw8Y3qSARbcu8gurXD6nN3hq5PUqmWbeRs6e0atK99eHoty2YR
Po8ZtUt7RjwipG+tqgHc3dqJOXhWkRjy6J20WP/6cK5hLVJYVNpfxwwAbb7F3aWRPzcshbGSrs20
cSKVQGqt7m30CZq85UACSzOgBnH/I4FHx0JEocg/IksKKrzcBhTvY73Hze1kb8OydumNNXQAnbFO
XpijQWtpFeHnB/PwOvmLJHleLHmHkDQ2Zl0hLZvxDCxt+2dw/JXUw5cEmluTRk+yiX+89I7+p0qv
6JYRproojJA2Yb1hSVdXMZ1/sHzhUS905eCdSgU1vb2V5VYMM5niMF01+bcfzOg0MvCII+sBGIKh
IbKe6MbjU/uNGhSTVcdw/fGO/3Kr74hW3vo27Xg6pn/I5WtF7Q23EmTXi10Hdu07f9ZGVlrgvtwd
2iul/ECI/jjO9t5WSVpHeH4dAiSM79Q1AXX6/1SICvlLKhEyhnc/YRyBpVxddYQsjkWlJk9bpwbl
on+UNVx06Frt4sG4A3Xjz23KHtlNVkTZza2ku/rHQsqhhmyu0XOB7MOJL//832bHg6vsgf50x0R7
bnxVpmAV+hQmZFHvA7u8WpAbpiCD02j96VMjz2vFc8WS/bt5dLJDvx9ZwB2j56e6RpIrJaihJon+
mxMN7uUKgy5fce4xMLBz5ftobX9hPdgMnwieoIepqZwyIZguVwfb2enEHmlkkYA9gLmLydd//RWs
npaDzbMEx3RMNjGUTnXQXSWqHlVmaMHdPg4LT9SqWMbDfWXCURbxAkbJJdZAleOYZ8tokl00QL93
RSP8shEeWyL0QP9kkNGbKEq+JC8wfbt7h2Ujug39WaBC/9f20dVK0cM+gLQkkq5i10e9sCSTyrfo
TQD3b2TP2WjVhcIOFL836rzOf6y1trAw4hlJRHCfZKK+tJbjzSy/P0qOyHbR5CAUq2PEBw/TEO8C
HiluSxk9IhDaX8vPwEbQNgLNW4fZrB9V/C+PV5JMo1f63IZB9YRBOdpvaZRC3cj/0PVQbC+o1QFp
mNln/WfYcd1H5w1mqs37aIr9mSEMvpXdz6qQniu/0CgzVX3YuCHI4RvoVBEGrF7CNhrdgBufQTRy
dimLdsP6hvtQwn9W8TacmYwipc4dKiSoJG9Nl2k4MrVfZ8BrQnvKn6YISn8TsdoP8r3KqPfOIYkr
ZH++A9Nofw8G8lkf0atix9ff+Xt/vOPFJtYdKJ86e4A7+SvEHAOzvsl00virWJ+AU2d/7ss72MdK
V8C5OXEbKXSZvQUyQtVFGQ3KKg57QZTr3D0zZ87sTEBIe2PA717U82D90W0wp3/dCDyBFXFmJ9vG
466pFZDL8XX6p9PgRRdVUmQyerwV0RjlUJJ3+I2nddV65/JtySiOpfrp18vGGaQgrhMQvhTG/JjY
UaCxKLCv6vMqGav3Dp0jQMmAo6xTEGgSMTWpWs0UfjiyCAojnl1031XF02vPs/ayUfBfxqXWGzp6
uO+Wv+xEdas33XRvNnxHrpXu7duVszpZ6GkZCh07nLY9UuZ8dLbcndKkIknW55K/+TME3ko85xi+
mznpN4QaxjjmFhWz0EqvDBg0GwNBuXSjfiZWfBH4zH3uZCNIuKu0yD+FOfWGxtH0xQ3bYcWCzN6Q
GguT/MhyV6r3pep+5qX4KiuHZcYOVANK0c+v68Aw3fU5LhV0HIb09Pg56K8HCs/JKLJPgYsc4Cy5
Np1+oJ0kj7kJkcvoxSxtHy1tulouYsyYCbulzBsD0Qz8mKjSVXVfBLwppP7BXmWOzW8wrzsWv/ei
7E7AJsuOle2mSNi28klWcNtN0xtuyniV00Yo01q2lhJ5L+Qo+ntWJ8N6r3HVWDUV021VqIsH/y2c
Yhq7WrnP5ijmXXVbsHq9JojhDQ6xn39lWaKMSmOYlq/byjnCeq3VthGYOp5CtksoOZIDHQr+wx/i
eXn3VcNGxalwKUSsIdVB5rWfd9KkUdX12UJ6/CtDFfqsW8yPbbluLbvYCp220eCX6x4aaBTdH15o
wvWO5IoyTcZIyz6oHLCIVRN5EbHJqXoHGNMvA0VtGn3c5jrsqor5wDE2ce0NWLxC3KoU0ux/eAf3
Ev016fW4rtRYuC0K73Gq60a5tsJJg38RATL+AxaNC/lqq9eLTFl+CZYS+pgTuT9vUP8NuzoSQL2o
tY5njhrhu3FaZk3xj7i/4GC6WdPJrzuByWDBR6RO2t0e10CHdg+nDP3hXwWk/SCMujsYfieH73F7
B9Tnwz9gvwVco++VXe7rBvwfXMk5uKSthbsmJzqYEidcWj6ADHqMMNi3i0TX41NrRgbli9+qH886
s8MtIEYxuNoM6nC1gw3n6Wc9iieZXztHW9WgMiN1Df69mwkeQ49KTbfTaXyNNV85vIy9rimuYf5A
ZSpcXUVpv64WcEL8tBOINC4gMpObmooIfVV4HTjRTLEA1qNP/gatxSl6wXDpv/QNK6v6EmrjlIHH
aUUfxgZ75wpP/iE5IH27AfMUeCWC0egq/AVZEl1zUOJdNGrn1FCR6hZB28gxyN0hJ60kULcomk9r
ISxZfduGo2FmKDPDZWXmTF+KAjRebRqsRPDn6itvj/eV7eG+N59O5mB5IeJEtl9JIhFHmoxpYhi6
EZUHyUk9QdxcwETgxZnHcaF2WGCjDsW8QDIx2mai9XfURIrF3hCoamdfz34bghovsblaR1c6wURc
xXJ7aqVWuQ9dsCkSX/z8B1qVde3IO1hTgbradSj4fGpVirntug9jBTg29F57ZamvEXlxV6B6bCNe
C3cNGLpIlbcdKsG1I99DkARrwwPErY1mzkJgcawAXuEH89I7tRz46jhid2pJR954VDniy+ePWsrh
WYZefL8PaBWdJFSmNCiYN1JQx24c04vZwbI1OTkN86Nht4XQ76XCMvfua+mMpKDFCgazJ9N3n4bO
+AJ+Eo4GTBJnKr9cmcfk1UH/OkUk5eyekun0OpIFrAmFdh6imdlnH3TFLZ6vfTX9y2SGNSiTyQ0W
/Ek3xA9cJZo+3CaPvxfxbh6XNNt7siFpQTwe40Vjgue2XnXYyR1jZN/blPNyztZMX6QF7QxbUbo8
bWED1MUcIuKH6h3kvrdFzF7wSLbvLv3NmchpgeaAQYudWj9WhtKwUL24xsJY53cm2fCNOoOzp3Ll
lWscVC2GMZkwKhG4NZkPdKdUa3pMUMM/kB0zxqpoXryniGa9HQukPqU/M18E7i6RWVAbP3iCQo0s
+aD/ilxl4BKv4mcFNfnS8xPUP3AZMTYxFDKp6bCo6Yt4GdwjCkFuFx+yPuuxbHUZRYrmuOeUFTdD
2YLKh2EeORQ5eiwvY4m5HxJvCySq1aLb5PzJgFcuNBVuZacAnjZuETGy7QWxigFq+JwObo9c23+h
n3fcd1XxhB4XnVk4A0sgjSkQFZj1GSH+1RXyXGfnR9t54uE0CCvH2MIbyVPP7rm6AcYZZfEO2dZU
e9uT2Elgip5uv5RQQ2FRAwow0vPskzUIMLqp1RgSZRDhbSqFXVnpMWoN22wnLZhSsLzzvqJpIqPk
Etnxc3bRWFmspHB0hsOset/luBZSNc9PH/Lqa9AstGKIjz/QR76NCQ9a4rgbbsVUtI/ks5enDt1Q
xHZq7ctlzKRZlFI483+oPH13lPlBbqgGYEju+HYFsDZ5lgICHTHGReash/loWX/PnNtkrI8PEohk
Y3jHxQ2WmFRLbaeuE7twzJ7pwhrKiauaSbTSMY1EKRQv1Ntaon2Y48ukwgXg7XCJd6Y2TKSiGm1Y
gjC0+krv5UpdZkRS+0fZ80wuZD9doXW1pJuOZxxwOfw674xoZBnOs6J6ahoJQdFquvWLe5Q/L16u
xNyxZQJRMHq7hP2T8Q9UI7rhZNZ6UUXWHeKRoAIhLGhQRFQ/uKiwLXXDWr1hpMIWf1m2RM9ntML5
hZM/E2ygwnmmIhdJQj+9mKGFHlN/jZf+6IlWx2SP/yk4xAyBiEhs5ZegnoJ4VF9zCj5aqoGO2wr+
5+n6TgxqZpxq9biLZWIQzpUjlMXAlhYi/RQ/B6wozpxH3mwetRESi430axg3fwLHuKQQOgc/v4cB
ZwvorcNxlXSkmmqbbxx4mnAhOeOJxvvTmw7aH4sXSib2cbpcTIHmEkmDT5HYbEP/zeNtrVUUrOmM
jLOukp5Gficd8BMj3iVAcGz7ZrG5Twux9pzYOAZL5AK0LVX66PU25sUxpyOgRsdJ9yewuIkSxQd7
gy2LpSfDvLRGdEBmNd+UK1tl5NhchiBIV9JghjTE2NpD8mr5+vFubbD+0kVPfDN5Ri0H3rW4kIk+
I8Rdh7mVj2wzq4GDIHrbdz/yiBQ5NFQf6zjdH6COC2TmF8GCgY4ANYoHHpf1vfvYuRTE28BCQ9Gs
RvMFRmgPqt5pzsW9T3eRrjec9Cxqm1NMDwN5IsSEp/d8UGM+bdcVkZu+iXssOrc6moqTCXPvpMuZ
Ykrl+XrG44oTI3pPLA5jVyqgT3K10FMFT8FVbLAXiYNevjwvVE7pBTTZikGi/JvhwrT5YNiENIFm
5Tann/0wpv2mJytqfER2Gj7e6nlI2p/ckKcpB9lnf6AiRKo3C8EI0kOypl4aOLurcwRI/y8uUcqt
M6jHt/uBWO8ToYmP+yuFSvAl02BWb+3eR34naCfjdvaFYOh+Zoq0O0r/cErUoSDZvmxkGAx9eH3i
kAfUyJrHsMzw6sogWC/imHUOb96MzlU+ANNKkGIm4Fm7AxszOyhgSzlIv3M+GdBCeZpIQNiHMKXb
EXoiZXiQgpStqnb5DsVXKLz9flTQJoZvsV+JyJl7t4INGelfGeaBOEv0UQtrivfY5HhH7a8mqpBQ
sscyH3N6BTKSlh6IzHQxcBdLWf4bWq2eWWnuwmn/gIJAAepQ/T6LdTizLHe12nPWmGmTSzpd7PQl
lAeMdsGC7wAcg5YXVAHumVKTowpR5fsl47imcw8gFr+kMr7BFxUDXVcbRP+S3Os3Z+I6+bft+88y
zgN5JlzGyNyWSiFqHcSCpWfJfCx3EEAdH5Nm6NEutanajhx6A0MUJkH+E8NWkS4UFxN1JHs/XMR3
Xfhl4CWC/VglTNMkwj/m94xrSIIAO6cTaDMCXF83sPu+KXLMtz2Lms6qdsHUls7bFjndWEWmWO6y
EPzZBMM1j5949huarX53FKpLM40fSfh4jLg0744i6UxCye3V/nvj8lgNjlJcN+4H4CdTONQodSVZ
MqqHPrQIr6LQIzixQuZn39S9t94owDRI2qc0ZAQHdP3uOFepjjcy4W4SeegR3l87BbRdedl43I9+
dxw9obZDu7r065L2bOtawEtRxYEapPOGwc8b4Jw634nYdhd3NYSQ3rkBMr/RC3FG0BkVQQIlOrPK
M7aCDrNXSqQn6EvUzPWh+JR7XEy+pf3waOYkiU22aGO3M2rQyVFrMq7S98YEwl2wlOglPXZBnYYc
cIIcagL2WlreqQneKvFSrtiefOkDV6KWbP1WOa8z506nBbPbzw3s3UPrWWXKTGpH5DXLxcWWmkyt
2D/8Xl0C7hsyUKJnYPvxlEGy97wwiILUDste+sTfkn1G5jxFy2nO6TdN5K/YMZQkoXz3GCXdfJ8E
5kY3o2rjb7vFegrUbU3eDnxcfFsv9jOYnRT3JD7U0bGpF0KNaD+ESVxPrL3lqEw9Oa9cCSbdwEXe
XIlB5AtZDF71PQsA6oBrzPJxXxo/gN3cvPg1ZEkJGwnQBeSzTKHT1dQaioXVYj1P5l3ODRw03DfB
r3oYfXOe4cyHli4YrThYqgDwSxL8EYevN2mLf775bqO6/KHEzeBdao4aPDNTa1XajINyTjMey9Iv
kaWZuzduBZQactbcMHRQspBVd/SShGW77BZqWdYaKLEcvETcN23nj2AludUu3oxtkNrgau00TsSa
M+Et9IEt4pkEglPyyAt5CUDPbCwnrvr8+xdNe1rO7SNOUPnXDxixZEQdWDvRUZbxArS3XmZhciN7
wigV90dWmKMV40+Ok9OKpBP4B+qMYJDbw6P2+UoNOBuVXB7BXMnv0rOYCVRAj49q4Nx/vUc5m6z6
lltSu8qR0qcy1W9tfGdiEkgTWS5rbD3F7SNC/EGD5pBmrIMfLxWpo12E0kRGawoL3xrc/hCpnNR2
paZ4lNk2Di7FgpuF9kNiY63nYESRukKZ0B8iIigyah+KS3Ll6vsn2mstBi9+urNxuVVmwi+LggvK
cpL14nNjCke8XIJAr45pqY8vXNoY9JIPCneAXxXD6cE/LLeZF8bg7BCEMr8eWZFn1PrtQ+L3iJ19
Mf07kJ3A/8p5VUD5hBvyaewh3oJhyTGhokb6BX+pbd+abVlnYNKX3koNVyEAEpmC1UNRXXq00EZe
v92xQKxSdm7M/aDp4Qn4jr3T/G9+pDC/6cV1I+CIn+UMX9RfXQEp8jIi/8RpzFqxL/BfQdWmwv8Y
+CRTLZ2y7vs/PspxHrsDo9NO/aBZaX3MNx88fEDYUAs0SMiKgbW+ilW1VAoUtk3C2mZNX7jP1QOQ
FNFPDQBgjdWWl57iOb6mgbFzLq9gvbhRJNSgQrjolE5virKkPLUoIw52I65ndzDtJ9Nkx9oBsiw2
ktdwwEcKuVhBA0iQBpbkfESPgNHxyM1WJWJB4qzlSL9cdxjeregJn3hY+kneyoVuYBWCd1lCudGV
WQNjHukiYmrX+NP4P30WhvzxC59jMkuHf29aT8HPs1M/G45uGDvZHb7ftAo9SuymLKwuJ735ljkY
pinFVtOxhLL/2o61Ms22yFPj9ec6yZHpn/mcqa7SfU8jnItik7D3p3zxuYO12mJaMPXzqNmShslX
Mnqb3gWxnGANJYP2qdULOTVzLVGE52YJVYaZfsY7EWpjofdCMitquA5tPH3RQDd/UFSX0gslAK/z
wyxSbN0lGrCjDcinm1FNxkVjPRbONtWG7Ltoi+Eup7cfXh/R2vPYddXzot0C6KVibb1USxQgrXl8
Wsfh9yGNPz01VE9NNthDlNZcNqTz7Wb9s5fTjmDgOvkDaHQrdUhwRb2QIjT6vsmL0jgpZDa75uCg
gC4w+IBDQspF/LJp4FQhrToPjFNM/E0P1TWOBpVVSIYajtmpVqmsDVhwi9vNxrp+O6KXidkQWYOJ
NF6yYePlIv+6H4ni1hVYyZwqDtGbRlx1PUXaYDtNN9obEJxMYjlWA80qeddSvdS11lLv0BjIUa7N
N7qk7DHrwYmj0EL4wmRvpxgpwIgt4KLHFQyMUnBuqSmn4Wu2MaGiUgkLTRQKCmmDQ17tQit2T2BQ
EqIVMxqcyhMWEZHpT3KZM4u1OAvRGlc0SkGjIkvyvByEOKYLHZwIUZexYuaBS9NwRgTPSvmatWm9
1mTP726YLRjwC8ddjJ8BDzUd5ZJ4lEveYw7U6nkXm5dEI3rH21EFQYOPTClbs7s4e/zis68Wby9c
RVSmYHWI2DxplZBN3T1uWkmAq24cS6BUoN52V8sONj6fCsPGWtkhz5lV8QLLUruFK83EL+KQw8bk
SkPat4WCI6Roog9GXfy5djwG5+j0lNMzKOIcnhdjJpYOCClW7fegDiUvYf1Hm2e3iOft/yPYOdmM
DkxW+FrAQARaMRwEQqR5E7uPr3kmcNCNYYk4gZN9/KqGow2VHfD/IBnDWYY1SVEJPTVniUsMBAnp
DjMnhqTWRYVCZ8jRsnH3zBZ+PLc3v17g+5mYsMXtml1/D1s9YM1l3O8dQ4R/PYG49nPOFWqKt59Z
1uQKc79PYKmwDq58s5dtUbcrPNUzKLJihq1zZ8qSZeL/C2H4KY44CtO9OuO6Q/GsSlDTmN+bPtsL
s0JH7tqQri7sSnT67A246X17gSi2mQ8y5h2Mm8NwAbIbpZv4B8VC/N1Dq0RYnzEVKV3bsbFplVe5
2RqypeCAZtXFjukdvLFxFcofMB3URqsoUqZKpVZP6YpUtLG1BSvei71CUylaN6bKqIO36kPc57EY
bPjsxgi3YTLIxfJ5rc/ArD7cIcyQEHGzHAiWB7daebKG1x23i0MFH8bn+LrLfmoIzdw6zvSqnhIY
E6Wo6amsqlqF8QTIunF1wu7kSrf1JC/Z9Ac/zZyw0Z5uBeSRXEm3B91iBDVfdt3/jV12qdDJwLSa
0GJ452w765doEsxfaC2J20dYLY/faVt8gXsn/psK3jXOKWgEP5Je5bttGY3I3kGAF4kyscWavc77
wOEO0TnFnSaMk7kSj41r+c2Vy7cMwvuoOUQWibljyQaSJIqLXy9xQ3OBhVKvsc8jiwxf/XEw8u9q
SUK2NcX69dSib/N9lM20B9sVm1pE/xz+bi5kKfIAPo479fZHxkXqJc9Me1/Wk2YYI3Pe3A/QflY0
KgDxKm0S8YWsulaIl2LeFMUCbSe33wleZQkzqMIZefLB1VxU6whTgBeZvaUCkRTCwhw7vuIzh1gN
7AnlYhnLKDAs9w3djg8jvtvnPfMqAd+uQTESiVwK3rJoOqMnQHg3kqD9aKtPLDUXbvHSg/7qAclO
4BX40LeB3yO3SSXUMtINsgekGMMS8SMJ2FWG1lijQa2dsVHfooklzEz+fOr9rr6L2tuzwX/t2uoq
T+iNRk3eSh58Yj5RUnIz89R5tuRRrSYgklcnUtPTl7uLfuAF0iFOX1rNCx2EPl1r0myJmwjWOBXH
KrVbokU/A9dq659b27F7ShK/ubs4xiIDl/GjCttxG5bBKXyKqKiaeiVelFKoguZtyE2af3QYXs2d
eoD4Uys9c8Q817HwB9hXZgQcejHqeN+Ql38B45Q8IkXxSfZbVUe32UuF0ksLf4XQMq6zXZlPzNsO
TSHPuEWNikgzqDXA6CflzTT+0k2qnPIYrGsk/q2dFcawVc1JddvCyxpN4kyxTpoe3fWzYD+i7UmA
S0DBIorQU55miqA9Epmi+6+06rbbGPtXdaWOMCnoHItjxXGZ3CgtxtO1C37RQpW8VvrB4yaxo2X4
CnAaLPgqfju9bdd3TneZNz1uudIp2UozyUJpzH7UXfQrLwC2bjwOMquLKrG7FE0xwdSJEto/c7XE
gnvMZDoDzewb5nW76CPucLtY4iW5yDv/lug0oThJBH6h4TiPJ8PAFVF9vA+kpytB2hMR0pMPJkla
xmMmunkINPKZKo6++jqaEbTqkRbSevvkVr8VU8Ei/xlAr8Xx0PQw8HH48zXiIVuc3Fdshi1fYsTo
qtFrQUK2qZN/XTi2zV6gjtgiSB65EAyDC7GFeV0MgHVclmPYzucTspXfpzKVqUcrSQ+Or0Pywj5f
anBWhdNuJfPMBcjzNMMJ7blIoLrk0J0k5YbVDJT3Llo3odf4Mas0L9oiC78cD62Gzz9vJeeyQ4RH
TCpuV/1RH+om7af3J+zWz/2herAKYYNiYt+8GLJeuMkkrxnIIJawInG/d+1+1Nmpk9soG8ObqG21
nEmYzNvoPJG2Mg6EneG0wuAjwyIWXuOfYYmg43h1U1iLbOi/AkiNeSB8AupmWyOL/TlCfaKVuMJP
0yy+ezMGrquulnmj0DJvrdC406hmA3V5/4JaxXMLrHRy9aYNdFHTRDrJD9i4UtapX3RBa6citjS8
LJVpgrmhBSZovoMYWM9+ZW0mIGVwy911DzygjdOdIxx5xg+nmIPTKs0Grb56l8f/DQB9Db7fm40v
j1jtOCtYICrSLT0w/+VUEAZNNiuqgzRW548MRpg3DWZyT50T6aSENTm1mxJPVwyV5/LsWNjZVoDU
5pLF6Z9UTQorr1fZDy4VQBGWP2CUaW7LrWy33kO9A9d8MFWOSmKMvLrM3+SumBtu7h9XoNTAjHPB
S49aaS0UAMuMTc5ytiN9C0nS+14Q3tFTmcqzFyBLT/+ZN61CW6PF4r9W5Ts73VS/z32EPBmw2i8d
Qo2iiUr/mnJ5ZGPZ4pnSK+T8ZOIACDRyyslewArMJ/GCaIB/2sZv7d82HsA0E4zbagrpSy8QJ9qR
pWJQqabw51j7Nn6rgIdsokOZPOtxZRbh7D+4Afb1jwsVB2aeZtjRhiqZGKQNkp9BG+kGXfuJ8bDt
YtL8WW7CWMd+df9dN7LpKuvnS2n7rfEKrCqV/hslXXOsaKB2HmM21Drso9E7hieSmwCikrK5WXqp
GJKghJ4Phe+vEqzYfSvxFs4Uy7gwO3KM2vHeX3QZpIUATLtJOeUrXHgtBbaEI7rS2b8S2AgJcjeo
6uCjy/J9wMtH4Xda4a6klo50iY0dGBfH3NS9f1X9oUeWBkiPwwVLMd7vCjZDMSndS34+W3J6icoE
prtVw+nnN7yxLTX5eJyFJvv2nzFqDbxOmGpsnzHXr12L7V2CksAo0kw5y+dPbU9e3KWCWLck3s8e
OwvN7K+BHv2uqw0RkAcev2YUe80aH4GYilgxU7BpRoFQtzVmJi+yfIzcHXPAS9G1DtT7GWt//F79
f0xwk6vKMlD1YDwmz0kgXAM+jiAnn/Ii1Kt5R9lqXVxzINBxoNfOCNivSEmNliEscMn7sPBQQ5W8
gHEao3/R9U/FSDGTvZNKhIH0QXvXdxISBdBWMD+WF99SKuY7Cr5quI+Y76husHs37UEriGzcOxVo
cB8EfTw5whYjCrUVpNwTyUf/NBfnZunxpC1AsuNgXR991wtW1Czk/NGaKoHG2XMRAFQuGTXxflns
0vgqvfr3RVnM/gHNY/w4P12gk6+FSFeb/mzGBxhHL6UUboAGqBrZJbX9iWFz3pUPO0545HnbBeGc
rTy6JZWgpWtiSK8oHbZqoGjy5FFZXb6ZZd9XHuXRPjfS+VueOvSqW2LQLrc2F96vPeUF8bvtFFFy
OcVqew0002Xqu1lV7j3Z+4bepHX73cHiozCtC+gZtrFGqtFsDnMN74kxxCPoVZEM60oc4IzJArhs
sl75v7l0TctNe/4fLGuBWv/0AC4GRoSB/5bB/pQM1GURZ4t3rt7UHCky3Siy21kebPmo/TjJf7vN
snx5C6wJjPUKWbuCDbsZQGLi7gW5UsN+jq4z5rW4Ihiy59IIjXu2o/ib0bb+Aj4L5Gy4UDNAFkRZ
Ayf3xxsVGlXPhj5OIffYInhCwTLEQIw3FDjQbONQ6om6mGzUkfg2Kqd95KK8jfjM181KSnSdqdbw
a7bHDKeZED15j5ZhO3zERkFtltES8wkcbNH+37khK1c4n6+jCAm6dU+aLIqnIRl0wp9w/fLIddBu
MYCTC6pYMAK2mNEU1xx+H/HhQxZ13MU/ML5UkhYnRqiY5X3/Lcoy8prBaWL8dqQcEj2KQADKEwio
AuNN8gRZHop0S1wXpK5FCF4oUvcFNkcZnx4EtgXulDAFIGNEii2L6xhSJJWx94Mo0sETO9qqFHzs
iEdkIaIHvefqmgw25tEZs1Dt42L6WyGzFPfJ7CwQSytQVkKubQJX0CR4W0jcCthdmUeGwC/mKcG2
wILoaWtAmSXaOu/ZRebKsFAuWQPK3aUc19FalRShgxa0glz3S/SWmkrJ9kAsD69FUEu4zKZrIyHB
Ow6QoYD9kjiRGd04lahft3h93DeVbx294dQ3Acb8kSvnnATMz1/T9IjGSwdwyJwdRyQtm7Dk4ACw
lent1dO2SMBWaONFv7ap8SjZyb5MBEZ5A5zoqc4rh6Khp6RYKlbUVHWXeRKzkthowe2L+aK/dU0G
oFNdjjaxLg8NkRpRJQvI+g6fG/VRj3gSFHDJxuNjM6IGo9bHePpYPhR6vkfy0rfFQ9Io+fU67KlX
3yomW1Ic2UxfSjDLmJy761ZABj22B3VTdD0tPtIBH31A7H31RzGlB2NuwpCiZ2+hOC/X8WGCNssB
XoCFvGh5l0+Cq+MeB/juA33y4/2gKBT8ZIKYSONwZx4S8AUu61aSpPjX3WIUV+n/9n7I9GsKIyc3
0iMN2yhVnh2wutzvVDZWfGwxnRDte8j3L0Z8D39PSS5ftA7qN8pXXfFg8XFbrIDOiZz4aONl6WGu
XqtEj+sVTArjnPtrrb20YClNJZZOgBC/EAGdgi488tdx1mHPseYchLUgGqThBRc7umTSWwLm7ILk
H0egCExNklQ5W5s0ggXWhUVZFkodAzxFEcyoXpMDJ767l5UpnD860n4TE2TfiLSlDhqpXt/H9PkC
S3El1dRWks3o/CqnEGIfg7S1cuolV+bkdNDwvci11wUXork5G7OtSwDVfrZlc1sUx/BTueROlRPI
nEa2WsEcbw7RT6bIn3TSZaJFyW/cTIHM+l9jWhgXbnxJjchmgEfgxSvP2MjwvSvl1Qgz6SeokGJx
CwFK/0dh2LbUkaGVc/PRGUoLKUuP1+vMDjJXRqjNzOnIJXVKHyadlAq/9Hvu/iRnmgUbQLo7Y0ZR
NFZvMeOa3dSshFDl1SIMkFMrrtnwoCzdpwAh8SiMCGEAQXyeAjXV7t6U70F1lv/GuFFO37ijXwQ9
hoh9n4nODA+BcR3WtYwO+vTJmE8phoEcUScpxJhFZoWm3zf1eF+1ISs0CN13jJ5nvEr5h1Lw2ovw
zyCkE6KDdmK8M6yo8HTE2Mi14FmORJhCRaY8E9yTwyWbcvUfTrYTfwLibHMKXYRNn+4RtSRLN5yR
iXuOOzDOPVPMwzovXRV4SOyqZ2iA4IPorxEIlLbTciVlpvWnR4kbLN1TkAKm5CjJC3qGDaMKek57
tdTJvLqTidFr9+CtW3Lmxc2QQa2G8tiKH/IODIXz5H9a7qGiMfoaa2l6P9cYZGQjFVIArYuRJG3b
uzDylm6Rbul7gIoy0rNKXi0gNegMBCCH4vP0PyHf1r53Sdm8Hq9DsgUcbaFinqfKWF307DDr+jU1
dKhl5Tps/IxAZ2fA3CottNiW4bqRxx17yQoEv4BYDZavXnHSilJdgZ5C5Dk+s005Q8/AookLiAuS
J6dz6orc28k/vZQsGi6A/zDLHHjymRLvezqFY0r1k4OfKlaFABV5023LFBJWH2yTN4CFIw0Y3szu
ubN0aj4VeUinS6LTxx5ipuURg9QLEo8v+RlEYWRRcxobKPsY0IwRcS4LoLDALGreBOAciTmFX9uG
sQ5rt7EHEQtmHFuj9eWdDiYYzxBwGiwOwMybu2VZb6gSuTxMPVpYHJY3e8PAyVRmb8+doJ05goHt
nqdaTNILZjAZhRusOQqs2dgJMloMTnXtN73CU4SUIrqO4JxJC02UfDLwbKvMAXxkt3M5ir5RCJof
WZ/dDg/Qyj11nmI+GTgtNl9p48Fm2cnICxMTQumgdm195VURwmpe0nfJ1bmbv3sE5w+Lh2spCgdf
iJXZJEzXn5qbnpps1ofnYlCuojFKb/O8R7wznQCS6jFJjLyqWiWuZ/TWYQAzhJyleZ4kc68lsv0u
AlSTyhL8nsjH6hCK4AKdL4ylfw1L/GSIUm2qXLshx4oa89Ami4KZipT0r3U4nUOB6OxsCyvqQZyw
hwTopXQnskSWiDZKnePI1HrPSJkBADOGswJT4y/MxcBrnqTfckKKz7KvcyDuwQEqxHUvJmyeU6zF
F6XKaM0j78WAGxopPHV8S9vX4iA84J9JS9uUY79GHevB+TkbXwAbcJpXRd8DqWW10MvVCB2b/bqD
wPkjE0OWVi7CEPs57rpSF2yLY9Ms1UOtyFQvQNXg5NKyqs0RN/jIgTqAtV+tWYX9y08pLcTXVSYk
UNMQk4ASmss8dyINROQeB5s6ZxBISdZDHnxMyz7g+vliOHbrwsPmugXgN9XWOHbm303pgPATPvtb
iEqO1pyPrpo3lb4zpL4xcE9GwbjEG4Fg0U5EqelJuqUnl9dXWHjq5Cev1oQ9Y02x5lJLKUNCdykt
Q6Sp3uBfkDAuTfQksz5EB4+8QtvP8GqgG0H3keZN3P/4CIICD9CnvXPhrgaSRR1k3xYa/CL+mYPV
1B+lYoJYOmYEXvWI23qoZ3sgOvXOIq6PyoGIO7HbsQPbhcX90Q150I140e8AcvWZAi9ooMBThNnV
gwj3CReGxABgUxIlqhADYcuC61oH/lF0hmkSftygXyO/kC836usx2EF1eZrNEas4DnxrDBjiR0/K
YGEWWTxvZc1KN00Us1XMhxO9CBUDy3fYs69PWkVmJiIt5gSS/PVkiSnasp3NNFtwvAk1gRAAM+Me
3O2X1+mO0MPsgF9qdThE2pLwgYjiXYiaikxn+p5jdlr1JovdpkjcN2f9l/QtqErm2xWdCTWYtfAo
noqT6r/BpmTcdibhsMVkAoSVp+Y2CD85TZjS24I04KvQDKkAegapCy2OUWXeV072qwu+lJkoxKGz
/6Wu/xftukPTCkHwQJ3QFBodRWpptXF7CLvT/JBya5cH59q2Wgsn8qbIH6KT+GKiBDgShMLtNZ4F
qzOqsRlXSjVdRYLD5qNOFnp/T1J4Jff1MjdOYVUXpDXjaEIzrLw9v2wAQtNxdXwYA0xw7GskwfTa
RsY2palHi9xEMOb1yjg/d9qhf+0rFy+o2DENhZT2HWD3+K4GH4ugQH2fOXeFky7YAMZeI8TH4pFy
boiX07AbK6NcR3ZFrjJj6zsW966NeRqXaUVe6i+Rnvx32QydPtWnR4CgPET06ppOEk1abNRLshht
t3eEd5UGlsv7GiCPkHOnuikL7Pt576bpYySnUx5p7Btb8tR0RCSYFUj/VlXykxn56Y3UpEVkG+gi
a+dS2jVOrhmetvQj/BNqRF4ya0/wrzWsappgE/ygKVb14JZ+KvDiwgQ5iTE0LuGkYDT3P3OxZnZ8
WLM1M3vuU8UOUi4X1Wdx0Youa76P0mpf0zoRkSqSqtnVBXRpjRj4ZfF8unSq49ziBleOGK0ww2sa
X66BI1b8vaqyYpl2GJuzL+RmmquLP/tlsMyZtWe0gXolpVCxNKCXg3UDnGcm5t6t0lJ232/yPXgB
gYN8l0PfJUbA9q3LY2ZK4gpxS4G1P4LMea7WugPtV/wIkEZA2Yu7O7dCIN1qQNmli8OSUDw5T9ab
dPH4dBQoAHiHZlp3jSxyryR2gaX89rMF3ZOmUCNfTXDOYwdX1Ifykk/cNqxYacC7r9I5U4Da/IjC
gc+EoStowGZx1pkChO2TFESuoYqXNGCpQ6ZF1SOvE/1KjUYp+nXzP8YL/GCNMy7mr7NfWdBPNBvD
TFw7y01lVhZEmXv1zgzSPAcVYcq557zIgeMPIDgxieCLIlOf3l8Jft0JcHsaSTeb7S6iQtjGOzBv
Ub3NlqZOtBW/W4FpNhoyw0jkiWJyMvjhIqkzs2UHWUNNFxsrSZBu8S4wqctHhmg6YENe8BBlhnNu
/Mi2SmyFQdjzsyHGNCkHf+vEAUYF4xWyyKTxVEr2WOleV7aHpRrEQXPmFvJtx4/QBXGbTegTdsl4
4c7TFot+sludtYDch7GSd5qnuBNNqsV2W5fDwRf3WflieoFuUYLPMkqaB2YaD+PophR0FZacTsSm
peTK175mxcYBCdTUWyl+NPf65XAU2t9bRoFmQPcudJtA7b2i9GgJKzVcJxGAksmlk+Tow5clLRxD
v3q0lih4vj7uLlDufnV4/tWrrDU7pXlp0kGq07yZdmAkYiBTssJbz++vk3CmB6dCKBsGMinfnZj7
Xijq+K5hLZsi9G2sDB+FKXNmk8wD73a6OvC4v3gX9bpwRhzwMYx/PL9lrqJf/woBt0SEQFGPJlIl
768ji2/HGni/xeIHvASKeFYmkQ9OYiWRx/XNcUt07FFlhfMngCtjHjr2tbJcjDdU6Nnh52kdk5Nn
PSOUdUzWjGh5MFWXlAKH0banKTl5AfIQY+jIyJM2NjehXIchJy0VJnfP3SHjEVQOHmy2NXkT12Lx
IH4wMs6M/MwpmDsJTQu9dZgmwleHwfuyWb19z32fmNeardifSPTgLXsSxF6o4NdJi6dmryuHpEVc
Xcm2RSO12EEr9CMdyHBDk+vkzpF+r4FxY8xBZj23eQalUoRXsMftceXCvS32PAa5lAKxx/1JnuXU
UmDA1AaCkWY3mHQbvzInpOdROQSqNZfeEMl+LqLWsiZmKVmnuL0hqBWV9jRMQUObtipa6kUmtHBj
+fAwJrCAel7A0twcD+qhF9/qYBtKP4LzxrGpmwzHp2/2OsmqPKuQ1K/FIPRUDW4RNqh4aeK2h3K9
6EkEt0lhLlA/RgZy7vZV/KE15nwVob+6G5IOXXLxcN2vfoXXg4AYNYQBO+B/xZTFaYFeRx3dTgxg
JX2TMkQ7oM8DOtyGRkteswVjMV+tJLqnIdPdPBeN1lcSJV8E/L0sKtsZnFn6O5yzryrlV4Cdiyoy
p3duUg4GBPN3lTTcXA5bm2uRYgYwer0/KTT4THwOenzOLC6NGo97a7+kAiTJ5dASpZxSe6drsNV4
ofrEec2o3XOScO2JMl8HLP3vYafZRCrwRQoPzPeTPMZYXFb8ksatxfxh7xn3vGa17He6oHpOCkUD
VG8JU+PcoxmuWPJuJjjgY5GrcjGoC8wM8FVF3oowc9V6QfaO9GImQ/an0LaJ9v81e0xg0Zqp6BmK
GrVfrA92ZFl1bwM9V0UCAi3g0WHvxxQsGVIVv3FAADOZ/3clTxhdyXZ8ruf/TZvBa93DkbQ0Zw3C
dLk2YHKDt4StPVGClKFV5XpQjB/wvKTyhxdAaR0wqX3VDg8lkV5LqJrZn9J+Rg/4cSD1CZvKgybN
O4lP2fDkgA8Hbu0P3HOTT84HYCq3fnUlJMdoBB9VhjB6+XgjSKZEaQUha2PDohzprmqyZRm/PS/c
nmRrlLbvh+7/Q2sQNbW5lSqRj2Mv8IhwK7VLcYvCtx3jngIY8fBz0mrQqDGaCB8hqtb33C3B4M6/
eE6wrfSWYVFnPPAIggEtvHpiRol9kIVp2DF4qJQwWHJv4S51aI+MHqCpazDSS/Jml8FCclnVfdAY
+4BaqFyfOSzS3WiMdCPGKYdqex9Bi5R7WGPMqwIgtDxemcExc2T0OYShFW+z7MFI7cOBrcP8Uipt
MjKYO5/Oa/cDp3FesEfYrsOS3wwmw4iHJjY+t/ukMP44TFjg0XjGpiikbVQvQshsLayYT2HUjd9F
RlyOqII56UgWLvPnYTsDkk+LGFB+mBgDspfNXX0fFQQ83hQ7rexItLQd0acojPCnOKEOat3Bdq0/
yLXtZqGnA/eEN1XYc9+doka1R3M2hDy5ZUCTjPLCSHRbrBKNEBAKwoev6/OX9DBxUwnOlYpWv45M
9zDUkunTWQkO1RKUBnjSnDBVBUj64KGbi7T/so4BOarEZ2L4X0lKhW/wfAZixKSthDxa8hUl/eI8
VfkALKzgCruNz+LrQpLcYu07x63MU/tC8+xYLu98F0sOfKtLSYSNZjYtzbyZ9p5CyaXb+CWzh62k
4W5WIOPJZhbBvswyvaMKuIIpDr2YvkbU0VwfBPvoua4DG42gRx7Lpr3kufmrrj3nMttcgIYXmtyq
BmWltyadOziFpWdeU3EOQXnqB3phR0Ybugv9TRZmhrXi2gxM+3xjDQQ5gFchpnuGepH38ND1ZqpG
D9EADvlS/XprHAJuJMJTGFgkBBp4mVPZiTCfudkCevW/J+4dyokfzcJNsa+IIiylZzJwiZNMssqS
TyVqYoSZHpgsQxi3VoEcok/BhrftxUuOQqU8S6rus84SoafKGY/uYXDG0BRNmyfpuATaQsxRb5Iq
8fY/HaXvjDh4gOoE6dLn12UmOvLLP0s9SF/FIHKEOLuSfhpx9VP5wJmi+MfTsQUu6PP1+okms5JT
QqXR1G/tr6HWtZv8OGMOvO4p5ZQviuejLfYcYs6x47uEOpYMwnU2vCA60OXiVPGLYkX7mB5qfpu0
RdjWvetszYihXjA3BjF7KApGZw1zpOtXQnmhnoruH9CGRJlVu/54E+Q/jLk6iZBZw2tfJ92L/A/1
P8/QRDfKHbgSXPihETNJqGRzlC0IRKNp2SQTuTvOZnOkfWDxz2aHk0SIsnc0WJ0OSuaF74CgByZI
emTDSGvDEKAqX/UnpUCfRdUNLYJd51RYB3WBKTYO33j1xDPAfDqRsi7eAgZbflO9mMsg4KJWKZUU
+cKdpk2Qdpw0g8k6Cl3n0krrJeO0jtWRgWgyJkz4s6rgJEb534/NOW6OcyCKca0f9iI85F0fGH/w
pl7kETkwmq0lPR8PIwIJ6B1WxA1pwB6NjnCdRJjNb93YDO9/+qbKF7JwFRuOcVS29NYO7iyUTOuu
vDfYorokEvuunCDuLIVpoo02ysNHRTl8yJWHWQcbVkgm2hW9EI5O4vbFW3FEj8p1rRzaObqQgXhJ
Ut8DYAmitg3bKRtaPaB+pDo1i37GqZMe+7o1TBt9Ggej1B/uGsJzBVW43pOCBQ80QqXPLJBD5Quw
XBD8ssjErLcCIbZq2G9ZcU2oOXZIGppGaQpdEfrJnTIsqqm1OHE5p8tbKP3zu9AIeWHAYea3FwRq
fy/1OaMXWuPXCT3xkQiBFtEIGuKN+Bz/3oCxM4o9w9QRuPzrGeILtK4gNYl4zURDU4c6V1B3fJ/G
Zb/MHHEejSiNZTel8JvEOC1LNSA6aJn3I0MvMWL+a8bqHEz0rSxmS87K6mf12iw9Ds4mzo8BRIGY
20nXsLVBDYGDFfrpEXkzOmHQkP6kur5q32bivstCrbAdopB3rQautVlppP8he2yLyhS8XLQBMCjR
+lFqQSwY/WUahqAjJkLWugBNxcMD2HjssOFKJiJJU5tT/rrMrWW+9lJEqQVQEC5kCCg6vdQSd0+o
IAgps6spo1T5TSDSwoCrtKMnzGKmf2JDqwz4tDY+soywIYOYXAHG9dETDo5tJQlt3v80thLastjd
23YAkKjCN+wCh+qW6ZjxGn6p18/Ib+aUDahSGh5lKzPkLtkKmleN+Qj5NxzHuJ69mN2KQIEzfDdY
6Sq9hM2nfSz+FhyUyNsqSEcUCskaFTDplcpyGRsSJpzOxrmY45+p200DkWfU3yAg69qgG7KAr4UT
Koy2J3vlEu2+JEf644K/dZbfZvS9aJ1VzS9uBiU+G0DCh8sfU9c0RIxeEBzH3x18D8wnhYRjzn0X
2mSgz+1/41lz04FkjtpgCI7Ph6LUUZA3BDlS4J5x9dRUfaHSJJCRwJny1yiHtoXEhQbBLuTtd9HO
ytFzZ6/BQl049HNsy9LgKYLD/rIn/0zEkrSKBFYUVtQ+Nk5T7DOihrIMzm7TaS8UkIDO8wKjRFw7
Z0npXOp0qzav6RBNYQCio8xBBazZ+yQ47fW/gXMAxScU6tt85D2NGKvFRdnI9ri0zTUz89e+DwV8
7xfhGmGnin9HpWkvPrHLrCN9qGRuClmbs4J491I90QMIYBRJfLnA/50WQiBtHwRbTMxXO4JgsGhY
8onjJOBCev3HF39RgE/8LzYz+2gzkdiGJqNAtHkrcQXQTvUh39i3QBvHWkzumBNkf0/QQchffkZW
ytHpaw2OPXE7sngtvKaLULCx18e3YyEHCAW8P7gKLBlSzlOyWIge6ariMho/tlpGlRdurYALUSbI
rhrT6i6Woif0r/5rgZrpHMpqE4Drphdg4AK7CRRx9mr3Qm7yRLiR4flxZco1vZLDVgeD5Q6pUqrL
cgvwetBT/PtjVQNQ8tZKRhbKWAkQ8b3lSk1OZ+qJ1imbnMxwEkpuJPviY6jH4sN7ZXTAu6sCAbFh
UZOdpn0Jmn3vmcMynSwtEGIofmmkkqMAXqdDfn7QKcPXGCi/6ZwsLE8WLNn+OCdMJfCEstwyFAJ7
cn7T2py5rKELo9oTw/MX9WGkRZkkHRvtkECDBcbK4dh8GHjBI7eW0JzGuUCKsRqQtkf8mSh9k+Vf
Byhsh353JaK3G+/Q1xW7ayTGtNvfUKbZmlBkZUOr2MPH5fbSk6O6AjQxsdi/rCWMJR7gxvnkFtGl
lGd9QG38vBaGpksF6HSujQYSeS5vNA+mwVkSFYSZTQBDvzWKTr+xLrIw2JFqVPGCbb52PrJSrU+G
p30sNFI1l5SIMkR6yvyMBvQILoeqU9EPiv95yhf3QiPoZx/w065ILRkQr5WU/d1kqNb4r0/y6wcc
JAUapJm421lgng0TE5psNu7RXW74k8Z0TWsxeOBSCzj5w/ZJpXXz2KyZlQt/0zu4SHMXf03Zm2Ks
b8ijVn72kiGeh3eJs4EobPrF+NOf2hLAVm1zEItzeugUogMEiVBLEoxa09ekJqYXgjwh8Xoee5lV
cjhsXeFd/WzFSCskwJN/PRv/eYs/Og1Bzr2TeDlxsR7GN1odG11X121b7zTpGoBUkLB7Pa6pR8LJ
qyT7vatpnzi9TbMz+f+JGzVC2JLGKatDWtPVgoPVOLsXSeWUf33KmqlPh0ZSyPZ86KkoyTV3g5z0
WEvtWaPJublpdrVOp2c59dPbEo2FqbEj0uuOxqsDE6r3CZpKyupNV55ZuHWBXUIZfMX3+Bs1aEhG
afm0DRk/DXmnOJCeIukDQ/nBLFpES5uxlHpX7wWZO8f11CbQBKCcoKox9Y59b456uEZLl+gUQKkW
+EVsdzhshuzxh3i1b3F3F6cx25qkUKnWUrS0rD3rrx56RMgO+Fx5yFrHY6Jgus3v1GKGkCqStHP6
rQvDxWmVhzYRrFbZwIdObBp0xmZ86P2Ycxe+cokLzNYg70IUqncAyVENxKOT0ZLACU2OG2btoCQg
PUTLuKCuKyfhuK0hfgO7Qfahdq4IYRS07H+gUdC0FbTwp/vSyLjm2xVeB8nw08kTNc4u9B2XnKMm
39FgqeAQrXsER4bRhzulvhg0TzQRKNgjxbA6iaItRasqV8AIUnYdIos2RmUSygydfyaTUSTTbtU8
4jC1STMig2O+HEN1ra1ZyIYUHVsz4+GSbKA+HQgchwN0GrdM1k+DDbKjiKulZ7HNqzIvAmIqOxdc
W4thgG/21XPJX8llE4yCGgocHZrTNR3XUJJ/w7+kp6L0kHFDhLwfEA/ci1VUvfWjyu6hfeIVRxEp
VzAlS9/GE5LIeSUs1dHdwRlTJJaA7w9qshzuMVpO4dKghId1p+1dlLadgXEymfHgFTJVlt/R/vhB
2Zs9Jy1Kfnsrq3Cu/WpUBc2n5HebxoiiFMWjxuhvdSMiE6edMw4XCT+BGyys3mM1QV8E3QNcPZ9s
xYjeEVJwhiCzpJCu0K1hhwSzuTa9yY57yALxKQtkh7I1ZjdPxJ/RnHb6prqWU1nLBO2e//ZgwQGr
fQkMnaT6FEHDvLeMC6mBKMdRiAjsyfZGZYhvBYC51usMLBNIVVp3wmgWxJ7LgbCpYdw6Bl+e5DYG
jLeMFcy+qF4iaP0si8Gs8zbVggVwMn3aP+NZVJBiM4orM8qQnMHppGMME4LuguSh+fnqfDa1+jty
Z2ePIafzKmSnQfomsvMShK3TrYLGmX8ne/qNeizpr1Uol+bVqruk3ikGYQHnlTdjUDqUob48fVki
olselt1lceV22DS8iBcGxo8+6SvASd+93DAfVKlV7Z1I+JB+CRvt4BuZvfPlw//7sOwN4ccPV/t3
mBRmUzLdptTbIJ+b+KX6uUxiOcL/s/bUsAtKMxHlbSdU83fnsubWqGouEyeHLH7nWvV0FYoG/XYq
cjqOgDGx0rIjXeNk69/h5u9PBQtOiR2jTCEaH7Rn+AjH79yhdxQmBkdoY8kMY+Vu79dHDqA+5VU9
SCeoTzGEZoJ9+FP3pcCI/przlTqxhmL2V5EOR2/fvTPThHj+WAxBXhjOL+S3U1E8b84ykDmxpovX
zGPGmqwY0EH+4JoSP1cBQsXivtJdQFXbzETHJuDUWimN48y7Gbo4cHRqb/n0SdLlSjNAnck1KnrA
CajxytYJ+UNrWDAzwJroxxWnuaCJakQsXQdQC5nZKxHGZcHZG9zwH9vjrLH82IxY+VDIU3h8OFhN
nmsH+MY/XOTkZXX9F0QelOzKWFp8Vjun2PO7HQH4mB+W/k+mLngEJTIoCiYwf6Boy9fOWfNDqJhX
QBYyeYCWbt9D4rEjsCHLn4g6vQZO0vZ5YbuuDa314QtIswqbS4YLIILua+aT0SRA5efnyKW8HFJx
2mU9RcIWtccScWCgaNo3rozIyjSEZB/qsr42vMXNs/AQKpBXOMen3e9THAMXNWV5hZxaIk78UDpy
axnnrWphqwRbsRglesDzuToo+NRtkSfy7cA/R5atIw5yZdJucBtAO9u0iGX6yud/sUTuvD/2R9cJ
UsKIcnFuvVBsSykNEoTu4HcOeGCv2qUh98pEW2gYef3k6WS+QSanjSHT7a6/cc1yGO3qO1Fs6urR
CumMIW4RaG+5FxwCAxuFOVucI9j8Semyzp5keVIolYSFDXsCJMuMyzNKv0MiuSS0FiPfa6rEddKK
nsxBITEmwFPdyWV6LjB+m9PdvYZtx5EpNkg5PsfV5Wmt0CxnUBgXgo5Z2zAi8Ll0UkNn+mZEtrA3
ypgUUotZkZitWMYx9HHoAAHojP9WunU0bZu3/UGWI54EKZCECp1cKv8zBguUo7xalc1CCQatVcV5
2FYkvPFjPijz3w1bUHVT12y2xJAWGdQkPgJjWY63s98+2mGUs5a+CPOhJolBBhXk1qEsjrUD14T0
SFXgok/OjfysjpLEWLGqV+kpOVJJZ4Wwovrbkrmlt6TOMiAHtYiAEOCCZTqCGJkjw0K8hoDXKJ21
d/IdsmMw/ovJkThSj9IYjI8v9e1lrt2BT8Wy4tk7lioSU4YtdJ9AO3NTDm5uSbPclI8s90SbVzlf
Jh/pd1CM23BEJqjLbaPi8x0Xi73oCfwaiuBBNLrgIe+yCGCnfwazuMImcnEjBy3Qq/MgJR5O/98g
v9qUQ6x+bBAktn08GB1/hEDj1Qk9qVT0fA2igv+9j3tpLFwhenZbwG+XdwtvYH6gmTFAXjQvt2mw
31IA5O6f6Xlac+qOE1bgWYmXG78JB5rOavGRPKY3Zp0GIBLEVp1ZZ5YUqZj7mDIToGlQ0amnsokN
f+sevAsD2mIfqsG7ZpXzMAgs/q0pZUEyGv3S1tVFYqtGcaLPkKSnPCbmyU/oqZsCDpQ8ypYlBMoE
UfKEwT+bs/DzYjeCuts2SrW8x+nOdwa40ilJC1dOpoAJ9W5yMxOJUfnglYrv3db3iWBRUAzEni+Q
GY3OH/Tn7MSHsGDuSswmna8t7qRMwDe4c4bBbZ0Bvk3IgyEcDT4B7sw9ALW28LhSc8S2dUGAc9re
Jx5BNwL7Rsgl9wIpdK7x9tPFOsMADlFk8Y9q68nmFqeVOjp/dsWA9ACpZP4Kr1IDdoRvfmAFWtHI
i8udhdIULjC2EyRCUswbvRBKmOT1aU4wG1KozA+eHkrnBlHB2VRO9OaCfkG06RkUoDPa1x9/GnyT
FlzzIkRCtIeqcuUWV2n6OLn8fIG/Aya2q4zNxBScN273lf7FAsk1jl0b15iA20HwDxyJ3WVSGylI
UBMmljIWtAu35FaNp/qVJ3unGanxw6gHSjgrY79eHzLRhaP9I8wWAz+F4aIL07i+RXygZCNEVjkl
BsojmLlGEqrqnlpLmKL94P0oOUr+nzQ2ZELN0EHnWpRSjcgkoKSGSVaOszfAy9J10VBdyFwBONPW
LhsaPp9JtlJdUXFFVpxzgJ71m8X9qYElyo1PLmcs2QZrq6+XiRFF2KBNtxHKUtbaAz2MY4dQmNdT
F94zUSJvszIf0SX9CTd/BpkUE3e8MKnJ/i6+nXrZkQdsVlT92/VBdYaVMMysrQSr4W/9f36p9RYD
EO7OiGvY1LXRkEfNHxr9JWbYJ0EzmWGGEjsOS+Qmhnw4V3uozK3olJPfrrwxR8nLJln6qAFMwvnO
WoCCkuzgLJbsPmDnURw2pVnjf14eYk0A3m/m1m8qk2n0WY9zIZo1TQKBsTJ9uaFO+8u9nn/HQCtH
Q5NAtKkMCwjxi00Ye2T+So9FVrWOUESqy/463VARVY93SBuo5VK7m6OaZKFW4n8ZYgpioaILftRE
mx39T9m2C/N071Fapu+k42OTpTJLI4xyVOLM0rFPqABqZUNwuvUoRaeZz7RaTu90HnF6ar06AIIf
mSiK6YE0I2aAFjMYei/bL2wnh3a3M/kct9O4fOc73ic805VdHYO8fmSiD630lx4mLzxegdPD16ya
lblNr/ypj+EYjQ00cJVBDdfh4PKuumGAPvUsd34TJ0YuPOxBl3TkelxeSwGfrC+Wg31bJCGIvPMg
lfZRJpr0f57JqdG8VsiymIrOK2InaBSIIYvjeunkaLxZIVCX98uWCcC5M3IOPUaslmCTq2aBudA2
FRKihyfeluYW3R5jLudfMMp8iwjm8XA/p+1394mo5rRLiRZdiK/3rbh2bxWV/ckSRWL5j2kREFc6
meP5ZQCBr1c6H8ZHSxQai69rTJJgXNIGyt1Y6qAUFij4sePfF1lz+aUlpR5rWhwKk5IFNOifmEMR
HaTC/y478SIxpg0g8eoHWVG8sz75os0V2Uq/0R5uj9+NzhaG4Huooix77NtZiAnDBk5Nd/jHQv/+
pXTlFjOd7GjzUUgKyccrTziQj0BinSYxfHL5kS6TH5wGfdkr0M1FjRNnaO3p6vDd3TG42XqvnmKX
xUfSiDnpTYIGlt+O5SF8krxom6AuCzzK8RTdobkQ428w80wWII2abPEJneZQtdGs6yiB6xUOT+C6
PIQWq6RriFqWSmsSEoOC1MMlrWK3eRafinzU7ROf3XHJXMpvfvVNFmwFhqI6UnVxzpbNEZduIdDG
7odFKP5dnimHdpj8Qd6tU2mdXI2sJ8OMTo41TksqePBpqI3RPanNMkjBCbI9b3UEw8IGxq3eA19g
t6QM4j/2was3Mtz2hCUi6wWiS5WyKFTOt4D7KUTBkp67EXfbW3Tn5PCdkB75BYzwkzEut7Xts3l0
vT8THSKtrg4v3esXBB4g7RMTFK+UyTq1dpymSTCzgNBMvhl01VWLjZ4cIDTVydZeWuLkl0g62yN1
7SVDpMf3tkSx0/vw7B/z8EGQ/OJ/ZuDZxVPZAnf2B11ISIXzrUN7GtginJXJXV4u1p7g5Zm39e2e
9+5RQPMDNrqFuvBjW1hApg4XIEjDG81iJS0FHdz/B3G9BffmtlI3dP2i3sZVdYRGyyzV/2BAcvoK
JdZpkwwEKS5sONZev/4MO0bdOyY3/hVlmYa2PiW6pNIhacfiy9ct9jz2fOdtu+kxk4S9mze2ATJw
XFW7pJOKa5pMQk9hIQnlPiSLkyYjcF/TVQegPVw9FC9eU8TZu/kC5AxQI+bKX07PbFBgYzamds9Z
jMuO52qaYT2hEHtrNM1IJbEMlVvrs2xsJL9+xaYWUSbGrxzNJUYE8J6YvJ6P0xXUWAhHI9TW1qzS
lJtNWBZGcy5YD4xCeXrhcaoE0BM8nsPrfXxhaae13kSwSYubXp2V1Bor4HIiw0pIie2Cm0ejI5F/
WsRHydD+AdSkreU11F8hXUxLvHzp8+yYoXT1WQdTMaLf7z+kEwTF7yZQp32u6pOsq1zcKeMcofVo
Mm4CrcmqAE5RVfRAhGNwJylM/+7Ix6nCF/720PRQp6GKkzX4mi3xTcnD5vUiytyXXBFUtQaoaE55
8P1znim9JDREFPPT9Y0cGvMVa7TCQspY99FmNdqjmfHfPljDWs3TQeN1rZPD7pfRYOoYJcQVGibA
bCugmL4a5qIrUzcSMVC6OWnO+sYqWqw2c5KLQU6jPSPbb+tYu+Es3pa6AYMSF3Iptd/kDE5SOwtI
4gd6gJsf5XZtteGQxGeEbv21LNghFSzNEU6iDWSXJNdnP0fRhOsdL8engnyMfGb+bw+kvX0by280
W9EvJF3Gm77FbKuqbFAzUP121NjdpgJuPEkPZGzJ3Zz6029f57oHxxEThT0yGIvwAk2q5wCTFWl+
Wn0f0qxGKUZhplzUYLLG1Gc/2aGiCHoSJKzDqTRWcf6NCfjWfrK82gl+X2Et8nLgZLqhxOKgarLm
Lj8jXsQFzzBFNoEPmp49DmcQsTZEd7aZZBOGU81hMiFA3UNj8faZCGTY8K7C5NunjQw7A1XhMWg/
Fohn1SFAGkn//Q1IZGoswtxPrghMI7t1rHnV06JOsmrgWX8pHcmNMGR2qzKCtmDA8Gb9gnba/QsP
K5h4e1pxImGYjGFQH/CFj5SCKMlmPWuiYy9HHcgM0FUwrx+3oKrBQXiCSd81bLmudz1LrS2xBY3L
VpOmLwqjfyCFO+6oGQfRjTmBhQVz9MJ+OvOU/H4eMsctWdggetCBlfcCw4fnmVDT7iMFpiSzhtIM
EXHbcXZ6zssW4ncRZAi2geDNQGXs7YeNgcNKERZe4xq5iWP4ZqS45AVqDLH8mJzF2XgU7Q7WlzgB
aVqkI0eVnhs0qB0mOYsVrmWbvVXBh0k5du3tmIay3dnWSOQq3QJ/lqZC3h33z6Jy4NksTlqwmBSj
q4fecx0aQpDTVUGBr0wNtmMLY0pfGfq+7d/geB9H3ajsFD3XP9gKaO27y0IpW5y8u8YA5uH8Zf0v
6sgQwhQvPnuk6DWh6W5df/u6M8RrgRVq2pWmKbxnM0l+V+mbtlmkTSjtOO3qO23o1JkSzrUUBlYA
oRfPf2h98E7rvxkuXERFxTyzg33XNXf8kiKQcLq+rZt+/W/fAtZN8nm8xEX41ZNt8lUIacQxM+TJ
8LHZbthE3oC6+2Zld+O7toil73dNp11VaIQdE/5PAzAjftASEhvpgz4lKTiKnXFawURDHvbXnxMG
3xFEX/tEZvV1R2Vb/AeIVocqbhXlcrake2xP6e7RMT9KZPq5qzAlmC42YvYB63Oa0Jb7eJF3Ttng
OzeSSGtE3azQrZxWPkmlZ18n/8adw/J/I8BZpoa1FQ32+M/5+nrWVSecXUhCJY7G3mvXjeXrmcSO
PdvOX9VdQhpf3H4yE/4ECmIUNCkpsQsrapdRCjL54VBwa+S28QHPhdNS9ObFsGhmvOAf4zMp0H+C
d4zKhSVQPJrvOSvbVJC91RoAkGriTd7gk/AdDGuvI6PukUWrBdl5pMQAuT26cApLLGKCY5KD3LJh
mnk08q2jLiiInP3+mnU4jNaOAxvGJ62Nsp371n4VO8ZWjhsHOnQiRofxzZwEdg6brqnacywf0FQr
i28R1szIbQi3nEMDepqxBt0QAKl7pClHlvrPFU3JSKhwlLRfY3LfulLIJ3Pd/ZwQsk3uoKJ9vWo4
FM4g/zTxzSC20XjpyqpfH8gLvbo94oK3VyalWoIE49HKlnesL0LHDQje47yCir+1hAtNFnlY7et4
6+zrq5yISXPUNlLsRr8EVwcVeoWBvNXNoSMpHHaC3vXtBzZ75o8Ns2eyuzHUFvpVN0VarxWPe2Vk
Qt7y2AKMJnmxEpZkGGG3xcsy90vGIfQCvQNbK6p/yaxFHSb3p2BnE7jeSYgVrC8RObBWxcNkhSmh
s5w4yFwiHReRFXwoOjKb6dO9uOWCgrEnJ0rWTk+oR1BwcGwzkPjPb+5j1tsv9en8VqFNnxMI1Ukx
mbe7CIWr9IinKhquPVlkjQhpHUJTSkcfdRSK1cXfXEx1Z8iYEliAgi27a4RV3EwirWRJzRAVr4jS
ClpIuVQ9CN5B7JxgfRpcOPSm9igdtJoldBROmAfSfGzCKZPQek626saL1lo4Oa1zDK5z+WlxidI3
zpgqK/e6MhNGe0ng3Y3Lr1xCvyoRasxmNn1Yl1S2j5czAFH0gkjln5mThUCFiz2rQ4lr3k2I4eI5
Vas0fD2Q0hLcycEbSYmhGyRQEM5zv8rbOMAKix7cCtU94cnELpEeMF855GF597ADyepXtOT/eGst
kitSHQOlc1vo/66rE46Qx9bEV/g2vYSwFPvEpluNky/LYYXfyZHvL30PkyWDKudR+ChGYpxXip+O
2UrJhJoF3jqfRwm+0kJXcYjPwQCAR7PcssDlD8zCgDGKSy2lvy4ggjPzlPJtHMLYBRrGzI3/196/
f3Y2rrs2ZpH/KE0cXLqA+Zgdw0V9s2XcVqatbTUWaUkMuwy5GwO959waaGPFH9FhN2pI82cNYy2l
wmtFbbzk38XRgGrGXkspbzzha5sNMV99JBJazsjFHyTuTbKkmTAVsBrRvwEN0sRBZHX5k6Vpqt/o
/UIGxkbLRQb1DYZsHJqBPwwCLyNe+l3qsrBTovzp9XAdjnhK27yCWUmP/18S5SAMAUf0sv1aqidE
fgZgDnHsu+7ZqviI/+3E+U50I/92VO64CB5oIeAS1BJ27w5Xz4bfwIHMgSmgNkaqDCuzPDBBqS1c
2nOrNNhIpnDtB77ZSUmL2u9W1VFBBM82UeuASPl437q77eGSaVIEkBSOcGRj1OBUKeI6ikqmADNS
Og5j9/6qquOjf8CBkbYIfw37MGKKVgM7cbEHp4uTfnHCkBE89ZN2tJW8W17LTmLe3K5JDPL31gPm
cVzeZD7O1HkXf3Qhad3oklZC77vAyIfUOrreRPT2zxqfBHOPpx45Fsyo9T5uwY5xURYbvGp1YtvC
pK7jRFK288RkFgRm03azS0eN/ZOYqQu46Rn7JuCnJZe7fssp2oiqS4oExUYALsk7V58WOZbKM+8W
a/e4S4j4f22Av67YmLjU0PPj83UlTrqICU4G5xbT6leeUdK55pIWuBMrctHn28CF9EG6tVy0jx6T
8La/GFhdIaR2K+PGvhszszX62/EaistkDIJ3O0NZK76vkOX705bIoFHBjpgbM17msn6rZFsH7NH3
8J/HNwlDG93Hcg10ElID+dgYpRfadIBdz3KTCfouQPCxltj6DZCD6tqBrWYxFmq6kCH6rqkwojq9
pTrGhmybL6wUznIjfKnm7zRPvVsPGLQEUXEy74klD9E0NGnUkfNX2L5YygoxikzPy8RKVHXx49E4
63vx7FpvL0kb0tZktujxKNvtNOD4P0iFFurTnx2c0dYRDvE0PuSk5YeUUfAzn/tDP6LZ4R6d1ddb
urSaAEWUJg+Gme7ddkQ2o8r9RiPDrVCbL0kEoW2LwT5SnI5GaukE8g317agYyQPEW591uee4Mo8U
L8a5bfQOdK01tJ9tSSRjdwTGxTEPBWSDLfW1RhTCKlZJajxmdp0cVhYbEjWhi0Tzm+fe/C7Ldq3O
1bZlI+FsFIHWIPiISNXCanRNNTRZdrt1UJvB+x8R0/AAiwjjXzWk9LLqeU29Po3axbg6H0uHD8w2
hdrG1B/6venuYF16PoKNoc275eSCdYWLC6jT26hFGAqtPRj0U4ZEKskLzlI2VTrMPoc7gFWKhhwl
+1qnXAaMHfBd3BBnZ5nAXwwhBqXrQdbTc0jkMzORsLPuBo7N3/54Wf97flA0mN+HOLdtue0bt8X3
ORY7h+ImumuQVdz6owjlNJI9O7dfmUhg0lpfM7USovlVxlWetH2Q2USNQVKga3wLrAokPsRBVQfY
I7jZHrvTW6LIeOzwJm3cmfeiRODdIoo6PFFHuS/EIClCfc3Lw9xf8GIGDlW39IIXw63RazSGeZPv
4q9rSZ6Wqx3FcZ0XAJpkgIXNybFO60J9OGmS3T7Bry9uYJjYV677OpKI6NInDQNC8yoqwGn3A/Te
3h0LOPbxTLWcrcLCJ59yxNOzelQnVHl1rPK+V0/iCa/Iidek3CZfJY858yMq571/y7X1dnBipy2E
MZny9CRn8n/LmmaL5Kk/gZPr2QxpGkBhT8U48EVZUpCVw0gbSGKWjx9VMCyR6DUXQYzJbgfbClhs
UYBbTHFlBKTFx266sjWnLaxXbX9n6/c8iePgpo+b8FDt1bdxyJwFjzC97HHYIGCZM3oydnND36rD
tNnAAvvP5K0ChVyxSUlDFDa5xCFxWUd+XkHsWNRURCljlmGoI7WgH4WW9Wl7+SufWabNn9Gsq9/A
KVvZY9bZDelYMZSxXCUmg9ffnXuJn6x0KSqXqrRQQvdgDBPsnUK9PBoOe9VzN7UzY2wlOG9dCruo
65tU6pnHKNzIE6puO6yOzJkLgV3UI7IEGj1DnOauqjFdVKU8d8d0sltXLNRvl2PIDZJ/3iJPgBVp
E17gH27FmVEvQgzSfjb78Pi/6pRgTs2srmsuO6x0I0Li0/HejfCCLtmwOZo9SO5SKsb0Sqi6P50A
66dNYT9KCKrkb14zRQ5cm17CKZV5bIJaO3KFOL2uccDtOQ4bvOS5USKUfo5IVeCgHSDue/rokzU2
m7SZTkcAq4iF7ePDegSlRj506IStyRewnTIpa6PWuluD0Abqcmtog7UFN74ZQezoavbewwoMxmIM
tGadoqwL+urHWc+x65CLSITbsA6r7wQ+6m3m0dDLmo+Px/lw3ZixY9CRbol+ql5gu8y8QBlXKWzJ
BwnvO+cY1SGEufotpEN0iPCA6fHizEHcikPtSx7O9281QSBSr3YP+mrhlC8O1IdLY7Ws4OeCcuM7
ZOq3zoqGE7Q0v4aFfS7/gLy/h+J1QDuGcE3pgAJ41toHfBtDFCpyGpe8nZtf/V/Gd96cV5cofiXN
PGSx1rR0uB5l86R4nU/dr5y4eBYRR6bqeAoRty+bROZ9L8nbcR/Osr0T//TPSIR8kyT1BMkuohW7
Itc+5QSj8q7bn9B12Lo+2t+3W4EAs1AZj5GveGXHn1Dvvn4W45aIicQFvLqjDUnNROFeZDX0wps3
OR+xwPs1ud1+xlLJ6Q8rSsDGtSeLRduJBHkBS6VHutG7dLh5bMaFtAR7cl1N42UJ27LVGRdqZSbu
Pzi00TAdbGaBcaexP7D27SyA5QfVuNI1J3QU8tkTzcC1Jq+fVwDYN8Z9ayCRFZ4nuheMsool+lPX
1l6pivX/EFZ6PZ25onxk8veOk8KDXUQAJMQyfTawYXIU4Q/n5f1isW7fj8g/JRCyJucjalHOReL2
tIykcqIlzgnxsmQLh6pJZHE5vWd7igshtSo/rRrLTnkgvJkYDtzxS2RsOKmQEuigZ4OhzRWjLwg2
6v91ARRrKuNfcybMi9qR8cEglxGsgGzTqcgBaGQNZbGeeFbSpLn7xrNZX2ArDovgpF9r75bXKUs0
G+NqAD867jabk4/RqtdHlUgnP5zGQWnfnnw3Hp5keOpr0Ch/rU15+/7HVmP7gs5NG9C8oryLyTvX
bm81auofIceJ9SQ4ocYnuxmbSKzni4+0vX5/ZJ7E+syPjq1M/FlJv0qqLUsUb0lHE9XY2CrXL/+X
91bEeL+m1IHALOeEUuMUNHYXBxxJWKhkC8H3tTo9FMgpdmFZFp/fzEkMw4A1Fx1DbDPExdcfFThf
eGMVLpZwgJXM7O4rUT2pJ5i1oNc7HKcdowd6SnKwfTfybXzeGL6YWMtY1aheuJlWcDiEVFxO2KV2
8b2f5AcCGjJOuIPq3kXduQAK9QEcF6gyf3EKxhyjnT+PawC56Q9F7UWlXZbZ692eTK9dDeOrhWEM
jZAq3evTGDfVGUAiA8/2h+jYsn6BXhgb09B28ooTvhEQdC2JB4JaRQv+eAiicZ6D6vpgwE4ZsRt8
z1hjbrakO6SNr/meHhqTpBhJAYZVHbnvOi3O+okZo/BKlVu2BEf1q9MNt7/nEDETHGERQssxgIeG
wZyWYFz7M8Fqi5XEowadHgILaCYmNB7j1fS2lpWeQnXhchEcOZvzeCUq2DgssFOC1o2PmF6NAeZd
+Vxl8gOCAQ1lEgHPoGxbk98BnN9JaJw4uD6xFXslNE3hMrD5TUU9t2LXb1vzM6zujyjm71fvhYqy
0zfE4BujL1a0+Q3tiGdJQ/L4TnGUCPYtuh6k6uciTfwmK1b/T8zK173mAbIDUG/WR7gboC3DGN8D
7RFBDT0o+SHWKf8X2LcCaidb4D1vsklERs9VK/djj08sdK5l6ePb5bT3B0sGrcM2e5Zfwi1dfkbB
Ww2mpFLGjxm7Id/O8Oqt45OIJtbArd3uQ4htCGSOr8uHyrnL+lz15LtNX+7XAgcmfGfBowf20zPa
GhMm+I+6SiUa7uoHLQlIQ4UjBlGoJPphZPkz/zwV9D+fdWhmBRbJ+rvtOlyBhS5DNPkDhVJ2/nLY
MqelJZlKytAzutqlIDpyg3jU0KsVIUUvTz474wqHQpPkyvwGm4Le0zYmVPgzqIz+SeJpMy32WwAD
RIGHDRJ6ZIzduEMt6YE+teeVzpGZMFhOWuES5qHxzkzlCYCgCupdV7YjRdLczAFzzPH+6EcPshHC
dRXaKMuJwRWr+gW/9iD5/JiL2bbQgEvVkdNO4whn590Rdl9N4MrjKVmQCHifBlgliP1b62xcpusN
L0gxNzsaSEqOjHNkU/+txC/SUhKXsnDDpZPyeXouX5o2VHCeW0n+yCU4LSxvHJ37TMqnfn1KQiDH
OyxNa6LHeEdFfI2w2hY/FHg+AKyWSGhHHRzZpxK5qpEG0rgaDYjHkq+S7WRqrVgWz00ecnuAoEeg
JWqM2deIVr3VEqM9Zq1GIKMUwtQb5GND4GybNKGISho3IIlFRNQTJB/901R/njCTwIHEjsX2vg2W
d90/2nTJ652+F+uvjK/x2ax0IeaDrMLXjSJB1ERNv8qppNUxSTaeC6DfwkAdr8zp5iJcDDfa0Jke
D8/xNTnyyj5TQW/g8VBe5mLprWZD33KTUpp0QbSeK6pGFIbokp3kpm9Ll1sFVPlJkezkv+RomZXg
DXSuVHQnOIAYn8Ad9PmHpKvAEaBcj5loz1FXpMEf5YKC3Rl979pSB2S8BaHEQmjb93iDXx/Dk0yG
ZRNs38/FvuJTyOCFITALdup6m2AKLNJoAPtTSG8jo1i+ccSgOwbvX+WW3iwHw9D9A/XATcNnTM4k
g6jguC9UrAtDo9GW78mrjBnCQ5dLNX1OwDmgYeIf8Es00rIIP67fpjF0JrunbjS43iUBTsITd51a
uobPuobZFVNpyxzvOs8FDGWW0DMBrMf/orSNnRUj5YdauXQkSUt502ou1LcNXI/7Moo8xvI3zN4r
525eZPm+dfxiaZwagrKZg5KWXu+J4O8HqmSMflo4QwrQJILFSplkBeTB//Vi0qwGqphLGo6W3FFQ
y+gmgS6vuq3gz3uxJSx4FgOX/TwJhqh21F3X72aJmohD/+j2F/AeJZDVu/wDnwk/BsBfAOLP9fWB
0bYcgEq5VgId0H2PIH2r4zVaef0eXGn6LM8N0qiItTZkiu8HwjBkXyNCfW8gqjlJipo9adSkckKQ
y8tflhZ+BPMdqXVySCEvj0pK3ZqmWdQDJNe2y9RQ0bLnWWaHR2NM+D5O74nVhjfD2+pLPPdOtn0u
QkXyCEX+ZpI96+BUoZvH1CyvPF0DZowcodULsLul9VmFCBRYWKLdA2GFlZFUVHaDgNc+UoHCEdhy
XytMKmVLrYh9cmUl66cKn4TufYHhCtNyYapnZPysD5pU/s9UDHDFBGl3SKfTRFh0RYhIZ8GC9Yhi
DmWB0wLrLkbvKxs3YWRaoCHzRdMUSC+e5EpnktKRWb1H3otw19sBedNcFYjHi26UBLqVhOFrFprO
rhEnGvNkT4MctmU/0/TL0Mq/hHDT4c+xE2Bw2Aa4a8pSLw4GO5XMS71S+zPvwbpuljJeIbSWn0in
M/N9ZUwALkW3nyNqJtNIz28EfuKtG1gntGLBTvIC5Dp8EvkbXfDkDxN0UlPenMYV4xVN5JYhmdlX
X6Yt35+U45KoG1kqNDt16SDvGUwZ3mUZeD3V8lSqr2UhgmzdS6d+Mo5WBEiFLgX/o3RqVVsuntIo
1+07peoYyfNWpMkxKvNGN/Q4/aimCL4Oa9+9qPQMmJ8OnnLqQnK3pf8Du9AWSFe0wnB0cG5n0AzW
PGJhX+DviW67zY0t4z/CX1PfnncVAlqXAOgfrNDHI+p7uAGa2OKqE4+XIeAdBsR/+lSBLsg6OZBc
U5gKI5BwmYVoqOVqvt9Oy7QseYvO6fdRodzCIyZ++UkAWda9svkVPbDJbGCDANy1TutJaV8w5pzD
GI9tNO1KrR4z9ZZPpXvKlQezwFvsmp8/xvFoOsJHuT86fN7R/cSvNjxHTWDSUib9AGCuFZOFgE0n
qWCpauiHQJwy5mF0pnhpKIu/taPA3bsd3m0JmWSstTLRpNRTfxcTmN7k0BljYXqBF8mAimrrbEfD
NKbinq8IJPsiLqYw/sF3/gQ2lspBIoP5JWO72UYCk2RyeoGQF96T43hoBmKs9xdrWF/Esz3WJuUE
67knBa+2btK1lBd7ZGuvDhC0nWNVe3gBYwz0PBWG0dOpUuIiiKOPJrzotBltHXB5mjdbmt1KWFdd
w0jE/JIMZ6PMw/JZ6c4VG7VRNch6IMpehMlZt7dMZn/5faOt31XAarEYddBZv9vYN7xnE7gqjFQk
BTjeLpFk4ZOWIuYc40ioDgAdXiIjbHEoQiPN1+qiaQLiHlH+PXxf6Qucr5U6CP3GuYptBFvlcMxj
ZwDEWSc3ak6X5H4dNluRSzdHEXFBytnBtJwqWX1cSkV9O86dvh+9EfPEv/MGYXY5yKjqhndI2E7Q
WGMvaQY5p/ILY+O2m585yfbth0qvp0B1EHbvHhm3kexuObIzRUMkcCb6OvJh30eumqhfQdFeLIa7
p0Vfr0c1RPf0G3WR9ceG5NPM5YNKQaURLmu7m8mbioLe1eIRQARcMawd7MtRtRa/E/7qNBJRxVV0
8DO0uYwkBtiiLD8RIf9/NLltOqWXPsAo3MZrUqOuSmRLJDbaGKZ0x79u/f/928clkV2QWKEa9qtS
wXsqOxuWmSSJoYMu0rPmEJH8UqS1ThhxbU4cm9o4RaFqXTkvVSdvBMBwwqsOiJwFlgbkvfNo7ogS
K1NbPgfk1ZbGhA3W2xFpLtmhGJAd3zh7oB15inKiPs0TyFUkNIQEW88y1/6MWLjyQZbnxL+wTBfG
/BOXFeceij+k4ww3Le1r6gOxhXuBiccNevoaMj2l9wTG/XagZiUdpUYwPwrVCrkcoRG+szN7l1ht
V/S+q8qyu+VS3tVNxokf9ZnYC+z8h4rZP9eG1HoKARbElcVX9OdPLVSjNXRKq/queg+x5ziNDLs3
fDCTynbdjGUI34UZZpgQfVK6zgSKLvXCzT7VX9DWGRuXxqMYsvpE08e7zKMbbhIOpvezugKCjauN
sOadg23AIx2s/Z9iDc733yL7TLcuK92Mrg+qafQSYE+zpCMvH91N01RIZBIX4GM5C7zdl+jq1e/h
vnLqQbuquax2T6eHjIN2qyMtaA77cxZHnjSJw0X4/hyuFYnlevgA7cXxaH5+y1LgD8OEeFW6HW6R
xKUVF8WO9PWuIKaNzph6FV2z+EFBzI/OmMkMqKa+vR5443isDxsttyXx08fz3w8SHofHvM8Pad+y
s/f11GGI+F/VFecgrDNav/iN8EvOxxntS+qtP3AWdziUocjmYbpZy2XB4T8/omzOBFWHFKW+/Wqc
zfsOZX69WpbLZJKDqAPIDaflw/IsVW2SWUWFreCRGhHlvS7tcs8GEaTUOQDiJ21xh0Am3+6DZLK3
cj/j4nwLD8rQePCDrnH2Etm15cubhMTlhe1mdlVsEh4DcVqSJCBIudPlQhBpCYQ3wHy3VB1JgHmn
KRdo3zI1w0ACn9kPkvXpeJAb3cUfu/ozaoKbiduU+NQKqRzm7iuloJ7RqdelbuV0EBHfcMMcvmRk
bzxHFJIXDarehvrpA1bOWrRTHJ6sU0N8etUjKCTwlpw/3s1mNLaFa6AuczMpAQEdA3XhMcGpnfY+
KIK3djF//Y97L+e54mpGL5y5zsCK+ppgFMbs0USu1IqjBcwS3Q6T6U43zjPysxtrXzQpj741MaPU
nvp/W6bCsru9Etp2BYnZle7ch3DhjGg9QRTt4KhfVgB/2MYDowsMw0TNPhNby5gJyIOY71s4epBp
knZN6xLEEVpkVj/z3UOFSMPUb+gQvC6PAeiQTi5cfF63SR61ygGMMAVmZ57AVWxLYCebXA+d7FmQ
NbPERxe11+Bt8DdB7+DskSPHi/ZNjvkmEG1Pqip3x9Zk90K8E9VI+VicRuMAUDuqKdwOAsJIO7MD
ogIqNctY4YE04QSlCw61xzvLnVLp2NT6d0mvOIu93StDb4g5/3J0npKMZfI2z3R3JjhHVGjJ77pk
xRCvftjSAvvRFJmLAXxuJxspWGlKMTWXeI0VBl+lz6ECm22DYiVwYzwewCs1s/RbC8GGa/8s4jy1
RqDItS0nzUDXEoxmMb1x+/Ii5VuuGhgW19UkDuGC6RIesIgAVj0wufikTpFlevNUc+8NNXkDf8QC
EZ4K/VSurO3plwhwD2Urk+SsOnNuk5BmBfUGIS8YAAZYsMzKVSqGqyKbJJl98yDj+k2ARDMH9JRQ
0VM+ZMA/6siL1/7Jqi9fNMFLdgoQjGDXX98zhtVuXn5hJ7YfOmEz2xBYnXTv8g2rls9aZJcOxifQ
t5JemVhJXusxa3jtgtZRDG8TxyKl7VDu7PHrfD3eLgKQkj4vZyvrgJ+XolojeKPzNTRQusJXo4K0
SvihnbZPqAz3DTfNz+iyokR8E0CylQq07X55fs4IrvKaKYj1JYKTDAGsmEAa0O/20Fqoq61Jrzj3
i8rL2xGmxuMTc+8rr+68o1YwSCyVMSL2qBJ7GdEWLBa4SWEGljXL5ZzSKEmU0rjXgOkproLnQ+MC
xHpQFJo8B/h39Jq1DjzGlPXNnufIX6LCF/yVn2hdwiIlEed7Fktl8Iwe38qrzvlH7PKRYqqoo4x5
khAXgmqkAr2F8d+utYxY352Aqim34+5zlsipmHef6ru1s7irjcTq6gp1pTJAA9TpqOv0ftkwlxEe
fsQtX+Y+7ZhVv2NhWIdoYNQ5gPB0yJoSpbqIRG+NLic/IDAyUipzz+zakbuJgH3pMIGXaRUxXwAg
sAWcJeFVUkBVYQzwTm3ndiRJ57SrzNMEjbEx/L3QAImUENx2X4hHpYG02t5x46S3XSPzWQ8kYLjZ
E0qUpBsKiqt59U/sKKj3gvCVSoZ8TrAFnrKzJ5529PVIRXYVIg5EDictGgZTDqKK1Q1ZsSruQra9
OeK2BtW56LT3hqQXKhuiWEuW58s0z+o4Hj36cQhX2Z6F9wY8b43uef/azmvEyYY5WBjwMVGu/GF+
DSpDJyCk7jnDLuIvnOXuOsblyt2ALblb6mxhbtlWCoAl95Ipf+xAR3OT7KbGpqHHCl4gSqwn2pFX
hSoNRiuWso5nGjPm/RiOq2+2VCVCtvIbCzfOkgHyKTvNxbtHyog4y42HIYHLG+9fgUMxbz7rNacV
uoIcHRD4kXQsQ/V4WPGCvPygaB302DYEWqUF/P3X+ZpeEMcxgzfgajQ902mXeI/dedq9H/I78u0o
wV40SeTbXrwPuAk8lROf1YMyFPfv3Xzt0qNqTeFJbo9Kq+EGdlzUQRmqrxgA6F/WVgMg7KN9nmDG
tbfG0amSE8FUEFDycKer/r9v9ZgekMvhr8SZ1s+x6GBZ9FgoiEApF+WtYm4VHbw8GcxBpBmgIJna
M1paInWwlh7r8Z8GcHJcuNdo5fWNzX4fGrN+GpXkNRkrTNPuLEs915S1oTsS5/cYMSSG0lDRWnfh
W7mdPxeJNuym1nGSBHh9qiuL3kToUwhNIq3k5L+oUIPUYkQjiMyp7u9yN+5HVdY82HYDXyNPF5/1
aUm8BWZBoOKb0ztlLiiWQUvxOx5DqoMGRfDmgdThs38dfrOqrJbfe0uz6duYPRa1IQNwgIr/ig6y
y2IKtspnNIziqmMKBhr393mjNxuBxbF6QvDfESjnSjyB4as46o714msHs1JSLbf/AuhbtzRgB8SA
r2h/0bq4pf8WhNs7Ma9A4vP/XnWh1AYFJXneFR9/wP+Dd1kwxxb+WlbVtvRHYgr5K1c5/YXNXHY0
UmEMdgEMzMbeRNLG9qRxITVeuRnmH74DsgQc4Iu3dDUtsupAUawwypyAF8DhyuvSonLvvou1NuMp
SwLFh9Oom9LjOthX788bDFzRa/S9TlDskmQPRFho9/Bzv3zTbWnYXJ6T3WjrJLFHRGi0kSTbGi1s
xyKcsbe+owry0W9IQWxP4K9/Fknuj2kOD1fcQxFYJ195SYCKt8hFzsAfTJkwzN89kCNZX/Ct2x1T
Hm+FS+/gQZTNtuznTkAosD9iLz/6XxuJEc9PpOUpVEJEOLaDlDlXgOLI5y7MrsroKp45P1u8vZQD
IvhXtt/40nU2qiwkcS/F6udQ9e/WqGs3Sx9C8TpqbKERTjv0Cz9RZ0yQK6m66Amr4D3ad3jhd2u+
9HvUMfqPtt6Mgcp5JBf5yvQW8V83AN1lG8MH0jH8iokpczuy3eVd+s0qGMuVjlEoLq4pWIzb0N4k
gZS+x3vWVPyTluFSWuPl4i27TIw923sJmp4LHjDG2AXiz6rKSh0PJwuEllwyErnQf3utzn5Fb9Q2
7YcnTemPtQt2QYJA/sn9rPAhc6g69za86bLdCcQWc+5cqpi3NQvRNN6NTXM1ecVVkdbAm1xRIuTp
GeWckbsT8nmAyQLngei+JWW60Beo1Af+J8KlTo99puXVhUupPbaTjE/Y7SX4Ei4z105TAWLwGxyW
VoIlSK2DRrk1gEJYehQmDuBUcMZQifMfvXLPvhIquBf03PoBkKxCkKYdU7o2SuY/cnQbZO18ZYdy
KxcLFsMQeFPrLPa1+L6S6bJS0L/9+qU2AI4b1Dx7GEnA13NgpZIAkeGrc9UQrJXakFGhDgx0gDPR
7uxW+uJIPJlFBIxxCfm1iWVNm31RAOGJx0Z3DSIo++u2u0mJrwsILA7ZSoisSwO2vRdpwj+28h7E
ZVQ2d3QGVdq4KMeuritJ535aLNcgx4CJch/zUHr/r1ck+pngpPgYN+2iewRfzier5HBwoYDfribo
it/+uxZiVl4WnbZZqvERV2ukq1Hf4cQ8FBy4ylkZy3RLM4UDYui2Y1hw07ajHmGIdT3Z9mih6GSY
lwfaq8nHErz4O/7WuNwfwovz2RAKRAm6s+5o08gVmmmX9HSMAwq6MGMAIjIhcMAOChuIMlKXimp8
b887Bb9ngiAWLkGo77nACxEUolDcxozSewYXPRap3jVDPRqtZNJPlkOaXudrk/3SNYbrQpkSPRNp
sJOtXXbT2ri/546ca9Rik3Kbe9qJHUz3kGxme88i/zwCotu9gn5VMWgHNUdLb2fPaBU38Rskx3g+
jYhAXcCGMA7EJoaEHn8Oa1hgweolAs+x7aDroZX0tiK8FDQ28B1ShpIVAdHg0oGfWemlFeDsYvUR
rYHgericegjJAR0q0z1tTTDT0WbfUAKcioqjvTVF0IsoT8bWkla5C+3VbyiLTCbiPCRe1JZyPGG4
qKTZ5ZaR3re2t+lxLK9xfXve8jSySL/k2guna5ud1etfimmoH1pgzeBqtIVErWGnvIXMLM+zp39s
j0lAwHbIrEz2j2dIyxGqslPPrm8iLE2LbTTd04aq7aHjkXrp5ARMfWoYLrOYnEGRAw58FWbS9I6d
j6/8jmXzdwmiGDR14ghxc2o9pYMPwLZZHKVr8xD+Fcr56oaFgfPMwwzStzkpgnqjlHeL8FdJvNI4
aSbvn+f39MexSFmNqnS3yYOEW2w6387hJHGTFFY6P+ikcblbRNmLfs/jRW4xC6IXHcjZl1x9DCvY
y/CZUdqnidjhMo4fmb4BTMqATnWIGTAp6JdnA68QkdIFUbkqKGbE4yH1xZSsWK3swHMguwdyEHVR
FsGBHknbGQ5954MM0Ycpz6bw1ZQHh0hySeSSanCr9G9YdAFw4Kn3A18tcv/DY+e0lOt2H+wOJlC/
XsNs5tnUHOREJ9Ba0kGKzc6Azji2sOKjiW7E6oT1+ixCauFsA4RSbwLtmASg+VZybECwFPewF/FK
v69BgR4WdbFLcqEhlo9GE+CV55C8BqNq2mVE4n6lFHJfvNyOJXKDl8UrI/QkveqHR1ZPmNWjsffn
d2B5ikcTYacs6ZE4bYaObOcGBqZolstq3WCiFaReDmpAQ9kyP7dSsGCsTwCqBK0Cxkwt3pY215WU
i1ohv4Yq2M3NlcIWrhd4Cw57a7m3ugfLDdfDlD1UfghMH34iJFDlIdpZWHqlhzADdUIXdh82U3XY
jYitnUUbREspEhMB58+JX8/c+LuE947HYyqnDKVH0aDjbC0DCvzTtDJrHDJYXWdRpdNB7YXb0Ihp
uYFIkZlagZQpj0Ep2y1GbAdLWro/slqTD4xye0XokD/xcoLIQEYsaGzj+lFx7HOw7EWH0n9ZeCRV
/Ma5SFG45KpkZ3vGHCUBnqNRC4JuyMZcFrrzbJSceJdCQMoWTgGt8F7aVrr620s6vModCNbvI85N
yRhbKQpkNenCfgSMk/9uUgjxSe61wPe9XDA3x7nNHbyCMTTcvt7vd4IiSkDuxIUtOQ4YKG62BmxB
CWGnyfpcU+ZtAT67YGdwzveLvvSzYzU4tKVp61TdT2DSPYn6yo4RjzqTOC6NQrgOLHqqvF5CrOBb
+e6Sv1fE7EgeouIGe7Ah8mJqra3vuoHdf8zPYxsrX8SRHwiCpKhwCt0WetmvnUFAEtaqi6u3dkIL
TCm3OKb5sDL+Vo1C/pgoIoYtvRv66UR/BqBNAyTH1Ep2b39cA9JHTKTMjKVkKuLynkgYqchoAuCF
Tptz2Uc3yjdMOgw1kmUtMuf9VXcv78TSL9z9u8nxKrnii3BSwwZpee039bjTHDPcqzhDSLKWQlnz
b4a1ZJl3uJUmFA9ZebGkp7xpZLa5fJKu63G4p1Kef3BWCZi13E/XpzF2HX63h0zrlRumT18f9rmY
ilrWng3kKQ+VY7ksvTwiIhaORH1S8jPyFSjI32I4Cir8r16fPf6Q4hcAh88aqGnyC+cbgznqL3bf
8uMlRFH8QQ9QWqXkfEPZu2ECbomBCwZ5hj5l1iBF7v4u94ay05m137i9Ejk84IRO0sgD5rk/8/bh
UIVmEupmS5CTp4U/fegNOc8uNpqIN4CesgS7y9c9/lNg26zF68FUFHghn5Au8qGo3oxLN1NcP5fw
dx+SWA3269E2KmriP8pl0KEnqqM6M/AeFd4enTg42O5pTpgH4TYaD2BB8KrwGiKszR8ZRsGRK4NE
t9A/u+tk5PgWywq6SAUSnhpeWG/1h69nQZ9Joi4CKcKeX0qRg19iX3lN+XYwg4wEJfMu+ByXE54Z
I2pyf6kUE4LCAtvYr+Nu0sloGNla01fRm3vHnPs76c7DWASITgc9fBMeQAD4vIABbAUaDSrx4le0
qkyinGgwjedVzIKyLWaz7eQlSP5bXBOh6okDPZdOMAXeUxQsyAt0dNxmmq8Lbnf5N7ABiJS1nEJr
r7Jtld74fsj4P2zhjMhlEm6vabUOVpCgXF5aHkzJ9E8YSKUAjgRwYkcscpx5VlwLVNRIVFtjttJH
34/Qe3o5AQDCuct2Q5Y6JDdC6A+f/03gFVAN5IYTYjDGgcSByH7U/oYhrzAe94LIu9j6txrAe7x2
VtQ0HYh1gBYvG80JUj3hxENZdhqnKzOSUWbQEVEPHj6t9TXYLHGN7CiZXTK9zZgbNu2DwaKI1+eo
mYLfxP3Dm2fBEfn+4/rsCtqBvRYuxx6asW2myx+yPm55jFf0aX6Uj0JuAhh7WERcNvSdtfBDiKdo
3hqkuqlg5q3Lg6HrbUSgq4VrX1aKgMELRxFAcb4vr4W2FZCeNv0/82tx5NgCcuqpNwtcffHT+ZtH
/MEYJyJzus+ceTqP40e+E7auNxePT6uIRiOQz7nF7fc7eAhXOxgYDA9ERLMox4UrgAJeAioX+2Yu
V+02X7QzwTDvmP1D3mVqdupRQCnxpLTbhM+IZ+CNt+roA8BCEPGtZe8cKQOhh9l3nCvLb732/ZP+
F5CuDd+x6q1J4W1RJH25uTp8bqNX8DCtBilb09pC4A1w4Zpe0ASzSoDbv850oVjBiY8JR5kMXDd5
lkAGKjU8swDnfqaVDY5p7NNG8L+PhJxVaVq6KEQ8B9RGFURohkX2i/iVMyH8isx/GiE3UaFZvUJu
/UXnXyNmwiNDulTuOpjP2oL/dQQtU5ZGnl6GRoxBw9SFdmg7Aov1XuP/eB9eIAWwTJMj7/H0ASwa
cwF3/nDMozHOtJL8VaDxhQBL8/ynRcMXsGHQfM28C5Jbz+PeQsbjBSlpnlLbxgxRYeB8I7Brah/x
yynybPGcBxU6ss5L8qE9tEaoZjHBgq0xx59ivRrskGDN/7PfQSk4qZeOAqz8IpIgcapL/FJtpJBe
HYCxauOBzRLv76p8OsjaLIJJU6o6jWmb3Lo6xDfSahCnlRgkSUZLp8QI9UcPoalghKLD3Zwsix1p
NmPDqVQj/CeW3ah14Vju+vIOgrMya/dUK57OaSiUyrZalB8wOUcygsYiBxEsJ6C5CRF1Gy+Q2GBI
z5i7FyofCDSz5WRVciABIMrTL3VDoNlNy9qTuMgRNWK8AwyoBpjBzrHAtYERKD75b1xtwKAqAYh0
5f4T3ebq4QHHFznkhyFJwImh4ZJEEapDmqopjCyUN61KCuXR5Cg5Pg3txDndlpoQzSVnxFU7V/I7
gaP1qYsXy/FkXghNgXin1Gy8V7afjigoUcijyMgXuU1Cfem9sZsbUCy5NTCtO0en3XNLyy/iCxMx
243n/VoGK3ERK6NDlOBpGQs9pRUkBgUyigsCxT3/CdWAyCW0DddWYJlGYGGL0ek+g2SaG/AUAjmx
pflmwBGmCtFMjA3ibsu/dtN9cbD/2XNlMM5J6JZdaTlmuqPu93FzjaJH/eDJrZTudy1qUY4kQAZh
lLodMgqjqjoMrsoDUi1uyOJG48UVuDQTp6semsX9XZ+hifgl2F6dyZnjVeBjbegDfh7RAzjYf/wM
clYhEw7+u2EAbz4iCDf1fs/EbuZQNo9+6MZI5OA50/PCGOLp+3Y4+n15jv4cdi/p/q/eShwlaltB
XncwZrUxNIpMvUtCjaP/FxlGw8V7Dx0VGf5ftk13o0vPBquNLCjpkA4+hQShz65VtK5RThFdkaJT
X9BPBLPliI/3Jh/gR+ahVSS3Q8ZuH5k5h4r778tgxnH0MYEPO8Z/faYgz5WRm5Ha38u2C1yUgVw9
McM575XG6CiJxIPmEWNp8w+FrFLCiCUR5NfNaAa3TOT0SQsIvhVFpD5Sga8Ydenyhvp47pXP6ANx
546TMsXiQeqL0GSJXFUHHA0uIdyDKg5JlDi9+GtPtkPsNahSR8ngdLo5NyP6cifjuYmnT8GN69km
4vPLz2/LrL5mMUhjP3mBL9YtWID3UPFbjULldNf1SkqeDVpvkZEjrzplC5/YzJyP6Jmzbu0Z3iZn
W/f0WJdJ7F+66HayK2IibbowA7gSgtYL/VpJTzRd6FA1syG/7GTo6vDY5JPMAf/h/Oz8IonDqEAI
+6nWW8MfkKCgKOI3M6y5xFpGP6yoiKUn0cJu9zDEk9qMUEX4s5/t1HlpmKgsd1thRVjMyRoaUurG
6wnQzlfNRsRF+1e4oE+Ium4UXGH/mRW7tf2c+KiLPcUuEC584MOAeVGBdDatkBQNPeXsOJWsQq1L
Pio8EKbOsXPrm43J9StcOjGMM1pAYJmPQsIoVzIqdsEluS5T8m8tA3CMdWMuXCNJ8ly0XbaeY4gH
9srmRZt1NNRoot97vGBJI1ByVVFZCU1gbax82ctd/DM7OF7OMgJaQq8V8gVcOhjDfEaslJ1TzDGK
YSNuAASWaDAEFliQ0VM+670BjM4G2ei1zyK+JXYsLIKsNB8Z7QnABVI/4ksRwP+Vo8lTJlxpeG0A
oRrKprs5ie1ec6akCPM7GXfSV3t0hu9U32NRJfXqKLM2DVrzDFaSiYJ1SSYhcdxay6QIw/AUkjUf
/0F1tbW3CAKHHrwUd0e2zMVLtRthdkFjHMTNoYMzE5xsG9ddE5WX32uqmUSZORoJgW1ksdKn60BJ
c6Iz0LlzGUxekcbMJxsS5Zndc+uYitxYu8xvnl2pNk60SXLLT57Q0rXQFnR/LFe30ZGUEyC8MQXl
8kbxA/n/W39qmN1espRMgbMP5nhx5BjVa7y3pvxBeaaFAeGcu/xL+nkcUYMa9ky+wo138HFuPhVC
VJbjki6mnMBagbpDc4jrTcG8aGITgC3pOBjTSUCgCEY6coran0QWLFGtxrQ7WGADrOQmOMFmNcXh
TnKFYtBAO8VtKRR9sDGW+PWZSwIo19yNo5nzPMrWSlNEzPHzKpnYikgazd2t918TPywsZhxEU2ji
bgT7x2h4BItO97JKAcTYVU+YZmGw9+WPDExzHP0JNW8IbueOlniv+++axFAw1/BCybzorUpdUro3
zBtquKzI1V8SGQavVq1TKB7qq1Z8t3YgFpzCsrAwe116YSuBTeQKLIjqj4D+vGuPHeKGoWYbW2zF
+17TFB9QDTKZ0PntobyF+GEddrJ0ezfCKQN8nc+i1wukjXeq/lEwH/t3SkArZeAiGFSAB4+RZgOk
OIqwpLmCGhzX00z7WbGlHGf4sOm/wy6QVNbtg3ttjN24N4Bwz9NNkPJ0NNzB4nLfu122u00gfd4f
2LdIvtchS/xtBir7dQaaa+zgTI+e3UzeLYWrgw/0SizNYFE4xfSIDRROMslxubhPJVl6FrhKHOC1
luszxHUiExa909316X6pzvGTI3rKzAlWR9BEUWsuEGEl3rEZYxnN41yAxMtjw2VvwcvpjKOWyXvX
18x+wJ0FZsxsF2cvjGyAGnq0RRvqFNRmFAyu+I7jwSbgRFv/KFH85xKbfNLIvZDK3HfmPEeJv21B
YxFjo1aw3h8l/jkZmAyeF+dXqW9WBke9VyBlmez6lWA8d6c8nsBhPjt3cmCWZsI1YfItmP4KfsQC
4aI7zDAdsibmKC/0aqAI2D86FnfCusqdS9cRYhaeO4QPfoeTKFaWEMnn96d6jJHPo+f6RiGlLjmn
HDn3U1769FHOgPRHo+jsbbsSJrYhZaWESJnCvtsNUjdtqgV4fMhlkMB5DOIaTSKdH7sI6Ndpi1Cv
otT0wx6at1cXFI+5DMvFQjKD2JRPldhuamgC+pW4IgdlGPwKSANGSprinCyszPI2fvXhwVN7CgWC
1RJ9MxAp6uX4zN+m2PP/ae/Q+tveqWow4JGXnDeB4sOTn64Byjj5Esc04z75qFSCaOFy3gQPR3k+
dZAg2J8U9YYHQNa1/LWDc3kVMPeRtXXIQXDhbq7EWTcEtZXnP8hE4F3cUpi4LS3qfm6/IiHqARDk
sGsvRiIU3KYCA8cIJZHP8DyluPNkGdAkPqJD4N+NGtwsVF4keC22BgVn/ywZ00P+Ggr5KpAhGo1U
J0iLvpcWkpIBf3aSUKwfYbnt6O2VW5B8wCANvqEeUELPdhs5U043bsEEV8K1A/Gi2xIysUoSxgKQ
ZwBoscqVa9eoV4hR7sY+56w2pLcflWvH06erTDbkbe+TkFEqfGX6gc/PcFWIFZ7F0YjfDU6OV78G
5dHuXNP13wv9ZSdqoh0uRnSv0ds2HQ6aqouHKHSMv3i/zzpVvu2/mi3gzIMdWsvkd+a3Nc6lbi0D
aIOcs/nW6YK8BwttVj/wjTb1PXVPswY0Qb6aUQPLgvL1/BmJGZBZuKLVFkJTkld9qF6zsrAtDCZg
96y6Lod4lBHCH+G09O2aK4PJ4sOjQsQoqfzfODcfEjoDGj/0pe13wBAHFc6rfFZWjocYmQyYVYgf
g+3gPufAXIpupbdZdwPMg4uFctD4kQguXDlCJfkfPraWNX3v3dJoaw6cGQPBcRWVgVedSwLqpbEc
fjN4pRrwZRIj/So1sB+fhPQip0afsEtXhJZoot/ZPHDb2OeR2gZ9ugKEi4eO3X4f6YTexMVjVgMm
KPCYio5WR7wnk2BHU1vygMiSM9vutOtepKPiRB2O7YCAlFZWassqW5iMNHs0Y0EbOurwM0bx+gcG
xDpTmfgt5h3HeCYKreLs608QLxWQgvSzK3/htZcM8+Evo64HEN3fpY/6edwNOJgF8p1FsY97lYAV
cvYHIJe3m5VZ+JzfGNh5acnYR/YwDpa0d46x46ufyn7ytRILhRN8/XCrZwCmjMdVDp2q2Epe/6BI
QsOwzWRCrjvzn5yOsXTxj/BkhFe02SINW5/KzWIjYWDNBjyKuZRXJ00V6TDAmJ79PZkI2f2R3Q5t
QN20EIc3dg2FMqusM5cQNN0cYX3K58MU4EEtUkQ4e3/eQzvmvadDmmpL/yAt3jW6twqJzqj8mDpD
8T1rvWW/Uc8JyAdYJtFdYxKKtjuuJb/fu9YA+YKMWb1j65PqwBO7/rsesW1O892YMiIEfjg2vGyP
lwTvH2dtrtOnmqy1Gl05ZLVGpxjeh/7s5sJ63ZQe2hQko//A/2mVEUZc/Dy1ChU/82Afo07Tpa4n
Avyhu/wlvPsp0yFIRgfv/aBQGzgzF4FkJWef+LDR/fZkDz/Vt8H23RjuWGbcDuobuFHjsUqbp6Mm
X4cnWcMI9uN3kg73VgqA22Zh1ZtPejDtQbQB0iArSUexB2+R40HiNl2ippiiYTxKkeBYm3IfyIAP
7w86LCMyX7Oc+PC8pDz7BBoEccNqns7KjuYnOoHU0DJN+3yIUR0z57+jtSAVD2XWDpw+US5aUI4S
jOo/rrlA2+/uOcreC3zUQjZSOh0MIxKTJ3Rqrs4NoFsBX/u8DhYNfm+8H3rP6DhP5H8Fa27F9ic8
CPIgGmcccYSffgkHrDsuM9z1iOwZs3sXwKGjena33UcuezWKql4QIBTdvTF8DXiUK0WxnGOOYIFT
ujwnqn2Ob2tY/9iOcoQFnv24S+QSjCnYnAidmCIMsQt0K3kLoPah7rG0TaoQgxHtx5VpAcuF+rcP
ELqZZe52AhbBAxDBBAkUGtmN95pbYP3UogHIjFxiXUZ8xt+6vlxSszP6rGbjAblrzFgJL2ttzd2M
KwMW9f7aFwQ9D8oc9shJ2Fmv73SZMZROwjXpMsshxDff7FlPAidtb0CNtL1xp6GoKhrMHY+/bZwv
Sbm9WBVsPClawFQnSAz7Rv+cQ4ut1ciEbgoPUkOFKFGlIm1YWUjlc8hR0xNYcqZ+fVhg3h5MKM8+
LDAV1Lh1bOENxiBWzU2i3bIOSp0J4wEJpo8UAt0mzl5xbRtFgak4zr9Nxa95jlZ6LqZZXMlckzAU
hYoauTKwYCdItqfVXbHeI/9oUd4wyO8rcfQJ2etDF+a66LQYGhbWLtFJ4tP4jRZS41GYOtQlZy9O
NM0qowrEOylWMqdv3kez6abrdq5lNMUcJJmeZ6OOZIK/gxo0QgcopS6SFfbQNJEMsG47GWNPEcW2
GlAhMkcFlQ5A7HQA/TdF6AjTeIy6MO2bAWMhK9vAPI6Oxl53aPi5qgmG2RH/bk90VnBJttUU5hpO
7tjhieT1s13M/BWZLxtWrgnKlWNDPI/Vji/7R8NovH+IdOLbYfa2A2f6Bs02XVgE6TBbGZ6OiwcJ
67qH5vQ3HuA5Avsgi93Nr1BYwwdFKFZ4qqBZ3o7ziVuNqcFLRyPsmDOdQQWwRdjHgP4kdrYqNk+Y
OYyvb2f5Nuk1cgyGZxGIlB6BwIeDrUPcMKNFxiq78X4LSgZWuvazGvDNohj8amdWVt9xH6zzED5h
7KsVu6CfnIU29UhIgF4qlGlcI+OP68vmTzK0fiFqVFYrNfL3BYkdonel16SbwDwhrojvnHJOO5ET
satB4INouuMqHSy5H1hJT7UekT0Lidl+qUPx1dyKc6+Ib91Qt1jgTAR+Yx+xzfQJamZlGHHk+A32
vycjbROBfo6SguQ/t7xsnH3VXJnAyCNJbdMpAbzB9aPSVRtuMT7NXFjkpZ8rlt5BzhPrJxdsFBDl
uNX+q04N/xQFS5IGQNIxvX76Hkn8066+XnKBhDje2EUqwOAi7sTuFtdYrvggV2fPrh5yUSuao9F7
NKvIHlA1JGAL/i3rbt3QM4Cnpvu7m0eSC5rJj4YTf37fXisF/ZTYtJb/WdOYgxwuJ/F8yT0DxQxx
vVSdFZ3Rbbud1af0SdbPGmtNiCik5IvT/gbhxOMhRBhzFN4VA+He2JnLW/gOb9X0nUQdus/GFMBV
bEBU9Kl+4bkpgR6QUc2fdoMzv/gKOHImt4VoJO//wQJfBrm9BNNYf5tgdT+Nq1WYax631wuN1UO8
Adux3yQDbHbzE7xLBA3pMiw4kzHTeqkqbHAgxLMZRSsUnfS44kRTfIZacnGUtJ4gHP6aVQaSI419
O58HJPKybyeDdDds1AaOzRA4mzWlSMknsWNgouOH5Pqyl4YOr/OTV9uiuMp2uz4YL6BNZw2L0Tth
bSEhGcsVi2tM3vENWZc9eKWVFacNG9KuMJLPJzbflOqgGUJtZ23SzwEwawKXlG4nM7cTeV0VEHZc
g9wibkP0TUvfr0ryK3jmHN9G6rms8zzlEIaFe+5OOBYwzytvBPwqvJyx6JTEICGz4drXEP5ZsAv0
yl4zR12SkG64UakvEWQEp+vpfWdZB1tuSQO6GS8iVtf5x42AAntKj7ytqcuRwYr3H8SvviPpTfpV
YlqAmyi/7dVBsTDtziITXCoWsZ+FCvhPQWy5uy2mYkAEZT48bzC2wLqKKONJ1+WgEeZp7PA0uMCk
W2970o3gVKy4aRrW6dM6iAJ4fc0a8nWLPM9Uk5EzE4kJSEG2hGiJTtz9NRvkY8va6RElAiLSCQlK
b2LoXoO9IuW6vQyRTxNFW/XfkmlY9Pv3t4cTDWAwR+DaD/iWPjISVnqSNDI8UMtukT4Jlhl6ipVW
kG2GOe/ece4HSJKUDQq2dsTjnd48lBTgmgdjfpUod21EN/ULR42saDOzh4kv2NQQU2kNbNPBK1cV
3zjnSgFwd/DxG+AgPIPdHqsFl/s0b2VIFEskDvy9ccCbcRJCeXRnRHPlFU0C+8yWl3X+cdP7DHCB
4smJuo7D2jXSR3G7yYd7sbIIdeU+Homw22yFyF4CPhWEeJg79lb+I2i9mrSSwohb1KJ3ukeGhR5s
0/CUGnWsRpyNrHrJv+BIOTFzE1Rgz3J2zNYL4IZ1RChx6xkg51p3BqF9B4eGjwjOfyLKV8GVBYlT
aqwRYkA+mBJGjNRMArWuJYfiEv9uPmtBCPWNpw36BQkY/h6Wg0kICr/5x6kJShuK2MP9LVDHwFX9
EUdpu7Skt6J9M7sH9RZD6z2SJf5MS+IvX/vR5GAdkVwNdJorIHzHQMfdjLuOmG+rELiyILr91yVm
gqHvEaobnnZW8aRNWRFAa67low6GysxJuhH6R5TDdlC+LvDSAGexmmmn/r5eckVnYqVWv+5lj7tx
Ozbhs0k5BReV/kH+iu3ZWREga+QUFC0iKUw6F8bPPVsGfOePQJ/N0t/NrFq0xNIhFTZS6/h9w0tB
+r/ZpbWhNXsKFiQeIcGJZ7yZ8VmhAoUGFtrH1IaWFrSY4H9i5hH+zp65QuPlfXkTVZbh3IoDTWQz
z6C3O3O2+4MHgzFksHkoIwlxBII10MBIRzLtoSISPSEx55AqY+sdycvkUkmmKGWJ1MwYIxkehFgL
dk2GmPPlOJaQFJi0gkl5srFhzHgS5Om585FZjeEowomq0GCa99+L0u1h91ZSalAAESzhJM5/LTpy
0+PmaYJ63l1rInVSJ3CPE3YHEDiQFQyzPLXb2w7dP8iZ+kssXk1Ai8OzQMsTth9t3EdcXfsOSXIB
V4zxjCD3P3RPzYDz5nnJbHL4W9S/WF5k5XlwoyTFR46OjVfF8XxKlu0459ZrziIy41dWI8QWk04z
dewJZ5IUAfuYpjIAdTm/q9qpsAsu1sXFUwx91hCKZBN5V6BwV8M3knkczzey6gwC6z2IruPneIFX
JpwrMua3AZGxXmXjKCAmp1WS5dWKBlSEAfB+I0wiCL/P4psXVi43mGEsT/SssGp6Mf0IbCiX35Ju
KeW8Mawq+OYIFgUVohQraPp+ExfvcVifdiI36UULzKVs7PUjzpqAFGylnV+LRQHTS7WgXVDh1zAC
YA08EhWvFfyWYTCwBNBJuO3CcrNLtZINQaIZD4W1bgbcNNicEKhA3LiD+UrApt2XNvc/qW9jDt/W
iS255bOWWZGOqQU9scZAPbtQ3xrS6l9OufDeL8GwLPo1uyR27IUPA4EnCMR7Ic0QhTdha7t3xwiW
f08SFyZd7JUjNtDPGn8nda1sRgYCiRCNBhx4uEgFoVdzmcQGMz9gSgEI/OFmJtmeWXcMEjK6ff/i
bQPyt438vJzEaK9vbL1zp6bf8lRKhp150XFP95mYVT62Kz4zc6ZMxXRe2om8X1wEW+DgUkWsiyWG
GbBGZRlrtrrDeJUeLOQcDgoozC9sE1jqap4R80Y5Grw9ceYeeb4Whq4Qwna0uj2sBxYIF7ecaj+R
Q1ZcbdBds1D+xPA7fd5kaviIbBxcNEsEAkZzKKmZ0JT3Y8e3mHu76bR9y1Lab+jxFOLNCc5Xw56V
T2j/mF5e/niEOZSsJfGCf1H9pDjyWjeIlS8iWnZjOQ3cidbcEhGtE2XMl9qv9aA8nQzqyohBstfN
nmctxsfkUig8D0ELe7J48BhyFwZQRgGUkgO/SExq47DHhGoB+fM11aDzUyRkXGwd+BQY2osDpr23
Qs5LjTyrf8WUcV1vlJa6W76e4x2qvJOv6sM2OXN+Q/gQg20DcFB+/sTUWh34poEcnM9P+p7+XjKD
ybYSZ3V51fd6jIsCQXa+S2AB63BexmzCJAjRaIjY7gatbzM5g9s6OYMZuYt/6Tb+NudoLinVaTHo
F49Nz3HbLfVDUMuYsNoIk3QWYKMEAl14ykMdfSr71J9VK8240Iwh6fvKndRWndKbMstygm8NSoLS
OiWHaEPHG10ZXwttgaphuNH0RB9ZwD1urCvERiOmdeK7VvcO2g8/6zd3zsu1IYE6LVNW2xXAyUto
rSg9vdSr4XdIOHI9CD6aixakr694i+Y1yZpyPFNftsDY8B5+3geAn+t5Xt3oetdJdhlluqB9kHI2
um513BSmA8hAF3wYebU0MDw0WrQCAyyLjUxm6dgwI3Sme1vjT+KGSyYwCLeKuacke5h+2qOsK3Hv
tw0dEMG5yxJW/XQf9naiv8JzDjhIvLHoWLO6epCQzoITGlivXW4CNb6WOSDHsG845vEDfK3H9PTI
GkrfSmG7FhgihI2OdfxnsD0N9afJjVD72DCVWTAmTbfzcNhh0N2FeJx3W5jVNCFiIgv0t8HLUwQa
wItucI9nc6NCw3m+OQMKciMmbkv8mS8BmGGlZAS8xbGSZ2wBFOwgTEo0gUVyEbNEO2mDW7Z4WS/F
l7GCu8C7ZmZ0qXERDaNxyx0TT1Xd5gC7eL0D/bHeYCTbocycKXLr828t7xyh4wFYLStisb5reTOw
xZZ15FeX09vdJZeZ0w2zwiVgITAHW29ktMcUe79rgW0vAe9hCLpUeFtVQYVJuum394zkyGUV2+4F
PcLaaLHf9l2iGYJxbpEDBuK5R541FJXo0yrhyc2AfCwCQ7yHDZ6Dn+0fB6zgUVM52e7+Zkgvckue
BohCs5wGan3jJoHSD1IrgExh/CWguLuxG3ZdXJN9HOkkJo8Lsc4oeu6dIs1QuAXCmP5GZly+SukI
PoaI3usIU4yU7+nZdAoLCFbRQ9b1Yo3raGuPomIfBUoCN9wV22b8NTPaRMijIhFiNqd9sOCSElgl
bt7uqGMuXIU7tp3Mh9nhmhgKQ4ba8skwyzFsqqHpZNm+D5neq5fKoSLFUVSlJ7FAYngylaSjgDBH
kqMW4Jb/NYaj5r9fd6tG2MLbGiQu46PG5asR0qKvUS2GQkLOst1fXztvRlQlJUn1qTeUfwudLzmc
XA3gfbcB+bYdchhmMcvMXDioEeVVcEFMPTUOGxrrMEMvr5iNR78JT4BHYM8hKjuQ7U1CI2ZRRs1v
0+kHTR1miGHxxafnzGp6gffI8ViFLmK5yz0Aqzyo5Tbwvhz2ym4hFCkoPng2PgfXixY9/UgDSwr0
3/5u9BDuCJS22PXaY9chKJoiF9YoXsG4lmAT0p6WjmcOXEHMNC5Wae9RHYtKL2mWdiuzE0zjrd6R
iQEcA0DrUJLUQgEWa+ijKnobi0RYA6SyinobPmV3JJw3BbjgFDwtaDpBfQfDBwwa/5DgENPe70DD
hFllS25tKEk1LErtOblSb5Y4PMO1C7t6KLygTsUMW6K3wWYM37Y+a7ueEQidO5F9y78BhKXvQorV
0Dq60LiYLFdIchU87L+Di8XNIyyan08Yi7fNf7D5uNf1uAvwe86J+9eK/6/lmR2RfteGKpzbgEcj
jEtDBDb8Wu5/vVRuktKtM1oLI6Wp6JS9FBqIkNBPeq/QejSs21/FQaCYy92mLE37lwhwwQiYdD7k
e6ns2T/v5ewKydxBNNQh+TONWUZsL+vlitTQDOggVoNdl335oYIE3Fv9+LSc3eY58djQEYx6M+5d
WixSduceH1sNCKkcQiTUtuXkY3xfJ8GamwYbWfdcYKsm/+OpisHkRQjbHsiLX2LCE9ISX29mLhZO
Haqs8HcWpASTbl2ewFyAHGuQfNa6TA5ZF8EuD7JAGcuPaiBBfyfyHq4R0DIr9eKdu7JjFdKa3x28
DCfiwPmOsh9Kvn6Du4UHcgSjuuDVUES8K1CJNth1N1yPi7kTnps0y5mqt3T7T/COE1RVLvtf0jV4
YIbH05d66MShVAHxlGI2tiFUaROFUIe9IHCDdnWWOE72OCVgyw+LmepgOLXhSZzz6e5Gbdqbp2Xw
7Zc/WQjHRPl3So00oUTzdKpXvD7NGpduRmmGj/K3/7gQYCfnQHTF7NWnA3U98jNdjSATalJ+5IO6
Ju4WewZoGFxzNpn6e0Yo24pQNr0fPUi29m9VjPHP/E0YZjkh6A9UTc/HA35nmTA0NSoNrU1nUWBC
y/uz/F4s4q7ap87vIwkKPm2ORkhdwEs2u98nGvtFrIr7BvsWO9glzkPCaUQ6iJtAJtk3WqOvxChV
EC3hEX/W0AaeLVyvz4DIs981grtuNLKEKM1hXejhq13Oj1EwNSmVQikeFZdZqx7/+v9nr+hPnZ2O
QkhhG2n0R31hPiCpKVAKsUArWFu/3Az6GgU0+Xujv8hnLjcr31cQBYcH7OcRvNVw756lkihrZsYG
UiQXr4bfD1MNNYihSn2lO08TpZ0Ujlz7lES93SDtmc2SinyEMrecmUK0vbCKS5Wq6X/Yp4MDjyrT
27SqjTwVkw+LWpcqeHjTpa5WsE8mZeBR9QewkI7vy0DblqtGgqBMGOqBJCq55UojKQwHx1BKETZ4
yF01tWRbDfQ/sewMyq4bKbzpK9A+620IzGDXsFjaCGBCP+s8gp2AI9C+iiZDmCVLM5VOMYncDMHq
myj/Xvjr7U6k7Lqz+/21Tej3mqtny+feRCiVynvz0mVH+ees/qu2OSG50TLYTkXTHoBhLxjHRwxo
xBCJ7aW4TuIFgMtbniwJs3HkUcIkVll4AM4MI6V6Etbx6kA9aSpw/pfRw2yb/y2JT4Dbv7aq/wPN
m4GroPzHMmigqHxZsRw+V6RGcAcUrUsAXgWQbpABzOK7WSoz+rqlsddX3qWyV8Y0YI2mHmXtdOO5
GXaWFThEQDIWcQRbUkhfJgkhtqOt1p2VAfIuJSh/NaT285/ByMZ5YbCGs44ZonHwoL0xOljee3bT
xw3v5LRmIPyTKjVSPnp4PZiD+CdbxqS1MaDWbNvqr4wdj5l+IA3udGHVg+S/jJ0YEyfXI51wZTB3
q6yrb7e72gX2qm/Z4HQLZJ7nj+LLYFDVkoFcFqHsSumyxdCpin2Lft3dK9q8Xp3/U65U1aziGpXh
fZZXzRgUKO0c1+vPp6auzxVCaoJ1nrA4sSwdthommf1NgV8SUy9xVSkHoHmjbjMQpVOLHXncVRCL
h1f4cVQJ+gES3exEvz0AagHT3cbdgstpjvIUmFzqch0gBvpwJa06UVhDnvDfd48IRRwLhBFbCsoX
uqflNTn9KtV74/7XfBtQXWM3ppMQkPIx6UhpyNV+Rx5wuxZ8KoXuhtr81tYaJO0R7Ve5laGXQgHK
BCzvaZEqn6GuOuzeT7ztxardxy3VJ/7K1vjbG2CApaWXgGKhcp9runwKXy3SaKuJTc1aycgeXwx5
HeSwSQFJQHFRrqXVucPFgb7f8ejDWgSJuozAt2gDummiNwXq3JdXEy3z2l2A5mM2WmL8RzO0NaSz
jC+ywVqAsf4Bx0hFylD7gDkJIBmOgzD5tKA6jVPspn8MUUmdGmSeoxQCLKxmA0h4NKZ+LnmsSsoQ
0ntsjX5RAMaEDJyCvLyAgymt7rgUTNyGXoulLUmK/I1+CHTqI1NNnTT5nNyqWEDel3XNR1FJpxqL
3oWDt/TZvs70fuxydc9K9G/Y6V68ea2KkMPRUUzV6oBbyipzQNYRhMOO5LOg1qED6mF/Uz6H2I4n
C/Jj8H6NreVcMoBe/XWEcmGtBvNxRUxfyxKAwkchJcZnRkwiPROKnWeRmFfveWXvRNYJthVBI+lA
IZVR+rGLhcmahzsuha639VQq2Or9eDj2YjCFAO9FU5zUCheiDAVzCyVs5I0+BqhB65IATCvJv4rj
ToWpkSPfKkQzn5JY6jh0SUA5HzCo4qtf+g62W8rfF5nwGppsxxhtlRh949K16I8BXtBNT1XSKJ+1
bKfjjQVFj7qRemixkYDAlzWAuUtr2JmYuU4/ViwPPTfa8/0n3qVkz8FYcj1HE/BeC2KiaR3YhXT7
UaC1plgIHp5SPWICnB3ALK7tSfUj/mcbJALsZUp3WJez/fyM7OKk7y/Ej0zvdy4qJAZGT5Ycaj0A
zclMF4/MQP0xzSnU6bPHOxc7CH5/7l0ono3z7gmbl7KcFVlA4Ajc+qXgdb/r0xfzh6arHUuGFuKR
ZKXG7VcXMufWlDFravhDnONKpGlpWa9NyJUP/WFJoLyqao9k11cjL+0WIhVY/mFRkpDcyun2993M
N4f/EOtiK8xp4RKMIvHTlICrLGJePZ9ienC5vj9nif3v4YWFKHudl0bs3Gvi292MaJ2W1690Wrcn
topNNAv/kTcY6173CI10tP6TD+GbppFYekyQE1ltaGHpO4t8rVv1FDBoO/eLbOJ9c65FEgHF5eH3
o+00w0JEDVsPjMVjK01oJNSxmdsnEb0Sp3g+zGL3pjXxo1Bz6p9OfYUEwWzmgA4BZt3/kMvqOmy7
XJ8vww5UtZ4LAjoQL2mVOiVs+anM2DXrsPJolOr4AXuL9OeUghQY4ztH3mlMg5AWxS+3KYQDusJP
ajW6DGM2DvqOGuAdxqoYH/JCZvGMtSp0U+VYDzyP4ovlh3xr7+eWMGAAtakRZWvgwjMTmkaF7Z8L
NwHoeBZrsWVhfTQTXQcmiVj6PAYxGrLHG7ixTyXoNZSt+RvNRjc6YCutoTIdBLWHcJUvAbcoexaW
o/EySybepjPHR8Ev3OZAFVM7zjg+8Cwy5x8Lujz3D+8aILnjPyixIvvwFE57++Wi8+9LY6mCWvl5
fdc9h5Ar6nL9Ku7k32m1bhFhtzRn21DbRHFS+1rlM+LtWERa1FeRt8fPN+KTf+QDcV9j3Rk6TesR
5GJ6H1B69hBGnm/Lu/YsKdvQPlyA0cnbQA0sh/2ekbmbYrEzI+U8m46lWe0PgyMHA2r/B8dHXjCm
OseBoj1q9p5+mm9DyJuqc4uhDCecgljZSlEtZhXgOlC74H4qkSMtNP6gMCjWhyHQmqOtM4Sm88kz
jUV9PDBx5HHmnBrMJ0VO7mjFj/l4uVq1YffHBDnHQmBObTpw/RxUrCTpZDoMhJe7SNEkQkmqXmpP
MCW8C89G3/X5cnk5hYTgcIPfkApkkjmDs1FGfpK1Z5r3IdhnuXTq5gxsaSmcet5bv3FAdNohlHDU
67t4yEMZhUoC1qkAyoXu+2NN/wBBrmqHcC6jn7rCpxl4hjBa4aaCEs+jj7tkL8b4fyNsSa9dckfi
g+J+VMVm/D37mSrrY+nRierpW0fYaf5Cns5FcgjbACnJp/4xpIJuxtEOXAN3z2JEmVANmfI6Psi2
9AuNkNfuKcMvXQflyxRlAIepx4DA0gpyfLl5TdhRp0wnNRV6PAraxk4cz/sNsQS1FIdEcu43pDru
1en5c43uk9/jxP714y3db80KWfKhv6ATyV5IcuJaLS9LP0/5+/8p/CEbEBlcCJbaSY5rNzt50YhH
uG3IU9ybicghTFG9KqQulWORlmqwcr/DLpdhXiUuZop1hObnLwf22oKqE2k2idbD7Jw5ieL9MGMP
JJ2j+oxAlhqxVtmonz/jpdjd57FjGZY5EJKWSLX1ySZNYQCI2NWBi0B6SJOA53aCy8JgaUZh5AuS
dOjR1RQZrNHwuftIAXOC6gAp2bXV4gZjnl1HUwMBPn0/QYzN/FogTVCKowJpyCJW7BPZkj1TesYw
9xUvVPWwhlpglguWMLN2EqhdsWydpE+Z2RSUHbd4BaVTj+QNpdmRPbrdEKpRX6oUKOBPVHnFNSf/
oX4E/ZSFBerhFUo7d4X8mK/sladGvwTh5pWj2goY+bl9uFObh/k/iooc0fWuBkUK7m5lZSSz3p4J
F1rEWZG98kWZnuXc9QaLx+R0ZR/Gju3rq6GnBUGsA1UpPCqn2mnGO7L71jsKx5B56DexSF+pNTgG
GrFncsYTzLyXYzm+JgTmNG/xYpiBmisHtOUiq2A0KfjS9vPAzP7wnIQGs3DdRCTpFlHEJh9sQOXi
I0aHEh6gjN3Y5tmw4GR86Jhg+QDTBu5vp/li7ZzcoQrOaQUbm19nLr42D9PTbkiJoUkRQQlyGfuW
LVtZ58rBzqo9E0jFwh74mAv3nFj0ATttb7YvgvBKCjyGXWPKxnF/V3RIfeYn72tL+Dix2PPOHGdY
pMfzD0J7XwiTUnjpIIVGRDkvgCf+QarEtQU9Nv4s0txDT3MchPa4gM3JeQnYvljkB/i79mmPT7u4
FYS1DLojzllNlohGoW4zhHcqkB1UipEGbhRU2QVSv08uLcmlcTPd5IVwKAEEzGP7LObDOUD+Pp3p
GBYoNB0nWXZOBPYoU6KwTU0jZ56UySHwazmxEQkipGt0x7lFcxGPpl3pQD2mP65oIfs3l0+M+to/
ktkfyFX48VeXhxnzVRAZ6V3PRmPjpgvAl5zjf/Hq71Qr5kkzEhsUpSlYahAU9ssZtag4d4v71kTz
M9oqU1UbHPxnfW+eGWvP9MRvJ46Hj7vOTqHDrwqPTi67yImqFOJSXAkU5LlVdvRCmmsgY+Umfz/x
WX5D7LTHqdH2zF5HD/K2n7Nr+VRx2ixscAQ7B2z2O45yDeQ0r3NlHXGKwxtLwbAcA5jvq6HYWHAD
YtoMc7uqu+Nm5o2e8VePG/QVW24bZXRNhQbqdUu0zkoFjVrXDCrhwYMxHUexZ/1KGSVqDX1hZjE+
RWu1z3Wf3xd1Y9bpaRs6kK906OyuD1iNLS6ZiI03zV7q/a9g9IxyFPlQ0wAMazNtPO1pyinz5KTe
oozLMjwoTgcPMurfznjBATwU81XZebbdSWtl0xF7iOcZ67ZpF0j04/70uNsIEpc3H/HOhFdYE7PQ
YqfHlPCqmkgsMUMiZwR9+nvP185KXj+zR+K035KmSkMmSCnazI32j03PArkkxbcM92SJC139Yw+e
jP/sebuMAYkGynk6qmme9As1/rXqiSrkoSj6Vb9i128EQt/qaU7CHuJda/Sn758rZynORxz2eE4E
54Bo4iLOBy6l9K3DCaYxX+KosNtl5YIkUGkbpQbc0zNroEH3ZlKHydLx/QF71zz5QD1old/GEmZd
7I1IR6Hvlf+tg9z3xvmKrH9PSMesDQtDUP6jRCmS1V9r7r509urQVHXyicqdZftmsmcDTLNFDZoV
vH2w41L2WMBP7mq0jv8d5hmyR7vtadhT0/moFTfcS2C0flcQq6lqKAWFJyT2yotu9Bbo0mFA0Ur8
kRJMt1nmRnHvKxhbtxOv00cJwKSOZDBAbl2b5cuBNmLkEw/8yxJ8u9q+ErjA9fooyX00nHWZe6Ks
Z3yIl74PnDGOrl51CYp06iUDkn0rUt/eUf3lX73Y9ljs+f5s4EhnWKn3mVJ3AmWeR8+mj3rdXexy
aQgBkFs9yKbTzhS6HITnXb+0Q2mhC0AQi71L/R0ENU6O93x2br7WN+ONRf3SVbYyLLQI/mao+NY7
fn0zgBszs2vHtjDDpR7tmbPutp6eyU8YPg+rqS8IJPAorvH2RXU8J/FEn98TNg3c6mwsTvNywa/M
wM+yTCLwuJAVMlLHcG/xDTa3gp8Cx6+s88oGcXGdFIqIM4BsoHFtZRzyAR7EcPJIwQfXoRpwOxy+
5hrbJlfVFttmtxEuJb04mtdMJNZAfdMf6TYCuU5Uyz0yxcDY50dT2z3nFV1ZvaCrUdtAFI2YnVB+
9ZdQQtk1fbf1T9rplftjyTJCrJOdUfGVR2j9RrfRsrukyGD77Ki/uqFURl8TraJNtTlUq97uPg6G
JvApeoJ10hOXxXrrcKXD9tT5vzXmhjURwn/rH27GERCZZfglTXMQuzOwsrZYR8LDtrRTbFEBE2qA
K2z3LUFPXTvCgcMm2zkQ9KSlmxS3BGaIoV2aPxHTIaQCEO43RoOYGOwNh+djD5d8efx3J12lNGvn
3R2FkCFfSwfU0HbKu26UM2N1IQVfJlnlYxz7uGpRJ1P4lnLnE3xajdb4Z2TmqjD8neUnZGXNrTHh
EPjBmJR1iscblEQ8ylugN5K/iYhf5RFjpYL+glBSkME9xQGITX/kDLGtlIdk4SR8fLWkbdTMv0ua
BB1U44lsmqoKqgL34JOcNlKenuZ+Et6WGhQ2ILTU6TeOc6lvnS5ArrV1okJmPI+scqvhas+Y+db+
yaXl6W4zxCy6wFfyOgCjjizR8YcPUTDZ/rB5+k9MtWBix3GNRGvec33Kc9R/4V0mzM0eIi8qbUbm
8CNAsr4E4KYA6zIlAs0RCyO957eJyDkKuqewVKvAQBLOSqlrK0UCrnntb/FFMuNC0wXSbq4rL0Hq
ZJuOBDiZLoFZKTqEZtKmpEspAb3aVueDiN6YbldayPYY8U8pHZMHnhe/NRTxMjuLBPVA10kNYEPI
s/2IGaVu2iCnl1LtszDzYoMLVTnq3s7mxXDPt2AnR2XobJYbkH+B1Q+jBmd9cqkGuWBLgP/Q9BDt
U0Yq1d8x3Kaw6GN7UHNkhqTAhx71k2DiDAebRdDmKkLVt0FfTUED9xF8WIFecXI3i38JbuNH0FFf
kclCUWR7I9sy+VB1LdHIfrNfcpcc/gK5OjZ5McxLjxmvrAOE9P+N/iWfBzGN6VtY/uk/eOrfboXT
Hq6gdPJGjFTY6nCUqrIplhlIOg84qcmFJ6hRBJ1s5cHyuTFUvvF3xK2Os6ZBHc8Zu73o0vGti9Ei
sFyZZk5QWgjlzFJ13ZPMO+0oi+3B4/6zbysO7sy5/dre2aqQOPQ2dHb2+F8Zktgw4sgVJczxwFzu
UXscRGuoPpQQMJZL9SrSTZFjW6QPVp2/fbjSyccRdwpW18vChdD7ndvU1B9Gs0vlHJ6XP4SU7BBb
kunfUeRR5pdOAl2q66rouWeXxJL7SEjbw6fnjLAJ6g3tXmjM3I5AtC6I9Zmvf09RwXLhQAJ+aYdc
I7/gFoH4GrZvvsJwasWzre8XZ2qagOV7c1jqPUlikyTijGp5JghiQPAhn/hop1P3tlWqVO45xSYX
ADzZIwIKbm5uEHerO1GeLhTq6yRDtdfDJE+qGcLYVliHF2YIHloI9PIkHool8hcc+JF2LsmUCjcX
7kKsqJBXCMgvM3XkN9F08HIX4KRvsZdpQfOzAhysa426e+64Xfkq6oxUolofIx1PYs65bVtQeABK
72/whoIfeiFjUgS45fi4zPgsr/1WBCQYB0cByhBXeWSPbmiFZOXPZGzQTNczWSv5rTKBaxEabWwM
3dMZkyIuIjd4brmmfZv62QjxbQKwgL5GAks24E7GAAlCw7ceoa/d7HPQXI0Aoltw7B2K6GanZhHA
pGeZpozk49LBfRmy6QOQFrwPIxqmLDieCVKTZU9O1NsIti1jzavu3oDyG0dJEJ46Zg4LH91vBvMF
zewxL0rJyHCA6m3ckGz6eZPdbrEvU3lKc2blYxpZfgGIfq2y4OfFQ7oR+DGLwQyAk5HAm98NQ+C9
7o0BE8wucwTyZES+0Ce2YUd8rg12nw2kgstLkDWMzjoVn+PFJXaVpM3sxRrRjWuzp0l+ln2LiHo/
5LeCF0wZb9omrRdqvyDKc8oOxK0atwGCfGNG+UZD8IdwjCU7UiR8e8YzNL0oq/0Ji3AU0vg3HHau
YxAPSLj7YIfgnbtxr1sBqCrPgarvzEeMyILxk68FucQxJ7K8iqCsBWDH7zkYP+Oh9sxZtQCMm5MD
KRxT/P/SqdcostheGzkAld1OYrDqXsALxPFl50eYrxC1k0uj25BArklrzzoEq3vCh3ZiH9rZVgdW
vzKgxV9Ey3nxqddzCZRpwinVs623i2TQc3nr7jjcOZ85+3IqAF/liaxLEubuXM8tM4nr9wsRPJbx
GaqT3y1uJiFo3pRQIW/VlR1JptB6kTKPAFXKNT0Ay/aiEfFHzzEzx3FNYjdLvIbX6tGtlbr6ycB/
61zGFUiN/pUQ0kpR9LxV+VMl0xlXzp07dJx3E2ldtFV7wmAlPb7xpRXQ8N0/miBQk+OVbTmKlbBu
aapbtz7UtcyyYudbsq/v1QfjjqeFU4I3DW2E8ZbrWrphD8LNlZuyPSrHkam2YVVb2YhqVcRC2X9M
C/PIMshXc5U9rIZWoU4hyr+z1JpZHkyNqaPBIz+rSWGj0Ff5MUd/tuqVRPJqxa3pEZ41lYFKhQWK
iTEN5VZfRbcT9QTkKW+L+x66n71Z98E5adBAEO/SIFrg+3R3L94E5K0j96C3BmVYju7wNwGrB8Oi
wknlyPkYQHRbheJyZ0OAeCQC58qQNk11EVyQcIxD0juXMOfzhiJodtyA5y0xbuSh1frJtEbMazFp
WRdObDV2AiSZoCmm4NuEPr8t2P4lOSgzcCzCHbLY7hCU7oRFqVCDf6e0d27Ve3Z93exK44dNbsGt
+YCNHHYsey67Ox1dz/9EAnjTYxQTqpCZ+FleyBMAdLu/dBc+JEH+2bziLyDFcBeE9DU+DCAAFOqj
cDwbzjFp4qcmSO9+11Nu/440HI8K4IK8tC6WMenXeUfxOzwVJxiM4g+6t5w0BeRH7e9uIqK4TnRS
JVHrC41pha9nd9uAu8EAy61/ojt2aiUHPP5EtxOxcw9enaVE86syz9XxTGnKfsEiqFRvDHm237L3
f3EOXyTG548Ush+lp7iYhj+d1FxK2v8Nk9LAUWOZiZte6ZWcIMtGmATK+E50hVKvhdu5s8oyw2Ks
YrgZPHzlUfE1uBPpEP5IlBwxGrXKHUnIuKWaxU9m98VDTWYBfWCS2jIn8gjKKLv3UzjTc/2j0U8F
3TM9hSDUd9u5YPa2G5YvJIVtKEB9Mgo5nm/F0gemDXttTpf87a0C3NmA4CcK2lj76i+/bAyJju4g
3papfV434wgiqgT06hmT+5sd5hciyDz6hLJlwxSl5Dpz/8jIJhftD4gdh0B8toUnkjg11b1+Mn5C
hHfYbQScW/WwlJH/IjL8/sVySl2hTwG5ZFATyUZLM7y8Ydth1GRq1I8EmCy3w8NxiBcIel/iR0y4
2hnE8rDIagxjt9Cc0IZO7F/rqFxdT0tqkYzfyfALqSGkIs3UpUHWW8yqz+ImQaLLU22eNZybTvUk
5z47MNiV5d2BGfEJwvF76CDQCVmnZQsTMqAUNYj/P4IDNSTZBCMA+Phuh+G8f537rM+cFvrO4xNI
1p413nTCDeRU3DEXEP5w7eR2V1jepJIFE5UmMF+F3vgJwBh/4sOrD0hoK1JXF7anxbcqUyZe5y9H
18Z9C0WqZfr2i8hI5TCqxIRKTZq9azRJ0LJ+NnDoSi/WnGSEmSW2SGWrIktV5nz5/2xQNaPAlNY1
qIsE4dWMV8K8mmxmusBPBrOueEwXM4d7PuwCQ78tSkenpT3+HnS6hW+VsIVQV0mE7EN1iBPsJJIc
knEvAbGKyaImZKmYglIblQb6Xfs1dDnkHAIKy1mZA88htdsDkXTsp8Slom7fW3JKUqUVX6PG/80r
x8rvQ8NxX51tnu5l+KCv8q+I9bicr0PCUEui0g6XBqbtb2kLtrEfRcGSgvHFkjZs+H5mHySZmimz
kZFoAlqDkG9PzIruAcc7cxhxQPu/mElwZPy6qw28LyjHyn7Cypjv9PrwCMAJ9T577HbSHkPiLTuA
J/XdvoGL8PBnSZtwSnafGEIozreo2c2HjqT/pF5dLIYCEuUFDAcq8EJvIwALojGyDpDuDqCYW6bh
rLC3Go8ykaPdMBGIXG9JXAWU3midR8C16MBpm7fyMxi6eKfGPh37VXfcNzwBiQNWxtIvnqKw8spv
L8fNGb0mGUhHx1RRCrG1+1wOt40LR8Pajm8o4GsffjFcuTV+0WAYL+zBqAfopgfB124jTTWr66KP
Webr1ZhzqDbTGqjLU29PZRDto2AU3XhKLt+sCeZaCyjkQREWkRsHlEyQtS6Wy24zkgm8fAh21GeS
9qIlgnqAFR8A/hd7x4XnoVtKIq5vb1Qt5KC4X6kvz1d0rxGnMMOGVGXvSI0WaxhZJTLwqatW+40H
cLsV9/8F754coggUO8qQm+Qyb+wH3QFKIxYAmwd/GGR5zzubVqkA64OyX1dobgFpiR0P3o4IKdGT
1Ih3fVmYTjRLjhBbPRWVvY5vC+m0ruWvV72BGEtsCQKlP+OS1rLys0BxrTu5lKqNDXzX2CACS7hC
lQDvt2iuipyMXCP0Cb5eUtKm1xW3B2q87ERu+fi3APrVbjPWO4jhn77OzoCveT+aWriGTVeXVe12
NT1Svr09dprb+cCUndI4ra4MSKrMj8nSdqsmvT1KF1YUaeryEii1gfl3451EOmeerzb1MDpoK5wb
/SI4BB19hKPT3/exK6Po2BHumk7MSeCQ3Gou7oLrYO5ojsenWuOVtHDuhJyKQ9xOaXS9cpjbxmPV
RkgKndXZTKDvEcMKN2QVEIWdX7I7TskYonhVF+GmnWoOBpTk7RM03gBlxCqJaMB7MBHx6Vv8sHsN
YAS5s3tKSfZPYV3P46iTAle+pjAjzi1Y92YkDyvO0Zaf929KJBRZXWLuuBjv94EuzyP9JAz8lEyS
TE8rXFQnmHEkLwCwTsLAOOuopzs8kTY6ra/PNArXvnOOD3570Qlu9M6u4DxrnMWcQyOCCZlHOyBl
rG3kWy6r26GQgrK3ZkDfHn0aLH3dRPE55ffZIEQJ4gytEhRoKN7WHAHhhVdoefQQujoAy4TGMdA9
ZWGsG3GM31G3Koy+i3tBnnJJcajthIxO5nEM3notnDMe4kmKyKQjElDxZNw5/NlmDLGxPnLxOCHY
lIR8Ng07PsYKpeWJMJMs6xS17VOXpXv8ypuMhdznoZQ4h5u+YuW/S3QgMPDzNbrLfY+pHrsnNaZj
gCwDN9p+qSDKqS26eUqRiF9NCo2g50kxe6GvhyxPZScZtjlnBEd2vD4ntDHqkmVGjXiDBDYh4hqf
n4znAlyn7z1v3CrfVOeXvLeERE5s/HezmwXQ8qcEligQ9LBTT+ZOy/cMc1X8Pcl176/K25f0iAQK
+cfyaod3ILGcPYM0AFNFTynOlx5ISynLuV4IiSYXqops8wa6Co1oukmM51Orx/FAcHBa2xB7osW9
MwneauthYROwgPVe7W8H0A0icCCLe40HY/c+gRQR6sVceFKRq/XQr9g7ygyI8Mh01njqpYuXcDKC
7RH8AtoPG6z/5MWXqMzKAuaCJ2OnKFhnFB5IBiLVba1ivf9Rttef0yOfB9XmVrc67EQk9J/KeWdZ
RYZ/7e/0qGYH1WAjfxh55yBP4zzlHM1us8bMNwAancJyGmg9XfV27FHDHdGp1x3oX0z1rWtzGUNr
dtGdoEHRJgFCu1qjZmmFkUH4/rzbo6JASBh2T+mqz/6JUQik7TZ3LYwSAGY69MSh7KQ513SbzpbO
YGqJqmEjbvDXnB+sRdrSmn0XsMKejEBv1mQbHE23yTU1CpT44gMWBwXMHhweLv72lGyv5B34i32A
Tzl+kjZecBJ9UVjC/6Gi/7di9L3cxN0ZuBt3TaCyll9HD245MGJN7X/mnNIJ/1Tbd+g4K/RIMqhY
5cqcVd6QwkvqjWjWns7ya8LnHw8D7Qd+qrVECW0GZSs5xEQV/mnBY/Ost9+g8AiNM5ryhKqJv6Fb
7p7wz6lzyXM4E5jrTqaOVPYGBZAMiZ5J2E9L+Ei6lkwtSBaaiYbLDuUcJWYBFHriM1xKYPD1vnLR
9jfqGBqTvtw7dG5KD4TvOYzJj1Si+p9DXiYC/4w2A/kfBs++qpd++CIhtYiPkOx1NKr6VLMWOhB7
/J69da4Xx1UgzYkMTEwrGS6utIEaYYpvJEusjlGHAOFZlQufertlBITKL4WEbLNoPf5BNcod08YK
bKJjoiYeblFb+VTLdDbieSxO3lBvqVs8Zzb0/Vig1lqlI8N3kDdUjiAVLJye4lqD1BtB25BnEAg0
Iuvf6s+7vPoLDcEJL4cKAdSRlozI0kclKERk1M+T+KyJjzby2dfKo2UUTP7GLz6KAa7hfrVlHJso
DSxG1mvQlV5qIcnr3b3ABpDs214EHbAjQ8kpvgb6L89tYPK/cZr7CuxRD2PgBvNBzOMxPAgXX5S4
Uy6zqkOxp4Vz00PzSKem1Gtmok7+ckW08qCXKcROKYJ5ztHZXmFI3RLGy6izvLAM88YcQW5DeCry
NnCmNgjoJBZq0DgvUC2EEUlXYelvgiKGkzW1Eb0rr5jYGEChNKgGIBKVlBhzKdJKCKH2+NYqhE3a
qtvbPUbGZxaYh4YDnN2vtGhr2OUkc+RS2igcJ4KiD9k/iLBot+x6VfBOAm3RpQpzYlGtuzfJ7XgR
9iRMAjqEZBI670y9HzqtGrejmWjxcTBIBMUrRgvwAak4coalAgEePUl6Yj5BMr39hS6hra7qCchP
GZYRKW0LAIHQmqKf8Q3lIM79fXn3c0sK3FTc3AcLjl9rpjxOMNSxlrifjV9u3bqfsjTvJWITUreT
QdG4rMtr/DLxvCnKaJnYhNhhPuCN9z6VM9fit8TLkkYWR6MMZCNVkbkn1UUj0q0HfBDdz3xj0rIE
pGrKraVwX2sybd2lXqql6/vc3eMNEpaNDOQLwJhMjWjym3Vifibq9wczNmhqD++DFPK7btch8OTz
FVxa8hRnBU2m0uJ6d5EsRrRnPBg3wNpTyFzniPh75FT1gzY2HA9ccBnGnXOf5ZhIq2hgky1OZ/AN
pr0Yu1R1BhrPBGPHFxPT4yPAmvmDpxnZYlP4eVoccBQGGEXB4WxSfj+IpVBIS8MsLNZgO+ddvPR+
Uephx46c1/Lp6LdBkMogJyusehw2wHLisv0tI2RFJ/k5+NTyTfQ3+ZuA0lL2vAvktgUQGrEV2qXg
V+YpMAtzD4654iddhH0JygjpO5l0vUqcCxBhChVlSU0J3yPxfmBIqLqWRLa6pYpQMQsVUAI5bYui
35lFXs6DvDMnCi5sVhOVOGhuMZznCsL9Xs7J3U0L87ybrjEG7eSfSSUwnJlxEm5BLUo3oJ9dbhNp
iKWzbqGO+WbrcrNRXuoEOKgnj15kfx3g0ljl1W1YvTx7MJ3qiEm6xHLsEp/yBk65HSUeB9EzzOJH
Fb/stQVU7yMYrEQJ6YXRSTFGfvKOniwFZx99fYTPLYrc26h7JtTa9whNW6uu8BlcNlUM/N+Jqb4L
BoncoiZgZsJZSR1uoGs2ALCjPC3r5klMYcoLXaHKKGYjoTtwto3pSarUZFuZoNrMbKxl5227s2uJ
n4s3EFLuwt4nKhn1Qt9QUXqfpkXoZQSUSZqsOAjCN5m+xbYXnRcjkH34nF82BajFsvDUqBoPxb7S
3aYEzv4kQVTTxL3CwKGS9UDhjvDNqylJ5WNUNsZe9Fwy5ZmGkY47TjbUcchOB5rX+ZxbB2iQJImT
ZP6PVoy/4Pm0pdejSn9Tp91JozU5GQL0OxbaY6GxbBAmipV7qdZPwmdteSqnmzHTBMLiHeOurNVI
tqK3jFHAUnkzKNRg1uAaip33/BlF/+0GSfrXQqjMIKTr1ybUYWUzItR4cDwt/DkGegA0kNCaO/Xz
xzPLYpaBpFhKsNSNbyxRTr7FtDAC58Tdm6oKzObER5JInfWx285WqxMG7ZsoLbEtmVjRPpbNCfRU
SwWAf3OF+o/JMpbHjFdGFU3gd/Ko95ugJzGRK8hOlm31KRmmc2RTFqGavUv+RQ0blSi/jNSACJCq
hUAM7bMXQUHQKMHNjrWxIydx915Mlj/bNkJ5oIpprCTmVPMFKzWfvOA0zU4ygDlnzI6d3t25mJe7
/lZZrd6vFJq5ktagIS0Iwb/5gNiycbzJVaGlShLpjCAS5p3cGxJAWTZVkrRJq7dif94PrG/pLFO5
z+MeZ5dFSa8DZoG/NYW2b1iy+VKM0VBUfm59BwwEh3tug7llWnCKvTlkpI8ZSu14MapYy+JEYSOA
4xMBcBekGupXaKnil0fOLDYwp5RHWblI7Kq827EaJVpgc37n/ZLRtVHP4TkSAs8rTHX92E50xVdA
59d+XIi7dS6tdVL1VUiUBZ8ib2EfNuh0HxXDVNC8i2HlHsZkheq7EvJ4WJ/nVkIIyjuYHgOX/kjF
NWM61wJ53nTZ/k8Qmif+L85F1IUhzKsomRhBEmxL+MDNr6AChN/4+5PNKpdsMtwsyDTkxz33Spip
rgdvIHAAgbiiDLx6zq3uHjO9wFZK3QC9cOZ0AFqToTYJnyysg1CXf3TSUQIneEA/Rgd92rTJ2Vdf
qqNCQV82kt3+Nz+te0qyPHumGyrcBlYYatLMNQ2eR+aSdeHPcMmMZw6ienNjryAfuDtLklhYVrqG
kJgziHyEIG+lOriYOHPE3ic/S7JFiEc1ZqMkeTBdQlH62dBq6JTOr/tM3DIob24Mw9JbFeb/dxQV
vjfkJL3CxWtgx9FsJaTHl/KB1b4SW7D1FQhrVx3cqv47jcZbMM74/dGLvhT7UcK4pKbBH62u4wgB
bchh3IWSRe4BrazVE9cHNS4g68ndgf1NiC7ascnIXRGqvaGR1hqZbaDNuGRblNYYOggk3r+Zzni4
85MBTZd3gIih9WViTE2FnIvPOZQ3aKStUHpuBnzg19rO+86Lp84MGQlMQuh8wPpqOB4fJ7d/bNGw
pswBn+cweAOu5NH4Vc0vB+ccqu8vZcwPvD98bPa2+fRbXlGmzWgWC0FhHv25nb8eb6WXGDlHxLDE
a975Qglq2mpJ1r9KMGlf0CH9UfPk51wLMaGLsdTp8qlsCivRThZHh7O2e3xmqolB+pcgX4ukqm1T
nWikiTBCaOX0aZQcNldEe3aWw/DKsZmA6eI7bJKVSJqkm5E2rdz1uRPwyV9Zej/p6SopOgw1FB0L
19Wc+a43hDCpWhEn+rjiA8VclXVTQnjokNC1Mtyae6e6S6GGR8baRyrO65jVofKbbu5S/7g9D40v
B1nQguoJxCHAjab4XtsZSXKs1RtxmolZYzSrgXTlQbz2si8iKsktN3wguzZm3wf55UXN8a3QRQUC
uX1u3G+cFCX1BVZqdHzKU3FtkYMtlAS47pywIFdkg9XclcuQYMzXxKiHlDdfULrmA4sb9iT7xEx8
373aZ46rdov3w3mvfr5OV7WDDg/ZUktsNR7JxWNA3lU5XiVmnDAoR2yQ40o2AxjPS3aPuCdc761y
8At2wp1YAf7+aOqrRj/3vnZnldIJa1dAH0GlkqAQlVxoGGeazBezIT1B59uxueMeLesDJ9HpmAxa
edWzObkgfORXNaKYGAqSxSgk+pndZj1u7IN0QxIdIetagtlEfGMyhPZSKno1rtnhd9otDQCHO5dr
vkmxQ2RO2ooInLTfmdnjSmdVSJi3JJpV66W+XJAxXv9LyCrwgtAJZ/8ypR6dBD65Jd+kpfoYEtVS
b9gfcZm9pMwuiFaHRFcSaktA/VwB5mC6cBLuXKrXid+gKqU=
`protect end_protected

