

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ahdDAHzz440n+Z6SrLNKLMBChQ5FzHxmtmolGyaGzRzZ6AsdM11MYnHQlmkXolfzuQvsH0tiYFpA
bdhL84ynJQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qd5Te5HYUFbAOVCK7Nrwmf+xhp7iHLV1qESGeKRRemMuPlhm9gxKzGI5glBpEm+Bt6GS7xBHPesU
Rh2RxY+9Nst/QoTZG24XGDjT8gulIAFW/37G7vhPLNVOq1gP33zQ0iNDRVgAsbEBqL2aP8fzO3c4
Dl1oSNusYXsdFmxhv/4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0n9Q8CLs0GcRArqoXB7pbLNq/7iI54QAnaQ3YfVTrcoLuaPhMipi/u1YxvxCeQhStE/q36RmAWKU
vuVvb8WRD5dX8Gc/5jIRt4ORXRhrtme6cizBVjYhymzdNTAgbAuH8k+0No3YXlnw3iXuB/bUUXlS
9ThgyMn0i7erFTJ6h/eogbI8EG6TwEBPQ11D5xXxMjzz9Q1WQ4L1w3R2CAYnCrSSlQxqvapc2X6+
HzE5EzvdMpbru1PQrGeGwaFtvlT4dq9BRwJcYQeIth/77QtTOb09uuY2bIUtRjnczrx+97he8zc4
F2HQqnZwdLvPbSwwqlsUdlME2ell5wSO2A8Cdw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fXi1UCgHICyjHcoUzs2uXfr4QL3Zd6fFq0YYnh7DHj/Uz2hpTBP/xGkihvbT84E9/Kgj7lZnbxyU
NW3Mn3WgobnvsYj6dHFEG2LfnPYpGw5nhTQMawWoftBXy0o+AjB6W5RQ99l/hgORyzZ3gEP6q1mQ
SG+9quGTTiRQQEHy3Sg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GxP7neU6pelOGsRYeMpWhq9H64emJJW3ch5ZqO94Ja0S7m2rL3jKbNa/UebfsafxW/Jq07+9ZHQH
nakVk5fs+waKW7fPdCvasFZq3bHVoH2M3uf0FMGIXnsyGlgHQ4qCnawBWxPqrfn3SKY260XmNThN
PHkcyDSRI2OjZKzXzE7AHiKXBnUYqYuy5pZkIRpG5KuuXSL3l68wM2qwWAk4Dy7OFak+VRDwWWle
Ve26y55BBWyX0cVH+A1y9sHRRFBM6x678gQjaKYO8u10cSkLQEatg4BKcHaSLpXozsPkT0ktveBN
etZKKhExPa6BnJyzgqh9xypSTFtCXtbhEF1Eag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22208)
`protect data_block
qByBb+9osJlT47Xa4s5iJtRattP8ygoWQtWfGy7JKqAOYOCts5TQ7/st88g55jqCH/JVRxOiXR7T
ZIb/xpADzV+FPbHrs0iVDYs2DKdD7Dwb1QlDY4osWnSVA7B4pCvrOQJU/Ta58vQoIDh7w0DN3all
XZmBL5Qvbzy8Gldf2O8IZbJRYj9xc9FG1elfGtpDMxIcSubivRWgsEIpdY41wuPYSPrFpHWsG986
3fs7t2EWulO2q7JnF6jTDZjDs6orMjPep013Euds7VR5U2h7lGEuxu4+zXSnpnSNx1pgxOa4qZ0H
l8ucEWoEhmJzu7clwZ9mWJBCeZKGsaa77NAPZ2zvKupUByBPVb3/9BM79xhRLLbi4DMYsL60kjBo
oOJ4aumcEwi96WnwSacD+wI00dh3lZBxjXa1x29QDcoObQfYMdAmXBuUWhHZTCjWtZOTb+mISSNX
0UJfDXNkSZ7iL2qt+ohggNqzOVZxgvIguSFvhqyW1z4gwPuuu5Nkfrv4Eogy5Vay37QvTg3/ePZ5
fXwLTbn1El9AvNnYGtK5HntYFPMtke3iIzk5x8PaAT4BWBr8srEs/LMUabiBWJHwgRtaiW/XEibV
apE28Sq+Bh69kssVRxOYql4FpuqNBZQ0XR+cVe6F1v6Ev/pvjCt/dHRFiThaK9JvmvEB6CpXDI30
u/qe6e2c/6oNjMuPOh6O80gt8I1L7s9Jtg2rs+A8K6vMxc0txu5skm3dMmazOtUT3tRVQnwVDnDA
ju3ItS0Q+S8U3c26IHlK5ThUjKjVZkrq4Zy8XU+893Llo70NB+Pm+5YB4DNEJkJecXqGZ/2YrK61
P61eQCto3LkQrbM94ze1Iir5/FtG9LxJ7AbEgwSTweJ50BwvkpQBRkLxYkGWPWw08W0koHwOH4pz
oW+SoiJv9FLoRl92SbcmbPthwcjU82ZWt7qaTaPz/v67U321CnCPC89W4ZOt7BHF+wByfEnycinY
iWKeAgBwK88qPeyme5QoGecHmE7qM4uKCpg87iEx07ETelQB0rVnXl5G0wNGdu6I34bFcW3SorHr
Xsd/4MqKQ9wGLullUkRuc9IUUq4977MGgoQjpoQid2b733zm9JDrJXG5PKdcV7zM86dY4F2kLXyJ
buGK+7I5qfzfccn6wrsyfMuy0fROBy32qmR7Er9MBZxCbatTYKybRgcjEKyeq3RRPrGLtzLyOy1e
KhUkgB2yjIc+jIrIP1e+hBU0vzs67nMx6SCGXaSXSMi6P+9ki5Dt9wteEnVcval3aaT1INb2WCo6
szzcI2rv2lRYeMPqxHfR2p5v3WS6BNafGOgtNSEBPfUH2s7UShLnvPraEyH5CswVzqTbPevtWFoL
Pl/DLXTFJduhi3AF3KdWllbMpO8oOVp5e6K/Qr5WwvIxsm25N7A32vbO+N6BeS1tSGA+mr0ezWJt
Un73p/igvD7btVn6Nh/C36rBnSc18AMcaX6d+DgvEZ0U5hHkENlFc9UNxFw4z+4ctESFW2nOvse1
8VnsTo2Bu3hGLBMjPwrMvE5MITyDAXSNRY9T77voPZr8HzLe0/ZkVlhJYua3wh8sTq3dbegbmSa5
EUjNIdDkK6G509YrncaBbTHH57p5Mr6We1Br9D/sUormMrZw6GVPMvwuftNJoO7JtmTT51ZO55n3
ce6qIskeMuZHOB18cs3qjwjpT2LGOhnMhR2EiJRIqwYtPRC3Ge3hJdTmjIJphUmJ4QIL7kz1ZhnQ
3wZvCm0Dm3MGNXjz169zjKThe2wmKtcu0B/msxqKiuB6RHA+H+pJU0Y7X2/aUDVceFaS0RaTGjfl
+BT+VRrCctp6IyyqsAAUL2ti0nyjCY7oIhgvOAT8wliX4ONukjAr2cmvGnSLHerv/QeEpQ+AAXiK
OmqpZBtyqjxE1f5f3lelJSS3NEcUFv2rjTkSeuQRbZS10ejKpIt6RWVX4a4SsSbyE3/IFWyusy0F
LPcsMQeqE8osvxVFn3aC4rpoHkyYwYtupmno3Q0YNvFUKIXmJPIIrYV0ma+8vDTJBXPTTQEumDvf
aYmXMfMpkRwcG1vIE4GLWfv2oL6AV9mhFzXqL9/9wAWBgAH94X9tWHknWNMqoPlaE46FHtmxrwY3
+Du0GDuqWxtuqNzax0f9ZGeAvT1cbZIXDfQbQniGt2PQa5aH5SRXR21Hy3IiHzltSPleNz1Tuahq
8BYmuhXSXmiNBNWib9tvnFYxDL3E4M4esxUP3SPxjkQvZJVCTOTxF377l+PWpeQlvsxpXz1dCQMH
XngwuZYoWABgpqqkAPIqCerTNmsfeMCymft5YoHBaHgtsuHjkRRgVJvAGncI8ow0gcEXbDABPoxG
HFo7iM/bQcX7JcB9FZ9Ag/o4S4RJutP7hLOPkm1bxn0a+Jmj6J8yv3+c32n5YZWGttmrxeHdwhTF
TBGbvDgreG68Ue297JT5XeV8UfCZj4k6GjvsIV9i7KZC9+f2eod6x22sFCoEktJHZ+ux9iVp16g4
QCdExwuzxBaTzO2SEmUXHTjq1SxOUz2/hr+osOUoNehQTX53tZ8stI2tTri+SDO7Ob9IPx7sqhCa
OKu3Lyr8Gmk24Jc1I9gsFBjxqOyOosPRD7XhnnEqMJP7jasJrTNhTPIpsZB7eON6qKwdefxl70yH
US/4VLcpbCA6pP8JP5kmq/RNXmgOYhAWN4yZSXgXWpJ/9Deo3WGfueqqIZGLm0fWUuI7zhkIqjdy
eY/BB16jHJMcG1asxH0EDiLbKCBjFIR9PEExps8CLIq18PIk9Ad9pjd4c28jiMG4xzVR4og009na
5FC8H+IjNVwUonBSoDWzyP73KFilj9tG0cuADCN5qOdhp6uWyeuV1MpgypeBNrImc5nuRguCdwpU
n1Xuxb9+78ca1r3/QMnr5nrMbjFnXHgbXpTvua+q8NBbExlIQs8lRjAnBJg0amXM9slzy9zs4W9O
TDSygrQoQdwxzSlpniGn9QRlLQ6lxSyXStM1stxYODRXkDYPtnKR/fLsyeib5wJGBZeITV/QWSMl
kToAwPy8Co6mLoDOCNPUI04Hd2sBaOwfXZNIlrVk7EFCj3syOFbFwoBy3nSLcXyinPB5nnz+LLH9
s5/AWrfbFUIJwWIU4dcmvxMwD1DhHY5l0cHAfbpIQDlhLJZbwD6formfUFpXt7jXei0kJQv7YqDK
pn4h18PNq0Nhm3+LPcQbei6KZnYEZrLNV67CWqmWR1b4RXThn/Xea6LIs0qXMU1LyaNJHw7ZETwd
RSK3vrCw3CltlZKEtqV/5uaJzQLOQpPTgcRTGb40KXBpg603lPqawqt66GiRbzAuu+NNyuO5OGPU
oflqov2nmMF2Zj0qiN5Aui60WATHLun5Yi9bGW5rbqlwPNC29xUW0pftGi4LhJG9xWAX9jgysbXR
9lwW4eBXdacXAgZcUCoEUg4BEtLjHZSZHqjhjzYzbtSWGd/7vPh5OUBg6PzY0QG74qA8JhkEnzoU
wfBK0aEiXOb8TYT9AAJU9OA809V5mdI4YAYmI5zz1rtBdal7mw1X8TptzP8krZHob/PQW4xwby7C
vNAUj+tCdHFnq/CbyIwUOsQkdXBwu90/qAh2ngmVlp5fFrKpLMNffLU1HM+VOD59TC3GFT7KVD0g
uIS79tobF/V2x/Wna8D0zCCtCyWkFVEaanApWmAWA54LulYE4Fd342K8fTmj6kjmXTA8nhPF3jbU
g+aWZwpgVaqsoEQt2cDJu45KVngDmN9xJ8eeqUdzklL0ge3f8Ep66RsZ/FN+NDYHEnP9Up5oem0B
6X8ujjAmxwGV6ZS887P/rb3rvOgkj/ToRrHK6qvquqiq6YB9iwbcsHdcr1pBevL2dewakJEUTYIt
R+N/6RaoZEVOLRxYJemtcs+eLrubSs973HTOqKZEJtqWvFBFN2iR/K6ZyjY+sTOAYaHhZDca91es
PD8jNbzb4r0yNsqrsCK4w2t+928iqxOeHDuqcRY8YGmSlEQ07dgrY0nvGcUsdBTUxO+cFZXecoLc
CmgR3M3M0N2j4RXg7zIXvAU+yvM8t6h7MMxatpqbLDO5FNAY5ljnb9RB5Yj95EMz6LWrESrthbBx
r3B9DMXnCDT5AfQmAYOAFjDVVDnlopLR6zUEGFcQzmeHWGzAvLk67pQpe3VPajnM5StLQYKJw+Qs
VurMaUzmq7WBwAKFgCl2cd50O4z0h/p5/LltrwEyE+0KutLU9mn7X8luZ3laOwLOQMcAqoRuUl8Z
DHlg1SD1wUsa3QzIglV37qrvC5kpQ/Afmy8D1ufhPLEeLnC5y39ALX+SsNnV/6AOcPK5G/0URltS
ycTLAlbgNTzSSZuzFdA5ziIcycMgnUyUM5qX1XuWX8kMkd+nSGdHvhthz8uv00Xu9QUcRHZbJmDx
L0Y3di9byDQAx1TGZeRC2WCZRh75azu9Oi3Rlpn/Twf+K9Sk1rFt6hQE+sQ2xeQ5ZNmm1ESVLBVs
JJ+NMZ2mK4HZcoAzvUuA+FcRFbNKP4NG/DEOFSn02BgklH1GjmGCI1fTbUSavqx4dbD8rG4izdLV
hAxbzlveuUdHPshpUCKM3X2iiFC8frD78WkLUA5E8m1gLHhNniy2tz2H0lNXzrm4n+qvFDY9jynP
Kk25I/vy7aMrgVkkIU8/5MApEKD1PN2FudTlSlqXnbcKPGhHzzwJvy2Es3d02XLAUvkLVf8wrs1W
wqeXOA5XeHKtWSmxLmlIm6cBtqQXnPGaNGRE1RdPHf2UszkIkQp1xi8OPx2/5wcUrFYjHkp5JIM3
kVMV97V/NsZbjrwA/qsID8EQ6qtFzLmkz/sdtKp9nNVrMOFh4mf8n0rCdN7S5uYyJ35mtMGFy7XU
4qejGHs5fPE2p3YeZ3rCb/qtXoFCYuwK4L6Th+uQOGe4XCWSnQWRUIliVvhA93DAAFJA0u0oWaTT
K/0c/aGBFFH6hhbXyD88XEqpt8NjotYM15kb00vFOJ/ag7i8PbgfOWskipvrF0TQNsT9Y7SFc/Wc
fvwB8tZaGUI5Dwg2J0y3jDNbYVC6HagKogWbuuOjzVw6uXX+Vet87rTVx5Cbyet/ntOsFkTCnuCw
IG5qeo575ASBALF9eFW8sW2XONdaNNZwr76wRcM5z/qRAiHyXyWFEnKjrtGR0xgVjb7z7wopt6lC
gWqn05aUTiNbrKmyCdnUgjPQTdWp+8kr2RuG75cKY45bysD0GMahOpgoSm4l0uuJdfzJJ5SvS7qq
JUKSO6TnxCw/NNxf3glkoM/NLEUvFlX+qAR8xvK8UfA4cADpdpfQEJfshJWF4vrmRUU2RZYd2A+8
DjVToIBrz7Or5Bzci9Mp+j3STdUGmcKT/T9BW0N93cFO4P/AhObwVnR3DYTsN7xDON4WuVr+odin
CcRCL6L+oKnyXXyzCIyov/vB4xR6YfrnhMgh8tS8PzsshGM0IMFMhnw9gHoRlMQj+uI2oE42U6ul
cLury5xY5AGKW4yx9BjRw7Doj8hCGudWGaS9eQhuHKzOeWK10w3TYhtktr3knRbURxZ8a0AozNrj
9PFyi6b1N+/UY8PrJESjJ615vZaxhn+4Ocgdooy9FaF63gNx/nvGd2CC1//l+pF52pGnpQeywFTf
VP9GIomYqMOjvl6Z8WPXZ1qOHp2M7SERkyBeny7EpD9z6tT0KPMjLY9ktHZ10zokJmCgitTewOJa
cVE/XiQagYeaGq5QnZfHkM32Y+m9A4TL+lvF+ZNsqbUEGaEYt1dUoRrAY0XMBByTJ2GLbBrJT1pQ
BgXjDH9/FIlmChzHDC77RWLoh2p4HXpjpkUJchR3J/HMKIPWOCZ2xfuuij6aIJ7E+m4F2FnFN3HO
O2EXSjdWDtfq8DEOLQdLjLx9wOXNNMw4D0NgAj4RDOA+gLhbWtAhD9LwS4oaxeqfAZNWAVb0apsh
XHw3lJVOJDycy7kmsDo4GcsQ+I3vcF6SgpEB+rct+lvt6ytY509WbXVm3jUaSlBepw79JwH54iX6
eTkIPgpaiAyIrWs5sGwJ0t0ZNIaTZx0/NUSryQxhIJfbRM1K4yh8TRiTAwvvgkkS8c/Hh96Nb6b4
MdyXBE7PwHt90sk/Kl1dwx+he8LlGfU3W+f0dEUHOWTcqjF388boB3J+EXwFkzgRugmQvTlZaD+e
r8fdVf36ZdbyTZ5LgUubxS5J6CcIRZiz/Yi0S8kO0yyX9TjKzv6fyrYm45eUXuYgf8iffir/rNsg
sJKNpiHYoQEujzHNHLrc9tuHbmhwB9ZvDFpw5a9agRaJwrNQ+hWufHE6jJs7UYHx4fSmLidxLsR6
DsYB+wxdyXM4wpHu4+p259JhHTNGMwkuKnC1fpDNBy7vZ2Gnthg3kO+QJ5fJKUbKRA4xjYLJJ4PM
Zoh00dqJBCeY7xiU0PFCkXa+88SlM3krjLLxQdktdJb0TsIDL9fP7IUD0pAv6ky6Uc1HYe5QL1tK
4TA3IDIaSDkZV66GzP2JUBlifssZZ77FVuZ9uX+cXOTI1CJWxix8FSDKYQc2gBcuoBc97TzDbYV+
MnDyLpXzh975em1VHExrLWd/Oug3YujYept7NquKBZYpx243j7B+gvbpQy2uIkz7cBcnP5rXuzQf
99JewIsQGf/6eeI15q3L9teBsT0dUCUHGU9+xh9kMO5J2gp1p5jUQAJv5IVYYbkb8AEqPZCWeYhO
kdcejPbxNc6pxatvQxh5+ijsnET6E6EvjSU5/a058j0VXAt4dwznv9y7hrUkISwOAQ3WLfBYb4wP
N01kvMjZ5DrF9JSanyhqXV3Hmp6my9pv97xt5hQwxm6Qqnc9RpStZwSAMQWpNeOnNol9G4AjxOJq
K3URlgZvG8mCCp51C6HdoEk1Y9FTSyA7NDtAgdQVb0UjbONgRhKRRmBuQ8coI4uQ6U9Par8SKXyx
k8ST0EfEaOZMBQkxn2dZL2fnmFgRaPE/2JNzWQzlbOc/FmGOUDE0kWfs/YhImkY/mNJaVBNHWJvX
hp+dw4Vzq0wPkDZVqAATmxE1UBP3+AUl8nW2/iMn8O7znu5UdcrgX5MA8b/6u48k9pV8xwDZn+wt
UUUMeO0OX1UMLuqlnAe9ZFYbq96Jj0phVm/3EBohzKSPuwLe1GDTlIuj8qKbuCSDFFrHfFKX8rmp
QoO3spBR4n0XO0GQXT8T4Ta3CUZZ7ypBk+PdXvcci/zzn1MSANx16lfJEk54T5LPbknxX3Qakx8J
ncnyGGqdixkVbxioN/5sQW4fuAg6LmIsUz7qgwbAjSByLKKgQEJh7AFxfSi4ns0mR2VjyPKQ7FDr
88KRiQRknrBtxapP9MFuz8WnsWv0xyuKDBANr/bq0RIsYnUlxjxJfZERAiEKuGsZCLFSNSwYkblT
O3ah9369Q10mFg0wUh8VxEXwtNzt4wxvgOLcPa/9jFXxE42VhjnY/rdqhPX+iLL5PkvgNVLLmx2+
gmH5chBpQbzbKeX2cjZjeutLBzim9qw+YdzAU/1C1X98iQ8VdeIgwSYJCPzcgZLn+hhQDTOPlXWs
dAaZh13x0Z0p6RdAz1BbawK9rnQ6GnLbf+4JUQAZLmysA3B89gQiY/Dw6kNHkmHUTX7D20GQwY5W
m0BM/evKjHIzZpQWRrmCnNLoM92I4arYasT2W3hFX+iokjJORWs+ckR4z+pFVDJYqhGKMOUBMyIq
qSHPPihi1cER8FFhuBBkkkL1Djuf1A2cXIuyANiXuPEP4v8s4ah9g7N38M56DgUWjUUZ4SRJdTXs
tcNv+zeQ24oa2afhy+8tQN1xDrC/YheGCeVRtcjA5KbeuP6hoCpg0witBU2D/2EZAnD43Ve3F5ME
PwsQAYUm1ajNbs8GrzR4y49+VpHUyWHMTbDc6Tcr0CcVcWh0QRuZRdNGap/AbpPOWigrSlec2b/r
hhOiNnw0NbtEbkfXGlDt3j40LgVSmSqd/9WWpAmXDk+d/ItIIBPiuMnvagzgiJIBZsOPoWtKPv1f
3MpFE2ISSjaET1w6iYb/B15DOT1SbPA4rUbkiJNhC2mvpG20u8izmDigXpmkIND26eluCQlc/asj
ZXXKVeQTajZic9rwICwez2ISb6XcwGZcpO4tF4tv7V94Y2aIZ2QB8eq590bZj7+O+gnW6+p4QuQA
aBTfNC/ZWhyEGe91I4keN07U3qmgy1kqQkP1+MOP7Yi7zsfGwfiV9iu5qQHGqRx6TGZchbQntn6T
/vJOsfn3SxfHWXZVzj2fN4FLrKqDJDZhOV/1+H8Brw/IV09bcbwucRcF+FTE2cnES/8w1IAGWu5g
9lDM+FFz27LNkarA0KUgdDxxcl4C6er6nBtpXt5Czd4UBx+5G7xADyyq1oZolx+8QmnqS9GeqEsM
UUA+Y+k83v3BvDIAMsHDB7Kn1eZg/eBS7vEMtjYwiJjC2yVKCmV9eMXr1/r+fz5tzjlDHfhwyLd3
9jI0fu6GJJvdtX/cFNMgOf7EDXLGlTrMWW1sN6HrANsjnje6HWrHV6Yaz9zsDcVf1Q1fLtklgIoS
00xIuTNh4t5wtxHcFAB8DlOD+5TMna6H4Z733rPbZRWMIwzSkrWbAP8ERgRGEpSP3xYJkIlWkyWw
IlVBgWC8vLYCueMnGvKYB5UG+PWSEbE8A4Q5/3dKNk0IP2yb2i7ZGNVBxEbtw2j2TGCuTrw8bKWv
974ps1/CbztmxtSaO1t5RbzZ/OL9mI789meVr+YuFIV7/2kiuGqyXjOmzaenw6LUBPntyRFY+eMr
PkwI/jA8L7/fvzQ/nvUhYNg9Zs50DpnR+zm8xkagdd62yqOoWbtq9mqqQj1YCZU2liPlCtSbrfpo
R7YvYC9d2UAaTdE0go9vjJ08VM1xnVFJYFhcgJT1UpWhRO03j+2Zve4BZhjFubWpTaj+9F2y2ip5
9YbFJplZ7FAUsLoJEDD2UpSfL3dsc6wkj5B6VErkRL8r7LPwumIpyuXbDDE4R1HPpcI0l5ZG6Aux
davLvB1xIoi9uQxG+PNdzJzJNh4qVD/7dbf41BP2aZViVCMXbFq3B/ePen/E+1zLA+rcNBgcks9i
rgsot3piGteecwzmhJz+Jb4r/M1mIsOi9vksJLnTH8LAcBhxjKjEIivH8ECzJdwTKimOJ/+MQuax
ConfZBA8Ic2IJWLE9TmXpr3SHdUB2Ic3p1gnINZx1ziTQhh1nedJLyLU/pvetbxo3IUGSD9XIee8
1ayAXqashhKzCp9NlaWpwVKBGCIZQmbTwX69nKhYYx1Mi8q6985OTBNb9jM1TL85mrvUEL1JAySJ
KqmzU9h53SUDuPy3MyCHDHw/KnztY34BotSLpXeGTFapo/IHjFHE/cFU0iVCplvvu/lGnD8mwI6A
+gcLMAqXMh3Q6BlGXqDbCrFqKDXmCy8xNSCQdP8Web51azd6Xd891bb9PPg07dkFSSwBaklQ325Q
O5SBxUw8QGV0oCkb5vozFQ47VSnHXEokDWnbuktDqaE3awJ//6xaSbWCzwK0ueARBpoUZEpQAHPb
fl5R4gU/I2SiapBo/Zfkhg2emzXuTCij/BtDnX30uHOHQX9FR3CibSlb24NVe5s/ARmjlhBekyk4
OmaAoZFqVIWb3v+NTGkH/k32YJZu/UhXchbbxgYAteWIDBmrnfKOYQLJ8qKh+iYNiNSBeg+DklaM
NjIaAILe1Lp9vFc06AUXC+aMVz/S7h1+6iK7TBZteBsSFOt02vT6KGaDC0wP59dUHHVh0NpliC2p
+4oI+cbLErB6lecemeCeiTIDvYbS4MkGQAlwYRLlMzM4dqmmVCnIITj2bwnjGE10cvsvc36EK8FE
iA6PvQzS8oh2Zrc36Q+2LNJIlai78iT8Qecw1eMoa+NeloTxLDv+BjdeGSBsuRdmbvjrDd6T1b+j
Dl5TBOjTHToQiKS9ZpQrUdT8Nj8DaIFEzRCuVu7qgzhzMgX4fogsZlz2Goir9kM0ZzEkzpg4TXrH
Ql9rL45150w1iil593ckxO/7GutsxHDpmzdazYM37Q87ZtWPaBlXpgEZuSVp2dxN2S4TQAq6pvLT
AEGozQhGyYzMOyE2opimx3i7KhkbOlD3FW7ngO6orcuwCyy3+VEWRjvOTSQbkdc3Zjc4LAKrglEy
TFWkvSEJSse9Xr6cft7Wyc9kBzqgi+mUFer0IcqxkaahAn0FcIgyjA6ROa7uaJ9rVBc8vQGprfhM
HdcJ8ZYDNxUYUF2AZH0WwytntCljAuYoH3bpdj0yO3I3bp6Vo3u8N200VSM2cQwMhl3qCJS7GRb/
f+krICNcBDtegX+pPuaFFJnABSm9fReFGD8OaLNaX2DGh5oUmx39njOwkdtqfij9loLL8jmVdrdw
RP2EogrzmPp37JpvfpSfKhh+DHTNEq2CXz8u0WwMXIE+ujNxLe3VdZAHGsQJ/rDFkUbT2KImjzRl
TF5364lPwyHenRhiYHCeIvTGcwg77AdeFcbZW/QlhBcyv4nln2o1ag7DacbCW0sATnaj2Ps+lLA4
rf6G/zu3LUMKxtmaB3mTGjGgy9dzCMMKDyGbkPimG9fVvI+sxDuXvHcMLe/g3oZyfRUIy5ncyX10
c5Kl6W4so3XjzbOv5rzgwPetWu76QUTUxhdqpp6kY3O59isFuxlTmp+WlN+KzEI/4DuZF5TnAvHS
TDM+yxSElHbp1dt2d0p0HHtA1k/kPizjLqLJayWph6ylLjET9C2h0vJqwh+csbGl5+MUhmsLr1n/
sr4OGk99j9odXIUufs27vy2iVpuzwK4goq/bACXMTQwo4iER4U+Vt/r3zhuHr/IW6eyNwkAJilPY
NoGMuemVvFM/bA8lKqAr0h0g6OWhaVszY/+ap/1GyFiOUQQECzO+b8zctCJnJ54o7kdPlhPWZ4Yi
2X9cPVX2SUIT1upUr7ogEmCLxeN4gihFC1LQLacC8XalQVcXOH+7hZK4MJcjT14GocceDRnE8wsS
ymCf/O6H9BGr2Nxo/SXwrZPxq4objSDRIY4EnrRf0ynzDYDZA4cCRzE3FOnf2vMv3wREO10enX0Q
21DiNIW7QozQaBYuHGVnZhmO8R1tX3EKeU2Gr0ymPM6XbHjzQKEMbBu5rqQridtdU79/x9CjksrY
O7gm+r1H4LMzjS1pEnfebV80ixr/Sq2doxq+AVffu+Rme1UVOSe6mv2Un7V7Xmyc3m3MXz9YNNiv
lC8Vi8cdxVQH2N4s4Z9yzI5/zDwV64zNkOQ4SKiSisWAWQLWvKBa8H/NyOgpwGubeZuY9A9/gJGo
Gt/NWnX+vJDs6CQJv35Q1/Ab6BbSZJ/bRNFEXxr9jANvcOdDIu8nccu4j7oYbHdXr5UIQyPj4+Ov
GJAKGFTRjF0y2P9Sz1ajy0S0QK6lz8tzJeF+WdeEM5fAKHIGEWNjTYynwRnE0eUgT1xkjNsujODb
Q1JbSnLqmkZ7l/lbACMfasdAMBsXBPBAeXRQw3hOaJ5rwWSWyIzqxKZfq2VVE9oEL/dB7LcDJ6yX
Y/Dr9oXcpihT5LKSLxE/RF4nftS9dpWYTo1kTOiM96Tq4QDb5OUEwu/QfhHpjoo3FusuXlxcn4iQ
ALbbgVTYEqhBogXKi5TD9Uz4vPpGJgHgSYqMk7B8ewzaIfxb2dr0h/S4vxGU7lVne05VRsfQUw5N
B7TkxHaIQ4YOQZfp5+XmNClp5Equ3FqxYIiOJ/JLGap212d1cootH/Na2pz9FHtVAHLQu7TuaxRM
b9pO2gLT3yaY1zx4vOY/ADihwCEWa3P1cYODaYC5K9TZbrvaKlUenZkc2SbSmH4WRsff0sH0Vo5/
W15xX3po6wtuej1YtcOcX3WtA+Lq1M+HhFNrCDkJ8bg9OiFc2GALO4dQv2qt5zFC/MVzMc0tbCcO
GgkZxLdoSa4lItnu16cpt+d8QRcVwupNs/7g+G7/R24OeY16Dv8phC+7W8hhJY7Gqr1fed3hB4hf
KM3C3rGy+FKnrPownNphABSNgaUX4OPeeO79jvCaz77cliF6c1fiiV0C0EnvYC9LE67wpux9FfRg
ckcbbdJRAJSVE7T3i5QGbvnQFxucD8zt8ygcuk2zkNYGIuOBFv83gZBYXIfA64GvgosfyxXI1qeR
83l1aJrYbsClvGW1rQJh1Yde1fpzLjdCfj93HqzFJWtQLJNwV6ene2cLT9WndAf4qUkJneXlyh5W
TUc6KqxyCNuAN+SFqo1DfUHJvqCM/wfU3aPfEKXTBOIdN1cM8uL7EIUKSI4Tls+Q7jSJTkYy9wU7
8kUMS+w91NzI9WYQPMDMjt0qVcEc1mRcRh0sgWG/osXW2bLk9RveunY6p6VuEIgFS3YEtdwJpgiP
UiZaT/JkECroUVoog5zg0gJQH7IejMKeimucotFgTSd70jV+EIqJprwDFT1vB1QSZq4RFjUjZ+8+
3InlqrBt4foAE/HYepzWrXKxxAZiongWqQhOe+MSnVu3W59dP2+UGkoPSwLwp7Wvcd/Vf5N47Iht
YuO5/SpGS6FxIuEgzxdz1k/HDvFDQfz7ie30p6auEXNVwdfNqUTL6sG+gan1R5HvKN4s7HbeGfga
Bywh7DaB4bVafffiPCJyoDTVikKFj6dex3JkYvH8ti8b9hM2PcG/duN5gBzpSk7l6XBEFwxyuh7G
2xqV6VPJnn/M3Hi0lDZxOpT40X5h4IKiNlcsJBDgLLhDuY/BZAPpqwmOgCBIEnJ/d2+VCi2yJ0+J
e/E4m1Gp5OFNwfebxrqWLLZ54mtU6+DvrXjGUcJrUOhSYJwQiSPVPxXWTqptZaQE9emo9qL+/u1l
+poy2CTPv0UiwAwFZ1iRi4bL1fZg1KUywrQ7ZB3ky9a5D3euhXTPJxoKQtBYBcYD0FHx59q8ga9o
h2S3Y2/MB1uLOZUCBTNeu4gyLiD5GYp/Aqrah4bdYC8Po0DVegAEb2/egSmkhcZECHbGquXPhWVQ
mqewcz1bqMisiTuk4iF0FwVn4uFVZgpmlzDJksIRuIbysp8RdYjdCrdwZz2C3darHqL9dIgBFWM3
x5SK9oNjGjVHXMofsNkCg120+dxiwhS24akAOocKEVQmEbwa9qYE+LrwOM0RL484nYcVZo+QSk1y
/vreJkLqLjiNTNzJOR+QUnvlrnnQQFFB6kUkGF8FUwKMVYoX71e2Ivx1kP/8eZX2h4hx1z3Kf+b1
AzOvhxO3s3f5wKj36k/zOUE4X5S8y8BVQXtnqOwQteu37r3y6LFR77z94K/zvjE0kXmmWDF9n236
5tCsja3o37POI6UGak6NTUNgGBpaiyeCZJCLYQd8vTeL/cAoJ229N5D2VExdBhBxbbV2nCkgBHz4
BOS9NNa5yLitNisL9GeIKICkETvxv6UdwtmZVZYonytOeXOiG6B8+FCMn/ECxckO84cPuLu9UDRA
BJffqlc+ygrIIYBiRt1A4M902obVXlL+h2UkNo//UVs4OeLYRMuSl9u641vbSoBT8ztSaSIViMto
g+sEUkcpxExTthhRESU50NTRf7Y7X2lAGb4khVkGFXcGl4M6+c2ZIWHlqhhsBNkc5dfFPTORnete
2laKH1FdyZ0iXpWiEcLm2hir6T1lIN0RhPzjngV/M1/GEctVUmJW2d6YJ+l1bPss96kO1LxmPtwm
icf+g58Db5bT6mxPGKCgqtcMWU/2YTNOjwd+l7OGF8NBM6cZ6/HkK5fHxtcvteC+v4hqK43Uou9m
EsGJwP6EWgavx/kABZ3rtWsEIEBAS0BOjPN6tVc5CCPasBFlzguU5JhJXOnzfTzyUpM9wajwABHV
pQmvZtobkjLd5nO3NZhH0ldyz0LrsPszlj/8nTLzqu5mpZ50cqAzXeyRDilBaRDdzZCsLtPicpbO
Aga1QImcBMsaAASWf6Jt10d9coyGpWcaWW8HiYHej01PBzbJIGZZOcioOeTd4f3VMvTrD/ct1UIX
HTqAfR1kya7JdE9Zy9MkIL7zdJALpDaI7ZnX80Kadh47hnfX2JJuCYiKud7UdINxlY9Kr82IFwWL
r9aTeg+Ly6DlCFOdWeG0RNjS9sA2M+sNBKqVjyyNY5wvOMdYfCyWOgcsNVb8Ru2Ub7HLIURRQD4v
qpZzv7iRgqvQGR8akoCpQiDkb5ZQ56NE8PWnyRT/GXN+A2Gz7UMjrUXQJQzMs4GC/HGHguBv2/2B
Kj2D2DOmNMfnVTySqmuylT9N1UODViuLnRpK6C5ECXFNx9XHbxYVWmhc7PuR9NeOvYLFOKy2wa9d
2vM4IPZxCphjxtP5U03q4CCfbOCbZCDOn42OfK71VfpOiSlPEpgDA8SHXGFN6j/s0j8lOnnUvvLX
4hC6n4EUL/rzDGmmVSE8B5/kdc1SREFyg1AdnAEIseOQ+dp0rz0hFS9vwIbAfuWW0IKfmlvw1dUy
e1JQQnGa/5Xp33nnF2yrnQkQqyKp0Ou6gHIKRMP1mRanyoPFIS3ADGfjCz8tEWyHBOp617t5/Zhp
hDEollR5mEeTx18u54+JZCYT1Z1X+ouIevcB8MfdKGwusi0Hm0M06i2XTWV35DtgEOHb1MrVmgVD
RY4+r/Q5YPIN36X9V7AiNpxgD1GW67s+Smeck4ZVpbFvkofcEYg6RKxLzBTgsF02l+a4W/W1mkGq
TLW7P2gOdTdbJR3FtV1B7eLV6etELAOA5yDZ9MyvadrbhBNRXcmVndBcE2kvRr1e9yEm7SqMhQQt
9IPx6zEbIJB16tOJxWg3BkJ5oy/GJLrXUKbCf+/Kmfri94Rb8dbiHoMgIC8GkBRSm7n8iqIg9vsU
GKyM0HRIq0irHb0NKdpCW+d7QMZEGIDEdJsU9u73BgAIvJS8Zbrj55B/hCgigpUXWbR0wXLsneqY
OZtpykUvhYcDu52wuWQSpKhgb4o8Pa9ZyOdRjZHoWFH9bV5SL2LBQNkfSpOlF4sHmvY6IdaJI/C2
uJ5GPYugJ7wF8oQvHP1iG22xybuSibz1I7SeeKBcZZtJN/RJ6BzTMd7a+F29rykrnRhlRKKcRtQ1
VGnehGGWqAQGv5Y3u/sW/Qlqy6lWhCPWaGHN4VwSBm91rImcW0XBus4rWm48+50eQ1Z1vK1IJ25C
2R0CFPFWocr0Y60uCfM/5sZW50llV6rPfpGwPgJhbD7vc1jCokiottL2RC4AOFgDMMJv4/xvs9qG
X796y4ifgiH8jhtPqxpFrJPf3YBMczwPrs+iIr4kXR2oziSfeS87ncWBdPWgSY0/NrZScy6kTx3L
AeBYFe9d8dFh26/DgiRoBambiwzLJSFReG7BHByglSE8bjnWUSPQguCqM4CsO4VtaN6Ray1rg0f1
B6JyqRLTDsqopg4f1YVkDa56T12iYIxZqqfxZkb32AhI9edXakylJ5C7DTdt351vIIHIUlexCrmY
ectqzDW6LIA1liEK+R4VEncfrk3W0RqdqrmVBQO2+oysGGTmMyozoPPVB1gUUqoQsN81XmyT6Uwu
6ET3QcRObbUw/y5+FNJUXwizrScDCzHYNzKDwi8HwhkvlProzFXHVlyhZGymJnAaOG8HxYeZe/2t
w7hn+MIt6awSqaHDoYkWIuMc3BNxIuNywlrE9yXFLskZVqxYF+oOQs3DQmi+FCYZlLmRCTinqAEO
MK1BF3KeTc7VVYW94TPlY2gDkxHliERDPw/cq6ZmeUx1i+IG2bx1XK9+pmkVn8AjoFh9Lm7YaM98
XzdyEENBvYbBDJyei3TPbR5ZVKQ0tnDwaMn05z4VbC/g2h9zYg6EgS1FhxKgDxWbFXi7Mhz3Poar
eqx8TUCsLQtWW7b1iRhBy4I2mmUHV3LtNTFac7xZ0KCZmA1RLMwbBwlLXz/H0g6kQyKMFGUsjabe
JXqVO+3p8yhVprhfMkL9ij7a0hnNKVfb0hRAlLK55vA4ctv9N92OWztjStKXbITjXTZRwbkJuVqs
XbXMxrG4jmtTuwCrCPUAmV7Lt4Ti9PhbmMIKe2gJqZ+KYXFLXx7LzA39J0thGkBcugneqZ1bO718
Q3Yj+pSJXQ7yH97j5C/VP0/FhyTbisc8EavIoQE0hDoc0b3nAYXkCN1OQHZB5LCGrJRJIJkNnYZT
8RqkDb9CoSCRzfj8hI26ZhcgxDXqTkX0LNEaqsW9Tkm/F/nQ99Y4i7WY61pzx4rkrzQ7R1w5fC84
ChHH2PcgKQ577BBj9RImVwQXyW4O11l3jeHh0zul8i1k7/iJp3hZkseCeqwV3bp9TsDDgLqgQ82Q
y74mY83PBWH8GFM3S0EAE4xodTvUZaIthzMNIhK6OEWT35dHwDk04TxbrLRDNmkHlowMsC7l+GjR
zq9dZubqh+heMdAkOIVb88sjDASfSh99J7B0znBnyQHT5sZdzX+yBWUe9tAKyE15yTlTevXM9Sv/
eJRAfO1GzL5vB1B3EaNEYfTta7JdvJ4xoKzk6bd3r0vGPv/cMOuUjgM4BKzATj881s0Usokq1Q6l
vY2+w8f2YlZBswM9BWC0/IC5Ciuior4kE1LllQjqw6lRKG9FhL0rB5ihx/8feOkoQvV/jY/W0pQo
WYoA5y7siyQtpEo9DcDTTAmJ3lN4OH8jZUeH6bvbXKA0Z1EZGoEIIu88x9IWwBds72ZLPUgs9l/V
crooWo7G0tEATUZYDlx7f5968sUibWApnhVg165IwIARwTW1Y6cy5y0lACh1YOCKI52Nx8Kd1TJ9
41GYGn83QtXOpv8D56m7tMQmWR8Y2NFjQ7gAwtIOBPP/CBkQWdo+ENCeD4tE+q/eUXrJ78KlcF/2
YtcXfsPAwJz53mHiuMFEQ9lNV2s63EB4T6KT0VrAbOnv/pWC8U3lj0vMv8zleMzkb2S+UTdZEYS9
LIcjkD4HFVvApTgtuCKJsnagUCRmXPuQq9WpamQuxofOkCAE0y8sS1VOqgigewyTmKRsbndcBrZ6
RCo07e0eK3p9H/mEV1+tns6SyJ2+oA1PaT6/uMZSX7oWSBDGU9etU1uQmgFy8OratM8iHaKlj4ZD
66Rl6rmnTkk+sqWZq88RmO/SKpIvTqjHKyeG+pAFjwIVN+fSBrD0aqhhvRKy13PaUqQJ5OVFqbHH
7kGvfEGOjVDdpIclRcKHkGQ78fLUPWZgTIB45+AqAqsi3B78dHFkuk0rKEplKNBYm/X4C60D7P7S
fiDi3I72GulKr+9uVJ3otKzNT/k2n+f6sUMwy9y4+3lx44nD8xX18+Rm6WKGG4fXNqSVzdLOIoEY
//rbhIPOoNpZNnlD3VcVSxgnSe7D5Whiw1uhBJ8ZRGtaxX5hGjVMAzlNWGKhouhbpBzlbf/QkQ5J
WYtLdABPZqymJshgroPpzouRRB81D0RTG+caCLOhSpUzMT0i+7K0VCsAPXo8F/Jh/3A2sm3AwZGj
KTylBT3bwWDMj+s7/vj5QC6WiPlTeAIjSMNf3l7t5OxgvRBOZxHjyL13wcjJ112RA2EXo8AupPD2
h4w854lAqqVRZO3wCZkpbbl59dpev80cqbNKYCrtnD8H4rN6Q2hgbhs0DxmWLEqSjHHFdGlm1Ad5
kdGeSUytnLBlabyMaH72hXSM36+D2JORQyPvU++1mThPF+TrJvDm6ueIOzu+ug1B5Org3uRFc+f7
5/cw+X1aZZwUVvY3ujjOHvrnzwwmc+tzXA4oKFsXfnrnsZKgQVgsLW3WZToIsmIpOhGORfHH3Utb
XG8Uu189o2X0f1rxavCDjmxaXmBI3t/1x+vdlhhctHh+Gck9S1sM7qbLLtbV0GAIHkaziy8itadA
TfCDlgeDCKxW5L7J686+OLrBefvc82iwiWim5usNI7yYUdot1dBCiMPOLF92GpeNDodwGRlQ3pne
cNXWlLGBJFn/92byE3nzW82I/c9N+urqUeVdsuH98o7JCtd86+MPKKfiZT+HioNynH72vMZfbC/U
jmUwURrjl/C6UkfRnjLSAQm6TwXH2qEFuSo3ZUNAWFpm1NP6G9wGQMzjYDcu4//GfogsTrlU9DEI
xqIH++HbNKvpbom4WF2sfHPWLQg7VNzLZZ3GKq5w73pyNsni+Pz3SjOOFSEQFl6yNmXcoxQz92f0
gbz/A+9t297d7LtyQSBVF2LDHY131XzfOW2jM4meNoGShPZ0W8ZenKgvgNxevDNyBYaofyGw07FY
lDdUAUUR5ThuT6sfmNpRKGIJOtFps7q++flMHdP0OfSyFWi68L84n9FYLwXmEWqqBtbvHtq4Fnqo
GNABJITBvhsnx/xwJG1sbSA7uWJS1wB53FOe62j3h0wltjCj3iUx1gbX10nYpsthxSgc/HlGI1yP
Mka2aDR3M+JlE+T9meWNNtju7O/UxcmAV9a74Vbf46HcuQvnOj47pyFVVNHdTnfvuweImTzFXj0A
xNYfjlyNT+7l9e1wPUUgr2GSCZtRH9RgWIbIF1doIJ1fgGi8ZLoK/WAHAvA2HvQn+zYMB2TmSlbC
KXwO+7HQiwEfyezK2kIib96iMYphF83wRVORHB1US19hk4If9L/jDHzE4QH71f+ae1vofHQkeYde
eVjbaJWKpVyTLiohhsKsB5NzE2TEzU7M8Q5mmYf5tOLn5d7mQS5p24M19KgEklHqsphIHuj/oKJy
dJiootqRXU8YDB6pfchCQ/a67Vo2iL03l4uE2ng5p0w2Os/M4pyUh6ZAna0erqN6hpSOOvOEXAnd
mjLOnAXsaa7RIUwoPQy90xDME/4lqYV11sxU303aDXMSLR0rcWnp4f0OyCnwnVfq/taVUvEjsmTB
JTE6/P54wZqgp6FFmtCJ+zr24V0Sm6X50ydKgKE3Cwen/6fuEI1nR8K96nHdvEotShYhbSb24Chh
cc4aM+eg8USqVlRKeRJ6W3qE9HabAqvQ0GHsti0DG9HnUvJOdYoA2KLDPpCvD8LVmgCeWV+bliLn
QTZIUlJIrCTk35yJPpVOQ/gXH4qHqeX3XmXI1s0s8W2SIMFUAO87VngztsOS3XYN+Y3g1U8fqswa
H7qQPk9HzJ8SlLmTCx8HSONvQDv5n93SAiaJ2SdSNjCDbT77RHBxfSbERWqjHnPFqdYlIegvRqNG
3EU8Y19ZSeGM5lOiHIqQuKakyIJPA14RzHTkwtxGwczpYwCbYTZ70fLqYk1LKmimUIGCuaziV48m
UQwEIuf4V0oBgV4FfpNOp479H+h4f7e19qOoUULz5G+WJxhZEA62TU82w7a4/GoeXYIgYWYhnNDV
Sc1OUP7guBJFlI55FUxCS/QpHasGIcWh04ezFiLaJ7JjtqhAezFvHbkofx6yOLWLO1Q9LIgxBgeL
wsKKIbcb+E6muMD0GU40jBgYAx6DSh+XuTtp0b+WfJAFPCz1lJ7mQNL5cp0m6AmFAwLLe+BKuejy
SqHIvR7AW8bVQ3QUUxFrhpFW1Zpm5UxD321XaLW7WYLJuKUeNA93114GftaIQnCaOduRyuI+F0HL
SH7Ej+gTE38o9QgQXii6PxixepN6GadjZUC3fqQMz1O2o4fdFZTBXgZ6wCxAlHVUEIfP5v9FCQ0F
m005cpxORH0nURw23XTs2KBvHBeDdC/Jzo1fd32nXVrpm8+8CBQBAmfAvzXhnUe8yVkpQhJGGhI0
yrjknoEDMCYI23zlr5geECnbsnoG5M1IWxsSU2K5dfsNmI786Kv1XV4pixQ5qCKuqiSSgZA05t21
XCR24FPdUPTsmbEBWHDi+xy++kwTCPD2WF6/XIoXDtvBc0v6xGzeMh9umaCN6OYQZajIDTaIGCYy
86iIDwDzYWQoF5Wx34StUlJzm2WqFD5scwUGNbP+iyTnDbztLs1MPv5e8TKrANRZDWNeI+QXxglK
2X+h3jvBpz07Qd3wl6wYKTC9GAIsNg82fA7CKdaRRyi4MSptTds6iD+ZixGjH2pZzemmwwg3jLi4
8Q1Lwdcnpj6MhgH27x/OwrIhWJtOrOIVGKJfiQ2rQop4OHs4g0+KYaMtylmqF87JLcnOM/FeFp/B
MT8+uqrd5tcPAdjC4gqh4bXZOOoBubhQR0kXCZpXBRaCSsUu0ZZgZTMcg+6is+51mZ6dMqsXkbUD
1keZuHvelRQpI3UG3h0dS2b1NfFW0QWd5xYh1xxE0sEPT+NAh5yE79w3wJe9yMg4C9HQzNrSuYkE
t5EzNfLeh8CGP145YwRpG+QZQ7V1lVl4s/GTXSaTVexCMYFUPVcFQSMIAou01SV7ITFStXV7i5mP
vM2V+upvvDoXg5AmbuMc6j1NLycXXvM0GCp2QgynPDosmy4ZUm+/x0+F/zZsx32uVg5/cCsNdG7a
frdtddN0L21jhEX0eqsDWf57HjGGZ+hTSOz+uCqUmGhL9kkmsnTR20fw2XZeBGo22gVbPgD59DEp
/bJAYxWzmf/3sDdjNfvqlekoHF5AajwLlFF9fLjN1AN3xpyqPdqa4l5lQ9eiEJLb+7UmRLsnl+c/
Did4Wl3SZyXDVaI0pTYbxM2Ajo7RYQDW+nyP+Mu/ulfMkEqHbdT/2ljQlu9YHSQ0UJ6iT8AAEgPo
JGCXgUvTBqkx2XD9hh2F+iOrbKWkEtOt/I3POnPhuvOjDG+Wb1zaUMjIpMEUiNwwpcx+UAyGaJhj
Kb7eQcaeZhIn76jK95oRL9PcG031iW2NMqIeFBo0uW3ecN+YJICXLXAsc+bKqugRUVCGmhr1TluU
g8HOpHhWZVycF+5xkoVGllZjBCUU7J5aQnwDm5iYRXsvObYtbznhTs6Pp9bA4GsH8cBOuxQV6W4l
l3iDIOqumGNc/NhS9RgYo6W/Aa9G1rNc6DN3NaRkuAfMv0aaBpWEYM6WP5S9/2urJ1k5HTV3Or+v
cEwnMHDtiqMb+CdHb1nBkJ/Rs3vOTLbjqHDB1pTaUyHx6uYs4EeXNTRZUW1rLzmuY3rD1m+RVIGp
klesjo6FXGYnIEQy96GoEuMUY9VB/GSI9+wYxt+LvVRBaJ/xGoX7HKpXHwz6K/O7lgputoUR4c3D
Dh4JZIn6zNupFhnb43uO3aXB+4epATpau3JxouUiUzvDZYtT4WecIrthfy1/qg4sWg8AwvYB5Rzd
V5Pq2fB5obbdqklpHcJ1f3YMirOKUjrUV7n7e+tvbUDfcjiXBT6Sbuanlix/pjp4E6A+UKw71bV4
eQ4dZffpn2MAHW0M2oQtZVUVWoAVIcBsp2dCMjrA4TsXbZURYjdcl5ditktreRr5YsvqR8YZeZiQ
XRaKeKCJTnt7SYI1HGBjueLOM60wzUllWhtsdInwuVEax1lLyq+EtZttW1JoUsq7MFh3J2VtXPNh
xfgPLM8dpN3EC70T70X4448p4Otze+lT/H6TGs/RcMg+98u0Ueud2dxLDNmHCx1Y3O62YgfGex2O
9CfnP3rM/lhdXhZ13k0MICHJwyjmx/BpMtW1EYEUPJ02gn6lJump7cWwJWQBK9okk71WThD78X7x
f+1vER3PdLIL5eV+mGFnRr//YaFi4Nxhf0oJlMQRE9kk3c/KPX2Dajz5tSxgXQ7/z68WfjuEJn2f
iIGKh2M7WEf/TUZxAjaUdiBzhv7pQ6pgPNH7rsgN+7hiogrvXMHgsGBHYuM7rv49K6Yp8JZ9myCe
8yYv7FGukMoau5Vt+1rVZpQk3Fmc8z80ONZ0FMMJwmdcbSvAwS29ucdtuxUUNuesyw7+/G9Q7MEB
mzzFrYcxmpNdP0mZaMX24vg3XIuON7FKI8U6CMWa0qX7wsavnwX9CTO/GmcefgETzgcVhwf9LQfj
ah3S3LzFRampIUBkQ8FoDcrqvmTqGIPCMy1V767p5vADyTnBiQ2pBJ/z5lCCmuIZGUVQhCzYhyEo
SsIQIWR32R+dJ8SUlObKoIbIyEQbZfhkGVK8Zmpas2oy/YeB9NUP36qn96i0C3lCF96Ocl24F/2p
LUad9gZHBzEJTKyMOLMsq+R8rgc/UJ7CjtzTJkEAad2Clak8RTvlUNblXjltU74WSotVSTdFNj8V
vtAd27sXnMMxXQw/vpvcVMatKTyKKNneO2S4LGq9CBo26jud8VGggJOyJKS/kZNCLy2Y1ttn9Ww8
UuwcUN6w34oJ6Caw3JF8T2HA2YRb96BEbxDzBA/LMDNDDYep3ymrIhTFud38+AZTpyCYCFjHAGZc
Xh6DeQyVIDKNlp8P1fRa0+ZZtJhL8ubiWfaimgbgsfQgaX6twy6yTngDyxyppw+wLVlTpvhuUTMO
vYdNEOLqnX+5isKuVdmtUmQlmsOGTM09TGi6rWSvyaqZ6boKdUaROSBZ4fT+kZAKxsLIjXu8ebxM
NyK2550sex5H4ycUAXSO3/4riRkjK00lTEZZMuReZY/6lJ5fNFIG+GkS8Z5RUbcxuifk0tFDxpP4
9ZECMFVHadIq/o0toKwLKggq4JdL471z/M1Xl01NEI4cgoRcI8Tsz16HohOxNTDe9TbGrAUgp3cT
0TGeL2Ry3mWjEHx1nY20hJjjbnRrQ1lQTv+IB7crAWjLIeedtQUTA0L7jp0Sf5sflPR5ogIm0cnV
qcDt2dA80vXLliGXznrZRCgsoiLQY9/+3A41lQNqTZ8OvyDmksR/Mf2UjOf3vQb28I9lAle9SqlA
C3LF6m67mg0DtBSE1OnXDbnzkpvpmt4AEXH5Vgtg4x42oOu9liXFmk1ANFB4qnAo8c2VMZFqoBzx
HCxN3k/PqrZVWttl4ek8OhBgmlUH244YaI2A7LrCNNuUZR167F42FwF9F5U1kpGis/HgQkz+vVa0
rGN8b4ab/pFhda8NjXSm1pr8Iq/91Bo3qy50XVaZRNAHVGeNTNVBb/6kWrwih+BY8ARH8PJBIyau
KCsymfAcDX3hZIhMj/juNTYjaIMayheIpjlBoeVh/FMLUNKJ10x1k4cTmEhBKsDe+LMd3jyG4sJn
xq1uQnDWpWthDFhYUUWaNX88zkBkk91HW4Yf1nLT15+gw/XSeYZ0T8v/RawhXlANJ4Sxvub4+sjr
S/YWtfu5YfpT34H26G1iPs6GzfwAwGD2rqM2SGGHxUBI/SdYijwLJ4kco1G5wXUVS+7llad4ZjeN
MfwvtsDqyTtRQ1z8sbWLvbE0SfZeBbL4rLvyDsWu85r/5iGo2FICwMvrYQ4Tm5Ns+ha14ZvDXa9K
4X7qyt9/wVjGKSX1uBzmYm1UZbYQduRpMArPbESXDAQP31g4ft84zYlFWSMOJpsbtM8+83I0OXcJ
J+c+c5c3ldin5k0CGa0tw6KsKuLL98y5PAskpziNgLcyJXcsJH+Xvg2cvltPivg3Kemewwc9bIof
zKdPPVghejxurs/uwOqFqrAXlvSfipeX+HNFnC31xwHOewHmOtpHUu+SdfoV8KwAJWPsZOkezHe1
mfucz91sqBuieJd1jaQhM7wvbbLVjaspl6si8xDceRAsmaMxU5mG0QFxoaeAOCDENJU+2pFXB9cZ
Wh9GGQI/zxbDeqsDC3dmbjMCjlkGHb+mngumPFE/CkGmoGim9qGWiEWFDjc183yOiBUMImJMGZ7E
4Q+4wu2MjlxPls4HucHgtUJWBx0Bd5WQ/pVND4LNLK9ALokXK7RATZ+sVIzIMGkOwoqQeeB3Xz4o
e7BEfvuvhqFS/Of7g5xyaX99ZHtdbfd59duYMd+XwEGowq+EQnPJBGCoZgj/+5JdRUP/7OI9F6Ii
zs9qkjtcmO4+MbcSa7rQyvQBe4ps9okBnrk7ljLfQaUUFRvyq9W3DLsw12Yl/ERnG8MuGQj6y3by
hZxFwPFDLkDUVYU0DXYJ19bdmgb4rpfyIzTkzWU9TA2paTkxMwBAnAT+gNKDGkjgNQZxNKys3uZF
qNMiqxSjeKamU+R0b5y5ScmN8Zdl7OnLnsjXAX4gbBC4c8areprKQNKabzZkOCPmAJ5fmvtEVzJ3
nqt79MVQ5DRuq3tj/AhgqipVymuRDt06a3cJTKhNI02wHPtxf5Hn22jF0eNRo0J4gPh1fulhRhvP
D2CHvnNpUwhMWnfQ/AqY+oBApkjQwwmD69K2oZvBK5JfrBjT82MQN9mfViTfUSdAtvD36V9uEwVS
AjwKYTq8LfObIh2SUYxYceM7UkXKJlBsoKKFNpSHfvHWqaopeK4UQYANCncnSCLrUBmizw8qk4JY
mT7CdMO6xxHZ3YLEovSoiRgNMOKmf3yXxSwriiTnHk6nJUvWoqjvq9AoXsp8CelivBu8i8iQLt+P
Ki1gAottOAPTMsUxZTaYGbUxRSfUVuhiPi2BfoHHrB/MyPk+PBk+UmVvEpQxEKpQt/TvaOrm0wsr
nUapfz7z524OgzPfvkZPqhZyLgEnIObfuN9AwG4mF1Aqp5qyquuhcrUEkfieb7AHdaFEATjOZKuS
Ujwfl7Qj6NwKqXZXXUmUAoG46CwNkUgPN891gCdrBj+E3tfwc9yuz6PF6nrE4YRzQyB5pB6vbEEb
sH1TERmE84txu+G9E13Jisdllrp+/rsDXX9gs4xbWzd+8kV3hoojiAMi1vCiv97dYPUGVYKL1QsT
apgC1RhA5eIlZo+I/VJo9orRuKtC86GV4NxUBTluSF9B1S6mPXMrhUjDAEgrzunKjRiMza1F/un5
TTF1MlpeVAnal28KDqITeghWb7N2xLa55X1XVcuYcWSM+06tOLl+GMvCaH6NG5BS4UaI6deZYVHN
5CdzfVrAcQugHIzqUjHfRm2ovbgP7lWAgDlF4z8E2ksi2ZsCtbSqyHMaW/kHWzd6mJnNFK9dodQL
NmnRqWIBke4jeScGOHnSbTPmEPzHOUCGvWV6edMFPHYjQvohFLmXakMLxfkcyaagO6qGuYMougca
S/2ahT+U4TjDSrQF9FX/3YdvKPBa1d6GSlDjXSkIljVtb8/7r+Dxggq5PlYsMvN4tlNagDRoZdw+
rkaRTScS4JX5Z4Va5Fq87FJMv1T8D/XlNNxYuHk6g16o7Hvh6MjDINEAXpD4ZJnQTen6QlYRGrko
rPBtBtdZgkKxbS59eBuXYf/JUa07dPr1gVmASCSPFtEfxDOoCTcYJdA0P9APCkFroPNJVTxReimq
mHVIKgJcMzbSOmKXo8L6cno3r/VgkyZbmGigYljrlsVOL84TFUsxvzELo2Gr6yAttwoKpsmOn2iP
d6UW1FjsL1Oj070246I8Gpr82XvfDJH7G5kmCARqW6haqTOvpK7qWKYp3+SFsNFcnMzHD1BAOMfR
6SWUhvJFc7tOnPXSFqUmLm+xlZpn8XSOMqsfW0QW2+vNm/6pKpE56a84UrJej1JeDfYNJZmHnmHY
vmvbyJSwCq0P789zyh5fydN4oOW/kIwntsRShP+gxHUu2P5cw5Cg4eY2vQf62vYJ/XJT+sc7C+2q
659Cv/WhkK/w9TDSOAazrm1KLeO3bZYSi92RKxS+C571HwXLlOUTfdfDhumR51PAn3BZQF1uclzA
SXAF4UyOLQL9bfu4a4jvlzDmqQHQWR4AwUx7dRXUrkqGODLaRC+qt0Y7NmhNQT+MD0B1Bnr7BBO3
jb/baIPkLhF4Q9X6yN9dEjrq1xtmwVBa+amg77TItDwmeSs77XPzL3+nGXwn4u5P1lCqPnz/KLts
jE3TFIMehl6Zswwzh9jVaa5HuoOpD2gU7aVSPFwJ+WIX5Bc7bN5mSS2x1Mf6IJ6pHwF/Pm1qPE47
BZKBKWufT/oxYavqfDbIm9PTBbLSw3IKWmJgKIXQbHZtOlOj8eRC0Q0p/dJX7tfdNklggV0XtKu7
xLtJHpCLBQVb/6wBZErjGs5djWeIIxtL4D/0aL2f8LCHQTx4WYrM+7FYD9ifEJCFj87cXkz09m0G
VrAgT+v2FyphDGHwyEEbxwj6h8wRdqJz+1IQea7gwvbJvQYXsSHop3fzCIiXBrYneHML29vfqP/4
4YM3XhyHVdUqwzrkKO/ZlBJJfdGS8UtwV/mFG819yALi+u3p45xGAMqv3wcYdSXxOTQaqTLoJ9BX
WuxeXgmyzcO+lN2h4S7gphhn9TavPSqeCUm/kVg9TG4U+At8J1M88eN0k9UeJi/d8pVFB9gU3ai0
Cfpe36EcDn86cvHbcC+n8lSpss1JX1eWMLjd5ahCKpatlslhJolQ/3CeD62lCKD+164EPnPdPu+o
fsT4h13Xf1F2D+9IrSFJgfo26+LMtR7G6pRBaC0YO0hkek6lGVcdnF3dmoKpkaLBjdO9UHK6irbP
ct2zMNFzr5w5gbQAKR7IWv9eHsZiVTu5esVXPOk+aW/2zna8vFJczoo5UUYNt1Nwx8Kpiu9XuOVW
UEyN+58oJ+RANIbMB5zXT1fBaF2HOmZj1zskOnXRTXxRRqzWZRSfMIi9B5iVQtFzNAV3/iaEdYSD
0xUdmWF4HZLbN01wKG6nrKb8juvsnECTTfT66FnPMLqr5ZSn/MIEozrZS3AHqM9YsVBZg+RjC6ba
vJXfGgE7U6Tg/7ViytpfJh9swUI78AUWnKsVGXIOsV03d3BfCeNQZNCbg6AtaxcZfV2rzMugslt0
mIhgvqvK2h7oT1n36FP92Ssuavnt+0EEbOBUbnGV6dm7H/aYivBEKk/+gA7g2K25BzeMfZlLZgk/
2llz57ByLnpwcx4F5HwZfLvV/nnM1Y9EMsKlj+6o1XhztROLv3TomT2+t967jO7KCdsE/ynToy0k
IZvVMFCtX1L3Qwy4c3O27IF7thtOcguy0Xg7CxUV/T+pboKo4un2ZO/b9mDackSnBgNr7HZT+F4B
Vs3HUvirTkm9nv9znwhtdNCF3v+5TganSt4v+D2YiLTreTfs7GpPOaIF5Uq1u3tDvZtxKgMqAe4e
Et1cf2K8XPpqiyWbSS058ZtQxyTdUG30sesR7CFoTRCjGBhnsyAZoDzzjX1UyLrl/RlXjKeqlb/T
DttMWCDGYEOTFevc7s1ZtOQaQhmPisVEUKEYPHv1y+sB3dDybsTUnKZLQCSscHQtLa+Tp6Sh5i3B
giLqoggax00UDoVtiBEB8Ors+okZyNZg2owj0/Q5fiHAg+aFkUedi1scXhfr8k0qL/FX6MWiJWJ3
Z7bhztYZmeKFmMarelZsWANZ3QW2wGJyIZyXeJyP7nvgGVFiPIllGUgwx984zxi3ngamQOp0TRJx
qH69pvbNvyRA2oZg1NkzJs61uisBKHgVy6nm29rGC1Xs+HRxjS81ZU034+OfJJrPSOUbZpLd/23H
hrLgCrJbY9W176C8DsY4kM0GsM4Z81OUOMEbbDn8BHFo/9VfuV4+GNU3WvcDIV/ilcFmAIXmU6S9
kuWG7n/czQ6LDuES85gcfIGuLaTyIGI1P9fVQ0wwEVZ0aDVtO4WSCRwf8zUddZXkY/wAeGGEiGhG
R4MYouW16tZO0gE1p5VsYCuGPlKSnKxVFxG19L6SCjIIH9ObEBUxmwULED7Q9TsFQT4k2gEcXkmK
Vhp2zYrGiA1toJbhxlwYAtVlfeJbSb6fJrs/28J4CE0H6lQf8UWt+XHvEp6wd9jwNkqA6ELJPN0c
H88oRkB99kxqYzxgbPtRBQ0USgd58yxt/R2yCw0gtcH7RQnOWuWZvmrJHsmVUP1HOc5gi10Mp3of
uwgQAEKrJ5gtAc0I2FGKVdib8TEj4vQxIgVQW/BhEzIvVjzYlmXqw2wi0rXafPnqXFjLfRuCVmeE
yMDof/vTPQ3NjDmho5c2dfOu4O0+sQnjI/CgtYVF0jK3OREfageNzLHjgyKmKu28ER3f6x63o29O
Z3KRpmuq9apHhS5tKLGUMr7ZgbudUP3JPOJerWJuL1+PFfOoleh9GFkvENGbR7uwsYQ28fnJStdg
Ot8SCfFTA0jTpvP35fYMKqqxyH9svtXz5cxlm6KPw/A+/sX24kZHer6fs+pSOa4CLIdBlFvZR7w7
1VtmK2WCW7OvR8Hyetu1Zd4HHluLMs80tFriIASLamjFxhceqHRbCMqXl7kbrxd/cY7r+R574q6I
Hx4RGPMMWSBX/5LFmkGhFAsPBac1hPKF8+Z1CVmZdFpmrxMQmWorTSe5TGCnxKUGr2pHBGYHIWVA
uc3vSr+xcmRgkm7C0DDCd+iXbKUfWdyqHBypHt20qqSdufh3IHhaEJHAfln+H49+HHk9azet7X5J
PAT5zjPFoCYOlXrYZKrAOtStxBsNtwsQ7je2aKzqtRKEAtdExA4KfJdi4ygAQ/dcGEIey1hGljVJ
JJw+wGW3m3IRPq4Gqz8p8Pl3FwRtTWy4A6PHkanSF5rl4ZH6Ae4lXpbCC9hycDVgxKTzxLeGulQd
yGmdCIkomXjOYqOw/1TYaZuaZSbGoPEe5zT4YTORcBTgJG4k7ZB1Pgu7trlaC5hmx6Mat5eJiuHl
Yb5eEXLGIcpvCGQ7LN14FidYV2RjYrN3AMDSNZxfQzvdvxNgDGmkwTUT+ePG1mx1/bs4n8ubFduZ
Atis9B9GSyzoKoST8kZeZNnXCzhUzIz+FcrXV7yjGRNCbsAI4Fcm9+CmFZ3l44Q0o6XT4snwoCSh
jm5WXoq2zAf31nZGVVEjUEwKy5CWmM1Eu32sxYyAa3rI2aq9DamTVG9U5D3tvew7pa/RImGxDDer
qg35fqP6MkYsrjJCSfp/MOG4T+2oeBDf1auVwexEVsUCmotQuNZLaXf0PE8fFgVx2SGyMd2J7Xf4
Mb2j7tvtOkuBPRVhlJTF4+91vohJvmM3XbFmjiAMW7fIenRy5N50fAbKl/02mn/wy5NdM2UBd6g/
3pDjc7XCCCABw0S8mouzOrohgqvz6oFgpoke4gN0q7WERp4yVab6108qjmxjSX7blpW2X63WbKMG
8GuSB84N03gZukUgLb//ZHjSqQ4VbCfRE8uumbiWsRg9trveWcJiRCOi+KYmCWZrFfqwDNLK1HdW
2VIvM4HxPQNjNWG6TKeXGdye2eOnHf3KAeudJUWOuY541VCsrhJCqxlxKPj2YPuRQ6ZvGjLhMprP
OhEIwMbeQWBzZII3IOVpehbBBpJLBEMZtTosRXNcJIKy6/bH2ieZe+nEf8cS0brX5xw/h5BV+0en
spo+1M8gCEi36G/4Hkrtgv87c1R9tM5VeVZZxjuGEX9JxMe3d7Rcbjxc9HvjW0JQb074TKyBshHa
MKEHw8FAbLWAU1PfsqzbsnEgBWGw6a/QmUtP4e3YfKFrQTVdZOUHqMFxJ8GFkcVTlwsXWfxK+2j5
j6xPBagA0Y6bFrM9D/uGgN8Nkv9TCo/divafyZfoy/wcBZVJ0bi75BFxLA/HU/U6ywLkbi4+pH38
XRXDYnj5aoM+nwbVkCp8QCDrDBqz1/h1YwafIqnp+H/3kUnukkwIEeO/Qw3PrUVxqEMTXdwjhaSU
VtLGYAVYGALLOcji4cNpucOpvgyl6hYOLLBuMYe39FyOnP/GRNDC6w1UQBas8XW5hGZjoIk8RVfb
2rQS/HYC5zpSC5TjLMPWWD3xS5rNnQBtgdwa1Nq+zRHELXuw8rTDRCxDcuuGYnzB/wVKm+SMqHtk
HU5MqXqgMeLqu3ruBl0hbWTGgtfHBBeJHf1vteaMz9VrKXxfyud5xg1NzBrs7I26D4pMIJzfBF5r
nWHAotxKnsvnvj6Du6G8Fxkq8EmAXY+Or2MVaxJzAjrfyJjs6eL40jQi7M/hZjCiMmsteOf4Bi3H
rJQe/NITb5B1V1iayWsvsfeo+6j5HbgeUssOFbhPUiUj4dv+WlSkd1C0lbg/b7Yeabu6TrRl8KZQ
dJt96nLXnzB//krJQRKaj1/N4TlCxSAJaRxnhhTpwvFCcvE=
`protect end_protected

