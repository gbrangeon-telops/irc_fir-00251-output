

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JEmZWuLCZazscYOT+xp8tQcgcJoo9xw+tt17VTk0Ee/cpOS713F8lYXKKz7qKA5t3FpvNSj+LwOT
FOkmwv2alA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IW+w81BdrtEdSrXT08IyeN9itdwHkCyvXK5q8xF0K0oVKDwJZ55f8rUD3UDvvDXIcAjvU+645JL4
ch4hQtC7Y2FokqIuMtHZi7cNrCDQXzP1bGPJjMCZbuYkodHhhDFZq0vnJHG5npJwjfiUcFOs/BD6
321VxRY2LE90m/fkP5w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mn15icVDdA3CjzJnkJvEX3d4TytP/AnBNj79QG+E3lCes2UF2pZhqISOBY2uufaQ44Iz0NeMSC9n
+tRGbjECz4+Qnwa3jPWzed02j/IF9RX7XCNKwHKcmJw/yHIa2jnhfXGycV+rW2BTSaOcvd71AX8c
xlCKhnyKdiYayGwfRy3hMXLuu2cdwaKnu/UJ1yLUb2SMopRlt3x1/DS/ujprioIUaznXnUPKvPI+
tY5o7OvS4nta5AxgAsVoz+HHq/K+cZ5D10lOXIDOatM1ESgBnEMFZa0ND/EVV3+YXn7orwuIkC9e
CVEV4WCQjR+/QOWg525B6zV97OAe2sVt80NsNA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3K+sUBRgBhLO7z4XKbbFj5Dm9dnCnLXJtz9DyutJQ/EYt7E+7VQGJ2l3bkkVJ8bn/YxKZD+Rqqzl
gzUxIUqSuvPPGmd3z16szdtLqj5YRAEZVXdNbeQ6P/rYfI4kn/0Qw+0hS8K2lRo5EQLrCely7fSf
ojGqs698Kv3dVxOM2uU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EHFOd5L9tY2zUSTwaEQFpNSik2aT5WpldK4px9GxR5cWZzjNzosBm4ckg29GsE3hW7YJVXJwn2ft
qvaRBZQhqD+DF8s0vynZ8IngOkOgp968BazD+XmnNms7D3n8pwwWq1DBwFf103zHNgk183z41Fww
ghnhfPrVLnkJtKMArkX+0VsxpoDgdODsv3fsT7CkMz19ja8WwHPQXCAKUD3p2rptjKIU1LKJfHEW
xgEccgVmdaHJ8o7kwvdgJQxZnf2Fl62jKVF8AJCrqXWKtvakZCxpEqbYNpoJ6R3Ns/YvtWdsZkRH
TW3+uPSDGYDVS3Az7zcuFIC462DOhpyBpwOGGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31872)
`protect data_block
HxUgl2Y5IrqHkGfOOFe8JdHr+xIc2BYoOJVoLBrCAA+svGl0CDm/WQ7fQLnwfLnPJYf77kRja9PK
TWcGXvQFd2hwkAw3V3/2vk9MNwxWn4IzGc1GnqFgjf92cDlK6ZbawcY/WCEtTYsRSEmsbvQbzluk
F5oAtDXCUK8C2G1Xkw2RP4SVE4O13KurSmrzADMhg64ZOVP8uBHdjXA20x+rN39t3V8QkXtnsPeE
dDgE/eGjbjdSk1gCSkGVS6EUR89iw0DjjjsxWiebpx7lqIEVMvi02j5hEsnREkbF2YduQcG5Svu4
+MgOYCAqLRwgiUP5NbxGc6Zzmk/sj1TZRzxOR/+yFWpRzWECuDHph9eFMKwjFJbNSCXJRUgNEefc
geLGon3yd78FXoYtful0jU7Y86vjNBDHaYSbmQU6FGo7nrqCKAxMI3uhhIoV1tsKXKULPUQDTs4f
RDAMlcFrzjzCyue/a5/ZFMCocum1KwD8BN2lr2gWLELoli8d2XChApxCgovek1T6RgwfeOUEK2Jq
7vGh1t5UigtOuEISMcDiRQJo+N+RnefBaqEg0tpA0SK9G46ymHZ+0DaxY248ou9bYQ346nrdMvy3
mUjjL66mXeyeOgFAf0jArSkYRMuS5aKcIuavjhTjUV3HZg6bqTb9N3b6GLa9AEn9BbZjL6jHQrqx
/ODGXYCJ3CCP8A4jfddhHf48E42mhhBXyXVX/X88Y7LK5NUIV+icTt/ImNavpfiitkVQC91O5+BA
9XwQyccZ4kPAELMfRutWungSi5BZUqrZPTXOrII0N35VxCs3n2YlwwU4f0yLYzWrAqBV67wkKjci
VlWVSMiww4LcTmcI/5BTzHQU53pkA8TQXUdrsgtxGUcDjqL9m6YVi6FU78JjwijBA9SFZb8TKI+Z
FVlUhk2gNQ6snlm4VhKnQ/yWmVp6l+7Nnj/6vQFcIjRq8nSWAjyQspCgh13kqvuUnsjXOmdHwpu+
FGJQJHgmWZjAjKr3t0Q7NEEASa3Soua/UUmFp8RwBkLmmpSOrGX223ShDxV/lDEZq8d85zaHgUpo
uPtQ1fSgegJxvzYWibTGGb2D4bffbmNXA3kEk8k5qi8QYHW2ALaAh0hK6vb/5mjndebMh1wXprSw
aj8XvNS9JZOHlvw5f/9XGW0c+LFdAp1JQt5Zx8JmjslTml/nBQT89DL9Dl0t136xmKf/f+ryZ41Y
DNHV4y7rWeNOyruHPpbIW66EJWhaBFr4pnEgx65GWTOXfoei5yk3aFHJ/V8d6qOmPRwHYuKF9sY6
OC/QJgfbtmaSWwcuXQs0cIvV3tDsC1lpREo/qBshUi1hi2nys7V2d+yHa/m8CiQg4qZh3f3Ec4Q1
kqFHx6XBy1i53H+ZXPMMBR3fpTHepwWihBvanl3Ez2ynhGpMzb7oR8LI4LKepwNrn/8lHdV+8DKI
TwAbznt4+SubOk/T1KuqbNY4XM1/vqXzXR2h45tM/JHhhSpzelTNcK0MD6LgPjkVhJS4ju1i0xV0
m5i7+ED2DUhbPdWFyx2ZvondH2KWGPmUEQCoujqyrWJ0WMMNtrciOEIwI5es3DWLt8Xn91zsnSWg
Hp0DbG9nZBx8TOvQza1OF1uhGLxCEWUxRSCRs2VuxlTxoRhZDPn2MwmZ5ZNba7Tcn3aKExEHj5S0
oSLwGNebRfOZe1AaID7ses7dB32YEbV9dkY5sWv2xNXDLZDhk7RE/qU94sJwUCSr3gwPmZL/cZki
5GJv+m8G27puoPknObYzEQpdM+vVGpTDmwPr2y/5MOQhoF4JSigba56DfzwAevZUHLI8vufDbhdh
rNBK2aiO2/zPfqh3s+t87uYlnHeFeJLtNnJvPUQhpaGcnQf61jMi073PJeUGOJnsH50JI+rDn+mP
RhKd8ZOBqM4us7QEvoXwh/Lt0UvD4KYHDV1USU1amB5n0+WnnyqOw59JpcTf7xiJRBSIESVmZRk7
xX1+aXPhXeWyR5BQ079Cppfwu3hGuD93gt08WasxG/rvCgtCL8vMjWqUpOqtC6alF+SBWVcWjaUe
9TeKQDfKV3WIAmLozmUbiB465CqZfrMk1FBdlYq0TXSGWXHBtajzvu855ICRKSdGpIygbRxj7iDZ
LuH91gR6zv0hZmGBtJ9N4LK7DHRrv0fwGwUj9QKQJZOljCb9SXJ4pJBJVDiO3jZBLsBw1wS08dZ5
nJjhL+lfLzhn5kyGWfwUWc1VuqZYhlg/LH5pYiPGnAkV/6zbJAShnaK895IkaUr0hgAxN3cTnVjE
BsMbAns5h1tqk4nCPei3NWusTaOn/dqguRJL1egleOZ5CbOiWxrJ2TESX/abc7qv8SBeOtX8bx05
VJZJ+b7GhHg0OMqgjJL/EjtNFJ+a6jrc3+A33D/vJ7wLuwLCrIwUBFVU4SSOT9XEtBUdSJpzsuLp
2BXGMhujHEXlu+mpvCdBDErnD2Q1QzskeiYWX5FDI4K2ud9p7MTI7QFfX2aGCc1KPEsEbZYKMQmn
7MY8ZazLzyMsKDrYJLaV55DwPTDCUP+9lCGnG0VqregdxYW/WXaKxug49tHpY6USsdScTIv4DV0p
7rxKuEONLNmXjWNkKHVlhzJ3ESOZswDxl5IyDtP2MapOtjmaoAx9gwbwDNDcCpQYH/ImxIt1ejsf
2A8nzIFTU6rk3fpdZJiS1nww+pxZfwkU6YlwTpmOXHp6KMXtCXbq/RHtvecevorou7faC3QAsflO
BeUvhnR7CWZ2xgdoEeHlqQw+sW4d+B4QKXKFUnhz/hkeh0Q7SiSVPxSfCtQKy1ymsnymh+UzaEbf
lYR15dLsLzvIxWB1+Jc6FqkvHAzxCt0+D6QaCFBxlJM1zsjVSUWWHIT9ocKoWtzDKPm9mIss+CkC
Z+2FEViikRG7zGGYo2JYxxDeCaX9uNexb1rrDz3qrnQAJSshLF6CzSvreUD4S1Cnf+Is8taaRd7T
FXcoaYhn31VQDlHg5sh4K/RfH9blh0AVsW2GfRBSld7e6LMCETGA9yfg7B9AiV8JmUtWJtXji6jj
OudyDO8yoVWxP+15pCSsUTodxZ7tZ2H2AsvJCmvggBDEb3AAVWf+XbdWG32QbyD0mXBveMRK5MOD
FZgmU4Gu2TcLgtebG3Ap/u/ox0jRSSRflOWRxxyH0fetSSMkm/IetkLWQsS1AdY11gJlNU+wS1tX
etzOBfNbc9j3m5AyG+zkkyKAwxJEN9xr9rQSVKFw4fphmCh99Vc2O7vQ0YuSZ82o/1245benQB/h
KMRm+4mjPvPH3B8DWE2MVZvO6JU17Tax+qRhXauICfYcK3Dc503pX5ZsgsBQ0GeiHIAZ2Fjq5fyV
e+xV2f3vYsqqP/94Giaa78NDBV/RhgGN74JCMaG31XBmMeQhQXf/01st32Tdd9grpCxNFmrH6NAU
4jMEndm2j0p+I0JzeX3poPFDdp6P5JieQdQ4faHRJ5ayqPJ7X1SVYQNtuDMfbv0TwSnrzAF9zb2r
b7IV72Ctxa7Nm79nw+/MkQbE9YhEjs4dQw4uCUoR3A9Y81fqbPu7r1QRQvxzeLrZgpRL0dPK4ToK
TS4pEe7Mnt0iI2pdCYwYESXy30GmggxNS3fH27Lw9+smUD8KMHGpoSJofhdFk8ZkdyDfisfE6ZIf
HYNtpQnzpr2eATy2MRVN87/yXAjaAJkjBWUgG1fesLk9BEiQs/WoAaIws4anw8ASN98PXVKTHMDD
Onn0uYcNhuEUhgFPtUm0FkWe7dnxjhxg66v+/eqpo5cV/IejVUCekVdhM8pQL1qsK+9gIBT1ZtkZ
6P9b7awphL1tFVLLeUCEzvES/k7URMxhhHUTpTVppPeOmVz5x3qx+MsZDFlnKgIDP/2e+oUTuETW
cS1G9Q2W/v3iX/tcGRF2qLECDN9LEKGqqVtfrble+vt5ozwgDrLnSWRcQnLddEVFmW/7m1hr6Oda
MfSjn3ee963iUZ+uE1C8rrm7faBXke7LXqYRmPFKCnENtUzWxh6mMhN+hhBEo4P/BQB5qoOg3rEc
uFDAgwM0fNm/lEkgLYvpfWPUiNzM7IZCBecX058Ifak/kSSm6e1ByLrv6eb/p49Ui4OeATid4ag2
0vndl7gUlTSXchzClQZA2vlL1jdqMHuos0iG9sKOI/AulL6B0iRrHncXaEhepFhBUBPgWdlquJvR
ePNgBTve/UyodAzza6h+K0Uzt0Rif2MjNlOYKv5xLv7a2oemmAPn4HpFzKDWAJTOQ/fXxtYbax45
SC4pwORA4vxpHliRPkV+NKqbOzbJ3MzElroqAjvvJWLP2I1IVL1stiAsA/80aZl1QHViUi3LRWFC
ubc6pWcfc2pmVlyoNBc+Z14O017DO2/FUMUKh26FXMX8e9tlrGDtvduxXBqmKGP+42cTEiIbJsBU
EjbjSHc92+fcwl3DVJ2HscAWXxur0XpMzh2AzdFUx/0qUsqPeafH0D8nOJ0JiWP721RzSwLZhtCP
zQ8qit8AYXbTuN8EdgW0yYAIrcnMamFNuqE/YeD9kKLv8M1YVGvUAoFtx93yC2g9HmWzrNqy+NzZ
Ak/L3+9f6gHesP1EposEqHzZfTqSpSa/oQFNRmb0CfdjiXmHEUlL65d4JEzzrR/DX1N974Mu9XKV
lYArbnA4VOZfWzuSF1hP3EAjLL+KZUA6sD+5dHPUyfwokMOfl4IGinH9YbHyE57pKhLt8P2+jrRw
LDpc+Ou+3TVutMIotGf6zcru+EhfaQSx7+m+Ja+Vxt80hRwcfE5I8AvfueR4wTK7Xkop6HAQ6Jl1
tzbm9rkwWwipRAxCW2/W4s8xRl3dC/aD+zyBw1pGi5VF82rS150LMvmIcmPaIoc7LQ/7Fvz7WPMo
NUsCXrChm9SUMDAXjmSvPxCmQ0zHf45I/xaQrUK+IXGGmyA+xpfxtDWpnH6/YqHF/T2aHMapDM7y
aO8ysXTmkNBcYV/pAK1oQpD6IRh1Hg9tKzYWxJK0zX8Ev/D/XuHrWyG857/lm11mva8J1IJnLjeP
27JoEn9RT6Jo1paEBMNh0wvYjc/8tva0lm6DJyeC55t13vv0HMmiZ8M7rNYKiPVpuTKw60GGJgUX
9eW9TmmD/iLVphjfPRLQCWuV6FZVZt3DfPDBuY5WxB/7Nl0Qgmd1ymQ1JFjHfwqTUQIEB8J2qYIo
dMA7pqr8/Gl96Ux8RQeo/oh9yyE52rasew+skqSAgW28GMZLmoNE5+8bNxenXV3yAEgJcaebcqCM
4/GbmVyIVUAN7iTIjxXxqvL4hYZ4WezqXNM7bk1OMCBziQy13ENYaKvUXAUgUcDM1sD7BowWBuMA
G+gVurhOBhzkCWz37CxYPnMKkM9DhpB/xrFAsPfuHhiOETyPzPJDKiViE3W7oFkWUdlqrWy/q+Ab
Gn1KRVKSTtZ3fzjPYGom69uarY6IE67I7k4gEqfEaDdt9cVBoIs6M4m6jfqPf8nTNhwa3BQ+IcZ1
GJc4fp8P/JvdJR5gRTSL1uwVBR/S4UsEwTyXhPZ9JqJCHbu03Zs4Kvkex1kKp/hMcSP9ElTo12D8
ohv9kzvoSqtvmMvxND89k+ErBd5YVVVlOh7Tav3NUECq6Mnz4H8hpr+nGY/0goMs/ZKYI2sTsLRf
IQzghD+AGnOhoMPL/6UfF7Owv1E5UIDhHoixEhWn+hdv0yA5NlRCiqLqGqlAUibKj5t9wtiZ2n0B
AifBR+mQVHO5Bm60BRFXru2VB/v0u8tMB4cGKZFcWJepRP0JSevRdTKxxtsS9FUPM8qq+MCmtOsG
cbkkqdo9QfYx2yABYxVVsFyJmkIzVz9tjYWDlENjwFgiXww7t/vhujqNziid0H9LVb2PgcsCJhpz
i9zGx6mnV9yIIraV+LMPoU1OxQ7BE5zkyxg5a7HXpDiUxxkitWff5oyl/xWN94Rt4dCPalFFTJFd
2bi3Y/ailvEzSFRXpcLIzbzp+h3+Ckar7zQxNhUTHng6aalE0YmxhBfcEfqEMXQ3HJ7Fr1JPqt+E
jQ+7Xz/rh7wubI/hSOZJqQNW/OuMweqGMMQM4xf/fW8futCNYMnKozMiq9P0iQ+jYMXhBWkul6AB
fjJRCohQsKuGSQs+Aql5IGh82jl5kITlkcNmGr9EFexMn72lMOhrCn0XZuUi8rdl08LmwRe1S5Tm
TB/Vt/5X6TZsz0NazdfEGM1XKBKCgFDMh2DZxQvmJQ/HdEE/YpvcFgeR9r8HMas/Z8Dt0MsYrjE1
esya+842yYd83v7QsUgFLMif041XTDfhlHRQm8zI6i1feiq260QVfgU+0PABMR/EuuKHjgtAQck7
/rIeEhvWSSSK8KxzMt1Q2oyqykubeYa/8aa9C7R+WwxUhA9pom21dJxUb3qETkBXWUHUAsatXcqj
sgNgOLzXwA2L71Dgy2DLwQivWCdelOO+XJUt5NhfMNLn8rQciuvczBNnAyC4TVc/nBEGLllM/Yq7
If5/Ocx7UF6wwe/ker33ev+qIg6AlDZVtS+J0DSeHUpzB+nxrxLYZbq2nQN05yWbRyytYeAeEIYt
4lRJnU0Nmth16dpC18E462NgB4k79uHAW7M+bBqYmOs3cY42rrdlAGUEwAO0qACe/OgML7k2UvfU
dcD4zP0fj7jDRyUgyaVl01xFiXAjzLx4sO0HJtUpuRdgRCxm+Y78OF01P0f3JQ6TSLd2AKSK0/vK
bMFu4rAuuawnIgU0RpuwUt/fy6YIT4L1PLXsdnH5QlkIAKPQ66/rWe5qvLckpwq3lEHo5Jmzh2tJ
kxazHtD0FqKDIuRvxyPhvdeNlRhtAgY9qK0WAuJ6wR/VMbL9XzA6wvEZjfKjhgEXiSVocFqDEu6L
wB9+DwHlR5WlQGahObNQvd6QBzS/Q4SGMzfmJq1WcWRcmMjplqu6vXQMhhsWUqR+5ZX/CqNyL378
9x+HQ4oPkU/c9A4SNh19eVWuZjKZ+v2WyFr9/Y5B+7Hmbo+QuRMtW9zUOeLg4HQqdvrSgsvxTex0
N4msB9qRtTLMARE1xn5xRA1TtzAvf288vFHUVuF4F9istgDVaZ02wD09rRCoQyidHfCAgddkzv4+
x3vhZMjVCg0gnOiRafjEbJ1DdfwyC20uh6WJZ76ts0imK3R09esG9FH4gl0mTZIExdJCdPKQHP7p
NBgymoKqoMRFKx+8EYQTot3/gQVqe0wb+fN6y9RB2sNu8GAFGkL7zVWFha9muRyS1SnmoCQtmUhZ
TrAcbWzCMwPceI8N44qcTiGUB+j2QMmwAgwx3JdNl1V9coKUnKsmGqyqHtxnBCFblOjuBaYkeAAC
/28g0RSqHVvXtu8S5O6dijj2pra3IK2Xgj/eFHTMq15aICWeywz2Spux7R2Ib7irEPnOyfm2Q7Q9
MjwYJv9adkmZ6R7JlNareOEXTDHh9utPUHr5Mlvv3RQNhsavJQrHLnTedpIm5f15Hl1vvdK/tdMc
wamHDOTqGj5Y2/63eAxKOYW+2yw8C9fygJMOWd/g7e/e0mrzYNifNJICa7smCUzLM799/Nbl4GiF
Ey8dY9kk78vlV9kkQimw1Yw3zQFcNJcBDpXX9X8asNAnL2R0mQr4M1TDAiTvLgku2tQQywtJEJ9X
86rzrESwqzNXaPUDRzFoNkt5RWbC6MSSgiUyxGpqzyov6pYQMfwj8jFuRVZcbLyphUnPDvwCJTDr
RCg3i4XhEt+4kMRMtuZACMK7yDckiarcZQOG/gE0n4KTxt0YJlQ7JDptjG1GbId+9ipT1sqFkI6n
xyyVyhXUb+ay7/XZKBsf/nzJQoF1kXNdBePPGnht9+VWgYU1/MIMAiI/jjYliEZAYQaewl3WNvca
8ABZ9HOl78ejTK1Nim6zCv1Vl/x6SXHAruMR9YL9/eQaq9OYFyIVgx6dmajX5vseqT7pSONvrI7r
erymhJAcBFaiPl/I0QjIL0QPNFemMKPtGFgNEh8z3LTkLu1v7fTDHFBBQ9RLsZjurDlTHaRWPFxY
VZpRD4KHyEh31bvJios0lNsRx2xUhMqHtP7T6q1mtmDYImgWnJtP2NvYlLHYodlrN2H1Y1Qbyp5v
xqxByjvYontofD/KlH27QAlcUB6w9OCxc5KBLzuLCw5G/lQdNU4GiW3x6z8Y9Qk+zf7NrtoWb7cx
huefuHDNVzg4Bh5zZDpYmvDb0fImo2iNfzaLbHOCPaNG5Em2HdyLQ/WVW70y/D/unLRvxeiO2Z9o
x8nB53xoS8ATfFVcQv5HFWf0Ze1UnM0zN/LvaVL4i0LNPaa49XVLNrs1ZG+WeHjkwFaTTL1WYxwP
JmrhwP6XS+VQ8LNbykyQSM0nayT4WIXOjoctVqiPeZxxxowWoBa+Tze4rzMTncav55K7ZU8/GpTi
jfhD6mSxdqKJlAGsm1bFjz8bxffLlmjzXrRFL2ueLn3X7neRnBwLu4E7fYbfM8u0etuEN/ZXbsXI
L3uEXosZkeML75NO9ekqXq9+f6Qv8y+bVf8tRZk0sxLvBZGmao0yPLRPkZqy82jknePE6dIHmre2
E9YUxEWRZYYT+xDC1PlCbrY3Y92eBz4x7HmaWw8cpZmbh2z3Jr9+pRXjJm8mg9vZX6VUvkLlxxoF
Ei8Yy3UqiVopCFEM5jleMYrG5XHhwWEXUyl82QkIC6uYypHRgmsylv30vNsyYq11xfPX5ts9BAGh
rBbuL1/7HxHlWya5mHSoRgYnDD1Q1Ak43R6O0ZHP60lm7ru2Zuvqtq8SaZ5p/ZpqAEWUo2+r69ZB
uMoavGiww5byH7xu9qV60S94y++9qjXUp6Wj72edjIWJxDiXge2mEhXXThckxxMbFFEsgaf4jLFw
vM4/NLChD1Fh9Fw24n5wqgqDRIt4/FEiEyC5UpixE5jV9iEX8eFsnXcnrKx6SAKyl2EKuGGGrd4/
yWO9Zf2eNFa7VOT0tVUZP9y5sDragRp+/MEauJ/Duq1ddgsm4zAE9uE7USr2Y6fIqUDF+hdVOPTb
gDHrqIJWxwqJxlq1XHBP0zP7l1cKwBs2zX5UZnHHW9hNuY5bh/YV5rW60Nrq4JXMwBRkufrVhaGc
uCYtPy80MhwNzt3vjtMW932zKP04f2HaVFO9lgESbj8A6xu7qH8LFI7zc1RAUy0/lrvy7JpRkqmZ
yNJ8TkG3hnj+yjFxTeQLiLdrfSqvzaCWCTB/gxFeNn+YuU7+q61VbTLJrcO6hisQgmjPPEAuEyrE
VHYB7qyy0J2Prak0J7Jjz8FjGoDGO4x73Zsb9prlbaaVVg9dhRML3dlr7rvnYCM95tcy0w5/RQdH
QTd6YwpFqzjoCBFzHhgSUQh2MWTgBdpAjeJU7eS6NqDChS7R5YvR81QCWm6iDtG3+QeDu9bjT2eQ
O3kNLdQt15LaZoH4un+xiNBqbIy1UFiTz2vLvLtkciz5p6tXV+omdgZTqNT3kIjNAQrmX910dvHN
Wf4y6yFyEha+/FBoX3ESIQum39k8g1gPDLTJ6PcG/7zdW9oxuDdQRSB/AOpUoXmEB6cskoE8iyCF
vhUD2VzIzRjcNGWzfvzptK/M1p6smbEnihD5uLgfHBtktIq/onjbKQEcI+nRsLxa8OWQBn3+oqxY
tqVLJH0zjRbac2JUB9ckaqwUbOZHXYNgvXfTdC7Alj9uUCqUEIFH9RDJqLcd4Kmgv5W+kfLTVRw5
7K5j26BHx7naGbVNjCHfPYa5I5YAuOryfjLQ/ATAf/MDs3I8Sn9FeAKIKheVI4BCWGoIjzINlz9d
ckz2CzRMxiJNCzwtwdLtWA1SQEMZT1IWz0Q9M82n2V4gffWQZUSipx7gM7ai3SQqd1JY6lNuO8ij
Vn5f0+A7RBhL6x6Y3pvJgawbshJX4/JpKD7IKi1GRAOtZpQZjFt+ETMJvR7Vn7bYHiLtAwZVxo5q
/T+SfnLzfGZMkHGK1BsQH36T7JBArxOSsHzEKHA+mLBFFoC1Fh94JRblmLmx7ztxRyUVbLccIudp
3AP86JRuNR5uWSFe29mSoBLzn6XIehdwgi0g0d/oFqeqwDV+PyDJDfv3+fTBjAB/fXMyXpu7YWMm
6znO33dBp8dQEYq6rpa00M+DqwcZ0beQROyYPb2Pi/H6ic1cIcVurbmdophY0HQyQkpG0k6CEy9a
PUjehfUKtwHUOEGWjCyqqHSAXSvDOE+EhzQk2880aUJuj+NDI2FQqDspoic867YKrFA8leblJ8pJ
EeHaUEZzzdEkuPIr2Z0KNeYRf6SV36izy3ZtrtfcjbwdiI1qxMrRfKcV2RCMLBoY/xlEAJxsj0PM
PZ+N+ajHt/mzNQpu3cpATT+IDLWylOpHlWUuRpUfHKkF3a9chVxultpgrIKM6syA/O6FlnyuI6X8
wbUEsi2FA9Jp2fgfoLCAda4T39mnxbP/jxotDxzdcYqT16Na6zBVBQK/h560XBdts1f7JZH0U79Q
d3bWHFpJZTmj9fSFHQmhizsWY9GWbsP2f6DIcZt5KRTc4H+64/MZgtqbZWvs0IXFYjjy6+tbYyCe
8+YhAFf0Iokzvix/0bEpkzuswdFxEBrHZiPgGlGGaTLLRBN5g//azUGLatnihpp3aSJxXSMPmfBU
EIrF+11MOoy6LCiJI3d1QulsbINrZ7PO4vDWTfnS1jGQPKtmApn+k0JpepNiRo0uDxjsf/zHLVys
askctt17rGbQXegh4KJzNEX7F50N8G7VXSPfpKVoigSKAMcrAUstI+aSxQ4lkloX8mR44TgRudds
impImr+9PU+ZRj9/lHroPIXj2cf2fBUaA7ubXJXWCSiM5rnrn8zIIK43/rH0UOvv8LmPtauEisaN
reuC5tU8jORuJ0LICyd3fHpqIj5Aadnslz8TsqeR+mD8pGB+K1Me8fbdMLZulNxJ4FkBlq7XgKXM
vk/37zlLU9Q1rUeFR5j2Iyhd1wm2Dx/pWF2E5zPrXXNnLA6QEeNUmXzYwjT6tSqT0YIwA3/3CZqM
9JKoAK47SJochhDjQ40b2CYAwWDMvORLBtcwqAedRflMKwhZ9wF4UGAkszBBP5zcoV+wkHU3zijU
er0hx9Dw3Ud2syceKOrlywuX1xvLCBaq+o5vbArQiOoyZBFVKah6DGjQgvoRSO9KyGzMrSaCjjbv
7W5svq9XGfQZopFcMZCJeO+1evEzgJnQndiCr9fQe+DdqgNKxF3BhuPJOVw/xbBAbIAgzK8U8k4m
lCxereZr/ldqBNR2PEAiu4WwzkyHZTfthGTMKuzkmMNI7as1wgyEKGXh6jpoQPdGxK/0FZj9ZmOP
1572LbPVhT7EYuTBmaFWlIrucPDq16qQstVrQIbjQA0ujzj6kLIFtF1HFX/vQSv0MTeDlRZ9SGhZ
O3dABHogl4umigQE3P13c2BdVWPAQROSTme3fegBF359vWZ+KGvzT6kk5IPxbDYAOt/Y5v48Bv5m
X5x33sNKkSBGMclfdI9TkgjHzubGjW+kTQkhPU/TCT2qa4+jmQJJkiLLoVbieTBcFLLsEneJRtMf
pbbKRbESp/z4acOGdXIF189QuLsHNSAi1nbPRPyaWm4S4+9gwxMoTNX8zIF6gpNHvTO4CVzHOPkT
r1fONGU8mJtNcDwM4D5ajRDWQaLD+Efl1GXSofaZgwTVYUr+8hqinpG63KHFSapNqcNbMMFd4c77
SpJGokj6Typ8YI7ZyMcJ8aOd7wLm6VQOlFTkV4r4IT7Gdv2MHoX4Egreq8cp4ExzZSsn5uAO1bwJ
XgINH4WfA6x5aRzSHN17bEVjagsRSxHbLRhBNQd4Oua2nlrS1S1+SbEIQJhTTfwkmpZYbY2bipmY
+P67HJ9Uy6NId2TQDLO02bs4Mxa04mKVJ09ZG8f2EFelYfSxJg/U5wLrTUg3/Y1W01x3Xm8kBCaZ
aLEB5z8Kln6Mb8LqxVLNsZLtYjX+VeYi/4QVGhXXEr71dEDPtttwloHxce1EXv+039NsyXg6BBTR
T6pySVHDsxSQjhgM88pKN36U/urOXG2+7jYv2Lh4qETiif4aQ9g5Bi3/CDhkm8YvD4JwqXAzK3Af
jqkg+wWik3DblSuvCTGPAVd9fEBsAHQeVajIhB7Re3H0Ni/bm2+Hwu9IV+HILOM3nCAXXHv9Lsnt
Sqp/7ThiXpBGWKxlo4NS+4Sut5TJqAoda6Y8hVMDFqdx3zhlSFTTp4/uGjTYKr3ZZt/ddnV1dX0w
bL0P1BLgPD/l38X3K5bk2inWwXhIO5YEHnuPxBOB9OGLo+7FCsNhV9h/2ICbczxYET3nqe0S2unT
4K/kJa7R73x5VpswXS4iusCTA368sZSZz3dmu+sQhUG5NLTnVVI/MlMi9YYJ6uUIB9PgB0+uVFhw
nk3iYyY1sclGaPKYeWhFyYa+JgB+MoeJ1Ua3WeKu5YDcDiNjGEB2kXHSLQz2aRMzLoDSwUaayyPh
azgeyaQdBSVNMN2KbfL2vPal19PVCoUIOXXctQUQZOgSbkxBfysVgaKDz7nshunxflCDoj5z2/Cb
TJbSlP5/vSRg+KPuaUoNf155rajqPKI11Yy/W7TeZCtbcf/SzXYu5wsa0nCCtz1j8QvqJimD0K2b
37FVki2OTJza3Dmv+96Y6TIhFApukrpeYn+iv8JulxVh1X21/afI++c+5DCUKYOuABVAzMDd6Oc6
gEiSQOGl3YMwiIzFEjhckeuJAOKdhdZzNjwrVje6+Wugp7PTGSZWX31b2IqvHdTyfLBBX+T1v33R
W6bKcZGobGL8ZmAqHE6t1JQk733bFLJpZCxCy7in2/HltjOor5mtgiGHjOKpAGPkStnvdEwaPLKB
NdkD2R0CR4EUH1L5RL+fqvmf64yD59JRBoslEPaMP3kBO9i4K37hiNAo/rKFYeBYnICE3TOw3e9G
QpPIrSSkQWPRgzS89ct5air+d+JW/DYR/9T62mcAHvCZ+eRxxH6IJkhdyh9FacHNrDGj0iH6E3u6
9vyjGvfjIDqU/Kd6v+ecRnebDFcDdhdAcizHy+0CYVgNKo6DnXuwBMYsBYV3MD4VNElkxEga5oK2
P7V+p4TG9V5bIGNJ3wADDSpvzWJg+dZW4i4wUbNlzRlKZ0m8q1T6qgAPF/0ODm0kAHKsSUfngp/y
u0jCnUv++6OeiB6WdLYiMdH20a6da6lOVN3WOIKjSTrU1jfIhtVLZIZFv2DhYbm5anao1TOTWdvq
0vD6NGPx9UiH/qDmxRMVAqsT294t+2qecPV77pxCq25vZffpeFaIWq+XKnXfLUD0TZNtO5f0o5pB
ynvPB7u+isfJLN1wOoqXT8YQIeS7tbOLsjmYmrNo957yggQem1b7WnddMGpgh2KVQ7aRvara8oZJ
k3gytzlbnV+s/O0tKO9ynd2QdyN6PF5PaLeXpqKVkSlE42F1wgv7PhtdjV5WIFLbfYo4HG+7zvhH
975wYkpcxRg/VKKiyt6TsOVPkabGJ3XODxYCSTkrLoxEBxgLBk9RL69BQ8AV1A58Q+iFduJu0T2W
U+zTJbC0Q/Zh9+Ua6CNVSX6DhpabfBo4a1+L/734UmASM6/YLshs1+rF4Brmr5tIZUvhCOlJTQ7O
bUCrKwadyPiEmHE/SwXEdh1lxGw03MsDId3CD114ii2+4oJKvtnFu57WjJUN/anm5PfiMZWi12tg
QF4ANGZ64EVyz612G8uV9LB+w7ibZN6GRCVvnPs6nov4AUdPlaLKiQJm1c7LbQMq4TG+DzlMbT/Z
cYakURz+mepKtaf3Iuz4fP6SNOFra0T1as8SnLDMkyWCIsYWBOMI7coSGcMTSTbN+f4m2qmwqIQO
NLb/auG1LBg2BNfjCNx5yfKSQsDzml7f4lY1z1yHq/kHQzvPjz//JtvfIbV0M12UPDKiweSQbc4K
WCerzZN+v2wb0trNUzohZ15n+Bw+ngF61CgqkxZbYSCbdXbO9gh8WVCB2FeV0fFHX44zUQWFq/z2
rUaeUw/0McmIbFwshxDzsVJYpwLBwjTDTLWRYBYettT50AOkLDf6kc3+CydiySlUO0s1xMciMiMs
EZCsrBa7AQNx9BaZLwGw05a6ymjTQdSYO7slcdHZ4dJVsgOgtWbPDRyp8p22sZcT5pK0l/Egbios
18UuCAANbZUaRjKv/+DtFotZYGuGeHH334xzll5PaAL7qNyn0i3mzHAUsrZST9r0ythGEKNWPIaz
Ftx33ACyg5EpBfIrFfsyZJs1sKOkULlR3VTXNbrUQirMwIp1gvr/fmOqWDK5dOFX8geyzawG9wdp
wiq8ANOlpwZ9fV0QYbYbUMa2CBnvP2PJXD22n8mkWHVqr/Q7WgZBk2CFW8ojUD+jFAecFmYW3M60
EhhA9x0VTvR+VragQAQ33AOjF0HMVmrqsJxBTd1+Q0Flqx++PRTDV5t1jfBCMSDqQzlLbPp+JL+7
0rHHgBjYbk/vJIBowhl5p+HnFp9iokCiEeZ0jfKuUy5w1DozDKOOUbZFHFtHePHXTx57whlGbrWw
DnVDdO2DsPn77LwwFitV2ve4WXzKGZzydB0rrVhuxUOhUFFHkFWOts/xlspDkcuL2t2syteiS/tP
PbZAluq4jbmBQ3tzL5LYjpg1QxU4tKd4vRRhThDRk+tfnccHAw5T4iZVGhjRhFNG5Axdz4YEAlpW
EmE1EVP3ELlWtqoNC07qi4TBb+ZxLiH4dALi91mTykagRv7nz0y39howyQOK3jQZKGhNiJ3G1ejM
8NeeJC/BfI3mUtHDfogRTEtxeL0Tko8fRDL+MxcqCGuiI/N3rqiQb+fjKomRdqe5GegEoLWZhO1T
BT4AY0DU5XOOYVOla0+qwj76Gd7qE4pINZVaFThmaacxDJ+8B66ZPIvY2HjJCLc84fEq7YVs7BVT
RjSXgqdXKlGK3lQMljRUjAyjwuHC5FiZxENihZUfCEtvDGgudwMwgoonkk+/SZ+P579F8rF+ncDJ
o5Y6Fs8IqsqL/W7kxTdf231h+Cm1eq9V+nD14661zErPrmtcu1zWJBZ2lym6YCHkPHDZM+B75iWq
XO2LYaO8OJX7HqHd3pujcj1Y90uLBcv5qHXHQwDWn6/gnFLlid/fbkzyjdhYC3oKBWXTDh58GMTj
eCYsT2I69Mp/L7ikNmA8Q5pIYi/lmBJTjAYG4OqSuqNJMKygb3UoU28GrbeLIW5L6806uXfitZ22
zdfr0dk4m6+VoY5HNooxXvOMpYLyvOfSnEKuHfPNBTuWcWoYt1auvs65PzJ6B+aKryQLBeHr0nST
QpnkmKhQucOLaOBkbr/cvGHRRPLL1zhdYmqQYqczF9LGsS4+dQD9KwuGM2GnJFzt0FVn3Xud3c8i
b5Fox7mEdZOGZKf7ViYIUfScNewEX9f0PfrfsDX5ZVrDeOQ2Yjx2y5JuJzpiox0zfd54ZecmmS/v
SNtkKMNmAtUiS2XqgXtuTZTiWPj1wnfNdA0A58F5q6dNtdAEDN7fEOVWUBiAGvKT0HLXLg/sPcpX
ffdqyoy1EI2LfTzitYrvTxcrasCSYYGm9dSAyMA+NCsaaedOnv+jg8S0PIwGsiTSWAHXk7RTcfcs
Y+Ta5wWOC1YahBY0sNmgYINcUhdjh3MNu/ic4ZiDE/B8rA+xwmVeNo2vQZusXBvc8+6v2dKhryCf
1X4vAU00kIXwfyBDPkfw+NHANkWQbEUhmWUizsJsmjYCmkzqB0Iwu1iEGmaLH0yqSpet1Of22ae9
5WG0lA+9z3jCpWKkavJw0eUnsH8oR9dkDeji7u/Kr5gvXTkrjcj2PjNXcZjy2Ya/ls+8Vhcow/PT
hSVf+naLMOryLgjLTROljyi26pV0qNOkZsg6/tVxim2nL9T2rA5dFc+oHz0XG7qs7myDh8qXoE+8
kv6RPjVmf8DQldVted2/zQwcOE2V4sliCuOO+PNLXOkLqfFnlZK5CIOBmUm6wtdn1VFbfFbi+Ja6
aq9VHiRLAU2lptl8WJ+3g5/KSSIe0BhLA0+Ebw56OCKxESBIeDvmiXScDMuuf3c/0dxAi2kU+TyI
eaK2gxLytcJhioralT+KFw+ssNcBF/i9SVoE3Ci9EydrjxH60YejdEcFct957WeK6RlskyaD9JJ0
1VxYBl/wOxtnSsYSsXI9dJ1qGdSFW9+VbDNc3sYyyVEsuaTJC1onJjDqKxH5dWuWgUmEkoyvXKpT
BhkZty9xPWGYSu4cuBxV/rVqAzIxh4m2yWQmme39jmRxrq1lZu21hQMmCi1vDVynNmYIth2AH84B
JdXGv3uKkA5vU86YSZZ5O4M900qsu86MSgCwosoO9SWaT9pYa2A2SXsdpV9x340t/9Lt0IP00V38
Out0V5M3s92caDbIkwg0GgJ52hYiyawFN2EzGWaiqWQFR/2MNKo4667lKcfIpm5HLZYtgzQyvuu9
P9cSAhIEvGDwQrI3UM5vmfTWI3H9SWnwjcTDmjxxsGY1EQp8zWD0bt+bH4Br12gGC9S7uHWOPYIV
5uUahz5f0UDxCb1jZDpzV1XWEYwgwo0nzSR7kcQJgNRUb1TELCMAA8jH7yqmAXHDZJFbj08Y8UAw
GoYiC1Ev/dx6GJ6icLeHOhxgUlMl+wmf03rmtYXjQ0b4T7Lg+OezZBUUKjCXQ3Apq8wAd78vb//+
3yi3pHVP0oY14t1YPh9bp70kRGK3dNv0uGehXIhMSk+qkIQSb7x9EBLsqic+jDF+TZFBFQzpiHm+
KGZ3Us16WGF0P9H1ddiWTtLGVLEez5HAdQ0YMtgLiZYnUKhAl7U3WSLIZo1jAgG9TICOIuGSDbBO
8gYqRW4XP+XFcZ+nbs0fbY2DB3Tvh8BfvAtPtCinpJpOXfuUXDXGocFiUVc5wDkc+RkL1fTsSJhk
KOENR3ORvLihoGk1/U9Ve0iW7/Oaz8a90uUluYXWZvnBmomJC8ytAJ7mOIOyXDjQc7xcdX5d6Blk
G5c+PGFscr8/Nz8Dl8uM7oiKN5N8no5zJ6EMerrHwjG8n08FW7rHpMgCfOSrRBMQJ2oyCiSZT+sj
mJ4Dxtr7quDJ0Jl75G4NGEtWNwKAD19FpBHXKvelcf5ZNAqWhBc71GCZjGGjq73ThXd+yAUqq85V
i72Y5JbjQcv2gtbGIBMRXFzjOXejir5RbFHlLwL/6bl/Jg5B4MJydePKU/0mZ+bY79oKxU1gVsAz
axWOHezsBMBoHmeY8M8ncYI3FC75t2L7qR5aZmpNiQFN4PKx0RI6H71/vixyeCGnRXGSCgLwoBcV
DMDQu1Qkj981CZ+Tgxnlq8piVfiuyf9fTxFNbBhBZJK7zG+xDYWXI2u4nNPrGQknh7YU906lBc71
pSvXjSQb9BxwvkYcBI6xRimPcGGaW4mHcNOIo0Ss3TG2Hu2kL2evqpRuZi8A4jd/4uzeurLEujzb
c0NfNZ80SWELGBEOlixZptJA2gVcNY1BvnifTwtU4O/wGZLnybMw6Uslzzz9zPBY0v6O2RKqLNkd
rNQVTjB8ly01SDxXwpf16At+7kSbee09l36wa1PW9MH545rQnahyJE120SJ0EtMySQr0aA09hkZV
t3U7MXSAoy5Kd55qbQQyRbUD+UXO7LVBqVZ4QX7+I0dYvfRmv2cd28P9xCyc1AddFn/4+E6vusl9
sGsXk2fqqByAv4zqkwk2ToHWT64EhQEw0NPJM1TrCgtxIwV74zPtAs8QA5lyOn8RNN6DgrYaEwwc
wF954NoXl9Ly5K9Kd4dcEsWvskpzWazhbkFn7SniJEOiX4nH53H1KJ5wdGJYEBDBVGylAGtXNq82
ATYkQDe+D7Vyug/60RGysecHTCZe+x7cE+OKxZl/LMesJtuv/l13Yjj2/QUhPSJiLqplFuVjl2nl
uXernNjRdprwbEbNSYCDnL+US+LshJ9a1QGN/qWLcVgWdyuKLp5EjcZteiUH5pFvXBFiPCxT1F2M
38tWVc2iPINPiL7zTZRBocKhuXCbWgo23/fYmCW4wMve2QRZwUQ12U3hT5FzS7aSQQxeZ2J+SPxq
yaaL2hafuqGsbN+/gz/PjUBIKdDzmVSgxPJAYn6Qhj/hZeekRc1Z6X8yZ036QaYz8XE0rw2n4RMX
loZXiwIHIJe6PAvoKPbvDGyZAnaR0gK7nqAvdVe8nVb4L8bzIc9B7UwJRhSpkA9DwHzxpyXmo27Z
W9cGczOpNyXb/coC2/Eq9LPTYmZqOAQq2HxNvVyxohdMAHFFwAGCaqoATNfVY0bP+BSZIFGEkcUT
nEzEMbo2LNtk7YkpFbOhE+UI79ruMY/5UGTE9ruR8bR9TIda7t0WZwpPmzG51orhKZTYBRHuWWQu
McrPNKRW+dbNfqnNzLtqoTMsWphkkUhRUKQbXn/X8UB36YZLj2K0VrwuT1m/o9vtbKLShazziWRs
ogsmwxlM38N+TyOPi8CPvvrn6M2DjPw6hxc4B/08Vqlu3sYXh4ZFzWsaj+X0Yc2mpdHL5XxpNGZA
SmrXYxrVhIW1hT1AEOlM/BzFvpZGYao6ER81fp8IbSuMqCuur35cX1nId8Kx6WSgmRFxdjpUp3HL
JhoeWOUU2J7MAXk7GUzf8r/3V00Lc5KHqKP8r8vuqsG3QoV4dKQs6HVbkVDP6bDMoiaykWaMKzZA
qq3IW6k1yhkngUcbdzdwgrf5w6t4cW0K/Iw/zK5h/U0vDU8y8xTaQszCinHyRjh7n+a/dOoP+qlp
oGIfb/ICldZm+H7WNKL/rn1zXM3HT6SK0Q1zcBwNCw4xidnCKMlrIpSvjtI61b6Z3d0IJLGqBGE7
ALywgCjtQtUKskE3dE4McP2hOd8CCYISYVzsfnQiFqXjSnK+fc6keNERqn8sc/VO/wOYbLQkj8nV
lcKfv/ex4xsxF62KM2olHOcUmlpgeYccOygUbPVa72OBoC4kR7MTIhaGu5jFTMZiF4wx5HAyRFki
shi7sMc7SSkx1CodylDksE5MbeltKDrtXWW0Fft0FLkjLoNLA3YqegTCwB5phyE9HDS9lVOQ+mX2
3NpYU3LhQ//mKIte/O4AJ6BHZorzuRCch7VIKwbQUVyjlQPvlxC5qgMmXpQVqsaZiUr55WA1QoLO
4b+HbAE51DpAbXLdycs1oB3nQPmmiG+oh9xxAxU2MqF+UF6gz7uHvVL96MHZSSRHdiLSBMo/lJo2
+7AQ6XFKCqPE52b3vKcVWVjxlFQb/Sg3VFSrtD/gLGMQLImP2jcXwxIUaJl6AD/QdTl99350BTxi
LXeGaqpkb2RQFM/4VwiouNfjeo7NmcdBL50TQV8Citr3vPXrqKg+/HnLr3hAfYiz2K39nw5HNjFX
AjTXLObLGoxpf6q9fbu5QD0PUglZ5+0dpukKpd3wMaINNpczI0G7CCjSRsPEcSWIPmzUvjFrLKFK
RyxdlNBjkZSyG5NgAT7P6RUdmuzZ/6w5hR9R2l1x5ONLYqxivf+A62lGcj7beJ4UdagasvCE4cRu
+4QX8Duvdfo27Etoa9Ojma0l3lRF+FbGJJe4EzeJmH0AUbCLTCOgEe/1OBBMb8/xW6g8qWu9hit1
yEtsq9Mru6YKOWJAQvQLwJspJANevLO3zqvU7IaFZQV5YHioUYGejSp82+KdZJVJTQvArxhXlf3y
4uzwrXrmG2ZZPa4qY69gE8WiG72t2zPVqdJFMilR1LKAiY4q9OFVVWc0ELv4u8Q0+Sl6y3qRKx1w
L6Vh4vdztA7lGf6DUHx63h7sNwbSWAh5h7dhD4ALWRnMn1QsgswHXP7pbfngC99++nNn4q0Hyngo
q7qmItjG9UFkkNB9wV6rWhZcHpCCSjoCv0C6cZl8XFKW+bbPwyrcROVORxtl1fTG3QboDZwlNR07
tD96hjS4K82IsDemdTnkPHkE9lWAQqSQtqyrYkhS6M9KLXtNzcYg6S7BJcr6QfOdwbOHmfqkmYOP
d4hUjUqZqUi1UQyYm9VZUa9bD+WJaoiZh4oAH13IuYk3FeChGCP3kfMaZJD3Fhlfm8QzzHKM7JAd
uDuy6QNO2WazxXMbXGQnFkHFoVmrtVigC97M5pj5gHMtC4sknIiXM37yx244SaE3cCAeacmUX7VS
HqW7MTZBgwIKoQyd/YWYMZO4lwXhxcqC4+PJeLo/yYFIME7NCw3Uhnyyc9MZdxZpCjAz6ZYTsqfZ
ZhJkrSFV1YaisBYzVkupmQCShiKlipA6TzbwHC8ol7pVnciWOg4MSOkA7IPVi8+PPf1VfTltJ23w
NvcoRuxL8gfnt5fi+dAHkAxwtPZR6I2HN6cH1n/A/uZ/aeGyssvZPG7rfGqkqXyIXj+M9UQLQhHJ
nkEgPC1csrXGUunggKwKncWfzqcMNpds74rhZaZf7ksNf59cOcK9IeM/Xv2CJ0P9HDePEQnuZIok
chP6W5LilJeh2ZPDD7I3zL+y95INavkHozZYMyafKC9seOPi4ORORBmPnSuVLNCte4pBSDTg5dwr
ZqeSZwvkGDo0amFawJlqcL1ck1QXGJhFHcUAuV8iHaxuqIhgzBPxxM2tj3l4ehyVonv7B88Vmp92
uvGS1Rt80xR5GS9PRB4Yz3inSGVHjw2T+bxK9JkLezC87PWmfkn50CJuq0C0y8ksMXbd21l8T9L1
ZyIopwiyTIzCJP9h78OGrAK1BRAWr3vLArS/vHH+ovDa0vRADisRn2F5ftpgpU0Vd6yx7okaAZwd
bX79fld7wxAokNw5TdCdpC7LZMih0M9YzIn/NzNxyWfuLU8WRXfyWYrO5H1bV8yW4LB8UYhgItdB
49lxBPDhhktmpJW3MIMOrPk4cW+e9QjzWX1/d4TnubCvN4ZlSJzXLQlJOhMFcatvERf7ZnjyCmoJ
03QGdQN19Psu74yah5zvkBtchGqKLKZUvKq547ZqbOV6q8UfG+eUfxjyYBjnLvnLaf1mpFPE0LAT
SZq7B1h+12ee79PGVStup767HWnxrVxUEmHJkEOKPq3hIs1TU6wLpKfzY7fFJrdBY2oys8u3h5HH
xqbvUqGWiysmw5jOZvYu1KXQ87oBwwDVD+08C3D1AzkMbQ+Ybmxhga9oo9xcIXDoTZowrF5FFAT6
UrmbPGiaFrJ3yd1uyIqwn5J3wZ22KPu4wBRNOzq78Uvh045fPw+RJhzbxHM5t00MmzTXZ/+R0C3v
L5lgg2mI8YjSGNjujaUm3Vt1LCq5kjSQr1DPHxRSsjPJzRB8ZUY+e/S4oFpY+8Lr9z6ebuxTY3UB
NltSPy+4EgRBvUm3qZs23cQkz/dhOAZ9oYkltdxxb4b7iBGn2OI+NA6JMOy9vq/fD3Q6fQKe+xX7
69M/9DxdyH19FSQI39p43tAOt0DS5ADmA6J+DFG51JQ2goDP+NpY8uy3hatsz/RM8A+TU+HOBOUt
wWR1d3SHJTc06O5acjbqRTOSYEjeeXqx2bmcy8Q5Rwmc6fz3wvTb+w8vlEfMVfK0QEHfHAhvrAvT
SO9/FT5JrGrj5zEOEFsVJ0pVVOjcNWoZkSyWENz/EDU6LKPJoMLL9wLyd0rVuFVMFgnUjMxVDxcn
lwTRu1KIa8XlGdkZNTfIR/AsKB65WwB+43Eu64V6K9HPww5doQqhf7Yso/pv0+AqJpMONTOwu3hv
gFxhpf8ZVaWfOrAiWOz8B/dg6NbZFexozJ0INjHdjIl5T/5O5BvBmBtEOfliwOd6L//BjPT28ubK
/GkqFmWHkx1HWIAjMMdi2zpzAMeGQMLvOXKgd9Y54u9i8slmTNJwtzbd52GX6qxsi+5bgEodAP4V
Ga9366e/uPWu4I2tPET7zrgHhOE3Mkvqt9lUYUe1wmsPktcjAHI1O3Hj14YqJHNMY50RaPBheAGc
fVgKXAy1D46Dr5RI8rJXTJRFPKTMaosdRZ7LXT9YCwhfs9y/x7eig6WrUkA13qz9fxKi/CATJbwJ
drvxg/kfUGI/haWhsoqAKcez5OYDbe0GRdN0IivMPS+ZEfTQfwbcvXnpq6YKHRRZ+td7OtnBLD/c
XgJa30KZpqlwmpLmE33ct9fA75hUHQOMXZEEpI5cPDtf5hS+oOzIYObwWB1SgogUk0jwtlMHbsJ+
09cYdTwk573kefqiK5e8UFhi2mcHjVdJAFNS3KyDbKkuGGnHG5DfbIlgpoFJbuI2P2ce2nEuEpoq
f+DiV9v9T2hdgbMoQtJBOf0tz3wmlOzDsFLo2AL2iitP6JK5z1xK1j4v+2z2OARJ3vOWItAMuiHB
b6dNhn46p/8zXr+ITEXcqAQ35dwc7ns8bMWutqCRy56aUvn5vD7z2P6ZFFxiSTkUgCWlPlMKLeVo
7sKF9gCnHE2qM0NP+6AUWf2SInsO3o1CV5mpi4X9X8DyiU5LqDYsYVRCWREDfArIESxoIZRo47Cj
tqs+qofRVLSI/Qwn7vctORNGw8N5HzM1QWot9PlvNTVSLHHwsAck8uzUgWmjdfGVVsGyikz1bgTV
bwIXS99dI/FlZnpkWFe5YArfA2zly8y1XeOs7mHs95LC8QY3pcS9M/HylhuC7o5bTcSigNdAR7yI
/cuxvW8M4q01DYREgWonDFT/7NKd/Oq/opCRgYYRQymJwXjd0diKgBwEfkHQ5pWC0l0qbC3+b0/u
E+8pz8wTec338tYgi0T5XtbTOMJSiLZTXh04/whK48uXHgBs751W6k4aNQEY3aIiMpaD0V4Ke/qo
AR7yZ9+eN0Ui5aXisF6ysMnXwvtkGb+k2opiRPtKpiUJNJBiu7Q3+kHPnJtPd4UrC8TZDHcvVup0
Nwfubt4qRiZWkVxVxWSNdE2j15iMSu5uYkyjMDnWJnGYTnpVWSlQfBmSK/u81jO74Py7qf4TGiLz
pXXcLxvAPpjqvFyTpFrbPO+Rdt1nKYuKczjr6UA8+7ReXZURMuBWyfTSeqhgCslxjIN7q1nIVkgk
dBup08JbvgWPjll6NmZlJDCl8gAlFOozOsXkrOa4PTXPPskjczzVu/YiM+cwDs+aRNg8aqKr1bPm
UXIMuXngC6oZVvBixBxhFHDvnjFUHJSIMKfAUg7xBBsBtLxwSX+riA8yAT68zKZe8Ffh6cKIu31C
vyKvRvG17kwHyuzjNdhU+X4BLhexGRdx03nuwVdLhgjX951pfvNKIS/cd71UKDsMKbcgGu1DJFwl
tygpxpuxI8YYhssNDq7QrEARA8jVSC4dN2kBb+HBG40ftYv837uob+9x+OfsqkEA+HRB6I0k1UCs
Z54lEp2mevP9Y2asqISBpjfYHcaFSeq6I8JKv8oOffcdJd0v1V3lFpNJes7d48etQqAK1Q47Rq0n
Q9/hJY3hAvJFU/M7ypEvwhnHJ3MIuQ5vSRd05oEudRrqyxSypntX77OGnm3v+i2KwRssfPGKqH/L
TAvH1jb+0Z+HGMrzlpW9ETGdBVqfO5CHeTWuj6A9t2gV/d7SFL2gmzwIbA7d8nCCpiFqPAROZ/fE
eMtoRt1nKNI7Zwf0cbC3KT73wRbJlSDK+a5x52zNIIa16CW2tvdlVuI7+VvBMfWL72Jvp+l9fudj
chBhM8TFaJSl+OhDNWUx/sK0/HLyvWyFs3dYY8KuwFsJ320ooC5+foUAOD8+DFS4HTgAKS4QFImj
5cGmDHADsZ21SJ5cgIa8UvYPC2eHHAi1mky2+6wULNuEblTvIMswkJTzT8Or26Stn6hsxXjVovyX
CRdx0KWEZgJxHOSAOmXbEWhizIAbp+xIGBlFFUkvN8krw3J4F0mYYcNiajqVzs8bwDd+zIOgE8bZ
3vUpVpIMIdUjxiHHvykJhSzam+rXfzLUoqVSEhd/7F08aIclflZdsAx+oJHqxzUhH35n7XXeSJBR
6wOUUQXtEoYOo9W3S1toef0Uos18o2XZlNLrDjubxKKuHtPRInMjNkKkFfHS6ro3OO8dUiNcx1If
yXeuWW/R1Kpvu5SrVpTv51U3FwMlqyKnziHvGosLf3fL9Ba8niQMzEq4yuw9yOCOym9M6nRl4Rpp
DdHxzvlCca+M+JKYnvgGrRywMVTP6ALnB0J2c/Zcy861mmAWromQIkuD1oxdtlbuqmmpQi5MuPl8
c6ojrRrzSgEn9TqErCo40HA4mlVsh1s09is/QybZIKdZvCaURMgP8asOoaJ4I1uwNpe2KBHdLSRR
JiH+2I5OADsD7xQEdc7OGYO6C9YOfa6kN8vXyX4jaIvwNkuYtGk4TzA8D8nzLLwIri1EoUfse4Rv
isibJDfDI49N16Dzdalep3bjGA178RnAfIkSVyUpuP9UtuxrEmimJtnd/UexO/798xF1dDU+HL+H
QQI7bhH5XaPfJ54lM0SSBL9TvpSUAqSPslA9gZTjGfjpXfX0Qf2PBFMI0OxkgIOajdWC++dsVwIr
u6EMNLGK0/YdaZEt38opGXnHM5sxlRLUaRTiWkTUMFplAXoH8025DhextYbS65cQPxq8pB/CxyLv
G2vSLLVFWNmzKxU8dx2CRGM9covexWGVja6jXb+mayCO1B+E5LMCfdLN217jwZhj5VLu5owYgMKZ
nzmDFbcF3VHApAk+xce745Kl4CcOx6baiGNnttdtWs/nP42QV67sEYnYhyQYffuDpKgZCC+I7sbz
Tavh46Q4yO4ihXzWg3lk7Gw5JbAgf+dblZj7XgR48qwgEolB4gPN7fng5wVaFQy+gd952FQJejMB
SLJclEz3PyA/4+M2lggUzUDY1QYLMgvfaxAqim40OqpsEtGGzFGHYimkf7Et4oE3tsT+P3pDarD/
JzWQFlu4sAasglwdKDzlbLSt/OEDYtqzoAtilSO38ji8hNgARZiBNBrGTk26iLhtoDPlGPuFqG9o
n62mfJQzarxMnhmJfN06HZkCg2rX7HTbzrF6SQbhdMaNVt6m2FLWqjEXwsPvTv+WPqsXC5H1wShW
+iwDxnyBYynT5jPVJAozfrsLtdJ3CQlj6TYAnuAhonq8UHqB5OOmkto9fOVWQJdo1JRuSuIB9b/v
fs+zohfH9Z2V7dm9yBQHM3cUVL6WDVyffj7fcffQrqS36VjiAi9nWe8OeREuPpRcyIK/qimyKBUD
lh5T5EBzkrQXblyLZz94FOGKbi6fTlBNkyL1/ddDjZa1F74H/PVFzCgShqOruQuHmpRE90Fc9cKj
Z7XjXpDs4zyoK6/9Y4RgnxSmOSKgrYGGQBFA01L2QEZJgA6YhFsZzI6EjFa3qFnKGEJ5B0VcqqW1
WPTiEA4M32vyTWUbMnZ8iX9YhYYxSJfAAAS0KroksNRGnjD+Jv8rSNOgXRl+kSEwiHcSEhXoHeVR
PK2zJzl1/gHuHWKhSoK8Hz7+J0B3TGtHfyv+/LbhCloXMJJG0Pt0UlN/j/rD+X3eqSv85i62QNpG
Jb1cxQHQE3tUqg8GET1BTjGJemWvh0VYc8txVmu2pfHfcSMyd6y5zVFxus9SV/ddKi3pj1HSeDjF
XRfw/6JzBLfQYHptolIQDv1dlf0rAuUSRx2GCdXRjfE6T+CtrBzAVJKGH1HFgXewgFqkW57YCJl7
K79esiZ8U7QQgxN82kDy10OdhMp8kJIwCssfdFQlacAkusjv1eFeg4+nKIG1zH131EUuKx3F6iCi
w7nyKDanDREeCAlxBB9VstmW7oinBI4gEApJ3ltK5LHwKOnh3uX4Lb/ny3PN9403NzjsMQNGioTk
oXXe9Vlu0qvba8TXWovsxXmNMLSyLp6aFxkYI+CF8UYuzMc+ycRh8Lfxr2GPUUug09G10UwO3IFm
h2QKjpiwyE3xzpnNYCWBBJb+mx2oR3PMAG6ASJwOvqwCOU07/BRTLebDjCqK81omznOFEWYKmctu
0jAPi3SgIlcK6VUPdjAsM4Jh15vDSLUAiNw9Pa3rblFiNNIx5Yhgc0bbOMesUS//2aSDWS8O3m6P
0CY0VCanjE+V+WbzUQAypvK+GAyea/eY3QKH7lfjDqMAcZkEkdmDfLMwDw8phMYs4PjqnY9od0mj
VoY06nPIc1rjWGaFpjxAlEJGoYDWr/ZeX8ejy7z0PxyoMzS6Q/2FTGKooXaUjO31VstT6wCeoJwX
NuglZTuX3xeKtGSEcF2eq5bQWUAK2pcd2XOA/oOcRjPOC0BNQYSMoxrSmXWWowjvPc+4hH+wya59
DUJX2SxRALllDjAr4A9AUxzn0Jw2qn4zwWW/mIZVnNdJMGYtq4DBqBs8hy5kbgyzfWJyX8e3Ojqq
lmOUsUjGxlO9nKX1YH0HTCNZNyk6NMrzfF0dsQi/MNeNTiqosT+LgDuxZ36QmwuPpGn99RbYeDpd
AczawVB8IQsdtM3UQM9NvGutUE+9vhl7CDRnMyNgIIHXfwKmgnIjBe44QsT/NdfXynKtWIKi3NI3
qOWt+NyeuZ1GjxVyQ3+LfDnh0PsfbiGnUTOCAN0VBMLvyX+KhZP2hVuI6PI0bcPck0snG4CX3tdO
jm0BTluw6Q8Alf7GYZ7X0LTcBS4jvH18Ue5+peKbIm5ZXXqEeakEX/0S9I8qRVydmD7ZliA7JEjp
gcd7kM8rPVEEJeKHNkLx6J0TWfe/Vk6p1eDGz/FLCu7tLc4gy4biojOzjoswcfE8MIKlhn00H1b/
cpxrftIB2URkuTq7Z/77OKYHjCiNb1w0FzxlcyfVxYsYKJ2ccxVARZi1KLwfS0jmZCAME8lvgvOi
UTJYyz5000YXZ4b2NxrWGXRXpuYwiC6PEw+9+cW15whkLyGBPf4Ih3/W3xcxQ5jKahAEunmNEdCP
onUxYsI3cDKXsHCzSLdSWthtQxx+dQwsUjWUpKGh4DTpN3LgVIS+0REr5HTsZ3ld4iiPg2ln7o3K
Skz69CF6FH3U2gku6m2tqWOLZ2kaTSZM7rvuPzXmUPHgsICFyIRKmHN0Uy6NqW6a4C7+QGx7gs/i
Oyuo7QW1GFPxdM/V4HGRxV3X/0HGtSow+rchcvavWoleMvCSwIk4v7/Irv05kYwCRwKKBHWRSxLY
CwqnBDOAM/kS/LFMUoJZKaLTS56TExnC/FG9XIeRj6uzirVG8RLkqoI5u6YuXK22FXJ2c9aU5a//
g1LKCCw2M25MHXHhMvAZ4fwa41nHneuEwf1BSCftHLhdYO0aeKPivB8Nbs/0/sFywaQ8cAFA9FUf
GX92cL+2rhAKwkHxVNg4WzL7JfPBwz4agNFyxckeUhXNHQzXQ4jh/46FV3L4D5SST5u5FfoMu6xF
HuuY6duDdCXQ0I82WrjPEVdxl/Eziwwr3CvjQ0dR9RYZWfN1wTsY9q9RSNx8n+qOX1mtDkrnIDKk
buSLjd2TMJtTGdOtfHqnjzK4ClcVyeS83+fF3tmS6z/eLGp60bkrLi9JwU9G0hqnYFsIw5k1CY5U
164vUfWuZr4dGjcYc2aOi+1+7zqJLDdQSHgDuUGpwjfwLbSTHdgwoH7I+DdkxrfXLQizRGGBEiZE
0T/98cGHw0z6HQbtatkhqwGN3RSATAO6J5Tufp1BwagVY9OXiPM2xJ6nIyHyXiO5s7aoHVj8ny6r
eEgHzwqXZAAbeIHI+8fKp6Wsnb/cnS0CnUs2lUn2Jgh8ML1n2WSSh15q5xPuEFWG5jMwxxmG0aGn
EkKCxLfNB8pRHqw4eFySyz1NTmeSjn9weIwc7fNH4CptHwg538hqkrOU79IEH2qCXHNMvI1WJX6j
UzMkm8LKqMctEsm7fX2dq4FbHrOFIbu1m/wrAkb/Tw387VddVwaEBPpdLE2AG/eMZDK7oiAECEhP
c9cHlw/J0x7NjWvYuIIGwqg14epQDG0cm/2O7rsRG/kWjOLdIsJwxg96olImXfLqbkfedrtu+XsS
aHTDwmSebcbjs/0c9P1yuezGXminZZQz+8CiGvRTG5ScDz6F6ZAuaDgYn9EThlsggxleB8Wvu4jB
Ajq+2eQdDR7mUddBEl0f4PxP5JnpP904Wyr90YSRUl85mZl4H7kqUWYietIFxkEd3hRm4SsRbKEr
TTtzvK2GVJA1H+Xi9T1f4MGUMGgg4PrJ57QoCKkGYxKlkpbsedj9DXz1cPrh7CCcVpyiQ4RIZIP+
Zds9ZIwXib5QweWSGKgeumXBYJuA/h0I/UIWz3ZKOsEDxavJ15KG1Unxles/zQwJsoFBoCSdSDp4
vwCRcpA7LZQzzuNNNGyFqPm9GLGCmVmqyDF3GZaod/O74bRPckUM9XGnZ9D135VdAJvAwYp2wP1t
K8oXDWE8/yayUukdCUuvhR3n/eGSq87ru4KY3qC5fC6/6rbDwNh6xtYElkOhH1dgJetmUdAfms17
fwG/2I4RZJttMVixeUOJUD/IRxjqWoIS4DdnyPnfyIi6e9DJ1AEqGExLu9oLfdOtuOuU+OfyMr2m
iPoJU2OXH3nB/oDWGB10DoIfbQjJk/ASrxlOaJSqn0Ia0/svSEtXwNgbZS5qbmKyuckBi3uZDsQR
Fz02wE8l+x2n02zkmW5PKDMoue6VBX6Hv8t3MlrR3ibq2e6p2qaRDuuUIjWuBdzjBu2q+QF9k++L
ElM1pOkQpGN1oUFVIF6rC4Zz4htkv8rHw6XNu4oz8oEne43EYLCnHholQ3Zzy62B4g+kpwFOX9tY
XTS0zL4pXOT/KgT0tquJM14syi8WLyMWSrXmFe9DNCv6nozO96FeL5ZoqjTzJOllOMIiD9hi87Y4
FHYcLQS/VXrr8gS5AbLtYxI5IunMvAaCHr10xJqGztZibxX8PbWjMneQ5+1MeVoNfhB2K6jwRObQ
iJ3V6vwXTPkCF4wwahBINRwh32Sgrn8o5kZt9xpXrLz6zrdoxjE5VspgbZ1L9fOQFTLnFjv98d6c
NH71yz6FNM2c6HIxe2fcofV7P2ThgenVURyH8W5rIbTQqs6T5eL8+3Mjv5bmEJQXpjgvKVgwb1jB
KaQElPB5/drSAxDIgfIr63Ny2SnN8Lp78nwBNTCaYjOIgvjOT+gjFKXbA3dctmNDvkq3tRSx/kG2
9SH4bvcLUThgyvfNt1n4aZoO5TsIvG9DZq+XJgoAss60ohdqz3Yppy0cmJr5wE/rofbvPwUxBklB
U3QEFVc3IvlpK1uUrGMkehkCzW/RwD+d4ynopeOMVI8698a/DUGBv6BGOsXBJhMDJwKZORitBf2v
BASE3vJyMXYbYP9Uw0aVzkHSxSeEgjbK5NlSntgQZIOSwpWd6kfK1F8tJYpWwHYFX0/RYszvdDby
I7BMXpI0peqUk8ZjzuhTcyUmwao/Gv5DqO7+HmVTe8f2o7j14uSl1siOC7wB5olBLba1ZZ20FaL1
sdWEXur+KKESWROxZLL+2KSsEN9OmNlb2TMJfVnJqkSWGzHUIdZaq+mQP4GxJgpJzPXcw01DMqJ6
yQ2E4UZhdLQ8HaPTAGNetuwB8SKyVUvwMHJzVhfrHai+vlrGSN1vJYBxB+RwavEjumSz1HgtUtBX
mKoNyo5mCFoejgrWMTiB3mkEoZXyURIbMnNdtWCaz3vMdRpcYDQwrKWGsK3XwXyuk4YFUDXo09ec
BXggPn5JxdpBq7ZppBudpiCer2cSf0cj43IHquY9Be4/4vzXIIqsAeBFUiiwD/0h6kIKuaJgxHkK
1wMCRLk5kRVraocsYpVfEiggVgK/ZirRJwdZld+UrWYUloEU+JcPsXO2mCcaxMos0IP2c/aTQeCb
IWaePYfew2DLMCngblUhLgJm5VmR+epXERpjgFfLbWzW9HYhBTQ59ObM3vexgP91HosSCZsPHCIw
cXLKnVwZdblhpuTotjI/NNZlYwKDbZ3+bqz94LD+HT+VlSMO9HxbavewFQUMdDxt54/e42CCBJuF
AZVuHqEs+vZnj1ApcqhF52hascNQrgzd9oM3cuHKBhuYWJhh/DmuYewPywr1S2/f394DIvDFVL94
6gm/nrP5cjsumH7NmQcFwjAQjGZcxGSvCAi8wHv4dEJpTz8Uyi0LrDeaOpC96pXxk9IytZ/ASe+X
p3YZVneIufrdWdcFMTO5Iac2xKCFkkcnTs/krgDE665YeBh2xQJw8VToMqXz1nRuLkpcJw+y8DZ3
b84yVpcSgUOAwlbi3mK68HkbxF1YJssX8t7V3ikG5nPO783scFU6i8GoaVm96Ih18BudTObGHCcb
4wAg1p59UJEMG+p80SfcZMd1UmKAVYX6VjR44AUpAjuH8JBSpOrvMeIwInFCwhme8xBEmgvlPcn3
+2EvZUjHwbVC7Em8kEUcx9TuiDo0vJ0OGRC7kG8IlXouD9oYBqXJpGgX3TmWbrohl8nJggzADMho
Y8tMRo6zPeoYWoSs+ItfVI2Mz+E5BWT+JtksX20Cd0+bqPhDsMOLZaxOIvX+ZtsjnA+VnHcevifF
rhcgK9d25KpUAYSwM+X2xgrU+NpdbbbkHnI+sn9Bfy8wSQ/d58wgWm5HmeRMAim3zErwmpWXvXPX
iVFSg63t10XMqD5eBtqe4aH9pamQ9alJWZr8KuGm6S85w1cY74oZnFtdiOIPbSMwaW/DiQjvWAge
86sPPJ9xy+tqvjY3Q8TJJtXZfXUex7VKIp9BTsBc83BTEF/m47f67L/OcHrg87H7HYodcoM5FMSi
mziAoO3ZKzWNIipZgHZeizlCEVXUN3Lz+oDV1zINuvL2icz6/avtHhQnedoXpksG9R0jcKGmQyCp
+K1SDnRZaxhQ3mruKAtRdKTXV4JxwyuXURbTEy0MNEkEI6AJDxbJqE/wFueku/K0r0FHtGP8leBz
mSeeTD8cf7fUaqc5RLEkJoIGqA8PR5JWIaHOZ18YNJIzXIoa2RP9abFbHJ9k8rL6wS1Jp0rJdvif
JpkE97xG2aRHWS74ToMURYVH05Z1brSSDchM6pvyjIuNUB3JrD6Wcp95pYSotAJxCHbOzq8jF4/R
lUJN9O0jZRaOaJ1vzule9dorjLuYvreL4Db7DgPvjKK/jx7iGEwpPX97UBddoomwDcVpLNjh9ugW
A5e/PDVDoWyX6oI49FwBzvUxPg+HmrhM1LkCPaVRs2C6eHApnP6kobKBibx8Bz0J4TFO3k8mDxBr
cCv2Tqq/5GBiDkb3uEw/HZDKqsFyCuWJ4vF9+HyUULRw8aNCh2QrwkF/y0yn+TqYXWm9XV4nWN+v
wPVhmoN+em5qRXktBezpas4GL3Le7eaa0jPzYUQ6mnoBmrUA1NG1bNi5Ix9b9BhE1xiE31L02kpW
xRVR4NlAYdZIsZ6q9L8Xb0dvLqngE3SgnFWPMbZ5b6Y9epV0UOL1nWuTJ49J1TBRWts98m5+0YGt
Vwqnbqb1SfPsrjaUDBkN4h53wXAHN+CXQkXrg7PykCOewSWbL3Qh6NsT6zhpN7rO/lqcvZVdyJir
E7ENemBoxEomJxy+P2QNlvxOfUrfH0jLgeG2SHqLeUs48PfBHNA5qEC8d1mTEt3gZWvdQBWh363B
IAbhmZj8skWxrVvAJ/14Ct4K95X7y0HnE0IzTBRHydGm0WDUy9CLvE6p9PqA+t8Hv0JI96HgdEcA
M1JU6QGTxJCyNx4pfg+Vvlga4q8eTaoMHCtB+J0l+CD9O0ROhfQWrthqsKAlvgj8xN6HkJLgg4gz
T0W919OLykCVhS6MgVw7ZHjCXmR02P7iZ6H0zHZTxzAJIrztidxpd0eObY+aD6c5VPXwtXa4PWi6
yCRC+Rvc4Iw6+ZYNUSeKeP7Wo48VeVV5KXGhC1PrUDSqnXJQqe5/rgSEcH5XcUu8LXU0g+hsEQ7m
XWHS9FvWwPWmR61Jj54qfPPs7DKiTlqJfBf2amDZuVtcSYhFSGxwFLS6QrHumrfELVABdIkc4otw
LeLKhTodciuCWy7fCHYBlOalBfcqMLjZQ+I6Qftbcv2f4JwTLxuio1aF8axCOsn16dnOy8wY6TTw
b5w/EqeSM/8vBBzBJfN4W0Njb9A0DZIRrucLvFJ6/LImTDkWHnfeR4+8GjtyxPz32mBybGNSnYhe
9efvYWe5HSOTdFXaMIWqsg335z13WOgWRuT47sEsFDh7Wpba6FAG2UPCKs7xw2gzzpS/7qAdJhcP
Mx1GhHFtRvU19dQ9Mq4HpeC33hmLfd7ikn9mfSKVPehAR7KTIAivDBGAmxB+GEHMa8MIAUsBFMmD
OP16UpBqV10PbdpGt2quEsiMFzxnGnoMoyjSbo0FdtRgOTCGN3sL7fcEjSb9IqUoyBQ6wM7RlRqE
YObSlQ3uvDfSRajad9BSOhPVwjtzUGmS9kTMTIrYv/Q3dIEitZ+xJNagUxlGRkqRAk8jLhKAHIEd
4fMlRb1ICP+XTUBgXs2OIveSDYwzE7TjcB9hKb03R0cjtrixGfFB7RdgT1gt6FGKBFRqGjhez2MU
Y0KM5kvNjedQHui5TUJ8WhDwdeylsgH7gYnHyLdjA1EBX5uxLfU0OcpV+9hE/VIbPNqrKCj6eRln
5DJW7xiOOXk4XMRP44SV4LeEDm8NDdagCeBtLSamvRjHa3tWPJNlp6qwXqTJfHp2Gu32v7XZu2XW
W+NBWjP8SoH94qDVELLM6AKJEFh4HP3AimzUCYnR28EaYXq4y4OrpxMcpgMzogvChsjtB27pJsI+
C2y524vfNX6D3IfbiXxFgF9xx/u8GTohoeW1J0BR4vjjptm4IeMSX8eVzbESQraEiMqKEnFEUCx3
INOYRG5srpvt69udYetLYvNPaJ1w3e6jjqq3sQB8hRR0ynS1FUr1amuNMDdrskLwGEIIsINFnVHN
vg8sFoF0WHFdKjLCWB3Zp8rQD45sRtsMdYWKyNT26Y85x/o7kGRLKuJyHEuptAklb1bWCKuim+tk
zuOa1NGNp3GNAlHxohAvRF3zb7esvYyKEpMUjhw/q7WMG4Co7Pxra3+DYxImUappHQ9+wzaUdhpn
5Bvc/jUDyAq4q1OHHN2pw3BXloCYJ+LcqRbIiZOiLKEl3phQjg9zvi7hBeWWUHBqsVEfpYBfJnEF
BL7giSpJp9QgsqIIwkRAErKqmBYDZ5ljfbzg5wvp47aGtZMJuPVJSxBrgYhNokagm1c8/nMAA1tv
3+925M13YwPvf57kSFeMM4a3tHMjOu7icvd4dIsopcNQmazRe0ZrrUYKFsEamtqpVKMftCKF+TJu
bHi1Aabw5TYbsFERvVctAMvYTyOpk6+QsqTsueZ+gh4cG5kxtx2cYW6scFml04Yl44dbZPu1Xm7z
tArj7X+QE1q4AhZiN3K1gqUAhchNw+sKax4olBpDkjBT6wa3isSlU/PN453sAh7aoCuMqe6p6Fky
un3zLwEmczcusYD74QmSA4+25oeQ/ZKincD6BNR7ichWwEuxNLiFeskBXwzF9m89OMC6VrpmX4WE
f90jLWIjelq8bAJZh2l9Vpws5ObXbh2PnsEImFAmc/4Ejac+8peiBz858TgMcV+YuG/ypzGZU+b0
g6sC8F+sdY5CPAtjvBIV+N32adMuZIyzMeosVNUrZ2+4LNrTBvfgOWFdXv8OPVpFxEz8FGldubAf
e5nrGT401xZyCx5B75U8FVYBNpyvvhmUufcbP8aBdJNSkHF3/f384ZtNX03tthz+VhLGyIyJ/iA2
BDBbvKcjmSaDzoebTVSU5Nc9kL+N9Mc6EWQI8HGpI9IM6IEUZ5D4euCY0LQhDpUXQ+cB9B1JNVE6
EgLfrJbUBX0o45hCYw3UOLE3VQ1JtXGo1Id+Z8/4r69tdTkDsM1eMjOz41LinpT47ZD9RuTY46BC
tkpBhtBC+py1kt5wJ9Ir0yPGk+tgoqnZtBWuvnKyFezJXimm6wJQB5HX5lC7mqeZlUlGqKEr4p1i
sm4xQSs6cZV/EzpE2o8c+xdnZ8akI1Y58aIlnj5EJY5HlXdG0rtXM4PBZnG9WCLeTloMJzMBvlSZ
xk1ro03C6fdbya82057nYJs3o4xj+GwRZ8lol4q3VoG4nLXyrUlmfTRv6F2b4gmTSoT/PA/Atk/n
8Mlgh8gCEB70l0smWGe8/i6LeLIwXdraurfL/RjQz+SVIGN2Y9fxQXUjumJ8R9CqGZmrx8Mvbttq
LffKrJqahDXP4y0Shd5vy5vxQOK9QkCgHEZ7z53rtkZT9W08H8sG5R6oVmNIJ0vuJ2RntaVFHIei
1cDA8giPT+03LskVrDg8XgZYei0QbT0G65va910xUkAyrwzcnnHZpUn+zXopTG4ym/C70BpGUYgi
GgeGUYNFTgoG8wjn78GtJQ/JtCGrcgkkbGBak/lr2o+76NG/6xX/mvlbfvdoSeS4bGLKyCUwctJW
Qtn7+6QXq1f9Kk7ixr3DEqpaLpIgP3EiC5LT57rHe26LOPhKHJHrQgEVmAKvykO37fWcpmXvI35d
6LKFLSSUo1hd025X9qJhExwtkE27gOE7JA8m5TxmqghQoKQMCZ3jeJg/bJCj9zmaMMk6hFRh9iUJ
vr0HqYjoDQ9Pw9m3iMuVyCDbUSA/rNWp9YtU0l4u//mZnDpq8DS6UVppRFY65HbJveKjlxEWH+ug
ZeHv/75t99SPROU64gv24fbdsTnfLtRSjmlS5jF0B4BrwjLcrloTmsb3F5mDJtobSyzjzhWnhJDh
mtOnRE1zov3YBvV8XXJCcjlEL9a887fm+qcCahKef+FHKAVlLXuV4j1TV0IUSXToM9od6hSUR1Et
9FQgGu9s76ZjtMW0SabIstsO6PzB8n+nfbT7fmm2tAMbQh3VuIB6eYT3/UwKH5A2IN/YpTMZMfnn
ruHJbYzyaE7zEzLMi4+aBlJOSrWWt4G8cjxHYhe1iiXeyIoMvMvD6fEuixeLme/bELGBuAfahrhd
Fzd3nHsfFeXVriVOSkTE7lbPLUGyuZCnZeCdCIR1WMLNr/jMZyjPycQKjwurtiqdy7WSUzFUjPOA
Cxr2/KK9Vef2QAaF0ibWZPwZsd4frljsrY+ndrHg0eqtzOcpcW+eJSccU3ASOFcclyqkxGOI5ylz
XSABecFlPadyyCY8eK1rb7rgxs9cBLj2Fo7pFmOG6/ubzuQB9XFy+tXnflOqQMxQYmoVeXD3WwV0
TIS0Tp8CmMvIcWG6LXesaA/Oyvz31hy1N+wZyKBexKqQiAWO3yt0B0rfE0lK3lodX+553QvQsCsC
5QseknOF7oH7prjUHLqzZwP20Li6norPAr1wMNThyrqxsSTKDXJyCnJEkEb1oQDRHcd+x8DUSv9T
Us20ooL1VOLlm/EIIqwC5VWdCxMAnic4wTmHWOPanBjS27UlIhfJzvBYxLW8a8+2t8rDJsgR7s3A
OdBQc/935YpG/lrAz+hosQ5+ZXfaH5glg+L0a0khxO/aXsTKraDlycm/gIQj+5j81BGVDnzPdbS/
Yh2nX0F/KKRkyaoSf1NfT2PxXR0B1dGuuc1AROXBsxyuR/21q1eQZA1FhkPCp10WNitp1pOoaqOE
jbc8HlFf0xxyLzSeCzukbcdw12VJbTR5KB0nm1sFo6EswdDIVCdQVbetOmlZBfsv6slB/VxjUVhr
uJtfTE2ulcAvKHCrVAuvaZmwX2taJwpj84JsNE2oafgx+Q9h6NLuMbulfK3NFa7q4u/wFCdzi+D6
FSZgBdMMXkfvE+BOVD8bF4CySwslf2/PXitjxWiNoMPFc2o19zv5q97Tbh5s5k35iAwC3E07pzLC
ocgKXVGbMX0Vdjd3yyHdQ/Uaojw1iibo19aK8L3cw+OqKlpcq8TblA0NkEmMpME0ZxQEbEmn47bw
m+OXiPZiZu2fH2ythl+qOsOZ463FhHGDJQi1SyD0KAgTLbfOKW3IlQ6a//VYXdr3kKk4SVz2dg8f
DxFjgiCmgtAgAoWWPP3o7ACbSpJ2q0ZUlIAQlcqCnRwM0cy+3aiLiW1GNTB/Ohpd0dOFa033cUej
QcDt2tGE0u6Yzf9W0e3Bio80vPSmoNZs7CKTYW5pFM6iyaLeOAvh8W4sF4qOMzS6gQ6sWKdu7bB3
aaqTSYlxL+F+qAlZSrUp8jvjfOooqe0JTK1LBLuwhKDNRiQDomyojlOtbbwvCsPvcIpTePIw3P2i
U/GGWytGNRUuSNPF/5lQIpyHi74WC9P3uzQX2lsnQtkXjX6r6OwSbVQelelb+YgleJOMgqeTkWHj
WX27/b/l2qZ0iII9y8XUx3irB8bcFXFttdQnQE6FcJpsfnru7mB8HEiDFjIrnt0cShTWAWDU1coc
0NXPutgLm+4HwOuIvpfaqp+0JP4IappaisQeGBPMpu6PcGfUQQq+JkcRW8qGIaZTk7Up4gcr9Z62
8Yq5FHB/r5XfmFWs+G+P8p7ElQp2+hDwXVJwfjY9q/lt14gSS6Z4sj4omS9vNVsrO77Frx1OHd90
qSlP/F3SCyelJeR8W9fgwELKn4pZ0uuJgRjPm1n7T2LnGjW4vud9BTci8UGYptsb9fUgS/9Yp4bc
nU7VSOVFa0+1WB4OQH9JZZ/Jhpds/l25i7kUpDzFiaYSh3C/VNaO9kppKae0OemW2rf2SA7v32DM
+yBYrvgHx+596bM01ffjDxPulnaoYJ+fwrrb/1EyrHNc4RGccYH0l44vhsqYgrk8F2Gw22ShXUQa
+o7oUZnWPl7eIY+yhaBJq7LFHU27L48ri4YPH6K2Hn0gxREN9Fv/MFv5XkFbwkl7yYPBTAQCb4t/
lQWRt/a25sBqcbosRl9AEqQbUKcuxvWIkL+bTUd2JFwjeuGND+6rOV6cBb2TeT85irf9ylskm4X9
fNs087JOW8ZasMqfEcAoh8u+eJz3TcBwLtUfaus/5OsI0URAZksizU0I1cFaIkvlQ1kbDo/EY/n9
leVNWxX9aNpjeBqN32qYy7FgkX5qLyQr2pAu4ls622n1v7YMvbbpfXoD1VcHzmbr6ipKT3z3f6Q+
eaYxtrARtNpGjfts1nO5zaBFqQSYn/YuZDVszuX5GzP9tPKmYbHIqozAEMuJTi5zoSSsjp2AvD2D
COyTJ2ZIC//kFcgU63HsIFhtP4m2TTs3uBMeQk2Od6/IDx6j69RRg2m2avVxCF2bQB63G0LwFOkx
Tq6JGqZbNG1TClMFdkCR1f1m1rHNh8Egat5E5y21yl3ZcBX1AzckFzPpAGNt+qWeBwvZFC4qY7ro
FbQ3Q0wTwODZMBiZYO9LixJTuPGuYNnuYCrHTuuW8yOqE7RH/jNXrueOrKDv3bRuouwHSlVvWGC1
A/T4fiiVN+1F7gCwYNWzdC5yiUROqKPusXW2DzAQ0pAt/5VuQTKU6TpLzutx5kyHMy2PwvlX/hH2
xR5KDTFJ4C53aeLeqNLJaX1HE7bH/FfiRh7bZc1fvvX1pOw+MQQSmEyhKLbQtHW1TvjbyEA05A3m
JMyuE03W4Vo5f+eAQm7DMjLao0tN2Q3vQkLuWdm2fKbneTHZY1HLp9ff4F2pTpCmoNQIT6uNdONG
q87Xswyi14Llu7H0N2ndL7R+CRkkRz/O/AprOUkofNNdrYcbfHDzT9V8TdtRujYEacJpE57IFxLv
W+k4ZAX0Z7e+FHcUouo/cOw+iuiryix8fCh7sj/UI+Gp3uRFgEUhoGDQVtGZIZgSVRH1xAuFHRAZ
DYphZ7zkLj8IxiXVUJJIdcTXNvgcAOMFITjtQMwFxJThvUtM6YQ4tjuogKa14upzkWbDVqKqnhhp
3JAB1t1NQG/+YgQ85CxE6rqV3Yne4t+LRCXgVUvgI+F846DtUJPAHxkNl9/9QyWON8YaOOjscZ13
DbIH+eh4+9YwuFJiDNLtR6zF3jZ6p+0reAhR6ObL62OoFfj2xTt0z4jKxdYawbBu1HRx6pLLVRGW
bn87rpspAUPQjqGuwxZnP66vrkesSlntdgY2WXWYYmyM+7+ShEUefrGxtubZ2a6pNk+DT7kDvRpv
y0rpVMim4VmIPc8SLQEgIle9uthZynzyJTJ/Ry9XoOrc6YILE1brs8uEYzFVLPl0wCNZ44lwT7/W
3LnZ6rRBbotIwRAwNRqLLpTof3UaUC/NW4C9035tNTcPkTXuOvZCu2U6NYqiMxTlfCPKxiTUPRFj
TOz6og1nvtMP/ogBnKuNvinXxVn4+qOlvtZqfesmIK0Ca8TWiJKaF5bMp2trdFiDLV1+G8z2t0WJ
YP9zV1S/C9unKl2wGC7w7tX0I5EHjtlhvL5YHy1IFC7/CCDEE+ba6/UchM5MTFnOm64elicRZcLc
F8U2F88kVxQMfF0oRPA5TP3HElSNo7iljMQ4BK01o2Y+380ufHP9JIzfKEz/SBlzVCHmdTDlpKMr
TF0qAwY0mpC5Dupgbp4weiyLMN6BktipYv/Fgg16tIW5MbdTdFl1nZl/uwz4aKOIw+RvfllYdtHa
oDyNIO4omLXckYUO86m28tHZPJtwtMY+pjmIBCSq/8RO1uYo5IlWsfVLNhZTBZhnIjJFCgVUWaTb
I9yjDVILVHepSAl1/RX8iU23aNM2SAb5rdqjmmus0rMmRFehO8JSjI+VLUbd44BUNcd9OKpTLi79
oV8HG2P/08JM1yAxVFD0xJvro6DQDbCrlXxETPCpJeznycF4BFShvW9diwD5pRDWQH/wWhB+ku3X
T2Yk0gS74Nukw4FSR3s1/KHTuF3LXAIWIGizR5jh8Mh1LWwuJK6Zm/KEGjDhh9XFKmTUAGFViu+M
urExagICtLw7BN6Urq5eqxNYaC6rMRnglRIHixkZjfsAJz44bThN8gcZ854HYuBcw8wDp31xuePb
+bDefzkx4YSmEt9t2xR6xWjSU+C3cRhtHYlLm/SKDlu7otXXYYfpdomhBq+Oi4hLF8WAqVo5kjhH
gCqUfYP9RREg+Mpj8SPf/RuQo75/yMwmG035fWHMg2zQy33aUjO5TwG06EoM0PU7Ii6IV5WYYVG3
Kpc20aQcijvGF+0f3f6/6rdIUIwSsgADNJU8sSoUd0hdsiyBGf/FognLGrdX6mFfbwiDFBE3dIMP
tVVePXH1t4nkZ/0OtH8u+5I6sDHmVCBohhVSk7eYuRE03NfqyTZKq2IKkcGh/UW6Kj67B8yMbjnc
PMR2vQqPZ+2//HrKYphKgPD3LA6jsAv+uqQm2/WhuEKpd9oDmAgp8YvnMxxhcCQTrjNQYt8Os6nd
x45r9ow1IHDSNzQOwN90tNNKTgWKjevnZ3zbUXvabkPJ+kCMsVDqVIZM+Z+kuCrifTCLT1MptqTS
8mt3SX+6nQMNNhcBIHAWXTlRMOjSAr7rDxiMnbvHoAdPQF3XqPFJLZhRW8sm9BNp/V+81YdLyD9n
W/NFMXHB1JcGAYUn9HEE6BLBtWp38N6vmdJnos8uqDRXDOdki4aWvzR2j9CDVVGfjtIUUm1FObNb
aDdrnM+ZTXqBNRMzTulB8uypvaVdfEwRuJpoEaMu4g2gQSIoEEuAsvhIKp1OxDwwCRbE9V0D4V1d
7ROJqWutTgKHKbHFbEtqJ53I7/c3YulSXJXUHRB58yEn5ECbVxy2KTQRgmcz/LmG5ZQFviTmMdBH
TkNdkaOHy+fRnlXSusNvzeHmOj/3t3kW+d0ata8S46F8OyU6cmzKVZqJgtmuFteqpuyxM2hmClye
om9E++I+EXaSnM6Y5IpBG5rsZpaxS2YakwPAtBT5uC+g5+dVZVyWLp1udXNfb4GcBLbArKQdWA4G
sewvxoFZsgnElARRTFKpDxndw1hC1x4fJHDUQuJsv2zvBZ/3F0oBcIwDOMRiuvNqcjbX2jO3a0/D
D015ro4/kS4jhkMH1OMCxicJIr3ADOQa6DVX5uKz3UgV1CuVFYRo//SejSS4dw6BAxZe6JzztqhJ
RrvSzK0sIfLQ1ZYFNu4ujO7YJZ8hTACzsmeZP5QFB+hs2Zv2uCeVJ60o3grhLUyLz6fYNmXWBtxr
EoCaeHgvDQIKSuJY8vAfSnLULyQE0aOhCif1wFEVegRha+GBBOMKR1h3pRkw4tYLerBSsMwZ9QZ/
G4DHPBQPBjXbrXE/UixyfkjK1tIYT80jv5zlHj9urOjnoH7lk5rbU67HOM6DlQy5rlV+plJeroyc
DkNZW5OFGfNJzhR3ldYWuJCclRKgwpDonncVXw1yVc5b7FNzpY8sPh+g0kkBoQ105+vieZU2mqn5
mFBi9WWgAqn/PPI1vCUMzf0AkdjDDbz03HPgx+MMPYi2ihOD7hdf27jVlws5EfoH1Hy8hZ0hu2bj
GcIv5HNq3t6D4CpvDZBUQSwxKRLuha313vFZmKrYbKwRbJhkBJiFtlTmoC0D4fmikwpcJ9ZOeAj3
Edk7EPZywmeOda/lzr5lRUK6zYcHoZ4yS4rKPmSmXHxXJ+1ynKVAUzWEu69LeZ3zUbZgk7in8KIH
HZlmpaULZToLxZhrUqQrmw8o5ckwBXJYocyd1zd31FJ56M9fn9JDORgGeLBwMn4MWSHx0eq6xRRj
MRY9sVfhk6Wsc44/QyHs0OATnPKkoZmu3YzkekMoQWhMN/cKVKm2C2nbA+UZPSZGxscNR8UbqCUC
iJiOyzczcxBXeRWtjzt9Vr9qcw7hKER8GE+Tc4kYltjYDMLpn14aeimKLyeojLZNnkfDUj8wj/nO
bIPp8zgv/RnjvkFRVFYKN5Cb7QRpwbstX4Wq8QkidfEfyA7/2ys795q8p5kVt+PdEyqbklgnxMah
sEfS5DyUcwFBW+L0tIiSWPBSG3/6Z4mKKboiVXM9Lv1OcJBH3ZHUvz9of2zOCb1jISPuSQudXRyB
n7ioXKihilJzYe4SLubvy/XY6nkRNXSe1XSbc4+283EjzYVNeTZelEU1EWBn2Gg0iUOpYlzW9nGh
TxHWMNUrWbOpFdM8dHSGS2u7OV89+WrQjFzcPN/Zi8Cj/anrFZWxNg4EqZvr1AUDwyNyOF5gHikV
V+JgZ4PQb8fJgOPY8pxpLwFZ14zWqFWOGXFA8g6a215So7P4hRSibZMoVltHFdk4kuA4NVlDhkq3
BePxKcJohxMOungvXYM4rQ3yIrJYaQvVPsEquxEJc4twpJ5kpdxVy7xPegPfP4aYYU+ewHorj23A
S0woutLtUgp7yeZZwQNXSzwUcp8eQKAPD8sPAZLI2tv8o6yXz31dfsh1IeYQFnMfofqLqnWojKiA
Znz9cVEkNLl3StGr4gxoCrdh69Z+lFX2ziCCQjecKL5Ib4rd0JZ/m9BiTnJFEksa5a5ZYe19LXET
jxvHMHLR7CX6IqtfuqO99m8z/yGhgVn8gdSWxOmAuPCKRjfX21T7t6P0z0/4X56/JWk1pqdNbZci
avknWPZInS2rRIvmKtE5gpTjiLZsPY3heNn3YfAjdr/rHNEoK44uUP88rJv420YG5SLZq17NZsTl
kSfKuCGDINk9oMmEhlVRndfPhlhn1RLrqgP2oAqXTH1ZaqU1lSVtdmycyzSTeWFTM7R7039UJrcV
MEaf9LIoQO+mck2EeMTUuFhUeLlB0PPN41w8IGJi5qy1HWdu+vw0+/wtbeq/sSrPuLd5gqrPnGJe
lDU0AcSgzJC1SmyYJeEZ+w6zxQ4X1D+Ka+XIqyPvCoC1Ffw65HWYTiVhHXqK3Zcv1SaoHyjGTYC8
8geLtuoiSNiGHLUpUfsALfvhguxDrAo/WmQLRinNlKfKBjQsxcTSNx4Tge+oy7ATQpdkI+nWpjTO
FEFda+4Pu+sNfRCzDAR3V/9a9Usj8+LMKioaDLteaSbsFbf9yQM7EbTyZXqHh6OiB2U3Jx5DI38R
9vzk47ZAV14oVi/bLx1jkeGydRqk8vqZM0/TUh01MhzfjFw7w2XTMhOTnSxffrRxZWqmudKoYncM
sQCWg70enOzd3ZOW60EPhB5KNGOmHBv/YqDcN+kalywCAa9PI2XoBuGbTcXp2VvpoHE6/ZRhOrlC
V5tEuIcHtiAa2VLOdzT2eZezOZEBy8OjutKb96+SRedao3Tq4e/71JkpVJAQonYiXsnQUCsyZg2o
OFiE7O3tW2erzDitMiE0KDzqOKY3mwwuYw95DBntxL//WwxTeCJi+cgxNnDOrduZT8qwfJZ9xBxq
W63+yRXyvH+PtsSSgUtX1gQkydaYbKB6H/sT2LMVViN2lwC6H0RL0rYi7A78Xtlbk09OJBJZE/mr
9RaS67WfDMqWeCxIf1/iGSgo0t+Ai3bXkud9dy4up2kfpjEB+i1oWLCOqd0k1kk5ZwUn8/FNM7uc
/jcDTQ/Wq91qVV5b67IzIX44ishQhmbPOwF3EZuMgK/Rcwsnc4qJNI22iLdBDS/e1MqLFAm0pyUa
KzFtLIvC9kgrTNkdIPvhU0ecPLHyrpZuGXEhKgidQn8j0wKjo0+lPRfHkG3M8PVX333XAXTFYxC6
JQdBTqMxQM/qZVO3qMVA3+g+kOL4iIb0Dy5+DmESjVVs7jQjBnVCWFzBCuxU2+RmWBDP3AOiHM6f
QL9YudrUGEIUcViqSd8R1jCcJ/EaRgmzUcvJRS3IxgQUmtAxC0owwGml+plXQfVqkQIjH27y550x
EG3SjW4wR+jPJ6bY3anj36sZ/4v/K9QCEhsuK3BHzD2jGctvzPT6P0ZMO+50Sk8v54riGcqdpDgV
Z/4pauCGNoDOQnTrE46pj0Rm5E3LvKe1+zrolNibtLI7SUW8W1w8uwu2QCaawCgtr6V4tFWih6HN
Ssm1a2RT5T9pn3klJcDcqq2bMic6HcvSGzTCPsW6N2E9WP9oMC+cPBiraXcWF/EiVNHjG4HvlSCU
eeKQVp04OaoS03eSrBKvggbQcMR4zXqBOzWWAk1VB6vcUgsPFVgfkq2VczCP7jdSs3gamV3bsT8/
h8s00L2+7R8v
`protect end_protected

