

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iisr0ydwFOm3eepmhOYSaxO3flYpViRsLN97vKyw+ai+x1TubmaH8qRRwK/QFeVsjlGTFdxookcr
olQwv0bmdw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dJvTzz+PoD3n2Ot9SgKfpEhIshJxklhDhS1tYcrcmprfs5wN+lN+5Y+o9jEEql61IqDkJEIGu0xp
zaDWEeMqwkFuovmZnp/AnbrHb7R/19zPRtwSyZ8+VQRLsRMgscwutXu29fTUST6Ribitutae85tQ
1okc5mYK0mcSMIggcMg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZijKIWnBSOuwn6R4ZrzJp1qaSPGZMrP8GTp+SV+Sn9xEivGxLJtGM40xMLXxiYuxIopDD/A1usG6
HkSoNT6OzxHJWKkUEyyVzrZuJdNHJ5q3s3y5LSNY7eMxN9lY4/gygh7aVIBAO9YWzsWu3HLtrHA5
2vsUFQxQdkG5OTLVP1rH68P4j/dhqr/LVHw+9H76c/knGyalpHLRC7tnHQcfuezFJWlkzaNGHfUo
b5cE1YTvtdlZVmw2sVG/GbXIRi5fq3+Okdy+JgckZ4dVWbI20rfa9LkI09/kwD3anyrnovVQVx9h
F0AxolVKVVyWNAaSu1fvXllqzrdJiRLbdnsq0Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LUajPw/jRTLlmEKb+9YylQ2jxw4jlSx/1GGaY1wFfWFdMwK2p0xvQMjui8K3EqJF0fnb3QNWuQDl
1vTtf04vcOAHkfRCeW7Mbp8qeUTtAsflGIPJDxHfVU8ZKprwANsENc8LVrpJ0WnjDFQIzJw7LDqc
Jj2TofWjKprdxXsMnu4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KG6kiSPrd66zvVpG96eKD+783ebVLVFNF7pXgq+rCyBBRoa0N9Hp3DIWK5125mkICodI82zuSq6k
C8aCiPbDiv4tiuIn19WDNNPL4ncknL0KLZTLAkq0BIQIsnFNRaZegM9aXOdMYGKYLpnjSD9KRWRt
WPXPZfwprSu2D7PeDZMiij3MY+cixttgVmNfcx9Kkmvg+1B5sTSDTVs3fqpJBBO1YslTmxyJAIC6
uDuGqvQ1138z6f4f+f8vMXratK1Ypo3jPPb4FTNLYJio5Vd1Nbpl9kRRtj801Ie0GGhbggK6IXJx
785o6wX6g3tRyoHXGJ4DGUmWlIHATg0KIAflYw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13424)
`protect data_block
Pt36rSfu7xOJeQqpJCiuGjlOR4l3jw2H38hGYRduqV8CZAaofHispGav9tjKUHNuFuuasAyS7xHb
Aa6OlozNhunUS5ST6sT0RR+CGhqZkLZymltE3Tl/1RWhk44WrgiMEXx1Z0dBxmWyYCoIHmUlUeaZ
+w/OagclM7EmHO8IzG8S85UQSu5YU0k+t8Qkihx2Zp+y/veoXTiYOuPjAY9wwGpjfOZKnLex7g/b
a0DcSJNcMj+sr9Xud5C2cZeLLV98Ahc+XsnGQ/CeWQWW3pR5XqYJzf2N9nj9W+KJQTeWx9OCOUZ4
VUTgEjDjdo4XepTJ7hWWynlQbslYW/PSNCMVVj2xAkWhfKjLxdHOa2xbkfyjV4iGyDqCdXxNoIyF
IT7dJ40lTygGDH6JWJEax32itPY+R0sxiEpAunLk4UmzkpUXlFa1zM+SB/GgnAlvM3WStbZCUBU4
hbIQFL9l1s/DfPUxxJ13fA6JDpOh73LLAv26MNIhFgPxq3Ku1MsZYkVNGRQwjFM417HZfMVg1JM3
ES7YLZ1blTenaLs5cbO4EPqQg+loBYTKiPoy+qjKWMdCuONrs2wdhWu/aSP4Tx27WiP5U5YGpkny
5cxde3I0Bw0+OwBIYXMtFO8lrxSIz9KR7KJI947CInGBoNT3KslXf+o1wpVF8w5QhlBzA/UKXYUS
wJUjwEOAc/eS6vzaqbTbRBx6BPsjXndJkNk9Uhg3DZQxfvkPaEPATHpIXbcnOe3qiFv/BI1MjEWp
ZdHoOcS9vsFW92rl7BSw+qIaHELiwepvRpBf/fqfFAN1+JybznBQ26ZkrfhvtDMI+pVwq/o5XJ0N
owQRWF7VM3YZPGF6FyYeYNUgEnkEnscHEziLSjenmaPrj1AckWyzLd1q+0HKPrcxHW6PCUdY+nlz
G5XyQqPCG6ZgrGKB/QDrnzmvJUFQhxoLIp2wvwMKcTa/rBpV9Jg7+DcF4RmxvPaRGBlHgwzL4yg0
BDkKAm4czkfIuIQk+MtkGactQfUAPJDt31grMSnGCYRM/c66M4g9CaSu1NvOVqnIJx5oOiH4o/Ae
e75K9kHsS5lNTY3tcYt4Jw37CxsTSfsavPcs4G7UncQJCpokcJb1uLpbH+KCHBdeMWblM2KK6qPy
LJADciqMp7PfwbUs4dxnhPgxWf/9tRqmY3hJn3gbSXDNst/xmsDkpmfvIJ4jbHW1Js8m1gPiShDL
XbJlz1mBfs+PDB8IC9pl6lZtfqUlbZh1i+CuLp+DtxtcRit05qWn6ihMC7QWxsNyGH/gMocsay04
tmJ9IWU2PP++nE/cKjvFt+UTEubqStnBUkNlgWZiqxC5URi7UQ6BjTaBlBeFAxKfzDfYJMuc96T3
zzMdd92WFzyX16o2+1x9aGWXw2o4TkFeMwLWggDwQH3qtw3WyfepIOHrp5HbCUSOLsTswh7Ry9c5
m5CY9Q3gijEI/zRT5WuDsr90B+8eFXGgatfDn0zkp4Znjk2j6MPYyIUC6DGz9IurGy1TWlb1ORrj
HbRaLbaAE5dl4EwJKZD9lVFZqjYKGkqmYm8d88WronzE3SltzbEOsdueFfzlNM7kmmPAKb/gmZOL
116GBKyOinqckHFoVGIzn1MEFeZWWtNMiZVX/bNuDqCWnRWRrnlyZJnv0Afn1khx3oGImQT4RR+R
kqjlKzo4VU6PPHsc5UYr0tyhG0CQp0HG9vQl3doPVm8qNgjlTiV9JvjNqWSkoz/WIf/PtSa+qqKk
dJ5nlqoUJQRRgv2chYZKPKOWlKRVkhinZMhSu4t/qXRkAuG7/uY24KqBoSDg4znmVTQLOqqraIMf
bGrHwNuyTC6TA2gm6aY1meDTFBaeHIaTtVtlNEZWX1k6ZiwXMrNG85YrLx2FHKAYIL2OCxUZFTrd
jcCMPzHl+KODEGj2KBc6258oe5D/I2vs3FWce/CK+CaRuTt74k5FvX47JEazdeYv+Qn/NxIloFEK
3RzSaD5tkc016N6+eKrFy5m5ZneDvv6LZ9EN0oRttUac17ytTbMXbLW0CLmkigalyTLpUdfywsX+
23plvA0W1pba5gxI7zoaabL+twDr70IomsfpJffzJxsHztFy2ZT6RaJ0tdPvhYejyKbyWLQ9jrR9
sMpE8LQ+6kHP5LSl99iZisUH8/eMvkWrewBWOgJezMjCx3h4MX0uSGu6d8sr/MFfj2SJWO9NWeuk
qxZ6IA60s9grqtWovliog7v/JKnFJlkzB88Hgf7JY7WJnQge3p2qWeeWOgGKFbgO66oocLmc2XEI
JoX+M14HHVQroxa+iDN8HuZi0nhfsQeK5HCc7d7XJSeGEJrmsde38NkCdYAYce0I4d7GuSoBikp8
yjMsmDVu1P57br7lrWPNrnYOd5y3Z02TO+/+NhgzTzojCAzEh0sqqljYuQUc2sNVxUWelfTDDDvn
Lr9V1iP6+RdkJDlS/Ff3joj0HxJ2fK+QreVK8nigdE4vf85weot1vI2lM+P5YPRu6cJO3oqRw5cG
zP3IcAeKrVSai3sFDkqmK+cBBbL3qbobf1hm2EapE+IhcYFpee/yfDNnJsP6Bv7Suxd1/5EqimQk
3tSUKvjudAeU9m5qT4igP23tIU+U/hIRCpKopobBtfZw3+6+UYd9NXReioP/CDfk7179JmUcIljt
IRyV/m+dw4TFA4769uw4hJjCwzkFa0lgnZIzkAczpbyyo2M1Vn813eLjNcCFbhgjcaVWxpWTNEpA
YSAcky4KkCJuiPFZ4fggsqv7joGrzVHMSFbzZKom/kMKPdJE3jeHhl2DLnRgPyCjUYIIyvqeN6JY
v7BHMH7+Sy0W6ZP0/5elQvKs+bG4JILQAkkdJYlEByJZWF2r+K0H9bbhAjbgUuFI5tfUy5zdC5My
kl3KK/5iMDNTqZPm0N+L6LnlNNdN81Z4V29UziDfQomXoyIFa+CuhEfIjj6sjrSaquWV5raIQM8p
FuBvOzaXZE4fNSqpT7oWMQymSWVbHNYxQmnPwvcJoRpFrTKvh1coIFwpVkRYivjj4tkVlF624dgg
3vQ/qIqP/qCu7JpaOBS355xftO8s//WMQhl6Ykdq4q4fR7vMnlW6Dphhbs9HhOlOv5oF8vsqMI53
fDsBUwp2AI/RjPonjD9j0LEIL3uvHoTFvAcX3QyurtTxqOdJdvkFCOXoFFpqgij8Csdf+H8TAT7t
zy7hka7rrftU4A+hWiXsJFPTF34r0u2W4aPzqYVdCTuM7V99dDGt9dXo+JaU/wOALLqUjjQr32LO
v/Fp7UqXzF06D5knMKHbfKBdrNlw8kMQOlzw3+8hTbiRaW4LGooa5vQkDB2NWntobI/eZ9KuBTqI
t4sZs7u/J5HkMlOCQxkF4UCGL7xpOTWTFKiCu67I1+4uDFI4zPY35XYYX8sDZG7McV5sJOH4CnC6
9VjGWG0ORxtXVDRFohRaUtgVMT/y/thBXktzwfka7WOdvkpRgddA/bi8Qd0DVI8lISjLslSCn0v8
Ne9ZS7AgmjFQIQdBnP5Zg5XIVjGZodLHYwvmQP/9GVanwbzijn6ALS6loayVX7o2jXgH77+BtqBJ
AZam9osSCI1Es/qQSLHXmPIEErjvaqpPAEYSXqq0CIGjabOf71ZN9VQ48K+QqOcBi+eHHL54Ym3I
9kPt/W72HWCyhzhFy79jJu6NYc10yc4j8AeJST//kprMOaf8BpEh84bAZ4bKEkHkSvy9Ra9/Kczp
janttveiWezROeD0CsWBdhWIwuF0hvOivhUrKEpISSPcQqZ18+GDLA9vSJrhcdktq11SyfmSIR69
i6fpbKYVb7OI1ol7L6t+sl0YCg1TNarOeoGh8fhDezd2xrCmjGzbN+lAfJioY6/yVzPP8mbIMOw3
yFwp8+rkPo5tdwjZP+fUKS1J2zhGaofz0GbudGfSUpgxs6J1y5anwQQlWDzNVhJNAYUmlsLNy8VK
wf1qQhpgfXWyRfGPdmBM4YFx6TTEnAgq3Q4OJ4ZgTkSi5Cno5s0shXmbRHY2SogVfqfl/h429Zn/
M8UPLFDItp+3bgdcU0MBbUx/nY6AmQRZ57CkNV9fXMCji+54gQr0AzZm/86bJiJ2TTCmQ/RYSDKp
/voqtYuNv1bObhuqlX69lqS+r726FLpl4sF1Ou3qQNfCMfFZOSNFoIWNw3j9peTVAG7ZH6Uc2JPU
QxilnxkvMZiCMm8PWuoZi7nm65A4RE6QJkzcJ1MYY6RUZttey+ZxyvGFQEWVDCxKsMiBey97qP/9
lhDp3cD7n6dPPEIA+SBwjWhEINl0c+urg33uJ8ll1eBp/K+5OsfzhS1215XwOAWiCjnXz32lcj/d
JkyMpcLhHOG6/VsLrK4TqIHQFXWkQaaPJPjccxePDd/BqHtDADtdDaOcxF78qBPC2NPBaKHI5p4f
CmWT/U9KAZ//dGTEMkp/0d9TnZG0qYkuhGuZO2R09mVNwibvNlp8S47P6xanp/dBZlpVCqQq8tuO
oSbmzCCqMgOj46FQBWTtvycwXGwAQ/Z1inYK4rB6KsMF1rCwZ0VGJ69TWJHmj1AW1k6ePPqjiu/v
6ut/Nk6ImBTMp/Wkcz9UmZLLCxDxmXSepGw8iFDdVs74c4wCMGECK/ekmj7ZcI06aDTeHQV3xJDj
Bnr2CJeuL4Bb2nB9RvzsOscRzTP5JeTbf612jigayfF4agRXLS4WlqD0O2URTQuJDj/mUqCIwO0I
8kHIpFwEXTiMDRVavqXoIHz4NYSjEOY+JIXRwKY37bfT6j07GfggxgNAC6mUG8WzYAaeX+crp10G
Yzhqx1wRZxcfaUhVaI6whbYNRqSrGW8dLO+KBoiJGNpte9ro22E1lhsiOdY0ixjFvWKia7HgxMtX
SbqmS8hXcqnd5DsvY21zP6fZJ1tSP8yyHRKYNEAXh9FbsZaOllTlPvQQKAm0Vd0O+8xs2EmkZpoR
jCzWIzGLdDV89Q8g93dz7xkUdOjEE2XN1zS7FZa438mCCUvAjrYD5vVa7RQRl2ItX2aPKyHpyKJc
QQuxdf9VtckZK+0x080XSPJWTeKTgq0ypWS4JaZcCjalgBWX4YKYFIF5Gj3sXZkPUwMDCq2AegOa
7MWqETxWPJAgLHXNITlRzAf986EvstYeFZmLN6mWnRyYkXc3VfPzytDS6AYj2/vqo9FJ22pfGpzK
hFKgU//0K3SRMXKMUa4Gm/Cc1Wqb2x3P2Q+h7pVxeYOs8r0nxiucOr71VA8c8CVGOzoN2Wwg2z1D
cNTdL/QeYOF9ILClCR8KXQjGvqsX9H/scmthjtgLqQSmbUVY5VzrybdgM9bv3VDwxtYXOrUdOOJF
rLxZN+rzKcxFFfenA2R3SuYbjFpJYykoaYX37OVVpH2UkEkWaw15Y5rsZHkRJHz2JhNNQzT0wf0l
kg5pGauACeCA/b6vY5oT0pMYB9Yts7M8IOiLPFbdha2XiQSp1ohNf6m1jcnUtF327xwvFcgzDgsQ
0Rv28DyhB/6Qwi8h5oHIv/eslVnGnBHYlqhsiY46vVImk1FitqYRgqIn6v2nut+JlYPSU+ND3zgW
eG/O8Jknjp1vOGmSkTfoacb7ljTwP0U/WRZ6ljinfItNPW4agVAccpFxzOYCFBdUiP4+K6Tf856q
PuH5QMQ7igL8B7eeywC4gJXH1/pnG9vEjxKjQul9IcYdq4HVCuKCISUCL4niNB0noDCehe7fbi4I
sO2/ScGYP4q2p+6dqudkhseCgGHh5S2Nle6ArDZhp3GZ1jHqZHef9geWlcLKU5kdCTb4Pe5gh0Ww
gtEHpq47Fw7uzHDUJ3OksadWLIgWBjlf+X5Z3KZq6owvyPN4DiEl1MpirHYweYYHXkng4VV4Rd2i
ebV0Onou9hBkIXIrXkaFlqzqQLxwLFU8S/r4ADA9YSmy7WWFZoGNcoJBfL2wK8PawfwQE2sJSokQ
GYLPGtGbGOl8PmRtR0O6G53BTSBRcFX/B3oFvlIuXXXivq+YuiPgrCSucJiWzXWLm7aw+UoUgY1R
zpovsv5es8j6ddjNw0GWrA1Msp+GxxYnFsSl+vVAVEe4cMjBwsMutotiBsloeXMM9unxshiAdPHB
5kH/B26Q0i9P0FTGJV2+smWh2IehEsfjhnzqMXh+GUWgTOn2eSawnO/lxtubISM0MgM31FBQoKMN
tHmaQ3VTGaA6BWB0lKEiPNfVA6akXP83WyPTYzyw+1/u/KTWYCxRJ0yZJTXev0lUck/8t5NybCO4
URNvrVXHBc3f6eCB78rCjmYc96Sw8Tw2DDFHg5naZwDKY/MkMbB5tGdkhfe/6pjUIpLK9MTZcZQ6
SaiW04avRVRt5nIZkZ6SwldR3Gt6KhCzPhgpz6SPtym3jYs3Je1gTj+D+Ok7FCxsWwInHvsjnyz9
hBOyBIQZ7OcZDTtQ5a/qSsIeBHRRb74iXZ7phe7o14Y5S8HDOeoyrsOBxa/eyCCvjsjgYryfe9jX
sHOsYjv61a6vp/u7YtINeUdXyRieDtMZ2QJi5AiUKOAcERUrj4X5jIIeSA2sugtDAaYeR5LA1OdD
GXXPPl1Un5iY+CK0pyj/mr/rIrbp8XsjreaGKw6PVD+NeXSYInWsAdnhbMfS3Vnd/5B2HKIWuKaw
/smLLBOe/irivCvBF0VimsXhbvQuGTsB/9hDvSUUGxsLdyBQi18yZ37OFHHJiWz285XZUuO43pUy
pyN7RPvCtoHsyWkslVUcGV/rCRjVDTN1SNMaYePias103C3zbDJ/bGXE1CDSBHh8am9ij+WB6zlW
1Nr3nlpNqkGFzWM7+Km/KCnq3Q15D0iPJSG8Gs7y+h8fPHPKpFVwPkxzwrHkMeLDcYDNs0fgXUuQ
juR76JA+KNj+ZXrrAfr5CCYu4esyy0LHXAKz3kNoaeUFB4Vz4R1a2Ub7dAXHI+yaxZ1oMxm2/fh7
l3kLCwLMLdY2iEkuKTM5kCzWXJ6uUOa9N//MOjGqMtL9PIz82htAvLe6fR20AVL/L3+XzJc/Yscj
MmPtDZf85DWApArUo+LF5hEnmebN8jrxc7MR1d6qtplxdvkp/C9ioi7JUeDameob6W3d/mOAEp5J
mLNh6Spyr4dxKIqW4QP7y1iGB+sFyOPkIx3JkhXCSwKwPidJls8PP4zI6sWtljgftkmaew2viaHY
KsSquSdAbB8a/5pwbDK5QTVUXlUcmx1NR+8cGtC3P1mTnSInyzmt4GttKT2SiziBrDYCZ/7LW/Fu
HhJAuSMlICSz19eZHGMKGL0x97FsybEpAjqqQXOV62U+TMAuLrlrabR6EwI4WwBgUwgvE7Poak9+
Mpk9TnAA3GEccSvavrrzhPGzpEXcz0l3rL3YjOc9poDj1TjgOMBx52J+UobJEEwcjtWoUDQedXJ9
Ohq8a/EsXaO73cKzie3W2+Dx7N4eWP7iPxyzcoQr3ywlshgaRADi4Iw645KPMy9I7wk9Dm7TF+ng
79QtEsWQIMQDwPsXlP6yXdYIz2ZnVW8jd7ws/Vocz0kJRoy9yU20STA0Gojb9MP5YeqUPQ5qgv6E
NU+1CI30VCJPMWwtrihnopvJ5+YDdWdg/SQgsKK3gg50geZwXNHFdmtS18jwLxSL6oMdmnjE+gPj
f/fvN0HmYOjwIZLYeb3CaH/7bGFbjpBygO+iR8sTq2fyVDUMYL3XxEu1c83yT/TPAf2CvDtQ6TmZ
e0Bkpjij22kE0Y6CaJhd8pFeW2yZliNiYNXDmSAQSuK2+uBzrjD7wz6wNOZgqhZfg7gK1mpOYtNf
7s7oweJfqK/d1NA/cozltwXQCVwMCRHBU0iN3RC+kN+fX09IuJoH5lXlw8cwKF5LJaWsm0Y7xpi/
nmIIBCkP0FSLw4woRSv/e1E04G6BI0rUitk+Ub8/sY+yjrntQO6bpVJelzabgEd3IrNkstVQjBcj
JR6cSqRrA+Yusq+NmX+JDM3uhYZsbui2kGaDhMgZVNvuodsS6UhHpKWu9rqTbhm9a8yw5/QIRiPt
B5wh0CpmiAmCCkR8BSoHmaHT9rSxNGgH7jbVYQ5SU6xG5fiCjLhJnCp+CXceury+pvX0DcKzhFJp
JXrux4dglI7na32xWYCEDokWTSC8Mj7miMPlNtm30ybHn4e/glGz+j9ZvX9aShJ2EK9bfZkLI5Vq
Ltf8oXOWmDdLkvBgm9lSNxRWvgXbgVEORSfNr5ULTuhPiHzJSfqEPi2qXOPz7AnV12RafFo/0JTK
pwpZLtxHC/fTt2bvD54tN4smhb6ZBQwmYTYP0rBNuFdj43Koqy4Ne0NfXq+tAnrv3wFbc2+eZ+wL
ng36niVCQLil9dbTDncfBAA0Y8oy2rl/6MmuJkr1Os83SzmenIaza/kTBa/sljrc6JfuDn0cAvGV
5U0iJTMWLRGdydfNWg0lhPYxUKEmIdHpvA85uWp6I/iet7l5AllhvSoyeJzQKZevDgSXP2mH8ZT8
pyx5YOoKhsLbnPdEqZjqWLkJBSOLaVV8ajPqzzqf73KFCQxi8tEcw5szRYcCCfDBm5qXsDWSqvfz
8t4ws8q+Q9SLnpqOZk74PCGHW4T/GTBCkQe+GtvEj9F0gH3fo10DfpCwqAJ/qsdhVngcFDJ08Des
uCVxKHVpQ4QCoLi1Ko7GoC2Pk0+mhhL2LH3/AQIrpgrsJUs6IrACOW/is5WS2WNUsXWlrHvDyTlN
zkphb5+5dt8AZsGssJStiq3w7ZfknASmQPYM6CAGH8kSImbKYcEUN101+B83+6n25BSTVULHEKxC
ffRSzOdRKeFxwCPDLKXvLuivIEr6PfSdr69sKJhk/ItZQHtEyCUymQcQovfmVSY1TwJ+/SSEKW2U
eg83v8Q9FySffoxOG1anYDmQ0vuxqvJq36kTfnWEAUg4/dTwqWv4ytD1hr5pLEKqYhIq7bq2F8xd
FcNNUc6G+PnnZ4JjmXVtxqpNNLMxyxfEsOsU/XqbSPhgIOtM4FBoTo7zmUN945/mQupNw66SIoWi
/dht2fPjuKjhgp07pc3oLuoPc0hahKZwD4tGgn257/d+mrvlWBpAvHVx28ziIoALVj+CqDKmgKnN
vfHy+R26qxH5Wp9LGjuZUdL1pFMGLuI6nh79Ggdk5pVe/mg5wqQZ1u81+u9DZzxJdEkN2z+9HXMc
hiOnTliynQii6pl6n0lrvH671R2/VN3yRBTHMyHmG/Lc6cFWBPaJqhJr6jYRcM4Bt4B2DngoBO4v
KgwoAupw+vo6HqFlGWqz5rekGBXTnS4ZmFFhjfijGsNUNHfEWuwpJ2JXT+5dcij9WI7KA0Gp8e8m
RL+BsR2dmcFglpRbY5Kpia5iuP9W7mlCA4Cbp5W5IOPSTJ5UHk2WVGrBuFBpXWQMPG1wkraE6Tm8
sa7uJcYPdwWPC9W3cnCxnlcf8BZ7ewwsLqFQnSRH0ahs5j7jgu56Eyd5qFMFGp4LlfmMyevuCOko
pgtBKBwb4NOpg//o1WwOKB3IExclMdPDJ5XlCauZzxgdGPhNUED6iMIfJfv3FKF/ID66n5/3aKhR
ffROTQBHUS0Tl9Yqj6A33j7Zp1OZzOqE4rHEs3c/K6caqQWMfarDcTKRGdp0lXEP11aNYzg0dvmo
CfPtPqdxNahGkehDSUR3O9Tr/K2sUp/o5xQvY/HvRZ/oRz7qNAXLeaMfPM2ewYbL0LM29aAYml3W
uRGCkIvDFB7HL1oScoNVLvAuvI3teU/DMx8tXar/kz+3LG2KL8OdPseG61HpJLsohrPJ50dB8sme
jafXyq6WDqASA1HXQmiG6rP9svrgNXarlBFs7i38301EL/3pCXB5PitWuoGBgZ/n9eiDD74PUbaY
pzOtJmMrve+MHW2FGlPEarwOr5Kd01v8wga2xIMm0HgP5XjdLF2IE0t79TfYGMlrlDAZga7KbvZP
Fcb2TO6rMR5v38nCcLEVwf/vR0kUWPZWQIKtGd3H8vClGIdS1txq/3IJJI03l3Hll77h1cUQuxrL
VjCFCX34kx7NL8h2iQWuAyzUIzu3kzLPb/q3qYQPdi1VDzkCsqJgDp4Af6qmxf1K0zdnJbh3t6Dx
OHHdQgSzC+x786uep7xmpLTf81J1tKUMAUdedwdaXZjbS4Yqx1uaSpVUGO6kueRpAv4TZLuF0dud
QjAA3h3apNmfVdALlT7z/xn7mBjvjzBYU7NWQmPDUwIDhZaa6YvsAOVQ4dO/6hb19sw6l2tcwm7V
lLY0bJ7kW2XrYS7sSodx5EjrdQ5Bw6jFF8kthOg7Qlz+XmV48QmIXJoQk5KpeMDkeN0OH4APux0R
mh2dtksvDrJUOGRcBIQ5aegC7h70tzGfjs0IcmTXL4dnoPxod7Haomd89qE/csra+W02LLE3BqwM
9ntpz5+vnPVx3ck4JfHbDoEtHGLBDMiw7orNamugaC+qd+smlEowSSEP7iFhLz5ewS5EmNml29jv
R5sYWC6v3S7OfQE1gOgadNQEsdIDWQ0h8fFAyIS6+nRKLlxnlXx47KZLbeaRv5XpbkkmDasxkpEQ
ZPej70lPNGXiDfhekbznzz/iukcUOoqPS5VNCZBYKcWn3Nei/8WmU8Lb9Cdl/5LlhcRXghqBpX36
Cd0Uh0OfuGfcZM6CscaUeWBMPJa/sdYV+x7yYl+jfWI6jcLSmZidA8dUBDojqXJUgzKmZCooPnC2
jB2S4dBa+NNgYpeO9j2TJfRR5yf/U2nP+p1PobF0fc5sx94tS+vyA15cQJgML8RznAJlNTxuMGLv
rMwTO6rU5wCCNYi4ABRpX19siIS7nYjk66aEzck66B2RnHwKmLBa80gKax1oE0UuxYgJOr+tweed
GVzdIO0t5oK8st3a+Dl1K73u/6A587T0bWgUiw7KoQRd/acMMnwYw526UH3TB34XAXh0DXUWatQm
As5yrMMqhFCKPEqfmHjgTJ2npI4aNj8KtTMIRB9Us53vAxYcHhykESh1IwickeVIDdLF1nddZRsx
EFGrF+stW22ZNXA5gUWBD3zj0lw70LaNk+rHTukx/0rOxUn10ZRzk8k3q+sTm8wa0Ty9NGKJJOZC
ZoUtXm1Mj+Zu3beCDIw182Q8LF1MmfAiAr8Fx/IO6uMA4DAStLVmWvkfjIBi13vQGrv5iBcRnZ92
tmRusdqpOCXqZDziXxuSPJOEg6tIl8+G2YR4kf9/wJtCatRR4LYKf8I9SamlkWpwMq8W5feq7WNq
XLJBeumnDQrRFcD8ilWEGn+cuNJEobnEkTwsidEephZODs3qgpzNeDWqfxNWWA1UKL0LDNUg4P4J
ZAQCL1yIVoGHjmjOT2+Ib9V8fl4VSFCN/xNYQ5HWPDzHkDrTcL6h8kRu9qfvEsF204+XH9lSnypn
vyMe8fTNcaQ+7E/urJ99BPORIiyePJ0tLErvw+fDXxUpQSUZ8CHle+gePSTeHCQSIUrpYdTOikB/
/jgoVMnSoi+mBmbVj8NR1b1GwVPzaX2z6TDqREU5ZMw4mbFo2jmdRWGNPuJXUjQM3ngDjEN+1krq
xcs2qAKGRpYF673Axkfl96kCMF1Q7JxeSRXKff0EcBRzX5HnRvsSB++KIlaMLRRDb7qHMN+J9IRv
5tA20lIou/z3dZDuuUC/LQlxQqXPNL7l8NH965hIJ80xkmFIN1SSSambUUjXJWxWhH56oWuYH/7G
zs7h5YFRKzZHOiGdjuJvWVnEoboo/Y56URFf5secQroziD6iGQ3otKbgUyGXQBFVUPW2T/K0x8/X
FhnZOnHb0VBScTEbb19gYJawZpB48bRXHhh2UKFNa6EO2t0ctT8MS3NYgfNZYgSo3yv/EvEW0Yr4
4+s5gNo8yurQNCc7wCyUQduoGueMRw8oxed64jMmKrfQHefKvxR3Ffso5dg8rCs78O0PNBVA9vDa
10spkMwjhd1Jskl+2/VGNZKq5COTgfeM4r0WPxc4oMQIiSLQr0xLMg+q3K3jUtO9+2XixwrjUbR+
FgR5pmMsj5QjFDNPyLGa/ipXdv+3+VFZC2T/hSyo6MjP59pQqUOSVY4h8ko7dXMRF8KOhJluom+t
PZDMRzSarlcZl6PheR4YuIQH4gCs0OVsSwpSZku5VAmBa48/DI3K5xO9bCScX2us3+nRN3qsYA79
/taOvHI52a+tEwkpc6bWqehKrRPvogAAsZ6YE6e8OqkpUaFdBgn19F9QboqjOStN+HbFqWZ1T9sj
LA0+ikwweaZa6CIVjC2SmewrhOgsDCGleVp6T8AgEh6RUuk5+wcii8i7wVf16OsyBXZoTOReMSSv
4sywNPaBOlA54OCH7nXppTpGqFcwcN0P/b2ZqUVKfI6XniR1e4ht3rixdel6HUY1AVeThGbHCuu/
9cOuVAYwkiSOn2e1vlXpYLlklOSJoAkKlTR5Ysag0IDG+4dN2WKtpvVj2yA6DrCCJAj5uOKZIBLM
KDs2wlEIue006Ppt1gWAvsz5ANnivIDUUh5m7HzppFPZzxfTHpU2LlgGjTige5j3WmdhgAxFltRY
pRV6ok3nNzxQeM4R6801PMtssLq8YwDwYXT25zLAz7l96zI2PDEVw5DwrWHHWTWRkz7ckWgwVwkC
zJ+3MgF/Gdz15wckLDPICbw3vH+I6lXBoP8tUYUQsFnrxnLxcf4S5PXX8cgfXICRS3VBmcP+b5gX
qjX8oj3dWesbWxuaQGcJbgvnsdND+mk2HL6G2qYGSn4PFc7VhKBR/Id6yFT5+okHvw+CrEu73dSs
623TuO7a3zPgOsfCyXtwmsov4iwv+Hz+UfA6WVDS4UcWTqb5B4Daf6e3tsQmQ4FoGZLU59T9YLM2
/IyQGqz664KEw7FsTyVYC00rsO9zOwEy04m+dpoDCBmYHHtGT38zlVxVChVpBaT32dZ9XBWckWVY
nQsgYQKXYaQ1hts2LwaS/oYV0/pp/bEu1wJf/pbqbA0HniQQONEPNxaW8QLurVStsvAAioODfVoL
Mf0FKfxJTybjL8kDiozOe9IRJyzBq8XSEsMu308FT0IVC44PfQRm+gWqhLhJCDQdiI2FizYZPjzu
Z576pP80TMIkNMgw/DK/B2RFBdQqt6OMFrWIvNUV+fGzPJpGuxBT6UQ6JunNA5Skr2W2hSQIndXq
bOhhrpQD0Ua9n0FjbzuPN5L8JeodPbatxfJoHLcGQUNcvywywgi7ZC7TqfHd0149Nul2aI9+cayl
65P8GHQD3v8uDgt46PVCcOhmXFXipK4XKRLUljvpBFlhHoBOlJzWNpPyj3uASEWi1tNcQVF+o31S
qpmTE1XaTIBQXLpiCKHvSjr1JlIH6L/SOI+lHE57N3KXmglx+ZPzQPkA8GJmpuaEI9doDnouAlff
YjbJmbtIYVmgVqsIib4d6Ee97HX4RTrhcsjF3Qz7uEQ5coU73/vbo5iPR24pyC1XUEKRIyH1k55l
dy8ezXq7B/BPuu+ESDXqdv3xU+SmNdEK12tplOO6yXIGecvc0xF8t/XoWp6oYkHcW79gnswFX/jo
vxbpKVj7KU5qrV2uz3mUtbvzQaS+MjXqwNs7OchWC0kob/Iq02VXsYRpbY4DWeRLJ717B4JlEu9G
WCj5gjEiqnOIEf6LGWtxpmhJx6rses2bXvaPXsaYf/P76JU2L2UPTD6qoLlmOk/OzzV266qdMzgZ
+jF08IUPQcm0dhdVSIXTkEaXrqDOa4cqCvCfiTfbWdw8zne0k4v8r+M6zXu6cr4vreN/bAaDa+nQ
O/RDZ85TRVZ8QtboPx2Rpft4Smtn6gB5/EHn6yc9Z1FyFBJFYhX+daXTMg+FzU7U78oKzD+UGGj9
bnHza4g4qguINyB63euGSeBDHJ0a8LlT1JWG7bRZr7tG1QfaRoBMGkpER2sCi7GBcZ9H0r9K5Uin
gL9wJGlQD2PEQyx+4R1rQriWxEAxc7GasNNlC/Ex6GLmbySbOXlx+8UBA5JAYXZwWQQFh9J5zG3z
MB2nMM3DHcnGzCCiHQk9AnBILI64TbM7yw8nn91/1wt9zPsNw3aINeeiB/lC5970zsppE6MGB5s8
3/7rSpXsMHThAI4lDOYLe+ao5mitCxJ1tzvgTeVcFiBl3XIfhLVY6Jj/sylTVw7XwtJu0kHjSNH8
czGFBvNEjquvtvFV/oNxXFTDI82TDUyVeYuh3WijJMwTxnG4BD0IOZnXd/1aQ7dXDDoQ0k858wYS
9yvzFk/St1GoCX0OMWHGsncAZI2NZRzkpaeNUlpjz5OGv9fGBJSvS97W+0gXTT1Ttos5NTCY8f+R
xtnXq3ywa1deI2h6QCr1Pm9aMO63SIgsEWtw0L3YyLbY0qjGLvbF/uwSHTIEeTVAj7KEO4bHYUs9
n0vmnCOZPwZjNcjHFSD0lOb/MMRdNOuLM9dIExyqwKe0wt+iVaWxyGOivkeL+2F+78V9Cpgzp0kI
ujVyGyBJTFzX2RrzqpWi5Dg5ePKbqN719wksmGwvTF6170iACUHkD/Ofeq/VP59e5mzDfDvaVXdz
DdFxBowBwIZZWAYkYwRAv0eRMKwBEXKqDiIt9nozWG1TRe1dy+EWrg4jSKMTqDjDbfvRuscaJCKN
pDtHyp8IxkKD1Y3qnxK7zFK19SP9G+UQu+yvu0LNTrOHoAlWT+VgXYFh5kpFsKwQ6G94yc7d9TGS
u8stUNdOonLhFDobkUNLwEELLMhtd/ViFiB+TAZ6T+kjtoyMtikyLELMIKyL6R0PBIKJXMF06h1X
t+XigCoqhb3pd46GyAMnScIR2cdDhaj5DVJaqrBHbo56lVRzMlMsA20P+/9c6V1CIiTqZsEfclC7
/ehk8qmiDFxlUYJeKJSRVB697KRIC19eLAlBRqKpfCkJ6kLWL7E9s+E6Df27kR01F70djfP8sEQ2
sKBBN033hKSyTmk7n2cFvKzxP/8I4hqWfGfJeUbdqT1bc25eqpb+eAGTnqkBeMX28Uqh7axT5sYM
8rfHBSwfn1982oAHJe1vKfvnWePYEIWvs+8SwkX9cOshFg98mONL4/fwYvDxgxKeKIeNbIHQe0PW
N9ytX/szbYzY6U6z6FedVBjv8yPMCdgm47PGav8S3+v0zokdHVaoV+Ij7SyR6tSAJlNoT+wuEtck
raFcTE0qx8so/xMarsfviONx8x20K0yy76ZyMsi4R4P7Q24CiJTMt+muNEuVjsOVGHbNXn8CsLdm
URVGrYSCrxhXuqb2U+wVIPuc1R0pKdqv5XYbU8w2Z9I0Zo/3yBdRj7YT6iUbmH0qdrN1z1utJbld
2EUGfxYkJSpi09iRCMHd+pPA6IUMAnB0+9cnKEoOrbbU4XlbYvQAu5BP2ROGbtVsgM3IZg/1E/Af
KNb8oNN9mUROMe5IWW0DMOJ5JWA6PUwnG+lr72RxrE4aM4mGXHswTJHqeBqyu+J5ifiIXLaJWDFh
I0903b2IovBfthQFW91fDn0b9pAtdfOqpDZzlgU1QREMEWPyLKIKLWJO/wZWGuVDM6mHdbHfrRbO
CBLsm3ZfnaBkqNe1W3gbXlmtYhk3ndiBTxn9k+0jp4JnfgzU8kqy+ykVa5j9vNxHRfE6OB5Cx22o
C8EGX2xR1FfnNQqe0up9bXSZCOZBWdqPQBfK/UN4mu2UcdcW5E9poajGqwK5DdNkL/Yj0oDH6Rpj
wNoM1/Epvrnf4qzpPSMfc+E5CizcpukDI+1ER82NuJhwZnez62f7MuIX3/eQtrQm9x+nrSBVSHaQ
UYxrtC/gsJEI0EvNDcoujZejdp3ZmONmR1iGncb11NcDj0hjSueA5XHFWfJPgFfkrXttOq6gVeEc
vovaMxVC7p3CUlnOzwrjLY5ftR6mZbmXbBiGXSKQT2YBrEyI6rp+hxmVAXeMnmrg0E9wqKd43KQA
c8Rikl5DmeRn5whX0p/nWcDxdx6EFgMt3yS9Y/5h4eUj6rGDrAHO/DrvT/SgDMxUXC83w8Doscbh
DRhNBTooC7iQOCXtrrbczimGuCVPIbEg+oaPxyEZCeCNUlKniJLYan4PP2c/ZjZO/q76/tpBU87E
ANDCBlVhOTG6eNSDiX1CddVFijbsGudswXNgFRBD0wf2sTVkLEHa+ED3gjMTCs0r/XcPgYI5x3dV
LRcnkbZ6QXHu1XvZ/Fl8tcrrY5bFVKTtkGJzIt1IvJusi39WNJmafVcSFH8RxbHBbzD8u1KVrevh
X/8HqmFFJi2oEUwQH5AAoX85f7ZhseNzW+8nuFNv9wEfZlPDW7EMfh9eYsRiCvogg4dqtECJzZ71
Slq7379Oeif9c7G04p4C7iJ9V2dU89e5poIjf4Cn59d53LXLiDXDfGjeX1bHSiKXSjDawZidBoW1
bCFJebEG8vBRaDzL8X0h+JFVrgCS6At8oz9OWYdAW38e5E9Y+rckpbv7r3//YxSaW96W/VGWpRAg
f2tYlJSP629e7Or75FlbuIhn28EHmLnPdgZ9xDgcjqmtj4i5VvyhDonsRTkqW6Qq3jCV+CtCxpWu
7WNxl3EAoQljCWWS/BFJTyrVQUKI02oQZl2s595MrQ9V+amx13KMy/DNzyFfow1hmFDc735aapXN
VXwsDZdge70LvR9g7l6aaMw1Rr1WiJ1kaCXDLA4aQ4w2oj7Ykjp7klwH7OhBH7fpctw7gfVyj1u8
G2OywA2HsLQl+rgZhNQtJzXSZixxU2bZdRmXRtcfROQJlvlAWuviHjAnsM5iLPGIboIRgK0gVuYC
YQQAL2r+lsvrnw4ol4xq6ByQm0RcYD241dIsmnqNm/CSlh87VJwm5dBJvuZeAwSIM2pSnUM4G/jI
0PCMLxJ4na+Chf6Ytd4IB4IqoI1G+eyx/jif9FU1mn5oojsky8STBZJIfn22l2v85jEygA7zP38R
ArmG9mIsFh8Iy+AQgNTJKU4eix8StnFimJzmvf4UoZDbLqs195t2CPs4F9uHWGPrOa7bvZySsljl
5bBv5ea4ClLjXnIJnrvjji9UK53eHMqpDCekwPx4MmxPlj2jVbdrU4A7FWoYSn7xmL3sLB31Ja0r
1hdRIwW4ZFyhVruv5CiGb8wWAUdt9hWI/L2KC8YhxR5pL5AdfapPgq7uvwz5YHYjydQsbx4UGtYm
dk3GNljUsauOikc9OgUZhylbyx91+x3niNN1Nvu33IUge4EqnoISyuK9XNQW0lNKnQrwJhzbm/PZ
7yc6uVvODlsZomv5e7BU+sGvgdkm1JXcLQEEjclql2RjmYvb0OHdR9MNzENX9lKYSBvDtjIn70DV
K/WNjgb44tNjCm//xX04pBRYYs+zKiRbaOUGRqWJpwV8Bz2P8ZglMcA4hgUUJy2YCozL/BmfrsE8
XKeeGmUqGn2CdZPItCR3pf322DhTTSfi2fJPv3jaK07bfBsM5X5ZSUIeUQcW1H0yvDhXh9bmf1ye
DPWDrtGAaPE96kcgL7eiqsqCk75E2F6BkJIkd7ALNoDTiD3669iKBpafrsveDzpEfuSXZFkZR9E6
XI/ScsK1c1DoqKJL7R9y2KRqRc74LxVK+QoeFnBU9U061p5lGPRYNlNGYDe21ePCn7B9VuJC0Wko
4wBKXgTe6YiGmL6bSCEq/nkrTaP21PBolHpGsfWOh2y/oVwpjXktmCvtiQNepjcn76D8XBNceBOw
Ep+VMY9aqyPbq6oXP7PYwe3ALMgjdrIpYaw2Lf2AHdeZSXUC5aICg+QX7Di333l8kjPViBih2Gkq
FYsw066I/it8biB65VuQv8XPR4cuZYBS6rK1haB7CfZcjLoIvyLA1W4uM52O6x1KSkQCW0U4BYgn
rieW9eU7OuNplJ27X4w57nEsATHOzjDg8I7BUD/5D9MyytRgJGBFQqU3KN//PSXDpul9tA+d0B9V
uAF3mdYox8hg2iBLHyn3g0QB04+hw1GbzgIlnYtH8dLV2tGjUukHg2cRGw6YvK+fa8E2efm4LYIr
4eVg4Xi9SqNc7/KiyDd07eBgVQRqfHIeiPIvqkA=
`protect end_protected

