

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rLWvNa4xmaUmUmTsHaZZpmf+vdo1ZTZAwtQ7nnw7ufjv5GWZXhLdNQy5Q06lrQkoXFZkjYTdRiP3
F6m6R2KGJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hpohmRSyxraB2TfGOSuLyUSGGabJEMublC4fhU+HZ7LC068YGUgk2aE7EHkl1WtDE9Bb6v5v3Qg9
2I0FD8nMKFfSIsem6wrqx6FPpal5aJB28sq90dkao5/Iru4xYelKhv5oyEvq5w9fsErMuciA6N4Y
mVn0CtqFHil9PLQizOk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e2qQeTSxab1fevbjz90nhYXx0vSvMvWBAXsx6NPtcQGmGbeJ/S+FZG17TXPSmNs8pJl+7MKHcPRl
s4fPkRF2q+UUqzkqGrUfIOlc9iDcSV3G1jvuqC/KwL75+As0dV2zHDw3g6spyRgrF/QyMSev2EDX
wNjTOD0D7tDHqk1b7PsRTM/m5LabqbFbAoaZk3OIm0Vx4hjx1H+Kj+5LKlzym1OWRKYofd9Pxrcb
EMUCk84oHB+E99UNC1xkjUMB3ggxmGGz+tj2pQbz0ixGcWE5awa9i3czC6zJ21Sph72Xl+p+aRC5
JcGtcY8i/+JbJchaWispPX8x4NW4FjK9r8JxKw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vltTKSM8a/zRJ1QJ/9B9ijVL2/YbgBrtsRTG74WarkSfaW1TYFA90LAMjfijw4Dh6V3t9bzMVLiX
18WW94nb3vnRj+WAyEjiDaLRKxJmoyxgwsVe3baoS8c9YLsCvI4C+2FRQmKh6kD8j1o6xfJUhYAE
QHwYAw6Gh1Fc1rWYuMM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jeozeC2hZr+0l/LK5n/W7u82KI9P5tCxn4L5QInLhVBS1ZXkJv19EUcHMrHeYhgivoQ0MQ86TEXP
Iah9T/vQMV+h0mk/ZiG6XOYby7qUUR5Ipu6A3NdkCDCZw1M+w2At4X13RPUlLeERzh2uCLeznee9
UbtfGUHB0e0CGrBNEj1LzA1bbcGeOcLXMz/DrWLUmi+Iv7nTaL15UXhNNoh+XY7m46jwFf+dQiLA
SkppMG/4vt/EhyL+TyDlc4FcuyPEIIJCq1gQ6KO1U+4QL61Qp9FOEA7sAw8XZEnuD8uyPmi6wlXt
gqJWUq4qR9zExL8yZmy88nYYAn2YB3+3OVd4ug==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 123472)
`protect data_block
iDdFRnNFrBGaUZ5YNW6BvHInjsZ31I3GqmQx3i1l7JtwLILh0Bwj/rTRH+sx9hhIlLvjlKeXOG7c
NhaiscwUCSzN1wwEBsRhrifWFOdNp0WNngSr1Sf83OX3OeT/k1G4ovzzrqQn1HvXlhPLJHYUCqLc
gmjikR2XJkW7i5teb3zcHN2PYDkOCNqKUWet/Zd5JL7txnw80QYvCtUIZUwXZST9Dk6B2C1M9u8b
zWdQbDqsDdrZ8el9Vw8C/wM9yG8W0h85qfhKHQ4FhFQ3AhKwNRvm7M7stdmM/36tVhQmji1a5Trs
IKyBEer4I2fwDF9FIDLDFA+npL1Q/ZKW0RiNY4XFlZU9adUueAelQOS4oqwtxW6vmSeYDV+OhuVU
39ybPxYQ7KC25exUV2HrFTLkvY+DdvJVnMzp7xCfQcKVakngre5e6CTURxcp3eYbTguIF4wh4hef
AdiAreJzTgct/Vuz/QyIFvc19sg1mPv8xLiwM0Cv4i3pSOvw+OmRYPVX4tjIjNDuos+5c6ybAS+6
Lr9b2zMpTMNGOv/f0TZxtBy39VbcN5OLtfnmW8WujboeH0kJT0cMgHFgsvFeJbJ8nlDMUCzICZkd
9lB68G87vq+8Bfc+HqeEHfjwMG0xx4oYNcqUWUO2WWbBiyRW59Yc471vkvfohsKz6UEUHeYoaALg
97LuWK6fceDb/9DU709bp683dh6nDt/d38sEM5c/waiyyZ/CamxiANvBNI0zXIt0HJgFQ09ktr0R
+QvxhvfkFIHq0EwAdWC4lM0L8JGzSVIAdyernjYaM91oc7cwxODGBzdNikVuQIsnldKwGStIZtiT
BQ9KUbrr6Hrs6snQUC7Qbt35aWuPZ6CxwbgneXNax4NrJqeltx+jLkZn/U0p1JDpWpsSlFtKYQ36
7c7ova04fTPPR+xByiuxT6uPru5fNBGb+lrQGMcSaniF/KYx7Er1bhVkNMOQ/wEAiJoVO9tVcqYW
Jjn7p2q1Oyj2rIz9O+RvT27jTa3CJcY6Ozfx4Op/6qv+DlHfjoMakKOsn5dH21cNG/9bFNWzsdce
HNfnpK69zDjuSfOlT0UejJSF50U5sj8x49IiSs4cAbksIuf0Ya3fK/G0xfJeGr60uVRPsnNoEk3V
ip7wfV8RUPpaT8koBecMlzN6U/4zPwgWZxdSKxo5sJ8yGBqChVrBaR3c38xDxx1om8zHr37NKhku
orE2StngtJb0riLdZ5NrYYrYcVGZRaC+KC2rLJvXOVuHjnbgan4MdI80lh4FBvRYRVvvuRHX6biI
Cw1sVh6cBpl4t7xdgmLy54sPv3yb0SLWwowwhVs7ZgP89V62i0RJeeM/V11jxWFUsWjPB0DFwM5w
hxGnYK4v4YJrbgD3I9t8zW4+fWGjszE1djdWUw2o8GdPqjZ6Z5Re/bj+DDB2C5Us4JWAqiCmD6GE
jEwm3mqL7VmsA0ywEvOjVZJbwD8Kol/5yC0Mn60RKMfJOM4cGsLyHBTlwGCRK5XILNrg2Ov6CS9H
b7JtRgwOChnlN7BGIrBY2cXORwPI7eNNWLQj/2kEVrNVRBTcynkNTkk0idg6oByL2rrLTZxf3JVM
bPMHOy3w8E/qwsXm3NLx1GPaBCoKP1KWoJRwhaDm/KCNnJStG7ZA5rIUqjGKJ3faKgdpsQb/RXVT
opjCor/XT5ms7b9IDY4JXon9m2kfcLzuZzKHmSfyhPj2fpTjPUVDs/PGi9QEGQALN4NceBqjvo7a
cz6b1ucSYKX+8aWigtl2/oia2o/vKN0T0MzZqLA99rLG46yqiayXiMXtHOLIejqLD9OhJnCIhrE8
X/i/W8Fhfg+I4BtHg3+Pw5wjJ+Aa8SYUyencavyIksI78lXqSIODAwrCLTG7WRiMkqXTmmJu2OMx
Zc2erH8RdApkO6m2DXuoEww2zQZVdNbES27ShR9nC8RX3o9arWKKuUwH+XcULCi4YSKgEZC25hpe
7ndwHdIT/RmCd39H++DeNxbtKrOZ8sR22ErSZZCwts0J+aj+UibDCva4lqwgSe+NLa6qApjYUw+z
7jqIDbCvBQGWj9lJIuT+ERG66uoIoL/HeOfV6Nyunm9AykUzVLZP9Pitg+Ob+r/qhdTYk8GVFhnZ
9QeWlDBd9VeycvR4wyRNsDmCusBnCs4BFRVS//8+Gm3Qb13nmU5ykpjXkc0iK/5Jgd+jSAZgOvVB
K4YglC067ZDT/nI9GcTKl3amsivl719AW1eL8Lt9J03J10kj1izwosQFR5fT1AhBTHfL0aVqYnra
mnZJPvEauiB933Xh9wsb2v5CdQtnYgo5ZeMsPTOJuukkAtLThpPbNSNV1N/KS8AU84wsWJfzh0Wd
d8+yhTdW5Jz0FUYGo6qv+lSKEFtpqmYv4FXIU7402i12ilTUR77rIQvtjUUYRoNSJO3KhvejdE8d
pJJh9H0cxXrjUXHX73ch9NiiT8cBbg1yxcrprAvmMlput+ijaeoPZ90yfhVKb8frqqjkz3eUPTBJ
tw2pAnYAUVxS/zCMLK4MsiAVYUxH9rkad+VMsiQDlLxq8bWMIlkf6+QZJPfFZy7Lo7GIQSRFRVmK
7bQkJx6baHSMJ8dXwocA/y+/rUi5C8Ql9VXZXtL5UiNx33MMem1oOZq3J7b36Cc6ifmKg8SqYXS1
xRfFZcqitskM87LyH3KJo4WxYihxxuoIm3fCp09hNTacojKxr7401/LJLVuALgfv3q+9jSVfmZKh
s9zbRYynbkfxRPBVcSIx6DKzusMsEEWpkQCj1MWmJRnRIGntoB5GUCXgQfPX7qAX2ISaEnJNLIiU
e/vJlIu6VxC4tfxptFTiCHYtA+xsVCbKmoafRZOFtso2AHdWsxZHI26MEWZU8krh/vtNDMewhg92
qRWl6DBYswGbTwvo3+vmtwXqtwT0vA/7vlp1aj4xeoIrrko98sP6hQ+amffShoHd+qXahqp6r+tV
fcA144gwMwU/1c0k2IoD15aXI3OlB4XCBF30Yhqd09tv2LqMJwBHymDI0QqAgOkklYsG4v+wtkpq
gteR9f4eRjtcBtbXyURFwy/lhklUWwuZRrQljBBY4hP2yLDEZuURPyHmBTflMXQfOdB1nMJs+PTT
xz8UmhdMwjLCq57mdHyTrGMQXCz6LGY+sTTliddNvlPiP11/7L4lH//uzV7cRr5gid689CTu0Jf8
1VH/4crc+X+kIDrdJ2AMmNrGiBAwTdbC2Kq0HswJ2K/0pStMO52Twjr7M1flKktPO0A+UVG0zPRh
HRbkiWVulqDTCtE7bsXGHUISuOJiN8zy+cQkDHDMFWj7AotiYNDi6hJOuxYiuRUS2VWWVtFW143D
wbG5OoWHiywuEzcalLBR4KPs1Gd3q/98o1GFx89kijI8zDQ2DjsqSX8YEj3iQWRAgpa+orMP0Ubj
nWxpZ0UTQUzGj5TNrlHFsccCEHKTI2FhZpPidZ2XtsqHIz9rNT9B3n5GreIHoTh6IJvAWQ8yvr1u
OLcrOtHwz+ZCTI3R+k+qoo3oZk0yHSo31uiJ7JuaKnmpMJdkb2Sr6XsGIcshQSZYNqZzXQgdO7/k
5D/R1Nc6Y6hKmrgM05Z9kZu96gzfFeH0//1Kzf0sWXxus7+ZSzbJ2cRNB8ahmUlAgOuweEOmbXZb
a9yqA2/ixDy2oJOTz6dEbARLsRUbDeZUmliulY/WK3lMq25loaQpVFJ+MCm5rFg9iozxIw3qH345
bagq6DJwew8NYDnP58I9iobuDo+nBbQ/6d17Jh+lEjPch8r0kxsCj2e+3ncSOA4ZtRB/SHa5GQzJ
YOcaDT2rlhPkGxcn6axcosGLPqMMhrtLFuHCdQ9HCm0+X0RtCFS2C/kB1xUG8VsGTgpCKsNY9zbp
UBQlpDRPKVPjwFl3GdJRAvasKI/PlLk1bhWXgzlT/WGFvOUkperSvgczjRk364JXeJ9Ric4Kli7S
h/eucjo7XtrEB5dQ6wWuuMdQrJW2Dp0MAbFwLxeVfQCsIxs8O+g91QDzByPbs4hCQNvoy+QR6R/g
o23LHBC7qS064aTJqJZzU1sO3R+QAWiIrkhzUJBcb+5B2XH0r8kZuU/FKaXosx3VnrwFPp1InNtG
lbsaAgFSz2jX8t4Q+J8NID7CyYFBB2xATRqlEXhQpt5tNgDHmMmcY027nNKpGZrCGQD/pK/LjMKx
sD7r3wzb1jm30qITRnS3pQP7bbvOkSpJtgO/ZJ5uUVKKT7NqTzVjaZba7nzOU5GIYD24FaiFaz5J
wc33NEayNczARrYQVRRMCZG+f/7APux2GNwtNfxo5kWbj6Sf9OdysdFAHQv53dvob0BHEKOj+rN2
M+Eo1LvPnKH6v4qK/RieUaqUJAiEkLLVjI4D7sLrZCp2eeIACahPaAfFnSOXJIcg9TXv98Q41Kw+
zYYgTJirTc4AUBujSegcFnUZBWILbS6oHUY30d/RVqdz0VozMmai+HTcifV26XhyVZJPoSTNZkYT
Pv+b/YRSkbjAKueccMgbhN6kXtb6pfgVkjLrjWUx7XOK1Mx5tamvHC6zhmnS60wLqusG5tRBnK1L
HNz27uGDXi/ZoQcVm4A3/9j4s1Dc3k6ugtwyj9BxOZcIt5Tnt0XU1jnXf8amyrIAfwZjbnGXQ84s
B4xeeMqxNBvbDAtDB8lsXLDUjOhLWfO4wFBjgpX7U9W7thT/Wu/uGMTZ+uPwmcavKXrm0xu+9BB7
Yci7cqCxP/+W44nX/wOb9ihITUn6kou/F00ZDcDvvSlVPu7Ohff6Rgr9wo9+utiLQ3IrK5VRuJzI
whQSUi2OTyoK10UxkxNy+5YOef8gi2YrkPWkCS44rin6BQGns69DBBBDW8a+B1PjD/sVI0Ih4nWL
enrduq3pLGwenhnjdgptjhoYkyr7EU7BfegBINPPRMo+DN2d3X/wMNAdGIlrTJOmm8pvM97wT1Tj
oiC5P/X3aXUN+F2mLE24SGVsDRUHQOExXsjRwshgZg9Pyc0vdR0A71rW5AhM30XqdqADW20d8wNj
Ch7Cz3fDaqaBk/Hr6Zk8hhSephMV4GTtCwh7GknymVtGeTQ26z96HOunOhyPKiMop1bMm9lWADaB
428V2Ra/7jX5vGtxcwqI2+PWhTp9dkH+DSJvQVGcgjxNDD+Ej3vW+XCBQOKHWzvaXjBR9r+ppc3q
fVd2pC2x4bkC09zYbxQijxFX1vhmNopZUUPyvwnUEDDy92nQWHddPDB6FAE7sFItF8CyVCYdgtip
XaJIUOlD85lzIKFl1BMkJgo6rNEuU2fi0GsY++MeicF3Rop6PwBbfNZSYaMe9vatzSKNVm8o7fRX
lXuSi6eaKA4TWJoSxeYNB5oogkJNVJzRVLBmgVlWhC45OE6OTuQnO3TNbqYjvHIhkNTaD8aM1EUp
UJvxq9oe66rXeO/3KpMy8FEzk1yRsOkDRWOV7cP+LQah8A8BFAU6OkpJW0qEwCWnS2ctwFKvxd8B
iDunj8S08QbUdd0oFabpyn3dM2Ny0n9it96KFhCa18KYsF6cghgts8yRrmGNXIFGoLLy3QI9dyNX
QQt9Rs+mtlt+Pi4rjbNrpZq4GcBGkxqjzFFHP9LotAfJXGCEy7YeseREQJw5DxaJH7pCkGuDUcsA
53qi18aBk+aWtLOBCLB1IiuUHxjtxyhv76Nq7T8tgqv4W8PGO64zrqcC8pdjxajjwbuKG5my396M
IBqJichg3pp/FRvURxVKgreE6JlvFaeekrFhzHhQA/Ux/mgLwFANDkdY6FXbMcXqCUakMIcqxKWZ
0ZgeX8d6plPfa0TWwA+qxsMahaAE1k5GcWizxyU4DmjCoyUE1GC9wgXN27owBGj8MnU3QF4cOLE4
dg66/yWT6Fq4K1Vo7TSjO56grKgZSWup52O0Bc69rY5oib4WYY0WUCEtrA6rXalXOJKZIhSBj/5q
1UF0HI+EFIw6JrZb4WlYk4pXm9gYgS0gkIPS2ZuSkOsBKkEyaJ9q8m6AJO+Ijv9OAjA4z8RLyaCA
58jKZrKvO/++xVlgH4VFDv39YBX3DSUZEA/hvojMuJ+wF5L7z4TUPqAnp3eL2jLJ+X+A54Jfhwd2
cHeSLMyEA2jB3jF3lHOg9YF3qbiwaLFL4xSMUgw6cAkQRvBNObAKFwD/503m6klKhoSWoPYHD+6l
6bE9Q2BxFXFC+6joJRuaRmkCkDsLxtXwIwv6S2ZJFLkwYRw2rxiKO8oqJh+YKr5LGJ/j19iQHsSS
Yeg8hIzYbFKLdkuqduyWiRwILnVkQQuiI/7s8LRYGz6H5WeDIHaVYQMoWoyLn4AcKhf22pENQ/iY
Z4NXaxERoEeR9Bi/pPHiBPXz5xPJNk+lmU8VGUuyiTNxEqoc4sbhDWRvn2x9xUoj/GrHk/JemtiW
+qoW9OLSMQZn5ZGd2wq10+eLbGPQscdE8YPbZXsu2XrPj20zLAp3Ahjy9yIM+QqGNb2o9tWliUR2
Hq1FSy8kS5YNsjCwWUph08vLMQz73QKkoBSQMReqqAH72TyDPdqkuphQcKrR24W4suX4fZSx3Ru1
98DaS5FzO1xAJ0DdxwqyT+Ky8tU1yR9x+tRzRfD3276Y6NCB+UESHnaPArR4Qal4aolxDaVupnVr
1pFTvzdva+WS1ZdWppQLQBZYGJ8dHYXNR5GM+It/Cyzokekzwhy2OxdevQhVse/YSP9zz5Tn/ww9
SD03Dr8S6FBGJ600e605Bnf//8g8Ko19NmP4PCwCRue+71ARyRNtHindzAUrrX6ks8W74+pmXF2y
sW7L2Jl1Kt2p22TnDwbmV+1HTLfadjk2w7wfjPHrFq8ubwv4JDrcIGCGA66dmG0ZGb0VySOKQQyT
6NnIrrXotkEdHQplPfKPkcG+fjdjbzhti2HTr17jf5M6BDczIXMTmmAmq9GTNFMGqsV9dxGOVOgm
zKNvkdF4xLPfR82IhvUzjZFy7kyaR1AMk3qTkJP3aKUTx0eIiiE41KZ7Np8sYsd4DiEMrsVo4cfL
MHSnc45ZDszK12T/dYaP3D1Ardrq2iaRBSJFJJSgrm6PSGyh1O5uIKNA+bfQFYP7zaS1GxA8lPMl
/QM2pF6iVWGhBjtekwa0foMYQ/dYsQYJdOnsgxYRsQb0XG+hQRqpEwYA5oANw65a3+dlCP7atYNe
aOPktpVJgoWeu1POKXSNv2Ng5T3qHNPc5Ceuhk/vRCLqFI/HCYtZMoXVa4LO748fxwaWLuSu0pq7
n9inhODGMO9KxzO4W0cfi5wkElWaJTJSiAGAKXPu8Y1y4dPveZBsgCLcTFM4XFv1j+caKYJ0Ft8K
d3+VoKRXr2pRUPoNEDAxdxFTWyI04O4D0u1NmVE06OdhDn3IOsYY0nnD4szMWHF9cgcdq6GczZRi
64QVLYB3ZyYLP9UQ0L7vazZ8N8kimKlzEsFxskb+kfoNhTzzKCs0cJ3Wv8/BPiYJxykTp5LZBrfR
0aFB5PIp8cAgJWXDEcZ9IFXZAo0ud5DUC7J/wz3SLaPOImMYHiWSWZZ1cNqSmdWuHB1hKdAVePTO
vYTx5LxwcMj+CPmnvrzCvnvANTyGK/GHG1Czz8QAR1D3pAVo7/uugNXer1JHWMLjmRJL/1Q6Tkgt
jzbSzJNdlTrBPn/9Eq76f8qMsmAaleFQVmoWhA5NOkLfVZjm7z4tcu07ORaYRzTwSn6fTMeYf1jJ
PoibQfKhIaIJT6dwkyjIQYw4ZckVklAWTbLNeOw2TFlSCxkIANDafsoVwtPHR7klVUoEJnBCdeUz
/MHrAVeImg0ZL51l4kYwa5aK2FLtbtT8vmuWlBqysUjsx2NVGQBmBuB9AOYsPSXHhvvn8+ukkIth
7cJwUVQgq463Isbs6HHfck+WvZMav4zx7MEXOstlAx6DiqwvEskF/RKN3/dQLA7+K2tWBtRmMS7k
4D+kX7wtE2BA9ZSTqqj3iIkKagOdOBYXjYOtPIewvKClS6M6VfRFdJ9ZEzx4Glk8kXcrmq4u0IhK
m1kTkFXk0gM98ZOsIF7cwHYgXRj/PRo21vVHoYXKClz93giITnjxGqzGrtZcfopvQyuCU0Q3qsHI
8tLIlzGm0Z2ExYjYBOBYBW2QAYTvx8FVdfSCbxM9lRVA7l5zdgYSY1DiOAe/6eHmOhSUsNiLWbOQ
vI6/5QaJpTsmRipcWrYUnxFa2alUhU8mJi28w24+smx4894fEh4pjynpdtv1IIsvPHvLvCc5Lpy3
6oCpCj5J+Hx/VwpeP+GIZ5FKERVjbpsUNaFglfi1P7mMcHszbcXrKEKzG78JXSfFs/Dpge+JQDWF
dK2nVl5/DXry2ELWllBXlKgCgDdzjUEvEDTar14ghEK58BHR/8ycPKHuZ+dTAzvV+TAtzgZFmbPZ
q+Am4kIT/kf0wRTor3OPiIiZYLcFaAmY+RbPb/moElZSbhYSX/RE6vG+r3p6CB3pA5P8dAVFxd1W
a1AkW10RTZyiUzs3tSFG9tIGPy3d2lDoJSzJyKofDS0/ATHQDLid7aT+VFmik1tbYKtkyfrKH1JI
oIN2RQqRnT1IUdAiYX99uvLgrQNLtwtp099YucvoV0lhrvE4053xlcCnY2gkWuN4Aws90/eDBv0X
2br7aRhRveaUgy5JFWqUtj/O21qOFwc6+SXOz+t02CZMy2C5iUO6g49TLzgBTkN6+p0OwLQSJiL0
AR/LxvW1m9212JPLcrS5NVQaaf7kTJNChXWlYN0T6NuWiYHJDdmnwDjEwwNo7EOBzJ2KcFkcKGWi
kc528Ic5T/gTtVmJ1DXH3M0Mo84gtMni8L84TP9MCzwCiv69WgfxD7cSnbTRQeATeip0y8MjSdoH
M/Cz3nhkPFY3s0eBTSGLYla8xbnfke2ZvyZWEyapfJfBdZnHKHBY/Dn6PYgWKOpcdUbD26wAMFlU
T/hjds6Xdk02sQNv6Q4pILwGlp76wZWVDy9SCy97YVV4BJHIvcJaoaf/O4wOotdNulCI3APsqBV3
00k6S2IU8AYnagKIGPQNu8JS+T4HL/eQNaxDr+8lsUTxKZbXAK3mIJY5O3m+igGStEDltp0mAzzp
e9WvrW2XWcjngb5ZbkfNIGyzg/RHGgtbNNIIhxco9PFGKFDYAVsrI4kz+c2KVCG09TtPEUSzCrQv
UJ+wP26SuGPtou78NF6ekgw+3y4LW2KL4UUNxr2ypD2qykr5TXWkRVxE4Wxsa/uJmuWAhKxFQufu
Omr0fTE9sl4kCAGL7S4FNT7B8zmNRJWbti289zkZGEfFcdn5Fjuv+UjFb9z67m3oFfbeTzzDGvrW
cwAt1f6iEDXoyz67c7wD7inrneintIO591tyDj4KoR9PGEl0HyZd1iM+MhJSE9OdpDznS75nvQws
ShOENRj55hyubgk9/cS+KrkvHG1LGaZTFZ9jXY+nwl6Ll7CzKQ/EomKaixv3JWrOpNJJYljcKwJI
S4IK21644Ojez+vJxczWV0HqcsUQT+erffoU+dA9Vzt4KuhZ6HJ837+/tYNvHBdU+uSEkeIPqsN4
7jDPCJi4nzrYDhlaUg+X69olf8TULzxpvNYPvj9z9zuL06wZRu+c2wbHL62fngls2Whr8rfgFSqn
dVR3Q+pIbyugHnpvSwTgg8DDYmboOlGRn+VSxAEVa4t0lGaZzInYrFXtao+jAbz40TpYCfrrCc5q
KwkiN7aHDE1s8izD2q5Fvye5+W38oZzQtsnhc/rmcgmoBWg4zYuOlpiFHn31Usfuzp93hauJCtTS
lPpAw0zM6RGatLE9QsTsAFfLgyxCrOdVQWC511amqxeFhnO2yqQL1HF3Hq86fUVgUQAmWKQ3z8s3
/LP11V7uih54iPlB/mRny/wccf7QbJgE+6/izgffgupm3PikCqFVDDY8kdkRQb/vSp/St2ZH/8eu
Ya9UyQIzqmgnuHTrWeTamRwAmE9NgG0jYsdXJKrAO1SoIXoVR/1o4JVvRHtInB91He0dxptO2uSX
Tysf+xwm98d9kzDjY5DD4eypVlkJP+xaEL0RELpSoxBPOOyb90edP5r3sFGRauj8Kkehwwqzo4Yw
jLa2DAzadvXNAJt/f9nHrluxpJ9yxcSkAO2omVUsrJdXNPR4hlDgB1J+VC+jsf87hY8RdBwkeAu6
QBwzBPTzQIiK76Mhc3YCam4yrSOQllvf8ItbOgkQfUQzHj3Gd9mvsqvyMRsAzNHTcfTBX3u7lKPS
8EGsm5I+78Lgsnwe9O8fmCUMt3QgfuZejgAF+VaiTwOG4qzK2gL3XC674gYWuO3YoPKyWEM3yqEV
FTIFV+B+Epx2+qh/mAStVhH3Ir3MAh9venoTPUeB1z8Uzg+TlcvcKMQa1Kd3Gbb2hH1KSZIMiEzu
c1WT7ZNp0e4LZ2dHtLyD1heRw1LTKcX4VVlYUWUd+uFmuyHs065/Gs/yErlzWtXVvTgTvJQmF9w9
uChqXH6p9Cc0Ur5gAKUlp71QiRTkUgavyNmrKY1EhvypnUvfuGvT63jyN/NKrWujNyG1jrhUCXdO
H0TOZMDWQ+SACg2VUwLIABClGwmGgp0JEC55/rAAeY9V08TvgqtWeedG1n35gfQvswmVwt99tB+N
CPTJl9xCUWWkzMKdKnEiAGKirYoogBTt1HOlv7CnnHPmdflYx4cjYZoAYDxV2/7SlMWwEeptePAQ
dHJ7rN+XaTEIfRmRJLVJO6ecAKaDAcgOVJcVyRuqLgRRRwHvMOFw+T7vo/qquuEJwpQ0dUGavVDP
Nf6CWtJ6/rnIXRXJmaovgJMpGY4XDE4YHp0a227BInyf5v6BEmmGab7S+OxYk8VIAn9kL9sxwele
ZXK/GspIUqjd6OxCafg+9FFYsgf0cgvZyJXr6tF/lTYLAXFwwK7CdBH60Jy4qFJcNjz5XRYNYlGP
M7pHznktg1Fu+4vtkW3cZXblOQ2SvuosrQjiHyPGkt1PWvidKlIudCGH7i8jAbvNuP00DTGyckWH
d6ldwGFj9B54groypjjhyFBGZeLi1ypNWRDQVMkXPtqMgc0UGfpVQoQpequwEUz04WtSdaZbJcs1
bmjstfo8oLCzWLuzag9d0+RLF+BYWovKQfiuxPdgdh4xKItMWk63pb2vrqLq+LSivYIeywe5gxS9
frbpoDVpr9KWpBOw3kFXszeHwGt/KbguarCSJp7r4sCnRU4fV28V+LyZ706PCpnsZjAJtQwUHGrq
BUhXVeRclAabQ5y8bj6XxOGfEP52Ni+jem/8JSm1Wlj1WIz7TMOjT18Ce7pvarw9lrKsKjDpMnpg
Q6yr/SBY2D7YFdpF3HHMRndc6qGS3vG3w3OVwadNYyQzHJZL+2D1qhkR7GF8A4UnHtXhICI/A0On
qsbiI1XG9yoBIzOYSNycB/6MkF7GBsryVmvI5IrHYXa0/2quKf0buaW3TpbiyhF4/8Z+1CN2yk6f
X14TXEPRCOMwKqdK9NE5aP4JPgUY7cOg7pTHJ2he7kFGy/y9kHGJ0eueTxXQlOJq4p3WiiGiOsbr
8j0HyIGzlWv1CznrtWz00p1fFPQ3c3wSnWvd3qtdHINLtiooOT9n7rsTsNYK9MQh2uNUtstZopcK
Ibl2qKBEHTB8B5UGRyZu6solBBlAxEbTdWb+j0MxL4//V8yMoCogGT/2rxkW4JTPrx/BExk01DE8
qTZ7o1ruSZAqUyqmLu0WHxSqMq6xSL+elbjOb8EFAxoFN1pMPK+YMiQDn1UVB4olxHj4hLc1E0au
K9go0sy/4uNfW53XAw9DZM3beZP1a8hEY4YEITbryoN5fiv45eXxqsFHOPSRJpjUIQD7Mex9kZ/I
OTW9HJ1pTUMH6s6A7sJifEW1I0LHiZJ8aIH+qhZiQ9pG34rGOj1LepHFgwxvDPf1/vS9t0xgGizg
y/6MyU75bnNAryu7ZvoOQ+e1n/WDQ78Jx7CUq+RXZmEqgdIK2VgqkSXoa+rM9Ibxs8wMpNCxzUjY
643JFvnr6AecKRIFFaURFAx2e1xQxnkq0RaWyhZBeulfysNalx7uqNqsRtHspxt4yA5lsm9KL/KJ
0xgxLAr3KgG/j8b+5o5z3SfLeN2w+IUWZg0DQethwUMIf7QOUZjFR99sBulJKEAFqZRdSaB3Ybxv
zyf2VCAm/Z+y6Cot8GF65xZig1a4dt5BS+oCYc7GIoBdIA53M/61Muyf4j3L+PVuMoa7yfFyCenV
jnd+E6FuunM5Jshu2FCb11+RUw9sLHAIma4ItpLgT0guaLVBZr6vpZ8Ux2hRzlJXKwbtoCesVuff
w07sSrvzlASOJ7w5TAXBZEiiRoMUdKZYwkTJRJlaSD7MYD0uEV0Cx4X/vLd82fAm2Togcte7zrMP
4hM2F30dpqm14tDuG+OLVtQjW/3APKHLZcGztY6f2eM0lW1LZTP6uLaFN4VvtghGXGz3ylgeYc4p
G8IwUCG2b+msiGgqXD8WJUAO3JqV9BPipvbo2CEAsO5iWKIfwkxh3NEA5oZiP1IwNy8zNbGYuofF
WzYopXpA+VX6qV/uJKqiXzOmJBt7WSvgFhfqxQpVlT/6d9dQGql0CH4uwTTRK0p7ZbVq1u5SfVzJ
q8r278YFhncQRrv7RhUyx1qle4ZCLkxMGbyJkMXd7NQanPkN4VgvKOnKs3da0trlZmuOH6Uv75FT
GhoR1+9+nHtOQGKXr/LTMa3pcmcStZiRKeJRXnz1+BJTjhoaRyaIwdu1od4VFOV6GCFXAsn2vU6+
18wAwk9Gk3TWUf3wslCj1ZKThBONz7WlmayJHQt9c/cj9MAvf1zKaKueTV3tU2r0tKuPGK4+H6se
lUFNUqnTg+0me+1uR/m8hF4v7JZRMDa4L28REbChbMbTYEapbSIqJuv9cEfhX7vpnu2LbsQZ9jhw
l4yhLdtgSDTb1Iu++CaDoiUh0m23I7lP0pS/HZB1uIdYPyQwLpWjmY+2A9djVITwJpJbn+BpPG2L
fCJL0CkLeWyIkbK9ewyYmZoi09LQ2ACGDxAMmWAs2iOicKj0LtL/dGPr+vH8RClDQhCHJ3MoYvNO
l9vvfcs2mebIQH8CxdngDXYHC0IfJ3A4sVnKOvv7eZHylcvpOf0q8MbwPX3Fxtl5ru3GpKajcRYC
//LIaygGLmgUY/ICKA9eu1v87wnF7uonemrY7HoDWWi8002sfqYe7b2lo75ZieFHcMf+fhqcfj0o
PJekIfP/SVbbpJS9l+3UztaUnXL3WBs4jhQTMA9rqRmTO5N2qULud5LAqICEsoefPHuzUbQLD/TA
bgpX6Kv7rR7DmHZW9yM9+ojx9cjkHIwdQKmHqrgV72UtBuQQdzMJTCmeDNxzS7Osf34kuf2SMuLa
A8T6crLAxXYvs2jkA+Pc5Xp3EqcoZPKXsB9uB9dFGHFsjZ+BlsNY+2RauyJIdZIVtfYkZ4X0TIaF
ITv/t8x2hg/PUNCenq7guyO/O7L7wI2saKXOQ5mKE46nDBf8rOOGdNWcG4F/NdThPW6fuvejqani
ot9O29ZBIfvD6YpoinIArpAJwGZennKTJzX2XIgYIMkl71cA29efDv6uKsPvIzWr5Za+dLqwWd62
qHnCWFTSkjfNodKjHAU5iVvWxfxZRufXTEduagciJ/SVY0213BPvhqmkU9/LqKQMIu3jMPb1w+Yz
4/+6H9k7C5z+/a5dzkB07EHrCSbvTf2PhqrD8icsSJzGKViS8kaA5ffmbkuDpK/dGy1xg/86b5ev
shFfb16TxUp7fMQjN4vFXE8kFJ9QgfBnfxntEKuHGgB6FiYvRy7bqEvz9Afk8w79Kgv0dnuP/d80
t2kVGBhl8vVNJf/Fj/Rw/u+o7wmXyMZFMp5bLIesBFl/aNOu5F7OcHsRT5FLBQYbFhLX6oBj0Qb+
JCgPgnQ+3UY12S9/JrXCcbsrFeM28iiUVsj+IpMZmRoHJbjaoVsT1vGRXlRjPASQcEqSaP0ZBGjs
xXfw2blDxqSsMAc0FBayyseTLMu/XdvO9EkrDXjKMuI1ahgwVPCNwb9RRFqNJdidXw9FkqgWquQf
sZCebYX50TVUfoMuBzNxyZ2IJHsCD8wGPU4L6Bjuc3AVKmGX8mQRwNFfn2l79vEPpsB001ogxJB8
ImGzl9w4wPhFDre5hdN1vli3uWuwdhjzwHEre7WML8MGgom5nKaVyrCBGBqvxCr12J1LgFOWhy2w
lbugZnGpmwDiwmoGhXM+ouvC+9HaZD1zQi5wdEIynvIPcC3tIcDDdxqtNTX7csghYjbmdEOG0iHq
ThhAx9BV9FL3WpQJp5BrUjGfMRHxRw3BYlvxd2jbNuBaR5RFJKOhps8uT6l19tRMqCKWuuGiDO6W
+kjJAlNlWHL4GPkN0klOaD/VEEA3IAlfX6s5OGeoQ6+bUf+JAOJQh3MpRmesaACr3xL5xx+UzKm5
WqXkqvPzKTyGm/DNEm/gdhMJIa77wNya+Otj5USi4EWeQ7dvyKv4SRWp9CQTyZ4FFWZQdi4O7kKt
WryBbGUa0o5K/FKlN+WSJQve/48n6bL4bj7N5Mc17pKQbmsCE0Jg0PD/9TEfcYZG6LZlBGTM36HR
mKjcnsraojyh+PtEMkLc6XyHV430jJWDhbN4G+gx39caCCnStmvi7WH4kD7NezhnGcopX3hY4x4K
duu9zOkvTSZ9hH74Y0Y4W8svkap7BhQnkOxMO9PhNH4FJhjWs4nse4eBYlJuFCn6e5svjBdIUd0u
khxr0JAkrVFKwQllTVDP5cbNDIJw2es4tCiVNlkv1ACbqWYqFkiYo+AiYpLBuDGA6bvtammPCuN4
7Xnv9m8JIIPAUGUDrsKsCmFe8CtREBUALPDq7wQ33bTBxw15Hd99qcxkxzZeJQuCXPlYmuNFfFYT
dBSc0E3px3fboJCdCox6cBt1cosT6yB6++XznOevtIMHcbcNZ2YXpGnzcAxtQXTGsNkUEDaeT8qe
szQ5NAgRLgvozHaymB/ppm8ezHMeif2qpOSdJqcKaTcgVxJK4vE6bIEnDBxKIuHUUwepKYbOF8U+
N/B4eh+F34uPmzeOeXdIMyad/T1ggj2lbA/6VgomxEK7Bec8MSiUvISwdEalYjTkfB2f2P3E4iad
uaC/jzKqp1Ot0f0kSr96R9Mo3JIk1k7RXR7iF1rIv0FP3X4XMbKo6LztDk2Yp9mAy6tiAnPPcDNv
7IvvJr+yKn1VuIUAEsx0e5jN5oTjQrfZhVwHFu9RsMHmYyrqKbgDicfo5LjQeaseFu3khOTDZn2E
i/LB5QwSkJJvKAYlb+oIuTI+CQauC923hGo1d1AZfwvfEPZs7nYMsbQnNTBYS+WAxo90NB2KSkJg
aKpVPT+lLcQcguUcep/6lM6XHIc6Qwj2fqaD2DQtdNacx8I7eGypY/O7MbskjQhfsrUDQKhVAuvC
ms6lcFvt9RzZmod5gmLfnFTrgTXc0M7RuEMHgNKvzxQ1A+HoXR1QRzDpBM9QywEQtVlzTfYxroE9
PHO3O6tGdXYfx1DtPnm/TrMgEsT5ee3Q13n3QCH6AV+Z+BizgIJTj7A3qFMLxGuqQBe8YmJrG6XI
ZuSswYXhHKOHujKaVthcgQsDKYg4STrxK0hMdu3sVOqW4huNQxAXQ7cxf1RWCap3AhEc6LB+r6ci
weurGXuSm/r7fqKI81ck47ugns4BqkXoDWLmCJ37+U+uILQpw8ccNJzjPw8x9jD27OWh090nE5X0
cEt76CJro9OQiYSNRS2Z7Y0kPGG+U6anrf/5cJt3bQT/wD97TnH4qB1A4lOsQLq0rNzjGl6VVqXC
3/jLkuFdKJAeoOEFLz6KRjtaE7HMEF2sSPG0DTNh3wbZgpTUFN6JVKphCCK2Uej/Kd5Bei7Kycwp
m00DlXjyHftGxr9At0v5rmBLfrLEWjzWwSE3kFwRVjp0wruzpOT60OKoYzAymJ455L/MdgqZiJuP
FtI+JiBbokfWxTGaLE2eELo0S7LMpBS1Xtcq2jGypV/LyLvUwg3ELONpw26cm1e9yw/eY49b5pR1
uBbz7M0A90v/33y22NzQgCpiZ4VJumNmIh8qRMck3KuOuganiNd1i4jzugkpPO9SI3CGnh4BkqXh
SxNI2ARyTppmd7hVh7Y+HOdDk7ik0crHRsFaLPxHXts7lKAaWvNAUnXX+hd2qQ7vulC1WlLsCBPl
wkh0V5JNNiaao5XkdNihtvx+iAOUR3+lQBLtLr7BCTDKlinpjNvSLDA3pXr39KIWnSzYkBHaoXa6
/5IyTx2o84hpxJ+oC6bj27jSBvUu8KaAY47TInqOonORzGLJOM2lsJQYYlxRYjrtlZ6xqhs4fZrT
roojS+qLDboT9vmXsuUY/l3tQNI0E4MChiCgzGCiHnJ/7tMe+Ype/qe+RcWPuSRQjgqbpChL5k2U
RbJOYWHHMSbtvsEItlIoS2H8lssdKu/OxJCLwUW8aGDdgyn1fkM+LaBAAWyIQdPEGuTyYR+znJSH
dml9SkUBX6qmmS91oGGE//STjMjvb7vTx4XMYXJlXPVx7whnGuIR/RtRr5ElJEgeO8iRKacN8M2L
4SPn0f/SgFYaxifBqXr+pU6zeftZTdhV6w+hnPa554p0PL5gNlnrcZajkn6o7FJ56etzxbo6OBzS
rvyhBrDzpUSM3SRJ39Mfdp24Jl9ylpWPU8ShG6F/sByGfghVCr+pRKdM+Vvzi2yV+JJ5SNs5sXOS
qCUPU2jIPC6JtMHzpG9IbgknrMUzI7ZS9rWFdLbBBJ6NbgQVFztbog/rXjA9GD7Wf1lTDZeUnQLZ
gHSQQjknMpZ9wcJNU6liOI+aXV7HD/vBD3cbLdWm8NgUuiOPCkAzXrGp1C6nHXiTZX3o1TQVa5zy
8GMXhSn6qC4hoTt8jZ2JUt8r3vBepQOzKCU2BxcYLIB78XfdZOZe6Xgh/SUxcJ8Hd48GNwBfmMXL
KScdJb/GREcyiuN4jshMBcruYPJSPOlGKnZWbgR6RSt6wIiyXb4Lvm9T2yjOwpYj8IwIXNytbwXJ
8tegXh63a7VUqSD0prtSEPeDLwA10I5vuryUPGMX6vZs/HkndlRHiHYNROS7qGgCFonnuo7enm2r
8wO8YdYn8KhoVFbAXo/lGIeASxZyjOa19rorgDrc66fAI9XOfg5TtDOUiJ/JkHcRh3wkmdSCAC2s
HmMThVyvJ/raTcNMhvD3gkPih4xzTFxDWrCkbmX1wX3SRmPOAuexu7e66Tbuwhc0FFoeLcZmMLCK
72Wztt3dpqsIsn9PF/c5X4ZFodfzN/h0U4a++R1jm30LZ9BV8ea7/Kv/YTX7psM+UWbbgoT5kym8
wmB3ywIQfTxwx4BKgOcWdSki7MWHaaYW4hgfEAAafwU2Y98zhjmrnkYck7jEqBs0G+czxLdjbraP
rcL+vWwtZmglwzQ0y9jSBkju/qiZXXlTRKBjEZ2X4k1zmBlqE8/SN9kvCVxoeLtfmE/wATvdq08m
PSipnI/BdajEWXtavhgoj9E7XTfwjAkG2qymLuTcSy/P6de7wx9kdfITPm6QhrkaaNSazbzXP5y7
sJYYWA+xyqde2fSwk5S8uD/qABs+4zTkMDJMGqtc6vMq3MM5kM2wAs5WVb19+pS0NBbqn3s0UvYD
UgzdyXWsJC4BJwtseacQ6e81402dWAnSCfx4QWXAirzuGZ7V+tz6e5tf/lXHTdkACvbLKOROT+Cv
DaCqYIOO5WkyhgCMGh+OwIY7jaZ/2UFKTG8eLA2+G8jYqbaNvV7WbDruRFlfSzwfvazBs690VR1j
HC+M8rhHM/0SckcYOFtYc9Iva1Y14uduwH8ZZDCFA44Uu2FzKZY4crIs2ln4EElwTKJ14oyUKo3f
bpMcNFgjB3Cq/6Py5o9npG5eMgusylB47/Br+0OULKaMP+JwTSnuKuQ3gf8mE1Wp5IR4DX35LnsR
aGpCm2/PnpgA0nSdp1a3QSVYSkhJF5QW0hg+hkZvbKOKuNIZK3pxR7pro+Q66zRDgnHy3f1ksfzr
/m+4+M2J3dMLnMGmobkIbbUVe1PbBQTQZHOxxsdnizRlc6XUT4znYtrXKl9IOEfQmSsfRY/Bnm1m
kACA82NCGG5s9yc0wf5ZBS93s76YthxwB5ImGxaahxTQZvvSM/pYn84vQX7CyhGtllerNidydVIC
3NcBTmCZcirqJnMD+CEPbu3c3TuCuOdaM9HtGHWVk6SEt92h9/JhvfS92D49dleAovm3Nj/Nm02h
O4sMaUk+X9YYCAgcSabB2pbTaP3MYJLl23Lv8DLlwxdl7iQr6HrK2tqaFsVlvtTK29PwMt05lbmo
u/YmfhY7VY+8gSrFAHYAO554abNfQDqkVeQNGYQO1jPxh41GSIwC41WxDflWIAm7xPXFU+QXXh4P
Nl5Mi7zr7jE1ZrNPcuK//l6sn/Wv1FRWhXHPKOJMlTQzKzpwdiazfrGd08sX0NUZb1srvWLYTcPe
yQneHsh63jCIcc9Laj/0uK517vDPMuLj8A8Y2VmGTBA0Dgf68xklgiIXhGkuNnIRjMMbLdhwbkrn
vlY4TyP2CqC2UiRMj0cxweVa1xcw7twVzwnhL5VuREZsn0vhJ5RsuCebuzBOz3Mk9t376PD+K/ft
KYfr2DF9aNk84Rbcbqr/uMQynD/9j7BrE2+MMhVa4ZGAxtZ5rqfg9XI0VnE9QSmQXeAnW+9Tcv5I
Vx9HtrNCOzBNfS9ZhOsIEjN6myS0Ksnkmly0yJM7bG81pMTa6zbHf6gNgdafyavSHQ4boxJka1p4
VJ8CDfUBVdo89QAlu5lsK+nGkoSkY4+ezYqe0PccfTmWHTfcPJX8sqpRcK9S28jsj8dfUKKUrimE
p6PydwVNj12nzSXl4rOcu0Z/HAduzKQsrtGzNTMrl+P9g+80rBzvjsPKLnDG6PadoxD6Ut6ZZfEL
AVkPtEX7ugWAXV/p+M+SUvDSZwV8XzVBH7+gGYB5W7RkJuyDW/5G65q7SDBKWpojJXHUjMz/qo6T
Fw7skZ72uweJ3klTr8OVgbyzvK9W2hWbm7K58f6SiKXUogc4LvYawQCc+thA60sng9J+FpH611dn
HINicVYz/D6+wNyVzSk8fRo/s/9csNoncLdPBdp7ipsQ2o7+1VPSrLD1jY5RXsYY+WHp0onnvYIE
oXlmbSTQSQFp0FpgGWFU2ReHRDqKY/7ZVl1TPA9K2BlUkl1EX+sdQTsM/zPV8vrcz3JYCdN4Qq6s
wvdKEg/5RCbaZmi49igu/p7XbakUeB0R/4ZounkIIgzDvPiBfg5nfZot+Pna+cIaxqStm0Beb/5j
0vbajLKWqjha6bY+syJAzEcebeen93yf2VlJh9uAfIxpYfxHx6Wgj+2rt2pqFUovoiRY/ywkeGao
Kj+cDw5Mdgl4snMal5BMEnQSXisKgpJoOEjtN+nMvo6U868eKO3aXA/2nYqDflI5kR57ZAk1kxnG
yFX1DhHKBZiDuaKHct79/de0SOuuVeWGD3mCc59ESixdV6Su2HPZxQv+o4tZaTq2oapBChnBNEPF
cOSRViK+scXsxxjcdg62QdaejWXoDmS73405m509Zfp3AJZbyBrq2YPCBLMamHvcfgmOMMXiw46L
RNQHRcq6FZ85pKRXVib+W/pMOwlqqxbxm9aY6yKw6KT3FniPliuiWWny/+g4/3xiAewFJdaXjuaF
Sc59/nV4dUfEbZX+WQ7cBS5+dw0LTXrYPu2K6bExTlCoK1ndN40o/VYPHuQ5d/+SfjyzimHi+JfR
YWX+En6zfw8lxvImmg5BVX/f541k9cktPbiivqT/fS6wL8TtAiLg0Eto9fM3+20X40AClYeLMjoz
Cr7nRTU3kWga0Eq9qop7ZtyfzijYKwriMBu6Auh5OfvmlklRyBjB8a7tgyh8iF5x1AIp3JrAWp0Q
I4LC00nooigKQvSwF7LTDP2NTEaqsIfymjV7yIQeQmHATKoUn1bdt9oz3HPTJxVEtWae1ZTRV3XJ
/m+LZaDa3HYXr7ymwLfSgcPVPXb3cxp+zdUpn4uhby8yjQTgA8u5YQ4O7F1Uklp8OSZsxWoQ40Ih
YQGij5/7sH5YreBJi+TTBW0Bpfs2rn0ODVarwQTG5V0DiJYczTPQjuuVdmov7YV887RYrc0lNg+L
kfn18wS/GHAwiWzovcvjSm7kqP3PQbYov4qXrY3Xu3DOnc4SluIxhNKIW8H7Rb+GXFsAXCp1oIun
F5ccFYz75dTA2MttulWZq1xMIit3mgteP5KjID+ZVCM+iFT4903h2mpKkm68bZzpK3SOlQeOIXyz
VRJ7SQriC7nDdOfJ3pTEGxghYjZIeBqq6oaRLDCoiGVm8iCbDAdb2KL5vZwMvD7RPINcAS0H81Ng
fjeJITT/WKQzCN1wWmGo2oQv/PFu3CEqhS5AV5WcD3s5N/8btADwuwx6nXY6RymT0BMP7ApKOi8B
485CZwiYJ7K3RTGkcQc2owJI6RvQ3hH1gHL1b87c9KD3eYDTUgEYp1OWt0zARPJdV32eb0QurKhM
R1sRp6BQTO8lRKdeQ74DoXj9XvR99boo2+GkZrz5aJouW/MZA1rz5bu2ATDqNgbksrnq9z1et5RC
HOA507/wWWMaxkMml95ctqx6ocw8FC2ISjkSyBT3PQIx8CxyBp4yBCfeVak5qIZbXTkHUzs6N5xY
xd/Nq5wklekwG4sDjCdywR/EbNVGxUym4ZM/Mde0Y/EqAj/+DSMO7KqGh1FyF832AOqKgXfH1Zm3
RvkasMJQhgBzrd4QQVCR31WlCo3uyEUztvba8iA9ty+1asfu9Sh2HkrbinIYPZR8m45yTXmEo604
dCRc2MYqo7jlADk15/pfYHZUbsD0c3TObxIQdrKxWzQTLYFxCOiLXj7N2NkDgMIsCho4DZI10/5T
WJTkbi0LUFM/7PFuh4b1g/2RNGnQV/F3UQ50zUPk5dGtIbDv4RzQn2tQFnpFQDi/+DzUj8HPX5Hp
Hh26N5khcLZq3mK8Y4tIFRsDH/EJVvjmiUm8Mrd0Hu1QtzroTRFPDhOs8H4TCJmIyK2KHGaPYruT
xOLVmNU9y2ad9+qMJLfvHDQONRKJylQQ5qS/DaX7nXqqvvS8WLDcWOXYdjE/HcUoGx74fAC5uT9s
1utHKdtoRIzp2CpDNgpOU2qBA0IQhCLl1doAV8s/4R1i8sbu02UKStX7ytJYVvu83IPSrrZ1Vm2y
1caYCZgLgN2u8IVzDWOQvHAFsdag4XQNz0BERWB8eNhP0MYCUwx1jyEfak379HauhMOrhelIzgDt
P9bWYTYgLieN3jw872BFvcWJH1s/1GEFBYJmuOPRwstyMSTt1zUzFKedEBDb5Y5+jPPM6aXj8Wup
WPjmwWPY+W/SrmbxMC2iApJrW+6oX2oorinYMAXfRthfbtVBGSuDAGECtA3MYL1ksGi3upo7/cSp
zujZf+Mb6kiv0mUngCPR5+h/9VmCdjZP1cfN04nLeLc2MRsVPxTiOOvFf02OFqFzKa8TShxq0TMq
ykxmGfV7hqyrS5KAwOHA4AmHDg1EN95Z1viU8/Zffy0pl930dPHZcnSJILom6gu42wx1pFmiUvhX
se8YP6Z5xoyP0rDPWdQBA2LRFAmixnCNEpNEpaNXwd9ecZnM/jXOwthcTqUmYKaXpnFg+3H/VUTV
j0gCsnCJt0PYnWX64xSWLgIpjgQLJXHrvOSsNkIZZP3xzInvKQNCXc3HYZzs7dwQOD7MTOlCG7mC
a/MG9FJn8ipR9NCeVvANIUcOgOWsY5sQfMUm6Bsn87XCT/ShIlcYtCy5vTvDByGwlLUslTh1um9p
hTeeJdsZs4qwYd4jzGg8yBsFlvQj4VJQJZJJZmZWDYGrIBN0naY9xDq6v5hE8ciLnX6ih1K6x+nf
id9rhvn3JlyVT8fEHuNHCaMUMBVHmf8wsybxhIAjTJggWwtEqd/8HXZ84eGsuuGdFIgnZKinFmDY
J23siJO3mBGqF/KQHUDNo2rKM3qRVQvO0wUcIkNMaEiKSK5+sdAn/M7NGbrzMYrgBp4EwXvCvc+H
2cEu1fb4cT1rlNI0PNtuHuS9IFu8CUWRiQXlbkJIQCgvsK2X/5PK/yWfRgbeGQny5aqti3K3l2ia
bfas3C9gEJAMaGfarU3gW2H66wauX0+ypvuWYqTxqDInhi9p5R0zGULCQw+VajZBH6j4NetdPZFG
ur1kaD63J1kWPOkvuTjwmM6KwY0jfkxx6jFH0kiSIKoVl7JCBKk6QqQ323ncTXVVRexjdm1VtaKp
vxl1Yv8VrLBffsTuw81LzmNDRk/T+fTEmqhfxiOdEwx+1NhCSQtrDATOXthnFliEpFTLiAOoqB7U
fK/yUTohm0NElN+8H6Q6gzPSdSt3jBIbFS6tFfhJdIDYx+Ph3irk2lO8egQQHWgPAACl1sMytHMW
nJsT+et3ocXBbcMJy7p9d1QReF7lfNbfEUJw/xMmDjh+xyEWtIvivwDTAwtewcBWu2FCwPt4vPyi
mRxaYV9gNJDHl4r53cChuv2LGYjPTCJbS0OWMKyV2yatnYUxf/DIjCAB8BaHAeMUHutZQ+2yq/sT
Yv2Z391HNP01TuS9D5pq1ZA4TiCqXtsofaZv+7wZqNZFYzNPJcCwEGVff81AglxzYG7pzObJKHNe
prVZaCRncTdVAAqCzaPRJUZHtjkXkQi+ndeE731rVUp2fnuidlxdhyRFXzzta3Kw7d2t5w/hTIZM
jZjqbjwRwfG+dJtaLYB75JR5UsVZxOxU4u2PfwCYYu6LOWbqBPm/HEgI3JX6LjIPLuzx+hTT7rAm
n/iRLvsGgB2ualn0N06MaqMDFiCimaG+Mh62faIjNBdj+8G/9VcGthiXYrteiV5v/qdD/eq0GJtg
Qap9aEmlkkOHcfTM2hCjqALsnJEVQRH94g6/2spiN6HoVEZPXbxmmZKA8NRuG8ws8JuW+I2DahCa
l+pP4MKg37jht6hh9Udp4bqj+nEMngL5+pQOLa6pE+F1ZHfOi102SE3vE8obu8JwpH1g+mbCtWVe
41MtnZXhEaTR16oLJcAzw0/EQ9xzYefkapT7/lK3nV3eZS2dj16EVbWW6sWhgU/TZ3kkcQfEIbID
WoZyaFEf3OjStFtaZP0VNNuVBTk884B9D8w26GF2iSEOhkpJdwHZ3Ey2Vg0c0GTM/jE6Rg2PnwUM
eyfP+YqXXxzJBaVWbWGjK4uZG3qKxQSkZf1mS9x3c/QzuTtZmDs2cmF2qpM6g6ys+98FJKFAU5zw
uU7fil2V4nVr7ix+D8GCNMAZFW1Bhon4PT7YGuZ3Q3IkbrNJdCiwK0oXulUiIQ9YaK8einWl0XDC
ICveT9IL50p50Qf8jSLcSml3MpTtxE5IzUUvvw3TqPzCqqVq3uZ7ZiC4a3o9auG62FzduvInYdlw
pB+f0lD8nHTFJAZMVQ73Ip1Ek/M45Lot+bvlnaJAp+XQ6SFUPf4VR9hOUoA9uPP4jgohO0VfuFdk
OGWzYoNw45XzvXZhisQBtlJ0HPope57k7sBavBTlqUCPeaoZY12TRlo9PklGB5/ANXW7il1PE/Q/
zAre72RplDZmkcgFqVP3xORe1qMngDauFHNzwSGzkIQ+bmJnfDH7IwRRw/gQ3RACtAJp1k/sJPz6
Z3d2Dh9pG/eOve7icMnA5nklc+8iKrTob9Khq8KLztONhNg/UfLUMTRALnZDd8DqxW1qQC7D22uw
F8EUU6n7i9BKswMpIrajoU6EyOrIq/NXmvmzwOHUv4aU3Nm9uyeBOpeTqD6x0b+E5qmL/MYQbThk
zevDTd0EyCmrxOT6ZF9XWCyVbVzD8woxn8bhK3JHk1ykgOPPcib5+HnUsRQI7fstjzK18j/zVkKA
8XxuUOke6ANvDLIQffbCmXZhm4saqe3Vgq3KcqPcRgpHq6QWqmc78Eiu9qbCL147Ui/kJupseK0f
8wgE4n5Qyy5u6npJfzEomhBUnxOKMuuqEDRIMnvuUgP0iIV0a9Zd/RRssez/ZFV/kgib2Oo8XwM8
FeZr7dU5tNDsNUHFNBYgqmfjqNzNJMnL1vRl3b1yfUNWsTLxmC/B+lf6+4/uZFJaahCOLdz+oJSq
SwhV08X9XHkEYjsGbJ/xJgH8Fv0ZIMu9iNlyf0bpamFgXWWrCuljNK8/7oKxuhtm3yAiVYunAauR
A5ZK4ZLp5Zwzk0avHxLAawk6LpKedP6PRYuDJqgEUkhEQnFZAbNieTkSoTnLyojNM/2mEaCH9YLD
C+LfFf5qxvbi7q4uk4LZ17aJbxetW9Oweu2fCqQ72GcrS61JkyTqoZP/Sne6V8H+w3Fhh/uqxr3U
AQINKxbuKjK5KUQpIxWi6RXGZer1+t+WcFT11PrqrjGtdocFQaQe1kZLXLv8VhNWjW91cOOXRCHV
Yh0DKbqXQu0O3WJnTYUQBGQj8lp0tgtKkpQWagFD680GGqFJztgZf0+j+xN5ULL8R64Hy/KFtcxY
ULknzVNIRLFgmUqA5rAwKoxM/XGiagagXKyCOES+Z8ogYx2u50yaYiOEahPq/iGx2mbdDdqocJgK
Je+viYy8T9NT6B+DeodJktApxRHXdvVU/kQWozyO9d84PmmRhvSA426Zgqxntsd0ouX8a84ljFGB
+WzlVPADQn9YdSmloqEiDiqkdip3i24jij37z5TNxn/E3LLoGDS2H9DnWjQGa/EX1/TCoUVK8sj8
UuE+miXQeLc56Oz0xs9F8YOzno7CaE0lqAJou/RjHchnKQc23OGL0bvMX61BSTntq/naRAHhh+Gq
u+wbq7zdTAFvoy0y8O6C7CwDsVRSXRv3ns+WSp4D983KJF86etBrgI3WNDGspMPEaxQO/NqoEdfq
KMmqoomSzHKrh8YXqBEghW+Jg9w3PfldjaFGuvAwNSwFdReEztfVU3P5VJyJOBwb6njt7oWZYvxN
r7mL6c7ExtIB8bJblGvM4E5QYHF7igyVK+X3nCP2WeFpTeLSjOHhBRZ3jy1AHLb+gHXN/bv/qBgx
YbAKNiYGrivRvWvNrKAj9qhnBcjpN8w0DQ1NodiIP2+tyCHjYb3Blyagaraj6kKIX8WF0bFzRAlr
4+qLxEDmLfvUhPeOVSxcjAI3RurKTV5oRc801i2P5zZ0X9zUVkBBYPmo8V/BkyKKl2RbteQVTR4v
aTN7hXLOKoJk1uMXjdJY4fB53baQg7geM8VYsgonY1gEX7bW8o61o87CnQ4LRoe3HjCA1bcBKB9P
1bq4n3I9GgD4eNiomSe9XaD59f5/s46ArM7Bcq807D3we7cdrgjKlOpR0QqyQKc/uACEntn125+t
G2k1rEX8/ktpxgO/hwJqJMniaO4S9E4UQORZggS/PBoFrp0qM2AMrxpD61+JknKNXXY/ZRBSIipV
SBNOxRjy3fdmXxnfZyFLO7SLt2Ly3gg3sdaoqpZorEu2xAX1vOjX1PQKgRzZwSxF8aDQa8xTLV/z
MYRke78eIJMlvXB/4d9z5Uw9ttITwSK8Fw9Zwb60ulL+8S2XUqgB7emOOJfF7K591w9x0sGr3d/w
LfX8/A+/WaPMMzwnj97HZJCdN1dT6QhYlRxSbdxfCjqdv0io91ihoPtYcZDEy9HklYuLcil6fIdG
6RDsT+Cz4U1NoUJBwkrVOBsz+FOIc3RizidIadUuFc9Le98VIyuSdnhIsDBUM+E0EORe4rl0ZpBy
XXOb8q+U0lCuL7BjHI+OVlu7gzfGecoRKxT4WGYnWLlGj7c7IIo4Z1n7xc4BPkNcYh0UGE99K+0n
VC9nLOwTVQEvBp072wyrejaJf0lBBsJWXgBMCxfjU/8gXglcVuWVz39MLMclNWXTT5UHs/PFJpW1
MOkNDTDypNCb3zrLUrXKfBAfSQgdKatCdNSIJQ2lfOKpIKnJBgen+DFKskEqEJE9y2h/aQ1cUUYU
c3EYkP3QLYE7oIGAHLu8DIcA9aP5HPEr64wrq0nBR3UVxSI/CYacGSI0zuk5UYsWYLk0BlhbyjY+
DTlD4BQaIHED8uodL54aTo0Fs/hXeLWDbbyZ33Zw5IICrZ9RhPPFcHxmNYyPmTTW7l4KX0hAvWkJ
Wle7PUYxCWtoxsRpemTLOCG3RDNNxSwEqpNYLaGQmn/BQss9GzD2ShmFuGojZnoown+FOBTvh5E3
7yPm66pfXHlzEJ6h3oYYzxxm9dxK3fChgJ4BcSuyG10Kaz/WWwEcAc2t0TIqFFdFjZjqBmZ6MN3r
GvnMGAs+6iWAPUPl7QxNey0JxdeKxf87QdQ5Nhm8dTl3tuPRzcAA9XD9XHToWNu61UIrtiXEjYBR
7+36oxhGoj/c3RCOwXbt1ze5+TxBlNWiN7OR7yawxwow+hbnY1uBoDF1Ro/hJe916jcQhkfzTRJA
VfDayOLGqA7oaNAy7J8Yo1Z/0SYs24unbWNZmshCSwSPPWfIcYbIBkzGJb7Cx+Nd9IAur9pWMTVF
8d9vXq5XwS3DpwNVxg5MM82UyHNE2hxSDp/xIAWJU+G9R80cdeYV08ixqUIeKiSVM1t+6Tzpyt1x
WlxKl6SAcYyELIdXh1Zy0ENEkYVvLhsIUE2R9ecofKoti83d/6kiFhnfH5DLpfotMiqXBbG0gpPs
Z9iFg9HCPTXmLqg4/QqV/lWiUXnmLqGEjMzy8J/xv/IVM+UauayYlvafnaQXDtG7LbirNS9wOXXu
ZlU1IROgWDJMoK2GFhdtGMYR9IgfDOIqbQqFW/hmqtVe+wYGtZcMq84AbEJofvcl1VH/4cFA7N+v
FAbPMXgtb5N7QEjVzO8segB6A0sLdzxh3QnBodS6k/V1MUl0kWRjGv36zil3aRO8jUeMR0SA1aH3
UTMGJUDhwog9FCO0OtNJ4a0B9xPU4hxKvbi7wAgOJFaBloeQF8IUh54VJvlA7Og80VJaYylx0jim
oastQw9QAAn5Ixq1rOwibE+Nn50c3eV0m5xj3Zi/bClUzXlfwItyMtpFoTB/vcB14C55Omz8ZDwJ
S6a+ZHQDenOVxCWZCCQgDX5WOjkBboukqVv4dsE1NpPvZbeEXWIgGFlrhCXaesjZGRz9I8VoP+GS
ZKEvp38IyaiV9k6l7pMdOvRQXJsCh7TvPxfvpI5HOr0H6KQ/4x1bwpoQpyc2+yuO9VHDh4w9GmPV
M08cardLJDaXyDAdbmLvsdXwlzSiM7SnjMVGENErLtKjzNnE+1FmuDfbfmjjkwCpTohgAdndiZ49
ocbNh3feERwUg7luG768XOoTwl147+W4ob4KaTNkaY0cMMlV4INDzmZJb/9UFFPUdi7iWJXayzTE
sLn5pjoHw3Zt92t+5s6oDjx/g4M5CCoFMGaTobHNTBMDuITRPCQFGWQraQCT09STJWM8xM99BQZu
/gY9XHePf3/2kINn94lJ/QlyGXK3Tn/xCBCjpsV9UWZVjYXEhnla2EQRUOKFdQxEnfDMrfKZa6Yf
AVGuo8EJ67Bp/koSlY3+PzizSj5n6WEQoz0LTzHx1aXK1PHadQTMFtNmMvTBEeCQtUSLLNg2scnl
ToiUOMtfFqDtxb0nuYRiExnuUJrx4urEP8ImtAV8TpNiYJhXj9P/NUBktnCXL5NH7xfhkdx7rtBy
hQ2BFvComXqUHcbX2w9L1hEZGphzmsEBs30nVLDxTfL0LJt1nIvsIT2HROFgr51GB7rBbozgikTP
94l+vgAPJGkpAoGMOmLlKSKVv8ALe/rsUmK8BSy2kheEFQGUmOBWny11BJ9m4Gh+whuM4tUwHwLo
WPo0DIjDgwDMTfzE3i3/9DppJbMMMewMA/aqYySIuecFJ13SDmEFYrNN+VWPMCpQfqZa+EVQ6eiD
U1WowJXh4W9JytayZa1sEops32F0tYUby2Rvko6eY/3vJ7iKiG47uVguBHiM0wJ7jIRC8kroqmRP
LyfBOiNFwXBhofr2VgwpGzlOINZefJguHfuz+Wi5Y0z5+N0gsbUFvm+SSIbAHf+Yo+YSq7uhmwHh
fHddC4KiKsmBDuXV5gqd7+T/oL3n8C0+4VTkgAbGDcVcNWG0CicrNVnK+7osV2+5Qp8tLNK7tRZT
ogymmHSDhcK8MfguQaTht3fxBZGYYWuZsTQsvjmCrbxKDiPb1iZ4Jgc8zNCDI7E0/WWJU5OWgt0k
u90n7zMT5/E4uSy0303LETfe2PqgCqFEQWFF0bW+BFg+Lrz/cofB+2NWeL6CfnSTg4WDumzAR0Rc
3vNBwgqERulp0YuxlSWWq4jFbdcAicTAR1EKGzQi9JinD83iTI/Pu7YqZi/r1bHoRt+oXo1wzYKl
hEqQtqqVX3FQkOWCNVRaY+fZM2+Nqc0DfO12Bl+ZdS5cT85mirdqQ+dS3/e8k6jK3b9CF0ATc/FK
0q3JeKfav3ByZNu8MAPHSdIj3uhM/Z5MsPgd+Jz7np5+mfOhY83s/hx3LOy9h9pYSMf+/KmjcJe0
ifRaNILIHpSWXfjPF4A85sSWEmbGDyWUOp3FIrS+T4j9Xd+GX5bWwJ4UX1mLQRUM4WtUYeb5JJZE
LwIrvhpM93EDMb5wOIqIHWv8Orh4D86xJl4FDLqJzt4k+M7g0gJoV4AYRktiyVj3R4HCqnhjC2yW
ozjdSL05bWqWTPnrX43ebi272yehJ3uhxaLwAnm68t3TLFqlzJmApFmYUnil8WxhhFo5+3VxSMVY
76sXnfQHt3wA2cREIDFrAHgfSRCMlu4rZgYs5PxFmXx3MADN6GVydeI20dnTES18nFDFEf868Eff
q2g6/Vk1utkZDVWrdny5SjsMf+DotSSUceWuMU2QsRItiNSJgftwIpW3S94yzkKv2EvOP6Ax6rbf
1U8tiQi5C4p/NXBEYnKJ+lUtGEbikjcBOEbgu1fPdVb4JsxWOpetogk1ETS7UcLj8J5UMC5QrlT0
Isz3kUtPA7MN0PzyWqDbTAOdNoufxv27BpibqZlOGy6PzK3E0w5jxRzXWOGHFrq+YIBPJkm4ER0N
cWUeIKsdGL9nMUtTZoXw12aCaMnMkty+Ifkn4Z06N6isZHrXOtS0y/vO8trrPHvlspHNPFE3/OoC
qSgp+wb9rrOn3/wzHIJ1QxZusJoVsmTMO+n806TVCQshKvUxEyzM1x1vu+ZPg0sn2awqLeKIQ5tA
9iwuAOliaacWnV75DlxTrjFSRYuQFS8e8jdDmiKHajHA3Vygfh6g9kFfBw/9bpGpwDJtNHm8+VyA
S17Cm0mUNJ8wRXbw9lE+x9CHQKfrd8MHUbN12lrLyBaqeQxaR8gyzwkg30PAjP0Aj2YPtBZ0ajH6
hZ622LY8DN7nc+oV345j9X7IJ8yAt/5D/ZRkBLcuSwNHQSk60t5UnJKHYLzeb5WJ6hxCK7+AGdbs
JOSrl1IcjhGKUT5jCu/mn3g/nX37FKcxmZJmuBBC+zCXFHZI41Ldje9ZzrmRyFQogXXile/J1iXG
tLH/R66xFXMRSXiFg7W7NETzwnrQFgxHWdImYd6CWYsRXeE6BzY2L6aH7LCL7oR2cNwC4dUaWYGY
o6DMQ3DcI9ArTCv7cl9f+smHAnlK3DmE8wVWVHi6f2o7u3lHs3zpknTwDs7DM9aoVZdpGBeXwYQD
5Oy7yHsnqblxvd1F1FlEdcU4miCL1Km7MnIYMPNYyorGTaRRiISCCAp/T0jze/SF6ijyYEYmXHws
rkeCWKpNKyOHJf0vCKJUh3t3/Jd4IyFEaG+VzupNNZAEeCf+9tHeAU4hvdFugMNC7uxi+PT2e9AB
bGncZ8WPE0xk+9f12h9+X34qwjI138Y5jQqpw45JmG8Sfsl9rF2ov7jm8XIUqfwo3oZtkgCl4wF3
F9a27KUikkD4jE/A0uv2x+ar3WYGbWN4Zwn5WogioZHmJPdC4UX7ARbfdJX7pRiRV+n/7keyDuUT
zL31f4rrUWe7tpc/0rg5Gn/7y+xzPG9SJcMPMivERamVL5lwEzD047q6h0SefPCWySc9aL2aHUWW
t5/lE76yzk193hKGsfM2mDPhJWE5DmCCuYoUtm4VSFfYzopg85GwFZpB7hzTAkjfBKh5t9VUb6OX
IttPmDYd6W3CbfoH9Xhfh5JvOwJvyCUP+5jIXys0Fo5NQ3XuWPlMU8OhAOcFoCjnfTbjMMAIKLtd
ZN/UenF1FI39OWreTbS/z8TGb4KzJaPsYyF9Zwqh55oMlXmQheT7P9vUxodbcxx/Xxah09jcGq/v
kiWicOyjNd2+fKkj7M/uKPDiNrVP5b1gAXhGByWt8uSllKuIQpvX6HXt/jD3d6evw993Kl6zQ8Db
m/6SB3GRlek/1FV3EXoLN9DCI131WSJvE8t6T7/+NRv0E4C6bz1AMGwTMqGs361oMDzkF9RsnzjQ
eQNa/M5F+9YrW78sxEEEF/0ZjIjW1Pu4uB400mmg/G7vYOIsFL1aAFyB0w7N2+g9rs5BLn4uOqCX
xSZKYo1bwlkTk6rOpM5Kks7nMgP2EX8ZClaHNQlj7J4gxji5ZjJmBI7yo8peJq6QrkyZJP8wYcb8
4noEEfdiCKRakyFeXvAz8J+f+rwQA4f/PuSRyqj4s6IvyAR/3QRqqEr/lBmYpTJocucl939OCS5x
B/54pIRW4g+oyZ0UmaCVBdbTPmCfPu/hMnSzUkOYqPojKG/zEvkUHThn+x3tKNk3UCVkV34j7C1n
VUTJwnT/XShY3NYEhpM68pcOTGief6rQnplZ3YA5LujwF7xMevxRu1TIXqrAFR4Dq2gotbyt1qeH
MysTRXY/84Cs0td3ALblnIF7akCbimmuIXNgh3xb9tLXf97HqJyKMvr7FmJS7ZQnLmIfhS3sK7qh
CpHlG90atD1HsTbm6LWz4NoHOUuqJbbZxn9Ez+XJ6jkDHwDKQrTcQnatNU6YvuuOb8Cck8QTd3os
Xtm4YYc3yQOLxsQ3kCffvvUUuKnTh1ohwek0UcIMAP7ILeFZnuVHZtPK6WJOsN2/jwL+iZqAYCr8
6P48s2NP65OLT/p/HLmsMPqoxFvV/BdZehC16koHv9hzKQgXm+E2cNF3T9Ka8IgQoloszXCClLOG
8mxLYzXWH4D9m1ZGKuODgd3WMjqCyMnGofTktIqdqRPcc7QEL7xbm3zunh3M0p9u/qr4qUffOXOo
J/xZ9/lH4Eehnpd24w2WKjX0HXTLMtjhlvNsW3a9JxUtb9OX6bdXDNY9NnPd9eSd+BD9NVdx/TDs
yvmN0yLK2Sf2GrmMiR7r3WmNb88jLJNAJc3GTyOBJHRekjzAAg69+2nvNA9G8h4Q3zkz/i/yHj9U
e7BBrskceG+COgMFbfjiVoSSgBRK21qkC3CVudxwTFu0KBblf+JfIYYEDdVhV5EG8hTola8Asm3d
vsMr7JFMB6a48DNNPJ/3dTDkp5PP3dnReZAp93u3dy24qxtz6Lal+jletdlOJ4HSgWj4zZBKE9j6
QkYz0kLYKnZXn0jRdsJ3omMq6zqZFk+9clVHBVjp4mUKYDNyZjClFY4j8BBlgMCJhLz3eg2aDEs4
1cuzhk4rYwuNFqoIU3zKzao4daMTjKWwZIfqBXPGljFwNnX+lYT8Lqranqyr90OV+oDQ3ddlVdyw
4umYM6vt5OFaP/5F2KRHYmJjjucGn5F5hU/liRUiouPII31sjZFIEis3zx5nB7cx3QT2i88QEWXO
AQOPrHDw495lsFJyaIehLM4VbPvKb7NJxMyKvuTunVcN6GfO31a554MyyWNXgaksX8o4jx2dzZrn
1tfCOpufn5UuQ2fd9jXfEWid2sjcf6kyJapGNbJ8ZzFyR15JkXPd6xZGgrcdP/J51Ov8+0GoNe0U
nO3DpIf1MPHWqBoQ0hx3fIVlpSyX3IeYWphpwty2zqeOu9Ba3w6/EmhMOLTauoWjUTW4u26KDcAE
n0OVvafIp12OQ+TbKVbFNpPk0HKO9blsIEzIE4wGhzxDPX30wrD8bRul/TfT5Bnqxjw/c3DizVNa
+R7g7UDYat9Jvf6paFIIbPngUGBSNhBjobQS5DMWivIKgSj+SXXQM9tODF1WExEeehoAI7Q/R5P4
EoVs+W6341+u3r+6LzMgafmrQWeAw1F1kjZ6/4GLyP1HeZn1n3iZmjeDaWogxKZgRAPKnW8skyiS
HQoEEH+Hrkjy+SOyy3YKlLrI/3SWQjA0x3EZ1s95D2I11d/27F44K2cJ2gkM0/lSrCHbbB6eGPgO
zZ5+UVQJ8+gCsKCgpHSeYHFkh58jW9kbsrh0IDSDZ3yvMsRXZJ7ML7cb/oC/phdmz2vZtovBmgjA
oteZG/IdD19GCLbx2tbVNfxkjjZWRQEADH1fOKHgqdsHcAlJIKQjLz8sNGNFYkg3da1gggWYDtVz
KHklPzaSh3r/bqGzbNfdNVDIiPgf6KexXEc6I+1WNpAe4es7uEBN5/g/V/mEwlUM6aceG9Xr39MQ
EKsnwrRyHcwxg0bmheOlNg2LOjDD3Hiz8dYoBxxZnuA7FNrRA3HLBhlozz63JOoEyoOyl06kYkOQ
x8qeA5ASpzlAs339jjyLJWN9dMf11T/wPJ0X8bTPmKSO+wO13grAg1e4aII/hG43sPLuptHRoOQ9
PwrvQUlzcxWu7vZv8CgHC0hlKuhSLny/hHi05IMFU6V+MRvRn9J8uvYNq90X8bsmDLq0Qm/GMl4H
nhksj7ji6q9W6VIFHSk+pUjNcEXukhrmxeA1iuaUCgC3IPCowFcATTP/wLjT+ck42N0SfDJs8qzW
sVTRMlUyTlDi79oU5XFiPbF7G6ekhc+L4iK1Hsxqhy3ojR9LAv9BPDQu9h9F1O/pH35RC7dwlbh3
zplFVAraZEVvFdZ9TTkmrydiTwbiaC7iII8zDnmRM8VEQZRSNGQ+WGf6SLYM2obSOI+MD/br0y+Y
1Du6bES1Hf3gST4fiRoJ+qljYMXBG91Db8KOnlAsWfuAg/hVTiRXLSr+Wou38dObDGnSaysHoEPc
OBTKG0rXKQ2PnS+luZLeFpBivyPUGqcVSQ30GrMVPrMqW3/5/Y+vOnhr6T5V9eJWpVKq3mqVUHr7
UrCWktcjROWCqMJikZkLEOc/+xaLXApqQLMnrDD/91Q9i1ErzMOjNzlZbcUNlPPgLg+FZA3AGkDO
bHEN9pVPFMjCK4djxOC3yWzAHf1pfCSgGGN4t4VZVg1AapohBLJjTPFkvw7511pRnrtJrYqzMfX2
LW+/EjGKNHjKof0uwxsVbEU1eQpUG0tQdhYy9Msg09zctSBwqzdNbJAbFnR04MBcQRvbwu36Z3SM
5qNVZE4R+9ZHC4PqLSol4t/3Xv+87R63W9NtV/czwoeKMdk1NLwJOgFKoAW5+A/YBezqJYNWYzpA
w6qVnwhYF7C3JvUmzravhJZ5sHRr1jS1m33h5w2GCovTzvyS2bKndeA3u1RdG+6YB1j3jVFHRsjP
6Jirqmc9f0rjL38CVHVkSV4O95+zc8ZSnjXr4/WIKselTgiFlGmXiW/fH0qsyNHdABgZ5eZCGbXe
BBwvMoShKYj3lXzNliVgpJVaMhbwYB3wHNmx6XRI3Qfb881FiHx1L+G8swf2r3Wt/VQZzQcv5mdS
vPfdZQQCUKDGWrD1HiX9JxeDcw6ReeK3AxWhuXEHIpLzAvqnd+hsQ9Rh9Tro11TKkZu7BAdOJbRM
CfANfOvZz5AXs3UYF6AUHq812rMyPnohqTCVMFmnTIm2yhUFU0pFvl3IzUuHhY59NFQ4Kk7cdzzp
sG5b/SaUhmFyk0TTCrGD6UspQHISg6Y6aolnD+2caFyrEt/CY+4sE1fiWXS5ZQOfbLdyco4vhs3f
IM9RYLjfHHfHBaZQcMYO9iHydcwGUGrAMumYs31N9pdmD6zcKSK3pENhSle0Wr3i5C+JO9t+7uEk
Zo96bGfgx4OMV/Qq+uQTuQ/iP5Cj80EOIFDXEeZ5MbibONLVW5yTuqok/3o91unf7PONO3KYQJl4
0zxYlt81BaUlssjnCDYbP7F8pwJmMrDwzDgsM5e3Wf8eXgrkH2uxueQyWWd+DIKW0VxgRE2haDfr
sS8Y43ZffZ4MdIHGiA/Q8Er5cTGe0b+v28wQMFTP/FMFHgmc6q1mXQfUL6AeLlpAj7QpXcvqPpZA
DHWnjLWQoTE2eOVqMxcCVFgueDgR9uQEj4funL7+7qdQlW8vfe0Mq1OYnETCOD9iLaAcxWEDnYNg
Xk9TGWxd3qqtZRuHHwAGRb1k1Vgv+nz0PIPKduPhuIzCxuIdm4GejPDuIEU7ZYPOHm4D9x9a/Dbp
TNzV95KaRPqKzFzZPapg6/qbMg/Hn+foq1TiurO6fq3vHpsW/Wl8+AwGAf+v3lrxxED5ds9HJ+/f
GFFRVooI5vOoygua1EpcGnEW8QUlF5JWfEJOJ0hBLoFtqXZa+7ROVfsMQ7Tea4yrM27COE99g4UA
JpJPijxacNTPFJEBqsZLQS6gO4i4ofmB26bnPtLPvN32PTr1B1z6fjGMjzg/0TLtA6t+Ot0uf1nD
tTPKkkf55FbVmEKpQLQHpeiWBIjbhKGAJNGHhA/lWdJyMPCaxTShOhwODYt90dZ0RjBaYkibVknp
dCRBTJEf0WNL6ARV72FH+X9D5GuO7D49QFkg1F04Nc/h+0uz259LYwNweOJj95pHTxw60Cad9pad
iOvjGWbbyiVxolximVUNqnAEmFBPlsLVFWNQf7SKyAstBcIDR+h+Akqh3S/4GE8dFQXjvgKndvCE
Ki0814//qrSbuG1HEyTjhxEIJjTsBlHKfsPdR+qGXgkqfPdLOXYRlyjOMbIqmEqRvP2g3kq5wxRq
V0Iy5hwj0xiufUzV9t+TJdXD0w7dEaBQxDJfBISAraXTjHrqIn8tYwCQaS4j1Qf8jLeaKCjhnJhN
u7V9CDiQ/XAPHKbRZeBiOsbH5WlvOa8yrLqN7e2OW0MUYd9e6qe/UyiHV9DY48P3WdcjD8Z9bKVB
n405Eu4Xgi1BeTHTsFCXqrRqMPwaq7wqKd+Cx4MdhTt7wfJdIF7ybf9+i3evHzlKjV2Yadj+DGnK
eIAVjQZVVb+cHyUiF16WBKtch2RF3aL3W7iYC7URrbgtudmD15xpSfVPw5fIKsAg9+18HFSvir81
2nWNlyJdPk+WO2TvXBFvOFX7FHZnOGz08bZTWTwVD0a5AE4qfxQHsMi6zvUeakxKAA0CJ/H7zA08
KDsNP/roODwUR7Mro9oCcF9zGW7AQBaqzqqlG9b0dMJOsAx4zkDRHX+dIQAjFQxM+LVuPKQYY+u1
zFJlPFcc26kp33e69cjCgqwwB0PnifSPaO1SEaCKvHgX4TgzbxZPLobwUWvWd0fgIkwaoMdT+Bug
FPtuHS1tgtsxorlSbTgt+axLQbycUtL7rh6F/OH9Bgz2+0sYGFSDntqcpqNIm1c3FChRugxNJMdE
4IueIwAtAexVwKbVx0tf+5gZkRnvJVYxjqO0iiRH5vRANrbnWaBkdj+5JDew/9pS7bQ2oV+4bgRT
KPpxzJKbhaAeCWtIiayIW4STko556usMTdpAc5A15YfacRUNwZ9l0UrgKxYhUNDhIxw2sX8VKhcW
gFrRPQxOncZOrYRIIvT3XAyka2r5QufCsa9Yi8Kf7Qu4re6TVR3WmzNWOiz8rUjtzxgj45Rw7Zz4
JLlKjs5yg1Zb0EuHGenSyA0fdWvPF3todFTLIuEV1/LcNm+uiDhgcKyRRYtqmlLkpZtOcdvk9BrC
y/W4sLRdCjs8Qw9Dy3ZEyZ08ptiXyDLj5rpj53HuET76n5JdsyyiXSUF30XbyMzO8vPuJqGJ3sXv
JJ4folldK0XS154tM9djI9oi2pvGPT4p3wEHugdy8EHth7ef63gaZU/MkGvej7ar2DYEL3siPoOp
lzqNMn5hTJLWyDnrwIgo1vJ5G0JiLtoSrCeApEYEW7TaCroe8X1fVkwpUhRF/Wgc+NtNvhsbEB/f
GT2KkL9LfRJDvxBC/KJ69mNiWf7yz3dYRcyksadlCNLD5+J9Ixrn0gu2B1oJdc6Rc1rDcwrUDL6u
D/WhTIyRIua/RTUXWIgQ4tDjI1zquX4ris7SSIaue1HVEkVi4+lt9KUMIzuHD/K3JNBpUEEEJUt0
UP3KBlY6TUPidWkMCCk5QK7Z8lXClJMkGqQr8PtYhiq5giMyGc5NCv0YaPLE5Z9bv1XzDHWVAZ8f
QlMt7zr0T/c70eVjRUq5Ai/5oFZrCyheS4DD4ZjxT7kLilUattMFJ37RhbpwLG8wHZwkllkhzBkR
p9d6PMclVsJQ305JbH3Z7kX+gmug8Det5X90AYV6KQw7ZW8nFWeayBw0clchZWzWC346YM0qC1jH
fDXW46/0llCAyE2feLZ7Tf+S40cO8+6Q0SlcFVFFJrq57LKzC2/ia92NKrQQ8DBaHCjMDMWhQVFM
BD9eHfTT30ON6SZSxOFsSWORlDHRGF3RhShZzBgdwPwCws/aD7ThMTZDxUZNl9jc2PC9dIbthUQk
V3FGRNbOFn7zPj2WWiuJcYeo0mIvvlsyOHcnhUqhFdy4k8LtkW8A58akg6Tcui0rE3qCEBlLxfRA
aipyjMZC/Hr7I14Zzz6/11ZUtjMeGYmKxcum6AyNykIYQwEh5Qq6IExN3+X0158y2FPLVQvDSqMq
5KMLwlD2ewlPqYhIeHV2Ll3A1aMhwmL1Bu5uAU3CuCgF30YPnMVusGJQW1X1Co18BDWvyhRBVjSM
zaBG68RfCXQQDQF53A6KTtv/ypTDKrPGED5ftGTINUbEjX522XfPK//N6LsSFBbTu/uUaCz8rz7J
epZ71ePkqAOxVO3NE4pd4jjLBu8QL9doQtLcp8XaPzZdoQ9OORKHZmOdx3c9IB34DYNH1djqgjfD
8cKpioi9DzwHZyzZN+rVmeC3OhtZZu8HfRWI+XlbUwPEgkAv5UuIjewbW7iTgxeN8Aipp/A6ADkX
dB7EUoYpzqxm1/pSQisFw0iVLbWCNzowuDmlNcs6p83CY7jK/mfMEBN0vw86xY0ohGp3kLc147+E
63SlQUPCpW/p3RSHDjACPt7vuAL4btnM5xSIuAWEvOREznoUft0oQmAbXNzLU4k6yUfdLVt3dt3Q
9VmnoFm2yisVB7EEz8R+bxI8MNyRLpIXqd2iok5GqByHHOEbrHem/jGJyzisQzRJqZM1rjI2Aulb
MLwoDfM18hFbSlzcE0iDZF30fRoN8rMp6LBwJxghvFVURhwKNDxGmx2hUyyn6VTZwyYBCo7nf/My
Qmc/dk7z9ca2RLlnWw0pvYzmVmwLtkzhPEXwrmghNL4Pod+YB5ky21Qdab/CZf9sEyczfHeBx9NI
uT1CSpBkUqsZ+7+lGmxUDJ9nKBvfmbbv4mY4LadmQ5LRf3BqXRrr6QKHGQX+oMYsu+YXf1gJFkqZ
9kRe0ue46yCVhTvnwPGp8e9Flziv5jCB0GBTc92HyW+SvQhUKayAMJvFCvbIZYoiZWy8a5/U9ypw
kt50gRC+yJJxuWf/ysD/kzBHwVn/T3VRD8/sorA4xTZ6X5UJy5PnDjVzaQ4/uzBlttV17h2HJlDY
09o9NdIy2NbKoqfHXaO6vOO2Dl6DEB9WCnxzzL2r1v4zdpF8O3gjOslQYjC54/d7OHlFmKClU6ua
xlJrwQbxrTR/j1O50nV+rol6HET9ydJY2Z/1AvExw1QXoZM7B+vJ0u+gS82APGtU7vthpjtcCS00
WpmpEqbh+0SPTlqHU4vOcuoTRdrr0rp9Ywr1l9VactIkLMRQiCl8sj2tDwkzBq4H7AvhICkSyaEr
PnyeapAtsC5CtjiZjIGqoVelwKQ2+N97OWfFNls/4FIPkKxgsN+pISTTeDCtSkcbgkAyOoLSASb8
cU3XIidyn67uBUSznrQAAzPAtxIk5LuR4LwHyBCULntibgzFN6UTlJvMHRmKZg+Xy3OKTgaT4UEq
kX5C2uxxEmrYVqbQuKiTYdSxFujpjpZATpJ+v0ehQbRbhSBHH0vkvB7f0MdXGvCVnEeJB5halx8k
PcDRfQ2aCDlSN2l86ytR71Equcxc4T88Ym+RpAbZRUaG+Nf4e+j7vYy8IKJ8TpclJuCJP9R9bgsw
g7SMlMVOgPR1WuyduBqXFlwPpDxocv9v/zc0nC8U39aTH1l/zbyHL3+qlHRt7VRQ+Q7W3kTHQmx9
RjdOGhBVQxzFRL4knaV1VUWOBi+2bmSqHu+tVA06/RLCJhb7Xl9KMqcAghiSGKkLp8hfEcJQQGC0
glf79W081K2CZbFtiEnbjbmyArF2rPJU1Nd2sjFW/Rvy07MH1in98fWyyZS+gfYihNYqT1ymcTmg
Fr7D1Ud7+ldjqx20cOLVtUkydm4J+01mxw6zmDqAVGJBVP6aV7T9qkdw/U9DeCxwLXmG4Q/+Cy2F
cfsTsUy6Nc8u1Skl5cVl1ZzpI9ln++/8JLNf+VanR42fREFOQTDvfC3nU7WSoEZfhB5mspONUUXt
eiYoOwQo9Mj7b2XygfyyoygXvkmRfJbJimZrOP5x4XaxV0m6zZU2wBdwzr6DbcPIMxef4UflchFC
Ex/0CYsmGkHnvbzoP4RHvFxZUjNMdP9Ni1nuL8pXKdBq7914nN151D6S+nt5PSqDh1S83eNoo8bu
Xh+/AZhs0RcW34yBXm5GgGsTx5SZuj6IKd9ZEF6CMCTTQ6crkOs79aVnBRcugl/0Ju1m47vPRba9
VEGcBRwq2tLcjWghcgVx41zkMboBFYYisLTtNEX8nYAahokkVZAnLoJAF9TUQhM9j8/djILJhxd1
QzGtG51CyLV78KWIpKr9JPItNBZqjmoJjUht5j0bm81FLpulj+6f5Plp3yqHOfZeM+t209VfLFg+
KvLywO2KFbGLw3PVkiyrNzYV0hDh8Jo4Ymq76SMqIIFwXJG8+Uuu0td6C9qJ29ncLu+9WfN5D08Y
iJZgkOIt3Dw6i4h+cVwiA56fo1ozm6SA81HlEosaVK2TWPmk+C487SYZyW3fuoKI1ywec2FOH1Cn
4QyEOeq7bg4TvjoCGllVf7bwW+90W+agSI8NXKXnJFYz4s+pwkBYP4zs4WjaAdEewUkZdZ5IfDPv
AYhVQCL7HjoNO6hoWlITcrzqV/NRhyfzB8F7JZabFMSqOAb2SUi9uU5iDjgLsISMnJpmnj8twk7b
p8FKfoekjby9+XRCZX3F9YAPk0m9unO9EKko68Lu9uB53FNRHyZlb7DP/Jvd367xZ9BUYW+Jm6Ky
yHexejGQxZHOshNrdJatHxVCqW/UeHxC4z+fhfh4d9J9eTh1N9GbP4PBbHQJVQvQnx5U9aDM7A5B
asCAzI+UJ0uqOfjXQGRONVytQ4ISGDI3jovk3MPN21h27d2Obzj3tE/XXeKW16+SiMTQKp7KumMR
VY3Yy8Z8nCoKDSHmyg4Jv36Fosn0E1Bo610e4Tzn0/RO9PGeq4WDRAzTURgD69fFj7G3xeSfrmhE
+b/pz4yT+vX1E33EAQdOoFrRvsSIOMavpNs1i+y6vyOgyFsn1joFxq5S1zTWvgYhB6+1nER0U4eE
tHO51pwwTskHaK3y2XHROUzDojsQW/0OB+fTlMsCLp+xQpWrFxLWeJQgN/Uvx5pYs2KTXaR+I5xM
XZEK79ukVCD4u6hFx/uKT/FIH2e5uQ8N75EPTaiTqlDMFAcKq82QdgGw19DltK1M3eLmbCkx+PdE
u8L5z5YSISEiMdgqP2tnzy/2akljrpkm2OLZFy1s9l0zukuBUvY3qAuLj3954R2xeeXH+CiGilSI
pJfyrQ8GJ6LUFj4WZ8Pb3d5wOh6I8A0zhxkYuvbyt6ZPwURzi+duFDgJyoBLnQNwwSnj33XF8O8O
tmhURamQxEPp9tkqk9wpWF7lWBVczIiu4PPmLgZq3CfxG4aMk2UA6lzYbjHUmiPIN7jLrNxf5qHu
bHmSDtXh+LKj1iDoOiPF6nu+j06WNibVvvLwiN4wWl+OMbGQ82lx+Mt3plpG/2cxk8GTqYRbEXEn
uczo9cgUkti457A2EzWIWeGG7JWTTKmFCW+tz02/S1ELQP1RgF8rfyfAaGjOjMz5ROmRKkVXJ1RY
dqY5os7wodh9O9XTWOC+nnO2oPwycjHJQkTt5f5sbHvTzGEvkB4TDeU3+fKjoUEftXoq9vQgZIYN
DE2rEb33ZhJktU8c0mL5VYRJUnJU4tBQ2gzsymN7Niga0/rLZiAVCJOjvYtEdXP60ewPTAVltB21
51c0w7E7U0ghj1O01WlgHCDh5uu9od8LtIQGCiPMYCjwrKp5CtW9Jdxwt/3LFsaol3VaS5QRlf6O
50rFO+3jCL+sBWWx8f1OunZGErY7c/yq9Lwp8WxdN3qEhnPgT2P9dWIowaD68HjdalKkR29yhN4N
sAHyUMhIvszuhmwNj7aZaVBcGBwKLcJWbS5L0Y9gxhDBlGs0B42v0KyMldRakdJiElLrEQVH9I42
TNE4Zg9T7f7QRW0sHAcOEpMrgG8w4hMBwFv2M81OdsqAfdTAXWYhZbAXtrdag2/apL/iWNlEmSrz
1jhUXIoH5TOvrpxN+RyC5jdJGyZvRhpysKSZC5E2wUnrBbjnyxesAZHCygLC8VAJ2+P6z2c2ZxC4
lry9NI1Ls5fVl7ZiOSx88VoIRgcjoOGV8xgSAm05aeDy6GZQ1CI6YZVmGAZroIoYel6QH7UO5Lz8
0CFLES9G7YFgYxZ8TXN2K4tobDFpayJCkroK1TE0HG3mMZgCK8lOyEWqORG/22Guqjo/3WbCb/5K
PX36kZ+yk0OCFuoxNQ+T2UD9CwvkTwnDKbmlFYvTnxY524x8xRkA2lHBaDOj1IboTrrBKBp5wAsk
3Inv9Vn0YkX+dkGjy0DBlSSBzPjICuCeafJe+p9z38uhsIP3wl7LWsEsTn+Zke/yoQOMe0VUBHhX
pu+Lg+I1YqmO5oXdOHuSmCnn3FFmABm08iqeMKBF3kV8WRnt3NKlQ7h1iAQW11KNNNPFvEJKHgKP
V06FsTVGetJjK+3jdwpkP7YXdU2ZE/FVvvHI/qJjvLm6wTO26uqczWDogY1F6DXTx1XQojsplchG
GRE97yP44NrNWQGHghIPTPkHRLIRndlTXC5MjKti0y3VMcd3By4gCYage+XOr2DpeIT3YgvMxU+9
TXvo29vwHS7BPOIBTVahZuuR/9+CSsVxUBR7cJBTmDaj63XxaqfFOyvycKFXL5EN7v2Fbtr2DBIe
gBm9314dyv30giO/H9ShA7o3qP5euQss78G4w4XWIaiLDkg0t2PELQRrffJaCxvlS8UE86iX3FIG
0nlQzXbWhh41GRU9BrMvvfdmT7t0VHH8ca1XeovK1aodpgHFtF2mfeIceF0nnD+vFn5Uz/IR4khH
dZoWQdiLs5RcEpbAexG0/ZCLonrRBWLTw7jKN4I6V7v6vwYG6u0Ax375YmB/7j8LXt0FluvZc6Oz
by9luk8Ra569ASHf2uh/8Gna9A90GhHVmmgI5p5euvbdkKQFAogK27UoJ6dtXhUz2fwysEhrRYPC
d+FmF/ilKWTLE4KCx6/gxHvoOiL/Gi0lHA8OJMzmgYh75cbx2FQxjiQPFcMrYbtftee/8RKZgLVC
AAilfZtI7YTgMXzujYqtJZHSfXjnZ0vH1EExKTQPaeFMzgC7q6HYVckmYfT7OrLMrG7Co7a2dAke
cfDT8zTXU/yrS3oruzpUFbr52w+jvIPyhYRIvFX3ZgujkitNplpLS5tJXTbN3sCSuUxUoZNNlFjk
DahmMOxaBbEY4giZo2JFgWSivo3non+ZJZu92GEsVTcLu2UsRg81Q4jfCt+jAvcFZGCFLLUsERIZ
IfZaERcofPu7WT0cxSEJVare+iy7a0Cb/sDU40l0bXyj3jaiUSALdpv7ntXExUiVWrQl/Ftl4i71
oN/XQhKYBrKH5zj84MQ38olVXIePsmNbSMBzSEZdRnqve08TiQhceTqzyzauvFWQesuKOAonkz1t
SmW+CWzbDyuUyxNy3XVn66FNzUlTY+7YDTCElLs5M/22FgdckAIdH7+n9FOEtm3C4X4uOyXBWstL
eIhlBC3ddJbhTHs3VUJOyxfQoggbsbR8gtxPREC2bvtvbnLpag9GZGUbsZUhmPoezuvBZ2NP/MAE
Y1chTP7KBAh+SuskCApmdutEdBt6Hl6CbHJ7rm2ZopZT20JTH3qnC9kx38mxaZHPaYHtU79BqfLD
q0AUpMkhmzGzfW2mAEg9cX/071qK+ENHVplYX7XFa8ZqSvjAvxryMADzRoq58Cfq22Wx2sQPNm69
sfA9keM3qmh7V7zT2tkoQuf0H840IiVtr/cCgooW0NudCiCQqXMPGEnFo7qfAiarAkmHJULuO5dr
5cilj1pUGj997sUg7rwePkaSjdS4BX3x6np+YR7Gc753amyImHdejfIYG6HXiiglFXylxKO0rujs
PoeWS3z/tDgoDuWG6UZ7fU9dVImIfUxtISR3ZeWzA8XqYFx5B7bNCcQbksQ/fzj+NC7njQ8BZ9JU
FTlANEvb0ATgLgBrYvA1enSNZoPHwFbJjXICYj0MPebT27vDDJLy7qbk4P3uAPl6mHbR+wGBw5Fl
YHksnppm1uTDWQ3hLHJQc4OvlJJMhqeLrew7Cn3rRhub0Ha7iXx6/gVnEvhdszaOIqKJ5W8y6bZw
H3w3luFp+xSXAiTS2+LOwphfYpqLSeNMUxUyIUnDTs2J+ScAmNQkSPhqHneReJsk5y6ZpUrR1wfv
q3XsoV7RhIvotxCcmCC1d4VmzscOXHA1a01Z0EbTpg3y0DGR4WF0ostR2q3LCSC474CFUyP9Klle
TLI6i8ni/iL9/raZ99f5qLb/QJd7mRQxRXiAzkX3Mz0N1SEC51sk6myIOlJOlE8qQe5iQQ/4j8T6
X+o45CAwSY98XYvRQt0gw3MGkX0Lf9ywXA+SUlsiTiyiac6TNTBCsVxastGUPbCCciO3Buz6H7WP
zyCchRE44nWOzuJHU3NwFeqNl9+DnLEXqHaM/r33PatpOFhFkd0cY2nzK7ZLzR7QNSkuEeOvKGvT
cVbeejCy7557Y8cuxQiO2rpcVl2LDuZinSxFaDluajvSXy5yhv02BqDoKMFcQlsYg/DuLMBGkUo7
DctbZOVhNhKPSUpE8ENFOcfF0HozFOCLCjayJYBOjwEaVmHPuenwRAyxinTSG0GiMXOPcRUt89Aq
9/pagAUXeQiEcYByWtb+//OPIYNnzi2orfCaJYOXNg4c8LgLQcVH4+B096lBK4b0dvEPN+C49upV
3X575DEuzdEviK/ghA9RnT0/nurs2A7WhGeT2br59jhqrS2d7bwNztKkpZG/6A9bvYLNcmhazLKd
AH6JsAHo+ZChhdmPiXLdqP2a8Xl029qD4gCTvtBaPuwU3Lco04WQVYHLG8zxlM5aHPAsCRU97oYX
TXiDTlSCcbwioCpstGyP++0hxvDneHLQamh5hjU3k3BbaIXyeq0yQOcsHTHOxFXC7N0BVpZT7J63
ereBJvxdPEredXsXiV5Ci1OxY3lk6SeSYjtS9s22q4xbIQ+qDTW4+Kpe7JU23rs00CJJIQBYFOwY
LT6hkmbjQPsp+nLjBBYlVCxxbtajPuH8MkqhvEB4WgyJ34L6+r2TZzP2rZvmjvOmsRkFvGW08F82
S29AJiLeVvvkMYzd8lPzBjEsAsN9MOazKP6VFZaEvx/iN4Pgk5DROi4DNiWrVuoTv6qo+2mP01La
Otg2/QA5dDA6r1N1T1B6nyOcPZaUSz31hZSQDOYXaPoisRkvTvHirsCBkaOHrj91rmNDm/0PcMvI
80forZeCV0fxYpJcQLBnT18XTvtHDY696IUQ9IkB5bib51u7Y6nRy2kyhWBYa8rvZz/TbY/FVQQh
LoQqQcENBxyPdNOZycl4sIpq+ASth49fybR3aD63wA2wT5kY1OisPZ5LmBa5YBVJzvEazLN63JW0
WmrJl1ox3u3zpwiDFgwH+5DxUQpKCNMf7PcjDxRP2TJRM/zNc/3wCNL+atvLdDpU9Ls6EHc8RgjX
sxp7zmSWFWqrcF7GjsjZfZfFHpcoz2Hshx+4Lap5J51mcjbyA7rXPSiBsJyfKM8F1898X1xQlhgv
qBZv1JVv9EyKqvnjgupbSFzTLj8OwBVpYYJ3bsmfiid2aQoK5e4lk3p18LfAOMsEpCXFPiJrb0nm
a8i+9UevcX8CwN38ryjcGw0HSsCjf5aLDSPQ5X6B5ElVss6HRw+pzI1QUzhC0tNQCNhJIWkdr14p
yDze6UGiricvClfcHk+uuJnugj7vrdjt6T+I1n9oJN1GjHo7xeUl7Ee73oAPXb/xGNI/AtMSupY2
SN74Vx5lPETCFM/rsgMd0DMPBYBGSybYKVsUirQqfd6MJq4iDYJnXphdbxkTJRvMZDLHdGbdGmmH
hYHW8n0n0Q6a+OAviDXwHjy+WpCc2K9DloymMZhjOgz7/NuVf5B2FGIIzuQQQHm2n+zYOT40Lu6y
Klb++KgIn5gO0tmM9Kn/Ituphn6/nu3ib6bpvDj8Ly7AHXzvKqtmTX6XFFZAV64lYutQW2SCyZQ4
RyP0ZnZ4IpMynDLeLXJwAYCpQ1SV28t7jguJqMwUERykut2NgNLHCJqfX4uFN0WWgekDcwq+WlOA
EbxbfJC+qN1S4XD5oGvjPkHSD9DVDHTPKC3v3sf2Bniu/IOuBn9uwoTMHJHplldFmFy1f928+Ofe
pMHDiKT6ZAtmCteo5TBRVTjPhJt2ykozSCvQhW3dpjwGaMtjje4S1vxPctl8gplk+fW08IF2KrOb
z0Xszy7MH/L8oikF+5YSD3UbmhFdd80lcw7j+DW7XrREz96jQv0bHZ91ryDSuh60gzrxLdwLY6fL
9DDZaTIVvGj8eYcy2Vc1BclJzgMPTXjDz1Q983y+tKKUcwKhFa1lcvr8+vIfm1RQhA9u/PSUIRLK
gtWMu0kDoN96zQB5uOQ4fDWVaXkaCbBwfrtkZ8+DDMo3amTgRABQKLdT3jHkN50vGptVKfF9xa4i
I8AggxYtmRdnI1DHtl/gPEaXQ8jxiJ2z9gUz0AOBlOPc9mDT1JuwvEysEKIwSQXQEhhLGwzuPIta
Y3oz+8DYtdDn5tOgmwHTgvWZ3F+6TawYF34r30fk4wvtaGpZDm3ytSMNe8n/zAuBLPJ2j2QW7B3f
R1fWI71dSw2IFyFb+SwL+i7rHh69+JJps6o1IPXLrLS9MxVEuqPDIqw3oOZDO/amfLDE3F7pNFy1
GrIslLqH32tIyafUwGPp+XgLdXIQrJZKvWaJy2STzpYWt7iwmi/pzJMHAs84QGN+KAyNpES/GemP
lD6Zcz5HvdsazrG6DluwvK9eyx/vRYLy8iOXMPDbcpdunSEP4kIvB+/rM8TRJhOvLASlCbWFG1XE
/DEil35oLCuJNsEombot9cHrZ51rE9Le5TvIrE5PtoG8RdjbL2XLw/PlcDiH9OmfjczFf/CuDEAo
PthB8GD5GK++jhztDrtTH9uMVXHBsz5RNggV1Ovh3nV5YjSUkvjOGOtdeHoTNNhjGrphWNoYmVSI
I1FyLZlIPPGYWdlYG86v9w5iSEfIANbN2W9azHf+3d6Qp23BCMmyt+7HihsH3zineDdguvpG42TS
/Ge/n6x/RqBdkM4EasSvlnWCCjX/nGJRkpx+do0A1P36IMMEJrt6ItesMfc/feaAllU5yyziXBnn
e8RSh/K1Ukz4UhBqlfUtofBYZFs9G6f1hZ1M706LnTp5+jiccZSaKwUD2eLts8tLXSQEPN1iAiGR
fOswZkN4Y48PXydgxYVHasnApK8nu9m8angHSJ/K3mcDpxUZvlv8rad+j/2z9rcGKg8v0wIAex+Y
iHy84kMhn3NAddi/QIwWSeVdZInFVshZDkOO9F1Zze8LI7PlpLCJmlpafo3PKpI9z+nSJStYQoIu
czyeDxfkzXHE4DKOXxkER8TJyR8TLzVlneo2CPQxPMn9pgqpl+BAnGRJFlVUqNfWodDj5oNF1RCv
Z3VZEJh7bvvOGCZYl51kueIBPVjvXpWTgT8z6hMp+HYP0pYIywt7r8s4IsMQgLl2zAPLpdPQc/Kl
Cf6H1rFRty+TPq2IeEdpEMRbdokKBslHD3sOQOXesGOjE9uduXbCvzXeOjCKSgxAnP56NSZJnDLl
+kNXwKGEi3iVVvY5IodBiGE+9lOpsAewhPStIDR/MX9jc65oUWSgicUsCuFPaxA5KkdhUeltGhyI
mJSu+eHD9vL5oeX4a8LSrfYISJUDKrhoV/9Cf+hGzzrStHTvw6nkvJSQv8a7e8ZEUBFA/HzFb5yr
zCp8NQcbcJlqL+o1+qrW8RN2niZpW9wNwszE/NFx4pjYZoFxep333hndgw+ORBCsIs8ZUGBk8nIj
6tPXiucO2w/HV0t+OqNmELfEE/FdWE9danQimlHDPZHctWsxNBIhQoPwxP82cpzgJdJWS9an2mhp
jx/N16bXA2qVOYfV6yKsU6XLf1jWqskO0QyF0NXRyKpZlvvvcOOJYOojsk8LVGt4ZnmtUfvMcgsk
WiMIjMXzyDmeP5tn8TP2z5BbhMHkLV3rHPukzHHis9swextk4F/Mar8+jKuaDH7TK0FFgx37S3ln
W/0vG9MVRtM1/zlszkiJZ+DDh6gPIcSgxVzkynd4/k5aioCWXQxrj4xkyQZivoBihfFpLvyG/kGu
4DcI0SiKL8WY74FdACfjw8aNmhhX3Hx0zj3bJaGOltksE6xfUIz4nN07CZnqVnXXAs2K0PdA0/Q+
owamwRWwVnRYHfHzmkhfnC2EW/B1PZMfCIijxyhx3wnNxREQU0pr39vdKMHn3mbt2upOpGcXv8GO
1cGJUJ/VvivNA1FFKCN7ce/P9IYeDj9MkDrwydCAU5wPlMOlUrql+4f7huT5sKHkzP8ZNuVbF6yy
iIh/gH9/QG7FPMCypcyI8BgOIf77cQLBUgRJqxrJJgVhVZ7tyS/+Z05Q4fTUY+fCsFzjXDT22Z8T
mA1rknOm6eMPpXbm9treq/frjytIjOcNrJnQaXxga/Hys1+L7z1Ku1uIYr8bfW/25fzjDClLzpXo
4vQVd4fXqMsr9ZOC97ocrjgwzAacgvj+Gj9IKVr5cPCIMJTdi0E/VUXLdfFG47MKYGwzGZydpy1u
31POekXKRxnhGUzvL3Nab5dWV9KJyO3yCzd+wV5DHCiKtsbuFB2ZACj5R1AKid+lZH4lR6mASNT6
i/y2gPYceKJzUhiotroDjtvkWPQgPyiLvDypZI3rGNCOY9gDyWiXSnzf8LyPm6q6vEPWv6lEf+si
I/Hv8ZV970f3Lg/DFia1UvUyz6/bNCRYt9mfWVndGTfKHc4Xv2DuErjSGWr69Sd5TrfoYj732bdQ
Fl4VIsAnsNKG7CnMcCrgI5xT7AFUXrA4ZQWsJ/lDfEnXZROUg5Mg4clgkcRjZwgQ6qdm6r/f+Ojq
/5hLzB9TBN/aB/8c3fABoP8VlAMdeAyjgLpH6q0cIBhLzeh08z++3N7Q9mxMkp9WKr7tLVZt9Qg7
YOUhj7CNJJKMRl3+mS7Hk0XLTlIrJ/144aL9M9O8wUj0byWLUevSUVdAUljROpJRtqwOc5/qr+0f
7YUgq7Wkqx4uZfQa35LJ3NF4PVxzR0xYE20/QWfmHpQ3dihibxff4VysGEHSynguifsYhmKHoUSi
v0j+dzmzkJxIWH2aHLajFTx0qlV6BgJXzSHEQFFRbMakY6w8hp3353C25qE/5Cjhr8IRKN4+RH+D
BM8hS1dPxlqSOCHAXEx9BgUlRmdvLsigkC45Ya+qEuFs0e4A0jb/lzilHaAQO2eWqT0Px/bn64iY
hIl2kYNjxnzMedNtjq4vJYxUrCTRU9MyY9vt8Duyghe539UtubaZ3+QrSA1qJBtEukUncD5KDzlt
NVOurs5PQCV5DFtzMUApbEUnWb1+9kDU/lZ3GP2NqaRw15pp5TEnDWXCVOjEgr71PHiWmyqCSknC
yTHGAHrG9WflC0Z7GlejjWNWqGj1NC295XUzAvD1qFVyF4OFhlzZ+PDIHhbcsLqCnQ0smh41Q1Oz
BsXsF/uU3n8namAR5GsNzofSCZjrp0je/j+sNOwSsNxPxGiuwMT3qdQeoix75HU7C4TCbHtO4II8
1/fzIihGbP0WGGJMmXQ+uD3+wXznlbTWODK3OIRAjUKmFaKQWljOGRBdXnPsmtnJxyJsdGM1sBve
3HfPdSvjDt6Z+KjA1ESe+xC+bauy5IVc0SnS1CB7ZSF+Mqn1As2/n7vi1cP0CCfHRDneVlWdHoKI
JgTo+zPI+zZBQKMb5SA/17tQJdFx/Ry5+HSFRTbtuF1Mlm0GnRvRT4QSbz7DP0yrMzvqDNvbIOHh
hVVPdasEnHNmGM2hNAF7Ap9pwCfjpjEDpT3C48nq09ITQDMGPwECVwdcz+GMF3YMPCmqusM4rQ2V
tSbs4m6MI87aowVLVhvgZoSzDwz84AZA0OX8WfGgTDOClEhB1jF4bSmtP3SeXcAw/rK5ulamCut0
Ml7eZrDTvQV1R5N1jurUl6F6Ei1fTkfW8efDy7LATv5Cbwf+4L7+2CXSeyzb7vypB97iGDirPcpw
PtI58VxjMzC78qMyz+11FZUJ0gIp7IFCUof4dQ7Qe7pq3sZURDhk6M4mtLVCb8cZfW8tnFWAjHjn
9Lh9Lq0dHsjcxWAqKWO+xtgmyUbE7t5OaT7kLqdXNjZ5Sm8Eov0XUdNYP0zCB34At01iUBTl1t5b
rpQSlORXNxZUJ2INR2PyAV6rip/Kwpr0Mkmwkr2AIdxn77AogOcxftTtS/pR2c6rl2S3oVCaWJDv
PtcvcZ4F4HoJQOIl9S1F+zcuMiTGVBigszTCO5MbcVC0Vg5TETMALHfObaMcXaYS54uJoKYAhvqE
Ape43IPZw1hWeN0ryh/l13LXHn1EfmROxSyfd0XX83C2eHZYPjO/WSeGA3U93NTgncAwKHKw98iw
Nt0c2127RgbmbZGMvQmB7NSfadXqhxw1+seEPdeF92+U4K/L3lOY189kjfLkOFVeJo2Yx0W25+Py
LBG9iD4fiCSidYU5YFRYB8JFlWFhNZ3WHaz8QphaqVXyz3QCDErXdDujuzpbt2C1xXznB7nAMRi7
IDAq9M7xYh08xz79eSUecNg+fdWJhfHRXAEqjXt+k7PGFKLmTNGlwFdZGQY+6QQGGcHn0gIyza8R
miiQKZDPd/jQaT8kIy33Hgh3LskE4RYfELQpjae0IhIiPFzfOYNpQT0bzQjiqd05lOH3NSLB4zKQ
UUIJSlQOF+IdXbZcJfKgLk99k2xghSnUPdrUf0Yk3G79yVVgs3YHzvGzNMeIQJpxFFq7/hh2lwRq
3m1oIP5OJco2310vB/PJ8AtCZBOg+JVlhT3OsVPYsHkND/65pRKsPIi00V0+VdebcLZr3kbb5yd6
mZWOsnmshiKvaPq7AJ2zG5ZSpE+TbsJCvzUtcHD53qy4web7qiO02RQNtnyNam3ndfe1GmqpUeTz
nb+MC64FA6K1KLpLoVSzcJU/so6oh5nGmiKjURHSIam3OcvS2ZuU9QYQoW8+2DFY+IcpMSs3txsV
gX0XAj1RcUBmcV581t2XdB7S6LXiC9V2pXC6bVqhItWIRhtQFXYOCWnANM3Tk1+rkoe/jMGPZ4ik
Qa4F6w5KLl4vxwvciN04vqh8ZNjMLRMuex1rpzzib3TETH4lA4jtUON+nr31yk097HUZoR27lRZB
Y4fPb7zq3OOtYX+cBg+W9piLxd0r7PFYAto2MOKuGnb+8VXsDjTLVRLSi1lto37z06X2OwgAWow4
vYAWXTDV41brszvY6rEa4iCrfEGiZS8jrFeXMWzrxHs9ek1x6P8yDl9zRFb6ngUkqLbMIKmKUrSf
47J25bBHKXDPeQILCQGx9UWyzFpnjoY6NsZ4P2FaFJaWS50wSMEWgO7MCHR3+EFbNbRP+zZwal/o
jCfg60BzaO3QabeumJ7Ac5mOVglk4BoAMaYGvANlqYRQ936SWBNtMeqqMKLkuYw0lUhwXLyAmrqr
dBoVLUunR+FvxJ3ZqIxvHFez7o4e/+lND0fH6IFS5XiOSWWvawARu0S5Clo1Yqc7UFA28YKEy5YG
c+YET0maPx/wcgRuHYWAv1LFt6sgNHGO4xLMc3TGkNj/JebjdLufYdRo8ra3ovNy2SgmRP3evlDf
GFe8b4xmX97lvzFTLhS/fEE3sxnbMFSe4oX8v7K5/ZrEsi/NpMJZc+XayMGQihe/28QgR5jYfX4L
uLNcvLa1kLvnJPTOQLqKKJ9z+PDsueMt9PT5MHhyjQQJ/4DOI6YOt3ZzQJtVkXcsx4x+Bq2piJO0
N16qJZp3qgo/mqXMUVCOY4o9EZXA7rGn5JBB5gao9sa40MKbNgJpwsYUmrp6rBBYIo/F2lE8KShF
htjgCPQHKzSvhcrLOGiDTs7d45/R7pMvUqgibK65CtZjUuFCqFgGN2Q+MoCAto0AM+R13EZdGegv
6/c76tzy8XL70LBHobvtb6B5RGY2B/kEr215fNCCbiwsu+OA2qvxBiebsZ6Zgw5Qr5K11DYAbyJd
DrHi76pD067+hwSZ6DhcfjgyhJ12fxXImBmaF2pYcMHqDY8r0zVu5ehpM+ThvOSeUEbz4+KuZ5xG
Mos2kwnQd5SVzinOV19riLb3wnaVmxBrEXCVQfjm6y7ohVCycDRH49IXQ5Qdupih3OwGlrvDxlpo
n98EYSkKUkljjtbIvLdEiAvOEt1DA8SomIjzgAbkKGRrCoJwysaMlwlXmt3PDlEeN6c8qwzx5TXa
9sokA8wc6yW2YVtkiWe8P+nF1jXNzKFzsjC4ZY3ccns6RSorXxkJq5/8h20zNPAx5Fq9M1+EK0w5
qvaaMvHk17vv0W5YuxX42DT6ePqjd2dQXai6PZViLynoMXdRdYJzLhVH7VZ7hD3+URvEiZsQayV2
PwmgQjPGJiMqjWOPYyzt8HsfBryKz+UyhVacm2Xli9djh1tp2+EN2a3C52kodZLzdgxYAHq1I6Vh
WAmIk+HRUi49TbcDSR1yOm5yNZ0kbctWQos5MRL+hyeQOhYhFqPXNjvJeVhT36gG2ILWAwXtbRcZ
gtb9+bziJpKkBVnbBbYNriUFf6C12Fk1LHEqmtYeCvMsXUCHu1+zsM730/GBFewX+2UhSCcHc+sk
G/T2MfYt/rZpf04JMiYyPhEcCXxQidDMOWwoItp1IbrJble15SJ/1wIHHiUI70+4HllXXiEt6gUg
4eW9YhwAcXIPCiAfwgciFjTgw1nYiKNwh1t+meR15GT6N/PGeazI4Uey6tFP1lKx75qJgLG24I/Z
AQUMp/+RswDt20QPXIPeWQLSRMlxi94j2crdLbhGOQKghezilqm1Qwy6uDcmMHBTA2Pm8+Aq5/eG
CZ1U1ncOJQqGy2/bqlrV1tvi1ssGheN1X8k70BrYthmByX9tS/3Bo3v/8F2FGjSokSfgMEccy3T6
MZZop9ni8PCLHrHY8be3uUH1DuO76hvyrRNBT41WWdGuS5n+Go5RGXTlqG2RZJOe+e7DyOZymcAz
Oqf3Nht4GUn9tiSQc7qUMewhKzdL4ylWDHEhpin49LOo+BEclIWY284dW/hefR2EZ69AFGKJyjkL
WWLCTWumi8CKAceStSItiXYnXy8KFUJ4i3TBl60L0BeE8ltIjIpCQMtMnsKzKsolmRFlJjNygLn1
xl2pl+cVzkD2KeC9E6bSSUJjhyG8iCDEzahS3fwWVQ2GnTJqJPRNagqjSA3GQ2Fbxhc9bFObAYbH
KXLtflW5JMLhyVK12kL/X1TIVpusrc0QRa/RMOFejMG5lQLLJfIGsxKiB0kTHy1wRSnMZZO8B0/A
JF4/eX7Kw3MS+AH84vPLeg+6n8OX/7Mw3ZRSV6xTWmfm1Wj8FGqih0W9NUkR5lz6MHH/eYcgl9Kg
JY2K9gd6IBHelKC3y+A3Wc1Nb7pbNPPajah9SF+xgeFT0ba812DAkisJMwQdScLlUXTQ3N451nCm
pn6a9lwl+uh+twfTDuUry3DSupQeeBgAiC+S3MMqAIivP8zLlwkS9Xd3H5tlI6EwqG0QeuRqbFI7
zM4BgEQYRD9Cv9HeVSfQnvwOizDfuO03QIqoB2596QKnFIwJY/fXWy25o2bOJl6GqpTEM+4DCs7i
nKNim1dhetc+X/wqUbtjHXd9cQaaYr8Zlb6H2G8MAvGBZItMraZyr7EY976kq+DjyuNwyFGMMiEk
CLpq3glzv534M5hcjMWSmXgd7Jb96AMqrreRhfo6HTn9IKv8hAucPpCw4yp8mecC2VtcYjbY6rny
TPvn3ghg79ikrhGIE/U8ePzJRbHNGQr7OVMo3hg/FNKgsSJPMqetMgnQ7cWrZ/b9CZ2dZQScsiXc
xi0/48lROmi9M8TzyGazcfRAJ8QZsV/JbeY7qteI21tna2Bk/GKcw3CoZEYUkQDRZXYml2Wq5n7r
F8vIYF5EoanJVpflQBNT8hF0mrm1vg7BHrMRUMfP68WqBi36RNuIt636Cx/bifyhVZMrAKYRmnBZ
v5/unIsSx35fzKxSDBJCKQqI7lNzo/j9N8g7AqozC/F3jB4edRb28YLJGaGFWaX92rfruPFpyMnX
VzrUYDYy4dqojBUJOM85hUAM4KWSYYPJyrVP89sMI0NBpabUyZAveuyMLdbLP+/4sq5sSt8CaW4b
NHO9Bitq/r9hNmSlCjkmxJ6vvcAVJPeyF94yNgwWUSO8PUd4EyMZHeM3rMr1FSbCKwI7Qw/p5eYw
PhlDjNNPCE0HJ5xb8RKfpjlh8fZ8CP7MA1RUaY32ugKK1szM6YM0dVlvj9I6v+4i82C94A3new9n
7Yf0CprUIwJWqrzQeWOOjkFYHPJJPoCFRhF+rcXgQpZUlM+iMbTfWNfRZzQ8+RVGzAbKbBv+eEzh
/zKfwthC2vujGW1vmU9p+AWnPcZv0PL30a/NxUCNsbghF/fxpZWHZJAwGG+ZwiLly2DDQv53ynJ4
DjqZXr7g3iU+c+aOUkC0TOsAqRhhnKAndemdpNdBjeK5X5bjrsK6yGcfeXeNQFYiw7EvR3vk1vBX
lPY8mUUNHOkTB7fnjw9HCLrxT1IL3wR7hqGoPvMHfZAEPq7LT8LGLaiOjQ2qJdjf6hN8sNwK95sr
Kzpud6ZavytHptKf745FfMMBxqr4Q1O3WRFpiuQeTZxA+mwaaylT5xaIGerYvihlubcgL7I3ZzAn
iSzr/iDHlRphjXU9aUr3d1sZxuQra6a6Fv+LFA0BoYYVchzU+/9qLFmjs3PUasyUpSeix07H7y4/
AQM2eWK2qZe28r2fYe+qQzNF4GPqPt/KjbcisAbskKO3MGDMEFI6ia5IEEM3nYfeyjDQqhFlkFLv
5E3owity9/DPd1luqia6mZeKRpBJpMFeLDMsApNAdUxgkQ7NeAC6j0ASKykrpmqjH5+0/pVjPC9k
HGYvv+KquhC/L3OywKxXxKbJMAZIO3rwi0HYFiPD1bWHkISlCpbXwvU1/JM5qKgp+CHS6Qrq8eaC
BGiHjIKSbsGrL85MWUfb7VbMiUygGXxVWhfbTAlWtl4c/sRQWnMoWs0fbF0o/ULmZtcJ/95XuXqa
+htxAPrSlYjdiubYTdOJIq7jsHF/rVG78QNLNxapS3S2UIovZ9AnV7wejhQH0IfI8W9J+ur8LW2y
WJMCGFA5wxep3eKMFrYQfveCDoccvp+HeWDNJy/QRxL/YCgZdtr4iITOd/2lTf3SlV9STI29Nihl
Pgts8xsTt5yFLDwKjQHDPDh3JmSs7mA3N13SaMbQcuTqJ1k+n9CWtbEmeTVWNDY2jKveHKTwKhrl
+AdAF/ikYj1VlOmZ6Jtf7ZTQIWuvS0nEvejlVIf7EjC5f0BrfYTEUrvHmyDzE9GVrJIbFfoTblgv
BAfAeA/qM/zZRyDCogUHxlsZj4UinW0yyJYcP2fB+fRdM+GmGP1VF4XahCkAAeUcJdJ1tUhgD3Lh
nFVH1nqvQaU6W1ehtTtEb96xRKoplNpHvXzcjbl5laYOQy+lFL7xznvJjDrXjBYF8QbuZPcIN4k+
CIz4UWHZxnAQPDtXxlFFcsgzlh5ltbe9XMAoHGYj/N911j3TjBdC6ePRQPpVn3hx2RJGg1zm8cgg
frdggVQP3nGTW4JvEX3FlzRv22qHOqYxeN+9h2pxr81FiY0moQKWV1BUtOMkN4XQAycOv4Y/c4iv
U0JOr4G5hSRqGXKSmPeiCecHvrVY8eMJ+tlyAhcUgbUDpGJlxoDUc0BA4pM1rC4HZXXeXgdwrj5I
GjkgbSVcQOldg6dOWuBsafQh0alAD7aVDEqc6jh+iBHMO3QxwvbegA16Q5MW6jt0zvY26j9wK/8X
+S1K4GXjlloUHEjXNzVgMWuhX+fnH081zTZ5homP2jE8k4xQKoG00oXcf5poz1hFf6G+Vi7mlBD9
FR5TXHuTEvXvUPTEnpc+WyROCnQVhI/t2rg+lzKFf/EBqymeiiR9Z4HESzzTK4el316TqhXANfdx
nJyJg5QMPMO5Pu4C/14Ib0cH0EfGz2R+5vIt5bx8GaqyKnAf6dxraHCr3/sbF6asei+WOMxNyIok
5bObomwnjYVbGNX9freZ7UeoNGF8lmg4Jh2Tu2kuaBPBudLnF533rnSmer+i9PrWVtIOooAlBYZH
UW48O6bycsop7L6s0N02MAqHsRe0eH/uF8dL7viAdw0zdBJBOc15Pwx5L7tEJ96s+W6+YuNO8EZm
hoPf3oQfAKbFu6s4R/YT2s7F/SuQeURo1MMnXi6rsoOsGvu7ifudpf5LNrbRMAIGpnMEI2QnIUeQ
8uziU/N+j4JziSo86DrWr5abvKb/DUtKa7YSDP61SD2Clle2YOzreRMVO65JNsym5nn4ZClS8i6i
b2UVXdJ6cvbdquaYVCMap+jTDfuaLsVE9pHFUAO7esoxwX9m3JhYmUjqV1fRyCKfsGUYX01jGkAZ
XR58dihzVG94L5Xb9FWfxhxYX7shuMJkA/L7oHluuxuBp17L3tc9dBJbLFu732Idg5FNMFPgeHnv
x0iY+/VUw5n+TymnCJi2PpDEjwRoGvgY2fytKgcZYnHb6cWE9f+bXuTvZGpiw/NsKRx8CB/baCi8
65WV7+otiUdt3OiNIetUKVuth4IVP+LqdDsJCONPcGomgwioL1Cz5BDC5epsGXGT8q7pUAdgQuQr
0IGnefcVPdoIKsav+nT3yXe4P/qkz0i1ysVioaFdUOpkE2BBt/1XIa4l2NDTEWo/VEkNoXo+q0bv
bFlLzf3/poeKXvhq7++Z9M0xnvFnzLNbL18rXL0N+3ZJS70a2mpkL2McusIS6iJGa+17CpnmxAme
lV3iCd9SoCinYEDqvtOUSO+3h+S/FjnTMAq9l82gYQBDQJ6aPvXuxPOFyK2+5jmAjMlsqfkUiSbP
MYDerToUphftDef+XQV50LRqR8OnIk+b2QTKVbSonjX7pUomEziaRwG1m4nmnZZao4gPksXjVsdy
rcG9S+FHt/WdgVlOc/N3UKs1tVSEpzJBjMWv+kIaOJwup7hu75I0TndeoJQ+15jcoATJ2c3uySeL
OtD9RYzuLy2VJUVCD3sq6J2sVOKYMZuV6XtrmiV8Z5jIcaSA/KxeET6I+xofllcoxCsTdkLO2jtS
wPrxKpCXGzL+blFWn0lwLJCWFovOsHNi18TAkuqtCi04rIzTOGt0NBCeW6Lym93pdvWWmpGfM5CE
1ZUKDH36pPqxIegbPysTG2ENzfndVugjtQyocr4GaTGdJaHcw3g14yu4YGpEAAHEtdzGNCp/lhuL
41vd4k+pni0Cyw+W6hM3+7aDc7B7/4ycigbZIO3iMCReJX6y7g7C6yEjIvwnF0NEwiliNIWwlei9
QwX754oYPBGWlUO6T2F/aFJlYLWtlYVUhtQYHFcOMSP4BKd3mKiiBVDeJnqVtl3kL1/PMOSlHZjy
6Wz7zCL0kl9FrPL8W9n/wy1VIK6wjVNBirVCV4iV5f46RSBAuwNARTf18Cqx9r8PxtGiEIPto1YL
ag2m4jV8BbGQe6v+fiabKWijlzg7q+nVHlmoqLIH3mbKZ1cpe/4lcowkAIyogKUOHqQasWwVvwa/
FnVpExYSjELbRVY/5htceSB35JVGvt92kjByWGS7fRq4Rw4RTHUiHyn+8j3t8RLoUOLuFQIihtxc
RAjm1LLTChC8vavjt8AB8wuSCG8dsF3NUQTNLhxhDOLZizP+gsXKUCI9mcs4slokYZBn8C9jCyP9
yP8LvYwu5A7JTeedc6jeiWvyzMo0Zy9JSoi4rK7/0nxwnNpFHpzRu81jbc3WI+6su0+UZnSVqG7g
HCmZNe35sDH8aERUWTpIxRbWNKOMSchLUI3EPyy6MBDRoA2F3YLSlxqrNL28PvHkQkSZrNg9EdCD
JPwUou0mglIYn01QU5U5rEkrofMQfUqkSl6ShHOcU21NzeWdrY9NE303A6fo9RMC1ifGDmhZUuX1
k9GA7gSd+y9TXPDLT0HsDzf/k310F60fXTdOIp94Mvnns7h7jq1t9/zmr3BbOtIMkmc+MhddTSJC
hbEjsL1jwHtW6+1AVuV5VvHjj6bI2C6fkVNlwna0547sqC/Fpjiv6MvRJBtQGlrmRoI7RGXbdI9S
CazBGDlVOx2jsFRaTu6dbPRIM/somJrSSmBGv5iWLIeyKwDLNG8zjPgxxXRJmcq9C5l8w7ylreab
3ynbHgp8aX1d6yXXFWUIQ9TembqIbPdxwcpNA8DcmHZNITug17t6zYTHn9wwTR5m78ESABStXTe6
Y0+Ubs+aXRT4nWGsJ2UzAtdxXhAUPJBmxPDpS4rCsCrp5e7MNM/FNIjRYvuS3t+J5oBsT6uBfhoc
I7gh9XB2e4ubmooi7DyQ//zTjJW43f4JmhJ5VKT9ePPywVI04Y9iEB648A6OAez5lQdVaOpWYEcn
dft7s7oqYUcDeFx0Mk3VQwgnrD9Yk9JffPw4bL+Uabv+495kmmbBWcCCrhbYmumwey5aUbjhz6Ex
I4BRHzK1MSW0hLSWZ07TWHFyYlY9ZpPrn4XEfcL6xLHq4DZO8OsOdGlsXxUzKhFJMgNGMMjt61Qe
33BY6QOvG43bx8S6+MN5MDUKktAAKkTFUHQMlI/FlQYmXO6UI3SMWcY8OvXif9W9G4+rLAMUKvIh
9HDfh/ZJWrrEQlnCnNtM4TSZS0+qXhOPCFqHG19ez21mHmoupYHFPEgZ8aelBIiIehJphnJmClY4
HdZ5E/065WQRVFcRkYtQdGtz73aEqKR397HPTGwPM9AlzmIJXcF3xQqX4lZoAhJckU4VMQBBU9CR
6TJWdHDB3+n9qKZL4VAkBSWYrc67AThDabzN9pZtq0j0+vNXzS9hLX8SU9MDWU3q/k+lnFQtjVCz
64AXNIR1Q5iuWLhKK7B65/Dut+3xOjuja469QjZ14BjimRVO2ezaJe4zCaX490iycLap7G3vnbKg
T+KGvv8Epy5oDuXn7JKhd2cti0yVTznO1tjEfs3zxcGi2C7hERaqLPGgz57U0yWNvnVkyI0RkTBz
1bacDss6cUaQRKWWuD0Kp9FEw4+/sjILkX5cwc6Tcppu7qREkmQV3Xth+hoqOlGKkPgC7yudRRRN
v3j5tytDjMHp6eg9px4HrwERKYeV7J7uyBgRclssm95N3R1JBEd4qdl3v4xer3Za8Zt4B9luTHGn
mbG2v3EWoynHmR7ck0p5nvp8F5pZVGhf3d7+ux6c8IAmLFuzwf/T3gRn30WRYMD4Qu28FAgnXnbo
XsJBAQ4DvphPUSKZHiq8vZ0Gl6JkXknPREyu+euqNMR3XbNE+ZhtbM/rpL4k6jldOr2mf5Kh65Vi
DyoL6S+Z2q6ZT3ZIr9WsdeHfpH6nD1amB/XMgJChdqVCay7hZw6CtGXIiBH9hZEusoUGHJ5vj6aF
d1HS/tT5ryFK36ExmgchqkCj/H5cy7esXIrJ3al5OkCAySyCvrd/MCuV/z8RXwfSK1XiOWaJCbox
QGGAoUSfhYRTJLceuESwjIJkw27Mryzxa27E7p5c2/3yQQzR400VqQv3ZlNo48/Khmwi1pQa4Lwf
kZ9ifrZkhTlbG26DGbVEBOx7IaFLro62qyV4hE6CBLnkJvfnxZnOQVEwqWW46m67bKOeliWAItq3
QsKVgE2t8pG4J6kRuJzsQhBy8SppMyy4YP7yrC/YTbbCZN5CDpMLAHPP2RAaX4vG+Q5HVqUzYlji
RjqN3Yjy5cGcK/K6dEepwkwaBzT89O+/ZWg6cLaIONuAtiOAvN0yhmlZXMA/ZJp0AYTSCJ9/rwvg
x7c7c/NV3ZJ77VgU8zn36V6/jQU0DSARR6ur2xy8UriuGrGhuGsXB/l0MDJ7Xkiw6lLAkIbrplC6
Au5v3aytyyg/0LAac8QDnuY202f2zN8iRScTNJ0BbJ/cwcnrEGP8J3hBuv01eC8BfxiapwnorodF
0/I+Iq5+MzQlRpVMQlWyVhQUsBSOodV8VKv3BcPdjOeCbDMYOYKFInROKTqS4aYFYAQSlYKJlK8p
TOJpgT/EXThQWmMDpE77i9tYgZ4z7iDwcWiaW8AXCn7JA398BZI0C2h57Txbtw1aheEShvntXc4u
RNVMWncQ3Mq2dobl0DrPGsj+5UBDn+kjNPGpvtRLhlC/CwsCiIlYjXZphTpt8cgGeV00QZJdB/5s
u2NtXBj9NuDrGCCtYfrysyOn9npz+95OI2OE3XnmGdQvzRAmHxUB2ilNh6MutUW0cblLEH2I+yUv
x9PHkPI+KqtFDhWhyWyhTbUoH7Rkq9OT4ch+XocGEFY5s+C52Og/Ij20gyz4djMQCJYXm3zyiSLb
u1Rq/D/P6aJrNgu/yonRkWwPaFTuoUwta1pD4QzMHKRzXNCR0MWeiZMsQ8tbuMKlML36itmOLGAB
tMSv5o3ljTpKZQ2r3OZzpUA3emC6wYuf2qffh4YyZ50b2pJMqibcmgtFMSJaIr+GpUHbBve38akf
lg17nOHUIkCS9iCYzpnuJKbi3SzhcG7+m/t6TbYllzIfwG1goOwcwcb7bEdbJ1xLGHvvgYrdqo1N
uDjFpsiWhW+vI0PnBoFIt8A4WenJEQ7+vUKTV8Q2vBu5k4yF95qyFlwMvwqPmvcHc1E9+Hq8eout
zUFGY/iZeY7+yypa0+Nj6EOpiQ+fyjVImswY93qReHf53rmZC985yLK5Lo0OwB+r1pq9eGpmPESI
QlDXW1ENzFI1e8B3rss7MLiyaW2wLSWbh67C5nfFiEXauAuR007HGDc8/mDWGsubPJZTj1glfqa7
O4h6lH83FHY1S3VyxX+D7SXApGWIUVDb8OP2L/B0VBrmuvYgrmZ6yzhdfAAyFgxXjo4uKhXslogo
EO82smtxup240xZLmTnZXD9wHGiOSl0CRfb1IajHn6A6ogFTKqEAn4cYw1iPAdugerXRigtLYlVq
epdf30/+8+WR4HMGyqQF3glGbSDbzknF18/BF+OY6wet2n1JjtlVINdIyQx51GV1/vZz/AiPk3Dx
lZMg34fTXNaafACkPW+5YSoO7reqdht5Z1t0yDmGfsvFlFCq/8VFZmBTkGqgQKk+zCqPPW2O9K2v
TkoGq4pLwFhalE9roExd+GgntP1zmu/yXhF9cQlgR26n27nrzzqW7YGDaCt0341ySaixQ8hpFoA9
cbKiAqau6q1Iq5F77SIEJCaIpKcI8bpGi17YgvRgNEaapABETjkSLOgPxksoa/IEqH7ClJGTIL/j
WuSoaxh+dtuVUnSK3NX/Ke2ayD8cgEZ9z7zaADiolY00WkfyY15cCpX70KvHrBTgk9p9OrVsPHhO
KKrzGui0kel55KXYzaopqgS5HjLL7z3CMSa6jQTWGY1KrbqeYPe/hYPIzybbirB1LusXlogovX3y
JVMSltQJHJ8TNRWW87iBUoET283BiFgkTFymP6x4DRjzaR0dNg9x4OkX0wOPVIZZQzcq425RtSpa
qI/UWEOksUHsW79Va/MPRBMHa1Z8RjdJy+OCK3RImPkQZl2jm1lkPEkvIlxSmCOHVMEFv61RkGSW
d3QkP4KQM49m7dA0v5c8iDPjAj38JbBQHJs0lIMrlNwAPABDZAnZD6UXwLxkagkY1bN8sDQmh+0T
hlHTSkGA+JwFo12LHEhGepx9ApjX4T3x5m+/Z3mVuMariuukj+COOALHUcJDy/gRVk2EsJn9QjAz
YH3gNNCjefPJlhNoSQOWxFtjBGqyzw9fT+lpZ/DnGsEZnZSdUQQHguVT9U+C40m/5/Lj3GB+NPXE
cRRdyzMgu5pPkwz6fbcrVW/7H8pm25qLnqe9vBwfIBNgzq4qnJ9j6XQuFuJFksZbVLGIaaSNiM+4
LUZJt/znw7WBlUkqm6a5t5gSv3yg2OqJq3HgSLaygJ+M5bpgGdaD6cACGZyejSsoUcM21troTWnN
AoyTP7vD7wSC50m+mlyf0oTldPtpe5Lx1wsAXxXgTNlLzRlSEOCxJaa697BlzyQV8wOuqU5/6yT1
ImpAXddTcHlhlH9hRS34Spb1Y76uNNJGoH+owHbEN8GrOZVXp4PRwy1r6UfVi+3xZ037mE8UNiK1
FtP4Y41G5jNd+d/gQeuuQw7LpmRVEgzzg7/M8eT3EPLviCubkIGRDzL1e1x59L+f+Dnt2Pn3xgDZ
oVdPW2owj+mXw99VmLo4tME5t3nLQanm7kWA86xC/1RNG7wrrUVRb7D4JQ3zPf2timZ/Q9rcRtrq
e2A5OCoNuIH2ZTqRBq8b15kB9S7T8yjCW0I7u5USueCt1OCbU6fOoSy0hRwUlUzAD5CCJbV+ESn1
8t32JwZdxMCZZJgwNpMunT3VMpoS6DEuov7wVfuC7bDrFQNcyRmWMj4dAQuuBWLcps6lXTvfVc7n
0f2xpvgKZ22JIft6RhG7khsrcldHUhSE0v3DSnn60E2LeS3MLF1iwJkwK3Q6TkU8GUz2D0YV+GpU
X7gMhHaCN8ehdBIeWb5did162bXtrwYAHMdN+8CrTYxU8hG4y3QgZFmtQ6CtN5XrgevXw4weE3r0
qM8uxmUzPcVySRaFRJ/Pst/KdgR0pneszOkKjYpmIVavmRRQRFA50vpdKW3XYe2mPTiDSMxrYwEr
qj+bNeX4vSkNlKldnpWEE5zw5NjULseWBeBjEObCLPrL3+ZpWiFuzVVa96tzMa+9Xpt8DD7z9T2J
8uOovO1g2Ph+VZTXD/w1Kp1gaPwMRvX4fXO3rjRQuwtf3zmWj0WAWm0yMy7r/ymduGeLJMAf7qvp
9viU+vdcKTecW0TrkSphQg0b9JjcA81yHP1r7u+EtxT4p+py1rU47gmoP2k/N5aeF0OhuvxNY6yp
SiY95BxUBQgA3AFvesV+6eT4I/ipO4XTIwp08a7dA4a2BbFOT8nYYCyceVjdCc+nOaM/LhGNEB8F
n7ir4LKY0854Io+gRo+na5drqctLYrA404CuhjjeZ0yaTTJYRXMeuVDIs6WAZz54Vr9dcD+dHMFb
5pWWJr5auZvoWlW51NgrybJ5iEB+ybcIAUWLcaHQv5WtVJAD3i/Fpxkwix8vHWi7Tp5SUcEoDfHk
X+ptvygMKymP6Caot7CBdjSR+cOVi34uQ7tx+z8h0TIvMWygx/RfXnLZEGtzP4UCgXPT3xpXgBAM
s/vJUtj+cEskOlNPj0q/R/R4/8af+7n0Q9gXTKxdlm68Iyr+lzXKHk1oaAzyZdkwJRmVbPHUBkgv
N91N6UkfuBAihVy9ImgTdA9vLSM90suPByEi1o2L3q6G1P0VTbsc28av91mNuCMAuBe6xYuFSa54
wHh2gnUapUi6zYyh4uP8UXYr0QwwVWEbX4d/zT5rZJJsauZ9KV7W5ejaCKrkgDlpcbg8kVOODX/v
aHxZO4dSTDt+UrXsu6ihi3yivnmzzVPvJ3z5Ybo8It7vtxrVj5y7l7LoOGNRuU3BQVEO+G0YyOA6
qsfh0tOIas13siGc+5qSpJjSDhRgq1NPHWW2OPXGVVqsjgAxQQavX83jmGKDxqLZwhSzSn3JJbDp
Dr9TyEviWDM5myLFnEgSP/kdQ0G70Kc7C2iYrEEyv83jyX/YlralNANL8A88YyxtDYpY47D/JEa+
Hk3L4u/WkZ3g9WExsLfzZ/OYYbCN4LbEgFzOyUzzFLQUbL59DTIR0moX+qunTb9t0qD8ER6UXnF1
4mV1OwIS7e9aV+DGtJEUbO8y7fV0lKfZwyZl71QxtZ4ZIMjAHbwVz/xmsykzhB8vbsjNJWVbv39K
CqC4xOIwANyzkfMkWInxlHIOO3CBGS1UuWGUWheEniAGtDmY7qBoXpVVM452C0b1IEjFP+tlysog
NcdL69Z8uH7oXcXrRg4uWqdMtbUgA9wffnBIRpjZ07a533OA4+j0xetbM2XaBqyUkgeV74Ztzcd2
Cn5HLApTovbIYLWx4t9yTXPBCjR0CoRmvUHsbxkCvH2IvjATPg5joC/hr6TxG3lAtYHfotsVKFiF
htChU9hno88+uNa1hTzUnRntvuCqXu68cHzoiRsNtv1wlWnvuXvCcU4HA0ZDek6pVipsxaw+GyWl
0m0K33h/K8u+dAtnyny/pk2J6deHOGn2kJD9txDB8fYAWK+svPk1+PqcAgLGBaEF8VSyiYyB6kKw
xHiDIeZQyel3LXcEnhAkLU/fS5Zb8L7WQ+IPFgiqreMBP/X+tLQZcVZbtqegFjISebI0lm5xk4PP
yrKcqjQKeByWBu9m7aKg3OUiC3DuUgF0JMXvbWHmyB5Dyv7JfiLCBviRnPwITfKhKylTO071kM6Q
QhUaH1dPhsh2IXXVwR9LbC9toLiRavMH0WD5o0WtoFLZtIs9lG3c0seRCdZGsAeQP3qf1z456Nyv
cabRqt1WRcaE+/0RD7lfGgTWDIuytaedU3GP5afbWxO6jsxhxtzIvHbin/alEO/Kw1iApXjUZa9c
p3ptJ5G7pY3q+XBk0YhO8pMrj/FbTJ1mEG+wQptsW4jGa+ta3Hj2jcIXxZyKyxbvHflT1pp19MLq
rOhzLeSfJzIMJKCSIlWdicDB6cxbMErptGu9lDWF8TPoCeKDcV94hMpNjhngeZ+vJP90I4J/K6f8
nXlKY8NqHq2+nqU74hhZt4HbKi0j910btz/flslc/s32GOHPKKJK6hmLhrAor+5dH8mp7GXxIDtA
4X3YS9V0RxAvE5fupCynonLnJDIwb13aV/vyzv84tBkxZQmQh/iYXoPI4GonuXv0k6TreUWtBdO2
PDEu2zvOpOOSPiwXSw2N/3tG6MpAdbGmf/hWM1BcZdt2fmsJUIHiRefqJnNzCDTxqai7cHOnsJzn
lywjJ1Of+h0fogfRf8p0XA2OlskAMKRPzk9c+XWcA5srOg/FAGd7UyG96eQvJatEwKXY7FFeg0jV
D3i0LkE8lqh2vNnCPLT8HaDee2l340rZFCkWX8M5+uf+fWUX0ZS+LCdpjZF3buOCc4zdKHHZzObX
RwYDt+oehWO2tMbBCHWW/0RPpD8nX6W1lAVHg5B1cuo5sWBY7V4EBAmxZkG8UC0EoX3CPuBOpD5+
sx7Z549frqttshBOb8sp9i+OxPVTeeZHa3ZPywQWwZRYC/r5dkp9XlnZzzWttTrbVsDBw/pi6KPA
yqMxIrNSDsTiQPbfgYsKF+qWqbgwXqFgGMjF1QLK6bln4TQ/n1aqlA5AgKpZs+1Agl/4hxFOeLuf
RndKjcP8XM82brYJPvT+aq8ZJJ846rme/0i0kLJvTNCe2/ZFV//BSMd3qfPiNCRNEdo8j+kjPMA4
UIfJimTH4Ym93079031cwU1i3yDBNr9+2MY8ymcQ+Y79TNIrEoNDRxrQGrHCSVXILauyrI+hv4BT
H9jPWSL+GliZxc6Fp8xYmTTXtOqRXuAGv810bt87TYzAy2j8er1mxa2Rx5tXkDfV1sscEWzqJIuD
f4H7Deein/rfc2uZbAAi0Vdqi3Oq+s+qVyuMT7CyN5f8x5ZFWSlv/ziaOzxZJD0OhCK6tB3n64wh
RnX58Rr51sw7P91afcCuFVRjxy0ToAarBKC0bZmKnnckQStViwZam5btxESWJoiGKU4v5D9M5HxU
rnh0Pe3h7IbJtFv2DQ6AhyeqNQ/pxa+JGSycTRehNzQzEw0dKIF2HZL6dW5uDAhkRn9huJchFuaf
QXz8fwfBAzZqAF5JY7J+LNtbuXLFLrckR3NzlS+NKV/+yzH3VbTP3BqQ2+5vNGBU/YbyoLUgVbQ6
nC+HhdCpev5+laJMzHLEaald0fCvc4/XQohVqaEmjXklraUwiQczIbAxo3y8aPDAfq8UhJ5m0H68
W5yL2yo5DTuKnMxrmx8NFWsbr1ogLWLLnorcAbG5kIZscvztdIiMFQPqLKx6nakYrEk/SkdfNvt1
t0jLtQk1m98rr59vsrv2p5VwAbhK7jE2ATAeEhuhVIQN0WLQ52yjNwpkQZj3nr8vba8NcOylqVE2
Xay7QtBI2SIeEvdbhjnCXkMhHAgAPXGpYJ5hQPlwSfj+PqsVxwGDD0mleq/ITY/e/ozVCgVUsthQ
mQzmiT0EI9mkHywj6UpAi1bsD1jXWcJr91BL5Mo6jIZ7ujw63iWF43Zpox54wkGoIxm3n5n+8YW6
yEQRK7cZEEEVivbA8rZvsnZc5dVnia+EHHaA2ohy9R7Ncwk50NVsDlB6C515/nEkX44WfNZClIEj
C2JcB1FvYpRDFSiik08SjGdqEgmDYcyP9YOEF5GrFgAKE1jW2DV8o+nmI1DIZWyGdEE1ThzraL1o
j0DPwImaKGbTPQZolRRjLlNrUULQ9fXdE8hlC2G4OlVkKlXTo3a5WGg6m63M7qOHkA6EJo3+15AP
YAvlHlQAEz266JCs/Ounb6lrq9Sg29LBFAdVm5OZi/r7sFP+S2HSAUikCOUPAMm+QRHHpWrraTFb
plzSXpVPSTwa7RPKUp5VDWty3vvVV+uXbf1x8NQWfF9ZrR8eHht9pbU4syCddD9EzHRzpibs2Nb7
/2xMtIXhkdDNLtteMiKnzL+PHIbonBipTCvG4uDRuGKTD3yVtkXW4EhNezAF19wC61CXv/ARRFTR
MnPCZzRJccHkl4BbR9gDZjI/0Qq64nPcXhaF+SXAukC7U8h5GHBzkqMS2sTn9MNtT1nVRUhnvRN4
VWWRx18DWLgTskzHNQfWHELxbCecxGxSK8KV0BcyqolOK7UfoJGsjDN5JxRcWauhmSVPs3FBuHhD
lDMcFYfFEpBR8OQZcfaH3el4+32I+OCoPAJyQoxTvIiVpagSEsnoW1rDIut+hA/p6TxDQCkYXfBW
wUTTY7ZMRUkU3nbzc3Ru+UmirwnnhBXK5ItceWqas3vhW9PhA7NCxrJ+cMFqMI1yg9zkaM+Hd7Ii
VPRnebezdxGnFGh3pnCq9+rYkuvdEg57s2Cjfvcklji3r4etC8TXeExpbMUzG1LKRc5LjR0djaTh
ZZvthJe1b5tAUWlzaRfF7je7yrN4nLGgLyXvxLEJDpFSZ2U+7DU9FSsotD/mpaCjgo5zF4a8vUrE
CAsHM7fYbSS2DvhjjwqtV6+WzYjn3B5hn44zhA2biDyg5nh/KV2RUZppTPhEG5dBFoyxiGaZVHX/
VurjNKU9fNQ4YJppvNqCfo7i8mRvB9JbR/liYkqiS3m5ANikYa4UH0j5uH0F49koWvEmGiKfmu7e
neimETZV27x3oID5Q+B2fpWZEa41TCLn9dBOsI+ryv5sfgDc/Ln1AN8vWpFJL1hayBDdMH8eeWuM
kRKIAqFMszJFS93e5+OAe2XOaYzw4DCFA+ffFQN2Nybh9vzc02c/fx3+QXOERKyOmJ+ryBi2ISE+
uc9CppfTDzdFJMoQH9qv1YsIldW6EW7DyOzPI7613naZRdZKLA9UXPjQhgnbuq/j2tm4J3WisPZk
LD4EVl/JDdIis4O9Et7+i5z+Ub7glNUfspaODewfsnhES7NTPtUFOVt4vIVfSYkb0P3ivtaCoWT8
ejZeTMw7QNhY/FPqO5iZUzWYy2c8QZrANuND+Xnc073KSIzoqRBhgf+e1XCqMY1bCD8oH7CwZ+za
1tc2A+7qtdQwAXO2TgxP/8VZTIAyckWQThOV4Po9j10JdYnLeq2a2gt+OoWed0RAiGesprpIuizH
o4z12FdnImxCUaY3xtGiZjkua16YzdDokq2hWzZS6bkUh3cTavVA61W5IHVT9bO4UenbUEC+TC0B
9LLIIcUin8xueRYc1iSe4Mq7YSwofShfb3XaDK6c577SntHVZO8RvkpyxszWZ/is9r0Vx7bmjOVc
gAnee6/QZD4MQfXUGzCPH54FhbxmTW+N/Hrk+0Fd9l0q7tueLCQq4qPHFrk7xHQQEtctXhVuN7Zj
mOnDonYQByxpXKUR+rJ2dH7/LCxK3iXJnUgi+26kEa3j4iRZ15LpAxrwVpmih1BDuUhliw+PxWZu
S0pn9VVyqHd6v0MKZTuS9Hckes2czd3xTKz+5pqdpbJ69P7JeI5XrAFIYGOnKr6iC4l+hwyKYTJF
ZJik8BdD4N8OBL8Q0g4p1tqMaKR9oS4BqPGOE/g2gNCR6yw9B6OXbll3xvxM5xgsSeh+PUIW2rV/
2kdm5tRd7MHPPpy9qhE7hHc8qQ+2A5omcy9AuffZicLlCpDbmSDUlKWu++D/w+rA7eyTYlFjF0Z8
w6v42huemrhj781Si14Y5h/Q0nFpOvQA+WPz/f1FAtE6ajZaAorMYqVaNfLfuVRAzx9XAkpt/QnJ
UL7jJPwDX3xCHUdObpTNE86M4pnwgFYKUkOaVm8h4SFw29lzq1ewWFz+cAWiX+Dcv8xQwubMd8E2
6BYaHGvao/vIFlN6jhY70thP34+KcRX5K8YBbgO7pq3FuufvMHItGyx6gesZNoN6RRKcIWq9DczA
9sppJ0LEjTccwhx3/PvErWatLpMP7w1iLxflu4ZOxOVbOHqzOMxDqJYt02eHcMyq8jzu6+QfwD9V
oLg9SBVSUc3il2r/PO18vZIZoWO0sGt03pwajwBHH5y/+koqSyOxPQQx1Sg4Z4Yd9Exn5fJT3+tA
gtSoaInXDlVCcpZEddCvw7HIKWF4tGO3Xu8ZnN68woXpPlVl/F5KXSCh7R+ecB9PY1spfoIMne66
AMWMFC75wCHV040sW0u4PxQpnEOWmFH+AR5w3y9GWitH8MTXLaL6kvWh4F1UBEs1RI9q4Cruyao0
u+XF0KMyMgUNm+lLUndxl5fYBKQGL7sjYGnrNXojigmgoV2l5TA+QnRYVdeNsCEK08Y5dEb81GEl
+UqVHe547e0+UjKiuDCVCPjPy6zCWLzUD1D/i+R38wpb3tPkGCd18Y0CJimQRbJz1SEkaxWcmueX
zUlhbWLS+wPqYiMm+385a2Jcnxgkpa9gCl6yp1UuJ//LMY5FzWhDdS6jgdfq1q6JSMPj7i/c1xI2
odoAXt38R2vsnWxh5e7+sXqgVMxkmg9EHb7WLnvPkQEGkIc7eyJEYI0bP6TQE2VuaJdQH0rW0Yvt
8StwB2qvJWqMCgkOkGwAehC4i9HpsaWr4IkxImajPwULCRy8atidCXPxPJ2yg/ZpD5M3bPfFVG/J
LEreLPRB0Emi5fdbXTcVIOpAWE3Vy57+7vvTbggQ8ILK40UjKsOvHJspKSTAksGeedttCUCe5f4J
/gtN3AoaUyw+pJqtX8hm+K8PapMCM5JGLtLQEk60aPAxERh1HGYUGXOdV2U293gDJ2wzUhTIUX97
bxUgb0AoqUGGA7VhFzBhumXsxw9AZKHbJPK7lR+NYss47RebqJSAGWbjt7w+gskkcCdS6JjEMXyQ
NJIGTAMKU+xgUaQSM4fS7HO0Qz7lZqKJYsIxH6ezocCZXdABTaxkGDtMYQBdqXeEmd2ta/HKyUag
fjPVLXeOmEGScmcPez02RRf9vVJSsGYBtDFlpUCb7OReL9S5qx2pSf8kA02dfxQdW24EFtcqh3ts
4U9pBgO8L0IPtZjYwGGNXBoa+4WcUnNzKgJio+uyXEqpF6ITftolEh8PFV4teeqPrXDdA1e22HIi
2Qr2yO/Zwni6L6FJvylfU6onTmvqP+6yzfIvrR7VUdiXL9IWjlPUXaftoeuWfZWo7c9IgcKyjqHT
T2Wl25IxKfqTsg+vyGUO5aqh8c1h+2L7MXPXK7zXVpcFZHvv9qntLxahk73UCCavAJq1ZfA5fqmg
4ORloBCpvzjHvpzJX2qCh0kWYL1ghu9g4QMdtMldnS94+iFbY4vrFWosD44Ee2wMIBzi4dbrtR5w
zSaE5ai62nIhBYSpaytq228woSVBimFw6My1AEsUs6L7Znfmui4W4SlRF7DGbj8hb7B7YtUZuNbg
TdtQSIMXvxFYqcLtupFUZf7csWB9tNnHsiEb3yMn/oBW+1joKgof1RQh6YLcpHQQR0YSoybfT7iT
L5Q1ThuiYWKkJxSmXOSVcQDY2kK6GcrM9encEj+SM9ZGkByYfQHiuiE5gSNQSY77IHFlqCyJwTP4
ZQoJpRZq6z59Iui1syZ7pa40UgIOeCbYspdegI1uO+9fpEIFyIygDGoCLBTPezRCoyPLkd9IzAxU
DOPUKkaSXt18tiNj2SmtFlOjpDOwlrpVq1Dd0RSqK47f05Ru4e/7DgA2LMu+2Xtf7JWvqmUC+fcm
+tpMLPqEu3Mqu4uRyVweG5pOKMnYfgKrUI1JUPT/hyOcyjf5h3oK6Ipah2/Doebj5hqOxUWkRGRj
B8zk65I/JtoGD7jOgx17WboYt2qLR028MPvksBW9B7FxTSahs4L/k1hvVtHBSY0dDCd8D4ACozxv
b1EN0+8hrjyB7Wd2JwV8d1tFRPJIs3fgc0RhB+6NijrJI1ym/qZRcj7RUhLkvXCD5Ez4VTjwLbMi
BIsLebZK/d4W8XW4NXSvcKI5lBu3y2nMtxFCa2SGTfaxR/xFWZA/JLvTPECG58zsNcEfzXKKDwIW
G2aYRUEYqJk3RKwR4ZelUa+bUjVK9kA9V7A6SYICG88+EkT0RWl7sqRTZkAfFqavg1U+cHLx2zsy
oHR3TDh6O3srMyv7c0dZB15ZtH86onEeZO2OixkvbVDEGz+3lWexQk2W3al13vtDe2Hmca2GTm6v
xs4DQ9aiuNT9Hsj2TmPc0VzVuJBw4Wi/HbpuKm0U7V9nKXlDzJlojB8Zq4Cff8GvBlEfv68OcRnX
qFaRC2k8pwPi4pHbUzust7lgR2+WK3lAt+YC9bsLnf94muRH+FYcC1eYQczF+PZUeCFfoPbNHGKe
jYRaasJ9U6y/Rs5/6xDj64xMgUfYHVXhP050PYwE/N69Q/8Ky9z4RUAJ1CJFD9RR+g51I1O2yneE
AmtVjO/NYg3kY6vE9zj0e1CJb/ckr2YAUJsE717ZCV3sk/SGbcVGMnl/ivnixrZSA2AjKEgv2CpR
XyneBy0iOqg+56D5fgU3JhMzqvW+zLZhLs3znIvJzVPzD3/RN01jeWPb/lR7cps68UrpQGR+sLUc
SN2ypJGiSKAiDTx5JZ/EddyLEezPwKyhaQBSOsk2KfA1DVbtdENWnGzNkDXW18kQDT06Lhpyeqh1
hzRudxd/m3GPyxwimo3gAKGoARlrl2oFP5twroQK4MdJxkXmh4DMFTSzS7a3CMPReqyifsGjjxz9
XL2aoPIC6gg4LXcABdUvjbs3qoSWylRLYR3HTMbY0kjGtKD6tMXL+xur+EAHkipslGGMRET7lNev
zNxp45bekwvQWO3md1SrdPRz7X/WcU/fE3lpfFL/0IqpY57U+dA91rfl2D063m5pJ9m4KCmDsi67
I0TOlaEwciJfigqkeJWLCOEjdfof9C9dvehTnQHRyTaND2hpcBo7gOkcCH49NLhDawEDu3uqgs2i
pfpnVwotFtXoKZqL3QcHyhcqGI+mzYmCjvYTTWc//m2V3VrtMFYqMV+oNG/rLwy4wBFKfR+lgBAl
AiIgP8luHcbQcKgnYL5dSvRa+7nwqo8FxBWV6aNtU/cEFFqv7Y1RVfSGEB8PUWz1GNUixotN3dHk
fSM15yk9NSU8hCyUPlCqjyvHvtof+N2xNqvXjMSqtb0IwZWkiAeukdAjA7yE7a70k0i/DnmBxxkZ
ZfVBvhVTGxMgw9sNUOsRHKn5sI0KnPuALXoGmQwvamqWPFWFMrEDzTbx5ZSj8zKZIZvm4yRUImk3
IYT0US0WcfZT3GC0/4qnIJqBi79bbpPBdv3Qpy11RyrrU/+4ge8YyuZrhs9GAZW2RGpUGxYQAG9/
cUenykEHrhup7NiKWDxO4Ydyt8NFBJdP2/ILuZ6A3N4WINzA2FKPj3fG+/xu8yRd4jZsWjj6bxXS
bksW3KUVXsuXWzWjIU4Btfy9fdPUK8QkbxJXu8N3NR9DAyyNKkbtCsDo5qNxaqAv4ceSm5uMZIXI
9Jd58ltji9TnHPznuaTurdnjrOyLmNFolnSbzlf4NCP9jqHjOSYt87CATfoFkcRb0wuw3MJUY4xV
x1LQFwXLx0ug7z1l06BLI1EaCbyrEULH0f0qGzwMqdpMPzS1OlZUKgPaRKMgsm9Wn2N0zZGWp5za
yZJR1gR9050GtfKQoqvFGHFPWCqZxy48jme2JkqLE9JQlM2w2JLPwYOfz9Ew8YbgYYjTozs9DxlQ
TefmsWzD4aPuqpEVpmIrLvSQD04VW59S0nzEegumDOKLpCOjyiJZGNNsNcmF6lnXJlSnnc+jLhKz
vkoJXpr/l93O09lxPOk/eJ6roW0QM38jwc+5Mno75RbOJ0h+PABx3MJdqB41yANneA7ZYY4BRbQH
C5f+LrlFzXSUrwzOxfngH6fkLgCMT8vGTdfsj8CeHKmvX1rjDYqYWd9HDYcBw8Mb1GHEimInKUUY
7zN465IBmNeIq9+E9hQmwgyrpl2mkP59qL4XRJi4HHkqHoKAMjnf1JIjBvs2ZjaFDquKg3CETu4y
HpeE2nBg2qSiAjDwdmtUJWW8rbMXuq+8USmrzszPSqdG4ste7CwS3SiXbpnjue1cA1O3vbUzL/bC
2/Ti6cJBHK1w0gjmzw8n+sCvR6PFWmwjY8y/l5KRLZQWySsIixB5UiKQxFeMCLHac+jIF+HnmKQw
DCLfiYFuExgiBIWRBA7evifLtFQxZfcdYyi2KGhV0NOssxxyRCJlk4MhuMds38KpZVva2FOgFBmY
hxouf6dyFmZskB9VRPAK01M6b30oAOP3mhDX0DjJBzw5D5R+S9iw4RlEWxQjmNnpClLXhGffpolI
3J56APWRvZNkqYGIks65aoMA6j3/pQO5Ziuij7mzn5QtVS7NyKzohLtmClBq0YxMp5hPHmxzm3Vp
HCKrxvXZ2X8eKBSD2Q46eyJ/SNblwwAcOajUrh34hl/blETG8xxO0391tPyMu7YEGzjO8WTjURhg
iXK9JutQSDOkXMN7eZrgELQAyiUixFW1F/Qgk/w20tzVcfnT3QnpAQuRvBz2Yvnm4DgqEKg2A/Le
KeCx/uEi65Wy/K3NSqZ57ujHJc30GpQ0B/Hm5zmT7u6JGsrtZ8Z3D/m0oV7yl5qCqvP98fMxkurV
Mh7VteJhMHYFr6BBtS0GTNqAi6eZo21WBnczEFaGNfjn8tszkvqPeMUJDKod2nV5LvWoUt68MfoV
fU5LdDpE579zo007p8Rw/CSHrQ5CHo/JZj3TZcUfNm1y9ndjnua1mEEUvc+cl4wB+qvaCS310BNb
bQDEprpKzUUuwT6OwZ+ij4uLt6IPZHA0MGK0Bd6OlHNBgzKeWa/iylup7s6WO7Jwlpy+Z4X6I1D9
DMXcA3+bhAn8H0Zl9kxSNfOO6Ovb8AVHvdm8sC2XKLh57EqF+sRx7xOxXlUNgB3yWh/klG1n4zAU
0VD2k8NiftL92SCu0EFVOttWtIK438gfr82BVB1ennRjgEV7oYLknTsVJFrlkOGcq37nYSuRT0yW
BWJ69BexFmT5LZS6ncyGKF1i6OhDYJYesCeUX22m73CMsUJ5Yq5+A99Fv98x+H7lI4uUjph6FCgk
6mZx9op4arvO0cM605SlJBuzrF+2hRe1pV1lWjzlnSvCA4mdFnE2rGMOwnHXlnIoQB0Ml5MPxEbx
L/YFSQEFR5Ro2/zJPqH2fMdPn8+SpCt1C/Hxl1Aq9Z8ah8v/MSbUltOM7Uwo7iPzcjcSybfQmHyj
TihIAZ4e88yutqbhf/vWZ/Ab2DoNetleCIGVc0PhiYQIyuYplVWcASb38QPscB3amfDWNUTJYh9S
Yl2fl0qHJ5BUqqB+CSeo6maSn4XP25arD+HxfclP6QPfdRM9hFsmJa21dPRYvKzcChGyKZCkXgR3
bZHS9XQfjLur1ezuZpB0LM5JVOVYWyXmdrK/L9z5Wzvefv8P4X7tH2DZSWf/VvHM95W9eZv0WOdR
uox5yXYO9m1ArFUFBp467vPqOuwAJWLEcqyhPdW3d/UL7XKk+OmSIRNZqA+S75V4wnSRqxbl/IaW
xCoAUztIQWoLYF/TfABAhmNiJEMqm9V26LS2ZNzabS1q2MuwO6yqdpBAKHtZtL7LORSq4XOYPp65
CpBAXl42rdWkwHcmRBaHpBBokEMU2HMJzo1BiE3L8T3ltVD2AADhHgHgr97wJ+UeiuHXO27WPmni
Hb4YPGyeFEBEq4vdGur3EIMI5L6OWswGmOKM6Csl5lZv2okXyhBDYwRN63SSrpqJVxL+f4GskK8+
vUIBSwB6iSoRJYSGTmb2ssr4uUz89GyifKY1KiDLcKPUiMtujWmlI5Rtr2izAkIFNpjrtsJ1WrAT
VUfAeZSFNjHTpTBHwrheH88UQJQKV+zq+7OtiFZjYvv7x1ORwu3Hk3NIqxC4HaflN/I+YEK7mMNQ
FX9rDkDx613epLWiieu2E+BiAqwASSHisrZ97HaKNneUQXqrwjWiCL0Da4W5rMqJOENho9KT5owU
HMik1ee6PmOI+AwyHrxxeROtCk6Wl09dkCdCxxkvCxx1NWxOsYBS3c91+mYMZwnplwuXDCLANISG
rtf6zPjQPTcTnwMZp28lKCnWTteFcAgN19+s+ozQOp6a8r20aDO13JdKDjNPjWZQR+ETJuotYNld
YDFItt0k9AjTa+/YIan8LK/9xovAW9KP32YKY9wFxR1i+HC/8FBc6ovjx509RuyC3TdQszL6u5yN
x+0VPp4frDPWIzXOTx3u1/Q52wjNJDAYMoggNSnnE5zfFwwoTXm+BwuwL93AsfLw7p1AlpJjlkAj
UTOQqN7kSkFswwkO6G4FNiXhbg/HJWA4iJqKMl/FrMBAYnU1m8tSzZEfIn2ZpKs1LvY3HYBAQXQ+
cMDvbbIVCyRQVgDhSHHiEfXLwyhnQPvVaYFtGFPpuxoHbM/cTe0P9r6qt/0gYG93SyC8wKDiCMC0
dwq2jUaxSJTdbe6L7xKtlzkU0DLCQvD+a4tB8layinEGIM7jtQuPZUoCIVyDm1q+zuosf88DAGzV
0RofKfSGpu3kdmWC9fwLCAizT217lbSPZ7QJ7AR3ZIljtlz3RU656/kk+cngd0Jz5BObs88P2zoB
pGM+hReQiMfHqtHbvr3XnS/cRyJIiKmdXHmjusDETQVq///Y5vL238/u5H2aYn7mFxFxQ/taTFm3
MwRy8tzU81d6SWrho+HMcibnZRd0zCjbpagURU3aiEJ3sSpd3DO1JfcyR1369a/5sNZmAQIrWNEd
JyztEKkTpTsHs9RJcrCW0asjRvsjXKsW3KmkCzaFUhDVjUlpuJVbYFHgwZ4YY7WkYTKP9HcUS1LA
oBsUteB5v5riSnaY10BUy1wRGqjpit5Fyz/WUxK/CQjcwECRTcfNZEvbo1TK8NfsgXBPmdg1gpb0
z6+SSJ5BnNpyrJEDk9rIeZ2hSzVJ34SjL3jFpg0kZGNunba3AmkcTtEfHjatJSWBx/8DImoFvzks
/TDo59HiCYeKQKzB8XQlOeLY22wdRN1cLl8H8+DP/zizEQwd6Gol4WdNzYUStoQznyOiOhu3ccta
g2rlv1EMlL5MMMARUK0q6iQEl/l5V4ReMS/7rKb/2CsuFg8pm3MKp6Y9USu8KOl7+KajCT4FeOrc
K0vX6pWIguq7h3iZ/5fHHl30ZJSL7OplOpBPeWO9LzNWBipXQrs1dZl8mOBysR4AxWvb12jW2An6
OhWC9b6Mp6lo7XzkZukeTeOESL2dddHpFI6CYV9rqcSzIbi3kX6syb/eaw1Qk/S3kClsbcx9sY0X
IRDnX3r7b9emzp1p1vscFlmnYB/u5JWakvQFXpkuZmM7BrZf1IFTiAq4ypH2BWa4PRgfCzLXP2lA
xjcnWuaj/2dHdwjW7wnmYxVHiUtWSsdWSkGIP+DUXHowhH8fy5s/E2XaVZb0CEVGTLtFe5PfkfM2
UfQdxdYyIyDKla9Pdyda5A+67C+cmboMHT/3HqqBbkzMF19AGkbwuZchqR5Hd+mAHtScxSFWR7Md
FMYKKMb8Go850pBNSnYY8hwSYvKly20uYYBUY4K+rSt39oY7krFBNsBWe2/aei/DU8t1kkD4QeW+
inEvZPisryQh5wydY3hUT3/xrI3zMlstQE9GD7OeodnI0DKBEEIcrX0RELB4t/0BiyNF288xhM7i
g2cTXCH3etVwQnIcZ4ww/tX7iLcMZzVebFjO4O4mXrRzP36R8ft1DtMArkL2xwrqyRoVzZVvUPo3
pr+25JbxUbqWSbwnSEc1M/4XW/+AVVT1BCtE0aaGs3YLb65S8Ljk0Uj1zAaV08q7r4KOYkKzYuOE
MWZJ4uDqsfiBM76v07JQ8kwk3dCBvM+Jka2djZwheVNjxG7wSvqzI8TsHJsnR1mrqK6akCMNnN/m
lC4X65yxEvUzAxeChWIgLCNm0Fe+pSYkSPVjSXTtTX0/1/OpnSaOMT54T/YpqxFV91lDm4q3F0Yi
a7r/Dh9AZexEmatyEWUCmVTd6vU5CvZOH9/zbT4CexOCKZqSTHgPNtELv9rog3SxI0T1zc2Drn9p
zSGxxoKf1hLnP4orVd2YJ8D/7eMG+flxLcDhhEwtc1lxpjGHqpDgLCRL9I6TB6GsJ5UQ5wYrOYCq
DIBymzi2bg7ySL0EnwkaVTD/jPISxcmhIJMXr+fnjKvdwd1b49CBdV1RIGOX4fLviwL/tY4Dz9L2
icqTqxgqJBpPOVxkFmy6NpP7ZcLPPOTrk62xXS038Vhq3OG3rMh5qG71bPzFAu30no4TtPzbazk7
OY5+wOEuadEJw2ugnXQVJRgEhqGDDY8pyISsDHXT0z3QyAUiSP3gglJ9RB7T7Y2ub8zzN1E04TJH
h3M9xq01oEy6+EhmW+t5RfiERNsmAuWJGMFWylhOyZvQ7LQxVnqDiFOIsEKZK1sOBooa9nd2xdaw
b1oofToKDk8/PWszoT0Bsqu15WZ9qN1O+un+vZBjyWekRC0jIyRvJ5WzlptWhbwEeAj7TEVNpb2E
YOfRaWeuB/Zegz8vfF5dKypC5nTG7ACx8OgkaMzu+NI3w6ixYs8jkeFY5BZATRkq3hTpTd7/AdpQ
0bN1+Z7WyqWv+fnKSjzPwS8pShebn2TWW5Oe5N3c6xeA+9EdN3zq5l9Sdm5/kkGGp33Mb4AdclaB
pVomxIbDHKyIRPgSSsF80amdbxZvNQvF1S2GTh99hkTpIiRtCLDbGYcyYx8WpOga9xVtKEboA1ZD
cIdoQ/CE2qOJCaJN548fySXuPigR69X0C3/ToV3obrhWh718WbcqEZf/hy4pmCrnTNXaTJ78C+ak
hOtZl9KUEKklwcLaNhZopD4zheBS9Se8mlNO1NzJuoTwNRICG6ZbsZWm9O9PNFoL1AoE7gitqEHm
oC0V2ZL+jRYv2iHi4LGYSPWX+Z9N+1d7kP6RrqMRbQGSC7HLVIX+UiFzwsWti4UsG+VLAh1seYPQ
VlOwDZ95H3yHPKJoPTWQ2zQPS/+YuaIY0VaoCSAJowg194XHyhuw/JZoWqVOO16E7yNkwhScs0sk
XVQcK/Qb9NcZfTFaqx/xOcH5522WQHqGdBnjRX8vRYI9oBS6XkCG+lpno9V+v8Zhkq6YRvsrHiNW
myILyIK/9iFgBSps0bR1I/0FoJxtkv29HTE0+RS1KkuwLhnTdCrtfUP4zIRZZtI9A3URp1fRniEo
LtKqLAkuP30eww63MZ21UvnHsyJgQRwig8XW/GBetA19NZs8RzrGNPR+cRE+OlUkMlSOmnDtC3wT
XUkf8xKa2rWr2FUuJ6wISb1gz4iFQ5vOGg94Xfu4qONRHgjAKh0ttYMuIfcEOMoXGjDQ3TqRnBO0
gs8SxkQUo8JBGRheuy56v506k7zNkoZZzBqyem+2SSokXUsZ3wLfFtGoSg/0rcXZhcSIFyOUALcH
x5W8UqUFPusciD0luRyyRaWFUqoMPqYRIRrBTBDh0g1y0l21QLTWRo8Fi4S4q2mA5uy9LW3I3O/p
g3qrauyilmOk9nre8SpSTPzHbeeE5YilGFH1wvLL/8B6qD9hxj1hLx1mvQ/4r8cbrnDWGuGigP1F
Q+Ap/BExduYCpGq8VRxDn+Yf5sAazESuJenPOb/p6cmshKnTlOxmO1zvqejShKpRR7OcI/pbed0r
ppC2n4Rt/bm4XdrtN1oC0Uf1I4jsgNCVz9zbmSbWJV1+PR09SOxUMfXM3XFzH85maoN6k6bd/czb
fQlm/ntK9M/JNt2eFRsHbCfJM9Lj4Moy4uvLrHDx2dbVOHoIg8CXiefMLZnmbDhSqCezw/HuQoD1
qxNEe9VJFNNONLQdR3d0HDOZgrJezs4Q3CcNEQa1gtNX9W3HVOZ/RG6Zhj9U+XxFlKdx36x4zF+E
OnLw1aa1O9j4I5aLBPD5+yjAG9hj+nICPVHDV/S+kPpzL8Ru+G462Ac1ly2bsPYaGl2tXjcb7Wo6
KsWT4N2wd3RgtpJ+Si/IPTjFewsN8bKK4Bs0N19W25/CBR1nNVXDWgKdcc+VjL8lxePL0upkrKbu
SpdzdzzkR7Nxl2u8LeSLAe+vZLotzH/u7nrHjlZ7uyFlnItAUFCcGAPy1ViRdot7HpDPgqg2LsZJ
TQibFzluuLqyrRwjKOq2SCeJz4/wV6Y5D3+9M/9u0oEa8Ks4wl9fRGysdrf82MVdcuDzf2iVY7rU
GydkRvbHDgGeBy3c4wP9F3LLmcwGXPq4m9cKaMxNn5v1c4TCY7Q/XJ3tmIeDH8foDlOG6IH1oNf4
Q6nUBdHigW3puVZEqQ1+d7ThUtUEaXlokWJv6U7IFn5t8RIQDlfaci5ebXw5lIIYn7ODcyY6Yn/f
xDUhmJqT8HCmIqSZ/Q+qWAmunt7uXq/2k7cSNYIQLEiiXx7u3qBa+BHGiMKhxw6xBj//bO6Rg3gG
eN/H3hp9KA0Av/Pmkgxulrqs3E9djn8KG9jRZFh5eKg+/lXK1cULpFGx41+Lswa0TuJBTMhC0pGK
9urT1AlClFi2MgcHCYdwxW5MwSXGJlpuBg8J6sCjEwsstIYc/7t4kQIcuwAvh2z1GMjfwwkSW1UD
sa0zHL8ddEX2JOpORtRjKMEVAoe3mZZDT8Ar8iy5mIZBeOVwiZiqenS3SmYT034K8iafUhrf/UGV
8/Rp1/u/c10sNFHDP/b8QxFgg+X6JHWtgJUF5gD6llIe+A3JBmdgOjpiWX9bBDv+s7IydrqjQ0Tl
DJ7OTxO0Bd5a0XuMLpDAvZR5/7Di2zRWA3dhf7nqTP2y/MvkDdTGHcQEs6M9MdNod2aso3bzHaHf
c1lSlS407Hj2ajDE1oRxU/ghfeIHl0S53fyV/YGsrlT/SggAYSrOf8RGhpgbXCgwxfVLx7sE+p3u
vY9dg+M2zKDTsfQNFkDRofpFxt5Uemamu1wB7DQcmBt+Czn9aOn217Qjoc9SNiytcp2WgPweEE4Q
ZBZp2ZQT1Zu2UId6vBaIOKK2ScClsXgacBHV3Rk7WXkAiCvgkAtgwjQ1bwJ16yiF4P13teVh7vn7
gGGyN+iAzSQIO5au2K5ARKZJCKTZ7RKsUQNH25HWtw9OBaM3sigeFTfWdCqoiygb7hyrh6QK9TmR
8FMesgS6M/pyEZ8MEfDO4yYWo+cnoxkPadveS/eJMpShH+DYw96tYrzqkHL0RkvAWGN4cQyp/T/1
+xaZoSTaF35nOcgfZ4tS784ZWlWFvMTTXu6F/Am+dqf8pyG9DbEtowoyp0Wed+leosMbzhtpGaSe
3g0ngOSDSVnlANwSef69YhsUqUHmY6BM/k00xrdnFpwZLdbNlZLefnSSMOmhd/W+HI24FsdmptvP
zJjtdoCT9M3Yy7lRgNG75aDMOGNK+NaUYHQaM/KEUF8F+utFBsf5STfALl9GaH/PIQQ00Htg08wt
QVq0uHZ5MFLo/Vdqhj8uXzsA13deELRzMvtn5mLqfbgkODtGy++yEcsWwGjlKQG2RrgvO8sRDUCa
tz/axznDQuomT6D2usynPOS2ohX8T/yeVaBw7TGhSLizJQZA0tU3XkYsWznAuvAl9pnGLilyxfEA
eLidbSbqThbTKdfa4ny6ug3V556bxP19+uXb+5Z9GYg3Sxm3f7zV/TOOL68EHy1+3bI5mQXnKi/v
c/l0PIj7gT0i0HZWQ6ELsPWD81muRYm0wLKrnoiuLbZjQcucD/t+Dv2ecyD/1p9Qbh5j3/uzCvCD
fadMs0fwZZuNcfjjuPMhn5Q+T6J4ziPIbkRH0LUZFBOUc/YSBFEysFqabGHjJL6j0DtMha9sxtpm
jQDIAKGRG33nEq1xI5bWDK0FmvYKJDq9DoZNli0XOFoJr0/36LhZMEeVN+zs2HzMugtB59UgNBWC
DnOUn80OUJRLV5TKsImK6oq5UPAvLOr+hgH7F987M8Lt8bUdNnj2fxplEGGjrAtlaW80KTttOzQa
M4xcaxDp75HVjCZ1mnbvzZO+dHSiJ8NVa3tknNKQGRKOclS+LzEhFnlBh6C5JTuPZWyBZqi2KuyB
YOd1GCztcukVRXTYeRuesvrOzK+1NoFvuPz5Uxfh0TIcjEXUdNZ1P8gbwKM/XZ+XjripW15wbFdl
ogJJhj09/FqeTMXyQREIWlbn7BB1YGIN0C0hVJi+Z1bqezDpxDvLcDOFYe5IxAoBNvJShKaia2Ja
5vor40E6Qwnsl3b17Qj7G9c4qMFagJvo6hAgzWuTbQQvZXY1K31Q4mBdywuXr35j/Ken3LW36Y41
B49+trmwbmzgQapFPABLde3VR+a6WF7CFMDq4tgvjPi/hl/QF5jHxV+bf67a/mH/Zs37L9nWC/wu
0m7Cm8sFqxBdxj11WZRnzyBRIizqSmZd+Am637gDIf6vdaU3aM/Hnv/bbCeYcGuYSqQ7X0KbaA2R
IHY+papYwFBovcpqwGB3M9Q7YVbYIO91TCXmYiO5k6GixTkijCOnhPs2+V2cTxlABYAWV2nnH8CL
C6T3P/pE4wCpxe8uqqCmsp53bmZ5WR0cb/Ey02RHYKho8Xj/KwPXt7RUNVZvMRahMkjmKlYZsaKR
PEhqyooIOYWIbCP/hEhxg5sYM1Jyz8UGYg++pIyb4Vw+xojGw5pVNWUyvohkIbCAslFDhjjP89PE
kuFW3H3SuAtrFiP8D1LFUUQTOPrT4b3MLCUkGOaOGmDY7qR+dRWV5tPo/NA7WgIqLr5nI9QaHPC4
G7kvc5Lva85vIjqiggb/p98ag3VDARoezlJWOBGDG0xftUiSpeFCbgjQqXzjplskV8xvNjUzgj2w
mGutRSqWttP5CL6ZbS7pOQ5VrraAjC+DKYye73DTKMJ7aYH9dguywLG6lth+XwrAZENeSYpZ1h3X
ksSs5qDDLak/NrpnmdhYbcNcPLkYdXToC+hVUqWX6jA9fyBOGNo4KLYPCxaS6JZMeKcZnE5ls+kH
3Oba87WbJpPnw0DPF+Wrflr41BGCuecnz6gUN8oqfDhusgzhHx27XC/aQY/1uPhcWiWGQvlc6yfc
RUmAtB2EffBe6qiLrQiwEsAFsJo0gvh3RCvBIJXQhjbYlk95PzOs3AlidQ8nfUxWn79nkWth5pGS
cm0RSWxLwJooAvIJIul/FYgbM4tLw7yhLC6nyKbXm7ve7rd1uUEKmanGjLZ0xATuamOe8XWvjpHN
qls9ua8THZnM3I78k98eHYrVkvfFaxPBluQVooN+00IFDkWtP1VtFCGSYkhbD1Ew98nITNyXr5t7
IOXS8Dd14P/IyNn6yrGGeC6IOO0NdHw6BxWuyCFG8OJDk+9XbujUWIeHYgo9vU+5kUZASNf/Q7zt
IKvnDDLhMyG1NM/X8ySJPAfLNmZj6olS4sH/e9CK5JK6NOgGPqHueS5XaybZjVBKCvDWl8wavKcI
ODo54ChZl7TbmCBE8Vjxlq/zaRSjfKivKaiSvcJgVFty7WUppbilqv9sB+i51rzOr9dn0Ci6SkQD
g8BA7J9cuR5Vu5UkryTbAObqokAkFx4wEgusH9gFgKEFBeD/1kgKEy33ITyDswBwatHZy3Vbh22P
sLnLiaGClEfGS/9m4Xa2SkNJ+R8wu5hQ8MWl+1ttUp8T7+IZIBNw1/4DsyZipmD1BURCsCw/SyAz
StUrr19yeemLuFiwZ235MOsoIO9Sl4xFNSqc4tF0rNXyWpOlmNtJRsxlts0QM6sRFiuGznQSexJz
ETHhd0btm96NamnlmYOdmEOU4tm3mQcf7nNnNBchjNqCN1dnaY12sy5ULFvzc/r1pvcH7IdyZ3PL
ZLbLCejM3OHMMkpFbowNmtGW2kDCmQOMf//jL4A6B4VWBODxaP31iEVexWNDUiFps5VKvzNA1CVa
8TYWn7s32bIR3DBLsQDk8U8RRiOviS3lsL34HE3NeGhzRxZLmyVpfKtE0cZb11kSzjPzMgoG7HSt
j8JXUGCotdcySmm+t3oGIaMCFMvlMhiw2jicEUEqjOD6NOvadcj14rurUlIUzcKdZZuXJxR5N4rC
61dzRyoLil/6OUCS2SMwp+VtHoKxFGdw0gGwx1Paf52ZuR3mVW/lHH6vStw06/ddPObBaNvFrAbc
KUCbzJA4KkuEuhr7MosX+l69wyiTQ0KHYoEuXQqZJj2TGVOPUMskZnIxKYFmdvHgMZkTmYswwfiy
r7Wau09qycruro3EVBbY7nPrkL1YKV3mqmZHM776HdusYuUuNFgrPJ1Pzn1m3lGA8LENCs+x3FpA
SJSpLEUn890tIK4wP1Z2S6IJuxahWAdnCsmJZ6ycnQRz3Q8m/SVgJrIo+pmNpUcn0Dymxw61iIoZ
LKOKtTtgRZC9NsYKXWa6gU2wYFNKZ6jLmoixFOqYjyqHPijPNeRffa0IEpNGmQFy1KA/X6upfKqg
qDUETqOpqup5D2HRWmb4a4d9XtJ271PDxlJM43pVKaK93dGJ+M0WrseejCE+D/PmR4T5pF+HPbyh
gay53YokYc6DBp17lntJZ2kHTzOtwZufoQfYWtJJ0DwT+2I8690BoI+I6NLVRqlyIbg9ZKNT2EpZ
VhBCqNudVkX97+fdnXkGgm9OXXbJwofn1bd9sb45+63Ig7sPZegWrrYzvxEpAiibrgOD87nSyM3D
q0vUR7u1kNknOgCvp4Wmej9BPdLtJER2wyFk0AXV18qI9K2Wh8VUKQe5FcAVRbvAn8FDkju/Gn06
zU3zGEEJKJ7gljCWaZDsDZc6vm1ef8be7k5XzEcZfbRRk7EuiaeTX0b0YtMqZ1oaBWR1ELZCS9AX
uGryGelzlFpVNUWJkFt0/zPRqyd8OO2Qy4bb171BWBkLqavweGmUJ9SDjoo1i45w9nx5yEY2hCEm
5rB2lG6Ov0VAEExGpnF++4exxY/zal/HFwamzuQm/GoanA3NCIEdPjVg2uQzGEW+YQfx/Kbzz8L1
9r7b5djWwoHk3ZJm1hOii2EknhRQwU8dToOCuvkmQRlhXdiCiYRb6/QBc9Sceuoj+Ei0aXP9qFYI
Im/Eh9lTzie7XukD52iK76P+MA/aZ+ETqlL1vioVxzZang78ZdJG7AnO4xdNGpXtIl1Iwpn3S/Rp
saMnRWwMa28sWU04oxbByvdH/AEgAHP4XdmQtM0nHTk/0738hq63Ip3IdMNxsT/mlPtBxeG5jpc9
HNHrTjmwz6ZgutZbMk1o1XcEHjbfr9OJRAbAIQc/PIQnH8ZZ0OEv20I9RKXq8oXtmGEnp8l6IKSy
5iwI0ur2BIumlZYM8ae2ZNuIZe1EBGlSs443/X9URsxu28FxAtk6Ievm7pSPFqb5aYKpwx5lM9al
baQIAQmU2tpk0JRkVvZpradMSiI/HYM0U0u5kRo4Ydvwu9AkGVAqKKa5YnLR9R3utQej1T8mFXlX
9iCGTrgCb3SLai5hkxPTNj7107jArxfHCBVQv0gx0kBOpZhffguL1vOqihCgypMhKH7W0g9YQuGO
ASyy6HB8r6AxiVcBR8xx5m3I/EQPm93oCxO1sG7dZXQHjIINTsPKuEh1BE4cOmgXqclmJuCZIR6C
/6k+b83cCJhfvPI0IZQGacsbNqBfVbanDtKNbhCEZUEtHrvPr4RjfGLVvAv1SdP6a7qwrU4IErnc
IwCTfNDZd5KILJIZmP6Uaj8sqM6PKMZFrKzp7L6W+S8KgimhqeWC50DuUzrQeQfeaRHzrXDhTsCt
2jy8f2V1TDoam3yGPFTpRT/FgGM47k7Jr5+Xj2L1VZc6xC9ijR5Zo9zB/AgAEC36cAXtYcQ8sK4I
98EMXNkN2Ggc+hz4oPrjDIx1mGwghEAWl+6JrZy+rYvO7S1RqujewE84nYP87bPFgdEydhuOhwno
iZc4rNGtfKfxb7u/5e8e4JArPmNXHKLFpFBW3FOG/Pa9KT8Y3DkwBBu4cvgrMU/DLcmjqJhw4Vg4
7pr4LzRXcSdi24rH7Ptwe3vI8AjHhL+j1DTS4ONQGqhbuOFfFmN3W/tOI1kkqRDw2EVsNKSKpXKY
MUmIXwJWPeocapauIrHJnW9f2YoFZJTWtgNlk6AUeNBB1TG5VGUmAoQh+WGW0Nlwwbtn9pP2LvzS
qEQMz+Okincs3v3Zu/UGAju7XepLEMQck0JfU+GH2WEWszG8IfIlOzA1El8+ky1PkFImnM5Qf3qw
PX8R9vkL3I5PWcI2ntkPho9W0TUV5Mbe706nU6vWLNa7Ofwo3Q7JCxIgbP3GX7YRfZdAE46MXrXy
Df4xLwUUGHwPe9PdKimQxaIEUINGRA+ckY5vEKKKgMhOvkgdQcEM7PzgLiJwBgWGr7051OFJ75xR
7/FnMrV5g7O1f7UdLOOtz0STQDJHh7OCkkvau8sJkEnWvPoqh/mmF7CE9SMsM2DUmn63l8UPWsIA
ImANJNkTN2dNyBC/hwaGlWBZzODwz7CE4nqo8gOdezV9+6wa47gDrE0ub8cbu0x6QxSEJGnLelnz
dMBqAG2up9DhNwmp6j/O/LAn2AW+naDgShLk3s+2wH/SbXN+2QBN7Iwp0stI7XcLxjsmrCkDRCJO
We0PlG27NEV0tleq45wl0sV8UTSKIHd3QEvSRfRBo1n8dIqd5GUfksp4emITgr4lML1AIvpPR2HA
nlgWq0tCSRIR+8y5l9UaG/1FhgAtZ+XIDVV7QHQOvoWC1F0ib5rdfwy6g6MZfZn2/aLtvFV5Kyug
X22qURccX/p3ghQkOQ1d822C/qJZmpxCWzaK9yVZWMjdFVnFFYXwkeCnG3tF7ITMgLH1qvEgIhMc
ES3c6FJZoEPDVThvh2DygaAkpYgdLB5CZR+Pc6j4/q3/xlqtl9UrgKRdoH6mnGsKCsgXd3Kz9Z6a
NxjmnrU9orv5Ky8LKYW+W2lay4LE/bXs+9U3depHDQ3txGRHEkLWW+WozUXi3Hi5yqY9QGvPgpwH
Zl865tekAgsCwynVMbYFBMKi3anxR9ytSpkolv8dVF19HMMabxsAXBtkUm+X25Hfg36vTp5MUu+q
oMXnJHl3UETW5Q7d8NnTosv+yRwUQPmSc4Z4vtz+k7m1jODtyyoBBBdmZCQGu26y3SpX+3OFrVIF
Sn0S0fgxJT0A+RE6zhNqOX3N+Sd3g4MVAfu7uu/SI5uz4lGj99owZARA0UzFo06SNc4M4bgVwcZD
zFDHFF82P5rYOFxHCaycVA/MKfMfpTwwAS2BECjVAvxELBbLACpPkkaSW6jFSiquj4YnFBU1+DQA
9Ey3YTT+yM8hrwTgd4EVI43YhYIQk5mQiPlzNv6UwagzebtTLPojilgiRbgW24xB4/AUOvfjMes5
XY0s8SL1yJ4rNxbgTe/0dTOOCi+jRXTVK3AqhFnix0k5YVIGG0Ppo1yjF908Bzvj+00pwT6c1jhx
xofp4P6u7RLPpjytZK1KUacv5WZhlsdpUnbW0YYtwYnEQuPq77WjyVbaoKl2oKx+ITpGe+kmBXGi
gwaQDyXc8z5UVHVfs79bpW3yyQgDRvaWY9SWZcr48F/GCSbgfeNVG4RbTZdhKVtKilF7vYCOr4xh
Ag8a8gW4dNYWNeLg21bATgKbBPwlUbkm1F9DVdwDz4/1zMs2j9++vXa+VZ7PDqQoPXNDs5rNxYRI
r2tn638G9pz0/CG/L6hjiEYKJ6YnmwpAAZ9OIhIWlsWhCHoGliUV8UkPkrMR+nGVPYAicpKQS1Pj
w3bygl5p+RSxNE+zfNgV4LsGmCZg/n6REXPDLicijSePdaSjR222w2ohBuRqtU0bp13v7dCY/7ph
yM365wUdIcytK2NE27HyLnqR7pJ89p4NwVw7Tb5D7DheSsUGSp1lthzI204qhJu+skAWKnxdFtqT
xcR/tcdwb11UUJoSsGh97I0OTtAwJp0/hZLLmUw7PoLrzixlU5B/xw2x7N1s8ar3vIoSqK1F2Z56
VCIei27rZ4lKQu8Qzn75/ZUSOG8UaYPCDN4vS5sgd0xTutaDtPZgH67dp2GoGbJy81AJkt+c3fqg
dyFTWYjt2IQB61rV4OKnhmqWdWVUVPzaHEBKcix0fY+GsUqrXnsjDm9oXwKdOxe7+kFVAT3chCic
/Nc0HC5MqrMBdEt/15bX/Jjf1Qio8wNLrGb5GrYIEwxLt0Lpsux6n/LzNy37eVGlQhc9pyEfClOy
u/4BMJGfLIAIifOVmYsODL/CUWwh8kDSMcc868bLfZ0qpmHglfkelXAQc3WsYSfs6rnP0/W144Z7
7Ji5IjqJA6KOc8hYPoBQoS+VN7gnxnN0p/KJly7BCuVr0cZ3xTWpabxjeZPefsV0NIhHIAzvCD/k
sBcm2GepPAZLC3RGjf12/dH/gl8Vnq0GfcwKC2U/ZP3MGzerN3o9OJsgDOs3aE5psEuT2xJEpSCN
ss1Vo4+o9ccH0SkhM2fgkC2nIB/93zbBl1TmrSLQ/Vd7IRBiJ4AP04d+wmBPQCHzeP+ptcaO6mW2
Lk3T37jMR8fWK8yUUvX8mlYby+UhzKGpMl8KdMYjpJCBqsNyNuvo9ZMq0yGctApzIRLdoTiON7F7
PjwruOIZSvnpjhqeod4nOKs08MTvCeZZhKPGaDgZQEfUnGEumoJ/t0kVgt1MjOrIG8zezw8U4+d8
Kep0kUzd8FoNnbkEqr/Jq7dC2Z0/8RmGT6SB9KxvBcsy69j+31FhoWiMy/5o278wvshhOTozYTAq
rCl5vPKd3qLB4cWPfPJovho9wLMDlP6CwdlkDxGMo7Rnni29oQdy1wrJuKN0EfHj0FBFZaj4qeQT
fl747/NnQWiGpwTdd37ucI+JegSScDo/fLJ5aIGj6/NWVrm1DGO0+xFZ4SjjI5SyGyDiPwTjOaxo
f0A9X08vI9H0l0fmqECX5WId2HICRG8FDC9HuLY4CZbRsXJg23HhqRd8jSMASVuPWj2zvT3RwzfP
+AKqv9TVlv/Uksb20GQzc/ep2Xr8G2fGpApZYzX6vgCxjWxaCawlGEzK08i1Ivzw5USeHq/A1U3U
+qeOoqeQhUb4ZbKOYB9PXHgvUN08/dLtSMNNVOx3A7hdbOl3ovPuRyGROyoIbV2DWDo3CmxegBSQ
FggmDlwSGnfKGRIwSDEO035rTyIPuMBmm98K2Oi193qK8su5TBxDhI1VEHwhaCvOk0VheTcP2LnC
qokGnizEFrIdHhMRAtGBVcC3v/KaZ61e6PIS7RRkzKKIG1+j/E2HmCC9c3q4cv+Latb/1SDZ3fuP
cfyoIZf9RkUlXNfGN0MlMh4w1U0CIP7/8apflrvWImZ+Ubk/JTQGdOfyWnpndd/TlNumOGHI+xTs
6clgej42D+6TwGhYo2FjjZ6rLXZ5n+ByRkWNBg/uaN8EcEzdR4h1mEOXKjzA+GW3eD5PGJpFGerW
+YMMeSfc+jHxgkCe3QdnjFR+vp0DNWhUurLrosdLxH/HvFbQhqnML0eVizr2R92ft1Ofgudk5LD8
Pu+QAO6dmZ2gv1Ml9sTH507ht66bhfp1wLVDQq6zieic5JxuANjdKiRE2kF1kJgw7qnJaJYeQ0rS
e5DeDxfuNScbMnJFyQ2Bz4bkUs5mbEPEeOsw2ONGzsfGWS6SKk8ApDCTwX+Hooh6oypUWOPBoT7q
vpmx1ix3tAIQb7aP1IHVb1tqvsgx3bsWK6DS+N7Wkz5VrxYxbhBdl4NEnPSZ3cv0ZihPMRDUYuUw
bfnYptzIGpnAQSVtlw7u9irKP/sXZHYIHZOO3XEaU6CMgY3G4gEVbxH4KiXNLKaO15CsSL5w//OW
9tEbv5QTs1N+/+sjcuiSxbG+nrwht5P9RA1ZuDzuZNTnxCmeSxp0rV2zxLVoPJl4jNiX+MqOnb/p
jVCGj21HwjMPU7kIcZR/givG3GKlFTeD/vUC3qznOHMvnD6NRZfCpEX8OdECI6dpg17NYd5GWY1E
WUTSweay9okeeN94rZPZffLrbuldTlN0ZP4y9dcVDK5oryI+3p6FhmJ1j4SBnsmPxrzdT/XQBUHw
gHp8W3GD/g4XAmXu1pJlazE/cKaG7A7gKdP01Ls8iHn7Fst2xtsWdnlTeWWNjUYgyU3hK8/A7mge
kUDaLiqdeAFtbGU0LRdKiFwDKKtgjSjan2PiZU6x5jGtOu3KI+vym1xrteaO7Ict90eSvWPspukL
lrENF6NBBZm3XdTducexw/5tlliyIAWK+4VRVwwc4fnCF8GwD5yxQXDXTYjSBz2m9r0A08klyKuX
LQgWMiMW3tHskbct5mLHegxGa55uEfG5FcvqsDU/9Kd+tg3wHEm7CW2gGNi0lbJCq88WLarVeXCm
IwNbvlgd3FqpMF2W142ikpI3/mQenMHc2S2adLu8G58sXL65Xi7zm/iqiP8deyCTKolh2/Wj/RdN
j75inpeXAvphIrckulfC1OnhYPXqEzVmm0M44QHw3giOpxoYaZ0t+FF+N4CX5gLCvC+CeQmPaN3Y
00VjNAwUJ8QV4i2zPCSOFMvCxBuqtNASJAdg98Ib82KSQAhyGSa3Z0uUp08YAOX79SDH9ICit3Pr
RXNV8XkZ43nNa9vgSWOH4mNHXIpBWPbcotEPd+uDRVkX1jx8HV2qBL5kQuIxtAqyGG/UxT+StjSV
KCbd/AZFKFi+/T/6ozcrkY1X47nO8wZpdo+P7Pva94iunZDAf2gDd4WUyTka/ACw2er0aCtoozAE
Ur5L0kdFl990AsiRUxrZHVEMwsNG+a5ABW6EOfolO1lbfgLQ9OPJ8jZNlZ+8qgLMhR4r/NDp0Au4
byQyNP4TEtVCgo2AG4zlBJFoqdEUg5Jq/i8wEWDF3JNtjaQdrz1JU1sojmPQokTTcmRqjdggFfiA
c/l6L0rbVlDrAKf0oVPISnPUV2pZ9T/xleMVnHI+vZpr2344HPyEE6Y4dXoR7T/FMCh0rUNKAACf
X73zBBNNdK/Gwc9V0IdRcZlNqtbtMWpSGoVpmWLH4ydboS4m/tggqqCl16pUon96bkVfrIXXpKJ+
62ajuEMPpZUkF1Zj4t+JITOI/lr9zruPhcR/1zUC9RKhVFcrBNjUtwifMmrdOBMPLrtt4xZFttrg
q2FpKxmawlMm1U2lzBc6U2jJYmXpJRVnoYOQNMq9Xa92SzJySLsYE/zNzSkIgq9T58XGj+KCWIA+
dX/ZyFlxUjCafsgxaedZm9kMElfxTl2CXv8AeCFjqxd/ROw3mo0o5kEk00ukhZl3vQ8uTdjptVyG
t0Sk2wECxfGFMR6OqtcMIXfrpzQrf5GgROIC1UPlTzwY0nQxjlWuGaM/7Q+EplEWlTggB1YYRrFL
dTw5II9DW9qHKkLKxzkk4Q+eoj+bI4YRRolTGdeKkrrazCDIme4ekZ3csC9zmCa7RNN0lky4cHZ5
94jdYrNqqgbarOnZPvImBecqyACnHwOvN9U403JhjBIyDdiSI/Tc0TOm0dz2AaDqB31ozqaPsZ0Z
0f5C/Hk/TRpZF6G6KKHoQcx87tmAdxcsgb6fuJ8H1vEesgdDh1VexvIr3TvnxfHJvjXnyb1gD+5S
TUNyoRcAKojdjSasnBMwLz8sCzjeRDy0assC6qEJg7s58wNJtPAKW0WO84rVPSjZPxwHwlGs7r0I
8i7GJUZykZh2Da5Liyyk1eOzQT5v9Rz/ZUGgYWqkurkZ1wTJ25sbv7mSdQp6daQAauSG4vjvKkES
U/pSeQ8cgIBWrCPpDFMVjP2whyr3TJS2B5MTbZUsB9U3mDD3khfOWi1wdpOR4+FZis13B2EeoRKX
0EufpDeYT7sniJTmR08kKP4LP/kdbQ5VWLbXZ9Sx7zOy/Jg7b+5OoXPrqHrW+gmrKPhXHhcuThW/
M6EbaE8PUj8JlboxTP2DVOstOvKohkaigJ5vAq129Kh0z7CHBr+Bb0LWr7SgyFF5g/3tDbXbLnPU
YFtUVQjC0WoBQ5nE1hMmyBF1PsL84YHKyKuzDfxUjCG9RKRWdnR5Gv+fbzpOldDixVMe6IKDXSP9
W+G3oLhsCSE/Yic8GaK1VaEP8JDABO+ffs5tDP/sDeQlBkkptlXKegsIHdO6ktxL+Ei9N+8s+jCc
CYmD0JtHmSe3Ff/a6e08dVPhLuhwkC4sHEgq9IuC8z9uCIJw6/oFcCpKd5EgQNOB0gdQzn6VRcIa
4do4OZGY5k5HYTjpoxHMnwP9FUc4Yq9fnu4TDoURqT74T20yJHMs7ojMhUnIK6jaQDJGH++9ACIl
tOQY8+Ec1lfbYtzCgm4yiufZWgYb2ZTkLdgyNVWrXIgoP5DdvcXr1qwjrV7FpTOafXXEpEk+YZk4
dvh6rlpKGtOso8fQyEQBfiwH3/KPSJs2JUSAjtFtE9HzpqU9OicBCZqCXZ/F6hKXzVCo/tTsTxwJ
tBBk/a4JxGjggkmPUHCqpmg0Nuznt+rwXhIEK0XW+AULRHG7+sMMP3MY7fvG+laNWkxNSVJSGKuI
XUWbGFKXBtQJC6lU8uw9vz1pSCqlgQSvuwOcqKYlZDBZpP9F6zh2DHQhvcJqnxLug79EnH82jIIv
fHV6UQRzBFtjA8xQhCOM0zG5le114b3VlrAyt3Nqv1/F9RUHDdctnlMWUCbUzuaIx3d7vZpEExQZ
a1yAMSTyBLtgzvOERTbYhb16N5shMF+uKleZk64Wp0Kx0kSiuPHuh833ygtO1AcyT/DgD6yFGlZu
n+LLmY9UniiIBKvQcqs7A06ApmIKq4Xc+BrfLamxH1BhoHefqP8OaDfndRVFpZ66aWBWChxacA9g
dEJOSod702yU/E5OkJ2qWynIuQ+pjtP2O1MRe6Qro1/2vJcC5k7kM3xx2atCl7eeNWoap7ctiaIb
hHU0oRH6N8c2AGL+YlD48TdfdhZ9eIR5K5y0uxBITQTT/Wyg6tyH9DnYMzuY0a7KyoojpaPlaNn4
/Ju7l4EuK0R5+mSxRhnnH3pbB3DKL8H1Oijgg+Ge+PN54azqms+TaHp0lQsomrDGg/trylTG5FGN
9chzLALpMcEgv7Q9gcuRv81XDoUjhRwPwDQLA3YKzFVQ9QeoxTPwDCVIvvT0UUDQ52W/Whh6QvuH
sv6wY6SkoziZ/BxJHCzN8bS0vEVG3zkTp6azpVjixiACaSHghBv7kk7cYbr4B9lp5nt60U+rbGno
BEKPASWKaTlKwmJhYl8ELGcDdbFcsPuMpBxYjxtXkW9e+tCZiRJC26KxQLp1+w23lIbYzxolDc9V
gy0oH9ruEnby/rCC7Dg+7AYDxyLAxJylQ7zwE3zVZzkIR3vt9dd7Ox2qwyy+5Biogy3kOOiqj+Ro
7rIX1v2eYCfSIwPcPbR1CfG3uIM6r6B22x4f/GeXPB9XB2bA4lE3R2EgMadZQilAUsX0RmyhMhYP
aVV3R/z3SeHe2mtgB7R7wUz6SdBF+P5hWD5gby4VENg9DKxHxWigmH+7LBzQeuu6M7+KnsSLiy6Q
riQDjW5KyUBRqtptp6xbF94+bTsb/hQ67xUB9np/SkxxFbtyvhCVYWPyX3VTxRd1M3+gP4cghaZT
xbHiz+6toNmrfHHKv5oizqv1L9CfaTTZBECKBk5+RLBdZfvhXb/kDmnAz2jiGF1mrrWU3apySTbF
8i3lTrYCuNXh7K9IfKvNP9ihhODQaooaDBq8ADCS3MKCZ9ntCuHrLlovcU8jYSmBoi4gzJIv54Vs
vghYA5F7lnWu4j6CkCxj3srqR+YRR1jI1OXQs/SZcECiQgCO7ARf9tctfn9ohS2VuCFQF1kJFOBi
3TScqMwlIPiV7lybSgDd0Kzau/oZyVRCFsefu+/CGoLAEqeVJdRULViJelqrt2dLeuig91A5dUjw
H0YTN4/hy6TNuI+hb3F6UG2AbZgyG8xoCT/B3YeZfu6idoDh+RLH+yIn2TFFxHZ8tZj53bV4mvpz
m00ds2UwpKYafOVWRpFRXQOJwBxPeyegySW8nl5PhcuMO3n5Cpo8HfpqzsCatNfDwhZp9sMu0Oy0
mVoiGTNSoKWs/OC9P+hDIbfDb0TQtdj5EFMEzXfwV9Pv0oFvG0p+0rr3R9xa3rrmhuJL4D9srNgO
DBzGcq8KM81gxGbKK9F4E+Cr8NKWKd6Vv5w0Cs657b7w6dV8ByvlOpoI1pwJO/YcimkwqMOQPNF/
rOJZSCUP9/IcGSnylWEHYwSKVnC6MBUJ98tcY5h013D6GNGwRS+65ecZkJ9CFKZhX1Wm7TSdAlp/
QkFSJMxo0KOFk2dytlNz3MQK0xubd3qJzUP8zPSIFzC+c1Ln4exLttUdz4yMWDxwG7pWX1ZmXd+1
kjgreQ2vDuoVEPQfwIhUahOQXiuvf13QxhzxsjUhpyVP9Y94WZrt4dMbU4hUBVBd6uZz2a2Ofdrn
wwSUqkPLV42dKxCwmuJn37uedGV0QQnIMDh3nLu5dPRWtlWaWfnYzbxcDxkB/24YNKk+Nn0c3maT
vk5O8/gy9psioo0I6Yqwh1YdkbS4YmK/9WnHHvWbQrVLxpI8uk6+LtjCQ6csXFi339F7Hz08uy9i
w9xu3TzfN+lSFV8ais0ABIRpUeXp7/NF4J9P2gzxItSM/ngKbAFHtafaafp00fj/zR+ao+yHGlWT
Y3+we0vsQ8Iq5Wby+v0aiODAaZS0+xL0zngxKQEc+itLRPij7i5k4el1vO4Vq6N3RBbKugONaERC
7i7YIdpydXiYPCxFCizEqGgUnLaYcDlSw4NhDGPLatcQY8yT0b2FI8dd4IXLLSbC3l0JeBd4A3V3
QMPDco1ENT1TkpyTDJurO094mIcdqnPFXH1Ie1OIR2kQAgR1wSwcGcGxUEXgm/P+ZEzP6KVZ46mu
kksjcKjerRjSCjYiee0zqfyfmVJ05fKA0nE2tKgSv369Haxvp0Ba3tVEa+5A6PY4wvO5tGSLKOjK
CLIwK0ildQRHre0gUBi2jYZz1XUDzkqJcU9s+4WODTtS5J8vQgh5EpTWrpxlVX3sP1aXkmcPBeeM
rGe3GOwl0cy+cDDKWN6LbTaIyXC6MXUqIUtBQu2fFa7riVnN901+dWYa6au428DgAFASd89/4brb
pI9DsCTGZY24bWhf1JuY7bh+vXdzmYsw/RNOkL1NQaP67YEGHMoQuDNwiIUvt2RA/RSvfHjuTcKo
LBm1p/dcbQHWfYsZGDYgBCVKhLS9CjnC2o98cL5Ol423sv/fod3uOfBu08I0SPU+XIqaN5yQLgef
DBViZxeER30fFCDkKBD9KZrWi+NIdwgSBWcyvRE9c3hHP0v9Pvzu4slMlDJN9L6gCTwfnldMZu5F
Svn5ve+Ji2XVDsdrDFNrGl6Enz38NFT+URhB82TusbPjqQ/xx8FGyS2fjB2PTLeFZMNv0TRMBUye
USNXQfuBCcFwOV/VOJGeACmZxQKPqRmpbPnk44AX1LYzdTwh3A05qVTjw3W+Lhi2l9uaa3f0ES4m
7V+ZVo4kUVY6/6hhwPjpSjf981VgClk42/COwqn9Tatj5CxYDghoqMn80euVFOn7kRRm4IkkoCrX
IbvqDlS7nkCN6J1qqqpv6BxuSw8t5ukCzlAafT/Gq4ejOBoNNpCcj/pmwJJMlym4wV+WveHCn3Ou
xOQQCbmWI1XUt2nUrt55UU+NIlC9b8GceqdhOHrrUpqbsHOT+L6nBrhZGuDoFQTJSVr1jUOd445K
PaeLXWSxBL1cTmGK/UACxAKS4VwXFP8broghjAroAjGqxTR4EQBvk203ZLQ3JdzjfQUPCCuHlZ7S
7OVh3KS6X6nIUh0+sz7ZF9WW2OcHQQnUz5VMEpN1XjW8NI0fNFdJR3qIb9k31khMJ/6TZcIVRvVS
lAPIrMk7zj+cAxCl9gpeTRkKAdgYUmaHcAPSoAaa1ekpf6FTuyNenuoR7F0FVw0jGwY6BjfRXPl6
IRVvSGW8KF0nXN7bt0UOBSxb0C/5jR8U53S1H2VcHMcraaK3gvyNPeZw9YQDOxxGwMvOjHigxpPG
Y38Ks1Rz2IaO4AyWCYIwr/GuEl3u6MHCTtaW+8ZQnVhso2tUlZ//s/u4YOwMRxr+j7dDVXRO0Jm4
YoFOrDFANOxqmwBj6mGOQJGxFN56W0ejgz7eVcXl21VAhS1b4DN4FlglxGRYCa6PpGKLR44X45gD
Zf5SSSvbz6HS1fGPUP6d1Q6MHjct9MCre+qk9NPaw+Mju9Bba/gqEqXaT0/Vyvg/l2rDjWK26pnS
b2S0fkU2Th+dm23v1CRCkASTduKBtMtJXZM1+JrC1c+hEppljnVRoHqeEB9VKD2dcz/o5hA69/QG
9DBGQJZ5r7/XlTrUE5nn4J39hOKe8U7IdjJ+PUDFi4kbDXuTL7cw/QZD1OluVrNUzkynrkNMgvHW
pbggrad8N1u0Jx/29+l/k6LdMcswSVwoZHr/L+BcgBC31+7AnSyfl4fNVJ7GDDYxG0qeYJtPmomy
TVW+Cq0hdViGAYLQKoTXeyqNprcT4T9Ut8ejtwj6a3aGtmQKae3JiznJYMs8DIJXGdN4dRw5Ozdl
wYeoDtqC2Z7ha2iH09q0jObWfdHAtWmT0NLk2Ck1suW44dh1ncbycBmJaFeHR2DljfFq0OQKEN9u
nnoV2Wa65wWA/hlT/7/kn4GKHG912AP20oeP6cicfbQS2S0pWum1iLkxH0Z0RtG3nluhJ7ZbJ+hL
O3A72sr6uLTQeBUTZ+UHyEGUug//8LZ6TetzpQIiUQ79h0ahN2RDDw0HAfOh5ZoYofGI8Rqf8XIa
IjyYsPAUWHGeMrvS0VnN8awbP0vGabYXYXDYO9ie6g3HaM42FBUX2YnLQM2r3yMBbLt8xYnfSeF4
/hWNmsBec7zmPeCTF44rNJyqcRF5HYjpj/74xNZQkJO6fc499XGbY7ufuR3VzwcsiPexdtw7J2gP
SaTFw85DxEpCEHGPkbjGFHSdRY+YB4YWPN2/oOj0PPhN0z6MPrDnvTPtwvOXL0PAvjMRSDtyvetN
Q0VeAq8m+XUv9P6IbA9CpVeGKUpBzOY6C7zjTJ6OEkmfKJKOwJnieP03+4fukZFiDkkqw1AxQBXQ
cpx5RsmA7X1PuvQrsJaIUQ5SP1UJ7GRskE/mzpdFX+HGlKUG86mt98DZcF6RCVGaIxs1/kiedE4T
dwGyeYL6QN6nHTkwmV7ifvbFay9roN2vi1hSRR9xaQocOrIIfuQkuUNXrfvrFA3H+TVQKEkQvZQz
rYfA245y49HX86apx01z8TUmZ2f+KJ7lvKKYJ9OffNM925V6JgT6nfAbH2MdDran4PBM0k51mHrr
CKth6epsV2jvcM9A0Yx6fHcq5X5nHf6fmEUvFZJzWuSveXw7axb1ihi5znOJft8OHEjuh/cRdSCs
38GNR4rS+iaCNRoLtnCW9Vl3/9m9UBKRPJHUhHcQpU5tRF4dA5AiEcDiLLu7WjAU1D+EOzbF4/fU
PrH9YiELg1JBSbqZaL05k9P6K2icnxDzbybHMJpk5YxdrQ+kKYRFuKvTYZj5drcsfj07znzsJ15f
yIxdXPDvikoQELbjKGaxU5JWdMeIsSHV/Lp0mwi6o6IH8H9NRSnO3fnfBp2ocGuh+5YxsINJQ9qa
uTwXRtsQixTyAkSQzbE+Gipj8zZv9NFBupbM5wU8VJlpAf6MKZsV7DPd97bgdPqDlX33BE0Vz8BX
RM4WNIAGRHqas5yfka6vK95iV1DWuXu/lkereaQkAgdIlvFjUYz9thybDcw9RWYB1IzdZRnQfNi4
vphzRJ+vxxAJTwD7HwCHRFK9LE7dzo1XzcZYSKTOCy6quuDErNjVXJRO5p4k+kRO9yhbKdlwNLGQ
saIBhBF1Nt7srNZV77ytn1BzC4NWOMFwSNnAqv4dFwumfzjR96C8H4oS2LqtQRhlRGZ95OBNrW3Q
8jkKlfIdpE4aQ7TA33HdWax4DLz216iwRiVn1s//VF0N+OTGTTRxo0V2qs4iA9ehW6brqBdmD6ni
nCUhsJFAXsuptfS0aWtMiXXMj/8pi/gysduCyV7CgsoBE5385JrTEhMLkMqUU18YM+Cr6WhyVHDv
zmNPz77Kvqc+xGqeca0mo/aF8QIouX8UZXjnSK2R/xERA6eaioXZfiPQl9HYNvQfQiLfEFiZd+jS
6fxubYa4OlGcZ4r3jCcEh7we5SLwnEtIchDwSiGL9NJvCDGwpabyzr4QSXqcdGQr89aP+mZsJKbq
FQCfGnHJcFUFjYr28VPbCHo3aKvfOqytn0TpBCIIBfDsAJsx04UD3ogqqgOmXHkC/pYXdcsODBGv
Csp2mGtrR8ei3zxy1GVexIWjUyWRMNx/R3FOIzKCvQ3swufHoYn6AOhOikfwRwloh4PkItq0JbZN
XRnSRQe8M0INu4nHuldtuzoqDsaIg+asObHfox7een+f+UKTMX7ogH1CAd8QYDWC0F3GrV0T6U91
xKdi97o2MLiWibabdR/wYhjFXZPNVje+zfVh/IqeV4Qf58o1dJOYKXSPcVIbxmk0BVrWWYmrM8OD
5H6bdsJ9+Jb1Ic2uz/epSbm/6pXXi+ylAPPoa+48p64sa8AVQMIJeCgPnPRTtioiyiPfGriKtJ+V
Cn7uyTSxdT5meEXF63sKiRSQpAxgejt486NstA0QuCsddR85oxmFaRdGWTwNSghIvqVUZ94FN8Fc
5yigIsgYBt/iDfFa05ZLy9boqgH4QkKJ3mj7lS3ZH2X0XWzXS/DzV9pHOChp8L41w1cCU16GrqLr
Ah1vSIMfhNmWDCNbQVs6dHaAnFN4QNiVi8mYJeaMTtOjXGcb8llFXa318yf4bZviVYaKK52gUxVD
mDvzX7L+QIahQUjxnDnK9C/YQgCipP487PtOAkrm9+rLfM6UvualJLEZMFR3QRapslfBqbXqYDaf
DfRqd/qXx49jQ6WWQdO+NkuAFHC+oJ9flX/eQ/d0VY4WMXR2no3W5KLZK+U2tdpFn0VkjjLwukKV
Jr0LcVIn1gZ8y2vX2k1X0J1C0Nr+AJe0Ti3iyr89Yy8HrtEPJGZyI9vGuaBlNNXWSWvhdXupD4gA
92aFs69KueNiQVhjnjNe9XK5uPfuYEOxqoDAr6D/D9gGBkK5+S4yM5hWNIqgBRft+mc9Zdr6OC40
1o7WnRl2ZsFVFKPWHu6xBR5ueZThdPLqjb84I7ObXkvXbMEkHztkGDIHRWck0rFDJaPvWZ8xnWCC
TC0WY6KtCpOU+nhVLURlkIF5TTUbOLb8P1eEnzBBe2Vi5G63yU8QVPJB0VRJk2pj+WVjjAVJJr0V
xD+ESYrVfGyDf73MPvNKg3Bq3PCht4sjIJWtX7X2LKGCcgGAqOCW3A/xSZm5MFUohHua5zqZzk1y
yca41NcWgLH5IB8Un2zN8wndeFr/WGIjqreoRuWRwLkXYZzpQClvtnI/BZQFbvy32rnWpCDV64/o
ArRkjFBpkwJjn/5jOkLcbEif0SI8QGhvB1l4zCbSVx4mCWBUD1Pc7yca/idu57VycDagC/F5k7RV
i1iT+ra/d5F+Q2+znG74pL8B/ZM4GsIaub7PMF2c+ByPPwZibR3Yxnlks3BXrPw0yaOSdv70SbtK
mjYEf0FGL9YBUk0WXo7lN6SziD/FflTUdrRjMxWQgJCOfdovA1rsqRANxIvUgM16pyGj0A/KXyAA
wP6P+1FYuLmcA16tV7Fqwj7YRxm3ih8jhWGfHeFkrrrM7GE1tokGwg0o0QcQXpzLiKJkfjMXI+4U
p4pJjTdi7NDNNv132HpTYp9/t7qKaryuDF1CKnGCEYSrfTpwDLOVquhX/YB52qvygBAVFjieTRKF
NDnJgUd04ro9fQ5+qSEOWAmTDX23KC7UX+rETtFIGbNZVaEqtius5mnb1HsgyVdojBpaHdq2IY06
Tnk2w+AEW9fEyruR8RYlO9x2lzFxK5Ih+7QUd0GQjhUMoUNB918ukKq72aEmX3JQnf6FLMygF3rk
2BFqyfs0FJo5kLST9OMP1gTS1cqUod9Yr+XDa9OybgPEvQMQF8wOTCTLCloBZsDKC9U97vQU+bZ+
YHT51ygg6P//QY+MTyucxAuZMjySWqaDE+dGlAXiZzdVBwZJ2peBc2azCtVgK4Wj8GtksskaqZ05
erPIxGkiE+ztZl5Lac4p4bHx/2gm8sPbvjfR66KKySBVtUlPBnoc853w0DwgUO6rBFq6MhGYpAvM
SpnTEkijJH8jNMdOa+I34afYSIiK8wYBVSnpLNwFKMvPTnlLo8CMjmENLIZl8ny3EnnwF16ZtYHr
JOWu5MtJzf3CDYbjA3VVn+ZKrIEbllc9oNUl63pzboxPuH8fr02pCRnOfVjaAKkumxeMpMj1fSD0
72oOcconjxa6zSyqKZJBAprNLX5SeiTRB0g0fmU6ZN/sp7SvzXpCM8Tp8HMm1La9cxk3i/OfXBmQ
b0MadVIwVO74jRFjnpqUIl+RWYcqbDTMYbqF5bn0BZwALLQNp8TSPWwNg/SC056uUfw6an2fgszX
cVWnoG1E1GpDQwT9EkTOwSjbBLma98daFUFfsuOlzc+X2kbxc8msw0S8jXPtdnS/fSoIuX2o5Y9v
dbx2Npi4uTW65sG/uwbFcSfc19kqH50ONoe3fANBMsBKDR3Y5g8KrZCg6BgYYFTlp2tWqiK7Sqtd
W8LsmSM7va0xQt/SEJMWlvPGOgm9ap4HWzDu6BJ6p9+pA9MyaX7XrjGKIyxvBO7wJ9a/Sb7jTQgX
geqFT0D45slD+QMUKxp/7BcaE/AmJyPgJosV95bPlugZkHDGP6ehI+6ttCR44Qgz7qV6xVoJfuly
bylDlBYP7zaxW3HzHQ9QwL9rNvUAx2kSXlF1T3eM6p2i0OjFU9pYpO/KmlgXlAf0bKHWXEHIUANh
N9uUVC2wW9KwTnxXL0N5hs5ZahmjQdMUW3GEaSeVgJXXSbZ6ATtf17AJ99gRbsIenCBzyr8quMDP
NBYKw1eiBFVkdB3pKiw0oHXrbAl01Tru8ug2mOUfBM5OvPjdrIMrJfpeX4HwePxEqmT+kZPLMTYb
QFWRoWFqFavWc3f2CHGD4hFzvNj8nzeX2+ijn1rODsGydnoqI28C2ykoOcdCjjFLpS3yuCfBUiUf
FKasnciqKP5VNHAlvpaT4DoGF/I7Y9t0aFfnBx+pPCeSH9VunMzbIOXeFDNz68YZPOWhcOsvVdOv
f01nLMvf/rla7/kufJlgxEs+QYMgKLd5akQb8QModXb4El5smpKEQk5mEUJpwgdaC6Id6DwNABpz
zbW5ujJRpdB7RFzVneaY1RmY4KT3Vu6rdG8OEhLOTREjqGkKFT/5LGIopXH01VWS52J2Dwyxs9Q8
L9tXrJf2WkK8ViO95zn31WlyELP7bODW+lzqmxAhX5ZqjRaykS4YNUYnCcxFijhnq8swkcCDwq+g
U/kyR0r2PUvzgrPxIjf1ONstC4RCCmSee2WqUPOMef77ITxAevDzbAX80WY9epTeeBDw9oilWY/F
JN4AG15Ou71/vu0cvIkRQU9QUFf1xHy9kfkoSbKfYNrR2kaz4cLHkP4ZqJZbAKekAW14CH9xixwz
ZUZBY9kIrdYQjEx1krHmiTqwg+BXazrBiSHDLkIql13/QMJJQC8Cbkn//Dy4FKzN2ShwoZfQaeZc
+F00N1qzgWerij0h7Q/LunBvDc7DdmDt0a6OnQrcfuG+MqsV1mG3eWdNfp+IbLpal8jAr0zyXk+3
dV1wP7BKmK4pWzG45mt+36fIeW16Kg1L94syQL4RhHiSK7VFtQscMPziJE0dmcj6yGQUY4h5F0i3
ZcsMAEt0W5Wwv/l3ZKVxq1IwfwWf0wnt37EvTOaXGeUvJdLuiVzmEzMS56qgrQJrETHlwDfU72/Q
mOgU/9BkykjGEOJUAhhu0xQzMWev2cZSeN/3c9iPJeTzpAbccDs7vBjbA+CVY7qNWbmnFQezOMB+
wj4Q81oq4l4WzMUWbwgmkj4Iy/R4T5lpOUo/uPKei4MmHyFUXV3g0lVYH0enKeJSB242FTpWrNm1
oD16d08+OZzY+QAOXHXPCjgnwo+ZekklOpOS4EMxuFG4Gsw4D9BLkE1I7GQtdGQQ8PNtnhj2q45o
+WVI3CyinDHCl0qGW1BtCFmI4bzt7rNasrBO0bswMEB1teD6fd8KgQcEgBobWn1HbO0IotINVOQ8
15JlauGDEMpQnZ/GAouTu/niaAea5nYxzv8rMzrPR7B4A2NKTIkr2VCm595KFgynW1BAlp2MHrDE
po3hs4Lqk2/j/3LcWthoCtOc6c6lGhfYYgSPXUXOvHP9bjM5b1oKwo6/uWR5LdSDtWOSfilH9irG
IeYlagzWGICD+ErGUlRjo3K4GbmYAVedajK/UVUUppMBrlLsgseyr6N5i0WvwpVs60z+GFafgd6u
XnLcVW0cNX8EscY9YhKMPmF5wjy/Psp8KnqDxYyVfC/cYMqjWixzaFje101My7M/QbvFbN4nYiwb
Xecqyl/EqeAnKW3ISAEy70CXifh+JjeMgFqucIY/RoyRt8vgKSu9EhtVckzVNGm79IST9W6K9SEl
nNfRAfROT046uQYpq6BNYGs/J42G+dj4OpEkPlda34r05SCsecLvsAbHbdSULGq9uyKRubVZG7Et
8uIG92poTbYZZitGjkSuS5dlDeoVOw2i9FvBPyPqTBDs4PgTpgEpfIE53YXoPEuKun+vxmS/6hRs
JNWkuH8Z3ewuZVrwum9lcwH92EZ922i0cxmoiCkz1AVRuIqoFdDTNoFv+l9h9YzKfXEFutUYd7cf
qcbW05U/LrOLnr8sNA13xiAsGiUTR3fpR4G34cNDfey7CB0Nm2VcX3qg4W8qrRIVhNBMNjIQgVU3
xxfo7gi72EwUxxHNUNYWYsu64Ty0cSIT5q6rwJ18uaUh7WMyxO7QALYai9AoXtGFxb0O3mzkgxv3
JLH/L/jBBOQLegKxFC++Khx040wrd5n6OMMmrzXKSZ3ULeiafmDCOtUnj1lQg/GWOD6MDEe4YfDw
QgJ+XC/6W1zLxwwSzi6XbYy5RZ8QUWt+jrAE1EJJLnEFI/zbKBvwfNXSewhXqEOK1tug+WAleaFM
pFIFZ6lkgQUMQRxXOzqNiwlX5BGrbNIQaNjiY6NJ/4YVOomRyXXjD55iFeds6zG43I3lcTYsG6F1
xaGFU0Nn58ft0s6mBL22bR05+l0R/vQ6rw0ei43gqXIKQkU2EMwBhm/ANLtUGTQc4tGNOhl+84Xs
sTG1MhTV7d1BUIRupuaw4/v9jpRIoVozpG1ciwMMcbo4/PS5Bfclv8IIp/u8LWbisFSnW4Husyds
IxNPa5dpgYbYWXh+X4ATf/EI0OAQLqrKVU2NiNGh4866xEbTaXWmdzNUESrbyszegw2Qq6kY8WHj
u3NMVnUsxNBH2ck5kOyKmtUmg9W0ymemjQTjlnUzM5MB8OmNRvS/0D9yudQ1lzsJwSdRF9SKZRRs
ad8dgmBESMbYvzcbhOHlJjH0CyTIOAh3rdW0y9BxNLnBxyCL7Gybc7+OfVHtuh9FXpk9Zg4hSee7
Gi3WkQXeFzSKqo5I7sBUUV86WM2CzH2Z+VpJM0BonjBXMf0cH0+ScwdrFWEibQKVaS33/nhdrwKp
yQmdPbTyHyfVctN8GLwx+YDev3LvXsd2yepJ/uXYwdHhr/Xq3IhvlzO/rZoReOu8UDy9FeJZWhpF
e0S1q4wY99OvNBvM74eEjD0SDukDD+VoPfEUO4Vo8H/ZyXErRTMb4GyL2kMQEcRrZambyTyVNCDi
PH+pmcxpSQiY9qQLx4hG4RXLY/XET+Jl7HPUAjubdAqA28tAItXZnbyMRK54JMqzWynU0Y61OS1J
V3wSK1NR/rmOHhHVNYSYkL4ps6ecD5zd/nA4otassE2Nh4FdFJcQ4hV4oSrpDanrr7L7qnoCYMr7
xPD8b+gQAkc88TB+CCNppHTfBk2NR1VVymZ0Ap7KBf8joxDlBHif9NABEXHZOKM42BCOdyKQxjUv
WilMQjKZaCLKQTOST0UUb0v6vDJUBEQ5HGkXdrjRTWGJD1WW69/dRO8Ubn3ScJUO72LvNAH1O/w3
JKec/vwR19Gh3VxIKvomdwrZ5ChTtUji3Yr8PjSErQpH5Y3VrcRF/VWIghLD7qP123eswWK/KA+9
VZtphq/HSkbuY+p2LDKSNG+kQtGFkDAQH5r+4Q0rIysi7lSB9H5T1Ny5fx0/oRTE/IcgotjdfBxE
9XwP0S63zBinpBjk2kAOjlTuZnL0xF5QKzDhNyb6cO+6PS43p7/TuqAz/+dfXdZjOvLkrbupW2Nw
b10LZxcZvCZIwJVBFX25DpAdGYBM1tndAlYkquWjJ0z3x++T5zoGIF+hU4T+2i0FlPlpRO5WcDJ4
bgfdLz8TdapBPLwQhVjdz1MjO6FnRPv+8FjoxUQXKGGTMW6dFLk/U0TcB8v73dJTjNJtrvaKDdu4
aMasz72BULyl5+5/PuPgMChpoUSOKL0g3XtmIV2IH0awlsVQ7Lks6MZ5wypw4xcp1Jel5kNYAV1I
JDZlvLCvitYJULB7El2l6A2qeUSSV2hpbzeCIkr/IcN4lVRMINWa77EAvrLKgNKq+PwK5aB8qB6P
6wqeWsvtN0xCbMbmfJUnBarniL4a5kvE1RVmpp63zNY+ORBqMUELfHkLhoaFT1drVrFhrR8KuS9q
XO1R8q7iE4z6W224Bexm1vbIAgIjPOlGb79pkeDctwMtGC0+DShTi/ohzWNtf9VZCnJmpN4OjQau
Vtg8n9CIjPvCogf3HREwSIaee4D+BGVPH/7gye38KcMZwGgAf/dRsf7tkri7LNAsIAag6JukakoF
H3ttwU4MPHBQlS+buYNKHzIX60oekpHi+/EQhxTchiCiZ0kQf8nWfY2W3F56Z0sqY62sMgfAU94Z
vokJoqUBk3A3F9TTQC8bS3WBn2HCZlhrNBG4Q6TYiilaRq1ovD9q9Y1G9KnbwbCIupGmyNSxeU5w
Fus7vqBZEbf6kjKoTWpn3+ULkbDOZDj3Qs54wX0NQUOG7BqHWDbWDBY6Wl7MuC1oQ+AtpNoF3uDq
PmgTBK3OBd92Kz4ro+Gfb/sArlclonVO1fKw+fXodT1LvCv5ForuZl0HQUSJ5uJVk+gEU7eoTZ/W
CCt988kyUWrVV4eWbG9dWdfEe1q+85TKFypbbsX9r3ZLlvYnn/OLDfdmNmq2htrSuXbnjcZ3CB5X
b76jRDv7DlyxbfcUDU9u0MoafZy5DZGpdbx4+dlkQyVAWG417nzgG0NwuZ+NjSMtSEzTGFsmOms3
P7Ge4uHdIfObTIXX6g9oykcKmzYMiDN5W5R90GhRZSvW2R8UE4XfzEct/v7qyCztGde+GGP6Mrr5
BHDzbAXWaNJ6mMxBfLVh4m23pSlla+EOh9TOte3CT0fHqfxy8C41i6cZZgxK1QowKsMYdYpjQMvd
d2WfvVyIhwBV2mtUZ/d4JvQWl2rBahClVTcNbnaabQx+IjV9aVmwYEnPPlWSw2dfMrV6QHJZO5x+
FaFmDCuZs+drS+XJN++T4gagoJFeAQj9ec7Mwg80EhQneLwZnZGUSt5r6PGJPKnEqkXpiCo3femU
KESc2pYcPdS3yCh+mBqvA0f+iSQmqhn7q2Ra8dk9X/R2ulmf8w0MEJGUG1RvRNdzzuY2olDLJu04
tgh1ztMOMtS3g942GEW1mJ8MjSMWFdx0mmsTdNnYQpzUrMbPWsiVl4Jj40qZw+Xp8PZihby0q4/7
S2r2eprTGMqknrDia6V11/ElhmbzpVtqKc3r8c2eEW6EIcpAHKfLER5cakN21f5LHm/arbJcWJnd
usxwTruMg//WhTOe/+HlNjZ7MyUIDnZ8X/HJFpYhfGAeILzbAh0kgQ4gYKlYRRcz4ZWpDUOfc9RM
DJ2Wz9uOIF0xmtZY8j7n2vEKyk/N1XNP7rsFoi/xcjbj6mUGfvfQhRu/vu1uNhoKXm0VqTo+n9Da
BkNqM3vWwKySd/Gqu9FdR6BOTRiGbQdc/iyWvNjOJqplKRypkLNwAVm5sGXyyfA+o3CK77ByQx6L
DdNvpaqIsYnh6VxMuYoDE5uDV1uP7Ai3EeKLAs/x3eenulnYuCzRfq5qkItIjBN8eQCMP4keFk1O
K4+sz7bCCb1Na5Ghfk6q4b9vWXlsP5KHkPktz9QnvXQQvs60IddovD8k631ZMM64ZmQfldcYHD/Y
8KGJOkunrYlZ6NNO3uhO+/hCaNRm/LLTaOcCVQwBt4mpLmxPRl9IsUuAirmj8tseGHWlWlJBxMN+
jm4Yr11ROn0bmT4cITQRgLHWZCOj+AcyUVRi4sVeLawVxxfyg0iTbldSTdmFnNr/Tz9BbM0S5Nbx
WRFACV1ybCGOP15Q8QpxSkmX+hdOwaLZcyUqVX53X+lHcGfoF2QHzJuStz2Zfea7WXouUEugUHoO
op0T5A+dm48ymcEUyqWTBQG9awv1Ls/waInh/SKdKC9WTgGNRhmOsl+g8TT2D1NbNnlvYVjDXkd4
tqyS0vRhZYKJgA46sVeKHSX0WUD3YOmgYg/FetP/YoUKe5E1u6g+PLczfQGoa5yKFjfsqBVkn8dO
9ubLqT4XRwr3dg0Veiu0wueaRIrXuy12BETIcAFK/ZwqAkxUQGwRi/nNMNtQgifz+oFEUFbMB9WH
zN/fVObMsUuDiQBBWK8P6ZzaPTs51yYWkNXyqMRAlIzjCCaxRE6EoHp/hQYDDlDfZcm3nIbo1P7H
Uh36DR4DYboMX5L/+EDsKc7YvQ6waVZ91lfT7d31uHvoeWnrHrdPJzad9nG5OS/6eil1bmOfuR1b
qSucMEqSJe+VY8Ctqcx/VRnca59V7LJExbDTGQACr38JZgXZnwQU7nWjD0vCuOXwH5RpHzUlfkoz
DKyFuE24HviJh6d/PjA+sQ2LvGgZv9IW/tlr6jn3ck5xXTkuziwG7HNDeGnwY0sMSyFLzguldHbI
dcPd01hziF0ZJJYU9UHdoa3KiMFmeCn2BCbdeM9v6B+QHCAFKYUEFe2v3uHOLr+r/7/NgJK6i0hD
g7Kg6TgGAlo685OR6Q4jV9N5CHHgzYm3PgorBZwaEN+EL8YoUNFROozwCXshLfrf/nDd7NctcMuC
KKwY81cVYxK5Bdqjzr+5PB5J6qo4KFxKBiWbyYiuxFRIij6sF+s2gMtvHDiDulpV+GvMbyoPhbCW
SIXiaoNzyuJ/yoEmLcqxmgoGDOygyTT2LVV02cz0bG12idDC3dV88dsW29xRvZwUI8LORdY2glKp
jEiXs04y1Fb0PMrF5kYDG6Pw9fl+GG9i05tldz4KDDAGhH8fVcK4bJBMmOO2BG5y4CEfnf2AmV+a
bue6n/4AbKBEd50DC8FmqA0VGDcUER9FI5RpKnwTBR5j5lMiYWVGsrK7PXgBWcONNlQOzkfWCrCd
K64dOfu2UIBUaWuTQT2dF/qQ4rFnsCBp4lOZMK9ZCjFv1uwRxCE2nQ1gqgV8WWXMifCnVhJqku/a
9XzQaHYUlzlRbvbu71w4mgGzFHnxWvNePYVT3KqJKgSU2pquE+WkaZqx5HGA9+DgkogZZvrctBsx
utrKgOrl449kPR1OSfzT+wi3FfocRP26GbsppFZGiHwsJUoLgFpGG+GC8nIxrX4mBWnv1BXeyaQA
7SiB3UIkdfQY0s7BoBWjpcE55Db9bVgUsSpnlOonfCDy8s9yqnhtMBj5V4SpV+a29fqtyYho1za6
lGD8wM/zAwPpb4dSqcNQjPyPUG/ettE+Ar8tHkSd/hhF7QWRIyLbeKsMjMXidSoP9jap+Az8aETU
l3DX6z4Du/H5aDj0G9KnqbwNAmlfl00nFA0doD5a62vR9WO9UISWqdrfuT9R2ktK88BvfKM+Aj2C
DViqPca7QIB76yziq6tZ5pk2WPlja6PR67AXEVG9DvtoWSKCCNwbecn4KZzvCmpAkAJn8SkFd4Gy
iWaIaUhXrSKKvokl6jaVsrAuwgX0H/W2t2FxKVhsFuFT99W0gJRsAn5MpL/eMIWwnw8f97JjdRmt
KhX3857h3JWxjiEp1uOcOMrFzO7+G7ASA8PK/fvz5KppIvXEs8xoSbRJuoMbJ6ZrNCsLemniteQU
j3VG5DmKwJoG4S1hpW3z4NVFgNM+EjTgNm4U1YjpN1g9XPhDBowPOy4u4nzDRUym4p5gfgggQ0hK
20fAQrQye6CVLPUuB4m2rbkaqP9cR1xJnl4WxKWEojciWWNAzw7axvb8UPS/plswwCopNCGZ+Qxd
b+Eogg4dEg4WJtgXUwmyY2OUekcRJ4lB6KRyrRmqjvXyB3TceybSWliwxWKLXPS2V9gRYlD4dhQR
HyY0vZEolp1RtK++abDtDIhAj2eVkpl16dSyhxow+HtVv65JQc1vC+mPFxY1JoEf3f6qIR47u21I
VZnROOiHqUodOygYBIBOMTvhbzetMeYYG8tQGXMcVrOp4bE5ReetHansutxm/5jL3TsfPcAgCG3U
KEeu8FqkQMeA7BGthmuqL4pBpJVYN7bdkLD3yRWcD4HPgywsrGYY6SA2sXdiLtI6KtN3yOAE7ZXV
b0EBgSJrKzyoJ5y2cGqgT+Z81zqMPPf4Tk59my19ax0kS9lEaq4OieHzlh35z/YdCSbQsH/3FjAD
33LKwOieQ0/Q8KT8Nef659A8m2iuqQty75v2gJ5O4y5RwcKcWzsRPwMxpR3zfB1uCePwutSv7M6I
XaleiqB/t4qgbdQtVn1McZF5t9x9uUyT/3MO/nQ5VQNzKl9t6e5Ie2yLBCdanGkHGUkFXJs1I/yy
x6LLtamo4/01+/G/cehdY9fCJUIjyA8t7PfjNiWeY/5c17iEeB+7rXQo6erGzaxeXKaEQuTPbv0w
RUnZkdIxZsZbz9CW6CLbzNGSOcR8GeORTxtgFJmqbq+W9rgmTpS9ElsaOeUYWSDzycK8Kni9rDsR
yA1mBYWD+8rbLQksbedk68pTorIGsBzJ6XL/onqMvr66+xwb4HIoTDCikOa6tT64KxhHUlmhhdV4
YtI5wdS/LM7zkVCXyjZG5YJ+5xlKB+bWxJs23QAEsU2/9my/6X01dnUd0cvluX9JHiuMztlGBRFc
udc/Jq45vr7hGyeE1+fsN+rkMILwkji/wGEwfBTiCUcRtVwBflJr7irjRI7JAFHLeW+n4e9PUEG9
HqNcAPewcDBD01lsfCcdmFScU2cyKSz01fOH/VRl893wrtXP3aR/E6iWI72Ed7wwQZ9mCLSUS5Y/
ALSyoTC2U9BCcV0WK2q+9UfIQ4P0a5mcY+7L3Bw31+FUt9DRleGu/8+dh9Q/WU3TcpxUptMRaL4O
Jl8d7HDRBkDg9wAMwj2L6HdCGFFMTVpmlesvJqL+1Rxcuz8oopUbFp9wQdbKjqi4zxc95NoznNM2
5wJswnKhDmoHnv1H2jIgnSIcaMRPcWlRUsYyQoJCDbD3iBWaEVs779zmG+9buL7cklCAUlnpwk/9
usXLQ25PIGmMkm+X+JJG6wW+HyiUJMWG/zMUmA97OqL0h/G4yazUyuFwhg73fgXym1ivFcAkA5I2
eaGMFO6UTZp6nv2YLCMZAcDIS67pwnCb/52itKRJRqc4r/+8ZOcnBcZ82sCBhr9eb3KmHxUckwev
nXvg3RfI8PxNdVEjRwwVu52F+0uNrpZms19V2F0nNsHiKsrKx2YXjvZUU3clm23Wl9Y0991fmjBa
aSKuAuLnw5Crezx5SplhJAbbbflVlmqp4qAhRH/8e8fC1M8+fKCHagwPRhHQ6FiVOhHvc21Qmjco
TH5oTPtKyzS5cN9lNgY3hITco1r6cAiOIo7ts4KCYryS6czw+nf+mPbooEJtnn4Zhs8yG0YmNVKw
GzNwzaAsOo4Zv4h/p7XCoBBlx2neT820D3bMCkrQnukzhIAbO3qZ/CK11ytzgXUMyMoKu2KAIXnb
mUk4Y/z7CaXWZjleihDH1hhbtni/XwgPARKq9sBmlsD1Z1vQRMNFbHpZISQjLyiA9MfWUJZC8Ifr
Og27P6o4gkL0HNb5yNhRY/MDSIMbI7JHafAvqsMr+L32/YKfew2I0nhjqpQz7CBz2/4PfD7V5/iy
zR3fUa3DpxvesLvdYHWYvmpkOfInB0JL/bnH/vEpqv6Uwx81p+GN4e97qzSBeMs7xbUE8TToubQU
DFewA5QfASzWojYUcWkwDonpOcZPxA1lKaS8KDqAYmgg84YX6lVKiooBSRNjuggb1w+t93maShxs
lWHK+Vn1gg/F3htmeSscFP1Ctg9SN1ObF097md86QarLTmPr4k2zW69OuMXvxVwsjUsRYaZYcv9z
1uyusqrPmKSEgt//mLB3kiDhnazjJrlpvWlwGRAwoACr1zKToBthG8+Ivk1Bc7KDhSeHTnuTsvl2
pgFZUGz+EzIn4ZCgYVvZnz/coghucAj1ICga8cNKDjejbiMTacCpu9cLHJt0Hmyu/uPhvm27wcWb
SlsLgqCXATLmC+kGcFt4+5vO40uB3rk5ktbx6p/bR0d3qvt9el3dpguT+72WfAOx/sK1E0yQTIJE
8HcuZxbc7a4xNKshy+wnIP36xhjAB8OXXgqREL+4E8lLUHso4nWAXWWeEj3i8NBwSxaFCjzaakhX
tEWCb9+VtyN01flDb9DESd4S9Kmm0DVU0fdA3u3kZpCZLRa0RrWMMi84uBl2XN6xw5cP1rrhsK0f
MsqWBuK4RSXrj0fuf2KoRrjjPM6P3MswG16Y48r/LBsvPlPDmKCs7iWDLEV+/9b6rEph4Pb8GK8A
4Bj58MXOp056TrY4+Q8cfROYIjvY5Lws6unhyKezS467/ozrHteiDG+3929Or1bslCH7xQufg9Nd
zZc53QqLnIKXd3xrc0zc0dPFTjze701hfl/z0Qofk+Km/0lic0vRFn10CCyW05Fl8zOnmmshJRmB
tCiws3SDp7pahmB1sd8NmU8+IIyjagGgi+KBQox1htiZEo0WNe2hrOXojXMbGfoi84LOEJfTOaTD
c7EDl3C+4ymS5tYWneIdXQ86gb1wEsGnXOI+D+YGMb5evblGCWmssjfgnt9tm7wO2QZGy6bcFYQJ
FDA6el/8FkgDpPrW0oP++0/b5/U/woN1Qpn/a5NL+y6jDzTXRosxGJHeUFQhmxGjXpsK2N5Hkp/q
fWAoG079rh/1ucCmRyAwCeYwolMFu65Xo5u/qLAO36BSiqPJot15JMQOZ9ua0V9At0byOxjujh2L
3afoSneNpc90DbJOu8A+WJhig4cIl7B7NNUAAipN3nPSGQmxdTy65U/vMc5DhtDCEkWVERpCAXOU
/7ZVoemXDp/SWNuVfhNdLg3JUa7Vbgrp2iOiRDpP5c18HWAP5YNDSmHHNveYBqlzcguYvOPaoZ3J
8TiqoR90PlUBhmfGzanyORDQtPTsCgeIjyBCj8Laykbn9EBKmSZKjleme3Wm4ctd5Z3lHTGU/k0X
kKII3vy+5DsUjMXqUjr3u/fAG5xKuOCV2qI9dDHLFygA5Kfo9HyRjyMeFk3s4tjfaCElRscYXpeB
VHhtcI2NcpIrybXAqNNM6f5Jj4h9iMqXrTwMDbntzdO1r4jHRGi2tfuijOjVO1TN12zXEL83Vujg
3piKT00blNoGLErhceAW4t23cPAWvRXrcjDw38PXNg1B7doqT0zQ2+61vWivIt5Y/hM0jnVtCbdM
othDx23Na8YAJ9sP3hKmKq+djY657wsLKoZ44nPUHQh3I7dblevy5lIpezveFm86yuUyDmaUC98v
zhCHOOPFQF3fotjflfHjvtj43gTZ9GOPayvzZOqCzqwhTpgzHQ0U1fa6HeNbjXUjorW9XFh3f4KR
/1KNom1jGbq+Y5AIacoJx+K/h106yW3gLAt2Wi3LikBnwp/cELO+F7d40bfBJ3dp9WT8VxLQHLIt
t72DGY2+hOmSnz6pAT1cn4L7UWDSQiWJEnxJB2iYER40FqOeLY8+9+7YLdpqzUME+TebQMbd2wtD
NNFWPKqxbcOWVP+p8FeiYffMHyZ/D7OeEBaTB0WC4VWRfp0iN9HChvDXEdD2lwa/ll7KhiedA0TH
8kOlgiDoNiDgOnINEemn6VHub56ViGZXi8qv3sogOO0vk66m8Tj9+kePn9ftLNrn/dTMT0mEIyqR
3ibxGA3jjGy3GZyG1rHu0xxWozTM/tl4xsXBvPmDHr1ac6ODJldOxpI1dJKyfZ6hqfNSKKyRbJeg
VCWw/YQR00jSyUVmh8SlXG3c0+zN+6RTksI4lgdnbz+mwv3YMlnPiCLyK8O/5KXJYpPjRZivr03+
7hHjoF5ye1+k7LV/Yhaz4WbKl7oLws05gqk68o3DHiRoVYvQLqoxcsAXlO7oDXkuGRumlJDCNXDI
VoNvNzCh7qSlTjyTyG2vriq3eLJWmsobt3JYJaMadEz+WwjD7QlKAPyQ5DYMZcFobaZ0mGKW2Z+w
+/a/+BdQVdQ8NoZ+7+wG8ZAcD4XwiplVHpx7SDcYkVkx6dO6ifqW1TxzeMtZRsnl5ZOR+z44BFi4
JW1c/yKaodQGkeHZxMdggvvyaIPQSeP6KVSEhIbhCyGcH/Lx82Kh2FsDFuB07HBiywoNzPZpd4FC
YAv+6rJZ529ghQHNaYxvcLbLD6w9SoNm1+bAvDUESBu8sOcGAjhKbIKnpDP2thjqTV0lFGqzu4fC
ozJcnLzT6rARX6t6nm6unI62HP/Rlwaotus96UNqaGYuQfhYGpGgtpOGn9wwyaugHrqWlNYCEjlK
BhgkajXOsRwXuBRxZySVS9qHp4QTWNSEi1ukE3SYIGrahu686pkqZt73lD9kKqBkeFTHMaSlMwEe
EJ1OYB6bDdxFaysItrRIPMGKxOKH+RCAjxjPbs92h1zIwtLshYItZ8NafDK1vQMlxUCGwgFEyT3C
lyZ3t2peQfi/JdzDAGpcFKkAy9ZDRkoCckOxqiDZpufsvnM9jUetf1iYyEh9IzZCdEhW8Fgg+jj5
esvTu1o6hhu7HTcT92IQ6KNgMWLBFKW11Lciqbp5ebO93RbDUkpClA+NWAvo8Jj09zPt9c6PBIw7
CGuyCGou/CHA5z+42/mmzRafMkgbCLktvFl+jwttKp2TIbB+44DTGadyVqZpIGWJhU9pI2Suu9+6
L+c03w/zV9uflExt8Y0ManAIqFwo1SvXAtUkg5P87qxfv8us/7NvfR+O/rOydxXdMjq81KlyG0Rd
DPHCZgOk25iE3X4QUVYEgy/FrIH3ggYNl+Q5helVRZMo2y+xodnKHetnE/BP/U0f6ojx3684qHIU
IH2a2enLYBYHIYmXIi/VkjT+XRpzSJhMlNagLzfYKbOmblvkTXZHhFHvifW+uh9Bq/5yrCZuBkuT
Z4myIGxzkn0psfNumck/rsHaWNnvOmFHGfQ7Lh+0b0kUFxuJEgVEgaN8mYuGnporZOeGfwSIZJtX
yT8LeUj//RxXUp9pZBT7Zqzh13UFoLj6GT3wnxVZzH71gvONl8x25zpDxEDE/MxYkwbcwpZzpYdI
g6eYXZWzyN5Mij8XnW8bHvOZnlaxMpPjF1wqGQwLNWhKrlS/TAukTKiPC5xLj3AygofXwQZbZv4e
GanK4CBRR159lkqyeKNd3yy8FdsK8dxFtgp7wtt/021hkTSAtg6Ukb2Om0Gs+EPIEOA6PJj6kZTt
dW99l8QDetFBkB5l+Z/2ZzmupJTvPPDl9jFlTZOdGxJBBiCEJfQEcblEIvDwT+TrdglNomaQ0QpK
Xqgy4fTzpsld9hB+uf7FZEDELmOoci6J7neI3Ak46Pf4DonK8xBsKurI7eXmlC3W6KyCn3JKZEee
1vnyW4PEmYk+PadSJrNktXX35EwlvDMoegwsdFrsNq1WwHFx20VCvshYsNjzy0oVB61qcKR57hRP
AdZgeQuRxuP32vvzkWsZmgiFnW0cBHEEqyaMPI3KgZO9ttyEWOo5Mc8sgb2Za36CWkWKyfvoMcjp
xoPtSfBxrXHXFKczXxp6XfUF0eugjW5IZsN5Ir6H+AaImSwRRczKrmDfcsUmKk1+L4Cxpg7oZMVR
YA0Y3AG5GiVgAfCHxzYajmFm9+nkBMaq3WN8xEuXipZbQvpxotC5xxZ1z9KaWHy/acirmf5XrZ+A
xyUB2dqt174EttOAGWhQ7m1z8WbQeM3ohmy8T4/HYgMvTRTOTPhd0VqieqzOdF/jmpyAUS7P6ZYo
qr6K5fQ6rIXBg6vF9rjfR8J7XLv40Ih+7EorEbEIe1+HCuG5e27v3QcW1DxaW954F4xFfGv5YCBe
EIgXYzuqftvZ65glReE0AuKXy07OB1RTYTh0ihmoGm3GuK1xce14mAkyla8bgxn1cqW6ECmRf4Md
9VZ3vTv29xPz5rPlsZGKGGRJjUkgQ6UxnbE1XpIcQIe8aUixnjv3Ip6gkSh2iBSUi8oCJn9KyTVy
FtWeRARctui4CN4iiacDq6XrGSZzu60vK0ffin/+lkF0l9/5xWS7/EKCIVcS64JEOOXvsDh+s+jm
n57OBBvNUjsd4A2n/MMQ0QRZ0pkDvZJdtmrZbwcPPWwzrU7WAZkMLe12tOLtQ0Y+26x8vE3mv4/6
ccgM6j1Q1ZDPo/RjGUfPJJgz4oAvZRWGdACZDAOsCHwaSaU2ZEyp8tMtM5I8kzJ02jUMKJzabbOE
ZdP0zMapyWIfvkundb37TOtcrWh4nYRnsUyesgt+N889hsFnkOnBnZy6oMZdS7U/GpC/TlNookqo
j2CiUdG2DwQ30PKuASbA4hkGdKiQp4y257qAthpgo+NB8idWN8rQKBOFI5bN50u95nQrSg/tnJSF
Y1Lxfaz3/d9YJDS4C1uvKwCK1LtlgF7u4qnRrOxQKHvLBQpgIeFnnCcXeQwnC3eeLjH2mI0rh96G
FpqeORmu31MWF3RQYBbZkevBYT+2O/MdtCg2+lrT+Rn3KhkYLyDF+/Gex/HGrypiYRszRf4oGZWm
jocweM1Fyl6FZ/WICsoxSr06KZxjlmGWSTSJ8+UrggTSdbWDuR5y01CFihJiZBwgjz/DQMl+4uJM
YHe5EO7tUABKraPxw3IRAxjUCHuqVxib9cBINE/7cTX7OVBZfRktbnSUAboqdIQgkuN8xBPDQTVD
HECZLxtzjs2lbja3PtgiHSkDCSFjA8G1proqJnVwHCQ9JfzsU+LD4MDBEt1bRmfF7ukuniSmIg03
SuKsumuMn7honxuGGnpD7k3qEpvl1sCt+2sh+d9/3RDHyAHHiz9L8lGHzxOhGCldbaOquXST2E5z
qoNyoCYPt4zKZsuNtBmLAsYuyGAyFmDsbu/TXNcdpvvQXnwFSpSW3u6ohVbY9ilToGTVnXzeg/E0
QYyDtc4RLo2U9TgDMUsPCMvTJevOj6AaC4m7OIbXRrF1WwowK6Dc6MOA8AGkIaUVaiLWqAtFpcMF
9hlN6iXg3G351wcI1cfQBX5g94Y8IbzoOhJtYaPmyyFnV84lx5WiK+Y2KxZwI/dEx2Gb/PlVwOkW
Nhf+MCpo2YjJoF2MILl9Vh98UjDPCmNnG1WDu5L60Ox3oMfstyS9COPuhC5S0MW262y2o1DRjbdQ
4L4kyaDDVk9ShujTrIj0a2B9RStjS0zwDpv3oD4P0+uaACbJz6s0jxSIhDVVj/YEO84ZJYsGXn0P
zut0n2FLoGusQphcCg9GZRCpr4JEM/GUjQToaHJTEfTvPeyfdjLiis2ZyFyu1HFOIO7tqDL6OsE/
EXC/HG+y+ILS1xdK7ERsoj8Pk9G+OFaedjDYTgwm4c+yNtBkE/bmbj9V4stzkBlBaTjrLncyVCk2
OQ3QbUVi7tDOlLdOtcM7JsKuDeTe1jUWhqQIDWV9twizoendt2e1AMpJbu9/swwhdG0g+75SG6IW
icIvAgkuhUd3nI7Grk6sfxx/oPy/x/3wKUxMLEK8a/JN227JV0+lyiJ4y6UOJKZUSGO/oYePODDN
1X8z5f1PbpYOHLVQ58z9hCW1fRtbHIOP/WkAQZFkMV7u1R1SPf9jxfn83lKSO7ZJ2pvhNSswmZY8
d9lL3f/3OLtw6sTQcdopkdP/aPHZjjesYpxqppuQDKPetrJEcdS/tqcfyv17ebU0eFjxJfoASjrJ
AORrEkbLR4amSsG6Z9jPQoltuSlz+hdufIJNNYaPmo7RIU9hVHLJhdWXAw5/D+MU0U1ppDO5NjDW
pnTOkfS1iHAn3vb68hhftoRjNlrjfBjCNxa9f0zJBQE+vH5w4xfRBWY4ZOewKc5Oyo/NfXtP57S8
LGbclGz5sQbVuugRKaB5yTvAeLlJm+up1UiDNA2vHXXgKBFC5fnPQF+w8Lu1DjrannWafkJZ4Pam
6IsjrIgsRg90ent5UiWuVAjcljM3KbdChafTi2zAPdLMFGwRCJBvwtulBXXhfi+k6OjpUztV8Z2J
mhoL4Pfngsf2f7CdpJ1Zqh0znzxw4xzCRNrIEm0sOdjrOLKa2PZmjBWea1AkOfKqsRGsBT5tbOIn
xWNdvkvgqczJg5ZhVELwxvOP1rX4TW78GB1vOxrXdtDFqBfBu//Js/wVtwe2qTMI2IDtRtibrvZ2
FG4J57b8oPsHcA5EBATmbYiT1Yndr0ijUDD+UiVrYrJUYcOo241ppUOV3COZPQQSG9Jofxw4MJFL
339jzhCdNt2DXBC09GngNNbC+2UOqrtCSfS8qZSs/Fjqu+7i6RWtR0fVLERnzsch/7Y62m60OKZf
aSzWJGk683V5IPvH7pLRRugSQbZgThzNdp6v2HRwd2oi/7EhRL+UFrWDIWlHY6y+Crx5adowLe7X
P5I2Tv222eeBvwzGlIpzlNqyF81GM35WXxe9QAk7Pr6gmwmLMx4GjDXjlwHbgC8e/0d33HfiR7l4
XzQweZvy52YGakjTHEao1k5h14PsEn9FArqT8eibfCD8ZJbhcEyncxPuwHWdMT5dpKnopic1L9DM
E44SjgnAhfpolqyckwgbVaqXePnCvmQkQrS/AwaroEeTEC3OBugS4ht1dG7/I/PUBRllGMqiwhX6
DtTDMJAkLFBiFSka2vkLXEBgIhgTc5KUUvfISM1EKII/L4N16daNgfPdYWDE9obR/Ka7G9YGD5LT
UYCERqq3ZDczIRUMUOtuMez/xVBdtZxO/1JVF+ZOpGdrnOYN+rWc+Cw5X/VMRebEmInMHw7DkQAq
lwpj0H9a2COp9/1pMApKOlx0pXGX4t19rHzFpIgLZZvUMY5L+kvXKILnEaHbAn8sCcKp/uWHY6Lt
0UOEHAUXgBN9z923/TkuDjdtxpCqYgBmcJAeZrLL590Ifv6cqPmz524FZtoEjsZT8Dbzj5Rk9kLq
2JIGs3NF6mp7sDyzQ80DVv1SHMiPgU9ehp+owCADuO0dLOfVItb9+4Gq+zIoBot1BpHbQoWakpcc
pFKGNYsDaDyePVWf1W8zBosz4MbACgxh9YzHL4MCIlGAoH7i6agjLkvSEbTfZd2nySVQrKpBSsJt
DpD/+Egyuc6jZvvOKRn6sreOeyXbs4zurtiIXi9zatolZ1jBTGf19BdVbSzYfq1H5AS/kIrucu+7
AFRZMPfpW06Lh4hQI7l01BQJw56tSR1Wbvg5dUoiNUtN/fgnwh2KV6wL74dV46C96+au5409/9n2
Bbx7EW+NP7340TLL+FAsdIkjjS4L+LazMEJDP6VgiprtGXowGOnKngWAc6QbE2iarBYw0boRoek5
0dkGJbcINqptNApiO+ZQ29XoyiAGOXkgyOEgMA9rprgkzS8IlsA+bbwZOmz6xEdg+LzwlCGKBxPd
2QRUsjjClnDLdIAEW3Sgh7c/ji4SOqmntnCiy2lI8rx8a/IX2XHykbGfNlDzg1NVf5EKVCxZUwTf
eZuisKdXAXYTqiLB3FSKhLh/WBETBdCL1jWeN7fAPZxQbONiCDC1MwkueTc2qGUbD6EAF66Q/0lk
S4fZC8cGgN49am3rsOhqDUZVJokzIZA6sL5LHnj0nKWKo0fv4fv1Q6aGH89a9XGAfmR9yeVWgwvc
IJcWiVeYs9r1/lx/xWsc06V6T5IGb2ncCLoTdTGJuLrrSlId9snPPEyaJ6hBKVX9y1yOOrzG8z+c
H3mGApFTm/+LofmCwnOD17sSkgMgC2Vlvb+FIUdAuEIJjR1AFauG5AfE1JROTr1UEyF5VOTAERL3
JwU/l1Bi29TMZfGbGY/h/JTwFLFtYtEY47oWLA3LeoM0us8oMutncTMndLAvPFMs/OfkLpwyB0Du
ejI1ol5HlW4G9tJxXuAJVYxbtO57zXw6BRXSaiGq+jcFppdNJAqw8qmXDX2AuuNPkpHDbf+ChHuu
FBbtidPeC+1TCETLmCOkEoS6ZsZfu/CeC0xHmIv3mKXTIm8p0EYZv68L5+KX1rf5IeBzUc4FZ5iY
uCDfe30HeZybli6Q2mFwP2Jvm7S119W+qRcHE5Nfgj/uQmRT8LbtZQJGtPoy7m0+U/lCgWAzqv6W
9MsmQ3CbzOqSbL8dtbdBBbkA8qA15scZfbCSbEXJaR47cj9sh4+HAydIYoyc8NckPn/nCIGi75Dy
LeQZbZdkydUr+AxZGrsBJme5GtghR9ab4j+Po8cvYuTCOHlJrqyflHny330rPScLX6x22zecWhuk
tghLN0BebO0r4/yK44BvivVUsdL3MTAhkeAXKsUVmOaN6h3rk5fWzOATRoXJEC9Nis7jfefJB7iM
uysqAcr3BGTEbQMWgt2kkXau3Hu5Dc3XacqpF9HWCk5tM2CF5dDRt6vxTrz6eI5RYL3/EmRUNO6c
8Ctnp+HtJt6UdqrjtEZttMpPLDexB+bdNxqcFNIAfyYedS2W3UW0jDORge17oP9J/JQ6BKqePx5T
zfOxK4naNaqWna4f3vH4wcVAJtqwRIoIo6MheKREnvlgBBbm1NPI273DjJE90ff6BXyrO0MmkLTL
doI/U2z0JfbQitI84bUimSdZPl5sBWlWoQUm69ic14LkE5s4uLwsKX/aRcb2tAzWUYtVU68WDj2F
lEsKuqniwa1mHufBEy9acG2+mXms0JSTZ1BvsaEHiaMuJHBSjM33YZQnkfEmKkgg7M/JOhxWmRto
2gkNQoSgTOakZSxsF84ggECQpzVospWOYQaL1x7O9AMkVmVbG99KQuCQr8XzlAJvPqtmHWOIUE1A
fnSxfLd3UgVJiAXgXHLTGugU+xTkLOwk8wYCGSrU0kbrhKFf+d4V/gHCvTRYIeVAohmx/5IIF+pC
QjO2KDoCE5OkHILfTh8f0WQEQ2F9ki8IkZZnd5/Sfbd5GG5Sye3tqtiUVvoZKUedXXaeCVZotZaD
mBzQiIHP6H1c2gl6gR9kG2gw5FtW6T1FmhqYr25Fgp9+CbJKE+uaN++dCA07C1jKc8xF6Lm1vIde
8RRcynFWNWS4L3QEMQBajhUqxgRd8n5yxX8BbQtnkST/s2V9WeG1mZxK4e0D72den6hQfyd7YF3y
qabeBavrsj9Qx4496wqmgMcgZ2eH1B33tzUDKoZ/WT//r/2V059YXc3SyixlxSGASB/unu5zVeoz
4vVvqClsbdAGyi754oOW2GA2XZPzOu/A0JEBiZABcyV9W2j/+2c2Y8HaH8G3Uyl0LB1RNY6GIuM6
yJnh151igskqSUHXrLk6KkFR8HyWf61TjuqKuKUCnKbOX65GavrrxEV+LcQeIDCgPj3dCgm5p+c+
nKdweP03iyxBlHIJxvQ4Y4/AXRvXlTEshoOIJQQi/oHv3se4n3SutPMLlZWI4FkMZc0/nDCnDoPv
hl6gsIhKGfqOV8Yf0u5p/wlXXMdlR0KBamAaTwRGIGF39Nj19CrR/dW0hFd4AnDaWY1G15RhJtj/
bHrEBYcVEE+M6Acd0QegPuo228QRk2p6eC+QiUlGIiA1EDtonuaUCN08O/FTFnukd7tJmBaAkLth
bN1/RQQKQMeExhIZmGq0vcXkzUT16EweDpZJtKm82OwYYWtH0cnQWtCLS+M+kwzA3DdVxml0z9oC
nid0suMmK5JIvFy/P6HVsrel2Y4HHyaDwzJ9nBNw+I/v4EL96sqWN5guDHXZ5V3rhlkPdEU2CeMz
rTZfTk4BLhIzQtaxnBJEgFVI8G0qLnKJPSSrEGaDu/XHzoyRSTizO4QxhS0fdi9KcDDkGVyQZG6y
sVyHPeXbX9fZrWKeUyNICmIKRWPcDKhzueJVyVs7eEFaj0em/mpTNgtUPZ4jngoj75H04iSEvkwF
4CgSPEoxsB6FpGnmX+2uRjpu56xiNNQ5Ek98pO8fv3fPUmTZxJJr2tK4DSbpBIYyKbnO3GaJ3/0I
o0utH1hSt73h7wWlpqS4z7LmtXPeHGxDNFbGJoDdya9H4sF6y8mhRKBwZFOhasB2etCd5Ip8IO8t
VXbB1s3uMxtYzKc3FIiadX4bauzXFdE5MmzLS0ZUJi0JjevY4HkI7VhEVOcqaeC8gJm7Ko8O6ygp
RqehssDuLSKstAp0WOdT1IkknIeF1YptvbxHSnOHTi9hUan0vKkCjetnZytQgoa+1jl9X252KtvA
WGkfsmWlAJjpCeGRFrWn3WFh6z+kQpKBBZcvEUl4cduHds9n9+NwqtXL7QV9WNIHH/XkeO6dCgDC
73S1VRIjw3SN12QQS9WGmTNA8zyRnpLm7U4gMbCfOH85MAsUIMc+8DlDM8IiBpDdGWXPbqZTN95S
VcGyglC04cmUjhzV9ptv0dn2pxUfpRder658lyfZA1f1MOKEeN7It8Sx9VYx9Rtq/sDxVxUYc4PO
do4No7z04IDSQw/Gwv4MeaSQ4kQ9o/vlRLmY7I9hXz6HD9KqzVFHkud6Q4O2BwszGk8StiVnbLB+
nMHUtUoIN/b8WtWysqilKlJDMz2knwI5bJFysAZ0Fd06CbMdHkRBuVgHdfB6oSFPzYN7BHl/Ldh0
miMXojEL5Ugzo8U6nBhNl9HlddNwBHM+9zZaPum+0NVgbuuECVZC8aYY5d1K8EYc148qMxULC61y
27lyD1knlSQZowe7y/Q2/xuA2/DPaKx/Sn381s75CoELqF80SiN+ySSWm7fBQo8yoEnMRBm32nTp
3wX4AC8CIipeIQDbl23Bs1iEe6YZ6djxAV6kb3F5XkPDH+uZb7iMetufMsrullq8M7qa4TXoZ9ec
LqvYhAHKWuPfhJoMQxJw+xo1E8l77hKRj/U+gWvJCj4jDPUsb3tLt3vYoVc1MeBYxrIbaS7yiIni
WAUg6BMB6la8fSqV0OfBpKqhNfhJgMX6JEmfr8XwiDCCpJaTNkLvyagfg/FIH07d/KvkU0rRuFXB
Mny1jf3sSP+euyzpBYfysXYWTjxk/bwHWhWh4xK2YFDYGTq56t0OGUg0Yqw/x+bO4WQad7QmlXSu
yqGvCraq7/sbKNM11/viohGRJOtmZd3z15wPJ2AoZCizff4FSPzRIAuY+hJsbidYGFM2GFb6YuMx
uSFGfuwf3Qfx5EnTjfcGHAhRTG4fM7uT/eMflmFY9jxs1m/nZgKqOyzl0KqMmDPoQ74u/U96lJz8
XwYI9KTCKFJsqcZOAydd2vU5Z0++Czk0aHeBY7GA/lH2VqPOaTDPaicol5HbGkWB13FDYkjRtW9W
wl60lrRiuJF9OJOY7gUISHC7aIKsTWK4Qqe4fvNAvNV4KN7b467IfPpiqiuIU+uixL3Mfp5RpMkH
EyYKImHtzeF6G9rhmEgeNmj0UvE9XEFFVQ7O8VjQgS2n4dkhDM4xFkCkbLDgdwdOWzfB51+hBoms
xBDDHDJaHAjPobEqC5Y8fmpFYaz7Hh7+CtE2vH2AKyQlykO/7tEOA0t3MmmrGqF7xLgAJKzpQ8P7
3N9PfPq3qrM9Wj9O8MrhVQdTky7VcnDGR6DRVS0AsI/8+Nc+4bEJnBA3BLml25cy367gOZnX+30J
yxDgBuc3mSNqHNia2T41qIkHIYiZiJ2GrWbKg3zlMnl91u/cm4QkwdPQT5mVDJoBSRom/ogKrSDT
O6LKEgKQnt7ywE1pxNNl3/Zlhp5dPVZn4SZmboWMQuMypnAkKGdj/0+zVBxkgeunn6NJrJ+4RNo2
Hn9CWhY9iAh7M0hI3TebDq47+RS56M9Ux7Cmv8wdzGF0l1PL9YEBZSpJRur5OdAhTaL7RgTXtEE7
jRnF+XUgb9ejJQoU3aZrvnPnQWoneNkodPuYkZJ5XJD65TmqLruB42CbGlDr69ZRPVVpQAImtJeB
mAQT7/Z1ZxF4qPu1W/zEjx7eYKTgGZP+Q7rigTeuSIQuPKJUkPYb/8UVLQH37h3tFSQoIL7ID4oo
HYTu1KqmRU61trTdc8VFnVkKyYLmrGdmSop7eew1b2rp4HP2h3o3e0Qywu9I2YIX3DoibWVC7JQE
WpWqI48nZx2QGtlwcW/Ff4BOlN9Kwqa+dOnlcMhC6LagRp6w+0AemPb68raf8WJxv4qtrR39/joL
NMGOCJsBVvvg7siiakCFFCY8DR6aasts/gOp2NNVJpbZwm3yth31MY2dq2TyNpQL55WiTXXG6RL3
dNcuyGdU5Kae1rY/Pam8MxlZQvUuPfMnuxAoEhMGCUOx8saFtjGEREtZvWqwqewnozCDkHN8CWta
CkexPY54f94QRw6mziSp2VFdOraIb4KFKIfJcdSKwnmu6tMqi8wesqM3PmJCgykh8TVVOuv6N5D4
AtZw0DMq0WHmLDh/+u5ldGP76VQ12He4JDxKlxVr/BXTgLssTeqA6HQDXlkKt4HlTEbsA6OFrGT9
KllFjB/TemxZux4U+nPIxXvY3gXoLG0uJYNMzDet75ygn6LKqWNEWrmgeZN0D7Ko4b5HBPb36Tfc
MLR5yIRr3P8qkvvZp5UKZ3cPdRCN/ntKb2kwJp9eA0b2AMxQWrqn7x8UmCpYtEPnm8g7F3WFBe42
6ySW1/dCUILKi+fAkdcCTi68v/0x+OiyFqHGf18WZlqSA7mTyQvXxrYR6YeoZ1+65CWX6p5q0tQR
wZiglLveUwqh+l6+O20Ch0KGNaczJJyrKwHz3L989Pg2Mxmb0sbNDHWi+ISBeY28wavhnk1wf5kY
YFIebhS6TOfE4MHrguNnuiAy7ruo0aQkUirliEXfFT1nSZa7mMbWkcYMM5t7+fwW6eR9lWWWvWcO
ikJ56uxYmzcAlAQuSdVCNMyObQkKvbs9b8QLJ3j80IUezifzyYIcLtxq4XSt4X4QUZbeYAENmGXw
q/6+yAFEqESFG8v8boaBinLi2Hb0XpTwTQ+QonUEs5yrpB97myQZoGcaGipshfQBzm5UsuGRYqWU
tsHUXsgBOToDC6IUS7Rrv+xUyETXI63PUVw6p5r191+EFAcAchioUvY1IT45GOcFUqNxeK48AHG+
JYfDdBacN3r3XI2jhmdGzrvfhBXjrkUaOcZgeTD2wSGic+c1brpfIMJ/kMO/IEFYJkKx1maNO81R
U0vNsSftxWXN/La7jzbjepqrde5PBxonB/0EqXRttPpXodeKyQYK/EAoqahnuPHVscjZfK9TApdT
XScHySYk2zp7k2RJgCTciqZdsPoNa2KRxevcJc+Fap2yEpjXaUAI+jcQcRB+C11mbZ+o8lbTpER7
+l9ImNm+MLtZPiKTEIrI+TB7oMRmwMPpelXfF/LZakw9jPeD05bDMm4/pOW4/wuhc550A+N6wfRT
zwaJFPyapbgP9dXPahgn5smN+wxhfu6VghJWeoNkWX4itnn2lGYMMEx+ihdds7EpsEgGBxA1DiUE
HRbry17A/ny9HdEfye2BLq9+j6q+qmLFtmY9GuS/58Sevb9PVfsgCLTxkfzeF/d+UvEgEEPhQfqf
cdFaXXzP4BQFvAFpdS+HdvKyh0pDQyOTdOl7MgZ84McXSGFFPAxw+W+UEth3SlyihIExWRYZ4eYd
AoYqSIYxiydU8YUyKmJGAzzHFq46SV1vv6JAEjBEyf4WeKnda66A5NVH/ietIfKytRpwARN6QJxQ
+i0r3HQppujcXmiKqrTNyZ7X35GeQ/B+Me62G/tds7ynNQAs5BEZd37pdHIH/XNsBd59AddTTJtB
c1uOeK0/ioMBZ92YR48TIOdUKT3zrwZa/BYLwPtSWK5IwI1PSdJu6aJI3zNOZPrbsncxWkojAvFl
jmvx2cycTG3sU5NlHTC8RCDd0aPhL/QhQyFHl27v3q6oOwKHtTOy8FRmYRFLfTkcbPtsqFA31Tw6
WwCABU6lSjCPooR5j8JyOVyujwutJVg8TngWaHiTHV6kmLuPsDVMgxHX9JwgndlP2Xdav1twXcSx
DeG3QJR1GFqCrBJSl/J/3+XtWJSdSzf+iO0y+IkR4ltpsCSse1fac2qlONPkZPR7e6/HyoC4PGR2
pUV5Qh0a+Z1IWsYwOoFIS3jSdDYUQTJkM7SzruqH2Wljkrlz5B1qDnfI5sw4soophyVftPmxehZ7
e1/2ygh0rIz+mlJDUg48Z2V4IFRILRnpIx7JvkDD2jZpBv6flcscELd2PBDuxfF4MDG4+Ruw5P71
jN489Hs9OgGFAqs9T1Gnd/S4vU2Z4yrl/WkikY6ux1o8HxbijF6iMoDzdwPeAZ/7nptKHImm9USy
DhKsNFUXdW4ff99YFny7Xl401NO7VIq6sOmBK2dRq6Qm2VqjKakJC+t7IfXnGWNThVJenzDe5vXL
SMYSTlhbzcHcY2EVvwLK/4p27YgfOGEf4Kk5dmR9LELFehKon3iUGUSOzlCelY0po6YqqA1DbTou
eGgcAtljo8HGb30H3rrym8XZnuYBz6nqHgOmDYWOX8XDd96/w9SF0mCQZF+3IdjNOHGGbQoGsJLz
RPxlkAIKnp3E/Mr6qZhlImokalP5Wl2HucojhI1YGuU1YWaTlSStrgee2kzjFjJt4rkT5cb8Gx6J
tv980w3TTj6osaxfUZFV6WSBMRdnJ3hKolNAYSn1WzVLhmIisOiEXLaiQpRswSiYAjdolpt82auy
rVBMF9ms6D2ofZt9Pu9zlwQBh02pRK21Dv6/O6rjeRMD7mNu1+Onk3Rq4qUt2xC7ri6q0h2DS0dS
QFbCO0BMALntH4uQo4tVOoInYD5mFqQ20b93rAEPVA5UMF/T5OGYTBQ40RFWEnyIEQv3hGL5HbN4
A5/HXRYX+vIo1P65+XyTJeQs4MPC5RdT/q4RcA76BP8CI0UGKAKayfqe56P0Dvnnfia/jpQCF7D/
8WkFYaLUyQqIFbOEJces9y2JaP68uNc0g1KCTAuVT7mBjg+YsLuW5ukaB8FlstPQdTCzotLamAYG
e9jOL4JTe4s5qKcJW42uIOZY0mRU+INx7J+JV064Qmg3e0HfEvIJ+t32YAKA6NDbJqM+GnGG3SOR
F3iHxObTtLicfWFb8GqkK7bCxu0byS4rS3EGdJJU6ajR3Smb2mtt3Gj+SVYQd2HKJHhP9lViLeBf
nwiDTBRP7Spc9O89h2lPOj0AOiScVHRmX7mv3/5Ka87Ng5QHEjG5/lXq29J7dxakLn8ocXHlBKis
YNJKOHjAHBf7FaVziEjwLFxyKcCJeVDMKKTAVzIZdURgHVMUWmV9RBcmjnDSgkxRYuTHD+eWERw2
+/RaoKZefLOi1Jvt2w9NkKmC4+PLPicVP7k1D5S6hQDDpmtfkWnEd+V7Kb/RVmQ7gIwbCyP4fWKw
LFxoo7Z8CcG0CBFghnr2hCUzzJrWFawZ73gCxee34aeHcbuWxncKj9Zk0zWyid6QChXil5zCkXp5
Qm7fH8mXe6UgdlJ3odFqcsuJivCoYnOVlNTMk2RaOsCeZJonO7gOkc1fDZRZHxOQnC/1q0vbYOtR
XSQdBKLd35VP/X7WivjWNSD3U8yE1axbyb9Huc9J+5UoXeamhvrb1OzdrWFwAxr7XCIDmXvI6cJX
+UIa1DMoCid2WzJOuiYaUF5gjiPGidq9HUYAtdSh5cK04CcNLeInBN/DW2yVY/XSS/fYlWQKMllC
fgcs+iT/14AES8+YmgXCteRg2Rf28wjHsi+qCm/i2h2vz3pFiVj6BWZAueL47oO3GfPBAPVwwoHh
5YwVAPiH1CcKbtODS4Vme5FBTtP7azznG+9HGDzWa+O3Ka0rIF9bQ1h6H+CR1zIzugcN0lnqegsD
6lZ8CIMX6YhIbk2MUHhurJ7Z+Mq988NLT+k9MwrM/2cc0in+BFRTzmJLgulqQDOB7jIbJ0EblDPI
4HLw+KvTahhp7jh0BnRDcT7LAc/vnmTihFLpLPc51A2d0s36ojxzzNtOYTB8y4m4v4zyQQ6RyA8D
OrY6tjl9uriCkkcOcGrNDi1IvLfcGDjxG7q3UJMzdM2+I0JNUyLxpoW8eVxBRT8kAY18vjouvSXy
cE1fABu01d0C9qDwM4GlNXv0AAjJvKVD+9rp5xlEsSvf7CaA1+gW8IJamJgwWAyOf819kbNyfgaq
P33i+33PqhfaXcKaMWdxMF3CJjlyyiGgp8YzBAgaQdqBGivLxfqIrqFqlb8i99TFEtkfpz0kWZXT
diIhPuELlZsef2UcqHntP793Dy8BPpHHcqrPpMBwsP1nhrboJWBZLGkpIi5TWVk1+Z7sVPLxx+Zx
ISJmpJ0WVheBIl2DHtK7GkBV5SPlLZUA2k6gOx4RZNt9SlMHccvmvQpZ6OLaIv6+9ssmfPhT+hTg
EthAIE3d2Ii6FeeS4Cj9MDMqCnaXfSHQkEaZE+b4NKRUJ2rZf85iIIVpNB32TPb3jKVuV9fKX08a
qlw4BBLxsZLXGOY8BYifXyNfqUB1E25UYAxgn9A8INCrU18g7bX02QuOq08AkhlEPvVrfSZqasO8
SoKfzjpCE72N3rJC4k1acV+v4fcwp7WfsWVLlStfygi2l5tMRSvTKD4rIvg2JAzFrO7D+d4xzbIu
zvV4p6vv1S6uP63GzMKJdJqYvW6WRaXePjjrI3xsAW1S3f2f6RDi+9HF3H5GWgLH+x1urWykRtyI
8NDhiMLTEfXmRHCtoWp6KrQgb5UhjLSevNuOM1rSC4ovXNoNmoUozuKTWeT2gxjNQWbKdmcIqJ2D
xBx0Pav/Gg8YKQVqGJ6Fz40tMLldfwQ0VM9PL0mhXumYrHoHZE1neb258yGf6ngTuGL9lG4TIKlm
wEBRdTGYNT0kXNja2Vvghd7bYihjOjenG3Zg6GkaEXDMrIf8+EVjZVtrACZ4igQ6MZ5wrBxzUMOw
Cm426DMhMUco7HYpUBwcwpJ4ZU9oKhP/Lyo7bQO77v/4cGSM7ZG2cFH6S0JPLRtceROrfq0xzIGN
bTmGPEfpVkBBXx+u8rgoL1mRMSdin0BLmjNveXnjXBkRDLk3bKEstArk8yAo0cqcFovlPx6YuxEY
cLiCu9270bZfzvx35mYGymZvOiDpaVp/YZiTeBmrIClq762pee6/iT9rE5R4v4oxmeMyFo3n1dbt
qvt+U1GIOhPvt6A86bsHvv9YuEjhOK48i6SUuPq53F3tdisjwjW6izhVDtaYbd0G1zA4V3ysKGsG
5ofwEmqVObm0oX6RsBT26CWMePJ8QDzQ3fL3pUPlJ4aHxtaBEs6IQLPPkkljtH58j9VHInb+iEoc
knD32f94o4ySrMo9KFIagX+3G10b9gvmcY0IdYLLEv32vVyKepxMnfg/oO/5c9I8TNYhXdeVePJ+
vatAFOPIhPWS1WiXnJdiPU1eyAzZ5kMLN3kfZKVyfSTALkzATaEE9NgkOlC6I3/WGITylnFbwwCZ
jcdPwdI7F7vLb7uPqcDqsYE/bGVE4o/Xn4g3q+b39LWgZA2Ytlr4TYLtHL1gIwDBecXFynnKtKSQ
apOoK/qrFqPKQtzKYftlNbKEvWbF9rdomXznLnwXZNo6fBWjqK9mNa6khN+YLa0Y8WEtkzn4myBF
aP1mvADVCOSBO9ap/H9QbxCstYFe1CIiEouPka9agZy3SmZ6f1i6mvHFsDlfJ4deQ9z/UWb+uBuz
e4ZSMiDIvAmsY4TniOBq5F1QkhGA5OSUVXtPby8NGp+zqREA9lat6ULVXu8axP80OIaFPeQQBaCJ
g+CydD/rzmI5o/S/OlnUkKPxhM9Xtr9FqdnSwP+4zkQAUXWvZpxihFh53qwXfIv71xMmONebn8qH
wpVQtMcm2sDanVV17rr15OSxSCwAUn7xuJUS4QGjpnxQIjKF4sDMd9mWxtomutpQj9RNk9HSXp6r
lVW2sgmbbEpvvLxbI4OY6Ww9ou199DUtzBdLAYGSpQPI1uNRx4ujxOWi8WQ186JOdNGT1GujcXJ0
U9q1ZJVy80wz6o9Z8d2ELKCv7iL5IGqD52fZg2/fZj/Eu4bjbdOYfUVf16KElGZAGMDdezywatEx
8NMsXxDA+UGx6fTFOUganDQ0kS6gAdg3WZYwLNaL78mO8uuWvUIqzMGYMvH3KlQGN7RzzIXRfPzE
wyfv+XzitYjhA12sAZ749s/v4ESmN2PT2cpsbmkG60B9ff75ai9VAs3dFmDJWKNfeVnUroxVBeK8
Z8O1lg59a949yoBPdoYPNC1+YBNEvQ3t5dk8soTLs71vjDj2Ax3CGxu6aIBQgK4XIaCsSVdH855s
KcgvGou9N/dCxNfc8vY1YWrKSmkB/s7ysLQN7ncdbunggGAlmXF80FO3WitO2LhAQapP8PDXlohD
WgT0sD07/CSI0Bab9HSkxxqml4hpqZlclKErWpZ1yLf0OrTfBDDB28X5vbfRi+ywaoPDVbXuHR2W
jZVpg9mnHnJDlOvH5NvRt0Q1wh9PEKkewV9RWLWzBVQ/170Q78zrqcmszzvQ5TD8KE5KBjxeQF55
rdSgWWv8fiGxXspsy/CxJt1ivEz7Pc9J6GPgq+r0PyOTiyHEEGUyp6WzHsVB2ZRYRM6sPWcujV2t
GhIKUfEE/MxMj21Mc9wMrDrvuIm9QXITZvXD4RE/MjZbgnr7OC+c49bTzzmd4E5avAIA+REGhvU0
Z0AH4X8IlaX/gff1619yp9cSnPpgnW5KsnlIyjmO9dVsYDJMK/vp+wg+ti3GtaYFe7bZc4MXV8fb
2JnYSl3wQhlmjFR6OBWiPmk3PGoz+5b6H/PwCxdf/YBbnrsJVnBoZ2nM0SI8Wn9G8hDaVFum7+kZ
KHAXxOTRWBt6ZfxYyuf7ITY0BkZAJTXlV02weJATcrLrZWMceg6XwNrGgPEdfIac2zZRw5klY3AK
2bLMRdc9erY1HDGgN2napJRJh4hO+vJJ4LTVZeeXlkVI0XDJdJVb50+78gPyRA2GNsjKJNDZZ8KC
MlWY/xSjmz3NALfoAJ6qxf0NSUHo4DrNk5RbRol4BGLDPD4Qd0C9EKED7DGfgGiSYup1Mi75jmEo
ySKtzycSkkaEOH8IiCx6hSMhdq0TlGDztt1kMf+e1ge0sfeJO8yivabMVdAPp2yRPmUYYdOU+tY3
r5RSFJ5vpKjFuIJj39NtdS18tyQvx5nQxqPkFEjlRS0/JqWSEcSxaYoHoG5QQt65KU9T5PnPIkJu
ugXRKTDGwLiI7IfOYtBQ2wvWO1fxVk2nA0VqKmJtt0ZQT0OIyYpVVBK/WAYMiB0L7i7xByN65yDd
EmlKUwu0a8SF3kFR9R2p82fDgGR3gzuOCGec2MK4k8g3fuGQhM3R57cjzDCYqAtsJNxa/4nLpUym
7v9xO8tyCK2RMUSIdE1E3Au34ABsTbqwSKnFhLbckONkmceCOKJtf1HW/UKBlz/7u1o/UWu4gJGn
AySNm/NMKchU1VXKwl/zFclI7/XoXwXym0ucQsxaI9rrIrlyFQyk9fl0sNGe/lj2w0ztcL8CZTeV
ukj6ov18uMcCqnStNM69tyx8i7MdhkRtFSyCVm47eWnD8XrmuhB3dZiXEk4JgdAjNc0SCx0KuPRq
PLjZly0OXHTYVM7OaJ3aUAaZ5TJGPkIctzEPfeqN5Ekm8vETMUo8Nqyvg/6mD/qptvJX2jlmezFD
BTaznLbpZHQzLM4qhTC3f0NbS4XTBNYqjz4oeqoQBsu5W9+ZLophwRy8yDc7jpiTcA3BoKZ55ygf
T/PAMH48EFIu1E3fFKCs1/S6+SU+r7o+MSha6LcqsHGENYCYpTGw3n8qtDFENnvHfQQFULjz+cMf
+6H60DuMIK/kb28ecPcifDZPbMm4mmDrIBPKsZIuSySTfo1LeIpbrnDz25LfZReIFMYaUzVHDSHW
xG6wJh8podV1Um0PaAHOwsJc149esT+fmwcq9eJMwfrKka8Lr3OgfnDWgTie9bjGtSeB/+iePdxj
A7elVxP0wg2JdFTXMpmyoP+rLgoNVvaTIPr3nrvHFyu/n+cs3NgizonppqyKiH7wrPmlA44MGw9h
2xPqTny9A9KyR/NEBm6xaj2cK+5QgSDcQ3CUP9NhVWPILDMhc6bqCnzg39+4lBM9ObNo94vZ6Nu4
tw8vUpYpjVdIr61mkwUEDTBjjzALYJMyDi3DK7z4oR8Zvxde0b+9fp6K5hpsfSdmBaJ9/huvi+ds
xKa3xZMjVndsPh6s3cgWO4/Q6MF4F9K0xSu16WEj3jxkj/7pmGBsk2YtdGFEkkyAblJ5+G2qqmDw
sLeoYDBxGKG5Kqe5jW1x2R8dOLxedf7LeoHO8/HWmbX9QYpH6ZhTn/y20WtezY08Ol7AM/9CouD5
L0jgawKQykm7c3/WhTaYt96CqJAtsL9bE+unBeDnXu+rIGBhon1R+4ZyHXjFAulQAaiKkIwZUeLo
I2YDwpJO2jtUXhYKml5E7lLpL1F7S5acNVfl/Us3o+HoopXpQto45w6ZHp7EzRhBx1v2LNrGBnKg
eObj0H7BA4WXlEgNmAzUosSv6u8nxRVwNcumMmZIfAkdgDIonxkoasAB+Rtz4DoxZw24wbIZ++25
bnmQQ7zB1Rbemb4sNhY2PfUWK7rX20dZgDqxgF4YKelVpVT41HHx/4+dT+g49duZRcMK29zwHN5U
lurJwgbxF17lKcNFJu79WdbHk1ac3G3dveNE2Sv+FLdnPBmOZmDWuH364otAVWUhjLqc6YbNRDgg
10hX7NsPSmtqPSZ9W7ctUEi0oqDHS0Bs3dMO6lk/e7qnGgGFtciFwpCOlX2mLIxr00oQr60OvpP0
A0+l6kCrpz7TPqBDwTrW68FMjPC9BOdR6xeJhPbEX9iYR5PKvEAyxIZl+vi6xN01ciOmdnyxLyAY
k++JqeF8xmRwzXuyHeLnD7gGJKCrmIO2kqHlkZxuU5U4oD6I+ViWoOP3+1VqJZGxLqSUOzi3oKOY
ZP24PgLO1LGykEbE10Qkc4b/TznVd3UnZEiLmWHhQysdt25XXMwbc4IUCUjjf9Mt/y8vNxYGeueM
qrb5vcQt71jEx+qRfPID3A1WtNg2PYagklRU92UYs5kSuHD1BpBAlJWput6mEkmQwkJyoxpD0K05
8dhzTDwDnmr6g7DSm72lnkWa9Te7RAPonRxuE83B6ePIBHnegucYF07GV1lqIpL4Jvi0y2MAzpEV
q9A2OirF0CGPVAbkJtV/cUGGRmCRcy0BoHKG+PZJnET2X8WeDXQrdE0fcqc1A1fpseypDN/TQDYR
AgzZSntde3Ao+KpuXAbhEYWms+wn4cWbaLsQGAJRK1XwMHLRv3W7VyVaxwZDt8+atJrBez8aEtyV
kYI3L7QwwAvw4vN2oOL13Nvq1PkEWyUgThn1cgstpzRkhmuYuVLSx+ssinlodoCm82A386Opv4Ab
ZDZtWkcKwHQoo5/UII/1hEtLJVDFUirlMnRUGPjOIoaHJbhdqBqV225lQwcpJl+AuDv+67E/YXIA
MuD2pnjUdyKQRfnf92B35kRcr1oL+fcwulvDudsyttkkPd1DkLW99NSF5avvR479WzEYKD4Xxhex
Sxa93KHUr3On2a6jv+FZnh9ks3DvGe5vgrBMGZFGCmTtOuhTuyeyjOgEdExXdlcedxvRG3ktUGGs
eTNnLX9jckigE9GB/HvNq3ItraZaBtqF9ddy6dHbAZWZbKgfxmYkGeZBVJcRhxZFyMjMPdm3UzcP
BA8fNZ3Yx54rjDuLVA3whI66A5YzDCFRuHwr+Ad/vZbsejJaF0pJ6evumLjt5uJQCEyXDQ6O9oPJ
WO3x8AmwvO17pmrrsmwQTYKzf89smi3yTX3vHmJk6UG6HFdeJJ4n0v9kuLlFvse3k4a6M7l+tQEq
A1zs0P4lsI/FJXXnYpKHJAJEB/0DcrfcD9y1X01DypgrbMwSEnMKZpjGfTj5CuolkDxX9Cc9OQpZ
NzxN3yFNVjYTEcK1VUjezut8TjlHY+5C4nuHz0mNMd7uz2pAVLOKen+qehgVNNBh3S22IaHJ6r3u
Z+GI4gH+nRnx5WYvx/w+0OY/UJnKcMKfmAD5z7Um4GaWhB5JayF5p2Wwps2Iw1sETqgzZTQg80SV
ntiI8yJ6NRwDOPxnja2UrDxLObCirLpS26g3AoGtDIE7tHo/Th27MvxxkEoxpLbLEciEZEoRwlzW
tbXdzxTYDS4OI0rbXFm0lBVwniRj8KDo3sT5HnasArEDM6YZEZhR1tbqqr27Oi9DC9LyNz6OsEvo
P2K2dzN5KjOhIVXWv8fd7htHVwH1oRxQC5MXL1GIArOX9nKzIsEPQwSPqcBxyAROK9dxehKEU84r
FR9CdOw7UlFzj7lqLsoybQf+m9OOOH+Y9rlfTCvcM3vlIcszKavtjZT9NuKjRoEfHbdET9PH6p4s
n2UgoxDxKYOSb3cF0OvlZhwKuDg5VKSHHZUvvC1Jip1Ecll+msRGIstFxZXvEy1SP756qrvI3Czq
Hj0eoEkgzckFBqf1GqB82KpjEy5HL12bN9I08hZMo+Bhb73eqYPLSS5rCl4OOyCszXSc1WxuRZFj
GxHuOIWHA6UTCVrvXGUiA1AD0CdFtoV5mGK3Dj+C9INHQ0to+lf/gw/EwKLvmnBx9hjseNFt6l8K
7USNhRaPUziXLzh5lGkFLPIDUHuodEv36a4HhDDwulwsYyqeVGemTv0jiRaUsT5o1IrhuWi3D6l7
6LvqIyx47hD6Y1t/Nm5zAfsCGuJockNQ78oX854Uxj71cuO6pN95w0ZDC7f0fY96KR77ov0wvr+7
lgHWUussCAoEBVVkMNfwJ0ZoDbPZ/MQ8OuXIsikK+cK3pyqX6dCSUrFKoQQNWZhVEj1vYMLvPnfZ
s3krFSVGo7wPlvQNx3QR7aAsuTOvVA9p9KkH4JTiRSeZZDQPOCVGNLTquuoVLnamv0G0gedkSq+v
aLhvjjfBul6fjycjSebCNCzBsuguBOQBIc4U5IWn80oe60jygIxYY4EwxRhm/K2PnrRDvBYFPNAX
nwAnx7KLiTnYfSplfHA3DCi64JtJBUBGjmyz6W6G27nKgnEM5T2BEjjzTiUNmE1MwjeLJ1xviFWT
GWk+tvRl93/dY3s/OJE9mDp1UWh4G9aqZl5MAg3DcMf1CeWRB8Ls5KXxp2Y9BqlHR8LxU+S3cVzG
ISRoesXcGzvJaBWB7J7HmcsKJtN+ynw0skUmWeYrlleJNABQbgHlEuivOfRW54dzpFroiDjNIpqm
Ztxav/kMH5A7ihXjLdKIBE36RAT753x5dFy3bpXZavJeGMpHbbWIST7mOELGItCxWuVmOCCCTI0h
oxrt2qyM0eenef/bybCp8XqUd/wEvSxrW7UswZ2HKeD2r5QDq81pi+LkuOexSjxC8H4MHihcCWp+
LzdfZsp3pHwKCxiUy9RyfQubSOg8YvGzZ+Mi8L8jNwijbl17b3ByPlmdMSjn0cf3fKROoSFT2vDP
6C6Yd4OxqQYpY50p7SvVCowWHpOtMzglPsv8nBY3/TOSwA+DJ8mk4NpSVy8UHGr2kWpw3yBgwLXg
+Jd+cQI1F0X8aCj5lqjCrS32c4OmN18PEd2beLnH2ILFdgOGQYFoatiDjCSFBuzNZjL3lQkHYyTV
TgT7777zssZbXBUReX1+9zNr75gIMn/X8+rIAUm5MUXWLNs3kfLGXQFIjfkqDnX9q3TjJFYgGKle
tw8ZXUiplaJWTEY8gwKhbiUtRYz/FzB+3y5ITH4A5cl5F38YIV1Jneu8xzUIMEFynniNA2JuLFU1
5qaXsfG129h7RcydcCSIBuFprHOSicTSYPo7jdQxNg3JVVom7KAI8Yl5QzGCyVSJcQJFQ2WZont6
TfKFs5JrDnKx6ohi6mU08CJL1WD+kuPZinGWPL6/FK14lDymM5gGomUFRNOJip86SQ4oIOYFWM2N
FexhtoW897uTKyn8D+MrAMNzlr6M3SZr6kJ7udczsyKWskm9VVJsGKcz0GVcQaYvSvXFO1TIjv35
INvroKIRYGteRGYOgkRK7kdiGB0xAhgAmYgVRpkS4Y9O1169ow5QrMFeIt+eCxI8LufBTkxQDZnL
QcFDC46eUbs4uw/Ybe0k4MQjIjUeImpO1pU9M/Z7f8lQVYqJIxXslizJfaf4yJPS9n2wU0PsiPp+
HRc5hSYaZWSJ7jIT+Gp6Y56FN0ki6YEE6hvewK7gWCRxQiyhr7bVm92v+kMQ2Ix+cgxggUHZpYUY
+LLD5noq7eHJ3CPNWBtIJGggLgCVvnFpEVmqyQTEuPeeO4MA5ViCiJ9PdyaWK/Wy2LwZk+AExy1S
49HEroe0gqwir5XfpvI+rg5RYmTy9Dfv0WIUpDtMP8UP+fhPdfYHQzcywgrqcUSsNfW473lZbCZd
kWlXmAX9DdL5Z08RlE4JXcwXU2icZ8HJjZ2t1ADMQvx72L1rJMBhp7WmAtgcIGjR6YAGCkwaDkh4
PIrB4dpNqe2MMyF24YmoCKIkK4x4mo7bEdVtez24XEKbyFoNa7kCZGVru+9UNHdr0aIFhvoUPHn9
kQJlTyRLEGzgo92Nz5HFdIkeYdYcsTsz1z14nXQWH1htuEDQ5h/HFafCl7pYAvdtyPe5URvwarzS
8thXOROwwPZgDbIY+BLQgVlWxALVL4o2NaazN11VCC0iYcdZxGhq2C8MGcC0tShoAZPtGLPUhPYI
cHLJMKY6NkLK9PW+aw89BXMaF5JUQBApjwq48nk5+X4gq9FUoJigu5wvPfrIzn7AFEDheSMJmYqU
+9gUgaZ7mpTII82cPhk41nyn/GDmGAXwDyyLLhM3yLtvDJAA52n8P6vuf+cwUFn6zzJUnvdp8ENT
/xRMdSeoqqUk8z3fHE9HYZNehbCuGzluSb1vylimZuXTmXbrubopl+krZnEV9V1C+xquyccB5rTA
d7Wtswq95KD0UJCRzYgtWV++AGbYxjulHjXWRSfQrEVL570JQ4+RJbe5H3y0Qd/7N3b+i7caRyxW
U62ln4eIrVByvTTaGmRsZsWSadF0sNnW2RzgJwdoHjm5LqE14mC668NBWky44K8eUqkyTlA5UhQY
CQgoL7Mhq4OJf/01vp8H3sj0WcMjXYlLT+wqushOabj1QzALURV++REdr8Yb+/XslvBtTepdOhYG
9QN58i5koutphLV5uTIeZPl5bp1y0VELQVocrnvio3n2E2UzbSz0iFdHqWiQqQ4zBlWVPOingwHE
jFk44FzgU3PEIW4sU9ufmisQo4tebh3aS7Utx0C0yWhrB/ctkZXNfiBMRoFeEi31vM89wRNjkgo5
ZzybI/BaDCcOkEqCb0M3jYh9lN1zRsAs7Y2LeSVYDmXJbriRAigU5CJwTbdrR4t+ODB25RyqPYI6
fA4YwTvkZBR0pLjxTTwEj1VTZTkGxcftyvIxzxgydlljal9unaTUaPXhGEGYklkvgwMQ9dklkDMr
q7cenQSihV9ELonlPbBU641gtmStEgWtXqm89Z4Lu7fC0iCDLuxIK4gsuQ7hku1S24pX48ZDVF8w
tG2i4V2rEq/y6IWB9uLQd/J5Y9cPNBq3xghbwOBhYv3aL/7yzHuhcerKn2pQSnAIVCZ95FgjKsvT
e7yC0iI3fIFseNNeKXOWD1h6GB5ZzxtJ8CqG7bagXJvgsLAeF/2OJ/saIWE8KmU/o2jN5zhkamfw
CRQ5v+jTrd2eSeegHGg2KJ3/EXgoVdVqPBjcHId/nxzWky3F0u+MIIhKjwwGGDmJD5clHDqfltkL
y1q9t5YFdtNBka6XG0AXvXDty7LUH+S3uxhcgUC8piVW2i6tsAOSUaiEA94oDy2SJCg84E4lezEv
C/vhy0lsEYlHN/zf19N8MVtbOWmie2bvYgs6dDGVBnoJ96At0yqm+FHtiiJ8h3GpEWnOhkJPwb+V
RiQltQUitnHLLafamNLPVeaRXeLMcxZPGsbTEReHIUoP9Xri5WSMyLxe3lZHV+swwkDdKdqsRfCm
GYgZxi7hls/CvlH4d03xrS1N6XlFVrIBlWaPBnFrUwS65Y2+7oxL4qXiXrpnDWi637zqwCS+Fojk
6/JlPNavBOiT+cXn7JQhjkeBYlrLe0MMc2IsubSfRovYE0LR6S4BcqIFjaXqQ4AhSR/UdzLqHMI8
cUaPEE81q6hsnIaQOlDtCGaPStIj0jvOJ+L3l/F6P6UUMwDc2qtqwMgglBAi+GoCzDf2fOzXrleG
unnyWTz/jJfgoSTqQ+6RhE3vRcSWFSVKwXzZSF9ze5AUEHw29Ujc4K2Hkva6LfDtmRSXku0lJNVH
rMi3lshwEKmhc1eddHwdQoCYwwbX7BBwhAgupawkne3A6zZKV0oMaZAAfgsUe2eEKD5ESXOaxFyS
tngJhgr4/7am7De68m3CkHYB1wmlKlzUx7DHlk9YXRw4jCHqEp0m9pH3Ori5hHBpS6zttDlpwvTQ
VvBcCJ/bXnb3CG6MpolAVqbwUuSWl6JaDXOcZ8MO9KOYBHMF8QV56vvCS2Z+keupM+7jsRJ0c0iJ
t3wElCEeyBkIRkzoFk3/7XYH/6z2CqfYYRbMKxaDaU6Kjji5ZfIYLK28Q8CPgkcNhQoZXr8lzWLe
t6dSrnd/3NKJc/Y0L0iOc0gRHGQ03arQYKpF2u0jxNr/oImG9fcVwkx8EI0Fb5xHz6eM1BAfXLkE
m7n22o9WZCQlxK3UvehLANaGM7b871dBaaM6X9qsGpXogvb5c3gCcvAx9qVNDRNTC81z0Z1rOSPd
YMWhHuaIqzF5vLpbOILtG3vPDU7J8FS6K3CevkfH8sPLy8oy6gDqqN0lq2+qNdgJYdPApsVqsAee
rsmw+kAkU+2hHTejGik0olyS2lWFDkx7qMqgW1pd1IWDCsoU4BLq6/XBMO45tjQgKJK0EIeq91Pd
2V2B42OXD6rMmuFJdSDoQTY7FZQVH4Ox8zbQ4819CW1Trx6lg6Vr8xTRQixCjAt9SqEEQz9QiDF4
nSendgDerqbQiGkuJHAer6Xp34JDgI0xc24EPzWSnJPu18lBKkl2bM9SKLf0V/m5mqnBKsjgv+gG
iPo9ZpFU0wDRcC/Z4vVFgspxGExMr+FP/kRfzTRo92RfyukgBXl4y8j1YDwK+RZKrqEjakbT/wpj
IoxCdkCeuhkeM4QVMiCKURUThh05hngPIpPxiVMb4F+M//Ocy029sr/mg5UrkxkOF7GgMmxRX9Bn
col3im09q7fxcCLqacqEr1K6+OHWOmuGpLbpl0dua1TfbArq+ekZkNI805V8Iy3npfZLvQ8nb+Mq
S3mBHDYjZ9A/WMGjyXKgsvUjqs1eklKEXy5pbj89Puw350Dprj4/1NFC3CVZxDwTKXF6MPmwM7Wq
wGWtlchpf7JUD9wKa5VwzoDMJKcHE1NI9/vitu3s1ftqHAj/sMaxFpTza/qP5Y0pqutTdA8dD1n0
Vfiny2ORXbiQrYkwMMNPrRwqDYX66uIjrzJT9cNb4zptcTtIzNg5GOghHk3jnEMkT4lyksctlcIK
UR7+j7xCa9/P+PFMBz4W+CRs9P2a43W+O65UdGrsBsm/+sqOh6b67jJqKxcOpRh0a6bzMF1TFJ1V
FPwSRgeWF353nh5MlDbmivHlOegBIlV0hKbeuH/t5cJFXlaxP3TKDYIjwmSHHbUvZ2Ha5UbH/JdA
EYrzqkJ2XabwVcGFi94PcX/XLbcrw/yuX920QG975TWq7vGfBAq2wnXjsX3SZex5QDYMIaMR+zY3
yfUQ2GhhERyOuFvL9SzxwJErmsdsx9BGK85V0qpyiCrI8LVbgmhOaHC1DBd5kND/giwWOGhIm0Mb
M9InAZZGwJMvLCMAR0fx/m/vgewJ+qJn74ZINIl1YtGZKg/konayPoAUpN2ztfSgMXZPA6PezU0L
aVWG6W5d/5C+cQrr/oDajEpurJH+nHLQ23QNtNAAxW8ZfrQFO/JErPAGUfqcho6VKXAzBY5lkh6U
ZYUrGIGYg6PdcsigKcFTXSxcrViLGZTDlqDXO83EzdiaWObcqimsMFHCRfCi1CNaZVDYg6w9f1NI
rWWRfChgzaMjtrQKXYWNsQ+kCWuGRU0SOAJ0XStGCUxhGVy2kWVyJSZsIKyebaxUjE9JKhVRYARm
evl1Rrk4ahECWFYcTyob2riJGAdoB/lUnAm9OpB5OKevNTbAWMEHx9Ar8DD1GebDHn3V2vdQadmf
CjFyvDOQW/TyDlM9igve8IskN7/72oRziHvkaOpTbHDZQeeMsyk+HYwhGpx9poq5Nb7+16tcBN9p
MfqTabQ0+v8ePwctOh+w72yTY2bqwwwjdRfd+m063ujcLn3NhEtDZlE3w8RgIjlls5LquwMkF1C7
4tGSgkko09netbdeDBA8UFdBziP1nVGmtGAvS2LGKxSS6GC+abCW9ibOx88LktD3HUlhot3gPt/N
v5uvI2TNv3LrECaO8LvvlORqu1ZCbM+MvLTXP49bT/f5mPXYnNd4JCEIalhJLiiDbD3W2V45FFhb
sm/uHfqK4jXL52AN+TmHp4pANAXMoLzzAuaebhzX3cs0zpYufcOGcBC6v/YyLWuEpeLcz4Y3sAmQ
d8neBWyBhHs02EiRPiC4EhyEmbjsRb77t9Z/PqP3EbA7Tqxlcyr9t47denDSgbhOfE46VnqpzuSU
zdApg7IJiYyqUZ3cDtBCnt52IIUzLdiL8663M3gVc1MzWsLQTc41RbOJkMqNnwZVDtJfRZX1a7D3
Z4qs78IhyJsPOPo5zYMFzdyoZlCKmcdrz1EkW+3PkBhsL2uQ9B+iDFC46tN2Errd/+oo+MRZnWNj
xSbr5SPXeP5ZF98GrlyHkD4n4c2Qv/ZeTi6jVLrno9mXt06pbJQTVh/mSP07eFEUZYUQoi0gbK6X
D7cf7vwKmhmtvBmCaboda6gPtDt7WPSFoR57yO69BRJL6zbRobzRw6Hg8+Ja7OD4stbaFEDsV273
oYHrY1jTBDIlmNm5ljQegocCGgPxTIAJzDqDhEwakeVgNl8EqeEdF1o+punhWwaV+vAelhnTuL4Q
Of2gNr+/5aLwfiu8Txlfx0hrgwdn3CtSVr5oB3Aitzcr4N7dR8yVHIyvx1pOHMU72fnD4B5byArz
C+8ImcGGCF9mCfMYsYpZBg9T/ibeB+SXd8s+gL7Ut5k7z6erCdbLex0JXcliuOvbtCIxKRXFOEXq
IJBXAw5hN3M7eO7NQm89iRd54joPGEw4oZfq5yaFmSzVZJcc9oZ6E+oNrD0xjikrQC1TBKbi4bGm
32MijEtRWzaNBpA8OCmbdY0xnILqlXBtblE7o3W1DR7bAOUIbVNIsJKDb7HE7HfaDoF7Zn+Vp4eP
nWfj5bG+S7m4E0NyMSo245ZUmAKxrIk3BE+l8qnYJqgL9NopBR6czcZy66ytiAbc8YPs5gWGJP+3
kL4jBAU7eSL8RgmpG8gpsEx8ncxcyX4aQscz4shidq/DKB/G4Pkv+rGlf5waagD32/Dt9eCoPKDD
wt2SN/x38QSbmJYkTK7UDwqvH8FnDJAjT8U1ZEEB6WAD27e1rFQ0XfjMTtRltBtnzXcMZmFaI9mu
pdEEurUSWQiyhKcoOLAEVWlE76kv9VbLwRls9EO/OvemOCk2TS8cgap61RH/wMhytKjwD6bvhcjr
en2IHIkzGFM75fLwALIaIwOkAhxwP3Z7uMhVXNTuzhtlAmOBS61EEewbB37PayNDcFlcrE9cChXu
g6ol7ZZrxGOAaVujJgdbRAw5ZiXbj/ovLOOTKFvWTsXBGlWeCVAWN6i54cYr+SGgtggcBZroBAr4
F1/Ls5A7gXOraeQB6TlwxFTLPF8IdirdklcM9kPUvAp2DIrMMTQywVgLIjaCl3p5dOcEHFBtFsNL
EmK42T5NxqCINu3NESm8FaAEdSAdtwnlr4zUczToQXkQw/gZliEYnxshcaYNC/tVjz9T3+rEWORg
XF+IqHGltyn04h8No+NJgnP1P9lMiebqhypgakKQy58ut9wdUsLJbM8ujRgk/3f/bL4qJX8FmIaf
wH/nubOYa0qVd4KjjZXDQ3KHQ46ItGUCh49ZbCh+Ll8KrV/DGUNXMK495NailBFvL477DoM2vgCJ
iFcBE+vqNy01iLzzbJbsCc4w5G0BxF1OexZ1AroOGsE7NJQU6Y9C30IwinS4tjEQ0Sm2hyw+FII2
5TBkAjsIvfAbGUoAvhBzY99cMj01VaI5+rT5PuBEWrq+o99kZCpfu+Xd5hFWoeaYwoZawIzHNXGg
u3/Jk2nO5DLUwijNpKkDzIhjXPM3DNBdBMpu3r7xs42rNWGl1Y5zqFcV0Q4Sd3uNwa/S5mbYA5fO
tkTGJJPnD7EuE9FU7GTg/nutFYQH2Yciyzky9r/+bbwDXf1xfn//HvcNO/ZujP1TEj9It1PoVFAR
f3e92DjYioyGhLGOmfhcy6aI2RQ2jomSoLuP4pt0medulFv77HIYAPRiL1pFK+PvHiIaKv6Wh4ql
q+wwhoFqjiSY/ebTTIq87WkI0DggcgVabV/Fr+ffzbeGGs/8JoJNuzej8G5sFpuiSJVeBn+dDVW8
RaYsGhM3SFUL+7YgkwB/ouvQ5Aqp7Mb102VzTyHbsUjyJ9cgamyIxnEHiBuZDOVB6sPwK1fFEPt2
sHJXQ/Ylm2tI6syQIk/1HeU+JXyXnYYhxn8d2toFyuZbh5qN7g3IjkQ20/kXgSDuWiR9cZd0p9tP
yMNGXTOHhY7XGWd/LsR0H3vzECJdlkXw2RgkB34JQ9fQZVB8f5d/knu2+pNpk14/MP5QNABrfQF0
ROrehTKEZCX/s8GoMimBaU33IwO0IUkmVPA9h8ZiLOJg8BGgYKdf/84cOZE0KKlwmHn5H3P88jHO
l+1xLn+QZ/Pmdt0fCMC/uzgTIm9rCvI29RZ8JZYdyK/A11E0SAgqlPzw7v45Holbu242HLQl8CW9
DKmUs/H5QuK4KNl83QV7jxF7UnuRe/V8TIi/aQXJsdGbrln2O4CdU99NJZw3Ib6eswd3JMMBXnUy
bNyp0tTNZDLsYcqZN412SpWGwWoQxbOgyTNVMsikf90pMS2kfRBKm6/TJXnMngyqXHXJM7S0glQV
IduRV9TDYxWv9DXXhwy5qe1q8Rx66Mr2dqs/qyactOtqF+q2D+tT+EvhgU9UHkM+aTY21EGICAyR
1Q/cr7gLIviexyHAiTwK1XLMDXMLMr9QpTJDC/KpLaktrUEUUoE3YpuHfdfJWub5pPxNS/rItEl6
dVH3oKZnG8MmiAiCiYCc5m6h9VuDb00agWiCoY35qUqsW03F7EMoXaNSIvbuz80vpNymluyjihoI
LPcGgeFpikdJitipxdV/Zs48zqO3PNENjCl54uevshIGSystg9FG6nuu2Q03JDyRRK8Mo3JALKMD
bPft0pdJ9/onZNQpOP4f6/0Ccdc/t2HkWRMsGUW4ItKMlIffaW2afyWCGBb+4Ufd6SYux4LBxpFL
s9ayWtH2uzjdHsNZv0L4A4OV5K+ImtNfAtJoJ5ke3YpGsH7K5KFZ0tQyeMvV3KgvjBluATO+9XSs
6Th56Uuk9vPUpZGx5Nkd2v3GAmiVLEpF6EyAo5u0hzfztqbCVfx0rQX55q3fVhGeKiVyNEYVkisl
3+O32AlwulSmuibHOw1SRAEahXoQc052Kn5dD3WJ6yHW/nsnYVqb0xzEmrqko+O9s7ED0FZE36/Q
KuqJPKaK807DYZ8TQCP2cbDBXrRvBqvE8sm3iacpcg8Ok4hg9d6MDIc8LC3ycHKpf1x0jC9TpAbt
L9gsTYUV63yBwf3XJ+x6x3YohpbM8lGJwWpxXECkykrfzZ6gl8kE1qYgeFymoBBxTL2dEzi0MIYl
RuKvrXR5axk2CHAcHzRtb0vdDE8TYgp2DtcIsA1UH9E4zzH6sEh8/Awx6MF8n6DTsnhSp62eBGJi
BAu1Uv1b2jd/50rWhF6HVDaCZWMxnqxCaR+YFtwuTp5+qbfv6t+Y6U/oYAPNrbBP7f8RBNazAj2F
bSXJ4VgJYhh10uMpw69n1q5Knzh2QA+DT9vLS7TedjttK7x2XRIvvOCKJvRo7Tkdun4HiuxvrFQd
nV/aF2Yj7WcpGVy5EUGl7QMk1ApsVF7sBGNq21PXX8j+qKS6vnor7LHsW+9hzj7hkB/uuUHNASLJ
avmenozXXHcv29PJPfQkeIEPMSSJLyCQL6MQGCoKkiVtsXJ1Uw2IqGFhfqIMPLneIfi4VFYr03ZX
jyYORrLifezucBQXRPyYoczcU+Fx3rZ1cVgGna+gdBrYUqRmepbp2Rj7pVzae4NTMP1SA9yw0F9F
T0bg62JG+C0qVi+nxNtbD2AQLshNmUxYJXafFdKyp7Ft8wtGp40In9o+StNPXbNKaGJgIo6tgn+E
6TW8u7wlLWu3c6OCwYZnX52SvS1FoKqXTEl6311QBuNMlJfWv4zyBV6djgVo/Vm9s29gW1i8F5zD
PCSTCmD7eaBTlBrmEi5k0zP7SCHLzirSpefFFZj0pTBcYmIQSw92uzX5OhO+QNnA+t23MnBGnav6
1H9ncFTVA7xvzmpHoMK++K3kedj9mjX4NLcvr7pbAJ/t8EsTdpm+xOOLsVEdnqBgCVCRTtTaRChb
GcEMW28tHxy4xDMVn0+EMSIyJi/TmqSdC4BfWlzFjbAjghXnTkWJQyQR53G9twLir2R54bBkGGca
+1ZpLWDI/IKTeDTTEovWkRNMFzUMQ+Zlbmx5hlVzP2LLOrvvlvct8dgvOLgdYSJsGa2664BbEH0s
wvviFYK7UZwpwsrZvwJLJ6T+lAcql++8SKAmLG5WVtGcd9SBi/+PEdH8fa33BccGn6tXZGAyPK7V
U/mNu3QGJ70sh54y3UWuINkspaW0N99osCmAUqUcoT+mLHZvN6U4XI/uno4+BU1TREmUIWAtYnbY
bki5fg4f71ak/MqhlaZlqvdlmmOuhNgSqdRoxTBjLkxZEUAAFm9VTIu4Mrd3XjUFPGpXBzS6fuuY
hgaTjIEKGz1si6/0Klz7pcS3bcoQ30qmuabqWiPcUq3d4MyeLYZ2QL0pTVIXaPQz4V2g2nufaq96
LkvrmrgVIC90Bv+PwP3YD+C22+I/Nb9CKCIZUt4tH5onv60AF+o1J4QaCRohddLnooJtVjEalwBG
aF3KMqTmXtytGLdf5yV246d/HqYF2qGtM/WxVDWOZh+4UCyitrRMchrhDm02r+DmCeGfa8Ndx6U/
b01wJa/IZ4JCGOxgz/iyy/FQZRk5WYv66Db7mNWsY1jDLC6CeFQWKbZ4CZATHuA1xQukjIJ/cCxb
mDMVS8UqXpYWElyrYDiNiIpWeggGJBCZoXO8IickCDvpIKAHC6IPBCeu9vsEnPKVO+LVPo1QceKN
mAPh8schef+ANgY8DyrTuGXdSWmZFbO30df/Ugfg7LmJUrZpEBUp9eTgAALnhRHYFqq59G3gOkfn
cJHD2tf2VOZ4s9DgP2z3ZZ+2A+dlw70HKX6UHvJtcqbdYVA3db0bzI/xiJLSp1uZBipWx684BKAR
B9ALambF8kde+KfQvDKUPR9lwNkyXZLM6CyEOl2eSFLmKDKtHElD5Bu2lpmg+aXE3XHTJOXMKOG6
XanXCAQshHaRI+vc7b7y92sF3JfDDC7e1J8jaghWVzUZpp+hg6GpLwUFo04et+R/Bsg/8V08KKkn
sV4hh7WH8pse0fCte7LTPw6AgmgwlLvqH6nxKbRPS9ZNJ6IzRVIJ0DPIcvw/B5MHFCoNS1CL5mk7
13MC7/eyy+SA+653KuVIEDhyds2NNfjcsEgPCbJGWhLamsUMeZShdiB28cVHW0CUiNY1D+HgYEeS
b0xq4VZpxbfhxKOXgrqQErbPKsGAh5mTw842Ajg0801cwQEobJ/u29K4bH8D/SoHgwfyo40GKgx3
YW66Ldrxm0Hvbd0Uol92pcKCvN4vIgrjICef6SLU0HINUaqLUNmqo5LKDzuqgZkKpHGE+djw/bUY
pu8J2ho9A0w/kebmN4liDnZ0gP8P4eiej+dOcrZHpPIHifi9BnlryKysLrfO6VLGj3aiJL4XyALU
CwZaLo2LOxTHb61cLJsXEwUAovU28qh1cz1mFgddVC7B9KgzxCjVm9sYlD6a0xrvXJmbdZI1Klpa
ZDumiNH4JCNsIhNcPMo/9KwdWIY/NHBQHkbxMDWENxNkrRRMUK8Yx9Duq2eCHzOMR4VQLUKoEVOp
PnsAoLCZezQnJoY9JNp5aRhzwfMp9gco7XBk8hGVUDAzhIpGGbvwh+JDb7e3Iki7yTPS3/1J2Yjz
kwqxIeAlQChlikxc8FJhKbIsRRSVATgyvAN0cK4ojTwpWGE7Q+gqdOHXwLm6ufUocdNdIbENTGC7
oZyxgKsWcj/elAc999VoexBqS0hcN32noaxli/qa+r9DRFF+vEhaZgwwUG7RGxcA+hLC/4nHTZ35
rDY6760WmnFw3Cc9MbvnpI4n9b49ui/jnxAb56UIGDyvU0mN9uIomJfF0pCul9sEHBp54o/dhZCw
8NeI7uH4V8EZch64WUHqXerLn8IUcEpXSV7Drprvupz/AARZxiVZxMCPvL90njAdozxyEvni7Dj/
rE54DLUKrR8xRCbc8qk+HAVuxOYVgmn6ZTW1rrlPYYFWaz8LxrB0du0xrqh9j3kS9fysQN2F4WJk
DF1aLxlLQF+sQpBP+Q4SPvbYLRr4PJ/4bgwfga/nPwga985GJRkGH2Xm9w4crTE819eWC6peeCs8
uwqeIfpqpAJgpsOVLIWu1ineJtAikRsoT7fX1cEn6IYVBbhOgfpXtW7mIyMDjC2VCA8tbsrqsYyu
9VQBxh8nsDFIuNUfHLPxxUJnwQJSa9vz+YUDm/OTuoF+cAsKzHAz0WT0ExKZbyObISmzaDMGeX/7
NeAbhEhaAIKzAKGFS2VaO1tnzgNbVVqzuP6d7b8eLMSyyFaF0IlDl1BVklNZQMpOzcawBv1mqmUC
/gBiKE3q7hNWxa6qkQmok08M4b+4FyeHMtH28V96nGHH5BmNbWe69VuwI59/oIwPxyiEmGdSNOr1
ul576lwlgJbTA3LfcxyaGBmGf36nQc/Crxq47JOBEoBwySLEYYj8eqg6NDR9/KhbVrKFXkG2fRIc
+MlvTBoT1mFmwXAqRuj9CIVfm6q5TsHioU686gPygvXxXH0D4hO/+ujrdF176QxKIh8JWaBxYnxx
BGivho1kRU1gqlfAAXx4pJooPmIIE95BROc22sZqk2B1pNTmSo0hCTA5AUTYG2si/NMsBM53WCnH
LNUkAx2SRzryEMQzBuRMj+pMDPFb5dqhOo7iU+hIUuQDbvTt6FVOdNKdPovTJcwZbK+oD+6ugshh
WnX0WqzHlmBNInXhkAs/i4htFTr0sPxipn7PklvesJyAAMWaut9F0d71P9jQWXz+qJDZNxgl4q2E
gEKRkBBbKAoCvJd6QiC4/5L16KTtEkd+9Tq4U3RjtrWSL9SGlnTZ2EXlE5cdglvcAoJ0L2VEvuje
CjsFDsxgMKiP6FexNtvWyfSDJry+nOswHpf5ZnLrORv1afyQWkPk9xjuUesqxKqtAOzzDjG96joR
Elj8/ul3PXTkjYEmIyPSaPvPNF4thBuXfn9Th4eHZpYw/xw5lkZX/Vb+8HeHs0asVGHTkzmmcDft
H52QlHZ7UtBiNVzDW5dekT3cKfZXBHjS8sMFSDY/dkwXbzPzx+eIBwLqkXgw7PNyMbcg3dI5n/uW
huIxOkEu/Gg6xzjnAVzB8hYXLCQ8O1FJ8ITjsgqHSwvxYRyGtGzaE6VHRJoO+vVNfSYlVNyVTY0V
XjRwOxG9T6Si7nwTF+apBDD4Ea7IopraBHINdKCmpg7yMiQkBOCLyTjH/K+k3B8OO3x5Hs5Qjz5N
sgjrAD53+FUmdlEgCMuOVs/dseHUakydtiEVHiDzDqXC4itb9Gn7giSv7EKLaf57updg1fhPdilD
dBtZTntnzYaGzFeWXO8QmMJmbnJ/9SJ9ae5T4MgquRLvAd0fOau5s2q8oSMu1Ebp1RmxMKpe5SN+
yozxjVPBo2mpwbmxgnNp6ccL5UlCaz8NO3Y+AvHjjc1U13bLWTXAv2yPic7vgW3s3hlPeNTR2zos
F5jkNKVzCTwy458kvf1rb445X3zm/vBhqQwQYPf+5Cw3UssVXCCu+SvblKNIngjeu1bMvd4WVqfw
3fywSmtjyP5RZsn0WyB30loX9aBazHdfEKPfqEVYz7SRR6mEkRlnc4JL/3qFqMgqkKlInh2HBiyR
eR6QSvfa9Iz22qCAyHa5ZlcQVRvK/uFMY58SPeI46x98nRc3AwO9uh9awFQtsEygb2LYCiuDx1BX
MtLYukE74M7qhpL7o5kqOpAe1svh/+ypsf3O9uHwfrnsXiDsZ6zwtAsPvRMdOOxc4WF3bMHJGl4+
MYVA+vx5oPsWvv/4Ul6IECMMENRe3vf8EQBPAwe5CB9jizm0b/yYCQV2AqRMgcGj2RtFLO+NVOaD
vpetG35ahfhQCPo+C8uOf/WEcsggm2rcyIOk7ZvvK932olWq4KfU7qBSjMGvQ0tY2XW8mDNYm9CX
6b7a7i9LV02pCMI1eP8VKuVGxk2tLffTVSMzTnU61jBaBrYfDWKyfJUjtXw8Dp2S230J64OKP/HT
fqTFxLtomH0HGDkp9GFAheX5ABa36nZ8K2+ERM2Bo9YorPQ4pjdssV4SugizxLk0jb7HXSBtmyGX
AHqoWOHJ5bBRDD/C1r2OudY+tZdm35PMjDJ7haQHjwswCxlrbIu/e1NSEaD0CCo7MCh6TpfIhF5v
0cYRVbasx35NZJslsnHyaq/qcRcwd6X2qk6a2YQFPDp+rUEr1/SEshd1StmRvWq3Ak9tiCau5bsM
pgpTGESafkpKPN5ybYCOVcUCT6hcmNk8CAE0ewaUrsyWNgNB4hK/lqW7eB1zCyXJf0mb9sj9euYc
8lfUUG9fHvKvTbdGmT35a/+/FQrhl6JREpJGktCwcSSNSQXHLB5CCBRX2sgOdA+avp+RI0WVRHnv
gT6q0wjkbJzhqxpklDSZp1EFpzf5R6AZADKr33ShCW2qEKd8sfWgTKJ0/xT60COavOnSt8wzMYJ4
OeDwFWrZNAPM6EuCXO/sv+ZflCczjAbq13k3vqD2gGjSklGtRUeQZ/gtAAdWDaPSNFbltG86wMDh
j0liD205FmXAeDEkUqCzO0qapZO5t1lJKFUpwzRRh7S8gT7sdGMv6HkypzfOR4NjcIOREZGUJiOQ
PvNuA0tD4qEiZu10JIdJUXQODNNYWQHwPSrTi/aiqdfqzzzU0pWYdgLwfIyV3kqt/Ftm4UIptzuR
1kfpCxE+fnkFmQLvL96MIDs7oJx7czeGvzS2g3qc9B6JGToYoRqCzB9pv1i8Su6d/SrP2E1AxEQ5
+bJaWf6DgGUr23SSQrWuRsAPCaLwtSAW75NSCjB7Qui0TUA+FOodp6hDjrRyYnC/T5H96zmMCr2g
tK+wd1hU5CPqytFNPW0wvoO4NaTGTp9sOYMCz5JuYpqVzmkdAiDcPpjPX1wxH1JfZ7HZzsWiljXE
No2ZuBOd8eHdbMKigeeUs+XqgpLkX7uvf9QcIdp1rix47c39F+VyiSAXzT0Rseb0s0LjKKSA1CaX
gCKJHYlv35VerFTkuVOeVyiJsVd/OXYLBrICwfwBCEjLsDfXK78GnLtN5GCarUs6wmaR3sB7NNDi
SDdGtOv8lz8clxtjr9kkK2yRcwl0a6UgF8WwzXwjI9t7/rmQNHQZlZY3r1aOX6Gswi6SrSzWdTMF
DrTj2K9tdVKt/eS6et01Ezs3JlFIQzmyXRoFD7HsiF4xQLI7DWBWVDhBOtkUSdgv6QHeL2K1zvYc
to/Ke0aoMcsylBbhU8CEN3KmPcrHmUcGE7XZj+tK2nuCKUcWwhWb5c0v44zXdY4QLpVeeALsrYNF
rXaGv2+aegy3yc6E0piRPnQSZcJpxYBGd0fevqb9Jzbq9lfTJd7bIxAdZ9w8XkrOQIz2qxFLAQqU
sVus1a4FZx2Hf70CHlKyN8ZyIHcLyFoxztsJ+O9VGLoK58tc6bOtPP2NIUfkDGvIukpePBRjGemh
DKLhn2N4HsWlGyqvkQPn6Z9uQkAgtE71WFVpGgphFtTKxNBdGwCHVsDoJcyNOrH1WXzEA8V+X1+8
mfU0j3CtSmRVfVHB2QNG3THbI7WC9u4ij+03fpZFofNPBE2Yk1xh8IObSjioyDoB8XFNNyI00jR8
RwZr9IRmYm49K24c07eY5mEhXdSkp+dP0nQ31/k4UwbaFoK/kkZHMiAvKw83UqHLn1ylxyUzjZiM
uEfGqgh8YS10U00pR0IdZ//qLyvg+RNUZCjxKDwFS2YgSFZCgzlCKHI+rjjG+FjF3JVV/FNzv+pg
115HNSemvkmcVVhY/ucXhrsy4Xfp8ijfcWdQH+ZKIkK8f2SmP9QR35ir5RX2ZDdqWfQBIsw09sAm
QNoqKmqMrkzDqwOGADpC8kIibgteo9mfSPunROJXNXVLidPRP8Noh+b0z9Od9Uu/tXNex0FW8n1N
GQjqRiA11Qr+P46kvCpk79m5dvwXB1iOGBjqCSSH8zhoF/qXUn0OCQ4NDC02pLW9G2ANKyM34W9k
RDVdElTpTQvXWCZe2UK/ZSWxA62dmEqmQmNfoWcFB0cJ3+QkB6M0XHS7wXOBw5xfusE9eqk7+KGy
qsn8ZQkCenWunREW4aqjzrAHDZxzn7Bni981O/xynk81e2CUIdnbfmLy7qGFI5ECeC7pA17AMzT4
kgJ09XLX8esdik/qHSRz0vRQnwaUc6xBSlEge+4VR3sOlkILmvBSEVgh8e+meb1v/1EHflU3FS+s
nRNBQHWO0mqpxjtU/qCRTRXz0l3T2Agkhk8MMDoZzVSUWXzxBnqRnWDO4VbvYTB9t1SRmheBiu9p
sC+AIOcd8KH3qccbYJpp1OLLcFyelSwcaaAPbUQ2p4aDuthkiAXgPaqKNen5rbd6mDrAeYUmpnT5
4NmO0VvCrVnUfiHw0pgSXLxVCsxuQSJz42JfItoUmY/jmWrvQ6P5jwb8kpZUbKaMqd4WAWzr2+cJ
/bAkvj2XV8Q62n+sepDSDBmNcuQC7GipBAVNaaBEu7jtcgPCZUT9ieqD7LXVRSn0plTbfZR8x7qq
rOafhbd4NOx2yRJbhld/TH3BI0sa15f84rqMe0f7ftXNHovhmCmrADrjKdlnsVv7cDm3wmNqVfk2
uYe1UwHOLSaJKybTPL4fz5pPRTYqoMk8+Ac1igOBG4TcHfkzCWIRv+u33H1/k0KphT3I6YL8X7Sy
IozH5aPOCJ1NW3DH+K2vGxdCs+8c8kt2IZZJM74QtDnq8ouDqK5WPt9q64nKJfEaB4/tgVzXNaYU
ArPJ90Z7B1O3hr71dSPWEb8OjMSHhPvZWvSNlYAnnegafzVq6ncqEvsGSp6lb+GFlRl1SgiBWnxs
u9Qob4CiUYbyaEaPa81UB4aV4vR/Dvlfc1IunsWDYUl1t3dRoivVdanT6qoCeUD0rdVw/r1j3TCk
eTRTv4Yk3rjxemazFbJGawfhOvM95qIwCDWIJ7cGHdwBsbobF6hSkdt6n8foJ33z15L2rCGjUTW6
g+9fF7urYsFJvpHGL+OZm9OWmEMNDZ7xjUQnaiUwfDAHupNNUYVXOcOJbRfnktEDFW/k6RyIS/qO
nxxJD+W309aYREqE+5VMVLgPrprSH5HZ9zPRMZ6NLJpxiuteKVD7gBTCfyw8WdEb9A+yxyeo+2pJ
Om9PcQJjYS5icLIPJyLwl6CjVLN+mvQ4OQoyY8+BejoDdhlquxTdtIdEJo1vQlHvNu5UjJUZjUKJ
Swc8XhF+524Jrxob3H6/wrG+iyT9gNTkfljN/t6TAtujkm3IaVfwzDxIM0Cv6waLyYc62vbjPPID
DBmRwflykTzRb8v466D406Nq+M10ByBjQZTHEDCI3jMGjDd5sP7E5w7MRCDbu9qi5Zgtixtr9lRf
yUpASGbyhRAKlpCQfpOsJsKk4kYRybAnjSIjnzRcPMgQ+IPr7qMAEBxBtxgEx7mky5znvC/m4/TK
+DJJAyvonXORAaDXodjMi7s50psNlwbHGXwG97swCDbDTOlOq01OAfZB+tyEqQ3fWmC4t1W55tbR
FcSCcIJQbjPENUctYuZ9nQ3eMDfE6hFeWbxteUJk1ffWqhz3lOqPqa5uyiwnil/1kHSomz1AiJax
RmCzNFYGXfMKkxuZFeWwRuT5cDffjmSN3tVz8p5uvG6SZ9FSnsPJSG/TTMI0Xm/kcPVk0o020KqJ
sWPN53yyYMQHkEOycK8C5hvuw5NoJz2t6Y7GQRRQtTuaLSUr1QfEhSIN1HJqZDwyRcLig3mZFz9H
+zs5S6mKMdNPh3YFrOq8QgOxBMzrTcKUXH7SkM3uTXgxF3ghdTBamzlEOTfGmCVtx/NaPrRGiGwH
lki/AO6epfH3Te4CiKV9tHt28aTwp9BBTfJHuHeJCDEfGgm763TyGHsBOLlqevyl4NiDlxvPWJTy
1BNfOcoY0hSqWsWSJMO5Sxzw7phd2oSHqdEYcuqtjHum4z4kqtO5hQJ+koyizvwda64dEtNmKf/r
ywfQ0GhnKJaiHpGciaDG5j7tCC+v6txZaohlcPpkh95UyVkA7FL5lbBeBZHPCgSUk03fxV3uhoVL
EFNeub0krb1AIjHb2vaO0nrsi6vNq7M3VpeyBjufuieQgF6qjV+gC4Dr2GM6Ysf6Sw2NnItT2Gsq
aLRVs2tzJ5YnyXzqpESrC2DxwpL9Fk4l67XzitZabKYlHIBb23R9EcktZheYR6g+JSeS4YbsatPk
ThJqQa7OmEEGMib3ALrgrfIH6m8CNAFjBru2+NOmmVWPnt7NjS7b2I3wpX0v1tcultc5EXfJmA+f
3bVoaiYozE0UOTq0CMCADs4aBfQtprCtC64wGOweTDI5zB6+MvL1aLbd3Mw+ErRHizdbnzbWFvF1
9kJMlUHc/e+GC/1Z7S5ypyVUyyOwWypbJ+SLjdZzhtotOjhFgW20A3Wk4lJTBMS7knw7go+Tb3JP
GrMpBIpxzWLB76t+kcjo7CM9vukU5DaDhNHRdWjZ8vlb0+rHi8BfPslkEGTb06iG2+u+H+yzedqG
E72ORanVYyYuwaTdlQJXtanYZyeou7LbcsocL/6uVJhmjqlKiarnpaZtn6Jz6X1O5JzNxtZyW5mG
JueBtWlenzHegAUKOuuBfOsP62GS07P2go2S7ZnXAWkR4J+MvxgHNBGBcpl3NhIM/yd59f6+QvHJ
amiiYbBIIdh91dGK4MxZ61K91BeiiLNg/Gwld02YOdJ7mDzdtY5ybil8ODa8GnFhdMed5uu2kIRf
Q9SmgX+EN5umyUkR977Ag4/+fzpMtRatplWYHYUDQNAscrXJDbvfjX8k2Tkq7eS8/1kvY8KRyuX9
EKi94DG90wBHsbUUVTN0nNDmuSqs9byapYeDaBGqpw+D0QNg9WRL4bSq3NwxkoJckhupGgzesZ0q
PKCevUl+2FBAbpw4lHyQrxUe6sLb/llmuYjmNhWdYquY2qzPc/mJiVxFnLWa1yO3qPoJhb4ylro+
6+8fCg35NqoKg+iNfxL55nlEMYS9e1iAZVjoe4Q61VaFcvNzdXItz2dM7ju18eXzIQuvSPaHhhRZ
ZsdCfm1IO2GXxXavTDLImnPdW8lVEpQrifnHOFOUOqJnSs+UZysX7cBbAWEmKakDVSpjONP3HeYF
4OC0vKZ2H0EkBiVyN118kNBHl5rwaFNrNT/xZX9GzYiMBpoq1kMa++07WvWB7jP1Z+3y6195LoV+
VNrsC+qmCsxs6Ei7RxQZlgwc/VX4Su93NIV6KdQANiV8DhW+1u3+4V8koMeYm8GBJRLhq4q4nGgj
r94cM1/b+eDNKQsRgZ6KBc89xodgE6IDNnfS/VglL62JBLeF/5wc65m6mTxa38TecnUdq7hQX6ry
7VZW8LOQlnFTTCUlXA2hZFYvXOaxlSGXUZQU4K+1YqYQkkLg8NYcK/RDmmlnL3D3XRz6TEQc00po
oAVAkC62FTeJkzv8ob+OUB+j+y9MT1dXC/WbmZ8dsduN0S62aSWb70w7IWVva/xATOusnkcr6rWo
vUjbSCIrtwSi2/lsHzjRo+Ximel9gbQMFYxuVDPXCFBVASPsZMtRSNt5/OrQ2OiFngmmM720r6H5
8rkhtJigCAX+7GKM8EXD9B0cSP/Mmt3LB+aBtAZiT5LpEB1nWkQeu52Catm7eN6Jku25m4mbQFhm
ZgYkJt0uxuGAhP4aVcvOr7RmUV2PI/7/eNRm88pT9tzSwtV6U0GqJ42fPB+DY2mFMQwpOjLWTep0
o0Ur9819DIKwCAVhe9z1GmkVZTrRt8PZ7OFxAxIjUrJ8p+D+6+i+yOE1sVcceyYM+rBkhHd3kN77
+SbmW+sJST5Z9FMV9C3mhawRKyPD2bzg7mDR5ubfbC9/J8VN0kDtsWPjqaYo82Jm+ht4v1HwVuBx
9iosrfQlRud9Zyq9TsibDaR2RXgBKCA09bJtrb45nU4rHAaFGZoXh1pXl5U4e3QO/3Wabx6j2Nvk
jaKY2YFuQHi8GJws+1ZzuuX1tb0WSCSOS7yMOtX+TC4aoOr61Q/Jdq13dx/N8pO8lOihZB9MhRlx
uGe+UWRIFIl+P5F6NYoEC3iKVeiu3pB/HpcgL1EpHYkgiE6teskW8PpLN4j0q7s8wLyWM3zSoq1h
eKacv3xutd0xjTwOmP1T1SEpga0+UFT5N/unjlxdzo4BSlEOWcejeQIzkvDwA0G+bx2w2aIfLtL1
7RpBxeOwg1InAo1WrcVhs2ymUo6s87JVkb0DL4nGVkQGhnTOuQ8MPwsn8cqVhzpO8Pdj96+RZMll
1QDG7p1Oovk9cQXnHJQIXgs3HrXpecIVzsBaRDxelhzH0npYtgqSQx0HZMVdvkA4+yh+ZvGs6f8O
4S+SaWlZJZRlgvHm969z2b73cHUPSPjpzlMoI5igRdmHc9ZivMIgmWgDM45X4ZhhUNsRD0JupUny
fthkMLjuVAYViqcMb3PukPAvT8m8hvFZRGJWVf+bhTMkvyTXAvCI2rC0pordBCCWna05mn39Yhk7
GptIFzbO3vNmtHq0JaK98sQegYY42l0x55SwPmWY4wi6XpIbN1C2xuNCnCOZw/klGBdxRtKl0SxH
Nxnq2gYHm6uYuOtIMht5I0rPljsWDI0Oid7P7YGmbGjLef/FxbZl69JhiZRqvJa3d8l03OPIVcxX
ydZkvgNQ7BMGJK1uc0RZqtOUWdyCRFo6qYpfxmI/WyKusm59uvMuX4vcKxfbvIDSFPm/jdFUyaxM
HZ8hLOoCGG2w350eVqRRjcTxwllgN6/K8e8MeZEfcJNJg4jlIxazKQRI1aqWMXw9Z6pUzBY4o9Hq
MNu9K5vpcDfywUeHtItaThYn3VkdN4CSmEPryFwinhUvJVwTriWmZY5um2saubSfywI3UQAhi+3G
ccNCo+HBcrVbqtv6lQNnDUWaR5oOjQ6AuS1amP0r074esuFiqr1ZzK5AAhzsZCBQ4OWU9urYE7T1
8TZ3kGGrdUxlUjT8iOILDNV1vXRPS90eHVcYmME7+er8b/rcgYkXy5S1SjJCDD2fkaT5MjeOajP2
Sk622yeM/vJLWvlDVYMOS0qxDdAiadb3/2vMyANsvbW17qjlM+chaEGwyEznMbJGCF6xj1A8uJG8
MmYiM2PsINThx5IS+Cb/GV0WG5m7x16N7wdECNGAAblt9IvUeqcAqT3D+z5xKuaRFpk4WclF0oO6
YzGbD1ofEigB+Kn7TYhnj3PhLEgI29JrYNjBpIxL1r4GxpJznAZPMbwH0Ey9w3WjhCSyg1UHYH6R
iNOb48NHhnWadDzZxP0HDz1XB8QghfMeLbRRoMO+vCVDI7D3I4FIe5qY8lUvo0BMwCQwqNjciijE
uPXgVPsJ2BY3V8WBsOUWYQgwgcBLKhpx43y9oYodpUBa/BI9K8DP1b8JELO1r8giZK9O5QRQEyWT
QrAqHCbDu60QFfNxGA2VVrhZ6k03NKwZ8aM7dhYCzKSJ7CgiCXEpsNqZD90if9+9rKGzwsUyoE4d
hpBC1FLR7TmYS9i1yeGnLqe7gcobm7Hu996LRT0M+o8loUc2g1iQoX9ger20CtgmHz4oVuhKv8ht
+1vVRfr4WHrxk9l/MtEfyPE2L+DdhubyOCn6g4lRa5v6C55GVWdWwo4yG4AX9Qqq8QETerOfA+8R
hwMwjymNPIvin0yCf5LvuDwWDWW+VYXt2lWKdkUnIzvNBm+QxuX26agshmHaD8iw9kfRVZnA4N/w
4wHM0G4ZbBPRv9qEiXtjlrHy6VOFmfSlwwbJdcFwFycs5fSl1RNLM/yetXUh0r4khxvPCsDmf6l2
PcZeKnCx6zYQXg5maX7z7Uz3xTOOcU4bKd+zzN3Gj/LaVpmDemqf9g8WaiiaIA3FGDFG6aj0jPgK
Qju2ObLn/G3/4iwoyJOeKW/yvXMYjBLxQ5jWceDxgIKt9iblDKmHt0m8CoaaQihYOZsFfrmDcnQu
IjWdF9tg/Uqgnz990gc6yD24faZaOTOlYcPi4zUQigrQY1s6ONvcJ4d8W2Mv6YsWIx03YZxhP/QM
UNQ0uOrhLXSdrH9P2sn7O5fm2yPDlQcPDIC2Zve0Z8aNWhae3lTtVSVXSNpAOLZtbPdukBqj6iwE
TDs9Kz001uFwHeWorMP6yrZYasuIJyEP6Z6A+sRhUxylje+xnazEHAe5Broz2kLhA2r1L4KesL4h
bpHooiJeVhgElQT013IcrEj8DweSm3LKcFTcl5UNG4/cQiMNZ+7AZvSNjpcsb8paPYfO2bW3nfzL
0ejB64y4otKe+hiVhZzrT62DTTZXaUr7Ba/MkV5O75UA7XatOePRd0RZiQuhkOSQmuz0Lc7i+PAk
1xbD1+SDPFZlSIjXsgCCZcUlSjANTV+WMOFrdn73ZvtOJOWTi3BXWQSJSF+K6KfkLN4I+306tB8E
IiOtdP1fXDjffjApYhZ9PjDwIQJZg4bG6v6lYUL6mi9lHXSGNfGSRloquboJtdCFCvIRHPp2zX8p
ZecpLTHDCL2e4Z6WN0pbzNMC03pmGrxjSKLlbryKcM9eB1PTYuKeCVHFlimqaLuoP/KGqRea6a7m
DCOsDFIvXFr1dq+S1RYjJwf3YzFRW7+O4JDqke3Btsi0CBcWeme2uLdVVHjwJA0RGQMkOoIPHmlg
/tJmV2GLPufdhzmuWmyRFG0b6VFsqSPqBJ8doBhty66Y2+8HDept1zARWDovGCxi96qLrcpqd1Ki
/CteS9YaS3v0zQh8LzpXuaHmdFsutKd5PbWQeCADa0FkQOEol55jFGJr9QfeBMDVq2zh8QC72cd1
5PpNbvfTqPFUgJXB+xCNaPtVK46fMuonGKbs4HYbXqI9lOpHH6qgudg80v2yM0bghcy1eDZ6OyeX
dQbYPqH1taX1wOf7WuyQ8dBv28XA0/WMEqjSThTqIBJiclQJHol572wwimq59T3xhW4moUPhoI+2
qCpc+DCvLWAiGvxzMhczjCKwqbEA6AVPDjl3NN4Z8muNTU+iKbmAgpsMQo4LrDRzQL2Saq8TxE2V
fkkbvmJsteXUvo2OEPq9zW2QT+wu8IoR9EIm16KhTvGtNSbcXDtZeOITBTzgQnZLR++daP8kmvDb
EJ/YvopO3bAqGYiUPHb0TVZqRhwRhMU6NH1vTPy2Jz6eCXYFKIItIRNjJryrAI1DUNZrPQSDUq0P
o+36cSaoTT+Nc7gMDN/N9Gip8T94sZVOCiy38E8rMdOElcGaLcK0J/RfQd12uxmynNLHW5pQowri
hqRLNjrVdRi9BhU6KvoNR4QUBC8ZHBbkQOgpqWHB3SNounzM+voofcWIAonkXUYcgwhmOz8lZn3d
UjyZskbd4vPsM/nUw8z3Qc1rc7yBhCgwbCWxoPZJcAG7/6jUxQpNHlut53pfVdhp6MI8dQ1myFYR
UQCzi31YU6uHbS9YuO2Luo9BiQcqXh1ENmz0BV/pgE5+DUdf6jJxDQ6N06Gl3xjcAflMu2W3SyVB
6A9OHIvm2veaHZ5sC9X/+wSqSRyYl7mS7bKQ0nJ0FO3CCV9JfmwCyXHa3idUhjXiNpK8Pjkn/YpT
NuK49at9QCNxJl4y1BtPmrAi73wWiRp+nHaIfMZSXbzLqsk+kZwFnW1AEB2fGfD4B98YlHHNcgjN
1czz/CdRInmO1asrvmLBb1IvR0OW6sUelaUODYnJcM4ZBLYG2NsrT4IsBpijg5zS3HYXxk7RsI9O
bavhr2bRh2/uCM1LElTrwelx+GgSeP9ksC+o8Ke9sKkEyBYiZGCQd377WZqXcqXAVkzKbV9ZP8ie
gyNsrt2S4Y9B+gkIPBlyPAd8JEa3QECRz8iSCJzJ9NciHRaMNPEvJMevEYeeSCBIqCgRAgn5AL5E
PBUGZcP0G5OL73jyACh0cJN9+GC6ylnwdLj7SkB+hVB+ll5Gd0XfDbvi93b38rfVYsoyQUwHX4vZ
nnQFae7bQIy+VPjoqdRiiSLfz39FkuJlp9EzSiLeSUNF4Yzj6yTuxRD8L+8sHxTUFXlwPMQV9LxC
TOKN8bLaHyXWFPKWx++phTdsY5YZQtFTpJMeIpdKC/yZpngOtazMCTrS8Cov/5oogH/PkPFz75Ry
/StOwpxV8NHfGq30isnikJHOz/rM2wspv9Xjvpbg6DsdzdU3WaVPN6FlLn4WMde9C/GWZCqxznRd
evxG6GAPcVgynDiVb5EC60aDwlNTZLyA4Yiiu/KIOXjarxUiqgyUBRAAAN5j0i5lSZ/AFjPabc+b
OMUeGjT/FuIrd/yxFQ5WgyNHlSWVq1ZovfeI0piCOxXfvt6YPVm9RjUdU7fWy9h8wOlwDl0HIExN
/l0OpNcuwwTNRNtdL1HCYwE4AqzeS1sgRoqE1ZaoNAjW9XKNw3jJ5scQtQgO2jRe1aXvWiJ5y9vy
USdsXWLOyY10Gn8r7jm7ZMpNPkALPWSjxaNITKcokdZXbP79EZr6afHDDZZri8tXPKuCL12DuU0j
G0y+ly82Fr4r96TDs8S37uek0QfIZHAYVrlJM7PokjS9g2gCPn4gyvxt+1mJxcn7PWl9M/WSM8V/
B/8jzBc0+u1gTAEDf9PNIhegUc5uUNZ0DVkUKI8WPlyN+KkBRQZVuU0OY7lXQ98PutkcA917iB03
tJTy3OJENudO+5c1mY/a58gXnNwRmHysVU5QbY1XwU0Y34mvxJt5mT1uh3JjPIWPj5Lp/h6jaAnt
YiD+mXnXJlvQX0U10ktI9F5HEk/+CNKESzhrQIHnl092guBtnFGoCK9YCik+Ep+mRPCZy7Aa3U1P
v7caVP72DAkTAvPyOhFRu0Ga7xB6GR624990dunA05FVkEvpuGrNrNeMnbr+J7AzFBrJtz3NVdBQ
8PB1h93CMMJYZ3n2fZg3f8/QZFhNNiVE4byoAEsElCnwrh44DGHq7dKC10rlNmzTohGSDvobxyaM
Y27Sero8Io51qlXm5yhIRHgQk884Ll821sXLKm0a2c/E+eNzC3Z4VzVwXOYujUJpyTwJ/YkbhQnQ
rEP9lx/dxHFiAO+PEoipNFH1JkBPM9cGXazsnIXJN45OFpbK3Dah09R/X40VE4EO/GjWrRjas1cL
a+hxw0F6EsBuNwdf+PPiMCZZJKva6t2TuQHtfPYZazgmOk99aU4spNPwDE2Qpcxzm59pdwREJ7Sv
+4USLSWnpKMYX2SQ67fnGRtqQLeSrOS91AyqljIcgLRyOur4piDImeXBYD3oU5TP3yTFnUNHkIEe
Ipv9wUzsHbk0d+vVqF6WnNEjGNuW8n73J4NEdZmTYYhfGj18LPlJSkkMHMOYWwBTehfpiN8INhqu
hzzzWhmyBteDfbBXcdgF05v9YvyBa4cd+aZfYZEc6GvRNb2AJWswfAnRWlTfuGtwrBBEHOClcGOa
aFla2GB6X/XFcfDpmymkZiL9RyFuJ4Dc2fYdGXlYPg9wWjajUMIWVsQaWeENhKlyu/IDQQCUHqBs
gFSWkNc2E9TZXy+z5hgXwGkjIKDmyDrmLe22uaQpdXkihWdyDyuqpXUlAOKTtbASXjmKbPkPcH7w
yYOzAQ2qDqRPJYH7HCdoAWBCF9m2iX1vKWQ0eeovxPhuGAUAddDyY7ux5niw+hBWv5rYlOGnrab7
+i2PgUoC2nZJ+QAv3fSTEliL8OALl/kgem0xgHtdliIZ+Z7zANLy2mW8bIEiKl57ITcbstbBxidC
eu+nln0p6vvP00pNUhnXtkkq+7TdcM83Z65nZ+xoKowBB+K77QdPWPKA/6Si5WLwCXMp0IWGtx8X
KSxp+SBNUgvg6bpmc5NU9EnCHqVUr3JQom7Tsbdc2cN0XOPNgUWlezuH19hgyJO+zkxytOYbTIqE
5NTrKbVrA6z5YWZIm15fz4iB/ihDbnZn+Kq4ZeLAtGl/T9IaPbSFBiyvL9XOqE/PnGHZgf02Dqpd
BZaunpB89wz6ZZn6Xc7diWSS0RID2pUz4ehVkXKQ7R0OBrj+jxUFI6jdfLfL80Loy28yujsAjsKp
HnuVEquavn9ymvAlms1iLMXUT0bIcshwEWNU0vUMQPtpJ3OgRNRnhFVOSBUlVNj4vqpTvqJI22qu
HXuH9BinIoFeK3wsFdtJKKN2SWBJIoYJPP+ZaTgj7Q/w17X80EMftK7EbAiEjP81zdxI5UB/FQ7x
hodIvHgTqlOk3A5GaP8ayKRXwv1h0GTNvmcHvDxafZUobeVk4JUPe44BArHNCNCcwyESt/NnxRjG
VM6q2a4iWlg3Kn5sXw+w1j2kcqKZTIDqRH1txyzoQ3RTC8QKWJ11pOnuvwMN87pVqhBY7zES9cHb
n9nTLYkQJex3SZC1ckKvHNrB99nojUOdcFaOvwPFPZPUG6wbpTLkxuzJD98p+WhBohQz/BThJkhv
FQbwwNzw1AZPvVoMPcP879cKXDTmzVpSSjYFUXNaKGvxR2jimm3ZcyWQoSyO79IL3YQ6XzhAf5KT
uCWH9AscbLHQTYXTObZEi0PKi41+cPgh4PFeC0GfCRfsE4GhhV+rpBPt0zue+yyhP7I2idDxYa+l
ST8PKcV9oJNydQIPk/Q5NrHEmHPHpqIuyH70tA+5pWYPB3xlH3RAn0v0/kOds/y/D3E3mFeJp641
vfbHFPOteVGbznhBVDDqwdFTmwP5B2c+tKiih2hKPTe/1vEz4woW/+oMBzreJ36botS65lIAabyQ
ZyKwwg7s/zUO8hEPuEWqERO18hldELYRMUblgzy8m3nHuI7OBg+259R2ho9d5+RsWhhoIYZfeLyQ
BzpFqVdNR+hpORCLYPD8fpINy1iEOPW3Os+pjc+0tNBPJD106agbSQCww9XF+vPfxFItkNMUqbSY
x1AoXaourOWB0BQVs02dpoN8fjeH+ujFSr6wd4WKJJFb6m7smIeXOkIg4pq2qiMAPECq6XqGOOb4
+3jcjXy39vHF2XdgxKYHzLxVwM6XnQ7gT0VSRPbm1rL5/XwtGzQC+YzYGiahUpbAhwoySfmkzufh
vR94YtZBQhA7UUT2gskKRBok1zm0LKsSWfUitufL0QjrcKDCZeXPtETEvo3LmKDWI3DyKXY2neea
KO9OCVx3VnXX6VN/R5oA+Ifje1XtLFPlVSQyjTBPVaAC7s4YIcp7AuI5XKKrVVRvBZq1h0X8Iw0v
VJ7X3ipOpJ+n5JvjaCuqTznr1zMcv3oYqjs5ADRT/0xUTISMzajv6XJTmWHif2Knmbg0H//q0qR0
WhUEiIqdY23F8O6nI498gwv6tExGTnxWWD+NYzPvX/CsOZ1NvalWsQlrPv57xbwDwkDJpSSJpFSm
xNU0cP4TWESoOsrROBwi6L2695Z1TYWqO0a9gySXwzQy0/gpo1sONTY1n99TAk/9uFP020Mhjjb9
Ye2iCZN+bSoPSzH+1zAdZz4gXOz1wtfSGAOddkrys+5svnAOrRdVmYV3MOiGHDbWtdl/uE43fZ4L
ZP6XSIzI+egAnLJMIljfBrkyABvXXwoDlwmNL8ghLfgc1ECdnR2EfYxUuW70N2gNwlYGLr+YMVDc
OPQARRkfCqhnQiitYaOkpOzBNseAvae/B+eKAzkMpuKaH+Zh9+G/uP+BRdCukjBVFp1xFfH4FjCh
4Q9GzuopYOJ7SAO5LXKhc8UmKLVeM0+xaNBK1GXdR+qoEvBrZzRxPO0J05Fa0ffl9oSsCQpOsoWn
gDnr/Fz//lJ1iIDK49K9iDQlcgELcpbFhad5uFBT7B8zRYi9BxEQtsgyn8HjeAMOSOajqWWlTg5e
AVRlPA6O8RndF6kRcagjy4BLJG5ajmWFEVv0YlhzJmI5WeZrz1iS296DmQMDzmPOP42zy5ShJWM8
7wPiq40nAcjELts4EGNKCGiO8mbpCLNotzXqzZLfs7ZFDfY0ehrnoh38VgjknH4XKnStfLktI++K
i0cadfwuXYpf5wdi+ngj3K9Eh5vUX4fz+etJZlvr56Vlp7nRRdYfgYGRMzcnv27dROyBZ0EG5w6o
HUOf8O3d+5Axa1kAMp4Z8732RXS4PDF93HorNB/0NAclRWq9uBgsfwTh+31Ao1FBkCjGjEvGOyoi
CKg7VwxSsGkkC3ZA+2hUO2pFJcanJsl5YHdW17xzXdS0lZNKEy1BeqVhx5x5QNN2XkdDCZ+gj2nL
0Bh27wuaXNBIuMA/UG3j6o1weEYYzEtMRunn41IhBlh8Cwm8MSUVBNGIQ0Al2WqWyTgexA0GlRUS
EC1OtnmR8/NO97/l6mhnY9waseCj0uVbPgf37pgrp6/leqyYn4pe3RpC9fgatxYaG1Ub1bylc9aE
bXilsnYUgjhjveV7b9QCyGerff8KY+FHUqoMeCj88w0fSm2ReY9j09lsTDJga8pr7jYlZN9dHRBq
r2sQ7FQJFs5XMk5d3C49YKbBG5E6kUTY4cmsr6M7HwXHs+MEmOh8aYfh8CF7Z+OQ9rQZRPjBmLBU
4QYZg2kGtLaUo1enbogaVfyxSYm3ZVILsURNUSPtWMDHH2Kj5IptMTsevuoKFL9dy03OR4HbeB6Q
IQSre1AjYkKZBwUCkogrww+BvA7Z9pQTSGAfmHzTfsjRY61X9T13Gsh26XZorkbLKoWL02R8paBK
F3TlhRhGRI5VQWLOpGKSRIIe6fUDV0xktmigF5yjXHxnGNcFa6oWrPTuim0o3EDMt7X+AyANbvAr
iGAeOq0grsUtYvuU0h0IjGfleOsVXMotJ+vXwjgv6jz+iIzaOQQCHBukNUiPtFS1Xif1DiahANya
LYXIi3WY+aSakDmwV7fq9ACJ0c5w31IAZRYzIUq00eFuBsuZFK4wcXX6ElHbmKPZQP7qjp1l3f8E
MMqduEdJ3aruZommFsGzRrmi26GTrDmyA+Il3x34xm1pEmjyQHSB7oGbpcRB3od84ysjs+QBRT2a
OOU8aXXkUKVCJLpdrOzbBevPTj7kN42+oMkDBGd5KsKEcZx5rGlEKKqBmKvmgsJDM741sKK/0C7/
LhglpsMtrQpq0TaHC1Bike3MHBFZWbJbLIiDkNEJiGJBwaCS06HgiDC6anUA2dI1w2jPjUSdf0Wr
SYOy3Qh8uWNm1mEO1sNC5bPxlnOlYPbjyV9/w3SX9yhwiBPUSxbVLUj7Nhwyo/CqYyMmL0KsAYmC
gooqyFMXhpsJqCNhs5Btc2+CbYNyj/FRmOBPsbFx40bCrdcTSxXRb2wpNdD2rx9fRCBC6C1h1dua
wfBhcMGN31kBtDewo5UloZ6s4rqaWX0YkPRJ2bTWmWq4MUlcJkgjfPvakEMlseArDHX2B+u3PWJn
L8pQy9CeMratXmna7GY/Yi8IHFBUrwkrofTMVd8oPzCQG19oDE7FHNeKL1oZvbHS1xRx5ExOAo6M
nCMuBtLkK41wpi3v/lrNU4dkvbNqC4VnYD2ZJ0e2dpZRBqWkp8W89gcqEyr49iPtEsWv8hvNQ6BH
c3+SjIFt6x3EV4zd++1CaU7ULqV/kgFQUdCwsWM6wY62zn9Dml2kVEBnkQfVkjYMC56nyx8ZZU8y
STIUXvUcsKsWDkjdggpug1uAZOwYvwvMPjllcaOjH52Jonynz+Ieh4N4ceVFrnN0DTRdsZ/yFURQ
mxqwi+6jovnTfnwMKUW7LrMP0j3otibRNrNyS0NmsB2DpotBMCBzuo2hGR96xb7Bw57Ph0PCHaNZ
sEcRzLjTZy0eWNd+EtueELPArbE3psadmOZR0xI+d3YnDsXDzrUDwoDj1YCC/ObU0eFj1P6lHtMu
NRvbC/2dtHWsl+pKLZD6Qpo1gXZ+cKVT+h6QPFqgwUWd3/3c1ga25mCALF3Mu1drsT5oJxSfJWwg
RLPGw2d/7qND6X74UZp3xfri4RoGUxishqgNnGo98v5XY1xeZWQi/6oJtUmpnI944kIxPtA3TFPr
i4sYHjhfpFYEDds9Cwcln0ZaKmBnoSPdOYn2WPLvwDq4S2wxOdBG0xZd+JJp9pP1go9KqBbweFdZ
jEUBwwzl1shUTMM2OwvtwuYAt7BzkwAa2K6nOqBgrR43HP61q8I7SSt35eYpIlxu/Y80IpMGDQZ+
C4cwZ/Y8jbUMipyc95DcyBR5r0axxYPffOZJUDiQlRxIBv1Waf98B90GhBEDjLdaSBr7IsdGfNSz
qiZKk3ZTtOLSRGNjDkNClCyEww3tD4FFReTj7InnXuVRHItTN+YHJHyCKlhhI5MdcTNvsyu9KCtu
7xVkJdhPJmLh58utHYIO8pzViHzvQCymA9/ppESUbF7N8lG5U8+C3IYCpurt5g4ct2lE7w6qvbNg
rO6ymaWi8ybZGeGl3h3R5J1IwD+tCt+SIems8E/W6tt/sWeK+qTVy+uyyYUfwY7/7Nzk4msymJl+
HZKoHOOwZ0W9zVjxNaYmeXBujpbcXkcLUqQLHQ7HCTIWYXnMW8+La3R3M+7uOzUlxzSu8i3DgZ8m
3Qqnw51IMIgGzHagK6ubnKtLk3hhui+dyLXXNFTXW4B2ck7cCqzv3xUkm1GTbiYgTazEyfQRjulo
IMUTa+9pJ8KnncdMpdetSSpWz8oODWAIXNFpHU4lYz9yrdUOgztsGAOKQ1PDAkj/RPC1heEXuXoY
pVIhherJ9JhKirq/EB+up+efbN7YUasDfm8Ue/p0Oicz80ssvQRTayJDRHdxuqFNxwj0V+uzYIeh
RjTJL60A66Uj5Yx1WhWTwGDGa0VOa8KrSeAJBkww07iRxPo26gMs18cAR10FVgsHmfdfwVr78H2x
syz9pg5/22yeZx8sPjvr9zM3G4VNECTUy2NRSyE7o0OTf+BqhvB+jcjgnik7RRUn3tzwUk0NhKPR
wayAzMvgU7HnVb5BTDiu0jHrKyCl3WKc0r3UX2YDMseTluz9giVQnrVU/fd4Wx1iTijbEfGvpoaf
MGcqWKWoq5H/BLLMzatOe+kQF38/S5Z54HrTL5iemP+ZyMRu2j2bclVJUuJOyBOhwRwQV0nc+2kP
l9qiF1FVja4lg6JilJ/uj4S5JcB8ZkUwY/V+kCyqcrVZIwf/mjDFxqVmQTEq54Vlx13NcJic5yla
+XFruaAXkOc5komoohtxMzeyAo1+HM7zSeDoXRBm3pw2N6g7VRwcGa86rI9+0XpL0TjdY1VxNm7P
XobZMbP1jG5ReMF3HgvUJZcJ0bmXZXK7TLrrv4XCgtd1hUSfl3mis+kWzyFygFlBJXBFOIfNKH/H
uFp7aWvk5YpbiZMJSPOsG+ZHdC/x7bDU28v442n5QvK9TrQdWOBSxPUeTQAb3g7XQk8vD3YRJz8l
nbYKHsDhNpfDgFXfw/I2Ui7ejoKIopB/2trM1wV8i/5sS22HxCz7Xf3YJ/fs2OXb52u682Gm9ktm
ThjVMZgwVFBDWJsyWSxzavrAIQTi/MasknhW9Z3JPd5QH0my+EQi1Ef5C/gmTr6PTgP55LZIo4NM
Ye+F02fwgZ50rqPiaWPTUkTyJ/U192tioTx+MkKaSxe3rYeCpsymWmyYTECjuNARE+GxTixUV0ik
sA1fYLmdMLJvxQ3wODwqJCAtio/uXZu+7TzH0e2gXBk3Kw4efQ23cdEuRoFTMwh54FYp1Q4R9MkM
8ywqpmz/xwYW7ffddKcXpmbAXbG48ks2F+f+dv3B9zIMYg7OZxEprTgzL0i8LHpJtBzLZXLaTOW7
TOr3mwQFQr2Z4P7exLimvcRk0C8do3qm48jgUQaPnRIid7lyvdPlA79HvQ3w5jU8SaKDOCmcfrhQ
z0k9igZeF3FiQPId+4osVh6wU7xses0mz0A7dUqa0pqyPMmvYy/4nSlIl2S4d25fXmvL6NiX9f0K
L7h22q4JcHQbv/nYyyQKB7swQ+kNdmrnny8bmMG2bTEUbP7AtYqZK/VmxmxtJswzhO9lZkGMaxVh
0xio2wZJR2LnlX4Fctk0RxKA9diUuerHt2TjeWsOetQzeVbtrsWR23ba4kZ/Ae+pcpNB609gt/Pm
Vggjv+ZgXoXCUPsWrGlsm5oAq6GoogZnrqkrj12vf0EdeCOXXPeJT6NB3E6Qv3lz9bvqmHKvzTqC
aiqeEGK5rhSmQxEdlLiT84nRPkeHpEVUKzNXv2sAggXgatAQJQSugq/XeGaP7ZjQU1u4t4Fo9/wU
vqr5DSlE0PJEkfkHAc0lqEiKIpQCOamLqxCW6RGfBepd9trNOZsL2RO6JslKXz1mDaGITiNsdEHn
aHEyQURnFFeBFYiqOiAfqVCDioBrMXMjy88sjUGUSguy4rec8l45XoqZeu9QgESQKqdhkXT8LzHQ
Af94Wr/tgGSJEKaD5abo4VNPX9GyzqhmDVQ3SevJfcUBmexl0u0/iO5NASvz2riprnj2nnyQs8YK
pRNxiokowkLiE64tYYRUT4aikuRoQLM1tiKiLQYQTPrDz5FqiBuyAarVOOOfy8yDWrsgdemI0J75
85O7uRc2GpGSREiZvRiMHbIhuluPrTuyLaEmKE+7XTioC2r1X4h6FVUrTlaD+zWvT+wr8KMkBkdi
DeINZqK3uNmBX6Ljvs4S0+YLgfHxJAcGav05m7E5I860RkkAURew4GTyJLbJJV7d7464dqZlVzri
Ql1+WCnIg0CSPMWVCANU0LjPssy6N888wnNUiif3Vd7Z/W/cbNl0HcFjAGcIFYDz6anGrssYSBZk
zqZbGmPydXlbN8w7PwQ8EHk1TQXehJK5AAlIE0w5M3fEjIrWqn5CwHyRcwQd0uwxXhm6Frrjqiqu
kdr7eUD3vfFaecOrRazcnrmquZtBih2zNaQKfT8ekbxItDHhREkisOtBTyE2LVneciYjMWe36jaJ
76IXr/mDk0phmyliiZSs1R8ts96lb0413E3OJeURI84HNVrMOHbXh2lS9LTa9tQcQ5sY2Jy3qWnd
wFGZ6WGgCJc0UoLS6DyH3izSI3mNYYBrUsfJayzeJDsfr8/xh3tfn3tpG9u0hh+QS0QYzR2WFRnu
L7oSAkfQjiZG5ayCb14G7wb3LHCjkSqx/ELh/6rpH8oyBMljYjB3jCKHoE66B4bulUrJJIPNnzgb
7sU52CKZI2sJ5oX0iVHSlOUBFMmhpGrlj3Ucgv90djpcF6Qyp/53V7C9nsnBvg7RrxmmSFvefpfH
uV3TwwYw6m/M3b7xsmHalfGBVM+6DfqTAfcZoME3syTX4IuBob0lPQuqgkt2tQjLh9ASuPd+uezT
gSEqyQ++IuXb8AnSyFTi5OKA8vIeuZUtV3/i0GcUioTJnKelFoAJvIFtl4dON0TSViYDJsxIACwM
O/YPe3H97MD2nnvhkhi4qttlCcsjfE5lz+RbTXH0S12j/AYmUtlxEq/hF6f784XPmKpwSLJjbkaK
nsXKLfNVnEnZIXDqB0ISRFUJwdOgg7WiAj2OjvySEkcQDRxipUSrvPp8Gvprkr70DeHH6Vh6Kbvl
VWFx/pCxeF46coqMBJ6WxrpsJD4wiaQRJnA5FBT033NJ8JB+E2DeV8xXDTzVwu5mvBZVLO+Xo0Qy
bDq931J9ZlVHh2Dguh93BUpRsQa4jQrjGA7LKuafCU0iceEV5hlFVkXzIbuxg7UOpQ/LuNkHiTiP
ZpTKB3ClPEDqzhylHwX4itD3aIOJHpsytlzRzfbns66xV9EzgzkG4aUZ5ocwK0DJT/WLEPfifznP
d7qSNPSb8hV9PpLDC785uCG1sbwfyOWXRXi01BugOxHwdjnyH40nJLoFB0lWxoRnakGfhxWZDaaW
QQlRqY4prjyhLayTTbEDNpDzTYYfRpVAR6k4CEGKhOcPoE3+SBnYFNBkt2zJriRILFTbyXioK6pe
KrKIUqKNQW4WusaVqD2mQ2Q13geQaT499yPxjEfh/RAolpOO1DE0HwQjf83Ooxpq7FSw+qIl8qVH
wxvPZjtnf12krwnNWwwXxidop/jsewNzCr06Db9RtlNhKZy7z9dTdwygRHtZfZjazHxUDPia3iaR
BkaIDpjwXA/Y2YvI3DVevUyTtJE6HgIR5sWi8y0TbKgMyG5N35s1ymLRIzY/TTlRLzE2Tr/6nqbv
GkqBipy55XPpA4gI+CzKjZUKSAZfmJx2Iz8EcMk4VFypJMkeLZRc0tZodKF2eNWzu8KrY6sEShEr
kyuRjiRVHXvMmF3gXeCG7nHyWorL8yQRpI4tDu+FL1RXeb4VKNu8hJrgPBSjTiBslsRF4FYU7x4t
HUG7sP6Yb5SoUgdBkADAAVCojlWuGUACWrQvxymeDec2NXW99k6hyf5FP7V/3uZtZ5FbHw3r8ZMt
KO4XfiXB551BJsQrQEostPQi6Y6YA8phuKynRVbKOfohV3SIoVgILIJb3ckgtQgxxydK9iItH2NQ
kUen33iEAwGQw+8g5nl69/7tXcDuPljHegCGmqmEU57oXtwqHe3lvjLJ0cYcCMP3kTmplu7ZdlKT
nfEC+F/JGUlQDyO57telXghE8gsrJgszTxKFfJoIO5hxlabb4322JYHYZ2TbqfcBL6GlSbA937YM
ExMGsmC7Y1KpLxfH3CzNEzWdHDyIW5sNLbyFEnJqIi7N9clNS4o56Og8QfgfETJbPgE1xxQKE80V
x5g+ln3wHLFF7MWOafpKoRmGQ2zkYGAOh+rf9D2jBzF5xC+mMK02z1pg7PmGzeGaeL9+ru6IB2Vs
frzWWWYLcvNZAHxecniSm3AeqOBPBpAW4tGA1uyeqcHzZfu7W4A7yaJonmjUjpQxK+SCYcAgFb9W
zGph0JXVt3Aan0jnPtmLMnt3zhdvdDHr+QxnC27IhvSt6ok2a4NBftOk0PpSvZVVDunzGMKl4+3s
0/I7eGmEZS4F7yeZ/JJSa+XeMXoyh31yXx1Dhc0Rn+sjTmaJ1AlaG0SMRBaiZdFokDECF54IZuqn
FQg5qXrh34xCHTSIZuuGovSCFvlnX3NbfOTacEISvLv97WWaC3uqPgM7u36WJKiKycwPGAR/69eD
If/1ODqc5OBrflvNjJ/1xucQuB1Y41aHyqP8yZFyNT82L287UwEpNqqanBEGPpSVb9wZl5cgpQku
tAEaCA/st07LU1m5DCes6Ftu+YCe/Qh16Kb+q7OTF7BRyQKs6N5bWcxsT+yNHzDE06VF4kgdHkMA
bNnbZ6evbUUe1Mu6IyK3f6Z0Rpq2R8/rMs66JqyC7PwxXveXhjQG6ejp1vk17IIWV972u1HbWOTO
EqebuFFp4fgZJG4GdDikwZIZiceOBk/QNRjWISbSIy8diioUyoHdeAFnEaoHWyHrTHrnhf27t9W6
zf9j/qWvAZFrsKSn7jLfVWg1hzKXvD5dGHKcKIRmweaDbe+4XaCkPjMUge0KZE7Uf1iHHR3u/XFO
fmw2eFRUJ4H67UHKHQK5se76wm3jPg9XW5uYJTJnUmFauPdzB9UOSXzM/VAq9jMtkW/whuKcxAbd
mmC4h/rE5wKu9A==
`protect end_protected

