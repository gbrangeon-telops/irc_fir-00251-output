

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hezhI5arYh5Ll2LsYr9SKRVb8M09iAN2m4JSbciXeqmprOA6kAYKyNVYZrZl+7uJ9rCbSy2t8SS7
C18wuehlMQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iG3qoWxeKUs22C9+IygRgNw/Ob9GNJdHtLxrQAtYdMzP86eceFi53EP4Epvud6QFqZ+YCcJAJz6X
BiP6+zFZ6SCjFFuXw9pefFKNSIH8+q7UF5dPb1d06lbHzIZD+3mRDkhnSZjrqT/zLAUZb/IQ1Lbm
Z5oVMb2d2CoW5etMngE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lCcH3M3hshWBn3vT8V7Ds2ckpLb00IXg/NREvwDTgQ0x1n/TYrAfJvH7lJwH3QNYGbvde2S4oTtp
dxVz5eb3NKybz4CG1wYBC2N8cyfQblBGlezgCm3PFTB/fb7+0CJP6o+JNkedc2s49uA9zPZB2axM
QOZ+WiL1UDOqHRt1CYUPiwYxRC9z2R+kY3HwbNnbrtScHXOfjyqwc/ifFZR8DvMU1CEJYRjuFvoW
cH+V2gM6YyOHMcuZuaYjA16MxseT+50plqCZJKvjkYTDhSYcuZeDAun28dPbdfRu3AO52/Kq9gTu
MLy1G+7O2B+746vqe0NC8W62Tyb+rHxVnOWRgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NvvNy4fG+VCfM9NYumsm2clZ8IZDrJQ3Wi+cnwU6WbSkr/joDlB0ZRXsdo0mhVbkhlHdY0OhRpkR
3RYDWBuljULA6BTyF1sag+KB46HFjV7grhZmVLUbBkCWRKYz0xq7bDcNxf7s4evpI4rWpbAGWyJ9
TlfOT5npzM2PM090g2k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KN7EzciqITw/PNwj48fL1Z5o1AjZa3hMKXx25N37JjIMxkR/++b3PX0LoYvLH1v4MmFRO2F2HE6o
+A9StU1NJwej2oLxLD63NMJa+VjJBFCfkNayO25s8BHSFsZkhjc8mIC5S+PHU5t+p8zDOXzJvXOx
j/qM+zNzxFnZOpagckJWraMSJbbFjRIGq2RuUI6DTykdz7949XyxajpE+pE2TrgIaNudJhMJkV8s
PmKxeai9osJTVlAQyTdS+HOwcKIcXexlGTP+JSkiagntbBuHEhDR83LTtvkaJx0GY9b8oHB0RXsI
Jp2E0CkC4MgVpkaduxkwBZ7NjlyO6dFeIGiehA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35376)
`protect data_block
lmd2ETw47noblrZdq/6xzvbux0vUj0I2CFYsvBt1n6AOFSWjcRaQIQ0TS8s78HO2Xo2zFBRp+I8n
emq14NDEg7HxYoVtNsvuPDeK8UYJL24Vpo/KY+o32HcgsD9emPbzTgkp5e/gpnfxtfLb6JCZAZiK
kl+oTBtVDuzgT3EKuE2jYmgZaLBh1S6yXpEAKxMulh8/6sDXZ4ePCqjmy2iOxN4BnjTsTlTxyfK8
ZyO5Rv31CZlgh26O4FKBiaxeGua6w3JgsO4jBg0o7ofPFRD/xAdATRJxzsVwH5vWc01fAg5ttnzz
tlZqisF+9y9mUWStjmRgKxEU67gHbOMcx16by4UG5wggc3IipC4yOj8T4yr5HiWVAzjXSk+78dSD
OxNvWh+W6ds/naYcv3AoxzsOsODVgbqDWhY3QI07i7NqZ2ylwh4SeLYgqaBG4DOLnii2vEXg9UJ0
kfnLGCTCeJIOrhj2gZdOuplwnbiQ52HLmOW3niJJWEoD4FMCCVghmBiq9pU3dfsvKZAsZoPkCn6R
1zV1WnmwrUPGp9JnzSKJQ5aLl5RkWewN2ZZHkhBZv3HhQp9YpheRr3J0Qt+nfW5MpQxLaX+W/Ceb
J3yt2jG4/KglF/HSSo31SqJh/NJ7IXh+6weP5TD8vEVn+QYaSIo8RWrDrih7ALpgQ3PzO9u+I7Fb
M5lCzx80u4Yu0XJioCt0dqcXoY95fT+slz2ktq/I5FpXRKQijES7NuY55nv+QIwz3FZyZvgqUo7f
fDAVNKTdvgmJrlz2smCSyCxqezvXVSjGQUy6OfaF7RGKP5fsFWfwl6NyoH9vyjPvgtTlM5MiPb2a
W78t8FnuGZTI4VtpaLUc9woRduFhkQ/g/W/18R4E9+qIhmQ3bbr8NPPbDOP0pOecBd+pCvsUsZlQ
C4K9ThCLsIdRi9P+wgKlI0vnHqb5aspjIe8zlOdusVWMKNI2KLEHeYChJ4jNiJ6jtrVrR+cK2QfP
E/QnMkkHCwFlnguMGslooNmg27/R6fZpSHs70OzxzOd9pgyDV0uI2gUAh8vf64sef8ibW19eOWYo
nGYYPHBoJ2WCE2Bi56sKvhv5POiLlY5wQ2gHGZe4/w1FZiu3u2icL8wXu6LAUNCJlHxfDlF1LaGs
3mUSjvdoS9aLLij8YND+JafXASbDNHc/CbXbrO7PweD5fLEQCu31cL8et4qOBmRO0IbSt/yfbFXH
o51EwZP9LADajp6IO0S1UuFscLI5shMsurZTWuLDw/nPMiIuW1MXyO4zi8W9858OA+Qk9vda1vIy
DOD/a6gKxs2tt5omyGKl2IUuK6/6QdtjdFRxXRDZBQB1XrjRx8r3kQpW4e6Ko/LwR+femXuVmteR
Q3quRtbaKLFIkJD604ns3//kEV4ZCNO9dUw8iMG/VaLCkOw9yEOizJpjrzd2ctItnFB2ImrxdJ6b
8hLQDVIvb0Cw/uqWJebpljO22B3H0fI1GTusoEf9FiKUKBQldJym8xUW8HLsUF7Q447jEZR8So8b
uCu126Ajj0/QSTSeyQcugkpAoVJXFj9XdmMpWkeicgjGJCqXpaXmMwxY+JH80Z+TDqodyyCkYF8R
IuwxWdihv81NuwsNP7eYA8uPTYBEBMTqNQ1KMAq4Ro9BusNhshDk672tRvetwCmOQiQD1Cp/IQ8K
V2OLkgQ5rxqcMapcEHvTEUPCh/7j+/SiouHp6nQ5TpdalCSvn3HKm05P+osknig9uZYBrLBMkUl4
rc44uP3rMimhbA3nv1NrEnfeBxiasfU2d4kvavjd1ZOWjSLd12UxBF6TCJxuZ5YV20up36Gke8ig
wz7ArfpBTVvQIwD29qYij94Unmyc11GdWu79UdDnPFfiaQQYfKb8AXDr1XU1tJhUrubwzMVsEYen
6c4pCAyiPKRAAV6DYHefUKVDlSxWtPBHcir3dPCeJr3j2GR3KlX2RoUPfNk4whNV1uCyv2S9/crV
hRP+i/c3d54HMf2RS7A0P7Jl1zI3WvH8EvLvbOPLN1AZO/R5t5ODzB+jukBSC+BWt6ASmeeEq9zO
rlv6OwMVr896jLKNEvLdO0+Db3tKoGx421aN3xpYCmn+o526xMKTiQNCHfFFTTP3q7Ojgtf3V1Sw
HAmc2pr0r1mFwI3Qb3gt+N0KdGW+nBDJn3vsQhS5d/87sACkK0SSOo7Z/sjorIJ4RRLaW7sdvv9a
laurk65YXLBv+yAa4DeBc/u0WmT+RC3UCC+BmzUUbPZuQvncofgUPJv4btCz/xdm+8EbNdGSDyoV
OcQ+pOfn18ENx40oFY0g2FouP5XJQoBLgnAfBmr8IM4190AZ0is6TuRaPkt3SqOUYQPq/9ov590w
mAMlzZAUVHPvjRIBVQ0Qx55088vQsNb3RVpOLsowxWsFbqKlyNebvHVV7UQ8JSw6DGp9D+ZPBcR3
WO/DPMQD/WwurvVMCr0pYnHL18v0ocQegotoC/w8ohh9aDi5F61P6Su96CBXXBtxh3JNBFhqEmLa
vRgOQUlok83DuDibWVsL83OvdQaUCJDa6TzkSvPMLmy+XEm/YBmbZmv3bSTerf7TOSYa66nTR7px
1JLGym16iknEC52eW6vY2uSso9XHSWL0XbLcDxlsMhrSvRRGxrm+sEvRWV1YF794hNQC44ML4DEK
GBKc40jjMPMXJebuzuar/rm5Gho6ZZj+b37jNDbSfVZgW8qtNfp+qo+neDtVKg4Qy7iQLQAtbnX+
SBaB6fZ2nxbOXhdxKwsAdo0/FkzkK1m/A+mvR+jr3tjMPuYQ9AhS6WxLo3Lhw0dZELWbMmFvrMH5
Y55kYnSc3pf2VzTtJPX2j+AsoHf9P/ZPHb73/UZjkqa04SPwrJSbw1slIJI91WsMfSgnhn6ETf1J
QHzMT4OBaOCB/RBgUssA8ine2pggXh7vx1Vip9i6fwY4e7D7h4VFvmKw7DSbacnwRj9uUWRa8oa/
dwDaulZ41tu5+3JRCyTKPrpJorKSMgxdP42NzgJBPdAAeLAWdmW2eR6oI5n8fZSOwtUFaN5Bfsge
FhH0xJsFf9RfjHrNCmfwODnz5ZuHLpYTJKWjfFzIHrCkX+mGg7ohnw9qFoCQf8Z3bDxAvy9A+4fU
BDmr1JQOwUfz3pDYjkq+ATP8pyOYmKYRYLYeNLDSeZeeTjbm2DUCT5aHGq8RmHOE1x8o6dPjIE5O
A1h6U7GzZmWsQQSinZsX/DFowxzdKgybujSe1q043b0XyvjxaJX5RRBHeLOX/aZkCHhXZ2V2nwfw
qBbMsIRsW58oD77VOhCv7JKNuuIxbpbWdW3g1egZgI8wYjy8YHp672oYpfGhddfIJmJuxLnOPxql
7VPudE98dq1hHTNi5P/fHzSRGD3LKa0EaPxeIYzU0qvkR833Ag6O2VlKNf22D5c+kGkKb45O5c77
j8eVlRZwyfHpxKjuQUcEgvdjrIxOiaB0YFnWg1LFs52yGeACEp3OOvEcUyWWOpjHxse+KjTPhDn/
4t8pDFXdvjA8BtKpJlxraNCDBBs/mQoi5VDEwABu+oGrS/uYRv5KSS2zt2vplKn7aufFNTZtwAG8
W9MchON4ZJZc4wdDJsxI3TMo5bj4kw+fczu+yqu2NoHbD2pgPbh71WTk3ICByy/zMmUHiEct4Mdo
e4nE4higfdMwL7hDSxwMBEwpgMc3YE53/6wWhHjkK8qWimKY2YfURWyCxf4FrlQV0uc0zkgx3wd2
DON8bE7liOnuTZ1R9RXf8kNa3lsAeey9GW5fugj3JND8J31qfQQ0T7Ca7n+unOlyyPKP4xvSc9vD
qb6T53JlGzL0YYNjQAorTFIFfbeDerX7/UUsrRfzEWNnhWvh/ROTOn2o4KpgAxPLRLnldhtenJEV
0s0aM44soP3QH4jToM3FNTdkKTVl6rVvPCeHmp0ZdimmUzdY+S3jknRxUAtBo8VmGla72OcwDMqR
O2F59lJGV/kGv8+E/zKOq2VoqxELlB1Nzbm7COMhySqL02vShjO8bD6uSC1KsY9CoE8XtkyhBYds
Che1Ds49B2FmhNGoIiZdjFwotUyFHiJ4zzFofSNpDq9IwfksJut7cJ1TMNX04yn1Y+oc6aU46rby
nuBUjsZ40fndbw0Qc2A6avwLKjcT7imI0ntunRK7zOBd4LuWdaTEXBJ+OaGo7glxy0buSPKfTAL5
XY0gFPtouWdQAyHxSi7LxCSP1dS3fUc8iPvSgNLRJy8n7wpIPyYc+z7dqUVezm74lKv4tuRBO0Qd
fW+4d6ifDXWSQ1y8yVu9ayp+VD38XIyXJZgOWmlf/1a4bhslw6au8acVb4iQ7ZOvH1zY7nUTM3t3
Xs9DKMn452tYAgHY8UQYGNXuD9L55p1GDE5gjOrn2ZYd+1e4BTAip/+M0P6R9JGJ5LUpJHGpJnbj
GchpdS5j4HnksnHDRD9q4U3Kuam8ylm9a0htW6o558/tKoA5UaDGqfp6He3FKRqs6odcweopVhTP
aPTJeGOvr51dD6Zo/jn13qcFIpo+zvhZ3v85jvvbm7kMmwhRBQZHuakyDtPSft+sHrWrQk1Ohhna
bbUKA9gEYn16fw7GsGYgJD6TvX2npVGT0i0dDef79moqCqoQrK0fUChuMRMEuVFqQw+DMYoAGkfU
hXj/yWg4XoVVK4pVRMf4CXTEPfPaVwSvVnInHiNZcm76bXaD6jGSxMGjgtww2k8+v6m7IxJDF3bx
eN2Eir9BE7+HT1aE3w70Jdf5CWTl/bEH184xlk00DctB6+AkXpGJcg/CdR86uAWdQVj+qTcK/OKu
q8se+moaEoAVvAptMBxFmmMwpcqOA6khhm1XZ0eGDYZrmxi9+R9E5BS8sNEj+ApzVyLh3NXIlBLh
J8eQPhR0o0qO6TuSnDNXySr0jcNYPn3A+TF2qwTygrEmmwBK0jT++8ngZoez4H0yFDNlMLuklmtP
X6fLwZvDEqWWUXwJRmx1uTf16AkynvWs+mHN7/pw9puJcXRcDqqpHuzw6W/GzqnhI2n00fTRFmXl
dkAUGyMLVSSsap8qt9puQi2mJL7BXkYmRbbUM8EjoYE+jxFLLQHECZzgUHQbT/DawzKC2harxbFV
e0RlaB29i8dvV5gF44uyMZNWoo90sN2gCcDJkHwSCPNs9+UX239iHmjShm7MCi7e/oXX0P9B/gv3
dBPIgmPppjmheZAuaho5jcNvYvxNUGPXAnZ6S2/MmrOIo/9zueRJwM6pSn0GBXx1nfdnI4zdHEKU
Txl0aaa3IlmR+VzFGZDvjakXepRRtTFiueBmvGHTp+R68wtQynTWHJcfDxmntSSGynp1QUMpnurP
rDSsCobTLGv258XmEcAEQeVZRRg9+NPexa3RY5UW2wepIQmcSfvVJboVbFeQv5Elyttuc/WmMA8a
nayjCdzfjVhy6m+6UqXAvV4yWwY/9hR/Zg5AqeqgX2qAvaB30/fwEr6ajl6tFXmr1qWpo3QcoYx0
JN9tgcSpxZ2rqE58llxgHAdSXqgMnWkHIaZcDsnVH2QjF8G7mO1jv5EHE9wrgRwuh8JGWf3jIXAm
ejHNkPWEkfMgIFXxg6uJQFKtjY+FjOxvUm4dkg52XGoXNrbPjA6RDXIvGwQoCVnAg5T7DYhnRDcq
NM4pupSGfsLZidh6PvcgZHstpFO2NhwfxUR2CPC33vJAh2E524YIeMk1evgHfIMPHJXwu49GImii
zCrpJRc5hDbnT0VNJA6+XLK3Y2CaBanesqfKOYpnIValOcq7MOwMOzD7RKiIwGinuAW3nDR2IFhI
MX0q4gjx3KLfQudhJngcWg9lJyPExCv2VNk98uIugmUHHBJQ46apl3slo01kT29FooPiXh4LGhU5
sjv4URWuTm0UCwilkU9NjUYiAenClpYQ7y+iqjtcsh6aKEdfQWYRVtoTtOmjyOqUmIITMj9HxJhR
bvBI/TUKhm6AtqaXLxKXa8RpLmEqmtB9z/S0BLCR1c/WTpiDa5h3hHHKiwX+LDG6gG2ZjEmkpzXk
OInp0OidPIojgd69JvfGuo0unweBE1zkXj3FgfabFB0RvwV4RfYSnUNPibluegO5OycUuDrBupwo
X7L+kjo+ADc3aEoBSzR1tgoWG5kmKT4MdDpZzU9RPRmksSGPfqyFgddF/TAC+0uQ8uFC/lsQXkKQ
jh9riRuHYZfwnwpFYDhmPe3kik/W1kI3wmsnsEUgewtRnBogvsHklVwPrdnawEgSzhUqRft9z2Xb
VT7Fu6uzlp7iq9dOhPgmdASH3GhX1qUtpF1DWWjYGsK91lOxIdNsmKpi6NSl952FxE3S3gX6wnLZ
cUAH/fR1b3oXMXnDqWHtx7HOuv5boDsTrOUSCzSmRWMw6PC96g9aC9o/dJpwUlMtZO7QOOXVEKHH
/zhcxPQt3S/gqmHDa8ACzPGB5R1Se7i+XYuPp9TUW8Y2o2NIYqdI90cfVA+ovXWxFphmsNAo9/ru
ezGnLpIF6X88Vz3i/IFPBbxJpBdO/tXxE5mQWoQMNp3YZnEfHAt5zf5Mu2seu4CcBgdkmqh1kXRc
pjYZsd1CWtw5x5YCOz4Tm9czxHTCqQcgU2Rgaj9uG+zAtmC1tsfh5/WRPzWM/ufqHnFoiGtjfR76
sM6/751Ni2eybYhO6YlB+OtFtSd97+wxarzJMEp0kXPN3cami7gH6a4f0NCALzjde8KnOm0NY/qz
6FvrQ+ZnfmGpfv+HdxzOZcuOaWg68lsht0/Eyar78VSeWbBgVf2yzEMdctIxBjh4b4GdxpjtVz0e
wcuX9ViotUDf9S9goZvaaB+GjzXFer30osNA9PSzz2JznMbjIy2cE0ekBl9yawpMNq+TT4dCZT5F
IjWfODhCH5sPXsrN2G5KfhBVFEfyPS0M9lJbZtlpnGomuzHq8flQR/Jo36/Jz8ZibD+dy6km2eWH
age3L/q8/dWY1oE+HjuJQyxkE6PGcHQ2YMGz2zFin0BMRmP2tMH5tB+ObNwQm1K3PORK9XrZCt3G
bKVKyZIubG/QfIs6EY2OoUa0XzqnopJugkOeNAB95RmoYq+zFjYJR2AdoeOcsZwqjv5doNjOip6L
hJvT2/WsQkoJf/RITeoqwT3JtlUBr1eHpwPU5VCML8RpRIXoTwHqszt9XTcLHDkEan/TFNkc9KmY
fNXVdXdP1poST5VOm8UDFeTftpd1FA8It1MArWPfVAC1d+KF/qzF5llr6WuWO95j6Hc26gOXGqMU
KCBfcBZ57cCkjXOAZTF33og8f/LjYN6gkFxT7FYrPT5agswThP1iVzWlqOz9RbJS+M88lSfNoTx1
+gz197H72sPH/Yyb4Q2TgOW8qbkodIg3TXcVHIZ6z5vhVJ6uKNiCuuN5UBUwxbWPMWQRcEqa885S
+tKIGQCnPsdCevI/DNtjFfcuOC8Qbj+pIV90AKPhzJgYUCobecsSrFWZbZasSin1agJx0aZUzNP7
N5Cc53PAl1p7PW8Ptg5o0f94nQYLQNC8QNuIQNY00gAJXWLUhWf2ysX4bN/sj0124WR0wR4M9l0D
DDFZg2nhMaSfx09eMDc3UOKtzqqCBcP//sSbEUPCHKnMLb9Iuqh5JxIRR7Zuls40BOK9iQNdRa3I
5nar8Z6RW3MBu1B2Yd7FpA+Amm/YtR9MNMRp1uDx4QhZalual9/lvM9G0sw1VpL5Rihom8ECVhsD
G8zv+beABNoQVKnTPjEsjeyBhop/z0RfhP7WNM5jQQHk9CjxETPzhkFWFMtHAf1mvr1RWj+Ha+ND
XwXE7+f9MmRQeWoUmZnYOicuVOql62J02mWpD6eZxHa7nq0tilyefH5QYEp6Q6C7lid/0G77d55T
L6iSR6HYGNDf5DnP5dJT7HJB5UXehzQctSpMrTTOT4n+Jc2HdL2uE3Mg6nrgfZ/zhvZzRUk9G5qA
xMVO6TvHbqVVvARB5eIcRvroRYicgUJmeXL0+BCzHhWDpDNi5sbLOq1BpRIi0fRoFN3EGuCojqk0
3pb5d4PbVjHGki0mJ9Ta6RxSaqw/DdmdJNB9uja9OJ3atBn0fLl8CtY8M42sucabivzFqOWsYpHS
LvkE6/XIJaSTUCxd8tlC8k1Y5/fgVgYAv0UTpI2GlsQMfUp0MXzUnVmk/PtZKjKy3VaHTzbJEcOg
41/PLNzvgFZd5BiSBWMAaPoXWCXhGKivor3inp3ATVABGlUE7T9J+cvS8lLuIVrS4OF8lt4cHBra
JJQfVBoefk3Tn+K3yKnnTma89N5nEWclw7VPouCKyWEquJwLg+/wXuOdD+3fhqLQ+WwSPNvc/qii
ozmo+A6bXvJ8Fqib6UZPATnDI75f1ChBCsK4O7PkGK0AmKgpp5ISFDj5IZ5xy5UlnvMNSojWanOI
M1V/bbKHEfD0KtIvxH30d6zbd/UdrjsfDI1bKU3X5fuqJffh7h7NTbmnTy5JSBf6Efrxqwkjdq8K
UnKNvuOx960A/h6ckS6k14u56KVG5nErpc1OrLN7HgYnV1pHzMv9WI5PA0NWfBbVVIMDXDFqWzsW
9yH7eYod5iIW+ntqvQO9dXr62LMpzI3zjCFYwOBFBQDs9VsCqiGUWUVeO1dbe3GWwpY0IgAr7F5C
K/yLjYjAZZDhT0urN5ld6QEOyo6vKKlHEnjGjo/tkUakQDYAjEh7fCDX+oj54l4u8YCaRiRgKO6M
mBgrRJ6viWi6pCdAWuf33OruBgh+VZzGSz/VGlrQz6+0ZAwhhmU0XFjPpE0iRZ/OWEx29gJUTnMb
VX8typbSUsw18RXzdY/xUm7PXqkgWqv76WYwVWVtwUTjr4pJ6rN6+IMGujQuL6MTUI34VRf8W4NE
nv5KnJPRAWdGOiuiv7qXzmFpsV2sQ6JtRkLHM1qsagkcWISCkpjHUsw6pqLGI6VXwUKmh+YDjp70
He51Di7MeSneQmYYla5STtltuK4AY50iUZOEB/+CJn49lPUtJOOI2nmUg+SobE8kz2srqwVbxlRa
FFfslKQ0nAD0Xl4WPvaTzwb2snZ0nEvLV4cz/LI+8QBKwfIkhI2Ly3w+qR0wGw2P89v/i7JNNJBM
GE5j+U41UBoqLKNxQUuXi9vdtzIfyA6SgLXGh8WFftrCejGYHpO3Qgdk3A94C6zOXX0Wf62CgVs/
ltr/j46CZsyjaj6vI0TT5H6XYQd0kXnPn2Y+MQZIRW2l9TKq2rrT5zv95JvZLhxe8FTiGdYk4QQe
hIocsc3+GMZOMvYWz8vxfcWoC2Ud7jMRReB/yz8tQ+Q0nUXrwRcSaeP9XlSJfITru1AG60crPNCB
ZQzyK+qnZ6hftgj6UceIKV/qEuvIpDzav5/duZRozOn4kWYDtaz2Ke48NrYolB4nqwIm82qIQIjf
LkiimeUd+pbrPd7j3XcHB4SQk1a1uWyrSWsdIAXEI/PndC2YuLIEnZNErmpI9LG8PKxvauQzxkAk
cQps84Kks8MUSOwd8940K47ZeUM1JQOSVB4EtzcJXWE2tIUFtTBp+gA5GnYM0+mx/tZsd5zmR1NW
g/npSeqYOKvYP6xTlTOG/eDiKkhW1v4eWOFlPo1gpuWlbCFtggqWG/I55sSG2o8Poypz7ETmxwoR
hJM3H/4pOEXr2usbyYqXK7Fj+nsK+kWXj9+M8j7OEnthLUtkGnv9rD9hAnbGSPyNFY3/44V4IRwo
kbtSggexz+bdLB0Y0lau759t66yiiYt6W0UUkX3UB8qvMHRcrcRfEzrQh494+LsI8Q086XFGrciG
l2FMz3MAG+1Y4/EeZCzzHl12wBKJmITYHFy2DgoHCeFTxrW3WJrJi5fQFEAXpjt07tfHulZUVZ3T
6my+49OByY38Dozl4wHUzdjAyM//JMOGjdjF0ZuVU4ElcbO4abfWF7gtZ7nyLRC8nRvVLiY+JXaI
b+gEEeLkW4fzrO+OyVhoqYiQL6gv0EzWTKyMy67b1uGRBfeAVBpjolwTZ+hjTnZXgkiZfv+Uekba
Q0PfLasZmmA0BZHwUvryuxd12sUY8PmGdWVQierNPV8gSdUH1G+v275C3GiPdqEI+YQtgA1tasnb
vaRt8kPoi783Y6JAIA7XsqB5z1XhQOBaFJ5vwGh8xfnFYnZLfrFHCz5q8Ok6W/3b6eMwK8FmeuSH
1y29pWyrM/6pJqfFJydz5/u6PA3+ex/3ECxUc5YD1eg+XfnqqmbumY8Td0zftx1Zz41b3pBNuzPQ
uonRj1Zl65JnGEK+m1tVDzJQ8lSexW+9jq+3OSC0akI3pgbwEP+BQiNeHysNAJTqcvpyKYhx/06B
e0DI8KbseACSJnPp60ayhgi5IOrzknGKHOgsofp7lypS/etJnFZrBg2mtc4+NBSsn1jQTRNr4mSL
JcOMu7/3qN2ZXkyS5rHD+2DpfvVBIhbjfbEDfEzI4ON4blnx45MONfL+YZ5D7zMcCp7n/gBx9CZy
gJr31K4c2w9BsEYbUpDHEi/Ge3k3c8Hb4ve1QEmkmrj9Jl9b7yYOoaY6ou6/QNncptoq7OTYCaS6
MKOlUq1fOM8osrd66zeZeEX0GQ+YoHNTHPnKG4jhTje5c0fdUef4buHNGsiOy27JKfeV2xN80n3x
0cvd49EfFSIe/9YU1IZBpr6Bb5ULHtKMvSM+VVZxS26T6/g4BGVaO6luH1bqSAG4ICtlLSQEJy7j
Z5GGQlQ0Eg8H6YJOJgd8aBxpZj6AEza8uY6gYb2yvcYcqazxah4gH/qwrdHXP9djveO3Tl0c8ryh
7k3DVK/eRRyd4i/ojpG8IcYaoVQf/9N7w0PpnyPs2petZR573lSL5vjM1cOmSR6b06K/gS3K1WxA
DhB83G3B3l0gts1lyIsgu/n5pXHk2uG3uvzJFaP2KiQxBpWsQStAc+IJEdK727BnVytR6Ad3S7qY
NZTQQ4/jBjjU6N+oehN7blkRrO2rFHEYlOYkX1N5S82NAGomjNBXuNqc1jzvw5b9fGF5IM7MGBze
N9Pmzhl9Elpp4RFaySpR4ZLa1wgiSuJiuIdYcPn7aa+BcBaheG2HQYCd0af2WEFt26ZKTQWtgcep
+iFGYKlXONw+j0y589Kqf2XyCQu5B8wasXqZfSPfAgDEWmxx8kYOaX9+qX446cBQEEyzHgMUS2Kx
/3iS7ijAdHEax12+9FrLWc6ZiP/U5/Amhnvbj/tdh/Uh66IQe7gMKFIs0iQj2tWL3h5Jv+Ly6D3a
OzAh2gqoiKYG/Ta8MQiZwX6ai6fKZMMi6aIeoRCTFwbUinmQ6BWtkAvUItNZ53/tDfnD1iR5ibyS
eDfI7IesubDIkqrSLk214dUBph2GNiEFQ/3xFLO4MD1Fcq5woSt2oi2BExNCUxlFNLkV4axV4s4L
nVazYt8p0o8tnrr/w/ThlOD0dZdFrP218PHmwkBj+qlt8PUKVXM9rGFPqG2gGBz1tVeaXWvyoghU
tlPaJ0mvIHU1IJNxAPbza1+2EkE1F3PtiJB4CQE8xvGbqaYj2oTf+y31+Qqfrz3VxkWso4eVWz6K
0dNukThAdI+J6isaGemATfzk83MKic0umEKr4bisb97SGh2Xp6pLFRIbn/AYdASSUXyDJw1B9Sfg
KBbCAeiM2oMj7byfj/pHykVf0BWDdxR+Y7p+x2wDQg7h3o9VCH7nNF2SNDluFMZt2Eu1eCDO8dEo
pPSqO4limgHtBZUxnx4X9m7U4C8gon73ddQOVTUFjhDQfR7o6fbus4a33x7Bk3h//Gf03bmYx6WQ
6A7tF/7PgFaZUuSz4KXOSVsuiN5B9X8EKYE8tMdhUvOm7UwTTUATiDjLyXFZ2n5t21Bo6DIZ1DqL
wjq22xkwa2MPZlvbpW2ZGOf+E+9ZyGB/0WPw7wB4Fa/FYcffV6b9bxEu9KOEL/+ljgRHdOgYcpM2
nqBF5B+6u8O/OGhbTKb+FNMOxYCjA7i0tEsiYrdlpSoClY4HAGLHA07L5wl2lh9juFUBvbtTdw1V
dPStmP9qOtKtpko/goHPn8D07mR+FQ8uP3ZbHFlDFOyrufOmYQ1wh3nQ92kPvuDZvakAJnu2t8Tm
5XozXsBrRc0QeaXrpOibzHsbgwc6HMn6z/QI9uLYlk4ylI/cndMOb1vyaFZyPMNB8+Eke+7xCd28
sfcJedyhyXO7WDEybSN2QH49SHRoyEZZP0iFi+B1tbyWnvhdkTdGURq2GEPyvdxscq95HVlR9nQK
GCndz69FrAX3yDhso94BysQTwXcfVCLrbPm8/gmNWP8OoL1B7UsTfClHHsUiBr9pUF5qEpoXRr4X
AodLkxHXZ504vYCui+kIhzsiF/fdQR1sSqsVeP4+mSLNVkxDnTDzn7AGzcLEMQGqX5Wdui4A7kjZ
1euRlhq2tEEdeX76kYlgCeESOuRuah004Wd92kzcH2UjSyuL1Js8oGVP9umsIFuxDg4SiOsKUGZv
WZIb1loipT18TzCjqCRIzh30VjwWECxe5lRnkf62UDIzdl5iJnaWWdU1lBosjEvE6JQmjpKzFjnP
5GhlgN6OCiMLeMs4V1IwPtc4CpJ5NJotI72o+eDXrP1RC/7CpEMpbf08RaNh8EmCQQFa9k5OAyN/
uc0AVvSaJiI9HUGJaXXKUrdyrFLG/DlB5ZYqTn70ih3dYw4ZiL3bOUBsR/Q1PkJovS5IKi/yDS60
WfLHKAydxjMqbpAExaRTWHAXWwAuEn0/S3l5GnQEpyf2Bk3A60VntNkitlsMxcUJUwulvMUQyhLl
9y9YWE8n5HbQ4kvBBDJyRYh+5k3hqbs2Eilp/0FWGy9vjlPRg6i216H6BZO7//1gwlByYUDxtcK9
mzDaMSdY71+oZe3lRfUSIOcEo7z7c16A8hxhF10AHBvo0YbloIu86lbrHlMbhauNrgYT7ebVH5DK
TUKLisLUPBAb7RGE3tK/amNlLLQZ/tIJ0hlrLSNgCdkk9HQRw4u/D3ND1DLq50YGJAOGRMCt3VTD
UQX7wkBikmnxqzW1o8on4Ohll5CMSNiUaS3ROO51LnDzf9uwS9vQpfTsBfTtfc21Kz+mH+t/rOOm
+JtW8W89ZI4kXxRQJodZkJyOde2tO6uP+JHW0J3szRwvyWDaPulF6IM8un09nDavJUFhUX1ITarS
hg0z+92Feto1zWdQI7dYIRlgwb+cp5wGIiKqIEWlVI6FzMY7dGM6teJNY81VoGB0xOQ9YWjdgqyD
nF6HAQuGQPb9X2SKXOE2EbEAZUVHbLN4XjFqFwZULnfyKdPcYwYZzuw4WDSNO6nh+WfB+zxXBfxM
AXHL1bQ+nIy3CsqIIpHvUJyHBfbCfCj47gVL4tr4dc6gVeU9WjZiob4O22cur8RJuTTDiBB0a2ZR
ylvmVJtO0x6/+8wAYWk51RJr3Mvefo3E3EuQEunq05GqGMstIIOrK5cyGUx6ElN3gtXAdkc9z9g+
vI1KiUB4lKTWAlgDuYSlas/HGH7fiy7HUuUYBVnOeV4jDJyf55PkDtlgl83hLC3rzMmUUjLDK90L
A6STw+j6Fvxj7tQfln0lXVGrWs5GAppfRQkQVKDiXz/0kjdOcGGFUZ3AmU/UWhZeoft+pp4a+eoH
cxuB6OrLsndPccxKsDaBVOaJrsIrwbRu4VRgLkf3DMwA6oHV7uQiu8iRXjidYEGxbujyb1hd+4p+
vKcDZc9QvLQmVjAl6R9DF43PRq4Wy5OhOpEoJ8ys3vqr4MiPvVg2wPA8PW3qVmnARap7MJsT46xT
aKe19nA7Zw6bNlADRI3sgkCxlxzM2cIr1utaHZzreCpdxJ/yQfiuYWBuaIYyKn9zCOVg9WOL62yg
uY+umVBUaHB9kdOefTox0byvF0JihMXZJsPpkGQIhV/iL4vLyeBcB1HVknhDAjJQmKqOfuJvYrd6
Dk/1T6refmb3+yxq5rtJXb0NwLx3XqGYPpDe62ytPqfjMIwvxebZmce9wc3mcVhOJPL4vObpU3a4
voVwvba9wRigR9uZDAI0aO394deS4+ikCL8iHlA4913U8lKLfedAhkYuWbBWAyelFh3+3r/a7vyy
bvdCA8F6Ch4wsb7OuzdTp8x4isDIkfumNKmmfA8eoTQ5xgsa5au3EDZcspVNGPgghrc9rDY4Y2nB
fTp4IJywD9aDPK+64mqd+sW4mZ81+LCk0cOI3sqzYAYOSphBAmcgwCf+nsxpMXkqCRIUBQ2GiMT2
hsgFfgr2dBVrOtTqHuFzz6++f6ECR0it9cO1UZjpmycuh/5S8FuVzQKDd8PZeE7pVQg8ODtxZhSz
aSVJ4byhi9tYP3p57e4DAMZjXiqd61h+RgqF0kaweOejVGBiSfyK3idBNNIEsV4cUAVdbGJmoZuJ
r0r9za8SFztZ/M47XMhdR2zTPd0zdnmpOb5Eo0Fdj+hDKraYETEAuAkk6F3gP6bykq+RGtFmb5i0
7eEmYbIZSK07nIHdJSMH5N+Sy35Yt0/SV6WKIYfQj/9/ZrZLwJKDUrqBKAx9r0uR0fMY83hw/iSg
84h++H7442LWFFiygl5YiVBcLwYSi48KVitXJbViQQhyvzTXqUVUKQio5iaU7qGksY69IgUv9MVn
KcbaDRm2FfJWQF2iqPa0WeQDSYSfx4DKWujn8oINmsO7vMRBaax0bRIVsGESnTf547ifFLTfaWTs
5/4zQieqzcqtd9EOmpl8+fszJdtddKfI7R1PP6M/J0m/EGqtNdLiLQm8CWa3WXlHmXTxYeZp38Cc
tYZVGm6cxhmRcYoBU/Tb8sMcr6bALBxdRuNIoaBKGS4K8wdiBP216XRfLI31SLO1oQpBLHR7WeoP
UX7gzASDCMch2Qh6zXYzQojFSYm2z188jNh24gW51hhZE8UvE28bzJXyzxkVTGo28BPH4c+jTFxH
e3vo88xoviing5c8o3h49DDEz5tIKCORYGGAN+vrDKZ5TQOtchEGPidEHEA/f0gzTTb5hu9wpcCf
MzUCAP1uS2SoZSgFi/WeWM06TCaonxaaoMjSF6l9efy2PwN34+n2JbGrbca4A5m0Ylc3w9vAz4hG
hqbH6d48PAreMj0fwtFc2s2zNy8ilzYWa2cwF4FTD7D3/S9QWMVxqkUTWRuvW5qqKxtggwVFfXnz
eScuY0uoxwD2Uwth8MeVbAHFaPtsu9BdaehErskMGq+hThwKgufQ+2eNaLBezdXBaEGcJW1y4dVi
vTd9rRyuECEffu8iHgla1Vvmzw3GIiJ2Z+KysQsuG1TFsmY2Ei3ZK7dXpOXuSgi/nDjNENKI2uqR
UiOG8kUE1FCHImU8Bz3nMs2Wsxsd/9x0wDgkc6srC6atWsBov/rw7cbH9cKYDX2csJgiET6mKTdF
1kC1gugIVmpPJu+HrUuD/UOUDKaE19j0lZ9kSPd5D1mif5hT0sX7aeGYI85Q/69QssULFLaXOxTD
JuaNKiN7DYVNJMuJ9MHuXqWrheJ3PsmaxJi7Zs1dMl0RMUS24l6/LB4JBQr+FnZx4H8nXSAGmtZR
4W1k81/o8xEYnXf9ZXUUY042gUdE8pggFQlez5lSEt+4fThGZoiV3R69SR5vUwbB8D2pRyT/YObk
4s0x5mcHwc2uA3S2+CZAYOncwNSmsBz9emBf/XcYYOk/cTFk4v5zeSJMMcCnf0unr2m4ZMNKBTGD
irv73RWXHa5VwK+ROIDIQ7iQEYX9QLnhYT0StTQsLaswFlji/yGOZlYWSJJowI1qMUdyIs3Ap3TM
39S2sW2sEHq8/vOxI2Bj89zYKEwbfm7C/0dNx6IIlibR8WEs7jpWv+DZFo2+DYs99M8S94k/bBaK
Y/0MsedZDqgD7KwRvLxNSdmFjZTN9EXDB2JF4DB6iXU3ezhPfJT5s7W+On/kMopwedV1DaS/fhVG
j6sFxBzhf5j2tKOinwId2c4C4suXoz0+CQeiztiwgIqfeI9hf6dC8ujylwBchaQd5+pDW8I7tHdJ
0Lem9U/ATk4QrwRxWuKxepjd9F3GVy0FAeYP0cBLcGirELWFILrqHSigqzESfj9pp1Bj7H/eAoQD
jyx+3ToFZ6STFBBYSoJfIQt+4FXC/7VODhibwADS6kXknZ2otin4KFMkbhcQm7/NDzuiWMBvQgeU
xjnDE9d/6Iq0o8WqZ/hxYYmIan/4PjBLUsZiRhT84mHpUL1wcO20lMs1emX+HMV04NHVCacT+VBu
MSSkktRC3sKxiXZBWgJqYVF2r5svH6a7krZWQntGD4mOB42CA0D/EmIMTz9if5W+j99TLnPno8xB
odxbrIkL1A62yfOXoGZRVOtk/1cQKUSuBSDs5KXK+pmKgpLdFsKC+SQzjIDXLTilArI8vqZmxqIz
UG3yVACWJLjJXAsmopVhThl7XbQn6siaMZ6tlosPH8xMiHOmPoh5jtp58PBjgNt3uDH9Sj3AxVCy
kEo0JRjNzEx8HQzgnZpm67ScVBZOSwI9ffynBzJb4lUqaXrxYClKg7XXs6ZaFK6o8b870Bl9zQZ0
GuPrqioYADvrwCSpBXTDKgOPVONRuJTRCZLeEK05F86f0LDtWgEnMjJKcIxpXin3kXVzH+UgqotH
PQg3CBub4KNtu+xZfexYsU0e/eCT6hk0j5aCY9c08jduKcmgPGlMjNc0gaYUC8asH50aVzf6CZY0
u8Bh9pQk7VJAmhZ95V3QIeCBcfdfcGtw8rFojvqLrc390W9hdmK4K9eNHLDCJwQz3ceD4Ec2XttJ
YAV44Z5K+yrE4S9h44Wu7ltIf+4lDK6Ajt4i1fxpbpx6noHjDTarK3IJjZ7FLgafZbbcbTXLpTEc
uIuRrxhrMM3zE/I+YflXujYPF7D3w/WKl9qaYhhHNdeN4QB1dMCTSr8762lVlWnUEiuB338m2OL9
K9uKRGsaHAmTZj/H6NXmRqKA/i+Xv4zN+vMM3kogre/34InINrfh5abxoSHRZHNkfdDynwdgPKPL
GN7VJ+W1CAd4placTckHAxLs4GMg8KB1wGVd0ybVlfcF8jeLrsk8OUX8dzETicyEGIWJZxYkrMHQ
+amcv9axOE5TgQg1jlyqQ343+I8rfSPFgYXhfhgiVF4SXSbcXNz0MQY8GEOiCgLZhL0VBOlq/CcZ
ZjoVqTNGd4MBzgQnFffU+m8ANXeih5fg/DqHz3H42/aV4zAkq7jakfjIjCLiTKY3kSowNBFjwRBM
sHkAK/rsSHdceasQ5ArCfU6/vqkFLSi3B6C/pKjpwsyugm1YPMI2P3DeFCXQzmWukf3bcu19EC74
y6/9gdkdq2d6MaC5WirDFfPMI4POd4QOj2ka0NZUd95/JxEHGnmgiCo5vlieStxzjhmU0JeCL6DO
RlPBWmGzOej/Tbh5lf6xk2+Csq07ba6i4vtNGhfRgaUvQebt2mJHbXX2+atvsen3JYsvon3UU8ea
lBRdZtbfiwlT7vFMa0uX9sFOpjirdY6MyS0lgQRI/qRGTnsvdNPjkvm6MOHmN6w0ZdyowJ7xKfSg
cbfKZQcqDF+tJuSi4jtS0peH0Cjg/rbTbpPi+bPZPT/O/kHJOUZlsKAXzoIQ1gEOF9tHTGxYAsKU
KJriI1M21Ug0vhi10RDjdBeKwp8bYXl5rnVcwnNJmd3ZqA3JziHb9wvrS3j6G/YkM/LDGiKXoXYH
faMVIFLxOx4UoOiWwO04Z85EEQTneb6QApAJmeDPfbWJQImTe0eBOM5tNsapHftK0R0Nm4uIVY93
n7I7K4WDVGRftPoyh85pSPzIQRkogjzzaaIcTj7Kcau0DOMSLWZ6PMbZ7IqxhhDT/SiQ5U8G1x0G
SMDyZn+als8elj2ovhuM8BcUba6S1KTJGnLNL+zZjjpW3jWQ+PCQ6/zSI4EFUEyEbAHmTJ/V6zl6
vgeeA/jV6Qh2xUCjEUZwFxxg++PbXQkdNe4oo3QH4IFiGwAsrPWt9yW4V8ZaG1eCM9QZDo+65T7G
WkIwfG9AYL1r6F3OSlGEtqyYTVR7spKWPmCt2lfH2wHfBmLCaOaClZCCVTwMQ4HTzd99x907oli1
2+9qqlpoiI3Ai8DOSNsICJ+LXxWPA2yBKnHvuCbKOGm47yO/TcoS06Jgldxxo6d3+EUJWNW5S9d9
bnKqIVtQk9k6Ueikae2pOEz0aJvAM+RJ+qcBaNDIKFtEldYjADuckxxvckEP+Ps+qqM1K9o+7mA0
nN5wlxiWfXGN4oYrCGAgFDxDCjFGTG3Q0A9iXo9DRqVrz9pQUI35CbwIBygkmV3mmnvyr/9ejZ/4
m3BXkXtWJPvhpanfGtlB5+gYVew0VHD1L4OSzncAI0T7JzbBBznH2XKWjU8bvP6acg+qTc5fj3bH
oxH0Y1vWQI/iQLhLukdZRKfrSJP89XRf08QxrDfyyDp7mBpiGSmkjP4CpODnDbSoCwUxhXQ9uu9e
Y5ydYBmT9fxwSua+/U5Iy0UnypGdHxL9l3EmTp4+Ng8nLW4Si+R3iZYZv92AQCQa4wTUudJn9NpV
8zgREG+hfbR2V1IISRiOFMjZy/pc1niuQeZrHSDPV8m5BUvbTWXaslFImvZowTz/rDCj1pwqEwzP
F1i7lMILngoaMmdl8Kh+Q57QmqoMdiByJckAX+29IantqucEHRAtXDt0vIfoQTq2gH8CF1HhK6Ht
ix6cyxzZ58dmNqjqnEcUXzPvrFovwzXfwuf8MN2qTPka5QgHIdCG6O4LFjipGldiH+SFs42l3afl
O4mKxbGyNMTNK33/LxgBwK6isxjS95N3+6P+9qtHyj9u8uIGL+xgem30TYgeVL+txKZi661PgsTY
XMAaFUtPLWiSW2SsHG5KB+lI6HvKNIpEPPeD1qJQ0hOQ2GqM8Nlnep/7HvxKMYz7Ms6KQrUhbZfW
VGVSqw3xIwujvxjEJ/EU4Qie5KIa8TQJUmIGgKWD4d9psEsIdD9/6fC5UKFBfXf8LYvbtm9eJ6OM
ow2kaUs3ckQMUsXn6hgqUm8mEIxcOivK0ulRBnTCikcPCpK/e9sSHRUs21GHwG0mn8b8EY9CALwv
kdS2AtaPnqjKDmvZenFC7U8yuJCcWUPJXjbof5U9vFcIxAGENFFKmrTnm1fGkgzg8J6B+Heb4P/C
zaM7pioOefT13TObcPcb8RfxI6LItSVE7LyKb1xG33TBN1qinw4+i8FVChGUY3rc4fufKnU3oyH3
Z4ti/4Z7+WqR0a3uOvAcqrf2E4ZGHIDkwBAk1YxX2AgldHaV6R0qXwvJkBnr5ULlyuUAZ6DKNhQV
uusCcYpoKYCLAUadFbET9fJ1idIr5+h6JexmU1yq5cNGTsxSkDCDOaZmFJSsTGqZ2hU3l0Qgqm44
jaNKbvnjXjJC3NiSJ8D3WATA6Bevinv9kJ0tQrIDWaGsL/dYrYiBNQmP7kG1gcGAYXY1e8ZJDhG2
Q3wA+v4al6oWM6VvWWS0MccODIvGIH4nBVJGumq/VC7NimXTMislRkBw2YwYMQyquoeTphOhIonP
MkkcP0/pxbXFaZeGTEB7fxYGjxy2GSjFJemE98g5c86AxOotGaGPdnf9wsaZ42GqAVnRkOrsQS+J
7PfGmSJffcdJC/QSYd1qT7XTrVnIxpbDdd/+hzE4+/Lz1o0SGPStDsELhz6cIrVAzqDxqHFQ0Xk0
cHIkQA8Gs/tehps5AgQBvtyu0PRkD4Ukq5TFVXSFy3lTtT9UeFgitiaWJ8/rKUggXZ7J1pEkQSP8
TZoaDzbOwP/Ka6Dl++LajrJcW6iPNzp33w1cE0uU6+C3IlwPPhvQKmgMMO0q2ifGTrJeXx01hWQ0
TbOeXEH8A12kw0ZmVQKA0j+PDNV84jJ6H79dSlU4kWVVUsi5MSQoyKFzXF1q3AblV3v2GoTRePSb
qZuO1rRHwOwfNlGKY6GtjedLS5DIKgaZSd7RYwtPRiYO79uvHPCPJ+VBPdrmQhwC68f23N6Ec1v8
t9rheRAnUm5W4Xk/uORBdGDlKrnFnFG6uPL9wlgButy0OWP4EodOzl2XkNjQMLdG5qL1oPzUScuB
bdvgZQfkycNh5GKCwJ/TV+S/umn17urCMuZG6M0X5IJcGlqAUWztTDPyWwgWUFmG3LlQZGF4tWWI
j1ZexTjU6sI5hti7KygAdXdBtLiSpc1prK/scXjcKGjqvx6BSZHQ1EMddLgDeguMSJr2eZbKdWAX
f2vxANpFbLM+1XhNqJrVymCMBoo4oN15JEIoeI5MF1qSyw3ZjQKhZrdrA/EDpz0LIVoyif+iGOL6
1hS5ndYcZDS3W7pvXbFeuk6xYcELlkSLxnWe0OVAqReI6SmTd5lCGIzNA8NeoPMa8dnxtc+BiE0Q
B7T/xijwMXob3RkPCW795hd15ePTCGZNXu3Idm8aQfwRLPHpNNIlkizLVPXju15ZASxbO0F4Te3z
BA3ezW1wYYWuaF6bKXFgiiQLqJu1GtSe1MtgjJtA3Ji2E00oqxTsx2AsLxRLXOysXe3hEGNkgAZz
dmp7BdyNwZCJAhXsmVSyx5mkx9aJSUHqkFlhtc0MaDdtRPhX4ZS5LJP6HOMyGvXbkanQwXETB1z1
z/VmOy5rhhkY8STFe7KUegVTGmKDEsW15xtCBaXJt+opN7zTNhW/6U1g0l8RC8L8aB9nmokEty5+
2PyyEmqnjGI1urGWDx7lp60ztutecRs+i7ADmxCvELdPB53ITTRZgxNA0w+AqKjDeZqDKdsdFYZE
BqFe98IKMA/BY2zbXkhVlydLMm5Zil8UxBgpTS2mqnXm0yh85RwAzwrNC4TTo9TFUI4t6JcFN9a4
H7Urx94iLt3Ck03/wHclOA4Fre4TWVjoh7O9kaCugYAvhzM56ZxZ4SRqPqwUtjWGD6bC+1kFf8Ze
eXJBQjebQQcqKcddTWPk6Kh4ak58MWkmFwH1vqcOv+OhaQzaPPDl3/tUwDDnam+W6u6eyrSHd85V
QdtKS/YwPtsiEnYvWxzi063xCzy6HSfV938pksWMYCB+NlC6h5B/tyRy4m2DqNjBQiR3eKOdIsXn
T3nn4YvgosPzg6OiIOMJXr4w1dql8iqWpE2q4mm2mrCds817i6aZ7wJ60ej69/YRGw4IKF/TNzbC
VwpBGMHn6nksex8tOihnWHMTXVfk15nODcXhcP52g3bjTMrEuiplF8CcAA9wDUjt25x+LUfSmpv7
ovmyThpP+jwOdKEMlV+BO1T+9k02ZgcJZF2BcwZOcmytKIvpLiAaucTko9tTwxIu6O2sj+JRtJT4
KXSt3WfbU1a7gMSUPXoWev3+/RR/HTzmfIK4UbWG7LNKYJhW9kyN+zxPuGR00VyRbw1MbElG5/2l
ZOhuWyyrAl/dKjIKc/L13S2mgkWhP31rS5uKaq4u6SLg3Wu04hdmqhMbMkAL0QQfGRmDB5Mdwxxg
W39oBvgRfvd+ZkPL8eaDigdvu67ViQexuzAHht6B72VZrdNF0igbMIHz3TH+082xNTMb2GtehIve
PRvEKPSX29nNGUabEByEEw6mkiORo+8205XHeudos3l/8K3AjVUTGsO09Z4QrvUDj8J6XGXUs++/
N3bU8Zy/uuJlt91V22ydKn7BenyH9+zWVN3wG4gu3C3FrXnnTx6+rtZnvjmtBFyUUDnlkmlALdpQ
4UDjjiuR8D5EneiUC84bN24L7CP6Zlg6z/nT4QGuBqzr3q7NXSnuuMNmbZTDf4QxJrizNtVk5sDH
9ZwYueHrA0Fau74QpyNb7uCuJxe3qywe5gC8EIT8c1gV2jrXJb2n4BaJLYhWXMd2iB/whvo/N4eN
LTRBV5z4TXFFEfJjhQoaUaHARlUtFn0IfKX1HKasctThTX9QYx/EMdIBGZFeb0dBHOWZRp1ptes7
wPHqlJPEAzSsLvvIt4aNnCZGXzL0fXwYGmes1c9kYvqedNVgLG/nl6eWxiNcVs/8813TeRmI3svD
BBR8FcOtmjX3wo/1dw6GkpFlfgvExOoPvYs2ru8/dQlt6RON/kwA886NTjNQ9nQfn/cHtp3C6lih
ioXuFFes2djHFI2S1xre9hTeO7X4/uCYrimH+OlVNNAlIjvUICBqDjVeoHy5o8DgfQfAUGBEGocX
1Mg4PxUNIHTt7t+9JphV4alOJPpgRM2khZ8ETI+ZsYgie2hUQjHRcPwAqdE6dWTiuwhbZb/dAW4w
j9ZjxpG5DH/UBNotxmnSarHvgd2aeRMit0F78lLLJur/8CBqAjG9nPsAy3ulsPf8fNMi3q7ONffw
jBQR+slBf2L9hx6ad13gxkmHysh+w1tcIXYd33X48qhUNerZK2W9Jq5jpT9FmjvQkhY5g5khVC1G
1h2Z1Y9XBysoTIqU3LqmtLkbo6VNLYbpuxCWHktiTMfv4pfEJ4Bes/PQ7py7ursftLVgtIg7Q4mt
69QtL9YpZORXwei5wFAWFgG34+T6knWW+VJGz7A3AvLePTvH+tahzEhXVm5FqmQRUARHciMTVP9m
wXp2XjoYRtk0y9DBsV20RSaV/sFKfPxF6qcYH7i4yaFbh+StTY2B8BT3n/5BhrS44TMUvhUY4oZM
zQUJuujze7zv6gRkNKCUzQA7YiWGvCwIpTju0dAAMS3ss8KELt/C6Ue6+Td/gK2NOHxjKdZP4yqp
Zb+wI+h9oMZofeQNcQs9daPoZH7UleId0ym2wD6BzZhoEgTNlzWZTzT6A8l/jQ2LFeHMxfzE9cuw
0xvmTasXk7i6Nrj4a+JxKe/UCQSV1a4097xKLtVX3EbYeJObGJNdMMf4mhMYXUrH3ZU61hbrj2P1
VIsTirNjtXz+Qf6nJG5XodhmkZQDXC8o940dI75q1OIyqlawZQEXhUT37QDGxr7ahL7ZNw2BN1SL
y4f215uSxpEv7HvQ87FGC3V29zFXDRP1XcpRnUIuqgq8hcYaT4mgIM3knaUQopKaVfTFQGNuBlYK
moz0lGQtT2XyTMGaSfW8k4i8IQKhvwkz4eRUW6B6lPLWS710zRtppk4qOKf4mARV3wYhle9+YIXK
8B6twTT7rcoRyKMSzagP8AG4Vqd3WOQ9bhSoEyKwGorx/Ri4RTLd53odsAaVQyGGJNQVb//ZhnsV
UXDTvS3ueRHgFtYTKg0syHB8yYk4IrsMrAXbxVVaTSF568B95P67nQra8g178IhxWuKe9XHAp4AT
0uJ/yZ1UwOz/VCOUbQU2pzOQCy7W66h6jC6ie/STO/t6EFhhEQeXkdkutxaeB7dPbUL7E0dy8Yqv
2y/gXb7G2MoCh+HVAQJoLvY6utnNpLrjV/sgoIvdwAOQoQ1JZmf6DH3Mq5JtiCW23kSEb+Oy0jsR
gC0Wutc9fD3e3K5eDK57KjAvVefNISzipiO00zlZ+YxndRTdlMeCebjWm5bs+TlhBq/OCWvu9HVy
bVvS/hIUbpydCQ3WyuMqJSe2m/o9XSlVwUbD486rWHnslhRIo88aC2SthgpZ+U5KfBvj/IFitcan
UvzYZ7cohWovoOdHkxoMaPSSb3fh2iwJQeQf+vPKetWKCGit799MP6EIUiyQmU32A6sWGOq89RhA
E6OTCZBo+EuZ7Oiv87iKZAk09eoqj2iI2PUI2xPl7gJ6dqw1dGJ9wBBTSBmQLIpAJW3jpxjVCfTS
raVcT6HGyHQVgk3mnlCfMlQZplAJqReVbe6yif9JmxIW6jMVKej/uyu58zIAaxqUQGYx5JhABvKF
FOAH4SLQym+8EVhVbQ4WdS82fVQlGUIaCwwUGAGd7DPOPTzGpvUl8QpNjajIsv6xU2T6nvqHrT1R
XjISnMustGZdlRq2ZFVi+pnbQPJyHs8nRpQKNKMy+n5OG7ksVHUREnzMjDFfOzfOeVKlsPB9fKlg
AhtI/RV+Eo0StgLkBETNuS3GEIgUYzhIaGF0buKu7tOX1pE5ztrJnzpACfBXBk8jbhbakQRa8sbe
ahmaZad+jwaSLQWcewrZggS3Q6ecQg93eQ8EjA4ChHgh02jYLdx56HxDFZPeqNJTeYzff5N/8dg1
qcna/8bBzM+aCIrsQi4vv1npFN3Yo9/u//N+x+mSs10wrF19oLDItiod3L7LjLW+rCJTQk8rXmkd
eVfmPMWM2hZIFu/CXAREE3qZ8YEpjgKqmckv4dfqdl2jT45gm8vubGZPpjyFBpOrpt0432U/M9sx
+RV4DNnJm66MxvvCE96J+Y9PaWVji6Yq/8n+fQ095A3Af13+N6hOtRkiUBNJEp1/agYf94C7KdBd
iZn5JcPhzik2mKWw82aPlXKx5pC8xxIXYwKuTnoWDiIEKVXw0QQrwKMpafZCA6hdTUd7fXaOMVu2
97JjnIJli047rAgGKdgPkE/NsOa2ki1cKvQMs9ZBfY6KrIcilqid7AOf6zWCz/ZEDpiFYEVHtg2l
8wVqZaLL3lBAuZNhaNlNJ+9f8HJI2r2VQWifsmAadlL0Tu2Tw+hhd38gIETzL0amRd7DXezqPljj
9OZMPfRVViDUe6mkGxuvGI/cprT7aaZvDFQvlE02FK5SRHg2Bpn5dsx5lwBGI33fwJu0+fd3LXGN
MB1uIr/yWlfpLiE6R8VIKzQsmgnelatlNrd5OlQ2kruJu5quI16OfJFtz7EUaeOnlrJpIFI02nAW
n9F0TtbIXxBxSLsC45mGSQTZNTxf84qiRq8WPCks0ZhsVJjncO5LE3VVBfbh+Xyf/QHhe3H5BSKx
Kx4aOpAMihQIyXmJN8gYVDf0O76bVByCtqi9ixEM/ADlGiVnHsV5CZw0xv3D1QwADJEzI5qvlJnz
l+f2Ae2xYJMpFZc6GnBR5Hal/8CHoNAMcc45K4TXMgmoBP5cTYXsGY8Q+fqfbs2a+oseHTkjYMYL
wADftDfgiWCazJ//xbmNxxKKAiku/AFVsU+I3IGy3PxQ0/xCIqf+7Tt89EndwPDPTXPfm9O1jhmw
26bIja6q8St10p04CvPTrJgj4FtAxkE2VWpUWaAVcmwkfoF8hQSPsaDi7jSAQjquyqnhTMi155F7
BrNrap64SWA8t6UiVUmI2pBSmgwmRNuLtfXvcvTTGi/nJSBf/fiP2EuUhHnvnjQVOTLtIIm4pt/h
YFfJz7u+yXW+kRjSjFh3Pr3mIeZvy+AVgd7Z1B8/e0rBAzHnfkqNnXp/bswaVR79FLrFvfqD+TL4
7Fnt/GHYLjsLwqhuVgoqOrGhprSfsfg12Dny7lI/slzRbzbF9xinsnSRYScX/M2AlMTPmScm4eQx
UXm+oIEPSckFuitly2J9jwqI9/SwtqmFoxcHh0J5DgR4i97gG2heUQU4aiN3JFLOHoJkqv7B916n
VdC34TVPHCdKnWtjESmAv/d7JPp9C/LmoBOWX+3GhsPQU35lhmAorz0BIH7w+/nIfzlZ+T4JDFLv
niVUU8e9dr2vp7799ih8lcNM0yPgEkXuDsBXRe8TrJLO4N6EGqdp4u3JuoPhKEOT9RrUlC5ZT6MR
GpF9PxKDMp4vJLInD9tdZ5u9oPZy0+dDdKZx6/qhTv482dPqgSdGY0S3mBMGYUr1avT2jVV4C4+w
uOinDjV+cb7UexXnjLkma481M2Yj5yPm3TDvM+a5oW2LeI/BtWd73G1qt60K3fnwGqnCHmxFuKNU
w0fplLcVKeacWlLORdRaUMG3ui0yOu5Q0ePSPZFXEuI8ZrJnDkl77ZfDnraBfbBPNMmy52rGHdmX
yD4O+WUSjjYbA0g0dQrKwukvy1epB2mQAJXUIT36OkdYKj15W1FSQKGfS1ZKwgSFWt3mcxvcoFaU
ORrfp17KZ6/UhkPhr0WhbnFMjywNCkdkhrgXBIwE7WPCkiCPIXF0aeCHVROIFrPQvcL3Sn88kR1X
V15sQmS/251f/Oa+OmA+mEUs7RAy8gkpEhOLQUnRjfGNV5+U9SOFZr7rphnzsiamPlWYwkxJzCCF
n1bP04onkN8YIkL4hPOz+mSfKVWDPohxIqtIfTuVPOPs2RgV4Kp28D6ZEDh4ELhj9YP1ghtw37pW
ZnLzaRIgEQAYorqSvVnwG6xFh6dPCE8cN5DnJ39xWOrPcOHqUNpk33grwGbSIqvvAebc9CWq+/yZ
EfA5bBRTSZ+hSI7iXiJogD0r3pDfPrfiIaJuN+CYqa8FWvRAr5KxlTAjukMQaZBAv+FG3iCm1PAT
qlQqeLCYTTzQZM2NFpwt0rXa0x8OKC90qfQ7PyM3rdOOuxnNVdkaCVffjcAXXd9or/agexkVufb4
+G7xawB0sqaCQC47BLMNeV5nle3irtn0zQ4LjKKyCVhwn5bwmZ2DyFdEDwbRUky9DjZWxf1kaG4/
2cagLkjwGtggOv7qF2ohHMQOZJS0TfE2N9AK4rVP4QWJrs9W4jHQ7gIYxZOCqjoRPm2R6660dE2s
U6ME8hn9RC/u7tRoa9U+IrzzlGZIVP6OZ9ujCoAGGeKfeiYUPhOWRL8YN6qGmBQQ/htLOPxyDwsF
k43CDaLHVlzLy8n0QWGsiGTgm54G+j8XVn6kj2LbPcV7ItUgYGuXZ7d0qAz5FMxLDrp7GhyLcp3b
LJIJJmdL0V6RbRfCdzOjW7HLuQ/3Lg7X6Ww1yYikAPszaSaKDSQiX+nshr9/Nnmn+f5l6kbkz3ju
jFslbi8zp3CeHffCsJCAn0JVkIvSqm24aYTPGUMMJlMts2NLymd/VGKPn+6md8vPMV0yviLD0aFb
9pf0N+4o4QzIZcbh14uJb1l+Nq7zIDIuF0ktJqsMBhI3eHV9Y0AUNHlEVaN8VfiTqoML0YmWLqsP
lC76hjsxe+HoQxmEtJTWY+cdjtdxbDwuus7PSdcLBfJcTuwhnV/D/AF620Ud2lXc2YA6F50pn4dv
9Qp3qAPvbc0bN/hNodegD6/YU1NJpLtArXj2l7k/iwJ8HZcfaT920Uu/RCpFG4Me8EVfiR86/W0Y
TifAVoQ6l2AVPfJy1h8hs42MzVjDg1fq2TKdsMY0VGHXFLBhBZ4763WjnUBpdhFrHMHXxWKsIDur
QmUxbKr5UdfzAWWXKSiJ3Z1ViQwmlwuZyJb59j+jKIcC3+iryRvQ+lxxCYJwnwCsgFDpe4XgPG3X
XsOPufG0W1n9uUQLtMyuhMzPNopDO5YyHMz7tzC4AUHtOZuPkPEVwAPc3SrO8L8DVvbRYS+ZKeHx
Wk0rtOAO3lrq9B/MgHRpbR5rY/sX9DzjkXp+P2HyI8DB+ZAaeamAkDwHJzCtje6cArO81Zjr1Iln
XdTbDqqubIjlJBjtcVK2Fw7jsEZGBjr9DeorZjcCdEeMkaWHnmcKlxcqfAeCOoIQ1EYSsdmyr8B0
5L/DuFi7opTx9xxtuZXNhtphAZSeBjHIak1FKGYPShS2sWrC0a+QtoOufcwMZrOEugtDDbu2BC1G
V9WTUHHEUtl4lU9YiBLaCumrPMzjASCIVxljfS3JT9A1FIIbzdSWegBjEW+h7E7OvIU77CZjUTeG
iSk49qBlXeecBfMH69xyUvFxyDuPJOSV/5TjqhoC3ciHE+UHG8m0lRGJ7qPWIY6aq2DfyOm7QPFB
7jLYVdj4PnHFl8wQukylY0EImsNHOHQRASI1r9j+Jy6k9r+3rhYng6BD6Q2lTSn3TeBDGN+UzAib
qnA/zJRi+Zrb3Ka1zT5puWKCLT4fecVe8Z5/Xs6ZUvSw/5GyGnR0JsKDLRBksNlW9CbqBAlB0Jp8
JUSFY7T/XBrcsDdsAFBmcc54QGFd3Z/mzZp4urrmJ6O0o7V0KmbTlpWLRnTD3a7bDQVZ0EH74rWt
2WtW4ffDFN/RDmrPuaJqnPXthms64uM25eEtc0FCNq7qkuHqimVbsl1Bm5H906Db8YVodmMb5qcJ
clwUBljvRIsColp39Y/wEfw2f83OYd/AszVy/3kZkbxKidR3Lq9qeVRCE48pXoHP2TzRryLbetR7
4XyX1UHj+5FXEjMPFAr5KUA5P6Z6RXlfk/pCs7I0vsjodbtfVw8JZkvE/pMmAib0oQIKLThDoODE
zU6x6R29xffHuc6kfHDy/id2hmggtQZgv++Ty3dvi74YoI6AADs4DpQp1vxI6LnyN0EPDQDOt7Tg
rBgbMZSrCVV2F1jNTKRNfjF51ge3uFi5+pmfmc5flpi0VuovzcdEKP0rOTXO1VfVIYn2UQ6vI1b7
o/Xv7Gdu2HmZvrB61p7V4A79lbE+yB/+d2MQU21wgxV4b4qX6PO87Gl9NH3t67fzG1Cx2hd8j9ds
DNZLWMG30N6K2nHSJoW2cRzjID88H8FES5gP/b8zAJ9W2nO2PrFi9Lf74Tu/XDoryS/9VRRIoSV8
xC9lNygL1FP7+KJAIRhV1SfI4DZuIoxd4VYGaKoP0ztJnIldwaFsLbJ2t2kKwKV35gGtaV3245mM
PIjRbjalWcGjh9G86tdIgt+Z/7DJhlMJOwuL5IbsmueMtUeopA+9Uzbr/QOob0Ndy2Ec11UPI/MC
fMC051m+mq+nOwuWDOX/E78EYT2XXVsK3h2L9WcpjHHveBMozRGwi59LLselB14itJ0YazDGHj1m
ebCm2zpLXNDX/19az7JpafIDEASJtbzf13m0V6naDKzt1w4y85XOtfa7nfGpWn91aZkvvYK9Nkgj
DFZwBZuPKbn68kY7VOsRSD4qfZCNyq0u6dISvD7k8JOPJ27L/cLligQokBQNsHspLv5qNHm1xgRH
4gZCPyhakZnuh5wdhJyK3E4fx6sPSjwOkGWfLPirOhnP2vVgdlrXQwWDa8rbblio1BuxqURxs65G
iaTIM+84v9k3UVAKn8dRh0TFevQQnJLQrVNQwc7+o+g3gqvlljQ34fde/wKJOcOuEFJCma57oaXs
x7MVwzjmJ3/+KpwbsVdBJMnxaj9i69is0yNbN0x0pYMr2H/EjNv1MW74H01mHIeUwQOgITlzO6fO
dkjzhgwqoecrIumKwExpXVD7vLdwTYMAesnMHN/FRxmTW0Qubyvzx/RxlhCsp8aj4g/A+KQCYoEu
b6D4ADof55RTbxIhk/LMBC8V1ZJQ210oQHK4qcGdPlh6tBD7eUSeZ2Z1SNfZomEpNvo2GkrQw+UL
JK4rS9ZvIfKEGsTORb1tlvl3gCQnkmlSVyGa6ZRzyE96MhthP6HwxiRF8fPplBOllNi6fRjjXPC8
M5GkwX+Vo9v4kEnrePmGZwjU3LzABjXACV/xgxHmBATz/hAeAq2ZD+2D3Grqjvkhr1OzKZP9Lhl7
Y8JGwozR7jOOn3jDMZy8v6hHvTCp0Jr9kpznJ4r9GzcmisZ3WyAV3gA6kTGsBiuuP9X8hQItY6Y4
9HkM7cij8UpYl677sxOTZMVTvvD50OmY100MO9enIFhSGl8UWdbueI03hOkXqShk2mRfGQle7hXc
MIWEOaZ5edq8bhO5OaFVkk5xktk97obXrYo+OqktKhPscLD/3LkLCEl43cPrdo6bDGiynoGvbFPk
ImYR+HL4QOVByrCBvymQ5agUEfwcCu41LT4Z3u68X3slb4Eb3p+bhyN4iFbK6iZnEFDN0azRBr2n
uE7fyu43ZZwtW+rcDYLv8MSyV4goxS5A32ax1NgATtvQ7MoOpq5Qx8gsA+PGm5nIZkCYxhk5taAV
TUcdRwL1UrkV7b/qhlWMl/vQHT2p/5/V5W489fhGrh/hG6wJZy4H9Bt0qvgS4tX/Udu4UMypYm3f
6s2Zp2OylCbbYJO0EFPsp8JnZe7vJe8ds1EjdzVLTIQKf8smXPhrv9hgtPZELP2Q9HT0paxVCCGY
w/dwlKYk30zA16snNAavMTtTkb4oP6o1aXRIGkCTgJX+934M3hxnbiBIxapmv9yedKUdheu4gZj1
bEXcP57iCLBG6XJrcstkB4vklqrOfKz6Theg/hWlFbTefTL/dcXMC2yz+O3AnmWMxE9G9i2Fcr1o
YcDVJmIKNU6GLQEUT0QEut1uTG1pf9QBGMyipOwa42iTrx8nguYrARv+SB8DLN72mo6HdOdkAZ5Q
UVk3OW9gxVUUPyEMuLTIwB1RvkMVG3/Nly/icLR7H4efnBjNez6epZN9ZWDzqD+0JwTGo9G430AN
LFv1GuSBznUBmc+05SLb5FabaIBEf1NvREuC8/yY2WXZaL1qFjNnn9OJVerI7XEgg7mERbQa3csx
KIe/z7nsOjlUsmR9qmOUi/tGQk0l5tPdDZ+dquzZTE5Odj6NVD9VqJ/JnggfHTR1Naa3L8HJ1aVz
B6dX2ysa1SvgtZyKQt09VId2UjsYRr/oiAYXpFlhjq0CMsHBYfGC5/wARW23LSPYyzUH/3ftt+Ob
upvADt1cXodxR3ruLm6NzTvhY/SDHgNQCG/3IC2paicbTxSK5LvV5LyP4Q+PM+avDhl8iL13JJgq
8+jSLTzVR03sMcXQko1ezvFVPAY+qtyeFMyXyGFPqcgJZaZhTcU2s6zk6O4udSsJqwv/FF0f+Ydj
ZaBG3TQysgAIl3NtlkXOgdILazlpkNkiEcVmKJuycxMa0QqGycr+MkAwMklvdWnOnjjOYg+3olDH
QEq8rOJJUqGCUmq5w/DKfHaMD+ceiIMZRZxiz8fH0B+pbPYZkhqRUCoToDNvoRLizXAEruHnrZiQ
AE7I7akt0ACrvO62A2tMuADi0JB54MHszdLTC7RpuCPjbGQ1EKAqo93BV21q5FOJeDLtHNR5zufy
B43LO2FjglFYLd4sUXbYNaY9Q76I+oFOvuVy75z4enFJOOAKB82o8ImDcGZD9GTViDrnwOvhCebX
1yl/hZ3nqTu7Hhwn76KnTGLzBGD4/Cu0t6CJOvUWnJ+6Ks1/70FIIJhsybuYbWc3+oHi9g5BH8Ek
M1n/jPlmr0H66Ba6FKJt9NR4wNTzxkk6arjmNbgITvYFBVyUaqWYKIUSLavJF0xCOA5BvLoAtE/d
bCXRebHuX6zmKblM2+IZCtlEzul0Np2w2Q/jHcuDIvO+ywJlrKYQZwX6zGJFBmd0SkKpozr1xoxK
BgQ01/rjnCBo5mADMgDkKmk7JSWu9djUpzBOuNEp602iCpscIBvIWb0OJvG4wdgh2nInNekrUOFB
pm71Ylt/xGlfTkl5iqjWiA2PFf4jeb522b7gTaRVs68a5CM32q4i4kNkSP0nLlFOtUrnTAYp0SM3
MUvHHv1XbENcZXX5Xl8fnV8FclJHrebdtKIvvtDCywPL37iPy0+LV6IJt22i4LwNeOSRfcU9n5H7
otblQII4QMRi5lPkiDfA2ZRa0ZJc/U5ST7F411WrpfyhAhONRfPK8Q13BF92vl8EHPwNrNngX0cJ
DQegj0z3rZXtkTrbpjYRsTverjaxykMEj8MUHTJ/qlwId15+v3ICx9YnV3AeAp2zVGOsvsWCP51T
QcS5KsK9dBvTOGLxCXUX2WZl2UVXocQpI0f2szhls5yzeOd7iaYCdOsfwCcu+2UjiLe9TU9KoLdY
YcwAvgLNMjXVPfF4XpjQv5a/bq+P0MgdIZMCo5WlIqWQBDuN/IgrMoXfjBjxfBBzQOx2slzaIi59
8BbZLHI7tHh524GAhKzy6TYIUohZEkWKY1CXsHWTc9txkgXUjUf5QaLFkQcgO9kRIgrPXWf9gDAX
TLKAgfCsvn5SUxPnrKQKRSm1cogAFcET7HU7icj6XTrFzjHVD7l06uxVmiaNiWOQknHEwheJmj3K
QCzmX+3b+ocYdGAFTBxSSycqkqKTcQfLbcEwbQkcyKoSDSDaQzCyrxwGG6I1TRL0K6KhcDipRexP
+KILQ3+yncgbO7uUqfj/yMBWPkpovDNZoVqnRUnVeeKMLkgnHqRpge97o8BTAdbQpq1WOW8tpijA
XaFKqwbtnmUBslqDisc+N7qU1zIH4rT05ZZFgxrxIEfs11y1iyyDQaNr/rtqHaiZVfRWrkZtQ5W3
otSngrXyoQ+Gf5aI1DLreEeyT5jbsIdDaWxRp+ZgUONWhSeoTr3cS9Y4DFZ/ceWjJGnHzeu2gYRv
nxAe05WZAz7Qth63TwYzgp1hkY+uDh2+R2FhvoF6lOkE0NbJhg7n6FwHqtuHgHxs6ak1g0LIlXuH
WESTA2H4njaJaR4bKlkkCt15msC67ibpapNyNzY3xslpnDXi/c7GrEOCisLVp6eoom4JjhFyaSxi
2txjNxBJfMMYEWvmGxoyV0W/OVrnW7Ef/2Sa4BbQJ52M12UNEY1jOAL3FAsI2S/PHpFcROpZiS6B
5hVlBeLutYwBeAsTAjD39vXHMxm45utbupju45liN4lho4Jv5xaWOC4XVxQ69M4jg6HR8FkmDDdF
BSazfrMzy0pbZ54BQooPlB2JsN2cgC1Ukp8WQ3IT8xf4z5wxuLV9kpI/ynaJLS9399GUti6S7zop
Pe9hwi4UlZ/hFfelal2pzwkkvGltrCushpP0QZ3iZAW/9OtPAwCNELjid0r7/gHJ9JixwnDWehAw
oZ/jgy4/AtXNTn0DiYouM/1G7jzxqqwadWQsEPeo6WIJZgj3jAAraPVzcChFlfcDq5ePXC3lfIaB
+fMk27HfwOGwqjVxagOUGNj0lQrzCkIJg/W/wxbkRp75OPaQv6bdYZcWd6ny8Rmcz+O9xSSnlWnl
BLR3EdKaQty+wMzyY5Jl8OseoloCFg7qgrx4WaPdOgHKGo5IBZoAbBZu7xxoknvCh+ySz245D+xz
x61m0BxSlylRCFaZJb5Wu3BMEglG/vnrTi+9jNFJ5Djrm0VzyEYv4aozT+75P3RdwQlPjPh5PEhg
ox8QAfSFRrZw3/+Pb2PTbwEDbnT4q84Jr2l6iqtps1/ygPVEJa2b/LJv7xuhmmLabX/THSwD0NGD
97WnC+qIYQfuPcFdA3aIDTZn1ilvYGDCnHnyUPC3GB2zvvRv2rUs8H7M6gYVAb7K46lPhhaFTZUX
SwW7Qg55RvRp4BroCJv8xZkf7ECoN51fekAG/rRAG3rlqWW+FwJlvEh4JFmdNpU8upCGw10m13qe
CzUBWMJIP912kvtAaXRrLh0oelQS+lYnZJGm8kYyLrfqzN0AEUCnNrrbyYP8wFrx13RdqIpl+xhs
IrTROGGkaAskq2QUZLit7kgDAQrMqB85oGVOleNxyxwNn7+wPNaaF5gdsNrdz7XyEiDyMyVZRmeW
Fxw+JteWb+agC7sgOHUFj79QNjxZcxT5NXAaZyamQBHZdo6AyB4sWhmsMjc3L06EFbMC6qmmXKfL
VuM2+uBzBy1B63DTV+uGhrfsj8Bg2uLQqcqFnok6j0W8knvKUreFM4Poy4PLK2iM7wS+b3qU9zmJ
nUngL0Tnd3BPtSM0FuSvcrEmqGQEifLC1isqp/Fziz3zpJ3ANyGpw6L2p7yJ/6IJfzBVPkNJXZwP
TWdTyuuqyEKbbs7bR7Xlk9faWQBLMmlMGjBFbqh5BHQ5xOq4gTumPRh3aM0/WGSDsXNiCQOyOzCk
Gr5B2RWJ2GptZkLVnY1jdE0A5qRorvzQ88F3t3avGrKytnQeD870Df0BNB9v9M53pRWXVowrQHLn
dQRUDHUP50HIe0MLNiCAOz4ba8/9hI3/9yK7ZTjBKXDdSj5eU0+VYCxj1uRtx+tnM69TWGQTy8cR
QSeNN3DrGiG0AC3r452LYrMWKYIxa28OLDKsYOugfbJpyH5x4UbNu+W/b0vWs8YulMkuMOoP7dV6
hMsQ2kL09Cm1CbyNfKPA2kip2eG4fuHOQnkBlingMw4jYqvXM/TM0gWii9XUqv6Us8lfhcyQLzpY
iORZD5liO8eDGwgkPxrGZHaPyowa9qVFtntYC6ZgljOO25THZM+9WNQM68SSVik/gMKEY69JqCoE
b/vwYm4RwSOtZcxfbTBYgw1IZ1iWCtABOqRUNta9IkVjJH3ybwKd0M8lcdwAXB2TAs6z+mOZ57ip
JtlM7T/AcBoGr6RZM4gME8BkZSAnErId/UpGrmAd1n+op7MWS1jWbdxlaZ34KtTMaEI7POfWMybX
E8IFzFhLLbbOCimu7LUx0J9w4u+bSSji2K35JPmVdXVLK0Fl+fSDwQCWSiPtRtVIXGF2pRQsQ7oJ
WxI+BdxnAQeGokJz/UOlO3m8uWncVr3KJgtRSADSNUWG2DQTkoGiSYQcNeLVFh7naq4xe8RJ6jR5
ffa7/TjC3G+i9TDbMarvqgG5IE+iTRFoqbs7WNV4uxjrS66V18Fi0/CX4JBjO7v7PvxRSmCrm9pC
7+toCEt0KNp7nukug6l9tW6BA171sZULzECnDCbQCHZknlSv+LtHT4zJjw06MNm2UO96rt61JlSb
JQS7wEKheh+BWigm8wIrv8yilco3XqJd/YigkPEvGODpK7dGcbpzQqADMYKhUCr7QfTSMvANl04s
fk3fgo5CTEB+7BMJZWHndZ6CXZAXIzZ9FX/dO1We1+dvZeK0OYUzfxo3DPbrxa/bEZiD+IiYLvEJ
Mzde6PuR1t2Zodt4zP7o5RBDAcmKdF69r/XbqvDLNE/X9hzJmeCv+V/1gqC0zw6B76I5y7EDx3ra
4eHW2xkE5B9CjfpQ6dJFrZgATkdS6La2hiq4ljhJi/vEAgxvCQ0YvZfujkLLNu/Eg1cdvdRtgfBv
YAYqD9xMrt5HJyRQ9u6WIW+4lrIaQJaApNkJBLTgQMpJfvwUDU42wyRyEAY2LQGBvuQ306mk5mb+
zzNRhO7mevbbpGUXkiISIcgijscdVQq3FQ3TMT846MKlMVLF18gBipjJ+hiltLB53Kl8Y75Ac3LO
13yyeYrpkAsN229C3vblTfFDFAAEbsjNBGtIp/d7YyHeOIcfdf5nh3aodjMPYs23/6LJL+O7Bv2F
svjayn70343ivKwPfE0Vc89095GD9Gh9o9lbcr/VEolhsAs4dTMvgd4LprfT8c2GgTzTwXdzryr8
b63be5g5OyESsspEl7g082p90gw27bkvNqvjE0A1k2i2uikGX/K96YvHv+nhH9gkjoUCeat/PGdp
CanqckGQbnjhlP+fUREPqupRyH6Qd0v9G2pWtfJlZ7CeBCL6H/6MO/+XZCwTv9nzUBzMqjPHyx9w
Emy0kMpVv8wVGM7FzX/KjyFCs1A2It9F1HjzS0gn0QQ7KweT9TyocMMNpPiW6LEZDfjrLmIm+w3l
fTRiGiqyf9ICKXoM3pHZLQQB+HnvwGq0Wtk28+k1RxvvYvmEXkrEkpgL7O0gvRaSHkO59/sm3Bi1
Y0AgEnWI6BYd+fukJihUw61cEHkd0PdITJHKwiCrEilvSG2McdwGoPAs/LCeV51y7BwNgVZOf6kH
HROADy+cCFjMxH0FIa4vsvmhrWE9enefzukoGl0XmTjWwx0QZF5plKYVbmFW3MhmnKQN1+3J9sV1
lrDO5hjC4S5YjTlE3GiOCrcyWTMLCWNy90AbniUwsctztIveIY+WQdPKbkLF4el190GkXaPec6+G
9KfkexW3Btlje78oYenN54/SiRdcZ+zEOs/s6gQ9rjhMlDV19pCdV9d/T+qk9NalQ/ZaX/enjTHj
NPA39k7cAS26SlnHQG0oE50k240j7sDYu81sfw68nmNiYnjmpikiMrhSA8+pxdUxwBvwz0laXbI3
yp2lCBEfI7Nbrj5oo7a/kPqkL5yd2AYCXmMxjh03PWX3hb2L9TQ9BHr94qAhqjU6BuSoUK/sKrOk
ogV6xRh0lceM8gWDtu03aGHsjNCUz5ZwH9Ey6WNgQLJvExfdeoVcVfSxoYt3/YlIFjcrFTHsDVvn
0K7Y66e633bQ2NYq4X5BAkQFmDjYU9FxBb9GWK/HkWbat92Ju6I7W8xzZP1xJ4ZHzgfbiJpeJFKE
xZsncv2AKhBuXGZkCYeUpr0HbBJvNM5veBX//QN2mK5r40giSD/lcAEB9mg+wo7uDzebiYxHMkvc
ruZd7J04h3AtChJoGmQ+9HMc2YWXeWbdUW0KXM+wOrOGO+CQluehZ7ev8leHRsmqP1k5iwT0n6QX
tbn/4zHVdwu7YQ1AczlX7z2qXVhR6vsnMBYIPjV+82ilbGJzYg4ZzP83unEZCzvRp4g+eHlQDW20
qyVqriff0dHkmX/icsaKl4Pv/6tO71CN35AFD298zUZIeTrqF3gy6AsAge8Z7zQIL333Wip0CLAN
QtsQcXE7Q6TWcYVIJIFcpTXIuEvy5xuB9TIpJpTqGM3kKn9ASBPg+OKzB9spMeTOZhUE5kXYJ6g+
A6PED58lEbeZrnqeNj5EM3DZCCddGtty5apAMrtJNKu3jiuGFhssdSfrePjvuYIkpgf0Wu1D3tN2
iPayoCCDWKD8xk9vQb0/xkbFNBERIB7O805r4XzDzzBY+bNXLfC5Esof8AW0JkjyzduIomb0AgIi
JgGIHbArDDVkDTPlU9gW1QaLJ3bsr1qu59poNwgx3o/TPpku37cXXPYU9nc7543nAvNZTimhp6bJ
9uFzSAmYy/Fdek2K2ItaxUKst7EDePyXXPKDjUuoJkRzojhFDFzv5wZ2cRhz896cSssSqYTorhRJ
130defqi8FNxQltYLV0SvBWT+4EBktwZbbxL3uAqD4oZrFu0u73tUGtIjqhrDajQixJTmEEg9gK2
M+PcxAfHCos94mvsy/Y6rpmdF0SGjhmeJ9/dkBeZC+8xX6SVs9Lj1zoiKv7hCkVMeJ1CZuBSXKop
2Bxc3+/bfHnDKpG5P2ZdsbkeJ5eQ7Lhmtxdq+iIWqxj3Cvgr7InIy74ita4ZoOm/c+vUQv3fB+sF
BuO2a0gu1thv/Jutuq2vuv3uNZZ2VSECYms72LfoZxsGjk38BjCHTN4v2bugvJavP3VRU8Yk8zV+
eCiEVRGobfMFajP4+Sqv+K4IYazUhYZiqwPRUYKGWGexvriSKWRz0FpZmwYvOfEqfp7h9m3Ih2FJ
S1jJ+yUzp9pXJVqtxGmEMKpD75A/0uds0vB3bsn6gL7mIra6izfGicpGpc6Eb5ZF/2bvXEaKI+Rf
eUDpL1NwIZBXQkQ6SybSvLrPo0sH5k8+5bkY7uHTC1KLeTAI+e4nR5KjA8kg5foDeh9O6wgShZzb
/2HXSbi09bJMFnPX7SiXsxdWxleCDM9dC9BjSNVIJ5Nldg6/brrlPIkVGA3Sur6/wfAvyPxd2jFH
NwaWoqH0jt5iFdhqwxCGOxCXfhaZse8Se1AKRasxaMS8+pkC2bImDeVUnORhS6ratQA0I3JHgZGs
Fy6hDDY+XfRaM/T3K8c/ppaFTdM/hPaxClSG1p5rjx2Wpu94bW7tf+w2uhtpoCha8++WDLiZ5wGd
Tv48Ng+npKD3oatfl2xH2M3OOx7KqggREEFaC73bTMBULuHfRlHVyak6+IP3SDu/feL4mozP+pkQ
7Z8Ptjm6Pzqv5TYJ0v+W9m6YcS2nVmyyh3jSv1pfRLNHUjnlh+DPr38PF2y4lnGJobrNq/HVV3u3
zF7Yn4NsPbBYDQ31fMBSOfYmDoyi6Aq50hBnKp0B6pCOemkuCr5X9D4nNXs2/3pTGl/K9w9nAsG7
99VQ4HzGFtp3k2WSJic/7R8Wj/4ej5tziQAXaYSh6XeMkBQKv5q1mgQHjeHGC07+ClnuCTAkTISz
1kPgLgnXDR8BNuEi8HBjMjTNKdOHqQhNppmCNdq5OFYZ6xGd3wW5IBJGI5xZ+eBYL3OK6CsGt+9S
zfaMW25VQorgnza2fMWhDgjs4q0KnwjL0CB9zqz4hgoDYOLztzRK1tTTVk2GF02wWxxoqacXeLCo
9FIDLwscVgj8uN2Nnah0/0NECWkU03nWo8k58zfMcXP9PcDj92O2ovP+L1XZDtTrIilGN83+7UvY
MXDvjehoKfSa9pu6nbIWFpZBVBcOWnoVM87rDLPpqLJKhLzkmG00mn1XsL9bHfWys4UzqIUqocWG
OcSLIXt7tpEYPrexwNMQ2gaLa/6R95so/NHw1YRSyoQuGzm1a7uLpzIA2ws1xbLbIpyQ81AJ+pbq
j8mQddf5rAQcM8jKfMrKWDaDT2/ofprvYFw67q9Ft4Jpt7tzx6YzZ3Vl77LjdCoz5T1OHCh/re3U
o3TEATXJ4nV7g6VTu6x0Ivs24cir3mafb2yVKOmoq4lx1YWO40dxtTwQ+MM7fNgc0FOz3qhNiknW
0EoqBpp0UE10CGjWTrOQa9wpmp2hrnVyianhjSU5CvZjxXUsvko1fE9USmmZfQbBllHSlSrXQTR4
e9LPmMS4yDBr8B48YriaaAPlCgcSVxL6KnoA7H0UD0D+qet8g9MNzcTzr+08ent9ARwU4HfzU6yF
O92W1gYls41D3nvf7x8hqhlQnjpNVUE3+8GIrQEeE0osKYQx9ULLw7dHmQ2JTWGFB2o4ZocMe8pN
GvVY4H230dFq12kbhw5ogm67yxoiIrkBZ5jP6E5aiwrz+TuT63WDJjDW63MXJxZtyxWTaBKI3yzA
PORFKTJ3q4ugqXqTkfAOL4/HgkEJ16v1SF5zjyqrKyIyWhlxOggm/eRvqh/qN0aGKgh9dUb/RhhF
Hv6JyElQAeVBjqNzTYUeT77dl6b65wxAseMus4uLrbNue7xgGaYMCxI+BCRoHqx5XTye95dOBZ7D
sFBAfQ+X2X6/xsnl0C1Kq5QiwM6pAVfIvtXNc0Zq1IHfFWIA40rScA3VQm9lJ7Vacp1ej6k7BOoY
zQFZyObv2z8pw1GHWf8SXWcRR7biHH8/ZIH924TSMLHY3pdwyjGuiS03JygRDCxGuXMdqA3hzOkh
LoODCeOw28LLwJwdQAdv2SdIXNFXdes+1MyHjkWvcJJ1C4RXbm55ne1YCFeABEccnb2yKABwVxJE
/Dp9icaZ/RTjnYc4YGJzkg5TwkLyLwzBQOq4J8fxZYwNgt54qoSkYnDNyrgu6kApUDnQw4qQJkRF
nQt2eTyLK1Uoqy8ayzxQj+3OVMS4spKt+E5xrucW4ifhwj4cQEKIms4BRPzkcA/NYuRMVQozBvYG
EFTGg976Un0DykcY9OZe0gYuWAi/nkJVy/T/MMGzvuGVIXxvTkBHSSoCkQ1duV/0qxyGU4tnlHPu
DS9GSiQmn6WPA33o+HoASzwWC50Hd4hmJMXaILA1E3bvhEP1QvPOPqB23qLToO1uzv4v+tdcuucO
DlzZp4F3jJ9YSIVt6OnJ26z40i1Pv/d0zo/xpOVnnu/TPs3jjJAfYnrk3vSxFlTm/YFbXR8MTdsl
+zZ7MWF4n6qlL2nCKqap8K6HJ7+xlI55P7LwN0gob8noEI4sXEVd6wqx5ojqrjhFhWLfBS0JTOR1
tFKghlAjQ/TUwfOtfIrZt/Lh0myeRI1utAlldwEcgUR8ED9+gv5s06gqv6f/sUJc7d6eNutUZMFu
P0XTCdHoXucxECoNQdPKdpMfuS4eDqjyfhLOhC0cYbonf4zzne9pvd9Eusg7s9ezWTSKSHgs5i/D
KK0tS5niBn1hU0bpre0fj+gap5tVDisml7ZlVq9vkIbvLeZY3yLsrI0G8se6jyMN/vaW3ofevhQz
mGrV2ogEr3oujaN8y1ZIUGdjrAeCqoB1Q3Z98pLF6zYWoJmrFfpOdYPCGZexcLW5VvCW+1JjNhof
7/GAVp0FG4hSRc46aloLO5cnHcbsUpjtBbdxEIWBlLx+06e/j6wwIS/FaQvubnJwHpypmC0wpaFq
Zjfo51dDASWSUQ/Re5SvJPSnTlolo9BvK3YBWw8LdEuWye3mck+PdmW6aAk8tTgQwSOfgXKxl9B6
zmkmt64rr15e/RiHmFlm2VikIUyL+XA6ddJ3ai3WsonSHdxQGR/HJ/L3JLunE65qbHH0kOX7VwPS
Z+B7BWmxdea35XOQfQHnFAIk2ZXoqKLRkneTZ22GWXYEFBpxI5qHXixPfFkOlxbosqUNQWqOmWRz
MuYtEXdZDDvD3B5cAsiItFoiYs4EbutJsPvzT9ed9v/yG3a76T4bk1iJ1B/vyEuDOXNIiw1c89j+
2AT78Mrnv/8B8ZHujRGkGBs9Cwba9c82lyf73jmjrRCjWKXkUNF6MR6KoeN1zFcEDRYCOzgo8ag0
ND6P811dRv2nZwNGMRcAu/EadHHtsBtPkytL4AXA4HqSYy2+Qsnhel6m6K+wjvK3uWc6D3HuaWDk
6oRMY06z7gV5PXloVcVmVndMwcqeiOvnD/lMBvFWviKw+3+TmRZKfj3gfiYStvvuI2TFJah6wyGr
8afhH8aCSGFFcBHlFjuDsAMJniS1kmByrIa4rOx0lBjUQFpJ/Iip2Zqu3fYNXTrgHwsplGexlq22
7oHfrxPgx5h1waHF4tr/5x607MyfnCjra3o0+8Op7/+0QN1IRQ5sP8nD+L6MzfcBfrIt5d5YendY
kSKrmeMmbsDMM/FyR82v7Vn9Rw5nVuCu42n//aHTqDbbpaU+A+C1rirVRGvOMdpXkHFIY8PeQ7RZ
B28XtH2kHJFovE/aGVwA4KdT7pUVeVtiMWeI61zttdw5zGBg2jgRKkWrvXoxEZgep2R8tN7Yd2he
EGHff9Em8ztyRp3SWwL8EbFdx4HgBUJ7WAr+4HfM129zPndiRdHVtQSGzX/RiJbqLo7k9/Ui3YIy
xELger97i1Z+Q/tKamMdlsc7c+PUOVYdiv9pMIbLSrqWQ4rtiZwXK71cKjW+D68EtA1LwsUncYrS
vn2ZPR7UTE4yZCJd/UE5A+VlXP9lqxr+ZATuh8oO/5ppvLwHviNr+SkjAYhNFwdOUS7zrHw9+SJz
T8TZXaWi/+7xGPjeTrBqTSQvPkNO/chUFqTYebC8SfDNJakgjyyyAU9Bdxv2aEYFCIEg6KC96t2k
DAvVEGXu9C36UPtEE9kByvbN91aCfY5qFQaBsK6OTqGx6oJQK5DX5EmOYb/xlQB3Amo5ySgmBZb+
OIu1zqG2pOo4cgbkqh6GNvZEjGa1eJ9NfDop6yggzGEJydkGJLEWYlbPvl4DNirCM1NMP386A99C
0nsNINn5AtiGJFYWBlZUeZxEO/akAff8ocktTV2ViisAIjIbX9/t9Zk8eYX1oJgs7T8W5ycig26e
lKZWyfH0ysXOgnXtx1pH0L5pmv+Qz7JohLDGlQuZPNYD6W0pOAnN+xctw/Od3+QGUpLUotFAFnf6
GBhiWFJQ64zvbI6FLxEg1qsSzwEKFcA2Ke5Swx0gsfuL7FY3TatVBilxJ5M+rFh3pkZ0qTVldc00
IKhIuO7lqxhdXk1/5zB9suabq/p4v4G5+23BdY5jnA6oAMmq21HkONvgpfA3eoH1savEQAaaY2Yq
Jxw4Nta0jYIUjvb1ZdodDQNY4b4FMovcffCUotxIdD1MJJqLZ9gWowTRQMyAnPVx2rKIpcj5T5AH
s0AcD92r6TrNxuXCu3+12609F/F7HrhQiYyYI6w+nkTf7T7NSKFDA+DH2vJ0UDIT4pkqrVyRFloQ
aAgLtVLw4h9A1Q741g03GF5GSNIyH33RrvSzjNrU5IAb7eEUL3CVqkngl1q1z6ZpL/dH953Kxvqn
gqepoMmetCgyjCEVMb0TTNKHrEtXN18cGOciGKcn0Puj44F0vutaMVzyNPbdnabFkEvwXjivkl5V
jLGLG/EzHDet5u41ztygfYtt2SPmCSpw5qlMuXYR0M3u/VqJE6Cvun/c4Zre9FfrjxOCIy5lREO+
HfEXKZQVWvV7g1UiCqeJN8J3lo2VBAn8beVx70oLAVeeB7sCu9SADkHK1R57VT4u/sSeF0XWuzLx
Yh3u9GVMmjRCRXcEANcCO7Us8KdCR1Hwrd+FFRwrAkDIYCmdtu2ovGJ0SHZhFZGJ7dPJmxj0aQvV
7j0wic9ZuETYN/AKpgME32+acFfC3JLw7PoTGnkG8uEAiLaLnhVFZJK+1hOiL/iBfTwBy2Joi/NO
cpRcMR84MRBwuTqFXSEuLXF/biDNxanlUOEfSsXMYr4Hl5K5HnR1m/cFC/f4xYuB+HoaHnxRhsJT
QcwBNf72F/c97S3UAKiX9SK5dkUxT2O8JQx22+IBjwGzA6WX9LpzuoEmSxak1OQHQeoojGsuIwr5
ZigDnXMy/2xsnPJ5ToaINeeeqb8kyvB5R+YQRTRXJZH39A9JO9LMjMjM/l5hTS6XCECPJt4Q3Wek
7SegQwYjLiYi3afEKuf6zONL7OwQKgZCSrOiVttEXnA4nCp2NHa1Q8X+ob5dDrUvTcJL+xwYxaLK
1/MPgVdCHinHtIy9RRLZEPkaXbEYhHJsklTsDb7WjOxX09LZfTgNLkdfMJqk3jidup/ZQbhvATyo
AVfkbrGvsMn45q2d/s89LeE6+tfCWy7SNcI50q1QSTNb725H0hpnoJDV1LGHZcU6Y0VQ2Oz2KLN/
EdvdMOL86wpAt7B8F5COCxQAf6bM/2yfAMHi24+izUrWtU+07YFsVQKB0cGwvSEmivPCADL64v63
zrHJc8to1YuwW9xZOjxEGW1dfLty0VYSUhx7+hB1Gt9aanov+rKeFr0v4EIgRJQfxvajrVQsEG90
+AdQMbTmE/ApGND0N3Kr5clKZvvznGUjiOxwUft/EWm7pImWR6aq6/twgH7sF5gHVHJrY4JtnKee
zLbKNBF0UPFUXLno31+MRAuxaTI/f7e428khqBUYZ7zEQfnzTQe07VsZkFa1IbToOqGY8aorExef
JE4IPvwliBdSm7NSjAYZKBJu1oIEV+XCwn7jBcp5f8mFEuvyv0Hqb4j7pncOTdkd5JsAnWc6EyxI
jGB2iZ9L0ZA2Mx/7t/IRKK1n5D4DECK+plBWLYwa452/hgNCooUM3tHc2dn7eJdeILRADexg5yYb
M/W2Tx6jR97u6DkoEokFKy0SIeMqSDNI8QRGDxWIvvw1z3imFaiXSOHz1UfQF2oylxydc7AtYwgi
c1XKg1goU2JNJUwhujytwEDUl6fmV54FRqcxBfeCz2t8DJf7MkBC2Z/L7/nBjL+vACupUyY11xbl
+z9vIdxfbpCQK/NAWgd688lPu9ygl9ow9sO3JMnxTcOcbvQe+K7qZKXMcqStfWSgt1DLHJJT5IaA
N5NbAzoL90u1UPu+fkSc6RRSIaf61Rseh/sXEfl38fSGfkDRZkAN89CY8tNk15cr3UKdFzLWQCO3
dM5Nd3sWCJLropBs7CnWd9+lgzmvWY7lkFTo20uBaN4V1gQ954jb2h/ZngkOy5DlZ/vwDY+tiwXz
J8Xr4Fh7Yl/5QjvGslUajGq7GLCUlCS3MPh6rfRHwtayMY3hOr5K9S1iLk7Hp1BQo0rWcMZ+PD1Z
XRMFi/iChC5ldcfdd7HWXXIKW1eXNbQSBGIUnfLy73sQex3Be9k7YYG6fn6tW0+IpBG8L21ENWkh
3RXU2EoiUcwf8GQAK3sVlXTQDsbWEittqRWfo4BVWLZyW6bTHxSJA6/wVF2k7HLWei/TP+9HeiDZ
tBBQE4BAMKTvGGLQz7oNYr2HXZ163dZo0QP4yE9k0fQ6DyudDu5lcRJCDJJQ1L4UxVefk2zVJ7iW
uAGtBPqPAkHXhVMjILg7mpSXqbKjbEJWiA14+Wjqtg0pcM1dzirlEt+yUyotEE97o8DOK3LBrf1v
kYhKgDpX57LE12YZeTKTCq6ejXaff7eqxYS6FfCMyhhRnqpfhfYrpbKgvMDXebh199B070gMWBCc
Dfiw6ACk1+ajkOiTiQ52JXZPWMTAixJbtjLyuJwZoPxy2tUhjCnHjONp2NrrLCgKMF6wlRiZb0fz
FdojgEmCbZ/BRx697VQ3vHgzYbN2JDdSalWPrUXLdNyKqW8rHLJeBvCwwRfsYGY3kwgklszUr9/x
0mg62oSvlfSKeWaWRo2K93byKmLFtgg+psegnxvxrVZi7yLPiFXt43l+RUz8rqjPlJPP7cVNklIc
kYxv5WiJdek97CEHlhISxgI8ZMI/uhqnugC+E5DAFO3D5JVsRZtVex3+u48lRJYvpZDUf33vsxpS
gaiIqPKLHm28XxAMfDW9X1fcvkn4BZaPdKSopxGh/cvV+z87m26ButlNtrcrjDkFpw3AD3VS2QCk
aQJW/dyme26ve8tc/v8jvMN/tys1tHjouTcqCy84xb0pWUX3ve+nulH7QL9nQyLvX1hevjc4Bk3q
/sz+SUmHkpwYcGhU05bZ8RRs7uVwOVfe+KxJY0dgzzFO8mqCMKifwTk3Gf1Aj9I/WB0vSkKU0wTC
Dsea7+feAifWDTuIcaw1LVCd5I3p3MbgQhRVZSivmqHBqqC+ynxcvYDAnnwAZ3wwd5epreO+TBVJ
nRy80vELvGvPBdIdQEgRGGEf7cMQIhyOImWEmlwsxVB5NDIxnk7o4y0vVjzGkiMNSaOx7X83BxxO
ut/vI5avylBhJRXqnLiP0sIdr6PKTUxGoOKFzdnguf5PQFaZ9wSSGGEiGAEcvhbTdHo6XcEOIfaa
OYvkWFierT0e7d+Z2OrrEeA2bCMXonkJHHWYxZzeO3iZ9f/E11Wp8yRKDX7ZS1opW5x7zKCsrm+C
ubrrNV45D/dzIZ5bIMjccaZuo7OrfKOMLDfWFaOcuUcUiQl9tKmxcJfXpch5yg5t/Wk/Fk3jWcUi
HGvkMiEdVzPwmwdX12WdWQAgqH1HqKvkWB3+JX+XCLAjmIicCTDeFuVfbOSSRJSnK8nBP20WHS9V
t5648N41w2uFRWo4JKsOfRL5ezjg6o58eYf0ipHUQjg//75X5WF4w3azqP6T2S5QzGN1wdt1fM9T
BFwOzxi5RWjdeu+uXiuDfwET7qVjfczQR7VeeSBzWr3nLGX0uSA3mitg3tCIHbGr+VKIgLvQl8j3
1FaB+jjvSe6enPZwgOAie2knoVpVt2LEQ7RzIOI9s/tfIVht22dawGegfm01BXChO9niC8YE4Au4
f2DV7n2SNu0NKTjUz2/DLiJiigv55A5TrMwfcyoRy8lXPc7v5xvMnHwyiXWKQgDx7YNIdQeDnuEH
UEWD9sFrS0Z3cAG23/o6xZricSd2KYJnhkZ7MV7Ep4LfMUUou4Qc61xUOioEzcFE0xvKhmv3qVZX
MC4UskH59CnQUBNH00WNGOuLxYFesF70ptEGh48CTel6PgkEacDN40UU7rMp3Mqy4yz8G1p3ojSF
34+EGmVWdd1V11AE++HkLmx0xPhMGfhBllwITncCD7PvmvcE5hxydg2DUamfOWFx3jJ7IRGHZeQ4
oLhl4eMFoGdIPGLrhUPUVx8RtykiYGpIj7MM6k8YAI6gbKoiCiy0Q/O3fyysv01kqt5IWhP2lISd
dxOOPP3tc73/mEE7qlytQBIzkUVT3Vyy059AdfPAqbi9TOK6UzBrKk4E0do2beQ9vOemYHKP/z2t
jCQLEOj/DllPCgbHsEPoXCc2TX9Vvq+T6RGAHShsMp+OHetkuL3r0NybxyC8AYU5+kVS+csjRc3P
61UuxsA5OCQOkxZjI1TpYLDfveOc8W3oql25hgp3YexXefNVoD3Q5Bnvi3H9jkiX3Zso1z10NKeK
bM8VSSwKCLQWKDI7tTWysoJBlKa+MBvQYLghfaOZSAs7qrSL9ewXDjTAR8lMMR99iQL+/3g2AGcd
t4yyaf0T93YzI2Zzgu8MP6PCzhhri/7AEWm9vmxkcw3DHcx4FsUVBVqdEL1QLvjZ6g+x9dx4SVR+
vwqw7z/PeKqVxHFi3K9T7cQWw5y7guxZo1iYBQQ+Hh3peLSZ0CWCM/7OV8Mr2eC9gbTjihFgf9xN
2+A7i52FbfUeIbl1YJT2QWItg5JE9AzXq9y6IxOGtmOnjA8KCogYZx9rmogo7AH+Jq02NdiE5T0C
5YWvjfhcG80XbcUBRCK45jFLMxDNRK7WHUiXzBVIVil5uXB3UqBVxl5AHQwBUgXm5SilTEb6BWIg
9bP1bEC0SLDzBjBiDIPcoufasXtTsv6znDFqhJiQ2p5u1ptKu6b9dBZx3b/wVQmufH327uV8Z4Vt
Jvf7+bA1Neoxs2OIvSgy27QynbpkjBMvH+ArUHLhBNvz92QRM/bjeS2A6hE3sDC9TElO8IOI28Ur
33l0QyrGWVLFWFsb/6urhnwLXDyM+lBoMkRLGlnx2EG1ku/VF7TEleDlZAGBIPMBsOVvVBM1AWI3
oia2E1S0QkETrjt0of5gSvoS/8Pka/CY4DQANZHe7IJw5vUa0uI8LLZrDjp07D+yalCh7D+SnmM2
LrUZIaqOYkY850h7TQZXt7oChkihwmR0fX1xoIKD/xvPXZ5bGE2WWmiKMWSz56SZ6nsEH/RyWLee
o8sATsvyxaKW5yrcnb1Os5hGIQ7n3AVXzU3OCKpl84NzXq3Jp5voLiVztR3rR81TRcAha2TEsJ0t
yZnnSOPl17gViuN94sqcrmvZEWPl8oVXasw2F/k2nnhv0yxacqUeIBH7fQwplOpWcioocm45hU5b
3L+zk79yUJQySgbZeJxH6aWdcWeChDqa4Q7CULaTq0g7oEBch3RPBkkLIdbXdG0dpsMLRRRlUG25
pLtyJS4/WYyOdgUHuQvNfEXYXv18NbwYeMOiHqCL3rpFoU6xqF3VDUe/d0yUv2v8PI1WtZo5jLEO
w381ioXGjF4tzJpB3pAnq4Cm7VkVXYYlZ5wg85u59VYmnWosnKnq9TD2RgvWzZIrTCKsaO8nF6jy
FEtWZAQs34LE1daAM2fQMbcFeHth5LzhUfdpmcDDKj7l8fFcGowBxYX0SH+lRC4GBLu6XGE/DHnF
vd1uqM03ObIPw3JXDTI5bpJTA4eaybsMEThLTuha9kc6ZSmE9DgFrZCcjzklpT6YnUU14zUe9q9q
XJcfKJLSbYHTm0xfVK2bfYqxpOg0V/9TQ1IjXooqyMubSDUxQJqCivr+/nfPeshDACUHMmJkh/1S
YZTDBtjyAso4vOYkBfPhD9+73QkRhM84k/KNa0eCDjOcUOkZPW/qYnxJWcvoiejiREUOKIlogX6m
WIt6TW9b4vZEY1CaxUlcJFKm/nPIgl/NZylSR4fTp78K9NUlJ+AjhtVQUkAPfZ4NCT6O6PgzakZx
pg0AZBFH8JT4IUz/yduL3qrunhqWmSUjT3UuPB1vq2Lcq22g6I4upRyrJaVWYIPYfOxj0m9nmkWz
7RvGP4j2c1+KB0iPNuM34EEjBq/Lf4inHNSj+ezIOiEUOGaW4ePwKU7cjesr47v9uLxKlR6GFDG9
y/N0C0F3HPB5BUAmbX0D/eI52SVV7MppaI6A6j8Qmq7AG3bv/lt6hJCM/YjhDAz+PPQdGNTsYx5F
jsl1UFL6h9TEdZzGMPonJzds5exZ5gb4SKmbQW547rAk1GXAFwjYkurh3MDg/9LMWuSWy3Wtl21S
ISZvKW65Bc0FcMvd0jqHF/z7+g7OA8ngmZgWHaXnQ9GtfCBjw9/n6sKgZU4+etoNVyo0hSZbVkCO
dgkMd5pTgTw92Nxe9A86Q0SaYJaNIyQ6OiaEdLR7LUxFHtU5hDZiREkU42Z962bbXpER/L5m2Ncq
+aLIynZFR3ma2UrN9JSuIsHK4WIa36Ui7ueSHXOMNgM7k+rS
`protect end_protected

