

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jPOKnt2dHOagW4dFov86UptHPGMdrE6d2ZgqMnfJehhzqeTiVLl89did3kf45SSrRMnQy9YGjxY6
jqpfslmzag==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TbXlwhQ0d0UG8+CBDSNOnRgRBfh1oNNVi5QwoMGV3zJAlkTsnTywwNiy3IArHTxG6Niq+d59upyT
QOuldsHqtyc6KQBpxueCYJG7Fv1OIOGGq8mGjrkLmbJVhJEwBvPv4mlhsXKQ+/UhmQDpF2ZyKhkK
EbgpRIm7ap2EmEdPduA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iaTK7nKuH82rPJSrGYALVeHLyxEbb+9Rh0wJiyQuCqzY3/f+ne/dT7ytF39Hm0BXD9csWKwQp3QC
vOqzo1FyLi+w9Ik3lkb4njvMdZauHueYbVoku659dslyFGV84Aivwjcg0Y5de7FqsEonjWrVPTE4
0oo4m4QHuK8VN0pa+LmuzTIHDEzIPM6IMp8H0IstAk4VaGHg6wlCrG0u2kbbhcyaOKk2xzxiDfSu
gcUy11TT1zHFME/fHUU4VO3aHMSGacP3N+kgMah6x7bBUjBd2rfEXkVcl+/1g+qp0xW2BzItYrMY
Q1wtoE+N2GipiyxU+AmrXQ4zQNqO11zaj/N6Ig==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QkbQ08NIPb90+bNjwXDlVNk6WbvhfydYhJZqryulAczmjZMBvdwitIPmanwzKj9BPStsPNHXyOKf
9PFA9l/uvQOwVNRTz3G2U0+6+YFy3j+qj97mRopffETTpncxm/BoroKpRNN1DrgSjygcTkfrt06N
1lOXW+551KWRUPA+fGE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LXGnS/C7HF/SjGcWlSWMUKmilNZr5UhJNWaaWr/ybus0u0ctzmNkXcydCyfmEQe8OngFPF/IKSaG
XMrlZODcxs6BdW6TBJGvkBlKfbvIYg7iCmAit8JvgZpuYsROJrZ/IapJ9XCUZT5PW0Y/S/PoGs0O
fXalNP4hoIYlP5OYjMaSowkFFmCMq49fHUdBBmi6thqlMFhrdpbAhfGoJVYkjStWry+O4YcFvpKw
Q8WXsOAh5J64eppUG0x86EZ8HpsK6EGAeT39tAy+jNSSIcnklat3mhXxMF+BE67OS/DRt5H346yK
YrLlKC5qbVgH7HjzWMBFYeVVtUec0iic45xLPw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11232)
`protect data_block
ulXutbllu7LLWCfiVDkKcgV8xVh68yAu50PJ6faUPmfA1sOLrMCi5I3QgX00q0u9wch6lOpgO4E+
VvsMNbMgaC18lZzPMieU0btyfO+aRdl8K03gAnY8oGH/ltJnxl+4D/EiSg3YqQBOIRt2Rwt+gXLN
e3lYHwNB9cKZipaBvG0+Hnlf8bV3LxVUtln4pMppMboX7rfGk2EsMW1UXxkrKO3AVyYRGRejekOJ
gyYXuJdfysOWkBmRrwSLc4n70IkGBtVPE8XRcCPJRgkHRrlHwwaYhe7Oor2Z5WZE6OdRfryJy9I7
8zH5YBfr+Yo1HRWbRp1K+zk5f89eZElQ3yauHEJw2VjkI4msh/NtdZTClFXzQRwvE+2DgcSun/Z4
oBdl3FmVumxlD2oYugQWz2IxSFBvfLy8vyNkOUPWCtcJoaPivCb2PcJHaRiPbH6a7qzVnbKYsPMD
NXMR1nM5IFMCT832JCY1tJOXPr7SgiYcz1uqEI1xMlFg6qjaPOnlgTQf0NnDFxi9okpk6B24N9O9
P7eY+WLLpodbjQB8r4YI2Bc/H/5Ro0fWrsetZcxKJ4oNnJ1IxU4Ha4TmznFDv35ix54CdaWaHovc
OS2SOywKAJKXZxB9pNSsEZ2gWyVXXy3mj2jhjfzjZuanLiWHvenTSSvyRoNKT4o21d+W1gl39SZ+
57dmGhYuADpg8drze1rET01rKFEMbVr9HacjBcstR+XbK6i1du4lJqZX0+hMKtCOBwdXWj8uDM4/
X4zoMrD6LW/iLE+7RBZBwAMz/cFYyK63Iwgq06D7DmKCFCiOQxJb33ZRgxbJc3nxDx5Gn9VWYt1t
ystEoSPGnPYwE3jS9geoYEdIzOdR+DtYSKEy7pE44/ICwXtVtGtL+/3VEimjB7d7JGo94aVoCc36
RULPOm5GOCrxnez1VW6SyZwdul+TB3kcxQqsU1tAkTTRiF3/EfKtROk9XsoYRwb5/zn0n/3MzRLe
m++DKhYFL2udNF5FxF9nSyhW/QKjsOdvDwysbabTGo6/KMilrZ9vbuKwCd3Zx+gyy0G2/pNb/LIw
ETbyYZBUFLluJIeebp5rChiz4DHUbVQxbMD6WAIKEyTkqJoOI3YH4+NkO5HSFgm8y/ApAnU/1pDo
a5QSX6GiwjfKl+tLsuDjMJN+qtf4vz6kENDE6SfthsD2MqlS7RldbuypZH5ItlUbxE55iYqdjd9G
eEqlSs+LkEgwn00AguO2RbqPhsri+DyZy8ijcjKOa02Blu2LIszydXrza+4AhT0Qi79U97uU63oP
glyTZEagBmr7P/yoPboBPS2EZRFOKw2g2E481kzgYdLZd+8o+X1vYOx0hhfKnw8RotXxTFp62iJC
feXY5pCISfWlIeNaiWmMhoW11GldrJDligh35Zdq+NBIkAQKt1/NBPagyX2jn7I+tEFmAzPqknRi
9MUruVvT8hXqaViJSl+Wgk3805O1CzxQAraq056IDVpYFTsthyCtGN8xTFO0jiwqAFGKwUZUp90h
jrc7xj+bxS3O1Mp13KvRl8vk1J28Cs3IOht6hMBm2xQhbSkj7EwSCVI4hUrf7WgbAZMCY64o12FW
iV7ZawpT488JiyVgLsazumU+mXbG7T9oaOFRObyN3JUXeE3CntLrba240e+YKlL1wmJOXgfrWZzm
KMOzEGQVg57DivQDDpfch3C1xHCmMAX9jNMfsdkMnko/ix11p6j1Aymqjwfkk90tkkj03q0rXNmH
AQDQidSWkeQvP2XCeM6jt+bHKMsSTaofx0GGQzM5qNWLsrriQMkWlnKN/1baepVGfPhAC3JddJg+
h0zKsvn1oxPxCMnwJjpEim7rUED/IfUie5kRjblcGkVdJo3hHhtBl831+eCCd0CnAlJVUSJ7XxbF
gnxRT96fEkiolERJ5yzX9887ERnRN2ZvwpXEW6wtQgU1moI+pF/LOZvBXgvu88SbKcWO6+tMpGwo
06Uq/JcXU2iqjbwWMOIkcqNoDm8dVQotpV788zrmvpTdAS3V+fjfe+iM6+dNhJtMlekwAWoY/y5P
ij+dKtnXKqVFwAwKn2UQICS/XPxyHKbVjO30Erck+ZpXyoo38mTa3J1LCOuxiYw62YTMAOPlG40h
QHlM2s4Ah+7CICV+PHvABGcvhel8WSztYFM4QIVAWAJo9D626P6o6MXyIqVs4x69643jsLvAF+ga
Zz2DLhKnIIH3G3Mov/1ArdNFxAHBQfd/d4/wbV2fGwmCANbO30DQBhJYOAYApDd2cVb8QNnAHUI2
iamAIdjdFck/xpIw8QR6sSxJJLQkrl3hS4+x4a2n9WBj+Dfg+99EVsPkQHV3tbmPGlIAjbdXjdeF
eQC0O60n2bWUYCDgAuSQhULK5h44AX0CGQyX3qrYSA8ad7IDN+LI/rQL9G/bWC+cuyaRD5pu/KQD
IG2ba121C46NpXtE3OYSixoKzva0y88lLAfw99Epy1pzWM0GEoLBapO2MHr/cACEW/pxuDeCaudY
vsXmMST44YLhl7Lh7LZ1LzvKTn/YuWVdigaHAamL/5kgdZyQ7XeJBcFlKFlFBO7YmeDSqKFbCvZk
QKvc4cg7p6QwfXvdxoISXhcqkqQ4kR3yzyTItBPwGp5zC9+x0pnp565A/qfGGrb9iTSLV303i5FI
I6axppv3ICdQGpOUmQIRQ4yQ49Vq/J9FpIwAL27B6HLhaMy7qu9BFPUSo9t1z/6uz0LYmzNb5nmY
tEYY+fuGWeXldxsNTqVNgWJuLvy8P0Y59nMfYyymwFcDtAO6JOMJBeIEw/iAcb8qyP4RYhcJP2d3
hct8jWSI4UbGMKnOVBZQdwk+KgAEMEiDHT9sK1RrqvwFtK7Fv21HxWMGb9EUL5f+SI3NqQhrj/LI
lEVFyMtoRFCnGwSq8shGjGpL67JRUw+b0JH+68IyxJ9IplvnKqcBMdP+8v9erRIvs4WClkXRbzIF
66YVAue667PfX/88gkAw1pYjdFM7zA+CxbvW/XgJIa6WV754rahpje8ocP2MsQlX5coJW3favf5S
L+2Q4ERDlN5q77RNrSkJsa7h/9rVgWznmnC7c/SPU8OUYRtsgPcKi3vPZOwWwAJTHe1wD1N4k0Gn
WASQ/CoBv4sCToqnMZU9qraWpHAprqMcYJt4iPGozYaLL01Mhhy/82eugCdfQvJjq16G2/R/1KQ4
jGRQ2q1lf93DL3fFm3qBHAoc8gzs5QXucumFmcBgSAa3WoGrfoNEe9wAKTRSQVlfGqZz+GBU+Wi4
tftkFoegzkNwb79vhbcSaVzLS31840WUVW1jSqnyUL2LyCzjEKgW+tJiY3ulqZBHqESnm+V/FPFN
QL0OljFgxchjZqxYyebgtlWhev5skN60K9A04NG1IINEX+dTTsWr74CHDHW52wadyU9G67EihNA8
k0I23vDRGmpQW20x1+EBMcp0yGfHZLzQGR+v13/N0N1yYBR1SiystA7hy6J4RoguRSf2r0nTZ7VO
w2o8LA5rzGLx1OP8kzswIhS9Dsx2xNJ3szFbqPWZsfI8eoQoHGA+nAZoj0PBiPH8TwK6uqfQAKV5
vQp4xghUReT515e7dq8J3YVKLlwl8hYPabl1lXgH6uuOtvgUkqnkvTxP/saiyII/mHMA17/rCv3t
PTPvC080iE/au766x3gkNeEc5uOizHKN6xfh0LT4NMP2H2Ql1wEAEqCYfIOXCl9QBpwGrrZ6wFPG
TgvELVLkNWkSwcpOgSrzfB+Hfv/uBc++btS4utjqb/3LXRjxlQuSfnUv8XvvisxK95j3tZRnnjTY
PEhdweOmqTAv4e+coOmfxkoC5VU/q7Arr9FuaAQ1d6EY/GEWDeEDolYBpL7YPfMiIlMXBqTeFR4O
MkpjsaDcyCF1yJExTrKPDh3bs4t0hAEH7V2pKoqnoGWU8yUCe5ttA7Bil3mLJotJOe8FcoG+m8VE
nUThz5LEiqIaMMl8JDGqQIjtM4ICSn8jb+WOM0u2DaOO/Ck/iz+z3SjE+tOCddrX8MlWeTSOa3Ff
EggNT3CLtnKPDMtXoToU08RDG9r1FZf3f08r+eiShORans5dK7Ok4yqP6SN1MEFPdm7AF5tff4h/
DNyFXCrH8HPv/G/YxZpnZEc+DkXnOx2K15Qha3vvMtG3M8uLxPTL1PEXHM1sOXXPZDf3iIXrAaYH
zltt82gwIJ3Sh0Q0xfKiFrR36H93PykIpnnRYego/0OuanNOQWpn6Lwhl7w6Lzfqiiyy1H2SCcqy
AM83IbeGs2K8gymYJGcMuo8rjgWcWcQ69btepwntrO5+67NWQCyNuDdH3oPwrwR8nKBKdBP4oMB9
JDJgYKmke5boIvfc2fnzVZexidZD4sQKPvYU1fAZI9vIW0IZm6LTP8wpJFGBQkeZbwhsQ2rMv9NB
CDfTaGkRiQW3RcKTyBB2Sm09PzYOWSi9bHx2SNICbMYgke5DHINg00kcCh+LaZM27NBktyr523Yh
syP/t4/PVRygtM7XJuBmea1JPL7BYy41v4VtCqehFlQfJj3z7YhwWT/w51+zPzZR6ByUoT5wPsfJ
VdezKwBqq0Sxev5uz0ahE4FZdXYRY6PBhryjP63E8ErFmG3AmaQi4hSrQfhqouuEeK69CxUm+t0Y
FaQcXVLTJ0cCCAHvghYCuWjI8w9MWJGpacl+bOyc/r6Ddjw9PIa9lWcFWkM/O1COmw97IRLINzpO
MldM1mbRrQ8D+WYF6BUyENlZsQZh0FJV9pq72T1VF6INBeZr1dmynbRaIrE9F2ZuV8SVZ0kKwUK0
gatKrNRmmTcC4dws/gEvM/P4DUpQHRA8viuWN7IzeFmMBV+xIseuLJSBS+dU8W/FPQDxTcGAzIQ6
t62ZCjjxAkAynzSX8yDGFQnU0zpt/1Zh61kyZvEJUoPhNXnqTC/XLPXgSWrLJilLCVY6fdAcWpK0
ecNPCjc9Bwh9Z7fT1ALot+uPXXpWaOrMlrNpTxC8GZNl8v+bNYfC4EnPcUXxWW6vYbEOOQ2Ufg0Q
Mx3aSA6jHKAGU5PIwEnVPNbtMpe4nW06DyfMjmssVaUpQ7oAoykEldOFvlOYLsgV7OCmhUXgBBnQ
hoAjoHdwqBELzOXvXebPK9o0R2ZZmh+/DMF/esFlDew0+ig696dQsYuhLxVO/x4ZsdsrAfZbZ8kb
TOwHQaF3kay7CA1BTF2c1YFH/K8J33HzNUFf47XrbXCOY/a2Dsn43Upy7OKUr2yvUnFIAKLhTpLF
jG389ElGzS9U6uS+sD82BleqxnsuBqD9f9IpNYr+MtVGZKQwlhTTwNJnOgQS4bNEkL+QZrSLGTuI
qjLbpWsmq+OIDSEP+4QkEGoKtC2psiscsUwlJK0sp1cRZ4Etn/gMe286+SaukmTKLZ6CNImqVomB
57tdyMsdjeMrobW2dF/+N6qD/T/itxoFpTC91TeusNLDa1ZvY9Z+wUXfigOvbks+dfNp0/Do/3R9
0QgbgiIrYAA2T7KcXx/NeqA68onRDjo6CTXBjGuT51Dy20PY6275zloMwRf2YN+jnIqCcA9nZOA/
vwESEHyS9HzGXRLQ32iIzxy23l7R0x4i8TZEy4o3O+HGYpDMk/1FYhv0t15x15pIL/YG7ioc9NdA
j5ijDO4+kvc3trXk0eTvcXw6k7ouF/5okYEMmEntI2SOgvwczUTnykdftFwNJyDC5PsV4wBkinbp
U73aSbXYcc0xUBa3jpfXlAOIkcDQ1tLMi56eEcaf/8WtUcwrjmbkfh3zDyPo8u+fgiqo4ifTDHKB
jYXXVtvc9zJiwNGv2W1dxWoNbQdFNsbA+K4cifbFul58VzF+iZxA8y22gkoC1IL7xRPqiy5nxHS5
u4pxQpHAlIcLGvLitf+V5wJPgnA1aIJ6BeBbh7Fu64Z5WZfM0OQ5DooDOW2xPAxuJlGBPnoYVlWe
CJK9KsDikoiiH951P4QqOq/zTfqGwIhB1vCCKDicm8DjOvDjvSrvQVrAOtJp6sUHg9k7welpaYJr
1B6OVQmkYZrQ/4JGcby2MQrAfMQCjg3dccq9/CHMq1ayKv446IqbivIt5L/WEfXEONddclubAL6r
BKY5WfUXUGu6DjD6o0t6Wtnd69KY1NC1hg1Ra+dM1T360nmCLMz0HXa5v+WvBtIjhiixWjUTy6cd
POy7vmw/P/kTk5xaV6jMci3SAvL4urT+E1xFI2AfBpzhNdCCY7DByssYMlmPRrlIZpCw5ZD+4ALZ
Mw3LSA5dfSp1nAoz+kDgLXG3e2/c8fUh/53Bmug7C3k1cUsj5Ln7HJ9K4BN61x9YCIzFGeEghELA
xafcDrIy/mmkGkqEEMgFTla5J80eaMkoqqkuF6w3t06prZ1VCOzsuT3HYYZ5IuzBqie8p4mELyZ4
0BWfKhLwLtlFzhN828wO56ahPUPUCzxS+4DPVXvridg5BE1hxvZwQcEA+MwX/lTUsn8kYRbrqLGx
n1ODVpDUlbM4C93Hkz2UKzEHYxivnFSnmB0QT8IqlGuRFapqOymn8sadnUUE6ZjIO2PITrYDIbz5
fdl45v9P5oE25dllbv6qBXHSQAn+Nq1/Dcm0IZqAKmIUdtnCDL+TgVt6D8ZtMM3ONZAGzt8iu66v
Ns6qC9zQDkS2ebmsmntsmBeMNayPwQ9/THf9KEg3i6D1y6Byhnd+D67rv/aJP9Mr15r8jy7iJpEh
iQcCjyWygaIvGodHbFj+ZNyLvbxz/HfPfMlYwJn7kOckmNQgGPwZuSitBS3CCbewTzRHY/GYlgZs
iivIsyqcjXZji8hqC/gDtej8Pt8nlAwfl8+ivcMxgg9TeduSjOUOhqHEXFm7NVSLR4Y6NAkgJS0K
v8bjkmdG9qloB3ojrA5cXjUl7fUv0SjJM0Z7z8tI7U2yAQEaPat4IhWv6WmcLAuUkcnjcvhvGdGC
yofuMNd+KyMFw5MEqzZQFTCkbIkN+4pSn5bFVfFmlygMGQbUZ7494e2pSm+TW5dipw063tfUBu25
kyED57289+FGUqIfGBJuTw1B42QInznh0oNurb3t3QpIQV4YTIzSR80fGXCcIhihBMT3ORQsMt2H
J6vxC99fOBaXhvHBXbHt8B1ydT/Q5ucmQLHaBNJqJ9H8btAapV/4EJG0GPxNiHCc1ySqB6aZDtwY
8lkWgWAAobOZ7m7xOd4rttvYx/xbQItUkhY/Clh6rznoCyJndV9on8mhhIvhzKHdVP3xgLV04wSV
ncsKCTYzpAs23Ae6JgXiICt+v0n4K0BU4/mQLXa0WQmjh3BoEutzpfCgLGUfCVPih4oAKIzUy8EX
yXDj++Nykff7kTKzXS7gK6zY97fYZIYY6nTV1Eg9IKKsSWKd1OHLmJ0HiheLM6sNeKNXlNuU3V2v
eFNbNQZFdSiRYhd0JiCrEj0zPBdBIZn2DwWHOCqaOLD+iDA7wVuA9P1iIduETkZ+XS6BGfL0kW0N
EPRQM3e+OBpUIdxJszSyeS0DknbdG2Jqou9+HpvzA3dHsUhmrVc3oPS/xZlpWiuj7ymO2h9e0rTd
f1gUAJxEh10/MpNzHVszgNWK/X5Kbl7euLhmRmSU2dlw6WnSBA1A1HmTPsQDrG5YAaHBYxkc+qqM
wXf811n5C5hwLG3DjGdcS685S+nG/jMbwvUayuGpJTh6K6Jo5uGvDbUX7GV6CQBQ2REUaYRvpE5z
sDSnIwOB7dw+i+gyqnt8m1gYw6o6UPyxDdcQZSWVvLRI+dipSc+5hNhqKL3SrRCR6//d8U91TFgu
xV4bsIsn7msD6kO6jS3+h81a8cItz8MgzmZIQk2PpiScuJyzJpHQQlLJWpzY0+7upYPcfDvmfjes
SioVvLdRvTSRO35LktMAl2mAbGjfbLIXwzcKMUwgUJINkaVau4VzcXaRQr7D38h6ozlAwC9yACna
YravQTT7LJeK9GIoxg6x0mg5KCUmjDz7ELcsngp4CBaCZUqe9iUiwhaLgqQpalCBOriK0pxG/DWX
A8HSx1WpXdV/ndFNzypzHaPSxD532jveQNLXOWSVlbRZtBIMx6Yjii07Tzms6Ifa/hpE3FcU7pxy
Gicy9AqPNGzHonQGHcvvQjMsdQzIO84h01gtsQZYdlm/fuZ+u63dfnQ0qwRns55QNSo5/odzJBBL
4VGxAZ+mck/VIov2H2TfhP6J0GudwRiClVwZGU9CsPz/3Qt/tgAG4c5R1W/tF2XhgfuDPRA/NRxd
EFFW4sFtzigUM0JWjD1bW0i3gJ1wbWUEz2/WGtuovgWOUEbQzBq1pz1W7up4n6SVzLXkQ32GuEkn
tSWnwD3L6A/uPmAWyVqnBunD0eAPbhi26MFPMaTaUrM534SPy83eKGqGwixIJmV77r6IaBuxtoud
tE+d9plCKH4WD8QnZGytkpiWM9w0qOLU6M/jl0zGSyBIV8TLyKvkPF8HghKG7MdTpLIrytSGgoQU
6gA+desswpPiVSfYTmlbV60NaHT+n/7U1qcabZBxYm7nRI5BWc32ZYIf8fSoTgAu1gCAuS1eR98A
MG1Z3bTZ26ZaUfkDC4dF87jv4E5f0Gppr/HVrc/ITAFKV06YJPSqLM++hi/9Od9ZStQ5L4NQqMSN
9gQ0IZ4nb3+58g9oI4lKAAn5RV6UUcEGWRF0QR8LnN21LRD17pVSPgOehjb6BDc+vBQ81KqltRmR
HoMQ0q+NxibapZjQrmIi08f4cleYno3RTfW0eSwHrshmbKWmfDtb6vJH7t3GX+xyG1TN1bakMIqH
Vz6YRpwngHiH4VQeAxLR3d3DTfWGrYZQFIW3tQBWfvvAp9I79Y2Nsompp4sOmkZVjN7376Zjf3Gu
aT3KiQ0dNfWjqYrlUjGAICN5jePcnAzkCo/MtXLrpswnLX7iDVw8loMs+dvutWMWNZyfNpDfPlA+
YtOzjMYcMAHTBOARe3lGWbRC/kgL+wi74jdVyKj8WxrKViYw3r7hDp8FJbo/ZCmZOpxZ9L7/NgDU
3LyPPh+ATUUdCt4WDjiivso1F+xl1ogo7sXCFXjfOzcGN/xdZXYP/PNilbpHH8yO4lvgBa2cys5r
0ZG8zHSgbhoWAhKy9bl2RGBwh/sKOEeD+22BvfujwHfpMOq1HejG5xmSGQZRad4XfNTtQm10oV1S
myrGUBMW+NWFp6xr3A473KCciteAiv3Suc7jQGmGGLq+IrUkbqCVnRBCC0kLeKrAaE84D7R7jgLJ
b2fqR9AOi4+E564Zu1rISvuPLG4+qNcOy4z72+qk+60hirdlmMb3L5Pm+hikIbd5NeNxFRnDi+9/
3uGsXs06DL3cCOsRquMMK/mSBcc9dXVcMpdgPFOuiTav51PRAQ0qkFZ6yK9F2B1/L3g/rS15EhUI
7ndFa1NvGKwiryMa4VmhQTWQJVGKT9ZxLOu6S4QgIYReDaSc66o3YIVEXEF7qPAoWxtsIhNj/j68
5R7u3z8zt6wUJlsbjDEWFbdswCOly1Ju6/euELEle6eFoMl+RmEkJOEhF1agykGIb8CvbxWisSw+
clI9+95ChiO7LGDG4IdtaSNywrfjqVmH+Yz1B/gVieAlvK3F8+NzsWBmyOKIJPEkUzQaC09bNuAw
kKL66STM2e4NGNvLY9efyQAG7AnN3PPx67M8KLsNDG1uepSwK5bnGzGUnTp5gMsqIZHlVW7166LP
/f1vKUDzNLpU1uJKlFbGNZURArcBgyDiOvAQGAgWam38+DH+EW57g/Ag8fxObOdVi6QUjvsHNc46
QG4USrWc3zGm9peL79SC1qUGI1GRiOkUew117nvaQxXI1o+0ZgxqVR/oiBMd5FMViM7+IVG41Z0Q
nfiMf3gbK71jiV3GpDXAOmwzIyTKdRKW6CEaQRJO/AvjFGVYZ/tbhEAxLTn64r89uyII1jT/XO9Y
1iKjiB5QRH8iv+Zz0ZdFvypCmL2lZyrrtOMuXXg9cDAsjXqEF29mgVuRJ0Nc0G46naSlj1Yfccge
HaQ+CqV36KO0oxkJZkCS0qlRdH5FBF7IEBQQ7PbqoheWTHAlREOqUmQ5n0McSI10dzCfFiuWlUby
UlENKHPnafM+oKagbyIU47N3a+BmkSyz3mWyNUN+W/NaF6UWVig3YDx6uCL2rCZwu/cqMw2UHCfx
QoVezf8m28/P72FULatSx5XaUuLr1f/tkGzp/EkFxJphcU7TpYBNo5EMfxTPwuvE5tqhgcvfH9uy
/UyYYGAwf5hEp+Rfp4IxXAlH+ENWbbWcDOORCYl+sL1AuHZUMiM9lrp8+jBgMZZX2atXGA1VkX3U
IaBnrAWBgckc2Hxg+Z05PNgpq4uypYxdPlDbgIvXXjc0DKPnlndelsMa2RGh0ffA3P/URELQYeR7
FBRToKZ0SurPQcJqJJ0oLIYHXJa/4sWG+GBHacjVrO5vhWEdZrUh99g2iw8/bZH7P01mVZb/mcwt
nEHcTHtxiBmdhZaF7QDIlLK03jpHaJcy1LD7n7MevcJOo66tL0wXh8uWVDU5NowGVAvFVz8WSkt4
vk/3Ah0iS6/Rk/p5OXldxGM2TQm7Srty1N34QqzdhDEq/72RHbqvy1BgXCoWFA7GJrjQ79RNZBLE
HGRNHjJDxrGngLJW2A1E7xY6ykfEG0B8xi+ZXNa3EKk0qKdAuMcU4gXJ2uVHLRE9/EJHXtotIHh1
ONOMa92udX6V7lgWnn1I4dg91BYr/wUeWY3wAB/iE07PNDOw1IRbjbmcToiwAP7WE+qA/ZogoW+k
x5bujyvYCflDqoLPIa8KIRDjiTwVWMiXpSEFFf11821CXzP+110+AZCpVW4mZfPzNJ14hiPc9dQn
2D8q/RFu8riFY77Bthg3tiydFpGA44yXOcS5Uib+PbP6rzK8IoKCFJVySijSsJkR17dHFapVj/+y
HWF4KsfF/T/jU6XHgnMWykjTdA7l1Ets8AdHLMdFxJxZSzX18gu5Hxd9/cDRjX53A4p8rxASOgBO
RzvlPEc+oy+xgvv/QMuBwIRjy4HcrdUP9mo78hOi4Opez+TI19tcXwCGa3i7dE7SUg3T6OfhI8pi
819ahFWbJZPh+RqXvvEtVVkFzA/wDgbMRLiKUwYeHVwOY6QKVIGDDxWuvvf7x+c5XD6ozoSY2ph7
lRLZBAYoVu9J/zPgj/da8x1I12fTwU0u8sVOgRYSyLylre4qVg5Ta66FOPvf7C7mqXnMdQn96qx4
jCZnhDKCYQGGhVEbNMmzlpvIh0xtXHcvK+IAJ5z8P18p/HMmxuqGyC9aH+d29dAjB5rWZj9bmLeI
5luFhFEQpfy6Eb5G1Kop4Da7vuzqssR3P1sc18d8z0Pf7kG/HTUc9eQn1BYVMCBfryJ0Zdpa87lH
MStl6qSmZ907rC/9co8D9iga84yn+mMH2uQJS/XbqPeTKhUMSFg4FPqLMi+bUpn/PIKJO5oBPUgO
GHDLY34Gc17zk6bmQbs8+HTgJNFYl58jKbukMpRVMRB9tXuwNt/DUo3MPb5Z2+lLiChAXdKH/R7k
+7VlGo1UM8cCGFvKPJFATpYKDTl5IHV21PxH3ZeXZjuUMOyV1Z27iJVyg6etlvmiDhZMwu8aEsbl
kvcSeAPZiweQ2l4eo81Pq0xVxFpUpm7kXM97JqtZ+PYLJrUlZlJfL+yiQxu6NOm9/HLqv31JLuvi
OHl80eNEEJP0EUnypyKmqWMMZsmumz3FYw+72RwUgVn2BrG1FAlCgJTia01BwCX76fuq3NgHSYOE
uLRNGKrZeamJe/bt9m/WWtPD9ZHuD0RoW2WfZ9pYW5cU7qsnAkZqECu8TzWtxnTfEeeF0tteEFoF
Cqcg0u3t1WK3eXa9i2QdzBlGjRsLam8UUv7inTYKe3+g3pNQsPCESEqpJIh7z02wxuylRJyuvmvq
RMZHn2dYZVxxxq81Tywf4xHqjTh0EAb1f5lYH4z4H/CS1sF1HXBkueQcdoSI7jVB18EBsgTKqFsL
jXiSeYY+8oqmTl4arDrbWgagJZ9NTF+r0wZY3KiqVDW62L+IgxRUPRjoDNMugndxZfvZYE/ppZBH
rd5rutcVSpWU3wootzDJ9JD3T17vtnCBe+pT6+InLE19nobBcdhr58Pt9UsxISLeHiIojIqrU+pS
RiSxfDHnKOLzR9faB+TOp5D2iDEhQbkpOtZqEZ47xApvPrjmGxbXkNEuBBxyfsBL3hB4lnJpZJe+
ZVW87zzcLlaNjfwQUdq4YpJsyS865+pjQrBGvIWlppxdM8LPOT8xl7W1IvsltH3esv9GbZEnsMjf
+bby+28bLScgKu7SXfxlrKWFNU/EsIgljD0kRCNEsqQ3D8GJQLwNxiqXarZsEAhQ4x44WIP7TXKt
CoBOzxRbBWI9Byu4pIar6JUQPRN8laBVcIjs/bANLN4ENDc8SHmkoDDLeACJhqlBPc/4YmHKWTJc
43l3QfCVO+4q45IpEVvEA47Ta6YBRbz0BCY44KFT7VDkI/vMs+jeaB6VmH8PxM8bEYM1sqNDlwli
J2e24FCep72i4CihrkcTWl8p98SX9wR0POJ4+SYw/Lb2gjSsE+8uMSoG+HzppxcqnZTEga3pdsY+
Xiqhal3BaVpLFzt3+BPrqUDY0BLmBTper08M5eTYMIGtpLGCpXjGRU/JKgRH9cvOrVIsI1zuPiep
mlVBkAwGCR9yYly8gspFaeI6KHEb/zZ6UaLv2nvztjn4b+q8463tz+1lEHdp6X0ftxAjZ7UV0OAZ
aZkE7FHdNeS7pvbPOXQfN9k1WpKFkQIcx94brhHh/zHoj1yIKrhCLJMJRBhlydMD+/1wd1m3zaYb
SO9T7ajfx5UiPoM9NL+6qWgtwEpWWam3mmD5KhGZN4kvv0bI57ZpZFH1PswJ+MGUo1VaLhVsCC9S
w93eU6UKPo1DYFpiq3D5VzWVW0yN44NSVbE58jSD9h+NWrAnslER7pxSRTSU3xwbmEeS8FrhZp8m
ovtwUZ3lUjfEnau+AtumheJLAWq4Wlh63y+GjTCQZgoTNO7ECgioFLOjR9d1NdofNhOpC0PS8FyY
FpH5+CSToxFjpTgD4e9ChrX1aIybW2WtEmc5I7b4w4KWm387xBn2BF59MMtZcrdCiqTtvd8r0gK6
XFxKqQJhAZLQMHehk2miuLzcGhd9j2LOgoSUiC4+Z/tcKD51Kb40KnnXuxUACfU5vRllN03erWgh
K+JUXXKGcf7K81a6b3L0UoS3OUZFVOVo3VegapGdoHJDlL+eifkybqzR9jPHpbp/NBkvoQBabZW9
DHs4uEo1phVlReLymC4QcTFscDH2Rx/n5V2ZIDWDDwHJBamDydDoGZ+NoahQlSxEjXMwZgK/ySsy
W5ESuy7OhAbjftC7/BEcD8YwDeiJAPfzeDzM8LWA8o8I0hfiAm26gFczD+WYHlxvefaS8pD24+tH
eIHwm1/R1gNoCx+NMEd/82lK7C2nyOlgcSaBWupKB2fwwVLIrX04OdPuhRkSFBUAL1pR1zakHAm/
ur7m6azUYQtA3OA48pSAc0h6XI0l4Pkp0MYBeBBsodguqowKsvvgBTNsAbWA9717EaDvNUZSDyTS
Cf6a8DgFvSuGoSg1h2MG3et8m05/JI85aXUPer9jwccZsNLWM1sj5iRsMx5qip5wyht+ykBBGzsX
ArnBZ/OpEhuUXiHuCT1knh77xlQCxh2gA/ihulX9fAXCcqpHlXrHqN2usJvT9DjK79NbPQyKII2I
nd/Fi0NL7ef6sm7SzacmPeFkQ1fIPdJu/IaDcirp5z4t+jl0KiW5NayVjiWFTzHTR7SQ0tMBrEnP
UpF9P1SovOxZMeFtQgAwKnq+7EgBBMYwid9b/M7DoOPHUAcF8OHUQZ4uJigsRCf2E/Nc+Wu0XFZe
Sw2+VaJ9+SRTYgKjKU57cSGXj7WDDI8D4SsdNGBq1ecEROKYds5/mi6O+wbwj6gwIkk3qk9lHS6S
qEdhfyaSaAmZPV4howU8Skj1TngIKiMxZrwJBZSQ/fAscRBC4580BlCA8+p495QWNcxhLgrwXSlC
prZE7tFfBbjU8j4dP2Si8MUYpnsF516XGWcQtQQYMloyLgpMcuIxe+6Ozs6M+61bVFOLEdr1Fo7L
l13ZWlTq8sKZEzbGGBwJ07qxxmaKWjn90AwgK7ufz+D7sTH5cYBdQ9+0KHiroZFd2Wiq4PXpTShw
E2G/kqvdVWpt3xd5irYpmkQYyCD506B4jZMzaBsltrQcMGw8UtIpL4bsFkIL0ZVSDGjSFTa/PkiR
kHRUbsD+F7MLINbGBfAXDROvvAcXGVaofvh/UJ20zxjKW3zDOJxUHPbm0nJWmFXn9bJP42tVdJ/8
0xoubBuiMg9rqXi2imC2xM2ihLf9hTlTsd++9bKJi4GJcVL+bffgrMTFfPeneiG90fjvUK4MLgQb
IxdP1JbVkXjBZklOhJJga7SMkC6jux4Blp60Z/HQ6TEyb+lHkhDMbABxkzAy07wkDpSmqPBIpak4
IdRP86K9BfGmzT5bTkI755A8eu3bUfCIi4r9hkbMbR+I7vyUVtJpIRuiJoCIC/6pPnqwVYxSNZcA
3+FL4affuxWqnueT2uGcRJMEUVSucPUmllmEKOvofLm4AznXnn9fAWeCSji1XJiemtljy7w2+UCB
eWKgB56Wup3MdEjf4U8/rXtCS+3cbjJ9It+3XGTxiFG/jUfwn41Jf4sLCtaYMI3fzT0axKASZKvw
cwS0pL6sOLte2bwqljRC81BMAWa0fwdGOQ83bGyH2JfIka4djqqkasuWP/2Ro8Ps5kZspNJ7hkmY
tdfLmzJvxAyx7wvC75VBg5lXS/bkGbrw2lSttsOx5ccqGoUKWTbnW3Kg8QdIyOkvkEO2P6KP3m55
EdJtPxDhj6sHJ7l/LpX8YlLtRk3/uJF+UdbE/cGuU01R7j/my3PKHN6tqj5axB4WcJyVdflfSA6g
bsJ2FJzmAJnfgTvsxxDFgtTc0jpLcrs+zypC+FgjyeoVljCzMQ/X0ZlNO1b4OlmAC747iV8yiHN3
XeRZ
`protect end_protected

