

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DoylSncttFMA3kx042gUfpgfS9f7wYF6CWxJheifm9U5oZE55E7a0/gn13EV1/Vn6tAoLpUpkm/0
hmdlNetDYA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nsjL1A4AfS+U1MlmYTovZuA+LXs5hJP3SunimigW7xSFqc+G1o1qnLbV4BnmOncmqUv9X6mR1dbm
lvuLbnkHJpdv3qype+E/DkwUU+uuHlSP7/5qiYqLK0/kXVQ9CK4RGY/33UuCkCUXhFP+4VquDr0Q
ctFJ3ADjSF9u4KfkLp8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e8PwETDI60MBXnrgCDSTetYRVktLV/+TTSXZzS5MByZtHEX2iao5JK/khM4FDpq/v0uNsNW0rhjn
1dIPd1mlQZEDfzGgZ7rgxmjzboNMUH8CMdtSuB8lFy7Tjd1hDXqhliwc0PhPBGYBs/YEff98J5pB
EaQ7x9e3Dm3lUX43BX76qZ9cgUsaVwP5tX42M7Z1CZ11+5f7kvoiSco/DGzJuhCbDcHoQ2NjrZeO
tRQwYWFDIi7vBls1ETe/q8cjQLCZThAhSFjjijV74aEYat0gpNy4Hxz/UN0rUMO/XCqC2k8lo74U
XZlHepR+ABhyrwVFzKEwcRDXuuh6ogUCrZ1mMA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YvHkp5oDmh1yxPKtyY+bCFF9nl00iIDnF4JnEfzCQKeCjt2Tok2cPb5/9L9T+H/cQ1x5qpJZSOJk
cf36KzabCPbu4/9VIe9vwmzzbE9Ndy2Ov8q4+HYXDGn/u3gDUJZcIYEnVlc3E6se6bxCrEZNyRYc
iuoolgurhXiPk/HMhX4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XZ/Rjfda7p8W+LhE3BcXwsLXrN7RfTJezMmvWQf9ZKb6JJ7gmlPk8WkUFEwjbu79kr2SMWbEP0wO
UouQmHkylGRubs4N/1VfavspwJxzO5pggGGBLKHkmxqVxAWJEQ3Kp5uoaJSKWxqKIRLzeGXsW4p5
F/e0YM5v9fK6K2B07V0FxCP6WuqrungKJmSTj1Ji3gWd+VJATYp+hkh4HPUA/aDTgCzwwIaJ6QWy
QvHMQKHrEHbRztbzfLMH3RPC4Jl5v7PMeYTnCv8UcX2dwujd4zD00VIt1jMD19vjN2WZ7U8Tl83Q
sPvYlUbNQVTnqIBf7mqYAoAlbAFXbg0t5zqPAg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
W9oEpU7IlhRHusaPI9ql+GNHIwm9DVSC2OAzCnC+6IKJ88uwjAPBVb1ZKFg9pCzQ3eYRQQgZr4QZ
T3yA4Jbm9Zefp6xRm8Dwb9bSpfWex+HHiGPSRfQuN6S6KhnF8dxMOg6bu6naHaGedoe07qdHfpHf
LS/UCYEKl42CQub5OBX8k3rT2d7TIg2v63PfzfhqATfkbfG7KyXrM5FdmH9guPpByO4/YHpt0aYc
E8BPN4eFMX+DYth68CceeuLDt08EI3Fk+FTw3MeWEpINPJRBypR98Y9FSLbaKi0Yz4PijjsLGFY6
zc2azOwMT9zLuUlDXDMNsKxPLWF+DpAUc0YZ5CENdyTFUvDn0HjHbOdmLAYOo0OT5N8aUgTZN7fc
DOjlmxxMjdN8+Xecxr+KldrUCmWrf9KtJiLoA4h/XhLyc+oFnenmQ1m4i9sW9eiF3hROCA+kxzf3
RhO9eM5E+RuQpBCYnLRB/BF0/qP1uVhuxvVVlR0FaBlVrV2hEX/1LxNlLmA6QbpFKycubbsEKDh7
lZ4OqLabH4qTE09HNuySPErNxUMx6CSlCpDH1Vlo9IP3TmNKSNGkVppoUq1LmjqHAIGZvvJsvvn0
+pWu06sp1hBSSR3n1XR9pZpbGA/kTZJyW3dJbTE662scANG23oNNDbHUraNlEz3vyU20YnBsyf7k
fRLr7NJXtSqbHs8TZDPIgVwczUvua0AQZVxr+JPOGl8aP2t+IPsgfqd8Ng2zHrBMKbIgONF09Quj
FNHzh0o4dedwkRIKTm2B8T1Y45s9v8iELHHgETnynP7FMQU/o5PwOCaRBaXq0Fh9LSrSRgnkcMLS
WMfGGCt6POF4huL+HKgmGhOkYa+z8ensy0JzoBTDTyBMJoXhjEKEjExiF8dDV+7RYTS8oqx4Cf0y
Gb/KPUlgRxyGHSNh6TRWNf3PUmnj9f5E0XiEGKcqLBihWwFjDGd9Q4/KSzAzj63yCZvg1cmgy5rf
qt1cy2e3WQBnuGmmjg3b/0m0uKQdMCJiMceCLkBl4F3Lv7/Rhhne+xUef5Wn6PyAfyDw7J3zhLZo
2yvFYPl00EWKu9hClkMR/PaNdUY/BlPBxuLZTLGueUSp0JA3hK1gXGG6G6CqWH+xmMNgA2ROXfa8
naG3JxCuLx9fZs575L3KIVL0vY78ssCbnMuYLL9mia3L/DnvrLmi93NVkzbpCIvyjJSfwVwEgUZz
P6vG3B/L4YwZcHHocq7zxbYF07v0gCUPIxbDG2md+DquULsRc2Hk9vQ20Am8Tlodn4Cr6ff9R4Vn
KGFdJw1dLIgiiV2ahv0VwI3Pva5O8PfA9Se2446ju5eeROlwmuii9MhRk8NPw5tu3Gt5xFhv9UiS
JroE8jZlWboQIFfEVfNAJl/91/0yl69PePTudzxiWhVb8Y0O97iWBGmduw1xGkeDZjc70L0z8b+d
3PTh7oaPnbWqPOJknaC/V3Wpufw1TW7NqTChCAeYAYqtiZuVC+CVY3+opegZbvvKXNj8yQZNwUcz
jqHQ4R1WS9fSFrf7C+xJTHZi8oFSE0SRI0Tvzdb2u/dr1uHZiShUiLpKpDmeRSAGL0Y+JFjdU3/d
iMmd1CfyGHLckxfErRjzQ46iSXpo+vsESEciuUE8m8zNytoSjDyDHOQluy1yswugzkywVcBobjRP
CchWiM1lfj6NpeqIjkj1UEzLlCS1Rc+6u192/fo8xptMiX2s/4v/lQEsRHFw+0DGvxzlQSaSHkIp
q+G17jF+AEkZejA53S5ZmyJ05h3RFqNCCCyL+ntHlSbmzjikrkcSNTe0Ewtg2F/G9U2G+4RjD5pr
IBIRgPXT5twIT27zfpE1Rg1ZiW90LOj+j6/Rc3IdNc0oLYE4Qg1N9XAsrwgagFHNFjnE38xl/ksN
KSCGppLQf7f1Mq1cHCyBb/AInRCA2tjbfYOu/1I796X8GOUo5Mjp5SpdahXTf9DVMc1RtYixp9ZZ
JSwv7dv0yiceusknusGlbSphjCH7fP0hoLZAMeRqf6I4VvRQ71qzQ0I09Od/c+R8oS7RjlIgTGPP
ox5WhzXLcX/uc4kkF20GhSh/XloaiITSfEgyEeAZ6tv3IPDyLaG/3onChaxFtQK1WLzEhyut9Nau
pApvg3IRc1NMyh6sAiAJ1qHYaM3uBSAHrfph/rUW70EH/09Zl1eSg4g0sxUt0zWOGXjikKNgwGbS
y6drC3S1V9PoPl8nkWCN9jGws0ZvyMWSfWYDU68VEhfyj3PsLDras1qqQ1QzWZ4+b7thOVTguLOr
+zvXohqgwxiX7v7vGr8dGpaH387mBLJaLhDFLbw6wCWFJYfsgsrfzSueTBuCXqeLYiU1Ou7EnNyc
W9X0DoU+iB80vCIOgrSrDlrqBMC8+8vCFrSMFWiHyw5OMbgxCWVuh8gLuGBs3NsK6/gPwDfzlhE/
RvARttKJmg4jOzrAsrqQCu4BsKpMEB8w+HF3r+YTx/G5p/qJl8e+J4zq/f0YY/2uQYw6BiXU6O8+
7BLiyZpUuHfLoRtn5VwhaXNxrDFjFybnJpa7nKwe/zYFpO0kPYslmMF+LXOyhMWGOW+TE7ec01Ek
C5sTxuFEgol9e4QGN4lta95KWTnAx4QIpwW6h8b2IgHOvK8ByQw7/HUm8Zgvn5R8uV3R6xDKIZ7n
t8dARtYUNNGLd4Km6g7OIzq0VJo9yXkqz38YHgi/NZNioAzu/ZV+o4EFEQ+3AUeGcATzPMA8gJV2
gp9rl6/5AamKvl+DnKu1zWCQeefDL7noW1a6t0HmNz6vbaf7SibD9TU2EXAz/9sHL5jSAZjhN8Wz
C4nHWAV4wnxWs1Sc7BGlMomZvCd6tUhR8mejMLe9yCpHIbEb43bhYlDOp+kA9q1vc01FlCRzDeBz
mO1lX/DXgWVdNinyzXQvORh/4nkCG4xVUuH91Lx+t7n446tuTkR9FHTcVpi3lcXTUoWw+JCXtVG4
dFwZ9Vvt3Yh9y5wtIc0SfQ54jipYqjCLyo+z6gG8DdMmS3t/SB64HuYKl02gNqzk+o5e980KnpMD
a2EpSPolCAsDkVXV25jU1EMQBAAjdVL14HSJ0FctU/A3g2BiuF4lFVx1axDOyLIFmoPTA4sXO4Pz
Qtl0ngcKaetpjUj1qiKqPuwB8jlGNUxcM6dVDzTIqnlpN1sGXP6l7Dn5rMyAyD3vMt2UmN7qxVtP
aN4VKyoHioZcBEMGB89ANHJJ5jozaWa0NVVWHVAalU6BmR3WdSPIh5ceyyfdOTTMvfgN39Oa+ErH
lVu6etSzMM0e+pVTEi10CS6HadjSd1uNMgOGaefrhDdfW6jZw3+7Mvh0DmzwrxXPhYjTnNu0WYmB
K+1j+Y1ZHlWrGumFeKJsr+aUL+gmqyEl3RVMhaVP+128yCUrEdf8qX35hz0hLsGAR4e3aBKeaZmB
zVnfUh6RdFlyQd2elZJ4PCTeMiAceIS9iIh2ZxPtcVvTsJGf+YsVXsoqnCs6CW+KLUeZFditxetB
EEaZAJguSIB9Nbv+1pZVSKNGT97GyjtCqI2JKr+WvKi2qvM09s+Od7xjgxPfs//q3KbLS3Uj0EWu
Y9DtvEmIBlyL1m0K/CugzZ1Fj9o1YhMymfWdc7zP0psvzFnHrQyYKUOXQT44wlFzjlQamIW1x5WH
44r9RpwUrEnDux3MKORsiUxnx8eDph7F+3QvL/4H8/EEzTRbEsST+T2qHagEAXC3jefK1Ds/6wtJ
FR4z2nd+E3qpi/FU54vkuLbF/hdExorHc7jg3oc7vM20w1qF88iSaqflpHcD+Qgra2ZewMklhVsb
XCHsO0ZoFygdHC7vE+oqckB70Ba/tQUJ/EaeN220RFJ7czy95CUQwfl3n1mYb8jWG23h/+WJXJMi
Sx/2r9zUkpz/gohyNCbqlZWN0IKtUGLPy9oSODTUcCHkL52S7UCn+t4FQY3xKn27f2V2oYL0GnT9
mBdQv9rcdMpQBinbKV0Fq9uezLx00v5EiPyozSraIBj3Q19UWldXGAj5SewYQBu4ufap9QGmM9nm
p1JntWS6g0hdSehcTCFarnn/n6t6akGpepxmC6bnBfzRhvZ5wHuDk7fUDqNv6lXlPQH9TGhK39RG
gUcLz1KZdkCLDo0apfIRxyRBRejBGRYHTpUN896FHIzGHwYUQbYlExqSdbJ8rJP0ofb26tfaDSop
YdXm+1Q9ujjE6rRNv6Wx6OfCT1d2ZjXo9NpJDNW+QKD15utIcfEob7YCHtZaM/FQGfMh37lW+0E3
i3iQP6YW9aDgtriPXwXrEeekIOxwmUcFh0fswcSHH6F9hd6PH9Fv60zINW7OVSaHp65uOOa+t9Em
dhLKsFZMvTVkFQNgicZEhVjmmZdyDa4/9nToAl9gciitncQGdwhruMK3OC0nCquL9VeeeVwYnCQV
hgpA7xGhHAehSAiJTP6AjROIqpL59x2gdPebdcA5Iwqs98mXGr3slifr31ySQV1r92aRyJsEzTuf
DKEBBR/LlT//pOvIV/sh2rIBK6Jc3LbL75yH+UOz5lLB1m2R94idDtlnP7iGGK7VPhqhhdrT2jJ3
swPKHyql7Tb64pIupmNja6x+6QxbibjV4CuI1f6GSWyqO4HSDoy4rmOlLoRDAh9isrRaNUWY9xhL
KcWj3GJPR3SevcIjSN/ljytvZYFsQ6mTBoQEvFqr95uC7AWMLU9tDpptUwDul11OhczbltsCJ43n
y2NBby+5033y/FwJ4GRGK66tLT3wpnunGRXxupPneMUWo0+ZuYRKGhAyURC3qJJdjXaJK77Gzp3W
jvgjZ09t2n1mTh59udR3sv//amARVDmTon6lZC+l5r9s3PxKZCcxeFrCxcUBNBdUmMeBKpsIHqeU
hLL7PXXcKhZ/y6HVBkijP+XYyX5XVxSfpAQpfTVlvwWh8buUFzoeiq3zHeqFWYF8atXsizOyn4Cr
HE+atENG6kXnSIZRIlplWloa2nxsjX+E9iPG3Mxd0AvfM8U9MMlIAgA1aOcpEcRQoVdj0x2xE/1q
9QXU6eC5HnzqJP/A0KFK/DC+hfC9kREjJYJTznPLakVFqYbmBKBMkEv+6FFi0LH5U1Qi9xWoIGxc
L0rT5XHDdIOEL4XW0fB3PPWOSQo2tbLHlz3sfyYzMlsxmHMS2y4X3NEoywb/dYzFAf7pVRRz4Mus
NYr6SMHHBNvKFopqjAolfePfkcSWvrD9myiV5lB47Ll3xMiDwle6+GUh+s3sVRZyRB9aRLMO0wBk
eyEGc8skGclDM5J3Ybid7J4ul5NiozwA501/E6DQ9ealOMOG+p3elafZdLx7b0whhntxew4itHqK
MdxU1cBwzZtvt6YyM2KRO/zKj/1QxRUKDx4sSutmipggYMHJuQk0gqUqLJYvsx4hG3dX4xdSNz9K
IbJBVsfG3IZolJuJhmSgzCdcXszLB8iOZ1rtBdhKvOa6U4DYu+N8TasbZtH4ZjbFbB46fUEg5tlk
Q+lWCi1j7vl8hCUXQ1WQv/LF0NllY/v+1IOBgxitYl85PQhCXg5TXZZ4NtaAGeEPwcoU4XmO/pk7
oZDcUR5i1PB6HXRNDZPrRQZeKSpSbGQ0HyvCP2hIenp+2nQzI5E+KgfmvnoGwRZX5oP0V5fVme7g
DPiB9jIaszq/+20Vhoe/eSbi2gjC+4JpSgqFA1vlMvkmbp2MLiFjKPWFWk7mTpzqrunIAx5AL2CL
6ho61mxxPDleki+KVsCegMMcY3COwq4qTGNBHx5mmz8wuuLHBH+QAnF13wkt68vEKWaDZpmDlyXF
saA+8ynbHVfTS3iYia0KdgxLR+04GgNeWAwLnPgohCN2LjxDBhQ4Ew1ZY6xFROnX/fkdiRrB8itQ
gFUU4WtEBu1sQ7dHwlEgPsNffChlc5XXfKU1i1kqDBoPHNn6BwwG0a/OmJoU2IE8dDkqrGMxp04w
DoKpLRm8xFB3X52y8MyVtGuKfH/81gf+O62lXLSEIPlj6zt9Xph309vD/mssxeH4S44CN/xhc7MP
63OdeK4R43i8BQ6lWsllBgaFUTN1+prUL+n3+tUmmeMuBgIO6Yz5hASluainAWg/dakB1fc/Di0y
0818oHPgaHbHrSvXdcyeHOtZJcck++LKbI7wTcHN8phZEsIwDs+A/HAn8+zPUIy2BccIFMJjTcVN
o5nL6p8mUGUzv1bF3gj7VnBQABIblkf/QbjdVmbdTDv/NhixwJ18hYoUMWUCBf6yHyxWTCUNFZN6
D3wTKWQlXhRxyibpvPaDY8+0STiYk37+GwuGnac/UvGsqUvJcLvcvYZw8WKqFFehJWURvkjAvYlv
8t51OLARpfSw9wKAawvw1uR8zAVXJ+CbApbU+nHlOMUkHle652xy2yWeG30rHoWdwOqsKimSU971
bImAinOYkS0VEeq7w2kkRDaqKs1p54YrFS+7P7kbZPdDeOcsmQD+jKoT6N8CLG273LZp+7yIwtiU
xlQmNbPkUVqbtvaYTWN9m1elU1lsSiANwkqYgsgbKL5GMQVZe7L7hlf8dhs9swQl/MvUjc4gUu8w
OpvRMYMidCYdjc3cfe9p8iFZYMdpHWJIkHesVzIdjwrI4eW+J0zX1sqNILNpD7cqnEviEGCoSe6T
VdVmF/N/IwrKEBQ2+ZFaMEjp16zBTkY1yoFVae/+I4QxL+fufY8EPje+c9HemfvwUKh4p5F/iRLz
5+7OxyeNukqAoQd1DW8WVJ5ypT3gLdyyhFTYJjw573BNHYZfnwtEI4VRkoLQYy1E2UxtYbTvvDOK
+WLJXHqaMWo887WL80N0iSN40fR2fxLPE0vPGsAv43EQHROGq/gaDUIDusW2K9EX3n49cmQdc5tS
NFvUbL3AeFUGADIx0KG7WgsyYYoF2sHmTMUZXJUpnM1CODO1CW+bKDBn+iS/UVWuojw3PlWq/y+M
KQ150MJCEvgFyN9ZIq0vnv7g+pr3qoWAMPbRRGqodBC1khMNPjcUgtfTQ9rlh122zzq8lg4tLTZB
Lj6nqp22zN6clUgsIYbODImIteVj41JDcR/FQdVVGGAEmynKKylnQfpQbYefzCOsl5t0N92db1dc
WnX2Ul45Md6eMImWg3ge+3bRmzH+ahv8ax0gQo+jG6t99bUx/tJK+sfAxGH6MFunDvI5UY/9/Nl9
YObjkKVauPadUMUaL9C160J3iVxOmnc3/0YS6WLttGI44lAHFhRUJvULdU4ePiwZZAC69+SVCRDI
AtiwN/5tgWTfH5GqqXWblmdTJJQ/sKo0VCwkVLZiFtkMNCWd+I/aRPoz4DZ6iCH+Om5x62Ya9/Yk
N6O6jscb4KhMHeq3AAl5dLH9YwLeYLTGqcn6ZKkxvthxzaY4YpEwiKZiGIWu1tBx/OeQH0yJnOLH
pRPbEMgiIKn1M2JgMFYadml2khyg9qJ7UuQZ42sKhd72hzqgeQ8OwikGoMT/Hu3RpoIRcck1L71F
prDnln2AjREB7MxCV5irKznBthdKNaa8bsh7o43eq+VIxOl+JdmSHbso0dO/SfE7WXwtpEHNuXpS
fysrAaPHMZSGN2Ia0AfIy8BquXCFBPAVc8DBxtWbO6DvHaXyOvCn5tV1DHJ8fOe7v139eNW+Gq6w
NewVdZ0CZMUMsrKeQgzQnwyzWp9olYAKvDopkJbGpseuPkGd56dxT4FKoLEhMoyuojCW9oHGlVdN
Z64ciPqSeeAKUjrHfQpYLITZeIr/5xAFK1HkwxpfWez4+tCpi7JXXBjI6ZyvgAPYACDiCagiZzOc
95/vnb+MeBdWmMBJpT8WMW8ULfgGiIg7y+HYO/re1VLxDtlA8G6Oj0AhX6wqScxmXhYzMsL0WVXI
KsdMoa/xO3mNi8PVT4IjBpeLAsxTZ2V+yBVfgL4sS/YKB96KTzoAFcqjnkKzLNgPnUoq1P9KG7Yi
14BZOcHqjrlDsmuAa391eYkNQcd98reBECHvAaK21OKlPgPWutF3J8voHuEYtfnUcD/x9+wo7+x6
HxbtAqfZI4BV1TiqBrWYcaa0SmSrTv8gfZ68eqqT48muF/HHHkXC+eURNizvcoKjt9Nei+1HQXSc
lnbsO4ojv6lkqxliCpKkgbAni86w3144sWm1uF36eX0UuepK9ZUX6H9vXDmC9xCBAc+XTIbZTcGf
eQeAPt59ZR3/C08bkGJ3t+NCPhgZtZjnVgMNvC85so7DnoYCz81ONre93lZxFCSUxlPUsVstlYk7
vfLPtBm21jkjx64QUYCDnOhMDvzyh6jOExJG2k0A/nqWxbi7mtnKZiu5euqF02WZJKjWRxFR8wHr
QXWjNxSbKM+4joHgFkqqHfQmwU/1vPVVg5kizwX/y6BAHnYAa6ZYMK/goM4bL/5qyetLyWp2ID+a
kNt8Dte6jP57b6hTgP2k4+7KCbOSdmkzTeZmANIStIQnjajngEdHGEhyY3b2JKMtw1lwUQEcaPaw
RXHmxTBQ7qDMiWRuRW5ZTgb8CAswKuVJPiT+cp1xLx7oac2Bcw8Pdaf9HsFtDgrywocXcmuAOC0l
XUGakmGa3GpQ/e6PF6lF9lHyZENBe03oh+zSVJk6+xqUYv6+xNbDQWdiCrcd4zG6itJ1ZZdgEQcG
p4iswijRKyFpZA1lmtDpnhW+6foCMUHC8OeC1vU8iWHAhvrzDxbnEu+hSZ8EDvW0ygYPmNW2TLiH
zDvJYGZ/ewPE6v7jXR+uuhLQvcpCzOVz46xqh/EwLmLfbXHPw51JWVMfOfMCFfynATfvp+J/oWFA
KIrBmlCtoTHvJTa8msZwNgVZH+/ILH1saKd9fUebzTmSxjobxFqWYdWqmK/+6EekibxXhHdyKJiB
uuJqgGZDo6xQTRUBJ7XtEezd4jHHuXU3fDsQybJXMvoVKHjsBzkRpuEnGvnCbxQqWpL5qsKKYmaF
m8nsNEvrXRtwWqkjFC6+hVAzgVcUqJY2MjZmzn3bl2PJ5M2WPS+IQ/OwprhT94f/Anqu8NhDsHP+
A3etPOzsRWNi7gz91OVx1C3qfQwDxmBi6/J379LOfQzrfoze1GCxTr54Sw1K7Q/iMaR3I61kyvgh
0Nx1WW+r5xkc1wa0f9uZcyBbuPXwWFtxNjSxIxCyoIj2DYAr3zwq17LENSa6G9aL2vG2DR0Y3nOO
AWb8QDi2I4mEpp2BEFd5it+gw90qyrdyvJSY4ncc9ErmTCwBaCdig/YmnRqFP/bgq5gcVqTcjArL
Xpo5LdNLqnD1m7PFsm2Yki0ryE0dv04P5Kufariw0XsQJfQEyNJ7IdXkmfh6DyZDrtKNLmIaPO16
p0dNIHlGGBcoyhIVIc32Eb7niAejXMtjNHzMJ+veLxzLeTtZJTg25DUf9MvPlHr2oibTHVMmxc1U
bm352JgEdZ0FhR1Ic3RLOMalsmDxtbHl29vrQEjUHxrB2MYR/Xg/E6v22pFKtYQ5I/0PeA2LprFW
1qXegDB2YTbGBrqaJMaKATR0WAyeG5sJpTnH2WiTYBqRrUZHcMKrsmeiTwXouAjpbDA/aiPQ+7k+
oQqgTEsMlvrpBga+uyRZYSETv/Wl+5sEvIzhjoyIbbUF01xV0xvjNAjqxXzrDAkzrnGoJ9GVJNEW
ugYS1IAHi5OzPAC6n2yJ6vlKRZpTvxo4LbuDXN8dbQuoBrbhBVQNjXHsoZH1uRMNNpZsVbGGnR0B
wGHyq4rzC6cPxgVqItm6t6NNua82iJrtKFBHd9AFmlZhe7ptk0xQvzsFAPQJq0kbW34e+tI/W5lM
0ROBbNIBcfvk6XZ+soiQqHcWGBN4+YvrQA1i5DlEQ9Ti5AKriZPKRANPZRXYoidRIZETonqD6SeI
IF2zif5mEc6+0MVTajqB/CbXnrkvuH38QLUVtXpwEz3csTRdY2NXY2MjwcZtb3X+Zs70iv06o4ny
r5u8HsObTcyuApVspDKUCT3Oui6sdi9HVZmRNGXrLuFjMJ3omaqpKnsYdtDYChbrhNBDlITgXjVb
baqBI0wSf+zyANoQWm16zZTIFWYI+HLbF3+8UjsHHtZ8992B1RH+TPX7gOiu7Wzzf+zD/F+LGEoV
eDnBLC9yA/iugQOtmuAz8JULZIreV91YtDNUfcFwGFuBKM8KKvIft80C9wOu462ZlWUwq/mKoEEC
GeAm1R/otANjpFrbOcQ/RgwfeIDB167uEnIErknrVtMYjLm4omj8xuKDqBMl+nJoJGvIECVELjYE
XuXWreeFNw9u0O7sQUcjKkSJgnP7VXrT2FZWdf1Ca5P2zpYMgZ1oiz01rJv7fBSlRC1QnMdxyww9
1MwMSirP4PgjnXdk5dgU8sF+L2t7XhsusMWuUTIVvtChELBu0plA7LPQ/e+6sF4MsBe09DVzvUyJ
hntv9MR4DAlVDG+yI0oJV1pTKUEPHXD+kBpghjuogWFZmfFUPJr14qqMSkp1meGH+aqBrLmqN+HK
+MLLDMKhUj0GKhKoqVb+bSRxRDpkYEW/dRjHJxmIVrhLrnwllK9Uz3GaOjj5glZNpg5SKVUBj3m8
KizmidiH8K0Baj5ustzk7KFnmLjzJZxksQ9MAg2kh9jnGb1aXIHD9sWc9BlQ60HjpkM/qm712aR+
gJujQyXcONbGCUQFU8T2cH2Ybp/iILwpAxLKa0sSbRIw2EorO7+oPKldzcWxbZbeoXac7pN18BFw
vq7hS+eGqyQBjs04Pg726hr3fsLr7MqA2Ig6olcl+7vx3/DxZiMOJQLWYhD9fnNKP3ABHfTw5PUm
XwTft77GH6e8n1Fglfw0iXzvG9MLxYlM/gla2INNltTKcR5kFpkQKRuMVvfeI51tN6weqe/zKXV/
HXcsL3AFjw3QG0OVjV60ub/LM5vAup/6CRQfIwVO44qYdOvPJx36XUZj/ED0nnU5xrmXPk909bRB
HySSE1nFINOTHOL3e6R/LLnTXGIigw75thlDA2KoprSF51shCGpCIBOWSkc4jtPmZHGmEbtV10rQ
SzXP9s5mQN4vSaYzTN05DYbdORsyUx8ZSufkT0AuPtDm9OyQHTX/vECM7L7EqkmSdGg4ldeV9Nth
Gp3v8rHMd98ko6g+5iEbG1BEwyEXd8JaWpGBPGClSrsHEtfGOvG7S5DEeyVjpFeO6BZ0dG0TSZr5
8tKxxzReTyt1ed37GcT57rfbEI0rcCic1EEnwLoGLcRNBujwt10OzmNQW29yby6jC+l6dDyLwwcw
rS1G2dm1c1j0viWwFOZ/JmjTtp9n1+3OP8g/fvWZ+58g8VWdLPCnl7TCMyGP8P447OxMPBgwSoNY
xK4aFlitzn0w6bVWMU14f5OTdcc+c12AJNmDz1wOSY+9LWhf64q9Tg7RqzTQz1KBw4hy3ZfZuky4
P3i85LmAnBPSPAxw1ZBmVRRjXyu/mRxgXZvrIH1EOv9WkxI16C1+VJWw2Yh2GegaZU+S8YI/+9f8
ff3ZT5cWr19gwGFy52ebCyFbYFM/ONS/J1biISphJGM81yALvJSqvmA0Cp2crGyTX+hUIgOTr5/u
LAL1Fa+LQD1Z2z93g6pZ7Q4VLCcJ40VrE4mGrIMA+TUCmgMThAErP3WuHOKL/j4c4l+0ZHo0u5fO
WAoj5F85ZhvU6HrXvR92s38aA1/fv1FmD8jhMVdI18MdLLq7MzdUnl0oDOAXYcXjq/Pwih/GGvfP
rb8mg/euRLafueR4pyHZGaUlAa2k0ULqUgKDQIxRjZ4PXYwyogBVnelsvgEKr5eMiVxb8iPGJVsH
7BG3zQ6yKmoV8jnMLiiCsORovcUH5aSvKKeGvCxhBVUR0qVub1nml3dc2GZ8idTFzC4UV2Dj2vAw
G9UcdwiTRaeC7+/51+G9DOBpG8I6k+BLKeFTYOWDMuHpr1d58x1zqUTbbmVem3me2fGQg6SpgpBe
bJ0c75KjLNuP2TfUQhG+qet/ax8MRKC34feZWjuV2WwdKOcMg5mDWpn7Cwdow/9UZjRO1sdojIBX
4A48E2tuMCuT913sLxCtnJvKeQ8QjTRA7bQMNT27sWLIEpGJx0Q7e+9eyzyCE1Z0AYSxqXfYcynT
WK5vN7GkLs0/SFDZ8pkKLjY0Ua/nv62WdU2L6RuzzeZ9JSE7b8PMLaLIfVjUuHN3M99K4ImFhEzx
zXZpLc/LMW34T6f+y3DXBL+9ilnLrEibZboYa3DIDDqquM/nSjVE/ngsvywLblWyem7LFpbG/l5B
DRsmXYyLQGOGrBslPIKG7d/qPij3f+YDBa8VwE4rwcQko06zNPjlE42znwtuBPLKA4UOPaDtx1Sm
N5ikddGLVrq9K8OLSbqDLYLnJYokQ4MujqwcrfDCjSsqGXDXQFZK+jibdBgzOj4qT21zMEOM45sI
7v6oXvaE5jiy1/FKh9QV9l+PM99k/SRp1mHN4VS3GQls+CqdOYUH+cAPwCA+dcSaaHYGgd/xA7Hd
RLYLa0HRr78oqd+4Zs5/2KzgKHHDCA2ZI908ZOnHW007UUxg84MVCImxvJKkDXsjGCWgxznMNY2+
jSaA2pjjf78Rh0MPT7P/LvSMO8vW2lIgWnKC1YtMf5jKrjlIs/F+FEWSp20TOfHz2w65Z2FGvz6W
ccUEKaJV64UfksHRGSHiSTSBhcM90UtRZCv1MSHVEs0xpyDon+w6etstvgWUGkGJ3s5DQ1B4XqVQ
vdm4SRc/3QpdSphZ9rz9uPdlzYcHCII4mAcAPehzFH5Q+ry9b4U4SmRZ+1XxVEJm7yK//4KeYucI
tE3Q0ClaJ5KBrPR3/UAd1pGajfKdKqc+epooXSLF+vWMjX3eDRh1HyevLLs8NwrB7axxKBicZvoR
qnsxmzESRbZmHnbsdXv7CV8zkc6/Nfirz9TTlZZpwSU9b2LfaQLeLTwwCX+vxgaHtpqJXsOADDyq
mgZhcULr3nTU6iJovtID6fx6jn8BSitZ8e0n9Mb0Vv+r1vwzD1mw1NvgxJAzK6J3RlqgUiZmntrV
zDGrUkyly+IgduexKKuw21Gkg0KJXXBcVxqlH8bQdjTBoojfUHJUjVej22Y3/eclFQFostRkDvnq
qcEDu3vYjsp0mMTAYzcciZkxemGgFkDkfnHfotHrYAfHsEcNgNduCCdbA89APQ/8rBq5sdHXx/Cf
YHiqeS1qqWfE4lr5IHacs8NWekpPlyUnr5PvZWwU2HJIGZPmlLq/PiFfkmlrh1Ba+7GYRhkjN1+6
B7E1qTbZ2rw+TOjM7vp20KkJIeNALKjK2jXuGjGp5EIAwHPUWC1UMRW756qumWdllm9OiH2VQ6hq
5GyaqgMyf5nX2bVVExxdnXHX5is+5zlg+yEWjmfMlkT1TGZwOXjECIOM55bkC9hOkmzZc9nHx9sa
Xf/xovYPka7TljhEhMC+uFsVCJ7EHlXCjGlSF0VcqKovJUNZBleHytyPVBixyWWsHuuNN284T7F1
U5b7SNhufBQ4cFI3+w0ziOZhxkF1aor4lYr2u9PuhtOMlLREhvTbHNPKkStVaV63x7VvL5SUIf8a
NN5FdO4+UBPYWyjWZEG1v/HZlrPM6BPx8/mQfrwA+sH6L232PSVX3TSAKzq0D5ZOiXBVA4/qfuiv
jd/qcDVOjdYMZI831rfG6w1kmDSZjBbdSG1MqUrbTFDjzhjksZA6YVQSMN4h7HVcX28zWCLkd09U
cJnBitzY3o1BFfQviR/qxwHRr9PLCXGa50oTk5g02KNtn9/PHr2w6SJjmdMZfWcNXOPz6TPIBfmb
3flfmPD3PI+qX3Ch7XBr9BCPPVSw0xOeq0nu5EkFDoH/ioQEgu6utDq3V69GJ65ufmjLAlwIK4f6
aY2AuIUlBqZ1s6CW2EVd6Ifeq1cETt/0Eyq02x0b50jdIT1fihMFmAgP5X8Yp5rV/S5j+6BIsvmW
aTBxdBJ+9X+iL35NpeKzMvSneE9+S1fM58gyH67MeP2uM2kDYBMkCkbnFYXMvdrf/sMpPqkqFw0U
I4gwwRRd5LEp6JK7yqSGWSKEhn27tcirTT7UZWe6kTjn3Pv1l1pGRAY+IrtgJwKtP4t1rzpKAjjG
gZ/D2uxk4YY214cx99Wu53TeJn785zK/1jGMI7JLOnRloWMYUshobDyTL/2jT6/9rVinViX2Kjfl
M8PkYd99U+L5DhAmQaWBj9rnbqJL4GLnnc7lFrwfZdWPDeWx1r2nmlQ6hNCwllzciUgQYe53+924
N2ubuOWwY2ylLR85sovwN/nZCnSsiLQkKvqgubW0gnsbcQxhaee6XO/D8P3QAPNSO8W6zd2egV7s
LklVHJ156uXlPIDizJg779ujtrh8jiohZlA2Sb5jUGPwwYxNfSyoZQk/X6+DOy8JzUBcVmPVr+hR
tkzQmQnRg7KCuKNLfCZ2GYZur4+UG3Nor6Wdb08V8as3id57K5zLYjDUa2nd7QyA3PZ6k389VdWm
aMjts/HfV03ZLABaIPPOu9fe6/KK7s62bjfGvkU3GLxBtlb0S2zhXWP71KcMSQP2fuCowbnCLDna
GQ8Rffppa2H9+a0tZ+4CZ2sP8jqYydqlrwP/dfGEV7mws5gR+h0tSfhutof6afE7nVolcdESsx0H
W5b4pLNZHVbiutCltFC3T4MuIOL0zQey2WQCgPEvlu3T8Hf2oKQMkmBwzzC3NK7t7L9NQCyzudxf
MAX351oyC4fHNNVZ4uTUw5Dn4hnpqREjR7BHChQNDOldx5kRq+ywVNSU/ApEUvG1gcT+cIUWAmKc
Kp2+kI1Jl8gOHVoY9reVknnp1RbRh8yX+EkKI+DTb2rDqnUYvVry1dSjImOJfWAze0PPyiBitO9s
tJknUdKX+ZEsrvYAqzIQY9IvlVj4xhwIGQVNsDp37hQOrpAP+71SrNMDnUZ+uos1cD/ab0elHJMw
iPPPfmuekGqtI6KldFs3YXliemRnc00n6Zu2z3Csw/poU1mwfJGjemzFFBxpaQoOqLOxVkPCrAH6
bcq9tOqGmV15pPEUvaXHBVVcqbmiCOWptJ2QwtcB2vMuHtg4B776Bpg4A+h8s7qwGSF1BVy84on2
LfT4vKBjUr0w5jdRJgfyg+jz4fOe9BMTuETQ1uHIkmzERtYL/W4aLBcvCrTfGj8bqJJtQ6r8Xmic
IwpwL2kFTDvXCA+DBA38rl31WUd/E3D437pXenvcVLOGDWmZvDrceqH3wiGGEhDqSKllXfn9XMsd
DcOJQoXl7qklk+oGEx9c4P5IuyMSBbwGRdDUQvMhp/4mBkrbKoYg09KTaNs3ya4gBFfLDuxfo7V1
+cCtBZgaaWgypz5UNFW5+DneKZiD8FpnigAI8N65qrTwYax4wgHI+J8i9zf/QWSzOQh9c61/Yq/2
/sYtWvBZWO/G8ckaT9U6Ci/I6Z3C9Pk3J0H1j7Knm0JHEIE95JJnN6wNshMgVDtjcKuYwl3vPboV
suQMr3d33QGCBZXMp5bN/2zLqIBYtNiBH7Jvkom17yeZE3MBows1W6vdDZqWdfQrfw0P3jRXGzp9
8AiGPDqw9/UTkMlGJqDOkm8WRnDq+8k/etEOgpsYPXiNgzXOJdk3oO2rceCosAbpc86ylarBSthy
gf1RcrBdlaHSYh/6bEYQ7csR3CGs3NcW2aYYUjYFbV+97h0MftXxYQgs2JN4rpl2OMdleAuIIQDK
ZBuTY7raXBPgdT8tbGX5Jp/og9wYNXpJ/IDmk5CuAuDXFisTZiV2Y8z978Fm7AtMlGlNhqKt8H0U
hZeOt0jk9sBhCuuoEq4iLUD7uVrnSjf4Q3Wm56KGSAIlLPOLrGhqE7Kl38lb+dnyk4tA0QOkGWAl
ti67JG839qOhkmV1i0sqv2hulZ5LzCoHSazrooRtlC0xj99aAy6MIXydR0YMY9LuOvnbRbqw2GYi
66n07ZVo0AVzlhGY6TLbYx9lyrdwfryElutGwwP6JjY8bFbdLKLlwaWXCwnTtV9H1OGNnJWUfKjy
j3bRQuyGL+7C/WKjGusq3tq51IYQlhnqeAom6nxxu+iKNk0cOb/k4RCx48SaoHSl0Edb/VYI2MTP
FotG8yAeo2JwkYL/aAdIICMelIWa4DhtaxOEYiuMpx8Kq7bwlGQnmCbn1baX3yq8Kc9+OeSqXbSp
HnqfDjUU/Yfya6Te6phY0BCZf1+oz7dzlELW1E8tJmON9jkN/sBKxbIS3IbaqHe5iWHsIQrQiEx4
dwVOKLykaM3Upa9XoNDsGWsNqtClkHIk5iB41KfuQZxWw75b6hrbYTLYf6f42bGhq1zdgnhni7CT
ye5qkHSszmavkOKpyKUNckhk8XhUww25opRmXdI4StJ+5oihnsuRxjtAmgOTiTaEnNEmSzdhLUx3
Q2uUYpExmXGRAz47HGV4ULrM1YWmi9LcPPFO9ppvB0Sd7QXN6kxVbEaV1VlCcl2BbJoWpdcmR8Xn
sENB3lRGuQphqhn+TwZ8K8XoNs8sAqoN2+zHosZ46JMDg4qagwG9oGKBT8uiavd00K+qHKzL354z
jKPx8xFhfFXBAkPSL8R0nL8GQoM1CWSIbzda9wgAT/8yPY3MiangvjXdSqxd5Pkbf+JbmuDsA/Hz
BPMwcpK4mtZS04jZQz0pgS3NKhLA3JVY/1XR/BPGD3HFSfqoufFdBbmfQd/GcjmyPIwJl731yx5L
RdKROSMn9waJwTEM/bzGq1IyZyy/DO4/3Gn+F6U+Va/Bou3NbaP0il0xGAyu9RSNFougJw05JUHC
KdOLaSeb0PZB4IWfzwmNgihSKR62vmbVorqg6+vpWwAfc65JQSqoj315FHxYL2ULx8Y816GNXrau
cPapRgWQBKbtDGq1rawJFDGELZOICEt51H2fYwpaKbrVNGTlheDJ87MpaxQGqGiviLcYasmRvS8U
DxUB4VFqYcWlJIMKZL4EkVop7ZpbktrwJMhju66DuMfk9Hd/whiu3otU0WrVlr9pt0mba2qXrjIA
lFix1rZYV3j2xPJHZWRAWu0Wgfxbwmx8dlI86RZ9dMn8JZmdNjnXLdRG4bWhpDQilp92NdDWT3mY
FiGWf0qTJj/8+TECt/Y9T5+QRaMaPEzC8q2cvTujJ3WO0iLIsEwW0rSp+WUwOBit19WrBhstsmTR
wpxyrd77PYN3ABkr0fdWvrCbgiPotAXC+dxPtyhhX9LxU7J1JzsES09nO6o+cB9vKgdEHRaiAqNQ
FYanVln0bt8j5UJh76zWCQGZ2dwXvxQ8d7sTOvBSJLQHMvYRWdJfE+mlrF6XuXFYsk9rMvPEUbDp
NqMurs8ABXX7cviWZpnWD2fJCgy2rPGL3H7RJdKy9qlAL5VgtkfVamRcmBTOjAM03UH95p/gzEYm
u0PdnEAEANZC2QitjlRUPkHQgkIwW0W/1FXpDLBrjGUuszb4rhBQaAy2OZHhHnlHkpW8X48Ft+Kn
rfD/y5gJZFFxG15nclbgqX+5C0ql3lQWkk7PjaxaPf3D9skiQ9VxERvySijMLvR8Cc+saJYGbpAl
0VkmYgr5GdL2FQzSOV01esBsp7xU7af7ql5xiLVdorsKFNudsMSbMybFi5iySx4S856qR9UrT8AD
h0cDOdYWkT2rh365KbN4eQ2AGDZLsxJ9EyN1sRMgTIV5KBxo/PN6yUjJCCTlItURXmennlmdvzE+
0PKPlnMqgBLJ/TU1geqxbTRYCoOVHhk0n9DFJL9ot5isCZQVC53Rf0c76fKpM7+DnOBIZ1uvBnIZ
CSpw4XbHboQ8/bSPNgDsox70DDNeatnoQ/JggGCtP8e5O0fd87DfBLw9lyfR0zscNNM33M+EYHRK
Gfo+y6eYM5a9tFmlHZyglghnkZMeG1c5DRchfvMaSyFA5egWEd35EuTcPSi1L8T1nv7lV7aLG0Fb
hJt2PELEb+kQkIx/s6J5pQUIBCJlo+tRouwTGBK7XGYAzckp0yR2UPbwzo7VTRNFanhKqFmTWUvf
1sMIqp+wWLLT13YJjfFqMg7Hmw9pXB7KENlFfb8TFFDtBTu6tOScAmyt2ocnqCOsEVpqo2U1U3Np
gf/APycmPVAR0qDwnHQdsUmKYpthm4midPyXU0yX8/QU8WrlUf+/9AVBOkSfyW4Q76FhR6s9BVjC
Twhf90apgS3PAsvLQk0Ly8fiZ1sJCRP6DoTaxiMRNdP+6i3thx307DSZFlN7U4018GBNxCjFGZaB
e3cMC9ggeliNhJ8Fwl9QkNz2KcVV1Tr5AnvxNL3LVgUoeAZuRiTyGZnuEtgVPNWZZ5UDtnNdkadk
wSxivJCNoewryxLeqoOIUxPgZjzi+QnEOOPAdbm2240xd5ZjMHXxmgXMSqUqimSR9TACi6SEql40
K3KBNhvoFgyL883R7Teh9cihChT5TciPx+iXe/K26x/fYcqF426RuwyYdvWx3Z5ofqJIPnqyKGTz
IdZvYp7d8lEhycvU0+u+PWr9HLHc7RxjUZkMrZ1TLcwsCv6lnrLpUvRwz7/yTrqRWn0MpBMQSHyP
4sm/Fa9Bb4jjOM2hiDhLVuZrO301D4zlhjLsXdS6E/61mNYPQ1bnUhPWSAEcHv5igcbjlDTP+UGT
K0ZbOqK06Q06J2rfUDN+imwlnGBi5olm94GDuw43AdUwLzskt+dO7RA/xoOcJJSG7DFoqH/lkPJd
q1ZW3EOjziuKe4qVmWeznkJbbH0/cV1Gm5iw7I5GwIzPph/YLn1nXKIKUFhTTKeHU/rIzxqlMcbO
4Xz+/qXKJO/URuYuxoOauriUid4lIaj5sOf9ZHvUILe03Vnzz2NJKy/dk78yMPMKYXqP9lr2FXYP
dZWlhE77D13RWxfnMFlH7lSVLVFR22Yig7qlPrFeazv0fEfdN6UOnmqGg9tcbLTJzgyGh2ttRTjx
ybturZwnHbTLU6Cxgcu3LdOAy3BaJm56Nss+ukB0ThlxOkRW/64ckeboobS3fkxEnjNVGlVlwQl+
n2iruqI8ZUsABKMqdtIZWAynMXbUqSBV+myI9IlAPQvMN5gzu27QLg+75KgiJdY8Gs0QVe90Qax6
ZQHFWYofXHhTTsZTtFT9navYtb0bRxZwxCvuAXPYIilCx4qXDIi9OP6ELyc8w013FtmBDQwJAGn5
8ip5L5uKxhmuA2x26pQhVN2Yw7jLQf9AbIaievhjRCJodisKYBr0kaJdHVbcnZ24CaGiZSkULCtj
Ee59aMeaUdcbeYUz+XvT5obAGCtew2BYGwKpr7f8Sd0M/6Kvd97iCCjhvdS/3N78lz896e2mAroq
acdlF3ce1E9wvjXWJ9t4af9rg4jAoEBkAKmMzvIy23bnaQO9yAoEaAXVQPUar/jeVzVw8L+ezEDB
69eVzLPmMu3FQT0sEOesj6c5HYEw0RF4tA6Yj1OOXbhpLogmqYtOh78+xa+DoY4aQdhCldw1RwPD
m26TyusrO2FtZdT6NQof7utiCQVWON7Rkjn7cLDatWrYm4iIVRiXduK5u68j3T+ikx8PVtJOICA6
XazXICno4vFkdmKXh9E8LR2eRJryllyow3R/F1TlTRzmqyhIIkT0w73bGPTV52eaLsvCv+BJLIHd
mYLc2Uvk9kV0hRaOrWEf9cTqyqVqyNOdNjRtcaWboBM1qdYUyT0I+AOt3dAEeJWmI2+H9NUNlIy8
NxT+GJiJYz8Xf61UC83kjIj1FU8hjT8uaDvclYRCaLOND9aN78lfh7e+v4d3s7Ll2uAzBIKqAAl1
XvpYPDVnLP+JgGhKmDv3tuIqKN0CGmRWv6OduyYekelTAho0JOWMGzY1GHiuvfnaBxVVT0wVEuJk
R/dY+EpUGwLcUE+D8VN4rtwHm96IAA5xCoOjol4UuS3i3v0WH7Mj6oOxzDkL4QnSJHA4PwZuvEy9
Rnhrp9sU5W7bo0fS1Rolfs3FRztz2tEJN3huumJE9mpg+eEvtE3ob27A4mPzTgCfiDv7uLkLI/5T
GxnyagIBaq+h5FNmKaqAinLMRGzbdmTUUXJFDSdGNOGoJiLt1p2ckCl9F7SViYsFs170+wFYY0r9
eoh7qvY8WLuuGzrnAaITuuiJziq1NQIdYrqDEBdO25HSrLgyh1Quorvfe8RoPHSMUY577Sanr7sP
/BRidrhjuJ4ge692AO+c1ytAaCpBbbg8mYf8wMFcYpnb3RfS2eThv5s/HHaCFaSSwFUN2h1KSdDa
QizUk+zgOTldJZgn6cy15+ZwKi0C0Pcw/qNmQlZtIVhdyBJkJBEB4ABpODDjye2f5xhH++Hl9BVG
byxthAOYlEu5xfLaj6lFw2YilToe68NG+Mj37bBA9sGb74uofLm7rjZXDUYWAAHDRwt9ctK1+w4H
bGQ/WfAzr/C0g2N/KS6Y/xPmDh5axZ6KRPuQCIE8z7HTiKuf2CVyBAn2mXEiRXlm3mWhST8ephwq
OI/CB75FL2mNNSyMJFnCnbOWnkj1FcPpK/aTFtZ7mRfxmNW0l+BBOoeXy2C79nOp/30Kk+hhilfX
4Dd+gneV5DcaZeFkiO9OdhroVirySKEUGSEMHPv70nWpcJDRkg6SrLs84Q8TNqI+LM1V0rppVGVl
3ey0HEaqmGpmw3VUYAlDLwE1mHczTdCzFHNXx3djGIzNVpkJ7OsPZFxm/y3QRQYQEBYuAyRIJPBZ
a1lRVY+Q+4EkCMSeWjd/42mG21d6BK/vBArhySo+4YiSJKmNQQITfgqMlyqHS7StiPyJMBt/t7Ys
HjlfQPe/bx4hQB32/TARKzmV6F1CTgyJ4q94QKsWZCYhYagcUCri8A/Hy40qgt+IloIO3iU834/s
4bTro2tSTl2DtCqe8+9AE8UKCFwHuO1pzpx08C7T6I+nVKLnaY+iJhSUwI+rrlWfgLa5EdlLNPcM
ofbI+u+etwfpdsY24jfc23LG0+W9TLTVTxo/0J/si6ISYyy0FPF/QX1kpGxZfhuQXcZc0UYK+MlZ
Xt7r+kqbv/hH3RMw2juqi3LA8/qH0D2eCqMMmR8848TAFAUck0poln9n4r0MJx5WeIW3GDbE23OS
1HesoPPlpinpWbVvOr1T+IZkfDJfk/YwH4EWrVl8YWR+WzFuFIhaVSx7mnDWj2I81Ne6LwObOE0c
A2k+Nq+tDtP4/UYiipyz/nIZPs3LksekLiutYAdDVEgXMQcyZKO6KcdzYRbM5ruSNjG9cMuyaKet
5caUT5/M2y+Ew6t+7ubV1WpbSnXzTyIWRJqVmokY6YbHmVYmVHTOJ8HPwkvwcmO9fhjUvFuW6nZl
GmSocB27PecRHxfYVE04eG2vtaoLQ7VN+3uPItAnhzv8AQA2MtUeQb+jtZ5efBpkGAwDbqUFsCPs
HjMezigDnJ7G7XQr1pJXL2jkV/HVBtLDP5jpOyoLFoBMUPZGFeLWGGHWbWmr4ResESeLxf5Qi/Yi
NJHBvLh7M8NPH0/sE9yWqQ5p3DENmjGT5BYISr3sm8w9fAmp1TOYR+PNBWT9mVTThk3gljTUZKLx
iUk/xMKdGXte0F1wwKyiLhfOa75kss+QR6x4OPtOJOd3xVyHG19l2YHQlidx6dsm0jBCeHA0jHJP
IEO9+uzbPUV4z9AK/U2pM+j3lpNyaQtTXNRxM+7JL7eGkGg9Wz91HwkMRdiSiycqzuQJ1pk5Z5UM
TrvpgSD/Pqh4jBinrILPyKErZoTJlu+rLXW1l4g4Py9zFwdxARy+gvvae7lQhasmV2kN7Im94KQz
VmHdcQskf/DreAv5Zr8lIDC13vT6KE6rWZkl7gN2I6yKrWl6cua7Z2Fy7UW/0Ni+yN8kaVkDuhYY
vkEXvIIVqJXX1IkYdj8u3WY4sYadZU3r6bv/RHEodFjsfG2gMLB6TtyOq3vvTdqajEYxuyB+L+7C
Xd5OW0uKQW1eJIMZuc1z3wALzgoKE1jLWulHex21DWXppfXFARHkc4+gnDY6hK2HZth4j/rPJhiQ
rI3md8H737bq9OsH+9gQ5Quf1a7fQA2Z9+G39/L+ymgmgNiS1f0EF4W4l1scEtM6LXxQ1PWPuaIa
TbUNxXpCDqLm/yR1xAkJfJDLj4FzWu9aeNqpbG20NLN4ifTRZoaUA8+xIrj94yId1aUK/NuLgx39
luvmM3x5kBApdV9aryGs3BzyWiP/O0SBcbS8v9ZH9DxDXSmkdHsTqBsoZchUIHm4xppTFnJzg9GY
q46HBpCVEpOtBL/qdxYCTc67KYzk5Ty3AXWUFgQ1IGoSgmydvv4SV1DiSdI/kk89+iBNjTCB8MP+
gtLj9SsDAgYwdPrpKM5lpr0Ef0lt0kqKvQ8gDW0oCsaO2xbrLpnnzeKLy0M5p+BrKqu81ZFNTxfU
ZZ9KCb9cDd51TCUdvrTarJ7WBr5a/ilDBRVQtrxJO57MWnRvtuKpylRO791TabBdQck8kU/k9vVv
avtwOXonzTMrPP/wyUZI3XDZvbUBNb6RJLRneNOE8CbOpQ9lIYK513zLdPh1qVbdzOgmojtIKJT3
cu65aqjqznCsPLHOH1KCaspzslv2eHqsJLAXrcGpZq9tSEXqyMK94jOzNVfU0Ym4AjjiuEjK8FUK
u7wSKQE3D0un9cOJz4jHgOOg7uHyLI0pUJZUdv/8ZfWwxYuIImPgOJTiCkq8vJepLU+4LqAGMVXS
RAatxEVviQp1UjircFHH5Xl11hlYkEPAt/IjLVYn8fNzRg+rvxnqeta13xAWPkfS8nU7W/GD3X74
mrW1JSDYycgF4TZTq1DpIlockfqfiNHnR2gzGizgW2BphSBpiFVVOr7A2UImdWHk1gyQxN05YHy/
S8OSRHIV0kUVTGoqO3FEgWN/BkyKlcATmSUnud3WuKQ5sHkaItuPnP+54iiQBVGUpOCLjdcMYzcn
+PWhUQ8nEpV2DdODBb/9D+6FBYfnsnINtc12HbhGD5ZNhepzv2SInRWK/LrV9wNt6gKSvIPCXQfF
D/J8MoQnOwddtNmgEAXovb4/zf3ddNjmiG7AI//HCdIjSuhkEf/HJK7XNcDZvgTeazngAH9eryoG
m0eUSUdnKGzQULo1euCCYCH0v0wGc4kOOj+zXVQklJLaZp4/GOV6Zd8gsMW5qAmWtbSvdvB8JnlK
dlAaK/6AMrsPZviCHmvyyAmURer7NmGjl7ZoYWUs6Z2uW6Rteb0IxfLWjzeACHRH15RdZcUPHbkr
2FMOqt14zw3TsK7fK1peDb6Eo2ncf3xt470vjgIaeqhGnp0dcM6309LEMOpgNZ9JfpXhXcdS/EjM
UZEA3Vi7bBHtacDAXTRXNkgeBi1AJHQpyl5t1FAa+nsSfTcBGHBIhPk5Pfh4xvvfW6jEf4c21G8R
x6DkBpRoNAGEAehcXCNo4ff2UI1/cfmqzC3474BrioFme8n47l7oJBEcJvalufX4uMja5nigkHC0
AU3LAdvk6Yx4d3500GDgN4IGPKzG5lbdr79Ni8OurXL+hYgp+NivHC4NlywTZjnsKvj5LQEBhi2y
IDcjoI/aAw/cDbA4kAIg+Aynai0ExIIzO7YphMgyend1ysfugFy9oELVAOqjezugeY3scuj/kwIn
WxsNFjy1YAhAF93oBYceX7h7xCbGF1IN8lCh+aButNYxi2wUMQLrcjP4h3/tnBF9WNcPdqEI0xDE
EBnELrEG+dzLKTiCCByu5eOIbPU5xo+rCOQ9a36hSfQmZvEmZdQaaIbPWQIPyWCvMj/3umiF93lL
3IKU6H+NoK2/hwni1B2MeaNjXGS+Ri0QNeSwjO4YF9rnzf1Ua8bmMid0z/woIftkBQW6AcivJWU+
vocjOYIYfKqK+eltO37rzEihr1HVEWIB+wj7T8wlWdaj5Hvg5EvQZ07UikZcwdgFUdH93Vy4p56a
BBDUFBVwPefLiMbo+xKUFXgP55TUqsIgZEGjyV18ehqagQ5RITb8i9mISVBaL13OVGjoEnW2CUf1
qQrF/ZK6vIX/CmGSTbtzZasDsG6vLOOcVF4uTPVryvFdnMbCM4nHARbbXnOdtDFRJYvOOhl0FhrX
gskmvOOfptrFrRj9M6ikFKa+ZOFquQqkzle46lsYdqwomUkKMRBpWdek9Jp0yy6KR2TUOTOcDjGr
7PRmOloGIn48SEXRRH6N+c68NNqS/gekaMysA1/KFUWwOylF9MjTjYGYpE/n9ZNEIhqN0IWL5Tje
MwxJ8NtZzy477uvTiCngYVvdMKupTTKH846Z4ZKGK/5f3O8XfLjiZPkIjWqREHhgCgX/0UEGfFLI
yQ3rkLrIpY0y5ZyeIB60xCLKyCbMG/1PVlr6AeOv4dsuO81kRezw8EohY9Z3KSYjCxWciz+NksBW
zXzr0hjrpF7HfplSnLRuYQ3SqZvj2auYURLsla9KD/9KL0zJEgVdBupTZoXfOqj14UBDOs1YfxuE
G3qKtShAL9X7dyOxb6RrW0qCZIP50vbOAt925h86ZW5f89XunnsfzLI6pzBtYKUkXEII4E4XptgF
1eLC8qOuSwi0Gvx35Wd45Nl+hGZWNxYc5JtDvScNTTPkX7b+fbUSb4+fecDtoOJD12w3bK1l9T76
ZdZVV4eKYKh8KSjZyBZuM+HzbugDpnVjfyWLDEvgEHapi7CNDFs6PG8Agg5WzPq7ZaOLwzHl1tsZ
Cvk3TSUDt/QiZ/0pZp5ZvD+9j1uDNjCoL3acl1bEcg79OcO+nAFP8UVSaKLYjF8Gah4mEY4mT78G
SYtqTlbu9PC8ZDQzQjwBOpRNyF4djRerijhlUmiN2YuBpOYMZaRD2TfwEaZQ31ZKPAY+322+KFg2
Ut3ACuCLiqh8d3Gy7bMtIP4n9YBtYtVpm7x5rCWdc3hFv+Va5HgU9bH7qWz7s1u04Gdhk1EMedxi
XnsnG2kEiIP8gwaqJarqd1wecjbTOdCgropHG84TLT1wXJEuDigti6nUJDvILg+ZJFuYWoOqjqY7
eFRIgodEisqXulidjGB1AgWTYYrQT3l0nqhIOj9Duvhzc6OzmmKqKFb2ejVIyaJ5DoXHwLNyXKFR
tceNfQ7uoOqSDjQezGkziMaB0BzzCOyJN/ZG7OLcsGynjmv+mPhknnTTtVSiHBH7ZTT9hEbcn8hw
RX7tUYsh2Ha62Q3IQByNeYzfV+hGZCQmEH7+N9DfP5vijwzochB+NOYPrOJd1ZQH9Qh2JHQlkcvu
He+B0wfcfdTXfxCFQb6XOwEaEiEJztujGAQoLPg32XTnCNh1D3nuNPka5Bgub0t9ddPVUu3MbXSq
X+Wg64HuIBWm4Zi7QJlm4dq8Pw1nCObRuabrGE/sySvBOvdi08YdJbhlBYNqHyNgokUq77qKWmdg
Vn0Gbey+9HhVbuc/B6B8KojOe7Asuf9pLgd43bUUt1Cqxq4zqTheSKRww5PzVhdWMIejoS2GheMb
SDjWs4QxZHqGUmUYXcvFDbNZhKvifhZmw2FxjR1S7zRJicXObKf9BEWptET+P+GmilKTMWTAQdTi
+rCainfR92tIqRur0o3+VIw8eGikPIX++dwS3/FGrgLdGM3Nc8Ni7UT5MzWzAkuRqbZF5CV2td8N
ZpuZk7SjFsarQRRAgjaReS9fC5MNY4RzyZZVd7VizDZw5DUmILBNsuZvPqExNuGz8Ai0Pxfak1+F
WRr8fX7f+wsUHD/jYpGkIJKdTT1rEZ+e5PsC/ckAz5foXYDdOS/wokoQiCA82v1fIoouc/dJfBW1
XNjsDc0gaCMJm5uufW8AqIPjNkEwVud8rwdLPRAPa86moNp/t/dpEEPn8uKoTBFl+AL5MCwhpzLL
EKepQlXtXZBbbOVP+5pc1muBuOsVTSvCyHdXon0gXztaUPcab+JQX+flOk33qcaW6VlnPhDttyCF
9C/qMfrAnbfESfFGKHpFckizSPi5mfXR9b3ZkdEjhPYlBwNGsrC1XOV74Tuyv8riVN/1NhN3RCIE
yy9lyu/cYApGbCe2+et3dsUR2Vm59R111Cs7UpA+nwu5XExxFMcmtc5Skv7+OHrkrWw80ZXN/zlh
KyG9LOFUGRpLvfKDQI1JyRP2LFDZEnXIuugI1HfMzdKXlpmTB0865mziL0ei3U7HXoRze1w5SUGu
KWqGZH7VFbM/tu4//VfFGYXRe/AnYJDjMRK4DnlzAG1O4BbMuUF5HyAHAvHHMHrwy8vGZBjPz2wq
0hRMbZ2A8aBJPwJxmOo45b0bmcLGCseOe67cNzVah5mXtGCb+UtekpUojq3x0VWZD49Cb/ClJKZE
jc70oANIxx/8NLR33rAl5WihagIp3Hw9hSIne8SbjJVGROkqe2Pfk82pRfYhZ613IQ02QIjS4xVJ
+VCCq20repwPQwkDJO+zr6gLsuy5aigKyMbiSJ5KItd/UPw+pn3jDEcWAvn7/I5LwkT1aF0xmic/
pHpmJ+BaEoJMAYOW6vvwnXDlkf7QjlJLwdOO6UU4lwLKUzeDfrJc4NbVD+AxGShGNjvwf5Nb5ZMQ
R+FwWQJVgSm67idNYEezDT+hOrKAd3EFOB2wZVRv1bhnnJE5WfkKJ1frXb3PXH0Q3D0B12PAN0eX
7qpAz/Jwge2J7/nysiFoMbHqo3J57NCE5aqXTg5RmR3xa4F++Gua9N90nvdGGGuuUgp8TALh8Vbb
TKDgcqaHLaXRHtUQznliumYSurmBNrC0O2BVA2CmeBlNORIKf7VfdEAQD742uR6hnRfrfeZD1kYY
cnwsZlL5c6GWatxdX2HnEZfPaudUcbo782PUKyqvfCinfu8IHiYChD8GIz/bIbSG/7drxLAXDi4f
cSCOPvNo28B+lbiyrrhrnA1C63yrN/N5fvjrqmOAISI+C30r4DLaJOUZJvfak+uQmwhESC1cmXSq
oNm5Og6Isk/2hzfvmvnCJAbDmShYDqnkUWkpejc86wGP8b5QZ5qbZqaxfYV0O3jYmvTs6B1JVW6S
E3DX5qwKHWgCt5mqv576g762o6S6+dMfaeWBk++1UgPU/+ill2Q5w4b9m0tbXGENPYaJ4jWgtAL7
Q0sTb6owc+WMn8k6ff4wOTBLyxPg3Vw7R8wvP9s21u9+qOCzERISdytVBbWOjNbftPkPE6cDsvVr
Ulqt2Gzb16AQjCzvYi6xDH8hbNSU0xt6mt9WkhhrkyrA7gZbmnM2QXX0P3XzfOA1gr5VjsdLuVls
vjH3qVAE/iuT28T7ALSf7aYGx/ylpqLGVMqxm9YHgZcaAlB5mCAWnsu+Z5s1fg8z2gB5fehLTZRC
x+TAa5z7+QmbYWC2kWN6GBi9LQmiJXjdOHB2RFL43/GgsMlUz61hKUF0CC9mFlf9gdfafAjycGFf
421U/0Agfvggz2ndeV9hnzPQYcCEOoILaRGlqyuIHgI4Brs2+S71DzTdEimMgzSXwgxq6Xs1SYRl
w/X5cfIU6fsH4TtXrk9fGn6JFWbwR+djlW18UBSIib0KgHRgtBp0/zme8Ww0e+rgs+rf17CFo0ki
9X7+WcBIwgugvRNW+SxNTj7bOHjxZTSK4yRdnOZ3eOVRHDPWQmirGXpHrSl8iHTlfo36jcTGQZVP
mV0m114NllBESi9g+XCGg64FgGFxM3+OX9989tFbDKk+vQdk3opFDUKkF79/o6CMjmJP80e1FC/D
c/9k+h5+/bsaanwsCpVlsZbzPAMf+vLhSEJhJSg8Kkvk1U2AUYiMQU1Ydg81/MvbReiWPSFKaJKd
4oIlZ7knMGcnsGqTYrSfhM58Y40Dr8efl6s9SZkDaIkbyAEFhb2vZvRxJlFluy+jQtr/ND7hKtQM
L7aLoYepFSCLfvcFCC334kM1LltR9g1G/TtsLAXWeYKq+bEOU5JxxFaCX0v2MOLJRkXZqmdYciiX
j80vugKGw0BrKaqdIPyeyq2HBNMr7xQa8KAVHAzc0TK50aF7sSTZwWXnNbeA8g5KNKtgPGoBRD8/
cOqvJqT0GE36SkCtYRL9k3MfydZ4b2Tiffywym2PBEq/ryGe2sPX+TBv9sE3G4br0TklS6SSKiyo
CCdPwwubfA73wp1ap7n2SEQIHPvMTscE2w6FdREAQmY5GDxvsHwRz4gqAj/Xx9Rt/3HjTA4L44AA
J8sXVZW3IkV/wZkSUQvSP+kw7cV4Zz8sr4V8P55IoleR9P8bt8xQ4nQWyj3x/ZB3Nt/+scgFCYIE
mJ3Lh39O2oI9PezMXoU1cEBp42n7ME6/hZr3Qf5WvEO/rGCuUZl0qHlXk5C6ytllIbe3iOtTGCTz
AZuP1tXha1/01QWapocH8EgCn1yVueJ8f6bx41hGPET7FwI80yI9TpaekXYOLqBEtiQewQkwMhbu
S7hf+mJS+CSAelZZMEjFv61OCJq/qJxbquhSvVpR+5W5N3c1XYx+nGfIFd6bNrVgBT2Ethb7mf8M
B/gCTGprOukmX/WMlWaqYRi9h2p1QPekNm8l0qDHewcqOHOkQp4SSFyX/eIWtF2D3rba/vSN6IH9
zmuIMDZfkV31t/PWDTKkNDKAha6HKlbzmQt3pW2CXoVLOWZHG6Lxiq7WVXZXwJ5ufy19zQ3GuOhs
Z6PN20waatz/rbCCQJ9jJUx7lB/yGHgf08gI+kSnTDdb89M/4ZDyiMDlpROWv0yEbSQEQ08QqT6m
LU7jg2UjIfFxZTAZAbYjRlGoMlplVN0axdZAVi5Wke9YLPq60e3JfhkF9i+u82cku2nBYh4cjC/g
1vyuQQzLOZLpbGhmfA4Fa7siTM5JWNxYxVV/KPd1n2gEx6pSTfY8O0KnRsK7+Coyev93//RkcB/7
lyr4og7q4u/a51yaI91SRadOe5SuF3NaiDWjMRHxoX740oPDEm/q1ETTAokdH0DVHe4jufze3HyV
Hn6+/p+jnWyuksYzJvPxqiQ+igeHKQwhnp75RwWs2nL+xuO6YvWDuMpPVCOmBgpGpF/Wyca0IedC
KgsPXtrA4e11geRHsKq3J0AX2oxBG7Q9dHu40HFh/o3yavfBk1nHy0ZGwo1GvCiNHSFLY/XK39bD
TcnTnVUFJHGDL/wAiOq1mgXiarAdCetYjIAYn1k3E7hMjpJWVdwXrIXR3hPKPKSHX2k1Ch/dmzdc
CRq5VEEgM7JQF4itJHu1DJE0yz41oKbi+ZYmvxPes1ciA1kUvPKpybSHL/IAXR0yyPmJskziUDFu
ZeNtvLRJKKGjiC9WLaNcQQ2rf7knHAak/0BzG+nr/ZwSKpIwCCc9DwaxdmtxnyCw+tzQN5jX5/J3
rEqBHx5WbVF8DsRzNv2GVggQiUuHPR6kzLQJKcKun0dvuZNJq6kGS9iy/Mqfo8T9rY5FiShZtS4E
/6MiRGeTE3cEHOmwHwj0fcn0y3nQE0lpeRYsjqyqLC/h9uxy5/bOkxOVuON4+lgK/FqUnNJ8kdPs
bI3Hv2tiui/J7qi91q8jKuCQXsTngv1WiXb6rGHMzNoI25j/iOG/FrFutkjgPgu0pNA7B7ja/WWM
B9i74M1o8DQE5B7aolXnuQNkZHKNYhSDEjU+70Km3mk/B5IDtF2QCcYNWU/haylB3o67vUGxFTpR
rg5bKbenwnFZ1fFX0lBmXBZMK7Oi09h3QkmkCtLtbXaVcpyI4gIZflKzyYcZ8igTFd67bRzM1XNt
WODPRmT1BbEwhOk/bRA2ayv+SDsineM8IIVQkRYUwufbayTZyuXeT+2c9uEEeZ4odnednQ6waBCL
c7F19kgdiSRJV32wNffkOV22lekTWtDu3qoHDqkHI0RoREmD5EHIQWcFXhYO9Z7Y5xyNFZ4if19A
1qGDWRS/wQd9Q2QJndpin6xkOg8GBPR7Cv0blbEBL5OfS/UdQcgT9b0lcuORTvRqODf9Ta62PGCg
T7l44XO77fRNEewsRpzOKJc90pzKdXVq8ZlhU2H6KfEc9j2JZn9kk5MY7lFo28ZMKVx+IoM+p4V4
Sa+PTfo7OGfGrNXA5DdIwqZZr7YE6yfMZ8Q/fdVTPqHO5LNofD08GCYjMiDC55Ieyq2LLsA/8eCC
YN9wL+WI1Kq7TIP9qe5lk6sibHlhPz1HQY1Y/4Er9p/ZigA0U9xygwrjKmaiod/qqi6tciPZN4sU
1s54rwqAK3ywCQ7O+hDPsT4Br3aebI7KQT9ujYjHF/KmuIz/aoBcxAp/xPR9gwS5di/B3VyLAQTR
txkoW0QQmEak4BJe8n7zQ3+GvfYjAr+61w2PgCu97Xx7DbpK689VgYlZWv2GuBDewYsE9aqlxl03
pMn0F/6cccGZyOwgi0XOgOWtYYhPQ20FX8cr2UncCf7qdC2Xns6uULC9Q30rJ6DwPnLWtImUYQwD
0awPAWZoWS2/miV9CRVu5/7Cht5eBf5utfXzcKf0mut2e9RKQiz/lgJMJiocEKIV0GiO/6CGWUmB
P/WZaafcNUhLAbigvSHCWS9vpZXhor7ZBvXFSVOLK/Sl4BCdUvKrGiWFV2apawrwDLfZvZ0EdZdT
5YmGaTDcSssjC8kxRmIbIdnmxeXHZNxwSpxZ1SUMRyn10gYJPIgXsYChFB3B8B0Jadz1qXcm4cTp
k2+l8hvDuBwIdCf0IImfFoZMnrt6Np4Gq4b0UNjV7GaU/so6wI+jnnHZuKLJMURZ3NMWyYABu8xX
/VGx8h+fCxxzJWmtr9pfQwwVKgPvkzCgOKLfMGrU09yN19MEf1CedzGFyWDKgmFqJAVI+SFAumtx
8WEAvUQlBJ7mjZ0o7iPmZ5UyjkeolKoeR+O0RynDpvfe5YnYkuUv4YRti4U85e6L3bGkAHO90qYs
EZom8GDzkTif2+HDnVj+usz+Sd4iCuuXuchBt2gz
`protect end_protected

