

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e2VQd/JkHeEe4mr54dnWM16g2399v0mhU+1ZT8oWFJUJCdyMu4+q7oH8u3QZmAK8Rcnxp+2SrcpO
m9pYEpjU5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e4k3IaAaNAlNFkvmIoO4qJK1gZoF/VExyr/L2EnpV2zV6AVGzYp83eEX/q7O167vsBLgWYGwRFsP
yi4sfYl5lIuJf2EmeuOEauZwESJuKd6uc1klxaADn7CdEBB8W/rBSaqjDoVCuWxTpK1As0yCX9BZ
RkI2Kfe6mL0Xs6sQpTo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IbtPpkhRONJmgAFUIssZ5lSlLGn92JCOk3a/5TU0b+nZGM9b2fJWwwoGbY/OL/gG3eCzPWC2mZ4Q
yQHVXagA0da67WaW3vnZMDAL5frakXXSrA2s87T1FAjqJLmQF7Unh7546PBsqL3OQpKa5tE2Qt9p
EVAvDXDTdLcKhvmEciakrtXwSTthowcA9uRLxUPk8f0EUO4CTfkvluf6ycg5PO6pxfumZFj/0WGs
vgTtbHeVNSCwdx/DPIPQrx/2AfRxSZujtPeD86jE5AaqkaHPmVodviYONlhtWin/aHIYEIBELmjP
OfgBpo4y7pdG2K9gwF+I76hLDXYgXkS1E3SJtA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jYNHOo/XTSvo0oBfqkgIM6041mVNycidzkShFA7DjL3O3k+3PIOaz1gxN4XAJeVyBTFZGUu9UNpb
lLYIK0sXIcMhzqD/csYXqYD72yk+XSADEYXGdJxFpJfGamCnDtSyBZIo7PBWUINe2Do8h7OVRMiK
aS7bCOSSci8hvDiZE80=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZHkoK3izETxxNJyR8GdmtFOEPHd8+4rIb//gPmmS/L1BfMiycMWs4JZ0IF56rYeBFqrbQeNtD9Va
BKnGrhYVPTrxcjX5+asuKlu46CBX/iIHEmzrKpr/LAUFIgJgUQFePcXNFNPZEAJsYZmhuSrzc2sY
05sJlmShgR0KVQTbBUWl7mt1DY93aBIhdhmiaHpULcmSxpAU6go9uAbU3jUM00ZMhYA25YYv6AEb
gg84k1+xXW4rmxbK8BWXOVrPImvNZoYgt8qi2fdGpgMvgaoBCq3Rxxbaiti+CXpWZdQ5NbjWArUp
y47h8RokwLA8qG0K8OF44wzHSSkCcalfq4pG0w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26336)
`protect data_block
nWilA0E3yfTYmg/JFefSfscUKBcsZfRLCzceZlBe9xN4aPzJWM1e2xanIDW/5187u8upx9jmwWa6
C1X1NpIYFh0rkXBOelG8Ba664NWJlm7QBO1Ds0UHmpBYJV5+xYaeUxs8rLfKqP2PfwS/9dqoid0e
7vx2VL8QvgSMUTUAUu1sBowj5M6i8HOWMPr+JH68fOGi4Pfwj+/UhuhDL8CGeLy6ftaA/jpYR+Zd
wauti5VR5ZKoHyeUhc3MvGGPf1zp+qzX8YBtc8w3Y89TYeZoEiKEgZkqRCIXr9BN7WANCFHj83Wf
C7coXy2RvlMl6TZ0Eg4rgf3QbTkEMWdUqaKi+OBQVZ9wLJnAVX9gVMonrEomC3ULaMn35Li/dZlb
wfOaIKpz6Dq5Q7Im1HDHRPwl/Eh1GhRSvTIDujXMdlBygHaj3mPtcOM38jPTQKtH1cinyWv/M7ee
JTS7teQgLFwLlbvibFASU4aCsAoTP/kUowH5Sa/c5I59q3ePpWnKiYGFmUh76UgFtcAk0XPOQlMk
UhbrKSwL0MCyM4dT/67pLBRM5Qdt1O8y9zAwypZ5gDKTukywGmy8qrMxs74rg36mUEyNjTnPm85b
u28GQz1pq/uwocEjP9GwEhQAF9wWC8BTYOPXJVBBEYrIWDWKuF/DCZLaQCDa8WJ8kUpzd/aPjLwz
65uKqP+e7BdVUDgAHpmxvLkn6SNBbsVJm72VlG/WcEB2e4To1vfa66mWDTenMIuR4Knfo9HX2L3D
3NgHznKJQVdMZ5/olxJbyt8/JuVkF8lbOssQOeV1pZcxSlFIOnmM5pIOANET5U6MbffaOXwpjWe+
qVgUCv+6RQwPlqinXigeQkFLfB9jiEiznthePCQS92dBUgyCLUrU3Jqzy4Xdsgq+mVNtaYlRVQR4
bZQ/41XBSSMbQgxoUhTmAgMAzsNrU5O4KMHG918VbAQhMoAoGFkPYIIwtwgJzR56eGKwE8Zccouf
QEcCIQm/Zkj3JvTBr5bUlqyvtWOtW4raRshtW5YLXXZtwmPrb6FHwO2hwWx3CMfxstgHcnWWVRj/
HQxxTgBF8/JEdKjVE1gjVKIFoIS7+gRA2T+oRd4B/2TI/0+7SXhazfT+aytRF27EKO+n49OqZBx2
bmXvDFQkOp8x3y//ZlqNIO5DjzA8t9ovhmG7HPlJ0liM05A1FNcMw+LD3Vw6h13DbLgWfCfXn94b
Datywy5/z0y4huOvz2e+jLih9jWTWzi34/pSlG8WE1N//R55uaHf0IkCUIW8dOsmzS1V8QxVyfiw
LSnJ19SYpYWrVr/xyLLfUkXJWV65dTy3anaW6Ohvcctk/ojJyuPqvHduJ0IcVmy0g5Oj1XrVez2F
Cvr82CnD9uOUESZtlgasyM85mW5CV9n1e/nldaKcwg2MSDNNh4B1Dm2jigYn36AB6sQ3bpYozp/1
JloXnxgz+vl+8VgRwj5YVW/QlJQWxqr2QLT8+T4EJDA5rRg5QCQqobpYVghRddKZW36jNNjcrELQ
MFHGdzH2HqlpLCuXeDEf429YLZyCeGU8Z86ZClouPFSaIrVgvcljsDi1heVZs35wKJUhgbC+T40g
ImnGGS/tytqiuJlz/Xe4ySIj5gLI5EhQk/764enid5B2jdaIk0JY0rslWm6nGbPFQcSgt+tCPT48
LGnymbp3HBFxDRHN63AtoTikKF5R4o+rPTlW+AzIXl/ekrvbX4+XBxzkXnr2PoNz6Q/IykCZKg6o
wXbmL1l3cTUVSZoTzxo2Y3LrKCHcQ13kd6pT8AGqG6S8B/UsxyFD8HW+f2LwnLNFPT6iSD094IR0
jhMtWA4470WP0nb0tgn29D/f7TukwRmPwYoNVp3rBqBavlgoSYTiyGKfcniAeH+ehpacTc7TSG24
SLtW/aDG+6x0lvK+sINDE/S4Glr+FYKiG9hVeeeDlmyny/ETKK7PsX1Q8gyz0LAAaiaJyEqTDyvt
S7lneCXebX5q5asYPLmwqsvq6duawj4NOm87uPBA3buPbq1ZtKqTbCF96Ux7mKKnDGd6cjBZl9t/
BIAsAzYA1VTQxSdG/6A24uQH/ANruPIPeQcAQodOww03AufBP8nGcsWbOK6n6YpIO/ClLvJGf9J7
mEW2gwZnzbprnAwIIxr8ZhfaLRzpqyPUZDn21OXF1AC3tm61BNr71e/fUw6sC0AMIpWOaj6a+ncP
JBg72DAUENPZBjejDev/dim+BlWhoJTeyLq5kUBlFtocSnJ9iJ35ZG0M0wfw300DVhNH0JSsplvf
y2YYoHC9gJJFx0/er2bH90BHascQjsCy2zVPJOehBpCU39rDwoVcqYwUqIW6+u2cV1wiszgrQWl8
k76Duw8IQ3vHArnFrP84Xo2VsZvhsQ1b9WFlaoxmuJj65EeIXT44cDgyIAI5JtHLbd9uBlFQXoZ4
meYO2Eczuc2+hBlxkUpunMtg6QmefsD+cgpdncVDLE5y5eYqd/0gQHKbvcla5R9auRDTq0YjwMzD
zLXGpkEfKj1FlBb+hydUzSohC64w84jgXZ9El8WEuA0+1R3vjFG2bogtgd9azDSXCEfl0fJ4cJAG
FRu+w4faaI8W/VOiPbWYSzDVvGQf6HnhP7QlVC3545xdAocr72o2qSTAuHFeoRmRe9MJ5gYKOUsD
ToPb8OpENPWLos8QwCBJ3Oph4xl/Jpd+DXec4owFMB+2BXlG2wneZOkawMCQi+X2Q7i2lKuJ0TIw
xoXpdCVKaonNydgLEMMUZIKrliX220dQcbs0X6o7aBA6yMhvvDfnbxTThewZHuRxd3qJoQ/cAsaP
gWE/bnx6hAhhTWuDAPFBcrMCQKeJSLgoCDjM0a7fZiu2CtHOl89SCtjBMFSZlTMKC2YmMC+CALDt
V9tkzrXmDaovpckoFUAMk5+mMMHmv/PNNkDyL5I33UYnptM2FFi5dMbQ8fxD8gvOApJGOTJTqAoT
uiUAxQViEOhQvmo9XYjzPD2wyaV/NmFXdiUB1py7nKZhxATqZCmUJVBkZzzomE1Vpy2/U0GvVKg2
DiHZHlS/Lk6ESkqG4HfSedBDAcsPkiKTXGFU7waYX5M3JXOsoMPdCwZ+K35aSD6WLkDyPJeN9+5R
BuefpfHck/yQNdHD13UGATxj1t3R7GjfbBBn8Npul94aQpjqowoA8jN2gfKrWCiImA6S6uZadlTo
Uq7y41X5y9bXj8kT5k91+WGHuDay2cB0DDXe1HXKWZpZbG+8bzjxBHT9CXJLiWkGiBTw9mHbelIp
YRenpbyDMDznrqJCBzHbEIeVDM2p6nnH4cZw5bNK8ghFBvJfDVdv34zX9ZN/IOGCLiAselLD6a+7
kJruIY552NUB+53qsFSZROLLkgySZo1KJYhlE9M0GOb5WGDCuwAo3WnDAMByvZigj4f1+X50Ne4z
5urR0My9QorhN5xXS2mSktEr4WlEsSwrGXx0xgHqyNNDkJxh2xRpXSoMlfDl4EUmy4UyUPVIFyYB
NGLV2FbX1ZtU7eEoqUdnGL7F30UVsxmMQ9e2okslnMC4/dL9qkhu/bkKIRKzb6lWkKqtIXKP865g
lmw8ce5Y0ewMPpiI8sxqjOIh2OQ0ohDzsR8BEnPmWaKS30ytWP/+r3s4sGGV4muvE10LOowWTM3w
BaRr4NsJsJxu23XZnwdfgSGoBgb8xVeYhGXT9HVYKFt0z4XY1rUiB6GdC5vONkjEuYOEsHoZ2R7W
360h2Qj7sBqDJFPuI6MzvPLWZ+KVWtu6JBxRMIJJRVCPCgO57gz6CFYRBtap5mM4BIn7Eyu11AZx
LUwPSsbWBYT40vpeH76rKh2qLOe4iZCLaQG+ynIRUvCxpEvGLXpWrHSM1Qb0nilcRXtDiW1Ptnj/
4FVebaGv3LVs7fLLt1sHlXrOonFDj0jamZlWZZny9ZBxQNzBITlgn8sfpAPyC7O3/eR45DYObfiP
Y+Oc1hEmd42pWAb1qnr+V7gRnBh4+1VgPpq+9E4dpmxiuWiiyOXrLd76kctIA8wlPbof4y3gGCkD
XoL3WCPk6+zYOPP2NlzCSdM57ROb5iqP77FEJSU+j8riUFjJO0rJ6hRTEGrWFSQlcb9fqxcmXoai
q4LECh15gMPg2QWX9unW8tafjj6boA9MSzZYTNh1NpV4Spf1Et6ansjFmt45zIFlZWYvOWeZDumo
PlA8WTzSB+UtlL4iFlUMD42YiC/IWnp4fktwjubJ22RUw8ElYtQcUhufXBiTXguAVb/1NWQMrE7v
VfOiaC/qlOc0yaTphYxFs/81h7CagIJ31N4K5HxfrdStHeAxMjuSdUv/1yQEhnGIS2Ny/h8K9yUP
oMnnkRLPYIvo8vMtE5nlmY1rWH3yFbvsB2BHOYsxhUid175GDhXP3HsxgLlxWSYgqdpz2j/D+7zD
5BQnVJW+e38WGTRT4TZX4FSqHSPAiQMPsYDJaK9SxZyNAhUOSVF3m//P3bbkLb3kzRVbJFN4LTfa
eVi8kSAyWzMRcdAGlUBsYr1Pz4rh77ueH/YKUMqCaUBDB+Kz/qpqPSpQNyNN1SrMPSMBv/Ue/tpm
UkpQvuaFdIzdqomkfsI9YByqSG8NUiurll5kyfubQPzYxH/NAl7HEyuiQMV+i3E8F6e310wFmLGc
SwILOGzwtbNtKtCBTE9soBYGsxNvJKrX1gFsl9M02FuSvZB21WjhII/0TdaOOoTQgxWsc/V/CzxG
tvLwTDLlC17d+T+2nf055K9c4tk119yYwwcd2pajV7pRagEryMdj75Ukkq8PPtpND0LG9n0fdXMm
ctFWAGs5oGUTlzZDIvoecNV3KHwt46IGatFL+lwAZMrRahko00yr+KeBk7yJt7OaEtmmNhDlqcGy
Ay4+yjq7WwlVvsIsK2VsZPgkeE/AM+bF2T0+Oxm3q+4pkPXVPC6X3dxjwBh5honLQaOg0RdspROJ
pO1xbVgessOVnKC8vMOnec3NqUKq9MJS5hic50CNvxBf5p0DxFIrrwebFMCRFGH5774p09kSp4Al
RNO6p9+oCDrsbfghq4svzQCjvu1NDAmnOpdym8jhRbaFvfzXof7wTiE/TiY6uus0W58W5SgfdD6o
ol++zh3HtVuj2goWfZAEK0SS//MZXEPcuEfMa/KdD/cVRClunFARRr+75ItQ7ocZ+WlbvPytfA0Y
p5lK3h6em6N2eLFSLPSey/1Khalo7DKCR7QJMe30lEi4lRo3q17qF861a0wAxkf5aewmERpB/dJ8
XHadeWuhvqUtSZWd8940xbrXvRYNT5T0O8KcU5rqgmcInrMMuSThWugUZsP+Kj6yxbh5qKoEDxOe
E/HM838eRBIthN0N99jF6IwY5hm88yCvEnFFov306iPjWgObqNPpas8cZtuvAjFYHSt7MMZKLY47
xLFudjtFwXPuqy2v7TjfDScOjkiYH7yBSzG3oHmETSf6M6Z2acf4uGjWJ8RRnz85jCVzHSS3uU2/
O353MrmoGdOWQkwzgQxLoG/Y+iTzNQBetx5QwKK+qVH0ufrvt0u8kFsCoVySjdZJ4OROv5ptxcHj
7TdI8o2hMnw3fr4HFqsAMzA4PETL2RFTIXyRfQQztd//YLYT6Ap/kplC1SMkhIXZD1GFwIhm0ypG
+VbYEo/9mfw9OStIFNEYZYDJgAuAa3ibq6EDiobP/y5XIVsnN8Jb+gWBoVEuF8gcCFA4oz7gr/WW
L1WUe8P35yArRQlVfnURB7+j3LiSP9oaGPVXJlyp40WCWOx63S5fp2mCKgfDGr45PEbBSV89DtoS
7vx63WERro4T/Vu17u/kyPQzYcpQZr8oGde9toN8wmVtsNvsfWpVW+HHe0cDTwgVCZSJADUSHbTy
QzjpSR8CQEv+V2RCQSYN1ChHGX0zxlybxNsTcpbdN/HxVSQiEX6NUmI4l9hsIOOV+6UIFrPqeYO/
gT2Yj5a4rCmSt9vhX1TMBSGRjJ794JQMAVVYzgfSHpE0s4OHmLxErZVVpgY2WJnH7MQC4G/e4Gfb
wKIBbvm1S48oFrKceXEaQjPZwgjHpAHgit1eojh/OrEXc1lmd5bxHIC/NV1qe7W2HJdk0P7GjOyI
hiq56bKUdnS291gcgsSZ7kU+6Dxbxu+DmyZgRSe8/LOXmFzdNaRCuSBgXQGl9GlWMMxOdWOVAs1L
FgrpaGl60qNmfD9+Xwi4ntFxjo/L1TfhnKKPWXizLc7DpUVt8nE3y/yN/BFiyOVAssmH9kVkD3u/
fE1c7UNheTzik+md3xnVR1QIkzg94xtJ0RIDCWfTn72Dwgrh9cFYNCymHIFy1f558QuVclO+harY
3O4GpX1SvKgrOqQyQLxCKGqAHuxoUzVn6m6YSY3XijGka6DNbS66Hme9Q42JDhgSg8b8iRFswp8K
02o0BuCteegNM3W+TnffzSuSCh1+mDqlsspjuHcTqW6V28C2SlxaLGB8wYFTkMiLXVgbhp8bUdmh
BEKsBV1le8aF+CHCNXASAiuzc2P5ZZ8UzRH96jcCYC6O39VCEcJ1WJtgaHjx8pSpVinfVDsYRlm9
nemAEa2/gUI88dKIXLjWetzSCJb9mSiP3vYjFTSb0uDeo1eA45w4YykyhEHk0w03ChaO5rvULjIG
Bg8xNB5vczi1Nf+ppaB9Xkz6oxGSbf+rm7I95dHOwPmvoBLIGKRBTnG7KDgFSa5ZiwjualGla856
OCjCZJmJIrHhLywFk7Rb2+fW4DGPxNu9RruO4eRfCRlL/Vun2Pc2meMDYd3JZD+RJsmv1pjV7O2+
t8fGz0nfBHZL0XlAAa7BsxFdf/brCjJBABZav/XH0Fw2kgmgxIWP4kRcYs4Mzx6ZiPtt/qK7c4CS
+ILKo1h+abmkcfYsSmLIeDMv6zZnca0nG+k3i+TauXPcwbvo0/36pUc7h9TedyWvgP3Vn2xtaNcJ
CveXTfgbngv+oIcMcFz8cEPbAF2ulWWge9DwLhnbry5Y2xf3rUsMkgK44Re+9wUAZSiSju+VFa3N
VkvqsuNt/LzT13EIrUR7DwFheWZxzDsNooigr0/i7JtlOisPUAmmO8ShI1Lo72sOeC4dvoG2wRfk
thW1g3Rv4zr3hgpEwL9v3iKgjfGQ0ArWY6loNC0gpDC+haU+vHavX/Md1n/4JXc4WlSi1jQrmajL
IeWh+tqi9/QZ8zIe0h16sYwSJI8PLdMuzQ6ijFJp+S0b+jIPE6nEDYT6vJwAxH4kmUyNUJt+L5dZ
5nZ3dLnajczxjbe+UWVAZ/hGPhxdycirogmFtJkaGqgq/ZbYdZppZZbTyhnPEixK+rtzG4p0dBO6
/LK2OidZ1geWO8cjnr/BdfWVnpMSv9uLY9LZJE1b0xTdtRdvqWlFzgLeF0sAeHbK7vtHjIIiUOpY
dNiMZv1xDCqqj06+PoReJYOk70XH2F/Hc1qsnmwvyJNOKXS+/Zj8uug3DW/us045oUvoO0xBe1+l
V86B4VeKBY+CuHM5Rgw9rH2yP/9UcyoSfOqqKCVxKN4PEzFdZJiWtOdvi7JSDrNAx4FuENFeGgYm
De7Tv/Ta+Gh55yIlf4zEz4FDxWVeJmNpES+lTvAsrnnFEiHoyig+x5kR5NOFOTOKbOUJ8BI7AG2F
H6utTAGWOIsff8NYEQuYgmFxsBSxbUtgV0IWslnBYB7JwhEd0CbP8cYsxRrz+DgC7Xc1tMYjU2NF
Lxh5F1Mx0wcYveaz2o9gYphsMM8Jg3+qcDNuhlOtTrbLpN4fosIq+/0viRM1IFaYxWFR7I9wQYxF
WH6jeaYPhm8FMoeGsowtsFJ4KJ7NX0SKnmj/x2s4fvA69g5Fx2mFGTBFEWrt2I01S8mlf/BsurJ+
mz98hq/xqppD9PYSlFd4ZxaEOB2IICndR/5lrqqDzXLSheikyRKJw+KiJuXupkRuNItkQxtZauAa
zzhyOK9npY8ZbdDTMHBFBgBorNURbB9BbGDrPqQhHrH3JsKizpxXlVTp89d0u1TzwaYg85amh5VS
6UvPbZmoVxe2eYsamauqx61y1Ja89SVhUnQVSSo/SdnJbd1WLdwVRc4I+I+KC8fqHSMWBgWMl8sX
3Ck+4NRYuTKslLnt3/r4+YTNspbAkh/HYcTiBVO8qQberk/A603S7AjI8kPOYh5YZ4xcXnemSeXK
lUOpyK3ei9f8/o+UITYAAkAL0A4+dsFNemovNZzkfXVBTwcd2tnu09zlwR8diRNxvFDLJ2ECtBDF
G1Q+K8zV/kqO8K96zgI2TAurcyuwPV4sFzxZzykGJQVvmPSSQ1f3hF9HudRQldRWz/iwF9hRGWFH
p945CYUlssxy7zAwxjPXq75GA4l9m2v/Uga6fIZaGHIYKdebXhrldl1WXFix/9spSgeQCXE0ApHG
iExnVnZXfXI+mqEQHyMkSvklWtBv79gv3o2H3v7Ft4iwwhULK+FdkGxeIqjqmJYJyr7kPRaRBylk
qcAYpCTj1yg6nb9+tmB9lQRfJlaCtKq2mRoQCVNggaIe7nziNgvAlNwmyWnNVXhcL3o8MYyKovFO
Bn6awIMJnYqYcf3JcJ1HCIwivHaWt/0I6gduF/t9F1YP+Vn6v9ltvbKmiAHQYVJdsaqbspjAp8Mm
SOEPAHRVPIS3pQZknuJZFMWaV3llQ4DXRZDbwVgyvdwayMWvMNwujnRocGAyxSzatfjxN6NYd53d
jJXsRgVuY5lNZfCUxOVzK4y9XiyknxbrUuOJkaQQUEtTo5CJ2xXLkydUAXgqErhhcH2gSIyPyRpr
Egw00Ew31Ijjfyq9qIwzxMGZ1KEKfcjpL+qqqFu8qsfyj96F2o1GdOWil+oaMClrFJkiaEfx14sv
wW844X2zbqxzcxnGZ38A6K/LhbK06Rj86SESlmleNRs9X1TT3BejL3w+9nk5yb0pwt/R6PVgtCu0
6kZUsm5j10GbETaTlk4T2RU/iH/wAXpQzcMs/FCPLCRO7lR5Xu9ATW8X/qhTwGFLE+f2mi1NcaO2
W234KbbsXdF7xiDuw9PN5Y6oZuVQaxdIx89ybUR9nEw9ej/HswLLRDc31szrjrlfDnBe0v1wSJsi
sNQY6rEwdCTS61/ENrYd4HiOz2izJ3alCu7XLeou1wnxbjOEdMlZP0HTUFgp6nU84zG5EdYRJkcf
YkjyAoxNmvYQ0KtlKNQJc/C5M9nu7dq57gLHzTAeTlYigGu5m5ZSwucL7Qo511DuWotK6AOUEiv8
2FRYZj+EtjSTK67f0sXMuhWZ4aAThIToW3UqhPPuM8ZR6I5xaqSPiZnPNKsQdw4NWebVzAUBC/t5
4yNuZy0Y4H8CIFje2AI2gwc0IAoPhMZ/qAfnyzF/m/Mg7am0NEQmNhY48QPCx3iebfJrxQiT/lWR
W20q0SEkFDQMyd2eVmuntbqn36UN6YTi1GbdRykH2jTA9luomH/JFMvjW9nHR/gOpaSIhP3Nnte0
6biVHE2+zLLlDkGSYNmldiNNzVKM7B3ZyCfwmKn05l+P00wkWyuipdRtM/zFUQMz1z2Np5FaSpyF
NVJ/1fIbCgL4AjQHr19DsnWhffeO7Kw+i4gWg+poNlQVwhpQna3Igbq3jxfMxVfrVQLPH7F8y094
XCmnu/UWGj1ZHVVptf3YHbIhvUsQd85hbHnPofp2FthW6GonSzBCRtS2LPd29EG2+hG4tlssTeuT
nVrIoTdOVnYLM4Sdo51r9fpZTbiDaqyEJiJ97BRfh6P3l1c2m2PBb3OnuyvgXtCOrU27DdVdTNEy
k4kliLv6KmqH7ybaGp/9FXOoy7wMrvOORAy81n77gp53Do0BEjQhrZspvuu2HrFgNjwiYvYxeXSu
EKlZPmD3FKfsuztNzzzYjA3L6OyX7yZ5VGnNDybFSWYHBTXMaXjTEGMPmKuAcE/BozsA1bc57Rw5
PAgBkisPH/nhubaAvABmGeR/wmpCkoCx6pRFLMpeCXdbbH2ZQrcRuCNqOlvse35IYd+kiBrSHrJh
9v5PT4bBN9i1jfMhUmA6KKCS0/fjlvHBSZgQRs/VhC3x1FDLRmRrI2pgFhvmTycdO119ESr5RGIJ
Miv77hoeM5A+tr+Fy0DSmK5VgBKGNnLRx7oVVHlr223S4th7w62LRfviOpsdMXsShkZvQyTowuQB
Y8DM2VKqKEiV1QIr31cJXe4F1uyKLWYNu9noLtE7SC9iltaIaYULPVywCSWbVfexaP4YV3QvNNph
6LI/RHGF+fGntRnGNKPMlry3qo8Kq4feTK1otgG3YMl8Gp9K4fTMYb1OF4ehdBkr2UuxXHCFS2ln
spR96Jkd96ZsMhRJKQkLykJngMBwn+gnuxu+B7Fav7wDYkw7/GksA3eBgFGwbpUg/WZoKawAX+cS
/TTmNnvXpH2d2llsX2/I9aXrN9SGiNe5CUv83DfOKFdWeKwGsQKsQm8PUBRLEyhyIGiRVgjEl+qp
rEHFnOdAxG0LqgMTyIH5cUGJwu8T4lqBYJt7Tur4m5NpnC3qgmb1c230++xixH0Qb1eQ17i4sUdI
xKK5TyVQg/D+8eesGnI36+2ZGY0qOzQzqIVmiO8jXxUIGbviu+FG7JMXWdFv5QeXwaCrLrUgWQqi
cxq7GOlm3Z0maPGkNYuKMGyZ6C4G5w8/pe8m8mxHFI5nHiFUq31zCVwYMLbw9L6iBgSMlm3QfjSx
HhXYm1UZw5bXgv8lz//o7wY4WgQ1NEArQ5OaoKZi3ugSyyxXn5ImdOnaebsdJhbMa3rg/w7JIxwB
vaEJQe+oK4Z2/WpGmbMaLudaj7WupeUXulqCRynDrpNEuxueDhyq9WcGSt6GyS1qTQNcxHIO11TH
1wGrCNVBG95tt313aa5Nm+6jdZCntPz0JwOEigHlqngLOEkPDwppo4X0mBsGVuOEg2us0D/jya1X
sebWwxN5KdJOtXrWxwBpb+P8tzwNgMXS03Z0+SoaDUXGm9NrFI+SRKK6t1RjVNY+Mr8kKzPjykg8
doroSmiNFbNiu+diamAtxBz0SVv7i7u1NRAa2fzBlm8rBX3ZOKryVbMHkXUU0Wb+vrkHtJrbHi6S
pOYYp9oU0oEO51zUZL+s/7OIkmBYFuHwIg03oeAHLXcjlIx6+M79E1MOoe9HlZm/AdGAUJzoJCuh
UlB30ebMRgunAEVvRxuIr/CKBsZKTAX9qqCl76QsrbTBsy0CHYsgPe4CDWV/KWmHvEw06xCpw7ed
ytMbxX6N97lMTIziDtM+lOW7YGpS8Lu1O14MV+HtJ2Ame0vYq2CVnUCtLnj+PbIZtxnuRjhjb50i
GAoDz4OAsEF39+/ZCbZorhWoCh+/H8ZbkhzqoDsboCtxiDmmeXwwNIIC661iHwa3HVPReaS6w2YK
0y6El2gMJY07kUjtYdt+gD5BDjQ15Fy5CV0TqocUoBF+423ILSvyqf5RP8kiXCy5tgmDqj7wuYnX
VU69ws5sr7UBzD5//S+l+HI7ULMpJ0wcmkSQZVWZbOlJb++DA2eI8GdM5U6fxPM5Qkirp9e4O/tn
HxvvGPyAlQUQBrCb/Sc4vYdnNRcnUijcqy6ar/0RhycwUV+mbvFgA23P5dVs5x5pw3efyGtYM9ES
g6fP0YwlX8ZbT5sKGd44F9H+5m0Dg0mQi0wltHgP35htH3gbja48cV7pSm10R0uVOz7oW9U+MprY
o5cJTBfBGiBfwyTecf72p5hZT7boWKH9H47JFd8ZGfJ/0HZCx1e9e//PgSLeYVQeCzuBgpveimAW
k5yDJWSJJdDvMBE+EWfxQOQ3tyePxeJCzkhA+2xMtfU63CKs9aUC9BTwAR05DC3yeoI9jmOjul/h
N65K7Z57N/WN1hOnVp7EbgNK99SLwVyTGlHoOyXWGvF6qpyhflcKEJA8b2RSN5UzMD1o0UI6z6p0
wjCXeuvDDNpjlFAzUtGr3gEIIqggYMvTN/MXBFCptGwqL5emjAg2P9uITjZyXRofe69RmN+HesJ7
jZRDHE/jKKANSMVGEPxkIC+4ToST7Pyr4QwCug5CyK13SL5h2GIg3M+iqx2oZ4/m8lad4PfTvhdk
uoDVLrW5c9Xnr0azwzpuaUD0jiq75WcxQCrNdeovWthCmdl2yvEgqeOgwC3lY7PyrzUzpqBh/v1b
VQCksyWuTov2CuXVwPnNJO+o5qQHICz4QzBcRPC32XCNL+CMWZSXyHqJ+FX7qdWFOaJIl9PEg/Ec
VMyWrNalGQ5WdWwOKpRqJ88GY2bopI5dtkZo+UdyMqkYlYJxDh2RLH7+jSi34b5E+6POo2PjHcuB
Xt2lDdXydeX0uqM+qmgQ29cXYM8W/cdRKBT02pqz8jiwMBsNnuSr24w//Fj5tVxa/VpLfFDuCy4E
dbmTCgxmwz3f4uqcZhIopSPN5vaXLSDn7d/L2OU8Qo0uA+suqExrrqJ4xAujyrZOn0TZI0y2sjcs
PBR80Fia/GwgGqG1mk7OxNOmmPhTeI9koWAfID/+9PRKCKIHXfT0BYTL4kCF7mYs4eumXMzPWcOz
pNPKjJLOduVxERmQbR3JRdWADZdFaw+f8CXbzZndEcS/Wyd3Rc4hBw/dfUIWjwWrJ+RoBuoFrXTD
rfoRctuyX8wxS/0D7Z2kBE3HdbhufEUKYqLcLmBQR+qiMDl42UqW+H6D19/xrpEFh5krGJCTeQbx
JMCpTda0a2CuONDA6NV8QR/66nBrxTz1qU27Q6qgxnLokqInfjxvLS4JlJan2VQOzjSmPgs61B3V
joI74loSCvV4tHc0WwzDFsGceUsmqnO8XUK3u0SPBi83jP9jNvXCDg5Zqlcn63d34dMl4jSXXdph
iYwp/Xz5iSyyXsu39PfZQgNQIY06MGGzE2wbAFa7lEYFMcaQrGpIOoGWqL0/wGc3Afc0uWnSy5yC
5YsmvbyfHh8mOVKc0NK/8GLGwZ9Dn2DORU8hac3yQOhrZgJIU5QsKEEJ3BnSU+40LesBFPHKNpy6
coDvxPHCFRhfHEQKo1ZRY2+bFb1pxQ9n+zjm21BIO+1kzyQrfJNZTOr1Dd0m7pu4Kw/ys7T8B+In
pQf3Ewc7Ri0M1cR58IhDLB2nPx2Hh9ayayp2p23Ds19Tqcs3A6IfjG4ICQcWmBMkJ+lfrh9rlhD/
ILujYXFEAUSGvtD420zGyBypLbgSbs7h3Rajl97VgOJ0+uz5TkcoG/HKNGBsCnWBQk3sqgFLt6eZ
s2CsRMhtWR1J53mxKYrNSFA1VFGZelWyaw2MHq24l/SG6uaomXqEKjaI/Du2BqyhWPnMKnToCOwI
3nMstXayHnxq327dkyvzKCe3z0XhvxSmQLZ++2o68cUiQzQIVAkJ9fB+i+sWVzDlPs6v6RDvPQTf
9tE9osMqF59rddMfFRJiduicgGjwFDY05m6vYfYos32l+wifYdha32osPpSb7LUTR7RC6fnP17kx
lO0BgMkaI0B5mQVDsEuCq2KVi7DM0EHgPFuWSNwv/+zj6qhmSApsymbtauSe74W5NwUr+OQCz06H
V32fqaH8hPH/GJyhvfnFGRrmrzNMHmPhEXyKmLr986y0mHBaMP3OqsaY7UwWrqsXgy2AaFaP+2iN
7dCBLoEqB5cjS87VudUgR7T/My1vv0RRl/oIVkcQVHp00G7fOEvoAP3pUpl6YFAJXeHXHKCSlx3+
LRfc+bOaI9bxZ3jga+kKcCiOa2tLcmMt4J84nSAWyfUW60a5reUZ7OtsiT5L9wjvRPfylX9Wcpv1
jCyuiAEh0t92mEqN9khrqoQr3lWGDB6aJ8xhiOQB8kN2blK23Nfyiw/LHm68vSbuE+opGTDuwPK9
Xfp56o00SRRM76bOaIsV1lkkRXXlUrHz8qWfdpz+SvsW3LKbcypkgAT3TzUUXNnjM86UXg56r7oe
wDRWtCXDpfiiikyvTqDzPFDfX8JjsitR8i+lXV7TdbcnTqfy74w1kmjew/xEPNyDLxtJnCXcgzSy
E3Qo1K2qcrq9bSj1Mq8O28sndPudJ9qtAnXM0c53w8opNhDJeZ1aTIjZrlPacbB6VtY77JH07r5L
gw12rMjkQFsr+of5U5nr1Z2CW7qB9NWe3sqximkh+Tz5Q2UqKaYYH6ZRTWz7w6LPZrIL5BoDwrQO
JT9Cpl/1VQFoBEsHpuzKdFrr00DTQ9lnrQFM65WrXPsqTQarfOvGJVGl0wvEsUVsubwUKRbJTMzF
33nmmL1JLH+bssQRHuPcP+CK4B4QdEzNccVqyw2HxwIRkPdMmkx80mVCp3XF5licOKp+RF1u+9da
/8lnmCi7FDlRp9mPCvJhLHfdT9C0FONWdO7JcOyItWRUUo+gIH2GL5PGK7gA5/rdO6SACT8F1c4V
lD4fRhun7tBj1pGhpSQYpT8m2HPuYCL5vMxmvfFCJHiwABrFRSwIXQU2mLVnPoBWf+bU52XEuqcN
n5bqkhujza4sEOzrIcSOYIJ0clPyhUB+6XXNczTdH+acWrfg51JsgPTqQxRl0k/xdjpePIgHxFuF
Ijx1+8Pdh+PBhWCjnagrONknaM9MFKs7KJ79G8b8vRpwPXgJ3IOEiU3+ELcMGy/QgCNyjHcfnD6L
0HqE5KAQ8Go5kAwLq7OMrprkEjVVJM6q4JHZZkri+/cJC7RCcS6N9LNiOdpeMS6gL68KEXx2AWfP
4Jgtm9m3Vp8T7cyA3SHGxs1SLLTsxtOnT45DBUFyXU+Xq3sUuzpAfKqR8oFEH58pJvLeMYfHK8Y/
1K86zaRsvFVeS6K92zbnai6au1pb0v6/kWtETxf9XK9QcwpkqZvw7gvh5MBRP7tinSuWsPY1p8Er
tEVjuNS4sQdPK5EGGh9t0zyPXwDBO1cetFjpZbDbnH2bPUmK0ciYex9YL0+X6qHS2KAtRKYtUXhl
+vKKUeRuCET+9J5ZwN/g2CQk+FxCwoGpRCDFRlhauoNWjMz3yOZAA+76DkOgXQKTIMoQjuD6v9F3
We+FW10o2h3832Vw4KkEOacZRV1gO/fKpd9ZOPkhKeIZwkVAsJTMTXH8LPJo/XFP6ITXkdwM02ee
RTJBXQCipcd5vWILECxqnhdxMM7DZ+D2cbqC2LtVHtn+q3WbooBPh45UEHp4NR0N4iFZ7y34YBsS
YwHa+b0cXHW13wR4hPMR0pnmf+KZFWNNOEztfnDxGvIMFdY9962voMxJ/9HXKCvAaYFCnL8APAQ7
ODTNc1yGqsVFjqjPAFtlRHGb1fQw4q7IELBOEXWGolektfYQeRkM9YMjUbHePjz4zB1xsnSsDcaf
+MK3fqbcxLjvDsZ/qgGDBfIT41D2oalFAIjQMusssL/S3rcH4DX4K+FJKDzukZPvzQOsM1lEKiOe
Ohs2cTPPI0eOZhsk3IS/t+iL4sqCs6odH/4UWX/yptlhVgcTjknsUc4wknnFNnN51UEGi06ddw/N
ZRaQCKL8TOaUxgJPWkI8xJ/+OgQSpoIfvCMOeBX/sx/2t97TSx6z2wHvkOqAkZCso+jvjaFjdiLz
nf1iaeH8EjtEogHLYIsdgIn0eZ9LZRQm+ajKN6SqZpPkFRw1xZ1h4rlC4DZ4898E1AyNAsa3pm+s
bTWuG3ZKt4eP8GktKQ4PdvPdr1sdOIqjWL8yjh2GX89NLLRz8xXh7lfQ5S99/RRUdLFOER034bNv
hFTTmOKlMVXdjcjNyErgr+H2ATmeFgzMYFQC0proIYmPBXeh8vDWS4AwEswM69fJ2gH0dB1oQJGa
8y9tlwqWC4kgYBfMCXumKcmC0fl8qOW5m638WdzYImIFkSoUIobdIWVhSpTVd8O5BfanOmHESuZI
h/ms/7fBHuTSmSg1pCiBzRKAut7TJqtZEcgw79vodwVYKfHKwzwBvwvqF0zlpsMbidYEml0xLkWB
v3YJyruFXEIfLCTHX9pTH7B9iHz3A9VL1G+eZOOCwoZwbG9a1Gr5g7Xw5Ivp1WHiUFXjR/mduivY
sZTFIqPSMol3ozacqF8bCD6imze7pe+ak8Qd6Skbfh4qBRE2Rr/FZcFROtnSCjPqzHmD/4yQtnF7
H1fECbfhvJJoaetP3DsMfdTStTRa66nHeXQ53guUpdar7baxs8GXYe4MpA2/vKizJGB9e4vdLEI5
kokQ0jTHaFUm4wch1LXlEqCokVZ7bXGV3dte2VLKQ5ZuwKzhNAgwbMHkOxKroYlFqvIYmS6hid2A
S6A09J25246YgazBtz9b0orMcxZNu7e5QeZlwmYmxgDfu3QJo1M9Yag1BDGb6Vrj57hJY8JKPCaH
3qNp6LRmxbika8v/32wjNRHIw9pHMN7JhATZwC5ehV+F6m8M5qq2mEdoVedeOFjloGiA+yJ3wKTv
9BwAAo8FkeaodGfZQU6S8fgZXWlQyu+t9hKwVmA+fq/IxklskdE0Y4pWrJo+L9ADcDMl7BwIpBtG
RvF3MWfNf37r/ah9uG8ZUqmLTypCrGt+a3Hgyg6jz3dn3x6GVcZWAVTmgNW74ShoPb4k6G4kwcO2
VX8asvBfY/Qc0MIUY75lQ4cvSmkOYb5Yk/+TYlgTXEr1ydHrn9dA7oRnAdemVViVu4AJOuTKHWbu
EF7D/ps8S0EhHc4MWBnAmGbs2wRP5as83sletYgPzk1JQgBP6Fs4+Wzt/7ML7Ce/rQhc5sUDfgJN
1na3Ys5wm+vw3O83DV5yycIHPpD/2WJJevHWWSZIpB/Fjp6rTIpQkmTvqaN8kTpsYR36sWJhhuAH
utznaHtBHfUpdHQzLcNTrypmq1g+DJedZL+jYvFwDYzEF2RkUP9JQ5QuUsyXavK5GZTyO9UKn/h+
f7R1/+Ajd/ddYOsXildj8Som0jW35cP3UEDuCEfHwAXJWQQN/mXgOOHuJgfal0K3ueDbbmtWbSnS
0MiLmOVFluQH2fZiJXaMtXJMuDjlEAaHgIeQSKewABvo1SvMo/fHQr5YNSkjLEt8+n/Gm0dbLXfq
nc/W/5U1TzOTKQVjaDYMib5S5wOSMerb0ycMfBchbIUkHYtnk6MOaEbbV/5oECqY7b9nIXxpsBnC
wEjxG+C+JS9o3ctgEhZcIJ21jOz83yMHrVHuTsbjvSOc+fPxk4ShOdBCSFAqyh5RP7tWC3Xs3J2/
PAhBolHrw8nmogacjD/Ay88xUKS5Lzk/+nFvjwmJFmHQsjKxK4KLVAvaBBtEBKFCB0UYkpixFuhz
ZYSjKfdCVSV6Loz+wZEzl6xGP1sT1vOoQKoX2DmNfZw/NX6k7r97kjAZkvdmZV72C3DApCrwzOaT
rhVf6JqmgsO/+JP5BvXZ+XACHAnAGu999lZB5mv6bF+tkDp2U2jojM1BBpt2cq4Jb19Sh8rAew5/
MEk8L6yv5XmamHJgfqAVYDntNYPFbK6CJYHseg0Y7j/U8JjWFPXmoO3hjChxOrXPnCD1Zv63IpwE
QHJaIV1DsScW9rXBB4Trvnz3pE4/rJy//v73lMgCkqTWpMNMFwl16HZeVd9ymU3YkIej4saFxW8p
NMdrtjFdgLZXrEDN9qriOwKn+poTwcGJbb19G6qNDdZ1B4ktyV1f9fNJd75preLady+G4QZVERGf
AF4pgVzi/A66noox9niOGxEeourKN2Q9TrfSiCnrrx0BJtl5UDtcll/Dfi4xGNqMPwU78oBtJoeJ
7fyXO8fw45RJpqMrUNSvkXjpgXviYMPy29HgLUk8Xpwyj2TLFzaZNVAqhXsJTx3qsPGsoOU7DsBU
FFvX0AoC2a1IhhBpmYmxb2WCntMDFkJ5kNwFWLekDhnUlR3Z19bTEs0MEjq5BSRpox7LlysBUMhk
x+6FfMWSaJ+X2sasHNJT25NaZT8j5nqtiPy04RkqiRq3eTH5yNNdxQz6BIg+s2BpIOhYu6htk+zM
dyh2Jld0r4VMNG7iYp5NcAYfpHC2eRBTgyna+gn0RnmmzMnXBOJgSZV58mFxF4mTk9R6Jwe/kOPZ
9Ge+B/bsVC3LMefMKajCgJTDWi2kmaPCIGkU4mbK8Lxxhmu5cQqWlSfXIKkq9lS81C3lEgqOnIfc
3e2B6veoM5LJBDstLlJa5HwJLPPZpZKwR4Oxius1Xg8f/eFS4OB/eKYvGtcpfkaxU4/WpXD/lpPS
BIUomWmezcnR4yaW+sufMtVIQyCK5F4xcYhMv2XuD9En9Z6ExhoSE3Y42S/sftFdsVK/C/hTKbVd
baS0+4uHYkawGbT/iodlw8siY382O8TqvFbgDEsDAkPHVmDR8eBAKuoI3FjzGCqB5mSVTeq7gPIY
ctoy3YoetjIdC+qLSWMQfOhKuU0AF7IlI6t36+Nueh9wIXYHN7h0Vn+aAQvx0SGylSfLAaC1bh1l
GYPExG7RfYl2eR5a7LmVFUlbHLbuuB8JqzpTrnX3rkYO1WgTQx8/KkJCkX4EuaUF+V/o6dmHdWsh
vxeJsowlFOGzK5to2UUB37HnQw8jiKoMTCw+llMVIMH3mSVXtXfpSHn8x+6lwKOzaYqoXYZxmXZe
ZFM5ZHxFONMEsitc4GYp/YyM5HTZsg8X+pBf0MRTzoLQeIollvNslZfXhTGLWEmwoSaYd7f8Ccle
1gEjBOCVWwMaYhbUTfuLiqQSpyoJwrcEuFID8TmZ5ESgZJrHC6cwfQVGNHAK8UfbtnbMEiy52C/4
pHkY8jx4m6qTw4WYO/168jYea7oTd/KUpU2Eo/PaVrOFpcFeIrtLGantXkzfCaFo9lCQN+5EOIBE
0yIs7v9ukgKKDLnBom5P3b6qE0xO++/dzjR8aWRQgkYGWjaXmJdwa19ZSiYyct702Vy9F/7oxoOO
oiOXlDto6x9efDxd+tMB6OwQhKwQr3ukdC0jBB3P1tyWDXGyurPG0OUGirmVt4IxOdSAg+whxnwd
1wmbZgEX2tnydWRfurTdzkhlQrG78NvXkYX+T29DdVn8P3VYqf937snTzzgGJuNzriwvYteZCYm0
biuQlQLP5F8L4PKIQQ2IonXqTVdy+CsYRi/wIv1bnVKzAFoE3oY6zaLwrC7281hDkOQ/aQ0SglmD
jkSGqW5IOouG87o2If3sqcTPAUQH+OlRqCPxjmTC3mBN2TQvBldlIU6qMr01sVOgQj+bU2wiyxwi
lykvRAtRk6laYhye+7AV0QwXVvyd13jso4JaMMYULgm9vxeqFXdg+YsIjwLLJkrpPvophntzeFu/
biBSqTjIeMahMeljGxW82NkHJGRk6nvqMzpAtqz869L1VoxC3z+P9DiFIToCqBHA/zKrDBL8s+D2
e2YBGIZAtf02QfrxxFr2ve6w+hWWMYK2R+kqaYzQcTJ4gYaIyTX7Fo1hUif2x5mUbK7ZKK9GZBfZ
1eO/MnyB9aGv2pLr8/xdLOtSoxUdF9zb21wQDDVQp8D/AtT0XH1LruY3wuO3TK5WblerNj/t9Vv4
AvYrEsS797LTcnQDZqqdwXT/h0qNAph/bgrxp+WdmGHH/mmwsTbCiJCU19zgrBaFDt++nDx7olje
uaX6YguKvgjEMvf5BZIzdg9BGZje2IfRygn9Yk4Xqwgm4Gfmnu76TisfzqS/sjhafHBsKscKWn+1
jWWxxf95u8Tuh/c1+0AwhKPwW2tdeCnWTG2WCAwTv8b7PH2mPyZAkVP+C1rTcjpGmezMhNZxwFye
Iz6BHFKN6QFhZ+OFwGVrRDEJ+Z///1NouPHmgxGZBRsuINrVZyyT5P6aEOtNa/u8TRG2GJAM/o+v
t1H994tX6ZYzyg43uLSCixMRua3C2SSqbj7qJnZcVyMQJMOyqy1CYzHZWh8FNRriBHCYUAa1QJeN
QMyN7g9c/Owex6td7T/Z6W06fvmtSJBlAiL8B+uBtnO9HRRMZej/I2n1I8KE09UO6m2hw6MEeXiP
8ow4kPABuKoYY/Uqh+aEsKg36D6Hiyk/p/y/LAfcYzI54n7GeS5gMsCxWzX4pBx1+xgR/2DxkDnm
MaL1iYJcUEYaQjHRjQwHy+QNIjQnOwpAZ65NjTwGdcJi96CTu/QaSloSPFOKxxO0JzVQtrsKhfHz
FaV43JKiWmE3bRrayfQW3gelNRudyRjFB7qx9jveYivtTrWKXJSPPDFckKb4VZxvFzYK3QDLJzCX
+9wMs9l/d5t96yfHy/s16xD6lT2yOLMs8TB7LHMTydxJ33Wjikhj+zb2C1zsW3q2OOenlk6BQDPz
UCYgbzFFwsQkhshssBW4FA+E8mXgO3H9shRSJam8ch1+F+d3fzHz/Bl/1SBSPOpb53OurcB/KyQo
5YsoXHz3X8v5HPe+XudrH9TkRcEW3D/WCKAUofRRVYp6lr00QLFw3wA98yyWWRidsWog7OV1qRmP
69w5SsVu6bWiltZNg0nJ+to6VrsUxzcnwKPikrFrDDna/zkqTc834hyrJdUqADrM30m6cJyDRExy
JKFw4GPRHLMjhDzHiBhzblifrhdAtfCrtCSinpWAzn5kZ7wLf8wTyOXMDmgsle+7WgzysFR9Nulm
MnzDcgx1YvZdSvkH/kWw6c9hyor4RF6Lf2c+ipvINfmBLJQsXdl7/DOVwGU0EIfZWKdya05+TDma
fOMRZxYPufR8OM1fwhaB+xd+cSHcEesYEaRQcZf/Syvn3pkBH9xzJc+dIeVuplfBJCJ0ffOyzb5Y
IyDNE9cHqoH+rHCoK+Na2wnOXDBowydOl3c4CkeNgc0APwDFd/K2h+5gC0I/sWIGGFtdoiEpC6Au
nb3fY2fYEyT9rR92gPcDug1mgL3sOR+cOuzgVnZyCarzP/EiRUsptWOFZnMoZQEFUYeKYJcjOdmU
OTaNpxP8aE/1VUTNqBINrsxpFPtrKrDZSdmfXaafmzTDX2Q8XtVSmAAw9mov7xRKxrWIOpgonnmc
2vqmnBw58cBx54zTL0gn0GTfu1hIMOXqKIom6GoYrXLmKQP8GNM0ZFHYPODhhbcCLuDPRX/25h5O
nW2/carsiJ+ScBxlPh8IO/d+uiQMJnNRpcgX8Yc72dMKCLKP67OC6U+SsMevJn+ahSkISusnNR+d
qGGeFzF74+8IV0Kbzpp0NHOnICkvAUbUIjTeJj7hD1MDRiqHKRkaR5o15uI/3Tvoovu0nnYVQzqE
hE2vBjwVtEmWkn5m0M6sKXAgOyTz4xyqfMEC1+Px+GUEi31fvtTPDMXZP6VLRnt3Z8Jqa2YWk1xu
K4hm/jW/AqouYONoN7lWYamy1k9Q6u9I4aNqg32kdBcl7aVMYiTEmHlP/Fxhy+MIXROd1GJ/g/Dw
b9b6jA2HhfwwHGPFfXH2QbRouxeT6QVGVVu7rllhgPUXZQuhIbbyHxrowEhzFq15xy4/bJJXfZHr
tRglNfOdYQRvdh5bS6eHs5XxlfOTJkxol9mFo1q5LyAH9t2i8UFM6fzA30jDPnwK11NMPX35P335
ltZGwpDEG7fcgq18bLPKcl8d7MRzja6r2oiSc0+pdCX1BIAfiSL/h2OirDMsReMHTt7idtQRfHY5
Dsnb/qS9a3HhB6w3VN9nd+FsCSIY1/fHolllU6l24JItcwUcX74PRPfrGznFs7gzYMdCTCzsSg4U
JR82EgbsHkO05scEt5eBjV55wrn3N4jZaFWaNPeNtUgd/DOHfvPx+OO5GaVlBdzmuuhG+SepEqd6
TBFXngQ0C4ZZbdVMX9IiyGFQn73yJ/AGmOi5AWYR9mq439IN9h+Vw6FDQXJqJl2cF0glJwPbiCNb
pPogIQDzpixiRXsnY7BDBvsc28FxpLUtK47AOfs1qTKCTbYhXC3AYXNjUIsxCgf61QnYnouBVNjc
kc1FSt6MAf5Fl9o/j5lDJdwevZvquiKVV3airn7jNJyzw3YZBTmhobewQ1MKjQ4C6SeA3aFSA0Kq
jWDmmOOKm7sY1RjS7M3+I2Ns8UVvou/0GMBjRRv+dup6cLkOgiwY7LefbHicG9yuLO9z4cSm/+XO
oaXDKoRx3ZFarpzdBisiDiB/nYlvvDdogzXckjshPbG5l1Fc2GG80Do98SgcjDKlXELN5YgCAklI
vcI13F6XW0L/t5qPVSx5kN4ceUGExSm+7onxOrQuA+YVzu5Acr91CVDBrfxGl+4r0dRmYUeR/WXD
1UH8nvGkmq6rrcaBoBHVXaKhrg1xCNBj3agDNO0Q0X+bFU63vOG9ZdZ/RXHYzGWPV6K/A+lBMSJr
1hzp/8RRr3Okc6Zor4tIEatBlCfi6hAsaJiP8sV5B1jkCuDL+BejUvnRbEi8HKbmKp353pdnME1l
JfjcqCupjJYotYkn6Ut04Z9DQmnwYF0xvnJtSsvKzudJ80a6tMINIdVHMZBO1uPC34vEbBSL14fj
toWcoNR/Uc70igaywqHNtNbv1hBbRLwypx6Mt+h9gvHqzLPpYasbMLkCAdVY2m59tG0kOvNTEQVX
TW0pjJNIzIw1XVsNE6KLltNAQ/oC6QynRpqPaZE3j7fUxD0iWEafmzRdf/UqZpiXlEO8Hrcz8iz3
8HL8eI+6fitHQO88U80WyTUnGgr8y7ZQBS4ZZoi8eVWeNtdam+s/MmUHVmHQkRODJ1S6gB0juNfc
PFKelws5o0mUlnuDW854zUZ5wCppz+1okbpc1RVL9FnMZVqgpp+6JC6oDk0M96Om6XCPnCSK6I5M
Yhz7Pyx52WgEogm/Id8M+AXevOy7MBwI1gAMNMTSQb31CWlv9lBoaGfCW6wPNq+hk82X7a0wwimL
miCwLMDWy8TNVjEp7rvFqjOjgSqxU1s/kLuBe/QYjCqHrQ2ZjZ7Bvh2MUaGFqk85KPYhZxLdY59E
Xq+YG0h6VNsUNYbIQJ493nmVCPjnRMhNR8WfGUgqCCni8g7t2z908sjLhW84Pe2QiQ74FfpF93QX
gGhLXLFdFjmuAKm4quOvVnrb2oV+73xFibverjgiWEfSUwRzqQ+V1ysV016o2xEI4mMqpBaFUrkw
Bu5JijAxJQA80rfsxO5QkYFmYa24eT+iEBxr4wCH1vKloKY5dQX0KQYzhKyIe3BVhIq7ViGpZu83
8IIslZskG3WUTU/jc2+YkSguoBJdqrFhu+m6pBR1N1LLS8wbgE91VxRiKCIic1bR4yz0jonHZvf4
IiUjpfvItGQ/hDTFQxC4gZXtPcW61DHYvr5E8LvqBlIZ8i+/B1VXrklYACDxSSLcqC4DaqC2/82q
nyPSCrao9fgyuG/3Mg7ixxkcaK3Js2nIKgByAkYXr4mdsO6IYZW3+6SWaZQpZ40C8UwddBsk8Tqy
eSqgv02NbhnGElDRkNw5fvXymlyCdFg+54FW4z8aXlqdm1UyCoFgmHKO6vrHA+7M1ix7K7r429hf
xSmBZEWH1HYfswrDOfwCtkfj0fN9evngAzK/FVNM3Ij1N8TMCD8A1EA/S2X9KOTPbPF/JxIyeRjw
KN3tUBFFg6+NTw997RnTKD67gzWnBeM2LPqVzkGNWEDwyV6jdEtSYp1vBCixehfNxmYNKqgR0TTN
/N2vy5vZXGpVVBQN47SYaFD3XnujqBgC6u/OixXmHKA9DHFFGpSjztihYSs1RgtFc1yOx2qK22xI
JTFh16ESavPAe7kceHaQB0Q0hBsV/ePD26dEgaQBQCEi3nl5gFNqAZBKZudlRqp8YzFHLSKrT9dy
vb7C24Nrg2u5aK2AebNnYm5MWy5gW3PJXKhguYurpcok7h0iRNjQdVBtbbQhQimlKEww2hvo4H4X
LYRm9Y0z0oxDeEHqOnnX9LXV11nj7XQguOBbEuNSqcJc2DrmzUvuOmjTGpGFNTb7k8ATkY81K0Yr
wGe9jnG8NevNhOQz40k2ZhJJAvPTtu/RWf0IUbxc5YB3w1HuQe93C8PBkpeWzhwzsXjvklT3gome
5sk5eBye2SlWJEvlDVQvZkSm3O2AlOKOr+GWbyxI3EjLDEH/BLvtSq4Geh5j/FCi0tk9+JDUVxI8
X26oL9ouwOEbtdjC0EGdzQfoCikq14wg1Q0VSFN8ITuAR/cZL7bnVtc9Vmj3KSH8cLWhhZL3n1do
qo+AiPCB8osZgn3xdcifoo9bg5L4/TTe3o/CGE0SnR/u/Pgu4FGPKraqzY6wocT2plv9LBTKGZJs
b7ZqLpHQ8nUD6m+0wxwCtXCCRyWqLRKcilaKNr37j7/HgtN7wttOxTVSsU8Hhnd4XZT+MTFLCeIZ
mydrW+cerkxpSUFvIsS4huYYrDkq4xe0kCDKdlb2BdbuUOgWIYkXKFqJ7cCZc/P8xI1yR23UH3or
t4cpFlcjozX5SFtm3/8Iyd800RYqF88CrerLQAbuhVj+UEP1yjzpddtCO+yttL8QlsuaYusvPUs2
vEWodfFhKmiSpcy7Fj6Ynvf8ty9lubBB+k5qqCsVFMMPkE1MH7wLovO9MOhdyaYcsImDStubKwTn
151lqoY4WkE87YcHWljOA2veHkThr+kY6MzTHusi66xf7V65YYyeyDvtWF4Qx5bcHJ2jEOxbuPmw
pI0C506wl7XgPDoSoT4iIHqRWZ6Gd+XBP8b1cAJQgrDIfFDR6I5XlPmtRkcnXz+CBapl4w4korl/
Qjn0nofBljWsDbT1gqLbzXd+Jxo6iAiw3tjPvTQ5PX7TTFx1ta2pbjVASjQnAvYbAahniEjAD6d9
AgZuylFPOgPBOfsOgjfKetcu4u6DbEavj2Yq0+Ezro+0wNZCUYr4sM3qstBC+o0OC0GeZCdZWcQ5
nfak3jbhzmoVxl839WMA8h1+V6SVaVf6sK3YXMXyZWcGXzRGIMpHsJe3kcFaPY56/0KrJmdx6h+3
rrKnG8itbkUxfLlsLus2zIzKV3/UTvvMFRE4NFNi2OsPPww9Mwx2ZrKu0SYcqK8PwBuRXQxEmxZf
zRJEvDGQrh2GXImncRYbYksnDoE2r4owgUnhVDvSqBRJODT31sgMBcbMh0kygFNjCyycPwsEZb9G
fbu9y6bE0z+fyl4jnwZ1ozqEcLsFoeT9LoPSHzv0qJ/PpeecWlBB8P3TDOuD/kp+gMpulk9Fv4qh
bfSwq2np95gyTLwY5hiV9buLGYArPXkp1tk76fjeo2s3w8S6OU2/Egen5TVNW2GrUEWB8oYCcwwu
v9x++zOqTF7pu1CY9zOAI97vQP0+ZESpdCR3Bq1pUarj+RxI2x50NDwuweYorOmBQrqswZdGBNo6
v62yo5SaWvtFNpkxTpffv0q4V6aBqB+K4Rvv0J0LKqqSQ1qkEoxa/Oh5thC+vRCaUOukML5PP0hF
IcwAXEV3W8ajbD5bnztrA2l5fOa4rbCvXj2mEyz6Z/ohI1ZYMulskmCrIdYDj/j25Fnac+mAWuEm
dODE90jjf0nVXZhBBj1pp7Iw3+bMfn1GLKGAmc8dFfff49fzxwig8E/KG0Vb5O4gaFEYjuZPImTc
hLBDdrHpkD2seJ/lcKLD4QG3cUyO5B0py511l2TwWqQ/d13jY2GFmg9ngrLZIQuuzcHK2pkpMLPa
wJ9eDUFKDAA92tKaKW9sKdPeNIMRtF+pjYk997d7QW4zcz4xXOPh1bRZm9OCEBDHXsr3CikeNOk/
KQCw1sZOZR8/61Q4BbLAl25bQfjgSyGsnqhQPG2LHuWbvXlVEgeGYqB8Wt5wU4TVY+fFFwgF+pU9
5qxhaCzotb1OmSCGci1etQhienAWrUZRE6l8z+E+DZIr0tnjOYWoN6CYFtBa3wsk3HPbnafiOO1v
nEoQdpayb9IQZrtQr/IUeptE2XSgxlH18NDJOpDJpl2WIBbLZeN7USmgaKiHaNBwAyCs1qZgneJc
ibIFzod5nE83Fq/mWl7mLoAukMnLhEekNOWJUElQNxPDxpQ/se1bBs7RJTbNXeQsvmxZpR6qk2rU
wj9WF5jybGRXp+IWjz7TZSVucXJl1mG69qfVAd/8rINzVobitJhD6QO3+CvVJe8pOWrFIMlOZ1xk
C+yG+OayHB6VQaH+cLYVyeMzFJ0DZRxEaPOVPdQ/re7Av19RVb4S9clNMxsa8YKt1eKpgSLToKEt
vhfK4XH71uDEBJe5wz+daMJN/Q29iB2aYnvNQzPetu2Qtbdcbn9JhaG/BTW2t83EJPhfsgcQW8tE
BqxSce2DUrkP+oHaedzzrZCOoxD2A1qkuYnp/8pKbMKZJNNqYBkY/WhDRuRNZ2A24S3UgLhTF0en
XtTDfs+sETKqHp7QSxv4x01iBZHlMok0+hOjr86w1S3wY+d1hehNmUSykyKoWO5y+lAnXfHcG/2W
VG+Inm7eATvfDKn9wwydvmFmHuoMtNg0jlvGRL133GsNXQmpzBd1I9tPe/HNvhXr48WF0dKcIXdg
5/qBbZAVNWjP7BqONPSEsIGepOaf7bPYC0NWgQuajAvdwNg++++Z6HgqbbUDbNy0cOS1SPqXK5nu
juPBWJD8SKMs6wGlBMn508NeAo3g0xp8kVYsleWXRn3G7LUg3MSw18qc2XGgM/RnDPWg7jNg/Pal
KfnEVc7SFpZjm97oLLG2hWz9aQkhicfSgLYWr7YO+lOVG69N+tI1nwF2P30RCNaX2lsOp+8yZyfU
p9K9t76vEEHt4rwQclWLsCx1wv6vOfdPbLvHEYoVfDIX2Nzem60lbhaxrY2m+0eplZGY+hsUTJhT
E0f0g2P12YuS+DXLJGRHLLqtMVkboOHltHcnTWiV5nmzq3UJT2XW+KeDXw/DGRB8JnHPWZbFziVa
NGcHolZeoTGhToFv4t4KIj70s3QHQAsEHXUNbtjbA4h7ioaHa/ETaHYcyJK+ldmAUOcIErvkTYbH
/iFO6sE5qXsbAhfivYkO13M44D8LE71m9/3ZuIm9mSloFxUyJAHVVf8RfJDhfA4d9D4aQNKhJFeh
NM07amxLOvPR1zeidrH4eUX44kNenrkD0dHUHShwHv8y9MG/TvStMSxvqHq96YR+ODbc8ejJ6uP8
U6hkLDAz3W+S9ccDD2DjrgQoa26fZYlz39EAJZPsbZpTc4NvJ+FGDhWC+MTP72MZO6e3CGSwhLMo
vU+L9mVkNqOwlOdse8mAfp36kNkw+ZlFLSsiay4wYfdh/itzOQhf+rPmsqHJmuP8KLmW1wmmkYrV
5jBNHrLUbeAv1cYPuFSuIgkf8kAfYMAw047dauIPPsS2KtLCQqIfboc770Q4ijM+V2L2Q/0EYum9
kMrgA+oyRwd6xUHeDa7m/rFVPe0n8cfETZm24ghdX2VYN9PwfJF18wBsZIG1PzU/O4CG1hl+W1UA
qNMi9xX3OvOKWLnsfm3s81FG0rsf//GbRNNIXJZeaNFQ0ERqPIXzOSqI6u8X/v3Y4aT5V9s5xBag
yrPnwyiLVGr0DeKfNwwNGKQl5IvarKN7qFK4mzimANbXieVjTc2KCYZwohlqFqQsqawDlZkkEWE5
pwSB9jfTX/2FqVA2HgDWDCnORh5E/bCQfcaMuZSXykqwTZDayPl/QMYHh7jpthHU45hk7Gr5Oj7a
9tCe3lWmqZUF0mohQvosabvrlqUdGPYfw0AT4RqV2Y2bm6BNtx9sFDM0d9C4RRf4AR/5zWobhyib
p5d7KDe494ZUsjukN4WkE5foJkErBl6tjjuaYOwNF+9/LkvueFhSYXzYc84/CWOhrdCyV8etJqje
MAGEDgAeP05/Sq0A/OxGTOEJlqKj0QkbjQGX4sg1qzK1sR6ZYURTXQyUkkj1232g2OeFLqFweAkP
0E96FhdaQ8DgrcehViyrGUJ3wFPOAZBVgwQpc6TJ7N4mtSzbXcSs9jgLk8rmho9r9x6Qc/zIZ0J5
qAMEXJfQKk1onOyqoW7EcMdN/bNYOI/WPgizxPYrv0ArZwFQXAydU7EtV8b1oXR+PZdgJmbsGm4s
V0ogAjZYtTlq9ShXqiVpILlTphRUYLGos05djs6YuEUAbo1HWnfq9Ovw4nKXvLmCQgSMQiMQ2WSF
Fggl6uworlYg8sQTdgmUZ95mBEc1+0RuuGfffzlYmUbpWNa+4w73hDr4aOSZILIAx4n23G13XE11
dU6kLXOyB5dP8jDRTSP1xRbDc8mdIXx8huB8wjSP4ryiGb8W2S912UJYr3KMLwTY3Z+K39zo81Db
NBbJ0sizGN6i/eOmwxI7RnNlsCfop+CVeJoyzNrsEnYGQWUdQw6NjCCtYq7zgZNhZ+OxkSR0BcL/
Kp2G36BxA9lOwurSGzI4qfZAdBykaSaE2Tpcy6jjMZXYE6LPE67sIelXYFiPDtVJg7eR329kYvRx
LlkaD7Ll+yEUVpcH1V8MYkR8xgjQjG7ksyrxmtfL+zAfFC4KQZBOAsYpd5Tms+CLQSYYrm2i9ACg
kAX0Ouc7chX7m9543Nc3dQJOQs0ZBhzWUa2oObmPMuuqNaxNLFPGQvTKHiP8soEuIqiUFzw6GsZ9
vF3SwJ5iuCp8O2VOpE5b3ifBsF0GvwNeYuLL6a5hyGSmyYM1tMKst5aYWbDHsFT6E50xQS+j60ao
IwdT6j17Qju6z5RSafI9FgwjyTexHvZurTevdYpGphHxI0pj10nb+gk6u5fAij2tvsN/Oq9K6WOc
vQ4HPEuXG5Db3dY3jtES4QYND8nX61nhMRV0+8G+JjfEQJgm0mFjfxZE3fr79jq1PHA47VIHDfGS
DFXqkbzcWi5ft6Q1dgn4mT7GF08mG8ryjXYZ2p68GJrDcmix8OAA/URglmbwHWcRCyoqmgYFg8Vo
64wrvz4ow68QukBOjsV50JV/Vovv2szcHB2sP46p92dt1Zlw2eI9x0MUVHofZ14FLF8zxN9wTggj
3Jdf4QhxrQCSmjTGlT56Hkt7c4YaCcHTWCu5cJfJIZsEGrVEq5OsK1za8NdtvMRrDC4CXtEnZKhm
gh6yDaUnZHZh+RmhJJEVkLC98eXSaffi64dZI0I2wsLrTRW3VnBlb1T1soEVwnmxEgF4tuKP2o9L
4rv0Ed3ru2u8KoD4X7DnNUhaZlB0VzC+eh2LrMekr32Keq/NW4HN6E4pmHPakgsSo8J6b7jzSy0l
ChKCsNzaO3DzydBUgTot5w2QB/a3UdiaPONBVUNqQnrPMTmAMvjxypKD3m0AnsPPWNqZtK4MpwUe
CjcOfld7jYnA05vlhvo85JcI+/wrWUo5CeSKFl0IaEje0Pn+XqK+CRwQysWk7W0a97z6g61jCGYW
YiOkv01X9lnlTwJsqhewD3u/Qd7D26bfDa0JfNr4e2gszG+5LYRFOuaEZ7VB4FNVw8HVeLOerL9j
Z7sCTMOz+T5Hpz8m1ocreH5VRHa452JC08s+YrFpocctEBuYxYXwdPsiSCFTUl56f2V/UDVx0jdP
5oT5NNCvBd0bJDyFxocvoJEMWndVWzlkA8RtaxshLC3wL59HAQ5Z2uaqhLcaXyr7tktNnNQrsajX
bgkRYuC5iUIPDL8ooFILnZchi+TyqQmybgJrcZgXUvtUeaGtxvHFUCJaSdWFpduJ+anjVbrD4bwq
PZXqCghJXzXoIQk+EKupathTm9NgjABGE9QQaQWQTmBPwBlUGpfONlp8YKrQBogwYfJD3TeN4xCy
CbyfqF17bPE4w18ei9vZ+SxTxLk890hwMOJknhIVUcmXk1RnKtQS/FKXF9JXb/R9VgvI2cKrFiTO
6qgBvh7TE0jUGj+MkwRL09bFq+SCgPwcJnifXblpP1qBl1cbfB2fyTPsrFrnSnxNBibNgE3E9VxC
2ESIDMg2Dpg31Oza8SssnU3Nqsw4tokkZ3U1Wc5STyXLm9RDJe4xC2ZkdWhOe/PqXz+J8kW01iCD
d2RUksOG9OnNMfXkHxsNDJBcn9Ww3s2IhAEqD+nZVirAOsBqgxT7fFqdJPpDwoYUfu8ETsdHrVkB
sH2u+eiWtii90r6s0IG6ZM14qJuJ4xBNClR+9axIRxWrcPXUPeF1ehTHUV9QqhUPxx+qnTYf2CVp
kxJzPahxeEAduiDoKTBtUgdxpUty/6lPVMnzezU5+gG3MeKhVQ9+0jyWBjHXs+UIVAj3dB2omQGm
bvwUFehFWeK9oElAwiMYH+qoU6mpcFUAfIX4QOvVo/D9pNbr4Jhwn8zM6J9WhSdnk9KVPCQ5pwIU
NV2/lr1VtEUB8WoTKS9ynsP0hBEECREXrydymYmSqSf81DBj64erDfDRqkQADv+BKMRU8TzSGRWS
3f9vSd99KbWGeHv5Vx38nzBA+mNVpOFZEyGihXQomMZ3quDcrLn1h0bP5IZYM4EPLmIiC5gfSmtU
c9IMuxfyyNqeMj7CJedlPFyko7ZoE2I7wtg9DybH5gx6Im2j+GLG54Oyf1DFvF4ui6sfF9iV7oPU
2GI/laxjByiAcTjV1EFNjlIe4ZaOG0hjXP/nt7d45//Ig5FKFI5AA0PmkRrPcDjY469WyqMeaz6l
AJuKkxELOl2Bv+ZNDdKnvh8oanUQWc9m/Wv8zBOdz1j7aD0TjGP+dHJU0Iycof0Vpe6h1TPL9DgB
Ftd0QNBY9Ba0J33tuv9bmxOg+ZqiivLI7IKbDgkjBwNrzMp3rtiWgCFmf28FMflVJ/+5QZK3GjFA
35/E5/QBBHbfUL1ByQaVwx3x3I7RtEOgdqPFEXaauvgd0E5yB3gS6czP+wTXT+oG+h2qD7rtcV9o
Yn/o4ekYEErRT6nTKLPgqXeO8BTmCelVfHfV9u5Tdl9yLC1k6qycSMhmWWlj5YgHsxhP5gDMwBhd
V6Qv9QkHq1zo1wrtEog36CjYQm78XtASPAQh10ielxENNxDwy50hPAPCH/dgTte8ePVc5OXVWngO
on6WZVQ0WRPE5ufLu2cZwADJ45h9ueXvTF105heG5cuKEoDofXOUrHoOeHJB5UQoO6wgL21ZEimd
8EiouGr6bo4VzC6TphLoUMUhobCOnX945aOwo21QlZPFo4ODVGjpMQaaw00bXMCANCjrIiqahYFQ
KI2u9MM6tnz3v9nYAGKKzW1f3Hsy4tb+9nARPD7d+tXNu365v65RA9Wh4XwPhrQM3Eavhx1KEnrA
2fDhq4MRPpfRLk3HKq8Sk/ZnB/v5HdYpqNLZ4gWskwNAUmMLo8h0lgIySmKLGbPjnqfYLfLjCoF3
OD4/I1L3dT6hUqbK9t4pyhbf7pJguTw78xGbryLafP3nsfl4ttnZNkUa7Y9gWMAtx8qxW5MKQhTw
UAqJ4ckG+j7R1jHYHbChmUhaFEIr/5H98DIroosY4kffjBnTw9lCpHmIxst0ATW0T4lsT8Q9T60F
bh59UlKNcnQn2YZxPslthuENiLPWlv2K2qMChFgOgz/n5M4Z7M38LqMxbnPvqrVSlKCv5S3+ZF6p
Qrx2E9XXkec4kB6xqOV5RERVNYQ/6cGmQ47GvPkNakxUP2F/nJhzNofbQpaGTgJ/GSMsZgk9wC6O
EOgrI7wTMq9tPPy/l/qbIGVdfLlOYh10b3eH++NeumeyhWfqDJewGpV9a5d0CL9QsUnsPAs8p4Ez
EckGKoMU8h/LPW3xep929UiK0TkJcBo8taFgB7oB1T//3aXCkAXXeCMSO9UU/GFvAJmF4BVQQNqu
kXJ2Aqwj8SeP6NBy/dtjlGM68HVX2w11dmOykU1YKO8z9nbcDs5ND6IqSu7vI0A1o9U+W5MLiQD0
0p8KcG3Mu4AOqb/KD6riPn+h6TpMrrxdD0cfWc5QXvP81kULdkiUsTfiM0lnSmSfAsIKDL0MDfuZ
61yWnSQPbFSGYbtZ9xO5u1yrA2NnZzFTNMSbleH4OcoJh2aD9s5bZE9iNcJ7ZvzV9KvfgNcE3ORq
jdlcnOro0QzoOF9MMcqeSdO/v9Q4AqtOTZ8Kdr/8UmuT0kdM1WCsWitm3NC5NnAivtiGPAoWFRQE
r5SM+gQf4lbiMMt295BX4fPxFm22Y5g1+bqEwGCFfNHcHKH4NWlP3g5tGLke4/FGlu9C2NjLJSyY
R/AP4abm8MdpZ7u4NtCyJIQpX9RFFQT3vMNXaVpgNSSsKN6plBwJO6CKf42BjqgsUaAjzHeOZS9M
sm/et3Drgh+B0Ck5Yq3Xe39MJSxDC+k4ZmbU9/GWnJodbsaqv30MN3ycDybYmZKGBVKwHf+bLBy3
d8YRbI0NH8bFvjkCmEKUXy1HOfIqWyo3NSG0Rq6csNocVYnR3Evlz6BlRKTDROPVUdwXB/AlSI4i
gPC+5BXS0cvYRFBgSEORpdgJaJG8tHHlzaMgiFHcFT8MmUIH1j+BF6+AGZAFA0U0UMhXRW6WEJW7
VqHHcvpciv5zbB26Oy1CN0vmPSFnSgLthI4Li3XHQ2ZlI9aUMKe2NTAyXHzCssQ4HUyDOlX3WNCT
DKWVIlHw9ijFWvVjzjRT3zUEMmTYh2K6FJrLqT8fnFNp/BRlqTL9sGolOCMzmgKC//PdYT5DoBXH
N7TiOsSA/kvnhsxaJJoc7r2tmqjibcCLxdUL9/CLykiq7UlHwGgwggEfXjU7FP/F6k3rEgpRf52W
Ban9i0jzibkfv9cLPLbabffmDqeE4Mc8XasD9q8O6ES2hzs9AJpw+B04VRyizKfMVOvoWx+SiECn
PNFml6KlFRIgBDtPFLx6IZvttwArc0WSawsygFl849s+GJl9k6g4HWTuHGWYugmVvqDq2i0xfJQ2
i03jn9ZbgZ9H6YO4sTdUG6aMIH54kxLUqOsPKIRV6Q5rCllLVBy0iRoTwnYpN9Nw2L7/w6YmWIXQ
9wQ2RjpBA0exz9i+Fr+NBC1cTlPl9QxVKfM1KPBKgCl20Wq2KTxg2EY5/V8czN0anQYWnsoW87Hw
lr4wykli+1w89q2kh/EKkdhrjndmTEa8aDW3SvohpR6kK5U0pgxzrYMgkTADQrLvipiTJs6iDulr
qhMAQ52Rth6Av9qpUu2n1eNQ9XeQj9jk+RheAB8is+KhrtOpcTbMhZgQPSSQ3JmngvB58nF5lvC3
31JdMImjMtcg1Fi/m/MNGpx2EmpAu+Wh59InIrkwRccUc466JBEVaXvRm5wI1ME6iegjEC2e2GWm
iCr1Rin112Xn98hTStrUiQWr54SP8ktKOsiEbFhC6AaC2w7hMsSsPaP0DP0fgpKyL6OsAnjS/fAC
66AfoTLBOXAP2RSvso/lHCNeEuAL0nfbQk6bxk8nGBY3LNpvLHyF6c0+dp14k14GAqqtC2fIaURP
OLuUjTFlg7Wq5nxAASKZ78wJ5ZNjPj7V6kxlBQf1mxRoJDuBTnNzpar1eIucSM6M4OmfovLw9xQx
20rvBSg+xqqqYdsHN3kZJNCv/mq8SO4S7WD7NM7VnNjxfCUxqOHbjdbvBKZY6aAbxpKmdxZLiuFx
K850qI++yZCu8oPKZzGyYkxxWIgGK5HLu9FBLk9haaP2s80jVxsOHGwICpHI6nZ7MU8W2pQO4DbC
D1rITtBsvKPYeDQeX5tE/HhznIDsW05866mWTp3XqMKVKS4ehQVv1P0e4qD7JnIbpkPLyh+0husd
bQNnDhF40lGy3RQzHzkm9CpWwbgqwrbD31WAtTsBR9k4tcnOTUj3T12mnvfGIJvUCYYSQJiP0XdJ
pyH7surlBiDMxv+odGboiqb8wwNIQ4S0qr//FXj4YwoRx7xA7HGqtU5K1MO1Do+nxwN6xvlzcnXw
Fwn4KCqBBfXpDX3PsyCMKpqRUjA0ka7mRE1TxF+FhbBKSMJ7EXJq8vaOMhOA/uc1Rv/jvktWtSPh
vUrhNJ737MHtmBmgxNoD08QgEE8rTIsyYicGDW6VpZvQlwueH3xryOrc4gJbdQBJX3rWCD+KN2mV
h/nFFqzqdBrS+VS0oopCErOsI8kqC9J50YM7/Mkoljl9r88s6d3zn2uPYuejf+HKNMLL3qMEs9oc
sjxSPFDmL5Cc0vDFh5fiUqtvIigd8BOQedzGg0nUfy+SrBQ6hyhiGbPk7tbA8VC7Edn+Qmj1oyMw
pPZLyGvs2bUbfyVRCXl6FRGKqz5pqJ7O/jY8k4Z8GX7ByZGc3QeZR7Wu/OJrhWef1R6ROWs8a6Kf
okSS9J8UijmH5Ej06MgJ/P6Map3Qo4WZVvLza8HUlYFA/tBg9unDG7RF5APf5VFiZoJ9//yeVIzb
oBir0pZKkqLePSP9Zz1s0yQM6Ne6RI1qHzHcz+9q5QzWqoGNcdnFmOrpchtyCLkM4qtHSkoYSnsy
yv6I34tnoyZg5X66KbYjnuCnqfGOHC6gRZyfWNbKvgydsPyBcGXtVPV5aHAYwPpqE04ZidW0h0yK
ByXyt+xnemH+bvT37E1gLJ7RnWzylpH9MXBGSYtFoy4KFYXFjw/Q8WX9xbv7IyJhO+5oEZFiCftX
OQcjEi0LnVDBeQN7sLyPMCayr1fKewf5FuEt7SONHgmgQ+Uv5c9mF3Aj7rvTs0rPq1WCif5JeAbw
0YPBhkWelzOIh31u3KTUl4WHwHlcHbFICh+3Lyd2tud6YLN5T51AlgLXDPiTF/k3x4glpRahsDGS
eUbjyFODGzOQ81wSoANpaXNCQnvLQlUpJgAPHGwAjN1iFZGv+aF+OyhzDtdtiQnXxBiGCKhjQSRG
mSLAEC+8QX97jyz3hKXU+ndiEXhzjjrNReTKdLFMBKwYHal4V6PQAAGGuDMqbblIZOtl3Vdz7Rsn
UcFsdcDB2b5RowQ+Gaf484wPqyd8kgGVY3rz11iftfEQw/Gtf+DIY/yMXjBEZm4b781ptdkIIpj8
OgNcoMfmDJ0hSdSDmKaHB5t+Sh46kTE0A+G9uX4m4O0ttLR5CnReEhtQCl7jzLcQYs+CHS1UQVOE
nQcWGsP79YBrrIGLH8pXSba0y4u9qTYdhsWdb8m6Py9g4LLkqEAlO7E+jEJ3RQ+hqoJdU6xrwuYB
kxKEE9qNZvfhb7FZUN8VzwGENO2MpnMl+lZWVzflWKga2Z7QSuHGwGpwZTPx1yJ7KWEFhrXxATBT
BnOAx428qDyy8W3KFbroChyqQLXvCy1QBmZWVlrkDTYekj86DRdV6j1jy3uTWwHVbwSXJtpXVw8x
B6YLa7c4YlF8NJcWa2ULGKblVgwNnVkxsczfZ8OviVQRT0tJK+gTsOfvtfxZQusmrV8qH4pA22Lq
yhXbzN72skzDR4hf2U290+uYLmhNGBI70XIziPm0tIkAJNiLhR1pI2L1HDYTV7biZF3BZlPFxJia
GjGb3ZjaQEJ68LI3h9KpJ4pXB246cqOYuRSaytGWJz4dsN+hT7hyQK5g+U9I/V4rsNTQoF5Z8qQS
Nx/45RoDjNpXsVRPkTrONK0e5XrDnlQfEaY4stMM7zF/w1NBOqMK/w1W4mgtNeb3qXB5gcDiOk4b
v6eH22GHHx22lodBMxQFbdqOQBib6tW2EgaW0DvLI8o6knpS4OdzD+VcF0OEIyVVzNpCB1ttAQiM
7tg=
`protect end_protected

