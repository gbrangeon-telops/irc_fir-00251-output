

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OHeaBmhw2WWXga/8pOVTMIzcYutI6Mhna2kzvZmeKvttg8GRcsMBDXpogvkdmdxp1KLLzWXMAKSV
fUAOBPVAvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ao3tKAmGrk9jDIJ5tmEl5p3MIRphIc7Vg/SqO4TER/rFDRMS3J83CwQ2b9YFrnde65FSvizCvsTV
0Knxkw8zoIma+TSgIxOnivhI3WBhgKeA2uGkUI4h7aI3JKyXt+ar8rATgfMIjtkwwZmXnAQdFAm/
DhnKD9KmESp1ihQZWxM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tIRCJBwrqw861TllYkYZisN+3Hf+P2JXRGH4rS3/mIyKaeRa8ciKvXh+DuDwE0CQ8FK1JKt0o7Wy
5niCab0pNdgMIWoeJTN4M3Yv3mIYHhxe/uhUY+qL9dbTdi1peu0ypGwB+pCVAaCMnYsMP87ovoxG
mFxz/aWHoq6z5hUiOqs/8QctFGTu5uGrqo/fDpwnQByfUDzc5kOGUXom+7Ix+u0CBnUzxUPMVE8H
FW15FWlEhZ2/WOv5odw8POvTaQir1St/I4TCBaM8Ne779Z1F4E4v1nyrImWHcYGt30Ex/kdASWup
x0rIb4g/F4zfpMwk2F9PI0IRzfsxsXBx1PSZmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vDR9iZfmcKoc03DxzsUkjAUcoXZpLGp+jz9oB+bhIzk9fA1B+YkBJ4B6wGhxOSVsIGzj0A/2+sve
cYv4/y/PnMWoVJu5GAXMXsNWS0+yhRlFm65eqZTnif9T4BQLUfDB3Poe8t8+8qJraoiNha1dShh9
FtnafnjfaWlgFCK4DSo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5OVsGiC3k02pbA8zjICborh5BXFBySD3cMhIIsNr8DZdx+UrjbiVbqZMU9Ry3hJ/1iX0Q8zDyFo
F6W3nmvV82n8xeQJN36fxUpz69izOLDYVC7B/XqC5I6fwrewIKThxTuK9lZtFdQHHrzj3T2ZDLDy
Z1+PK2wQ4cNjjft1DSS07aO+6gcWXb8X25cWmNGk/P6Hl0pzIcfFFHwO6Oq+bJ671kKmsX3jUKAg
DTTCgxx1Ex2XG0j8cWCnhZjmetyd9o4fKBdb10goxmIXB8/8Sn+4BcUJVLUQkMnRwy0YJGGtpiHs
ZxxUU5IU2sy5csUBb6rGbP4ap8jLGVFhtMQgiA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16944)
`protect data_block
xnBzX5JW/QdFBnU/72PLxH0SrVjQqnm7QnR05nNkgN9Yuh1y9NI37lnkIcSFre3ENMOcnbyazmzT
xnMtwPedZ53Y5qNZxdMJ4jhKheVAwnyMMuDbNqY09cxZblJDRBa12RoGaIoZkHCBqF8nrHvsTiHx
Z0ephFuBogCOQvir1OAjnHfiJVzceZUz1wBSWXvMhU1l+u/MetblR2WqITGF+ufGMaYWTqZIGmyv
ZKDb3Tk/TSPzt3lJidw3wmzsz4pwvmzAywhdLbVSexuJrRqJnKYlNvRByIlZ6tWJMExKGM9NgAG4
4LOmvX2u2CBH7fd7iw+Cun6d0jk0EuSENMz1tud8U/l+hMwFltV0e+ZYhtDWnSB8JbWXi3tGyfnL
CaZRFZueuI1x+DXphvAYwoilQ2SF7cEszRCSY9c97GmmNBEkGMaZQIpMIZYNXblVq2KC77AA+Bjg
kgk0lbsAK7Ej2sS+l4P6/BA7iOsMmjLB1bT+c6ciAYwB+7PKFhbQU3yxNvdsyDH8Fj+ONZa0dDNa
ZbX70QO0Z9/63Et04qJU6Q6yIEavcsDWa6CuZReP/8QWkKNGI+UmPmGeBgnzS0TX1tGf8e2tiPHO
u1/Orn29vSASYzJnJ4zPPlyy54+QAZJJip1kmYOqGsitctvT9E5NKJPSMookr+HXkZdH7T/Tx/l4
X/GHxx7yUS6qlkM2jRAkEfOkgbYlz4c4Aqhf4wl+V18nOk/BuuRvNVBR9sZWdVjRh30CekTQ+YXA
DdrPAfzs33lB5f1KIbHLN6MbbHEeOWNmuRWrLSIxXFNZCfcliPiBg9N755e7muo78UVU0U3Jlsmv
dfvK74BWs7kWJcjm4Fg+NkqGG3AFRRtWXD1NUUEfFTupO0sFa/0juz4T5lxiSYeWVsd/mc2AogZI
I4upS+D1OSRSJBbyA1r5s9znWuMMRz5oL5uQuSK43Wdk2ggn23JVQuKwwv1QYZZfKE+KVE8SRSCw
GaVGO0YsWiMY3BrF6Ca7lWQJYEG0FLs8O0jCp5/UB4R6NVx5PTcaSOyiwB5k1oFi4Sti914FOYZQ
pno87Xl6O1Z4sKsi+UGfs6RfEdyQ5WkUE0JDHop//Mj+7HwjvGWA9CoPX9dBXxFYCNFhfDsLz/+/
3ZWRceES6QpIkWVMkBskHLJHLMVsDPMr0b7sPB7BqpNt0cgVE/xi4ZJ9UkIA+Ktd/KWi5j/8GDnI
JZyHW232+/lIygYrNR2NDC41QolmGgG8P2Q98/dVyCUvVuf6ELNKakvgloISqj4qXphuASVTzhRK
znKuxta+daO8KS8iwezD3NyrPyPI4Si4xNhkexGq87Ph1OV06dVTQCfeoD9co054F845VhW5v0+9
vLpNvnaoswkcX5t59cHsCB2unNm1K1N2jWAdawazsGFxW2pTLXok46DGjQl/Xf6jlbwBpwI59/iA
8lnLYxi8XRQsHzeeAnO9aFKsYowNmTKRqm9whpbSWohNqXWXI+zwW9HuJyIFSCQ9koGp0Uda3RQb
LIJyA1J3oRGQr3YrDqNJnz5+SX0bgEKoXRV/xBYzCYzUxN6xmD8ATNdZ+nCDfqil6+lQqRB0Q+1t
uLGOVNOrrUyZVT6udPBetp6rbWTA2d6WdWDltABSGMjCuxvg/tyTmJcfXI/1FxZol5/BcXDWrRUx
bS4+KtLTPypIVQmo9KxFGbD36FH1XmabF9FqenqUCpH/ZwuH7MeVZHLcoyzxWbqG/C86wYGB1ieW
L3jyTGE+LJ2KUAV1SISeKKFqYyFH4sS7satTVco3d7VQljeEDy/Vgkm8PZI5OzyYIxB/YVFXGIN4
bTnZnGj2pWflDWkM92j0+joGk06w0u+0as09O4KkyUWtYPdocdz2thwmbYKvxCbsdGh/ruuJl+3B
+UbzTtNt8hA0TgYlMznkbwJD0TxFbvIsIYeJ2uT28rMfjcIM22nByvaTPL5EZzlTJuxnlMUDwXF7
mVlfzFM5TLvrxubMu3Hjzkhks6zzE6sFKMi8Lj86JM9g/lyR0AsDcKa64uzbOTIfI8hYJhCLOMhm
I60uh7k0FyG2lmzH5ZLc1A/dKkcg4x/SFwXgn48lIlEQP2IUfLaIQCekjt5BnhWlt2KqdZnCX1UT
cHOg5B2VjmwnB7e5B7/0sLhSxOLKOupdErWcNk2b0z2CvoIKHRY5zYxvojLhtVdYPJzeQh+gYsFZ
20gVQjWlkp1zbVtJiu+2eMePIi9QJbWKj3rVDCRUU87VHq7nwmsnlJwNiyQVRVcEtEWJr21JdStA
kCpcXb5I2GXL4P+la8gaKNM2UILTrCXR9mVRO5jRmZ005As/Oi9UwBHEn9EkORllB+nPVKamaJi3
TWroQDuHFOBx2uUxz10lZim9DRyDklwCqWsBh9voclhdthxiRY49mmsbRD7XP7UlHf0sHzz0P4Pd
2o/+Wiur8byUCbYxfr270lh8yEyD4sm1+Kg0xaMF6PWmggeBMVsHgXz12gRhdxtJ6u137A7B5R9s
05cZgNTOfz0dgnDLQyGFwQhVKRlHZKaqD3DZ9ij13raFjfAE8yOJ9MNnEeqRiYHB793jGTeGIVcl
85z1aoC9aoauc6LRzqdB9KINE0NXKZLV6CIB1iG9xTUNM9lBaYuMUAwiEw/9ixg8PREfchXSrMB0
PRnx4sHYy9T8ucYsaXXLQmXoZRpzNmlAPoEMqMUTLgCcAj/V4YawVOGAnwLzxy+zMjzBwEbPoyH7
xspWanGA4LP9LJIsd0s/wBtgW+6BUuJrUwVZEJBB2wmX8DhnUV8hrHG4tX9V7RVFpuyRcG+izTbt
hv9aoKX9ZtTAvx8q2/ySN7x6/Yc95pydNWpFeI88YQBZpnC4a0qqkonzU+++ayyLtZNYY5K9Pb/Y
uqYi8Iyj/NKIc84H9cVOAgo2DZmj+HCNDImDeoPBeace2jo7QhpWY06xTXOBeL5gacNmz+i2+5DE
JhbLsuREK9xb2x4QoL3BShVbWWHOWZ4G+X1yNZ0h4VIzCwsKuXFZjC8TCWC6ZrPawAua6m1oDBHc
nugyL9J4s8Dwt6MW09PksZf9uK7G4cylKLPMaEQYcUv/Q6RX5MdUxdn7C6u48WEff22Qi7fmKoEl
ImBzTYcc4CopIg4b5aZIjXQ0W1KfQmkB13gdVrPuCntlagJuVTSDIr57C6iMX74WiWAfPNC+H4FW
8GiUPiHdVKitrNAnUHRoZBr2heGGU0eX5OvR39qCbPBW7OGXOHu/SSdP/gOlZTHewcIfkxtYO/iH
VC04iNPmUgl8K+AT4+I8RaLMq3W8GLA66zo7IEbCqL6c7YnSS8PpW2p09drLL03rHHnYcker6loS
tqUpyJAeNce4vPwvAlxSV8a0eYugN84xAn0fNnreDiKYWQRzMEJbNYlWgJqQMb3xYv9hAYvmLQHP
sf/+W2Z9mxFIp9PyS3ywi6HItV1liDItkI+BbtyIvvWoweuigxbYFk8E/b/MelQmFuQ6AL/sKfYe
EgbGTOLSlF+vOCnN/x9D/gP7FP4niqKqcifNybaF33ffEsZf9C44WKGdml6iuweL2JEK3cuA3WRM
Y9ZATn6cvczfd+l7pu4gO0rH1OFAZzvbGWVB9G21frgZsgrRs8jX44bj/QqO9+1Ytm0Npqigwsxz
P6qAizXKUhcI98ZDY1Hy30Id4uIjyv99YD6ywOrphC/xSevaIb7VY2cUJldhoxXP5X5nCGq9o+q6
VuzJptkgG/rkesFBYyJRkVxU5GWDVMVaqnjb23EOv+Dz8/eSZnQkjumKHhWjMU3YIesWtYL9TARg
eaEqrzCD7QBFiqXEeWmP2tvn51QqZoN5csZVgmC9aWcFl5+9UPWvRrcBOLgy2tt3YzLTbcMQxVYs
/fJxOTl5R7hgWGVtCceKQjdxKt838wHJgzZv+4mIo8kMkSzdsQSiCC7rZMGu30Dx9VosqF1hQMA8
ErX4fIBzrqpxX2yyB6kDHYfyBOjf/soBxkANgXvgqrLn5px3GGTytddB9GPB6suLcuGZBW5bUdVB
0M5fd/Ggel+3jQYNTHbqYlVDQv3eFekSXpWzVYR6F7WkZzMCGSC0kLVhZPsV1438vQnq7VkEqoER
vNQcxBbQ8IHnj6COsfUq+TT1gIH8//tDOWjz+TSTURxqZ0rVJ1LiblUykvHVxyn3SDnAWjGeLBOG
Wi7ldrmF7vAIkfSSnI6KFiS0ACyebOGc35Y/Iu+43Uzi41M6oNr+Icwy2rn6nHp3Y9x1L4qSFRo/
A0gOlfddkPcmfDRy9IkVhPuSAO5DnRpUS7YV8liZOKXlzz8Tu+uM5KBEyeqL54JG43vR6nf3AT3U
gplKJlQ98xrmGleu3uXCkhYwehjY6GWYi4u5Z1iX2NZ1058L7+g8GO5CbkwukSXFHY40gWQcZMaY
1S1kjCZVwWV2RKHDhEg6Y1ahqkeU23ugp0Www649O5nyOTnEU+//jbUI3KATtSaWa9b5v64tG4/k
DsyTf7vhXlon/FqvzyR/AIMN6E8uZbTfH3B4N9ndW3/notXXjKPv8NZmL/ZlZrNuz5+l4A/oIZfe
3Ab/fbIwwflqtdSnqJaEvOttChuYay7iWdaRnlQg2EakKt7Wus+6WTWWJwcB7yNJGwyAyLdZhn35
XAWxAf/oGiPFZMEJXCZp1Im2jPJ9IgWcmB7hk8WXM/2/nyEF3SpmTxaMgzGm37htFabfsUgAVgS+
zUFkDFoRfPWMS7IdqPhhyvNUsSmEmhZ58CkbIoNlIhpW/fExn1x329xEQ22YfPieiFeEYXbwAwAJ
2kIHf/4jqTOct4rPAVqfBsnKZQolgOcvJb6R1CXWtXToavXHVfcjbxvCQM65qXfinojzKsPA7qv3
nThZeKaIXZPWu13Gf8yspOee73jZuTBHbYjU1eOAD48GgRLd9cVfVbGSQZ64vtO0r0/1+sT9dIrF
84V2WygLfLLeSN6EDbJB/L6wUeW/7812XjdRjkYK/utCtz+S7JxPh9i7R5Z3+kVY8uK6lbIqrwbq
rUcs1QAYTO2BRBKRwS3YhqC1trYaQvS34urHKffD94H2qKkyi+imzm1MrVOGZCeSYin6x79zkTNZ
1Hy68DATgUR1DE54fT8Bj13mcRgfj0lg1OekcAOkwwImaoj7aKe3eoGEVS/ahOpkCoqtNgwcqYGa
2vW9XEj42DPUmS27uvwgq14/wePXX4sVRz82YlfAai2pTpzGguefOtOSL/fWdintLFFXzmkezjKx
/3RLgIJbRLRRHSPaaH5/fr6um2KdCFeaqDUs313jHHiSICq8rYyr1//M1bW4ctonTH1Tz6QB+Beg
MuuPMa9jKLaXGmLxjDa+fJ5sBR5t5vq3Al2MqvHwWwj2NxyWWGAmVFAlQkQSkFpjwYpg8vl7Nlls
jJFRuAHMXixsNwoPbV6eA7+ttDoNwaPh06G2d56iM3VFix9iJKj9jU5jFSxbZQMoIrGveuYr1YXn
6Yb1Bws/M2XyCzTQwPvfBMOr+w7lPC5aOmjR1KedvgyYtloYFO4Exh9aRZLKO1pjzIZRc6UED78l
UW6kGfdUjWQIP42gxctxQMJmKLofDfOOkIEp4ljc0CElZ9xHeb+zFNKOiGTCMrY4AAz3fcNvmRw0
nxdsYdszMXEMn1Skq7zyfSMMEBSz1daDb1aTRB7XcAtbhotauytitRIB66tdGpTga2EcxiF3hnY8
ob+Qo1wpitlGYzlcs1SyKagUz8UXBzpywgn/7KsZmtRfP/ozCCtjz3xvJzZgmTgJShM+g/G52Awy
0PxaAStsw5kGl+gvP1cQIBamMAtgt4n9hSyukuUSV1eC7LAaC0+kctm8X1mZfEkwmdeFV96XNsbe
bc0u/wrX6Hb8Av4m4tA114NPbkcnD7Vk0w7yx/GYITXEXrwpQk7Rja19voydKJJHGvnYH53i4k8u
HVE3DK8La92zHeAgjHQFicm4H9GuyTEdVUU6C4AVK14lZ2ZBPVGL+ecnYP3sVQGexeAz4V38fghM
eJTjTbAT8SgtiRTQpg3kWGPrVkputyXnTWeoAFA9bae9jeEUhL5uzPwe5ByopHsp8gVQdSy0Y0/j
3AU++5LmjZ7D/+3a4ocTUirCUnr3MozDBOeYhzajisHIBdKagQ1smFmlK2ZHtT+dQe5S8kyIc+mu
bWy1hjq88lYwzukoj6PtlTBq7o5NsyICkgc5C0xKJh9LJi5n0IEj9udb+W0DKHVlR2p/yt9uo26O
hyE8Oe5VwqlzeiOiLnX1At9bW/bnSTt1xQFnZ7jzCH17yVectXqy85hC4wTV3VkMgNunWz5O52ME
QA2ANIO6QGsn+CY8cPifpNhMoAykcOFA+0xNJSKNvrBjuOcH4AumpBRqBojyhmXHd9PcKt7QWZ9e
Cfh0zo/exsM/76rpnWxjHMhBl1hpEnkmdi8vn2XfdoKVn0etEMeOqftxM8YC1Ib4toDK34W7xiCM
gqk7HZ//NG6dBAIWiTCd6PnBPKrZwR3771Z88+ogJdJFPF/Bk9F2vhNDlXIv9k5Zsgck1kDzRwQm
kgVz3mMlOExSVyXfj/hxFPjtu1jEy0KUDMGAwM8DCT38IWtqWpED3/Yw+OtMO2zduycsCMD+E1VS
yfwU7xK1SISdqivyUMKzVgdiGYuP4Dn5DYgUlQTOhA/eaCkYT66MzbvXx/tC8JJT0OJF3IIUdKXm
0v2i+TBiDTB++IHo3yWqapXa7On5c0OjYADrZXAI0EOnuXeCLfNq6YVcJM5bYqZf0fRNCCOFNvCL
KNQ0txgyQfPo3xVXZHTGL6mW7bsAWdgJeHGG7K+0RstPYPdqJses79ZcNCX7DPwhPd0CU6cdL06C
Tp7bhUimaLdsCavygBulktd7fIlnpwZhbMxRJ3oI6AQ5boi0kM8u6inKKPc90+w/aM+zwRuWtU7N
Gvt6XiKoURvcwzIZMDwhASKmvCR4mv6EDJoQtql3uKT5943z2eGztwLMfZ6gxmKy0+JjX+3R7n40
g7hb2zAxGqKbOcEShyokWk+CJcNXH459RSNF13G5pQczQYoGm6+9OJDbAFL5N/iVGK1CnbfalyzD
3T80VfhHnSfi2R1RgpTXxwxAfurUx1TbgomCMjMUNDRyT99UqyKRuFR0ZmtJbCTO7anzTB2KVj9R
2keizOB6Jq/okwNNmapRVF5VkdEeasdoOBViuFdo8a65DzgdvY21k4eQ7i83cypY0FruUVx9WPUx
Aj6bQLRY8IkIyB3ACoAYEu4n1BC06sqizKkhPPH0LEPOTfHL09sRv4RuMXyNnbtZvhUQSOFVu66X
/Lgskxt+wtLmh7G//KKL8/ZnAoE9gDy1MkHYBkF1SxJChintczdbn5fHGUMvIbf1V3BfCYCnJGWd
zVtekp5CsGUJIYP5XushP1uxHOjzSk53ooE54o8kvoLw8dosP6UoY7qFqFl1D129G/9B8wyVg1u7
z4rSbST6IfNfK0ShIuzgKW/aOC4ECl8NV1bU+WVbBPdWjot8ie+/O8FhTIxqXURuPP0i1LYcCSp7
oMkI69pHqnAcB4FGQGdPRz4uXv4mf6lcjMV0XWbzXUNTXPOz6o73q3UKYj5/gA1dydxRF294bKK/
U2ThL9YWlxTF4lJOOTp0mP00gjo3j3YVWZ7w2EezY6tOs+oRrEnGNSMj2xYqkXgXB4V3tbadmW1A
qRYo1oxbyislHQittki7viYrzlJ4fGvgylMWyOFfhz+cAAMNCEw2QTU7hn+wVAJ5Baa/Lwevn+YE
3XZUftiG411tRTeqtJrq1ov66tKnTNf4DWnCRhLTHeGjCuxvZLgLacNXZ06VrVMxfCH8lSk/gDVv
21WzDaccfUwwrwRlnc6mIV0c+3z3SO9BvZCDAwud+oYeLrUTI+RS5hhpe2YHL/qo/c7JADJGo7F0
3H0zEIJub72ckLvvnar+R4p5OW6HDytrSLc0c+WYzHZ97GSiGoE1v4MwjOA1h2im/9g4SVkehsWz
ckNHxChLzXbodTw9won68b00qJh3iAsfqvjI2qVMdtdOmQuqSlDsZLUJxkgqI5fmx1qk1CpCsjhI
SJWA+KjQv3mwLAbRdMkiBoigvYeszQW8HS/beRBtjS4icKGDh1fb3L3D+WwfVgEjueF4lb2dwL0k
bq5h8nJw728BMxx7VOIF5H3BCkhAOEp/AhFRV326OHkDuSrBZgoHwk7gJ2hiBDEshb+KsWcXs4qn
rCmqIkOD86p/nSi71oFAVlj2XJochTZMVPO7qOfle70d8sd3uWkF/qLVn2cfXsLT7+Oppot4NI9P
yZL94gEPASi+n/enAXS6PaYxPFNuwMW2UOJcNmNGNagbVr9zzU6+rcqSJP9SLxXSd/tYT30XsKBd
hX2jmUr0ZtakWD/hZEAmULLI4oxsi+5yQzvMEl0f2Q6WJwUbAiuWutAvnphvDI2dHA5mNTq1VwRX
63YC3o/de7HDSyq6W5OFdk333bWxSW2mNQPnQ7q7k4b5WCLYGEn7hQ2ypFlB7+RAWWv8I+Rbw+Tk
ZiWCD0v8pZrkz89XQ7g2sD9ifoirOQb3k5OrS3ngbq5qw59qoGrXONGt8t1aJaUAYFqpcJguMm+p
rUAZCavg1C9RAnaXL96GpHtJ5AD++hB/CKoQPhKu40tLDn52U0hu+Ws4zAFKyzjNHO6+3orrBWGY
ypmL4WUyc/+1a/yhlgxAzNh3Z1mYixd+T1QAL2JMWZxrC4Ajyg3CCMt97Z3bJUoQwtPSGR4Rb5w3
UKS7oYE+JN8nEkJwnuxjT0w6wE+QuBabXc/0Vm7z/8ht7hSnREBCX8hVHSkJKR+us2b9nkSyyFaw
2CsRwFN4DknnDAs7/Q2C2qmYJob5Eq+F7mbSL18SzFZze1G479D5xryyI3Hy6DPHRyNUiDmpoQtK
CNPy6S9QxN+cGdPqZobEpijOFdmfLe8QB29ws/HN85PkrTlYozfbX7Xx+h7OKqc468JUpP1b7ys6
EvvbUEsvQT7pAerLOJ5EFAqSIAbsB9PuNFOGHDaePe4tOJCJolRU+lPeM0SmlpO1mfA+3Y3aUzpX
yh+8xX4AN50hi/0G0HtJSgBxalzPqGp3e0l8+kgEp4JoRnYZO20m9UWmp/9A3GNzpwF1zdfRCS3D
JrFb/YuP6AqUYKs3CtQ9VX8vupFymFlSfhmUNQUsxu97l7jS7YKq0i8nofP5+jCzmdniOQk6iJpa
D6Bk1kLbANc7eqjvZpXy8E4pxhgzxdhu0VvFrSSmG1AxeawYniimDvVoJPbp8rj5fgGEsOixckhE
I55IUz6TGFqyfJ3oo/zc2IZTEmGwb7z+je86ntad3wG2m6tjyaUFZrGa4PMEt2i4t9fmkeGpfMgC
P8QSU2c506QkC6eTE7pUKD86cb+R+axXHf2abZo+PKKvnhqEuOtkkoFYWull8QRztrumtm/fL0C/
Gw1IlR4agPObAfvPXRHhfqeAdoXlicKQ87mlzVR8GkLPSBdp7C/WVFQQvXmeD2FdfZasVH1C94zo
hdt/KXY73K+v57LwGJRc5Eij7RcjL02O5+i9W3dpBc140N9SpKRfxOeHILSnTu3LYEQonAk4zXOj
8G1dOAB/97zw18OY0Ab1D3eh/vajSbBYxbZQRVTlv7iYmGyauowrH73dXD0xGar/FE73r8PkMNhT
nOR40Lbtx/sorGGSFp0b5VJJFZUKD6ophdvrF6HLz45s6BYY5RtaSBPe6n/jEcTgwL5Bx72a/iwr
sypmQBrCq4Px+jNM7uh7B7lDi9PEqcAJAk/+dW0fPRQfRwrBO1Qr3OxkfWURdTi34vrx3aXeLjqG
U2veDTRMpMvPvmpYf4AZV6qcg157GyPZogbF0qDc47bsAevFA6V7SQU4vK1QRvegpNcR16QnU/4Y
HOgh8QjQ6DrJQXiQBY3ynrbSp35Luid3VR+oXeQaN0vxDo6d+kQlKLAuQ9GDtvtJ+Trrcw6wxCp3
osOP4GL27Sc6awumZcMKg5aZgbnHAzwTtxhOT/T/poitR1G9HiWBaTwsFVoB1/NDyAAPYxKv2D0P
9QY+UBWNyjEvHeLfb21fWnc5baKAZr1BTpreaIPdOYvSLN1/nlawEo4uHtc1qHj75h10ser/r34n
teXtfIOnRCbqMe58b2oxuYfmMBy1umIcejtG+lMdnlXBo2amy1YbtPQUCsI1R8Fqs6vordKrzLjA
jKwM84nyYshdAPhhVjWUXVqNnVMJ3Mn8GlDltYwC16DvUxNJqFicYKsd7XEbWxQd96dcjE6KWB/M
S1t819VbZjF+pgPG7hDjMp5q11o6niiRNUPgcSz/RAs0EpQVKidROlhv+Cf5Khz57RyUAhgjJcTy
z2AwVUWcbZOTFcg/5VCTAx4yyw2Py1Hb88yFUbP5M3WSOBaUdcILXgLe2RDZZZGtTQhm5Nh7lz2R
SOSGTNHN65AEXcQ4igniXIWlQYp8a4iKXg6c36oI1NEdhqatzKecNEG49imRJCswaoJisw1SCFM6
rwnpfrBCG46MmW00OnXB6LDEHO2RLs89SNZlm0ZTA58A/9h+ZfMDh2NWgMRm6X0SBtjF92ugDDSS
PgRPzQw134JmpDB/3PPSnRSCxJFtbHCR6pq0fSz4cQvwvYu+gL3LoILQm6cZ33nRnAIUJukSZody
ncBuyzx3EbPsBE9aqRHbLZg7JBRyszPwl6IY+At+rS90sD9rY5uzEIiP+3hna1gGVjv5wKPeQXzz
0eFxs8xJ25MFy80jF/cKzp4/9Pxk+2aKTwwEFZbXkmPgGIBXlZuo7nrvUYPZBL32S+e3NAHHVmn5
Cbm+h6Kn7WeXOFGbndj5gMiYNB4ocG50s38SQiaP9KY3Zc2+KcEQ45JD6r8HgvBCC2P1W8FGStmu
tj3if6KBAqZTlcNAZDOfHxwg76YfxTmS9BHyu82LwcA/gdU3XD3Gl+dxCscJiAYxaf4lLwVIUYgf
GXwiMNzQobUMmFAuCQftu5K7xr+3xvw4zUFphSSxNvCL4dxV8CL+FpHQZiRp/mwqwaVTFxj3P9o3
jtniV71KdzBKvTXsMHKXt2p8ILIrV5Adsb51oW8YKhYE6TgQlZOgeI3/N8oklYWO37na5h+xppO7
WEFoA3Cgo6BnczzfdUcNytIwhyZ95dKYGUvoadD+HhkCyDz8jSZNmu11RhrxILAR/0dgIEFaqtVv
UZZVXosLwIowwV/a/IK+modxbz3PKJSI3ODfDtiweJvfHMmVNrRFgY/FuI7nW9BY8E7zFlKIH1Bw
V8mRBiSOzQIIgnzFd9Kfar1KymUQXWWurC7F22IRXafn2x1zr2p1J7K8mfcWqKa++RvKNMUX2i1t
Yr5y9IQjp8DJE6SyqaOEyvZJxKBmLiXlTggt9D87mD57ECmNqXecrG3OfBKUdGYiyG75e0HwubV7
Oib0UiqO0Xlsus6pJfyWxjXzQfswP6VkVeymW06bm2amygEjTxAnb+cgar0mB+i24huvf5T+rwsR
rhPvFISCm3J0u0nlSuaHPTKVXDfbM+KpX5rRd1gaTuDC7/qidaoXbrpzVy1wyPY/soakGXznhUoL
my0FYP9/Zaw/EY9frU39ibHuwyKzZSAyy09fsEstHjOHeB1fFXycEywsNZhBtb0AHnK2hhbeERqD
Gvng0CyGAWnsm0hfkGfdcsYb9+VcpheSIs84KJ1rJm+xff/O1nwXppaERYDU29Vl/LRGCgL5BGTe
SKKfaOOdimO/ihBOOxsIlqzWcGxTaLcqyfhCONXBjInMC0qScs3ISL/ZdUIku1CBnL53Yztr29vt
sSCEbKJn9REmW/EMMmQx0iWSYD52euJ6ncVWMn9fm9Bv+DT14NYOgWHSRrkASD18mYmbkyZfk/eJ
wfqX70FPfx7IOynWIsIb8poYm5BcIdnP6+bXee/D0IC+i/uZhIK2POowLP6+z0mFhJ+0Chhw156i
DU2VzikzGfdCZu8qXh5vWd+nUNOZWowJMKyWPxOS4NdbW1SevYUVxkp/yhnuK8hhQnit9SvPKj48
Y5cor7dTM9xW3zzZW0te1GctwSuPL9IHew8qpbIIdJgfOaxkqxDtxBQ1dI1kg8NMsSjbMkbkt+dU
UpXsLALQbgHGpnoc0a+R/w81SmquzfNZeVY/Tyvmq+kPT8QePfKn/jydEZDIeYHQY/k2AOFk7bw2
VKcwl04wYPonYoAyruh7pPkpwho+TELUlC6gjFc6uc6GsJcT1w/ofnanVvwoqOeKPnmXgFH0lvNW
TcHqAdiBScbZSE06EiGh1AEOtr7YqlLiM8wUBUN3n1ua1zNsKs9sf/vb9DlI+VfNZsDBdB1XHgaH
zxvgQPaBpej9e75wpeaoijzRkgbHAUZrEljT2psn+hvSUQd7mnvPBGVCS+rYV00IpTx5z8zTecQ3
uncQfRAs8Ygid8buwKoHaSihp0U7oWBl6HsPt3puc9gX/1xSdZMD+Hg77d+XccK2hRUMVuzhUCly
Nty8W2zVy3EXpDv5l90Y8Q9gWGQWrRaRkXP+Uy1uiRgXgYut7+bobxyiUxIF2XmfKcirolzXUVsK
Cl07SFQRkwN3CLpK1yyXNDVZ6WkC1QoNJj29HP0wwPHqWNWYjxqnaLAIaiWzz7MC1gGaJMRDGibb
Qycuh6DxCf4J91w/Spie6a8BFKI+QQEP4D7pcM7fjexaqsriH8cdpLGQYU1Wh/1VPmMeXIGIh6dq
BQB6MHLLzUfg1D3FyGag5jRE3529W9sxdFv0trdQVojFHH2x+Jh1c0SYux2dSYkQAY3D/dOU0qZW
Curxs3l67ySnLembaBvCHdVI0dJ7SgXcpO0u4Je8SahP104ZvhBQv28AaMWzl42Y0nIWt7RZjx2P
UKOnkNUn3v7fnqC6rbvmQT49rrrZkLvUu23xYT76vCYNUa3CPNPOPDfofa16wE/vEsLg7e/MjCQI
85Tm/7rGsc14N3fB98oRzl/X9EB/ZiwtGK5vRFqSjfO8ussE/5U/sKDlow/s2hU6ygPBXIBTsRHh
+Dnmz9DHC9WuWl/WF0RVRKlbHUCbGIkIYC2+xxnAMyH488ym38Qu/Fo/K1GzM03P21Emo7Vt9d7p
O/XCLxIDYTW3sJcUB/2ugYSPPa9tmZ7GNmtyV0GrNv8qzgjLWSKibaDkzE7oLHtC40asa5+HTgJs
FmkWkS7C8JIjZBIM2lBTUHu9e41Sf4/a+qxyUzVuU533Inqt821aIw+WjSXkQXPhVYRy6ZPq5ETY
B7nHM7zdvUlONNq2IXM3kt5qRjfYeQsxTnfnHYeWjLDwQlg7NLcv9UdxgPhfnplMvtCp5hRFqg08
hFZ8dR+1+K/EYs7SURyT+6xO15rDEkGLkBNKEdyRbjZnU/7qtXNEhc4iY/nqpGJ4mCi0QY2MvibX
TtEHbDO/XCgLQlasE1CpfnnR2slkmlHCv104l/cMpfpQWLK4GBMyyCm2HTdJh1fLYGRbQ7qoCOTF
bvF/fgANMxYoaiCPBT4g5NvsscfTtF4uNt+NumiHrfNg+SorN4A1RgiI5sR/RVBLBMJ3uX7uPOjj
t28Fd8fME0Rg3RzOy3NgflIKX5Ep5bUmgpwU1IHVmETo/nhQ3Z3df6YEGb+kUCxQBBPRu5J5pH4K
qM/Icca6kQ2oTxjuejLkW26DVwLA7RMsVD8SFv18NIVL4lFVkkV/PBPRsnWYpk+tD65nrZLhogfc
jmXqiuC5xRiEdfd1D/mKCj4xtJ+uX/xcxUiTk8EL5/FNoabwi4/IppKfDrR5XIayWToRcg3M/TYX
idyeiSYYhMuRxSUTkC+aIIw0GuhjewDOdRrQYazXCsvsUUwp0aHV/juTMGIHyJDTomyXg+Mz+Cs2
pxzGootStFIkFbsD3MkIozWg35MR0Mj5NtwGcAkPMXn4t/kWEleaeCyZ7go8MaufOoRJYZoG2jp7
rd5c2NEYmcY25S0gbtvBI4DOlO+QGNgBTv54s8A4zk/KcTklRbvOw4oZziFxnOUj7/DTfDc1sweh
80frWxDbcwM93SplEedZnWmjzAdLaUGeUXAumQzc82ke4bdol9Xq6rfhPdZ0Z8dFjIX99QzUFKfa
RtKqvg/qcrjAZ8JLvXvlqFQ5rH2VPMWU8w1GSDQBq3qVYO4Xhw8mUzLbzqC/JK8BXKB4D7LcfPgk
yB4VIb8r31UdfT1JDFXHYNvrCAZNN0hg4gFjeQwK0TtNDcySJ2UiOy7zkQADTfrrC09Sc/MSs7Ei
c/phA42dPMX5ePiDzqwb7OJC+k8CToC9dovsRCEsoaWyAjEI4ALhdrHHrhXQiQ+KXjXWrZUY9XFM
GkW7jkTMJFenXjlhYsCJ7biF6C64hV4EWlQiXt6xBK9s/StaDrROLD6eOFH8h+/x9PlpCLgLJdh/
tVTZSaGI3ihnjIGyPNQQcOcDDLKh3aSe2+C7yrPTPbjQcuHM2ooBIHh2DNWNRSTNZhgVQFZYYfVI
T3N/Sb7aIL3JhssAgeUTd//sfEjcZwxPTF/7U/MLUCfCvDjYE135RCvB52DVM5JQy4a+VwNO4L0Q
UrkUAr3IAprvOHFWE/MGdmvimZUPRtvQ6ytsTTb1FSsFM7VDejWKrjpO6GILtyzj5pXmBTr9snNb
GgkcTnQoOEULuYOH7vPIVznu56hXIUbIDqOG/ffCfqJSYuBhIKsTEHhcmvPkXOt5HL+6R3KBHe+5
7jLNCTJhcnM1loj1gp0yTVO/Wgcc5JBWyKtZLEKWkqsWvYPLE30MP+hWm5v5SVeGetOp/gunIu5a
fhEM/rZJZt9lv1cLPRpKvOdEamujtuFVwM463uXw/cduyfDcAJEY99ohfIqGdCg5cxkP3gzd3o2y
YS7R75EkZ6I+z2W9xddcgbsSs/dAegBrUna3oHZKiTCJ+dOHEP5ikiQasEVGbO4Bb76344uH5FQR
uMKV+Zrcv+ZF0xCLMyO85T7BomGYm3SyevU4ildiUCATbKE/mZVnFYrz+Pg/kMQr5CZLU3UJTlvc
U+wC5yDtqoDO+u84h9ct0TIY+j9PRBB3/CyOrT/EpVR2ms4FArEoBlTDIxmfdblNw+NCzYgDSWVu
YXQJPRg0wEU5KyrFwNrrz6Mg/lNwtalzW9mL1etgqMk0H0Hep/jiN/o/O99MZ3UWTjXe3T9N3ASn
MWts6JkAwEa/fzO2FO/Zp8Y4rdfMvq/GwiupnfFLntt27TTVNtjU7xHL6LOVB4qI9Ugkj2Zb38dM
lDYy1OFbK43xywiZD5ubI1joPHR4pqYx5sS9+gS6J1QfuCSolVyRv9/23z+BjY1VrqGXJV8tEK/h
pQYmqEW0G7AAwZZgZM36Uq2kP2lEgss1bqIJimjSgeAfiWAGuOfUUNs3PtLEJzNQpPM5GLuHvvCq
BsDoFBZ7e0e3UBmsvUWroh9JB4IKC6pPg/bBQpyHVuAAnwiyyN/NeA398GJbLm+++E+BR+ZXLpTf
gGKhJ1JRavXFkeR3SucahL6ty3xyOLPYnKwK0kfT01PbxWr0rG4MVZc6ne+gVqemlxb5Bc3YKEPA
R4Oh0t8jNwEvOkgr5/zYKx5a+IWumChlgUA7GmTX6w57HKiO1NYRB1L//Nqo1nhxoJRCIr833ejo
Oz06D/yL0NMoMq5psYynQMPp+qsXJlrITDyQPNf6wyNqtEgWH+CONssmLeMRzpL9gk4X3rBHHk4Y
H4rxmNfC/zHKutbVIc+0lpOly9+huBX0S+L1mdFF3dm7MGzsW8yrURy/7nbu4521BaIfyVyS1QOy
UFVct3kUnF+lsNULeavoRTMxqX0C80SAW84Vy8DO6nQJT+fsKrqDZJyDuClOezbZqp732NEhITvr
HxEAdpnuvATpXqGbDGsVrY/c8jbF9Uf95pxEUduHTxqcrZmQbCj6aFwf8qMfRXw1FUeZL6G4oR/K
hm3+2CQPiRG2Cv9xAzNIaoZCUmnLfd4+HGKbkSg9s96gHfZPFFonIFH+wq3JlJzPr3K3Nmwshbz8
yT+g7bww7yxYSZ697qWstISelBD49HvBQc436sjXZ3jn4LxzMwQFVMDM6dBnIFDTgJEyUMS303El
fFEsL9RzTfHrp0aWs5Xu4BK7ZlglyQLn/6dcHDg1jeXfjVTQYEvIXsKyIP0/ehUyErX9oc/I56f3
fOrb26pWxXWBo6GmhIqKGLuurcxQgxUUCUFOS+1/AirV/kroTYKv+64FD6ExN5gJkHMnd2UBZZEM
8r7qtA7WemkUYB+ExEhXbjzVaWMgJXCIbgiiDAw9p+SANTqfK5MVU1VXm1xExLBFX5XXNgPnNHuw
ZnF+KRwP3j094cOljMgeIpo/swjpzo/RaR0QmUjiPJJ/s8LKzv6pm94Eew2vJ0NQUI1CQthWpqO9
2EDJ30wp7MJ8CquHLzxi4U4xV3px6isKawY7pH/taBX+nyReZU1mMwzc0mDm3HJLyZc85fsJLhyc
U44IE4r8E0U9mUmduoR8YbIxpnS9N2ADTF/0kke4IVRTg2vGKo4qoIM8Mp9VssjfktVwAF4HvtvW
D7rpS2yoMHVgCCEnreraK7Eabdj5nUv85WwH1y/TpcLkSLc8/hzbGJUWde7PZvOCEbh47B22BWfd
76nFFvynJE7+9N+Du2hi7go+Nig7tst97yqtA0cXQJNZ2GS2X8bTbJSRkTT6c4ZPAHYNDh44PWPA
2RwaJtrQKX3+c5SyzMQS+db+wRSKl2L3rCvBCEZ6rZAmWRZPcJ/TsjXlqWMYCAWszYaNEaiX4pPD
Lbxn2eZ3qSpxYN9KvXe4KmDwkNKIsdyPSHYMVi26pnBKEeuh9L5WpHVWAei2qzkxVNgun2SW321i
uPZtC8dFli7u8t/H/5ZBZNpuXRI7xN0IgIHGnh+RyMq7J9lZExGOjMuw6iEk1C+vxNcaZF6wBUdL
0YfmN2vSq1POGgM05GJ92uWEhZdARXFkepdwxvJz25quhnbayVmcYs3UP6fMaSRLAUXMt1NFB76u
hgpziJ+ifLatCLjqaBCUAS4Q9y4wHp/jWOlWVw1/RxQU4B+0OBF8EpJvUJ7XSpIAC6WN4vvSHm3V
8XJ/XZ0VqM7RfAT8/p/TKx3ppU6piRCz84iBUOvtVjO135nbGgjxwuSq8IlokDo23pMNSNo1vixe
UM36RB88JuyiiVjOs5zNMdOu9cuqeCFZIOvReRzLbkJp4hP3jPNmPboXpKvXcD2DH0HRKqmA9C+X
I5+lJ57kDVuG7bjE+MjUKbkukMq09nz12fpw+EY0O0iC3APQJ/EW78QMsGH2yPmfByDEr9HBm4yT
MfH6Ay45uQeFk7ZKWwP2kmKMi+w27e7zuWTn32b6btz0t0SkqdU2jRWbIQe3RP71DwRQ33ror3LF
YamqxK87IsUODN/4tuYV0XparnpbBPZnmQbyHL1rSi4Y2RBWiMrKpZu8XRijwlwvCgVwrsGdqD6h
W5ctkPysJtnn6T28+6AmCtuufGvXl7drPc/a5ovqoEEOtnUSPrtk3pof/aWzjJlzaNk5MInyuUz3
spYhOExzBL/xOyp2r5Z+cFYv6ZhY3KtLd3vC2wnAgOmkP4/YYrd49IGzwTxnPAf+Kgc3ra/8GOiV
M2D1RFzDGuauMyno+tdD9hgHbba6vHqUkdnCBYHcgad168fuFDYFQ3n0zvusQSQYUFowCChm6QVz
1FyHqKXvaPUSEkgvIaYwwUYy8mpT9MSwCOopGbBLUHMJHkEVxXHfFYeyT/5bwV5C1WuLw4vBt5CH
TX8mfFBucITL9lLOgxnsCAcQTFuaYJHWj8jOfOhuNpOW6dVTaw9rIL0Z09ZdnWidKaZUJHyleEFB
oSLxLR4jgmC3ZEl7n4I5FgaqWtNraZZs3K+Q13JX54Iy48K34vIKmj58ufEHXLDIsKba5cGcx5ch
6HMAkOsf8l5ucmiDl5Tr9lO8e4z39mKwGKXuHNl18pE1T6V0Tcz+iK5ttIPwXZ17RS/QXpxMeC3w
g2n6qASo57zKflsOhovvffpxycbgk9Gu720gKU+3Nwlw86tzQ+7fEr+yKopiGnR4bF/ZRNk2DTto
Db1ysQd6SHV+oNE8QoRU9eKaqX3pWdFa20wK0grPMmKm4Gn3gC7xJEP6Ckxi9p7l02stUGCx9NVe
fQdA8ijnMSWqjEqTV8GVBE0T7Ke4DyHK4sLKi72wpfyyhKJmvy3hMrF25LY6rOr0dYKYlfGcRx7Z
4jtY79j/XW/aZzvOdMb66LPqyBblL4JsBzN3zEn0J1omDh6aJNGs5kyJC5RmOx3Cu6IZzbDOr7JF
BQ40u2+p9zayVatTGWpjlybozTHw0WZBLu7IxewGmYSmFbym1BhWsa0UTOEzmgaUGjVtYeaFqxnt
4Nj7FmGyhQjOUPpwqeEjCHYwxR1fVPndwTsww7hRWA0hV0jKmlHnJm99JXc9dngQyDK5NcnOjmyD
AnK/Ggz2K8KWB8AEDx/Ms+5LibWcRu/9AnR9E0F4IcAjwZF7N98PST//t4Ydwbe3S8CRjblaeOFT
nGtmiy23rxLKXhXnD6kvC01U36fgWa9/GXIO2C9d+UhYzAVOONSWtFzGLP5wLX4A1fRMV8xRxoFn
ieyK143/RXzvuLQEsVhQUthVMffeKfVfCU1cmRqpDd9O3wAJhVQX93LGpCFbHZ9DDFLU3zTiiSkA
YNppAkF+uYqmd5/Yhn3FF/zLXZPXm8SYEJKoSXEB1qj9SNE3WwAS0Gaw4uRS96Y0m3gEk39E9RDL
DHo9+2VtF7fMZOctrVS0DaUzVlwl/6ECxF8DiNFD6vyI3mM39Yig5TUA0bn0fvTWXSGD5wQ09mWE
NjhKGaxt+2rnpznhFbpoL4x4g/IzETK7qNy+I4hCJW1VQBQXjuxNUOycgVmmsL4AAy6FN9tQcov+
NqHV21jl/vLqP4IWR9ijSC+sK5s0J3dYbprLAW16BBMOlNLXnsWJEG8r4otMr1BCwEHAJru64tVx
kVJ2YAcueT9fXj4oKvOaeGObZovsgt6vwWDbTI8lrqlKPyCnlXjMuqBadJO1Of4oZdl7KTyd0RhH
SzOJnuEmVXSufLz/fO/F9teDjNzfYl1J12NgNLk3FLYSFnKN6HomF6UvhOBhuCqwNAIWzb6xbjJp
g2KosNquheqLd3nBXAutGxC4kX2KNYepSBUWCTXZz4VRHjC/Y5OQ/vG8heS7oFSFeYzvn9zJwxJF
dSI+LnFot7CAt1PiKHQvjl+hRPe7++WGVQu4r09qZD3PTWM93nm2Q6EXccjwOso5X9sCsqyOp40+
bx0pGp66TVzz/kHzDnitpAHvu7+Vx+kIQfV6IHUGWsfsEnLMQzFJmOqVDCj8cXV51ahwCLV/x4wj
uM88eA0TKUHBHC3iH7EWsJRw+tYNKmITdA155CNZrAUeG9piGmK2HWMBeZqWZNzWQPyDZU5RlIxz
0zQxlJ7pffEKBzOV/xZw4JRHGkghOvpNngDK5EXCsqPEsbua/0IiEpy/vDeX1fSKF3t2TQEw6CC6
Bf7MOml14qFoEpmQ32Tg19f3t0oGgXUBqjoDSpuM9gThRUrjzh7K14rbzEPE5777XtPTUJoP4vsf
9y5/TwuRKQ7yJIdUcXX3ytN0LI+VNZbSjhkaPSYWqMW5khOeXLHfXoizcMengvuci1aFdYAueRUK
eAUGGkzNvrrtlt/+97G168sFlS4xvR2IfKtRanNX5gZKyERlc6qW1LJPx0QW1fU3rOXjaQbLzqeL
nQKeJcMjWPSb17etxxIpq21XEhLIGSisWsfTHSCh+mS9QaZZeJiII6JakqcRLwHRljpIIi7XCAXX
Cgn+62GY5FECHEoi8Z2S/lT3p5gG7X4U3DjkADbBcKg1liYAhugjEATT39Jmc0Tj6Dob85VPIJNd
L0A7fj4Bx5Fhg8TJGpForktI1/E+hYc4upt6j95K3W5HKYYXqNT3AMWpbRuNooEroKUM8bRXYyvf
PY6ai7/gTKFXgYmAQHm2SmrN8rPluGLKU/IYMca4bYQLLfWM74pKoLY+IgSt6onQd+2krFVDlJWv
XEij2W9hDu7hEAowNjPbBmuk7kfMlYUSonwLt+1CQZnWuRj5MUb/mzZVNFkRP7WlfVzq1WkgwFT5
iKvSe2mGLnTxZZTSc3FsTn5Ersq27LJJ7+m/spPGqXHyVpxZQJrbUKhD+yVF72N5HkO+g2P8nwDP
rQ1ABDTOstACTSGc8459yZG1jbkqu6nnnghmJJKfAu7WYX3N+mp8VrTIZ0I4JqOIyWH3YJCDQIEq
JJp/AQUTxP71XTJIQlmoBL7xIXwULdcBSqUXE8ova/05CKhZDwVq0PVNFCMQ26QP6VfE/psETq/3
EcTZzWlkRk/ypBBL1n+Bkz1fAJyUrItuecGT8GmcrNOHJNc5PozS722a6BGSiEjWFePI0a3gEep1
R2MjR4G0+73ClRhhzgYnBJkRgtw8s6gcLCQ9T2Q35L4cz0ZEQqjy0wkcojnVPrZAE+KjkBDExQJc
AlEdeqG7H/QYtsxnruHEoBs4wXmPsFbL8AeHCdE1AM1jYFAptaAOHXuId46iqfBGNI3HSsx+Ezt9
+lLWEMPrCvxlmBpm4OM5qE4Bku/uMaT2NJmW37FtgRJTvsljvsdLRIRDugoiiL2RPU0I9GFT+zHx
tSfT8NE0R5si+1Xe39Z1jrjPCA7zDy83JAfam33u5n2IKFAMzvsE8scV8TY+ofpuGE583Rc8auCw
JiZ9ylK8WSrfsI1HHBD+a/dMyLHhI6n/jDDVYdHo+s+zBmHH2Vo0xuA994dh6ErFkElaRqev7mdz
xFCpWvNa+QHF/oCHaPN27qP6QHNWwesWM4TBRSiJF7NgQo390mIwBzFgFYJtUKYYTdTrXeRpAcxM
GSF1W93zLm5iYs1e+6ioaN3tb8oxZR9E+K3aoKjjqnYm0cyrHIJ+Pg/NmURPUVOkmComXu8PqxzK
u7A5TYqXGmZtWvEBhLiNdV3XAPRxgsjTtcWRJFE5VjQD2uTQI4vXT7hpmrGTY11mkv9JCS7Sb7f5
85WiwWnslqo1ARCSMvqAzLVeaLAqCkWqP9WmQdJwSPXf05QMujBCFA3GcjNuZqsM/hIb70JDOT4v
TBsgi4ibyjVgyxcBdDuV/bwjZ2oi/kOUAmgkv2Uy18m17oHEEdcIHY0p8LE9g/aaWVAjWelqLWDY
6px21C7ESb3T/+UPLukQrCMzn8s8ijxn2aKjioJSV6BzVvfQ+D9k/EXtlsSX7V0wHCVVkPwiOeTf
Dfnti+mLBlRxaBzy9MzDY/kn/QjZnsfYR+OcF65JHNnZhRYgtcNqOzgal6KxU0JqbI/OwdR1gvu1
awzFXbCLkEVZpKmwtV0Dp95dbLGHjXebZCoLAakWFpHC5H4va3tnGwj/uzo8NfEUEfg8kOgJDKZ2
GJtOk+DIHV8msbeKpUO6Hc8pbPEhY0FAieYyWthMBDs7Fm4gbOPqazEEaU1Exg+Gu6O4pEC3+J/e
l9lODwLxQO14amCxKiJPVhlGFIq5uzW8vU9Yr4QTzIPy8CW+BeeU2B6NmuWGNcAY8p/LBERwwlMY
rjUu1p/OLGNloB8MEcmwsvyYdd8K2ehNI51JlZvzCZNXevpWtV64ViZoWmXearQQMp+tWi+fMF0C
MlP3gQSMwF1lM9TVwgAJe7jK17mABtatDl0sXaSmbLEL527sp10+phOV8w+M9js8HqxlaZ9CUXYE
3S9xxRfMCeAWDtQKiK97BbDwvUwJ3qSuj6l9B0dVIyyZUuyCLJm3Nm0KZ2LDY9aUyQWakUucYYO/
1YmLSV3c3L2KrA113ivHf+QIJEupOFNi0wcAVes5GSwNCbGDSkzc1GPmNE4Yzc11wPR01atuQbpX
UOIPK799A42/LgI1nfcO8Ek2C19QqXHjLqk2PpoCRMnIrGisQ0M7H/NrqFeedvT9KPLyffqjjGvA
5KLXyjV/kiRq73PfeA9tTqPmI6sJKkYUDyMKcxEGMXwJ4zNybEhMKwajxOwqwYKOjc6Qimx3p/Vp
EP8jiOWp9J1otpDMpuMf78Br4vLW0sbLs5wLZwhFAGHpkpt3UIzASwSkEEiFJho4efNWocW1C3HZ
FjCbMJm9US9Kf3TSqh89jCEyAFduDJqwNYCed3Bhdm9/hhXGY1FzRMVqQx6yCUJyuCHlslvi9GuW
efl614er5ZUIuXHYdQ+9xJEyPeWT7o5qCghSsOwoFOvHemws5gsM0LaLvOclQ3HWiKiF2yuAGQng
wW9ybnOXCl+S+Mq1VGc12MmY/g1bCewG6oic5IN7StlGdOVnFJu6OD4/7jKb5ylG8Vh3T0EpVxdo
84U9W7kQCUYrWGUZsD/T8Lf8tTNv6naeemJPaIERD1oPf4p6fS9fRamLbOrNhqSxMTP0sIDl6Qke
MI8A+Sr2O5kythwf0NaorassMqkYHhIJ5LK5jvs01KlE0nyPvR24El1WoIiUJMP0k5qfXPc+tseb
osZtcAeK7x+fVkA2DY+UmHn/AahyUsqIfUM4bzOjTxDo9IBErX99cncjJaxKr4iy3YfIJvWI1aJx
t+kKsF+NkwVXGZ7TT2AXBJOUxGf34u2pJ9eXDO/ARXtVwylkOoKxqU4o9QWgSCBCrTrybkrrOOzU
93bbjRiZxuncQ4s0D+vT
`protect end_protected

