

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
To/0Y2C4coh8VFh6WzI2wbA/wXer17nunFaUIFXEvO3kBprRAlXyefibFdeqGdMCN/jPnm1lnQge
X/HG5CdHuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nnkNk6e3rHUR8DaNj0C7aWkCs5LBgvWhHhtsF0DtIcgM1egO9JMHLS9VXFoTsIgw40ekMylMZAif
7Mz04TLeS83J8LIkLQIVFCxUoXkTdVbP2vwAOIuzbV0fNimpIIdRDB4Qyrb5oJF0cClV9EVhM+PP
xrslkcRoMPftZWbNXzc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fa9acIf/jWyoTf/ZQQ2RdBUZgeC1x0Ej+f6KiTiJLxfGAO1lB8jxkDwdqife8FqrZb9GuA0CC+35
3eXgFQAQNKjhv24q1nYDvGkg1xQe+JaS1IiyitufBE9Oqujx03ehRV4B4wJ5uK9qxFjJm3WBZQeA
cWZiPDwrU8E27DqZYUHGXiufRSfFhYToep6g7NhnZGCmAfAD7Cg9pLa/AvxaXAS9nnGeBo/RPlyk
G/XXEB6YF86+MUOkeRMAxi86Vcag14njI42hNh7J8Lfa4beMq2Avi5tz5eGJq8y6uRjal6wz33O+
m0Nk9SOLFKAmJ/ib8Fpq77uCjrQp1T7Cl70Ebg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h4sQ6/cKFAjr6toNt8WCtcnxvbT2RbQqvunqru/ZMP069wFljAWXbbabme1u0tsoVT7hQ/OZYU4t
+qXe0sbPKDx8M0x1MxaKDasoQ543qKQAHxR7Bn28bTi4sQCu/+YxH72mTMVFjRAGH6M6e+MhTnGO
FYX19oeiewDQZSakDrY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C8DUdaX7Hd0diH5RVXOZCPD1GItaWr9F/mVcGAwJsPm7j/BsnnF1JwcYxytFDkPy0E+fcaWYKz9u
7/hZwJ449yH3vkp0VWbVjDe3BqRjhnTwAc32kEGR+a+f8HB/6hGM+mJkcuw5DhoveoZqvYIICYqz
iQAjheEs1g2k4DBWxSdaCPNW8fXVd3J/pZQSuvaNRnCtPGOVMt3rO5k/WAzjiaWwDL0KdanM3fU6
uD93ZtkLZCLilGdf0EAax4p+pGVd1C8GYV4+XW66vJmZoT9LNfQ7rG/mL7dKp2aZ5DJPqw3W/O9c
HVwQSloSjbmiN1Fhr9Mdj7iCZycwuy9BYtMK3g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24720)
`protect data_block
dvSYnDwdZozislvFckge1Wo3Gd+jq0ycGWlMojp6/gMCT0EyBJ7ANBJwIYS7fQLxhIpiPw+B1gsP
T8dMWkFNfR6rtO3PHWSgtHAUwQZjA9C8Pjgdj6ibdOsGfpTdlbGULxwfhn8bpj52UktSPXhsYLx5
OA+/JdmLkXvUbz/+ughug8+hhGQv7yoUpq7zDCfSjdgxHUZii1CHZXeWMVp+ip4+V5VLY1x4kvY8
XBjHrB6LFN4cCL1D2bdqRnZ4+x2owCG9IsWdb06sRHZX0YupN7rP73UfqTjO9RxGhmUmcT9cOBJU
BpLzCMQCJetwtoOJoQ0C/lcD2x3QbvwKqf7kzWbC/6pq8ClF3btFN0Ia+kq8BTmp2oySdNfUbAsr
sJHX4jZLlforCmCs/M4P8JzpUxHzUoZ8OpbvCiq3ODvKGYWPndYw1mebWeA8YsC5id1wJtj0kJ/s
4Hm6cdc5hqrC3NEtQxEg89gbqdFTOV1tGtlSlEhpVu2Xw1B5tM8MDIBhGPYmH4pQEnIIYk3JiMNW
eKHdBVlQjHvgelqi+7aHCX4wYe1FTar4VDB0+oZDDoxifoV94w47CyR7RGzVf695mWpUyPgFueTL
vzZrttMMl+pfpPMERTDCaJvkxyHc4mp8AyHojN18nOpSNqyc6BxQoTeryBjgJO3GeETEiQfyWqgN
rX3qfa8LCyypTCpzRls1AwTUZQ8N1KJhdgBt98DKjaUji88C0thvEH6baLr8X4KdeZvSqF2UUTZA
3fuV+wF1MCapCPqeFxExDW5VwF8OfRKWrvmEmgxPaAGo0UKX1kN9G/3BwklkN4yPcG4gwwL/9igm
a41My8vVHi0XwmZX7w1V6SQ1KFRmPqd85iJolXR1hFpQNTv5IIsbauXvMBLg5K0nJvSY+H4aNOzT
GCHLYl1JqXI1L+h8mFFDVWY0FtxSkg8k7vyBv48ZNbx9TzKKV3zsEuDO6qPPGb203Hv7KVgBqmyd
OTW0g6QrJvTik2YZdaBhckz+fkdLyw3DPKAHBqA3jPm7X9Eqyli9+TKuwpPSBKRmPVW0HHjB3YpS
aD1FhKtgCSJpzGNO1IlEtAuOtCrzLI76JgTatijnI1360m7KGwgXTiXHfPTYbECGfDGk1jMk0EcK
LEjWJpoDCFvPCP7nCGUMhjpO3vmdQafCZzJLzmO2E3J8WAwlOKDM+pRs0X/Mgtf9Gz/y8DtLQIaC
d/OfqS0dqQv012Vw2JyhOHwq9h+p1TiHkJqQN378YBNTsNJFoLmvyfSNwqn3jAUBrBM5hPzAcCBa
OSkfRp2I/47/+RmCATV7GEPHHqHgxKB0DvCaSQpAw71zUYeivojzJnTYMcgkiYYDGIAOpAhoj0p7
mcOtwX+114nHqqDL6reBEb+YTIdTfQwf7wqNbkldVb88Law+FRH4gmuSNxF+bl5EleSDaBOP5Fhp
LzYn6v9e7wAv8Fbygbx9/zth3jblDi98mSBkgbpzvCCVKZhPIgdztDu839WHDshP4hQfzyMi/2+A
5nhS6TKcA4xdtvBbG/ZbiX9psrswlc23H2BP4R/vaUTrEKaekfslBnkbLvE05B/zefBTaZDjwSmQ
2d5l+DqYSpj7vz6979BOSP/OWQ7tHNwqwDrMMnAbpllGzThf0kIqzF2RFKSDIMJP0x2Rso66YyWO
j9+2QtKUbINAIjouNgsMB2kULWJvPyLoleg7TxnIWNp0eMxnKyGjgA5bR3NY+DvDlwlkC7amTTdR
QG76lw+ShBaYKZ0ZBPTafytI+K5KMjVUpHVBZL94S2LbDB/wfYjY3sf6kXqAyP3Z8QzdHyfqVksu
KdPc4AC8z20jML/49qmYUpXy/xFcEubN3s7dESLPxDyzmNZAAGM7a1fq9+n1gmOJm2X1b52Lyak4
srdg/Q9iw+ykuuSee5xUxF2rsmSLdZzSMESJVyFF+HoCVMmtghQPUkQcbV7M8MybRERt7Gff1XL4
BvjANoDa3jz+qBJP3xjcHcEzRSH5eLA7ZaWq+B+6odwQh3EE+ixkMV3MgKZ8qwmCTxi34yickoja
78JveVmWLC+x/QlIY6CzN3H1oQskc/CkjX1olmbhskkIsEr6S9znbI6o7lXvN4hMoBstC4DJ8OCv
0KgPpz7viEOUy+BorJAYumWuF7pcYFXUITITF98gE3Bn00e76ojaAxgOZLzIBFvXYeuCEC6hs1mR
MO+RyKmhlS5GZpm36T6okD9VBmdBa1m1CH2O9vuiG1z75dAitnZohrOjJaMtoEsyLUzIK1mpdp1e
4mmT2Y8uQ9vPfyleMFAUGS8fcILsu+sa9lnsMrneI34PCf9u6V61UnQ/eyy160klNmrd1eF5IHL/
CO2RksBD6HftkGA73lzXWoyserijj1MulpMgHM6ZX5OIK+dvq7bm8hygSCBhy3ZtSftxb6cmmtcE
IkZGRc17mIa8yMJF0DBJ2jQMSAMsIpanLC4dpFaiGVPREMp4ODthbLCwr31LWxRexkr5oZIyowTJ
7gN4YBI09O+EGOUVWfuuFRxhVMZX1tipZdauSRhwwywyKfug7AZDTGyC5/y/7GqfDR+KR79Que8d
SCpgLW5h9yU3fLQEKiJYjnYxNLtBlqCrFulBL01Y0XXLV1D3vNs5q4hy0s9XNN3pnI8d2yy+D18g
9A3Ec9YV/eFi59CZk2UqaA3zVzUyZBDevsrO6VwlFNdcRcICaFh5kPF//5bvPfgZMMltDdC/87Xj
2W+hjjzvog2YYBzfHmFpSru/uLXzlG+Xx95sru8PF3E0mO8XyjcRr5UOT+ryAbEkq3Fd7t23xkZG
vLJuljnRzPFepbj77XNWyPg2PZjZETvRrpirsAYxbef7EfJCagbFNxuYiHoo6/8JTWiMQCL87qXu
t7TrQgR2udM5QZtTjlH2OV4t4ubH5RRavZweilaW12MilBXVU8S6tgCXbCOwRPVT31+zCG3PDtyK
wQUKidhS8xD6n1d46etFQjFT5yRNHSOvKymQ41nH2Os7Uh/UW4qqdcG3TC0bwaXqhhr5A5cHlxI+
QMsPCQyCc3ATImpCYV71Ug50ZJnn4aj/q3l3PBnoAKWzsNGjv20qmyguEPCqlE1QTieAQU/qyNdC
gW9AHNoMdcTqq/RDJqnqWJsf7E3velX3BTKPl0J7nc5HihPnNKTFbK9aXckAF1RfEqqzjeVsNm4q
a4Vv9Z7EDif5YYr7qNMovtJsUKSDG0D/9i6tx/y+ke8oPXEnLr3NmR8Vd5ICGQj+7tiddRBxiFyE
V6MxVj3CN+cfTeDz+9X9yINdtRw2tBwfA83mHN1/KRMkdzS98FCr3dWwb1+uNCUQ0+cJHAnTzfT2
QqhDy4ItTJjVq659qbuxN/nsUanJtwmslftJDjdCHaaTjrIrjh+S/iq1r0p2WvPf5DjPH4+wpZyl
aynZ1DQFhEko3gAPajYOvZ5sh1m2Xc2PlP2YzbI9c4ojhfIsJTUfJiWnx9yK+6RufxAzY0lbCJ/E
8S9VcYLNxAFj+LUHvxv+UXAJ0pOa83JHPgr7RWbCYtvWbPOB7Z1BYYt2A+Gb8xq9mng9N3751wkF
aptTk5AT1VFZmD5IHVa+jvPI2BTjdyl2/GxQ1Fn39tHIdu+v6yWtHLrVCpB0nahok/9xBlz4hhpZ
Kxa+EXryWXFUxVEc00OvtkVGbTeYTuxXqwiv27mSxZZcCpKWMKDtmyulNkKLw3/TU/+yy2C3Fgbm
cynB1M/1A/nQpGZHS7xQlK/nHqWvVesG4YRtXbK0eKXlHcGca9GSwRO8jZe7kracY6YPXRvPOGX7
Z/pl7XnAzfECEPxew2pA/gv81COpj9DBBAt26uZMxaEF7gcoBQZiONbTAYIVovY9rhHKqwugys0c
o9crppmPTzJbsVZxtGaw6TuflYRLqE/HQ+6FjtZFpExIPQhBvHEUehfc1Ou2m+ra+6ULbxroKJAj
Vit4/pln6KJ00PUyUtnzp3acVQsCeykp3/6WEcprNerA69KoRl9ET6L1YmDlOi3sbpnBITnzYMrc
5dvmpp/oEvZlzIdCREI32hj8W1TX8UHqcXjApMNWGOEGdYVubtBA61HOQo4+/MPL8cyrrtJV7yTc
lfghETGFiMuFNQu/eP2lGiHVuILRQ9dARWtWMatRKsckptJ5jwQE+zEIvQbqfrh0AjX5n9ZYil6H
3qGlgEGwWJG3s3nIzr77oMb9lLSSBsBBlCWRCZhRqOBSWBjwZAHEQKtj1o0kfRj8jaf+iCIlLHp5
r3HrStkTE0aFV8DRhMLz9QLDDxn1SaAtMpbb1dGrpTivQhua6YxI/RaMh7PPKLNfbO5EkR1BFpRF
7YoJuoEO9j7gNzHSaPgpF7lg3j/T1fh7nYJDpxGpBejZeTkCZ11bSMOqpwcJJHykj8+1PlubKlgI
bJftzpmzR6MDuYxFViDGQpdwqp90PEatbmmG6xkS+D8RmNTHXXnipUGVizEa2lEKaLL+4i45eG+c
y5Cgvp8QsB1swdv0+KGk0NlZVgDFbU4ZzMHrQUE5zXkL+XkRCrG64f0c1vaxFyUVvpgALgYT+v+j
VD/knE95qe+5DJCV42vgGFCuTYZvAD+lXMQSainWlN8/aQ4ifE4AHjsYtnACaua2vm5G+1X57VYs
XY359oOGbaETgL3MdxooC/1ZPnjYqXZr37V2JUlGZWQL5wYHphxWh5jfyH96lBuGp0Dmo3+DHtKD
I8oVHi56hpfs8HURP5OwGyQsK2DRZTW+49caEusSX+HBRMMJgov9ekopEj0MdmnHkzVeV3htWL5D
F6cJTOXkSFG9KqJoNo2+WuRm3t8JwupKVauNBsLY5rPlkQ636riL/VdiJA+qjngu9fXfaMJHnLQI
TDjZxV2ugiRAd8IMr2j52zMMQ+O7xb50yY+izwejgOmN2nbENmfv/bsOQQXqM07Zc9B1XgMX67Ne
i00sNNemFivyy4CyuxB6V9jgB881l78RgCCXc7ufJtOkfMSUX/MBxZUv7oX/OoDnIKjJAGcmlMmc
BbUfSSg6j61tW3MWUZdswUaEBswnkK1c3gYuCLtEs4CGbk27+BbuKzfPAxqiNN652yjQECTplgOQ
uOwIYHb98FejJDar/zBX1dpHIRHoTD7W13a4W1yMfj4kgqPwaJ7p187Mlw3VlMj/yEkfjKkHNpU2
evV0jFcFhJ2dGvrLqYRvkf6kvcag0KFepO02m93taI0laSBvKkpt/esfZCVB6LwSQg3pLgKR6Etr
RYc+l25hpYyBo3oAcbQRSQ3m5fmeBoiIGNsomqIzF4yheZ99u8a8JlhfXO9dBE6CX2QurODlYKDn
VlVBduBfRTIqRln4paTjY605ne8zHV9FgkHauXSHfkQp9vHdDOUyKgLUtbzxIWR8/SNX4AEGu8c0
dWK4c9bXm8fivxYATJc6FO8PrIpXkOqbipkKrib409xg4t4m3x69TePpeTWZ3fqFYbf4e9bEhRYq
DJLD+Sob5wK7sWBiduVt4nWkpMpicwIfZ7QEHG97XGfNb0ikS8NR/VA6y8Ge8Bl7oGexrozb9FsT
zc0h/GnCuHDvKLkVdIQvzBOQbjo09LRrAEIlqGoDmOUBIo6xkrFg7IvLuOnL6UUhVlOrg5ZZijp2
HXR2EYNjUqYhRkcEQQBIPdh7lscMyCfX3VMwHb30sQMpzKAdJCB8tWm2IHCjncTTyK4hSsln1XBo
pNC7XoiLC+wsh/ZOUm5lkl6fCm+FIzOGAryjjQ4+0h7foOoYak3Z8NolMWSrVheqSRuYpKk1ff2M
y/wbZW90cA5i9N7OUCVLzq0WiMkuYVx+a6O7b+u/TiVQILkAmJqc7TwkU1hODmcjHCJ6qsFoB8mt
TfZ3Fk9yz9RFlCkQcZgFlfJmMKNW3VPsiDBarJOvAlqWi34jdBWQUZHeQyLzpN7zFwWuOgPCiAAU
+IKn3lvcV4rl+0mHH3MO8s+SUsV+0QnOJB3axSsy/sa20QK2rHtBOURnAwEAkKfE3lms19B+mbqW
Yn2q87BQtqggtNDnIi0zXOYg4zx48VsG98Nogk848rppO7H2JVHNURpobIZ1apjLYLdYpYFOiFPc
fZz2IYfcWVpmZZcHcNMCd5dWaxNjQ92cI5iWNKmJLMC63Ul4RGhY4sYvCjWkrIVt2+qg/Q4F/6cU
oP+kbFX3aoMUla4j7T5f27XVvI8Z//N4pWLnpIAU/s0eYVlgGtet49Mp7z4OFE9nDTgOqQoR9one
ejXUuGp6yoE/fKSojzW+ye35Y2C1z+HlhmUXHSGEKZc3CMnsElVnF4qFD2GS8SuWR3UCe/+c6hGf
hkelPL8jLNFJWgeE+9EzjlddQ0RRa5nuyvdDAB9f67YJBJ8r81ieYvkLC5l4C57XapUlaEjxXTkr
I9wMXmps+SKNcZJzoYedhCGGK2N+gvbKzw2ATz3BfTGqoqmQ0EQ/WBWGMOrgEsXMkfkKJtGOm14d
7wtfqOkMwf0rkJ3mkqRhzQ3uCBwv+Z1QZvOltCFWNfEtHlwk8crc9+sryeEQwmL4pKER9RU0OZ2r
5jlOUaVl/DBI3ZdQMT9b+XAvK3OnPltA/e0CCZm0XZk+5VCZ7ELEi6lGY7zhTdomT1dj+ZhGeNOt
e3FcgoR36pd6XKNbqpITD63brqdtwc65jHC6p3DapP1x2/lW+korbGP2+s4AyHHutQRPBIKS7P0i
GQIGyY/Vz7d8k+ZTTu6waJefkvZCOoP5/qjG8d1ftA1AoVfaXUW6sSkLI35T+qUHoiAzrGGESZes
p7YY6r93IeasH6phRX2zKQaE1oJ+4CayuZ28qh9rSvrxWNnQJpxMCCcsJTX/CJ7ZPrCgYKRhiApm
JcTqY8oYjKdEnhkzqVaTxaQuAzKjzm22HVR5sQU/nIQCVRDM7Aevdh1j2UAGFF4CeYJU+WwDmbPE
UI05HazqCSMaJVhCubV85q3UUo37vsflMc/mv7ufPAdISVWdLN9wJ5jTYyJf4hTqdYFbc5Dlrj/j
okdr/5MW6envoamDJT9i1cdkmv38o6vaJJuD+l9s2TO8WzFrUCxAdWdjO+5wjBITf7N7Zs++Yjx6
D/Cdjbzcm9gx8CdcbqsIyAq3izJ6lG7eQ8LM5ayqyjt8nhbM8CL8r7enat9GQNMXC7zDppbkUqJ3
CTGmed1TjpYgjZSjGXTmxT5aOqoYiprBgVQ8ObvpYLcaoJvNkvOFILW8HL1E3WDfMiTCOB+giyFt
/9XAYTUefCrEru9DNYP98L66YmRudfnQnMI5plx/x7uD4qhhKOZ4W6bM8ttxyxUrxnVoGcl12Uht
59RV583s384ZiFbwGWE42LZAHNUCuzya5WK5t+/JIdnQpkSVupCnoJ5Gqjer5VOBVQWWw7+oxX2P
OAoWad+4e7oFAWumvZlrMh00GV5yj18F46KCF7JPchPgz9/UMVJDx8sLGEuxK+24UQWuLvJ6aIFn
M3QGcGOdxEgTmLKI3sYYdY2EfLd32+mICEX0GcLW8c3HlNcOOmbTuyd2N+eH6YaHP/b+9KU/WoSd
/yBdsQSEi3eO+BXUEwKb2D31ab5rLRnYk1c5Y0RiAG29cbGuybAZNj9c2zSZg1avtwabubWacjg5
1DuYRgfb1zd4fLfZCFOOrF59yz9/75lXTMvHa0mXGeSEL8TT162bKxRThrBFqwGgm6WW+XUCLWQo
FGEtH4jkz/ZhxVcjs1g+evadFPJK32NZJO14+yhmqSlwisSelexYsSN5T98OpTskEP05kuhscg2i
WF/yiRnk2XJGo5Q+X+tFvpkkTNsCDH54CAaV9T+tYzvc4STCt3UzMYdQ8tS6XD/gxXZeiTMfhRKk
68ecwOFb1mL0cK0WBUJD4Oq2AMgGRDest9Y3Y6S5ao2+hIyjc7T+3/B4U8oMcaM5Gsm34lGnXKqS
aG/vI5xMEtLZVeNVfXWztL5CtuybWV7VvdohKG177lLD9QVBkKhbfP22lykfV//PrUhpAn1apcbS
1hlLohPQdvraU+HZwq7cn1O3eyqDZhCpRxLGQubeDbV9G/guVxm8+W8B2hsCb2El1oifDQ+DSkKJ
exjEYSgKnSO400ukxBpnKtC62lCkalCEbRNJ8t3OpLI7G+kFsQK66mRO8VJqhC0Zi6jU4TlfoUqN
gzLs6MsjGQCqPoO/2IT/3HputWfPjXfFEp5oBOxCpuIxBJ4Q9Xkz2cYJgTqjfpLefssp5g4SZzSq
dV0qpHa0uiOLHEXQMCR6DAxek7G1pt1fOaDJ+mjRnjDC5wZky5T0aijCMboULYEz+Dyo9LQcXRwa
BGMRpcDkwV8yK6a9coyx/ukGAjOk8K7KFh758krqenpNNHuQ6uZMTMSUGkdZPg64cU45a9LdZc0y
f6bLhc6o9zLjH8j7jAlMmrw/raUciHAKpBkPkSZOkWmPZgE73Rlf2sX4rFYwbmdht8aP75hn2422
UM+IKTHMoIuzRlAumytbX/JfEbk/wTfnnsgEoT5MewaYPoQD4k4N2qLs7J83iejaGvHzBYupAPnj
yC08o1BlgNfxDglFSrIu7qhD3rGs8Z8o68yCuq5tUfYTsnNbdr8YLkmVJ3WbVna5G39K7pXn4NlQ
TC1M/9SGQd0/ROxVT1BgydF5DNhB4g1aemFiAmON2ksA2qA0SABx1+NeDCD+UExJz4KeO9iYgey8
4Y8ho2eICDgMpW7LWZ4rFyIbnqOjAokOs4qBh3BqyTOAgq4N4FQjOU5loA4BsqIN/6kmxIiXCb38
BJfoHti8vuqaJAxICX9ZeQ2r97xmZK1vP/+9Us6hvhDKL7e3BhJJyqKwWB8ubpJXZUjKr9kDnoi7
OYJcdXHe7SrwRjkR5MCfVHea9/5kK+UCPOYlwJf+Py4xEe9SALwE7LU7cqTGCcL6O8JtHuLOjBgV
7w+65cx4CgK7rd71p+zFHQ8qwoIt/J4YnsNlN2FBbRgbNgC8rW738WwQw95Ps0+Bnou0e2kVc2cl
+r/u0QaxQcWc3+oK4IRHwANlOIC/x9Okomo5u6IMw5pYd+9iDLny4ZUM2unrjQlNkszuppGrsdYA
HY8vIHjJ/itEvqrmkUkHqpZHfqvfa86uO8dtN/zgRDmVoEBIpPjuJxJSZc0GXzmJbFp+zc/v38ci
tjVoqQia59xc6BXZ70Bf3ntSMaUHoZx2UpI0UX8LercGCA/KHOlrxVsf5vnIWQdI/czBt3V8keA2
EXzpXK/AjHviieQO01LYoXUqC5UirUu+8tg3GxkJb6npgsO5clTYspffPP48k4am8CDC7EnKIagF
1MTKx++F0BPnHqx+eoHpDJYTHxcUBidgpdt+91kKOGkq+ebMkXKcZ5KVfjcdidb/U5fCUsF2k0cr
IuuzMVD/9urZoeM0Lyn//PbPy7tUgbqP/MUICfW1UwlKfC29cWPl5Ad04thyr55rls1VLW+L8Pns
USgU8YRQ85OedlYE0f8qLASwZZXAWw1kmD/MFXeSxCp6Gff4bivoaH0P1SpbSn3k3eUjYB5t28BU
OmwYuVo0+2U2eXEFy7zpIr2MOYLFsWiJHgFr9D+QK8ilPUueqI9ENoP5GcO5aeI9oxvMpoMkD8hv
wp4IrRNnZMEANbdWekftDQQ3623eebou3Diyh+U/gL6yKYXz0Du6atx7NbnvSF3QtPCNlyPn10ZO
jnvqd3Epz91qpMbZzg6cSiW/araIkYykbCPcCY5AGvNEhxaZp+/ihJ6iS5xypqVwMNoStl4uHWbj
uvimioUhkuRdwPRX8utMXIOAX5wiYWKfjLMFsVJGul0IITM9vbc2jAOUikNnlkdurDmevgDXES0E
Oey2AFKxRFpVjVCohYvA8IqhrcKNGJvwIubxX11yCCyHeERcNYLRq/sQp7mxjHZXvQhxyTuI9W1x
oqhFM27Tuszog6fuaRxWkDmPzdfHHAL8lUj/vTsbSJMXwDgGOaB+QUqi79fqmEuh6EEZKQ1tM602
uzP7eRxp6/JE6pMV9j0gMKrCIFkDl5maQcYf3SIcBlxF0Q97+eQ7byYRH5u+rQoQ5rZML0ov46jB
y24e02h/qJ/gG4QIU1sIZpyDtaH/7FdEEY9DMA68Fho2OfCEuld+QSa274jIoG1YHa1mvCqZyObI
xfp8fwTQ1pRo1FZpqLqlH/ML5KIZ+ZNjsm/22HTUBfz2Fb3jZWS5aXYiG4uaDD4CDZlPcRf11zCp
vGAdM7M38Z3mm2nxTPJYITsStkvaJRwVHiAiIT7eKw/HfIwchV+qAB/22FwcgeFYAQL/jeMvt19G
BA9SXAsdZUFjChmTm1rRmHBgy2G8y8bNzhe8Ihs0AtrTg8PjklLlybJlxfsmJRj7zVNbeZXSnGje
XaZlJ4m424t/hUxi1JandmMQxlbmzpUVIWVLcJ7w2qDv6YPJ8rnC08Q+Bjrl0awAvrVtVdEDtobN
sqFYru/4tAMsP+jVcj0RT4ms6eNG1k2EUS+gjGitA56cz1/2gwHl4rG+IDgs8WNk7dE1yKV93z45
9X4G88Fx7Q+VfmCcyzJqZykas5J3odGpczDeX+Q3nrs9tHivMbPTlDatdGkjZjzjZV5JWgxcKXJ0
QPVA1GFyls/+kRm/4a8ONTMfFksrcz9UgOOzf7RKHBBShpXajeAOTZcWM0avvsqadWmEjBUDQn+w
eyTrfqhxVAKU1gsuxc1hronrOIh5GoZT43Ge5cwxx124LnBa4Ae2fiFsjBwZ4Y85GZQPMTvuWPb+
x3eFQFxH1CYWcfhuPAD3jfdG7hrcUIwRdAINjn2N2vRIxIp8unjeL5qghc4i/260KjSoma4abOKZ
ZXg+litW3WNIy8r5uBZZRkkMUSA9H8M1lDMMbV3qEkrFzJu1NIYS5SmqezXlw78ZF6vdhvP/Ozs1
KcqkPE5aPncsSSxWic0Vu6puhtL4U0VyhKGjSjgZMV8V+qI+Q/kKmHjHRjcaFbUy6GKrF91CLQqh
VWEhX1j76OtJSczLka3s2GHuPjQZdP692Wk3rTVrnXBCAPDRHcOn8A8gR6W1VRdBUvQJuv6DTQea
x7e1sfPZ9CZldYr4NP+gwMpjeyQVW2AP1IyPZNsPElF2IN1vChbjJvdJ2WxXOTEsR/sIfn7e+EHV
pu91GCzfsfGLeRbjVkrShr+YKGbcELKlx1Fwj+u9/xnbyPEuMpPahCFb0ATFxxytReKPuvT+QmEL
0iqpBMFGSsMVEBR+QReWqJ+cYt5ddsVaf+dIUsr7Zj19EI0A/2ISyPzueQUqOolW7q/brCGEYfrg
YZVReqhpetO16FcW8Oti0L6whcxVanr6EK5vzcIw/TM+FoIASHpam2FW01OuzPmF69OO6m9pXqZV
yZOAcMEeRVVm/YsaleJSw6K9klKj1xeKqmFFD5MEB8nVkL2+YLYJMg3OeXHzm0tJLyOt2wRNGpjw
Fsa8Z6YIwz/LRtWwx29fSl9kKN3tIbR0aS4dEDCa2sVVmkUVemTTrw0df5PNO+0Pi91fw3/xA3eA
pOdyOlQdoavI1oxBQDK7t3EV9vFIVIh1KlAIyqyHJ1k1YtaHS8Xx1XhhzbnZt6YM3dGyuAH4II7p
kxQo496MZteEcnatV4M9T4M+fZtxRxRPav2j+5pJHVdhX+0wD4fwIrNfAPTHXZIbXesZvY5viD3L
nqSNh9CgoS1UN4HLog4iPByQ9eO6SL3A3BVdLPb6JodvkhbQgLPkdv9pb6AKAsUHrr4j3FBCajyo
U5L+n8jZ7WqRs+noVyEgy0MvHpXiX7vVvmI/9s37/vytgeV03jYPtzWU5TRc3RIcmAInLVK1m98g
+XoKgaOVa4x/IqljGlun3eBVmAEgq5JspkvWzlkzGycDwgJr3lY7XBD7pah0czj/yNqrgsRIle3e
8SQsK5TJ5k6msE0Zbg9fyUSx8jP5xIdgVah0vlenkbjxcbiHxbAPMiuwGn0I+WmEAO2EqavLg1Ki
cY552I9C7eLH2H+MrieUMeVSKtg4605Jm9CFdiSjkeGcKQEPt3NO3aFNEJYL5341yQqwchAkdPzN
cdN7xqY9pgaChu8R8ggZmXKIW+JjO3JWCaCDQeZlIWG3CZLbVyKGEzG0glQj2UwYAYQQQ4CpqW6j
dTqtNmQ3ECu+/s/sFIguNXA196dL6Le1TDzfTBILwy9tKozseaLx1G9DU5cpatMcx+5SgthgJQWO
RJvoezWyj/qB5LXUKbbx+DSBBZ4R+yqV2GPULSzpfUXalQuh03l3G936uc1sBQSVAJz5ZcsJVGpK
Xw/Y0v66NTQ1xfEnWeE0vZK8xQFAB828KqHi0AOAJ77FoqowDc+I6ZHeQKel2kRAtbbYJXK1vfw7
E2PYbD/WVaMS4o9yl+8CWl+QVSUAZZMNAm9tSj3ZcV5snIfFXxGQN5oND7sCNXCiYvWWX/z5Qowj
IvTlGMBHTap8YV5jIxcaQt3B/8npCTHo8xjnTBMTjo4C0sIwU0v4hK9niO/7HBz3Z1vWNYrHuWmo
in3sofgbnHe5WFndperEH8kWHCnR0nEqqJwCp8039mnnqFVFz5leajZXXSDNtrjuRdv4iOZqVB1w
243a3RlUi08d6b5tYpdWhaEnkJCd7kfJQovlO2ZWzYl2uaMTBJh/i5fICw6kB8e3bjozwAZaFMqj
3FsC1+H85OYm2GwvYgqUB7sr9bL5xAyqFGyKkzVfqf84VJJTLfPxkwqRRATqlryaibjfcMbPCPiK
8079CNKivItTMfkJLv+rbbi9PmPljPRrTYvTJVSgRzeWVbHItTHSPN/4vKCQkcgaqChQP/kyopdy
6OXlpghAO0gUbLLK+QtuYppayrEBC9rwN/CyswnyAqsme8dpP8BjlsQFxZm5XlxZ+5g6UPXKvBBH
7Q2QnEe3PzTkaKyPB/TfLHuzPE8CIxCBwT/opt6xvF2gH5k+R6igWZkRnpyVMorrUiU2iAiCDckT
wyrZKr2k2Ih4nDoNyUz0lXAU2qWUFZtqHSOmSOZwNZ9AkZmos6eq5Fq/7XwP+96rqZh6HcybTtAq
9O+8MejUH1jQiX7XK4vH4JpmtzkvzNr7Eeznxu+Zkxg/W34CBCO2f3ZVaRvm4PvOoP/EXxlUZWYT
KQWP44STFhmHXj1tKAY+4fJNq2HtYOT3i0a4ImeA1LajVljefo6uUBjhdEosY2Ot+kMjP4xl1OtP
Nw4kPwpxStO+0+BaXsyDWowl4J8c6TUKPVkE9o4uZuLp5uxnI2sNcYuE8sR8g0FeaD4T7aVybQX8
bfvpCJNWTHN0Tr9foHcMb5WN+oSvXJQYIy3Gm3+xsv+yyJ6eTeAXinfNaBXNqJDZ1T/UXq69qjiI
4xk6OH8fmBien97Kx1IAUVPjp3cfW9rjVs7eqchpIGmMNOrE7NOORmLyku3vVMgP0rZ/gRjoArq3
iMNAo42Jd7PZNKXtB9PFm4kCMFusUWan+DyrPj+/yXDbL+FktHK2Y5LG9gRsWHg0UA6QQrk681wh
ZMLs/49nzKMMCOJlsMeOrkG6ysqgLUnVKGZq65P6VnqLsnYCIGCV5AtqOdasGm+aJibLxFhs7v0F
Toagffe5jkYy1yuwZKn43Zdaakkpe7RX0I3O+qRyYwcILez+WC0LglH2vq7j8JnDvKdMSxRUfhwK
3hJJGSUu6mNTBMPh+5m4mLejDVIh9LxZOgWDxvV2Zx6/C5s3XyPLC7rkn5NrPd1k5UFzPcOBPmJl
lIZ/2hX9bAjoLG6pXfYRHFXOnYwL5HVts8S3ZG8tPYWl0l9o2CzoTtl62EiNNJpaDkEC79v8IsPt
FYxbAffgQZdqQGmA+SE6A+xc7RwhTclbmDtGn58eXR5Xaw+w3DKQ79UHQlWGKLgG87lytM/No/kr
G6+n5iyaetFAdaicKdiYEMy6V733Bz/2jgKGFO317hFl/KvHa9IZme4D0oO9w4p0mWP/aHBMOSlG
pAtygO7PhtMoHGpJigumGxgQd1lA9UNlCS5Xp6Un7HM2xhOq5idTo5vXVAHR83u3F7/1/NivOowd
ZoqiaJZab6YXsuZU+SA0bUDP7X5913Zk+h2LElxApxjMpmEZwnzicvI2WkB14JiXfqjjlthWBmT0
U+QZY5vTK/WhVZos28pCZCMFmXNIPCMQ69Z9ifExA6BXclGZhVtsOYXb18lTORrercS4rGLF9/cd
prTz3VJW/oUdnyxC1B22LideZ9S+GgHCfiOw5xc9yymRjCn6JjAYLuCw72xmVp14AeP2tp1vc3w1
pLsZzDymXTKMZcThstycEtZSxWY+duiKuNSpoWDywgeH2KsxtaIRyy/AnQqeMFPRQkRd+rcjdN05
oQszQhDGENoAZgxY3som7oFW1/o42je0fz+IxD0rT4yS1A6iTWGyFJJrIfj0OyiZnIZU9Hzijylv
G/FJSwpW3CdC0zQoPm8MYT//n9bSxNZ7KZK+yXep7g/g+pJfYi4mtQxTK7MleYwiqBrSxlp4LsHW
piHChJG7GBXVI5oCzi8twUwRUkXBr3GeeO5Ri1LuhTE341eQlq8XaW61nUsX6oHBpBOy2Wv+4jCc
8juHdwucCxe8QWml7QuubS0qebjlV4k7HuMdATBVbw7kkIJx2D14B7XeDeUqzHig6mqlMM+P6rDj
+QlMSFoAUwzTVeXzw2eyvEoMybFAUR9PKKAtWkumQXcemf56VA4GQXDXa3j/rBOhztT8JUMo0cJH
2esdVSxHa74zLipJeCZrUtPVXhTB++v3Rvf8g0eq/H9PaM/okA6DLwCBGw2War1nsjJRMtxEW5Sr
EW5KPEsFv0xgMn072LBArp/3Ujy7FOr662HfF3ijDV6n/LSh5A9LH4So9XcvLLvS9wLhxsfbGbvW
NeqSyxu+TSxWEGe9FhOejELwEb9GseeGZ165Lm50VcRAI0mjHljqh20VELEQS+X//oRFk4hSaBPn
fWnj3uyuoGbI0RAbtDhRj5skSL06c0/xZ++WVsNug0pvFNtwoP5ASmAei0pOhGnKQGImPSBaZ2gt
4RCjjG7j4AdXx9cu+vozzruvQcvALtB4j/60Ue5tRMi+k2iu6T2A/MG+0MIKd24ctiAvtFtEmhZY
uxoU8k9vsw0frHKCF695g6b445qufAs+CA+scu3+H3ubwuWKgtZgk3y+hQBZCJYcIIIcbaJbU/XW
fQbHN6nf9oiqXX0pW2EQXoQce/1pzU7c89Ofirfx7xo5mNw0LegxgjhVsl30STmgDICPa87qsO6N
zVrME7nLDrR7YOr5zFXr6TKX503ZdKVlx/F0Fviavpkn+Q4BHcJ6XCVBX8ZEyzpMEe+CZ7yPCVV1
TtR7jkxzXzaeU6v+sOz1D5r+2pse297/cX9wDqlBP6N5BGV0qATQEpm+4vb9xNTfEttpGsRqRh2P
MTdoWe7D7DJFS41TtK2vZMs5OCzzv5rGHx0gZ++ztFoHEMKlE7KjX9qJDvlYUncLEvfvRODgKLih
f7i+5tKQnSyksTFnxH1IX1UsNpoT1tP0omewbKS5GLWGhP+RrRclG2vVhgATY6orn3+aHUKOxXy0
Q+kHbZOraQoPUtlRZWcGnkCr8shiCa/9MPb097dgWveqJA0TihwS9qwbHuu2U0Ihr0H99p7z9FiI
LR8Z4tI1PixL+C3nq+xjlTM6muIkyE2QkE9TLJ3YoAFwzT2kuUXOexJ5lqhG2OennMLLYCua45aG
JuRaFtX5ej2/xC/waKjEJLOS1Ys1DFQG953XF1P/K/UmadIDREPOug26w8TlTS1RCzoIwH4CpJHt
P2NDrtW1fkrRz2FKXP87LFVTMbLNtcz61j9bNdugwEcF9HpzAr0LCg1wfH/e0AlnNyqpOHJMxh2E
2UXe5XgsLXzzv31DUZq8rZ6Tezwo+4uHa3kyGw0On6Q5vAM0NjxW0uk0FK2QfIMSW+gESEVPApKq
i7JAx8wmqBJ3zTLksv5NJc4xTwiQ2Ar4Nyuw6YpFexvaG98+RZZZhzDBb+/gvTUc4MSVlU+ReBGt
P1KFyVVrKyD1hTHP5MCQaVD68kAPAgpIieq0L0n4VzmQNIIuQxkCmTpaENmXYSlVhToXM04ahW3E
WvQa8o51wt2VQCz9tm3DqDdr+3/rlW7+U/sREO1l3PChHJP7Pb5idmvbkS1FzvcC6wEt1+r93/Jq
SXZeeVOC03WbCpV7U3fOGia/e5Z15tX1r1+9RGbhymyvQmRuFWwPUqIXD6CTmvJwCMEOoh80mZ6C
XT8zj2cQtDj8U3lN4niZFnxahM3cC85Z2YNVj4JN7aWIpuDSDoTHz2VvTkZB5lQGrFip2Cgik9j5
xQkcEj2/pf8PbW5556JyzRETPiRuNqemgh8wEdb77ldYDGiQIPbuSOgJDbr6XBDAm7RBdZUztZVd
bHDWqfTJ00Rw83FV4Qp9uAtbcl1e1lUcV7roFLJsL6+ZKzy5O86p3lznNA1dISi03Lb6kzL8vHni
qFoENrDeIc0dY5ptaVgmFn57TKlesnltQ3Q/h8pWe6aDKjTtVzucLaelFZIS181qXgGQnl/fyeQ9
VOqQ8X2cdLTvbOvdxp8/8mw1MFkVwIWzAQwaMnkuRTDuM/7OJ72VvAC4lRvXNx1ingM2Ky7H90Ov
ZpEXCHExdzGQLghrShpeLXi14QrFBGY8LRcEAvEc4kDjgYT3uyPxG8n4Nnm1FheH8Jfe9XZprH26
tE21+OOlkYjELJdhmE16EwSPhwE/NTLdiIu/la6O/1tXjye2kD0SGrQWRxTFhaAUxsN0535NVxTC
S9/ajrUlze3klIhVnKbYNCbmCMZRAQ4eIGPROvRl20Vjs63fOVIoWh7TANc1+Mjjiuum3XHUcQzc
fbRGysSAh0WInvuK1mV/qdFuaBVOGv2KCuIFRKvEHXwjlbDOt04nuICyL3kgy4QOlpLwPYE8EbRk
sEMaB9vuhdUDD78lps2Dc2p9FvT5HQz1eFp9wxk3qV1n1Jr7Dg7/tFMCBsRjrv5s9vYjas5YNx+Y
G5QWR0SCAfUnLF9Qkiz6KU5J1RUqwFK/8ouhfihtq2d3SNl0D7TD/en2Zk7xR8wlan/J8DEA43X3
/ULLpFmzc4RPhMimMk9OeGi5arS0HflfNSCUX0gj5xHo4TFoh9C+rn3EgMfRx3qGULG/HN+duK2A
hZQW57sorodwAZKlFGeN4QEXlYau/yx8k4U56qu5W9Uy2J9NYRz+SAuSML1aEa5Jq7ZomlOhW+iq
28e9XbJac6cik4eUNEnQ+jBiX8oGoBWofQ2fVDtABstZhRPh+X0PHz12L4iC1b9c3NZuKc7dKPP5
PQpDbKPmhFyKTlNtPbk7yVvJ2wy+Jb8oNPgJwA3/PFYdc7PZ4OABstlh8F1p3nccLD3JUwVCF5kX
pbYOjQA/7VConvtg0wClhVFNnxo4VwMLpPWU1l0cAl9cxYbIMxnMFPEgFzHw5RjAnCNKQo1QWyMw
/irM0FB243GAaq+eqrfOtyMkn/52d9jz8yTVcAB/8OmLefmxDEQ+WgcVqFbiPixNzFxqpxNtBJrm
eHXvtim7kqH0inlNOTe5DO3PlaACIGkS1HTuLeDci8BiehkJrJu8ZkPv9XVVFyLhpXtDCwQcYHQd
VEMHk3ClktaeIyYF1fMGslrqWhtR5Lc1R8D5fnEhwf6VuO7pcmtc53TtrSzNvMfm5UOHYIUKHDPm
4UJuExl2UjPIOyUIMyh0QyKnHGfK9iL2p5eCXIYf7bfsyB3lT5CxuipUN3+yx5tpU8j1i/m5/VLZ
5zCk5IaqxKrOcPn5wbmkKErPYKlWTvKvpULpwK+ijrHszrPYqzFOzPBkfrE4U76QRl3aPhk3dljj
XVJNzUtK91lYWb5+7XQdIOUuxP+5XR7AfMXU5xdT+R5D0UGCdJM9n+7Eu/i0OY0JEaLMYuww1AHF
46woJXQmfs33ICZdFeXHMD+fmBWHcKojVNfaqQHrq5G0qp7tPSlwGtZ5bwxbD0p/V+xQVCUqm5eu
nkTdFxNEvQovMbT/lxA5g30qp4uvVzIKARVhQHBU9vEu09qBim+lIKmHRlZ9MnonLkq//Tacs6KU
pnaXP80BinYW2Cip7uTYV4eonlHTx4F61fwJJEN7fGwqCDnFeE1SQ0dcAtIypcWWg3QiejQ96wMm
zkN1weS6Pb82s4wJAyNpahIFg7xBY/5HJKNtSsgFE6MEiivaWDeboar5G3dydvJv3qByuqBW4YGS
7lju/zFePrszBec6jQB+LeSvIeTb+4rnZi7VlHZQyJiL4xVpJ98IpIiKd/9I9rnWuFh4319MXHQV
m4jDU0U82F81VtrzVWXHzTtRXrAnbvHAD2nzQAyBUnRuuQxmWIAREaYEz2Li7+PGNw4TuM4VyDSk
2bcMrdnr3dEWEG9+BoAbHELhDEkRU99kb2AUOefCWr3+o682gkEmhrsVX8f9Tib7MVyK59xDscd5
ZPla4fW6a/f/TjawsB4ze9KNPWWj8V6oN4ve0998tivZqQjgbKfg9KlCdAQkRSz5KLKUXKkFi6NX
9yqCxCJWH+BS/2HnqaeBRuvjpADrtT1LRGKfhFxef+LZAl+73uIesf7H6lHq8FbNdCdp6PyLVdlN
X24zYed0hZYKn8cQ67id8Ce87QUSlix07mkuj4dXnOige/UzOJMwOYRCdMoTsgJ5B7RDKz/eZKB8
PjRFQblIKzsxn3kCOmMOBhGJJPAygDLG7hLotPof5dEx1u7BfOht/aCTbrI6vWa24h2IgZOlewz9
bgVnMZfeOEXxY5eVwchRkz5NJZqlatc0RQO0H1gj+bvPlLEZHAAArSyU5lBHWmNFXQw6wjtjAR/E
ETzv3U+tM1261/MsxmwF0RSyGKWzCZ7nFGaZEj8o4j7d1RiN0lKXYdEgttA8JJiIjK3UwdsggejA
fjpCBfOQnCP4LItnThqYuSCVHX/Vxutgs3942yoVdFnFEubu7l74WY/wTAaakfCGvKyeQ1HpchV4
C99E92b8PAt8mvFyURBBgv32E5apMEth9BjDl2XmCyfp84KN0Zpj2e9vDJRgH3xvVD8oDW8DVbbP
+Q/DS3TOZ1FWXPJRS5WgXyXBgPYiCGbP/vOG0cnlPDbPdwjy3h+LRd7dVGgoY19D06EO0Vm2rFil
bCqWROvy2325oodWtiJICEEHoObY+aqYA65HBi3GyKhW50GyBnUWNm9tFgFkkY4GumgzhSznTot2
7bJj085whmVbbbX/hKuSj6Kfq/6q6Rp8G5ilOllXVY9L+t54F5wKotPB+lmz8mtRYDH+NY5g2n84
3imkNtnrlRegi6i+nfhYJIG5tqrHTLtronmnroJYhXmRsYDmYSTm9wv/n01Z//ytDsqAPbibXV+9
sUy+WhZp3Clxlu/qxaicCcwBnh8CyLO/V0OH7AjPiT+H7w3dk8HrO59qRunQOZ34E4IT9uQinHWY
kbh+cgQF6HdLG+dsi+tE7injeAeGLOocN23LSxSdGxCa/mabPGL+9CjNisTjnkLAUAJg6d3xe2Kc
IB/EmX51134E7WXSXgZ3PQcLILZ25jEOMMloxZqonw7MfDBOCYI9EfVzo6PvSbeoZEMHHBlOr1u6
mgzVzG2vNd5QOuE+8G6vaH7eSgNgkBgRxesEYuCS2fsszxOuR03eqWPuBdTbwxzwgV5zafAxW1p5
t2q+VEkEbbQIUG3Spg+FFw/hZhNWpjwcTrJvoEDuKmd2bj2cxqm4BkEIdqAmhTCWxqvwDQsPXCRK
IFwZ5tRPgG0mSHPACDqZ/G7tTUSdQdTCX4YK3DzNdPGIvc1sUvxgZLcrjCobC9o0G1W4fkyPgmav
gCzVTt7yLBYnop5Mxmxj8Bp85hesqVuu51Xkd57FYx3IIOJcjMc8376pBLWz9PjoW/s5x8fo9n19
N7yr8a5D57y68ThKGuiucuy3TQF0AGXNmQ1Mn0E6Tv9ez+hP9iKozgGbDvUTqrP0qSomAQ862ZuF
lFqMogDGJRyDWfTaUB5JLRP1Y907JzcTtEEJQAgNNO+aEj02AZsavavFv/AOHhGAxUMuygAJNXLJ
u7xcQHThYvcRGUVPnmEIwirsnlbmBv2WMWKRMe64qF07b8A6zinLZteGAZUjZdoHB3G9NAgShie/
9Sl4saIqHYLiBhjHtHbEauohumx3UEUbC8iQnD+hAYqX/04sBujFGbNefSSCNLNd5WZQe3qr2ZVc
O7tGFdAun2qz9Dda6aZIbxa9bCQ0/vPu2wh9NvTRV44BEolxUJHwGThszyZLskwN/7ws2T/Qzc4p
K5OGmsUX4byM56rqkUhPRi2wh5hUmf26CnIg52POo/j5O8OWgUkg3T2YEkEjZ+oXdC+gqS21MVYk
ZAJ/gV8WNokSRxb6/i//fKHN3J1nMMLhWOLtug6KbmYBX0bWy7S3geaKVBT23YehX0Sn602E/ThY
fRbDsa4IkqBUU0L7EycLON31dTFRLdrJS0rIYgBPCG+2jvm5gzzeaeQbZhptoA6dzvri53daRgc+
DsjonwHdDJRwRg7JZlrreVnaFQ8tfeTKFv0DHsEwerm6uKUI+xICA/B+ykFew5Z9ApnmWTv04ePv
Ep7a9CTdKXsbDrRRDIJfbIuOqvWG35uEhr6KpeXe/oLyJ4OGATQlHlitGkhaPhZBWeAoFOUby9aj
3zvp4un0AIJ9gUWPjwWId9gpmRDnlZlj33pRNTsioIJCN+MW4/K7/U/Z+KKHpzYavUCA41qFPWde
YzcGqcI42W7Qmqv4v08xlP8l8iiQCdgpKp3ITQ9Lc8YG5DhOyY+m/9dKsf6NGapjqtQgrFGRh8vT
CsnOfqBU5/cSrRsn2yl5gTVYhR2oKuRvVBmUPb9h1Yg5X+Y8RenmqqJw8EzatIA933IB2UrPqmut
V7qg2WNXQXSpUHI5j2FbH3IMSZkIOZDpSiJtPbiPYFe/7IPEamsHa7Dcb/xeBUBi8/QGnTDguw5C
fGy/VfZZmrJ1mlYiDGGLdz0jpdm6yBNmme8ensWOcbMJZa5+CdSry6xxxJHxqk5GS1JMhKAV3hT6
ISaonJT96HhpLYVGU6dNs81Z98tQwxM3txC7Ug8R8uRpW2nVqH2nfx42Gx5gp2nMvw/rmxOJTxfa
Q5iXxfW0fbqQ6daBBdgzZA9MUz8H24lm+TgaCp01v+15S7ermfVumiqEunLCkW5cAt0UIoTwnuRu
Vft/o4sDTdqGJFOiWeli/ltRHEMp/cFqATRZjnS4su46fK0zeu5CEjhavFwQH4GgkOi5mea92+98
7eGPwk7lciAmCdE3FkKpVGn3UNFqXXOW3XJS1pBM9vqU6zfrDaX1ZUOpci0QcWe6+AB0k9VpQXla
F5voTnjB27RrjA48woHeSv+flHKFvjMdGtm4crXz11XTZCcEn+oDGKOge8TlIggQNmKCMEiYidF4
MizKiVW634Og6syoX65Nk3FGGf7nfSpIwlGAiOVKTOJ1I1FSURHIdhwjPfMl1MjZ42w4fcO6wawZ
TJIz9/iOImytahJgPCeA/Ir5pmPmBPTo3U6CJU16ZPw6XSAXD+ZzEP23MnPLOOIldQyAcIEz4Elj
LK91nkzrRJSlYSgmaOnIqbY+CoxoIWrgDXoyy2oAgUlmycO0bOPEo4q0UX03OKJuFKNIDGDhRxvz
ORkNBzkQ2IzfwVp5shxBJXyTvF+jyoBKJMt23UpafGeUG+kiEqxDTEpbyyJDZIOFABk8O0oCksyy
alPrvKzRXcrSy8k/KTjbbWEAM4lMMbk3bxivpib6H/2L2L8QdLc2eFjLsFZKPolJkPHZ9PwoAPRN
O2nxIUkIFOnoDTt9DagktiqpwUZxxb4tbn+2Olmem1a2O5KeEl/2kKnEik3L0A96q3skitttGZW+
p6o33HpB6QTVaFPDZmZwPlPn3FDiA/2DGTpHNUENjWmoxkQvtsTpw3VXCEiqu2Z/mhdS3FSAtpaV
kFjpMvlSF3qTBmshhv8b1Ergiup5/F8Mj/nAn0ti/K1/FH+6hTyXFIlmpbNn4lbfZ+3m2cBKuCJg
vGx9+vHlAxvTMLf9XZAnrIcTiaqYxltu1lQ072NLiP4jGPR/Kh86vv2/YrhV9h4wx39LsZN2a2AE
AE8E7vMS5PFDpIojoyHx3wcKjbY2h+t7Z5iTlDub7ckqm8tGTfWfE6iYBoYUlUYPTmtUlONOPGos
7qWh7zcEhwRPkMfc2R4X70bPsKSsdXiJY4Th3cWFUV97d9km61xmSI51e+oDjFahz+bUS6Tf8o/C
T9pweOQqGSWXkBtFkFWer7DiDqjja/MJr5yD9DiH7GvgOqAd8aVJ0Rmn2nOgTy40kvRROhfowCm1
CkyTRzaEeDoVQBnxcGbMeJsSlI1Je8XIM3M7OOSL5NS+g2u9BwJWZLTKqiW0+mKoX8vK2oOQRwuF
ajAbGAIfJkUDGW9KbZff1t6XBL7c8hm0asgKfmiVW94iDV8elMDosTAZdE8PsY3/YGM1y8iykFo6
ay2sSTgyq2Fp5ZKKnFms4YOb7vuNwmG3KnfHKqliMKulj54JfhV5dOOH9WUaWTeIPEU5fxzNhjeA
KUnrYW0LadhxZ+5C1eVt8kYF0NfBDdVVHHnflXQ6rtCu9uhOdv0qzVpzCuR/dj+ZaSoSWRRy5zL5
RXqn7yZXXQVj7i8JIh+0e7Bv+eZ3wkI+u6s3vdZou2m0m+yYLiMgNcxppGBJd5P8K17xXzMmiQpj
1i+lfhSEXETmp3FmOb1GvN7xh78R1SMwm+ILSB6G18rsEr1xt8O/5eTZxBE/YvFTHV/uikNwGZdB
oLnkM/nVtRerDNv5+0tEskR3RspqFYJwgvPbwndZYiqrBOvA66uwJvpmbjxxkYPsOPLyzaFzSHjQ
nw7B3IoP1Qikbo47bR4tBuLT1sZVRjS74PxnwjGgzUEuGRzW/5FkBy5hzymFfyx2YYTnNmKKarNw
v9L6nVuqQIWJdZfALpKmtWtV7fZnioN53WxVWD01tqx+miY7BlkWOwQwdOlBA0gkKqKUExtFSbtq
r64VtZToWhcXu8AUf1WU7ePO76OJhycNBDHhw8YjSrzXcX+nhNcXMbMtt1TrR/h8z30J2yEAvJQR
q5eJCx+Fn0O7dQGg3Ts4bOH9yLB2yzrEqPnI7tRMKxD35PVQwZc6Pm249GGwNtJ2qJR4JeoCzYCy
s8hmBwwXfYee8iH8Xf/hx8LMy+/UYAbTHy6+H0uQ+f76JcjCMg1wBCzSLgOrNwYvqwpTXAk0xHVL
+KVsugCzr5Sx4AuAPHfFlQ+AjkzyCALRntXmXv+JrsIof2i0nQgVP4uGZ3SQjnLGI7LOvlNcbOFA
9wLP/mC56ZR9wY0y6J2sHlFXCfssrrd1sl4b5634Kuq9JtEuoit0GB3icgEeUhpGy1tnvZaYoY9m
WQ377dQ1/67OZVFLqvLX7Qp2BuajrA5FNqQdYJ8ZNGEDs8Sk8PoUyFzWLAFBEFs6nq1F9Iu64kgy
rzG9Gr7SxHKkhGxPVwNZocnUQoR7qMp6uJCXrbnaUUjb8KIk9hodPM0o2nWNSiCdMo3xhkMLWAQ3
ctBE3OxHvnuRhoVEh/cJPcio5JsgKsPEu3k9F9zQZDrFFQG/3DdGS9hcz86TAF4e+s7Fs99IKwkl
3VOi0XxXF6+AItOyurt7zdT+BGOZFbKiuOp031nicoNWxFpyksZX+NYoNXbO6o/PBZBm2MNf90PG
pcyjsjW+061gHjADvdOB5pgSBZuUen+y+wiEzgUVz+KVK6LdoEhjn5IjqMBRKsg+4Onjs34O4uCB
IDaz48uzrODx8KQ9wRS4bU+qaB1/neYPGAviuN1SgDfm+MLcM+Vxqyy49ELWcp/d8gLzcb21hE7H
GBBfwuRXOqwk0BOQcMt2vFpcb4ccbmVxZWMSGbMM1h6uuabO59Os1/x9qgLtk18d7GCL5dTUthCC
bLUtPcAK0cVANAO4wipzPQg/V4nfZ2K4ubLxoMejmBvOr0iR4L7RDMeFZIE8ZQK9W7kGbebj5NFe
0UpfuzetH7hYerWCbRBXqEuoEMv/2tw6LJeb63ryhWf/1ccMk/7tSO5IvjV3jQwnuNpJ7MfCZp7Y
hHBMHVU/rGJxvdeTc0c4wlw4S5cevzH5i5krGWBIjEtCa1CHtr2zfjmAE6XnMTc6QFb3bwiyjTSA
vuTdQHUkg3vu9lOiqX6q5NpUMzEj1Zi5h0RHc0Qc2DpPB9i0+B9I3UIWtS8xeQ97uuXweNiShAfv
NxMQ+egIYa9f+LABQPnoqLk6FuyNfKmUB8YSW706Tp6t8iR5GqcFjypjS78XtAjLj8tHyGFr98Ef
l+3msqdccz2IAWNLD7KLOf2QHIjdJ7FYsov11OoA7/DF5mw0hlUdJeSd6GA4AZi+N1V8VrKJ1mcc
jXBlptCHfUEmRjeum6qVONswoh0imexVfcO/9yA0ScfCDilhanS7Jxd6U1w7TBXbpdZs5ud40q84
YQHBOZkQGIm42LvyOoamaTyftuDgk6+5ZjmS7g0608TWHfH0DZt3APgLqB10FaIgQCrVhldU/obn
tPigJF6KDSerNKFEV+Im4DCI0x6UYKM8IEmGxzLCz0t64N77UE8xYISJGEy9b1Bj+cT4Ug9HPxwL
pDdnUaqtkOzIrgmfvPg3KR/WgIDtICIuHzJBFH7XgSyLf7S06D1OmWMMpurtWBM+FUUOuKDeK0DG
v2uu77AFjzUrQmdEStOqAJ8sdjYWUVS8KwEJMJrW90nai2kGDA1YPSTxByLubvt6OdBpSvAjBCrx
TUVdznfLjklmLQTvvrrfxSRWpP/VBfrQcTY6ZT6tcN9F0AO5bxbAyQlBuRgWA4AXKJOpYunL8I7V
uwhrXLIJPDRloHEP5dtbxVFh3+Eid6mcBTFqZRVOb7a5qprV0GaZVnhlFp6oX1Xqz1LQLlABQAzD
znE66KeLWy1q1lwwv5dT9P+/EN/3LYT9yJU9fnFLuVC/0MVlR6i9NvMARZWlT04Hl4Z756PzB4nn
hyv53OkTdeh6O3KeRGsh0TMkSgm3snNslPevnrrgW7OW3Ye6B6dVdXY1Tr6MYaEqIicyWe8rFOT/
mEpR14hanYFlqwQbXdiPV8bTYarp0fB+WNH/iKLMORTu33pt+P3Imd8Z47M37+dfr79B9lPP5fnk
4sXTOiucujKTeazmaHc+TOebpOwn1vlgeIGbsbZjLYFGYO++yy54oXtz1OF11JXGdHdArx01Ii8m
tIrxtjGIj3UUo/V6KT513QqP7oIoC6eUUOub4F1hPuPu/7+lwCMAyvkjQ6e8ZLCUP1nZyq7AiK6Y
bukfmHr1xyYA0pUfQmNgvR0oNqRNCGlSlZ8HxSK/UKJh+YEI0EYmH6KpxgeBMKkVKHH77z+tFQYZ
i8g8ix/Sp9aVaWyfo/NLxCwCetK0FYWEIWY+PXg51WEOXbytG3t54377bmyHndoVGT605VLBvmM9
iTmRJcAlN7ZsRs2tH7Q5LuUDfpuuGSSXsz1dj9MrKd8WkhyrEjVjGLx2CrJfhPymtFNIMspFon6X
ij/7bMz9y17FRyIa8gBupNKJr9G8UcQGB9+Rlf93rK478oyIA3rzcKgIS1CrIIDBiF7ClCUdrJHD
UC0q2gn3ClOJKVLLAiQJoOAqmbaBt5/1HS5gVoE+76z1rfusGd2lXLLNQMQt0xR2vQ4DcFidorxP
jZ6wwM0AYBecUOMJA2ymCxml++RObohJSD4KSsTJej3cXAYujg6SwleDQwv09ulfL2pE47gWChx4
1tUTbju5GlD6ZIRkKxWyhisvIXjKvB4xrBU5Q9AEP82e1AjWPFcF42S+2WgqYtxcmC9D5WNi9P73
JR0I0ooBqCkcT5ZNGlKONv/5TJlBLd5QgfXABFnZLsyu8BIFl+FTHAYovwYapjq+IdQzvZxHfwDB
eUjOPhe5TiPsGHf4IhUPse+ijgLiu3snaSAyhFAKgGvgubaByvGO2GDrufr9fHNr6nXkBPasyRvP
oMf14eZm7h5K2CZOT4gD9PP2s7uNeO67nVg0AVwC1LCz3CNABQuGi/uM9P0I5pK5GAh6tKk/gPOm
PUAkjarebLKogvL/1mRs/r9Xzq2DHIehYHEAZE2sJ5e27hVM8a9TMq1OQKtxVr1ATZOfnBSDBObv
V4/mkiMMzjrD5vjJ1YxIMHPmJ0O0wOVDQjkLVc6XNXGNgx1wPN8FjUSeUnLK8slq8lkH3vcDUG/l
+KXnVNhBvJB4wMaZHeuTRH9cIplPiX0uddE6B1x8o73VDYRyolEaNd41ZRCiTkV9WHG5GB5wKfNG
w1reTucXFrZF/sQ7kFgenOMZOk59ghBn18NDAM9LyPGgNU8Dw6N7eqDVXe+eX04DiPG3DS/IpQy6
dI66jWY/1YWFdqryCC6fSyWOoheJ76GQyzPvpQGfV4El2DFVO8crzg2ZN0eZbRnGR6DwZ/cuW5/L
OwMFEsD+qlEaGB/8+npc5wMM1rJoNhGrFJoXwSBIHV5vR0oZDBfC881xhG59vba77My+/gfL3dM8
q7GhxVtw1OGR1eGAKTpWNKoirhDGFdnNDe6vKRwLyFadOaRyvCF2UXWEXCKT/LFbUpTGiM6UeNAR
XSTW5v55SAHHzXSsnBeiGpUdomxS3TC8/dcFAImu6Tk/l2whmHzXQB14z08TMIfxGzpk/EggtC1G
Dy3y9HH5qkew3lZlA6NGwsyxSOfnppllDqT/INfNQh29gR8EaErAwOq2upZmif62xYYApeZCAmpV
ioBmR6G8uW63vds/8wLJ6vUMMVOKkEDUlP4LdQ58cnne2nodvUMf/eErRqRwkNL5iU+IKZmNDrek
5+O4P4/Hsbg8x/DntmDPdrZAiDg0bIUTqiNa0Vl3SoHdACFvhQAB7K/go+h7BKLfY2zc0+c4vPe3
tlQRAyCokpTtI8tE2yn5Wya7cTbjNZKPbxNiKDcjHIIgXTtPVc3Uwy+xGkFPwJLSjfQZthLnOFD1
nNT/DEARjYWa1L91Jj7pXJ8wKeAp7hsPc/AAl7sVwRSvg0tcb/y9obsMJTDQBuVXVY57nSaNEAWF
DFXrTiLT3jRyeIgOrhKxwsB2keGJIQUVs5Em2UUAExAlXpMGsDJF0kBs+wOW1D925S6qvYGWBj0V
SBj7/URgEBIKf3pgS5KOI90QNWLGp5mZiZzUoESY1+Gao0fSb2W5a2so72/J1RkwRYNGnsf1EM23
FwxabOfrE/3K9vGiJjH27WxkDUigemBAdnKgJiVoBgXXDrgLdGIRqjzz/CT0SkW3Mcyn3NgNmGIv
HVNCBcP4BdbB93wvflprkOvR7Z92vtpf1RDn4JSP/gnd6yAN4FQF32iAMFP6vhWEbcUX1QUBJ4oz
NTQoZK1Gqfew8Eavjclc0ZsaIClEdv5NxyQVXVBzKOz/CtWQUOGNfZUA2hEgwxgDw0vTj5o95kxL
BiU35TpTSSQiY/bYMAOD4CccWp51v8onAxbs2ycEOluqxQTrfxiLkkNhpOx7M6sBpvEV1V7Fua6/
VizA0fiMntgZaecTwLm79Zvs/UV4R6Okcvldyn8e8Y6qHK4w9gngu6eTpHSsvDFLFNdyuK+RREId
uHzHfddszR2E+JvYOefx2ZzwrImhpNK8pJnPm9yzGAwvPrhqLLSVvxFKNIEH7T++YZdFBhkIdbgC
ODiolJJhT26T7nsv6ja+u5djML1wye0crwBCC1oAQsuhsbE1279bpTM+Y9xe83liRX4/VxWpQ0xJ
XO78qh1S2PulpjHybXm9grNQbrHtp3XUpH+n9pY3uPbkGVEQEBQXH5w+Pwt59jbn9j226omPdwJd
UzinYaJWjur+4SHdCqmnFyrBA5doPqv90dPywEtWkqfhJ03n6z27LL4RPtT9xeh6ndWQvq9c929L
cWD2QNJl0uuz03i1/IIR0vXt3kBJcEVSdRk36PoqfoM6+7iJDlFmo3mVMzwRpQi6cSUDCrIo6GLp
fGTWZfkGijWD0sP+K42B6jZua3kfjyKWYAzrBRFtrBcA/0hV1Z2mg7t/sZFnxFSwomHuxhdul85D
UKa5rl8kLS07c/eNdnfKqnwkI8seHoV1M9uD97x/T1Rwgo/iFkW4Xxd8iPrNs396K0YaVq5aCCC5
bsEJ6weo/6z+KrdqHCmX7bFHlQ0rtSdmR7wTgnu88QIbNm4zkj2+S/M4ZCz+tLCEzXWR76U9SdMT
9mlzt0hmIniwCC9jMig4/QJauXs9+z95kKaRVWfQ5yo/5nLJIqKI392pDA6E307wbKCuYsaaJ94Z
AHoRGZoe6axSd4N4xaJUIMp9pfY9Wt3FpraX9QDgSkqTB4zGHEG1MJd5sPhoPUx+Y0zpfAmgL0Ry
yYxansPUN0brVVC/GewHL+X/QPnSBO1EUBgCZsEvdJT21TZODW7rq887Dvv+6Dey+b2kLB5uam7q
QvN4q/K2r7bFl/5vj6qGhzr2dSEEYlh6knb37so8bIS+st8liEKjHmFmhjHSZzPB9+OKbx3xYSe8
Za0fRt6Js/9mjISC940Y9NZ+PAhEntcyY83CJ5WRvn/o5pNlhQYkWxlipJTxahmqJHUKvZ98K+Rs
niVC96MqOzXhSMAYIjRiuOsxbS3rlpHdDv/gVsA8L5BChl9zP8bgPu1MGx4sqZhjxz6XzzEtdkHG
g9hXV/rVNRhMOe+bjDcCeN1NQnXFBaOzOHn9oXmqzKdwOZdTzFbpftxa95bylTVmHjuMQ86vtqdB
epjdwd5i0zQANSEgsK54Y+zjKwwRYbNZk+VXPdqRqS/pEQbyddZn10NvLOL8SMBea6/+IeYOSWuE
cfFGSDM4uQe5V3w3WAmj163+qJ0MVHRAUFZC8K3kAKGd/GEi2KgolC+VgDHt5wjpUUjFcYQO3aX+
ul2QTHTG8w+P350wwJ9tRI+qqoCQJO2XC+QQ+VGxt81yEoZiwFspL31RM/A16+FVB8CFbMjxBYPI
7AgIyZ9MeJFyXGqTnOlqnVjIfUUav6oLax672VaBRj3NrEA5SMfj8FTDNSs5y3ecJ/pUBAUbN2hg
u3arPD7GfIZxw1MYQlTOE4Q94EpOx1AcHBJEhq0vIiAjhGIPmgr+VJkR/WnTOd6XvhrAkwtJi8Az
RcFSv7W9YCYCrl/sgoqMSD69d6vULdlv7Mzr2IKR/isrvMtHpOsvkWZ2Cu6zXyDmXxe8wa7gZDpF
GZLDB6ohlJl5wpKIqsgzojBJFv5y/wn3KMTemswFyGjeTiDPFI7B45/sUH8YYEfFxP2s2rwDomnM
XX7aVyt9FsrEO90yoRBjCh97q3uwt4KNXX9I61R4H6FNU+vBTFAPdz7C97grM4vzAjdJsEXQtT/B
EnXBvXfW7qOOooAl3cuoKk03XfvGtfxp5T0zLLvd314nA4caD2e2PxPse1pijyUwJUl1mU9fZrXn
Z9RHd/WRfR1WMV1BYawnnoOfrD2hkFsNGPCgtqJcQI+kqoavy+/kMzjM+/NenF46Zqm8UBlcGTON
+ulMNXYGuCCJiVMUHBqeeZqvtc5tadMpSwK0QAUni7P4q+UuspZyJUFmPsdq8t/NnhetUV0jatwB
D3NyXqZs2JAZHELxvErtYH1wo+bK+xEv+xvAyVkxm58hi/gW+tbJMdLirJ5CCakF/iHGsEDoG+b8
L9lSAfYaP9uo6HV1zYtXASzunxRGrLwH00ypggjBTtUcuoXN+cISN/yOFWuGYjZTM28cJHtNOfRU
yfuXT/haVOnYGmGVIA+Pq028WtBgkKu8IF5tv2wPQGTLvjMUNTPzP44iI5tyXKp6MUsAuTsMhbp4
/qncp4KpcKpUPSbq563WsBRKno9jJGrvPyvjjhWYA7omrzygfjTLRxZdQAIF+StzhwRtDQCfITIq
BwUEhCcWuZpP4Wh7ByAG89h3a+15OEPeamNzkyHgHO3T2J+TXvrJsUa5QsLAhLqM8yoraTqPnoOZ
kLCUwQRhCSz2IWSg1tgQsNAfy00N/ixQkKwCYtMjAslUHWRaiu5zN41YnLAtlBaA/Csg+AG/j52p
J0ztcOSNdbldbl79CqH4mXR+oR1UeRhF6Gh9w+xB01Zb1qUFXJQGcR9wsSKf26+NA23Lr9DDFvfO
Lm843ZBPL1is9uFE3mSXvhC7IdRWsDoJ/piRdkoFEHZ94s54rbz8Z3V3kvz9W+KiS0NKYHZ6AE/E
RJFEQmxXDpR74cESrTWhtUW2hv0VZP/MM9sTu76kABQzFbTbNLpPv3SluAMDr2DxgU+bF9dO8iFt
l9cWIQVMEUSbPPzoxM33/C18ZBSBQlw8Berf79fJtLZWLwfxu7cu/9dyBprSPssg9eGcg+bHHB8m
og0snre67GEqVH6w0ggjttrBqigPnZZXavs0gndbBaELJqIeekiDu7QYUBm2Xxa5PZTKsFAYew//
7Ioe+UAL2kubIHHHIQVdp/yCyoryUgZsfGHVfk+H8kb3lmrM7WKxya9ek9e9dRMyetuf3jpVWkkz
WfAD0Bp3SLHcogDugHJO1oF5MV65HPzAREPKVzAi2FuASerdv+EurxzP2nLMC1BRt4LbVJ54Bxrz
5Omj6YtFc5zsmC6B7p7tsqgjUaXg3jthu0WAXi7ZTq1l0+zMsim0aqY40kZ0BGBPIQvHm+ZjgTt3
da+EEdFOfhVScYzAf/Ed3rcpVmrgGwAlgmjTPcC34/8LymeQ9j66Sg+9I7uqQNVKqBQC0Z/i303e
rl0NE9/FT9K0T620zs+lrjSu/CK+8Kl6piIHDBE+L+vULaVl6NwiQmuYKHCqrajgMow8Xia0SY0t
S8HDmEh/bX2OuzDwkfXqxY0BbUN9nCOHpMs6EafqeGK/gU7s1DUoEMP1vYRnvcGujWzPwN7sfQCJ
31lD8sBk9a4upDIXZE+ZKcn5hmdgFD4vw3z+sQE2eTOs62OLkxH2VM304z16Fvn0ZfraP5IbJSrN
dVwjG35mZGwUnKETrhPzYB8ql44VWa+RG3UsnvVZfxnvEygtsO01UBSGRmecAWwLgTvQXyWUXS0o
vTARq9rn4ERD1jC8sy1vknpfiL9kuvURZ4cKWb4rCUQrFUSF3ELR+43qW/J0gxdC1MVMIhmTVZum
Klxx6olSt/AxoWbAi4n7sEyH+kVU/rkdUdN7iPliecgn2bSKQG1F6OnjKvBJxLG+RRjPxokxGwhq
GKtLABSF1LrNDYhZWF8RaAS22Ox3ajFnPruIrwOBchYA4FnF28nWNqkBZBcsqs9RDTUzLGl0EkfO
YkPHYkBlrywiLPyoKaWlkibQ0wQ5CHP48dVoaw4YMD9Yir40ITFnIy1RlUd6EEQ+qlo12A0xBsrt
YYKWooksEWOf8dxmQXplClz+nSAjwB09SHOqxwqG4eBQPpSiwT6cJ/C4bc+kVWgwh8SX0hnezUkC
9ZBzGSr0oGsbsxI4qZTV4n6S4edSTWDNv3a2Cj5PAhaeCAbFjgrYZOoibuhbSY/zzM9FDDeO9woR
gKtN5IOziyEaMHmRc9JpGWsiijjrZdsdA2+3EE32Wy6dTNsp2G6jdFPqSJJOCJNqHrSuAr4kuWik
DNSpKhWjpqWyNJRosnoJuf9V3kle6tcl7hyfJ0ZJ+G+P8nH2x2CvBcfv+IY6eVdPBG+ff8i6o2+I
VI/XtkMD/tGos3mKHT1LqFYMjI/QMng87A0/dhBGFUpWcx6BZ9Q4YFbfVgzBmPGfop//mhn9O5g4
dB066gKg9QfIwDKnISzXWSj+PXkXJzMqsHcR05CKEXzXf3pJuHDswGTNBkBx0zwhel42z3gUpGEY
XpNFC2f2M2jUEK7nA5qMBKaLCBhmAmV/FvoHX3jUwi5dIb0MQTfyO+nlzeJVygeJEDEHdjr7YEcK
FzJfaejuy0DvaX+LxFK1gHVPiXSsQxPCZuATBHNJOxScXqzI8BOptPSdRLUbx4R2InqrvzFdxRT2
Yh2z/+pGVC8mdiAjSlgGVPs4aPhNRjL6sxvNziJ8eyE9z8uZ1mYEfz1MB/B+xOoRZEaQVCQXBtFq
nYmChMttwGUTC6p/2kVU0Y7YXjdEvUTO+IpnCoNxINKNI2GQMyetYOCm61Xu2G2uXCxBzLWXnxCw
m4wA/1FAb1Tw7/OUkamnDZvyiRjGbMOOMfYIQcCgG16xz5PuJwSELnVSj2O62L5ilrqEghtnOFrS
xUCqUPsuKUOF3y84eCaPlbk1fACG6/wQZQgYFS3fPna2g2ozulZt4mqVjgNbSAd/0XzUCvBrGiZY
f6BO/FlWRebyhjs+w9t7ajW6rHO6kTrjcS0eyieDPigklFA7F/GtR2AQIupnFVj/MUyiJO73qtZ8
+VI0amRLyMQircRjvx0lxjPi15twoWnqny6o7aRDRxpV8ecoclcCcqafTQa9C5V6//Pqe9+cN2nX
B+z4Y0f8UXhIzzVc7/t8azdsCuMZi4c/XQ0cYDPVPWq3pCQJ2bMp3S9W8hXJzERrEzY+i4AmNa0k
nQK0cbjhnPntVUljPS95huNaiCcJhhJ1wsMyLpYXGFW7Jr9ocCK+zn1zs3R7aom2uwksHqM9Sy89
c/9XGOyE0SBZh2ywGP1f9eZdxsKoAK+TAFMEJ75Z7afSqaFFRJ24PrfhK/4V0Ca3YM0+k6rEDvc5
VAhxedlpJLKppjZ7MLRMW2F1JBFy2IW/5Ovz7kDNaywF/qgxRjzjR2ZJBnIObZlYJcBgB927JFer
K4X+Ow6q8KZFlYCB4mJqel/kjj/Fd9Y7efkQeJfhkziV8Z6zsobODW8HkzvsNhuwm1lIaFKORUC1
yf0dzPWrx9GsPcTf4dvNrvX77xgcShpiiYflSb6aOJtbEayUlZias5l8Mulf+kNdKCaOFOsN5vlk
ehjFm5ZNrjlRVelmcrsqJy3TtxQQgPs8cAua5hDdrFy7CKNWY5rW5E/YHrwZzO7EDx4SanVnduXD
vn3jCSD5nZ8yAJXm2Hx0kbUfIbA9CQ7o0GXuj4U/tI5Di4VywR5gJlDltUjibzTyxLCgH/w7YIXt
EJpzyPBgcOuPJUnB7qJqWztI49s6pv/+z/+lAV+uOLLh9szaXzw4
`protect end_protected

