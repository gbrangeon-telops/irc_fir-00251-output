

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FZWxslbw+U6Wgup1K8ZmbZ8ZvAwEdSXoQX5Zxu+YDpvGpSAvyJJdij56SPMVKmhf+X7kxMgvbsEm
5B5AiAyVHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ntA4Op0vLLt6gLQbdMxO+e0Bhjub4O0zQAgtU7SVthNE2o/5St+SvTkDoJ1ve5MFs/Rgt4JL1gtd
IBaLjbwdyEGV2JKFzmLfNOLgk4U4bgeRTGAx1e+I5wKQlcq6qarG8xv4yuzAX6jRFWecgDUKdkZr
uIZCcXBmuErGbIdhFKI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I/9QBkeb84dQg6xWUGWLN64S2R+IIBcNXAJuDMwqYLTsejjUFtntzi/OgGH9xu74CzmvMnJuiSkZ
p7NF+AufXfE0LUxVeYNmvB8UnCKeswDMIWMuVEpX3XPk8OVFRqBWCRJ5c38XRjldLuPPEii8dq/d
MjasuPQowI9n5pgL7s7SczhrYfNu0A0XEQTAwaUPGij8aO4+LpdeoyqZwdg7p9EXJlysFsw3bvdq
qHiouBqf7MqPbKppmCVMlrH1R0q5YlTlllFEZblTUq4IO2ZWi+5zgGnEERNaNBZQ/na3tnrwOTGu
mqAR/EaIPbn2R/AR26ZYNuBuu0Ym5XtWJuqzJg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jRGmdT13qAzfiT1K2NPIFkj82nI6QO0hHDoQ7U+cF5NSt11k+3KuVBnDKOWta7RjBJSeiJs3q5WV
MSQx2R9/yJGRUjq6DQS8PVF7sqUyuFjNc8w4wdPwxcG0hsCFj/tEGyFHTU90BhMVIeVjf2WlERXd
+UzGn82C1ATZxC/M3Bo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c66DzsXEGPMNOrzYyBeymw4AV+RpL9x7eTO9Hf3l3y/JxC1wwEbipw1XtleybcrcOfKY/ACDBUVi
s9qFxHBAPyb46Eh9l7EGLGzxXJTWMed4eJI910mZ+WMPkBgIF1jvUqr1JGStUHDdUjBjqP5Bbe3m
2g3HBNLeS+8Ciq924vg/jBwWCA+G1zUvjlqI48sc1XMFszL+AzQf3r5t6tBvdkd9goSPiuISrM7C
eaSWriX/kCtr9jogh2EYVx1Ud4JT59uRVRlS338jlkF39xoR0AXtgdhjpZa3Qu6PtAnEwyq9aWWk
FBo+MHknw9HNH3v+t/wWSpyyW9f8/AhQrF1o5g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12512)
`protect data_block
AUtoJsQPmb4neZzBt3u0UEhpZUSW+OlixxVxU/PaQG5BMuTYhZOn2mWeKn77t05b9BRB6RH0DDss
Vp7I6TOs6H+D0M7WA1My0/d+Tzb9N1cUhiAlJIpbg7gKISpv9cJx4qrm5qex3f2HmhMjUN9zZ0Hc
6DnRPA4bZfPE0ygrU5KJEoYwblhsistategRgQntqE35VGWE00YEX30aCLWa1V9vIBgTNeWqofWn
TyZ9c9QGuUybvEG1z5BwuWQv4GR6iPu6oI8lu8CSbeszKZTF+wFP/IQjfjYg7B+cpHSzBBBKlSIK
rQor2VrzOgccIoVE3aN8oDelRkZrQWsaZxRarYRRyPr0F7BeV3tOW6Oq/knZEImvPIr7QvM579n8
cXwocRxUO/wvXcobw3zPp6mpIiW8Sy+9YTbbEO16bZbHZGgYz4CGLjSCoep7jrtMCoXJ+lYRL6wC
A0N3j8QFIjRxcPBBXNYTUXnkrRbOtLmAscyZF4f2Dx14MGQ3xZhSsQHZI2DN4OUUWnCE9BOjBK71
WugQd6EMqaHG6hI7PrRjA0RWNHeidx/ExmqrEeO+xI/ivf6bfY/IZNRIeJUZxUjDL7Fh6TS/d4o3
Tq9sGwAteVLmAVudTmQZ3OEpZDTYXdScR5H2KvqTCUjUipah1+1XH54Rc6yDNkTpl/6KUhx/+ShU
l992/RF0ijjZMu9c2Jc0DgM898nkto8F+ujADor6jfzChuOd33g0qvOw29tqWfI5B3zyJ7uvfpUX
xTIMjvgWV+uJsAT5AnkfXtd+/I3L641nA7Sz5jPPQIUDYNHJuMEpppMvBS1y4bN0oWNCt/C+4mGg
1vqXF9s8uMOvw5/YDiBEmOXFCEYoB5K+0TOhXpVQ22X9ZgUahPQmS4uffmz8o4kGuyDJfqJH7plu
Y3RIPObmwThol+v+xQm+GBD9Ic8yQriftSZUTcARKfuPYBCfkNXKzp/mOg/7uMyL8u9LR+NLUiXu
bM+AJymohoNrxtxQO+O/9es1FU3ptwxx7N0ilvHJgvNuYrAagmqyV/gtmDTMNL8bkUwve88EJKPw
FwR/XMIK2CH2t6bGuNJgTnFR3wUkQsmUWdlOZkHCJnKf/29QyML3QUxTlTfpVpB45pXJrc6FUbsw
JGth3csfHNq1+9BvY4nhUqtLz4fg7FYRMC2YgP/ub4bmghuQj3TklhLYbkwxsZkwHzJkrmyBXaRk
npt/iDukvHxd1UPUnwfxHzaCgUZORE0edeFND+fLpD92RhTpMBVW9YHmzh8Jw75sfND/w8EMhUES
ppouhSnnUY1ayADSBw363r5g6BbAvWQonKepFvCywuEU377PqRuprhMuBw/vQMi2MOyf0CUjGD7f
P69isTWt74WGtB/J5NcQ4lqo0RcleXqpWnABVne+phfyyRXlVOIWVtj9PQ4JYCzDR/7+TfKGlFgF
MgfqWw7VGBMSC9GVXMHIiJVtgMt0sv3RBbDJ2JGkOUx67nqK6aAEIwuBxNSmYzuXe9LENqUeoaUL
gM6lRJx43P4GYMTln4S0MV+pYYhvLa7PYXIHZKwHMKcOAo0gNaU7YYvqs/ZtN6T7PdQeSBjBiSqR
k375HKgMs/QNxuoFOkaadZlhO7ckmbcZQXGBjDgRaHmgeew//7xph+eiOhjVwJuBuNbGp5w3ZA0v
ch1bK4wIKpsu/X+IizcCZ3Q4ve+Qx4yMYrdJxhQfNRBfTgaV5Ep0flUw/gwq4Dd690ILTCnbURB8
fre8yVk350iSWM5lDOoenG09UEYoKTOKPuDlWfbDG0tJXXWMMs9dtiiv+FC/hFhT99I7cr3gZetM
0rybplXqXgRMtzlOvq+yWVWtSK027rvKS4gvJd0n0C/fTLXP06CnPvUAl1ZtHqt6O5Xmhp1p6CC3
xTJ0DnGKvfxU25KdXuSfx0AQZpWe2ylRSROrj2O2TlRjY7WYV74lN6ztoc6dJ2Ibtizhq8rJaOGp
ViPTD0xz+k8IVLNCMuO5uwHZ7xFMHGfWs9LjdYqhyRPPaNpbkowj45W2Rdj8lp84L7+dMxLmEw+F
biwxPmz8cNThV6vEUEiydZifvaFu1r80EUQSH3lVoYxDBGpuDfA0m4OPRNNCtpxBAa5wLggo7RCy
FQNC7uvL8YPuMCeTsvNVtH1OfnuhOo0BhRpuuz5oP+HnbRDIB4jhvYcxxTbqEpR8bWJVK8IsyW7K
nHXPlUdypo21qgaRIWTgxv4uS4cf01ODGxdvE819nMVM9DMW4uJzSE/Fj48LDEDxMAWmuIUXOENF
SxAhe4GeH99MPD41TuKWlw4dMyx+dz2K4CmyjNJPmQ3C6lAhrefhUW6tcTf3NwlW/Z9wPsWZW5KR
4ix2W7n6f00lq5lfMfN2qP/0T8eCQ0tb1+kpdOyStha6ID0dNepEa9Yaja60X8RTRcOQ4qFP4A3X
gph/SFbbUEtCQXaVoENLxOi0uPHV1gFa0pomNsBemWlrN9E/XYvLMvdwgwnYUiuoNCWvxtZbAw9r
T2+n1yIq/vs5mSM3TMSh3hvhvXPEd1a9QgaWGybS4/K1tF74C71TjY0Cru6tVvmjpBUMNOa1AoJG
QN9ggKW0X8HedBTzid0IoY8iaxeWb83MsxnLUh3QgamGhxchU4CRaNAhjaVPupzV1dPrfGA2mj8M
hb/BpujvCWBoPNfWNuD+dT7OTbBbxAa7yBF0o0A6esTrSsWRDxkMPSsf5KKw/qP151zFHXMYdMSL
vaXw788n/dlGtq3MKWuHW0GJ1R/2xjHso5vrQiAcUsVSCgJijiWHioBx13qGfI8greWpz0peGFJZ
AzJZFSlHiyJwg0BkVTAJhp4pg6JlK9g5rPBeVbQEBnf+NFun4Jc31BuGkGoipMNU7Xn4rcav89II
1K9VGdspz+WFuZ3aP+RvnfvI0WZ6zKvJMLAZVzxL5yoqSv8FV0FsVJGAy/PjX+u/8gC/efoZNrqt
mi/yw2DyZKiN2Bu4tLjlqR33t5yWva3Pb2eACripDeEQtiO62vangVvTDurul4UYMqhkOH5DGoBK
w59JVEUXe/zqfkYaja0pSa/umYVqPzBC6KFLMDUlyvXXvOLB0necQn2nwON8HYko/meKfLVx6I1H
mnQrw9ikHWS2vnwdEf0ogxKWrjcQq8H6bzPU2GR+nhucTkqHP1Q1U15qWlGSCcfLMchO+ijp8JNU
H6axyrPuF+qId13wVWtuXCQco9EUTJnLrFaB3kU1MobMy6EXRg6QCq5zz/hIhHi7n1KqgNgr6yUP
KSUmyAMwBc3+zGhDjGFpOEQ+JfrpuTHsl/lDjqfD5ke/LHh2y60Ks0fMHMRRYfGCuVj4RlCnCGU8
QPFdJgMRN3M1Du5yOFevwUNFIyYFkwo/NEG3zxGqbjNKMg307lWrvPxtz48Y5DXIecdPkeRxD8zA
jxAeYK28QzFa2hZkg4BQsipUwPmjGcYNfs4noekep0O4wxr6/MzTi+0Od0B2Bdz6v/BZsASkNFO4
uRAOLIfC3aPoAZLoKPlQJIZAc3L3eNicGqwVGY33+CcxkHimYZjCHIX2zCzSWuzAX4uXj0ergqkv
JVegq9m3Od/ULYZf6rQbLI3StdBmt1RoRYr6N0tfSaKyWGyzCuxl1cQWqJGjXxX/grGmq34kJXQN
3pIyjGx61qWb+7aroUCLfWrfFVLL374xM2qGE3hKisWovJ0+oV0UPS5TZTkev9dRdlO9zErfjjgm
2WAlzQiIJoaa5mpijRn9viKPmKunzZYDl6vibppyu9IR0Ph5ayzungSEEQ44O8dpYMB87R0GrOE1
1kz9h1H923OWzjbHXs1V2BKT1rn87hxQ/lcxKj04MkU64zmibzboM5xdeyMjIaWbZBQ2ZTiwmNHC
FKGS7HILiKTAqcvvRmbf2sWMUW3Gj6m3jxBzkHu+EvQA+WV3rVNdF1Q3JfDNTw4MciQDqArPQaEe
A8USDTlMHI7hobwjKTi50lDJi7Q7nPsFRcxKEQ8EBW3TgjBZZhQVcb9DtPaq9Jh0+XwuepcN57zJ
pcPZ5OQDE+S4qZOG2+amSFH3qUoE20Y9VfuAVykAhL8LmC7lEBdSAjvzlSDEZlhVJ3ggVHHSaDjV
E6pnSXz1Cb8p4++2Sf/6SuMSesHoKnEq4biyZaqtLkMB9f566Fu0n0dBYruvgB0Ii/ykj8xPn79j
B1OtTaKj5drPnRm/l5qhcUEQTXi8IlCIKwRSJyzg7THW+95cdhCBpmvoM+XGha8d1lwBJ5r0QWYW
aiO1Uyi57nuwDoYA3Nywt5X6D/UhbhW7GaQ/rRinrf4RgJHtYkpqNdVjkuirNleQFwP4mkLWZ+mD
IoJ3EBQqjr9VzSHRryQhtCNq6OXXbAT/psEFO3KtpNiUDneC7gTR2WM0V9xPgQ3XwvBzc7szEnXX
Z1Iau5tBfEwEW31zSY3OO2I6FOVURTdrXuq039uSTvvEVzBrkSANzuKE14DrCIzV7OULeIMEI78N
6Ql3NS+6ZWkAhKaylrtuAnvBbC6qAAGCIMIoLdJEjieSUy8SjMN6kpeX/UWYsPNvP90T4KsT/r9k
E0RMlN8AoLPeAz1JWdCu+JvhErEv1fd6ne2cKVxgxfL3HM47m7m++L7aYbqkjurQhHMV54mKTgqg
X7vz+XEj03X5yb+8oujlpT2mki7Ss3aKud8fpetfL0QIcJTZKXFPgGzcv5VAbuIUsdLN8yl3TMBB
vZiJRbogjgZlXKlN8uOPmjz0HQ8fNbpa8Lt235J/0IgeQZt7qd8C4iE8dMtkpalYCGxEqeW2lcvD
kKEsIvuxrayi+fk3c28QncoTJEl8UdsLLXCydOyHgrqVGzz2L1MIUvcPw+y1b0kkFR7emQWhlLaz
xrDnjz1ChS8zgj2rQXP/qiEl46W1J2xVvEHgV9FhiH4pm9CP4giQ5dooai2nEv8z2A1onSnCiyL4
cfSzx28wFXpE6xRsPLmbBCQYCF+7GaVePU+AXprz+oTvPaM10FpmjrsuSrvL7UEswavl+YzagBd0
a9JqbwRUA2sY22UEnFBTuLCd02V5yXDv6UKRQGD3q6WEV9se5S/UoLwBLUA9n1WRc+U8FUxqhVNq
Xe78VRosQNxOEFVy8eLIrpzgqpzdk4eXSjjmxdDqwsi+weag6LcmkRnoquVPOGlf7uxcXZ/IH84c
10z1NciyxfbzS6EZjjNI0XrJu7SAlu/TtXDN+jiweH1k0F3se3qHXE1+f+9yllDW0yJlHqrOfKwG
+L8UY5IcefHc3QxVHaS7Vk8cShBSgH3T8sAP6BaOfDGUPvkqIF7si8eecKelVTqAXiO9+sZdo+gz
qn6RUvH818eFjL0CK1c/FQD0VOHvfR1dyGGPQFpUbSY5A2bOmYmwwerJRvinzMRqsxW1TYeRnbuk
XJ8l8s6oTMGxKMOZCkGDFPPhCiBH3zGCNH1EOjePoqWFaGZX4ECGJdSZ2G4ojIlO9UyGcT8Ff9j1
eVW2ycML+8gUbJedMVfWGQrO+3GCNOBHYVsZLwByIvtbqEo0/qlf1Ypn80rV8fl6kVdHKY/HPC8X
qsezLhEvzjUMKTWZXXxWbp3+qn8WGLtEeaECgQQ8I4fQ9FKFQsz6KetVkVnkra8y1M/ceXHuch1Q
t5o5Tot2kj14lEoK4Gx4K/Y4DZDpFAIcVLoF3t5+LoiErdzDOZ9JSNxMDwOZ3AO8Qurw/lKnb/I2
AoKT2eRPpcdSirkn+Dn32D8X6QiE+kkME1RyTmPj7KL1ckBKJHSOJcKU+oVUPQ/ohLhVZ+4TTBxv
vyLbIMMcweDjULjPGMWLQWxJEp+1CSAzvrVCvnuZhiNhUWkQcBT3TPAz3H6airedHVyV1/k9eqDy
cdr3Bf4CU7EBeZqzpAx9CXAr5g9NHIxbTizIL+E9S15FgPkg5ZcMJsqDPurB5yZmgbZakQLBbXen
bFvy9s91Z9FIDbAX5UXCIduasY/oFNXX4sCUjGlg9Yj/hO6u3I9DlROci5xifM0AvZG+1Hr8B+eA
LXL1v3Ufgw29ARkKZzhfeDzSJguBeOBb6V13CPQK+wLavM83+KAaqmHCsiOIxCZAeobMfdj1Jv5w
r4iCj6a90NLDP7aMDXt8qqX6j85asboCMnDWuJ08kYU66+K8PbXkYZDui7110Qp6DJVgeKZo0RqT
EOtGUX16tmGhQo38SGt7dAuhd86+s3qy08u4JBUeLVhN8Bt3/orkAYlUBk1cQz61cXaSbO+jUdCb
j3urce9RPRKYLTpaedrJDzJAKkWS7yDm4A6PA85R7D06+fmeAMvI9fPBSQM3ZyuB5wJqWxeustc1
6lAi5NhCWx4aTSr9FIzg7WxMpRLm3PfKWRY2dOZvGY2mY23aoYURTwiMjQgTD2K6gcdoJLqIaGMK
LGdoJiDc4iCBQJVAKKTY6T0UGP+1VHiUi9wssxKShPi+f78+d3vuZUYNbGw/PvaGBqus/kr4egXo
YJYCT8jSLUVLzxXVEh8fyZ+J7L3uL0Vw6sfHnZYWqw2owlZdPtufyfKyeSiCFHaKqUZBAwDYPkwZ
m33HU4GbPHnP22QPigsa5w0pgLTHkC98TK/jC3KpVInr0I9uOow45w8RTO5GO2thAoVpXDbWzSC7
1A35XG7iv1dLmq9jB36ADzst3szEdsupSDHFwO0WJ8p44mTOfinGEcPP7911cLT8rf+2UtcVwIT2
wD02Kk/kQKn+jxR8l0Q3HBYb9cuQtQ8Bj+yHVQmfj3ns7vGZUbsdBs4wrJHl97s8cODa9NcRWjR5
Q/MUKAYv50qhDWeYaJx79tKhPBDUvA84Nbdz3eXaPJpoCTKjvaY28Xi3IAOEASJDjHIHFqLEToCy
EXs8vSo2abfjqmEP81EdfhNIRD5dVjmHLVOVXWt/qJ/pxc+mXsJ/lG3ynTpWDe4qBceJdARruErv
qAwfhhE1jHXSV3OyCgjnF3w52WXmZNuuhlqQsWqOb0b9+j6JB57NF9kqGcB5LNEFsTOZkO2z+9ii
ID1wFer4U3CIGB889Iw0QdxmWDe7fLvEukSthhFycsvX2MV+eVvaQlbGwZPS6604mLJLyIgkmlz9
AikgXPdPWHKfJIsYuvtgcvuqhTs6aD2fg/WA2NObLZkYpYamKKPBcfmlQIcnVTDcSA1K2QI6XUU7
CD9RoMDBIoUSg79e8t4tdgZcp3cpah/pxzgxPxo3Fc7nw0NMf8pJe8VUr/EyHpjuN0kezXDS5oeJ
esFlBEeZlEvhjs7oKZNbzHAAgamRVBmjgWEkZq+enNs61Kukd57mMOyu9IoFJO8VIw6Wmsx628J8
T5DLjihTFfbaWw02Pw70j7rF3nEDKfPXhWV/xloid9NvOYlPP2xuIX34krg57tJ/JK7YvlBGLAPY
Tb8tBOqYxyk1Os36KPK4hHrr83lqbQw1NVXMs2/CoFdxgO2vYEUYdTHXAxtmZwKejNy3HMCIvwK0
N0QvNTmYqcvbDPvwpijbjOoMzAe/3dcUJY1RJqo26j96+SvEU/iA61hZbfk6p0sSzXjGuWtSIfXn
QtFYXw6Lo3D5S/0bsZyvs+LsHT/T4AjaNpNtNHMwjcie5amHJ6mHG6DDZNTCrgKWGXjRXKobydrO
v4b8c2PL7y/El18FHRiJyU2jyr7UAmLDoB6hD6Nw5Ia+IvVjb79g01miVZFxEaGzeZGxcYPLJ7iw
zKCZ0N5FlHd+McGLlfswZtQEdnG3rNNj0EVMUxE03T/gytV/mlze0gfNxMECdRdrXcT+ZLIUgaLG
1I7+TPxVbGcmyAlghX9UsFYk0bgAhG85OTXJuY6aiSffM2tQ0b3UE1l54RmdKS76l3Sx3SL57MPk
Y4c4O2HkvzYaHUGksX8uL7WGJE5Ypg0HbRsqEFE8obTIzneroa+yUeC5grorq1PlGeYSWybujfwd
LaaICcrAJZMuV1dTHgyHg/SRC+R+59rGNE+EjNrPGLfyna58v/gGyDMtRLRCE8CQKMSFFqv94iky
W3CcoDgMrlvUe0mwtk35mJfvsw7SQkq9dEBvc6KXZ4gRwTT+Nx4j4Ba3BzET+VEnJxFqfKCYU3Nf
QV0Ite867hosT5RT7oVo+5eVTDVOf3HluCy4xWVF73wf7405LR0R1/WSCh5mtKYBaE1FXmbDGbLg
6q96b2XUJ4mH/o9mu/Tzu+K/O91th/x9li3YUqsquknkTWB2pxpHivIlkj+WauiEC3kminPxkLWu
eGJracNrSdaJ/WuyKMGgabDVyC8p8Ei1NxWXgoWSzS9WJqS2JqRbN6eRm8wSSPG+EVbn/r4bFWqu
AiM/TTCGyMhRIDBNnmoLUUYsSRlq53kjwAifFyYYmLPCUmoNgUFMG+8wXD7L0Wwrgo6IJ+mRB7dY
mS3OkYCUph15HsDixkUJzB2zyXqoDt3tkCf7HeGfv66WjaxePfYfBKEBEmDCeoS+zLZtlYnutnTN
AJUrCqn6lPNUDRVw3Q66AnzHc3MEeMONbqYdIvQVCJULHzXpVVdydge6du04ZdQ/l6BRBk2GlOLH
wFQ1Ebo7JDHuAZk+kls7DGC6F5dgDtryJqd8Iibtek0iLtsUndmAFU4ldO/VRHNl4mpslnRbn73g
0pFhsUE4rVRQYQTldeVFO2QkNbXyCX/UjQkJTCux9whoXCmL0oaHbnDrR2owyoDaPgEABcq14xiB
XohIBHdvQ+PhTxU4V/ybx7BQ+/8Z4DPErFwv8WALUMy32RcSVZYTy9EcP22JF4LPrE+J4MSibGDL
/OJkz7eprO47crxY58h2gxSu+pxazm5Ii30xVsp9Yk3lUcpW0WRiXIN7WeVRGaMeIbdR7QXdIoXe
iXqPEkrEm+7cVRrlMer88jbNSg877mPSYp4+YEHgQ/woo1BSnNM62S7vVLGUSEc2McHtkjiQIcTA
lvFAx8NHuHztNxHqBoVA9nWMT2h6KbPi/l6XHrRiyFrb+kdztatjT7XpXun6M0el574ABJP1X6ci
V6CqD8p3SkwI0x5yGPoPpQujgLFYwe16Zoz++FRyY0/FAYxWgiQMpaqTbH6HJbHlH0YlHtclOJ/l
1+mkjJ2No2G2JwHRTLJVhO3hV7X/3zN+pzdOfleXa4BzF28H5TFdwb1OCPDi0XszH9vbpi8APTdJ
HJbtZMTozpbzJV+xGgZcI5b9tkW3fZXr7IwEBkp7l0PllN9jwcMIhj+7284KD7mVWePPIgk7hAKJ
+jAcsrDJuiyNfyZ+rPH0/+cTrgWjeZXQtb/kmJ2m3bWESD5h4j+DVTMbmRY8+A6wwaojPAKYql2O
l3VkqekvVEkDH76KAjODY8UqF/jdiWvRjoZg2KczPgRxWiaL3fR/qKxzseaFenIl511+0PG3NDv0
rDYT6hSjnH5JmGd2fI+xI2AZqQ1Bp/F5SX1KLKvHoORqfQAEYD/OOnhBeDC0LIvIhkufPKJMKghQ
4OaAHSj0obPGRLKYFduYJtBSbzImCDQAtQC6SGlczWVJVNHqXwYf6A3XSlNCrz+GMnen7MSYewCQ
09fVcW+k6DgW3bzSvt18jBe4YHl2aino7ErsLwmLGHSivoOaR6sjvRigbdg5Urt1OiBP2GJg3Csb
A8zv98+ntCKPaa/GlWDM05hKnPS9TyawjsjbNm2D8iOh0LjzwWmefpaMx7m1OG6DbtU5W4QHnNEw
qQ3gF7rlj63DA2Ewmh88JIcBCw0THhbtRbfmMRezD0ZquMMyBEN3ALWB3Thnxl+XvO/IpmTuIJk3
mHM3sOFMhU4+HG28/GtuTOeJBF5SnrSWyrLKt9gZQeHR3vhoZHzWN2Om0m5GMyV1bSg1bMHYYRAZ
En+ZdaXGn+EbYTobDdbVB7eoX4N8LRHOAJlu3Mdqr8/4X+olhvSUCFyY9f51/DtRYlEjn8misuS0
fv1TSCXCaIBIUb0dPs4VoZ3eh6qBWHHFSN+E+NUrq3R9b7a9Dg1M5s8HFujm6xWWIGn2eSjPVE2N
R7pA4+MqKVgbikQqEas77rQedYxmJPZxqN9Gjhax5akqBneqoFMeYaQ05hxp810lEpmzvZLajzO8
nuvpj+iiu/QeTLJPnFn8Q7t6jqz0wSC+Pf5fv5ASMJT7MVZXF7UIQ+7kuPbHeOM4ErCvUi04Llzo
VPteTSwnGMeB6CPof5YU7pfOOUk0psKJ2zfU8bqZ0lNSbHvusnOJBhLO2utIiqItGYssrX0TraYc
a6W2+BX2X1lNigkvQsclSrXuEBUM5tV0ZRgoPwITZza6VwVrFX8GJBwvxkr6WMQkI45IhXHaNvyh
QTfpnx/JmG4Jmeo0T/QXAYqORsE02WzptJ+/gCQQB1x0NvPTS39IK7bQ83Z3JcjW9tp4ifb17LSi
dIsfe8Dx0a5fzYJ47Uz9CSMiOcC0F+ImcgJEDzwELEN6cUMM+dlSQKVuAwzobUqaQei0adln1nEh
C5dSBvY7nkdIGopU+SLb4u6iojTMO9WI3EypxiCTtuOAvfgg2fAbIDR2VzfxhJ9ralMBoskHWQZ0
XJgBxu5WWgD2k6BxdzmQi4mEF7s0ej+rb1bFBZjcacN1xU1LYqIv7bkouu17sYi9cqO7/0r6s5By
hQy8XoArXpLbshdU1dW5PbL3LXFIXAuwTxra0EO3lDLd37l6DWGlBmdmth4sEFt/B82eS56hOny3
2D91z7cH7oUCE0J9X8vb7WovguyF2Sf4/vS4q9ITrZ25sJ5PGX+F5rGx6wH4iT168LPqHW6O8+zI
QcCBdhbp1Fs5yZZo8TthoA86y4VSdXbRBDzGpJqSQ8oE/0RQ7FGzSSYEYvY8meXrPr0YKMAuq8zX
/+ys7WP4cdpz1hpeQvysXnb4eSl23JO+m1YnsUyLceRdko09oJv9hxUMZgtMmoQSeI5vkEGCOLI6
Y2bLuzG1U1No2ccErWuxYFd9m106tiGqmM5pk9p4m37ZXP0+cGymrAL/psi0eDb4R6gzF2co2SmD
baK8+AtMrUwXFQDsOxhUjxPKBtXiUI5xVmG6loFDXLdWx6lVYZJTjWQljVEtB35gYzp1h/hicwuW
n27tirLnZ1XUxZ5zNGZ1Xc3lq3T1UCnZKLdnpTRLQXyYFjCY90U0Ouw+SnBjNs9zjhHcs4/oHndF
svlv1lL9QvwERvYnUnfGIdh2ECy/SVjpyPzuGAKioyucxbci+/7n4tz5BhH7vS0FUK9Zwi7aTmj7
q+gXGHDvwgj4gwz+LqpXzENGPwTZ9+gNFnHODMq3hG3IpcJhZNDHSKQG87C3vpV2fUfr4RtZsX9l
WZTH/9a+lCYCDPG0FVrwpesHC/1NZH2HJTXKq25K7O6kiC9pTTM5O8erGeXN1iykHV7Gii0+wMRt
yD6d+XFqPlrPOX5Vbt+ELw0YAh4qyvJR1ceBX2Uh9UBl3zy1tWFPoD/N47MH4nJYUeaJcQfvKz6g
kBsmKLHqBLnmz8o6ILMEm1t/f1U8p55LYXay+cDgAzTfO70eEprRFWbeDh6n/GYljydwdkZoM4gu
OzoIytRmgrjw9ujLB6HyPrFnqcvS+fM6qWA7L52AK7GyCGqfaUJSPA4S1zwbTUex4MYNBfuBXTY+
uj1zQ3kX331nom9od/vJtPdVrpqFBFAgePe4M1AYFufmmy/sRSVgWkbFpzHS3CuVxnqvYsHrrP6X
d8CrXRSqS2do2+cNhL9B3fCg9C9UNWkT+4FIsXGYSEKfDnxMkGPQjqBDCMpwjZnQlqPykFUxd9o/
+pCDfG6VlniHzXCtl6RITq7UoebTBPC2taAsxhEPrh5hgHmM7mf94WAuLjmQOj1o3LkE7WiFH4SI
vl15GyfCoL0AlrxMCCnnNQEV+hG7/ppsBwtQKuL9jc1qSKmY9jfgVXDtJoo0+lnQQ+cjZlWHmgRK
H3OE4ONNvqlLV8KmfuOsJRVYwIyu1Wo9U3f+PpXb1ElA9aUDhXxaBUYKkTB+fYVxS+XdLfIHvRtD
XT0M7EtgAtEIT0s/5hBuIOHgF0ccZzRKUG8dlkJaFfXGx69XXA38QhdpCIfqJqgt0lv70osZl8mC
du9ZmkTPU0/HUHOgpNw0y6Z6SFWiGTu8rMc81fuy6/zw/RshqbLlnQ2Yx+gwCoQWNq2Qfaygt+gJ
1GItk1tV8XN99xHJx141OQiy5JjRvFj23UGuFv4cj7tJsVjRP2pI8NBvoojahAbTlsSmw2oEaXz1
0Ly/F3lMuVMXlKdPJhQgpledw7uLdSBuU+rS77zUKYJ/6WupWw0Qi62IMQtwpVQqPlAFrlIw/3d7
otAMNOwpWsdXgELZjNUtp87YfQ7ATTvRTXxvUZjLlsyDzIM5760XGT5BK8TBUex8prESro2+m8Zs
qRhg4vedBtkEa6FI4crKOvdxWcEcfPnFdOFKwxr/Xk0XnYtlmbtKTpvzwrHgIKIW7khLlKMmtk/2
ZIi91ndM9SiWLVLM70L3OP60Vc2GUHB6zoWTeItkUllwjxStuZT3BFpeoWAtBCfiJjguKufP+bLi
Tebyibl04V2+Y1Ud3uDU3Lmd/xdaoIr9BB/dSoOANSV45VpnDLFajkbsVGjSied2iskjcDvFY1TV
qqCeC7QjsZBGiq3YHUL+b1tKr0Nqk/KYIC23RMPipDeyoqn5qwBsOclEd5HDNbQCApGp6zu6gPYR
rUnBYl/04ltX3EJetv9ksyWsdHV8eScZvbHFyUFaAGCYS0YfrsEOzbboNcFMrD14/FXM+kz5o+w2
w2cb7WyXfB6NN2gkxztWMwBm0d3HjbHvEGpfC5DCINW+HZ5cQJu0GzEV7UVhGf9ZSRCC48v6wrzf
qwNDT6xuTLEr0APfiby8vtQhS6m/0Vdq9+G7YtVVS4uMsWwonWoDmqW8FhTFAFpXMH4yRByBFXbr
WyTMExEtWJzdFM5vsbGRZeuJux3uoLh0kNi20uWoer74i3wt3dP9lK8uxYeHtqjiNEtn07f8RrI9
DqA3jvWixasXZf9L+McFbsC8O9nmx987B1lP6UkDZSRu+dvA5f/2ZhSSl5X0ihLZ4Uap2zANuZcc
SasD8msSEA7ig2AeITeI80DHSr036pSSWCt9AXcQRu2P3O3ldBF47tRjqlndlQU/kqqQi2FMgijw
7jnVJh5kxSO/FnyMwxqeS1JH83eH+PpoUXqyyqfok5VrIgfU7ebtIllN1LTERNxBE4cDL6QKtYyU
sfbnawSvNxt7O6bHNuWUY2BwA7VpZ5eohDAQhoEBHePEPwU2OsQOyTdFONGDluTHhUud5fQ4L3Zw
iuT0VMRQzdmQ+W7Y1xXXxYVSvujzkAuViBuM72uSHOWbl/wpoKePnqdpcmIWh7JG9D3OwdhHXZat
+SE/ZwzbFwueKLv7ryJ2e9EXjLO30hNlfQqFYH1suZ4PgMJcbtoM3vu/8aVKV2abEyRxJVszxRGC
4DaJ4KPO1cIU/xbeIb0QnfQScCUk6Tr9Lk+fr7MMs+YNQCVStPSrp/pkXnisKzGVmso6hJnePDu9
WO7osorMxS1Ldqw1bhmAYrb/0rriu4ivMlFZadZ4skxRYAD/CqMAcL3z95J9BLc7D7emOyR5AfsI
4YO+8FSIxS+ik01U4KxDhVZRhbcT9nM5a+mNhpxO4a62ptETpfntJETEWyKFP9A1A5QBO5WYh3mF
VTFzgF0LJ3PfZ0arw1cfQK3UshYQO2klNP5LumI4trerCvGoBF7gd8AWMJvZvCBz11KiOSarJzmR
pp5UfOpgl+y1gVIiXdnZ2InwLzMlEAylF/XKdpGXZGXt98WerFgdb3G+MWPLiMpuA8nI0WcG9mpN
XiZ0vneFEtnm6MO0tLykSIqEHpSQRVfXZQ+Ch4ABU+llbA2uDBjkWMSB2q8ai2/3lfQ4K59RANIC
7E3dcIrxyDpKYWQ5wIyR9lp2FIpRONkeTxg8qvku03J1CCBeijI3adjaQQziUP4KR16ZAqznUuRz
YXcFpSI2iTL2X9hdowW6mNlCoMCqwKcbe05drVrz+At3xDDkdYFufaHhHXPSGYgtf4WAk2sOgpZS
HQGGZcd20Crml9r46HTGsk5Ff3NqRfDWXvg00uNIrxw1aaJlUfbSgrLvS51Ag7dJ45Oo0wFbmZcC
i1sXvrfz9m0RI5bEinsl1O1HJJhv6q9q16G3flCjt4OXkh0kHtd1NcIzsnYaoTncb2QaFzdIokG0
R49YBZXAgBPfvvBpBAFKLXSdc7vxM15N024koBnaiHCQ2F7erxmTfTK/XV0aBPg7PuGaUPwtTg4f
lgUA/a2IMz1dt5cxLcDzVbYZT9XGZkQL/chxjY8O1M/vIIV5AyUIz24dVVvuRmrhnHhAzRcPLJfj
2raAWvRM/X/2obyQZnrzj778XcGB13qGeq4S9X3rR/W72NKkGi278NrXTutPXp961qSQnH6Twwvi
1uyC6aDw7QuO3FgpkCk4p9h4eLJLWCsE+8pFKhxi33GoBQx6bKbuJlaMRYe0nB0H4Ds38CFjPUpH
KLSfJw8rl61jheQHGQUYvBFo7mH1cTzJb7HiwP24HOaKzlZmjMSK/hz7oZWLL6S2Rc8qc4s7Rp+t
VEmm0EMuFUim7+lAIA+8wfGWiPg9ghsHjYyx+wsbVofrEwgaLi7VDNu93jbclJWRPQx9ZllIc/kG
f0TeBu7DIcZ0CVcddtdFJmbAI/t1KHK7rj/dZZjr6evAVsqqF/DftqtH9mh51GvtBD2D0TP20WZb
bHTwP65XvT/YX1QIe30ogQLYhSDwE+k4DR3Vs4exsjojd8Xpk7Say5D9JXcFljRFS0Ukw4sTrdR7
XHZsjzM8w286JwW8qp83zl24c9Ib95LFU9pfUEp5aV1fIBiG5ZCzubZrgdBrTKC94Zho2ng317aw
kzWZTUp680F/9+KTgIRZ6xhHpmiN3/tSHOoOqWqZsrfno+/Etc01mJilT4Z1R+Z+zu5UV5q2vLxs
hiPobKpWywe1K3BiFYm8ifxGGUXz7mKTXIOnpVLocxBBUy9OjjVRbXxmYfnvBVmcpQSNu2xYPlWS
HngCpIrQ7tprTzRlDARRejDcNgNJfkypn8D8zvQhRo3y1whTs+adPwppQJVZvlpRvEvGi0s1PXXQ
8qpX4fqIg81aZx7IeJC8+FN0RiwWOjA7NyIAGTTznjcUeYFtMMq8Y4g6zl3Cl0AWj2jSwYpAD4sp
Lwo0e6o0UZfBzUytLx6Jp+KrpW79Ddh7PkYr2qmzoHqt8l91MfMS3W+LlnsFRBZnDzt9IVzD5D+B
YEF94I0lte2HoCfUKPnyWL0iJpkawBIadnXG0TwNCAj1+LLL4t5dH+bC+Fitrdm2L7DyeBOlvbUv
t9phqlUi4akwq+OW+L/Szk7fMce7kN9uAEyBV7MqKh5zPZCo5tgTrMB07SP8Es5m4IB34CjXtZv+
WHRjr9YnWoux3229H03E8rscTUcF7myALuOVPDixZBFp0ls+7NIpW2S9fypdf2GmTUS8G5yJGdzh
IrWha41HRa3BaeiHulgEbiOEe/j3PVUr2ydjRM4UQ6iFyRBfdiIbT6bMo2G/6aOCn7wXZodu1xN1
ei40d9EXPWi/m7gKNyBfRpZ9aWdoAV7qAvpwcEGtJtr3I0v1CwaSHxa3OwR5sSVT7L25DDnslGLs
RL9olsqPm94gDkQFisumH9FNOd4WAD+cf/iTWEULVvGfsIq3Omo809h+aE6s57BQHJP847TkqAsK
Dy3hLCVeONQBtss3CmIpafmmOh1tF9/pkO/GakMAijh8XB98T8dW6JP6QQtHWDARYRlN1RaXcfTe
4w9aKJA85n6f3S8WtHLkkCcr818qMQGrdKEmPOxrhrPZhrZpqE+nCM5zUVrzARxMBTf7XSdcDvtf
OVMZCEk/jd5/VK50mJbSlygpPXHMGupAuhwOx+XC+HOV6KDuRoTNGzTv8GV1Ieau7ZKbgVjY/bbT
dT9Wus+WwciEmm5V3dIWP+rT6qyfa+2IwuNil+wqG5TqNSHvVb3GeJtTdbyKoKX6YY348oOSaON4
z+N507uP3qIQ5fLh70vR7P/4FTEpMHsBgWMEqsVuTiM2eOywKOcbztPK67VXmOdQAp9RknPapHEK
/PRrm4ZaREedIgaOlmKMmLwm9rXttS5yoJD3bOaRkNTsflgJDFX5tWYa520LvjnTTErrnszyAz4g
OkecihcLlyUA05/814lxTYa9Eiazc5frcAtQvemgJ2pafQ7LNl3fesbX4sEHTrjPUE3J48sAAwET
GdzvMrxK5QfijwwMjdVc4p2yneIBZGGSKimfyRdOepDR0sB+1tvSa1BpQ1ReBS/7JXb4VVc/WYHq
dOJwJELlFPlF17ziEvxo1fLd0SeAydP4b5Q6IklZhfA2ckc13kDQT4tbUBOa1Lq2RrV4FAj7VOn2
GPSQDYdJfhikQjnfl2xz/mejifyelzOR/wyjinTan+AoFZvweCuS+kLL68mFM9zDKpjBZ9WF52tv
NYFsOfH3J+kdrqFYvNhkjc5CxtyjyRAEDxELRpMqqvy/RIIdPjrfmnbLGfW5NIfstg/vCjpKNQr6
en4eMDnVQLocvcRS9+XWxyLHR3EuxJHPGWEUxvEy/dRLYs4gteOLTven/R8znDtwYiT1tAVDw++1
rEx+HiTYvnRLLwG/9igc839EwT34TwGusw2zQ2+fpFwq7KuQmqhna/ij+YxZI4BRaqW8wh8Kd0ly
Rz8Reuuv02UkF+xS1iAflmWe24o4hp1/HwiGarU=
`protect end_protected

