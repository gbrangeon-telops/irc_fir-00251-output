

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MxpeY9fwU4EddFSpExWohS5o9i8UPinR6kQv/f7rVpVjW9v1XPHFNv5NQBBqnxbGk/3GroOhKYHi
zeZXd9sb8Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
genV68U/jEyVif/FXdfTRcDdNLXMaB4JkzDnEPHISJLebDAxHBqab4xQb3vzSMzS4EZxJxM3czS7
l6/Pa+/lUNH4iHFgH3/d34ImoXy9UrVsNWI4O1k56f8CO5JZkX0ENM2JUr2+jZNnrmepHCpz3pyr
N2xknPLUPWomWT5p45Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
4dyOi6X0ND7jxJKLfQYpMzBQUnXRUvqhIlWd2qdz2OgGY9VUivCAp2239OkMu2rIWSpkdV3gd8Tn
4E+XnpveIi4nHAn1AdqR2yW6qJRqYI/CpvcG8E7ZhuUiWSAPiQ/jcxRmeyzLFdVhgEV4hed5vk+9
Qi0C1DUHqDNPvc06f+xZUSTzBSqXkxyUqGIa+j3ZmCrjq04hmRDILUEkjqmR0K0TOLNdsLd81gAl
LqIfeuzK3hLcVWnnJG54RzS/q6bahPN8UaYhtJREcAC9BD1S+QEdDXRxFczj2T1LQBL5rSryR8bI
LV6YqNl+85SCCMZmZV8Io9S7fDVIrhzNm4Kcmw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PIdLn+S6alHzFt/ir7zZvMPdMeYQTL6BrWSuIGxsOazGugSdn7m2jtyII74LXXAGUQ0h11spxnUf
W/HpoHHxg6pfmAZclwmfvLsFiVi0w0hNMmIWoR8TGPdAC93Y5+aRfoAJNuDfUDfLzdBM4O7G2ZFx
YGYpvBcNhzcFFuSCCK4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KkGw0OOEdMUjhZKEmICwPPGTbEeQxk+K4HH0ah7Z5cm5dbbyDDJyn1CdBy6WY7ZD/SXDbXp0Ibi6
BH7Y9BzUsE3rhTUVWQo0OMHXc+hE0CnmrdIq6Yy3Wkf73IKl+pu+66Qo9W7SdJGNPpreGME4X4AM
zBwAv9xByRwGoY45EIIGTaE7VL15piKgLihjK8Y2Ee8q921qHsI62b9osdj+stH9M0nIgGIwpsIA
DiUOa8Naw0kRMS8QCXDqKr1fJ0jPj3cnclvP9Taz8J5tp8Sf8I6bs8irg+MGD1MgQIfeKkimA5VH
MerNz8gbn3+/Vz2X2+nKanM3LebAMLyCO8EBfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35024)
`protect data_block
iVXCcowH0097HjvwyGC/qUtYJSPNdazhd/DGKBDMNL+9hVm5hhoaKORpOthcKsPkepbj71KdikKo
uUcSBY5BDjfqq6N98/mWAnP27B4QFo2peXnv6r2iTF+j5U7DV7yA6hjJVebWusyDCJu6Ys3sDxOu
4Oe3hqiNTFwCWDiPRzoVF5u/UjphIqFjEepci9C9nBpbwVa6KikSYgl0hwK46/Qs/JzxmXH96ASU
aKQk2Z0dA9i6Nn6XKbtFow+bjcQ/uQ9NTp0//KLqbJ545ws1AQIyB5KWK21TA9Cyu5UUzYvBMmNh
/p9T27qXKBfIY5U8DxAyNz9TFNw3CSfNo37OFOoQ+Gq978C03kPOKgdOxSxeTRT4HpyBU3d1UFKU
/ivagh1uk0yCjKjjJd7PlAF8jczyS4I0jP4okT7VhCGIkAy9B0HH2um0B+5K47jYyU8Lp2Mm4axM
AcgV3B/G+MchWpLnoliWIg4LsaWlIelzAd2swSwSfRDG30IlJBoQXvElyhMHveuD1CDZDI5NSrC2
444NFUKrgR5KQ+Iit6NIdYY7uZzK3RlyntLs0tSi5lVgxcFG8eUpp/msQnCD/n/hM5sVDhttjhXT
rsSIwhkmR1Bw7wUsjze4C4K0Ta6SDOPVWGtdrJWK5kQbUp0vSrjwqSZ2mqnuM8d+7/BwwtFQb5LF
x5LU13KixdgpLvUG3OYRmBQYtHip1tf++H0/kjCDpIO87fij+fkgnxEIJl8ShOHTz3+X75IWiQrq
k2RZkv3bW2qJJ6oaZQQv/od11euLtLxuwuB+iVWIQ/AG5xlZwfuSFGzulsOlI0xom4rACGuxOrmu
F5CcThPvh0LVXJUMcCo8LTCAFwgA+o/H1rXpej8wgwWstu0lz43GenIbHhU3t2xWPSLs30E7k0ux
2Tm1FvJAgPWQW5hkBhRoLFHnxsNcdIO01bLiT11n08yaDWwvZMDAwlaDCrEb0eg/N/W88eYEBZNY
nwzvaSZG7S3gqJTf3VyE70VAffYDBpXpCUlQ1v1shCSCcA4Sxxbps4qNr2LCoTUdMSaTDqj9wvzd
ximRELcuaD12TBMw48/uPO/ewdPsKWyxmXnkROz129gll4ddeHcAePenU15PPZ/BAPejHzVcEYUH
UPjN8nnDhvbLnoQoQwLOKOKDrr27KEkW2AKMv30C6oRsg+wBt2pEcs9VHCdsmi5qGy7u6pRQUzLq
Y6+btRiB3DnW0uit1FaQLmjfFHJd6dyWncYa5DU7c71wQyorBFRgD4YxLvNYYyA0wVehMMqVOiZi
ImxTnEctf2X0yijaqAqO3SknCbZJwXy4KchT+7WuDrnm5B4WgHasEr14qX0MWKv5y/VDJrI9Ffhc
UdOkDST+lzUXu17d1G/JOU1BEMsr24xZbv2nWdmsFKxIhDIIaZMFMfdrDXWl8Gw0gUjtW+SJ3nSA
9HyNop8CIQjg6tQBUN0ShzTlzWJrL9LUA/8Mj5TKzjo7AytAdIdrzvPHn+SSeJC3YC53H7jOAMfK
sFUMUsyCfitwJTC5KE3EAkEKY8DMt+MKiPGhqHzhaU/BxuQDGUuTbTaImeUnznPYoDOYXLqvqaNF
VE8v42tzSH2/B4Nezh6J1vsaSTt8FXxVjOckA7rtvu0NEXKjQckAQY1BwRrk9xUSnwyeOEWRYkYl
0CAKTVCZ+6fSl+q3HZ+woQeFCfoWt99xJnLCGT72SecKC5Uux45aiUdsOSPNZh0AgKpJGH8clOgm
+dHI4tr4K43cHOQZnFyNVisIp92FKRyxFbHszNBeTOmWQEpsBNL4umo7y22IZJaXWOG2w0eOiU3Y
RsTOYQgog0TVC98nc0QSWa0rekb8H+KrTDCkxDif2j8rKe9r/GgFtcvO8KDGeHIBgSJP84MwC4Pp
n5jB+OaYs8K6GzJKXxuYSiozUpGQ4Q+KvwA1Q03PCG58j0+Ygerql8sE+BVWTYpcuv1BAbuKFo9c
Ke8LMc9ztUMNXtTfGhU8Cghnwmwgqn6Fz8bXf7Lh8UWfJ8QwMMnSeBCdTLy11f0GQY6G17CZOjTu
dgnDgtxuy1U0UZ1LTvsBubIBbG4DvvtDtM2cRyqVQ1z0KoCqNrD75mYTrkLmOweLqgiU4uNyEBoB
1442gPMfYy48a1uG9t3GgS8Zc0vuKxHEldA+vSmT+5Dl16OXtbeV1ubm8elPMK7eCPk0MY8kQHZa
sBcngZabcfMyAJJ1O1Jcb4porJAfperfY5SfdNYou5DEdmOKQpTTQ9KwlBQqCm/bAQMISZZesV2v
CbVIR0PmF12q+NTuQS/SI1JtRVG/NdrJOK6Ld6APWUGmTgmM8ebA52dxWrb/C/evrbrjj9L8oETC
p6tVeWT4rriF5vqOrRGIjSU6z/c3W60AQruIaEHodIi8aSvUf0QB33Aj5y8Brl9nimNW0ichYDFj
TPMidQZ9L4wrH5WJQj+VCMzkC6U3QoRdcU9EzxArxnLKHxwt0bxK9iNza976CeVyigWwd96/L+nG
vNwepUo2lnMDuoq8x/r11l69oCVMZQjQ8fM0X7WMhHMBJ86Zt/yfeUh7oWezkaClWLk3IDyIN4kK
OvaXN0uy6SdhdrGJReeckLqymfEoJrnVgPYaFvJ82TlrhR8n3u27rZfKomJv1tB7Sow1PcZna/3D
2bvmAqC+egw1RrpKY4p1wy3Cuy0pXL0RC8j5PmW0PivcwbeGDhxVNTd79gnp91tNkmbHhfqbvQAt
NpjW5ab1ygwaIJzyhQYutVVgS6uVtorDB8HaiPCdzX5YCKAEAk9r5n7WZ/h6j3j5gj+QfusM1SsY
NdhtkZj6p3dc3hO+nEUvmGCvg383Zj6HGH/Pw6mZm9WWf0F+lUaF6OVa1J+bdKySivJfqMiw1Rj/
KLjredF8ohXFp0jcZHzyMQ4j1vGXJY4AYw3NiMYrGnYZ0dP33fC22rs+MfT1D0hRAyPHC8NmqWUh
YDC6MOdbfiDSkvIqBSJrfTSxE30iR1uWrHvYJWosYmRwOY80ighHcooGkjwmZJA3GLm6Vb56GwfA
MnIBgynU7d5vc2U5ZMFJ2g3/oLPHA7hE7nIJ2zG6cD++urGq+Uj9/anqTEH6NnRPFrqXV15RTTDk
IcTqOtkO0aez+5cagWzJ8PYDhY0IER2T82OtNhI3w9BDVwlfENDCwSPGlHvHA/qEJtZEvl+cT1Jh
IVOQcxyJdBt0O4YGushZvnkLzxHkdJg7SCN59NR1p4IXfLJaeUqcBOfqfUnr0ryg+1mF1d/2slL4
F8BMlCeQaZqTcY+6Lu81BAuoV166Gm1FkrVPC5PoPvvhpRd/5uETg5jcCjPkw2kV0rhk3JrBDcW5
d0drDPfLsJEfT7JfKsHFnj9lId+WE9qjipLnTQjFHqb3ByKR9WmQBisK5GzD/ofkg4ZftpH/xvwq
m3fAEy7073DC0xvgXwvWaTv4IPGuefKy/vwIYi58+cNXjpSurvECu5DYmmUGNaJvqUmbHMOsFFi3
Vvi6ML9JekkHeGAi9Rqx2sbsHAn8cIoVKHuyw55SLBAjtVS95p8JifpFrBb7a/y+b5h1gWVqmYsD
/MjXwAZCkU6vdfj71xp27HZ+B+rJbFr2SayLCqXKFyDgJsNwW72aUgMcMs2meCXkS74wtfAVQIRY
4z/7YY1W4+8Jp5GGbev2MZj1TZLRM+pnlXZcV/ziBWMvtKdQ8qg+z0wvGtX61zwDdOoa8ic7FFX8
ydG4xSozgF1lezvKHHhdU3MN2qRkp301ii2Yuv7Uuwb+15fF3i69ejOW9snF4wDVNA8nvf1LGQNH
+aow8SqO1fg9Hz7PjNomxt1pMdqN5FbGIeGNW4FR9R7U/8q9oM0O5Qc48KNtjIYCYU+UkUdX/Xav
iuC6t1CpNw84iym8+EzG5aezqsvlV3sF7spEUMzFpoTLg0CeWeBGXpUYpNiJtMYvgSMbC7bx5dnf
kvmr+2WxHnl+Ml7n/gPiuS4kk3UyGdnikzLP1hbWYsRyYWEkoESFulQzSuyWMOKikxWpSpyj4mFU
k3FIsdGXst93pz3jtzVHKjB/M4kT/ZvPwDTZhUB6kjFHvB4gEFPXrSQLWhCds6xZ74VBFsKbhPi4
Emfz9zM1XyAJuXcnaJ2Lz5x+h8NED5xXyinQrth65QXY6flExPO2bloTWsmBD+TG84t28n6suOqr
mBEnIiRmzjQEtCq+NInYJm6eu0X3RDMqijFzUV08s14WPgoOqwzyFGUzKW3Sbyub9JVwaVWDIkOw
fRYRwCQg+2lnzQUzgbQOpMX507aKPfHWUR+MrwchtamO0a7g6hXjhbSn9fhTwDXcCbyQHBrLFfI6
17h3yzTowj8Ix81z7Cxj4G4GZ7l1VCtYoDWySPpkfAY0ZaFcQhmmHQXaIlutp1XTO80uuLmzU3mT
jUsMfpoBkTHY1LhYgFnE24s6VF0Fc8I2kbiLcm+7ewMIKnnVHEDDuR7BTi7T3nQV+VFJMmDMrtP/
Z5QSHmIIDaqMzNsVwyYJ6yZzvmf+sAl8DPo7PTTBj6ZAcopaM+r/G2x8j2qgSH3PPnXztxwRBTpG
9dwBsWer4jgjOTR1euGPH1zk4VVyfCu7vDH6uV1Qf5pIRjiWfAVGiKtfdQPYoIpClfGZnltkfe7/
qN7O3zu+oBD4vWC5IHBRxRIEwow4b5AnBGwQrMFTsj2Jko78SqzSfVY+sdYdFDAzseGCVoA3aZEv
MFwalgfFbWeIkQhlDvfCF7mdfd5P6ln8WaiboJ5TwbEQ7uBOCXX6hIhUoROVYS25ApkSnKU5RCdY
1osWOY0LkzOMJkAMKSvAg3GDoockpVJNhjpmdhMV5SeEwy4X5kMPHfGahs47f05cFWaRxW9IKXRP
bVHqln6bm6v2OKXqUUP9YIh1VYen1jyqUxqMLEIL6hmspeznDOu31v4gxPipOpFqALS/785FKogE
VLW6bLjyalh2UHY5+QB15JK/c8+HauyoRHEtJuzKsFQTQwN2Jvg04xUVtwdvasjNzXyp5sBZQAau
sxYrfozyk2k9TtKHRZjyVLswlHvCr1tWzys8c/ZK0iT+hooaEAsv0sMsKW49GfM/knHD6tPd25bP
rCvBkoxk9Uv1PJzRQBi+7bek8uoRahqub2CkxaZosvWTEMIK+ka3QTjnqpsIpHYqCOuI86Oa4Tug
s+gUb8gUldPTyChBjpOqoCKAN7OHHTd6404Ev4vPDVBorSlTcCTi+m1lLGXL9jXym75wp/uUqYEw
4kHUSh+JPbGfjg0Wk9oZE5w+9SRwx/3BTRf6w7bSt/E4yf3PROu78l/8E+MAleSesQ3lW9Lhu9GT
PQlak0afg/cnq5Ing+DPsrkRoZWqP7CieP3spEFcULJE4+ajCSdw36o6BbII6mf4Ga1RNMksSbpI
BqVNI43e0y4W/VurFAW2j7ADbaLDYZu0xnaDqehBPec1eM4cw83Sxp0wuQEe4x51EzSwj8aiQmEm
VwszTCAxsiMqVyhA3ouZknu5LCM4me8vckxndz9aokc+ELo/57KLJGIibwuGeXbaz2RtWE9tOgTR
eraPDYLp0x0FtPhfC9d+qhXqMp7af4OHX+s9VtCabKtzZeZJQzc1EsmlF99uRfGdvP/ldhMMRMNM
mzFiRd/gPlU0JoViff+/lbI3bXItonhhjiC4Fzl5Lpam7igB88TatUwJFVATMYJ9yPXbka2A4Qvq
c1pNS+dTwN3IxnAiHHFy0syk5sbTBvyu2/f88aetMb7dU2dHWy6qnhS3lgim0zrkcMly86ziVBIc
ioqYMJavo+SSqcVylc+rwX9I4SCy2tP2mT+onhRu8t/xMF5KHwh5E8OSwMOx8mxyIkSZnDbIrB9L
XmiZOGZVJzE95+7PL2Msm1k4hUCAbIHd5OvO+nV3Y6RB0AM2QgKO4E0i78zPlQkFfdbdbY72Gh5e
DDlAQ9DNX60x6I5yoYPHya495CWsvNOuQr0YVROTWx4h4Q7FGF1nwm3A0dbIO843UVcqzW5jvjTe
AE2exvlyuF4yWVFxoiQ4ToulosFDF933+aNImW/rsSPclJRHdUFT0bH/QtQD5UNpiaTIgAtD1PgQ
EMhpnVAIHdVO699d2feKsuVswOkJUxhYSuJTOQWyc+H/pdiBShV05tXKFaQliiZVmSqzstz9vk5z
SV4PIZoXxgo+z9i+tuQ6cE10xMyq1yJczSn62tKQW4UFLu2l4pKtd54pNXVbpLEO1IC+Fku8Y58n
oJJ4ovReErQ8l8HEuiuI2jx6FNhLPJ1duvfXQIPhgjOCZlZHf/V6EIvhZgP4p9dHGDsaxwC/aIbg
Er/md5yK5cEfqCgwaESp8bcWEw42oOwIoK4Bfog5KR5rhM+neWRyCVyKtsXut+RioX8+g2kQ7HOh
jAJz+8V+uBtv4a0OTYEZBduVVJFAMPyRZNgE9a17PyEuW+AjCQkybW7JQaUaM9gG2GSeSrF7YNTm
73bwI1Im9QhQqPiyhqp37tX4ZzVHMZgj5g7tgyHmNRBDWzuIdm+5eIzIHtu5imJj3vSEnd75SsQU
5TC9i8C/IMVFu4C3SEehrbolpou09klBZpLL7odWJ5DITR/N+T9XMgpc/TN3EfkWFJlkNBNd81Hv
jfB3/gKSmscUoDV8t1icesCjh1oiQwtoAR0CX3QBghO/L5CLFztWeeAzg9LSOH3xvOtjSaE0PVd0
R6eFS5MqB6McJn5aXsbQN6Wy6LhL7zm3h8EYXi9bXbjHpgwP6p+T+Ike7hPD3jpHQ7n9VGmefQW8
LW+NJPWbRnwbulp0Tfw8RY9+oQPuOxCp3VyHY68C+8J1kNc6Q/6YgYGFLf6HYbNCmnlNv3wfoRBC
bdirDYfA0Oj8wSl2dnkBIcfjcoISFOIRlwUJHsLdi7MdcxZHDAMZ6e++g8GsCogsFXyOKdJgHbpv
ewtYYMFfxXwP8XoqYOLJcgqinKVxRQP46hItoPz6SzCiq4N5jwxj7XQ0bRHvnCiRg9C1DN9+vwAD
E/nqchO3hsYXWVE4tcWQ0bQuYgqULNA4IGRSTMmDBEy6ehvWTyVFuZp7b6U4lyvsapWtgiT+dBSN
uLSBknn/8XhNlm367ooeLz5ide7BkAefZOLFNkXj69GSuXqfWFTKf+KC7nXGMeRF51E28ChcZAwE
nGA2SVfrEgj1uEtfO5Hs6eUTYaDAkEiYg48/cbEJomwJIHW0f4LdZfpg4lvRt5hZNPxPUhHaKM3e
0Z5z2WHMnxQgsy8uY+6nzsdvpDSl6pvwYXN748tejxZVGanbAJ0+A3IXDhBPaPav/U0pYc+gYPST
bfxc3nQs49xnvs5uCL919iJm4gNh5JP7aFNalcENMPB5VK6GL9N/vcy63Gc39PgYWratxeJY/ZtN
H1e/+6fYCA+1gfa239MRWmHRO7VKBpNfzd6Cw9WklxURVSedHrJj3d4E7OBWywy4Kd3gZ41m5+uS
+1KobdDHKiFHussktypFuhoTe8HNUhd+JeTWRvjlhMAbTQRBU2LrNuWvymXkQlt4oqaDF5dtSoeG
8yLeIUMDwjPJKnT4loRhpVNTKBAzs3POkod+5Ct0t3vmgqdEx0CrR8NjTf9Y+9mP5eHZ5n5hzEVy
QXyw/8UgYBT1BLNt4HgDL7U86Diq32cp326J4tT3TjksdVilSPNBZ7EOkOwbwFDvjsHdV4Gz2WSq
ZSK44PSnNWHv3NyhIdB5PXSouymeJxbd+WYbortO4cWLTPoUAS4UpkCRVEYzA029IPz7clHUjjxA
t7L2d1s4nOuu9XbpbJKpmoWyPiYZx5yzkqq/m1l5G4nbKOFTLIf0hj0w9iVReSu7JAagnAT9A1Ay
8qogN6koC77958EzUAWQMxKZLTdzNty2FiyM2jjVkkI4l0jGI/H52ABWiAH1JtDbvwljvJ4AgB0r
F1ANfjUeC+PiIY80MccZbRkUd2dNP2xFF6n5GbbFThypAfKjFH26WuO9SY9GADu7sTdmOT276YB/
ADOP4hHF6cKtC2+Swrne0H+mjMwO2a3QQUNbc5Ok8dh9zknvDfatBZu14FZnyDW7V6oHxeD7B9Y5
4bkKIcaLKxRSifI5aPhcMjAq09fGC2ogYS/WOMoctL1fbhbpbk98auSxFF5V14Bk/3jqkl0yHA8O
wkPX2d/dcEItunrSeTPA5rrEECu0v29g1OpQUng89cn6LtGnoKf6HiKdBFWe9qFoXbnp2vNMY89M
G6KhjO20jZZPKj64530pUBpTWp5dQSpYSYqbC80VjVYHzritedRu9QsLEb97GXVCOR6JpBFeGn8R
BTdBOK/PLvcIRTlkFtNK7IkKbiq+LDmnr2g3oh40ywEwYY0hw4mtN/u+c4+uspxeTHcslX8Q31PH
Y6REKeYgX9vfxwzb7pic5UjH2NIOo580LcbBVAi0TzM7Mi71Jm9cmt6wxcTEFF+Qu88WGbDf/vOi
S25EVPT1zGhsfvTEaaZZmwPf6XpMBI+6no5UoCYM8Y7NUsYN7t3rfPICd/60EAEQViwm2gqxTRvd
HCQcN4ik2hl8ddGWhq5PHLOxXtmXtHss/hEXYfe8QaWPHIX4uffCLkGO94DmWLkMn8TGHrquShmA
GVPbelFG/kIU20Opgz56fO4a+gs64gkX3b2CqqobzjmoOnmRbUc0LBNE7EvGsA/Zfnxv1f0yN73M
2z/O+kZYGQXJMR4bRTwktIGI6ZmUhWKG3ZPW7TM64UsxaNCR+3tO6KHuZuL9pu6hLWY4Gcl+M+Ps
cV5YSCKNn/80C5F08vXMHPa6b1akLllnKHstFFm6O3iJZikm2rVszummyzm7TvkXt1ZGxmPQlasA
axcqpcJ5zWANPuJA7pFUWuHD8hpeylt+Lu2h4qBxSvGK70iMOHFnrCrYiwZDqJIPsR7j66QW5qIT
FtpdLvLxwl7+HTkDS7iQk/EequFpvcFz/5hMF3JqVqdf22WVoX0uV2R/45uRnLKHa6ayOG8aQkQI
xOA5P1dT09ToGoyckJ0AGbQh86e+3wGnR4FxYN7PcaTPREoVTvH9/SxEqCEwriAe/Dq3MVDCQtfm
xlCkNJY1caAmE7Q4qAwmEdy+yIJbP1ulLIzsd2qzjXaWsUkRVTk2f3JHD8uxtQKX0PLGAaJoe61P
Ixs47R9xwv9nDs7zZrf4/zwbVpzifJ469Kb2k7FmuC2kEtXepyuhUImgumzy5L/+XUQ6NKMvXtdW
gnKK0lsBKqpXQWqG53iljZc09vzULixqCE6jLLUI/47ebfwMEtAlO5yNBsb5VrnaoLkwDeaodvz6
Fzxf75M0EVuEdJ8QqcIsB/CGQWd2/YZQD0GH6rz288goqdZLHkp5coR7KjLkYSYl8JQXrSmh8HYk
R/oXZDu6sGc4ekhmHkLxkTDMXYT56suuHWG7FCsXg2EaDvnkirF4x/THTQoqGXhVxnavi08oyZp8
9QZ9aIvLgeAcVpnlzP4dzAze3LdFe4GzJ6M0yoMW8a1o7WHRjZ98aZW7u09TVniJRDLSt5Tleca1
Jrxp6jakwRtDrfhmBoUkG6p+Gkjr4eJyCSzHUxhzIv+dsv/nS3sKYjM5ihN8+5n5TXtTVao9SB08
HEgHzNNEqopxZdS2gesFU1aCa4buxixMHj9qq95H+1LrSEmwAaVHVvYvqMJkolT3ixeFCOVPUIKT
NBO2CtjT/FoPxLTr9CskPrKKAubSLVaHRJINOtoNFi5kbvtR85TuEwZJTUbWiQZ3aUoR41CNGbUE
NycjdXt4mTo/tQMVs1AJfwtkgfcULfvwkPGkl3+dhZmYxpVZkdPmTqe5zhGrOh7FqpO+W72fFQmg
sXALYCc2q6P9rCnUJRETZVRX0/HNMgj7EobtzNbmhS/mmVPs7yp/VqpsiMTtdU59qR7pQcC7lHwp
Uc9iuU0WEI/NEly4L+nlNz/eSTI1PvGZjDl8JMogixpo4RUzKRHbZ0x2mYuqIDz2ggsD/q2MjTkh
40Hp2i6qRNMqSXZAfinXfp/NWktoCEEUL2eHQXIVQ7sZSBpBCN0R7k/AfmRevyu9W/AcHhf1e30k
MsA4sUvAz8B5e/yGyTQsW3hYXv1qFMeKUfVmCjY55JuLTH6G8DorI4SoZz0Fgo85rN81JOEpHiRm
/2gXxLEGU0fc9borwDqsrcku+xdhy3ELnCMuvdsZDrBj23k1AsgaKvLou1IGYeK3GNhSW2eJe63z
KMuJsIiwQLi0wm/TRa/HKY3NBVFrKYQS0mGKGkRh9rLarYj/ZF3OghwLye3nceERlK8Ix6fF7jBk
n2DdcKPcNmipbETCnFxnbSWt4TZElYKnAMUmQnh7l3bXNqUdj0M/XbTwztr0O3XlKTqd0xAhu9Dk
/BE1ASPgvsgLYEz+e7WthpuOLMkdVcmsNf34EZ6PFEDoFAIi1lDICrKfSw0JcvnYB8LqdjgdkUtA
rjDxUCSgRz3/xv4XviIBFpCKnBdjJA8P+dzUACei2YLR6z5XlmBersobiVtQpNPsnxBFc4FODLRg
L2avgiIDmCEZEcjCl1YUUPNlbeWwSFHD/E/GWAXnbKUupMxAOduXGZoXW5DrpzVDezMzNzBVcRxE
PY3tbv+7g4vEJcuSJbZh7qTK8esXOOL4D680bv+UGiodp4SpSqYwBJNWkPcqsDVCG9m+O56xsy0F
Rze50H85IylJsai/Az3lJg/D1YmF2n98Yd+EScrbeohWOjRHZ7qFCw1/pgukGPQNn0R0YN9Jersb
b0EmCpbbFAueoqyMa+RUBR1qpPI7Seth/8JlbfwvqEGm0/R6BxGJKkLg5JxjhywZS9YNDXT8Zd43
oEE1XkQhUSRw/4oteZE1gfZMm9yKTSHc1YSVuuYle2iZS/vF2o6Y/5bBFRXsaoL2xKRe3XdV+6IE
kTJE/xA9Y+7rzJ2i3u0rNv9C9LrPrG0CBc8OlcGSEhsE3pEKSo30ZiEpNjkDN8TEhEMiVHyCrnsi
jytGN1ZnIf3zPeCvZX/ZkAtuZA87e1oxc0U5JdnFdTvy8d+Pg2oi8CJC/hHjUaMNVTsR2GQSa5cL
KHRV1xuOmIRDJlO0BlMBZOhqzbD8UiY6GoAWFagThHy9olBTufaonPkQkTe60+5fBkBfTHfkYDCM
EsQbAZToEQohArK2/XQ11jiL3ltLdG0OTdME4wVGL6IxnZesV3+DyoT1JfsSiXE5JM6bVsoVw4Qw
L1PNxgkDRVzj5FEhhgGyPlDUo4Z3Q9Bpn1/ux4w7HPQpXN3BXlcH2HQu2RA4eSRR3b4jfN19NC6J
StNleKq7BhE6PtI7dAHfwG9gMn7u9xP3ULZznAbb09s7GagOhNpnvSoYoOT0hG0ZG4F3Dm7F52HX
zbNJKFvyO8Yq7UHKLSjlPKqZK66NP1CvGo1aY7RQj0+yMVkKuWAZATEahIc+Y73F7z28zeZxbnCt
BabPwwRMcku5x4EMcRNcs6No9W1dsK3mSAqTfmylbneJgPaOx4tnRssCFLn7VOhR/irxG2WRxr3y
8QqClSDNz2uXZsM8LCtrHOIc9aHlv38DlNlMe1eujyL54yzFbRFp1++PwBe1uQsyVzBaQspA0LUX
CbomTVX0XVb22crMgSb95L0MAdQNANR5wYYSljGrc5ec4CvLGj1mq7JARdfPxzdNAikSu1IOgeBv
2P+jWVEd3KPN2T2zSm1flS9b1+rbhS7+ShBCe+93Jw8U4+/zT2pX26oGNZqa9O6rhsQC1O7oLNmT
HipvPDdOQDQ4eThQGrFJUIlgefXno+yLDrpLtdKLlyWy5Hje6/X8+8FwBHr4yYyvG4plQHXrQhVC
LDBTBhblBz9r9zeI+rDHsHcjPYpwXJibmRSu5/PfAMUbLjqXl02MntR/JpgI8/3DgkzCNleVRn7O
Sbd0HufDE7DUqPTvJL0IozFtRb1P9ZXahPYWbwNoRa5YAfdU2zSd/xRHgRaJP803Kkp+Ry/bBDcb
ccUYmiFXu9Dt2teEVkSWnzoEd6qwBfK6A2iegajdb60IYow/IB/uWV4+l10k0zXiiP8UItF6IS1J
cnUZO6JctFRDuzXhFJp68inDPkees/m4APc3vkitS7AEQPi9+Qou/Qjzdap0gg6vb7Y8Suq06PyW
+uVnA1b94DFCX59O5hhl/kGFsI1K1gIoB2ShXS4PhRBQ2TmnXjhOUCjFB7MZCuKlenBnfcb+Xl9/
kEcNsf8YKpucTLo/wY5zaP3xLHDjc+748srp43SswXHjXS8fTT/Plve+3V8MykDQm+x/00/Ewg6A
WZUfUDSzfXGGdzwpuQoPKSFM3dgtyYFB/cByVq7h/lmzauKbEV3Nga4kycw0PWeD2zbrMcYGD86T
3OglL1cQG/hYmi0izt2qrFCfgpNU30avxgdRPMrYPj3uCk8cwJGEJqiMyEttUkJdBrm5xSKRFvDz
4Ee96GTzHZ85Q9+GqFU0ouGCM9RjCFWT/zyVOXCdGHy0EvjTSYmY/3b6TJ3wsIjM8r41ewkRLi4l
KeNPB3px4pOoSE8Ihvgpa76RgCXbxIL0fj9ADoDq4rFmYLV+2p/ZwwdKfhUt37qQty1CBjayKfFD
5h0zTp1uXLvs60wbgnRlFxbQFllR1V7gNSqvlkHrQ21q7u36m5PIbuTAhVo1AUp+P+rfU50dR0Gl
o2VSz0tqNMlihz5F1WifVQ9xPxXFJ8QffWAmOZzhJsaJyFsIDXDaygQJd1V4nDAE7gca/dJHQ2di
GL+aFuZTqOd6faeKn9FSf8Vyxs+2msO9AdFTfk5NK2aHE35+su0GalCCmbV+i4q8H0mCoS1Yg4eZ
+pdzKQK/8CLDletnwZ+c3OSAkgB4rSWcPjk+Zvoy17d2kr23qcvJLX+KE3w0tEHvaYNKAwRKXeHu
Xv7AmtGJ1926yu1Ft1XVaJHukQl52LOB0nrJamPn58r0jav4bFafMP/3HWE6zwevVRceplumFYcW
RTV3tytyq28T/VcUoQdpOuE+O70rSKrm0vxtTY6h78w1uce7Ut0qDtpZV4t6JjnmNVXUmnXGd3ak
jRFy7s3hewnMODedsWY/xT7SlS3XCW8/9Kp3jIgBKbZV7+dJwVvOyYLbrlEhEBCyJzeM/SFZilkq
JkCxPkMTNDVFASzw5/qNcSd5ho7SuExsQfWilwVEoXvyo6rdf/se3+IO4T1m1FXgnDxcOegjJHwy
NVGiQ34KI2k1LiEIOGBXm/kuSHvUEa3zE+DmtqZSi5S6NoeHSyHiG7PkMjctn1NG9KyqppartHOR
qqPp8VxDg5+9Xg97SUhRPyfFasjk+25DyIfOitYm7qtH+95iAfv/g010j+GOn6XGAvkl/j8UV9h5
Eh7iRlN5mYNOd/bvYQmtOe35GNhpphID+rII566OFtJLgp9p6XbSz6xA1QdMTZp3GgQ5oGzrfXn3
OY6y12uowZirHxp55hNwtkRJ8+1znVG1Z2Gyy24Gxdu2DlwC4Whi+hF9mmvOVeVoh5aNJ6BqkU0M
VteBxnW3KFMsfWPwQvmJq887daXzKc5Wp8h2ZEz9NUjgX5vLLbp5RzAN11Sl3Pvy+vb1PM0esRQj
+uFf8DfLDEJvq2CWKmYggVPTkybi4eoR2rSP3DI89j8SpzmbhnAFy8US+wS6CP/+p45sDY1lRmSX
7EG2gVg1ELJ3nEdj7IIBqLyGgsgNOQjysLk5HuPxd8CwIZeZ0N/XdeOFoNHcVYHHP2PCXiND/JKI
xZtrHHDZ0289rrgvCjkPxsq1s1ZZym1d4DSAaoViTGkbyIdfq+ZLe9NIQ7/s70zH60tKlAPOCkVl
cGxpdooXAb8hJyTYE5Zvv+9Nl0bD7NzxKjE0CD5CZQLuU3VZ6QJ1BaCxWX/MPm3qZNNjxMLZUo3D
YKM7V7k60OCGGFdk6cD7Y90YsuU86wXMcY+0S8cueaYeW6wzTy7dT54DAu9XOLhRaOuOKimYYcAl
a0wlogcCIK/KNJImQCGj4SnHAUIAeOXqKoKq3b7S/nPVmeQgJz88XfSa3/1EoftgR6Fe+iBE6dtM
/tsBwaWjuDqNOzWR/IHACPySx6ViNXZwk8e/AlueRSMZYoUBmafF9/AnccYU6OCcOtFkOLyKjeg/
4OpriXcMnytTRiMjUMPGOglYcIasTVGmHTowTXjv4k6U79WiwY8uRx+Asq2FRFPnkZXxgVQ4Qno5
jF22L/05bGoGoODByinf5AHN373sgsu29hd1FG/nT7R3GgIS+BOAKiqo6Izy5OX3EyEkO5lo0S97
iXkpABIDZvE3mgy3w7hedcOQjsKc16U1KNf7X7P9YuD3UiE0huh4VRrWEgqznGLWG/eaMdbjoRlZ
quwYVGmq82L5dlojUB9xET2n4knilq0WTQpV+5CLy3fVSOX9iuMO5h1ihYYmlj73Yp0PpTf5wMen
X5J+GCkNHMTC6O0cwblGcniLn5g+RgTjYs5Xj8e/IfLrdb5sRPwQPlOb6IEq5+VnDFbG5AFW8k1W
9ia2qDlj51nGyjWZH7kJoOveXketlC4HUUmNMDSrD/WtEtmHubEfeSMwBQCCU7hbKpJN08l2pQs4
C0pJdAQEGWiYJ2xz37s0pPtv0xoQCC6+Z2jP3QixuUYMu3dRBUAumZmNz6aX6ca7ICjtNtYrg/uN
Pz853QcgL9ZYR8n4tUDWeASiO5V+vTweuyCJnWXOMBkyd52NJ13DbkONTD+IjcXj+GfIV2wYDCt5
+X50G3HICH+IZF9oPFw913FjK/TyT6Q320+beg4d9twD84YCVNsYo+35b0CB6gS6ZmKaW21LNRhD
qj6g0YJOsjMFUTQ9eOUwW5Lcu1cXYDTdeJnpglf2IAxb/yE1FbYiZyNz1xKJKdyuRwmTj6ZqozQP
Rrs6KjMfnWx/vd0VFQyeIVzBpTd23ZJDx+JnTvgfqYeUOR1oQh+8fDZ7DIf2oICnHmRTAYHWXeTw
1x/nxpEdyozFVhUwqNSyWSJBQc79vCXnYWb14Dm+q01oQbOkiWNvmJsXpwyeS581E+Eo8vhb5wdx
hnNWyhc8Ovve9YRAoa+kHFoTWqEhBf7koslbt70urD1KVeLe1PBjB9jpwsNTPD6u9CDFiJYfPUSW
fun+8XO86P+xx+Z6ZmUy9mkXVlvxgoUDmggYETXnRsHyRfSucLoHku64mOVG1h1yJltb7DEO2W28
u6/0rnieMlr7efq2jam7pqxvKvlYB0tQaUwQV9DxbWmYFJSqffoZSDHfxh+4OL41pOxkxOjzhj2K
HKCV6jdZobe1KN/BellHZd6jf6dQZ10dZWjayoSw48fbCYGg88+s3e3pX+KpCQIsbPLG8R/pmvoS
YlE9jr7RMTnq1IfE2gIlRQRW8k0BT1fwtcKW3cbFYzfFDC28vLpfu+DHtprafBs64L4P9bJ3nDfY
JgF57qAt9ch5joeK/kgImRI06S46Y36KhpWJBVDXlduuZPnU85ELexOF4nyqduML7+IdFgY+X2Em
/wrRxLkfL0nHvom09geQ9b1gtI0SaGchllbUWObmIjUCnKoEvEL9YPeJG1OvC5dE6IDUO9mZI6+x
pzSe7hmvuN1kdAv2/CXsPP6GygXY6X1vMixoLGzOJOkpkAIF9oah/lDy9MsCTOMdM5wGuS9LiKbP
MuHVYBu/NXvGuUb+BxF3YQEtiyHL9tGUycOwqyEB9hq8lwVRYhmOK2+fkwPdcij2naa+6eeQVxMW
fFCVN9SDgi+SgeZJGsHplkNXM2XKblTAW9m+JHEWNv88bIiECrE3yFA+JylxmuXXMk65Pc13ujt4
9zAh1J3qu3HfQ8pYuLHa9fguO9bgHtNRzSWQ22dbx8cx0gQ/BgCJfhBqIVvfTOsiYj5tW2LiCeXn
lmHBIdCeHLcJLJz0rYcCB6RsmT5P2+ZC17leTgWM88cc11TQb9/6K2bSJkyMpBxhnHC6MHC9b0u7
5ItlSTuG6M8MaL+/bJ3bSSkrKUpMXOKbzMp3l/cdTrZUNlydJoCzWoxdXJYvMhb+GOt4NbVjdbnB
70n+kgEjdXP67w+U8vv3diUe8RqQpAR+hlhwsrpuJ0IqO6A8ePLN8/SazzpxHHOmXPDlrehusDKS
/4/WFC9AcBViJhlytOxXI3C0Tv4O+WATBSJdRWccuHo4rjIZy/dlBcToigNnhO3qT3xgvI82u6S0
xCIjsQDO8jPcEHK+Q5VlHAPyPYcx1eU23wT6cbHE4eXuneQxZNNx54M2/nj2Wk/F8p4J9+Zt6R4Y
fqQedGPIAuar6qT5dDZq0BBV5TVGugZib5Hv7NegISxSWnv79RZNogbiTn1CbTpPWx3/OzcTMyIY
ZcjZK2/ZV/5IWplgQNuIUcArtovT+uR3zXjXZOlxnHzYcho9dwFQBfbMR/t1sN/LULrDV0WXIqlO
Mcxb1evA+f55MFdpKQ3DOrkB0+K5+W2O3m1dCpocssvpD6nUIBonDpSmclRAzN3z0n2De0wmWkLH
NpCWpEUVbD4o6E8LP2MCvLivZiyx82B7ByczOy5ypLBmryL8LgeUsFFnkH9Dz4C5I+G7wakYvGZ/
RW+BkMZZdNxqK5c5FHDOhROgsgBFbUEXTxW4wgTGJKY4y1Nse59RSAGyzrFeRKwVtskUZpDX7tNl
xruktB5TPv4I6lBond2vdsDpfIC42dA7RouNGYkwfoIICinSC1ChUkSch+k7lfsXybjxhbMIy4GF
DcTZjHGkmhsoY07irKWA7sXnURAr49P1IpmE9B/fPO3CWknmqa1X4X+Vu1pmOtyLEc9Cpusk5kOY
ZC4mk+XB8Ag8PgX59FLtVvX3f0CDSjWSri8Xg1ILrX0XQ1w2nl4P11HizyOd39CXgDOh3d+CeD2V
pQkTqhsalkQf2Ra/T3P8wYsKv7VRKj/IPWwEAWktXh1HVyr/mblWiTRn03AdBWdYScDR26zVoMWN
YagY6v9URsR6+NxQQ1t3zLTEY0byp/bMsH0lvqjvMicS3CUVxPIy1lk8WTRlbdNv4QKvfOoSkXx6
wVyadFZoLqulQAwf6NunT1NcYZE9c5jeATH+tdLRcp6VieJRREHw0Z5RiEUVroKXJj/t6Nlqfnp4
kDYzTRa7Tjo1wK6WrUU5hHhmrrlfIRH6sDKOf4n+CkQWiJvRVp7tRkzJNPLRv/YRptEtJkt0uugp
W5QBvP7UMusoHjzgpUe6S4P4sScEVqNM5IOglTylSszbOgLjx6KSdEaq2IcIh18qw8UMZqzlWyzP
199eBPJC4mxvq6hb/F6gBA6XYLpbUYMj/GsZm5yxJHL28EOWBNUOBztIiuoMO3ly6G9Ib7U72fk1
quNrBQtUozlU3GIK7JMbGleXlIsNFeny7zO18lm5yd0lIZ9t/57YNKod9SJOclOwcecNjDlEeljI
Cqdm2/qj4JtcRNsa0wiufqq+zvNhuM84NMbo3GphjHqeE6FD+GDKH2bppfSY2mzYlLnf3xjzRe6x
dXYQbN79bFQIZR9fl+7drBPVVTM5wr9NuFgNoa0ZHHLhqh/JW3d42dSa08JdCcEjkQ5l18qk/S5J
oysBglfDGX6AVljF55NBPu3kqKJToircZayWptPKDJ7z5Plh+ObW1IhyUlkT5Cf2BlRlC5N7SQyO
fiaTGYGqJOXV8VyMVdFHXPToKZmWUJNIsNdRN6ze8gMGczBOHpkj1SCy2XP6eWaVVIn/3fpCO7qr
PeTpXN+m8eeqnBPuG7dSL/g+1UPgWUlSSWcpDql1bPD+GxQS8PjBzfKC5TARqAtLfDA8zwhI656n
W3iFYhjMhClhy4PnsSK7CnlPGpHFi4cDLsDyHepxjgY5kPZiSaw57dURDGW4tqv7OL6lWUtD8GsE
JtTRwl+3b35HPnkR+V80m7mHaFFTe6wCtUDz97FttnypBKhGaPHEy8cqafFRdPUcYOzFl6xRfqjC
r2y/jMj1yb0Ux60I4OjEEyElYU2EkODyjUq9nv9FtFkEB274XNH5gAb1M2z0uOTGE86EYadQqvpG
aLV7juUEKLXR3zwt44lqZecmfDVgepwg6mRSj+XEXJ3Sw7bkVeZIKeslQrj9xB28pu0MZKWhzwsz
7u4JwLESxhFaxJJotJ1sH7hrGkkbNK4Ym5x5AG1Mv8Ehh9e2taekgStI/HMuHbKpnI7Np+UhHpTJ
nT+OwajYh6HXtypSLahMlarnh0Ki2v7euBhHltwKKsSDlbUkzClF8aFZWfl3jwUjjNHPgc6/O+1F
QnCFZHnQifvzFRp2tBds//e8bUxJClP9xTCc1d9sD6Dj0wmVw9TB7QcSKOQ6oNhMXvwBUTtEDExZ
4AcK+T27sIfevE3dTP7WJmsmVx0oxgBCoI5AUlsvZx76IZfrXmbLDrsjEMKEwN3k1GK+LnssuhZe
9Qok8x9eYgqep8BGJHLOc1bieWuNzGVk8bH8LV7jrjZDmHZLSgNAOF0Xqud2nxdTC6FuquhPlIiA
0nteaq/UhESChcrIS6Yb3N3qlLT4+qtXUjJyLULyyUof8ux8QQpejnxNjQKdKEnTEBMqWMcgIIkn
tZrRqsb++HF+SIiM+vacDdvdKNndBKC4rq5RlruxMPUfwUQpidOicIOSq9nzkWy4a6ywLwRt7gJu
15I6F41HREYYPqDdEf03M5WpadslUgF5g04V9WPs+rhNsCNe2kbkxeWVvlmCu70G+dAVXKxHkCfr
yvx89tA7oi0UQSnMJu4YDQK6xMzqsfxq3UsUnw6BW7F0ivkwHGQcFQXZCUmnauVnZK8/fPFEcCZ8
mM02+dU8RLWyYLTM5pAxdsINbXmF2+aunR8m5PW5FB0JSqbyWGwzL6KNX8n/ubrVNAhBE+K8c1PO
OzJcnxTZwTFjRx6oj+MfSWlcCpuIwtoKtINfcqALVrB7DOkRH8xqDAEJvDhgQ8hua1yZK/4wJSyQ
1SK89GEjk57cF1YKjd/3V+J6TchQy0P7zjkyJbeew3/4jCxUqooiIEzO1nUVLT3z2OctkT8FVe1L
qi6HPaJMillRZA//VgM9vwFPc/EhaV1aXPiUqJXq6aiRSJrKglA5yeA+MClao9WeVSkEyCc0ALAO
fJXZD5MnfhXYpodVV6pCmQ76qweOYDvtY5fsgfwUs3rAY3nA+o0PA0frjL51jLGrVbKYgYBHYvvR
dGge+enPo+XL/gWXRE89rjlzrQPbuPZY8RAHksxoqk0UBkei4CmLWqOx6ZnmQTG+jBNBgRfBDItB
gFf5I+og+ZxKQRgWBBL9ysEARpcpCvonSLto+7eTXdMpajE/G7dGEmDnY0gy4cKaHf7LklqcsS4j
eY1A74hKNSAEGbZDOqRBzjbgUTeyWB/Xi0QHVJkD5rSija21yLLHtNHORfMcSPIgNq50+6j2Prlg
ej3gEnpZBoLikgWR6aG47wwKLYu0zmIHavX2tt5+ZMYrLB/dRSuzirbeiPubdqNuCrHZV03uWfGH
bVUJRi/nu6/9wZp603/nOlH58sGtwTEGvmJzS/4QwK36CGw+8TR9P0jIBkOPrWpwRSlTip1C57jE
DXv18+cvyx3Uyc4AgttKXFe8l+oBOH6fEyRrrwTGOwgj0eTOpuaVefUhp6AC7Y+fS3u5kt3hQh3G
anAQl+sviuI9Ii0MwH1FeM/hAXgW4RiSLa+M6N5jxbbU+CsBPN9KDQTedqPC0lQz09BDiBw8tlhX
KTqU+whBKP0UK95rOIZdd1ix4JmZJ73jauSB8bBbTiXGkYNcZmzk7wKALBgYFW6Js18WufeinK1/
XmxIxJv2dpF0Lf8F3kkeNRpusXkiF86dkkCL+3ncBIOQAFU4Pd42WlMldD3z2KD96JdWQeXti5uE
fh1sOi6AFXYT+kCG96IzhhBE5gOIZw67JqcgJXphi2aPWM6LxagIYeEmChfXhwvoXUeZ3JC18nvL
l9MWcpfVBghFeTawZhQVwGsacHlqlJSFPEQ7MTn5Q6soZMW3XDrdWC0exhaPCfeX2yb/0eiCGcOa
LOWX6H6kJBrMJ1J/GZQDG5LsaQfhSzNkRj8XVH7XQJbUwDKxJzivEtIclMNaqfl7mXW3pIYYkI7I
Dnch39kvdt/Tm8W594t3msfEtpoJgQEkClV9sKXmlUWbpqkxTlPdADHpOdi4hBfUXdKPvl9kFd2c
Pp2ah8/LqOGHeBcB4yAGLdbOcAukrNUIGD0F1UeINK31yQpUbMPkYof8WpdH4+aEQb2K8WbO+5nt
8pGtiWZxdcmarQWjFuZnbgo/c9VJfMAT+wcXKi2YQw+3uyrgGc3+VXCsucrA6Ow/62MfB68wA5wx
aLGrinNfrywZlX0VWbOfulmdC9ieFDEa+DtEYRKyjqQc5amnadYKYoX8LAmHykAM7zSeRCdMPsLf
ATQ2XXjKNwDX8MNzK1QUYoh+iRO9qMPcYue7DW34bhvdlclVvMHXCp3+QlzMhF5kawlpdYYMC6WK
1SBURzopyyo8/G9DD1OJQhGMsdQ372W3UPs5701Yk7rDoYprOGXJQL0AeSiKEaJwJsr+tSLb/9+B
Gwyp1f1vuFycxWj3f/K8YL6CuQeV8XYYVVvIPtr6Efhtc27dLYdxOg/m65CbxaUk+sBW7O/30i5C
AdzweqI9otbpiQmNyKlJzQ0L+c32HzEAI446tNqzwad0GFvs/ordz5gjIhd3C4TYHS7KgyTCmTXQ
SmpvgtQn0cIirLdciowUo+lgtdTGrFVifrwSVeQpvd6XykbFguaF1PWaIufyOlLe4DmnLB/jaAgF
LO8+V+07hBvudyuRXaV2rqqZoLWn5I9xGhoO94coiQZPiDGmDiwE3MGk58hd7GzNycdiLN2yi/PA
gF48SGUmN8fpkJmgY3XMqNheUFWqiDM/8OVYj5/8c75+9HsL09NYSQ7Obr1WgZ1gIvz9iX7fPxXd
ud9CsOtWhgtNTHZRr7XImGlrQZXZbIJ/dmAdVBRb1cV8KiPeaNnervGOowDAydHBoCotiOOHVech
R+tubIZTRNDOmpQkg25ISnaRuUo+PpRHCHFNYkPrDJ7oR8hQ66HocoA3DIYPcbh6vXeBbfrG2VUI
gJ546lsw7xclAIduwxBmGU5EDG6sI8M0E6moFU4k8cugqYil0AYE9uEPQOHDZ5jTYUUHDl9Wj0jE
rGVVkvivLT7va6vAXuQD5PQIIYFzKKDFBjExFIfgQ2uXn3WTNmk+gkjHnww0+N8YpvsojcD3P0od
orn2YROkdiohNz3XNv/aorlZB4TeMOWi1DZGdbgJUqnEE7fUbrDVpLz9S7sITvJXLUnmirt74Jc1
SbkKMbkLL8rGQfnAfJOdojAC+JQSIQQoUI986F1lLwMpFR5h2MmiiiWLDsQyXWttqI4/stLWt7yF
DOuvNxH7orN01EyTkPIBrJ4UnJzy+mlMguzc9AWVqDnxuYWgI+meuWVCEoTELG++kOJSJTdYqSF8
4ujKN2tedw4LdlrKzNloTE5vULCr42BXsGBw28CYRAG+sxnj33W7PPH8V3o7WXPZospulXaLSf3e
mlm4sdJTM1BrcuFbVKxAdOxJXnzjOudWr3CqHbmhi72hUt0/RlUucXUDL4j16VCvAKi2KQh5YcTV
4sKwKF48EgBwJaE/5sOmYhn4QcUGZ5AmlXLblL/NLia3rYBiSCDD5Bvw8x92cwClXel+ehqr6U0q
8RqfZF2RsNjIbpvwEpZqdUNVLnZ8r0kOrPDVKleTqfPoWBOf1VaQ6Orj14pPHk/HDDuA07a7ZkOC
XGmCXHk1YaQGohHEdN9ny67CZmTl2uQs6F5srxwJrvPDJ+mqzcxUkznC3id8pc2D1B5z+RTAStHD
I7ol+vxef+Gj3Ct54OMelBzHbxC1qG4PpTL9zAHl2OM205Rf+smP7hV9oQ9KGXVpDtyZYgBGd7jb
7kMB2XwBd5pXojCHVPAUsqikp+PZ/HeubyU02auSNUOX7J9Eh19KNtCl9vWNY5Lf49zvET4B/rLZ
vIsnZ4g1wT+Ki+xoxLaPTJ9+SdxjRrXDxDW09TaGk8kXajT8l0K2znpMXP6qftN/u/84tT6TM2Bx
AFncuPddY4nZ/eEHlCi2SgX2bQGEgOjv7PlkncleQtPyNxR5XLlddM3Db1H1vWoHtOc5Rp1c+EDl
i1sxr4gTGJuNpUGB6/mgg5GTCoJCh7tEDo5vyZyzdWXfhcZgOojqEYz/jggY34yZanOlB0Y6AOmX
cxyJ52AD1u8qUqXm6ymCuK4n1diXlOO3Q+HNNv0kjWNXEEFK3izeeBav0hg0sUSmelMX+8fOb5uE
2+UonqaPuZ/GGRKGZNBi5joJpbHw5DG+VA3NqZHtK5PzuSTIZZVN4v+MIvgvtxme929CI4iawFJp
MITWITm3m7NnTsNvIA5AIBAbsFcQAxjy0FD4gPwX5XfxSy95HHnq01bVKptbYmBt/LQjFRMyQIG0
/nd0GZqcTvAVKyFCSpcnvgbsUQofuSIrHUfAnT+etj/713O//j5LByEh5YmLx700Y3hKPP4BRaom
rqyexLfcZh90znzJqdnWUs0ksSYowSrn7ZYjpy4sUiEiutUYwRLdEl9Vpeg8dosz6RXqxhnqxiIa
nQVDTaEM0nH92GueSGv8JXMvuurt96JcSaRd/SBRhvKlALjRWpIqPYHPqt2cEduMad5rElanaYlP
QO0POW7YKej95DeEham5ILSMP39ErIB5DBZxW/8ffxVlCuZUKbJMuCIQ5u/TUkQKF9o8Bo8GD2wp
iDyDI8Mhig/bhf+bXBK+nrdExSvFyTd3sUPYVoTzpXqmBs8D44EVm1RA5ooZaM/1oSLrBGaSRE4o
7ptHgwCCbnvfOb8GKGoy3QUmrVhb2dKmvS2FtvI95ij5T+jJulF90yyVOQHm4sw608CyUxUmHxGU
faF1n7omTM1Bhp3OjqnYPivMJOq51SnJePmCO3w1kGIG/tJ5xv9pAPPcEAOSbFNJI4mGAQ/c2vUq
cuWJCUxl/RXLmBXY/0BhX/zVH4u+8+e5JeXtEp1G1B98FrQPYxFm9CnouevRZs+FdPIwKNVSH6w1
wsqjWwqNFeVavA1LgPyqcJPjS3HHwaV0qpa4vgLD0q/ki44WMvcR71F9E21WqMUhEc41P7w7m4ZB
FoRYSzahEkzrOti3M2LGW564C9wTBmO3hPfLc3UKz9ETfCLXZDew1Fk46J+4ZGDPtPR4i+dCfofp
xKvRKoR9L0OMk+KKPTCHOrkEFG0BHcQXUTWbTLhm4yeXCRLsdE3ufffipnynENGXmihhdr2WRRgJ
vb9kn2R0nAxBT0rCbfCMjD1B4HcGGhx/EFT8Y7gsS96J0xs6dkoQvnjDxHe9AtlGIVYO4Bso8vnX
7Sms4WoR7syWxRrpQE/YY1v39kKHWxothDA2uERXefw/lCyJNhJ/Wj2sE3NFgqWOD+vzq4gLMzVz
rMC9p88ArLwY1BE4/0Y2JxhZ0oR0QnBb3DmNnWpZUT1ARrF2TIJHdNV6K3DHPb449Du8ne02tdzt
57GJXaIgeUbm89n9YNz8kOus10nwkVEtLsiI7TZsKuH4YVFjI2WKBHnN0o4bG8dnLRGoxlIRxbM8
SJ78wHJBc6v1AAuWd3KfEwdZ2PV/vUW9FkhpbYaxII3SOydXxTV6dsxr+/iY/d4pC2D9DD+9KrIz
G8ZEkIU+Wo4Gt4jEQfMRw40Z9qWsLqlZCzuljNFxFG5AmUKSc+JyPLyyXyHl9NI3JUqVoaaxuO8a
d3OpKGXwDwwnA5022D1GRYkC+nKeO/yYzs7LLvKb6cfwlZfoHU5PL57FewLjNR7DKErfXrI512wt
+Oi5/QJknkRSJysj1Bg9N5hBN7YjN+RRG/S65Y41arzD1aov2fhBCLpJCUfzzeSL/P36KWaGiK8/
8tOOkYgRPdNHw69s4FGiv8OIzsmhnNpOCY7aT4ZIFibiLxg1trLjMJJGZt04SdDTiOWlEbRkx1Zj
Y6LmM1/HIM49Z0xcxkU9Zm/6bNNMyd7NE7ycq/q9oPGA15r/EarrSy4CEyOwM0/ANp3kxiQulDew
UNqbefhdGhUQ5TBramxbS/UbGPULORiQ3NrMi7illYOow7J+zi9mVk0lq4bhjb6jHjSkx3mtVvUU
DE9JhKf9DMUZRnTVKf6SFCRzuBwMwvrMTrzspIoO7gdTfApAcrvq68XGUFVYcUS/HhU6M/MISdXp
KgFZwZOcUoCYxHc4fjRMtRLlLLSjpW7cuVEZBcSrPM4bv2v6/xf5CYFOAVCIZNtn/t07TN9hqP4L
P/HXmdhi1mvnJtsE9bOk6gJLOI/alvMG6X/qCaGglJcLiyhj/3wEOXrAWeNpSbV1pve9sAVDOK3i
0HdlGvQjq9MrRw83w3aSaQNSuPPze5+FCMWgDYTpYdYXNq4R1bYmNOvyjPXA2b7ZTv8rNlOplSHH
sc+Y/O133Qv2xSI0ZBffPShjSkNnG4/kap0Z6il9/CehJo2UtD3RpERRRV/b+6ergKj1UIIyFz+T
eNyzuP93zt2Xjd5JtyhZE/TcXFS+1QaFLhZDJXXyckT3JmaXW7aD7qw3QHAK3TQKLWX9+5IHOWA1
JdgcezrLFjIUdl5Sz9PkEmhfWpFtHPpCzTMVLfmeX/s2t6zsJ+PcvSFL5mIrxRcGbkU9wYOlpjqE
Do4D0QilT3hLlDDXA9WmEiiiSWu/Jx4mard/kzSFp8XiBKrBMofrMH0mTT6Xa9WmUAKHyYqVtxA9
uIEjWi/skmrHvAcqtEJm5EWKtyZw5LnCwnyMj96fuZF0Sv4P9THsQu33jur7ssq+2U/WoFeulzwg
SKxtboSNTokBUkHEkbd2AIAUompFlbFUsmv4SxHO+cJU8Ym3uw3b4ehRj9GOKjKoTLnXJg6CV7Iy
Ysw2VL9be/0htZ9pDe89KQuBWh5+i6PfvuKKhuJScxToB7I9kEQgvkZC0qiQ4X3S5u45zlgDrQIw
lg+gOD9HaIKMo9UjZJJOrNVvjGZPR75MNc6FLTKXW6z5DzAGM+gprF1YhcVYy9vdirfzYX8ca5Wt
T6ot6s9rsfebYpYUrGhe7NjmQ24dVuTCSiHELVU0SFmk40XZDiRQsOND5SHcYK3jMMczIQofu5Nk
sktu+0hSOvQQ4mNAoC5zqqKrlAaB3p/EjfyZTTqqbirr3ZV3p4kF+/S8MPQhoFIiSwA3hT3tZXsz
xPQ4YvJ5agR4H/1JzkTRNwD17/7VEBhZwQ999iXt8M8aBuqoeOjQpwkI1BZAzFiGF4RDKn1Gus5C
3vRNXmpraO1uih3LCnwpESacTOBUYs48V79rdHQvOzZPKVPRiO0hhpOZ/p/98zsW7gBnBBLtWWvr
iOyYOC80cCFOC4ybsQGK3BAWbIWOLy73Ley55gpbZbD8Z2Z7X1xZCGZrMoCYBlzgpiKhfXainXoh
zLlXOKlu0KV0c+IQr42XBwQeF+M6nfKni6NuH4JxVqcV3eoZcwBnytBw7cAJ3OOZRXnosO7IxuR9
nSN1qPeGw5opakJ/E561yp51fcI1syN0UHmU1yVayhye7WPIzlPUW+8awYYBHfngEDLjXzfQfpHu
oFND34lbDAW8SxHdTkFTDNIMUbfeFgZ10Pfc/J6EfNA3kN/kZirXsFaxwr/PLXDzj08et/oHR25M
Z1z8MKEgQfLO6IPRYjQn/UjUDX1BfkcqAozqbP4D85HxuFEGpzsCL5KfrgVHsFMVrb3E+UDMbGVb
OWmi9vutUrNJM78E6gItCRlkUHXk9ulGD3dkURko06mEB4krgh+eKjuvfsDY/7ZJBa4aLXEZ6uNQ
Qzp7+Qx4pl2Y+gPUdbGOd8E42Osw/BJCH+RspRXkARbzPLoOtx6iktPRx+R0j/wTS3ao/tmvSPr5
eHnZboVyOjtn6bWmlw7C+X3eH0A6fxn3ccRCEjfVZ0fDERu5gLAvqNfnvN2GtQmk1yUSL1289KfJ
CHyZfH97mOexQDc8RmCL6HmPzrdmbhFgYmX14F+4ie1iV5AoyL2cf2fNnhCuexXcg3on8DuWxnoG
kPtrtyBv+hxIIEtM4NFWtHRZviSqD2YzRD4//IXdzBQbpaiitAMrm4T1AUkCs5uyV3YJ90VA1rry
vfDvpuJcFNQrWbAIw/uU6ATkW9KyPJoBN0buZx5dGV3YjIFjnxMmSC0+Bunzv8XmYjK6WLBfVAZL
FTUzyM5Vdzcp7xoVOD5RGyY6EJ+836mWCllsHy7DaEMvuQsPTi8sP0R4eemLiLeDvc9tRaWvj3a4
cSAceJy07O+dphcnPEtYh3XQcQg+NbEDBZmdKheuT26Emj3NSFNUdPZr8+17RIpm17MZ7Ko6Z5mt
3N6KUt6HJbHLUdXGSV6iknwRGodY8Hx9rHoXUkZeuBEOypwRCqiZ9V//MS58rXIJ1c2JDCzW4jNw
Ad7GjqMp/v/9W+IMAnW7KaYjZWtCdwOFufWVSjC1sjHwOfI9ZHn7/JQTmTEBmqEbIkea5uG36aKK
Mu8fZ/oaQ+RxsskuVx4fk7qoffELzl/B+DGsHwUdbKkFpBXkkizj3RUOpAN9zzbJkerGqcsI3VwN
KpRNjrkG9DDRG8QrZz09SvAzEUnCz+yu+UB23LkFHbKQA4/8wLByaKEyDs4iGFqXsB8S/VzRNBBF
qIit8jdS7/awT8UfxtaheinEsbqNJfFDBIxKwrN9pAgi5vYqWCumRdMSCSB1tPU42MPLBGrH2XMX
/68fVAU+Zp9FW7UagnRPbDiigQbCe9IeDYGKEHW3+SrXFIGkTuvrNaPy3z/Y/2ze4uPVHSSkbcio
5EY3ZMbbSQyya+tWc6YGMOPfAc9PnR2dSX/sVStK78xPao3CPPSlQF5LcLmOzKQdgPvRgM2aYOvP
M3jYUChWSel5okJFyUgXd7So7H3wgq6KAOdMYjvM9xgo9Y8HiCHiXfM13BiDmnlSvWd/4i6bbm4P
JSWdx5nH1P4sOKJsCaMlSz2vsvYwCVF8NMWzbq6zg6QN8gZOqR/EHbeJFCaVEhFml49o1oUugda1
4jdWqN0UDoEDC2NesOHPsNfWpyd53gh8RSZrCm/L/5Cn7MLJ1MuQi5dYfDKguYbXCiEEDm5UgcCF
dD9IT23ZZwVRFQyROoDCse0eN022clm+E15tSGwkDRsCZ1qQ1lW5Od8v2S+fy6DM4cnuimMnRxwP
GWV6NXqS8YfofpEhgQ+HbX6JTvvNOYEJQANMZqxFZihcAbAva6XwnMYGDjSYuxedJ7Wx5UKwSnum
xt44NVQMp0USRCGB/CuYemFVEEAVdrTNWCN0zUMB6ANDcevqItRZmB0Zxfs/DGS6ocEUk57wM4pA
VUfhgMdKNPPp65H2ASDR4r+bmA05x/zQSPWrA5iM7zXtHBwqBXYuxXJyyixXYH9H+0Mlr4DMzgTy
NRzWjZgizftUtT1rJv8QfXMi6qjhE2tlFbfZZAdRxjCGnZwRGPpTIn6Av0+eqQseFE1QO0RPycHN
C7lvt98e0rf6E4gJ6BnrbfqiKeGE3sRUSW9fEkroVPN/K46ylI0Nw1Aw+euB8kjFaPdUlGxj8dSh
3I1hJ4mAfZJFipgEOaCFlN5FS78UGF5xKxuJwLHBIGaZMmQU1IkvVuWkflm9iMTEdTWMTMA0kzeX
dRV4avgM19lh8gUfbdgi6FXhWfu0EqNIEzbTb9axt7lZCu0rO74ciO0GBGj/aoT0HfyyjW7cumr8
Tcm3Jw5O07zp+DdmpUfc+WHyCNgTCD21zjdAt/8DsXiMvO5K6+snVuDq0+pDxuL6AKwF6r+lanqu
needVst1gg8MMILz9xTPVVvG0R2xA6gpHLCTXkxgd5VdT5jnRrtXzXUbAM+tdrDZEGZxLlBq45Va
/PaBgF9pa5adislgbrcv6YshMt+nFiVEYJ8GRt7DOiBhbx4h0O2l4ehMAMVbus1qvVrlkIob4MWz
amRVm2W3bSNxDPzPWDVTgr8fKAl2WXb55DriqrNWLXZFtKI45reBHtOpQn8+EXZBR/68NqFaTyw0
eZT7N/KUZYRXoBs8MNkkKRD+d8cPCO35glhqNGBp2kdG4198dwegf77kjo2y5fw4Wn42sw4fp/bs
o5l29bZTWIMy72e0r8h0Hk4PLtzJNY938anFwFqzajTJ2pqKGFMqn7YzZh4y3Rdj4SEMa+EuJXBT
1sgEfRR2Yma+Njq2AkRtQ9IakjeOfXB5ZLABXmXsfz7xvRErAt9+a7VPBEo2P3dMGyIyYirZt7hy
4QyZOR3joJvpcVGJTjtHPge93pP/mOOlurTfGllPz/3z14nla5jmwcNbiTT0ZbqmkeijvHHWYEB2
eNFGkCN1FSQSIJOs4XJjNrS2liVWBi2sgaZoY5EyIksPTeI0vt+Kf4MG/4KUi/T2KDisItnj8NZL
+HdDYFPQLI3fp5lKUHRX9pFdLAEKi5ffPiNjN8cnV/LAEtS2ptptn0QPTwW5V1OFDZkwKb7DSxIb
Ar+Zx7tKBfn8N7oGIUYC8qdONBG05WNCmOrt+RAlLnjr/1TxLbmap1mUGavi/hdYlUsjMwbz0M2D
qQWU5i7scs/JtjWXQsDi/XMfN50T2uVQGYLuIenK65brZOmrqlWNj3Ijdhkb41L5qAqiiRr4vYN9
eRH3egIRz+y44tgFqTOCMVjJPHH4vWJmQVQIartrliS/3cLaSiBZuUz8e3G0/pdYOzghcZbLLx+b
2gMQSRMQ6Phv2hLveRqDOD9im7dWvUTv4u/e5PS5oRb/Xcgb1P2hU5YLKWlGMFsxjjMozilfQrgL
8c9sYih758lmwHwo5onGGpam1DVR3H8+Ufwnntuo/jd5sn87Jum4VW1HwMg4y1ORPAXjt3fQSdYL
DYnik23TvHUwrPLWyiGWKll+L+zhagI0J7JRUCpDYXFXPAecP5H1nNj5Lxv6DhKCgnwj9shzrMAv
+fkfcw2Cmd8cwfIyJp/KloisE+R2AzxTVhT3a0iGSWiKbs4SiGYnHEytqDSUbXar8y5iCcFKE52q
VYaDOtj9sQq/GoEY0A/WDTBHJkH8Dif/jxJqAnmS6sOSuvdmX9nJjF3qpKobNcvgqoFAwcc0eIa2
UFIaINQGSZu5ryntJ5J3AvOcBjf0+rB8pfGYBYJS1bfFnpiKoqDIBzZrsPM4ptBRt/T0Ulwn76wf
ttumlLIktq1VkEeADGGDjKvHxRuxmbcuiAX0Nq25QJvLdfcvZG8Zb0BwKV6A76vGNdJJzVTCW1V9
oSmwdqz7lf/+9D8d2mt6OY/oNjnvnuCh3VVxHuKv2MPtCrNpBzsR7oOix49d+3iePYfFPJG0Rf75
wODVD96LYboXJb9QymwSI9341yjR+OHKYEPKrMCZ5xqB8J+uqVZLWcYkiIV8LeIIZRjdVcwhKR/V
2CF5FsCnQb0Hws+BbOONXsbznT+eSMa1tgpH7Utxk7S9HNYGPGZEzeXJS/jxsLvTBeK5QlJPo86B
n7bxJpLv/PK3Qi9QqNAWjG9DQFO4et+FAZRKhPjBSfNcjb7q3SLnT5d4F/2rXvPO/TtBDQ6zWWwi
sJSueo9o2FK7nmx8m6oCldQdbVi4NZsD3/mqgV0wKg1drA2EBqWAYNnNu5azvN8wtwPVmdB9xf3n
gMsx/UHHtv2pJbqIifT9J94qzfLxDCk0HpcxZ3aKm9kkTG4sTnydTX5070kfupP2XjSLnSOomkub
IjtAVJ8+xb8HSIElZfXdZsEkEEeMOPGtggX/rxRayoVmtepvL/iKvtPQ61wD9Smx6NgW3QS7RyiJ
Po+StBRE8kuPh7NHyz+42liw017DNz+0ydL+PD3lhj5IoSMbXjLD8H0ep9l01O9vimUklM6NKYrV
PTs196hv3jCfUI4j4o5BmnFY2N2ncGjgA/UWR9til8T+pqq2qMpo51/quxtYFI7Fk17mLOksa8/V
6Un23+vDtYNE9osnVK8cn+k1hT+tkDLqg4TxtHvsHI7kj8axKBYVMbimsjSOVRYomY9n0aauRpkd
U92e5JH9Ag5hD0F4oOEL7gTfm3hxQOok0PG9P/ux54s7dHxoaBvx//eGUypH2SEIH2dVlspku8OT
FFEZXEBv8t1GinIRudjTtL474xqxDAzbKkzqfrt7dKltPjxQuASOUzb5yo/hWjvErt6JJnOXtnH9
CotGtUEvMrGypyjzREK5G+6Q/mjqbfKhxstC9l/ZUOxjjoumuLn+RXW5faigP8uFxp3vz0FlJZ6A
cLuT/PL7xZo/qtQnsRYjFyMDf0XD1eALHIAl3CM0CH8ZDzb6nk/9w/IEKGYzbGymOquZRWcPPLaG
g9H551xd5Vi/ngtG2TywPVTFTIL+FCVfJlHA5ZAfs30e5q7lrAaEd77V9LbDbsgEhpkX4tRyWxbP
yNFN87ijSMZLZtTMaLRSyz8vGNv+vvsy4LYnkUpImpNz4/q32up37MQLGCbEY4tE3P2HFzu/LUz7
saT2YjCWzyyQRf03FOuH6hrSy1wwqbILsTExW+ACTQ+pwcJfbEq7xTocr7rGZP5vtRk/WJm0wPSs
KJOdUcZtpdtBUl0JLKfWd4Rrma3dZdoa9xmU1XuX2ljEyvqdgprf4kv9Wt17/VNg4UPdyB0n0/E5
SHQ84K7kj+Tr5yx+unBgpJyjQ6YDhyJXPfon2rqv2n8uB8zluKWhWAcE923VEbfUs3KPLec/gXAF
ngsDqSinOSAvvmNd63NO9wMANfOAFpHHT5d6q50RUYw3KN1nVLdAef7K3ODbdHrEFvNap5LLZ/DR
7Xh7oWhPjTLxmlaYsafE40nHJ47XEUI6f4kuVZKfIKqvzscMTeVipaWCZ0m/lTUS5nZqxRTg8Lv6
s512bjyKGKm5w4+f/boeoG7jBKVfgm1VJYd9SCx2zU8eEJnv8b4W7u9OoF2LfWILc8ZMgr/mNTVP
Ux7dxpdBNI+NTIau0Ogj4iPevo15YX+ET7eZHEcX/fwXawZuYoS66UBC69tCfozCFkvSvr7OF5iD
OFVUJWeWm5EMEc0jV0xZN+ozvC3ZXl8aKWoe7opGDPzW/IglK2yr6NY+3GJaVIqjQ+f+JPBQy6Cs
Ho0VzrRhkdb/V981VA2NyLCP5amZ7St5elKqx3ZgTRVT/Krrb8clPfTF9wd/tIW8P+4gy++UhP3X
xPck1CDViBv/FFL+d9cu7hAV0wLiatzNomgc1KjDVQXoF6oMLWlcagBldUmjA5qKC5iQGdXgfkQn
iaYPdwHptsgJlGh65EzuZIMPmhSoHBEdQQ8e7Hlk8qrQN7/8ghazyDhhaA77NoQ0UoBl2x6lrz+9
TZb64cHfJ94bmdmUH1wsO1IqIJAwUXOeGL77j8Pe2X4thHlHYaKJvV7lVb0KOGQzRNEQCGiNwPAE
dg9P0ApT7WPgwqWv0Q13DeL28OwEK5wWAdiMNNTJYqKeyy46afr4AOKdiLjwkPAw3jdPhY/UbTtD
bk113A5mg10IyKxGYCCc4FKdeUCcZR20hxUs96PZYraelplBOPiYbW5pK2VS5UlPbl8Cv+9ISBPb
fH1XDACMHs1TBweFYSY2FJhBK4zUiDpd9f3MDeamMMPakcMMFmtl5NfnCx+O12YQg98xiM9hhqw6
oLMAiBtIn3eWqveNGdamwp0SV7gHPTzJiPxwYLoWBYfFlDg+g1TDyJt9/lLsQjuLpwhpBc53R90W
nj5RhUCZT4UvZ+Gw9sJoJUmsBv59D1+/s18j+fFpbd5vaHT+sB+dwgbogJasepiwFqGCMRh6V1Um
ATD5IWYPx5YTCHMqvM9Wc4NiEFT1ijnpX0WuT8MshBDsJTG6imZn7lJhcyj8X+12ZfVLzrp3SJrp
NHO0iPIqkhuGT7fGsxmBBj54BHYr5Zrns4uSoXgzEtjtbj+BcYjdE5sEhSAX4aHefDp4fZJpV9sY
RzhLS5a9AustoKU7TImgjkxrocSqpOxxLmwNvfSB1+/Aa9nmrhCsc6qcFEB5kymgzizX5quFTDuA
GUEmui7l1oVAHrgoduxiU5veelRkUXsXpHqADpR3b+tVB4R8KVxT12FfVZe+FfRbzHzQ8BDI0tCT
BvsClDWNEMbcqUKlQPlPnjjXtBTs8fCSzEuDdQj9sRskcQ4leJjduEXQEvU6Vk+KEb8lMKMzxD8e
tCMCEubDjfpyNtomhiNhG55uq1snIzR34VUyv/QvzxkDODz1DOV0TGmXwZMKCI05vv7ZbHYhT+pI
H5NX8aJ0oVMdh12ChV3HQJluhnqezbKDyY1FshwTzfbI6m2wuy3nO/ISp7o0lXGFClMFhbFpFk8v
6dzlnROENqKgKVKUlSXXKFE4ERQ61fo4z0PojvdUCrA+6kVZmM5AqZt/6Yzafam5Me50NNANOthH
wKCiEyKu77xVxv6lhyUmKqr6yknl0Yp0YsgQzv4Y4nHsn7h9V9oj0YTw1l1njS6O+EX84HQBEXXL
DDHS3UOPEUVetPcGkdImda/NeBAE9AacDCrcA62a9CH3YPYlgwL6dl2MItQ7IeYNoJTi749IvtKr
LebpkIhXrV1+IoPjUknhh0W0C47WImCVJctycPlWXcowP3OOMRD4ImkIng596441TDblGLKUWBa3
kziUR6/oQPNjbk1JwFDXNhV/zMFQvj9Rn4H+ZrUWSalKmMxjU0Eq8vligkoe2EfSuWrtLTXpJ7th
PuGmjlh8HwDTuc9P56zp+vJ4aRkcT/nY6NrLbAv//eXooy3ffBViRNWQHEe8KBfXgYZezEvGeWRa
Y6Mk7jyu2LwoefPqTFZNzLrKdLUVSrDCcVfP1C3Po3LtT3YNabi5FriDTBlRRZocXijUZAtjQW/I
lT3s5/7/Ai42QRTHchDlt32K3doFQzr5GDxre3qav9FNOHnjZ6bIMNcueyLpPUM4oUoX1h77/ORs
4+tpSJhE3zG/0dXv7pR8dzBh3X27EhjL81v3eYGRxpLULbtwWkiytrr003vilEuPx7cTfd3Tzbss
5IptGOCwQpUzB4Y+cDrEq+L3ljtoUWXK+aNDqlnuWd9AMxwirZfErzlAh3FmYDDVapSM9xSLoPCi
AAz2Bmpd9HCFlvzo0jBSJXqTLqSwTeNgJR9j4EBZiQbotGu1EyAqCNPHTBSS7qU7Gg3BllqNU+dv
+tKmvHoZePt0k7bTlrIjuJWi8KBzECF0Pyrb7MKpb24gAk5VVeDzLPElqbodBj6QMY+Tq14ecXPV
tu+Og919KunREL0NhVHnnHHh/Zkh26fHmZP3E3+GUjV87ayx/4C57M/y+dZKuCAhBYyecat3HxFZ
STdBot9443pLfBvkEH4q36CGe5wd1JU7bGzw+F9WiAG1mn0yl7WZekDkGTHzui+Dog1cDLyWv0FI
Op4rmz/EvvHimoX1XCv11rtma4l1hOepxzIn83Gw8ODyP6JMuu0cpx/ZemdAmpZ6SZGqmspKGGC2
YJJtLQ64NYUn8HG7kd0HhAoySkGCA5Ldvy8Zku760uojthWJ3jckT0wknnozLNtChFddMnvcNUaC
rj72BabaaObLPAFE994VtFM6askoXLCtUKe64ZbvW32443hk7d/b4hjO9zXF5tz5KX5gAaPN1KDN
UuzoVmDcav7BH5vvGx9p5Gc9UT7LHHg+3JGh9mqyvhjuPug8X2PcO5SsAkGan6kjXdKORmBstXy5
JzidGpaLWNXMuwT7NPU5wkIIOjbr/0CRLQRvIPvcRnDkaxzny3SEtQ78CTJS0b3+RavK3AEJNps/
L5U3tjR3mCoEvEtR9a9s/ceFEvDlv8qjbeJFBDEnmZ7W4K9Haw7pBKuoQPASeKWgXKXcS4HzajfE
q1f7STpWCXRvduzLZ7s9hXZ/bo81iIOVRTS7yMqWqyHvj0UMjw/K1riYA0uBeDUIMuldzjU9LvWG
1Y9vK7G6rN+Yte4yDeUel/KIs9xBGlhNotWa1Yqpab8UOLNwnofMwnw1yzogVsPYltIs//hfBJIH
AGWe+xbmXz0JvGy4vHOS2970UIdFUD1s3fsvSW8bVYpDj6e9V/C3Eig9tgVl4pMt9bNc3CTni2LP
f4dhhYIZMsgbG9g/wtT4uOmpxan3orlP/xj+K5Iiym4K1tOoHYq5V43fVEn9R0Ud7kVaLdZaepod
4qraTstT7++YemJit7aD5yAN5ofJcdbJtdw/Lvh/DI2SAcfyNfbOZjTy0tGj3N0OJw/mKBSGKQEH
aUXuLOYwbzr3JmYBewH3AOnTmX2On2KuG9YMj6AJO5BhauRkhte56Az28lGqRD4Trs4kXD3Q0yBH
aF+zcyxlocZqpcVPiPE0GLaUdi9KU2Yas8ofXZG6D/UdQTIT41Tel/aF55ttUgdspwFDt3cpDLuS
8HZNHoJCJ4GRYgQgSoZDC+7QjqYF5tn2yLzhVj5i3pbKa+dBqnnRbnGYehy65xVzZ8el3cg6A0l2
V/yxiYqu3HPnTqcQhaHTwR/9FJOYIgaAbuyQX8XEmR+8fZU+2KZZyJYDb2k+VqXS7aF0UHKb6iO3
ZyXqh3hPMEqnKXeK0aa1wP9WOskJPPDK/D9hG1uAU9qMnD1334kVefzvFzOuG5FBtnorG7ZIf4QB
txU0zlGmEzVkVLHcqnfWgCQnlzLoYqPJE/G6L9Me5u05G3npNJR2QSVzhULUDraDzcSat2ZtAY47
aBmVG7wC29jnl+NpyA6f1akMgx7A8Sil/o+rbQKYrFBULD0Dou9YZBMbYskx2ka1eyoRDMymYxo6
63j0vjgkiIOEl0YF8KtNM7H23GvFDw2LdXflN1QzZQ942DQlANX1YPCFkgMyC/dFV/qScmVHZo2o
RqLlxWkobaeEpKxEvwEBB+n1imvwsp+JAMUK2eP6zTjLKkt+kvmRgRXIu8njEQEjk7VlcHnQiarV
MT6gHzgI3EMGcWP6PnkYP/AnsVnSPwtTaXhAF3M78SxUxEkpEOmd8e5u1nwDUBVsaw4F9y0QPtFy
nmk/cgLsF8bMXQmbKzJlq+8pGYELvRf1/ZQAdyvp+2x4x3xqu2QC9aNHH/5tBU3MWdSGPQva9QRQ
Sws2Hr9fbT+Bl/9usxuZIF3q4IMj1KliY+sMYrGSgN5lACDKxNhdmgG44aYok6m13CBIdn1H7Cvn
i7apb0CJaK3tXsGAKwYkbHRsFpgwYUYAJHLRQp6zv5bIXbcUfxkeQVmEOPKJcaHb2msSKA60ypym
655t39x0mFmWJfDkb9FaOdhq+wzTwbdTf71kLY+zS3mAIf5m9p/VOuxzCYY7lzTL/KzxQjlOaKlg
XFUcmioABYoaJpYWGvAV3ADzkW+v76iswFsiMxl5ctWp8uC044cX1HQvIhjjLJTsxiuyPtKjGCfj
cnPPwSpDO6npDPQKnUI8vugvLLd/u30PNwxRZ8O9RPstlBVYLV1JlJcJCivoej5E83eEPGA6BPEz
juJg6lWFttV50AVjniDtiqMBLqxzavp9doBXvbw2jclxVZzw0l4WpfuxhA/9/f7zJ7AjKxBJgJA2
bMRcXJBWBnNz3RjySSXnK/WurvjuTazAq77M2Ib+3UaDzwVsVBxcbYfTM/AHM2APr1Het70dC2o+
zHHG1ryZ1H+XzCqiHWRtvG5n7XYQLwR/X12kaaByprDVGUvHysU3Tp30SW3lLXoLh4OayYhAZ/wh
JHRX0Gsmx1feVqwcy6hIMjAE+3bm4AzA569aCrDkZsPJARtMFgJmMiZs6A2Jp0z6uCdOYWTK9/qG
YfBl5n094iBXhHEP9DSwN4gIUxb4TNv7Wa7Lm/Q27wdPErlQ3v2R5KRAnlcLaxsKJTilMiC7tQCz
V2ooydzrpX+ddNh2agmU1jI6Jg+2KchRVrZD7jwNRAJtK3PLNPBb8dYA2HxvlGE0V4g3VhvnL0Vl
6dPauRJ1+UqRF0Lj38HK5XIVWqZarqoiOm7nkBrGmsbmEJvLgW70prHF4vAtbVGUovdKIMzTxbp6
+Uso83FZF/C+u4aHG6DktPwgxJ0bW/3tDBdUoPbDATPm/GVAldqVcnnebbNPEUVfTlKCAM0Wv3Uq
OrtRYuGQHffuMHCxe8QoyvYFOnbVvHp/6fFAkanSgm+oOPObRIo6qFvXWfgHjCXHl5/36ozxKB+Y
UKZ7O9XMSwDu17NYG9FFNrWZCaBrOQrlvD0TkkusKcg1rnBGL9pCDdfFe90Abvx8tB2l/NnwW13i
SS/zMRf1wdEMwL63saMWP+2xLLH69qFSXYq65//AxzpOKGNhN5GyS7l0ffS93OcdHqJU6JLxzjfE
4cYGV+NZSfLH6zP+k6MFjKYL+X/+ZOGlYCfPEespEHyMRwdmpqSZoAIUcsv6VDUNZDeLlTW60tbu
su9dz/jiiBQwwUuMFmCJ8UGebwTZNhDlA6MOu8KE4XTm2SIwXnBiTEiOb5hOeG0v/Iwf8zKf8njW
xLYLgGsgF2bDs5n0jhfsS6hhk95VGPN6iK74T2acIdIHYFAG2bIzWha81owLfCYdlkcUwhEtz0Eo
fDkzFEp1Vv5VWCpSbB+sR6xhZv8F4HhOgI6Pp2m1srBdxMiXoGQbA5j4zLi+9DU6qptoIPBZqT8D
AByfkNgfX/DACHHz8sAr3gQXyeMW2u44fk2s+Zch0EEz0FNZg3/1KkYOaeGPIBvUbRJdOJ2J2hwJ
wkLGnjJLzv9jTeeo6gj5DktyPlBAKZoS+FL4EzKbEvYOIi943T1nAd2lftV4xgvkJFjHgpxBCvqC
vDAKRwMewYZDFVOWMUPaWMsKgx2mi+t9y1856Ibg5FQ+eLw5Jmy7bo5B/I1Rc4r+tf5LMBRJ6ABQ
BJRRoddBE1+yv5LG/WEeqSLrtQl8f6qgK38HPYxO2wqzXYsPE1rT26xkeloOdyqMUMfcYYuCNJTI
qWWLHlS3MTf05bdYUarEPI1IvDXke2P2GPZhKeDI7FpTUQybTveAZGHmqlaYxkgWh5fQMOVds6ru
eR4oTdsd7uzBhPDg2meOV7BD473qJdirsQvRogROmS6jsgPlMjZR2XgsAaU3YRN+2jWeCIzmr4ZQ
HiMhRtEtYayKo6xA0O2Y2g26QZWfNui/YyJMXke4erHBlxYGT3O/wWEGgpMW7QhfpVn7Nd1SIVZ/
yuOglZv4P5gqyT/5rYfg6KyYkzR39Q5tCK1Zxi/YX0Ff5isx98CzRtoSaUsyq5BtkS7bb1BPN/C8
HyOmAOFig5EoJL6eemr1vGGMDKRcl7eAcw4Cl/PnZyOvdn6cNzftXjKzCjPpvTdbd1g1osv7nrLG
XICuAt0B7g9lPExZjnpvln1jD/kNaKW8+98AW8ofxzATVZgAmSy7I2ZsCidfdJ/3zkgcENEZ5OBN
rPIOe71LVZbxqIbJrRK122b7c3A/olKp7hGTfdIkZmURZcJz2HPIxWAEwWdDzQ9dA/TUks7rCU5m
Hii4WqHEQ7ef5PvhjFqy78r1caagfjsywVG1axsD7fPf/O/teGcetYCr67FW9nyQr6jiEP3ha/Cb
gwxKfsWZSNPCi6LKQs+DWONCRUd7BzYHXevIjSuUXVZebnijiop7nxQAl9WVg1+NgdLRVCCqFyEX
XcK+OkoSCtzveWimZZczoVWSCujQ4ym+ayHCLzFvdlP8OmNXZWe750OCrPZ+KlWx7k0iheSximUa
BJMYDRUgCpY50r42y0Z/+EI5RBN/bFJcRr4/Am+m45WXheYXeAO5FJWhCbMeuGedNJvjL2MgNQF0
CeADSgo1JV2mAfEWQ/dWCTsXxR3VQJInPh8rm/O80+nwFanGDr4JBdBGkODROTxi6cFVYrAIOYFR
Lia57xgCUFvVNOkZFvDuvZ6Z5I1nxzz0D5KpO4OeXFfEpKfdZDFKRI2jAhlPkxTiUWHCV73Tjgrd
sUE+65+pN530734/5K9oQBbg4dgWV6eyYpaB5Y1kBm68fspXjhqr/SLo4tdzxj8fmIy0daLvtzBx
cKW6E/jdxX0F3oNIcWyCv1GhZq7Jkhzc70/FdnvZ8nsBNtHznG/Rvse1KmcsaFxLiNvZJM7FW5C+
VnEXhIM9jMeSGrVOUYauaJcRK1KiOTPscq3m0QxVQP8dl0IgMpW1f/Zea7vdZpguxTy/cJfiZl1W
27OiCyqCe2ZhiOE2SjXoRQKn5Ubs1WUzq7ZXiTItYGnJufUDg6eouer3hMRvTJn9jMEaNKn7vw3D
XnVwY9BB+ou9H/Mq5fxNsGeAdP6r3scJT291uVlpT6l+LDvIjo9jVsaBMwmVaU+kCTRxJmalOURG
Udwj3l/fFGrKkAb1ocTo13uj53tX7WvkaH/hDhXjnZqYNM6xmhgebLQvg6TMenT0imgRNCP0TQsA
2RWBF5vdsudTSPQP1jFJgp/oKAVVZYu+PegmX7lNrOI/aMw0y0nD1bGQBkRyAg5Y8pDREvhvh14s
rHYzbckvxQgwU8mQCIwMCoFCGm0FZfPtvyf/6Xe8ysOCUkC52LRnvbVwwW2HvqPyMmUAeqc39CL7
Xs8jLQMPPb3WnjX4v/dZF2pjO/VN6SMGiW/U+8z9Fio59igO9jNTP9UFmghelB1E4IExcdiMiAdb
e+oA1G8hXGFP84Ntox/aL3SLIECtG0AQLKteVhF+wDrQgwed1v+yPjZwEoNWTMoJQtEbY7RxnGln
wQUP6V96Nm9P01Pl0X9bp6pzBuEYElyo6VLhpHsA3BzYb61Vqte6VIG8rWfmdZ5AWakLcxXjiW6J
opQg7JIUq88tSckZIq8dKu6GoB7wqEXHl3v6f+CJKaIJGQ8z5T+VU/K0pUJs6subY27LeHHyAo/X
wED1Lfmkgle8ZF3v7LQkz/ZgZn4hhpvUGq2AUoer4Tzd/Y95T9LObXotTFKhVJZVh3sQsNhLE2nL
KOl37eg2n6sZnOpFt4ldChGdYp+sJIlilHGccasxL6NOXJcSf8aec6K+Zhc3GoRmQYrQwOq8RbJ2
q68un30zrFGnE6nLU2jmyiiXrlC2qFARcNjUp7Pfag2vN80zQrRt6PnBfcctNFU+UlGZNWL7umb0
mgKWGMIltkOtyQcjxhbXngfIRraSGAkYXdLnEPrWLyD68ujcpUICbjhiQDn1XOJ3VPOUTMMJb1rM
6SZfFkPj9KCgUPGaXo1NcdVjw+2Es2Ajk0KZYODplzn0rbxrNhoRnOa+R8Tk78K9JbqEzgyGSttD
Afn9Ng2OkA8jMvkz5FzV7AoWfFbiwOGYN6/8TG4xa4corv123fwsHqZGaXh8UJPDQ3T9MXGKsSkD
ck3tRCe2TAD/4ImgPAZMiVJnsBmMkaN/05chFevSBmPJSE6h6K57LcwLjMkOEKjlnfriaakBfkZh
rahTtrJm6Ni8iutIObGz+SLUTlZqxh2AtysGojU51N1CNkC0uEU9j6ErPH9TVsonXKAbD0wgXWJM
KBEGDOsRN0tICuzwIX98mfsn+rpy3mBGhS+XvXCsc5xYzKDvl2hHIE67YKaHMn0HRK5uV4Z9dzOt
HGovmwJA4dxiAa5O+2ILaeOJPG1SbzCAlmAhqm6NEI3ilIxEcLRJDch99clEZBEJ1JHk8C5WU7K8
ozQ3N4e5+rxPFfa2SjreTVtVbYusVHuGz8CA6TkLYxSxEwQvxzupbRNBK5WBKLeoL9EWSsAQ9k64
ELa7Mb6q6L6dXHeiJktUaveVfpUdZpcMqove34gBhUrTOwppQCJa7o5qDHF7oCLmgoFQzbR/wTVL
chkyf5OtrcJW7PUIajC5ZnuvSkyoe9p8vbLa32S0u5FrL/LdHOdYjyBMzdPKMQJB0kO+AnpyQPGJ
ZLHGmCP5OZXxlm8qwueofEsYa9Z0h1mH3AjDsBGDRH9nAG4933iQTAES8YPkTmb3GifwCX0yiLH6
2X5pX8ic4y4TnF0JQ9wsDuoh/DUmYOz6agWIEkIo7y4ccTEUzC3WMvR9AzivtEfmIem4XG5ktBbf
dscMKEXDg7IffHlJAY2QoySURX5BRpG8MsNty/asDoNWeraEJ4P/vykUIHYQqmyKmSNutRRi7Rwj
P1nU5DOzwrF8vgZS2fjYm8RfG3Ih2Z4fOHhnnBTj2G/XmwGtejNWGXccPT7x1adtquhnkEdNLcg8
s3Xhs2H//DVcECJJo7rsu8Oc1cWVIS1+jwy3YV+DU4GWIAgOGkfpn95E/qs9kVk0edGHr1rI+1df
amc70YrTHqo5oUASyPoMEhuWcc9wveGEZSMF/6pJlkiUE+1/3vXD2EOY55me+TYv+cpgAn9Jyw9s
Jc9w7/AC6xDoGuoS/aeZx/Sv57lPNR4t2Ng1+sv9a1iYKRmzL150K5htuBzFgeT2KsFkgIaGxtZI
4uvuCtK+G1Z5D7medtRt6q5JI9SmeHE4uze0z0WDcl7iZB1sxuPcCcKnetixLfmSNsE0FAdBiIhA
FggVfJvmuG1QbaZv4OK+9rRtD/Uko1dKO8aY+xVJOUuA+ACBcMw+wIs/yeDrZaQTeHIs0NTTlcKz
4Zdiekh2S6chceWbgPPDnHhCEa08+7KTCjL9IJNE59SK0kyg9cg+kBfLFCYTXUBoL3zlZIF+i00y
fl3cig+bg+45PZ2MK+9uHJYhYuQ1Xajr5FSuFu9QvrWO5bKEryq368ACmAKo/2XxWSH3PAt7sB5R
VsmEpmz+19Zuo49iTcIgVbWMUChCscF+YupC5e67L9l8XKbaN5VIR/28zuIw1rxRvb81tfCe3RBw
cGU10upc7xyj/+OieiRKjY54/aDMKDV/x5u4PPc4OkndImoXbaemDzz7cFG4UYB5cGaRxPIPFiia
tUONS527RQI+jq+FJ9skiPI2nJIaEwj9pYyot4Yxtuhvuu3S9A0L6eM7ZEv+15FLqNihBdM99fFm
m6M3aif8E1An+Vgut5ob/AQ2nyC5IgaqqEDfpSlp60aCEqdn8ipWXTzEVgipsWbASPtv7nd5SeyM
DEPw9990Beg/Bczc2vzXs6LGYIu/LMMc8OR/HpoCeAtW9KKXOXmpFE1geTQfSSvqynq89KH8zarS
zVUUtj6A3f1KxLwAbN3gI7kk1EOLhAP1XJ7yTco6zq8D0nfSNGVzPVAasZnyXBpoPVZiUAVrpB3E
pmgG2QtAR9bYKfpfE3XVkwCzoahaDV6YYUCmSlzWXKcMqDcAKyUvPxFu5dKrWZzhzapc9Tv28/5J
4g564Airr/rpmeSBk17C83irKqCikUtooc8Jw/jBNa9SSIierYYobs3B355ZqKJiT3fmOgQMmeXV
6p0JTFQJXyFoXt1YDy2zU1MVSXR0nDzNgsUuVbNHM1v5oFPGhnTF+OEQmAAFXx7/IbNHEBBkvMv0
595CtRNe5KsGRjtTsXx5XeNZJKhV1liS/y9XAY7y0/EdJBeYuJgO+uKZOeT/nLXKoGfVxVeWUia4
raBmrXQy4uiaVQaggcuv3CmkhL2LLVyaEMlhMWQLEvf9a+vURA4A0NKqSGG6cTUXgt1Bxh2/Qccv
LbFXUVCVIU+chzztcv1VHwVUH4ibymjpvUfZzqbEbcwnmj5UV9095hPWPbjdJZ/lPFByDSP5UbBD
kV4QBoVjEaCaALs6ONMYilFFXdBJj5jUh9Kyn8uSZu2L5hPdUpV6QsfpzIgzyW4No0Nedqht6f7B
uW9wR2u0BLVHLS+wWBdf8Q09gIZU7lv0N/WqcumK3q7jqmrpfh91g/ige2I+kp7XqGLCmpEXhq4+
45kZYOJ4yEtiRMGvkw1hzAN6O/ib3c9mXmIyzLauup0pDs1mOq/nLrQbftq1jaYtBsDKoM164L0m
M5Uw/AzDaPmS/LNivIrpAGBmVP7pMYHY4Z07L8Mh3fdhd7BPeCPji332vU0w8nsyEmssIT8gnVoN
M/PPOkaFt9tUNazxUNShJNfESjPohupYEiejgRS+ZfMcZpjdsC9SyalN4NtnB6n8lB4OuqyADQ5Y
w4fgszM6nxgmobriDM/Uacg5y4DdZC1vHi2QWeU10ExBLM6teXI3Nr+CAi4Cch5Bc/hC7CX9Mng7
lewEQ6QtPJTJuYqxh67fQD05Yo0ITBkXsWcoHuYNqNYDO1p2mWbosbaHGNcLvWXSQ+n89gtAitgb
e9UcSVnpdcsklw8jl36CilazpzrI8IBLILmoYelCtQMe+ATE/KjfSRChpl2F768BOY93WTmn20S5
eQv6mgvJ16qFUKZ04mPWGw29Hv9LBCYeB/4DDgcEUGUBG1Py0mJ/HWJRssVUJZFMsq4uPuUvd/Em
el3iV4GgtJzDQGjF+d1m5zCN4stiRtFTpHz9Gc8k8t3KrQ+JoQ+HH7cCFPDeeN+GBuGo6JSDK/aU
WG+EYz/6Jk8oZS0O9M8gbpFgI/DLZVe1f8mypk9c9045xByBvPFYk+aGShoGPLxbhybWWnvmohX6
uHwtfA8EFp+VT5CIqjUhPaUvTyQKWy2ZbVk28C4e2PYRfpebIdA/lKH3cC6+nJkOPIKrPiIPSXKY
4XjhJk6btuE7rdT9SbtlY6eSV4AIaQS577oFb6J4BlODImMmXxYP8LecYQLQgah0e42QH1QKgGY+
bKAAUt3x1Tkyq64rBIjp426N3gOS/tFkidz5GxW0GsckbvGcSvmnWUcNy+AnNa5TsvOM5Enetolc
Jdt78aEUywv6NBtFPRFP5c+kVg1FZndV7cN0cbK0GXJwzJV+lcG903xDOWqR+agvYzSv4HOPriUz
P8Wi2pqGx6ped/wsDAYRIOvdEhGtNkOqFfPDB2iaDx+ZrJtWuO1CITvgkWz89CXwkqxZUurF3XRM
obu+ky4nUfSdIPHwTHiRFXlXLpQrUjCVpQshvrzPtbNgbFkLS1Vz8YXkyPBlOUwy28QALIDDInSA
3Bv8iQzMHjyve1z2j1ZSR+fKohkinhsC6B6ouki0A6gjjP+JPA5TrNMpZ8R0h5i+/AQtVlp1Pz9r
cNekVdK6NHpE2tG8ZUMgb5LaOS/8gh2FWsLWvaxxxQOCzoYQc0DvZJrUOi5vz+dHzUjUpMeYmtNY
o9pDFfaKuJy01IDzJEEmuQNGyMvyPByzHcsOXQ4f6E1VNZGmTmdOLnnzb52OObaOVrItLpFiHcoH
D/uvw5GHWKVCIepoL3Cic2SCvYG4L/2APiD3hHSH1+pmw5uHEmM3CXJbEZkuqW86nWwCe/ry7lvf
L6Me3nrGdEvEgeMzIUDrGvribewCloytc+VfugGajeYWpmyFp6bo6CfIpbUs5OsXEJM7wmVY33Xq
zW5ejuYzUZDWSYuICX6NxkJedwEVXpFM0eyap8Bw/fmmpvC47BYjzpvKCLJzUthwGQedmGyRRUdG
HBjdLtEsVkBmEVHhcN/5qaASN3zMtsJg6J+92wgI8a8KipimMk94yAr+x9gwB8ZwwdStcejZBOCy
4sEhZX2ZSZy7lyEIHodgdPJVqT1afi5K2cxXQnodNxCUEDn+SR8FEEfBdaXwRcc+5Pi/QF6CCIZv
T/qEk1wP3eVS/sZG/yVAsugMapYwj/XT5KaNJJLs1ND1GpQX/504jCRtR7hPEYVlV2fItdxql5ZV
FjrJnRCz3RKmfMQ3PtE7DuK/DREQ3Je4Hvv82AEbNqakWivhLq9GT7b+rV77w56gJvHOUrQVb4rX
WapvZLHJDtgOmBDTIuqXVV7yNSUAITCsWkw+bQ6UAH3rBjKmTVm5kyF2d5ihXzXj/DJKUDHyyGiM
kpdzR0cm9o10HLW6WmndamZMpxS1vXVr3Lxpbi+0ysrLt4eyxWRGcb10IyETnEjxZLmEclzvZfzM
pNZ7aCz+WXJxXt0J3VxN9rWA8uq5qFNvUoSOT97QzzVrakheaEz+3PRmbLoXiA3XjSuJwQTKYcxI
Dk6J2F3+LOMjJYNuxi1gbva2ubjsyZnzVmaQ2Cs6vBJZ70QQ7+Msc4Q82C5oXL18jHdzihIinvHU
ba5tjTYH1irL4jqSmFrWFwuK5HgUeMarA/vd0jhlu6Pglh1x7YQFpmrOuj+SN+C2B0jdm3xIVlxe
hWAH3JL/yDE9u+VQy3FSpCT6OYxiViodtg4XgB7s9iaMmFbjiPS/ErVzqwn52aZtuVuMDZpkTmOz
ndInyL2asHOQtQawpGecRfTUtxNExbnBV5p90lwIFMrZ1PeM9KKz9wbs+mHGO98evRoOaUyyDSRy
GxlRH7veMlpDlUmrL8Uz8tGaPvYyxtR/LoNE9WHFjnov5itbZ/PNhfOhfqKyvp3ytl+qDO7sKJeg
OQd+AgvFC08EPoVsiBPSe2mrvA1ZIbK0sb6QyTTaYR9iNX86smH1hHsZE4iXP3E7de164sj/J9YL
DJxqRPnjsVfp4hVHsO4EUPyRXCDeONIUK4apaCBfMop1vZ/ZSipNfx6YG/Tq3T/uYoWDEwMqcoV7
h/iKJkXY/prfUj1YBzlzWauDVa5nq8eiFIXlZIs07JtbQoq++ec70p21lsX9sIMqC9OmHP+qrfTj
r5aXbZRsjLk5nWqYwofYIr4XvWTuuSNktYC4XA74Ei5U/KAhhpSvVlsc+2txS7NoGC6l9AsdwIIV
FGzClN0EOZCs2+8wM1SRrOdNFg7uxzO3QE6eNLNK16cJrsARjGMQe9l1kI7wAZkZH5prX+32lrRa
Lr2Fsy8ZBT4r9tJgMqmioZCm3P4uURS8Q59ZzcYZyzrmUM/5JQzoTX26Ni+h6W7YhZRvbKpvwUQ1
ytTLNmU6RD964Hdb3xY6BDBAqJIlH+y5UYSLOzGVRaZs8YL1CiIOzSy8XQDdeykralsym+yENOzi
HVdPb71LjJAmioL/lu6DwG1C9YrMg41WG5Ub504tCr6anNe/n8dNjvqRoX+NDIm+Acaxhy5DvDVu
Hw+saZrKLtvbfxakzSppKUO7mEvxdHOU4GKb4nwBM2ubci8m7eTz0180yhEzMlfXLgeJ/1rK5Lla
lv9YVlxNiM+mzPQXPBA2UafEn50TM1dxIx81fhuUZNtlsmIvK+FahJm6Y4kD0W8FShl8oxgBao+0
+iS+/R4R7UP3Wb345wC5vTGekgyCCzeRmmnshJ7PbEHtM/s4FIPAmwCea/39IU0LEP77O8Nmrvu0
Slg37f4hBn5LNi63BT2v/sYRuhQ/OOI+pculkRLj+rMNqg6eXtl9RFOg3KFEHi72ip7tMtYi/NRW
2qylVTX/4YEcn3EO6SS4UOoiBWmc2ZkuBeTBIA09EDrb42xvR3WmoawW5uM9VytV26lC4QJE+6X8
MXw8T531skhyCT/YN3JsbAX3AEvflMYJ5IfJiB4ZP4Fe+yyD431U50sPl/TwPqFZdfp8bWLTfHdg
kQ/rQpgsLTW9dZaE36X06yrd+K+ExNjuNC+MVbwY3tMhyD8unwdXr/YEAXbcrBX9xbE6emp+QdnJ
8YYo4RUHTfbBopxP2QG49/XV/NLntf5PUvrCBt1FOI4E2sRZg6tGoLQ248KgqxYFqIo2aUhmoPXe
AYHCjdiH8784npbt/zKhobDpjtGOMel3z182704WCiMDmUipaegb9tvX3zpT7bHvSQlypq3mHdY0
Ms2h2YvsurgHk4RDDtR+h9tXYGLWVPTDXOhsfWdlPmPsQVYMyIssyg+ZgNpMECmYJQLRSVWylmE8
Wz7LVV+/l2QL9oSWQBa5g1QpuFsmCMGNW9G2AU3MIRRtB9mJQ+TtzmZphCObPqpLzhbzbXo58Rzh
wZLvyQbl8HdtUl3yh/eJJd2dYz8dq97tv/cgNsiDt++eM5nzh+cxXIAogVOYcoxEfcbbfJqbrEiA
IstCELS62flWh/hOvSead8G9ifwfGa2dcLIkhV8GHsZLRmnif3yBrGGnfPa0f5KOgkP8JI5ZN8eU
OuAGs0Jz3kTSUTeliyhZRLJhscrkbXW+FBLTABbbKAPwr2V4q8XnAZZGCrkpr62MbVYQ3bwpJ9aL
PDUsvDKpIvFUIpHDYQVEcDvXdVnSmIwAuoxG305TtjYgwTnkfOJw4HI8uspa02xKXEDKwpLWjIG0
CIXEIChQiI4as6SScEL1KkDHqVMRSS4wCeoXdQCNy3xe54uf36SKujXViX4zkfMGmC9pgR6P8AlU
D0pvM2xSvQpKUVee0pkbCtfdXGvUtKJnxnNIjaa6ctB6akaswcvejh13Sh/C3VuQPZH1bcu88FUH
G2yb9+TTqaAC6tdU6z/Z9GJy6QEaYtWj2frqQl1wdVWN6+Jdgqbc3Wod0t8tBwuVFzRlQPMSkGvb
ZaPR1yYOEWOYPHjyZviHrIjfsdiJk85XIyLSmZ5yBpf3fCKPhdyaxg+Uz5pH0UKQ+8e0SXkMkKLb
XmLDar3p55a8OznvHopcJCsUn71ydBPTBi7qB+vIkO/vWGX/oVCwnUAGSTPc6v9IzlUcY3TM8LbY
5ExEk7KU+I68lybAhDnzETxMuLXHLF8nMam7CLKbJ3lKqozKjOdldaX7S9fj7IJETFYoRNoGNiaM
sQr/RHybSpQc9aKRKWlBv67oyk/QKXpocT47+NtIvU68toGo/Ew8QihxirXLclfOYcH2FJj+eaqG
l5ALv7pWMgn0CwmpdUuIRJzUoDkzBbv9/GCCiXl6mXC1scjWaGc+u0OqJ3uYUprWEjoyLYXoc4GC
0rGx6BjsrmJzRrBq9+uzYEvQAiBnIrR0EtOlLlIjK52cDd0fVV240a0Hvi2dBDfXWO8n482Q6fiI
n6q6/OmhlEeCJrQ1syJQt4Fj9F8s60lGRBwp6EZy5x4L+qSzt+WTXvwPllpCNSUL43vs4I3C23ND
UtGNK8GNDF1ZOknFbbjf11RT/Qz3YVeA2T3PuFdomJz+qb5fHSspF77t/9r7FbmD+7a6UNtOxt1X
7KQn75g4cuOnfpX2ttKjPt//BI4PWBNftNrQDYEaRe7013FIQMDA3MIPeagoun0LVkIuhF+Te0wz
QSe1MF4kdpsD5SOVZWfGngcRbPjWJgxRcLU=
`protect end_protected

