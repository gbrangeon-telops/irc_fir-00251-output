

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SPpb0sHtYr+7D0Z/NdHkBGKHFj6bPnAk4zCT9Qd9jSi/NZdzqHWXjKwgFh3NrYG/AQMVJcT4R9KU
T1kWm6bsuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PM0w38wqoKZTqxD5ZMv+He7u+x4mAKOhS9vNWqYsLtlMu2ni98hkp4Js0D7iFCQdcFCu3Jaj2Vqe
E0m1H+UGB6We+zPa+TnTKUC9+mxtEW7xpi8i+GVKfIfe89n3euEibIBIS0WLtZypuPRjuzr2TWw/
TpBFYS1oUTQ1qwWguI8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OIEbVz6QJBHT228fhImFLc7Q94gbSg/QOSgeKpAp1zRCxot1azeNL0EHN3pwZU9Qs6kuTNEAn7+w
agqdilWN9rl3uQlRBfW5KbIj2khza90rK/4UYrbcPGQyMxF8l/LBS9RaSzH8pqlJgQ4YfgwGNaq6
EHHkNL7CBEprP8VBO3A9geAIYBWstNirz3P/01jzH8PT87csZHkt/KV+1ancvBdl8zy3Pi5RrOtK
WdR5qLkbXJ6m4DjaubrW8HdK/fqusuCVkVGxmajuQw899iRpx5AiTEwKYKOor3msJGxdK7STL4ZT
S1m+Ec1GdsxDwYBgiKT0A3c1/unIYBS6y17V2A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y9qoE+tEhAFEsAZgxeFxNUflksEoY80RYly6rjz4X/QwncMYkOdY5w8AxmW4IYZfWprQfyfkxMrN
8JuXogLHC84iIPhEFIhJ/+RivFHW4gCUIf9NTOGEkQza7hd31B0/7LZttbZHcfTR5stmYGMhB9xi
VCriwe4C9iR9zFvOJxk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eCcOM7HngIZB2JCDRQ//SPPOptJbtDQ6WJM03A6xR3t8OhM7+MFavTdB4aR11UrppwUsYiZCHTBc
4AdaSSNbTEcILhRaZMNZ85hgqiNgFb3YTJu8ZIWifM+Ad5U1zkzbH1xsVssRl/Sl+cf+TCDh9Psd
UOpjIzWfsyGgyfaSSbczC/DMklBqFcyspqzOP0YGdgI4It3e5xnwDvYeewRqIZggj0RyjkJH8PxJ
o1XlyTZFQZIIFN0x8sDbcPdsUekU3pOCvI9JK89jigNzKmLJRotLEgZQt0B8gMiz/gm5u0+k01OA
f/7Xo9TSexSaZ5evmswsNTBQhg4v8j39bgkh9Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7744)
`protect data_block
a3VgoGxV3FEw8g5rUimxj6V/GbMnaTFVleX8/8AY+3JjL1ErwFMX+XnADULua8RjGcMuAgoo1L2m
aUQgAz5BYX14vxYozA2+MiX00oCW+TMKVl1YphmpwJe7UOYTL7bvZ58lGw5vwVQFMry4iu23PMRw
PRSQplxY1PtvFKVbIODLzMpfZergjeaul1rWNdJf0eKNqRi0RSAz42rfC7FrVEENtER74FO4Sdnr
0n+QPXtBoJ4sFeeD8w0KK2ov3i8VLzehHjoxzVLuA/fiCRiiE1TmZeNkmmdhf07C7rjNgyAxix35
kW2LqKlkkCEN50tTC9RkIsEJp+0c7rMtaC9we2y+0rF/Hujc9viEjZyiZfPuIYUJrtzqxdNBWypU
O80K46G6pPd+kxHyWmlL5/0oNJJ2K0AfhgHTjYNMgLscU7mYMsUA/6LP8nTYA93XLL/Rx7871hli
Kii/Zqb32xxQ11fxFuMchFYHTkdxPR4JTO214NYobFhUrEJFWUWG+InUEDlNvpYrKTL4aqkAxMAz
RnT0h+L6zRpTUQsjXlLLWhkDjOwU5mg1L2/gXRjFlPfXQsm+z2cFcpQ4Jdvo/y60h8haQlC3q5oJ
/q21qMa9pwvAd1rdVRYKGZI8NCJfHu0TpUYiGQDSM85iBk8PyGfDsDZ5dLxhLJblxasAlLjqEG7R
kmRLTlMkqtHBxJq6eyMTMJGWq6wcwyly1+WOkS6d1/O9QVgiIBA9XIBV+/fmDclmQdLo1iDqvivj
PBhBRvEPpgQ/zUodncw7CyXQ3QFUigHpgQY7wAJ0lBlczeZid6AeQWxQECuoSh8/lmxmtVrBoEub
7sn4RJ4dyh1UWtGKBt+So5lG0md69JGuf5F63keRpFGUGADxHsz3mFBo/ksgmbt8eJOLRU4kaDZS
3v/uJd8h6WivR2RGyJB0xnUuVPgyw5qVeiFrye2XZFvU41Iu11TH9JZ3rbw4kkhHS8e6Fi57JO2u
+0CXqJZ60kxgZK+FASTCX3DeP4nvv/AHbdbyZ02bL4Qy1W8eUUXq/ozHL4KLcqgWUM6bGCl437Dj
++gOs3paYt3Trw0zvRPtRYhhDeOKjvfrxOZ9tlOA5bG7bLukx8TxMKxhP/tQggEVBSAqJSBoDUzV
iNkRZTanpBSBya1rKcQPvNqyTcGvRj1Or4lJqwa3Cqjg68YAF6Hb0yqkgMJSrp8ICgXjB9dnET4t
Mx6+9hyXtKQqb9UIgvskvU7jFjng/VG5yQYG7yVyDUORrglPii7dRm7ao4Z897JwSewXRx8iuT9z
7sXCXk8frdZNI9u3a87fUCwMvmITMxxqTtyfjymMOAlSYsKEVplf5679Btro50d3b4oGNd6VDmZu
GG2ZsKdXdMnaxWWP+moqWI/PqUMsTME8pZ6D8aPZzXiBkKUiMIuf2d61v3O1TPkiDaBD+jPeWjoE
NUojyF7VjR1pZjC2MMrDp9sVB979AedZ8KKBahWt2pDGppm8OcQyrfmTQr5aJoDCCfzC51tGzSo/
qOzrEfefCeb0bZan39GL91LxeUoDRE62rZyyt3UWTjb40L1guLIBjPq75Hgu2YDl2FHspxremiJk
mdCFuIuT8s+WeCpK3YPDFyf28cs5e8M1BQbxSWU4StU0zxcgJzEaT9xYp3FVsrobMxBY6jeVamm1
PXLLcAd5qx4KlSaUh3PjR9BizQPIChB/fNz2b13s/XdfZg8TgXzRjVF0k275esG6MDzCH+JofMuD
A3F5rrr4M0QUL3oaEG1a4un1Ghg1oHmCFhperCr1XRqEwqicsuDP/mEfBUU2HRI+cNemWdCYMb3T
YTcro6AsGlrDujSSsvRzDQzp1E6swyqZ19iuZVoaVcE3Ah/SWEXzzGuXSKoDPmOzw6fW1fZihAsT
0otfZ4RZogi34/XNPOPxEWZqt04E98YPqfQiyvWqB7rY/DDMFCVkdLg+5VdaNrHhQ6eWqdM9sel5
Ve6gCKQ7E5UnbeA9iqnsv44hUhOlf1qs9beCEtshHVf16Rjb9VI+js+OvgLtsIJHZqBLeHM5Sx1a
88idhd6c/WVIS/d1UbzBUAWPt427o6ERxF5bLzHGo9Cv/RnQJWfdnXGg38WaXIWsYPe+oJH2ZhKp
PBqI4VhgcAHy7Sc4Hw5bQWHEGodFXeYsphPfbLhx8OX/y7T+RvPzKrd8W7489He0xY8H9U6/BeWk
QGdkmuGx92Illseo8sL1ohpTbygXNav2i+fwATalN68R2QAuHAE5UNPW3bRWmqmRdOQtZYCDwbNx
B6nhuDBqVgZmOv6zEI/MljHWMnIyEbvSLw5sSpqfbOlCny2dXOWJlqF7Pvllv2JlmMowx+mzRvqk
AIE0of14U0cBFmFVKtCFlbzbfdX2JUiBh+RFnN7Qjg/k3RXcgCcTj6wsLoORb98HYUqcfmUukYFt
R3PF4n7XE3Itbka3ntr0eA4Vd8hTybu6e88dcXVHHLTSu23pS/aE8MsTrGeI8KQUl69KkdfX4wcI
YkcCwrSoAK9R08gP3ZlHBzn6Id1sZwiHNPJF2ev1F7Wrld0Rp90DS4oqgUiAKyEIURlVpPcr2arn
Y4pVrNODHFmqD30vCB+kaAtgBAiigx8a7lvvLQX1oMq7iYJUEcCovqolUIBSaGHhKr0zKdNxDMa5
e3yccfOpD//NigLjemgmYD6NDCZfRwX/oZYdOjSCmR9dHvBcFGEjhrJZ/Rj3o2/aE2+wyqQa2sUd
wz+ze0wWyuk/ryunh6FKvkr+0hXnDF+w2e6SnPw5MeY2T/EBzcv0iiBeRnLCEuai12RY0jbCddoQ
AZhjfXr7Ios+OYYmkz5Cewn4nevh/Or8EngN1TGbtKH/Fo/1g7zk7/O7+o/LynWDIIrXsLR1pZfC
lVrbdtGbWY4euDb4RimngqfzFYcnEqP12ilzy9MqOQyQClbthUFPm7/6GjPVSvCuHji5SHmZ0uzb
aY1SZUHvY50W5HwlqFyBQra5wsVp9eO29RH6EvO1E/fJveeY6rThjNtb4rJ75mE1KHA/j29oV/rJ
aeS6fsTMZ4hdWAo4ZbgReShRoTDT6kBgiej7BVBQlSLg9sY3thBnq/mpXOcn39ASzBA7Y91pbyXr
Px/CgYomCoMCWm2EsunjpGdhlG2NRvZ/Q+96zGxJiTbLrDpMkFfll7kTTSpnPqu0es/5h45jP0RW
W+kWfWwj++mjjOlv5GZ9CPHSgfiPgyjm5BvHXleRmpStadHkwbuNpKN6MvBCML/Vi8m80Or+I9Nj
QDAa+/ACNXiKJvWvpo/6zDA73/TA6Fgm1orFFSWJo93qhZpIbYx0b2U/lFrCpQ8hmUvdNP4o3Czo
qwNX8Ndz7zFBRyMyOiuOuZfZUL3A++EP1OgUH3MWD18lKcy67VXrOOFwKaEiO0IUBoR7M3epkv8n
tOYzNvxcSyspp5zkioleAnq0mSeC0l7x4Rmi7P5fLNMIvH8LxNeBuQHPdAvdegVtZPKZYRbtes/e
c5YvHn4gdmeCAckQQ48JSVwPL1SpKfp91E+cmdAewAXATvvuEPwxzxGPk6rtNh/d5rYC0AliBnNX
Q0NzbjFM55AcRrQjVX48woVUwPamzbAUwMB6fKs0BocLjEKv+1uEcytxcgbMab6Av1d0yNrKMwu2
UC3f2iZz7fvCCJJvLoYPTCs+Ys+bZ0+FCtOqmsLC1LM10JrKgAagQ0Ds2WtCD7jcd174VdrEIQrT
IefPE5b9NyOh7IMCNXS46lYPUHUFopwQIuyllbcDADO6ujNN+bsBlMbwMFzPr2lfRkUg50ukoqSe
2mzxNoBn/el5ZiPLCfWGgwnu6rss2pMdmezr7lOmAwYbkrUrRrKJf+mHjp6EG3ztgzJiIl/Whxzl
NfP3xxW6Z1PNWZPxfulDMTIw3eSQFC/46JtizReyG3fgId2dBlANe2M5V9q9CCXMat4dY+jhvOqb
jm9cWzDfVJ+bynroKQz7X3X4ztZuScwHFVJD/UKbU3Zj5Ujns9j+b4qD0nC7Bp6suLsb727yShAB
HwH8yV9J9TxnFuBEvA3W6y8a0OznwPTPLr/ypFW3Vy91BbduvSd7O0wlyV5mOA8+3aeqgqozMzjf
6UIutOM415qyUPiZLl6EhPcZfxQWOF7a+vWMx7e/MNFebIx9P5/2XL5MH2fSTTztH9+B/cIT5e7V
2AZqAoXDZ4RMrKZZ5cAjO/X8BEOsBr0ORay0Yx2nQSgF8WRar/QjFN8I4hHviBXFv0i6u5K/hH/b
48CfVC9FeV0qG9ZmlBc//b4QaUHbPY2fr7KJR2FCpX7jcUn5nd3d7wlgq+clZ6YC0kzzW8EoLPjg
HUiJ/JqtfutdAtTjdvvmo65YEijPxQBt8QDPmOHZQiBYs1g8xQsgCcIgV5/DWnUZqgC8TlSfChK9
b7prLNGeWHMb5AVDeL9dk0PghjO9sM5dQqP52Fw2i9BUEkvxLzzpE1pyl7jNLeleA1Y8IJqykT5U
PRG9qaGWti+AsvWAWV3ozCn5GljsXTImdlvJsmOYzFBC4/IJdV24oL8R0zHRUBtooLjKFz4b8kpl
Psx8Glmx1UGIUzXyhg9Nsc90bKkGJp2LrJxITgW0+c+puqer7K2nuYnJeMPpc4RjBTfwbnjW2y97
YuhxkuISkp4/LqE9GN3vFgHjI1w1ASUhQHmfEkEJojDGIGi/8yRxLnHamxxXJA8+XvvxAXllET6d
/amZny26l1g/BVMqq2laihL1MJroWiu55QxXTiB4ee9PM0of7lon8IDTew5pGVdi+/W9m7XJT19m
TjgkePBQ4SIxfMb+5rwkmAzM4plqCSBA5BtJk0wfQjmXFIxViD17UT3Zn3Y/IifwEhctz0dKDhDh
0pvRpu92WCaWQ3o+EWW3INhUtFI6nADNsaOqLsMghf+JTbpenJYW1C/gLUO4PBmdmbbW74PquGrq
/XGb4NUNSxgMN0YYuOrtgeDz6Gc21uLrDZFiZzCOvrazYsWB8BcymfErduB3gnpZaQLwRnygYS/9
8svE/TSer0RG7kc1uv2F6kTdxnG+dhVfmYLbLKBB3nSv4/KD5wFzH+3HHeGw7FEI5EwY/qkU0td+
Y1McxLjtc9NU9mtR9TUO5AnaoKZYgjurUGmTfovJvFZbVAu5PXKsrIwgJm917TjUEV00NT6A8TVc
fXDOhcgEuaEJWlDLGE9AsqKCodfD8tUb5cpyuxk+gQryk3GIISVc+L7V2SJkMXPRlIRyING47FEW
/n8Pel/I+w7i+gRIYQJCujHIDgU/vBS7DK7zp3ghq1pB1/MHGCMqTDKDy8uVUZ+H6BoFV9QHW5wN
w0JNB7Fkp43xcC67TNabYLWgQEo7OQyZsj0cQ20oLMCmIvs6Tz0Zui855To9hhg1NGmGy+3g+tzk
PGeoQQ4+1SVfPzMx3eb8ef7WTFpis2IYc37QNiFL+C+QUXALIL3Xn9un2/V+NZZIYvxrVyrsckmX
3/gIh8CJiu1wXgK4V9kGa4EiAnXG57hxQCV9G9TbupAGVOxnwLFE9stSMYi8Bgv7cf9i6W9kNjre
PBxU0YkZOgX1UkQus/EN9jrWNtRL6/O7ChrxXg0ds5I+jYO9UyatnESx3uuI25O0sB1nRddqmN+L
GyALLtiPZH0BKkc8lNCCKKCRdhhUtU0SyAwVJAH2N1KvHnk3HnDtxIUYqBkkWHgWcGDL2rwEnv3W
7a9+ebKzS4bfFElD7Rwhd+00avwyGcpOmn1jGY/g3hD/chjn5ucNrIgQ6ZdtYZqGS1JrsDokEfMS
/hgkyijXC/nadzXJD7ebsOopKTUsXOBs20DeUvZFsbLCKI7LndS2VLKF4uwJGSnwhoITU8wPZ/1W
uLpkBral0YWnBmv3y+dDSO4kV2sqNAcai5rPmQkXYUjHKF5SjJgeYoG3e/QQXM2vmtILXIXjuBwO
nKT+hwo5HeGekFpJ/7ZM7aLbJcb4C6R877Jo0ynmrnS2cTDg6JgbQ99Zub9P/K4krCPZJe9FM42J
sMeFwyPoKcy67Ma7PdiSC9BYw/xNBTs+Q7ycdj6Z1H5o2fW8dVQcUxLzcewShpISIDmlIVI/JeCU
cxTbb4keo8r6FtWn60Sem4mY9b1+VdEEyS/N5Qp+z8kttL8CQyaDlDlEqy48ZXAFKEzAOiGJ5stn
QDewBG0rZmdagV+i7/UZHcZh1s1O68XF0RfFfzOM5iQfcg5Kls5rU0Sn4OpeRJsBV2sG6l8fWSZK
4MzZMwLtj/w8Qt/tX1jTYIGkcU4VddSqNzd/ZB0ddh5oIWVX0iqlyMjTEsHSLo89RbNnZEjHWa2d
9ULouIWHGSf3cRBlK/njTkq4yzijALnXN66dd3OgPvLcgQY/CxvTnz0TGJ/eh+y/AT97ETOzMtZR
J/lhVzfAdYHd811bGAEWgrx2eIJ3a+riemCfZVl4kcy9xx2cxINhswFf/fNax8uJduAxC9CT/nZ4
5RDytUQTLk8vZTXTmvH/j5xU5cLQiyyQK+HP8PotM62e6QKLQwEqc02SqInRzuMm+g51qz/hwiGy
ss3ig8fM75ECBdeyfucHpMP+3NaRvtxaHXMNKn3ScPwOSoZJ0RoQgMuGpBxD3cMkifClG+r0OdbZ
fAkPq2hgHh0f2EARq9bCxJX9TLKN3gppIkNT4A/N8eRwNA8uxujiVaCqbBBuBlR295XCvVF4wy2E
VFKoSBJ/IRQ6lRxDbGNHRxwxgn1VXHkwp5oadc8IXDhwe/ufv3n1VerMHho/nb+GvrvNb9pRsZx5
yN/Cg/EDhoStfpGMfA9WNAyeI/PDEopCMLwOXYlv5W6bKRT2z0FWrBY2ny7XBf7whdM1v0g4rNGr
5aa67ytctk7/1qu+mZsYjRRXHnhmkZ1C4CdJYxCvEX/WLJXs6LVWmBWIfE64Wdc4sibfjjhvOabv
6ZyXq4NB5iPCmJ+LiMYvS4YIj2Hn/EJKmgjsRKWUs/yJSaTHmX8sO8mZhNWbvc4KLZINCamToXVf
l5gXySO71ErInPoXL2NGW1NGlfU69GoWj083/YYgE+43XGpbpmA9m3u8s52sl9E/EpASHAgKzK3v
w8OOoLEMt/x0JTtNBl8Z4u384ti/DxbHyweqMRV58ZZLDCZEcPj/eLe1n3zlSq9kMaljRyt0SM+A
L4wfzT3HS9L3XQsUWykmCdHKphG0OcChkQrGXtPq/RT7npBZ6mW9Li3fZl5kw+f+f6ZrGb39U0Xm
j3I6D5Bx1gegNxEAP/dnxgkf2eih+zr1/MPUnBGTt0UDxkA5PuWRU/8fSssNGh8APr+u52ru2gNt
vueIS2lSWEejdrSw+rRopj7a/VEPbaUNDwcH6MJPAsucY18AHKvEkxf/jPiJf4k2bGn5e88bpksf
eyvXuRWDFRtOnWN1yZ9qpXApb958vwSQ87wIoJB660fGRk5pQKLUSE6sk7bUWYpqrR8/6XAibrVI
IlPEdbUdtRhxt0mxbsjuX24PU5B/DrAM048xAE0sdxyR5EcSCJD4V8GoNCup4EgpSc6iMPJ3ijnp
P1EfHxXfiohKb+Rvs39DiRLMfq6y3XImJxX+43lK4OKM9sW1Wv+3h9ubjPYsx6jQ1g6SR6hYYoir
onJ5i9q6RC6Zpx3RbAOlSYwzhij5Af9cqMzKnKiyPJDgWuLNg1Z8XrVfU/1OojFyOOTuVAtwx3Ye
I1SdcKvAkLdIJb6QivcJdu/cZKFu6gwVaUes42S2AVe2NLSR4ps0Ngy1egO4TFGWd2J5hhGGVhHR
oxGodpQX+4hmSjcUE3P0DMnKxJAYG2Xv/j1x80zpBvWLSyk1tLe5Sj39c+6t7DZZY++gLL6sy90r
4cnI1YC3eqv0/hzdiFjaH8U7Taz+RCxmO70SwobtlPQg+6hvVkXuAd03AJ81VeS3WeIBzWaAC5kD
4isq8u4uu0Y94wG9SbytjOcPC08t8cvfzKOJ7jYQrRpJcp58FnGQyQoECfTbv5mmj9okWOwfXWF7
fohMZxsWywOG6Jzf1UTyJcCHWhQ7ul6kkMITQkP84aaDrw2eyJhO4OVRGj22WE3Nv4MiWLDmPVBo
MFfw3p5Z8tFKvQ4JXygy9M8cXoVntBG0j+mbj7smTGVfc0zfn+tH/nkENExTTm4pGmpXoKaJnmSD
b/Y88PiXlpv+6J8OShYwB9hDn/e+5VY1aoO3JC/R7iXiaB5b638LAGB8z5nUe3BPBv2EcRJvnpSQ
wvXzknTaiCI1/EFBogRKSKaWXAT1CRhoLTQJ4Oz1gJHSF8Z0Yu69k8jw9NdBIpg+RggSKZo9pfqr
ew1LCkfv+b7OaEPV7R21shoFK9lvtrZMmXJe2PD4VxoM9EJEBtN1PHY4ei8BjNhQs15mULdNdXdr
ospClaT4nDPclZroK3HQfwFSwoQzxix8xFKxNw7l1yW5hhs5r71OcVm4JThUvBbMBKVPkQcFOKcN
vpQ2y1OwnswU+xVASco53XXtOM0KxBZJ2SImpfZGWxykn7c1iR87VWqo8XOkBFcELEKPa224WLoG
yWlM2wLWghGTgADcAmKEQ3aHYb0+05Fr12MAFivqnALytuqMeE5fzcsmutT78xT3Ykw2f6krtq/8
BvfOkku9juvf4bOE0xYiiIjIkQdU5qV4JQ8y1aZdvGkvljaVHYNEUiDHF3fwNIMRobAg1rs4fEst
3OjjTJhzdDjzVxRWps0+Bq0+iwIJ47zFu1VViLaZv6rFsGgV08pmwCzhtuwaQvZW1s/iNBc3tkJX
LGmqSgXo9vDXK3b065PK8ZGKyqHFmmYwZkUU0eHu+h1IkfCB8WxNOSFzPrrYzW3AlaRA4J/Qtp0T
3ifRd0gFz4Q0qjVk5DodZ+rELgxk3M6YFRzak+QbeGKtgGHYDoMqO/KdnsIA0jtL8ekEzPWsrR3G
NpIzZ/RFtOK/lMsLN8E98kiG24oKiA6k5HWu3pskkuSHNFFITwKvBo3FZORHKWmKKZ3bcGjdktaG
qjYKITpG6SLySII6aAUT/FNpPKstuvHNuWjTJa8brvaEVSwqNtUnBRUxmBxiN3Oc+D53UgRZHTOp
SbmeBtuMkW+8BPKAYaq3Q3huhjqogZY3Z4hk1BaBvPtXGwxVSm+vOeJ7c3L5Yft9bC9/Cg4CWF6j
qBsffwMfnLqKs0SlMJwa7S7mGsRiubrg3obSH0SWECScvK42Nb/e6h0TceM/xYGehQG9+BVwPlQc
oN53st+Un924W4E2YfG6N3qnumJDNaQDR2XyoFajxjfE91aQ38818q0GGErXs4WUvXnLc6KziOrc
8iOQKsKC5yHOuPT3dYSS8bYMdkxqh2SVY8KvPFpY2gdILVWWMegzXXkOyADiP/ACewX2Ci+J+wX8
0tXUuWfZ3L4LYtRwuo7wFKJceAxl50tEXier17A8FRkQ6T0xGXdJuG7kPn0JM9sza1LlQF1Ivt+Q
oNlHeOFV0oTWtKRqTZ073XSTJY68lrEnidc0Zl0rn74IR2U6FubwfMRFXzlBGFZSpy6KVhwNSN08
kCdHUGlSlrGIbOFsLmImNfR5oEiJu4ZnM9ADcoocWAJAGkCJcXacC750iJ/bPJz/JJop99d8YRmq
fb2ovjz/ukbY7k3XNvo1wcGWt1EKJUA+dcYS+GNkpXdoaH1swndGzN93wn6Xzn6++vcnou3Lpbxl
FnQ0gftiyONY52Be+NJlUSXm8QtHooYKFiTo2TrVA4gawdZ/5tMPv7iiC/aw95wxwK6J0IrlQHVl
4Y48qkuAU6Hue+SW6C2/TuN8lqTxDLTFwsbECISugHjDwbT3dmuIdzy4IZeDI9juhsM04JhAXZSH
QHTh6L+a8sheUpn6LdQ57gKZsX5OYxUCUH0L6cJ/3GzGqOT3mT879AEiIvr5dUjNeuPBz9BiiTLO
Dq/rsDO1loosaB1RbrUjYeA477jbgM3416d6hAAYn9VlQcY6H4PwSXrl9EtA9vy9ty01pYVlj2dF
gv+s/+7XczSWPLKzgdkoD0U1sXoj8M+g3xO7cKc97k34Mwgzkz3/JNentdazLTbjWawBh99lFs/C
9es7nckns0LP55nBGUBjVFBHaAK/J1ah+fhBoA6QfAqzpoLwVxydS60xMsSPSskMpaj10BzJPCDI
gv2v8Yr3zbjMAxbB6CpjoNmwP5UCcwZx7H+2taBszAWUYoodL7VW44QhB4aAWrvVoLHS5S0SzgrQ
UcZ+fOTzpgRJPXw6V5IWuXXKsa9vwUW6tFnsu4GWp1lRDW9/AIjCN/mXwxBYxJow2USpzMv0JynL
mmSGb72BalrnRedzDJZG1PZ/a/ITi2D5UftkneFrsQrbohJRju5NP5huJK3PxZq0Mw==
`protect end_protected

