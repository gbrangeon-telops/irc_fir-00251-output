

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jmxpJaVr346lkZ1a+LoDVE1gRSFGUifNjtRZEnGV0oAexMx3qGrmrMofcjVsktZm1VmWfXDcztXM
2yFG9i0kgw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dOSbcKbKyGmwastHjwhWcvg7mo0iC7nVbxSBuuKDePvzqRHFROAJKKkq6GTW/pekpDi7EYOWgoc3
vu3a7xd2BbB8KPxJrQPbDcHKKLsfi9Qu05pG8kNfZPTmVPdeph29tJwJuOY3Bue31aDGpBx9n97J
il8TNCf+vPPl3qN1O1Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oj1u/InDUMUdQbb5KKzCbe7WKv0Q1mJ0hkD57NzdtON+OYFVa+iXuwhtetuyEkD/RFkOZub0bzay
EGz9mYS8JrDX4uhqviZ/lNeQvlGcy4m3aXFV0BaNm28dZ3yofXU/BObQHMb2AJcvSvAG3+NK2bRe
O1i9rDUCI7L9zpBAsqwfaKowW/ytJpmf9i24R0N1DPpd8Du0b8109OjIyuP0B6/WOaUz59+u6rpk
YBt+RO2we5Eynllzej7EOx457Zs2AfpyYb/scT1J2gg+ITQOiXue3l6rpuOlPDO2s8UVnv9AEDol
dBES1PgrY5H3iIxtkySbQdPn1RgrbUXGoP3Cyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nf7SNu0SV1jFULe1qPx1Us0aK2tBb+6HkavjcQAOW7vm2bkkBw9TTTcBYW2ZVktL2qtI4SdzYqok
Ur+7+BvPVL9Si1NxET/7Dtm+YCiSnZRDjVxRHT/nOJoMkCyfwzbKJ0c94Mhpx/IIVydS9opk1YOK
norD0fiQ9NScYfnzaaY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gGrec2cOqGtm9E1Oi+bdp4JmEjroHrWUud/ZaF+TGsozi+qUj2kRQyVPKMhdue0iIQELWZ+mxYUS
eLZifl90wtAXYuJxD08Z4LzdxHrYp8+GuCF0avDcKZR6UMS6GdOF0ZR2WdDmkxgQdaVnCHNmLABF
3DC4E9wBUl1YKYXSRH2xT5Tm/cD2sgS0Uobvp+lTtO/g/wUBgQClX1AYzm6JvXG56K4a0tlrJqsS
O19bJe8ailtvTRagvfU5lh5iVeppPrENq5fwhz7scUcyvohRe2r5jixGcPz5bVE78eEpH4EwzJTz
GDGFrWw8qJ6s5hJeVjOB9tgbpdnAFcvyrMEGaw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16464)
`protect data_block
W/ERjDkAWBF9rs4eYcPWPQRu06ckRwLgY/HxwRC26dYsWoYzZrE58He6yQLSLA2FGAW9sJsTmiTd
OVXoHrmo7esJcgePoCH4+1v3jz1whHaYGYVsBe7peRp/+B3IVkEB+NIafBcm075pJTBlCASnyefz
bPo9Ro4FkskZG1HN0T0SBbT3Ca6Nm+aKwsJDrUIMPm5QyGTSMdpjyXXO1FPWBvHpI7KsL69Dy2a6
4hBTS9Z1r6OsdbRb6+Cp6kBT2HB6wED/dRiQa23VLkuIAh5TJ7YkyHclRccKb+PDL+vLPBMnlGwY
LI715TvZMINM+Y7Fsc55KegxcR7TRZxFFwISn2gM7114Q3I8rYVIkREJzRcR5tVc63mAJkHgNZuo
n7oKAV7aoVx9a/17rH/xQP4wwC5YrKySNvPu94dBFXNJFoQC7PaWf1jzpGw+7Bd3mNmh+Z+qBgEf
lc/xUiNfckoe0Rmuy71XNgPO48l71LZ6dmPxjt4PVITRrcWwKFW9XgCK+5ac8QS9c4j5BKnlDaln
kGFCu5Ldugom9MdB8r6Hbw1Kle13lMQ116diZCTrcKQRyYL3Mt2ouWRyhxklz15EXYCU9D6DhNsM
pjTDNGfW4Yr+VPaV4g97EXVHeSmbrf/j/K5PEGDKBBn5gLDsVEu2DrBfZQuWMD/sXCbqBEiiowhj
q/fZWAEJybbhcpkgeA84fPk7mfKKdNnAnhqWTFCzQx/LsoceOTE9uaCRz733zvss2NqhRMKuko+8
jy1xJrbVjz88x+sezel7On1ZDqSv0rok2eEJVG9fPTvJCRS1W/5VMdFp7ud5nIHlgNdM3wLWkEKU
6n+v0E9/dJNBqgDqljcjCK78eO7rh68cizcP0I/8hX/AcYrve4aE8FRIXGyFO4oSkURGCgMncn4Z
Q5UO9CRFcTIjxkNnPoyLfpanB0rFc637HCuxp/xqdXloNp3Qbc1TEErUqFwYPTsdOrZMHrtBYaAO
++Mhe6V/UDd3Q5OypfWuXI/1vY3b7qJah1hXIN+Kkc/sd6Ygf0hUaeFgl9GFcNVBktyUgahR0tcM
D5ftQaW5lVMz/GdvuKBp96Dn73AwB08s/b0U6VC5oYGTpChs2srQrcgnxRw6OkuUeUReIMBuCQPP
2diJRgi6DhahAYoVoJMV9ZHPdbpLIAnyFuO0/5oiuVVu0aQQixnccgiu6nvLXWkwvFe98+980Uo/
RV2uOfVzHDtZR6pQ/uyeTxp9PpdFKzu2l3Avmp71zoZ3zs+CN5I/G40r6k9WDOSCi1KxVKOOeDHh
zKXoSzkKfpCk6d+mOiYs2obsAebPuQudizKOkxMe3fVA3V22P5zDnoj3CKC9tRqZxzqRP0WpzWvB
AbYg0tuYEGTQ+iw5z6CuttCVqpyLmqv2ZPmJfRvC2w4Y/Nt5xiNm0PKJ+9YHgeJjS8OH4YSGx7BE
t5Ecrhgxw7dJtLsyY8td5bRHlDnnuvmL+/Oi3Xw5M99oy5zb2GGQ3o73YWvtpOV1x2PZFJ+EXdNZ
0lcgwGFCIx9XtV75KfmLgMlk023IOweowEbkaJrEl80zG5J2/RJ+PYS4gsQ4F6sDZjnzhvJV3q/w
z7zpImux6+8qxNybrwr2ZhXnENvq1Gx2viXILPgxcu8F8/u/bKnowI5Q5v4Ud8R7HjRF+LfRtE0n
09SoLJ1DIm9LRHjYFeC1EeZ9tM27gVEY6WElZnVEw9eb5LKK6ukETCDwb/BYqkVhLGtxQyT/rh2k
K5JL78tLJrxlGsuAynUMgC5xH+4ydRXzsDTST4wZPydD7SpttMGjeiEbsAcktSrRKFMyu44aHurF
OwlXYbF7yBAD33Rv6t0yPcKUdB/2VGDre37kAdkwkvxWMZqru50YaxRPsQlq7MFZI++9On32FjuZ
j6HRa1ph5B9JvICsbsR5BAEEooA9p+3VWAciDTqm0xBM7gMftNxq43v/+Gys0M/EOuGiZvkpMX8I
3F23XsvQSFmPvlr0fO4UVM4CdP+EpGruX+J24f2K29p/YpD1qr5bT1WSS2AZvCz+JSnQz6JKJJRc
0/4KLZgxgwwTZdq/tKTcscNaEnd5PzpU3LB5Tiom/0VvqrX068vy7mmaNEzLOGmYsHM7TgOYm6vU
4ZSS4zLaqjjq4sgHxTV/Ge/uYE9EOCjBGVd7NPONCNiTGSJ+1RTFE7QmUS6Fo1Ey996W7945Nl7h
ufzr62iVlny0+ol+3e590c1Hr0on78ddrpJa0uSPRnJkbJDZ5UrAL20WX2ylooKmpyoYsbdrDdR9
fbe2Y8PVMRkHBNiQ+n8sQcfFRy8lwAZy9n1Y4+nsfWpeXS/1yYACaISXm1F+aqp3aMkPqVkia6Ux
m4lkIa4zIGbe/lh6H1A8RQLXDxpFvzeXqWy4mN6i+7ZHXaVB9POcprKJpWVWMINbVcvGnVGoCc8f
EGIbrBN/OwRN5Dx4Mb/JfmnxzpDtTSXjUZ7o9IZT3R7Q1MJqo03BXg5I1Ddht0lZBczo2rZVPkDD
lF2Zyybo3VBgJZYE3p9f90sDK1dcoRkdkEhA0mwuLAK3o/Bd9aQ2wuQ/yp84KIeJN4cgoW8zYR3L
Lyg0+UUi4trhQerHybOnQQZXENBbTujtG5RLnOCPWM9gc6hPqAUFNT9mZij5VxlgioNly2MtyipI
oSjDNnW4k8NYAqX4J8uApykI9zLUrafHdDNQ9coTysZdifSq2PiTMN85aXcL2trXQ1e8rS1aQKs4
SJU/yiY0pQOP7IBvqi38qESaRSfLgVQHHfQgUAax2sl2hiIQPEeYhpetLqm2TYfvp5eLoso1vhvM
zyF+NA8uXdH2C7dDmfJcK9pBvJtaDcmYWZjXlbc4GK0kpNeg3wTzFOH2sxrqwUUqjHWef+kmA/T9
I3dGzGQtBStF+IjkYV/ISOw/CIoXDlGvBYerWoqh8+PtEhpZT73POvsJwgFn1j6cZgAJ8TV6jnt1
7cKf1oXKRZ8XCEH1mBCZWB+T6BO1STBL3bIMVzkQziylfPIDJQPHZYV55B9mHVSTbO7cQ0Xgzc1h
nXewJ6kCnPLHjcjpZB9sE3YBY3eWrfdGEhDRBCRLsNcTAmyPKogRHdvKSr+2OVG4sm2g6dWQVXI/
LsHGINaYy4rF43+L1QYcc18wm0wiUpLI4xSrdVFBOqi5ILRtFXMEovMdMx2KkfiToyCTX7eQuye4
jtCW81JGnWRdgSoQ9OTICWtenZdYEb8ij33hFJ0lPvAftmYLdME79jDv6+EzZiIlwsXXVePQ+IRw
ZWy5hgNYbhQ4TARnuEDxokbXDsy5b10TnVamW4A7xm6tMAJUylT5ZoBEkHzDEFec9wilNfIXsc13
uS0mWfSvqimRap1r8cCYlxuWNQNDGw8w+2klk3+hJlxDaam2LwFlVii7ihd03QYPRssu0S8afna3
u2Zc3eyY/6z/T5zoEyXBbFFEcFHyrnMK713Cny9omuLoeJdwLAniNQ/mYTRO0A7n/tjzsf+YEojs
5B7JzQwRWvy8nA9E5h/XliguqCnkyw0rvLmJX+2uhV8WRvCU0UVrFHtNNKeXddcGsnMxe2rhLwt2
QXoOQHqAHEYmM+8tdlWCEav5zau7A7edvcW4UrwQmt/MRBG32qNDQKBPWxbtPlvaE5+LwahsS+0C
JX4vfoTBb7oQL0RlrlO+LhIWIXAcnyGW/Dnxu6rq5KF3sB7Gu8RjIaL12/2pRzQppS0GR4IQ2hDn
Xh4fo8AtFR9EO4K4ccsGWzfAiekNjeEloIG/ZIhl2nVMEh9bfpAFMU7mZvWlcBxKtJEwd3lcuewh
Ld9mjkcEm4zpH8uo1aAN7yzyb5te1F0giKVz25CmUCVjvrJUU2Vsd644osIsEfZ92tUm04F0xUI6
QCyq/ieURmgBTY7G7oZicrFimZnPp+25KBwpgDQWA48wCdEpFopRFpWtxt1TiKBa7Av6hrAewTin
QZ7GBVOdfXj/46CtsTGzi53mr5Ic0FWs6L1E/L6QW0u+dRkpwSlGg5hkmYFXAxk5oiRcYNw6Jozq
3Itpf2z8RwSC9IsW7uD0lOrOgd2O/EReEJGeL/IC0+Qp+fTsGPiewDP43p6IXIB7V37+lnkiL0mj
maWcUUL1cNbd5Iy+H2IZ/kQpe2Mg1/UxOmoOMwXiuYySoA5PdgVg9jwBW7a9Oi81xHD6Wm7Iz0gT
GHgLkP3VgDAXLmN6K/JuT0ZmgUyJ9GUDsaXkKvBDzDGavYFDnUKglvzYnNkYLEXjVyzlwwLaEb+9
zmShPZjBPKJglMtkr8PKgDUTck3kFicbsDG47rZrPTGEbAGqcJ9T1719DwClaozN9Kwnpx06wL7T
15V9FvQkPUc0tNmQqtvP0A/MkKbiZZad1xhGU/QN83k3MGZ6weYawbI1+chI3aelCn4LEYbuYQ4Q
WAC+h1GGvmyyo35XPVYb3+LVzzgkgP6AQfTbDH/90GFrZKHW1n034NWMbm/awGmq1WgrutRgsTAX
o6xIiOYUssme+dszULCeEVaMmUDQWaNhvk47fgXiPB0D2vWy5xxefuFT2sARb4wE9MOjCnu2iW0O
lXaqSjITOWa/Dbkv0+XgCztGulcAvSef7PcdmKFuexUTRnwgM4U//TPR98BsJESwf3lX3uA2PmrF
FLz/iECM7lw4mioF2zUczS+H9DRXbP4cMyDtPq0kOmdvCDltpgX5UhFN9nt5e/k4N+f14xikVPQI
mSY+gdUxKSzojSr1EvIohSTAg+LZt/3/l1J9GJTfwDyjtI1J8LeRYUP94Uefr0KMaz4zyylS0Lak
LVMjDlntNsuRO/19B/Iafy3IxhCYGa4aRLpmFy2X6WSoWwZqoJGoX2hTXsyFUZkJS7/vCfD5Rqce
Bt9NKsBYBFCEZtt0dxUA4s0ZaQ1rETc0e8h3LCnhVLHDyELiD5I/FPXy5qnt7D9ja/FwLFnVTGYb
3IQ5ntWve4aifOAnifXkBxrAU55pV22zsSWkiS8cqt6BUZ3X3ukSuO8ah5EAqkhN1byudZRK60Xl
pBuU8afMZjBKmVTqOvz4J9LG3FYNegitbnnpkOIXt/5t0BV2KipHIaTu5pMtnj7FoIekhwHKBmWS
1ULCGuSELgU9VNTg7EacP2webd9/QsdmGqsi8a0w+Lqx3vmBRGa4d3mrPgLKv0zRfwdGDVuU8r8G
C7DIrp8tsEm2gpIJyCfJOTnJqE0gYVUXwKuQQT1LURMV53Lef0oxN2vVelF6LEAwnsN5Ezv7IAWZ
oi2ZBbMYHi44c4/4cInJ8Iva3TmCy201a/sBLFSbpefLW0AsvKJ8EOnJXiGKFaI0GxS1XUU1GtbM
wuXbgdn8MwLNmKeDWmg3uGSacjuBIwBPSXWNaZ//ZibvEhqEoKny0KRUBEstrMByTo/KbSmh5WeR
km1k/dv2VR9FJhoC2JEoruYBunsuH7cyDjGTXQuDgLhdnOZXHmjQASYwLO2d5t2Dc49RBNevazHv
iIOGYEzGsDGTqZIaz+X5xcHKXlCgHmLqU8NQzt5Iewi+DpgpFKmzotDVDgTKEZrt85HIu7US48DF
DE/QR6TT0vVcq/qAS+Kd4kLcED9le5R4ERI29GmTeiDKaa4++zTFyJ7EkYlMQn8sJ0Cho0Yx5mcb
LMewKlpzixP9AE72LDqQ4O8Hws2M14X3lzXzMbC/WmDXS8gCN5JVyUtkykoCwwJH8N8S+mUWsttr
oB/T0Uw+nuwbHFL4PnScL2wG0yw6IgBRibhd9I1/iad5SBbYAXMTLFuzHq/pkdrGtjYDFdWQ4y5i
AdIoVbeE/G559OmmcUbx/7RBO1xRhr8JNjT1xMrhX2SmpjwbECVw7qFQcnMflmpuK9aRSCEW1e32
h3W1Qr8fGv4vziWhPAE06hrhuX4S94I1M30rPCyPHCVLWqMkU1RU1SPFrE5L4cIoHcqzi3VtrXAS
kPsHj/f1f06AiKmg4b0LCfk7SoeibdGkYimunQI1X4tJIAx0jmS2N+yWJnvsrLlQRA9C1ggwEBUA
jh1JafbZ/ihDFh6T9Ryu+EUk9kBsa1S8pFj46lVG07OIxaALzBp7dAwfC6LAV2zxeK1C1N3E++i6
My4Ereuj5fNG570PFOeC6YuK3JyTAhMZDmieBmKgGk9hNk0h4bxDkJC6rcnhWqC8phiVBGdV++12
yrH2DyGsGQKYSLQ0gcoEeBL9JrsMt7LLLvKdLbbFzNcl633EOq0tDggocwQbLSvZhVp3KQnAz0w1
tWz00BpObHHxpZsl3G7HUCHjlpRBpGgm2dRxI2BafFHFMHMgQ4LphWAj5ezV7lh3067dol14woWA
bd4vmFUCmTn7dclwXXJJn5YcxnEMwDJYuX14gCwZpJvmTGH+WuNxsWSc+SEtkzXWee2N9JKEdGdB
SbZgoUB1I0D31LUDhHa/zd0B8GiRaaEHjRAQxANGnZO+BN5sbzuTNYLjU00+s1OykZ6nvnWRoRlG
rXD6wW7jAH9M/3LL0j0QQ3ZdtoAaRR6mbBKaqdlKaWP6oRqvUyhEdmS296TxZTuIlHHZQLFqQq1G
1Yp8j+Eklh0bc0ge4JfqJH7uKJeky6UDz35q2/9VWIbb2LIVacMlNMB6+8GuzFjkBVtWpW7/SnM2
i6NuGTLhLeUaNQmYm1eZuEZkjMljuw8kaWUAAwMxnd2fvmA5u+gQcKL+A+43kp4av3sz0zSIfR7y
bHj0GETZBPcTZmVM1MRK145VnF9kPWuSYOyoZCopTstdtndQ0lghwxFxrDerIwqwiAITbfMw5YIb
yDWKdToQOGL+iUz1UzsAH45Y7QseQ0v5c5R+FljMTdmjjCDbqyAVLqnuK7SLtASPGzz4bNYJqM+3
jPIG+jURf02UxLTXwJZ1ao/Rw1qRmldZl3CPidZi/bsKPXPd8REPgRY8pLCZ7Idx+kCUuNgBGtde
2/MLdDW2vsX6bsCJ9WsJD4FsMXh9A+DuPedkxmRHBE7WBtjXLc2E83V0WiQp8ojTlOqvrI+RokXE
WiEPqLZRqakydU71nr+plnVXVJhbTtPnGQEVN5g86PTb4R19IksmpPNI//ZJnqLH2nIe3HsOXrDe
v1lSkoWSQw09r/kCKeIssg1oTjXmDEb8zeFgonQ21oZNR5MVIRPee3SpIjSg/xNX/WeSVTkJjWTc
jM9SZ28KoDGd0mnuScNyZdh+0AQiXTfqU3llLO2gt0wsSpRQyUhi3zlrhAwPvdbGLN5FRNjdlGL6
093JI8FOQzQzIrF3y47RXwyN70LtUfe+AgHTkChY0qfFW+zxfG1ebanSP57RNuU9VeKF3P5Cd7+J
DLFDJM6PGSYlH7ZOJRerXQKp3Uc4aQmWL3BuCGzJNejOBtDWcWwOJDjWHeymlZaLX8QrRuppL1fD
6pcYrEHJoPH4fEmuF19f4x93YxsRlZkPCIZRvqcNKb6IyhORuPBzE74jMVOF51dgjZHJ36a5M/Sv
wjr3yhrXO0vriy12IyYgOgtZKBbRyHGrdmd/4edFNJm2RljKS4hCUpxTqdW3OPr3pe0hsqQjIgku
+y90PaVxWzfZh/MdMhCtydfMUC0QM0ibPriZXblEJ5CnF22f7in/l/PdDlzYaxa3WqX1geRczBXD
T8fMCfjRUlh5s4fazojIc1fVT/WV3wSVrTQRoWrE1WGEOWrKhApSXNJBPVWumvm9tP9+Vjo/sisS
xtNBxcqxnlUEJbv4JDIdfgeHjumywh4WRejqIoV/aB4DgPOGLk1XzXWpLWpoyal01+G2v+WzV8Jr
JPHV0cXKccuAq8qF6YBSfmaHegY+Mtsop1hR+iVAkLvPJnW/evaRiOYzBEDPYkRHEby1dnIFlsb0
OA9rIXQ4pcEuWWISUg7KFSw4Bgkim+yEM3g3hIgP0SRZFj5hPgmHn5Ft+qqwXucON1xRuB5fpOaG
0X5FufB7xpDfBsy/v+hEn38oIZ+hxziv+IGZyjp9+V2vBrraIRmrS/wMlrpYejkaFG0rYQ6b5bHy
vsVinVRd5QtiB6sJcAyb0N9ItIicvVA4Uxa/ZWpcOFCQLhZlK5iYei/mLI08fnswZjv0BMzrPkUt
/Q1DYI7v8J1BSNC+BbH3RLEPMDbHjUvouS1154UZFrsgdSZP/6nUUYi0X/JbChtzDxXgLFm1kdG1
wi0qk29bP0dQzSEsHrVso7rZCtS/ZI/TijWs7FRxKykgjoVHqn3lkp+/RlP4sbcfwNGk8IZE/DW0
xjw4c8+Bb2r/qOeXa84jBgueVcTBCHeER+O5s5WBvzz2p3DbLnlnnwv1o5jV5Cj5zg9vWvq54tk1
87XxmD/j/K39wqC6+ycsqA+2i5NuGdyGgBC/RfaEjVuYk6dmgOj2MddX1LPEtZTr12Rd9ZxnRNp2
7pWlKcCV+B5ntFOzlibXj6Gmjl85fuWGHABYHV/UDE9NX+8DAsZXeESX7a7m6w+7VlxFG2tHFWts
Lr3+W16sbp+zPya/6CDkKNC23qsqyV84s75tAfZVR3C4tVKfl1VP1+KglvWIq3FqesfnGUp5CAtH
f7C6oDPcrsLtHV+HqH2rwi7mla421REf7RQ2rkYRfCtnwebKe8f88H6VOiPnGSOdlUYhTuF6Ga98
C8KJAONmsdLr+4SvqpCIfv3JFwxom+0pnxtWPFxmmqT9WJQJ5R4H+WerC+TZc0tESlh4dd5XtYkA
QycGzqXtvRjkPbSL9wyzhUa8RvpqsU6SnkuR904a7H248mLkZXhNrWjz5dBOi70Hmz94iKe5FG1b
tNVlA1ifoF4iEYAoVwIxG1SCKO1IZqx6MalKRBnCPEeCDJFzVH71stOU3SftmpZqatzj7KGz0cby
5I56oY6x7l2EyyqCUBs9jOZiD+SE4Chl7ErQtBNSc9O94DE7iCHf4nNMuQf+nJw4qVXoLb05vVI0
WU3I+y+u2CHU9tVuw6H19fs39AldF0CQWFkFKOnS9ogNoFADmTvQNt79gye2JdlOobLC6x6cJMqT
v802Z6HqXb5WGO3vNHCx7t8FGdGuSvVXClb2jlhkC3hMdihOlYjKqsIceLGTMbrIzW0EeT9kyUvi
irTCrrkjtnwCrcNA/UJcbncAW0ai7uwYjduLsQPPC14YauXPOvUswuQ7pW9HQqR7uLqW5zwkhhA8
Rnnmn/S3rxFuj/qDrflHqAQTBzs2EEhgNIknoG+SlCf8XXvl6NLVHhvoDqYHdYUR8uQHkRBMYCm1
2VbHraMX+6N3S3eEuQRF9bjFZ7nKE9oeGKgOvYmX7IYR4Ly6++Yqhgy9S14spqYZC+ZkBuIPlAWf
hWCpyheuYbSUmz+4c3O2sp3Mo3X3buvMjMno3LbDVh5+YTmooqF1jXTQGW0VncpafaK/Vl9JVpcj
d28UBpN/3XQ6KV3JmFfgpYgkga4zidKTiWMjmnLkKnJvJ2sRzZjIoLPaNCd6uXd2WE85ciSwGTwO
vkUR6EjEKXGoTIgwIUyNJ/91rZf5bwilsl9D1Q8Uo8jvVTmbge4pKmHZ3AP3/X3qCwbzyEE8vBQW
Yz+Z/+UqZgWSBDCAGWY/4mQDei9H/KDcYKgLUSKpvNxTdgq8pUbNho1nXRWoA1YnCTjLLUx+IoXl
jiz7GDiY3YFsEKDX/2ZYakRI/cp9AnqDwr9/PGhpNBBGWx+8EGs2gxhNOCx4g+dBw+PKrw5iE5wp
ii127VNWp3/U4HJJhuUHl+RqjPR23VK7gRm7tx9GaHzEifxB5/LyMh4ouKpjq6HZzYxBMKnQJiPx
bOHGhZDLf+LfypA/jFm0vgQg6ALhW0dtqAGGs6XAALkDsozIVJ38d8DeKHPX7Xrs9CXXFjFOUDuS
mQhYJ2MidFDNnq0NyD/VIsspf8OjwdPjD4dO9ywA0RaL3JfloRMVzdVr6B4zpP5ClvHmaliaA/bz
dI91VDzN/eSWK42qLa2xr3C1C4OlgdvsukZ0NWsIeOdQyjJI7VDnh6MNKotPeBhbO2ljrQbqaVRy
mRtrQEAmUjnWbEcKqsvUssMHQa07/jk25bHqAaazhWDE7ezCboSKTZ3aQn/nh3GXdo1AH7Dyg1+N
ESWEDteeexaRa7e85WvckTIjHmVBShazVzLtr9FQ758p4Z03OmYk5l4Vv1xN8nw4n5rN2XXRdwMi
ZO/gpCLif/+/aYdTzoDcwg5lRn9vsQCxEHX4NfUQ7gMQTf8klta2j/N8dTGwGsk51Jv0OPEtQX14
gzu/vfN/RmR9CgwcN+QRRpBUVGjwkQncVGqITue62s1/h2ShBylP5B9/yQVOXwtGcRP4JHMK+xfc
FRnbWPd0kyBKmFnsdSeTus3aTMZrlw/rgqAZgxS5yKpNvcSBz7RUs4ztnQOF/YzZiPctJfX7GJgP
NrAzeEzWyGGGRCOTSdS1EySFWVgml4cOzo7NbAOnXl1AkRiCN4lKQ626coNDrjon54wqD/qMcDPL
aS68XyP46vhWdSx/QBFSzedLZAIfjsaA6wnEjTPE2WkeMv8d1eeBsCu4Zm6VT5XyfLUvhEwpyQEK
WMLuvXjmXSBOH15BFzdvB6vQg+9L8TZ2cVGnrKd3ADzunZ0FKZQOnMKHaJiZxxyib1fgH61N5ijL
g+3ERv7tY9Spua2y78Ryj+nWoFE4u8ScvBe90V2OPcYCMtVuCt029ilaiqN7z8pm/dhoj3qEnTIs
6KmurO2NmOzLJzVo3neHjDybPthgxZekUNfLsgEdbIeXA7qpGqWLY6GzSeuxx5OP/eDylAvu+Gnn
Wob4xlM1rqHHA4k8CKIqoBz8sbWlcqozibsiF3IX1S8AZm6ZdAMDp5zSUZN3DkCUPY/2d2s0QQGP
8zF4fGcekDQaqz4rwyYjv7VC/tLQehBYb1GxFRTa4oj77+j7evpm6nbywaHFHsYc/cXRwCTl8y8B
Rl1oUcJWIfYgr1e6Q2V9HHYRhNn15WUe9C0WbQ5MAGoyeFVe1HRAt3qPDI4dfqay38fMMM0J/+n8
putNgF3ksR1mHZze4rcCs1kPV14sxYX8lkzMAybe4ulrwUitaEtvvrY+OHVHQWlzbeWu1S5Sa4Yp
qBaoRuilTDFAdL7sL0dRWiZub11MeAHwY/nyqQnHuLRZSWKr/xNHgQ1pNIVf23qjWymQTbOLKbXb
1QUZkukOKlbcyKnLeqffM0AhBC5mAFqcueluwdSwLaPYfdO4w4bgKQ2h5qy39csSi4LFA+rHfuMM
LyUxs+wzcn7L9K0PMVWFNuIbpERmdwhEyZAIBvwdQqXkVh3ZvEnQO0OUi8cnBjcyCJNbarSNF1W3
pYbPXTHf4QxFcS0/g9QlfFAMfR/vnKFjJiPE1b0x+g/mIW0RxKRtFcv8w/ceVuK8qscDJWW0qGC+
XSuRj96gEjPCWp+4i0hT2udpcNuR7Vfw4RZ9KcO0kGTGpAifwU+YyOEaxiw/FdQB0rSGys/sKa65
dh9UsehvyxDzpWDTvGRBXwkvOxu0e8EDE8SVaDu6qkUaxqQJGS3tV6WQU44bU+mu1gADtZpaGcp3
eE4bkMCjHpPMnn0T3mFMiM/KnIr11T5ITxqUbIThJvRQudoZFDTjVpDRjtOSaUdKX2D4ulvdLGgh
8KRgTdKFRS5JiA8m1n74P9qlpQ/haKmx8GeIMziRDqnhvcxMlVwnPSHiZGZDD2sdCUUIA2j3C4U7
P0uZh5OKoMRl0DR189r1h+rDi6kPTdsBhmmIVZtyIsc7AoGp0lIDCyiOhwMuwQusU4mSU92xy9gH
/MBY+CVYPG45bOKK8loHqFbAMEdSB4HIzxOaVacxCwZe/yDbkt9DUc2L7Fc8KdM4z/xfg2SAqtGh
209D5fSpIHeDowglN88ls8a6eIXQa6amqMldOzOqzZ1FEvgtKX3H0GqveobAtvwc2Y8Yb7MTUCwt
g78oX43258jEjhvaJB+cO5AzKn+KlbCIzTzP/JlytwlimWA9zM1+e8PJ84roqEz6TOoKl9Pth59V
ip8qs6Tq84P8qk+pStSWgIGrSpgBQJ90zB1uF3wsxRqegvmiKF+JxgW9b8mgZwhbs+wCD9vPE0AR
OMNjQlPdIpwkN+FjywvPN8LBC8NEZi+mp8md16jbzFuAFR1Pm/HaBowFX0dESSljgNfWWGBrvHBW
V1IY2Iroz0Wsrup45X21h/iOQ+5WtK2ZnlwzykLYQbDs58HeKCriLw4i6sGmu59jzZz1lUsw/fOH
6r7qVsXjgRdpKNu9fzWq5rWMBDKEuC0P4O+ZR25o93oTewkfqN27Q+YFf3q1XNOSdg2eh0D3dSa2
mGIBc1b7WF3KNfBMLiTyhNC4LSc+Zo/yiynUUt98Av+BMpI/Amh3wMYDqFcexPtVxhQRimb7TwYH
Hes/F8gjSqSh5CSVpv6b+w6fPXUZ/9Pcvm+HWE9AQoWtE04GSJ2vxQnTfAvtHtGO9vxshhWT67b+
A9reSm0hPxSTreEEy9F+dYD2URILFpeDh0w6rLh9uJWQjd5regRQrTnOpfdl+jJISFgxaAlqbJ0t
IloqVEuYT+Y7qejIugqYHl4ovuBZex+MJPzb65mthaKMLH/cVQfuZ5jkoZslNqpDDZv2yF52uqwW
q9g6bsn/IM7ALyuzafN8U39Hd8m0hb1hOO2sHbY7mCGRjnQCK0TvGbLlCfAKAIkva/Ndk/D1rXz5
waysqkQZLsOvjGSfBafj/AmG9j+vNAJY4/RxPe+qFoMslrxnSl/y7hzu88cwwz8m1eQ3lAgBLUyB
F+58sA3PcdozR9FnuwvzXiLOnCUWuDfcEAWaLLnj7vaUD5IAd2KmlPjcJUDaw6FR1QC+EedjtR+D
6y0zmfIXgCxQB0HyE4I0L/xDSjTCS+GkK8lb/jmQQGWcaju2TgmcBgTdgKdkeuhEVsxgZxIIjrH5
uY/Ts5qVnzefcCG2PTIyxCqq9yyH5cF0SL4OLqnk/trWoBH09w34C1ZiJ78WOnT7L0wTub2cnCHA
Mr2zntYZkPSpDo9U54nnGWCzc7GWEZnuN7b8zaVkQ/y0OU8wvr+b8Atgl6r6JMplngN5Caq2sK50
JvflyqW19kXRc2Arh7ODW31dUAeVTTidNIDFwo9p/0LG8vULYmuVmAR9AhAGFDD7vi5aX2H9p2mT
B6fhbjUpGq5ITrz0MtiGgXPcN9DpaczOJGiZ+1IyQnDTd6Iy21wTwBZExgC2LulzBH00CKK6iDnd
nK3I6unGjqGlaEIkr1qmOQshARI8wHnxhbFHdtXWQZjQOFjPouqOQon+pTXNmuvyQkVWrofgGr3D
FHmcX67OSwzBIRBcGfnJupO3ILapXuuBg0SR4Ra6Hs+eE/yi2FfBcV2p0nxkgWphLQkCfM2uax/A
nSuMhhqlBUm/eNgKgVFimOnKLipbZKEYkl6H/haluCBdhA9JNN7k6x07HEMph1JX31+rXRliFvpM
E80u0gP12TKKy6rPUxcGrAr9yQmF8asMDsq8aKeJHty+SmHFEUv8vRMm2PUuwAFWUtmra3jZJcpH
jE+6szx2L3uKheOQj91hP3f85AvhpSSb6bL9jjt3GZ2Y8l3xAXQVBNN8FftbB7fD82V+id2Khrnl
F3pLlQT0O1ofSFHTszeCV8MMK7vR0bD3RRNttzhXMDGvmJqF3mUYAUZ6Ut648ygJtGKc+CTpY97q
VHXz16XPsKBrJYh7GhCipkfiVflFrAn1LCG/ULnV/41QMNucaPPOm+z/S0a6HgxNpPEdI1URf6AZ
bM/exYithPJJslGoxnUB2cV/CNTQ7//S+v5j5pupPK2KXzTA5rcDnfxZ5JHcu5Z0Ye0dA3DEUViq
oXQh2dC+iaUNM+Z29UfH8yAuVBnXx0BGRUwoi7UrZ4hYQYyoejN6VaGZ1p07CMAAGAY6hUO3lGVD
kz/7/Qo1CHxxUzOM6Aqh16XjPqpm4DJ6x0fpMWgvqWynj1Cu22s+1LBDgEeoo9z1JVbZivs87oLH
RFbS7Dk5IX9i0oRsl4oc36jn5MnICi6OJqBkDOvu0ApncLGDt7WJIYuzDMjDN26n7uGP/7Ket/og
Ti+ZNNsK+7cWz8Kw7sI55Irh3IS4lDNdg0G0IW/wDcsQdLTZ4F+A+11JTG3fisM7E09Rr6OVv4pR
tcj4ecSajHXeaXbDzaPfc5pmuzCi9OJJnBAG4kndh9NY/pE38BzrpvOh5amBOcWqPr5r+eG6Md0I
xw/FZoEdyU67PX7+HZxQd264HlNNRlwX1iYKCYh1age4iO4MIgxigg+fVYk+hnvToNVYlvL6NxYj
aZOYq/1cGpAkHA0JUcIR+yGqKnot5vnNtlInQnRq4uM1qGYU2sS2sEfQLkWXW36Lkilk6e0ckdzO
OMXsOwmECuyD9C75cnkwbITR6bbDgw4n4ObtX0s7YwuIKUAtuW4odq7WO2B4/M2nnlNivOoL8Dul
2vsuUNDqDdCuzdUUNK7NrGiiwT9ND2r0ye6kHgmcGk4hVnTxVzlmwAxqxlhXq9dcDolAvA0BsTZe
yDJV45QwKgpNQPg3he1jXP0xliHPpwkclzqwaBx36112dwqPHa3tGSa222ojtVDwQvl2k8umWJbZ
5xpQp5iYjQ0XMR8RTQ9DR/6wq+Pv4iUXsJYMs+1u04Lc7h7pvim060OjqsSZO2HJZh35DZ0+DGU4
j1KeLaoCt/eFvfO+f90iKj3mpjNSq7jzthFGhv4IP1N/cGavE0wTNIQV5inn9pmrTOcIIep/KZNd
R9+hNESN0KbqUVWi/hgTA/qIGxnRquiIPkpEzyV5Z5JrZdTy8+MLe10oje1jf8d4EZkAqxm8B7dz
rnAb2dnM+EE5uC8QY5xV3NY1YpntI/53pae6Eu3+oTEcleGv9Szjh+jH5P+a9g8h0kzJymsCumZw
3cbavbcKy+7p/hQw11jxYXs+MSbI3PcWK6k82FvtsDv6uKruHv6XTFhyinHAOz5ILpxYv7u7AJgW
hP8PkFvtu8OBU3J/0iVTVi6lLUidET4wtBbpvmviFn2tx75WW0Vi7ul6Hw9h3uXrsI3FNRFbOqZP
Vehz8+wrJJ1C3JXXt28kJylbeR325R3+N9gHf18iAFhDkZSPuHwNspdwEc2b2HbgJEdN18Gdf6vZ
xoGeyBpr0P7OOJ9VinIHv5lnlqu/PbdqPFpk9sbEvN0oTjxK2fRtuaXGPM/kD25xflovE8ww1oN4
Bc6VLdJC6Ax1/0aZ2zKBk0SiL0BZgUmgKq4TMBdVHSuXMKNMsFCOUOL+lvlYCSafV7qZr+W0huPT
r0nYbh3KxjoPezQhiNAxBJRBT+bPFVuFiE9SY5+ShRzCw1lb+cAz5VnhxYRfKBWrcvfkVYt5euRt
8RNm1B7oNSPUj+KuIP55NYhdyNlMZ1WFzH4qUPEqiJlUqlCuWfBGcqXIjEtEMiJPpf/jLLt0j3IE
QpuWqbiSQYf0cHg9QNmQMNfxY8MUPspojUbgo6SPqe9gS84uDnIP6y98qoTsOEfZC9WD3YlYXY/M
MqcyLV6usRXDOsJUW1f2CBAmPdHgD7c3MsLTTiu50VuzZn6NxqC7y+ZmQ9OpebVknLmKidVcqgBF
IGVuH7dEiQp841C5ZX+QHEYJFEPaQqj4Oacdnf1S3p7ftj2Yy2FDK11gIO5oZV3bskOKOjd4yjIw
8UnQV7FKCp5A8vraKUd5bIkj7djZD0T+OHhuhRX1HseAJkyyBXx+ObhXyk1tRMIk4+GB2lxfYuAB
7mACu4jOeDsMRhl+LNr1L2k3M/XFFuw2HwFXG7Ixr39K//ZsJNaSUpBXt5gbB81fkTPoJTxBBAGV
a0B5YzpLm1EBgKhHBWD/eDSyPi97M0jV80jh0H0paueMBEfkQ5UrFlWM2sv7E5brxzmFVmkywQfI
+6Cw6z/qGbWwjQ0z890i/qPITUPqqRVgORFQRxxv7iSsoWcJfDP3WFIBys8IUybNlvpcVBmx0XyY
AB8rHQGjtNTH9D+eUEzFXMIOOHEKaxsRgI+hT52CbwsacfChZSyIVQm/6HWODEeQM7gGGxdJqkrM
zEBqnZ5fm+0V+Spv7Qe/zDLCP/TAYEejuCOPGJ2RxD01t3qkUK+zWSyW9f9zgbuMOX2bEPIpfZrs
GOUT/jpE0dhoAyIQtmek7HPGCZhu5hW+VF7r3xnw6/8jYkBDq5LmrFPgtgOg8Fw0fSSVrJ0Nj2Hp
ZYxi2GLE1IF//heI+6JOaCHMtX/vvhQhI/X4ENDGH/EzE06quxSAG/hOkmZ2n7p6U7PARVV/7UKd
+PbVm9kkCl9Ve9yi2ZD/ZSPZx7xKHajtrq0ENX5ghokqD5Ccp8omBmVgs+y4BG3ZthnT7s0PT1d8
JQBg8/+zDBtwtRpbLEfgxuvZq8BbFLoHYzOrRsBkIasBNX2bMI05u8gT0k2i+w6KIv2R4Hl65+NO
o0hQom03eonVQ/eTjFgzuxsw++zknpep0kF/V04fZC1tDGr2hQVlWXAWcuYFkfTGcDlcvD/N0zUN
th3Uw2nKof+DyF6GHo0twOAZyzkbD/DFdeY6mfTIdbsa2z+TJ8oC38YDlTr/cVgme1Tfyp7lF3Uu
rUkcel9lCCe7Or61zjqGHVvGQ5EYxtX9k0R1Kzf516GWzKRyR6PtBCGkGy/aQz2Mc+7iREH1pHMM
O9zcCkfKjYwzIxJV5qYE4Brk+VRFth3fhKr+0CVd9JIJTWz0O6fMcSJemuprOpuX4ThBhFUJsSZk
ujfsGDkq39bk5Q3nmgzvXEJ9etc8SbN1nkQT9hvFmIQl4m0pbwYFrTQH/iuWFvD0G1aehGZAWCpu
JQNNFj0kjYJ0gRU6OYaxc6nrm6PC5x3Pu5Td0J39FS65tdbSMdh+vSaloQ6mT6IHmjAo7wF4aT8S
XgIJbAVqzHYX90deua23wRek+eHlNKJ5Vys/zLhr6c5nHWJt6hAhHjZjYPSKwxinxSDtUZOBpith
UCBYphqoPGAHMB6OxfcKmJQPRaueoLRERT05180M6WgdGhu7w/Ko+opjp6xldqBtjU6ecVhe/SNw
8Tbk0zjyKpeVliKcFU8sLxdUgx/lfTHg29e/cSdl85ks8MlFUQN4vX6Ctt9BxAlC00Kf4+RZwQ4G
EylDtkWCwaynNgjvdUbL5T3qe6r51OCKe6ALs5JSNQR6FeJiC72W0Ydj9cPs6Hg6fC+AdtXbqfAU
n6nlitN5rCLonNml9aVrJ/kp9o8Pa4wX5mmLS5w6fVXPbQDrz3VqW/qUncNfcUk78DlKRGDOlVs+
LEohka25oNyUYLqtJN7xzyJY+eOMa/WPSE0+0DmkH2m0hqk3WRUdEQ4oKvYEmal/t00G7EeKH1hW
MOum49Q6ecKWowZOKOpMBFbJz405X+gZSad2CgPOYRrdV1uLMsz7wDRHl7Jfl5B/kpxWEmjSaNiN
KoymoKa7M6X6QWcKR3A1OchOlHdoyp/R2J5MSsSftmde98l/pY3GdswO5lHXjwxDiHLYlNI46GGt
s3DFUBHp9dGBBbqfEoFUdVBNZexBTQEOS899QCnGeUOCVtHAxVDd2OaYmMy9JOPDgtLKKZNlCxIe
FxtNG7lgcB3OPPQ6WhJDfyfymI1+PHcaUBTotclrrxZ23P0dfpkf1Pe1Tdu9eoq0kQrPWgLskcBF
b46WkDzDKXNgFCNrZM5gHwFlaZ/6o/n/1BxoZ8g+xkZk1Hbgw2dXF36t+1IXed8SzniR7Tp7fW1F
QMqgIQNqFFBSKlKbgbVWgofyIGmSV/dEmfwwM7d1C6S+hdPl5n5wNKf/XxycQotltyoDSjIHdac3
8Qq1jVZWhRUnWMBgGeE9YrFgE35djLO2RJqLdEP2NxhkUfkMljXRtny7xfx/wBIIePzVFdGvDMsv
h+nbpeOuPMo5YmnYAe+NsQneL58V2f9/aJX8v2tI0ekbzimokzTIPfvNajwELVJmamS5+Fn3nXDJ
eWLoOQehCoz8PsXxy0fGsp5LHmyszCLS64WQlsIcLoZO2j91SDrMKQYtzjEEJ93I9UGiCfV3QRDA
I1TRquJketsdnOTZw/s1/OMh9DxGjzFYPEJA3iwywuhDAlkUEr1TyYZoo1EdwHl5PteJy79Ohq8O
flP5HPeOFNfVZHpHVOo9PhuICZUk3dbA3q2n6M58W6YWfxWoX+mAoOg5gUgIfwWRX7m7MDvCC8QL
cstqyEvKZ5N8LvXVYdIgaOEnVB9WIZaXqaD5a0VogcWRXTFcJ8pDgASeMS59i4AHG0acpA9nj962
qUrUXUczRbVOaszz69sckX8ixBkSkrEIFDY103ax38s6V4/WIGYQFGzFLQo09zwXi0XFdt+a51/b
Yw3lict0R8vEQVMVuIH7mm9MkrDKsOilh6mtlsKyZVY0qI0kTxFeICfgVoPTMESgQMb5x6AbVjQF
T/eYpa+t84kHJ1D6AvubEJWvvJZEEOXs53d7POcnCtyoIlCDeeSZXE0ha3wrEmRPWVS2YHfSN+yI
ziFxU5GMFhAFntXni3OmBSkEw9QSUcnO3wKG070fD+4FhXVAt84/g4bGGldYIoj37SKSuTIFD+0M
VdOWT+ErfownxxvWU54DF23EA2je6EiMRtXY9dtYYe45ZYoJ0Hk78WvUeengNmM3nggXdd+2FKET
jL98UW9pyyoYHEaXXwTpv10Ma8soMJyZjbcx+uO12ZHBg3+CPhyy27VntDhIec86OFwVVrOEav8C
fhgPLcW4dDaTegZkdgxhRsvUg+5F3JaQhq5CxqcVa0GBWrfB4mrfAer4dH3wlLaIT4syLOWekbcT
ThRmYHizdaEolRhYcFGzKtVIz9xbSSuJEf+yK+/KKbzYhEqQAxeYWqSjGB793tgJYfqxWoCHvKJu
ggONok6ztus740fPu/Y/01eozsCOhF+hfw0It40mgvMwiEefsEM+i5E8xQ2HtoZcaMlEyglAIbZr
X2w4N8OoOM8RTndViBpXQPxPgQF4Cd/2yJNsbLsPyHmJqSPxCb6x4L+Iu14jcqvb6phpTEz4HoqC
KRXkqG+uFOb/4WkktUVUpbGycj0sx0FvSeD3KMrZgslaiHEej9ELXiiDFVXRj5MZXZCxULvH8IBx
kwYc+ayLQCWIm0X/Mn5d1iVCgQ5/Qw6S1wzrbLUQWHA7ceh8w7qcNnGNDr4WKgiRA7lpZ361f9QA
ulzJrFkEHgUhFUpigJhTROnFfpGQ6fJN/FfulGNq+91yaUL+dR4BzfQJ9WEbNtOLu+e0k885tY/i
NzeKquTcbKjD4yyZq9tCWnx5zg2SmDCjCb/HRCzXpYkRf+JhFvJmZAq0ggXuKOJK/zo4ZjH8F7Id
FLPmCV5e2eodrgdWOyNoGYwwRPevEdQk9ZP2ehUTStMStZF8TYqgRd1Jb2rrmvK51UR71b0nISi8
aMnWclYeXtNoyYjG+/X1yv1BvTp9BAK8Gv+8roVxt36SFfRo5H98wK4zlP+xJgbwAT/TWuzHMTAt
dWCqw2ybLSxS2VsTBvrAVEicsNmCffP1SyD2WRueFPmYOKD4Ge8cWcgVAB3Lw5IcVQuCLYkvlldG
fXCFA5zJCLLKZtKRvVEcioqf3mT7Q24D1XQ7li+wIX5w3rrbytNX2wE9dli4lm0nuR+Nps4J1CM8
z2KP1R9Oi76vyAyEv2FJQ9l9P1cxYUQCBmvk2jyzdRnDhU+bkabW0a2XbMxWichKQ+9so7X4r9NO
Z5plQUZvl0Gj8Fz9+s33IHBU9ysULwD/XRPtjnbwrPa78XzftJ1+mxcbBhZKpwrMux24Zj1x2S3r
Hczh2O4IW8pfyWmZRFrQBd2S1in/i4qiH9JVj/Z7mqbRQAz/nkJkLQcuA783PN9CWBkYd7DaGGPp
EF0u9jQqwLQYbaPe/nOW1YT7ygwmjcYJeL3UTAeEbg1Dr6NQgM41MFvLCde4qmRqsKowr8pAhbrg
zLc6wlzp9A6w3K7zXwTjEwhnGIf1dot24AY++enIpHpeR3h3VWSpvW8daKboKNzhvYIcnhARVi1m
QymVCcnINioLZDfv7+0AkxY3xwbY7CSo6foyBqfK5kgqiDjvAJQcbEOejkEm6LraT5/aL6NRJxZR
dUdTGGhOnyLeRHlWhj5KMcqNwe2HDnu3AHLQVCwF2e7x6BpOzVp+xdnCktzJwAau7gpJDfXs0TQU
smqyvRxtSNovtjsc3bWXGYc/eFXGpuLLGIxrxNnH8IhMiklSNUXiyieSY7U/OrmL1UPlu4a6Zkjs
7RK/h9B3zrbQGG3YNbObSVMt9hukBmGVdBE2HYrclSa/+0SUEYzI6uEgZKIvGAnQIFYrdpoKxq7n
AzzUyj/iF//jxa7LnVesXhquXEikUSJeW6TSuxczSZqIJM2QQ50zvQGf45Yq7ObOVuCxp86R4ejP
1BM+zNCCacvTHbALow1EukPLxlBLtBrSAOWtHnXrKmMb+rF0VNHOBdvQ4r75Xv6U7IlmbbGWkrLN
h0aeTsRwcyN1OS9VcfteKH8rtocdNnOgMdyDfDehzf3Mofzgl3fUE2IOHYt6UkSwWhBuIeW84f1S
uZttFKk6M+lMJaSQ9XGbwI8HGWtnMX8kENy0XypgkJ1IUHmjMVa/8vEMULvfGGoGcHBXDoduDrMZ
MwqbQv0WiwgEsmqi8tt04prAnvasYrEWftbOjSN2u0qqK7eIRBKDt7dYzIki7TTmGMh6zSrRe6xl
fog+EW59b5Wgf0VSGgwgrFXCsi5gI9DO81YB0jLttY8Yy+SwxYdHoJA/2m1PDyAl2o8NJ6buTFOA
Ittulb6l6Ec6vYBr9zHnZaET96i2oRT2rkXK33fRK5yAx/zQ+ySS3RzOIz48DFHEPXZ6jCExQ2xJ
PllkLVC3y9krNDZJw/ZIAnx3a+KZ/Jl0AHyshJBvkEaBFAZzfJD4bCC50AHWDBmVuOF/GvanVWw0
SU5nuoNN0J0AQQcbuMc8NjUiTcAAfhnEY95oBP3p1sIBtoFFCFwQ3jhAnppJgs7AtgTkn+wijhy8
kDrDvk1y7xmc1OdHiXMcPh0WeymXTbR4TqEjA6zv32Y5jK+EY2lMLwAuF+vbQo/+vKAG7ua0po/R
LsFN/gNY37RWfNmdk8XJaQKcebIDEsWaLAwEncqtMWOR1QDASUw1zYLtpq7cGnI8DBNSkwASmMoY
UTE3iweWD9ASIMEISdzJOTirxe3i0tDci0iup+MjHIzYN4IGzOOa+2E+fyiM1cekE/W1H+hcaH06
kmjdem7Ajra9goeaAqdzPFs9BBmYbcXcEyqGFmHkU4MfzxGiqaCXIpSFQppMX+A7Kyt3qYBiHmys
9exzfbDMAn8CfIa2zDBS9syTlOe72aI8mlrSko7y2FGVo501vygcfDsm+Zzo3UTJdQ2MRj2NsAnn
4mhv1BhmHT3wdNcklnObf4wsAyGihy9YiHY26Vv88KyX2JK+MgcyyFlsR91KcBKRFeki/PgUufpG
PW+bjn6SjEtT5nkbDqGc2YqfDzqDtm7OshHJRbUHHkh8zXFEjV4hPdWeaK4JeeHNOMPo/6PpHYUA
ajNnt9Hv1E0WunA3aJ3UKFixPAaY7VaO4t1H5aAgXZqXyE6EOayTUnryaFie3EpQUFL21ersLsV6
hnb4p2MXyK+RV2bIQhsiI0IE491UBaiFOTUpz/6GB8nqMy8jwqVt77ArCY0viOyVqLmnjkF8WH4s
IK2UEq3jm4ukrwL3emM/nyCh196BRxU1GtMuCPDw+Xp6BLzojKc+7hIpAS3PMZlz5OvCQ/exvn0e
73VHd/ch1FnDoS06gU9EjggfuVDDg5OwotGgw8K4Dbvx4wawelHF4Pyr3dimUQYCCfbsC16HVxve
klzd1OZdOwzrhq626pO6zf+qylkBAjUQwJCw0mWbEocOScfV0a2vT9ENmaAElrM2oVXPcXmKy/A4
jtZv9MJI3Fj07eC6ZezNhG30XSpsmdaIkqfCmrHk+X3bgLKOYI1WL3Ch7SiPrgjNgEJ6unTdE6RT
aykA5+PHFuLk8RX3pgeICnOlKEF1rHkWu2HqGRIoJc+l0qLnWqsHfOE8poDWlbHu
`protect end_protected

