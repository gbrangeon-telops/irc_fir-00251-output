

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Gub1VXq/9my70IMNYnI+loF5VZ7ee86ZBpAGzL5j+jwLQfPXAWQ9vuaGimuQWfCvI177d9QCmrcK
lRbHtdPXqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XCHJyRkscuJOpjxAlpPvd15b2tV4+cleGX5HVVJ/2Y6XWbVNSZsCQSUsTkLA7IyKge516I1wj3zW
vSbDpitOXWUELSO5CG6d5r8ZVemvSn2BJybpLquf/4fVeS1c+edRHNf6tkj5Q4P0LsQat4mBIGGY
5hCeyo5aPtqLWGIyMEw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RqwoFbaHoCNWZ4v1HvZQji+hXgCjT1Fmm8RnwPGBKk3/N74/TfbSFLeQsQ92UsPWvT9gifFKCg1j
7eGei0ot9ncWAfgeoFsw2zoynofNtXpuT/2o69ZZvCyc9OMmSHilEDslciAlUOrRZtsCwGDHNVP2
rJ/b+v8vvCejKLtIXh5C95/DXV+eEcsjEVRpSeKGeZ1MtzbV+fZPJnRzoH2U025UhnP55OgE68T/
nVfgRgkiVFm7ZUA/Q4uTOx27LPbQmDFQ6plepnrYm3dIFbr3WOiv7AWG29Y9MZiC/1j4MvPp1qqq
xE8dCNkJmOz9uD4DUQoSIb5VP26bf6BmGLvFDw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uV7zzv9Zx+u216Ml06an9UEqL4ajf0AMjc1K2s6n9qbyEnUVTSm6yFZ0M/IFYGglaG6jdDDlz4rd
W4zdLmcu66F6EUQtwXBmHtk4+/Am3fKB3kIu6GlcyUoJhx3DF0omCc81HS8JxypUZEAxz3C538KP
dZmq/6pOZleIRCziFs8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c2sM3Lkice55qsGCUzeim6Qm2yWa4rXMhx0Gil9+l1mRl06adQHebvNeaVnD5l4UfTgDiNRnixMg
t4I3MixM5k+/dqMphg9yh9uQH4HJHJ6CTIPJ7b0uq0QUv2e+GjaxWZa47ZVWMUHJwpscHTsz0hs5
a4sgfCiRr4cQxV9i8u9cWFqcZ4eu+RYLEbH+mYK06INaK4Fg1vBkwveCaGhKFtvHtOBXP2o42BPE
2i+HCKN5sLyGLlDI9h2MogiDBJsNAtjJ9geF4nPG0e4nijR/pyFXErJCeKppN9041em95AkpK0CN
GYWuH0jkznlTfi9EHnlKl7cj5ibz763zI0uZLA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10784)
`protect data_block
qtrktBBjXo9WcUivlxWLssPnooT+/77/bfCaGPVcAvDqm3nzx4naKUHBEMZmkAJFmvedijIGR4TT
KXID2NC/7yjp0JZeoUHJLdpRETWbaRTjwuL8Op6P/+dbWpDEgdfxufs2sGT3fqgLAg3zrf44NZA1
D1Snf4b0zmERZHNFA/21+A2h2QSajCaMChKZR+fJu4mmfYRwE+KbL4GCTks2rVb2TcqNVZl25c1y
a+R0WFStg3nPJxtbtIxJ50VIoNtAdtUvJU16qdfuKn+6uY7VZgwIHdeBk9+9TaeN6DlXlooY5QLG
6QO7LrbF1jelbT2NFGex3+KGCzZBXE1rzmrqbLkmOMlplt4kS+9Iq4npcCMFNdnf+UjEcQF61bBi
uJWp42x0qSEHtZGVLC0NpheHBuVXulbUp0KE99gR8gWISNk30acUNSUfI9mYYfvvgPTjJx5MFVcS
I3dWSqsrAK0qUTFxTLepl0JdEE8ZpyYVMi5iFNaeG/rQVglVPksIgENndB3CzwIrL9fbrz8m6UlO
V4sDZzBo97rTWH2NGi2iPDbhcMg084+nnDmOIoQWl33zzahcpuFZHdtjb8sr2+Fp0HMsy+w/uX/R
8ivFgN5xNTl4DkBUkyHf+Kd1DDGLC5xfEMg4QvudTLQHETMUL2QlWuATsNJMZ0Kqttn1IoUx4XtS
5T1//GuGQI42XfvdXR4AgpzWN+fCkq7wt3Fsf+lHklkdnIJ4ZUira1fvHsy0G7kV7b2LavXHmYCY
13xZcpuA2EAlpTRI9pz/AYjWJeKUSOCUTpvWSVHKTd3dEA85VhdfSCxGJDHGFDIb24L9tabcnkuF
GRZPvkYet95Ph9FAUtiudv7UHeHhlIDr4ENuOv5U+OVIWSwpmjQxsU4dDaKMhfO/qPtgNtEghrAZ
Mm2mMZfn8JkZV+RSAfAs6m8hhyO+PlL5X0iEajJIiMkPM8cs+dXqZwJ8i/pZtOLRU97578uDLoxc
OzhJjpcpA2uqpJ+o34Bwo/LgnOyPvThva/MnsQ+W5+/g0WdL9KvgyslsldyOpfME5Q9Z4FpH8Qli
auzMcYcDRazbahT4XngzoRcoq5tylUVq9noUWl9+7O6VyKS/pzD3GWoFLideKpE1SECwRNYUkH2e
G36wCHJXl2Ntens0aLkk0qsu+Q9hBUt7dbBUh2Od2bxpPcckgQb4ES3mIWXgcOiSKvK9aAQtNDsd
7PdyCHcCoSJVQkLwc2lawoTyPwJyJZs9UAHFnQYt6xSAaCXqBL/PAxgvuEbVQ1Co1j1hdQnzbYgU
PpblxDhmkDYcM9EFbDJxEFNptsg+h2XnCqjpnVo/4OPGOZ6yeEeh4a4xeDwWB/+ez9Z2x2zkZh2S
uq3wTKrrhBltadspS1V0nyMIM6ecZU51hjNadgUdlxQ0DF7KDfRYoTtcDKXwDHp97xfqLvhVNIVY
bgpHLNwkv84awOBxJtRhmDEHddC2TRD0Zv1BTw/mobE7id9zMftlfvmPaWRbsZnhSIMsiR6hxf4q
/+xheZr7xSlb1khJAVxb25m18JD4sbAH+qr+oVKWVKFNV3r4djxbAROfWQDZK6XzxXM5DO+MHi4h
giuIihBCZpiprjVKOORsEa2QG4GjRBBKt7l7hQLqj/+Jbs1AqEbZu9hZ410rREe1KgemUyrrRcu7
7pwmkRRMexKWEX10i+zu5U8eVRnjWPt0Y2DUr0Jx83IzcehCwcty45ZYIAM3WbARoOgmP8uCwj9n
4jXdhguCgn7y+mDXdBsne2V27wpWkySnoc6RNnfVdbi3P5boJPZecoZ7vjhFdUoTjCmjnTk9vCo9
Hcq2iIhYNJ+kmSMV4myblifWboRSOXXCOhlck9C8QCtTWwBR+QrbbdUufeaP4kZrq7HyE8Q8Zltl
ZpM/Ip7Gf2E3Ghv3kyPz1wc3+S1FQwL3xpxxHbam5UespQQR//w+JbavBGNXJ8KcZhCFbNwzFKWe
GWTO1YAx4sIYBCmbujAc4EOsuIgZJI+Tw56km+yps+hRehf42lbmhayFIbZLMSKHgb3P877cZZDY
C/wpizrYeKXaff0x4nraeHfrg5n1QohMUv4e3PVa2qIdKotdZB7HoL+wY6skG6QpZJnOuv6TwnLd
n8H88RvdlOzYy7WBs3dcJq0KnyWIHnmIFIcBEbPdS0XGSpwAM6HQT16QH57a6+btLTddDDtvuEFT
ZQbhKE8Bx+kaMDhacHt3wue2+SrcaAeyAQHTOU8L3r9OtM/prn0z5W4aokyb5R56cBI1BLIQyBzv
SQoMRBeSAnsejXBkswEdv7eJASoS9HHqt6doYuKl1uzyGQX8wY+/OYjbQGupDBp81a31AtDo6m70
gpZb+uveOfsqpeKyLnt6y4M4QOcyykMa3uAXgof4pLmphKz718LNq5CEeAj0Emdudokk42VzoA0i
TPdYbLvqUgpTxwWPum9XM5XMU1u012aFKr5Vef8iTXJILXLY97YFalO3xAaO3fLYqmV9XWc+w0Nu
nnnTRv+Agw9LjzPUhyd5UJuqHK6mt0TyZ3bqBHgir6wZciXgJ/dN5Ep5H508MkMiAanpk3a1tIVe
ihTrKIUGw97Prg1W8syv1pAYCINmAEWrqp/iPNifhhjebVrmTJBj/XOdDlP6HRy48BnY8WBwFXFu
2nnQHq/nWVr5tKgxCgdn6ilVtWAU3aCcXEwW7V3nl6dL7AxUlvSykYsARr9Ym9I02W7izURLQr1l
KYqXVSkToIzcshvX9sid1tj/4El/8sdrT1BtalOIJM7kIHLxaheqlogx5tZWUKemY1kVFvHkM+rN
jmXExnF+K2LsnFNV0SNmiRHueeS425Qq4NDtyUJkQyFOEGCGJqbtvtgEuXwY+iFxDzNE4Vfh6mTN
28CXc64Usf5p4HZAAN1EblmgLJkYKSMWY0P/oLh41utjYt+jBW7aX4CyLEzRDYA0CSZz7gS2zwTP
9IdDasqjPnRe+/jySiOT2o0z+5RTkLKlxrAqr5H8p8iUZ+rHK8dZz/Pez+Cnf1CHbQdba2GGcUUZ
q6Fozyw8nN8EyVYCvSU+qZqfkfjgDcjkll8ZruJ3pIPGoRADK5bga6tnaCgkmhBZsHEHCNTxzUv1
OoFg/N5BmYf53oYPcJc8197OEJEPLGbOihy+ZifJTqTKufMakabW3X/xCc+QIVM2Lbq5NOAve2wE
WmD8h8o/smqdvKei02oEMjAWA51IzkzjhVm5Z8MGvfLSmPGORv/t9hh/79PfT8Snb+IrzeCBS4hE
JhyVtAPWV0ZsSSb50lgRbymJSKJQjZ5V/TqHhZTJ4NGgPrAdfZJbOjpuS8lzf/TDtI47cEQbLEFp
leYc3GNr5s022rtiC7Hm7nPztA9DbYfah1pFSVoo8Uor+g16MIrulVBmgHaYSoc/QmQQ90KxpVv2
J+68E0zqh5PQqCMC0Ak9KadGZ2gS57xaBYQOY2hlLgiZh3AqVPsvg3ArZRKUHK6dwawXoZVZGtei
+KocIni32cJsB/J5N0i/UfB4JnHiTAYADm4zpc3o+CUv1m/46BUkS9ftCi99jHAIOoqeklpUqTtH
nOwzEaWaYccyHjO+OjsRrAjhhFBZsVdA667U1mNaLwJq9kby2LeS/OZ/KKlGWU8Ec1T6Ml7+/BDV
HoAkBWz1vQai0zsEjPZeYlF8s3qpuesgx8/1iuOY09eMn7O4qyQmTfv6kZhcl/+mhdVyxreCrSTk
H8ft2ymTr00IS2VIxhSQXHEKYxfZYD3Js4BYCGmxMzsvyFXs6JN/dcBbRpiyV27zEHAxhktk+p6V
n1Jyna61ryU5PuTSUy6QOVUKg6jVlWeYcHdtjylRMS3YyH7NBpzXNCdU1EjCWpnFXKoApRpU+9rP
3z/EWhS46dr4g2TkVJUd+1lUdZsLAqJtFMaf5l++Bwhi3UgOqCR9pqxcWJuaohh7xpeK5oBe67Dn
H3m4HAIW+GPVZzJ9vXXqxd2WqXm8EnaTLkJewqnm5azjUg3xBof0yWzWrVDgcKs1mj35cNxXEjhw
FezmBjFxqT18HCGAgSDSuHuhza+2K9AWZkqFZ8/Guo7NOFpWIsR4+ElMO7/Tc2pFgqTNNHpv3Hx2
K2UpfdBHEs8UT1sFIUOnMCe1GYdo/w43PIygnT28MWPSdudeBng9WwE9DImswaQWtr0pEFxIN/nn
ceGjGfggV+M7xhqUYHCvf6Wi0ZtOxExhZw5WGgpJmOJJHPvihi9Jt4OUAOOWQFM63MMvxpiTFkHC
2PUFh22eg4WlY37VYxvnN1v9c2QdKkp9Rp9iaHFOT+XuJsP8unpkbCyD+ZVz9gH7Gv7Da0c81BHg
gBeB0y70nfIXeaqIYWIrPXxAvN68xAP9npQU6myJfM7+SA5kYuFVoYRACBafmBUMWzxCVXSP0iAs
Y2k+Fe8WBNjOrl+zRABUQybJY2uN2QQHCc6ahrfFBmSYkeoXFz+QNPOp4qoX93sK0TPha8F3u8oj
0ZaZ7RYs1FMy55DhqZkXuLdEtJ5Ix0QCOFLC+Vn1zSmqEzGxxAQh5D2kaaEpC2L0fhs55+52Pftw
88oHekUnbGZOAJkNgM/ZSO5rj3XCiNnpheZgMuEOXy8X/IvzXX//sYF116qKrLgSQB+h5SkEy7pU
Y3huCtLCOUOD4zKSsq78UEPg7iGGwZvSruUVMV/lodmdy4U04nCmlOzGCfdijMzUa6gxF1MrYXFY
2YfVQCnpmovVDhRe5euROn049NUj6l5HFCTc+VnRW9UXRrIYxAHoayKNuL6iBxV8kUUId8rgBRhg
4jXIePgQKRZi/mcrnPYyvFp0tuyu+l7QOunGvcwnlCK2sgqXmnA67iBcgsfvYT5rU8OODbiJcncW
3a3L7C7kwN3v00zfrmBJg8hY7qlQWZlXpkDcpzHfL5mSxcplmzGUEt3lQ/KPPpdyRaT2gB79NK4o
9YDjia3zEvQ+R6Tt/PJ/RNNvETxl6hoPlS/vLL3WkDET+WCW+5KckvifXFI6SnE0H0gRjZ30CBtx
Wa2Ctbk9ycqFVGpF3qvN3EAXn7HCJMrl5L3lc0o1JAZx+7cRWogy9kpwBtQd475cRuUgyZyycil2
SxJ7HaNg3cbtXNQ7Fq3CFeajKLMNWDxEIAVmFEIRPFH0DdO/8sV6pZxewfNUTGNFQCL8Oq4zdX6G
l+/M0W3QTiJUlJAhCCr5QDPKieGQeFwDBG5lnpbkGfJ5hM94KDXpzdBNEdwNkLr57YQb33BAsosr
n8jk4DkXFcJip1J4Psw3KTrZwXjHAxQJj5zIwUzgN7q+kM24LvI02pcAKSKIEy98RMaMCdGzeqzS
+/DSfTG+zEILPDz/0JHJRIjzS+LRvzzHrheu4thFRW7TKhhwwzM4n7Y9SgS8TCuUEF6Y45W1jw7h
eq0VgGlD+UShM8c5r/kwvUIyKaFqqLEDKjSjC/Ahjbipgoqm4hNxYkq/K9GydODxNL/kLGRZMO7w
/8Le6FKw6M0FJjIkjmDFXt2ma4OdjqfynDi8x1WCOBvm0+cm+ys8+WDkN+HhB1vBmgX2vFzf6zlP
8Qbtr6VTYwPzRxYDohFL9l4twW8gEjpI9DPtG17SOFIVzu9OwCkM3UCMRi23MFRIwvCTZwdIOAie
lFJM5ZxMrn+oF2+gdVX5QionTMZwoxMbuHgMU2EXBnAvXJPsggtsNAClakhBXRy+dbOIaymcCy7X
G6kGNjnfk0g09+/ET/z0dn7JjN3YXr9WRpFIYNMN8x4NnA3NUJucc3x1QAB7DiONQelCtlJYH+ti
VmFcHngu1CzE/IZ+iMfpzTjsD4Af0vMZhszGofTAxCuAHkc2zATpkUcmkT30W0YImOECblHaTL3D
lVIaPvjCeJj3Qfr9QSPciG60qNKjK+yJPzSZ8cBfBNOCnMvmGj88pxS/5dKhJIM7FE6J1Y/N5MsY
p7k7YWO53mb2bRcSvKtAIDwMkrFDIKzflr39DvyQOoPq7cdxpbdO+helzw9/7z0GN23tjgd1EKBz
zD0qI7fYIdd+ul3JmsMSEpzUuRekYU+PDRTvylZ7NVnInLIE8BcDQGt9EBSu+06SeE7jfpLD/6Q2
hJ34yDkJsu/bNTIQ26vhzF6+eAYJaGA9eRptgsKpEuUTScP6RII371mWrJ+iS7jX/rxZ0bCFsrZH
NLSHUdQ/KV3YQpzJf2X+VOUnLV70kwl/OtzFQc8Wl+RsxppwBMbUsYsh46naKkU7iCJCkphaAGeW
MtgBdERs5IDboOmYT+BWVJ8RjMBAEhXS2vsXfpP0Wb/SkhWWpHmkqZH9zNZX2yALTYedJOneZV9s
y2BxkdAL+coNuWBHJHJUOlNoZpYweQXSHt8K49/B9n5m10+mOQ9Y2eammHsPPnloD/oEDj7zLoAx
dHmWU0OBRKGBIfw59G3CCHZFee++pPU7BLLjVcEVxkiz56aNBpI0Ra50ztKyRKHWzSY38zO8l35/
kBcf0QQI6s+cHs891tBwKSYFBqmIlOV/b9izFZf9peT5N+FdNX/p2oEAfrH9L1UyiMDANKH+jRRn
KBeuUEXa7JUflnYM2Yi6TaXpSG7rxWK8HTX7Nxp0X3W6m1TudRr4RuVTYjtXWRAMrWgBhDt5qXxU
+It6SKUAtmCrcG1vDgy/aa5nbPAhV2K/0LpIinXC8hrasT1vMpQ+bwwm224lF7axNJ9vM4NwcZ18
ttKuiKq0NIHdBD/fKGQLJVThT+Mm4qdih1DIS/8LK5U/s6LnTIznwyTqtYztQ7cfJl63anXy6Gup
Szf1wwWtsImQT04n7BBFNEqbUU/mjZpHSyT44PGpoBPsh+8G8DlediGJVN6pWOUnp+Rz1q2SplL3
20EiaX9RSjxC3i694Is6/E1pqi2ofhmPFK/HfkVZkuNUsU/W+aaseGqDXGd5CqOJ7FwGja1moOhh
KlxVTPJlMtF8ltlxxKDj5hd3OoQ6nJ5CCuQvfk2fVldt0gnUN9cMSxOSFZPSnRpj3fFz9bAZctkV
gL6f0vMFVVT5aincmIm2VMzAa6a2UncXqk6ycC5k9vRp3ehChKR4/C5xqS+mFfnRDDxciSCRjlgq
1CI6cF5DHk0hP5EEccLW9gaU7wjSNwreEH/CwXQbsJ12Xc2jidUNMtCbe7TVpR8ycPouFF+rI+3+
geCxlrA5wiUwFg1UaRvZAxqjjbT0n+LcwOPbuYJu+HlJKhZUkLT+n7LGdtFQbkSoreAP7K88J00e
EZ68k7BG7yVaXhFKIAR1n2jjcU3DNfqFUZRqCboI1WDHMe2YKiykRa6+oOwKo1lzbY5dt+aexA3+
HQV+SwYGTdOnk95fB1tp/MSeQFcdeA5Ij5ZrW2XWCraWQISD0+zyat9tYnn7H8VHeV66PzNYwUjD
mVYljEp/jlA0ywhKxSCn02fJtOjfzk+RAbDWZR3kAt3htr3pUK5H4xrRNZS622j3H5qitAEDOi27
hGprWe38lvSRC8XMEEpp609lwnumJTGzl9nPUGhA8+uDbJdTFtC7J6XMHhCIqgxScsdwHeu8GNCy
iX7muH/fjFf/68b3flw5WaxIznJx68qdL6uhYoMQRhPkGkMjkwPNjRgNiAHUgpIVQfPqRE2DvBCX
YZJ1S4nipl6oa+eG+LD7Z4dBfyFO27NNis1EhAO3wuvXiRT1gZ06OS0/wl8vNRitnPzWm1bZsX6V
HO2CdSC2w9xNcboME2ecS0Jm++UCR+KpH+Jsc4VMJEruc+SfhkuJhbOLy0fghWTLKx7+qIDvky0s
x+cscmcShvlMdHQH/S09xr2emlPkC260J2XJYeq5s4nneCBbrOYYvS8eBuNeSPYkEF+jxJv891PM
euidYS8EBjgGlvSPA6B3biuCTsdmPAS+jIqlNI8uwPWhVHUR9iD9p7eF0PWJnV24qZZCPYprog5j
IMS1xXmyuApppOd0MeMRiUMyd2i40IemvACuRpC+oO9xtQkAYST03S3ua26e+qlsN+3a1myrM9Ea
PWDn4hkdPoLF10i93vPBnHqprkH2ZF1+eL04n2WuyLQaGeLsj199FYddl7/UHI2YmVknLdEQ27R2
kMTMeJSxKSgzGWPxtFRu5z/wHd4pqi5Mfq0nwoEcF5lqpBROslRa3KF+joeicWfr2kjC0Df7VPQf
/qTY9PF+bl4rIjWTETIBhKKHm/byik24op3+knSywrishxpDpiGKiakWmrgsfSRrDXYSIBRZVwLA
+e+ORm9bj8HNLz1gtc3lzgCQlnjLUtJ51cadnlts8REKEs9HVeAA5bx6gtX82Bnv1FPq3jojluLh
eWMbzDKwb1dDuEo3K50+8c2v02LDckMgjwJ0ZPbgv9SFrXJX3D+FAQ/u+jbgMwSIPLAJCoU4Xu/T
0jqErk7NwniRfByZTAkTBwwY0YKoG5X3Bs2YwSRbFec+mRIEebfvsR+cQuIgn+LU1I2qJVDcx7xw
y2GHy06MD/WHNgZMqBE+0HHMpPcR2TJKRU7fL4kSXBpA7kzvvLZX1a4WzNiL4ASkuGWnAo/zq74o
zujEBcaM/vaGBP9oWqMXJkat3U2wDURwk/g531HbTmMPzJykCKaeykXlDIFaOtV1VRJpXI7V2VTv
sRMRcIIUhn5md3o1PmXkQwpgYKfMVpOa8Cx9Jurl9hrrv6fiDfwVMHPTZGH4CB45+XF4/lVqV97n
wXaXjdptiQlzHaBHwrxONZfbp63bdArHE77rtDuw6LJHzT7LNG8BBfd1dFqOtTYUWq0WKi17s/xr
G5VcyA1RlrSTLr4+TlRFRvV5ZRc+0F3/ecLHAhvtTvriUMknh//DIhoc4E2NAw0xBSKl/kXPIqKj
rLPDyzJNg1DouXl/Y1cDUIQpexuPnZleaR56jfO+e8pyIMHXRZLkSk+0cg5bFWGS8B+MMxyRwiKb
7xfg36tkDL9TnqOKYWzAw3eeIfCe+n6UCJ7OZUwyORccN0Zqi9d2+BOQm1r8VoJNf68q6o/G/7e2
TGfDbDQk9JM1pXMn0I4sFQaRhnfTlWL7MsssoMBp3nsD6r+wDKJF854TmBygtFSsjUZHsNdEsfT8
5BzjEDbaeUOVPTz4cFUGzCTa3DhShv5pZO+CsDdp4+wYVlOeDDhNI1d5gm2MNSxXmi0c2YJX6phE
vkLpW46PvcmSIj0Eo5ktNFzV8mHXhZNQPcX1E2BjrXJ4ieFzAY4Dc057l3JB+S71zYenBLoZkSCj
eUuZ+wgnaQ9RRCfBhkn27WB366X9D2aoReuPEV7fF1LIjMVt9FzeZ5nuUk3EmAcxrusF8NWLGpBG
b0hiTpK9AL+JVR9p9gCUJVTmVczdMl74DG6++F57WyN2oV5PR8+RKn1ArCgbjamZbyj+RXDjXu6i
qvtbyU6UnWmyS+H7ha1A7rBYpywYqT0Da54jKDG8/GXwz5FOIVc8gdXQ1XPR/kXUtKXTdlba+6y0
GwGtkXD1CTDo1YBroaP9ltiOF6DwodfooPEH9Duxp3bNul/aWOmrTRwlt4qx2WZQf0TqZP+iB/3b
XB5vPX/IJvJN8ERQM0CaFAHCnMUbbAB8GwlttZGBT4gFVm8YKtjs6vDIeZkYzxUTSeaYuqk3VpUg
Vzi+6dPA/6hrUbWQ9oetX30v6wGNEAOhF/jgF3BaiGyvm2mIitQTzpkfRLkkkzXvwSjOo/StsK8q
nz6KzY/vxmiHWDm18EIGyCbTI0uUYsA4AmYmePIrvKMWaFMkSedlvZU2yhktyhRdJkoGSrbO0JQ7
IX1D1yR82vGOOWx817mZ/F2ZH8QfiYoNHpf+ckhrWpz468IE8mvsjjVF2NNA2FHUvTX2qJP1H2wI
ZY6kZ08xSJ7PfO282PElHbOc+g4qL0XrPXOTynI2TzRCv+WuRntAI7vgY2gZ0vRHTwgrd4nfHxQZ
7UOZBAhsoS2P41iekpJYmLRVmfG2fOKw0cCuJO1sp4lD1yvpHXhO4P4npm7fNSyNsHqqPB1hLe+a
SEALyDD8IhgS6Ck+J+xhHjPk8Mhv5CfFtm7abCL7k2CPCALOOaKjgxpFLMyQ356Uda1UBwthORmh
ChS6+DB+k8pdvAW7+V8IU+RuU1L+rRLBNqcT7dPiLeHx6riWY0MAladZI/OijMlu9BWeqqkJDVYd
yiRScNzskhvvRvRRzzgwV5cew5lFrlU2zMrZAIAaFAiUEm0HUkVGXUB+HfMcKEDS3oqml0CEbyyZ
ThZRA0Ljhk2HKk61XopczAlJ3p5RWiYBwMFAgPtxBuL7MEM1IS5PI04Hs+wmrvddsaka4FFZDmRn
G05vUywQ0ozQVWd0XijLt0J8ulBs5TwZCEk6TpuuUItNbHTZViQgiC7vm2N1yEdheZ28YT7D3BqU
mxZZh/oNzKg/H2b7XW/ZhTfNOJnrcsKPv2hCofuJP6jhekq8eeueTuqY0N4uVlENxhj6m6ZFmXMF
gFbIf7GxciqSUap0g6TikPeBQyv/eB9FXYWe9cJsTtYrKeeifjyfdlRfGIJT3oNKuJ6wUQ0ujl9u
Cgqvf8VLvyfeHZ20Dlp+ybJcZOFa6/qFHwkc1XC7TFle7TPNn3rhsmH/6VExjX0H6TsHSyFanWGt
qBX+88Np66RR8jGBkORL3jhJAK/TDYqp8ZCKQwtdGOSyalYdxfhABvNOy6pawTy+9VzgIY6htMsr
PXtnvPCrJDUKeDRqAO/RyN+Uhf/V9EKfwjVvhSNcY6Oifd7A069fT0pXwxNJgVf63ykM433ZKg2b
3+WO6tDL+i1WbMeScDtXVN7CN37voT+XeZTDx/4WroFt4NCWaI0C/pq3oYp8pdddUktsM2KEkjGe
UE4tQniYDcKb1OU3x55V6bycTu8B1gpphHrP4dccfpV1878shBgG2IzUOzcqFJ46//nequtvObRU
SzIqsO/nFNmh8lRjPjtuPp8uLE7pwgevHZuPRfh/T+iZ92JJPLP6GwhhMB9VAgfBSglIOztqNANk
Qoyol62ey8Pbri5p/mYok7gTpzgmBIPPX230DF+zbbtN1EfefHhUg6jcwVGIDGIcHYWJYOUpWKdb
KKGN9Lny0tOjVF+EsnFRJ2CteiyNIiJAvGlnucrzH2YAsjGfF6EJME+mPJ5WJ0vGP95w0qbUNRnE
voSWnMbqVeiTMkU0R1h9z4uVLExcijN65wkoo3RR3g977behs3BZy1e8jBXNYjLob/TxHOUFEDao
DbccsM+yFW0DC1CcgarjZwTdVL5VeCkFxbcOYSeFsh+0dadQZfS2uKbzOEshn0q1b8wSsoGgEFcI
0IQ/XKNTe22ex2L/Qv9q+1fKJIQbkuh6PoBfAa3i1/C4m0DiODrhrqSgdnBnP6PZR+X4q/nY5bDH
BOjk3MX0sog6r9Xf/XO7CNI6Q+1tYw81UfU+U9Ab3aL61HgSCTQCscC7BkTyot9RDNHbuy23T7Dj
OiWRm+dItudmF8ggxqTVxSklRcjWhYoERu/c1fnysBfJ7MWRODaaP5hJkolgU2gbNCTE1b/U/BJI
votu0GzHCP6tVrB2Cwn/CKXsZin0xsXtp66Qygiqs+zhVQ/80bJnl1VbVA3mE3LT9KR9O7JkKatb
oN/Bof0oJaEH3ZVlESikFqRIIGvrld2gY68VhePc4DkmEvyB9kbMN2Yo2YSsbi9Sy3GShOCIsmhp
qIylcHSrXsOgEg+rQHzI3chEpoDO4HIbaGI6THh1v9F4MIgtNT9kxWP/mx7HPUzlHNtlv7Qik5Kv
bQP3ZPo16Sr7Km9GsSlgICunB5H271w014qg/mduV/pVS/vT1oEsm/oCHM7M85m6eXAeOfNOLeze
pFX8xFJFMUtaIfbH/nys/cscSs3kE+3D3QrnPTSNVmf1XjKQg5P4rPx1HYLylJ9/sKtAqQjkMs2I
GdKvlUv6X4YYh9/bESDELiyBhTYpv7fWA3MNdZEnviSy8AByfwHOHBfsJgLV/0SZdEbimOlKIX4I
bQnuio8E5cu5R5ZJ63ZIDL6m3D6HMfpWtmdDqI6riivIejgdyNLfjq9qdiiSSSo0nR8YgsHxePdX
9vOxy5eB4cadynlnKAXVfr6RxknfxvbOGHeJTpxCvDwC2KuRL/XYPiiNMc57m6b36hlqyqzxvNKs
AHSm0dcFvwcaa/19rEuhtLN3zy4brpFRs3IE24sV/EHov/vj3Eyvh/4E3FOEieu3P9CUZYVhXIR5
XG0GS67ju60RC8UNsJtoeaR3eSeQ1yHxx3wjy0h9sGHuV2p3q0d5691L1g2x6lllK7EGighzn27T
8FUUbscL6QasZenSqVTGtfdQH5d+Ac6CnQLBBdV8K8Y0dEQuSMGykvlgG42Lpdl8fokKKrk9iFod
iuxLteuDQmQTsvpS6I9dh8AdZCeevVgVZTd4lGZoTjOYwuQX2sKcLSL95Fz+wMket+vaVXqf8rFf
jzr7ei74tdsPYLgri/1fmqDs067yora/ETDK8/aKBtn3TexSm1LeP6tt2XJZWkDOzjokDmbph1Is
FsRSk9/YgBnrOK39KhTVvTt62aOyIc6a2oB92CmpPKWeU3UPBSJYgFJpcy4b5iOZXbpXSF21LCiL
dxa5/dT9VvpkGcLOkgZ97CcV6Ks/9SqcfWuX0t7RUOI9Y4PLYHhjsAQVoxaZu3QLvpXcFfXuY17p
mCShqxM1kzPixm9wfjspyUJMJSwAvGplC7Fcd0TniihXdFN6KcpcCJMSF5i9BlRzP1hp9Xfx1OV/
c72etyX9fNvYBDX880yUT8lIsP4Mfce3Sf0ovbXi2qE5/719KbCCrB9B9U/hxB8EPT5xDGMu8nKR
p4kiOiPn8HOHDYFOJjVtIuASkRHujh2uYRJ8iDWFAuK0N/CFI9OQ6PTIriaq+WaVSHXqM+xAm5w1
lHWnkFPEtGyiphuWZN9x5/N4Lc/7ZKDOncHeVuUo4lOJRaxzy6s3a9RKp9MaDJGW55XYYCSuw/3A
Uy0IFX+IACXKA6saxaubEwywsNYLfFY1B9R0DeQHaNoMbOC4OhhwK9N8MdVdwNAiQ4BhqyFcrXs3
/5p5HdgX84jt1u4ZHeXhkWY0Czsb31tldTZbZLZnhBuHXWTJ4Q3h4ShG/BKpLcshMJ0W4YhoGeNs
M5HWWPcXMoRM/qIkZ7i7AShqHHc7q0cZMSVt8oYMfimRT8CzjaZUeqMGS/O7YMiYzmmbHNVJwNys
rQqQuvzZAGVYQkeoTYMjO94r+DNMhukntjkjOxv60ndUIJdMj35+KkJYALdRHSF8n6l6VKepCKDm
wL83FtYN/TIGkRAgFc4kQH6Va3kgjIARryq2WbediVB6o8uFiacQT6PYOCROosDff/1ofTa0q0Ds
qAxju1KlvvQZONbBdUDPBXBWC4n+OrDqZeuDJBFR+zV1mzga8b8xaTVUWRM2/4jSaxdOeHdS7+eW
YsXJ/TDLeXmBDo8Q8DB6sNh8JF9ZURb06IYoxAg4UPVAWenGlQnVX0klgvyX8IjwdyOizG4NNY7U
GrPjvNS8if300ZSUEsH/5HHHBNXFAPnUkEy+CvRXZkw8ES7lQPsypGQDD40HjhTwhqbszYWze4hU
CwmNkJ+iuAlqnZOFGV/LfH4Ro8j/YEMqAq6EA8LmUd64dMhzNMVBN7HXDnEMJhh3GQPoSUWIk0mg
Om3OSuXFRDWJmpV7/L+yqP80dMbxVNhl8un7cxr2+ExSvJqfvUyXB1YsdW62VtzD9DPBVtEJcEfe
gjjUcHYXCeNwgRWcHpg2RrJ9rX/bNapkceifPgU/amMIeVTD3WW2EMR4Afy70p63QQRzxwhkDewP
karUaAr7yGEoE0PCKfhOrjufcMpY4VxWTbfyXmNKVSdZffQt9oSz/SWb1XiZdCCm1i3qc9BoJ2/M
PKGmTz1oywWO8nCnWuJQCY7AAVsMj7QqnSiZ/0efPlV9ASFf4YhDROsfioH0OnbX6NldAA1uma5r
5vlZjljnYScRH1jyQWODWpie7hPpSldCyuglCPjpWQJKjPtdIZo+8Qw2k4FqfY3QN/PkZZDIw9HW
3iVLkcu9eOpnSHvTqiY1ppk2Gmi6c7CHPhknwewTFgZqHQWjPjteoO8oAOD8rFWK1WEVlsBxku02
4W3yVmD8jH1CfRBvrs6+PgrltbA0kopxa5FGO/vJcS168X7OgGZQKpnlTvrkbae2rABmsbM2ydkm
PmtxHDC6EJGXyxoAGdVWXnjSSmAOuNZQtCEvPZOgPnBfwhFwyyf6OgQ05ly3Y+vxU9Gtc5EVP7CR
QdQSVjH5unKnSEqvEfgHHCorfDr8wj1g8++3eGHHEhfOJt177rz1TFZP2dVn7HfOCb3PEpt44vVI
E/X2KM8tYC3iv8Vz1qxl4kMzcdgdh6D1HWz/FsWGstqUiHkc4B+r007jYT7vhrm04ZOVGjNHtZqW
sp12rpPgl36IKPo=
`protect end_protected

