

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bvOwtDo+u1XQuHmmirIW0G1Eep8h4q1lu6sagQVNOpqoo1dUL25zlZCKWpryXBrbavlsSVZj+/Kj
u5U6Rqq3pA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R8VeuF45EN20zhkGmJksRGl35KTSV0YbXBmOJfN53AFOKNxf64co0R3kMl1KH48vuem/BXWPzNwW
17k9On+EP4ryAUZ6V1YvtlO9Er2xv4nZefuEO+pELxS67R6s3b0HhdPIKa2fxDF3e7AwjfjDxMiG
HOQbqK01rVOmqe+2yps=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qqYTedtVydnDu0uy4wgVS9xnI5W4e3CBu2tom9I4ji9x6Du0u8YzLw4sHBXlBjTr0CIBWi+453uv
6i+HBaHUw6WLmgP+uD0PvRoMp9iMm4rcTjCZCtUo+5bxaKDQQyKy3VozWJN9cYsOEXUyn41sbHk0
MfnFQ231FTzHKrD8+sW8iXzJhrvAxVZSOCQNc8FKSuvFHDKgrQOZi/Dde7fskgmy7Y+pQzZQUv6h
7xsxzMyVpdCwJjhjdow/xj17Fc+yTtNKSxkHMIxVK6RXkbOidb7jBkIw+8aEzlqsG5f5vpboGqLH
6uQ8IqqBeKv3BDowwIwUDotWgCgTdyFmv35LwA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xgoCG0tChkhv+ljdCxpV0I73D5nOgliZqF/G39R6pkQNEQixpt7jSEz4sP4s78dR6d8BiB9A3KNg
s8gNghB9SqKmhRG0Jvm/hSIBQCWAqWOwg26IvTnT3j3MalMVsj1r5WE9uyiqdJ+QCTo/Y58NBx8l
pM5ABblrTJM59LnIcqI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VTcA7V7opij8+vJ+tjjgJGiOJ+o6V1u444VHa/k01STvZB7T6/Ztq4KXHSVmD+driESiC+2EQRes
dfVcUifCMaPU4kNZrlpS+Cz6GGzKHuujVBDhNOZum+ncGM2VGmayYd6F9EbhwKFTOVOkQmEz/eFL
4IAryyIE59LghhLnEgKJ/yOFNS6XwipLZ1ztAAj7QDruS/h8wJcmBcjwC4vXftAO79YXKmVgRKly
SlrrXAPgfawAm5V0hj7SI23oHUFrT671NQiN+jfhZylivDC/aANQXHsoSuY7NkiKvHESuXKmJ3iX
cfk8aGjoqSspgWZUBuwV9vfaTHDt+AtBbt97TQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 174368)
`protect data_block
ZHU45LnwtmkYkeHHnRPSmWYZTfLDx3z+h6gtwQccK6PB5IqSBrhayLhBnMXkjxP1Zz2wFFgnZfQD
A7XvGI4IpI22ULr7cAPmcLkRA8GYCAge1CyTZLdTvjFEbs52cVHJe0yreyc5y7L5Y1k7/KQlE+p/
Bx7W2rf0m2i7AuliXZp9l+k2aC9EKFlXhEQPxieTOtCiopBXihl43KaJIjNz7VgckNmGTlVLvGCx
pgpYOPW/kYpWRz2vse5MDA+MNKFe9ueOXXKPKBTsI3ah3nWo8cuQBoIc5y8pZyJruxHz2jL9iGQz
SmT7vHxFEU+vE3uaRyNam8B3U4EnjAUxO2IMTGkCXo3XfKKozij6SgLAhywfFXLxn6w0WCr7M5B7
vAvwAq0ksAxJzRqwz4tci9+nV0SR7warUAn8uzXf3JP8zK/c2G5e4J2S+q18BFZRelejI9hmd/hw
bAD/9BNIxgUrFG9+ISJvAQX/gK+PzYYYtaqSWLRGRQtqefT9jrRzXe7tbYLdhajjIg2Zo2ANuSWx
nbk9QYIvGAIMYZZWYt3246tohrAY15AIwyD6ybDvFs+EcGFxONrzTQCJNzvJAbTkNzBfqXJA+pEa
BOeQ13mQLUFPSR+trjqM3ItS7N/Wff+T6+ATPD9EU2QWM/rcdz9ms9/8/ZU8cH7Gev7okQpuBgyt
6T7xhqKP/0cz1STzqSs07zKbZrJArvj/X34jIQ3q7s6rYHRR8GLLBtc+WLNPbuU6V83v3CGXoIPr
dTpSnaHM5fR4Q2qlT2ZGbrBsnjG+KXZOrBoY1mxG01fde7qLr6xIJoBEX9blAirBOt0aXsTjXV4u
ulL1dcCxbt8H8UTn/fc/dNM04QOKhPlxEkPcFUFTNHuXLLP4ae0jfvt8biw48YKMCW19qV3Koj/8
wZC2R1i9h48Modb3ZzCbdl90/5YSwU/gfvkcMkLiLzYa5oGogIorZEJwVrWGqrtDcAkUyy2rsoeA
Vn/k+lFM2qJ9rb0KEggp1tHUir5NIAjUxhBrvSiv/NTJ0fB/A4COmzv7lIdytkxi4rk9+pdhpHNZ
E5kNYzPKwg2ehtdsXGvKHft83NaskK9XV47H+kTfWOynyeo1PBt1gznVxDbn+VEsaBvcMzIkuocF
McyckK15lQLAZXghXQ5nlXo1oxZc4jHQp3jdTTKO4UC4k0mo4IINoqZfqjBYqqRrySFlklbcStQ9
nvpaA8M0f8iRVG9yDmMio38RGU4Lu6enyam9tVvK+k7HXuxaceZT3Zi2QYGis6A7EoFRtXtOK5Cc
SS/sDL7IY5KgPIMZaB/2nC946HKNMm6OD5KbV1cpvMRMLAKeg1V2CxPgj7DuoXMQnZ7gOCmoV1+s
/o818S3jBIqzyDRUpWNWuz5/RFKZ2nIObbPcWxiotwXpFEdlHtPIUbRnFamCghSXE6WiIlFXlPBM
Axut1rG+aY09O06WhnEe6FzjKQc4jtSUVxj2oF1xufO/qo06Q/q8hrpCGI+//9XVcC0bFXXmF/M7
DT8Qv6qt0LufhjRsOcEqvNdzDLc8SSGQjYeoWCjAEhVxw+llfALI3sS9dgFgRTjuo1RAt09SrOGk
MEjVr1Afmxs/h/Kb0gG7LOpK0JMrz4IGM9E4TYrXl/1IDVvRxsMVtL1HeZu101ws36KBXaykH7+I
a8ixVorrvOQmLw/ZIFQ/kkSmmLL5F/lkKZVXSrF0L/yA1OdvhkmRFsooryPpCvsBLf+Ptvgtnzzi
mSksdWiF3OO7MrQRQVxZN96W3MOGu0ad7FhTqa48KrzafpfwST3bgR9jhVSSf3UXOu1uZ0R0o4Nc
3gpbsXy2e8nSPSxtJ68OyZ4alFXl59TUrG/TTxBFtt/0yFYJREncjqCCL8tL4dj70EHF9vVWS7mk
pU2DUEZgn7gzgxOU/wDtk2We6j+5CTPpMUqqxtWgQG6EcAvND2o1PDA41AFYy1B5SdnYgnZqCgeQ
UfbWkn5XXdrl8LIKX1B6Z9MVnM2vAXzuuMUI60ptxlGQv8lv+GzqkCBFSW9ENepzRYpfJ/dROdZt
fDFqcWe7Ieq7GNneJSDxEJ6oXsQ1xd+WUAxKvO1tF9ezidDLKfbCd7hggKD/LtW4GQrXkM0K07gs
lQBEMj+0l0EdNkrIV+y1Mwd0Z9lsY1olmcGmVmLeuRVYzu1e9TYIjFUFXgAWzv6TcVgaLFNtZ8oL
3choZ+A/miRNjna5AVY9v+dg4dRv8acBjcB8rj6SNIYGaI0BLD+X6G8O2FAimerEKs/ZyoMZ5MHz
dofS6gKSxHekI89Xa0G/2OMdNo8OuQc4CgkjyUgkd011BS0H6Wapdnmf9EVbWUkoNmrQbwcGh/oQ
xSUtBPXzikz5ZdibMao0eSGVoGkxd5blHS8h4otkW50g5oIM6X5TYBrU4/VGFHy4Mr0Y/jtaltld
qbTSm4u8+XfQABVpEXVqkwyhC6B8Kh4aNEPiUBg7QSv+5jqqtbXpFEttE39Hq+WwbjRFSiw6SfjK
mOyYK9nTiEsWOS731BzHvkJsl2d5V5IZCYSNVNIdMk1xd9A73Y7SggyiUg2wuOWErINdTbi4Aby3
zA68/l8u+BI3BlMrXLivwDIgyMlC2XMoSHuEt6kbI+1pUmDGu94KUDsVrYE0rBxWTUTuV2BTNVm7
tPyjAjBVJHied8IUlQLng6E5uhlUbnchVf7yMGCfrgb63xkrUGFImiiKLexel76quo7UCX6DsZi0
Rr0El1AQ+pXY0gleO9u/YkKo3bIWEPHMqWU1ckyfnGFgKs8HtWlRt8+gmfs6maeWLSt88GquHS2A
NxX0rvppEofMoes7rLrKGP/GODHLkVAa8quCWNH/OqlakcMsskDUxltoK7tyDQ/nNbk+ns3nVV+p
kXztuFlLL7TwlYnyd2qNwbqUr7/ymm5DtnUSuMi8hS46zNj1bdIcDdeCRpJOY2QfQUNoW6IRH0EB
cQAUe5L3xUGVfPmQhVRTk3AW4uI8i95bdXdTIFuOnfh/h3r0Z7AbIjB8U32QAWyCXDq9tLoFT0jG
xu9KJpijYLEPPcac+JKNNVtBoxD4tc8np/xlLyQTvR7FGqt9oNOXaqsSP4piptmmlUyfDzE3OPOJ
KTOnAgylyp+mq/R/jQZBWY8AvuBiOHTpvJKFLMDOjvCKRJ/E91LEHnOhyAyUQJ74Dlk7dPVfgAnE
xF3aZxW3fjFZ+WQbXPrqBqTQmof0PaKUzXsHW9JS5YnPDnVZ4+cx+vJ7e7Y66TRm2j3yn1bgXVKA
bRRCLGIIC6nkg5hOWTYjVzylHH2l/CnXmYoZwRVrwXkdIJreQerFT7+fEOa8E4olhoihnw08EJg2
DbeyJB+wRbHmsggkm/sq7gZcRwycaV+BS7LXb63kkFpaChOQHGKJFQMogzlXjRqfj3lTgi+ZHt48
DXI8u/VahNvELHMbE7gjxYnxTS7snmPWEkUMX+LhNw8FYBWKtwuHd955+HbsUpZeXBHmtnCfU1Hf
GFOHTPaUzKg+50qrcAI5Oyrfo6DwESa1HmzCZaG29XIeLUIMF0CPt5ouMQSdFWAWBa/aXVmg92Ij
hHIzTGaaNSRVfKvWoHgf9RgUzkm2WU7IafQGv/GD0z0YF5fWpc61L8Ew2917QbZcHKyE42VLP/bv
T4mXtmfE58ysTBMOTue2SjNnk+gHbcdNpn0AzpGEBPSB0spz/l/4OEaoDKCnhQRmz0jGYURHqOKv
N7BQYXGJH7lR60D88/pJww45ft+xQqwuhHlb8eLlp6yjSdWywaaPGJHbAX+SSTDYnA6DoqiqRa64
UignG2AJW1/27i1wi5on2RBYYMy2PBWaX55VUlrm5of2OEDBuPyn7uEPBf/hxPkg7yQPQ+QXYGNX
ZDn7gzco+W7ufjnggU1TWeat6IzI/7i6w9PYBdeq1W5xnpeJrjEk8290794Mu+kVpDJ1C1NAeMrC
iC/RSxEUkZjH2hecqvR6O5TXBm6vrsWHm+m9kedqC5yooY/9fNR1vuzwPOzReFp2f2i0AHRkp9fC
XKqnmSzOsioI2yUGEhKTxkcUaHe3cDFTtp1YxRsEXlur28FwpQpFIDVptkbXGdf97wFLDo3tJP1u
4uPNGqCZ4aVHo2mDCBDBsiSB3mGASaUGl2JvQfB8XXilMfRu09iTBJ7osOOlGgaGS33SFqpZLQWY
ulh5/rXJU9o3vcZkQ4JEjcBOCQcY+bR4exgPdNRjuV7RJ0u8sssgUqUbxgI8EZN6fj+6xoOoXmh9
FFq0xOc8ZteT2LEfPAvsSyQsqkCpyl3AVX+BJSzgc10xTi0S1idl9n7kxqSl8wvPe0JzvLFEHvNV
HYnN+fKZBrJlOymcEu55kRi/tt21tA/o4rGUxIHSbdTE76amY6ot/3ntbSB4NpCE+EbF+x8tnwry
OZXinT411gES7xEeXFIbzcAs6w74D0UDq1+p3IjFXUCt1rKjGbzjLZILxsRS2NnLsHdV9kymrvTm
F1Xslmr4Q04nXmuMQOAbwijVKmjgMyo00lRX5qKNLhD68mE9I9IHldK9U9PZXM3Pa96EHU+LrLg5
GWslnoI0PtATGpQE0ny6q4AUFieW6YVZPKmisQnneaT5gUYrU8FvRbllLpf2SDDU8YzEfdR+3srt
Z8HeiugwRUoguNcme80UoXxRR0xNlYMOUPW8xwP739ZwUzs2KFfDdgCkC9Fg3fSHGle1pklpYEEy
nPges/ZvTjNmIdRWFONFJ1eEh8nb+vDh9LD+prOBHKbIDaMI7p9fSXpUTGiKGD5dr+BbtAgW+QYT
0LNSadv1fEzPim7QMf54Cw8JWWv3gXkd2QT5lszC1RppdkVJ0dFN+i8PVYQR6cc78Kk5mhXxn63g
tMXU4OVzLv6U+NiHSlfC1heQyiUmYb3Yxe2nlZeEzKyhIgBHzUFnjw4+GkTR1eTgwzXJnGX+WzWY
HS+6NL4W+NYD48hnX9Xct09nVh5HBk6HAro0pvh7fGls1sZ2X87Dymtp55ggYT9yTbJVYJ5lyhm5
e5062JXhtbThR9HoTIoW9YK26Vea/dkUWSGGhsLvwikiEYg8ccr8B+hvbpJqkqVor1pivuVRU0MV
9eojBE+OTDkEqOn179gc5EoHVfauRYXsmCgwiTgzO4WAI19XL90LLq4Hagflov67fT/g4+N3FsV6
QuVK8UnJ8kX0Utr36FC1Jqhs8AFbNR1Wd2gI6wXeU6eHukZyMNzrPmKxUZaIfhJ/SpN3txKvRBcS
+5XGYaANNekfQn22guqIhvw7gOfSMmSWXIx3DEpDXD6ZzY3wNLW8StZ1ddrySjkeJ+jQ+JR+vjXR
2AJhaD0C0idulfnImG8w8dpmxGjiemjhf/1AhxIbOzEf/hAagFacNC3mGHuDo1+aLtFojufnzoCj
WT0af26hDLcRgXbngFDs1VVhF6O4CmWMBS0BEtLnJPn0eqUit9dCpQzMJ0/h9sGsYkkMkDCnqBd0
Q19NDQd/Ma86qqRTZXGjsMkSiMc8SMKqfpWuuxTaIiXAg46mdrZ37KoZLeRaWXoEEqJ7X0HtO0Ln
4gUXoz9NcYXgXD8GSfuvXsO/9Grn0hbs4e3AGAMkMG1nQdfoxg7ij+9pNQlJVfwXPlirJ7AIemG/
hiWJtHrL9ipsVsel/rM/4B0/we777k8GRUq7wJcuhxjBsYB8794ELvFXaEvWnoislax6/wpsCy/K
zxv91wGnJqxVKS0wsS15BVQcmZY/46vBy+duDlVse97Vzlc22yM2pedqMFmGWYEqOoupbYfox4q9
4WeDHOnY9wtLVsf5CzhQjOfb9eenTfNe+2U+0SZlSzYdHMJdMe4sfU5CZNyvuE9X4DhNsTlCSPVG
+kd8eotubMAQbfb3zYylfwV5irCzS8LQPcJyg4Dzk+G0ob6slbhPgqjwRovSlWU/s13/fbbtxcbh
jFsAEgVtaP0gwn6Zxvc+Z3lE+DLVfiqPMnEBgx59HCWLTWpfGWRSGorCfwqgQ9r9mNPAPcKpJRUW
PDlCNdFwnj2Q7Wwgz6Z5iUpUlT61COCviNyCU7mM3RAKvLu+Bq3Io6cbRUxfjfSeGQARh8VpkYtk
RnKBc91DDUp0iy4awXoCVoMVpV0jfYZFZXVWCcEM2UgVq1Vrlbu1PzepQjVtLNFuujCdmFzxjMWR
xdeGpc3Z7vBsNjCocodc5znpDp0bLAls9FVEAkASu+UN+FI0PqmWVNBwLpFoNqr/BVWUYHc3BrKb
Tc8kRXReD5zmQCYfowoH+sKLeuw0GnPe0DWHAzj7dZCF4CmkRhA5gBDU1klU6uZYVKq5Pff6UwSc
5AbWr4SnBSfIu0vCwvaF2ndrnUp1KgOSq2p09uZXNNQzdeZheBQUqSq8sp4w6kTqN2dedY9XYsdQ
FrUBgHZWVmQTGENzbg8l9MP95mDbcagAYQDqUaOfRG5oNCgcyTG51H6CZBaqoQtvfyQowA1S6izU
dGRnAxC7hZRiOVXyPI16Dipb7x7bRLeY0c8UdOq0eCXbHotky0GIqGJZCivLl2BMNXDnM4jGx9g2
4q4eTO4D2ZWdtcJWeXAluJhy1yPqRFAcZeNSTnODzYbXoLD7QwaqabU5Uub1Mxks6P4syeBO5Vhp
AZ1cPCKLzsliC8sGQMhHv3bivDPmDPdQaJ1iwKgypzZ1EzxNsrfgKwLoaGOPlmIxnFnXqifudjmh
K9FCfpyWkYtzuQWr1zcGusAHDyLxN0ZNgiJ6E8BkVRNswaGIBwCis7oGcv1ZGmbAoIvi7ph8Ku66
sbXpVpc3KkIFkFY/4VOMIS/lHPgnOvexxCAiO/LWVSnf+iQ+F0g3u17EUfUBTTp6XKJf9n+BVyxV
Ci1g/NXkthKXNOPnM79lt5Ml27auy981Cwqqh9DbVmXg0mLxDHj6QuSBZo8MWcuHbtpjaP5XI4RR
q/MsGH5aa1v7CDY9TjCJq2veE12of2RKnA58PTRLKe/dNFhmG9O9hr7Ba3T339RrK1MkgKYp7s0h
yW1L44TGYW9Wbast8Ub1P+u+tj/nFsJWDBeAgS2qZ9m2CcKTt62CUMy9Eg5GovuVoq/oh1opefGx
XosLscpKdPWFjNK4/Pe3mdSKOqWqUwVKaqmumGfXs8j/T+8aQEElFn0jGVa14cyef1dQyVPrQGZv
3C/sHmekc+QuscJAMbU/y2YjCuJhE3+eQ8/QCfIFWlhNqEnU8NqAwzwsnVCrx4UrqkkY/pTnNJN+
6AOg2y/gtkNZqY6lxm4s5WGlKSX3acRxH2L6utB2wKw26SZHstmNgrBoPJkb+xKjBAtPqKhud927
cqGXSCpslGTVXjw1NcRA8w+4eqBMCGH0oaKz3M/e6WDbBD17AVMkMbSYxoxJecg4it0CGq7LTerC
vJy5wlIYvA3eQ74WaS3jfhfBWuHA2zHj1qlKLXQDUrCHE/0G98vwewgDXJTBGoAea1d0i+1JZya4
eLMrmHusTcFK4k3AsDYNxkicqZBXJ0uEY8nckGFOcx8PDHS/eVRDu3ehUFI3/Oi95jxm+WNb7caS
kso3MXX937NheH9fWnjDEG4JgztfiZxqb64HWS3WYeTDvwsuxx666JX1dtboGQwiL7D7IRrwVRVN
mCgEo3QS6SGozrwzdd1lBreXOXID6jZ46iAEVFkvUSyLb4dSj65oilxViYe4BhuGL37+ayaSDxsq
N+mG/HMlQKSLKUC0Ibtm1P3utGuIGkVigA9wK6qmYJohRYt7V4ZdKN40HCNn2eI9+w6+Hqf6crDX
YrPKnuFHKEsyRsiEKwYX1HWduNqqhz/vrUHnU9O77lJhLFCRlOdbXmUuZH0styexSM0vRDYwDxN9
85jKkfKRhGkyxRVWz53P9DUMw/iQkD6Ttw8K/IsZYGF6F41/HyRHIE6Oizv1mHaVF31Iz5UEqdUB
shtawb/R3RazkZftzuVOmcDfc2gJsjg7wgegqD8nF9QJEYr9sznpDEvelTIXnVFkCm21y8DNkyoX
jRfYZohOQnku0s2deVW9AkHhx5s7qvSG08avLoMB8cVWz0XGpP7haTS+OvZt/3ghZYvPhY1t8FpJ
ZRfonQzTKlGqKZjn7p3PQnNwK+f6wkVRNLS9nPl7SjzHje8kYRV9RntyvtMXID0LbMIy/0rx0sZP
trIOtXh9RGEIVT3lUwo45GFb9UOYiiiKNJ2B7pTyBBHNcEn/Z5ZlHdjkxPH+IO6xbdBwYbRkCgte
oVkS7Y1ctbnPIFNKtyyIIm7e6UBr9gPLB8ocCvdSHuV8b6a1bUVkOM+IQ/XvVq9n41muz/lisHOM
jcUEja1maAC3TtVqRNun4axXuhM5McNH7BWjR/GkztYgd4139RGeS4hc1fLZJSmE8Zeuv2MODiem
gdsl2QZYy/kJ7FQhmGJxBU/PUMI6fX1T9dYAhrL1KmDOZKKsiYYejwt0h9gTn+o0RNuZDua2UpPB
N1uXm4NI4Rj3KU69dN7k9hBAe1km+ei+JCo3k24nog8EKGswkwBsqM3cvJZfy+MKEwP2Kt4wHwE3
P7n7wAST2j4kHBR9Gh9sr5qhn2sZVRbsWAVP6ibqFq8JsPh1UqkHEI2oXNvf5tzWBD1cffqi+aPD
ezwnp/r4y+fr6FLLILRe5927EWpnHad/vFKG4ZU7+dA5iHUO4iai2uoiS2J41OK0OzdsMynD1f4+
i+pOW/5iSFO1ofNbvdOZZ0td4CHLliKmvCmMxZNvWzXQKpWkPPhyb4U3Z0lhBMmp7rZ6ecZGibDz
zpLnQXkSXv7LTFaE/BbqNQqcvOhvUxAuHnP2UGreNqNVbec37iHvkt2mnFgidj5XnmuQdjjAKo3a
AmL6YmBMsyEy6LY6tLa0nDkFeoBVAXYlRa/BWL2R3rTb3fhA5p0oX+oLFr4gkLsT1AR2YS5ef0+j
XcaCzBeqJCshpPv3KE0AvkWJx8xw3Zf4gi3jkJYPjtKnqMpzk4DOMfA5uoj+VA8qONx20nnJMVXp
ISyFWXTJjwXbFdDLXdizsr7ZjFy78/ZFH5saffTe1F/zy8rJ3JSPbuEP/SCymxrVZF9pUiLEBwoi
D9piyq2SjYdAy1NuV/bVU26dLT9/ZDZzVtfcB57yteUk4vtJnqZqbhKvjS3A9OCvq/HdqXMQnMcY
XL2VTPwQKOHp8/e6CryDfXc/LsEJlX/CeOIrTdV+fmZRSm+yr4DCe6anJxBUUi7MrAqIQ3lYHBRM
4M3PjSCk1htMkaxVLd0ojQn7inL3qBbk9Hi8tiiYNKIjQK8ET+lRFgKqmB6K/9enyAFuNX/c7GXs
tdVsvqptSJPUb/+P9CM5wf7qPopu+ecSagM/LAFSoXrFH/yYbmlv3mtIVIZj4BI3jtP725QUndOe
Hao5jZKOuZfqhwPHYM+4ylitXaar1pCcd4+v2hHJMZKEo9Ux/vSu4OazynrSGlYJRf8yECzSQkC0
6r1d5Bwv8wxMUODGWx2XCrDVThdbEFnU0jF9c8Vs8n22RttuiPbl3RVmRR1/vJ0UBjaCzvrsRoht
zmFB3e0zmMmMJ3xankECyzVHzOFjjp+BdUP1JScvJEfe0LJkSYUNMm299qOMJiftGcamerP9sziS
i8fF0GNH5QwP5BqRfxTcldiSSS6KfefN+FwVpode1w4AaKuD14MzvfKkXulY1EJWtH1KW6Tiy96P
+pPl9l6oQF7UF5bQ+kPPuTjqYAXH1sjfcKtBC2ISWJSIRlTVHNY+iaQmQxk+BBXMQ40VWvt0aT/a
eD9E88bbd6qRx22iCZzgPDVPlT0TAceeSP+XkDEkbBQXuXvr/KP0H+2td+bghbnTcLP6P5DJIuw7
czd8wvDm+PH1MiEUAlZe0VJXTFlPjn+4nrNNA/q0LWkmXP+oefLmx0D+GYWgKjDYi9BNSfu0VYUL
FcGqgh3PueRRfzarqGvYHmTwuph3UFFBcUt+YzFQELjWuVhl8eGe9Jt1Ikn9ywKPzLRAOvrHqmd1
UxBK32ocJ2rY7eOo4D/tIS7BaxgryoBOY7tdbNA6rPNzaQRVt9XkTOP4VijwJgzDD7NrDij6S9fA
2A2ULSD95F9XVdb+pAbnTaWDKPjpwZbgolFBXjYukQVnWr9P8z1Cev/PDJ8i5S+i1feBpkUSnuw+
tq6sJM1UtiEAZkzv2BlrhyY6vw7zEYr3t107IgigAfff5sTMm+pHdc49xBYsCK69QjNxtamvnoZg
4zpgouwvQ3afRev6fQGerjoEhOfp2J/aIF8JgG98LXDYGY+qE9yNqulykch1T9iS8UetIwb6Y0OB
1G8FmL03xh1cZ8v2XTm2nBfTxvAYOq1KwarM4ad+VNoopGlw22cPhm1NFPgPNTSmQTESt/igCVFV
KdpYggi59Jd2U4h3+EVS7GnhybaaJwtmJaeF8n2z9msJzssZh4X/iQ0de0lZfLQtEoHSqBSZOCVU
xbQZeYe96B6uWuf/AAv+iEltSbemh5/2QCGX1UbxidsturxVSR87lrFN+BSj3I8UZe8MFg6BPjqN
bR9uWpAMQzEsbefHsskptxs0CtXhfDs4WTF2U4pc2aITtOWEZNrsHP4WmNPCU0YBvUchFxrIEs0m
h0S7lD/XiG2Pqd0/IpX/+Kb2b29ap5gNzGtl5NwiLv6YBaRgWjysuogTDy9H+jBurqjSZsozDl3r
sLX4E/ZWfmnJXzDOAkI/hycXtEfhM7o/9E3wqqm3p7OFX9k2FvIUKFarKTdNytCOVFmS9+ThpVD0
thh71uvNbjYLVRYXV6oVSL5DgK8AmYfMIz4l2NQ+k/Qx3v41816fS785t/LgwP1R7y8kZNJNcV3+
mmCs8ScfATjD6Ls98TYTqlmCmpJG1VajfIhjk+Kce0u0egyxkV8I277Z0iUgS9wlEjcFtpyoBFU4
389cGnY/YIoqoAwVB84GZHACWcVvqJVlRMvHt9YmKkJfQKvbYd/8M4ZDhbCvEOg53txYJ14A+bUW
9wMgLvR4hgcfMKbDIVgWNBD/1v0S9bnbXxHYWo8tPWnk6+5HFOzWoI1SRKJPQiM7Y377IygSWVEN
jzWx/8TbZw7nAEF+bvxmMNEzqycjCh++5z+vEpqBVBupGoEFNrGHXE3i1nm63MVuPJfPevlifMD6
YfqpG+pRSul4rIHchey313hpcSNU7oBhRHdJFsPxBrY1spFc2gpfASe/zbmEp5Mj4q+55oto722J
kxo4eERmWNzzA9wk8Px2bAvyy847D4DCUao6vEwclJUFYit7pBdYCouB1pl9BN4eyz6cUrQpwMbj
0hgozKqXbCc8hQD9ybbxdN87ex+YH1MDsWiFfeQ9jfcBgBL++b/Ro72pDhtZeWGedCUa6Zbg8X7y
e6Z7u8sxOh/Gjj2VmV1p4FIcjLSqlQnVmaJWfwBA6w8z9ZpZVX6kEUFIT19PP3Bkz2GbGBiV+mc6
HcYN2Q/yP1kH4VFm56DNHRPyr/oxo5zjXC3oJoOC2TL3JOTdznFWn9tehAp7YUVR8x8oMLMpRHFV
eC27vRtGbD6b17DwDM81GADKbJf6XMkbSdv12+bMtx1qHBOZ8C50jpeOudGsAi2ZblxPD1B1PnQW
cjF37HRkrNyvLvMfSO1sCCcBgJg6rJBVTOcbO0Sa6Ot1uuC66Ua0ufalYuG9/22Mu1CJqWJENR+I
9THJPb1p8fpLNqhuiYGHdT632xjaLDz/kA2z2ZLK6L9N8nyWOMrSvz6aFUXivZAHzFQtiikndPEY
F8PrrwueAv8eRwDEP9I3kcEGB5LmNLqqRuv7TPgmk4lM3o9cMnjXsZALaKOXPOky+9LoXftcitcZ
8DwjWT2s8f1d7TkzW7Xtjg1riGtR40zkxUoAzhaJss8LIBndWYq+WqLcuBg2q2Iq1tO8BobFb2xj
44BavxbkuHVyYjdNSXV9QdqOyH/k+IwxeUZ4loa5/nna0QbkGPzg6PfDmLVPa/t7NGeoieKz5W92
47IEHg3hQwgaaFW4UFVqPly4jlBiX7YMRe48dmilvNdK2+DL4qXDWQTi20SCwxQCKOt5y4nxw2lL
O0YLN5/F91PkpRctPGkCkm5tyE5kOR5Vzk281rj54VIEJOWQ4yRFrBAKJ2mmtq6U1PnddXilFcCw
37FICl3LCpbwDGdQaeeNrYEuzUjAKyN/N/ip5V0Raox1+hLMJsbeQtJdLukjyD3XcPf9ZkF/7GKy
40cczCZkEZh7yJW9jrTbBRnHOOGRMGtf9AC2ux8j77Moue79pgpoeqolgmSOGp+H7Uen4kA8wOVU
MySl1XRQANeJTuQql+EWH8GVbBlr9vlbpaVhPOmJtFabkCe5CWiduwKOQuTpkLzrw8rGg/jdglhU
elPMStG491oGJfmSOAw9kbH1G1BEsTEYjdkjwPoVArGW71O29JS43VYAn/X7F3rMDh+a17NL8Coh
Qr8n6dESLXagFXNZPLhKBqPDrN9iWBRLAynTzI9HtoWVKv2ZD/sII068hmfxuxUNfjfzY7Z/KRaQ
Ujy6Fo+3/yXO+Rq8ZbkMw9usKWXVk9eTFaJHVjsmZ0C0Z7k54smRq6WvmbBFSBzDnBLWbdyCoxna
eqoiW0FGtUoNw7LH9v90mRl0Lm0GSTMzgBCZ6VDZJhKTKgDl0/HVuaz3AqyBreJe4tbv2Kha+DYc
yfGM1P+zjR8TXNgUv33d1Ln5ykeNYQ407EO1+w+aAmv5yzZZDJMt494meeibtTpGP6g45qGeq771
BK2UIS7Odjd0qTxbimFMd8qdkejwzOkSpQH5rBHVgBBynUA5rS3HpBQd7Aei5FggAH1vB2TWeOMu
kLIppZzEZ7WORmPI9DWy+AKIyZUsu7S8OmtT3HZHU4gcEKeGY9j/dmYI+R7XBuLBZLqP9Zxk0pmy
/udtnfzfjbHwmbwCGEzuNBeQCVzBPwLVptBRQK3gij6AEFIU3Hth24XD4X6o8al6g8Al0Qrtfrv2
ndsaB2YRksxydGD5j8gNnjfYeY34K5okv2ftazYvGWQPdSGSp5LYrgcC+khpV8v63VDxkJjLKrlF
5M6P+eYXa8EIdUmgbRflz3caamljhAGnHFvpQLY/EKFMekL10Gd/OJF2epINik1UnOOxlFkv7SVH
MTSvEP1Lqs0Gmji2FLYvTIXOpbPOLJZLMUrdfTESA0+0nLGBL7kXwU1gEf1aXMsCynup8kmhbRmg
ZudWrvn4s3KRhHRuS4I84PzouM9/PqzPBh+YXuGgP9icuaVo9evb6J8zwzIw7X0P1Qe0grau+M57
hBX9Z0RWi9VEsZtKc+OmUARb7ZunN0Jlw9vH2itW8rw3KfKpVu2E11Uy7awbGF1vVCO4gQ72WJqa
oh3Bot4MMGQrVrEKhQWkrBbLTeHzKoEC/cpT1y4WQLivxa36vL2rHnZT6FS7oOlCrw9QyCwNuLtc
yzzGmOU6+Op1BKQJUYBiLO/MmI6/TWBjRRrFo5iybRH8ACV5do2uB3ifLofc/opxFkc0Zg685gGS
+XUkcBg7ZZret7pO1IP7FH1HCxk4kbg4CPlYFtJUCg4zIMuMqpB9cK0BwBRAOkUsIdKCRq4qf2bc
xq3YLqklFErWlUYdsNSEvYU9qLP5XD6Hlyw6MXHtk6q1jg2D5J9iyGJ7IM1lu3NAQSKScP+yLw5W
cqTyTTyWyzd+R6a0tch1ipudFhIQMwUSGPi2ugKSBNZLdR4aMsTSReh6rDnKh2SiDuMoMlBeMuXs
w/EQXyrG4VSy/1MHCHsQ+/Z7ayZHSDjJMH76uM2EIkpRwb3Ogamvhj7Mj+AmQ15MLm4inmeqq2ET
y4m0HhWJw4NXGBeM2EYdcmbW0zUfTTPs662Ns5vviymR1U+UR9Eu0TlW1KoIvoek9YCN9b73avC3
wlJ2q6p5ucAxA9DNqUKOYu0wJnTNU//xy4ypwjJ1/RQoBhxOB5xHdAwtejRkkMAqAOE5d5OEeiCN
bmo5tpFLvqC7WBXDsW33Drhh6N2Ypxjr/VD0ZSw91pxnHhoT/t0XUYTXT6uHNDAlDMo/FuNniyEx
D2YWExRVY3fHNobRkTyyTz4dcVjaxNlP8OuBneZuB9ClsPNtcv6MNeaC/hSAVx0OIc4TD35hPw27
twsOp2dWadmv9U4dEqmfAJ2wbEikpDg9vgG8Mr1/KYZ9UmF3tJzPF3lRZdg3oc/APmElCCuaRIIN
fPQCMDAbKbaX5efXrLZN8YuKtQ6zfRm0KEuUkH82V6OQV90P9texRBHc6Tq+mbru1SVNSsQwVY9j
VL8KBwES6a3D+wDztfLw8ZPkH+Q+aV6ljfvWXtfDW43YrLSAW9kNF6sShh/VLYZh01Nm6ii5NKAh
BeTdOGoltw6D1D6TRtgQnqoMc27mZPk61+JScXwPrf2QdlEiktIEUkmk0oakxwZLk0R6YDEE5KPg
vBgsZRPQrVHhpq+ReHALG44KuCdc/UR7YW0+cjgIn2Cy/Xt2uornvoaRtAjQDTTDtZN65e3LK/dR
ZMjhmCgChYPPG4vYFI7olkyLpjNVPUUdaCqx9B9zZqQ/6EsvPsrhsWQ3lJV0TdjcOi8pz2h3zixy
mayGz05MilfhDBJqPmewTq3jxinpEpuU6Pv0ETU2Ho15Sw00viNE8qNgCpK8eAp0vg+x1DKgK6Ec
5ygKQCQ82PGZJTm3Jubs8ymni1shj7jE2M2JHKYQR6YWF6+oyifSzOJSnK7nCuIH3usD05d8GoBF
r5ZQWv+0IfTeYpourkdQ7sja/6JnM1mFKXceZL/YMCvhv+MtPcssHIpSXk/ckGJEeA8djfp88IAU
Cj7MR0hw1Wir2HfSJDB37SjSom5/AtdZNcUUmd469GBMpOosvsi5ZZF7m45tOTEpM10PaGsBYa+D
O22C58gFpHDwP29D6q9/nC4SlEFl+kiFy1lJHbz4VpxYI4w8qOQ36xQ70oKtN8CBd23MN9efQgCH
JrnQWzZnuz5nYEOtBdv1UYBIeumg0+7RCAPuvBGpnW7o4qJMOnYNes+hTVVQh9KN8Y/I6V6vJsuv
iKgw4QS5iCGA7DBMwqFtapCE4R8t9MpRX17x7jadosvcWc373df//nrB5uP6KgJDtztXh35gajt1
U2u2I++CdpnnuW7ZHwSEvhEBe7tAQ1Ad+vmfCIHjpAosJ9xwHY/9r+BPZvfM5F+Mt1QzTATrha4v
0Sjh8Ca28C+/hYMcMlycLI6mSf4PGhFunpDwWxkhITFXgla+2xjmbzrMUp2aeHWoy+qjT8vAzFGQ
iKBLFfqJaCYkP5nsBW7k9v3EqASHA5fhbxBH+MyYE580nsnl2yTC6GPeSiVCrLBsTp/HTm4bXhio
CP05RRbGPKEQRq9yRoF011uS92R9OIyHZAWKi3sBEXn0KUI79c67vH+A7abfouYsYJxgo6GVS1NE
qw1tZs9IEdcjUz8/uXpLfvWi9IsngrXIsb68LMTYlhy1moXB7BEUGZhaZywcpjTH4WeUajAEKuKn
gqzp9NxNvPreoX+ZUhOvn6sDQGr+vgEsLGZ3c9b3+st8NAs0ZQlb+nOqSFjoA6ByjVny3jp3PuFb
Rnug6/vQYbhE7Lezkr5ccwVZ9c8PueaSUV9WatuXAwR3bURJReA2pcqngp3oVtvAbRj2+DuqN4q+
IGLRN+4+hWznkVGdd+r3ggrLp52r4Nog2JOV2YwT3eoA+E32ld3ZorBZImDZMAecK3VHU8Z+5VWT
Tzs9vC/HNq3d1bmlmjqfnx/56hp1NKQYWxFRuqby2dQUeesY5ngZSiJBe9t21YPSMJKi/EMly3dZ
6VkR7UjVQq7QYIhTKUFHbTFf8XeGdWiZEfEj7wenIm8hrg2x8nI29TqdAOx+UE6oH8xHfcgibxPZ
EqcOqYcWMbW2kOhd3ezWIeumoOKZMniFchZgSBHBSFvOf0Xnvk/7LYG6r/IEgVypKLePpYqRc/PJ
i1FtH6ElLfsC/IA6KD+F6E2n5IE1gfdKPijiAhgvqRqAUjsQlQ2Q7qL94VQnYojkUfwyh/WtTkDU
1mQ3uMfv4cVCedNQw67xUkm2j8TyTxZRLFZcBoaDABi7ezxzlps+63U5+euiK81l9CHjt+lWl1fn
Or/nVyOiJRwYkoyp1E99Q2vhgSQb6eAgH/CLpNed0AQyZbGmYyULrglmcPRWKiL6D5n7JdDZEAK6
M8RLgieCZ/OgC7kK0s7eojqe33WH0VrAwAlatN88gM4WyW/93S4qzHquCi5wP/Ez76Bf0BLZbV3q
IbkZGaESA7/j7Y+etrhTod9/dAcfIpO5oxw1Ughd/G62RNq+ijyQABqK96Kq0QO02SfHQEl5l1lD
zA6jVPALVlKDHlarDNiBjOOp6HVrduLXiEG8iw/PytMwyEWmYhCAr0zBDHWN2Z/EC3LQeFkK7IvD
GlVWQqAAauRNGhSmAdbqC8i0++J1DD9ChvKXAP4ZWbHncw244CpkNPy/G7vwFq5XHvoTlTV1avnT
rFMU/yBDtsDCu0rxpIXo3IsuPXO4fsn7C3SlvH5QDw7SXwAO/fzYPQ1+EeCHuqWGXIC3AlVLyqcN
3osUZhJIIy/Ec5w9RLNE6K9g/N+WEfFBCJ/ge8/vPRHf6TPJjf+VgaXVQHemJ7yoHMLcMd/fJtTA
DerkEx9yzK1sGL8Pm6Dzi5rErEUdhesCwc40gq+liofZtrz3sVuRv9cUdMk/p/YT4ffn9Doi0CQI
zP+AXis9dkmdQ6Tq1fhijMbGN13VTF6UyP2hk85ypNlZD9BxTlOSYGovk3jqmEadJ8ZKV9Y62/O4
aUIyaiA5U4eQL6maKkZQtTZaZeVi6qXRzucQ5vnaBfg1aOsmjV+28oDAKDRfusb7wxHqQf5DjMQU
r9NEAFL3WBOwiAOMbfXLKntr8WlK4ZirB00ITWVdZ6zqn+/dR+w/GIe6BPSEf68I2XecQcul57cI
HnZmWLjYKOqMk9d444y+gi+3nFueaZMdS9e/Ds2O9Wzm3dyc51eiKr83io3u6D3Jp/3oHJ0ww6oM
IPbIZtUC0KspuXjrj6qxhWThBKNGDyuaBzvnV9gAISvev3AgZODRthdbLcYvLEGodRwybBNSxZ9e
SGfWeVCZIom3QoLgujWm9WU1zym/Nx6F0HE+WwWFEAnln2ApkqT7kpzeNxmDSy+rRCgtWspNq1t7
mZj8wb+Uj9zg8+pW/Smwx4f+WP98IBcgEszEdH3UC5EJr4RreFHRIs9o5ZxR7EQZnUwN0QviHTT3
1fKGT3xZnMLxVEM1TxbN/pm9dvYKvfLCKbKhP9SHfavnm+pexILcD5XAv5ZIF8m5aQaMBV5uRLrL
NvRIeAcIiZPw8v5TtJSPKpMPdR7tOFmWQQWnt/W01paVPW7XSDMWYeAjCDMwQBEXeY07q/tJPe1z
5cEKHHGwjgHb5y+EJT2jZcT79D3wCRNpWQIhabwIH1K4ZsjjVfJ1dw95n8hWSro/QyzndsiOUUR0
lp7bia+7eNO4Y6uB0W2cUgNZEWAxxmYEMKd/PLxuXsCvQyE92q6isYkQo5lNYwcvJsA1dPQ3L3FT
Sq43JxPA5y5GWaUMsGXUFfnGTsilv8ra4s85UcNfBVKf1TmXKjgr7dGbtePeKvAVC6D7PFtGR9J8
nQfgcQvv0uEhu23WBTOBhLEYgZNHTRqawoJpOnCHxiH1n7rEL/mfgsFK8E2H7LWjlRTFgppesMGL
LEP+XZ6GC3nxNkbLuwyYDcfoRlbMKCRPPv4rFqI36TKMWyD/1sWdYquaeq5bPIXzSnwF9dzlnN3t
sugn7mH9OJgH0/Mn/S5LCDyqTtN9uMpB9hspi47nVpHWxGw+3NtK9fGb6xa3SG6qfObmpzxYVEE1
GNy1Vefos8thsd2GYOt1aI+zy5he2ux+ZZCtfcTU+yZrTHM3sslbw4PNWdwBfsGyeBKqGr6gpF+p
BzV2eXrcwovKhUWGEMyoAANQyu75k5JnBodT507ChBFBAIKqXHxHmvowi9AKfrJcZ6sWeBmsmZJU
EbZT9fKeUtvqp9hczgp0WnMntf3e5YFD+5HJ6uSOW+v1CaLUW0NEAGFV5f1mCuIQ/WoVTWv37TF5
N8/YkcujYZfPn8SLlzdqiVzk5BHTpWIQJtn0jUW8Xl6k9cQzE1fLmArouCKkrCEXOxquypAmYY9s
JXmEFFt/vtON6mZXToJXIV2SxSgPxS+V+29I+ABADX+UqlzXa9vA3fq/0PYeQODTPbjV5XYC8waX
GQs5PQZWi9VEUB3WOgeWcW5Xlht3nFNtpTpa0MEFylfxps7l3GljeMe0uMcFDT4Q860yY1t8Yzjb
E2xFmslJOoWmdzvEI+KQCtlBYmlN+l2PYuuzDNjMIq5+mPM7YzoRCDPPK+iHPjSuBilVHPlyLi+K
EC/JvicSXsuMtI9pmOY6gw2jZnNb9Huchr8gp0Qbxgk1eyHHFWBhq58CiONMwOqp7qq1bRPigZFL
qqP+EO8s0qb0NSzLAHhWZDjgKbDsD/ffpNovQcimx0w6K3lkPg9oDz2OKhEtcTo/F8VTgQLxACys
O2do9fkuEpYjDZaZFb5ejrqNhqfulc0iqkt32oVTHTimvOspxwOfJDXvpN/T4oZEtXGiSHWjTvSS
viuJiZ3HdsU+WtSaJ0nJOGzl650eJwW232BpbZmdXE7HmPcGSUrFMnPD4L5c9QgiqJTXT2c9SHdv
XEWhMnLQmDXSHrJmdFffKbazbOe6p5rgTGy2dKE0Qu3zEEVgTa25r/0yPDa3YXv1c1XM97klm8MI
bMhyb8RiNYUb5f7zkBLbkEom+SeS89OvAIhvz3DTj+g9R42q+QHXGbCh1jUhYmWkT4j9czDznILt
khObzFKKIBhvK4k/U+L16gJBHv5viI22Q1PEPE7r4BPFpud9vtZnTb0Nzawl5yTnLsgzZ6MWv1nW
MfS1x5pB+het4VJIze/HI4q1cb6np2jEbl0EVaLYATPRJPNQfJ+kaajkIAlieTDIrPKa/OdocSPO
eY+sCkp7h8M8bYIpABbNrQPqHwMmwT/NGiAqn7R7Un9aNU5dGAWdGxCsDqLnk+szoHivTYDSGyg6
qeaI1n/8d158BU/Q99h/J/OL9UXMDJ7ZIDedf8YKdvQV1YzXK7LppVp0a14sHPRaR92fgRSG8+A8
KiO/I4lbYqImJLbEP5whdQBxO02vpvZc3/vnHccNnGWXXgiZw+n8cp6C1nMUL09qTNqg2yQc/RHq
D8MR6121/WI73Q6JE2TnqxSNS/bKI6z+kZpvafx4N9WgqDVbqFg9Vo4gHS3gu03GBX9wOU3PZxai
ucB1Jz6ClX60QfY5uFoXzYww4rNW57LBl5qDGQFYXo44UETMsJKvqGpy+etyDaLETWhypvTEuMUE
SPPVOePmfyf+zWFU/R6i7fB3zKwIYnrt+HiSsrqdQjq4HQN085CxjogGFDMxLMyF5EQSPD+bjDzs
0TO6ZkqoZ0+XvwTOueKjb8NYN9F11HoU8ZJ7zWsNaEstM5zFv7MIMfBs5cJJtBrjittx/RFjAHhP
YoGhoA5LeW4amhHYiyNKj+Cr/Mbv5hyj6DQCbe9jIBe5kJt1nY4wyuMZYVdSDFoWDydVmbA1bxI5
DwUjA/o3FEUeFMdSZknETx1Mewh1ahaa2gX4j1C9N3FCc+Oe7tmo2Eds2A0Bdga3Cviv+WLSKBzo
neNJ0osJ9GKUkZqSut14KvWbSla4KElvhhnO+QFgNrtIbAGriwyBlGj1eO+fEqHzxhZX6HeXUJqA
U0bM5WAku6KE9LZWC0H6L+npQ6wU31Uiy4QMVCK3gCES+5sBbAn/f8YaN7B29xb2LHr0qNXpMwRM
neJH0h4p7j6BGnxABhD6eeu51qrZ4OIAD6zw1qsqrBkVv4hZN0tIRaGwthFQQa24fHimCrhnLr7n
GQ7W1jiiKXqhEBF+XoIkWRw2hFnmOJzO45VC6sXoq9r+dt4oiY3pvjEm/n0TGLGQGBfWJaRqtHcF
6HaAy8NjxUz8S1Q2aqVtR/viD1bbtA8i4yxnZaNlkbdnuKa+jlE9EPZhQ6Bgao9IN7P85ffBueBy
axDUws4wshZMLX9Ka6GS1ajxrnuGJbw9W4ZC12lweoeNpdbC/8CxmbP4f5aPI8tAyLxhuynS/A8T
VFhcGvUcC1puJC29euXjeyZ6fMIZqtWkZ1e8TfDy/eIJkl7gftH685M2Ta/fD3db670TwKfEWxbz
iydhFwofpcQroUJosGUpMnQOh1GkUA7OQBKEdQlWhikJOSrEtaA2SnzyZbyxREqbP3Ucz24BacLE
jO2JcJiRhwnJvZhJo3oP9t2cHYAEl2Qu3D9PcP/2txXYTddaOauDoC3koWpuP/PxgaCPLBEo4Mut
+5rSkc2eXaqukwxmPScwdylXz6RvkaMvdmBe9GaghX7APZicVx5R/9Lr/+aOsqSZE9P18WxHQiRA
PD3bGJXC1XAD8YF9jBlPO9FVvBLRiUphPM5tDBvgb8ilfNRlpdRhkOv0IgPQGiCocIzbxaUaLIwg
0M8tYkLqq3UN0SpVcK9POpG5JusAfYvKNkvSFB7BrWU7tyoA1l7bB6U9IPLpPrhXJ5e3vbu0rpSQ
OBRItT9pejVBqn+caucF5FtP6/bYT8mDdcCzgc1LVEcNSeweg3ma0vQkbY1s/BSrEftjkpRKkn4/
dvP0DJF0PvHh5mlFvfy9AgAOr4+CM28lL5NuHSrfBgYWHnZ6Nx9alQoJTjxzsZ/XPeHDAENZNrAf
67rlYHf4eUsKW9mjZgNrJGJr4trcnycvbgpw1d3tAhlatJT8NAcTY9+lc1+lHkkch4PjjaUOuk09
COMst8pNImf2oh/sUVomhtw2ajCOiveE8nGKwptDGSXqq9Ep0MbRMA3igQ7ci/JdSvEhmBL/h8ev
+jXZvqrNgXjzADTtQn5I5mHiC/OqofPVqdPBd+4T+2VPh2hUx3LRD0bjs3A/t0/Ds3fkcaT9Zmil
p0gq0GUgeNON8ZNjwM4lTPhP4oKyjfeRF8wMqyXITZbRCIuv5HunhXjC27vSaBwxZOQGJa0GWfqT
gptHJli6vwWEW/0piiqx6fKIFbh+D9qbzUGyhfJYN1TsrHmT5aIpKP32UjwIy+ZAVcK31shNrYWp
+loCkzIPTkJfSPtR7rpwXtiJvf8+C9zU4BX+N/BAOqIxO7O30uQFQ4Yxv93XP9z44H1tEeC5zjWW
aUxKaQX33aA9m9jc8KsDmzOmrMf2ODDjQLwhV2k/X6i5QVj2//sYvcIOgCRqOHfWf+vFAdtQy1F/
NXnbBWVoI+IGI+aqNhYmCGGsoJKrCL4qY8SMaiLCRbU+9KeXGFO+CTaNsw+GL5Xv9cnszcfBiQZb
EbC2RsDO5ip3e3KW5m0jzVtlxe9FELkXcB8o9G9vNce5JxY/tQBsX371ZIvnIXhnXaDn1LZytirt
vOC9FYFJ7DnYbPy5JEANeZ2ezQIS1L0jGddBwyOnrQMGtr0wIsypRq/gMgt1nxcO9L+RN1k47gSh
uLArwJYykpu9XqFVWgJqrNpw9c7sz41MkoCnUW4HFHGApKVmOlIOv1xz2un9d+Rj3997Qh7rv0P4
YgPdRqE9VkGDHxgwHsNrWfywqZiInK7Efq7213gjfGHkuYVyUfgCXGLOFjRJit7UtBZkJQ49kDMG
zU8VnAD6XRBkk9R60Y3Bp6pRyA5BUq0B6piYBH/5y0u3Y8/W4s3aMQ0dY182cv5V4ADv7crOR5Mf
CZIzz5I/5fUwMUrgQZVjr5Rh32y8v0qESlU4gn/se3nW5N3iDMxXFhmqcKMetQOx3pC6sdl593np
bQr/+7V5PWlYkaQE0vFYiBxTXcUpZtUAKv1buRV+c24B/sM2H+3Z9EWM5dUP4nPEn/g2zQkzPoth
3k4VItVjy+isW81rbAFd3KWvrYuVlxuFEDsZz8QyNEbxBf5bVtff+lh2y2dtdm2d51VUnyol0ykr
36gh0wR90NUiQ719sjHu2vPEeVCi4BDcA0ESG+VLfU6ibuprKASN4vUYX/wEwqucT+1grN+wuLHs
CCvdpgMWFsonwVbekQGBdCvgyCcNiv9Q1i8rWZY0SmSOrZn6RI+mJVBGULUResC/5JxVLdwhsevO
TP1UHMJ+8joii+GW+EsMFtJgVroc+MFeomos7faF/O6T/wN+v12SFag+4yLlmKz2yLqez1nMWSI/
yW51p6OOqCusKcoAZOi0hBgHvkjoBU8+ewPxZPtb2Kw62eh15vkQrLuigKiRu/Iz4GNwgae64ceD
H9dGq3eh8StJ8AikmOdHENFfUoR9kBjNyVJc+3tDSOcMwuqVaAtDphDDmjieL3m0TMlCRDj74iBC
sCBS+PgauhDB8Mc/TIFzdYHQ1HFzW+i/bKWfHmqIwTq3PC5snEGXxnFUSU71c7LwTN1wltGH3Lfg
LOBeQyiqA2LFODwJ7b//axABM4+V4939UzVIxgFhiySp6+PtwDbIg/Ft6JiYlaW19/h8u/dXCntF
DTjsIFpGz7yFYXi03MudRKQlzUxGyplS1BjcuUyA/LojWOT2gW50pKSYPcexj4DMV8ljJcicI2Pp
C4tfdrVBhzHwayXHEEShY78Iu2sChRNfCKR8/cQGy8rZ1aFNftPs89jSFjwUPE3/7ZjVKL5U33zl
x4wtr812pQsSTI6KDA9c+UdbzAPuYkzTVrDIhQcWTO7W2/0T22M9l614b96FgBczZeBC3hLaQ39E
nAUcRWKd3Tin0xEsK4F1OWurDjS/9TUe5gOZshfDTMkmPKsBbRph8IhxYu8fFJVoiHxqdntIfvud
eUtvZr8XWMQgxzZeGTozC1mChLTHAomLv0QMwbSz0V6vLJdDiWfyME/Dzsm6U9L1ow7r9cymRY0I
XEKACt8Xl6df6fc++vyKGBVXCaXgHW5NWikE5XcjaDmoLcSiMqi20XOqfc4t2Jb5rQOBmr5AYTEF
oPKn0PoFw7p1zbhnMubmEguo/p7JmT5cFld5vGAVa6iW8wO+wvoEtlDybam8Pe8IB8OK/Fr6B3aR
+Y7EHkWoJofNAymJpnRS7p8VqCx5FyPE13vw3J7VHAUPH2Ktq0oPt7HFFTplLZIojnCQzTdP9BDP
wxJly32UNp40NYRsjDPNlfBQ3CLgCiz5xifeIS3MdOElIwNKvg4PJ602u/tAuCulFGd7lTWoujIz
vNveGDcDqje6M9LKiW2o35+ayXcFTZUiTw88cNtYBNcQGpsYRE2afWvKF/peaQFuENdSQxSV3Eev
/AYTvsQk/EmD2vVBt63mqQOqzr4IbcwD6lYr0AvSjjSAjJTuAjgKGX5+7N1WELQFhDLJfNiOvVHS
HuD+eipSyQddSCOfHyCXpfcnnpoxrmgPXne+VDL1pH9ung5dZ415/OX/foMJfhDTFomB+mH3aJPy
gCFza6D4WumdQ9KPRiN49kzZDWAdZW2GWBkZawB8kWvD0ub1Xo8K23x4Nm8hQvAk79rIvUxq4vs+
DtAs7b9tvcl6g7McxFgHXUBXHJkAFE0mWae6tMCR5SoQrh1vSiQsaIfRu+TM9nk00hlOEzIYhMD0
SR0SlSssP2tRnBNbUmhwmRU1pIXISgOwlws2aBUjK54jOv7Bnic7ht3c2mUT3x5G83GmZtZD4jel
QVGTkCreXJs7CvajM4ZCucHRzgAkn4Xya2T5OusLTaIA2yjUMoP701tGoPo8S3x9jnp95VH6rU2A
3mIiDNBR8eZUEK07gjGGDpyG2xklyOgCrPHmxkwXZAzFZUkqV1/bHtYS8hEsDhzxNkGaTOTHXIl+
ruEzCotOGn6KULk4017UPhVjZGgFzEfPsQF9GSplwcR9Sy9i+WV+gbvr+BgIQV0xgmX+cDqqGY/G
73O9BoUiyRNn9stdgNxPxNsGIXbM0w3jfQzmpH+rxiLCHI6YF9jMETNXZTgCjojv2QRdDZ3I4ZcD
F1hH4H7hjh+0smNt/AgYsNpEPZRjV0kUxItgN3wzLojGgZTddYHw1w+8nsFlp8H4Wrw2YGRFNAl8
5K5M9iNjwS4/h5f9v5BWJrQVZ+jYq1NyMy12t4dZu96bME/5zYJN18SS50OWbefjk7J2pFhQH504
PcsGY1fukjY7m3vMwsEv7rnxAcDcqgJmgdrZAGFdIRZd0mpmbBjjKvFotpDNI0MrRN2TBAVJvpRx
cLXejGMnMnRU8+nGvQZd3rbFD4tfU6nqnuzN+x1Id8v8IbzXsbIonw5l4/7C1grnQkSEVRj+BUgG
AnNnxGXYr1bzEzMZw85VsneGC0NkB+uLy6feoJ07TQHWuSh1ysKPa5nIBqcSMtd/1xk2EVD2C9vc
7UiuCdt+wfajPOF0RELx/SlWLI4wJb9HhVrugudSrnSmzx6+BaouR7Iqp5tUrG6P0Hx3vlwFNtPW
Auo+BoNKJHz5MCfmizwnZ8JqjC5qt+noW6bIMBKFZ0c+2q/xc6KnQhhWDw+qpdyvcXyWJHE03X8f
mjlQW9tA0kPOs9HU0Lf8dpPCQNZghf/zC++o5yGYmEP0Sa3tEA8aw+AGU0heu8N6iGLPRY9E2Msy
sFuvDiZJfp4m5qjZULLF/Cs6Mmyf+yDa79x4Tgq58T/KrWtmVjaRK089Bzhwjd5u7UAcqievRcbq
58wk39FM8hVIlEgGYo6/A/+zDJbMfJ/vi6Ldkd9qIA9wuL/pI3UtdCy09kCYLQX42NH6aMpVcJ9f
DriLfiqq3Sqbb+tpaPA2WO5tTvnj+RiPwkY57ZYCcAORsMA5lFhMKt7j1wS1FHSuKM2UztAFwO0m
ZH8L7K6pB0bouztiR05y/KCYn7YobFrqTuSc+eYQ9obto3bN9zLCxMoFAlqrtbuNIEkHNFfpEaso
+wvLSb4MTikaTGur6ftWH+Frb2NLlVHmMhT9I9p+uVK5FeQUWd7xBa6YfnucQYGChXwaamCiuh7t
F1XSgKRI2xdkEvQII5vIQsGdtQaIcvvjCmN6nzENFKh6mW5Sx0KQeHCBSkNrDZV7BgmKJGLkZqZH
jsAEObJb+FjVjBm0MBYxherWucw4QHLegw4n7SpAbs+O0DDt17PtqtC8l8XaYZzS4iIKLOUP3OXH
BOq2myGwtRqwFX3EKHcXW9H1oeNY7wRd4zIM2RcvRbkZp8hzmi9yRZCJ/yqst1G+CN4ko1NMerXM
JtIO6jS8gxAlXV2Rz2r6j2JIXqBH5JWh7TpOlONsyBulhPjicodSLjP0swW2WAKuTD1agl0zSmNs
rm0gI0Z9r9KTanUWqQyOJVQE0SlOVZy4ZjIW3c+HPHDyjIX5Q465VwB6E8jipyDDmLGpAreW5rHb
vfGuXiO5uqQaLQynNRcfz/tBNqgKFXGgjl6nYL5ruS8C+B9Rf2C4FTyN+SbPADKtC4lCsU3Bv5Oe
anFacUp953LHJ97LEmRPGBW36xGF1Q1qAJdtuBzZjZP1a6JVqW2zFZoAw3QHmYF7EVIEr6I5TjtW
cUcF6kX/z1M7wmpOmO2bVU8xtw2l6i/5IhjJshqR0WMaNnziqgw8MepIJ5RNX9F6rSXYu0xxNUmo
eVszJlEbOJK/lf4VRw7wzt1f7Z9dv+lpS/b3XGKtlpP1O8eNtgCjTRRFHJP0Ngce4i7/JjFYst64
QZ1mxp1hNDj0OJNYzM2OJvokNPT96bmvujqownqsGFnuoHDhAJ2pTXA/oiLtFQFaWFuWph1Ks4/N
sl/9DrzfXSr/qH7nTsCAa2A73S4k6uv5/7At/aK6j4oZQjlSG4lINL5QVwi+YazZ1aNI9hA39/FH
fA8U8OHXCKYYurjhUlehY1mp3hU/oBs8ozniIpqUEvWz2m3/vuIy0sqIn4OC4xeHLyc6N4yBvePG
hbNq7xdA5oHuUb8YJDWTL7SezqsptA5Ckwj/zBlwX5ZE8n3JrbS9aHG7mC624YUtMGIwwib1zNgC
yj4q4YY5TZgSoCL9HJ1h+IsPErz7xcwPFTYW6cfZuzjbs5ibAKCs9/CEeXoJA54r5W7AezdCp6Ne
adi0UHrJiPdyOHJlY2oOQLcpvOPVC7bgxudf0D/3u8zq/ixhF/B8v+fTCHrpDI0IVYNFHS1nTg7I
P2NUuuaJ6xsPT7mJNxvAoxY19KjQ8RdzzclOVw5U7KE7LXBmKSCG4VPXOIT537z0J+urmBy4jc9y
t1PmRVH2DqYp+i/Sm4HFW4mAwfDl/UUxoZfHxlZxBwd7ywBW/J32MM7zgfpiE2emCrsA5lOZhtRl
L7sROx4vD4/S35XV6/bCruLRNiIt/z+3BMvW1kbiHBFqwVoIbIruzf5l98gdRzDwmsd1Q5PJRVCQ
p1koIiGLekZXEkOmqqOVb/EQPbv5nR6hor+ExqrFD7259eSQNx8gLQb7wuYJ9bvOtwUe3MDnNVos
QHJ79weiw+4weoOmfcpTv54yVPBToKj/MkuCMwbtd0IIzmm2X5JcbuqgacN3wjADUyyiVUwDQJcZ
98UZJ3Rdmpjvy//759YhINhZQjatgGPFF/GhThvtnnRhNRR0/kGFrHglt61AB3OK90xblWZo8DGz
jYV0SV8SdTdrFiAEhbROkrqa0RKaTUNrhfq/8ZMG8j//6uPiE6vvYm8t8brPkyWYWIC5SgWHFeM1
oCxelHeFS/0ol7Eieg9e4S9wjeYUhzvdYXuJ57mJKeCQU2Gu7ttCeaA42+SMWCvrfObta8S/WoC0
x1svfwdblFbZLwmzMPYWgoqOB5ZvZ9Tj3t5K+E6eK/+B3mca7ksdcle0u35jRAKH+v4ClWYRBePI
1K9p9pLkQfHXRD0Pf9zx7CskUu+qqBn5/N25dF+Kps3S35d7WzUPX5Y6d2vO22PKpZ9uzqm30tXq
KLh/izspe4bSO+kZUA3DVvZ+nc5dujhaiPgnSnJzksQxFAjIUwXR7NFVYXZJ2P86Zd24a5iZnGUK
jbgeEt6UATY5wgoPK2u/xCAEkSucDwnCgSvInPPEruDd/m7diKC2ALaP6Upbszu/8yyx+/zmuOJS
OBXW841TbfW8j5vpacqQsjv2/BwBuG5f3cP/etQhJw2gazc1U2eN/vyF6RzJ44gNagaibbNmPtPY
8k335E2Hn9/EICCObIFMUtS9SV4HGoMgKV5l+nsbfCaq/6QURmTBZA+DXPH1UEyiRSt4mrTowOH5
xRUbHt1aUQQlpXvN6CwW+FCgLpKVEaa+Jbd3mBfOQq1byKhJ7hWqLH9nQ1PzAkiZBCWq5t72xT2Z
SVyNKtu7JRVo0wuHd32/H+8CH3cM4IHWRHH8j135vZi2+vhfsJwQAr5clQuzF8lvziPJUHgXgDWT
wFVaN06UQlH6inWxnFTrgbQRkq8ts9ZtBdTdoR2JtPZr1ovmzNhW1R4FxUgUQZLuA+t7jx7MFUEX
KxY4euCeDDo33+ze/m07nU92j+WhjMDdM++/SzegP3v4+RPEEnmg1BuymJTyEWNpDRaj9X6YlN7o
hM+R5hj38JWy8m7AnOPbq/X2ADki0zApm6LVmy5BbNSpCzfwOFL7onKIrqVoThzXOed0Q/aKXCxT
UAYruo5TUFuejsEKJBqtrHxeE6hNmFyROiYDEVRRBrw33pj5RXXoF4mfRdfNVbyQmN/eoB8sYwrA
Dmi99jCwMEO1TH+5guATb2pQ29gNMJNBi5p2lvbFzbNrDwTSCJjh+KsVL/RIC8Hj7zDKUbJYMRFT
oj/OSaAP7VF0qoW0KCFQR6eCUT4/vwzkmPMudu6DSeMvEyS8or9F1c2xvKhBRwcgyDVwNxgu4Tf7
d7T2K+5NV631Qb0+HLzntppKs3LUS2Z/3AobQIVe1r7xrCMcfybiWsxJydVUifhxaHz+zKoYdc/B
EsOaaWOm2MvqR4j27pT0fkzYS6XwCbwGtxwzOV7rZ12ccs0Ft7jRGAWbRrbRLbuvA+mVHH0a8alD
dihE6g6nQeos1v7GMbcb0/ph5MH5KcTcRCwLH6CJswacu1f5B+RBopQ//s1SY6FrbyYI+w3JY2mu
w3binY46ISOqKNVCGN1y7+EXx1D2UCGStco5DM+at6Y6EBdQUXU2MIGnbHny+np0RyzvSTwSi3ZH
ywi8+EmP+voeSxN6cvnNJX707z+Tj6IaJycOm5u1jSrUJvicjTrl7QKO1Q0FjlQPu4rU7Agx4ojA
3sbqYyamBBeQ6dLijlY5qndefLkx3JPfqpGBoNt8NgAmsong4iSbYOiuTEOsGo3c2FkdWHms0jYz
Ta4pfa+k9yY2CjuW9MpSkAlKjNWYEnWJmX0OlSLsKBdnsazlMoW/KA9J+Yk/2MJxa/7PxqUcE4RC
zT0Y/14RP+1QonPgTfbg19G/SARYpWbaXxSw68sCSX80YVlZVP0m1oZrOzrBjHAhQM7OkGqXiyhn
ALCeCx04Spc51OrvDr4y7KwZ97wPFOIBTClBRMa0wAqLR6o6mGkDhllbD81R1ClpC3ZtVN1Ea/lj
OPdbwnPkJfsGOmg3yzZA75CiTjBs0/2I5XZ44/6Cu3No2ViSfhkEg/FGu40uP5lJwSLHFizu2+4L
MdvVrNlMLHC7BJC+mU4vkpkAAc6U4gmxg2RoebmcbttoUzHSntaYwqYpL4R/mrQDCDHR5TvMThKH
u/E3MwY3pvmEmnzPIZ3MwyhKI8vtmqfzXgqMPCh9LIzHJbNGMMN1IH4TO1fl4T7sKvhHohvZqQR+
/owWNKF/mxP+F+n243RKNllflGV1m+9VfiMhN9KGl9Khwv9X7Paq3kai8B+boLh3MVyU1DLnUo34
EQA6D6ZZjZ2e3OvTEm7DWJOAXinLI1Un/ya8WPyh7C0TEDKxYtxnWr0Tvi6kd7grmFLeY7SitH0O
nbE2spzmtuF1QWZnLFSV7V+zl9qvKk+MLlPZ6DoKlwrtbWKGFiIdu/3AANbwdo84I2sypozwBgPF
YyilglVBYttbuoFPXuCXbhDqa2V+JvvWOYg8t9ZDPSvLpjIBO1EICgO//Krq5SjkJWQGUQyTGKn0
oG2IfZyUTbAEH/97NR/6QDmPoLwlGYEIfpxdtns7Ja3EccYDmvrIJj5KtLO/3Cw6tVC35uD+6xRc
8kX8ul95PInRMb8t95r1AeeZyW1/7/g4qRKQ+pw0hMKiv8aTFcMLUTrC+2WS81soIJZemEX9zu2U
di3MUhn2N2uOzG0XZn3pGZKI31UlcedxflREO52PzvqPVPUs2yy4vYOv7We6kesEny2BcRZLZxpC
lrYCyCGpnFrGIvBulHYBQKUfT45xjAD7ujgKUG5WJarKiD7GTXo2sXerZm9l2KAfyWuTtplJM+6Y
offYsZblF5R7afvYCxSPQvif51j8DlJduu1dghrF5m5tkgi0UHWxEXC6paX2ovBXGa/pHKL8eNLp
hNRhNS7YEkpZm6+gFsO+okQEiUSRSisIoXxZ4uvDterktfp/AquhC+7i2lCg9PzJFQQCOXJOIZgZ
WQtA47gXNupx66fo5ZMPDjlNH7488I7cVoH2peP4/Lc8V7zsaIW2likBf5I+DVaYDWVD1edGd/tp
80UwhuQNwvr45aqtMU7Ar+7kK1KfnBTefPiK85m7WPUlhg/RWyLXEmksYit0v6TVbM8eI4HmBZmh
W/TH6RiSy6KbOXH+ags46PXfPo+SGvZHYq4Q7neliLbejd5Yopc4mS+oZCe9GW78x6BjBLL7a95z
ex2fXX7+s6XxKoGhqZ9sqtcR9xhHV0tNSx/yW6EZKXeKU2j0pXizhO8fEufPAUKG6UBu5CUVNt7P
VTMd3CqTWwCq7gqhkUoSIhv1MCNJNPAkI15Jc4i+QxOhqv3DULEY3G6683qUwCpaMM3IwE7aIxwB
wb5P2zzKJ6HSE+TLMsBG9OUoN0DPlY4LiezoHY6oJXmjXEJ84W9kq7nmHvas73tE7RVseWtGjlz7
gEDwIaA5NiJSAN58B9rouWQlymRws8WA+PjBDF4Kh70sjnhZluLYEPQmLq8nTHdDdDeY6GIwO0LH
05GE+rdjaE5n5gRDXiD4BAqhhY8HPkmjskcukOEe4gFy4ProoqckWuOW8iKP3IBdfWn8+U6R/bMV
ZPZTN6Icxye6Y7fBuyksRKGOgB+kqVzUoN/UaNdGFbNpvche9oDxbPahG1oFztD1KrQKXs74m7lo
GSoxLHmwQgbbtV2Mwfq2oMZ2IuoiMiPd70sFpLc2ZiKTJPF4L23c6mZARBYvJIEfmv+rutzSXm5P
xSeDeU8fNGCkMAXa652qm7oqGWdNu1zpgGi4r/SLYTwyM8+cY0GIE1ReuOUa2anlzF8vHcGn+TZS
EIPoZrh90KoOuWRElWkCVL9UoR5UWW1GZo54PIxXp4TVLpRsdKJYRULX+anjaO4hsCjkDD2mW54N
xVWZc1IPaGvy6qtEgjdN8tnG0cagdI/v/3ul9AYqT45Nm7DOSCbALiHM2zr9R6Y4Jdd1c1L9ZmSy
fv+AryVUTEEs6SoDw8qcUFSEroEw4T8Dv3gg2Of8zf1axZt5jBhp5frIs3oDxBPkgJcGJBYyLGTY
ELhHEuzs9XrGnp82ny2Rfq5ZjdUDnLz4hTRYX+m7WC1p5yTv6bFEtxbPMiI93Bv6v8WyWjGJyGo0
5FznMplq4RD31cJLzGK8Ejf5kFKDLuSXl1+7J5oKEbC6kOWJq5AW02E7wRinL76eHl2BZuPyohNL
lart9U1icujy9iNWKFXiBqUqGIKdUdchpQ6agBcEOa4M5JN3p03IIGwJ8xKGgRF2asRVgsdXycAU
u5RVg5mM6izY/ZBaSPTuEmsTQplwiQJAx2sqVjntwPOeFzXvbvdDwKLEdR9EcrgOA9a8e2yuRWbS
fXUqLnW5jfVErWwOrOJxjTcJNLddwB+Q2BYGskUQGFuKIQGb8+MEW12MNKTnnRjc8nYFqFzJlWmo
PLcRAFZJdCVdaMHr0GMIyDh9dcAxb03yPfGqfhQmSXKTOq/hI3gi5xD8fZ+gHZPLmCp1a0FviAKm
HMTmUPQWeiDOBGsehmvNfLvLpYpPYLdDiL3mgRndQhC+IxWaTZfG35d48jMfBCU2zC59rKW88Djp
VXxHzKbF4ZJftTl9FM7YS6vBouwSwrtbveGtbaQ7a6iaqchLpbQLLpAckCxIpw+6CB3/2r9TxWbp
dcqefAbYBUhYzXMYlYE9/DeWNxJdGNTEVkVurU8HIXg69Fp+roBl3F72nYi2/IHrN0feh/q9A233
zrPaRh/j2I+wM9m4cJALSKXsbyYUWhDcVShWbAb1PEcLUGMk9pXpFMTCVTqulesiYfrajjYegUCx
W2jLEAekBPYYH4C0ZUqeXWZqwllZhu2xRFMW669UgqM1mFGn/3JOmN5rME6nfbTkq4+vk2f4pbRH
jwI2ERh5xYtUL2sH2A/kNuI7tQ8K+uMgE7lFFbBc7Cm9hZHLD2hUgB7eSqtNhap5b5w1w9OQKR3j
f1NxWWM/OgDarmtEeS6ygLBBXsaDMoTFKSqryxIsNlPZsN7I1Ah7fmgOU2qabsbYxl8jlGVc+nAR
0bpFbdtUnIqje/bh7SJLMb3SVfzYzFoIfotbsgePgLlzDQq8bjBKAGLc0rFeK3Nv4Jkap+qP8EnX
FILUm2An4Wrto4YlmmjD7AjU+TB3dpjP846Ee2BMVs9F0p1rGczAVkQVxbKExtzdYgarVMJ/tcmD
8lNAGXNPadCTKky7CSV1lCqM11kAIzSKfBpxAhPZ2VD3xg6Aouzmw5aw67/Q44mL1XO/UV9J0vbV
LOHITk7XQdEHIsYgHPRCCG5KId65hp3fw0UDm2RyMhvNcTA7/gIXqZtacIciaPUgU0UCAlc9wTJk
o6lOFKJEvovlkkHJKnBwzW2bEIjAKKwUIxAdIaXT/Qt3YniOfWpHel2dJvVt84Isxe63iMHrYTo0
dLdCsvknMeZPPJrfQTZfOcP8BXtZcGRP5wGwwmrIQ5XoEwyrn06FqIZMtpxDIJrWA5PpWyBpm8AX
9TlxfTPTZ/Wv0XZrwQGRNC18k8Eu7H9bnsMqExwQoWXYH1O/bYPuQ8PizJhy23NCuTI5x6zZ4EXS
2WILnms7rcROwGQlHMq5zdH7r0ru0snpLdgQUUFtGemBhMmlv73x0gs+muzANDd/yRfRWjxnhjPP
cnDB1f7yxn8mxt6sJ4S0XShKbiGtjw5y5pDGuIfgIHXSioqQsH8xWmihfhX76V9n2Hfl4S9FLUBv
W+diTWedfzVH3Nv8fsCbQO90Ofgt8VTxO6DHMxYJbH7S0mAHA2TQkuzT0dZvT/AJRJ7NLNfHiGuq
9Uy9X8jD5Snn5XVkwWM3sexA+1aTgF+7hQO/OcCQBM2gccFyqxzEvOZ3RwWDoY3T5MnkbRwMHTyU
UXhlrq2WCqQpmbT3s+82KyixpP5oLcI5jeGGG7MNCCxkVBMfQkUSpd+LB7BoFVd69XiiBYy/hqLq
u2Ssl0T4TJuNFBLg/LmxwU95EthSgbpqRv7I9fMHdJppwUCbuLXaFPx1bX4f4Nnse+cYwwpi0N/5
p9MHZ+hJ/1aiEQzCiYNNCITKjx0KR5EhUmKLnF7Ma8DAhoQSbMgbYkzuMIunMvxfhJbn/Tf8INXB
jAJqCPaqiaoIL1znfZJP2+AQ7fcAUCd12O4jD6dlNZ3/HJbXRvhBLUr5hIfmKJWPZqdob2NfxoAK
UK3rgmNnOPzbTV3ju8PC8SNlT9wj0/AZuLPUarm2XLlEgZngLlu+N/6zJRHtbZK8CmPzfm3Gibc2
d8ETpXEZwo6iCvLFS1g7fbGJzqbmP1PISOsndO72tSZWHJ7NiFpZ7FiQyu6KS3R9449jzyHg6nAB
YhpklPoySbXTMatHgiWztneI6opJSC1UlD+C9qjkD9FC2/uhTdmEtd2HnUhe2Nr5HTiYGm7EV6II
PlOnJ+yJ7AFTfnv4G08Y0DZ7pR8EyJ4Doef/vaNuVpADsCq5+lUqsghODTrPCwjnzEd9udXiqgbm
R0jGA3BQn0AirPaPyJMhiILdFL6WmQmaOegIix6roHXy1bSM2SCxSl6TW43bF0W2/IJxmztW0AHz
7PsFb7zxvQuiRZGPkLSLcXyfitHGx3+R7syIRHiCm7Hp1V8TFlkiS2jlRNORUf5G329PncJfDxaw
v4u99l4uNXH1DK6jFAtgFn3LJLoCdlTCG6Kd+yF8CaFv982D/eayUuidrhuBdudI0vj1diqmo0Uy
bnGCM+EXrVloGzz1yXRBj/HCyqSB17wH4BfXq703aeNqoZqB/+MZu1DFJYZ16kyTmAWhHuVzrIUI
sx4nLlIavp3qaIPJI+p9P5t3FoXcmwasNSLe7vw/fTU/c6uxs9zEoEvOVtWqZFWcqM1qkBTND+Qr
IRJE4iWed1q8xiNAEoZr7rdNRHeRn09ZAhRj5rMmBXcBPd4Mc8nRknboxZ405Fr7SMiEW57kU9KS
UXSTh7aJSyLb5bQ/tTNpAW8HzIEjY+T9+6ACBPmLC4O9XmIKcmAYA6+6M/yuzjdOiiuYyMCBPy1r
3ZJ1feoT7+zmZ/8dpAll4H9lkKfiTIFesDm53OwfkHcR521oJuPLaLkWVhMqvhBg6C1VKiKlJ5IC
iXqavRI9/2t3tiF7ded0DWGF1SwEymy9ygI4Jt6nvywMLRUYYRt8jwcmWFNReXQL3We8NGeTBkcW
Pa2dHBxHe2iv2rFPwf+k4aoHpnroJy9EKoDI1T7nVRjbApD/XJ4eKOwWwKHwwcJUGScXdIxypg8K
6QUFox/k7L1dumABea3KhWOHNGs367z3qVGtDq6UXj4TS82O7oCPUqOhVANsksSPolbZ15iXGPdo
GBPYRZxVF/r3Ol06PtTM077sIxFUj8jk3wP6cDyR6NCK+jIXOKi6iDO/V7B6dKHuDuB0xvPGDDkR
q8xrlXnRrs1stCIEc89Kfl3YeAJgBF0e1WudvbaIoRWJ8LtAXydkl59wR9FWL+7tFqYORkf3TtbP
GCAT8gV1uM4HIAhPDmRTdL7BitJf5nQwFVYJqhr2vb/gWJnjFCfTYfI1288mfBBHGH+pB48BJduH
JjJHPLJMBlDXEq2GYpEBE6LWuRohQ/BlPCH5hj8Zk5EO3RETvM+zYMnnnU5kCIVilx8Ww66AyeZa
Qwka1MJ1Z+tuzVZbVibNhBCj2M95C0CgeuIY7198tW4t4cRJ0EzQPxoQXt+yldOmQ0eyAumUzF3g
Zw8/mc1/Ub9si5tw5+UMl2zrhJ6XpxHN72ROoHA6CoQQLJXi9gPdItGR4mb4qDtoQAiKG2IrJBe9
a8A51OIiNoMnNnELcBkDJ3h3wgb3OhNcDMZVQiOHmprI/n6b5VVVfWVHy1onlassvos4dgOQLUkQ
AqjyQw/B4zp/EQgPC2jIwqIAMerRidKbLQH7qOQXLxsbeArZT90sWCMWKUMBmRXRbopAHAJ1iNI2
B3wBfkCOifQcr0oimyLB7TjMjxFO0TfncMjWD4MR/ywgEeqFhQa0HVq5c+2iEFjrvZejsyATYJup
zUYddFxKyWeNsGpjrKMIt/HvnEnyFeb+zoOEIG8tlF98GO4w+oaJtXKYW8H8IJixmTWt7OviILZ7
Uw3hi62m08Z//ulfDAQgMhbFTXWhw8XZboXCVxgfykdag60iaVwDy4KLjPblQzLDSd1wshEdQxos
sI57Le+MkT7D17x08AGtv7mAbdmqv0q2he7u1VxlXmgsZemlIBLOuxxuNP6nIeKh1Lary1GXqBv4
zkwlPcnvo+u/IRLlAbYU6XO7K2BlssLc84ncj1xLPXrPSEUqHilO8RnFuo9xtrPYsu4+yEk8aWkV
2YUZtjVAmDfyxp9+P0L3SX3P4W0iAzpwuOXbu60UUtiU4NnHzH297oaSPQGcJ9tM6BnlIsn5GA5v
mpkrdnoVVR510USOXwl5Kc8BPP5CHAEI9i37eP6LFjfSmG9dX0JOHj0XXACXOc6w3nsXjNLPsoIo
mIWcRk8AMB5r5LCuv6fSXU3XALS2x+ngIYUamkR9sMIYUhSWUJqndZ349plx4YFPal1AOIhWZG8y
SptSlMUInc/JU88MAO+y/nH7CFax+utsHGyCq1frrFxzuPYhCR7JaUPs/1OaT8lTRzMjIv40/wnK
L7PM6FvNCEOoUuVexF3TWRgnajzY5zAUN/ImnbkL1kiKBGJAeQwhJrmWyeZek7qdS9kdlZIHQAj3
VAjrrZ33y2KE74+AhXO4sy2LWsunOVsobMGZh8SgkTwyC/Irv0fq/E+fL46yarudt9c++73476SX
BsqF7Ln3+0Vfgg4Xh2R7jdLw2+ZTm6haaI7a6dGybGePfQSyltzTB5Tyuq/alIjM1O0ZobSVw3bV
CYY//Z+CAmPbb7LtwIRi4bOyx+vJq1L+1fFPf1nLPax8ufqU1kkp10Ab+NMIua7Jyv+eQvpMCsH8
fZSDrpFRdeQuIH/w/AtGwCVO07bqqGQQria3W9KS9yeQKw8FxuotDE7aI6hz23v2pITWt/UaD1JM
l+KFWS8GSaSg0ARM6C31jga0Lrms3YSbe2Ae5RnnPQk2rTHhNsPHg0kNOM00PxA/IPfz5Z33cnEv
NUsAsAbqnMNU+QM4UUiSLa2BCUPDgn7hLhYeF17qFm0e+9lbHn6k2XvkMnlGypcf+Be2GcMe6R0B
o4jsYiM1kCgclJ/USrmVbkeiWH0+m3SwxGM4wBFc0DLkOI1Wa1h6KnV98DpINuVQ8x8UcxLMyc3/
GVKiz6HLnjed5D4bPCyh3WioQ5s2j75e+73QJgi/t4rN8rJchShFCETPwO5r1rU7GRMbyd2GmNsN
T1A0Mm+74AA6EBAzQpTKJg1gNjSTh0wXbt/dzmXd+SS8xX3r7v1qzFPWB649Ghg7MzoOzf9W8SLA
h3IMv5gmtCI11/OUAc7QqFHiFkiAjFV+VtlANv85Novb05Sz4OfauxE13GmUXz/v/r2m2ixfj8OT
SDuqLz/X6juDq77EO1Y/HIpXQh4pKOImHZX/VkKOP59tbI0DJjDHfR1ZrZ5RUJSNVm8ZGKQ8HI4W
ICkwsSJ+UchoNzz7h8Bs1gIO2hhgp29ftVnFU1uTJEWeJXa79SiAUqJjfeNiYN0TjyF74XBOwUi+
vrMt4NzpXcIZyTPR0wQzmD2A3iGiOBa0XveL5eJmEe7IBLu/utWsT7i6/LbRaiSOr2/0asu+Fb1M
uJQPXtzKzyDRDlEOlzmuUtP67SiyZmuryrO6XKxLIOIiCdGMmoQlOgZ/jF43YNKFq/jXtnMeZLbR
sTfaEm/T+53ChRI282fPR8K4on9R0vCXsA1+XLW5usDRBpBmu/JiHZrMm7bLRAo+xPhsbsiYNPhP
teYSqdnAQiBAC2oKMFmazuNXtLluYceyRS80AXVmDDQ/Nc5rTF2Ybxk5S+wh15395iLOLlkd0k3k
BL5SrWQFRSgQZnyXqnOHEwxbCxcTmrYFZpsYJwv+w/z4ENByFmBhwsbievD1MaiscOh/EWNZxkmY
B51jwvu6NE6pU5z/Q7FRKxXKjtodaSMGY5exGI8FnwG6HrvQfOR51sCbs0V1Iw7w1nLtJpD+FgF8
/vmDXYOoAa4au40CjMG6ARqEbhKqoUlGAB6XQxdEmQ5lrXmJdcR2jUwUj7vOY+kyK0+ryGZm9Cm6
MY+BGygXch7HYLzLv6xrrl3ad+Byv+Kkc18NnNM7x6AMQbvkWH2ebkvcTe160kiWfeLhHlVWtGAg
92dXX361Xdwen2D+rVmJRQS0lcrzaDlA/BsyJEtq1RFJqX6WmO155IwmpHZKNvHf0EK+OPqMtdD1
+z/t26nPafC4LTUY56kXvnDAQIrL70wLW0SgUDcGy4sn7dk0zQ6A1J4G7TJCpVZtvHwXtmFZXy2Y
Sa08G6/th99XjB39eSc+qNm1usJCFZQ84R/DFLzNO0ukLEfc7qcXOQjGC3tAGkjz8V+01dmcQdq1
hDaAvWszA/DRc1fT1N/WdKzpnqjEkbFLWX4qb4mi3EbOMIIgX01DbgOZ/Fgx3VHdtIgrOtGdchwv
I9zn8PEE1ejkouv6XD9VTX8TdOZqtXYqrauDH4guH7qtWnRZlPt/4eWzcU3X9bgR2+3ZcUUPtRSQ
XmtS+T/EXLr2wDcsE5Rqv83QWyxVBWOPVzbwyKlY8wCuFVWCcPkFWivszW0PubeEXIFGuNKqjOjf
3KZdXydqzgfY2gZ2CfPRSimGIde31PAmCJ9808E7EA32j45tu/AuHgt2PQpUbKhBLqGDInElvQPa
HxAYgZcICjUHVM0haiEJtnYcgqD87HRyRlvP2xsFcaK10vn6jvSd9pUs+cM3Ls6VcykIEh8P6IaK
cwFw7XrNE80Kgw2it3VPRtkltvlkvRzKrDIBOPbrN4UrY9eeMYKO8oFQ+XLK8zxMTLGqz2Sl+eFs
/0+Lc9gM9JBeRYnUZQTFhg/aDyOI7n84cr6ObJq/yhCK3ityX5WnlXe8eAA0U9QADhILjPfVFB1e
ZQ9+sqCbpbnxfi8JGRH24mogGBkVdUya0++rxXhDPp5cO4+cC6s2r3Jx5SBm6rLycA8Wk9zLtKAK
kKLFlusz4pWz7hgnt3huOI3pwdzQKkj8oofhYnDGVbfdbYdVX0xqq30Rw911+Eyjew6X4l7oX6Bk
MNAuTPyxdS5vNHxwMJIdBhxVFkjWVs4HSeNnLYdIRYXkaPDWDOn9eSnIiCPTm+X7cwU9zaF/OZyj
hOIFmdyqtm1fLBZO9oShtYA0qayhwz4qHj3DXym1xA4EWuotE4EFT2BTOAVXn5E9miFBEG3lL9Ls
8yqSRO+9yUgo86IP38QWO+tFQ3R99Sr5SCYeGQPVTvB6jKwixCBdlPRS6fM2TfIf9Y9YDM4oJEM8
Z393ld4fY51MYsCxb9RbDK6TQYIrvu9+uUVBS8mEBNjFVLuWNNoTmzKSeft3HcDVBvSZp5bHYpJj
aHlcnYQ79GIHrg7cxnxGz7CFZVpKGjrRHalwgaJdV6XetH5Vf1CPttypfYdVb7DVYevCvOqyosKw
y8NBG6WGN8lIT6RB/NzA6EZizgt6A7TDfyHZrZ4eY4uwVDFVucNWAF/Dnj8EyRUNo4Wr/2pZwifc
5+WmlrCRSWgrqVjb4i/BJnW0haFGAymLfZKoSz5HM7Xev2kDjAAGtVu5hohYXcO1jfj4Lm+lRXYg
kLW5SqX95K5tNRycs25HrkvMlVSow9xippXmIt00ZjyjmNg4a2ALEVnNNqGtNsqibxVW6H/LeDxE
0XVpbM9Ycx302U0MhUaKQjjjI36JUFUi6lOhFDR5TIqCwvIm3sRgu2DBEVUbrebK4v8ofe/324vR
EZ1bat/q3XieBf8YXePjvt2JiSBqxrMUkSgFcnL0pXyybHE5Knxo7jMrTYAjOAJi1JmVmTrMRZEw
5n/tdbVO0c26e3bYBgiORY1lVjhL/pWOm7i7erl2DcJlnsZDS0uPPlNqsNYp0dxmuh93M6Krc3gC
Pu2cOd2AoTb1H4I2HOZZk/xJ2UCR+hg6zndlx1O/izXkOoYPL8PVZYVdDpyAzMJyasyt3YdJMr25
jxQmnES70oqo0V4VOPVtXQPEWxsywo40XqUkxFc0Vchqy0NQzUEGpEx3alPzUcEcckPqg9xE0+Dr
39WXwdipKIJioMfJ+X67V8gi2BD/RB1j2tsxyRBwwjcFxQ0W6s6Uz9WT4xDplO9ywVZ7XLRfE8NB
6ADXJue4pzO2r0fM4vRJsfD4drIyN23FFkROgLMc1nocMZ5S28U/kp9Fm97pBWn2tBVvjOhYaa9u
vDp5lf/941lOenctQYEeLbdvktEz7fAQK5NmNgeF5s4J1S8wN7RevCqoBwq+Q0MEgPdtpiWf7OHs
SPZbjnmSsAshgc9g+7FqHPbjfACMNZTRMCSrQA+zprWt8fcKKCX6mMv9jqd58e4VqzmvlGVrXPQr
cnzKtsR0gOQOYzyX/xc8QMH3gFLosGIJr7b1AFOQVSa/dQbhZAj563OBL8uTzzQna+nF5h/+NHP+
e6fuMvBlQ23tBw1EcAgA1U6Z/I7OitAci2q26T/IKN6+RTWB8p1J+7zwRM+c6sLFONaCVxX90Ks2
cEB58VCYJG/0nXHel3t5Qosgio0+4p+y3nSuif8tyt1sWh3XaVe4jv0yhUmcxZhlmoJhv/kAMG1i
L0uK3DoPQqN8RojY+BV+b1tlYW/VULY9zUgGHf4hrA6W4LpRUn10w9YZENAj1VX79/FkKrYyIrQJ
dHJ5jlUV9Bizx/fztrt8gcbnjnpu0owyC0RAYscxH7moVNcpHfyOT8YBxd8tscAKOnAeUFxD8uUd
VckFjyOomMdTIeIfNVIU10+ItiuZwjU4GBd9nxs+rXD9jcXPVncpaQQgSI/+JcLPbwhsKe1ZHp7u
GBnRLVko1JofW4OaZRYcBYpo5F2B/MrvV8GPHivL8ZwY0LJZ1VaVg+HWgputzY0EkEeZo6mLs9lV
EQcI8/kfOL6Tm0Pg8quZapd+GNqUILZ/7e3fEUJkr7VzNzI6kzg39PUfFn653G8+LJzJ3+902zQM
caDaSIti/ycu3Wb1cOjcugriMQebdS7gvLmmN4C1VKeuPy7+0WsXbOaMNXwPsH/hzpap7KAHSQOv
1GvuUbtLNURdRGc1W3xoA2QSUW8iUlMihcwBa0iIXu0TFeFPKdsxnlKsfcY9i4tRzCdhtBg0numw
PCExBIVp1My3J+1+gJJc+Ks1agd2h3UYq+YSr5IvFuQUPj1XepCnDYULBlVRZgz1U+qcD6GjvuAj
RKI92YDImiR14uJw39fgqu/8KCPMl5+a4ofjsNG4siDWz2oXGtppCRV7cmz6QAlY8I015lgEk6BK
WV/1jshOFyMrtoZVm0Zqho39vdrR5VAO5pkXI/by0edE3twX2zMLBl7rc3RXKH5J/3rJGTx6kr8+
1HAvbIeYBox20v4bCxh6aC9FYsD6xK1VMlWzJrUSmutwuwUi15vqqp+RZtaB/I6Fpzc0l04YKYHH
1jaCFobQK3sxtT3whyuUIpPVK8xKqOXbrA55Gpn0w/YWZy3Gp+Nz29r1iEitFo2iNkkPUMFJENRA
5nSOeqDCcvNaTJLOWvlVHRD7N3tzfnYWpnZWZogFeqH4Iphon9uEf1T1D6pi0wyoDFpJMJoRoGZy
YdvsLPR6A3rYytEggItk5GAwClE/s4Qsb90YkDQ/hVg6qm7RoZXTSzmDjFErgTRG73UNTtfM0OTK
SIDdV2igahUB2LfPgLm4vRKlnxDfJqDAMCSyxUJbccPWWcJ6U6BzRiGgOKsAZCB5VMwx796yxi2G
u4ykE0VHDcTjiZx57hR37201UBV7xXqy5zhXoj8B5VpTZ92I6dC11vuPwSCSMajBifsphBX9ennM
yBFwwmAFnkrjapdDDjfvfr8qa4cpNkEGsWE8CnkQH2pbRW957ZJ1TEX4roeeyv621iuWzt46A0BW
PES9JanrN4kQXq3aIY0LlY5kslM3HtSooNRu3FD23Ofpu553cj74UnInvlZsxORu402I0eAVcsBi
GByfMFdk50scYYjXQrHAcXv9BgpZplrO5iltloWJm/YeKw4G7RaxUxd73A1CK0yAlv9L0v3O/dxp
sedvXX1N9y2N1l3kc4LZwdcHhmjz1RzVDL2gzIEDQWAD/q/CuueiSXELOoVG65CflmI84rYYL85S
GtyDV/txNHkN2/qqA4DdmI0Uh+Gq/LEOAIV9I16vc8xCDKyph0sXGovyB23k7L0rEj2po1cBa1vT
WtCn0zX6vIRtlsu8bB6L19EtbNgSm2WdfjXyTrz/2UDHSCEDUCHjWxxAgpeuV9bfgL2IYYC8F2fQ
Go/RZMq+DG5T/LLW7JABk4ra61+cEL1GBq/hESaFJ8JhP9xabWDUTuQ3eZjfD5A10D81bjr2QoVr
4zxs9aJ4MfCzNbN+y5LHA9CE5w6hq4svtb7fB1W35U5rXxFVrobcOqu0CuT/V8o1qlJ/dOyJKFsT
vESjAIn0pa9kCyaAMVXVmxcJzrkEp9Kva2OvNCvr4m5bjaV936QQ1TclAL2voAEMipCbvRC3qeHY
vpSULdSEzvv/f+h2PN/xm1V+46I3NAOnx0GfvfjqX/FbChQ0unPpx/PuG6z0j6sFLF/FzjXPdx3Y
DNEbKwov8HJZzN0+/YPeRWZvuyx86BbvEgHypyZAbEFn94WDspL+XTErNaI9alqifP+sMGl94xTh
SZA1uVD7s557nDhJZ8u+FiXZVobmIufGerpTa0Lt7FMRbnge4/8CELRKXWaFhUMmqmnm4j5UQ3GM
70Uss8k7/arjw/MwZGveUmJ9A8FqXCK9F0ABoOUUtIblHFmwwoW6wE1g5zRRP1pajaLiuC2TkXLw
bsYRfXMC07CR1B+G7t+Kdj1QCn/V6cYHDmFKoJXQNxVP3K4yBQeOdCnKIqE/hfFlrdoOy3YAg4bp
KAXon1SZD4W0HCGoaeY/GpcvYP3MqYlTMpzDWZkYT0CQuqIttknZ97ihugjCV7qjzcwQUYMFA37w
I/jpZ1pxZ3w4HjQT97/nkwFfnCcQ59aadCzy2c4lw9tLkDa/4CleQptebP9ZEmbMbM6bL8VqYN6R
HNBuj2wUpUpgsbdafVHa98AcxTGTWkD+wUgGf5t3eRp1BtAaELAoMth6ifLVnqAAUoszdhrjT/6E
KenXby2kco/CTeEZP3sLRdguQIMA52gXmndZl+5uWSLUhoGCPffsb1XV68d307vgY+jG0kQ077kh
d3Gb7PCfz2wcTy6xpgCwzBuED2/p60PGw9d6HaKBEGgn+GmtcJ/7NOyK1lXaGOkOPDtuWU8/pbHI
rLWx+GSTHicZXJnaJ9E5p6EtbMKH2HepFFMNTNjymB2i7wCkMA9sgMquZiBBFfcgqTXy9nsFx2W/
u+rwzDVaWzkH5J5AbN9CYe/fvRUoO5oewk0ABiTZoY8Uo9ACuPQO21BT994FD1eyu3PSzoQHqWA1
YYxBT3TvfFR9ux/bh3SpeZNzrz2oU5YnS0RfB+cqT5Mi7FyiYcFZ3fqfD6BgKRMk9WdfTUMgNZWX
KBxQ93xHkGbqQzYxI/GZJYNsBVlp7nnLCrijLATFJ8yYlf58vg0W/+fq3jlNW+XQexUCFH5H/TyH
VKgz8EVcwdHMwyPcWxGCG5CSefM2y9WJTvegYIMhYq2DuxxjHyqbVP5+l2GjlgROkF5M3NW4DuVE
xireeJsurJ1378ARupI7hSWtp5T+CM7EQw1AzQtZx0sLQtiobT2grWZsZR39ArLrEweKaJDWnwbE
GvXFqwzkEF01ghTqcB4LmboYJy2gQ8q9ywi/LqXvNTCtFQqEGfDUE682z+63LnzVFNXe9uGH2/ef
nY3xyw0P7dWus84+znMX5PoOE1dVScbDICnlUM0VcjWdIA+InnosAGuFDlfn4rszEBMRVuY785mZ
ZMkcZrRqI9avKU3eKdQ5Ui9zukhtpnnBfLTIC0FNteDJXeIcDFbPXyRD5hZi21SwjPZ20ld+8SxJ
Ar7SPG2SLtryOjc3TMzZmWxoET5zi9UO4wAep+ljUC5q1IMRpEnwL4okLbILFqg8CBZ3/ecTCSJy
dsOU6/mSabQKoLVpVPaRBpQgFoPS5ErdbJTiQNS0w88gVpYlg9woh4HSabhLBYZRhNuT8MVjkol3
Ni+wruWEnW0pCQwXghDtDXV9/KqIY336P0MMzBDfUdbtfzQ3MwMb9bYRP1NU56FOm+H7aVO/yQpx
8zn40edB5WK4vDa59Tv9OXTvBnWTpZq+ICH0LEPLd2Aeb+GIUvgnNBuudmJS/UyF4TuDPaC1TQ6r
nS44T7tK8GTJlap65KRHP6ODBKiRaMaz1TkJLjRT/I/uFzamfoVB+YoZpcdReZdFCDZbvOYN5tM6
thqBETTZ1LhGwxu6OWd3N7Cy4Dx06vGc9V3ZsaO/xwSfBkBcF7diOwp7rEd1oOpjXm1oI9tTkJjF
pmc1/jKhpGRKzsSMBdtzlLLOzzQfc/VkVc+aWYF4mHCXei04Ts4+HKazEPgdRYb298U8Jt0N8tyv
JNWrrc35NbWJDUyfuX4cVtAqwp1iNgWOPaCXuSQtW4rt+9z/Ujxdy7mh3Ix3eSTr/ZMZNxrOy7Se
c5itrftue3pdjaKQ3vvPBGAANEWMMPeOSH3lzuOvYqFVO5uUyL4nBQfdlgmycuU6wDiYOrcysnMO
QYIlusdiU/dRplmJ+cadAGnwfndGSwcBsc7txrQsB8U5YBFjtXF7YdOT6N0xuUt25iOKqqVKl+hf
iNehqcRQ9B+FfEyED/MdsK8hjQotfeoPuBz0jF+/lbMDcUZE9aiW+ECZGIWmQxs7ZqQ9N9/+vtpD
lqULuuYYMs2adWmHDCXBMxAGsS6wxQprX5goY3+k8saaDm9ymtNWa59oCyLsAsTut8bjm/VYdiBH
/aikgsLQ4QUQrnyCVgm7ufDkdWsvFmTvW4XPxVOHYpGy7UtPrlo1wdI6f+zZNPeuna4GkbnaE4kU
r0dWFUjiPYZW/ikt6bhAnLb5AZCpIG1FkpVMcvWUznE2iLq/gEmzTlgAreCEgqfADR5MgTxVx9AX
jGUVJs+zJymBvA9xcfR/dynJ9rdQYBhRP0WlmVAwWOv0Qad5zsSq5hmOmSCifLVY+a2Ecudvma2U
ySbKAujyP46R9Kl4tJSn4F1J9dzaeo/YFjQBFrhToVPFwqjJv7JESPv5CxX72WVj+HO8MJLJL9tj
ioPxc2g9sFn+2kW/oJ7pd2LZYeagE5uolWafjyUshiG9QEQWRnZj6k/9KTOnKu3pP4/rE9yhVgXT
3i2QVqZvoVVOwLH3eP9V68mZFzcpyM0TWwzICqVqM2bx9ezMKZ51VAZltxa/APyC2S5FS2H2TPaQ
nHoJLeT/vwxVOSwIai5iPF0GUNwr1Vn1hVsxza45ijv4w6p8mlOsBSQc6f0rLesgefaY8umT16n1
kHFEYGohK+aGgvim+Plmc9hm/UJZmj8MvnwHhFWLmvd7nJ5ByxcxXlZmwk0cDU7GMU9K7eF0ogSb
dZfFOP/Ma/mBwTrVIXgKBCgAGPvgL3zb40lWrFVwZYk+lox6VqP8Nxu6rbXggsihE+428/seIYoG
7F1eK/ywEHl+3KcFj53pFrdaiBsr1ZGgQnjXQsK7FvV1c5xyoBZZyE6XkOxE709OxT7le0p9WXcd
a1IendvVyrVh5TuqUmZSDei4z37+wTCmd8UoloXeh4HDwD9r0coMLBxk+Dq3gHqnHNZTUul5GFBs
b4ijyDYxBSzYqDKGlIdpUxNc1j9gb1gMvcH0m6Qb6qdEeepZrONY5xXZ4We/vpYbz1iHONkx6y24
OULob3nlFsb61uFIT9hpeeB6FaLq36bAS4JSPiGPC+72YJotmjKgIb+G/jE09zLx3pz/xGAoRmOf
QT4WAEGYLg1aCndDEFtS8Bsm8PHhxR0N97L5qbPEwtxzxSgq6++51djWTY04JD3QNHoxDq+lt3d5
GDwzi82SD7C1ZoeyZJKXyUzgxzJ+MqI2C0U9kwrSW8bxuAvJNauWoRsRYKbdOiD2kwdZaKQ23nwg
hluy42KuBH44uAMYnomjdBW5GAriHP0ELH1W10cFAyWp5zxaxXXc03HxoTZuLOSH0uClqMXDT69q
ZHkgrVbEx26C1ZeXkDvg+/Uv6ya0/wzoBTcgYWGewZatwo4pYgatgJvL33asuQh75ge7UM/PS89l
Btx24fhblcYOgYk5BT9815KjYQhjn8erDgG+akjFgNE62f9dwMV6efmrN55nOZiMbBEbS+v6H/7r
Fcp++tQIciY1OZan64PuhyWfJvOKmfnBgZBNL4gQsGLAU+P+HlUh8BrOIldeDV375MiBUE0AlUxi
4hqdP9VrB+uYVI63ynGyzdOy3oYOn9BqLBGkJm31VsNjN2eIrC/k9nvOsfXNlSXd9ECPvL9GM5x+
XnZuENv1Bo+kVglsloA6oBDEmzQ4UWAlV+Ia6jUOY4lV1WJ9Pk1a4qcRmcQdoRwg4fCQTipwgt+J
dZPJieBYqDPNRH1m7TMhJpmYCT7L0xeETQqYplZoOltiHS6BqPsIElpZ9MqjE2Qh9mkME1mYOgMQ
QZxTLm723xjWoDV/+5on191LpqT0bA8luHmr8QrsPE5g1uYHWramQPU8wgYdYKkDgK6fHrv2BwVQ
71JAi4/juZ0qx3B8hkM2kAdm8lHZuG7IAMcZngJD4FMo+/9Zkcjx2idQl3Dva/Rgp0Mxlp3FnxjJ
UKNJeAPbm/GQoruwkUanxsq5kMbfLVQ3TAwbi8uoc3Zw6OSpvz4F6yDGaihySVXxuRT5PW0G73DG
elpcDgCGMelrD1aHrxEkp3zgcaqljSzRar00gCAFGNp0sxTFj45Ev+VYm/MKkHRH8WkGpg0Wxl9S
h3JDVMBukHuHf+esIm/qMWHjLpOqEt3PtWUAtq37TyrT/IYpQXMH3awc4LrzVJ5O4CaFAoq3vvZj
AThC3ux74DM1HPaDs4lajw2a5FqOXPXB0Fdn3DClw4ojQUZ7hFDjFg0EknDh+X/y7wb43OnhOlnB
mBmLNCTQv8eUWtbUbS0rbz5waT81nc53TFbcxsUdYdEBm5M0jCSfwVaiCyfXLN6HtHPJEh+oRWaY
cAG5zSAwLKRkWkzH1ilnWip2y4GB5t3HhfnYqBRRjFu5uH1niNOrIDyTFCMXJGSfESwNzbZI+sj2
aU0Ty3+QXzUj22sccncc4MbJjgbAI3uGNIyRPE+b4AU3kuHxenk7FIAJvlWcaBJ62Jy4yCYbXcXu
B9ptcsdS8xeta1cB0q7AefEF7YEoFq3ZWUVXgUhdTkX0cexCGBPOBJ3ZIarYbYdV+pAU1ZuGr96s
HS3o407IVhWtItfQoT2L2W8lfmSdQAP9fSzvQB95KVyiVzjczDzx3zewvPX664DyVatyIT2PrsVG
lFjDzSWDy9VmTZqwYQl4iIDHNykGMrUEp0pPThEZf4DTI866CnJ6O3VKMcN3IyfZ6xvkjpKt03RB
5mB5ugkjUBucRMPnOfZeqxrubFL7xdFO8lE9L3xzJLS1aSVeYWf7t0mxm8AWbbRxz8wQTT9FC1qf
qFaVkVjlUUcxu+9BvUUfH+zIOAhRzHM4jGoMVVxVPOWslgYcXqOLODLmOOkCqZDD07v3EPwIgImH
JGUo5aVeASC+dL09MWso+9s5afULqmNQsDv7Py6V1c/UzuON9bgzhO3dhehIsAGzd1xTmT/ED5QB
5FcD4NVVRHwC0oI9UdTz9pFIrsos7Vg3r+HOpVQhwA2bb94GBrVcKe0T0wKw576WBCpPLJKt3PSS
eJp4dNpQeQgbF4r3hv1BlJ+T8fTV+jQnsj3wjYMlFG2ePh1IXG4Zr1N8KpkGcFfU7xITVaKr604A
BBSgdQks+LzJgJ0juORuKwT6UsIkjj7rn+DhcOqBCAIZVdWtN4b3KZdwLV1Gmm2uL6DVqeOJdGuh
B4qd0+cFq2R6pK0N3SSNApuV2ibpzD7ewDKZzuGdkTvoeJHC5YQZJNdOGHMAqES+QmRviPVLAwyR
HIu8rNni+n6tnqatVgOSX1/337ibmv7x0FU4ZYsLamVLaXiX73hBgGIo1pHxNeCgcaZChSEG+O6a
L0l3b5PkqDmGf1PhvZIRgpwXQQwxJrzdyUhPnXXn81Aqqzw8rwtb42uikPQubGwyuMBFBvgp/RCN
JEMPVraUiPGWZK0t9TQHGD0izb6hWoRZz9b8QrdPk7sXKJ2ci2INlbO3T1TNfG6WCpfTkW6BLNgf
TXExLHdOtyilZ8JuEdGSWa8dJrgFeOLrqtWIzeQGTw+rEWqzBXljImWyDRN918jTRRBbiV9Qkeb/
fzm/ZxU3IM6bs2Z0cE83sLKaDE/tkveusj+e+q/UHMWQIoQPVGpGq1MSdKA7f/863bmTGxytIsqX
XLp3eGbHgCHMblNprXjITEt+6/MvG7WxhR082cNkOESyVSDFCC1ClwqrjB/TijNAPcL7j0GaaY7+
vbxB7qb6PEZ+SntYT2pBCx3kqu6E+LsthIS7Z4HTmOqQy9faSubH8BWq4bOzSqJUGVpiYfCFZjpR
cZlugPJacdwpTJ2AyX2JPKMakuLEiq8g3pRRmzqg6NjOlG/a4g7rDZo1KEQFI0/t8qlCb2iy6wn3
VzpBDKwmr2YL6uJiMtgPDgU8Xl52fHF54g56hIoJMXEb0d4vukujwkodeOYtGZjxQzeXS5bd+E2G
HZzGPr6HC9G+nuk0WNIpFdMvk414FsiKZslKO3VP9V1VTJ5TQZEem0TLd8lIr1Qdp9gFKAYdXOXc
bhMWW+7k3Y3JuUuiJ2qLtkl7EPUS3qbSa7tYEdocpJG5XJR/zOtM+iKpbwAwvbaWv6xvr70QdFQ8
v6PFBS+cYPQ/0B8/8qcAjXSfmRwP+0hiUkMdMIOc8hCNydaYBEL/Z2k91f1awE9a35KHAFCh/EaB
j9DjPH6fdoKcAEZ9NFV7ylYzWbOv0pAu9TTy4PTSRXQHhoXuAry2lkY94f4uTaLoHOGWuKIkxZLz
4nXd0F+po1A6K96UzP60ygSbxlmHsb36UZj9RiyJRCt7Ms9e813Y75sxgjoCEAnuusQMH3P3JRJF
aD/1610XRKvCKDOf2u6PUlso2JNhqyDNBtz2YsjRodY1oe+68s21/QBYKkJsUDkE1U7YjpZGjQb4
3da8xajjJP2eSrAAmLIdNn9uzrFxeseBsQ+NqfcehnH75hpjuv1mdxBJmK0ng1WU0rfyx8/xIe5u
BT432yNny4LF1tTgdRiPvJupG9Y5t4NDyLwmCjoHa59MzHR9e2K6lXsjOs0JWQ61LgkULuy9ResV
RZrVYvf54QWBNpmLut5FkXcVuWRPfLwttolEAReFHrRLZmGmneCq6fhVvEU3273DC1r7vpLIZY4L
2IUSSrKeuIp2V2hYaMVOwAmSkMT5vTnrUwHo7+oAhZAFTTZRKzB4os9lZgI8j4tM9rB15nHmwTrU
aAoT7azP06XA0nr7Sn0/tQEfoWaGPL+ZIF+EcqtakRPw3hj7AHodKCf5bs1lqUYzvEv2qxOsi5NM
7cbPtvwGfQeAyl6HWmBXvOw2/ifvMc2AzszTqifmCF9C1TYuP3LVk3GC9qYIwvyzTKUN34TZ+fYM
Y/Tha3mq2XH6j8HOoo3qg/2XvgfG1Pltvxhi9QU2YfbjRmJ2a6EZAJL3yZYC+o5/AqjMzPNWzcMS
9H4U2OkFaA4RzllaaiLBbbvKhBNf1DlsUaBGMotid6yaIrOHKhQTVmr5/pG3eJF/dhZDxwajaw4v
JApzd9ZK86FH2+iI1ttb/qaBxgm7fDss9FQ/enpMWRbLHmzotooIzoYKoTfvlQ9PjWOajeqk4Mc8
WAnWJT0KKBaHoLQbWhYHAqzTZcOPzdl+pgXXtxfVShA7zUFzYdTkVx8hamk4KjeWoTr4nwFOx1LL
455ODu6SLv1P9hfLf2x19M6ewVeJpqLR6uLBWxFkhmFIhzgpOiE8/qb5CPuYHr0YG4k6Lq6cvr76
PMHjvfDLBjeqUAco3q15Dqx0U7tM9gxYG+J//cH9yiZUlxI+jYapWTOu1mq+5+koH1yFrHBDRTIj
KB7KH9cC6koiphlL7ovitHRn25rnfudDLs8tVWfILbgjlX7g/IGrf886pxtdR1V5unnwAReKMOy0
q3Jre43Hlq6xl+5OwMSVhoE7B2zOXHIUPabeOdo8zq1crDB+FM3zWqV+HHnI9v3EG9m80nXgsJHt
ugiMhMTEoi4oILpdHnpVFDL9CuuUgCVw0Kxfgy2XZ5UFtMePUb6lQi/yLDNjBprBXKxTD0NkB/qu
m3YAz0MDgDQ7J4k2OLsQobUr9fNq5eatYbTT+LAwUZePNrW3bpJmfWruTurLddtdSm55nu2Zayd8
D/b3W0AutwWtAPWQ7p4rpfNvW/cd6/7JwKxH3aLfHUOz4pQDdr5hRWbQMsfwFZMgTaZeAdFvPxjX
dQ7IiSlqRjVfVIT/8HI9vo62GGFKU7owV0o4iN0ugeolwG2Y6XvZHmqwNbElPjbMHjyqRu4FLXMP
3sPGM4Z4JYd1n6C1itecXCRrlse4+0XrR59qEwB5xqbjC3+1RB84hRnE+A9IO4LTDQX+gm0VbGxp
GOv9BMChsbV3qzCqC1SZCloxbz8RwR3333Z+6hIFf1QwN09eAVuxNlfy9hPaMS7sPYLNsQ00Ocya
BPyZK1vV2NBx31pc7ay6vYbRsuvpZG8jHFPy7U4quaICRH7du1Xa6l2aQ0hP3T9ZxcrOxkiOAx38
58uYa7gDcCvRZSPJ4yWL572VQlQ09tJi89ypTDzsZ4sK3IwbgpldHd/KxeJvz5FE/m2pGr+uA2p9
2VuPt9Lkn63Nl7JoGB7YkDvT+Q/841sltZMz1c52G9we71eDWZ7Y7QYyCQi1yN3EkjYDQM639WKy
OLFnQO3D6kNxEHkcI9v5P7QuUKqGAbzgPY90FLXow1fwGbaKsmkyBspwU+9uwS4uMcTYmV6f1Foo
VhKbGVXdyNvDVeyX4Pl2KDPEAPSDyVxB/L4qFvg1NaMPYYB8N05XIAXaQDn0QbbkSTzLCRcRo+hW
rbgP+c7NYk8MxsQQL9BP59cHFGxzUWHDi+N85s7XnejAw3zYZtUkOTTp3Tti5DDXmAwKj3rFjELC
P4xg6GVS6RGFbDQvon4RNhVdZCYbHJhw2vPO4y/panRxI63abm6gFk5Y7OQ7xCS/uNdmIBOqEJNq
QG8ZAZQ4DuDpeLSEFapuPo087oZ8nzaoB5Ke0KdoLa0tft4Brbmx9ETkY7wX88lRHzQAfiPMAiFz
4wvsznSClEAfZPh5FXa0WONMMS5u07TeUo4ei1BpLWvZvd6XSZK/kBtu8YY3qOcTBmr2vhqt015s
UbQWpTQKXyOsMWALhkmMT+R5AN76SUP405IMgg4S8wvGwkGMfyOvKFupcaB7tuwdio3OTQbIinar
llQU5mWbLB4uXzXJSmsp+3K9RtRQZUftUiEa36gYMuoZXqxE7p7Mdpb6ZrQpmkFRRx4TggA5TwkG
4j+dttYk8frYU8ZaN1GSZHm+6lk6hnze6dGdPka5/XBWPqSjKVRSHjZ8XWIb+moNCFbR6/yxoi4f
wCM/ZxFgbjMH3jKp9Dj2I9mX+rL2rp+n81txJ997tBaOvwlQJyt6UjyUFtCiVO4y4oQ1mK/eRQAA
IWFv2W4V0wCQ2n3CSBLZm4pjqVLWtEeClAfgBtR91mlr9ea457+tQJNLgLotouWqt9m0oQzu55VF
fML+ge5nBZYxATtF/KZjyTXJ5eR1FIRjdryjAxi4dT7zy2NmnOMAmQcN5u4lUvmnjm1Z4tzLczKb
THSHO1E+2y1+uI3TigLNIP7ZTeJV6c9iUqBe/drl7uhbJ+3hnlJB1qdoZnMlzFQa1M4S3mehKVLj
QjYaUOkkn2RGyubSF/xFytyaM1zQZ4/jf+iTp5O9tvXqAxBROOfqwCKkzF7HmapE2RxPCHQkizDf
sz0kUFQpR/38oDlljxSVoseMO6fCiYWHBwHDUxiWwGu+ctJ1IuxM8p0nNIoySu+sDQ1D1mN50ndq
jCi7kcFvU9cudR2lDgA0KN9WAj/g7PO5NubkDfJPlS2WUl75RyHFFVyVV5jT0MZxN2/61AvWIR/f
yBcU+FfctHbrWNnN8FDSfrSUKJXCCmD7mSFN9OYIWMCqvB3ygp6DVp1DqtkYs/4KZDaa1Cwv3jbL
/XhE/rXrB1qou9Mdzp3R4M2PbYgth3+BtOoSCYQsn9qu3sRpqgKybUBqs41RMSLR+ERPnxggyw51
+wLfa7HKbNuIzkPpnDETaDhu4QOxIXy0g8QtOuJmrsRBp8TcIXX3/yps9rxgZhQFsR87LATXXx5i
sIAfRimaizUiym9ep0BksW12+N1VnvyuGiNNHUTmtFIS83gm7635aEcUdEOC89px4lc3VIhI7Hda
vSztJu61R8IuEryblfsafm7JMkY/fv0Pz/f12ylwhvqIr/+6at9KyYytDZW7b+Rb5g7CBk/p6FIn
DMYWb7BN6JChU1PO7vGW73jT9jBvE1Ak50DmNTbhKrrWBR61qm+yKvGPALlWU9NJgWJAPNThKNNY
I6kQvDHdslu2yI95EonwhI4+cy4p1MSkUQfOHw65KiqztkBpEGUGRNUVJmbmtUbksVfTs/Iz+OYb
c6yqV8Bhq+E5Vnqn187/YhrZSFNidYE/pLwmYFzZqp1Q9N/fwFf4dJK7SavlmukoG+NCGuTxL1Iv
sxAGPK+x++7nWGOmqeXhUhg1hFnavEXTJE66u8/RZYLjKKeJyRF09S/yI9+3MyvmY/DP/smIqkTA
qgsjzJjrDjUs6hGsTog1Z2I/g3vcRVTfTOnkXNWHAJmfiFEN8AraOH/QgOUi7Cxp3ujrntGEYER2
Gews/Pg39OSyfVmibnGR7TIni591sM51rHztTbejYY9oAUKp8sbbTfKDu8igqO+vk+GQ4z/0yxL5
J4U8+CU5xzRIn0ACgYKFQ5gr1cHZDYzCASiqp3bJOA/p58ALQOV7OF/w8PmN8z1+Ruof6e29EzYB
WF/9zAhQvct3sZlxBwYnfVhGCikGbY65bvLyPMQ1xRA24CqnPy6V4MFdLAZKCagCKOHR1w28V54x
Q/Caypyq0XBMcqTYq3heoYigRl257CyUkhw7si/6oRlDSTwQi1oCpvA7RPTMd5LHQBsO0nERIdcT
GBGrpmyIRB3DVfPPH2BCgtSSsq2RKPykHxsUkvP2Q4fs+yf0EC3gsNaoqibV8it+OapYIxMISs0M
NqZLakMwbvPE4U4yEsZCLhKwVmu/RiVBl6iHtQHKmeRs3Mm4vOLJOZrrZ1vEnsKk5F/CfucE2iuS
vIKy2wmmdN8pdnk3PDgtzmzhPSoVrUw4xQAI7Anh8WM8uL8OofWuYcy6vEjD4P1pJ9+J4w2tUQlL
lK6AuREyhE/J1q4REsEZM1hMCecL7AR+eMUN3iBOvXkYTC3xSZ040/52a9h9PVLzsUylw30daDFY
0tluL1Gzox7aefUuPG0KgOy8mZPwcuTkvuDBAjflkXyeXUWts6o8APA9gnEOHnmrT9lgx1W/ejVQ
boMJCrIhIGSYBiy7R/Rt4dqIPw3FyJAUdQpxAWP+sqANnlE6SxnfYxk32+CRRdCivjUlAmhip/UL
NZQy4sr8oQzT9U84f79wApGQ88TsnpIyzbKA55EVxrAggQRF1IEEmOPD+2f0nMH1lt0bR/+V+ja+
GeObxj7u3EKrcW6A4DeBFtZGmMsY/LL6kX51q/iA+4wALLyeADGPGTtjkb0ZVvMlJJMAIm+wFTaZ
D6Vv3Tl0KhMCNwJsZ8/K8Ybn3B/TeKm7qiqxsEg7qM95pTn9x+5priIGMiJJ1CoQpbwequQnnjPK
xw1UpgO1L2IH+dnOO0RZVxfL+QXD+lcivKFUQ3vhifw2vjzGoxTLM1eKJKMaejCxqZ2hjyJl+UtM
h7m/4OZrUa5if7Yd7P9pwMmQwyUKrwFNoFv/4qVkJtyDEolGPFEek63XeX3qdJ08f9EDoqfdltlT
SBGF+fQHCTg0NyZLM3c8yi98r+DMlr4NPfvtVbk/1lmJ3quT3un03GeyZPrFBM9znIkrOwMrmCey
+y5wsIE4mwGtNA3bITqSWQk1XkhMW/44hZh5HQwFjhgUkUIzfc7NVO59XOj1VBr/1O1nnNfLiEsr
ZpB7ovO7JMFWrw6rxUXQMHX61fz5HLJvRpbSZ+LPtjvzjuKmEgoc5VPksFGypzhshgc6x3XPvgEy
hiCZMganLpXSsq3X15eo2s4mDf2xsQNVnNbjYAKjigeQq6CPC2pK7R2ngNkG/EfU5k0beEiiHkSp
/zS7F4Gm3Aqp1yv6qNaQ/uS2eeAzxdCRhVbgPyvnFaX270+DmGyWoJP3sLxe0LRdFuiAd2Ap3/kx
nbzoPmS/GvIxSe8PVeN7CUPorRD5ifZtD2c77FzEL5tbtX2zQ0uqsjEdnxYXkHzMgeBEljsbcoXc
5lHqCf5Mih7s9Xdw2hBlxAhOgGNg17HMb09CRkIusvc0xBAoOMXg7A8zKZOZhkHTZLn/M9RDkt9d
WAclk4UnmtQ+uJCg1iPPKlIRmgNtcXRr/PUIvkgrcOtUSiW6Vaw8Zc9ACeSKkeLc0KVm3h/UuVjY
SsfU6EtKshUgOLTSfo7wQor9F7oKP2U+f4JJXR0wXHeIdDkXO2tYMRh7JTjXl9ZwA2AYYblQQ27h
EE8s1XnXSJmJXyxs6aOMpI/hKGlBO9fXJyUEjRBsWTIFCf8i4dmkIVuP3yAuj256cO4o9BXWqWFm
aIGxc5XFkvMIpnx/6+DMLD5ixBW1ZNmdEO8hSx5x4aq27k88ZzNSeyJII1H44+vQJeZxwQAseqx9
vQMw6QA5OSyr0I8REY2UlpSYB+afeINAvOKpDLoOf1i4LdHKwuaSRyY5Ik4CbYS8KOAI6YvEROXD
xyytPV/zg+zbyiJWBvaJW14N38SFbzkGQEqMJWlZm+FxjDNE/EB8BaxKk9oSduUhZ+jFq6o63+SM
jNQOxOhy2MJt1415Xhib1OOOEYifHPP9n7grd1Ye+GarieSiZBRzgCA+Refd8uoVWH+tOUIpAQil
XgH8wOk+52nO7/kmceXnDspJqHd5j0C6jNN9A+Rpm/8TKexDXsSHnVQ/t2wUOwbLfl1q7L4eYEg6
d8n3dd6ZC5eosmGjJbQAotA/0XPwMm2nZ2FdaY4kQGND1jsODSydO7scGTAYOGnFcQ4xzywuuE1I
+i0h7xgDHdfPg7k/Csenxd6BlOx43DJ8aRFileUGHjhdVSLKPTlILw7/KL0NGUxqakwKuWGUtZUo
7SnRPIZjMxjw50nAf++h07n1hD/ARd9Z8J8U2hhy8qwggCkuMd1D2s+qVPwg63zb5tzIJQfT9tYI
2u9u2PPZ6bRSnKZmIVpAfuk8ZiyPWTJTms74Hhv3KywDZpLywbSQ6G0GTWQgtCjwYtQ6zWhteOvw
Q3/5iYXgKul9/MBI2/Y0Q3qKdsZXTM1IyGBn/MHD9Der684olV+yr+tFPXZwQqznTmAuLjspGZe8
sCzn/ZSosK+hiZ1M2nYa2CaS83DgiXLkrIkZAATTby5aE72dmC16aDXP3vnLoxsbU4mOJDMXIW1/
QpqimsRTIHC1LsCGSQTCUV0VccG6p9j0NPjKRYNPovTtGpaeriCvamC/+WAanvoBN/fPE9GXeAdV
sUGWsgAb1x4g17yxa6fKuAm6yVv1/SbEKGU90vAp7w7uB62E4r66sUqUsPnnzoSVAbg2rkf7R44R
ZXTC3fCRzW+BeiECMH5SeWo/FBP0C1PBjk6t7G5bwb//jMLvPk+F08MZQD+VROkE1MgAU8R61Lzv
dxrrUb6t7EdanXbX8IMoiygobKI8DJ/bnR68XChcqPtrkE9q2H5tcE/PGZHjQja3S+jgzdqfZmTp
5gGwo3jWZVDaU4Wtb2ylBtvxwFR+Dx0O4gA/cvfVaxu7c9P+OMzj4iY/y4mDm5FJ2fn4ci0wNtsK
szA7osJRxcmHqjiESVdPKl/qfrmGILScIngYD44ZC7VFomqYTXcZygh7wunrFGmFzWgNCYXAYqF/
NTfKh/IfHKlfN5VnsdwTKU/gOnKtb6JSGBlrbug8XaAiUzp84mrPFD6QZQI06q9P/f1QZnuDgq3i
1gr/Fd4KfvWn7XBTPOkyleJPw/g4+4IZEjkBNmsi7unNAzfDWh2hgmCI9c5YXqWjf62Z3aDaFSYb
jrIaE70TG1m6G0v3uBl/PMeYiNN10eaRmVG0ViyEH5kcDKuXrMuvkvDNX8N5Gi9Dvo8S2IqQiCtw
tcJ2Jm3R/f5CyK3xID50XVCX52sPDRlk4EV7qbzNrNv2V/+7HM9qJFEdbu6HoiIOjghBViTCYISh
yn1EDafbZyIlV2y9JclUbfprGZr6nDqNFCyNRW2J82YRYrbViJAannHOKPny7uUNfTor2nMmuJp/
OtGW24QQlvhPv16nosWF1hNyXmqHfar05dFhu1q1g+Rrr69zXMVR7GykA9FNmWYHWH1xkFBAWb2+
RLWnTD7G+rXF55nHVzTXsKRBvFtrg3OOdh1oVy8Oh/GDik0+Lr4lL1AC7lqkhXxLig+/N0XSDQIp
5BXp0UhTHSOP+YHZH9kyg+XRBsl9OCA8Bi6t2lCekUxkBoOy0wrYezrVrX2drRbzh9nFUIOcNj7o
mQovWCq4FYRVgJFUn6azRuchIMDPbuEC+arfe/cfgAJiB8AOVvvSDTK+K6dq4WO1PI1Ta1ydMf6w
T9Sim6+CcK2betwttZGKNvhmhQ3/xIsVOX95OJvL3vCtYNiAHFHZMyDYbxMkDE/BjL4SpNX/mb4r
O5klPeCtqhBcZD5N6aHS0lsdvyjuWub+V2H19B/mA1+2Z3+BFa1aDRZZscph9aJcnfWsQiwf791o
Eyzy/iGLdKSpE3r5RTij0h12KgsFdlvUKldd9CSa5S4XVMbNz/FpxolkYty6e39nbti1oazohgMN
MWx4C5XqTOIGYHKhKzqFBdWhyN3NE5nqrX+cXD1+US6+XSJijafcW3DvtHhDOTfKBJ8eMR3PRBA5
cb0GdaX+AWkBhbvYOZzl3G3YcrBhInc3ZgTu2nCrcdqbKpnXnKF2j5zRNX3cfX9NmOrDhSCosw19
Uu0h3zOtBpodHFvvr/h7SQrwYyn9LcQfyGhIM/I33MuLTB21SNGJ1YxejGS7MbPVy8Te7CJBmFLB
avNV+dES4MbZBCugljpnugOCrzNvOsSPCAQmvYmH8GtAnGS4WAWCYO2heY2g17bFVDiaQ6/6bryf
cbReNrOK0+l8ydD+GsQe8aQ2tJyYeN52SDkowd9mU5IhSdoQyDvnqz+AiWU23NnoRAjrU72i4bGc
KFewbsbzMbSqX3KMP/bQhJzWC/Q+1jjWvX1z/Mp/EMoIbGEcER+NYBo6CJRZaqc06it9UUCuQa7d
4TAV4VC5C6wkbIzLynLWyOr8o8vwcPeZwbAYe98oZsOBbzYzxeGx/IKCDBJCvCaK9vvXxQRfDSrS
vT1+zNyj1RcwmvxX95FGWhKtCeHhWNR+sOX5vNJDSUThr1VQZEgUpdHm502ewRXFrzFf5rCqgXt3
txAIA3/LV78SXgS4CXoP8e4itTxJw+iU04G3ufmv0bl9bfCo4rqGvcFvAS2YZfV1ndxtJQmTNTNM
TcjCpIzjCAqGDLXHBo7/3sMHEFqdPnLDwammU2pLJg2ECl/xnpdoRCs3vYRGLahyDzA2+Y/om2Zq
our4hG5eCoPFBp9tg8Cf5QXeWmBgQcYDpEDtwMzx4Ccjk5DDu84GXkiy07fTGfu2TcYEBTHiv41d
j9oL/XC4szd1GFTsp9HdwnQdCwnvZTB596qAdbwGEsbblgS9hSI3wGMRwflcQPA0P/PcavwgBQyU
U/jy6+WVssSJ96w/7g+/pV3Rt6KeC1vPDDBTuKhyqBlE6soeXFw+FKKgAoa0zzxOEC9SjhwKNOzo
AkV1bMvGByCN0vfHVHqGEMvAYusmpp/+GmmsHc4JWetp7PUYthjlarlxiFzlgCxuc9sIuilgWzl7
V5lxLS2tsbIittP+LMZLemGB3tytzyy45Bfv97wC0rYxv4182dP3aG9qzp8nMnj7+W2lp99zNQOs
1baIgIxJysZjLRgrQUuw0H8wCgE5WJ85NB7tchn0HE7FF+EPwmSHmhqSxj4+ieYgruwckjLKzH1m
e7nXVbAa/tP39BebTMBPKw5/Bes/PO9DRiZHbfVZdALctfYe+f2XmCKfBZcqKziLdqWeHg1QZBtp
7E+pXNavB7YhC36xnUk1hXklTkm1y/ARNcZHaXBNkCdEh+EsHkBiEBzsfFP4bJQ1AeY7ZqtwpL4o
jqdZyi5mO4fAilUhZ3qA9+553Wygg71Uk8aP2iUZmrp5SiT+pcgCezxa4LlxoIHCrVvPAwgtuAsY
oxvxoHIkKwI+eErRnvlTKppaQP6qUyug87O2Oei59VtbYB1JKraZHVtkNyhiZ0hP5QOW/ZvtpX9m
sCJ/sZvgN6HjsGW208k70EDyu1KBfguzHG89Oae00+f9TREJWlDt6qaQSu0CoaeYeHxx+cxxrIC0
RRQfFY6HaTwlb7vGv1EZlc3/iC1y1HRaTWXrBMgR08a3BZYRDtbGHcgvSQRX2w2DQ4QwNyLF/8gr
RruJNt11GO002a/cX8LKXV47Zm5UfVE6NNYykyCjWDAUqtFyBc9xK8hq87VQyuSUzf6bqcWOuA5h
PeRqPLjFq/jrqeSIr1hVZ9tNepPrSleLmcRY8LR+1/5uqXMPlqUcTymrXkeC31XLwQh43zmm3kpX
nhZTYd9WDsyg308MfMgaGPm75R1pYgPAvedSQbaKpcFiTOi76iEUeFhNO2L8i89poVKxKWTAg3fo
p+dgC5pa+L3CxXW575SdfieHne/tWKetdMYSIpcC2WXaHH3ow5Dzq6r/ItNOs3KNQwRCu9We12nl
euUZ6B8htxDKMuXd9zAN2S1fgpWEz/k+ml2Qv5RYMCkE2xKg8TlNuFG79qDql3CDFnVeRSC47cTf
A6ItJwYC3TXQgM6t58a7o38Uy/DA1bFB6H/OrwiHE0Y/QWuG4n9S6cRzqiz0nTMNWYANKqNgxYtz
+LzhKxIDSbv7HGh5XycYdpLN+sKWawufOfVn/XNjABLSdNN36/9qa0Y5AvQ8z0MoqvwJJxZGDmqG
nl+sEoOIMHu2w9iM+fX7oZkeL32FrpOxy/g4AL9sdvBbmDCFkzcdY5MIWKzWjPBQEQ6CIyVH6pjb
yzvqVPnBT0CoKJhk8nnv1hFwJO0CGyqdfYy9AYDzYcb3V5hNUv+QCXNwfFggYPY8N9rV8g1l22VN
jvzCcX2owXPZiFhW+8//URdkZNfk9b7yvuYEmAsV/NOWyOBMZ33NAxBo6IroJSXYYFERayYJzcTY
4fWSt0ov8Lq0HPS+P8gvxQUNqExqfU1SGIacujx0d32Y/YApxkhwX6nOvACXQW9/WHG5KZeNddUn
ddqWrm2JLy57gCLTDYjKz/2HXJ72xAF7V8FvJ1Z+duzWRWbyOv6y6p0pgPvxQeFoLC/WDtVkdhSF
vkoUAvJd5x3fb8YsIN38vYdpQHWj/rTrVj2n3P8kuQKHL8Rm7X0zvQmy7oRyRK5k+/aJ2rga9JQE
CqvWD0uvqmtzQ3PqPPQjE9QTygf2m4Wrrfp4eqp5gyuf0Cdui/CveSnlVfOcIPLGS35jy9OJQuLC
buuA8H8v1P5lmth0VSrCVvkaxMoJTie5/jl8lrM+vO/k0ko3TR2+mNrg4tMVGBE0h9Kc8eZK+IAF
mhwxBRcr5rw6oyUT/MVeHP5V94qGt127LFncg/VXuBe1ffSoTvoJU2x13ZfTroR6FMYyMwjZODs4
CZUnhnyQf5Vr7PpU0DYJn5acxd0sxj/ZpFez6n16ICGsAfHlXqYtgTrEPelKMSkqPnQDZ+wmYW0N
mtm9M3LTP0dwBn9kiPpdU0SjBcw+nwbVjNjnggDGP2cDS4feDHVj02W6k8AXDKOsXXlDP0ruZkhL
x/ep/MV+o7XZPmbUEbSrH2weC0bVHCAtebtCL8zGUsz63xf9CE9HGqS7Orw0Ceo1PTPzUFTBOpZt
m6kF9GuN5HlpOWVhzpKvnh94KTOxEcJuvXVz4mW7TJGThC/KtVaaCKAoa6edbmnCGE3n7JnWt/OQ
ng6USMNVrdgbfS5gmllomqw9UX4CYCGhMUYAtkmeEABDj45ZrgoJuFoY/FLVwEX2kyn5nvCCtkOZ
A+xe5LLQC3SJTZpkpB/+fsl5Ez2Upy7b4mMvVcL7NzZQqyk+bfiU5k2Q9CJfYxO/NdtWBa1yy2ha
4uQrz7meuROo2Mv6KQIh4T+ZcGMLvnyZ5aZo05bZ8IH0QSHd+2YzhS1zhoqJR+fYcBD5+LF79Ukl
pHMv068nF0lFDhe+0/WsFmEEiaIq5EX46Q6EAzUKpmq+WkwwbL+wyEs1RRNiGQwjwk6J2coRE24B
lr6bbFWKdi7W4RV6y8Nj3NzvvgMiCMOUPA+z6utdhAz3FoyEYBCMeWbLXhMnTQLjyDXTXrx9DUFS
1lk1P6Vg3FKryplK8083jN8ckaDTD67WxdxqyEgi2x18wGOPPXMyMNclmPXgj5s02P/x8A3nQzk3
nfeHXddJDEImey7PgG4C12hIvgitbWqfdiBCnBou6ljAAtdOcfo6L5HsO2XHNlfmF2kn1OrBwTWl
8tChk3uosJ0F5e6WDMScp/hjcEiXAVKbEKGw5JkMfyySm94aL/ZfEpfrInBfypMwJ4jeLxYMV9Bt
ZQTgB9iGSCQMvtWRYbS2s/1hdgXFkUOMolCQ6wUignDJNl1J082VEoKTchRZUqWDHHhHQIy7Ggsu
kL1rMq/dWoXFzPy/HM1nGllAE4/2/k/g/zbh1xokIOXnFci5Xay/jyusRLVd6f6gnsKR/RoFdNkW
EpTdjWvpLE2oVJ+sdAUhMlj942UNXMoqaJbwXsSdZLLZin/fTTCM/0a+EjQFFdOG+Gq075TJgfz5
cCn6uC/XdBf2V4VYHDwNhAc2p5HyLErI5Am7WCcL2rlifyQ9Wj5+WS88tR5iZ8DM7lyDkSaNvmoc
iMvSeiOpBoy0szNclJOnVbgtiIh/LTh41lGBEQfLPGc+z+WR+IpjLpoH3bjGb03C2uX0V1rEXmBT
iUYKiW/fXpkpaX+M4IMhq1BXzgWBs1IiTTVti21sbwTyQUlf4t9T2Myo1kEWBeEGrNA7mlfdAV/s
ZA1xS6mFv9XdGOv+Rl+PLSPttySkLaf5c/YfuWKDKBaPXDFzf3KKnPZYEaVBSNDPCcV6q3Onh41p
vgH0U64wd83qqcIubJjUn0jOB3KPfNCl38CkMaNhMZqEjQT7NGjSYbDWuAJkaqOQXQ63UuXKmL24
4ijhbL2O8Pg4bG7VFyURCvqQzaHpce3UD+Aoe9fZBSC0DP3syleegjQ3vT4FeQ4nCU7fhDQEe+Le
twM4GWNlmsgeSpNewx3koWPo51hMaS9flAVrZ/XZat8UEgWL+6seLm4AyIRE0W4LhLK7g2pZrQXP
MJ6vAq9EdXewUt+fkUWmNmt1Wz4wlWa/c5usT+e1rHOXpVZcJGqEe8u/nKuGgEdFw4xfbDqg1GqW
5nKSDrEuqcC+LflcUow577DBhuelCEfHrqq1E5Cs/PduDKwAR/lnRrwbPUuDPec7PZFKxu4/+kPQ
53UgzRZl2R9UVwgK/N3f8JeUadcNomPQs0zwiwZqVmwoEJ+eyia1DdO76xjdF54amROlU6sp1FH6
cwTAVVBpaau7lft3spIvftVJ7UQG6cKhQm95XtS97tir4lfGYCppkQ6uP3+AezvxrCzLK/dOX3UX
Kmg665/4Wr+n8FrfT6Y1jJz+oSRhZHn5W1cnijaLliAquVNcT8kNz3YDtUuPhJpE1BxtfghqNhB4
bMJ2sRTfi4ww/J7Y5AAIc6W/0fIAL5VTWUhIkmuB/enjc9xn9F2q766CWml+op+AZpN+Cl0+n/rH
i/Yyge5rayBQXgXjzPngR0tffF77WJgHQ207tsfSLdiHYDw7hmPxCOMSpwsiEE5JbliP0EJBFIkN
OCe92T26Nf+B0/RFu9xPpSyXwyO0Nv/n8jGS9BGn0ewW41qUndANOLC4xJFI0pljZgr6WsONeduP
2V9ZEZJ7qtq4Rj/A4UxsX2FMtV3CE3+jDx4fGry/rnJ4+DX+jFs1oTMqHzKyHXtyv+LeO5R+eQDx
Xs/3n1cPXjQFFW9qnFx333SaiE9LpZgluKiF2pgKTtWMbj2gtTMbVwxC21fH+zeXXOhCVABwWOSo
e1dL5BuyL8z3kE8G/ymANCLFij4mkKreBalnzF5LL0gPLRYJTUj0o59zI+fpo764D3I6GA6+xAmx
3peUy68meoGCLqkvA7lAj75Uz2cndLZbpxhN/suvK9WM6YfEz95i5oubgBHKT4503xU1Kvmd9clM
UFaPbwM0VctHxZedNQvofG+jY4z7VNvTcI7GSyWJ/jfjKyIxiDfDZhY+KD5gg52WkDaAQj2jUqzY
YepbE/DnYCcKmeu+/gEp/n79hpabEbbyejMNhRnre1gohIBLJkrAbEMIIh051XYadV5J0dP2tMCM
hkPOv2aZYX11pXJDjmRznDgm5e+qV9/esTA/CPTeQXacL+i0OdpHxteTuj4+jsdkGXO0iEYyEQyx
P1I/pknaLrC7PvmD1Mus660Sif3andrcSlVQHv2FSbRqR+JlcssMGEl0CBAZBmTwz9mDgm6t6lj1
YIR2aHzexXfYds9Jur2PEAlmxL9gLFOSw5tWqV0RdUweUAU3pE4eCZQSpbwYNDnGk3lRLTTpV6Y3
t+oSeFcTj92U1d9/+PBV5qF8aJFxy8KZlD77ni9CqgiOqj9DjwON6H4Q9Sil1B4TPk46EgwBchaZ
X2/LcwhJ4DfkjLG4o0efw6KiYQESeMLoI7sZr3xVdbnRZf+4Q2zVg2OdiaHjy3uaHnHwT7C0I0j7
SYXmzOlk6cZ7bmQCnlaiRkEvsXwwxYfPd3kq6o3I1Ql4JHO99LSbDOyx5bi3kB08FxihdpSPeF/F
FmArpp2EtX55cyuz/6NzUymi1EzhPbcPb+8ghM6nrURiW1YopHFhSM2n3p41uDZMCL0KJXjPkYl6
0whTM2WEQbbnFyWkMMS02R7EO0XZ940RZ95k5OtVLGW2SsjsTCQvMkamtX62RqcY1jfmNsNyHAoq
Aczw1Ip9uq6iZUh98Ht/sRd5wcjc0ji54BQrj9fUID6dCe2oT6mKS2a3KA3Fo3K6shOVKJnNHXeK
KfeAbihw6cVBoZ68he0aYpK3mG5ade1z9U/BeVVMCUzElXH80BbL8eBvUmtnJIZiAfM+i7pIdwYe
S4CJf10pN+RfntOyo2pLbByxNfxGqTWoV7s1Kd5ew/rC7yrDVnRDOC/ZO1dwiQqTvzvHtRDuXbsa
keoPmB4GJgkoVSvZFvcCdkaI75yC7xnIdTyGN+pZ/SXrdb41mE55+JslzRDeSHL/cnqs6YfnbV+x
z8ET0xIulHc9eVLMCHcaoUevnWO9uWg5tit8QGH15Wv7hygCjPm7T4syyZpNcDrtblPIkBj6tlds
eGkeaThlwS8yNR1uTEiKRwNt3tLp02EeAntwo67A1cDvnbhx+sZjSn6F/CJn1l4ovcjN5RML4EV/
PUtKsPuA0bI7aZlGmm8i0vQqFplnwEqbqbijpYbr1WaNyr9G0kZfPub2Km69JEIb6FjZ3rNReAHM
PKbLp9bZrqu5mSzxLmcgIo83HBSL6fNrB/R2uPBrwkF0/Fa4JMP6J+i4f4e1T5VchFxBozA/qVZ0
bWI74hC5TJPVIe+gSsuzp6p82CQWzs8UR6BtRKGmeFTcRIuZRrzusmmdJHTukJmSTCdOpn4YpZhS
5zaDeUYWUdn+3U0NmqFdm9hXpo6RlOekE9NdFawqzb4Dtk5ES+Rw2YRve4sJz0P4Cf96aVg8OuG2
J/bYRKPOgif6FA85MdCfSD/emAw1bSdi14Q+c3v/U8nX/AQfWEICrQ/vPF9jX/XMsy9JDULKQUaJ
FWjchMRmW7hR3UJtVAbzZFJ6aq+E05la0QpYLJCA4Lm0bdRszYtAINx/emo3JlRwFqkoHZwVBRVA
memYY24HB6y+Nu6OhFxN9U5r0vqdkn5Cl3zrOuhqSvQG/KDNY8VT4EkX0omazas7iuU4WdLd0i9c
RQnSGpRMYTOW+cSwWeEMPSf7TXqlrX/9h90hqv7eDOZEYIQbw2UKlg0xOzPg1XuiqfK9UfZ24OgP
Y8FVFVS+msfyx8c1w/O2qSUVTsszDcg5Hk2kefDbciPL731QtQEnmwbQR9lANTAUeYVkzUAlgjNb
I1o4Se9h/pwbBs6ZMn9ihvfxRwRVy/TTbC+yYsIObsnx8GlfzUs4H6tqqLXfgDWHS1u/Yxm7tWXy
6HZtOdPc4liuDunELjky0VcEqBEQKxVhTVgeq5tA2ATulfI2hgwmmaVTdAhO1OGd58JtrJgd1kAV
v+iw4P8+697HPk7MBbEyBMZFJiZRuXbdmLebCbDM6f7lArU0jaEQBAX/xaoVy5HPX4RMZwSVO7rF
7p8e6+pSFMPuB4b4nNEOcJlPbvAnId3Zuj4nR4FOHWHC1LUhvelpq4FaxGFhG7bt41FMxCTLGRCM
s9PRnIsyTNyFCXVTqOOssejvzlrNwXplvtnhtRCt8lZ5PyRn8R/zAEAHcozr0AI+FOp0zIcF9g1O
yI5zui1F7Y5daUiSlA0w2Gd3oIg/dMZzkbeVmJkrpe4cXzbkQJfziZ4Y5vSBHBfOHzjfTXQuhd7Q
Pw6YYLmGVYf6x6CmMvzc/nGUyHGCyW5iGIBU3ZbeOUAzXVjPsfKyl5KMqHfMZPwOrpTKSbgDBgwf
h+X1UsvnKoJ9pxiDodptZj25lbgxMLnh6BTkjvrGaZIjN/MkIDSi/ChD8SpshyW+N6c8dDNAaUQZ
CIRPLToxs8Mbayf3RGP6fRdcMM3JPmOCmhNhQU03sPyR/Emufap2XFuIRxLuFZ6NgKRgjJ86lWaH
I8/l/FB0kvMOuUBTcpA+mX2ocn0yKU3yjDVE0hpFFgBH9CjhstDMr+QYQNv/uRfl8Jin/DPtGw1A
BMMr0zWuYzXrlmiSD0jpg0lzpBqkKYuhJAUukk2Gqi++a+x9T0i1fY9LSEL4NymcRS1hO2JqFMdr
Arr0YGv4246r5ugjJZmwPbTCdIfL8M8MvYUE3XpzfLx+simt1o6LSYLrHPhCELStUxE42vqzwG/a
oFGGonjSQ8uJmwftMKTjx3JJ6Zo4hqjPy5/17jTeH9czY+9J8wK3W1lwgqzTLB3fGomWidKFo0uG
HAJ4/+++d7Lh2B0+u1pZ4kQY9yMa5LAXI9Huo3ExFUzk6h47AfFi6xWknj3ixcuGyywd4p+zQ51z
8gIzxFJF7ZrkfY4lVFkcPOD/GKy0lmzz9JUMxDvhepxlAWTptHXguajLjAlG3Ip/mNdQFZosoie5
NjFWHzIyY/lBdesH/0/TEQ7/DIcJv4MGJhvQoWZKC+tNEoTHlx7ZnGpCTHi2x30prQKHKMhxN+x0
ZS0arL0sXLfirDQyRoW6gQKdzgt0d0Exoakm5yGA1a5eeqdve5F3yvjttw6AVx10RsPCmr7YW1qA
rY+Ve73WRnR9ND5fjwpF/H2nt9Iy+BUNe4oBcUqQ4WgDADPNZanoylxW/tq+G6ZCjdi+3Mo2+b8G
7YFkFrdj8rlyKNr4ZK2qIRT3bW3qRCQGglfBptLFnv1ge6uEVP2I0l2QV0keSpRw43vMbxrqPOw/
MrZvubWEOVJv5QAvkgn0lUb463xukgfenFBRmt2MgA432GUTVDTrcpzLVcvDE+1YG84YBo3wapO+
UmEC8jVzntd1pBV16CQ1/tTYPlm9Gv+2PU8s5DvCFghuh/p55O21F+bN0dM5AsqDooU3iiXIKvEs
8rnQ0YT9HpqG0OxbWT1b+CG3DIPoh5z10qelSWE2TV50M/XnVRwojLo8f8hG94uDcGx5MHmnFRTz
Q+YJSkP2MCMfyBl6FxSX43NPITFM2ExEcDBYlVbSFe/I/2vPSP7fNLubzVIcLAnmYI1iSRX2mlBl
XnWq/2IzijcxVbdoXB5K7KElhjUH/BqpdDF9yp2NtuRkFrsmSDrf6Xht5NZux/p2Lfo34Es7y2v5
bFhqXcr11HJ0gWqexaXzddYXjg7vX44kFAqtSFKJm8GPGemBzhnIgJF5TlvRumQVPwDaIW+4uX22
86xv2raSxjtBibGbIWlxvWN2JOA+HUigzTIvxM1Pzh1FiEEh5UWf/RhL8/IRM+EQQHl+d36vSf00
TJt3VE5vZ4Xcc2Wdqq+2DQ04UeRcAC5urVfn6pQ5Jwms/6RQV+s67JYtjO+LvoR9Xijk+taw0fY4
VOlk//JLI1xD9TBRsnMYUGFc+XWAby5v4gQiqD+0B1EhbmJwA3GpTk3ZWaXgM/If14cj7mOLlEIz
M/HFhB6XQNqtFfGvolDXaVOcQ8uf+fjUqJIpG1vrMTQEGHIsh3+PbRY89sBpwB1GV5LdKL2JLSh3
3A2olefNYAlh3tau9gsUnxD1zNDRR8F4SpNsZ1kwhHIh9/YJWG1oZnXfU7AtPRzvamP++GV4QHPW
Qg4pvYGmttahcGEZoQhRHYpZLAWUchlWUW6FioTJoMxtSAM08UWCWjziYvg5LvZtiS3dqCAEUsyU
rZf+XaWItaIR8JcAsqFjXZMojihaXiZF/jZ0T4N1dEs6GSknPHS1B/au99CXgunILHSnTl+eX5HS
5t7TIfAGf5WVofE35ptAKPzzqX8Lkn8+XddfHZrWZD0ZEEld991TA319imwuIS5L9RXnslNV+Di9
TrPnUuk2kq//qxIFu4SN0NLftO1gzzbV0FdZTvCNwU4Kdgvsdb2DGkd4F78Z1rfGoKIjErF2WM+k
Qttm4cZguF38/gKNy+dSGbDjfoBfLtMQDbwZFtLVC+mJOrawYbyU2RaAU4Pf3T76/cKJedcim9a5
3EPdECDaujbAFQj4QjSGgjpc2hQG6MRcWFf3/pIgjwyzFM+C5sqUqu5NmkQVIAiSALNZr4UZiBAG
hnYGI3wonRJdgQVEfrBap+xKUCVU7Dicv3ifCjaGkopCtnKqPqZ2VmeWgMmud1tI9ZD8k5CpShbE
XoYEN09kCt7jCTEYs7aidIdmgWnC9ydw5xKlEFPonhn2Fo+wGJist2GlNA+h2dvqx3jrpSURVrL5
8caBeeR/uT5xKRnkNQ45YbVcTXFXd3NBKwg5S9ITS3fX8acAeBz3lu29egvFllrlABMNCjT5fjUr
9eMo+0k4Rvyl/pC/2NLOXXJCOpO/3IrkU+M5kJZ368KoReCEozjN7FNgcWuNnpfOhBR/6ArMgLP8
gK549vujXDVDatJTR84Zp4K0n1ywTS1T9qLMO4TMFfgAwrcTICx2eDN99O0cT90haVv8m3JBqR+/
CHDGakn5IT4/tf+hcDk0+riunoe0abS+k1RE+r0KWyRAcX7rf6qh4Eitm7cWvhz3e8jGqYHVC4mx
4Qjn6o/gDTGTkHfbOFrbQMuMr9A2AAl0YmULN1Hwdjv8Zs3wzOl9pRARGSFCrOTGmWsNqham6JKn
t6Nj3+XngUO6Xlao0B6+1iESz7oeLMKLOEteCQu8WE554eEBp+RtGTfxy25DyMYMvg/1KLIHOuCe
xAQxdvn/h4cPiIw24jmPI0JUWbv8LyceI49ymmgvi45vDjm9P0NRwnMB7Eas4TqGJhPLJ/l0bsco
9j0Wtow0zH2wwq2zO5LHh1dWRNL1IoY104LIHBwT7a68zLDSNTNLPc4T+fE8sjCuUGX/y+RArOFt
BZLuuQS+UePb2MflLqJg1J78hkR8qJq75bcyc8BlAVqLZWvGDzjWpaYO3Mr6x+DmalGtZLa+ASO0
Bl5Awz57oSyr/Z6TssbyjLmw8mgNk57/7KZhXg9phdX+nSzJ+mAw56FMarLio//nNLhVojiQBccn
Z5uNZW+6Myt2ia1LiqQYxu10lGQ5H0n4B8IgiElbFGv7fbgkm/e4v6Y6BVwYnOfF4ARQR9Ui5DUL
APIeyBW8AiwLNrVKq4PCyKpGhinz/mRJws44gMnmi7bTUTLmbDCUty/Nf9Rd0nlzPIRmhZWBBylm
y2RV4dq5UGX76vZR3QpBBUH7ZXcP5AZw338Z+zTtM7cFJVKVukORbzucpXxeTzkEqG6lzqXMiihR
V1UBWE6at7hRSBMWyfH2BS1S6RzKEH0JL0MEhKv7LNZ/SCgkV0bzlub4Rqsvr1k5MwJOP7TzA0QO
q5atk1dFt/KqnkJDa3Kkdr/LNNzG/t1LzHejFzlmzX8X0SEXz5YTmnIijk7LkCBAN6cZ+N4T+rtn
UxWrxOBXxbkI9T2z40xbIeu5wfMmNzDmm6oxKz3A8F10lMnyL6lFXxCF3yXPJB5E/R5zCzuRUrQH
7waNVFEZlsHJRg3PUhPusk6Kma4mqpItomgYNkvg9wRfKZYoTKCKgO/vjT8YeaEZGGzIYt2eKMYz
APXFqxU+c59vT4/ciTRD+sxd6ho9vvQbLbZMScja52Y/TxIXGzXqBxezSxlmFTwSCyIZhGOgh3tN
p25BvR87lwHb/p5FbVP8O80kKZRtyyND8ITR5e+q7yN07GlOmCVI6k3d4prJax9s2teocq00JGLe
8IeZMMjS56+cyBaz/vEBKFcIh6+pJemFUPUcr8AV876CCHSeih1ZlR8Dc9PlJ6RNepBJeMYSKLWB
UOn6fscg4gUv9FIfn6YGEoiiNAvuEKTQ34WCd2sjHHrSsM0yhrM6qbFj1zpCL1uq6JzviQse7RUA
y8cYI9mMeTrPJdFpMBWYZNNMB1V/zOQDsvg3L7O9931INZ4ezpWmO1T5KcdI+r2HEi39nVBLORUb
eKolgiaPod6tS6tIyXWhpgkSkVfhtr7oj4uE/lh9VwB8+h7ov+Htv7DbGui5vLYdbW7jJiGAnRF4
jyFJ3Xa2AsnbfloIJNBjGyUxsv0F5wls7raWxn4a2glWB5I7EpsH3J3SYlbFtzV1Ho5+uqsTXjgB
MOUo93coABgfaQWZqCthaDvZ0m3cvqkR9R640D5/yNaVMCwlSF2k4FsiOhgVr68JzTlK+VO+XPdv
+kGgr12bhj42dJbD8HIQ16OZ99xPq1MsOLrM1pvNvfQuu5V8xuoXArpNrjDJrv2DxMKgRXXFHHRM
t5K5SMoYQPdO7l02E4BHjGMlZh6sDYRS+L+SaevQL7zaKaJnSDbA1r2sf2HJ1w/ORfJFlknMhnad
YNHQjKiV/loXnV6+DJFrIg1ufYHXXFttncq41LjW/foirMYxC6W529KFk+QxEG3CptXTdMwoXksJ
qh8CXW4vL+AaXhDEic4aFhiCJfqeR2HXjcydyB53cPAdrTVq7psdwySKMcN784/608AMuCoMbPes
2bRLawU7DyCFAEXqY0j1i+kwyP4V++a0GopgaiJXpYd3SHYemR9OTPr3W7RGfYZ5PcT42ttTX1pH
so0ylzkA98sw9shCEwfFR1ad1dZAmEFYVEg2oOW7QO006C4SZlSjwPWCFxff7dtKAW7bXHbcrHDN
btIynYqGka8Ixs6rdmE8I7pa+lGbZk1Cdhcb5WoogJyVNsDhRQGia0GlU7k/1MhUnTosFGGbnmNw
KMlGs4ZZE5B4yHMLlHIH1H0HmkhWF3p5VVXVKjHXyYZxNoyfKPHGNntLcqsljZsFShKoeZ8uLjRW
z+U+7WFCcCchlLU+mQf2+rVHuexsbEonnw3VTSrNRNvDbY6jBij20GqNiC5CKRX2HGRfXqu56a3D
Kgl8EVRFFiBt88CihC/lmC1yC8/dFQ1o4Qf/7d3yLnDPHgiCKag4QrlTKXnZjvQ42cjTZWcqkcqL
BTeqh1yhpdVf10SHl9Z4BqVf8cftOS35q1Fi+2LZvfQEcPT3ujDacjRS4YFOY9R9GaFAJvl9qVQB
oAJjeCKF01Cnn6P3TCXkf1PJr2Dyr+NP0FCvaNknAaOPkrvQVjZTygDSz1rQJ7F8U41BEo2EtDZX
oP950AFviAfKoHOY6YtGIXEKdOZjLva8kq6DzoKK56/p0q9ciRhkBGP4Pn3JdRYsOFx53RIxnQ9B
aUkIuB339mieDhD33TnDedG9dSsRuexFLA8EbMm0VZZbmOiDmmp36coInoSyxD+huuO6PgUbhhkj
KigtjmlwtNq/CeAXMCSHgjF3mDIZVBjIaTqM4UdeXaXo0fFAI2OXnBb6rDB8uxRRZZ5JJ8iDv9at
kcIn8QZY6dSWoI2dps41OXn4l9GEhKQso2wtDL+Qpazgsw86yB7L28rIKwPjLITX1FwUKrZAWHkj
5Tyni+Othdete41SLqfHC5iB848BFmGnJCelUhCrBwF4Fx3r8JB6yIOS2E+NN2Lr6RO7ZJbYew9A
68Bgzvm+5CTJRHoeX7JEzL1ChwQyakfRzWlDrWGmLUEFGcBH8L/0y029+MV88GziqmiJgc1OjRVO
ufbdwgpOuzF1aVVbwCPDctOy734diVRNSDE7Bh/mmGZqWAp6v6M1k34VU9S6N4RtXlQcOlPN3UmR
uMohEgKO/+695kM9Naqj4qu9x9KsdZQOwerjNryab9FH7Vi8Z3yEbqS/E7A50JXtLJM51bWNqwSv
uUcdbeeSgNB1dx861uQxANRkf5nYPAkjz3gZVo1IjFZ9tpaj/6Rw/hhP59oa/HIl/J+uK9MOWt0Q
A+cAXVN7AgApuRjfMulfzC+iKYmUM51DMLe805cZS190x0fF2zfJV8qH8Dwlga9bKOFvAeVp4n+S
R6ff7Z+KbBcdD/OnBk2HeAWEof36FSineTsveXEwoyCFkrlpQt1EEiLq8CxSJfJMafNxuaaAkqdF
OKmrGiKELMg9othS+wNi8JPsjurfwMkSimJpm47kIbOT7m+g6Syll7cZQaTwffv5dxQcGZPmFQFK
+10LeMDT3xm7zbUCyiPKOsRnhmbn4sQH7rzdLq2mwrVLOOOWZBrwb3q/UovtJr004Fd5vTd2Sv4g
pei1+IO/hQUZ8TH6lZTvFZvAjtfunbYB7QJrj9c0Jk62cFEXLV6AZVqIz9njKdVUkjvjqNogr3IM
zeAINROr6lPgiqG4ygxBxBtHQey1GwlyIa+SY0VKImzqjNC1TrJWu0e87o+MAcgUaWcfyIVxFYEu
UHP7BXsV5khvUiiGMFMSj+ePaoGZ1MK1JUa54xxpzx7CGdGmGFXzW7QuWOYakbOclKR/lHOdulkM
yHUFOYcnPfEObU2SZ9N3hNX5zx8n7nUfP0oUFCMrJz0tsVEBPgI6OmdH9T9/WXrv9nWo6S5hfHT4
Bp5vXd9ofTV1Ox6AeUE434jcCyRQbcvUsLJ7sg+AGQob/jfPBRxnLeWaTjpxvwKZ3+77grPjzy5N
kr0ByL9e+UTzHY1U/gCzDgOTZapMyrxyCwj2e2sMl0Yi2ZDM+iakIxpe28cf8YSH8vOsd4xAsF4U
ZTjmTI6Sa+cMmh4SO0ZBd4UUe8QQy3CO/bB4hrAzLlWsmi3mEJZPLq+dEp01oc5NebsadT79Ada1
e/xs6q3VqYG4Aqbd/RFGgDwqqtz4jCV6U8loMkwGqA5NwijNx6Z/i8asXWMjAAqusVnlYQQtfgAw
w3QlQWhDHLS23dZMQcNSonUP69HaeVckw4x/PZ8HH/hNX/cVnLtnqB8Pl1SNbZCcsNakS9RR+Nzp
bVA6+lpq2wMFKyFqIIzyjw2pOh1NBspNyoC/5wTe/ekwuHoPGV668hWcgsBejpdDdZbZQd178REo
AuB/FnLTZ1ItCdFnsOU5WAso22pTevbyDBH+oS9j15nZDy6cGl6McK29cqhbRsfKVeFyT5wBujL4
HcLKm7tJfMooaipfh9Nx0vPsToV+3DELumul7nyBWioP1jGsxsvHTvwb9ff6MqTRu5uU67d3FTuX
zXoqLHBhBQTSjoxTKqxCZ6UwoNQ06jl/O40Yz9ExC9O06BAqiUuMVNkDzGaBw3YGbDjyJKTdaUKR
9wAZHKxg/7EZYTQBfYtkhuN+4aqnoPLIls7Pn6oK91Mnkt9JG8EU1PLBxJVn+wNJysODptEzLhuR
WAt6phZXMsWDKBYnDYnTMAU+d9Yu6zoIn0tqqw0VQgs6y8uANoSS8Sam9jmjOxNL7ng8GqweZj/v
DrrYUvyTbEXigd61eIxGiLGttvWmhij6my3zlgjzz+UcHdNQDXx2ha/3pOej0Qfxkp7Gf9ZQ/aZT
WzVmSM+tH8C9p6+AmHo45Tx2M3lJsLQOPh47NpVGa2FESAWyz1/vOrt0Zm/oxDJ/wAeDYzudLzjL
Pq5ZLhWyyU3LIitb8XnIzDxcyHD7ejQ3ZF5sC90l+bv1noZohXy5EUl9AcHsz3rdOmWHx8J6V5cB
CEaPKJk/FDqCeVPpqEDGeQ+3TX+AyUcG9RB2kqXAPcHfmFXEEw9Hy0zmC4oiXb6t1CQfUay7ccnx
OS0HiluQJBU0wR+oO6IDrnyButI4K/ygqICi8MUYFtYkHDPZxby2igJiGEnuC/XOxwSSkQiWo0Ta
GYOU3FlgiGLciWt8bWNyA3MPsupdBTVA6as9OjXmskQonTbhTrjUiwptHviJq4EDDjdnnUVlN1sz
7GoQ/wUYU/eeF9aOyAA4RHsw+Lp1/fcR1TJkYuuiEb5/Z4+vVaIq/MisWu4BHthrlgnUON5pN2ys
7Ry0W/3RBJJ6tlI/racFIRqOIxsMdWOVuMUKaxXqHAiWonyqUmghKMdCdGuGJOfKSd/5xYcqCPy2
rP2ydZ7vL7ND4ihOpnzNxvQsAmyjAkyl7a41MSL6F+a+X7eUqph0hc9ASxjbL7Dlva1t9AW/YeLO
LnmYEXJy3N+gXJ3+llpr0E1NDlze8NRLA07t9rPQUFi2hC6NdhsYZlZVj52Iqmi+BXKPhkVt0hCl
EJUN+UyTJ+MnLclM8H8aWmj9QICsB3KuEtZdOIvcHwYt7mXZYA9GXG6L/BHaxMYcOyj96wlaZqSX
cBI8KR/uNLz9b1dmwqpCR0ECxICY7VynSX330s7MiOxJrwdoJeTJyhT4zdC4amdQacVXFA8CdlAo
vIIuaQIva8Gm8ixzSBnspSuM3ZL9ev0EByG1rVoTDkO7a793l919kCD5BsAKz8Jdctd5dBYY3tSN
C2BipOYaiA+4W8J+KtSzK82mhTPkn7h2b6EpKI5Y3ZyFMCx5rxynsxb+Fn4LvK5n1du2lxzKwg1S
svJZyuy03gnaJAfnraKPNDulTKQVnJEFGXq29gQO1Mhu8DzboT6Gk+kXpZtdYllG0rkuTFvbg/lk
MuDe1RZJHghOQpt/7BcLoBYkTNDu8eu+ftini3l+JKXFAVu9ru2z7Ruc/7RGkilJ6NF2Xz5FrBDx
Fi6OB4UUARH9Thonc7zFazNJBc2MDeCmQyPV8VOetUyJcYByl1SJ0jZTU2WTeav9H1GS6Ps/dJMj
YTzO2q9PvC7EWqwvv7Vb+Jyyayfm3MGobDzmWOO0Lp9vXl6K/2hf4F3bEQjn4qKLNe0c8E/3t0hH
kO3WP+TeXVNhfJ0PFraPAUnqe9ULWvU1mv/6tf3N5nJOfpiT8zog8FbOVMfXW5cbU5TKvROu8RS6
HksY2WwXozSqRKW/QtuC+dDlg2pOpmuDdygM6gDOLDIuOgpTOzt5MVNpgqPLl8iPU6Fo6a38N3H8
n773JI07WNlwuWFOqBsdFe0Xy0AQQAuhjCO9LETNjSDAsKTubKBZdFP3ZzcDoFs3vh7I9H4so0R6
HRlDGb5Tj/GZMIa8GHV5DnmfV2/JKb0CoUr3Xj3VKy9euptCSlHA1VluvkGpZSeJLO6mpu/d1V/e
RIA6v+Q5HyBxNnpgWHvtKpF5GlAz6HhbwTXb1n8qBCYM+rGxsLepWPBPEk4aBMfmFGyVKpdMDyzI
7h8EMV7YdywlWVxone6y55BkxLP+iMBU2Lqkz8ZkBqXlmp+xStUTET8eZovBXpc8mPBXrachFYfc
z1nhccIShUKrZ1PesQlfFCIUYzWCR4pYKP4NJtX2ONphyvJibsXpy6iwG4NPOkm89he+8ODRarAj
XPqEXkCImcE+UpGOtMmSpQUdVmhu9tKoIVw+I9dL+EmaT1BG6W0pwGgvTSNcI4X/56ax7ouGyscF
RzNh6YHNI90yFDS2IdJgjb014vq+HTd6LCw01Ypv+kCn1Qm91Eg/Ev+Oz5FTh5OPYzv444BuR7YS
e3NqK1yJiSTjbcptau1VqkuC03s5rmOx3Zqgi1C8UBDHj5J6Vgg2KcwrMXHVUc++fWQueB2W/mjU
QhfaIZySJbHOj2EMzfjmCNiJgaBCL6WQXEJEZZfUpWbArJBu5+Ni+MVS+RTLeWVbH9WsugSjgsDi
tOi5pZLLmy3F/W0btNIKuS2/ks55oJzldVQoilhGtYhd54UdUtpBvOv0SXzrcjIVNQT+TJwyHkXk
A5b3Wq3m06JnlSFMKnv6CYL8/C7zpUZZ1/K1MfPG1pxCpYUAhwhcbLyZZnyvdP1k3m8tOVvKTLhc
pbiqRpkMMf+LJU/VJjnz4OVYvoKXdiHh7p4jWCWZq51so3eyRvmFvMpPPbTWzZObrs4bFoDQ+/iH
z4mJQ9VEDncodybX1NPMiM2yAxA4x+HLlVdY3crb5QPEhF+j30qYG6VJ9nLqUO+ac+iBv+gk6m93
bJhMu1JT+eBmsMn8STrtMtnOjE+YNh5yLQrHsm1M12gh3bsfo2hR0fVQp2t1GR2GIh8pHb5qGpld
ee2H5bBUmz52Tzb1dFxeiYQredIZJSfLTAV8s+FqqgSTNR67TvJM+e1FHTEIEVhkd5PctIIKy2nG
cbtjQzdxQKwJt544aQEPtSYmzieZJBQCbvXzxm5ohk4waJ5C83gNMqzcLN/6H7NZ7erQqEVG3Tus
EStCz2lOeNK3Q2G16ayLutzp/RqvkqOfGPCe2pidFPVYHg34oe1/a/tf+YaoMSLcCNcfQqupe4EQ
DqqW8wDJkjKUk6uxM5VftEOBxTUDhyVpcqrpQUQAGbo74nTOsFowpwaBb61HIEmjoYbVlf3jTDIz
xApCPv/s9zfgqpJ77lUeTFp2TMK1HUXfMSZh+sbiyiQmHJ+aJathPqDEu1X4M9j+diPzUY27fM3Z
CJv9lzspIiD9hVVjFCv0AuHxTGUMci2uxuc7U9k76VMZynYNOj1ZZ+EqyV5AXttS0NvB5+sQJFJi
h+kWbibha3EbrfJN+G7hi0xhXf4POqTdKIJyvTsGaU1EiE/cFIPYCC4aJVndWqqevrmnN5KdzZnB
NIIbJ5PPO6bvg4WiPysLuHDX2kpPVQQW3F/1bwAdZf2tdBoM9xkXq0EiEZmQeZ9iNn49JMX2Aj4Y
ZtzS4GOj7/KRhbFHSnC8cARxnX1lDU+CV88TeFrGazXZT2AFdpVgVQ2cb5/oJcjnrffQ8o1u9rJK
l10yDIhwiDUWk+/eutyQ/TuoDXnKDpVmHpSPAlloE5TwovuqJqUYMtLM63il8bo7Dx9M1vaInkMS
o4w6+BUh5qPk4Cbcw7GY3dT4AToV2NnHhRhEyS4mFkVXffZr3e1QNcOEPi+ApTAd4l2jPozyjmoM
vsOmhgkOXMvihEuJdf+INSgUNpW6B6rEtVmRTafDc1WIyQRx416LTEJlIYnQPkIMIDw86Kz23aC6
fybCnyLjen93AexYDU4/qMqiowISU8q7UFtx7Y0TlTCBUTBWsKhgZOPwrEpNGuHsuq9CQIz3PGoY
gwZYdjdFZ1WW5dA74swkSB2/Gy5IGMl00lZMYHcIgEcXT6WrX1UyZddJIh4Fow9Zc/o5rgKMOmnG
IFGA/F9XuBEUdySF/Qn6gQPww7GA2O3HJKbqZe99jsFTO52HTnOU+ciypMYs0xmzT4YGBSUogPE/
qde2C7bSNTV8MbYFweqAw27V22fu6Mbn4MQuZQ3Gi+iimN8t77tR3dw/baFgdZxkKJc08GZpUOXK
QAWH+54cba9Rb3JMBSHMJAF0PqJklq1Se5fl2NfgUHRvUa254xrlyJOyvM6HjDfP2IFnsUB+tC2C
9/nOmkGLKoMUG2ojRzSflK0dUUwLZDl5VU7A1cOh7t/iAt3kLkoS7eKAfSV3uj6F9H2SxKsyXVfe
bTqL6Cpvhrx/qGU6+ixNAhzc9ohQJjrjto0WQPbK3n5Vhy9i0aV6eTBhyuocvJYs2jrcgV5f3kDU
Mgj7X+V4UcIJIFu1T1C949Zgiy6ylt+fHhGzkqDJ9QF24eYQLUbyHZVa9Vg5CT6pENeXrZHEcSWH
SXw1X8HlT6jwJKF5Cw6P7RdwkkBz4msgZFKjLK/R6Ah1do47IdEbJnSvoi2IV9zxoRzkLkKmygWN
5Pip23q8KNxfOURKqRnvt/MvrRArE5Omyj3KW+hVm11EDsTYKgoXfkkLqM9/sR98L00IdJFMoPy6
VTNB1QCkI6+6/ZDf/9lWR5QzmbHrMmH10txugwTwLxCa4nUr6XSeOPG3OIcAWnv06zA+7tp/wXXs
l22XXeDkNtVqqJqsDpr4iqPE3ylmXPA1Rk+EJzstofTMc3eq3KIS85u86K6Gw+/tNyNy7tOYBH0r
vuKOGGAv/JxLohDsk32Cmwy0BpPpyY1RzN9KttLrpyPVxYvXGeeQ3IosXJ21NshdlRkdmu/6tYeg
Tsb1u5/+O+ns3f55J4fAj8lNgHnQi8D4M4dxju61rPp4jrTbyTBTtKF/W4oEa7wZ6R0jblUXu0O2
Tw4w9AN7w1vSH/PSsQw6jfltEagxKM6fejBKWTuAXuEqp1fpyjo3cAkSAlxVc5mnf4moNbKOO9ZY
M9E5VroionDw/XFHISF9M8JT5Kb2K05KW4CkB92SOeb3SqlNQCTFppxBotaRP8RYgWsBUMwlcv1J
o9fUe7DB9f9k4BvjCyB1E2bYTUlHunB/ey7ozoJIRpPKUYS4asZOcSSZAGQ38mipUAf7TH1KujG/
BaWtixl49cvzZCOkR1rcf3ZDZ/gH74SlUGSchzmXSbCXp6bJ/eGZAwjb5DdBnMU4U6ThTIAVwOQF
sTxQRIJlGbWCe/wYd7ml3FpTv6CahFVfLk4uakPAKNB59nV/Wp44ct4hBFF6rMtlEiD/B3sfyV6b
2ASDChMvqKH6oG+tglCzzTIdGxHYwU83tzu2st46h8u4a1qM7SiAFo9ntlnWBjCTNjZ4sGOgAl/c
skufbhTjcY1WhpmNvD4ulOJdLY5HUrp2bhZkaVivJ3c/SlW7J4XkUJT+oGK9xmh+lnn8EcstEw3m
ZYPf5LM5gfFD6PcXPqdx83+zV9/RInd4on5j95WrqQwfooLiAif6RCSDe/0PmTfrXW5T3nhVercl
ihwDeO+vPKlXmIkcQaQrt3f5s67zaVcvkreNxJwtO5DSGqLMqo146ndCVbarKJFxOSxB979Qel7S
W01iKjQdWnyZnG8f2hhL6FY9OV2u1LgnhZWv9TkY5TKbCRnkigYwGV8Zno1z3WzHcm6ABvt3zh1c
Qv9KESAe2/HCIlEIthoN6yK6zE42oWNGvm1GeRta4BHwzsSXT+8EphxBNxhiIXjHXu8u7PMWoU2Y
VgV5+R5k4nvR5T1uUZ1Vxhhn5vWfoe7bav+E2uO7epzMFZ1xnstgTL1AL+ZTry6z/eaHO00K9M0I
jTql7Alh79NJiGQAXplK1+VCvRJDk9uyTI9eHz7Ucpbfzvx8en0/JUgLjOat+M5JN4uun1whmEep
1I8IMt4SyvCp7ErPpOZ364pJtAumfepIrEBu1yByGeNDovjLlIr/+Em/bYcy5uS+r0LP1PCJ+kml
2wd1mvnRh9PVLFgxf2Cpjzp4S0yKzcVRDML/tkly7GuHbN3Nyb4KVCSQj8txakcWvusgid2OYOsA
jg6XiLLEQERXPEMoSQw1njBXPWlU9aYpASir64xnMN7mWHdyakVeBxzawJGvJZ5iCgImhaZ6P8bG
GsWWd2MJQBFpmfCCIQDYFIXNe1n2cGneU0rToiU+a7gLdBAUfwvtqvPPIdWCdCGh+G1b7+OndX6t
oJr+xa9LB1zdwfm+0LvjZukrCl5Vo1bhqFoqwi5g3t9c/TdUHw7gj2YdX5WV12zzNfrUNd2yNkKb
WH6DL/eBpNG0vQfMzFGjDbMu6wqZlbupLIMO1GCyqrFyEyg8rl4/LDrrMXfRj4R23Nm+nSlArB+d
YliRGWu7jgg+uyRFOQvl7xBPyycoAcCUAoMoSdmxMKztBdRvzFbaPQtGFnJqJ6r/3W2QbZsPb20E
dBPD+k0bPL02nM10blHu7kqll755oOZ2g9+uJ8PZYPczjdk/SUsU8ki4VoU82wgpsamHjjPClg2j
RiyiIEh//EskGMZPoIBzngdKmNX+VEXbJmkU8tytzQDP2qLtq68eg79HZvVAW+XNpm68iZ+w2OGI
fd/h8xKIwAw/CViRKqFDFCU+rcYsV9Os6Vb5Ig3q0nKIM577L9jby5WfMdEa0sx6Xegtr1kAlabQ
+9SHtVVxJfNBibUQRy5qq1y3F6/S9b93SvTMdIqS94M3I3LhZFtOxp2zIEXC2/lKETFVTVTMWpd3
YFpLuyP9c/GRCR0zO+RnjAbQ1lrjH//oLuGz8MvHb1HKIXU8aKMTcmDPfQVLV2WLjHnw9av3Jxge
rxEY4mzj6i3ow3wJP5HaotugfeDFF+BsIln9ML6vuXkZA7Mmys8EHqLx49YSh2PewnRI01wjfK+5
I+xdmRwsV5gI3o/nqmKzQiF/jCSC+pL+4lBcCh5v8wtFj5oVj9EfZWiI6hfn6TzGvLiK8JqyWfoU
ehY58pRNjV5rCWyCmIHtObkefs2PKMa23nL89ADVoZzCHjk7Su6NOeKLVG92xT7chwy5wt6mn+tr
/1Eb0PiMgHgDg4bncseNhMvRSdtajkniTkwmqTIEMip7N2dpZOHXijGx3wLyfANyYyJGLRPYD7pi
/voXHebskxAzqeC01f+rWjkLol/emOlHj5zW6RfnPT1pGD4dL7/37hDYV6lpQGUxIGzfJNN3kxaD
oXMiPdTgm5ZYxb2beOFYD9xTL0cWNBcLof56x9qZz5ErjG/jK9SkXRMEhG7C+/H3U1zGutlbB1hd
vmYviZSKvvdQi2vFiwOk3IC1x5BwQXoYO44+JogQT7FFK/sLpAPW+9WKK68pY+e0A9iQvfvdyHE6
X8/NdsU2UOKfinhfHhvGrXAmTkZZ3gKfwhhICNvF2PuiJ79RQ39ja9r3ZYHeeQHX4iNvvhkOkFFl
vG/PLLKjSvYNwlTfI2eCqzQuF8WZCEUNCBPQyds53yjZUTifjjUpKLzzPlAh7Z9GpRqagTep1+Yr
fQR2LzfEFd2iMiV/GiO2bUP1gIOPOOIDIHT2Rpa8hhNrRX1CY9bDIkNU5KEWl2P86hBhSZlM9po+
GFOMYeltcOtRNWubWZ/8HqBu0aDrBp65qR0g39Jrv4nVRv7cvtnjYLPFvxg+66SZrvKTbZVGBJM6
SYX58M/xo8gDVptO4EWqGO85FqY1OEDfSB9sAZ/9TiIeBUtQlfjELv+vs2I05DaLLwK21/X/Iqr5
tHNkbWU2yBFyTuTC2HP23tenISIs8w3lOLh3/Q5VwVB7192fJeV27E/Ic32cF0322FYs7Bmy0430
kqvS4SZp2+UqUYy9HunEHU0ZZf085rMQ1imYQ7H7hdQlS9/pp+DeBFol0zvon40kTnjubuuemU81
/jyjBMkCmeJL9hVSa9egLo8zIOReJ6KBfo2vHR88ps0g558JygTBo69oW0zIp+GnTyGswmRdzWPH
vCV5KhFkXV8e4TDAZc1DVlYIz4E08r5BkEKvR8QrCdgePfbdORYq6oqpP8/PmIvbr3Kb7cYsTeGq
H+p/CYgJP6DVpeFrHsb0JqchIGRdNhUD5ddwZDH3KQ26z5kVDxVTuHQLRlqtnLY96RfrWEz1d96T
C8kHY2DnnuEERz1c0YDQ4fnkw8mC5NFpXbNmGOFONTOYiBDSJZVuHGrXkd3PEKbC43afm5JxHkea
1JXR83/EzGS35CyQWna25tachUD6njBOZsvE+ajqfSzcMhF8Cxv+OmPmnFcmV3KDBHEFHyvx6iNE
rhvEEuuuZ6gJOnj5hZaRPTPOFp5Fxw9tbipSO/GlNLSo/jA2DbLYX9RWC3LXGqzeE/oUcNxVL4j0
IuMvTMmJT7ghEXp6+k/I4FhQczsObq4wKMYjrYDkKa8cTR+TJLYMFIh+cWwWz3xFK4fIlP4O0weW
gu1sLndINWZioBR0mNUOgojr4E5/Dwevstq4vpbU9MqP9sbfPePd95tD6HYKUveHMHHxpNLYhkxf
L5AIlDSlJq2BHfhxvVYjTfoxKsncz2AF+JqJ93P3bVPF0JSH9hXK4mS6xlO0298sTWfsyzDdivZr
U0jfnDqIjYKBqZFRyOg3bmyWAcl1bGaoRtibC5RVrXtMvTUHxN3gEyNs3tCx8AuQoL5NI/7Vvo88
37C5ML4ITQNDH1T1uZqQMvh8VPrkPHzscQnzU6GIR5TQ8K0vIsLnU4ICLTMTGVYvPSx99cWdhDwJ
5tdtVGUhS5oQtjczugYbBZ/9+WqtsDkJb7R/cQlivL5Z9jGQ5ZucljqjG2mYnJI1IlXG3BmqRGf1
e3umACnzsDajc228qI5T6s5c91DC5Uun5jwjcrRqQ22UpI4xVihdn0K6VveBs4kK1WvH3aYqTZ+f
Vdd/w1goCiV4KyZSxzIgEfD3rv57w1j+tDB81bKLX04c5oQCqJPn0+kMglfio2swC3bVqaR9qDO1
AO2ZjESKZ/OFy+cnvM/PrdS1ggMd99+4uB9jUzyBC0i4eYLNQ2oHRGRNj4KDTCa/QUraTTGWBv4Q
f6lFsAwYM4Jf23g2E3qjCOhNhuZbIs/StLUZaIUl3xL6EShDviBVii5lu5cUHZUu6J8Ourvbx0m5
I44dE7CHCPe8o6ULOLyJpY72cNbGxfC6K9NSIwRFbyw4eAM3q/T4xoI05Gpxw0kRmKHdoiQNpxtM
FkM3f1ToRW6R2aqB0D34vII/eEHL3EhPP5IL29BkXZTJz47VwsS285HRru+JBTEFPUa87FF6gDtX
VRFqJ7DV1VTRFaNb+Mgfs5aI6Rjl4elC94mJ8JfdR17+P5Y9F+vD7gUzFV+aUd735g+wDED4RYy5
7kC5xyqD8Xzslh9p3OqheaH/wZgxYu8a2wWa/BmwEAcNpoDxu6A7UDk7uDaMUCbzsuRCZDRZ4W6L
434oIFT/8K7c1FecrzNHFeanJBdwX944ENWrPc2k8UQf9jbvbu5ervYZJL7BafMYwP3UmYG7dKKl
6ahlwRG4DeMyeB7JKv9YWUqIIjnWe+iQRKLh0wQmk49fHsQYB2d6kbETaSqIGmOrDIbcV+xyYAt/
mc8g7KQ7b+EovUtdwIl65c0/3oOvaszr7C+CNsRx2wT58f9FP+c+xChI+xzDp8bdPeoilJxBAra+
aj9hNL3Okc+UQHZOCjKgr2FEFcVDfKxj0Lr8yf4DFXkmzueDeOJLsWCyU+FM8K8jSGAL+de2PccH
v09j+4IZKxDxeiYui8dyTk8ko/jAb2UfIrvOi9c/VFU9+H3CEvaLWhTVCZ4V6F8bs3h7XbQbHis5
Z4l+KJYhemSgj0uXgDZInQK11UKkDViifrWGTax3gGMoI1asMSX00aUSF6+o1AgwvmFC2CVZnNBk
rfZcOEpcGWJnIKtMG6j//vCpPvBXG4KavDdB2C5OfUhQ1HYZE3bXuPSLg1fdl9+/3AdhagQOm3Op
ZjKVc3hGIPfIy4CSuyhkiEgbKFxQJf7IlvXSlIdf/CV50Xshlh49c/7U92vwd1W0PabjUpn6lCKP
TJpOQcB6d7Yc0yF1qvx8CFDft1JhyMkiGKqMCPWRXFiJS/prj+LFSy1+IZrgD44vmN8apk36w8iA
NieH+c016UUW9k/qpwRISX+aupF9ktO/S0t4rgmDlqp6EKzZ4B8Wfr0TPIlV6n9trxO4i4ylK4sj
eFeHrIPc1uiG0wXr0SZz1iKX9CY+oF8jUMxhlCJnRojvF1SDjh5358nQozfv+CC8QoHJjifXXofk
VggLKHePMnmQLypXYAgJ8uJl4gQRnFdMsUABQ3q042nz+es0BZTsPxLYnHmjeFn1PHyTGjcBTjmz
B60zCAbGMnakwwBRilTGISuVrw5hXjsWxDcP74NhvEMqtXfRXIuw58SvwRberQY3Z3O3xVF1Hu1R
fpRL5QwHO/aS4Y70t82pyjGlzdlZyIHGAwVeh4Xu1xcAQ/gkUaLzSNt0qtUORQkk6x6B1RbdBTOj
UBhFWWBy6m7FVxd6h/7PdB9YWC/53f9EPVhfWxeYw18U6uyclP+jmLkb4adqvYs47o/cMd88/vSW
RSRmtDFooZKd6Sq2J7Jfss5YRH+KAROeI9Oq1o8t7SlcUtyQun29OaE4vtUaSp8iOUFhNcTQehlo
oIpuKp27JkM8Yt00ddbkzwaMTod7pVYsHyxfSt8qEBhZ8jeODqyLHYp/tX3AViaUW98Ba3FkItf1
4RngLLi+QUKg+9DzFE0lv87NMpUvJFgnm97KbJx8dHX8HGg5Ztu854acDVJgjqxuIPrtA8vOLiBw
0Vv5Ci3SWlAs0ron+nh2x6grI8fg2IclpkMtIvl9deZeloBGDUcraq4ChnKTXIIFJXxYCUMpvO9r
Uvc+qvBwMBTyGeDbqsr0CgNx3uNmSdSwB1CSVYyPi/RZ0NvJRgWW16fZm2moMS3iJsFfq3WYqA/E
iqFSLDs4vbNEBAthL3+9tsQCese1pPpPLIG5QceaP3gSPUk0sn+6U9C5gJ238eLetPlgcXA8QVDV
N0tvPMET3ux/H0wE0tnaDMjRHLCwkcEdP71aigbztRV5TtQ4e/dKQtundQop5bW+c2Yug3cICqzK
euwHqcVrNg10NzjEYPMInUl2VGLawIytMgVk44NDt1xr9mMjFgm+JO9Se+Z5NuM4+wULFkB/ZOnR
plP1L4Z0CN0ZPppjKKyWtOPA+yyz9XCrzh7PIg/82CU5ec2fIUK/6taLbfQN4Vcp9N1SFs5aGsVX
rYAOHNbi5xpOGaPvsJjwUHl7DB4oRbcuwvGnuEGy3R230CvF2m8BOX6d2BsR7gR+WtsqlVDTH8yb
pawtB5IxXaRyjUYg25r+Ka0Gu0mQ+mVXQh5lptwLC5zd9zGsvdsW9Y+83Ih0u8pFbT6FaR8MezE7
wjf4DiAKvhurAVAHFDsG84HicKqg3P2dSI4njmZXOs7RxMMYckKciS7bS5EbaoIHyK4MYHrZ/K7O
0DZHyHGmJIdry8wQCiuF4nUD+/FA4a9UC3qqzZ2pGNYiXzV+d1JRvyG3TV46yYYpn+ILkBumP/lS
yhtLjWEFeGVlG5Zhvg5do0EDTK24+BPaNU3eGYUvsW+i2DOJURlAODDJ3rpg0QJYnqiYvxA4Vyum
ZVqrJpH/1pbm7IzUd6SzfSOgWkcbMa87FU9gkaLnKn/9hjDbZjYTByxtCt0XLltYj4RXfv4V/hB9
ciVROLQGcUhVrd9iw4eCh5Z/cIbQ2ehXYG6FEiBRiUqLvCt0ctFwAkuug0yiwJepg0DiOCqnBTjc
4y6ksxPywjpL0rwOd7T+Pik15MhhGa9o5GomLO1/cU5nZimZr9mLCO5jDJGCfRQ/a+aK2MLzMUNq
/i35j3Eyxru3P5/Q0U54ApFXevF3HHn1Wn3Nl82ICTNZEtBVGh74JRklqxfxdz2zOUx9QxpXq73n
xE6D5vfn/JVWlE/mbD9+6aANzH+IqLrjiEinp6AU2/oZXkD0Vqg23aR8TDSUqbJyCsQX8TYvIg9t
EJXTwxNYUQDR8DQj45wyfRGFRfwMzk/J/MtmBa2Za29/hLH+tbiBddanyG88isVihRPNUa8yOUKj
3znSbx2eUj9dEIE9/jsinSoLlPD1yIdWUFV0OJocFl4KB07KGS9a74NLPj+DGbzUIm1VTMKGQJJZ
hnPK5c97xQoVXF6SNxwlS0gaNDFNK9apM2WnJHrB5pYDNyRaPEsre7OebytWiT2AuIGddqWbUCrA
EcnkXJPZFk785lQts5YtjjEzfkA2c/tGaRPuvRGDVKWuw2GyR2G4x9s+zOo58U/jmlrbIIAnBRww
TV3ecnY46zZ5RwpFzxFAOtnFZ8Lo6tDOkeISYwgo3idIKLPVjKZF0jWon30OMlDd2qqxDpfjTE/z
puGmP8xrkudsP/eqhuUJCP+pcEua/Do7DyCKw5B5T7Q0UmVcnpBJGMala+CuKfepSRxshxTbVHAX
kP/QKdVSoUKGGPZgPAdjNn7ARXxZ8sIzfYOJroFzldfU1wA2rRhKG+D1Ev7Ei5UPpo5iBxiublOA
S8l1nu43dZFtyg/K0TAc9hPswBWRSukDul8KNJLQ9XA7ZHLwvuWQTliz972YVRAvbSlQMS3FG1Cr
B5zfWfBHMIFEYvgC86oSmE537BMERMy3iueUCfZfhOtxMh0KEnZwFoMjl/Mt4vX4MBKk/RI2/xwT
3QLQu23I18fN12PvsJhC+7AifY7z0XOuSQHS2GUlIYTf976A6CCPAASNz+7Gm7M3A8nFLG+zltPl
bTYv++hI1eoynivDeIjtxhnEhU7v6nIfr8q74zY/s23c7/e4m1FdqQjoZAZExNZiEaVnYWLgtnan
CG6ncljLWlMPdRrxa4aRzEhGC4qLrMQeOA/YJTXEE5IhyxZqz2KiJto5IVdhzclgPGTAgYXul8C6
41rGNOVzUxrF0+qXMs3foMzPChvRgk8RQr0AoFYPAJwCefeUy8JUwN2bMwQCnhR/psYnkRHV7dkV
/9izX9Z7OEzZ6MNiGTbiPWI4Ze/jISVUJoGOwef9vdhZXinPFkPywm1pOUDfjhofMp+xsF2Gx98y
wyfKfRt1P9eJRHLR+5Q6LZMxqWebBaj6M9KBA1cnZ4Ery2KHAbX/63dMSSSo7M/hT0UzFv+hdhbU
abQTjz5gcvSjPG5+7zFkrxMOaPIZmhdP8FwRnH/UrQuEnwfS9pbtGGwEz8exB5ruFbaTycQ5m2FO
CAqvYuPVV94WZcbwFCUZuLchE7m4fU0ggypf7q/mwq7xJ6J449s7sSWKcx+iucTH1yJoFkfnG+Vh
a4UDer3N7DoeV1M1WnV3YT8AoSj3b62n+DfWBtYSmJAVoG8ZgCI2pl5FoTkbLZLEvd5iFf9i2abg
t5oHGR0tYpvd1ND9RKNTcTSvIWsUr03IcLZp5/2/PJJiRbqg4kFcmTUCGh6cZ/O8FTQytAETlDEq
+VJ8tn/5z7OyrkD4Qv9Lk19WQIgufuXRz7d/abTeegasbAXWcdOd34oKAeGlzJ63ad/3fWkW/Gl8
Wq622EnkPKmhEyfv6wyaqcjhoDQB+PTFvPLq7zaP6WmSGm+k66o4rNkvfJP9ElCQJ5pRkWlCOkZA
eNBvh5sfnJHwtOkHX6CKgyA3pySHdpzNPT+QmCtiA/aTHWQzE6gXpdAEjUyL1zXSgBIpI7yAvi1y
oXSn9zTr9d3VDGc1+6PIDuJpybHPFjLlg9P7XmQrIApHJBRZOY1VThEyS7LCHx6/PbaMcsSPaRdC
feaFqT+XAOWCc2LJzuGNU0uVVmCLvwYUgAjO7UjTo4uRUYZlrJ8P4LBKIR0w5reXIptPfAvtLRRE
KoOPoFB0WftQKPBd+HoPMTNT/XVnQtYzzesj2q1qoY4cKY0OXoAupv7bB+Qmnqnh48qLfeLjjq4/
+EcjEwAVgxIpPd9KnAdDl50briwoEryPKtlmP9LMkZm6g7TF/bmZT0Rug2+NjxZvlVT2+6Ao9DzH
CWN/XyXMz6lTr6j6wo3pgbbsjHqaZ22feOsjG9gIwipGbDF6FkO/X7mAhlFqoJpA0GIDwm8XCp6b
vE8uB+coIz9B7+u6aE8x21PwD5UT/Ib1C4IZkTJqYIO36buHe2+fJLOnSg+poE9KdTIE4nxK6sni
XMhLBcP+l9k90nl9BaDdbnJEtc5ffpANaSgdWtKhRKiv2wVoc272zfGqKghP1Sara68fBQ2471lz
3i6iK5kRZY0pw/Wg3Pkz+bme+3Zn4FEW2GpFkvcOU8ths5ayMCQLVyzjUpNCr0NedQamcUzMC1yM
tAja/6TfL2YIARYVQtOEM5XL3pS3/6k3Z2Q+qEJ/wEzgv3M7CxKcIVu5PBJHZiIyhC7utcpD9YJm
SM47X55HWATIEkB98fEled7QfMase//0sUGtfaGR6IwERVT9MHjund4s4xc1nR30inTPSr1/C6b2
dNoWaR6UXVmhOc6+mASDNQvnHj1vdCY150j30I9XCdegAsgdPTGQn641aneM2uGkqWY8MrIMO7dd
56GWZ3GcHJswzn9kqITZ3cPg2KJWym4Ko/SNI7MJXqqEzDuuvzzMnM0zybV3BWD7OjAPRdGIXV35
pOouHc1jNztgblQUfcIf5ZOXlZMDS2YxV9hf9867EPwRlJKQ4htXEDOi0hXPgcY1stiiyzN2QnEb
8e73EwyXY5D93Vr3fPATx79LIoZwIqcnvl6EEuorr4o8sx1dJQNn/2CjO5n1knY7IifmFpN/pQJk
oxFaFFPo5sjS2AOVO0e1HHYvqhtkPkUY2Wk77r/Q07Oyo9cwweq8cP79G3z2lzPOvq5H2+FyqzQA
CGE8bOUHzDoiZalw+kp/74HOntaD7+BLQbsgfw51mOmgycP/5FASLUWAmjZom8qLBNYaQ3iqSGte
9O3kCGZz+jnfB3mgD+QI+T2GkKcWFiOOULasub1dLNgkIqiXUFaEUdmlrgJSEaykZjH19AFnXvnb
N4Ix76oMwDncKrq4bE+onkvrWf9V6ptnFDNy4vR2ndKsU/gBlASEMJcbx1e6pdIP7JF9/LNHRD4c
hUQ/ROSYHQqcxodLsLEHy2hk/WYUF7IgP+IAYrg9V6zwrrzihsgsaAGi3vv3MX+t/Da0Cz7uhFMN
VCK1Y0ZUfD1VlVbXLKUDfcypNOtQfaqsiPhSGwxgN0XEfjE4pnhqrmjnJOxZ0bG1/eBzyAH+vZO0
fyPovjvF+w9mZ13NN8O80dYIpzTknZ12bDBmvoGM+52F2mjoqDKMDVNLZnojjWv3n8ApeE4AF5O+
aNj1mPK5sxyO/AjaJ5u8bpj+n/z2LTp3VrD9yOCV4K6uzdnomGrMusyjmez6eQJHBWugqVsKlVVp
75MbzVUPdnwrti88APu2yaC41XZa1RRcZbfR75Sa1BpcC1P/imcRSxWq/1nrDCi0coTz2ZwZ5gAt
JlzT+rWsEMElH/DJITD+jw2+8vCIIrJqNBhE8aM4VWyUNd0asnjsp7CuYEWPxHV64o3DEuT8/ciu
rlrlU1qhYql9QOU1c+ZQXysU/BaTn0XNQM4VxiP+IghQP9A0ctIsbTrWNB/XtQ6cDS0QKQgu1OnQ
hWm5JgQFsvFNo1UH/L/HQoTbJk8Ttjh1lRrlReTsYpGo+rvTYQNiTtWSfKRRDLgj1o8IOzvPCgsZ
wIRHxPmLhKwASGZo2vAbGY/sQb5YfgJ06GRbUSxNVuF9yXuK8YU3LlZACYIqNot+TuX/coGUUOsD
WxNHmtKf25RiJBIPAN6uhBgciuOvfqenOMmf1hajhRbSJnZKbXs5uwlKeZnGzJdbieQ7Njm+djCn
pD3bd2CZRdEOcpgOTHjNq1khQoP+QfWAXYLBmia1DIX8bkRqO2AdfoaQULXvo7mmvi/nC+2m0FjH
7s+FCwnmnBQbbdajnmd/2BN8MY0povp4xkfTTRCM8TXdW7/0Njj9spEbx+2r/5eYZSRyH05FXwP7
7gmi4/Z3TsDnDXCsphbZiex8jNTnuquVhHGsf004IEmZ+mlOMow7kX9+AzICyCSIWjSGTKydM0wc
GnxJtFH9eRTb6UNdxNChcaDHCpTD/URMLXUo9HNnafP6xIKFvh0gYuITiRSpEAI7mzZSpRMQBhTI
x/YumooeiW49AjApynbnrfGPtA0ZWzswRidIM8haC8gEDWO10hVRBlpM1NclujWnNqetmLjhKKUe
VAQXfrl1vLKt4fz/a2ikXCEk4pqyOMIJ5dkmACkXGXvrS/eK/xavNnW3FdD6SZ2TQbSXO0+Upeds
ZY21eHsB/ca0cTmxPscY+lvSQXVNRCJ0NpGgKOj46zPzH3+K8Q/4NshROzq2ECbM6l4+ayolXLZf
VtfGEyCZCLMk1hs27wFwDZHRXGXt3CF/9XZ8bxvExHtBl3VpvhiR6KyBCyxHuEAMQ+Ma6UPXJgRM
ITuh0Pl5UCZpK03KN8VztRF2WAoULG1Dho2UQUQXHAh+OfYpk78RkyvUfqG+7z33+PRHQvbzUmhO
5km9rs+XrSwNvsWr9Po+WcPlo+E0ZqY48VkHKQgTawS+qbYYQjybNjQvmPaTQ5RVgd2I2BtKOzu0
URYhapIst+kIBfCcmkcWxkKa/6EPWXZmyG19tBHgycqIPpCXn6JqnmU3Kin3VMm4reKIo39bJH1n
zgOIJT1bV+GDjC+VKSS6LwxFuNzs3t5uKnXVdKhVtQEipcbIcGLkJBu3mlI4ueOaDCKmJ2TqOuKw
dTMEMH4KURNHvyOvv7B4YxvWFFI+zUzzIP7Hmkswvy18jt1oOv0WAtW0D8bxnMP8fTHN0K/mAaEN
tAmTfaFlY4kiYm+qcN82yLOT2br0B3uc40Ou7acYoocrYdNBkrI8kNQ7ic6U7U18F7YgiELeFs/g
tNk/1rCjeZXUvF4VQm5/lhxfLIqtFGUilW5ctvuAX/GLPsIVS/dLrBQxIwmrTSo1CRqY4NtZExJW
2rXgWR8PJymijbGKG51XkqVQRRvdIhVnYBgnMMQw66AhPi05DifAQIvoCj0pv3LXdFBrHoTMYygy
j8JX43yo03GerLcP6P8YKfMKXhgs4hd1kwMnRQtPUKWskNuXNQ366enuykGh9Bh3/1KYivG6xQVS
bkhfHMsal358JYLaYExyjD3YRc9WPtQJbjomFugDlpw+0ygA2wq/ENgGD9UkeNeZmzEoP171yQe0
dPJoftLcxak/7xtB2ypXtl/JL44XkpiuYuGsSUQjpsiCKgKJUJS/ZG94BgiI54b9evpKT9H6OP8v
2x6LFo6tk1k0JLNKX68IC9TSIqUb5FOtH5jNgWtcxeCM77mFvzNJzU4AbtYNsNN5dWrwSIb9oBom
9RA7v/8Fi14CmxaD7LPV4XkVOPkhLkiUBxHcCaOU2Jsco5H6MUmNjG0S+XTvcjo+pOCoSdTGEAWh
lxYj9LTr3hKRHLbh0pxQa3KtTaBwxnMLj5UUuz5B62L51X3FO+27zS9yMRE5vbugwFIVQPjhkghp
BeuRpBolpSTWOD+AxBa9kjSFRLAOuGrtXFH4btvjBKR0W2Go8eR69fR6asiZM2zwDmNXoG6ylbaO
vZyjvqs+ky492hMgc33WmhEiR+gEeLWioIXC7wTSmJmIOAkwSSyH+bfefieaHpqVpWrN+53+4ePo
Jztp0N4aeo+jNwTvvWqJOcHGWqk5QIKHrWls+/jeC3RaRdz41eN5t3RQoFjITdlKPvvgP+9IJLSs
9CxqA6zg9QrHzSVdVnVIkFwrrPLCV9U2NTXyBhCveY8zaQ2PoRrks9k6QW4yDAtPoiKH3U1cdd8Y
IpMWPN0tSQ3RPZTF7x/lrL+sN3kAsYoC5iTV2E5HabhiedJpClbl2bmXy1RFYhCRHWXw1NlPLKyU
PAohU/LAD+lkd3yGlEnzJrC3Oc2eVMqSraBAm+qJyPGHGVUJkiMi4agArq4RRWy3T2dvbik9hVl/
YGDopgnVyuZ9liL75u5b8I5OXB96L2rytGD/7QUlVp+c1zzdgSLykTZG1FlLZLz2B79Tgzeeu9lh
3XMzCzUZH18h1bVBRi6e68fMvwpZlckE6eP0WWx6JTtnfyEImJjQsrydUjsk38UtW+SCv5Y2axEw
V+9HRv6QNrSQOWyqcIMQW+LGH6QBkIOgeWcsp7xKlPqglL0R/4ZNrg25p75dgtrKyM6Z0JxWk3wj
aTxWnK1N5Be3pIUD5bTuHISHRD794itu7Y2NINf4X5zPp66ExNcocDzBh/G3RcIoxxXewvWQubNl
Hgk4KB7PzX6RiPeo1SBvvAxEReCvseeFiWtFR0DpnY/W3Upn4cpyc+WF++qmkP+eOftnjeVM9t3j
JWxFcTAzThwD6VZ81LUSEBK/wKb7OUsDMOek5PDizJLmq0jAIi9uDgzrh4Q+YXTfSSZpP5/0oMA7
EdlX2SCh0DfdukhvVTh37mZrjOhx4BtUA8bndei6rxUin7V6WTncXz7qvZDcAU9gAvwmhs7b/ARy
4+Ae0MJdO/1hdjzcakJXpba7vmYTE3Q7gfhRm2ZOEyxNrNLPjpoFkS6o4Hos2KRp3VRhaVqCXGE5
rWBehC5JSJNahpNMs4fP0+yoiqk4gFaoLkBuicMdOmNbCz3N0MgT+ztncuvReBJ31fT/HG9Yr1dG
O+O8rWedYWKxqGBn+y42Jj9M0rGnVje6x+Gg0aLHB54hH5zXzT3s7Z/OGEarTSDAqcWI2ATciQNG
uHP7uOZTVt/YHBhLUYC1EbZhylZ3iEqJHyYPXEiYkjRWQiIrUb6PG1586YIm21WoMIn3N0B+5/+W
jnMGbNamQPiHdysWG/aSYHwafdqdwAukvFxovpIg74zCwYuo2m1EJMWidzjXBaMlbi47HDKXQHt+
C3ZvjgTqaCIiY+Cc3+8/avAgxdR4YvQKg/fEHPLjnJAicD+Te7EEEBxbg/HVwKJJ+G6nMN9hRU/q
+NcVrkUeiI6Vh+6rZnwymIUABANOugZqPtJmCY40exGyJZFSZ9jYICD7kfAv+wHm2XuC11IbVn1t
rHAWKLSi6eOsKaohBslPZuFw83VWyubT3tE60T/wykTiAaOtrwz995o2dZPpnkwZqOYGSwAgelNN
Gh80+DF3JZz9x8ch8uf9si+w39EY39Atk6IJYVv1lwCqgpKqJJiLtqgIK9IKWfhzQBIA0if8A2Ab
J5H0tCBXFnhtqGTAXGstQ851m89lM2jBnWCGVgsLjGeeJAw++cM0oSn50qKvlXW8+YLlq+G7N5K1
NZ/LibavUOsaYVveOLWH/3JJ+tMKy2QvOwbMAHCKORN6raJCqtFrLKwcoS5Hwxx2b2mnrJ5uD3ld
FnIlg0ZXIN7iLrIFxkpNKdvSdn+zkYrC0fZBQVHVRb09dzH7ubHKKfKMJ15Qy5EXxMZ2HHsoRnLh
l7J4d1GrHjh3/+ofxqvP4IEETuLfes5SmYT5p1/TqldRhL5xt0rwe3vEWGQj4oTBivyFodniWZII
8aXNUDVsd7oPRqpqL/sOk+aVGF3yeXY//kqTcGLbvINQSHS9R/ngO0XSKscZJUvxUXNvwGDs/Pe4
EZjVw2HrH/nmk9vBYE6wf7nGaCDgIwmR20GqdTYc05k11NtMb1/Wt7B9jtpZTOMtGsWlUZofYxXj
thQ9++dsN3g2KPXZb9J/2l+MJUeAEO7RiOmoGC4QpeM0OjFjxs+rtsdyc+3xfTEizltdyJ0uQVPZ
H35qnyw6Vk+zrBpQV5tuiXV+CzZ6Us3ay1pbo5lnm3GPxaOuOsionYV/stNs/KrkJqxoC+PMPtpE
WG9lJk/pdeHlx00EycgCu4RluwwUwdrwcLveLL/AVHtlK6pU4L/sSUicEHJBO1J+Ib8r35ijmbvT
9GeCb6BbJ+hdzz6GOVRAIWTbXBWO+lW97SlyB3HlT48Srl99ex2xLI7/RBhdpmuutJrmoRu/Tko/
CSTKEtQJKuKaOXNdUzmLZkiKFcrMkEhngpOmifGbi/y1oFWtAxQQiV8O+jF2Kak0wbDhNzWp2sWP
ATmnZIykKeXqud9GxVXtPEkSSgwgmZs8syv7XsFtzbh7kN+TQVv7A39+nWXKKM0t0EB1YgrGRskR
3NwZ6qZUMypUnBLuAko2jvzdCccLX2y7fFg6Mmm1A7Ap9ipexaarEb9wNN+a/kc/OU73kkRt0V/1
Gm4vAPbUDazi2MLUIRsjHy3nW1PlsUO+MeqOHzqXT2jM8JWAzZ0wxHeRKFTujCqGvQbKP0lZdSZP
HqiOgrfKRzvCaNsPgK/SH+RycU2zLVc3RNfWD4r8AyE94pxk3EvrWE4wXHcqnlAdQPCB/yVEK5PE
gsYlkrKptQQZpgvh5wjFEjWGMBiHwV0KgpM0mcpFMMyHjLHW56BHne19ByduonNoaVSJ0jclFsY4
zHrUivph3kzZP2cLyiRF6dp31Lr2dINJtHCksaSMAiSwvkAi7NQ1fKvCk7HtTzEdI+vwQ7rRZAVo
N4SVaL39IcQbvUW1Pe7bjpO3yweZm9QLZBYh9hVIzxPgoBAh+/gC3caKHPPylqKcHOPGIU1iYvFR
BLJwXWvHpu4CHSqpeseiOFCfqIZJDMNjLd5+ocdHNLtH8JvZMv48O2sFfHiTSx6SYQh8q28S4LD9
bInGaS2WtFxlnx6iAiz/fyBRnKXRh/0Y1lQ+Tgtr6vFivsEjV6Y3ffyGU0WTJ44vsbILKvjjvZ4p
OWW/qajatvJlOufvQWocASZQi/4+T6ApJTEjBPsa3K3XPsEI8ZCsq2sEmnnBb7H8hsWq0eXNgquJ
FY9VnCBl+sgYDx4UvKb+tTo5wIlr2m9wTeJLo+Rz7xvZ8oPOCFCv+9A83/dKjPnDI6Cn7tcXGmT/
kC+hzQdLxe5fw/uM5wc6sQ76gFJ/d1hANCfMwE+JvUoKYbKpt7QTWgE342pgCXGkb5t7UnWQ0soZ
uTu6hE5C9OzFANNMJDZpiXtlKG2u0GvJjSIZmWCI9f4VpeRwvNjyqxLThZGTCO8bnF9iVK1fRpRw
x54IGK4DgcXYu0jwBhTivm0hz376wPp4OtDbj5k9qVbiooj7+o8w/wAB9Tyuqy1g5aNiSw0ln0fr
MUJuORHbQqHg88QxmDssDlqqJ0PI3DJXY1s15fg2E4IElkCe00HA7madwxiJsKR1vbdf1pcs84cD
pKO1mjIjOspG/t42yBHoB94+qE8F/NG8Cpm9sdFmdpuzuJfXQGqp/vZvlSTGEU3a4MbANxrWzXCR
ZL+hg52H0NXna1e7O1EbkwQVKnh9iZDh6hEgRpm+Ab5uwVPBgQu5o25EyAcV7NcWg+b3c0i/sxf8
F3NQxvp9l7ZRFFTNJDx3775ciA3E9zj4+SGLfey3r0/vIQMcymLhBMukBieaQFmKWAREQ5qGcOBT
rcvuyhTTPTSyizJy+WUECQIvFOCHf8kEuOdJNw5B+NXDhE1S6eP54ysU5f1fcQ/3jUgtEclenIt3
YVLM4NbNB8bZWoCMKSruJtk0nABo/3A+oJN0dcdJ/Ni7Wnx+aYHoI3ervqnOxjMmqCBFkBRm6eue
Zs11d4Q/LRaqgO3pH+GuRFlXkiVLv/rdrzdLy7sT0XIQwokpCZmWtYUScudeBx/UiywopHz7aHTG
vcdbvhE/RtclXi0BDR0hc0MVIJ7YBgwMqvxeFdc9PMy51wgax9s6I5cptr57nouF66RD7NlTkzhw
5gPDjJ1nRUoEDT6m6PUt1UY4zw0Ukhvzd9Es/6b1Ao6fK0AkxRi1ZSjT1pd3Omj/w9nx/yxPmugU
Aqh/ZT0qDKkC4O7gePA4tVZR/AgGYYvG81T118LJ0fWUja9PuX2c2dsAPyjI3bM/qQV65kJwdv+l
UB/0F24FqY1HqFxiv9BexXFOfqXTjCUuOKXKPTJvT3C5oZTMLT+TE8bB75Fj9aNzyiWdTZDD2sr8
IgBUbD5tRE++zMANNMZEEYYPpJTZLrEkr8cLcqW4GewvLzM5DYMwV55skRN+qUih/NlgKrvkeIk4
xIoZEHV6HsSkWIp9Bc0Xzn+eyesTCwpBQ/UXhKU+PxA9pwk7s80LrxBI4rZpf8+f9mbooYC7W87e
SDZM1yPxBZTEQwdb4SJAeL6fegANePNOHCWXmFdWyZZKaCQlu92+F9vQcU2wy+vqj8Rq4wtDVQdQ
HNuCpTgltLo6U8CdItVi8iflx2691ElDQnCO6YqHcP9xueaUIYtiHRwPgAk0WwWLr76aA7QfFqz1
eMr2Ie4ONpcFBwjxkAoWIOIiNRIVw8+HkT025YUprZ7QA3BzrU9yQAipZcrvYP7upokE5/yn/GBq
cEDtZJo2VZREAuJLI7IGLD4b8VXFVngsX9c2q37zCoPtLsSyOxbRk8jGehR3CKe99UG/LBENeSea
8FsMAJJ0k17GDyPb9TvRS3yOwTqcdwURpWknSYRBuLn6UMeIKDr9kTlyO0ksJwD8Hlbwm4qJyCSq
vimB6D0um6oL7dgdfOrB7Er6j1IFMg6lKySpqI4Rr8h+qmmr3xreDGIOz5xdohOIpyQrXyABRf0y
8sTHtF5DtC6tlLpr2oSu1M4luHLjFtwXCfB+TRmIEjkLJMOPN14bHSMWw2YkQRLKnVEI+ona0L2T
71k6TXo9Cql2DYpylNdf3gBrPiVzoItVwjGk0ns95HQqGZfBI9xOeeVR8619kdBlA2jauO7jFnVB
btOThLOKXso2oMNxGJ6LDoi++yiTONTfgxU1rqM+zeVJXcHO9EWpVLUXoTXEkrv0CIGJTg1DHJlg
l5LlolYrFotaU/mDtUSi2+dyDRaZzBC1NUvy3B2kYfRfVPss8H0QTYepO65+BoGWpkMCYoRrvBOq
Hqx8O25aKYkN7MTsCXd4CDWzuMYTJKswNJNFgdmXmK2Q0r/3QebC9o1UShjM6ish/JTgX5hjpCC2
MZTdCHzWAMQonlDQw0b4VaLmS7wAA2FNqZsUhVty5/i8gjW1PdJi/LRxpioZ4CwbNIF7/fWqzm4w
2jzq6rQjos5DFCijTHSFK5HQXjkjLm/7OW6f2gEAW2uXZvvzfQ2emgltGLzoYQZI18TKki9Yh5Sb
rXPVbseYlalA/tbx49p8Zn03SlQyQHRPuUopA5AArKuuewI7u4/d5CERwXqOvIzeFRoaMPTr4kYJ
gvjQZ2opVBc5a+vbRyG1EU2mHQeLH9uy18CypYmy7zp7sqgwsNXTR9O9iCXSgyOrq/EQMscDllsH
A/zn6cKdrOHc4JQ3KsNiF8yI1yaloN6s5bap1IFNg/F0yAvfjzbmn1/uoos+eN9yWei2U0zplREx
/lTJjH6hgkeVjEmta1ciU+5ym748vQuEYYz3EZmY1Ga+QRkW2jdLSrnXVlm8Rs/0NjxuOHuZLrTf
er0jOklKRhjJwaFE5oz/E1XQpr8ySGkX9CHnSsecSpIEU3NEW9zmt1OdfFRkbGzAQIgBXN2Abnar
c/QlOgka+qpF3oJikGsBvIgTE8EtONU4gyl5chrvtTgWh4elexiTt6bR6VQZMr9iY646nq4MAaQB
3GCZcuKrRLcdnUID4+W3F8Nf/+ZIgxBDylmqW1gYPiyWL9dGG37lWE3/SEvioYomOdrIa1e439pr
aUfFK4MIbXWzFfN6QpRavrPJdXVT5JlPfeRqxZ1Cvqvqcn/ZvwtBvLoxQgkhGoYNCpWFonCPe38D
d/aQsuxm257HJ+WJKorrnIMzQpjO5Z5snD1KajGroK1908tCF5pU2ftCxu21bUq7qFCHW1Lx+BOj
/plkrAFhys1cGHZ4jjcfx6EmaqqjJH/dpZot5IHP4Hh001b3LP1T1FxqmbBRuwbwaQZm1/2kFAq+
OLwmoL/WjhjvfDrOkgrmLyaY4Q0VCEn7WGDiZrwZpwGPHIIwPagnbY0Iq0MyQlwyzf9SKJMvsbnE
4KLq+YEshdiaIuPNfJ2arwPE2hTv7bbYjOLSBCcPnClZd9r8E3XCtI5bPnJGOEf88ZQ6KSfKWVZi
o3W5qawW3ZUECp7rJ57AFCof9I0igzQr/fshcPsrdLOLTKeZlFuJeBkaF08t/udDbAY4+8aGaDOZ
BrjFzPPQg6LCRDaNC5hdeNtS8IuWZE5aWMsQu//ktzJBVg2GZCk7llhlV1kOIOWkZwMnEsQ9MryP
jfamS5BjcGaajzvNCixqFGOR0XyZjKUiMCTn5vGPmkDtnfTfUTxIscmTHuOU5PRlLn7A940wxoU8
lLh2RGCg79/PW8060AdGsXjtoqs1l/L26i2jhHuva5wuLJsTT29R6xUW/E4GFJlW73VIIqOYTrvy
AU4oRC6T/w1tRdr1PsRtX6RZ4gg+7Yfs6qasoyVvrXSlbBtFbYD9f3s298pMmd/594W4B+F9qay7
yD0QLrfSdHGa/8WVMqeGKbNYhiX0IreYQM7dJoZ7Rty3cDIHYD5QlX2MLGPBa0SyTbmZH5acplRW
96nJsf9N+L87rBENKq1sWpqROHdR7q1JaJ4ELkHKavUASYfPs20VlT5L5H9vrtAdq4gyqgwsT1Z4
1mSlNC2eG8Tj5IXYGwmC5BbImwIhLOxKkQNlPg1PBV2OdGZljCR0ZT3scfSPjfydITv/ACzisfU2
IVsbkfojYyo4t9pTgLxc6/IK6kR7+bHdZoVscrGca+B9JbW88RVxAxrYZa8PVqFyCpKYeIPzACIZ
6B6ZBAN6xN9/17opp/XNnR8ad/Cql4ZGC/aqVpjw9v3JNkuhmNopsOiDzjgAJw/snMiANXewv64+
YXSa4sgGf1cDHyFMcyukVE4A0pOTkmF9L3hD0jPec4nnqzo1Ywh/+MmbeWseN7rC+hAbk5nc14Dc
edFf00QVmHvPFISGSb+9WamtTcGuRi9b+fzUDqpo0orqdxvtdGN2B/tZsG7QjZP1Gb1EKePpqzU8
hwoaqaZAkclprhVjxy4paGljUxGsFYgjSbn+wqsUewpm+FZsQ9rf31ZzW87hmJGX9B5LFRTMofY4
e9VOi38HVkSQDTcFg/Na3ZyA+gFtdL2ydT1CSM9To9i28uerEbSSix/gAyBh6G5SSk/0Q8Y5Z/0U
6Pv6cRy+1Hq3myN8As5vhvDnCURyghAOA1sLxSeuBDCtCdpQ3kFQADZ/axBllW7enlVCLNr6cFLg
9dLP4nhWXyeWXU9Ab8TSFcGRdMlItyQ6dsWbzvxvgzm0cyx/JN1SBtVKDnD/1HkN3jhGsDM9BRoR
DQqJJ23gZ1HRy0/qpOqmT+rZ573J7o6lHjo4v3sJ1AVo4Vs3P0HNS4ZEyDbV6qKDT0/NnMaW7zho
IDvuXIZgLqrALwy8f94ZUQk1MxoeSrsCK9Q5I2f1MIAbW+iJkCZ2eQvcYnsJqDdkE5g47U4/fu5f
jc1OC0AtVHpOkdl8wGUNf5FLNKeowuqI8xSJl1L4PsUBNDutQzxhzQQh0zEMjQN0Irdd/o6W3XeQ
hYk6lEm2I0H5JKyvj5DOp5Ze0Kyg6ps2Q5wRs9PJYtVW/wVhWwCq3DkcCSmZCXTRbv5LiZCR0hm3
PMcNH1dNar59lpBG9fSyPoUPLTwxITW/6xLR52vJYQYj8Kznleua2TIUcuGbL1nDHPX54vjNnMyX
TiCzO9PnFpyxAOdCtTAxY2ZCTKzz7uHp5egVJolobNY6clF+qP4FTD69intZN6iFFdWZFDahseFn
qtmF6qhTaOEP3j5RP0sD0SKBPO4C513JlJWUolZrxIiZ43Qm4caWuQu2tIaZLkFWYfM5Z5G40xvF
FJ2jDIsCE5d68u8noe7H2pqxHd4/y2bQboFb5sEWXDGNlrmb47m8q++juDNoL7Ri24Az5LE2qE2Q
8zgym4/EBPKnnZy96NGmR3dyCRD8WzYIRGsb3/EYkDQKZvZY/mDFIT6k0T4ajWN84n76Rty4VOBO
s4cfciue+Z2k4N/05G1Aads45HTOU4OCqDGY2Neim9gFb+GUZn1KZgiIbJV2dam0xBuajnpJld9l
0pVxoAYIi4+qcMYxhX2/P2klC6okBBOtvZJwn9A/HF/h3m9B1t162/cqdfm2cOau6NlxjBGORa4V
aKaVXX0RkTdyzMREriM//9SHVfMuVn0y2sIt86uo5I1ZwYnLBP6sSirocBVmceu+xOrPLvJOZwtO
IpWpyyAx9hZ8MJ9YsXARzdUpayZWQ7Yta9GDJk+G5XQhiZ5/PSikurAwPLkTJdkXjY8w6YW+eKpJ
OGK3oUIvPR5kCpu3zcITgkdtxMUT8cp7tY0JJSpmCuhKgfQeAk8wrpPIbeTNu6kv8nC5eZKEBTuf
yMMnvA/cpRAgKMDXEuae+p+GhYSWMHPTQUVq/QtEG8d7y7aq7PgH95UowBJiac1im8ae5pMc6nqS
8MwsrPhQwqPXGSaT8OQUNIN4ROhBmnH/C7jvksjE7iFOhmK3sM2gL1wzKfDL425xs2qNkG4b5o2b
q0epaP2WXqKeXt2rOkAIAASoC9SBUb7b4tSRsKBnhm5B06qvjPLiW3WkmfR0AjrNnJbfWwuIssxK
bJjV7BgmSeJu02mUPrr60e8wXNN9hk1JescKk/g+AVb1cWKsphI45EOk/ZoV3iL+ZIN6F9zHNQiA
SVPOU7iYN4FUe5OPIHqS/3Qw8cIK1i9tZeioXlBkh+C+wgWPUcAJcWV34jbIzqsa3L9/JqXowCYN
mvQ4AUvltMoYYxCfwjBR3Uw9DMJjyQwltbSkrv73Mlt+vWf5DWE/KCOJL99zk8e8mX84UD8hhRbH
7lBVGoqqE28Snz9CbaxHUd1tdsrYMik9BMa1X+efzOZ3C4j5LE9lc/AYUfzmDnUdSbqoUIAa124+
w3wk5cdX99b09RCLjnHg5itrE4DEqewpUIFe4gJgT1t0E/2Qu31Z5h8F/BqMlxhHMBapV/hbugx9
xAU0MPr0QU+mkjiSaviheirEWDxP31r/ftQCjiwryjJBGW3V5XjO37NEkXLpoqCS92epdKDGKckA
MWP0sJnEPZEWZFRU3PWc+4+9RZAtI3tpLUuzBwxygSyIepfikRRjCtPqNaZwSmcDhukx7YDC2HgX
L44iZJUwmFtCMx87HsOdM5S4lsIFwcXP71jToiXuc2DL6K9jXI6B/DOkfbyRvrpGfnMBEWYT6Vkk
D8ja1AbhVcqNKxFnaIxSqfePYzuS7MRqLLipGgPJvPcmUBWJYtNiXg/xtJCLesMKxLxHj/9wPCVE
nrI/v0MHJAVSaL94wjhGhZ1KeRHeyAWyN3IzZLkyLFcLjYDsSNeLb/V7QFavlXSpQsMw6WsiACs4
D+4xF3zTJjgar5tFs6ddt+sumVpnigPOUf/8HUqcTkELuGMrHeVUUeyCsOoqj5Qh2ZT6DqEXpYRq
YB27Jrnl2q/LGFFxpATmqMfmVONAIaszKkp2KZdf/B6v+7l3nP6wJ0Vk0moB/5PJlr91WGOLcpDi
+azkMYA37MV7aCoEgFACDkkEjI4yHNmIxuqiCcAKcL9P5oElSJXnTW8e80COMb6IXU/5pAo1+tLj
DmvJzwvprvB0E+e7nxUiE4LZg+IzUMsbDMrBnjIkOwPjh6p4EyeyYItdF0JnDlpT+JYcmNTiolQh
YbuhlHi4I2R5/dBZdc60w36GHvhZOkNHA+BJaxjwl3eW2Ym60TCxk8JctE/o/cmP3navYEGKJ1Vh
1+UiVjq3NT7eGyewyiyYI1caQDhVZ41fudQDgpb2hStBHkBq2nMLLJuL8q7p8xzqRj7hCz3W6l+t
+8FOB6uibGpGM6LvZWbN3/VuQLb8Ie1/ugtAxBJXOqe7vJ3K3lLQGbydhCTi1h0HWbSqitrqsEGJ
Uamxn9jVeS6nUVDZ9VfMjH6U/RALlyLYEZVCHKlvsFvzuJxdmOxne/fjmnlyhBo6DSMy3L1VvPI9
RX7bFyXmlDlrWGiwmtTbfd1dOFSC5hozwjKvSzeygebm+Ld1Wo9b4+6Rk55YuXeKJnWhw1eLS8T7
MoN7hx+7L7YeS9WdAaL2f9xkH4hapk8fuiejNwJxxhXxOysTzymcfJKq57QPOyXhKPb6KqbrDM/I
1BOeHqpt+uopb2HZITPONr+GKn7PwmsFAddYB/OAXiKtW3aaOnljDeY5SuduRiJrhWnlaLbIFzXr
28YDNHDZcrkCr7UkHDWoIwHrSIv/FyPm+6RvvKxOvYQG1x68aDzYwfHaSPTUNrDhHsYWpc37zr5e
FjK82ISIy6nO+LFEHxSA/BXxljWx84SDqXhTsw2XAvWxoztLQq3d/+i6Bq/OgcqZocOD7P03weQS
Czr5rFJzVdDbqnuLVrxk/rw33TXHtUqBzSLVYJ28Ns2wEb0a4UQjEaLgzlJkpGo/nbws/TSromSC
OKGAZURBy3wPHYiH7gq04E/A6dPclXy+PI3vPe0ESExcQYQJlrSzHUQSrcGNkoavYxupQhNJpV6G
gN2sjCkapE0cTIsksTRRZ/CUC46hf412vna89dI/esajM0G7kJX/K1nBP0M6mYz/G0/regsRoqYl
SrTFGHm+tmeK6XVeL6cMGwzzY4x7XQcaHvy1OWKuathRy7xcAEBV2gcho4j4s5tI18RG8x9EvkOt
i8uiqgJSlklSOJ/rS2TabaFrNecH4OBdFayt6Am6vXZunrJifqEIndg4x/swVkBv6cWEe9qUc5FS
CaiDQLK0cP5hZOlhrVE+Ol0hrYrNH+J9jk+jPjNzuXFRefjEeFkw816iYBoqr5Kcf3uuGU4G/DeV
rsgB8rtWXgehhil/RANNzCQ7rU1JHcGqk+fhTG280lkutC5+0I5/ZEB4kP+v9i/MP5rsbHEPhUuq
soGcLak8xBYCUssopJ0kIFpDA+sDU4wHKA7HI33V1oOLInMXNlqzDUZrY+wkujwwJeG9eYSo3PK8
gDFTkxR97NuB5/4cw5QiwHQrJ2zzyyTq9kE0NxYTXA5HodJiVSongaBd/tLhaDiHsS56+6N/AHQ7
qEC+37VTTWN6+5/wVa9eojLdTwA/HvV+JZbMGRW1lPrZCgXQrD/bSQ8IU+OSzEocnqlcC+SKKGeq
cjCZDsPvMEgveYQw/LRW9buJJbiT3f0RlcmEYgvgo0mtrBcjt1H1xDnEbvih41BF6YiQAWDnJQQo
4ApD82GIBT6CGaCzR4ucSL8r3AgqVBwFxu8Pvs0HZcxdl0Wg30+OnWRPOXVg4stOvr5zDT/Og21/
VI2HFaq2l8B3O8FyEa9JFt1I7NlXBdut0oo1oKPEA443yeL8tqlPSkBan89H6OKwcQUJn8aANHDV
5V5ZrrGqxgucYsjh8TtUAb6ruJgqhjZIAf6bhWJoYIv+/8GX84MsP/BV2eIG1ar161XPBsPIyFSK
TKqwMr6jxnd21oBm2xtnryZtymv2IG4zTMQas4su1dbFUxtQVBoNCQEE8bWV2qK2Ca4+PWp1oad5
U1R0KqZxFQUb3UUi6g4NmwOnd5ZAQRdlyDm8Dw3iw2mtCZbfR0eMKYUd3/xMEEcNlXkHBEafGf5y
sSbEW4cqlbXgr4tJ5fcDiiuIF/kj/YbDnGvr42vhYuZlU+aSuO3Xz0qDEQ8VTJ2klkuVZqfC8L78
AESKFuJQHibaKKlDqc6Av35Rnkz7yPZRW1DAgyHBoC3jqbtMomewLBFACivRbQQiXn8KF8peA6AG
+oxw0fdk8GHHHoaYe0psQ52rHz6szTRTIdp5fNuLHvE0o7gnfwWMonI1I+SuTowJS/CxBv5ir+P+
Z66AN3uOjs+xUfvMfkYABHuloZjEgsc1QWC2pTZaDVA7W916Bvxzdr8z1zKH8DeR9K+cltRwfP7P
ujCJrTGg8otpE+rYfMlKETOczJ5NqD9fbkmlSI2L9zoiOSIEU7nbF+29UOFNFQTl4VyquMoMtryi
WepXQgI8J2KicA1i7v2TCfcenEeXZpUpNjLiemWQUcNG5essvt1PjHbJhGEtLPFO+ES83PSUhtcP
awPS2z7fwK6P0VwYT1ZzMxjGJturoDhZNt+PgFw1fJS//6Zb/YrgLURjmRnxxnswyVzuFq6fYysF
/AEjxnirU0OxXV+cVOQWliwf5NlF5dqk/Y6qgbVn7B6P8BzhboT5K1iN+ABe38YGZF1jawWE+sKx
lwT/DP0B0i26kQR6Es+FmMkI1tQDRFNRQD64AtCiJ6WPElNWws/qOneRMLZ9voiM63KQ0Zny9q4H
QG3MlHVEuxFQSrRAFWnRcLIY357gIOCpCY52AJEceOyVY8v9i0pbnYvJIYJeN+oYXkCq2LVVGcPV
Y4JNa/s3dA5+9yV+hZ8RTtt7dPJ6xbf2oESqDbvVLjP1oz5oX24KhLKNkv8tMdv4ZbMcMBC0dQ6t
KYsbiXQY8AIs9BOc9icS/yB0KtZxSPP05/O+dZJw6jIHiGiYGjYsSvYuiPh0vPu7tcMT6ElQXThZ
yxRD268kxGMH1XicWl01/FVye8WCbp0vyN1oqXS6bUXf2B+C5gzMu6RMtVBqnA2e7i/K1KohczLE
t7lRZYjjmVVsqTDbw7PgB4ukmHlsXATJokb++qmcNSh7pFlAwuyIB2hniJETnnegmNZbzo5ds6yp
wGR7DO8zJdPqofbWptgaSAdgM1HMrxuyR4GgoZiooQptmEgdh3jHok0Ts4vE9uTrzxRtfmsTYb1z
ua/9PFYZ12lEFIptdu7cBYug6XW61g66emKsu9+q9cvxunZWbyj+fllxFWW0ucDT7IUUh2vP7MzX
Xlwr9g/cR1VSa4RKAUIRrvfzxcA0DqvmvdMnD5gQWLfJDzty3MbC1y+zO8ijDIDSpACkQLfEK9Xt
8yhEUjxWTQsShfplwdBz7tx8WnFWtbdLV7Q7GTlG560uZ59V78lgMWXtvPaHfKx8DlBoBNf/W5uK
xwzrOADTATzQNvP8qe+zAta13kfVvwDe/QjFZfHbkfpdtz0xfu4MbGhx5O0YF3Rw/wh8TfSObCu1
Mr1CRBO9fJFnfgi1UbvIQOjO1WrtnraDQ/0VlVMyuT0ZCe7i3klhVr9gQq9xOosb4J5Ka46M5mzG
jfHSMtGT8PGepUysO49c+nsHK81DXxrUglYKFTgxhaoKtlyDmOKJMqb265DTaMVDFb8lghMfchyh
gL6wJY52G5jr2v7ZHV4vcAi/CbspGeu0eMojT/mhDACAJZmcI02B8UI84+dmrtv7t5lisDo2HZNZ
iRkCgUd8AafDtTZlOOnuSRrB09CWrWGmJdh9mVnkk33U48tPsmbKY2TtnFghhBd30WnMierV2tZX
aTZgUKdMwzcLP1PtrEHT83BAZW3tRoQYfDA6vTKy/ySUK2wZT9HzTKA4o7wM3HxmTF8tIoBvS6g0
77nsyNik2KVktEu9tuAtDa0UvKVtB6CqoPXM6wYSBTmBh+Njj0XXu87dNj6YAfO/o6gAcEG5AsHB
xccbbuRDMbkzVwxdau5WKCn6baJukCCGGEN41IfPng99RqTb9xB2cU0VZmYX/K8YWEyOXBmHkd0e
cZwBEc1qc4ugtnWaCLKlmGs65x8zOFvqyIqwp9Osyt186wIS7SWhZkNMwIAM4b+67uArYek7SxP6
1Qq13ZhgEOa1h0ZNBrJI910HLfXtQPlaL8HAoE8tIVypwfoCxwm4l3YsU8Lbe/lQ5+hx6gghUScM
2dEquhXk2A2I4NJ5lY6OGLDCa6RKEq3EC2imOMABqSqAHkStcnRuQrlgF+fQu1QpNGzjZ8NjTyh3
X/jkVGWikIeu9LveUxkS2g2Jd11aeuaBOHmlvX1bU09uCSX7+t+9ktNEAxgtxuW+QWVAjtiEtBzT
p02ncmaxfu1U/XWvs3E8eG71m9XR7uX6rswcCuPqkjw7+jdtCSXpeTXxe4+MPZ9+gJiXDBPK3gVS
Qq4MvEB53j0wF/o2NDHQ66VmZYsJAj3lN1c3j5pVP0oNh3IGlTg8kzhFVhHvy0GV9+TcrWV1GTYJ
Rrnn9Fm6B9ogOo+3QAorDAmcEUpiZZvVu+miuW9IBMtluhKPDHBYavO3wUsqVuslZW5oeG95DO1V
JlRYyYti/VwYuDYVU4I56CTmfJjOSqbPIK/2d/9f+4Fm9lQgVCwloaZ1Oi7zWTAk5fPkchi79QCP
jJmHl7htiezIC0MoCYuezQmnT/kxbEjJ552L2maKcehiXbrNeBczxOxTDo+Ae0YNDJ5LrLbci3u/
iftNFZ/6GY/uO+msO8/wqS9C3hwuPgppO7mkNA8Lz4S1oz8cBZ7xCOj2oP5sTVEziuNaA44IwB9S
lrpyAFX0C2wWBRbaRavhnOWkkCTduSkWX8exE0sipK9Z4pRacgD27G2PRQ5lWC5+0EJFxuaZNFes
tAWA5XqC5B37gQtFP+4AbAPnrdN8noYWAsolTqkFzaPghheWoWmO0lwOni6nslGY1mzVv56MyIVW
0KbmRlvY80MX7QlMmKZ2V39ISDEvYoOGODDHh1X4z3ClFglhKUAu14kr49v97Gj1GAP8aFIcLVMB
BwGC9bDcwDBGiUYiiw8c9lf/kXnB29qx+u+kktUK15NMG3cBce5rrdMpB1ULmEdSz8nxeWLPorEC
Eku/PaERsQL7GZrf8vhyUAK+GgWxLFyIBIt+eaXwDdVDwHcmhX4qJp16Ji/WgE+3GFlkqnKd5GP0
oepK8rnXa7IXG7Ov/vMwgjsbbi74RhKzZniZWWwOpnkj6qtIzNuEZINXPG7P9ccUb2Jut6ONMYx5
ZLufzZ9qZpB498F2RgNxWPxxgs7+wEALDxs3PdEHq+lRRR2lXcPS34tbjhfMZkbUwQdANxNZk9WA
Y/PgxzoEYzuO4KR8YgdxnIas29bLP0uOGBYws5H9aTq3iQ/akqBOKfe/e2Wz01PWf2hdQCuDFqhG
fyokTlwmImDZfhtSCZ3SD4I+gKF5mbH9hlOSWNV824SNCtNQVvQhdF0QgRo8IiNqSDvicQgf4EiY
VKR4KMZFX1w4y43kUvFmTzhDxTjSrFBzyBc4w2T90QJILOzLrNrR6umdk10ImxA1tryq3/2GGubH
vFmycGGrndLF4tM16QCyU6IV439kU6Xa1bDjce8z+szFzVHjri3llemhbjS5DM4hXnDW9FnwKK1K
RgSgIPHYa9FBIzk3lF/Of6zu0qyGg/O5QNXColjvYpPUf70P97U96VAkKhr9dIMvwT08D8uAMO+0
WCZA3F6vMuMJM3W9BvWWheKuOCr3hWfyxXYccbFf87MlN5wYkbbndrjrkXxQs8/gvUZxxtiB5NHB
W+InJEPnOqjoVOW3yGzQoVyX6L+cOe0F1idLGg7BkbuhjYtDS10nxEglSCSunSp234OeEe2XL/uv
/2gAnWX38GUegmXwvhQDab9qIcGTG0vLTFCmG7hzCY4vssW7fWyeizRO458FPdiE77vYIgVgNw4Q
MzVCV+REXppQQ+2OU4mslQj47oFicFvkdGE3MIkh/D1M4zL3LlDB8YAKMDRy4xsJ/h8P3T7dxILL
+za/F3CoWFPbJa71U26lOpglBn3ieT65mxVUv2q9JobMFSaMiuR+AyzG46i8yAFGk0HabCyjH6VI
0iAEflxbg81CD4Zf88L2JqqjRGVOry1VwuAjq7IRngS9l5xIG9tCpUvud/OUHLesR3p/G3PjUBUF
9ga3t8wOkcQWgE0OzV4SIFfKbJVFXfMXPbNfsitEfV6l9y9PWr1719UAfQBi5CF5vulAmZjHkecx
EYK/xfMkKZPxuiDHTABfI8cjWvVmVATtJzFKNZgM77/LVq0q1K2XYjI4xaqAcvzRUX2STLOkCB4N
ySZYdFgpaHTmAqtLCRtXnpoTe56NyxFJvsyMvyIHgz3yrSTr1hrlc2gxGkdAELN6w1Mo+uzljyoV
sem29pvI3pDXMcCAKtRbGaWGwzJWYfXb5n4A1g3B3nUIMDvuEQtTdgGL6WCnj5OLFlBGDAmwtT0W
NqUQt9lbxroN8wPKp6DORcyDFKo4dJ4x+ZG+Exf1m+2WCyajKCHqSgqo75hw0RK0RfXx4yAPTN1A
IFJVa6j1pHg1vcxcBfspr85Ap6qBaj5bQ9AxltZjallRzMuG3GF3Ncc4j+6XPjM87h5aDhcVBmN+
V9oRkvguSMvUv8UkmzJChdI/HQ4I8WF+ZESFFObCmkNIGTGnCCcavLnEal8wlUteRYNEdxwBP9v/
TDOkOV/adlUyD2ylYWwamNJms6zP2Yh92ZGbFcAfah8miEURFRoUQw/B0Yzw9A9ehLPsvUB11IOS
WSd04W5UZTAnL5xZWixeSzELuOP2bvyTPr1FKaHkGkjcrAI8JencP8LoP/YRzsUNVpkW94Oe3GkW
8p02J8+YfY/D2+yhEbaoqlQdiZVae/qYjIvVtpiXdWPAQ/Kb+79cF4v6mRDXC5xeU7yHwRc+Y7Pi
fUHOvZFiBVWC4z4gABMz5VjADMkDs7nXgBLu9sw1D6p87OGGlKsH92Y3KiPWWwBDK0gf8OTrXZkG
T9pue+wBOyrDDJp20fYQ6koO94jsA7dpNEYnwqs49MNc3/lLBQ64a0+Amrq4Qn+xf7SmqjVHIZ8M
9y51otQl87865MaAPIaE0tYpNYXx3apOdDaIPN3Bg9ty8a1j+a2xSY2nAiakgoNKlESZ+6gcNdst
v0zaJZpFl2KpenNqgqS/nEI63KTCl9k9vHErXNiDQRBh+YH7+0M6VSHEnP5LeMbNSCuKPXNwLwCO
zjevonBZqm6qNu7exNLO3wokzsceYnKEt9ikenLT+HfSS9XgN6EUU72mI5OttDfqnWLYU1GTbFMr
aaYG5zHyuhjIJN7K3O4S7cr0bC81uTlZ4876CUQVmw9e+pKrClkDwvF7J241V5tBn1OP2nmxvNmB
fJyhOufrf9FDwtMvzL9J2CNzwqTEVn1cNmRsZactSC5nm+9Kwh9bvnorjh5JSS83sysODLMJ4jTh
NU+ZhkNfycoqQK5ChAIIZ3UW1srlHPEXXfrZmSw3MFQ8iD+3yG0SMR+gKugb43d68irtTN7rDhPA
zfiCilZdrwKORoyYxoU+G3Lep8jlox9YFfXnEwgQhRyy46+L0bXD/DrAq1kk3EB0/j3rAXxtRAi+
DIam/GRbYVALrh6GtRXAuYYcL5HiENlojexyre/BtsOjg56e9HNYKywhU3+3Is1F8OyCudlN2Puy
xAttRjieaJVeLmx6L/WkD+mbkg4Pmp1ZIzwsZdE5l+4d1oBOAxf2LLgoH1b/quQMTJ55HXNr6TG+
bLT33UunjVmjx2bglDLHAxnQYuO18pK2QmEZFhBJ4GNmt0W/dIdRmyxkrQ4jqRIwX9hLmNnQQjo0
zZF3hO1P5SFOBIAny1hHc4saB6wzjyqtp6XHOEjmmhSNRcjUd4ETjsUXjDas49gbj2+S/sOx07L5
IgjOgF250Q03BouP2S9EqIwIaX7F+a/Urce6HzYebxSldtUpFEhmOh5bJKt9+1Xe+ZhKQGHk8d2n
odsFZstRAf5ZWtAGj43JuDHAtTZF7U7PYYjLlzq9nDF2kPj6enx/YwBBytlxWta3G47g3rulal+s
OjYKGa7spcTePogO0c9d0w4dJQifwdMyDexYmI68oA4xP2lTB1cJSCufKvKpChOLVlae63bRQjep
wZQkcghfeAr5sCxu+XrfnA0V6Yjq2TEVCaMy+XbgP209Bd2GTsPZkVSfx5OOnU7CCn74ovuOtIzj
y1iCVc0avR8lNUEX0moVoJHT4g5COjmSllQjUCJDBhajHUGe2WwUHN2M42WkaYeGnoiJVZORebF3
pEnJ7wbuHDvDazMvjVtCB+kklcr+ysO8N/XgHkvWV/PYF7F3hOT4tsmn5PVL2sgFFsNwZ3LYF7bn
wFgNqQnDwURbnDNYkoLSgy/A+ll+JDEzCV6VmTiOuid+l+TmSE55KTEajXMAZMt5zeJpNEYi+ZgV
gsJgbJZKpCUzxJiKmeerR4cQTToNfbdRqXLGMaM04KTEVltvHbwpIgyH0o+JdSR4anAhm5tSYME7
0NiOe4myRijEAc2k4AI6tl5gM3YCWboLhbYqCma8bWJJpS3O89oQwlq+QLGGPzRdV87znYkD9906
4T9Eyps4UQRhUwyddpINJmyQ0UdH7a69IdlCkSqZ7jXpZETPJDSuT28KGCd6Aad0+eabgoFQs9ba
GFKyfAGds/tFX8nUP475StZgjj20HEQMjUo/y0ifDmg6mZqWGSie3tZuGBaPLm+RR9QH8wTTO80C
RUwBcCflqN7WD6f3P8fU85qsqSBax6sP5WXsECmKSEPDoBY9WsD2R/Dfo7Xjg+y6G4lT1Riz0TaZ
gG8dJVVsBdvjmhMRezmX7ItGOgseghdFamkqpSFMNjDU8JsyOwNtUT3JER/cfqMLeKboPE75dJlW
IfAS7wGDY/TNEZi1md6GUadnUp1P/GFzTvcLR8RYrLevLLa2Ee5eoX2wdOZfWIuI3o4VVuWcWcQG
n+u7u4mjV74aY6PgakqLXcGaqOfcUHhFiFyGQ31rsEHwgoUqyXX4KHpfBjTRK7hR3pK966qXPJa7
wm6uNc1mUm08YZFDvb5nrgoRxM9LmG2+rXwp25g4gSntjQ1wamy++NuFJfrxeAB1GSp6oIKj/YY1
G3+gsTJazXiAd+aq0gmADUTYvRThsNAnxRE2dDtO3jvV/kV8sNBSyQCDCPfmNWaMNodkhVrrO4Xz
uOdoZRHqrtH4vTRwMRbti7b+WD+sdePtIN6hgPC1++a1ALxpAf6IFJ3NP4naoZ3CXMMdO4JUexx4
2ySmqA0dHtQopkYkxdlop2QhypT/4XfjBJ71zRbaXZRklHY0HZQWDhFGEzpi3ZGsP0NoeeitAxuQ
SMvcgxQEK2aKC5zUL8GpPbif4opW9GciKyV7zrfIwExjJI2uoZkyQPAQfOLvqtTq+uyH+prItQ2R
7HIEBoAQXQJwvmDWo7EgiaugY2oOZXu170jzI5E42UP2A1zyr4BwJyPxGGUtd2ODPoRwByN7TzX3
xpvhjHMiuA2Tja/HwHUmyssi6jYvcKaF0bsA/iX1qrL2n1P0nfBeokefn3l7/ocCAcqFBMj9fCDs
kF1HRK7tPZR3uPkSu8clgfb/EZfuOp5CTxuoqYyij7/RSS47Fjsnk5WfqaDYZW+u+Ecd3/l6ICbc
Y+H51W+Q2ojP5AqqvQsqvhXuKkHGEBGwogUjfj8zG73VrZHGKPY+t8U9ul7DYc71dJ7YpMHfOOi7
YsDoGfOeZ0Z0o6XAk5Ct0NBjV1Rbca2eIu0WHMKQM8vamIHiJ0OisBETvt/TiSLZQz8mmr/RE8IV
lOl6YDBP7q/6e9buFknNTYAdNFxKUWlle7hN/tCQBiYUjNHBLAb2D5YQB+MhU9tIaS61FNNC/YxR
0buNhCHCZ3MxKgo+NYunRmy6ekociz/7fuJ6GwhbhYBfo3p4uTwWGRLkApRhXMMckzS8RQaxSmtb
kVV/zGB4zFBH9Qd8Dsu/Ndpmkr+h4Ge6geSY+gS/GxO/7ds9kQkUGY2XnGUeg3/LcBrUuKZuXWK1
t5WJVvbniD0UfVKp1uj0Mw9QEPW7OJ6toq7ZReTDAQ9gl33yk3cI9dS4gN5pXx5UnWhsPpC0riHF
vBHDyVk0kWUODPjtkOlLUFu8IQvyJ7pTGnocMP2d1zCHxZ9niuKCgxbVLKzI/ELigpQyKWdYFwyU
tO0jXGViOzWk/ziwYHZ2YXncZjeTTDEPclT/RfXOWJ8/i1u0WYTzeo8uxxPqLSTC0XaNtbd+tS1z
GOKgc0LsvcP66XcUArBPyczTNh9FOi0wka7CuSuvIkKRqDRs4z+YI6Qf9Z+9igINqKtrJ51uInPM
2+dldC59FuRNW0+9Waqw/Ivg7Sx2fuaY979Dlw8vTQk6Xv9Erg0YZ1VAq0lgUoZwFmrNq9tQ2kOI
PK4Q3FkwuiiuJGImwqMhgNlzpo9iZLlos3+ESvf6SNcJvVYC6uOP8Wif6GxrjWVA1JcWIo0J/INv
+NtLamTkY9gmFlOED9iOCEn2v2weiMxGl7PYlOSYisXQleyCQKcxnUm8qJHrhfhFGDbl7tQmTwqA
ZzQ5HoN8nEHl5ndGvwcu76uAtOmC/Z4+g+ewlnwY4bfMhuHAFqe9RT8KtKx4S2TGQfQIoHt0mDAA
sGxFekMUPs/hxM50JyluaZD9GMwJy1iUBSMHl/bVR/d3JZcTMaX6fxNoSzkW5wqRziD02Pvx84B+
fHIrh03MNTlIs+hvpyRz21wYDcZYgNUEzOcTTRFd+0j2heY9B+vzz1jJgFzrxVgtuX3VbLw7zZfJ
JuniwX6rdTsqiIcjer92tcmeCZ3mCK3W6U24l2Z0eiG88H0EKKAkgW1rO+f+EUgYNPsWYZ5TBq1/
3iNa5pFF3ywhYavc811iTXsvvzm3eoddD8atmDupwtobfGASIzlyKidMaZjAhd9AkPW4GTDalgI5
zNVUiHU0SOpIpmP477fYW+UR/q9JRxLXQblgx302KFAwFLAoKM6ObQ8jz7dqzoK9uNZtL0kQuPB+
x9HrkIZsb8MrtWvMffNgPjILCt7OmM4lt54s1Iu92VMEJDA3Ina+KN9Vju1HF9LCijyoLtwjOxj8
ZX/+MlN1Am0zPuqu7zYIpYZnsKiAdii4PJqbsszJM7qSn0Gp6bs+r71AIKEENUDEBI/UVXVXKOqy
Yge6GsImZZRP5gcQk+pxHCqNlHp/wTc+uC0ccXOCKGo/7fxq4wfQ221652SrKz9ya3X0Kz+F0JPD
6jG8uwCXe1lwd7vKm6KDwClcBNTHWoET97W3gNk4e+c+rgjcwKzSsaDYL1Jm0PSqmK0ici6FOHzL
z0kOkrXNyLT4+lddIHbcLnlA+GvmXcJWjQ0HYiJ0eBPyENKCJ9seZITWsIgWkSRfXmvyVCMWxDvx
xzVh7b0TfVkQrL1mToEfdYn06qNWdwkb72RA1jMFYPCu91Bl7sl20XU4tOKMxv5p5IUSws2BDuqI
9eoqoyq8Yj0RWEEGEs5zH8s6ro5j71rCg5DiBnz6Fymm7UNzNVxcX+aG0jyAjTi2QvzX9njS+yXK
L17R3RlBmgulDw6W6u+N/voSsqVMgeJDAc3wECrlkrvNpb3L/FzMHoe6cIN2wS7lB8VYDd9yAirz
EVG56I/k/ZWG8zeV/Z9JtL6FLIXLkVa60AvhbKHvTB7C0CbyEQ22UaBiIGDbIxELKyRpwx5q2bzn
Xp+y0xJJaJ0VBS3feZQkEKzsPafSjFNIqvGmeRCUn8cGeW3lOY1kMZQNqYzR3CRbM7Z+vIDZqcOS
z3PQCCfhSXr2rScxaWTzx8YS5/Mxbdt4EKVYnH59dJEYfbFQrv3IoZqcka0oLEr49tf3PsUTFAV/
kKjNKMUsEsf1k8lJmBZ6+9Vm1GjOitKLMeBxBTG6owI/2c/oSPzEocrXYVh/TeBtydlEieDLCu0J
ki0GpEqCXL89K6ZmCES0e/J0Y1HVt0XRxjDLmk9P86N69uL/9wqsLDep7jDa5IrFaV/wwHy1s4uL
ZkaLbe51SmSgLZAAQfwmqtWzOpVHzGbyrzN0KxGTLSsOQSp/kBoUDKoVK+EJm8owgtoY+oQHPWyx
TPkYR5mOyYX7/5ACsdbYlMCE215kUJ/4qfJ/XQulQcEHE9yvS/3FQq5shHNbce2MFRPt3frnrc2H
phv4MYfD/CiEYGeU55gRcnsEPpa64i4emHuoGLYSUlfMzhX5/ssVlrO/gM9UOq00mWhqcO78ljSv
jaCU0AiKEY3igrhX3M4v5l3J8BSJUy7jSuP/cV7TblSRh3fokB8TXmTbTFrumMovL3GOo8x9Icwa
qg/RKmvjQTjMFzZmYKJjgSXmtA2pMP/49IrDLtrI67gN498W/PyJCJ9suARdomlEsXxoMFqe57n5
4wk4MAILz6P7PpQQJ5v23NEwcq5QSW7/eprCHno8ixsiLXUiG/iK8awBXwWHoOmK+vhVDOqYc73H
rfMCNdSg1pyIQZ3bD8IWASgKo/pKP3iarpUB4ELUuGlcvulkaHHRzbnIxZs8pIsuXWtgXJtTOgFl
w2YsW4v5ZtUKKHD13vPaAPrr6E9+V2cAMFmFNR3+GQ1YDdXNmJ1HXM0CG7nzqagXxb9uFJB+uB8i
kt6Ml+B2J+bRtyeQDqYk9owTxN9UYb9Xq1R7tKlp83ck7FPsjCkkyZ7hcys50rHJGSSp0OQAn27Y
6M/5ojqIH6oLntpL/pYitCy+uZgmpl8fhGXt5BrnIQ30g1fnkCUvezDCfiIYA0xSaf8onRwp2ZdW
2S9Cnhbic9dk05YokD8LptY7mx8XBQwgkURK0HbrNzBYnVdDlaOxC4OdVngWwZhtZ+aPY/LLZB5O
oXirM3+tehB2W6G4GfN4SmWEP21E4ut9BFQGZbRNsp7GeXKOek4HgdBgBH0aGPhk2OU/6WhjqL3m
oYkHasrZMXK0YJs0bUaWR7oz5pfszGFOGuvs/kvEre/zm6bmuxvEUJA+Y/UEVOVJ+Ql5lbKCCz0K
257leLFnl6n3OsSM/K84bFIFRPwyj9lNTu9fBh7smNYMPAooQzUo+jj9mO5NiSrPlOuNkM+m4njk
GFGGCRDKSeq+tc4L7ZNtUDPaV7B5JVPb2crOQXriJJT+w3LotR1/Dnc6jSl15B5jLZ6XLb3ZHIjx
joPNgu6wS26iO9LmAI8Ar4vWiY0HMT/34vgWTHD+ZIrfheZJ5R0lbTPid5fGO4LwfQV5l2xkKiRf
e0kKPrqGDnggpuebUzQSvhvkapm8MRO3seLwKLySuOhh+gELKyfwGO/N2jps9CI+7WnoByX2svax
Te7grf6RjShHzOlT6KKsK1g9nxsiVDFY7luv2baAl+CDm1XkyDR2YYc6jml8sImXqroLbCpsfKKn
PWfENFfRZ8MmEBWMyWhr0zFSNx7h9AZ2nQVek/tULpjbaj3McdgsEjLFRaNHiBT5LIm/4A/5fvuP
G/TAP6Qf4xYfivAwBBjPByXYI9m+fmdWyqllFWe5dAwmK3hSatqwNO3yvVB7uJ17bDkZ77yemdyI
+LuVC9YZK6zWPeW7bXDh7ki2h8eYvl+UJMax8vtu9lUCF+0MjwtHSDmMwfLmS/uaMauJoF7LVjZ7
TVQDdxYqc0VKZ4HuDL+uA29yolf+A0iMNIMEuoSv9A/5pNzk9wf+9gU0b7ydiGA9xbI6JWAJziL7
PZLwf51/khsfAK7Q9wXZGh/AQMp85g6gQhJ8Iq3idZuJN+HlSb74PKVkvl7jzZGNJ6ho9XepB0j2
yhOObe7EyO0wKkJ3qISPo/OGRbHEm0enYyAPa58kyEwPlZN5J6v7majtJcMZDV4uIBc69jxIWCIz
8wuRduYVPDDzvMP8nyGO2E2c6YeQ2+nthb2lbDVjc8LVA2juZCBbXj2UEerpHIsMJqO7aU3nXZjY
o1Vx+esF12L5jTWs7ESAHmQd1XPWSjpxcSCsIiFY1aXT/HAbyqbiWsWrh9Sw5Vmvk0LDrf0OWf0W
lDw1vkQFabxQ5AYD/SIyFixP0AhQgIsVkP2tXGmiTfYwY07g6K84dNzdXztWCxMBwLCfg4GCa14A
RFbb4X3kUENLFlQ/HMdFWdcWl/5Ue9saiTlshKmq5fg1jtpCE692Kba1/6b19EFBacUv5t62cTxa
URKb1OcirDM/FmHZKtRW/Lf7jLWXIa7xL+16xHHvpPPCcGxKeuMTPPaOt7knhFCEUvHuZWcEjLGN
4h/AEn9bnsxd+2Iv0l6325uoTXXC/qhll+0IxlDpQhFq627XyLZX9yvLW2e+aKknaGUryXDgeldH
UulW7rWI83l0WfCadW9CJglNJUTUyV8kb0K1HodaGR2mfv3RM8NeUGfjFNbiUFCQ4czpQkAou55o
Sal2jh/AcUbVm7/tg5a+B1a459YSKxqFPJpalOfBnOZnraqMnx2roPCkx6++rxF44oPKW608vr8O
T3L4z89VQ7j8Dd9j9NCjR1Z1QTfxS8DNrb1EL1n3LjBCybMsZpeahsMvjbJeXcgeqnbRHO2Rinzd
NXvU7Ei7/VMRTcNTnnuf8qbGBbcKZuJzzDoMIUjDTON6dOKeXaW/RsCId4utA0ZdQjSMUADxNRBZ
Tis5xRNU5XMo99HGOCejzMA/5eyp8+4yZnso6KSm+Tacm4TJJNYHKqIeFPw1qW/8C8Oa8OL3qZUS
TWRfFJ9L6vIEJmi4Z9uKeA7mssxhQN1L4HdGK6sTBf/zakWOHO/5+pbMPIzOaWQX6BVcDGrfYxYX
Wm3AIQ5AeJPAOjpSX+bAW7Yic37sbA4A7sjX1ip51RTc+VEgemdW2ml5ijLuCm0ztIFGolPrlmhq
e5ALaRDg739sGh+PTbPd93gLBteym8Ly6REUEoyLbNV46E7j88mygdg4gARVCLCMXEzKSejj1TOR
M7Tyc2EgNHrEp9ocA1ZczPALNpyTIy7meTd4NcdFJFlC0xs1vMi3KkjTGGgrM+IPaQaHEBcTeTq5
clL03fPHvw9f+UWeaX4GR/+Npum1d+TmsWj+YzvT96a/3sQl7obP5KmBpZpoLX0ogDuaeTqS8A6O
HkGeTUX2iM8g2t3ABjj0KX1Ge+5cffnODygPloMff01l/i25cgwNo3dODTdjJ11woYhSnOtsBwUc
xJ2rwZV625iadjVpeSQRMOrU/mg9CjSNglQBWWlnIPZc+M/pa44tnwKmmyPdqw2eoqzqQnd1lw13
ecO93yr3pnO7QcR2gejmUyro9s4LGU83zyOsClwozBM20dLftkcGwpkfdCVJu4gHjmkQFPNMVsJp
K2egkalqrs/Fctn3lUzhejG8D0v4fn+woiR+Iyz56Xcktc1AV3u8pRPP86LpplANNNK2cue3bL1j
oClE4Jgho9GfM3gCjeKvNdZlfOx5iobG8zrl0QxT1c5Jru9mq+T2Pcl15D3QD4zPq9mkflOpbuhb
AOjN1jMLif6tlpqwz+LORYNb54zbKD8Lkxw0savTh5Zxw50eFNKZeOoRMhWMIlQPSOjjjytS8ayF
iBN0zL6CNpwwmQDweHkJJsj5fCGZ/+XZvM8iRF91kx59/gpjjcCFt9BeAoSjfwUBVxEprMNHBOAm
Iiu7zsVClzcTJHejfG1EkR/fUVHeLMd/zEfPRG/6Y8hURKxM2omHa84abf/G/2IS+GxBvv9lFMR3
zMgd4QYgvzabjZhbD/J+49c4slNnNKmH0g+S7xwqXtVOETnv3AGSBtJZsR7mQlEe9zzpg+9Qib8N
WtfFXpVB2wuw4JY8JQXhn9GlNDaRyqucLwpIAgyZyCwiu8811Xyj9F0Ipz9UNnuNmktWNQPuafxv
wO8SQsuFW9JTCX4MtabUb5bhUjfenxS68fR2bn9BWC7BoId6T0LKqNODsX4ARGAVCUpVYXT/ks8o
+I1XN/k7k08FI+iekgrgykFKZvW3AB6lt1i6smV4I8crVkmdT3dV/HSS+o0XBI94OM+2X0HZU5l2
n//ZcQqhzym6dCA3ID2PFM5IGZzubLNmOSCP3xGIklxmFbJ/RR4sGCPQkZp9fGO27ZQXPdRpwoDg
oJTfpf2kxaYT+tgyrclyKsz7Wtg0CTMdjI+gpzB5wYa7gKhoVppZUAR3RCmQc+UYd/c4Kxou9sE5
9VSHpxAzE67BbqQ4+oawrMnu+MZVvqqyBQAZ9UaJlx1Bg8XIuFz9a3lih4l5cJNTkr5GpX0rfdmB
1uKvcET1X00Eqs3yn96hk3eK2JUfT1IVK34joZv8Z0ZwGHOEwMDGJAXmxzltcCj7+qyYtfDXJOZY
DWv848S0PS/Z/NL9+J3iUiv3/uyBEnQiQRXpWQoksusgajOiwi8It4cV4ScsU6gG/bqWdSVkDKn0
fLynAKCs/cM9PhguKqQN1EnbbnEaOosIOXI6ZmhS3rnoszUpOhlVrMiLGdtB0a2Wc5dULOTUqXhK
BLa59i7/K6DdksPdcpI9NB1dUV9b0WHbDk8+X0BU0/pt86hI2JzqbPm0E7W7Sdj5Ox5tNscf7vHp
e17Jn9GOiYttRT82RIt0wGsXDC6zmKFqoW8xRDrtBBby5nxMWU4haB0k2+Pef/CI93Tab8wDyh9v
Pmx6YKjYtHWMhNpX/044UBVinCFtxHeT0gX5yZhQpSN3toAvcyHbM83lhXN9i+iTn3t27qhWPBiQ
KmyvUdpXIMLx83eeCjiBOq6kavGmNcgDbzaib9LNOxLoTlijb9hNoGlsBWVontfOeglQcAPemm0s
5ahcWWGIV+/OhzBaH97UCyMBgk2HWQyOqQVaqR92ef6QFvxrLOkxyX/+eYFkdQLXr9PSwFCORau4
sGg70Pt05Xv+UOmRl5xOZzuknWA4fVCvER6c+NR0WpHp1X3/rpQ01WbMxlqCtZ0t5A17uXDuwuvX
7PQikEnF0aQuIP6IdodLhJZmdgxWAQOn/ah7bpf2k/b3KSQTC93rbhrlKvC+8UpQl0XO33zlCY7i
/E0G0S+dUwW4XcIS4Fk5/4Bo3FYzrr2LlNjiuX3UlxteE6YGfMDH9A1bzUUQCTsBEXvm/aMgCRmX
Ng5U2jBZtcwBKEU2eLbLnMrBtJoPE3lgArcyWEsevLntdw+wRCzaNBiiOjuVPfJFWlLWB6wmzL7h
M655b4jzuqmxXTl+DTvtoxXea5ncQ/s1XbTOxs2+4xbCF+VM/eBULcKhpPomTq12cSp8eR+J3pzo
D3sfSWrIPmBkiqHLxf0rmmwnK4QBz8I9GV7k3st6TYxxmAwEF2xs159teeiiKJCrTAu1U3/qyJXp
P8SmqSfEv20RCAKcdlrLDJwV6qtmQsu/Y5iZ1bCAmMaI0D3LKOtTI177Nq4LYKasXbpA0QFPDJC/
0gCOSyLUG3RrnDaJ7oAbcHdnKZ6gmM1ox2REC0Y6AklJENyWAn+Ta3EOED5xV4NPyvnstFKaFPDG
aIhIKmhnfB7oNPjdimvt3CA1nt14Yo0kVbomXMcDjm+PZDoC5OKczg2jK5toQqkvlnT+BxBB4I3x
O9B5p+GmK9LsAN7q443+t2kr3Aeeeb5sOGJm7JZrvHP10hm/wcJCDkzZZknDGI0/9LLGTXoWEUiG
uRfunkmCY/TvnkTqqQif1UgAfs9NTXf3KvJmOYyUarQO0iZjFSVpeNQgDTtF89oCMfDRmNIdlVZu
Z7diYCeAnVTmoLWKj50UB+gZCLkrWrSYPn1WfpyE0WZfbera4AzHL/qJlFkWALFgEf2kdGdThsfT
ylZcsvhlJhnVJSFAWbL39HnW3bjU1ukIoS03kRi9+vcQREBpG31i46z7EBwh/vGus9wweTAXqEJ5
0EaH+OzP6i1n9Ii1DTPOOKBfrBEj+p0oeVw6WxsB4sHybrJyh1QDMdjr9oG7CsQJh86BjHHFdVYf
gA50rjObWIxktbataSyl6v2dNsL9DvbEC4QE6JFNks218dv1TDWprznxb4eva6Sh7OU1vvwHDOMT
mJVDOpHqXrmfVKR6BREL44fgA+3/4d54pg+Sk0RNDYt8pY9ISUmJS6T1vW8WBsLaO1ZXUcblcJBy
XLBxcCRGZl0rVpjlnalqa33Fvqr+n/JBgjai8SsJsInhksUrvRhT2+nPFrSIVP/9vaZE3Xm0aMrH
mEu9YBsD+2SnHazXjGbOn2yXorb50rQg1tGMziR15w2cxZ7jFC+Nfs7Co8Tb1Ni1rV5JbpQ76DTC
GNPmCFbiRBFds+KqbT07ydrugbPD60wKMyolhLOBxKDsTxYls3Msc9fPciFJ+cpXHzdtrTyXdH2d
PigWKW2lublnYMSfmHhlu1vNyT9zkt9ESbzCyvOWwij2GXaSQH6e6h3OQXNgH9CQDr9OAv6V1mC9
/MoZKftvuqECCP/2ez7n/xd665xWgEMhitRe/BiOPxnza3of+JCRZlsBmHdxXksWSlYWf510Is+9
8Cb8m5RyehZBZw82odhahe28Q9YyCi8zolXqua7df5KWz814as6vXQsV9D7MKelIaNg4DrDSzhta
Ou8vRT5u78EKe8ngkqoyQg5EIr9ZEGR4Oa93ClvrcDFUrViFx1CO1xVUs8QJbpxBaLbG8/2MlxMg
wWTLc8OIJYEiSLan6OmNwJyb/pgL0RGyTac4ZBeJUIoJCNkcCj4WpVOxCH6OAuR1iP/pGtsJzYf1
uzh/6IYvnfZbZCl3NnKYAsl058eewPvAhPhtxghd3hSk60dVSrOOjflfZWtu9DCmiWLJgcyhexZR
NKJgMqT1kHWnlrTrwisnx/lvSWGG7xWFt4qr4Io2SgSTzFNlpcVWyOcVwtUVj4DRjQDf8hyfH58A
Og2xnM7rRE5LGyfWVwDip7izAMWhbi76YKUurXXLq/RT6+4FW9EA6ZbSYEcTDaj9+92Yj4PfII2E
HCuA+BBEDDqeVJid74rGCQRP65pn2N6jET2Ny3lz4AwrpZnCHaE1BAYMEWvDXQQMpJFTohTKGATv
CjPRoyH1nMGlTlKS8VHc3U3M9yxbg/T+LONtXOv7skYWzNwGr3tcThvwaZwu0GwBzscXh7Iu+79A
GuBUjgl5d98EzUvOQD+4frATCrkRcBbuiTYyGOWC0XMc7iR9w+lviuXtRBk6y67SU2K0IDoFilb8
rL3c8IndpHOFvtFf702vbZAFgC+ONSatlel2k53RDkXUt7Od0/M4SlpLFmWXfEvc++p1YBiiQGQG
wWvBiLrzxz0KDt4apYWUGJ0Pf+khvP0NiFBE7C5ZvMbbTcEhNp01kBmorwKG8oqwupOKA8aND4qN
SqC2ncQWu2whysWFCV9Iv/aHNhzZ2mWpZb1yv4PZom6T8mXlsM16NYsEUVnNQi6f/mWJPzh4MYuy
7iskFgCHBMaEd8T+mLtyZd5dBA9A/DZRa8xaJGvN8cuNUc+I8XHCRcKEg5kgnX4iPN9hu0orQdYO
gVJs8JDkYLlRBUieQ3m/65tKvr52KVBmiPZGSkxQ1mqfaUtLs8dn8r3zDAgbGcGWjAWuLAN1nZa6
nLqy7CBY2XllphiTkMSOXZBdGfhPEM+oRKe8RGeC1iBI2+VGVToZBRCFsfDoWqE4g8tbD247b83U
KCFxeHr9admia0pWnA/eBnroC0EyArqaVWaS+XElx4xL3GdulmW6zRcPVdLlGMr9gpNK3TRub76c
VHoMgzN71NO/2JXL1WNrMXmkjaXJPftfvz7BuJL0HbRYfqptOzI6TWzPKl69T2iOCUyuKupXKaTQ
ESM7VDduxCIE125PfCIHmqABgWjjYcz9NSYQygsWBvCUimQ38d2q0/si4tfcFIIKZAjQP7S89Ku3
4G4w5EOYvOa6x87VwE0xuN1dpPiWu3r8k7x1wY0vxStGWvG9skJDwAcXpVDxivlloZKbcVY3isae
g2FZUikxAbBGP9EfTGozreFOTWc4uukKv3znLJJXUltmMcxmj2Lku9NXpC2LxbhmA7pu8rF/P1PY
5ZHSAyq6UlRT90bmxpXe1Qaqq74mSksOfnshcAJPeWXx1UptnoqRucdzxtwKbRZxPacAGIAipuwD
+dOcM3p33nVbn0zCtASPesxP5PIOqR+G7q6Xb+7yuN4v5RcTbc03nYcnA+suPoVoqJDNcSqpEBbp
Jav1G+djbGgVBtICAwIB/obz4nnekbJpd01vVV8n1EER6e/tTLfTXkRKGCq7s111+WfrjpJS7+Q5
MN7paMyRHoBufG+bslbfi4V8Jh9qL1uYWuzlRLa4yR/k6E9rqgWMwWl3Q7Qsklil/U6OWIdlzcs9
4PoyrZXqNXrafe92vzUeGVvl0L1+VfjDUkTXwDgTD6whl8RJit2fWagRpLcllmruZwVyxdZbdLcI
3EVySOrHeirIwoTUPj6syabAPiowmHavY5lKD+uMuzkecmoNVOv7AExZDEVgEJ7xY4v+nI5ZgZHE
nploZnQoQPu37nteBrodyTq8CSzySLM+9/zzrUwRGoFiYVAPIduJwuD0/kJAebR0bCwKu/8NTLkI
3lz7QBh8rkLLKB5z549dGvkYo4UX0cTdFepJDA18jnmmKtZDj90unlK9VJP48gI5yLvfoom8EVmF
4qvt/gH+7UO9eom7rd1EaBAlt844slJAOC0sKZrxIxrLaK/1/jDUACPNDn8mIoNcofjHqh1Aa4au
uOJU42PwCHX/RrcwIF2LqRzGcQgFFb2MxqK4NLLPq+HBbDmxhU3mYwCldEy+GxbC/L4dupBesFai
8O+vNyv/rGTq6qJ3r3XFjm0+Oi3VDhO8y8CWXQQMn8p3UeFWtp/82XaGmitcTMqBqsW50BUwXEMd
N1XqGdDlESuOa4ZV1rJn+2m2OrQQcJJ8fsPELHAtpbuzhSm8A1GZwbN9K+93SYEUQbegSdmZ1vGt
2nqUDvL7h9vHtl4ee8y6h89WfodJjbKcCE1YZuKxIElSTtmU/S7XWgc+5YriLk+sl/Tb1qwFOiP5
ytPbjYP39mGBqIgAN8prTVepa5oAtYjaUNmRh4XyWh3koNsVdzxK4UnRDFtl2NchFhyFdV7YgOOS
VQFruXb/mFXRPTExB3K3zoHPrCfaD81dDpCjzmhHO5N1AmxHKnBv6kC7ABvuISM1K+Sm8lJjliEg
MBR8wrWjl8WYDUDO6Ga1BoNAr6WJYrpKnZVrmkQYffkqijEKZnMyS0exNMIpYgvsJX3mAYBxoc/R
eT1yDTgt6VjyEcOxJz02eKWwMCGL8B/vBdp7vfYAdOSbQ5pDlKxPB0F3SjlnEhvb9bI6wHt7vudJ
KD1bTHlc7pYuIqpFMtREZ7H4QNJVD/P06pIfgQXSvsVpFt+UHDSI0WUqWtSMBYw6C24/Nu6FuU6m
ExdAk2OwDyg/cGC1CzEIYtzDcXPWGcIbgEl4uSh9XJWmLzCiai8EBP6ZsEzfmYTCTIQscjuGzxPH
exnW0VuMpKNhyq6ObSo0O/MHvpIzxPhmfKxDSmIpIz5c+L/KAQLD34kmmbXC4GRBjhB4LermnBzb
rKZ53MpwCj7UrmYdYgbnk0pEbWH0NwBQ1Q7w1W6eoexIaKeEFwTL7GNNtWQ1DuI1W7JSJdjK6xPW
eRONGsaM+pyy0yOvG5ehL6YSAeXqrkMYbT7BaPp+EF+kHhA5oxz80kysT6jZImZLRESSWtzpDUy0
60FFX15A1gNvxjQF55NOn0+dN4hp6450tjS9sGmLSS4rK92MeBkXV6TKfZFAk5pVmHcRzVTK2fAD
EnLb5FhAvTGPGyBy8XSfrn/4VlHCeiAiFXpyhPNDKXKQBGq7QsPedfxQ92VMyKvN91Kfgfc3q21E
Qj8tZVhsmygX6A44znNk/Rvkr8SMC8V/r0qCEhvAcQO0HqlfF/ZWb1b/9H0rsJMo8IVLS8sye1HS
gdeLsWPMBNBHHgZRJNmjzsgXJJhBhDO4exlhUex3saZRs10F4rXbHgAozRLcnZYc6NzMNvrXWY/+
T5Cs/6+LTUhL28j5wiAiXfhQp3bBs9Ks5ZoAbLz5RFVcDtjUkrJKRsjaeCdQUQubXtH77g9IkgXL
fSnyDq9dAIFRSBOPoj7DG6t/8Ek0ZCQi/rs/f2i9+clLUnFPbj2CAZ11GXHpf6l5wKom6pJs87MG
4L/SAUTi9deMSxC65yKcFlIu6B5FFOnMMmIhFV+GqBtr/5Nsk9ZuTGM10VbJn5n13IYKmQsbzWvc
Zd4YQqByGGOrEnIuzwbl2r9R1CrrfEQjUbJ6r66KN+e9/CD+yfGQwjMALnE71W2ARmKK8aeiBfKR
JcHPDEG084YvPXDerX3bH6cvyU4NHH9aAi0Hslxl9OAwcyZ159aKmy4KogCOZFI4G0Fv12FXUKkC
FY/RVzu7wCAE2GLA2hFYQFlTmkoyiWceeiWLtnXcB1/schTyrF/JNHe6h8JVuwOj3Ta2KvPtXH5Y
UhP57GwEBqkhhtBwk8iUJ241bzAhCPWTetT+aFtiKJRv8eRMO2MtTnoC5HzBgVGz46cAGP3k4VWH
WYKVeJj2hgrsAUQksbTtegXsqA5mSZ+RaGGUF6F04p8fNVk77l9hYMw/8PjZK3bZxuukmX2/vPUz
w4ZHZqI27SRfOHRRSYLaknuCP5inHRFG4XR2upge9x2XgmR7kN7J71Z2wD712rBzHgXmmQPuBBBR
/S7THbReO5SbzHfUFhkZgrDUpPWQzeqoBFJjjBEWx2GBM5R7CdzTgmBZ+0wI20w8wt9O8qgprfUd
H39AP3j2Do8B/qoBvb6lnROfrjkTHr6LzBLfW0mOZZi6iReGq9pLmLfB0vvtaNqFbFnuzLRDRFpL
CDjKskbzbiiDUmZjXfkuIEa7bKReK4BNKpvFatoyC2ch9Y5r/gWdFeScQ44Wo4fKwdlZqZEzdQ9I
ZY1qohjg4PntoYknOVh17lueEB2IZtS/ZlmtvnuI8xmiZEndKtisGM5MsSjbQEwXLLM/t8HOn30g
r/4ewdQHQrvc2cluzbaJmpeM2/Dmbsk1sGEhDXsl12CFK9UI1XzCN0GR84joxx50YbXKnNe44EsN
5xTnahtPQyQ5ooo2BHJSiWfF+9PAX0BsVt+0Zvl2UlN50yhfiqDF9QbtBU/6WJy3XT03TQZhmYk/
FcGjHr7sRsxT4dU0zCRi+6IeJykVZyi4EQxW+dRmtbR8HJsu2+qsqI/ntNJ4UIc6vf1IDtZnyP+u
mu5dHORieN0M1YyoSukEKjP9QTmuQxgOxvtly3/J4no1A8fxljQWJlDMIM1J6exFeJA/DhTXCGSX
oM9Ql5d0UEi3yOxClPwUNRCIrpdwPVr5/1DcmLP/dNCJ66IuRTNqVKWB+LklPfXLZPhD7mEcZ14F
mKhNlq0XOdL/JBne/fRVZs2F3BMQlYTmBpQso2XOKNLf2Sy92fzLgBIK1AZpqCvwDP7ztTKuT7+X
SebcBHIIGq+xUmzZLPh7lTPh+apJ28HOlrDQksSYL6li+/TfG+1rnOjn5KF8lLcBfluxmw1+Kv6p
Yb7imUVK6O3E/8zpblziEz6RCRf7h/tBzh682RwsDZ6sIJh3NnGoyTnedDIKGNa5Fu+fvX31BsUi
ER/eoiRuUgWzcrPNNkS1f6FjOPlta1YdWr2w8mX6zVjs+56BXt7EKyhN/1ZdQVT+oHa4gAqetSKJ
eb0hAZ6216ojL4bHcUXC/Orop8JXKUot3X5pV5JDZjQ+bd1UeTzAQn20N2U2AUlM0OeGJ92xyxDf
3Vk04lfxh9SV+vggg3rXf6KmzLLarqPC7N+J+/cU8FHJAq48xHZlmSQ8/w7059MZir138PY0/90v
sLwJGioy94ByBPgujLR6VDy5emdub3THv8Y0O1Tkc4JLhqxXGrwgyTX7mLTsauLNsUqpaAEwWHRJ
KdqLvVZ6RuI8RHaLQ4DpaGSZYulSAUYoOtwDK84aT4q9BMbTqquTeQAqkyWB4BHOk/zH4B7rOOJQ
Bms5snJxBEneboQmAY4C+ay7BWywpk8oi5KcXKCCxK2/I5zDzL9o6Cdn8PXWvA9/AFqzwJC5gXhm
h+mobXBNDCcoJdD0LR6jmr43G1kVv2CUICntDsj0HDWm7YH5iBIqxCk4VN5FazQC4n/7qlNMHIgj
dByA5NDTfNzekxxQyML6sVb1qFE7IQV1I0y3ptJpCExQUrpDHpGCB0sejihUHMIezJHf9QuSV+QV
QzrDrhGBMePNXnIzqUpPxA3DHJbdvszzt0Mnant2JvBkTBhDV232ITu/pskyx/iY/Q06fKphyvwS
wevxVfPWemLA9fLLvhmTvtjrN44p3GrWC2KZgpy5oPs4kOLtKXMXOLG1MUpVU+EqsneQIl8Kvu92
qXfM4pSmKSD7M+P9O4Uwy2FVndXCBYbXTNW8e5kxxBrnwjT90R3LEPiCUw6pU5g9SilnGZ/IYxsH
ieTOA6pVQdeUKHs8uHwP1ypjRzCW6m9cWCGTBNA20fkfEv9yTEOphNE96lOlmmUcqlhp12bvcIab
z/sC8WeZRPpro8exmH426jG0I72VlMGOXsAine7XdtUlTnO7/6iENuFZnsMtczc6fzsEKhiKqw0g
BIVeoufatv5id0o6EOU81YS8v9Cv0nsFn272EK5MJ+6G4/Bzp14D4zvMzhZK/59l3bJk4v/giyxB
bX6v9XKyUEGeXuFH+R7ZlEbKtDF6ATz1swdB4XQ3pIQdrfk+UN5c08aqPwPGUcmrEZwV9gLMoWvd
XkEaX7u9TZp+9CkF1G9ZjPMKs7WmKKkcm/BASNIpzLhv682/9noLJomSPQq5TI0FGbnCPjjaPSRG
hIGGdxj2L3eJcUuogeWnCBQHLVBrGYiun0Tsnh+r84DQ9C12V8Upnr36b21XJrp767jzTDDLcAi6
XwvKTaYsCtsWbedMQrCwpUm32yARZR6R9QEWsAHFURID7ayPr3Qj2YxH/R4pYBMUe/avDzBypXVg
rMIFzd7dSGRKu80T27ObVAdeAutAkY32FWdI4brAPlQHyb7XFvSHXa73uxguM2HLGFNXalayqxVU
3Bg5nhZpwdSJ7DTQ8RxnC8pfQnnKwl/jx8wpcSMnxz+zscNF3ZrYccxFXTBp9DKkRfxbNPUqL9Gy
2La8MHTMg+hoMQ2A1hkYyNsyFGRZR6vRlpZ1JBojUefUE9BbLw6p7zMre1hr6p1tn+o5Il4FMDof
GW4ejrLTGFSP9Dyzf7mIL+U59sV5Lj8Z6NrQ18XIVLN/DzR4JWHK4UbFeYW7znKwBy8FE0OGWeyF
wgaGgbTrRGwXtlBIxxExXgxJjZ1UO/DCUiuWM9xmEAAJP4lbpzE5JZdjA8BlX2KP5m02OakY2a/w
mOIY1ptgLKmoRNEWvtl/NPlSKQPZcUsHpZOwuYpfxqoumk+t9lk2Y0q3chM2r2DAhngnZ+9nbux2
y/3G8K4rIkajK3fQcFIOMPMWGPrLWQ1Z1ka0DyToXtfguyAQeTC28A2McJPSjVkUjmPrU/4j2N/H
PRQ3ecWwPB/QcPy7k+BALfODHygR46okOihTcqN++Q60sLi1P8+8aSd8yxZKGkVPVDQY/gx9kqXL
XGz//ZuSPBNJrJI/y2osMtHTojHBK1KtvInw6+3yBD5Mu7fRhGr+P3wGDUepWq6lWKqdgPWtJGwg
MLauA3VYfV+iH2XbuswJs37Q27FY4cWjCHOqCH2crkQUNDAve3a9nuNdICX3bIfIb5/Ks+dgprp9
tBDODs7ycuTaRaJzq095HA1p0nALD4RUJ9eZIf2UEN0ik5uqKIYIkN7jNac0yrpC70wF8KsNrcFi
+uCUrxdYYSxwImmUk7OgkUnqeUlx1RCi7XBBl2CBzGbLyRESgaM67uY/LWYW1Ils7tFCIlLphLgz
8kYzZaGFOpxRM8cFlu88N6AWNI2uIfRkcuz5RfJLHtcmdYznbwAhtUTBngh5dm1NDxjEbIGLYzzu
UciuAp3b70bNZZ8IqaPV1bDgTVRT+NKGnRcKJsS4e/l7zSqpAuT+gx+9nT2ZLJfg/YKI5vm8lEmX
AS4bxbzVbsWHCTs1tL/uL8MtXLYUW1nxsATx42IXNSOfvkyqw5/iyyVQeF73HkmVdETTXu2gajrJ
7CUhE8wRdHYmHsws8xXxaVjxH3oTKHJx0oFauvOLA/06g9MhpUUV+YsolCdQCFMc3waLot/ZeDVK
H5jLjZfQqMD5L8qifufUu40tLkwcz5bSL2C7Ch3XdwBGfr8IoxnvapoZCJ/iIFDIuhfbIlCWoczX
fMzk9N/iEV+b5Y1udP5l1q1XjdKsttiTdOgiXZ31Qc/mGTsCOv+DxnbpYTXLSrTy07zgurx38/Ms
62PK3L1Uh5ScLSa9mUTVuG+ndkUxfvUJCZud8/nIZGLLGq6isagKB4G6o2bSVG+vQz8f5gDqf/BK
FTEGrtpim38QgUHbAdekq/GIbL7yJGjXjhBdpxBptVvwAJTsGN0QQfjd+VGhKeGVE/AHeJuSepbN
o/CkeUBqsYUumoGELtc+SUcP1yTKhqQxk3byGNbv7W1BPKDHlBeirCjpQbVSHFsweUupXu1MogWS
buT5HN5qG/EkK3sssf4yVe9F2XrKeXaIB/cqhHmC1/9w/Hjdoy2tzKcMQCr+69ed14tj/CUqa0EQ
8eqvygQXQIWNpmT6OpoMgC9bNvS2SPfOhrh3xlVx73pZspZbb8ElDmdjsbEvsMoCpKaKzkyhHl4y
FJ/iLzsWXKqkrRFrlmO27/vyDwKLvlHVNsX+Hi1PR3NU4g5tOb3T36C6UiGeV7Gbf1yFfriqewLN
UzvT6eIYU+cufcSu2pkf8pM/0z5gBpZvwJ8cMkI3zOLZ6PEOQvS6J+cNRy2guQRS1jXT6dikhjF9
rZQm/jbIRuwwH1oki0kJ+iUne+GVaEiWKxH5odKBBeED2h2vgq1tQAg/OqeJ4NqILM+6fGSAovOd
NnNG9rQmQ5iJVfqoFpRGmmUFwtr2uOnyOnTSnvCmCdS41eqhRjkL8pN7YPu2ZsHJLUORTH/DrrPh
y2BHm4b5Wxj4xrr/MHNWXerj3O86ruru9Bou4moDEJ9Tp/lnEOp5zMY72zWS43FTT0Qt9zKCRHFV
fi5EKgcge9YMdbIjqLc9pWvt9CAjcHYhtkHfIOKLGA70SkRl2HJ9OvXzjTYxI8E3bmc6/QpwxgT2
8ml1D8rIrpjo29NnC85tA2QoR8a6/IRlDz+KpfG+CHxMf30QwP+KA+TxMX29Cnx8aWrGNED1Q7yW
dAUa+DzXJ6ZFBd91nAb/J0VcrFTUObvS7hkbIDr0ZZsLKYHiE7JMqIletpiW2Lbt3d4K/IcDskTu
ph/u7QbgW2CX1RV1gisDCLQ0IzJB+FgTxyF/hRAmb+lPjLJIq7avGXQUQMdsCl2e8YecywJb/cTw
F6pxkg063KJSLPnspj6LrOXUOkbCcCCeZyO3eEj6//XKtiKantfLI1knEKErw5YSS156571udi6p
iSwDrMnrwxozDbvAqkkJA5B2z3LRNd1zc9YlppLwJSJC0gKMsHJO42EymQJx3KlgBAEt2J/xaYwU
O8jcB/kTzxArMp7WQ9tI3XP6WI/xQrEtj/oklXyXXqTYiz9HCGi6HC4MJUwd+WQwwtobe4ESgq3H
5EyyQBn+JtovuyN+ubydzvOCw9A/o7scvWuMJcVIHoQdnjjw6jUqY8LJlD/n9YYHkKgOk+c/OJwI
/52Z/GKxlbb1MndTKWW4oRkB/Quwj4+/Bjbs3XvdNW2Q8hfFpN9DiFkGa4mQnY5CXIUIRmFJMkn/
fiMLM1Hm7pfJccDNAhZVSXzpXKKYx9OPEEA0uR8RcMDaNDB5Vn3LG1ZAHIWj1H7xu6cJad8o/O2l
7aQqCBkJNi5KWzARsSnV3cogDmp63DkvfMaLNjuCfiFwrligY+4z5ijReK1amVb9xS88nVIGyVUG
eK/1Tvri6D/zgNvdQ4xDGMhXsBDdgN1DUpHxemSDzfW4jEhLhtkJSVnvY68cy31YE7de68uBdrmd
kYpoNeGJACO0FhxozJ3uCtAuoYepBmninQxr+oA4xyPJjC6g0ZInpWTUXd87pdEdD0UkqcF2pNCV
tAuEEq5QzJ6aB3WRoubrihb7gHLuvcIP8NWR/Ig4r3wcwAz5/osfHlnT602VW2REQsSzYq+ddqrO
8IlVXR4YafAaz+5/FF8fffCKZo6WOLafNvpDiu3t64Jx/8C6RODLTHndpa4iTyfmv57nR5qYvvuD
UG7Zr+Y6m5FQW4+LZv9w2JEFaSXB3WXW5kBNqBVqNhC0vajr5idOploaK00dx4Nfs9OCLkC9NLmm
Hf+BM6jvfiq4hn5KAlX2PWNcnmC74TgACVAOJa+fBbZmURwmSQYrcw1KWqi4UFAOcAs/qjVaRvKa
4HchZl8CaYktIPOn8AIDA4itTxr1EGQBLNIqoMUWf/oo+p1xfMJyEzGIAN3ihRIhaaQ9bRzSXrBH
pFdik/f3rv2ugRMTUfximRAECMWfcTsZTloYVZxIa+YfjH9J/ZzLGFNAOJvXkg8ov+UbEzDCgQne
K/0tHYFzCJyKZa1vxo45TSind3llckuTEEXF89l+QktEdXBBHF/TsDeQYB3MMCY/mxe57gDg8t+d
bM3mxexGX4YXFfxE1vpfn33WIMGV9b2wcku28XrIOM0fN0YC/JlIn4G+p8vlKY8LUTKvXFA8WWTq
TvCseJPNVtYfo4Ha4mZJotcIlFAjoNrcYG4Y9vmeUMXB9eCNHjlwum1eN6c/wys5QloI/zb1a1Z9
1UzNIIhMYIPnlcvVo/8febmpagJK0TaSucFtnPOnetUHoDTGp2o26/tPEnROp5QKbclQOxA+w4tK
PX4LKgHr42Y0UyD0HE+2ddgHjlIYILblnAv2tQZHICJY/EChbbKNT1vJsGl8vwTnLckAXPcaAHiC
njUfl08/OEqzn67UeftLDRfbUdbzwyDzcI3XXCczzBksS6lLc7BzKpJG6eW6qE7nmDpj/qcQH2rU
gYYsLrv3i0zKrfjmNPl3aDAfu2wKdEmCSxuLJVxC02ZsErrS5g1lE+xI85lvyoNhvMe+MGEtF4HR
CGUq3gV4OLcDG5uZt7D6RMEkF11ygoRItA2NCkmHk/1BEnBn5P6HJg6e8bwbjxz3Jn+hgB4C3LB4
RwdudvBfxEbCrU6pXA+F/OjGy6MdY9ivtJboUc3tZBEDJj/jry4sVoGor/VYrAPLgS/MgIWgZp21
ris/K7FmRVuc+Wn+upI41rfdxZx+05TaugKfdKk/hFkvJDQPSyuhxm+8O/1/5NeAhuLy+7hbN6Fo
Oz32d6WIa3akGC0phG/B/Asjxpls3NmQBQU9sp/6MkCzkfGerqZeJe9wxqC71GBNJ4a0GDW9fyNO
/jPRGUxVuqFQQm9Sz6ZbxxihFdJO52YN/nbtVKXDCodgIn2jgrGX5jfC36hiwQqZAenxmmYSQIGj
hVXpnVVkMgYD9OpAab8M66RVfr/TRnwXySsI8z3dGb3BbLVphv3jLq7tLtCDYAyifVC/YrfhRwbg
YW+y4jP0QC6N0+7pAwDVdnqk8A0tIos38HoJlEINHHzNyQ0aJaQ04xpY+d7LdOPAjrCiqSz8wzJf
9G+Czfdv1Kq7rbb6cWmhPfc6tSrnwZdOC9P8f6cqZIxG6hkT1qyVbn/SL03dTfA47/8GgFnuIac9
OWnBKC6TmX20R5BEpl43E2wYBiW4MpUvYtXjt1hUS3Q7LNJuoTmnrmNB6eE3lpaqiHeFS+BOG5yL
tCn2FRwRU7tGndUmPFHLvFPema53lDNn1VEsT+YecmbeuUyy5eVs288bUApS4zTOLorPP+QkYLAi
9lhc5uCnoxgncJFuf4A/klD6ta+y/00/JC0U2S9BTJ2X2TcpU+YQDCSuiujyWECkGHL00cXrmP7p
mYXu5UwTcL8FlXYYYddEHxQUylG5gS6sCXyj1cCr5HG8LF3akOu+F2+9zbCfKeSh/ueMvUVznhyr
e0E1K9nMR+tEFabMYr0+r2pStuMtGJizrSyTfJKiY1zbuurA9e/SBZTK/h0OxkQxNG1xA1JpJ7Gr
dPC/CSC2GJEOqI5NK9PYOMQzko8zaMWqQRzg4kzx2f01kFWwchCGfcWVrvq4oCGBC6BBkwQd9Q62
7LgEVoWeZJ8gOtD5dSxc9bzuqyXOmYlh6ddJBlaWAVupz+4iwMzhM1yI5EV3tBSoxer5CIyctSs/
pqM6RwxgeWNHKrIbgoVCvxBAy5bxpXpgLMbj+g2iGNNTFmpMOwLb3o7yTdouHnqVpRv1frVLqsy1
yF7FztaZDLLs0PtS8REvvdwjMt3+wwgjZLPYh7k1Gzo7EJpbvzP8vmVmxJZV4tEbiqTEyPFrVbYH
kXfjbbhfBEwZowPDybOiYfW8L2KJphh35CVBiSLmoOKWh5Rr5NcCBob98g6/YYTroIKMET4hR2qD
oJUTFZjX/cG8HKr1WbeDEFDPYFRsUMgiVc56I25EKRA5pKZlvlvGOJy2Lh6PulIvlOpwoLdlxBh6
nPkYY7Jc1XA+sc+f4T/3+JsfFYdPnChhQy7HcNYZVNaFz/gzEiAhTFd8eUbl43bgSDiXAjkIxmhU
1AmFgWMyQB8tumAPqK8rTsc9vzCwKpm84YPLX91+Nd7BLckcIiKvi+BqC/wgl47k7FlDdeK9vgq/
Ar/mM1CUU2CANIXbF59mgrNmR9/pAYvnd4zoIXirTIvRNUnr0OgSuEG/nLy94q7UpRznK/yj8inX
8SElEwBifTJ1EW/vEizoHjuZY5PnEKZFLbgfPrf5SJ4CNaW99iL1E/xetUBzzwBENxdjYCVpTlfl
dhIG8HllJtHOl4sTf6R220NWYXgZtbTtoYtCvWvIfRvO8tAvKE6BXx5s66mHW7MS2xA0M8H/vOjf
TwygExkTIIX1UJMQ46CHJ1XuPoNMF4V8LcWeEwBtxdXQCi48kcGulQl0CbrPgSqC7N0w0JENz7+D
0cs7IxaU5zJ/Ymdkpnx2zvVlgnVUIVrs9O7M8WqInfDhPROfGbGehQkLMlAqUMLOAfcJB8WRVRWP
jJeQZpBeHsFfNcl0194nVZQno5ApT6AXKqgzZ9NXlBiXuEMwpzOY2ldAjOle1hKIouQxZbAXR66a
6zKQJ00RN6kLbg87FZiqhlmvXyCUapYFbTd9u/9WzBr6fI1IOzpcgHDrYgUyL1f+6NQUPyahCxMx
y4gvBfx6U7C38rlyD+6e31Q22fB2msfYlud0l5tUc6l1eUqAkycmA1Zd9j7lRmK/fBV4aY/4cwrJ
3D1NYfDYITsQ1tkbpRfVkaumCruAm2zCJlryozQehg6sr2KEBoaNRILdM4K0QZuPGxnw65UJwPuy
2BpFj/rWmVVONQtMh+fky/oF2TBNoomFZ5Rn4HEutfvQuxHewYWlgsXgqD2lDz/8sswS/pSd9utf
po7W9GUw+uzN1mhyEzwRFR+drh4KWV4cXF6d1qnvRKel5BIbMNfxLgEDcEFGQAqzgE4XiqhOIuo8
ekR5PpR5zy6SFWNC7y2gZwHxTx46NYHX4RskI7jblQB3H1Z/+UQsgPlPudd0lwxhLlN8/asLqGJb
xGzobxiM4fXfe6hV2XX2S8v1aeFeXxEkBBiwwtS30F4wy2l/JCb85H5oNrjaOe3GUtjxeDT1yK5h
Dr9W1QlpEu/D5sFgDDKwK5hYqjbJj1mA95ertyfIPVM0awU56QgmTD+4lpvhwnX/3+8cBBXafBPM
VyQwyOV1mhnYQRgjIjMB3W1gk6LN8kPO31KmmSRpu/dU8uxk2ySXG7XO4LiR5yvSLD7iUf4r+Rt3
YiPEWTkgg2EPwVXeTbbwB7Nmr9QKpnMuWQYFVvHTasceJ+FP7fSAqX3beHN17JPq+p4UNWoF8JYe
TmVB+OkhjE9bNsgKsIpSG7U8gs5Jkso+QRTR8MB6uA5Qe1+WcvqDWlQhWNB72QwoqwHvMVS60FzO
hJzNXlSejBP9VMR4wlPUA8rc8QQ8QzYmQpRWt7QdBNixw3nhsslLGdal4PSy0AFEU22z1zVewTQr
V+6+IvZNB95G4qtcRRDZdqU6VjrOkhiCihocoDcM3uxQxPAjXpMQ6e4IKO83RnPEOcnfJK/Wolrd
K4jxQ3auaOd90Oi8ikceUaxlEVFYegcApm9Q5ZWvlyZznRQCCMzu6ay4UMxycaI4R1xoXA6uNrrA
9STync8i266eE0dxnQWwnX74mLvha67P7F+o6dT10QBQSc3DRB5bhKNmJZajO18Gd05CA4r/jVNW
+utIcgNqUXULX1EIlONYIdmBgn41OpMI4CBli81Gb1qO9fUMy/gvDS5v8q9uswauh5xHGBslM1y7
5ypA8u6nBlXYz1UP2SKWqTM/z8fvyKuOXb+vSJ6F1il1xYCMEUx0linBiynC6LETmo/+ohVjofJY
O5iioV0a4Yu3QP3BGG4Fm4FB3sl/67Rs/3T6l11/yXauNjVVQC2uz2757x5CbCmuY/Y2UYN4A5H5
PAZUSzJ39DfA9TKyrs4j9TeE8RaFf8jltrw0NSH7Ejb7JJN8f6SMuDgoM1l3qoo4lQUnq/HvdjNj
theDXPf+t1Sy6JkK9CAyoer+KJCx+NyJlvYBQpW9QjNNJrjBzdjovNwHyWgcYFVx0+Dl9aDd9fO/
oGjQ6BX1p27z+furKDjXkf+o7DU22gwk+9VEECgFk2EJ8q40vudVOCnCAUYU4DaxbDAEDMEUF94L
5rELXfIo9vIBP5HQGvEu83ksP6CEf209L57JHiUOMiDFll+drB9VIqShzhGlSLPe9vAl3pVUH3ZR
/HXVoh76kMCVG3XT7lgF6VpocXEujz0KRuA2EC+Hg9ek4PyKcVOnoCcj92FGn6iATRY0C53U1skz
q9ZoJqvKVv7anU9A0Xr2c49m+bp1+FwIY5g+/rk4A1rKwyGfgz/xFNctYRFXH8KrczgIT9uGxI2T
wUbbAQ+6Pqo/bp78ECjh9KUC75kY2LcE/QY71w1Js4mK/QuiORq6RmVmWs+mPorOf1XU4sx9j/xU
DxSCG+guUL76blgoKs+prbFw+NW4ElRrF+wswLJ8/N24lw0U7MQGKaMWnVECWJL0P2erotM6Pp/W
hKYbxK3GjHOWZNheaYwFyNNoOYLf4P+2tNXoLef4lk/EoFAO54ZkNd4KCSSkri+bJarhDp909mDv
G6KTt/Ty3e9uE76eNsR8j2U6jJO/mFC+be+IWoDFcytymB8czX3LzD09TOThD7+taak9CEUKL+td
xbeF8RYMU9qTNJvwCndmWWw5fgkTPEwLR+etOo/Lq5D54EpYmI2MttI8Bp39YYfogPPFDnJKSD5z
pEX9Bj1tsjwoa3uFVNL896a3N22grLgZ2g6g1yNZmDSZ9nKcDrXIjYXD8wtcYvCfbSoyXc5w8nJp
QKWkJVhlZ5fcMHWrQX8e5fyAiWPjmZSh3G1nRSvXYi82WjgPo9+qhaaesPuDOp+hXisQV2WMrANp
QWMrl5ZtgLTntfeK/H39lvQ0lz0kvLV4I7bVIuQd/7LaHLx1j6c5G6oS0WKnMhLTilA5QLc3Ja9c
gshNAD0S1QxuolZ5PYY68jqMHc2ZK5fJe1yIfIQafSnmhPvnKoULQU7/MGlWXFp5pH37O1ssWK2W
5w3AQaRQxQTtS0BkrGdVc3Ri0ADIwhKXLrdPyUmA0p2Wq+Grm3Yq3wUsEb91gqL2Ov88Z0ST4UXZ
xXInusXNw8/FMmIZybwUK+k4tLMCwNauKxpiVW1Z5Fo0pIpxIGEO0x1LB8ijVJrhrwjTGhmTONoU
8OuiIjXm1rIXgpNk7yzheUahOEIwIJdmMY+KVvxssBbaWW6ncZR3fxrXSJ7rS28I5AoIhUC3YQ5T
t/68Ft/rcLspQnKtTbPS+DLMKsaPiB53Or0KEYp2fyPTRkt1aHPXQjUlUZQ0G0pS1+bnHa8+AgRv
k9gkIev3MVfCvYL5jHOPp+RHzTT7aCDHgz0Tq2Jv2ks6gqbNjPeET0RdFcbjxrSD6rlm/1POZGaL
NYgeAADgtgb3FNbmYXxAeomLDsBkMS2CRcmytHfnnSXFCm1MA6i/9qVozt57ST8uDblLzy5Kgc5k
przS3YMB4qfZrT9UNkzqX7hgQFnDp7kUq/A2Un3bWT5QfneS6e4PoD7AQ4P4b1lpqtNjjJ9TR4Oj
ZbIXDFijNdMaeBykdmGTnQptUZEVJraTm8tqF5K12kJqP9G8xhu+Xd7exiRRvjH3rR/cU3r80tjf
hrMzXIwHPqVX7xSOwgbLbvmrWB9iy2F7cp7qutkbmzr6O19kcvg1qmsts1BJtAf0625aGZJR9CpE
XStsJs2U8wOBPrWIE62xxdpe2xsjbmBwg/iZO/b5Nv88gAlHysRAk/EkSNQ3/SC7rDf29+JmK6tF
rlcdRZVSNuePIMcrgFgYGleLxS1wyVYoUY2vCC1gL6taugFiGvAWbvozfz7VLGxO6qavKjp+wYJK
PIyrz+uQ+fQq6g2dI0QB2s0IxmAsBVREFbYPft6n0TmSVZOteXalAaYzq0OFgSwt8jb4iGGj11Ho
CL5XlJ5DRbDD2xT+QPIbuoSfBvKOx4cWA1e6ZnLsqrnwmvWyEz+OtPIydWIxnPig9za4jGkWkwE7
d4PzGubfgZOt+Vp1fCfCsET3WnDVs2m8q0eBpaRdAHNDp7ngDXdsYEG8ougt7/LkUG4JxiAUiiqv
V57PXb5eYiPk+hcwKQ0/aRPJ6h0hQnOF34mdC0G+3sDwBDBcljJO+Ihbna6X1OpkXUjbRclSLQd6
yGWFHDsCqXbaz8T6+kdR0cR+OEpIGoy0MqNoQHwpFEG/tEh642reHxGpTw2yMN3DbRiXebTGkdaF
uHT58i+7PkNlHvJwjMTwjC+KiQzq6dgQ95XWN+KeSxKR3ZWFBzL71/HaiZzFb2iH3eM3UmcdtRJI
++IZOZ/y14AeKtaa0KJ9G7w2peljt41Wqkbls2gazvlFKml5BfqcYEY5Nrxsuf+n4kgBCF57/8zW
wdt+bcXJIDx2k4uXPqh+888WAMrmD94EdX1WA19rGOP9P51cwVIemyhAj91y3dHCua5b4iYsa5fW
ag8sV6CsI8XcV5z/WHW+mT0BIQ80HKOL5O9C+Xj/hRABlftTdSXUgQ0LzxSKR+Bcu7Idru1PyHpn
z+KPHfPDZvZx/Wu6ehGjtGcCuDsPxZCqac3nwY/C5ogsnvwIbVbJ3Q9kt0ODq8VeUP81p2x/s0rC
7LYVdpo2L/icaWaHNzUrWGnbSQslVI6bqOZaqsadzHg68YiDfrzlUtmXOEHq+dosGgiRrrRaYqzE
8Yst32mfoQ5DHdgTzssGl27EqGhisNCgsoGa7jjS7rcibCh55V8DLZU0PlxTZ6zYAkS5Gj+WS6lO
8jHa+OmzFnh+VOPQ8aRnJh12xyRN1qFZOd1Qg06Wykun+wX/u6BmnYjb0C7To8ixI1VS1vRBMhuG
XU2xiRI5YYtu/HUTL0+6nxAyuHWxjiFQLePqZ/q1PLS9ZUkcWekfLAIW6J6U9YliP5Las/KHbkQ8
/v9yN1NBFJV6o1u9+HlGC7+qBbsUXXA8qR/zxf3PVsxY66l2GrGmv8qmZZyfj3iFmdiefyWhEA2U
vxVxZilhXXq7FvgZevFqIg4E7W4i7qi9A6wYXYVb2Op6Ff9PdkJaiRVEAt2S3bJrf+Nrnu24tt9y
0Xq0ddCVk/PlWz+85CrwLuNNa7/Tyxzs07W2FQ1ShFwRs9Y1USw3JtVT9bqvlOVo1UUqLhF+QARk
w/znYYWFzTbtNMUxM0HCwmnRtCSKbCXgmHdOmyUCKARbB61pXNgJt0ZfRcnz3q331ADQ5oBrDPiy
hgImLYL9IZWxxNygB/17dHsRB31SIrbMz2soGYeBjWCInj1xKhxnPk6lsZzFzN0eAEIqZneXDURf
g/2qiVVklpwJaqth5XfdYf1eOCGryJ4K+OYRC/9bzaT1hoEeCbAoh//r0wW7yH8yc7lp05Soxqnd
gVgp7SXvW/YChNFhxs+znf+YKxPEUwvXSLJWIUEnjZ1rdbDtReGG+Af2U3H5Vdqde6SsvGyTwl1U
DkwjPViy1CIe8F5YrjImUQTdTFLnHzrzccYJK6HSSbUEZN4hlo0BnVCQud0PBu5gMmpK99p6M4dr
8fafAMfoLa5Iuzr+vxsgDw7q+6lnOG7vyvFliin8rdcb3BrZLVx/MJsijMikP5JHpJZkMmiXp7j+
0nInwlwRLRLAzWDRHtd3l4i3tIpAFbBMiiTRq+XHYlT/ucSPuoM1juzUgqq4MxOspyWWIV3oh8Y4
XfySPycS4kGLb/ksa72tB3KoZho098rz0LqJWkxkfzRHJu3wXoA6YlA84VhXgFit7B2It7znWO+g
GtiJODTvoHxUJ6m4qB9hzV31zTW43d8C8GCkxoudmfhhDf9njglEXmkDnRwqUYt4A1WubZnFCRZx
OOmo0oAP9/mRCVdLbe+A2iCCQ1Ty55GkljoF/yrjba5H6C53JKZfgs52tcZOkAfdUJl3GR+l0kzN
aNAa8CzmvvZbRPp1SPfbj4O3pIcsVxtktp3ra8XgMUT3GdO9dFljl5c7yBVgNMhhwdsTi5Biy+ev
RKTTXBsnaVIAQTAp3Dmycg7rJCY7IERszcj3tePQEwtQsEXj5orYX8PNhwg2KHO0YtVtxfJM4gdo
rqf1a+IMEUphhdfYgIMiZUkViB3eRUSh2Au64t4lLgAOwicx/ky8aCL8EQMpob5u7wDvb6Tuzvce
09bB+RZ3AdSvXWShe85Mcar5qzkJlRjjbo0z5uN+yJcFSDJQgz00YLp08cgsUcnm5Sh1K9bOTx48
q7lA78CL7YwlFPQkVdOxlrADzrG1IMUotDKAbsD6g195E9/aTnFnCfVsvAkU6M6IhG/3qdda7MvA
RBXi+UeEwQmAKZZ1jFBFEovxPGPo3V7XnDbRzLVqFb8aXG+Z6sPvYolMitoUF//QYSXbojf4O7CJ
4HQLUE1h0x6M/qd29ETVf7zG/MT3D2OP/YWzjrNIQ6g6kd/zQOi74WwsYv/6xbA+0cK2YGxwWvK+
JSBKf4YSVgkvoXGGUaCvUXsxXEEQrJeAXOljxCq1AVazbSgFrLHDUbvtB/ao6AhBs0OVC+Wk/l2G
hQfuAoC2SGOroCWI06HADIX7CvfuajAl7iufuLXQjNYPwShuui1KYud6lpeDLNrcVTtUnL6imGlx
1DICOD1K+LhCE+PtxGHw2dIh5kB+H7sH7mjHwg1wmx/SXUvNKM4ZuR0+hZ6R7ihuTaIBuWK9NioQ
4k4LCZb30zNmS+2AbCqvuf3Pqu+0/oC1Elml5297b4VjGulvaZp48eRz7NnpduEfHvclL1Lt6pui
EFvJGqp3hZ1YoT8188+/TaLxJIdsi5clpQW08rWFPcezfwpjffrBjNRC1QcTQ4fvyBrpZVWqmV1f
i3x8oQ2UGT/hUtdmQ9JrbVXyQqi/gt85Oijlhcv74I3WA1n8aRGv33Eo5vRLp+CjfyqPLPky6sXf
/coEbp7CpYuue4S1dqAnailGCriYxy7HWjA5yDijrkdP/Zxq7/Q7WEpZFqEW1RdARD/QefxcoG2G
dS5Hhcf9730MthN5Z9lLixD4Izm0o+cr+ITnv6kUJuqSkfypj6L15LEGlB1+qf/FYPc3yT2ujJwL
nvljWc0lxzMwzl102nD/ZdXNNKOUr6uYmTMaDh6PxNUgD8MHSaNP0qSU2a43MtoUkMlpOB6M6DoG
8IiRvNhhIQDL0frWNTMr6MszVMcuGnjZRMb2BTLlB62+iCkyOq9MgHgkw2YxbumsS+Gu/GFSDqTo
RWl+1XxHMSd+ftQ7AgxNXivH4cTu8kBfZWCbifE6KDhVEvGMrmWZmjxSzkOi2er44c63TTD8mvBV
qZglLZAv58mnjM9R/MDfSQuAKw137PErR4vP0VbXC0eE84xK2e0wHmio6rb3TxNISbq5ZJnBfGpo
745m9PT61Z0tCMJJAlBRsGG8H8Q0j0tNnEay8j5BuykMVVrWcyVV6WRE+aLRbGb3TfOjS61FKK36
wUCZH8Hqm9LsCBXmqhTJB0OLkCYx50O2pg+TtMow+wMgZaCDJlBQba0IzkoNGRWhSFY+RBPJAQ0T
Cpqxj4uM3qKuIUb4mpzMSsOOZskVqUhZY3NgT4gpn1E/u3tNS6lCxwV+kVRGL4r8yYxR/HGvGrjo
EGoyZdC5emJZSTNgLd6cvv0RySSkREXyH3nudimdMDRm0Sgxs8l+SHl6ZhsnwWfNCnqDXm8svs6G
cAtw/YiRAScGrA8A81bDmBDlxP+J8nd1DnT9JEjMICT/9SZg42FtA3InqNktPlg7ezxiYPo8Mf9+
y1OkiMBD7D0VO6HabS7jMnghg7bte7qvp1QnvSn7jevJ4BUlsul0W1gPzEkI9vXDYpwhPtjTId4B
hOga6F6Knpb0ixGAAyAUEhRvquZ8eCwCte5FkhTMqIc3CKEkkl5rTvNphuqI7H2OvQgKW4rtAEDL
H2oTKKeVYxyOU0H4uqJS4OVqVHdej/1JrKOhbOL0yn1VPUjN7aAlwaw5RbOO+2hWW8n/hEglzxPv
n+XmWW89N5ydPDjeOUoz+IxwKLwNcX85+ytiqqrHc40Yoq60NEiw3Jh1zj1gYrweriyUHWl3S5IF
Pp5p0e2m/Hka9xchbnldgMSDUmYeVOv/1ivhJ+PP3Of+oa0KgQ3HLQW6ePvHyWO7gnI3+XLDOHuz
Z5t3tFLwQsgbagYj1HZmOcAOuZj3i9XBlPnt3I7Yn9zx6K1u4qKJvgAiPX4bhWu4BI3j6ZPDtBh0
qs6IeBEttmhozxAYhTaZwksoQS+q3YG5wqyuRHV3VfXBZI1vh0pOgAksFKN6Xflhzx9ERCyWWWk7
cmpHIczfKdSupYFbhXhUA5q0uMlANfJkDQNiuJ73Uaz7TzuFU4FbvoZmFOht0fsRM3FtdKckPe54
ON8/DuXiPo9MBXm8TWmlkgzcU8whfUFhdMtKdbX9P0ZjOOG4nHKTRFiKsvtbVlmcpL46wYC49QwX
RQlpU3o+Uobzj8GtdCN+HjBhBqN86WIvCi2W+NbuAd/wL9A+Bzu4flxOE9xqiiarc5KOX36kCOM2
812C0y+97dNL1JnCSqVrkHk6FK6+oItW+iT7DGazwt4T2243lEPwry65iwgf/twTufjN3vAhaOYK
PQAhon/wZsnvr1qjMqTa6Nveo5/ZWlpAybRhkgLT+cpun3A54Dc5DrQEL+FE6+hm8UlHJeqhmFyI
fZKtzOwJcsmGvq7NUPF0ULV5hQfINdmnnbmWXbFt1nZyttL1rOIcfLSgT8JYcnZ1gd5jDFX+440R
W0n85yhdZ2LRqUDDydEqvuVc7+pKwmZ3RbvM9q9+O+JywKeZjJZin8XzxGHYmbFfRBX/v1SSTF8E
M2SUxuSGKgCFE7vkfiqfBAfXv/zJ5PwCN7xFPI9UgKlKe9Z+wfmPIxoZi72R4VHnk1E8cyF6K84f
yWU6nJKEXD8Ts1egON5Fn1UoGU81+u7vTT+EQ7mSB9RxuWgPGTcwJQ//StrWFgcatjHiQ5ltxiRe
nMTCO38dEb3xxKWovnCcK1wKCUhTuduYNXLqEZ4nEmoJ4hbK7mTvf/84xA/2QA1ouZYoT1nrtqeQ
CrXd7F9oyUGQ9j9T9cbUh0w5fAB6i9eyEB6u0Lh41pi+wiXON/C/+S9QCdhiLmdgHuR4jvO0ZcIg
W3h/U0j7cJwqAjHUhNzVk75ElfXu6Kvw6qBo+kUCUyOFeyHmKsbwCuj5RLFozrjS67+JXuyERZLH
IaHNToHNHjIUlKDnFpTTRm2AjINWv0kb80e7OhMVHkGaH3N4l8gd2HzFsEHDEYQqL6axKK9IqsTC
bZMYFejJDjrO4WV2ytjQKmxYr6YNyM0epKJL+0g6fCLJTnp3wZAuzpH2QvxTdvsqHXrtqVOcxIJS
AeD2Kvm55Q43uCcxb4Zzcq7t+wStj1/K0cEA5GKFzCA6Iqf+6Syi+xpxQ9WHMg9hAFgmBVBH8yzN
lQISmcCyeKjObbNjPeiWD6ZuBj9cAp1ULC1KmAo4bR4xcVFi2zJNe82Be/jiOnf0OqMS6mCkoOEL
0wtZH0SV3a/tnSV9ppjAOKOtNL2FKnUpBNHJtP/P2MpGa7qD6TbAObeozzOGeiQUTBSqc/lKEuJm
/CrpnmignWn6e30PQYX177clQjq0VuaKDsUwkZiq6/AVT3yAo4q9n9WwcL5BXyg9UVGVVMVrBuMF
Ot6ydgr+mesNu1/xG3WmnQVccx5a2hNTAmT8KuoPIaciAe9EwuD5axcBuciBpLlpkwtJxwuqZKMc
6K8DXU0bbhej310mVJ/g7tcA9pK+CMxfq7fZiyV369+EHsJl8omdT4damDd5hyUNxXE90Kh2Vy5E
mlnhi+L1JlQaaHM92fSm7qDGaFG+lAVnwATJTn/zcXLp6/O/PWwDdYtMRrL2GtZ9bjas6qCvwZcR
FeUA23GfBSoac1jkwrp5uevAmNEXfMZ7HSIGrwJk/5xVFljvuD/0gXdjwpTBz1AmGBh4UzeiGImZ
8uj3vhfDWZH8/HRjmxXTHeqosM0JZDZfF/XmPLmMHeMlILKQf4EDMrPipxI9ZIjkxM7wwif5zhl5
E5dK+RHSZlFT1CmpiA4+dKWxZePNre25YhymIidItVX40Wb/6hCDlKagZxF9ONexjPNFFng2VHkL
jpGzZJ1OH6nt+pm4WMM9woTJrjCEPyk+S4++9FgLeWrlkndX3XkRefWD31jIZEW9KEY1idmK1XRF
Nm+mYzqhWAAcb3zxDckh6B/7l4je2Rn3nXr9gU53ETcenYWpvpOz4J3bYLpmzStMWM40PBOuJThm
VhOFc6phbvSsMvaBkg+pdENunccmwaG94AgczxY2aDxZTSCpGPXGrkDXtXfHuUWESG+P7sl77QK5
GaPwZZ3gREXsKHlUtATkrs7m/c6sw+hXapcSN7+IYxlam9NSIFG+Vg6/wordv9KvTwvEKRltPCO/
5vG/D4uUy9NBUMY8D8F3HFiF1T8LzgDDAz1YZQ15xfmEzFzmQylpEHgCmOvW74+qxRQyrSEhGBBV
i2F68HWP1bDdMZ+LIHL4NmW0ZYsxpThdHcA8ab8/VYqCtIUYM+4+k4t4LBEedc7JK++mTL6kqRAI
8F7YHdGNxbcn7RgGUy4so2SmlFrlGT6vuukNe9QwEJR7eUg6sMy2QswPjia0lDDjyzQujU1Ad/z+
7qUhzBs1AavACLT7RF0VRa+eXmlNXJqnuyScc3OQPtvN5jjCDhWJq256jKQnKvds/2Ox4thLZeFB
WOcHOjDLkBjPXFdgAesigBH8mnrEQV+lD73Brb3K9WHyeilU7RaF9Hs2a0hDTArdhJCHdKia0BJr
XIt4Ul5e7qxbaKOpsA9+2s4vk2lgLLc/Mbuu+7B1CPTIXODoXEbD2K/y/XRpWo3LVTpbFd1I5Trv
Bi0aHgxNQAXeNsUroAWNUdc2sPSYXrULvIE67P2/PFAv5vSt9zM7id3nVEXhwuACf97rau9zs1t5
gGeNbM4/MS7750mU7Q1DH/kwuPf+7E5CvvkikqdEU9M8C5XenQOCMyzCzaDlpU1/BpnXhvhS8BDa
W9JR1WMLNNpeLEuKRAsWVGxsTaWwu+e6tM5wsgTzDHJF8Ue4vd6MN6RRk4+CO/v03U/mlbCYl78J
E/5jfvZ9QUyIZdDqX0mvyKX2VkEDykCc7mqXbm35fkq87quafe4bAqAz2WrrQ9OdzwXpuiUqYiTV
FemPOmKk2GCdwf/Pje9XAoOL55v6c/KO9IGmhmx0gve2OmLpL1Nz/srCaxL5iUZqwX0df8kwocuK
5ZELXQC5ADr4pGjgsN2wdoL7IU4jl+BVz6AdyVG3Kcjitg9MAiLmFZWHW1INVBa9z7+IYFgu2/33
yeQOqoOIxVEtuD/nD08D6IbOe45/JPq6EYYdi1ExFdiOIbtLl51nCBR4p1R9gFfCgjGUQfJWdocx
awRujeR+/HmLnOPICrTXKfYdEmpFSK6ip/2gPb+l4UtyrLm+dqEH/BSzKdfjkIbikyxa6yX2Q2hK
GTL0LHQtTf1ycLXhmBIN4NDjL1l0mZaQh5jNgabrxy+WdPdrvQ1sdszmKi8tmaREx3gKbDHL9qvJ
BnaMJdtS3iZZ0OCJ1emo2rx1+vwbjdW0bV9RraXNTwZmw7/70ltxw43gsKoCarqAyp9fbh0fdmwD
H+vbegIiMfv0klKG8W1UkR7g947u4VWZCtaGsARyVZyslq88WvK9u5un9sJCKB2zHNcDjvQPuSTE
Dpl+hKZfHmJ9lfRYQXRKiv+9atq5T2g+ISJ1yTVRKgIIf96IX1zgoypKYf6+nKNhldp+AJjnAJmh
e8wFt2MeKSOEN6pPs6yXW4mmTSnPw1wipvAB1RQCbIC5RB9EB7dxHflO8dQvqCrNWQUEZlNPwMcy
vw/wuWw3vRr//6LUgimpLLb15t1bEx7hgtpLnO/DA5k8YtJ3uQGP4PxXiB49wWCxuvRe06ieGkdU
c3LpYZFDf9GgMyD8PCODTueKnC97GqnBkPAbzflrXIyUhwBXujYsHMB/FXN0pg6qrd2vZYmHQ1pZ
bBmfFtKG+Dg2EhLnni37em2dmevoUPAupen2VMeu69Mg3mD2vSeFccatUTOl5Aje9cG5aC+jDpLS
4Jgz4E1lYg8zjbC5bYu6wM8gl7nn8f55cOU3RSz/E57L3ErGHLE1WK4ZHzF76z7aPvVBVxLiXO+n
8TWqoU46L8Cpm9uBh8fJTNCMHWTouz4a6Oo22AMsA0d7QjrtvZpUZ967yk/PWRTN07MpjDXBaeXM
rqcPFbfcoPBciJqLxAMJuQR8/9wJNILn8Jdjl19KHfXCeDqp6JmoX7LKEI1XIhq1/fjJ4zW+NpOe
1+3GGnccdaz7oC91fNTdZY0XIPk5LUquUyufiN62ifwfso+fpIKZyNrS2WmxgkJ9+9TPqO2AUgL/
mUe9cfb4qpnrAm3tgBl7GdVkVBfHi7JvrqSSVxvVgZsU4tiB7BxidZv8NkRTaP/IBI0IglECbNjN
MocXUZCuyOWlpJlUrrNnqbLwqPNBEG+mq2cJk0lp9qVafQHIZLFMbTYVlNSmYNt0gCGSQsUh4zyS
+WET6R4hv6apOadZt4py7P8DZKMgTxDsBwumJXCd89bwg6m9Fy8bQiAU8pMPej14YgDQfHyjWJFr
nxzxNSl9Ta2vnuQWac7gPTP+WoN7Up6sAFpZVsyn4yAXjDOYBHizypoXH7/3MkL8tZG09Qv8bIQn
4jkUIi+YtCfCdWYlQeLtAZZJDNwG7yUs8030iyhLPH91emobGk13qbI9VW+HhYNv5wVoyYTbNzcy
BiovkHaiErFe5XZWWRMH6Gjq/463qsfE1TiNTefettHCeLmivhJDnnjmQQ9OS7+j2P3JEyXb0y5J
uZDH3HXdXydr9C3vRsF0WQy4SVRr2gjUqnBGkVRAvO7IfmStDfKSXBuBSgIPdssk+JH0M1KeOpdR
lb2ssKAxmwmsbhXdgNtG/pLhQfX+C9+o2wqCynb7CzbaCbQhelSWZyF+NNHHE9Sb4solm6x2tiOh
0pZGcJ+3Wd4OB0as0+rlYNZQe/UNTx72m3DjcliuMI12+HcBrr5C9DpLNKF7+ag/cdazBxmro1TV
rNpq7yYqHmxF9FEuy5jX4DcTgOiEu+015lP8sMDivwUUaxc7wyxuNsiyxHYsQ1VvoDUA5McX7heX
aiGRMM2klQkI/qFdYfm6Zq4Qn3CDwjyGf5dEvjcc2VH727knspKtAVAxT74pMEIa1RVhkxy8fo2X
P3vIimRSPGI4iLjBEMg40vPRJhYvSQ6SzKardcKHhoah9CaVsM0ICUghp6Aj1aVAadkXY4Jvq/q1
UfJ+DI6lLWM5apIbAyacN+7fCg1LDl3y1M8paYJYfrX3D2LQsl5Skcl4rCw/2ixAS7MNVMeiKBvo
djUousr/AfYXo0/UjD9yMfiydc6mpwUnFHA2FwK9Sd/hQmTmiNoNWow3Tpt625h8ApxcyxzolKAX
3Al84HLp5w4lpItY6PGkBett3kWwL7CrO0hMNwATE6xM2fs35vEhVVZfz9JxkGGUY110LoCCUVu+
aRObeb3swBITaP4O8h5LezfB6O1U9+G/RH9lFJRW8xo6UQiQj8jD11IVGOpBXPmi/oB67NBn+LF6
ZPA0j+iNnZFPgz8vnEpducq0pqkloPwXu179IR6aNLI6IbCv2U4YiqwIBCvuASNm+SqQbetfiigm
JHrVQp1vcUVqugeUQpc/93v7BABIz+gVb51yw4KRDW/MNd+lg4LawTMK82ef07I9dGyj5Hx7pWp3
D7DSJJGSsTjlGrOWUC3uncXg6XVIoVaJqXrLiNx27+kqKaGNMsIx9NnWYSuVmXM411J/H/zUZBmf
vZyx3YUuZaMXbvhaUyfo6GqEoH3JWZS/axqAzaE4rDk6OSfjtXwmByQc0JBsr8F2Y7sGysBPK5hP
YNqLtjcyBwWpM0sPY+p9YMjLWchIsOwlf96ha+wAV0zDtWMH7ZY6rHrM/8npzDsDWwjJorGlIiTa
oQc8eWfSNlxq4zEyeRhC1Yp//IlJtY8KLeUbQ7zxyfuHCUFhJX7w84hUAh/vlb/caPpFfDO3x9lL
W8p2bwtDb8pqcvISRYFP9X6vSp82y7kcmjPcPrhVadFhvmXRM4BNWw/SVBaCZ+kRijkIh4fxIf5Q
tSggofwGxDYieJmlZoFdZfCBfdM+F/rMNeGETR40bfSd7a8LclPRbkj6OrxEHeo2t9NyYuiXJGQH
Qee4ABDqPkC5g7iwFaLP2HPOTeUr6q/lRzLbkVHuzw92xzbDyh6a9WiAWcvnP12RZIOmTkxBNm3p
N9Py2FUz6nt1n1REslAJk5WPDoGz9I34ELxg2IyhnKhDJFWNPZ8+E39BtrwvAlQFTYhxplyjlx0f
eWgb+D0lG46Os1SIsgmOOioF0RY32tey17dwZFH8M2w0dMnAn+ChPhIv7oLcWrurAsYDQfIWy3WU
L7H1b1LmMeXM+7oylg3Gh7Tbs4siCfdejL/7vGJMxDElcUUpmQr0cYlr2w0MD6ycHcnxAodRSEO8
cx/N9egFlIXLM/2Ig3zAVPVzOuxgSedBcu2Md0meRl3ad8G6/JTAaHeXVhpA4qbW6RFReKObTbzI
AbUWbW7c3g1AKB9/B5Tx1LtUsmF/SoQJbftS21Q0/5Sh1Dvqj8qxNkApxkrqhE8NYT8og+xt3u+X
KIaIaLG5TSzg4vvCoBqolhJ5nkwBA4K2tEwAlQa6Vj3oeSqXv0mdZrobb2KoxY4LZ58taEpybRd9
WjBPPy7lILtgccyFChuet3cPP8lSZf6dn9lx/mOS9svgYJ53+99lvz1qIVUgjd6vDdPK25+uugOV
iT4+IGWCcOblnrO38UsofXn8XLOWxvbwCEyiE1YixDHkdlqvtoI0qtD8y5ZaReQXU57e6C6CJeAC
EpkiQaXJStEE6FPs1Y2Y6DTzfUzmNyKzyHzHiNNXJsEpytgfp90zcgw+UaffwbgUp/96psCRBesr
TStPcw3hZUebWWroIFEL4A+blkZxO7F8Xuj0MBLgvUzRtIZcyn1FqNAvI+3W++JfMgDdALlSMh/3
4eRe7IhUm5743uSTHw3m4qqiZuwW1gPTknbavFwKp3DZasaVDpmG8eLM9oudIhPdPwiRmq7vRu8u
Od6qt5RLvjqPnNELrMHjN95LKAaOS5LM/XPDhH7PkKe3eqJsnmI93Ac0Iyl+0QNlmi1ar6JCGtic
PrAReZC7Gx0nFxviO7lNIYCdtkzU4L740X19wem7MCBrGuZz4hxycRzGDZIurxSFkTLuQZ9CcVTS
6bQ3Ip4kGlnKmsbDCosfa6db2FKd28ab4noGKiRgJf0uUgqWvtrP0CSXeenzZWZsidRzAf4LoCqA
7a9V4mFqxU4ys4er2vzGBjZUa1LjQnfWJ4yj/PUcKitIR7W0/ZFrXH/LyDi+/0ciolTj1tIPKpM/
ce7a90GqFngzfZaIpLkzjwSZDEtBamesKAPfvNdbNKJUVkLektyd6ctYJLESRqMYUyTixzHOcr0f
Oo0aSsKJDxK3kkbL5QtqsfFy5hnFeLeZ6hx9suo2gNi2E7NixGR2qGAHWL80K24eOiDNhbQ8CC/8
WxsyPYB4vU2TxMRi0cDnpdkH+B6xL2yNeka4BPeZK+Vk+lfLq+DZxaqj7lJXHC32ciXYqBZ1IRGs
FdMvrtUEzzFJ5cPiKkPqJqzH8UuH0h/iZ/qqp6vUcDXE4f8fW1dOhna0i/Nqcf6pT4rwWemOjXrz
//djwDjMmPARxG5uR9+e6ddzMFylwnHybKPe6uorQjrA1aEmQJbMq6kMpS8+DMcUD9rPZsvheEtZ
haoqfpVAZpOSlf8FHMxbneKY2Nw0AQPpDRN/RPq9Uy7yU3/Rt3vDhvnKq7OgkZ8j5WW5cVEYTDJO
kS1ES33Xxt5pEvNzVt7nFr+CBJ41nqhp+8Gi4+SeXLe+F5yjwhgzbw8U4bVCgURWZPUtYA/kQY7a
Bw5AklnZncsIdjbO5VTucUS+0BZ1KmkATXTVoqDyZ6tneiVskwUNE+Hf4zerD+xlt2CoFssXP+Ad
Zb+6xgLxSi+jbrwqMyCV76/53CnhbUN/scbPd6jcEgTwStIMbIbLFwi+TUxZsk56IL6L+HUvOxp9
dkJXEgebFul1OB7oFChPpnR/49hal7XTu/1blJgpshbHkXMptDRgeI2wbfXPdM/QWyRifObMIKoJ
nrbqd7F7Mzd+oyFTtw3pLvMeep0yAAWF8gskYFe2z7mvwlQxxisegw+TDZP8UTu9pOb+TaWTxKO6
aodDWCL3MRqCA/pxjl6EMaL3zmMOBtSXfnTdl5KBKHlOZecgwjxtXRKkpIFogfoeEKZ/83IKmO3F
26ci4FuG1lhZLBr5DAba3NDc3PZMciGdGK5GV2pL6W39anp/mmGLEzBQLlW9gGLlHneDCLONb5OU
8DJjHbFUto07HTOnqvbZjPEm/xx9ARanj92E+tvZGCM+AMVvFCkmDfCb8dh7C18hap+4vU/kG9C1
+IqwaBOMfITz73vIc2oVNr1Z9k7UC7D1OBAr7oz5lxYeI4LycZRjtC06MYaYXninAHL1Tbgd0gmn
FNtvMxOwr4RIOXVM5kJzmv0S3ju71xE8zq+VtUCGupzVpNJ4U+M7itDKGNPAT4Kp+4WpQVYSlzFp
NY9SQCI9Ly6UwbflaPkXm+3FFOxNGIPDsOASVmvaxiwdhrtVhaNdP3bCqm48MxCess+uGMZPtZmj
d3Ns+xvT0YCiTcwpTj9CiAjj4r0ntK2EjZRpiRS2+ILcMifTsD+/oaF8jtzTvaPzczDvkk8SqC1k
qUrt0T58o967PU5RIoyYBTkgyCT/3t0tmY5Ax1b9RsxmBA8TrHrUYrpicZkvZatl/HnAL+s2nv6j
Zq76Km+oofvWz+bVCW+IyMOqSvR5ggxncDXRL9r5C3ZYUwAIgibCD0cyiYOpWDom/wnAaLsbKRqu
e/TtTQpsLBKv2U2q7EUmxGFeabdnVNzzjwS9N2PmK8dL1x5nK9/W0wkWvQQi5bs8Ubb86rL4D1hw
QPxWe2imIUZgCNRoHviItxmiTLnEOi0rajocYZuFCdCgIctXxJPy3APf22u/5K/upbY3TQzDV7f7
mfeM0eN1APPkWcL/LpphBTV7bARm2F6W7DXE9ys8hcmV10oM7jSAoSH4oRZ3wgh2OhbjCoc5RZnF
jDdQHmq+PtmYV6FkQKF7g6CmYnC2agtpGZbiEHOyCKlIqR3DMdO36P6onU7kpVFJEEZs6jtRI7x7
uw/D5zNg/yNaj7AecTVRl8+ot+tMurQwlYl+KPU0sB+FbniBKNmXbT9A1PXbvz0uO89GfwOTcDC0
I3FbWbqKhY8LzqViJuUZCXsbbxQtHtWraD6YWjC+raKTMeCqc3MXiW6Uhu2kvl9con4xKJmsK9VR
NTZ8OXqrzcDYWlbTNb3wAMgHZdxrLCg6nSM8SEUIap+jpMWnNauYEbzE3KNmfi0GpT0KdZUhGDGc
Beanz/uDUCV8pAcrVtF+6vuOlmkTBGVO/BNfHpzMhTRD72o/Oh62DyaYoNIdoKbn/z5YV08rf2sp
6NsDQGPIc7NP3r3fQdqOuaDlD6UZWsum4QQbNH5r9rngXMmzRirPLwY/ZeUgXf5VfhiT1xpWJkeH
s5tz4GO4Z0EldHrmbkb24xMa3U1x9dUWZ3E6g4TFG5cUKNfbYVtIhhAcbvjQ8YciR9bd7rTJwxqn
JcrEv899w2S60OYd+rFBQ/8Zc4RWhPcAOVTAbEqyDJxIKuJivB1kDzi+mBTuDTfGVWutKyHnxfZx
WezDnXs2kEpSmmh6JC2BtiPdDroSt4Jo9tKH1NGkVtyD5Aa22yFxJZc2gL1UjP8PFHbt2Sw94pHa
0hIB+EAh6DzoZnmym/2sqXqDRwJJd2ubaHsdYKoHxIS7ygYA1S21cSu46dbsjIptYvUxORB11+0R
Exz6oPG9ERgaDwlPgX3bWJGNBCiM5FMergvn0qqRRh1UAuBwE8fYyaIUEHWC5bVrg2DKpewCBMKT
MfzHc2/xIpVkvGWiMR8Bv1W4kaFSTzYQ04z/CO8Cgc1BYTa7YozaK6ebF3EBJBEfqEJlOunujmi3
+i2jcQdPnaA9GeLRSq6PRugDlrU64qXoxUXOImQZPmToFtkRsk95Yz5lstUNaH72729YYOhFri2e
+15uju2BBmsXTTibHw6ROIFalwdnmJlCgvJ7scy+KTJNePDlu0MWH/tC6iK2xjBg7pAuGkjm77pM
tR7Uq29XO3wATA32xic3KJw0lDKtkXHSZZbaxnHz1kf2Be4QpBjHSQtT0/iDNm3mCRuo6GGwcSMy
5LwEqWk65amczG6ZODoDPtIe5oJkdTfptvzA7GV3BORzzNbw2VY88JxcsP9G6mWBKqXkT9yvIOAX
Clm+udDsy74ETtYVIs3aIxCoKkzMOXZLQ92ErzmvAi3lUEI5tqGUfYLXXYxNyIhboS2xyaNXvBar
G8Mj1J8nm9VZd7w28Gwa3mAVW00PkYDNOW3mBW3tDas6a3Z9I8JNF+jlh6bix9r9HdWjivq4Tmn2
C7vdNaYr+ST6tkQah1xhR1x7gPZGX/DzSJQCR4P2exD6HtP+vCpPsfRgWeIBhB72NMnENSXvNizL
rav3K55Cb5E8CdvuRluqwrfp6heTGyv1T0BLEZ06MTfzCPnU5jydmud0Mu1HDfysR1Zwc+gOw9Yc
RjTXBCp2SkcrezbgEGS/HXaVvbVu8Zqnlt4ylNIsR5LTg7N0fK6+deaI9DN+g1zLe5+rZBiwurRc
NrFEGn6030oDtdyUamJi5oJMkcVlzFmu9dwTFtxYpOdAd+5Fyfb7mztH6b+oiRCTeNSeWeqmXLv9
SwB5abZ8APK32AI2HXfWZOevDRmKYN+rm5FiHVeJ2Q7Puz6XoVtB/c64ZYLLzM1fRmirpvDjDj72
0zjmEzwVEEqQkMxEFuWOV3gSKlvdGJGJz2yIHI4HVJeKePiuZo14WLH3swF9JUlEK/HFdBDEnSmT
sodMPVnIaigM5ggpc7zgZrwO7ddvFUBLIqg8q1bRsUbGq+aMD/FsX0YjIkfmhmjd/xgS+Igvk4Q2
uPf/PUk+K9pj9x9rbXQdn/t4DqiN/3EKa4RIkzEtQiOgU0Rc8mBUFDQvcYhTf0nVavFN9BAry8sj
8posDTXpP4r12bgUjKeV+u1D8nYNuIrvIfhD0xIzkN3M1EdurF8L6w5bRQccJ4XB1ZX32L2LXfg+
RV70ex6wH03HLjetGVTqswPIbQmhugOpPX19Uo2HqzQqt8YUtkGN6Z3GRg3pXAIw7NqMsOQaGyAM
JEUYFrfB2U+CjpvDYfW7AxPaJbkW6CbEANcmIUz2lN3IS4tjNCdK0RhweXEtnSkl3kObRT4Kf9IV
GayWEPpx4XAQrXg9JjijKtjwAwnf5ZbvsJ2fDzKnoHZ7yxNcDT6VhQxes4LXNNXRYn5cWEh7UeN2
PzedkvDk2oJx76CJA2FpaGsEKli5UWE+p+OYbreqk8yULsodgIv3MMgKztiuWee4MmeNmP1D2u9V
U6XK1DTXTsGN8XouTeQ+Dvw94ckOGCy0MuAv8XBJrwyJ3SVVk3cLkmiwD773fI/ViQdAynwJDw+X
9l6LjrRY7DhKrT/9bCae2zqrExXDnRwN/vPe3wfjylD56g4BiSqAuQucygBjDo+ti+lxIcV7WlS1
/CKdUr8+jd/ZXnU6e3jlzS5f5P0dpHtHWM75n93SKblYboFpX6+bTRW9CdWL7Ykxpspo8AkZfzhu
jDGtuvCaYLXfbcZO8OVEnrQ7f3ZkluLV7SCSypNdebDkSec+c7RXdb070iUd8v7llEXLNSmiBUOm
EvXpy1EMpYWYWVEPJ0PM8nPxXqITqrYNTCgMyw4Kko/yJz938lnv2etK5VWeqSnEM932ewNslIuN
h2uCnUvGsqKWwkCGggfpF9YElbo/Hgvx0bR//Sp8X44PvLyS1pV2GRqLYESqpdsY67EKancaBmhd
INlFAZOq/9FA3xuFPskUGkVxdhpjjZiDl55ZpgzteaVqqP8ZC1mSy5ATgYJP54kPRPmHR1a0paCz
zw6auE4SZqQu8C/SrDAFgXtFBkRn2Us/k45U64iXVYpJpKcwjESVOB4yq5Eb2ZQr4v3J12+f0rRv
hX6tk07koXoIpsNdjL0bwjJSGG9GqL+AhVwzo4lP0XBaIERGyb9xPWiR1gvoSXuw1Zlw/0jmF8hn
k8pre2gW5jZpxCMHUpj1f/xsaG4zU2LnDdwA3VCxNAvxwG0iFg2ii8KLU7iVO/dSrV8LaUXlo1Pz
riHcK6wivGLQyQKUoGv+latysuAKtc0ypQrHDThtMUsGwIsE6ZaJnvjx0L/dFxF+MtHQQpFeuYpu
ChqRYfOao31zJRIJA43VeqBUqhH9pqZ1WDJCzObJHRq97qwUs3mgwagyxFgjScgKJOR61XVFM4wb
l5s3ec27oO2zTATeQbP8WQmO/gXL9wAdGIUiV4FBSR74uLtrxihWcZXmutv1NwosVf7+cLPS+YpT
yqiNYFNOe+sTdydcNQjWeEavqeHj/lo8ASUTAUvvXhCu75q+NaG3GC2j6e9IykyNFaw+wmc/OV20
zIKfCtsPj8QO/5t47fXIMIvt3G4HOUco/kMGb/TT9q70sXFl6wfDHDTjpXiyn+mJTkekT2XH1TEk
9/GwoTvyswENxoy4XdQPO7V55IVP4BY6/Sp8+PKe/eIRWrS1rersMNjFBj/8yl4uJdPLbKKRGdra
Hie+p5RGRphnHnOeGEbJIg863mXiShF1uI/Jp5HAfxr54+xCHeyXlJ4pkByES9XBozPPliwCw1Hq
NxTUwD0ipJmJ6BoBIlZZMoh1Jy+aMKtSfdvFdZaUDQ0W5cqdvddd32qNXuIdoRr4ea+HxW5ps6LA
Vat2qUyV9ojLr/oP6OR5geDZsZ/0uvbymThBIizAg6lil3RNMLHNMubCP/K+plMr2NUZe5hJR1wh
s1o6pVUSne0NPRJJ3t7tvreA3fsHGCemb75dSRVXcTeGnmhW9scJZBxvhnSjqbfY5Ilp7PQmyoGX
YuUqlF3IWKGdPN0kowUQq9fAIiMkAaf7+I7C9riff8Yy7lnI2z9w4L6xcmdnR2ldIGCsN0RnimI0
9AU3hTkvX8iU7JqFONVZgsQlMoibRl4YhAcwviqsSBeQtEDZoSjf7LpLlieGUiYya10gxwmjMgTy
ietkzEPQFoEMTP7VgNzyvPMYPlPEoP22/j2FPaSXusWE3LsuE3mdX1WZLpaGpbRIT9R3fl9qjReV
IQBD7wJn9zB4suSbj/1eXOocn693aSfldPZskqH2WA3hOTNSEmKjvyudGV7jyBx8ofVVNJkCC1nT
hKQDWi8wlAs8yZ3LiJ4R88BHhY3xOOe6y1rvFrAzdGQAvgUlIaa7DOmIH78CQcbC9tLY/RFIVctj
qwxmgh5jv8FCrMxIsndrad7AfeVNpfuqr5yMqIjUd48sC/JE5QxTAZFJeOKg2Wap8rUFGNot0b1m
V7McO5+4pGMtk3zqr+6TuJy1L2B0oSRUfQPYnkMU+r1oh3bPADhREgUKDyjUMQyI70xG7Zok1Wxq
pmUO3Dd5GJ2ukyne/SjPZfmPNUr0MNiQ/6PQQgd1KJHnphaLu66K9FHMnXXEDWUPgqqIFsSKbdvu
8cDLA95aOO5FM6Lnv/UbihYP4LimuYWSKNDAJ0mCQGmY92ey5s0QEfiWfm2fLcvRY9RPnqPW3Ywd
Or5uwTZtHkAeircVXM0DSYoSnJz1P47r0xzekL2z8z9zwwBCg2Ak13hdVurrQyjt7uytGne6PhFU
BoI6VP5STWxcwdesBFe9ASxnPHeItnoxo6gg+prAB5wdomermkSeb+apBT97i8FEshZCrc6I7NBA
XtcT5QnNwTYJee9ibey+19oZjc+U4eQFvLpEe9wY0fNa/ULMOm1NY5nkZ22aAvKyw95aIQZuqsar
b9GAI8hEvJJcLLFBuZV2zbzx7AqaLwGmTSOa5jzUWPL34c+kHseJOwx79US9CkChkYxfqIiUK7ev
2O8br0HeWMF3qLtJnm+aaH6k7KrdFPKTU8dYy5wjDUPeUBQ44C3MRxvhD5FY4nfWan+i4CJnWOlJ
Ea/ojB2Af1+MXszOMHEVp3uB+7RcP5hCTr8iwROJYXbC+GHHw9lxO3yfF+3i6yYI+EgkqVPgqZBM
vfv1oec3KPodoVZoPI0QBYdCVQyGhpVVQ4p4RC1GynS4itLdEu4aCfxQPDTd2awxJXuxM8eHhnhM
UvGSR2d8l9wlagBvT6LTujPfUD8AvCKEkGiIg9HthisMDrLxXwWCo4aPNFOmNBkg9aVTUsDw0jgG
zKzgcu/cl8HvgKUwDs/77/QBxLmdFBf00BO6pPiwNgzh0hPa5BTQ1sbgG6rCBRY4H+KzF3EZwNwC
BRx8HZYftjQGhoMMxVVQga2B2XT8Nj2V5sVAgfECWqohoWOAjHkjrM8qbdD4KW+R7D2DyICexbuM
9mlQBdeuc7oHDtq1AZno1KjXUXcK+SlIXDb9RztvTDenl8KTYMnQSZkNH48Vafa5+N/J69Fu2vAO
GG51g/BANwGDvg5j7lPa+i9iZRZxyeGEExxUFKmRE/n6DM3zGCS7FpcXS8Z982JQTqBwMB+6DIsH
MvEKi0c37Dlm21pA/jL+uuKlJeXDgLKqiFuc8tXY/CV3MDbZz2U9G5syHdfbtGpNYowPWI1cGPl8
rU83sXbi1s1e4TZyfFMxCp1CUC+EN0r7l1+5hzQUjvkR3FCTwKB+d3JFAdqAnpcg8WD74IknpwzX
6hdjBC598p8zgaTprUnivcc22+dmuZTLAtOUmGJguaUvQmpIvQuAnEG+dDzQTaaVU5jXnTRcAgf7
Ly6xgBJp1tUtNG/6MB0ZtY6a2CCukN7F40C+H4Sl/JfNKsMIDLGS8X9SkPWhxfiTyjUdqX0svdX7
lD1uAURQGqYYpWLsdqgp+dMKCFKuhKavP3B3aWaWRdskLwalIOOf78yk6IwVEchsJ/oTcValTZZ5
/QA3qIi+ec0Ja+r2fhJglAvtkDjPfsDKscXr6ssJSNz37NhrsnB7RjJJ/ZnzB5zHNtf5bqwNXfoj
kcIa7hcsLxXIJ4gAGjNQQAX42Qh7D58dAfo1KxLZyzux+aVAFNNgRERfxIEzJcVOa+Eltr2P0iYK
Gqws1zMUvkLketiZctS7DxhaEw2r5fhoVxjubLBXR3DG/Gb3mPgemxqnKMsRioeKjlD3XQJWKanh
m2gnfQPH0lX/ezksdTXsnXNugUJws+8oMsWGjIjg/CVDpdcgMFu7FRrrSH/kFzjVwd6d53RL1BCA
FBhqsI8z1KWXEewAyHh+J3xHJIKl1nNlHTF4ZtrUkT8DPzco8ikXVwtWCy/q05X+qPB/o/AMS18Q
1nyucKhKTAewxCZIiNGKqLnWaCsORwt0N4VScthez9vj/wri4MI6usnxw7zZlXAUtcWBT5J36Q6G
pzAQY9lyZl+awPJo3HYrt6ywNqTtzGGXqqNrA6bXreUt2R/s5ZBU/QkVLttKAJJoA2HfIw0+j2LS
x9KBXoqJZeeVB2QuquNhI5oxsvmr+8Br3wnQluWxDh0muBGW1tbBO404UauT/VAi341Vf9soC6pD
6sbIYtd7zTA0gbsr1x9MZhJcYtImdpg16Za3ByhxxkV6knVkez6Nsj23vo/po7Y6/wnW1KGh2tZl
s4RP3X8pmtdPhXZyUyKrgfiJvclWp2nCmYoQw+O7nDC04fPobetOiruFjxUXakVg32p9BQM3VkKs
Xr8tS+5UYW8LHBYsjhFANbtzh2Wnq5MjOjjobBWRTwuMnwnJi8AnbxTYahXanGW6foOUfSvyRVEf
EozJLdIyjJ9SfrYDWDCDBeb0+DTs4HkQ5wJGlStPHsg+crEOet8Xv3+TvjigFKO6KYebZCrL1eqR
0mOXuiJbH/N6Rr7TrYCFdPWJOWOAb8C1qvZ1F/xzAX0I6vQJJMbW2c+WHS46YRZ2dTZSuf5IKQOo
JoNnovjUWMcPhzpOEBPnxmx4bjpRGar+jUiSezn+K4JDNwi/SKkskoLKHU9g5Wl4U8kWhJFlA+i7
6YiyIL/Dj9bXoy5H9CqqLafvtEUoyt7aiNkQj5Frh6osmwFg5VEJofKTU00nPbjXS1EoI9rJuD1a
EsjWkUGCcP13sXmnGGIGI+uJ2ef3hl3aKiWJP6BxStqKUle4mn87PEpge+b44tbafuUxSNAbk0mr
/JpuQSzFNiMGdVPAnkr8eWyGg73y1fNhXFiFjPTgfZsJnS0AGq6Gt44ig4rrEOcceNdkLrL180zT
y5ltIapLK+2sPuem6yjqYOEVrExFA96q/pMWN4IIpA+6YvNsieGmtmDKTpQXMCEz8T+Va+TNlgmL
r9QG7qE7lCZoo07J5BO/OHM971px5UkfTpmsxWv0ze2k0df47JZmWv4iraZuM+8q3NZHEQzCGwgc
NE0dEkev5CBxUXlX5jQXH0G/cO00m+dkTPalWgfA9khqowy7zWP6rfq9tCLQxTN4BvsmfxGcmaMS
e4xSbW1z02cmo4+FIWrKTrO9a9G5I+qzrjGt17h7ynLVpb2U6PSClo/Op9IUAmhWXMdOBUAQAtjy
yuTuYz67yFky6lJ70GzIe7+zikcIkO46+C9nQkKajc/WRhineKQbxEBV8TJqLGwGuHBhkygOM+6p
pVWCb9KtuAdQNXWuiXwFbp/4FyVUwOpRVRH9LLT4cGooqvtrGsp/3loFU/rv/VGAQyivfPMrR3ar
uesxuM4mpAGn6c3NARnyfjXavncxFKUzFlXTDvpSWFkn0qX41rR2Tfr+OWqAaecjC1rIiHx1VKsA
eU2rn85j4J9P3KSMJf2Zn1WfWh+Sy/ppRZHnxDPQuGYGSPvNie1XpYqJZRJYYamV+bmL78wfqzZ5
ejbsQLW3mKixnfyzKsDPwOeN70VKvBMd50GVJmdQwOLPJFOLTdmUD2ydBzMECy5JSATPo3fgib9P
o1ixRXjbhBfQHUuhkJPukkOTwoasQ5KxSuut/EC74DXVrGwE1zCgtdmxgVcBVpKwOZnsIgsBDTv3
toXgd0d6Ee8vITyKqT2CB4+awfn0GGeMI49jG2oWdADOAG3KGDr8gzUCE0IgOu0gGWlML+Us6q40
/w2y1fEuVPBzUQLpsd0IUMtGQk8ClarRyQFwOXSM67OWlkA7Pkfzl+ogPmR1fQ7v5fWhjb/W+1J6
+JLq48Eiu3T7xyL1/eG8GxjZ7kB3322MuRNAuONeZciNXEE86XA3ZKIQyVa8wtPWiH2IwE88pAyS
+tSCdK9RaBhLwQTfuQ4W8whvFzNzygHsgBvLdzJauqCw7Eqd+v5gWu0p6AWzIk8mV86GJjlDX+qM
tfCGEkOLg6d5SKatPgo+aiAA0FxV8Vzj47OsawCXo4o3oNlXwuU3E1eOqM/FA3ZLXe9eEu7G9/iy
gB0wQrpUt3fVUo0tLyJosutcBI+tq0vAsUwunbugG6P3gKszry4Xg9LqdisZXXxmui5FOdhbnfWB
mOsyuOBaTuElkKWtdOFZhJnXKxkTejeOdaginkC8N88BoqrbJIV0LPZZxjhKL2ExQwnudNWEW8Di
33B7r78W25pp1lmvqxBs5ZaxinxBkJx5sLJgs82hfQ02Yez8gbBagK2V3wOzFZzgigSqi7lh6YL4
2uviFHZye56Xks9/lSxa/DR6SndiBTv+Oz39S+OGHaGbheQ/xD5JUdemWBNzywqySK+d+e8deg2Z
wTvZ3putD1O3AJoYeCQPFVnH0ISk8teOvkUkUOKCdb3xZh+DXQHBoV1sGy+uwv5qQusyA+ZKZaEs
0EqzzL9ksptRz97RoavGFEGCj8gyi5t3z1trqRKHKjr3OZ2CS+RTaPMdwso217Aza7OT8zHlKb80
ERTvSMhatbMNA1ohYQ3t0crxVU/za+fxoF5wp43tmJ2OM0QH2Y/04bwfXnTjAC7rVfOVCCbV35js
6E/Um15awzo/6bQpA+ojQ2F+w7M3nrQ1y3bipYkCWHVUSGl3tyycdiKoDDIX1xEvGR6rF22BKL7j
xZRtBxNu2A5XhxCmnk4J+UgKvaKJ9d+GL3OCGS8qx92gTBIiw2KFdWqv1d6K4jEKZeh6GrAFm4Ym
agRCZTJToi2GqIlnj4DQZNl7i3MBHq/gQ3KoDnA62UIxQICIf0CvurN6ds6kPnH23Q0rdKGiyha3
LuIekFuf/yXVK8DzUkj45vL3yo/pI56bD2W25oxQRQSsmFFY5iKitDOpqdKWTo2A0qzySixzeibp
e0bKATuDPPtKGmqUd0gfdkCQA6DRAINy9a1fGo4eJ6K4X9OfaQD1JY18SXGltrFIiXwuz2GffBAK
UR0RAsqVjGdmEynL4DYGV7CM3fyQicNLGIxZM4fV3ZDQUCjdktd4slHW+Nd48DI7qZsekppRGlox
v/S2zxNDupUZZFYeMUTOv7f2g2NYTcI+hI6vtIgNBvPFaIAOMc944ysbf87q0gkLuVK8SF/XeP6B
JQLdwptsIQN0zIcGwmGKvN9e9o9YJ4cap9N96ckX3CvV+uXYnSAvUKFGYyoRcjGeRYTW8x/USifh
x99DP9r6CpYuACS8Bs+prRc9UnriAHQBJbeyB0j/xCJIj3e6lAo2xaeuY1rmLIvA6jb1qKe282+/
NAHAXEK94yY/7Ks1oWMO1jFTPbrN7XGaD6FHig0iXq4ZtVVUcZYuPTkG30vv1btLAUaZseTv5LiA
AWKRHwo5tiw2i8k/CGwq7A5Oftb3kCSbw/lJ/HW6aRygbRTwGQcmXCkQgq2kKeVo1rzQSRMLgvhs
kECygVsutGgLxxTjodyFm99ETOkT54+inl0sB3FOgRil9seIydy/lDHmW1o4KcbP4/kc73FlqPrW
edixdpMUc7Zww+9puGmIq4+ZXe7npt2DpZaM4g3m8iw+5sjdR2YswuHqQ+GR7JYFnB3zm/iGqavN
RIrFJEW7Dqa+X4lIOtuRSv6Y8XV/fPcPX2KR4H4NiZonLgEr+b0oeY2qaPCl4n+kPnJf3td96Yx3
6kJJ7YTAlASImetoLSokoqkzjhl6xE8jsYj+vKmMfYQ9DE1KHcBVOoAFkgcv6JRl4ldUyytdw3RI
yEHH8b+EG/y0sx7lQIFJpBQjD0fHK0oM9mlXYQMpo7IzxH8hceGsw73G3OaReKCZ4WpZBDN1/Yrd
iWnNQMI2fq3ZYadwNJ2HGiTWRcmmvtlg9Q31UqrmrPFnPJOpPIbJ+eWBMsH5gUMJriHX42hIDOQM
823C40WuU7K8XT6wSAGWaK7PfPbyF0R0ksYRpy5BegHL0R413qBHmk+UQ1aacXxbFHvgPyaLe7g1
TebaMiVPSTZnorDKj486njiDGkwDtnfEzm++zF1fcEarH/jnZB2uB7vMf4FMHzXC4pX5J93azQGK
pLoO6UoTc/aa2K7P7pjxPT59BSZprV0LoPqPdO6VKuZSl52R5IUPVW7WX/1RMNsRyhafihC4AAtk
tQ+eP3Lxy84b3/xPFLf2zrTTGRryCz4k5CQVUNiu7C2BJcN8bUsVDUIDelmRPA0DVezfjIRedc/6
wjYCXBS3ucdwnnF8DzwV7pBNfacFI0NyMtaMWMU/d1GZCRNrA91mjWRiPnNOIxyk/7WExPMk2cHK
miWdcbKJGpkjD09NowwpxhNRdcGxiuPPDQHmMVPXJzKfJ5/lXtF1A3hEd4XufXdLUd/rAPLw9RWs
J/3eM160WBeugOGhECfDNcZpeF55wICSajjKVJCtYTswtIfYDWOKy4J19oK+j3yxexiaqEh8Adql
KkZ3VoMAYlDQgpd0AewtQYHuCUPXp/BP5mckFcTgrDF1KJMDIGCAZi9YsnII048FxOGsrNSfMBzB
slvh5FwBNvcm4JiAdn+MocTvLUDgp77O97LKfaWPXY+CmrxaIvm6lfa+PR+NdXNGcDlCEiIuWUHM
bddjGLzXrfrkPjp7b5P+Ko+oZM0yC1ZGAfz027gr0XdZsQbWoCBzep9IZk3GfJhMDF2nHg+Aqny1
aiI0g7UVu0joGZeP5/V84shdBBb6FqrCd8KtX3RTcIYubaM8uB5VZAk0hq7GjDYDcHrXP77eJrFQ
B85oWpeeNnvpL7QX8P7ckxs2cjmslaiJnHhnUgS4CdaSjptSrl5mIfSx97h6TojcjX5RAWuA/UwZ
0pxwwmj5CyAFU6LTSriwSk2tj4q6ZFkVxi+tGTRo/kDXmyimFR2wnkqsd1L8bZsH4PfZeSr7IcET
bqDwEgg8rySA4FFLQATb0zHohmyl2GGbMlK+h7PgDimYgH2pTdVu/6tKVOAKp4qhbKL0MUNKcEYi
lLLRDDFjw/FhC99+GHvuTqhWs67czjseHTAVj/odPByBJS81Al0CzsIFN49rLZ2a7f7YgsZMQwGi
32EZ8wP0TlS8GzfiEZWn+pytS6Zu+ANbtrjrARzB7/vm3SBWjS38u5YEcFtZV9WyjLFcE4ZIeVyd
8stkXkGIzvogwiCBUdPEzApppPkU4AwenZluooeNxTniEySEq1TJA1+1V8jxxoIxGATObx7AnGza
MQ0P7zo3NQgENzq+uNDOY8P2bYZi5RfKMw7oPDS7ZW39L5ZDokikJYcmTYQSa/N0tPi3RCsWP7f+
guQPBABnn/A3/D+aeIzCObRrWdrOEfsp5vEzSn58QL/TxfklNGbJMnoOf9eGpv8fnq7RGsVpgvLR
zGYcUv3U0XFPC7c55Q+yArGUprZyf9f9oEKxacJJpZ+APXCem9c7eJFnhO2PPOROtH0m9tTxhziN
TWnPY/tUjVM0auJrQTF1zgNyhGcuxCeJ7R9BzFqAJLxbM7GaE/NRgMjsvuFcXams9CsdWovaMeth
slwUQBehh2KA6YqiHa7x611QVKyhJo2xcBfn+ZZDTJAJyr84qhymRZv8vfn4FESwc8mt5Zji9R9k
HLNwNPUXXOgd1OElR4Z5XwUSr4GQ1G498TrG1HflAkqhG5RQUfuGBiaEY6XRu5AcOAS2uGCqfC1F
OmFjd9htwwX5bj4rIHN446OXhG1n9NT84AziBW3AlmPmar15hwfWWgXzyNFZk8xCEgssO3iaAcfu
CfnAsYftu3JZksakv0SDpytC85jjiLs00Ig99mGIRuGoO7vPlvzQS2RsJK4W10cZHXytb6vr7mdY
MfhXgkO5OD2wdqXiqqOppfzHxnjeB4ULhiTrWaGwyDVkkAPr5LG2DniHFWsVJ4bXIvMQuP6WSAVD
gAsofg7LczbeGNO0fdYTuV44XhFzn1Cid+xIbcJLWfMAXCA/iUHCcKtcJHNly6WYW1uf8bIZ613P
nby8J419rW2TYRtjnhB6XuEYem+wgkbyV64H05SgNqDyw1qdqZMVe91mwRnlj/R5swI7fygoK3yC
aghmGW7rWPu8OhrlkDDwF89fiM/7V3QYdwNKX6fiKEA2yHDpM2rtleIFoJQZQ2bEa5a5YqIpIJ8N
UyeM3hGO3j7N/CLjInaiMICCMSTpYnYL/iDsQJajs02jMa+KFyUXWXSXXsRRkw4IyD9NfWnMIktx
wpPMti3v15BTPC4ZAArIgBh6J0qyNtT5KMiiZqqlUcrIMOTEuOndh/SjACKG/uriEehFVm0uVDkG
s8o1+5ugaoN1X5suteXG4Gb2Ggihis4s0u9aFGUA2sG7hXMneQHz1yRw3kqM7f7dl40iXEoCiCIN
k8lrXtNDUHPfm8BRZr3pum2FvdLeVDXcGr5KfOwbzAheC6dQ0EihhLiaGreOdDnBYaENk3F6t4Ia
G/VduYwCvV0Fcif3TGINIjizWjLueilf96MiUUerGNUBPy6BEkZFNz0rRsuqTJQkArAyLXxlmuTd
txvYYLzhgK6oRVFk3bajpxfxcJwhcgVO7NyTEx7AK/IWskwY7tek+l0rVP4spoTLBsMNzJ9upHII
Axf7sxOXAAGeoZ34HMKV9DQY8FHvFtVJ2a5TonQz/NaN6awmNRAIdcR9m+tFlR4fzABl8JelfBOE
L2f/ZZ6ZDNwMfyY37Kmst+jCiFtjVLNOyMfR6+WyAG9fqo3fmjTdugaZ1HMK3sXnbmOBbwlr6f+S
0QPhVvM52DvbpjuSAJu+b27igCZXDiPOfzac56E0qamDaw2+4B88udS1M+kyX0+ep6ngd2IhEojw
Cl1P025gWfgkyBSELVIGSU1Dw71mvYxzyjd/eUa0hbzbXtDoQr2dtgmcHXa0ifA7YnPayGxJXXiD
I2tYnChqKwvJcASDftrprdin+SiIBZ/S2I7f7xH1ncL+V/kbgOEmlFtGIvKYTDg4pYn3niRYG4Jg
ZKxxiHhrCyino6YlT/AzotpJq5FhKJzezJttJBmNl+Ttlrt5RnS4tMK1BpukeSJ7Ofs2psummKSQ
t43g78Ta2CKOJIOT3ntHSNrgu5CjpSmXYk9h1GODy1RDuAPIpao8cMQMPsSvDSlwXneUoD9GXY+z
PqipZhn67DJNFoL4+wmDzcRGzKQY8Dr/UjilEjRxivBjHqbZ1jjxW7ItDmUQJe5gFDDex0yevvqS
u4//Fbfj/jEdm+x3DGHGsz5hf/ODITUUJnHM21p7IPjpcP+rqfxxKkL7VsU+1njE8Qj3tKYsea6r
kBRdSdBiHFU3zEiSHxCXoULnLuIDkr3RJFsg0YVLmTk1EqDikSMMmGw11+IGRAyQ+SUGhOrYyTe/
PO9HPJONxDabNqmO1bvx8OnVZce1qyC72EKfDC6F+xr+1tzEJ9/dPr0+SIS96w5z6S7wkW8bneIX
egsvs7QnuYG4ZOxhUcaOCWFg0JDVUG0ShdiHX1Z4J6zA457ChijuK0qE05oY0rUJi6dBHKl0fnRr
HoeT/6r9oDBOqLy14B9m0lTW29EGjQHNpVKqAUPjT5O+yG+yzLQSE32Yl0K1z9QjBNUndTbv5RBI
0GRb3hDirlZhpEiW53bedLViCQqISf0J7oO60DqskK6gbJp8dv27XIg923EebBxq9Nwn2+WSsg4k
TsTHSCuo/zFmD0bsWGVajcMHJ0tZdkJ6s9Q97ipxu+m+GuKGBeuCvhsTwK9RXF2Sy+hOSg3jTybt
9NVgdRmrrNQTUp5qOa8tS4FSAFfwDIUwSbkrUmja0jssHUBLzrwlteoHFZEARl6VnvWSjOuWvxqK
z5Kinr45ge5tu6mN1LtgsdnGYY25LD6MQ5fhk4fAk2hy6agfz1LRKnf0AY8g7sLcm6Nwm4FaK9CE
pUOQs0wHPmWHDN4//3cshOPKoX9d2whmpFXwDDLbiVGyPiyPaUBTILtzXHx8u0h6JXuF49ID+k2l
TNOrNUebL9es0X+qXU78fycRcNmTHHVjqB3HWVzpXQKtPGwXNkQRBpFIp7RosoIt4RWD64OhVsnm
WFKArwWl01aZ+6N/xqjlLwbA+CN1KwNktsteDuhMZ8AzoyXmLHQyUXCzUFj4cLoIXL2Gy+gV8Qop
oseLtk8UPNpZYYq+waO4DUhefGGnJEAlStXrinDe/LnNbFTmDn9pciBl5Z05SjfArdcmAhbzTEbD
RpBAmAjorBnX5e1m2Q79tXWiX52WZxnvYNyDazWL0exbppZkEixFKJbb726tT5mt8W1mjg2fcasI
mRy+mz3rx86+3YpsgQdV2XYS4hFyZ4c/xPzq/EVx/DC6GA2hUE7n0yEmHZcTtnYSCKSh7LcIia+j
xGHhG4kwcflY8yBz++3+5AqvnN2+cpL2tybnQtGYhRJkr9LF5CUYc6JAHW4wxan57SgagNxOr5gV
Crq++syR4HannDVZ7pDs3g5OaoH9teATPjYyWJxdX338RAGZBER6u3hxDEyyyGitVlohLakdo3ws
R9UfFjpEf+XkAz+KNsKRcHPen9VnQgjSK+EMALgX7ix+D16Lwqza5OxEzuNgFAPyWCdRhSZUfX4t
1CAtzw34dBENxh743R3CPBRcoC2tFjAWwh5n3Z5en8j3wd9FzcjdV6TqTDIN26w2M4sZRjXjJxOK
MCVkr+DpZV1l+ebNdUtyTxIGDFQdsnWvCYKAJkT6OhOGKwm9Yk825WInJr9ykBqqC7AybyRgnfT6
SltoBPfcP3v/FFiH00eygPb37DLK3MRzQXwlMrKHxihYL9pP2IK55Iyr7BRqk3KA3Jygc0DznME9
/AoJ6JtknMvOzzCxNZUgpbGhkNjtWbQO4WE5KB8YwAjnoCO0xHXP9s0RirE5rUYF5dTBNMqqw+ZO
lZLoHCQ1RvxJ4c1iop9rIo5gDnaFeHi1bdTdmLgb3ZUCJ4cG6LjfTUGQaB9QoOoB7wtvS3qYevok
yordRYAVgVV5cP0uPVyPa8geNc5rUSGwJKasxVfNXfHeri1h8I12r2HXrZiHdT9aAZaTKquenVoy
T67TVgMZz7gJFpdmvHZn83EhDGlKCiM6xypejyTi84qCQ8+q1Dq3AtL5KGlrJzxHwBDkrZfRfnZE
XKdywplIxWoDbeA0CcD6zWTpixJ9+N6r/0DwzuZ5bxZVjgiHDAQcSg9XeTwezuYcC99vnhghpHYr
5k9huJQOJUMZh4/QZG7Q22nQCNumncET1D7y5tmKy/ZENmN5QI3j8IAYbv8pR+KxJ+6SHHNosbTt
xKiVc3XV/5ljucj5ju0DLmDrp6MdjQWkq3EBKI3o41YfDuT58wzdGjhlK22hJwzyTFDPBMhbuVcu
wXaR0mbK/SWEkGdAGjP5u3wVv8q9u1xqlL5ymNnv4zzFisZWO0bXYu0wdDkiCkbLhbt7cJFLZQuj
JAIEMKOzk+hFY9axWkYs4oPXM3TJbxXzS1zxR2AdLD/dwdf8mgPqBmKsNwwQFSkRdL/66LVPbPhs
+stf89ito1CqLoRszHOt8eTf7GYhbmvBDNvCZa/7Ax+gMyoWjcNdZPJ0I7WwzepuUJzlvhR8RnYJ
zjQYuRtbrzjsVwwjtgdrS5l+0K5syFfRdG91XoZSdMfl4V1zsqZfS0hPm5KoEoy4flPLHEjkT2c0
7dLU1JweiwxZAWaqROzMonNqFlK1lZ6samUTHm364wBvjY+VE48jeQANmDC2OYt6DDsyXVrQEmAf
vFLTgVa9yRyahnv9vSt1mlXtny4aXf1p36ipFzDGxmzyYFcR1pjN/zUmH7AL3YxD8vWZTj/ht7ra
6NRkyjB3tZBFKI7cdvpR0VUq/obXNMVBd4tB6FZiQKBhXtDH9l7Xah5WKLmp2y19na35Y02wB6RX
GYo09aTYimz3Wy4MyTUbfnCOAy3S5melejf+AUxT9P7+CXjhy2kefJMLaa2g8sdcg3s3T3ldbAcM
T4KF8q0fWnA45xfVpGJo0uXcjQVBpcFzOOsn2v82YYKCm3PzifLvWfmrMQg9Tp47boVkVZ+0BM2G
jA1CDbV8TkYEaCWKf/y0raZatGRkwI6ssVc64ug13W2/z5al5jd0gH0E3R82KfnmAqdUKn5bJs1e
GT+baL+U2jFJK+vS8Vs26MiNxlBL+4RdcwOSkOAepuzYcNPAuwNQTuAU8705+t1CRGPLqrKayAdp
SteHSqK/0piUN2MOZy5v6lt9jFp+vsG6ZellubyaKXJSxGd6AY4kHJ+yFTTCo5lfYmo/iWlypgXv
NUD8lYdTVX0O/ZZFzpAGP1xE6R8fjtF/9JhZ/apEUXxdew0Vlh1xgdwYiBtsK+F+N21TRVY3WcpO
kGwzcbUK6CQJh75OH5J4taxkMLoL8VwOB7bmS1JSXcSV8SzdUg+CuocuIqyssz2Ccs7VWkBvfsMY
uniYo4SNpSIK7fjYEvmLXalQcF60u4S/2nEo+1Z3DjxYZ2rOypD22+5pfEinDWjTRZ1kXdDGon7u
Rfhnu10eY+oSl0fDEqzcM9Lp8k08jfSMVS0b2SaHFToMFc+OQ8G/QOJq6g5P135c2CW+51rNf/Jp
DmTr7sY/lYeNKHp149JdmuJCZKq/BAl2oIHWj8MUm01ZQUzFf0w0Ghnj7AYFct9X4xZH3/LfTpyz
fsY72vPielk4vzEQ7woEZw6ku5KXEqQhboAvwNAft9+LirYTjxsPjZeH8HBDSDA3oKiyldhTZj8Q
eBzUkCy5ujVC73yH+qt4fKABrRlNzFT40Yc5Vc0DdowFAxGwhqpskEMd5siJ7Qu/POqIgIi5/03X
YJ5ShAQ9DXAoO1MxkmoblzbIMud4gbhWN3YMnV7TRkTxwaepIk6gvVRB7043dc2EeTkpxJTqyrZI
cn8rke8yB7EwrGC2fix0rYJNpY2H/lxc00t2f7EIPK4VHwo45N8Z6A03o2MAVJeG4Eu0E/m5fsCg
oMLtRGNnfcVlujCk6AKUJo3dNxIzY/wojlr41HH021N0NAUTwkH0es1umM97KNn2CXmDnzKe6ppw
TMSiHEfCUs7A0Rb/4HxQ0AczkaP7ck6+epvPAsZwq+ShZ/S3WCupEP671IrHKdSM5OX3Z3PQyU0d
CQJ5omYa/hBK01R732uZP34v3XntXTHjWdZwYSdFJRm8Bvheq87o6hLuu8UElH/7l4WMzmIzv/yt
fc7bCxospfRFczQew1T6xwJorFQCbvfS6joqsyyvPVhq9RQEnYsFasBewoLn+wwovw7S+NE55Wgt
M1zm7G/sUjvWtzG30dFA6i26wKGXIPTzuQlFYASOoO+1OvjNevSYW0BtcqoHNUyEfp/+/lB9bdyp
qTLT5uM8XTfH/iZ5Nz3WqVCup4Ss58nB2JASlyDk+kSNxNvJK1t6PWDicH2VH3GWeomnD53V+ndk
04FmyWw7QmcF8mU6qz9oBeftcLcMaHGnbuhGni2dSW+UfRvb7rkAon+JMkFGb0ILIfRCvhpL/hnx
0FAsbwQaPF3HuHRfFNUvjwZpx/QuR7W/NOqpepUd7q0AXCZczk2zfeP30dYfx6m+JqLIOCXqmk9D
9CTN/Ic84/N9b1N6zvVnNYkSUXaVbYcTAHD0b+yj25otKUN5dla0uX0lm/Upf0YyQuduRaz+ThBz
I2XXesGkhv/klI4+S7lJ7N25MTnBiRwqTVsH25XIjJiKO2gxQ9Qc1d5urpYo18SaKW7w07Qyi23e
+F/V8de00Qa2urc+bg53kdm2n0qmmw2J37eaq7QtxKbHiEI2Z+Vqy9WhoEJwSs63PBWaDwcxAyF2
eAvfxeNZR1MCBDzxA9nI92sR7Get3OZTSyv2eSHw2+sBnZRYAPcren/G2A4msYq/ESrhOp1lf+n/
NsHnoB0Bxjr6SX8XiD77AWLk7laPZwtWRAtnahyIt4v4UoR1pzzsZxo6Vb2poilqRJJGPkJTY9pL
8XpBFBjhW9IbxI1CVQyrLyEptdToPlsT6evG7xHAm/vlQ/JrQudRkxUgDPqOORzGaY5Mj/abDmwk
tkJPLKMRpHBjlC47IWJtcFpdKQIKMh+Zi4UjItTOahy5CxCBMA4OqEa8O/HenRethuaqn/YCD5KW
6/svuvm1iZUzFSSkg9Rd9fLIbZ4MDtIDY0MIGOduljC0UX9cEl7EIFBUVChkwwUqk0HI8yglXfTD
BC8RnrR0tbE2NtG6pZSaNoizIKIarOyWzMC8S8MZn+elgWw/3j1Uxd5WYo2M6l5B1fnKoEANOz2C
6xpmexMnFE0NS2RpLUZhOg0sjZVw2Zim/Jbdy/i+KCcknOTCv8nRmJc+USVgaEhtkgpaXAFpxuqc
LpBMJFc4lUq7oFMx+V1GMLaZORlCnDfVcT0SYSWTy5U6M6C24bRGVrc53NO+nbsehENTR8AHb+zw
4LDmw62i27oXVOg0+/fkpVNs/Cj2oEjilSfKPniBsFcVsKVHG2HNBVwPPzQeSsVZn3PDD12Jsg4V
3kkh4AyNgJseEoOvYpo5BtS4HO2Ux+pRVb04v5qX8ZiPQJifnLYewdv3ZkvRcoCs5Q87TOY5hSGa
Vz4zeC6IlLLgUPcT1Jy/spH82KJls6anjcUbvvH5miMwwMYkT/4d8MGSgBBoHeQBQbopqA9elN52
u+4mjU0jrYaMzHFbpGLdOjPtTabXvWlhj/bQpsn+Ib2M7H5hiEZxGiEmlceI/MUQBNT4MPPYWtco
yZCZNpRzBV1+42lXarb3KQBR2fjbBaj1jEzSOtVwpP2TgJvcXCDHH/KzxRKy7wFXQ6qpwQj0mprq
sQy5s+mGMQF6av8jCDUkYBalIXQicFALajyE0IdjZTXcRWl0L9C7wlBAwcJyq0vzRXK2JKzYvmLz
t2YwIHFm1jRfwSRBThq7nRIhS+8YCj4UUe21s/3M3fPWoeuh4Z046DBEpS8JvmCljd71uSZe5A7w
Ue4p61q5L0u/ADTb27Kq5tx5RMM1Y6CuCKVikXVZCOjqRaDOfDyVH/h/5+9JsyESCksZlvxzvhWu
HCjw4BzePgTVaHymMcHbjHTkC91aAQegH/yLzO2Xf1KbfOKaOC4rrraL+FEjLVpmlcA+avmsDatC
q2hAe+XZqu1BG1zkD2MvvJEGvrXtoXhN1xr6UDB3PoZTnk+nbY8+dAVdqztngRJ757Hw0L+aUgBy
56nGHxW+32ZZFP0u1g6Wam/5kfcKArGA2VMzhGEqv8LvGLPuxxzS1goxOxhNGw/g06VktNpPKTUn
h5zB2SBjz3jgs8EwLLg1udjSCaitv4VQ4MDxm9+k/Pf2XxvrcGmVtVkjnfuIQc/sKpTf/AFK+9ve
43En4NHkGKTnpOwuuDwg/yq1yUmYRGPtR7yCaoRKQ5LgZDG1tPmmKy78s/ONreOS8sxj4wzgv6L0
Kc5YTboqcXJojhVSlaiBTNns0rB2PlqjiNiJeby4uqpax2yxAy0Fn59sEJ0D1F3PdBKW5A6Xf2Kf
TD4tGIdnsKAnyGOJkw4jtxevUeD8vleI9YJ82ZNLmxQfqxfylsNvvii4ha9x9YpofjG4aepP1/vm
kibIAIBH5B3+s/YuwZRdWTawK/ngBxmXF8wONcpm+3lNjd2Tgqn4syCARew/q0zx5A7Y6qQ8PSkK
UIZl4Z/22Jx9BB6YYMevYoQJVCJqz198sDa00mykZk4sOCoQW42p5xOJa9sbYPN57u70uBFE7L9G
9iM7I/BaH1hTUdmJMIQONdPmAD+xuJRsWh67eX5aygkTqBPSTvwAS0+bPNlDqHmGjN3b1BzZ6yx9
ZdiIRXdP+kJtETshYQ4GXBpg/3bjsAxjmG/n4virGqeCAGrvssZgAt205BrHBA1eFWlEclTV5ahc
IMVrBjO9H/ZG1pIRDJWFd36BZaWqkxiCE+tvU8jDyCJJHm1xPYVh1P0r+FB5lMi7FBKeE30cIY+x
6NYm1byeLRLN79/2nAlBEWSdwcQuiYuD3bAbQv7RbOTQUZbDeGkHfJvjDFtJeIjPe+jGtZj/AFvi
tn5s9IoGl2/32PeDs3recIx/5ldUP8wjoXtLvQGOMOVzIePp4bs4LdsilC01WDW+Ypjn0TTtC99W
N/YnFKfrl7z/7OfdRW/zJAzJnfA+XpzN54uYlRIa1q+Rs43soek6WiLSOivrApVy3Tq5m5Jkr3mL
mT66ByqxqZWEML/R34kzoRwgYgYA5LzMlfiu4noI+zhEVcrINcWU9Iqyzw1kQsX94OQ5D4T7gt3H
uiJfEjLUrPqeb4KQwvrUE2JIvrNlDpPnKbb+fGHzFnYeNfs1lXPFA54WwWJiomzzMAiVxwNPj04R
z0b1/a9/3Y/JjG/TatGDSxRkE0XyEo9yaMLVOCrvs3WPqJZvWbnfi2/Mf26H5s+H950yKRMSgfBw
u2DgMJ/LILGLBThDXl1GtkyhhkvMAc1Q1T3DzBpgv7d/xnGL6t1T3UGlTEHWe/e3oT1ACdaW9v8o
b/qj0FKHypxh1ulr2ygColiirAvoX/C7D5wL6enodrlp3qhs60Hhtc1s8jxe50QSapF+1K8qe8XL
MTpAh/GKSqT6jhAy66lEExQNfHcvs7DfQ/QNNozA4YeKVMfL9ghZgqTB2RVPbmcT3aUtons8txcI
x3U98+SHkfNd1iKDdK7rmmenpaPnSM5kPWcFx0Ylo2SQLgkpaT9ZpU1RJhgGIndys+DccHixrA7B
AEezYOVSwOPt6u+EzX1sO+Hy/RxUf0V7u0yvk7LQbRqhQLEN1IGXZjHy6MMAjF1cHGmX2qYAuU9t
3TzPRHFjeBiwDhVNezSQAiShfVMfojvaZPoTlib+Y7cVfmOMaPsNPR70ihX0MIwYF7zWkPZyNj5F
g9UmMwF7b72xNa5gDd9TaktsLJTdajZ1XFTochyPSrQS6yEXR7oMWgT8GO+lgh1YRA53Rz2PDJ6V
85NXhc0BO1NoMxGOaNSajPTLD6b09nQ7tNZv4Ox2oJMX3fiHwPwakZbNwqXbppMFF4HPpuGHILVn
qq9yiBjy8FVsk7dJ2YCHMh5d71hO1dbAEgjSvSyBOUziK4EM2O6B2Z/CeMBXoUXxyAM+yvfKjYre
xZEQklahhV8NglBo3TDs/ftdZ0rQBZKnrC/xotTorbd1tSLVsjW1kiIQjCt3TUPjyY40t3pAVd7v
55IKDFon4ZuZl9NTPDLC4RYAf6/Arf8+w1sqItomGSopoNoafzM/FZIlsB1ZbM+G+FlsMIKa+r2Y
0L+WqT7a3JkDJmMcF5m7Wz6Keqs54j0rJhQ+pcwRUJBMbZND6BEXhk4hlr2tYGWojCiFDq83Q1IA
4DkQpK2k2SnioF37auO/fJ2Q3P9PBAZNFEq5h+T5yjd1CTUZcOmzoj4jPAtsqx2QSbsHSdDDY7Bc
+bv72gXsgilJ3NkWWXT6fKWJhx4DyCxQzrdVRQlpJbjLSSIn+vistwTDeb5KNZuU2wpSeBlXW46m
n1/6hMkqFu/dYqL1Udq2AZGa7IEdVXh7vOVChdSpzkjHrCE7W5Bne72ZnJbr+LSfLWxdbFWlfZaq
temqsA03bZpqZ7q61Q5q89sXMZkfqQ63iYKsB6n/uTyFRMQCI1RvdpdJCGvhzxTTsXcvAvWJjNnr
UHkXJV3CdVVxVSH5d5ETlGuxJHd2KF/PxS8lPAk26c7/QD2zaGmozDU62TazyQff5yihCAgB5Jlc
U6gzCnw8Xvd8vSXSdrdYk+kuq+e3Gyxea0b1U9WUDHGGNzaG5nAeOpggKw8Jyik6FbvEEXkfe67i
VEBtlnLklbK6Oz1R0+lUuokhpP92wo/wOklROR+TXqJggnyukx/8O7GSkZj7Nyacrj8CTKGyOGIG
Jc9IJfPrgukBMV3z6EJ5NCO13mhNmKKGubmomwQEUlHd4XZtZSAC/sOQZzaFkJIuTM8vvu87GCSR
rpvoZn8QnQ+dIRdhDlNss0M250JF4j321lZ8XnbYXMFzn3Y3/X/Drn46SK2aSARuWUnR3E/QnTaD
BBVKTU418UPNXR6cNj19icsiabczhL3uMKrqlUGW5qyz/hDkEbtNZuYEcoWWF1LXM4PJUdX8nzao
O9+BvpSB0eKRAX+zBcW1zL1ijjSBHp27jXpyrvRD6nrpmkwIGaYxAt8xjPLnrBgXt05CHLLi44O8
yHNjuHrbJGq690Xvxur19LO5+UqB+xDM0FaUF9b2MZBncGu58fDDxxwyjB00Y9rQZBuIJsIyCAMl
E4KoVWbSO34UmM1Hc3/ShWfJ+tOeUEFIwdI9pgfAqSuQw4tIUrOYYpj6VhAtT2531XBhYPpTi5ja
9BH9mSdwJdNWADx5M+kKwnn0RuBhSmxnk/RSAfFT5kGGDZvtNvl7buyR5lJY3TsklapUm5Evl1fs
HDCdLVnqOXt0cseUj5GNQOqNm6P2gBq04I9Gids0IA0YhWtMurFbhFU7uEOotV9KbDmeooch4leW
1F1gNe06X0HsirDil6CDMtt4UOJT3Tcfxaei1q3tgD/zFXtToAxS7LI+Ddu2rNTn79+gpdGlXczP
LenooRz8Zw1LwfeGQ/ZUO2GLM+pmP1BDA8MAZF9LeNYVZLLN1RbzHm54Zrmxas9L0Z+YZRkWHO81
TExri7ldnlWiHRJO8r9bvte0tItZkmWne3yXwtSWd1uUhROCAhCvLJ77fro5y7buFaPfY6r9Lwuq
m6n/KaIZsDbPXt9L49kG5hvct9xov+jwCKMpHM+WEFrEc7PbJZezJCB5UAg3DRxdBWBzt/k1smwz
Qd5EEPV3KUpktXvIY/VlqARFcW1wuPo4PxrkJFvnTyaNUvu/ZnT825Eczsmtzh6Tt3I+7Tlvhip7
/meiebPys4c1MxtbyQshNIyWKwNROZSjhcYqkQoWjlHdm0MfKimI+6hbGAsY8IrtQoDdtqNrI9Ub
CF98mnkd6dSywe4oO8+jKMJSSLSLzZW0taSWsosaQAcA4QQfXk4I5Ht0fWmBnwlczQKJEP9Z0Zba
JFg2m1yjhaMRm1Du8hR5K605PlSMcJiTgZG5DoVS9CKJe9180r+/yh6PBXV15GSn9d8SmXA/nfUF
u0L/mV5S+oHUnObykPDqnhqWIMSbQ0WhdU5Hg6G0i+OSrzY+S+RNPtz2RL0Fio/C76TXMNgE5shM
5iGTmTuEsxBU1qPGH6za3+2EFjYYUsYsC4uiLPQ3hsOsJN/RHdqrYqIWf3EDKadvIUsPjnlJqNd1
N9y41ThjeJTFrNoZOGpR/kb2/I5PbEqBOF9kQrv3QjNrLPw30D49ykgZchEO3upfkc8DHSo4LqPN
x9e6kWWAAZeDjprtFeseIxz6DVhWvyM/uwzPhfwGURq1uqFD4ATSSSCVsdvO4AvAjInuU6EGyO9D
yzpmiVJp68Eb4lt10GwUt+Fxg/Bv1xQQ+0kil/GcztpC/YgdyvEMaDNCKtCplqWdTJvhLGRMsw/K
w4Eb11Wdawns/SA3h2lxK8PyyVlr+XM8T/fWGOnMwuoxFCCiUIfEnqSnuOGlsVPN+FCn00odHjiW
F+GoifRJo6tvP7nxPPRSyTZMvlD6oVMShZC1QFnW7jGPYSYuNs/ZxHjnnLRhxCZRMAmHu9nzryfh
K67z0PyUcUf93iDZVPY8WhCkIWOv1ZlAv7KiqX+Fsev1esp5gySUMek7oT2jVqRoOmJjtSTi87Hc
+hymLjCZdMnZztxCLbFFFkM/jw5hHiBYg8sg5yJKwiqg/wKOr33UgpVqN+eYGgjMpJqoPMP/2yfg
aFsPRQadD9ST744jLjXi4DYYwVmRtYGvlz7ID5D4KBUleJ4xycO4OUUxJ9Enm0TwkyqGMHiJ+Ddu
AFYM/y7JjXmpMK6A0EFs4/yQ5EcqGpLir2ekNBo+hh3t0Ew69o7oli0qOhJKCfUVhn+VIBsqQWUV
0M7E6xbRtiLqnlhxCKy6vLT6aZVSGakWubcqnetBeso1plE6iYenp4CXLetutLagUZyvu+/4VLiD
8U5YvEILN0RVfYi+fxlSS7DdOSu07YEQsTKekIvAcgTzEXjkQ48rmtIG9jg4oo0EXz/FZnq3qSE9
Lw5D0MvUc0WvkZ4k54r2GfakaAljdTxvRvo6LStUz4OyiDQNYYe4pKrZpcMZXbpa4qO3i3EL4ScC
ZxrHXFx8YXrsgZLDqDvzMBdrmYH9aYYyeAAD2/jypyRs8JCsEwkl7p/YK0bf0Pd8EEbuv19NGx7I
hHNS8uOx4gzfx5pv8rMZfcwY4npPdyzJb4AESTeLmqdArQDY+o20R2Z0NGVDoonehc9XUhv8gBQ0
WkDraSWZkTT+q9NvBQjxffH87rkyoUz5AJLg46Mn03D57pV14mNqhh7nWBsjCbK30gZZsJZyP9/8
X55gLtt7+3gj9taoRg1wxnS+JL9QdZX9eSvcVK73dpTYN2hAVhLm0YXFIfRGlXZWq7r74cy4P+Se
IZbXg7txv6rGg+t1K9HJoMbi8EFuYf6GlKPc3kHa5wKOpiqkgytAqhj4yw+YnpIdIlWvZ3x2o047
iZwUjcDJnSUU9k1Np1anPYJRCkrJYgry8GTjrQH6QRa4lyyBRYTSd5qUQnD9jFtPLuAg+M+R2LzM
ySDZH+ywujvY+szga+K4xhLUFLLl14k4/6rA1jbAOYxIUSNcINjgiCKzfsGwoXzZ/Vad+VqpuILl
DHow93GIUmAy6Vrs3mrUGIN2xkxP5IAvj7RCTdwHDZYgQCz+qugg1yLyhDIeLatj6Q/TFa1BuDTo
HP6/slIqLeIoIiKsWhHo3Cuw7XxIfvSjjb7RbSTeP0hEjvu3mgwAhM/gI2PjlmYpGERGrFuL5o/g
LYyAiR8pidUYKfbQKHCU57h8+9OCtsVO/kYrOLpP049JxizAkF7ecqPwkLcuBNWqVsoXjcjtvVRH
jy1kbKWcs3IJqfBt9y3CLdEBWRn1fSkMRJ/yAED3vBBcCz+C1F9gzQowfBC8+EzkBn7gI29ZZU1y
0FtDVT7IEmEGPwztVcyzZF2MSJpmtg34PrhF2qGZBcWltFpy8i+v7RHH2CZiig7SvrKayKThOYrz
tbYPAXC8pbz2scZfHXoxAU4yg2wRCvrYhzyAElo/6qw0Agpyjadb98EojeSEI68DtYH+7uDJw2hp
jKnlQF5R834Z5/JvFV2aZWHCHnUOhEJ+dv+ID0SIwT3+GHFD2xmPX9zUcE6YeWB+BJjd+mFOTOlo
0N3i3Ia3KBiCJ/++OD+HZZQQsGo2QDW1hKb0B+d3LvhrBZszYtFbg2VmvomnxKnk576DwRGwDYBA
8DAHnRaVthhidaJuLVLxBrx6oVmfzHTU6KMeTYtKxumXHkVQoyhEz0/SzVlBHR9SaWK1JbFoShIv
YnBDhn36ZMTkL+BJKfFPAr/AlX4KsqDWuttdidQ3DCgnw/LBaxGwyE/YRFNhd4vmNUzwuMzFL5gW
3ByQTi2WonNCWXsxksEWS8AbW3mQIEk1g8RWOlpCJ4AbOcp74Y3Nhd6A8QSe49MsOcw5E3DwPXSD
Vqc2T7FuV7YNmzSznehBeBjJeJXvsYFPN3Yn5CkLIIQzTk8KGd+j9NDISFhLMhSMCIdlaSkE4nYI
718wtwc4VCttfGAc0F4PnB4zi8syfz9jKXZirvcr1HA9TUlLfLs215BhMr1yl49dR4z4fg3Hk+KG
3yJWig4K07wx4KiAdMNvYDyb7E5iT7hClEfPAJkaIK3y+4TH8W6N68Duw+SV0Jn6MmzDbODdh/Vz
xvBic+qtaKKrbQ0HqDVrssn2Q8U9PPpbiIjNGUKwS+Om8OtWbBNyDodMNPEairiPgLNTbM0yLJQP
GQYMdW4cMKQDClaE8m4q8CUjiVGP3WQCtxmExTaDB4Pwal3sxTzwgRBF9jOPsC9qKMCpnaQCBymq
YGf9PmPP0gSvZ7tcl4spF8ViIPvhsCnzoyi6qcWq7dbsglUYe+tuxavkt1bhMVOc4nQq502HsRSr
Fe8WrTBP9x0U7gacovY1fr7lZKbO5hsT9N5EjVljFx6Bbs1xAH+GVcIV+C+J0XBHob2teMUc/wQh
ura/zR/nxe0sjZbiNmS0FM4NaqnMnps3XhZBUWu8OPafOkrMFCGldIpYrwYSkdOup55awDMLpoEV
COib8OYwdWwOVvrMmx0aRvFqk5U+yM8ib3eA+Pl7mG0x9dtLmB2T6vYsLKMovw7ZF4ze5z5nNqrm
gSxgLsM0stBeriymhKVNa+ac2C7ZDuZdSk4+6vhxBVKoquoM+Vao9LHQNZYfmESLWZMma0wkKHNF
ZuajsFvTDYLpVqgpzVbTRwM5HoYVL803oEYcz/NVcobdpZvpVcLI0gfs94C6iMsaameBy/G2+jCe
7tilqF0cUKN69MQPqBvZ5pcSgByaj54R1GRBIhdylgt/Rc5dHxKwO3jFa+hgkqzJrEPkWyE06JiO
LywWQ6YiDc2ZIkKWykEquhDpBjbnQU8esPAalVEEQ4/TDVT2IlsR7UQZjP50SVeEevalKloYQcEx
YrGilxc9rSUB99T5Qifg8o4O1cSPkORLeOuO4BAmrCq4mCejZcHJQ70vTYz/UgAfmUXD+4uu+Owg
AHHU7wPwRMK+//+WVBvP1CtTymYr/rk7qiE4r4UZC2TdQspMGVj8hPleiKxxpEtZG5e8gjcBZojU
i97xe3tMOsZMv+Jx9m/DQ0DSoYaY1mWHped47A59X/gwuSmY1PajTz95qYSSAhkfIzwIEzbQcoM1
sE9J1TFMVklwWjrOtAB5uwc6r+IOL3Q+j5ksGZhJ1FjU4Alk0gSzJulqFy4ayv+wGSu4Q5HTRTlG
VMtDZW22FE3jU7nAS1fgN6QmW/tgvksvs4Ka/3/Au8G/zeFoxGex9ALtYA6Anh2ATP72A2psBQ8X
wcvLOPvR1wVmZfGVResZn39fdjCWrgeMp8Q2y654XGHHu1MovMNoJ0YVLfXZPJK7CKBCxtqwep4S
zymg9ZHIR9yszBoxDaybzKlK5AzDsYVU/sdS4DQEKY08ql7qWk6y9nzJxCM/dr9rh0bkfRWRaAjf
May7qdzW2t8FjK5PamnyH/p5JiiEHEu/zNG2byyQEZGNbHsFcDACkvea9MUkx/Ee3adUGd5EuYrN
HP6zlXstTKnH0pwbXs8c7EgGfCxfv7+cM3jN/VrDjfkzBZ/J5hMt564CsDVVYjWRcgJrSBypbLdV
gNlFyR6E+9aw1Ai3yAG+Ygo67/yVz6PYEqJspu6aCxrOWwJG+wldg0FqA8IZLcVpagahH12wd4HF
YJ7szvJGL+2TpRutB9LFXewtrMjo/LHhWviS+p9Vfth00F9+PWa5zOzGQNy9J9JXfFTC2h4W42+7
P8hYH7umOJU7OiRl9+TbzT5hqnx/aIUs9LzLdZk3UOqmcetIrBWZsOhvlMw4WF/DHUqhh+hQpMZL
7rLb0vX0NyyIYVF925h8PrlbhRRgFR6MSXAkrRIIzLtrMXxX2CVsDL7UFEcVWySO6m+0EBJMZFAZ
bmuiITsLIif1puC5REFHtxLrTmMY4CnNJlmPSR4IKftvyuc2/L2cAtR//l3/f1Q2IKNPaXF3KamU
nPuDmZButmZM+bGdJnDBhpRNWd7mDDfl6Y0U3V73UxHBCW9EwcqwoRL4eJ2mjSgSR4I7AIa2gx7c
U6ePof9EIX4uo0wThYmIspUJsH5GEMKt5pSo/2GHqDxhq2KHCmalkqt4d/C38KVOWW0UodkoqygN
sE0wbfO4ohEkCt9/fX08gAhMqUfUtrJdKP816seTvJGhO3Ksr5XgDtWrpnEBly3UujvJaFTv7gmN
/oJJHFsq1Hr4yhNrJ1i0Q4ulTeUOqguRlvEZKcCRITLejxeIYiDT2EKk7Vvh2Tifhc+E6XH0xE/A
uyVlaa0pZzHK7EDTOBNrr/MDtg523CuDA9cfkb9523ho97kEOuDaV0H+lWXaC41uNpT0sdbXev67
nwLmmz8UnAr2rU7XpDc1th/tgkePfqK+xcsfMXxoQEtdWD5avsjQaA7pjLtwLtiriCWUxMjG//Fa
5Suuo8ApPLRihIiQY3pYajGBVjoHXQpDKvSzv7uOrMy35Nb+b9DD40nIrf+dXYsPAd1VAGJdM7t3
IOBdIE4uGMU0vJH56wzR0dm3HOaUWiP58w1v+Q7qV0HTh2HnrRvTh3gJlrHv+rt6nt+qwkaXvlrI
e1EZpQ1zQ3wFnHnMWVmhyxHQFL6kNjkLxNKI3j64fQvXfKRknCsvZ67ojHdcsgki7xpeG1lqbZmW
MoH5MyEzVkwLpfQngfBTw1vPajlMee60JRaT4zyTt37BkJTF6asy5hZe/zYY7tVmHy3wZXecbn7n
XKMBPGg1MR1shrqH0hzUlRT0613FZAsEPYw2YbPCUZ2MESpU/AS8RaXcio2YZ2i+gRUDB6Z2aEXu
sd6mp6XabdJgv3zONc7HUuoMddCoGm8w6VKcFFd8abLKdd8cNv4rf1lFB+VecaMqfRWWq/3HLPDM
NiE3kLfM8FSyWxcgmVCzqvdUw9d+Iy8cU5no6ylpBD7pYmWl0nnFey6N+CwGsao2flxD3i2Kcuim
0tcSuNFWmo9juUGpNncviHT3sgGfy3XEMJtyBzLTXbA8bqVzfiKrplQ44TOKpfnHoyVkKqYrVTJw
HJVjqdOpUHRYlaI3126gNQLvZUHoE52HbCOfLDEjTZK5WVWYPU9mjpJu8k2GHsiR/tLVMA9aACx0
NlAt+wr56IS6MwStKDbyZuHnZyN+ucvOxyoL6FujpzeQ5tTxhMbTVjO3V3b7kR0ze/+zyZdB7hGX
DRMVerjfS82NcL6GPlvbBUszatzJsxWW5My1ddSVE7OIrd3sWbGIsjsmuTOtUqFhns6oXKQGf+3p
bwp7PvmP7M5tPMJ7aMd81yjCdrKdoj5dg7IhZy248e2trBykrzv6wGwixU86ZTUTAoymxeF9reIE
XNY5dIcASpdu+nN4KeMK0K0d0WBjq0gMmpzoWua7N/sBEXxSSzSyveQddMWQlw9qHtV2u/coedfn
gvj2RNAC2alJUL/PRSHHSvE8I2jlUwB9XmASCzgtleRKDMLFsFqlV1O3bSp+XpJ2KuYh63EspFaK
3MFb9mXpEtSCLr8RphfywF9wKDpiKHMcrt9A04n/RMluuHo6s02YHkohOvpFW3lyq82GVSTcY2gY
G6SuX7f8m9F3ovyICYq/6teEE+vccsa9EY+eAkgdQQHWc9bpv8fJcK7OM/JvjwXMovoM/vrm+B1N
5ZWeAmyJFSJ7tOXbJbmYvAAQV4NyRGvc2uPD6gad1ERxYtZKlNtZV6XOXA3siNsOsroNoZko5+bG
tHANxycHVKHgZC8j3wr/eRnPqSLVMU4sjjMNjo4nLMQJ4c2zefrcNiKF0HkjoetS2p2sbTpvJ86G
8ch5pXz7tL/8lA3KJjqtMlOvPUyxUFW96LXAQjmbkVK7X/4nHVs+BHeqiGnMZJdpBr7FkRU9MWqC
nvBZdHL0tq25IAd7zVEavfZU4mY72sMAwAFVwRBSaBxFkKSOMAHteBmZ0H3QRhRWoLPVYKuqQq9z
+PdopIHUuw7TJ+7kqJnztPn/CU9qV4HxqktjWlFE+Gwzrh9ILxKMOt2AxTh9geiq/AwS2EJ0S/kf
ZukQDtGd9B4hqKw3w9cLMG69kWyhG8hFbIYbqDHJfCwsxcn1+gUritFCNcP6EZlAYKoRUgA1Ld+Z
wEDbNXE4/qtP+N2B1BFc9cl4XNLdgPh1ZnEkWdLCOBTjR55PjyzGkrs52iUEMopcfWKo0NDWmetJ
OahXC5ooCPz7GLZpOboZ2HXhtIHK6zXtWIE/KUgGkhpZLhYVQxlc6Tr64GetjEWiHiFEzMD9UUxn
KQgBYuy3QLhpR3AUcYFIZLqKpqvuGUQdY85YHcBHzi8IdoVl0wARuTSYjElo6GVdCmDskm1UiLKC
XJqFmM+xUtuQxSZRzHmXnlyN4LW9OP8Y/5tptO7MEJ8a4yQFY1nFZuCUfnCLDfwE6phJVqImXe8p
R+iLk0CMLcVML8d6rIFgDwfQZYsdQOJJtkVwnAcJKWUvcTp7c32bPHxj18xZK56rozMYiDRDW7l+
VK3Amg+fbSnj4VJmLKEclBjzdkURf8fkFOvPpqMc0idnSllGC+Tg9XAr4zxcmPTP0u0kNEUpYoCT
4X9iJoeCy67LLH94AxEIxKWyiNmdMaIBaVuLjQvieBhk8Zp7Mq1rN2cWpjP07yk/k9ALqaDBo0pp
TfRzyLb+sNeg23QXgOCgbyT43vmzz47FUVu17onreUjCfTTor3PbwvuFTBHlG4+6qtmQ9j6N4tJB
YjD2zcy+dzBC35P0YYctobjtMAz5XXBqOnVku7lTPCr86FC9+E4jFKbOAROkaOR/okH6cb9dLYEU
dk7fsmy5aao01GqUmhnqIR3GbuBH4tlWEH14J8/4vqo6ceCyI3+BGue7Duryv4rAVozstdIwGXBR
6T0EovMI52R+/KoSd5SCvrLFVK3ffk/ywalQiX68ISN+TI3YNoDYfd/HQM/TIFmXoZijXmAl5BO+
M1Ybi0s6peZLlsNJoAGenLIKJWkCWbHaimQy5uc9OIVmVpj/+SohXVB4vDrAqehqkn8eS7NG/zsq
mnAaGvzt4YCzBCpCSpFSP4ZfAB3He3pBW6sxxeQMQ9LSYG6dBlZlF2YDrMUYDPuZgWc4fqM4uxTs
jN9tcFQ51PGQ0bF713BWCra5cucXlpBHJZ3zLOTFke6J89IStEqsn+ZY0Rk+Ha3u1QGBUUmawkRI
SnfR9cF/H/qJC7q4IDzx8ErissUXa5+Y9r5g1wKXQ+aeVxnnhgbrg4T+9SLfN+E6qfMs0P1hJUgh
ruyaGf308RIWm8rpydTq1UBBpYhs83nkpqOpyNX0kNIjanZdHcEdxVhahOOU/QG9hRzrtU8xeCGU
O3KV0BrrN4o6w6WZSjgNbJWCVH7RmH+qKXiBdqKfd3nY04BwHFg5d4PdL4b7vs/dSsCt8bsoP/vM
Ytpadsua6GQBM9HxqMMZ/XMwmhlCIzaLdADN0ZCRie2mRMEx0TcQ8ePQRuEtdFUe1g4YAEYsi5We
RyhPHokx7e886cFTMgR3nQ1+G4cncyeudUuf5ZjApPMIiEzKrjCiMBsU6x5VEB3vF1dlvgDbdQ3R
TOIpN+5YFoIERO9lS112s2ugLBg4QlblFEQ+/bTVTXnwLd4jJ6DHAdPHXAPJ29v4dEnNhHQaj5jP
lyzXqPxVjJxoukHgb5yCHP+r25EOXmyjpu8vqQW5lFs8LN0SdWxXk/nNHfMgl8Y801y0DuSNLDPp
jGwJpX65XJuxpQT52pFEuT2FH+r94VAGre3Ch/45scEOyXRdtxMx9QQddOfUYdqQ2qXZhOkfsU6V
9d9sFxVfaYIDy2+RwxxUhLJjuEp61MlYGBoEWiJOYmUMbDKImvOwU+xZ040bS7mvaKISyfaF2+g+
/KN74niKTCJhwDUO3muCASDTGf5mzEYxZCRbH8vfDYZ8/G2XHTeGAh7Lx4PSm860Ifrq7xKSaC09
B4MOkaQJqonA5XV1Qh+tqBUeXBk6/mzs82NwPQoKqmqCguU8Sw+/jlOANfD8s3CahYwqtuNNtIDu
giW1pLif/3HXZ0m2wedNhRlaYaxc/J/bh/0FGijP5GPOtKZSkOQTBPObV7IoCqEhNHMDdgIqVG4o
8brbUTMaUUts1/PApAlkLzigRr8m0Dy9wyCAxno2gUuMt4isth+zsiE7KSUkZLmmsrJ69IO+8qC7
M0nhHul9GOyvGx0c4ydKgSXuMVGnn7iUup0EsHv006UHh0MQ445ITMUbVxGrOipc+5Ljz9dRtSgU
n/HloiJvAO5csYqysQ8itNJp+tUFDq+bC76ILpxGoHPthC/aJFwfWlknLHBtnH2ESqIMPWlNirgd
bHr+8Bt6JunhyjmWwOXqrGs6uWvROkPbyrOMbiWC2yZdnmJPFh5lfqRVelfg2LABUMR/AkcSeCUB
AAJTbXHL1aLNCviWUbdTBeDx7AHCgYacqwXbI0D7URdng+7lQeNSM/5Q1dOe7+PeqRIkfC/QfQMh
AXZL3krlDDAhcgAU5IyOSb8IB5F3vhSSQHWg8+v09CWECxXeDeLfRvc13+r1a3Fc0JU4h62zt5Fq
KJ+YexInVhdNr16DuL/alDttGI1OQPkfnqcv652y/xf5WG38kPuuP7PSyaFY8Zt9p37e85MjAkD/
/AZJ/sSej6utE03ZaLtzNF/TC9Gm9lHaMSuatJvmM2WeXEEpNmLOtWKgsFX4xcPJwMcIvi/q0qFn
/xSOh1Ug7CI0oxB1j58qpWjxdn0DQXWAa3TaUZZCfv+POfl7lkgqpL7FdIBBvM0nymbzmy0ctyJS
m85f9IBRUPND0Drz7tUxdj6RD3PV1eYh8gzvGRnuX5VCnI5gcwUwQpr3dcvWZ+FpL25RrZnzsD6H
LlQ9WIh1hvNaKQTjuHzW0meQ1NXk99gqjE8dnZifxO4+6wTDphiKZjxpOkwioYusK448soKbRT14
z1+So0C9Rsy5sw0R6pxqKifV/ucLU0H7xkbLc8RPwlxq8+cv10L25etVc8ir2hDnrF6dZkI3P7kq
p5bvLBZ9nvqqs/OHu5K+yXh4dxR5l0venpoQDqh3xF36AGADpCRB/O5XWyaqLtE9uLUeD1SyQKu2
5UGaOtDdh+JDZIMCDAggvkx37dXcChS2Ap0TAHf49sQGDANxF740PsHZHQrVJmzew6bd6aNAM0sT
1DA6VaIvkVFrxlRiNj+13G+U0tBW2YpmvqPT79cRGmKuUdnF4LL3JlX5yyTkua+lXnKxBVxK2e7r
F7A1vXaLOb/7ErUio7cG4ayS078Ko9HKh4CRz7n5FduKSFCJSj7eqnV6e2mnWii+8wjS85HFlZO5
TCkNBtngqaTsnYDnlljLOnH44Jmz9q09pthzJoqsHhv9pFXmLIH/IAOZJ/P7Wr5KZZNldJrb/B/w
hG6EudEgb16r+y/5IVd6D88H3ASZuAwDEwR0y6npEO6fmgqKhyRHlKkMXTvwbN+c7PgY03zmljkS
cAkK+vLuwa8EskkNnoF2ZBxME3kh0cdIvFhcVC8W0ZLVkDROxcvqPjAaA78fdnI5PcCXKFsYmxEJ
mKQaP2KTxniuKRAZF+RKSmns0exddzMlf5QArLaOf/mY1TR1GQPaUCojLSztEtd6M6/TdygzqRN1
QFbe8rsl3+8B1EVaEfJlf/IkYUwr0/AE5LihYZpO4MnlBs/TPWwF3gU7IlG5+8qglH1yQP4/NTbj
fBV+aySLNxhv+BWHM0kpqfrOoP/O/2ZYMvYZi78aOOssaW7wQC+47NkIaZ5kdz9p4vchsvb8Pwzv
LToSXSK9wlW1P9AnysbeNDo85CPnu9GWJ2swB5Q3qIIXDoHktM5Iz2TZHK0B/UN7vZtPrJopS/NU
TdjSx1cZODQ/uK4pztVPEZOGK5f8vapp0Ic67Udw8YDeHepBEzXzvRKUMbmwUr3uq0CUvVbLt6cL
U3KLDsEzMovYppO0T+Vw8j1utC/1/D0BiC+eQYO9BSYd7j0FVPra5glv+Uhf/kun6TV/s3p64960
AKPlztSIncvM0Dj2i/zHNE5nM36GgpSHKsUaXrb6iVj6s0ML9gayaf5cwuJCNpRPsQv6Q6G48CIe
6WxFrVDCaTLJ3vQuK8HMLgLVWZOQk2hFgou28qX2HNqnqdyw9DPXrPnCuaexkQ2G6GkykSO9vNOf
kBfKsQRKX0Ykbcx2Rp3ciyn5knLWaqZlazRqzLwwDgp1pa93BvJyozj1iCH94HL83sI6G7Jxv5L+
g32X9a8dS63DREx7rLPSbc3TB7TTypt1T32vpmZgRa2P1csJDeTdwujGdNd8SQ5VvZQe8TM42LRS
MppQbsABjZQQwq45vWjde9XUYcJk2RZOq0uQ3l89o+J7od5CGOAR5CnHRCARtC2r/RDC2MUjRxZz
n1x2yBd/Drm+3TtKs26iQil+TAG5+ud+WCtoFPazrGPGqaBtNcFGpq38P8+YOADkoFP+x2ZQbG6a
6hZHyonV8WCaPCfGFlrXHVWWLp0W72f86JYxYYqsQAi8hDNxMQdyfqWBwiAcAdXBTRAGbxsXNvcN
DZyUK7tCG3q6gwXuymZmGkJ22M9jFKasQoNQ3t8LmksROgnF7s9kW9h9h8qnBVInrcTSurIRQWIl
q/fBO+XpaM7nQ1z/lHlODBNxCp6toSJIpPwQZeQ596HJButAWubLhGhDDtwcUpnxU26DwHazmzeL
m0DT9HOqzqwS4WN3XeVqVdJ9bdylKV48b7m6EL1ZRVez1sAe1bihB+zrjViYJO8s2drNC0x8i3Tb
UCR8Y4kDoma2NN0Bf+nTb18IFF+wK/Gts6K1GV12R1Wh3tEYuibaITSI9qAp+NpnDja44wV3FWVz
qVVEqzJwRoWRLpTEzqZyaF6oKdT6T2/WFH2ilX+EgVoeBkkJYzo+RnWJYUECslBO7cTRnc4pjbws
znvDKwbCQQJ2YPXxZa5PGztQiF+XRvUdDMOd3ye0qMsc/vWbwoZ5/+i0BuQpDfmJXkomNL3dgMxz
aajJ+W+w5nN0Gii85dY7d/XptOJ8CtHzcvueUDnIscuCURAf6/8e0dPqbfQHE7s3Fq0cj220lWkA
UurWN4OCJCQbBQXRwoEVTE9S2knb2oxPMCcyZ/uawVhNylWA/Jy4VlVuIYEqqKIj0S3oER4YPWZf
2hlmLNILDCSAEje3igiBW5AgIKxTMcrCIVAbKdOhlaNY2ydp6lxVLFK+jsJ/wIre+AQYUrKiGGjI
fqOPjnvM/R/FFYDFn0PzeC009c1RoK+ngH9qXJUaOjzHoBWH9lXSZgVmTxZ9Ftp2Y6lRH+VFRyS9
f2qLYJJzJ057oL1PilZBgYeeLEMdvO9dezhcNrd8nrfPCTQZlMtbW+Bc+QfQpo2eoryYDXiAC7uE
aRm7Z1SRpf3e02u0g2WKq6Z7nZjbJpCNx5xCxM+I8mOlFp2JAUthRiE96CPiKOh6ZQZoNujQ0esR
EoMxZFX3VQI8CnlZlRMarMbxXouy4EaS1uRqy6QB7YcRBXrJ01jBK7eja5MRkkfFrsQaNKi++Jn9
25pfdRlLSZnqOsdKwJ6oHpIiX8UBiK10pVJMDvTLnWP8cw6DjiG5gO5vYUhqgMjL5FhJEf3FY3Oe
MvdK9u2xY7Iy2oVpsLHvjtUhRW7CWy2Y1Rt1k6poXM3JncPUnUzpL7fl+/cCKjeSvB44wwxWSTIf
u/dZvwEEGcgVg/R/DXdFII2ruVRn63ZzrhLtsx2RKlC2WrYpgRWkUX6uSiZIQSjBRN6H3qV5cilA
WHdWr/8PkEc2fj/frMxZ+7gfDhLUNRTuIS8H/FhhiVLZEeu34N55L3YaqBicpP1/EfWPPmxY/n5g
876rO2xaVJf6LTq37A5Zfa/5cPWMIWISII2ihPpIbZfyfrhqXE759uEddUPS3cKM4jDsyg/VMpRg
dbF87aJyTrll/3vAdDDHV8bE6wBrE4A4Q36O1QrzsLVUA+jEQjACiA9qjkCWb7TsydhCsbbJjpdv
AM60qVI9mi8tAmMKnlukKSxviJRKAt49EomlyUZOovZzRZ2muV2vkjED3bPLsrmrV4R+Y9tSwCpE
80pr6UqDKnLkPvPVFkeRylMxylGcDwqKEMCslAKiXJOe3gleJM2hiF59zw1GXqPOgMK4GuzHfubc
AoWcVUTctbPgpB1TY09IBKcMkb31aiYcqp4LRUO4v/IzFvvQOuho/+G7i9g/b3MmOoi0oi9zyctk
BEHjx/wYAffg1Yp0CL8d44L/qfLCKz39Bh++/0M9BsZ8mzCkOJpaYbzjhqPqG9C2o5shlgTBc1Wx
lTru8BrCcJlM2UbtmIQO3FRTm8QuxL1XBDBdRawdTdHpLO7AkRmiFqy4HaCAQBWtCcguh0Us+dPb
nx2UyB0q+ZEIVEmWLU4Nrz2TybHZD1sS9EQoAx0DJpL54uZVJTr93Ctez3w0tAo9a2AOoYy8JEev
eFidDXQsOP5CVgCULqRk75uPvM4gv+84+Q3zhGpS+NLr4uPQHh6TC4AkX73kofCCxaOXgqaNPJvZ
S5azg4JwpAqfM5CNpKqQ/aSLKsol/F8D6qcA+1XUWaNUkndeKBNTHbgHiLy8X1TX6NAmtH3MIXAB
teqMCt40Y1j7stmunh3X0PWfNDrlbYAqCR0naF7TiRNi5YhTwErdflW5yZMR+VA0S6t38E8JbsL1
o9BHnXcRAKS8Kx2ha5mjKiVmKqZ7/wJFrHOWtr3j8HR+RMT8f9ndE2ZGwCh0s4ALDThxwaOFKixf
/LCPlpM/oa0cnXjthIyByC3wXToYpPlKQmIfUqA9+cdtuZ6IopsGnZ5O+hgeSIT5Yaqjp6epzOar
4a+HFNOaQQ8OIYDGhMXsAV4UzBWfmJiioKJFskYEjub0sx1aIlMgONWtuvmPuzi4q6CC+r+XQ4A1
GYVcsRllALI2vi2UJgy9p1oYZCaE54UqfT03PBgybzpnSx63TdE5wHmpjm80cEVq2dizJ6ucL9Km
ETcTAwxWPBeycYrVX22VsVTrPIjiHt7Rh7S1b2LAt0AAI7XBIpRupuon56oloUZecjNNHlUGSbM8
lojsiwzOfsH5Obg30r5HvHrb+1lRq8tJpIrbSTS4NKIyoxMskvCatdtfuMJVUBTIFFSwRW2Tvd+f
h9qt9bV3t4LgcPo7kbwjVDrneN2Y5PhtXiqw2EyuNRZPKB+C/aeuhaWl+VoMq0gdnNHMVJxS62sF
IojhI1u0KzpjUD8nL/IdjDGnJzt6Il67+bfKCPZPtEqMGR70m1h3bSgE/Tm7mVQLUhTVibtcXOFa
R0w9pdQrIbybo8K3s2yHggPzNlW4fQQDcGdSKUcKZz7Xr31HkYXbGrUL8D7Jvw3gK8zNZDy3UJjm
OV8UsrH2Ktp1C381JLUQlWHRPFF7GiP4fPbxfbcsSPBim6HQzjgJZnFv1H1tgRBD9fWwvas7Dlob
DIBQq6DaW3jCGoaWjYNmi8v/XENOgLD4QyU6CjUs7g+ExBKbN6VFpEHWUdjZ4dgxb57alsqcAN8s
up+ZAfI4bwkxAu11GVjWgGWZx0ENbkjtpveGmljwLhMIi+jjLp/aNYQA2BOYRhEG9op7tiwBGIVL
aunXk+oxZt1xQJgnKkpECbRzp9QtL1HU96GAXiBjMz87M/H1vYobPTZ79C+CzEyp5AYQJU4NNDcu
iBViK90QVSlKtoC8VeFK1YW/6luj5oX5tHjVlpbuiR0bItR4lohTQtcKiy8UD3LjyMqL7OCAvq+z
a5tumlqeINaIXyD6gvQClEdX/k6631UZO329R81MEMuLnEv7vJ4iDTNbs70lOVO2ipcQ9xuXsgHs
kIc1Ciobpa+WgxZF0H28wCh6dglnZ2SaEm3/5rkWJgfhy2g86CQ9IL8xN6YrBZJq7BJQp1EuKiMk
s9NawllhROxCV57ZX+1At8oMnBD+iu3JtrO2fxmwVaiZIx411UYDowBytt87ZXF6eHWQc407bZkx
yiP+DSzC1JPCLJQQ5TbUmOWdSMqC38YbN0SacnDaUEyI8yKdRq/a7RvC+zmkrvOUmhBZcxBcw4yx
IZKwvVMtSS7akGFNhbmzemx2s6Q3Ee743fKedUieK/+CwRZld0L4F9QxejQdc63tufl7nVvzILXh
VjaaXYzEm3opocvSXdUzwWiu1Ik31ME3tLHSS5DNNMWoI3Fh7MzvYkg/k4ax+dw/7EMqvXSQPbfX
fn+522GGAoereCB8pqkIwsiOoVDNU4X2vc+ZH63RGA1aBmkvH5U8pHlVjXO8FhXzmRvhQbBomSBE
qYfqhFCbU2+X2c4xDAcYK8fcIeFxr8fuQ10OWrFyevmL7OeTtW/sED0YI/hkoqpBmy71g7563fGw
Omxg8TnjVrL1zeRkZJuPDTKhVV6OXQoQwL5JMR7pH0FIeJVI3jyd5m6hYcySLwMR8lfR1d6U/I60
bF9OOOtTPDEw1uFvwLxioxD43/ngnfVyoOn3PaKGuWoId008ALilbRslWTs/Zy2/9YBZs6/cSpY0
eb0HIQiq0JMl09U/qpKTT88bH8Dv1L8WHDAsD7lcF70jyDp1ahudo1g5/FJZsx/xWGjKoGdrjd6p
fg6KpZh5m00TY4t4TolZ5KdYIvsQHCakWB5MefVZZ+cHtQDv1ZWhY90GIeks3QFxY38kEwV+R5r5
Q/oMKcpuP3+9mbOdJ2VB/lW782Hsp7cKqgAnOABzUuARvQquLPjMbl2NDpHoDorYS6VxvuwXMIQE
gY1aJkdJTDW2FpgreQJC6KoDE/f5PL+rmfVRx2flWFjXTNJkOBuLS6bwoviYrBl6paeKxM1gUBC6
XAIHOigbv0DTbj3asEhqGH6f0J7f/9Oy/FFNIQBZC9Ss88rzkjCD4kLhBNByIvvPtjQN2MDN3Iho
+U5TIFfTj7sHrxed8eOPT/6NKazWdXgbigxmHoDPy5IIFNofQ4c9OY0bcA2SPT/Zc6bzG5Uumll4
87G0NXZ8vpUZso0L/eilyCzJi7bAXys7qlqsPWF1opGNoN78QNaV5tDT1ORVAYxeJ05mk3Qi2Otz
d+4U9JPzI0Q/mISfBlpI3FPFAFNvNOsvwlj5n+yVCksECvH4UDlPzHnz5tWB3qVhOz2fIR374Zj4
DMifMUAku0s8dF+lEIHvDG+I2NqWGPtPObePnbGYI1e5D8NP1gBXy1wDze1+tfG7zzeHW0gjK/XV
GFz/rOqqE1wSrMTFrkRIxuposlMxLyfzcsrk0tbHq/eRwNUh1SuRanIB1y6v5i0Ek+aBXj7xYS0g
p8OLbZQRbaCy+RUzCFKkaCR5JmgVDnWXwK0NlGzeYjCnSAMnWXjE3WZ7WxxlMEFztfu1Nx13AscZ
hPKjIA77fDXtNfAHYKT+O8JffEsj4zBIRU0HmMycNfzADJnhmQTJ9uYZKGYnvPUQEilWyj+LsSNp
8ie/py9Gj8xA/y5HJBNvYFa7SUox2pIdFZSW18GWlhgSNGZTyZP2v+AXmmboxZuQmzKhuRV8KGWU
/s/G88oy97/UESgkb/qZpfkNDtGsqIGsZEWhRHQBY+oozHqtXb33EnL3jmjGum7ecFc77g46KGS3
wsMhGBeuTCxeeVD3DPjwzOvRXAac8nxnTy/mQ8LB/yTRvkhF+BRBRsFbYc2HOnBjpCAT7bSfVy5r
tLADvT/Bw2CTBe4b3m425cYkJ8oKyOlcwTQ+bTHlvGD09k1Xf86Sju+nI6g0FofHh8L7djV9tZgQ
AuR1lreGP+nInwuSLlP5OURGeo9waIwI1UjOjqdjfsfpQ0jWAmbcHobTKNz6phU4hoBvE7JJVpEh
K6Wh22kI/MvEL9hh5Zor4kcMpuZOmgX5vvSSIg3HOODrCl1BSqMvIMjNAJAVhiXPuzhKUWO9MFD/
HoffHDAiSYOnlwCUJ/IUIWVxIxBILN1Q3v+OtivSGWEOCmbIs0Y4QKuKOnMaSxdgBf5wuFmKX057
9IRHHDlNXSH9szfv9T8sR7vRu/u+sgibsPCAxjeV31mwHd+6KYEWl5kpMK/vtsGS24/BlnCQC3JL
7WHsI+f0eLGWUD/XaePy1ySnHJE3nySJ2sXag3debSHU572NTYXqIksM07cFO875Qy01m4yHXkXs
hZwH18oDsZ6nYR/uAtt6wejU2/B8+oayoWmoxWmxX+qMk1SRZIflgQiqiQWXG/Bos2kt5cNxky29
smUF+IG2G8739K89Ey/E8WO+Diic0+ur3apvI8DnOIjoYChQI1eCz7ST5NOM5Mfbmg+6PTBN+kZZ
eo6kvOzuFy7aJ1/iySUznKhfWvQpYI5FJcFQbXJyXHikUokEVtyWNf92EP0vZdQKA+CpQXb8JiGE
B6imu8g4yIo+8+Dkv0llnRh7NauR3ARie0+sU7kmpMbSItP72ybV5POXW1IWjPxLmnUG2REl9VpJ
75Lm55658z49zOW6e1A0SdN5zucy3DjtQF580X3k8lv0nt3FRvkitbawR3owQNsmCBNdmzagof4h
danTDzHJCuZQtAtNxTOgAmm5IpServv3NveKQULLuWHxxEneHdKYBOOsJOCovrCgptARwOMNtvdN
N0SDzHK4etYjd0efcJyeRE1ynTq+5rkKm6ThmMyRqVHNdHJCjnoZ7C5JJccHhHC+q/TFIvZ+NsvZ
uq+fJKx2L0aCVQv/PlpdYKGkYo/jcjM/j5GeWLF1rQfjtnzntxqEiVDWqAuoNpZnG0HIZgX3f8MC
N4XHcCyYxHq/+axmc9ldUiO+hNLZYLonhzYDS9cf/1pyDz2VmJxwt+VVml/PDjEqu7NxkvFuVgje
hIoF2RKlhM/z4/69D1RJs5cGCxzZYuVDMXIpPPyrynvlMWy/6VL2nvotMaIbL7bTunBqXOWG9gV7
n47H8ZtwCgS43L12wi1uv4Zpct/IzOgq8b+I8AcQkfo0XUWH4m2rp7m8NoX+Bbn87CNhvmHlzewX
ElPAhrpYkN4tKVbNSeYFLxOtD4aw1DDJUwtPmr2JcGxXb6v7pshh1PXLTr7JDel/scoyWHTk8hFk
gxtePfcO08Hjms7ntdwdkuFrf/xHGZj/WCsEZ7u5kPFLBlI2rLP9rHiNyydEa6fEjXScXc442N/2
yr72SvcANfe+L2twsOryBCZcqpmKC8Mcc38aaQH9IsJyPBNu2IS/ADkzds4pQZb3OZjxaGQA+eyp
FAdii4VpeybP53PBIICpR2/IHH0WiGwdH7b5pyNiQYEyzcPWsLGsnyulAJQtA7WWonid4p7ktSQk
qTKUtGrGDK/yWZ/c3tZCJoUddrCP6P4dSmQj9u0dW9AhX6nqNt1lt+ExjCkkenVKPm60LCrX9fdC
Mi884UarZPs2jTrjI95+aplkF5We4eCxzPNq6tf1jWfz0CPq6I0zF4b/rWf/f+Fn8D8VCkf8JTA4
aBv7Qh7YQBr9tnVT2vrpEiq8f0RqAu9PLPs2DWzcNdfWlNErj7bS8vf7p7QxaLYdpq5G3m++ul8Z
bsCBbiRoTWO6VGkMmK+zeXS8x1cMEO08MuIsITFWl/NfXKgFZPApMc5FnFUJcmIkLmcpU+gjmKxL
gCMzUpQuZnFa6vtWbNQKhUQt/0pdxpQkhjSZdmqT2zvgtbLkXlvjRdpMC0EsYpYxdK8ycK6SV/bS
jQYcAWtiMZbEWXjeqnQX6DplCdY1WSToL7yljThgscoFx5VRwhzOsKiSvf/BB9mQgxZlyy6c5ubD
DKEwSS+SQg/sQiJMvP2ZaKMcm1e7ux2jQZNDvh4wSr5axEfpo5cRAxLrQipFHpRZC9omeB7I7Reh
Hq/c991R/BmXb3L4VR7rYUCc9zBm6rywtq279wINY9GzmWgwtvvE5Ek8imrOhvE81xJuJtko/3RP
p95B2SY5EDzTkvxcGkiBf4rtv5Yc7e++XZNpd+tpf9mZIvJTVs+VpZFnR//2fzV0kx3LxclRHINu
veT5LAvzN5mprNjHRoVB71WNJUSxII53pwGky8l0ZIzQhNC07l/HaGRfvz1GiLCJLxILDR9CA3nI
TFcI4MnWNh4BIhQ48xU1k+Y2KjpOz170L9BnP5kLyN80r8jF1aNPZHirt1sOPdLbRIDxfKdOHoHM
sg+4i3LcuGWiGQP3ZX2O+zctyHNxt1Qjp9KXGPDNhX68eDaTdPZN91mwNzG/0L9mHGUpuB9jtmgT
bFGCFX8S3FhsYf00UNN5xXlJLwztBSmoarTCvpvvF6JM+zhQltJwtvm+rCDb1+tHcxOZSu+UBiOV
8EtR9HtAo8Chm7i8f8UhWme15691ZoznenK+llQTOp0v8EBjvL7ASYnjxTy23R70J4MFX0tU+LGn
IxYDM1yRgHUFOF3xVi+Tal5Ey+u8h304e3as/hYMWkftZ6sk7fJb6wAZXHBnevjJwrcxt90GGVfW
ja29tiGpyh8sPJmx4VlmfhNhpvypp/Fo2yBMsRdjv2ovVFlicoyiG2Tg9SMer3hiqZjR3/4sRlB/
0qCBsoBQn+nC78vZR1wQWztF8sSUort949tBNp9lRf4SP7hWwVma7IynDp2qaQU7a5okkz4doPwb
sRDjuTyt52Uly881IFrL6BiXNjG/FAeWdJOTn1ml1iT8uj6zeAYkUSDpiiDp3ESfmxsV6wQlKBt6
StB42b9eLQZ//eP3Dd88S3J/gwbMCfDpqACE+iUi4nKoxzP7664J85zTkSsXw04oVN2VH3YvEmTM
UBlOYD8B9y5LTWRWZVN1TTczck4alakPMLcqabAkFRMRZyL8cg9/JgaShrs4O4I2RpH3C6uiJuIe
y1jXmR88n2PGhlxrkUJDSwuAO+DGFacrWtp/XtXZsIh+PtQmOVu4uhZ4X/0ys7HUccnijr9Za6tY
nKLdD/iSGuWwfyVB5nk7NAfwU+MAqWsm+kT/fmuijBSSKNn9XgZ0SOMtbIxzzAJp/SYeH7xg2hIp
agNBZfLT6couZjGiVVY5gmEeF86V8avR0E3m8vZ1xT85Z5gzDRW2vK+6Ijmno+EfDim2Zc/AYnc/
Mkn0bdMIhj/grAiJKUark5gjnSRN13/bqjgcFI/5tVF3G4VX18zz2lhtlUeE3NJhzl2/YJiJeGKv
ue8bYStFVL41+W8kHHv7MRmOoUFsq5BG0XKqtXBUtx+Xt1rXxqKEwSLGc0DRpnh5KOK9iVzyWAAs
u/NpqjjSxmhPlapbtgjOZqzxGfpTVcn98OBGh87IKB7GKIyqYso+5sGZ3gjONAPZPoJUVTdFqwQS
optb5SsoRgCyr7treJ7e5O3K5nq8oeP9WdyZG13eaLSRgizjf/H/n5NDf+MO5K7gHFLu5S661hqr
g2kA55aWAtWm8Nxmjd6lAEtDHRGBmshNf82A7ckub7TOIqo94CdB0lMaLtYxuijHe1fn3MzrFN5d
jh6B2vIAfz9AZgbRp8mnxIXL7REKeXYzf2TQf6oR79bUQMdHHU/beOY4c4NrFACfETsY9xb2y1Eg
xwsJrLLxlFCSRIx6IRh+P0rbaxB6DTdnVmEpuffyyPuGMB/EwTHGF//5dxLE/ZG+qgR9Tt9mFUDf
sea73uCPUmW8zYf0yYfzyMlMJf0ZQSfdqPhw7yDIpX7fLFiBPNYpwiMUoTbT7+xpHnlwIfuQUMPf
t987jGAwkgDOKsLaUcoDwK0cF6Zz2qFStEicF2rA/jL7kLfejzjnF3uZIl17Hgk2/kFnhTgIUPaB
aqMfKgW1vNWJhn0pZFLW59341GJDvdzEgeHsW+1HnTmkXoaPReldGJLW25HOPVXE2472731V77CJ
FXLamBUjyYFoPpTIeIMgQzjw1XQEJMMAcSkYTz2NY1Hl17QvpdT7FGLRZ6onzWGp0Kt59Q2rZxam
th6M8UecyFI2tQCz0aNyISLSt3//eyN9+kxhjUqo6QsRHp1z7GTsf389lfEjdz8McRth/IwQ3KF9
F8ina6Gtb6Y5kxnTyP1rLjayohfZD0pN8WPeW4eCczHczmd+aL2Dd3PTH9HRxgmWH3dvZiiW7W4z
uYXAMO7Zw0Bg/jwqf/sZKhpXyFP4Q6vPHHHlUkyuvZkAQulEDp316jkoYAgXuQu/sTU/CXhPviD0
rx869NXfyeEwtfBtQLxRTyM4AI42eYwrcvaoRC4GCEY9Vs+z0b0HNW8WuTPwoqE5k/bTac8z3JbN
b9PbHQ8YAoH4YGFIhd8H0nJc6+ovS0RZWQyM1fyou0WdoMWcS7NVQsKha99PD5l+9crYFocmrQIV
5uXhnkw+mOMj/Bz1WBIXb8gEtN8o6r9keNxhiNRwvZ+/HW/IGYsuYAv6bcPgcb/rWMqSbgWeIs4I
ay9eYtTsMP2euhH9YVwNFRAjl90s18gAf5uigOo8eq+smDoAPWz7cNEzP3kh2aLGPtbZGPsVswIv
+74n2vh8/qfPTU/1TgNnyezOoh32yiZV11i7+oVGthjbuI7Wa0W0lpNFDZWelbWIywLvFWPRA6RZ
3JzwTbhXzbDNai8TfPWDrL1NnqaHsniOmyhGU86BZLRsNQGZOSZ4ca9/PQMyW6/T4+NbTrQqGgvl
MN6Cc/wMSh3udReM/rfz0Ng2RkwxjKTHviWEV+J4+jrxJdzGR73/3bWSWplvhz8XZBkaNotv93uW
FhlXFKR156H+VHDkbuMrBHfmMkOweXkbGG4tYktqyaHji7B7iWXY/Hn1YFPjjj61/smvVhDKUKa3
T43ufbLGCUrHuVUIlUxY8/Ymdmqcp3/czDUO45Y+X4LGFuxuTw91a9h5TKIq1YQg6OjBYaB8nJRN
9gzia89pmfyTjV/yK7VoL21SOyh9m1ckZy5hqWIUUSB1y9fWVgr3dxLn6LDJSG1p8QTvkcu/ACtv
Jd7JFDWHJhaXu5taQalqyXX4dOlbUK2z2aVXVrxv1fqAANrf05kS25gaMUr8YyG3bAgY9I+wLjZt
NCMXeDByFZg6tFaDl1DV/ca1HJmsUT7ueEjAqK8ORg4GAN7ff5rD1UZ8rtX7u9qMBTqUQsdUXfTa
ZUzPrNPUCF6w/FD1UEQMyX0DF1i0m6TItdhvo0Xj8oxw3I9zC9wAIq4+1C+cLUZDY5cqVdy0TAsV
dt9tdzJuR7r4VW56Nn5fc0BB1yR4Xulxgaf5DMf4Vx+hcnuz7PICJ/NSVOW4JqUxXhwbvRlKDCIj
y8UwoxvIn+McZWP6FBW10uXJmgVxlZMYT8cWw1B4nDyPsj8a/7DM151MWWFjgWjlS0Ihrj8LLwU+
wx5YewwsJJv4wJzvWsVcwEYBROA9nChYdx19ktNqWW7NoTnqrWrdh0Cs0TtmKBv42AjSQxR6mnWS
3V9eOWK4gVDmjmf3DZ80yv6byKhuFQ1mHXd5IidnmRldqtEAxz4jRAMuqq+RTI3k4H6qr+WrwsVx
s+WoUOiTOPSUECLkYxltCO4CJxG/L/NWXBKPEvWI9L3P5WywyD/SLAIIM12TPYKKlhMfD0rTNdVd
qYmVtQ3VJCBOV5Y99Pmutq1QNJj3As6exmTc1Q8B+KhDX+c+Is9Ur7vicFuJsflkNEXoPf8MfaSZ
E30iSUAthMXgJk/t9tEH+U+YPzKfq315jHsWJ6vMo1lWKDSgtxlQrI3WtS4rRQuxXMPX0PeJos28
WQge73t0Hng5vQl1o24tqwyR27dx1NCxJdD9+q4TZS31BzyueLqScP96ydp0xo3WKIxoCFlKN7r5
r5OqXb//23Orlxkj8DBkhNnPvLSx8y0PltUDj10jfnHXypKLQM+ec82FLgroNbTdgia9R3MMq2Fl
L7zq8EjhYQCl02q63wwGKKf4omyJGmaF6uIkpj/ZXSoPEyJJZfXrvMME/fTHdneYiTdatwArGUom
suIuDF/M5jHqSEroG7XbXkjkjqIW4S5ZIlwS3eDA8C3ffyr+kTyxmpJBmUr2n1TX+aeicsXChPJZ
j62G2wjmLmiF+ymoH1tnTAYAUe5OnC5pi7hjzdjYTV8kxoVTP7z02vIx++xfDtX/2CQn0dMLVg5N
5Hrd+Q3+7ZNHC/HRYtp/9+gU64+vxni7A+FzsNUDGUfaaVRTmwv7MbL3fb5GR0ZbCnMGj/Q+k5xK
uh75o89F3vjJfl4cqGt2cC2VaTFMYlNFZSBcDanYf8wlxBv5iXwTfgWlAYDH2h/3Wa1dFr9SFTL9
1Mam75O6tFWt1HClWqcD6kl8+h1VeAoPzHTIU/0is7QESfEthZUIqGKJdxKbwhramNQw746O3XCH
EIJtDeLhlGvgpLe9LEcIJ8W2pTc/Yu6zMxhfrNBVuyY9wJndRHun5jTOGDymqsudrxx71ccXdZ4p
/E/RGPBGNA0/LZLRPQlK8Ay3TPTWeOYENBrDqb4Qc34CBXKfELdRv2Vn1MsdhHrlb8ZMq28cbdlI
KxQmndcdNkyHcNcbqFrkKMg82sqsyfxJQ244KBpy/dAQHWItIpIdHBw2UmJsx9L+R1NXGY1dDIvz
t/6xeYMtaj7vn4Ia2GHyS781GqlWb0hphTBfoo8c8j2+1KeS67+AE+t3E4+5R6zw+f1epzrPh1sS
1QXKGxQfwDlnB7migZL6ZQrv4iX8COrWrtWnplpB11wK5CWiIuBqwshQMSZ/H+GVbpWBLHzxqBg7
2bpeZozQwyAtLin0x/kNL88rMVcmnTzPSZ1ozoYdN+w0NcDYJe+4g4rUJCo0N1ahzezstwkMEn3s
Pipfs2fZnJpcEMAkM4vXneHwoLYia0twVfxmH/Knoq3UerqE1ZHbrp+30sP7zNcFBr6EIzPGg2Td
Nwj8PeUV7Fy3yq3qPBctkygJE60vlayrMxXs1qcWI+6IykxidoCSH9EN9B8mTq0VvAb0G095s7nb
sei+i37//ilTT8Y1OsyLARsBsuu1MGO5zJ4RvavqKiwTcKks2FpTOT8tvamWo/1vKldL4eYwpRwf
G2Iid3MNoRC4ra8oamvVNZ2Uhk3OOaidR4+mHg/9VoS4b4U7LJ1OfhWytu9QbIJR+cqkRqjcaK+Q
3Daaa3IFtD/7eB/nioZIZz3iGGbpY/ET41kLon252L7WBOGNrYa24umVOLfJXos1w1O7liHAh9bx
1IvuwhWeuC8NAfSkwy/CgEUd1hhk9kXQyrMrTvPf8engL4bxEi3snmn0E7emTZkqR7ymVHjFDTPc
uRtZZTtR5OPwSXgf9rWfiTCG+kg1VGeaJxH/gKeWDM27IKDTEGIAqSFUUvShj5h+8s9s4j4DAnzz
5Sz37ZcEQQlJG/AOqfQs1k3n/m8wBEFpqdfQDep3WrP04oPMLCh2FmHRaZCkMtICScpLPs73WaZK
qALxTGZzIzFM8+XZ+RHU79h/9xTWbEyiYnzReZ29WIQP2S8AOkKDfrMr1WcMzacCw7g/DyL/9CKe
xoz5ZEmXRUAnq8c/KCKBgmektCIqr9YVaxF5pJEZanMgzsA/sJCK8tag8tT7Xm6gF6eeUt+D2sTl
NfxFA6YkfAfAwbnarqZ+WMGedrFIbDVGLar+N6wnsdzQQHW8jovj7D6k34h4UNfLOCFoDRBU3RgJ
7GMXwOJM1pBUW37cinjMPeuJ0yXUKZQc+khTqkLAtdtyPq+/0uEdxnhipKG/wiGG9De3QiMULLhI
SBa976VG7KNg6ekcDFIcj2+1vaxzqH1sQW3k+T/OyxhuxiZR7PprKq0nPCHXeV6BNdV88Bw/vWTK
dMQCJNc88TlHyAYBrYhJb1QzLTGZpUeoJj79ff4i7nV9MCkNzt3XRF5qKfYc4BfkxdiE3P12bmVJ
agixWHAwNJWjpU9fyFsU0upgllpho4qbKfG/cmFriJOprgPyiXzgOHKRK/6scrzqMEUUXlknDxk4
R56cOApik6fQCTB50YKGM5sIm8lAkmyopxGeEsCva0e/9Dbx/QNcdRId7C9YCs8WpCqKCLryB8Tz
rGJ9NEDhWcQe65wfdgF4xxVWkuoNNPRTTinnlp+aQG8y0G3s2qb8cMkJNUQvMfioIRvnPGukMybT
jOB6CfFqfWTm8nOSpaRY0qExTCZIQeGV/yt3dNGA8CC+NGeT6bPS8b46UzcAbVT7kuyHNvGLO4wP
uIqn9ILgK/ijY0zJKRZzPggcPCyvna5lQ+FISTdDJFnvJqvxbZlJJNJ4OTr09qiqEbuMiwrMmY4p
51d/K49WowscbTFkgPu1JKDJelTx/nmGmFrGAc6+oaJ5NKX/Zxn5M0vWMCYXnKbPLx+66a/BxXRO
eayaVNYhjMyAQFV8SOmJVlVtUhuAKEyFMacudJdXMNPLoNGIfFOwlP7efbLd81eQ1onAp/Zh2/T7
gd7mcQMFU8XqCv3d0vDxPumZ0hvswjGLA/AsJ8XWsngkxNii3Bq4voSW8FGB4+9+6nN2OekA5LJu
hnCcL8gUinj1WNvTCgE+4Jj5aGSo7xjlmWk5vAFF7FQZOQPkmSSDCH6R37F4w0cfW0VxHNUW1NKY
3AzBOnbXVS5u8zYlg0HB9BmIYSFzc1Jle38LKdTnwqcvkPh0rKghMhmSolWPFy9NX6eMHfZzBPm6
uMQ09OOjFjlgfMnv3fjZx8TTUXwspLHBBN6tv1iAwe2m4vsu+jgX/oct4hWxPu3JBYjngR4G0zz1
3i3VIW3pWFeN1d8rxdfAG4wcLp8l/HKwcn/v1iuRYPxix7S4eW7WucYdVMxhzUE32bN7j2DFppLE
PAN8ryMNQJeeG/pJ1Q/DymI/zdtzXzxaWMhShEJsV3t5eQq/7oXgddQskP502ZzYEtLip9fgCiZa
RIFQgrH/7auRUxI07fwiaxcxTYvG9hEIslguVW9sK9H+gHVBRFElvDsQSdcFZeP07sT23srw/vVe
4i+l98daTWC5YOUNbQ8wrqdtNr5o3CfGNBlTv2ExUwvgP4GTxALSfdziHOwUyta8bCRRggWxkILK
stcgS6xTEZO3XFZbWR4CQL+vmVYOBIBPkGFlRKJAO+BYJf6wdPjdvuKJbOPVWmICA+UtJ0WVrwF8
Z1PF18jqHX6rzg6PqWQRbiPR1NUWx+uSA4BQeQZjtPV0aBUofFf3xEyLinUHkXWtbezMTRS03yKH
6ukbCWdabI9L9ALl0UvCIeYEtT6zOK0/3D/duBPYb0NQpYmuKEc6R5H0Imq+d8yLaVx3hVOwOK6i
0RBao80B/51TSivj3HPrNC8EN0pQiRHMKmtCxppQiH2jIqduuk/fUGJBkD/aZRSfl9eIm7gpOLZ7
Xqe2W4hvQQkYYMWL9m7KLG5zi2wQhuxn/oCNamh70PVp1HteeYN3jei346s80rrkyA/12XkU1h3w
27XDwDjUw4Q+PjYLmNNy8CNzLxjbHjjGLnXvtTUf3VHb4bNoYhJ/MlGTGBA/Sq5XGkb29v6qlZUL
KnhHnmazL9c/I8VWYgCvIvWihUZHl1+ylTe8jGEhXaj96NS6A1+f/YSO09yeauDsWsyg6epmqaSR
M8WP30qtYoUcuMnAxqQTgqmMm5sb8K+0ajWEIVlOhePuAiNuiF7ceVzMHJdcEvazVWUauiQDqXRZ
2BnBqPYglT1T6HE8GCl08qe46COaALGLtnMnxniVD0F0pwRubvdMTv5kI3mqeNf4jlgTXR9sJlKS
EVQ96ZkhHeoZWaXL89JtXUbPE8xG0tI65Td/pZQrLlrVBoya58CXv8186rpN55sTJFQ+fisZB51B
WNmP+BVPhBychQhBX7ivwZUF5kXsugAcl5hzNiuZOVJqJ75al/Ncjffx6AJSyRIKks8n9WCxWrLY
zDG5GFmEzkfh2UKheXGynyl/I9f+OrgQvbuj8/ziCK/v2J3009ZB6h2JYgaVqKlwGBSDYBEi3Z7D
I3uIehz6TlpAhRB/WuwgXYCtYOcFBZTiELh6LvPjtjYV1IjyBa+EwkP0qrZRyzgHHm0Or3m/iwTg
ynuPMxgj9BbwExz2PMLcANSZkOoXUKTB+SZEF74JYcg87YogZ2jPfSdKOgn+oRkCrMAYY3gMKJ87
KIobz1sjsznB0dWTNu/BbqcepOgT2cmqh2WoYBHWPzh2cowWwyQp2B0IaDzlOKYtFgloZRSlz/Ma
7d++g6Nu40ddcLsZUYUtn6M4HvBmvg3Tk79Pm5Lh2o10bhHGP0wyavbyanhlULcrEfydGMFoc9nz
e/yNBhwiAgdEABMd2jQw07KUl8+m2gN4Y2J8IzXI6+fg7J/mRbPM+4LDQ3TnAUi45loD12vznxIl
foAd6eObLOxfKE1Smp/7BGu00LIaqFHk9VhieWJYaH4x615+UE2Tm1wuXOadC0VXpVA5UdbInqBS
la+SpA12Xv0nHb7S6AWBMbcY66cxYYqKXyyhgF885SbkIDulGZYZAVSvoKkEluYrz+U6PTRqWEp4
hfiFVhKfJXP2hYhQEjp+h6UhlywscIgOmrKWHVdaeEVPVGLsrOrhqVt/kPBvkSAmO7HTIXC64foW
21uXcPLdNq/Ph9h8bgTUWMEoCvZVcINndMGdNWJcWtSaYfMVX22hEwmTouCgFRNzYCKv775Vc/D6
WGMQ4UXjaUbYghaiXsSTa5Yl2NtT5mNWugWS5fvUV713lQuiU8TRYfiQCiTT1bzukFemuAr7VM8x
uHM9+7PlCkY/wN2nVP/tG8RI21x9v3ZhW1TIYq9m4jf+xiGuH32NB+XKjb9BZhE6g1Z07t7tI6ow
E5tRZh6g+pfk2B/foYvMhXfwAtM8Av6fYyfsZO3poUON276j9SUojKw88ThPi0IbpN2KSUYD3KiA
XoOHaZl4yF66w/RhKMpNO75dljpo5r5tyIR8nWyHL3LWJ2KHeCly9O58xhkezE8VhKJy64Pu3bGx
zVk11hJrqEdSjPJzXHh5jUCWw5Ra+8mXlSBU5W2iz0QDpSMrsE7zZhdHsV0RTVB/nLKN3LMfqBOR
Ezyb0vTvYUWUNlc6Efk182bnisiKu/WmPK5JQ8F4d5+z30Wg/WrHPhoY6cDWKsOrnegjvNoGCDbd
iorZILw18Tpvpuyp9HuwUjOWxiUeBv4ppbPb29oHAOdRYq92fasP6kYRIgIxr3lPT0ZM71ojgstG
CAb8mcO8ZpDt38kyGcC3ZxxIFjg9+fyHvE0FI+1aXlZ6bXy7K9Z4Syi24NfbbLLmU6N+gjvvKolH
5xacu5slKlPualq66wT0V127NxolxbBxyi9hlLONYQrCD1xzDrHtYVlnCIHGh+Bma0vFQz6E9ZM+
EACrSwOtLFN2GFZqbrptBYz/VV8zERtLm3vrJqa5XqNK0redE3PtUbMNorvppnFEA1fqof/rOdDr
UG02sAi3IVfveOaM8AlXbhHbQGljL5ATMIj2oNwe7EEc0xzTLpwDyxqjd6Dv7M98ffHX93vl3Grh
TpRBaO5hSGFqDhafDVpSgwNBUDnLb4KshBpA1Z50Kq+ZRQ8U4qbUbNLHv86kZWjDpZ7EkLuquqtm
zkxr6j2p1s1VLJN9/nL0XAkYG5CzKJbdvCr1QfS/HlujMnFJxS6hyp6R3kzjBIhHKVEPaZPIn0XY
HkIeWdF0eWmE0iF2EPipaLwSv2EvX6bvkmzkUPP41pTZ+gCgz68cIFk9D0mK4iv0ghtsrqyQwjZI
yI+aGRZGY0Rju/uPYy3Mu6TQy1oulKuo4ooQDGsKVhnZz/4vau2+8U2BR4l6Lwbn6M5b/OuIMYHU
utkQktikRx+npFos8ORveMuFWAHnA4nWfdF+gjkTIMJzRuD1Jd2Vg+MVjXcGGhhK26GiH5F8YZ++
o2bNRMIwt1V7dUuMXg/RMtNjswQeAUSR32pxICYd0k3wOpHVWTyw6jKnWSKxoSGUl6VKsgIGp4C/
0R0lZoN9CVB3yEZd1TaCH1134QAGq07TVdogLZgxKx5KgMx+kyE0WfJO/ttNUGvvfJnfk1FdQtBn
O3YhnMnSdVqGrEvtEDqvPlKZZohxf4RoJ8kJtrvYpCt6FwAmZxgYXcAEK6DJ8pFSagrcnKDV5nkc
DGTCBprohO/BQm+WR/Drmwpol7MzjH2I6aSE3W0pIeONTZWz/odCrLnfkCKFRWuMK5PdwleE9e0c
t98txawXUpj1oElqanbHcQAYrFHLWrBzKoqdyW3p2uWVoexi70FhiMyYFHgNco4hR5No6BHlek3l
li/hm0jbn7N1oH/kIs256tBPSB1rQTY6ommqrwMC2aVKLUMMzgDIgjmWjZwEtSRUaWsQTDt2JvfD
b1nunEiW7DhFmYgJVteaU13xund67K/GCdnQz5qePULRp2nO2IEz9oCvL0CVj/UvlF2r6IkGze+J
tIuX6LviSXbjDq1ezbiRO0Da382tUxrBcz0dQfBe2SiXWz+SCT6K4CVye9lXve07kI4oz95qBo7S
Qvag8QoU/WzIEhfA8/L8flhpO4b88gZgNBxkhHVtlVFe2RFDWP+Px/pgx+SiAU35AmLzojPLxYx1
OJTwLavewUl3iY9S2RAdcphjAJEz533bNQHxMKcQYgLbT8c4PEEGoesHxKV9qVXAV7cK+T0kzKZY
TQ2D/QKBI/1hsOrmQ8uC+npcP6jForEEjoRnSBOwS2l7g2XWMtrpncBotYM3JdBtRHKtFRrC9DxG
0lU1BNc9YOP8Nd8KDiT3IIH+HxrAJ1HR/rLLXFA6Au+qiHz4Y5edCvPLVptbwrRQ+zN+TpsuIAE6
Qijpuwtw9MYrQReV3bYSmXheQov2G3VmWq/c1cQtpEfnkxed4T16rWAkzFQIoQchNp/4uOuFTM0O
z9OsfLW+JNFC3hl5m7DItzAjAdTuRiFrKf739Luxadech503AlOia/r5JbnhiEEDp6YWGlfaCfeu
QeItwvep7kcrUPYVzzaIFT5Eq5Nk6cnpCHsmFTD3t4lqd8rV8zi4doZ1TJdX1GrA9W58ng5gq/be
CfoaPrJ8gohO03Zh8Ir9/WfcYs5pWU4HkLG+yPg8X6KBu/Fi4v6fgugIZ/ApVxasheewvaF5MSrE
4dMQOV53GN+hqci1GyG3K//S65aCQKaPI0mRn+9fWvKeOJxgBCU3BjHIz2jd+AaAREXzsRg+ekvf
/xOCGda1NyoO3BSyJ7gu+m04ha9WHLzr0NXKi6oVIRWuthyhyPdXM2nD7P+O9n1NVbQzBuxXR6XM
lM5DWkAlWKVGitsFCe07bxPrnJ3ACM7VS9F6k2MHaRg1bVI4oXvM7PPzn49uEOLleos69vR+9Plx
YFC6iDYcpZHuOp20vcWH0oChP5kw8FggK7paYuC6Oupq822U6x55/Qkdu/ul9xR/6RJcpdw9OB9z
rp9+Ae/LZZSdzfho1CzJd1htXVr3Yv5q+jP4AKdK9JAHyDXzZmqe4uGcZmKfB2yWemNSe2fZeplT
YQ2OUgBEy8S/nP1pTzIfcrhpDiAghX6HjZUU6Vzg+HKYnpwHB+coBcE/Ek0TcRQV9p7TCXMh92Dv
Sdyz+Lo0dJfqaTmhAHw3F6tNMagtpVFdA44h75y3aneXheEXo7kbtwiwNwpVHxrS2lni85+HazSX
LEcqDAmybMBzMx7iJB6PPsJrfE/R8auqVEG5rwaoIgiDx9R2qEHZenTSL85Zo/obgGnCxMxLfgKZ
QDl9coc7uQQ9sJTFnHu/2mq30FKEerL+15X7nHQrEfxv0IuFj/FomaKiD9p79TcGJ1kMjOuYozjz
v4iBOKhlav0yJUUsV12HmEi1eeB6NzRti7Kasx0rOObN/gUhGyIAC66pw1jvpRHRx6N8Lcb5B0w6
ALPZ7WJCxrJfPLPyVyNAhy893L33jv5wmXT4L5f2IZpCGOZJQb9X3ie1bBEBJ2sZPetTi6MXPi4k
tbouRcHwgwKMtoPclnctfBPn8RmiLYdMQ0/JSWe0IKuWqY7CxjrByoYrr6mQy7IixLYAGFRzeQKc
/an4q0oJhxMaowZhFDmduBO5jY+jHpI3bHlKTM7xffxOyV2a8qvnYODOuIBM0jGUc2Sz3jtkPlW8
gMb5FR2NbWooUktAEQschy65fex5gD035lz2FZ5SIBlz5Jsl3W9uyPQveBVtoLbaySBFE8alCupY
rSZ0V1aqHQQGyo5ZvRVuQOvCBHCQzZ1ZNDqrQMC98xjZ9ACHNlZsjhLRlmA5baU0DzxCfQ/iiXKo
IXRSxmx1/OKolT/NPJQo9AJQGWhtmI9+sZ78dEwi4wrHeXheIasYhf/PGMR/1+0E88d0xdJESTBo
0y3poaWkLgnSdxehRHATuWbElWrQ0GypKrr0aHpP74t0neS8rAtBTCuLtokbPh9UQH6YumoMGNUh
Z9rzZlxE0cNoVUJb/1scjo7DSD1MFU4aOogUn5+ic2ciBEN0din2vlIuK5QfZcOVAM5c+UkFr1ou
aolzEaSBsn+91ASokgSAdb0JTeLQ+iIKMuzT0kQckDlmzU3w02DnOiVz4X+bgjmMOwQC+4uTHtTl
gAXjSHgyQgQNxIeayaPEy4IoqH9Ujb3e/NE8qDVyskcAe7et4LGzdTLrAMP/Q5YATTIw1pU5KDCs
C7ceNoAgui1q02LPWZQWWzSKdtcT+YB/7uDF8CWj1Ks3EBXJlHaxxcKscdOlvtTP/ZHFXGf6uCrB
vO8mcwrITkx5A7OvqFRX+KhYQAkF1AczziMIaTSOE5s9sUjGxpZeoBRb4OlylRKcYd8LJuSpRETe
DP4qAp01CVpPucCdGxxNOvqRuaBTecufPfHsGdRSA7T3UcN4LW2EgYvAbZSCowthrGaSnkFOKF0y
3Ua5r7vJJYAdgLm3K+tU7LP6RjhtCys+qMq3Ikexk3G7r/2YanP+GFrYManS4L/8HhXepmCobRQL
oqW4vtObb8n/pZ/8WSVtvaaFD9Ynn6NFHLEgZ39utjII2B3pc5SxiZp7MR5S4JRIcz2gJqr0a0/y
WpLJQM+isIIbx0/Xgy+I615JRJyEtV7GKmuZ+7CpgWGw2CaVsaTmBRpnqsmqnZIWNLIGalYPEfG7
AfhfYOvqsS5vBLjkzwWjFpArFpInTnTJj/s2GATVN0bGqjw0jp7buq/8NCwsgoDwmhaErV/CW8ra
npYxBeMjwDS4bPkGuzCy+QmRkEP0QWRbRcOAiI4Ge/uAVmpch6vWVQBjS+bKWPx6tGHUsfBSpuBL
hnsMwNZLh6J5sOIXPFV4mp7dMbBCCKIDnyH2HJB1ve3kjK19pknWqSeEcbvw1aJui93i9Tmljj0K
uVnGItbrh3P1s7OraQCGWKynaOsAi1XdJjQade51uRxPe9vP5gkpm5peDUs95JTB+atk9kNlHl99
Mv/ok6uRRyQwcTYDTh6xYudy741mpdVB/uCZ/9u92qm28/wHDPVK6mcSyqkeD3f4kXfWjZKdILhH
/uEGxaMUdx7u6zYQNtB+UwK7U1+hmuhQXwLN8gmMBsIl7RFPA7jC4jAAFKlkDFmNKzaTovyAQE0w
LoxQD6fnwteC6y7CESL2qANKY3J9cGd7RxKH2L+xCTyDVfMkf5ayAnQsaK0gwyaJUJb8nivU09Gp
QwC6Tv6rRSjwdqUAKVIlAugiuLHbtQYu0dB6FQ/8n8tsaVkRvItS/XvG4Hq5xEO/J0ncXTIjL66L
DSEnWmyIiS2r65x3l9QrnlOjTuxFRLWOoQPbCLAPfc7pMfgczl/VZr+uvjUqcNPnaT2UBKVEt8GJ
8zBQSdALOP/BDUpijKNdeh/9bluAPc1ouDirYfGt0ixxCdS56LurjEMQbpCc6a1+M8Jxqd3ifSVh
PaiRuC+UKGtaptBCbwaKADK9vy0w061pf7MyXqq1PkICvYBpbH16HqNE1AZoxQ7hyR8UCjfyULfw
LDyN/lUh/qOLJ2PEwec173txOwF+vbz8knV6KvLsUVzIhCrMnJEuu3IoTKuvtaosl2Y3cjpf2p5a
at6idWWUrmlByymyx3XPeuaL7Y7h4JXi6nNi1c+2Qd4HuNjDeM7W0fgjM9EBYmmTui5wupgHnUj/
kZGrinCeexQmiNob3nmFG4QTqaWhPUpDXKkP7kQyrrGdfIST2kRh7shtuJldElVqFwJ/bUcMe0vj
taGbyrkB9VOAep/391QTeCiThUL2Q1itumBWHtHKWANoQDCLy4yv8ze3bLj35HBXZ1989sD1VzKe
p1V9ss1q/LB2Qn7KqKRdWEXWHlEgdepRSb97rvsuFa8hkP8UCrQJEOgfBFoasGx4aU7RS/28x4eq
cgc3YImvMn627jVFcuXej9SaoLXwX6Y5eihySsECjZ+x2mZspZuAAGCkJTh4Xc81sxpM5rJs/OpU
fRlA9DKcx4fYf0RyiFJWvR8qzlwZvmiLVexga4XganWIoNAUc7Q9fptG4tVRUZfb71zDyJ7aFZF6
FifmaNZZPr//11ovjeYwKaV0ceX5k+HbvaPJnvs0O+IQSIjoQzR2sf5yxrTwQ/zud1/VMlKaN2oN
OhMHa0u8q+1+aAHrgJOwb+CAA7ZRH0XJNHDMuiAkgeiJB6gUtgzxprp5tszaUkok5RkZ1Cwpio3Z
HhY5Ttivl+bhBgJGzhU6900UyNQPP6FIeVMvMGYR9RU6ciuEX6Xt1sMuIzP17hIjiOyxB2jnJP0u
mqsC013h/+lq4STI8L/nJJW+frzcyrzEMuzV2jr/Jlc5lA8zK0ZDb2tCCU+rkXXxFnvyAhisEwlg
7cCdPpz9UzM61HzY08VPKwWb889zq9VJA4pTf9v3yzLQ4lYpmqcYB2HKhKp2gOwVh73ozMmUrQ+L
7mRqY0oblumM8G2A0ueNVIamf5hr4i0RVdC98wIwAi4ccb257OVsO5rKPQ5UYc5YEIEG9twAsrf/
WzjJIbEAFLAkZlvPAMuqaOV6Ea/f4VqBte27Y0T/3USTU9CcGtV5aCsq+yoD9davDmw6jBCJLx54
Y/tWYdZODEA3BkjEx/6MPDXMAOkyctu2hhl3gFY9onQGzwn88dZsue9XvBdOf5dvV3E/pKct/SbK
IYHRASakKeoVPUQ+yBPXbDrIYdFuO/CDOrZDy/hZsMklrGUwE0C6bk0rxmb8aE1lkOr3B80bu/mb
+/TgxUe0QtciEQFWo1RFujmezR3vdzAuJkbqJnWsgIHjoTExL50cYpw4K5biD50agU5cvbRaDLpj
Tu2mCvbe/n6afKTGh5ILMs3l6DC6/budnCAOBLeb5qJ4bBggIZh9g//3P9stKtEuOPwDRzO6mfMI
BSfQBTB8g1oGz7nzXbrYJ15Wd5GR4JTyGTOw7GerMqr449pCONX0Kjpg/ZmLKE1Uv/xnGd5s279R
5AeVdauFqmubsPY8k1+zLKDTeuYDYOqev57soq/Z6ILWgIkUjx4V01HZ4Bc0UiskBOWV8a/oxJ7f
b9vS4SRhErhIBayXheV4CFmn5w1fxsQ1+W8jlAngpd3gSGFXIoWw2S2puQ7+4UVm+HoNt7XqCyUd
MqZaZbHZp5iqhP2zl1HydIu0VcCFPUDnFZPM8xz6/4Ue7Q12qa674VoSdjUbv6/eFF019xPY+X93
ij8ibMacaBX1JAYUI9B/l/hC5f/WjcB6RSqDr0uPSk8ZfoIeKDMiuxZ0MDJ7s0S7a9XHQtbR5vip
ntZZKjFDgLAOjHQTHVKi/NUq+Xke7bzXqMF+hNaVzJNYgfqbjaZgnH+7knmm4luTdHEabjV+jioB
M+H2+eUCqA4OsLzqyXdzzVBDqaTlpO2NxfYGEmxcj3KyxNbUr4xb58iAD0gv6WLL3shYlu1l7Rri
jJBpEtz69noUC8Jkea2QGeZndk7jMC9v7gx9UBSflqF0yBsEtFz+f7CdyK1fpphUV6wPfztoibu+
VWCKFTN/A9zy9RrGIwFa84TqQ4KEq3l8kKtDo2P2WnbfZVpesCZ3n7UQiAEIPvCbB+TK5gRF9hYb
j6hInbC4M3hWHX1OK8eTc76lCuNCw+JTy+KNmHA4KBbYrZ6CA6GOBOGHiJKaNUbJtxvB7lFXWAuM
bxIDkxpO4g2VFswGsZJRCvyrUwpUNVV8HDpU6E/fzsFcslL0DoRUxyj7DrSZJ7O2FXtdlPCPcnAf
wFtPjJI2BRXB6d9sPwoXNKbmlAdnlGG0fnLdmBmcJWOMDbG9jTFt4AA8GLewHMqNinl1bAbizE3Z
qjyE3Q0K/XvDnsN5RLBdMsqhSVQipnOIjmi32+A1QgIBgli64WMiV2T0/2K7hjQFmT7dcR88MIwc
p9EaaJQKPK/2MgKpAyi455Ux5JEDazvKTok+uaC3rD+1GfAqDgfK5yUVjX97xojs6P25uR6alFdu
Pt3qHy+7zRsF3GW5v786QCgtc/sh8GOKtDnMoN61hY2TE60JdkzATBIa3hTX2i+KEkhQjGqM4Uo6
QFDVEbwYvNeR32GWY79VpEu4ietqaDPz/3F+Edl0nEcIH61J1na8FoFfZsydZaVrbvHudU2obFNJ
O5kPA/c82APMORkGTMfnA5MHD0C6+/WV+LKudVxD85IJhlXYo/uxPV9jP3QVXYphfBPzu/+Rxstr
hqN7TKS8s8BE0UCC1GSMlomNZcyWXqiYzNUjUPwERK9uN8svLHAStLO3thWjY4Hk8ACAIo01SUwk
FL1jr6qWwLTBq+szMIaglCinw0dLF27zLjz538GtwqbJ6Gj/gIgG4Ode4LeGj5enEqfBeC86OfcS
cfEgZi7Srp/ApMurCguipkdXbJ5xXWOvp9Z+lHXfxfFjHTWbDinuY4HUwelJ3Hu1l6cq8SltCbTo
zoU/SDUcbtqxNeA4NdBFLm5LYdyGpYrMQ7IV9lpZxrJT6nYYyV4MOB6CYyzsaiQfZM1tmFI9Ej62
LtieTvpwTU+SMQjcj7NdUBDh7go8c2N5RdYehvg0Fn8Pyd1x9PSIMibgbkPk3CJ1hEWG8bZIb8j4
r2sck/Hh7eQAKgab6vzAQ1vSsUN8tOCUZYZQqMBf+Ys80SwIg9Htx68vtdS99gEg6kK/p6sgHlNY
ZXGXw6ftJfchTS3T2eb7psr3vAGFC8HwP+HHpA8TFqlG4G/30WTAi1V2Jpmd1vHoTf7dgTiCYzOR
P9QZfOD7i/E2KBK9tG2V5LstQmf+lQyzGiJk4x6ixxf8WfKIzL1qWm8f/QjAHNJkvHCbFG1y0cLC
/ClbfhhlOBPf1XHItDe4BTCFjgL6hE7o/S7WW/32UQu9i+I75a8omlhrhG1nQyAKEonfvbJntcT8
c8xN0p6WuxcH4UwLusbSyRFpBrhPL3lw+4eogN+FoUQ42Ba6km/+gTjhThOCRR4B2v0nSJ20OflI
vJcTrXjBTk80/9bCiIV9lJEOQihz5aqsnojFDcki6dAdEaKsTX0EzAMluJ2sjYj2vXPSAgdtlWyV
7IWvN4JZcgBpQ2pcav16LdzFleWeeqqzR4J/Nepxm1L+HxPNZhQT/fPH303holkqs8hfFUMoabWb
YHmHPa1RZ5zWj0iqzm/ZtSQtIldk1j34OLhAFrLIzJZ24P4bbP0bsUVUsCx/rTLe5gjtI17FgbaW
MQJkSgtbIBzFGzmLG3zypQe/5Gc/MxxapVdJyjct922uwRbkLJUk4AWSOt6sKDuisyMLPd/BKL3I
YgE457YSyUFpn5iGLG3HWt/HNak2ft6W02L41Z2oazcPL7EXIy9q8O+P/R12QpHc+uS3DcNbfsp1
ETShnAnkJUtGwpxRcUGi0fupR+bfB+hIUKI3oomHCovm00lW5B0qH0GngU9OA/9Nd3dz5pFSOH+e
Qj24wMHbLaRBrI+3GKfk10ioDhutQ1Rxhc0oYRQ3C57QmHFr0xiiaBANhI00qK6tV2i8KnTwFdue
xTZNrvjDirENJZqRiY09xaLSwNXStjyOSlW/DtbBXy/Sj37/GpOyK/0VRr1WfAkg5iQxIUWIrRoC
NcQfGtHl7ItJ1Mw78mBKmf9Uihk7nlJxNGZj9evYj0x+hb2hGED/RRl+Mpjvlv9bliLe1MsXZAyn
9MfcRKDZL/Lnkx/C5c7kcdXOaUYFwGGH32U9I/n+QPXcelDAYFEHV8+qCYbwSkrijuSgzfsBplzb
tEaFm4Y21erHUqA5ELKsCerubUooAQ7RFtCUsQAWFdssuupmJnBjAXPKGpB4pxHhLY7kwzpdLbI/
w5/eMv+nSW6rNTMeIwS/K0xrdvaswQ7u5LjZdUJ7T6zwswIpGuqytGmCgBd6oRGetwuF2C8VrdEy
LE04ddSYph4gx/7u8JIASV0SPeXrIpKVPMnXlgJmtAjie7cxk1QFHBbcQtZpZfoK524YG3wRY9nZ
6JhAqSzP3rZM4emlmMOwkMRu1eDPTWgrRQlk4oXmJ/f4JrBtxlZIWQYKmuFmjp2UwM5obo4A2Yq4
2azj7MEZA3u4shFCM1Ff/gXCOfl3qiVWkZHbgrodd6Q6hZ/a/R8nzgxAIXy4FMpZaiapynE6OcD3
/rR0wkSQrRV5hpkrdXIDu/ltRJza0UE9MajkJt+A+6nkNeWyHzn+j5UgNSJTAZSE2xNhYCb22IWw
4FlMZld9Pi4/vAjNL8dXTWj+hjnVDsT+yGpFLMkcNZFokrMSBTQ2czvqZs4TyFLaj1PAjbZX6wKb
58ng0JrJYwt6sAotl8xWk+vMRnBQvjZuVMNAdlejP6bqJ6/YcVmnHuwEEFqKZ1j6CenCMUPSAdmN
QBJLFdSlopVKK0GDrJ/jXUh+xtXRXLCzGjpzHVaQHGQEN+WlLr6YD+6ANRYdf2mp7LmvnMeAly7a
kzdcvyt0w7WqhwljFp7U+2E/xrvE5B/A8J6FACScOLX0tZHDmZyUCKlpqEXZcvsK4DX1SNGFx3YJ
j8wHOAjibGc8ziOqY906zMCyVxFu9fDItfZg5dEnZXEV8WJ0FbnIuR4Devp15HjxRIisCdUyza1Q
1FtH/ygJgHiLoXcyluJGKBU4sTHF1ciGMl5HHMlxyo+kOQx/1LUXbzDD0x74AV3gIeNabyOba2OV
umaxisVWOkWEuy3gy7iXNdb1CyVoI7qqyD2zUhiUqLJev5YqQJeDxdODKJMuHeUb2LF/rsIUUL4y
k/z3zGdLtiZCLHtY9NqsWJ/SWKMVMsyKyRPEstDD6URn3F+p0nXEz3xXixA2SauiMAhraGffamxj
BnTezjxnLjJH/NuiQ0bo9u7x+2Otx6XAT4tUpACljaPbdVSO357fIaKP4OSt5HX6/WBtdEePB5w+
dcXUqJl7a+ouBC9ACYO7hWoChTt43xFp0Xh5lBIbuJ8y618nuy52fvgD1cey0qlkABQhfZbLbhzo
JLZ0b9sjz9FrFq/1Vj5+4tK7o44Dd2NKgGmNnLvpY1p8R2uEnQhOpz4havgdCSPW8HwvmvzM9i9Z
oKq+5ce8kDD4sc6lvGbFzlPLfE1tLvFA0xMU8RVOa74xpvLNqQatvyjHrqYyekBjLj+ah2KCTahC
pQ2MNFHfwL1N2369dYKAFZLnl8SrzewyQ1e+oChRSi1hNW1GSO1IGUFfPx2ypuAi/5QpcW4LBk1S
hmntIuPBn8eXi+90j8hlfmJ7iF0dH5PIu/s93xabLl4uo7h3kkLQ3rm40VTEZK8F+7CFG4qkKdZJ
YynNv5w4VGmQfQ+fz2CkPAGULWFH9cp59lymBc6diEt7ZncsaGNLw+yESbRuo7zoTbXwXYuN8kRl
M/5zfDvx1wkhiW8tq507WBy6nNwYyLteCtpqpm75lxjyLENynNaK1n9bCN9byIEshq9Z0mc4hno1
PWTKaHYwnvx/kNOP0RYQNKSP2wbeqeVE4UbywbJnP8FG6jjwyoaR7Tz2qKWvWtlC7EEm5qbbnKrj
boRnhXImA1jI5byb6Fz9vtl4SCNJwCtazxYPq7a5Q4nVLiRKsvq4T2BZCNoZWp0PCcJATY4+gsYI
G7jnPhXIxNpM3aJGw8+gq304IakYjbThuhSNqWgA1OIQcP3FtaWMmogKF89V5AR5Aqs3JPFA1cnn
TL6LXHG3a0i3bF6z4fZ5s2x1MbQGPhJbenwFKpk9faH/vhxMjqWlMYAf0X24Qyd9ux7PdxxIhzm1
kGchzRjfZ/RvtDYMXGQ2D0SI2PpAG9QxDIFIzIkc99OoK6/fejjfJDPt653xALhzWLUz4iQ3phos
dW3bUxnhUH39ZLcrY/lPZ487+BIDK4L8PaZ6ZOw18qYwjMvxtYwujHhkWJ0cGAvRt8TrM3dCC12Q
HZDF5HDZ5lV0JJuzcwzM9QwGGFUbRgi3VEi9b74oNFcdAFgIAQD3zdd9uRpcbqoyhbtWnWxK6bKR
zmD3ZTuaGPfyCBp1eGVC3wsU65NNskiK17kfYBx1zwLc2tMquiO3DtpvVWcJJO2NDmbAGsKJ3IIq
lzNEJv6QQyslPyaKOX9p84Id3D9g0it2FM+1OAcEyGh6+KLVQSquL+lVfG+tvidDnF8kpBuFMUaI
ebmWC8P/+CGTb4binMsAfhQ/KXUdGMXsANMdq2cOOKWhSNZHlEBAtKE7u14ULdQVLX5xa63mN54K
985/wxMv+pjgrwVMxi55PhiBD7gvqQ/mvOH0OHzvZUq9aOlemXBD6mfBFKpbVREN/15zMxhPzmRy
dnfbQRQmtTVQi9PRWI00CgLKptKttzzZZ8tkXeYbBr6+l+lY/0s0aA7DDB9xdio1iMKaiFbOZwNu
Iu8bepwgES1uDXLH3E0+KW9ekO5vTcJU0kX/Hxalba59TnC88Z90PfNKc9K7D/eYx3j0cyyPCHqm
MdBwjz/ji4B48IbYk42GFDRApkPbE4iO2Ar9ViJvCkg+d7NT8w5VgitLSrYjuk3Oc8ErvSe8ytWx
5U8v322dEZyrfEPfbnJmzRMqhC4CU3k9X6wKhZBFUEHJ+bGqeXNKvBxfV3dwGiAh5RJobwGo4lAP
WApjv5VPI0oJli9aoazFUtiZ8wjs57mPxBYEKO0omln0mVB2K5/hqZjgC00SvJ+1KVdc+P/sseIp
YTkWa4/vFGrem18f4LjI9pkq48nj8Pf9FA7/JRWbfEADMlHtYf2x8lpMPojhyzlW68YWAOOREEGG
Qd18cwi6eelAtjTR1+qZdZpdtkk7bA4T2NJuYJClW9nEPTXv8JL7ZW7HjUsjU/clh2pZs4QvRk/P
MC9oV5AyZaC+id5gpo25d4hngugG9GjDYVPfSJMAdUjxGZdYE9+ZPjmd7uJRmMevTP4QXTgIvhjC
5yPA21Whi9ozI8ey0DTSTIzSGY2IrZCeJehpG1A1jHn3htq5YXNCyqN3e9VbGJR6UIcJTlY/vQSJ
pIfKZ67ju4MJ7xyaz6QMBMFV9ftdvzuOI+B9Wnn26xnG6JZY61aWRx2vV/789FXbAl/FMgGK0cnR
Lri/Km0tbg3bLnrilj9kYVHQnxoHfDbSBYGOCyCELMI0to/xPfVxTAHx8UxKdkegANxFtWu/IfII
B6bs6TdHfrRxzY22bUc0r/ocYcuy+0AhryJHKgY7WGw7/2QoX+0ClNwCBwrKdDfj3gXWvtQ+xQn/
CVr+FYLnReVROjIs/c0W/DZQcZoKTStZwQoI3eCCs6ybNDULdhMMV9TrVFm9BYIDpQUJF1Eki1EP
EqRYhR315yZbtqK3NDBeF7jNWeCRvQZNbwcZagE9PXONyyc7dZ8hY955WYQtZknWRP5Yn0/3Apfx
xD7gZuTzUVk8Y0lYg/rUNJGfnKBn+FGpLytIgR5u7TzGHcs1gfrI8lt8YwcnKkiuP+5V3guMxnr2
pmm4CoiLEgAyEQPjhx/EjbmIohVueY1KRk9D9je3LMM9njPmZNK6v224yr1StPPQxSVY2j9Py7of
UfU2YRpgKW5LeyLzW0Fa46iJUi/xF8WMoguzMGPJBVo/zl8bHTfVt10+869/yjkkKFhUDJH+GE5O
WRbnVTsuo/FVmDdgARnIQorMFgaMSwKinyGRYBL71BMK2OYWbaAL5v36O+kx+1w/28xlFxahEkts
ywIyVjofSNcHSSev+AVkW1Pdr+lGAEWZq0gR0iJDqgNVJ5HjtxaDOd/JI8snWkTkwGwgeEncdN2X
wjkwASU8BjzzQ2MmeZoUJH86QpSMZb8o/WxaHMi3jQxxQus6i6P1HE3xkkSYk9l3iVTxC/y41RH4
qRWIX19mNMDhtMiXiYgXmmAhIcNJUW4X6qXxTTQ6E7lG/Sb4bOD576w55CIFhaOiy1OhT0aIbDAh
xP0+8UEm0/yVoox0Lx0eqvclnd6FeU10IoK8LRdJO/WAuexRau5UngfJvyEuxx+OkujNO/Ym6ZbJ
mG9qDjBlZ10DVlZ08/9YzTinjet/dnW9qPJgMKiUJRvY/uAtN+J8Cfd3Mr2Br7yESOXrFnbq7n1p
3OGfEzwNF2wodNhpPpgTDGYuJHszthvvEWUt9b2kGgoY09DBJBIlFZH2JApzCcJ0c1j/kofW56Lv
BE2nB2x3gipcJHr1nZtfAiwGCC5cCKXCNr3cgQW+mcGmfSXnRdbD2L7MEnreCuD24zNFlwtLnDM8
Oe4bYet5AOHbvLdCBySjzQQRHExe64VgOWBxPaNo32QwjA9ooQZLnPJnPGPbtELMk3ZaqA2HfZwd
SRAL/ONFKx+9jm4noVngLkoG+okE5dWBydU2Xdo3T1WVa7zErsDEAPLooPXcPrN5SIOuXERKSZ2t
amUW2DUk6iqz8NfJ5BHCKdb7Pt6ULVKGNLwGCdyEMr6jl/TPtGmLoWtcPDdV2UtnK/iTHxCznn8b
HVr36dT/9/UxFWIgj4akq+uqSNGaQ83hbxfLi0UWCPLwWEMwqoJ1AnlsHJ+wLfaYMoGM8kTB1aI6
BUyLdSy2yVlOu6IAxR29bF49OmfHzWLUXXNFBA3WprWkln/j5J1+UH+kzwhVWz4KGNvURlYejgNZ
m2Us3mc0EEjPl5SFW/kxnDYpN59bWO4sQwEan/H6Sax5w6XaoI06IMxOPkhFIRreGQEtJYdCqq9p
iqI89AA3ELMcJzlUiGAkjm0dYs8PRH8oR8cm8oyNJyIdu6btVg7p47m5NLkT7wd+zzH+tDhcF4hw
ysqxHiJGZpoV5qxomyY34Z0wej1Dj44GfVmntHvAfFTmn7MIaZfqh6WDwCmJ3gbRT3sjZNLVTY2x
+OkKmkG89rdodTT7//zUfALDYt8xaaTQvwzQzL9eb+SpzR63G26VlztwvuS5TFShr87me1Pi8UO/
71VBoseJC8qtsQBZfQ4PuXNM8xRvQsL8ZBduXi5YVPaOOvyMKyKUA642offS17X+l0D2Y1vnKOoV
Pezbp2Mr0+XSWO9nujqpujt8+cppNKx2l4jBMu5H4lKOkqR2zfUhOfHGi1XlQEnthGEhYvvogp2M
cpcIOlYPHELFB1dHO8R1JpnURsdgFEgEHSRHogtzUqiuKqgGMXj03tNW0+dVqZbsZofmnjEmBmuw
QjDgQ9DOEtdbmBLvI9daJsMEPN22Mh0+yEuqpwou9tYPVsGoo5TJdizfwuJjd3WeksFgZ7vyZ+Um
8XcDkAY8ZzjnxaQYyDDta8pwhTMPiOVzkdtpEAO+061F9kcC4KJF6c6QvXriargvLJD52QNZ83Ne
wsP2BQxIP6oPjlbBWgRGFNTRY04ioUUMyt1awmI9noGrbfOovG1k1rTa0tQ9EMzm/DpGMtR8bq8r
j1z9DjBu0DA+5KKlbeTT+/mTy8rAaO7ZX6DLJW7/L43KzHRpfG9zPsdQLawIuIkTtVGhcBkSnCyC
syqAkSL6I8NS5oCu3QYkYRB+Dr2YZnRqAV3unMBPeNefd6+MyQKuN3cBRVJQ6l+nrWrEdRvQEdsY
sjYBvNf8HCYu/eFvl3J+mg/jWTZwRsKUgqInT1bNSYPv1oJ8akrHYYaSb/S3kLyG7YAHSjvRavqi
YTUsFX+MCcLRFVm/sd6+jFdjIPp2GSOmkzXZgxxfhWT1RgnT5yvpZDIwMlGlbAIVzk6ygKLE/Wgz
w8AqrxPPG4T9l+JX2DXjXGs9TJsWapL1Ss+2jjgg3RpyXhOaxcCeBjyWyiWFCxBIuYHbPzLNUYbM
yvlD4GeoClcRpMeG9O4/G67tLkjWAxne0NkjpiMqOS/F08uC51Txhm+4AgVcH8rahkEXRdZKRUQr
uZM/EKlsBINCnF3RJ35N3KGfNSkRCPn9XLLzBtTMtRI3DBfj6zEE5IuC+LIwkpeftw2gINjYFCT/
a9+F2zmMM8UX+mW4UQftwlWdBWyX05gxLt0RqxP0dTxF5JJclg+THx/WoWVH9tJ1455JmaK9CuxN
d7jXI8Rj7OVlIV9j9qN4B7twALqHPlDQZmTJzMEEOzs5g3nIb78zMBh+PZr0Lwmrmz0LYkLz6L6+
/VuqShhZwRtkyiaAJbunI2jXthcxCV3IHzN8whBmwNCnEO+Hj/zMvZE3/kA9N0uaZNpr+u37yP9G
v5xzMTbGz06VZ6Ua/0v4dvG9DWvqnDZ5JUzlJEGErPUDY1Zaw0+X8EzkHLYLuxeKhiBuOd/xt/oF
Ikp6HiFKX/HUdDcu1YvjD11qwOAnHO0A/kaEnQRhppYQUXjMWAQXBQtrKxAS621mByPg1ONYGVZ3
0QwWAjLSVz3C/ScVHGJh3GhVOEe7WJDr3+O7lmiJoMRAvy0YyE1cx1uNyl3zLSZaDx2C39xx12m4
PU3/9oD+QkDbCCTfBhk+bzfFhTp/XebL6NFthDFReXX7j1s71aIaO9L19bGG5ol6NllEfgbQ2gym
q58cHDCV++jSQpa+/pMAxkH4GNA5C/hegIl2T0eZRz0Za+oH0QFwjGxetL7fFaxzFN27HpqwaoRs
aipBaFFH8fJw8miqgRBJYynLGcigWDxZVaZkJDjhmkoWgK0B71XPGj8fS5FsqdBcYgo6tOlG+m5y
njk6zytE59XQKRymQPf9kwsuCnk0tS5VbT1pp59XiyZh67debmpWdkwzni4VMByANFruQflvxz9y
P98hnZCj4p1F5vTwrnntagDEMsfkELms1Sv/t0rNOeWyLIITWT6kvMCPSp1O4q//sYcXbXFO7lYU
NTpy+iV9SnF1gntYvzmJ+htJdN1/RzPjZXRHin0QjrJHV9SE3BSmX4K7HPNlukdONJmXl6FScgOR
LlnkYxXXlDFNcthNZ7McwyTXzVXxB9oeT1uIZqXSQoDsXpr2lpUMrL43McbVqTPospCE4Ns1nJEI
AJHb5Tpg7UPmoJF0cyFrfZwJERZHEJkgEsKPA8VSczeiGMkHeb/fnnaWfMOJ4hFUcH2fHNV8Xc3+
hV1lZ1ECdpH8vol1mIgWhbJB34OytY1lcnskZuDe0qvrTS17/ginLHHQy7RL3EfTIG5z3yKq8OKz
z13UhQMw+FIsqaDG3XJI70nem9stke3/I39+XjXOV4H1Crc/DQppsF6LTDgNWms2n9lp0VReiVNS
p9Dm+JO+MlEj5qlKaGr/NaXHYS7HSanVYak+qLB2gS8UXidU4l2QD22V55nrzyR2KrpFZQ0mGWmk
qrLC9D0gqbrRIawjAdVAc9+Rgtkhe4W+ZgW98X0vkPxr1VuaVjE9KzqVmzAwvRWSu0bzFGdnEToR
gh7YOPqQ3lPl03su+JboCqV8yPy5O4IcX0AOOMuArMoM5AIqM85xZQqKYJr6iWoqXRkw3SyQLcfu
Hp1wcCNeAjSnTmEN5m2Ju5c71LcxwmRz1HJsz3HQD0lzHOUMii4v6CRblL0EofdVZJjOiK5ZlNAN
QT7UjTz52ybZ+bbuW6z5dVi/+6JUr+MoCGkGc1yYjZifsYDCP6EW2txTxhiFfvG7ty8nc8EFAJKQ
UyxGv20/iRwzNfXTEC1uZeicY/zeuors2cnnRgMhL61FStJVxxPaaBOjnD9i+DAT55IIRKh/tzPf
9TY5VP7HVo10/S2P8IpNKflgS4j3DMhiBa43A14uoKhv1fQn5hnekP6qqU7gj63tnJLPsTV/fi0N
rTbw9MhXT8YTM1lMKU8ocTbBz7Qh1dzcaaQTERapRP+p+2XVBG8iwRDX3uxYu9xwrDo1HatCgKzq
3nSC1UjbI+Jr3eQm24NlPar4qokklCLNmlNoKe0QXAnGpH5RJOG/Lhzt5xPv9mVfRGsJwc1+6UZ6
jqQzNywl0Ad76ooCo7m7TBq6kIDRLyfdg/b7rGWEj7ruVbVcvuo9q1oHZXEVdXoSPlMIl/MzgIKw
MNlP7FLE9FGAlAzaPbqU1DH1UbLBn7lNIYKt0wuSa66BGc2p9A6JBpNnp92KTCL/rtbBfermXoyN
JuFa675gmeu/TwqNaul+H7b6woYI4waIKHjOPyaFH8jL5AmTD86qf5VYSiZ7+lHeliwLmUsElBJs
oLI9IVeN8Vjx+KVzGyXYUxobpaqumLh++jKfVmnDz7AAUTUT0pGbWU0hQEg+ToOl7dA7dJktMyVV
VeQ/60xlwSs9vfarpZ1rySXu9adrNG4ounHIKy4BSPTlVNwznMWlZv+NKZXtpfIKWnFMCnDRF3Dp
Z8tRcEz4O+ZeCCCoOVK5CyAIzzIvXVMyvg2xXY3TRPrgsXBBCX37OYqZtY03MwkTOz0cd0QGzSzV
TSns5PZ9rOheusTIYTlqkQQlOxoygOQxcS9RNhkVmhFKXbRZxxpElXGU0yf6L131BNuy615+N1Ve
oOg/EURZ+7gVVap8LL1ASWKFfqVHwyojZvWG5UvBkXmagI99uvhFmx03MdQK/LdtRi0B6qHQrb75
wZwROp87P9X1rx7A3PNChfMEJc1i1Z96yum/3tcFsoxT38QZz3OZR273GtRXJZ+iwGY4b8YFnFRg
sZJ6hkvrL8YXbpWPiSG1ZpsXMTWm2RmrZ+rmXrBYbp4FUoRZEqlRQzOjbQogzY0AALJSETLTOscY
t+Zhv6+zMf3u//m817DxFh0TMD8eZqk1UtiuGyRw15Jr5XiyaIvst+VUuJjrKxJ1ojLPMPQzAQlc
6WHkN859J0YKKEicOdwfIsHT4HR7AnejjAMbRExld6SdNn6epA2YObgbSb6tNu/BX1FhXmNoKFO9
NKHZXY7+0xopT6YquMSs5gp8T9CD2MJOOJtWUz7X8Bk1o0uysHsRrku9JryjcVpVFcFC0t7n3uEG
ejXArNEJSMGjreN21JcZRCrqj1lm2wK1PkPP3pVWmx8aYTs1eXFN56rKOjTMGPwyXHGTMfHCVK/s
4IywczPmYzY7Jsgy8uTb5Ws0OEyKVugeroMfxyK8eyIi9JMWL1GYXId55avcoOL/ojv15P1gn8E0
VnVv8TzEq5jH/2LyyoyyDcVcehrWqRWLXmQovGcj28KSiyGYBcPTSVP0U3vMNON/CDsu55bKAVLj
Dt+BLopSaqPFL8xdUwOABipniBHuMuIBnbYW0t4qbyBZ+OKs1N6mJRfLemlgsTPgOEzzq38yo1Mn
1F+aienSKe6AF8BycSESa+iFhpTI2ZpV9QQUw0bA4iJzUqNLJlMfHlaUQwJlnhSRnzYfXmu11/te
mpFO+injf21suaS9Z1UBP9hwLp0z//O2/tZhgdTXwSPyJcVcHeXWRprQUKoSVx47z01SVBbrrZVD
EsCcIlKUEsd4hBFKSRX8D+Us4f4VWHZtHJ4QI+pXLiJGvA637eTnk7uHZkGE4pFjnt2amQhwZZxw
5w9XSCWqnlZHCqDqALRxBYBm+bkRPr395WzaSXkhcF+aKTwvYHW2bP7xBvQgTYBITOICK5Vhv6k6
Cfougwu8VU3ttXmDDx8Eu6aNvFLjfYe9j4Az8mDEt9455hcojclajEHcpIgy9z8dIt1s8KaOqKH4
eiSRJEj+spIjj7EDQDmN5FKK1+bel3/2MfDVcsqt57IShed5o/WSvBHiNTcwLFedwsDqDgWOgH/e
2A7jZaBvCZDNrB7tBVdS1Td4/WVJqIwvfpDjzI5Y/HlnlwZmH7PtKD/wcaAczCfsBv2XGIj1msue
F3pAjNM1yGzTxfcX9qYKp25Zp1XdZD+2haO2/TX4h/crDXMnc3Sj/k5ecSCVYw9ZnxEaP3/iLNC9
2w34Y/IiGdcAtJ3f4L6kQ2z70xQHSnWY36coJASFfyGnLPUA+iEB6xiAHpZzNVw7UUG+FVK0Rccr
GfO8m0rSqdkN+LQdchXFOAmQFozFa865tQUU56+xi+m//OjqUpPgu2BUSQZQfjOQ2nhbTyOJbRjj
NHQWhPIndHPUKCbEoij25uZXwWUAjy4FGf5r6FwTDBQFMFqY8aJyjZrTtOO3o/puh+45YULnjJ5n
NFISguuVp4mgnx07bWhipjks91sSO5wQQf5L7tLA/VZ60oMYLcRjiNVPFWo2b0m1A9PDiouQiO7/
z3tIlAAtTz3CEbSrr/f+mgODRJ6u3hyfpP1IMbibNw26nza/t6uJMR+aAGEWTZl3R/pvybNkC1eR
g8K19OZelmuzREVwBvlx79kdUUBcJ4KvuLD8cPWrOARAOZwc+qBJUNU8e/zP55ycqG2QIWXnCH7S
O+K/P3kIGk8rKOBp51LOjTL7JDPS/baNy71hg3fC57nsOgVDXrLNPgJ+m6sdJDPxcuIdS4yiVjv3
/vH2ZwW2eLckyoBDreymQrHvUhgFwyMvA9jPsgCcW8yppI8bXFMZPnM6iCX9e6PGOl34dkjyfKfe
Tk/sJKP4h8sSsf1iH2QBv9wPonWNk0VJFuLR3kZE9o1JqJru9CdhcgHsal8k2Mxof+DQse6T9gaz
bt6oEKW9tqkLTVrJYcIVVw+6OnuOvHUqhrvhapvMOk/9n/tPzJMSzHCqil+C2f0M3ITtqr2qvDM3
qQKL6e/gA0J1XdWShx6QAWwy+fEK6CAyumRKyDF1lawSsE7ej+BbkBZbILoldW8qRrEgAxaQiCQT
YdE+2+wuehG8c/hRSXrcFADEENGYf2SrEIMqvxSQAV5DApp4DEOEYLtg92R8jCNcUeshicqFC4D+
GXeOpVRa7AdB3Y0H+MhGoLYPlISH0ToGpeuKhDHJn/v1EGEiPHg40zn/QhbiUHwfsQvcFNFPEWAq
uIVZjTe0kOsnOBhmGqnGI3ghyRSUU9e01Kq6yg2MQ1QkI9iptkOn5h+pyTuMuQiZBBnr1aRlZaAp
kfL9vBaIoSSKJen4W9/UAUb6wxX0ewpHAFwmWCPgXjdhg4Po8HSOTW4fgig1tqaw64dViKUb055T
nAkuBPOnXsPfoe7yc3F/MhVIzP2cOGg2ox9jD8ClQ8aGbBZf6lTKcOlAyEYrpVaqfYIzFjBGeyX4
kZd/Mk3Dde/AKBsbpwfSRkkaiWP7/teca8ds3wKld7v4XdAVX45102USgm7NnEMREvvVuyTn6vuA
4PaDjZK/4UQFWm3k0mpZnKzSf4awNz8acp5/nDwgQGu/mLnHsfFkGVzRHMuMinCbzM1YbD3nEBXL
CBtwPs78t5S52UcoqOikMUPFvu2PqkJ+ojaB3zH9nEN5NECL+uHsPQZ1/jjm44/IvQIqHYvtG8cn
Qam5hHeRQJY0J26ZW9WRdeHflJnV9QcJmoy3eQW0OBazKkIPItK4Hwfn/PGBJ/569MfCPKVHjueD
Juq9QW6ZYckkEqAfF1p5p/F5izSaYohWSwzpk5ETI47mKEytT7IlV1GVq3Eo1VRShJVwzDAGwxsH
QNcBx8TJy7vzHTJKH85gBFe7nlcA8+OoQsJ9pScYrmCD0ELDrnSwN+aDNV7PZKcOZ3AQic+qo4BQ
5YO5IuVqq5KocxmWDCMakCTJ3foti+xSyxx3qbf2gQ7FptaDnt8ImLWI/5OFXcmdY2tMREQxUho9
oCssZTg+e8CNuLlvx4aCspx/eSJBMk6CYTGYdQhbhy3A5aafl4LXzqE2KWB/Sd944NSqemMCm56M
aNn5QzNsOnYO9RsW2ubMjJdh54q2wTEIudlt2OLakkYu54vjWcISqHBAguK2NYiSeucbBy46tLBP
v+ReF7pw3NDb0p/8/KvKBonRSkE+wstFGZXwZ2YPaNkqFAPiAWCFUva9yuYOoiuJdJ9bL/6eTo8k
cBUOujufvssA3vxMex8GpJZz/YEV4Ob7RaKgb8PT12fJujZbfI78HjSgr7XKeFcF90IXQs+NPdCv
iQ/PrAzggOzTbFkG+c71MBuZviFWX7E2l1RiDPcf5WlOL/kS9u12ByBQp3SPIxMy2rUi9XDwABes
jSmf0ORtFLS1oKfRKQV7AQ9Tf7eQigqj0ioVquzrNWvOOTet10LJzc39YA9m1y/iaUj82iOqxt3p
DKMPQerL2kM3HQbSu1if9AXVYNalZATwYLVQXpz329VSnZfMXMPIG3fawEM6m9S2xmwZwI4Do7On
2YztsVXEI4HPiJ00d36efuREVUUYfw7IqxZjnwzOrH+EGTgpvR63qGSMS4WgBCCZh522FRNM9zRr
HM5wToFb5lm599WSvtNTdmmuhkolcoqOSCb2jrnDT4UNQ9KL6IgZvlXMPwMjdnjqL+WZZsOlVpW4
U2d+6yOcbkFai5j/FdYG4TM7k7LqAoi+i7foq3G+33auNg83jlYtZzbOklewmNXoJHpPhEA7YN/N
nV+yItHvl0rCBdS9vDZeSqhDDgTnwi/56A9FL+QXe8NlcEXTdfXofisdZsqKvJQO1KWmVykQjc4A
IaDOEzBENWc6/4gnUx72Gg9JvHFze95xR3ljtEeDJ2kZsA8DS6CcVRja0xDNZAK5LQykTTwMSWyq
9FBATvCC9kl3NCHp9redAgaVARZbJw1Der0FpnTMEf/72eaev0h+PdzHBVOyq/w41LKs3VE/v0r9
fqF+zRSFAFRAr545n+MCMoIEl9KHFX9Sh2OqKz7iQ8SQQhUnKmh8F3E7Fps2XXOfKy3ou4eEmGQk
nRJBhvoDXv65CxZPyaU4QKWlh5sGFSTNab+4cTwZlq+8UxXldpEmKErh0jHIftcBoWkledpoYe2f
CRtCZ5l/AYcXU88qa/axHlhpvgfPNv2S9Yu1tJ8OQ5zLjvF36DjkDprPlIT3wq34J2l8ahq/UC6Q
yCKt7AfgKsA0mcPh4HvzTaIBq6eFk8TMZYMjXkw+X4OfeDhi98uWqX3an+YY6d4WX3HnoBrrtE3v
iMZUp6qSdeKZzgP6yaZr7Tp7Am/9+0L3SdChtoohQrbAHcrL3Zl9Q5Ez2GN3rSMccy7OE92C5Hpk
XzUcsSWurGDXt7dBzxtECZ8wJR4qQiIm/o+myIQ2AAZi1QGmqYV7dhIolsF8HENjZkbYyBNrFaII
xSk6qQQPKEPRAfZmNIvs/Em2yGPq9niF5j3TbLxtGvSsJm0rcMCYYkwiuAtIilT3rBNxL0PgNQi+
v53R8Wc9Zm5rn0b7sx4smhbhMTws40xX/lOASy7gXGPjAvJnqYedECdkU++vKj0SNiN1+BwuujQA
gj+CT0punj59wpXfwzKiE7fUzV5HCOPXdyAciFyAkTU09nuJRmESYkghLLESTspm//dhcxYWWGzy
a+ELeUPtJQA+Qbw5AZiNQ14VS0zUQ5ngpQUygRvKKk4mt54svmaJXf+ZARE1JQoYO9P5x4ckq3AK
gzTKumzeLDrvPkVqYRtveH0U3W/y6mVcwtwlcx5LJ9e8kfHeSnuk3aZVZt1OlcO8m8HIaWroj4JL
b1JXptSC6tLe9iyKekFjx3M2vyxWCMsye5fvSqVCv3HywTGvCFsr21XQAVNP9m9AnFbO7cr2PksX
8bx6yPsDEqa/4FGXIH2TRAmFZOegRtQfl9b100DAOs3xDo3qyGcfJltub4arkC+eyh1hq1gxWmxo
DfilbSxtv6xsaxnrDVgCkPqoL+xPUPfAeDJeAu8KJrFC3nlJWY47QCTo7gumgF4NEStJsOguYQnQ
vXIqyJe3Px+UwI2IBvVEu3Dnp50SbB2+7nFiHaabrEUCvLX/+nb22ntHy6MFGKCNU6m6Dc0P1F66
GYeFWP6dLo7lZZgDVr1qj/HkDb67VzXqQYZJGWzGIpMo1J2B5Bojsh6mEeuxdL6wxe/hW9iWuyMa
bzywtBfrPcMTHnyi88x2d+9MO56ooXsMxvCMhTuxA5lxoIYtdcAEwTPUEMT+PxpBltwM/M8j7eCn
LJwewv/bXEYjzcWCo3qc1ReAWxmNlXCLzggNcsyvIyvW68jmfgtlc8P5eH+eAfSWEh9HwwvBsLfZ
WH6w3T5QqW6HQWuywXrpHgkvOtYWZzsVTOfmdOupllBXo9GcNZgGhYSnFVmgNnvh0wKLSF8OWhE1
u6wdFaOM3qOVB/5gDgNm2vx6MYUKKr0lC62uesH2+E7aekh0ZZeKUhreDXgsshMPvLM34zaSV/xg
6DUxaqlitMv/RRCCrBY7WvV+OQlrnXF3uhqChRNqEosdl+0a7q80azzxdUWgEfmwLUCMI3jFWtv0
W+96ozCuJgsf8swRbWXH9XODwNTQZ9KVLml2VKAX8m8IPVQhSOECYqwEbs8a7wCWEqR1BzqFi/cj
A4JDaJb8rSPAwGbdKwy+yWsyeG9yP5RrnOmDLwWSZGWmWgqnXdo4kG0w9RWZByEKgi7vb/plzDYZ
Q2WsNm66Wq/HKwKeRHJg/7I1nobYzLWZURIq4JpdSaueVG3DJ9HQP6AddPVGgdEXPxk7Ok5LDBWc
hL4mcWe4djxWqu2B9Do1lHmxrcZqeX1E6VY6mupdAkbT+EQ1QcX1DNMQReBX0JSZKoMlokNyuK5j
rWidXMIqsNr8UyFCrpvM+SlZDb2+ZVdmyyBP7235uP19Jh44JnVwyd/2GJ+FR5K0Zu8NqeKM0kNf
nOd/Dz0Tz8DJubr/H43FYSxk/eMd0heNFSofZVduNl/9ZI3J1PCEXPoze0961gyRqZarMuZQ0KhF
HSrOc+gH1/e8Ld2b9OSrVz4M13/Agy8A1QGM+D7buZxUs/+98uxnuop08h+0X3bNZFPQnlQE/evR
udrg8PBxV7YeKdSSL7UglfRP/hraIhbGTyCgSEEr6FhnkugIPMIxElmTzngO3YIEhvmwPYp3+omE
cV88KeLoz2VZQ9MmEuBKhpigLB+jvuJqUhxItGOoUbpI2I3IlePoczRYN+3oX6mzdinTzRBr4z6b
TrxxhseejGdtB8X/dwJwfTPR7Pj+lD4IpnmGT7TrvGVgs5QlPdyQsQ1JVZWXFBWvBKCBePJUQLxy
qNn8fXuPXFOAcSM89xC3zFv4bIucAnGaj/uHqlf9DPWyAy58FTVdO2Bi6BJ5X8PfO//Pq6e5ccdZ
93hzXBIzWt04lHi+Hxtyv1mVIkKdGUFfKD7u/XFQvxCeogNy1g0HFj4umZY18ngFvz+DOKRkDeen
LdUuApV6Uzn5zxLOK/xQwDaM/AnmcQKkCIp8ktW4gHR8VPtECsQjtwBZrEwLCgWiYiCxqIe16XZq
atZ7tlkwHmCoVve0TpeZbAvvNUbPhAeOuRt4UoQXkL0n7VPqzQEgw0pZZ5bqHrO0dWHMZlGaCm+h
oMSOucyBe6fk2RoKh2IZDXezK0KViBk9v+eVqH3hDSJUp+U7MjpDJr//0eZHEp5K8YozA5t01e5i
uRW7qEf6H5+FmOY7W8khvi0Cnm06k3NH4z6AJyFicO/bQpX0kbbu3KV1n4LPxfLz3TkD88KdX5wa
rzT3AzuCrsLFJKEqmNm+4whO7a6qgUAfSE99RJImr8qyo1cnA4ZqbM+zY52DZ/oPX8HMu7crTqDt
Qv4QvvlF380MtIC2TkJA+8oBNDLGP6ULzaeCy2vf+FyF75KIPIzeXCWjXXF5o17pQp1NV3CY1S0c
oevFEMT9H7gpjnbE4e58NkuNnKaQeBcbwez2b4QH8N6QdeLgeoiHvAZJ8hZ1KkAYQXiq2DXoRAAo
P40h00H6RGlZk2/om7vBewpF8V0aC0J7hTAnDFoViGSz79i91JpGumnd8aYBOxtv1lslmI4SpALc
nuaiRHZRIJWHfV47xoy8trlv+sfYHqE5kC90TP+z8jOrgQ5LjnQGSZtQd1OmLb/GxAZcV+ixdwET
WxVPM7MRClbCQTi/3mhKHG3y4qfrttt0v+wU2l+um9wJohA+cossBPm1TjM6ThoqHzfsPF6r0470
D2LH7pKqmR2MSjjyX7fDdyo26z+9SnLbC1b91+sDKh/oBolPR05fUyaCbdkyxODcY9OpoJ2J/IoL
T8cRcBataoZkMdq3H0ONqTV18XahGpzRHJhzhZv/XRpfGTWorpOd9VRRxMlDo09aSC35K00j1ICB
0nW0keFJXvhEiqGJ5DRB7TeMK4jYmGmKVJWboLtvpiHqdsnv9ttF7cVAeSOhZK705VQ0kTiPtNzj
nCE0sD0AaxjizscvuYWPQdtpYfGnpRxn2U+PcoNZ0d73ZURgkPARymkJMvAhePPB4rT95l/iOpJ6
heBcDdr4/gBGvS5B22zs042zBaKWchdnAGMT/Uo6C7to3Skt+7WBnrY/Byy+d6q5tubnj6UNNvJO
tKLAPxLwmqz1Brpc5AIY+bxRK7T4foo2zwrpL9t27cabLWcLcZNeYkdXORQKJCakNHJbft+hqauy
JQLxpiSD2CLYpWPoVthS319x7p0APEnNE7LWRlCaER8kEUPmMRJzFCIDSALBHTTzMQJPS+SyF65v
GZ7q/yNlo5d3wYmxW2PMu6Y2WH0DRa6SL4PtHyML6ilJxN5DpZ/9Cy/mM96Nz+Z1dR2iWIZTyvQD
2uONrWgc8ihcIHS36dQhXGrpaKtreUkeP024DDZYS6xFIe08FJdnbghzEM2GoB1493MrIuoxPx2Z
XSl1FhFF/anekwf7cPDls5SY9K4Fo68OiBk8309RRW9TvlZy7lrD2sZH2S3Z66wEji0uzDWLIC2x
GKigND2JqFYchYIlHtq0nFalu7PQk62koN+1xtMLD+PKJNSg9tYlCJANZ3iFUk2K/1kV8C/yWu94
UfykmOqjBTy52E2Mg8dchS4+tud1cFpt7se3ek/m/DCYhZzYGMJxWsxnCubJd01J1GL+YEkZDGC3
R0LwaS6CLlqt6ceYn/nte87dtomWDS9mOqRZcGxBNs8mh/ywf65SEG/mPvqFiqOu7PwA08PwBq34
Jpk9cBFlW3IKvbjwA4jZNYxfv0wvCz8jlq2jHHusdHxE0/V1KjH7/rXuG0cY7bOPPNovzZkUABSF
fRCnX7Umjf2Xgc/Lpj2/GGdDLGMHAgm3/CzI0QYpSB7jnKL+FQwgNIWQR8kdH551aUwVREATvgVQ
acQuk4S2T09izvwbH2vq4CqsJTMiXnmafNVVtR+7m8Vp7ZEeL5q+abTn6/9POQyKZWU7JdT1LDRc
ul6r6TyglSK9b/SVmvaHMxCAdgsP58cThk8DiW6g01YXyW/igxSCrwsEQeMuJR2d6u4GV3QULpdr
TuKMmefdFtKx0QPEiWi0Sdhh9UkQcJRgC8SJEWpY7zhlGg6/Y23rMX+olbcSOm5vcQpnCj6K5EOa
jQuCsjfqm0QA2XLwmsssnaBAzGIq5j57uKJN5QSW3qGJvPSrtUbd2Wwu+FFpbVFwYB46nabf6rQ0
Yf7FXY/Dtsc9N0tN8Dw6hXvoKXQ6GzlfkTyPdSsc2reZPkvxvY+7uAVPU0FIZELKN3KMkB1gJXRg
M944tLUk5Xu52UWOvumZEW8BeqDePoXzwky8hfayL6Zk2AMJdUcGW7NGonIOvhlocAXnkFmLLAtI
+ug3KLHg9vCbu7lnKOm2R6ZhzSqhQAMbvZ/cLISq/XckFCFVBNFlKaV7cRxOLkezb4ysU0dMKmqa
qo1FiESFKyuT6iKr9G2Zie2XHk+A1SP5u6EH/z8TfXrTiYeraj2vmoDjRUUpP59z46rEQ3LdN24p
TrwFIDGCanpQPynu4hZtQpRbRHTg24S9oWCJBB0+sWwxonUhCZRI+VrEPfqhabb67ysMT4GgIXzT
ck3BF0kV0G6yqZBWG7rrCOCNfwhhUKiEmsaWS1SoEvmtr8JEVKHlaUimSTWV0ZWCtiXHOEPRnEGr
98VGhJ9fe1TMK/tGWlEvGQHw9UzEPCkSHzsKCWP8/RUNMwBvMlEOAN2wu1FhOl61rgQiBXBWC7Dk
ugBCqo54/iBWcsLcElwiF47sbdglMZfbC+r/aUI3Yr9/ro6kbmkGeQGxmELa/kCGWcMDhvkcJzfj
YpW1ydo3KcruX1TG+9FWnNB9PqYof9C++voej63B/3JVIAIR8dQX4xz2V3dU8/A1JPGevF8B55BP
pTX4v+D0Jgh+jCFHthFHpeHkuv+s/Dm0bBDLU6hMm+zhoIc6r3FWEjo0WAnsAXcr7XEJ1QMpzSH/
dhVA6spAGORFYCXmrRhpTXd5EjGbehdXBVn2xTvnZ3uZguVvtqdPL9amQYN6mdq/jeBG71HNSOHe
iA59bY1gbD+zH+OyBMyl/z9W4zrePPQFuMv0AjL0a5fJKal8Cv2xSj0v9NbrF2ahoSpZP+n7iqYo
gc8hxuiYJXN4+d+/zx3c21+1AKNiva4fMKoocfgtCD/JDL76D9l7JxB5LZS4RnV3TuRDcUJzQh9B
p0oK185owg9qdRFYLWLBCXkKaPeS0f3SQCWqigcUk/f6IdJjEYuRIKArXVkh9yTtoqbOCtG9bQQB
uJ2CzNfDMNOEiqjX4OrKMLJ87fDYlHlc1BpN7UUeRaxglPc4jyOnAB+vJUXXGcdelccOndtINlI6
NlyetuFmIQbIwPA9OLYKXIj8I8cYuylwH73JkrQBgnHvhizhaLY/3VU0A+eEn+YiKN+FnyQBGI4d
j79XBvt/1208OMjrWu0L1F+ikEAjfevQO1ybwCVgr4E3VqZpUlyXp13qZPkPs9MQDMyeA44bKWGF
oGj1/rPpLCowqBRaAFyoaFQuXlHVZV0dzJU+Rhtd7tWGuKWKbR+zgVyjzXFCB+7p/S4XEq+kMB06
jAarL2XacbYx+EzQJORhZGAoYTxJ3qxjSrkbzZcm1P8sND2l3sqeCATiLpDPfrTUnlRGFYoZQL26
wICF31dQaPHESGORUMgpyKgs0mCH+YsNc3S+JTJUEeKGJvjovJ0fR2RASa/bGDYK/u7StGoL/C00
07iSCAUWH6ktU8NDOHI+o6x6xSt4SRT3/3PJNGsMmPwjHpPfKA08074+HF/3sLMZc9kboWbM75NF
I1MUuZ92hZH2zvdWMqNYaO2qJjKOx8rD/UcPXnwjQqowASwfsXvk04eWFOViFPNJEI+OKhze6rwv
gAtq9xUzSNckQhk78SVhb7CPjFVMYL3Uu92uQK/SXldFLmStiBw624Q/C/2cLxs5VcsnTXj535Ii
T6v7x8PBsdGt7URXShqT50w9bjCtbXUNygKH521e6y7aN+20ixsFISLI6xlqcYM0xGmZAkCE9ylI
WIfoGi2raVNWlsij79S6WBISsNw5imqs3B4M0/FnikH68fXU+Nl9r9cea8MUETh71x5yL2KAomJD
bocOnG6U4OXC37FpF6K9G4ku8dKGRhT+TtJDSuE6eSvQIpvHMb4ni6f8gLFN5Ccas7v2JtqeW8fA
2+/olJ5zcbc3Ij2NbBInz1WpbIrxYTA5UEznLLyYUC+a4BhtOAaLNUh3RgtMjAJvcPi1py7VfOpf
QxBD3USVmrkOnbs5/JjJ02LjbjD2hLuLNxYJR/k0cHH1b08O33CWKT2/vj1NNHSgIBoM9btJomCg
X8XnhiBBg7VKcwrzLRP94fZYatlnZPVGnAnEnpZP8BQLMpNfG8VTDmZmtRHqRNRBJxuRco26rOMw
2Vhcw5h0BywiRllv9B7DX0pxhYJToDCN4W3v9qCiG0TT/Rjupanjfy3lNBYxM2cQM9cRWA4GRjam
KGBO4f//hV6r0AwmhmzxwucZ1NZIOSfto4CAqd2XU0Orc9mt6qaQD+54w174gVW9mH2tCCFHSqDx
Cox7N4nC3uMeB+NcGMF4dXlgvYTaByT0DFREK5DkfjiGrvV1cuPBEGvjiSFi7bu+xReBFSCxbMTv
rDOnUJ5y7/pDjy2ghqnNRD+SruRcXuAd6UUzdc6Nxze9N5u7MbAjlBUJ5sVCHaF8Lj2Dtw968uzE
PC0m/4PiTTJBpoQ9C5VZGD54y9ObfsoiVWO/vNEsVsodewlj1yt73dAOY6ssiBP+uruQ5ntCWtgi
CNHe1yiOXVjQl/bhzdFD1h5afkTGkvnBJms+UfUGPaq41ycxh/30k1663bC1MH0QiwkvR4bqKY//
j+4Q5gKC9oyout3FNqZ7wcZ/Hs+N1TqlevbV4eaQG2ITtzH8mearoo82PHbshCt8XRWXbEkdJwGg
e/fSSvxc+hQaQ02V+53WZuZVt5dCbWThMkuO3RmboMIlkgVX8C5sT2kaHLMC7ttWnWbmccJ2TElK
mK0EcNhtEGJRIuQUOFx5JT27A1LeqGx5g7brLGzaKJTlH9Otuizc5UKxb7gLyGrLgzNHji7Bb02f
Mp6dVo1g7bKrrvKFQtxu0YlYH54l438X7cOn5s3iaeSK2ht9m/k3J8nzps7EAtpDUjdiskmnNM0s
phKdH8vxY+f2L6wKmdAWUrNU5t+w5fmShO5T3z73c+nMg6K7P8RqX45kHHt4DI8LlS/2MsDyAAQD
HggzaqMziR59BzeP1eCiJ9R7/KZvcgZHIHtSGdSs0/s9D3ubA8H7xyidLS9j7S4eekuQ7lmWW0B4
v7x3E+QVtcHOSUFnA4hlyNQ2/3AO/7+VqIcmtd/qGCmJOQXV9bwqqZAOjS6MFCC7AO5aN3dRwFha
EDC4p6L814qQ0rsaFI7m1sn6kDa/hqzCErco0ZBkGKHHTvLko7Lm9AceIsnYC6l05z3aFSEPLdTK
fqk5XSjF2FeQm+w97wnkcMjnZpbNJ5A42OE1h+IUNYxMhTO0NBVCF1voLwtq+9KXlUxFlLCf8fDu
/uqvD+5u26XfbdtRmIbPm5peFxEPBbZlT0NWxqeQZS+VV/eRr9qb7zrwHu5jK+KOTaHr4235Ggbh
4GNDrlgD5MI3HCPdYWv5yybYQYnMiFiOM+cVChzMlrv2UFJSFadJ5VljjbTymjIrkyLc8RjeL/RO
NOVT7a7KSELjgDRyJNv4Mvm3cGZaMFMarObcKaXLnQyvGx30OzhTtMUgccMNA0abhP1dLLC2frjC
ECejJpoH7CdcY8KZ7+TIOEHEjMFqrMp3pqhTQrfTy7QuJbS424KD3Quf32/7zn2Ff45PF8J5C9fe
Ze2wbyXlv/WOj2vbwrJPQXuvBC0lHnlApgtAisieTmIOPgvpFLYQIsrLXvgjmISOj8Fe6moZiBA/
73jh64hiMrOhQ4qYwzjw8QrBGpDfKbnvPnwgVD4cyPW12g05otVXaOiMOTzJK1HfqmfIVBwTBZUd
vGGz7t4/K7MacdUg0dcsz6qWBKi8Yz3frOyUp2+0oEMWytlDGjx5dzB1Xa/w7pZN0fJz/1fRwbJf
BGTswAFOu1gVXJyk2tBm+GyD5dbuJKPMC1QS0gVQeCWfulvC0FofNQKC9V6UnZyhdzzlirHpZ1yE
vgJdnZbbtS2/uKpKTX/IgzAaA473rRsImhkT5TVp88LDNJClOJOADYno40rvFFOiYPoBBi6Fk720
uBfIEw8h6k6WULhuc3VsqTWPGxqg6hBp8HPBdz8G8iWNjgEEwPViIcUlUoAy8gusSU6ua7ffoTdT
L8+qvgZlg8mvzQ+f7AsLMYKDv3P4cV8Wr1vr0GScGvmUO9CSublWLPrQeElzy0suRRN7ynsflhmC
D05fz8GS6nIXsZwN+C12rkF8OqR/WNJ/40QGGaO+R2+GIbRFXotJ5JRxKSrr6x4SfxUcWVYF4vDp
WI9Tkgkr2PYmRpO9XJu9AwD8Swm/fqI6vb+rrwGrgvvUVNjiBXzO6PjbRrTtOc6EGZg2nsRxw4cV
P9/GeNvNNb+wIgbQdKpBQkxsZmBtQ/70GCOxB9YltrKCKt4exDg7QLAhKDQH7hBe3p2BWJpaxjiV
FKy4kGAemBrBYoRtz+1zVmeIYKEqvVlAxqen9PSVUAW3t/YEb2U2GYWV/MIlqERnqvXzeYNixaob
xuvXbjCqwmN5DpdEQIjgc6osalPMP3ZVRPUqV96vRH/3WAOsvX5VVhoPkLtYeuWWZY3PILFVfF/L
Kb7xlv46+SjiNpX12QMLHcTS1mYflJRxmyX/LZpB8ycOJLT/4NBzF6dtCdqfNFxmUBNql8l9G/WD
sWNpADdPA8JiVnyqXxNT88xp2xQURSuQbWPgbrnykvPDfw1nfyC6N32qIm4BKSftBeD87nagMOKQ
rCaeUmVbKL9hD3I6EOtQQvuLJGw0dnnhzZE01hHZyDBEQ4LW67hzQR80pM+p2TxFQ5OCpZv7ibAM
LppqtTCkLc2TPnN9MstOmu4mGQ483S9F7fpnCXwdYy59pCotatsFyti8XXd5r0LYwY/Jh/VYgQ1A
6UVGZjN6mAFxlp9Pz2xB81SD1i09CsIM/C2Q2zmf/fAdkSntB8e3haNp934pnQrNyl2SEh9tlD8z
p18je+YxT5RpXJVf2FLolFkW909mPmz2cBeNhHJ+EuJNJIPn2ct3G3vxrkluAIMallLXK1x1EeYT
nAkgin/7Jp4oYKSwko3szjxc9yAEyVyQEM0t6/eEAXeRAK5qm+M3VpNoE4pXkh4RlUKmNEuyK+RB
pkQgOvmMhMm4CpgaTWpiYT49aXprgK1jzovolxbTe5/4DpHTPyp+/8s6gTvnNR52iB5LeRGsQG7D
GZt86YLSFqDzXAIajZXCzeBkWXTo2W9gbMw0StNqT6d+pnjbkdg3Mz5zdXMGzPREIfOLwFP5mR53
Ys/ZJJF9w6siC/3Wrfis7PveWsQR10n/PUQwfx8VSCSpfSkjEJ3Qpvabqqx+EAq4YhgHVatZ1aey
1aV0tQuHczbP/11f3qpguoJU7F8cnUitbktEwUhjziL2jwWVZINsqz2FF/XrkvkgHRcdTg2OnNEV
E8+jR/GSHVzVf7oBjlzFINu3xdPqrs/wUVJsta1z7vMlrfaXDMzgtzRbIRqgDxFbG8CROWK84liQ
rsnG8o8hGOL0oRv8Mi59AY5nTmvbubKJ79TtZ25PwYgbeZkevJqlLWipx/dB1FFFiEkJYbX2kUm1
jmUa+kWcj8OHInSpp2E4FO9NXP+SeaPuh71AN4M22oL/uFzqHtcx0Iu6e6Q0UzvGm5J5c3CiGB3h
5hmhiuw2KRyEhIfthk6+5M44JSGEwnLRVRx13kYaTfc62SWz7CdL5wA1qkQXqHCFXp/deYN4JLYN
daOnqVvy5evpDD3HydcCDeR9G1jixJjU+d73MDq+h3nOFZbY1pHMVBRgBMIFbPdAAkI/4IYEZgcm
d8s/2DhTBmk1OjTpxPgEKNHeiZb/Jh5x/OwBHyStU50lQ9o0E9nfsyNUN9kJijrZQTJgQpvSEka2
n50Iz1kPI53atU89ahKU0pkwMv5yuM+yLNKlkSBbMLBSK/Dg2z+pR5Hble6WjBqoe7v5QXBgzZic
CgPRV8H2J9GcSfIEuV5BjNdCvVezdMOG1peCc0WfnuoLubElJ4XsZNw4x1LaX/lFlfGpTaQJWbZY
AzxmEtrR5SGBR6LKoem8IZCF7Of70a9cO9xR9FqJryuXnRVUwnTy7ilr2C9SUW7SLzRZl6R6I75v
low6IqrjdTHw4gq2vLbXLXtQJ9nOXx+LnTlWcp9anCVYzU2HNyPC/hz286e6hfdc4tZKxMJxfeuY
SqBffqKnGcz9pWpDR8W9DZZi2TQq286bm/6oa14RBOY2fuaO7LGEOATKqf4labd583EZ07eAl4e0
OSg3LV8MfvHry9a3194R80WPi64xD5h7K5jYmWw0z0JVWFWdekcwUghU6202iOHCA6dgR1VO6KRT
ZB87mDE85EMd9mPepRbK7DO7okUFJtF39RuadvUuV8ewKLUXtwmJXbfOcsA8GbcMyjRVmu1jYeRc
HNdbRyMywwmYXfdkDdwg7YKonNmeYoRmgYWMlKT2CWF9aTzdYQxHOanJYQisHTDgWIve0qwds+/v
HNwiT85DTOlt9QsrPZBt1p8H1CCNeEUwfHek6yW3ZsHLnH3vbi7CdAuMfO2aZz/3R5Xu+Ls/jrOL
4G9KmJkN7KQI5cVR/NXl0GzvIBAXZ+hXHBkiutpVtJEJ0FvYgdA2W/GeYsjilc5bfSVvA6O8eYBA
qyDPMUvbEHaUQ3W42CbNsyhUARm7hD45WEDenhwGIJX7Y1ujgkgE4QS/777KPUBmhAj5K4lhBPty
Avb6UQoW9qXTgo7TsDwYse2rA8J0g+9XZMyGwjYPiEP5etHG4TgPG8m83zA02KfATn3k0A0VV+Vt
VIF8PbIRg+K4cYkiLNdrsn/9EHA5k/TZGiQ74w1VSldHzavq+Nc+q9G0sLkSl9SohNgIDvL9MAnM
38oaoq7Ir0f1iaI9/91f2i2NQMqsiIg0s6nFYiJ9trRNmsDea1AYPrwsdFx5QfmMHSFc9JuHPLXL
gDNPDhAAgqMkZysestzRx4UnGX8VnMTmYbPaayOjziU4wTtOX30e8OqWi1EhmNlAJ8GlTaiVggie
nWM+cyegZsrMSKSXicCAHCvkTC9U/YFdyVVtThbwij3COF3FXW8+iRluFjTR8p7BDEDaLBCBTY7V
M7n8L3ONIen4y7ODwv3xyAKR96gyuHoC/bnnckbGGQcafo1RM3F8JGqrDaF2Dj7iW2CmEd4PLP34
T39zr1ISbDFgyIRzVp8KZbu2AsFiJKVZB8TBp0ZHnkVQWd9TVohbDNVVoVY7WttKRFru/QT+ut1N
C/BjGwhuEvt56UYkdIO677wxqFp3TSW0b1RGUntdtucWK5j2ScoOIorM5oU0oRoJW72jrLKJgkXj
ml48oY/vXjixCImakfJStsPsbetzAeiW1EkCqjd2WnuuvMjecl8Vo36AQ/tXs6XQvpvbLLsjKg3v
Lyrvr1p9X+22oBYfvEiwFPb/BV09j715dT0Dtgv2W9seopdSC4hOszEAo8LCz2rYBqZEAc7AtVOR
J2vJ/glH16hsUbBlFcLDn53ian26yMPgTSh4pFtRuxPesKKXyTgS39q3Kug1tgbxE+XOBiCeQO/v
a69itXO59ZF8v6yCr7WzAAw/tNFflYdRsd5eTWLLkaL5trSbvJGgNEgWndCcPvRrE6embIRhrEMT
jsjnAUAA+KS+DtvsooO7WCbtryc4R/VslY0GAYOwBt+HgpN61+Xnz85ltZXTrxQGWc0HfN7bPg0f
V3YFNuoid9YdIZevUQyEtFVgZ+I8UlgIGInTtzh2WgHk4sa1GeMzK4EE1u9YeHthGVlkRe8/E2JS
yUfojjmb1luODweZ06JtDxvjjag7vCvdRcnLmIFCPq6WcAdLP3xPAvDND+2DSf4vgu91jpQpJtw5
oo26gY+d2QETCjSI5lytN3Ecwk6X7xF+bO24eZsEjVykGwXx21VGAQO8GCPsxTaKpQs/UCa83G86
YlUz5VgN6yf857C7Uq9xSg4lAN57uU23M7eVlc09M3l1uvMOf9pOYjHKHNoeBOAQgFnGWWADE+5k
KLLZpmm310iZxKv3WL7caOozBpj6sXQFEQFQPS5ilK5NPrbEBSuG7M7Jmsx5jF2NzQMseA8DxtEd
HEbWFQ6abM/YcelRwI0kwJHHv3QsiXHZlFCMqStRuB2qhYRVEhq5QgtsEQkuHSvct8JTAb++4G6Y
QWZ2U8FzFHd3tNMeVVWCK6kokBDt/CimGxvC5WPUJsaHithFUFmNE9PbQ61saNMzi2Eug+6bmXLE
sD5do140dp02X9jVJ+vejy9YO1clNJBeQ+OLGoGWNYtoaadU2vAHal1YscDSRnSBiYkW+AI1X2Vd
Vt4Mnxbie3pAFo2jHG3xkUsyvDDLW/FDeIlB2XzWqbki36scGwGl96gAveeT+FXMc2dpcZYzEJTx
2cnz6wEtI1h9/vdtblfKPLN0JUhbUnQ9mn29b86crzwaO2pUBOZapiLqrnVl2FsNsD+QbCxmmFdt
mwCVsXSEU8BDtLWTBhUP6GEj2ffegsTUfsuh808tK7CVEmAD5jFyaWvuPAWSbqmcnuPIG77DdQfa
HyL1vHAhZyB4C85awXTEsOXT0Hk8BFsR3bEId64sYujg7d4bYkLxwZ6qy+uRhGBMbZnyIoHcE54K
exvydm6jShQ5V4bWvsVclRiXs4nlxLKfaytipLatRyFGLx18TQ9xKBg8d1idP8O67sf7nqNMSexK
gC/1UhgC28gAFJl894mI0GV/IFtAVhiHRC9CkgQEIEIeZC6VRJLLizB2gzkom2GsiJVL/zS9Y+64
jKvpswM3jxrHoxq2oPnN0lpqMZZnxI6LJW9uQvgxq0/9om3/nFdCJHXy/JbspuWZ1VKnNw4hMJ/U
DGV/G1DRHGT/Hr5YVEM8o+lcweA+cQpuka6oTM8vQE/+4sL9XJdQykYLsa7AaPcRIVUYTmzHYczx
48tqjokgQdjvEqsx6m0jYKNstc38BTLFeISvj1aeMABh4JsQiUDUthQma78dI1VmluVuxgAPZviT
r78GB17nQ6kuCvuyCasYNjHLqUfedZFrcQR5OWu1j9ZFT739L6YVwihUl/j14aAVZ5UjysInI0qi
i/fiUjjZSku/7LEZTh8b/fGmB7OfmMUmXovU9yAm8bLlhgKDBSIJMWMprQpu5Awm5d1uxxJpf5wf
b+bC8yz0kMXJNTjXpZ55y1gcpAJSJGrAc1na3H2nIN5yqfGgp7FUuRlgjXqHbrHp7OYiVuV45REo
diEafhJ5BY24hiHL4TpMvTqKaneQPDuuInfksOhwiPork8vhasvaLDZfZ+Tq+A+p/VlNuYBw38uY
1CXGnXTq/kiBoQvJDFLn47s8MNBQOy6RIuv+rtvdX9NPimn5BDpewNpkrszUHKRRHMGfyw64z1sD
7Ve0gM5wLPHIlG+9WZ0cjfHTH2BVmV2vuQgS73pXh3Xr6JPx9svQqV9eDneTxTssyvBSpdWEDj8p
jbBSJhjeR54/HAjxRFkIxqrCEkVUB8hFwbImHbPqPZ1wQJmUY+bfgGpXmjowq6KvQKacv6meUwld
OvMQohgnEUj6taljlsla6F8AjMyDgBjY0/Bkuxct21nxQHOlPK8u6rPw+Us63J6JTztiJEDHjb9j
rFOZ2SA3Oyi3FKS5GKQ+JLqigN1mqf1w44CZBjrCrr4lhnommdLHGGe2WuB6eHhwcikDgXajT/zw
71etOAg3Qub/CjIdxhBCdcmbSWM5xH115ty2vJ0D2VGf73aAhNbFujX9AkvClzg5mqxQJzzZrWKS
gDlIHHS7p36LrjWdkYloOUJlYtqV13tNWbEZ9tZM0bvT/55/NEfHdOBcN84YI0pUnDNYnaG1qZX1
ZO4Ez4szLirHZJYBwhlF1RHsy+sdAxFmfK9Gl0AIqPWOEpOA+lEV3xFy6U2kmsDJMi6nnxrkTTHM
aPmT45y3bpAm4vJv/XWtMRg8catp3ls2+Ch2FyV1Evu65Be1BGOKSyEpuW5dDGaod+TkpUrUhhRU
9GlAH2IQHwBE5D/o/KoGYD8dtYdAw8zzY5SlAu0S+b/pqBiWkKedrOh9KDuJgW5VCTOpyJQ4mBkg
sM4EfKnOhjxSt+ie0i5sbhmDfSasitofqI1JO3z+pDENG4Z4yvjGDwfzxPanscFyjS/2C86OMqS6
aX5yAVOXyzV01HTcYmnTK7XIxL6aWT+u7OPEdktnf6+h0qqJFK8+oWZNbcQBGpdju6JcPmsq1FHi
bQFb95O3UgDDm2gl4WKZcjKCwe42UDfHvTdDqaU7Lxj1/GTgaLtf0aJenWm7nfCG8itRJSely3s2
U9XYbvFw65CdWY7tO2AZj881SSFy+BblAeDH2ety+hPbppeZrYs8ODL8Er5rIg9hIZjCOkfw1c74
4ZSiYh9WSHTW/k3ipY/fxYm54GGKkQVuh4Gpg5dNsk9atUmLz5HZYV+J80BcWeSC97rJgok/YeFH
/NScV0qKhA3Xi+92Z5PA1vyTTKFOr525PmiIbsW49uohUDPPEJT/kibvI782S2/VX2Gg5tsRLUSN
oJUA6pU=
`protect end_protected

