

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SYUpj6do5sFTflpbsRmqzQKFPQDYrJyRQArefGItBrRpeTStPf4iOexrlL2KuY5Tjxr42gzfz2no
s00d/SuK7w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NR3ykkYMNFMRKu0xHAyt5DYiOktc2YTf1JOlIURJ/ThqHJccRXVvH+Sc3vg9x993epLj5za38fd9
R5dBjv9keX+G5g1u3CtBsdqXK+hNOz/uDIy23yxr7rHw0ImE57TmiDkVMvMwv3eYKhw+6jZKYes/
orVUKkqCIC9qrUn5RTg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HlVxjhtCNCKKX+WIZOv4bglrDneJvrVwpTadJxqH8bLj9DfFux8A76EOB2zOay/g3B51jEHFXs1k
cSPeVifBOPOW+4hnoJ3TimbzQC2WXDZLrgI3HV0zvi2+v+260AsNylQU2ks3dLwbxExBHvawkhdm
qLdLQIFdyzjRMD/G+fo3ZOpvx7tOdM4iBWXd2qur6t8wJth9ryhPu98XGfaQXlmJP7Tzn+0ub08s
DCWHug4G341eF+dWmcugGtWe2Ca08XjibeU1gRioez7LDJacBlMb+me+eJNl34Hg9trbjeo+4u2p
UhjBKGy0TbAWhSuuGKcCtfIFOUbYcwT6t2Yt0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DoI+R7m0zbJxCq9A8c+QbVnIsy2kNMG29/strbjpu4rQhHX3C2LKQKMwC4UXbs35yFBTN82oCtQE
LCzB557xK8srP2DUb2FdCBqlo4nmLOUDlZKHLRnMjMktj2MJoV0ExtbMFAErwe3zZqIBchZgf5Be
0C+OuuK2xw443onEGyA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jkJi3dDxF04M0w5noeJKvbYmN6cGn5suzWOH55jYT8k6r3UxrWZdHPmAWJgyGzXTFa2rcCzw1zFN
8CUT3mqhUaMicnmv3k1IZXtmQp8LLIMHIhFQWUBUexg49lQQHlMizPzJBAEcyMQJQl2JrQBPC4y3
FtPjOGWfsQSXXVoSz8O8MOKUSTmbuzqKeAR7KYOBiW1PqJBZo+vP/teWIw2p1h9/ADBVH7fQiL3s
cyUleDPcPx934u+grxqX5IGh+uK/gO42i4Ms1tDDhMblp6piYQ998xcC3XiMWw8hwmR+KGnfqU8Q
VD22eRbZMxNB+D8sxEO3PnV48eApa0h9wT+rpw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30848)
`protect data_block
icomnpvP67hYg7e8BrEWnA0FftuqvWeGYHCNdx9zmAZSS8/PxL2tFmC1d1fvMeysKIuMkSNjkene
g+U23/eHRmofTajIRqkOlPFlSnbmVA4q9m1p1WYMtR2/wMDsVGwqYNnICTh/8sBnu+jRG4n4dCFa
/2iki6YKKjx1jWdzN8qBCClcrWvv3nqi+AT5bWMcLf1c8uCw0Y08EZaefumG1nwuaGsXemIz9e/1
vGNUV/JYXPrCra95Gyo8S9UYDYoJ9suWsURzOyN3GrxivvIB81vhV97z7aIHYhcP20Qn4PoVRMwS
Om0M3jRSN7xZ3uafxAgBEMScz+L+xWhnV4s8LqMrDSGxR8VFI3CzLqA4KNC8AHU9ad5fqC8Ah97f
btBELfIMCBEAvpOKfl2qU3aFe9jvRmRssFC/kP8hZcCZD80hE9gQnuFyPpQ3lr/uyzQdOlZC/r10
REtEOnpbNXeebshrlKiXdLtPW/EMdTSMuuU/sBVqHegRROvMETmSnug+YBgKpe7mpy2armDK3yqz
6/DIt79MZWn4TGaeTtcUdYUB/oRCQUXwA75zKs7GFqa0sWislVDEtN802EVgv+HtHL2H8uLObcmZ
KHM8EWIgEy9xy/Ji+r9iB1GdBq+0Oys2wT7b/992/O01OI3kvCguLGyH2AjuBTnaux9d2x/02RIA
Fi9kLjfhq1dgd7dCfP9S29GuZg+2k2BK+JXIzmM8jvjNZL7n72B6JL1k5KHE7dbnuMcRVD4nqFIM
CVsjbm5ShPPFoCzN1iXj2AI+62CALJ9NplQBn3IdaEtmrrH0PXHL3EMHkrJMKywKHxlC7AylfR0G
9FPqAw36h4HiKV8J+xAk+dL4MyAMF6wfmFthu1xpZnmdK8IEEkv3YIyThGSqL805q00Ih8fK8tjw
S/N8y8J1+WKtkHm0g2Vc7i3bn+0Nxh/WZlGLFAVIijz2LJobJjcLklrvzm7n/ZD0zDjb4P+MJW9W
zMWI0JpcJgRwGq22LH5k3sCgTNaXiJ34e/AfuyIQfxgLo6AvaqPNmrXVmsaOd8seZsVw2nXRH0rd
r4RENWzFMJ9vQoWMazukCeTPT4rG5lajeP+BbLz6rEtZ5v2+tV5UlZgy/65XfUaFr4v4Te7sLslf
IexMqbUANvHWUFBxiVAda8rXFTVbIjdK8fueVMGDwKGAK7pFaOeDgR7gKOMn3Ym4H1iQPlUu0DH5
F/ezxB1G/eti0Ds1RqyYkbF/mDErOEFaCWx26aYy9Oktrt9Cma/8UNfcn2iraHeGfNPiw8C5EPau
nqndXKMvo/mlyd+O1PojNwuK5PxBlbGnLeEAqLODtatwjgTQLoX4+2pfZFeiIhzL8h4R5u1jpYme
7m/1Sfmj1VDusWaHfFLI00ZqSITgCgi9LlcDVG6U+fNyIDLjlff7GEayimtqjw1hraOap0dOePo8
SE+g/JpLt9dCHlrSyspJoT/WVTWCJ/T2HxteP6DUSrUqlHye/voLb56ILDqzdWvSaBx1msyctD1O
c4rudGl+FKyv8zkeE3BsmgBNQwrkipiW+bAYP+KGdukRxzM4OMi5D5MbM/uiyn4gWSmkTObf58sY
an//ly52nvHCSKjWLnNfh1a9nJjA9OZY0qiUszZtx3VTYoIl25ZJhQcoQmTvPYQxvU4K10LdV3ga
d99zT6A7MzqFwDf9yzVr0LMNNwzA/KNo/ZpKJtM/uLaReZ54CUeS2+T8etqmqo7iYjbrWuk2uoDb
OmG6qfYKmeRWPRVKWsefnD2NYTkG3H35ABLMLdTge+spbypiguPaXLzO0+BKhyJoYu4rjT0+oSHd
J21oPI2BfX+NRpX5t0anIk/Vtvr9mxPMOJo0NWon4CkEKKlpXpjGBUSKRPCBpIC4alCdNnc8t73g
HJ63TOFy3GuJRoTWoOxP2DyRG41BEs5QlJussuS/vbaDpLSpIn2HNPLVhk5FAbt8rflIxmYjWmwz
WCYtnpvA4XOPiiOuDkWZHBS2WZryxWf1XfQbj0H4x5PhjA/Fiph6a5ptALxw9F1Z3IzI8vRb06z9
RaFO7xbWoTPfm5KE8WgE3qzTKXFcJC2r8HmSBg1d95ZJXkMD+4yVakiVD+8wEanOu+7ZvdsvCEUT
9eTXJexOdTngm/GlfuDXYPSnaH1Yh4IgUJHcg3nXN6zFYhPVQecrgieMFy0HP2P11NduXzDMmG/t
UbkTCeiIuLB7kPlGWWgF1MDavLql9NFPuUyc/h0OfWbvAD1SGqNnRJt2kQP5XGw8ZHHzjQ41wX8R
daCDz6qVH49Kjz9IKXowSl8thFqmXqYhbzGulv7K1/2pk6UW1ZNhJHtdE6fUl2QqvhzYBdVSiZXw
PDAiTdQBo/1hsFFo34IQ6THuUPUm+ZCrgtL4/Blz1wjcdW7Fri2etM73kUE1s0UQ41fM4+jNURIm
ltAQAlKEddQ1eHZDxnjUUFAom6lGIVNFLx1RZ4+k642R9aSFa7cWppnBe38KMnOmhq3iUJnPIc5j
ICsE4wpkC/Js8DZ2rwjHOBwxKVmIkSblVMty6uvl8ScTCKR0wun6/9Q7ArHIFrnnoMiV4IDWK5SG
FfeMqVo0uBjvFbwnL2VXB1HGINgjYBIuigpMB55g+Hjirw7oMOoECzXCsefZcfYj4vZ+BsRotIfc
dLyKLOa63eHQ9abQAb2IJakLTi/GtInPLOLrl5QKABwLGcdSTA4k1rrv0NXZJRFYdC7Iath4RBJw
9zw4bFRaMi9hC9F61KOatxujQRIUFJc4U2BZN1iTaTqVxWjpYsXgrHZWo2h6+5nI19dP77jr2hqm
o22CnKQaNNAiUaAM/GCHe2IiOgtj3B0che24a2gIkZGPLYHSma6DG2z3eAtVzOqf2t1W7J0qdkX4
Rv0Bz+XUqOKG7yFf2fx53wMiW7I083ofF6L+TtJmey4+3kz6f5g2/iOR3eBZjYEHhx41BmOcMOCt
To2Mq5WcsPlsY7T/jXUFtKCZUktCRR6m4pBuQiV657jsbBQYR3r0TsWIgtc4veg4oKW9Xh9WCG9w
RvRGqB3ANY9pNu0zzbddWCOS40y4n+3a6kq3JVuDMKj8Hk/EjjlKpZvLhwqrC0DuA45iJmR/tY6X
WTi4pRc/MiwrsX8bl0p9k+H1J3ty4P9lnA1RTVjNoZh7/Wvx35V4shROqCxG50KV0FtABIFB9N6H
qFgGQbmfvAfTTC7tw2uYakWlUUbtgv5wVG9ucIpgBqRz18X1CqqZzNhmmumpdYvC4JipBgAd3R2j
d19qHTuwUAUj9ZGcEfVUEP49jqjuWrwDQxS4QvXtxVe3zQUFPhsXYUqE+g2qP9jTG+5Du6O2HkN4
xcAOxEWmxC4ierX9copUtKyHhrDJ3iMvn9FcsvmIeRu4HPyUxoIosFnNyfLDJFGGK7VdbrebUFQa
fPKaC2GgZPGls2kg57DeWDgVluELstY+MFHZFW1RfqJ7W0XuU//fxoTzP9Z3Hqywrx0tRtaJRkk3
XFLgrbqRYDt1kj6owmd00scSRvqNchA1qFYt8li5Pxo7np60lucF8ExNx6n6anwYBjc/Gkub9fno
5nXYUftaLV8+EYTB7QCuh/OVL8XEzqvGZcOBc2O1njKquwMeUpJVFQm4jVj+wv1Z1ogzQtI+Vb1I
7m/35Sr1AXpZ8/Pnrz9IG3lImhKgYOQ8IOkLPjuzmIOFjInJYxa9opNSP/MUBeOkxhN9O873s836
zWevCM8z3zfvvkJedh4r/Ri5omykEMwqplOBkUHF9FpSLBxXkUotqtMud9qns0jZvSfdTq7/Nzxp
8Xv5voYmVRyS83KpvJfp7sNxb4MXh1C8m5rZIwfkICsPJbYcDRx79EbCFUD89sLGRaDudJzwHcK+
bCrMu1UDCztyZ0DqXjhpVNqUZkihdaUXaHdW1zGTP27vmQmoJ1VQqVsaX7LKkZmaBvCSh+/12+XK
WkPge2K4spaPf2YTMnuwZQOd/ushX4h3wYPaIFEzhrvoJrW9DDwQifhi/hn7ePbiGx/pVPElYczG
5cUU9YM6i6RHVHS/v+e7lTi/0yVxN4V3ktwk5cByhCRitCoZQen0yz3Qs8qkDyAQ6UKLnwFnX65W
rYIWAzlQ/GZmK9rtAO+fNVOhZIg3fEO+5tIbASrteGHPGkKbNE4YJa0WuMp9KpBtkKvZmA5Kbrbx
9v2wUl1wMeroz17GnGcWm5n9tl5FjTu98+YnPCE6/lWqM4dwbjW74+974WuFR5DDox5hpQEV56yg
2LXQuDZAmY1PIxXOvImLiXNEJvORVKzwLtkC+o10lyDs3YxlvCRQA1wSUqGWJmSBJzeGOvyLafHV
T/uWBbzOS1BjgBq8JKPjA24iSh9d+c/YP4O/kTxjkUSz6ZyVZ3h9G8JikoYn7Sd07ILM2pw3C2ES
tEo0zBqCupbKJohW/4LauQlqCEDal5nwHPYMyFXFm1KOAIwrqkpO3q0MNvXGt2iKOA5k3vOK70K1
ttoK6uIlrE9FypfP4X3RgnQhGXPFEguygvqEwsik5KKi2dBz7b+kRE6irGl76aRBFpqH2dwLQPqI
OBkRfhNJi2ZZxZtGuhZqyrhSqZV5RwZQkJDc7kgdq5ASi3wKcyUnHnpX5bSbTjT50Z2Z5GNgV3V7
XlKE+8YB9tpklKvUxm12mzvn8r6WzK3SjgzfVhuqKZeoDsW2iGeGveEbRkId+OQGVP450bojgXlG
gGqgE/ul5Vi3V0aryB2RORQXCm95jdGfM6pb7rpSTb5XmKHZiaSD4a+Nlviu0nu9oN8BejlgIUO1
ihs+/kC8gKrhwr1JqD8Y515LaLtfuTSx4th4I8C0oZ8N8eirJNDyBpfliGgJPZUGnB4jsfwMCtkP
rOJSnMFBOvNXojSC5yoQRub9MHVN+m2s4jNebf0xwzwZta8XlMttqbmWGnLR7v+cQFHgvZzILDlQ
Gh1BJlNbkSykL/JePiNBkPeF40MyuUnFXt2vnVVLfMVHthLIQCoQZq2OFFRptFOkQ2YBD4sLe2Hl
ZOE/e0X+NhTHFyDe5DkvRHtzC0WUpb1fzoXKnM4JyogH+4Oyaj9QgCUNDBEQ8x2Y3V3RDjKA+rPU
UHHiW8TNiD3TwoCDkp3e6oMIjCrsZwKO+mmMIDR69cjGNxE47XQR3Aa1IQBvQAQOBIGoGyAyHtui
3QJVhgZoysk9WdKx9oLjDGVcfLNzJfL3XWb0xP8eP+SIRkVz63SbeBOJqSfJZ9+ea0g449QLN1Oe
xObQ5vAfAVTd3dChxGEjmb8wKWXX64CHyQEqoVy3KVD15r0STABJU6EV9oZI1wuGBmEdsWFwx12a
7etAtLaqEdWQt+4TnIaBwzsFGxoHb3diKbnk2bG4qPlhs7woeIZWbJ19ruqGfzyvdhNjfnuGVquC
lcbWSqiSMiq7rXqL8hhQY8sCEVUoyL732YE/Vi/ydK8ilquHpJxrBl9y3G3hljuZAIpMicAOPxf2
G8ihvfPD1+A5Yog/ZUY0AhtPnnreDMbh6hVx31uRlTa/HeVQDT8g6MyOa08TNDTexjqB2BqgLe5g
YP7RfCBGnru5iMcWDLCcAy+f/ZpAGz57PSAao1yyyNlQ/c4/nIJfnTi7E0bHDibcJ4mfmN81uoIq
CGwJr7/mvb+UX8zWjeW2dM5dfHQj+r5hz1fRx/AFwdtjXw6HgqMC9h+iguJeLdzMC0Cn7I13/e6G
zY28Kq4P8edr+ASz3YZd0cD1TMDBEEN8+4izHe9riyB293Ek1/BDh65vbNdxdtXkIILa8U1O69k2
cFxpVvkSziiID2+nYVk1+I9uwp1kpyKOOw4EXYA2eun/lSbWDC7Ofu9fMBywGd2Z2lWUQ9fk7Lby
NHfedAUQLPCDFoVLFA9yTQCzvOJahLUPOOYvT+zM2rAhq0u4w5MWiyKaqHGIqzImQbAW4St8aHDR
SPfMe6CKriPrGv6UlqxzhhfD8S+Wxzzh3njxyHpVcSe0VQJ9C9zms6MD6ly9rOwmajjRXEmx3vY+
X2DrQSKFPw+xOCnTY47H+be6YeiP5zU/HvFVWxsnD1FsT5/r0Xeq4HlgbNGbo7oDfdTN8NatMi6r
1AIugob/4zZu1PARi1CDz+OJ9d7Ca694UhN0KsiuiSNNf8i0I87+CK7TczBMbjF9EWxxa1JsKrtb
DGXfaisvbH89LuGHdyt0droCYILZFv5ADbedyOMWfPte0j1TFZojmaF0EMlDKGoazPcwzBDPe44X
45VK3HGNd5D/yVJta/DaF87xiXV3yzgzWC3qfmx25R/VwqDZD5CHSmOivKwQsG914B+sl6ccOt6Q
rUaE3LvpLrYsOxXZ/gjbnqaLgYsRcS9MIAZfZ2X8SUobs1iGMSszIWaIIdYqIT31Isg0DBsackne
fWDVBuij8lI3T/r2ve2XzA1Qb6Utb0p2wMvH0tq9phryqMD/XykHLvJ5OZ0p3i8gQLf2CzHPRnfi
A06dyVxQdMoGjrRH4l2yPCwV567YN94BPZ5dGptIzQjqeIXGCzhSHA8qVTBmMaMqDFxtYeHYtODr
K5dRmFTHm+2lTYYLb1/t8gEHVtgFOmWCPIcnPiF0BL8UsCCWj72Aqp0bGm5VB1tCGoils/gC2wsg
2OErIS0wqUBjUDk3bCvBDem1qtUhAPC5F1ukXq5X6HdxTmXrBFpdYZJxaV7GH0iZ7MVW42XR9bu6
AN/211813O1pqWOaVbLrOpquyQqUNPgmaRlbanYKK/RB80m1fuwW5n9fTb4fWHZRYRaDtKspUZPO
03z09lQewtRiw70LPSXDcNyGKUfc0hdfJcMg4yiev9Bol3mYRV49xsYBSk+/Ss57at4G9Ta4Vvk6
xqTgW+2WdKCJ/dU7/JdiQH+k+d1I4KiACVQS+vt0q4SruBLz9QyxgKVIku20E/izZoKeja7HTRXw
83Ai4cgkt06Xi0TvO6u3fdcnrRQyEFPkinV+cG0B4k3ZwdDI+iiE6t4HM4b985M0W5JjoE9E/lmR
IU4twBRjPgvETl5gjA8Pnblcj4FPk/mdrIGqlNDTnCd3ejKI+U7sSjfsCnrs77LL2BvT1H22FtoV
KO25hXKWmA5LfTUMuPE/QV2pQbhwZuUsze7XRe8jZVtFzFcHzGsXvU5/Z4EVYnIyuTkF8/sTyhNT
OpAyMaMpvm0wbfS349ptlyCOrmhkGCNTSeL8B8stS3lIsHzETWUU9WcuC8iRf9ONfAqRvbNmSFR2
WvhSto1RTaoXoQdLCCivHOKLK0QpoidN1wKb5XvSpkmhxduGpSPxd+baEovf48fKlMbN/Jis8cLH
K/gn2XzUaMhnZWwM98jb7SYYz534cVnR267woddnhOlVsewHl9sUML89pk/I3YwuLbE1uj5OeEwG
zD7AxWy6XQqLF9HbuNgAjtJu0ml43w2s4SBNq3sV8PToGLxjhDMprcQEpZ2ZGwa6H0N5v9ixV4Bz
4xNBzb3Lwi4NQRi7chHIlL9bsbgSLkCke/LbIz8sX8hehS3bQiF/0hKHP1H7nN4oK2wAtZphS1qq
ItEs4MPsKVpKnR6e1lKoO4l8VehCWAe6jdjgGoNiwI8EIo0rVFw/+o4N5Kdyj3ra0aR0QgZCt8rn
/N2aAPzNMQQnnMNH2GdqkoiLkcKArQss4f0/BkUzhCT5cV0Oawni/A1mvs6st1P7YMU5wgtY6Zn1
Wb3eVZvWXAy4lX8iAIUxuL7VqM8jVvmvcUOK2Xg40SBho7hfPx5g/WeSvJS/nJ/IgUq94e4WKZdN
LgzLEP8aQuzoW0+6NTOqdkBUvHn2mySWqJQ6OGHh8KBkV8s+0TnDqoEm1lxbCwadgARmhMlqaMvs
TZ4a/vgFjZ7EGN8E07RM0GXHQfebg0SxXuoatqcH+Z6k8CvErtwbvMPxAJRs92tKeLylr7kYrO+7
hxNceDfRWNeSuuVDMor0WcmiMC27OOMFpd7qOV5dCk557UJoxTjxkmLPfVY/x2ETn/t8AY/IKiLn
knhHZrFYdOlNlRK1eSxvV2P5k4zZnW+4G8qYc/zwzXt9xSrcT9ZquDlLIaTbB6N3ecAq+ahDmoqE
jjWfdQACXojtjhxzFTiXFR6TEOFuS0z/ypPgPTuZCnURAogz9a2TeXY+/ADUDCXzrpYdPGeC2osP
+IXnkWBDA0xhXHY0ul7xXNGzZ0tXV9QNNzK/EHLpqCLvuugDxTr1abf0Ua58GcAw7iQal/odxRRn
/Wl9E3qLnVDm8s+iCnOqzqNro5LsCZwN80NDebNDMjj4NjrSAsmCqbQKGj92MngPuFQ6rrziAZEy
tJR/aXvhOTE/3sIj70hfurbknvUhQRjutLQL6aUOkmouiqcTDHu2Sy/NvZEqEy4gnyG2zOcdyJfu
mJ2jb2cBb93fffpbaPJy8WJf2Pc8kNvaem0MXezypk30xKDxU+wxSIu9LxIBFqSE2SDI0wFFk9Vx
E47VV09K+w89zGNH29H/OxdWDAbfJXJaM9Rxi5KaUHL8mOOn+SXz8nqpaVo/9cLQauLW2+4a8TiH
IbeWhR+NUZqkOdC6DV92EZGJp2ia+SLvs+0XuaPWrpLnG+n6d24wQrA5XHyZuzmlvjujcPaIXFqo
7DGhNjsMjBZVQ8eKroq9vipD/zxH8XVMzoLA8Xy5VFWQDeD6nItcQFke+J5sRBke5jrjM4/6wcoj
zLhIBMS1pTm4JgQeOa+WikxW2rvZqc73EsnlEAuy58xT+YBT3rhJeeybZBN9XAuKiF7r2siUDTCN
x8mPyxkxD2/drrDcvWZVqjuas38xAmVWZUHHliw7g7a8hhfTtTenJeASTMNMMzabsa9KhH3cnF14
9TSYs2mHBP8Nu5+MzpScFTeTDsVzJILpYXDPgHjA7+ZTfU8Mx0faZqQit4XzqmwzbZOlmJhp6LHX
aS2HLkdpIvWpZqmeoh657GANmTFAy+ILHzfRqHwgu7i2j/ClKFVKfNtLHbRaaL+q1FXPrB9E18WX
AawnGF6xeinbQepII9155L8ZOQRdDVdM7iil1mK0Kc3qMHsTEviQDLo0GK9C0DkDkfRp+wZKnPQN
tZbyqBxufl6tFAvOUxHoNjBhOB5V1je9bkYB23xIo+PwbkmET8Lj6r1SSS1IDaiw0tOFJy8eJNO9
NaBO3Q2Sdy20FivFTgs3BKtHmEiPhdSP2SmBXDCA5Zy62FmlT7SxaU1tjp7Fv+eDm3GVH5MmrxE2
XiiJpzWWAGWub6z1T6wnvOLeX7WI4b5EhVDcwQHzyaX83/LnhJIGf1A49Km5izHzBiWjxpvKO8N7
Xpo2O80U0kKPWh03nKg/zf5FAhIthsT1Si16lVX83zIyLFpIc3cBkXzDl2S6jFUGQgwR7VUj8UXE
MOhlADI2AG4+Q2vVshU51mS4XNDQ+0Q388zjQEwHs8d82ygrVJ11SNmn/yi8jTZU+FShHj75Xovs
HQ+Tup8DSxpTuJ0N7ybHFf1Rd3xMzEhbR4x0Y3AU1kc4sYJGdum/F9z9MbUiSdMjqfuw0GULUOPr
NylBfaXF01opDRU3n6wueCZaUbJshW+fnpGtDH+KOum+P/slqQbLSKGgEBgjOQw50x+kgp+QObOT
n+y0uM01QU+mXvAmOwOq6+kmRRClXVJ9wRzEWIAi0t7kSzqPPJKcmxC04RgzI73tzGkzlitbu61x
01PpZDyToMA4AbXCnN3rwe+WMka33WZNwakGgxoD1qxHvu7PgVEN/Rj/wF9nVU4R3h07bpmR9uKn
Bo65Gho/i6Bf7JIRRSfaMS4z0oTpyxPcZ1OX+IGcAn7N3kugaN1Ka7YWVbPypYGiQTrhRTKFaYNj
zEk/mmQD1w7YaI16LMyXgTLqRJxgRgiDGRsn1xtYgpcviJlXtJrll1UaURedthE9gLtF8ywhtmWB
wuh6dQzUAH9ya2wbJuWfuywdR0OciN1lLqUQPuUf9eRu9BjB/32zDZYR3S1wGw1s4Xm+Lx0Cqi9p
2pnCObzQEmO6umV+Gz5QLB2Dbzi4aqlBMMRTbvUT03ZO94f4mGJAYofyZ0Tw7A+TV0zpw49WhpTD
xnFuDK0b6G9ZUl+dBcZh01EZyBmxthiyW6+IsqBKWoh0wcmw2YeZ2rwv6Z+ozUMP2SzFys1yGAi3
BPLxujwz8unsi3z3yxwZ5yE/Nblarr54uKdzD+RU+9N+0ra741nXPQCoKdF2nwpfIGtwZXLcEWIo
pQATFfZpvmVNg4zLnmFuNqXyz88IfAihcNUoGOD/why35NGNMpLagyPsYmiFMFr1U44Qluzzmk3Q
TYEHyGuWFo7jQVP32YHM8ClpNXOMFLDgPXz2ozUGg+8cfh1rIn6aCMvddv8obnWSZTeaUHHXuAEg
HcOoM9mFC0KGM0WMO+pzx0XL771X3R5xftmJ63o3p1YeS/iVYDjSkqUeoX9Zi1yTXn3j+SDlgyFl
e9792kGcsmuaoytcKxwsqHGiz5aIL30pRIU5Z7nsRRbZcoZ7zrtGjAJ32bxRemk7C3EGfaVed9DJ
I5dsTfCfU2VBgehs09UMLJIaZaaIb+IKNFW70AqR3MYDpEEJa5qcUZ/QRpvN8kPyASz/wiKwKlYP
hwN1RKGbrynXwCcyWLjBI2v1M+HYrPSre928w7qsLgNj0QsiMaG5UMsBN551jH+Nri4FGCwjIUcI
mG9hvGmkTDJ0MLfY9a/1eSFvUt2RS4HkjOGxOoVagAJiUNpXP7P1BcvujYzqO+iTQguOYqY3p3Eg
koqhp/p1kGr6TEqZEcxv+TzP1PJOXaDtVymVm/xLfQPuywhvA3EhL6m2hO6eVXU032cMpDC/o6F4
2x1QgJBp5HbrXvKLmPMrwiWWwl2ZVe3YkBKugk8l8PUOIF6qeyNs0PEz4XSFiaAlq4ekToLo5JMl
CIL1mQJeQRcZPl/Kl64o9Yu4FTvhnknlozde0WLJx95xAjeLoW4pP4HLN+aX8DAjE2JRt8goC59r
+3l6zAEsn3zY71Osw9YHBSbBaKYZpFMPIiUe41oNor2tgawiqypqmew/VXmg7p5pMb0SPATNiXeA
IpNI53SsIT/qJyTVlBRrew+72cO59h6Fz/xEMq6M92s/M8ph1aq079IH9TFp2lODhQUuxsP6v9wY
ZrHxCr5Ip4P0u4WZaJY5u24ztxobyGc9dBqmmv4TNqNfTeWnzUjvVWT3KLMaTDOdMylgnZGuYtyy
s1bNQP8LrJsCglT5ZEd3r9tYrgXwe6G+JxggHDgIytVpVVQXvLcdEkgSVb+8JFjC2uD4Ce0giLN7
g+js09/KOKY4ZsIgoF4m25vii4ffyU7nU5tW+PS3VjoYNnjPiNHUU6BEHsHIhGtNdTLzGiq3H4wA
meIpmERoqO0yVtbx9Na0XJwJBWCuJWnRiFEYJKXblD7aj2gFOvHm7U9vs7M3aHFfIvo6ox/AUVEE
3ahZ7OmdSfbXANnU3eYsatbOD2LOVSe9dZE06oXP7iGrkjAqq9XzmEOoxwPZZhE0M2qmDKBYGbyB
Dj24Lk/A6e4sFIYHVpYtW3/aH/pLEopqBr/E+0xdkpeGpZUl0f4U+LXkJSJ9I7/royLez/LKnB8M
MD2WHO+lUEWNuAxhCK99XOTQ6H0jbY5OyCMdOnXm/xohPtl3INcPyJQeYkmusRpBT2PcyHoyhjBG
C81IfbismQZ1S0B0bWZ0+0DAMuQKQ1bnL6HwipAieu21wMowHy18cx27YnVUjpSqMGOGf8DOPEwH
ptmkrUDjBWVNi8xwsXnRMpB7KyPBUoR1Wg+pB7DOC8BW4w3xBxpF12+AGbdSLmv93tjd8H/ojtWi
WXJORYYQky0Suq/7e5w0CmIkryG9i2COwuGAWVRn0E2BuxqB/ULKxCTl4ePAayIg5OY9SXENho8B
DUisROnETnJH8Fzx/OOwJXKteXOOqmDp7kcIfvDudNhPEoo/r5mYmcjxSF00graauuk0NTPKbI9f
RxiZM4T/6mz5I9pGpbi2uJhP4l/ah7CQhBTTC2KFwEigcdnD9cpSlLDnCPBGMjPQKFK/QxWrm94p
t3XB2JRj5wwy3qYV6/3yzsVsgQ1BjZ3T6xg3Qk8QR2JwfrESFciNqkx4M02RdgBtCHwVyeL0lWkz
aT7iq9gpBcpRiL8ZlYT/2ZmGYEqDzSyHDEl6/4l+RTPvrfgoCp/MPH2zXpaISfGG3dWXwlbsjN2h
Oigm9HBy/1uwUm3rHwsubAzF3BGlCj0M1oaeF5SrN0+cvy/Zmi5NoNYxkL457hx3yOEluRP8G7aw
mCobdSNqNvlu0yKJQknPDRV7jibxopZbZQZ4Bkqdp1BrhdbHv5+kOYqnh50Bj+wAsI3zvYDvlHML
c2urrC6StSAEasoejfIDtwNqIhlAsut7X+1dqlBmD6r0nRarbDWfzm40hl6+K1k4PuOtYExPwB91
I4QsqFdCxCP44tWN/ZJB+JyZgVraTVi6rzGGEk019N5S7O0MhyQVdODyBVMpugM1RHTbJnlR2xBG
j2OhCqLVO6N5P3hGkz8j1K40JFRlSUmyUsPkje1lxCdZOkkIA6I+jBib3MT+4QdFrcBPhhR/ugFz
OiXR9x6yXmswkmKGqi3UCwcABSCeCQhPwdstWjyzXHzqfl34PERpQM7tD18NUy6ufa9T4W2doTl4
tIC27BD87jTMqeFMRXGB4p8sXJG+hwh7XZNjHV3UVA82Qz7RE0Qfsc+DhsmdNM7N6b6GOD/2VSR9
dgNRkMI5sJ+SYhMF25ayQjGi7X5YYs2QhKa3xslTSCZzuEx3o71URCdafgvZOqZ52ehd/hI5OHtG
3BX7djS2Tn7CE71szYjK803+bD7CkS1w21KDk6Jcwsfmer0Xi9wE5mXTpIqMJVVIIc9er/SduSWS
9h3iPqwMnyMDCdYJBqvQ9052Dz3H0ZyqdsojO85KSeWuwMDN+GopfSYkuteXxGHgd9udjT6WWUOf
83Q1AQgLQmr+wP78Z94XFtiwgMn5V5kcH6syWekWnbu7/xyn3oZdyMgMUZ29QmkFPpNvhDDyRgnE
KgVB/RysPnznGWdlCIU54PhNlAEqAKoSgbsOt8VuFrfkyJJA0tFqCuMpQqWIflQlRID4I25H1pE/
AT4IIZkUAJxgkgJL+6C+MsitN4xOEmotHraK8SrCeLPUJXU6L33ndET8bDKNDkkDs7VpeULNI9Ia
OlrFY/kUaXwxZbznJzGFk9M+DVDsBnj5WOKWGzRuAzze4dF051dxUzEW9W4T5SiKvXvKdS9h7R9H
gFQAOFvsMzx5LDpYzxPbFzksPNTt/kluJji1ZpHYNjhEoxdEmcK5qazn29V8iP2fo+Q9LF2Kvv7P
Akad2tJWeNSiqdKPTgHfHmnbMrERlGFJGBP8wimAjPStimTiCZPjzKQlchxPfJrdYJ6Fqin6/p53
aQGa2IM3qZ9PSzEDm0ZGkKM+41jco40/DWzWuTRDbm1hMJnHffMpqIPwrY9nWPHIdi6RlW97NACu
T2BDwlV96e7/4N3sO2CgG5BYrnM2ncRaajiXRH3+Uiy+xE06hLu1mz6CT2K8rJTgCfH6eRJNW1kU
9gm+Ts9I5vKYuXhHe+TNU7T/yip5wCeiMxelOSx0VhTqDZKago7Qp6MaDyNPayfVttf9p0OvmDIH
pwc/TAjLYPnRophwtFUJH4JAoIP+cjWCEl9ASZBh9qk9zeVWNmAZfs7MnJTBy8Jb6rb4KHb/BaJ2
rWeSpCdnsNmmVUU8oZgcVNfYDrY4QUpO5WZkK4HTc/a8OmWjsMMg29+zmPIVweB2JRmfXCfkSC5Z
fN3WRpNh2Q7mU70cll2Gf/MdkcGlTxQCsJD8/LBa1MyasufW05q7vdGH/nc+c5/fUBXVR6vY4VMy
AWgep2zjhGw3AzgTyxAndTg/sXA9FVvl/j83slGOpbdmhznDcY6xZAHqQ+anVDtFoUz3tOxCpIir
/pxrIVjc0FEYXf1yoVQ/JSRvbNSeyOU2cWCT7uqLpWwERmEflBscpEFdTH0u49fxcg0J5psW+Dzz
HW3NqvT9DLPA6QUgGOgSnwyVqDAodHKxadvYoee0gEiTH8uszIEfTFiXLyTaokvWIrOqHwx0leqk
smvs4QDXzcU17pNSpvaCmIEh+Ahky7BNpg9BO2sPj4DQdnt1CFCbQgCRVdHHt/RityXwScIUaCcw
lTSeVKRFcSDOqasenElNis/SUI9lJPqUTDMpuRJuXdJMyHiudtdd7/2O2TdBfQ7KZL5/rOwS1ZCP
MkB8Pt/hdRd8m0Igx7vOV3+pA0pS5mhoZOsDuKEeFs9CWALNc8aPCFoaVVUpJn/zkL4NzpAUKrmb
i24AJqXL99ow+bnM6zHtXWO3UNFehptA7RNtV3H98xdSNyWRDE+9/ohThawbPH1BFXMvTJLGIH5n
ZjIZUA73peEbXHyrwwlFf4IglAw2WOMR0gb8v78cs0aMb6H2o7lDPR1kx5j2+9ugjdLedy10w6yu
KXuVB8xzbx538ffJi9z8HnHp7pS07OiH9Fx9KFztDHBDj7YP7irPx9Xhaa0q+FpN4DREqbyC1JEk
aXArBznt3e29qaAqbQk11VW+zLEgW8e+78N30W3J3FX8bPwaaQwcwpMSiK1ESc2gnsA7E6XJmUiK
ODFQfjcZBdBAsFp38unWsyeuPzxyhYr4IeGBUGUII4jwgLNTp7zCsOICc4PGnIdChxzW5eTjM9dI
vzbavwP7vs819uxafvLXHXaKiOysSeFMuhp23WnRYZ5TavpPGebQCJ9bgE/lo9pqvN+/2OpKi48U
v88amZDbiRcvWGcva3yGFoMQufU6D/aNhv44RHwEIoMklc/ZMGGHiZbPJBUVlfsNxnAM8UyDJP1t
YpHmo3mRjLw8Ih2fWu6SI2VdWpkl4BDIQUEJhj/RzzjVkd5o0RzDUw1fFgWP0bv3r4c1ZUswxdMz
RIOubwAa5G6UeK3jEWVZcl6Gx9H5I3gRWbi5ndW0r4XEb3PNt3OpPeP3A0AaFCW4KInvOAt/Nc5L
nSdemNziT1Qke0pHAbrrhKmKYU/Leqje+p4PkUZ3dCRn490CtrqrNgRDNO4JHWWO1yrar7UJ5FAe
rPHMtBywK6E5jHB9Zc+ajpU+C0xOxNKVC3RwqmPgg7UVahmr5pTeyKAFMDfgEwMXcf8D0Sley5/8
nCzN5qZKRk4vmcaAgZTDd98/ZUw9aQ55zlgkEuROTl7A3OorZJWHqe4YBYzHKND962EuWQK67EFP
OPr+VmH3kwkqUqZUY3SS8CngmODdi3+5+kbQH5IKAI3TpFwrXzxZLdGTwRHlNZlBdrtjEynaVQXY
vNAKnTaeHN2WaT3iV7YvQdn19sXb2rDCajPoGFF5onji+Ufl1v7LjeXKNzPCNAWRybK8gD2GmHlB
jXn6aF8IlIHtIWf11mpusRWqUz7K9X/r6yNZqqZwcYvIHabodJnzwZBbTK5qKxg2nzb97v0pzvev
yg5F20xIe2ECC03Gz1toFVIS+LxBzeCwVssyYMEf+bTFVLScuZQcReXdaQwzAefr8TYRZhLiL3o+
vpltkoRVqWfiSbg/RXVbNcsk0QT8f1c5MqSHHhdZ4HCi7xk39E9NgTIV+ZUXCIp8YUT2jLBCihBZ
6PT04qVf4p0zJ1Lwt7OdchH/W/QNoLDNar9vLz4+OTxcFZ1G61W+TOSVdVexnARai8rKx9rC8F/u
jXvprzlKFaSgJUiMgrus68z63VhYZdinL64Qlgwov7YqNw9fPDLM3cljqzuLfGzhery8FYF2f8zX
0Y1iL/G21L/74ijBCPL/atyH6YhXxZmGR7wurwF55M22eykDxa7DVzFe9vy7qiF4BvSXV700HLBq
B525wY0uyh7GPtNua4ToSlS1F2ZEs9McYPCfMFrOXRJRDte+GV8zpujiGzIz9fGNzeAA08xrbGO+
mDU68E6ge/htsR1LD61sCIJeOT9Tv2VAMTzLpwVu//yITwaI8ay3SNhUQLlIGheKIg4QLHr/Knit
5QyQHw5DXmZsG4nARP169EilYeUoecoUDJIAFaP6VpPfjNzzSx4gjhmKnn1gE/f/7SdLNcGABk2V
rPLFloJZN8iqHXntykXO1lyHV1ifk+KS2L6KtsfldyUq3LT24fe1qk1Raqv6A5eApS8ZXeqPegh8
jd0qntDSG2QavBziXIkvB3DCWdonnzb5Wk6LS5Kfz05ndYYAXOAvIVbc5G11XpfIwq1joCpLbsr0
CTwP9LCAKnQbUmtaLF1Wk3TINC/mFdnxHQEFF3b/xpH7Kwe8SXXLgKy5ewDWGmknCW0hjFIgb/pi
HygFjtQdJN1fBNg3Yd+NR00WQdMeUJLK2dKzL34rRJBKQ/K5bwsZ5ytN06lrRTutLDtvJZhDuFTB
TdXdKF/hnYX7ff1BqpJ99OiykE6XaJZzExa1eU0Tczxw0MLgHzmKWCo3PlGk42r+12CyYlL8r71o
0NJNejKAOf+6TfduYXi0FL2XbPR2P8vASGHGfEkfgi3po34W/VbuOmP2sq0xvBIHl+twZ/kfXkL+
i0JRbneOxJ3uf4rDgyaKk+feNwJuUzsa7/Fsr7ynSxVp2bWuxWOA0hhcBjWqy15o83jjUHxI00VI
/Em0cpGDFmZUUSgrJ37BrIw5O33sWa7ylbcuH7o31MttAondkyOQXdD4dXwR1HDBdsVVCSpvQrBE
gdO//tzRWZ9hNHzkGTuZTe5vLbFFeUyXeYmmiCrlRXxu/Igo39Fro6ewZz/tFf/A5c07FIOA2EpW
L5FT0GBhMLgtyib81OfC5NF8CuHc1bpTJmu/TN7VXOEuswGQxySH0coXU098EX2yDPb8tXRGOmdh
aOa6jGdKwDH6FdjIWPyIW7gQ/DWN0FA0yWXmMgpw+m/0YSAP9xZqwZprsVV6kaLObrdl0voAY3y9
jECVSiL2y85fQdJP/VgUZkuBWEiqVL+IBUDI5p2txskb0S/eb0JlecYff0FyQPjOJJl87WcRA+66
o95/BnfrqWFuMx+iivFwGX5MeZz6TilvH2BxVRXZBibzLw/kZkZ8p/zd9KmDqMbMIOWpbriIR+/5
Zjsb18ewxPt3vU08/7DDLhIiSp1nw9w4r6nugtCO86yLXiAPEwsHLxaBNzSOQMng6fCOksR4U6JF
iXUaM4EWG/92jbPf/cYz1uo4lhTiAwOxr/2Dy4+iN4Hd9uPuHQLm0PLjiZqSEMHeySJFzXBRNznW
o8djyijsOhSTh1DNoDKwnEoEHfKs4px5vJ5yFewq2FgLb13owF0PG72nJf3gyiVYTWAOSPusjD7S
5vBf3+exU3SniU4IBELOxrVkB7Nh5yUqm7RHXYFFnqavpJpYnlVRIqPd+/tlYn7mGs8B5r3WL6gB
TR/gg4mOlQhIv7rqJ9az0h4Rxqk51LpRokyrER1KpuVwa5U2KhMY00y/SBrIFmuFgnHQ74ju/wGf
7dFhPfhMVjsvXtRA7N9bR3MrZNzegh7CbvVRvA1v+zqahXLf+eNtwTEtbgmt2KPgUGsjFWyFgfdB
9ZzGT2sOHWNReuS8ccJbXLaoDh2ENPl9BdHpkU4YmlahB135Cw1F2sFAbULHnXcN+vJEGzFWNClc
rQUMsPJovb8sXZ9J7nQQ0ryV7m3QWRd9ndi0tHRM5LeBLA8Z/KvpRL0PowUtDH/J4FuiA96sEfRv
rLkZLFn2NGlxaNRlcnlkQzA7gjhFKuK53Tt28WZMjV326TZmSxhFPIyqEASmRWLbK8YaaRa47dVV
JqXM+JH9QZJ8DsnXqzJ3zGESE3063UC4HgCH2LOu2xxQqDl+1TJSRgs4F2TNbeuC9iYFf2ZYHI4I
QMkChGNliFGiRCaZuzCTSY0vwVkNY6iwIPHdANEv1gNkOHDWZwhfkrYelb9md9vMfxABNeFvGHiP
yrW9Mxgc2mLQsGjy9/W5614h9u/1Pe6qxGiT5eXB+vTaRbxeh3erc2PwwxENU/xH6CaxU1jF7C9Z
oCe4TJ2gwVhzREn3OGtjthfqzHl/NMy4+z8s0sVnbKt1m83Xs1yB3Uv2H59R1mMJFJVoSLR0oq6s
e4IyjcjxIbxCPfnySihA6GVDMIedqFeCSYp3vxAQKf2Y1eZ7Qy4DiTObZ5DeehzVtcv+BdMEKqXg
dn2UcKqlGthHlfG4w1tlY2ERjMHL8I09h+0MAiP/ItmklYKc/1nSQd+oWfYUtHvYYa5YCA3D6Xzu
N8VS9ciNz7oFa7mI/fvPqiSv4lblz2gnuo9ahZ7q+GY0jUPaLxJlgpLVWADhOW4Ow8LsY8pY5OLq
5eCBpPfZsf1457Ijap0/o+pN82Ph3/lcyQjUjKiROhesRy62WhL++K8mvtpY1NK7L8o02eCB5OXp
K0ReYEsGTjwsa3giZh/PxWX5V7TwR5T5z7dUdn5BGfUpjCNxzF0HP4xzCr6gjdguR45RqSuvxo9L
muV2p+vh3EvaDUTfiOGgh/Y8eIwmkTeGz8BKbUc1C0uQnr+DRMWMnwmSaAQtLDB6+shHog7bXRbn
PjUIsdH18b0QLrrrbEG4WJXHCVcOXTvwGRAfXuyUVhzodtY0V0zU3PmPuzycUf4PH0BjUjqAv9ZH
q+WhdtnKGNVqNFDBTM7K21aIRT9jWNwmZe3HoDEA5rIzWjHzH6RWNtg9G94PpBu96m4DehdblMEa
6IkFXwNCfUl/OMAcPQR1TvP/2eucAc0pKInmiTnsIdF5jzpZuHKMrhpu5r9au3o8GFq91mz/hvi3
FqCGN8vO2W8XB3QV3kFb+kUZnWpHKalyipHYNeXCpWYSYLhcX817TAZu5QinUm0fiPYN62bpDyVd
XvnAIS76VoZlAL2uClsquFjSIQq0x21/OH5qaGoG5bQY40/90sr+Zfez2aXz+Xw0zudqduOCmbyj
ZwnIwSFM4KS2Nbc4EYx8/Vp6R4USfLFOs6xEG4IWl8eEsI2x2XNrPt8EKisAG5NlGCejjrfbfzza
UI2I1zVQJGm/frDB2bnBb7ymO4e3cEfxQVYj9bLOqObe2sKpUzlqb8mQTIBrWD1ntVd8OROBT9Rh
u+aHQGua6uEV3k7Z+9SYdHfIoonh+M3Z/H2XF77lRLJ7EGzm/VZW+UpyuGtcjKnHO4C/5dKQz3Iu
pTIRqqKKtzqg6YvRVxvZxrYLJ7g2jQWViBEHbNG4qdKbunyDQ+qCcFGLYa+sx8lavSXykFVn0Ys3
JeL9+SU2a1EtflXL6qibINDKDhDBqWcFdfbVitGnRZzAGppG/MWEZyTKmYQp+Q8hDs9o+2TdT0cz
D5vPofm7cCFRGN+beg3WIu8OO98NEWiFs1RXdU3lgGVFx/NOaM0OSVAWZp0HXUP83lElmpQv2dcj
v++APLSnQiLTKrA598CRUOduIU4RVgaKut7W98znNS/QYrXTm4vI+TR4ckha/EoN1aWmhTGtl95k
LSXomxP9dGG4pATkNhi8FLezx8ZH439ydB7a57E6+gEHwCGkYgDwijrFQuOJdkCRyB/CeqYfZG7L
o5UZKN78L9R5/h4zThbTTbS1cSBPceq9FygAhtUmxit/iLCniPv5P113URA9ZH1atIuM7pXzVU2d
yu1WIRf7U+4oePzFOW8kdCQsQ90/B1lVkSye3QCvYG44vD8OO1hpKXooIfjqgdojxm3LOFh2xcVV
ICBa5s57NZjq/2c5fWQk33y6cmCZHShEVbjpZUpjZlZ4jv2ISnL3SBaVtZXevfreJtXy0gKdAQT3
1TST1djN2X4hovxCwn8xKwXKe+sBmCWEeUWlvG3EO2unmnNbGI5wQTG9/E64HkgWAoDOa9tGZ29K
StyjI/uSONrFMF1IXzchu0Laz2du2QTbYIU4pWXRpiDfVLu4lg7Ffu0zxevI7YlQSS1Hhio9zJKn
88vqwvnaNdTzGKv3U9LzTJG/DK96OvTKC3sfV1Mu6WMzYaIrZLb8HIpeQ1G2C5cBVitcFTYVD8Ds
DoCCNcOSaG6539dI4BOdMWbUKn4++APInyDCrSpWfyBMQcM7us9ui59nTytPNrtVLfQ+6nvAF5Im
XyMUt9AAAuojw3PlzhcqBwlbo7xPKfr6m0XXL5c435w9E81Bi0ScUCGtTq4TKjlASyg20whp44BA
i0W4dOWakk9os4bvQazDD0LpJtPjnC5niO0vA6IacB+gscIKwbf/GcgbCKgKM+Oc/B3VBDr/cXrS
MVxV1Tfz8UTik9ZiclOnVKtdJ9td9m/nyLTFm8/7JBAPcVjquZancRB9GWnOj51To3HtrwRvQrVS
LkU/kialK6rLexzHUzoSFYI/5qwOF/uEV4yKlCXXRQhlJcP5EV20u6T0PgwVjOpJNhdOUcttTVlr
Bnd51jdwG1kxeI4ms1xqUENZvWJyVtm63eNyLz6ZIKt/HSCBSy214PlT0rYvt8vE6oC4hnZD9dJQ
YuDJzeRki4qUEG7dApM5FOCDhgrsaRDGL1lQ+XgOZsKFdCi2Z9jGGQBt8EL6Grof6mxiG/tO+S22
1nfnFT0bAAbdKc9dAUBSmKwzISvD74fSWg33yMlZlnuYWPPdWe8U4eA/E8YO0AzFVrjDxYH19stu
f9bTTL5m1Zl/ABTmHUYU7RT2r63w5WzDHY7BbUuw06EFSPqRPNHYktOJ0Jq7jOoSp5bqpehvEcPS
2P5oOmqHBZv1DNcxQpHFCDWpW+CUchZCxEBC4gm29MKEetPxOu9JbChESF1+gIFrFyhjis+MO/Ry
d4hwjX+gX3KyTlvXAlIn/ACWzsbAcI/id8emE8perWt+s0ALytjsc3RBJZ5b99zkFXhNcbm+fMwC
BhYOM0jw2wdOzz6OH4dSckXkDNNmJpg0/rWB0Iar81swQFEI4IDMjLfkA6cdqhabeg57QpvZJbkf
x1/nAMU5FzTSJpUC9LtTHFvxzEBRvVucAEmiCY4NmH6xP02jDM7OsaD0ByhOih6tCUDG1sFRJg7y
tKKJaYVG0q+arUUjtoFW3uWna2Wyln26Xw+MNb8V0eBMF45DOx3t67U66ZJg1BTlL1nyFHTF/DiK
wMdp933oAMuRMf5hSMH6+xrgOaVybJm0VBXRhlhdCbcXQ/O9VeJLGME6kRh0CO/k01QWdVry83XO
km+xjvDG/9XNbKs+/EPJw0DHSAUG4gZs7zoL4hvki1xyCIvTP9lkSBj6VkxH74QxiXqZtEXrhmiW
16yqHCO+/O2Wy43Xa1S1zVRObsm26Su6zeUiJtru0V1MzHD4jpi2tvuM7YAOxJRmgnukbQv1YEEq
r0dk3r/m9cslgasWfNDvs8NZfnJHE9PoiYv9kN1JGbWPee37JqrSnxR3X5JTXErNo0w01H8rZ+zz
IJ3i367MKmUupk8iPpVGU12IU6R5kL8dQRfUJ3aZElFbydfZBcMXEcCoHRAbBJT8KcwOFYOQNuEu
d/7sMXkwzkqa7BZcqiQp/F0kDXsS6za6POWkH6Jr/vyLRreanAl97C+R+iNLSbJw37g7pnvJciTU
a1WRaNKEOSnoLiFhQtC9Iv1sVXUlRAz/YZ7QEkBneyCrUBCzDHaBDF0J3F6s5q99+RvTRGJyUc9/
mxyLFy6zpLK9eisvsw8amTTs+mxdT++JJBI0SB5jHdYnqyGBaOMD3jVJtPTiGMgtVd7xOVnWRcoU
+76g/2zOD1q6GTpJgUJnpUevtzYuJ1vostrQ8n8IPif9ogKZbp3xfLKMSMrARMJAOFNW2CFhCIoz
+cRoGd9LXXIibDiLv17HE76PSLrjdXDLOtg9LEkK77KH1NjjBJ1gvFUYsmeNbs8nCo79Hf/51HTF
qGCLjfIjczOQO+BPmiaGp4knNInRZdD2crfa7uNcVfopBZAschmJHClieEoxAP10NoCuEr2x59r5
094eP8YQ0Fqr739jyms6q1U0pTCpI1lRr3TbCt5qB1dzH3EPBxhEwCY7tcqv2/DSETWzLo/00ug1
nsC6OF81f3CdRT8484HjnFJ98Z5GV4ibmlnJv1uGsEBM4mbB9AHV64kcjAg7NqYgz7DpA0zUHoQw
sBtHvio/0m7KwCwg9FlQJyBT62QTCTTFJXIBvmuH3lX2xP6SXbr8krq9LOlz2pWxkIYM7CkrfDIr
wKTxV+QtQCO6Pq3bbWPgNPpZDWFFq8WVl/sPOgJwyfK5DCxa9zRA8+b4oOZ7a07o42R+16WsgUGx
6P0pqVcutd7mKL1a9Mjf1/p79So1zx6xHOZTNV/Pwkrs+36eLdB6uRVs+FjkEnTkzKT2Euj+BQnf
Y/qRf2GGpeiee5UQwYR8qwJBZKGOgoUOq/2CiGIgZFW+NrqfKMln+uldvgtcZ8aDKZQKxA2HtAsS
cf5FT34kxIgfkuv6hleCKH7XDtE37YZkkaUnpHKEznGJIXbAWasWmHuIO/vcn1Xdu4pvzyZ8zBt9
NYDwx8dgBex2+qk79CmiDtMHg/EmchxoFirpi7nL238NXGsOFEqSlO+G10HwbiOwj5i0qxCRoZaQ
hRaWQAdep1wzs08CH4ArJ199O0KuL7BGfV1QcrV8/hvk7pmRRAjCCZDKmwqILaXEjCZn7BoCx8IM
rpzAxYSfUFvYHBxiup4CBu/3sUstQ6ny00THzm/5ruGtGNnIUzKBlQ+N5nX9nbiCtboazOgNkke3
pwl5cAEp+K838dMXAhZnL5w3hHICblvA+wlN6ddMqZLtXbN/KEn/r2n/adwyxxn3FqMMZpdNn4mw
xRxExHM69FRXfZThGi7J3qHVqL5SjsEefymIE+dOdwfJmlZH+EWNYCgwGfoSwqOFxP/u2azc+AWD
fT97NGS0rwPcLub5nEedI6xDKJXbiT1PlpB/R4Uyk/mrmmC9FnEkmE9l+WdftPpyCrfEJIBCM1Ab
y0obxozskrA/bw/dOuXYWb8RW2VfLvL3oiA1ZxL2EEAQ/TJAinufAhC8jyrQJpwpDLI9eTX7isXc
TfZWqrssfPPP8MO9HvC280bvGWbqOB2yT9q/P1z1TkeHAzoibwomLrAOC3dJzJpEhd2mX1LEuaJt
HYv/SjNJwPqXbrpfaX+jxvBeeHYYlWs4wAQ6j2FoHcYDcO6GZRzuUxq2vrAGe9pRVhkiLMftWx40
8ZfDjVybuZnpjCLejFm3ajvDAhZQeyY4v0gLOJZIkzJY4CmmC3A2pucCk6YLsfOtNSZ8S94/Xsva
FyJKDetiVzCOOV3o4kDJ2v9NgR5ufb2VtgygrdHsw2kGocRUyByH2asoCSs+z+egYUYso6kqc2mt
5KvDR3TLnUyN2r1okLZX4WacrmZBELXPgeJrRyoS9hb+QV+5983slujOpcbwHjbOnHELD3Lb5sV0
ATt3od2StGTHzgT0v3XMVDjkdgJ3wo/o6QkwF0KlJvG/AzHiCacJe7E4xiJqmjQE4oLO70vLKj1N
HPXVYh2vPO8gWNXr0OHS4sgMq2mJwobPK11usvXI6bXfflwk/aqgn/YRwdx3SA8Ss8ikR3vTy3kK
ct9BVJ/OfEiHx6Je24lkR36bynxvV8FYrrnzO7Cqv79CuIBk+urU5C6VZdGdJVh5P0tZ1Y2XhCMA
vY7n7iJE16mNXnsDrLFhQgh7hK/G2TDpRAaqabRomRr/JSo1eePqtLx510qNWj8xlCueKhwcDluh
NTMClBPeqw2EbkhVGH1Cuu9PEVL184zaFQvT7E7hBDqKozBgNVVGAhjZaEFeS+1htYbdOJQxlLa/
rHxdxtI+soRAV3H+zS5+k0Wbjn9t3ALu+9jgtelz94zhbn+iDlAxe4WrMNXTtdRVwRH1airp6QYe
EbeQpvlp7xwGfZSFTmlToi4qoU9hKcY29NzksNuU02KoJAwgNQ4D1QnMdlbTdB6PpKk0BqwbmvAi
vI7SRZAOyjbRcgmWYM2zgYCfcnrJvAuZcAzDGugMTI/Qf1uvN0x224ORsq7eFjQf+1ACIvyhgh7a
bauzgGKPZytmD4VktSxONICUGl6cwwXa5rJVBvmWNV1nfimSPsO21ZBqQzQ2pZ0MxOVCtkzjoyAH
vtY4xooQNzWaSPQQdizecBSU2W3xKJS+7vbelWTK42c8v7OKbC43+lL/MlkKWYefrWbQFDWeq1+H
qogUCkGRfyCNICJfiRDre4dGxBPaSunJhOAULBsxK7KdUCdLXoNpYesD2ZfaVda2KnumcSO4FBOT
7R9cYUjiLG8xRdK1JcWZ2YX8o0Mh8CFmbqE0XBC0BedXBKgjrhwrOLWbogXBrPRI+NqH14nXRhbt
2wAIgA11TnUDBV4W53Mvr1KYMPMouGdOlZGx911esFr5GwB/hJk6rmd8TRjexWW0lF9hVUV1/M72
0TwLv1+AUrbT0M8H/myDZ3XuNi+jNxQbtBWA7yDhWzuJaGwcHsRV0gKLX9GlJEjFcX0Xim+4iRsS
k4pkHXIDb0ZUBGLmVZtyP1xd2CXIXnl9dshsplHDwUrsgDGCevkQ6I8218OH8TKBWIdhz3z+GFEQ
5qxYx0JQ7bAREv/ttKqhw3DtvxBaVf9mEEg8YZx2hYX6SmGqtibCls436KKNgHm9Zrfyd1HJKGIg
4HsL0GmULdXQXG1FjU2VTtePMrQjieYawyJybWDgBJGjmxBjl9VYeX9hB/B4pvPbHhhQHWlA2r6J
JJo+XaFolIbIbSF7xLMtdx8W/lAqnlws00QDsVm6pHn/alsSYGTE0dxpEgEnaBsNlcY4sVy+rhHR
j593+jcXcsjRxB880RWxqH2CT7oCc9NWpKePNBbWEdcYM6WZLrPENJGJW06NF/GJFrezYUWxFWdL
a5lsFpcojl3V3ANbDxW0zqsMLwkhEWyNZggdQYwiKFWcTpWkZS5zpXOKnWt0zowA+z/0lgzjt3nM
cUdjbdgPR7/ksa+ASmV1fMn/pPQSYHNLofyl20s9Ph2vN3J8Z8oidsIMlatlHRxC6eYYj50AE6ei
zfwlfNznnKg/ASAMyBC6Jsa9+dL1ColE50iqRLZEITsX+ldsgbdsLu5a8QS9RwVkz5L5F4ap1mt1
hgg3g3mgbz3ofX8rrOhIXdweb1veYbpPHfxGy1sKJogx8QP9pdXNvDMGzRD7P6GYNXbgN0SsdnY0
9Q7S6j3IRB1DcLv9rxoreIsCBGXrvxodaf6lQM8A5pHICWzRl5nYkJTdhqUI7v9YSv9IvRtv7CE4
VIqObjhS5uliNEqn9GQD8LjYt7f3bKyo+IuvqEZT0wHqS6q1BRTvDRWlXHxWs9tCKVaEz0ya2pUm
rifM6cYwZ6FZlaIEsm+I2yQwCXmzVN++T3z04iJuvqdMB4MDNHgS0zAvnHlV75IY3juiETNI0BVz
QR1hxnDCBwHR5Udpzr3zXNlVz6GsLnVXYI+yTOVpubhPWHeEqdu3Q9AIsUiiwxnTzoV4WxZjq/y4
HeQubOES2ajPKmrWbNhJV/jNcLgEs4/JTTd6MInr6bpBbkkQQo+76GVVw78TIYeysCjsdnenQeSl
WnanBegAMpI3Nro3rpsyIv/fF6+SIVFbFF3MXrk9eG9qLVB0AHst8/rgBz3nhd13VbXXhOf/LGQC
lggmYJvw1s2PJXKO19T69ZlBG2ko2si54UIR84kb0Kl5D+hbiHxhJSj0jlR4lz0DUFIJSecsRZrH
Sdbu0Fus5b5LxRYyBACUB3BRMMMR9GIC9R1neLHnOQ+LfQSH58i4WQXIcqZJmW4NsliLm5bPX83+
JH5diSbfryj7nxLi6ztNccdwV1Hrgn1CQUmWFWnb1slmhANifnson84+IztmVHnluzw5tprvj6ST
9KW2YUDoWo/VdvlQ0vUuLkgZVGIvdrPoUWJPGbWBBSWnoj9r9x7TI0KRVMMvLlXfOP5uqpUdChpq
rXVuemt47s2ijECozkNpn2FIAm1oBatJHEi7WGbpFuDoKlAFPGiJMUlv8g49+XfHQAg3tRbU7z1+
janEXxRWVdwCZrMhj4Yh2XTSxYPBEM949GRmy57EFpYpzHjsoxWMJw5MUQP0rjC2PvESLKJ+RSa8
h0qfFjzmsl/RXRadja79OMXBDQgTqlnu5OFhTAwv8qzwrEZoAvB2Ljd5lnvfWAt8sGc3ciOtX21c
8Wh3zN3RTugUR5zfUjRY8qAa8iSU4XAA6xZYxrgNqobjwNXXAkGiNljIhtlr+ghF8gg0rWJ7eXyy
whUIPjikUflDzxPL38JP19P/OHZDk9RuNHIXLLBf7KxR5Qei/E1zIDlAWYduiCaIdU73oZyiW5pD
UOfS3nWUnChwgnL03VCSN3yWi2Ubbrc+rJQlGSq+IoKqU774AVz2+QLDGlUnExuSntEA1M+yDy45
KxASv2kiCgiTaRk8ITBED6HIsw6FLPw3UudRP3cmHuY4nr8kmqW47bZQAaVIKktONdltVyIjD4Xz
z40Z0YSb4+/4Ku4mlAK1qzuJcfMrdKaR5zVyZl5P8Ynf1Ypc0Pqa6X34uoQnG5Ur3COXunqc5uzX
37TaKAZ9L4zuX73jfyQ+xlbxqz1+RV4uHnIgYsrEnF0RuxkB3Jcv3Y7puecSdpByqC4eC0u+w253
CIbP4SB8sygdWGc22ovmlutRbc6fhCAQFAyNc+1NbNrkJDGT3zD/W+Lb1lybooSOiDRX6zl/CVEp
E9PtK3/3HyKGvJN1FoOJP0HBg2mZ3vZ7rbW/kW004ufcC7GoyridjPlSLmwKnOB3ggMiM62MQuE9
/7QkGMFSijZTITv1oXSMN+/0ZilPnycHAzIgh2bYAZlylccQjtmS9Yxgt6iOk5263jip0aOAspF0
nVboHZCyimhwlK0femcBTjoIOnJ0R0CabT3x3jBZzzvAE8yngYVxvcdFDx5soWDE8J5sTvlpc2S2
NOXoFeQ+Nlm09fUV2eWztrYVfLfEpfiod2K5HupcEBXHVP/m0uqQRle/JVPDS/nJZqHNC2MrWL+O
6Zfpvz8i3BtO1sQVI4Imb5nbKLnG5iIqUihl5KLnvquo26qHnSIzHfc3OjQiqHni5hbVVuI7sJT5
mvqiZTG3dwGG57hdDxFUponLiKnKZvdx2hE0NDOodxBV2T2PkS6TBe8F03quONseMWIn0SEx/ncY
n2AHpR1IiIFX+zOSoCvK+YzLrWLFkQZDWFAMB3cDU4NSv7FxN2WsP+HSqJQp+9jINV+hpOBk8QXR
o4JDV0EJIWiwV2BGK4oJSc9PltWnNj7KxND3lUc/fVYMiXJFd9bx/rNH7zmDIrr7a4XzYokQoZPL
LA63prz7URA1C6P2u2E3TTludV+OZX8cdKfIWy8s6HZu7oFmS4mgxHnt5Rrz5PyqKfURhZ0wEigL
BjXg9p4QbhBrD3KwcgAvCpdiGLGqwI+tPqIjDaTS64WW2NWBgzLVJJF0RyIh/fzjr9LBbItY7Bpv
jZ1T5WX6QG7Iu5EzFdFKezOiI7oelOo5oe3TDh7ikSoXagtBFgqN25kVCfpiNSuIy95OUlUXl2oT
zCBLKM4AASnGswENAsC5aqSQjPn5QIDh1rIPuGBLauw/lMpLR9Mw8scvLhf7Kx5dQcrwOkvCuM/W
txo3jibsnxUV3drAmF0tUCtGQ99hN9pITsBztzmo14l4fqhLMvGad0h/ocoLsl8s8AiSYDj/tf9/
lBZMU2iCTlXwsrQZ7XffP1gfz3W5jKGY8uDCc9cTePvbIfU1tNnKc9VvVI/UuzVaFKD/gzJ2IQ23
39NNj9LMsJTDydx4VRy1DY7i9k7Y4aVWlGa1dHQuGbPMuW/MAQDfLM+9WpdiPFX1ioSmOLP3A0Jp
QP/I0DclL0m5wUQ9kQ9OPpWhn7eRZWnjI5lDzS/xZi46WMk6KrArLNt6aolSqjFwodd5qJW6EZEs
W1EgkvjkDT0cs9fV1b1YkIT+xwXY1+2YZj5mtR6P3h7GBxz+ihEXCKMZbZbSTKQET3ruitbjwjOL
Ni6j9305rnY5Fkca7jYhOMp+cae7owPctGY0f452RlFVIaVPttqlVHK7Tr57b0sNnxUWKPpafqBX
UHcHSSZ3sZmHA5ZiPHRhniLb0XU66svPvntpA0uR1T/2RpPckUxyJu4GNAx9c3z9JxMLf5efO8He
GGJ0mmVPeaItRLj9XTCt2/2d3XBbweEZTzppbJvMCh/1HIBS5VWB8YjsCX18hYdkQgWtHu4SpxCS
Iz4dytPU51JdzEFjJJSdeJCCcJus6Ko8eEcYIMjZaoAcgR12mk2z5gPKcBdEXqgXJp8nHoRC0MLJ
XL3mlW7FD1Ii58paEJ6hwJrKlIAkaPCwr/d7a6C4o2urZKXYAa5Ueb3h/IaQGK3EdoDw4zomgB1X
ZQyLTt7R6qo3Tw5GPNrl6YfinNCA3mvsWjebOrxnKtfqy7BerKpegBw8ffi2hAOQKGiO0C6Z4Rce
qTXdf1mmctRFZrBUtFTMdLb53bsOmHHaRJZJnt84noFWAVLETCUg6xSvectjEbz0JZKHIp+1fViq
mBe10AxEPR5br+jPlvFLK0hGEZpc2ufvpgWu3I2yQdf1PMI6QwNHjRxU8r5nUMHgP7jkqRq7aLLn
D6zeWNJjpm3fsAit1SYUTpQkY3td+31gFdvKhqqCfQnQU5rFeqtLVYT3jeD89P7ELY41Ywbjhfcx
eakMO+118HY4udYIWhE+KCGRiUAmrM2jcOK59RTEft6cZ7UlBNQZ+GCDMtUiVL7RQTSKnsdkOYUl
VZdCmcRfsQ25Ptllm90imM/egi5f217Lg+Xxw2vS/Whw0pOzemnr9I0z/7GhEyMbZ+lEpOY0GDF2
31uN4RUcmJ8fK/t7tH1bhEQsij5g8Hqt1jVuFIO6aTkxnmDsTH/EaXf2Pj8UWojLu1rhEaD32DDH
ZRv2H4m9AIel8SpX2C/pqg9u9lOvvkyLcz1CWS4B+2LZ2Vg8oaU+PfKqMzcNcCAc7iuW2Igni1BI
zNpCPtLbecxFQxiYsNaL1b39/QLxQxSL9aCPy1/M66poOhblEqYFG/cNc4L7qkKgnzRgsSbF+W8V
JFokxdWoakPd3FnkdjyQxm1JERS7bc9GwecNeimkpKHZH0UnXuk+g49giD16aafzt7fOkGZBn/q3
GtjBInNjh53uaeaZ0qCqqhlX94Fbn4EpQSUo6WSBHuLnCkYgpmVh4ZXhZ0aeEAW0ogtpWBZQ9COs
9TcJgDQ3an/Q7zp8eiiPIaFR2cX+1r7Hret9nvF+rOdAybg+I7poRFzhrTOqr3VRM3eTDRKwvF3A
WFYG7XY2h4xRiKHnw+N+VZteeRzcZ53xf6FTDJ0CV4q6ogwOKUZgtXeUeXAc4HmrShLgh1llTeXr
8jBCzAwtzRvDXHi5T9y0QGuWgcmsXgDUoyBqvCrJJEO2FALMRYlGqULucv+VSSyquDZ5pEh+FWRK
7tsRptxS62N0aphBkV3S5YEPjq+qqbNj2kyPsvGtMQRSIMRN/jraM9GeBh9W5yQunqbnLJElTXkc
IuKSdmxbKyFjwVg3ms/l+/krJGP5imIvhIPYsuhhjaopSZagZdDDR9wVi8XpiQ1wkFC8atH5uYfI
F+TTlf0bCJn3N53TrQ6kJWEjBNHbyGa5w8OVne+2vSFyAJ5rU2jZofaSORTI0uR84T5mdXhWlNJ/
pKiS+NMcNJvxD+2GKCZz7CRyl6lVkhPX5AoCsji9ciHcCUezeHdq3aAdidaJr7rj1Q5T4f85IGdG
E1OgxF0Wp/31uqSrLSSWMdfe4jZbJuTVm3H0JBNYRVdF9I6i2Mqf0dJf1J4ILB7vZ6NI91gcrCTL
7tGMwhO2JOkaRQftNiV18aMjx0P7lnCkLhbue1GyPGJoMY9rP4koj/GDFkuXbx9v6TYfdVCTrKfu
qwPPe8FLJjX+DkEK0gaUGN+1p6I2li5qQT1MO/MPonpeMNGrm9dOgwWxMbGZSV0v2LlDNJhOYe5c
cMzF8WseqJrsvdhYdcSDn09mBxMhF+eDgAdVxW8QcfFdq+i3cwkakGGwGNfsp9DphNBekKq5sxul
X5fn2bfqKm7Ugx012GruuQUh8G8l4Ca5LbV9GqbEPm2kQLC/GCIN0F4J18NgCiEmU3v4pwvXMX6N
cryBQwvInOIWL/wEfEAAGZy/cRcZIyCRMO7YKJvNGHHcSykm2+oBSZC4xaRU7ntNXAOY/bDRFmr3
D0fi1AjvZ+jnNuwgYjYZBwXMavM2gJOKpELw+YXde3DdsNYWb57S1bVBsnq+PqUDRXZZiSrYWkMJ
s7z1tDuLVrgXgn5dOu2KQSVVO9mZ/iV8VCQApuk5Z0U+jRwaTOiqIQ8CFrfr4Q1LFTSDKUz3NKiU
5QozEaXbafSCZ3hEGqQgf4ubNRlIUUQtm5EkaEM1lCEBrKpWdVL4LeCjeSktbrwIA1jvPqYwzomt
juQ/CnhnxRVFSEr9kToW7RWy+BBCWifIqNTj0pIgbdL00dEGes0ElnEFd5F/gx3rIkUlne/EEQsO
cV+G9hGh08GQXiFe+NJrXMrDC6oFU0HRZRAtT902QF+jK2CQ0eQxe0w6C09DyzLX0DOdfXBFatd6
KXviBof0JHaR81lg57q63/+sPcjkV03NFfuQ9RJj9q5xdZQiQgE4rboxFVxoA1DmXQe7/c7vaU62
ZCKp50/t/cdxHXEWhLrl5UjaOETHwywPl/QPZD0cyPMZN2vai3kb3z3VWe1YDNr3CL7Z6WNXT2Z7
+BNUaKbQQJUnUrnzL9O8rQiKvAw++dCJozusGD/5njSLAMQBkL1vvbMfQMop5N47Ik/GvAfGfcNj
aezREyMJuvT7LYDLPb6LaBBXhZZKa/4dTlOXWtFFNIfkgp6+WL0x2cCmT8Zk2LqHkqFgcZfKNTWi
gsmUUbP1/arz5vOQPO0SIOIYVuFUB5DpocUldT5paiW5qB47sryPE6G7z8YjREO+IhmqmnSrEZNa
jlJDDtHjylGlIVqwXHq0quRrRIVKa2sl8TQ4pU/AjpryZx17fNC4O7PgZzqbKPst1CP2ImOKV/n8
DhkSG3dZzmzSEBXew+Idg5oEkYs00oX7V15n+9IJ5TVdkdm9QSqcluRdNUVgL8GS77hjcYB9J2Rg
kdRX3YJMfYUhcl+YlCwJ/iQxYiAxVM0YmtZMF6vmnLJ9EBbDcri/iHRgVw5U1Yb8MkxRI/uLBgBq
GQAJ67KWD40J4SCz4iqc86ZIZdGKM/ykKcry5xg1HvG+e/6uVEnPsliKY2CzxpfL9M9aQhS6U91V
PusUYQKDp151Yx2pojLr+8o1U22ZltrfdT4FXGRoVnl+SS+pvKPQRPxm6sYYxqLRv3d6l9G8oJx4
huky4+4pyLivNzEEA6DTQUlS2YCfdOZF0jXsWU/gEGDrUhdr6bdNzxXW2WbfIpqMzfhSGDbjcHmd
WzdbmfKm+bOIFMuva5Ti88uOPH5/wDOc+eamGmruP08Ycdkz3ArTzs1QTbZ7Fz+ymnXr2+AwrJmu
B3PPjBXHa2jnHGui22ZAu7vEW6/woMZfZyge+BMJJA7dFj6dSU+TrO08Covtk0LRJ/udm/E6kYho
zD9OF7+ghr923WiLJqi7wxIW9sBOIsDMwWNHBm2lJYEpdSLmyQaP11L+9F74Cj6Na+B5/kf2fUJs
MNMCZAgCMcGJFllyYZySQaM/NMA5TKL1sV89yijjEC1Ww4Z/CocCtgZKL0egc3cMk/vrMAyYUjLE
lk1XHm12ZiEegbGlv0NWXcrA/rYNBZwJ+HSxS+jPbSb/KAQSehfr3sK387ApR3x3vNRGqyCUh+Ev
E3HuYHl0+nvM2mR36zKB7jABmV3gs9SU5AvP+TivZ9yxdFGVbgQeeZxfPijXrUoqv8BBvBQJhzH7
6XNYvz/uP3c0aFhDQXvXGgF4Pk3Ly2pyiHKAvOhAIFoe4xOHjbLzrfptaRpk75zxQ1zhvsSKr74B
B9pTi7w/x7XkrAeXUdzJQuCQkMSuyLUQIK/jP6H1pCkxkwK0l5GxZs15dGo2gjh6wMiJp8OcQp3J
fnbOpK38Z9AxZ22bcZdTWm2qIkQiMp2uxWVMzPOKyAFRSH2BDG3lvbn3ZoJDw8OPAurn1VFQQlGg
ImR4UDtH4qMigtNQ1g4nmbkbEW3eRlCZj56PgxpIXPOLyqB9kn9+w9Jr486oFpNPXy11qx1EXEVM
H1ioFlwjV86ucAmO7HDlkEET7FR6QRndsTzfSEfoHH5bGWDiWUDPGtZUYZOMwK27aLn1MKD30j5R
G+V+i8SFvls5HJ+wliC0rk7KUXFaL0v3wKvfcKJW/W798AVzedDFofWUeXQeLNn5PNQuNB3ChD8S
4ABIpz3BbeHAiAynXDOmU99A84nOE9NK5N8Ln2WjqgvJao17bMo7DiDlZaKZncmPmG2xv4evgbjN
p8Ch6soxuuITjsTPu0gIG3aIah1kpsZZgCjpUhPzA0zT+ugKjeQU4ApFHiMakWqy3jAKYw358LAj
f8BcuJ07vo+bbBR+WplwEVJy9VMP2+UUejZ8aa9f1ZhZlFctE4nduwgNRWPgUDxWrb1ecSFBwRRC
96hmSPjGfgJ1a74xukaCehppUaB8YigfWND59Mg2E5FS6A/oeoBn8Vnda25AqXyStcIP+lmeLhPs
9uuYdebmbZocor5NbJrgKfPQU0VQs5pV0QWnKfsh5GhVJc+7o1yf0r/IoTpMkgXsNJ/VTs7FJWXf
xhys95Z3/+aTSeugxCEFqfgEcwgWDHXA/UPsicqxRs8d75UloOrO97oVOpZr+N3cKeh4xs7GKYiy
gm+1MGYRVWG9cCIl1W8p0VX/qNIJk/s8feuAhGI5btTS/suMJx01MgVGQazGYPu1fKVWyxorJdhu
jtTYX6r7QwWD9CUYuGabU44rG16XemwQtzYv5mO+EmJG15qlXrnYBIeLMDPzem5c0jm7QUGV2rcy
8ydA/iH6z5zhhABUXtJ12nBZ+X10r+fx4qcB3FVJMlyHXRsMX2gP8w8ZKhjYcjXbhF/yw3aSUSbD
43BBcGsNZk291W4zByrCvt3oV8jcocN0iyWrBm+zohVx083JnUgPc/dZEuB+BYOvutyhm6QEhYRM
lMsP1U/2ezbipSmbrcS4tivP71WIMZGgYRLw22XUH/yovZ7EcFlBjKGNoHcpEKXIJvGSeToV1v9I
R+fD91VcZOGAlJ5tuue0QQxtTUXL+lmaqaDfN2PKMZLJDdsBt/9Icfq3A3kf11mEXAyxOEPahJLk
jKOrh61/bwxFT5RRNYTNWcdEk8y1zRdCcRhYilAP5Mw6xMoMGMe9VVAQZ7e8dHEHJz0ASnLYaDFJ
jr4zcbEok3kV1xg68yLwdnZPKmOR536nem7SFNIeRpF1DfDNwvojFMg8uqZLUFUZXNpLry9DI/jH
REaF88nQtj/MHNyR9JT7d7WvoH5OO3l5eC8CsCNF/H2olk3QkaBJabNSPDD5PzhHCFOSXo3M5hOo
q3bJlcAC0sweaH1VVfOqXOUxY2QMcRgsdnxYorQgokleak+mbfOxti3dvR48UZdWKiswoTnjQw4t
KnMSO4/yyOoBrWLsg4qF4Gjm/ZtXw/evygVPYHPRv9+a0lhl242ovNW4+ij7UFidDiY2o7UnWYFP
I/gFwOhHwHz5gmo33LXLj7rhT7B2VQXbN5j+bJLusr+FfTSo/EF/wkhBq7PA3popgk/4NZkCAmvL
M3lFFEEb64FZWsBMKkTugsJWmXlJrFZUbEfA+Vgoftf3/5qCqLgM3S6OPp00dWJPH1KS9IOhNZ7B
Av+RJ2b9sjNdicx4deC3lv3kSDdj7ZAaqL1grOnFe3O2KUntkOlGf7KaGPsIieSSqSCGnzPT3mSs
/70UIkjfsdQbOX12cPzTSJwKkYkIVlMqxc08hPCKUz9cV53GwzQjon4bxJCg+mzXsf48GflVSXjG
Guyn9Xxl541rsudrqkVCz+EOSCDXWnnfS0YW5j38l0Egrx4C1yuh0X9LjAaort+APFYItpS1XNk3
iV66fI9nfu3EpPqfOF/1ZV8lhCfO3TAXzzGNjMjLcZCYsaGsC60Oqg+Pp+xpl2Cqo9nMX6MfEJbG
XV2hvGZUs2MHKWzsIKJUqdNZGWTRjwjghP7B5iFnzPb5/3VQ/P+xuAePf3PhP+JPprFj2+l+EbHv
OLCLslvqpUQptBkWf2F5Bpngg0ydF0JWOeSgKydnpCNpf20XcA8XfMpbJxeOy9J9hrD6/M8mmCYP
k0Vl5IV8qwH0IHxoqdH747nHR8zEeVfxGLFfEgGF9HN+Z/vbGCnk8xGmij3Zew8AtszZJTbErde5
XCLUPhEhEWEyBXhEZhVXyhZ07y8PuCqJmfm60LqgySvHLnoB0pXxkC46bMyfMWZOF7dan4RSkZY8
9+zB8GTmJ9+43cm3pEA2J+E1L4vOK5ARdPtTXuy8ElXooBSKh/vZluxogV5uS5UOK+dQlTenbti0
MToH/JbYvj6B3i3Fl7PprXl+WvSfbiFWYoCkyyrRTY/R4OB3leMkVjuHSBK6Ap8ms6mhfkUPcOCZ
785F0nmijDSSOeGjDaGp7CO71L9+cGmrEBZeRbcoIUHTKUG9uzA0oQ4H9fIx1NLssSIyFhidBHw8
089OIfs+8nO4SSKLMl8Gy7Dk8xDqbq1aD4xJ6civ1XKQYazfbNbEbKYsNFUG71j95bc8RUkMDydK
GOGU+2L1DfjfAP563izYTduYXgYW3muIfyo20T/4NIRtRQwPP8HExYiBUhj9OsdCyJD2k6lflRMs
NiyWe5/SXH/te2z8g9eNnfxjr+4u7hpFoW1WTVp3IsW9sEraM8yTOt4yXwsHbnUdlVaXB6TIXw3u
KHIulf7x+z48E3YR6oxdIQeD86/OfeURRR3OZXXbxxgw8uYt3OylmLmIxXgyHwqXMs8fwfBQb9aw
AMfEBMIyBzqeZWSy2wAeFhB+PMo8gkuo5jXk3liMFm62MYVb9Qd0JPmzKeWULrD+0d/3hyvgWpGR
1gMmH0OucBnsxnfPu72dwKTEQcsutHQW441PEr5l+oQ1fcGZIthT5ZYgVrhZgahAiufZa6fNX9aA
kp3e4FmAQtqOi3FrLHGxK9fSDDGbe+zkAMYNKTHPjlVU+ZJqkpkpyEuwWrXRYAKNGF58hmmKCX5W
JObN0R0qXYarQelVYS82TdCjYf2rE/B7K4orQ+t/WmKFpzJ+y65e75m2/QauGU7Xj9kUdvLZnDFJ
e10R5uVYTAYkOYWbIWWx05Gf8z82yflZPVSfFcjdsw6kiY/h8+katZ8U+hyB639u1TUt9naejSUs
gWTSrJYPQ5XMweR2j/ja0Pf1YcZyOBxlC71jFTs1N1P3j8yoG7ic/AqibtNChVGqt5/OfGxP/Sgn
vBWoIHbTvGtYJ4n7YXpcShvZCVdFHldsfy2eL7szP18+0hHNSZK18qL96ubs25qimr2nTmPG8mG9
xgdVsilgnyCsayQVzMrIgOd3PFwpgp9XwSxczI0s0OU+L5Seu554BgdTSNauMV6bcDa2nP0nsJ5T
q7zBKQfPqg5vqpZIeTxcF0nJHaFa4owZGoy9e0RQQApIk/O52Z9r3pjXQIGKwb8lFav0It6WO4Uo
LhyJykR5tPfvWTiQJFluABKOjMOveBzSx9ZNwfIGzHnZExfk5DOYhyvtqlX9zi6lHoCpFW7tfXpD
En6D4Nl0PgVTk87N/X5nuZsWLSFu9AbSnqXDkGjz3UHs+tTajzVuNrIuD71FrrnpvnKG4dlqDkUI
+omGGAkfr/GLGF+yocSjy+WnNbHw3GxrU4fMrAw+Xlbkib1UrmusQGtQh4F4G9vTEFHIlSkvlyz/
Q1Ds62R08SYYKbcO4byEy/vt5iruUpzQKkGsoaUl1ZDwT9eUUQFuBoVi+t+RCKl/qwlSsxCn2f4g
YQtLSiLNVKQohGhVGRb9nJ1n/DouYYRhWmsh5HV/kbTGFeDisq2tNh/lJZlBHaxJWu/fXUFRxeHn
Ues1YMgicZ8GRUWlmO4C95Lcregdl7tLKY6SCs0AjzsiDYJR4KCjKYeTvjY8dgC2XWNH1F83uka6
ExRHRiWK+r18sdI8yctxP2fP4VO37IFnpzP7pqCuyqG9FoiqiR4q1P0m5TCQ1oV7TL/V2vWCKU76
TfLVZG36Fv9zIOYlg601DWcB9tKyxeARrU/iYwkskERgUK9omB/NVazMfUMAz710ERiIv+yZizSv
ProXqhqr2Ym+fD1kZskzEiqEvMCbUjL72tOwHM4F/qR4e9XdoE4i3i7fKHBwh3odbq3pLbYVlwlz
EST0IGcfqmQWRGPXUI3P2rp1vesOyMkgUle6OeFnx8NDuj9TM8BtQcBZu56WXKu+CXSorJSsCFLE
+UNnfwpTmdCXdHZhQvoCeeopWIL9i3gUsXxahp7xmyxuII7Yv4jkS6KiJ8WaknoGz6Wr6HZnaj+w
RS7t4oiRPnWZ3I8QG9MKzdA5cserJG62E/pPeY8uf+qfSdUXgigMeNH/E2wq3aK+gTlgWoIxOeH2
38tR3fpZ3sslx7s/L1F8ifs8lcXZiecf69kgth353qLlHkO6ijZdMK9meJzUKtySlg6JFtM57mHH
CozplsWhLOOdhjkpRoB0YAlVK4lMA3gnBZuVEpLpyx1dyTuyid9KKrGjAQnduRWPV0n+qWDBwzFN
h2AxIyjFnPMbVC5eO5G+UAEYaQAlxK20Et3XlElp/qsWkSPut2v9Fe6Hguu6j1mlUrsBMSXsZeVC
rrSrJvbCwNVB4ALBGzmggFtyKKKzrapn3CUg/7ys4p+QSIwHRrqW6I6CtGN/SxiTkR8omhLigmM1
i9mGHAA0NmySeVtNsg6kj7zAxELT0uEQuZnyZnah/oICcWndnHPYNBE/yihdZXHRv/KwfOyf52hi
Csi22JdZH0XRB48/Z+Wskh6B/4XFDjTC2iGDZfwCvZBs/VKpUvqLDk1hnCSPyHmiO/iZT5mx4pM/
MQGw5kokutDce3xx6k7WtXeUP5jPwrJEz+SHkcanSPWvizjXoNsp+o2k0JYcY80PFEzazdn8u8sN
5OR0yjMnNa+3/V4itDE0FOgAskowHPjz8FKRtER9AVvs7h3354lGHwzrfSlVW/EjYP88glHaKKK2
MBt0nUFJJcnseahbzLC+b//zOuXRCK0+4mY3kZDonBDTVXlQVD5uqbUOweFiM7BbcVRimLVJ0dgb
AcLB8AVv0T/Xcf63uwl5gL0vaZ78LnozqAgwgD1vua6oy9DujxUWZL4SI9+t4ZkHkI7JRQhANQJu
O3zn716vV3jK/kOFo6QIoLPHMqu16YtInpLzout4MezTwiwue/h4sD2g+OQcYwlRkkWk8ZQ91uLL
0J2OT7/x7WGjYYFFbQZ1vZiWPmd267muhcKvoJraqowf3g5st+dj93voi3zJ4X6aPXgvvBcPKR+Y
j0DNbr+jw5uNxm+SZtfT7J1MicuMTpmoi/Q6I3kEZh5SgLWV3s8RlJiq4C+viFvZPZaG/hnx25am
vm7vy8mpzaesH3JJXP0KAOjEbP5ef8mnP9Qy1MfoySborq4zOlPy3PZl3kwE4eO9MCELOz0RjyFc
SywHAf+BEwXcmjCvwHgHWpneab0u2GQ4eI/ZqNPGghDwODEGzcfAqZSX1euumMOt/aOvu/TE4QrA
OMWMPUZKv51MtNGuLiVTUlsCylPxnnnjG6vf1jZFpcnIUU9etcJ/2+bJmG3h9su86nfz8KMCS66H
r6e9PDgua+0WOf8rWch8KbXykLr5uUZ6Uze2jR6nMnaOtVZkOpoyp1aJl+Yt67Oi1jnSj4gzTatp
fSWiRsRp7rhVNSI5DV4aGsMKCbWVsD0xE03nzBgSd3a24wRFr2KiddroPimNS2F4P3ybxDWG3JXm
1EWqCpBEXLYPjdBe47WE9v4vVYvhkw2Yn59TiXSNDOG+8SFDIiC4P4FikhHhoBz6/2KQe5LF6VWZ
V1kRL4Fo+dfDg8lSAbuTzv/dR8XhC8IfDN17Gh4W6AyILEkQlf0kBj+sbJUD/f+7jNAWAt4rSp2m
U0uD2NEl26WlVo2AQa3pwQCVjdXozlJbU3k4NXSshsuG2xFddVN5MSiQrsmYFSDyUVRGCOSZ5Y+6
/yUGwRk5C09PtWM+FrPMXgcxOeIbNSP6UAMb7wyhwXdrc2bpFrwmzuVDU3LDcRX/Ml3h0OGyWVjF
LiBuFcjoaH/XWKCNLGeVsfgWjWAloJ3Luggn5q3+9vyShzVr03h5eqo0S1R+c6MqwiNnccplAfnX
hMV22Cz6zKzuTYYbw5HOjUHBwVgXdKbfttV+PG6pkaLD7j+j6w6yrcmj+ZhztA9FwNELM37MVfSn
Qx7Q7I2tfWBMKPH9huDNApncz5q0EtdSzY/e6f2gifTvI+Hcw0CuE3WqJ176z7RKBABA4ekJUVvT
i4D8PaQ4nPGL/tTpY43zZOfHEhcfFXS7s/+6zV/PyiWzS4e6tDGITlzVUqivK95mkQyT/uWJ9HbW
286c/xCwkt5hODbF4IDJq0GeMQYVFz2NtESo+4Tc6zG3R//e9q+W2cguh0cwYxhvLs8dZQv1CXEZ
9VE4JxhM3dY70Ls/kh5K0Gzpi3fx6sGvuKyPRBxgAz5IF1UG05P5ONLV8w8xn8zZy05fOALd9Qvc
GHKXcQtm2mF7t+gHon3fYT9bZJlFNQhpgRFrn4LQfX6ElEml+pv2X+9A/uZ0HpbsnaTfy9WN+XBg
PKgS1oocsmOJKzIm5+Sp5KZMrVbgn6cx+qFBxiPr2Aa5L5CzwgKpygKAFN1TVBgieiMPhMTAFmvq
39o66TeqwoFNJ5SFDcVwkOC7MbPRqQT8j/+Kul4/rmwuLY5kP2ltwvJC8+TNm9XWNilwETtVAaBL
Rv+3X5tvmu+5FXmZs+RyTdbxaRmjKzl72nQgqQQIPxAByuegS/grmpwiY0AYiy31QEAA5KRdwgBt
afAHl1JYkqFMGoTSRgzfqimj5k3BDJWR3Xnr1aogeEeam7QDVIhcknrtCmuElBoU6UQXvgPr6ooh
zKUywzj4MzWNcfytSJyfmZZG114li6PtizCGdGr7/SmQC4Wye4m8L2xf8u+MMY7+4q20wKq59kIO
gtU30Q4ACoacOSQWK3BWVYj/lQxxed2L5kf7ne1bznH1CJbauU2PqKM6vvdJ1Delg2vlR+o4+9P3
KT5n36mHjmSTgOXTJk37lIZSDoc6W9TnO3V0k1oMHNE5wCOCCD79gAj3R7DpQPTLKpM6m07b3wIL
p12RmVHd26YNOZv9ef7JZ4qqRN2YeRhrjLx2qbTB+4Oad17vnGE3aG3OSC6a93q5isezeNVs3ZO+
QNsgpA7dKqPc5Ewdaro71tj6+o+aYnMmi4j6bhaQ73jU5Ef0DoTaBidxMYubOZnESYz39up2KQbJ
gFZ9o+xY/VQ0KjhkMo3sb8kw5YJ3LZRMUMVHs/TOhLGL0McCq7JM3v0aw8Eh2Ug4wwYmekZn6Z7R
7rBTQ0breobqujAVmsp4xWrrmcHbF7hbKPWx6RV8I2iyCXAJsuzSKGM7D/ONWioLagFlnsNV5uFp
UpE9/4pF06OKigOgNelqLUy4oLWt8AH4ayYPcPNRzJFiVDdweTlTOW5jcoq1XmReUXCZARzJ822x
XwdbYovYZw+DvzjK1xcz6QbyJ9RiheKFU7NmhFux62eC2vUKA70tvREAh1IpW52mUTooqH8xHi7V
lrjqHe+OZ1iH9qKw63znw33ztrKSUqHsKAEQE4yGoS9s4SRiNejK0S2sgpdC6UuRaTM2q0XLLASa
eYe79wpH3u6XbQQE00AsIY/Z9C5NsDpg0gxYw95413ewMny2vdg86gKhVIYvdhHkCucJAqGoOgbr
6h8I4p0YAF7MdDTqcLer0ZFIRRvT27Ht3WeE777nRbXZJUCMf2IBH52co6OB3hnz360WfsFCgG7f
7D3n4UnlWEwAi4aLLKma6ZYWUmn8TE0Rzw+edFRWQvKhsAMQFKBEuWlWXr2lR/C3rKwY8n1rs0IC
UbhStGK5AQzUZtcKbkfX68tN/6JE2fn2Qqf6xFjioduui+gjLNhZteSYFFeX+SqgBw5qYlXA8Y4f
4WSZtyW1Der8lM8CkK6bmFBQsmIWzcpu/NHoXfyi23LLedHXxDaDSm7G6q0Lg7/KLxX3VFDv/eg9
RaCb7+vCWuR7sSHgIOmmJ5Sy69+Y+7EYROP6qa+Yg4eZ3cFK0ncYxw6+eDfGoYBcgxYXDS+mVXcH
AZQsanddaBrunso5U6qsIM9UwZV4KeGaXgPHBI6gYYqM7zcCiAhZQnfksgja7EVRgxH3bvsvfCze
VnyeGDH2UB930iFCEnqjTBVS81vvfUjAAURM+SekNCQUejVfXvIKU/XGb+AbQh9BV8Y8jNhh4LQj
YE9qjtbl+7+UYSM3GAJWhvEk56fZAiNEuj0SD8zkH0jNG/P/kXfLrUsmqAXsqEJEi1Ee8oNDpuED
G7cEXcG5bKTAfsNlxI6lO77f+Pi9fueyhVHDJsx9NCIzyzuNRkGVyeU4a4YF5lYyCPd6PAGoxSey
hXL36tzwG92VN5NAu3dpnlZgMlVrnCcRWUtpbzcCwNGuftw2BQVqXBp6ZwTRMFjhQw0WsLm6S2O8
Rszsf0vhevOHYtQYvK5pmcgN6WNboKA0NcCDtEZ5xpyrwUN1ZUOMk+QIckh22nI0BbUa1/cylDnr
BTBv5BoCY9gKUhqe8W4wHxCK7TKbkqbicE8m5N9jjrfggQaT6+B126hDWqg7YhDfu0W/JTvXvqqL
R0Gq4ZAuqw7ctT+4VpXjY++/SfCgWYL9Xsx4bwgxLG5TijFcvZcO/bWfA7lxUYLcp5ouM9Gbs07V
6b+o39vl85XVLRTUx6OH8huJ8zjMQGgzN5eDLDUGE+Y19NvNau4f6+Jg/JcaRPjbaz2MP5/Cebis
WAklNjoKQiklQiXE0v4YlGu2rmWlAeDe7Zm7bD+6dC3fGLJy/DsPBNi0/n9cKlBxSN+O+OVwK1Ub
TrA3AvanBnsCZKnOvsfWEjo31TA1uIOFQK+dZxzK9EVLWVqCUacTAIXOWYY4Iu57RLLx3Eox9msj
W4NMyY3P9RHG3DoDA1ovOsAXxxvrjGTS6DOskSIDYoVqEcCb6n47ALMjFY0oNjFYgjPZSzBXGedP
cyISQUwNko+ubdlB/XPQt3xjBjtCOnRxHiIxgVr0BiTd7G3S8SrvlDF0Tc54T8ww9I1VFiZPEMpF
7AhnxafW1rWA2y9i2DJEqLYq4v3xLq/f8CLdd3ll7E7yM4Mc/OfLdZJxP2lYyGHl38YkBpvWyclj
VNBsRB3Uzn/rbVg=
`protect end_protected

