

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H5lQJsJvaeLLGFRhK1oe708p9zTtXNXItx2KAtknEaAF2yq8IXwKFiVPbPTO8aJ4G1wQZMrKgMvb
6zlyKbmneg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RUvUfs9jruf9OSb6utxk79ymugfgdQ2mgDnw22tbcF4+w9YY12PtlphQ3EwSjE1BR+YNcfcg2ppx
nVp8oQrlHaYHLiZdJQiFcET810isTDBwI9+sjn4Ry8+ftUrGRDkzGQghSG1UFCnSyA55dNVCduAa
//ZGtYPCXRggO0BwEzM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GRoj0md2TTeeyD4XkfgAjr1JI8z1r2plHgATS4H88EONpa3oaJwG10L5TE6c5MDXVxHb/m1WeMVh
VBt3w5S8h9pf8c485G3a+NVnNsA2vHPB4cEC1yhvDIpNkeqj7HvAUARW4zUkp2MDiimsNN00ZMVQ
inLzBlDW8A6T3Y2b3GmoYzUXaMQElMyS/PaVNF6Se8+PIRjTB8Dv5G+A8K7PF3j0h0gW5LdMZrCx
isigyN5NiqJ/3ZZGLkd5XiuLlr0DetrgHdwfifFeF2dmLtMjIx4kUkMG45tToYmkQS3jwm191cux
eXIUgmzmvPZHik85i0iZegdiOZ1LzY1yO5OyEQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UnEKB1f1t5V+eYV1nijBv/smbMsJH58WebxNSKYwmtj2m6R5AlGEZE0haiR3VYCxPRjmiopDDdr6
uBQOF41DIKvZSm6YCypTeVt9WvkLpXTJIiHnLWz3IV+uvKXohhIry2Pg30NMC2EWPfi43aTNvtNH
ROJrUVVcDZeGvVPmgRI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U8EV7GGC48XxGZ3G4wShg05dze1bZdqSUw7dITFWVJl+2U1VEqYTGCRl5zpa3cGdqM2+nFugC+BK
YIux1TwcaF2Ng1I+Bp1k4H3BhUPfmkZlNiGri0KnFOiDYzBROYyyiUUX4IECNCLZnG/OtNfakQoI
AjU6WqtEEQ5JSpZpL5mpGWt7jGfdl9gqPeY88IdcWnasDywKSPqo47azQ0KIzwP9UejnEHChmHgr
3Gpvmrmywo7/+/EQRujU1oGF+ysfAmqchOGtHLtDFJ1h2OjLVkv+puXArlpXpB9wZah1XCGw2FON
8d2jAO5M9wEJ2bQpFyxmedBeZ1Qj0cJQKZW3Gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51344)
`protect data_block
eAigmRBLPk3QddJOwFHV1Hy1OrU1ghjQ1uM2jdnbfZ68HOnRK/oESHr8ma2IGTSEyuU/qsa0YdbY
oNSTC1+byGcZvc2m7Tn9afK5RZqinuvQwMUez+vdltQ/j3NRL1LYgsiWCr3GLdGmo2tSJqTLxM16
LW8z/N0AbaidzhfPOSWBTu+b5qpFWrYc+A7LQDfBwOgGxGyJnq/iI0ohtt9Eh3Hzw63Z/8bd6DAn
YXPPr+ko0FF0ZqHageGQm+hJyDZMKBHL95ElcBzmjX9GvuQE9dIXNpO2lqS8Zn+vEgNoEznAmblY
61ljATp7LWeYtgaEZ8WRmyKvZnDT/05oX0umFCEUU5Mx2o188JdLRqf/loB+2OBi1F5YcvH+tLKy
nVYWWY4wqWsmAhqU2D/VFzAEuO8kgitY/EhJgf5iyymDMaHPVQXAxM7vbclX5FMUc+3dCk7Q/z9J
SuYBZSKHpoFi7tvuZmmSbS0Tj/wpkosffOskNFr3Smr4XrjijisNW/ek7YjsgwmtSlLAW2H01TNh
Z2j1wcpm4SHctnl7oYysCHdTvWzS/dMshADgjyxrIYuGywgbIkL3ixPGRAdpK65rBoWduV5plDG6
ZHsZB+Ii+ts/lAA/6RXNkjZXK790uZShtFAonm0UaWi50ViobWZ+7UgtVLO2vbXO2X1lN9FhvoDc
sy8Mv5NHI77f56cO+HMvlCo0JaCL17DJfUipaPyHW7grP2TxSg6pwMMExgvyUVzbgfCKN9SGig/u
HG1xBewE/czOJGdNQU23+C43IwBQUNKYY5CIONfThwp4CfA+AE+gaG1oSfI9uKopmKcXrQbHobuo
g/gLc8M235Sh/YvgkLoi6OmVavj6qDTOmES/T8OFG0KnoK72MGIqTVV6CZVrFSzBh4LIvw4zGoe5
unUinnRx41zA9iw6Mkf6WZM4Ivj4JA576T6fKZAcJJuAiwmUEh4hUQqZES9ec0tl1YfzYAz8SkO/
dy2jInRjuDSkEKLIvSSrujFgrnAmYXBi9AqrhrnuoOs/pnOs5vJElQ/3YwzNv9UXV1/zGKqzYL+h
3BpOD9oiPT+WXsloZqudMNlmr7r/PukgtPClyNef7Bw65I3lw9BkPI1cAenazPPwj1FyY0b8iDA6
LKzUDJTE+cZ0uuPLGoaWsiBIkGRFr9/4TEVT3yvvXNxptdx5x/ARW20FvW4OZuukaPyGOQaSKYcq
+CEuwNueCxTf0zmBIlMPMvEsAR2AeWy/Iz7Fj0FnFSI5+X12pnBvftKT82dS/YOrLJd8SH55leu3
7MmYl7Nl5eYpQNBUum/CGCFUmhL70QpihWkxT9C85OYODIawn/wu0nFF8dZPENW/EKkyCkWDnH+U
QUtxelZb+KYMKfbIZsbq39a0d9TklJv/O3SdMHlR1R1yc10rFCgcS7svciAaAl0YZgB7bunBTbO0
OBwRPAH5Mif3Qroz7ULyZoTDcvl5agzS/G1brfwMa3TRDXAPUy6nOHQq4hvO45DZa83smgDoj8NE
+5Z0/9V/YbaFIL1dtWMg0iORfpYtQ25jVup09ASw6SJ5Y+PQ4hR2T/jCetXRLgNSAmrfC2zMF+Jd
IVJhCQJRwoh1YkW59dDqd9byv09dkQxJYCO5BEAgP6zQAr2U2XskWn9utPzn1I7yZf+EmNzQYs0C
2GakIfozx71PBYdhvmuEMuwpe2IuWAbdiweWY9Q8lbKruceALqEDk7DsWL4Jf6yNOkWAEf/thKP7
zLFNRPp0YyNoSvuy522bTJNoV99QYwhcpTmAGDfB7LcWpD25jQExC66b6UvXdjGgTfZPv3+ZgPX1
nULGQyKhfAFZjbLDkaBs6HBBhQMY7Aw0STaym0a58AiJx78IXq+yhnz/v54F7+bDxQUr4H2/uKII
zuN2RJtvCB34wxGqZMwZMIs++V7k4sZRyhYpO+MQUITzbZ9TDLKUCsTm3Demcg3bm9+CPvKNrWom
KxDOyCUNeacJuD62nB/J7rmK1FHjq4R1I4lzz/LOr52/BdTYeYBmYlQRTglcCORrkS01m8G2iQgT
PU33homq83o3ezANrTj8RcLFiu6M9LQi6/HMSrhw3CyWM4adcJqejPQDbLhq/hJWay3GGNtGsG6M
uzN9T3PXaPOaj0wqk36bqJZ1Ovfbmmv93lhoCoNLhYYRJUFlZ9+Wes14jrs0fiMr12bu5nsB1EJ1
qLmsoMRMqGP6ub9ZdEVcJWhXvXfTLDKKpk47MzWON+8ieywIH/ZsU4WXTL0/2T/oRoXQ6X7Bmikz
QaiBaVK8PRSZPCo5fbM4rv5ODBzy0bA8mu5VAWlqGl2DxZZYFAFW+FXWa5gunX25k4k2rFIAu3n7
TjZ4rsbIgL1eCuAoVgKw7v2Irb8D+g8Xyr9L8FezOQ8/IJDcJpQeWKyiFYlG1IJL450XNC8luUdf
+mtvpoxzWEqAbwxXR+mXlgW33hot9XoBffn9as610lNs3AS5cNhJPNEIR2oRxeEwhxRtBlqcDh7R
0ZFBh7U51c6ekgljvirLLI89qSqTH5AZmzsJ4c2Y70zxD5ImoxjzCFo+draI2iIyVjD/stPA1Zok
a5IeP+bgQ8EypZui8OvFySG4AswNbtZ8mUCuXjE+aIE4+GVKELyv3IdT6+vqPewXChAu+Z8oFZqc
V+2v8gTWBJDtw+s8FGcvEVwgYx/BJEPaUYG40kT4L/87RgPuO3DYl0ruo/Qjdte2FtFI74ERcfXw
sM854Qr4WjAHFyCgZNpBwuchL+ABZ7m9ogYSLH+L+LD+kN6Lbptk/LyIXST+GYxBg6vD0msDz3sA
PngwH53azC6k/PBEGhW6WWQQJ/JLMjYnG508YtY8DJ0B82kAPKUK3omukdSYFtUmajjabp0jTLZB
4OvheErGn1B8t042WDgxnU7Aq+QYrQaSly2nIZOyAXdRfNLFSXvp3+FMiRmCPtWP6A7Wg8CMIqrV
d4IJ00LTIz4cV2ie6XR7ltP3BOei97myiKeGx66ewbaYYM7moG9t0kp6h6mL3xllkpKLDOAUDNmr
xwBzl7e02XpL0WZX1yTIwrAaCoTMT3rAtqM4IQ3jVvAMadt97nQkyuQA+cOD82gmoIT/a8NLCTgR
5jUAjfwafXGRGiRe6xkD2fHzWocxgt6s2MCnI+MkeDrl2DNgYmq5stf/h4uPfNASgLhgPLcdheoS
xtmibts6pdLeUdoTzs17daL/5xIUTRDcewIvSgKE8Rifz4zDtbeWsKLB7CxhjPV4jGwFneIOx2Ij
DdJKzw5MW1gsi1DNujIVJV49HNtnyuGUviHkfRx36OWel1X2+k5heBdtftog/9EDNl3XG1UUhFND
Gz4Jubo/kp3kanx2zkGsS1RX+zPoB+Y4a/kWklXfwvLd1EApscn/RbL/93YRieoBAsu1dyvcqIcX
PQhWF8Nhl/p+LA30IvMWI/PvwvJg0Xk9uVrHvpBMkCNmMPi1We23wD27VmCkh22SVhQD/hkVxvuD
zVk2/dlTPHP/YYLwcOSYDBxfcL78/CLxtGbdzj6sJBuY3aCwzSAFxEYqzSrIARPxsqbnbsHS5i+E
lczEwHAum0stCJk20yDv3fdsqF3IPp83Q5f5i4JNX/eIjtKGEN/COyCigtC8CswpvUYqPrYz1DBR
5I5Drc9NGDktCFTrCW8LpSee+Wjf/EkoibpIKBDWhf6SNFtPqmaR9pZSJI8c1jNI4fIVe17j6bDT
M5mh/F7mSqek7F7+IO3HkklW6sX8M2Jzb4pFm0MgPzq3exV2SFKI+V8VrEBqqpou5du/EcyOsZgM
d9fKzrAhYDLJWGcwP3barbKqy4LHmvJLHvjLxd3OOELjwn1dTJ3AEFfwtS5efgfcEBishbDVt7ZT
6DVGaiN3iYcnk5nAd3Zu/6xm9/AiSuyrzuCwgQgRlkN4EMKVRqOEINRxEd/glGC1cYr3+GGH00lC
JNXD9A9S8Br8QcRr0DcBZTPjGtpMMHaCXxHBHjbZP6hYH9k4umV2s75qAjON+PReHYt3eGnVgXfd
w5ksMxKMiRyVL5fnl/un8xmXdtGkZ+V9NWXIHYzzH5hJLO3MfbEafTmC9xmExJqqZvkecfuf1c3t
4hxNyC3RDaQVwrvWRKeElfD0xS4k/kRsx05Zx84Zp4GAd42YwB75vtAq9jCsLthpqac+tx4ywLkT
wUQIvEy3D7BkMZmxOuxn7pgs+FkdZtsxx3wDdZVzYTeonUVF4UUIu6dwvw0QN94WBE87YHv0uSv9
LXccYwbu8URS4lIPd/KRSPNSyKGiZWzTAvuT944wV7eBmY0FZ687xeloclJgPYNAQD+RuMz7Zw2E
uLeuuAKStvo6WTVFZeMGny3CFvonsFhNOvv7qq1xQ/efVV4FTivl2ygoF5XTayTIPIJBL7QmLOy5
QRP0QjKN+6cU3/sTTxMDoJQo4kUYgyCjn126ENctUzfIyhRmqtmdcdJdIQhImbcX9bajofzd5dY7
+ILXJ/CLOhFd4hiwMkSeLfjYSYryku1fxhYhenkgQOe1bHKJhVKjsQJd0Y1tTo2s9l4+WQmMuIIt
K2Xd+HI/TF7g22zht6NuvDiXvVDjCBGhjEriSFDgTWUpBi25E18O+j/IfeAmTvMyL8x4HXG5bQVR
LLK37zSjBNSmyvol7x1p6uyEr3EQaLK7M8JSCdaIfsFJV3SmR8VVfiqCaHY73pJptrVjcjIktLwA
XdKLDhcHfnulz59j8fUcSwRSOMYdt8e9LHhj9TpCw/nGuUhmrX3aFpqdZIUYcECVBejZgG16U/qI
Uzyk8SmCVI6axaaC0s6Oeb0lAI9UwPnlXfOZN9BWlz02U3eM41T+5yMZvGLS9xkG3f6WTj4VeMtq
bunJqhCAVxvcCsQHHFS/4ps+I5lzKPbPwjHcCwESBAq0XvXi2RjaNj7dqCMh+SCvLdloSj5GUSf4
1bht+/B0K7oeFUZsWNcb5cSFKw3l1gHhFGUIQnmGvWgWXqGe7ZXOb13o9WBqmLk5KfD+MxyDtgvE
aQA0I82oWStA7INzhR2daSufeCvniGWPhgm7UazvonHvewYE6kWPam9j+sazxho+PqMZ440I/bY9
DVHyI+/OkThZuXoV8mVeRg2ay6r9WPoseafynR18P96EygRz3g5OdjogU/GSNqQ0ob4Fnj6xrRMk
FxroaWFCIFBPW4NCHpodTz2vElIwJjaKqYYGDJMxa+eabp4wKavU0EwK0IXJFVV7i48ibKRVlLk+
v4fGHGFoOFSdjvnv+StCPClLEUurzhZMW+PiORfR/DTC0LrwMpJVWb1m5oZ9jHMkVkryqDeoQaKb
YTzEcP2zw8cTHMrzvy8ATYqS5ax98iyI+g5a3kI9AXjaSmp1i2MbRhJsKChS1lv4txWaOV1I+Zj+
oYWf/fRSf/NOCvZzCY+YP/7Q3TxRmiHoSfy88CNT6C6dijmkhKajgRVij+0VfeHygF8Ax2rNTY4f
PrOJGRGqR5mRp6qrrzMzhyPkMOqcJU/WLkwr9c3ARB6pjg8qk+ojV71xXSvYf+bPly5zNRbCvfma
lTXy/PuILQqd5JRJ63w8k3/Ndbfo+ZYB0JJiX8X2Z4N36MUfhsiMc8CcGsKwRFLYapBFRyJppcR4
fslo4LmGmD1Z7hY3kzg3KYJlbESGas4KBC0shjqsOA3r7fffSvOlXnRP9FmeBoZQGeyjGy7suHw9
IpI8PCqddjT96x0HBgO8J+jeLFmUK1Zfxp0TKUBag5GkChQy+Q3gccCOSf4ygLcqm8yTXk91gOQX
Ch/6aaLVGXr+TH6qNsvdcTzbDBU2GB92gqyAfDbE/Z3F1xt708LZ014Qp7sNPqQBsmFi6nFDCwcf
Zgdlv427syJP0QFfyZSDtc140z5Tm6jrjKgbxKl3Q4QqYJF7npiGM4WyTXLrrVC1yBhU5lzq1eKL
Io70s21vPAhA78OEYVqnNSWv4joxC551I4uplmkgfYkb28RFlCYl/mKxLZEdZ/4Phi/MFa6djtPN
kkz2BqBgjv0n87j/kykVGd8wvbHJM0xTeu1PgAmT//Fjnvoh0/81XHvRzmPol9q0zHyIoaNyv6tJ
mCdAShlxdNJ0aIz1pBSOhTElPuP2JYjrsZrC5wz35TgZh8jVAe/42lUoaDQA+X1EQnCIVfdlhYkg
iSXTgFh3Iy0FZi66RS/MM82d5VH3hrpaWSLO1W81QoK7SLplV4RgI1U2UwwpcVN56X7PSoC1MhQS
0ngmydGqIYzkMgUJL8zsEm8ru9eqqQjxfs4XjOUP5FaCYFOshkMJMVVng6wxm68d+UQtn45ofVPi
prMb6YkHPNRPNRWqNcYm18YarX818jOF2cJzMucXnZPdQGibiUHswFfdD7heaFabY7iTZZNTvmax
qnsvgS4m0NGvQgFw7Y8Yh1T6Hc1WScNlNhMp/m/E6g5Joy3IMeRAz6eztEc5M+tNK7yGdGo2aCPt
OEsgXHDfy7zVSvnRk5cMe/eurCsJA67f1nWZMTWSE0rClDZr+/zQ6nIbYgmQ7pfAuO4psWhcHEcH
HLcFitfV41NruG/DmikNBVP09KsfLSAF9AUWBd45Biurig3x2xkvqwP2x3OLN6efQqHgF9IudQoS
BPQs3M/M8nXMVI8eE83QsJFbMcmOctuD6qZKo6w5zH5zJW2NFb3s/mtDcgqGb29uCxvHZ7nidfA/
b7RBZ5i9ZWtB+KcQrgzbfAUAR3VI2Nm2nBoq2m4Klgfv6kCt8u+qTc1tt0O/Nr6DqKJTfq1f4Bg1
W68x1EfGNq/ucqWn7wY7AfT60cdOOA7jgvv+2849LfQ5tqjUyEoZj8RH/CFTM/FF+A6poFFMuaje
wxTuyfF9dJjq0cde1+ZUoRiI0VMDJw1x8/C27ExWskhgfRcnQFXU6PxS7mZqoh3dALnnXp4t4LnK
n8Yz/sUEmRLdvuUwhdWTt14ldz7w2vrs9E95M7VE9ka6Z6Fvw4IH+UxTodMVaNgOc8Dmpju44T1R
s1Tih7NByVoM+FND9vXWpJsHmbFdKaX0SmkI2QSff7bF8+LRH3E90UQkiHEVz0XYpM9tlrz6Tvyv
gLqk+Db44/RaJ8c5s1ZnA7xoSpQFuCRGGVsJZxRFnJRm5oJiUmJNOVFa0Ne0WuyprUtTAsWiG5ie
XWm1xFzPdSi/EhyGaf+cYP7hRP1eJJh/VPl6uqsr87IHCqm9fD5hlg3x3efkjlH9X0zGhhFLJ/IL
xxUDOYp5IZUmxnDy85GQXRBhWLvR/lkdcTX11TEPuSgtshJg+JdS/sTJoFWgGBC8uPbCNFlhxBm/
i/tDojv46rjUyM78wL5cr8wZggZsOAsecJnKc2MojXAArglSR9BkcolnNnTPEJ21EYYI+ofeflzX
RvUbxHs5Vex62senuiHNk3Q2lDbiEWenXw9GmR1z1HIivBeqxmkROS0ZeCaeormm8UblYoolNwmC
M3+5j2tekE9sHwnOxJ8BFooFNmoJOKw2XTU6TavR7TBPhOoxCMsG8NvnY/xtlattvGYx+M3yLyrg
A+rYDq5jQGvJwUh8EdxwN9Z2NZt9Cp0VmBHmTJD8w2z/QgLqi64ELmR9xUcAXdk1iqfWRati7Iz1
eBQty37AoXiL26Zk2K3dLahuKhUuF4MXBXmhUnuOkYZG/cSq0Q4AGlMJqZardg3LsYChAF/imD/w
OFg7/NAy9w0GCucUmea89aROLTFXZt7Lcznr9W5RvxOKla1sbh5AiaQqWWsOBBrjenQVFmkURqO2
gRInR8q4BZJhOxLQzYS8eFGVXoHoDVAr12/wqPZD32/IHs70fzJKa1wNqh/N5D9fZPNDDfwz4Gbm
kyUzRePamMQ/zKyrzN38EnnHd/fV8t54cgrEwHvvGcmhrl9NcqD8YHzzlbk0PvhDoyMKHC5zNyqI
WcmVDWNHAqdn052cUjZytzcK9pGWg+jThvyCkJQ7PEY0KrJkBys/rmfPhS/i9EkPg2IMdkDO9psE
Opn8iH31PA26iMha1uM0goOtGUW+mmoqGEW2COk6PvK5B4Dqo+J2fvWQFVh6inb9qkbyJvk4GbF8
x6/m2DwnKXYcbLHbsJmGCVmNcctjUfKgskFXzFrRkV/Xriv2tCO8BUtgixak5SzPFqyzm+VMSknN
F4IXGPyZdVwI4sNs+gGlSIOyY2j0DgtX9mfTk8XBp4m6cFXU8qxllbaONjZnwzBt7PJxpG0lwUmR
SYeNeJxUBS5XR3OhoBB2NajL7xad099SA7BhvBCANgr5k4/6NxBgZWM3h/RgHFvpXCa+1woP47pe
RCELT57YA3Ig7Yq+FxQTW5h+R9PodRZ9GXqyWUcXMuIapIYeWmEwtmb2bntA+INg+6hCPdBLue4F
vkWqLDWgFfOYBp4HkTqp8qIwVvtTQmrta4hfqs1cvASxWmnoY8lLMCIUXjeToHzyG7naPlo7elih
U/2tPfjQV+NUuR3aA9SxLWAsriVfdIJeAMreup1m5JBM9aQSj+vWhfpAeZj0duIvxsMvAqiJziUH
rDyE/5IzQLp8RR135/sUJn/SsyoHLuY/0trZqLtTtbOEFPyEw1T67z5qQed6tMvn92DHHx9FCcUB
illtYcU/bDCa4u+mHD79okXf7ww8L82pj4vFs1Yc1zGsSdN+BEH88Z3WDbd3ZbXybRnEoakbW/Pb
t5ScE8NVQzUulQn8c+iR/FGwRbfe1ILLVyZas/PNaNIVh+pCqTqL2insaqwfg2+zo3spa+SaTTtr
pXGEBYEdtcoY5SEbkL1ZWk4HR9Qdwm8gDxFyJbS0cca23anyivTBv8Qem9w+EuUttV/ZgPBVQtZ+
oYIhUiRsNjFd4HORGG++iInHeLFkRzTljL9aQC362ad5UWGDenSg8cpwP/kGves6XRtBuo218I2j
gTMUdhOGAGmKAbVWAhD+9xmci2XEYE0ey+AjO7pueycyrjyljJEPol8awWvKxcbbDPiJVJrHx10e
m9jnVhKmbeIK4bNfT64S92heIae4DhUkuKUeJAYJlDjAFRN0Mb0Nqy2z3s+VEVH+m4BJo+HU8ASx
5rrNqCOVghFnnfJAnVod8X5C0SnI89x0XjrJdb/sA/yir9dhho8CmMCMcbPd8Z51eVnU26BHkZcU
GJ1tLjPnS1IoQ1LCI0VOCbS3hpvp91M0xV5LSdD0zli1QJaRWCHmKS3BMEVldI+LeA2L4zB1l1NQ
8KI4ZvbgYtd2Kue7A3hZOm7O/cxBbAa4M/vXlEp3xX8EhAPOSfvjKZ/n8QKr5eOgqqC7gifhMDtK
ulgQ88riQKGxahXkKx96wGgEzA4yLdb2X0ugdlOPnmMCkVJoSu81TUf3eJblkuv/bqQUA8QSfzc2
D4IaQhgFSIcV6AD3pROtYNCC4ltuJy/VQ1FbN2qs3jbUYGAoyUpGUNTd2816J0ocUOKoOLNmaR/G
C6v45d7aG7XdQyc+pnt0LjbACjEdIxliiLdBJCA7xfZ/7X7S+kwH81lA7Ud3JLYZ/EvURLsUzvW7
xnrIX1/AmkH88cm/cZloKucoYzjW6x/WvXDRbhoofd8kYgX9wOlAezmqbEwF1c25rxvWH2WBuYBB
ndWVyNK3N4hvpeQ+/Mgd1XYS1wVYGpJqAh3UNRu9PZHOAanE0J4VB8qz58D6mwd2PNFWrzu8qaZp
jbevNplMDD8L89qXjPFurBDoByY/4CUkZVnAJIuXRDOz7u2EoXsHfOh8XtTU/3Ldw6vfniz2KpN/
Qiy6CfQ6E3iairWFzgS4qF9Vmw87cIx9ZS6QhFL4R+8Aqvf7XcoWd3NiAD34yUQm2Bri91f8SHtg
ekMy1b7AgmC+tmwTWzpJAg9Le5CDmYIW4Ra5SQ1SnwbdENc8aV6/4tJUpslkjSur8D25xZ9lLy2X
N6Dbp4l8a4RpNFf5r2rF7oVV1hX6ozV0pbkmCUWep8PNhKAS2pii1cOu3jOnkLpPkL2f4/wePexg
WRS0LGi73Z/mW9xro2MaXptNbp5wYxnS8OS+7IDSs0SmS3gTHZsrFBArZz3moAKNtaHyKWPr6srk
DcM2H6eY3pLyWBCqHKrhYj/voYJZplyFBPseRdcLN6a4xyoon6bvIVd2m5EMK3QGGT9d4DP04rCe
ORoFpHDigaJIxMH4wY/T6Xg+fc6YyyDPEm/Js1tXi4IIi0PuHFgLi20+11HwIPbAAoomEZcR9iSc
m7O8lj7+Peg+LV9y3K/j2Vzlc5Xt/nJIh5KusdKfBd/COBcYQKcSXiIzp8QM/GTawu81qxN31e+s
oHyPeByuwiwE5hAUgNt5fS6KzGYiX/DglZgZFObnFHOBFKvT2MdkJNzyOEiYbi/S0EVluMVArN8r
43XaMTUK5az52kMXAekpl/gInKigM4y+GEamIalBHlRbOoB1yvYxSHZuiL4anBgvckHwGPUW03sF
mSZBw22Z8jVjbS13qZz0UQNgDRf9nQ59CE0rbFF3kOQUuPiJ3JFyoLaHU1uyGz9Kad6dKuImxLMb
qI7SDjJ7pz3hRb5bBOVZ47z3/oaCzxtnP6JBkzAg0vPnVVM2tjbh+5H9n+lnHXQnb+FIQ1j2Xz1T
8VZHFymg0t0txVlM9yZxJKVqDbxUhZX0uciqWXUj/CZFiNCATEpEqK7BC6lEXh/BPJwlu5HNc6gr
eTIGmtJ5XLa8Bp/qrmfobB7W82sRMlWHlkSUiRfQahGdMNFpy0ownYnFiEEjFxel7I6ORyDjlyjl
+RoY8LVFmVp45vN1n5zdD4kq5yd6k2+GirbnZfYb7BShSl6cbi2Lc2xUfzZsmCpmF8gTGlBg3rUG
L4/Gv+fPwQQkmpFYJR+Tx3IvOUkqWNVDtPf+jAw6rZKVpfwI+s8gDyx8C3LIJKOsEgGaqvE4P8vi
o90KgsJXw0s4oSX/76VY+7Xs89jnCLQ+moRMIwGCrqU0iKV25JCZHm/Zj7PPACMI/G+tGMPXfslo
9xperiaV3uPH1GHgaaIrvRMVvecMmz9W39BaIOjidBVd2WrElf1egwKUXQalNlVPsq5L0eCWFG9o
j/3g5JaRNXnpzKY1XLYDX8MP3KG2ZrzvcbEvK/xvSazYfyNpxe/hnMRCSjDIk/adh0jIO7PpGZTw
eoK45DJ8PL6GLyIisU99k8Mzz23tq/hKFtvYTou2YuMIXXosrLe111Isy+QIYr57OyZ0FdGStYnB
6yKG8UH3BommV7qbnnoyqMhRr6DktsVHsiC072BQ2TDbCF+2/kclWLGJNGcJK6t2AlfbJHUFFT3r
Fy0uRmBtDMed4g8p4VjeClkvnbU+HaoGzt63lPiwRiAhCyfyUZDDsKwO/1bi1hTZxbTUQESTAJWD
NnzXbTulW6xVi81vgtO76DHldqEgvxCAXYsgdo/lGstkbQQKz0o2Z0c8AEZu/W5hV8IKGH2XEaW1
kpashnTZYO2RtUMBbDSIpUj2gsjCcaCwmLhOutLIkoQUwgGoI3Lz0I+P9D9Xa6G3qr2d55DpfiuP
ZtnzecsW+b2ja44ZmYelg9PAd0+jHBLVhPlDqo+7JTBeYoMBuxzvQr9mSsd5qAlAy0ykpb7CucD8
ksiptApCLKlRA+Y/DiaM+tt0A0tIC2Hb831BiAdkPjFF/FphYDlqLJcYvIS/O1DDgjXjqWdlZ/Gl
izMscEd2cgCdPUx52dGl7u0/PiTCpcbVT/m+JT1MYqby+H1QdOmC+4YP+c/LeS+3Tsl3yt9eLg9F
xylu+IPTWP7DHok4cEsfIyXS17krgUHjPN0yz/MLhLJch61r8aWRvkVUchj6IBeXWBm4rXu3ZUSy
x9xnxgZlogRjSfLfU6IPUIVlspenTyVqzO8mixAycSMSNlwYUs81i0e3DX/KEqjvOJsljuZM3G0X
X/nWOcPR3xF/aEn7ijRlOCWTPru2TRprwUJoqGV59S/x4W9yvWZBdYjClWMzJkYv4M4d/0HUsg/m
jSPtoDtWxotHRhIIueN6l6Qvq324jb4Cu+Oz43PqZut8tdhWxd1Z0B/0szSiDa+7mzfLxdK5KazE
+75NMW9SWGhojQQRyPYe3ilk6fWrRHHIENwZb/P/tT3I3mcP/n4jbKgQFkwOmvZmgYbIYUaZoUp+
xMxG3m2jj4Tp/DTRzgbaXyvk/iQufJbbgDwaAgmunBR5Q6mPA+Y8AOaRNyqEQ+Kjx2NMRH3xBA4q
YRQGkSTblYtofIgsY1oDk/v1PqdWYW0hrYuUhAtuy9PdwaFQch6EsOB3bN20zN6Yta/sclqXIwki
UuL2qYc7sOJUm5br77zrCk7VETo5L0GPMIggPO3vwCi0hiHbL8sLeiOza5pVHeNPbl8oX4NENuUt
/rBxFYWbq94r0h8VWjakNtBq+UZ+pVS34RPZBAq7VvfVqzL/1dXasGQMrUw67wfF58AHBMD88r0A
4AiY+1L3CjD+hdTnx3C0FcJawEhN4yGvBI+soojIftTnBM1+ovdNr8P7772p/eYnCQCtssc7+D33
99Tb09Dzw5WUBwR8vSbbQWyQPwuVC9y0dtEznUpoMQ5p8FJgp/WaWVy9y6OFnGrFyRDhGlqg/0hc
tsaDgzL8hZ8SzMQUXCuBNA9NnwY29VfjFA3EfrPayU8oVCsKik0UtZaQvCtl3sRm8IG9XiPY7/P9
+GtwTdmrcRatDhMuKe4ZfW7qAuWHbDG6nhyw9qrQX6rcXkL6AcKSCBeDVw3I8mJR+DfItpHNjmjO
0egzVjqcQ3YncoLlV2lT8Znf1adKII4NwV01quHTQaHaDoFv1OMHrfW66KUeRfrC87LNh3sU8rNy
afP6u8XE1bNikOLJytGzmOXFjo9pKhIoPbFgGMV9eiTvJY/etFJZ9acyFBqpy9Og+Uo2u1nPeJP6
3cExruXZh4RJX5X4RL+S370MeyBYZQyEbZ3uLV62/xjr/j9RyJutUFGNqQ3NoExbIT/luwQMHBAl
7QtrSacU6ZvX3o4O0YFW4DktU3VgxdYs0gLhfw+Ca4nasP+3aH0kCNXTt+c993IhXs7Qmy11LX04
Qe5BlHthRgQK82+sMpbs2566co1YbLPs+o8h8+ojrarDE03XUvWoBB2mouqXtGTn9vs+9FVoMfXB
VNzD/iJ7Xd2AfaXIn0YhcG4MuZjLIjhnUcQLv5Wx8P2i9pO3CP5zHkwH/dSJZdA71C300HXurG7+
cXa8+2Wg4yoH/kLiRWjEGjhujftcjt1WJSEl9iIUrQlu2s5F255+S4voVOegR4ot/C38WAR1A2UW
yrS2nk/v+eHQk4mcUZ14IjSTJhYnku772FMOMBYRGxm8p25Oozx09uyAkmvdNsdrpLVCXkl4RQ2g
EQ0MrLB+mFauSUJPxCrFsxnFM1fNl8ymUqemvm5hOisbHTvwEe7O+cVSq4iGCWRW6mR7zdVESxC2
2vK6aBRw99FHT8E1tnIK3Rima5kqhWInaffpM79TgbPyf0K51JAEJrtnojXMoTzd1zFyTueOdFd9
+mN2EQZ9140lUobcaVMQyQvQ28MHci6S9poe0CKoy2WkbaxNSSGIL4tqrfFZs+DjhDRLVAuw24QR
Is0YgsslYMq6pcpoSjTtslNGss4TQ9Euz5cwZtjuVLHiLnlKVLXJm9h62BfwT4WZPjZUv0bgaprR
pTb2KYZWp9tyaot12z2iWPnssW+UisWxxAuJlHC9ULtJzaBSghAelX79peRDkPl9yv97W//Cq8jD
L8oSF632dQlvSUmBYjlc4mMoulEoO+iYh4jbueu3AAiCTXMZjFVdcsf4LGsmuj6Po0seuIloVXOt
h8z+CsgqG6x91pWrayR9qP7fjyzoYumhmJfw7QwIbV0I5SDAl1xW7J4ReHusZpt1HeogefunTtEC
ZLxLbHi8ribmpCZwgl9b+0KdiHNVdXA+Flcft/1e/lctLjWhzzw3svWwpA/UiV8/XHsTGTphXtR/
9EU/KM3wAh+3X+pxGYovldTQtyEtQtv41limJ85hydZS24GTIvrI5w6YKBPlwfip7QKDSTFNOt7W
KK7N4XsTIgxdlnYOmDCdZ9NTs+JBu91sYXmmlyNYHn1E6GIEwPp1fnCuQPLVDx9755IkDyzdOXGV
HGK0GWockwcZV5wDcpajHSKDbBGl8KqA/p5/xZn0jgluMJ23V1H7lwcXEEnC/3QxGxopFHKoEmA2
6P2xPO67s+UZ/35mx98jI7RSeFhS0++t/nmNz1JuNbXMVOflWECWF+JWGndUdXG8PvA2TR53PoUh
MTn43eB0fPqfUs+i9UXsLgrfMIbRpInn3fyyPgS07K3Z/t1BWQaDL9A4pEZrTQ07ffvfHqEY+dwD
YQnAwurVIy7C/wpzZscOTcf97U9sa8aDe6gi1h+xFSWhAOHP2f9gDYOZ2zj0JKNUqwQzxfTkEP5V
fH7GE9IOJLKEa/T31RdSHkl9Sz302rhzxTG2xuDCMONlTNZ6iYc7BDu0WHk/PYGEa3vgtpxDnjo0
czArBRR+CmKAOT+ZVVAhxJ87XQ3yJVCY2vC27f1kn98NfnsUunOsdyWJZAPGZdoW5H3oJHzZMSCn
L9itbq7U3/jFf00PTzLYRe6kYVJ2cGvqaVXfIedfh1UQZ/dmvPN1TFQ59Ame24JP1VSdpJJT3PFW
fXJuVXZupxmu+p84/2NOIc/fwgSBZ/2U/7IV5FpdeASLFZAPrsBYYYruIWeLifUyV5c2kzFGNAg4
8hHbPl1CBAjQix0ADSZgFT258dETOqt0tv72NyqtIqfMLq+6fn7pSmPBsJHEuLs8yprpbZKoU5Q7
/KUXfH0iuN7GNIUB0+PbNhvxu6aWwjC3zJYFpicHindVqrj2IfzeoceLwDL4ziUR/eaQY66p82ru
Gu9Y4qsWQRiOQSBcVoCfJH9dJxYMeljqq6ZCc2acw2WOsu1jhPwSw5jY16I7HpKOc66YyYpwxeE7
UWWUSBVD9V1oNNf0hLU1jQSCpTImb1P7167/rhKkLT59sz9zagQ+0I/LHdZ+GHtBJtzKJNK6rz8P
zSHKqxIRpbmxENU4ocJIwc+m1UYprpmpg61c4Y2r3IaJG1kGh+Ai7XNUOl6M+Ds3MMkfDtbVQA9w
CGstdXMpyTOqOXOYXQItvveIhfZUTqdAnsl4eNr//Xa9DixeYuov+qJ/vm3HsWYr5BImyUOjfYI+
HhbiKt8XHTLh+xonBVxTl2r5TagENiTdMOKYR0apUsDRwwuTgrGHv8LcyIszvg0eaCutPl87QZtO
Np/sCK348jiwVtJHIRQo6QJ2ctdY3J/3iMS6rfaDp1FCq/rM+PB8iL70Gic3c7qqswQk6WVLdYTI
HOCK1s/tNk9xk1Nm1Qy85c085jML6nHPx95CXxgtfeTEZ9tox4uQwDEikAM6Oa7ARAFGkguzQGfw
oOjZTEC/Qrfq5d/b/at9iG51I+DdtFLxZyT6RXJCuXiueT4CAyJCAbXMU0NBaZq0+rdHSU/E6yao
eoq7OngkPACLlgOzsdZJsNzWYyBG1Q0plHGUIScxpg2dI49KGxST1gcXn+VdosotaPhC2FinlCAM
jOWlxdtoidzjMhCzPrJQd5TtoGh3ioACcb9HgN4Nd4Eofu0ANdeDGRAWt/siwbcieYUnbAbFlOoh
v/Xq+GzPqVDx8ZDbvGVVrNB2GyGt4KLX0Ce/hFAtWooszq59fU1ksxCoZjpEQGkC0KReRz7e0izU
z83HCp9YWJLBMyDRd0SKqxY8kJfr4PfkKJVJKvjh2imHJH5rcFITeewvgiZ2sFfssggzrJ6PJZoA
4qGHMzq5gUluz05Dp7lkEIzJq5Ub5yo+eWNc4VlRJ430zjyuI5eDRHAYUUTtksEfY8BT0EWfbXRz
0FUHfijDejNnsRzzfaO2SdNf+08lWUxNwAaZtLaM++GGTbQQyeBdRQYuKY8ObqZuiYz/qPWVkKtd
l3ZVg6tvVzevIsh8bOZwaHpXvSFnq1vYCIHpwcucyKX0iIU8jiSALTXWTovE1HJxl62PEDwAZ1Qj
FcHAKStnEMucyq/B5LflcwBQOXLHQ2GglsBj2byFmOq4fuTYaTX3Q8TZdXUUfxgPpFjw1385rLDL
dC6j/JPAhlynm/jERbLd8ySPEz9Zr2HO2n3KCWiLR7KPzv06kPTB/IWbR824yoC/XsBsuylUq278
mUHLRYIHCXL+M6oKM7QuO3Nd+BDNcHotETYD973+qXKGes9rWTsVD+iN/n6bjJkdT6Y6Ag6oU0RB
ClsDJYSukxsBxlzaQU96E/7dJyfl5wBgyRVl6xAdBjVGq2u2edB2MHSUaGgK5dUT2MQiotD1zSNq
T5C/YFcXNfKhGM+jZwk6Bvs+y0X8jI0Ixe0bneGTWcieL0zLgLbVt+NfA8IZdC3Fo4I0YIKG5lxS
3GCUbFkXnVeZLrmO7HVWIeoc4sg6AMmg9bsVxsQxJYoKyiNhp2qSyZk1HkmUkx494MijtKWOQrFy
DC1+mSE5NGn8RHFt+co3TJIu88q1wPL22V4vVI6P242m8GF6GlGCGBCqGKn6V9yjC6deS5PUxrkM
xX7+ltOkGZtJ6yfBkac1F4cm+ugQDCTq5lsonDYlRogD8RIuZ+wny106MX/wNRp3uBSbuYX924Cb
9Pmrew3CdjrKKoI/PBgGCdlVNt8BdbOk4XDOEylIH0++L7e8H6knBdNA+R87bjNgHuIa0Cw1DPJS
rbJOArzN+Or+xNl1KWe0YhWgl27BBczwfWpg7KEbSS8GLSBnXQiAjgT7lH6BZXKsxerCe/nbprCQ
zp9ST6GKCJR1v7lskZDeJUhfXWr01YSLrBHANPtnsVxLKHAE4LIn+/GGvfxBjLESGuwvVZxnjsI8
Wob4fb3BgN02eA/FzmYII2Pv5D/VHDBsCqn0zAdZatrD3PY0Nmz3NAhNm+gfJLzH8wGWq3unGpeP
Oy2cE9tcEmsDwaE5sYcYgoPWvIVK1WCHUgzHmaAhpYZSO1BGoum7yBUxps1/ssXPRYQSKQCJlmBX
wRhLG9iiY7LGLDNiET6i6UVZmLHFpSmN6DWuxhpT29Wl7NDcM4/N5iY8I9yxyt/qbWkTqRxxBUSM
7PiC/dd3y0RcJqmzmobREbrSDRoD0W5XBUxMvcoLMiAJDYQjHe/I1sTRvF3sPVyzVO4M7to/iJng
20j8bNQieFDponDOesV+da62M+FsMjeTcvN5Az4Ww3TNlKtm3oMlt2qcboyYV6vtjSB14G3uRqdZ
b4nGdOJfpJUu8RUAlptPxw3UMP4jx7rM32ppidU3TD4ZxXClNT5mP5P1bMDWXavpI7BUuMkXa01e
rgjr3Mo3ZYTIZHJ0Bhe3WARBe1AxrVV1M67A2V3oRbyTNpYK9ziwhkfOYLThhIaCSGy9BYAzHXvM
KpnzfX81UxVV4y1nw0fEB4X3+zo863bigTXCTvLgZ8V8Ou+MUPylcaDbkg+5KryGxoLCI8AHfXWA
OaSmv7ESTU/HZB7Ws8Wr6PuYFK18r4GwRI4rwDF3INcsX/W14UZOKi2JP2q/J+wfH7dDjAFj9Ydz
SUMjNda1MCaVpq4wGz3bq+MyH9WN+mU6R0QF+uQDdMW4OCTRsPXwNhIzximdr4Wr1hoQyKKooxwz
zsMgMiTJAGPLhBwrc4GnQkE7V3ZccejgPPU3dO86iX8hFAiRw/NWG0fJzW8u4Aw+Z/DODyiz51Dr
k7GD3/L5/XV5DjrEHe3/pR41WwgZ/YigMed+Xb+1kfeU+g5VOPVtxvfSaJzQZl6pUVJdpsGIeySy
xCJ3csQ24RGXEVudxbXtQAfTQgvTMiIXUzF397Rr/LOWE8IPtWOqpLuKvBLE7GqnQvG0vixmyKrl
srhQVA6/mnQNpvQBzh2xG50lUFDC0zE8Xjj6vfIn4+l6z46TrEPvFNcDai9CPQVBspqLEZAMa3YC
u6qaXkaE+miUegWRw4w8NZVolnW57NvtrM3pptTIEpsQZjWKI2O7DYWj0IWgAE6n8HD661OVPDQ8
3jMdE1oxlNVR/9Se6Z4eQ40FQKqpRkjVBk3uHdC+c7yzs5JIsB79nh0jr/rNXnhXifc1NYkopHsl
9akIGeM7QyEcb9ERNOiuwYoSnMlWG6oJ3v+5lcKOWkzt2/qoO/zS0A6lyRyfCl7HMcQ3iFCUxUJz
vv+JI+fkZ0g05EY0PA3bGrAyemPU3iUC1DhGe9BA9PBItcv14HDqJIxFw5t2D4joo+AEa+Yon5zR
zTHHFml0KPraiplejc+zzfPIgFAakqwvcF9LYpGRuloIQjeOi/tl25oyAzDwmLsYidA5gvcdf576
j4uQFFTVVzAAKNldr1I1JnZ4agtfb/seGCzRv+lHdF0w0/Vl8YmU1VHksiVo1dz+Y5yu8aLrjySq
VKfygRpnZ6FhyWdW4gREAMPNyq3t1cfR2S473Vf74/ImT/ertSnFvq1INe9D4eZKrpY9SJsHXVen
DrBIQQOq7xFpSZc1WA8n3YzzSv+zaNuWUB2IV6diNchytBHDTryNAZQ9xsLLFCgFmX6R5xncEuMz
6BUf4BkswpeWrMpk3o2Cj9bQIDh+ODPpOaKX/+2Mjd9UNzHZyFy8lOPiWq+txkr/bSwBIqpIPBQ9
kej0QF1qEb/Y0NW9wPCZMsJqblVCPEGlWqmMvFUuIHg7XvMCcd9iFvLGXP2vhR2JLJeFkgxG0gFh
FQNjOilBego6XdEeLPPcGuau0ZxQ4zR9laSOQ3Z1qJma9Xbp+wOm0XvqdCbNSInm02bRoEexB2Ue
5bDe0egSL0TidtFWJ/3hF30pip8oLa2F9wfD1D5zy/1OjtEYYueuCs/a/W29SwC/uaET822rVGXY
/rt0wXJMifacpEsq7+dFHB1PEGdcroI0xEhcR39x/RwJZj/SJUFpjdbYEUyWMq9jWm2LY0nMSe4+
VErVDphJUfFPBNlZBYNoaPty8O2B0L4cPXEQ22DAmzecrGkWaGSoAosHninFCiJ0x3P8J0+coBkA
Y5slQEexMvJHMEBEMzGURl1Qkfc+JRrXD9L7i+1XkogRAl1y5wBbcZ+QsodwrHrvP/RkVR8uZoVI
5iks2s5sOc2OaJJcj/Q1umyFrYHZlgPDWXa0xN2Ps3IAsLAExg7+VwCQhebr6TB4Ea3D+cOVXeSX
JyalWCfIv029bp+nISCAMCb+knUfPri7GAV1PwtGmU/3XEKzq04QXNBiYy3Bsn0ju2lOL53R4hkM
+QzTom2MW8lkOdpGG4hKbJ04wEUutHw9sFbMhx6ZYKbly+C2ErXYdWx6w3UzWoeMcjfl5GTPheW9
Lr8c+oyI3cDsntUXnH1RPbAwEjwcNtvpxyanT/NL+YWo5kQ2/wikz299Sy698oOf3/i0AKAxRh2w
S3AUThzhWNBMrK/H5WTxvNEw0sjtAvu/D2/aSNt/szM0iisx9JWpF3LPXdrHv6NPJHnBFN4bsTmZ
LGMvZ6hjwVsFO6PzIAHleKXEOsdf1GEXVOvGo72PC3rPehxlAROaSqb2gX1dXDL5RBacyJ+Unuf3
mFFeWjkQ8PclxSWrnpNidTdbj2yTsw87KaSJl+kLoAuKV7XJaTPfU9Tfj9ugjbNkzBtGqhnzbqSN
lneAkWC+CW9CqAL2WOWF1NT34GE+I6GmgEyAVpb9eMUDwM4CtTFtb0po4Yt7crPZNLMJ8uO9ufVZ
3GcKVCtiBqlnjOAxZejjLF4WSGZr5d1N1ryzIgE5fmiH3Qngq+XckznE7qJ6P+WrKtnZBpjKU0I3
x/dLG422ifkcSAGgEjseyDJorQ0IUVbd0fneYqVra6RQgJqy9S759KMfIAgP2CWQ7Ps2+sWhlAOD
3qi1FMxsRuYbqeFV0agamS1lTkRBY2P3CjfgJqrzjGhZXAW2x8hJObcxMrZiJXAfhaMPzXLyrYv9
C/nHbjUE6nQaWDiRzYRobFAtQTu2WNwtWdc+iM5pdJE4Der8+k6/Zk9gwXuzzPTHcLzlx8hNGhs3
sdWSJgzRLXhHTS0FsvhAR/fTHn5xw8/QacDcyn5WZi8W32HjXF2huCeOLgmp4VXwKJJ5J8zbQwBJ
kpJTV8B1XYyNo9S6/Q0ULvwtlsAvPM0GFFg8r+l4E5FePdUuB4u5thekgSGv77IfVWkmDfBQ7ryo
AMr+7Chbf9Vuu8UJ0F0ZnhvyK2RPEy9bgdmJ0XhQYulgtWsOaS/hSHwPVusF9ghe57Ue7jPPik7F
uQwfbWlMrXCl8REM/GzWwld1rD2dz37KeBkdSfDeGyfYBwAwT/ptfhJNHgTcxbM43+bTqqSGZxTD
oNhNyavc1vPaopPNkS8ruNOYl7PZkxcfpCfFB5EwWYA8b4XWCQWR46b8Fxfuovs3zrr6WcJkn21n
jLuyTcaJJCPmgrDwrAB6gTaqlQ5QQ7B0CR4YaOcZU265uGDEMBsOndYUP49by91HCsaMKVrHb0k7
/xpq/v7BeMeXxhHIRMjm4/b8WujozW0CN7/6/J5Mxi5om68DG2a/ZramKPJdWqbMG9AuvkHOH3Tn
4C6mbjs4NpBscy4PaBgm4yQkIFDfQKxWhg711gKgzqV3fGqPHWdunzB8WH1jn2C0dlah5dKWMq3d
wlCOFlf6bsiYvTgL4GVij0p+Coz0b39nakU+kC6PJjW8ejTDKw2i35yyookAFtrgWXL/gEADZBye
yV1lZaK+DmJj8qge39tv/3EdGgp2Ll0+eq0x8wDu2OwUcupS1honVM0s4aJfiIYLke1PLCcOTbC2
Q1IOmcWFT57kSg4aX8MfE04jF9pc5aJJ8eqE1RipD5fBMh87RhlTN0YeTYaksbCDz67y02nbJHp+
YeFjghG7AsO3Jkb/UQBmgnfYX12x1FmI9QdH1FcMotdxkgYuUGmstB+hHXYY/he1YFHgVByMC78A
YsNBtgqKglAi784qS3jmLZioEut+Qujaqp8/e7hYBUxZkYIGpWxrzW7C/C7jmPS9Jx/6TmC9YkPS
AOn0CUu1YwLkdkVsTaBuunwRqBIp76DH+gH6Byezw7YRf48HvehFIh61OKOA2yykP92lUMDJsJB2
UNGhDJw3vMbj7ojpxkkjKLo1KPd6IfNTmiixIYKoMR4ZYQN7U2lbKO+1rv2GwzsCSt+AZoy2RVt5
lBdqo9ugyoLV6WnTd4MpK3sI4YDt9mMePhy3xUK6y8OP2EBzZhy66QE1QlD3HRymPcnzfub4GAbO
1pMI5nelGCby36dMi6356I66Ppp9vbs9bLV7MiYzT77XwsaBMjcWZ/dOYaFpRG0XEupMoSLP+I2e
iDDLOT1h/nbN7KoxA1gjgun+FcynOTpuGMUqBXFGkEGnaozDTWKAz62uwwucm/Zo0Nd+fBSYYUvG
MzFItK3rvaGExvdOknPwzBB8cGvRuP0hxaxaooKBs4cqlw0IlH2QVjoINYu5sk8Loe7qKMRszYFC
TvH8nRc74J0ISU0uhju5gS6fdjbtBO+lMzIOdF2XJKMkdowW6zjIUpiVHbZ5kQWcS5fA4YY/z0Fs
bme2zD048hfwfZA/fjDCTWq0kmcQq/g3HQpyGJcT6/l41PVajoCzdq85Uve/mQAUJB5sRKjSWp+0
7/NkUqI5xyG4n8meWABLVxJXRdqXRZbGbmSp2tB6uBRzytpjKxuO6duwgq7VSBn4fwgALJL2OkZB
7d2O5q0/rfnWNgRfRxXROIAdOt92rWpgm4NUJrSDJz7OOK1EaQDh07aGgxhCg4CROgF7m9X8pWu2
u4C/XaIs0TW7R22xk3lUcVqmuYW3F+KmYTKYOEMrqdoXOKRd/GNYJOzp14MhNegXOKPK1pH4lSGR
QOdy8KLvITxnPwDsi0ZaWzDOLV+xmWUBA7/0GOIhSEQdbSZkRh1QKz/HBt1e5f/aVE3HvDt9DsdT
wYPS8RHl7jUVCvvjEvzdF68O46eSDFWwfMy0oWThdNLV+3ocVMoJBzNxz07SA0fJpd7Ax9NfWDbi
dRP9Xp+9mRa+AD77yBlhIfTVxSmkQwqjNIwuCSv7ZpR6YEu4T54/ZSKf8d1LP3sl+TY8ER7+C7ZD
fkG6xsTfTaKIy2U0Nq1RpoXnlRPNS/PWmtcM1YlPgC/lZvCerqr6wpg1C48Oec5X87xDBh+YpcHy
nFEEyXnkA4+6/j/XN8UrCnR+P6azotLsi2kfmem2FOh0H1RV9Y10JK43k0RtEixwmx9PwyO+7pFD
fN6jC66OLPM4g2m2P49X+uXQgUMPZ4qn3VAUsSack9pq09D7JNc4BuP6ZmJOrF+5IF1ahAVPl80v
B6NzIufsqMPk/0XgkP3m8Pz83bQFjqape6DJRnI/WT1hgMVKJxio0K+oKVhKGjlQAhTnKQM0ZcGP
Cz44xk4RyF00RHW/fY+gPejColImhYqhcXW+ClUPnyWcZl2+FikgFmv8TKfGeM6vJRKsrFRTYM0p
4hVuB/y6GWNtSdMmUKFigbxbbX9Zqbpnpu+JfTiUcoYgKIXfi1kKm8w0uRhAWnbyFxeWj9nj8XXf
JxyOP5SCjQJNFUEJA53/b0CdcqCybEbF1gPu8KmNa1hqq9WhEPcEeVo5xlRTmsHxLshfrVKoG28p
fVaeHXXlelniSQOnJXalIuoSCBODaYsTKhWA5i6lO30emZNPT66eUYnTJbXsHjKY4TD15RoJqEaV
eawiKOQBzyLeuhXQ35JK4VV15nOJlWgyPaHMwR/RyxIQ4mg0EkuwYsTACNAd9kVtA3dBu701Tpvg
3aRpYzccgltW3pMdrTmHHodLvBw7/5ryn67m5+POEAVu+V7gRVpHbjAhMFXEfhVI7AHtR5RNqa21
tx39MVFV6tmxiIVYOODj3oH4C+Exrd5PzvijrMIU5aISWpTcjI/MsHqnstwFS33aNibgoq95Ce+l
dPc+oQkY6h0hShffYkiveyX+b55bxzbXJB0VaTOdmPLejCkkTlrsM4pTBuDErYg/ds6+m4JEt2gy
kOLi0+iZ5hRmSlJBZTuFogXY3LoSer4fXJcedLSZdg0tMbp6frJI2PIzHeKr0Z0wB4Ono1TP7s1T
WTa4uW27/cw2/TpJX6k5M3aDWtXZrKbpQepSgFg88FbATw11Oklce4f3f/msSquqShXE4Zz2JdJw
paeLsuGP8BSxXKX/UI31/3KneloLLQZ2A6z/bEOTW0HmD011mrAtubAFXUfc+fycdiST/QdSApy7
SuN5jrM4kOGeSURuPj/aYNHy8HeRlioKgOjEM1wFjnJU9ddhlIzoOyASaNw/G1taiw755qqwo2ug
S477PHZMw/G2HZP0cRhs1EccXCxWEpHnwdgQpH+LIJDcdEzQrm7vVAtx817zAV/bHdYO/gFYuzXC
yxNa/nrjxbkswbim4S4Xex8Ezw3FBZeXLH8SCPnwkEwjbRm/KTeu9psJWGTfHadqE6k1ku5kC1kO
S4S5lhT0PYoGihkBOkwQncsy08feCM8pS/uQO+BVNrEwkQu/chpr+2kKkVbU31aRenwBqIy9mJ5z
ilkWvkePCWVMQPvw4RbtT7Z7BPo9LuMj8AbQQ+eW3MOEggiinKKYMCFY70Wfx6GgpDC+SQ0Nmvw4
EWLriBEMSMzrTOFDPLpB4ZVwPN2hEXKwuz3+CxqesMoklhsTF+L9jEYga25MjJD+AAAjuFDU/qp3
cwYSsZIv/m7Pf08tNgrUTHIOciz72EQy4mITCzcqL66Vkq1g1q7IZlNqTZNO1UCjo37aBQl/r0Ge
t4Cw+dg+wSs8r1rKthQbow4ucHXJakQxxEttPiQ4UzvJINu2gjxhO4rQoRnrR+NVE7N1i/YT8bxa
YbxoZgfRygmDDMaRAqxguEvjVf8cz+fx197msuPGR5kXHzzJSvlg9LsSYi6cSufglgmjMklMgFrN
aLbsHv9BUrd4brnOwRMwa6IIBtczJLLOdzEXBsrhnLMraOKKUcSIS4yJfuzL43pSqjrr+Ra0SAFa
fd/9a0E++UNBM1q/tUq1JSPnKH45/EaQcHDuxMcKUU4JbMVSjEk0kd7GymcBWBhjUeq9Yzp+3A9I
+syFGBZ6BKbvUehDiCSqDRUHthN+g2ykfosfkdePkt0rhCpzWf1R3lHjgjrAP9hL9H6sYU/xOHOQ
KgP0y0lhlhQAlR3fDXMiKmgnam7SSxzEO47V+uypE9Z9UjUgA++t5pcq0fw9ZcsmbwEGivfhzq+C
1weA4R5FYWCiqqD0LHIo7MZhe5WH/2iDsJf6+Lf5DEES6xwpJheggD8SXY8jLRV/PA1vqYOCV1y5
572bFNCueGkg57W/Q5GrcLKR8hD73uMFoBurNllIq0Pra+ywHyYS/EbgIoOWPPr3KvPy7R2aOcsy
+KxAJaCMUuGFiL07m+8oNvf0PPu72l/8Zqr9EjQL78fmv35d7kdcdVqvxan+V7NQ+EOPBJLqdHbk
60etlLlu+fidaFQr94U09PVphRJP3z/Mx9aDEgtmsztRSq4QiBh/S0vsdCC7gdwKpgXMRAccRsHs
sXcb5c4vxySmyzHPl6pRKIEGpPhTGdN/kMsm+8wnvRXC0BH0exPEYiI3FPFZ1ee1uaYuafKv3mXM
595UK550LLEQEbEU9aHFV27ajfqLmo/sLnY9mVnHt6yqA+3sEqv+Ct92oEe5gFfFB8oFIjAGbiMy
V+QOD6UBJWfKpy1oJOKt7LqrbRS7F9yzmZMmUjgaoK4AXSgU40g/zsu9L84cHAZp2WA1bbxP+z05
S+pzYQjFXC+amC9l+ntoiqaK4paLlyzkfu2Q6msjm7OZiZjz0HMLkkg5SxS7bFKTMkUAodxXOe+f
dSnA5Hq0OU4DPqVb0bSBExNnGb4m/n0JFVb84zwrA/yyYJ2/DlVD0VTONITMCKs/92Ahd/6RLKiZ
WboPmfejYfDQM7eYsa+lEb7wn0yTLvX+AG48egZBNq8/ZiY+8HENHMV6C4dN647Qgrbgz0eaowyD
9vFMIKqlRirXTS1ciRFAKn52otE918fOSSByfylZgkKXPUzw4TUq5Js/Kqh9SKyw82RFdQFZngww
bzJuBOa/8iFj+mtRISR4pT3l0g5ulvCWq0SGdCZQ05uYUBmsIzNj/YZQ/BdxiJrntKNFmKi0WuBB
TPed6cCA2vCEox2z2aSJ5N3wGeYnD5iI2QDBvNVrvCydnoQJcGqljdpESG2pvYbKDF4WLa7ViCxF
JymfLL4PDe4Xo7gg3irIg4etDZug4CmrDaSK1cC4d/mMB1SLMS5UskCE6Ra6rwtA0i4MqKpr3aB6
tZvbQU9/zMIwD8b0G/71sgzmLQvC7jl0sC7AC/ChP6ZugUQlm0hZaHdNbqkxajXyVlgowdypCC7M
cOv/ay9cJnFF0zjLUkOWUUd7KRQP8htNWa+P79ncFIdxkPXLZPjXwu72f66FqsqCNEGCuxujE8iE
UtC9fo/KYFhAZVs8tRqxKZBOBzJ0AXcitmOj87g4HBr08n3tAIoCLrIbRQL4Gt8UpfQlsTJyOAyc
tLmxkV7bBsypfri3h9Nc7h2HHEWejqPV1K/FRgPrCdyLQfECE9S/avM4H7wnEJS3VYnx9sn2IjTW
72FBJL0tynrYWtVGlcNlcubr2ccVDAEPDrrLf/mv3I4nlp1ltjYT8X04PEVYLaFjX+hnLPCS4Fzt
qX+0gIr0Xr2o7FmkdoU/kSSD68ML1qmWhewrxugRowBUv37rwMhnixq3oIiy5kmnmmLVYn3llYyb
wKpFE4Jj9X6cl587IOavShamlzj3VWacqp5SE/LlDgVbl9bDA7shVcoFL//SWR2bq5E2biYDouRs
nPrgu+UiXrQg1Lc77wqUcSMOXuP4XfOzARS8QydjlaDTNRC8h0FCyfhUiaeVqzGGJqqGYt6vLWXt
dje9eRJRBg63mtl+31xRlogVPu5jJBOzBvCIZpyD63U26thNa1r3/Xzzj6xbn/tUIFV+YkxVyFYN
4yqtmZ/4p3z/9R4y3P48FK6WLmnY9FIritz4wDiOOXPYtMK9sgjQxPsw5ZNaNkImrm+2veVhBWLF
AjGnIu1kAL/wMRfqacV0jcSO+jDt6hpGU63SlhQFoTbxY/dWxxDkghZbM5dsjGy0lrNY3SPZbmUV
9qCONuCj/mNw1gceCAr3cUSYX+I9i0u2036BPn7qI/gWZ1LsxtIZD3ZwdycLbkM2p/kjay73fKIl
S/BfvAgUjN3ReVnAevbubioTWjOBDmxo5MILc5/+QsvrfhV6xtgNYFwZj+UrljBEpsdY8Rd4+9Yn
Te84Htt6yxZvoHKZQ1NGol90tKbBUIvXraAHabGpLDNnqw0siZFG85SJCGpI+WUwuOU930l0kv2a
5kG5MOmWVun4nVPd3QnGqv3rpQdQlCvrYyULHnqvcH8G6LawXXrv3Tij5zdPSWxDsKimLPQX/wZ0
EnxggF5Q/uPDuhFyhlOq2QOsEzlGRWOjwxat8fzwpaNmY/5ARpFR58VpRoxLGuuP1LDxTK62s5jT
AeZmDoUT2YxJEyXZLxjl/yV6/irGVwgmWF8/JWlJYXzWNXl3yFJweDsua8lMCV6qtWn88v2MbdDs
o23ZShb1e7N6Y6ZTzW7UWkn3g250kP7L7rxAoxdZQyJ2n0L3FgA/my1WThCAGevcDNoORqZd5XmY
YCkeLjqj95vRh7P/kzbYiQT0k6kW/oztKDMb2N8AOkb5lEAk4rTl9i+S8Vf534/LUjtbbvW+GXY8
ZL4p0VXaYNmhDejvtFUcLu+2YuCCLRgTgzNOnh3IqOmI+0PCpuxvft43H5IFLY0Wz6nxm14av+q3
3EVzJuw47VStEblBGxvVp+V70txwz2RKFn0OeuFimlZx2ZUHzTgNCHjKKT43SsRGkstJ8JVkz/wf
ANavP4Qxag+Yeo0gK4JSiOcF/wTE40+Gd+GMHGxmvlycr/zkDPVAaGIXXby2EE6jmXgXGbdWgP1l
icTJ6VxaU2TWlDicMVDuTP39g/kXZVZ0G9VA6uUc8vaPEawUAKrlnD8eV0rfx4nyFyOBG5SsqSD2
W97c6ScWKasKANjP29/Jl7Sq/+rNAk0Qd1T+F1eoWawbRblyk0Q4nhiE1GEiFqt+weZlvStfVgtv
1wVquIEJU5Gp07cILViMEhSgimx8AcvcQgI7gdJab9MfJ/E7BAgE5rs5fG7OLPbzVJcR8d9vUefl
mevPq5oT29AVV+jbQWgTkBgMs4xPC+Z8J3GBAu5N0TcxGu5SevpexJe4VAsoNvP5qZPJtStYaOiI
wL2oelj7YX2CMgGgR06pgtIDfERKgKdd2yHQf6YbnIemKWa2GCrii0cjVFzh7dbcoZogvR2pamTZ
LQYmNHGsV72NFezzA9FPFBO0bTWeVaLhHq+TM6XaMVY7qqCW567KeGeek1We8AnLevFrFKIZQV7R
3tbV18VEznKi022Bb3EneTlQAODcbdOoBOYu7XltW6667nUo4Wu7NA+JFmiYLFgCy4D0P43SUJBu
uVjjKuD3p1RBh7uQ21NH4sZi9IrguW6H5U8K6MPNV1VRXjfmRI7WFEgtUlPE1mSGmVQMfVO843v1
1Tz0/mpowbinNPVL+EpbQkWSwai2q3CA1cmk6i/ZWe+lsbzKiakWnM66NQKuDEOSwYFguR4G3Wby
7sbmvq1+sG6+atyy/uDkN7YmuL3/q7fF0CQk/KxFHozU1QvdgibC75nECsbcbeZ7kHM+7wdt29ro
Q+oVbLBtPFEYXeNK49tJe4G8BX8qZofh/U4z60OBPbDQmBInJJN5jLBtI/JmXLovYf1rEuh2kPQQ
dzhn2u0j/moyN0rJg1L5u2g7ndNUAJjMTBXSTt5yoBUAyGYCnAvrfUAmc3vcnjZ+obft5h8r/8Ll
P2ndzPlaeEtYxNklqdn8HOifGtg3CeL7GtLvdzDPSMEFvmv23PougjodVybznkMFqw9DDiRCBkYS
PV+lFVtpPpRDB9jnGtmw4hNrZWxVo/HoGiMZf1ItR+dUsA+vWSDmqPvQ7np9uabSyvChO4VF5umI
FttMGeMmtR9Y2b5Ba9xuaNaqqZd4lCiICg/jbX7EodSU8qK+j7fMbpTBI3ha+RY3tLefOlIikAxQ
PRiDDvh+rCs/kbSOMzTe00NL3ruHO7RRSDr0gXUqfCxqvGpabcazUiOKw4xOvyVJ+1dcgXH6Hld4
lKmB5rIQPfTJH4jxu3l8Bw2SrtIHFw3eUgoM3dMpfiQn7qeEXRc23jf7rY+aEUJApeHEe/cY1v6J
t5/jyCHZoSHzr3G6yr1DsFkSxM7rLC2WrZkIaedxXP8JzK9jtWzA3mlAEcHKZ6zNRffGTKFtoB4p
tuKd6enWi6f3y26lYoeiBhWF41bO9JS33b0iHaEWXd60V60kIdpQctUZyVikY7UqQX4+NTJ5wGfD
c7elyKyB77G9s2q/8VrEZvu+qPXwbqqMu7mzfDzSpINvtAXhcA/hKwHVHmQdLYG0HCPod8ExapCD
63Nn0lV+eMaJanBn5zGTBkwRC9Cl2HdMs8OLP6LvGwAKSimOJuk2kFty92tSGekxxrmdPKgJlajR
lg/eDeVECWZZO6lCrlrd2xns4p8OIRrN5CDgIlZYBgGOL6z2QTqBoIKXs6LS1OBapQnAdWWxoog/
8yCPw1czXTwA93dBLWyNwya1dFePxBmbgqx/j6QV0BdH4Ql3FaDLcoB912PjPZSIODty9OxBO9ue
MN/bz6Kb4v1z8EMPmDSFnlYKrK4tc1MjyrAbtX6adx3usRU8+MLivGJIF3aUj9PcMJbPFQEm/PdJ
nhktbgVsMu/c1f59mqtk+X1ZrfiV0diG/aJMEV8af+3KhNdliYIP71s28VCHzBhwxcrzykyRKnp8
rNcURjWp4VZLLaY2FQZ7bC3XbVTQPRL6E3dc0AH3PC+jLadObfSLASIQJJqelPVmhC1vbpYop9sC
rtqaoJX295wP3nvtXuZzTmqX587hR8HGEkBgyJBVCDfNy+b87DyuBZSiiD77TjuBa3uE7LfNWBXb
65G8u9o53iYysAzYPLdU1vEY53jbTk1jdAvT6YAddmMTEPOJ01d1jXwlAe6NL45EdJfVH/vwE1qu
JNNy31BiPgQGCn3QnUhhzTXtpcnkuDstErwcRQMrCkjxqXTaVdYEApG/XwjZneXjHo3sbbD77VJJ
C5ztfhpWTPV/dO9vOsBVECOCWa1S4ZtsI5CyX2RlyIb016Uw7SMqQrgbENEFlZsXFjdI8H6U2UOV
iRDUSStGxd4cT0A2i9o3P4wgMJ3kEQyoDbTFTI1f+x52CFq+TZUm+X6oW8c+4IjGe1KXn57t+iH2
r5Mqu8OgTKehlXlaNMlFg/C4KtML2Z+/LbWUfBMZCO0qljb7h/gceKi7CBxJvg8wm0sDhhamlHsp
SXxEe8ETN4i2dd4lHLTIwwymNuzqXZypPvM0Eg0SerfkfXQXtnT5D4zLZZMw2GcVT9IWqoZ10VAg
PAhaQmOBqmIHfTKNG+Sa4vgCBgUA1mMMhldeEgsq/+GdJWoNcK0jF36/8n0Tz5N+utHZspKB6wZY
PKxLVssLaBmJYZkoF9WgU2YSne2TsDBYnTJsKgJb+URw+um8vIbz6wg1m54TwYDTJgWV/S5Pjwo9
75T2fgH5WEtFLq1R3Yd+K6vfEo6HLX+jk4XeDiwjc+Kl8+zhjRDJeD5wfYQJdk1JQ4u8P2rdTEQs
iw4NkMLu092DUJQhLxm4S30uEjlxETOCiSpoQihTGWsypLgWIUqeuHFMOiO8EqIsfZyWlXTFnpVF
Cz2MS0f80bO1H+qrhhX9w/MqMsOlekxoqaSypoD522VR+p5S5bgv+DASlYC74kCnOSRQyAPoLSC4
T64cngILImxCzBNlXa9KrWqq05e9Fk5GQX+8m/eQpY5TnkDGewwfzBGcw2vQvM4ob6zs7C8Dc/Qb
3lDaCMyaQcpVVognpN4kuoobPE/XUSweCSEf/qaskQLUhskUmqiCyoy5CWZX3nCEooy+OYd7+EE1
sGRGnAm5Pfqqk0bVVAtSMDygfHjtXyWGcYDu/giK0/S3QMEEMdBbA0cV1Rbin07DbNWnZpIya9lh
RYVGY1A9jTrQOY7CRdpO6tngp9nA48wdbVWKq4fG1W88iNE8t9oVvow//xMUsbqjZ+379VuVRAVC
psPKSzbZjJsFsE3JGhuDFPFmMaDiZzEci0O9XcDrk9CKT7OoKeUP7SRqIZ+6GIJonWDimUCsNVWy
mB8pXhnVrtkbekmKWOiJ7u4gXDII1AA+uKSgzkgVTAUd4DuaSjh9ozriU3cu5Hek+g3DSknMeW8v
8Arv45Rj3zF4WYmvm7HuoIxNC7rnKr76mfyqq8iHvShMdoA4IIrry7i9fOxwUrkZuq/wh9RQ4T9p
tPiPsZ4saF/CH+b7gSU/NmaEL8xyljZOO2Q/2nkotTFLcIc+3z0Y1jfRI0OuJaFYS2eUW5BIvIFF
3ZvsF91THkJ65NhALS0C6A2LOmbhVWyS92OEh9iQTIvbEhT4mkPx34UMYMgJlRoFSwKIoI4YjAbT
+e4aOphYDByFP+SbVfk55IENjEoO0VuElWAXiNy8H5oqjq/9efWhjJkgBX8sxh2BiZ45MCgulpE2
HLL31/GbKg94/tArxZdlsSHI6SKzGur6872zEagfqZAb9JS/p2SJckLRbI31GaQhUDVWm7waudrj
p4JEmL28YWpV6I4QbbeN+jvXNEVDvwa9I9BQTUD0ghxtaYBBjUCILG5R2MtJpo2SUX93ohFxtAiG
wjN2JM6c+ttS8kq8ke6wavtIZ5tqgCbzIrRYuD/Vtt92IeNuIOFkAsGhUrWJpEJYZtk+ubt08hDo
2NXAydqTGtlKHIy+mDF6qndj3Q6TjeTu8YmnX4tG3Y0oOb6xLI53Is5yf8cqIiyMh+kjd9CsEchB
42FyCwnlo0ImdAXqnmVilRxr45x6VcE9sns3O/lI3yTCUGApWP9/5AoEHWGeignsNW1rX3T8lNuB
rM0ClgFOqnetv55jrnTCEC6l4sjWifYZVb0+i6cIMk5TqQAXyriwO4c+8Kb/1hdsJvoYzmCCDFDi
2J7JrwIoeW0SZYncRUXA9U++SK3PmkFoX2NwVWjXHkv/aUB2r6kwsbTYOqO0yRkaoKdWBGZGhBEh
iAqLGDlDalg6Eu7DsTlwoeNhHLouxugSIvqjB336VwcPD06EiVll1WOp3PJV+UgF106zFDhNph9c
UzC96UwlQ6ghsFsCp9KS8617xnt0DPU95zwrGF3sET1p0k0UPQHvSErxub3gYc6cg+3LYLoUKt2x
xXt4im9icpGXLb8pJ3TOteoB/8BmDvw2x8vvVdiOSmxVntUBewy4m28j9NMhewBkJrD3azyFkvjU
GIjS6oQF+PWm2LQNpfBVP/2OKKG4hQGpQU69bxXQturpN6l/oG3FIFJN5iJ9u94l/3k77ZT/2H7I
/OA8WsMIk0CU7oVpBAQOPx5c79eOCBqynTfve6lLLIM/Ral2s/o72TVKvQX5rMN3CsB01CPy+HdW
4S0kVwdqviWuwhU7IbW4mDIRARiLifMxcywRvXSlt4C9jzsbgYx+aMJ5tFflmKTfDTgaKpwIPttJ
e2MKgFdIC4qCOZaSBMC0svFw+QXUdnIXctrdxfUHIcY5flZlsGye/HWeNQHQIBtZ5qVT1FTBXvmt
UyKaYVUATLM3+HicB/SAwDnlCVUWTdt3betQTpY0YCeFa9/L6EZXtiaCjdIj4sQWaWaHVao55Bpp
hEEzWx6xJwHarGcuEW5nUuI4HRKKy92SGhiExm4t7sb/Q7TcQiIQnpFI3Wzt+Fe6R8wY7R/pSkcd
y5BBhvT9vcWpM5/hpiD1RpEW2aV+Zr76Kg4WquhvWjgr/+wZF/EqEbO94hoNUyUIKDsQ27+9kB/6
zwoPK0G1WsZTDKFHynUzm/PuYpbMv6zN1LHnl+ETPdFNmmhMmeEK7zDz2dn3+aBkwrcT53k7f2e+
U4uC5qEkTzbcIV0NZ8Ui/491OFhGKwaosGMUwc6AAzzqinS8uoYfRhvgEpU8TF4LotdbTDvOW7fp
ngrruasLBun02gGmsoNGtoK6nB/kvZJ6XYICfCLAo0JNHgkHOGYFO7fMUtwAw9nKFChq+JknO/9Q
lWZVtkWix9VutkaUCpd98+/mMleNvQKUfEuU40wJH1PTv3K1GwMROsdQeuo1EsNWTaR/JSzVa4em
9/AP1kD7AXHXMWxi/sErE2VUs8yvNtDHJieYnETmrVD5mCx71yQ7yaR7wz1f6xN5uqSvry93Rwed
bLx3/mdFGbfneyR/KbJY48k9C7ZB4WIeGrn6MRzf3lshhF13IAi1W1h4ndur/8C13NMRjRZjqZEv
k3LKWt/q012tVgq6LjpicpHB68K22A3lvApsqq4TizWGPzKvGaPqTOndwcGnCJvKu4DH/QNPfv3u
EJuuT61gCzdLigLWKZAdXLtjC3Q0cTkVv6A/BVVxVuLYvnGcLbdTl4kbnXZOEx2vQQ8TbXX/NlnS
gNGs4DY2zkb793Gz1Kn3A7KR8BWDShitqVGP2jlm50EbJPOipi4jRbpRpnTF56NLBkG1ftN3xGQ1
XxdEUC4ygZW9Wg2jgT+8ZD5Uh9wclep3XxQo0P2WqWcwscP0QdqRpzTw9H6PMzfUOb/okE4jpU+g
s7cH0zZ4s1LgcH0LCvJq/hWjEnC6Yye9Gz3soLkUNXjzFaKL7kZHVQbXCatazpREpX9fs9cVghum
I7xKQSKt4Ksn0VX/GXIeYYTN1n7FeW8k2t7YGIUVAYoi5Rhkaaf8cKYwFJ+0HpVVkFoBDRWcN4ZF
8uVCx6VO2GpZKOTLgughQ0zojYPzExXVKidpOnjRCEA9LSyuV0u+v/gedXfDiperkOxRrOqPpceZ
b+SM56tKHpPxMV25d48LYl6rKcZ0AhJdQczOmNdB37afLW52fjby6hxkMiiJaXY5hhNGqmkHAJ2J
XTphu8PTacfizjJwiqTYgOwVvU/WwWOHTXdTF+7O6xN2pPHN7TyNwoMMH6BfeIfweDeRlvH6uZoS
LynmrzbIQcXSFJMYm2Cmg3Xy7ZBHl+acDpFsly8Bu/kDEoVCZlhNbmCVv8LJrI25IX6n5IBlMhSH
xQBUeASQd+KbPDesvb3FPNOkvxmAtZOWa1uPVf1z9n9N+1p7iM3egZFmJcT1ZCVpqArylS+xDjoe
DAMa3zKNcu1HBBqlAvFdinJF4JsQ4EYgpt4MDyidWAflsrAwSjnh8OwroC6yFKT7gUTKm5BdHzfM
unQvV6f5XOvyR52100Sp8s7Ku6Vlwjkt+elbynr2K7UVoPtUqCEDZyvaQ6SuTO1KxH2XieNFVbuP
ommmJSVoZMi3C3TvO7rVW4vSCMR2sZ54iC0ewS63MLyFX1MRlN10yw15ufM+dq9uCZDGVCHmzcF0
9OQIMoJcwA0tTzcLfjwbQ+W+5L3A/c8VbbEfj4ohQPDsxtyyZoLf2Wg6wenX4SE4XdeDRAnI7jGD
HDRizYovmf2U5oDMQcUOfC8lfBcLiL24gg1JpXit5k+/xBp8SWxPEJDIitp+wutMEODh2kJrgYB5
oyfqQFyTterPB+WtPqVTdcJuqgO+S5IoB3bbKu2Sf79TWdoLqPxB4kEfwSgZvQdPgsqWlpXBra3+
xkbXVfwzKWmQBN7aRntgyaw6LYdzehS1FUTka6lnQ5QgItWQWQ7PfwrC0ssfUPenlKQe7niuFtLc
oWOZJSajCSzYXxe1L57xyWguzoNKi2DDeMnluyjpBf/EqdxRvw9kSUm9ZxPEnJxysh9hJm8qAtko
e2if5a4hnaGCYFZOCGoijCRl4GVcliBQDvJkDFgSFGeOLJyCjzsk7moYkgB+/NvEYcS/f8s301cP
moLHseYySzbok/2/yFXBKE7aPf7frms9oYdjWeZ/oKbk4WU7tcuPqUIq3u6pWp8ieJexT9z37GQr
TQ8Zm5fLngo1xXj46ZwrzonMzZ1KtEVthzmtWZ2xQB1DQvkw7bwCnr9I45DePlHjfAP3azLYfc1Y
EDLXD584x582XB2HS5wWqn0+7wXw1+zKxkBRiYAdBf1oDiyy1Q1oSZFUECWUJkmcUCn8Z9afqVJp
6+6V8ESCKuQxKai30Pk6h98YjIICsEyJsB1p+57yRpL8QYxN3ZJ9pNMf9RRta6ItEco2gJZXsdo3
HZNTMIjbw2AzOE4veQzKBFwqy8kSK6U53LidBovhlfQLJslgPp5dFCh5itL/JiAsgkbiitbQjxdb
ZG8NZswmKr64CJme8xMZfMQ5AlXxd8f0+cWNTrH1eM1p9fMG1T7IDEUASTZEI1uhDvrxo82Yt4J0
WS5mzPPcZV4Fr+nHA6xnokhN3ztf0CnIc32jZn0xu3PxaD45BwouHmyang1PDN5AYz0FoAWd1xqw
Dt2LhSywDEZTX00iW3bcBqCS+Q9VxDGCU3LpOWHmifXwt4IVXosuEFHqa2SQ6Z0j01u74E4D6Z+t
WCe//st6eSIOsog4IMW4Y1IQP4tULMCF2C/NipWjTwft6l1xsjVMaBPXEIVJsmgqsLzhamJX4w9o
hPi62yVhIf79pQb66iujBqOqJbjyrHZKRXO9ueO45XNISgdMDrWIHKhpKKNPF+5vap6+EYC8QfQb
aVymygTbU2+faoy0Bfv0JvSZOC8vMly2B7URxUKKxnDylA/oz5uPGuvCvUWnhF31b1uF+NiqFcHf
SeZ+ayd1x8HHrIXqssxAF2IcjRY7yEXUiqig4MGfBtx1k0GjDKtIvMQyLh0LYE4piYALEkZUU7lQ
Z0YKljkRxChwqDRgzG0GOOln+xzBfeCMYc/r/N2Hw8w2uiVkAIH0TqqI27hi0xskP6BuZ3WPcooE
j+KeYyaN3vAhE0RZ9DZK+ib66fmz9birpxPGuX0hlBsHFBAVLi1TxBDfxlD4A0vrYDbJe7a6xrHC
amA95uVNhWxEX0dEKX9/7RaIV0Kh4oyGsonQx0x5QYaWLxKik1dD49revEw5oznZzw0x0Rz0vNvV
W1WA3RdeCWl6D8HOkXAqgJJxmcwH3ybpRTKSuSBT+LDcVUERNATQNuniKJSJ52BAVJGmW14gsWOs
tqK2yXgbKZYqJ0gI8kon90aGvomEj8HH+sYiTyVvbu75+VBv5Sq3OvCcNzneQnGnJjeR+YYKHWpg
LeJcxClMnx8P3SzahDYgdidJo6ZVK6PTjU/x9q+nA8G++/s32V6plTbNWUolyGJ4sZFzFFS+mIrx
IuAZk5b73cGNDmJNsaOTvV9SZtcKjxHMswbzExCK9n4Pk0Ee6w/APY3+AcZjBoyL84q/zQcksGzl
CDXBaCpitNaPXQYMREdatJJ5dTMSMZghxxt0mIXXG2LDjKFmP/eNgLQbyt7p/OdKhd8jh6D2xTd+
/TuO0oOCUKkG2L+ATln6PH/Z+pS7HnD5kyR7eOdeh/DI+JrBO7jGLHlFSsjhdLWe0lqurLE+f3ar
PERsvkxYlk4IeF0B/tc/0UH+Wvgmvu+bWa9GjnajwYyKWR9szWpsvQU+qKlj+0d65zMqnm6QuvnH
dW1UEdDAsBfbkGq/kAsl/ywD9db88si5fMGEKnAwQT62BciA4+obI1pg9UgUEiHoc/lq+eBwjM+Y
NypIyIao7r0F0bKnoAwzfaWrtKsS2m+DTBu+7yfF3W/zYK/8Wh+NmWEXmmGWoEfl4oGm95vEA4VY
hWV1eHk0I3n0E+fmgnSL63mtWgRK4P5rLYqQX7FqG410fZPH7Oc6SIAexVhqiv3uSLHpoW0uvRN8
4FnVqYg15aT4ERDlkS8W2ElsLXC0QjXvoibJSmtHMTugsmukxdM4DH9IuKD0h1i7LtLhcErgY+8a
zj4ouqmddA0KIzxokPNsWNKrqajOEZWie5keJwJyniIwGfWhdrecjjvJ616Y2kET5CaqyPCFE7xX
jWtby6XSMnMwZ3xlw+XJJsitmxxD8Ok6fPoRy59/UOH+NAOf2E9XZXr1AzFY/QYzQH1g2BXHVjvp
3oOsO6YQTlanxOyd1YwWYWprUD6rHY/MuKdCMsXbuZLxmBT3u3o6r8VjpoaUlKEaVloJWkhd9cfK
5jksmrST4nkwF6O9mI3E4Sq55txfM33Xt6F9wrxaRAtX7v8Gscv8YKFP3BUOfoW3pyq6nuEoSyCn
5IL8UD5rbTXRLQS9hmjAqV4wYyRUi/zsXHd2YbRqVwloPNLlJHR5xoKCovOL5k3o8khK8LwOsiBs
VA2IJp4abHxCYADvL6fx+4JlBHYlGMnxLRbMXtDadRxDFyJu11TpUebcYE0plbbxKl0vBPirww59
UWxw5s7737DwZrlzp8BBO2EA37PSRptoJvUHKuH8VzEECqFw/gd+GVakHqiTcKWBI1ZvRT4P//3R
tI3AAbrUyp+SWCxOXfyDIBWgtagqZG1Z1bfP7y0ksKO+pWWP4eZPcps8jP+OCvW9T+SfjQJjlkF9
IWNo/SBrtvcjGJnml0+cpLHIUMH4HOAGMHBZjxg/BDm0wboep1nWc8jDpWWJWZgrDp3oH1MVkeYB
eRZ/SWqbgnkWZy5+RMx7SlBj6wtmFvidCRb7IHCAzDaCq2eq6mDyHpLDlFIcrfbzTx6DxKQ5ZsWu
FOVmyGI4FQkJu8cW5qEolbH6aLStkpVsj/C+Yfth1rYlYdr6r/nbKzCJlBx97+EOjdFFIXYXUhTC
G9Ox88RXo2SOpoDLIHLs/abrR9pvqDL3dZXY9JLAqgOnVOHC02f2/9sFE/uu6SJiL4ZJGH2kSpAf
nEdgWrBlbzdTDwkTWaUFfZDPGjovwHb/07KOLVrFMM6MhFFrRH9WV7/n+In+PQ3O2V3kjGfkX1ZH
i15R+bALSd8BnJaesZ8qDKABEXLZIVBaKIwUO7e+ZH5NemqsIFwloG2uiI9QMM9k0YFkWuSZyUJq
T57CXK7qLhfuXSUirGbbHp6Wc0nUZrB0OOdVElHvY1pW3NXydn4SwbNiKua/1cAx/3tJ2Ijbmw0a
s2RlHVNhmZpLjSAmJVQQUcKnBkbgpsVfPu2N95SLg4m3y3hQ3RWKLJ7wmXId4oRE6N1uckpRFFAV
vTrID8YfO2M5ywUotEiTGsPAkDdxZDvJ0Yhh8pLC1LK92My9KFDyxsvyxJERWGZnFor+pEnspGgg
KZBi77/p9hWPD61WeMxM0p4Nu0D1QtdU99t/HWteDs+pUFuSO3OHUbQ2jwt1Z8FN6hICBz/SGRs+
8qksPM1yCtGfNa6RsfpZNYgzWG1f4g9FXS8dPtPPnJN5eiW6w7JVJHDi3eqkUXLSkrzRNyAy2jwU
+jbgU4YDT+hMhSZmiZbHxyXCKQcF7U2Wh2yPd1V5i90Pp4enI8NCOx6ZOYXLz60/OJbtUQSBHouS
tH+9endhJB3TWys5ZnnS36tM+rdSAPPkRH8nlkC8R8iCuFUuwGTTAlQIIG5rm9RhOmRCOKMQFHWc
5yIVgjTdZv9Z9ne51u71GjwSQ3EqFt4foyxipdU/46JEtXDDJpCkYxnwQHxQloZP/QW8wV6Z0xyP
d4xR0eAUuWaFdltTAOCS+qZx69giU0zafNie40GoxehiGjpwPjzr23//0IppunMwu9wvUmStv9+y
WbnVbiOeOD9nCvvBp9u3OIbUXoD7/+GIXrzJMpks5ycWTq16/1DBKRoWPm3OVeEiGLPCKaYoMbyY
twLC7lWCSHql8Wd7dynkkV2q+r6/LlEsggq5EIPctHWpITkG8wdGmwgcob4/1i7TViKtujf52Xtj
H2flTAtBabtXhNxLptPh0uz/BwuLWnltbwDU9NXJlWXtyjKiurhmsGg7cjp2Juv3Bg+PM6MQolrz
zHTb44w15vMiueG0U+c9tNS6IfrNqn+qI5iej3NX9W8J9IcRT6acF8Y53fo5DId6cDvA61OkovUd
dGeW1Tb+h2Hym/8Fi72erQpxhaqZJ6PRXeS/LTejmQBe2o5HiIWfJK7eVr3JC/hI5pkZNvX4NWk9
i+/lFNGGRiMw+vfsNswQ6eo10bSvz2HcY9nUX5cG2190xczYqjR6K8u0z+UfZE41sWRantzxG8mG
OTqykbFH30WpLpyF0sYcb3pVuJNWqxr2sdr9DG4zNqiJD0MVf8gdk/paJ9kjt+MbpV1DlqdpNSUJ
PQ6tsAccyUX2NkCwTwSFtqIlEDpFrd6d+xgRSVXG6ATR7Mivby6z+Qa/ygYuBvrF3KuVgIX2O/Xe
NrmIpz21FM3RZ50d8oY2ewM5ZfCRMaFlvw9qjLadeMDLHJAMkJmNxd3bPtHYdqYdoCckFqF8ZXmp
q6xBW6kJlM10LDgTsolap4Tq/8m4fTEcZAiDpumkFup4u591S1azwl6QM+AX27xMoN2hFn9gbUiQ
GvaEsRczw38nddyVBHnu10wXVronSUEQo0qTqndpMW7jxVR1hNiiSw4LApzzmbg1G/m79/sIx10+
P5WZiIAP3F7hgqQJQ4SZBkolRlQ3PT4Ak62Zx0XxrJ4UrS7H/qUsToSZ5eZohNMj0V14AlGN9exD
dAI3I2TV3SItE7XtfdLBxDVE9cyeYF+PjD0GAK3212Gw7u+8C+yEE5EMumd6l4PQ865xiSC2TIjN
k71RaMtTdDgFd9iJWviPlS7kcUguus3IEJBn/vyb+vaGRDB62YBEPzmTHyV5l2WzzVRthzP+cIDv
Xm/IsBhrpmQP9bmOCj06dQabr1gVOS2VK7GldmRI25WrlaXbc5U7eX1TV0PJIIMl9SgPjY0B2ALg
OcqborAZhHpbk6yl9guHhQ5suso5/luKnxrIhaRHjFIZmaXvj7RhoM+QzE3H+0wyIp7Yhaat0PcW
AAzaWBvQvzMtEVuE6A81rLMshFpROnUTaac5mllX5sJVYv3HkUMuXUzlPuh4LHXaT8tXNvXWUNeV
no5UErl/47S4uv3b0chbOLK97j2ekntW/u9TpG6r3d3JHgz9Z2AQKP2QhZDvcf39LZ7NlfJMA3vy
Xq1C8TfcCC4RlIIiywNWRuRkmCuy5tTXcy83ozUqOx1gXfj+h82PjreCI3hm2i+RlEVXXjYcJnD3
qEuq2Y0405YL9n5m3c2iTqavDXMZY8mvsIcLimFOYntU1KIhruJySormOOoC2wSpAc4jhCW6ta7i
IC9JGuOiM7nKOCyVcy3/YPmq9C/kO4QLKgLF8Khs43z9nyqitByjoiBRwYodws0XgGae/T1sfOe0
/shShr4+/AwLiOcSLVIx6kyi8ObCkMniwUCDbVhv/T7xxoOdYbv0M1gZBLRQwJqgqlIfQL01bKly
0BOU1+055dgguCHXbMvfWNGhfTyodHSZg04mVVSWNAio9aI4vBrPshRP6AMTAQ7zgpeZt0BpR0uH
TcWmzppdXYDk4pT9hu6FFeSIIycsPVykFud3Ckm2qeDXjaX/76hoPmJe64vCq23CBTUYLUUK7uV0
aV7JV69VKZ+7OHAHGB71PTGnTEY0xXuiIrGvOfQ9xoiY/T8p5dxqj/kMy81Cq4tozLEMq1OdwuSE
Is30uMSurxKk7R4mW1N5K/+3WRUkq0tUTHbOO0zS9COa9AZttavLPQjCqATfrKa5sG7dMiKBIade
R8Ch0y22lUwd8HXsED+SOkoO3kkIL22XMMmkpctqmD6Jces1I9HS5hCCLh1ZLZLK7GZOpx/k/114
QP5hf9Ue3352kI9Jm4d3WN11Lk4olJDr9BFMfgXm/XLshVCIKBcDvUHPI0oR+Yi0zSUbaqvD8ZBA
dbp5tgHaiUEGi5qCtWCgLQLhAFEUdzsykOEduWHfKepfofeJf4Acyx2qvgS9vTYl27fYICkfaOvl
a7nQOlZSUwuQJvcfGi+mNbdhBAPq8w9CKrnrOr5fD+bk0mUAsRGqEi8RCfvja/DoK69S4t5YuPeO
fFDPORuhcmLVhoeYKqgtpFLlfKcCUukg+uA6NiPjK+60M0VGycL7KZNcFCilpNxtoYyuFhF8QFaA
6lpYAjQ0VZXdxlZ9ADWkhFPRF0L8Il+U0gJ/p+qzflKZn9sIH3edvd6TxJ4Z065NAz5X3hYGBOSQ
7GEzFUWKgXVyb6FDtMSIOEGyNocxEDFrpRz+NRFcEagJlBYpPjuHsV5Z3VLqO+dob63X75+IB0wF
s0HbRzwJ+GEyNaDhO1Yd/s+0+HWlUhiRq1DqIeJaVK8SHsxd4O/ytc4zXjiw0wFpfAYer0te4KxM
6QNyoEEMP94hgiMbdBlLFuKJAOmuz6f1x1c96juJ5m3/MhiFLiYopxKXyLBG1+IAK9hX03WpmtkM
sS7dWBQPJYRY3QLC6sCL7rBcXXZQGE9lYrKxt7mgxjrJpIJdKOPKofB08fUT4y1XgGRVI3CrdErl
YAvy5DYo27gd0vBHicU/sXmkhJN//y0oKE3G0L2HPSkcGwotQyf0xTz5CLhqpomF2K6ck0bGBuS2
J4RxWtuMGrpmRkUL2qOCmliXHn+wbY7XMsWbQu4ZA6ikfKq65swC+AqVK4amybg8kCdU0IqhEeU+
DUPxxxS74ldGfCuguD2C4pjNiJMs3xmGbZUkb5/cZZbm8yONViR5FB3JMe/H68F3+fO42serKMdT
IK3dflxYQcQ7huYg0PrP+fksBU7KL4gtDmfhUgTJRZZhD5VBqWVUcGwe/BzPKcmVYvPrQifRJPOM
qnvwKXZ1qZY++ISJzGdMgwyARzrA5ZHHtRQ2aIpOoi3yRq6f5wO5ucVUniDsFa3sXtDL8n3VLRrw
dbk4H49N/kewIloNaX8FyrtET/5srdAFz/i4mR02BG7wuHpQOqJemAPjyroEXyP2PH13HddOH4f+
1ROoFcDS3ku4ZA1pAuwta8VYHHfxOYoOEmZJxpw0udlE5LlgYXbAoI4hnJ5IXlAcNa1YNSUIE4BL
8ME476HunhA+vU4GiB56N46BoahJW/1GK1AJbp4/p1iGME3uNVJjr4P6Mk6qhn0YiFJxvF1m9kqV
A8VHlUhRGsb8QbLffPD5dAFdSoViJPPnAJMZYDO/VpLbMNCX2CU3t0FBGkW4bTwFt1t7CMLPz9En
M/a248ymGDaF87BkmR67TVSPFak1ywXTlBAsI+xBwxRwprBgHIWJZlr8bI8rRI9Z5sEuQilxV0dO
onk1sqJsvxLt2ry3mh6ySxJLFQbIpJS6WL9XSxWjd4zvPxYAZKMFobjp2oS0iZr1DfihwmgT8k/d
e14C8DMQoE1v2dQ3uOYNmrubEaUfnRGjucZKCcjHFUfEH+9JO8xRgpu0C6mTFusdV8a37UTCozWm
fT9ioDpMch4h0hwD9hd4q8Gl2NHxuR6bcjswD7BLqmsdudGsAHvGDQqLkMH7YAgKCllIm1kpaDf+
HY4nR143ucjnHA5uS61DubCR2naX3UpXPeK3YzK6b5tRmuKUWbHGflYNqrj5ISNe6h0517WJyjWF
iiFomUyJ/QGSKeEHr/gm22F+oVLdvwPw1/rOZcfXJ46vx3PVXrp6kTH2Q1aBrqXwBsNNH6s1+40Z
SF0Z15DWIu5q9Sssv3n5JxpnDNFxtP3vRIYIAJRAiR7+miL77DpSPBXYGpwf+7NQ8wDlkm9qkT8z
FxKVMGtsJdGf1I9oQ6gGJGoPMIRWtca26lMY5MxPl68RPmNjUidDmMzb3NIZkC5uw4yVmfotGUol
emyzhu/NsoNUBsZZgJrJMBo/lFGPNrbJfijfJ1AKAXz/2PZyf+hOtEVbQDnfVgIHNDBUwmaX7uGe
HhAG9GKcdRr+ttb2tywO6aJjGGzoNlrGFnVWX7pOVw6CJCU9kNcCicJ4yJyGqagjZOPBLXdX/0fO
YJSu/i8CBG1dkhlQez0TJvVAmzMQa1brK0/KEpsukwzoS8MUIiGZ3E21QP+F0kIRMQvr+nVbhDjY
/Y3kgoefJuwLjCfV6ubWNF2mA2TRu7rzE+9I0e0OMtoorauzFwTPDQiVnZzw9V1lEQ0QHUiqbfPi
RBo5v9L8lAfwFgaKmftKlDwDFTsYDhDRbj/UH/1TA6nDNXDhOlA/48X/E5rsXLhvK8Eqzjf+XDFr
0EEgnbu959D81TG5nFZsOdyzw5VHglMn9ExeVPkmBBUmFOR1FaCCH+JGmED3H9oZeVIZkPJkJRJx
p80+4Mjd+8Qlgd+1m35Wi7+4ppsxCu+ct1oOWQZdZdsJh5reqB5x6qyxZNN/N7pewpmIvEIHjCBX
g2SXb5Fbt1qjaTv8drXnuZb/+c+STd+1UWmZvLlXeClOR+50vBr2uYfqZigj/6OvwBYOQuvmfQgS
NeUyvruSDUwBm1pTG13RLQZiULJWhOh091EDzgbs2i1qH9GVSwF84IeysH1haUXjAeCuQu72L8Q+
uSgEj5AjBVja15TaaTaWFi8lkm3QXIaM2d/pcxI5WENlDtDrKgs1DbGz9MX6fgSmyJKwCQvTYk0Z
5D6/JckwSYsIRa4iVjNkClJjBaHhfRYG7B3t4I26C+uRIGI5Df7kmavKsBYTul4YdDuCKyXAZi9F
6VYTn8SczmNyUno3xrOuUVpV8Y/VJkGfSnJ+CpykitPz/yBNwY9Hyy9413CMNq1gNH/kqPDDRv4U
lumTlms8ecMZszOBYzyWh36iJxcD/LDWX07HPsPx+eu0PmcKgpirGCQixzqiEfw8J0euCJ0A5ZMU
oCQxycJ+Tc+OFFP9NK++nwtjizpGDNVEhZThPDgVduwx6OmUv2nd1SYaMcxSo1gyX11OjsqNmfoe
nzChHGyCnOlvOGKyu9/1m8In9kKCfUEh+BoqjbEVm/CMyQImcZshAWEe38d2btK51UCzlyFUTpUA
exgAjoHbkM22Vxua28MpfL3HY7QBPgQ35qk8SzMmfemCxB/n8+zvCnvnYbaIaPZ1WMWPOMUJmOCB
YqxFed2m2qXBaQ1pOHG5NLzoYAvO2mjBLhR2/UYX5LlURFLJ+RXXBqOYpZR0OTGWxvVjHhJ67BIV
BzI//9pbxgH6HZQAFW2xAV+AynP+fjLMCC+lPzP4iDe40J1G88o7HhpyeT0JbjGFfBnFjBFhNZ53
lRJid40zQa3/jIlA3UoVcaU0jpNhlEOpuzCIIg+fdZzzQ9BE5vRXZgv5O0pzp9nSfU7QAoZ6wOYy
Ztb3ftIw8NmxkXB7/nZFDSAVAMBw1ZwPskPziuduKnE6t7wag3UbT/H7IoAqpMrbf6Mdc/GaNQSp
sHsAPJvkb/R8oo37IAVosHlu4BOLIW3PdW1zRIprpQeb3b/wJw9+rzx7GS/dxIRvg0V/1Ohfnuw1
ZUbm5qgYsFskSbIP5Z1aPeRcV8kXutb+KlXOVS/VdIoDAWDcJDSRouTGUsubGPr+m6eJ2qv4aH7q
QFakjPe1wIEDv5zDaM3bd0rSQssL+PdB3+VW/G3l9s6ZHr0YHfWUzYZr40gu5Q+DTEq5pr3lexr6
OTcIeWqXIWnqnMglsclh9AFTWEErH7T26dSWQF1oauERzS4EURebdpXHxhP6p+5vM/vZl4gdJ4Zm
ig5PW0W+/X82+dbfRivqXLeRtyaBL5bcO89zqgsVXce8pArg1mtu0dUQllt2FCcIcDm6OjQS3Jmy
al48rQMFzh3m/P6JwK4ursbfFUh62EWeiCkwHoJd7jOmZq1F6ujpKGt9aU0HOW+5ebB8DHWqIXbs
plXH1r6/hgVVV7dN3DTARJ7XE5CyGqrgUaC1ZhgcBSa/JKDs/AdEBnG9U6C7JSCRd7NkWZXmjQi9
tGVoQgjBParDaGWyPIbns/cBRfz22SWzL6E2Vg95n933Av0rrSv+pQ2btfBvmKIWvsPSuhAeCuWZ
cGWbAO/+yBtzZBeAQeKHZjcNFT9Zm14A/6djSkzML1SfdT2qZj70seY1FypXS2plypAFC58xHTh+
z3fBy5QET/P9ntPeUhf9pms2E9kojnD09G4xS+rW1kddf6IkL/WozJO8bwKSKM3pgoy9S3Kx6C4i
S987q04wUF2djZq4T217NFj0XKYSzcovonPYgb/wDqrQk9sAaN+W2pTzgbkMwrEZXx6jMnOFUTQM
l+2Zdhbm5t+Gizl0Ze1KMG6EMkGAAa7I4GsKS2/k0x1jKPZB9bebNvuHQG3Q/m3i4zvj7889/rAP
y2i4v5StwtznoZb/cNToJoLB7e39+O5SmzTJ7uz6pNH4yILpk7cs47J9xpy1Ea3U3eAJj8fIOjmj
F0zZTLqKKi/MgsXqLAE8+jd+gxg9rPmqUlFm49F291uT4FsJbwnUKaQAkJb4vFaBCprW00KKBbRx
EMQobEr64CzA0ZqNdO/2dxAKqge612irFkEkf3XFrFamaay1zzF6P9MpbvbnGsC+FvdRhTkOxMrH
DBV26B1WjzjOIqb8DaIdZwbh7RL3UG9sv3PRKKDDgtvBzV4BPlcKfidaR3Hs/pVeGO16ifQYXa6c
JYuj38jWOGYfcHF2LMvQqfMApdAWzZeldvO/nVSuxILbMAntXcRKZHn2GOh3LudZRRZscYklh8tj
FeyvjtmmKlkp+0wkorYSdwmFXKLky3QjlaQGJTYDK1/xp7dQAp6dH1tJ1TTv/wj5r7+RTdhV/TkK
uiLNsWqaJ78a3u+Oda1TrjhtRC+25pI6RfabcGDa84I3aKgUecVis94d/FXH0PrXrKa4atB4y4+K
c0PSkVf7tqTQZW3jTCeW/j6KwoPjdLS70EKWu0QeH6rj717ihwuCR1asr4Z59Epd7RhC4nnOr98+
jce+byPw6SLSYfQ8Ak9Ghet1rjFFytBPHWrVwdydpRAQuoFgU0qjtJYXjn9b4k2k8piK6nvBjNt9
p2D5qn2VZTRK00v97YTPWTwJsxiKq8H9qIKwjf8dIg8NOpEU5N8Yg+n2unnYUUh2DExafPgf30vm
DV9802bneUBSwsZbRhn0sC2tya5YM/4m/n90LScg6I3fh470dR7Hqu51iFB+/Jz9rhZbAqgS8Jeo
UAQhMXgTsC9I9OGFBzkF9VYUAyxN9meTJCMVP2/MJBOGYUjtXRF10yLzNdfv1HcEjReEj680+U18
yfWkdK+qaeOrrxe0BHly3LhoFTPZST9zMYM9itTWD/vA2F/S7XpSxiLBq9uNsE+GZVOt4fI68BTp
lnXUAE9roZ5yCCMp0U3VqKe9c5vBlnwJZbb1EKGuoGW8Ye/59QpbAknDtYW+t0Xtiavj5+IVwFy+
l93WDMkU17u3yMgieJC5jNcOEsq+sh2G4D/r9dwe+rPPc7vCsPSn0cgLAV2Ed7XQ0rs89HnrqNZL
VuCaGMF414K/HLUkkSwXBFnMVSFi7ZEG37+7oQvUza+dyfrQXn3ru+T6oMTrHzzD00Zl3bvl3pya
8x6Yid/1OjA4gWijWZA30Mq8U1m8l5DXpRR5fhPBVUYts1Q1/0umLoh/6vXfwGqK6wQE03Aoc0RD
hP5yA29iQLPaOPzYtwA054Cx7XBYTwR6U1bgEmz8jF7ZoOgw3nFJtST7FfmccFuvtPy4IJTa7FsP
FOfTMvysg+drD95IhAHMmujO5sdRXBBAUgz/L+nUCsujr8HDMVYbAXkQ/JFRMMwwNQrbYs1XGV4l
O7UainWsuo/InujXWly4HCVDak/qqJrhO1DsXkjuQjxlcHujhAkVy6FzJECe81ZqKcU4BqvfhfcT
djQoFgIJdd8j4SYNhH04o4+UBLpvZyfzqo73yg8pUn97e6ybx2uH+HeKZZuEFQdMss3O9dXHOo/T
JDN/5CxOgrDAo4F/0/+HM/uuGOmlPL1QWl04H19reE097HJqXq1o1tx2E3A0+IjsPbrw7vOO9VP3
6dF2SGZYV65Uq3vJ0sO52q9znDY5igMtCBdRmDVX9yScKf0pMY+s6QCGWXDsNtEWRPOWkCwZxawg
7y67r1301V7t8x/Koka6fJdkTYQ7p1UrMRoIFL2dEK2l+OK1FjdwHbV3+crqwKXvNrzN1/3MO6rE
qRhuoCFA9eXDrKQb+8f8Yh6ppBkrhh6HCPOyWYrqHC5J2PqQKw/3BNAEbJXPxBiLRxWoyHZTtMBa
Ikn+UidqUg40FONGWt4hlzergAMdttVxB2hRdno55B0jJ9m4yOScOJVHauh4Qc/PhfAVvbAXzu4y
ZKFqWY+G/P4bk2R3OHWWcxrfv5zWhkmlDS9tKjM+bPMsbjUoXa3G31OoG9JIFgpP+ptmQkEPQSxf
lMGIKXNqgsdNCXCzH9B691XDvVDtb683MGkkLpxlHHZemp7JAYrwbHFcBRHT+0d7ofDfYsmml8Iw
peiVi+6sva+jqkuHsP+bLVICHmYZIV37ozKjpMZ2raR1GqPtIsaaH49to0L0/GQkzOMhTrHQYUCg
/v0ZQp9abV2E25PqNlrqeiXBDYeHMgx75otsmA1xOIs5j02ui6AghWo3e/niL2lP5PppUAe4u4rH
v6w6mZXkJJTp8FmMRqAbyi4IG0iv1/jjq22GAT9To3BPR9Ran+M7JCOufo9BgdFHAsjOAjm61No5
cTowppDlhrx6eu/PZhqGvLc4RWDi9P+23DfTBsP50JpdsOuv4+3oURh6zJxz/erL3l6Y5Wm3QlWN
ATQnXc14Sb3oCnCFknAaJPyXCK0WH+6FutdY8UwJKKStUPMZCSVulp6HZkAG1I4U8N5X7fwGlOZq
LjlILbZgVwR06MSjHr16JYVrC3dIdjkzz5iMgewWDddJteo5q6NiinzJiqtxGbAKvVX1nFIkJUMd
KQYHjZcNryIu89WHllMkShSYi5I1hUy882838ZUdLbwAxt6Vv9qYwu58lhNy2OLS8qvfsBg/gFAw
mq0WygAN/zoFIU1Jj0AV1EtIerAvsFy2NlqIbcZcOYUEo3iam2cGUXtfWoDfKmU5vzkcpLx10E3Y
CFz0CQM8+58Z5mqMS+Cxwt/dixEEkXnS6RIipCaWi9y4wTzN0DKKMPqbg5nJ+1lIL91ZEH77UpmX
SOBUW8OArHVo/qqr1JLKlwEmXjrdODKRd3riqpM8taihSM9ZLXBber7rmc2iEc1H4GKfNZRVPpWh
eP4ZObTPX2xxIqRSnDdYYOME6OH/JMwIJOwYgrMnCFntgV5fjdvdynZccbOmD05OujHyjo3idBUm
9Q0LDJSdzIWyPcSRvq+nL7TgcrDzLmQLnfqWrNso9JBO5dpnM9P9+wSro1R9Yp8oOeQn3GgYzTqy
DU93vcMvc85xErfjARlvL3j0TYR63tCbxXSR4IR06wej0maUraXdAGXtny6i57EvU+H44+n/vOiT
/WHCIHdsrxB5J4ASkgEFPJXhLsXqfPQIbC0ctmZgJUKRr5p4CU7q1aRMv9UCMU8t2ZRXCt227Fga
A4/GoDy0PiSmH6LjH2bDX00iQqkJxYsU7VMh5n+6N8GVQap4/DNdx4S/Q/Vo2zVNLSKUuFAC6iIa
xVciZY+6nPciWoLnXqQ1TOoBrgBGOC8i9TKXFSJko19OyQcgvAzE//mdOVyIXw5Yo34p84ZCiWfD
aLCszw6rDMuGvwsdAwHUBw0iqLAbMVTcEAqb7r0PsaHazi4aSQ7k7o61PrqpuIPiPAnPoPZrkEBc
IjcXoyKi/4GUFvR0+S8d3nlIzGA6a3CG3GGZ9vd4MKdE970+DgnxZhXzHjzJ5ZVYplpX0tFaMbQK
gu6hibxS2c9uYocssTNrNQZAjLSWl2gVgtJzPe6BepI1SYZfef79kYcP07h9aPXToOqZEdY49XI0
8b+puDmjecwIqPFZjtzJmDymhzewL2xeurWLYyMIObl052TZMKuTrABJVQLaLLXl0Zc8PsJx7Q0W
xB5Zm3t+Hv8N74YCSDMjB3AqTELkZsgGlQuRGGjEbG0gXnedxghh72r7B2Ir9kSRSIVBCE+9iQeN
24XLyu3/gnP5U1YheUPMy6bKiUBHjpNdui9EuemuKnuYta9bDP5/Uc1zVmonz062PZatHI6o1gMd
TglVU2pVa/C1+LB/NI/fD+rU5y7sRXHIGqw+nqfknKHV+JPqyUaoqNwrDYc51+JTg82gexmPD0rf
Ig68TUd0YKWSQa8njqf+LY4P5euBiFP1psI6GrPqdHutDLPZB9gT3mB6+vffveGFRFpPzTpSHa02
Xn2JwzwtwkctEeWMYA7J5sMtwsYVTc+q2MZm7aMU4SVW2HZTJwn4EYrOF2RNcxf3QIFSf4bTVWcd
N6mzBbzs2P4JBy3qodS2UT5U6aRq6reIJigEockWW2rMqRSm3qDfC5u1j0ZqLNLsd3CDrG3izCL/
/EcgxwDInQCQV/pmXR344rVFTnsmZF0kqxPgfZCiLOvtGOgX8C4FurLfpFP4g6AsSG3Nu5qAGo55
Qp46cTsXcaS3NrABwzaXli5p8gQbOTwVqgIZuugOTY5IClNXR8yUt7i3bUHIVGuCJ7GKyR6e4QXG
dncfkLnQEmik4zoRq4x2bEKFvxOKj4x7COeMRf19cJSXDLhsAAq51lDMN+eUra6Lmk64A3KICUfp
TkQTVurZPZwGNWdYUE3p2GdPz0eaPwrrYJ40yQ8uk0AQBNanSlLuYX8GefUecs2nttcIIlpJdysL
aHvPMh+TOKYJ0Tkq8kbCa7niEaNhs01qXMipLjxF2delZw1Dc05Sy21BFis2lQcaf5oWeuYecPpR
Os++8U8O7HdwT8yCKSgOcUM4nYVXD58MUVrQ0ogbSor67z3HZ3YCZUa4bTP6RyMZ1V3oWj42xv9/
mLiMABjOBYYeLqm+ylWG7yiT0mQLRimYb0HzMVllkLei1DS1vUFV2trVAW2RTvCe4LR6oKq3sYvy
4hG8wAarBHhIfPug6hdqsk6dm4cEn5JGb+mv6HpyhubJu3+4pkmpGvtiyntcchk3gZ8kVHr6y2QS
f/f1lkhXuMaFX97QC4s4z0+g7y0oc70DtOG866fWTEa6zEBjoMPXEphGP/Zfh5SXQ9SaUXRUIdEH
0TsMYjZAsgDtRoDfniwHggKa4FUIbYX+LMg0OswSIoroo1pmoR6G57JPK5vbYJVxwU4rSsHBCnRp
owop9TJMDnzibsmnju976tiu4fQ12hDYO4atK8uHF91+XmMIFl5ZGX7QZmgkRgmP5niMu/ifpXC/
Ajae7X8NZhrqEL7k7fybYhfE1XKU4IUAGXcJVa5+v3b2U0OdTUl8HWI5sXcqPjvZvWWm1zh8d8fl
6xq7aXlaKKQrz45kDhl0LlaPbwP0veOQzfBwa0fuo9d/IUqhA9yH1/+KbStciRI+nTunlWteBx52
/sAaIoQfMTSqSCHXxgti79297mQ/1GbwmTq0y19orqdpF1cDWtsGveIXwhYdvi7K6J6Pk9/kzcEu
Xs1EV6dkDiqQJeV462uu8QlqgW0xL6VcyEhf7HE2lkgAbkrIjTlkSZzgXCmDou7I3DnpAZrJ5Nuh
0cVsoANFLhntnensF2RgkgGrWHfBqxS7fAWC7lLuhkbGVCMNMzsPUvHpmh0b9Rl++kAaKNTOKJOh
wxoWdvgBAccmi93PXz5RrGBoFJH2UUoTuk7cQkkNKGh38/4bMaU4kGE/pl57qhOTCwx2+EDP5jrJ
Qn5RLb7mDAKoups9olTc3ORuTJNr6FQgIgLvUP+CVZk9fWPuglUgWCaEwapKEg7dYENZBuQtIvuC
NzoATbIkSajgginbhfy/fRbbWKjX547HYP1kCC7tWCZyHOQUxZ6PFUjHZmIDVyZOU6nQvbfQ0uyP
w4yRaf0836RAHJzRulK6N0UMI9u/HmfWs21Q4A0tB+DbV81LH6BzgYeWrPNHH0Xm85XwWg6oHalV
WcxAJ3xgpB5Zl7pwN4ukAQYDqFlcK4PN9TLIsb1/jnmXU7RbGKutedRdXC+OmiCEVwy7CehU0zAo
5DtEkGiornL7hOLNrFNoj4SNmdqR+owecDgLhIQ8+cZXgAqZHxxb9p9LHgVGk6KLQz/am73a5dOQ
woCcUQdSZ8isiBtCfUfACBZ/uOfds6HqOjMzl8x5X89H3diAmwZ6V2OOqOGtqr+QTjPXbh31pP9U
w4Xcp1fZ5u+2xAvBFKkN2qrJXF4wvJ4f4m9nZlWjVfJeiCfNtyXpH48Xdh20tINjzVZFlnD420ll
vo0N7mpGM9m2S/YDR+wf9JtLNHhO3tgSmzGWlhEomfx6aD4FfE5KRWpohDGkzZmIgLJyhz4S3E5b
GyKq2FzMdA7CPCSN3TsSjdeuqLlq1CwErqoED6GjlYtno+yZ1JnoOKLw3maOUWSEJOsV0mARcDTt
Es+9kYu9camRXswv4MhsJZhRRrc2DxvOlLNHil88/lbXPaEqJ8SARDdzgA9ks9Yb+1jzrP3jrkhu
4TZi+6RJvoTHVkMpmalSk8Kx7wC+uuzTyOkEOf3fYsqx5OZrMAaf2b34PC1YqV6A1ABZNNod62hX
lCe2o/GPRr/We7/v4oymZ6xhloMQVEa77TjGOcWnXCc0PrZXqfKGiyxhBJkaiVbqtWdPk+RiqGg0
eZBxlVEAXk9/2+mWsgNupt6ylgkLNI/f8C0TrAR2RcxjteWiZU9RNFU4f9Qzbfa2/pkZBHO4uyLQ
/XWL/NB5EXdZ0qwsuLzxTfrxYdY3pyDC8tW6e8xK2Ku7vqAvYO7goQKPkdipGA/ItNc0saDIHlgh
gYk2MoXMoe1iaxPmrhRR//aFj1k6rrw0nn4LJClB1uhskxfo4rNlfwtO9BHuXiTZG1cH0U3QEEX0
JZ2BWoV8NwiE9/39xNp2ifw59QgeoUTUtPfdMZ16afUDKeS5IBv2XpJDBtwdz/mYfKCPUB0wSdW2
t262BirXy6zYbCMvR3/JG/4SyjsVMw1dCW2IksPMXl2Pm+iHZp6tHosMpSgNgepVranGdh6/Evv7
v9Rr4Su3iQRXzTnv+YeeXxdsIO/txz2C3hgyZAdARkJ6gLmOwqJF/l0rdU9uzF0c/1yu4sWoWiRz
xzYbsL+fSlJQj34ZzT0AYggJA8G0I4qs11BCO+olkRDkodIcI6TA2hVBT5eJfeV0XIMLSVlXpVve
uYyyqBG9bF3Odh845wlmQmSy15o5XzGw6v5fSj/+WHaD8q+0HQe8KhWRgPjM7qt/CAs7cAuFn3nd
M2fGqj/FLnSOs9Qg/iq2XqqR//A1OXUFA4+uUZlHru6L8HCo84r7g9b0pa7U0K5HKq4fyWcq5giO
WizVHhC0O9yU78Pap3c4WvxtNyvYuP6yPOV/EmV0zSOjaP9iKe6Yy5RLzMr53VmXLU0lLwJGSgSx
6Uu75fRbwNE/0wrvi5Cb1XVdBI6RFZsFIvTn492vdwcN/8MM/8AgwIYg/Q5ofVhY8jCcVSm1rcLk
V8FiYGCvLQztVPIVCbAHWsGP9CsNeG9ap2f9HexIr7A7RLSUaYpeAqyyBuUZ0u9zSaSSv7giS+VA
0QweJSmQzBnQ2tNFo2SZaZE9tce74AeBCMY7xLfwSHhLJeguAa8r+4wNvkIgg1Yg8mhpTLahxDyK
dKsVz5GVA3ivcNStj4sIGe+4mDM+jPZyqlT0MuYpgpHiQEtQrM5rTdIP0fLbm7j/G2akpfN3xpyZ
z5EwVkLs4V/4RKoXm7BDF2EE8U+e91da/IGtRtjONxeZ7u7yCUPP9TsED8jcnrNUW+N28PqLNkTS
uGqMb9blG4NJIbpKKOso8l/HEDJ/qHVG3OazqlHsu/GIXtP2u91p68olqgn4BSn80Yok9eH6Dtu5
yeDFm5N6YgWAzQ/hrl+eimvP2/6g729+k4f4fIRlF+rjSKnesF7KNjJ84KsftvoFhb9bZSi2pRoq
wXHBfUr7oqTH555DSJClTJ6n8VQWBdJIHAM2gyDCiMuJIitv+DSQidtjVqWEfRHMFRpfmxT4Os9b
L1BX6TYttriuhKhHZ6pjZYGThJzpDg1Gpq76jgbCkZjQ3XMDSCbWLB8kixssK7uX4PGoSzAq4tJh
F3ZtgPRizHE1ClIKWqDH5/DSB4+q3OmtBATXG03j+LKarLcscxadxW84FsskK+5LNU8hcvBUNKtg
ogz8+7g7as10PsryKiH2XSmwJ86aSpL9qfPXay3MHzn/pzr0YnRDbhmzQM6TxliyUKYVQ+D1fUui
yjovIFVgFLU1buYQhW5n4Oz1HsBv38OEI8kdPd7eNgyiu/PBitWDNgLTfk8IIoFaOlUGbXauTURe
228R8WUs+5BzhDHhGt+yvLtbjkn9v0Lhqk2gmciAZsY5gkeoSIGTikNYrvLXJespSAbw9GMKtAXr
egs7d/nMUk8sW3b1jynLoYkFM+Azgf7idTfgkYLxEQjEPrgm2AzJnASkIKYg7ymjao8Rg9bpQ8VZ
rT3qLKT3SaTYMifXFYAva+BOTKQuwX8fWuljwQpIc3CwHaRJzlLb1u+oO9EIdg3mAdZe6c1aeFfT
Htr3HFMFGGe+HmMw2kWYWPW5BPnYAmD0Zxe8Ln9Dq0pF0ZYekl1zwQAlJ/ih3/N54fumJYG8jt7Q
0VbGgJMHf9yWF1fwblb2V4auAGXhxtCBIZL5RVY9HUxlAYT/S0FuI25VwjiD2eXZUyUQN3Xrw5YZ
GOTiyvL9UvdpDahsD36WqtDNUtJS9Lj2Dzaxl2XJ1HiCi46GyL9HyUY9k1PaC1LFb3f9qIVYZoE2
k5Yb14+4EuGBXu6OqbDH3HpHlz9N6R6FNMQnSwr0CdFndYunfi2m+rkkfNSQh9iDYaWTBdpPQuNx
MsCKCwbPRRI5Z1GPpsfQVHOhy+/CJLM7OLgNPB/j7wMtBgitqETKZK+OAY182gda+cxxRuv0BkAk
T5iifQc2122fLHhyg46db/rhm8MZx8DUAcBNzfymDBWbmyei3zFQpv4egzLm6PD73mrCAWNFshOg
l+XxoXDfiXATcIM8NmAxfteFUKO+cQosjx89HSkO3n7F373E4Qzefjtnsc58sWwoKclbz2+QbS4e
5ZcnVWvHY34Bgu+nlXqdw2gmMbso2x59AZ/pvGgcWVdAs4108T9NP2EebN4TF8hADlT14psWUlxl
cRDu1waxEIrpZvLAItn4GtB6MqResHlOfbnzn7K0JklW05mt8Hyhs96oz71W66vqm/MCAOjoWiEc
NXCErulIZy+y6Al43WLKZ+ZOz9e2IXntBe/a2KwdlZJ8DyHERmaJn7Afp42dmEXZwbFwX4IuNTYA
z0Tw2/6XmQbZo1jqT7Cmx6EVkhkbb9B8w3WKDe/r4NYxyFaQ+hBU8HOAb3pqAGTW/AdbacnKVFEv
TTO9VtlqrhLwvEb35kChT8/WlKgZGYCweqVYdeBZ5u1U189p5ZTF+4a3PZ8LhJaIVcFGVIVMefUF
hRDMpP0ajYAJVNsJVcN5Vp3ZiHXA6mkSOx1FjM8hbXBYilXQhCEgJCnMl3SeKrxdogXB760daFXm
hdrjTGAr204pey7ml6b6yeC6iabKSfMueqqZ1r5qxyBElm2apXw+SE/HiHDjktCjM9EIj9KnyEs7
LMpO53z28J8Lc5RGtKPD+NmgcOYxBcey0DWNP6fGaY7CSZ775ibdjFRG5auqeNvODFPSB2cxvPdB
FCGHJlJR/mjHdvI1pVQetYC2CYSgwFU54Lcoewn0K4DL3r/C9OiszZJh03lvZ13B0DXqfcJ9A+MU
S7OsGHQL+pV1D6w+JLq02I4XvvBDG5wpEeO5noQNRd06CiU6o8LxKH0j27XTyFs2iJJ/BUmRUMZm
xxwMHf2WlWm6QQjpguRIJGuJVgYbDkuHXBYjxLTYk5FskgVB6W5HI1XFgcbIsbna5GXoBHg8rWMr
HSQ10NXga/bSeRdYwCdFcG5CVN0TlFiMl9qwMmKti8rb6UhxzN3dm+mEOKrtbRATmzxtlmdYLq2f
+Z4JB0JNk/BoBAa5m9i7aRY+i6g8w2cODtkRw7V1Ki8m6zArRQWX5l5bmTb+AWwcoFGI1Ye7qz/5
SqoiMGc79LA3EIrnFdBb7ZvodvCgFYmrUQ3ua6E7f3rE7m4aZ2rV10B/wAD32Lrj8xjsoh1l9rC2
kS9MIJpdLfFeMD0TbxjKVi93oUrZ0dJinZ6s5H3xHZWXFdvu8RuZuTgZYAT0xhswDvICvOL2q4LF
oZNGV9fDOffCz1qJh290c8mxKRn1JJSoI7+sk25WLrl9GTD+crgh4v6TcVTuazbFi6b2k3cfb21Q
bh83p7p2l6bsoi0s/pTtWH1yS1K+HyRD0BiC7wIscctUhJNyHMaLAoXwcDsl0MgtFvXnpUfxMeE1
9AgeQsDXB5d5Qjn/Imnd9nqjSTo5a2i0JC9ofa8E2ydDNf6u2pPi7qYcRbcVZZEL0tgacy5hAUs6
y4Txam2akiZgtXRvXikEDX9K4EEs4wxIEhXg+bwdMHpGBAM8yKOMlxAsicjzDTw/Go2jEI0oFCpn
Tw5Y+dT7g1ujMylG2WLHDQJYTJN4ICevkwQIyeX0Q53xbJ5I0RinyyFH5h8xSbij1GcwqIp+kM+j
N1RYeJDbu6/C9aANWo2bLo4U/4JXpl8uDwNBOqk1xdUFVYvzcASSZhUmq5VyqtaJ/gjgLrPxeiaj
X0mRykt+Kllw3nPRr4C0AflLW5s6wVyQu7ZxEvUiLaeG0z6Wmw4PcNRSYOLxliIheW2zaFU1uvAF
qz0jazybWfJXGNr+Phe7lzR7P754wfrc33O9r1tMY6aG8+89PvP/FwmKtxfej5X6V4MpnrkWwiZA
jqTW8N9ZVGADw1CcfggenCAQ1yETB24rzQhtdb7f5AJ2VpmYW+uDA2NAdk3cyVWk1Pt8/wWp9oJu
gQ5QuXwYiKKav4kB1fpDfv/Jw8EUK9hID6aTpWQuSoQKfXs6/NEre0AuypO41EJ9xsxZEKVu3N14
mxQ1brhWYzMZ68ezh7qZ7G0OgLCc9LF5tBrRZMMKMnQTdtKLshM8q8IvXQDCJgYX2xUJwVk6JPTs
goRiFqyi64XlMTcKV+fOJmukybl/YUJFbdFcU4D0K+ajc5ya5IWnrA68Hgp1ie2F9IfV0TZsUA3v
1I2tfe/uDmS/x9Bpz/HwENRM1YKgu2RXmCzOdhj+Vt90oUdtwjzB+GHJZ6MMbKMflRZW3QmTFIS8
p4dICbsmI+NH1NyJ6fyyjzF3UfD04YIb7733KWZZrdoQBWkiIH4k9Gn3XXp1K6++mtKCurhO6/4I
e1CieWTHYYly3A0w5m63rREaK8jn9wAHmtvKTJBTUEWsCXDCOlSB7Odn9KlAzrzLq3b2pXfySFUi
0bVaw7aBi9bFK3am65f2wcBw8MD+8wAEZezmtJtmEv2Z2dnaBcUy/d6F/vXElabueAjntCjfvAP+
Wi1lajs7gv0foBXHYUaH8819v9lPaL6F3TedN22VDPdT6zyg9v7lkilFAFhx38d3lyzhC2HFfx1+
6309xSf8fjeHU5erwne6CEuEI20Mzvn/SshlikYfIB1ydFRrwLU+j3NVpSFACrV7R2dhh3fZH0RE
525FEn2ueeP7l/Tqpx9j8C5W/cmm5sLBbVSWHEG3BPS9XmrFz3O5PaCJfm5WR5j3RZJh2rw0v3+S
JwSFBXFzGHUI40Huq79IRu/+Y7pFkwoTyRwSj2zWruRXK0Y/cnmwXd9vIwp9QT4I5GyZVS71N6w8
wZwHJCoLrT5fPYF3QVfL8a77j8YAW/8YuHM8E8K5pL2uU0ChQ/pkt1v2w38bKcPSp+YZYmKldl8W
HDRogFkJ6yG8hvMzYfN7jD/myF1+75sj6cX1PTBCYd+U/s1GcQii/RA+iqGCn27/2YSURRgF37oi
JJbHJ9iXD5WX6NuAtRia5SuopQ7XpqmeDoJ6yqJSYqWsetKwlvEg6kA96WtFVu+IN5hJDz2mPfh3
l91jxpqAx1NtAUkhGI70uV5k2cz1G91k6XU7hUb1Q5g/T2xFcAjXuQXlRuHZvhIPWRm2thBHRQLp
H2BXW3hOeE792ASfzjL7cRuv7n+c4rJZ+ujNm5P+Nu52oQjbGRWaLLeCAq7ZaIHz4tkMkATZHCTP
VnFE00YSBnIB8peV0IJ+lGIQ6mWie1ONpwBQ/Q6kKJHrFcmHPqADRMfv+7rfRbId2oYvv6ohCeUl
GjHZ7fDNAonHcJJwoHsnTa39L70AqaAU3YGFGWlb0/XmwRnwvlTYptHbUDYq4unz66+5l0Ja/b+W
DJUVBK1THD14Y+iSg5tF05iKD0D6oPZk2pHq9nUY7ROSGmKeSYT3FuWMrvU1IwnpMW8shimBVDQx
bhHbLOvfTaKfR3+3cx9bnkDVJRAgPret4Kbg9uoXzcRkI6F3c9eh+YLZMQbAAbtUBJLCOFAM/c/j
B+jU335Fam5/xQY5bCDuysj+7UoQB7dEllzJSFWuxbWK1Ka2MmMDm+3691HQ4LfA8CH5AeoAkFf3
CsxHheFeRcvigUmfJGzJZF2NU9gAtXkHSBLnWwi+OhOhYUbGbctMdgNF8l1lcKcaPu0qVPZqTdLx
Qw91jYeMvLYNuSYlG5nthLKZ4+HPSVDNhRQYSk5boQT6uePPzO02xWQ3Nq40DyQoiK7PtSNoUoxW
tEfo+iO061fgQXWB/9O3ukHbeNu2PpWgsR66Bc22NEMNryy5gKgJSzBwWG6hNqso5I5XyCS75k4I
sDjcUaraojKBfeaWko/4WbAyOcPqDlr6Nd1RGGUYNh2JNC2KB2dMbO3OPYRDhSDMB96K4yuAyl7Y
Oaje+H8Tb/VBYWA5tOxZ0W0fAbkTPXRXGIiNZXXXC5QHbGGtKKpTlN+qwervH32eyW9yMvkXWpMU
fXyhyOoAxXDn71czijS5QkboOgvQmf/FoJCFOmhXvRKhRJrcZTDuuTkbXBzmaOkNF794lTRdANZF
tNXrnDkNpmC0Q4xAJ3a7BfQ3EipIAlnR/a+g2i+y5T1vZ90PKcmbW2Mp0qw2XqLjN/MGCucrPck6
g1mjI0gtQEODA+DTp0QNnHbN7Xm4xG+Jy6279/kblgzGd/J2yTwEzGuB8ltBWTDjOk2TbzdcDvT7
8bDXw8U5cW/cGsmi57b4pzwM1S8Gc3AghHImB1jjdBXmK/7KtxD84RNzoNM/wjnabIhkvccjsTSD
JopAo5Bg446dIV7NSv8a5eEfWVgF5dK4l/IJP4r3DDALnGNX0n4KaZJZRnEGMzX5UR4Gqg8HNP2Z
9zdZYDCrzr5HApZbsixdXWB/OQQHqpNr2zolRhb5thf/CJhNZ99nw6LD+yqU5b118eEsDZn82aY1
tjuHYNolaB4OaJsV43N7bVF+zGaZ/FCLcMaPsDNPZQFxO/ZEnnXAJMdftqN7OJ6f2xlDuiiulpCu
joxchgudLLE18Cjxs46QOGtHx+7wzMyVXlhylq72pu8Ai/7ZTkHl46FrZz+OKTAgxeRlRydAJ+VQ
UzuxXgpT3tKN3bCBXQ543T8zU3QPV63wiFfpsTGFhBKwoqFwEnbPj+pXd1H88pDkc2EbhjDxVS93
t+8hLBlq1kD0awr9nTJ8HpP9HsEPgdZfpQrmQcGe/XFsXbl6YQAjkXKwcGnVDSFsqkSn9t6LjH13
80F/Fs1b32rmwS26walmZgPtX3EEaEYw7IyGzPlbdvOzRBnjCPGotCabfZKcZIyFfx1jk2t1erjO
HWLh/ucx/kGQ8q1xOAcjf+NpuywGh+d5cwkcKT1/ZuKmX1HnQNCkrGqiKbqt6WCoGzNGjlZ/A89p
T6v3vPCUrCBeJGxumg/pusdlyz/Hu1Gw59rZFOGVTWsYX8KFuxsosSwYtjVJG0QOGeC7jB0A+Kkj
zmO4R4hyA75BilFpUCBNdbAem6BjQ1Z4dd282JHwglfag1ZCT0fTAxwRe7oal2WFmCPgkSqyWK6V
wybX1IN/aK1wKIYqGdL68cWsDzKpPYtQ7CKXNH0xTgy6GyiOZJG0yrV/Kzo2fBcd5QRMA90vc1nq
Y/Qb8uxPbfCBM45uDpjTbEK6vkIEHW57OSIWExfCKuCVHnm+5C8wudcwecxrDRX5X5o3mDl3bGaz
tjYmGIuVBcOTkKKoWbPqpvmWkYOCpzfAE74DNYuxImK1giWfHhUsfkmwuVhUpTuhRRhnbKi4AGZX
l3HU7EOPwbx1/c7AXA1xwv/D2XVbLjplJXWpFaCaTVbnlOV2lORKlF8eTjJlppSA1Z20Pr7M20NZ
x9ZOcAnBV6CCa6MBr7vyGXQtfFVS5iy4vz1zS38iZ5l75QKaXhCaEHn996NV3lXFChk/wLWmSQdS
0L8ButEypi1Eu+My10kWAGSz0DkOxlIFEiLcOuRhACwFr7qez0f6GXyQLi9IiXFgn/8ijJUZlXI9
v0NDVZQB7B5HQzN8E4eG7P+RoeSLqq2sdel3S07LLqtVtdR1mn2d0hwhW1z0k+dRMHY/Ei5+tRmj
PEav/RXdys0kcPG5DSjA9YfwdTpj1bCLOWKvW6xXBUFWDl2D7ZiYBgbEq/QXHBQwfBnY2zDuTTzx
e9+a1NiB7hGBEdu3uLm5fRt051qu2ksqJR1fIra0upx4/TSwySIkOBWtKRORTgL8mivdaqgUTwBW
zsN3XgcT9larZkE1wlL4w1cgfmdgosnYlkpCgpaa3/SGNFhWzkGg9c0iqBeIj+csl3T/WxpXptfO
uJW5+Eu3i7IrpIjCqVbcS7lW4wJfgxtVEJeCDCxzTrihpeN32csRy62MBJzJ3sDqyemqpDjPESnh
EeLav6bJVjtSdVw0nDrj1exWujVW4yZKc5vx6Yfe4iNtd8UQigI+zX7MEVUuq9ipTCM1Wy+hnPX5
0K5gbkh0OvfIU7h7bloBijq7xdiaAeeyi8mjGvJqvI0Z0YLI0/6LpI+MSY4RQKRk/u+CQSLGpgOJ
IzvHyd8MVu9kl/a4/wn4OT0Og/WwIEGEVEvjH5psoiCyv+/z6p2Rpw2YRYj3ZfVC4JwfWW813OmD
R/yt8ARZy1mxT90gu0MFChIHR+Ko3l9ry18XUBd35pS1c1BZR//xL7AMKY9tJp2bsvrHq9NkbEb7
dK9DryCVwLUHHSvKBSgfY66dHqV4uPXMFnicnD6OK/7GY/+2p5+nj3qt40ZO49XMRA36JQ/2+Exz
DzLo8L4H2waIGetthXPLI3i5zI977jeR16cY1/ltMSMbNrfRuii+25fz4uxfVtq21kaBSB6Y0KW7
NAdL/pTHdGg82smSsSyFCjymf/3Ve7w+eFq1mRTJtdx+Wua4iRyxvJC02FmdC6zyB83wIgkFLjbH
4rV6scq1W+rRRKWdkqN5iU0nYhvHOwn8lGdfgI6k3Y68HY/o2KgpX4D0Dj8OHKBbQ9Qquyq3Ryy9
s70jm1ziBSuUh4QrZ9vviN53Vcdy1rGJc8nxX8APa3ktJZ3yI33PhNTblxncMOBgknwvefU4Bp+H
o5eB0HxvoXWvi2p8ANgpJPnLl7elmV28xl89uruN8ql1LGhpYoeuMDs2aHwcgFqACSA6gEyB+nPv
pK81XdqLqCKx61EhxIhKDnqXyR8I7aY8jzGHWVnzJwm/LcLSD1LYm3Hqocr5UgOIWqpRdtN6aOux
MRdV5xkIhT+CL32VyL2+HlO5kZHKMsbGatLPgjhv4JbTKXPgf5Ylmjsc79Vp4fzOFLfYc/qNagHd
lP/StG00ve0AWk3wuue1FejOYIak+8OHoxUhKSHfHUiCJdkf280ArhKhzwqXbZJtetTDCAN5AdOi
Ur5dYsCS2JJmT4fieCD50nALbbD5KA1XoA5iztXI40yn9g52rgExTRcLvhEmAp7m6bX90R/Pi6pL
XDkIhXcwJu1ixJMY/CujUVc0Q1n89TO/kReInhu+Q+GpWHPmf1mju9Adwil/D2siuMJsuXZVQvDC
2nYqIpDIvP/QDKR8WrHkJLZ4zmuVwMNc3/ASsgCcq90E8kq0rQSa5PZH1eg0FjSgDSlMfrg1IfRv
Oa8sAvrOFS5RofyuczXZvG9zr/oaOhuscfApjtPW0NrL8CZEzYceilBdv3FMF54216409puCyRFZ
4d6cAAMEGmk+nKvwfP4x9K3Q6+bI4tfszY8apwyXphCZxrZsiw3fnkGy2bo8GxkEZT+KfGjKUjPJ
tLKc5z2romH2OO4cc4mkl6xa7pfgUb7BlaVcEidIJ0HZWuDAGREuaFYZRUApyfsaAnY+hHsXq8Pk
O1s6URsbqAlt40wnsBNP5XOvCKmM67QpfAsM+B0hUYiQHoAszJqx+SCnOB5KCa+8euHRaHNBgE1t
Q5TjtXHx6NWYMqkH2iQvfpcUfkFepsZmY0yauIHcBPgsVYZvK43ilVXWkrWAfn693hdR9OcmDWmo
04hJUIGBqBIuyqIm1cDK21eQmGr4i7ULbICRLf57Mguj1Qnz6X62Gps6jDGRL1rypsEM0utC5fsh
q7q8eB97b8ng+gzP0iYk1ZqQ+50lan5MmJRpvZP/ACqGrq2r+QWNvGr81NvlOaeqFb1UMC+1K5Hl
ITcMdt2W9l/Uk/WVHWw5CmC8tEctpO7XV2yf4wBRVW+sfZCfsVmVtUaL+YUuPT3E0XtnB8uLX1fs
Im04hF+RabqS8tMjc05OSv1ILyfZnW6a15/hKvXVr0sb6cdfngrbVNxIq30QNjEUqJOoMnG0cUGR
bp0KcVWirtq3EUfPATPEkbm1T1CtYGh2wfXucY2VfIvl5Pu8QxI/NEAwsLQ9Rgpgye42pBqqGlaH
3/7/Y0El9XOSoiyLJoTpeDh0i5qmRqeeqaXslayBtOGcKkbD6+TFQaTfIIlc3IpANDb2JDkDxJeW
QsdvG6wWA6DHo1tdkEJY9gIJliaHzrlmdh+C/DPIdVmskRiNtCVaQG4spOCJGTVgGKbRYiNoGmL4
YzmS5kztc5tH2e77eLLpJjKAkYzlGApiUona7WkSQ3lqkI3FARur/tfqnyHjPcV6cZnlP74q1TSn
1X87kNFfFDYcIv222plEwSIMYqo2chA2jaUQx3owxOCiaVuBKwTOpUY0/KjsyDj2GDgNcYA/VCgi
gdOKHRBS/zzvavqubbEIqPZKMMPvMMryXQojDu2YP0d4k3QcnpQI4EQGNJ54C1d4ATxnAhpUNGAU
NVIQSxSIVMKfkiI1eJwDTbguquWMfiBgHu1OqMsb6+SmKcHh85YphGgEZXPmFLyq0TezEgiytV0B
G+FwFx/X+bZdtIFRJPjFvGvXQh4rbrGmT7J6uzaxE584d3lRz8Xtkj/O8UiCG/aSCGLgxo46P6Ln
8B7JJl/HKmUzKLZW6lTqld7fkSFPdY0irEtkgQfPpc3GduFtZ8PTEf4lLFM16h2OHlA/lsygVmAW
58QVX4FydsDOBuEWgdxIUyfaNdclfIpZTajCocR/NhmeiB6UiFpPJM5vPpbevkNe4ocwuRPzu8m9
+EWVpbb/PilPrXH90U5zMeOHvLBEgGgvxZKBQmO8+Li2lLtCL0HDaLtrWcjAsrXvUFX7eueWHWwd
pSNwgfp2DGHzTfJRI4R+XVtoh9s7GhGJbgN17ySX8E0uzQCjEK3UOtRhM8fI/834LWjWnLX71drk
VlkQosp1R/9SQc3inHH7L+HzmVUFGktoviF17mFoD2x7VpjtEK/3cQCQD9FqdBhuFlchnqHgnUHB
jQQQUIYfkBGMrNpAidFEQMZ2MydfMpwQf4l/Jtai1dtVT4nwM2OeM8xTH/f2+RgvRfEL2Ddm+C69
kPn95cJlXEwpTnGwZSCwYL1wWS8k1cQCyHg+rAMr3QvaiTL0YPhzbQStbPOi8mennMZObJwBRLUn
rl6bxemiXleK/VbpUaDl9Q7WEcF6hv+CBEJPNxc7ASgscim7FVHY1M3dUC/dkRhOmKt4SKpsT29g
if/aUaG6M0+eNaWDxWIytxS6KUOcUb4mfG4gCMGamxcjhNniUkFbKUc8Kgj7mfOzbxoQ37Ydbus0
CDdps3c6JVeEJJS5/Be6R9VezJlcvvAsQ2x7CF3viP6A15VVFcrL/AeqhvOCV2y/Bb2V7WCerE4+
1uEjMfInj7sDW7ILR23yp8iJ6OGYypjmnVtOOzNjdYrKoxykMb/yeGxOR2JUL935vCwPtwn9T3eb
AD3XQt/Dygct8i68EqDLipqY2OuV2kSjj61CuF7+PnY5RLktPHdw6oD+4smfR96ThPwfc32qKsjJ
6UYFX04RkJbYHyytcYczzmZ9cmAmYfadRxeiohfmBO1RVThK0YWO2eDOuBFnSIqEv3cJDwUx0Xms
hGXXFu95RGTrDkGTZVtDa0AixmKX1ZL+dv87dlOKR77QLeoRsqUqXCZKOX2WK59hXWlC0vATtV/X
nzadgu7vAJxXjoTFRU5P9+yU5+zF+2JVOJXex+ViQIPg8gyyl3uwAI9Qd7RX50dyNKDRGzp17sWj
udMWJx8zeOPC8SPUn2HqRbUECs8hGfDCdohOVaZYWs5OOL6lT1ktFdHmu/xotxFxyLyOsJgSz4Kn
dSyQa0gvS2mBi3967ZuvlYp4a7B9W/YWM0/k6l9T0E2hN+QkcqpmXWTlgU/ZvidZ6vbCq8QZdDVf
FQJv7IOkFVIrUMCWPjruYQpxoghpWaEW72YpBH6cvHDSGePDgyJ2J1jZ0VhVUpoL4SFPcxzwnfWF
xGtcbGYwz77WsHC7G5dSRDiJb2AbznMKOSHZpYqFmxNmXEMv4b8VN8gi7NLxPYO757V+3YC9UQPG
93tRanshnTJ3TCi09blHUABqutLRk8JHoZoost9oOqxxXTCMmBiACEBVr1I68a1+fzXEZwLhr/D5
HxWpbHBYVtVQDjXieO0W4F68O3j9XTfEHib7GJKliKOCLlHd5ymMvZtIL8egf61mf6lFIJq76Y25
Tim8F0gvugy1L2eyOzLjmpK13w7deskYQYl1FGgVZJoTlw/FeWHD9l5aYbexXN7q9ccDYfy1JqNN
OQYD3p2Ud4kC9SS2I0IQnFabKHydNEfX/YaUed28S7TzIHkUu2f0+k/7UDH2KbewGQI9JOt+ojEu
bcHuPBwBOLKfwwxFOKA+hVKVCW1zISVSNJ2WfisGYBQ96O+dDee6CwkZnlxbTXnCkpbR8WoJ++LT
ytIsUfbCOmOTuR62tdCS/cnR6s9qStugle5cUas7Km36BMql0KHZ6JZqK6N3PPK8/qvuhRGC2JDK
QRThgco4X4azYITmA/vQkx0vCaUdGNTXS4SKVfbiZfw0KswgeOvg2zBn+a5fuWvuG+Y8ZMb+LIwT
7LWXgE2zEZK5+vyXhJSLX8yRKumDmAg8huZIolBYF4x5YnnZ5G7YF7YzOqIagVm4sHabauJHuaVc
FJk1sN7pg15qL3DueqcJhl5Y7KI8Kqkm32zECkMxK6+427tnLvrtXTdBzRlkbZsQBNE5q5ZZSRAf
wFAHW/1+nLpbXukAReOzu+4uBEfoQvFVmQvL7r0PgH+g5d2oYYXJrHhBfRzej5KNPoU0/qpos4Bx
wmHWtmulv2xh+ANlU5UymywVqlbMUsPYF8lrIRmxndYIxKgptrvEKDHBdZJIKaPUKvCCBxQJgjhg
KZo5Tm4ULXkYSRwdIf0HDLvEHwKDrfEqWjOlTnJi8pyzh3AKlvwJXbSrJLt/sRCrutXKMzqq8UK6
VL5S4DEn4peima+4NOkotHp0aBsjzJGVSW5OQAxUiWmmFmVrrf5FLQVovwJUx/c6pZHemzjqJvv9
I2SdfTYiKRx/44lrWFx+QH9ItR4Q5DmEp03J+Njudby+joc7h1z4yOO0ZfGDeji5ur3Tn6B6HPM1
nfUG6j7BFSNJCmRW+so/TV9zgLs4Txbsmc38II7EDhyh+BFnTk9nq2IgYYSJ8QOTTw4Vadk9jb33
jiib8dg4EUTf8rBYm1qw/aWenSNIVTbdTOcBUp/kOynU3uIwPvWhmMNkVVChIxUcyI4rbJPFP9MT
vuY+t5ucTwOjzEppTPk6KTi0DrdUiOdm1id5wUyS0Wi8Ov9F3z+LVKBNb2ppglfO0X0FDTPWkgXV
mnKelo9uU5JBbaozthZM9oaRHIFbI17nrsw9AftZAL7aYzBB5CNmrFC6qynaVwTwjtmsADk7K83T
iRz4XqeglPs9X0fonfQDPQHuz0o+DPQfbmG0Pal+nTPT9Odp1LbKFYOEbR8tLA5Uz76+w6DhnwuJ
E59Aa/fvPv36CgMVi/g1sFE12d26FlTedpqt1AsHaf9oTBUUhIM/wJtFfBlwmCsO+tg4cWA2kFM0
i/bRnQxLj0qEe02CZ1+ossQb/FrQIWe3un+ucpVtlM0bsm5BbjzCxeeViVFsWdS3uM1VmSSH5XyX
4+8jKkCO7pbhZhgp/YAAjcKXQM9QgCSP+F8CaS9wScmwwcLu0RJoeaFkmOdQjAghU6dJtrssM+fu
/I3wKq7mm1V2l8BEdHVxHTv+XRw2Vt0i3Twabq9nQRcoxUQ8S3UmefX/gdPCd3nsm7evWopQL5XR
zXQU/vf/H3Hmov84INJpLkOLejV/zTf9142FDcwkuUR7YwQoV2zrJGy/EpF+1TjDK0L1JJpj0jkG
YOZs4ki77EWbkh62G6otKxncZ+nrAlr0GAIlskCCP6889owQ7FhRMNqHwOzqU0gUCJLELeiFqYq8
bsEVXrrLZx8IgVR1vJeHqRNx+BFzFZiRqip8xEbNFkiHqqUrwsrhNqrBXZZQBiklHH4+HVcbeVgB
XbuLaUVCqk4MrH8BWRvCfGx8Zy/tCVwBpUsjAA4OnattWFaq/8jJxsI4q2G8lufsUa6lVMKnLhuL
l0LOPyuMLfLNLbhd5rdQN5iqr3uKuCc5HapGJ8XayaZphUI0VrdC6f30nIEtezWOJkCySoJsE7p6
Z9MJdyhRouyH0CZY1T/03kd5l2SeZZjVJLVlAb1NlpW1Utz5lXSp/MCCLK2keuZvbmRDsS+p1Q/m
qVdFbwmZUmr9j6AD9+QGtSbFYhuP1BoqaXGiKFVxOeVhbWe/vqWKXrvlw20mmDbT8pTwsok1x9Gl
MulYIjP8B7y6SuzJ3sAQpfyj6A2ZhPveHDae8CIpsTWRvnpPG36YUQBIVV/+fm+oWKo054nxo6BH
F+cd/e/p5zk9mPs2GxdploPzofk49Sw536x6JnD25r3Mt69fDFP96bPz0nqt5Y9qhBN1qjkTA4hR
Ju2DST7C3JASZQGjSzBNRPGXKOwiEWlP96+CJagx6fneb+5WHJH0+Aqi9mEhSROG/11H8BizcYRI
1j8MK3xaHhBdcj5d1RctWqLlJ+WVXPvsOxh/n+zWV2K7cSV5ICKrQ88XN9zmaJ1cTsCzUTaKCjZL
HqbESC0EpdiKhb2tgOC7+pmxShsjUOuOmqAgrQtFW9VSaIz344kBgqk/AS33R2pMsL9zbbeUNE/8
EZStGmCrJ+iK6yHmKFbH8ieXwTiMAeKRlqmOj6e+ouI6BT+5Ifn4DUAu6Ezlmy0wvcaMum2j/imW
H+pcCV8uEUqbKrRga+Teil4+iVsRGKaApkG94NVwLL4tRrPJ51Qp8T63kvHEQB3u4ZYj+w73whQ7
3ULzDjle3C+l2Jwe/KY7N01Z0F4lwSD41bxe/wkphSA4DOnejvLfJOGVeRMhCp+SpSoCPELwC93f
tcuKXnq1l7KB0abSVun19tC5MtVOIKBZ+Y72lNMF6jNzYvP+A2Kc/+vQqMobTinFpuYxjNtoIuCd
bTu+66Flfexy0U98ynhn2mBcP04xBk9Hkt9JSM61LjctGwxbio7MP8AG/EqgjJ2iql2j0TEwaxlX
04N0m/S6OrxYNyZZopkJYCauWcPm4X7av8GjEB3rv8W71K1kcP5Fa0JVZMO2sacxt+yjR/QeILas
SNgErtUQIXe2gMfeIfRLVZLlpdjZYiPx14tQ4ibe0nrx6nQzN4pxK+exn8D2fvJKswD4LG7l7QRU
3bDPA/v5ZH9vv+nEYT6BobJKjZfMfL0I7Bb1w5YKQmdbTX2NqpiAVd8FTRa+YpYQc7bfOqwRPFGQ
I7M4rHA1HYwAUOQv+DelYFAdFRK9z0aV0UTz2ltL9n/qrvqx6+66Q6+tjVO4x4QhIdrnIXoXgbgG
I7w9m2fvQ19Bwst1lMYRTvvqBkMf7lnz793TwWeqaomcaWDJNtMsBCXV/NSgDeXPYvd1Kzl+04mD
HOrI7mPnt6pQnHQqI4lZbWdR6cSx0ePWUBuSFhwHxeJAHnd4bwpgjYdbzqkIUJ5RN79dJL9Iij3k
QiZS+XTMlqPGLyGuUqTJ4DRa1YjLC31TVA+spHIC/vCn16WFHQ3vRUarihpK3s/awXrt4ki79YeF
wM2is2ER0kZXuTg2apd+4lU2JTvJz1QZ1kHBGaEanYezlImQyvBYvHWdcPcOF75viWd72NscvNHd
r5DNn3mgqTD0m1955pS8b6RTPH0JwWPOuDu10rNw3da+FyzxYtSECF4fR/f9c7tZQ/EVs2HHLl2T
nfvFWcvPjX1NxM+74OSfH/1o4qbYjFcEQTTQ1lT1zr+l9EcbEfVw3YuhpBnTXsPzMk7oX42ODRyh
MGsjke8tBn9Egtl9872MpHzHsjS9CX2YnKv5Lyk7OT1XW5PeiwKtXxQKxepdLdaCSx8adD6oIn+L
rbZ2dPXzqobyGb4uVopd+OrFK1wTJuot9FCPN3Eb9TQNtZiu+h2JZvIienx5IsZ2bvT8D6A5SW0I
uqQdLU2kapn2l19MjQYDVpkmoUgk7X1RngjbwZSDoKeU+ltByj7Rh/te286CDCnIeZQsvYvrrt2W
mBxUaKOlLJRWJOgFQyoAMxULU/XKtQl6Sz2bwNIwvHshHQfqRiuJesb9zB6MZrL2BPPpUoIpQKku
sCvDXr2z0TBEP0kXsEfaXR0Kp5FZvyVxf0+r/kDC6u88UhHUvr4lwY3R5CtfP9ZDI39iQq5H+LDz
7RDiqEVh4mWrrONttgQ781EO9c0OL1TulIEguOSTV7lvx0ULcYbTfnC3T/SPY1ARsiGsFPSflj6p
CBlBsPhitS4uMiIvZ5zik9U03dtlG4ubiAUl6q7MRLvJorrTYLCtcDftl80r6mEFGvVeh39WK5Oh
QsIBCxht/d+qkdNOpIAbTIm0CIEhaN3vjvjj9JG5vmlbZxhsQ7ZEpho7wQNQIqalfPMMmqtFhUUj
Rxryay9D+1SN/IqgKEA5xfs9j3OOwFFfxlHQTGFdlp68iXq9yhi2my2ifXcEv5J/msUERhSh8atj
2L4gpJxgXm7m1mrtjxjxGh90NhcMEE7kc6zaA4C7sXCPLM7z7YI55rkkEJc4WBZLrLlbcgIGeBWo
l+/0X+qsC4KewtQ9/92p92xCqu+X0+oNT44bSkk9oMcc+PIp7PoaXt8Kwwa7XRnyrtLRBtEmtd8s
38UFeXA22YM1/CPjTdiI45U3NK1714q182KLYP8H9gLnh1TlSSoSOJ1k/WcgTL54MvjoymDIX9IK
wgoVjLWKj++8I+E8Dn2/vXvIwR07no2M637PHJqDSaIpJbk10DOfHGG1NgcQ+wdWLr1DpyFAxqej
3mVtpilsHN8eJazN3JxY7r8LVgxEmgESClretbERdb8DFBspaWf63exfJzi34d7pHi6FtkpPzmqY
wWxZL+KzKRCwjqm1dUXn2eoQn5wF/nf4OgGpoTRdN5kuPk7yxm9Ee+bZniIg+hwPSH7Wxgabv8gA
ElHxsohvNarpPM1Idk22rmhwtGwpLBQkupiHpEtTaXSOtCDI4moxbY0587EfAWDK2voZwMqJSS5v
ZByj1uQL5BnndgkvsLhaH+1CqHUzyp7TiKZpJAOG/EYGleYDLyXt3SBwrB6RaSVm2SFN7qmjgLiQ
uMb6IWHFx9NzC8DvSH83gB6gQFS9Bg+SL2sZzll6olKrsbdEIJzlBgBfPxLxKZT17wkgyifp805V
zmKCuNg9CDlgrnQXZHMKjXjdgllhVAZApJLRLdushRRlbySDnTv5+ViHLv64hxLZMn75oXypYJVC
R6aBwIV/bbfQpkV1RxWP3Vcp7X/mzEUSqVDHPIdxGRN0g7+P/KcrluyITBKXFWzgwcOQUNGbY/qO
ap9hkMwN1n+JHGAUfCyvDgNqN4rzouVWuozoYJ7n+Tb1hX5L9qPYLqBEOiCb4ehElGNNc88xAG8l
Z+5p1N2JV1gw4X29aFi+iBf/2kfOhkcKzioE+jAh1jRSEEY4BIYxqawKEfDpqrykbGqRsKbvEZhw
zczRyIxdEHW+/Wo6fr5fXXALb57u2845X29Gp/xwDbTIxgPEhzNR2XjqPp8aSj4C4AlQNcEuiWiD
WAiLLyBtU5ZWS/xfN7LCvJYIqJcdHRHA09bxFHbgy+UT6Fo32Gw0UAlzfMZg4l+FUUML3fMciWy5
VQME1JcmlgcIr/PxFxxQyR4Y5IaAHMdb7Mc4jmVAW8z4kGGWMzjPFZfM9KOd0FpB5VbGlWO8ZBQ9
FqnDDiF0GyDdSGt13zF0aijLpGiKCS1j//9OHvoEQK3BO35LDwt2S0yll6lJFykT/lwmf7EHQ3FK
I1SmRLytrOpe3Wl0nQxHdAgtwUkU2JM4srfhrRM/Qxv+UhadwFsam95To8LeHJsEkbiMcpdRLqlP
MepavBGkGyGD1bZacGhS3H3YFTYeCE9K0w7RCDpzzsbUx69h6t4yTxkeWmjwFBJmUzjqYPh88e0h
AcY3lzr++75cTR7hFHtQawd5r+lzLmLr403SccdSXnShGYNTkZHZ7xLEF7mplvG9m0AZ9zpU06Y/
RMvTL1psOa/SLxO+O/sijXVZTR+ISCNbYjZhkv6VO7OA0HLAhbWfQxxAGK5+qAffIoROaNtmtqzS
ret+JBDMf+1x6KFxrbGLLp4uYbOMTTTJNo/uCvqdWKY/GUFJGRj/VKHrxCM=
`protect end_protected

