

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iisr0ydwFOm3eepmhOYSaxO3flYpViRsLN97vKyw+ai+x1TubmaH8qRRwK/QFeVsjlGTFdxookcr
olQwv0bmdw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dJvTzz+PoD3n2Ot9SgKfpEhIshJxklhDhS1tYcrcmprfs5wN+lN+5Y+o9jEEql61IqDkJEIGu0xp
zaDWEeMqwkFuovmZnp/AnbrHb7R/19zPRtwSyZ8+VQRLsRMgscwutXu29fTUST6Ribitutae85tQ
1okc5mYK0mcSMIggcMg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZijKIWnBSOuwn6R4ZrzJp1qaSPGZMrP8GTp+SV+Sn9xEivGxLJtGM40xMLXxiYuxIopDD/A1usG6
HkSoNT6OzxHJWKkUEyyVzrZuJdNHJ5q3s3y5LSNY7eMxN9lY4/gygh7aVIBAO9YWzsWu3HLtrHA5
2vsUFQxQdkG5OTLVP1rH68P4j/dhqr/LVHw+9H76c/knGyalpHLRC7tnHQcfuezFJWlkzaNGHfUo
b5cE1YTvtdlZVmw2sVG/GbXIRi5fq3+Okdy+JgckZ4dVWbI20rfa9LkI09/kwD3anyrnovVQVx9h
F0AxolVKVVyWNAaSu1fvXllqzrdJiRLbdnsq0Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LUajPw/jRTLlmEKb+9YylQ2jxw4jlSx/1GGaY1wFfWFdMwK2p0xvQMjui8K3EqJF0fnb3QNWuQDl
1vTtf04vcOAHkfRCeW7Mbp8qeUTtAsflGIPJDxHfVU8ZKprwANsENc8LVrpJ0WnjDFQIzJw7LDqc
Jj2TofWjKprdxXsMnu4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KG6kiSPrd66zvVpG96eKD+783ebVLVFNF7pXgq+rCyBBRoa0N9Hp3DIWK5125mkICodI82zuSq6k
C8aCiPbDiv4tiuIn19WDNNPL4ncknL0KLZTLAkq0BIQIsnFNRaZegM9aXOdMYGKYLpnjSD9KRWRt
WPXPZfwprSu2D7PeDZMiij3MY+cixttgVmNfcx9Kkmvg+1B5sTSDTVs3fqpJBBO1YslTmxyJAIC6
uDuGqvQ1138z6f4f+f8vMXratK1Ypo3jPPb4FTNLYJio5Vd1Nbpl9kRRtj801Ie0GGhbggK6IXJx
785o6wX6g3tRyoHXGJ4DGUmWlIHATg0KIAflYw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13424)
`protect data_block
xe1Ti0DRnOgz1/V1lD0S9W+lAsV1uYctp70C1VVHQvJ18kETRj1R7VpcIqt1SdVFYmpHlEeUAyPy
q+Xaz2MlsmMaH5tznS4AUQdijzMrqkREuw0wik4z4PASb7zoRgvKZzBXKM+RLufT8SkHlW4E6LQP
y6s66uC0f9PIp88VfgWwM/YtKOE5xgZOrc+waL7rbRr1IjGFkJoDL0qhHkrGtxZ/qKWu24jZZpyB
7WM9vFVFc0p+KlfTe7pybEpI3NqxJUR8Z+1ZelamuA4gV0qc7b3+dXwMyec2xtwKkDQjM0rfaNFg
6lvclkZeNtma8d25MQrdmndhzqts63xy3nbz/4wRc0BIPThD5MOlx03FfqrzVeTR9rqioVOCfrVe
V/tzNeTSJlEnWLCbGCJeO0lJcSRq8PCIFpH2VoAazdBc/oKDxoOyjm1fDOHUK2hRnZEBWOi+YppH
7HPmsi1JHoxfRfomGMpWM/FGrENEduTplD8VErZEOt3lBe7wnWIS74yJf5/viGmrbnWl0J86gd35
m+gaVLs9ADXC8DglLCeyb0YgG2u4EPfBtpXcUiw5vjUbOGdeADYHXfXknL8AcOBUNrC8iXgyqBPH
Vvnj67gPf43JvfT7Ta+YwqhHL/cbCkLG6O8w61NUIDF+Yg6YKGxslAbMClBK5VJOWnovKa/g3MoW
zpLmLvDxvdZACJEql9EdPkZ2HGIPFSjPnF/AWaNrvSF1Sd96a4nQQfz2BDLZVOcw59Z/a/9ZMp22
P+7wcYqktVnyaKPy12yIULCJkvY+alNzg1z4q3RVPL2i8zJBvc4NTENgSAgomblqoVyQOH8Jqh0q
btrYVf6ZKLy14BuqbZjyAPfC16Zh5chz7FMMRocjo7H1LC0hToIk0vBOaYQIP4qwGFIL/DguHfxt
byHBDRgNRnBaZntQCSIrCpSl0VQ77OO4cx/qGU8ruWZfg4dQCogaa+xen3/6B9dlYl4DvIX7jLKY
JRLuo5+YsCvGqhl4s+lBIiy6kiJTfiml3VdigCtNvDx9RGsVOY3YzWBjhd/pnq9A0sEDKYdXaFei
hGPZOhnc6W4bsNWVSIB0DoSlCVPT/dy13jhT1D5Q3PbueAy58vScDyQEj091O/IbGfOr1LyNQsNS
0Lnn+2xzVzuckAB2fXzXBEoI/XqFcErWOzeewbyVYQH3FrDCM4fUYy03nZRVdl971jr7GvNwJs9M
AWJ9MyfojP5BVKUPCiu8m8RYU6DG1xL83VlRdMTH/QoG6WoEb6C00vq+ZCWmrBRQqIzLI2yco295
wu1ONj6Hji90vJQRHYLgGJ8ZZof2xqCxF/BmaPIEhTtBvxTQEQCmOXiuaBwxbkUPtlQSQaF7IYk2
HRB4qoKKJ/866ldejQhynIUX6z6saN0n+mgk4VG+96mZXP7irmo3qKj3IFLZa1PsdXSXGxrF0Mdz
h1sumk3xcKe2uKjvEo8ORViOd0nN7E+DKrCd7FMx9digAL4pHK7Oa+2oe8duDPWxxwlUsp9kw4Ln
UpD5dlAVqaHCcOSS6h+J3jQebwtdkz+6jbTdt12pBuBt1WfLxzhUQe1pBY3kVPPL357JEnB7/sCN
HVnDEIfmtR+8WJJcRegVGKqA0QUgkgsLoVzsxN/pBMtP7XmOQI7eTyIqf1PEr6OIVr1M0DBa9tk2
kA/t7HyeLefF7lP6kUSOgE+Ptsj+ubAPsAjYUmyYHf3y0paXDpGDQE4kKfKKQWig0+DS2un5y0hJ
EzV6qIDr2eUw9ktm8k3FmzBW47CWObcfvzWisSh09XOowuK3vw8h23JTXGkjti5EQxHdeEvBOl0f
CtzHU2x+Htv9hg+Kow1W2XhJgnxFnFU8hmkhz3ZAGBT5J1UW8oMCaAkkd7pmepnJchll774QytXP
TuCSm5tb4hor4ywqvqxCT9CJ80ven5NHUabXqGYqGKMGXlA4qIEwM/DkYHxKA1oJI1jxVZXUGNI2
tptLxWFfQ/Oan1aUoFSW0QJULKa1903AyJFbpbgny/+3grU/c9IfJg16VVjFCx6VOYSij4iKcbJx
UGxZ3YhKBmFmphCsd3K0LFva/9U7g+Qq1H8NpfmNQEVzEbSX0VIO3B1neTdNBjXpiLiCKuue0k6C
0+6y9EaggX+eb9solWJ9Ofv0PLyUg2XM7vhdYGzRSCCgIMO9zxIY05coZYWgYkjtzJZzuXYI0DGF
Ikf2PjWWZ6qLEuHsrIp2daY69eWgk7+X8lF/a2kxRrCwqyzBEYqWa6Zjv2vUe4Ra+MDC4B2X9Od9
U/RdHtEWEnc17Z3XqMyH8BJHZve/TKCtmXs7ur/pWhHg0pBhd8ynNeXxd40xpnQmMNHsxvl2P7bL
rGvwY2m7tktmM1xyy8voUtI/nPAj6KY/EUlbA8gE5qCN08edPxUEv0sLCjURatH+pgFD6a8/yVv+
VF2mJIE8bXC9JqtAz04iIzCxMGcDAP98AsojD30bfHiCJzL6t3xYK7M8HWIJHUi1fZ3sAlgg6LH4
00IaJOFJzvxDPfnAK1oc8WGYqB87PaikeeCd1W2xCaOZbFtsWNHCHoSI34ZGSv6NyC1bytgdnqr3
EqNkLhYVbOoVnlVqU1KyNBizqMlIWDfuZXUNUUmCTUnLAmtbT+Ec39U0oIvvma2IL8MxPNeqU02/
dIUGAVjt3wRgBqwXQMOKAY8q9VD3242S2uPCEEr6ewx17XOr1euh50L16ZXMvf83Tt12+sPRm8Gb
bPydmx7eFRcEt2X/FoGjLTdBhWigm6aVPNluoCWWJA1EnuVrCuqjmuQjwNCJRoTztpZOyq+Jdl4T
0vJsa2WxDic1a8lFrGBW5L9AhM40wLLAEaNDT6n3+doEevOB32xajMyUPBGnFP6sQ4s+8Z8yY65S
JgW2C4Dlm4nbZaeSKlkPR8u7nhf742GJe4iTxBPtzO+JnHUryF7eSdiuB8kPSb1h4X/B1imbcqZ5
q5E5Mx1xcPoGteo5d1Nf1m1gRExveGzz9MqWivOtsfEbpJzjHEzAs+mlspQ4oYcAAkdvtsq+aZHy
R0gUU0Kg0FS8Vg3xjeX0n7BX6K9IrwXJzV9IQfB6NkFKQrMIRlAcrdMmuDS/ORdrojGAEHIj8fro
8vrjFyaE7itooVhw0Ky3aZg0Zel2pk1YIdPEaekpvxgdCm0W/bcmGbKRche2URNEq1r0uM+xOldX
UDzRfidTg0RSdl2/ValFxjTUll0FHCBde0EWYRirOgFgycnHh6ndVoQSv9wHqfpe4lG6oQRlxwjG
DMgvfdPPqe5TgkO3ABlx2D+eZmpQrkmxHUYz8xTl3Wpd08XPa35Wsfy8hJFb/HgREDfNwYClZd8s
tkYfMajcYBYmPX8FC/tRwXkW/mcrF3z8iw1q+M393TKEWA17OOdq58LA1SgbI5z9ScnRMVRrUMh1
ydEdHyNMSb8UXa3YOCxxhrFRlbZqprrvTVsvJ+fvLJxUo4jueg8nJBTWOBATwLsjpHa8NWSA7f4k
cLCMalVIwcknMliR8Z5APim3daczyMQdJ/Ne626AZXr+v6svWfmgJ0lVD0S3Tt1tUdJX8YEPYIGz
SYgVzmUSDfwDBk5Q3AQfkC6pKnYyutxp91yYY8shWC1Z1vsLyReM83cAF//fDinzPgB7LVibqTSn
/0tL+WMIEno+fVA2KBtc8UWXuyMgKp3e2OzL10+K4SfuwOlv+/0DFtLiUMtiPc4QehRLW71yu9/L
3Ry1NRL/0/y2xjurLe7pDgsssdNt2Abd6WqSQY+Qqzw3O+7v1/eh5ltPW/dTWVBJDur6CMg7PJc6
i3OKrEsUprCJXayTCpSDI/nQbkgRqGsk3R69p1Oaxw5Ul7bO/1zBLEkvyM2TVYDPPK8Pf91T1OIn
Irlpge2DmqsWPd36Vhm9+cZPMbM+1yuuWlekU1BG8i1dO3hz7+r6N9cqMzBZ/ifuTI8B0q4B8fgR
anGZOWDCFGkopMgH0iwNssxK2NAXUABn+5Hzc+sta8HWfktBRAtNNyqUYBejKEs8bYUkA1wsMPuy
vFpcFwJkP40u8c9h+xmXisKvNlwzaocU1gBtPNhF73om+YtOAGTgxLCtYI81AOFb54aoJEyRNJYt
AbncPrNuTstUXUd7GLmTa+kByMg7U6wXrtgVJ5A8rU3BS9E9utQB/pRCUhpHSK9jXJLnD3KCu2Tj
pe42FTrlx2NQVnSBf5hisbuNT4+2xYq9szoVakZhPTwvLl/B0DCWM3UfaciBWJCShSs6yXd5O8tD
d5CekJrKKtyA2vxAecKla1m4eveG3qWy54Q+CtLR+6ixgi+YLh0+Y6dvsSofjnSoXI4LJfHnY4hl
bnACSc84gNU6CGmD+ZXgO6Rg+EzqeVXLoqztW7ZPrYyGnxISDJ0nbtxKTJwZDf4qymnGcfmRcjap
DDLqnDoNo9jRG5pdPu1/I6RXFLqnsf7aVwQzb4APqLa8VlkdAEXZMEcPnnISweyNmT5KKCFwYMa9
jhHWYO066gH9ZU6las7Rgxhfo/KBntqHPxQVEJSow42dzqSQjF5VHw4mnldonlYapZ7hw92p4Rsj
PvVaHwmEhKk2Wd+2BP+gclwehrfNiP3b8jqvF+H+ppUpnBVx61iyM/fh7JjBAE8hsTZ+PINiw2yh
gEemBFCHNUeSzh5o5qj0h63ICwn6Uwn+hAGt+4P025mWsm2ytNqiiMEbMMO1J8Z7jisTCVq1wEzP
VLcRkkgpBlRLrzcIITls+fWdhNcyzh/sVe6ncN/u1qLi910ER9QLkR6HswGRJR2LwNPJEb6qwOaF
GgVJ0AoN4RaOR9entjlJi+7dGM6NxMlqmeYQj3RyCglG7SkQy/wdL+7k1DDuIWe7y5WonAWnx4p3
bo4uCugjdyaiOFzkWM6DpEV5+i6TMWYO3l0W2/B28cRaD2ex0uoe9aLpM4qAYo575CnXwL4/fSgE
1QS9957kOfT1ddN2+fwLv91ZVjMXopbjTZhEy0mqdXp7K9HAj6Pg6NKUYE04d+6Z9zS7tJ1ATfZI
CiN2JFNAZ7+fsrN2/o+5wJEXAV1TUTkbFXJqAXtmduZc3M/wsy9YqUNHPe3f1p9hax3v0bhAjLOh
10RgoCDacjtw1ZMuAa20V9ijfvsB1CERbz0brOEY6C1Uyt5iTmaNfycsLAyEgrEMEn8+yPQ+lufN
0QXaALDI3ZoSXZwMNzg3In/YsPZxuLOxHVa5v+DWQHqafDoGh31uKYS1o7EBGOChkglFnLicEOuC
KGv3N3lGUD5D3FtToiYGTh78hDorOo3qYAfXTfzpHx3uNTNzTdrdzUMR/IxFkQ7ACX1u3yFE6/Ij
Svuysnemvn7QmH7cYPhoQ+EnorhkCoO0sX1nLy5U3ODmq6GK0NEB31leTGxCkCXl+LGP8/EYiadS
FL1uknUTSiThIfNxhryStjnFKIH/rV5tmeLgRVBdR/Q8qrN2hgnM1MTk97KeO4RwAPCDx0auFNPJ
fg24B49ZA5j/9rkkyXHKq/piE97ksdZCTt30Dwq8HG3pI/PQtQkQzj/mSQ2e1vNgHGvKuMTtb+RH
v411H68yatp/BjLtPIWR7fGc7l2/W0f5YnVcNdEENU5V9BCzUHIBdfpm5aBeGMkvgeHJuEhRG/o2
4jEOBYRuAe59xODSNTo3lkJCsShFj1PuuorO/dBjlMje/BXrjuYQ0WVTKQVgoAOG2h1DyDHX/vz3
U30lvrx6Dp2iNlN3t1pwtvNwubu/UCIxSfDn2ZbFxhYCeRTgp9tYRkxgxhXKpGUshp6E/raRPGfQ
hgjnxo+3b4qEHMGMWxn//lc9A4qFR4n+0pipX0zubx3B4NObTs/ibk4IF/6/VhENotblU1oHYfMm
hShfB9FEwFKS5Z9LAd4hUWqWPv7+TWVvMU7ZTBew3oaCV9JAhrTHZR3vgXHI95hQcw/KzqlhiUct
pxWVO2SZ5S1MCy+yvz1GSx0vtfWckX41kSjzdacUQ8VW5CMEkKLOLdOyYI83xXobVUOvxsOs4AuG
LcyYgqgY8rSQzPLMZ/UnMroaBl3wxkrZNBHUj5cnqQLYF1TJimCVSGNsh5iyiUxGn/pk0LfL/hzZ
T7TbtA9lxMA3JfoBWyqu3boVcbUCl2T1Gr+Yy0DS+SFkaVGiUcXk9LSRLSDPuInoaa2972XNtBo6
cxLUaYKTlAAc5uQDUJjoAHSCaHM3plu+jWORDO/XldNqd59FDkzEE0hGacsj+Dw0Zjw82/5tmkJs
BNeMoouNO4m1z3lSfXYJIFhuicqkuRgIPVA5v211rfcBtYQFC3MaAcgfjwbkPddjTl9swpPL+r6E
OadjPJ9x+DP2Y5y/JXlxfw4SATeOtgplPfnRZpQiD5Me0AWSnNrenrXVWRIll5xTyvcHZf5aFiGK
fIRMFdI50WaeOv2DUz29a4AxRozMS4CfZ057/PILudAlosLZZw5ITM5rEZ3rE5QoI98dR6CBxn5g
xvqFjazWiJW0PzG/XzN3F3jVDy1ZJbG6Xj9CrSIgbNWYBtTRwlHKrJ0w9mK/887AAHwLiOGkqLu0
+Q0Z6V+viebJbjhVQdg1mmPUClAzdrZVN990cuJ3hI4bRtzwUhAoC3xqLnjpPZ2izxX5f4oEgUQh
EjxpmD1rmT9mIg7EoFk7E+kWuLhhu4wTxLF4nt1J9JXy32BVifRMq3WuIn87wTG6PJHfWT8eTNif
bJ3BKgHkkU9BkwmyHJqePQmMSDP5U/pRycHpIIjHiPPMsGzK3/8QLY0pnnH83Xo9qS460TUVeEJ6
khuuCMUzboAt0ZRlPX3t5+UD3pZczBVFfTiCp5pE5RhBv62xKzCeDTc10kCjxVCBfHuq9vx2+Fe+
taOyPu/PU1T2gSW4PCVyXBhN5uXulWpLFFk8WXhgmryDGxhH6Rp49SInSEhl4DNscWkXF7CjtxgT
VO/hkKVZMTU3FXh60J5lWKrhoOnavpFIz8Qayb034q1lRgQ/i76L6DG4b6vLDes8oQsZKN7EdLVV
y5Ks5F0rqsCsX7ldr34ZxWQZ0Z0A55ZoKPlGXdyX924wYC254S/DmWuV3oDBLmQAPcs723F6zaPU
xui+2bkzNvd8Qy+33U5rRmRu7vtvd23IEpp60UH5sgpX1BPscoFaRu/PHKVWKfalIyyfmiNQMxDp
iJ6CK69dY6bbhSjrrPcR0Xlw7NDJi1zMnoXiA+dC+oZ3P2O4Pxyd5yZcIK2R1cjGh9bixfmAbypo
UWC3dVP/cKua1LsVnqZjfly12IM/IH4VrtcKhYFNgO44i38T8BFAQXsQZo9BKzN0PgA56ocFPUET
xXp+h/LJSnkHYL81rMPimoh1Bxg6sqeTbvlMV27YIVGp+TWApk+B/iuq2WuMy0M1oYckEqLNbQxE
FaKK/1mDgzuAmd+Xfesj80HIVIoUZbXOdiqirBhZko3+foHzpNYFqc6CZ/adQpEGSMLzmzcbmjuf
GOraPrTxo61sK7U3LC2Nb7zAOjocU8uhFRV3fDwVVwHMe+PXv0kfzSqRgA1oJ1XcCGgl0Mfnz/ab
Kxajdlhx2w4sBP5ak8Kbf+bba5a6u8wpkIEDVZrRa/bo1Rwcd7f+pjUPp/hgxuYHQi86pajAACVw
tQxBS9HnXHjsIbB40nFVZiEln8X9sy1wTTi5rPiMDjB8MW8lb6Oz2ZkgtFfixkgqFZkytO2B2XG0
skLpQcrswChCrrQAC9K3hSzkZNmvyBrmolB8fYgQRGT0t7pZpZB6J/jNaF4aqS7pJ2rdUPA+FPIO
laFSBNMc1+SbHeWc8L1mjo8LG5v3p7AIQecn2Snfku4GySWClJCN7D/lDuX+gA9pP5LZqLhbq5na
m93refMqHKdNv92JzK6yYgNOmPnngYEGtmwGltK+72b00y6hvpzW/z7Q7s1374hvY5N6t11zjDgn
pSmFqmYe3HsXWRxeWCJwwERWbdxtP8NIBRaB4O8QlNrB2UdUYhkjqcf87NZ8vmQPcpsgAFysqyP7
ukHeouAmg0ryuUhLyPgpNBIYJkhh08nwP1BTsAWQbuNOXBPp7aoD4PefdzfxCwsR7fOqwy1aCIus
WVjVmzu5z2kKLD4de1b7h9Jx/X+Rud7oz9c/oQv6T5MdnC4AeFBnxYDhWBRXehU01LKY3a3GvphU
f4575wqfsKxYjZm3DLOafWsUdeudJep8+aUlookTpBqgkmYtWH9+UuYTQ+t+f6rFjs1Qk2VarE9C
JZmpheQtpKfwJJnt76wPQuixaoBHB+84IUvs0VKWRhAZPmtFRZon5P7tqOxtqeHmp0l1eCVDZ+mU
GIesg4C+zJWldSOb4ZPrlHm1rl7tWi1gs49Drf5ll5oiy2uwyx6e3GF7F/acmEcp6pDjSTw1j+Ca
yjNYVKdPG/nH6wAmJeAFTfijuuoAMaUs1rWdMnrn+E5a0CQr4UxpONqUH0ycbWs2Lrjfv3rChnhB
HL7/cgssuqR8poXn8XWb9Wva9ficYYiDtkItfhWuqMNLMltWcdo5ztQ0KYseuRPMWpab8SQ5svZ3
Y2uuZ7dEjC74OmEAk/CVr0i/dCvWfAaqlDZ7GWGk1hAQ40jwffWG5HrTEGZ2uVIzHQJVHrAZgm38
7PrhYTv0HHiBw+24wXC0CQvJ5l2B54LKbJMnbjO5sHQM6aT4Cuwn580wdWlOzyxsfz4s0TMI67Zz
aQX68QGezqY0avSfu1fLFftLZnH7LXacGh4arNSCugBjqyJqMljv3SDUKibYnbSwL8WMAOSiS00/
RsqpTSFtgHN6Jxw+S7pJLlVZE9tab5ncz8Nds9z8Lk2kxlel3HtSsdIEqUJeIGkcIn5ls0eYHRvd
KTpPSVbXtQeijA4qCqA35T2gZwRXHqtwBu4FY+4HcrWCsuPtA2uVvHtbpNPxaZBP53eyokEY9KfS
BbI6yiSYEDX6HrP+MVpgEm3kUi6mvvLwLs2xkiXsTpSVe8kYEczY+bDs7CD3SR8uZdKvG4SaI2YI
N6lBOjUttOC+IJGItveZ0VTsMd4YVS9+pf7IYEcyW7v0yuIV+4iAPf/VNj7VFhshjTdKsKnfDR9Z
ya9TGTheyEPTgNGRhMC20rKbbcniJzTFBXxpBLMCK0EwVjPPVaogLsI17/jKJgxQ+BbLKxAYIMPv
9R7mhspIc6rp2EPpI2QXciDC02OnEBe4F3Yk/NsztM4isIlhF6XCxZm4RfIsdZcqCEIQ0yyFwZPL
E7HHrYD9up6mS5DaV8ce4WsCKMXRzHY4oouUgTGNYxMY1bkSjPpvNyei9zfJsBVCqoPz767bycd1
qsU8HyC6JoM+7Fg6LMEoJqph1+IMkmT1t9D5kMQKsAx89ETFlst+s4Nf0OwQ0hYAkdVgi4eF4uZL
wtc35sIUBtr37QwXWMO+QPhWu08bC+gPAWLn519jnxdutTgRXcLaTuFo5J8bpbC4LanujQP4UmJx
V0NGHlQBHrdO6n2VzW8hmdcf1k7/W4MPM/WXpjU9ea2PFfYhf4R2rN6e3CqxXF4ToRWJO/6IZY1S
8XXSyTYQRKmPB03CK44pGmO3XOyxSsvExOBElLtW1DA9uhbSKhNfaYxXcUbtsKokXg7zMCWVJh4j
VA8BOopqdxxckJhRtUa9TWr/yvNPDnTMIPX3DuxTSxFdqukpd32MxVuzhK4uq2+r+BAliobKg2tU
fjZf5WMD+u8EEUeczdvobyGss2rd2s/A6NQyyd9gSjKM1IunqvKczYqiIqRRnBS0Mxfu3QsUaLwC
ZHUZD8tUTOzbEjv1xP4KS6baMt+J6wz1IHMr9nYCx667l3j6RdOpRpSDZh4TOUOm8QTedk+xeWtU
5oQWxSZVoyXQeOM+U0GbW51am5uLD4Yt9oFJNZ7Z85rRoLBKVUZPAehFY/WizzzQZt0NW74zYMGc
tlzm9YLZIUoE27qpLSVMDEwu002cYQZwA+Ov9bgfilgVW3rpJwnQSPi6sFMSGzGtFueQV42U/0aS
r46h0qYDdsYQVn4F2YyRsV4lxj22cbhkJwYf+Po8qdZlaQ88VD3bya7lbX4FQ/+E4RcLp3LwgD27
Ozldo2bQyuahPebl+8MX5CgrQFklig+Zlojyxzvm5T/s1o64kmOnsmAIptzojV1CxVXluoF9C45z
1UVqXxAqVDBO3Koza4ZuFHamE4la7OMsAM6ycMLnFfjW2Pjr+wdEF5YC7NmubtH6pl1255qlHflY
H63+Xzx8N5lu0SrkZy1P4NqIk1UknH15VE5V9FUWKmfyT9PO+Xns2Vz8heax5andajNeKZXyDq9H
Cwp1Zm1175X+nDIB7gqPpe+g2To7m4q182s+l6TTkCH4nnFtDwTP9YWtJrI447pGhesddHyDy+D1
fLmDnpSLX+ZPRQZ0tm8Xwba9x0kE++7TC4OGQBSYm9nI6vnjBeWehh4vlm0yd+GaWBRghsWbqyHd
KQEzitaIeqcw40d6mZDVTU3cVDzF4VACUxzd6z4Rkkbbwowm0ZA8UbeRqM3GSIPEzxCCdQW3S94P
8ULLiI4d4stMH5G1uothTbc+aShY/1+w4CdnQLvz1BVzwIRVNPrBa1qmbgR9vQsWu5gq/9A5tgbz
bU8qEJA2dGd3rTuR/sb0UC3ZwC02O2Ftg08mQIh9pegGe1qV+nvsxgE+I8C59nI4e7EAvMif6Euv
Xi1nc40XGbEwjXBj7tqk6xtw9rKR6AIBsjJy/x8C+HotACCdl4RrYRjhtEMWmO61K4Ime/n4yoQF
a+sz/SrB2RiJ3Mida/qnBkIRiIRcelR65Vv5SkYw/qI3o0F9kF8JAi+0tKLJxY9neIyKhM+PEcIK
fD3lShIaHCrbQR0EHje81wLeMT76aWH7gjD2gTVTZRKMv/9Pe6D0QpFmJiB4xf4h+1ZbAriMJXFE
c1g4tfq4plv1j1EKgFN1EmksOn9ufGnENYStCNoA32B+EvocYY2HI7hCFMCFu/OEcsrKTTdZcBLR
nFFmol6OpPqJqpHRMf+C1ucqabGW1gN0nCyFAfLDgfHRy0sCihy8LmrynXitFOfjeqd8ebU+zeqJ
iMsjkkc5MTBnn+mhZJS8ZzjGaWapbCDgdAhMemmsop/MOFsoXCm1XIbWuY6hnTIt1m8+7mFrj7Hm
SGjBAyd+J8oxyB/JqHZR3/mbuhG8pBMusfIvBfoKzSytoUv+sVRBD3NjW9tUEWTpzTXMRE6oaTVf
UbUcXhXld1ypyW3l0Kc91a6mQNSJA9KIq4mDL8BHkshmcAF2A0g1w7ooZk+kmzI4t9KQNsXrJ15I
nisu/2jnUmRWFHz89H60cw47zp2/zIBGZtiHnWJT36dOGJTZyt38hCISEwYW6zm77LHRJkrGSE2r
8cXrNQEMhydzksc/pUZD6dxF+Ot/QMRB2x/h7B/g9okW2JcDYI3yVIx+WZ40M+nXNXurWRjJb2pg
NqHVkR/pLt6ZEv1O3RG7t8oFU0rgUS8oMVxoTgqhHH6Ch4nkcZHSRuVwigaSBTKT0qREr+rxR0v0
qeXCi3FDlVcwMLQy1uXzrxvj6gbUhgEuWpvuMa2Bea7zI/Mc+JyC2WELh55dEtEQ1fZe6yf5408q
AjMmtpfdf83r5/hC5fLEYeV8fuoW+3ACyEMvnQIjq2CBT8oefPj9v/wTT4B9Goz9f9Ufc1O4PRiG
Cs32fz8fNCCtSpRlbOYTRi3Q9Broa3Yol6O34NGoncIyVo1nzRYTLz5xuQhkcJxv7hLK7IVHBVMw
O5IWGZDPUKCg0n6iUDrn8xQeTE2ECPp/Su9OSh9W979t5BUjw7txhYf8lRVlJXNq2xt5J95LmYZe
ld+5ANCCAGB+q7Goz5Hk55PvmXH2Ak7YMx2Gt1DIzkhFIa8qFNbPnUv3j2HarEILHNBXcNEA5lfB
1ydfpteimMOpI2tOlw+OyoUNMLdQMlbIrWkBiIOiut4dtmvnFeq2/H62+K1MP2bEGdTM7p9HBlB7
lCRE+gXR8ehAfWpedHIxlyJ8K70xCtj6Hgu5HV+URcADgD6GyIMfSqqazg5kQfgR6E1a5fStNEF9
+WrvteHfmxi4EJTfyt16l1WdTBcx2T+VoeP/kMOFSXMppuRZ3Szw6jsTRmVwCeYD/6P4ySVlZmQ9
OUbDaKOwVfbSO6vo7Xis74tc1S+na3RpVHMYRCCm+3pPmlaKdF0Ua0Lfbk0pwKnJ2BeK4g3XvyLd
PjD5nsavBGU/1NSDLmdSZ5mYF6UiIbykYovWgpLqT10LvyenPjd2dy5ljs4mIZmj+0gbjA8KAR29
Jks4anYsepcrmFKbYohbpt4+gq0oGCBB3GEiCyttP7a/8xANs90MdiZtHbjEQON1IW8iYEYzmY1q
ueNd+Nkwo5WuLK27Ww3lSe68fzt2viPiGza2FqcSvusplpfusV5V05hMTjgX3VC4LgV4Re0n+kTq
zwXbO/Q7nTODq2heC4CjmBMbHae/6f34DZ1F+AEIRsv/nEyVmXhl7iJogN0iqjoi5dHav1tI6Pfm
b55zKVxCHI4jvs74KGclgwTaTyJ03DhZfWNljbGi1DhpMAOCLdqFnKQJiGCW61BiPu+l0eMvDc+R
4bcaF9kc5/na/OWYJSvl4KFGzL5+mTbYf/N5408rZK90lAGcAXSvHDC25vfHTtbI0SXOHUeLBm4B
tvCFte/oeBQr1zQlG0LZKeSZDgtcCUlk/GSmO9s9xPJqUcNyggvoa9MUyQt1yI7oc4pZXYGak5nD
7X77CVmZ3b5hKlL+SFSM4g352Qr6dzwjcH9oMVKw3eRTlkBTQGX2bKkamsF5eWBKZ38p3cnX6Za2
MFZ66g7PG3Jzeidp4oS6GglUnArl5lG3DM60aSkdeNd0NfF3PKmkRQIRnrrEZt+XYjIShw1hynpf
/dAcdz62RBLAkxPSYCHMi45F11/UwQV4uPhWRzfsXCHfQu+klFl0Xd//WxSX+rLB3RLVCQ1qBNMm
E7YNCzkZr8TwHqTVG2n7E4/tFxdenNrGxanYfFYhHLhG6wI5nl9CLQXjZ3GhAN6Sh3SkCevqBfEh
5wZF6Jwvj5veMZt23kD1SfcaPlmX+IKlEawzB33tM89befkaxMCG8rE6ZQAdVj64I9NmNkxhEcXV
0DbJ3UMGSoenHGGOimqecUK7Aa98TbX9JfpaQ4stH53o4XKDMYmvBkcZPTFCb6YXXZw71cvOvQds
VAyKzQ58i0pxSf1NdOuGCn2pHttcWkmebyIzqaBcvFt5lN7A+wsEQSlNppt85FA3AhNt8BNitDnA
vIa+pBd7PXaJRNNQI+1xRcMn21jm5pHP5Jsl/xEVDwPnFC/Y435/UfsoiExvgqTMY749h1RFyzlg
lcKzpfmThBCn3PMxCDagbnINJElbj8owysiX8mnCBxLxglezsR/tk2k6Nwmj3j1qO0iuf4U4GCNP
7Y8KLSyIyEWh5TWofkDJBGv9b/GdCNHJEedhzPFmW8KLG3tdU4CpttUDSl/GBWddatmMdeFInUPo
Cc2/gsgKDyLTrBoaP8ADgg6lIf/JxFfs0A0Y7vyvVB13BgDdHOPlMCgs9bnSOEdKqPRJVEws9IOU
xRUafic6OI7i7jpHIXTqcMCrIP1RD6JSeeVZL9fXrpp8aP+U05bgPOoZAedSxEU9qYt1j8FdS1Tk
LN5kP6gPxzFhHti0HNvsOqV/ezrXMdxGQqoMuWoSTlssm9X4u9aDC77DmhE2yECdjw51YHfi5GvD
n55cI2UsOvPE6PlMgVBlsRr0BQNlVevskPqYhB9NMdMH0VTZ+QMPtxuRs8Aezvuf03kox8dJs6xZ
H/iSz0NxG+75YJDLbyPhMzfjpO53dc5XP8HxBMlaBi9LxpIdxuQQnwRC79hiDLpswhnHGorFnp4e
puaoNiUOmQoESUG4/a3vyOyidXgqEkjjUPao8URX1aI9cIACnlfR86HNyRlKKvg38s9Vpq0VcyYM
qz01la0M3f0WikVtZuJSukXqn6dIgN4CQBu4+NSgS2U2Zx9cwV2xhjG3m7ZOatDrFm+SPzCb+ojZ
0uDBQwcmheNPf/0uqzSaeUiZPPwXNzTUk6s2j464nDEw3vuMzBALatVzRPdXe+e8gq0NYDXVKm9J
ufh2ts0l/d3psq3W4Vx3wbydxNIkgaIITCZrR85PF6zHeA8eCmU7D3tZD+mcSESZsz6jh4HADcI8
h4GCkx6oaEQAj3VDmTgxKkvXdgLGSPyLotVyNn2D3yWuGMiGD/YAdomroScHT3OnFTA08SF6mbb5
JnFjL+C4XHILdp0hlHklPezzAfgbPA0Ko5h1iYmOjM4iE7Sw2f9b3nyWO+uDK/z+zuqIaiCFeF7r
aL7dfpp7AO7sy+aDlu1SMUtANgL833nmRQIEK9WHyokk5TAdEgl3Ove+pzofZkJhJC/1S8CQ/qtv
UkGZ973Ilnt50+cOu2Hpu4coUlVSI26DtFME9D0LuDkGlySZ/N+GsUg33tl7GAUVN5UazZJ/f1dw
Es1y1wf5w7Rm1lzXqCTSkpTGwgw4tPq/IBGAHDB6cVvfKuiRqIePVFQf/WlkLptfj/eZclPDbK20
aE3tmpbnc+wa0JSNnYDwG0Zn1Vx1zcV0uwLahWtgQwB1f3+N3E6YW9GvijxakOId6BG1zz8J5abE
vBinwKAteXIBgySyNHovd+cOnfRTiQTiJDT4/rkBLGQdklZ9NdKKPVSvmj98ARJpLoA2CEPez3Jx
uaxkR1ERsvk057+X5VSwy1uLZX0X1/GrrKTNtTURs1ozZ+brl1ohrK2GNT09Ky9kM2fwlr/PE2Xn
rOUV5TaJQlO7h1m2WxYAlhfgtRvnH2dh1xpFu7DXV9iMw55Jq868jOTGbV0EFjy1F34Tqc72bHkH
giGk9qKXvJyYmTVZV4mnVVMcAs3KsoYct2W2vvIzCXmbmr/gl6q7gE7dwqZRJRapcYRHFamG39cI
n1npWA1ivhDpdp3SPpuvKn8MgHKXiCuaGHSvDIuIh8FjyETpMV3sWAecl/Hv6JY+5Ub47lkkL6YM
lqV2XjlVBbDkNiHwx0x+ksJwC2osjFBj7twUNIHy7gkkoLxryJgD71uzjrDUwW6TD6fCJ6OWwwoF
lx1eOWuDVcCHys6NgQPrJBBDLtpRjCcN6cAA1nIBjK0mQotsnagMnzIYPK70PUfvzcrkX3xVGsud
pxSvDFkUDhJYtliU+jscMS0qZNGncbJud3gz5g53X4hj2myu7lG0Zv9ulc6v9khWz06tbYmLY+os
HIssmxPvHM//W0yKoQuGrop+T5qTlK3QodDmC6EXtzruxSun8zlYg3IfLToovp1Tf4R3JCscxusH
ySbFt1US+XEV8N3zCnLejymvq0RZBsl4AWv37lbdSp9Cjr/IXh4dSjiC6Q0tp7m9qZ2QHjsSHy9h
99wgekV/2Hm2ngS3a5VsQPs0yK+xbNgjfh4wMe+yoTNkbyen7ad7Ger8c8vhPZjtvPk5zSPXlkBv
2nN+8JMAEgiIpDRyx4LrjSenGkbESftvFMoCuMwNzlIcrkjbP/a6B1DwCizrAMtfMbRTbpQfLK+P
PI2wMEssVK5JMY77W5456i4HTURFaDcMdzBJRMW3DXmnNpB5//deomaVijnoHP6cnIMCkGLv3+5+
9h7s44RHQuDx5akKz+7h2pRB5FgCIe+ZKt/MmvpTNMPPk2anjAnEB06+KkYySUDMGaPS4aX/H9dG
OFDbh4Vp/WvuONecbDZ4aztNraQVv4mADedUQRtmcnqUsBUTeWQdi6hjzjPybqvvc7SoDTd3ACFK
75azl5dA5PzySQM23MuU0E6kOBQPI24BzPNNH6ICmxymUo9aOQY5irY/TR5em9VYsgJLOyuNNW4v
+uIF50BtkeBcNwIFxMnDS9eyd4t7qTZoCZiyiFCInIL9sqtGJWsSHixVf7HZzYUjhZSmvjFw9guM
Xv9QHi5QGSURTX+d+CvC2T+up9F4/AkSr2ta47nlcK7xOLUel7VIEeUFQY94WTgm+wi/xUIpiThr
/qYxPyWNPZ0TEa1ljJxV0VLEwMYV8qTA0SA29btbsE3koZ7sZwXoJ7Cy93O63FWWrxZrfsePQljg
QCXQrR/RHP6DGAPIqZAtIsUhvzNIS2+vR19HH3aqlrrG0wYFNFb7E24mPVCSvbHLCVkthWP/4YNV
3KtP0CsBoYE4DTfw4VDBJrqATiuYIVeESlZZlGjZAvIQVjr+SL/ahHSt7LdHoVbgQl1kIcvS0jd6
1JTG4Mg4i6U4MgOEULxausmGn/pbs0b7/h24Js/TcN7n0OL8g9fWndsEitPzeLL0m21wDKu0/I9J
dDBrSvaunMmbGTmbixoC9OsnuK1pwpRF6uWro06ESp5UwwbOzlZAJuJQjqpWnlwo1MjzxsMLEwTl
Vyem8O7C+bPREHxui0ukormhf/4UZQFE35uVHIzepDJQZt50uFoiSEmaBWD6DWTYBDRyZdbQCSLU
4jbuHJV2FWkJ8OPycY7BQfp+i70YRdM4drS4BOIyU1+Zf/UICgL56TXghcVbiWzFln9CcsJowNjF
dAZeGD1fmJoejvUKoNqTMViKhxejMZdhCvXWdybcRgo/epknoLkdDDe1Q0cks5QE02lKnObWLudG
CaiTogv6njFIy4YbMZkibBrCFG9Y1UbEKr51pHe2Ab2GPgFigVUtlDc1gIcZ7aDcCGO/L7gNX7kk
BuUNSyPyPIKdpWahhNCm20uMfHr8wiuhW8rnj/GcH9PedkpxAsRipH6BUJ8c7YSPtwAx+CKmv9we
E9USi1fJC9fGnJTtla3jEvnWfwQgfGeXI1VLOwy0CpayXtkat8GfOlWWyjqCXcVSIuwmMKah2X0A
IOj0Kw4EmLYDg6ovfaAhswp86OzJvKzfZUryt1zkzoU4lNbPWFjS1fhoqOcPJD87s33LL632Srdo
gbF1naSVUKKyvconeWFJDXi9ZTUGYjIFhP3PC0XPdG9xCX4gUyraeRnk86BU5i/K0LszrG1GjU9I
OyBoGfPOVzl6J3WN9LXeyb4ZC5GtrwCcv1vyAgXG7inifWGE4BCPTyta6OPvDZ93rFypD0RClSEL
0S8p6FW6+BZMTNYrnS5M9zYAxcOhysKUkTsxUnx0LKpnG6+5fC7HE5Rg37q/RPjkR4ymy9ljUamq
vRX8M1udama/mTlHHiB4XfUAQ02DlUf/DH/nA4mPlWuOMOMwtGQASp0WYvvbXESHc0CGP7D3zWTh
Z8lDf9Iz9CCX9Tb9jHP6h0nhVgN+Wxg1Tj2InVRrVNb3OBGlH6yBVH9UpLhGAgm/iCdDQIBGq3o5
9mCJGlenNmnZSlS6uoEn164uHAFpzmzoxF36tfCpUV+ivMf5e/0qyOaymFhynt9tWujzVY8NLA3I
wDu7MX46vXBX/VDkL9Kuy2sxvGtRBF7Q9mJu5rY/rso1kZvjsB3Rmg13d/5uU4DwOsWHSCbVxKTx
J6VcD+cvr/3QtIZTHcG83OTe2yl2pTEcAUk3ToM6qthGdwl3G7YZRX+1FdBvwCuHoqJOgtkhLjMU
s6gxykNYKmbd1Tw++0osOpPXltHAZBcRKdv5S0pl64zypcpfUtv9WH8z4CtdaCZVFcCRxUg/qJLv
DwiBnH2Qbh7lxsN4O4pi2hBquOfnKN4RjoVwogE5rCbyjcLDOmLHR3FqlFQrEOGPfYiP94DSBOny
455aJGNtlJdmVGJhDGFb6GzpphH2jQsbyZ92qm5M6GQV7GxDbPasnLdZXZYTs4ebIuZPs6K8LgxQ
8hWs/OHb56iZE41d6e/2qyBwsg4ZMByE37w6yJ/jmDDl7jbMv5O9rG21a/Olb0i279dHdjx+C7sl
Hb864jKz2rwl2F2ug/Gl89Oukvyv9jtaITumjJtGDMaGrrz+xgnC7F5MFs90rxrw1vpu3q1UhR7q
Y4sK52T2wuEKfZAb+ilHYsVR3YHHRSyNqiDQMcw=
`protect end_protected

