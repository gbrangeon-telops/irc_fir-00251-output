

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7Rd+JJS6BPhm3C8uEMSjtB2IOpOZImN8ABL10O7dB2/wknTrPPVnggIUugEe0Un6rsHScVa0yw8
WbsjeU4skQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bancDuzOXzE/C1Vj5QpW3wyih2C6ymZ1vv70urQ985WeT2kXc7KQyN00fbod+1ycgrcEzdZs+OxF
/cQLUqqV1PAWyHyEqXlxABFUHjs/nxBl/f/B9V0jlBhAzKCCHBVtW+DFv8KpHE75Z2lg+r4JTjg7
zQiXYHxUisemJqUJdhA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rZMEEzwWFXOuo5snJgtfZx9Urf7eZRBCxLhuSc3DgaT16zNB/FC6Qo2PLk9pQbhTwkt+6VFrAqaq
rIuJ+6NqrQaj6tzRnuILLQxRIcZaZnlaNGPM0QELT1/pgSpbDRVs/w+jfcFf6hDgLWdb7+lF2lZt
EzdkUS2z3RzGxMw0dEl0kPzX4BrObwXWpUb1u4DD6JMZb6O50zBS5jLIs04xzSPqxA3PuLRWpuc8
zAMmWK1PCPqsF6JmUA+ToDlUTA4DP+Qb/r/OItKXADHbpGUiJXq85NgUc8TOMYazRmcSDk09joNa
rvnt13K7ONnKnXu7DU1cLEZpB6zC/Q33/JmxrA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fSUvPGwGSOzh5U1OjbBgxWaXchd+ErSm3+d+gvsNPzEzvrhBDlsbz7cjXesFumQgP32hemPRlsUr
lFspe8TkimNAMoMtRIt9Rpr9MJxdvSAJ2AckK92TaQKYGICYWnAAwRZdM4hFhKQynq8onwVPOItS
8G6qhIBnq17qx8rO48o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MVMseSXR8Gidb6hUpBeQo+a3Ho0qfbo2cQ4XmaaPwOf5p+bpngyRNVgFStTGlS9V1Gq9sxZR8m59
KVYbqvyTG1F7VywlVWjcCzm53JiHqc7770pyh1TFlHFmlBkxaKOZI17/BbAJVPtrgC1AFUgqJIKl
KWFzGNfBnaqYhwSBpkZVKTp2N/RCKh6/dORV7jPLmH1kXSt5iI647oKA/xzmV2IPvCjRau9wfIMP
3BcMw9SliL4YOeA2gPuyEVJdJ+sinBGqyYpGCshGE4syCgACrJDHcCC8bST8+Ee2RwROkSw85PvD
RmNqdRJR8yBkuN8MggDeHwsPe2oFAGN33DaQEA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`protect data_block
uhtxmFzOzfwWHTDNIRgemryvNltabVHzw8t9PqIVuTJBiGc1RD5nTWm1zxCFkWfsTdqMTVodHoXr
cGZkdf0ZRNgO4bgaEiWnxfr9Xbn6/CdECA1SnIJSw1Hi6LjA91vYObiYQ4SkxwoMj94VPVnx8sfi
0touDioxrgDg64Cf3/ZSoAN9Brsd6qlHN3ur6FWsFqsljHluy6vG2U3/iPOxInvUVUc4ft4zSjRm
Fj/hNVpWS6mLczfwxVw21wv2BjulqEiKFAm0vm4mqMMbA62rdFem3zUJPZhQaL7WyPhI5ZzTAPiC
kItQmtNNwO+aUYk36ceq2RoV7frVg0mTn8yLTuuc4ZoI2dMVDLGQVZf0MEdkRjlHqeDhxVWCFiWG
Z0OnUl42rEkamsX/hP5/EeFaahKBZXYnzInuffSXGO5bvxEA9OITHbtToQ2S9HGt/gIyLYnavpWF
YrsdFKYkhS4YC4S20cy6y4gXn/6isUmJsD7thMowy7nqg+621ak6mLYZApV1RWagCOUlzppeNAmn
q58+WG++7cgUC3VZDtBgMK/aftfmp/lNjvQ6T+KpOoEfmQ2MTHj+wutf3FDHRwwVlqFaPZiQpJSP
gr9W4LP9eu4u6RS9RoY6jqIyrm7cCyWG2sh+AF6ThIQOH03czMWqWXaFPlNHGYQWMsq98MpmINIo
Z4zCq6Fc/UTVf1g3SCykbVgAnWSLDm8ptJwM/QNvWb161vBE5AXMLGQ6Mz2VR1/too23bDozytVy
4nIXSQ3XlKxrHSM8JAfnkpiKhQSwTnsZBr0+Y/hDQZiqx1E2EFnyHuSVbnjZ7sgoZ9sNsrwT5zja
V2riLHF6vZbP8eu4bhAcnSzHJNzHm13dazi6JOsYQk/L5InBhRxLTavsQ6CFykz7twiB6Elq//pf
hFFx9RlzXYYhukPxAzayH07jRt3cWgLSCwQqj4u81I9pldXg/zWSo1kDogXrdbMq+tW6tc+/8L5V
PTz+9hTCs01qTxNAzrALGxTk2KdWz4j3mRfLs405K1hegxMIkmPgiw4xAzAeFyR2LN1mA0bHurKt
JueytBbQoKpGMR25YecN1BJysGOUrJ4IYsEgHAV2YNbfXqKQ8vpFwOyRJrhV5+13PBhwmwFPcpvl
gxZpEAncoHbklApI+70YWHjG9MOhKJT23ptn/nvjnAfZr2b7OJ5zgZXoyBuG61bNZoP9fO84M8Rh
qeLZ50RWJVW6pG/+NhFhwdSyu4ntfX56fcdRhbZdmsoCYEZe43Kz8YvdxPYn0j+Yc9LBcSujO51R
Go9vQC9df6h8fN5bSIiHtq+1QxxWdWQh/iKypoGj9hXPGVu6oq9m1LbGLVSQqr49y4WL8QT4/mHf
QEHzI058jAeDzGOQxcNU7WZVXjNVOWUAwT+ApnyPQJA2rhCStUrIomWB4840s1uL/ki87R3azJRz
Zp2GARW3Wogc3GN8QYzuZRj+I8uLujfSVdYP61xEG+09P6qr5e0sAEgKrM+g7byFNukaB0KnMmU4
6NLAMxQCzI/RY3IShbv3KPEEKoC3p/kPr5HLCVXgDIL5RbzKtEy+RT96QT1dFCIpIBr3GD8vH/mP
F6X3SIiQH8xG5O0YlzjSc59H1WB9B8u26gnljkYX6Rlw4tCzKCMGv4ggSRdwzAesMWgyaI0HcPac
3YXAWVTYrO4Ao3R4ccyc7PkhPpBbFgDqLcZKCx6ZpxqgWvgecxr10j6PVUDmPiH+DqoEjF4xx9jn
uHF8n68ySKAJmGh3OmuJVp/b4MNbcIV1Seau6y3uX3gquOpzsfkrSKMz0eoe93Dej4RAcApvLK0q
DT8xE2D3mcpgfjTw3IU+4ibi/fzNesCzcozIx2BApgSju0KkOjKO5XTA6Zflxk1pVSbh+vwo2OQf
vOekObEOo7A8LvIl3LSW076iu2279Znv1Kx0yosI0B5I+97GeYOM8aqMEO5Kg5V29JavG6/FL/Wk
BUIpv+EmHiekTHQXeKybAYka6/yUUIhok1ygVoh1SoFZ3KDqe5jj7M6irBpGxyjZEPiRO6F5pC2i
mhFPVxOOTmwpKUsex8A3Ijyscr1LW9Af1JP7TUqewpmyXlooigZ2t7GMLi3/jRHQ3otYREu9DIZI
uVA5R0vSdRrJGyfsZgbbitEUMtdbO4b25n3G93KUGAx7ukQRdWiyj3iFER/+gATVHC2rGK6/18Z0
CtK7ZSt502HcapudWxXYkk0EgVY3Bhhp89SzerNDnJKMuQme0FnhsnntipVyBPZ3fYsTbrvecusX
bXRAMLIyNE8RN1rFiniROroHwrW1Ynjqv+hr7Z0r51WKyKy9lolYLIhU35QH9MGJBhwSeX1tU2Lo
P0Kyx2SMK9wC2D4Fm/URGN2FpcW2RTSdH63YHRuie5hj5AfUHZbjZM6YMfPapatOt1NNgMIAO5Ny
voa01umOYWk3FDuYEJzVdPXlplMWNNjL2FVhSTT2WVuT2foxstuReF9W4dO+gcJ6cQV5L4CsQ+7J
+1dZoApEUhX4HkwNsxBQfgo70TiDozBCs2laLdKIzgL2P9qagc0mYtA/TuBnddK4cxhEfbMbXCbr
8K3XSEFkIylLpdTtp0fCNelKcQectrxBdhxBZ8891AzlNfu5IRdNJzthJTroxkKOK3yiYAiPhHsT
3YJiq6o1Mr+Dy28KoAYG2lSLbv/Wr31jaMlhDBucEdNgZFa3XecA1IQu8cu39k6g2jh6toCf5Uj7
hfV6SL4cb8nC1C8X6eqMuH+FhUAUEV+4lpm5F+O2ABFSkD7btSCs9l2CpXyFK6qSmaFuqKZpaQfj
wxa/kXdMOA7OUwvotWbeEkhAwg6VCNA4xNJd3BuB6gpLcP0EWeOdLCP4aW8zkJiUhs+87z/trcbr
/q8SD5JYbor/+07L6uJfxDWGeC6MgC7fwD01U0jAaYQtPUmywVGrptVyrmkO0irlJHFTWuZldr+Z
tIGyixTkm5m2QR4pdiU7RrEhT1IJJw+93T/tpIgprVts202fT0MZQ82ZZGjkjsogZ/yg4h+uMf7c
TbtXhEGqU1a57r5drnCbNJ5Ly9vjQSbR9A26aqxtso3PG/7htKKimYW2RuxiGiOiV2jg5vfSVlLS
FUf8kocFD+F2sBUNfoDaTbULz69GCeDGLLZ1WBolYbTy7WGrMkesNloo/eCydaEpgTBJxV3frNI7
YlBDGgqQMFoLVSJVfDQ9n1QVDVBU47WRUkr5pVK1CUCPVM1bM+F5BWA2qHS+84Fma6ZWeDkMJpUa
I+szDnBILzlOTxLR/phFOR+m4tTInlSsOcn1W7Lc6D+hUmee83yyJsAZXbqvymShem9eqZb9iVXS
Jhxo7PpHVMj86PaRftBKjTXLSCszlu6dggIqBlnBNiVF3S6hhIJT3OT1p/zcMOxwh9rxCcl5NhFj
si/Ns03xyafT8kLwmfqjX5jI6BFQgkwY1kVIjeKDxg805MtAtdgK1aczynIg+wnwERBAUS21Blmi
NXkyNBQfzGHLB4ceOpXKWu/O0GKjqZYGgWKTKVONRvK2b7hEWXphonduRZ8ifbSFdUkMKePaC3Is
LFx2rwUoC6NfdJX+6k46pbL4OwgJwwKG4piqjtFAG95Atih48yps5B3RLIEMmurlS+92WcFftuNL
PiIX4yjCvHgNoD00PxDeYZZ3XJjgBIxhGsFmSiz3/+fgaPVxEfyArRCOt9t7sL6zxKUpi7BKpxfB
yGQYhflp2gBkMNRSNSRs2GvZKlxeLuob4OEv8LG0GwZh3Fn9OXfhE9q/FknH8FHeaQ0UHwU0CQQ3
Xjjew/uZyvyCvGOTvpoCAx47XisP29gwgMUzTf/0wCcqRW//rAyeRy95tAMmkEQQThClQaAvk+Fv
E4zknzMDfIfgpdKVEb/dm6fg67GN5W+cizOkWns5a7RWUdVXA3wVSJvTAtPXO8+z7m9I5L6c2sGs
TNOln1jm7WIDiVRZBiWGhQeOydG8oFXSWf7wRqI42s4F6hNYrBjR7vDALsNrZ00gmt01seoa1VLH
QVTAQ6Nokmi/WDfEH2n1dUeZa+niHyWvxw4Ftsoui3cVzAIW1uWGjYfDIYieSY8d4tNc/9Ml2np/
UKsvq84BW9WuJmjyi6DQcc9iR8fRL4WHSdeX7WX4ajIeTtwdB13NNTVRmX1FT9HQY6PfNp+U+iQD
18aqDz+xW30lLYPo0zDUyAuPwCO5AstWpjy3w8chfR7ccMIlPB/nTcGlg+sP1ZAqRwb+ZmrpqtyY
oPiaRqZiR10JH+ZcMAE9lOQ4rymsWXqJaS8NrRKrsub2yAiYxMSfkx0GAZS2TRDMPm/FeVf66Bs/
6AGT3OPUabe2mM48V3vdgPcaq1Lj78UfTgEY37iprTuaMdeXKuN7EUk1j9Ay15gQqFw9yvbfflpM
UWH4EL1FbbWexv4ZFJzzkrVm7D7eOGbuOHrJv2PShnJee3tD8R8kPYN+gaQ3g9pZnlI/W+Hc8o4k
qiAJjDxjy6T0BvkM0zKS1iqXAHxSmhFSdWI2QnL+OWheUZ7V53DQrUAqoGRH3VtcL8Bv2FdnBD6E
tRUSXPnHxGb5FrCSsPwb2tGVXYn6lVRmFQoQEYz3KVSVFoTUpZO+8DK4pNnfl93bepgCiv8ed6IM
assX8014B6SN0IP3YwsbDR0JWcAnNSGfhtwST+Bac/XX+pBzaE2RB7wLcL11cyFNNxtYTFMGyvoi
qXNsXrzwirP64bbhvjz+qxc1d9/zrD9UTU0jjHEdDsaaIJOueBxzKqyPb2UI5TDdg177/IkkKWNM
aLUNdgKwBSulVlE2py7AEPvO9rI895V0Ks3MpQ53NXCNB49ifvGkhPoFtzYtiXjtDxBJR6cFlJ1D
LmhcITKoRNEN7J3eNWUsBsl337X3AxVP8W/wwvEwtFVvfVVM3hrqYaUaxiqIjD2EkOj99PgTkHVY
KugxYw3zcIFYJekp8BHzXC89H9QVoFfuNK29VliZmMwwEjAwCDLbcfmI42HWtg0rXPnsNrrS3Gye
04u+6fI5LsN4HLDTCTEgng9BPceFc7JkhEwHrK2GCINYaJ0HBQqT1sWcVfE0iuKyXUvcI+3tKQJ7
5qZxjOHRjmHMNL8wTbdeyRylmJp/0NfqiZD6BKYd5e8/HLeU3NNgNR/TwqZsJ2YBBwg4W+b/7nls
NqIqytPp57qR5R0kZJJX7JvQDj6pCwpz4AfeXq3Oq68VkHeAGmBkFZ8xnaNdjhY9tmdeUUhZ/FG0
2d9fywhNwgxeWY99L1k2QTrVgJ9qH9+nYJyS2+5QXI/IZkJ7V1Nz9gY2knATDyrBXQi25HGhDCxz
btOEo8R0TywToEu7H+QAHqG+c3rC/PjtJKMwAqDTgs0cZukz8eCLLpcOKirbTP+FHy+m/cAZi2E9
dm/QBrMC1AOo+69xWH4eZ7cz2KTm/yvdTuNDZTW/NelKd8VwzlS3zG6b03XgrEtAVZfMa96d4fKR
Pl9SyA2MYzJJ9EcMuMgJLBbI+k3ka/8flumKR0P8dXHfbgY1l044DlaHoGbiKXbOA8yG+4gsmK4v
UTLB7U+0bts1xseNAWI9EeDJZmaLOPeoD2A+jAJAM3ursgceM/v6rkMdC92OJ+TSFEpOaXDsl85d
cUHLa8n36VaaPwiwaCsu5Vpb95yKIB2aQu9jngIN2eBiGWHzCyhADa39M8wL/MZVP2vGHDbuzDZg
o0Fy99CXdp7nEkA1fZ4gwTh32k7wcm3Bk4KJHAuoEwdWrgPxk2Jw4KXgI0nawBGR7mBWB1IugTjt
/mmecWQJiLxfFGsqidljYwIAYfbhYDBqQ4DrHoJQ3CLQAk3qqG5Vcku6hrOLlBOslXdxojKwEoEl
tj1/UKIvo+gJfQSThJ4vo5UBSyMCRWezPnibhdsnkt8ez6jA9MRDf3E8psO1iZYcqkaHz/L8E3C4
2pk11GpQNQlk24zo3mw3QPnINEDvK46w4VNym+ChZph22bogeo61yzxQ8dM6/zDvhOr0Lo+QSQMK
xWBlsKpZJRKbjwbwEbSucrs5hErKJx5WE4MnAjCnifQMWYioCMoobGVXV+pbtYTEgtOHjGct5xLu
4u213UvI4bMJJBNh8aaPrE3GhQXuijxPELEIMF0ZYE3uqlyv3CYK1DDx7ccgp+awBFHST/93KDsD
DsfkLHOHcsFUwSNCFyiGgwxR/PNMVztmuSvQKD2T9fgIy+M+DKUfZ3oCLdIKLXwOub36NGsvfUzu
Ps5SAfXPUlBmszHqy70E0cb4N9+f6Z/oF+kE8diCByI1eVkrprKBfh25lmnv7yAFuqo6j4YTuwLn
HfWbnoCzRDmN/SAOVoi5TeE7ZF7JFv2SYp/2YxSnFVYbzMaTgNieseoJUxmV2m6phJp8rFwmuFd3
ZE2MdBp0oC6tjWpLnOS82zUogFoUI72NmpFt3V1xVxMLrXouWMuBiBQxZSoXWeFmvCSCPSyn0Q9X
W6Rg2RzsUXhmsEInFmOANQqRv1tJEC17HvmRA1l24tiH+B8OBlbeIal3Ph1Fo5Lq1x8PwEjOOHX2
60NZzUb4clThYaZOSPijwOI3Iv7rNwFEDHA/6tY22hdUW/ASRbXqLCEDVnMpO3ObI7YzX1EL8ssU
djq0cDYmvXI7MweETR9eU9zAcvUlH23/7s13d5oHUneo2jkA1VW5mj2EoXiRE45ppKY7DpKMpVKG
DVOlDiQ9m2BBV8bnPIWKTdVQMAbT0ukMAwf7BZp44uHzIhjEq1YgfUCXLgWCDtuFDQN1oxzlhdNE
6GJxIdJwvBEYZ3E6ktMPx0DcEOIMFEJpvIvs+R70AA9/SpS/bcOdBQ8wfR6UgOk4GogWhuS7XOxW
YvXyzqhhayFv0+WkWUaHO7okWmczNMGMcip+vrAfQmpZsLoJwYYTnulcSlkcCQYPPmJkWzawDhUM
GxX1QwFXIHCFo/EfXnpXO21qELnRxdOm9gfyWcb0+OKYcW7A5wv4yjvzEZKR3O/ZXDvsksHY7DBh
RMqfVonN35SjhkYCRhepvOGpqxx/WnXIiV60l7pPqrnTxdlu5RcUj7Ta7QTaQ8F4T3Po8wHzBvjB
oQ1AQ+K0dg6oHmEXyhgrwKFA5mkIAAamXdbEe0CMXL6bb8YgomsrPTlx2CtORt+Ymxqa8VNc5ISZ
fS6MqlMq3XNJhNW6zxs3Gg7/xWaT3KsaOCohOibR0rUYSX56tHdqXOZesq8XGFTXNYc14QLh3C/Z
T2HezbZQx/tYB9boK+iJApS+a1EOQuMSTcZevcDnPvG3EU51Jr/xg1DuIz3lT3l9oKQ6+VdPn/vz
uvbG5LZbOnepUOAj6vNca4AO05FM8VH/Wb6gtwQd/UK1WF7hazENAk6Goscxif/G15rhX7lmSd03
fM9X+YzyjY17jiILJp/IAUH0r9mWQbZAVVaCK63wKLPwq8HH1TfABFQykYrXTrBm4C8jYCnngHmf
ztqTYLAxvYejnjNT+CoGeal3OMdVBtwZFlQhtA72yrliR00iGk0ufAZ2t/4kjYDUiBDTwzQ0Zya8
wHzgViIHSUFAw6xojj5qQVD7HOpaqHr/PJK6nsZHI3naKme6WYtGTI8/U8lODPoWpbnrTZ7DdwuJ
X2Dr4biVthauWq9zymteQvCUYuSfkkFyfG1lAFhV/a04LEY+o83SFLbrAWhn97Bo1H/wYUjfiAzD
kKAsH+ipODIY2r9jFLConZbkXJ1vLMcu7azdGFUuAva3JLwoST5xCDT3zjpVAhznzxpLxJ84ZH9P
q4WwhpLJVn5lkxPCkEcAKdCb41S97c3fNH1YWljLBJbyJRQYe9EcBfEOiQLr+HiK/RsiseDkCrIv
mlOzyhwGE/I/LEjJDrl0a8k8EutKmbmnuQ+PfECGv1BodTw18WiNA+QcFMrHtQasXwpXO/LQAgtB
UrsUAP8KwN3XRhXu+a5SNLZo2BDO0QOiXc/xGGo+zHlK1yuIkdpW02yYTfYPqf4F0Hf+T47SU13q
pS5L+aLtiYuMEYb5WIOnZCNr1eX6xRAnEEU5jcN7pwfbTNVDTHD7QZbRiSGU9yILWN1HKuNW0DdR
VqKaMEkhUn2w9UEhDJ5XFBZtNlzbaXw6TTUahHHSvbP+vE9cHWif4wWTEaUi+vYiKrBIEDksNfZT
acO/WXJE391Ex9cYKtmtl8kWa4GcEVZdx+ldfPCqYl1H8NcgRPpDkHYw6BYMn20jBeR4+g/crWDc
rNVo+OrR6blQQnWZ1Wzs7fCi0ldjqvZUzCvfgh6gzvrsePLu8TxtKOInTWggB5lKLRBiVRw0J686
wIy7Ovs3yY8NMkdeKWd4eJUWGTbVNA0SF8mWZbQMBy9/1HpxOQHCfkChYf8MBWU1NdWMIAL3fex4
C1jH7Yr/aIcPVIux5P590+aixh+OnwqbwllA6OpxeHknOmR4JM1XaXm5qEO/y+VbVn86ZMnx0fI1
rW18nYsDmVPloqo/tZVa4qu0dGiB5oN94sFSQ0p9xb033pV07KHVjZPr7cKHzV1zyNoTcaKsxifT
MlsSYl0EAucFpkFdbRGa5VHGIylIvv7wDvSbOwsCTTCit35/pKSSBsVWWzsSLkYdGm3u8vxps1en
N4nM26vPe0oZtOSlSagJ2Gl4IkzA1BROakYVSXjok7zxyOIKQMZBvz6szfTP7u7gCeOZkjiK0U5w
GHiTK+98+2zogh1wplNPwh6nLauLxjZicXewvwloXqe6tL6Iu2DDr09Re3KIOsqXdm4Sq+z/nwWU
vcdpSHzg9lcMvvWBqOmY2DlfqjmMBgfT7xj6MwWMmqY8FeZElsu+1WLU6HwiV96xF1Bl08hh3ymm
GsuILkFb829cdSniRT4XV+jKmLem1vqyVgOwTRYEIXq6pLuijHFfxxR1Vkf5oPRMXITqgbGAEQpl
V3aqMd/dojPlG4TtW7WwDoimUB7/uQ1GcdqPsZyMDL9YlA1hCsXuZuIU9dBqNaRwqwev/qQPPkKa
CQoWI1VIIj47Hv7KKEyma6JQh+WGk6fUY0uv4qQSwvCQxTeDL86KPLPv9pDTpFREjQVRjPYVHrpO
JfX8DuS1i+vZk/tzgybDRTDiaaukZUZHxVwn6biI3tFfQUH/VR17uXmIkyn0UboJQgY9o1SNjTss
S2sjKu8vLmjZ9n7emFkwBjuRnsHxPsRRshGf5jrnsJH1eOaeVaeMJeeSPodADdmyz9zzAFToJXiQ
de5JHbkwxDDcC/7WqJZzXnP8k3tbxED9xTMFXp/JdsP3Kts1vKi3Gr+QAyStBJ2d4XgiJTm4UUzM
2FRZ0K585pLhQDnWSkKaUcQqMdzyEdZ6PrJWeoDHRmzfgSuSCF+/VM3ScnYWBsIfZn8OLajIBA5z
ogzzfe4mSgqx2cqndIvlP4NrjFirQlJQOmQUhoGHw4uzg9+S1t3HocDhirn8zoMM7kzuhKeP1e4a
KVLAqRvQRgV+CTFUo8EuEf+BAllvTlvrA3ndQGHS3QVYCC0hQzIY93zSXNnCTpr2Q+eOEHkASJ+b
pebveN1/PY24jrlbAvj/et11lUn12EsHD7uIxAB4cEysMmKZK+tX6v6samMHDXCFhwuYP7lRMFU2
cs5lltu89h05AEGLxpJ7jj9LFx8bXmxLHoVYcvW25PJsBt8Rykj3uRM28q5AUaKEXA9wsWbsMJFi
Ghae+A3MoVut03JAZ1EsZ/HYUkeH6oodtQ27YrezLW7CD5pZN7yRSCJQlwUaCM85mVE8Mv59QVWb
vehVYhOr3skB6jBMIO3T03EzVBDcAFrSoxOskA2QHnUFzhEYV9cEyiRndb+wH0sGI20/b8SRGqHk
QlKO7Y6mJTHL2xBOkWmO1PtCU2JJMqmxufTVuLT7R46424NZEqRwWawum947zlqj/xQVbe3mcknW
DWxjCUR4gLn4H6mI/LiPeME/rjkMzQL/F0fy66C8rQVrauUxFVPPsgpB/3m2a92+LtIf5Yz+J2DG
CWe5vgdjwTf9GaLMhB10gxnuJxV0HltB9vy4erh3fbK1CVifsZrZhACQq6WbiYGJ9aqIxeTX5vZR
H2AdKONJDRFdRt/JJwa4yYQr1L1OHuLtYlqp3Zc73MkQAdiOsuw5pHIQiBT0Gi2/oYqufElTeBFF
b5noRH9lpfOvJSFtrvtLsd94mUqzxbb1KYGpzQ1yX23vQ7z+dDYJSJOHiJLiTl5rv0FT1WkH2Ung
1Y4TdE+Hh3Cghjq3ne6WLAQNP23J9You1uxQ+PJCAJyP72tThqTpFhE3pY243AIt4Lqpn6zPxT0k
YddWBrCQMKiHMi4Q3MLuM4d2I/6NL8cB43Km456UZLGfztKRWmv6hPy5fpo2QDQ0RKgYUvq3D922
8bd7zozRGs2eUhF954kjeiD35pIkLHxwzQD+lwgoBrDrE/qUOR40poA+R/3n/oMEvE4cOzIN3+/I
jd5yJNEn+vs0y2MXxIaNWEKtKbSkmagkQIvAXYjKu1jKwQhoCcRyYeS9wREnJqCgKGOZePS8zmV1
dACZpGx3B51PiYTSR6bPk4A99UevpXZlhD2PVFo0h/mD0wFNMx/VaiwUAAw16wmIgHDqcQaia8gv
aO++TkDm2PpYT+qtQVDg5uiNu5PjzUGBdXVxblSF4b4XU0lGN3aCZd8EIamek6hHIWo1iTH4mmbE
SDraqok83DmI/cn6AkFBP5rTwi6lqwGqM/vPGTWCyEHOtp6MmhZWxRHqj+CjIgxNzuFmKobOFpnN
hdFlvj+XLJTWsDqmOeK6qTsUI3Nsy2mfZWm/A2doDpKveoG8gIqAiVwbmnJkCNMomBHMmWDKgMao
4z0m4M5QcVSwmvpQ1RStlgiLK0vMLiMnaulx23HtYVu7/1s03YrhYYwS4BWEfDQs+st6Qeb/B3Sx
0BDSGXB2s6kKdzFfvNXFbLPLEcsOGZB4ATmIkxiMwR7Yiz7ae5m9UtFNs+uO84WzcQsGwrInFlaO
0i1i4apYI8XBtR0xe0WioR4Z4X4GX7NIbwCdNnJUv2GNN1hjKSv6XJ+7IqvhCMw9ObmPOwgKIz9l
awdYO+TAR+YB2uubvLA9QuHO7eck0yCtQprUExyleWLMOgHH2ZAjV1xOz6+kQF+Me7GVdn+9ub5x
+hApot2LcaAtfZrJ15UKle/7xQZbXipBJl4nlsu7uZf35IYp0fUtVBXQ4Xowa1FJeuY6F15VGxgB
coMEdmMsZDfNS6xBaabMg3RcHrjMgmaFj+/mZuYH9nfQ2661BtgPrZG50b5dCINetGgGgkVoreO5
/acTwDB9/WnFhVN1bD/bNbfnoq85US1N+jsx9Lt8bm+Vmx2BnQAKM7lKVE6Ndka01BSfAb2LqXJn
kU0hBTzUJkTNHkaf+4JT9W1NMrdzS3sb5nkYK2LlEOPyXqeo/hIzbxyfeEEDp+QUtD7dP33ARBVr
WBjC0ISwsVTDlYiVcsaDHecEp5ZEfMKJm3avxesRjsBNC1/Tt+2QvOi+KCZomt8rxSIQuvRqDCAi
JpMqlrysBUT4SCIxuV027M5fmppnjgfXoCcwz6ro9Xl4nJGH4wydI9t73BTGFc63D4qEc2umDI7x
UPRHEt+qgGusbFUS/QCIXcJqZ+Aujlq/vClwQzMfS04RKlGdZyimhS98zsMtuJRMjHLGTIdxXliD
tO58YHTh6jarI+GVbIqAoI8LfnB1vyP+UYxQLm/NKNWeHsXTTVFhe1o9PIAbTiT0jTR3wS6C0g7b
cx5TO48CqUBf8bL7PKTcoxiI691UDrAKDr8cpmCKINQ0f1TNTEYNmsqtxegqxqi8RQIVtkosMzrs
YTedTWJVHqx1GU9SftrYzQkgcILVg+mBakAI6Pq6etLbzYjXgHHY2Uv3+/s1Yv2r/yKnbauOROgh
hxx2m8UxZ91wxsdBjT3tQJ2Jqj2kYi1Y2dJsQTS8CEt9mSzkeeUhKR3WZsa8bKHRZ9e3RoHKB+lu
yCZ8thlJXg1HpyZEfTK2DELU0XGbF7evGR72aqwhmwTkI8Wsj0UNVEuuAse5DepXPBWjT5TSHV+b
KyyAptJ0SLnqNv9eEhWsNbSG0eDUoXA+O460Yp/xgP8H6EBEyK4BYtLcJyLikC0uqaZgTTSq6nvJ
fImaMopCLtmS0KVIcpbkJoGHuSMEWYzQx99qm/DZOunyA67a3xpdv/az/6G9JbpJnQ7c4tbJqi43
4GtDKEUZHSeX3odMTn030dLwURZhLk6bg0qV4CHmlIZwXpTWRHxNljfLLFu0b9UkBnDGoi0TONvu
4j0uwffnmwm17tu7Xr3gNeNkXC2mmSYPORYXSwBakNqIn4cmLMXTWdMAcz+4SK07WPpB+HK0wS2N
8RiQOXGFlrKxD3f6m1KJMajmA3Yc5Iv7n+WYK7IswoYimEGOUMHoux1WERWbSdlkY3u1eWwem8Ec
qkfetSLjRjup6CAqHKML0SYD7LMmSNJcPg/ASUEuhEkgR3d9sPhp82AITFYjt0hlq2M+8NuNZ/+Q
BgsLYFNUCi1Lkf5Ao8FJ0z5GFJWheUcXoyb8vAHIX3qAsRr+05bQBtGqGMzruZqUDeNdlLtJM9GT
CbWMoy9Cea9rXOxDMj2SUS9kZuy7dIBx+Qovtzp+/gHHUI0W4nQtqteLplQIVeiG6HhRwUgPVsKt
ne4sCikbrYmGZkyXiLJkOUxXoTYLhnzdU4kprvRw/i2juL/DgACyQQXVEyR+mGdPLgdsqi4oRydd
Hkw9agWwq7G0WbnMaFAFUvq+1x30++lgrvxUipyTmRNW83DNgUjGAF9RggNbC6SOA1wGW5nUus/g
398IeEQN8gh6Nk2ZGtevTNbwbrGaJIlCxJJYJTIGfyFaiHaSfIbnGeAxTlDKeFQrA+ZVCGRlWfga
2Sez5JFHfYJtRRG1WjiO9dikqfZ8n5NYBP9Huwr4qH3vVXNWdRnVtMAbJg3wu3d5zRB1s5r/+9aK
3+uqUNgKzvU3aondrii6EQiF0Mw9aiOA5MhjoH3q2V28HetSFXJElNBMRTYTEcMhCeFakUXAzew/
jiLd64AcvBN9CDYDwmpeoQCJ/83wsTnaZbExAWT2OosGLdZjrFy1Y6VDSYuWCKNdVt3VCxLKXjs/
nspQwzJ58NEfRW5EoECan+kdGtER/PB8MpoaEtNcb8VPsFaKovMi5cwP8y+YTkbruHMl+4/fJnyz
Gz97lRKK32cu14nXX0yhh6OPqagaUNu5aLAme9191fNtZTi7lQrKndBae8C2VloofHLL2Rc8ytRm
lEKqi87CGvGffnTnPanK4uyhXRg1ukR5ND20MBPCuUFnRPzp9Y3GmJ9JmQTVl/pHYkal+qj1sdKJ
YnfPjUZBVp/7SFC5wMm6zJjU8ENKP73RneEUX3x0rkLbpShaDKocr7qKaSY7o2H8gDDpBaO2xiJl
4QUAzA8pzUh1msintJW+WTvhi73b12Laxb6j3s0wAepf1HA1WZkgZnyrzaU6HWWYc1C2bBG9I9Qu
T7fYRkTWFb7W5Y1OsgYk0MYQCRGFw+ntUNrOs8v6ptsz2nFK6sE3bckCiWI9RZClDvV4hg0BtLKA
/O13m55WDzzY86zixmU1yShZN/YMLthGIu/0HF5T3O3xPgXia1ph38wZNRW1fYTO6shFGm3XSA1t
Rnhx4cO7X11XNlNCZp3s3wcalN149WQgry5GsVvxnHc5ODTGmXo+6/vX/wI06cjmfBd/oeIbU4Bo
zSbN/PuMyVr7N/25nUb0M5SDxEzHFQ1Mz7NPSh5JTVCK77KCnqKTYmW6HAcTJcqD/ehK42KtFACT
JsrW4bOLwKj926MeEH8JKsYYl/TAOwiYl+gIHSUf9JjirsZBwU7HTE/+xV6feJfkcKQQPxwQ1USG
2c/JX3qSfYdNrW97HwfpbA7qziqPsOr9cWzrdzyobEhS5D1tBChex/AykJ3m2qcq/orOENn17nF7
Z3fTwcUvN8CZMwhw7CTkP9ZuucYZxqVCxsT29Hxt6sQhNptvbj33Y8Ghj1KHKk3bJvo8q9Gpps2+
CVavzFzsOaHh7xz5X2bVZeChMcelUu647PhR+vN1F23JNlxXoqKGL43TcCOzVURRSzGYqzsi9LZj
ctoObAo/wTrBXf9SAeG97VnZI5z8Prgu4fw0cFzF1CgRwhq2AI7cYOLUDmy0Up8pT1QdIe6ETrNC
8ndF6Luw3oob7d0PW7SRa9yxB1M6o/a6WXFyoDzaAi67a7/i6b34FypXLd2UJo9oJOlBtzwVoCYm
EO3WruIbOkfq4QYXrUIHVUGT8xLAZiFoalSfqg8sTarkiIQn/+WjjAwJOuAIiTRN+WVJfbOLvFCD
pjrtdKaWgmnqENbr969EErpE9dDDi2iQuqNJBFtlgeGNFkAzMdtmdKY0eju8+tpd4qftcpNYSx7S
dyiblaJtZnLLoSa+J3acPBDDiqoOKzdrHQRIQ3m7bgAc8ErSOHG+CuNBJP5DEhMvmrclcOvBpdL8
0em8uPfff2ufKSIraKOdkrD4WV2kdx5OrglDxTl6t497e1eCJaCjFXgFRrFO8v2LPGU6goawPi0m
DrrlFVCQwkYh+XxGKzvPfZ/BMLWrcDSgrTBenMwQQeuvSdmEDOdOTdkVR/aQ4f/wsTts7CdAUew3
VJbkzytEnMD3SLxyfwvvGOobly+IWMBtbcP/lkS3Td024RN0QLal2bp2hL59QMdyOfnAqc5WSj5z
XDnzw6YhlTTCNtphEjsdXZp+q+tazMeIxOlrPyWkGUMHK5FuIRLRFxnQ5LNaVOvdw301mGuxaC80
tBCJfnCeDcjhVkL2RDkFxoqHwGnJ8wxPBcnWNu6Lxzqsp2+fuj6DZEPbD2TkSyCMV9A8QSX2td11
BEa6m7Uowt27B3xxu8fgAS5P6u07OjyfcYnGFNeVDf4C81AoBbmnmwYruTNwl6oBzFdtCpQIroJK
d/gAy50ybvYyRa8qp72ZiyRcESlRVmvTCYsoFlbdDWePty16jvHc+w4LMUNU9b88z9ULAgeItOzN
HBGvRdepzR/V2ED5qYQNEXM3ZNgQKf8HM2xZyP/g3cvK0SX1RNb9vdG3AzWPUiCjbTasvHokaA55
nn8QNme858YqsPCVR12yvo1XFTR+sI0o1DZBMhHLiufxqlgRn9Zh6yPy7AjvWXhh5q2vS7EhTZ9n
psdtk+RdsFUHp5u+/RmLn0ThcobygVnPsECM3qdhZxZJn9XV0lXzfczMF8pjspCxNuL2/93lk06c
8WlZgrzhI56f8SlsdLoFCHh+l7LUv9vSgmaHgImA1bSbBXuCv6DuyYUm9/ZuWYyHojT6nhdXyzuy
ru1dCRQfJX1x327pFZfIjZaZmt7nz7qvXBqkq296b5j5sg6MIt599KZUqQW88MOrU4c6vXx7S30d
d0nOl+09anoHarfDpdFJjvaFnDxb5vDE+0nMXKHNLuEgfDSU4t8g/Ani06hS+k3mVMWeps9xpUxJ
xaBlq6df13IXqrOdjYD3q2KibBY0dtE/id8skQjYQ7+l7XDUVBn6mFAK+cKKJmm86CR2ZLNk+Cej
nydru84gZM7FvPyJXqybYtR8oXfSuQA4tYoAAdZnw9eWi1UQIV4Yc0b3pduPlxra6w5MG08+aYSL
VoGA0D5kFWUqkOhyq+eGumuuQRngosq1geFiwC9Zawb0BQgfLLb+sND88pU7yRMHtP6c+O9f+/ZX
kmSpoyHE3bJVEOJION4/hFIFm/YDTMeEcqRv/ueSdaFn7funmoVQtANKTLFAmCp7a71AFUU4nllv
68ewAo6BxWxeB+aEpn5ItTJ3lhFD8P0DHZcJCZgz3wm1B2xRlitc9mdoYnU6QCIO3jfoWbT62vRF
d7hi2r9hCwB/zlG29vu/NiGdjX3ad2AVX0aHLLI3OzxvqLyXNgAt4IDwhCaMR3Voihez8LNofKcM
yCX/iE0Th/ZmJU1mHYkgt7WN5d9PPrLLz70IlTI+0wkZU9am1TAppv/E/1RJr7OC+2ZEwNfZlmR7
8hxkh9tFPvKc8kg2DwGRKw6TrUsBJ84WvgjfpfEfoDhesHzVSbwrxCb9FEQTHrHRF5pxFt0TUlUN
3jQXiUUT79tHfzT5bBgFIuyMTPSQQaG1HRG79VkAjpeDdiNiXmzsk/CQp36IxsSAcTmF2I/sOTTw
vVZZgDV9I4QBE/AxfzN/LjKcXVdqEA3X1Bb39V47WVlBp8ZwcClSpsUWeye+wJhb5ouVTSrRc5cn
Ba2odZJONjgRZA0z4X+QxQPN2TJxRI6DeUs2MHRn07OE4ZfnV2p8pe/Gj9w5J30Q3zp64Nsm3K0E
VcVECDWrs+2RRErr6zQlInIDlvWRc44QCPEo1PH1EWJeIgv/sfTe/ruikZt1psdSfbKSKhcgJ0ez
eEiRyKwyr0QcIDTtOkzELvp2YcuVG+Eh7MhMr4NUNMUC/N3kqFvJHZBJM6KswuG1hBUO0+qDuiJC
QOOGgJ1IKJoWkg/ddsfycUgn6xnZxzeLGX0ekV4U7j1xdAzOjhfFaCDUUZvfn8xea8yyBuH09ZWL
G2Hglx8C4CdXvFF4SuoHP2m/N72p15RN20xCZnvevbnIeCOekKuGDK/h70MEEmEwbkqqu5Bx+u1p
XwhqejzQOLWFotKCJyxGEm+zFsibwTEEpS0ZjVOYH64GGqi5Ydb1KSOYDvFgO1OrVvyGjEssWjOK
SzPsm75Wo75hgPMBQ/4o2ktbbnMQfXgL6UIkA180fV4BUQBARxPfBAl/tDOQZt3dtbglEaEUtpTd
rmCsREXE5tgo8x74OHXE//LMFjgxLmfoE8eYRmCpsg0/mqPBHgskbJLb1EWE9fcqQW/Fw7EpSiW8
51Tn8pUvJs2ZPaiA/NGrTa6un54p1Sh7TlfcqcAW6+CYrJUJAw13pji7N+QzDWCToX0EBcMaPAru
gVz/hsSI8OZZuHuUu/+QW9EcxnmEJ8Zz0ibUlJVXG6RUrM1Jnf/rTOu2qSc2kN/d8fEFCXMRr+V0
Sd4NmHF5cXKmLgaq+wHGyzWRiyPGq8GgvySAIpm5HDw/yAwqW9tivp5u9XzbtYF7dhty80LrrnJ0
vldtWloy6Ie5ZiIk70v4EYLITdmXYqOsDbTSgOqvTEckaesPYocRLQAResIxtl6Ih/aSz7fAikHa
BqDC+bjpgu89yw7L9t1G5dw1kafl3ci0RAEcIiX5wc1nK5tT2fJ9NFR6EzR94sUxXBDIY9EFjONq
2VS9b1amp1X18pmDhEjn6PUZ6t8PRYtPeZRrW1/YNpr5wZz510zgGKrN8RpePt6ma9Yzi97RaUCQ
prfdyu66ksnnviXM8D7orzKKBmQ+vaPDNnnflJ/66HZOihwhlu6ebRW+gdn7QegBGSbe3W5Xn828
Te4Gr7szFUJBwXPPvOoDSW8Tg7VQgRvOF4+lvztoSxK6UIP1eBhsurScvMNZ/UNRN9AuTjGhOL1q
YV+KrDstdKnpXEigcP5bbVpq54xgiH2lUb70cQJH2j9oYke4pdyJ4RppDoO/3fcEBzWoLKYPx+0Z
w7WIjbqnZFID3REfcnqn1JuTTXvX4fJ71ncMxVdD4KEsz/Jq2x3j4AZc2k/L3g58/OYdYs41ZkJ3
QD0kPEa6O/J5sLNzCeTFLjwafTZY+JvJS52J/9tumuxmHnxYLQ7sS9H9dawLCgBI0QfSYlT2CrQ/
LDbPOB7mo3PPKHVR0O+hX4zvwTGoDKcCnILDo7uoSEnzvAq4yUkffoc4UJcDLpXqgMZ0NWUeMVsR
uFMQwsjROQ+5CzaLKxeGWxT2RWqr8RIsZ5c3v1t+2+IoayRQvEQYRsg7qUONlcpPZ7j/8cZDjNgg
0U7XtWjd8KGvnAyN4L1n8S8D8iB8Z80yk9t0C1q8w3oKVeu9aVlMG0OuTs0pt2hqcd5PGV8nXucY
I2ncd+eakUViZMkw2JyzOvFL4iK02NeFszH7rOs33f/tLy3cDUGM6hJD27x79MD+BMO0gzPUr+/9
+Yvy1+MVegnP5S1GrwrF1zoPJ4GduOdp0QdtJZb5/JXWgyDegcK2bl3nLx//gHLWU8nt0AM8n1DP
APzgHw6/JJFkYmucgC5vQ5WZhbrpsroKp14ej4+eRii1CUEgZVzViVQNbVl4MQAaeyzU5bYDCUjp
nGXN6R1/+8goPzvW3JhSjvkLOyaJ29PiYoHY//7n9lGUnR6W40GZ+GUmDSP7HxRdgAPJq82Ad+xG
jUzllU9sApBrQ4fTgIqdHpDKarZicLI+FNmqta9CcnaxxS0w1BgpF1blI0dsn0k1k4MEGeWWEAFh
uZg+DsOMGG+YT+M2ZneN4v6rxeFLjoK8An+55Sem7PowDvX74YabIJYjhmk0OPKN+KZSxOR+QhV8
ezDAaBPdGSh9GMVlm1CfJuzZ1pDDHGfYOaH10nqDXVuLH3mbY383J4ZekenLnvN5md0u/nfLUkio
jezs+S3mOB7W7CjgY3cIKgQraa6ipNQ3LAdYkWVQVTDj+pb91YqbkMuqDpMueCgIFh1zsIrns0yh
5m9wJuvcPzzU1Du/rfy+xLnJFCN6Ma02V76xCjJRVVqsKiwPM5NFKRWLi3+RJwhdZiPa3XMnKxIf
kOI2fYO+oO+kMDcQCRgIVrLVaLN2jmGahXw4xCVrPNMni0BPnQAtndI8SJiQ62H5RFdBST+3QlhD
ehH1i4kMTLp4dq53UplKhD3WcRA2DmY5Q3vaHoBuDnaSJXt+ovHs/oYt3YtEW+F06UXW+skjW7fg
adQ7yhCD/6VfTmt0sCS9+Rw6C0FfkKMl+pWvDHY74StF5OJZ9q3JMx54H/5JUKA8BO+jkLJiBWLI
vVRoNGKU7DkT4m71XlYBPSrknESL+LALcKznm78RnWF93S8ijVrjqXZuHRgaUWsF/yK0eC2VRIgi
PLHDkzaG+7y1izWLKSOq1Ihsp5FZ9U1vrx2k8K5TV+WEWICeLJMrSDc4V72lyhtQ4hbJSbQuU94E
rYtq8jUb/qqHcXovpvqywjSLojE2n05sP3xtLZ4C0TtRqUdakYnHjkeK5T0/AYL68Z+9BFjTBPTT
WCWGe0sBsF9DGITUg/2w+GvmpQBShfac9UaePCiVnqIrl5U9i02DsE3wGrIzCM3k0/CWn4bFYnjU
6DNXM/53fmjsJqGwFIR4cWZckvtbqedvyPAvtIJ290Ja+oIso14gcvmJlrUfIn1DIrWO5cgeBjt5
s/Sj8rfhfNTc5u3afy8eyRuXGD91S1X10UOejdQjzwrMX+NCCaUnC8L2OV0y3BvM8B7F536pkFcO
Y/fg6VMp9BTD4Rw3pOiLPUeS4kIu5R/skIipA9xZCg9q0EwW1aTmezDyFJrTlDT4OodPnk0eNIMj
dR73CTp9lomC23/08SlJU/xALVkuNE2be4RCwQcYkLvndCCJJRdz+k7aMDvg/5pfJTkvYLFBzaj6
i1Y35dI4tglMhC0QxwaLX49j6WWW0FMV3rRHac/9rOtJcGZbm7XcJJSWjF4fbDYwAlC+wNzBChZn
lwoPj2eaZUVF7XFYXaaUMCfKpokmRjDZTEbGDmCYLLc+vtaX9kuGQ/L8L0mRh1/xIWeIgddvs94h
10oiix58VUQtDa7wLYb5sT3XhTamtK1oW666eFsdavMKqbWX0ETkvODoT2BrYr//46Idgt/v14wY
W6Xt0Q3DMohO/TxtKhlTzCceDtILWQ+tr1KZ4psNQYTalK6iWv8DZPs3tlcCOHxhpvf4zixL6QLk
buS/Qr7gzP9Z+qp/vCjEpS+YGLRJyntdq9xOvlG0L5Ngw0JAUjAqMZjY1s1ZpIG9u5CF/rwI1FlQ
niCGG4W2rccD2FCVLfX+tKBmlfrZoUP8ytJIOQqBitTb+OH9BdPLk3R2ZxuWKvw5KlvSKUXzFEUv
vWgBPmBPHGs53hdAQ8lBuCxqvHcymqJEy3FSH5ohu+4TyyG2EMYeAhrkeSTg4wEQ6zcKu43hmHIk
xHEf/Xd7AYzAOLp9RrU3icE2KZsvpyKrxLmYbeGteud3zKJU0mabQP0TmDIa5TkvgQnvXZ4PtkSQ
CSIsFBtsTs9vg0eHDfsAxHHFwdN2nHb2gxvBf22nLJUvLaa5zkfv9IhhyaDTVjmdexuhx+WM626j
PKDZHYwQxVXV2dP71fif6NKHyR4l/g0tXjd01bxLeIYd7yfpJFgtJYcdh8tWkEJnTl2dyo4WyxV8
li4hN8zk5wxORgZmsm/viiI+FZzyaOgVCJ6RCB6RAFaTkG/x7fIDBW9cwlu1QFutL+T5SjgAiFj8
R3Bj7TOxZ81QKSzi/CGRVQeI1NjG7SYx/b8Cz49L6itvRDTJcQ0d66MH43RpW/CFC8gVLJWHpFiH
ME95q7m/KrwfHJCNczruT06DSx0WhWbxkYtso4zV/tNi7eSLFOGwyNK/rxjcZIEPW1w2xjHCC1KM
n2eHXhWlAV41VCnPsON2mRNcVICi/IOb/AU+kutQ3WNHogE0eNUinc5uczMh2P7dQ5XpBRIup2ju
j13CRl8/6+b7njJk3PNSXaFem992Bj9Sw7CJZ+INpYdyFWysVXmC9x08Rip1/bAzFh0qCpZccP1o
QxMVlXXcX2H73g9HlT4EvyhYCbh+opHmDGb1NKTNOgcV5l6kvO2UGCH+n+yA8zKYrKIwuKMFjdvF
lRjgX7H1INqx0Jixf4j8MpWXS4J5MWJ0m1fV0oxu4/x9Jvdr7LgqhP7+86sUJzjZ4htaScopbzIU
NacMOj816TTtWtGRMl6NNCzfPPoNAf7Q6SF8x6G2ZWQ3EwskyzrDSDU9FOxjaBgZyQRUyN8083yD
NKE60mIwBI0PNtbAIK0h3UFp1Z1beS7ddPotqGfH/V4aQ0wHJji30mpNXzcX3mzj1kVaVKtHgONb
hj2bgRdnQV2BIhaOZPGaULZa8OUrK9fmuINCh5cgQ/6KyqaHpKwpEb+pavaq1F6SdRUAcl7W6QRB
hODQSZKAHwJIHBsC2T6ei+wQOcvgvgegsnHNv1MaTOLFv8kOtY/Vvj06WTtyXhfvFUoeUXVlM5Tb
hhMRZmIohnbf4J8tm4vNVgsvFR2qlTMEm0RoAWtxhmtxQOzGe0VbIzC3bzclHot6DFVPZEKoCUhR
RW2HzAhV7+gC79qW0BIAwjzuVms3Vn+FcWVl2wzJID0B2CTlbGZp7oXVJ2j+aPDIEsHS1udEJ0/P
yIh8Dp8zit9vYnC5o1N4I3kpSi+Z2k9JTSemsFUIPVhN7XYsdNNFsxa8CFRU+ueRAupjGW6IFV5N
vtRcGSiYOkI6M9gvQ8O0Jub6B9IRd2+xLuBoz1WmDOt2JtBsO32b+62PN6xacTb2W+JidGLzi9Jf
SFjNje6G/u4z4Ns/UrfsYJIoAqJA6oGeO+tLNJOVs5QPXemU/TFscG8BP8Sh8FI2goXhNEh7Dfra
PtFBLGFUOpXFGCs97Qixl4ntCmRRbA3oR92fw29aUcDyWmfk9tz2UKM/4KG3wEy9yvicnD02+tD3
rbNZpNtUs4eW/Yis04kT+E92C7GBrSzGQ5qBaVsxKqGibz74rnnD1nWt4o6P+vaLr746pGRvJ7s1
UUEOwpXi5DtTkD7T+88PziUMtZRVnKaZAnM8RojX+V8LBOoVw6fkzJD6TxqJAuVt1xOK4E5IVwJ0
zQ9D4N12K7yNMZk8lslVYIsOr2t5M7qRz8Fmm4xe7aom00hJwpwGHIzVIWImcnI34/45+1yhOIzF
/xqxjFbXAm+yYcKe4O4S1X9UWBlxx8StErRtO8zlMNSz/Tnm1tdQKfGlnhh1YfwyaG+y/HCU0cyq
Gs5d4BrrM+8xNPbotI4sDnJudUlq76mBRC1migbSgzOGDluSEvdvC/lTPVLdgkuH6PXNyRoxD1/j
PVgv01Zya6hDqErBT+o+g7dsfxa31VawxL1boOYJjaag9rAjdb8gdS42iICWDJ31rAOjidU3CABC
sAb3/eI9JXyE9xsxFQ1Qk9piZlK9p0c3lVeJ96rmUkG7XnbiVRUmnNjJUH07h5rsNAlIJlbDhT9N
h1arAo76POpZ3iIO97QpGRGf4HPPD2iXA5DcUzU1yqATYv1yu1Ylsg0yYoPJScivyEzJoxAt1/9Y
CgbTC3G5PV8+D39p9TKPwjEuwzOmOyEdhZGXBfBmlclL4+Vd0cjJJ2HyyXv0AEclmwEl7GJ2srsl
SbpoTJpzj8pUKoe4zbCgcwznWNn2w4kz1f80W7IiVVmf0T1lbR0SbJpznA+8RqQ/RjuWHqM3t9kc
hzNl+v5joEC+5q2wkWw552DlFm+KfxNFZNmCJBAER89EZVz679IMMHpMTxY/dPgQI0UGmeAjDm0Z
FCdBiid+nxJhgW1CBoNmvNudVwVIJd6QvQfENK7Rc37DK/hVg3zVHIzDho8tmKP2nV4PNaXspOSz
EDiMUsqoi2VUECSZyvd1ELmy88Jz+GnkY3OxiMRkWMRCDFx5AVC4EqlB0S4J8i7iVdh4SM3vjTXp
HLKARX/pciKYxSySPQpQHf49j4yB08P8i98zlaUdWqK0LG4Xx1cmrbkCtP4TDBh7Rucey+cyFp4G
TnJD9eL6jhgRaloyirl5OjZordH+krBCFIfqjRzRa/klw75LwHyxbBlj5vCj2rTPhR4S2Fjq02S/
5R8ikDMw2OZN4O1dc73NhgQ7usBtwCdYbQ0nQ2SGh3ElWeQJ/0Jz5qBdQIQm4LFbQT1WvJ8h6WLz
X6uGXjSeqWnAh3rUK6exBirAmpnIwlZ3u9cGGqIxQ+7HduwbmMMdzM/i9dvY0W3zp9Vf3R4UkvKG
sQn1h3IDw6BavBvo2xAZC2B5LnAJgptdXezeNXoDR6/lflJlgnY5ONCnUKitowgonqBTwCFHMJRJ
R1wuqC/WEP0+Hs0ty2F2Wa9iXhmpbUVQea6uB/UBeG4WxnMZZwGv7UFkQkXtc0qu0bnbepqYrC2/
/sQFmOt0BH1xOnGa0EtJun0Ymm04oJUDj0eE/fPzLTq/nH7lG15FOcQoiallNGhpaFpdUR76WEjT
QF+nHq7Hl6/9dYdXlOIQPFsmgbtbelW7mzvBMaMjeEomdkcFQX4U1vOWJYH6y1hNn6cQcEOQHcT7
5gKQJeVbr26xsr0sHUP5rvHMZE6hFa6AnFDXGE7It9j/h9HUxmZW2OWyUPW4JVONlEed7HQTOOlu
KuaNh7nLnlgCzPniCoQpYgmByaO865Tb+RmSqPN3WMrq48S/qSrpqN4n8bECPkLZbLUdT0UWGZzM
5LUNdUhYhzWOLjWoF1HHZraOIVhuJFNRGxYr7wA1VxLx+2hOo4A8zVsqg2jpHyFkT10hg6U1p9Jk
OqnRpVDHZBptn6vi6Zmxbn64ehOTlk94se8j4P7mpWDaoU7Mh3GXA8jgThB9gtDIi1XR0czR1Ckm
DyWrRLZ2F6iwvqzgz05LmZc1SUc7YwGLpVn0swKpJHHdsUpkh6P1tior6xEnNF7lx4sCMwoV8xLd
yWIEGxk8MqmnSXBJyzi/mwLoo2fBtA4CbPrS70qmRPP34rRqfE8z9CfSx8GgDOiKviqqgZSSdkfj
yPlOsh7FHJiN9Tq8rV3ymanjkrMCvmy9fHoLVJ4K4EGkm9iI+siF2Yk0FEuLM1b+ap7/uDNqRiI/
Re4DGcxn5DK/l11BJvN7kuMZoPRFrN8UkSvlc8bTbN+a0Jcl/zg2bEcDWRNsPilMiEq7wv9gOovq
G0ShVb2cqb32WXO434irOs+830JoNZoqSZGmAmYLwoXfPB923LewVXhh6Rqrin3TKhWbDtaiDSHz
o58Of/2/aAHCYQqYago7ng4y9aGRZ7YS9ODjQIBQi2iU/G+qzLL++CZm64EZCcICd6a6wrHmuqZQ
87BVD81LVzFkNgA73SZ0W0llHwfPBA7+VDYuJXoZaebmIpyDxyLNK5B+0w1R1JbJ89ylmkvX2Jom
MY6McyWmMgLl7RIqCRfr3HPuPZvXQLncybXIU06+06amaqybM9u9WZQoqco5S3cIuHqifCKl7FzG
fWmXXzGKjbRXyF4kO87+4BXC+y0MOb7HrCOTU8uzugVbJlJvYQGA41x4C8QUVOWduPnlTUFZn9UY
FZrXNTw81KujXkKXM3nOJTO2KrXFFUIMvWGwwtJA+v7yJWZcWeEhIWExHTYXa/nXeMp0cjVmZQg/
ZQ/TmNQD529kUPqXjkP0SShx7qDi1HVb0xdxMCAAg0tYj0yYk2wUW3nPDbp1p8+hRGrMCHn8VPG4
VA8QKb1EAIhBPZrF/kfBwLpLHWAAjgLa7goYgDZZjr3XYfHUAbfoPmwekaXVh/hm+74AgNOzi+2E
Xf6gqScjR4RFUs/b5ZHwm6JfBlXcRfM8GeVgoQhgGSKxZX9PoIYbY6SEv1XiQKxCEWFCcnZbU6z7
SbxPxn/Wynwem7+eSo0k/0Gc3Hp3shYT6UuVw2iFetIrtoxTSrYeOCH4QhTXmZGnozKQVH8Es1bt
bRMAyBXfonLc4LTc1h/MOvs0AsCuyn7zgXUJKnfkyZxvMQErT/mLomzx7wEE3FzmJRR+EA0ni5wf
ESZK3jzQ8UfbW/qkt5YFPsytpjUp0tOiX7YxMMWsOnpCnd5C52xlBkC/DNckH2Ff7WVYBg7wRsK9
Frc08JWSzMaqEdYUICLc+shRq+eYVwCsxOoj+ZvnEii4gejwwTa34AuIQQ5SjYJMsVVuI6ikwEy8
ykftpxxaJ1qRVNPPIIARMjqtci6ky4V/y/qnMwgjQfNnKVXtd04TRZGsu4rJ3F528yE9GwJKjgm2
v1SmKJtTLsKQWBjryLVXWPKyieCG7NyGaJhuHczXIVYl2UQw+1hvsK/6eikyJLgCG6rBaNyzDXqs
EyfqXa06f52mKK9y5SrDr0HlKnSMIav2VMzOsQtFXZfFTSmZGS7xKeLoWb3kdERCtVCyd2A1Oq7S
DEVgwRGebTdv6UZEIkrra72J9w/ttKK+8cx5fPHbmBwWOl42Aq1ulAcuio0h/i2wVGhZDnypapbe
dovcLnzWIZrl7fxgIIcH2PIVeAnoeg3vQGnzCSQ/ggBNRa85qpUKO01JWtIWoIQe0d2ulozj8kP0
8dYKqQCFEzneK1hTfz8a/gq8DnwRUTli4pD0AKhF/HC9/2AcrniMfeJqDQsDEJlLAWmU7g9vlQEO
NH8rSCgrFyM1vVe3CvpZfpbfIlg1r0FIGu9d+OeWWOYx/+6PKkh+UXiCotQ/mBvIUmyXLtqo9hVW
0WYB6pzVkiFzT8sHzH7WIAaP0fSjJuma/y9pduNz9mH+myFfd7LrMQHFjgFXeEGWiBpCdSoOlCl/
a6deWNHd+KXVZv2YHsFdBtzJ1elV7RaSralLjToNfPZX2v7vhmtxw6OrPibPSEocXS6LJq09oGQs
pqjR1nEoxNpUJDLelTB8C7sEFyW4jSjaav/C3vQ8BKsmOtn9rQgTlErE9nAR6SRtA2bUg45J5qRm
ZB4lL39EeslsQODsqnFbTrwOFIzx5QQ6esaD2L0HmdaHLBrRy8wsASzt7Zu5g4cSkQ2ehgSIZUjH
Cm9RpcmrLdW/UzZsDQN1rHPP7O5nHr1h3E1Sn8lPhV8gU3z51EKJ63cd2b8DPLHrZFb63WZ/tkHh
UFiX+wFVP3qhBDazf4pWBITMi2BLFINJ7nTFaJmF2GK5MkCAbjLD0zk12BrvIkh+KeTMc6A7xSYx
pjpElkKjQTWgcNi4TWUsF6n9lPT5H+DVe8FFX2m2+KEGNA8ZChMGoQCS/XOHcBSLP2Fr+EIDH6AQ
TqCsPv7TiXwWvGBikzLCHwP5Sq+osoBtuc2idDAwXTSOhWlNgMeAXRYhmI+MfdWHMKqX5Nth8x2V
YbEVB+aVoBwllieOb6cadagUbI6IKYJn+SOPeR78ya/nxfpZk6fOTwJLljMTcLFZGbI2INqjlhhg
y0FeOicpzwi1iLjJDtYwJmQKT1VaMC0lDVIYHvcPdiHwShO7wBD9uI3JVfPqPe1bMwcEf2KejW2W
MwmNe4M2iLj/GNHo4ZVVqp3EqbR99daWNCg2RpNO3oEtFKV2QZHrefeRORv53lIViDdp0Ov3wwVi
QMvaB3IkAk7V/csNaVXEmav/AkmrgSYoDRk2fjEQwyundjlwhwKuX/wIOd6hAvxJK0uv9nkuokOE
KV0hN9IMAfVP0zn3KWKdaMQrEHlzPkbGCVvcdKTwrnhJtE5pCCXh3QMDFrv3lwut4yzMcEM5gPEe
N/ICdNqz31gWuxfnuT9eKWWpIPqFlNgFAEcSSCoOTMjHSrCHTdnbbP3iojCJYhYQQl5QnXfsPx2f
1THGG1lJ5Ga6kmKI1oCXtccenOdSFpVAQ2t26eKoZpgW5FUmuY9bK+rwwxS30UvmRLLg521+pkWH
BWGmF3Mv5yTnafvGc3qu3CD/GGsb/pC5WHz+Lps8uRW5HyeTJSB3Lqk7sIsSTMSSo9NydIsJFgNx
prEUVVqiAkNnrlwXK9Am6vEUVmNr41YdU6IdTfZMHr4FhW/iD7pyKZErG/JNV58/RZRhDcpq4I6x
emureiJt5kWyZJA0LYn8WFUVYfQWwYf6gYcM4k2OvFL9Om+KSE55z/DnXwIu35z+4Q+tNY/mPsgP
pBAtBv4F2Cc1lH0AQKxxrDfwGJSi6jfPQMT297U8h9+PNaXu+jKtD3PLK9pNkjRoUxLogvM14mS7
4fQFUhRU+tLmoe4ujLRNM8GmsQEBNQ5K6kVOQrbmZfZCDbfzw2gpto9CEukhgXbcUSpaMrCE68jh
5/pB3zvmNfNKcVXNLkmGMcFAkg8TexCOPJ2WD14NmOaVVBPolhUxC+SDx5VI8l9UsgplJuCueQQI
Q6Q8DVAXVT2AHgz1+TgWM7d2AvRxIF/r1y5ZNqm7eVMS0+2UNBUy5TWQKwV2I9dBAOBE8AMK9zpQ
heIu84HJqJsJPwXOTNIwZSh7f+dGeqqfHzx6OjhXO3MMOOSayNgkbciuCuzDV27IzReGQ2IRbst4
CtECNHGmolZLQfobIxVK41gGcNXBT0xN3k05AtUYN4qoMA7hOR4Yrj1nRjf5MY1nIUX4WHInpGQy
UwCWr2H9xgsO4R98Ekaz4mEoAT4UVg2N9azarst8qiqu1CxeilJlXPcNi7uJZtunNdqOtMYMY6Jy
c8KokU9Pu8DdIJo+mUzV7zLZdD/7RY5NV6/EIYqGpyqJtnc+Afhc388nuboV6X+9R3ZYFGnd2spp
QT2D2q1557ihNiE8+q2p3c2IYfv15rj3Sk9qLaTfdIoi+G/oylpKtiEulN8Cqx46wuEv+7OmMB9G
TVF0Z6be3/dq7mx+EN0LYdOzzgSyxN8lmrGSGV+bo9M6+Y/QwsL44/i+JQHFEbgY0qYEl1orLLS9
XsgGuZhl1vo21D7lEpNgHIY9eeqEMdoxwhGwN/OCBmcn/I0Rxfm6wEu88Uepy07GaYDHPfEpLbp7
fAY+OXAEFZufsAoUCaoHRp9KwCg36G3RSi9Hzl6hjBgCcz8LzXV738pHQdLVE5GmB13v/0oaKMnT
B1oD05vunkjZbOZ7iFqXcV5xioZR0TPXtByHmhVm1sEGu6D08XhAyO/oby9ov9aQNwovr/YcduqV
CiBu4MRTVtScFLLlhzeFb7pAKkD5qvEuAwtd7kSQcxZN4nlOHrD0YA3eVbjIJSEhUyPdCE9H4ekp
h23lhVAyfPLcRke+0C+WohGlxnPYJIx61LB0WuYofekDTUuiU5UKw1RRruknDnH1iv6BO2DFSXqu
pdICLUIghAahNTfu2H4SYVR6uvs4CQ77GuIKr0SFiAf7SymDykbxxf/qEpIy8P5C1YUdhNzDyPRh
uUzAGt0uwWjp2vIttCqoxJKxwGM4IIRsNwZPdSzwSGxlzfQfQgeSxK1tOSX5EHnOeorGhaW5ONjH
uI5n593Z9saud3ED1bVRGjIANlPTX0ezMTG8Je4zdvZRWdkJUhkLbnODZzVXRDwp1+jDVzDJApMQ
6xk7R51BIplhKXJ9Mh9JoiN+UQAgD8gR7Q9SvBxgapqf+nQqffXafL4rNA0WJiFI6eUllzAOXSfY
1pEgNS9RckedffTVL7VCbzScyVDQwzOL4lFnIbo+AkK31HCzJlu8SQtWXB3s5Nmn0P2wUA9MzhuZ
UWXy0XyEOnd6LHjGEGaD4SGUQkR8VlhrzwJgxnbMPJ9SLnPXKx9sXfRlPcx3cgDyS2bJhg654lj+
W11A6leGdVxjnBRiTXjPuydIRiuHoin0GIm606r/kMJswVrQq93MrVT0y4RwL5foHOsuOBITZ4Zs
ksiCpVrAD9zoB+hXVPagazWkrwr0ioiOXRloYnC54ZeNBu9IvQ4LGL/IH3MW6DjCt33EHsDvfPVn
bumYi6uRsNFPIEJSlGY7Iqcf840ocL2qfRiiRJcDsNERisdSB57maQq4ZQkVqNHp1q5uk5TdXMJj
pG2xW808YdNVrW0LxUaWmyy0wyt8CyMpYcISFW85Rn7xO4Q5uyOhyLIjO84j38EaAnb7vMb00H3V
YyNoCOZAg5qieSVnlpdmxx4Al0xY50WkPaEw8XD2gikG6Oy4phmau6TJIaP8xTXmvobiRMP72/iL
mLePSDvbZ8yv78M0X/tpv1fi93EUkE24+yA6ZoqUJiegN4d9DFk6St3s/rJh8v4HfxYLk6sOfquf
7NNzHC/hESL8PUKBjOHaWIcQdvDG5BM5Tb0oszQSvbihe69kyWH3lciw16E//NvOeTV7xxnBB/nm
iEICoKUGUs73iNdvHKGI4XC6AfDBvqC3C3Wz844k9z1gOL418xXKdwwIg9IxfnPJdIL9PEeE2P6V
Hla3IpjbY9QxC7CzLrfGnKNggPBz5eFH8ylFrDqtt+HyGz7pXyuv+bOXEloYHkKCU50zMAzl4kDb
E4ZNwsxro9hIwkqVm06TzdqcCZj++qi1UY2Cqxh4ulOo6YVY5DYslCVuJnb3O7JFK/BIkDpf4dci
INYRd1skj/VkpXysGZNRbLiVskECMNaymPWfaDuaeLm/zMvMYagSimXdIH6VKslNj00p+fieON6E
eUNCGeuDRhaxxiQTzwB+1VEUX95TmYFj5aIZPuqkyKCtHwrAJC30Es9YGFjqbSOcmMRP7BIB1HQq
ixOoabAphQGEy/Kjfos/NgQRWJuUwOmUTwqwUg4QCLXXysbhRUholQSAyRKiWAjTEcN3uBMU0AmT
kH/bHXuVO0iXOBSJIziwNpHYlYOukr8YXhMbg5zzBc8lzGXewLpS/ph7UyK7JxuURELhgjCOkZot
2+tuFbgGU+0VbUdIQ34B68n9nvoJvpMzXJISrVXvAzrcJkgfiRpQyLLmMDNF7P1LV4o0FEIMyiHl
bMANma3l6EcEpfoV6opSurf4YyhciRrKbiubI1WmP8KjoudLY1jgMEG+gDFH1OO19w7vdbcFdn9I
+cKfaQ/bpmdxLXr/5FZZGxLjNBi6+xF+/pAsD5aKw4Gkxu1+JPO3tQclCATzWsfh5c5U9xtV1Df9
UcUZQWa3+9Vwhi5/RTg4iPMRAAhGLJxQENui3Y//aRO8Fwjrv+/EXj0/Uxf76WoVI0qNOQryZ7ai
CX9tNmOlBwHNHwCKKyinjHBsYD7rdt32THWJvRnGNIyGD6bQa33U/TpMrRarCV3pwbu+qz7XTu11
QzOSwcYf7lgJnnseEg5k7wTZ+OQz0xU8wnIgvk2cbvPgGSoQaTQk2+msGEuJZIxurWlmqePkp7TZ
rcECvxkvgsS0Vy9nb6hnVjcTCP0WaZuLqH+vVmiHeba7IpL7KWT8Sknj8zz+bZKv59dq3jxoJb4g
Qjrynahx5zjF+CcT8JiJ/jt5UB2bnNRzZI8JmCVmQVOnne3EmjuA87e0GSh07v+oJukVIx/kjPjz
Hco2yZKQXz2Erdnh4r8lMjLFF7nXgWENc0LqJsZtVVuBG3744Ra1/kEHaZiJXZHUzKvG7VoLhOOd
71ieXvgDHi2DfTe89IifDVNd1giEXRQnLDdlxq3xEd2ae2ssVgVt58wFWBiSjxi4PBaJzQedhOnp
tkuVcscclo0Rvg/dJURsVl82vW2n7a6OOK0iqbU7dn0U0SdtAx7rqel8EcaHZo2ucCNi8Je9ERQe
DUqJeek3v4wkf88tXOAE5/tYhuxDOzxsSZ0V9rXdHMkK/n4ruljlWlOt7ww8/+7Z6ylX0KhTxe/P
MXsgNwpughVdeGcWdLqr4Cm/hrK4xoXmjny2z4TbyZVBo5B6oeF8tW4sxrGEnEXVGQrnHVIEjSsO
xLq1IYEdUJZ9LDASjLK2PqIHEucAj2S4/HTIPJeMDwmg/6QuoQAW6izpdc5NHhFPaA5YlG63qRre
4I9phzUeBE0xuUsq7UCtIsnj1piiV9u0HKMiG0jJKy6yKJSpoGuM775Rv57Ig3+sK5o0tY3q2rbK
DF7tfIblEoo0OWijFwpJquqgvM1i5Qd/1g0zasWmKFglzik8S6Pjs8FnHYUa7irEdJ/eN3sbVvYE
aX+575Ds5D4StB97TqsG9t0hNTqD8qnoMk4aTClqAKqhC/H3+88tHMYYn5MgkFCuadUfrLLzwNN/
iXN+c2qGy5hqffLgIS8Hd9ARSaxi1hqU9olbLBjbfwnyfLs9XLy8aOWDlEu9sKTRc7lYkEn5PXGz
BTdVfdAaNyyil1NUHPYFjLdyN21PfcUbOXMnIo5efLaXxSGmX5i61hY0Vg3RsPy/RZoRJaNvbkRK
OYf9p2H1aLCmykwsDuB4E9RqadDUzp3/mwtEOAZYwzKOsP/IUgnkeBcRYiM0mILizMpEg2/S8F+Z
aLEcDtBoIHh9JaL3UUDFSAAm3gbcFQ3SXTNc9AEOPVv5cNe1Qt2F5C/Vc7NWcJWbtQEb0J7iofvM
tmgW9NqOAh49T9gEM5+iJ9JiyvDt7z5VHqHUdK6gAdkpDsAUAiBvqLhOhPMrOX1P3PBBWrdbOF+G
F0BV+ksKe6H4enGVjrQIbkBYqyQegJ41kNB+KaaB6EXs3snIZNslrgX66h1KDx+XQjFOhelfcYqy
HPSWB3GpaIHDJcvUBvZfSfZvrxWsPyY27EpB97JA0WSaEtaeFNvKZmp/uhKMDNGzymqt9W+qxzsA
QC5Pv3MY0q/IKRaKZ2/BArPo9H5XsF2ZZ2Q6p83KkqKDfoppdCB5Wu7j421SJkMwr78l5QTyIas3
7FdHs5kJEV6JzoeS1eQMt4Y4tnDFChh525ZO+sYrqK+uQG9kjo2/eqqpL4Nb1cnM47H85d5c0KgN
qKw5PPbPxd4APnHQ1OGLpk850TNwtqfiQ4MA772ju01D52dJCmkLGsYtjMcSrgJ8abFoXBuX7bha
iJtSumF4uO5ad/B7qTOUypsJu58yVDZM+ZaqQUdKRJYcXr0az5AeC7233PIF0p1xevIIFV2Bf16z
x/vnD+71mcTcJ1nDpe6Mt88nDChCPeA4swSlmHZBLCvPMcli4d1pzCSaigGmW8m5FATsEaBsGHsC
Iw308TBiFv406avSTFUapw8b6DqwZ95LgIW1lHex0PYqJTx/ersZFNE7XCMHEBmLzaPfItfDxqkR
Xy74prsbkhjYuY6Rp0baL0OSEabZFNla3o9AcvRWEhFtny9+UqwJBmn4wYwadDoE10c3iJAQLR+a
UQpTM6c8gU12E+9bU0cFS7deFVuTinZZ0o+ANRo2F6jcK3D3auZAtYSurDetGD0uU6qRmGw9t003
NTlBbQKbhMiSD4nK6k0DY6fi3ihDT3NUPOLG760rqb23jIaMxPWA6FwjZcML50u2MRqREFtsa65S
9G9X7BdtgdlUsN/WlRCjYAwroQ5w49/NrGg+GPnMyFskaGxfDqaW2NLuZnYANZnkGNxMhIGEgsQo
zMkcI9aabvEOuTJMcY69YmMNQQ8a4Yi+kJHtwFHzmcLb3zWsS140uzwKS9K0DxxjqjK9/LRGcSsh
DbUI7VeRf3VLVooWhjmLu23MeZBnYycdULpR70pmpyZlQA+LmxjcjolIPrKYig6tJeGMe75m0BLV
jqgnuVHuTFdhSbskQDIxDVxFGUMEFGlcrVI8FDyx/z0Pju++aJSs03mzJTes59QHribwGOodQuGW
A9emCMtxlkhwMYqQOlRqaBVhfkHneUUwk/yYZAH9xQXatNuh2I29Qzbg8kDTgBSZYbFAsfpMrpvb
jubxblPiIUIDOhIqJe2AEW2JJ8pea9uKnqPJmbECSrUOJNDGP3IT5rq7GbXw7FFW/07+ezPAbjZ3
uVG6Fe+ulCa/XEgB2cGoy3ZgOiDjeB4bUPok9QWmahXK+u716gtj8kYp0protxWdovgQpKwA6qSH
9ptTz+kUWz7Eytd+dJvwN0O+IAZLRHrnMc8ViOz7o9CSXqXfIvx6BW0qDXIzqnnDlwq+nXOx4H8U
X9lr5imqtGcNH/kxXnsPOc4yZWFl28ga1ztrWOglH19D4BWAAow1s6ftpDmlKepo8/DEbNpUeRSD
6eunLzAMPu9CiXaa/1/0dvNVtLvm7mjxYahx55YmJpQ6rkjsqi/ut/CbhDh9y8ul0gCzh1oJTS07
qunbKW0QsuZ1m0Sc77eCeWYu633cY7mM3Xkc3p7OtvbZgNmQGZiYJ60mfdZkO/mbYLv+SVUrfCLk
xgNSRoJR+AUMscezMqRyb1/hPOUBBHfNUejqnUSI+y4fWCEKqcUc5IeQbFRkQ2jQOu/Su7u6WFse
enuXMoPY2fa8Co4YIzu6exz4Wp+R+SKJur8Ag4oNPvSLNoH30ddxC73sCSyx/4NltpvjaZVn0ldM
Q3Z/vrOScb5S2RiilF4xxlyfNUWN+ZjmCpO8/UV05bUpQDE+pJjOVkW5/1j9Uc+WlvmDHf8WyK5F
52IX3icTgXvNvIcXjEIDUkSOKkHPWEcZxmXQDaauvmeATeAa1cOf33UTE54ymAMlpJ7Edpa7oa2m
h0/7KnQfKXCPM3FQzccXe4+K0eCbmiE4XMnov7PckGh5DVTFm8XmCePeIRcMhMhHk5R4aoPl5AxQ
nFRaAMKJ2gKgmITPm1nlTZ9mGCnIE9EaYq5Lv/bBwt5wboAxWvdosSrN4WAuPGb8+Lyo3mTl9uoX
ekyiy97SPZcuBDTeJgELzYsTH+Z6Q5miFw/0hl1U18ZTgoApWp9kwdSJDlbTJGrlRr3T0cWUkzME
vy0Nlrhdhobxuzuy6C9Zr9CZUIjCD+Me0wOD0+OkjnC1XUJqnaASSv4OEkb0y7pP2ebpSiOY1EoW
MMXqW4j9QynTN1k250TVl85mKeG909SjgS1i66qbmrfN/UaqfGGJR+qEPeizZow0yqM486SfO2qc
ETHIdMUqob9ngII4lRyirzU4VTIADulY/RiYyKjfAkOQgY6uyfUu5KJ9gtEF8dlKublEhl2VeSHO
2oLxIN7QVrEydKl7GP2Ubj+5MJN2VXk+rFpCVU5Q4QJHLV8dgXKuvqigpo/k9L6z/9R2vxTNHaNq
MwOa1l2QBu89m44Fj5JMsoA+K2Mh+cm/4zVALs/mEAd3Y3cAowwlx1xPLpU/GrE7gVVIJ0NmprJs
Hk6NUzClmmMnGYAk5QSI4yS2MLMQb4IvqYp/2Hdw/+cbSTJnkJs08KjblxN9Tpv2u5wI/NI0AdMo
Drv59KHGEXMERUW4iJPPjgPbNk6C3aHVFPbHcjvCkkdATCp3GWumXF2RG3WtUVMAbwXfRXYFIG9y
zMhn23v3khoi1FQPlG1L2ge3NiogaM9Jezi3/x/hobT6oy5B3r2uJICKRY05u8wYpm0UlbkWcyoa
kQD0MwaOjM85aawpR6s79ipEdkGE4ziUs+xjgJAo0cYBCJ8CS4aANTOXT8fP8EgrP8ptre4NZ2BU
CqU80s8+/6RO+gVBMO7AgUyUjP/gYjxAwPLLa1PGsJWjzbNJN0qUgGLngFRq3drDBn0B2UH7bb5u
kwEGin+oUkQFIfJ+ssk2yZSljo7JgF7vyt7urXgrUX3qbGRHhalf8AufR2zOcRhcl6AjSZbhtu8h
J/fNJniT7dXV3cXdpklfvOe3VKkGUqVL0idikjTz13xPB+y/dYjJzL/nbQLWKzd8G7CweymU6atn
NlDUg6ALxP5uPufESfloTfyc6Nuw5Kfbdu8mGWnPvTpXQ1+0akye0nLPUDenwr/4nV6PImCN0mpW
5U6SIada/Pa18vZpdKA/v/GLWVn6E2l2paROOirc+ExgsmJ9wewbMdehJHQ2K+iLBWca68SwET4D
u5VoN6oDbFwxceL1GX1wp/MM+0teN9sMMeleXhEAk1cvsHtTGVxKKAnvOpEo5Y9dKzRlvM0LyJ1u
Hz3SqBNph2zPZgPSD7ssPfRWXRDL3xOiZIQzprv+h+z9tCreUsh+tX6uNKdgS+vT55AdVaDDZG4H
MOpQ75/IAbFrLZE17wC73TQaRi6pCf/xWFEtdJdj6PmDMa6Dteewuxj+wXNP7Ai2Ouaelz8NHHRG
YFpRZIu2Ny5HYGUIutmkQBdreYRsY0eVa7XZOrUZm7oiosLWG7QQJsAjJF2JEb0QwuNdmZSKRVSM
vmIKbwCM5IkwEj1UqlIgxNtW31EEWJiwylfkbDn8HYWHyXc6x25Y0PICNUoaNSXD7c4k2jWuuBtP
xjkYpprp9OIBNEKmj1PNlYpA1Rz+e/gw1Wvcb+A/xKneXvkuRrckWz8RXrAmvq1ib2aHAzLhIfKl
4LLvVXnzelop/BbjQvG1VxyPFYi97aWILEAlVbinn7x5aysUowW+MD8vnFtfXjs4C0oyEyA4yNmM
yU6tWHF2D1XuFQ3HrQXCB9X7lQ9+LQw0g+c5KvXXMiIxZ4nxZVrED8V1lGcGH7Haj7FaQZEGTsK+
rkWfTrM8S+8XrnyGvNhyvuTezXDNOVksxFnuai6siysPv58HrnR95FCf5Ri1pqIgqyeMLflMpf88
uwpBsXtPzvbHvb+ELG7Zg+zit6JpfgXSYN01MsuojzlRyI9wgB8qd9RInUB1wJdQEECHSdFuo0jc
Lhue/Y4WN1ItLngITWxLaQkXId8CdYhbndgiZ1dwKFmBGUeVJbpxcbhkOoNGcWaYpLyHxh8RznqK
Fj6aCUpC9Qz6291Xs2mjQ/LLedDtRjyaM6v6MjiUlZGrS8xtGIox4CW7OgQ1kh57NJl0AlKrtQDq
QSF8Zs0HL/o9JEugdz/JbU1T45RPiWUCPw7JVmIgC7hraJp58ZpZWVeRjvzGpemhCoJn1sD/PH/G
TSfgGxNbfiPbg/P4lY2QRw9zi9ouNWiltA02LstsSfOSAu0D9XErFZvnB/mI+NGvGnSbtrY1uKNg
+2vfSI+TVKZQiwb6yJ8hc11SpvHSlQ5tA5kxs9dP0qJ+Y8deeJb793N8xCjj4WeQIVB2nmAcOf32
D6kkG+PyVUvBModiQ7nDmvum2b/TNpPWoVLwMfEJBV93MynCOVEVGGGD9OFbhhJQRpD7Ko6RM/MG
VIpcE+TX11YjszcCafjDAKxA4F3rO8va31rmiu87Yxk+h3HGO6z3diES46vNSw6DQnE9q6mbUi0p
xslc413BQoNzKIKGfUHMuU7zuCn00DcnhBElf0EWPuFgi22krtthTAQA4BUooQaMWYR9BgSHt07Z
w1QYN8VXqjuaDK+E3b+1QAe3D8DjtNYj6USIfKsqwseNwnZaqixxyOJMCu8xS77HKjMW2vEvU+PH
z6VNqEfR/CQO4Y5pd6sU5ubNWylfQ1mP/0NIMwociT8Cwqa8rl/hD7xd9ZVws+nlWqiAMtdWtWI/
8zycGM46zugEJcIGb4m/SojxXx7VMNZ9YLt8rYsHsiYyXF6ztzdI/0VU0zZe07E0AJqc6b+9er9a
twN1v0jTwoz3f1AiYP9a/DO5aFbVhNWaJKlOiemZ+W/T7HZHms1ygeVICiijYXyqfS62nEIkqwP3
X2Ve7bQKECWGyw2L5Bd/uGK1BQcOVAM7IXryg3iCO9zZLmMbw38o6SdUIBKiTE1Ya3dqrj6iaJHf
1aICMA7pSylM8/4K+CCGqCIFxZQcrJdchzRHfr/iL227pLt0qrxKcT9EgEZq1GjF9qDwUrGxypC+
HFQ2mqeZL923bkUK2B1DBoFbLgzKJigUWga8liBjtmcLVn/N0rG26rJrIkkF5sonCcn8iP1PBr+t
Gjb2fxaKiswGP1cH1zMMu6CIvTK3H4zrD4+xvb17SMr8I3oNqykqNHUKBQ+c6sySz57fMoEDbosQ
ngHaktnbPmRHIpz1Eagszyno3YF5mv2tjjeDbh0lJeTvj7EqdYi9QVMRuuuJ0+YZB5FHcjrTkwPL
fza3W/rHpwuv2MHHR02hWiQQZK0VjxCPbAGg8nu9I4+DkG83/wfFkmjyPxRA3emuyDoktl5mSxp5
COpu/E8ohhOpRpXM5Rv40XcAxMIx90VhmFOAbzp+Us0AgDmLe9SYp42qf/QpKuSfIeygOaFkp12x
zbAe/ld1K1hAn6tmqOilDcKg2AWxm2vfO4LmeVqUAlaCJot8Y7RSmzeM8HyJx0KFAE8HbSq0jSwv
1cSAi4SN0q092ITha2hmltSoriOZKyNFwZITzEcUhswpFL0KX8kfEXJVbt510ANI7Y6fxEe9zmja
B6dqkUJlFYTMTfRG54ixxuehSn0FAdWKdIInQi7RZNSWiDlUSCYTczO18iN11hvNifyj5bJY6YAj
f1tD3FKL0QzybpZ5FVetoYCG+Or88vM5lX5drpCLiUfAzJBWU9mdGZQGmm5lkKPDx1rqYyJkRh35
Z+/Gn+Mkh0sTjFwUD0sqdGGV37d1u9WiX0KoleiRRpSd5Bq9NKn6NbOkpqZ8PTzhPgtzTF1Ir9gb
GC1vNkVXXVjXwXhv9TntaWLOS7Esj2Viay1JU+q9ALcNopIvffWFUl8JSJzx+5yfb6emhqaFIBhh
YHD0SO89BaHI5d6dE8xribpmHCUpfTd7+QZ2cjABLWrBT04BqSE0NCOn8FXI5T3+pKwLliSHIqsa
NK+THQiMKn+hGoShRr/iXkYJcKRmPX2D3Dlysr2z0+ncn+W9unHX80yjCaCf/EpJ+4ipMKdDmAOP
VB1GlN/uvsgY1PRhzFLVfmhQNR+WA0n33RhQTsCqpl/HZUXButbz4kDUVFhXGNfm5bVGHbMuoaXa
C+8kQfjjQGMLE9mAs+SNSm+BtVbvkg5oESvBx5XRHIxuXYdYLPwj7OjxhcJLsMZFpYKyfIZ0A7a3
GdGBPDWyCC2fFvr16pq9WRQpsFP/GNVae0+3+cJSNfIZ3RTEwUvAPLbq/h5BVT5nrbk/kgLpW9/6
H3XVIeJeSWgFjuDXsVTf2JnOuyFdxg/kYEt85ZsBERpnkRA+VwZI4grJhIMfOMmJ8dsWFnRBQxtB
eEPZyHCH4EW6pb0gMXI7BpmlgjMFo6zwH6WS3lRC2//MsTrJUTd/S6VeYt2qsTIMAvuVENopTFe+
U+8XbS8L4B9kkAoSQKeW146Aa4xf/MPvwuNd+qONn3azvv6rOgnyZdDRwhVrqrglQmNGAwl9/bpF
rvlJIG0e2pqbrRsaEfV/r8pbQVodwUOPucNHCCKoYtlNx0OEHysJk3mE8XmZS7wpQL9io+6K0dIN
pna+GdzF4XyqGEwG6aLoUU95W20+8PrEMkSw6tI1yUgEZOsxXcLkSBBC3llFngBEvWIa9J89xT6Q
MMRrP3EQ5hMG5cPs6Rk/542y5SjVzhMFUlIJs27RDRzX+UWZctIVuZcEE/iMWoNRRUjOlZmzbb5U
rYWT6vfJ2v1UX7P+RvbQEncB6y3yuKH19Poaxh94oWeCMnvNi/klib8gKCyPfAS+w+exD2NOj54I
e2h3DWq9c0v3FMRXfjMn3deEXsjhY2xT5I3/wpvd4Dbf+C/fTduLjazFw4SbzokbmPyqBkHZMS0k
bBoRWpfYEKpdeeMHPqBZLztPauHUBRx3HXLDr5vrvD5bvi2oj5NtA3IE+mx3h8WJio5FeqcvLpNS
dZ8Ps8QI0fZE8+3Rzhny9hk+BK//Mgf47hIy1BDKpq1qdXc+0ec062wMHwdNCg9S0VM1Fy/O44/2
ucMQPK3A58Z5xcNT61dZoqgCPTKFaDl0DwFJIqWbsB6+8FRsHV3U/4wxuqj/eCqLMtfFXbcH+v6z
8dfRna/vVYSd3fQDhRmron+rAvxg4EUiEGpyp2uG6dE+WcDWsjKH34EidlxW3inBgtTBnrkBuZwo
z0lPDP9RXJKgGOxms8jErm/S3E4IzEXDoWrxbM/jCCrGLypMQsAsMx6w0NH9HrvCEqp0RuwTnAcM
6hW2SLOgcXYp7y+Rs4zlfZW3WIRduIhMvtvoAW7Tb284NaLNUprWh2zrx92NGi15+nRWy2DSLPTq
Qnpfvm9H0ROH0JW5iVi71gwsNpoqL9jRe5oxYrIpPCFEHidyRpjjVjxPSvDv9EgFpC83QqVzddCT
ha/c7UmNs/Nzk+GJ5vpIo+VxERm0tb5TpvZ4XdQRM7/udMsv6oPmVN09ouPx1WzyPA/ZymhXqZME
usn1pF0/pivJcafnhLXSrzFMXURkpzl4VsNTDgDbD0E9BZBo2a9nj14YwsEy63OpdfhF1Xyrcd6x
fILi1TMIE8s3WDYAZ2SR4bVQAVohdxMAyBc7wYk8xI0XldeXvofV6NQhYC/jEx3WnkOJi2z6qaDO
2tbWXWkO9qQe6hID4PehZ9s/uCGMkgVkNYaggz21yuS3cVhBMJwpueAdllKfJ9ZfvNa8El+ClKkS
3f5OUEJpwbVWY9hduLm4KrlxV+iY2vUUE+h1WwO+jyKHIUNJaGAq2lpztcghEP30DrWVUNlg0Uup
VLpBuAxgi5GudhQS9AYTEjCkCKZeOSHRnA97UJQGMwhkZOlUv+Hv6quVPB1AFf4ncwNDSYBmRLCb
5+ujVabFwRhGoQhH6HkuroFhvGMoAUGJ4tLG4uoA95Vx3to3b5YyFFaCScxbRgGaWsBBMo3QarN5
ItoyOE9WTm5WhGlpQoLBb5/qFezUUEoyBAolcgVBQCXzVjwspSWcjOma8U+nPeB0ljyLUZI8tama
8sab8EZZicvOdsg0VRm/sHb52CqFMJ36EH+Fp9OUm6oyxY0dKonQuiN9/b73ZgMNKDtxSNaU1tcA
c2RUxgiuNQF1bFiaXqaxAWX9ftPpx5BNDPq6Q1w722IVOy1G/ChYnt9ypyTlubX2I9N0mYQmWymd
6bcw6acJAwvOj6yd5du5J5QOnDg/FHnF4/omhgetX6tAawPpSl9lF5AdU/xVv1zddEBqLnStavsn
WtR0xIms/bF1IrHnUJz6/ZJSmARACxANk63t0onSq+UULHNLf9sTAA80XaVKu6wR3CUmitOxMDrh
rIZBXY/rzXYKzW53tM+jKFh367Xtgo5fi8Ww7aSWxFrnT8OKnltsMTwsRJGeKxm17gdDl+mbgS5Y
HPLeoIY7UilOZwXlh521Oi4GpbvPgJRy/kQ/UPxsSzQxiQFY4TOe3pTyKAUQyQleqaTbzJ/n2i4l
x9OWI2zTgZrX4zvuZ/XIzydRRNSSs2oxRz4k272ryoampJDdEfCwZT5cp3DkQK2B9LSwszf/xv/n
xClQXa13zhPkYV7C/mq7I+zwSDa5tvxCphPU6Zb87HdIpDaoSjxgxrbxjTxNiN+c8/d9Eow5XLxl
r5VTsVCefs/+6NLxTw3wLZbPBvF8mDvWLaVOSVPRa4TmrYwXC7LLm+pcMEHxfGY0Aj++B0oCjH6f
cpuUNP/ciInQnYCbb3s4EyflP+LpDldG6tE0YMzlr1M9IbHcFzQRrURXAqJFc6SPQK2yQoDLWV0c
WOqKOEK887sMfEPKGJ4qxFRSFAYu9ldiY/CBMlSmNTnY/R8eT+Xn37j0woChtLuSbDcECVR7LZJu
CHbLtNuJXKZHHNDxTZL2fehhuTTkzPW5HNKAywGyR23lCp1SgZCF7FlCv++Y4hh67t311165BDOf
Q1xVaGi9WnHOUWi+M/3+L7gq72DlKnZr4arzi0coUVhA7X+F20Ta/IHrIt1wXiP0v5AJfE4MDo2y
y717mjqO6jUVd7/5Fa/ZrpA7wHTFc5WkJlTnfBXtd/zZxRx7NG4O8nXoqxn5c8j1HclOfQkK26ym
e+67bDB+kJmm0AOsdKByw1tX2cCLmd52vQq9BiaZp+Daru4ilguxFmnL1/Bed/MqEymLU3GstkxW
bdJ08a0GfLe+qqinM5SwLLtQihUAvs9q9Bvbbo0BSj4yIhAwILtKUULDRkgW3a9KoKU50tVFnkuU
Ejpt/Dhzgo6qmtWp9efVRwnJVFHfYkmwbG4NBCSaSgGVJCWIx3FUB2ejzLgs/kknmjeOQn9MR0F4
5+LX5UbOiCx1puguMx8MT0De9efkdemh0bwAWwornPUW+sCocTfmnCIGm9xfDJwasXqxSzPlpqRU
pyWm+c7RNZ68CqJVkwNxY7SbDj9+yaNGbDOWOWnAo0F1rmOz/lfHDgRtO2h3y7KU7i/SaapQ0DWL
GrD7Z6BVWoJFYy2a2MkjqI+Bd4ie2BGdSihOcGizVVbTfea9+C2BvlkUCPBZsJSm77NOI7V/DT5Z
yE3CJPi+lSNibOxFybqU8USH7qPY8JdPT5rpYhp6lkaauh8cyYes/w1jRNzywFnwQy5lpLXDFzfm
DkLRfom9lJ5EyazdzkUH87n/GcMr2gHCIfcVaLTu7dkGkAkQ5MlWrONtBwiQ0aUujODIawvjI3xt
BXTpEADDAwNs+rH8luOdimG3aZu4JWeJCQMH6bhyYiIzUyg0XNJ8I48F39GuZyqsL8oWodAyvL2f
9vf6AYhPmJiqTbLSrmVNcSd5x/q2Qtjhoq9KQWX2LBmg3Ne1pi07eD/x79cCKxU5ZeSeKjiVQxcH
La5XjDUf8nh8wTLP4sSoWO4/dtbTGCybYL37vhXPq8sW4hkCXWvDZtDReWW9WUMiTzE2drK05eez
8PohV6tX1ysK8qpufXYJIe9QZ7h4dmrrBoLtS6M2WsrU0ubbfVhAtHJtpvl8QtZ1SHcYWfIPSdUK
uX3QNB2y8ctuh5kq+D568+dLF3n4GEmAtbe7+8W5aaFqRMS6coBxt/l+CZ+kpVeG0qMtkIaNO5XW
zAKWN2wciCy0Fh/8Dqn5J6e16JXNwxj7e06dH431qns7y6MSZkZE4MpePtBonMT/bkN/ne3OO/U0
NyiMDyLpQL1hZkm9w9GcIoMMj9lJAnv9luixaKVROrHivS1kHjRtxp6yPBqJTVdcAhkhpwewmX1S
l7LsSi+fdpIfXhC10lb9s+RZT0av5a/7cZhG8Bs/C/zyRe5MFeZKAEpGcGWNTwXfsIq/1HcYDZaR
5/Mg5X2uoRyePeLlkporuaj6H70pF6I8r9UapXehKPtdKDI/c6Z32nBw4Lj823jJiS+3bZkc6Ffq
/7io8S4jXVZZZGKFwy+MRacytzuENRwORQMBj507XUOdMM9jzsBQNNbNiO/4HCSgJLDUzXhHSR/3
SrwkmczRqHICgCxYxXc52Ld98XZpQ+rxqgJH/7jyPu+OHpdf1WAnLiJbSDdqDL8cIWGQk26STxLY
9du4mrHPIy6gpwDVhhRDFarrBomagOZHhWhYpljHLj/Zv/VJurhFWK238aWQiVn6iY5p9ny62Ts4
Zq0gjfYif2cJKXRiTxV9dawnzyrcxf9Ri/e1utYKGYCZdxNMEhuGQdtIunE4VInfMpucOa8ByZ5d
Rw/QfbNEJ1aJxLsbPbUzZATrEQWH2AKRwozPFTQGD96M4/llYVxRqoVu/Kq/rpuj3yDFa81tqwvj
JyjLcbF+VjML7D6O94ihmba32sJHAMVuhoyoWRpC6YfoWCWAJm2iC9W/MtVJUctZ7yJVyRbofrHf
bvkwC994EGShVRRR9q4f7BO1sPKUteKxJ/KS+hwQOT6f9eE5KjptbuCUs6E/kEDtKK2mKgd8HAOA
oQHu73LfB7YI2jd+Lx5UvAxghWCS7HwlMYKR2i3caCAK8Hrs4GyN69pWK65Q+VrKN80aV+ykpnWy
9kX4b0fRwWYpEHwImJQq+PhMROfpO+ix36YwrYNaHm5jby3H8o3ceK4CseGUtgAkLfGflVPBz15q
La3dkCnJnV92p+YHuoy1KEjXFglqaQC1rUcpUUskRnRLOmP52vL5XZQJ6lmTafxiX9FnYfBpOQ/e
fpnHKil6VPbyxryyoAy/6tAkSJZy9tcqytjQRBJTXpIEdjz541Rdn9X1Bufir9sHcIAYJs/iSTHW
P0R22xzYQSqWxe/IbX6tT3bjKTB1Os17YSgK4R1yUGxViFlCFV9paWOaA6w6u/V+vs7c3zvo2h1q
ErdizIAuGjqbgQQedBOhph4SXrxJ8lNUX72vhVWx2YMoAgdWhKEgQ25rzIF5ZVvjSpE0KruLIr0V
N31PAvc2nX90Slrlo/hnMPnjO26GMZbvXUdRvXtqKPo8jb5ax/q+14EJgMB/pcTlbM2azDJ0qwDT
b6nUNZEm1BHGd5CLCg/3n5AO5Ek+vBFiQjLKwTcNcYPtMOhdkLhYkDu41k5SHIkGehibC8E/X3I0
E/yGCNEntBP+fRxlHFM/ACgWfbf20TOU4I2y4FcAxIAuepruFpM1p76EMnU1UHbudoYBzfJvrzC5
jBEVvxzbNngOUbacKWSHAKg+nlJSSx5wzLXUgROD0d2VbUez5Uns/B7AazECjaajCkdvhZkibCsx
M/9s4kNqeiZAfjAKWWjjaJqeB2zAoUK7RqkhW2SEnrunt0fQYP4L72QJpkjCiz5sl4PmzyleRble
zGgOVX7QFDFcP7NUkMzcOWtDAeIidLIPG0m1RB8UFv6V5Bm9otzgfzF3ul9+vvq70SpWD8NN0pEB
SSlpC07DbjrS8js8KAaCTgebzfVPZJbMCrk/qY3xaT56VUN3x13VBKuYNnWNxG+SJQDP6myf8PbX
BaRvwMMEKj8lOTxaVcTzapamRm+9asQ3zgxHFij0mwgy3dRpZL6ELr340HBkhfHvb1i94/dxZAlq
StFkfjvYO0GjRPcpg2wZ/94Q7yF91nGA1curEI57WnAULSosiTkMxupSbLWFK+PTyT3GyBCMqw/C
6T0c7SyA9MF/J7WMILx6WXcvjshKJqhCLjIY391l1b+6APTYAm1gY39rkrnupVKYs2cJD7qsjJ8C
hDYhbxbTsOUdV9AZqh9zQCs+80Zh8p0fe8lqUFY6sjbgBd03MlMKygb2U+ROE0j0woMDsoBvliA0
5PRdx74XWzizOiBshJ4qr0iCLTF4ykZq8ZEkn7kNaIqE7Wrl2Iy+2ns4QNsaGrQBCd+Vl8jzh/SI
SB/HjMdXjaj+yPs+W8CusWfevMZPZueREUu2v1pCqKqa25U6vpcJv/BZkBUFn3nseRhSB+aTTgwS
E7WS3awkUdb/+l/Cs76ziCw7bLrjOQ5JdmsSPfXSEayI2R6M6SijdWB4lbGK6OqqTVjqZDZZh7/D
O816O7YtRj4SauRt+LDG+QM1rbhkEkzBLEfsLjYSqpstNnCJqHvKl+DlxnkePAmx5WfS1VdzTD7j
oZmHsiB1UnCTgQfuGenJZU/r1Mt/Aw/Kszph9I9u0NVxSWUveR7pgCMg1d8scJkx0765dRLamK/q
yQ19ogfBWBXZLrgwZYFb+FEtR5AWeWq3qq10Q5IIRyu3HJkcAUYbc0Z+iOpgjXm5zZefl+amHrSy
tMeGlfcI6f7J6PtkRZxQHfT9zso4L6Kw8vR0Hep+zDbSIda411rn4PAToCXGqbcHQxXaw1ILHF2k
x6b2Ydt1vTLyF/O+gEj/wMUGdlyPzYr0hsX/Rwf/hRf1j5NnWS7qQJYrE1loLnPOqg1BQbTcqI3O
fu5+Q4ANEuU5M/mqJZeaBgWgZaXr6Pk0sDfFwJzr7vvIYQjk17OioSkJi/gBwdCJF/xtfHtoP2cp
c7H/lfJBBuPi7I335JNrbQ3TXPI+X9RaXCUjbdw6ddxUHPzAel10ClBsOfgnS0Za5jyQQm8tCJbl
lvPG9NuGaHuxYvjaEfwj6AKOVMzLCTPp7QN0oofzsZcfcKfzML33s6I4Z0zLxxBPUkfraunvG5cX
hqF3lEg2zzww1r24ijityv5pxWsVdp0tltDp1JLQglT3YywDdc0dxGVlVVg4QYgyXqYgDkOlnMjN
1On/wbkxymP6SrOcd0etTfjWyzeUGdiv/2RngfeYbY31mTrh3RgBCk1fILcOI95IhbvaJtHxwiyv
YzXvE5qKNW+bO0tA4KZXUbBa0Yca/yRd7r36Bo310heQfxiT+teAFJc1NAEsaZ1Km7EAdLnCHaUk
6LgSl08I3+9TEPbm57Z3t9fItQg2iXjWJ+t1t+4kUeZbrcp6m8g1zojz//qy8wjU512Cjcnqgn5f
lX1G3zVySxuLE08kMoK7Ny9S2kt8LO+KTAn1ZLFny3CxjBZ8zQFK7v0Rkc29S1vXdJwZsEHcK7sG
Dsi2sOHOWTfrOCBGcsJB4Zu4f7TVjRkgcW7A2J/q5e3CeIdIfshY1Cunzf0aFqVgOAgv9zYuUGJv
4bEuBdvseIaPGB2RQ+INlwI7mD/VAE7e+NkEWPBKs6psEww5OB5+OMrMzPtcyIVjn+lTMCPLOOR5
Jnj7Dde/6xkR6Oju8V4sq7O+no3FQ3agaXe0MBtHBlEqobEUgMaPcmuC7STfnpB3Mx3Xa+IB6T36
WqMcgc/53ekvejENBTHDWuYPL467JQ3D54ySddc4RE5+c3mGres0XjSXjYM4djFM1m0Czq4W3Ppn
AI6qmklstHoVavQpEj6b8gPzBFT15qOdn/MQLmxZZMHWDq8CjsoNhiSWlOA+4dppytPbcpknhBA5
7fm5qO67Os9wXZSu1et+aVbooSNCUsbjMYkIKST1/nP5IHou1Ndzup7amoCsWCMCK7uyub2g92Fr
P5fOPk5ZEtXxnG4S4tZv71mXwWsKR3sOfCFHrvn2/s/nxuZ+8LSsjgvdntw8vsd423dPNjUkRgz0
55zEY5G5y+jB16F0gJfa6qtepUNiqUqeynUTu3pPux5qZNWkOfKeOlsdX3j3Jclo5fGakCiV8tWJ
klb/u8m6QHiGrrlI0Z7mFKpJEDPLEMNYk/upmJjQLOaIbvETdaqs2DsBD3TCFutjRYAmA0BCzm+0
VWkwu5I2Aq5BGMG4FPw5+hqML7LbMzTuXAhuq5L7ARpzB7+FEiRrtiakHrS6pIwWXv79TAEesE08
wA8bFJ4V0J3XDJHsPv/LK0wLTUqbLkSCpWX4RYfhQ7aLam/tXI5d8dXZB2Lq4zdjZAr1Q7hqlBn6
tV+yyeDVNycsDzAlbcm6yVrDEHVUZ6cfdtb/7MnTbdarO5DTWAMCd0WTb65CJFaGprJVAD8Zi8JI
yyG6SSUMy5hsc5LWyzovTBBhs3owcYGse4rStqyql2zAk5PzPcShMQY0PbKIio2hC/iN9RyZQcX1
hQEtu5Y7DJn4CLRlziI9/EYDaILK88UUM7E3G5j+l20AT1PjOmYzREm0Pkd2auDEyOqvAPuxLZ/B
YhLrtDc/pYJFQg2gZ+RG/MPk6ShnYk5pRfq3ujtT22vfkVjetgwvDDizMcM3XpcI95cJIkyKtfqj
fXzmflJD+vCRxL3KMHuUJ6xRR4LzVIjwC0fsS3QHpqhoul9bEXZ3cAPVqL4gVlOjcuvD3o5Vqk21
ZzOwOXD9aTAaIxYPJ0rQ1X2Dj0b98WE7DEKi9/Ycusijn45bkX7XZCB4C5yZet3Njuy12zXst8ri
IZ5Xyn6kFGkGWkPfiCAjGysjzQBb5oPDccWgZ5ZorsDvAJc8t+kdvEwTAf1zHomTVvzswq5VAI68
bqk5/xvXmcBMVr5SdSpbEcNnB/4d9AkJ+Vfv2ZkuQ55XKy9FCDrrh8HhGrWtfX7e0L9eVKG6oFs7
1Kv6otFQpyZ8VPXzPHAXpv+s4W3D7irr1BRxGySpd7yc/83CtGM4BQq7Yb6gYL+mJHYk7vX6gDK0
GYL1sRKCsYSkphWP85TmqScARyFM+IzHHd8IgsBMsWaCZZi736HL57ZR6Zvb+/LEj7m0+XEPbVI/
quaQ3ttmt+Bj3cpat1gRpQwagl/xyQep8qJuGEyxTkJ6No8dLkzcz4az8HZ3c0sx02wk2N8afb96
BoWIuHE0q/ZkffzbHYn6Y4mucrZyvfOuQCUC8OJD9y8U2omKsh83LCJyTQSQudNTcFy6oMmlenPH
H2EG6a1dUcVJdsC1BJpGl3sENc06s09Vm1hJ5GqgwEHCuhSRGr+RXvh6+ABd43oaV2AJvw96epYB
nbsBga4kd4EGHyc1kwD5H/yFWLPgEodTR5R6hHzGAauVYvTZ9/0TZh52hvcH4zogFoEZiUbvPK3E
GbcV7KVr0BJxKknNF4ACPLRUM1FUgiTTpRNpfnSTYeN+poweUYu5SEHIA71aHqfRDbTj0pZAgER3
bZoST+gZ4X5mS8usjh6IbL29CFxTGkQdLcZzuaeMiIp+BjKzBxxpwDwgKHJ71bdVhz1I4ypuXQDm
9b5A5aZtdw1ELaeKHbbjdcBXdv9/3iCr05gdZ8FbbULaLoQJn/7Y6Ws+2RhKYlO0xQVDQmwYX8Zl
qQvPq49jdNVJWizJV5e3RbGbk3380rvQ4q2wzIaa0UW9hLVwseQTxe8Y0latNqGDlA/WSrbeEd1h
jYwXyO28+L2rcraU0CkRLSiFWgHrnVnPn7S+TYDYWPNGJgLsQJi6ltllwwCf/o6giGumJzX8R36v
QvFUFZokolMBOQYQ7kS/PS3WFEx0WGR3q/YZmY+KgBKMZ30mwJq8FxZN/FDPnEleyZnrzl2gF/P1
hsoGDEfG+m2UEWY4EWxGeb4AAP5duEwWNg4hX0O17TlqrMGkwRxo4u7e+ZPpCD5jLHTL8u5wVndJ
vR2qxCKSnr8Gg69NRxwyIz8Ltbt2MlLxJPIHWEHSxs/pfvWNdcYGGM/84mDtaCD3JcinolD0fUkI
v1gl+CW7HQPR5WMtdNO4hblE780r5TYsgCY82gJZpWe5WRAKXtwrSALna1uJMrVpDpTVydLclMNg
q5NjPadfLLXKF53dpKPXNdf8cDraomjLr/H0mBD2HVMPyJKSvq4NqwBUsWFRE8AfACNUfycR14/i
YCyRxRU1Q/lmuJDL40SUmxPdgLtKVSwaF7Y9n9tbNj6GKTdUu3Imj9qqSxRVyQRyK9iFNxhe2nES
XwLH5lpJQFs+XZ1fsvwTIyAL5GPZIzhRbRe3SPNlGg+KQCB9Lm2Ha4Uod7nERxulVwC22A7xF4hi
WSjAu8VnuceV7jU/vYHtYPPSNZMhDSOwSQbVPllYXAIX6dCOMyllv58GscM7/cF8qQPEBwu1YJpR
JLsGGzgPovkaQf26uayoWkF3AVI+34V0YTW4p+u3GLb3+9o5m3wQmcy2JoXUdP/qiSa2HabwyFUi
4HB1aQs0/JY0mesSjkhJDNE9mwqz9mu7RnI26UXRyEbCnd3kkLZxdk01YhkqfRSJw+wlsy52laFy
61hVxbEDD4egmAOYdJs2itkjXzWSMrErc0P/+PdT7ah/4eBHkXEDdPjhrt0yMPskm4EYlgzv8wr0
uMmSpS8uttV7+lIcbk9udR9/HktONILDRVIMEzQ+l8X6syvdWICdjDBkcJFxPC9geue1V0rtfrs8
10MXBaWSKmEOHj0F4nDqvWDs8INAtJifMOdBigS0HQMiObDvbflB2qIhADkRokWMj0qKkstygaDy
Nea+3fusoJ3gs37LnKE8DOW+lOK1xru3EHhrMJov9aKaBu7PEDOTRmrQ1xh/qBI8GXkZl910FHLy
SCfUYH+1Ngx8b1cz0Oc38rpjMMV76RCYEEcspEyIpF6Em6uqP/K0xqoQ2LrHVsnNCru1XjMd3Kyf
E9DlTc2ffyl493u2J9MjaO4oQdV6DuAgi/suWeL+fE68lHgk+EkrP+thZedR/k8m42ePQ3SkDMtm
nmq+tuyo0mBdb+sT3Wz8MEKqEGKm49nlx89t4uQx6t5XMudCghxOl4PkqH8iyyVWstbXYGyr5vvR
QAFdAflt56rT4+mnwGl7CisHUGns5n1f/73d/exD2SPhYWl1Ycxy33l9qePZFMS3Y2o896TnxsY9
cdTi/Cv/K+rD4MjuSlMhn6ydWxs388soxRL+TtxlQx4lvDh4Qr2gM6EVTN1BJlZ/V9m6qPnHP4n9
e5k1Y9yFWiP8dLfsL57gffZXMaVLeFri2azjWzPfHu/OR+os+teV/4W8OVNA5shfgk0gtwOaMFAJ
VrA2i4L2CSt4yb5hv9OfFTMJyiNjA29JiLJnpmV4UY2zjR0sjA59u166EmJWj78nBTSAWueH3JWH
j5Fsn5ETo+7T7YcLxpmpKVOHB+yThGd4TjFefEeCnSp54VN0pdC6mTuGKQ01EWJLggcXwxyffbOc
R15ZxEyZAPEw3TtKvJ8ybM5nPyjRBtKCQ3Dpchlcp/fp/fc3roCCg3ScyzljCgNBX8ek88VRL3fh
Nq4aLWQ+yPNRAIiIDVPnROD7SMPkLz38L2e/5DW9qKaxMBVN6HEVfV7VytHyOiEBHPPU4uAyybrY
AUP6u2707kYIfOaX04TFsZCa6e8ejS5khrA/hrSc1L1QFLmRn2jAsjon31iMObvGAvw51AR0hZqx
xSJQl5iOEbyniiBz1WS0PMZzVD5WPWl+XXw+tXnVbR2BmiOkfYMkY8ZZ+h/S6yc00OqyVYw3AOx4
R8RH69GEQGicpSbtKUrgdpohNiZs+o+fz6obPAcCzFEObKYFvchcCX+uoB3Xb3uFQCiQpoTjc2Ly
2q8VRmNpvM8muuNs8PD/oWnWHNOJxmFceg+201Chfjk9h9z62NpDCi+fJ4A1B9guz0GNbMq6/C0y
GhrE7d8NtPldHVd8GGn3UWUG9uWjXri/CTYiimJhClshMmEA1DMebvdrAGwv//SiWlGEBuxPi221
dF57jR/AzszBuvsJJKqKLPLBZLXGsQCVHQFOxP4Mj7VGPvlZYI50cs3FA4lBptwOanmFiu44uG+A
H4Ar9+47t2m0vNKr+GmAljoXrfxTxjFWb9nT1HUmo4S5BZcIlHGzwFgPCxaWwiFYcEVDf/VtsAjc
NSO57PNJZ9/hMhMyF2sNB+3u6fDAbMImX7YLmxUaYcmjY1iT1QAFbbKkM00FzEINu058EGE8tPBH
cBuEq/AAMAcZQvVv/7wkw/syNERUq0R/Uu8vV/h0z+jFNI5L3bCKwfjCslm+kp7MasZ98ockND6y
vESkn54LL2ftQ1us9LKQKnbAE+VY5K3tiDVq1k9qfE6VeOjWsZGuK/uoN/VzDd8FLQNjjopL2GEC
GG7XhISUHguDFb0kiJhuJ7xH6HwKLpE8KdCOQfblQbUSektu3Q4wSSAVr93vwNwdg2CKS11EbL90
JgxGG+EHcXsMn2ZFKFwosoLCdwbUbu36g2eTH6W+GYLdw4bTY379LUuQCd5TIFJoxMJyKreYXCz7
zuHfHeEX8NwOqJqqTAbdDyQZWgbpGNuVvLZdI59t80ll9I2+X4OplrnggFYLkCr1eTfi9ztX5f4e
WbhvbcbLKMJwi/a3//JYjAs5j+MbPsPH8RB3ECqv4HweRO8aRMN10s8GdRzLMIl3v+S/zO1O/XXB
UBO+R4n2rJgL2Iakcyg9RxR1g/deZkiYU3ENDdR09nrNntgLp5jkN7ZHvFpV5H+ZoO7NFalbVSvY
lrsgFxvrSLiwy5pKoJOIlrM3Q2RGUJ9ipPmzroMhqa9PhD6j+H8EyEyvDCTELF8ycUl6PzRd6lmP
jGw00DZUh5YKNpgl4Ltoj4CrclY2UrSmBSO//dPlH9wmwy767EveHJ7fWHsUrg2Y64igKde/IJ3u
CQibbJUztzHN6uEzBTJMcHEFBieKEf0X6n9hcmsrj00HToVnoaLMOp8LCdPRSEOSucs2f5+JGPdn
Ma8FYTMzxUW9H2DNfTrtFRihLeCEHSlGoyIAMkkAl7zYn2qGO/JrwLYxCuhgC2iJzX//6K+B5fP3
DslM8gAfm8McTqD5UQ7PV3J4EjNHUPSujoSuxGIIe6zffBY3XeTusZTYmODbLigEf/guoPMrzD2r
DLdd10M02eNhGxQIXb3QgpmT1jYjHEL+KxGLOmcr39ywFeCA5A7UPAZo21fTTpT6WHvgtg6TuCt8
MuDtQlLBrG+pya0BJfWWvyyvByDLXbPl5TldWFJ4VA0xKHOLiSCgTcMhNi9K3VnkRoFkSzACJT7/
YmQtfe/uuDkNxDMmQdepxIm9hevg8vPetofzWJ04ccCwm4ynwEaYjiUNrJRLikr3Bd/FDYCXYPFz
s0+IuU05JxWoMHzsBVJDMVQEy+Q0oM0rbNNj3SjlEF7c+bbM2Uc9r78AKjojwDDhhkVoLZOiwY7l
hBoR7XQ+mlPEeb28HtOO093sHPb8RdCU3a4UwM561xqNc+OYpOmQHNCFR8OwUG0HyYa2H/yA2No2
cZ1LkcyneUGXI2PtKpoq/ZenBEOvgjhqTizaEJ+QdAKh0BrRSsMaPUq+x1eRs217WuB/09OzYKgz
NGQn3uHclFLmPqoXVtweDGtDsReBCe2MfffP5zFAQGfFRaQ5kxY5YH9a9G9CATa9j0Emhjcjp2f8
qWOdibHKx1Fq9o7GkheOUMpUueQBNVMBjfmS1nsRsgT6mfl3+e+CQ27+KoUA5yh3D2JW2L/tNX+P
oYTRRgcZN6gxtgn4X8Uxx4ZCsmxGO6FDQ1vqFb0MPhHvT/nk+JhePKgt58lUfYIxfVh5GCCKsJRF
603rycb+HZ7VKcSMu21QHpMpo4SIh+7mj1KBsFT/48ZZkveWsEs2gN/ZL/bVJ8E9v64zjAEKffbz
gKx3iMratYzVvsGXtnaCSM2212hJ7q7dbU5aee3ty/gqmNdgTFG0OiS1gkgglokA/Yqqj2mKDTOB
5lAt4S/z2M6igXmO8Mgp7CsPsSZ7Y1q3kCo62H1ZjuWhIgXvDoZPTdNCierjDdd60NKyG1KwjAcp
94QalIFZnCADhOu2947mVX4doDoUvkisCg/JYjxMOczYJqdnJWrsXF/KbBZhaPaizYJKyuXPNM6F
WacF3AAkSf2j9UXBLp4ovO6tyes+yGrkAh/wNAVNQzBUr4kblXIZGZmc6n0aTb6y9jqIRgBkBEuE
5nApbTA8psY8Cjt2+D9VfqPh2NMCsqrENXcOKOeGSa/kmRuHt+O6TFSmTRxoTk+w8UXLpMjeqF8W
Wc3g3UKxRrvlYjZrzbnlCFlPWIf+rILAU3LT1Zq2lfpemxJ7Om8sBaznXjqblDYOlOnu275tkwoQ
jqfSOnvz6w83/qt9HreLwRR2vAUjOQIcLPKHneA3aRnVN/aW61Wsp52hrIBXykvNbymJVwp5bbjx
jg7Go1Gs5WqRYFsq3O9ROT8/ELx8BiE/8U8DN21PeYXwI7rj22npYmw4BOECLes8byDcaRuS7UJf
gRKdvuwmR1o8TVtCkxmejc3xXU42miJoQ0TZdek0wJD58cLcDXJIzyq4QfdTAuCgPNOOmqMgI9dK
9RUG3+kciJ1l0ouu9hpHiar9oapXd4Yr13g++0bws56y+0KvdH0n+y54vYyOblsy/SohvwR0vMww
0A/XJD8P2kwPVZgP0HmtM53QHUm5BEcS4qsyww9LF4AG1hpRarjzGa8HOayT0alsmb1ZrmqRFHeI
vBF/2ZAxrtn6vxLyepZGqVngrGo/LKA3b5mHRxLFJjAX+6BthoZ1bFuZPpcHolO5F7HjMIubkMtP
xZEnsNNe7n+Kj+gYJsRODXWl8ub3ZVleZTAECZfsrRa2TsVLjvJwisZWMQ+hFt+i5FpImLX80d50
ifPLVLGehdKF/oGoHEWzxyKzoDLXZ/bUsRhf/SWFL5V+SlwOCU3ealQyzxGNCXpd/FoC1Z5t6w4F
x3nfAM0qlO+79myybohrWFDtlVN1lvn4ehF5J17tItyqTnrFAoQqgYOCqrbjSzRGu9+kIRcMPyHO
hsYxZfMsWElFZaf9MZr+dLd/mCjsW4yLamZfowU9PZqENlcT3WA69iYOA8GGfyMhbpMVnp2AKSqq
fBPqT58igVH2cMqKyTy5sftkapN6QvxMQj56gUtnIkZtsfXZWewnOuuwjFHljWIYUvwhtwUig6Lj
cNhTL4tkBACZ1e5KrV+5s7me/K1asxUuScgnuXeh71JNYF2vlgHxGXuTHfoXQ/+iA2za9nkMi3vJ
nSXsW+ViEU5Qoq0WWoG9gLD/zp4uvtUqGOh9S5GrI1/CMkg66aPlbCtLhtseIhoDqA57Rzd+o0K5
ASp8KXSEWQTigbNx0P07Hhh4opxLXV29LbosJjm6YYb+AfwKVvGRXpH8/VOsER8wH/0zCwxGP3fg
aSiglGr2SgSjgUVG9l0FvY3WqbCClXwxttir3qRkx5AFR7BOikOoHGm2tz+owRIkpgeINbZIcwSx
UVvUB9FONk8h2szVjd/WsJJg5mQUEXXrTLAPPbjR6PNyCbr7wz81PC7zcoL5xND/PP6LoF57w87y
2VPYWmt9ax02kP2vEr1UZJ9k91IEwh6TXUTjvI2KweoS1aR3n8N7ly+FJogdefJKSUneakRR2zAo
uVaScoq7E2Vsp4b9i0paSQsqWRcbksuyLr21gsp8w36otoC3Wn4TLjFasBxmTFS+9MjGQgSML1w1
T07+3bi8Aa3Bkkuyt3jVMDsWrD/idB8YppDIRsT8vp3Ct0/NcSqdkmJXrMTQIG4Sm4R2TtpZjbGL
ciK4rhy8Z4du2YUYji1pqUmH1e3t5jRaiHjLkAwliZTgJM/J99OoWH/mI5/+3+LHiwTRVTjTtkCW
bO26wzPIl+uWq6u2jxGSIBYjT0tGUTxPnmMHqq8hAtY1/Cr1BPbbLaKke74atQfa21y4kBUFF+Ke
94CbqAt1aIFgVHrc6JguzYUMULmaNntTQaej5xnCvTG1kucg6hU7ya4arQuYQku4Qbxb9LFLHZuD
TfzEmafxD1/GrQ8gSI33zHl1AndbTnd5J7wqFzLMOTJT7tOid7M/ZmMtAtEBqNSkkLpCjDJKsz8F
ATZ8pAOIc6y5emvvGT4PLsuTxO72fz84gABpwncl+oUnU2U1UeKyxo6sAXlKpFdnPaBjxOlnGxQa
RucK+RmXrIRdlern+jbujALkgdalAbvVuAcmmmzUFWKXHqKTWMffOah5RMz9Wfvdjwctnz0Nit38
Ws6gqgUi/mKmoSA2YgN8L+cJHRC/v0gLSY3lw1DzT5Cme7+YXAonTQloEhuJi5AhP7liQ/tAJdWn
XiFZfqN68rwlGpVT9IjpMSjrc+XONDpOr3fgROUxrsPKzDpxcGlhA8GqkZWi8sMkl0MPfv9dsqA8
iNOe5/jjSs4NOydkYEzPm6oTI6oOz4b7fSMBpSPV//U32hZTTODVF55dHZqoYlnbxk89AWtqYosV
EmR7KOAVmpKNTutAiB6bFlWcr4HaZlEFUxLJp2bbdMDHjgo5UiqFvYx+Y26LOPpypMmUBq9kTgM7
nhQS4yNT4hbDgt9djUZ2zOOHDEf9A5MCDr+cxnP5cpSvNbSlwJe83/Zc4CEI4g6USwOkzAe8aE3C
wegwsBBQxm7Yte9qoPwYWcrP+MRhJZh6sb3VRf/f0P0l9p/p/BfaWEQdBrsmey8pRrtxYgbAQ/H8
uGcrbj+oqlOUld5WCeV3eGaMxILNC7/XFAd8L7G+lvadbQEgTC7bIR4VTdyRDNK+wOft8Zq68y9/
4WgkJUkbZoxKz287hwob3OjeLTjtAU5k9LzLIzS5ezrpoLSo6f4dftkUWrIfrN0ZUYFE8RCfpc80
+N90Yf6ndGwtqgKWGdXIf/7Dk39MbMWPivi6nQ+mZcTf2+JewrhEykOapm+u9SE4Trs9dJLwZTWX
PlnlZId47UW7UI10FKmwV3FkbyuUAXJYrv6bR4xv3sFXF8uaWAtkf26YsjqYHh3pEJjkbbPLqziF
OjRGKTeiXvpmPWQRglfDHP8Ta91QwC4h48J9tju50zQHgqRUDzOnhZgqN+yBtxZMhItTaoyLvPjP
L2gZT2N/1j4S+NnZcmLOVxSfWuOlgwpLTyPQ5fI7pD5InUKhhRcmFOT5bWe8D6tjBtN+73aVyYio
pdC3kbaU/5wmJgHU8ITNlhs5iuIcZzBVSHu7CFLqdvLXNk9z/40q0O6kJSCpivsHMHoECq/vzRCp
qOthLOiSWw1kBxh4YOHlWHMEX9jk5/YSeJeSFTECMTHKk5vkFWIjZQaiAPwdsy/dv9rB0Ka8rCQ8
QIsCIc3bEeMi2UDh1xzGcPuxXH2shuKwVRvfVohCyexF128FpMYvuGvh1oLDI7en+ZUH2+vRsCnn
VUA/O1dPgqZfkgzRMRkVLH6lUwHPA0hj18LK5T8wZIb33D/wELw7NdQOuIsv9EqAuO4jvgwgAOYN
DLO7ODH8pkVlQYxK2Tuuu3/qdmCGkgM20hPum4vILew4rVUgq+3OikwtVIiRNzhLrJ0nV983eQ7Q
R8HPhNaWGaxe1hegxJM/X6mXWiulVc4KOK1kuUhspIawMGdMPV7FF1HOETMdDaa7MLVEBq/PH8Bq
2MB0FyzmisQw+NqLRrzK+/t88OHQACEpv16icaZciJKebqwT0xY4ZkBKeCRpdFQefx+VLDYdPsh6
ZHQpQXkMr3jFUOM0QnusjAYkS8MCYLL+9Fi8qEEwvbba/DypKqwuFROv6qPJqhHLaDJyhc6u9jRr
q5kcy32yWEuWro5mqVdVrHBI+3jTPk7zPFK+iAdiRh09sHuIroZdo0qabJ1E++MvBOSldv4iN0k0
/XT1YJIwM4tSzxacy7sfhWiF9msqe+un3mP0REeM5n9OTZtuZXDv8ClaOLjK84SrQ0JpY1WfZIPo
DsBooimmPjQXHxkGptnbFOiYMKIzfRMAAL/aPNH2iehEN2Fq+TAfR6/2Nn+Wsb/3us4VjmDN/NlU
Aj5RfiTP5QCBGvqC7HtMwBVA6gksheCZWr7o2Vs0itpqp6OI3ytoDCrtD7M1cEQM/ZnTxuFTTkX6
vMfSp2rrcOUFuqMIGlvE8yL0D41bKn3mWUi3YPV5Ty10FlUZQZ1Y8FSTbvwMlQRohoqJ+NoFSU7O
BDbz7hHcvod2lDuoA+c+v1gw32bVYZAtzv8IezFwtwQJ/3SJ1RTNFDvePFZJxqg+VpjPHOYwGJ00
hZAVKHdwVaxZ1G5/lQtKAyRXKeaznP951DQDi145Sbmv6hUthiaFJ7Vy2//uneGblBvEIp+Wh6wB
9YmzCZlXgz/6ej+YqBV5cLw7f80hsAeddsUl1g3LCo5sSvb/CgssdMcXkNlG2A4VnplQKYn7VPJb
WXEhW/zbrCDx/69a0ituzmbryHPep7J66CFfFh3MzWDifczsRb32M/sTmnv8ruu8jsSLw/NZxFEA
Efnr151uzSMz2Dbd/qHN4TTQTPzprULcaC/H2YqPrNckDuYT7dUF/GAIKBuhP6eqg06IOFR/Ko/y
gxjrRB7NJCE8xa1OZH/eItdL7aee2Nz65EMJarfMM4898Hup4MQXk/UHcpkrSlPxwhStf8mFNKZw
paKp8xwu8Yr9HXwWzQ/PuLbO3O2j031OY5SA5y3KLpjsg0VfmxNUhmhOGDLOh/sQ46CaB3YF+KVK
T3lv5/mCMU9A0p/Ia8X021sMmtlXh1MLWO04R83SQeZWCTvcmd2PTsFk//3ztBL27p7NeVRFR+02
Sze9Q7szWaMvVoIaPLUDKti6ux4gXFqLTAFUMmKbmonze4rwFS9jzJQq2EOsbNy5hfEFXfAQfGQB
lYmpXMZ2CWQaNKq25vwgAy4GYD4Jgo3xyrJ26vwEc4PNYpswvd5hR5reGGfQyoL0S+MQ1spNeL5h
+WULGa9r3YLUd8FK+ZLAWx0E8+rK3AaNHujP6OdrQGNE0gZcIwmfWOtbDmktmWt7F6xNYHN5pTku
dW1EdFtJ+4uNX2QaO5BxBDWNu922l5RDEUj0c3Mo+/nKHKnxaRUH7g0vKSSr7NeCwa3WiHitMJiY
4wX0zd2Vpqks+XnpkS56eL25nQ+S2WupQO6Ky5C3Ov8xCvEfjLHzLGZQqgFXtBp2BdwjR9vRnQQD
5Xz5te2x21z50nwbFJtsrTK//QgOkDaIHe8CHLHgPzM64z055qQ1TxBpsGTFqntbErRByJO8vZKt
Th9Xk2c4ZoFLSSMrBbDFWsMidpVbzqpyZxrwtl07PMB65y3m5L+4PncKodcWv07/0trZV0ztBS1b
H90M3xjP9YfVkifQ+PAjdfvNALiQ3CDDiA5LZFxR8dMb5EAiK/pd8bmgLY5khU59c0/NG1aogrkS
iEtlWbcoD8AycmC2sl8C6q69qzmaZqH3yIo1AAf2uQiIq7ZppObGUsFdUqkgxodSOR61lEf5Wqz+
krBXyOTh0afL9+LswLsZ9/Lb8MmLg22ObYWs4Y0S4iUVemWHAM+3CjsYamIXqxOxJ0nXvEn28SnY
Rh27O9EJTpgkl8G2TqJ6Am4kLv1RJ3uw+CUTzofmCc8ZweNDFU0XDfvAuaf4XHVU6e98ZJ2EgcRm
JW3M8IXL89WMMk/t2KiBPNjHMSXmHuvfN8J4nIcucctnZqNncKACH4yp7KjVYaklrBYeKGy1bDpk
IHWu2sW2zGGJC+PrZHp//oQAk1TSi5DMtQ7kGapF05kj6NdC6NhWTBhOmiDbXm/1tFqJBomvVyGk
FfZptvvFIW/s/35QDyuFIz1mp/RZY+chAyvr0kUwRKgdhdbKbWN0hiZSAM3fHD6PXqS/bKMYGz69
Vpl04byVbPRlV6BLUFZ03nKkmrnhia5HA1N98Ti/Q17r37P51Dprih8htlBTkQnUHmQ5iZd4zfO4
Fd/NMej74NDrsq8nydvYlsAvsudQTXR5OHoQqtNGe8QoTw6E32u2q3CR26IXqituIKCkm4REOPP8
4TVOtnNLkrsF3fWFaugaluzWm6HKRucigQ+m0IS9YqNrP2NgOBZML3DLvJ38P6zKNLoel63eFO7E
3n/falTP2W3FsyeaEF5cS2jgNJ0/uzo1xcmXLKtx/k0RrguTVIE2CZPM0tz7JpEH3a15R7dUQ9LE
JtQ6AFN/fM5Cf4hOHNp2jL4EPBShsmEboKpkfa6H8aK0s03PDXZKSUng/InbZZsdN+y1navtwbsf
0gl5+XaZsK4khE/AcStNaRxeG/cNpGA3pTl9q698akgMxAWaRDhJ/nTP70Gxf33GJH0Cure4IM8k
mwQ8gDWHvV0SqxIGIHjVstRpIEQkCgdzGn1n5XLdqWGjD6VsfntG2BwYupwbbNzaBaMchFoOwZFH
IgL6OTVNR9JX/mCLK+nHEHbr23lB71BFBgYhBV25f5MgM+Ekq9J1dKHmmM/F+KLCvPH57YAMB5jQ
LvVfLUD542+BTs3AIa2PyPMqMIFwRyHaoVwQML2uw9WtKDVM8PuQQTiCRvBiAHdQitUncl5KwysH
q9HLrJqwG0oiePSjNVT76q9HB8sKuUtGzLg89stO3VZ1E15FJlXPOg2ryqjVt6F58ifXQn38gBYA
ofVJnWBLeA91qHtwHlVGE0oorYIubpWbLWpF8iRkcF7lvrh9dHAXyEo7oU7EG3jpFjMmVvp3uOuU
5VO/xVzqTHKf6OE9Pw3YvKg1Bx7e5nvxD6RmsHJW6fRzO7ohjc4CeGsw6tH0J0kTzOj21Kl5Q309
LBuEvTLc2zHDf7TcdWYMMiJi9Z2EVa4jG9KLorrgPCZ1SPLgXnilKr24fpCXe9TUrb84xP4a2gtj
zMUEBzdZqJp+9nIZeWcugPqYZMGUzisGx/j0OgFopWrgDW2vnMKOjxnJQO0VMRFg0j6m4VjWHN6X
bnXLsFegXiZ61YC2bFTNu30GEuTJhGO6cV3ZAYuG200nYIaAAjto5rbnLi3AomTjzXPg7sZ3pQLY
NdsRvxW4GlfFnw3+SBs1fzb3BrnYvjBykFjLBR4Tt+5vgbD6uq/bkpUaZ97eU5QSF5cUEzjL/i6k
HM02WNKfeSDiBfoveELm819AKsFBawRWCgpiN23EUAaHzVCJDFIaPepEVMP21Eho3Fc/GcOE/B5L
uiB26s/7PX8kqsD1fR5HxXY/njYHUZHftm6Nl+T6IqFbC7f8agaYD/c6zELYoKXgMNiDViXU5Psi
IkbnjRgTTAc24lE3L0q4iG+glTSQlwLyEgZ2cnSMj3WTxcDxp8JA9+vx7D2BPcmZMwmt6mBtGk08
kC7CAZBqC0By7tkWwz7K41WT1g0RVPpP3grnbjMGWNt+Tbs80BZw78dCgiVZUyyWOvcRN7kqqx37
t/FdtAUlYFb59woDYx1St5CUP/OcT8hawtg/e4B5CrEHh+84FFk2kCCgqSOukvOhq/0KZQiI76oR
8POPIX6amJiKvDj8bLx/Ggq3SlkJK9M8yl5nNL8GMaL1UOrziTR1e8R7l5Bjc8na4VTfZjhfRL0d
o82Xd7sQbk3Ly798fzP7H7ZWwcg6v8WMRRhJ3o8VBG9441RuGCvaTSQ9V2ktXMWqorwXmd9W4Rh5
XguLUpVz5zaRIegmZ0Q/i0JJtm7jJxNYad6wmao5ae3PDN6eNst4FnTWjPLNui6EXiylAyuh0xsM
GIJrwXRBu3tPTVOa8UoAcC1PTytalYcAcLfq2L1+7dlDdIs0cQ+7fZCzhyRl+eFYYp4yws8Arjfl
uqO44P80Va2jmXJCK56gW+J6u1frcDwlF3pT87njtQD9X9VB2o+CynxiTQmH1UpDU1u8PV7l8RAM
vYGldQwa5HyU3BJqVA7ctCkxzQ9Kzff5PvPrtkB2+gjztfSI6bpttVKfQ3r0FBaLAVDURxhs50hA
mceg1lwo9SUYSXo4r472hMIsnyewfIBOt75FbglsI9n9QafuXuFt0y2XvYMnXCvN6lir3pqumZtq
hTNyAKxfdvIAK4j/IX2XiipmnUuRZ73b+0co11MsXJisnEQjH8r3ze4p9jAe047n9ntc20su3KwW
/xIQF+685S99GYUTsxMajjwOEtBKbe7eU+pIiFMNFAv6yYSJYKY/jr/b6KNxVuX5YoKHJu7Za4nM
APo5T4c+i2fWV7TKjwLCrNjhI+mnH8QkXaaRyL0zEuGO34sIy0nvHpKG1sXX/eZXCzksdk7SmqFV
NyTGUNmPARMX9F9n2TDgBbHdRcnmY0A18fmfyqEZWi4xSC5ieBPFFXBiMfZ/oH0kwgwJav9+95Vz
iCfZ1OpfLqe8CnGpHNb1C4LA33BsRp9xNjUVviuAYLtLr5q+EN/nbV2hii48GhGYdeSu1xJM5g9O
23G+iKU/s2pfAMulaA2GJLg6AFlCmpEYNiSsR1WfOzbz/N5gGFrQMXDnqgBvb+i6i7wAxRtiURX9
G6kbtXMUQqX6ErPrSOT6WA1wHhraq142WeGCNGgg2qSbu10nnfjVS9mLnvz8YMC23FddOUNr4r4+
Q3wwecwI0Gsbwhe2Gt3IGdPw5GroXCuLOlckOaAtaSGSE+ORTNYYPOSHukrJf/oD5Mzdrbr+6GIc
f8EJpA5hrwsCBYsjNd203OtfZu3mV3NV+rZwAwxPRodoWw9HfWwCfyx1wX/q+pLsK6Rzakxdr1X6
YjQdBWnyzrPNh30D29txqdNTMbiS1YrGlpVw3xxJOZPpi2N/xwXqhXiDTWumrGRzTsfLEk6ucOpD
9coFbF4fdJLtz82XbqfvceZZGEv7VAxcpLSIsj8gJtsK7lBAXIIV3vtrJp3j/HB5T04ggg3ntyC5
BUdi+5GQZcW/C9BGJ+y9w+KFQRRWrZz3BT4UY82m5sgacxvb2wFu3ywChECj1bWJokRRJ4lM3p0S
EUsla9yNEfenk4s1Gp8l4cqsxYEaJ1rQXW7hX8NON0bdS2DJ4FK41hiNSkS2BF4YuGSCtyy18qrB
bcOuyS/WJkEa/gubdLg32gOlUGpVkOlJvYkvd1sQoFGjW49oylXohwEXAN2jihMPnXHI9C650cRb
bIdez8r3gw3KnrlFi8yjuiXk/sZ8nRao0qgbh+6q6BXQMNpTE881VBU4dyxIbxZZb7U6urxS8wID
8Tx3bd9IUH9KUEd+2xF4BLJII0ICOc7DLqJ3umfaWhsq+/So76Go9mFEEmIWunp3lzy0QH2k6ULK
qXhRzM9vYTv3Swh1Go4yWBHqniImvIK+OKIQWo+T6pOs6OWvgrGpkw80D7cenMNO1qfTJ1Q7ll1g
gOQ8oRiukmwgTRUXVjGwQmPwspRMB6dDKkwmuy0cpm8gnaZz2G7W2a8Zz2oeFuBk37L7DlxuFQye
m7FqfsYsLS1T5xQR0rSXrgvdo0xENBu5CK85SjxxMbAJ0kyLwW4GtfCsFXLhb/5CCj34g/EQYtq3
5uyuwtpDTe0MLYBeJvwe+JYokEOEjDMI34eV/PDwJbhRi6Dl7Kug5Dml2rokNQQgSPXlETt/OFHr
oA34gVEmJzkX6UBEcwWwHmiUVlTFKwVsPFpIS2Dq0Z0BSwq2GycJ/VxlIvLxqNuVLDV4NCncd+7H
ZiBL+Y1zp6nxhoQbbrEYaFbZBKihJ54UVxcl81zklyx2CQWp75sXTXJxrdqbVrINbz1YitGFLAtK
yV6khIiFu1rPf1VBVVzSsxGaKqoIHAZPCOPK59KxRs/wKuztlnc0Hi9xHzp9Qu2G0wT4x6mWt5mC
VOjYkVp6FU0vd4OmSDXdoekDBkjkEAIkDMkuwvRhKFpy4iIxKlF/zPo8xT4JhlRq86uBHe5joGIA
Fxpf9wh1WXuIl20WXhGfJxsAMj3BuP1bzXyS3lqCoISnSwAz1JUaz9eaIBnKoK0UCGxB3Nme2WLo
RyNcUZFD4zzuLB8c+R6eaUJ5Kv+SjM9HzKAP8AVWJuMfC/F+n+1YEEUiiKUJg4sXY+1iArlr6t42
Iy18EVXrsBEQo9tbYh3HTMioRopjXwEntrpoQAnjbIiIOzkYX+hxcAMto7pi5om/2jqVNso+KagO
bdPWtr7xrMPyrurRyiQfAF4OsOVyYwOIm6YYgah3ocjT0RpD+Jm7fTdbpFinnveMcQvu+YUMOguP
TrC97v3kBf6esHCjI4rQ5tG9Gvi7g+xQRvj84IXNzkNsbJ+TNDCjdC/8CQmpHkkA/lv0+VGQL4hd
uOSXY/56XQklnqI2BdQWaR2gtDKw6dN/PpA1Gho5Wng3De59uZuVKKZ2JbYz8XrpPrtc8IsC1rLH
ZqESb+LrhIQutzJ8OdmeGM/PeGfB/KZe8zWOy+69MCVFjrwyJIAo7AeQjKJ+c21VzMY7ag3sWkAd
9cP+uP6pjSUilEAGpGn+QEGJ9TpEP3/0DPuNSm4oevFwKDW98Wgz6N8z1tiWOGVZw5Myll4SnvCH
VieBbVNP0i3jlGfm3c/xRQs/zrmj8rFSxCr5kYb6ZgqtPtpPw2OgACBvEQONzMqmgiPgiwReO5R8
POiwjLKXnqju+g7A3nqVTW0PTdqnTsb9IidTwbB1EIgi4QGU3++qIRURJm9AOf2bHmhq1/4B0I+b
h4mlDADKDQaZWOdxzWGE8Pz+0POmRvr2v8se9msHBeeNHojhmETrdIN7lcnlEWA0chpycvVgUIBq
Iay2hY7WowQlAQWCgop1oMRP/XTEg5JoeqNt32SSAjvVo+AFkKeBFSATAZ1F6dZUXKj+n7qZBz97
Uuyk1n0yc3x0dPoxeRJ4GWuqexcdxDfPfI1nN4rMzE2GpiM7cOeNXMfPX4N+LcBhlU7s38AgE5pI
5mfIcHk68c4lZfxmoxsu/HronacmKQ70cgmwF+wYucYuFGPD/wBNECqOfkqQ7/y9B/7tm0VhPc/q
vhgJIt+1GusRfO6xMR8cE00oMnGbMLNKyL7l0LgnOj/qE37bHEkvi9l0keVBOU3qJOHOY098kDzZ
7SrzepJy68XpkTljuVRIwFppyUnsXM1S4RHcE8+lpiJiYH2lpSkiQdr/tnC9/74WAA3kVvDgYIWB
KQ0TvpGtWHPVTA9sxLCJAGASdrs8WY72BZffIY8U9cEfBbDqKDAZVSRAUKJRzX9wKfEZV6nbjlCI
JMJAgHJZoKLRl92sMmIRv+m/1L7OSh3jOYpJ+4RwWNCNKqKAUfdV+OFQDNZMbEr3X6lAxUjk0eNb
Q+wAJi+u+rdNzwMuHnaEz1f4Q2WGHsc29p4KM6yYjWCvVVke1iltuSoaR6xWUuDgegc5IouPZvQA
68OK6f3IK+n7QotREBhwIm0loMNtpL9ZPknOoqLI2uHeeV8Co6j8Jv0kdtZ7mmFHLWoIXcuJIFeG
iiw8SiT4EYC9fRNGGLoAvRfmUvKtJoS14pJUYMBxEzs6rzcEIjaC6NNUdHYSyaj+dK7QP3MxlyWR
elh21iX0OcISXtUvMqZSxkm/VubD34PqEPFjsKme9m5ohQbCCEOOIQtUeA1Q6br5tZqBui8MOd+A
JMhsp7YVbYbdFmJP5Yxvzmt7yCmoVbDZkHm/bK/pDljWXs7pva6uIMeEMmiUvDJFGsiZY9P+f/kM
yi3CUyGFmPPXnNPvFWnBI4teNehnOF8Ci8i4L16l1IelaUDGsfFF43B/F9nj20w6zuYyCXXt446t
lh9gpQSK4w5OZ1TCPh5/k6+7XxqAtIjhmypfVphnadUPBbY/SNaSHrIiTiiq+X/wjR9sJAn2H3jt
4Tnbaca+ksrvHrKxZb22+nX7gOXf3hfRl4pR+nAyV3GJ2MLz7Ws/7AR56uLvQ3QTKMJbJMfZqVWf
xEdpR0JhAQJrq0QnIcDhA9nHUpslIoh8sfShzucvGqc1DycwKhNIx9yWhQxPo1Fu1yrihnrUUu4x
nYUGUZKWWnwgWCMrpqbFlnHqUpucD9NXeBAgeuS+gBY3qPgjxlTPMUdg0BtZ9NrQlXg223QS9dYa
PYDTvPEAxubHkKNrlSUv5FbImiRutHqIFtrk/LOGA2kImO4Zshjw7Rb+J2XtFVVBbzmWncjZaVcZ
e1QQnZAeLhZZMZkSeJom6xWcYoRnfFdNyIxoLzNp2XgfMqm4AAYHR50El2yQrHcD0nsJHLCzTQO6
arEn9yyRUOUxMTRSgoR1wjg/KS4se8Oic7X/sw5s/rmiRjQAJmmDgzr/WkOtMkmMX69KZ/5uBiuA
n351IJcHxQu4FQeHNSRp7+3xbfwbnWdrUVZcqCCun6DUiAjuKZ1hhi6eGBrKD01MX4M8pN+DKeQ/
vsrMdQZV1EFrCwzo5IdHEdZ/IXFl0UUsAamo5mTiVWzE7wIKxp6H/Adn6eOgbgAlevGLOC5ALEt6
U7tb1acw2n4ordMA21T4A8SXptJuJ8YQgO5lUCLUmIhkstIdpXqLvWZdz1Glzx/uXoaamtEoIiNo
QWRgn7mskbGmlc0Y1bFInfSyC5hY8kxXE1zO0xvHNkuadIicPuhUrhONGpEg29Zl3H9CTTCuX946
S5DdwFFqn7Jrsl53oYjV2jstFmFk8b21HXg1zxz++pygWsQiuP57nTWID1PExIQyFUkdJV8LtUFx
jh2hpENDXLLAAjkkv9gxJ+XImD0XEgGYEcABgN3D7YIbDvR7s/iy/OWdpqcpQ6TDP8dkT2NskB5A
NIPUl8x/BlO/BhL5y2C7XgevQwBbPh/n07uzfKkhpNImvRfpJ0PQxIZpv2fjUG9MYiwgniCCtx4A
6khkh6DUikTdKY7HUqksZcBn6/tQlLiLTj+0DO0JCUsfG/ehNKDT6ksV4lzpPPV3bCcT4ojcTO7O
seuIbra6qTFHzXLxR9ZgHUTCJV8vblF0Fboo1io7keMKWrIWJO0E3KX62uKRQr0fIR8tLrFvXA6r
tD8vM/QY0/9m+8Ov7mY8jOAjh25gJWLcSBHF5Nnwekt1syck0/lrQDfiR7kKNeUixnOtSB0UMTLT
t0stUQcv6MjeRR+zabAbTVeMYbm/ZP2YSHGSNHmDQYW9GXsva6UAWx+52RWviN/0WjNqoIyyTMA+
vngHHn/V9VD+ymrn1Qarpgqmp03L3aAYh15rnNSslbhioXPNlAo1KTU9EuI4ebSA8xOSeS/L31n0
8lmUvBirLOPFm0tX+KFDL2vTDQvbSsJWXHfpVkR888+T0UuDndIhDYqmRtehdaWwRsJvedL97n8B
nkZK+s7qSAnzn5DCVZ99N0q2NBXJRnCm5XFJHqWVzmUzlbvcDk9cd7Q/oHiT4gM+UbsP96pMqRXG
wCN7oCnkyYNe7DaRVHmAQS0iaN/GvPsPoPjkgFiIsYHcD55ezfpNTNNqfcvUrP4sjeRLtUJi5hQn
tTqFkuNB3MaInFLUHW3Y2Sa876QDgQFocizYE1sX2xCE1EYc+i94EymgaI6ffTuUr3urjdIxEMQg
OfFHGcTY/Oa2Tpr/7hNlOx9mQAaXMz+b/Jy0NoECgF6C2ZFTG6b6Wa5LpCWzA9VBwnfjm3S/z79y
7UsSPlWk+H+8lkdwrsUhi7W4Um2yARSF4P6xr7BXhkr9cCYg13YhqrfHLEWDgZoMo0wd8OPZZzaO
yqOgsH5mK0hFGb1JSMgNLw/jMxgqOk5SHb5kF/mZBSZJyL9bZIy19yKQDQMBOg1+f6+oHIP0BmPT
9QWomxGwGifQ7INjTQ5nXgTDkwvu1YYe5wDI5RAZyKd17BQORmM7lja0TrbeSCPwHiyJRzGft50r
ImyS1VXvJv7/6YGYw7fs2hDm41Op5s6l17ywf50K2HmuGNMQ7mMWaG15+1ZQlPd2T0JzpnFSOpuF
X1lhSQhzXo38ouaU54CrepmYbv8EF6eD4D7BkvRV1iZNUPMRB8I5xOp74nliKGl6he/mBuvTYm8d
Y7uDhFvhb86RPdusVfy6vG4NT5Djgd6EX/VlU9c30rpoIRNGODYenPJDv8o8q6rfbIhdNRXXq9k+
fXcHMZ8ChBnDhB+YQ+v4TCCHqY/c3x2PIJp0tANuQ/m2DbB8AfXccWdWnMSU/LEaa/x8zZ/JrHMV
+Oik/2J4OnrGftuaPb9K2aLbB5TwFatZaHPI1Q7oEH0wdpSxNnJLi9og8tCN96RLJg6QVmV9qH/i
RIfYye4/dWyZXEMCTDj9dnNkrZBZcGcOuzuP4xulZo4xW3FRH0b6lO4MleCcMPSE3Rar49LUdjrZ
9qLKczAxhyUBdlFUyOSnVOK6uq+gVyVqRTMpxbptI/bJEooZBzTNZF1DSmetAB/pAJbM2qDv5Lhg
Hy7ovMquE2BAaP7ZA6cKCdmKjqF/nQUwKwiskP2DI/7Rze6jXbokncjsp4zxNyTNrPWxaVMxH9jC
vkENSr4d7iR+x5eTM9JCMT00bQvEhGyXbgUfyO4WO/psmEOuF5arEGWpkXpV0tfMzeOWd9X9/8lm
Ib+YXFdfFSoPsIKY8sr7yhrz3yyrSWrqd/7p8rO3D4H3w2MF5R/kye/2NRDLxgYtT9kGWYJJ1IHX
tCjf8xfdJnWgIOWAi5j2xZaZ6aynKi+PaMWojOWZL7J8IzQIr/8eLaBrGltm/QIO7YH+vtHlVxGA
5atuLmt71UnIEb0WaWvdfQCN4mnvbZquJKUEfNj9J9TqyYupvG2wOU+Q6jfwwRK10X8xmoAHIvo2
ggxHcqHj6V4zSWpoxviGdU162CjmSjMbsVV3iaLAx0rsFC/2ajBMMIz2abw4t3GNfngKZcN1H1kf
rYcxdvlEzDaLrWXor3zUGlKQj5hdKP6W38K96/l3fqLZJCUYjhgSDkKCk2J7ovciuY2JCtCHTSMA
xzjDqOaNPyCz1cGMi3X3yNgaUZoxn72+9LrrkUoVaLys8dTQK0q7Pdq2rAaAGVpvXe7rkpc2imPN
k4V77r+DUpTcg1JNQJ8FdkaXPatDVihqJVDpj8b8Vuv7NBnmCuBEd0YRwNyRfpyioU1A/uAEE/xP
+/9SutgaQah+AXtcgNX+V8rFO3RsQaylz5IAFb7rvjDi/7YAxgmjkDtN4U6immu1bqr1BQngqami
tQJd84LmuPV5OCVvQN0NjnAoc2qwCUEJPGDT11POdHXVbigjtpMdbK+Mgvq7WnxbpBkwjTnL3AaO
k+X3w04u0aS378ZGTKpUlYp36phhmweXOkzzzd9qD7ZI02PjT+zpjtO/6f9rAQ/6K7VGBL9MO5Jz
hcgaUD11mVOFkDvElsh/AHduaPLlgWWT1Y3YikwgYGaJrZgx4St33eMim/wtFmjR6kDiZSpE0atp
TT5WwuipVWkpdiaRa0D0M2EVIi6FJJWNpzr2YvGKxyrt3IFdIZ0QgJJALUaLPTVs81fc0goF9j0g
M1YdvzRfW9mVv2EvKfaTaxpO3TbJ9rk0R66/hPdy+70iDApH/es3aASqjhDbrD0zPAEHX4U7b4s1
/X5HerMQeQJKNQnMvOwM43WxKguvLBQxG+e/YnLBSeadN5l2Bsdcbh5xEyFBbmAfmuXprG45Yih8
D+pCtGQHo2NjwRjE4zls2qjZZt4cBDJRQPBFioB8b9WZHzPy1bqbhRshIJcpR34cLRQBDRUOglBt
abVAbvZQ0i2tr39/pgMT4ffMfUDpmO68sooU51KGxqj20sGodXkq0UHrQSZeJdJAa2l7GNal605K
oq1X0jTwDlfkXqH9rZSw3Va3Jy9rykR5H1qHjJzj2dDfSitNFQhpB2BW8aqO8TyNjZ/RTwbAW+8J
45jKP+KbJbpyzWyVQAwus2plB33yv28+tvZC9iRHQRyKTao2P/lYe7PpxNmtAAbzDEjDeH58y1Af
qbPWx3ZIWfARHXH8/a1jIA9qPL7u7k9y8f3A307FnfZgwD+fg4CsN1r2DggDh0WpGlHe4cF8sU9m
RjUKjEj3OQD5i572lUfHGjG/7IW3AZMCganZuKW9Zk9AFBCvPZFmBzigsXbBnc/3R+qVOlYqeI/A
PdHFlY/gWIonB9TtCgONMP498qtfmSk1BRGt7usgSRspL1P5MaIoVAusJwpYfH5Yp8So1VwbpeE5
seTmzFu6YeElhwT3BbXXgcBqs3Tg7eDt+hU0uXuk4KE/Yf/5SxypxeSFspNVBRt9mBDes4zs5Gdp
iJHAh8XAr+yghUq5iydp/gmq5fKW5EPODL54P+b1faStnkgozymWIys7klvIEda9MIir0qnDQZh1
9dxV7/xldjzRN0duuWGQX0bQkGzUU3E/vsgua2RwEY2CO71I3Zz4qQksaQFYODFURwA1JBg7mpf7
32zrg9pBtR0mLh+304fAWSlDeaKs6hWd2wLIORtKVNNpsACA57tWMHpeK8jxMECygIxbdndJXSmf
JB6O7nFw+j09Cm5T2t9//JS9GqJrgXAR7ZV7UiqZdzqDLbZ5HYsyMLwW8uOv8W8dAAhCyfFz478z
b0t/VmHkhBk9/H62ltpb1pQlGEYu3SU3hlJlxsvzcSqEfdYuqsW+xvbLiL1xHjpdZPEnSAdfoR+T
HOFz+w0q1itL6iap2y87TnK6t0CE1OFw6uCpdIR8kuySDnArbEtgCrgWoksybFWkjJo1J3Uyd5tT
azg6a+VjDX6yBDuvffMSHjv9TdTGLpTzIsFR/DayOzSD7TVRjL2BlzHVbU0Ks5nkVf10lUpRLL40
Zxc5CDPEQ2bdWAZBBLujM/b4c2x9z1lataX89GdWKYmOujdGGhN9IYvfE3tHzMyABqJy2Tm/Xec9
THTptt6cmLMyeaaX7IIG1Jx0Qild/3YI2BQ2DfhlHzr92ylTG/xFEDGxqGLxv3pDM2bYrb4nqLgt
InxCFJUXw5ImsjOzVit8u0YgjLgZKWTeZv9s34RvSlTiZI/LY2z8JpD3HPw1ZSs6lLENlblwCVJ0
50GN7UTZo+8Vt15isU6M2u11YfB1Z5TrPZvTyZa1xVzTbFQUN8rmXLaf558ViJWtMnk5QzWUoPA0
WLadiwi1Z2If+UQg4b7e0nJraMTHJjho1ln8qakKgfg8Wz4Xvd9g+/9Dp2ccdZpHtwQOcd6XFh4Z
eGFecweEp4Z9QNz5aDDogZ+br8BnONZNe4CHNNfmlLGiJmmYpYCW+/hP4eZLxJrhUXWPgH4G1pNL
F0qeDKQEZpSalTYy7frdof2aCCdDXwe+Dj2WHSkPrPJ7WBu8iBsU0+njRqvpeqfvik4IUByPc2CG
58CN2XxCkxlq5iGZwQv+trQFS5ZMtyaEo84wN35dDj0u1UFpmbjZZ0Fy92S2MH0Gu1xGnpeN8Nw8
klA23uSYm2vv4yvsxJvgKUcjrQfVbob4IKDcHHR5+x2OfgmfkorFFPc8l6KEkG2inPu59Sg3Uzvw
sfwYnRWijtvnjW2vILUNSwhlow9bmZFql+tn60Ro+u2qHFZB2Rsx2jr9hTLwKlRVLkY+VlPpYo0T
ZI0XykUj6QRb7anIdD2ozvXHJs8LpPPsEOK1E6M9oAficE6HHn/AYpQV3RA9I89+oBCTEMA+TCrz
ta3n/DeM8fIZj3roH1yiuXZ787owunIw3joHvreIEjEHPw0m2bCmUEPd+vcO7x/avneGe/4bIvcS
hvw+nYSwud4X0E9lJeBwOn+UV1pH5bvD848bGHyS70kdOKKNhSzIk5Q8j/SuD3SJMv3arL8+d+kG
ZQUE4BjlE2MQZhz2TPpVfAbBUuDDo+OS783YoV2yJMaeeAP+HsBapmJoJj6fwTIRPKSYwJKnjiPe
h2eCgw3Jpnke5crCUv7t1dFx/FQVANF95wakAAoM74oep+PWmmVJeEZCkAluhWXPuBZKzcNnPf5H
q1Mq8+LMINHFdEoaXC3E6W0ZlGhzAevZ8anBbcCxfTfj4kSwJAX12q5ZBejz6i2ozCWvVtYA+cod
bQBmfCg+vdE46U5GUtVJMdkNXYJU/7qg1ou1MT3CetTfLDn7432MZA1BYQ645dzhKatXjHnhH92c
eqEYBmu1vu6GQXwoHyRCXcBFy+olb9xERzKo7braZ7pzgcMvtzm5weKmTmGMZfXPNNCzp2Jx71EB
1lb4JHq91hdzDmVLlzs6xwOzprAp6+saeQyHCX3puLWWLoU4GWv3kvcIY+0Gko/qFvB++bwMNDak
Bc+BCTGIMTWNM50K7QHJC1aBFJybgSAdOxVgrNvXGrI9+bBIxxM/bIMUjyvRZct3KNwEJLzAjozW
N51pgxHb6VzMsVc+SJ4jWhLH4wc564sBEDtQrFCEyz3JCUPWvsScmvYll2LsQYO9mk4y96UV/CMI
vxU6kTlFSraHBqRPHhs/64ZAxIBmeNPeq1BD2KyRGLwv3Bxm3p3CpDREGqRkyJFZ8F5OupUERD/V
/BzUBotGBvoVnPWeSKVRyrgNk2r5R3AYpfXnXVBy0Dg2Mcq2nk2o7L43SutDsfL4aS24KawNYAgq
toSr9LIgzBxYRiarAf5f8n6a0b8biHz6RovQIbQ9Cm7pE7YSBRVHtr5Ny2zsS5n3UT+kNXZoBTXO
GZVehhiuqALQj2GtY4n52AjWrgHWHWMET7uGznXVEO9X+I2Y1l1akb5WARWihfNXdeW/PjLI25Mn
rV7TzjIohPiyMrZyt5U+QStqEoj6GJQGxzu/9TlQPHOHQOaU/zNIFCtSWpwGnAjLyT3vKw5eTnxQ
fJ4OKs7zf9DvH/Sjq1LZ+yUSRiZXJLJ/jzREZ37gO70/jMdOtZrcdb4ZJ2FrFeneJBOkTVGdscb0
CqziiprtxaaTnRl0B5blAQW160nvZIifl6q/VwTHs1SWgWW+MKorks+iNqQXc8Wo4HXINy3cgR5t
rewHOE5vWk+KzyFDrThRwNHi/TNbZ6ote461/5Oc0LbQckYHAfurRFa0FMyLd8kUJN/DMrvVoG4g
kchtlk1FKLXhuFz1JwvbNiQPpq+GKeVuxl9UEB6Ux7eerYaebm8FPSWTrcuul9vJX+RGhrdzCTm8
oRzywZQ10pHIvbB0y8hR4Gy6cjxO37oZMhZxdaA2G8jqymQkaJMJmkQwEpt4YW3J9sVaKncTrAai
9Mhk15ALCvTEWSOTfwqB+a1UNULNoQFgPvenSIlxilUbZ8Tcd2iIJZ1EmgC0d61WSGxfIbUoEULy
zPX8B1nJbargtU05gdoyuasj7JXhhW2I3ZiP0b42VG+r6RSE/Qd3bztbPc5qkJwBNB7BQ5sGEsD5
AuwFjDMxewpW+3AT6cwohkuC+aeRpwHj6CKAn+9S7kiC3cF2rBVArBkOB3fIpx7W052dwPhP/XTH
TZdOiwGzgqzvzc0r0J3EGd6fGYp2w3rBGNk7VU/DY5W1OaquJOf6Mon6F60XFxKj7SSqU5HZATwZ
seTZ/o45ec4LgOgkcyBIDp3ab3WFwbcWzpOi0ciKCe5uIeKwoHcjH6yJX4lxpo1fbpaMYiMLCoLw
zJ8U5+0/Lk1gSgvpxJbede74um7dKloGGqC6uJI0lfutlH2r3WyJ723+HM6MsRxWm0ia3y3b7vNf
4+F8QVM8EMYltBTXQJWxildnN3Hnph/chVZt1YrXU5ClpPZmyAeubFuGXcegPMHtfC8OZI4lC1ng
eRPb4CbwoBb12Dd2OR+z3DfgZ+8BmfRjruYqcCKEndUyMLfuc+KCRQPwrRgswsKwuZJklXm5Rnph
ekeTqw0VSX1TkzCIQRsy2nF1K7TuRmwIhadBpy859xf7TKuNJbnDjOV0pG9FH9k84zfZ/I5W4HVh
srayH51jY7SVl51GKdgwRx4C0CW1O0U2QbTMR/X3GPUd1CFPMyFQ2+7HXnB6H/ahyOe4QqqNmt2H
7t6VhnHGKBzhvV5wKG+S8XC0HEiJKjLDQLjs+jIzeaaR/iO2VzC/bZPgxSnI+q0980JuySX1yMae
kcmCGMZqwP10Wo2Zm6WoPwcjHRKJk0lL7bg1sSQqFboR3xIf0NvrOsWBb+4yHX8WyGijxd/yQ5VC
JbatJnGecwlYWAhtQ1uaSNPlAOoSJrEqdEAVOf1MOIcxl9flUIe8m7bxOV2pQ6dBjS2lOIZu4ZRg
WF3ygCsnjuoW1OpMxrTX/q7IH8zZlXi6dGHKyxWWTGbUcFDHZp8SwtUcRJxxExbG09E+fl/vCfSW
NC+XwonXi8Bz+6B7x/89pLYP78apHok2CgfP8VmwF8yLDCCYqJplOX3YLi/uricwUkqeeH9vpZu8
p8V5WS2YxgZ+wBd1lpZjzmhCu34IUATUaVRNms/kxNQthcvpPQT7Fvxvl8EhE4nHBOody4UzHW5T
ccOphdVzUz0KWS3u5Ru7f7V7PyBOvSN81mGnxknDJZYNoqbsEEmbnkQllG4Sp6ZPmwnyb/PoUaVW
b4lqm/k8sUfXsx6aZOAzdM9c3FM8xZMQ14+YJQBLwr5GX6m+tLprOO/fjVOtNAu2J674yy41DSjn
y/eZ/YX8qbpsGI35uqGMjPBYfOS87cFCxRU1982MXFmdRTVjSRic3UpGCWhqOmLsE+HLB+90Pxcy
cSwE6oM00veMapOyXE/ubnIeBCwy7zPdDiBSEinsO7Ch8jK2t2fCbCg+v6+AFaw3HVdyqNdpYJne
/+tA5mh7iVED1yOjI5UYuWj9MKJROkXqZanfA3hWtrYNwz5HXH0B7UmX9naLBqsrWYZ/S2wn9KD1
Fsfh39jq1HbH8UGvovpMzuux9QXb5xsflgBFMk2CQDssIrnRs0a7VOwUKq3xOqu96j6cT4UP6M+0
jWFhGZRRYyRWRJ8ZoKvhxGhvg7FHfDU0iNG0bRX0zJOxq/XpLCxQ2vfnrjXec9O5NN++ctXmDwno
PoBONl7SPYNuljUiCGU9qFnv5XBF48uC0IPzlEI1Wxpw1NBUjXQtEibqnMa17LBGenYTVCkCACib
v3VXrEoN8R5c/psN57Nbbb3rCL4lI84qqHv0vwqhb3AmuQf4DESnODQQ/r6Glb4btthWhSgqEDhW
OdvkKWusmCzVG9B0IWiJfsI4T62Pm4WuXVl+HvEnDhlgtXxiCrlAQuCVGXIoyhXfzH8HMp9/EArT
9ih9U+6LWbuRa1YWfT0Tm/pzfQ4Q7DYGo7XXXXWQQuBMix62PmoPk21qqfjbq9gsGeJF3G+tyi2d
cBYQQEfbneAwa4rQeBcDQ4N37DFPljQIBKI1AQxJyh6r8XQjrZ3rI93H/0/Bpi8Y1FPFUTuueE8D
zo6luM4K/cmSOMfKr2/+ih82NB2zsbBAz5710vqs5T3gPAyA/iwNckIZaVgGGiIWWSaZHoYTfT8u
89AJZUNXE5+dN7xrwtiduFEjuhMh+CgZQVxr2l8hAV6MneD1mVjpHoEyUdER/Dml5igAFioqiMbq
p7KbFiZTsZGh11NmnLWHCKipk4KWwYgfuGQY3aEcQWL2dY/jmSqfHKJ9TxwCd/ZexHnhPEAKROlk
D92m11Jg6GpAAMZbn8SJ+Ul5Npk7Uz0jqbbQKVbKU9Ml0/br47QIHT/Ijfm24Aya+I2CgctS/eI3
7Kc4whLVfE28kB7lXFpCunxiUnqOg6Oh+RDm/R50c+89tSQRHumOvvD3Q8/PhZrSNXhuiFsh1Wbs
Ygm5AzMjg4gau7eh47EZ2UFwU2hivhDFb6WKrmTbWWtA73DgbdTNE5UF2/etBPsYdA9nb1RikLzQ
U5JKpQGcmA0ucLbKFl0Hnh94oLr6OE0dtUH9Jy3ZaW0TpNapCzpY2XF/qlaaBgNe6YVdZh8DXcRu
SXyQsf8nJKetNZVW3ymXaAA9hN8TRAKmQ3S3d7DfEfStp3phbmjYBQYdxo91scKVCAPdS9nDVkaW
uw4nLNrjqsWNabxZxOCNUgIBS4K/+cidjQWZc7d2sCUf6VKAopPFjfK7cFdmqCXIWoCnAXrk4a2z
b1VfxNlWHTHMQ9D+xv5r4RKaIqZZol+QkjRftWeMxCPg4DLdZVHdU/ZRBw+Wb22RsRSxTAPB1xcT
9hjwm8gbxoaoPmWHS3mnNbyXeHEah/Jwodv+A/l3dqGr/1I2t7+zB2nlHXsJ5QLoNRxfC4c3zyuH
aJwvrYSkgZnT67bCKC9F3gPesjQ/HsuJQPRI0e1nEMb8frrvqF+tBeOTR5x1LqzoCBs9CHRXgJn1
Hb7yKyDswlCJ5tP877vfLBZIwH+ghC3mAkIPsOv2u9FR8iU8uyXa9Yjrr3a3qSmnmEuMW0dofMn9
iZHRvSR9eiYWF25b/yqE+I6js2LySb3b78i1U5ncD/eJpASbuwRY/NdNjbXvuEoY4/yQu/2tIhAE
RuPkg6i4BxYPooBEDeGzMyV0GsbvIOq38WBQxUwyyf0kv/NBpoKh08vNG37Ur/c/V+ch1ERiqOQy
mRvsAxkWfBPRqW5jaMXgieP4q2GwQmctLVWB8LkQxiptvquma3w6Oz861Y7sHdexYBn+n8Aapq/B
/oZpaudex0Fp5E+/Jn9WQH8w8cNt84pRERqpziJf0J7YlQU8I3115sZt2NR5qhUAXGQ0s4t8f97n
+j4IAynkFowBSOmBFikCoPgV9uCF858gl2wA4hl4UFfGT5ktZFVVUU5AO9JOS/7GQp0RB3tkDKqA
4Hw0jfnsDnN1DCQCR4qo+wp+1TVvrjojQ6OTb9uCSLECjIcHj0zXman8rizkxCjCdTrxfCohSwGb
VU+/QXarOewPOgF1TLcrV2CF4civHuSteedm/AfwxqhBorZSdZsvjJBZRg02DE8dRob/LRqA4fAe
DpelkBEANw5v84ItYa853gNOZypTFPse6A0DbohzAIUvg+1sZ3LTVPkO6wdKNwb+ZCwWCqOXeuX8
pLfcJ2TUoEohRQSDYEhGGKMAnHQe5/ZB3gTLxTTavTKdgu0slTAynH+NovdgeIlY4lKuwHhxP6Py
9ZSmDERVLsNaSbm/u53VD/cCdGRGM2lXslzhC4TnD8OldWBHATLouuBC1eIo8XFU3PLOplL+UEo0
JHv12VSrToSILXRM+Ua0KBqHxbMAnLujxgheZym70e9zr+Icfzs1Dkxvcz0y6X7U/xzizXPCLyLf
TF1AYTWm5GU1ZN2nBl+jnoT6lZmkF5oilx9YVvh+aDPonBb8panElxsNJQoKDa0fxzkVPXdYUtos
EB6aHHJqu+6Onbwe3c853mpIrm06u3ESVRNzxGKrDFxVcwJGPUJQjmMTx/c7U2x9hGTGKTXmSpZe
7n9XhBUAXG7lTr6RtvdQilHNkmN23T76m9pLMLlqcnnmsiA9m1/7noKSd4LbwBeuM/Hoog41HXAL
GGpVX+FWT5ETWOpgNfdkY+tjvGLu+KA73wolrXBFW+La91/ozjUz7kWevRMxtioOysAJwhvgfOvH
8Tigc3qo9BdjBXJkJK4mMbi/31ydQomjOhDrLXNHOiEB8scSlZbeahpeSnXfG7ZLmG9BbBQgfXRh
Qsza4cB0nY0Fm3EGqOYnKJ4EseGqj8xLTu1fftpBBv/SVbjw9o7dNP9kHs7uC5a8pNgw0CoMpzEb
vP1cYJiRQTESlq4PEjv1uNU4/Ns4vopf8I1USQwsqmiYfyh381PJY0gMW4yFZte7ASn2NiuPT+Oq
rGWKSSGFh0S8qYxivGkPlTD5hTY4PCLqp7zWkwJ4sSMhoepz61uV/wuKL4Aypd1o2m7AW1EPDKVS
ZvwfICv8lp4eQ723UmaYJQEan7BMeW7uQlxe4ejpwsK5Mek6e/xl2uspncdaX7PQvExQ7PXudIFX
VPS7plQgcydezxAWxy0GQpNduC1a5C7EotWdTFn1v/REbeDLBqyDYrZHxEwazNpqo2R8sfXlPHX7
xpibvqpkToGvXaDjWQGPxGNS6CinQaYsKHnG5HCIy6esTE9BFqj34XAbVR4XoROeSHZEBp505111
6RhxJEImrTDmeGTGJAzyeIERnsWpmLWrtkd5NmihHeFjKsx2Wb+fLaN/DuJ/ruU6J8Wnd8pdM7WB
8soxsBqLHUack2UpPyA2FB1eStfDnc4dD7WZYv07CBuzC9/QmatkwBy5ehGxx//l2THmw6Ykk99f
hH0ZhvYpRZbjEmS0hP5YpOIZS2dJ1tUzX6sjMrWPpoOPN53bIjpQnFCU+9ur9S/vH3EYMk7kjwx/
bpaZsTUW9j8R0l6xvPGzJyOw3EiycStpfvN7EM6NOIjb0OntkOhHd51OE8AxZyocAvZjPJbVRe7Q
3zKK+0KbTt91fMs3bFQ5pWSglVstnlpbr4gMhZITzxCUk6pgBWchaaJgJ7e9eGWDaQlv4efwcRSB
KPLBZCEHfX59D2nzM2LNX1BehQ68w0tBiEeI954U1EYavqjpNaI/gyPp33uCIEze45yanOyEgabh
qiqDwRNtFytaYePJFVmk6N2H1KtVyeQ/faSI8BUYXX0seHZn+8Up9dbUxkQlZMpwK7KxQofQcp11
cVjKkvtLIdOWwVmlsi8h5cQPfXTVlqPFoCpFuK+9jhQs1wdteGe+XhK6P6wT
`protect end_protected

