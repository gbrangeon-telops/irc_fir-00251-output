

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
J8nZtW1Q/IGk5bZ13EIEEDntauAKqOlRji4Tz7aOFZMrRrl3qAAP4lw8839dxHbOPehATkI5mWRu
O3oQzXKv+Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PO3vY49rlamMYJ9pWAsIelQmo4roKT2hFecsbIIwc9Ce9j1Gil9MEDKbHqn/9XWL2CZb1+nggmfu
MhGokjjD0xhuA7bkrZ61EFG47AtPbrzrGJmyawEAJ1PNLVKIspuVYNxaD9rI6pyGoENRti8P0hyl
/TLRO8J/SzWO1wVCE+o=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lek8GlHbeyFgFk70bzers4fkqEzZWIlCFJLfSucq9OzFI+lvPoCv9lLJF6jbu+G/Gu5TV4ZuNXdu
mi0r5LAo17AD7VicMD+MhRKb3DE2N3pAEqyDrMS1jasKAHiVpH3eXVPN2AI+lDAVZoDhvjSuQjfy
us+5QMijcCxvAveyXwnL06kT9i9dtQ6hie8/MMqHXkiG7OYqxKm0Iia9+F6bzSI9YxeA8Doz1sM1
HWlzlbYLDBCHp8//PX7kMS2bPsw5C6UPaQ+TKox3agXXgpP4ea6EVU3GCBe7nIo37nZIVwI8YFKU
1lK2hwoX/DoWAQ9zzkBtnp8rOkj66EFG574xNw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H24CFb/lxJKnebrcZ74EB0cwdvz2M6JUcau88JBt2iuFL0aDDA6OprhhTeP6OvCciaaGRsBEok+U
cbANkg9G0zLP53/WvEkpdYtezlQI3mkakzT3UxyQr7e+pL5MFVi19R/4mD0m4WBOiVFQ4vPfnILO
XObce3WQbGcK+NGRsMw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RFnK9ETQkPWYtdMW+yKQ1MaijPhYXOMfuPVBKnsFVaRScaR6M3W3RRHlGeNOaiw0ukl3q+66K1rC
RHUWrifpwoSOSO54nuXmCv6joF0+cR+UF1LUkBtOigSpmJUx9SscdsvDcBNzrLmtogpoKRScYdGy
LrKeBNVoMEblduWARlt0XQCFRD4X03OLybCK5/hlbwAJA/OXY8QP1rB1MFXLkjS4zFm16T1j7dVB
psuynNAT4Rwsqrw26xpeXem+8Ft+gBzXVIL10rNKj0y4I07ITYInhk/p/CsNH9FgAhYM9jsWml7/
R3A8DckKe32XlGviTUqdr3zXyrsrjZFSJ1kTGQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 107936)
`protect data_block
pOymsE1uTxv33dYOACqqwLVWpq06mBDRzZcBsCONVFrBB6rAmYlZgAa3uJyjkeVJY1gy4LX/Oeex
fHtz1ov3sXUxCfJiB5/li2bUvcyzGNvGjfn+TtGSNWJbesJ+jlrk656KWxlEjTju6bzeX5RereBo
wAQ/edsHC46i50DIgCgvVR8pPJ/p1HTW1trmALLNDDJ6ddeK61tQIwg4kiRoJ1873YCoqshKfs1T
Lb6ynWK8Nrl3JT7QFGuq3IeqfoFqGAVuQIKJutAi40638ZgXcz8CEDGcBg74lHC6jptVwsSNvGE6
caPwAkQ8UkxTabYYeb/A/PVwBldqhHq7mjFchBwFgKx6so5ggcJBOMaSv0G0sYmm8bU22AKMXNDw
uEe4lT3ev3Rr3ZtbOR3Db4DEg34mSzsY3kN9OvWk0sp39fhpipVvOyoIoNyGnSTfEueMkoDPtWu0
rzFuOXzHc1Z9nDQ7EbR2Fbcq5faKRnMF6xsqrqSmADsgiwG5gtGjHNaen4SyeDtNtecaJ3fUHnoL
tELQx1Ha7WOAdJWGVKQ56h3FpElCIW8spuJnpjEIhASrOOvwVBol6C2I9p+FZI2Ey2vBrsgKbQQZ
cUmvbKWftk2bMlji/Bi09zSuxfMWjoRYQcHn23x4mr/OTB9AKUp588/aYX7hdfTsoyfrkhaAa2bp
U85Ae2LY1s0L8SBgYrqQrBM5SDx3dFc8H7AIXNPL73tWdCPFfFIkqdMvU1ljZqXpq4wlEw+2fiMK
4MHI1mD5pkSJayiivwZQ1xik3+jRHeedevhmsJ3DADnIWqb7LSfBI6Qtlcs4Cul3i6RaKHkT+D2j
CTB1/GmW3BhD8z4/FluRjU+rCMGwKgLvC5XN3w7i9x6uP9g1LQ5ZZN+wN2LAQJOBN94U09WIkQ++
Z5pdecWqXvmIRNx/O9snEqQnaXh2x6+vq/aG6ZPlliQ2qiBYR/mHczvcoHzTyvnkiIhtmGa30IJP
uXexVnJQ6P1NR995VuYo//Z9RQI72lAnW1DWu3TAARywn6GHEypPLYfGHBWsG/G+j8bcQ5nXSlq7
W0xfRKnPJXe9f29VYDIse5pSLQyTe4fI+/JEccELPNo9nL/MXirsGT9E6QiyVaT4+CeezVDtsuZt
J0NRVoZUnUSLXIh5bi9FsIHfpS+yz+XOei7rqqF3UfoUnNpK+8NJLMS2D3qWTL26RKQFVg6tvNH+
xfw+S66P6IM2KM59sJgsJK1lyvhB7LoV9zTyM9QdX6uCv4ZhKjTwV+kr1tfuUdbuMQlLC0UvweUy
TrTx24t13eelQ+w74FWk0tOsyyix0j+eesUVF5tqy0j6SmH+ojgljMct5ym/vCjDMqBLgAmV7kmP
K0DGYVPxOdaDaCuEpRKFOpg9YcpEq5yUnayxzp534tHxkpLaLSiKJB8OQMAeYXuzfCVFGWsBid6Y
QtLsOW8hWGsb/ZUz4WB7Bj1E8s7PuCv5ePk4UECh+7Y722qNJY3QMDDEON+tY8QUUH9mEHC8Hy71
Azm56vfbGFn4Xnvyn2G5JyPW181CBgyechJ1sKTgirF+cq0R/zD7i6nZJFR/LFI6iAm9eUXLMMX2
XIXYEFO/TqRCTZ8Kpv5DGy1hmeV03TLAT35tvRw7eet85sPu5wLl4LLwFF5JDIZCaj1igL96CWtp
TzEsnvBNj/uIKhjVC64PwNXWeOZga3q00BMTo3Vl1rxTQjNZveb3oQi71QpYxdv2diZH+Q0+DB7E
cN3Y/sq+4j3Pgz3PouJ7N+spLkQ/nMmRM/gSctvz9brPdyKj/AWpHH4JTD8a96XUGJ2imaVvOvdv
M8uDvwZ5CNRPr+Qg3BjQbFUFsXyJqHms1T3FMil9gX6fEE2mTtU8o5UK/o60WYbuT855zad0NxyR
W55LDmLnSjM/1xm3K59/O6mVSB+mnznYRHc7s6jqqaii9eRR10r3/5PZ/SpK++0XNcT8Jfstovts
GRw+tHzYNcxtP0sJRHp2bdxErdLeiGAy+3Zmvxj0+gTru9nXHn4WpZcCB9ZN6XbOcgmKS8S3inKT
G5xKVDDRoFUsnjyhKJCFsvm+S/zrSzpnDs95juBDGSKR6zo7AfUk4TmlnGKYsttcdxz8xLs/00fa
3yZRm96qZ36BB8dVq0sAX0HM9TwnUaZyhCW7z8ayaTvd+PzhcI+fAO47hh0R/a2jenbgdMqW0xuj
CaX/U7MPc7gLZSUkySk+v40Xiv/elWrtxiJ7sIkoh/HQMqPGRSvB817C+5qjLupXTJEC8qGIVyOY
O3w7aRse5+yN0XXn0589JnfDeTlzOMAWYO80A98z64LpZ8XH3dQN1dQdEGo/Y63Fznii0uCONp22
A/avQdsjkpw8dYziX6lnDBLjIrH44qcFzZcAp77CAx3sZYJd7EPK5VROL40aZkkbrJD/B0il+YUX
E7on7UtdT+dCOu2yHR2oqV3rjo2JqpgZcOrCBy/gjysW1uyc0Bj/dyW988OgNN8Q3OOZ2tXPia7q
4HeED7v7wsiIU2fNlgI9qyd7jwyrGEEamym9Zyu8Zqd1AMRpWryjc8hKgLKTTiyKNqV3mUSPBj7o
GJX7v+yQn+dWdYCjDdK2gbn4K4FGWSrkXUXAIgWYiLG89DrFwpO+8d2mcCuCcmxBWNv9sOXVKGND
195X+Y/Le/z3dJFOTzA5v7Do3urSxDWfsmiOKdxaHJLiJlIlT8FJBYEjv4sEXHBv1KkfaoSNY19b
g5yeaWkcfNVbpng3okZoGtcqf+edPfX3XBAHIq3r6YeXuul0JzaRw0soxdqdDT1jN1Gb5J6fmCjb
j/iV7PtmnnXM3gGQ9a5tayvEbp9GiTDeq5QxsTQ+Ge11Ja72+V75XZudFwd30YVcTpWOYFc9Nk6i
DBScbpnTsyGi4hRhiBlufwKl4NvlWfsGX3QaVpva1W+464bDhaEWMo5qj/rN/7ZRGRzUb5iNX+eN
KD95EnFaAlYwiN2cvVnKVBaN8msUv6OZG/eDfvDuUrAamzlhniroxBRNwxX+w/VODNRstsW4FPoo
BznMB6yVr21p2VkXoSADkRV2b9uJKFZUDgkfiLb+TwBq2dCb63+o8H0B4ct/E8dYZIJu45WG1TYJ
u98fQadZjE4Ry/rMxSpnt4zZuBQbwR6fA59OU5nXRX9rql8XnQou9U5zpQjyYOedLXqktkYv7kAE
udUYeDahGH4ucZUPgnfCA/S0qLJQtUcjl6vdTwKRrGPnks0bZjP0LkZaxP2D7EnzoDynnbX31C2/
foiTopD0KKGlOdMH5aoUyF6Lwr6fPoxGTu8l5T/eZQwy5hOVTkcJYq77xMcB0ZBRrbl+OGRdY4v5
10oPwJVZ48pt1YyaE33UMainLVbeYuaf94Vi6rICz6inVE9SmB8h+ch5JB+SC/7Hko2N7ZDoxlXf
MEJ5+XS6igoSue7DUdCCWib/1VPPGglzZtTzvk7zhlDYd2kEpSZCT//pYRppPTFuFlTx5MWkBhk2
uSHjmRThhO7mHi9ZXDskg8nhcFL4cr+l436xsXdFPBuXAXh8DrStC+9O3BchH9rt2EFCkSMjzfyz
EqEZHGRGNrsIs/ZZfEFSER8iAGv8YwYsJ2nioEsdFPmDZQH3thr8Gi1gFCQYb+wIKeekQEFYswbZ
oXfpYVJWovv/uY9NgsgY0Qb6qfXQizXvaGb4pER5dCJYwPT6RkLYX/XoHZU8dHb5iFILulPbtJ+P
0Wnb0eidUk+OWJeJjO21RCSwL+a2yqMSxGZrD6+hPngWxrizDOLkCmf+8vxtVDlab7SVc1gDkw+o
JiY870ZSbRBwGxosUV7VowW1WwVcYWF+qALB0+ydN+Jjxucot67CKJ5c/mw5hC7OCT7TsdGuR9bH
+iGS+uPRZeeN0ky9lxa5kFPEyKYDhciLZfFUv6lU/1rfYpDK+4XF1qZ3/0Gfsr1KuIBlTcechzDL
QxzvijNYVMD7W3/H3AZU8XS387fFnM0Dq55xICGMn6bBQ/NUarV7RWEiRcsCmIWBaY0aMj9KG2tM
TmfO8c09lc2fTF590GJKLKy/zdxohz/f6/xbtEzAAKaVQboXB847M18+LVtN9Jg6/kfQjqhoABd6
TYyeBXkJIZEH65xPl4qZyJCDXkFENKGSFZ6g+62bdRqc6324WxtKcSrwItbVbt1lG686t7bZTu/W
bmqTxkq/n4tgUP/G1U4Q3muIT8Ls4GnQX8f1Ojdz+MjKJ6CvjsLNT8g0UsqnBdnK9qx2tudz7vZw
NVvrzdmiVszukWmm6M1QG4z739ibXlMnjy5ZnQbCdRpP8aSeo+9z2LbT46lH4lksp+f41yOP7dif
gVL1T+eQG4J5EoIkuHyjf3osIRcwaAVdXPi3jHgkXMevZ6eoDozALkl+ZFRlya2vldMPiNKJSrFa
HN9KsSSDtKcNr9THMHurAJmc349JNTMMHTo1GcJdu0J4EoeEKHoE1jBZRX8k/1qOd3nqhWH0wy8S
4ES36Mkc/y+nli7+u1PA8a4HYqfOJL1OUtUvfB//GJMcAV2fjOt9iq1BulQ0wJBOOu4Pq0rnfDlO
S0HxISveRzMuRj/qF+Rv3JnGkuzQuGzKrFFnYSM8xDJxwyynYFg5OGP/80K2K3/PT0xytsT8wmYC
2Y8uXJatqWdr0KRfStAVTMXiMsbMBg2MnpK8TEtEm7RSJPhW3+h2tmhO7vm2aCmNJhaz25DdxClz
T2ixBUhL2ThQy9jQZC+b7GHQ9QftI+g0nFze+Txt0rSpq92zj4LAwL/imM+JYkg0KUC5WKd0J8/T
SnsqOtg/ArJIOQO3aRug0izJIL3OFLpum0UyASIEH4GcpC5+daFwSc57mb65nC9cCKTq+za1uVek
7rB7tXxiUQTOvkUY9IyUj17fcrwR4LX9uqb9y8nYhzw/3PUgni+hPDW/zCAzEfBFc2ecvSkog/qw
4lWGnsGB8/Glpfj160wKy+SVmmZHZjrWbLhd0HYw+fuO6n1x4u7z+oaN82W5h0lBx5O4UENb1mbO
SNwuNAaSh8I48lk4lDL4JkwDYtl93lSfhBLDbNnHbWPtNerJQu623DCn9uJB+YGBPdemzJ9A3zus
PftaWEapV3z/rO/Z9T+Grkki5ZGpyCGUxAL49MTLTZ4Bi5fj7FQph2+p3gYjBEuhltrKjzoAW+t2
RBrraM+cbkIKxMKQOzRWUCKyoAwrf+o7EYIFDWpjMeiNMtugUwmEFhd37pcpxL/pVmviYu2YHEDf
ZaHdnj4pVjfYFsDM2tLhekRhx8Ii+jfZLuigu4hC6c8MaPetg9oafaPXwJ4QyTrbLaUEay7q3U4b
zM7UTE4XCiljGk7ot+9Seh+kssyGN6+o2WtJ0GCclgkseFKdJpog65Nf6Lsbrh8IYaQtvqqV0xAK
NEIcZDinQ9SRhmvUN+KqPFvD6YKOIGXmrfwtybLr1k5gkriJpY0743xns8pbztlVxYRbVk+IiIbY
JlM1CGU/F0skL0aF0sU7UBtHu1ntObuDQh8mdwn3nN9j1ZCjxoW9cAKvKiRFtvTBOe7+9KJbiFfn
0Sla5dVRgdv15aCnsd4mUFx+nT8H73ZCZicobf5uKpf2Z/S4jSLy3wnnh2GLPf3UDsBILVnWyAup
QMe5NfhjDXF+NEq3Z8U8W44H37qriMVrqK5XuXgN60folB2bId/gRJjccPEFPGEFtylrT3ms4G50
mU6SDF6xYck1AGz8yG2uX3TvZpdYIBKPdodxMtd4ATxu+E9rrlB0nRitmQkNIMaPD3MKDbdoL31W
lc+aPvA2dFa1z7SSVfW9szqVSHTZzjQIJg8M5CWHpw6sLPSNx1UPxd3zfk7N0kBDYGg+mM8nQRum
+hR08fFsZFGLqVP0Z8jxdGFvh4Y1cu+9YPC1M6qgk/4Mb0sT9vYWhwpg+pOcM978ygXrdqIpxEQN
iZvzCSOKPzKO+CqqTxSSGomtHuFxL2jJxl23doV85x44yi/scdpK7/PZuA6wnPcxRSZCv//FT6ZX
Q4LfUylD/XhFG0SIkMUeLgnSRj/PiAFa906vic29ozjrl/soRgMHoE2gMkGFvuAwTWansDMCmA1c
ldtepiHNqiyBFnRdYMVrBWKYoUh/wQKf2QF662B336eCpZUq3sOztp93XpGmINRgL81tpf4mvKmS
CvesmhMcgfp+9S7WwK3MgCxVCYd1Eow/LLsdw3LHlxBAlIpxnHoqkZym+Wdo2pL2iMFLUx7UzTrZ
kEGnpOCeat7Y1mhkiRAnBeSTdLRH0e9V5SbC6vs4DeYAqbMZhne5OKfAjuxxHG6SnwU0UI/HtTDN
FVgJ3D3YqM2gaxE5dI83Db9qRrLBMlHO0OoM5S2ywZE9JliAoMC65tYq4ZynK9ihvovZbQK40gff
gQwNIwmOTm2K5BXTW/z4E/LiWcjWVrNHjubvr1uXK2X4atRoKjaqQMtLJrtz/H9k7KA/Rhbd9NAh
L5UE6J22i6scimOQvXWJyUdGukuqGZYxVsNted5zBcj3u8DIi19xPY5AvO0CkAIoYahg6ofFXnAz
8NL0SXStmR9C/jPAShSzqhCP9CFqypeW1gZSzJ6cq+8LORbIMmaFPhdSlNpahUIij0FkzVO9iuB1
PrvoCQLYvvvR/ybgKTHlvv4T4JJm8dXQ/WP9Jcf96R7j3q07lw4E1eRfQJGZh7nz8KVOOvBlF93l
1BRvMB8K0x/DkMgRsErB6jWOX3WAWodDwz85q8kjBNcWvhUk/HlqOYgLtEGGcjBOMSD8RXGBpB68
zmuK8wZBYgAbpqsqRGJY7HBDPfzHZI2kkj7C0IpZnN/xbb7wiVtxfW9pAP+SyGAVayq8NSMsX77x
8By57oM/aiAyomq4HUEE4Q6zwUeLO+5p2zLT463z+z71o2+9812pxhAq5C2gnOvO/kXqx7WGHCaa
THLvIeG2mgTHNfjn052dijoaRpBy71npe6VQf4bNh0DJesvbP/LRVOzkqHonpKgIb/Jz4Add6tya
lyIsbdc1vxaa5D6AP5Q9x2e/ucPIrdhNxqR3YKhxUIqU7nmHh9Q3JexBVb3cbAVLgSOvNTXaWv7H
j92Qi1VvG0VJkrkTxYNVG/UMpKiiG1TwvGcd14Ar7/RLUORl+TqmnW2ba8Id5euT+XrKc3kSBM0Z
t/HokiAcftAV7Eo776QQODqSDD+AaVXOAaaJWZdujT62fdXrvGLfhuCo6v0wgc6yemk+OESHnU1J
2T4u3XwsRCD7+T42dvX2do0hSCesUQAT0i4oOgcIiCaoE4yc38hrjOa1reBJXBBd4f5F9zaXSrfH
fLo45g+3UMxXsya3DtgyX/lH91dFlwWECsuya+EleAvo8UdVKFr0VIG4zCw9+xENmRYyg2alXTQe
3JSmsL+/vc7o1z5mqiCEBeh3TkWctsK1PMdaJ7+FB3dGZNiBf34DLAyVaTX4GcGy5blRigxui9gv
nJH+kdavcPBZVY+vIMe4nQ+LKxvwwpUu+2V44XHmBzfPXVVAF3AxDCz153IJg0dY1NukX/pMSp9C
IuiRtQ1Y6CTBGZzzdap9d4vLOCE+uua081kftkU1xC8thOsnud0M7iq/LlguPE0wElXWu52m4VOi
MBwRQdaw+DllmgT1GcTVoIRPe1q7CYyjjckP2eTK2OvfOD41b7IsXIdMbImSSAWmbX7sTn/026kh
2Cq/VrIzHT5CGPJCBPjh+CHLXaQJdmZFQ5mHLD6gU3WJoVYOG9Kga34sTqOmOGUUn42hey6k/9b/
QjjMGRFyfbtqd1oG0bF3XGesCvR/Bj4u6WmBg2rOnFP3UK676NlNDdlfWsoV+T4aqjLX1g1FXFKr
AjolHQ42qZJWt1ykfVGsacj9hPLe4oM5o9RIPa3Qib5++dpGOLUZsWrqVNGMTJxxGoZkVqc7qjqS
6pqdfQ47YCcYAXXj/aK9aN6WrAInK7Sz/Jff7IYZZcJizTeTj25LERfg/NPheaXb+kTau+bpRq9i
9mKGVyRmttyFpEcBiyo84fROVN5ijyoiPFXfQ25BjBelZYVpJzORNG5SimBEMuw+5dmiLCkiEElK
c/tgy74vQE4dN+PHzADoslMr01a33mo9i9lfA+48tShsTMGqISVR4G3O/E726iog3n0DOxf5bdtS
1iBwhHk4+aWKDTxv9LVQ9yHQPamHTf01JwL+n+E+yV//vqc7TP1C6+fcYWSgegTfyCKB2q7QBSV3
0pJJAjtB5JX6qfzTvfJorZXrF4rT4CSbfUunHzy7hEjQbWqcn4Gw0sC3Q1tQDvpHWhKDE0wsvQ+t
bVLYW2udgE3Xvjkam3ZWWgZvnKQnnXRNBMvRlm9wvBevyyJZ27lFVMWO5Gk0EmwX8JaMsJdTj20+
T0tTuzOePr8Bqsf8eZ20F6XuxVzjw/1Nd2bAa36JuG6F966gv7Pz+D0ndJ+4qtdgmOGamAQgv7J0
rZzUb8W4fUedHolU0AmG/1euY+b6QvG5uZ0pjq3uMZQpaQ/K5JOodGK2RbnLHAl4wnxdMZDHvHfC
1zpcSuJCK/KzvArf4UKGtM570I2ydS+3LNHusS+Vif94NopuGEHolNowXcTo/fDVclSdOGVQob/Q
+YreKx/Jdy+qjHvcPI/kQrkNnt91jNUSeSlC5r+opWtvy0wpsPTzECO0AFIK0UpKUaUIGWsBN+ia
j2hI+gqDehj91A/uegUz3CZdloijDzNXNV4DyGu4UIpip4h3/sa3RO34sqlxLzYfoZyotl8pMaCJ
QGMtZ6CUpGEPgV0ZdKustjU+hv5mXdxeL1C6MinyJZkKoCM8hXGhz9FJNkcyEZy6LnLj0PCJ2mVu
NZ1STwslOAUv5TObj+g3lc/PAXTnwCY+IJh1i3ImAbUGkGJmirWL81+DkkDQIDexG2+Ir9mfpSDa
QYDYZwxxAK30lIVgHSeMw3hNeDtHo58NHsOFwjajRfzIraGQ1LjbsSXRh3I8UORQPq6j12Yd0sJj
PF4VvIGgH1Zvs62tWWA/cPidkP7yRVoeNWC+avOGmTCO0ILX1wa8vtSQIkNinGaKkWT2D+vzY0J8
3UGpCvfNCXf7Q77OqkVYuZ4yo9EMF2XDincv7Hp/D9vmfv7KF5JgLTQTb2voq73GQzAUjlCaPAqf
NB0RpLCC8cabzFtNU2RPKLusz21s9QNipx3q/jXdTFYRraP3aGPqG0HWGbo6mfnSWr+aFiNr3KLI
sh/vcOsZiaigfRGp3iDbN04idZPOKoTUBvqS3VFb8r1bG/BZBskQJNAjVLs7HNN8J0vQIogF242h
KJaCu6i+l4OAVaJILrS6X4M3wk/+6Sy9h0kjPvLozGgJXS1aWP6wMFt8z4DUgtikmo4wwYNeWNEY
P8msIbCjFLUGbXMnJQeQkmlrly0aV2P5VYL/HULQ/TfVj/374CrNAAv1gI9cONeahSgT1omsEYXy
LYkG59Thizcc2997WnQ3vYyOnNEwpgfCpE3NoTbFK6mDymzRqAdgpNNMh06U5hbgRS+hY/g8t8f7
bFYUnZn5YBmoRIkrj9u4Ln2yVusoPgZtoSXr1TGwiCNXsCEK+kmDkL4orp9lszAvEMz67+HQm1oL
nzDM75kWBrMxGlxjOLRj/gP8nRcWdABoUOcVvhZdwy0ytLRu45xUmfDPNL4rS7Jp8hA2DvXMBH2+
ngsshl0HnCSmK6CeDVsgShitNVWYBIutSEjGRVC+xCgkmrjaB4Cap32nsbNWxEXkS5hTNowoIPWR
cfYIU0qWagBbJjtmailXwEgrq1OA/c7m50zGWx6cb8T5SxANLX7t2PBQfrVOnYf1Vqx6lmdt028g
ua3+ypucnWoEWkHukZ+8pmrhLyMQ9/ZLmG+nuJ1CKENDrDJy0uWqfk4mPbconbEAa8Zf/B4aMELh
PTKI1iR5dxT4eAQd6I005mnDDuUVo7UnxzppSShtSByVqn7qiaXIee5QRRjiDTQdXnbFYqmCR/CI
9g45/TnJP5Ed+Fa049WT4sPsbpyBc7eXVb5jJ/lM5TF1TJDJdSWDmxXVTTq/UfDfXyHMqZmkemxG
/Z2diAylG0VKBpLeYdrkccIVNO1q1P2wGha/aA0sDpKKUDx998K3KkAfMBIDeDcHqtJLIPSGOO07
r4HaPP3scNCkbw/mkAcU4Q64ZPxBZqvSoa37umnmBqT9D91ig93o1G/HvBuqRI0D55aEJbEH/ZYt
CPxeYhAWU38ThTwTfaQvZrrnsY1qLDalEofHDP0hZoXORaSv4D/c8OSezDaRQJ8458QjrWps15vI
TBOq0tPHX6r1wYntzU54rwBF52anJD9I/T/N4EjfjhBIswIkD6MPO0FE633qrstSuU/vQcp87zr4
rHDsyff79rBPDmC0NQ916DzttCqOd8mfcxByShcrCbcvAyp8+xRePG0BnPOcIg8Hn9K4JGZAV7Sj
8Se785XO8npJ74/BDBeKHmdaBGJcBttbVU94GK33fFj7OpTMQi2qwTuALk2IE0/t/4D6WmmTpRf4
JgoFy3rSQ4f0113uE5v0nUkF1QYFOIGNyogSu6C3UaR6gQOv6rGTV6NchBGWpEepfD0QSrkjhWEt
PNvViyyJVwJ66tHifdnriKLguUKUlNgM1iPtnc8e0EBnqX3B79XiNEUeD4ZiCpQpKyXrk5UBBfol
rjsG+3Yww885prb6MkUb+LNo7q2G2bdk+ZAe85xL4f9eGA1EpE7fFOfRiSsvkvBqxoU5uGkUTs6D
WWpMwI3yo3hWbe87+meyGTotquggIuRybtiL/z0VxZRTj9VYB7+sBG41yNEffIra7ru+P6D/QiJu
SpL5hY8OAKORyXnPilx86GwMaVGHaFH+xnxjM0Y6BVniBQcvCqHZp2WfTnH2h77IA/YDjxNQ7zMD
qocrTAE0v5hx6F284PA/jK8gUVraX7qxpkoVo9QbiOjE4p+pBtNJFibZuwy3yHu9CzoyCWPZJbZt
kF+C3De6LHL2x3wTNs5aDR6Ljbm1pMEoN0+cl15gEVs7Ms71ZM+cYfq3OSu5YwM5B7CA5/C9/rkn
u3fwpXMrbMDmNkB6b7qTYsJqdZWOa3wy1NSfsZ50Ivsa88SonEP2axbPMdBAGTJA9dK93cZ918eV
U4Ol2czUwylHhdCevGD9dDsYJlQ67J+ooTY9UZuH9vyUn7HSZuIHXXHIrFH3+iXm/oyEvlpXPnMM
3Blv94sGvPznxBcw/kqYlaBiqBwWml9MIWXRgjZOthSURjleCG3jOi95taQJ0hPuL2Zi6aHqKz8Q
pZ4InLWJ4Qta/62Da/gHiR0Onu9d26qQI6w2UiU6nASBB81v3pzpA5rGqhstn3X+s+iH2rELzPmf
aIsBaetgPuvJnV/PTSZ9sNVTOltkJ6wLW6xoSA0grzBQja88hgXGqLk8k3aXHSYAWc/gUDAtVLcA
ZweGpoyy+l58kznrwWdygsq6LM2EG7bO+qZGHwdDq8gg2kMbiAli7KmAUKrzKHp6o3of/VuSYI+I
qs7WAfbpGLoFgxDUzRO6ZRTj/ZJlX23kJ3bDPI65fB7uQEZVy+/ikwGa/1F4aWkZ+qBQ84hx2xzf
jMF00KDd4f5Wb/RoOomkiGRPP5zCx78kyIE7HmmjM3aJwZIVDKNSVIXbbfcbSHwzMi1nYGdpfUzi
BGte9HSlkCIHgyy9bi2QfCPtw5uAgS7A4+qZZxp9wXv+cMRM1CQ1mwbbkQaGfT5FFVHmKnVTC9Et
ulFPjz+ebbZZKlvezj9taNMJwTeaWlRwkmJmPHLKp9Z9MLy26agVcpJDllRKGRHL51bDTL2neaWU
6XI0dpi9MrJYkbCRR0sZtFhB5pFOngbesFat6fbjTaZAuFXlESvyH7zuDCuVVDlD8zoBi0PqUlFA
vKHv4zsZS3OGR92Qwji0XRt1OkbZ2n6qLu5YDw8HEozJ7YCm534/HmEqUqrYbynE3gYJWG92Y7Di
ctRDWaIdf0N589dG5VHhfdVHpvoNDXzY1uXmTOifvCZMV+9P7WJaY1glnPaPcW/K2QOVpGNxxwLx
4U7+LNGDMAfsehyjxWo5KN4cuvTuNbcX8v+wjvqwBqiIVAVoWdWMWbb7BbfpQDsuZWivoMEd+6Pq
zbYMyw+8YTwyjVRGv3EkgCp+EUOqoWZ71MImb/H1LpFVOw4tXi3fA83ZchfvtMZqKSt/JxYEEFwb
u8ybnxtqPl/JSjVJN4VYd82uQGtI/TkNdhJ9btE7Ar2g0MOuEWvlNFiBRRrTAt/MVbQNwD8liISS
XT3Hz9poKWt0CMZJTSQmPU3uTghoCJpOEisPZsduwmD2Vxp6PIpgsooyESneQ99SCDPpeQUca3lL
xnxaxdwG/0j5cF5DHCvPYxsdjmz0hgL9LJxSjAm+z7dia2rPCEhAHlVWWpSjg/bvLo5alI613+ea
lIWGSRYS+5sdoXaLSNtAl08Z9sSkKu6CSfIadIpMPYkoTYo/eyN7bvanF/ku6BkVcirsJBbCyQLh
BpxUsMSBCVgKJEaPNkjpP9on7IFhRIyljfeQ/49SsThlCm6aKvRnp/UjDIoNZ51TM2OuPRrl/Pf3
DFapCi5l8oAUdujqVmdsyp48TvcdPQL2zQppxIE5QiAuMbX3Erf00uY3RR/lVadyNtI603aY/vte
bh+GTzP7YvtLdgyvEUzini8s3EKQ+7gWgdDLkH4h8CtdgXPDCK+Nu4B9JOGk9UeHACEcOW5LWxW4
n+IXaoNMWDswvCNBgRhAanU7q6FK1GARm/bwmhiCotV2DETisLuKeOjMjGefzau2QLvAQg4zIC4f
S8xg+l7luraS83dvYihu42xigo2Ceqkncpnrgj72AxKLjqv1GRk8E7nprOStblbsqLyKlGKAUb6D
fSPvtOxQCeE6Taf4UCMTxEYHcb373I6dK8sOmVnHo4YTuSXNx1//ksjlEoi+aR+d0zuiGd7XUUfJ
dH0nCJvFAIvRLbj+XMUXmYFpKtGr2CqkLOQbxKSjIl0+b4+4M1SEyeI51O5COJTjnHt6AA8hcSUc
YNXbYMo7+jQ07TvB3GV0XYA5r/kR+QLGu9DTvaZFKZbPZg6a5otmt3DKX/k1U5tBJrJAkeVf+kTA
+CD4Qnw7b6R43uDZL0pq7HfgQVPbpdvWS5sf7nHs/w3aS4GSCDQKGVbRN3wEcxxPd2eaSkInjo6c
mqCk1M8jj++20L3iI9DKUQwN7fm3H2A3b9jsHBafCeBLHlLow10K2IxMmpViv0BV2nkRHREs/IfK
DxQnjBpYsva18509ZJn82+fdY4R2LVVSTw6XLzl03YsfPcg8M0KhDXGRzIYQ28hJuhqIMVjsz4sf
Y34ISM/AwMP5q/c4gOoEZ6XtCeqBEEP1exj/wZr6hoQRat6VXwgqtIiqWflB6iJBXdTuPM5pUpHr
dfjReHrQmphJtPtupAVO8CPLPxZnMGVndHrmvME2bqb932mjpYOGrn5TfgWua8fkJQyb9cllwFjE
wTEKRyPh3BTi7ypPTAtoQqvCPQH6mlbHJqmCdRgx39t4SV0uW2DUhrGZL64A3F6T+CdhQcN++mor
cTouaFrmq3EGM2x4/xbdL2lobjdT+2S0oUUbEDn8fWoGtaDQzdztWG1siHrTdxJKs3i/qQOm7zMa
y8S+G7b2aNHTvFE6KEp+HogFZEBZQayuetSCiNeVlR59DAnHNfsN3uvSss4/vv2HgFjYi4v+ryxH
gh+PrA0gTEIp9ELJuvuuz1hMh8aRY9DXJdVe0zdDlrLbu2xeGjOfDhmEMBF5DB5tHLgRsSdFjs9j
efiv6XwwpgK//cf/JC/C9tLkls8+bwvxe4rgOQxKjUzZpKcDXsUIAaIG/qggjieUshpYpf3O63TD
MnURpHY5+GQoBZg35/xcLaaelmwuLOQnhC2EkDqjOxR3hTaoUu9wU6Kjx0m96p33JBaNbiEadUFu
JMebSNuoOdpKPqIcCEKYBwctAyhx9xCjO4rCzDxLRbwMLHPhdBbxquqDln/FU7P5APykD4Y/VJs2
oTBHLHOceeyo6teNtwoIq/+Ml0o/bbgdkqp+Yi5pDbMSchJB1FcO3xJZlUwLgRStd2Gtu1Teajc4
SgMyC92ODhXbPKL/cMFfcoCrEWNte55LmwDymBBuFPTkELLyXMT7j7Royjb5QUkUdWryBtCfkSXk
VEh71gHcPgs8eZtGlYfK95/wrxejR5peXwY6VWGXLj4mAhFacrNB0R6scfE5HHnUzxs0TeJAOL+J
dZ/fTAXBW9HOQcoSZ+C5QxCU2lSiiCoVpymqzJEEDwAJ7ttMCA75bMIyGKyuThelsEDjNwNp5B2S
1iI9UwLBljTOZAHlY8k3232168lpSU2a9cTK/QgWW6QMYbgdcx8t1DceXx71VmjJTrGej7ksigJC
RsDAF3Bx193prHYTA7PrU28UpPwVYMHoRG2brY67UXujpVOirL/evjb9LjV9yjzcrTZlVwrBLr43
R/PW10TVdLWPtf+awjbjrdARuSBVe3/CVG6zgG2nintm1cfWq7aonzDc2qKMRbmAv3sdWFsqfVv4
FGFwq84xp0GTZlTQ7mKRzBOsVRTGV74XxT3GNFv5L31C3GU7ER1W1wvB6sGVLL5nTCsxKuAvrgd2
jSttjjfqkPZeuqmTi0xez4z9Wn9YpiIjT+PNUGLdZOtgfPUEBkaSakD3jS7PA5KtXeIXVbgxl+nD
qLOK40q0M4kykzyFF9W8gLnpf8vUHl8HiPmQeqse6VJ03AmtnALefYtZybyfWK8lq5h97mOCME4g
3OIpdq59MnmYm0DxvSfR3PKJnYf1hOH4tC5AJ8SaKnR1DP0HJhutcTxzjlH9rjkPFHXjrQZwrsCs
r2vDO7LiGCTRFx3Z6S0zaAVTF4eQk5BiM3/M3biwaRVPep2BNQFUrGsjRkpnykQBGiW7EzpAc6RF
J2+0JkD89psSSgP7RV3VedJVy45zXnysZfyKOuDV1xahbwuFZqp78Z0sviUeU+ETW8ZHlaEK+xt3
TMpYhcCnMf3ELLsCdKjuIQcFOF7RXexhvyhQNtiZH1ERTe5YR5HDtMldYDItIwoF/b+JAP3YhdYR
gNjpaL0+t5ZeiLtylo8t2i2tefrsIzFedL0HEQNoqQlFG6uYOC+pWfHizHcRcEnj6R8i4iK2vVpN
Zzkul8yvggFX6sFpoGx9fC6NJNL3fchipxA1V2gnUqTluBnEyMPHrzHvkSErJ/jpx1jZz9th1Apv
eI3mZjf9cL3se+ChVySJvSVgnfFvc1Z2Xtyxq9ieA1fcadUTaFZ/bApRvCv7EDDzvg6MVCUNOz/F
cN0MvTToxFLw/y3FOk3UG0DS5kJcxsYejrNcTFISVDQZzXj9H+2aG+VBR0PjFhojuWJN0HEOPHlm
3DWYIfuSAhoXmWsqeXEtRYnJ3GJqBNaYqdXmqt/VSQCbIa9D1cQNM0kV7XDHRM94pjZv7TmMaNdW
NgJKcS/MXVUEMUPMKY/wUD4wf4gyDFqnMBH8yTbzhB2L4kHbX+YQ5rcIfZk1ogJalveHrqJUIKOA
e9qXmfDhbE/HSPwKQKFPJ2Lq5UHlxtPl8QKiK9Ry04jWm2wu+QeF/M9FJkT+QfpCvklXErh4+dm+
ciiYF9i9uXsk2lMepW64oFZYDOF/fUFz36CObm+IvgRymvCVLl93z4TQZVQbgRLx0ZztHTq5DBtX
LdlqP/aaCPMnifksxkZt1qJYbOzI3AB1b/Kro/+UHeqPw6KyOOZBJqK1dmbvCEzyLVpbznA5apd0
ywUbsqJSKWw21r86X1ydcZhB3HzeFIG+jNPzcX7b/N0uim+2qz9dX0sEoFUF4BaK8qTrrmTJT5dg
s5Jkb0Y4AdlZ6PKpWfy4otEhFBFnT1Jf1pv6HXCyNLNTJ9cz+J2IivDO4z8RglWiVsUgBITxNXdM
S2bwMGgT4DuP4x25Vtnr701Bwq3oRyHjjY5Nn6BPzC1BrKkAYRY84AQ4cusEowgduOdb+79UCn9l
+W/3hxFwG1+vPScrdhpBf2DU4/ws4ydaHfSYXxTBWfLQ9noYiNpRBcf+VHmDhoYn70YzxYh+1hMk
3tvO/xIkeZeKuUdd+h319RLKda46oD7t5wADeIEeG1GKU7GtFKfbzZe1yl0Zso093/bhPmzBiIXP
PqmE26KCLxvhgQoGTf63nftFtf2+6mG+W+kMXeJFF12q1wxGhasrsG9U2GgeOBizu5bwGE3bztQV
D2Dmc28AqtVTKv+Vnd3c2TuZJ5Oue0ie4WFy14EVH013tRoFkJZFTy8b8Si4EspdQD8tP/8Irdeb
VHoUwBwaHGDtHhylUL4kUuoZL68KemvUF4EDVGeo4wWkfetdD2QobnxFe2MRumStf3yCCrdgXnZN
l/R7sXwxJp5/qx1XSPU5m/d4LZmWLSF019JYBhaC0m/TprYy5Xz5kOzfxUee1cpPT9fgc5X1DG32
YK1QlK63xzFSFveV3Vy38WFbqopoAuMKepgaMz5fxNQi0a5hL+T8+5DSYCzBzGkiGnm7fy3GF2L9
mAfXmSK9tU8NKbmC41biJ+qePLfxrrGrvqImrGubsGxiR1HwnvierR3alCxdZahXPJu2U0W2Bf0d
lug2saceVlktykIIwlhmor6LoHuFsN+BCzO4/9fJDPsbqV8tS6NI4rmVtOCOBTsFKOjiWDgxhEcn
EmdFKSVmS1If4GgQufSNgruCadOm6iPw+UOol//v+GmV6a3tEcUPtDV2r06dRLMBLhtpCp38RLjQ
v6N0LnMvDl4kSwIzlU3y88BNQ+YPBXvJa5Pdk5qyM0Alw/8pTpQ3DWsoMmvszIf4R70XQQ1aYfFd
+KaOzpNqA+5H1CbIzcYLIuVUxfIJaFOd/QLBPxgFvKzXsNN0IZQD293nbE5xanucR5RBXUvqM4VS
2Lu/ZsyLoy8gvKHp2M9Ed9vZbKvwagxxhpFqsOnDtJwakOWUcogXKvNHgsvFW4IK3aZyDz9AIeup
rsNDT7TSX5FVmyLgmxrwnXv3JvafGx/l5wFRTHSWp33hnfRfFAPvEND5xNFo6n0pyy8V3btJjKoZ
KQ6YgpbTxvE9K85/A9LxtRrLGE1c9oOE3J+gL9XoAWGs6k1mivAaDS5Jzf+pBY7heDO7A70YAy/O
/+O9Ur9Ex4uvHQK/z1kqKElS3wF2jJYS1D6zjrEGZgbcNUHVwRSlwtxcI1YMRCq5LSHydJmsH9aG
1QkONb/ZpbkSJehRm3cyixT0TSkt5P0Y5+nqpwy5zrwafkrUjS0wbn6oBq5BmS4KvdlmLzR+W80/
vort4WZoC2oyuY2548O5EXG+NGu+9KIHvnHo0HhxAxaHOKp8YeyZ5+mEW8RSGTnlFMRarJ3S7CKT
ZprfVjZzzXJAm3YTyWqI5aIIMZItFBmrCwd+EWn6g5LO6DXMEJlxuAz7uFk8Og2aTqVmAGq+INyz
ppjPBbkyfQDmU9kBz9orQdOWa6xg0sFTGR4WI02GKFOC+dw656DBZwFwldgq4Ks+g8qkx7k2HjzG
BQE3OWz/t4ysXWBSiUycybIB0rVdCf4L/EiNp1grPbZnOcGh8xDST5HUw5gCsY5q13JN/DpD49uK
qvHbyZC+9fJf4nrT3Aai4LJxMTucIKNXxmhHhLlacfTwD0D5T0h2HXCA8/RbDuxcuICiWzOwD4YB
SGymJ3zt2nxPrM4yOn1SrN1fE97eP1XvEUPAOzdNRCqIRUySnssjnWjOqvJusBH9USt4MKAf11xy
jlOsSWA+1Zzc2qfWW+H3I3pduTxX1PAuTyDZDGveh4c16wu3oQckktStwSrnqMts+VclaPbgGwWE
d3bKK9u91F5TzG1IBk0506ClqOjaLjpEb0xJfY5xjoOQHb9jP+DjqU2c564wVyDMv032PcAkjuI0
hxeDGHN77Gzawe3dbJSnpEsURPHQ60Mc8kBPi60JTz5hZc9BsuU52bRyNcQPIH4ssJXTLnjvQXxj
K0AfrAK5UcKOdtLsoFTAGxutmUwwJcOnG3IKeQHltBkwqePM9VPYNqRv02PZsWXNgwJ7F7FrN0x0
ewJSRWNmqSH4suDoSHMaeslA5g8klj/iXU4ZtnbGmtYDYja7G8wMK0foIFj3IfvikTfgPOVueVi0
lm8/IuLfCd0n8XwMtvn6Htz/zzRBjpyfnXb1xQvZcHXCOwku3S3xPKfRhN0GPI1CiGRUJf6TLjRo
b11SctP63Qce7++4UjFGnTMn3rp1F9pi3DuYXOumoh3XPMZ0zFlCTx9gv8+FRold/wbY36MVj5F7
1h5MEWJvCDkWMFLcKGhpPzNi6m8ozIro8b6c/fFYgLgtEZ3TQ811QvJgSIV4U9I34NVCPZteV4cU
2PEUnHPizertdfh5JD4r0OwjjXsZ8m53V10iNkuBmSUumHiTc98uS5iZIqafdemuX/gczUzEKAJs
U+59hooCAoyqdaIN5eSWDx+88ufzbhZgkkWsKhoTN9VmkZbf3HsbCcm/McgYdaQKKrZvOcGOl1EG
ZCbWMLMYRKYv1KrQj2o8x5UPoXACLqkYEYnkgfHPU8S35cXV5KCZjZ+1I9qkCc3paO0qckUMm8Xq
EIIO+qgn30zwfYn3+6d9DqZYgjQNcFnEB6i1sya9eEvgbP8YY72+JZ7u7HR6/w/e2iljLa0kETYj
OzMwWNJksJPugjPHlJdG9ON0fCNXIcaWGqPJSeSMZ22JcvEK4mBLg4DoYrHAYx9u6+zPwL+zV008
F5uRb4FVIQfxLg4BrpLTq0CXTy+HNA9NoN+2QXvUagjzodYG/ny7+bUchbDA9fRlywiy1mnSjlub
4Dk3ceURlrw3O+1W4wETMGB9ugCrdk7ZpSAFacCRGEbDVMf2gXcwmXkWWLCVR3KsGtbGcSlCqzQW
lbG0dAdfjLJDMMfUrfOnrJZgnDHJ5m43hz28OpWFeFikpL4RMZzmaYAh0sQSFkCf2I079gzut/Cr
dMSlSy4Zxx+TEopP2jKLvD5jDG7mh9oA2dNVbhMrzSp5eTnzpSMp5vlJHwxP5knDZEc9/mghzaRJ
ab+5pi7QQ6+4JsOuQoY65hIQTrR3dv4/ImJiF12Ec6xuFZtG1q/Js/GJbPG0xUUi46pz7uhB/IIa
bl3HZwHjDSUon13ScpidWdgbD0t1y5BmgPHZUa9lZCtArbFE+vRmht1kruOAwWAz4klg3IMb7SiO
nQO9Lz/TBRu/S2dpUeu9OGPX3P4X3TQrFtlwumny3KhGbhgDFVc05WqCAbRKs47HudnBtCE/RkPF
6mQKKrHsMYSbWaumJnqdJ35wHbaRyvY1ahd5EcQywnynBMLao70DdkXwis2FRfN3ND0uC+lPRpfe
wmNGhYrQUJZLxcOB0024+rWKCtEjXh6IMr9b8Cr+MQGppP8XilBS5Vory+lvr3cC6NybQlQx/WSf
ngMuesbo59fSrwUP1jd1mwuddq1IgKcYutfcHIjnDVkPQojj7LlvrNQGv+W1r1ZKl1XpCe82KjcU
SUXN5iWjetxHVA9k+t0aLb4Q0tXmhvZEahEambXYO+1rC3vArjhOvOrVbQadugnlSuEZTCe0LtqV
AXXisvQ1+mDa4eBCNqlzNqw0Qiuq32WMS+JUfDvMQbyKuWSoh7u7jGJDh7Zfo8QVini7pjTmQqE+
UI6SRIT4OuNAUjGLMWPY0SjmuDzKUPi7aXJp8xcSl0C5RvxY9qVhgkMStHqZuRrZsM51NQQ8wLpv
+PD24rEvWdVpK/DIq+m1NcCllL5DSJHR3xccqOVJ5xeXxHNbE0D590MZKzXXuchYRC2l7kHcFkTe
M7fIpjPW+Ll7fkg5LeEzKcHyghfa3JVSZFH2ff6XuQgTgdrS4bHdt4BEtiJkml6HiU/mpZWpPqNy
0ZGzP55NRv7cnRFhWw2CKn9g4tkoBni03MpgG2sd3Xa03r/ggW21a2wnCN6Pzg2mzlRF3aYKlQ0l
kjp5RXyI/ZVT/j1cYka5edw4Y3JdXGtxzF2c1dHSxV1tYemxD/FLOzlvg8HM0oXvW0Wg+VmUc0F8
6YPsG80BCs6IQ/dp3uRqoU5UJbBB5dKJoE4FtwMjMCYuqwMBwgH5ZByu4d3XoA0LJs37ZXKPdn9i
H2LvFfpFafKkXsRDsDJ1jsjkZbf9NU36Rq+F94PRpEniOvcpa/5GAnWjzlzHhyatYfvM45T55xFe
rHVznwFOQ60fht+km9KaZC1nsz8tZQfBHuoxyG6LlU6+TR5uEFD9cFmYNfsF22lXz0VTgaUOHUFO
mzixW8065PealG+Kpy+Ic7P4Kb0/JxUqvHAOVEjVKGac0jLYpgH8kl6hORoUT2H3+9H3zSGKlCor
kKzZztMNXaoq2tsg0lZRRMo/rAN8peNnahCf6Uao+KP2OP6pSzCiEGbsmMHw/mYBE/RMLuvt2bGg
D7FaEGygNTAjW8M7FsJHXdjHvnLxm6Gt2MXaVyTQ+mW10WRAGFBgxb0VWRthqonMNQEjx3IM2SeR
F7TFcutQOqz83+PW8rpruVUZsr3LohlGCCRzOxAePJwEMUUgOO2rWUy5vGJAO7PhGq4unYT6hOhp
xNi+0MpcpAeWtg3ICnD0RJCBzLREmQ59gJ+ANw7dPLlyVWRx5ivJ/qxdHmnKKvAj8f8/Xyt+5CSl
foVw29FIJDpgasCfTtDRgUHEssrW9w4oq1Z9IU4yfGv9Fi1A+IlOb9VjoFkERi2vzllteo19qKjA
N7HGnvQIpi9DZtCnmNvVPKHqlWnOJMevr8AQgAUwDL/x8dpKA0GG40wE7z87aU30lTjbb+mtavQf
VKM5tjxXQjYQdZ/SWJGqPSntgya8is0tEE06z71IpWmurZUo5NB6i6HYZ9/zzblLe4MjwaSXVrd6
vDL6zwf1AwCWhBJ9hLWeIjH3Rw7mSZzXNkZ98UkzfFC5zPTC8QjnF+oec3kH7JoLUyGCUT8FKnMP
QVSbIpPOah+LyvsqsmgeGMEZqBjAgQsZsX2ZGiLPCvGJw5ESxMD3BeqXQ2VGXtF1tFmIT35ieG1I
QJvogZlg5uqIITuOCHbTWawf5FMpfqyYuGBm6/R315ogfSpAJqJ/GxfplrmAGMYpxsChH4zA48GD
PcnfyO66FXeSGTiwgDDEivQEpEvJZ/FOBIINIWcDNJRbgeUxe35hpZXkFD5OH7awE0e7227vGu+V
wve+vMQ+4nh6fzk0hGQvT4yct6X0SFI7Rjxw6eEUqAHS1cSxPnO414+sUJ8qJyLg835rYOM+pBuG
7bbzXoZqT2Zwf6hEoIoBEoNENpJBkFC+FiTpHbJKC7hUWbkNX6fX4d9qAcy36hiPgbvH7m6z+zjb
JTlm2t/zZKeEDlvhWi9IUhEgH/rbMwL0DcncLuJprqGoiDl36z0fx4zFFfd4AfcCWew/v4ivOt9z
gbWofrZYcz5qG929yl+KT1yjxbQBK3vt6uQM7aXd/X7Nsl6m4sZi3qTfz4lL8VFb8J+zr7H8HEte
w35hHNSspjz+VAYWtCPFe34t0ryyed7UHTw3Hj8azwoXAyuPWHn99Dx4jJEkgX6+Zp9NN8gd8TN7
K55Z+XUaokeWpOZZhXq4k9NhIb60vmFnW9BuvJIK1291ZqR6dhcEzzH8aQhu2L1Bhl/hiLX6togm
rF76Pw0qSVHRoLiPAqPPVVZK/Li8S/WHUr3Qb+f7lZHtXWMNjbqgFmy30MboqTsd3fpU/CFbe9zF
t6RvbtlPksyLnheJ5mxNqBE9tRqFNarEorA/PRjRGn6hn+X73Az0bxV6uVr36Cs+ZgiSoCbX2C7r
Rgh/KLwnaUuzkmvjAUGnU4RXqqbVbyOth2ifH9+PKrfSfRXmLYJXRYcD06BRN+5yGGyQYOEB9yEa
2p01yusDeixDB56/S4+uprCf3Jq6WzZ2YdUZUMBla1e9eQ4I+U8zU9oiBwP5wyK0bf6kluS7uS/J
okU9v3zyR7Blerm+HcOPzUZArQzHcca/DyaAQ2xDl3JiR3uTPuQJMgEt1F3NTR4T4CWzBTMKHozK
mo8sflJirAtx6PIx2ybpAgNg0kB74iVn8oB+p7Ki14R/yvtb1WiaddcusBjVOaUQ8IJLoBUrTPV0
8yfhjLFGSvajqykFT10hTbqdMjIlRt0bpW2q64z0vegBa0Ubq5FNogyoTp52UcO87hcRDqVob95X
OTRn3ARoE4Pbb32oGVCuUmZ0RB2Tu2dWGwYlsWIg8W5k2nNVP9SHtRWTM8y0OgwiK9Gy30xFfeGz
hEEoE/RZhVz+iR8Fr4FGxG6w83g0qquIROk8F19/8VxxA4V4JYjkT+ygTlkxgx1Fmy+m15t+ptGZ
W7nhA7P1EhQ7ehRIZjn3BoLQF9niNJ+23eTz0K085qppgGgww+iZjiphKvYXnSRD92D8nX4YJ5QV
TJ58VUTTTI1aFSlzELN6X45yn9c2xS+LqYlowCRrVQTPIIvqHdp24AA9yb2TTq96SI2og48tcbSh
aF/F2UDcyYemtULYH65demBu3r6DmG/WG2LG8tmHfo6H9bYONecgeRUHpbDjEE+swa+VOqPQiVjJ
gK5c9csN3K1X9j/g8r8dVkzWc95qnhwLIoZllSDQ2wEuLXMxToXOeGUcXIjCCGQ/OmyANijm098g
ZlWQTjor9+Box2koqslDlS1ww3YW5ZxFIQ+lwnRdYyPogYZVcSxjMMYq/6Ru+7X50541hBJvL+ZF
kmrqZ/YoBB63jSX3hT5FsloEAqj+2vHunTqQdUWfghRrQtplSpuQqIpo2oVpzbzbyCZatEJbrvBE
Xyw7WGlAP6ZOt7hy0MR0QED/XNOXvlBXhmk5RTKnSFT15ss485voyI3jMTK9f91bChgTDFIbVTlD
Tr9x1XEcXPKccfMnRw39tRs4Juw9fhsYKqFkqvP+i9wzp6a/d9fMh0tACU6PuhcWsL5tbx95Kb8h
8ol1dOtUbpZIgEDa+8xZENPz9+c7TDSP5PoXHJ4onI3+v3sUPhNcrLf+wJwrV1whV3TKquf1zsoi
KcGfM242mjc6K8/n4DxsLdDvpLKdzwgYUlFX29f9wFI6Fu+IlAM2ym8Jr2vgKW3AmekisYkNMo7P
hK3XQEfEXfyKBC7zBa4Ha9QIqBWzOjZ1vof6Et9EtYZ8cfYJtAaq/Ta7FUXIwN3Gij27Z2YfH1IO
L6ELXi498iEPxiTz6bfgQ7liQa6zpnLl+GTkmRU7/5Cbo7WrQWLVip1wX37Ev8kddzeJRKBLqDpu
NrlfmjdKnTAPJBzW9TUC0YAPNWzfIewS5YPCN1h/ObVsmTqRStW4Lf/bJfDn28UkVFv7wf847x0X
fIlTU04jJ8ZZcWiHgq/DDUEhoajNi7YVLpES13dc0GonDNc7dqQ65qkQPrVlRlj7+MF848DqZhia
ffqZOtYgYbqPy3ZArv0Xs0iK+V9JXSjpkowWopUbYXnCEq8iKX6ysluBpDDI9oRvYClDxydhggxw
QIju7sqJMWGE61eAH5UIkPbOX4DOHdtKDCSwTiPMZkPnPXc6t3+VmZwIZi30s2qvIzlxMRSSwHcg
ZAkkQF8M79/TMLXFMlbn/ldvZ28y9exNyYwH/iD9nDcApkqDqjQWH7vlvClstoWj9ZOc4TX8muVg
2aDJUu+4147ce15Vi4hNgYX9mXtXl371e6AKx5nyZuxn+XJUVUM37nA+FjxuogHia1F+uAh4zpzK
M+3gO1osusTSs8G0MqLTwmpFn7eTOxI93S1tZnxuwUCYxkz7BR4CS8YMyKBTywuasKqZsj/7QPud
FJqJpfF9nHXL88FEG1Z0QJOEOTN8UJ5eBCM1eHw9HRXvVSsc9sN5FkW04QtVJ/TzAfyZvdpeDVaA
vfa7v76F8NU3izJmpKQCcbj3kHKqOW941Md9fghzNYMPfqkPyvVPIM3Fwit5MMbY/e4uHiNPUjrP
58fbua6nau4CtSVsjTVu8m9I2UocOIwi7ewz3wHJSms0Tp3r7zA0byu6k20cuDL094n0ZMobHDhH
Qg+jHmxgRg5T9UO9Her7nLdcboI+JidtbPQvPxMkvk7HAglG/Hz7Jg4zj5y0kummMZpginMsYaTo
pvlUngg0pX/y0xfNAcoOSLpvHis3+HJWHRmOA1UbKKVejZj6Vu4JC/+aB/qPUW1jWd13yRZsgPTY
yLL/fgnybbFOiP8yXP0ejERjk2duiN/qQGQp69DWo/3KPL1xEfQn61/PxxlXtYmlsXMK+TiKLjJF
SMxWMZdwJ/ziU5FhSpOUvXRMFulNemX5vMbt8h6E7b6t8OLcccj+pvuIKH88mBugtgFzr9gM4p9d
u/AM0JygTvTY8/CKg+b9T6E5XRyHeGRYKY4bpX3t13eEjYLNITrssOi/JoF6ZqA+4+OJxXnIINVa
mfa91GxEW9ux+8yAFeg2j/P5lwJ4WVw4QFcd4mu6qAoCt4zm0f/0xm10+C97l1LdDrfsDoj1ewCY
V+MI6uWrZbBDVgvMLE+tJxfgy9tyLougjX3dGtnVLnd0oFnklDZBFu0Quu46/E5C40/U2vrB1kzK
f97pQVmPE+ICQSDdXOGXludKrwVxh7P0wz5oupxTm4G+954dV99l5wR2p3sghUnl3HlQ36mNjCEa
s12vnz70VLb4PAw6la4iqoulnQhnUHmLArEeq9g5JizmlgHQRpbi7CaF4Z5HAe31/KaR/OUMURo3
S4WKd71i6/19cY0IWP/ONZfeCp7T0hXPku+V98Fp4DYJPQVq5+qxRX9g5HgMwgWiOukJKFoMCcfL
onGIV0PAedrCOl2XCp3U4hRAKy1NkcLb7mMd4T8qJer3z8KUu0uJP/GZ8ZQZnTa5AvWKuDcng4eQ
qQh8+RwbtHxzOyk18TM3MHBQHszkdHyNv1Ms3UFVlYu5yGWfnF/cJrrZQFPIs1vrwt8rsIvDR4CR
oXFN/DWl7AKgBygKzxTUGfjYRDvRv0swqnF1YYUDYPcK0hta2+gNbrPB7CVdv2vc+LCohBAq2uaJ
fPX+hhECuYflh4O1lJlFUXb/5PIEmbB0wICWFHOII9QcaBx3oVizjWrkaoS2dtYHG3FtUwhKDRIb
6NlTqIbGddFo/csKrX+V8M7vW9aCbU7k/dEACnMwO4SGnpd/gsT/ehAnsX3kbTdRLndejpkbtBUy
NijUvAM3c5wP/QroqAxqZftJ5tGVlcV9+dZ2RYO8xapqsQCuV1ERjqD32116hbKSM1sQTDozit0i
zeNW/jGZ/Msnuf4uNry/YDYm8Vd4AZYi6j9Sa3x7xMTWTxUiy+BtreG1VZL/2WLhNfCLjsQznrJO
TO3DkPCVImD3s2cY5jsyu0PoRsqPR5B9Tq4nR52/MoN5v5hwL8OvZ+sp4z91BIMZoJKZwms5dzIG
jJjyjCDaIX+tElZJjSVizQCU5eIamfggMUqCrTMkk+3cXcKVVp36eHi2+Ed51JJrREluLLIxx0Zl
LZsDl7Qzq58ipFiCcUeOzvI6qKW9DQLN+IYF/kEk8zSbnVAoeXNjDMHT+LRI4GKpjHW53YnZPUdb
zQPfMf8mnUVVEkTRYVPvjFjaUw4AFBPA+IdtsOgd621edvWdqTPH2yaSMJbevcq01/t9YCqFYcJM
GF51FZCP2ZMWi4562KhmNI8c4ZNTOm7DnlB1m5qRBAgNxc+YrJSdn9QHiyiBiveWgHACExGZOe2r
KZ3//jUVlPUl9LKPujA2tk7YngnWZ/3g4nDZ/hZXffjMlXaTGSvhOi4Vfsbn20ukXupTuVviRhRA
kEa+9Z3yHYCKM+rkXQ5VFB8sYXiHw/u56ou76O/Z/KUtR+K2w5IG2Rhr0W1VTXFoj903Ow+QW82u
+CcwDi/22dUO93SlCHawImM9vIEl3lsnAOzIaDHfOj8EvSw+fahi8gIp00QWNbT+2ostoNZ08yEw
PCKzb/6hFEYAvWmtYlU0ViP2gKMWo8Sjcn30sSryimmTLS71EJuq6kF1yYakUHaae/qWbmkFNGjj
qbfxkGjjgYXjqrIX36KPI81oiz+Kj/5xyjhIwCTeOcEHiTqNV+wlalRYgfAtXdEisF116Wizt8Zo
GeVZPwCuFJPEVMoJ8hCxYaUclANpDXzzUyvo0vd3Z5hFdQY4ccBZCboUTV7kws4sUiETGK8Tf7qv
T4sDaa0t0VlHZYx2AV7MpYz78Q/amGKBL8FN7UFJfGb2ir5+SvJkWr9XEFxY1CzChZryU0DnK1MN
grxG20pI5u2xBag2dmUtsLSkFsP8Gdtd9YkB+uZaL3ntzgI7oqjduMfbWgyoTxkJfnQHvnh+KvSZ
UmAYS50tXXU89CLzp2ikaADn88oYfffdO03bAEXLhGQfhNMz/H70yyCvqtFv+Hg537Zc6GWCaR1a
3GbLODlLhVR0+9zEq9glmQ8498b520tHDf5G7DtNSUZame23RLispvB58/yC4gEZBvWJnsM+2PYm
Nf4q9JJ+xocRG4Are64ggOu51k4GQjUSSRNq8WLTh4y/Zj5+Vlmx0Er8XNng3w6axKgV5ERhu2OX
pT3KOfi7N1WQMs82jQRcr5BlHVpTd/OWO0KbBPW3aVlnudQT0dSMoE/8fN8f/oIsyiU9Gt5bNZ8+
pQnTZdokzqQ89T4TdbSxegw3OMi9M1f1N2qPcEBd81/+T2NX3maTE8GxywcSo2FKp8D9LSHnVRaT
P7ievvz/vXNI8MbiowBdCy4s1rrsjmixeptwqHjaB6OM/RPYSqlKz85C3uKX8n2U63SvT7UIFs+f
AO/xMIRdgcFyr/jpZPQ0iJsHuD8SBO2pKoRFIIuFF4HB81JkuLRupJrwxkh4Y1pUo8UKb9z472Ri
9nRCfE+pa8LQcF+sAxBIHk2h+FADd9MeQweOVDJMhoq8a+XRab95/WelH7ZymS4qt5AxuofSkbsK
y/HgbUGdp2JVoNpWmPDURbAK1KYRp7erqgk/hIyjFpkL3+4wUt/j/09uv310q9Vc1A5ajs8XDOJG
9cpoXXZyKFIf3eMCSpapclEfZJ248SLRzhl108q6mxXHMze1IvjbNFuUB26imiugt2PyBKJA0TTG
TVxd/ZC++TAR9dN9svByjg+hsMcSDR1b9rZIPkycVcEcUTZSN0blfigi9AXWx9AaqzZBvu7pjQmc
9cMjrjHrXl/zQ/pUmfQtmh2ZAHf2+6yMAWS8L7Jz+37W3siNsHBygP9o1eYx1FsA0KNWhlekRwzY
E9aXYsEWpWt1XJgco24SLYM0vYiT1VpWC8bWubyLezBATyXd0tmTpQBEiA6v+xnMyCTdup1ORo/y
wUwmDtonZv8mDVQGmT6etB5Ou7qSwiE9wDiD/zs8uNUAJi9qbbLQOVfP/QLnQZOqwycpQ2Vi/XaE
sqaVSlwWu0X6IDipfREiwIfzAU2z3Scwb1KubdRHtUrZvtcOQXF1DiIj2d/UmWcPjS6H4mz+SSSv
umyXCzP35j+fb4dxHE3suffK3YoEwCGt/7EBKosHcNr5CJ+zNbfe+xlbdL265Gfqsz8N6ap0vKfa
SzbQ+MB0Vky3dDLaZnnLANDx/zWa5DD3ax7Yzzt7OCmWQIZBR4bJp/tOj8J//51hJC2W4PLf9EET
AstXTsFmAgsia3Qvj6v7TpfrqQmdEWIG6OUTejRESZ0Y6+otr1+A84l0GvyJLTDumq95hIgbkK9v
l42RhAHwx7ExBWU5dd2YaQVSCqwDqUmEScbiLpddsAx6PTo5wrzW6ftSNL1Sgyv9jsXS5KJXVLWx
bC6Le2FoF0RZia8sgTj1srkzBQQVR369rbtrxju0CH7rUYSi0tl4DBeDP1VUa10d3UDG1/Lc0Pg0
ef1I4HNxuWIL/gvQ2qdcwsNntlkP9XybM5i1gy9EoXC5FHhoXVxmr7sdfqMfk9SG4D1NRRiU3CAl
9R0kxe2IfCEb+j5UlXv5iOyP2SJu0UjLSIYMJnaKTQOQOEfOYIN5Aug0ka/mBBbtB+71KBG+ffqc
lOoRk8ldqeN8s6zEurd2BBdgnyd6Ow9Ma+iIO6TZvLLPeduiB+HzoySEGXOaTo+Fy33mBT8x1qaJ
yVM3J69If7DDnB5+HzU0f7Z9UhdhoHHnxprYKHbw1V72o9x4hAcNFghjYCRpTCNOtRZeaCRNspQZ
l0r7x9/VxKQDmY0lrgj+8Kee8glWzeWIGXtkfsjCndr4irCngY+4si84xu9S13KhCBIJbGqJUKN9
uQRP37jrcSzXjS3KwztArVbA9uJr15fgGS91xhkYwOrCAHjsGGT9LVOFa3p007qFH8JyMuOvLAYP
cphlE1NpURoXDKzNf8EoLx/P83854aPzBM5p6qZVt/SQ/zmn7EWTfhUcCTjIJQkvUcBy5+p5FWYs
x0uDKb9xd9ltQlQXbTc9ZosuFfiEuntR6EK142gqEsndG2CHixFmSxwWqqj4q5Npj6+DKCEOfxzX
3Z+1c45Z/fV6ELbDAn3aUcyg3WbL9xGnieSnMSoLpcY5bM8BzuubFXfOHC7bzGjzBV4HwkjtaPHl
cnmthrGfWMRs6f+yYjUTbOccbc31NhXehmS4edfghSLvPpwtvwWAStd0sZGxL5yRl3BMQdPnPePf
W0D1JBqiLbgVcmXpIGVEi269lcjhuk7GwSEGaeWA/nVwlylv6ftOLdIqynbRqf+JCnSiG2aUNT6+
tX9YaqtH2SUQOW8vHzNsaIfwitfT79Q/IVYiKRFN8UKxblk5k9pIT9aFP1wUiNt4U7qcgNXqJzrJ
U0EGL4eBgIf50OwDyTJPineM5R3O2pXDv1OkcLfW22RX4FyCyjD63Qi71TLzu7Nr3zN2DYlhbpSx
xIlyfnu7OMSWeFkgF4+rfdpx+kKeAeLPhisFhQN/PbM/e4rT1qLxaGu2MD0cMcL6eqZT8pQOn8VF
CBlKjoHb2pmikwLC0QOyoPIlbEY72H6UVgJbg/pFwEtapbu7+HIlkl980z7sTgXFHvYibVgxPgPF
JbMKEPosvoQak+lvWiw75WyXAgmTWs3ikZII/jbPGmitn36m9QO7dYS07I6PT1/eGFpEdixYjgtT
G5FFUPCUV4s7vHDc2HY//IoI8pl8b4dg0U2uaFNJ0Oi/dEC1jiBX/4vpfLP7WDhQZMl0OfUdFn+U
yeRBvxoPEGirJS/4zC9gnYfzNmkVeJKnQz2njf1s40IW3vdFjQy09K3smYy7QuMrYaMGt6J4o2iw
hKonr2RUr1oFfHvJM7fGVnuQoP2XEhBcHNCjDTzLp4wY3IVGNn3YYL9mbT1WzN0BeARce4Tz4rvE
KbvjP97y39n9XfYxQM8UnvzzBL9sdZHwtWQCm9X7SGqiZJeAoiSTNkwOcoUWbVCN8bQppq+5ZvCh
tGjNAKf6hZ9PwEPOl8yc0ZoPSPBIXpdl5ZcFKdBvmG+qMmOzY2XvsIlnwqyuNOZRH+LUzS/GCt4T
jrL7AKA6xqS4YX4jKdvmzMsWrqziByX4E3gVpQmb3jrJ4bgcP12is4lcIrGZgRfoEem8Z03VQARO
ycoR84OuaR+VxcAab33+9bc19Mv/ky/mIP9iyXbJG2ggMVwOs0xzbs+Xayjh/ZK7cPREsJIPj03m
yKO+etRCIDqJoiJMEAGMPTA1VNMOYTM+jy1w14p1fX1a6LfnHL74nSgrB91a/k260dbPZmp2Re5d
s/fUtD3rgBb2Er520ODVmWtu1d0WQZXtylCyvNffhBxx+jwXWI55QQSoRQ4xHa1Lxfc91mZ08iFi
oaiERau8P3iARQgV4zXmr82qcUDoTnpebeLg/c1mZ2QiMO47M8BvMw4krRcqlaRac3xMcYH8Ut9V
lLBA1JhRCLnvW6b3LlaWZWlpF6fkc4pCMpy7yZq/QMDHjA236rpWTF+s7AGOwLzUlvyOafvRaRXI
AixhuWqJckufe2o8cqKF/PHArGBjaYM7OTGjKMCZMUcOIghKSml5XQU1FYOhfG/E1hsmYzmvgQ7A
aOglmZjLZeZDiNGNgZycKeBfPBNMqVgXD/+LDyZalVHtJIn6bJENR+c+TyIQhSotdBIz+NK4e19R
PkrpW4RXH8Ole2IV0WCPpUxnlMgG/1xE7kFf3mckBfPOmoR7PPjYnOcHrm8WbHbvFYWBkGyXeCv+
uKrO958ek4/MDvpJAbAF4XmKINtRY7rFnTC3lujGeZhaU9gQgo8A9ytkIzyod46X6lJdh7AZ/5Ws
v2qKMR+VuTh/eEDtlnu/oc+WRM7wGFQNycirSp2Lwjomb2/x5bWw/lUdsUdw/Vz9DEMCseM2OU6X
YvZQUk2Es/KpNuXsGqOJMqFxCI/74b4sCyhmI6dh/zxZoQrEK8/J4V0Yi9SjwMC3yNelp/dyKaoc
FWM3pjmFVbFW/0ttagRVP8UZ9FAts9SjM5wryWomFtdGIPaoRT7BD1PxyRlbJ2WDD2TZ9wJ9+YSN
BMp53sFJ2P8adqFw5Owfar0sePWkqoTE/87p/f3D9LkeZ5NiYXQvwYNQR/TCZssESO1GjHscNmY8
KApuW7tVIiYglYa7OQJtk6kNgPXj3nCPjuDpXn1xaFENUREuS/rAbftKejU8IBEH8AFLKwT2RRcs
pYI9+xZhNhJ/LA6V3ffvrgeljiyMGekHx61HnPaxDucvbjBzM2JgqHZpd/Wr+g9VPt8Lp6E/3qdo
NupulQIl5nojdH8OpC/WTAfKJ5i/6z8FNumPkJUD/jIi2Eo1XSQN4rtdmJnz8EVcFS/0tdRVD+Ju
fd3Vchd/Xv+2pdZLxgiw32jURWIU7q3k4HdEBDe8bJmKvmhkt5btrxUgwFt6GY3AXrJS2d9+cDvm
IGJ78d5T1uhFTOtAmUnQx0pzcHpTIUrwVaOjUpTUhx4rfGKF9k6al/LYzi5L6qOzUoJvBLXMS+D9
FsaiLRT7Dc7FkKLC5KjIEDdDMnKQJdRY1uuMdOBP4+wIejpIHDhO61yVaIoGB7FHhqnx0PQ6Vv6a
7wI7qgsqB/k+sdnF7TceBP9mK2sCw6CIMRH3X6EeTr33JzGRRtx4WjkvqfwtH0w1klt0Cg7EQP+c
ERsdt6qIY5goylZm3Jxl7EvodNUOmk4O6iUpJG9UHvYLQtz8XJpeg9kvgNhjpNbLs7Pyb7axi+4z
MIHUHas2tJVEbp9nQ3/iG/Icnls3kPX8R4v6SGXqgRoKa2XnimlEt+daC6IrezIROusfeuUiZsU4
Eax0k3PGsOU8DYvKYcjBZ6WdjjZgPSIWLowIeEk+OGH8dclgpfu68RdsFXjRFRIW3iRa/PfHgluG
vgM58XBm1pD3kpFjIuoHtwEWlvObCMyPw/8IuCNM0uAms3iXbgpy3ITqEhkKBPFqr3Ih1I4g0Shj
NgTXS6tdEZNe/XQQxrPAO1Zr05sRyvJ3P+YmpqnkmFi1ueAF64hd22Uyrb0uLU4lx7j4cWP+olOS
hYQmlmn4wgkaqCTXDdyxxmBIKe4VxUFqK2UfuU/iRW9W0kkil9cksEOBf50xJj9F28EoG3U1Cgos
HWVc0gEETFkqQ+Z94OoiLTiuTV3JXKo1Ug7aN8aFYdw0/XOvevMy7CTKRI0Kxh3NqeOkb0un+8Kr
wg4AvhfodxTHxVpxnto6Ij4tXAM9UBJrQpTlP/VgW6XqCXovwdduma1W0Oe/5qtv3ZZ62J0efdhB
QvpqZD7MtOVgULl5Z+I+xseus/OVgNLFytt4rUWTZU2OOQAm/3ahVvwXfU3uuryMUmNh/ikp9zPP
eUtkUANvUSogu3O5U79BEwHgC/sBDEKmLT08hO6wE5R7E2EscwiB8wc/c+L0CetiTr2+8E86dUdp
KDw0kmTxt4gSsqAu3Q96iGIMXdYe6vQzVMgbUC0phBdleMmOA3AI4Wzdb6fmRnYcneyOVonvjisa
jLrxCou4O9E1BYWITo54Sc1C1hFyatLE+T1QLlZlE23R8xAInKht9h5vT7kwQLEdg6OHz0p4F57l
qPKu1/PaIBvuaRf+u2SLVV1kPqIxD7iiCG7uvGG3HQiHKnJsZg2tVpE4SKtRflDAUYLUDo6IjU4R
n/790zIUYwMTMfLSqqEsT5/8Mui50/jKZMqrRvPQ7vj/9yZu7qLTLQtNbIhOf56xLVNGPzv/9/K7
4RxlJCzdAtCimYnCsr3wdN44dNLu5ALdGC/0e67ye+StK8LfWHF8gD3fv73O6T3Q4JSkQUJgqGF3
BetT9zky96NlThOueGx+H5E1jjCtqM2l18KFY2rLJUA1vYc933AC7GehQ3IneKfR4UNcXBhf/5c2
eTncVM0DMLkt5BNVbMdSzT5bsFffUIoYw3I7Fh2p9mEER6RJ3Oz9YQfMCtJmmLxifWjfK6dyXJfD
LcpZGPczkUFniPqaLj60SCEvWQKs7gdh5qzlfTrWWKqAGwN9RbEotoX+x2AMxYWSI9gePuX6bfk5
znzBgX3dSFDNPBwedUf8DESgzS3nAJQjxzOrUtmU3tVga+na+OBtLY4E7ktst6WRggOxOoRfpDma
LKDTjKaar3rLovIMwcPIjl/IEUMCc5qqhWnIORRlTKFJ6j01gUWz5ascDuop0+cBrAvF54CW2Fug
vxsFqECUpJXzgFSoVOU7vaZxzQ7TesdLLHzxeervj7b1dp3JgfbSvt28KIF5umala6QXEGfsdfCu
nVunjBtmiEC2dZ+I6kJoDHGtdkeNCEHTgD5nVZ0qrYtFBJiIHr14FCR6pCmf32d8FLwGsnRGhOVC
kLx/5JTyR1R6xBx9CcWr6Z9IaCkoeK0O08qKyQ8kWqG6uf7OeFNaMpqOSySrM50IhBk2ug9Jfsrx
imZE4MXQxeJKGGIdoTjyJtX+iebhlT0KrZFueWmPJubjk4fg4Xus6aH5usAxqYwFSJJg0zuOcFo5
Gd5DaNn3PQ8ifXayF9hpYHTeBxOYyXjnTVd0GqluUKCQtVH0iyBxJyC4NWnVz1C+7j+blD7gcZ6s
OXU+JaunMpyS0uxVmSW/sYdhpB7zDU8Vio3RSMKJsLJkkIdOB6PYJ823VPR32/WRCxlUuwFBS6c6
gIFfzkvUjAoTH4OAQsgeWzl/N5aUi+uTzb/0mJP/iTbCYtYMYScedm33Cw3pbGw3yzXcl9dW35Tn
eg4qD75AF8gm0XL+lIxsGILZaL6prZ12PKnpTg5gg0aU6djbvqEY9cSjhbmac+0KyBsEjXjW0yL+
i1TiKfHwRPAvv2ZfpJT7nOjUC4Ri2MZGjAzmipcefUGbL0zUJ0191nI50WfqYUA6iP6vG3VXBLLC
aIv9Oybvwuw3IyvtwT/IWM0NYHjaMBzEoRmIyGcWCVGRUYax25RsQaGHDnNXsObp5yUZeATjRIjK
WhBi8sKp0UCu2nJR/AGUrRdMgjcek5TC1gIO9t9wn2RqrKGewZ4rPQPlk/dDehH6gb4UU4rXz/Ys
CbhODk1dK8hJxf8Atj8w4cnFB0C4FVXfvbIafJ03YdjqZ6iT21fqz5PxvPrzbWubbxldCo3Ae81s
7kHH5/9JZboxJjW5ZMriTEo2HxCF4NTyEpwV34jvFy4rOzR/DvcKoTErxa3tL5sk6GpzxJ2MAQmi
EazaBx+Ab3rDW+Z8gkXTr/uftUaqb5gqm2y4hw8nXgElx3pdtUQYUlmVicjPFsN6Ku49uBpRnaBT
QAwDGb7NMyEJrBnIXPWbur2ZSgS1owPf4NJAw7piubwC9zakksGCP7DFV3EFYFFbpL1c3OUMu8TA
Vr6g5RzPOFbUUQUdkufjLlxAVMXVbxCa6ZyASh4ro5mIiKp882OTPfw7z+CLmkCTKrok0XaWDRtE
eM3afo+1a3WFILXuiCD208MsCoWIi7jM+ppLalysC/gB0h3vg2V3uc2bs0VJjZBFhCpUKsqlihsX
OJXMCtSGR0pMUOVSqzLX/Fy5kPpgrdHm+fIKji+KZo8mboLKVZYj0FXvZu8hK+hwOXC+hjmxIZLc
h7v6UdAIs3uGgARhGvFO/ctsoZLaETVvDnN931a3+wCye9nXFy5aLEqQFyjQHiSRqwhnWGiF7UBt
3Dp52LEGQRHFaSc6+jZxnQMexuxVyE910iipqCj9SFtQXZNS0TfjJqTE7sqHQtQdRBofmNPl5Ezu
levSHv388MIVotJF/CgR9yAN1mW9UTuVC/S44QZbppdpPs9Lh6aXRn6UFvByO4rNTxCELBgVp5Yk
f60CxNuQ2SE0cmosenye+npGW0IHXyfNNVy/nOu+6S8G+T5PQUizMjRg6HS1D/oZ15WNK8KuxdWi
bH0ObqVMIoG2NbKoODajCUe9YUQTXztvGh+T7tRA04mHmkW11THAEW3tB9c6LkGWGbwinOnYSVsM
9YH8QrYm5mIxObUtL4O03Wd2PUphH30gX5KN82Xzjv3SjsGFH8+BUl6qyUWoHcl53RmSMmROnX+5
NPxGr0ARNGmMeeQyXkULmDsWWyp8+5Z2p7g7s5vDT3JsaIRTzqafKdTW7zLgpexr+gPiQagNBNkB
bZi+17jLlQtjc8jL4y+XvpWcsa/Odv6Q216+RaUAkhmClq2NAxObiASJpRzg4Xp2123+ZT3TGKWO
1D49w5YaWMri6gx5b1C7abvBKEO6CN0iFswE15lvLXEVOLAvmG8uwCxhdHzt5DAI1tkAJBoqBXeF
N+NwLqweBTYDeOD6q/8UQS8TbS1QUfVS3XyrXYqWztZ5wcDH7Z1ccVRqzeHtDKfP5RoEQ7SeTz93
mQ9jGzmY7QvtLJJnjJD00AjuTofGpQ4FOjPFGb2H+LJvVZy/ufGh9EVj2DMdp6Ph22LFG9hLB2tz
7WxccqD9hhGjcTHTPL/CohjNp2DAjjX6e+hVd9Oie9zxNeZpdMaTYXmT0zsC/l35p4OvWWiRPUIc
fW6H6xqWgTZC7xzPY7zzpSyMhCLpdP6ogqDiRXHJ86Lw8ZITGMiOxrYSFGPueNdfDaxq3fXPOJ1d
2YzgjAR5oQEfGxrQCFmXxxYS3F+8zHaW1zK9zTDNoKLKwqn5DbE49AtLh2XKmh/qvhP5c2qYVBJ/
W4siqjezj949BYfq6RjaTVtWmtRaWfFBvhUUf1R8ItFy7oXyWkeB3RVvf8LBUEty+pvkeIeI9NnV
8PgQD/uJKfCGG/2bkiR0d9K/Q4Kh+jA6X4BDLHQoIqxmvdxBkKVtPaPl1b4AfHG8/f3KIi0N1uRJ
1Ey2ziWmU8f06E3vALfv7D71VsKUUrelrzfVThM/kuXUHkw6/FfkGkbMACBn03WflZjiM8zOkOjX
K74VWB8JSkkfhMajg1PFZndgCWrM1zxp5z8dyegZJTNMDaOGgqdjNBwMFQLlBQ7rro9CFy50tNzl
y59uksUYR0lgh7m+fKtXBx28KUHFZKusiNSc22CaqKoZR4Emud0+lWFjrneuiudi3vn3nZXu0acj
jm+fZLWR7Ze6MCMNll8kWOpB5BgJ2Xc0j3Y/gfqHORYvr9DPJsGY2jvwiPxp5j4bh/6Yy2dZLzBu
DLLpfctsRBTx0HF7d91uvLCu5TzqPswqVwWCdqRnf9HYIkWiEeaWCPP8r5QqU0yanXq+ZJFBsI8n
rPA1LoX8bQuJ9wWXk27f5YbpLJfVoQ6kuUP7DdjeZ26JECGajHJfhQnZY1MkIDrTWU8kLW7DiTuE
HpzvrqGU2M0PxfE/sgJ9yC0NvfeuqJCySZL43QFTkbOohqSCFw1W9ML9vxECp4RXIRjpGXOpGe0H
mkvuwehyRwWciq7dVRaZJrQ9tZp8RrXgtujzOhAx1vc20fCw6+V/lN+F2NcfIho2jrs8LfnUZFjn
SyIr1+8zMPcQUK/gcv0zdRwotw93gdQWyO4HF5qSjosHeBETmCqDFb877Adu13xPwUDIr0wJFpXE
1le5WoY8whFGRb/pEoOdRpckZO6LtxHznWcERISuJD1XfrDl5+tY9KfURixHNQjBPXFJAgRBHbai
ld8M/Ec7+jwAuFgOAADrcLOnQKsCgTua6c1qkWI1DYY8FJ++Koc+FLx2C0WLwVY0T1za8NvVU8yg
us3duEQF5bVvphNBXf2XNMcMAtlkrXHEi/ojRqSrBgWek+4nmimuhhIyKtquiIEqUyI8CyJwQ3vf
1GRIaCLSrAEeMBRceVDgss2MCBvmJxmfeW8ZzkoAgEDTMQAWuDSVZAqGHbQkLpaWGdY6oNsYnHuL
6O4XLyPZLB/aJDAVtIIuxdKTY20U+PSDdlq0NFv7ZYkSioVCUun0W2F0FG8DY6P49+hcTh/V2zvv
BMM7sBPwd/uv9LIvTBw40efaBjOuq0ShnKiEWjIqdrLZvBwsQUlSpdfDzsMJgLlx1p1vpj+lRwIA
e5mZM6eOv0mqBUogTfGlliXNqxwdeJbfS9TTeN7+VPieMGN9MwdwEhmlOUKfTb/MLI0WWoVqolgM
8C2s/swojSenYiOOyiOnr+/mc6z/Ji6WVCsISP8Oqz/Ilb0q2IRi1VqLmLh73aO560uXLR8StWb6
aqcyMaSq4BGhY3CQz+zUOSg4lhaHatBliPn7jzAPVd7Zwds91I5boZGgdh++xkpBKYs3qCUQfpt6
cKl2XTv1i6VXbWR4SMHHy7MG+nGOEZCplRmqwW9wqqKfRDkeMkz55OQa3GhbiOUVVTVKGwnbRIDo
nY/DYWF4zihNRexWw266wi1d5AQYfxqKv+iRW2O6ta8zzRU4GQRmE2G8XahzS5/nqHhbeI3TEJzK
SHya5Nd+7VdVrN04S0poXBh9F+WwVBIncLjP615qPFGECma2tV2rZLsMkP8D36GAqYvpL+TDBRj9
9elMBbbUyD1TmfJzRADpq4VyWaodtX36B47xm1SNDt2vVwEbL4nBPmIv4VuH9+YNKAtpG5RxEXXg
1YKjfUVltgQ25v5aveG3IBD76tDjVQ3YpAS960mxuPG4wyurIGXdc3GdotDS6+/qIryDY5Ks14j6
ri/PhigphNgU2QzopS41R+E2kQp64HQTNhWQSTXniXlWI3qBwlsqx6K5d547UldyshNT/+mQye/z
Ferkg/myHCbZHijVP9vuBfB5t9juUhyZkCBqWgnqe6gnPIxr40DmnFJbS/o3BqJy0QVjmsXDLnnV
idIfztB52/ccrTytM/6QzSWzzYW+j4XbD8ffzYVzfrgJsZzTUIqiJuIw+hu3ati75zflLBiwAjEW
kxJMqRJ4jV+52572SMebLibpLt6lV0d2zg679Qz4+zVVAd2UJurxMoPCsEgdnzg6Qy+DAwSyxypm
jdd3/aDpcR7DbjBzzj4rwQODsTfDAE5ekXocwLBbknh2bUQVq7PxF3uW7oMO6hxMPCAOqbUdRMSX
klMy0sZGRO6TQAVSqLqeyrAWMAS8w+LbXhy0ISvHEhR9p3Oz1uuA813MqYWp24NIHwR6Y4PMhZF/
BbN6WsAeXM/Y9wRmOY2eSU5Y1Ki8Yy1AVsU0H8ozI1KpmAotQtkdvIorZUbhELOEyHJAAQMx3br/
KmIGW5rg10604SOH3J7tHS6V+FJjoPrjb12/41GkhM3DblqQ3YthNhrMb4h6b9YOWO7EfzYVgNq3
3O6h5vyKDS01qexJgtNizV9XcV3CDJ0YwBVuVHZbj2LTsz4lswmUd4FXdSVrJceARpjwOzC4/45b
eF9wkGUlZSupkIhuGSIyyRNZ5bQdxfXtZavI5ydUVx0tsLXbA8bp+zHMvlvmvPPypwKBmZgrR80O
+Wkx8jYp9DZWqI2I9w3OGP1EtqoHbXRAEaOg1cIrGXiYXIi93qsmw9Iy62iw3/ySojjhYluC/E8o
qowPfEuUTYUti3X7JxpVhVBtZlsb3W9JCfmjgcVlyHQz64q64LjpKMI7GOi0lUGEdx6Pnt3CGwKx
6oDksE2CTRtKD7hSVsdeB0oJSHIjG0xsHubDLLlV8Xdh9R5jiwi4grskleOJ9+aR24x4LEOUOLkY
Dx8mxXwfvVzrJi1CE24pqlGLZXdAmw5SiDgKz+CjnkXy+8B6LdJ4FjIhu5hmmOyB1RLkZYRHlm/Z
VvJHUaWRfvKg0J0cFFZCVCRHJAWNN8oUY/oqBwEsVBwmDErDWVllx2ZFcKBIwuV+JOytFR4pyGG/
kklU6vDjWTrLaCL2SgcSlhoxhIjKLbZbORZMwd0L/m+CBGSrQzmOcOmAZMurhAsvDgqywx7NVJJ1
4sVBNAfkUjnkuufX9na43//HJw4+LLC32bCRGT9rUAoAncfX3tmnq3xezCwawsaBOeoqgr5dGV+y
O2zgIvqvVC9Hv2kbUi4BCGkLs+xoE3MWmCQ6haPuPfd+XqwYB4tOFxFXnZu5dzZ42Cut2kCPgEus
3/yqN17XsibJF8+KD1gR3jBX7h3Hf5RcLbSDxSSotGqJW/x+nwj8kWILhAQmRQq9jFT4+kK10y8s
zu9GnymrAcY4/5Fo9nyocOYZY64Gp9dDuxZMlNlSsCorO8bpUQnD8lGONuyM2yOWyCd6Fez/Z7PS
n3/iXxt1YlePwW2u6FAm8mP7ogIWeKpWvLtCjdxX4kDPBxnsfdKNpg52RLI9tdq0S8oeuW7T1mcs
hqC14jHJIe4m9blLXAABBf/g2lBg5BDr60I0Z5hDgdG7mUm2hhs5lw96mXW3lY8Tkz0A3l3xdSCb
y7IhEZ9ALp7Y9noOnKvMwU8SN1WAekzrVmtTlB7vNN5ptFz5hrn46vnpSJiYNA4YQ1m3Vt68GF1A
PVLTTjYBuVrcyfDSkguluZ1bfaAQpshzFMlm/uOdy7/v9MHD4uMH78vZlFlZ/t08XSaIYuWCt690
5FavfdP+NJEdwZSmdfXLiPWTqG6HzncTC/JFMMFPCfmnLB8cFYVUvP7srAyJnNKoQFBzHUgZbby/
F5o7auVWKcprF122eYldlAmmJ8i6rekItR/RjTztU215FGuEJTXpBw30nyMccHyG1RDsJunskkFO
sVMl5k0MQ+bEqiAEkotWrt2Awt/vbAMOl2lnX4y498+GVvLW16QLnYUWweHm48t9jB6SNQsbeTf0
OLR1jx3b8J0s5IMkM9DfdxmIlNfMfJzX5jZIc/YmbvP7+UJFMakl/6p4QZflEm62iYdoLvJqEkND
2uR+04C5+xHZV5KIwFyF5o3Q2gtCk4h2F7Ro02ohZ/UiGNgYuoE3lYq++wRbA03BX83+HDfvDteX
IrVJ6Mzq03hkZns7cl19dK5RKr4waVUhF/WhU3aNgmLWKrVeogbrpXyw3F6w9Eepw/hQrBUfF4Zb
8TFKnilU6aeD6+sJALB53Evq6E3TfkQv7elE/Dz01yvS/G9oiJwQPNG4uGwaw3QJb9Ix8yZFpn7w
T1w6S4rILB2vpqhsqJLaqbGLUWES5Q4tmnW9gEAASGxxvw8fSG50uBU3dEmW8AtOWkxV0Jyq3NNq
n4mBQo+Q4Ca6QwhBNJpuDi8o7KV40rMH8P2SDF9kFeJHG5IEl/79dQ7pJnM6cJ4hh05nx6DpPT5K
rTKKjs7w78H3qNkQ6Y/XhjpYasM7T7cN9ZYFyDXvJk8dtfA8beLkWrnzAjUDpllEUUiNDXNQsOR9
EEE2EFTWV7HeH1/Rp08wCVX8rU+WV+pUvtlSYWuk2InpRVs7YOZ/pNyy0RrWrSFulu49dpXTn5Vl
JIuSChFM/nvnr4Pob/BBK1ng2tLIkIMgFd3TUKAXUjOmYijjLx9dVkmXukKZWyfhlywcAhxcKBi1
IPT/iBqRU1TC0PJtLuvZAo5GvZsAumkL0HlxvXWEJU9M/NUSIK3n4M/pDuly4oKlI+4ys8PjC7ql
YB5Zp21/40mC45Pfv86ssBnL7XL/4XRHpLz2Yv2HhyhEgWbway1PbgSu9NzCYJq4d1FnZ4rHFjeg
q61PY66zftEDLd4m20M5nkWthj1DVOVxlicl13SlSOrQeSX0rFf4SQ9TImQGKPrlYabVIIIAHGkX
6aj7AbLx/yNb6WWNXVe0WXa+Kw2vBqQ5m6wtu/xkp2ae9223t3FpcSS1zECqva0Z2iCHa6O9y1ow
Nl1Lbqt3RmWdNCoye5ONUq7ml32cuhHlhqNqd7K9ZCAk0MactclGF996gANEt1hO+8EazXjzyL8h
qNk85Eth15+GjymA+EuQILKirqpn4v2aByV/3GBh5xECjcmtiqeMa7VvdVGu7M9hlOy+RoeUAyg/
c17ynvGrLRh7sl6BQXtvHPKHjaRdH95rRiuF2GDOdZbpCpt4O+kQl0MTZfamQBoFSTDQO1Euqf1p
O5NSU/264Gl3ogiq9Wi+2G+ux6R/HV+zYdTQjveYBJ31X1m3RX0WmyOhvAevLBBxmA4euYyS5+Up
YgmLlbjS/oqfP5BiOMdtNAC8FRhCFvYuHcSfJHBfT9lKrR+0yAHf/nUfmH9aQKmeeDmMVWm5+sS5
jp64LffrVWSJetlxAIzK9zwOuxI6CBcm8xNAtmWp4Ozf2r8mCK+tJ7jXeSzoAXriVYzBBN7vHxX8
7NqY7sB2hjq3nbJcaM08Thro5TT6w/HJnFhsrcVc+aauQb0o/7D+RfkoopAKWLzew1spuCMA6dQe
76Tkb+gbNUkoFynYhnA8a9SdCq2Xau5EmHLp6RlxcLx8750T1JrLLF2uCG9rqh4z6mqSBxtCmFQ2
CHO580r9deNr0lKFpXUq6yBkQIE3glCBv11AFaZkS8uVXhvnH3eVGDBKbW2ukmhVYmeJWa9uwPEY
JcSu6/8kI1TdJQHamp+lS7/k9+lOEfXNnyjhwajJVNMfvEfY51cgP0VmX5MEoYV9qgetlgkJ+Dto
8ahRQelhWpC5wyEzGSTwFNixo8xhPRNBJxqpy+JTiQBQGKkwf2SJwLLqfx7PqGgH8/3RlVK6LH4p
+KxlJMI0r+pUrGcbpluRj6+eyRG+4EuPrYozZsqbqC72OmwPO6ge0F9PE1u9enOnVc2l9oAFnExE
35Lqb+3ecyShW9WbM4IbiQBZ1OUPXhH03fbS05lNZ3HMzgDe2cJYEQXAQK5Y8meKW1GVBZDBy6De
N268LcZOa2oHseb6GtTx6cdGD4x69VwH8CcxB9Z8czJW3Bx4lspFtESqS1/0uiRFYx5wvs7EgQ7c
IAP/i+cha+xb0YdiEQ3aCzPLIhGA0FvipwoZWFAxCH48nQjsSP8SPYqI4Oa7mdb0uyVVbexYno/G
kGD23LQhnIkXzPtVllcD/t/fG8hYiRXA3Zldf5EvJ2MiTuavikehB2CBPHjuEdlgXiAPvZVsrjAJ
2taDp+NAeGo93RZl9ITSblbAcYxTjR4BfMG3QXp2bXNxXJj1T11RPuRaVnh3wnPgH6hVspHAMUcg
XLfYec/ICzHh8pulokCwcE6lkn9VU1AuBjyl4Fka9diPxLQ/8UNBy9llXbGfmLqf5SMixoFQDTYy
R3a6qdNTAz8gV8fELx6ir1vxREg3jfEnbyTK/ppyf1LCwm+WASf/lZUG2rSD3rV4FBzfdG5FNgY2
FnB86klUzU1uxd2QB6cPZ0iNbB/BqHqcvpRm/qIR5VenwG/m4fzfkPZm6nVkPP6npL7uG4fe++ss
Eg03o91+eLCLzt6ZDWAF6Z6tSl+rfow5HRH271n7SeYA2/wkVGyh0wlI2mJaL5v8SWgcNFv7nSO/
iYQMIA7haVRd+KuKbbplOrUCnJB1Wxpepsg/hSAQCQ9+WhRQKLbhFsiEELJemeBddvvzSNz6g3CH
6+bIORomSdhUPMsLLaHnCkWlY5gLGf9OFvw3skXDWlwcYz/fHTkAJH5XSaJlS2PKOIR2WRqUAvXD
YKBmxymJSiamtKanrTXLN1v2qo8N3LYP+AUAS93msafwC8mRVo5yPxpTvG6h12D1ZrcewjmwwW/c
7b+0mZrtZI0hrrz99Iq0oyjxFZKhR1uyOv2ifb7qcc2IeQnglLCdbfg4XUuqvtJBOjy9f0Nh5d/U
KUPjvIyoTHQDo6jUbwItV5528olP6vdnF24HGHsownZjvcPJetQk8AZIRgkln0MVfgJnFzBcyt4G
UNQ8INU8cwewpIGRDFx3NN0N30oJQmSWwIARUr4VLDDopYM+jgWZ8UZcb9XD4caG5hFxX4it/Gso
KnaAjDtbD6ynvkEZHUQL89CV3ie7Tm99Z8yB7pVvgI37s3dSb90MieirBAQcUV5XyPEihJQHQkzU
yF4Z1oqWpbG96MFVq+qcGbFxjmNOJIBXM3J3H7RxjixHcBSlGWmo4uZcAGVYBvLWn7ib2OHBpJgZ
TRWxJX+61KZnC5v9IbR21jwIbS05ETXBRd0cpkvTDfQD67fX4oJ0jTVVsAauYQuh/ZEvuEepmX5N
5U9NHpQ6CYzN40pp0u0TZ6Bb89ch9FOm1lguScf+vZOCHqVUSrCxpts5NbyvOj6KnGCpAhu0NA7X
ItKQfzP50HkwqP+2BI2FetQLbB4Pc6947gzsXr54Q1IjBpb3ebpMR/UH7T1WTI+n29Pwz/6SSo1j
CmzatYToe1CkBsMXgXVQXNQy3pBPwkDmm243OV3egHQkt7V0NJZ1+FmlyUqzXbMTEMyC4aEXzLIa
GRuINU3tMnStN9TsVSfzECSOY2UUcnKupq46Ahdr2XMssAbLArzkzYbuN6Zb3JHDx2MFDa55wEiI
v8IPuQaNWNYWnEMEPjivqJUBi4ttHzMQACURPMbTwHqAo7TQJZjjM8N3DtHYWNGJnmUSvlygmp1i
6k1adFQAAf/dG2vRFRFtP1UaBjU4CYQpNhzy1rQQTBIUqb0isEweJS9mWGpxf7EjGC7Xp3poAzyi
t/Pq3dc9L3ZDqt3KNBFI5mKoE88/Mq2iKSzKawe8WSxeGusJGUvoHbvjV2UVvr80Z1/nHs3wqSj4
oTkC83fA55G8zgPZd3e4B4wf8hYtK/bHn/KP0Prgj5WA6z0AUsei/30FJuOaadFV09GzeRPwUqSw
1RxDgo18VP85LQwqx6unYxYpA9sVh3DmlyuWuaH8xZQ78LUTLqaJ2cMxhEDqsCXFBT3Wc7hTXvC9
muk3xOVsQYoxNLfsbueEyeL9l0Y8+B/FcRrPuxxwPE4KWkYgTDtEx850F6z/6ASp39BTlc5coEf3
2pfgppyK+GzU04wAOAvlzO0+pLuujGesCmeeGP9UrR7LhW7yyHtoqCNcFBmEKQB11M1M7wuojU49
ZKhFUzg0rVNbcFGaDmjQ/sjFut7FPrdcAMmHUJxmCslKCapNW+j5iyW2zNeczs9+Bo4u7Udp7E02
LKmJCRShuSuNB3nS4kywZm4xkcMvhwJGC8erL0gd6l/LbYki23BgaBnBwuXbN83bj6C3JIx6R5k/
3NLvlVlJ/PXmQlsJe4tAVT4JMwX06+NUsAelwbn51WbMcttFTRSqFDXnmsOONFywtBQK2xo9/yKL
538lFBSFkHEMXDNFEQtHwhTue7tOCl4G5BbTqODcs/rpk6HMA0GCiNBM7OZXQOVePTmdIcOqW4pV
ADiknD4fHHPx5yb2EkeYXuGpR/cshsDfv5wBw0ACItfZR8XmTI7PwLkV6YmCsnkbgOOgti90KM42
two3fNwPOTZ+GJ4V72O30DYtTORR70uyL6OdQ1Le7s2RjPSjWBy4xhqpJ9LHeW+aoGtmf4IlZIwe
QKs6K9Jz5l86B0QkHpa3/3V1OIlCECkDn9a4v0D3cClMO0UjFcUdNmtOJOYjZ5kIKPR0dthp1GNt
d5jOP98aoLjpLBVrfWNI2QbMl9114tsbzFUggx/eil1Zs3PmjSCHugydUbcvuqN5yju0YoEX4oNo
DwiUe7d2vbFgC7c+/f08Mw9zNElG6j/1liqCrTaf5YC+BIRWMA1wibzoC1Nepo9xZETdnkGO96MU
pdxjqOeWzB2s/8G1sf8+GzFfiW4MMVbXiqx1DGokQD1lq2aqLILsguILf0pKgeIZH1baaH+6hwaL
7UOeR06I/rIhs7xtnE2hho5+WWfsd28u8eOHFav0son8FqQpBJiVsVyJQzk5LhxjU0TTjFz5XNiA
qvz6eSWV7BHx6GWKeThop7gImXsLn+pFRxuot+zG3F5mg71S6lLgWY21PyrOblBgB949WMUjo6zd
pz2Gg9+KhvpMtemPcZ9rXSzPQS3Cm9v9a13i7ZURKhdyZxwV6xb5PdjGS8bbFVlqbz/RxovWQiE0
oSZNTjBr3tj7ZPsl97Hafw/XaPu0ltgBmXbnwAx48KQTh/llry/Ap0ICkUmO0gFaFRTLBtIPBCue
4g00zK5NLeyBILxL6ecfrQWnZRhbYMxTNsY9yJCI5cXrloACRPpvM6DAXmzlhnJlI0+DwN8rAUaj
UgFVeeSFwixHtdL9/HfcTGK6ZfVsSQb+/qUXDlz4NRXhMC6W1bDueqXmilq8jwa9Hs+zCtLQjVER
LVXaPVq4Cdn61MOd09w50/U6OF5uMophGkOgvM3F+X8ltM1bxu1GLyfSMRs0pzWZ22wVihBDWMH5
+szH7k7N7K0zivJqwIPbGbVxcTieaoHZtJQmCIAmU1imPwlmb9eeS89OwC/iumXFYsq1CrylodlC
f0eXksBJLeuNEYkzZJ7KBkbfKYQtqkZ6pcTrTj8hi0LsHlSNTAl3GCtgaR1vVCMGHgG6yAhjoL2L
Z6NUwPhgn3ShSSJhptYN7jHRLrGVzx54iFIOoqFYw4/j3h07rioquaSoaAjodQiVvJZA7nwVFiFb
6Ia7diM5x5ExHUaJA6J9zVG5DumIaQgdUuYGZ03qq4ECDbpnijP56ssPxGUa22r6T/h4Na1Ho3L8
oNrQ6/1HrAiRHmsEZSoXg+6IpKGX7mqnHBds49pN5p0a/F/HdqCOk/N/q1VzmyHjU4YGvG4pOdSw
YEh00wbrxLcTLWAOg28y8ql1snrwloaQAgDil24cM9faVPsa0dUE/lumLSZwd1offD36Z0ac1wX0
n8h8YPjAYg6ZqhQ7S4VAER7JDrQP8M3O+TGTG/uLygdQlPFcxEolGcTha5kDZ9DraMmbLz2WU5gK
sxb4PbAdGa+rW+H1m3dZeqqai9mQKEaUV0HmT6y31zLmDBJU7RIx1dtX15CGtoteu4A6BNqUFx7K
UentjXDTHWU76fZcG995qj3FRhOQ38Oj9FnVE69QKIyHDVFfT1aQU/LaTFAOD+J9RIb5wYec0ES2
v7Rj48woMfYUiNPDGCb+ZtSV1r7bYE58aJAkCoBdKu/hLVhDmIxnBAnu2zpcYErlpIf1JSFXK1Ap
qjhy1M/1PtV/4fCkE0gxIiUcNw2KhbOx4HI6bY2U43EE/r5yCo6qPOYxyARIcWI7mXNE1aWZQ42I
OxQ1lDHXUrnW3+YbEspBkf5+EG3+LAGC5zCQGWP3UNEdWG427R7Z2tnhdMTqVZgnK02c/a+Oz1V4
CI0BNkyKBzl1jKwjdHwqx7FJM+Jt0FpVBGR7jxDw90bb/ho5tPL/O3xOT80iGwNiAE620uRCi1Tl
cuMZ7sp/6sbBLa53eC+6R1JDtf1qowOUXa3ZMyqMBO/fOPbUgc2bT+iSVi4ICr8WYeHvFXzs9L9p
tD5cDLhGfK4l3OSr7KEBnHJlfvKy9V2/+rcOu+k1oH2htLe7cinqVadX83AsA6iEs8Y7FhctgNSh
VzHgtiRmqfwE2lhcChOPdBJmcpO7n38IGV2g3MNO9OG+j42m89hZFSOkgosVPsJsiHXNqjJYVg3r
yYB9egG+5SNfXPNyXgtVH+A+nC8FdTs4LU55WRVz4MNPCF1qp5YwzMBO0IW9RbwRNTZU9xbTBOSK
Tx8dAAdKo07umtU6CReGu/qXMukyDof1Mvjl7A2D+ooB6OHVan0b1hUps9/Kq+ppGigB2SzucxFw
S7aBFKHhMULWHG0XSnVWuPmsdKNABeca1mv/n9BDTlyA4fIDF53ngCZQwAkXuwHJRYuIb5umi5su
Uitf4iwv+ek5DcxOUjwTO2V801pdikjMhDGC+wyCBwZC+DUPbNBLTFPad6sDDvr4P+E6wUR3QVBa
jUqlb8f60uL6Trdo0lc8ib4Ssc4v6rd0SC/S5wbOY9bq4a2cvPlrLEa4yUF1hwCvx037vI2J1lOn
vAdhgl9YqkmY44Edr3VZ5Q6phaSONlol1jSAbv01vMfVnnWu2tHJUabUtGNQROKCof3kXd0wmBgJ
kodfijQT65iR8Q4Y37W6OC7dEMAQHpk5m6nIIKHWglcBKb2I2GXhg3JzqWq8sJPfFKxwRS8An2+5
kQV93U6VhofzlsnLgpIPdT93EleTFnfC8P6FcEUDkjONXbwKdTyJVMFtOFtYvhs7gKv9xRC+LlFe
JYqE86BBKxO4bM7EnizeiYGnRZgTmQnuPGPzD4qTJPrwodFgbKjIWw/+hmuNdkp8nd8GONQielB0
XwoiTFgpJlSe5kjC5jEzRtSrSvjtrh28k6rwrEw0TLZv4PQLlTGQfl6mleTbRzDZzaGxTIVJE7Nn
IHG11/yRrQpm6TU7pKIGgBsuvZyrgEmu3HVgeC5LPjRqsktK9ntaAyN8HHBf+gYjR/fD1srU08MJ
KGQH6IwyvvKwVRQuGoYDCOPGgE9SJc3ZdpDtaKOxu8/m0senr8omZr6BrR4TFBx0Dup+slLGmriR
W1s9erYQgcrpzowU3P8IlrZAF35NR7gzbvFPvC6p0rVoVrqmHpnv3q1h/qBAyitmKGbUBHTSU4jD
7SWWi3iIbwCXpUOPkdALrCVF9BhKLwWXu04RyJth9aZ50KxJ1pLsJmWKtDZWD5TKbD36DjtlY7Fz
7sAbBaSUjnIbad/EctA8JUhEjEpVyOdn6sN2vrf7w9emrFxmtd/xbcLVpuSwZxfIitDA1HieJDra
TpnXinN6JrkQFfVqZwYIjIdZ6jKOLp1+cP+L4MIIKsCXZIJfwbb3wbehcd36i7zDVsMyOeJPLpQJ
ymp/5ObVfFJ2EvDhriOITChgK9CKTGalekrv01A1z3+ihEx/19v/MXqwDPJfrIyL1z/rvzSEKyut
3+jLKcNRJwsmdFmTO7HbUpD/qnxfcIr/xgWK7z8bGylKWl9UPMUXE3gQ9MbtCerjcLKLzQFtZOO6
jHHPxkQLjPqNqWJx9a16Ca5PBlm7u31fivqThm1dQLkgescP/fyo7+XTYN9XBfNB8yQHdQ/FPVBY
nt6e21wIrrfWADRLDrPxiW7BTuWPAZxNcahuEQXsQx/VXfs4p2ivhZBIZFq6maCGPbuWJRqYRyaU
4nYOcLXkZAIlMrSPkyl3zrBrJPPVgAEdouBROegNENLHiRz19ALF7aa0TRkVZm/Fm+yCMl1ZCuMM
uib5hcZNE7vqFl4aATcrdqxm8quE//gewmcd10ZlMuNZ62K8QfO6422YvwFVQBBoLPWIFIlYxfwc
xJ8HFVBdjswzr4yG9GvBzITm2DFR4Rj75nlgtw+y3DW7zqMdPZFWFguC4bZS283mm4lAvL+ZIz7L
0LcN0/Q5CsooxtPhaHNN3PCocP35q4F2ngruXtLdF8+aiV++8/CG7YZX0A6DNu/ufceKrbszsB2U
unFV6AiO+6pPVKVPLUl+4/mKnGUEqudhENzMlVHm4k00iJMe1d6CVXW0U25T1PJ0bRaEfOAKT5YH
CjTxsz/i1ROnzMldfOqSUtzo2EqcY2W2n3u9Hl0KMDF+fEt4cSbfwz4Yhvkt1v6j05AHzLnJc3UJ
EtR/1mXO/kg+R0TvSCx/Lfj5op6lfojRRZwJq94m2pkz94JiqJ8USEmbCuKjapTkqGp+qhF7XFA4
+AzXeif+pOUxWj+wXc4g9otPaRJDaQBKp0c92kBwJCgtCd0rHd/AZfTn16+N+gjAsIDiwfBq4pbl
W9pwp/zVhDatZuKN17tmIvhPVsSvOFiOP6iAzh6seGXzJwkwJF6H5f93VcJGK2M9v2Jq38uzg6K6
Uy+YBTLagS3oVxuyfZWtJEOdSW6nZtggpmR/JsNnvchOUUk5nnyyZnjc4Ryjwhm3l9HhCdsYY0IR
WW22U60CnZh135vUSi2+3UqJE13onLN0quyXdJG5FDEyeDol2XL8w1YfPuk9BGbY5SlUwHQ3MGQi
ypMFG7YRwZwTpKaa9el9uu1PIQd8EzcKYuIS0RJC6vdDb8RGUXobW/1JhXsf3Y4zXfKOlQjn/Tij
6LHauo56F8/FZMvmi9j47dMaXu9BjbMLQyNnLuSVOW4QbrLdE/v2Pa6nR0/A+zzB1JECfOC+V4UH
5Bw0sdxuZ1VAcfGTMoUA668eqn8WdaM2bWuQOTNcrW3r6BLY4gDo248WciaVEhSU+xle6JJQ4eEg
ejqmGIF79Wq7h4YvjbDRr1izRPiMegJVqRpR/paFabIfONiAIl4KlSZ4FYaiBVHb4GK/GSyU9Y0d
UBeOgkuMii+IBTnupawVJ4xFjXbeykZZk5pDFoyU7JGp+WNx5pXR5x+DnG/+S/0zutku15W+k2NG
/tuSCx5OK67hB8MZo53SgtzK1ao3Qa1JWpS82OEBs1EA6Sk6zG8mZi5/revQOw1imd/PsU3MDe5Z
/pcCyP6e4f/WlbOuV14vsyXZgkfFDZsmZRTGBhMnjgd9UMiwW9ngUm8ml3Q1Zax4ei6ICw0D1Wn/
mzizgCiHPVNnGXJrngRDgFCOfiNvXvtmedngZs7/wK0WfnVOO5SaLxCjen6yyFJyVY8ANL+x378A
XlbOUrIJK/SBuJU8PklR81jRoZk/qvbNL0iWKfAGV3vWmL8/KZQRCMN+gO6uEC2Xwf2v5RIrgMWG
23cb2ow/jelVLHvpyVT90L5Lp2g3OWA509qliYQad1Ut2vsIZjYlKm7bb4PX+qAQi899TsCRROq9
u63V5aJjPvh57AkH4Cfz/RguS26CRcOdqYZx3d50J88sjFcJ/86UERkUpJ/YxKtlt9QeT7S+gt2/
rn6ew+EhDZVwMqYW8FG9C4T5LD5c2f8XeZCV28G0JHVfUfYNP565UbFE+gqbu0q7MD6AqVhLIBtN
PDhIN/abOd8o5W96vtMcp0nFXu+7hoJZ1skgEnKv1tTdW1cH7PFMa2dWYtjjd83ikuMTV2SguSq8
+UnQgglQn24Mwy8jOSqiJf8FgWkaFOMISkTLvOOqRK2/mkN5E42xJyxUh7nr0HdQGUpoUWI4EEYH
NPyqsPs8wbdTzwpGFxF1MLO8G/CZRo7acHxhnVF6F1/9Lk2dlx/iWwcE5+JWN0X1KIYxyFASGZIS
bC5glPm8uQYhVcLipDL//UXiQsmyvYcqyBGs5hoetWDcAHSaDODPHcMaWJz/FG5uvSnVy6dMq+Si
L6PeTr4GcV659A2LYNv8/72gFgZqD3yuj2LeHuYu7eV8VwJBVqADnQFwGzfZfg8AYoGp6XvviJdI
GojoEKhZbnpuXxoVvkJxYgALKSYnMbcPxYsGsOytVR3u7mQmExj4wX3RHUhhfWc69ztPcQtprdK4
glGV/mSNGfMc9WRd2nXmT8D/Yx/0hmr/vvzLRhR8QLa/MTY0DpfsGBM/o9XbLLoRHOSqVLVM+SzV
nLi0AjAPoMv3L/RTVwAfE8aHEH6xUx4qfs8KFxsFcq6jq1RRc0Dbc1wSOlzR03q3gOgnHKIasIht
xZrvKva46D4pdaXaX2Znk9C6VMLk/nHWMautdwtszkZxgpPlyI1BdzHScMV/2UfAKFgpNLBtb62W
do3z080zPlBlid9MoYsrb9Ip83UzUmvb123OjU16D1sqsCqQ7MPZcVoTSUf8XNv2ZjufKXbsXWBQ
13Hq4roMHhGtm0P+OUX0gr8W8C0qrnVTVq5lYxrY9PqIdbDXesenQgBcZpHe6yrMytJjt+GwhWLL
4kItb0SS2NBn9wk/GRg/7QEeve6yPi/iJVJTgyYwERtGrrr92V2l6jNUoCqKflmLiBP7SL/fIdht
IWHB5DEK32sMoMLOdCwHJVZbbfIubqHI5xXNTkXkL3uMwMdH0qLv8WbcPLWBbefk+t71MYLGp4s8
6SVDLT/YltohoAOI38I6XZ6Ps3y7a72dL/HjW5scOusCr7eMmkm3kECEaabo96O/o36II+NlrEMd
/fy8za9l8XXJjOiSGT3R1gObc3UzY9RRTeX9anykbJy9RX4DoNWmComrGC3xLwmuZLI1iB3FREQ7
1+6sdzDq0kR7zL8WtRwBPT/aui4nBGp8u0nqeDsd/BcoB8R+/IRsTHfVn2h7kcIK6E2cGnejkMil
JJDZZZlppxdyeOqOFhd9WGofXSdWCrSgK2jeUQUX4nPfgnRhQJ4/rylXAJHmZV7eMs5kfLZ9inli
dsA/FXPMjlHbOEDokPaG/yq9m5+AH9cNEZliFTyfVNxpi/PGm5eCrPCTF81iSdQt7th2NQeu+dsx
Rmho4tCfQ7kQmyXHQ3fltPv3nS/m0X29w0UzhTb0PKtvNlTePIW4lyuNNccqA83sc3AwAgwo/GiL
KM2/ICWlEkZe4Qu8PmfJPyAr00afuw/qkTgmnlbxp5gzwGHtXOzKRxmS++qrPojpRUOuOA/jX6rV
moAllIti4OMEEIQfCpiaRR8d1NiJGxK3/IsXFCLM+YV58BHvC3Ef2iJX1sw7gXTzMcHljGHCDxzx
daGklrNJj/BN1dWhgjmrt9KQPPhp/qacR+pdf8vBqSANvTFsHm+ZhCr1Ssm29HEu4UFvodKmiZhJ
kU9v09xr5zqDgG+W0qBT1pxh5IetoVUXg2/SrvPE1EpbGWF5+0J1/dn/cuGe/OAw2qBD4PIqAA2m
lNzecHf9nU/XKtHRw5fJG0Y514FsBS2W1I11etm1MjRjE1A/SehWmYdAOrtKmYdAInLczZw8mftU
nCqKr4WwUSH7hmgB42BG2kxrKpNov/eu2+SPVQncy95Rwi6KXgh+qIiOW2xKHelC90dBplQnhHNk
vsDvHJB5Uzwx/pfA7+LIKWNds6uP2fmMdEhBYAEWUpCZO6O5THov6WcoCz0yS9dIkO4KHW2ITJzI
6r9hyivav/GIxvN/PTO/NylDvUtlPmyS9TMvQbDf4P0B0n1XxHlYQm5OgMXfKDDml6BBI4Gg4vlT
NErqhhSOzMmT34fJYSMMpf9pMB9cmJ5uqbQSxFUrk8xGegPml5FQ6Y9080C6XPa/e7mQwcPliX9P
xyBPVOdCLcdrzJCTUCTSqFOYvnDPY475YI53r0uln6C+zwQDuaFXKACVFYuL7AGpzR1nfvEBqOGn
QpCwfbv+e5rAtbwlArC+1e61EKxquUBpSHAXhZYxaQaAHaeJPy15efVADU/UZQp2FRHKoCXKj3Nj
FUDj8WIA+6wKMLEYka4F8Ca873Pbd8T6jbHSHTrsDSMiXw1vma30nn5FcCA49zA1r5pSti8oN/9V
iLl38MDyZPFrj4c1XpUCIMB/eGAdcsYOBL11x4UdgHot4m7I3ucdNj9ZI4Dkv4N1i7Xw6GSt8mNN
ORWBpygoOhYpBfjzwFdfaZLLYE8LeqMeQ3Rd5AgbgZd7A3siFkHOENOTEfW8ls2p/ARKQHI6NjP6
ZkYP6W6JUBOJJMmhHrqXjFza30f+kRUhGEtozZpCg1cjMrf8WBPyG6yiLZlxuyL9YhAi/S90R2GW
UMWjv6ni8q/mb5d77OAV+nLY5gSEGs9SjF2rnPsYDIg1EaWU287WgrtftdplsufqnvHpTDaUHjvK
AvArCYJXKG6NAPtA2WYnvwB0CvxOfOtOSmpbPrDJoPul/yIkikrOzkuheKwigTI/tqQSrfrl8Cdh
XwCQDWlpDG3h0MekLURdnmSh0IBXh4KPQmVXCrWQqh0nCQEE9U8JOXqEpKvo10ze3jqIXKq3pXl7
XshZH/xpaHFupBxm7vgCOih/MtlzDLQXHED1fexXP1CK5WBsgAXWCTbt80gHrQpDg8rkNLNxaT9E
jN4nvHQUD3H0zWleRGwP6E/Oonrljwyk3IfV0ozOFZv+vosZfCrhL6oQVBwGfW04ZQikjsV5JbW1
6D4vLPixNDZhAVTnlxsaeXo0AIW7Qh1w/08Gy+bvWaKc+OzRTmu9OmGvHps/qBhm+MORSpfUDZBU
m9wwXshzI7rJXeUxz2pEeZFpcIcMShTlCOkzcYSVv/fkMp7JdWF70RijNsZpEU3+36TxSyy+UA2T
QWpr4IYsNmkVn86VY+WY0cLFs+cc3oGxUh3EUfUhejzyDUXfWM1CN6EsWmjVvG5OL8Or/tjcpSSC
qnBSK2MjEQnMvEQ41wlNQLbGjR3hQRV2UhdIegmd0ZZl3RjbMNm7CrOFSOy0ul6u5I6680bYW60U
xnFPiW5NWABCK+lITFGGGTAcAe0ZIWfTNvQyntaJd4pbw9h5VYe/vSVLmoFa0XbzGFbcVObjNrdW
Z5Z+3xRpTfO/d+qJyP79ynYHifOQZFlEIRUTIDocjNVXBkdcwkEYxeMcpHGvMMi5t6qu1LnpDB4S
fDdtDqDQlCGm+3FBpJRJxCbjAX+gak/xsxsriYDJrz1akJdX0rXrINHsLfcKIoNolY1t5hNHJ2PQ
+s+cK+OO1j2pMmksefVLm1dTpU9OjyeEHtyhmoJZCQPYz9OwmXCDJt4yaHmFBbD98VmHLn4rHkOa
mMA0b2V699LtMV5BShwZw+NLce9VJmp2hJ8tu5+jSUPNHAM6ZRA2I/PwIoa7Sbw+o/t06bMhgS2U
eJTR1z+6XdkLBj2OSLjSp1XwygMsrgW5PlOnv6JFPrMkVvw7ama8dDSyMDK5CEdYUeVfzyk1vxTK
L+e+cM+Qsv/6BnOhEsM6YG5ie+L5Ps/2By9XpekPn4Arc8E8TTy2oUDbBjCTesiicSGTycmV8K44
lWkUYSuyipHuRqS/SnapYXGravXxeU0DgdCyb/bxhjtg2kXSApnWLDo0xLhRiaopvbvL6v70rvH+
ocZC9zOmgOo72xpuQYVsu+fX6QbiqQMr2yhpcFnnBWZtK3P7AMdF1U4vbylN5REPuZTDpVwVkP+Q
4JXfhaoWGEoRp+6WPT/hsx9Q9NGcsuuxmzykMANVPWVUK8mig6n+8P10GMCN5aDGBjy/gHHK4EBg
+KtrsrHP47puAZ5XzhsMpz2lO8RkEObJFAn8xT3XI1ISmdYh01fuVyX0ARLt3+/wYE9gtwc0joAu
S7V3NkIV8eB+aWc2NakC10T5I5sJhHzSEoJZkFxFxRLWunRbpgWDoZk4thWVx/fd2gNUqSpbRpMO
1TddIHXV+bWU3uWVU4Ua8UmAUxw79A35miJYnskkH/WC1RQD63D1k5rqaL+o8dzq42v02c02rg6j
XjSydxmStZ9zhKMBxWVRN1CxA25/p4CkInz3VbPZwvRZl5tJSh168e5tBj+Mak8eXglLLC+oraM1
+9GyA5CXg1nGx7wz/sieIwgUsfsWNOCXGR7tOlHuwcLKwZ5UchWLAdChYnVBgY0VyoSgCKIi1w9R
u2jeMQE/m2MOb/iw8YhBCOpfxIlgEjF5xw0VGkZjURJCzAULdpwxAJ5mnjlQpjLlpVRwfLVq2a9g
z8c+fUvBHiFs5NfTgxdl2gxQrYOLHBID0o7QTC5a029Zy4IOsJBVlyaHUs5osZFZ2Pi8UQV5PhBz
74T0LYnL+Mf8LuEkD1+Z+rZ0wuBTh/sgUq7OvW2XTr/9k1hw+l9BwoUcd8OIxaTcoOQX8d7HIlQm
w/YXR1BtBhFojajYf75EYD16oL6sU8aEA4/dksq7NokcT6tgmYfcL7qHFhIRMT2WX+vxDvLMvIqn
rAqlf9ZgIf3JM3YLEa3DumkfeOpN1qE57Io8g6vPv0Lj51Gj0fGRFCnKbbsLgzOw6+hfueMCpQlV
rn6O8/7zvrQ8n2CNk7elPkt9GYz+p/qnB0LraiacGnlRd0TSINx/nR2yY8qEEOk4tx2XxFPW7OQ1
Yd3X0SR8jQTaExLPp+Pu2i7ILFQe+C0Xe4UJjT/wBPpE9eGHXKyrn0c/YJ5dHzMti1z6aAKwweRH
uFx7YJp0kn542OfRMaYFZNQIZ/C0Gk8JuF2G/583JcXDQPe95sWAGDEoXIVnVfL0R5LSafFw8A7e
UpfG79pB5MXcY/RUGqAhA4YJzebFKX7jYzjY523UOLPlMQra8p4IIBgEaAjcAQKEe91V4sacVxsG
hZRFFylxV4BErMGEJB67L7kyi6B2CFiez1/lsDMUvl+aF6N7DM461Pj8XCsvKnhXUUAW1I4yh7Ok
UNKb8k5ySQuINwbRuGxFP294+yIlWltjtOFmMwi/A4luGedRREFO75scVx/wnA4r1E8e+Xlj1p5k
PxY3vrsnETLXzDmiugXg4S5VOV+0ETODw3x3059+R3dD4AXXZAtUB6OSLh0M7enk0//lLdT4UqbP
z1o4NXfWUrBDTXVjJED5pSKSiADgi9ipk2QlXJI1G2p8jNgbZWPWZF4pZLidT+LGYiEg7JGxktvi
fGckXbLggUR0+W1fmV7T5cyDI9gd/Pc4mNf10Mj81+FVAOO3htvhWHCKDbtkTnRzqEjGt+6P2nf/
plTczzrPA9Gse65PKLG14r/X3SAymh70DtT88uDQIO6WJuicjAFEzTiRc5zigUpSXgVgvmrtqB84
DTYCW6OtGZVQJucfDbp/y0xoXWsO6hJYyqZZM7zb9QTcNU5rVzjNxqmuTvg0EMsbisbsoQCgVriJ
lmSeMep6h1S5OFQghrvj/VaS4D1R8ED9qY/gVV+06jolRFN5Fd1ed7pz1f1/bejWN8pSkUs/4/kO
tMc8lHSB1Xm9s8l7yAq42R0531cR6kslWdj65caxiVwiGf0WcJLDf1InrIw/Mv0Iz0z3HICVU//n
XAB0tWDuPAQytVMS3UC2TxlhUnD3mycAhS+6hvqNzBhWxtaGUaotR8IhtJPt0vnrgG3MwskUxfsv
e5AOhS0kzDjE2+japb2rtWU+Fb+3iuMinZoL1ZHZduN0UXYEpKdgbHbIyHtzYVOZ4/XS/QkhbnCM
P3IahdgfgYUbk8FrlKpKuvgi6X1AmxGHYkdYpAIzgoBNvFOVUeO6avE/vm+yg46IFbKLu18BxzNl
FqsipjZbuFt4x1eqi6UgD0nf3h57JHwJSygvcz3f6N7Wy29YpJ0vBRYlKQ6OgmSs20AAd4xUBObl
/BUG7SOWIP75pmAM4w76dQL85GFctZUWpIZP0vz4ehQnJdG7r2l9P9x4YENfMJkDbSfcNc8vJRRn
NpSGQfwsaTTCabUGteiI5cM4BndBNuNdj3S+yGoLbLvWR2TN3Yoh0oY8SsX9q8kFvJSnBgZXralS
eo+5LYjwmEUkMyqT45qRfdrSVB/euH1txCGA23Avn2EryuLs6clXfSaYDLn9QNwKSbTsS8qs3bei
CFsg3N/v6pX0LnwraI7mHSbdd59CqZDvFbceqv9DDxs+nvSd9lCAvqs+MZ5c09fMFdsOFYMORXLk
YTfvdyA1t5VjGYBr5wc5/58qMeoW/4gahuh4h6FNA+UwPd1IBB4UJ7s1iOh4EdzlQdDuERZNhh5J
AxKGQ19S2oWfmky6Im/r05z1sssoefCoYE7+ggx1iStS0tUg6r5rLYObbmLXcOxe3ygbBnaFxItb
xfPnoUIQQ3OjZi+QjMeeWuCNETJ7EOOgjAA3cOQLcr1v290UKSW2YLxGKDUAlGUXSWOssAcowsQV
P/p96zCVVsMxdOp1yE17zfzcNFtIk2OpUkBPXKHytdEx1Y6khkDg0iRYARjq4gjDU8cFa4mPdXb7
Kup61aY/JPFl9bPaR81J4h58GnfQiXJpS4WLgeVhxqT0z5WFP9N5XRBxe8Dzcl2D4CmpWFfWlK70
Mm3fi1KF2LpkqfnJsndv+tVV+ySCWSdPU1beA6RJgtPRlRxol/xOEbJ7dvs2E9G08HkD9Bm/PWEq
002ArRTsDI5PhQBZya4lMT7vrM+OeSUTZnMKjolQ+QEgJE6ozMh+1w5idyEG7GdT34GQ49Q40+GB
tofCc8MVXFehcwj03hBhtlA5+x8yKQ/usxpYhxykvmluwB6QdrMe/sHkQ7AbXi1q3bh3Aoof1YSm
TF/l6CYSN1afqddkAuNhem2F6D/wFzlZCyQbV7/Oo66BZGALly7uquL0I+c52VKXjbypgpitzAWC
kB1UtutxsTyV2tcOlmM/ET91+kZw/YCf2Y6L6oA89QtzW+PYVSCXbtTri6C4byJbahL0enyLv2wK
y2i9LSm4+Xf148ZT7jSeIZ4/9Sma2AbYmLqUMYLVz30xvgWAK3QdXKdmFnlg1ewU/ng6MQJdp5JW
BFOQP1IhPWLztwWcgq3oErga0h61iRuZWz7OusuRF3+93OJNcISMFHvBrNvyMArs7A/JfsdNsDaO
TCLZn22ZSzR72eyEPlDyCFVM5v4NEE7PKgIUm67iaAy8MFALrX16LGRsSc45DMAOoameHUR2Fo43
98hk/aQmn79x7ScFTsJHCjZjci8uN1IGbN9fcFfH3ZZtWcKZErAs39z13T0/XZ++MZcQPPdnBWRr
uGsh0skeRezriR504FsOvbBhVyNQYhYwzwrOzk7QBJUUidAY75UpmUOHNCEm+xhNx3p13/j1zH5a
8mrNtW86PuGai7/tgHRArYYkrhznjeKsZgvAS3mSecKZPuBEK1lbruCWrzWU4P8YAGlvw3CBlqj+
Bebn1sAIfVtplU1Tz8D5fCm6EOvBceSdigN33IV75dbWf3+jcpGvxKJ21u0fAxYYkUeax8PKJLzJ
AA3XafmnPK/dFkXRZ7+DlaMzjsyAq4jbirsyB1kdVHdCnrbXN1FmpGpAf+OO9sMNDFsQGpuPTjtR
js+/hdE2lLvG123NpTOgYq/FhApC2ToV/OBYAX9af4Z7Iin8QCrVNS9jLrZPuibl17N6smxW6naN
8KLmQ8pkJgxAC5IjZ8zHr79Hi5wf1NaVU5O47abDhRfIkss4T7dcxbip0m6J0ebZt4/pFD+LZBFu
hTO/3VHyPqEbggYSxP7wk7rafxauCGmtv3pOd5U8jycmgc+1LDNZLHFAmwnxhRXU6Xt/CvCJGETf
ssb/DYMfDCX5fpMkaO8RmdsZoRWfz63K0t035MFftIju1tXHeV50Vp8mfe6gTs44HfxXRTlx4eid
oPZtYaG4ZlrnQ8fDopJOt9nf5S0Ts555YB9qGL6/efvXT9xQd+KVU7pOghPjBaEJgeyj4gXf6nol
77hCuB5+8JIpOxcfjaxT8G0cPT1sEiIM/1b8rFbIt6lhx9VmKKBV5Idu3Bk6RfJsUp1vMqvN7ewM
zN+sldgXfB9jJr3+sGp9HbGnyDaHjSzvpXHqrdIWd2CXqDZkEdHPtfrQsrswjVj2dp8ekMVz/gBd
Kwo9v9j39a4JjSLTKvDuyC01VBlJqyzNERxey4ComsB509zghZ1npm++AFSbml1oHguZwoCHP14h
7ubY9ESO7xSFa+/7igQZhdS+cM/uMGm+FsoB6NVfpUJWSkk/DReOi+Uc1Nzea2FR/dUBN/cY30Ji
k35ViedxoF56kM9hyV9iBdgqIki+4nnvc5k69sn0q0Lxf7jlCm+OKFFMhBJRsTRvOuMe4FMCLsyz
XQPF503TQ4tVoBw2VKixbM3+mfkIQLQQLyvVHpic2tj5evvt63qqSKoR6Qgtu05UIB0xWC6YZJvp
OGoisTfIos0sYfuj62xrgmO6dqNt7a5wL4dy7cnYahWLUKo3Z0ZdVo+f+0OFztvHp0KR/MwypRVU
OjQXoa5FK3d6ss/fySn1ldAei5UJ8YNXXbHp5yEf6yHHdI8GFGppAJJdUms1nFKUz1lxygWax5Cq
UaiDsLu9nuSA8a1hWij7ELnbt593uyuPS7gu3L7MYqckT2hHH8lJi/sI5Gw7KQjPoLME6zm/j5qF
ndlo0AosaL5pJZLKPxMtrnhG/jm5DhCns9zkUj/5wTlDQ7KzVyGuIm1hRNzBERhKlJuWzBj4PJxJ
H68n+T5g+W4ZXQRHWAhXAF98fNP6OGQOTt41zZ1z7mj71B6hm9fHF5WWouvRWrX49kx0nN0rEmnJ
0Vjmd6u1woWwcpJ6m0z2DTQBsxNl1bTqCqSZrkHWPeB0t7Jcbu8NNRId/qqX5RfXrfDYoxEfQuAA
v4pQAm0GTrlg9pglo9jIImV7gRbmTocOe4CwfGCG2I/4OLRwhVhVXcyHkwy8yIJJ7OqOUn2Hkp7A
wujDD4hT1sNvtmsMPQnk6hmevVY+N1EX2QsckbGI9f15jqqZtvUQlqAa3H8GPFzNyB9Re0wQzlys
nUQOVHU0165Mt6LL+b+4XekeBtqDioEU7kc8h56GRIhSQuLDb1S5RrFSZQnoMmaKfuyk6jehT8eI
7h/utQHyfwE/8H/kGkPIkC3zVFiHYIUzkljo7mIMPg3AKDoo77uV30GnTDqjY8JfTmWA2wvRrj62
CNvwMO0jsrj/YGs+TU8QaFEDppG5aeiCP8xEXCz+qmaRP5Qo9yah/yCLuhfwI5cOpZA0daujf8Xn
dMsPBebBNyBLkcZd1Da/+y3KsePLOGU4VoL8GeM589bhgbtOnFs/OtO7MPaRO8146nFSuNXHEjEc
13nc9iJSeBpYlM57N3PSOBCTtpvmfDEx/M1GJ/DIlcCkM9JZ7w2TLuc2SAdBpI/7fRr77FX4Hr6A
ggFtX13OsYnc9MOFRhPGVgm5JO2c3TXf7fKM4T4cvzA7jQI9W1WCsljyv/pE1rOoCj4dNuSZxECP
A/8JWTk/2IZJM7laHmyta1nYtynD44DFOv4r2U7HedC06TInEaraeHxJHdcznI9PUA5enva4F8tl
+MInNQfUddV2/Vj0gqHuojOzzcf5GXmxMwy4aJ+0+IN9bEcbmgmfVznzGN5xyRIkBvmmRM3/qGd3
FhJ0KovAt/I4+gVa7o+GUGYolA3DQTRynMRRMA5gde4R2TZK0/KNzTj8IMNVOPKFP6xHsJqM7ZON
kFTzS0k0iMq+GYc58bXX52JNzih65w9qg8e2Ehd+P50lm2Fhc/lyB06RB2S6UMJtsY+fPiTz9Ur/
4T9fuFgOhJ183H353Hm94RIiQ1lZZRqZTb+akVHIOc1YN3OnVmCp0rKSzZHOWjzvwGmscbws7j0w
jlMNOLRFGU0kr/jAh2XX9MKiLzI8nuyCh2NTphvf68ONUVjQNT0d1geV7K3DQuek7z8Hm1po5kyW
Extz6VH4WmXSzggcGuaA86QP6wCVAYW3xNdJgq+oczXjalHoxh9vRwaUHWKuaU1Qe1BnNUlLQVzr
fMTVRRumE9AOo6E90tS55nOtbrFtnP2fZqeuQTV4HudkChjZBbRlym8fZyC38o0/8BBRrnhrjxUD
XUYIIjFaVRJjccoYxo0UsDahhVIS7kYSCZ02FPrq9idOVs5po6bqv535N2eujZsSZ+awyHNKKiKK
cqnIAdKD8kTGkZVvNQxQutx3soOKixQaVpODmlbgQgK6TqIES0Qnd+MCEMuNNeb/b983lQMJ/U/3
LwcYt9Lp1lZlNVsh1syaOcGXa5Db3UpBEg4qHVXXX24G02v7qMx7WLgldOZBb3bdQdU5NEb1bS7L
SC6ps9cOVrYsYZSXsVp09/RRvPbD9zh6NdNPYxomEg+cNhkKcc7cvu44jEYbrGARxs65CDR7Ky66
RSqaaRMjw5KT3JKoPlG+qKwzwQnDmxF8euRbIFndp9v1WahhCrGqlrZbimjUphOe9sCj7xk4NRU+
I2MQpb4DMEvPsalB5JBwaVENEpqh75xyfiKa9i1QhWMr2lFusn3LzApgMLAo70d3MPjxZ7NvC6W+
qXnqtWYf5KncOFP7P0mI/75Cbwl9PPS+zDloMCd1ruUGFP18kjFaUiPqkqJn/jVjF6TwrBF+vzhe
Tg/s/izpbaQ9w2XDxTJYK5BQ+eFfW58fqpdpHGsnuf1iZDYw2VcEvqY7t3r1JToqvVfH/4Q+yPf+
PNsVi6fX0VsxRukxCTOx6xs1b7yhoBj0GNIliVg9h53k6/Y1q/dBtw3cHsKmtFq2tIZ+NzR/z4ti
39cp35CiaxfFK/Z7yWwMsPHtQQcRfJ6KS20lvbqtKP9wfvGHYC7BbhT5LNnIRO/XmFb7BNis5l9/
bqmaCwUlsZLCZACsEccY0kQTqk/mwRS63wd1vw7l0pfYsOEfU2EekMTFasCpCkmJDZ4VVWqAhfv2
Vi1kXGGNdLl8FoWx0iAuLLnYDNHJ2beJo69Rlb847/YrG+c4X8zAsnG/tyDuAdSYz3OBjvQtWWg6
kKUcOx4U9nTx25LUxru+AqjjAsAfi4aCbQj1scezTYtTM0sj1F0JLAf9GJV5efVsKjBisUqR3TxT
RkKqqPdVB9ayqaTrlIPA6kZzuTdGNHI9487uEiVoxn7Mg0DFypm71BAcvPracFPpVCtjoFcRUfig
d1Zg6XM2/Lj4HKg9bh3IIKo15GD7e7HdT8zWnYhro0lhJA6x8PVG9giXiG5nGxergyA+XROs9P3j
yzfU9c7046fpLsg+B9bv0NBejL5uAjjeyxd4KANaAOQqmNneyaxgFSZz+pDkOLo69BgIJrRz1CTB
9ZQrAYgim/SSm0YjXxhXSP1v8xerC7mgholTvsSYAahwC1BysXlZg+G/iXCzAAsm8EjA0EFmz8s7
Emgdaqh3v8SSe4SROXHfaTl4VVLf6wK7oNiVpRxUXCI4I6vwILIaCk2znASrh+G+v2Li27XnF/HB
jw4MSxcUGPRty6gc5um3LAWs3zdw/JkBzlv9WUr15wqwmUG0j+uftLXov9Nu++nW6BTruyCce0zw
CQoBBDwiBB6WHullfUMrKsHqFm1yxa56H+VuypqNlTXlJe9QBuIikFHECQIa1h6Zkq3KwY3da57J
RPrxaBRMalAt81ImkZ1bI+LqhR2n9LKeI5wzR1NeyTY95yPGm4Ar8TItO35g/CvBigCtRUP6Xw2W
puSiQbCCn6AfhVBuJt3z1XSjUH4SXe4M1Rk6PSVGc16EHyOphtB4Wh/65VehZvHLxQKiIg7mQH1i
rEJMEOKvCiJxrgOQO3WI4DT11GOxA4TVUNagNdXnFPSBBjqE/r6ng0fLe1rlTeQxh9qCGgyg/mzf
wD2e3vaHLONGp1wGd2+sSrqzM/BIKIBYPl4YT/U0ANpFgtJZZfJBOVlv5Gf0nuFAdOS65Svj6FRr
zdisRTeVsqJ45n3jD9Uphl9yN0yRd2J/mivlciEcLo6VSJyE383N3Bs2secswIZ8WfE25pDQeU2F
EC25E0YtOpoHg+fJWJGC5xJ4l2rUL7umguVoWLtJeG2p/t1jTsEe6Jwp7G/8xr7tk83nfA/lmEdN
ReEiDeXr5d/XWTxO2KBTvvFIPe9bNd+RdzyuKKXTyCh9P6rDxm1Vlh66i8+T5MtKTzZiOI8jvDlt
45cLL+o6ewVh9dVr6CRSKhzSHTjbrscGE494hoGy1hUrXyLftNzjbItHhz1IE20/krPkrm4iE1Fy
VSFg+mNOn07vkbg5Onpb1rBkAiYs1a2o2uIM1iMMqPLwNAnISeTx5UCiMxyGC/EDsF4T9yw64wEr
LUuUbWKaEtTzCDA8kDnQzNCsZSoibPc78XX6A1STVuNafhxGpForvq9IdAag3ft/V7owtgQCxzM7
f/5k34AIezvOlE2jw+0P/F1rMcI/LU3CRmnW5JzW6HscIv1FCQCRS/OnbAsrM4X/UOfUNPECkmr7
w31ftl0Cw243tAN1Va0LEgKLrsPP3th/OF/G7Zrol7KJpIOdVNJX282htsaFcXyfVrUAVbkXs3cK
hvWnhwDDVMxlkrJ3NbI7GCQXD6BDWzgVhKoD3lWpNObDAko8bOYIe7NE35d/gXqWGLWj6ZW6IJyx
eT5SgskKVBccdaSY2/NLnDDmX8K5nAf9xrBEU6bp6Q/trBfjHYkO1idVmyT+dS+VU5m3DSLwBsOz
eS0coYLjb+L+jgSZu/xEjJ87Eq/roQjz05hp8DwHPV9uYERe6gQMAL8usWsGATd2PjIGE/iRecqn
QoMsizTQY6JpXHNkcz/a22sOGKBmx5OTGDsb8a2U0NlFsm5K3bCXL7hCBTCcoEsK4KHegCNcx5o2
WFONVwYraTVip1GoUDpJE6gQ8p3+C/mw+5krhrXEl2lg6fdXkntB/FEw8YsfJOCFQB6W0s4omo0B
bAeyFqeA+KJtw383MROJ8irIxbzyHdqe9mfmv9NkWFediuDwrogC0+v29JehnjoalhzhMDzg9ODe
Mdyln0/G8r+EYGySqUNuOHlVZsWbsUNYv84ZmNTQn4sy9eD+qDXYHYm3On4oWDByzp3UXkE9AbQN
ELB1G53qrJnSup4SGo0I7J4taFl0N3/XLA9JB1iO13RBICQMmiPndCQbpFSM1WCo4nSgHBmeCe+R
BLRTW5X7rybxrQy6PmfJU1KMTqhfk5sbBB4d7Pm41vNWI/vLZuZOj+g7moYJmwIwi+FiF+hAc2zA
AzNvGMYnwNaVcRTtcl5epRW40NuSH/xHcyZyOt11uBGMDI6J2YesQGJDrSbF6K5tkAf1aPHFHYur
Tuq10Mqv6ZoCUdGrNxnq6oNO/vunW4L9a1bGzx3/nYwVG1PD0TmBYkVRE/LRr4yCkvkeVYKtyNke
GNZNiZtBUemLWeNq9jbUTrNB6wrXdjb7sgmBf5UiwnsLEf3hnFjCMl3WxqJTzubvnv9jWHQuSHCM
h4ugFLFgmGY3jJGUvytJW6c1euSw1vhjdCBfBbdn/yUHX/Qe00Uxb2jn+XuIXHzAYNKXQwSrI/qG
sVVc2a5usZ//wrmuNpN3NhOKAQl3p6sFCkV22lKVthA/A+lNqxvhHHCwL4de2cLuDewir1aRE0Ae
Ycy9kxkLBqwEsCYN2a6ocwtdZ4i82sHdMNlumJvahyOzS3jeN3gt4SozoFWsgoWpWyfpW5IsPtRD
QMdtTvVxQ33d2tBjNfaVP1sMh2e0p6Nra6vGO79p/9mZ1X+twS+nD9i3t2FmSEWb8/mi1ISrJapJ
tI1fHoe5E1l0wGvZ11vQPp85QMXRc3vz0Y49f98Q6La++W6c7j7xiFFb4lc6X8/qw1MchkKaxsPG
yxEDvUO7X+ARqzqvjl7P/uDrnxyt1KFfl3ChtApj8IBOOqI/HYOzXL4v0UThSgtCEd0y/E3eoEVr
rILAXzSPo9S0Ct2N6ogGCFOPvUYDC+0fajGcsznKT5Go6t6RqxDfRJOinP88q58aRaaW9jV8iqip
JxgSOyT58zA6TtFmVOlgiiL0MLTiPMMQApdqcNfNIMuJNaIo+pQm40GvrLOlrSvkbN7CpNX8hclw
FV6hcQH0knXpQczz+hUBuaMZYi67mTEEkdoOU51oMZqJoUvY6Xob7pSEFEozAZZuEJ4q0mu51fpC
cqcGYsLsSyRux/AOUVAO42wKzdZq0R5O0IEwULnEfpp15+PTv/T7VrWAkI2eyUoM7dffuqXmhsCk
wk+tF7/+3b5kZ8hjmEUNuuB2df/81+QVNYKOpPSXiU/XvOZu/y3rjJA9wtOIhuNrNBt6rW8oEdJ0
kaqCF+bQ3NfZ3csSrH08FQwbcT7UIqmoEA8pkQE0jEVzgd8Cbt3Feu9+KEA5zDVu0UGg0nPGu6UI
+Sm6dUU45lJYlXXlxqAIY0+F6kdZ6v/THVdNPcpzYwe3nLgskau6vGImbc/GKgew0fBTf3U4sBKS
tZzVTExqS/pqWR/RfZpO4zx1kKaXiD0rk5ElZlM9fViKvrp5Xf0evaYvQq/vKM7sW11GWmunLCHO
cGcwUWbuZfYzhTPiSu7yLz2YjVpd376j+VfDZkTyF5HBiLQAxgiD47VKfJHizIe24spY4bjCFyHh
bJqm+98z1LKDRKX9Tdftw5apiF3BOMRKZfoYoayF8o0LRNcIF0SZ2D+D+2Lvx4rZPZJdj6vbu2GG
GPOInBfrwAGfv4XCfgvxk9APTMikPrtCKAY/Mt7xCZEJfLAmJo1rSusPTA5WH48sqC4EnvFYrK37
FCLj4uhgvN7Km6BMiBrtQ+GGhZw5GQWRnwjUneaprJDuE3S2makfPjHuDd+CYgW/ljEWmEFoQVZo
3yNoTbj1YV0GZPWbbRvD29IrnWaqF26phv+obHNVVr779YWdLjJpiKr1PUz0BaNYjqx59Iaj/X32
Jx4P2c8Jq1w208ihv+DmUl/Ir5rwPhAFd5mKnsvAJ383kQy25UQT6c0DZo2r0EKTBXenwDSzUjSu
AHqzuGEXq9p8Uuzg9s7ptwT4unwkbvNbtmPsuRd2yxXAjI7OnyNW3X9AMsrYmfilA7kbh/OZHC1E
poZIK9UuU/PUGCSnsM4z4JkvDGe6qwRZMRN6iqSY04IxPG3Yn6Oie2nCUsAeicAsN2wAYIFRLSMA
1qlalzefyCKsjoHw/rk9JuO0byesNNtA3zQ+kumZquySKzViiRgfl8cesEcX1X4wv6XygbQBp5gf
5qs2Uwa4IIDlPrNvH/EMmI7HMafnN17ZiLUVdBpPNFWLbRgDDAHFUjFIKt42asQNESoYTwR1hawg
5MsyRKAyzJ8uwJhh2Rk5JTgl4fZ3kmWNkP0c7VriQ55LLGdcLRhOLHE9VFPa6vQKa0FHfGfJ8nxe
9o58J8FLyaOOfmtGFRcWUqd8LFD08W3wFEPY0qK5BQZMLuXROfavWubm5T23ZlVZWDzKiEmP/J85
W1DxPE522jKwz/OUiaqHVfD8t6ZbU0pF8Tz4Yt6fHFJjwbPwC1fYL1SgN2vrwkzGJq6aVNlbjw69
MMsKVBp05LhKT1TJD0d+c7c9aZ26l04NjQaL5d0hya8WQKeBP/n363IlyBP1kLAtx7NryyVXSv0m
ISJF8jamN8J+ecZ7tmfx0wwZDDHn1KvByEXsMUUijS3j59pWMF95B2nUfNIqpJJ59Voozu0gTwkL
cQXhy65UUFW5QO7C5iW0utLJ5wS1ztIzwNQIxUcVsd04ZgH4rFtvwQoa2yx5pRjZbgzNskRn3iZF
RzECSNwcVicptiNDIbN1yci+JkfjshkKwaQx79B7nFBoq5N9Ru+ZWtGxrNI/yaLP98zAjuRR7BCu
uZqIfZl2DXIpHBQeRnsYPJuZQ7NooreHp5iVtE1Vn7cDPadjKVGPOPxExOcQygJVZ8TQ86uKYLBI
ZpLgxdHzHDXeJ0FMErPSqiJhkiy3nASbSglG1iWXis+kNRY3nE/ekEgVXhD2s03BHV4i9g5T7a2T
ifMw6ASnJUO/rlXMkEwvu5eGz+qmMcUL6P3Vqv6zE1pVcDE3eEYATWC4yrGAimL5vsZMvUM1h7hv
NX4khsTcfJiZGZuzBJzjvo3PeTKgErisrajCuUFJSI5OAGkcAb0fR6Gl80yWpG47p8Q+F/99iwK1
DrKV1/dhPVi6tmYUQe7hCX5Nh5xQK9HbukjoRpSQF5NeOoCPCZK7rQuVlPL4/dZAotG/g/gW4a7+
NKpY4vh4MgKxpvjxGnEEeV3rWuHTaCM/I1DbggGd1diMO0PeF2fz34+maJpdbc3/FAXOZAWTpYVr
9BMLv9CSvb7ULOoj2jCQJn10+FCzVs72a7GYxz/rzFOEcvDWrRyTI3Osxsv778tYSO4/g8KZJKpb
N7o0bLU3rU5389EiFSkup4mzbnj113DELpXcleUvGnqjEBzZKv6ZVfEe/97IPmqHvy7o9TIwnxTR
bfaBLPpZDWVlyjEz5wl5ZSV862N/0ZWr8BgWk0oo6U9ds89s6nB+WAzylRWXDTuMuTPNP9MVxgRB
m55kXktPiluYT//oVKYKyXe3JID/1WaVnFJ94iEQgp0d+DB1R+vagsLuV/hp0hB7S1kO0LYAW726
ECiO7WOSm7//uiJ6dsixRbpNmA7HKp+rhAM0xfsGOIoj4F1gJH2ORqqYcv/yVR64NhGeg7n2rZ7o
VwIAc793aA13BDzrSClKEHWixJhCKZZHIiJn7yHTjEU4MGknmxHSQ3XoNGuvm8ZpxDOSaqRftOxE
KyTEKE35dYtdwPx8rzuXFHsY2q4mX8c6ktaZeqbpv/1n4/ek/e5MR0uqCNEtED6TMxHvTvjRArUu
c3QB2ttk90XQpRjeLoOCFMo0ge4/ogHDpboe25vTTqRjHDf6MdmODdWed4asfCI5a8uXJhCcUu1i
1t9kLoD02ljkB/0OIXFA0gIOVFQIh84lVq44KRq3rEtznPqdntmCVYcmrdiD7NfWmznGMhDCSz7I
vTzozqCUPEBcDidYdJ9QCpZJSePQNdcEw6INfplNykooR1z2kx5oqYJD7dQXGjuktk3oOxHWsYOV
ISftCauqTveSmCxI8Qq4KTQgZkLswzSE/4kHpST5Qwe94HFwlK4mI4Gmh+oEMd5ygya7QNfyc5jC
NkME+U7zQHEa8SvBLwJXml809YzuOXgDMy7pp2ZySqPqJ5rzxOrzAF50mAEvbdzoq29ZNf3U/ea5
MrmhvCjJIh1M958cd8h5hTJdwO9gpSyJKffcJ7YF8PUo4ynY3wfCCg3Rv5Bf14DQq/i+NAuDYM2V
1aaH7LgPqaxenpd3FQkuIw6REXVlnaCnRBGZToWRFUW2PMbG6sF59pY41ywyi7iWzpq5FEbvyTxu
MYRL2yG9xqKZSlKCKG5b2fBGA0oV3TjtZEaEVuFj8G+8vP/nam6quAr2gG0lZ2CAv5XC2o0j2b1v
gHaM9o7Nc4qOH5Gn/qduFhRNtBmuF2rF/Gpj1zfJDOWEmY6Cl3LAdbiq+MiYCpHNam9DVBrFhXtc
S/pHov52WQYPGjMHem8CQGSpqT3XpKZTuG7d+aJONgw8GdInEgV1qNLPCHCxM1728rzrr8rhMxR4
TXZS3HgYsvscDDk6CMClA9dMggaiQ04zFPv9oigvi8RmBuwhUBJq3SLtt6c9i2Yuc3DI9wHtswr5
rXMSe9dyy+A72tQSw4SlkISnD4PyR4X5LJAnvRj4KOKVeFRtuzbzyIL6ChqG2z4aTOj7KL/+qWUS
tVX3htwrThx2EiDEMdx/vCNjQejh+tVXP+B2WpL4yQwkfqe28wLwxdoiobsYmi43imdDN/4rte4g
J6amWWEG1iuUIc68FmeidVzP2gjl9FJ5qhyfZny1R6SPzHC/5pLj55ilfZnr6jVtNb48A7MrLam2
YiRwy4C6CpAYi1fdmtrr9HO0WoepUpyLm1g10K1k06zKYUnuhOdOmvbamXlaXtEh9KHjNh45ILsN
BNFGtk4/LsqXAxOat+WvTMZT3xDcNfL3MPZU8MxyGh+Yh1Jz4BCSD4q99IrfEZbgTy/mOq9SIXN2
DW4gke08YHwagPfQ57LNnYK7lSUFRhN/UeoXQV4BDJOLxpxpmuRufHeFwGRUIIkFpCh7Jf+4KKQq
PT3HlxDqf9HJ3K9IHeCAlKOfS9OwVqZDvfJnw/bcMLTxO5O9+NIYm8ImIC5b55YN5qGiAJOh0WdD
TkxbjMVRHlirdsylX2x8Jv7sBzvIvIo1kKgnGK/6fQlUxgMBQ4QC/16C9iwgupuV/tiqyQnfkNur
qXwo1GriYPLjmRnXDTViDvdAQr4IFFmIkoKA3pA06xrlJlXwJIEOJUiZdqbXaPU+kXEsKxJ6UL79
zuimym6XRiOTW4V7wTePOce2Zuo7jnCDXVDfZDswG9cOFeotTzLqUavMOAtIn0Nu7DqJESYVFNlB
JTmjDoL1o8GXeQoqY6WfzTPZgzwCLfgtyVWcmiOsycTMmvI0QXx/lFBoH68k55Gc/XWBqTxJR8xV
nInDjE5S6SBHRSD/jLRfVTwDu37ZmvjBf+CEE2tl7DxxkbEBQRAJVJ3Cqvt73TpxNbLP+2o0X8rj
V4oIObJTdh4+lwcYC2TG9xazeU6yv4bHl7JcT6fSzLCMDckqtcrFyahv9TuphbE8rh7lymV0PKMV
R5ojDsZd7rNHI7cOntBeFaZWCRffog94NJa6QKiG49WOrfZS7OJy56pXKgZJF7juZ9G8Ptui3VWG
Vp2Lx3qpSw3gvFOMmfRF18EwNlU7XaDYdgMGNhKFekr7A8gJG4bUQL6T8wjKihmJqvDFpmeeJgRi
olI+h8Cwr7GtGvI2UBk0x/JsB2zl+ec+xlwicvoRlBrqsLmAVvA6uy6Sobu8tIA6sRZiof8XQ/v4
ypsUyiLxLjeGkNG++pXaQLrS/kEiakpQ4TuXQr+Z15Kb+/skqnrgzfGL9FSbmb7RZGr9U7329drM
05V5WQfp1rQrbgpCUVzjLBehHQZU1y+XERSSS5Bn4wOihwdf3fiEtamujd+eRoQnk9FwWRnee9wd
ER9Vp29dKBzSsXmZsXgCgLHKnMhZAOKr9obsmZUG3nn34UDI2TInOrmcVd/0XPheqYp+cu8zodhF
zX6uL1MrCxSYZtaKX7HDlyIjOXZVhM0qNV1E/r6A+z5iWeARTzgOehQCtJ2el3clusfPXRw7Ltle
ScbN7i+wSNmMd1YtVeLMgZ5T39I5g6CxhagXSSCYDkeqTZhtiynsdWWCUcov4m/3r76osU1uu2RC
MJUrewHYrdRlpHbU2tMgjzqhiBYeCkP+zWgPilua2pdyRAy9YsWvXwqNX9ICISMBkml+/rWgC0Ku
fNqBihY1M3RGfUu4el09XPC+NPEKPnWeXQrILjwfFeLqhVt0jYSiSPX6i6+sI/WiEs8tuU0rmFgk
T3mTEvVfbWPxa5A+li9Uo/tBxbKcRSrnE+UcvL/wjYyTltjdLWLHavwhOW1Ml9euaojoE7eg4+Dw
va0cYjNvqgrje2pxet6klKw0oqmR6FFgQ/BdorP34zhZT3KrcxInPHVYH9O2YzZd3q18w4S0fXvp
/mWNMEHTtKyaKzb6QDgtNJsqE+ebMxf00cQPPrboOsnKOZzlShJRoB7fZM6booO7yHfwa4PQXn2A
sfd/8v8jEvwiiQjAE4d+HTkklmyW+2+THzINAk33EjBa5ha11bq4azFf5pF2n31hXQw0U+m+d+dv
EAUBYY5SoaNvO9NLVLk1tQ6oFDx4iwu3H3AlpMwkbSuRAGoVBQD/j33vrxK9V2BFdokYV5fbOSRF
CbKxd3Oz8H4fQV+6wvkPNfPV+aM+ULb/R9Oc347TsNuF98p3ywt5yhd0asUo35ye3BqE3R0XoygB
aL4NPrKVAK+lP6nkGXFt8kccW5KeQxfgAixYtCGMrE5TjgHYCrTGtIEYW9IUXzs20DbZiVMSgBnb
1Owgc0D/R0U56EFFBaljHdygxxo+0NYO1kVsTJLljGTRBM48Nwa7ypzbmASocvp0LLfEttAclpV2
ctbeApDDk9O41cm6L9/97LFJSn1Ie6bYRSDzQznDyh0QDv5Esh0PVfeaXQHkwotRWXfGggql1kSR
yxDa36gw8L0mZG7ulvYlvbxXCs9XDBtOXjqGM2ffglE3N5ewwrlXwYD2OZzuKV+zflcpFBtHQK/1
1TFJuOOM+lP9XaYBTwtecYxqt+D/u8KN9MbCKfaVzeBip8h0KFRcM5sw+XigZ5VOQl6HbHUbqKxf
NRp5bKq5DU37cyYVXkJpPte47ZOoRGZWTN66fkudme+HHrcPQCJLS4e9CdT8s1QSPVshIqC2OxDY
rKmCv6IJo5DclIuoTW66XZDVf8vLQQTa/B6YpmX2DJTic1q8X5BsDl5A66KLiEcPVy7dId00nDTt
/LoDxEXJdbhV1uxSbpuQJrprknbN9D3hXwtkmcBZ4ghgQrHfRAUmGfhB2NPMyXGOuHQp2fpvF0ih
t3Mziz9x2aPJBDuJw+U9GO7RBZZR9GDrfEoUeVMjK/zCFfbZKFO4Dwcb9I8c3HLGFfRN/n2PFEJN
lV7VoxfP08szVqkS7StWX9gn0WLN1nVTx29VPkZXDPBTbfV20hE/qEWoXsD88I5ucCq3mSI7e9yC
B9NoPPiAAgDVR8hJkABDCuGoGf2O6dG3m51lWmLL/rZpkIhQrJZP1K3KsopQEfc45Vn9Q8K6cIb3
MA7WcMR76I6CLV0wihF4AdFWkkt8ktud1aPZbhToTmqlvObyJGQoMGg7yiDCfb9iWWYgLCCHLI4k
01dbqh3JXtwEi4j2asTFckULRJJhym6VZLV2UR3WUNmUCic+vmBaOXLNUDAE0jYsjV6+wy6b7/pV
bcpwKJy94GnrHlkNVznoaTiok/zzx+IMfaD+Z6a/4l6pPVFGxUGmYQfqidvLHkJ781SoPBXTCXD/
nri6SU4+WTnejK8uqa+41q3fs9Qq1Lezg9CgUqjcGLSEEEDRl61wJlHBunlTFGGwIEDM4A7vq7HX
AqimCzsBURqdpU4IZvKEBGwy6T9K6BOVuEo16iBDAXb6QwC11+JaoIbXFT4VATApb28K9rFsGpZ8
m5HI12hatFdIR2gD+yVuDbac6FGFsL5nvwNz9vub/9+WW+vLdCOKq6M2pGjyTHKu2Vo/4mrC20tO
tFeoG9QlNKk+2nX0UYT6K2KwOBPwIq8eVcDrJ6VW4X40ZHo5tD2np8JLhFxVYx8caB/vDiCS1thc
QoUG9RVD0ggAMZA4xLBXrIFL3eDzJpzdbhhod7xrKs+rVbRnPXTuxzrNBC7F7K0rFbR2rDlW0FbE
JHOtwPp/O7lp2SiblXRSwU3TD00YDE5CZdJV37+Oae44gNgJ88g9bay/wAOK2FJgBJ7AHiFhaxOb
Ugs1Rpwqu1byHMucgp7FiKdAdAyA+0LgW8JbqlB5IuwyQsOke6zWBH1CgGPWrcyYEtBV4OWq4zQ3
Z/IXqs8tSvbvu42kqaJA1Qb4RLNm/Hd6wNdmcauwM+vjmru+k+wh0/5EHm5Si8ArVSXhvmuJV7/d
SFdCsSxIuMGIz2BQje622vnRzquqGaJMgTNu4lJg/thv2/5e8bhIDRTh+KgbMt27jLseBpjBYJIO
ZKD1JIxKY+JxSsFrUvJ9lU749qLwzSdpJs9i2YRTn3fc2ZFu5cuBQN4q9089qDanvMneYYfZpd0S
R0VIfthLcJd2rco1j3z0zPCbSEv/QIB5cIo6/Gn4o/K9+O0/2DyzL7SANyWwTW/riVmiFxV61KkA
ptYNLjmFAOWCqEaNQO9OrBiLBK2Fp6Ba2mPfdbVLVVjbsH44u7WzY/lrKiwy/5/7j9y1XjT3F047
NJ18sSxYE42+a8ZXRxPUZvTBTrIVV8kKHkWna5egEXGrUjINdRyPKvoz+l6nkqcY+F357Ci6UHxu
gsUW55PZ71HT8WZGJRSdXac+y5VVkBYh7QmjlNqkDQ6C0j1w1AAsL3rDngFCoETata6Grve6IQ1i
vV+B+xya0Njg6WaTfdvfHMAWdagj4umPaHMSiw6oOHrPWiORZ/SrMuRCqrdGFpb37r/U8xMZ5cPO
KzWsT1pj/PzyJc7He5ToV31yIOFtnNfKhz0pp+ur5+oxGuNWAW+JG920o0Er/++rnb6yeXVkdCC9
2rGHbJAjuHhusLzOYZZWONtjCXsQ5Vp6RUfnNoPW1Io7A5q9ix6LtR8XcQCXSnQu1yPTq9TWFyJM
PPK8TXjz7Tvrz6nzKHSlFu0zl2tckIiIECgtpiX5H4M70fONNKd+n/kHZBXt3hmPS5cp4K0PrecZ
Kq888Dlsb06GN2TaTWIJg3B7qzQWkzQ4VFJFOOxYbnfXJPkKLur4VCiPZwLfETZj+hzaTduKg0Zc
hvP0aou785sq44Vx3i86EjYAu6KZodrEEYSU9Ezr2XO6a56+APESCITOQA45h79JW0euG30hcTSy
8yYfp2EJCyu2DBMXdBVr95d3A022IoG0ETpTuV3cj/bmTd71F8InVKYgYjD54U4HlPvCawk+jLM6
UTT4Ua1T17bCcw2rs9VKewYjv9B72xeE6dfgdHwKHTBrpJIcptx2vZDu+eAxrgyNYlqWQ2IGuYvZ
av2tRGj+/E9v7Ujl+eiu0CfbGZixrCuyA4Nw9fjIZDnRMfu8Z9YQ3wSIXdNQga78AWa0V1jXVGym
LhnHXVkEbLS6oMUI+iGkRLZXMc17mr+EeeupVqT2zfwLMm24oXxmYZtDaco115he3jvcNWTLdW6Y
hYKpUQp04EQ0RhEDCc33naRef7S3CREzKXwlpj1wCOGgk1WJCQHgtLZLVVP0gPQEGL+DVE+9k21N
nxKnMklOgifr4B35jLV3BK/GSNsVZIhSX5kcNZDs2koNg6NthQRDpTfYEZjbG2Ikiq1sIfKJkFy2
zoUVHANcKWMB6CxqKNpdM3S/i6adlmtBln/YcCqMP1w6cqK4dWELkXWuXHjwtYQSip3I5FVnNcA+
0NDfQm7lp2V3vI0+pU0+l9dTa+TBjsLiUy8kTZ20H68POz0o3siQOpvwrbrC32Tso8R0oVVbc2tn
NmvSL9Y+dWQz3uQwTQzfo0bdD1qx+Z+GN3f2oKrQAH0J8WcfGmrgLe7CJiMh6mHofgSRANG1eezH
arkUUdvxTjI4al6PFZH/F3VcpPrE6T9Kgo3hOxx4dciMWx8toX+zQX4dsIvrEV7gjhFkZExteNCx
JMdckrYDbCCRAVC5hXplD59NkD21Zoqokgh7gpsLLBgMW4RRg96XtpN/ISkmiEdZYB0IiOamCFI4
Hx10UIS3aa4VELzw6LVdcAcHdZlbUww9cF34eZrOG/wMtIYJSSKYK++BpMRfzYbMW8R4p+FEWEmn
2cWT0ouD3/ItfIvxV2h0BPiXFKI9+vjU+a0UjRm5OvqvmvBIZD/rpW0ruS9j8jlCarcWyZp7eInu
8aPhCoZBnCQUE+U4h1K3gMFACmavYqpPkEEwIPyjAKBYL9cZY/qgX0IKfLAItsiA8D/6lF5oec+R
x5EIdKk1GSXYbi/batMzf+r+lU5NEM2i9eJo2Eb2z78BXV7j49ip6MN1I6Yi0+KbRY6gt2l+OCLu
I5Do5eGtydSKxTyYMaW3mGzmf8znJ3O0OeUVvMXJyaoyyK0hGP5K1C/+MsFUTubAzUbhjyKVWgXN
y4gtkrNbF113x8DD/6MV1K4p7gyV1rOCt2W0qRblTGgrlw8HK8s7oBN9B/D/N4bsEkPSP/7m948w
11nXZGkftHuM7vX1D3XxA2Mv/tquCKWyMK3pGtNPAk7GRN4yjZbj0Bzddmp1XVw41E7WI82NvnWb
HD0nR8p85/6nJOcUj2ktBNJRKidNUJA21PtomWQkRslPE/JBeJlqy3cVoy7ITaoGs+quk5AS9VRf
fskmlyDx+gsJPJuTrxD0UimdP8jIXs7ckTHmPYIdRZzrb/rgk4cYHMTDKs/EAqZLOXH5H/e6/RVs
L03HBrqy8CEFkuMrwlMH81gvrIDzQmnhPtvPedj/WI5UygpxABxkEJCMOYfVXSU+NctlJIHnJZz5
qqU4O38UKl2TpPNJpMPseEU5ZHJ1aBO6/2jrvkGQUlUGtiWqQakEHN/b8GHHFOGAbK4q+ZupObx3
VAmLWIttZnP2++Q8uxzlfndFZH4xKk7o4cvH+Rq4l8jxxSbmKPRQfQqkceliZvrYKFfpBpZiGWqm
gcyMMrYCE6DCDXYO7gXwIwdDvHgC74C1lC8Zr1LQz22tAUZ77MfQ9xO/q2dPq89oOgfndXpa67Hj
Fc2HD7QVEyJbDYhAMMPsp/aPJ/ttGd8k2aLAE6gMz+sTST+FED96fhYqU+HESb11hXnJiYmnOqOE
Z1TdZRslkIIVyAp49xV0Wd+sTudyO5iohy0DmlGeiWOekD2kD8/SkKIg+2dIkP0PFMwuDs1uKVPt
OyqmN1q0/SobkkbUfa/YjsrdlSJPg1TNZLSdxJq4+vkJmkJorSRfuQ5wp8eXkQ6W/m5NCqu8vdrN
Zq8ZlDnAKFqmtXJIScxCysN3+N1cGKD3rPIRVJO4sO6qfPUSXOwMjO70Yc2yc/TIOY+dcukSogIY
ZlRyCIqm7IdtdDPWNcv2I6jxQGZUWwsK+iOTsk8uutg9qEC7M4YQ9Z6oBxvbAzaz71zGEwkLGoz8
Lh7biSspIG8MCX64QO8ndBv/hvWa8u8VIajWhyRR1nFG5n6GFRC1WVqqyWrpCX0OW9q9B629ug75
6lsWk2RtpfMhRWJzLP3obV/nZ9bFpnFlv8FHMfn1e9pBCyAM7g8NDdF9P0/+mfJanopuq3qG/cn2
qINf3+aSx59+mEH9MR+pRbfjYIcDMwJgLqkaaTxZ+KOD867S4FVbD1zEFGqtpzeuD8AWEcX6t4n3
ngnV9UzhbXsupO7yQp9YeE8MQuYB20xEwtWI42wASdL8Is4/ZZ9ts4vfGx1uEioQIKaaVnl3YvxH
oCmWGext9wNmIObQuMVhKpj4NoiWMnynmLpXgauqYxHA18tqwGQ5Dwg9X7XtqssgSLZOi8JDeznR
gQCPaG/6s2XBkIymiJQ1OnkZiE4ooejad/Krw/N5+XvA/tWtkSfEs/gvayUROvcR5iA3Qhw2k8A2
pYTzfqmYhHrpfuj769Zkl3Az6MgvX6eJOSgSstsekxNCgLMp+PP0ZwzPDt+PZCxylhLyffDLxbYk
OLaKfydjwHxuOJDEi+ug5TAEMq9OxQil6c/EjJ7di6GaauG8YntNSiRSh7kCuN8wCWwfJR9KCsyM
z8E2VRoHx2zVYFDdOinSOX2M7bbljLxOSIZU5rJGHFwMWdXM78NwS9hluRMy0q0iI3wmOl0QXRg6
/yzztvxE1L4QCJnZin2qKKAo703gftasYrte65/YALhsyXRzUbxn026YMs7FlPW54xIvFX+C7nGj
jfNxbK50n3UL/rwHGaaektlM/tKECYifzgKH88e5FEsrFYd2Nzw4tLpn6k38sv4fUrGzWg7nqo2N
CMzC3SY+bYdXEPA4PxYoJGXipIM578u2+zDKqfsgCpCol0eQznk3qfBgPQO/WNm0JhAXzC4Gdwbq
ZcM4SDFl5TGmQ9clmrnlQNaCwJffOgG+v6FuKauPWPGClretGAq8wqoLOw/33qtH6SM6dGoZ7pvU
jJL6zIjzOzDXWSLT0OQT6kWCzVvIVRTHG7lwvIAdgglnypUizPrVo/A6LUNAguzv6S4pL90r/E0l
CawtKtIRYXIJmhBIJeqSuiGAhLtBNUviJr0ZsyWiKQFMix6po0594Nc3vRjmi0NzsOdPHfV+F2/n
WnWr8oQwRhqIYFj9LPvlNpN6l+1nTGzd7W3NDi8jIjPbCEZdsDc4DrNruLmg7yl9X2qMPAyDI5JM
g7n5SCmVf2fQB1MwWt4QTW0iVkjNgxK3qfSINdk5F/0m8YH08k6MTiLh4ZEvavW1B/3N49vAaIA0
5+JW1l3gZFKVm56CVXP5hDyPcZhsSoSg5/GOltR4JNM3vYpNQlixZBJNj1ubpFg5oknRx4mlBaS7
Xwesh7RwjDjLs/JLJZKgzT+vFqMok/zSsFPGqxhoFx4McvfnloRacdv8KqjzVe6qXVq0qYeuHjfY
0FZfBytLwsswpPDiX5Aaaanr99PqGhDAF3SSIV3JFLFkAq4/QKjQigvzIpDKyZ0Y/oV6tdSsjP7T
Lly08xU9gy39W6A/zZTbdcg6wGuByROBGhnIwo0hemJqzp7TffCdgqro3Sp81fbTZ/vnzSXRRNtc
7oLT2IUQm2cXguLsPlFuDbKdrbU+zG5TD3w6l8J8ml4kGTQm+6/q6uVAuT9Z0Dfzm1VqFEkRS/Zn
fN1vaz4ueXom/e3g49112ELKXLz7IHZT+1I2t2dpkZahgRylJmVDqrrw/3k9t2ScpOCkqo/S+dFH
LHOh4n0FZlsS2WegrjndTpWDSr6/U9AquruLsWxhPPNDdGqlxOR8QmTzAOztA8CX98kuL2PBbXHw
MOfTGtA62Ws4gCsz85kaK5w7R+7yyBy4x32dMtKBSwB/B0iXfjaUgK3Wv+kuw804Ig/tdcbi7V73
nKsSN0mqaCFO8nw+d5kcEHvcXRBhEvU91u9TWVZO/9OCC8bG2mr31YZggeHzPjbBzBTmAgupTiQF
G1ulpXI8Oj5gImLI14rIWxhKuMU1DVZHXy6fT3VcemN+YUyVGPAfGbbfi3mmZwj7U6W4mF8wKZ3x
cZ8/pS+39cHbTQnoP4WOCRC63XMsblMiOqasF3w6hkmE2Kd9xz7vTFLKNQtSJjb+PfivedhliC1d
1FhELWCAR/97NBb+j3iwz0EE09MCf88UCIzTPzHs/HF+HahDWKc++r1oniQm5mSWoapuDjIun1fG
PFQU4Gy2H3lvE8pKtOleRooX5orark7ia5LCCn7EgxnhHk9r5eerslNskEC5fAQfSQ5KawzyqCcF
+E1IKRTJBFncthCz9Coi9W+lXGqfH4fG3VVmw0UHr5mj+CwiWS1/2hlmMP7BLqo0oyGgLwNdaLQc
w+MaLN0ixj6AiFR2bQguJLDbbtJZuy1vgNaSYT+ezPKA4/+rJmTO0OCRjelmHeDGrPPLcUNqd7QH
zT0B8/w5MnPlcqXtp2PU/MGycWRko2jFyjh/tjMA3BJFHhylaCHasaU5RN/y/8OW/VZ9VRebGSzv
gbZqojo2M9DSAWUlaIdmsDv7Lf28hQMvKVS70WNnFwptCw8AKqbLg+Xd4oWSs6o8GxoFxJBnetIY
TZ2ZKHv2zrAJLUJ6qZ7pbQ5oNuhR+nNvp6Yk2AXTpb5cxYHBFecUV2EhvondQ6hFLpHGcpAkW85y
W8aG69UwVOeKZlBe448gZGuP6jgz7BclqTaR+b/Q3lFMWXo01FXrdtLI+sJq+pOfNyAVc87IFhkZ
/Eg/f/VaAJ3AD1C9ATQO59FXk5ICaL4OCEkzZ57VsZmCYu4d+Vs4gKR6X3dUvW8RNVM0QVxLMzOa
WuCskTVwZScZfJm81Y6tjpeexJWT2BsFN1sArCPcd+4TTxwFaV9nz15T1NXIi7WC3X9XaBq5Fg1Z
kVnAlRW1F2Pbw7v8vo3g3G0sxeNfYvC/HmTQqlGpWVhq5teKN+c3cF3xQlt7RHG4JZSjmA5HgnmK
JSynR8f5xKurhTiwlGd4e7uyjm9ozGGSw8xZsdO6LXV7OurL+nDLQV1DMWBJ2/wBKCVv8tw41aUg
7KRdijM07+78Y2tutyEb+wk60Y+h3RPQmhaePmOwruZCWtu/Oyqg0XFfPV8mkhj+hU6otLjmp7QE
8fr/QTI+KF0rhvcWpzFgfF88e/3sIZhTZFYIa6SMOv05XenlAMIdN2IN8C8HcAUh0ryXpHl+mJ6H
p/e++8dzZ/G16yKw/IJASY7ys71ihOU+7uB1KPaLxCKcXVCkMFxDnCRj544mVbVikMvia+rqQkdG
PZ6ArXm213wkgBoWvFB2UO0CM7qjVa5w21AdhViiMjbNyEY6ZkPvYuxKhcKQwR5Gtr6SDZ3QSA6C
jcvnWR/fMav4/jyvaYFmy58V8OI5YhaH9h5AVZWANfnbFlp/wGd2h8FiyP2H9s3xMCGkEYWnGUWa
MzghxCg20x4QbEJLN3Ao836lIKvvGVwn5MO0ZOhMti0jF0nfA8enZma8qmByARTMRzVXbR0n2sn8
Msl7MZZOcAdnSeDQHjgK0+0wadA/00ZrRwXeJYlVxbNyRQzvT1vV15ZlY1PWNNqKiHCTPisDa4bU
sKI0kzJTN8NFzxqusfbmhhYnXU+fs52E8D/t9NAQnzE1wyxLn3L7pi3Vz4SGBlLeYWQgKTb2bA6/
9ZvNHN2ZkOBH7y67QpXxd7CUpe8yteugYTMLHDNM0rQTfK20QlLMsz1sL7kvY5fp+au9arDpEAK/
XiyAJ1y1T2cNa2Qsg973wCtQdxMGMu59DA78YMh6vCMcPnKa0w/0kQ7v7VtPmXwG1chrVquuU6Sr
OSiB3NkqTlZYp55PdXpdTfpH8PoS8FaRUdndQGRTD0NevZmzTUJTQEcKMYD8kxbKjziQrweV3CgY
dd1hJmUdv4Ib4xaJt0jPB9Uum86UqxJ9e8bKwwGAgVFNlzSJIX+mgshOFsupRz/OMXYSl63x184y
/UcvNCb/hmKCxE2k2wjuOxVlDEMrkfoAFETdJFXW7v5aUvEqMI2VupeJcbAa5PN1e+IkNyFMIFaL
gqXECLG5Zw8bd9XhbjHz1sbqOnOUNlQKseAF1QZSSVpGdgGAmzkNyxfgxiCDqsjuG6coor4MbFuZ
rUDzPVhnHvu+gp+hl9Litvm/EGFrhodsN9fti05LhahZByVrBlWdtPBMQH6awWiGQU6PZNqU44+5
PnT2ZWCpF7SqlW9aaeC8h6WEejrLkS6CXVzO0sBMvjNTFntsCa7aHX4I7mI0bjWplQk+QpSAv+FK
RnX08afq6e7QhML50cIwvSc5sKbWqCkHf45pE3sCO5acJLyVwPrPtlovMYcMovFbmF6wbTylLHU4
Cd+Sjfzl8Ezb8SxU3QVYdqauuM4OUFsxHCpWnJr7PhYeb3wGy53Pl78aWGKEJ7ii+F6gMJsNVUiX
Waf9jUC79YJF6nfxSrTQQJNlwu6svEAey8Ek+qhFEJ0rwbR+pYwp0OfsCAynlxNR8BsTZlL0GlMy
E3Q4Vz8E/Isq3sCxlzsHxXV9XGZz4OwYlLgKaO1BaGdzfesChMFx+C5FdCpazOttJEvaTRTvb+77
PyMpg2nIFCRTfm6jalero03s27j46BvooTPlPdaNPc97jNcpqx2JCH9DT/gBo/mZ7nACZihZTJ5l
k9Vw0sHqE7LnZOdaBw/I8aHTGDr0AGLLCgLGWxwsGOPO9R3JY5+gHCHWFD761H9t9mQ03dh6xBo8
9JxPw3JBUq4kdbnqVyZV49iIha2esfefIhjCKJ25SvSB9JYC1MXLE4IjRYEtN9K2xYVDFnaJQyb7
+uzR/Wwl5o1OTejsjTFD9dvy9L4AI1Tmf40aLFRaInRS1ivHxe4hkmSgepdOuqGHbIoJxrma5hP6
GlaKCFE1NN9HvPwXxVLK9gzkJ79crB5xdlwWyIGMvi/Mf7+GXGMlAFTXcYqjdgI8JOLPICgK+FZL
TE0vXXfN04eALpI1vVbVtTqAAbdudh/zXZoMS0UOwX1M1HffdcGndSYjUHW/Xdwj7fuJtcGErl35
UXfhnPpiGR9nvyc/A0QwGSltI+7X5cWPiRsoA7qGWssaXCPfJGQAE0N/G2ayt1Y6zZgaKNwO5HJa
h+8UW9o+aCV2mnSNT57dyHEP1vlDDRRtAFaF2z00QBsu2aj3utn5Alm7jsDUPGtT/9UPz00dL1oi
rc1/h0BNTh1WafzYQQduyvC46TTGlX+Q26P+zt+b4gv2LlykCoHe7gAHoed+e863Pg4t871V28/e
v76FvtPYnqwEK+fhX8FXb9nnXrAWiq4O3IMFhXSqYcWOQtXyedKBOVJ98V1vqJILHZQ06BOtWSNE
DNM3/1AFCExaZiF2AAXT3CFgY8OBrD8OHDXmuVXobir3EE7/a4qGQWo6oQnI8C0g2F5CfwZtvTgY
eMKZwONBp6iusGEA1jzdWNVupxKTUmSdOsNF0Cf3Gh6kQEXxH8FACQC0daxKqptE6xOfFNN1e8zD
z5fEejK0tUGcNYG559mXe6SNt8WWdXk/KHqsZYvNL0OpXiOjM3YjPK4wP+LggC2aRoUFjXrYP0ro
kAb/51Uy6IRUrixqHoq36ClUoFhhcKTv5rVYDU5aAUo+opLndDEbeC4SpJfRJOur6pUcucb5Oydd
mrLhOmkA9l3mxTPHZ17jEfceGK11GAMzGGACg0aSIxtmu6rUx/TPvXeWiB4BMdvZbb3umv7MUFl1
UHVPtmIOyySaLHWZwAwbr2nW4me8BLm9GrUFzG1MTq/c04hdyrjXilgu8SePk9XblkTtD6mJsxt0
TiKihLkuuOjViTQrrIokvjx/6hj61goFwQOxMR5j8c+i/JuDUtDAGZXTgoSRUtoUZbDqP/ERJOCn
8ZVRetWqra7Nl1SANLTAc0Dg2+xGIxYbZooYbWKc6UeFi3eeiWxUbLPJkLXR2tyMaNtxbSKZBY2M
S0UeZFpg54c/7IcWJLirEmSc31ju4LjHn73nloxy7XJJqdFjOw46upKO4iX7dffasUbPIM3qdz7a
H9w+NMG6Izy4T094pMYd+yZT3RJ1/z92lxdWhSHibHfP3wf9lpUvGLZ+hDlLd2BolsPQyMlJY6L1
+W71X7jLEayfq0nBhd4L/lLOrV6Iv/Um8bU5wGWE7K8Org3lHRSpAMZ+4eZyhXAXvgzkllP1w2YS
wlAuacuXxiuzK5bRyMYibEK3Xq72ju7ZCxFIVuwbM7F1FL4e9QVI/SmpVEDF15byI0mmAEZx/UmZ
vCACeGfhD207vfbt9D5DUT9IeCk307ZzlA3APAg6Evx2/r7BLTeGeuW8nDrGO/VtnF8nfgf1XzgQ
KcSmfjLE607zf0HpAlwPNQiTYYaHZ/8I4Yij3/gu+f5AXdugGcXDrTdqrHaWMmMdh/eXB2RZLSaP
qF+V068LrXBSqIlgXD7vm5myNvAL0x7gFQOQ0WIcK5aNv48gVomvInHv6Q7Oq1Os2aoo4mv/MyRp
RKW2awQnkPCjFFGnrD1SMF79R7b4O+WP7Lade7P+CpSO+7qOMvaq3Oee1RyWGssWueB9UF4DIw3v
EcJAVLBHaflvhuk7924g6mnyBmHI9Rhb+qHZwf1peKx8Nkq13tgtjmZkH07JDQe3wbRA/g5at4MT
/Q1ROeH/2AtP7EsGGwVEerbMRtgWIVzTRw1wnWkateNd8lVjQ/ms/xVAJFFE8EErgSVYKAdlCaqg
0VivgWv6AhktIa0tofT+hcNaFUOzSpGb+PZNA0PEofSHlgR+REBQlxrP6ZzfHNsJrv5OxUNZfE9S
Ws+CgysuAstcDe/yvdEIN5G34wTlmggSyKSh3AjSCJzjD8+Cl0IdvhadmuY+6igePnGW9q9Blifj
CARbX1tc82imLuplFuz37+L+HmK2K8jdMuODlaMCH503gB/fQoKd+zdwRlZzPDEhoW56AHzOdq1B
ZdZPagKQZPWoKxBKj4m7VF8swnF+JHUc7KA5zlNVeHIjGpFfCAvvJeYhjw/X3WyogA6L+CnruCz1
C2cCaG7Va0/umRHvCJv67OAAGH8FuiZ6amCWn3Dp4vpZhITqWaUWWChTTQclDsyYSyygwWzgN74b
6EXrgpp5qyNqZoiilIkWQwan/X5FxBw/ksyYIC1BFywKhxs/aXBiZmHNefCLZrD36FnCFjaYjS+/
c+fuc+S/ABDIT3YgwzEhfKY9srOd9zDDpPqqPeUtTqcIEBCF7OHdwtwPRNETS+ydi63NAcz7m3WQ
RpzCClscLFCCg36TwBfjrHdr+KIaWYfLvsFR+2hI/WdLGwuCx4Cx1NsoRgFrJCI+o7QkPcRq5wvS
VwvtEi4mU0UCCUcFtBclhus10ZzrZ/YZMVwBaL3TUZGQuoJKJD0+DmD6zheeS8usb/1+OthKFpXj
oe9p4D81Y4h5w9g+3uC1wILHwDgI96IIkLbk/JXluU0MCDGESe/13Xw8ga7WjHBDudANb5O2PHWl
pINSDAlRFmWBokF3OnKeq+Lfd/HtwYoer8D3yz+qKT84+YiRdNYjmPtL9rLVbnbNecfjw5gk6iis
rFp+ew8wdCmwsG/vIFbedkiol7ZPvfx/4jcHh4ZP9sTtlRCPPp3ZmWm7NMFoEEc7WZ0mK/K0FlED
whLKyU5vrI7NG7mLZLREMB4s7aCrL9Egv9sI8QqJAkqXickXx1JD68/KY/srISNRaxlV7ceAQAmh
wQAwXniULOOlHxsW+5axErg11HMU+9Y9zFwDtEuG6X+P90I0JNaE0SApywB7o4gofhQdGm1vNwPl
0q9m+tORzE+C1at8BgEXRR8bWECth3wsuyuXeP3XGeJh6rp0ur9YIQ+d0uf+iNYrgCrI64xK6XS+
/46IENrOA52GDeRXmbfOgVjyi+gZempZONYcEsT12TLTe7sGx+Kp5Blqg6xxvgRJxIHMxHQYILv+
7OhU+0kx52MK2MT2MJ4orainPykHYDn4x4YmfUVFSKuc9j4Vk2iKBGDnY2uudMPQY0eMA1I2E6JQ
U4ocSFt8XPKqngFRm+gH2KsQ5by9YsN+XGGb0w7rW+nUkuuVeIbLgIWctpXWlLGzX7gmmL7Ab+uK
5PHihSVF9RDYK2Zz160T8fpfWJ73aS4hwcZrXExupfhYXKJ6Kz37SJW4fOAmH7GwiQoYUPUAfq/k
4kMNngdr9KtSJK9USZH0kZMxJGAdNkFdt+w67ts5U7H1tMTG7JyZfSn4bgwPPUesLX8OGocqUmMF
GLQnjNoxyhjSmZc0GyTknCXk73qjRC6l6JVkeBjgBWMbn4SnSvZiSdlIp6aax7+rXaOvh4U4GepJ
hqbJsiDmcq303o9lB8mZ4x0Ly5sFmj5WYpoT7tgS0P9yp7BKdiwe/ZakSSkgH1uoD7oNMl3ZnvPl
OO5Q7XjSFXocUZr3v5/ENn/M9KbnZY260+wlcTNrhcFY79SnT30ihF7WUCE/59/MmtgsKGtWKBGv
J8+Kw0brzXirIn7KFodjGUT4QKvzlZ26JPbx2U/ARBhteYlxEUqgdi1yw/HRcw7ZSG15imkPp4HI
WuMW+U2wkA7Xuc5VJcBXkOkuiHqSyUM3ujp4a29ajt+hxxQZguT9Ve6+29pmalroSp6fl9ccXmNb
Paipl3/1YxwDT1kpHDPoJZAV79zuGGA3d0BcpyuHSl8D/p6xU8Mq0pr7aQFT0PBx3T6OLLYJMDJo
HvZ7044Jwhy2kyoEGDErThE2I6YFoh496bDJuTVBIrfBbK+F5KmOVjyaWu9SvJLwyKnbiFuqKMBk
lnVc3Gmp2KhTRRquCEKZgYpYNd1a2Qxfr+KfSbZyQ3vPMiWUklRLKX1TYO3LzyaPoisP6Csu3Byw
vuF/lz4yR+aT7DC0NriktYzfI6auU3MB1rZGGlGxlAPmyX4uhzwDcHP9TR7by4c3sfX8rePSAi1M
7Ic2AU48R16COBc+emI5c34IYxGJNXbLkbFHWZeck/ZvSJkYjNkqch/rTUL2vmy7XQrrOHdXDYwK
RuktOz72NYfKpXHnIAOR35t9Oru1oQz4X/i2x92Q3AWUUcxAgAiSnregfKm6qvrEMHry8qMNcfCE
oB+LxpAaJaiTRBshCVQqWKn6FALPv6NFHgqM6Y/+st6GFwxZspMwGgff16kWUwyUUKz1w2fG8VB7
T+PRX1PIo+TSRYCFQqYtT7BOsnRSSZB7VPinUXFJmkM0egVW21c6mlEAWHOJUQvvGr9cpCPSvRKi
M3hwJF2z2/QsVZs1P5k4Yjq/cPcCF+CLWEFbWjZ8IF3J15ZEVFlbRUJuK3L+EfVYngQc24mpesr/
ThK9kZ+6f4yduNbRjj+F7M/qkklP4kySpBPYnllccihm9lASbSrUwIdi7dUp20FtUAURaZq4Nmba
vPMkR1OkBl2i0VmGloN3M7MBfHes7SFsbB4K1Ku3j0k5nirTxenmleSBmWMeQ31GY1xunMMVVbvM
spJS1zTfu/aSb+LYTlZfPmlM/jZzRPCSEfOw/CQorBQqeic4TSEznKCF9X/ZjcBo5arXivSnWSZU
UiyYrSrRhrW7/Nef3pvRKbYeRvDCoVDWNQnvoBh4SygYvAjfrX6l0Fg9ZUiJcI92tZfHQlx0JDxd
yrBcgdcyXULJBNiJIvfHgl67CNNtRpEFi0F+g3fd8Bj5TY7+uG57f9xFtmsmYPBU8SEm2UEYlZco
FLcVECtT+MYJviRAM1HsSzT+u68ALw+o1JnhQkQPjG7t2e5goHAuFDFPEc0Xbg1Q4vqqbAeS5aEN
y89sBafIDotwbiri6Hwucv7cZ6RAtq89KH5UosikrAlzKUmOMnFs1LDSHIYzuj9Lp1+6tVxQs4j0
mvw8Exp4LLeK875E+HX65etBF5c7JnEaUB27jLdI1J5bdrhJ0Qul9Thod+Y0TmgXK0gTDmX59rZ/
zErqjwaTP2qlk1+6U5iDje8bwnQ8D2PIirWBmVMJ9g5UAbpMrJPQ11h8OmhqXTxZsrxO8i3VGmEC
uLNPIONrrZXGeUMB9rviQRyjnSR3L6SGOFEWdYXiybvhFGaqXMTapTCkADYxviwsk/evQLZV2R4D
rRBEAle3HQ5qj24KkyMLH44CUGy4SLhACGWEUuO/TKOGKXpSguPbzVpfXq/ZWdfwuBNzkbECKoxb
Z1kb1RRiXuzgRqzOXo018jxrZvtZmvJH7hlFFApiDCR2WJtwP86rZ6RAZRhkpiv8B0dvqX07STTF
Ys9hpa9FgYkL9b8b2DtZIgY8ZCBmQ32N8//e6Q11ThU7VBW5WwTRuoUyILc4ikuX/T3bD6wf6yNs
FJdw3iBZyEoyMYed2im8f4uAw8pdJhpXQC6geM+iC6EqaaBXKzL86fvJvVceL+Yfmgw248JC3Zso
RoQV3nS8dmPCMVPcDLojtHdO7p8aLtSYBTBEoE96D5jIczk9manRS9fmaWremW9biUq2TurcYjNN
xgMVS1b1d4MV8OEwXLBU+bd5nuTcf8EGPpbDxWPooIw8t37pLQeQsH3lRi1dSybWRkqAk0xrkuVp
E4TL29AFMbhvpl4nNYQt/5LSibUomLJgfufrO8phRcrAzR5HyEz6nI7XaoSNU/F/EE2cGpKDxz3n
RC/kiOX9gbioaAlmEjJQw6Vt1MQ4yhgpLh75WEYWgAbRDcoFRYw52h6E+BPM7If52QAqZEiLn0Kw
Ef/37w3LtEkwX4B2pjk6wD58mt1k72sWQl3TfdY2NxFdG4AW0BzqY40So/UX+5VkeVAZZb5VU33R
z2Aov0aj0cMio5nQbvpKdN9QNcAdkffZf5Et3rt6UA2DU6qwYLTgUXeVHgx80uG7fPrcLKaqwh1H
zEoB6iVBPw2XuItXIj+lsd3mbgs65r/O1CMTxW2wzUemNiHm5a4oHgc32l4r5lKiwHfZNbYxu0cG
HymmudkmbpcGfvpYtrIzvqegSqYOlX5bjay1SjjsgM1Tchr6H1uYgF4pxNb9L4fQS+6/X76Wbv1q
NOSWwvCkQ7gmMcqL2cS3OyTPjEKPvjpysIH/CggpxPBOeEqz41i0ebpaRE2iYiWNZpVC5QAY8u5j
wtShnf0liaDOkJMFzZHm+RUXps1xlF+wmg6vc1VIoipW34ARzXvPCdy1tY4as7DeMV1FH/z/hUNy
gLCC+WPCOkvGJxndzXsGEKTlN3iWh3pkq+CwIB+Hg2PXwP55kSpci4oWYLOsAidLPtxBURhuA4iD
b5nGsXTGbIxOMguyhHHEj3co2HzdAZzvlrZG8WI005j/qTmoris5+ihDdmgjyK1tcbDbmTYLLlcv
8oigWnAV0JQ1bTRDTqJ38Tww4G2J/7Evyp0MEq1dpe7FRvv3demxgrpvMSifGETVIT1//xN4LoAE
q6Had3A0QdhTm0OBU0wGlHPb5ryLq8JffgiOA2BkL7E5tKuzaa6PE4JEHuww9cbVM7iXMRAeJi7q
y3NzOd8EmIGNXetEX0xwIZRf1dUQOIQ3+ODZ4vjQvdxpixGInPjH1gy3PI0yMiK4Fe+zvFCQNTNY
SiTCi9LuvB6kJzEJTSlVFOkTXXMEbjtP7+p80xKFPOxSEpJl1aQSNE5EHz+rTrGjpb5uCDJQ38st
d1Xago5WBhd8pAofCaGeDgG41cjNBSzwBE2st1+RED0vP0J//RHBHiYhG82hn4kQG8Ze9+PJwbiS
ykl6JDrs/S8+AYMOLU03ZvkATuAOINMY6OpC8HaIutMgZeVrbjNgr2wup34jWtTJgPL+uF3eZYVQ
0NIqiMd2+NcvgN7q7L3r8sN9DElcHEVZMOakmPdJ/DEQwyoCrRr4HghzVNdmiqwiWHx/b4rV2Dv8
WpISGpefFS4wm08e5QWuMszV+W0j1+SbOQ6q5SK1XQNXUuSblfPk33+75rgFFsqLXHSZy8hdS7pG
QM5KXy/lZpizKUgGUqWHMlqX1bEKwwicQ3oYwHypiTMptL+ZyGAKgBNUO9e2XMZPflRzBv79zR31
K8taCSCHsQe9wL70c3k7Ml2h+2QJkvypGsH2H1Ks10VOzD5fDAbLdaqFzLmsT6SzHjqzvK6lZNUc
bHE+mHZjSrMHlmcuYBLyz+qWcbUSIwUmExvBJAZ9bjHRHJ2RQ87ocV5DoaFOCBxeHRU+11TbR9VY
kA9yfESUsffTIThUhFbpyoTNe0WFtgf90L8+LexYuFNmemSI/PF6FyG1iAf/YMhpEPQLJsVMzgra
2GMUPuMI1oQOg59n+zzqOD9EnL9YYDsME9ayvBbZfvglDgXlQYqNTWrQWyd4IvHWe6Z0liQzcz9G
CEnh2EYUYjNXmhstFfmlQot8G4HwEI5L4cg5XZFvKHSVcEcfmZJMFDj7GajPqBFakOrveCXBNt16
5E0dEJVoyA9DSZy00IhVDse286Tey7hcaN3RgGjg6yBxvmhlzdlr59HGPlNgst7t1CLq6V9bcCwP
OobUZjO4RnGggSGXGfs7JCzx9RUqvFW+cBJjG0XDTc6sQM27CA/qyuQ02XKRXE3lcn/0p6on1PRw
6e28BD5z7aOSni/MOv0+PiSaFodwD7clK5CdIRGXuELFs2k2mMrA6N9edPjWmXZbik1TOVtpcTy9
R2CMrHO8jXZ8BMPceLdtihCRcMRxdTe8M4ZHm86jtAVtJPNZV554s9Wm0Nfdy2XR6MU5tf+AI6EP
a70JKe+wCaMkPNEGICfu7Jjf9oOZ6MwHHOsmDKccpfigTRDBRrNO9xjZDOER5J7XVPmMhZj6eZ8f
SnwKFgX/lyqR1PX2ambY6hXZ6tkSAI9v1v1v5IRiDUhzFgu/zXQp4Im3QUhd5fw4nOz8rtVwMtd/
PsjaI0/Xrvaiv4Xkec0YiHpTt/jrbvJKr5FfaW6V5o4mFUnwi/vj2/terb+Jxs1VmV9ZpY8ksqDW
iY/JzNfdTZRrQdV+0z5999bPMgBqvdEJ+np24D2le1l/L77goSQGKCd1TrLWkIMiYmH0fU6NCGvp
jzGqr7efhEZkonMwgRU9C9ffQYnF7Lh/i69Epi2ZZh8wz269paqo4vGITSzSYPFt3S345U1l2qFJ
ZyFKe68n7JWySjNDBbQm/N3Xa0K+xRa81BpUoN8pgEKrIpTdNAcPnL4OajODGnMRPXAV8M/MJBYy
A2K8zvY4eaVyrdrf6HqzuB/qzlp77IoNuRXW+yvhzai0hyiHHIwurDKpoOI3TSpTkmtgOuQVC9ad
oc3O77/iBdabyQMsyRaaO0SFiM6Gw1Vft0BkxukSz5nI1QJAgHpjZ95Z9cHbpbsksNR66SUz1M+O
hiwW2QTARhfBON7cve6ioxiHXEDfM+95CQwDl8i2qRnpTn3p4xR1i/Sx8eOLRi4OtQMV2zTSABPz
lLYJBdHFPo+z6IXvUbTwGHhB4C/C8y6sna/1F6I9RpruXDLCbxz5MMGKWLzj+MdbeHYuu/uy2C2M
54c1vocUANM+ClRcHysBNSnwec35MkIVjBNnVqR62tNk2kihy9N75PTwUSSjosIfPvMF0mSsGia7
CbSON2KKlJDOuBassng6vrz8xisVmbFMrHi+ThBM/BMoux1tLiGIoau2yVN0lotepXXnfetTstM5
RZ6y2HbPXa475fzdcqd1Bg1wcilfnRWPsGhU9Wcc3FqXmFqIsGMyhg3erXk60Z0FvQHQovQf2hY8
sO1brSJnO0/vxS7AJ1igSyEElPWssKcQKNQ3wLIO3TbIL1Nod7mTID+5KPC8mbih8IPRArvFyTc4
ucYQSoGJR3/F68ellmWgMqY/UM1WWzPaJvPmDpjW9mph1TBz/cm+XXzjQZG4QYIz4re0gvKDwaqk
fEZ+ef19eJ/D58bVCrfkE0U9WXgLYAGqkWvwIZ4O6FQuDNKgBqOOqkR7BgLyQgfuq5is1FYatSQ/
3Np3gj2BecSZ8ZqfAmFpvveONcuWeb/Zp44cU2VZN2UcP6aRv64iRTaow3SdqhnEUuwSL49hWTko
SVBf3GVwzFu20Ez3MUum+S1AudX7ikNm7C2gaoSDtpHk99mKVQhsD8u6zpcquS2e/2uxQcYS9bic
IauFmPuf6EB9jU81uiGycdkrOfycnhS0USiALpyH0buwcYjyfdk+t3lTtzQ3kpxMsibNfpgE+Sum
rxn8/Y/5rjlKxJBZxwJxHP0gmKmUNjCz59Hff9TTRJmVffvABH/CWV4FBNELKCpBFofHqMHtn1tg
ih5Jj42MTlxh8N8LJubh8MKyPH+GVSEq1a/nvDr5+CQR2cHoIqTZGaxJPQEB3R/Cs+tdlwhVeXym
0F9Xnu16XvjnO4VQbesqpqD2RKMSpYsw6fWTOr8W9czWK9n1pPOaDl/WYxma7sIXMiVpbzArXvvH
ScUBC9Fr33dzdefbGpkiMBZlmclSrK15Uw8S3/hp4w8pfYhzJuefpnvpyFx1novGthYq0qloLt0R
m6bg4vVJKQVe3W38g25NWmrHJE7nK/rlpXm8Ehkq9dKItSuAwIy9Rp3TFCos5GTAZqaZwiZvGtwY
LHe5rggoF0vIdr5GqvJkRoif8q4JfXZNUmY5LPVM++IepH4pVXksshjomEpySjxAicl+SQ1OXqU/
eJPPBb73pSOTiP+8cSwJZFKyP1oDt3mm+yDwNGfYQsPLZOPjAdKxPvXPAaIzGDNrLSM+yPRxdLoV
skRI4uBAnxy1SwcxPfpkWMECL4vovDK+H+i6toWUM/vM5ntNOpbazzYo9K1mOaZGZHaNJrVYLZFL
WZQ3jds4hjZVzMyBaGO8Ajivcekai2bnk+oXa+GRAucKUgOq1tedQKjWHxk8ksxkchMSn+b9N0UU
pSNg47qhsU/Z9zOeUdn/uW+O4F/gjA5eYYAwkoQcB5NugWB1lEdak74teUhh4Y+s3GQEKXlHoyhe
zSJzDfoPaip5h/tRqC3pTfo26PyxHFbW7G/LGMNsJomeEeRSgS22AA6EjMEmvYwXYYG0vmycWn9S
swcH5siLs+HNkPS+0gHEESQNNnlDzu8GcQlQZk0c7GMLNY9rBwg53NatSu4Im1IMWyY80O/L2mQ5
6JTzgeqJK+zHUvEkI3GQJdYiCln2HC5XXgDX63ZFwwHqjNgOtq6tqOb7UBabKEl14x7MEdefE2ET
npCGkrsr/oX4vKEHLf3qsgqVxAe0Hnybje4MYmXMAACk/Dy6f3L4UdiWH+1/xzjaOQWtIBPTh36O
Aaea/PPvRFi9bDG6f3IsVgUjuxfLn14/Ax0060xlsO/4hU8mrC2lUwIiAdEqEI/kZOgaLcxeUm6B
OzOSibRyDeGB5/ViQ5cCtIYZSGQQWSM5VR21IHyA4zfOACftPIuIHPVwj8639XNnl9GRRQqtU79U
ECXdrDrjeQhvl+pRKgk/RVJcfpTlmyY7zO6GCMYAJvbp2Onuhu5PBbrNWkXLdSagxsQ6iVCxb5VZ
2b04Lbp/xLy27l/P2XneQkc/rF49RytZXXm4rY3QF50SNRA3aZzndlRB4z7qy0olp0N3z1Vy+KZ8
KKdQ00I6tgD8aOHvCvd7uBjt3K4cYNiwxDh4i1/d8d0ng0liHKoLvsB8ogVhwii1LBzJpzuuLL2b
JSUNkSCOVVFcvygnOcGylzJr7CfCC2qz8M4vJlnXSU//SLOh5DWGwttji71uNRkjHQppZN2Pu3X0
hq85N189PjIoTNGIdXRP5OmS80pNN9AA75ox79kqzCbF0fNetab+JCO7zO27XKnKVIt/NZOqT1l9
qJi8LDmLyzDU+W1GD+xY3B/zm0wJPI1Dd0DTI3eCnC3FRPEKOHnWpWEvRLeHV+lygxCOCZyvjgv1
cnStFSkhNUwoqSmKdNGRZUISJHCWwpyoXdE6wKJxRYM+j27tyLHTq1i3ygvtgXqnouoEuocprJoX
hVgtZG9IJNxCAQfb/arbiDoVRLwhp/mP17Cz0sNEhQz1YtYQwiB8Iz15883VTBx7/0cLuGiog4Ki
05LrtHY/RtacFaHGYcEOgI8TYaQn0/dObU1z5feWaV3UHV2KEDNwdCjr1XcbwXCMll99u9SWaoI4
8VsXPa/u/SExKlSlpNSudqge3oLNB66RDmU9jGeKCQrzjv1RBtg1lNM/g6r66s/2n3U6nOTA8/qJ
Jqxw8oA1T+f/JElpcroQMjP2yvsmDeZDTpFq2M4L/oSntMFJeXww/rgIP7S1GBV9wEZkH5X/Y+gR
dilScguN+/bphksR4RGIwcs3m2opkBfYD0r4aSg0UnGBWQrKjEzZcBIOdkXW8lfE7Vy4hUY9DzFt
LJadCAVTU3hlKLZLDqlXF4Njxm3+wdZfKE2i5XpEHtwuF3qldSq0LlN7igTDaaeliDUwR/cLWWY3
1nInWcdAvmlXlqzs695vlYkRcsPxySFtLZ9gBk6ykO7LBMdHDJjn3/VYgwTz+CrCAvWJDulfMUk6
IpjdXIhKAeu0Zxt/eetgPHjjizv0J2sawA530K147ykWTQtblsUMHCvcHp0Obwb3vvzmS4vTNKwK
1ZGzvifj+la7CF50JfySPxia8w6VkOmg12Yig97xw11fO3zM78CYM+PeZRATtXzmqJ48MVcyXmfX
qEtIaAWJO2HpFCFHmp1W9O2tI2KlEb49BcsueFW9f+cjgBZsrlC47fNLCKHI64HADMJ8B+4yhxfd
nq7NvoAFiC1CQiVTQqbWCYUne01xkz+PZ2gvIvpQZf1ntIr/crUhmJjJ0y9xhLAG1K421bOkDDNh
BOfk/3AnzZBjpGn4UcdPm9B+c4vnlbjlTMHNn8JHxb5aBJHSYepAsveJIhQJKW3+LqKKLSvFQpTh
+63fcJhznMKGdaD2VImwzgGG7y/ZAHso+/gsTdVgL01wztfLdBOJJh+arzUHeLQ9Qes7vlpNW3TN
oSqtGERZtv6xTnosnFZObstmA249daTTdQV3ZW2mi+InIWkIdwX1rl5/LaVBShPzEUPwYyCrCFou
Ktqo8srwnBAtgyXvPupn+EIhYDaDjx2KS+kT8EiiPdGt2FImBun5DqcAoJ0fmMkYYqZ65QGhx5WU
fkMbTtcLWYvc//8dSzkA063j8XSrY86trqkojcQxixq53sr8r/9xaZnVAAOGj+eHbH9OWI67ePOL
KJSgwXiDWowldnZgRx3S8RCmdLTCrelMBKhfthbPgYXNUBdIeuWnLQ/EMOPn8lMRkn6iP5NTcV9C
ZmgqrDkH3JlQ58bo8CGJr9lv34XKX/h6ONWgIND50c2KWmc8zbqzW5BfDN2jvlaCuLlktx7Q2emk
nGf4F+wsA/nc7BfBz/pfFzCBYPtgBJe4fKgX9W2r8Su7zG84oE+LEWLAEol/jLz2YHUPueyetXqc
fkzMh95QJvtkQwd1qWEP6HzsNkSI53mRCtKtiKwozIj4zDwmZWwQjCYw9R2S1LD8aZcqlVVKsmb0
er0J40pV/Zd8QMe4cA78x6BY9XjpWBXzvNWhDLu4SReLh0gxgaMrVDOMWiyhtoCROnQQ6Mijk8p5
8V9VmJdQKvIjzHC4UVDI2WsPqLV21lxbyp2RxGwqyUWyxcnIyMetM13THs7wl/BLUfxfOr5ueHAM
8hEO+KvkPfmJiCthCM+kQ/dhhtXWEjQqXqBCMzMXhjgcmKKIElaVVrk3h+Kj2kOHXo/Eqg1Noc9w
oOVKDRrWutLuqREOlI3j7aXsaRhg+iQ8LZ+LPN5D24QZccFXAKfqM/w8f4/e1LQvv12HrEyeX1ma
bIQoteholgEpdQXmBqfhFG7W+cwiZe8660HO2AnlbZtK6x0PFSUenLnrXsY3KcLUD53AY3z/v5QK
vghqjLO15sOJPjfcKb2kn7iGwENb+LIWf55jG17Eyh1b/6zI2o4Loy8X//bsNq5ttAMBbD7VgcN9
YMiK7DYsIhsPbYpnnTQXkH+P0fd1JG+W/Ea83tYJIw0++0RP3excOTydMHVvjl+21Ukcsjuxi9jW
8orXp9uMduZMKgnmkvE+raspnO5+H/r+4p9GhjnzXAWSBAsdZRQFZKaz1P1DquoCEcW6nkKAsRrm
pN62xNb6z2es9wTk3acaDU0+d87G8iQQnROtDNjRGzcQcSvAjMb/fUsYBmuIwmEvBDV+2Wh9fY82
Mt8s5otPceTeB2SHWRACuiKJVntAGXulsZBD6h9im+6G8HVcfyqxW/kSNDKOjfw0Ukt+i9cbaWlf
Umf3jon8BBaf467WfFJ9iyHKQhzlmV4OYIfH3/bLipW8QwqjeSXF5RZN2DAwfOsBmIIgCWTTl8dS
/u9OrEHnZE4u3QXN/thkjAJlJBkBIFguKdgH733NlnclN+jlZ32OpCJ3Csqeog9Gg+8BbC830u/S
e58xTfHZTZWY3QYMNxPpmN2+AltlF2TxvclwefDpjZyZZSWm0G11yZH2c94Uqfm+9oQmHvjku/r6
7VIz+3PFLwKYKR5hDhbgGVr7R5Yu6f0vNETzN6VPI2N3YGUkx0acCMNE1IfyGpSapMu8/GzD+ACo
gqaZCRjq9py60NN3Ie8jdu85NMFkHl8WoST2fkZTJO/bzmeVGH2EekJrLqWDWYgxDp1NEC05VWiu
MYnN7APrt03QgWW9K5XjCWTug2DN0cAJM623hC2alZ1eYbTvXPy/03sp2hwspxvzYTX1Drnv0Ye6
hnC9QxXM4n9pLaRwSapwIUAo7B50eaV3K0tIn3FPyJB0jOddu9o4sWouWvwioVJm7oPGoC4wfdJJ
Xs7IS1xa9vL14c7qaDu920SocrTxOEbXnJW8sYUZPw5IZmZoUeqhkKVQs/X4VaUwq7TxksoXMNjw
iGryEzBoxhMaZ1BZn8JbvsvjGTlOClIV/eB99FN3tG5IbVhNZNf424dngLbUJl/ylhNXZM9AI3/L
qu9kg5ySPVmkPDC+MRi3wVrqefbxKz/WN4+ExlwSmoYpxwVjzg95llY7aoIxIWBgoRBQo/sFkEFP
zgBrtOwO2bE3D6z2aQ2OmjbadkCiT0Ndzm2KWDixtke+GOfBTPIp6TXqVM66iqkueAbceN6DupnX
ZUiljHKMMUJ/qOWxUujF5HbnI6J/zdvSbOKGKy6MC5BmjVqF9KKO4Qnb2lvqOzcxtmsKVkNw8pJK
r3EQbQ1a2ZwqTn61hOXLDy6o8ECHwNj2BX6Qu87thhEg7pXFXWiSPlHq5Ibqu7exicue6sB/YFsI
+zZHMGNCDPTkDS5eEzyqOp5hgsUmFjL1M/i31I7TvyT7T08x5qPMq8PN+4Dz4Y5XW4u0aRYsK+3u
qBiVY/1HZ0gLtI2tOYcKQsCZcdXTYWd0adpMo2txd2QSPLu+15VTSGHXgCFy32N4IlSRGh6FcI4b
PRd2e0TU+5BLRdia4pIDbJx+d/Ggfbu3d297Ea+N664Xx74BWy7POZ8E3tabN4kQUgmO6y0WEOoN
WZTgHJQgrijn4F0FiBV8Bz8wo6WoQZNVyncyxFbgkt2cFo4rnR1VWWu2WZ2mLUx0XqhmRF5ZAiuE
CDiWb+Gb/Cc/Ir0O2sAQcFT9f5JHT5biFXk7Fg7/MDHFHWP63QXOhrM67bYBvpr70USvoFa0xlSE
Pa8rfslbkDh8j64jhXmpxRzeifgxLYgEbrvaUsg5Mvgx9hAwB/f3BE5ufcUA5xmFKltqt0dxsvwj
02CPFCPMzaCNwc+uYQV8wRriLc/XG+FnJxmdE9t2kT/3CfMVwYaejzqes7/S1RKRUsov5zLJ5gTd
T2ELbTVmAUfOwXG5V8xzHDA22at/Md8xf3QXVmGHXr34AqWsUeuBvDrmXpGPFPuwONh+YVfBXeeB
seAKwzF2RajCKUVvoRRgeWBbKH566tVZaO7MAqeXh55ZWA11k78iV5LN0LNsfZDVUE6xSgYqu8bq
rU4J14bb5I6P27kLZ44hRe2piMKZu0nXWkoZ42heG59CtRX4ZnYiPfAGJCLuWEuW7sBPPSKupUFg
nx/t7tJKzewrHgoidwFQzsTZKZDHHApQzCSquyIqrfKV6+56F6H8EgGculfikXODXwSq7vrMXCww
u4sh6YmchmVh4lKQIdNufLGOlgYyJEpEk0zcwfZoBX6dTahvdsPj3ut8FE3WBYkwS3T7gN+cbzGC
EMEjJQGgIcFk0hs2ok7KJsPU1oEKoOflVDnSnPbI3dGs+uZT8pw5i6kFzoQasfXcif8Yt0xWToot
ocbXyE36/gp7X4KXuYUtJ8madCUGaIzxXJWSFQgJok+kn76tg6LM4WrvcYTzCIuoNQmquLgEKj6f
UTbSqncgi0hMwh40Py/TcEPXjhkKgbNLHCV+Dynsjf9DLrLvCzmrFrMiNFRbS3G5twPFmdTrm8pj
C5WNJd18AM+sedDgY/KEujVfln8L625vs/sHo21yXEsu7+gzKysmytiAnNRKKY1dzceq6zdNGcvZ
2OD2G3efa0uxRnZ+iMuzV2s6lAUYclmUzYl1SwfrjnDmFqjGcbCfcjuZ7dl7MZp6rOZ/4HsKgvqu
/ImUrELjPj6quvuc1IbLxZbZAN1dmJTUwQHUyHnx3in6irf33OYhx6REQCWI6U610Vcja6Se40Rn
qfnqbpaP2nPWykmzf90GBp0yEwXsxrDZvc1rV914b8rHS70v6mgppRwoB2P+S5l7ppqRf9GCnkiX
VY3UO09jcVn/kd3Z8ADnEwMhMmGdc1QfZtgvZpzlhNhaxr0tcUtvEfSJWS+MHBkEzGzoCwgWbINI
Yu9Mgchexmh3wz3/3cVUcgmFBJWYtYE/UUXn9YAfONSyGkQ612mpO/+GMi5fe6jKt+czcUvB47gl
taWBCgZ+T6IqxzrObXJyq7BKTy96LuwBxpcqQmStNxTYxVs9OSykt9WBjKv7j96qf0p8mpIQ/gZ7
LagdvYyzaPrggWiPuzUX5t80zftHIy9/8WeLbjNR28NA4gHpy43Pi7qQsL9XYa53YAFRK7wqSWRl
GOjsrmVHI/VwhLVjpPR+TiunLBw+n6D6qTd/jCraR61cF0czy1psquhpNTA15P2PRa7yWtQgr/qB
CfVDSw0Y7l3csqc+aEr9Nz0vDSyxUe9qYbKDlEO/IuFO31lpguokTaMjNEykEvvHBJ6ppZuL/fNs
3BTS9hSpuIAjh+p6kZV51AnKu5h1gn3O/bVKicI+gYYnoSQ9zSxZquII4kKg75GZd7aJWcPXnELF
8ruN5X5UKwRLPvBVg2ZhQGIEYsvvGY8TUPq3fAN6f380LcKr+ez8afru3zqnCTcxkxfwmneVmZlS
nJodZeLtJJBuWramF5KhBBieSHv4ozWRejAU+IQGKbfc/Ce7kUVfPN9AoRgqzPFN3ETZLozaq/bG
8h0XYqksLNEPFCnGJrRiCbkPywI+WBl1BzUnzniKVLgnQ3qsx9xUKN4+nyjRBezKCq5gi3nktdfH
o21CdsxK/Nh9aX7p3ErG37+JfBT+2g3GgVhsaH1Bf7MRMUe7Ye+15hNLQV9lRjn5UtPdXkIwMiW3
tr/4tBl7HBT5Wif3eodrdkdWIjlHk9MZoHk9yR4rOi71OIHS5AJ6/370uJIn4gfDbk+9MLyhkQxj
G9A7oqs+2IVN9STR256lDEIGmhmVW6a5yu0U/0sOEdNjWxBMnS36ELCY5gNJ/ZMYmD4CsXBZqB8C
n6Vx8YomTUSr8X5fA3PxW3CXB9zUWtb8OCgwi64HcpUWGSghJ3a0GEXr2I6F093TJ7aNOC3p2n7G
yr2TzWxRtCuXmuj2Pj4v8NzKmU8Oht0dqw8lLtAcQv9Je3tkjg19wtjAN8YXMs9wRidILTJnosuA
gthzlOPXO5WTP0w7XqkEdQShiOZ0IHJsdvxIRPFS1UfZz4V617xTRy+821QiYSnJg+7muUrdK10P
4vyMSUd20XsluoF9mAAGscFEXR+JWJqZzcqXR8rwfM26xoe3ln+GsrcevF7suPJ52xhdu9me7fx6
t+jQT1dLf8uPN/w9aFNFC9pVYQS/XGbnbtKFBP2NgxMYHfYATYw0PJQOkjUknSzlFB3HoGAAaWGk
ih7RzQlU6aAF2RLIGqFTn+KuXANOV1iPwHPZsLQIm0yqoLSsfG6Rwx3k/q9EEOJRRn0O8riVkx7b
IC8PNpydalkGskgahIeZu5Efa1i2932iZbMurezm7YspO+2ZUDT3TN/Y0KzZS7FA62JB6X0TiBP1
MtFCkEZ3YGXh/HKM34Ih1z6vbbvca3N551/Fx9qSZuHH6P4iDN7Ors7W0/Ex4TFCHJUx4qGMJxtz
1ceQnH4qvMwTjZPU778VyW28iurAfGy0Z6ts1s1j5K71Rrn9lbkd2k1TS3XR0rZPhTHIi/VU4pcB
s/sYb1vMZMs4FI9mEqYx6USbaHaswgzI4sfa3rjRRCNewIR+UZ9zBXpYrd1hGRlEashLfBqcxHXP
YwF/ZihtWkWA9oQwwB8MXjoJtQEGFkOtg9zUEsY1ujpZ5sFfqTA1saMf36yHE04/OBohhMaTLt2A
7ONoN3Kg62Ov5OaAWpLLNAl23rFd0CdvOGbF02/MNSbEK6iL/nnqYI9dBhdMF6hye18Nj/sQ4JAt
9K8P5gsKFsGMxj1JMsGVfe5bi2/+pMTxVa3SvLNOYOZwv/lXRCfrF/G16OBSN7zLwl7Mh2gY4HSv
5J/q0nEb2rSVxtEs3DZeuFDG6CaXGQ4ElDdJ/B4DZQC5hGapPEFsGSdjvR0t6Yz5mrh2y2NbMpUz
XuwSpenn2AQyUO5qA8TR/vylHFdMEXK0q+oY1XKKFTopo2xIOi86fTwHUV0JMG8JdfSLWAlD2hiu
vc6ZlxtPCSDMXRwa6SbF0QjYjarae4iHHmtbiSwzY2yS3cx/tTSFD5eQGhiJXAEv3mzhHJD/WcuL
E+E+TZKOSOMVg9BU8/4FAzjAHKcN9UlPob1Kz2KnWYiJrTrMlO8VmK8Q17lqje4xyrI8scjQx35m
gFfzTRrAaGDsZOgIJFKnwYfP6xVrdFeCtZ5VGxSZSN0RjWcuUuyqX6eKiBYhftuPW38BEFdNlkmU
lSPC9u6/Ni4h1ZDuxQjgwjsQxlOlBy/Ck3ZMjB4hURSUak5+JrhQwR3z1r1kZZzRotwCJbcv6uem
uWoKNqDTcrf5u+w5YQZrUONXMH43+c3N1TjTOlGM0CaIjPeyYhP5tBawdCnn78FM5VbRQVfpiC/5
Of2irOmBnSpDWGiUkVMI1/ne0DiRkoFdoF+3tig8RVXH6tY5V6ecuprvaXk88hsUf1zTc54aY8ns
BHLygdRRapql3ucrtZchROY7hhkIyLkvnGtM0P/oBq6XOhhq7u+pubtcd6Nsy17Q53O80OVqxAZ6
6W4RtMSoWxY1DInc91FIgpjrTAKvj9Jdeo/3b/nyPm0CmRa/NrNEp+aPI8vLBQqInGZqBVVIEsby
YQZNAAWFrlsuASxgFrBV4KLepfJeOHjgMP8lzGZkhgNYZKLWvPgD99i9/jat1Vwuv/bdJrtfNYI/
hTK41Zp6olPsTEZTsjnC7+BvN+0TH3xpLcK9/Jvl5ITJFm+j7FhJJi5UUs1n5uyCgeiE/UM/aWad
fDD90V25En5bhjJiYb/U2Z63ojq31gBZ2Las0q9BnnaDp9E648m9Dzh4hx9JQBpEC0UqcBc/S+pu
TH0Hjbx4XK9qjr7FiYflUIdc/kCGZhpSa76yBVCQcAqjX8sisUqJ3i/YAPDcpwNJrKhePHbECp9F
qTyFdyDn81b/hkeG0hAupkQK7HL95mU6sBiMVfy4DHytG6WMBn6xyu6LyrypnGGOE/3zpvJZExe8
OVyXLZiMGX/KIQrCtKpJq9hB2fcay8v8jmbCYCS84Ak8DcuMZ9CSS6fEwheqt4R8BJ7Ci+K+IE84
PH02sAvmBj38zfTChV6zvv1Vxmrj2t5lO3I0cqJgb2Ichec3bN38nJ7sXEvLBpnBjGYX8xyCmpzR
/j6i3mAaMAVHfrZbu1KsyDvW7zzN6sykmveuaaimbIjiI/3RoLapw883PU7luN6pGTimU7YnChRD
DG9OG3kUcmCPkmzJlHnDeb1VY0I6BRzBx2hvU53S5mXf4mMXs7Jp4Zzb57ykhsxxcoiqp8VzTEVc
06+hmzHQwzLbQnWEUlygCgKrQpq1B7/PNbS31mh1qlhinjL3K4HSwsS/cXoteQKBGSlbkxNUGrzy
R1I+iaL7k4wahKEC3F4sM97rgTERDK4XHE6woBS318FO5+b2aw8aVwEViDdf/P1vUCHWGttNpQfi
oUSs9K8Y3V1hJdvuykcqB9U2qqvkMvYseDeI14KpXkwArMxW2wdEeqHAE1HIKAOsvn6B7swwy9u+
0RXWD8nien9dqCIgPg+DWvwSWqgT72i/EYJmxgr1zBIhjY9ArDyV2jBF4JI8lcuNY82SeZy633uJ
x7nRpXGfU7byWfdxnmYvaeW48vDrrKlntZ+EmE33/GRwaOEA+VEFBq2XpFh9vT5GFygHwfvx8KRH
6lT44KJ07PBxonTw6eGzotAjRkEeFPrDeKJ4JpEZvV3SoVqg+gFbdiILQAd5+80IBh2yXvLhwyrf
UKBzpc/69rHMwXQL8hrVYbLDeZfTkte48gu2Nps+ALd53mcyC7FtzINJdHNqnzm1WzAhWbTAFhQK
xSXRcVhG5puZ8dYh3/eqjeQpWWyqpq66g+Y0qZ4x0V6rQ+P7SrCjy/G2iTdHdBHnM2dvgExzoUxF
c9E4g6SHuDClYSoVnfgTR7rhavVnJDBKuTUA13cGAVPNvdSZeztmUj+Z17gIAMHXSLLi9L2+c2yA
nGSISqDoMCkTxS5tplv29plUof3z6BGw1mi4PK4AKa6tOUW8uIx9eBZSlYZocPt3hQEb/wLAcTKZ
M8Bwq+wiKpRoL3CTacqSXGq/CUTcCIfpbQ1eHImGtlGnEjEGiDr3FR8lTSMapWbXVmCY0V/Bi6iM
QDPBS5I3I9bTDURFWrQy2Y/KD6AymqseTeKsMHdNdpzRIoE8VCh8Ek0pePo6HYS1nJzlm7ltsvHG
nnYJIXcbEYlszCN1ag8OGYVl0njkfxYGOnz9oHeMDqgUOjZs+Z1eodXVlDvf9gcDBmUXJ5GZnwbY
e0unFQlHV6JZ/6LV5QXWd1wmnDYUpO3/7K4U18BZWQDlDqpKxi98HqY2y1AE02PRcAJQ9qOEyzXg
kNZfRtcduTep7f9e6tQ5GsSwK3+qAU4SwkK3P/dyfy7G7aJUol++g+vXcf2PCcdI4nET/N9ZwBgi
Q+OTZqA1eVozdF7Dg60JoxrH5+e6lLRwHcg1oKOd2DHIMMTZ7swKmVNOJrt9Tf1U0rlfm+3Dfb8/
6SwQYPsEiafM7euC5e3eKe0dcc2syGd/rUydqhkMtSs1NWsol/HLKucQqe+BEXCVjLeeG6zKlW0i
xsoEQ712GmSNsdnQOM6TKaBZSl9UxBeA3/QLg8lrvtScKHcU2nd6HvaxZf3Tzg5nCAK12n6vxuVj
g5DgloG92ONgAkzDy5dBD1/H/DWC4Jk/Lvm+uUJ11szaoPdTWAbfm0C4HN9Dnx4J0DNl07j8EBUv
r6lud+85AA17UwKCqrj1/XybwUL+qW4TyMHq99cOVIIsTuKmNNVK40pBXWg56DuBbjmGtJEup2ss
xefRLnKMe0rFvUh6aAA4rTW7myv9fzTZI9E2PPPcm+l08wt8jEyyqNw0TqPFGWOjwCDnEtbaXHJE
Q+ou5QxZYcsCOqtD59YxriRIeKA63nblhXsEAzAkP0S9mrn/PRMv7twBFDDrXh4aKID/ROaxVkc9
zisnX6JnOvWs4NvRiPC/30WaasuZWyeNWPJKuk1oj8mn7haNuc9qvNLfQ6BnLWZMWJObQ5pzCjkn
LxKojxUWmFV0ZIguMrOp1dlcADf1XaNcrnOAGNyBlCvIFu3sO6hH6fV9addMa6Dm/+SEeVJwW0ie
NTAJtS1rjXvvvgYmIqhwSHlFrUBPtLlDGRJQjXqxPr7wLtjLZD7v0111n55LV35kMVFhdrz7Y/sC
iSTpsTegr0deK34xMYvdK4FwMD62s1SSR/mMb3uHnqdrCo6EEYXI14NjgMDaefMqH45bFQ59uxp6
F+n9E/5CBBugecProl7F3dFr7bPM617GfA0eiDiw/akDTh7L0RbvleWx0LFSQ7dBG8kqDQ2HfX7g
bM2oHhoGGj6mtETFT3hItNrifEGRkLIBUvzUzYPhH/lpsCJH1f+Vk5GQ0Knm3YAIaBWJoJsq4V25
5vsED1i3CGOwhC6QOy2Jy8tN0Q+EmmSwh6J/HohCJy1Umo7M5iiK1RXfT3coMrN3onxK1vhxbK3b
JwDNQHftejtDFJilp4J23fGoiC9lyGrRLl6ENpRpq8FY/zpqnw3WsYZwyXwrZhujlWmy/xH5xjRL
ygnX0Gu3cUjypYd6BHAxPTtCGE2mUmEX9i+4BHQNCMLk4S09IyKju0lIaMEVzAJZlealmX3bsAQq
gBrbNlvOZMAjShdaEACWn2PKBXxITzVV7lfVqlqK8mTJ5iFfh8J6BQHKfR7Ao20lPtJBZIyxpBeL
MC0x1sNsJwJuqxMFa5EWDZEJbO6+HU8xZBxUJIOyyvBZyp1ey9dxSoD3W61g66VwaCJ9k8uYmv9I
oPbrk96W9vwvh9P+1lVJlBMLxYqfDXoJ6AQA2h5s7Srp5nMqvjhcPOvdqc8REbTnnR100I7fCxmZ
FLeiiGOkLrrWUpO2z0GrW5waf9HE56oVjStjuhVNlKpHWFI18y7+W6QJm2TV+hDG6g00uD+bcFZZ
70btr3HnV4s5day3AfCtbILeNtHjorsVLmMp/RqKQF8c9rp06NN43O1D/PkXbTAOuvmBsOOGuJMW
DiVLZGe9Xu5tIRVW6efKsR81K6/HgxvZbt6a0WV5jrvzlv/tKk25hPGyyx07d9qeyWCAmuWd/BzB
YK0t0GqgIXUf00AVE5GWP15YaCTmOVgy8giRIS1MfecE3n1zTXbml7/B165qzrUZav+OSi21X+Z9
0Vgzr2w4fMsSKcm8WkzZWRDYst4bYXZDjBrIAZkX9dkOkLSJp70R1WH5XqqaxciiRQ8lw1SYf6jN
JvBAR2Zixsj4jZ3Y8gdWApij0suByvWvYULgoz2EMuZB8tYOnfUh30uhGbcMPZH2b83hp1CQsr8u
n+e6sN1VSxwl+w6GV5cnUXdc0TYd/pFl0rdYU51ZUh2Sz0j8MyP4fFvZe1y/eaxEnnpUXuYw6WW7
OuKN/OGIAK4rI8OOXlAWk8SDxhM6N+NRJTE/06MdU8zoMo8fY3tMk6eMtKaO0+0nRWa9cAWc80fe
J8SVw1zGmevbbAISzrv0m4BZ6SuHUUaGhm/e0kzqe37pklU+wID3kzuKxqYNwhUIW9Zi5vmpIa4Y
vzIHBn8TZ6aBCz/117LScZ4Oad+Z8Ig+XCLRKCwlb0vEHy+42p4gb3R3pbPHbyah9RXtgHP7yalk
Rg466vvwSQlejqXvYxub62np9+8CA8/h2fENxAVQJiMUzWIwkgnbgyUJ2vS+tL3ZJ1JaYd8Pc/kY
ePn8nTmzqJidDebwAMF2xPvhD9RzWAoCX3jvWFIyZxqQtQHxJDlos9F59VftznBkwYDTbu98NYfL
hnAjQjDcHJjH+qiZ8r2x+dXHwoMnfAuj6vqjAh4dIXHYVePt3VY6Ob6RPkcOSHcbiPiuAxnLFCiN
gQMbSOnZIRrmD6KNL+ZoVAAlXCxWDdHfYsTgejGlnYypYtwWVMwNZilRPea9KQQGmR1f+R8fWm5Y
iLtVoDq5UtRHub/BC6IOxiFbGPlTX6kjPyIXudZ7wlaXZYRLKIF1CCCQHo368tiB/aa3HrUURIga
IbzbU8RS597V7BhTl4d/0B+hDN7h1LUa2LDejL/+i25+ll7I4PC5Ct0J8wOFUn1Kv09xWUcN7wuC
V12wfNnGDnhK4tJ0+bQbQk5C/rDLiB2tNu59AyCs9gK5uLdTcUh6Adcgwtg1jWGQKYkQV5Lj7lYd
yDjbWrbUKnfcWaeWfCaeLExbicgSEBKrrLbOLuU38OGp7bqb3SgVa3/WzWtYX15UQHgo1+Cv0fmH
q4F8xhwsOPx0qcoKGvSNVmvgVdn+42x+U8JSep/37MbJpGwQIQPgg4LsOuXDeZO2+xd88n4gDVXe
56srBIZZCghV9grCO9PyWJSxU1PmmNsjemMZXU99NVbNyCN9iGOAesX5S7cAuxwVdJeWug6WXfA0
5gm9tWDFLHt+RGWzxxXdG1Ltt7zAChqf1HGTqqS3COuQYsnQT9fLzVwzAQ8LbhakdBbtkrWa5QKR
6dyPxfFE+PwPiz7waMDtp0btvj5YuZWm0MZk+vbI+iLLybxNOvzwPxrle+0eafHRcoA7VULhaPhv
Dzljz496V3JqEyF7KGuNJzJliPimcttA1IGdUmb67QulhbGDuXRWTTNto3NWY4y9xtoe0mlEN79g
A7rv3sX//1Hu3VvWTYfsASZ01/p40GwhulB9d60he67ONpOxyN9uj2CmyHj3SU7oxY6Js8vi+kxG
k2oHWoIRqldvZJHr63FVuehPmee468/OSmZX3q6BfPRbbVeuJig83nXQfWP1X7i3uFBUwiFjCJI8
cAJuakXKMRD+qAWGWOsFa2Z9CDZjY40tRBW4cOapbEJUmTen1EFaV8XJvQE1ueikTSgJwgCS9llN
iV+YOOZVzU6EufmSsB5tgtJyTOED43yIe05PkjA0XWoBYKCm4AyifYbfsYFjGyw21Kkvmz4ccRp8
ImHy6CC5HfN8kCzTwspxPnoMe8e0lE34zgEYmDPNvAEMlALRccd9lRcM/qBxl10pJ37vrXVTZyFg
weY0+iv3h2Aih9KN578tKbKltgZr0ihXGI9LObjBusZv3vSGRAAYQ6A78DIFC0lvuubKTP37oISa
y9ydCKu4Mkxi3Lc507DFCVRSMjnNgw4am7jnPNRAgvGRZaR2djwAVi0UPb7TiYfPz2ekBlpEJigr
g+4mrYOJwikia8jcnf6n4onTPnbTZbGrAIATif4aktTvk116MhLcOxu8aZXhoIiR7lU45NakL1xi
ZDBHhJsQZZYzc0eHHOGXQZRgvttvO1HHgyLVqq6r+9V1btC9Bn5Dv8UaGX1b7r0R/uNTjuwzW7v6
5lauW7ONVGnSu1MpqbktvHlHYrR6iw/PRGtHfAvgKGZtaVkT36ARuA+i1gDOVXApwXaZUSqEqlHV
O0yfOgDUd1FlA1wmUecnKGtT721JygsCnb87lHyN0QMATPBOECTqNrm7DJ0OUIkh+WwYIocWYu7Z
xCKlIWIZ/o93dEoBjA6eloqHAPRLngz/Zpa1NUpgNQRSd+fgrBih8ElHcw/DAvHHAMVyKMMv4FOU
PHyiq2dYEBTs+/i2DUaFXJoH70j0y02mOAWhwlo24Q8Blqex8QYxY1uZMLYL2aTKXG1L3NcRImFo
5A+TXr27r19byanUqg/tD1I2JpxCXfGfFAjTBs0zor2PPbc1iH42w3bfj25gGaljCK4taJayx9LJ
cpnS8mfqYrn5l76Yz7CXxC3jdGUEVHWEAJeznwKwVYm75stVdK1X/lW2JBgGK/C+dtc7RlOsfqS8
JICLFBQ2WDZRo4wXpedRy6PlxKMi3qDp0nvqGebZDPnLg5C7+TEVKD+Wv1h9uw4+M6U2hGWWr4Io
x+WMQeG3Sacs2pddWy3SxzAzEEYLC91YoRQxKbTLH1+0jkXEcV/+d8YYvU13uUqwubPx6NaUTkJY
nAM/bCD91aKeH/fzxmS7JqdR2x45f+ueZOBNpQWy9VRzlcWG9Q6HlMxVP3szwN5RCHnl6g83zDcz
XQF25CdQPshLumZbxuwUgXX0AN0mjjtchhQR7Pdavzqdgj0qfnr81oNBaIxTMVXoz1RVcmZ3Gvua
/yUwdjLZSgtZoU+uh4eRIJ4Dsu9lL96ZZkQ4xTep/NFO8WIYIjFe0MUJCwg/6/us07oKqos/t59h
Rmb791U9GbacGWfwQ3AGYPw0PoE0ah/+9+W7CLCpowER2Jgf3/85rZs6srbjY54iyxP1JaqyG1G3
IzEzSTyWwy655dFnq7P6RyYnqDlzLnhUYuogwWWLNZUpUvH7pkdWKWfNJhPCsBRyBMjaTTpum5QO
QaDyvOO12DCVWvlADNunb0pKpRgcyQX/WqUTkaXcju9tnGjiDqLqBeOex7K/hfymQfPL2RowXZIl
gtQ9M2aFZGYSfuumlrprI0ZQcXSZaAF7W/Q58OdFJPkWEh0j4AKroA6dTyj5nI25uSTKdWn6ZZTm
BteCIxS8poDM0e22dnXTRSy9Z0VVsKcaeIAokmzX/BQTAh7vZDNsKn9Rop2sZPMzN8RCwiXTSBIq
+Oncf5trpdNuMo2w4JrnTNykkqoxYXpbYidbHKlpiA/vsppDLqmuUwPk5pmaOgbHjPPOevXe7OpT
DXkLgDEq/ZxPitptnfzPaxfQV2V9jtC52jGJiIZ3EqjzXlkFp9igl4UC4ogkog92RJPX5yXcqiAy
OpwG4KYiPqHfzvVXxXat+YmlO+8R32du3jzE9nv6wAHKwHSCLl+KnyWgCUyXaaKlIhRwpAQkPz0J
f5cOVkC0VUzglj161wbqGkZ8gdUcWQFpaS0Lkrg//AZ35X/LjhFo7lA6y2vsRref3chotCL02thK
nXgmsprmhoROW+9XfVvBXn23MobSRO1DWcV1iRzIAhsNtd2SDBd8iEA2ffqBurj7CeCT5xLSOCqQ
h2KxqbCARMXHPdFj0xf22ihhaPRY7GLL0nrCZGbmxyhEw7n1CF3S7L7gq7H2jKgNyN7Rz0KbCs3p
srsnwlW2X5jk35knO4zA7EbcETRldGqlSW92CdpyyljeQBi8ml1pvI9BqXXxD4vYdVO1mcnwwH49
tB0vt+G/nwnwqN3JcYATx5nPw4KW5T9XPQoB3nNNysRniWMfU0v4X0lEscNqf6Rn3iBfgMGff3QL
x3vX8GuUx8UVERo6cjuPCzc/MOtMjR1zlkfFHKltEf6NfZ/AdvovEAffN0yKMERgS2kYvc48Jmfo
Dy9riFVRaBc3CJo4PpefE0n5KO24Ot26sEj+ZSQEKqSDymhfyOf6K1DEAzj0HISD5ppvaIJHGCgB
88tU3cG05GGbul+s1GuIbncaq1T6ixbwBS1lV5g3H4TWX7QOqgxi3sJmX1exv97Hk92uGQPH6G/v
Rn6yfGbtPKXekVZX26u4SMu7PothSEYrAeCSXxYIjTZYfq4bIe617RgTT6fcxiyjxrTnFTNwItrQ
HyaofV2cslSNJYIK+WXEOmkq9/hsMPqagtu/Gr4Km7LGcCOGaLiJzfrlzuZ9gbd+gM5UMqBNmHui
T3pShgWbK+KDWHgGwaMEFAL0vNB/xPsBqqtup9cWjCH/4wbzF9b/VT4t6Sboqu16Ph2FI7fQCfg8
wY03eYIQXsD49Jwkqze3jtIU0o0ZB6OfM4i1XqkOwrctKWmidZKhjALOFCButlz7wpQutLDSQymq
TQmyXKWBiHu3nv03SptLvpmZj6JVgpXxdo/o3T2sSh7Z3ifQrhHDfrOSZvAOtR6jJSBnLt59q+AB
s12hrPsDQXOChUlg9uTZrKQWJ7P62F2x1YSz1PWBz4T7KpswxuPM/N90BL3ox9cQO1Hfytk5tHBZ
zOGx89+FMxod7TKcsG1pqyFnDGTZmm9q2mMCQAIqpZ/SHCJSyKTbyOQr8yed5C/YwQU9w4DeVS92
Zpvbm5jbvTAAUtoqdiiuXLi0wx8ZbWb+iCRl+DggKoODl7HSeR8PansKBTHPIjd0GWStTsD+vOsL
+GskeHRk3R8DklJOfHHGLB2YqqKaVkD4ebjkNOHX4dt984tLJtZgZkqK4vBN7K0r049Pdhhl1Niw
8cXLJWVKAyEw/006BKlL9BnkZEq9Ick8u3SaEdz1B3QrvfThqpAHRBXyCGemp/1MvsrQnuwdwRBj
fDOvsV8pmViCIx3nxqYswHeIvSsORG/vXZsAv5lRThLgxUep/zkjkvQikU0B+8dzoiciQpWZnAmS
87rIqnq787aS3Fr2ex2CKX2+NMgoQ7vjlnGLGuMAap7N3R/fCXodULpVlDxIyYwt/ctpaovP482I
AMLLv5ZagRPnZZrplkrhM07TDbN+17wNJgdotk28qBjVXrCOZhKPHUtvJ1ODDv2coUChFQd2nipO
JnD7fM23YfRP8DCGF8ZOxuwMZDylaEfxlXqeCDI0FHKwvzqxXZnRsptb2c58AzSFEVEJ3tYufNFq
NFUFM1s7eZrKCOkVImrXMusvce1qYpbU9bzahSij5SKvVu6IDZ+pPSo3c9UUfRvMYinqZ62xV/N3
sBj9vqJdKtIJSNxufAbhIbxjcAUMnIQMzm7OdlF0MRHJtdxFKbaBVaQYy9nzYHXsKG1mLq8U0SQ5
PCXG37VSs9tMmsMctuvgQfCdYQ7sXaRnTLULLLZ7wRZ/LTQraUb1lTxT8ibappoBM5pnDAxLlQOm
hwr8Zt3sGusqXPhDYIy9qpqxD76Xx/K8X9t5teOtUaR2i3R65fHxccX1okCjKwwbSE3s0Up3MMGD
DjiqvTPsv6rMDJHuZaqBN6k1wt2q8E7s8rKokA5y/NY2HpYJhjzi5Zh7fLJyFih7A8r+I5uFwF3a
mgqOFP9UThKsxFkjC3zsUeDtd7K7WYii1Dixxhf6wFPXjOGGtvq4X47CaVx+WMDzPOBvJA51C3qZ
Ag3VbdPmW2pQ/+cb4jDR/WNjwYE9DNGhJH5XJTjpTOnAYnfN1aa5qWf0bUlWK/gvtY/VJKJH6Loh
vYQETzeFWOnQdbAaYrXETlKQ0/GjEVXotnFA6yxoWKBRsO1nigioN08zCh5S55173NoVLxuzaFsz
CmDY8hvrW7KAbqFzKnHrxOIth0hDh6xSMSK2105GKJpgMY4uavylKzgD5+Oeolx2tc1lg5IsRnXu
hnlhdcSbjYVhQPfA+N/sIk2wAbZSy+nIF8NvTG+N6vOGG9paRUisW5Q3dVTCny8YbkGQY0Jpsz2B
6/NU0jxhtREk1uZbhIaS2LNvnYwPOAB6JwXhUSyxTNwoiGjKWsDVFDUrD8X1Wx/9HbdHz/rBOf2r
m73y5dUpR6PTh4zTOSl2TFbXFjQ5D0rWt5HyEXLWGjTyL25tk2VAg+/j9yV8meO+cbeye5TcXlPi
/co2j/t4b1oIwdInVEe6XZdYnLt7WKLJFbdVtdWNnDRjDEOLEzNII+5Nrrh8H3b0q0oPKeOC1atm
RggMxA70eALWDIMTvufVtOGJBYMwNioqkDTNMfC4MGXyyRyBW0/htnJAFT62kiGJ9T4plkpT//b+
bYVSZYC1XwyDb+3bFr8O+DdlzF3SVjW2iw3eLult+Zdm+GGi9zp5donSYAUQVV2iTU9L5Ebpv9+Y
aPn+ZurPNzB8qGB/SiXBOcTXL8UC1tfg/CjAFOHZ+L3Vs66kT23kGYgbVtshnSVVhqlw2U/BFEPt
Rfk4yAjnSHm/iaQn9oesNaWfsqb524d8nG4eClB06ThqaO9R0LLSaVKzszYDYLM/zibDEYj+Y8vj
7QDznqqBaJasyaOdGDlgHjnmY+52lJoBuRy/YyBeSUS6xNXubvr8gPgHWwGfV3tqTcSJ6JrRkm7z
mPt3jkSy0SdrS5LcsqaWI9nPQQmt/dAS7tzxP05exHBJlhoKt3Bmof22UiBwEM8RZJcTMBKlNqkj
0aWoQNIv2y/duddz0kUDQPFpmzJwo6OHBZYqonuhKk+2if11RjnmnGMlw1AM8QVNgig/rzkrfLDC
R8cmXHuTI4Nte3pyJkJyL8cdnJemaqAnGsT3mmIsxGwa9E4LdhFP/8P5YQpUT59J/l7IgVCIdp8A
nko2VnPsEJfbgGlI36L/SxGRQZTKlBaEbEXXgSchjDcLXMyk/ZWiPnTV34nokC1I2zo5T7CXKtUa
CoDE+XYMP2DnaWGrGjLVXHzP0Qjt2SEVC/t2WppDsNkdeiqrAid3b676DTJQTTMN6J8Euig4EDbm
Sw9AWtQdV+WXJgu7p1QEe9Iic5rphfp9+B0vI3/C4H2wNISycCW3P8675WBhsTblKtQ29IekxD18
kQ1HqCbLCzUlpfpFgDNgm7lMuc82avWjSuwN0FZ/uMAEidrxT5mfZeOA7lLyzCqWtXcF/K3mDUSB
q8ZWW/RJX/XTReFQ/IiWaCM3BXv1W/SebtaVpSAFSIUaey7PD/Avbtnj6AX+mqsBFepIiIQ1mpSE
2S3eV1f8AFmyvj8+QtU8cf7d8oSQ53QV7AY8HkQNyTJ6hIX7kI+hcsYKLRgKFaN8Eg4NX6DIXDvW
w1MSUZSIr2rybP6KSqxEUP4DA1kAkbW/xzl0E0zJVfW4zL6rLhOnUEBOHAEQGjYnvJvNydNs5V+L
+Fsi1Q0sPBxqbvoNikp6+1exn88ySGcuC3priyHMS6K3a9SFHW+NIloX18SsrqfDWnJWf5qjE5Of
djjeby/GVYLRCXWfghf/TMGByf5XM7t/7Cs/+snCxkS+sdUtrjtwa6PRdYpfK7HRklFAA5P7r2Kl
ZzIvN8Lyg6kEzT+6ot/lFO8qR29Uiij3eHfPX4Wavw9RFi2TcmHIcwV6VSGGXnopQ6yvem6N44OC
EOjxhiz3S3mCVbd8B6ITjGCMz5hHb3PA0VjHQI1b2kfzGccFIQLUwf5DnzO1rFO4Tc9IfrUcJ0vR
lj79WehhWaM0lAvywlKvZGyK9RcKpElGy7Tlqo022aiFy1REMWBk5HjP+j/1rH+4BwZ4EyO3UVtR
oRTEJ2PqWDWbwUQ5nsdbI2ScDmRXXS+vgR7BfgMm8A3E0Sf4jHWPeppgp1U2Xwo4j5Ta3Zzvfp+/
hw0Ft7dc/W77YhXVEIQlxaLKjmoLUJzjgDJaqQgeb1APotzi+T/+NGF+Z47VT1ILcy19JYD2HuJE
y/x1q3UXrVXqeI59ZIXi+S3G54IiWA1NHyBv2r2M/khxuuMXjsbpr42emrGlunYWSzasZcq8chlN
uTcKFUAu6NumIXkVzecQKRHPk18CMlo9cVj2RNeWwi7hyoiW32Op7mjI0JEUDf/l33hPFZNgZtfW
ZVpByxviaJkaNRxVARZmwtU4yqHS5DKdfIG/1XnJzMzqo6fGAgxkViUd9CP14AuIDevQi/uS0P6a
Jy3wAEeMEj0jqMK3wkNeQk2+6pISlklFO2pNAA0Whyr2RIPQRtyUUtIUdDuSE5G7ehDLKDlbmCpO
3qLsZ8D9nY+Cboi+6BQkhjtw0zsZEup4HM8PIorZeY6ic3Zf/EEk0PpyV3mrIKCIpy+VOqtxYfTe
n/x0xtaQH0Yz4ilJmRPGFQFgXNfLiS96Jkwa6hlLkGJySHObqAOpJg7JvKvffj/lME/WHs2jNFVH
NcmfTIvHAvls3vuRlZif+nmI033blyDVkgs9pJTsdNI3l2QS3MrfruTgk1XzmV9or3+szgsanoQ3
O4S8XVWQ9x9SOjuTIASO/RT4vQtLZftTzXx71G5g6R+om1KKp+Jux/PWOXP7xUHUcPPbI7rxN5rM
BHLs23rhObyueQCJJfGa9t8/GgHb3z8CREYYk4fWVARDnXZCsDSvB5Z8MibObVHVWCFlqno1JP3A
z7UYgZw8rCYUh6yCJpvLrMAPy3lcdMfUE5QPyNnC/SkWYDKzgISe3FugNYiuFoGXuqAqcwa6c0vV
OhJ4BUdxWdvnsMjncLiJkl0NLZeZuDrKf6YDAU6IPb+tcVG+z445aIiWBHQYq/nMUhNCJt8ayLzj
14EEE/QipBaHY0oJh8SIcXls8RcfVOwxbpkHOorwkvTrXbqHUMt+wGcFhNdwyDKY8TXZW0MGAC7/
0Jii55To1Jjd9d8cNYvtsS6GHZUPqv4u8zrMHnsC66dLj4cUeq5FYcOEbRZmfPX5swJKJgutvkRP
dynQao3PSwWbiz7GFmRWCVKU0tQwnGq7vGZ88OWmSuWjlz7XE8HsVawMnHmvBDY8+2CUuH/Vh3FR
I7yx7bb8cRnWpRwqLc4u9GtGMHgCJOPrNPclzoRijX6A3ta9/0ud2pszXu3ntmwdqhQPoTNXstfz
yfE7A/MHntj35iD1Y+l/gzubgq8vugb5rcrh3fLq49fkBzA5XYALEmOG5KzLl7KQVGEoRYv7yPIp
Yj2SJVMvCPv/ebfiSLrzSCtSgiqYHgzxWnaMRESVgpOar5vAD7KRQn4jXchF0PMfHBW0tOiyhR7o
nkc5X9MGmho0TdzJqN+zu/9+n0QJXTd1MZRdBrpwFc+LFssATgTeyS8a7hE+TFBEW11I6/GO6z2R
rkhlGigwVswDBI8Bwhyi9m9UDqbpEj0NoKO/FD488jZCm9BTl3kMVmSY78ELwSAGAAXa+YOPV9QD
GrSG9PR7ZxotKhaiThaYJvSz9VlKtJ2idTa5yliDhcHg3RLV87kZdCUyodN509C992RygKe6OuZM
5zU4KM/xqMO3CXv8uO3z31szwPGDeL0wYzp/d+Y60dNCOHZEtZotDP67n5K6EVx2FzwUcnyxhMSB
oxJAoQu5h9SpAVp4K8/lLxG0WFW0aavqbhqZlqiXCK91uFYwvq20KATk45TZG+E7FUJDqYfNhy8+
YPE62TBwhYgI2DdQrIhQK1dImj/UX6KUiP6UVAE/vdd5vJohlW9Vkc7r+B1ZzaHwvnV0YtHKqyEG
QELx9ORGknJSm6JLfQSjpRplEz0ELVw7dFFbQ157k5Nlcxk83wp0z37KjMHI8RuOYN+VC/PUeJBN
oLUykEyI9+FxTkbNjG2cBxXnJcTh0YkYwyNFG72Df9PKrFZEV6MrCPw2g+bPDOI4JfgZ3REL0crL
kKCJun5EyDFFbEeWUlsL770GJDSBfcqSV1CzMfmIwfoV7fhE3GJC6nUcojDK0fp7AbrwjQ5ailGG
a4R1Gm1/LkgaJKsQ62WW6F84hHU7FC99P4beXv0X0QKC8bhkQxZeZm68ZN+862Fukohtk6Z/7Ye9
zL+u0EaWIcP8l+5aqFRCmhTb1xoCQyTbvT+lFmatyu2ym0+ey68l6keULjafyRZPHeJvUdYJNJKK
FJUpGOL+FrTjCddfDuFOUcmO3mVLUqkJqFpz4MzkSoAGLaG/MnZMWaCtFOrKt+eDDnghybTebYFQ
50QjvmtkCCwhFBYopPVcfh9eip6PAVzf/9TYZiOPgK/YCnYdLxPKLiK0JPXizjoh8nnDZJ4wkv0Y
kGerIBlhKknBW3wpBnLmKaASl9z0w3u0XecgEuzRwKv1fB4yregaGa59Y47TWPEVn7soUkog+AOr
FX1NMgXUQ627hm5Y443N638sat86qYhByf+6KSfvIXZFPJHxm5ysKMgEsxnPpy/KGsmATKTFSJfi
D+1d9WV6nJrmnu+k9ve/cxdIfAa86bsiIG9zjqKHJjUiskbrXMLccH0AoLbZ5a3DyuOZ7vqFt7ow
MD/e+xjxOFimz8YAp+wqgPci+Jgm1vCrNgpT6tlOzkEl6RoCTh2AV1N8Q726LDpE5RIzAdWAJbmk
NhAga8kLaFGebhVJD5DVi18ugPgrH+vwogkT15DX2q39jrDE/Fnr2ccVIyWLo7TuyRf2vFZwaIT7
2CCVMLxo2ehaQa1xbPyLlTl5VU/N1/dC0SYgNwwbOqdEuClihwkp9KllRHsHHS0CYuTLNMHINPCy
IV0QNkBuHCkZQFBvHrZIyO8jHiLmvjGLAB0tltoswk0mclIUGUeW5abTycR6r6Qhy2bmwyESsJ1n
/V+HAR3tX0INF3snRTJ5qvXWeCLjVTFvB3RiT4BJvU6UXd1neQNRGKtGU4UNQdjbydZtU96H9wsr
+hMsNKuekv1JzG7SDr4HAthyttfZ+WR86d11cTOgPv/C93fFEx4JPTLKmaNRaoZNHCGuPOuMVLXi
2Z6t6vDvUu0Deu3lHm4VMbfn8nSMZuDm2RyUxJ7PvmjkywcbC4MOv1RwYh6OxIzOnJK5adjtm8k4
piEqMc42HkQl4QV5u9Z5UZaPYiZErslsJ4ifh044/LZ4Pp+iH/OLhWtzUHmjcU6UqZH60NYzutoN
9677YNvQAC2RmCSmSSLuyxZUBlnoVfupbMIewcwA7C3xBboH+IR9ZgHlBp3rGbUsQCCdn5pRboTY
9CWiXqmu6hbtekfA6dUHbr2QE1xLS/O6qPUBU8fq95PbYZg369v/qJxpfrqehnAWhhRGn9q41fm7
0Qb05TFAjzzsTtNJOtnNj0wkrlotTxIsgm5vbjeQHJ5BG/n2Cnbnqx1Bc+paB0TbBvDrjwXyQdwF
1dLDPQ2UQ6k4BUCme48K83S4DxtDoWX4Ysaxvm0R3chlR2f2fIBaTdHzDbP7K6JVtWwOwgLnYxxU
FiFp46yh5AYRTPeLbVAZbaAGf63i8MUhpgL2mWsBmVxPxlIU8PpYbW5vxBTzGaJiTk9OhUmkwDpv
9tRuy7mDTtiQbyuHIN+6i+hkJhO3urJ5W4xeMxdHq+/MC2lM5sNCBJktdtVYnLUi38tyKsEfig7q
8Rv7aZNou6mSMlQxWP2d8Q4gWG4poqeLou1EPw4oSp6fv3cIyStJzBo03SuoqI6vphpBsPy3NEMT
M27ifoT/Y8oXN8ElMAu7nZuH0DzDtjropgz2ZCA04dQHghJp9/270aoPpx24LXmk9lKMONUviZ3h
UWV54b2AOEW26Sj0JuEwQVgNJeycsmRX8mq24ecYpObooeVAXyYx+YKWoBW6ncnD9ayGGOE4swNK
GuP9yoIVhxoPOWnvxuiDNyepNAHECaP3SMIg9KuKXWKzycpBqFKG/GR5BHkVEW0gyWKbM1bSpR1f
ItHXilpSoRXDTF7mIlySoqNlYKZcIr3Stv9SR4VwymEn8bqlx74vuBNxsKeGPFRFeiE5CuUbDxJ4
1CaWJyIbh7l1Fz51uUgUeCskVu3JN3NH+Q2dZzF9j5DLLMgNSJQ41ZY685Vg+z8Uo+zP/EQcnMt2
vkMHsmGpJTHD5RtmpJzDqV8ufQ3ATm9ydWalp6Wjt4xuWS3gm3W2GTQpFE6D2yZIT+7JuFUaUV/R
L4slIYEOlTaPq0Q7eWLRsqxSF9jzbQ+i148nYRa+jxxjTXXxa8tkUX3OH9T2MNSTBkC9SIDlW69W
OnFOLzUs0UARZ7VVzDV3aX3hbkI5v3Vw8lf1PZ54Hxr/LCOewskLsZZVRpo0538CSKpKrEyN9LrC
VQjZVvN76PDS+L7ET+VmbBgbjEcSC5BosXtKi529LHc0bE4wkDxYhRT4DrE94mURXMluylT4Drcd
YZ9dxjt0N6KsLk32v8ZMIYe6HEmozkpt5sq2ZJxfxLH6mec8L4sgcn0K5oRVRbHUtwqP82RJaz/S
ehcRHcDKbn1WzWfDyEZBif5cwavx83pLg/8zITMSOmMbOL3Jwed14f6qflPMXYeZUJ2HnmNR1OIx
gIFSqaof8vu/Ex8a85EBG6vKPyL4yzqMxoiVo0SXVYNFCXLCEADrPBcBAUvWS/wBJC6cI/4D6Vu8
zfN+6MIHena7EHH79sGkhxwupW/5cLp6wTlZucqUdTw4eiK1nK9fuaLx/mJycQ6yiFSemOIoYZsQ
QijNx5qd0fXwgfWSrdU/Y58W1sm7joxpRZCDB6ggwkLuFAqlD5dLzYubx/p3OMcJ5Es/2rKvd+xA
o44mG5BuBRXAffdM4FiU0p1M/EMVr/5sHLDMn62QyorJaSrsoTcTHgtCVbFQF7QuSZ2Rh1IwZ4JB
q89JFNBH8oPT4JSrG6tgxBRAKqG5yHmHV2/K9P1CxAFK6m/G+M73O93Tw6dl26RUpKDAuIPBIdky
GY1dyavJ7VVwbUYk7Gc9Z2L78u+ZvWw06ghk7O1i632gbRdU/2PFLkrdyHLAcTGSmZSpP0/FmBkz
SVLYGxII61jb/fJIylGK8cqZD+5bjdXaqduZbuGRhwbt6EZ7U0DfC1crEylXX7E+EOf1kR7mDFdm
/b9TwX57VQkuXS13oebk3p66jNDOAvpKD1AqhsbgbNA3GPhUSR8kJbbmaW+sg+IJBPfzncrUbRvx
n0Tu3WZ7qfAN45t1PNBBufkwXnHZmzlwaDPiS2HW2YyPUJ/ypZglOtyanoHR3FZ71lSS38485tQ4
sz9uWA36etvYv10WjfwwjGMoTN3dCGBZ6xEDw39XFLa3GFYhM13FxRb4hnpdO4Tq4maQrOex5/Ge
91sVtpaQdnqF9IIqXIbc7xIT2KrNf7rcAkbpP7dtTIvKRyj1o1YOG0n/2SpW94RK8CL5lKX0buyl
CcWq8sF3BhM9VhZjjX0E/qX93h20W/ck7nenA3dj2IjddqXTThUk6foH94BiD13e9hJ/32kmc7kI
bBuM/ZiEL6mjDUii4H2AiT1ry0oqQPSyRKSHBVWRkKqAMHTaASBo5PFSUX6cG8atKXLwKOuyJ9RZ
pZbali+jLF9Gl9gHsECYTpTYSYx0hLgnuIw6mmkF4RY+v16kc7H7J0t/X67VqOE8DaXEqQ4iddGU
6eUj+lRAp8PqGS9ST0fCm2KQE3h950q/MnEj+wHkaryrfPrj/9kaGtT+Q2uCUTpWJtyhHguy0KVD
fVwJkBRFKnF5rIYebfGvJdaVk93P5klppj9f3X39KqZ0qNzs67LJKpGYsPWuQQ5oSMD6cQIWlMNd
yd9KoeTkw17Ci0KCiRtV78HvzOqefEs8F/kc9rJpLdyZ6/Qu61efmgBgYZ7raX5249of0h4UrWBi
iUGvtbLV+52vDyK4FOWn/4yALyVE/6k90KO8gK4JB52/orfB93Vg7wMdwpqsnodQG1m+ii+2WcA9
sRjcu3iBPIWDpKk8/TwVxYWe5hBpwdHtGBh+jgwAs8dDr1UCCO5aaLp8d+2JBk5+Dtu1mAyl4+m5
bKyDMKQvDM90Eawt5OGp3MASvv9W7Mb3osoLXVsSwiRgN6T/7jNL62k4S+o/CqIP9HA15x43u9oP
/QR1wPdUzXH4FLI9U/f6QNhEUdLSHEf0ymnkGzxgONlQjSIaNvGa6EcM+XpjE40DXi1jPpB3MnWm
aMsFdzOn/pxYSqCbln5aCmVve/rcnvJSANcNW/6TgBDQbDmHci8a5J60zSXiWtA3WF1zM/a5Lcrc
aDUV3sofKI/3hLkoO7CNrWNEzXxTB4G2+rZ871LB3PxJGdF4C5lcDwTMlC/HQhLUhHsXGEiVsiz/
4N5rcs1fBt8rjl2PWRy/K8/xgD+lVq+t/V0p9EFLC9h9s9WKIyeyV4Vsomz3oarAqXXBEwwb62cW
rxWMfU47PPwgSuDQzLZOVfFMpmqs+MoMKjdh6HPRIYElJDdH7EgZS659aVatiGnhGLX2Os0Xlieb
F0k2U7ZLHHpBJDDjp4mIrRNER60/UhlBO2wjrXPHuO9cqVSBh0HkMKswD4megcKfcOMarASh75KX
bqPywzhBYhJTIG52Yr+xhBJ7JbFuEP5VYLizWQtbrY0OWs7KGIpyVAkAYUi5p/nCWHSejg63hX6+
2uMEjK+pPqg6TZQfd9mLj+UBWvwFoV+S6jusMWMFRJGF4/4XBPTEtq/pEOveVIXOQtfLS0mc/ikO
aOj3xDOqO53Lyw76PE+OEhHiQV+pTDbr2EQKLRlTS0eEC9VmWjWQvMhlB0v7KSjye0sqmj7+xwMe
4loagkMOVCdBuH3BC4OOGktDJ8A+AIV+iCm8EreYwg2pbJF6Cibxz4qwE1TliG9yXcvvBkqHxs+s
Q86r9lmDtqf1uvKGi7KI/Oh2XaYouNTYwFezcR3pRKoqSO+/fU0jFVxS5yf53PnvbMJl4kS9TH6e
rhBBbr9/fg8cXXmkoaS96f3qPXccjuwzVWU6XdsBZPE41keExf0zZYbmELc+vpIjwSvRy16uQfr/
NwpKJr7Y9a1G5JRrpHsNLmFHlreA19IisvbYOSptBNa3nzg7ZaKb3abZMPXqKk0twuvDwowb5qHx
PFa/HHAu2BYw2egk/lXimAPkpgqd+AawA8FbHJ1LPaCbUT1N0xUkQNngKiARenW9Kt1J2DaINorj
k7Ird/Ngq28KaXmuwnI1AuT9qyoooL5C7pQw6dhUTab+6/67CcwPbGW50zIQM3EZguW1zbNrgEDe
YOl7XMNANnWwPFmbdLVGUN02lZHYSrqdXWx7BUEiMEWuFHbkIXkLTMwnGDIBlZDFL4UiOYVpd73V
SHYIN14NZj4UqIO33MHxEkzfsTVe6zksqPKTqafMVw3n+io3QFoiaM0b1YxhvTok0NQrG/Y6bw5G
spc5Rj3SBdnntPKBqEdVU/gAOzU1CVrf6pGYPyWn62Gek6bKLdvtAQ73lYxUAUBTTil7W9l/bWtl
GrG4tvpdwuezB1Po+JTrpz6d7QckgpvIYYCiCsRR9F/ix1PnUFafcxVil1Wmf7rJFBB9Y0VRTEcO
7IcpQeWyQNThzCRUNy+S8nsf7XpLXPDDiJWLysOysNIOaWuLtwYsc6gHSkFug2CWw7yq7YCO8o0l
dllCVHvCbUOTa1UMB6dIInxsSDip5fjzw2dg+9HyUf5No1V43YpuT/spr8MOXRvjmxEhZhYC+nJ3
CeYjQD7o24aYY4Iodf/KY7DbotwkOtgDstCULcf+ohABmd99OXJBcfzP6pS4lluTOkueGB7pYVPr
0+ZwmzoeLosry6A+FADaaBiEj9UmWkC78JnGYTg+6gSJ8a3SuuNGACxLa5zApwI6JFlUz1e31jyx
RlbLNsfv5R0OMDiN6AXPoVvLcQPbEX0kBVoBtaGxWn7ygUSHo9m5zpyg+6Guu5ia00UZ0SmSfcuT
fNqfP39+rxXKH4Veck27hX87MtDhDVNyy2p+RIM04LoA6TOUy28Or6knktdpQFODn/qa1nSx4PuZ
J57abf6OtuWBeUKbKwLTtOSGfWqPx9nRsxJVQVEVzANFjHcTHBtpD4WMyAHwAHoD0IIgmX97tzvR
zrBrmBycAXLEIWxC458BHkg6XdRZrtIBT4trs0RRI0jWatrvNY3J/jSyRGOFaUK0z0JMcAFS/M6E
4CxMVrWqs4L5Q4XNiQ2R59cdxpeLFL64oNSUUAoH1jTKr9dYerRpv8wXGH8sB28/6rEUsf4NHS2E
/YKBk7PN06cQQ0UoGS0tfCg00e1bsTJYsKOxlePdeDgAy7Uku3um/5eOmDlMEwmNNVxVHdNC5lNq
jLQOMzaEDh5Kyfye8rOC+VUXXvk0OMz0aMbxvqcQfQU6QmojuSMjAu1IDJ+Z/5RWdsM1lW1tu2Aj
c9ydcFRYUdUQZYu/zABKkfuysMNYmzo/FwjuNLgHlzGWmunWUsOktXbhVqiD/kclG62I/rZyNmF1
yOBhn7zQ0FyZfCJ5dVURC0H0vzmQmieOIaK1UDIaYv6IBTbhr16iKS79W6mIDUYjNbN2zKiBdXz4
lj5u+yTZ9Ea9bqWk0xa8LXrifWU5yxaVIl42E/Mh07tI6wP5aSpY3tBzBkNDvHlBJXXR1bPQACfo
4zumEqLILel+t5Dy4HxI8UwdbYKcVEKewLtIBo4daXT28HbKgbJprBGpAA3RMdNfoa6HBx4slg7e
V9EW8rjBR0rl+Oln+rCFt9D58nyWjP9MOsvFyPRaAK24O8WfRBEHs6kbCVAst2MTjl7vqRfSU8GM
giCZanZcifymdgBZbgOZIwfp2uD32jpRryPn8eY0m9H8nvf+DvCfG05jDj4hOjQY/ixo2UZ+naZR
sDvfQ5jzU7JqHWd73ogxf2/OVi7vEIHEQ1NNEE6ALSdZzD5h+9q2M/a3+dz/i1K36KnsMr4mAI4z
hdabdjr8YdfiI7YmpuwfUmbH54FeKVDvkiuYDPkNyQ4YZBMvv9iDGaEGYCKAeuXySRzvdC7LO14c
fEzL34wna1xjobdprUtQtlnr6K0s6CMKVBsn1E9624IeWtBYgEk47Kaw7Q2wBoMPPqMRqi0qetQc
O6p2dtV7j4GrmeYK9FTiBd9egPijBVOWQs0khbzm3UzfZRdtc3bx0+lm8SkPfPf601LL2IkSgq46
y8hLtfS/N1gAGkmiCkLJJQ2B59NDMPfEGpk0gIAqJmZ+zfvpX2USc68YMULqkuEcqxb0Er7dO0z8
dQO72l1NrAlPUA+r5gwsx3SpXnAidh3UwnZ/duxt1tGCQWiOLfc6QSHlIElfpcGVeHKuGmLF2JBz
XMokbL25uchLBqXZgjiVQjvpWthRIHS9wSiQ5v11HR5oZqhux4Ts6hmzGawATqTR9Sfp0xGY8uot
3qJc30o0kJfXikMEIXriyPq2ehWPeUW9dLT81w6LfYYhQclXLr9ew695VbfzHMOKKbPxGV+Dv30y
qasIv0y1W8T1jUUixNetFI2zIyCf5QOPd81K/8N+17NMVUQoTB7zIhilLR5WA3KqPZ10vEaSRdbA
/fe/IAxIBQDV/dn35ypfTX7A+AWWZdqbRFLe7MlwVu7/yOTMln0pNoMZ+lh2IdfMOGWS3BhptHa6
qk9rpRILyDxlNFG2WK8guqlOY/EnOrJR7F43sr/eJq06w+u5I0aFipDkfH8sIuXJM9WzDvk/BTHh
QU1X+dclXZFpCmG7HzJNDy2YWjwNcKQdnB/ORl7czlGxnYbPG2c9vPNQ9O6FR8lW0oc5PsNW16z2
eDYyZTxd83PQrKT+6In8Z/Rju8t7E3eYXdsoE98tziX33jcK7Sj4fBjn2m64tGcmj9pKvh55Ps7O
a/xSXN42mSQutyS9Rh+TI9m5dq7rXoXzgFW2pzACWwntSTvUqLvZE7kdq2tJZ63izHVldqn5GGx4
vGFlxrRjjB8dzcvGUMS90B+ZxB6V03FSFGD52cLgnxfwj8HG6Z0g8GrN4Oh/RUPhBMLJbv5uJYlP
Ke1LlfSOhRVOuts5agEY+rf+O1Q2A3rglWB8c6ob4C8ee+snNK2qmoSyS5nfR1xv3VNMN4WHAHal
X1+C3rG/F/2aa50GOUhXdtR/nWThk84g4xINtZrf1O9pkJXHCLkbH9BgG+HL4yF2JvWxLtwiAuiH
eCB1+Pz0VrRrXN2ioDpmJiBWWvszMyqypjGNvhrQTKRHmnJWSJTqC+4qlJmPhRDCIyvrcHUho833
G0yzFLU+Kf7OzOLQAke2yXSZ26UdU68OGQ5yuyQCK1AG4m6K9yMggXTviHPWrXmjgJTihQgZ/8xN
PcVZwGOuA7KnSQJFmxYnOD2Q9Z6yiSnPJXv+Htcd1SnrNHerH+wTubC9UT4LbtbxmxDjPdCO5T7p
C6O/+YdXtXEaUGJQ6X0dN+DIBSz/Hv3OztrU3c/c6GNfu9m3Ij/o8LZ8vsZjaYNfbdGIrwaTXrgB
i7su3kb1yeCoAuSkaXnq4Tzwqu0h6tyComRIKQt43YGE8AZkMyOopdBTkFcI3TKr7xyAB24UCgMA
f7GRCHU+33FSl9N0GeECbxE/8GoWzkr7Bmw1NoYOqoUc00yGrf7B8bWqavsBWWEM6UBRWUMhzNQa
Ru61LZdBlcq8MMyK62DmYJCGuEK3M74xFafmTLH9LpBeokjhTHcqMzbvUSMt9RNcKoftBtvW/eBz
7EuTIDZcejH2hqN2HJpC9k8unFdBNVULykskYYg3t6ZZeec5XANZmIUEUJmjxZUE4DaH5sI+s1od
BKBaoQlNZYFV6y7tPMXX0IGhQSBRtk3dR9bna+m9xLFgF3KSeoKFna+S71+LxjrUaPnWZOOITL3K
jvzPIWPAgRV6hUnnmgUZgSVJ0rrj5wcKAVzGvNwpjnKA2l3rnT/6lKgzEjdv8/JCIUtY0pxsszuC
8BFmXkZxA1pf6c9kQTYvGLLYW4RFqLFq6tSkRPwOdkBeRXKln3yU3TmEdOzektgZIDyX/VZS+H9P
SDzEkVo80OnsasSbIRxFUds8FA1fz39sUZBtEBFiVahZJ1n6omMiLQASKvBCn/4cFywm8U5AZyF+
PHD1IqXjX0dpQAJX23lB9CHQnA4LUF7NwUiqJY8lWUL9eB2x9Qprq4Pu+Gdy5nkNE5VNZCYhTSMR
cQf/7aRvinZXaak74j6nS9DtbG3j7oVdM52aTUXCj3/3zvsvol7lNFoP8E3H7qXAlOsq2sC7wso0
oMLhJ5qAoLJnS0iIkn1GfYqhveTXIT8MsZO8n0uA15lrv3ksM5i3hOlBItzqwZZ6OxoEvuJxK1IO
wkd84pUIv2TWC6nxziEY3igK3hG8qqXBIX+wNN/dOQv3tDssF9N/73s2hxm2+nA4ehfSiq6/cgcP
nBXHxtCbEi0bY3tgVCf3gablJxmkjwdPT7QrK3iwqhngQUpnzV9FqJegBz39gn+/E6g8OmVgNwYF
GRNv05UwyqobLb/dontT/gQJEFau63k+JvYukGtOk5DvfEQxxDP2G2uMQlFh8mZeMUXy+KIfrI8r
KggDTJ2jMiEv2wqaxktwufWMjFDGqx5RkS2IDsvZKEelXOFZ3UTiVyUkqD+ZhcCYnaVLlpMstUvB
omJEi9Ln9vONm+Zp36xtyh/lSdXRM/348RE9ZT1Otm+SkTs8VARf8My0TSaNC2H1v1lJvqnILm7B
FJUvX0jBuKVcK1gOIMYv74AoZv0kymenIU13Xb48irDOxklWtGQmQyqJQ/yR8EJstSlWC/hdlGEm
8rbTOxBn4VhbMt36p/M6d/g3nsXlsebtqFWSa2/lfbE6OejvyjamvPz2UOlc77WDJt7vntRyFBSO
TVEZvy2nnLfzHzak5wuMwSC3F5O52Tj8Pk0M1AQ941sRTQn2z5iwjJSHQlA/mpBSFiHfQ9ON33m0
/hv9o7yROuokN7LelhtKTkb0jhGIyrrAVAgnwyH3Len70EeADeszM30zIQ95f+jjN7PCNL6xusq4
5dvfkF8C2YWMk+QAjPt+JbC2vDvaGDlaHjPiNiTfwxCAYRsBECoK5pr6D/NN7u63ym99ITtdjrw4
HmLB19dcvyJLZnv/d8JEOzrMalssQGRv9KkbSDSfp+6L/c8Qc1/8fAIxgFeaNMz+1YsaEGtuTNkg
l6MJmvRaMWxbs9dtab3KjDtY1zFz2w6PoOoAsulq6u7TMXFNjSwQgb8cDNEvTM+apKnQ+WsMiJFk
jUcrTDZOGRXkm/YWiruKjOHv7XNrQWgfk0prDMLKUOoVbWDdCI3I1A/XWGCoj4HiUrwnUHGV5DtH
RVQa0a+4e5C+mAa8xQWM8STK+RGYX3QbycT9+4Ho8UFgqsnJjJRlQPMOd+2kf9UWMfW7U9M9ahuH
dU82gmwp6+ZlGQBkHCMKmiamxE0zPmQVgZAJqCQxqx9UagWf+EkEb/xqqqowAI+aLc6KuXAz3Sb+
8fAKWoieWxordqabd3KavEUGVgbf1e3mS9Q8DoYKO0W3yDSRNpMT/MprP6CmpgYK2uE2Lt7g68Mk
L1tYlL7YI9rOXwfZrsTRmVlRfEjI/u2MwXqA3H1nY4QO4MqAVVscTbwsRLXhvO4yTWTRzssuDRKk
/E31VMhPOO+VeyjWai3S086802QkMJdD3V4LU1cf1s0vQe92jKsnXCv36PNwxXQBa0PC5YoUtaCC
PGAh5i3rqtCIEgTUeEVbULv0Zg5lqNGSBByaEKz0UB+dP5CLQ7O4lMbbgtRPoPmD4YTqp+uV9FHU
u1FdHixCkSOfZNYEJ6shFQ3DWyCKIqib25BxgHC9uxwNwGNnZpAuqqZxtoURaqBJ4ItDdDzdjUMV
/WpgjmhyXo+Ovh7LPsXBYk1db72gOE5au0jkvUEKNIJUB8O//26sabRt04XvnYWsLaoew2ya2M9h
PaMbsN1m8sHaAf/gVmJMnK8k9zeOrdIFnWMsc9M2o5YmQ0M5OX4N7AJB5LT4vf4joCEEq/GfZJbg
GofPQjXcRfEFMCjZdNWUN5NtpfSoDEfWOr1h6Z+OEIUIjoF2cJcU0cruRCGpE34PPw984GLOk2kL
Z9OkN6Mi5nlNT2UOFULt8F5SdeJ9QWUBiBcb9X7p6xn1Hl8VG2csSBtjl7jyVhnavko9ltfAh9St
q9wtceViHOw/bOH0/SAS1SSqUdqMbMN1JJ/cVC02lKnKIS9cGSmYQrXgN9bKWQws+T70DiwZk5e3
yA0XguJtGaowKlcmfgaDk9GGAD6nNo8uDN4AJYrJYFRjrlFDFzy8O2T5b+9gCBtAEo5aiEKU8GpY
ozUtOE2X4dYF8zeb98/sPP/FfJfZNFdbciCxW/JcPy4h9mbCKonC1zhansY9QJZxTCPKqnapaTAr
vPjquNotZGEpn4OFmQ35jofOGbp1pJ4M/G+lzkdTXCQYhYIXipWyEkPsOxkG1lQTzlNZOMy02L6r
6fwG3yaDhAkdP7aAKmofx7N0/ulLVQ3OiuPhvE2Wwcut6mmuBzhfLwIi+Z88x6+6fOuDi8rvXzEb
IknVamA9Q5zXQ1DcQLdfFO5V5cUA1KOwVMpsgGK2R1sBvjxGZstJ94QUzK1a1TFALTVSfTWXkSVA
zXGqFo+csx+TFZ5QAng1O73t4HFW6Nkgf81Qd56gBhiKi6UtXDs+c1UsNxR0MKRG6nAWTpuqunPZ
cn9jq19uMairyxAJVB9LadI5/b5xoCiuyx8T1/LKMmyrd+G/pHuS+30oKgm6sYrpjBAq3mH7vqQM
wvfX2ikSAznFBdkh/puSmxLCQUKuiwYh3AhHuFBE63Pe7G5auT41xH0BvqEitWhJt7gx3+4BlEMp
JcruCNmvYvL1kstBSuNg2xj5vK8zCzFPZFFSmeUv9OVY60PozVomu5KYQ5cK9fu7VV+sBeVKPb0d
D03Ke4rly/XdfmHAyq9whxD4Q/cQAp8w162qp0qI7pR0GTz8QNqQM+XDVo2RCF3vdrhRImah2xGY
CB9TG5wtsz0rx/+zQfmPtYflxRGX9i0l9K1v6Kp4CnI4FBEVEG8QKplSzzzLopVRyH4j9ITg2/zC
zZDgGsxfJHmwPdCiZ9KYEra9cU4IMnOqP6dtoXS9TrvqahdZwx7WLF4UTA/J2oPoj3GBMxyKCtDU
gr+o52WZsQNU4IiZ/N08lTLVbrLMkJz8FO3w6muxa/f6fsQhRAQvF6dJp+HfiytzDQX3FjSUv1V0
mbNTIp/tSkAa3Ixnxvbt2+mkby/i6BtXPq6dhn/04wRVDqY8Xu2CaGljTl61xs+0CanxFTzdxKpy
rdleaQwi2CHMDBVBLq1qzwgrNdb94iCTHbYC2z+qlEe/UABSIWK4JN+NqXOBe52j2s+X0G1nGlTg
v8Egau6VN5BsC5MT6qN3n7iSkIJ63227HjDSQUaNTsn16uB9s7vjlxAI4H1zmKD/ls/hvvWpCQzP
cz9IgoaaAt4e4P6OvSRWqO/xnGaui1p/96jUv7KyXygGaZbxWKaRWOFMID/5s4PULHon46a3aynR
ViA+PfjognF/fnF9UxzvhOIS4XIrll0JFXATDH0fXEr5RJTTdAjFT9a5KxHExHuWVu2HzwEsh9gC
jHaE1Kz4szAiFWID2xpfMY45uVE7lC8kyV8cOo3SmOHlW4OtpmHUgb9hIJ9UNfYIh/ea+NZ3mSpR
SbEZQM9yP4zRFRU88TcP4KRlCr9L+sm3kXGYFauHV+lkMn/nYOCeUrB1hZ7GTtopOugtpHktrZe9
rGFHHbbg8ln+oJ4HPsEsqWwwd8TgqsGSdE1G3wL0nFj7xDCUBJmnujwbu65BRht10F1asSet8K8m
T1m3K9vnbs2qOZwZxugVcLUWL/ZLh+Yqaje0BNfirLZRcSMnV6lZuzpZSHpS1WO5rPI9JtmZsit6
b5u3eytCnmf1/fKxTN67RcJs/ILzHXSp3btG1sETgyr/b9osCyjHmfsa1U0hHeJqkud2rsSzLEVk
hIXWOZwux3e7IDM+2yATtUoEsXiUgDWU/qknL7pqIhkoQ2KkoMU2buEp1tBdJ3FmnYalcJdbQhb0
gJbCRnjDhlK0K7YEPI9zewDfGRvpYVMAKVwLrpnKXt6bV00TMw5tzJ/5hVr2zfeEXj+XCyoNlOBd
Kj+tg+mQ9doF3RLrwbXtyTp4PWiAXrilsaWEqFc5qJpWxMSWvGOo2jxb9+2pQfGTyVvV4OOwZv5F
yCRhIZCav6WyrVfPWhoT6+qt8RAStJ4axywlMVbwH9/pdMnHzfDaiip/96JOeIYX9cl2aITCNWd8
71XpTfOGpgisE4UV+PFLaBo18vzHod5IhUtL+i+cje83n1f/aHk3qa4Vb8oKcrWhuC9H2KlL4x0V
D5k3Nw7ejHdyVI0txu4JUBI6/WvpZHGTrDlVVhrnCGk474OJTdqGJfvauIXfY+WoxKHdoQEj8ny1
BvhokOnjQ2CBOL8pG3sR/prN0B5HCgt4aGyqWLF7K/VQew8+JvYjnHTxsxvyyUUatTCLNoMMJDrm
oSeXX3pUxOflCbUxL9KkWJwU6hBnMjJNvEWjoV8804K1xCX2xrmn9at4vNQoTreh4VFvoKtsq7Lo
R3kb4dp0jG5/G8fTNlnhgdDPohidcV1rrOemTOH9foWEc7NTH2pAm+mk9EWQgFxotFydYAC5hDAy
Cy9uPzMSrrv0/aZMfh0N/UbQjyRiVgVL3qsFk/527f1CF345q9haQbiB7fHQM4/QAN0xo+phfY3K
a7hlKYhufjdED5JEFprWwB6MIDcBPNim/UXwgctp3/5CHu6qwnxi7Z62keCMPl2b9PwHvIGr/LuH
5G6PXsSHG4XGDChTxgt7qo0cnXHDPuzH3lfvIXka6dGKHB6whR/iskod3gTpEze/gGZkt9VmVtt7
Mcv3TK0ZwInu/UFLgG7a9B5TVIyDnnUaA3kvXNES8VDV+tfujWMBIHWLotAlhk6BLt4pztkKC4GX
wfp1/noszVy99q8lx6v4dGVLDB+Kyp6Ildrfv50TzqkfvRZ1e470nM+epj6Bunn8L1m8MSXOYWHb
HpIJ9d5J9u+kA8B47NkzG+FsCnoqI9INvcMWLWyVPO3LUVNqrjh3HHvh0Hf84ZKqhVnQcTqqyj+G
2tFzVD7e8D9Tm/2DiOL0bSkfir7Zqv4zWzwonIZbHEuiRV4oC9Yil8tLWxSNrnz9qKSz3q/Y1Jog
ykIM6u/LU2UZ9otBOUhK3iX6srnUo7E8FMROaW2x0qm4pszrrJR/MYO7iq9LrlKHcY2EPct1NQTk
4pwYO/ekOHpnWPVoIejRlfGg724iglMZ+DyCwJRXtDNwIuEHXSADASdw1Jr0t+BotN5z3AcDFBIv
G7MzY5FnmkMNUK5Xvw21sdGrIolR1SIXgtEzzzs6iID0JAYbqrxfdmrch9if5Agqni/N7Sm8MsNt
B6fFIuRJlCH/oQI39zNdfyCJySkxGnvS7eiKOfAR3I5xpIFc9GsK3VMXQ8A+puwgNe3bsRgfxX+O
0c7Hfz4T3Uqz+QsOJYOCPtHcoFmnrWEKVGfAgpc8wr9PkeCXCWsMuTjdBvUwwVNW1t6UIU10NuQk
3bkI7sGpbG6w+p720QlHTVR8LjyWxC2klVId8GjzXV6HvugWpkXFnH6tH5G3Nb9rDf5wzfjFgYox
zPwF8QmBGsgxNsDD0HhXlhnnkkliw+VS55n2GcdaB9nzjgmxuN0tSBIKCiR4LMbF00iDeNHFChcN
BhAxO1gEFvkrPgR2J4lXp5YMFCK9F8pzCyMcnY9VOHN30kz9Qd+kC6adDDOhG1NFAbd3QMVdg8Qk
/Bz/IRTPmFzIMBhSDvUsE0JP6UGkZDpW9HenO0UhrwAzJ4TMaZ2ntZnKyMYN8wGLSsUD53IBu6zw
OkMaMacqtkQ+gv8QOPGIrGgym/kOdE6qJ1DgyS5Ju9xtZU4lSxTB/Sjpm5cai3Qc5T1UJjmMc+gc
h7FWsMylUETvDgulpAGlsXIZhBwsMeqcTLWsvDwuRluP4Vuob8Vm5oOmzPDlnisHBUj44qKXQzF6
+7jkp+GrFeXPhGQbRR7+ts2+jHstDqNGfi+HzwLW7wcn4HHdN9s5t2YUbkM+p/DUhnidtAzkUsoi
p4uXkTEO90XYztviG3ZWxW8zxFJ42aEpQWG7YbBxSTrwhDZnqtv1rRfWF+OKhMDTIa8+9xaD7jx8
s1q9Fe1jOtJr5B7DuSn8n1HkDoXX4nL0/ARNaAZf1R+4wzNqXKkJF4Vb92ZUzfSfmDjxTcmf0pNS
fI4QPU5sWF8LMCZr9kdhNfRkYhRjIitWL+2yn3T8z8WQURBrY/WkWKatVUbO8DxFzYdpdobYYGF1
TkWSNkJJ0/4LXYYl24wxMTESOOvDd+7MjBTNzgdZOUKh2GR43Zu0nKMyKUYGDyF2CDfDHGWf4M6W
W+cC/+Sel9hbU+c2DOcRgISp6bkkQU5i+tENsRzyrmRXlWwrONAXK5Bfucgp8xdLn6nM15TtVHXe
+bgS7vaHLRsfnyR7v+JJqj6IhD1tvgMmCYUV9v7lc3cQ5k//RcN0CqK3FWdaAxUkjd4hBjTJyGd1
VB3jFCg3Sb8AMto7VmZX+nhCYFuxzg52DI/Y4vcVmlwF1nzH9o7vAWZfxd7ICqvDby89acRmz5lq
ubz/8iXmP8PF0SEDB5nP3g4RQZs5VdOTe+7Pfky3VUGadgEUOlxfhwVsEs1AxZRUs30lG5+T51Zr
ITMzJgxlwMqhAIWar86XWNOy3JbIs6JD8dBvzwTEwkDaHiFvMH5RJfvrk3qD+xcnqCy0iTj7zfhg
sh+Hm9uiolINoFk3jzoaPloS9Ksu/xJhhnCR1j7JqB2K2XdV7ghwwIrr4xuZ5vkZvkty7j17XdK7
PWIYDw+1wn3f7NTVEws/7ITHpTZiAqspsZQJclSBx0W3htAtH72FYPHtOFIm+ES9DjAZQ2nViCWZ
WndkKDbmhYYTDe09Z6WlaULocGg2wEJcHbTTMCE1mCEzJ27GdjrK1VJEmPR9jA1TbUkl6MPwJuoW
Kx21jGBov0pud892DqbC5FaCGfyLWlTJRYNg7myHXthjOpaqEIJJz37vSg5LQ9RbiX/XUMjlw+u/
e8hdR+CZHOmb1oj4iDRRHukWsSs5KDosZrTVoDCFHqn5N73U49HG5/IUALBOkX/H3LovYyOfjbGT
71fZlPWdJnl5lKo/E0TSg5gQwUKTxb+F+KQfOx8UyAqg9xVZ73RwLPgQDuxTDd1Lcpt+TqErCAdd
nrFALgog+lXPk28+iNv+WUlgUe/bTt1Y5Pm1JtvmeaK8VSqZ6HmToRUUJa1CMn0KnOYIdYYK8OtF
K8h4ULm80NEt2Lc3VkEd16xWTHnuwA3gBSjnzUyi36vbAm+Mvbl7YDge6xKGNHdfbdNOJ3A+hH/T
gYvez2geOgKlpUJEo2820qpLp+S6Yc4vluVowjs83EBy35fU7AjyfpjKWRe0z9GFPNzahZNGQEJd
C4XxxnlSGTpZ04fz+f6WV8r/tkQRvO4iZ1YyDsqrDZp0/tuj2EIKlsj5n8VolT4gtaWiHIotKn1M
5vP6l3x1ICipLswi9FuCIgBdqv12Ec043ldHi8rGVYqc3W4c3e6JOEKexkufGC88prb4W0V1Qha2
DwTp7gw4IXKsYbjVseVJe4/dthQElbssyDsNN1Y0f3B2jSetFPDbb0yVvOHOmO2TgvwA/jKM09Pa
N2+NHd2NBJkQU/LxtwRLVtlDpWsSQzj5Uy/nz7X4jdsmOYkWx4BSo1aLTfDGfu9F77cJVz8A7Q6Y
DEy/Psdj3Xms9/RiVfbu+HkPEAaflHIOH8srTPDpQGDLAd9i3duj/a6uoEw0xvXFbBU8I2WJ2gK/
BBLpD5CXb23GO4FJ1oQQFYniYADZ3gdMQ8iQ5EJgygww9NeWceFKjDtuw2h3nUs5XI+8phRgM54w
1/5uErZbQ0bvsuIQ0GMDTooJ67hoz42J8a5rwHnz8LU28xxFe7F9Sl7hlxuTYtvkvbVb2mrRVtQC
fqV0VurRWAQolx07EhfEuDr3XKpgs6JY5QlY9Y1EPymPO+qlSeUtnYOWgXDyWf7eYengwMtf2aP2
jeLvnzvVcTGLYRM2z2ToEo54DgDLDKYMb2axVE+Ut1Iq7DqFz2heyBbPoScZvLnm7bdeAPt6M1XV
PIRSHtv2HkMqgRx1ZjcM14MW4KRVv2aamIPDcMu9t8AD8bflKjcVbXkRk/inOd3xBghKftmwFkNm
NgP4lkzndQ9hPkFUFIkua927pxwpvow895Y22Mnh9C7Eic0t9QzSc0Oip0ho934NNTiJF2RROke3
TZP7yUeyx0aXPjQKtgezVvtUmFqvhFbtZh1iQkg5mpK+mzYYzVAXCzLG0saqLGce/y6Il3/DXrs/
HvAPATy6u7kurEwZWdxvZ6g6onRJ/NZiGc6WFHdKQApKVXJIRIbIZQdJpJkXCcj8dOZfxsOMgCzI
PC//Y+i/M+klW1309PayAS/n8eD3VZxS+fD516heiWhPsTWHtasO+d/GcTyofn7EmVr2KnuNwU0z
+fgCorhE28I5cnSkHvwjIzXHN0rfsCuVoleBx/pPFs3VSdC+QzFi/kyy9EFa/4ef7/ekIOGtymtG
58pVYMjE/eASaAVY/DTdmUlvdp2xa72fsJpsFTGvxf9/tBrb7t3fJEbXQNof7piWypDs3UkhkJzD
t4CTqSYsP4yG4v81tSNF0OtZzKMM/I0BHoZgwmRYTYVLuWy6YTPstyzh/NtJqaDiguwWy9T0L5Lf
d+PhzvBX0abGy6aT4EFLclyMlqylnD2sMSikyNudek0xkxwYkkr1yUQgYjYMar6nDxFyw4xRtWNL
r5DNXFIszqFvdpe8BR77EKQdLtRppsQM7duXdPb0YsJWaDZYnatKEjblaB2b2aP2Ki7l+JcGII4t
1BuLiRUFEx44nGeq5a+JgRtK9NQ0pR2WVVvaWJHenDJnqCrzWtUuFwNA/bEF7nnSAPFLlUfTRZ8F
I0bRg2b0Ys5nTfKpfnQ7UuS2v8QAR8VThPRjV8NBAl8wCuqJf2PBjILzliK6ZPdGrqqtMxShl6Lk
1erAi0lDpMKLzqgQikTs/nTxhtOAVcAOrtwfLgkZetS5fwHwcjqSidPMlxPIxBamkPIvJyGsmEag
lIh5IWDQStbEHXTk3uGc4Dqek3Mi0s50y1zfafgy+2Yl8Cxlxv+y76rfOkU7Re/SPHMB2WPOvMYk
KVBryOsksMbwflzXlrfSmQdwOVjFsDiQqZfo9Y791aygfntjBMAL7iFWFbqTYS6Q4oT/kqZfwPVg
WLj+kvjSvrHRfXeuHCrfMUKJRkY51IZQ5wh6WF3PnQNlYi6M2K92+VzCrUcoGr9FuG7rmG1qpk+U
rW4YhHdlwbHtBOVGlXCHV5NQUY0dp5H6JcJaYodM0ROB+U3MEDn0yG0OsRBIJ8VnHJCkR64OMHVX
TpnS3kiVPkDTDF9XxZDwsATMbST7x/0vKEblMkPcZu3v16VtBgIzJ3H8cPEJ4NmSHggWdN3nc2+Q
1GhjdAmnAal7VffuCjE8lfFvMGSQ/hjpnlOt8RSV5v0S6sK/Sh2zJP71+APVMvUwezbZ269IXrxe
k1hii1Rsui6ZqV1ed5hsYhNODqE3YOvAIHJKscFhsequyVT4v2odT+SP5Dw/hHLE0xqLATCBW3xP
Tn6nKqqEawFbV8CeagwlvanRmXoJEraQ206jlaqo8UuixTWO1f7NyIBzqjdR6gxREPOdWYHjqfcp
UQLR3FC+jhy3qFDD3JNbU6VdKpMM/vSenwiFyAObGd26qwdtB5iX1eqKsp3FA+5orXlMuTNoe1fU
3bL7yaXJFWWEjFu/XwHDdO0xupKcOTPFzEpSW8O9hOXqHUqqtviMJu2zThdsB7ZDRaN6p8CSmuOk
XW707eYkcY/YGVZJBZtCDzvEN34lh1Mvm0Rz3pUULmy+uERoQUqb7usNd/z/Ej/54FvsEGhroPhY
p2DsXSxM3+0W+KKsQWQZNIK9xD86T3PzSFMYvH5GlRjog2+bkxB8Qg0G/SQFpFcQeX+g2gHNTzJU
DiqQArBT6Ez/84Yl3/zvKG1gQvqVe1G6nhflda8lJzuyFitIfX64kBuEg42qKGh3M5f9Bn/3ksp+
ox7Na26/YTswiBSqxICjPylg+wNfvZisAslISfofKOCRIbw78oz4dte7TStC+F0iNeGphkLwcu5V
3aw76JoCCldpzT+rXE3CNku71UK6Xf96iYSeqiFfK/9IDGdQ3Dz8CSa7Dc9E03lYjHBG+tMI28bu
grLVdLyfqGLzkk1uahCUjiFeggwcP/mgwZn0DTKjrfs4fuipSq6Ayfkrq2dVQ7k7T/8xf4yEWp08
xQkFd35S3e9g/E86nhYGlT07sNJfC4XQN013xrthIE+kORSKOjjLGxFW/SxU84QSyoxlemlp0kUi
2BRj2JbVdsTpt8Hd4U/AYe7/5q2TxTxCvggkwN4qvjfv0BJsLDbPleJqAKpXkk++2PSrslvY3o/U
bieOxAUZvZ92iWOOwzFvOTOlXs7vDMa4ut97CVIM82tOZ9dI/8Tf6FGT9QEvX3VhG+/ZQwBQBBYU
nVqE9APUZ0sdoyGpJEk/QCzszYN9ATOStBZllLYB7LnEI6B/NdqWYgmafX2CY/llIaCESIn279a/
UM8jG9nSREffynmh02dxZbgnlYvHQ4a+veRYpfaIBSJtXGzcKVXXMwxuoUgDzxCjKurOW8tcKaJb
Pg4avh2n4lqOEYe6In3GuRBbLaGkLdmm5wLKokjHIc3TRncRUF+AYP7zFKiq2zZ9A3XqrBNvsdT9
IgDRLxepuwL4rNMcWOrakK8tRW8mzj22sl5tkSRTbymvhh0MFvFL6779rwq+Jb6WodaA3bMiMYJ8
Kmi+qZNfesUc4MytjvPUL77xXSI6Cst3D0T/BRcfrcWsPSJZs2mCoCcJLg8dVu5Qmpd7BYiICIpy
AJiJExUb6Gec3c/FoyMYQczA0qIBFwuLW2gdRJlPK0UUBRVCX54rE489+ke9Nvpceh4a7eWITdxa
j3D95fR98bgn86+bpZhSDLPeVtzWHo34Ss1oe5UP+rMzoioenbj4HRJloa6RrnFT/59WaJpqywFg
BuRYuo5IGmLiu+0zk/5RO53DOlkbUdjOvZ9XhZEYWI7kTYKlGchxlf1rm8ZsgGuVpBDkom1jnGOa
guPfPNueN1K1jpUJ7KP9EnvpoT/qbDhNAWJpdgHQ8hz3wTY7P4aIKgyY9V+BZF4NN1B21xLLd7wF
1spR5KDWjWyg6iIurmVQUh4Jk7UaIzyOr+Od77EpfGA7IBAP9oNgBACOgeXWdPJ5kSCoJoaPeg/g
3KSAGCsQWKN2yEkHZXrTpCWM95ZXbDYSpxoqP4GyOTcmdSVzeNc0S6c1114QAtnwrsoGwqJilhTL
pvaMzlAQ/II5/uxWFIL28hYT2zkAdQUfMhdb30ii6rJ/HNIwULNXJcB4fw+vIbwe1SFpp2E9il6x
aid42r0owhhVBHRBWHe6CeqC37YSapG0hfhHhjCjo3+HNXgsudA6lpulL10RlRmddVN3CjUvbe6H
8agOEMs1JuWfT+NZ2NAXjaK7SwZhTwmgKqYo7O/JjwhpHH0ome5ObOAqAsQhVSi64h4vz5K9x5Nn
rSApzn1GE/GOKDo+tmsGCmGTp9V2LfK6l3aeOBpNmP+Xs4TfpSzHiw840elEjClNZajjwxBRzbaV
ELrI+0B5nToOoIkEZxsVlByh7KV/cXNY1+Y1vMsuxOJ3aA6weOrPJsom8mZacMOPK49e1B6TaNDe
IRIFvKgcAh76zwtFzx0bOU557Sq3vQARdSIZ8PqdfkH6mtvlA5qKtUO2KSRl+cwwytDJBa+4vy/q
KUcYs9FzvgzfFT5/R7wGO2JALfKTypqr9RawdKxidVeNTQsJoufyV1UFg+K7PFguxIURVYQAA5rR
ByVpeGftko26147TWmzaFny2qFmRdZGwPU5p1vKYq3WP6QAWfp9dpjct26CyTKqAcg504tWUOw0I
FfAlVp9sMazgSAskFSwEyw9FdO7DdS+UqGgoldq1huMXm8PhL4PF2bveS9M+hZhGndmtI/lj+0mx
jIKxWMX0x8wx93S7Ux/0VmMb5Q72Ju2VD9pcB6egAGJsyNJIK4qOaY3/uVR4s1+MkOhYe7I9i7WI
YzfPOW8Y0Eh465JfMXs1AfZmoT8466HyS5jARiUXZrhjpVPnm+tUA4tPIxbAT9EIkpPK+v6QBDNb
N5WO6DCrYyrsSAawSHpYS2XcNpc20kU68Af6pLNG8ZmPB5QCRnR4voi9XL+I6gt6DUuVX+GxO22C
XT+rUXMWy6DH4Fi1EaVXGzDc/q8TPdE1OBFCQevcX0rLCME30CM6X11GqKEzKj1Gy1VNEaqMNMyK
9DimrP4YlkGbmb3ZlSJTWdd0Ey5EMQgiiEULvD0SYWOQg99WLEMCiyHli7Lh8czWFnlMuLuvMwrf
oIhVepJN/RABVaM04CmQ54/couhtdcGmJzQng74YA2xKDI1BmuPbfeHwASSzCGViXHBu+rsPcGwC
Jx7voYBL3Fix71I7m7WZaw9IioysyKUVvWmiWPyNKg4F0NZfqRXSeVoursn4S+/Wx3fBKQEYlXK7
FJvVoI/7KdlZCvKtMyKgMet5WX+CRksdnbjAt4mNJcFeGXgJMmgQ6odtXl0fRXgq9JXhmd6Pxflm
bLWytGrRuSHrFwaSaLJVlixHHnTJ6kBtTZj5raWCcFL71L21MzzcMopAxSOHf9Hlb9JXpMet2hFZ
hs3XjE2W8PpXxbaMkaboOZDoN0km7VY/nUQ40Trjh5svbaIHbJ5hesP2PIhXbJRfgpm1ePVr7rSt
FoLJvcbzSHxR1gOY5lZbiZfrTQO1Rlp1ceAA2MLaSN0oFjQBj106ir9V+dfF/M2aFV1R/j49UD1O
alQd57Fz/ujGrm360EhM3c0O0wLq7iWB3KX645EB8itrqr/uTKkKFYnpNmVxT6n+iL7P1pZcvZah
lSugtYYtQcoZUwu3HMOboukw4UpBtdcjU6Mqmq13c+dX4F43Xy9GVVKmHjHTIKRq/QeMKNbjjGuH
mcG6Y+58L5rZFnnXA6WTA6F0n/6y65o7u1r7btUoTbzfEs8czEFq6rgbW95uOCFpqGUTVPtlLt5h
yUoG3QBdbWjWhqURX5JcOSUguU9fq2gyQDNcbwmTRSRRk6IzY4LiIjifk8ihGnMdmtP06qRAnh0n
SrSMxCwKEACf6u0KjQ//n+Gpy7D9HFUvHH09YyNmfsf77dyAzkCEDIK13b6gpASqQwHlCvvrHbjf
NYzN1qAlsDBKvjjZv6V9JjOKgvqYuj76B8U752J8DqsAZuRvyw1vf3MB89OCOb6Vpr978lRBdq8Y
0WHRNIP8Z+qxaN7CRmn+kb6xxs81xWqGW9CnTWg5Ke57iR8X4BYSxAi+YEr9oULw4kD3T48Dku6c
hLw8PwkfNuMx37B5+4TWwAIolG54TTNXF2msJVbYE9uEZO0HhmRqPWQDkBTsqHPbIXadkTBlo9Uk
eLsIf2gFe4DHp1N3idPmORz+XCKPd6Bs/7IeH5WqKzd1+JV5knDBRalcF0yTCLUruM28OVKapOiC
Ujt+FJgD2ACNRwQGx2OuLu/jjHGMcuEXtnXGjAW6d/8gOo54FYsgwMF/UI+hhWOvugZPcov6EsTp
bUocUxne88U6+kyziYBfU4EX72PFtvLi2v9NATqvwS7sGFKzxHrkZRTQlVR8/6akTgqEUfVh035F
xpkHumtvzkYeMeRnDLR+508L23GXt4hHW6/MwXycrFMkYi0P6XEwb+L2IdufzGzwMOPU9r6HfMpr
mX7CKHqWo7IdLuYQ17hppXeDh7IwSARjefc5cEGkoEwlU81cYVnFbjJyjthAO1PT95bra9Nnohc4
KdKBqIP2/KRMxlPqgF5MfyNNVsSF/gMGvhRrrylqd6DSlUE/wp5tmwXCA8LmG/ZTy+UpRhtR1Qpg
LpXZLy6/xv1RfivC74pB6BRS0fjfCW3c1iTw8htkbXIF+T7Nrfpwg6uGEiNFXLf9No4V5Udz12Sb
qcJqepjSUMHoy1CGbdzJ7o8DAdYY8wnCKlKpXsC0MRK3ptAr+NrdNsxLGeMSYpOujLeGPAs0YFfp
YtiXNT0A3HNSvT8iGYaa8PQEQrb1Ql2LfmsevM3FqExs315cCImr5xqg5QcetkkI4B5b5zZoqBRB
q3nCVSlTMqENL0VYDxoXouEQ/xJ+Usof4bkVOW4QOphpDhJRyRcQoJqeBHLhFKZ7WV+dTOHdcupH
OlaYsak6rzifiXuq6aQ0m5mZadKOPyxXQ2OvHMdHwcUrbqXxAyWLOTkMH7nI1dkRH4VxDP0Dw1/9
obAwG/Sa928T+Xel8I09MdJ4hGpD1n9UGNlk+aMooQAkoDQvvX6UD1IFhMLxMV/2VqWY6SeZoJso
fJ7Qqj6TT9flUPQTwySSlBb40u5jYsnKgLc8l6NOf/DNlXYDJQl7z6a4e8m0xAl25EOVnxLEacRs
x4MdA+vdWq5zeeaFKM/KDt1wAZk2jhouRMlzsiL+sa8dyN7JTZasxx+sr3uWcCnYcfKaV5tPWsiH
TkieovUD0zIveIUrgGMEuIMKmJQjdvRBs8sWlyxlMMTS17l23RRQbEgHWR55gpDks38WtWHTPI3F
18A9zBE/SG+CSRCeznlepJMpIwu81PQgRczrsHt/s9bMixsBr3IfO5Kvhxstt7mA8/CsPkAnVICX
BqRxgxJ9LkjWJ87l2c6uC1B2uou1B6h7QIAfTVND+1/yadiZR9HEP2X3Q7ZuJBCEfSCGov6vSTNf
YW3C94Tpg9bP0IUHRsNeBrgebBaGI+sfWlv8ZPfZ7DTVDeWjHPFGvn2SrkTgD4Asvq9/WgrnNtVd
BM3w4H1kufGw19aApDU+leBDOLnR6vYR12X6mIcgXy6c/yknrWEf6WHPIMjbA3GaNAUiPsmIumOo
YGIIEMjZdETS1xIA0JsevUsaH+11EMrldyRe4tXZs/ILPISvqLX/2xY5xbKyBpHlZSJCs+j8XDk1
9wS1pLYUeom2ryLfEELvdjIPwSFNbIAjg/WL6clpQ/047LVP+ampyCuVzuEtYsLCh7f9D6gRd5T/
a5zMm30G7wOevT39r3l2en6AxGRDGN4V4hJZSXQouTQKkxDXh+wc8/YSHDwOQ7326A2og3YEZPzD
xoTgWom9eUwrnS78hMDJ/miMBcl7khpgESV3LYYANy5uxiBzpqDd7MMHEYzYENmZ3nxxyeypnZcV
QDIB0p8WibvV3ZtXGrm/DLGdsMv982jZ5KAnvSFrfmtYZdbPvoS380P8wWvI8taWTUIx8oEwllZ8
9jeudqTdAj8dHgJ5dAzrezSFOBwqLDoPQqNT5ImYBYzETdheygpiaFeEgDYqNOsjoRGtilh36aw5
BUYLGrp0rmNf3dxKgAYIe4hJwEnQWkCnyn7QsxrZybYGTLYEBuiZ6YQG78qT7eRL7SPcNZ6Fv9P4
E+nWIIsdC0keAvi+BJNGKvpvtpq1p7mfqict1q149dyOsAclFn3wV+1O+jiP1Z/pSmqxUpJKe10U
7rYRiECBjT1yuf0UeOnyMp0BDkbK757cHXVMr+CrnPsShN/+7LMCbSuJlA5WwPtdLwcl3DYJr/jI
B/LlJFYqKG1Wy+TEj4Ur6R/ttQRrdLFV5oLftsVqG9ub0ObQzWytgCo1WQobg4LSLvo/FxGT+DyP
JkUlDdsxlAxZeg7orND+xsHP72PmcL+QU6RNjnYbcXsYFGSgVGEypppitDQM2ihNYE2/ctb/BBdz
YAmc0btM5YZslihTxNvrIY5E8mAZQ4+Kn588DEQnKKnzAPDPc6/OE6suLG518H2WHofZlnepEs36
g/mvFgrgiy+6HvD8ux7uXRcMiwrhd/WmHVVF1lnuy42vW44ZJj/1RtxE83VxycAxC9iJ/cyrzL+t
MbK3pJYUOuYlCdVuGUETdNmCOZ27SbigMSjksYD1F3UZm2Cnrpe8Em90V5GZ+qk6OH4BBUKv/8CB
H7RoNqCEWgF0XUKDcQLgXTStWfQSCjVYoItWU41Z9FQrK2QGdg9sfUhsyB9AYK8IZEQFMAU5BSIm
SA8t27k0DlOEoGEwsUtXWU51C5smmiTcudW1ejDiFb17onuA49bVshhU/J7xWqJja4a0EWD8oZMj
Emy7VfxVFCrI3fC9t/FsvMq2+D7ez3aIHoXH0Pz4qgGcy1li2cdkzRODSf6JAOQNHvVKpEbUDfW4
Yk4JNfnD4FUdFfE+rp/bgMmzvxKgQSRKX7SqQxBGKiVwFBtsbMAALbhGQ/ey6qdtfCSzrTzyOVpS
YKyzB2TSwiEW5iR3S6TB0RGXVzi50z/m8MImDGKUpJYRdTNScxYqJMkcIPZvpQN4IqQWVtqVcdm5
fCdLuiCjePdZ3w/wPmCEee9RG7mKrhgdpwEcS44a/eFMeFQ6aGyJOlyk9uwU66jk9tFg3AooC8QM
mJNShDaYBXoWyEmqce97Ffv7ZRVLMlHTq3LxynDx+dLmlXB9CzkQN8fXFYODGY0UZakQGvzs9Vvb
B8DLmEKc6WrbL5Aop7Mhhn/M1Xg3CfWfT8kAKomF2YkQKL8rzf7yFVQzGRWIWx5S++2tXHOhZW1V
TNCIWB7bklgLWllev3HSP2IKh1HLjgrjUTqRJq0ruNdTjXbMEr1dZyAVXX0DhnDGPnOAhUbvdD9N
ROUeJwAy04tTgvrgLG67OXDmIXCnt/XgvveNRbxa/wN41daMqyzUKW2ZEMaOvh77j8e3qIDOBME5
ucVvssLU3OewzTQnhTDhVwe7T/PhCFt6cLMncr6GfXwX3NbUnmO+HSw3OFy+sMvN2BlsmliOjZPQ
/TSHNrEPlQJc7PD8rZT0+qeAT0k6sbhGqeAETyxxQZKGnMaPTdMfOK8LjY075I22L/IeH5/1fr0o
l9dtvc4X0+YZ1MwuWLuHQ8G1pGg20aYp6ytI1RPLt1M7cDTpyOuU9v0i1D/2ZNApKvQp1ohCpJgo
8oV+oTs+yQdFmGAhvMHedIDhloyMe9DsyPXXHEuJ2s6ZhnKw/sjSS+hDadCxhn10MZN3RYjWyBU2
fbhn9YJZTNTWp51j8k7eLTi7OQeMCAl+Up6Ef9fKln+GQaFCM7m+jhQPx9lvQyzpbbrIYG0OGMAW
04PzfpCLM9PGMvIyaXzxjWssnmLQ5iA3cK4uICkn1RW3egvPn4TJK1R8mJ74TkvhlvJi3EQVYP+k
kxeCKyPUoakLoqOn9FUF419GTVysOJ52kkT3QW4T9N6gRzL7/8JIpggwUxbWZnxyTYTv1/GRKGVU
n7xFfRwnAf0V5xP1mAqfJGwGgVzaMoQgOyYTxAsC4SB7XR1APZIW/WTbWwgP5Bn3DyR70AfVaoqN
hbaLzC5/BRP9QV0zB79V019GxtvYgcZ1a9yJpH2B7gChArFAYKItsPc0hKNiMcYfUN5LrRVEKEDk
6olcVmcE9B1edJ7/3DhnbxZ/uZd3d3HhHifGeZr6XL3AD0A/CE4CviXA+YXM7E4iX6Jt2gIGTlHy
3mYTKLMeKxcyIsQbYkmjaZNdG94qU2zljhs9nM6bnBqljtJIrSgHkAWAxScD+LF6snAhDeKS0COY
QYBtkVFIz7rbIQOmQRNv0hutpQHi7p5t4aIw1/uJ+SWiyjMQzeEbhJeCoUcwukwo9GE/p9QmIaFo
xOzAZARcOki+UU9AJyJURK0rk4D0Nxl+naDQhJ8lhsRSXuyFvn/FiGM4AD0RrEomZzPGcvkePy52
Vvkr5zeFlQegvc8AJSb5s/VVVIox2LXHieYmTS2RQ5WvwXQDMoJ8Be5YVy58h89WrZl0ygJGoOar
vMh3IlfZgzalBtEmtFd1FRVbFKNtd3Hv3oxBOemQS5Jz6pEtrBzRf2jUXEWQmXsDDyzBHpKp+/eS
hiGHpvGCNCIajKSbnT8p7AseTOG2A7hlMhaGxBcrhlaQH1txFimPo0vlZRmFHYmPpXXk3rYDNw6F
ltoTAp7T9U2cFRqnlHuobcIgXqV5jKiJ4K1awIUWZ0H/dDFerrA652nGtq6Os72QKZI2GTOtX9Yf
4kWThSd0Tc3XFCLkhgIJ1c9TZSsI9mdk6+JzubW1VfIX/dNZ9YtYllrjuG0U5K/B1yDjVmWeN+tF
bqaAhlZXobEUxo9koxZMli/pfIos8BNkceTo73XkC1fb8rnNYjUa2tEEBsZdQBR/g5XtwiWr0mXR
DSUBXRDb6RwJDb/oPyORwOrSMOsZ/2pt1GVrOsQmwzxJ4AjyymJXsuAI+nchgNR/zEa1fxBLmE3/
AzaAlGIvP/noOvgA0AmGKYHg8WamtzeYIepIjQ/QOEhXbLhTNX1U9KbxDWpkde/v8fE/FwQFLfCy
vk19yYaOyc1NRxRfc9CFsLwzissbU8AaMzjiWRDXFrLR1osEdUb3at7MDFyE5zqBod9GdKHXci+9
45oM4Mb5rOOT8mEnY6+WZAcfWLp9hlOIbLa06rSFOiCAIE8S4ooRfjOmRThCYxdudkeUhiBj9IBC
0VJ3E0GAinzK/yWvsY1vK2HLp6pEf5pFFANO5kVLcmW+OGdyiElraLSODgYVTuN0FH0+YM78MKPR
fbhJzxPiAysg39/U2sdZ0iZNQWeL/NMzlElY7YFeF50zcfQ+LXMExc9XJ+mTG4Lvf/wNrqeXKpcL
CGkTclIgbt7II6AxwIkYbSBod7PUf2zjENfLRStZe5zmPtXDqLd/qyAJHTdOTHjjFZa+U0g/jIlO
2vRfwqDDz1edDpy/GDdyKqDdkdGLtMMn20eW4OqczFEQcsmy1FqXl5lR7XSEjdmLnXKU/cZ43EAX
P9pa5uMqUs1DjMWSOSNqngksV6wYiyAhylbaTrVmeq61iou3CsnE2Z3ANRCUuyiM2vULV+b6CE1s
rFPf7T7/8Yi5iCLIQJy9Xm0eAGv8YGxmvFhTrcEzXY3k09uZWP9zG091sEteslArWGJojWaR4MMU
mOaBBt1HkGfey36m4+oRmVvY2taqpm+BWcJT0ACHi9uSXWBtUnzkiTsDN2nBiXmHQrhADAzEh4IT
W8DQS0aM+L9UsjcsxgorM4bc4G13nim6oenzTSLg945b3bNK2WnSdDWgLXAp8+Lsb8CmviakgDqg
/Wn04hbbUI4HHs+pd1wLXIzdU142NZHfhheGXVpZGqf4HIm3KinDnhrdG1XRjQx1TvwKjqFP2kaW
D6WCDYyRlGAguJYHugoKdJLZzmyDtcQRhnCraYwcIed9fURyPbbClOMotvPFqmjQPzjQsr8mHx3h
/yeqBPaFK3Sks5+ic2r1Mbp6oYBIQS6h5yu734zPxEMUNjlsi8Gu6m5P8y5QIPB20EaSf6v3iJJI
+6R+aRVkTvzxZrNApop2iwPKDdbuknk8gIGEXZMESPf/TlMvdytlTnlkeydk2T6yQ2HwHY0lkQiI
PNTlVosE4+Z51mdFDILvakbiL3RgeVuPTsiCb2gNvePJ+7Juutga3PZ3AWdB0S7jZvY81A6fUtp1
LmQAjIsH5H6p+XdfPgVVjlsaXMbKDndDjGu+jQ0pWMkJ59KKTTpgfglcWPcI1OrPndZtzuSjXrNG
sIvFJpl2iag45wSpFZPtByKB7RSTSdix8etLUe0bHHODZ1Z6/KShJKrKd5gLvfW5i3CEX47vVJEg
NJ6HOefkAJBf0KNvXQrk+Ka20KBemKYAO+szRIF3PgDkfqclB5q4jNQzQWM1PKFDqbz1gEqM4GM4
ROyegs0m1KfLF1JeCGKCOUEwl8ONUpiZk45xV+CpTkvKz9/AKHyWBI2AFmPI4hpYeu2hzxj9HGsv
R1MIHebhwsf3J1X+djJLyB+hu6841vk/P+XnBajeXstzeENxESQHHRXn+Tstrg2M3+hrDYN1DZFM
P35aCyCoufRe5WF8Wyh3oCmfVPKe+sNzZ1J/aDAb1BdEaNLtzg8vGSlqiYtnuDIq74SDUev5KXGg
+Z1a7Tx++hPCzhlNImtkyrXSotSDPJgwQDfFuqygPlfqin6vKhciDwJxsDWn15vorr7Ms47S9Yis
WjKLR1jpFjaWep16pnqiniuK/98l9mtC5GA6IvHvRXYE11cW+vi8pQIOL2NzCAPqOqFG8Z3wHpAn
Ghs7uopNtnXAMUH9oPlZJPgU+6ZU33oT/32jmDwmo8t2ooTt6RA/bBnkiXo3lCw0pPiXH7MGC7qP
SH9BnXM7O3877vFEaLVFj+tRV5m8Afp2X4buzWTT9im/HgB7rItwtKWk1L/5cfX/MENpi16MCgYH
ZAAmKigKW4jCbIBUZcmomdB7rIlWQezGg0EQce5mIu1YO8+NA8//CKONn/fuFdMV4uOxoOeoCmfq
L36ADbfkAwGWQ/zrESlK42JCXqGXtEa4ZCA9KguEqRzaRJtheiCwMxCSPtE9aMFA2QC8YuI5YpiT
8c4SLrXn3BPtUMgtmCse8exeHtH9UtM6QLiu87eBm/qXI0Tpz1/L5RXbcbjrDM/4hpjs0Oy0ovrD
RkWP9SWR9UEBlGKHUiucDCY0ai6e1qP1IiCcIpF432nNQ/VYuVxuYWZ3C6nNuuKHR+OG1WGLzs8z
4L+ONyVhoBKT222vAlrKmV/Jc5sSjy6+EGJZF71hniff+LzztASubaORcM7mXN8Ss9jM+tpd4+az
F/0C01Y6tQLVa+6Y/Zj6AXxj8Z3lJPoBikM02V0HzJJii80nntS9qPbp+Qwr3WBI1RnxaAiWzFKJ
9hr/1ZBBiHLD413vNgVcDruWexwjBY8CgN6Vp0Jk95sjKhHpRKHBXgsvCNy5UnMVE10CKEjE42P/
diAz8QT8npMw5nx7nSc2OP+4Sei5IruBLLXxPb+/ZY/yRB9VZ/qLy5b6sM4RuX3pd2L1wMT+V0N/
/6BQbfwJPUsxdMIqvxIdFK0zzmE4gUrXu3yMR2OAIjrN6Xl4wKly99s2WRdDrs6vYTl7qIA6bivF
lzXfU4Ce78x2Oi3V3Kt2eKMExeXWeYG+MB16QJKthUdXunITL6bwdYKDPV+IlS8a/Fc1yTyhVrvn
GNRfkK3V4JlOXirXb1XSb4NW4e07kki0rDe2OZjSGWAyyHVB4OUOZKSSB8+LyfCxOGsLSDcT/5tk
QNpzglnaGTvP0r4Yi2D76lcdDAdUgiTaaKfpv0jiUUU5V4lSsEUQ8Qdz3M/XQQx8q2nGPLaOTgg1
XvSwWmzuk8+m45XfMObs47iiYvIZpJQrp1l4yTgVd3XMG2fD+txl0Hvh7fP/KaIB+TKkuQKq/WRz
nVbLmp/n+wJolVQzvbwu/KKg7/HGgDMEoEMdK8RylDW1sozRgtE/x+9U8Ev35p55qZpS0LEMVg/A
V0XYeejGltgnEOTy4E/FJcjGA/DiZW8XqRWNPhDvZDf8pDjHgXByA7jBZlW6UbpSDK1V9Ph/WBCz
R5a/coqwOvq+SUQ4Lf+BHlnXOk4pOlcsqpK1w1K6m7kvBIweVvDJsSVWqs9o4THqyJUHGBNIL69Q
ynpRIm2puB2AzMX71H/Dqr2sp2omfdNjEekEBjkGyVlry3KD+gd+Sn0ALGcr48vY0uCmHA9qkddZ
mADUdFcPSZ9FepdSbU0Rr6PUHroJOWcPhKGNEFFboDLBHZEaQ0zbfXm+ix6cfA4ZV52kSRg+Eum6
OG1MYk6cCUyQif/3t7yZsbBZe5JFCLdoo/7cNTgcmtVdqB0/EykbkSuoC8vSHs4Aon10vCRz6Zln
FU13Dj7ILDHbpUNby1W6GGCqObFkEWFXOezD62MMweqlAme+IbDb/e5vdhJymqHQV+w8Eg6MUNDa
JzbrMELu+0c8ST/KgM8fFc55/o6zdxpGhQiKv8hdI1aaNzEfqdPIm1ju7Hnvahac7Uyr8V9LHHui
2oeG34ZaF/ornRG/iNAL02yaadS+2FACcZh1cNlRUZqYN2JotHXPmRIilUNAEXyYWz+v7ROtiDNR
sjegF3v9kMT3BuBFEypezdgqvBCbFFqHA5TLABJHXMGgVfCIEhv7Y2MVt1GJ1LnBi3veD4a93Uld
upErjtptJ2eNebJs2LKkMj20IXsd5MvRcV+oaT870lDJ/i1U4N4+6YXlUyfGysxXbN87uimWfvYa
HivJRLClAiDkiESRnAlAIMV94o+tSF6ZQnsD/YjssQNA3KbRlV8yyD751NeQsTo52tfB4B63ILRZ
XheM1UyqHfmsPxgrPlMhNqJCz6N5Rhr1o9AaWgGvCrHMloQgIwCmSsrelYYzGsxPyHlwZ2W3TdVl
l6pQQlrwNDWccm1MiQxFdz8FaKbS6LNst8WzRqTv8UBGnx7RtJGD0IEf8GgvIDcEkbf8kdLpMfKY
jOHQv0OQmSdWwJFtBnVGIDzVzg2ql/8Hlfo4ul2Nl+lyQm7grWfACiotHOyDV55PDGN4uH/jQlPt
SZdrdb7mSTJ93WAZaL3E4cOVMlIocHfVuuTYO4x1Hca3axBNchVtdESiN4RDDhqDrmQM4b2YsQK0
aIoEgjIF82wRIMF7yKH9rgcLBNgsE5wQ81oYanLINR3GQJG8JYsxib5p4VvKLfpF9DYMHGRcgl41
hp0zsDfR5p19RfUsq8A9hSFLmLNkx8qebImo9/tzSbJJpeexajpbWrPRLWuWq7jwlGdK8vzFEYlU
CL4YtojXQwkamwUPCQ7BgI0DqXeYHqjyMmDTvTYX0oYmem51ulci2XYaqu+5qlPlafmO06s9kmzw
rs6bxMPiYyLkJEDYvepVvx8tKY1A/mttbyygExuT6MgXdqNtRB1lut+P7J6zYnbYkYyTn/VveTcV
wSnh3AI17lpivDTh1qYIlkt0doWrjtNxFTlsax/+CRg2pGjX22u3bWtQiOXveRsi3I/VS+uFYthJ
bXz6JcPQWo111pfaiKmdXuLSUqQP6JdqCG51ZykwpgTuTrk/F+kvJnjwHuzzZBWB1gQFDFdwR7+r
UTEVhbMWjUYJPcglOqgai1J2Rn0IopLP1bOPt/tQXrNrgHwbXWBnvXZkMae88DrnmXu6kDymDu44
fdR73uV9k6LdqI5a4cYJ84vArfjDLKAs40+MubOwHfkts8vqBm0ZPRGZ+fjB2Vhva3me4G1C2Zin
AsOd5gblsNzib6fsNSmLIUD/xmGjA1v3U9g335VGk3ZVn6n8s9Ugw9jW94VcfMh8g5s7Kpq0X7Fg
K0O63GbYS+xSwZJ1HzIBjUDLieaN2PlHTI6x4xpDMfVrnO87mUgIMVVwgwL4ClqFQ1/VkkyODtS1
a1IIbKQSso/ak1n0voJ4/SlkHaHnSauVc6oeJ5wV7kWJ9re0H1Fj2Qyzstj5jpYFSl1G09NYt008
ka5UviFABOqbX3WXSQQ1mJjL/PbMGDoya3XEEp/7nvtS3Z2eJhAHoF55Zk9s7QL1K5Lzq10ZLOne
BjnbYjGxKDArZS8mJOOStloEz0UCdQuJ+9AL8p0gKwROlrZmt3lo22jLEL+jY+KioSp5POgAB4D0
K2KswrzvczyWsvsOfxsXZ8Z4O9gtW5rvgajA2j2WaeXvSaf6NoNQZ+aVSaFT0R8C/v06RHtOWEuv
hp0+sjN3QUkiIb/VP8FNk49VROjPeuvTzO5AUQ8fUE9VaStGrTN82RuTjQYmuHRRu7i0lLOp2rQ6
+0n0UoUydoGK0EZvE0/0mkIBhoewhJ1cpqeB49OSYSlI54mlD5qy+z7VnnCw7qjferPhJ4Ro2SYa
uUarjJkpgBKLjNDrTI9NS1JYULHHPH4OjkdCNV+yU8CVc1DQKWvrOYlRkGPdZSDkh8BZ1Tl0pKDQ
fBMyYK4u2GSUpgOlVipliqDNozjrmBw8sbHs5Ptzcw+x3LeYn3hyWdXmQj+Uj45eYuvd4pJqp1wC
XmL3R4eOjwbBWBR4Sz9b9q3hoo104fpSQsWQUn2Vp+441yzp6gFBeWHbOqeA3Bxh+uHoFoySLo27
D2NkiI7O5/G7s74vQWFZ3TAq+rRugoi8g2DGCEWmV1KNj/0/SRSA5+mLBbpJ7JEjO1CUa/F+E3Jr
kr462wkKMjIDjTLNJg7PGOKRQmxZRPL8NR5bxLy7VXXY2mBLJwOMoke8yw7pGv86m5BF92nlU6w6
eWH3GBJbCzaW9pzx7vZVe1kvGWjSsuQBXs2MynzZ7my6M/2RDChCoZr5CXaDNdxMQ6rM2dk5WYjn
AWVvO6SQ5W3enAKQhDApiGqVrwLiusGb7PSKYXwTdGTc4bGw3Gw/OTiIPS33ZydC2rbmCgF7p8JW
Mt8yn5Q87lD/FX9qaROiQKzSXpH3sHApf/9R3laxf+zRQ+xUH8hNQDzCaqhw3r7flYhfB9DRJw5Q
XyYdqsmb6SOcBSiV9vMfay3w/nyL8BxdrTP2Db5J0cqhrmChebHpu/i6qE6dt/sZx9H2auiojkdN
SeCJuf0CHr6SSTxUx8jLTc54yCi7YmmuJIg0oVDZtFc1Zsw1QQNP4DRsE87u0cIP+r4WnVBLLotk
YdZqaldF772Y/WvH193+xokrfCIW0FH8zyKzF1/iUg7rhSEyHNJbGPxtRUD7Keg3dZeKHK8bHM7W
YyiLRtnSW56UbxxDeYv8bRX9cEraphboDtQBakuNdG0P4UntBaG4sX558qkwbr4GzI6ZnO5nZTWX
KDL9SrKkLVoyti4WajSOllPBQDdSsHFLc8DgAmv65sZ2wiQJgu1HbQReLrkS/vhJa0jPAkPmPysh
7TS98d4q5zqOZur0DMyRb8dCHHTVW//MkKMK6GJpcaOkJ6zBFKjSDaqsTM9ynckvYMKugGigVrky
pkvEtz/+0Vzwo817pGNT9/MMDMKsPiSwvq3lJLFx7kOjqkU=
`protect end_protected

