

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DiIoz1dwiCymBJ2I1DU3O4UDdOCD1IYbLUI0voLUvMCBbKM/4INC61S/TdKSOoUevx63V7g+6/mZ
lHiHKW9CUA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o/flwcKffhg09UZzkz7gv/qZXGXaahpZlLeLvCPnGMHOV0tl8mkXW6lQBADTMwmBGUm7XZoObamg
kh0wsLz7sz0k84YCYY3YnDkU0s6XZ4yFdgj38M8k6+BTgeZETPuk8RfxBp2vQOv9zQhlLgklCWqU
H5aMJF7gqYDH9lzMxcc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3XDlc/RrM6J+fMEvhngyPf44nazd8NnlO+9fuAyN3g8+0X5quo1/68MLGc1czSBp+H9Wyu2aBKOJ
b7lFkbCJ13UBsZfTOKvBryDWOFa6KdkhYbTVSV9dfXRZ8PoouPNER1m+r+jF8e7EermzCIExWInF
5NIain6XV3z5eFAoF9+1wNHgh2DL91NQvcMqUhxodAC4EBuf80hcej88xks12032BecjB+B/gAMW
Fju2sqB0/mqHcdt7IfTqsGyFva1zLX5LMPhiF5YeiK1qj1zrDwFPgvhslJ9mmgozdcxNrfEp6yGo
skXdLgGuFnqjmzVIe1RLirf5OErXnL/7fcq65g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DYSqibotPAlt8I7+ZHxqG1W8t0MXnDrQyejnExd2/xGgdjHg+z1O251s8cO1MsyRynExFZebXN71
+rcOQqj1RiIoWzG/7+iJR/rcMh398jmqlJyWLU5IbIHCNoZyFsPrWxh/+WMiLYcvsaCPV1/bb8z+
2IY6rcDkaBrqk/EwYjE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
otEsDJz/b2bcmmVLOLfSwi5yawHEPe/YwdeYC6bj4QnDnh7iDtRlCB8Vxsd5V0BfHeL/WYjoeQM4
255fcpmsdbIm804UqNFTD5E3bD+pXsp5hjDUkd5BI6UEMxrdFYZ33Vo2q6da9Kuh+R1oMK735BRX
27ixqS9zhC9yoKM5h3EFDD4lGv1ah7oo8vFXQVvAoHLV46fz+yTbcdnzjY0CBY6ZcHBHkW/tXesi
gSqE+UJ05pdgmjP4NMP/1EbWm0c/tA0kZtZOMcSt52FHS77tvDYPPfsmt8s4x48hzc87BHtAtJLb
p2k4Bl3eRbmVYlntF4Wojcy6kk0ClpBDQDcHyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 32608)
`protect data_block
NG79Ikk+2K8IyborxUW4PfT2rfLUKyacS48/VIENi/ZgBYJnxgllj7dxk8qeUk3/Ybr+naqoABt3
aEmapgTEChbfku4PlHFunynziGfJg5zEeNH5M5G9TMBwLBqCobugvVf4spZAyDvcEseEK1dkJtKR
5mA9xK2HTjuyHyhR46j2WUTQKHLRoDIBKw0eKbht9CiBGUH6klDhfRXXIE6TCm8QkgB14wc2VayI
Ks0ngvj87LNJiuDNlVcNeu6L/PVfXn+QtTWfjHzrDAJlzFv7uS2rdrqSvb0rVfo6WtC1Ma1lqI7D
uJxokDl9wJpD6PnU6szqrJSvDqLjrIwQIJ7SMLg2sPNKKdJiAxv3NY9e8mBA1otYvXrmKzsgNBOc
I51jEHF0wk+YkHdJmhGibjlrwuV7yb+i9z39TO5b6KMxTyUDzwriHwddtdlAkWx7+dr4u075An96
sqQb59+wsuofYnWQDDBWLPRyjx+ScGWm++qPd7YJvS3HGDmMwWJUxihacbu6CNyN+Brh1aquR2H0
sN96EmyqgJFm18GxNUx88XPKS0TSkcQ27+basKkQo/JA9GMOoZsUhyufui651YBKYyW6AyybMALa
A7G1Sbeu20k3O45TYHo6hCYfsxwE1gIrl2VLZ2oD0OOiKuHN1ggnfmXyUQhKgB5nWlOATFldODW6
PQMxfQt6s4+riJxCE1MhyT8k5dipI9YxN2PDqPeYSThJ+HAGE/sjewYfO5b/JKgsUpWMf31SlxXt
kqtOCdkBWcN4KQ0hmzRYr1y9oE4rN6eIDHSg8ZwFpnBrZqMVxkXuL3DC4Gu+J97dZd0BBd0G1WIT
vSZkPvktt0uhNiiS7uidzH6trcITrkkdyCXzLfbCUMFaC4jQ6Pk8FH4EaLlCtpzRF3tATJ/UGep9
mZCKJjQeo6zrI9n8ADys00IeYFpmkR+/dGb+T1zx3FcF1Up1MxY2jMyYitJIZEeyKaowwrGYxTff
+e021dDpzHks/ZVh7fbn337A/C+G6w/soCFF5AHILjdx9Z8xA6nHAKwTwbN7tDJmVomySae4wZfG
/GnhRdMF0mEiwndN/ygVMvtTlJ+LboHomISyY4yd5zXLx2kpxSQVl9lTJtofHzKhUwYrLaUoMAFo
k2NhtxM0Qm+kE765Hl2LT9rptflfmjc3Vi8F+nKcqjhN3K4w7SBHDM0sw62UU7HsjssLjkJeWkU5
Fz+2Q+sgIrYYdJytOvGMfrDvXmv1q9wUmk6PW9x54wxYNis2HfVOTqF3w9DMs1TTCR63VnDk8Gio
h4GPd11z8Na+BG3cYWaJVdS7Q7hC+5XnKxfEji8WenO4wmntXiaD2nRM3+s2hZw5CiUGlMjrnytS
Vbns1y0wK72VZOQMCNQ1DtG9ma05eqJDUK8s0hOdbySJGH+Tw0oswEywlm9gnjLHuGfAkJKIOIXn
QoFMDVUoQxW7KOExjEfHzO6Y6mfmnkmLfXSRSKHqdipQWG+VSukywFGxOmgDyUe/YR4Yq31mJXXX
XVm1Vtk3V7HEKvN9PwFdeRy4e1tIvKlSJvRghGHHq2GlB3wFAzgScERhnSFjNOYQH1vT/eYRmNx0
NvIaSFHcNPDRZP3zP93KeOftbm7wQ8nl00ZiziYJx2AJnJVIFNAkcFhqiP+8//rpJslaqLOUa1Nd
GfCBZWXXLZlTU75RSJKy8M9hxGhofv07vcJTeLJ0MlOD9c7FKC0f1njoOjOhI8ONRMPRvndj2GR/
53UZ6M6baKcVhfPYEVbx+QwJhti1VKRibHc5/KRCC91AnWidpMEcqGod2lP0UeW2jKBZ7qHKxp69
fhXeMfbxLukakTeiP9CYospetTBDoo39IlWarfvt5eUWIyu7N4lj7BnvUNKc2TYlWLltN7HFsPV5
qCf24zQR8StC9icbUnL5uRX9mG+zkvol+axq+wRbgotVs+VNAlBrN+q6zQ68dxmkTB8M7u7kmYKW
aklN8fRawqQe+nk4delnjiHjbcfQIL2OinihYmCe6WXtRelhl2WMLiuSrbMwqD1wXQGCy3RhwXDz
WFVippx79wEo7NhQgNfiJBwnlHD+sOh4QUHUOiwLrp57MkYZpdhz8UkzoaFoZhonFrd/hTZ2MkrG
gLr5rAFv2Ko3br36EMHqn9ttl9EpBbBYHwCDjRTelWXXsV1H8WoFFTQSPmV+Kmkgeiu4WEEzVecQ
xw0bldNnMEJ9dgVLTlxo9EgMERa55l813Ft9ief2aULruYgkNGU2YWDmRDc48BYt4lqXO2Er7eXh
lgIrAYKxO39T/yb3EulqEX4UrtWccl54VMbWwOU8SnV1LTdNMpoovEGvlPgJCLRv2KXAWFq00jLv
g0t+EMpC60v4+xPXbXUyQX8nQbr7YSuZ0/jIP8suBnfs2V52aokVBcw/A3oBU6GmXU2Z/HWjNKkc
Ufn9xYQTCkpjk5y2XynmGQMTvvbEtZH9OjFy/7o95je5kmqfk2qcjpjV/Jr2BXCI5hjEiH8jTdns
4Ag0/gppsP7n63YwTIgexC5EnFv4TLunmmc51XQ+Qk62D8PGe3MTA2/0BTftGCBryEOOqfqmB8P0
9CCBoS1qcC6bNB4I7Acve+CQgJQtPVjZD+th6Dkjmij9XsykBhcWth+nv+IPuSiKTfyKpa2jsz1C
VOXU5rBJsSMG9okGlYozlIov6nDftjjsHdz7ESSsRuac0XMlx+OayJpMAbOso0M9uKGw0/8BRKRA
7zRX/16tmhoBOQ4zYgH5+S18oeLjLmT+4PMKmrZA2s+bXjAezqT/fFmqm44lYGwvXrAGs/P5RWfW
Ol08o9rybPl0pQbzfUcEbZVssWYwwWRjDd5bVZR5g1fovCGYhZZ8UcjdfaCcN9q8UtscGaDcqXvh
JCiHEu10cojgbo35VyhG8pHO8LXkoD2oMIiSoHo1fhRmzQ4Sf6Rr7X2kKHuccbDc4cYLtdy5mGR3
B0Pfcj+sB8aH2zvpeqz35fllP+M3uOlX00deE3ZUfDMoe44sNBKXh0GZ64Q0b43/3L2fbKS3mWJs
E9JhfKBH72p6N8do4ve8dpidKJ4hX/rfzOsCpPUtEsERNPMD/5IaWTUy4nLQjL9g4DILyq/+aKSc
14Gbi7OyVaBX5XmfL9nXJBcmK2jAbvDflwqHnATi46k9wpWNT+YKzdYqLIEFDnAcIlbzc6WeTsR2
pMeyp7tNb5JGefMk81M1Bdp307GFeJfeQV7FETzymUSBQ1EixNHYPI18HS1SeLmKMiMz6AUBkrvw
+2klNv/z1R6s+YuZpUGwtBWJFJ4Bguk3YefN57z6dghjpOBN6B0KYbnGpTKs7alXnr344vRFHo9W
0Hxky43G/drWq8kVcx+WbITr4F2RmYpaM27O5a5xpMcF9zYKh52LIL8MSNocZrNQBe6gw2qDPra9
yH8c4RqD3Wx+uAb6Y9J+HZ77MpD3O5H+RiuMS4ykWOyk1vARoQVT4V1Ih4d64FLS9G/w7rqHu7vY
YO3jmP3tULV8Dgse5bIr+SaAE5+ClET8/rXaDLpkonb0dqmWqbiXgmbw0VhxC4EbOqbLuoX5xYQQ
E+xq+DaBbiGgLjT5zVZYybyKJGWfgK/vPpQzirzj1oo+L9gKUA+wr87XQNLQzvahkmYvkkqd17Mu
rDFkuE87OuV0+24NCb9/m9uROv3orpzpVI1ZvVaEWS7BrhbmVBgQhWVbZ6Edvxlb80xMuf1UreFb
JDhBBbEAfOIwuHutaC6C+ra8I+5fW5yuX5dCH/ErE6O78abx76Bcbw/VWkx7nLeOGKo+/2jr7whX
ZGGiWjx4BhEJOdIe2uPUUhjK+JOAX20aQHJBw94EF+IWFLiQuQWGiY9GnkbLdAg2GQXLJzaD2bpP
hRlEtOjLikVg3Rre3W+QETeM9WXGf0eP43EDWKBWRMln1oAZ29gAXq2XcDOJ8s7uC43FX0W39Stx
zTISr4Wv92d+eopGS5yl+HonkjOAlOoDoIXPWKqxAoeCZRdudV9FOfK5C2BEMegddsC6LJfw/VKj
uTS61OCkg7S0OxQfddFFgG5/npIWT9bt6s67YqcAoYe1kG839A5amBTgdJ7T2yC01tX/KtX4BTDQ
4A7pRqlhBZTz4IWAOe+GbNPclDhbBDJE/x2HG0CICqHfz9Qhis0cH0I9boCo6Cph7yZDvAwoWVai
P0rP/42/xu+GFMcXuDQUPpblNMGp8ZkIsdbokmBPj7TD1mIyAgO+U9LEqMBdSMSpkLdWkMQgtCxS
oVW7OZKMGWWCK1tyaOm2mKFhQQjZQLeppJAR2QzUDJSDCgnLq8daHi5im0mgtKQ4t7/4sQUySp8j
5wdi2RZRKzDAll2JMRahOemwQeZj6oXI9JGhA8dEIPPHrnwLXMOQ/LAcq8o/W6fRAw7NlMBst4/y
NoEADhjs1hTRsXqdOdjNC6TExhKCxtc46rggJc2+TobkBflyiDAMCfRDlpAKJro3UT41Eiy1pkMq
BKHhuRcXWrMT+575QrkzTHXkvDwGse7AfbDgcYQ4asRVAGgPGkBkx1nm86jruMB9mMUe4jg2eGWH
Hir5t3pDFxQGfsO4aW4F6D3ywLTf+hPCqJh5q/FFR72ID6Co8OBPvd1GejhXRq8ppgrEg8KAAx7Z
UVEbi5a6oVXQLUzIxNkGGCNYBS4O9K2zYFqW2VaZo8Zif2UyE9GCjkvUIK/4KZ8xoWTtiX0Y/+IK
Ay96HMcnK85Ru0xGPSeMJLmrsZqfemaI8qtuZIIZJeskyK0E4E6uh8iak5hcXacN0qIhmoxDAKo4
kxEjTKF/zKx+N3CyiPzHRNP0Uxsb0VQrWPFdbjGXWWqazQAnqmAu6QcPce8CBTh8cFBSnl8lS086
mYqQUMaOePv2thzzsT0UUQ7BPZ/8RuirKckj/AA5VoAzGW7r8isYlQJqIxPw6oyhQePC6K1MYaDe
okySwzW1uLzUqsTQbFLPaEmm+PxpXgNLRRlkXAI/dWci+EiGg0+b4A+wGqwCSbfH6t50AKbFDwi4
zTPuAGd1jk4YTA6xHNebbllslPHY/NpvwMluxGPa0JoH2dWeaaUORRZwO6gdbYDa8G6WFLAvhvlg
rNaRFuAlLWfYawr5WNIN7nLNz884utJpnY9OAyfpg7nWfwpt9U5TEgdnUxArs77u32rumt5hUCrE
jb7/OAQUSTUg8vJQ1/+H3y7VD6HLbLV3CN3D3/23NObI6aMtjqkgCVvxw3fwQ3aBgS7noCWCc+q+
0z6Pkifs0raEOhRQj9bNt+SgNo5MjoWuP1O+gmvGUzF1LtyghZdfJGmkIKubv1LrJbmd6TXw9k/y
aR6+cfUKwMuUHV1nXTNdsMnR3bDAeUVnmUywJQhCrSohwhipv07FLYztongHFVbeDOPyjHw3tFAP
tZN5PztmsfrkQUf2xaQ73MqFpGNgG7sd63LecNAWERLVsInDG5Uc/olAiROY6G6pdPb5mNnvkVio
rN0VD0lzP7Z4RMhO8IBDNkqbzg2KuoxhVK87NFwVvmwmcd+nks1kTarC0jymmADGW0Yuzs6n9LHS
I+Gx+3QcPPA3gHdf7UJp/kOc9aVJbMPf06jb28SfKb7b/pa+WXsmIwd4odSQocHvCxFkH7AQBojr
lhIk7VZdUwrgd4H0TZwclBIbcNjXO90osGnNVLo/uyvYZ1YwxIGMOj6viqlN391T0KfLxyds8DCL
JuDHLnSeuE76p+BHUa1Y15fqkZ6uQ5uoUlEO9zglNxwKoikzIhVxp5/RI69+9i6vkl0uKkWxXBkO
5lFy16nfWEOZYGkEQLP2+tq5Rj2u5vTWa4eUVpydWqe3OQh8KdHkh6GEhtb5zksVqd/LzFXSp5sA
NwoCUMadW+MSuldKkyA3ftpmabkdhqn7geXUS+mE7+9DeKuNK4ddFUBMOK1cHOcAG5WFxd8Fos+t
hXHzHtHTDCioHJfx/DLBtdmqY671nc6Tn7O6TCEGy+qhBedGWadQOCEKXhuB+/VWWAvh03N+ai9e
ArLWebroRddzntU31VjDpxYdu9qcKKqm6kYYNdOJE33mEVMOfPP2svMK6fi/Kcjyoo532UKkcwFb
6DSHLpMXN8dWUd2Rj7+7BqEaxtNruInphxjzwIWd9bCJ2VGN7n+nvHLccAtfyr0DFl7oakn+Xhuq
ZS5Huy3gmwBlaMA5r7kPvovxO6QN3kJYYYq5Wmnl9br4mD5PUn9ecJ6kSIY05qiAmQhXGl7+QroJ
xHZ19ilSCWhVx8JIQlyCbgqN9gQW4jxegnCINn2RLmmbH0eUE9mYmBpVTGy5QJouJY3mNOfZxvsk
E3mDVQGBcGvm4o7eaD4T0KMDzkxqEunR//zITihgXsLrwS9SP+ghEkhgYlKHh5SLFGSeI9Zmdh67
Ar794bY+lqmosoDxUoKM+wF8pJIdfGsoH12PACVsALRslVW7NT/tnWPDCkIvFoMUHXvygn5Txi8n
XblTgt1mfKDeWp9RQ+yGubrLU2uYafJ5P+aC0ZYmzWACs1Lm/ZU/F4UjMfl/yVT4XB40D/Ukcx8f
ou7rymQ391+pb5b+gGPEUmXgoe+lK7iMcG3d3JDiZoNtvDu2bpydi++mYZjIzugQsy8+F8F8pLx6
3lZvStNCPbxKr+A5bGXaJ7i5uZzvrYjv2PeoPh4JUorzPduWOYUMYBbWc+efKij31RjGip7OaXO/
jFKSeZipbHBcqagPUzft4AQrnT7X5EoKhldfxCGT3xi7f3hvEJCsvHqQ/vLpcp4h6PBRC1pqd726
TSRSAN9ySFYUUhUuZOULlhDk6Bk6CQVmthDKolQ6QRuVZPGP+c8xHNl0IzdQEfGvpA5IXihMTNd5
W3Qs8nP9+dXIeTTVHnTMbkNPOT/IL5LvDD9xVnzwk2bT3H3q26VHwSPG76kriPIYGOEFkQCBexQj
gHf4mo6Xqu8bOukU5A3kzArW5VQxOJGpc1WUHnS0pKISeiUkqZkBkztAvogv7tTQ0XeWIylSrmj4
jABeooGC1kKukTOozhy1yQmJx8lTODtcq8J6lEpo4cIR9levVbMp4hSdNMABx+LoOF7jMeglJO6F
K9VbW+Rh3gXoJIndc58zmu5yfIuWCTNh85Fwo5O/LjJXvZGM6PfzATmq+GXyvtN37j7jwih7qvDw
HmPEJXqmn5X5etyefu1iRrrs2wR10vUqXLLApe5c9PFNkZlVUf/JUWjBrCdtQSaGmJXJHxWX8wLb
DZRkgEfClImPHwmLR3s7cfkgAUV6MVll8o4EehdRXGO/qQzxnUwcywa226YFuPkcqUsinU3M11FZ
ad8Fhu8PwQmaRQnZ5YOml7TXHy6tcQ1xBzHO7PWe5MgJ0h4vm72KJL9Epp6gzw1MgXhHhEPngJ4i
b8SmRI6094FXX5t518tbq3yN5kCnrX1PY12vboMgDQx/JP70PKlGvyb18WC1IcOn/qBVuMe1+6xg
iBFb/6T88W9VIlXJ1XpUuj6/O0DHbPvKI7V2NNPuag0jFQFqqPE0wUkxTOF+KxYk7aLpwKIc3iAE
02oiWHuCjGCuVWq1QLXuM1w8uEnA4vFCh57feTDTzvebfuLtRzXu9yTjSiQ8CIfVFuveCU2n+YOD
yFp7bCxUSyuM5bucVqd2W89e6z1HKFn0myuc9DyHpYND7seloAnL4Ms9xeeBkZ8E8J2LaiCUUqXM
je3h0CEgFlXXBnSVYp45yEe7YICpuUA0k541hZGx620ISVT19yvtwOzQJOF65MThT7nggGWKcGHB
HVUSybYfmmMgTQ39KvMxprY26iLbkL5GNYDzCZVnMqdlQR/7DYqRM1xtGnza/zNLEBKD2zY6hWdK
3hOFSdWusa+KtX+/Zg4NA+HW28T6AS/pnZaFXhmDg4GpZsAOF5Kd8pUDTPjQ1QcfHGldSq81Aopz
i1NZFHjVLUocqjZ9zOuzKL0kzQvkDTeWlOLcAG4L7B/AJWOoQT7ByqwikyJqPWfXru28CF/BZ1AH
CC6N2XJFxbVlDfwoUxhRG7t8oq34dXkwOKYnrQxGbsJwAIdioXdyH6khGE7Z03oI4PKYHkkod4gJ
kXjqpDlsfXous9hghvSXae/NlBluEC/Z0lgxspyB3kpbqym+LhBrxpIA47munhEYWDvpijbNnpKE
/+TRBpRuJBoqeu/CsjDsLA/M00VjfnA18ngujqgbaizlJ06L+bYrWGYVLdktEf0ji9CEorGU0QXe
9wYZ+YTB+deuK6gbmMaaXH6UDtFFbOfflyrYJZ3j1P8uRUCmukK4+kB4sV89WkfUcrtkMYK9bUsi
nfH+kwqJCqGLBntKuM8dRXTuNY0eAhBt3ohh32adzpLQpZycZzscfuHWI0YFrt8zmvNzcgsuiTAf
2ZLXcXBD24H9b/jAYfnu/KECbIuvP0w20O0B8jBF2IFJaE0hFEFA9CXRlnInj+vFVcw+lfVsuk1a
Q0w35RiIV4Otmv0J6Q/nVhXBp0BVBeNeRpFvufQ6W9BLUHTG6owNI5b7fqmNdM+jppjhgV1uAlGU
i3HQjFVjrwcQTI4OmNGX4SL5SqELwf2/rxuJ0qV7KJKTK0KBT7F4LfZ8dQnC3Ub0kr4uF7Gzanba
KIpd1t4hFG/cDetLXz3eQTyM0DXQ57Ff836fnpMfczsG3bl15Ix4aFitxfIRVCjaCt2U9SPMqM/l
LvSTFcw14NsKW9aG9oNMjQkrV9h5HWjVZC0yoB2BSkTXHJlU8Kv03pcywLLvJc7Pf3AtHEW3mUDM
1tEIYnoMB2j7yeZT+XXHYNJmevSsCt1DllKZgMLOx3lqmzOCSuaBC9ZaflT8Ym/s1pjEIjALH2x1
kkTlThz2/nkvWRbLbXoY6LY2fBEWn9G5q8gCgj5+CA9TzjzlVlgoRtT36V768QhKe96N+xzK+3bO
yNZGTZkdZLPFsaH85IIfzdW+vj9L6R92lr2yhtY945Tsa4hMh3KaO/kTUSGtilH7e+Egf5mkn5uz
3JNm+8yhVAR9wlCoc54tRTx/nLOwdjLzUcxCZwyzq1PuTObZBvs/DU4aooGpdDfg+NWPQyRHsVok
UEYsvkBQ/XdbQ0d9SrYekadW66u0jprOx7VT1bYgO6b7IHDlfieo2Cn0smkNEQy9Cjdp2k7ayzD5
EhYmgWAIOSL41oJE2jSQmxpqijJ1Iyb/+Wtk0neHSVlKJQaTy6AsKy4+bEsgyJeF/IC7HRSwbGhD
d56LjZJsiUmFsEfgTQiX9f1CGtPQbCUsMW9k43FxtiQS/yxfZBD7AWWMDLue9Ux3sLdzggYcf+50
JMAc3pFrXoxbC2s34cdlMqI2BTZjB1HLKPohBWXBdlR9cgBC7bfQxoQ3y+TUrR7AhbJN6QSqiMHv
I+/B8DpqWtT7Vz8nExwG8kO/qH78Akc+BId9OdX10OWwyahz/d7S8UrVXq1bvshNf7qqoBbr5iNg
SwOOn96sTghX5/+xpLkE8pVr05nKEfPYeo9+fnnmuFFGmi+oYrbn8JWP2NdUOlVIQe6VLpZLhC1U
mzXMdHuztyrwc374xNGBIo3taTlPuOTce34RBSUt37GgOvHQh8Y0aC5oaYvd26sPYZ1i3MD9LKMN
HhBBd5tYVAKU4Avhztl5e4JuNQ1YQxxH9KOfup37NpzN5sGWV9xNUd1R774Irdb5ayIVzpwNyTkg
V0d/6aWwhBSDb/Ey4evmNmPmzzPIQje4pQOJhqnxDtaNUdCteGGp6zNukirV9yxqVBjQ84+gWa14
D369+9J9Qmq60RusotbythLAe8nDgaKvogZH3PJafah8/8nvRBpgQ4LPyg6VyG9p3AnMNT7trsYX
LKJ7ckxmcsdRO/uOcKpaURtSy//FacXE64umUWjCoaXD0j6NUBcKqVmAnPuweM/IJtdxNBtn2Bk0
YrZ2/zCRE64S9Q4EUy3Y63rEOqHSj/VZsg7GaEZOw4Wgy4FnfRBWW4YGcZ1ZP15oHF6mda1ZBR48
pjwx/hEVAH7AMO876KnPb8z7/OBg69Uk6satTTsq7FAI2PFHUrLQ1JDOjIZa+uK5o1HVyb2CPOAw
AS0rD1qGJdGpRmC0qgKZXkgo0aKU986yEKBpuEDS0jJASlEOP/URQ9kzLM6cXdFaTjo+bPfeCBEl
EyDNPLWF9eqOt4j5EQi2XOUu/pSy+YIg40T8Lfa38bFRYp9MCE2e9mFXRYx3MqIHjPq/wreLpRVY
QdV15UV2WLN3RK0fLtN7nOYZQNox0L7LSduzrlDfmqBUGPNUnZcKSze4ocStlvvd+oauT+YKtGgA
1WV9InNjEpAJmacArbejhsL3e+r0V0uAcpLolPrm0vg4pGVT0trXqq1glwxYS/lt6/OAyLWaJeUi
1Wsfaq+hSgKDevIY8Vnfxmy+iE9cm4IZnsPJU/LBqok+S5E7Rzl3XbPlkbl1Zd2cgZHe0KlaWDPk
6q+BPjy4a9Es4+kaNIe6OCV7ByG5G1XNcaQQWve/zJsi13giiw0gPUCmYVzGG+pbmzQ1+mozlnOo
JK1N67q+2KhlJOzw8bOkUXMLLVjEMJX5zMeZHMk8BmcOqqcM6lQQWtnve0NUrMoG1BrZpy52Nem7
6BptOMrPl7fD5RLnhZD8OO+58szJA2ZEDMPcnhXOiFfwpR6DqjR0YJbTHbJ0oX70y1lvIZk5Wnin
0pjeyMm0W+qT549Y9qdHB5nlebBp0za0s6GNCxYReigUAfnLlliQu/ha0W8lENPIO5vaxi3vdd78
4G7nWoIZukVz0QjS2XcyABuB+0VDd8Zqvm6pn79PClAO8OxV3lLhu6myJKpVvEx6z+9zj+pt//5z
o9/Rq30lGwEZhp8I19F2Nr8xtBkcj4JDWWZbPEelmBfgzYbKf4N+3IBIC0/Th6Ew1c4QRFD2FnI8
K8xZdzJtCt8OZBba+0qnhXrj3BISI3bkFjzF2syDt39EFCa8KiCeMflmmhLXN5+LCaza8+Lhmn5a
EECaILqJYMKqARhkD4AVgYG2DMB7xZw3LffSVYA/JZEz6iFFD5gZ2V63oeFDPXWSGTHkTh+8MlLi
bQnP+1IHUaCETEUQnZs+B9FCXDiEx6Ck9bXFgVFI7/d/qWF0alQGq0MSmOBUsAQ7lyX7e1Razq3w
tOW8ilrTRzRCY6H9ZLp7DSdcUsHSio299NNwQ1JWUK52t4RqV24PRuALpId8HGM96KW8ljuJOY4I
MwbZzwApXMTRmDH/os38FpCkoGCw7ql5BIfZcBdBWC6AOCcvHR6SWlilHAt75XfBoayd5P38cf/p
kGmOgypWAkojAy4enZCwGsOF27zcOBixMgqFwH2+ihHUw1qi8Z1BCY6SIWvDmLMQki1tEM95azjk
2HnXufCPTJFTWy5Bm/+SUwvY95dAoI6SWa9vdBiY/P2Yz8gw2tOX3S7F8B42AMjzk82RALKa+1jH
GiBvhrSbTlCA/6vkPWWiU17jR73LSKP47LIcdHhd25ApY3I88yqz/seDCcdPAUf8XYaJsVnauIQp
JwduC1dETYHgug9nhoh1/EEhMqZGGGxzHNuqM4nls7YbwkaG6RCR2EnSralLEjvWvM/LB9f8VQy6
A1/DhwAc8h+CNve8L2rovc8oaP3zkqHIld1mz0JKpyT9mZkYdJT+Na7m5KiRiOiJTIFcukDUVXIP
MJ5NjeboP1RsYNlwkiZYg6yUnTi46OfLeENojv/KidDPZKCKAtdspuC9jUJ3cFeiybPYNAAX6t39
J+7R/gsj0fBptbZLI5+eoGpUejcaLyeVxdhiZnsIUUz4sdfRgTB4XPMFT9t8+cnJdzxfcImMsinq
LR1gNHGM+T0YSwK5jE2sbBPKZqJNy9k2A6MSIPA+7B8F0W3vKPnStMfFhtNLyrAC32Lbg2DLDUSl
3h0mddlZSTcvwC2W+G/dY6c2dj3I3F1vAdJqEz8P7Vrqzh0mkayuRKE1QbWDTomN85G8Sy168Gq2
+hN53W3vz9Yi80O4pZOPPrWmKHskpYmRk2uQPd7toOv5xyH7KD4sTAGv4EZ/ECbWOovscCvYh+eA
Mu47d0d1e9CZ6spw4yUsHZZ5bLqWPOsZNoFy9a80OzkHvXOs7HS8T9qYrRVKsgUI6kW9ZFtR/ACc
twPGMI2Q12MYt7APluC4qG2NHW2AdouSIptYFca1LUvTs4W+1gWTAQNj9L+lqyUZ9/GvEP9Ql7wh
8AWLhN/WDn2E4KK3YJrwcYR5TIDCfo0wOepRAJh2N4VHVFbcFr5tEdn8GW1jxjh3fuSQQZksIyXX
xLlxK7nLQcZ4Qc4Mrnt6FLfwNxIoGMd8QyQcG4ZnNGWIKkDNWOV/p9I034VV3XkTc6fqmKulQwgo
8F02a91Fjsumq8/Zu9Ue2z92+gL31twfmtDsUn+iOBci1hcGgxYaFvJo2yqLZpGvsUj5Bpt2Q9OP
lvsaQEMcCZbhko4xOg2uY3pk69/+9g8I69m/5RZMjlNdhv3EYXqzRXLzOTe+erc4bfnmhPApDDOr
fghmgT69lESIKeu1sqZqUUZTJ67006XeMIofcOdF9bAi0LXz47PHoqhnwxnCP0v4r+lek4hFbQE3
tFi+hCHPvzIu4FlSAJXX7R+n2IJrIkpI8uLndqKWV26iY4rVDoqaQ+oOXzWqvkp4wWlDjcpPcgN1
VD0w6Eyjvl9xmAHdlIY0T7RItbiZd9ZMBExUbnPtHH5yW3NVQXBba13jCtJvjOeh6ihqoCsbmlYd
RnVg2eUeSO5EBqRQGmFS2f180Vh8ABbfVdaBk81sp1ozvUYSNLLN0BJ1DLLdq4ZSB9+EGQxQ0ODB
4y04okCBmUk9118IdlrI25oXOa1sWZKxcxl8gVB/W69tQdLeo+Tys6+H9JVyypj5+cT2OmfVRatz
PMNmHrjxP9G10f1OE0aRY8SdCIjBogk8IL1EmnrjAgSTcRpcj30HODwhordbQwZe117RReR7ywAV
KlHArNeHGsHoVmsEvuypxPGBzv2LUY/OrC1qPFdLYEN5dNUH/+pO3uC56bn6QJBfTOpG3+0RJ/0r
oy1qm2XccuCh6M8eD1J+agLD2YFATgEvp+JJnGC/oPIhlnGU5qAuSXAb4BNAjU9Tbj0pXFT8WZmQ
IT9mQznVnRuPM5yeLmvMXlhV0yqOn1HuwaPhSSyJpFO51Abs1DV4tYkXVhdGsLrD7HPTYmPOTs/X
lGZQTX2Y22pMOt4ZD5gSpJvYUWl95bjturxp9W0uo4dL3rooTzZNE5JAu/Ayyv7P0Y8cOrJxg8wQ
usyrXNe1oDxihN+KL/DwLGt2nkTRr36qzU7sjDk1WwH+7vMkrsgQl4wEGXdck/6QHkpLbr0GP274
CVJBMLDL8gB4i1Oo6Uco4aUIJIMqwa+JJ6dJAj+y6bT2sKSlaevcEwdPc7DWxFMDJxK/eUwdpTBv
OnINF0yoGHGdQkHkPkpSXduX0u4p0OR7eEqzDm2kVBXy0ZwfQHRMZs5m6bitsMuVcwuo5Mb/9Qwl
TxLPs0Phm06+ZRQB+ev3mC+KLxzCMm/e80DgPkv5Dz+K/rkuPR6eDlG8btUPulotfEgEnX5xNjRp
PQW79dNNz7NgRAaDkZ1D7oQ3Pj2/pQCgOr07RztqejuDIrkiEpE05Dne5OCGYnV6U4FSCupWDLbU
QLyKSKbia1PNBBH2vQmtbR9yMskxOFopCXR/L/mIiAYwhRAJ1uutoI1XNm/AwjA/Iyi/WQzyI8Zl
gnUD+brLxRXG0VJpWdX0zDcfr2poUp6Y79PAHTtvpb2xqw+vE7JUXzf9CDc8l8JIMDV76aqcl9Dc
BI37WCDUR2txbUkc8iyPnBhtBiUNMpCnGLrmW1/VfPKQbbQQkJiNtUaTdQ+gV/j9M6bnZGtg0gWe
5gWytauxnjzcP1O0ACz0IXhq09JGxRaJhKaCKCJxarQ9N7K1MzJFlmVgEQj+/XIWW8zeS0si6097
y2RpCHhmIRRZZ/mHG090VPvXCzpzejGWh+lCfP9iPTIWf4tqi1oRKeBdxqpL2Z0xEdbaGVYlX4gS
wM0qiFZCz8o89nb95DcZPiexdxkH4928KCgt2bf1NdMJJmzMjYBXUaRxrr3Rc4enosIhaEYc5bdX
rqbP8zsAAvwt7VdIJYT2ygDboTZBlM38xn13O08Hq/+RIItEAUJ7CwMYkezzvnodHzfhPBnmSQAS
LuZjaQNdQ4LWttWHVRcnW00pgizoVBOWjkCtjSZnTNOyjb/zrQWrjd0Y6nXMMPGz9CQoIcctjGRM
c8d6pb6VFyg+Ef+JoH8JczLn6t+sGtuX8qfpjmozfLUkvkG39w6aDkdH9PWBS0BEPLd33Aur/lh4
2VBj0eBAtXxWsomkRADAbtOezjEhTBKwICK9MoluszoAbEpFcgfTG1cz73L8++NQXkxuOnLsEfUG
DUcAl9dry0Mklf2vF+9pjPLp5Juw7NY7EyVGfNiyvvY57Gwn8l19NQyxzrpLAvqV2z+JUf11srW/
qYB/vHz++MdSal2d1YXUUsxFfXcU5EGUWcuQ80ZXYmkdrNiawceG2okO7yrUq3/xeqX+e3nNWbCZ
PnN3kg4CoXmtueTKKjKPWfDP6Lam4dQxqPFh+i1i4UWbguIHZyQ79tJj7U4D+TG4dOvvLKFq3iNT
sE0K65mHFG92mGTRea/zFIXq1QB7VuYZcudlfi0cfpAnYVKvN9PnKAyaA47nFCOOvOY4y9oom7PS
vdXMDFBKViuaBmiEcfxBsk48AW1Dm5RucGPbYxiyjbEpZzhRUtQsJDhNtcDScUEVUmz+eHJZ3NX4
5HzXAtkjlLzhzGR/qpRdsYmLPScU2gyieRqQAD36HdR0ZsZjJDTSKVR+q+nfpwEcfKzQZ9hHSSPf
62RSjJ5KVmXgSzZ85T4KqUXoihPfA3ibjxqRQzGIN5NApPP6njW8500QY+Qbq9vyXVbBFlwMOoEA
dmuEHMUua6/wPrGY4KfRfXxPy2Vza7Rp+tJqdoBvdXwTfx96b5TINLssAY9MZWkduGV5pILod3cN
qIs650DwsGigoTmxZxwjAsV6vo91XLLYS4xFIb1o/jt47RQIDI9gyOYdg6NhsFmmsW9edkn5rvm4
6UKUsHyONKZo/8IxEVWGcwJNHiw6UWivrs2dZiyQtIzUiYaToKeEggPdX6EuKYIx5RNGX8t4VOfR
XD3p5S5IOMUkl0JXTI8BPURSFblZ+/Zg8EXXJrA5N4jf+1BQmH7cu8+pp2HDFRfLpKojj4JTocEy
puvUxD4LskYL9JKluXSVn0Q4hfJlhD6CwVDiuwmLPgCRfo1IdDXuSpd7a5cNJlbScwKdtUW7MihK
YVqxhTWoYcH0ABHB3b78NECmsf3VSimt0g8s8U5BNVSbrQJTx4OoucWubFIHL4K6iGk8uZje/zi8
0f7+Zh78eGkxu5NzFFI3vQaG724yWPdxyehQW1ZteA5VfVgh2lxPCjJMNn3YJffsRJUKql0eeTCJ
urOLg3CMEKMDrdJ5L0jdJHEXlwhxQJvRYk75p2kBUJCUmKHqm1bAGKTc87DndYGbV9Kn4945/EID
b2nv28Nfb3xZTr/41oFgTfQOoDwI62B54B8elZQwCSRKZ010KOHKDOyGB1S11JxSBjzk9bh39VBr
T6XjAA6OfIT6mjGDcll0j+BLr0jF/Cfw9YZZFcmWg7Bw6huJeknMMIYWjsFJr4Kqx8576ZHUTCJ5
eTycv8PXd8yvsh66S7McrNb99bGGJSwhJX8TYL2ZtKJ7TRy3c1kRvRTK0KoS8Wk2GxzRLLOA3ppR
MpCBsCUXSAycKh3wtFz74Y47dEnCKat/Jft6sW1UNARDpFsgEinlb/V71NSN1cNvBgWvK5PI2Byx
ShHVAtFfOJoqALFRYVywi13Dm4rM+RlP9RHY6ZOjG/OMxA272f7Ig62myEVk2RluXXParxBkTBFf
H/vlKM2jBJTXQka/AV2m96YY18kS3lfZGpQd0j6k3leBfr9cbI/sEID8XRV++k+ELPKRtHrEBtle
y8+WcuHEVzQ48JC9qOW+rZtbO0jpMbFE5CHu7TO9gQwR2CjeHIH4Tlsr+B9ERnCVvF3F7+BhLDnB
fKNxR8RmwaKP61Ik5WsBSRuDQB3/COyCtcxeNKDIsh3cPhvs4uoH64cshG0g3eNVi6QsJHHMqj6y
hHlQjfbLFFLuTIV/BC0SejiFs2HunE8zLp5bENRxMruBh0me91XR2oCz4zyWL/wiiY7g9UqL5zOr
kDDy4JPNr/6f3UAHJ5g9aI/Pm190JLxrz2zPcZa8yFKI0zRTw0dQBltBAKKYMILmfBBPFurI7v6s
Y2x1WOWbFQZk4QZ8ZDRRWRl+LzBrwFSwvwFmkLLCghxMx1LgB2fZEknjtu5Q0AcfkHhte9ggASKe
XuZRwdMLic5ZPWEK3FapeuhFAuplVqkIigfkNOM0ktEWfLufVmXn2LPyqagQLjmxF8Edgvxv5Klv
zigNAcJXU7jiDKD51WzElIQwoFyEtiDCdBdYD5nJx/ZJ8QMVB6+jXWpkxIa3+InfvIhEnjkOd6U6
cIdu6ndoA34embmE0UBr2c9MWd1ilJGW3CdUvpqMmje+AL2rY8LqLd0W4P3nS+SnGqAm083MUue8
0VFhF5pto8gHsnpjOUfSSYbLZl/8jvUOZ8PYSpUzyHM8qCAnejSXLKxznJBHQt93HBTd62VsUuq/
QXxbLP5rLlmSpb75vUvq7qxN9CZLutTtyZuwf6qcaqnfQA1bvJ5aWBFNB8Doc+JKTAVl7bCMQywG
aJtoseE9BGtuXVJoWRv/zSk96vfPW6/jZzivmQ6jPSAZqnn9dnzUzdcAlNfTc5DNcj5Uy0dlvKho
6Va7U0SWjJEiIB35J+gIuT5g0JZtQbS0AC3BGnfXxXHbClUHqx3Flbg0lnx165l2NQm2Z8hrdOa+
JjuPfpGKlGXEWDvdf2LAdmV6eJAfNNKoNnm4Gb0uwJbR3ZuHK8E8V9wxOIp7RrsuD8IiK0InpjI9
XLf1F0ayJ2xaLPAfIPUPK1VrMsIrfgpKosr6cbSeSWSmMfV06V8APWcqS3+GHIsHTb+jrwp+14oH
HXi2j4eC6czP4JAcQ/qr/f75JNFfYRnF78GFJhTrNrsdHLPqlRSfvkFblIhMjVcR9q8ZfEE1QtdO
S0og12yMOZgJrDKR8kNXEOd1VWuq6o1D+zMXhJtBaiYqdSLhgXwc56KwocPJEqJ1JxWExs6haHdh
+mC0Vu4a0wc2lUmjUIVGsUAuLoZgL86d9qrsZFttK4Jf2+BEb/M7/bt4Z3t9cIOFhzyWRsOfqo3j
3LIj2Ubn71PZy6ClElSHeqpKwr4H3Ehln5KEY1jdL+F4lTyR1sPjWRsnVVlhWxubQwDc44GNS7nZ
cICf04uksfkQqu+p31qSxzZ5gz+XpFQduViCAFJt1M0LsBwMOnSfexLyXhqQzB/CAlmLCGLSvh8d
DVDXSKQYEIkvNpmknHGVrwSWXQkoqTf96g/9ZFO/3Kcl6FLhYyLRa421Oqek7rrMkP45L3trVqnG
QseL4oPRJZlBYeXw58hS/esWD3JvWj1b+4oDeuSC1HFSWXAfqlMxXasALIY2OX5B44dMQbGIt19H
gUvHSNwjsS+iU+qEixMaLMBl1zxafewM2s3EIvgXg4dmA1tqxwR/QJf2Oa4qIWIKG2JJIaHataoB
ZozyvQsnnqaJQ4jvOnAudCn+jGoxELWoYFAPrFn4NRplZ7E+uZtINJj4d8TRMchre4j9rKfqtHIz
onlVB25Vg1ZGcWUWsvH9Zzby1O+3juPg8b8skr5db/jd3B3RDYAVGzBMcvQE6zQLJDCHHZzbc9m3
1xyg9U0TX607tiryIqeL5UNa/bh2wi2laTNF/Us7UNPgrkDBEwSDUKDr7tBlR8CGuKkD/U023n6L
jfsfkck+Z2XriJT7r6DTA25UJWKCMtun0AvlTeF3GDp8emz/TmmvbPcY5GZjPFF+rN0EK0qNIFfm
rma4KRdst7ffVF7rFVIvQc/JqaQ7eH/G4Ja+8cVTsA2ROl109bX+n+yXACRO10nKgf86OpydxYv0
tFH5R1BWz4g/qR0xQTlHh4FE8swLyKsydKpJvpUgXuQWmcOZi/KUXCE9J3n191ATBarFgFyZcSsX
/SvdGUuyMY1FYoEH7YaFHMmqRi5tyh4xNiJDZhX6IOmDaUvIpUk3ZjjI0ymXdqkJ0R00oU0KZ5OW
tySyrL4MptI8lU2/DrB9brdjtgJAth3OIJ3gQXQsmr4Ej4xIFPFYsHdYWiEqmjwUSq8NFN+fRlO7
PISAkx6I5LP9uPEGdmBzn/882aMykeklkfgN8lFqYChSWCsoMHyLx5x3IPA12hk18ZQUi9Ytaada
7elkElIsmJC+2s7N3c5o93SMrNXxN4ocupFyBdjtrNnNLGGURo9DGhIkP/z2LAvmDIGS5xsKQLEN
4h5UmSQ16rBlWJ8PWkKz15fPGHTlxquobAdk7es57+R7Pi0lZ0+FuK6Sa0TOx0E8U80IwhqPav11
XURUIL2d8fRGGnt31fMKSqu3SMmAu8erkdhFfTDJGSzU8W/mY2jvVTWk+KfjUSFvx9sFNjiJp8/J
zIbB8A6M3kQhDmM2AjG+M2lLGqpfuswxEEq0cvJzytel7jCgt8sg3DEGF/GOf7IFws97TgCOjlJK
C39JeEuLD8MWnDZHIfs+mCPw5x5XfccEgyoRxSLUrMiHnv19xuDqT3Y+e7A5r70ONXDRpvc5IuEW
W1CGJSNYKvSgxUiV+MTYxHnYHXcFH/la3pvRu3YLZADYmcFJKB6AV/tORoQiV/eJ9tfeA4QX2LfF
W3k8dOAUk/Woi+swTKLDp0zd8c0xMdtGsrY/VawOt8UfUdthv5OjGpLM5Xw0nPWXlvG6HXOo536H
iak2tXfbHJTcbq3VjZTt1Xlh2IqhsYO9J46OH6QthdZZ9MTPrL4Wr5m799lq3zo0OfoN9hAhjEzc
S0RV1/EC654BN1bmW79vLNpb7bzLPvaoaoqg/zzNGDdRSZLLj3qmIYx1Fo+Pk+K8CxdsluZ+T5+u
Oz6FWvLssvRDpYfWWgIKOxxqM1pl2s/CfqeZzF9N6ZiV1U5ztpJmu7NkgZjy6wSBHoFJBQbPyiwA
st+JcAnLYxPOYcDgZFvt4G2IkPfR4NapIGBtfA6rXXOaziih1O8N53QpxPuZzFjl8+aUH5sYM2Wr
STScDmRi3jWtneqYmFceDLPMPZC6Hni5i7s2lWaICeF6tjGNyt9MCXREbOORM7xrNpIWgeIvnblr
O6p1s5/vPouvFN8OhSni9GS12BIeFtkTkDpPfMK7Xc1bnqSBVsp3iX1kdDS3y0CE2U6VgSPFV0Sr
E2dNY8uZM47CV2cPx15lML4xtEzE06WcJjNSU5/6YAROKXVIL9xf7fTJ3NX+KJQbCSLcOJXRa6fn
zXEdVX1EyFjTIk0RcEZFfQ6cSTYVDWaeGnsL0Ztd8lS/y73oOGGTyeGdPC6S726YEU6lM9u7LuUa
bCvyWdS6evamdAhCkWHV72pmBbdvwNmbSCKj21jh1B5sTp31GMP8/XQbPnRBVF/cYG786v+2cWyA
LC/8vh2KanDbmETn7EUux+Ot7wBkI9MQATLIOvmiVQ1zLqBHbnv5RSzV5pfi2PXCW0wKkpldtaIE
OC2Vjx7nww1JiqwlM9rw90/vSYeMFmHkwOiBg3WxnzUqPv9GAgRSAm+z6HyxoGHXMcwQ+ScRVHLG
sUlk5x0Xxzuh3wJ5rxBMIB8/XBUS+KiziiSFJwDX3sYOb2//FRVBBpovm3NJ7WUZD5WI8ev2+8Xj
6JyQ2Gp1IlPh2XEE1uybzAw1gwQd0NDpMQHek1UOdW8eJn9TbHQeFyFrBbwwcY8BjcV79Ix1erpi
59VxfeecPM08FmyhvrWzKSvA//BBixQ2F3GiqdW31StXXjG0zH2tmLza7WQF5TsYz2Vo93kl0EBL
ASSrSfwAOHkbvl86qWg+mSbraQ1CZdEPRcldrgS4ocM6uP3A0HpIXpdX9s9k2wA+0gpgiBjm5f0V
7k5tl9BuTevE6LDz3yyfzOCwVqGNIwecnh+w+UVUCZ82T5xGLzaIq4LMygxO0DZy1/dxQFVb8r3N
l7/SfEbgvpL9RB3n/v8TAphM6roszE1QEljqHFPzo0P3KUv+yFtiOPIf5cH0r6e1y1FqOJgkTll2
vjzqIg2fUTBY4pl5qwIyA19c1UxUzucLUMZD4jxPSCaiAvxryzusvd/SDBj9PcI8pGmi8/RtgDUW
2JrUjPL+r0KhSoXulie8IHknFfRxlBciD7eCmXyRjmN85rZqzz25s+qBvfwgqAzUm5tNsLbUhB7w
uwhOv32WyzfIKQD5xxgWjtRpOzYkaGC4Qw3TyN2w/84R7BaAng07ma6emNUg5uaoUkOJ0ShpWSWc
+si5NQCmdp+q5IhL1RY2zUKttG7X5RezXDV6gG+g27CYMvlViKoXRU2zsP8AIp/CbfjiM5nwP8vE
7sTcZX3fxrnsaQ6pd8yMx2WRc0ldHwWPBotRSIKAmLM0wX6TfCmQPxwOxdJ3kL1ca8WzDsEoR7KT
s7UGR9HvKlvTrGlHPvj1CWj/p1oI9PKcOjzS3yGu5nQH0Elu3Ubi69ilpsIBYjZmSaE4zINtmd9L
aUXraclYfeJW4IIfjutrBp/I/5UgOXmOmzvDjwWpsu2DYdpWtMPOT6Tp7K4bLrO6e75DOeD2xMrv
YXo+9cfzkNSZXB/3SV2rus8FzCder70PMTZxHDRL4o44iAjrAHgnNa+ZRkl0NH6zNvSUKZYiByDc
ONZPPzQxZtdctTs9w+zJ1jby/dH008MUcbMg67O3eVJUEi2j8VdXolFWTZS5rCkX8nTsxgLIpePx
m3s8rIYGPZUuESyRxnYgeIFwG/dMnTIGpSv7fqyPiijWaw2r2AFvGuRzPGjdvD5J+iKteno03W33
5PNApaaHmpspGhfex7An4zKLLcbFtQkQnq6lLuL+Gm5+5D4Wi3hn3W8UGYrfnyijnjSsSEGj3/CZ
9E7HqwNplYa3TnMzNNdUN2Ho10V91Klw3F20iawsaU2APM1UJOlv9vircfxKcUKguOLw48CKtycY
R59kdsKCMfQ24IDc8yHfgN5dp6rLdodI0jdI2Rq9kUdg2angEXRMj1Kioom1bWNB07FJ0v7itvbD
rkUT3gnft1GO6TctLpxJ+jFTXeBotFO+Nus2nnyYg0Fiqr6nSGdAzMeiEbP0n80ZVVXicuBSi79v
teXivYBUq/kUAf3AOn/8UYLc30uoTnZbCX4v2i+ZOT49lGZXKblIiuDjWdXac6tI8COCU6gIeYvB
6fHLfhJqVxp2w9B9BEvWcNTPi3tSyd2YlaMQqszVI62rBFyy3fplHzYeKtmULTQiCv3wQS+YIhep
fRsOhVVtp9D1rfPC/Aj1iMcNBDW347e1I+rZFs2dDNjaMTPg3zh7dFVkoL4F5k0DvWX5sLmkXKzI
P4PiN2HfuDuqVqQcNr462/QzAAsA3qD80ouh4C21BDyRi09wtYFB1gXEfNjZED/cc8jrJxc9Nder
t6qIZ5Acy1mzK1xDfNyArPktSoNxKQKB9JlYWoDYa9w4riQXCd1/RyEXrn7H7P/F+bVmi4V8yK00
mSxIlGTik3LUeyzE+dPg7jv08V0l0jlJ0nJNUjBRZMTnhK4UkKo8vD+9o4gag7IhFa5unn/QqluD
u9gyvwkKQboxqEYfcjnwga5neEm8vqNxaIrVeIKPgNvG/5F7qS95UldVw7DA8bWWeychG0Uh+D8W
QeA2UW5mMDYpZzkWgU350meWMT7xunNmB2JdnoWexX473O3HQ6r1v5J5DHBpR3cOW1C1It5h4z+O
s25Gw0sHduyjnRBQgA82ca3spqUqz3KGwTI2Mvc1BxWI4797Y87sqBrcseKpeNq3xC2bkOOckVwk
0awpzBbOeJYzcShCwO5MwEhxtVT3rhuYDNXxpGxH/ydiITx5CKtf39wTbZB72kNaE6ccZQs+YUgR
3YoyOTu8pNGaeyr+LeHSdamZ1Rv7cbPfdBZHaaeZpWofl0cCI84Qe264U7O6rg/8ZXdVCtgJdfwB
jluII73XwCWRZo+ygPG7yftENPwUKMT9YiNMMPjoVxs0MrsISIdeEALPiY7rfbF9vfnZosBlmSJL
IvdxvMGoWVTlMYK9jL2Xx/ti1hf+2HUfEvepxa0iMDx4dv6LsuVAsyeG+FLpmUf1fRZVEAICDWcr
w6uOzhZx7a6wd/69DgNs1t1IIH1Acf4hSJHWT2fNQ4zmMpDzuvTW+nrKY4VKfN8J9lI9rN6gh/BB
EIAx+cVm8mjkDxl9LPMX8ICbgTf45Y6h3yULQ67rtAhB87A34n6iVcrcDTG9pkDQRuaH+TxE6Gl7
suWxp4QOmqREK6buLRmrV5uLQyCDKKR9Poo2/VshT5ZH8d28oBuJspwaLVFIL9qnUp9Tv3iaX+pL
k9wm61bTQxkjY5Npuo8o0Lygltq/n1flU+wmVtvStk9j8tPNyA4lXRdh3jiMJ01XVWS35nUnkl2A
G6MYSvu04KsmRoamX62PIbMs8wbIAt/e6H47EIcdE885unK/edivi5gPIhtDGBkbXBQYT+0bXC06
n5eCr/xI1n9z4QUnZ4uWZGqPZ/U06nnFZjE7MHyIpAXUTseTmAVY6NK5VsRa71x4rDuE3OQcG9YW
/sEoWli6SZrRu4fIGIaM4CB5P/libR7lTDo7o2FzMIGnXIW2JV7A4+3dUUi+J71iEczqGQIb1c9U
0/+t71xsS/PzslG/wkjjMDVJYcO+VWeGKixa3WSdVyYo4eEMHGVFeKiWgch3PfHLR3laikLwkYS+
b7cba6ekcYiH7vX7CCqk28lLlN1d+Qz8k8OtOH4IOyYnL5IBlr9yRuowKoyV0VqOIL4Cx42tKrXe
nRcXdmxAvjk+SAkeeGcPFwD+gHlYvF4NwPUFGbmkXzFQWb5HPqUfUcGZh8pjS+Qd73MhIVuzgoy/
S2SP4dWdzgLKsQKdXCVBbmDLk4w9c3HewD8rPGG77BF5+e4yWCA8AnCr2aX9yAz5PYsSvhO2HJcU
LLLtxOHpDn8E6IZWHpkdfhLJWT0ls3X7foSyZa+gydyrS+8BwIKtUals//EGjPW6PBgkCkQ2R9T4
1ukLJXRDLHZgkDUkDLFff/iFUx3lTzJ7w62cCXzTkLTn8CF+Z1Yl4fqKyPwkeoo6mFLlyF8aLQq5
7VXF6EhqtTw1DmZ2lX90yfMC8DLBX89N/+Rqa4WFHt5yGbDuDYM/p+98O8oudoRLVGJR+oBfVEBj
61HVKi8WePYY2tjf9lgZ9svtr+gmJHmH75mZMcJCR3EmR9oZKr/MKggSPmLpKiZFJU5vVrJEb1fg
ziLSdyK4TLkSSjsPuhg5u61xzXWmme65gtTAuoFi9129guODPw0HEweRRZP2D5CtUIN9VxVL9Zbp
zAa2v7iKg0FEClub0pxci/QbCCKb3dfvDyz4oFeB6eI2Ve9wdP9VoGEvpJ/z/1flwe0n7j6Aw14w
Dcsiw/z6dabDJDBio1ZwPPuHOY77fPwt+aQYNpOR4J2UE1gE2Ct7DIAhRheIwYZYQByUFUCB3DzS
XxkORfdJOym68PFPbqBbHGzz/j80VjrDAZDwM5rGW35Rgcc4eZWfYtIO9T3pNtGbewRvtlLyfLYI
C8Jrkgn/oR0eT4/fwWN0d7aHdHiF2ecC41f1xl/+JyoiJlpsWMga4NNMbuME7/k+DqPiO4f8Eg4l
ZUDYPLM50nWxFrLHWV4pTuzTzTKV23LlBi0LS/E2WmGu9garGsaIpEurFr3rEpk1sTWr3RsQA6vE
FwxqG+hlpt3fy/1zePkM+Y3K1dNW/sMuIxamT9uE17c8gjvU+KjeIUFCFxGb8Q09YaTTCDcuoJsA
cwCe75FTuifu0hS49wo7wG3ZYhVgadkIiRRn2t73s1qp7MCOToLJA1TC8rqbTwBPQ397QeeKW9xd
OVO2ephl9PzqIsvtMN6iC0Zj2ZCTLC67WtCnBBSRwZt3xZyo/r3npvJrPHRR7JViE+Th6+Q2LAGd
3Tx3Z8u4ABiuV7Ka3A07x1fmOcEf6iuMHHu/o4OW1G01zH5u1B9CB4vVxfNLRkql7iZaUqNQtlFw
vX6z33+mAIbFnnFtKwzFQquedCvcDLbGq8PCMfH1eIek3Wdmb3E8KPkl/atCegKN+F4rNoIVB7Sv
EdCBtNFdQKqt/jkJVU+T1c6EZgjWnK4eP7SbRC79ssNwGIwKiakuCwNeMuF36oaS/znnLBA86MFY
Y3cpl9ReK9y7YEy6SMVG8gEQ0VmyUNnaftNK+xjzZ1mD0Glc1UqgtE9TUQkYi6jfpl5X4Rr1WNCx
/dJroudRtNqPe95c+EY6/1hYGQsyBe54upS15kIN566eB4t7yQj0iuOPXFYtl1xghnt5mW0VdGxn
XheRNjTxvKEhb/ppL6WlvtSQOsoLIqVLx2G6OZkdH5SNjbiqczS52NSzX3Ru7JAuTfLyij0jj8I4
mgwUtHUc1WC6nNWqRugCtyQSUttP34Pgxd3ral0njX7Ucm/NEf7dh3b/lKeqNyxv+A6agTlzGMxg
xmoHyW4RoWDAzBDDkhuCLcYDPnyQlKwWwNrGXMUxvdETaPJk6Yu9qa3nbQeq3aikDSAjQD+djmGv
qD6wVLvtcTtxr/KR5F9PPz/COCFx3XAq5EBd/GQO7nvFu7G5FJ0+wW7EJQdlSTJO2bBzHcU98O5r
CEHEPyAcEyAfrJT0fzejCmBbKhoEhC13h+gC/2I4OYskA1c8/6dtHOGNRlsPydLwe02xvNadhhoU
DnaE0eyM+qDDblXI2E8znOrjwQFCT8V3fHXv7RyLzLClYsAskyuzfMF7rU9kn3H5Je/jNCx1xyMM
QHk2bw7Bl+TefAjn+wiZgtOhMjjQfd6p5Eh+Qf9D04pMuK30dWgS8k0ueTZ/Pg4I48dCnWXB3qvj
wGx4S6STx7CgN9sdzwVDT1r2/qu6sRt2Lpv9kTb7j0aiWRz6TZd0i5jN+ZCVvU2dNVXmtC5pOX0i
IKxMSRAYm78askgmTIrunTEZ7nrYv3PM7dJ1PPLSHHkWNb+vjz5/YYUkWfOCfV6nWj6NSGJ9fFBz
YbenXHAZ5VmfIX4iiJaqn3h2l7IVgjpGPjWUzpTntH1hRJYg6y63up3xU+zE8CsEMyYZZZfXgQ8v
OLulFav3sIuHf+E1jb7740v6on06qNFBRy9CdeFk/fTDcKYMGw175mPE49aQNL0SGPRNPvtukxeo
OaOkef0kkri3wP4kqp8xZaN+lshO1zsDlzpuaaoyYTLKg+2X3nRxk5XAvHTCug97M8mAMwlJFD2l
iB8ZUbMK7QE0b6UlrCfde+FYRNR/4NEH3IynyfkKj6zGmN598A2v7/ujDImGzkXFg8Xxvpxno+f4
5DSBAKOE8PnhImK/wIC56olQcWwi3Ol0MpHaVu1590RxCGUEMWqt5MmXOsEnFRo9nnWcwoU4Xqas
FEQWbQoOXaw/gV237QsHc4XTYiSUHD/DslsAB2QpQiBpaLIRIcT0O+YddMZHFPFx5dDrqUvj6sYL
lrqXh9rzTEm+G/HSstMgnhpPNtl5Uf9tygDip8SZfdp0HZjIIje55Sn8QNhwq0QwQfxVuarUUmuU
2ev6dnvZF1DBhAMQWHty92L0DTjBfeHf/bz4tVlx3IPMsYfT/A3WkzYy2KHdiJ67OOTUHPTCBlTm
t0ae7F3e01Mkl7nYGxxEM7pfwVlZPWJtFpPVTu2BHqa4jkZhvNF2kT44pDn9MSSYFcNzwm3wDMoS
R+esSsiTqlZhDj0yaJHZxa3U8s+91hdbFgXJbhnb00DF1jQYEHCG4BggxKjscpEbdAm7eYlgZ52y
tn2rqO8VIc2M3b3WEA8tCAW5EtL804YTUIlGRmRt2RpdA99SpCHkvsjo65pRkkXeCDP10/31A/tS
PClu5ruR6Xwj/IDrXo4gg34HGGfQZZfTn2OaWK/aw+sKIPDzswd4Es8ea5texuT5IFPbzAkGkz1H
X1jOU5dUCnmc5lVo9kG7a1RYIVH3I8oCYNxpPDiIO7VOEUKMZD9ImJ3bIqcapH+zAN+/kFMBupGv
peQKJxcP0V2wdUUJei15271P6F0cH/WBWuo1D2J9yPv8yCgTeSV+6lemUX8LwsqCrNrajhPYvW3l
rfsgSHJA56Jmr4hPW5JKYEak0aMj2FefH2KslAK+AzqdOBijx0/dJEV/7X0y1V1cq+ZlnggaGUnK
zGrLOx7TB9Taw2kQ52DlEynBOaHnGwp5sTcf8M4IYOVreWbbZtkw92XcZp/VEMS90spG/n3UquN4
jRH8v2NT+UYRD/RzldJHumlBwRbJDmhkKNnRrG7AFJex5B/hMPXyr6ybEOygzHsnBYD3J4G4fi+K
ukWXlgMoz8RSwHBbbSHIVUwL5x4JMWcGIkBAWW3pHhzWAznk6mOun9Sulvv7r3FUI3Six9gvsTbX
y/9lQ2A4xLJ+HjUCPRbsIridfFbY13CZTXV4QaT6ogyk48z1CSlvN+H8UmORMNNKlZFKaBGPYoap
5b+bPYvCjkqW9N2bOsQ+zHmEUWGxMBIFkUmIf0YhN2LNOckfh0edY9ccA9RM5VbBT+pWXGwhMCU+
0ZsSX/eTQIknUsF8LSzQHcKzTxIREdtsjVBrzlEZWiGvwXqYuF59cbJ7OXGCgtZOa+3H9+enm1r0
wlBlCUfTFI/QgffgGMn49Ee1tRqht7ITOzdynOFfMy5iPTpMT7rX4MLYcR8A3d0HeP0uG4CgZIv8
5vmc43ZzXkmiR88GHV30JF+m81Hl12TLKRpmN3nC+7sRpUF+Kp5UZDTrilcKDD9JlqBFpfSJhl5L
V9Mb2HQdcYEgm1UO9v7S/gY4pol/o3tKPGtGCoqpo9y+3ff++IPo8WMfzYs3xbQ9kT7FPmLLtPCM
d5AoeOHGZ1/FCE4cop6e4ZBXXoYIjfbcK3Ehrwace7K8DgsC5YGTJ59CziMDJhcIkPqFwdwsDNEH
9wicHWcOeaAMibk2xsEo8nLOCjnk7n81sveSJSMJqElPYadzzwKRv01+lItsDxDkutGCZAoKIhiL
Zky48UMWKf7rRHn5zQv2Swfl5I9o7Bs6uM6POG8LSeQv+87pqHGtXglUpdszBVRkh1wJpaCB5bzY
cz2drxijjYMXanNd6NaINnfIp3QLQADtlGgB4ZED6l1mZqMWqhPXvN96SGaGrdY+eT/jwMPkXSKl
gbyAoJzsM2IrwIFthrThfrftF1r537wY5Tb4xSN1UkagDhUgc0E4N/XGNoShsJYLYMSlUWXfo8Ez
nfJhHasvSXTTt4x+WChfhAQPVUt0ZM6qMn9md+tMHnFJ4YWikgfxo3N53xQ+xwKZnMsWr3Ot0ZG2
Np7JvQq5SM/L62FaGe43RTZCPdUuBdMfhp869Tx/x9w5rthlewXK7EQ81BdlrADRAR3HiCymJCru
TyRdPsCnTUElkpmLBAFIG4V8iu22pxoOLaef2Cit4lzSlYlXIw19I/n8KA5l7nIj2hFFULyfslRV
jRkuVNa11IDfQl5nQSe8OsFsh9hUbXf18Z1SLXt7FkKQ9tzPxtf2Wn/3Kcmc6lQ9GRVmN3GMgGHd
KWpjPTxD36FrPS4GEdauZeRXogQLgxogmnFgCG7xz6zxjDsMfEXDaenNi+Qwldd0UVp5NL5qkEF9
KIwyBQeW6ZNgKs7W1OH0T+uXz0n8/+WkbE2OZ9XgbdkHHK0x/OvINLOJ4pigyPJCq2Iwpp+Ogjqg
/CFNl3DIgHshM2h5YxyO+n8o+uDrMcriz6uV7tdNJ+JGVLAnIWvrhneiXiq1/MSOqS4uz9ojthcN
NAYUSXvBAgnVRziEUGeXdwa9mvLWNk9spDXubu88ZPApURemeUtNvxq1ibH4bE80pXDEDv+orJDb
ZK37fXLc8LxitfAmIWOMzUMKTLJIAPJzaMVfyM74jPRTP3wI2cUUPnrgWWguXpen2sy94kinTpz4
hUAV5MXXgA9xf5gFFvx7Ut0lF7Ome6stapS5V9UqF4/515al6jGMBDfGZ+UQTvakYpvT9GKTE/EY
UIEW2sOinIYxYCOk0gaepdVpBQ/oIGu1SSM5CXpcfW9JDJGr297kV1YvlIKrdiO5ENJUDbA+yoEe
/GU43ZAE5va4CGZEufnLO9u1zQuU14mE31C+tDjZ+oYLEg/tO4ZKwivSXR6GUZGTKtanl14KaDJb
5I0uUD3yGizgHu7w80yPYqqjYNiNah3fpNxCp8BdVNT6fqYLGpxNgXVjqps0T2EI07SuZnvV41Ja
KXd3AcRO3Hb1MMFxsI5y1Vg1WsyM4grAZN3GdGywIaMpB7+wwoRgjSbZsA/RdmSE4iREIEc039Ad
IZWGES4DGexqNPG3O1dzhL39O/k7SUB3iwidSMWPGMdclP/p0AZPSakC/Lkj06NAabnCSZjzoyjw
1moEaXEy9qZIosLW4HlpN8vcg/CDa0gdjiVD3SYYgjWKnAQ0M5/5jcqYnKVTTIxg4odToKn+i/iR
2QXUhxpLSRxbecHp9Zdft5YGwB1wJGNbGf6ZMaU+Su4AmKFRJRRn0guMXIFx7FxC1x4b2uYes/TV
LjeM+OzFNdH4/Jzjm2dmqnWw2d6lIb+ufzGTjWr5kG7JbS0F0O0emqbjg1FyaALkiaYtsVFsnxJn
XG4JwIUFhp9uOil1Y2E3LMuGifUaYReRPbGirQ6j4QXVG1QcpBesBMeg/eptrlSP0UPR0NJmf7MI
MXKigNBKB+0+Xrsqj7DY/Da2vbBAOrunfP1ef8C+84j24l5TkLU3rDcYhoUPHc5w72OB8nf6+Aib
ESk+gO2+usz2UM3Dl1eIyWwwZ6hlWKAVYCZAYoHPhgoDIpv+rlLLROjh9KV1fvYikff9kwTG8RaU
fo9oun0JTd709yRqdD6V2+CZuT3scT2rvSERqrevDoWBViV2YuPYLTLdXb8bZaQYQLYoYiK/n/q1
ZIZ9Lb9lj4mV5Wq6YJVKVt1xbmswDpAfa84jXZYOGRroiFtuvJi5RbZpFwRNxdU76mkm+WCosBdF
iivAIslL7NhjTF/EQHd2kqPIDRIiGUaKyAojEl3GLnfEUUiBOSDDWnw46JBNDsEP3+utWraxMHcD
WTOF6ki0dIur9xq2hMF0/8h7Q0kZpAYOkox4CKL+uFBxjOik0lxJGgWKuN2cIOaOG+9JJe3Uvd8W
WVeXiTjM5efaA9VHYcb6yKvo0lipypFl6UewF9P783gwrc9fXVY7YjjlA4ArOz6FM/u5c6VqENMB
VnOsoC2ZcRx2aSkchbJi5+QNDCHWjzbHpDcukzkmbcwZOIaPjR9FiGL46F1kFXmjfd2dPnBPBkIO
DfyhbRjXBA9EwBVSddqAkpAdSxh6pVOteLmqcUBRleCR2toJFcIGct8+lWp1Z76AKdKCbTSuNgrR
bq2qdT6+QWCJjyahvXMmkWpyJh/ioCumr1kNl5ZMar47IF3vcqM/VW/BF7gtQVlWeVcSVjZE7Pwb
gBY8xpm6WKctXo1DHcjIRXe4Jo02EX7JnFRSjvX3jONd3RiESfP78+qRqMDMbUBAY/wMjFxvBRiX
UIGkp5jdmAgU9hzDo6p4eQ8cQxMUeeuV1G0XSJRe6xMhIUwIkVnGac2JNUMAcyr4240ZosD1DJMd
r7dr4oKWNEKZz/Gh+OlBEFo3cTc9ZqHLVbUEJVrCVE1YoCo25s4DNdDbMPZ36dR/4tfvIEQTkxAw
IPsgTVVPWh56J1qw9bdul28OADS2AtqiPPYc3gbmtlyh8U/8nXp0w60nCwt9pgDpe5YhNCPWm8v5
ond1FA4+oJOyhHab1Qd7uH6zbhAAx/QVASJpM8IeKI1PZu+RJwV3zSmLg2mQdkZopy/mR4wl/muE
4LYY2CURuIXDAnmVEB0QSLNSYnOdCHnmdwgNcwpaqpkFMrGE5iGdPakF1MGnzWXtZ+LWf0AF2YBK
vjdX8oAf2KMePdVxShcUs2+FmPRai6q3yjxRFiYp/6IoX1aJOQok5k4N6zYsFaa9M0urq7J6y0qp
OAunrYJAyi5pQ8sMnN/7SKrTUhON1tb3PPZis6cXZ0C4U02ezOP3iTrLJJ3/wFDVZXrp/3lfw0bC
xix4RZjIt0v2hrR+lAJ/hMmvOZMO4RFp+/gf9oj6/Ox7FE9TDFxTF4ZFts0ftV7xzyy56ueK3IU7
8yj27WejBkn/PCECSa7bQfTZaIS4tCdrIRpWnq37ux6qOHOsot8L86FDTrm5k9/zX+qevSqZKSHn
sUR9QUxBaKLmxF2C9/RNSXDYuA0bY7TZRGyNNcucDGXCSJvWj2Y+Adc7G9I0lO5P5NogBgy/+OQp
Ilfz4rVx2fWgwDrTbjzJuyJAeFAVcJHBl0O5wXoa+lKhTnxbYXKBA1br0zlXT3djka28O0zrPbt+
QaXjkWP0VlfA8uADALF+b8g6UGbjyLGtM9Oy2PUA9V01S1Eoa6tXAT5mB3Qm1vv8KTlbqPLc9Fnn
lsQMr8pWPHjETSSGykXrfTwbDybggTptpO6FI3ZMZActoCtuTYJKWrhkblB2YTgSgKGJxW5Ggm0B
/HJWDp5hroCDJddhGK/knxUochOw7KVXimt4Yg1zxhSFsWxbhqTVCeoiEzFZIh1nFJBmHrVR5k8F
fWv3CXoM+aB8vPQeRQ1jTQjDI4tLZ0BI8krAQVDllrEINczA4QbFssMGRFoAHJ/fvY4QNZSVivM0
TsV7nehTIxRyYk6OUyo6vew3lvFcLOExF8VDbP/7ZGHd3KSVhK8pHln/WlcmFKRZ/3/SOgn6pUuu
ovr3lKVcXu4Aw62DbFiw+HnbW8FcYZV3u36zfHp/aNW8ILpf6DxnkQrm37RATEJdlRlvMxf7x243
0uslO7NWV5WysatGpXWx4XmmMR3oH6WD+j8ZT0zdIXzBGTNVz79mouOFlhP1dplYYwk/INFenMDy
PcXZQL3YUYkikCB2jTEGhVzDPh71h66ud3X8M5h43Imy+pU2fBDa2obUYEiX+6luI/bV4EZkJ93S
BVLVplTNEODWz7idREDbFP24qjAMUt6benv/nTcKehfKbF4s6nsi5SHflRnGOux3maDbDSrenzvj
97sCgnNzN66+YRditN/zk/HUN0ezEMcnQiPjB5ryyX697MWFGHQqRBwMp46nkrkCSW5ftf5KDaR/
OENh4xGTLWQP40mlHH7puACNeah2vHkErvaiXgXDWV+iHThwvRWUs8VzoUERb5nIivlaIZ9jQlwH
fN0+/zrAh/5UC+iig9OeLqL45KfO5MTP/p8PgbSENJsNeJwx/R7+fGu2hOUH3pno5bNSRLUYs8/6
pvCcVBMvpuM53oaygdD/nriEEn3XWqQV8kPBY7Wa2UKzPO5ezS+x0YzdWQiDZFuRa1gqmxDG1bhu
TAiiO1zhj1WEtIgnz49+/l/ujsHyqtJBQXk5MaSiqUjZTABjmw357Rzv8OKhe4rDXHKowzw9T+59
KOPpMgMRcnlLI8QxdXChrNvaCZuT5KYIYtt4YsximpXqQzXyI9h2yvf+VKxYRFVY0cylY+Eqm9zK
OlUu2Fy5+4YKUonK3p8qd71ZEj42AlizJ0q9C8Q93vFMur4fTiuqp0pRiJg4H9BdkDABrJ3HkK9d
y/v9ix0WG8TXQHRLLqDYBc4KWEML5rHWAkZOPumKbkZc/Rulioiu/xfIQ7EP3swtImX7v9rKEoZ5
WLFGP6Xu/1dYZVv5NkvEzl4xnpdzoGGf9NxF2+yQf6noUrt77QcLg6qAwWp2e7f8soGHgTi7leD7
1oz9a7dXOd/nmPJd5floKdz9/ATJmbsDIhhGnSLKuAtQq4+7mAPl4TurKKqn9ZryA2QIS91ii3Mn
s8TcWB+VhORxnGVNCH54ZYlmIHeto7XuTsjV+gMx48hP44d860UMutx2cfXweFqe1oNEhskeAbaz
wcGWWvrqG8l26CMbNgyCn5fS3WnLY8aybj6Nz4JIjIhJ5Ca8MNDOvwtNBEZ92E44b7oY5cNj0Qk4
tVQfvNCvXarm6qeMtlk4q3A3SxrTNGgm4RgdFSD2yk/ou3FXRODW2yHVfp2tTQEsF4bnFZzZLnzf
tv0cQafgXdv16zAAJouI6htWlH0ILEOa0FyyZFNL9R/+tR/nNpvAQRMHJQC45Pq31OhP2dmvSBYb
XTMXNQXKBHwKxtvGsHQ9lPThM48rIGv74GDzvANIREzE83q531F5Bqg0jwOJDWL0MfldSKdOu1A5
3rCH4g81PDKsi+jFtCh7LZXv/8sUaluT2vJcUIyo6qFOlNagXJZ9NQOosIV24XlhWdUzqNxLaYiM
lpQ3GLosnW2DO2uIa90lgaawvAw4/qrQIZ79ZCJerPHUjALvbbK4QZdg08RrOjdXihdWzUNJ60XC
NA54J7XVkOXc3NOkdsbCWJZ9kNITU3q0Oyi5gMmWdoRSEdiqS8Qm2fs1R5jvA0HEKjoZ/bo94wUA
a3qBC6sGYZxjTOCAPVKZHKByGVSW4DzwFS4+uVa6T3tQcFJj7d2zaBpus6H1NCBN2VlI367DtDGc
RfCbpxS8ehUzsz0+zk2XbY+LhUg9EtxFAOl3NHwu4rQ4tx4eQowzXbg0Chs0fpKfKb3RHDvlpY6C
V1uEmhbxMCSvqnG/EeoOQL7uSAAbaN/z/enrNWidOn9ser3EhDLgL08rXbuVIv5CSCr9CEmRMpvo
3ojqRP6Tp87XqzrsKlPPVdE0m1K3gEbP4/tH5fdYVU3p0JFkDb4uS20FzpqeXyNLQP4K9qcrVuFD
Hc/UNdkGP3wt9wpzIm/YhQ1c1R0Ab2NfrQAF7EFgmt/7OrSms8+5CZ0ON2buHHVHWuIsrpAKFWm5
Pd+tIKyEKIhJXAMqEck1/JKXvGBQ2vjfuffcfxki6ycpPLBBzsAap+RcpNKqNSvmodXFEyzHfkIO
aM6Fnlweq5zuLy4bg8kA7l/oM6cUM2RmSQOwx15EAu8sNU6shdgjf1Mmn4exutPdptvNRjvM5MAw
VlquBVma0r3nocnWqp3JjBTPrq60N+x4PJOHc+n75gPhfa3wyq64hlVQjsJRwQPilV5kaw4Jg9bg
lOXg3YWCZDCjIoWywoIs5oM2bNSpVIXFzBgcN1jRePncTMYQ0UhxD51dQYXSUvsvpoqc6GwfjfHP
sA0GmZCWGAtUIM5Tf3DM5AiMcExOevmj6d1eDhs3GvVW6hFl9DZ72JBYi3PEnMz/UFjtRUtAvs+c
9+Z7CaNF56xnMCKdM5r2GbdHJ4qhiqtgQe/sgN6SAuKnCfd4TFlTn+/cf9k+70aNRoLlJc+GrRq/
hlAcNrM/Bk6tpM14l/AZMfbA3fQVCu7XzHwudVOKyhq0PgkC1QJUMJtkd77v9+VnD35965inV2tq
ICTdEFtzozsq5sWNnRNaYGunEHg5TCpySEhnwN9GWwZgxrwBUBUiI+JwjuWYQI6GUDMc4XuHTx5e
HVSvaj1miA0vvsbXm9oBlUXRD1ECJ23Z8hxHzQm9tmxToGOH9Tzb+9DYe/p8Fn80ZcQa45RapUmb
hNI2rinjqKVYpKsbTt8KNbV+HH7O9NHRGbQVhR25u9U2u7BwmKxol3exUSHLw2QZeys2jCtDZApy
/XNSZJzpXpMFos52NEV93rop1/Nicet3XikhdpjoKgayrNgXnRzPYxiOMC+jfWk8DfRNctYXqwlB
UAv9NjDWqoRRckkW1xo3K31dejpefBkYYfVM5ErYbR7jaRbby8pKL51gLwDws/VGF+5t72gASb5u
WoyJgsSXCQiL7mVGPi4+2Sk4NA+03noclEY/5uE3E+HasWpZTD94x1Dt9WFM4StY3CFKCEeGTtJC
7vZT/cAyxtsBKScXBW1NgDTQdE8IigZyRwDFnHjDq4MDP2Nlm3ZLLUQNonafoVgHQmKlEeh1mN2a
YLu1gXP5TW5HlEOzsFr3XJQ0QOvw/rsrJxlmMmInzG2qXHfhq/CzhJm2snuJU0wMzzjf3Q3TLdQ4
rH7z3FYJ+U1FK/tBho0yRK4pUIlaFcJd/9Me8dYbGdx2pBtDP8tiRlsVerP5uYfv0//XbgS2Dn5x
x/LVOxmrgCR9/fGVM5hoSEc+6nKDH3xdJ7Dt3Z9599pyGMQm4o4E8ak1AzVvicxV/dHA5DERXgn+
aUBHh6R5pv37GLIZGKK9g7Og6IVDX8WUzn8BcayUxSiUcGkePHP52cRgWXChH47pGpKWj4WXmrym
U9zM53EFoayr/mYzclizB1nb6Ei59HaT/NQCieJgCgZYCMFIeRgy+OUwBIi1FUSSAp9z5gPbIdZg
E2mOK9YyPYHT8DkgiaFyhPptedYEU7cmXOmjMXkQgNLPJ3XVcuo6k6MfOCwDnBBAlU8Jl11JTfyB
oxbKKels/bBFagS7KPqcN3GDeU6RILGaNkYR+sDGgRjljYLrRqDcdpxbqTZk3SEpJzdcGxCpVVLM
Vmyiugg08d75Q0guvAL+KbEwHN5OL/peQrD/wWVagnwLsmUswpdticD7nqoEwNWZ1eao7Evc9O5I
/NUSuWiuIE+ZRYsGeMMdxVjvDaDiTgQcPxbhL38QrQG3FHdr2QzrfH+IKOOq3oL3kJX28rNg6nIp
ATM0vtHGqtS0XSeUrnl1AGTAYfx/5IrrQuRxUvaHsVG191abLgGFboG8zPuomzmWldx0vbtLE3wQ
+xmsrouWJpxJIwJ62c5Ts/N64oBasCo8h0B4w+mXN/SxQ9Y/gdc3M4yIdVX4CguE48iFH7czccav
1rjegGcVYXcfIsuIH4OEdbIGoKEyi+VjT2X9AQUZ+FwTvwwnMJEAjyEx7+EatmTkLavh8Z2uH0ok
qt8xLqbYar+PmQ1rlAc7O42sITYV+qx0ITVDJ8k7Fr3Aaymbo+r/MOfpXjxIl5L925JpWxWcPyU+
q/TzTyJ9ZmmEY6ZlLDz5etPl8zdCkF2YHRdPDMMSFPCxZ7pDV79x7fShuuzMWM4doijCTsj+smPR
ESLjeO8yKzUPskLujpYLMOXs/eU14lrqkKSI1+C+WNDSD9A5S3+WBnPcdKrmzQ2t2R5injFA50V+
dL+2QSSwj4sY74twqwk/wRiKlBKAgXyrod8l2sZuwdijJPIWx91NRGA5E3+NV7bCdG5uLBcxYFGN
bUOzC8cWhs1yiG4Npm7AzBdqdXEkcAc5fR79ftirMqsqhNqEYxoYmSG100C5DSI48/wcdWCLLp5j
S4mH/tztxgSlWfgEowqXaxt0EecPURJkV56gvJh+kH/A68tgzPb+tAMvYcmAQdqnBAiFHm/Cps2L
/tJp+LF92nwESgA2AGnfK1vIEENMt46tTrj9OpArm5Zm0hFav373TNtxNzp5Iy8S+clnbtppZvO8
u14YH1+NWul/2RGWnhEgKXucgRzN8xLiyFCYs0ZiMLpVcupyRTeHp6o5/oFYVNSQ7p7Np/3sI/ai
SLgmY8nsPeHgmpDtjTvxLozoiPjx0WkKh3viIGUwhPT20Oc++K30wt/cqox6YcAdyMi5jp82QZQs
CZJQ2zLZhWHzZTG7BX/xctp2ION34hjKIcp68LyIq8/JvAT5E1KppwlM9I9p+WexkBJ3E7UUKWQ2
ClNbD+1hoPEMb8/2Xn+9/P+1dHN4Xx0KbJyjAsTKpcidRFJh/G97hqTzN1TAOTflfuGYs5iLQs34
2qmhtoc2vtlWfvQOZLwGiOdWEjxJjhmrglCIkhVMfLGXrsp6+99hKdU9Txu3Y2KpeLU24qL1Dha1
n37J1UwM9dHe/eFd1qrjxkIHPAYYq5ihIPjK4VevH6q8T7Uu3fPa4Ej72nkT36vEtaHyC91BQxLQ
5PN3Km0kUPc5uhGp6AO1hM5v9qD8zCYCdjirQpo3hD8rwL85rDIUfrdyoUIvQsbU2WpqhuSg4zV+
KXwfZNtfJHw2jm0IMnD85pPjnqH2FiU9+RPlAKJbDfvJIQ9w5GqyB9kmnItswvmaqVJX4Tq6j2H0
YsBbhdpDvAEc3E68RmsHM42bz0/7B0ehtHm0MeUyq1KxxmTvj8Y6QSqNNqJZKO0vzHXdw7+6mmvM
B5FiJDwHlE4ajinMqhYfs+o8nxR8XkY3cw3HdyCIAKoiUpLTu//WPw+xElhR8rDGCHikc+ke4CXs
FOTVRQRrVC5M1V1C9LRuX38FphNH/KyHcuk3WnkC0tpJmCoUyyJczOh1NDgrC98FRtF3Gp8zSV7X
7Gfz6oSNSAakUZAWzldOkH8eF5Xl8T66twsUKMF9n5wtuTgikva0uf68SKFYw4k86lclLEkLd4Xs
yiq4Ic33UrpAaYmFjh6m7WjbXacdKh4F8LS4tq2ScqogpHPUGkWqkHMEnaqTC02V67zjH2kDywma
NmWgl9fycz1dA1eT4B5wcGs9hXkc9AXr+1w4cx5FN0j7v9GMAWstpuGrKZVH3udp92o3cjX7WVXx
27VsnvbO5llDO+yX7/0M+1AogXsJF8pS0bbpCJC45v9VsbgI+KoU3zrBUUPOFL7KqeV/QyekcrkK
ywQ5ymw8KVe6eVO8C9pRawTap0R6vAV6QR+EM0KxUJlEhnWYwFMWRjcbew1oJUcf/Xcq/NI8lMgc
AqoCmIoN48ZORgsHYjvaG9fRTuZKr01W04+kyaAy/lNOjaryu5WaRQPk0qa1neuPeb87aZT97L4s
Gok02r+J0SVjV7i/aP+ul9EHetkCP0YV8ypvmETK7SPtxPx5sXWNXXjWJq1Xr4l8jzUybQ5I49CA
f72/I49CQYUstl3IXc6KHRDCkjDcJYy/rwtJIyvuRAliIcZuZP0ZseaR8NnRCTngaw52YO6gEtiw
U971zzSnSnJbSOo/uMf4pV4Q8661b2LuyIlmMnFUG/mOJZbtmCgSXvzAZd0LF38vJ5sDNX2sDxyh
qjk09QLavBVHPJqxPNu4n2vARALooRz8lxIzYHodhu4hULYHUa8T4Yi9gQxGVE5/O3RuU0Z7vv3G
C3OxostoG7FAaLZHn9cGTngKuw0PDaL9+z+WUwhjo0rvlYvLYewaO5sRZaiUCUFJMIaGPcZuR6o4
1yXg4DDnxgL/inZiRDnZc4gEBZccSN3P/k6UxMfXEdhyxP6SvpreNqR36gXkoWqDLLtTSnsqkWsO
TNwDSq1wUQ6SHNxA8WRmCvnOHfJaydHAAocNAQvuOlx/itEQ6UyErDFoKOGwKRH4xzUUwYvBnXJR
y7g9NGo8K6jieNcWFyHlDuOePH8UsOOt7UzVwh7NXJGnxOFLLRc+C3dW92g+pN8rcicbw8PIjAr/
ns3jFgzcTJ75ST+RElRwfoVdHK9+33S6+isCTD6zQhovKmAspe1zokLWXrWyszopBjxA7qk3qSRj
iBfWph+5+QvmLBGSAf9c7fww6cEDiTO+AzLKVSOYLT6VJLbi6+YwmJ1OzvvlWAZIHTAHMuud/KlB
YI7W1R4/9wb8Tw/lAf0sPEf1Fokzx8BMWKptxFSLso483sIXbdC6+3IKsyVDJlEOcxNMV66plb63
SnDHi46uZE/HML/bVhZcOJNN6Wp112dUMY6oXwnZcRulLg7lGS2eYWGXYCjBQXQs3B92J7+tNQcl
2GmOWHxz0npfkTTGmCUSDR2eHY1u0owkblpe17H45doWMNgCD+kLlNqqniDmhZMNeNkaVdUGUJU2
9fzkeHD/ELzPVhmjQwijThBwhoytDpkuyCZukxCmqmxY3yYaXccCqmPp2kZdm3OJ5mMT2N8mSgTh
RWMyed4nt7Ctwb70uXJRBwtSJBlSGCUHNDDkcvYNLMVDwnUKjvaBl2YBsfLDopDag2k1e6U78IEH
SUHp6OMO94ebpg4gpEN4uKrLC9vQucd6blRiEaCVS3BOCCK86nBGy5KO4n85b+fzNX0tLPhDRGdr
1UceucjwHOZFGXI0cQE7fGmJz7GzGKAgX0qejhJ2Br7XW7Hu24zpPTUPmwNbHxOpcf61UHGKminM
HOitMNMT8NYex77zXTOcO78OrhKw5ACFVnSXZOtg7pOaKzavxz9Ph7btERAACbqDtv41EEYFwtsv
HbKz8XQL3D742TTZF5gKtJ+CZKsJTCiXNNGJaoXwKBj1sarkRbsbsiOCZg9abdeSCh8rV1S7o0yH
qHSVDY+GELGBv70jUcUq1myTbkjRkHtAAUitdzyAFJvxXYIMrD0IqTVPFBwxLcZvlOf1k4C9MgKW
EVBZhlS9+9ssyoLN4lD0cMXvhuEdq/4hOKl0+jOHhotFR9jdF1UOpQSa+TAxmq7oiR20UuMbTAsl
rMYNhjaaiNX4DswqAaot/WuVZqKRZHMkL1poc9V6B+mhXpDNjpgOq7hzS/TS/fpEBxC33JuqhLMO
WpyNbXgm1YZX0V8b+tCgfL/Vf8V+AhN2dHtI+Kjqu133VNFzL23QRbXgg6Hb4II/7HPhG2V0n11L
FNFOamF2DRXY9z8qh8iBnQw3MgGA/VlXZ/QSM+1d509SsJguzKM78btYpMcbAhnKxV0SViRIADgX
HFnL9l/q/Qvpf6RmnFcqox4qfNrk8FNDdQ5l+FETUUtAbAX+9io+CkzgCLds2MDdn9Bm5pkzEVkn
blhRUOlmQ2XsUIJKwxdlb9WAwOLdYxfQTOfJu30b8fW9QwU89D2FFtTm+yrHoLnrEbw9FxSgrPTF
JYcr3La8/7VFZL6pCUNCRnsi462rStwWdRPuifSqgFXNSPDL4DdzBhLTRElLovu3G+DH2DmHWlky
pyGdIPXVuH7KASbzk4oc+2CPcCLh2UgOYbrkxnOu6tntysYevuPeWazLTGQZzW1PQpMK84V2Ayvl
1Y4MKSUmO12HhiDfi+SNd8B8kxKr2FNq/XoRdQfIVoPrjZRVP27bOfk/wFGwoX/Wf6Z6/zPm2W1U
diWCZpuejVTFZVSg2tH1cSEzpiMbGvygGhI+A0xm+D38WM/tosWmJzgGv805KVa6NsLixmr9evMs
gFq/mUkjiWvb6ynksZs2i9jdbA4+03euquj4xrwG5ic830ELR1uAgqMDmm7VRBGOyBGcMZek7FJv
7yMfgUNtBdPYyeUHON9piOQ6ozFZUe+iIPW7g4Gm1WfiBnEiTlSVDI8ViYi8k/dI6YbeiBgVl28p
0ZhhdDtUHh4BW5ukUQitQPROCIA74UYaewrObK/pmSUNNPQTiyQLmp5yNQeLuT475unMF7/kdow7
dz5asFrQ+1VmCV0Kn6W/i+uQsyL+WZQX7M1jjJC4scbci0Ol92l36ldDrcDhUzT5kBfFUXtrEywU
qAFt8KhZZIXl9VYmWGUe7hh63HpmzCy3te/V9QdBQEjcJVbUuVsQep6lMO+uPC/HKR05zSaTiHje
PpYfepiXwtchLsBYn5VEoqeMQSXLHg9M9Ifl8Ik64HU6hHvhhBFs65wetq4zjw2mNP0uBi3OIzxT
MLabJBxn9RvqbKbXjXc7b8sn02pdGqobLKEFXitBIt7sO9QSADAlyM0ob2iHfrMRDJudAg/JbH+K
ptJsKUss4wv+lUh2oyaXi+QNo2sfeso6X87NZX71mjkqY0KGeFiO0c7AqZn6yClzxisbidEb8fMn
s+K2Hp/uzaUo7QYNVdH02LIOO3nubDVKioIvNEB/LrcS8URpvtylhBAJrM3Wacfs+mUqSsqOsG/6
UCadlmhRxJoSLR+82lR5YtwP+bf24QJQswdhW8Tvvi1oI2GZkZEWuNWBX9l6si/wg37hKrDVhSdK
u9VyS/yoSl4Ernh31K64f8jBDMhfJ1/syl5941Gy0eA+wF9DCUs/fzpu+36TqXunbS5Bx3Gtbi91
rH5I0elNpTte/v75/OYvq/UiqlOqvI46CdMDWRFkS0nYhaxPbTVh9dgEqjMf579nr8RlJH0bqUNv
XzHVfMlSvh6jK/jAfboEKBxtLfs2owgK8mSwLEXhAE8m9XWeDUso8CIL/2PETW8PF4QTGQM5J4+U
f07bSxjp3Rj1mg2a3HPYLNfmzfoQYVeqmB3ajnO15pAXZllPCzbVin3MJQG1WI4YUCYyWUklXrUm
deAjRQAaTbpZghLIQTO/GJ7nXkJ3x3Ll+M6xDjMkLjkfSPhcu4j/H5dbMJDLFVL2maFSgRHApSLF
oqLoEyxx9rFS6CeQbHTaTgssY9NjvtYIJSicruLbqgpQTfU38AR8PviMgP5Qz0H5wD4NrOceDYUZ
DsLQ78okzymIxnnGL6FnmnQ8be/Ef31cKSUnhX8PzaNc7BpKcoXWtTcHtQsCQ4aysd+6PhX3Xdhc
2HMhb24AhIVoSAZ/mBZUzVraoW2i2AJw1tTkYIgesQx6dQ3qusYRP8AAqcbDb0WG6ju/FViaP731
CRhpnplAFkruEUlGKYemctXzr5WhguZgtWCZCaIK5mobJjAgCLsuYkP668YxrMlOVQ8BMO4OnwA1
XfF3iRUixv8t1O1s8wDO/3gQJgqJOJ8v+/yo3iQ/hkiJMcGNksgy2zAvIPe+/d8sbzPxAD0A6OcE
zKxJ5rcrz4ELsFyVZdRgKAdbX35+dSd82AGzYhK9n/XRM98XpMhuVQMK4mUKmBpRZVFBzHobgMXJ
/1YyoHPFcmn3gknrbeurx2l4epiNIlaEuw1uUrvdbOd/wdgnTYW/+wtVyW+5thHJ+ywbYHS4KO66
vqkjJvJMChOrU9bbAEOhE8zZUoIlRPYlseaXen0If4Oh/pd+qcwrrgGLS9RmFihNwjfyHnzrnDd+
eVipg7Ck01UE5WOFeOjUKSTy1QJ/LBhxifQjTaQ5UbJwyjzHvgRwu66H535DbLrY+3A9UT1fotMk
uAMHJqmse7ZPdQctSUqc36YhlOxuZtC7unJxw+OLjpP+FMNhpPCjSB6XQiOtF9fCm6QBr5qiswza
6roIXfJdcZtcLosqyvUW44fS1vdYC5f2f2xUixztdKfgfH4JzhOZlhiokAWppGWA7ggiawM0Cysf
K0fbYjAKHCmt5fJUGjahaK3gsg6XZbpZCbPmNKB2wnQL/3NCW+Jqa4pI/o0lE/eK1Pa2IdlT9w52
qHm8es8f9oSmD9t1gGx0WE/Vw4DBW93X1cyP3ZohYBL47wn0CTgPfR4KR/PH24ZJg93IVTd1wHVz
9mTAnXj9GSqHHqi767h3yg2f36JgcboXmVeYdC9NB0V0Hc9x87aegvWzSYojjPjfLvbvKtNu1I7W
3a1Q2JqgMGXTof7VkebbYC7d0YsPnpUEwi+vpWHguyPbj/iFaunMDEMDH9tyes4GdT/LJBOvCY7A
SBRaw5T7afTNJdynbFM6IB3KlxK1JEytTSdTlpJ1UMtRnaAVuvrBccAaH2lskyRl3b2BrI6fJ9+q
+2bLk0nrCJRoy0Qvdw/nUMZlLQW3s9C+v/87l1zFalz8oiDTq7yvepRBKcxvrM3zEl6DuuLrSk5f
/sifS2G0LW9XZ0MEkucnzd4TEIdelMQUVyFNA9vRjEJ1OKktbLntDEVDETsPeQWYTt/ntOi5a4bQ
rgspfTaqaVDdIeil7nvJRFLDE7OHYnFnli+gIqkSubL0XhJxP1SSs2Pgyd7TwLbKktrmvkja2rjb
d9mEZ9Dz3F9vLO3JfhudUycLWaksB+FsaJRzMlGY7vruZGlFfAYGuaKDMxGbymqxRIT0+c8khqWM
e2fhQ3+rjYCz6ZhdVolqDqScU/BPY7kruLWg5pk/1j+PKTxwsIF8RqLX8RohlZV7TlqBoPltKSTN
7dHZIXSZJibCRIreyTozBB68exfced3z+oH3uaVHblF0puSzSHYK6sLT+sQPxQsSvAhQXoRq4Exm
CInKblNkGG7QeDHPKBclGRLSII+HCfq2vxYtr9RYSyqp8YjEiU/lkaFYw1EV6i9lZiiaJGOkh2sq
G/qVzNvEmBo8fCd+gA+BBtRnW6gAvOzHGcc5K+GrkTCoI4t7BVpEx3mfJUfP+DxpkkyQ8SGEceRh
jBeq3IeO8Yh6n9shWYQ4Jlr8MY+4ZsCgcXZixMIJWTs5ZpcFFURO0O1aeA9D/uJ3+CFkRILTk1tN
vGFyJBRqoyBm3Aa8Yh3I+csiA/oSA+e8sndbVaD2lO9RX11DK6YTq+iCYg+MV19dI5C9odd80yOo
/Ytl4Lq9ABC+Z8DGkueUOR0QE7IQP0PnUBFqSZy9UJuwct83/GObMUOljaQ9TgQ/L5navsdT6WIM
B+NTlZbAPBnD5Qkz3a1Bu1zoaSv1SrDNRJZDNzDmGBFmaMnGLSM3Hqi46r8c9OPfrM4vXHC3Naqw
Ov3B2Tk+6RChmP+Tuu6JpQ5rTUSnPMbpa+kA5M7KeUxVNVIRAaNUadNBIGzxs7CVDQ5OuD9TTr8E
agPGj8WsdUDLZGJx33Ng79bc/qfX6akaSnUMt4noeFYx2H3ag7BcT8ZcDOqB/5f4LcuIpKhAR0P8
DZYqCnq1eSRbIcFkgkn0YDJW3qSZwffRINhvhujb/rdTSv4LoR+81N0D6OnJ2tGluPnwYU/2OA3v
p5eH4ibTr0f9KQ64nI/LwGwFQGT3EX0uMGQGiDVg2gjlYQltC0aT4ND2ot8d6FchckqTd2M+6xjA
nKPvuw/TYqU89y8WtaVxnAoUxsxBSW0M84r1LAJ9aW6pH3IYfyZqOZd7z8QI4RSOop24IkccKzvC
aQnx4JIUeOEbsTLJnj45BOaWPslStn/HrVosrBtIfWWEMqQs2qJrfQM6WSbn5Z8ZtsL0054oi5fn
CK4iJFYKghVLC6VUsjQ8WgcQthu9MvKIPbou6XePob5jPJWW8cf6jKZD2f+FCvpfDuA3i4eta5At
vU0XUngN/xmBjVmKvAf7Xbr4ULeagIa6ZnXSot0A3kzPHhz/ptK5x9BjFRuJf1Kfzk8AQtC4Sl86
9TDdmbMQcC01tlxmRahAcTMDvn61LZgvaULDn79eHtsSFhxxzCnlJHIXoWfT9B0p1GxtRwoA28px
nTHoIxU1yCdhp1TmLBVp4l3JCSvWSKTr7fePYzvCudgvrSktNyfpHyuLZ+CtQ9z6BuFl9uA0snX3
JHjnY/GA4t1WxJrVvFENQkOzpIHgQ1w4n+hA1M+O/jM2MrGR0lXCmO9bnQbkSFYhy/nXPfGpjuRn
tK+9JagTgXgajUY85d75HyzTCxxpBtfgYTzgEkI47b6HTFX6wluwrgVYnWjmxBB79hnT1k4cVRT2
fC33r2l9jNYdLQzreyOTLUi1uQpYOUiAtrZhrebTuF1eb/vDf+Q6X73LFkvkvoDqAdpPAlRNfIVR
caap1z83QNnUjx12QuEhkyRNFHaQ55XQDr6GA1LWq0B+b42fiZ4/6FA7vIiF9IdWvrB0UUtJ/m6Q
GaX42drcIT7R2mD9VBIcZT9DN9pAs14mGt11QUqMuzLL31k/fui/wakPkNWUcQxl7kPmrmU8zIeE
6BUrhostkp2ds4yVjNRNvxf9PAH7fCW9uWGNhgT+xtE/S+NW57h0dbWWSANuh+YFYwrD7HdcPB56
V9+WrOab3xME/HQ0mEgd7SLovWmL9KfJufepCLsXkUtelkmIrOL6BFfib7K8Ke6dqxrbPrFLPkLV
W4vGmQ==
`protect end_protected

