

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
US2mB3ZU2xYMwSgf2KG3QONmAU5qxOR5gFmXyP3MzegSXblZ76jq0dw3DGi2XivflSREvQG+tGNr
93kJJN9RHg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cVCcDe3dO8A3aQlcacvtDrMlOeMM3iFulWP1GnL0AstVpxpdCCRRxU3UHiCxbevv+1Dnaf6o7WxT
G4MiJBrZR0NZpyZrN6elCTa1aex/x1et3mJ/kXtaSnXZDYRGWgFlsFwFLktb6kdkyrjtbx1rPCM3
CfbtCvTObEIGzIf/FJI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ybpmXaWiA2h4ouUhToF83n5FZ6mSwY7i2SbAGhh214jlEV4EAw60pDdsC9S1DXRUJs2H5ijqRHjq
O6r3TnjNUgOULu96coukm/eTQWKkKJe9Aqdi1COsXCRXpY/qPst8iFpcYgvP7x9BLqj2FuOVCOp1
vBc1X163t+3g+Wnu5wdB02cYtsPg85Aym4KDvpdGC2+lcbTElJIi+JurCHNEVSPxn/s/byKj9Aee
BWqSso/XFdRP+TM7huy2D0efcTINLjUE/2qeG1Z2VdFBpyOvUXxDlOhNEr+qAiw/pCiqNyrHCapM
TfSbH498t2P5uuhd9n2zpj2CUOFq13OvODvHsg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o4nr3qLm7Rem+yVuZpGX2Dwzye61TgXXpiZsrYTQhxAIOttLQ5qy48oMqssSkd1Afuq4E1AgeeLD
pr9heGHoD5AjWxk13hv9r2YUI3BND7NaVLyrx7mIkF/pxjMjFTBF3rI5FZuYgxY00aftrEFjG/AI
XeOeb4w/KZQIUde+tJY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dHlANyrutuNgAtytsZMPMatpxiEBkM3u/gDZ64fIbSRqU16FBJ0WguNKCot1/TeXAq8CSJHQCt8x
3wxDlxfMsEEJdw5OF5Pn172rV07Ce6wZ30zB83ou1uUKjnNgy6pYqTworLe5Tj4SYl9VY0bcZ0g/
rN0niMih/6g+8XwbbPNRS7in3icwjpeqxdXwsRyEX3dbCrKVz4LXcfmP+ybNfKunFSp+imrzoFLt
cLJF8o/HdEoH/59p1whEdIyNin1+Ra+5d2hGnILLEgUP28LNS8Xr0dqjxGFNrkIDmtSmsmF2E1fl
JbLYu0fIIENjFn9nAJCzGQU523347ABwMPcyhA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5328)
`protect data_block
dQdruP6DW5S8uWq/FOvlskJV3Yq3ArKm1U73sManGSbYvw2yFK2/2sjaB0RYwCGQjThknNyTA5wJ
6Tq0RZdl4ippbmBaVkwfcl42q8RmOnyZIc0baMSOVZfSPrDk2TALW4qejj5q5m1wO4lGnAhbLjBy
tI3+66+A+0CzqdwLholLgW8Ymwi0fxbaV+CweWlP1zADsNJv4SO6SkNzJY/xpZdVjceOhQ9JGIEP
C4U1ExVvHTZPDfr/FAS2qhrsAvfBBskzpWexpUz+NObwUPCZyHYlAD0TTPt51FxG9jkTLpsE6XAw
Zg83t+2MnBkzrXzljMga/Q3DblReUuzssr0z4idADg+R0Cb4Lk3pJ+CoVcoDH+b27ma0Ko5llZb6
ggpZrvelqhCFbK7m6A/dpNCiVUTigpvwk6dQ0fBUcbZUnTXcwfvjqzLL+mKkmFNsxGk1JOCGKkDH
MccbWoq+zBelgOp+XHGh1PTkszgt6xUlMTzt6K4AlpED599GMWicSFcuPDbxQEJqK4ThZIfJZ0eM
NOL8oXanF/qmZhIk81YWBYO8p/WLkLMC/VKGYhXe8/5XQP3bG3Dd5qwGkH/Rrhd8XXjK7ItQ5XaK
8oKSkN1/5JgG9pVfdIbhj74VAtkROxaxjJKzXoc418CpY60sBfMJ5/LdTNRFnHwPrxvqy/ok5IFk
zyo45LHxO1eNZn1d+yvoX775pWF5C7XxSO1w5Uuh/Bvi9oNM+uiz2cR2O+5bj4cBx+3j2550mNjI
B92gQ6+IwjOYaEDhYepB2TBztwwwGOa3Tp0olIaXEqB31p2cTGjFLT/qWKKOpKalgOaowX5I7Ql/
695AIvUyRQbkZ5q+2a6iQuBu/NTKN1oJgGlVybdGiGLg3qG7ruoGQKYVjgCO6gmrV8ScuYozRdn7
diKhPHNKZ3C50ERgRIek/PZXrPbC9gL2o2C9JvCVpTwRn9bnm+bqker208+TTvEifKFUsRdtKZww
v7tqzobArBuYD15zbHfn7JRCvAe4jlpU4fe8/7rQw4oQgB3+qOVuJC4PQHe4iefSL4DEyES5AxBU
Y05bv2OGgaCuKuOFSy8du6oWZ/fQsK6lQXdbir+d8vwZle1x4vINz6AmeWXniuFx/Ed0vBZJLNAT
k6mhU9aCZP8vp1YpDEp2CV6YXKahWDYcfnBvM7Y610GLTvYLYy7RcJMmqNRdf3AA2iJ5jSXmsmXk
vgAgAFEqH1KpzP085GEIxMJY71C3gHrL6jBTwr3XC3PydIbbZaTkYnu2kL+wRF+Voc6WntQNmLLR
+meSpRCITqaADEbbANteWarD2v6Z4jB2MvBQhTG7bRbGo9T0DV+zq75u5k5b7xMsUM+4BbyC0r1O
ZmlaC7Hbk4tEkQ/cm/NLl0jqaGe4GNBDwIq0QeUQCBBVyI9W7CTOIDu/3W3coe2wbAIwucsFlTXR
iHAZgB0K631/xAgL1LyzbbZ6z3NbvJQHXdZVe6gjoIeWAnXbk5g+sw37VyrgYj8yvFQCMZvyaZeE
niU6AuDTNb5rVH0Te/pqLxrZ1FMPlOQls2lNSnJckh6iToSLkT5WtAM/4+qVaMHxjrjIOws5Zls4
UbVMN3Qwxsum/Z6jern7jKJ886Cnr7xIFEiWOLd+vxrd2tDBv5dBGBGGcwUYDdK3pTiU6PWVMgvE
51bJP4v42HeU8FYpFv9E4+97uAA+J5QUtmCXxZKGAwl3NX1GFJ9fjOykiRTurJYIOJ8/J6T9hDj4
gp9AGRvNORB+viMTXHjY90xvmCgNxzvaeGeJHcVwFylCavJdyUEOcmdMNlNlt/Y/8VkptMYUJdD3
EMkl+9/jzlR6eTLPv+nSeSWsp2Yk2GvYAvUcgr8aUszH19l8qra97hZno6Jts0W03gfieKaxFzch
CKgRjInoo1M9uq1BNJQB7PfGLHu9phDgDWWx4NJOUiHLwz6eiN1Xby6vB5O5uD67u4RP5p1jNvtQ
aFUunWec7r6YLCADR27BfGpZBU91kETpSR47P2CdzWqom93UDbLUS3uPq0Qv7OaAr0eS1Z39z2+s
9TPYOyZvFDuVfcznPnR2SOeDylkQ0+K63Po/e9unEuzLkk6TQhD892jmfcPa3x6NKPNm5NsJHNHG
La3gjyIOwshcQBik/GCRvu4z2xVv0ax4MSelWjWr0/J86ltpLIIoVAM2DHgHXjP7Fa8W+rZD6nia
igN1upj/0O3GFSzvILp5fpXqj+tnN4tlUAUcchwv8rAD1ItGd7hMw4Rqw7C+3GR77n0ExYMEWXpr
zFQKkZnUdc+zAtbNqXBWz7XNC59B3r4g2VPsI2Blcw26JtNNBfmW4GHL52xXQv8bopXrh6lFhiOx
Dpx45z4WnqBTlCA9QWkaJnU1iY4yuY/D2t4gp+cvgADhDOYoeV0sER1CVwmSERoFK5lXhBbvYrvY
+ct1HpIKlUvor79FVjPOVE2FuKNNDoPly50SdlOWu+stcB9e/KA57fwpN+OxwETBMaWMQiZqiRS2
iTZHR5Z/4OqzC4aA+k5WpNKBmtBeyOnAkI7uUin3b5x3D497LE8xSnEnm+OMxSLdR6RN1+M/B2zo
iEizPVpa0Cb3lRjxIPvMsK7tr4VCfvs7rnlcghqFFdd79Z3bq3qlg0udo4Q3bCUZgVQFmXH3COLR
ciDZySi33HK49C6Qxz8bWgW9vQu8Wq/G9EanolE+2B4H1LzXnEb8xm9NDlK5Fr/uX4o9f9vw3iJE
3+Q9kFYjfeMrR6Cpvw76Qhy/8SqbkXHgnKUEMYL4a+zX8qrPJnV+yPgBqMIMcVk5nmpyKqR21Ene
O7ITamqB0ZDS5pTdIs+JcVaZWA2mRr7Y0F2Ze+hD0cxYx0+X5MvUUnsjapsIRmL3lQzEfePc6egl
HCXinWeZZzzj1TXMZfqLlvkfj3imuouJrouPZ2CeBLf9SYylUDSIu8nAW/fahh/snnQRNfBWhYJV
jmu1olB23V/y+cxJ/2dTKXVqPjsiS9E4IiJOjoSeTsuY6DnoOHphE2m8X7p/m5UFoqy4JW9B58uu
/QxsFO4DQrF4bimMxHMI3y1HibgropdPTGelOMf1Y2ftEZwU5aZXKHRHFSfL/lAZkwWu4OAwzwk7
JLVPP8fC/qg/iY40+7zojmCdEEFvDICM9mmr/EwaXSw5FRQhYN4pi13kT/Qja+lwrVo7czaA5WsJ
XgxFeMRLkGTGN8DbVOrSIDy/64eoZCqSNn0iB55sRq2dBuQjul9wFxZ39mIWUiQPXJvcFc1YJLsF
nawTQ0O/5RxqRLs3QPXbjFZHCGbJeAJeGaNBNkTCBLo+8ObVfv4yPlY6oPYfXQykr38E7sDWAy3R
F0m7KmKqzTVc3uHUn6TmpuzOlUn9DGuLKqdPhW7jbZDbb/T1+mSVkugmT9AbKLrvV/QIycFcsLil
qpJlvkkcWao/ZYzgGUnt1Yz5KmtW7uTGVlJTy2gB8uOw9xMOq5dx7GCgZFO4kLDNvOc2drcrPVoO
hhW/lp1F6ZjBAclSo5+r4Si5F5aFJvEFeqHwRQc4hWNeX7/FqK4lekLEbZJD0UefQIA1wS5Crj64
Px9HzDqn0aWfDsZJFM5WwRUZjxrzwtJgslhm1RABsJUd91F5Zjl+IXS2EMsLF25Eg0blJuhUXYtY
j7G75vkGdE0vfgYNMgZIUj17rWLjwdG8YIK/jMbgPrK7Cx2QNz1UhteNP74UH7eI0/zrPjcDy+8l
/m6ar1aOba94v+YIO4aH/2exk1JUKKsPG0Epnr3bW0IyTevFcn9dH13r0SY72MpBlToyl0BCpoQF
pRQEEmK1T9gRFpBbuFuO9mT3YZzX1zMm7bfAFg7vrZZg2TUNgYcT0aus5htVOkIqRzCoTM4MLs/G
1WWMXzzazr9HKqDbQupnf4pq0lg0+t/c6RD+d/ZGd3ZOeCg2L2MOGXv98YlV+dNMZ7SppwNU+W5X
GeF0dP9DIJouYNTw/okeU6TF+vrPWdqV6PWBsTvTvqiGirj47HmP0dtevPWB0XZMyfvcpJU6ZVDn
s69iHbRlLNuY8NHd+wLCHtJe7o+0hfQkEAj/dG8qBzLmX0ka6eF+SC2Mi7hjT9hAidsHDDr7skD+
ouSCtrMqRZymznTAi1GE62Ya8q4Y85hjg6daxDUjM8am8BD7oBYZzD3SmboPja8PaiOQFgjDjHNE
xgkTCei6C9B5cC0aUxM9k6kZmfYC25Sw95x2WX1VtSS9AYyTQZkdbrFmvbIVpBXrWbXSiCB26OGq
wpIgqYHyl8F23ekQJtJ9rVIzU7bYVGYzNM8tatP3l0N8pz/XPOxSgOpK0kloWUhAbpfQLFEV2gCG
L5bq8oq5i0zD4bKQr+XXL4HJRf14MpPMPIQbxg+W+CUucT++ZSJfI7n4bNlHIw7HAzVDftXgcNzH
zHFVSoONAi+ZKmHREJrLAQgGS+Kutb9UWccnIfXY3R+SSeoLTdFnpp08YUSxzr45qJSJyG6zzBtK
GExBa3jZzj+SYf8LJUWbhUAGXZpd/GdbOtzLw6RSTAttvJIHo7eIoQ9GbzDuSdWEsfKpOP7t1tgH
zZKw6uV4ZrPosVhfm5TsYtDsw+ADXdANYQMkBxLNY2gCdgpcFrGhMcexSXIAy/xCaLB1QzSV6pQ/
LcFUOjksvdXBMiye91SNSYsaaNX7spCXzBnYO5I0QQuuoq0lvvhluiPruvn6qjzNpFC+qjXngtEq
Dq217ulg0Z3q+AGkWNtdNpQQagyVRTtaV3T+WFjePNl+et31z0jtbNTIafPRbDzAOwCvwZ5XoKj6
FiTcVKQ4XFIUaUO45JUs/1qiMQSgJnm+e5xH5aJ60bn+8ZVdBBtNixEUaMTso/dlnMuRuqK/ezJ7
qey6iQz8sV5T7qo34xgH63Ufgf4lq9Nj8hn9ONLhtDewYVnYFKMI0/EVBx+UydVUAueOAd6iV0GY
VN7e7D/iQm0H0HjOVs0ZM8T79/58IREgk8V5bIAV+nf0hGfubB+Y/fzCkd3SpzPBr0UHtSEjenVO
ZXPa6HrQ04MvIs83pcW80t5sgm4gfitxbQF5H2NXxvvZIQbqlpdCxzMN+yPdkPHRmafbZLGCt+NY
CCRIEX3uzC2dmZ+01n3dmz9h3WCz9xVpBhOGfQbFn03rdeYzKmX4j71Y4wuwhzO1HnJVdluM0Azq
Tk6U/LLk5uuA47lrd6hR9jpE4mS8dCueOMXyfA2gn97Hp4zi3cok8YZGWlcc121yIVWtzIr7sYhn
ODnvFrvTfqn92oxPv+uoVLcrmrlZJLnStZvwtLs13qds6rvJxiI6094B3nFvfRlOXzwUv3on9pmU
z5+nqKg5t8kEnzZlgTDpdoTt8ADfiyjYAI1PmY4X49fUNEyeVXie2sEs1y5UTu55HN/Xpm+Izhn8
kQjuLxho3SAH5zbR94tOppZr9gooRZF0q1M/p/+SsQJ5L9iMt2fe2KkH1HzDqXuIZxSz7LayrQZQ
zfa3SCn/rjD/f4CbsoqfuzsxYWXJTXU08P5dqvjS2Gn5FR6lktM021DbWRg51shGOdL/VqY0AzGM
i5CLOpcO4fgjFAy6P0Dyr0Z0980su+xT0sQKcFfgPHTzynRMWLBu/hCjroglG222oCAK8smfGhNE
WdsdYy7k5TbByaK+8klwIY3gbq1ZennnNXoIGwsfK+pc9xOt+YggVXwviArH/5FusGSHiWN2DpnR
d1bd97fN5n/SrYC840rpoQDc+7mEKflDOhbR1jxgQe38/WPn/Z1x3guQsIfVU7eZx6mcqiTm87cm
mRp8gXH8n4s0EpG501KYBzMgLu4Tj9McN/wPYYQoZvaR0OincwzCwUsfTj7ZF/cs4tqFxpOZIqIy
M277vTB7hr11VG8IJ6mB+Tb09fUfz3onI/8MIMlF/ocd8ricxq/58WJq4XLYOxC2wjKis/swwmC8
CIAAHHTPyHJZl5f8deF2X00pK6h0tyWPdGRxu+i8wzFCTk3u1gqwCmmJJ/mEdjcEn8lg0V3jB/3Z
bDTFFzVMDAkdkItiLbSFjsoAfbvtVLek6mJQrVsIVggKpJjuoowToui2YWfOu1jbzr5RR24rjpK8
IN4DYroUnlt37+mWbF+b0gSi5hRjnIfwCjK5dGcwmnleV8WwGLqEeiYcAiOVpCLW9R5P3NeoMxfK
m66l1be14Fekx8Dli0Q2D9NmixaTANO1seQtoMB1iaLSSA9GQ3kdzIfts+3KWju2Ucxa+67Z614R
VSLaPY2tQnbsPOaqWQvqKwmcycaFm6vMjIZfWpFGKIEeen9rt8mMyRewAKYCPTSD4vZnoNtzyCMs
R7x75b4zCevJhv36BUxXCXxMLocBFB4f4htLjYldBWhol3Pd7s4DLJHWByG2q2VDiM99bSqh1d2Y
xMMjDFUEBqcxPVBvJy0e3Ocu1QsYXOY/o65Re6hWwshqbAo/8VPWWl0RAzC99CE6o/eaf4QbWt7Q
dxH580P6OmUdMHV0nah5tCiL5DmQKH3SzjMniPm/HT5zALjFI5HQYKmyhWl2L4+9Kce65qWJk6kZ
KWW7SfTj3T1JXsdE7m7pHsK6Q403b+/sPhYYSQn/2+b04rbAcYLqAoaFh+PBjkGG5m4KE5ukpAZP
M15Exmt7b5cTVKP71FwdEpFRIHArjQHjVHpsGXqqDB1sW8CCrXVkkWB09Y62jCzG1afXyuNclewb
RfUTmwwnOOmLKt2FWAZbScEtA7Krk5QzIPCDOrtVCoq7XvNriSnEVkNIAcnK9LQWBrt3CPZf8UVl
6KXcHdeUFiCztyBLF54w/IdJhVvTy5IJ6oCJd+6PWn1bu8qursuv4YnF7jy9Bcf7mcrduKqODS3x
7MZTs0evmVi+CPG6xxrjvVvTdQmAQmeZyMd2HqrTgbRxfEW2s3rxg2hkwhgw9Lm8noyXNoMPexPb
4PZIDfJRRS98jDB1H0O8qEDdUfaOHyN7E9DGcetcq4WP/nxplDlNn+d+VI/EiHPbED9whvorBb9X
OFQerMwBD9e9r9AgcqexTG4Q/r2E0qaGRz3X8th8kEp0cf6uGlWqxKwqaYTpZml93N1vghbXWEtZ
hESKgA8gt186nhfnlI4fqHn1eDTKvP/Vg73l
`protect end_protected

