

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pTeL3lbzyXpg3zBlG8xXBsi5mPcSaOx7zOxONTRBSW321/dGdDH2TpaC43BqFdYZqpUNj4ng67vZ
qArBG995Sg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I0+MKhxg9FScVNavGFQn2xkzaE4/JyCe16C1b5v3ObJwo9nXDzI72pLgwgIfWMASSmFXtaAAw0ml
3uLnAPMYr1dgB/uJGeAtmT326qa5BMsAV4vQ1Yunxch6eAaFBVMMeEWawv99YiJK9jkH7yDAOpb6
smI54SxBdohXuGVE7bs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bDMpPv/P03hJ26zOMeRntjG40FHNolyY3dG2sIAWSb+A/C9vMJYUZduiM8NsMGgn92oqltQI8itf
kfh0mxfLeub+eu7+DutH/IonvZFuvU5PDOu5gXDe5IZcX7PKYSeWlg23QrTg/K5l+bblhZE0trh8
gSCxX9Y5M/tKkk3Ah7QmsxFm+D2iD3pm82WCrtLPh7JqPCGwGw7ZkIH+rqgZe/fQHahkffxj0VdF
wp7Pe3wFKtUoiMTg7uNHWsoKi6g7a0GVmS4unE3L9HQtqDdu8p186XHZQqxkv2iNX9KutOONjQNy
x1JPQknSlGZ+dd8WmzTlL9rwhQHGdMhFcdrMGQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CqlfcKpSPaBiicqGT47t9PnrRSQ8njMbqaZWYqvnT67KXQ7fxmLQJl9EXGvFoMEq5tU8J3rLbBm4
9pWLf80+KgxXgS9WPEn1zRTKt1wiye9VOUHfewp3QYM+B5lPR0EENtCdssVC8DxPUBy9Aythtbty
2YxNBkGFMjMRSnj+A14=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jiVIVHHI1er6oSZsM5uji5FpVlbZFUX1C20PfTXKPYBzpAjDWZhROWc8xFgszwvy5guzSmUMWOgw
XoJ7z9N2ElsO0s1NH9ojznzy4rNB66tyJa27TZfjI9UYZ/9rfTzXHnlr6WpUX3IChRrS6x5LI1mY
orERQz81jyLKT8cB3O8KkjO3g1Ks65ZIeY+E+7T5cJHzOHJQcoiTTtwLajrQktJS0RpyUJr3VZHu
CSADq9QNuiNkf73BoFHvperz6rZhWbdV5MnpWKfmllMNlSqFwzZuWbMdZs7ZNbssXYmUZlJVjM52
JpTXdo1N5lXyKjXVvDlv7kCHkBmnfQZM3rMXlw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17184)
`protect data_block
1epotjln5FK68YQyC5Ii8QGZyPc/Moy3rb5C+ujuQbWJidlFcPLxBUDaoOCXO34uV+hhmg6hSviT
fsLFVScs+yiTi49IeX7g/6IE40BvNil1cro+diO/+v1Y2XdNYIGmluWWphxszVxyjBPLWKhFUoBV
gQ6vBA1bP5CooAWDAEikoeE1tFOOHdmLuiLykK/4XSVjLorD+YgjhSjLy9Zc0bt2cj7mWgzr7J1r
9nBs/50Rba/Ou1IDqk030u+p1h3NAdGRhg7omNVY1pgUYK/bRXVHRDWo0ccqhe4XnB+PBXUwKO2i
vnPtp13wxmDWyzJ4jGTeZMsfIg+Abt1woiZ6esiZe537uRxAyVpYY03xw3gFhw4IBGN1oDeIgFcF
rk553mihjt4FKWFMAyuN0Au0MCjso9nQ8AKNMm+W4cVQg5cI54q7xB3T2mXG7gGkgDMILL1WMjEy
quzpoNVaQzGhz9o7ln62KtWeV2wBKzeiBj3N28yaiOWsr7kVEc6V4w73K3+YPqPCoQUZwxTIG97g
n/BX45rCmrJ18ZL2r9WRx6TIW3rzDJqmU9StKwERktRauccDk4RvGOTfYSDuaujKcxqZfGNGImN7
DxImdNcHHN8siyLO/bET3CixJG+ufzvqq8Jklzfb22iSrba6N2upkkkOk0WwbSqVGTMjVEXiN7MM
yNBL6GtVxrqkJuRHjmrPx20PFF2lHGJT9i+E/zGBuLu3JfaZpZXv63i1Muqcm6+Q/7KqZ/otiOPv
1IYx+18oVhqi1i+MgyviVWoEJQPtxJEFrVXuNy0ji1w29v5ae2uWeLZCFbo3OR0AoboQ0/0Hzv6A
ZwzQIscZUEn8U1YFXvvvxTOm87nfoposoZe+qRBOBsxRNEM2snCYrj3SMKeAqShBRydZU3ELnkoX
PsMHo7mh/eJsu71B7HGm8vq8aaB1c5zyphd1G7tQhQrB5+w7Rd0RtuZDuvqvNVW4IgmSICUksy4C
xM9tBigInd3Bt0+e5r7iP5PZpL7Hu9mTiGf4GDGsCB6//e9q63MQKTthpS7dsR4s4VQ0PPIplxC0
P7u702UuWuKYSuqhKlYy4JjTVt65fstt8dcVSMT727wWp0gbftozn/ErtLTExGwU2dqmwZYbIziL
SKBVPSwK+YoiqLthBUuyhl4BeeCvqPnUxlFRo4Mps/VVsZ7iuysVjTXhH4wh7EyyOSYGrrNaUvKr
Zpqt1UUCJ9BZul8uVGlv3l29ayNH1V4vDnVJaVp+2TZTP7+2HqhTHvEDIKs5H6Q+lhlYs4/aMcBL
P4OMG7bFpmi2NVjyy35UvtLQYKUSRg4T+2eMXYSQ8DYw6Pm/xJ/PdmATT1jPIKYF8v96phBZ8uj3
cRqd22xB5oulux04QTwQMK/beeAM63IJqAzlE/7vAGAPlCwoMW/4VloXNgbTo25HL3Mphpqdb4tj
m9mvtgFm/RUAUQBNgUgNRcQMo9/rreWTUz3OdoQT4zfSCN0Gql0T9fVxniJmAWe3kCdGk08VLQfy
SOqlEh6RvqLy39kTennzw544IZBcfPtScm3eUiUwwl5187sFWHqxHytcKZKlBPtf8sp9VOxd1XEn
dhjAcut+34yL1suIOpEdk/rc6LqtZDDMs4YQprhp3CIBfCPGjFJuRDE3EDKysl/GU3ts3kbFgt/W
fqqwnPb2zf6wVutJsqulC3JQjPTxFCHDHevA59POwgowckkraaJjsuTiEFrIas6rupa/fSr8K7C9
dPbhuAW12+ZhEzQSs5junTlkgsDJ2+XDBXHXHwk5ukOpnjmWsonVaORwHYAXPHBS93gSKg2sKMVM
u0OgvIHN1sM0hpw4eFNQR+O71TiWwvmpo+Vc5zMmBSlr3q4Muu7g9drGSLaypD1E58GXxbxAVvO0
hxKwd1JwtgkiAUs53YG0am5iYo1fdQV8YQc3eT/r6IddRRzH2IHiyzqsJtFqmOeBC7rweCXgM2GZ
4OM/NSBRJae3bX3vlO3vhF1B6fjvkjGweag9RDKp0HQvYCgs9rmvw5WpQ4lLBKr9u4aEkXU4jLP1
74QKL64iIRqxqwrjjKtZBWEzco6qhPniY3H+YX1d3UKAEluQ0YmhujuplPwIric99q0Wgvcv2XzC
N7edv28DQKBBsAARI/NXRyNk55pO8A6Jbqqabf7Xds61PGh5EzAsY68ws03uUPIix2SykISFxMGs
33V5o0ULTImv3902yxkkKq1oTOzNDS2maaizxY2dNGYXu8CZQZS6xMV8QKPyBwUQvXnxR04Ne2DR
zJ78WBuaGXjGge9AkuIzdilV8/9BeNAz2pQM+tb9t40dKjoULybKUxABgJD9tQdEION8voT9frYS
vU2f0/6ACqH1w5IPZuc7hcNSW74dXEJjStK3L9M+y7tioL0dcMzn6gzYAleHyXiTaoV1tD30wY/P
QO7GDDioSkflyphpMgmCjuxb2ddnkZuZTWqdGLWdTaWD6ZGaP+wFtyiaEboV9bjodI5IFbR5MHl7
E0lTY+3o+KyXjb+TGzdfU7OABT3EB/l/DcMN3ZVr14HrKRgKnInvkLM1yu5RIZ01Pp1hfnd6MpLX
6CzN5xZqCZ6fNFNDNt+XPWqS+zn7VO5IDvNfgeEUECXqzVyJa0j71O4/+x6o4n0fdjlRzYhIWdI1
XuxblVwGhKJu6HPQ/NqL77DsKPRw2HbuNJAawIRHtTYcmkyuKd1xr+6l9yc5nbSCZFNwZs1tfeKl
8Rh/kQXhIL+Ne8T9hcQhHR/cp6gq818272sgd1y1l7S1Hxw0o03XjplysJNK0kl98XsdUdZeFj6i
qxkP+9dhFEaINunVRis/r0WuKtqIrS+jiZLoEZveUCkJZCIz1xCaKRUekVroqNe1aU5jM7VJuxvT
SxBdJFri5qfaHMfRIBR1T0PpadD98HUtBkIFz8cLlfIb34k/VrvDmzEzHqNu5PcgkwuskKSfyKAi
+GRddULpfJkDDMOQLlEWTtAx/5YLf/SUrqrJmhNZVo1UwD2CHZunp821kEp+VrjT81YUXf++0HQ4
OPg3NUxN3WLg5Qn4GzZ1QonF2JF64tHTASLY398xI+JivW3USUJCQ6wLydbEW47LI64ro5VoEXWY
zg8CB+CXzDNkkp8PAzsVjeJBQ6EVP82KCt/hEdYbxDTyK/K+1wiNfIrQj1RuLTokkwkgZ7Aob4f/
RT5EYkSbRzCDMSCPw8M5kvyRbq68+WDMdPhqBPrLYgbO3PbKOy1Ydyc6uDSXB0xSVNeUlr52mFvC
pKuo12+6zgbUf/F/fPcTNyb+0/wXnRSZrB0HAmJFxg+dViIVE+WrKtb34nbABhSce0joBsUOzFXG
yMX0V+jiM+J51dowFVEYv+RZsKyEmdRp2MEZouB7Uqg3RdOpkGGu470uf962Cg5dZL6oqyDtYgdx
GHv2YsgVI13r7PFVU5tmXOEUpiTDR9674V8FOBMNuLSKIwKioixuaW8BWREE2yhBImn78Uf3x3rZ
IU9YPLJsJADs0k13PBZ8hV8bnO51/x2ba0cX6JcWagf/QTOmT0wNe4lvaglCr90rZqQ7qDnCnobs
sPu8RA43VD7a9WTAhqYbS4dSXcf96msEJIZr5VSgEVkw3GfHmtaIeU6T9FWuKTlOn0nOHrad4/7o
/hsP+n35PysrYpk+TZ4aXwHTm5nvCpM4Z/c6ubLS316ti7CuPjT6zCX9RtboUfi28jcak/L6IEtD
z0eEfxihgI2VjQLzZcSNTLlTAVSI2VVQSet2rM8X9uI7BeaA3sUb2Voou6ENkuHy9PUx7a4bOExF
N0enrECbJbc9alsA5U5/VfnFBOPuopyAUHWX17w7Pg4ufaH3wyrsqbb1Gr51YD7ZBGNVAucBCEAw
WRO9HEGhAIBo5J9c1zSM+1lb9ZEok/wlQO+wQdxG0o/lKTSKZPAkBbLyvg0NNt/WuA8rWKsMni9D
CJ/9B+81Cd/RGYwCnIb17eU7HQWY+8mVhS2gxko7NZPgL8SZjzreNupGwrifuWbvZ7UyuyUfzB1N
orWYdeJ8E0k5H3bIQA0/zzcdf/LB/evE1m/LQoyaI8ostcVURBZ4SLpjiH0ViZhULACKfs1cu257
C9yNTX4hekaMeI/C9Hjx2wITeuWFgEu+mAdHTwi1jBglt4n4RMtVeGZzK8dd9xBCuGDaodXAfONd
Z/Km6gD0eU5eIiIAtD+kdJXdc3EYzUz8AFC4yqNbLbhH5BCGdSsstiKlO2vlUprpKsSHO3JUC2YO
ZByJ4fRQcSfhciK5DS8nD+uUW9Xveo9qYf/kCfKOZrspZkx7HlRba0fEAtLH+EPFHOu4+vRF6xxt
hN0eny/SGbE6gdxkHpb1bW74S57geDzjfEnUTCG9cTGTOEb0KdCkIXH+lm2GtpFBzja/RuRoVkL0
XgRJ6esm4Hec/YExOF8h5vIEK2X/cQUum7FtDL725QThTIIqrK/skE7tyx88oOBtOKy63BmP3+9e
KcfiOl6uQ3+vc8x+apcrENJNi6lNdcvQg4JMmNHA5sBguicsHnNvBJ9C1Wjv8q8t0sdiTobQAvtQ
Gm8rW8QwGgF4fGO1dY26xGk1LO0megmEXOgrEJohwEa3JqW9z1PUpbV009O+Mvql0leuVtr9V1+B
HVgAEvbwX2eur1FRkLV0NPRQRNSaajk4s/vHcJlJFkUVraGRDmpu0ZjBvvgXSlB1qYpdoJVhTyTA
dAIVbchptZHSZi4Cr27MpzpoJ6lNdUj5HARNAACVUsEqA1bBj9Y7J4CMyhLwDzbp/q4mHMPIt4c5
yFSaNzcEhZ60L0Fdp3OhQZCUFCu48qj2Fj5iJU269HDTR3bhCepD9+Y3RMngRNaTdPqK2ZhHV6Ai
o58mS6PYA3fZPKe1wzxJNPfk71ao3rJtRM84q6cpzoqk405n8nvoTmFoVcqT3DkNXKA4gQVsGFCu
0VTsQX+UA+at5n0j2qsSansg02rMQHIvij5bTWUcqQbLAZXXF0oGncqPfFh8iO0v3rZZUMmW48Qo
XR2pwz1Oq6rlEIMCUB4YUnp4aTOTXxLILN2p13SjdUs5n1/EwhE5DVJYsFINrD+jreNl4Y5B8j+1
d2ameeXbksbF8NRN6+n6GlQwjM7TX4otcWxz2hOL+xlR+AjnKiQhIB0v9aIXSXKDByrUaT60zelB
aV+5Vs76Wxky5EJd7FQsItplosm8Rne/o3VYVzyVKITF+2WJTr1o4GHCwz89mn5MbiYb/lIviiWi
F/7WNnwQefE+PqklQP37AgOea//6fuhJih8hb6+1G7ernavwnuAdpEN259DvHwLoQneAo+pU7kEr
wqYsOpeDSe/3WBhWfVtt+GYMEQpW6nJytE0JCFfB7e/DNJEQACAqc1pIzCh19KfI1H0DKe6vIIC6
0JPlIx+V+/EBI/VoIKx1GcN0dWvM4d4p8v2QEC3GliWPHZ129iTOP688QrzoxFTfx1PszBHkh3Eu
2V5qduFCQn2tC5mZ4gmlw9jnhYIJmfhn7aWUMDjmDYHY53l/8Hagn/wUkUUQSXhRrJBNhMhHjgXS
tMqJkaKbRRFVroHKFzNBmxBIaBl0LUhZNNnQAccucGf4+D4VQuOlgHYqRk8/WjZy2k+DmbKL0RAV
4CsoS82GnWonyg/t/j6jB1bsTMLcva7rigX0viAMMePZLMXswzjfns2idOC5c5YIU4yo+A4fRA2O
uAEt2ucPtfv08i0lJKQo2Pl1/iiLRfhDM3omtrrOWTdCDGHoRqmSBvw/XAxqK8oaMDbRsHspwAm4
3kOUDQLQGm6m51qQe+x5ntl9eI1vBSU6HeUELmH6EZ9Cy/1H4EtgZnOScRToTjzLvdUywcg7Ir6m
ICoTV710uYDS+EeqW/li+MR6FFkVdVkWztEiCrCClhek5z9gwPRgqGeA2VoxWHPsNcqDCisWh+jx
pHCTqkWpmGolSB4nr7PU9fVmhlIGL60uR/xAGaXpwWbBivQEyZyCswZPxIAJrIgcCU9Ng0CqnAyL
EEI07dhK1y+BiClhF7kS+jLCjatC/Cb6zDU5zhfl4poaKyh5MteWmKkOSX0a/HFB5YpGJzlK2glw
h/3JDTJUQQ0VVN9kr1BLklQFlkHmt3y7lMHnrRHQC8QMyfj0LHLCkmDs70akCjhPLzdFB6QQWH8O
6xBd5+cB+IuqCDoyA4FE2l/0AxFLLKifUvgmoLT3G062ttO9Cpm1bGXK8ESTDWJIKy8qkATBKbmC
Yqr1ncsgfx1GLOnJQq2i83Gb6Z/BOO1owvyKv428YnaRdBDCKPCK7ryhWM0JRS6bzi5Oot87uZrf
2Wgn4EpJSR/RpyYMMJwXgRByiEoTbvDUSA5LJU0gE/D2InJ7zdNEpiTJK61ue9ohiJ+2Qaxet0+g
DfTLK/ZzfN4ipxqoPkC7wK9NZDeLh/VHzs6qJeC2zSoO0co/M2tBAAlQmmWm4pqXFUI5Kjd/PrZm
mKrsLYF76/jp9clHYIUlbofh2PH4gRB+6MkP1OwafABT/+WYwW42IkMoLLCQ1owERBEm3fAgOt0D
mdcjgM+v+Ixgu/cXJgyrhgr2gNmBnW9xVWDsujkK95HbsukxJKet5b0YYFAbyVGmtvjh/cS39dwC
24o2GjNfSC4uo5+iEbNRoXWAlyprBYngL97TSPax1cZEJPHuYZFfCCTLzQgrdiTzllUl+5VscK+k
XoeE6euapa8FNXkZ9PdBMqP4fwnFHzDy0AG8O3XSLqsUM8TgB9zKhLeMmwW4USfiu7ArPc5jjRdZ
mQ8+pnlPG5TR0oLc7LQVUH4gEL6oWHF2UTjedCF+Ut3ws/DO+6Gd2KNEam3X6kTmFGPwBverco5Q
Wzhljm+XGNDwvS+Wq5aUtz7M9sqAJv2+uBEaeotNlpPGX6prhOe9enfXQ2eOdJDpDvPP7OT5jvYO
CBUQnT98lKM3T13jwWcG1w1GbEbtsTteJUR9gIzKeAHLtbxqVZdr9aCsJlbgTUyc4WGO3MdUUy4K
aUY0AqnPn7VDOPOOVx9IA4Dafl8V7ymEVbuacpJRDcnqY68sRwsfeVjiUBhOEYApXW6sq4c4zF/S
7FeSluiCw9pqeStkodpi2sFQyC8uCusoFiEGRVmR+rchzbXsampN4hyy/BeelYombfqpQQ7wQONv
Gq6Rm65uWwJCzHFFaqilE41jkKURs/lF9GjjpNW8UGfJTWZqjBDjtyQUAmFVK8GUIAq9XSMfeq8a
1G7Hh38uAOduVVvLI0LeK6wywtdV+wYmQ2bAip/NEuYEf8waV5bTjBFlJ2FN6xmAzdL2o70ZjFHf
B2v6QLldDnUPievnjlvCsf6f95vMzXOUvm4O0fS5lVQxRl086KSFIza2dCadWo6uYYPYJkEfEsa0
XDWooi4mIKRUalFuOHpphcocfnQmTJ9MXfs7h2iq7DX8YQ/l7ROMRCXjCuw26p/d7Gdgna/VECKe
Svj1TS1blR28rhlWL52hfpROzmOu28K3PMoO6L4ta4cT2jv793Ft7sYL91Euc+5GGH1acDWjmS66
953zuMlOgSJ4vDzfyWyUB9mxsKc8pOWp8xBSWJKvVYVqkAIHbsE+dwQ48BZ9QNksLKLPmHYq7ZIW
7k2XbLt4MnHfZic85BSjDpSm6oTdEsNTJUtCEBqXKk5KvvWPXZjrhM0VD46AoOpAVgddCVYh4Mkf
mHNfr/InP+aqhWdLue8JaBPxfEc4rqsCR+A6sMSKQz+vcuxZzqBlwsc1/E5wt4hSjDjWJiprtbOa
mTrcnS99N8Qb1STlbIR3XNdIBuqlNd3CAIe46SGEaCZI02wnrdhDmgRr5ftOqqBgHEmlh4F3aIjE
Ts8xfFircxRqKDzhGpQ62ruvZ9qFlkp1CXhBbt9aKzntZAMbxQjtXvNbT4GyrQVQEKVM0ctxdDfQ
fSQ7YsxfovVVu06BMw6EW9F7FbvxfCHeb9OUoshUSlDXcGUZDUQC/RP8Ytf1x8PGbIvUfV5hG+1z
mlnKsOmF08vHc0KSR0xZMWQh4nLG8rNBqXWMfbIvD6LHoB7g+IGoYfcY1GnLpF966fH31JdSak7j
YwoqiYjD6PfbKmZWCOUhg5sepWIk8Q4lx7UWt46exppg4KAZhLZUNS8xwPIxxXFHRqkFm1cwole6
v7c4jqrczzRX50SvPVsJluueWitwGUjCFgrTktYpaJGUTZynfxoFZlJJPKC6dSABfsZz8UP3O0UK
+huwc+zWt0pYmEWmgH9L5b64qzrAaXY880RkaWooADRQI5VdMl324V+QRS6XpWBxHU/FXkqoefRo
heohpu0JCW/ImLmMjr7ZWqgFtoe2T/NjAtrbRS4FLBRTLSF2lwatTcJDuC64gQwimg3UlKouDNiF
R1mwd3bBbdzru64EsELsDbCXvqsapiJonWuKWK9l38llNoNJz0VvQsm1XKo4iU1eyPF2XnjdnJl/
KupBji6D6UcQ/KEK7wWMXUFgrE30qu1dIobWF/fu0bNg7gz893RFQFUDDliA2jRahhBYCs1FjDPW
+mIn1Oi4Ljp6hZ/K+00B7BTHkW1t486Cf7nO5zSI9alND7PkDPUm14AMXIaFMUlrzKyEKQ4BJePD
BATK2GbPAn7QKikRym1x28Slf9cTzsreXJptx1/PKQp89B4ddHVzWvuJETA2a5q9hlPrve1Yv9SO
rF3SqbMsKFLG7UcQf2vYdaKIu1wcTNzKRjoF81rioyxiK1tGaW4wUvwvmG+/tReSDHKZlndfKPOM
KStuhJf/XzXJCMG0OA6S7JFzfRzEcHUbvoqkxJfmdBg7n2vZAmoonV1DnoH1z0fMSsMjV702zvM4
DpZN0/9ySTkKF/ZMkdfcB0xMYW1Euof6+DedbSTxvmCnwwWayh0b04OH8+rmjQ+gWi+lKh4JGlK3
9KsQEJs5ITC1i9BZOkJ20NVj5IUqqo4qZZ3ZGbN3o69HbTVSDMPhMPACfqoDKV60bnW7+zawg6Rp
33jDc+fhN30ECMRXXamX+pdQynauiuHFZz5tP+2lDKR4vJJgN5Ye+1SRxy8QeAnI2mlQ7oJfxo3T
FVdm51ooMlrT4XDQqx6x5uHvDDYTRJVY94DjSRpFHEH5A+uPzrUdML90uELl3f3Ffknkl+Q44Njq
v+okgrZ8MLyMD/cYvGkYbX16RIW4ktBYQ/E7hZBMzoKzZW5kMJzf1bHiy+7ZwC9Kbyx3l3M5K+Q6
nuVzD4zzo3CBPvW815bXouVHN0ZBQ9w70Eo4Af42y7XpY5OtTtX/SYGYCPFyzosnzFB7q6OtL9J0
MWAqwdOb7CKEcMWJQ550Ot0gAApfoduW+EXKM5kbYy/w0KfesHoAOM2saiaq/m+juWAd7v+FaQNq
wfudwjSnO+B/AbkwNePuWuFfGwrMDFhZ/Yjodtn4PRKD9BNMDNURfs6zKtIHMtohVJ4FWDA3wTuQ
XlGaIAK+ZU8zoFcXckgQw73/tOPaeWbbW6710gp6rt7YKSTPZ/qJzXK0dHZRLnvUSoFo/le5BE6a
ef4/unilz/KiknO4wyBGxD2hquLG+cevjInxpw2vu9aYtybpdcnKTaTQWcEkvqAHOBjkXSRy92nv
lxDY8f3NEjwJ/WFcOUPQpE8Hi9MWiyFV4MlSiwoeyA52Wduxifmm0BigDP/qN5KrF6tJkZf0/LIc
MOJsvt6JIgIIlnk86Spzqqigc+uMcKqYbeme83HIRo0ei67npHVf4L6HGVsMCWtc+kHaIt9S2aRF
eAmPZ73+jDCZX+CK1SmZEub9zakoUh8ddNRDILyIOkWzxyibK3OurrvbitN0XL3rckNh6tTZdD8a
lHRjykVLjyMouvioaBThdXojergZlOLg9f+JeyiWQ+0Z02zOavTREnqX5EabX3cPjAS14lDM3sEc
IEY+vGOD04Qt7b4wPfxxguEZw5IDXAO1bbQ3HqP7ET9G5FveRy3K82kL/tUHgcTKM04U0tHlz8TN
6r/2Ru5eS+NhXI4eO3DRsHDh1OYY8GIOLSz15g4kHSFZI0kKLN4gUQR9VOQuwxYvLcoViwQx5PJN
Kho7RFgilOkm+0NOiCt6zxxmJLpkfUtidjd7wB7vquIGCyqiSmI8p+F8t1HKCwMY1EpX2z0O83YF
/U5SwyLKD4JgXl7+hlDZbQ59ON6GYuuT44/c8k23HHGXCISTm/zSjMc2/OBQ1XM5YGtUNQNUkjE9
W+2na65T2e7VtrK4j8eUfmXNx6tJo+cOsYYUpejamJkjZaH48pCr0r9EIn3I6vDOjzF/H5xkvUAe
Yw92lL9NSC1MKRu2AD26CezmL3ONrYSczKjV6UNGQrte5E44UUqXXMGokeSxoWvq/8oVe55uijWt
jt7rkiP4c0YskWyAZjKLleMEmfjxqt90q60hPiggJAyzCYsK+kMl8TOmjPWHoyqfOBBDP602U3Fg
i6QYaSJim5UhnZjb+cq0Z+Ww6JK/5hNNlX1SBtqPjvgEyozgUwZ7Ou/34rrOgfloCdFioBQHx6ws
iWpXxSrxnzf9IwncgtGM3kbZaiavVhMhqD6zyDrqGJpNKaKGsuzNuyCniBCcGuyHGzaKJY2UA2TM
POk+jpWLLcBUclztXVmi7YbS+OM8rbGKTAsFHW6S0u6QJII2rMfVGJTMvWjX7szLKUwFyIVO+eO8
cSXpAzLrVchXXjMTNBPxekh/Sp4YcKg66r/o/9Pv5yRFAMrDMM6oYzFLGsHBToD0fBZOEEn27Yn3
40KZNOxbdo5HYNK9DzsiobWLM7bbJryLP7o8u/nZVHWAmrk72fcXivYIc2QdvA1qTuSVvhSHqUIP
/hIvJvMO8zK54NehCVDQuGcDI4c+jL61ErIw6xjOmVQCBMp9Em03LMxSHBcw5ifShKUFUJeMwmPj
Jt1IiopWgjZ5jR2UnfNGuIjoI2meWt0MgHigIuug9itCE8ncOF+2lP+GNX7mxvUQv0bPhHbZaKfK
cfqwhvlrpTMzrCaoJYZsXK3kMIwYI+1lMvhi3tb23U1cBrorDudJ66pbYujkcl6496zHzAWwHvw8
2+6jLdc0k5g0j8AQbqqidNn8HjymNflPtUm3Uuy024xkxCkX9E8u2tf5NZN4ifuybT+35BjnYL5W
QrQMj/j5iw0JNujJ+AWJ8CRAvutOx3XwGQzqDY/SjyUXv6KL4H+sJ53f3EEFncw6fOxMaUZSFSAE
6ObQHJsUzJZSk5+6OBee/5rmMykJOm0imDW48CPS8z/4hjmJZmNm5pEmKRQVZvYZSUG9dY7JpD6Y
dFgOF6bCQByVOB3AMD1wX5vZBe8Xjj9SVNQXgKhnuhoAZwVbtlwQQaK7/L7Z85Lv8a/KUSX1BfbY
TlXpyVjKT3itas2MdVnwcgLKDGYorrtwgAUvwRSPcd34Vb/OvsTvh3kfwtd0zitIFugSkc/fgI2E
dz17GJ9MV+qP135B4TQ4Dezln+7kxfyixik+EEYFWKXJLs9eaWuCcF1PzQRtftvNORCWPmu3mBTl
qHYHCi5/loDB4CM9qks2zbTSir4LvaJcrAHOgjuDmDt17pjlaSn/8F46rKbhIMwAc4AQQ/lng7iq
uLINezrdS7BpUOJYyHrP+O2l667uROen7YT7C9QUimpvukIdB+AQR7ZOHyy5WZJyw8u8uZllZgeh
6B8QWgvOFytcq6yx/P0MTsLzvk7FGGXuMpbmY+HSZyRidysrCOkP0lrI8AnWwlg9DD11l+ECGQel
DwThUp1dyB0Ws6wsAgFxPyTIL+FfLFwbjQW960YLTbZ/DQZAmo/RZa/VPkn8nA3E410B/ECyewXf
ono0iGz1WXpIqpY7LwANJo6HwgvfGpYTnYGa5s5ijsJwB9vTGM8J33ehdQg0u7gLd1fn7l+wV9I1
noaWt0MHuVNmYYfWfQJsmguhskomiW0EVhpL5+7EoOxeFEROH4xstFRYicdt8vHCkpGxc8oHz4MM
TT6FIRgN/QYZCrocXkgqXTJAc3lOtdcNdXyBIDCupMB3ro3jB2k2HXhYz2h/xmm+Au1DvNJNstK6
X/cuQVRBsayFdp0Y4Oni5MQs6JH4iKrmwY//M3+Y7IlqcWSvHo/NubFujSNnkZLSB2CggkazbOfY
MwS+nqZb4njbGPXKpc8EpY2O+NGo54qe3HUyaoov5nRmlouriPAlYvLZPGdIq/4wOQgqygeWpWWm
4SN+vQ7JN47/6ZcObD36dLVhIlHKTfuAyZ99YXJoXz9sdYH4SqLrTo1dEKIGC8RRyyZyYXXpwgHV
YoSMPWMoq4GDNPk69SYbFe4ue0ezZSk84f2Jn1oDD9hST4s7VfuIRFJuTFcX5V8T7YtH4Yxes8pj
ORycOZlwQqxA7DgK48jkkCU0xGslq8w8ha08Z40q4+T3gvY/Zy4m8OJ9NfSzFAvM3/4KiieZuyFS
YfSmXcyJ+YQKkCVtLmWyxuTPH1C+jWpavhlAXOdQ79edxLUvVkfJa2AvSUCffNHkuuXmVtnMDeYR
ZV4N1+8o9ODTZ+auhYwqITZbXT0P67qS44PeKF5z2UXpL7o3nXUQBeLiz+KflMYu1yJd530Vyosk
DTyP79l6fZ3ajgoFtWHUpAMzvRtionRfgPGkzmDyFbsQ6Xxdb5YNdtcOC9Ce20Q2LN6CLJ9iNwwW
YyPJuqMFFMs8CqGECDXH4oH8NLmk3f2x9oL1HVISbJL+cFjquT0qUV0TrODhYV5qhiWc7ASoARl5
12lp+JKFBQDJ3pfgOG9A7Q/7IAyRq0SK3y2EqU7I10AZlNS6lRLVGQKjiNGDPslAQNGnZzOC12H4
+6S6z6naZGpoUoik/GDxoqaFOpYeSTpURGoOqwSJxPl52Kah97Yb5EesMlQNxaAv96gm7aJTb4Ga
1PDfdGyYnyjVJJKk8A8M+78TQ2lHkjLVOPzGUgKmbbyf1t68vLME+vu9zp/d4DO8M/9hIBPDKM4z
/L8k4vSG0V8IjSOkTVJdyelRjc8v3mqNjNPusWohx9mQiYPGlKtl+2ZZ6Oz4PP/hiK7ihFY2KHu5
/I9iX60DG/AC9kpE6DgiwMU/uCoVlqnu70sRFaUDiDMIXRhnScm1lCGGJ1E0OshZlQfyEysU/J2v
N3fncsUz6gwROIdCqmM8sp7omWeh3MZ6TDryFpvnjDyXstDME2bnaHfsnGTA+aNUu+VIWJ0PVQYZ
62ZQJNO/LspcwNg3PuHwRwbIEKWIEpOyU6l49gZJqov2iyU5F0ZuJnvfjMspYUEun4zWXgZZGLK4
c2SfGzmEFRkpkn0lxG9EXHodMS57NFyLbnyzc3lQjUcLeeuztO/YSI1A4d4s1W6Wvb2dOruby2gy
gT8hsx8OUszucXC7n47MqXbL+//mfTT4Q9itYSwnSw7cA/olAA40zD1L6vS6GgUJrm/St9aZrltN
ImQ8bLMqq1wXcH2LA51zNoFaOocFGKascv/avs/EKX4FDU5zMHb3C1oju7Qj+6skqaV0zCJHpvVD
Km3YofFTIBdaekq0nbrVWQVbhtc9k6PByGVJsCYKzqCOsNNBLckf6NIL5o+8+clLXt+FXLow8cJ0
pAEcdwgS+PX7v10ZtY4Ic+DPjYQez+mmqUKaWCryHtQDbRPSFeI/DdLN4PiWrTDBUlh4nb9PAN1h
WtaMe886lBjG5fHX5BlnLHIQfTofhi1LRoMkcPU8wo3kgsFAC2gyMe9Xv6FmvIKekURSOc9KWdyL
D3Dd5S1GRg7ni2p6B5aDHudVLdUZL59yl4NoYY6yG9w4hulEzJrfxTT/L4d8W47siC2lToftnnms
uO4DN274Nhs3yxYlHNy4WqNQ/GSbmmV23y9I34TncOqPtsUc/tQP9I/galj7rZlTiN4gvtLXPdfy
vSyiFc9142UbnpcpG4FANSpMT8wgTGFoCSqt3C3o+eByZgQJYMI96LfWtHTyLCXXK/u3/tJBjPyw
d78bbggf5Va9LyZV7TVyBgjUa4v4kk1d+l/lOhc1nTQXf3M0TdCENpqjzqGTIYdgvWuXfipn2C3v
N630dLCVUjsWzpJaKCVTMwirnYa6fV0NfR6ZEfSbJX1rnohynE6COfcVn8dypC3Woj0Zp2HZlyPK
g4ujScY6u+7lMCGRau5WzkyNLqSX6cFUhrnH0vx4V+j12GjRgpSJgYbzEDO+JGESFnn7zfICiQO1
FftDoKLg8fJTYC0YZP8YinuA7th0Rdhxne086Il+uZQ50F4fo9DHViuuE1B5nZ6GZPQITOjKmgkq
7OBKbqg2X1/esTVkBSBWKeo5/p50zzjRybC95CwoOun35gdHarEbgGHk7sC0nosPT8Pg+aYotKLZ
p+s8De9zeTzViOp+bDJyQ33swrc9/8eTpJHw7CeurA4jy/uO7j9CUR8pXJuyY2BdNDR8rU8jBSSW
guj5uAfp8OHYXAJZEBogG/4opPbCjTEPgtnslAbNszYjTyu9q8LJC3XzqJXYG+D722tTzlQrOhy7
g9cZJR1kp3W84yyM10mx0C5yJNFfATolX1bgvfa84uOD3KKa/TAL9+mQkCuz0Mu9nzjeRVqoR725
9mlKcWW+v1oHhlTJp1lhHRCiKKHLBaGeyCD0jqQv6L5+IwtJ/rB2GoUJnWBICvqTZxGB6z6ey9gO
cjoCGEqUC+sSZP9MxNFFdcXGCGmCZyzyVzcSARYPjPWK4r6lgzMKMj4BXC+D+rV+t3z0S9wAIzWV
IJzycYMPpYvnTZR2RUvGs90N8s8V1Am8h6uzI8IvNFc+LOOQF74sjSZ/Nc5dZvJUKci2bg+l38ON
+xP3dih4qz0mq3yLog4jJQeO19ci6nR2fH+Kv0Iav3OfT8uLivxc5Sb75ZGw2fYIAnOVs13TqtUA
O4owG9LxgUI6byMpn3Mkfbf63gFiBEpdiPaOpSol+Jq6excZB54ljJs35tAsWZk+pGj0Nhewm2QZ
KAXPGhyZvd7L2SYZs/wDbuP3/msXLesLTxz2Lmyf59hexVgE2YZz4hS54f9plLVlUjicE31K7WYc
PH7BEEfG0t7EMxSA3sAMe2ApTPLyGKvXc6wuJOhQ9KbpPdhuB4OA8WeA/xIIX3A0meHM5sSWSc7d
UMYngH87QmsDlgaT+QXsnVyQM9ODR4MrukiFVDmD6M1p+jxFKbmAC+B8pB6HBl0J0Cund6yOo+fM
WUEfETvrF5OYyaKQ5Tk4MYB4Fv0Yb0k8uWIH6YR/0M7Nni4GaawZW7ycZZhT910Mu0Ik6ysxcp3b
IrrAVXw6Khi3I8Pl3kX48bP1Dn4Ve4bphgIA7iSnspBvTULMYxY2eUx+32Y6vznrFWc/YlURz8+E
FK0cmzvJ7ZsJkuD8GMltY/qID/vVMB9OgKNYz/KsRRO8XGarpIlfUY+9rz9w1NrKV9mwi54TkPiQ
bSG7dujGvWKL4fZ18wzLOuD5dFeKvXRpvDTcie2948Tj0fz25LXNMM4MXPFC68ylJeiaEuLDUP3w
YU5/jtvXe/klOpL7cFT8ptJXgF8S0cVMw3YnlvDJS+QMhcYpgYQhz0HfoO1aToEc9fzWqThXDPki
ZcpoU6jAJEkX+nq8XPlUyCOk6BrR0ex3gZVFWr+uEjWNjZIYa3yj0nm5gRD+jgkifO78Fg+wHlUC
FL4kyAdrKDriL79s5ptxNS5tx9y2e3ZN9Am0XV7zHSkb+VDsR6otrqz3wW92HYGfvU4ld+wRiYcc
hlF+rKkIq2s5BR7woJ1rKVmNX1VLDL73c2dN5fA/DO1NUE9XzLcNcx+l0xw+LfhGcGOXCqaBKSOo
Tvi+9xsYt8PPm/rps1LZjwa0EISu01kaHSZ2UNOZTr5zk5Lm2ambgtGWQA6mjAxw1BIMAiSlmXxj
UsQsds90AWJG1ewmzuXvmUuSNBVrvX7BNMD7eeaiyTOpCsGlVhSYnABduIm2z2DaSvX1WguPXoTG
e2lrh6UTQe5OAFnUoeoVfpdyVUkvhF7CQCvLKoSV7l+lbaIGjLmUsathn4shiktRQKN1NPZfE5Si
UjcWfSQY1fP8B/0Lo3BzAo/90pbIuPAGk0ePJ35v1pazA26JsHYRlocH+Dcua20S6j+dtl3StJGT
9v3KajrfPNSc19Aqk1wz9usHPWiCQb58lHMHoTGKurWqlF8ZapZnYcR/3kKfdo/42WJ42VId1EsA
UnTj8/lnxgSU6vcBJRdWiPPBGIXurAa1eWaU1uDTwqtwlmlse9Nhu0hmE7D2UHKED7PcWOPBdBx3
7Ta3asolOU2u8PjWX0B0nO9vbshrkmBCCwpo2CgLi2+zG1+dS/8/qSXNhrES1hwzs+oIq0O2yNls
NduHX/ACCbd8vNz4dXisiuNhFCqdhKGGFpJL5cLiX/hKoLbssF6WwZvtpagoRj/WP6tfD5SzbS3M
JJqTLYRJSYT8NaV8/3MMJLEHNvyJXwrKVlmtyckyoZeY2nZsKgaM7nG8YdtohA/EKzAUR2Clyt2b
o7hNESyL2wxruqK35pn/6IbaHLaqhp+MdmqiouFSImdvuiQwUZslrCMsmyqqh0KqUkUH28Yk7bO1
MuEJtYvIUSKuN4xTwE/IzVkQmZxgUACgSGPLGU8xwT7zMuf2NSpC1PL/N9a1j8/rLDaqpwiWeKso
jKGrsK+SN/iyWRz/JsJHa1rbJkgFh8b/Cz+2d/buXcXsNiYByoRDSijywfY8iH6XXmhUoqXusTGA
LomEm5CGjcyTBkrc0hHYCOXe4kBqHQFir58bkDtkqxDTpAxXY7xnIfyjmUgVAIYsbsanWUrqeNVy
RuUMWBwNchmSpg8osrvy3ddeibmZrI89OQ2ApVCp9gZ3AU65BMRDBr/rfvsO+1vTRetY6B4uYE+/
oOhS6WX2CbDhHmQF++28QN3z/vq9ify99Rn2BSuvQZDj8oIpgcB4vk+rRXrWKd6mBfGoJKhU/l8A
NcWOa2h11ZeeijENWR6CG4uohXcxv/KCx7YkwvPEYirPZUDJvrsWS7TE/2QW0vgdKCzPeOj8jMZU
Macptmy7c1/QfQRAw3pZR3lhseYlTCA5LXPvIxXheeB04kHKcP33odh1J2gSxriZUlQbelfTV4fR
UOMA10mk9zY6QTGljU1dR2jrk+9+enW2qxKhuoiHbeEuIwU2ty8ClciIud7Be+RFduKVJwX/zo9S
msndayCdFD8JSRGwLakZJxKeSpJr8WQqFnK5bYatemr/g6f9HMFSnmk0eVVO1GDh3NqJBjOB4JdV
vAOYGkyHqJ6yQEQUX6IWTDz8W6MXFMSYAYLdLiWSMiKlkFP61DNsTZJ/bvdd239Wqs0czqhDQM0M
2hdX7W6C7bmu0PVPuebD7JG2nxkoE/uwzKyxQ1meYyo1vZdTc3G+xQ9lLiZ7b5Pvg4qVa/1N2gcF
G/7E0g5rLXaFgHkzyYurv3uXHgtu3mbtRbXL5o3m+LlNz72zkNEHF5n9kUmo3NA8Xq39ECxwZy7L
hK+moW9VA4Ku5logvGXAmPEzhaQEKDs97OPfDiq37Wphe75e7zi4cHdWUELDshAx89jFfvtCLpFB
sr2eptIc0e+xxdEKMeH106b3psp+VvZ4gwi1PlIQplHWQNVUrOdlp/s1+L6l+xCKzs9j/mnZ4486
kU3Kl/nf6/JkM6F+qLSjt1isVRZjCCqrtC7gsdDrjcJnNXWkpDuWH7f/Pwt3gFTn4upfrxJ1Y2sP
PhcYtdNIC46bpWlQq+Vqm9NlSfn1QTftPj8J2qO6JuDA/9aZM2BickWOOlRezwmb10NmMWESgE/1
IK1xzsNDrgA79W8lPmS8RaF9fIWYmBuMxrRaPGi8ndICYd5cPROxZpNzodWAQvds8lBBoczdOxUu
l88nuMr3zt28Px4+IwgfPIml+ZzW4urSd+LJrcyeY6N7pSDOgYvQBLjrBBtyDD9JkuotDCeU1wkI
GqZz3H1diQ2lBHc34WvVw9DGlklNcprXsMbat/Jk3FTa8y2pOU/sJRWxGDHI16NnGVB1GzEFtCi3
uoqTvk4CiiMm73z62R4I3dq5PMmlbOHXtLbVmMUor7kVlXbrP1NIVHlyIPNG1V5FCTte9JxmZnLW
D1F3xxZB+sWyrZCir/l7hN0/FqXWySpfy9KnAkBP9+EKxerUlbt6IolBabcjILUlrPqKBav9aza3
/Rr2fowV8VRzzg4Y5Kvq5qxWWdZWY95nL+PHJe1GGEePmrrwUiaIog6UBiqaFd7yjLYwWwiqZVyD
HwPNawSfpY0xiT3eh7GFKZYbCbgRGgbZPRgoZrVfYh55eYzwCBK1nmHdnwdGTJdz5ZNutRJGPyH9
mRVRU4teg/NBGns44odyTrmN6faPCqzf+N4ZEWLzb2IrkenMZuV8TL9zr60xMM1uVWlus7MJE7yV
yB7NmwAzhqrUrAGw2QPpg3OTlMvXoIBcY9Be75vmjZbkGoojyegvYlK6v0Zsld9YCcZ7uHTbhbpf
POzcAM6dv7HNhU/0+T51A3QJ+wGWxqY09eg+D3D/SigLhfldM23kEwQfR3UEyQs2iNyR8YlkQxTS
oHQGyU4QmMw9CysbFuJ+ydyzu4UABYtqsVHyg4s6wX69yOAJmJ1jMbQthr+WDXSuIRT6lc+Xm7uZ
jJ4pCtxxQtgF3cWMzCdH/fFV6BD+Jz0eVpo9n/nCZt9cc3ronod7dEPRGF9QDZ1X12jK477cI4p7
FiGRiH3jvHOJsfgEzgO34vBNDtBL8Vx+vh7z/+kgkjSPZxQMZF4P68eKVwpjvTbKZtilm91FIPfA
yvht/zt786+pWfGZNQf0Aw/qpmkrffooRpYFM2H0cmXC5jlzGLwaUpacJ2VkbRPvcC041tfzTJ37
V8g64NApXudf3bS5cEq0nFmbZHfRZVpzX5mifQQbitjV6euvY65wjgKb607L6MeOt/zxjvdlYyV1
GtSNDMaaHkfLsa1qFftuqPKhT9nMUXtf/0IjW1pVx8u57gFZlYbJwTrFk4z7n60mdg+0IZwQlV19
Udx0nkihlRnfvIpWHRVnbjfhFN4xIlec4uugV8WdyJ4z15CJj/+2jX2wDmdvntnF0i78Hmxs5WAl
9vEdDbRQq3G1zA0GfF/WnhmjvaKzm5lZewJdBviG5iR4wrIzuQqZWXyq9+KgKtRH3XcesIBoR1Aq
CGgCX5foIMtkiV0eafiXweMpBKgRLTqazyjhwZe3WQ7XDqf3cehi9aLjYsyf23hibd6ZzlmUMMaq
9X9dVHx32+4Ya0f+I7Q9lE1XnAtyF4Qaec4jnmPon4ztpLa9rd/+XDKhNZ7Vn+masYfgd9Odf2Le
BIa0wsUnMVfZMBhk3fCDb1yDXj5ozwCWDshg7BlbaS/rOnMtbI3Uh/GXH9UJVh6AFT23O/Tofaf1
41H15DN5/Q/u3zZKziaK7qYaz2kNOI86ot95CpGMR81MP0ULHzcNwgFzL3tYEh+XLaef5ldOvXkK
aTd9tYoBCet8jYghV14myBEk4JnI8VpKBF5S62c/amDkOQrT0FvJft0xlIi+5M3iSUbYDLQQkRvX
yGcI0nmLwTT1FNBTNK/mJD1kpdW3CuDX8c9XzCtNkOebopadLyVULieNtY4Qb/jGVdBe4CyadVNt
CpwjPgB5HcI0sjI60VnevZp2Q6liziBdZl1hdyG4gN5S2KMYbFnjlipYeByn/qR6ueePCtRNEhGc
rDqcEGq7ytBFbj/+0D6P4DoYBIip79CDx0E1qVVYCbv3f26vlk8SxwE7EmIUqE2xbc3rihiaDLE0
zPqqV8pTgbhBeoVrRl8LxJsF5vRgNACu3pKfDfLtjbgLQFexZTvEHeIjCB6GYay+lNGic5QeJols
UIj5PlD4QqcIzpp4zQax0PMjRZf9Gl5bO9sHCLVi2bOhpyWHSq4gCm07b9TFZsIuEOgwgGAWGvtN
PweMfl74ESyqPq4+iBqdugb19EKo4C4rVtHOSE7cgNFJPPFFDbodWC/+MEG1qVePtDarN417UJrB
ttC/Fm+Q0nuLsjNnvWj8bLBNZGRJSwEQjoWPDYyg6wAB3FBBqrQZAxOScs9KTEb3rFo0WKjxd7Dq
Vy6J6kEjOSdYGBXtgoEX2CQcAiwBkbpC4JTzbB/VQOmNpP0L/mpMYvVwJfrlOmFiUphY2+Ns8tfO
1+I2sgwEQ7NDiJADogj+goQUhpkCt3YsKkDx1hEiUQuuFtkczi8vSG9Jvrb/5TxkF3wCsp6zchTq
Z2YWDY2+xHZyHOmFLwFyIGAM5W68IjSzrnWiyPrXTPjkUEpAel7BnJ0H2hTKnjKiZnvzaoeHaYyu
fFm85muPckJIY8hU4+meAIPTtR1WaWt8En2QYvNQp2sU68K+ZIkTuxsl9Ti1WRfz1brTy1YvRuNH
LzG1AVoGFXWX4YGBDx46IgJaxaF/dAXO58bwVjAn/I/bSSRZJJ4hFW3wFEF0LSWY3FXL7u35rZ2b
zDlqXEKr4j3iSndAI8q579zXF8uhFl9LK7whiSpBIgF7l4VVVzSJzmm1f6K17ChspVg7eF7Sxwme
DWAYtRi0suHVyZpmyS0EOb8YyoLEZX9Dpb3xGYXXyroCe1OExJ5lw+/C7UKccdJRrcS5dSVLyJT7
VRHNjV6ENeGi9TkGO6lZIIHW3oX7GvGzIqSCt+0+/7TnjTsgw9N5r485ZKGzYDY0kZU+NdBSlMSv
+PtcCV/TzhkeKetVqnRUGCxi8na/CFSvQwLpAeiUSRMAsQ+oKkssvgxT2asMDYCrkyuLkFqN/u6x
d2ZiPrJJDaIYNLGTrWZtM5ygrp+8pKtXBl8euEeF48SF5RhOzP3uodSaumJGVDH6JvdwY75J8irT
NVVosh3cE46cpws/d91J+qhD/DiXUrSUx3vL2iZbhTVDCvJrT5UyUj4RqM0mVfm1GFrBUJZkeoo/
1WvX65yfO0lNgx+NyZK4xN6EerYP1L6qVdfy4RSx3mUpciZ+ikK7iF74VRfmtu/MeDyb2MoEsObk
UjZq3E+QJduQxjOxwAecqxbBd3QoQy6p56jieuvaKqLBrzdnhuAAzYRVr/eWoKoSvPqDW4IJ6fv8
4zAjAMoQfV+kuYzv+rXwIq3b+3lzLiIKoYkPQJ8M4nZURtJNTFeHwGj9efdNyludmVx/px8gI08q
qig0N5Oh8kVigYJ9NmI3Ej3TFRmXLIlgjEapOqBB6c5IpiEEUhLHkhvKGqrRS7LIcC2RxkTUltAZ
gpmEQTNYHviS49NBs/PZR68KT+5eXvnbuyS3OuTeshKAORs5djbH0r5Wht2iw2RyW8DZf2Fnn3k6
oF2OLCIvCyVp9HtayCx7NYDoKw1AGY6Y17ReFyLUSG54Ek/HoGeL0mmRdqGhPslpywf18CjlSpnJ
zpcTfRaIPL2QhVk4BQb4MkXcR4LydMPSRuUX1a9JkjKTA8sdCa8LhVAbx+uUnqMRJZNYZuopykCY
z269yQt3J5St5L1FPCUWNSXSV0yb7N86L1PAk+DLpypWZypdgHmn5JCdjYT3k4vJBt6v6K487WqC
D5szEXkU1wALt/JnISxTcNrJkbX+6r/dfiYi27o2bRbaI2gpKkaM6EYF3W78IHwPdXPgFb2PIQZN
y5L2TMBy2SrMLpghMuaZ2StdZKYo4BCL+LeP4jMCgHJ0SYzoZIwQ8fwqNphUJHcO+CPRIL1SL8H9
JCfNiod9PaKt1wu7ys+ixmFBHtTaMKyqov/qpMoG3vRMQ+CG+6Jq+bYoMgpXqK4jAyFgcWhZtkuj
zPnVFIOyJEoCQmufIGDgIG3sG5jMctUaMhvETN4mr3w8GU1Nt6mW9Cbo7NjV9h0OHlGSsOL+7YHY
NTnHojzYMIpeePfhSt7eyVn/v3GbNO3lTV/s49PGvdNHXHQkd+AWsaNA+wD1kc+kDBHaovwNohPr
kKfRGRVr+7OFEQoBmR1yCP3bwFpGuPVqpJnvxkZ4NJGA8wmdg++U987b5mh7KjPa4p/yYO/lqF/C
BNQiCWuxJxciPwjTCl47zq1H9FkjY9ZZ/JxhD1/SOT0cWWXv2rr8emWCYINt34u+deVoB8ToU3GD
0Sm8pGJZuW4ARba62GqeNe1lhWgb1qVfDbTA2DmFOxo1rNKNldCcUao9ise7s2/Td8kYBlp0pHgx
YQSpU/G5Vgs9dZhqOfQyV8U3ZoIrpzd7T1dSAgvbPrdzJUWWqRFqnNKQ7QbAE7XPWaKh7X2aZu4q
bgeTsF2ab0ZXpML/no5DdEAYJTf1gEyb+OwlSqmVoyd+oon0cyys1LJum3toWs19EC2Cq4+ujMoW
fP6JRMtdfognYTZhBFiSqDHy7xAaAXCVzwPYQRFitBL7Wgs20eGbrWdJPD36YzTF6C3NHc/gcJZ6
q/20gC5f1H6QC8tkHMjwRD/yFjOTLPbHuSfZRIOnkRzG9He63gri/fBUgF40PJSJuX3tyBbwPYZO
PJ9b3i0n3UL0aQOVBCz1JdXcT8o1q8qLtbiFx0yNQXPz7k5HKDcLhz5CH7NZgU4LHkHVQvR4b5so
nZls02VRPv0trSavj2XzvDVe7X/LaNdr5eQRf+CKwydgd7lR0wN7sHhqLH1vR02XPTbIt1PG2Pdt
Zd8JGl8nxUV4PhG5EdY9q82mzTCV+x0b5LRzZSJngoGmslYXF7isKVRDQXKukp9/Pj0CgCr7f6/w
unXyOS6IYMNEtxBJRSmdAQSGJrH68DGApJBG7LviWBAPqRRMIyPnJjGUzcJC8JzWrexNM4TzdBpD
xKRFjg5EGi/Kpfzg/W/wB+3Y3ZoH7IXU9jDgg+NZYSVrt/5VQxzBHZG4tEbpMp2Ee10aLTwCYjRF
FJWcKjyUhvDx7r5RcQUkbSIOYRLWs+gG5nS7KMuXBgeeL3u7AcHkYxsCtHPL/3UnriBh30qN35Rg
L9aMwUS5FtAQGEDeCbfeZsYRX6d6zzejolcO7vKMQwx7sZ0IGk4Y/obedAnDPP2qZWPziQFvqnod
2YNXUPhqjkLnQQlyupxcSXIbRVSuTs4o3RcF
`protect end_protected

