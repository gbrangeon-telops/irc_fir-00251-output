

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ISK+8BrzqbDVc2hIh4k9UuGvqsq6yFic71tfszsK7KRf52jFUoK33AosGVUYsGH1pmrUc2NUQcDQ
LseNrcojiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CxxZHetyKRTjg1ePIJzq+w/Yg+inN7g9nkhYUjpPSXav+SKIAQvdh174FZUi0SnoR2INo+rdZ3gz
yq46XymO3b/3npnRNCCU259giTvnOJxmkrtnjRyUpOg8jB2jnHg/f/BlL3OJUGGiFonBs+6rnNvW
4aiU6ycFpLQsNzqRlAw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HZ1Kttz7DNn3t428AVZ/hrbCqljpJfsdfcEo7T7pfqxl88ELioDFFp9rVcvvZiZMU++45qS8CpOD
SfwcEjOj8ndwnIsrDamIUHs+Qm4vUDDq8EtyiGhux+pwMtpg8rH6kCwLDCkdk848fWRbBOGctdAr
AiQz4Fie2ectzKGEhjERjquMNqkQkhNIuEu/CSTnyD7KnG+FK+llVBavN8lxjWeDvk+quMyk8Dbo
gA/SdzYI7TCZkNEFS/PvF3Z8fPBK4pBWz7TyfdHacMjMkaPd5zGsPBmQy77xwc4m/sfhM7ZX+YW6
VBTILiYtg7u194UVgu4fHE7f45jr0jTur9wbVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2VX2NPBJC/FYSjnVp8ueqtxuxLgenRIKbrff8tdhuTb77js7o9S4OVH2n84fEyvr3hl3lrO9ekVq
VvQQOlQBg7Zv5/tFAeI5YFisgygYrqeX9dQcI485CaCpeN9nanYXhtHWROH+ZOYckBZHUhhjC82p
LnYwoausKSjsi+rXE64=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HdQIwrCqCFDZv9OQZsva3DMtF+8TwiePvWLQndNAXK/1V46C6C4sVLdH6SK4FvPis45PZ52T91rx
x7mjaMnTgTVkK+VoFF3Ej7xzh/2PoR+YkiToyHCbvwHQXXvv3GAu3HyqWx9b4oOndnrx5Z1mco/s
lNgEY825qOfDqrTkPvvNBXThybVoOKs2SBHAdaQhQemuYVAjS7mEC/lA7vom+55/0dhIN44Q0vMz
6utkLeK9axPmrUz/LHNLm3BFQsfvacsQoIQe/Y7g5V8ehxANfnzft/Jgo74fJAU3odGS++0PsHF5
2T1joNptoFFljB/U6DScrAB2FxigoQal7I/OSA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4112)
`protect data_block
w51AxCtstcayS6nuUSL77n2rUzrLCfQyZltKSlIjCfLErZvx70Ya3ZOAEr1EIFe+oOqhRFY0cm4i
0Ze88F1EwgFq21CgzYsq7cu1LbH+7kIptOHVOsyXYZNu3J78j2cPMUsXIJAGRvPnBxL+R5zBiOnL
AUydGiOieMC54jAD/J/XmYDwrc+cLntayDs6eksz9tE4ffkTLvGn/8LQGF12wKqC5QOT7FrC4cfT
m9oQPfXG8aPYXE1uR9hq+bVsD3oTTMJHEfeq3qib7XkmdKgldMjRmvAbuTFww+P2VMf4vIueouP9
xFASo+ZszRmxSO9PFwNnOYVKTn115awINQU1FkmroDhT+spD9AWM0VBtgsPpYuL4X2d79CD/nfNQ
8CiWxEEXYB6vDSDZN89fmKK02ceKjdVf694/brYE0QsMPo4kIKdV0KgJceW177KGoj3C3pl5vRcK
+uvYNB3QWUM/hMjNUcNB6p1nK8Wujx3F3f9bVml6akPpTeBjQ7YpKRhs+75Y+QfKEOjMVlvsnij+
rFTgy6HiL6HU7nXvnD362BBkJPsl/bwv4ETFdDOG9IuG+Uo9gWBacVk9bxGLDrbMqTk7FW5FhgIi
5yT2B0h+eaclLiVlM2gheOCPU7u1NMUA/irLFLK837l/IhLvbmEyiE2BDaSxzyY4KlWklvBlEGAo
ivcwWcs/6l2kY/6uFEu/zMk5eLXadhhB9OYAz2NpnzidMWpmWP3YxKELEx+nO5+mz9tqlJIpXQeg
Y0DmA8zGFiQBEiesEaxNpo5Dqv3nxd6Uw4qdhD8yPFz9BON06qFnjlF52p2hCp0Px1Y/uMemnJv1
Or9v9Mu/jcA2+l1Q/6jBmiy7xfOU5+6a0a+hC3BzJh+1VTVmb3mY+CAUT8vaoVlNqEvUSQrzRVrE
zSwttC0kik2xrrDkuzCp6Up9Q92KG/FWbTTMrmKzTJ2BRA4hwskfOYTfPvBLiGLaG3LJL8i3Jm8B
DlHj2iglq13lZYQ++mwldaInAY12GtPZ4airrAEvpZ08q2o2sXbPziYvoRzSo4OOsMQYUb8OahlO
QNgVzvXRuKqDxSvvDPIpeOpUAqXzNbTZDoGit9zLnd9GyMYqjApAA2tDz5NnfxTl6vLZcdiTclju
3pWw3m9bNYxKPVWHE1nfMOoIC6i+Ao2a5NRsCeLudd8ezH3DiT+1G4XI8EvJiyjXVnrwAmXcKPcK
3cKkg+BRg4S+6O5BesV50sZzDPCNvbC4iX5qSRQPw82sdswz/FGb5IweDHbMnuQSonY76ajupz1+
So/gpXLMdN5zevmU3dbRecWpIQuTKU8wEcE3J5HdXl63rk88XqRgsNMRwVgKw9x2R9gA+ac9UOsL
ERKmphQL8fs5m0QRoFF3K86oFFIaqG1XxFm63udjnlQhXadikCbpQgGPJqxCB8fqIz4bUu4FVkTe
7kvdJ4AyrnM2tycIlQFqx6Y2JVw7BNpHcHBNBVcnxpr/J2gbT8zXcizPiYXIiVp3pzyyRWKHPeez
51AvBuZVo3wBZJvnu2hcWi0yZ2FbF4mZ4zOmz5i1qJ8K0xRRD2m9UD++8PfbfTX7HDvzuUNcCjdL
1abrIYf1ZJQyXblIdZDiCGksNnM5hvzD2i9S7c7i3rI9+gtvp6COT1RqKNq6eDW1tW7VZngeqsZT
fhJHhrOJrVGvA7xxeve66KdwDb440LIHdXjn6tKU0Z3D/WMdNagEjKR3GhUlBz0ICd5eKELPhcEK
tsXXtTvb433OZNW/riVXqU3OaHwS84h40BO61nzBAWOw8H7dltZodOJIxk1JtLabwFys/iwwJbnQ
1txEkK2B3nWr5z4D/FjDD+n4sijeqZOo0oM335uJ1VMSUAPPBjmeQwybOwqy5MEWGORvoP3R9p4F
f8yzGDs3a+0F7oqLK1Gr1e7BR7PF6k7I9ADxEcJyysjvUg+bAQQHt/01ZEIt/+XlV6qkDGSfw5JT
qMI0INkB/oAqgb7AcJ/Pk1J5q1KIZuH+lDJGl6DFCUr/OtYADafap3zY6xsXx226JIVQtTv6q6Tj
EH9/sTeUfvTJuUSzPN9nYg58fJMdRSmgajnEqCIO4puWzRZNvjn5cyLPeRZsmoemYqjXYiGmweN1
J3IFf/S+w/m/hm8Wie/hGRftPAmrwABiAw4eMTDaRDgItsJDfa0rfkm1IdhMWTvJxcS5UoqmMWpm
1341TgPq95WH5/eKJq9HehoprFsW3iQ82AvHkc4ak7kILEd6cb1or3vr+TRcvGAxAGLujCdU4H++
RlXNqmRpQ4Er+PDczq1kHal/Y46aicsOfxKUyqukcFjljYzYj3ySH4rbV5xudX0gIrrluBCKfl3d
YFUIjp9fuueov2nRvxa5QQ+ALwvvimAR4IRq7K48lsPD5N9VV/JAOWv2Ypd10F+Bi8F2MI7spZ+C
UR8oPnjPPa5U3DsQXLR3UHv+uGIcsm8LnK0FITEOqDm116kFKiFmlo0O6Do12ixJeynyYGpIRmdB
TAW2AdDTlV1k3OFk2HUJ8kHH7qai0UXzGGVBATYfcnnzh6UyI0OFCAFXkAAxtNfSurO2d09f/lOx
NCVEos+biWMR7wp2hFAYHSkS7/jpvsRiZ4Z29cVKPAkaF+8ou8B9dFUscPnT7Qngg2ZfMUuvIyEd
vIUB3/uKlG8NyGD3u9pv2QjJ6bpsmkKYZpUKMjPk1TBxuPTb9rPv81rXUjDNTLmpMP9/7ktW+fuM
N84QW5LMwz9Em6SVxhsseZfEKkY6mAR7wUOOCrqWMWUaME7lH9JZQCYHiA9KzrD6GcFYqSUTgGjD
GQ4666Ptoa0zaHBIeQji+Y80PMvAj8D/jbGqrxOUfpUaclelp8Wsp+5TizVhQEhawtVFzV0c5SMu
ncmiXBpl4xi6OMB5DqFoscqFcCFLVd+vS09OBTeBdKm9evIj086x6uFFQzwmEeF4DQBO+4JKrX54
rqcaxbEC7njOAR6OooZ9OjWW4xO2MzISfa3GDVqXhV6ZzjHSV+A1msxz5b499FHrj7Z7jrHA+2Dk
YgZZi65YxfWlXwjOier4j4wZPxOv/VLQWHAxcWfFnHIcZwK8UsbzI9pmiPXrL1p4zM9ZkOxEIvth
Wpd+sWVF1Jke7geGvuRN/RfomtjiH7f76lxCtd3fQf1laSNzpGugT7/gA5m80cFrYP76IuXGT+7q
wYYKxMjXHTIbfczDs2+tsZEhbRxWsAka9624SQ3G4/wnJAZ6iKmYnUaGcywBRG8KYu0RJUrVmyls
oZ8FWWiBffMrvZOuHo2SK+VjL2UMJeUb7693PwRXs1/ja5WwPM47TTQixS04YzXp2hw1HJSl3jTF
VfntBnAMWYj2SQ8aKSpzJbv/2kITz9Dv067NzsRR/K41lpwrqgx4fisMs/7sqD+XuR3qYpecWrvL
B8vyw+TG1hWhXMHrfi6+tGEuzPciz1Yku4nFZtqzg+tbBzmw6doJizlcMyhsga8RLywjX7ywMiX7
crBx8/QhA32C4pXKM/pqzrfgR8m0U8vhp+nZECdbnJfu3D/Zx4fmuElGvmXXOm9AtPO+02NMj9Mu
gGDAHbMrY/+rXqbBPJcle/oSRtTuOCkK197AH65VwURUckg2NCJvvrjjkGO/YoUu6ibaXK3xg5kf
v/GSZrpKriGp/GxolY6tc9bh3NNisLWYJj+3PXIilRCwodum7DjQRkPqENPNgCXK3hWFwf5ywIoM
eB5swIjdruCA78e7b3MERyyjspvN8O0qQy8C/9OfES4VEK6N1u1GFhdAlHI4VkjguvU2VOVb/Esk
G3iIWtQnP/f1jcps8dH5A1P3sPTFQZDQp3GMdmJ02MMhle+3YDjEVY3ksEdPP+33eZSqdxC9IFlj
WU3B3l/j8emlWC1zSNrMk6ybviylssnnHvuZ0d11/ysbw9IEeCH4vWvDAaYXb9zkgpn1wVkffO0d
zozAWqEwFRb1Kw4yBAHZnG8GiaxD6fnx9I4+vA7WHw98Ju671D7pPnv2yw1KldxIo8nofirE+MEK
hx7NeRIX+yCz3sOUr6bna31jtrLAqm/bQBTLzoQJP2Py7Pc3WmoTPJTvrdoxRWDUOmIpTedSoQ9h
GQn0C30mdx9fbK75xjh0iQCsgTEBTopSQRgxUu80b/QHPIf8V7x0BTmrOZWfzZiJRLO/TTqOPBbm
gng6A/PfBqisV16iK5EFL7ZllAbraPYKRE6gDFbvc/s1boFGBhRSsedmEGAOKz8FSC+si+kt9UdW
Gr8jgl/8OETqysM2iQ1am9xaBBgs0eK0lMDwVdLRYmZJUAs+7ceHLfnz0RGwBAhdw25K9UwOa+2d
4SqV2vj9fUygPnn79fYqzajs5HElnUKcJuDJDUcnXC/PgGZOFyi1E3bxth7tA3UzcfOgLNEAK012
9pIy9/r9pINQjY0iZlf2RUV/CZUDghKfVCrkO+NuyWEUDcMaVZ2dtn15fV/g1n4I5Bjh6ovSmLi8
ahAOgAC2A1lJrK2IcIG+ok9uxKzx7ReuZzdBzXiacdgPDBzoO2TU0mQCUvoef2UY0/auOd81xe4Q
YT282zJpxPYpAtBB98OsrddXBV6q26YSn+0uVQzWT9mozuXnWg30Ud4L9l15uIrR64SUozwiCl3Y
OMaGOp7JpfgMMasbFuvEq7wsgAH3tLWXSjgOnMjRfWBQRFWrQY9iTV0obsVI3wPAXeCWf2cPHDFs
CHBVb7UkwU8QOm2GAYSgCkSjTzy8eqCcFEf+kf+nGmGC/AJZGb4/WhPBL/K48Dy75vDTcHkaX1L/
25MsI+Pv0BJEaRzRwDFwT8Az6VGaci57iE9IcKYS702WKLuD6zhv7wxDlC+X/sy3PWeWxOwqSJfD
ItCk5WSt3IEmIYXx5M/DE9yECnaYLLLpOK1YFZGzh+QuTqR81LvJ5Z5WchTi/4o/tali53Gk2/uD
6xanUlmMpM6sfn4FLAeIzIeuxt0KtM2yp4GBiSRer1L8ZxHZRnBf2oH/JifE5FQXPFvQEfy5YHZ2
xvi2H6g81FkIbcqat9IX0xeZeX/8wLCJFR/RrPz0v7H4pzZl86rx7ctgQdUOvBGJlcfPvEAqUmW7
PcY3qc0PzYBaR+q71ze+R4wU+rk9YVMvkx7ZrwG153DM2DfyqyAsNKNhTjhLxUF1xG9lCddC0zlY
DgG+9Lo/zCGnkW5abCLFgipOBtuZbUbj43KyYBMVUp4ucKEU25c0l++WpUrOjvSioQh5DtIUxkaG
2G5IFaab7R56meKA+eBXOvRfzfSn2+C9dYFQYMjh0A61Z6ju0Kw6zNyUFIYOiyoYsFhuX0GvR4hJ
P8cqJP+6ZT9i9LLOQllzo6iA8oM0jficUC3nHTfM5tW1+RQJq4N0i0Ow36VsP07e+yefOL1njsDe
dSqdv6CKM3ywNCSqep4Axu2N1vFGwJ+PTBRdkOA4WQs4gePVPtgHEndoDW+6VUrk2FTBPhZrSRtc
/f5WHuXyPN0=
`protect end_protected

