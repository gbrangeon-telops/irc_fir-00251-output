

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jjl8vAn2UJruW+pwbvMAIo6yT6bQgTl9+ZqbT+VaAP/dcMa9HxI5w52bG1uOMJkKjbI3shaTb5QH
+WA4TEmwBA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jY7USlQiP9PR+LALAEYZsrKak9VnF4tfhT9SQb5jLUPXs+eC5ZbIVQkPjdV+4wzhB7b7ai6shnHa
gEu6kUZZsMTRIotEQn7SVZESTAIMCGAU4lDLU7RT30ySc+gN3y2heOoScYVxVF3kYNcbErB9g4iU
iZLVkq3ZU0fP1VLA30w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W97r968B0QPwlTs1emSg8mtee0qHNpQ+/n5wfXS0R66Akqy90VsNXhnqLJjbnGJNqaGSMTKCRNVS
ox1Z0rkuemlJn0dMgZtmRgHM/NeyMTSbsBwVvTSeFdA56k6PzciIIQ1S8150Bxbexnd+b7l/UMK+
JO8+KzzHPEIPqou3srZGn9dog9HSSfTUIqvBgloCeGmDxxwlsFwQ2VsrffuE8mB5Kk9lHG/A3rMw
tbJURgYaS/b69KLL9Kc/urEgbRWHU1HQCQDL4hSKE79WXE68MZJ00kcWMfNfAOR1zytQecSerjXJ
iVVvnEzEtzUejpnuhHCRhS+b62dMTzf5a1Q4Dw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l6IXa1kcvqxcIuqXI9bELoLDvGs5XxFfhbXxOKBitloxuDBS5IYgW7AXksTedGB5rM+6jbAr+PVa
4ykVDtx+9n1RZQ3HKQZNsRywuW0+Fcm/MhmC5isxnEClP56JmzAEyD9l7nmy9JJJI11qQTy86iSs
hkUJMmO3Ph4Kz8ptLn0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gEbAM0PoYz0kTXyuDtZRhRtQJeO0ezbVNuHzWd2Q6Djxe3WZnx453sNsfBBqykQPTu/zHrWi/wfe
VIPTt4c20XjDHHTidMXhf5YGMYpytIjNmzV4g6PhJehJgJTQj+T/bAmaDaXLcqMDTjUNont0w58X
XTjVYtxQgjqcVftNf5PS5GCVpRxSTsKbT4CfmHhBwwsNC5rLtE2tRCpmB6tKw/7xf8VLLD8a23zt
cVvVNX0bw3bWCGFmWZjC/1fhYI19WFrjQO9Y/0zq8T/b6JCoxXV2HE4Z2dJ8uXvV5GV8EStC7VCB
DhBS/R4IfNLPojIIJPxvrbzkKlmuEkhgwflRRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57936)
`protect data_block
Qm8D0kNVRwquphi5zPAumh/eB9rzYWb0qPrXfTnYrnv3FwAedL5zPVhx/xsg7jz5u/yjLiGmSD4e
/0N/I2IzKQPDN7bk/De+4v2speGzWGwhYb5CuBPxmK9XTGnYfv/bm5/Dq9Qmlt1RrT5uk3oleJ4k
AFcArMiTdG2H15HM7TggQFqGfuSmf0fmEYRy3IghMoGXWveEidcS6RPaowdHzkhXMD697isNKcxK
c3ZQh4Byi2lkQ8mVjJjbbcVXR7KXc/JDcJBpQ9NgJyOcSmhyWSNH/2EALfYdo1DRIMbjozi4m//0
acaKW2qQJsbcZOUb0eeNKyvLBXfawS08QUkMNAM3XOUIQgxWI/ccW0v54mXRKGpcsXEPSSmoBjRc
99v3GD+fnUAJciCithf66ev8bUjtoOylt80KSKFjM+XBk6ncIeRTeU3qLlqaU392XDDnfUZbdBl6
5t2OaxyBqHKzM3zNR7zrG3g6eJAus6XfqDXCaRhNcTrDRX2IJwja45VnrDDN2MMq7vcs0QovrKFJ
5iV5nzx1g0L9R0Z7hqs4U7Hd/dkNJRS1SWBspKFV2hQLsURH3dmUl5+mLvflTP4viYvWvZx6IIda
4QwH1RuvJ3pC2NR+CCH0Pi0HcSsWQu/VwbXWb08KH2jJgRDZnspUJpzhSeGD8A1lhYE85E8s0izI
PcGBbI+tJiqyWdD3FsRwwLiCkAwORyjAZPJJQCPL9VI0lXS4sDFg1uQ3Y9h7lGkGvI1FrGwjF0L1
NvvMXzi2NWEyQywCXiPGx0iNjZrX9wEVzPIujMg6cfyFKEHbbBkZje9Nmg+Qec+YH3tZJ9+G8koo
179DQp+KwNdp5QUa4OnSiq6w8X1Sa+CD4gywu5UF07SsGBx15MHHAsOXBm1nBWjVkncTyqgsdd2w
74MRtBAK4SPv1rPL0pkoZ/qa3vuVku700d/A/X94HAbFM265ZuixHQpQJJfU8r4RM4p9Bp7MdlBy
hTMdGKDPiRNsLnyGWQhDHPiYMzdwr5QXNcDcFqCV1fvF2/d2+CwJYaMvwNG7tDUfviu9pCBkKRSV
t0eHKebalPjcJgTnL1eZZNFN8OyGbFCmqzudpFSnj/kbV0TETO553gVXhJ1/6Y2CSZNA3yBt9X0b
s6ieogCo+7QEMYF/cUeienHl3eIPJguOuBfD5F8fKYRUxtNqNrEMvP2PuEjEZdu+GYU3reINdEU4
nISMpGqDvewaJ16dupS/fLzI0AbS6V9WHz4y51HclTA1jwPs5iuN+53Rwobq8gtxfodfzdbZP+8o
xB11GvNRaMtMAOSSVRMgSDj8zrzOeHIIQoXJMTJAQS07aIeeSO2RGr9fOFiTWilpxkh0S7CjYOcV
RuqEhqs+ysuxA7jpurw9iAFCJB7tCPrNX5A03JojeJXEGalbIc/cqvIFuNfoZ2LUUaP6rLyIu0Gc
R+s+o0qdMwyakmPZqrXCR9M7SjWltdcIq7XmM8HfJ0b2tRrhuGZAToklTQDiUUZGAP/WgKzwnLXJ
4qbiAnxtxbHcAVea3sAFlphfnjSIUAK00bFjKi3EgGWsY0C2b6rjpteTzCzIoTFwbhYRoRu5JpLq
VIrLFLjTjAhmSCg+iavS1kkDNdteHsMFzWfin2wUWDMAAc2RRqCkltb0VUiFxXQTFXZi5tZQe15C
c9q2V2MFCMMor5hyYTBhmVhM7kXmToKKTkaWYdadtWuOrP6BSjQdeSGi6f2NHoalUyuER51QeRCB
Tjo/gQqeys0ofuxrR24JM6xXplnb7uAnUOrNsRu6rMlwia9vi7pAvi1s3a6kjj6ij9EIbTqznl5I
xMiBESs1pKEExHPSJlmgAFMAWFjX3hToZ81ebNLm3eaeTVDKiRDHw9WOhbG+yQkDo1p+BZ5zbT1T
gGZkmkJhXi7wthSk9307DBiCufK1hJap1EJx82PtliGg9T99VRmt0bMt6rAjjVhyO8UgWvhdq7cy
udmVZwlVTc/RiDPFrgCzRnEFhV7jgsxb3JWBWbG2aZM4Emjoo4SVDFo0QfxDonUlFHXtG+nwAKgt
JekOJYgFV4HosWxN1jU2xsMvVKugQM4aGLzA7nlfM4IKlo8eMlTxHmcjI2Pt6jdAYrntSFRYWacr
GiCHCxRc0981UO+8PsJbnPSZlsKT7gRWEabvUzFd+FLP3qywi7eK8EG7oDAMlk/FLRybn1vRZwb2
SO+X/HgO9TJ4UmbH1ihCDCSNvnYhxKK2ey5PeuhdMaS+ENk6w31BVVdDkx+LIkuPv5g9xkY0sS7n
WC9kgqrCccoXjUVZRTlty/b+/4pKzlVkt72htP4zQopuWu6rYtLSLfiRqdnL42lesZTyXoDpzTtv
b7ttJA9Ime04W2XdAzYLMh2Rc65E7dTmr+v1dsmszj8wXLD/qE/ykYKWaMWc1KGin9DyGBrmMLWe
gKnL/WuTPuSoUV6UiP+amat3gz3KKjDSjOKKu5gOvTI6mCBCfzH+phOsQ3OPd3blre9qG3uBeEn9
acMBAj1yMKg3LS1WGDUU2ZvpG4AdwxQw6B2RI28xG70zv3RuxDOJVQAs6YkG2Ii28iC7oKJBlwxZ
fvFNJS3b6dRAzC3fU470VbIALQOg795gzod4rI87cBEr+ICJASDy/JbXv3tV7kXvw5LqvSNm+Vf8
hOcxtIiIvZm0H80TpxrW2eYiax91cRQMzAFWaNnBLEZrjfi9wAl1D3S2X592WwjKq60qGIBu+SXD
TzEz3KIfx7/VrRr8As+zQY75ZQl4l7R6Fi8gbivkwbm/lNM/j3rO4VS26Y6t9Qoe8h2yutXVi5uF
9Oppj+dZEFxp/dtDi3KCaAmmECz2zy8xcS5HrSSWLbUv6zuikHhrcgCNHjY4kHV8LCdblffi613z
dfjIBrG0R6pUsGMBjvpifi6l6PCU6kh/J2Ke8mcW3VJ6EWtAvnJQxbwt1eVkun+K9IMNbqE31tSf
/yWln5kw0W1ksJV/OfI7Bf5KILR0CDH1edhnAONLN25Rak2OME/W2I9Ve/VyhsuqPxWWXm5ZWMge
k2/X8+DP5u4ZH3UsPKaFRY6VJBespLbh1Uvyw3B20+lWMJhyIXOW94mWHazLLll+FcXxN8VzZUFY
x2kt04fsnHK35ndSHHwvjAf0ibwgMXerLOsTTY5es5fLwyj2dx6yaYPrZcpHCt72pENJlUoUyLVA
PG1LjlT3CBqH2WFHsf3ECbmxcOQ6M5hg49IdAG9pzDs2Sb2palmXl2b3nCABYVLnVdw0olKmRUrR
a4vP/QKvvECpdct1QfAyijEoXK/WxPnQ1Y66d4Ld2+JIHDGIsytj4mBnCLNpmmuZjgOU4KdrLR9V
aQv2uqoSuUKViAEUZj1uFHpajT52X6N807ZMXtkRw2QdBETbpJ1UxBSsUBmcy3hLAPsPbUt9WTFC
iZYJ3LkNcD8C2yyTe7CpWPLXnyYGoJ+z37DCXnag8EJU5dygXK47hAJLVsKpWWf8CJWewRUCQOsi
+s4adjJrpxfb0HNTR1Uyd7kFzjqsGcOmz5Ik0QgQQhn+7/zibY64igpunwgsR6e4pK2pu3qbPR2A
dtgcHBAXUJi3c7yXkqftTjaU+/sgmTkJCdSUHvdmbccsEGarscee033zdzwymQkLmCusqsEcUvO6
/75Lhuo7dOq2KzPzcicnm67xScOKWfGEawbMtmb7Pj4GOMLST74kIxWy8NtKoDaksYc3qcjNeZl7
/4vDrk6VMCECCnpt5buebqfPbs5x1p+4F1Xj4irrqWQ7YY3L6+O3/1OLt+aLpWUNu8G39INAI6Fs
dl/ZY5KzaCCnzCmNBRRN0qeCSsLnyyg7yk1tGkkouW4GckvbvU2bI4jiP/vNQ79vTLPRB5BzqkKI
g2qcSBSOVFzHwlINwn5FrH/11P9dTAzvxPUzGferfxfWn245b5s4xSNrG00m/SnlBFyUERdBQW8t
bl4zA2MB3i+C8bX0rASjyfvnXal3WwAhKgmfRsA+yNOUHoCpM/kldrlXAlmLMAhvWbilDrxTHaAy
2BRieB7IJKJKYRMgEYhtFExDm/pmv/z1lyK64MIHDONpZl3l2XsFWMLmoibEVDjOlg3IXmUiQb9D
vo8lZDWDmnAPwdwndR9seatklLjrpk2kjd9a49XDmefjWIzhq0il0gDy4STD0AbnovU6b42h7Vma
bAXi/wDDe9Gyar4rOmVToSaNgs5bBIiK48Mvs2HR34nBfj/AX/j6OM3qV3nkAangkKCcKRt98dsd
3/b4HKUAqyqu8SQVXRQo823yK4XowJVmmQsfpyBxv+hQFB8hm4AlTE8JwH4Xwoqv2RsLd8+9dFo9
DnV+h02+Cl8cagJdHiCllRn0cqpAw36QiOx5nW4L3oh9sIcEBQypwrhrpFsF/1nrn1BRCxTXsv54
+3dmHr6a5znkwvBsvT3DQE7RnmfN7BmmuJQMwHJZA5y8pcpQuY41eVzRgH/3UEAz8EsLFR0Fc/LT
SqbQMEfzUJCP5L9tolmyeFH0ceS5iew0GtbyDVwkn0RJk/ABDvcE4ri09APofvNveUsjG5NLhfh7
Y9Zb4lNqLKOMcvMrbIAaH24uVi0/pfwbXTWEjZpDXze2HgSx3divOLGsJdSsSVYCJdeHEgxT0rLM
BVTMtXW98HVkOuYK7Du3cycnYajmxbtVK/YiOP6UkzgO721mL3WAqc8nzLEYc19Q0brJ7N2fi7Ym
b597yofn1c5rkF2nnMmBYD/lsCJ3/0h5PubtZQTKPPpsvPGseQaF1sALirkfc70ZGxZ6izL72m+P
3ZgNyCqdY49JdlCxDaqjjpvJRNYNh6elwbHaErzbLlgRYu3JMXEm4sjgSdMPJyi55PzrBhlt3UOY
y7YI39MgMbcMYdnttrMn7leoEsGpCOYb/MFAawWyeObermSxe4joHiqk6uRufOwGgfFeII3QO6Dx
ce6Brr2f88Q4qq364T3XGpZRdiPArRvN7emnmQmT3FqPdXarClwdkizX42q/U3yh+4wQuOGrzl0t
vHyH39SkOLoTyuvrwuI01qAk4CyoAbKwHDZAxQK1UkLHCLFqsAAs0cOzbVydjz9SeCbeGsmv5cb8
Jo6rG2wattkpi8DUoYHmoIyqSph5IGKEcL3OPPoft6FAJM1cBvouZQq7gjisOcJ4W9pwH+cZMtmY
b15Uv9RHY4s+vi20z/7tpQ3AqtzfRmf8I6NAc204l4JdnZFNojMffQMKBvItBBB9FBIKUjG4cGCh
/WgICF6p+ZGitRGKSHBUod2rtI2LOVY/dx8up9vysd6ZkQ01EGrzOTJTIe97oRD1nLEi66AJmFSz
b8ILDcqzKs5Uxa8rNVLyMgw+Wf8BZkxFt49/JNpeQalFhXVEEIlUhKP/0amKc+ws6Y1VwZYC0p2X
hyDSynCRapaPVzRKeUl8GBiNplEppSpTZvoO1oZk4Oab6kCnwacpz/HvABkTDLH29TuGY6khUWx8
yaSYyIYdUSfCVO8gIhDR7coNuzrt9i9jxAEN7ClfHY2S7Bpnj5XuzsdGbWklwTDCyt1pypfAampe
XNZ/QxKLSJ/VDl4/Hg76zOLouqxuzn2gt+6tqwq+WhRTGRcvrencAgvUzoI76aEPTkl2WvYqutPQ
HGcGKaMYQe0EM90NitxawtrRWf0ik+7oK2Gp5fgw6SVb2KgnKSYYaI4e7xIZVM6OkyUHVSkbQ/47
vNDbnOG/KKNUNqkpbppEJlUuLpxyanEmvwkiLe2w+s0QvFw/fckpzAZ11caKSVpQTZyChQGo1PY6
Epx9Woo/wriMlnruYMm1GWrGXuToWcY/RosDX+YYuCSNgpoxVOsmEE5GsyjKg9r85Lpj9vEpS3uh
b8M2GunsYVeikT/O/vHKAet4/GOWvKIYrdbAsgxZC1XSnHkcwPK5+wzmkNJlHJfs6gjRW2p7lx1J
56omb/TWtmpXlVkGWrAHDBI5F44ADRac+XNspmf3Aax+E2v81MHwGp4koae9vnVxjEf1Wxq1aQP7
c7B5F4bsD1POZo6xecq3nyNKW2hl3KcBQxWEnmPoyWmzFy4oKGQwNfB+zWLr8zYM9/CkhkQCez7u
V8ProypojknTqisFkwPYvY+8fceU6yaF1fqFPXBUjgmN32vVHzrJ+n7XCRYwvjCLa1Ums0tLWRMX
P+LFNJC95W8nwr/pnX6kK1Oztlraebop29am91my6GqVOkTTb9NX+N2WIpTB6jlh31EIw8UcT19p
yfcOqA72XOEQqgp34XV8we8bpObjLIi9ESvDpgjHg0WkQlF46VP/SPMaBA5dn6mV6TQV2IoUVLhm
HsGs7tYpDOJCRfwLV46s6Bg2s5m9R3Ytl0BsKPmeQ/ds5EVI/juc9BPZoqbbJ1FdnHn99uYH+QTi
K7wAhB6iybX9JyGYjvBKU5Oh74ZNPZoNUputujxXh0aQCCsYLGi0jHbMk9relgM7X8o0hH+fPj6V
1omE0KVK6pvun2Ead7S5EQwfLv+z05oTryNkAkx3d9kgm/mlrjXUL3GQ4hpfGx6uO2iXUuhY0b3E
4FQ6oAUD+s/v9IXrs7k1UOdypokE6nnNmSJ+MSnHOn7IcRMIaPO6XXGi8I3clJnhvX5kfDbYoNt0
XEdRYtpFDNrtklRI0pFQO3iWlvB91e1oP/H1Sf4O9lFIjpJB3T/DOHjzOE77mYd70+z7Zu6seXes
cWcv0mxQHEEqFOl4TPftfWXBTI5OmNNES7RmsJ4Zz8DeKw/v6weZjVrY6da5yXntyAsW+TRAw3HW
swLefBNU4R12eClQRn6K2cIfkj0MPjSIwUU2Xx1b1mMpGv02LIqus+mbF16LHWBH1MpkjXKcCrHh
wCeIskaXj3r0GDKfpkx1ITGH8IT/Sy8Wqwunn8UljeCuFmWy/wrYaTZN7efwsAwKUMs4dMOJI4or
jY0Ao4BKzR/cR6wl7Vt7sgolLCEXZvNvHfakJqrEZQgaV4JO8VILyizGHeaeUQBZYU/A/MagNmVX
xy86GMMD9qlXtzZahFP++cqrTjVT9nNZnCSQ4G/3EsCq13i8Mhvjf1hrE0Nc0NZZt77yLfCZlGCp
tq/WIj3j/nyT9izr//HJmFxV1wxyLhD2L9sgWPOeylB4InVJZ/YLq0gHkFtjy4NF6rIa3IK9hSoG
btGFGzvwuV32U9eOLGRMy6lpaH1lZdUU0sqe0wZUX5SmB1GtNDv/1pEWKNyljeUXHYZD74+7P/9K
FvDCdORQDUaEiN7Gg/VlB2iLqUAvAlvMkt39rhlGGtvbWlMXXNi9igp8s5qsu8j3xG9aNRT/5FKn
EVk5BX9U5PjSK25KW4YDbrcmZ1Tp5uPV5fVRnTFue6stgQTER1VEhR1tOgegYrXj8ckl9XoBiIsL
AnqDGaca5S4mPpIzOBMmm/3j6ikuwqYyBAzxdz5j/bTABr9VQpEMz/UkyotbnMtB6sFyhRAIqnED
J/iKbw38tZApe1uzQFJ9mz6o7PLHMHmnOIvrK9cDmgsJCST11EC1B7vc6ZBssxgBD/UCuAGqKLHX
q/5dc5JKb9VsNGfC5K73o3RpLPzx9soQ2WqxhzTlOktKtioORH4I8fTXclVDJwpa9wqMrRITcgWJ
vi/jEZvJpX3iK53hwdrn8YVziEmYXJ+3jG8f5ONHlxK3TxLwNy0v5ipGiJ7byH4HscHnPd86OOUQ
VqIjsQU9E5Gz2Gy53IngDotx/nb4A+lUB/KBn57cXK3KEr0nPz1yeLURUGVQj4MkADuHo4L3pqBq
lEpiHMsstFwbNGBc/gj9qKJ4u3OAnIkMDZfPJVPpbTaRtlxqdyH0WrvaLOq52kP8bBplXDXXaVy8
BVY2xkX6sL1iemkP19ARb9Sak4dd1CxYN4EHMEBQjaEnE5y1knIgeSromixrKpKYtv5tXd2THaks
bRa8IJXhc7BotZC/2xY9QsVWzXjtFSlHc5rPSYIC2A//B9Ei7P6uBlOPvyPBs6j27DYzck9iB63V
KT+NHfPRoF3UBtCJT/WVMbILesb7UqUxf0Ei4AJ3PXg9nKtNHYhAQmwI8hP6vrFaIgH7PCQ8IIAh
K27Ek6EkSb43GuaN9NcxtoQ9dGj/niHNHxRvU5UoBSbuRCMCN0OhXkxCQeFm7HcPf8tjJmMHJEoP
k8rtKzF56ICftGZgNf2m0mhOsU+nMLkkJPw7pFCDV7nncafVY0RqFX1Tl5D1XhjmJ5FXXbcBhAK9
HGqfmdanOB4BmkoMaQvuxWvTnd0kHoixECCHMSH9wz6Ghusi6siFYiz2hZpHCgrbB8Ny20D1hx1X
Vs9f0fDJQSNloymSmJNftOB0zwsjciisuc21otQSu9xWXWrPmabJJjSPjCqy5tShLH7PxLIB09tz
840AQt+c/NcVaK03jK0CTZ415biQPaJrLaUWoqsE61IdZ+U/8QenXB18/wdhM4/FLg4MgmZG3Lwy
KqDZ0ONMgUHGmn4HFdo3/Hrt6LngWb3mX9gJ/Dy1+wJku8NNRz7EwEhrYymzssfRYFWN46JWRQES
OHsxuQUzSMZA1kg0Dgx/u6T4g1STgq9gnqtL/l5zbzHMzpT0jVqBvO6k8dVi44jCQBEcGn7gNNL4
jeXkAP0HkEqmgwtFbB4BgsP2skDVXJXOpsAyNPPlus5WWv0ovxIEk9c5+MEI2qIXk+RtcfBdPxpy
VKTeUcguSOB9VOO55BRf8kV0vgRme1fXNtb+dR1GNAj4nwNxY0txg5gW5DxyL8IjYuoOT70IpNmV
qes1AWSC4ii4UX6OE5mNoqeKHC3A6V30YZpQ5RNqF879n3IW8qdF7rjGhEcrRCAx3Xe5x06GuxYY
9vMUrobzwXS4bWqOY5JzGdGjYq0+N+3h8bBaXpQ5U8Y1fHKq0BUB0Vov0aVtYthTvFFhoKtjIsGL
AOIFe2vvB4FyLLyMgy/7tlo78e6WYOPfZzUTksrQFr4Hm2NCAALDONlqTLj3uFb4KK0ToHhr9I7J
4kJOA0JVdSyrPqTL/Vi5BZrbvXh4aus5Bq05+I41/sBMbEMCvL2hkSRDAMl2bYft4QYGFH7Z4SZE
QAa5pqjVpOUlzehXPEQieZMBufyydV+pXRGHVe+TiZ5oOSyCDDAkn2KYuEAkO4gc8IUkJupV+PlV
hAcDEpEPJY531mQgn4+JvPj6CYqQ06iWraAL71Z9LVb3Lxdrh/R9WnA1yztrLUOfJZhNFZJtePPh
FSJLFmQxmxlKcE0AjZl9IE6mupq0GlpLtMAeZrQJzebjlhFn1FGM93oJJTBHTC9Oc+zph0ygeS+Q
i958jZ8x7jHB1MNI69lb/e5zZG7jtwOgmw7ZqjqZkHND5jPME0uDsOD3yVPwAFgTEeD8StOwKHoA
OxRb51lBtJDtONv1fK1iScwmCUtBXrJGhXOR4IyeN522+futsjizom6Nd6NA4xbVi3Me/B+fL4XK
6CLmGvlZecD8XuE97ieA3NrrA5uShgDPM27Hpm7OJ7jvyx/6JghT3T/IQqoZRozEYFqh6T++yzTR
izv24YrSJ1Jljiamjypu4uxHNKL2K+eWKyexzGfTf+zKaReYK0lYyyB1JqUSqnsPrkR6BVQMMbR1
Vqk5hS+cCDT38SZ3PfgWItSP5uMQGDBgQR2HWPW4Ne3us+pHCiPPn3pvSxZlVSWtGPc7BmTwu5O8
4scbgUteUdMvqR3G0B6ty3KriXwkitFIWlovgfBSDO5JFUt2T02dS+zwHQnsGuhDpMHvP2w8m0qr
fb6oXJA35JZNnalp7qWemiQX1jDkcbN1v0duc8sstLVpUrNcrU0m/DlYT/kk6e+o0eGWoiBp4uZI
9IOJ//A8teHOYyHLPqbTloVt7FSxBY+EEqkBCwizhCnYuXQkKxZO8yvm7JqvCgWUAocqozc9T9s0
Pm7vq5A52u4jUo6hE+kt1MLbeaILoLawZGXD6QBiE4tvKQm/RWu7UjSl6V/plLItMKYrFLCLdBoe
JRzKJM2EolulJmY2nfpX5IgI/+Ss2kD/2GwWqPZ1GQ/IIJQdM1LxjQxkrm9eHFPr8OzHVHLhgDP+
yBaaJoXVfNv/jvQqm5okk0CBWIAbTnMY06fDkFKurOVrhiZjuld66dX8fpnq478wk8liz+iXpp58
rwC+loF8y6BDnfDtpHlCPlzmRCnXVIICo/ac9uvzrMVNqL03JtTN+v6R05DOrlIOYbdAxWPCMvHf
Bhj6RtvH4/ghy7W3hZyuacX9DBgvdpjHeWtiLlWcRdeqsH9jvZYIgc+vdj8vTJXoAKVeVcS5BMRf
7IPtXwFLvDdI1pw5qwb/FEIMB2xspaAx7Clojv3HSJ8K+16UvV5jJOEIWwyT/NudhO9dcZcU72Z+
YOq9HgySjoKc38biAhIm2gtf/vCEbgHGpUSQOLk0h6AKEc5ro400uTHUPqX5zjvczS51yqDlLkMO
PbrGDjYN9K9ynQgvbMOQtP0ZPkRUHIj4ReFm/x0H4M/Gx3Fq/nexvsKoDlzWFnsb8K0iDkxcOC5G
zNHR9UwNN0sY7fDHYLaOKA2itQbk6BlwDg9kn7LDC0xRZkA5GanDbP9YJ7UreIYihXuBA6z+1EaL
Xv9coywEhXw26ODyoDE0CsJCPfYL+yWBKgMdBIF6T8gsdteoszv+M/cNgXimyb6D6Wa1YG+v6XXz
8PMVm47jGRd4BB/LhlVdZKbFd05/ad6o2Mw9PAptqcfyJVwDxnV2k8bmKQV+xDs4i8UkhJ28UA69
DXSXzAB2BK8FljSjcoMcg1Tt72Tt4POqpM9S6DnTIPXWgIkYHRUxPOjf9ffD/ACwzBEjjfiFaewt
1A3rd4s4v/MY5avdCEDl+I5765CeJtfsaDXbTY6ZH3sqORo3xrfMAQu3scm0yfWgfk2nge6SzQwO
Xh2+//FQKL4rwhePGq4WJrSHjfPMUmLq44sgqZOB3648+S8QV8jfeeFSsFQHK4dRaZ4TRBjjtFRF
p7kn2WD2Q20m/2VR/LofELF9abWq88icuNwyQ6PkhM7SQYItYiJJKruGqkcMBeGvXnrz2QHcdZWa
54YNgWQb+DBeUSHqY/CsbQGBtpfNdKPykPG5eOqLzOLsQ1yODd8eTifaGOX8opjV+tgS50MFRGjR
vJ7JklLdGZbMyef88TxSU2auWxNXfAXHPxLZolIioFsftEn+7Inr+295fUikQfh1Kx2anNMe7YmE
3Qd8KmhaFZXJrCJdVpBtCKLGDmIS2QGJfm9KPgguWUNQb2kV3omBzMgI0ZZB5nkctv7wf3G/KUT4
ttnFtN4k+TCWswCs5ahVC6qnFMnjfuo3O5ldLmZq5keYkFJhFHn8cu5dlDKAp/7F/LsKjcSV1L2k
pBYIgZlk3sm0zjj/TRN7AcOshRGr+EsREhJfFc5FnbNyK1qOpUbyMrDlb6GQcMwqMqqrGXzy3zUU
u4OXENTh3fff3AGhqIfvgQrib9H3YDjX2Z3zJiixgP28mHpjLR4t4czYlpVJYYDgyoBYr3iq7Ntn
sASkGN/fhfJjmJAHRssfMeZ6Kcjo12GRkUEiUBMtXvj+lQpnn+9GvpvwxPN+90RDcYu1pW/sWNC5
dzeqDQpNtqt6+dzi3b94zWnIo0naIvlrvlhSXMoGku/smNFzfHVjMzMUiZiJFKo01e1WtRKBAbwB
QwdH/Rj6BwpCBA7amDrVfYmBxKPLN/h8KEL8kaKChEKZt1KuhwGYVGbTKa4EZ3QSUpQSLfR//jiH
LHB+3tSPHMXnsdoATapr9M8BcVpGw4wVBwR8DdUL4+T1rZlA7ZzpK5h+A5nX8h30yqQuYwhZm3t3
PZYFb0mtXLlBzQynIe76VDsSuMGIb9KV0kAzmUH5yRZIppgGQkva32Tlbyh2PCGM/NOGnGcRiexB
OXWixlSS28hWy5KPDM529c5KsHqX01+KnTb1tgRW2uQTbCOQg0O63CDWbCLoQDF774q2+AqhnSDA
0seiAhfc1Uw6mroDr4PTzd7Dia+rWIeHaQ4SLdwuDjYWrEriveMwMcpsaIj9I2/5Rhy+e/iFTVyD
YwBR07KY2YVSDJa7RhuhoZ/e6/BIKfdt9px4dIVoyX822pshoNnymkXaEO97mRwgJiTDEbtMULxh
NAKPkJYR/P3uTUNuDKND6pGwXNBoi4ADnyjdsb0WDEJqHwNBQHhY1FXZ5QPVxz64z58NYf/SVFXC
oIqQWYEPHrPqzsYnq0HW/2neJmxqGtk6d41EtgUnAGuIMAIannOkdVexWuRVL1TMY2pXds1Hb9ri
QL+yFHjboGAktKjRJMN5LC/tkW6KESAhLVmjpqSN39RL+r8fj+5YRklxWRryruGBbVqU006pSy3A
zdWGLxzjTxne5LqY7z+fzhlY40WM8nYfS4cD9izR43Q2uhJqnOglYu+GSOeUkXeN9sgLzrLYfxAn
h4vXgAb7r0W7j/3rCRgZOkngQq2RnhAvMoTu+i/frbxQsa3iCWxNjB6ntETcdzIKIZNCrsoQbuW1
MbMgk6X2cFA64RsZR9IHeidBUP4SotnajBuLC5IT3HL0YsehqHa2k55iD0m9JsaY7wpw9AxVx4uU
BX5RVkAWvOUfrB3+clTYUw5i+FU7+9eqPpWWlvjNymzWGbaUnRrEzpfNOI0g0UYXIAlPBbC0+SZ1
eWaFEDkraeBrCO8cEyMelryTqx2wVj2OEWStxwdco4k9wA4k8MIUv2/HGacc9vrOmRvDcfe4h5Gg
p5HbkAzhEglnQx9eeg6uRSsc5dcaLjzwB3ABI8pAoRQSfaAsbyaoMw8OGF6hlWN+HPWa+vH1in2m
mhUTuImIB+pxNoJKRNT/IkMuqiq5pGcRQ4nX/L47Us/uSQuOhNI02rqBS9AlNw7vIJEzNllFUcos
QhHvUyLg3QdO7g87q/EmhjUGaidjNBMVF1ETe81Ch6CUv4i/4TS4weF3eIh7FEOniATnpQo7AXux
RLYpsnyH9NBYek87OrKnqpRInSa500uSlbYRQZb7TYrlOC8cMtkLbwP8V2QTFvHc9hs+ila6xyxp
zfQDtEsO/oSnRJgBZh5/wEN1Ookxzdz1Kei0wM+7wcYwepa0TK6H+x5J+qr7qaqEEcSZy2Zo1DTg
capD0O8RKcwyDJujimeFwZi9uZ1bnYg5bZqIpAO+FveSXod8ySVvbEuuFeE/FGyRIXkAX4fcRh5Q
3CorFX8a3zZztcydm9ZpWTr0gkwL7KbablJm2/ezzbIHMqUSYTJnS7DIFBmLyEHKWZGH44Z8S9OI
F4tq9tBx63hiGwfCG7fNl2wVee63ZjYAfnTjxDs5nuT/AseZHI8Vt29jsRKBTJjSsa4GQiIIZlUi
DpyaCBeY+oT/nfrI0R03VCxl7ub0BMPP7dpHzcbDqqum0SpBV9qu57E5YF+IYmvEsgXSto7FHJjz
8ovSHLp7LwYQlcXqAuYl14nmh4s0awoWFijOxmUaInIJ/SO83mXg2L5jwTly8TT2tdq6WH76voUg
+XsqMMq48dVo49k9kMN2c2f22AOTop02L2xFJiT0iRLI0iNkFPyPcZkIiy1sPG/02VjL6ERQ3AH3
sEtQtyuvnQ0qzIJEU8lkuRbtrsvHfC4a0gBvoDv4DfHGgaQv25ISCqDKrDG7Inr7Etq609Ko0rsZ
GGIqV5zLVG6LS8/paYith/3Wi5+Az84EweIAKPI95DynemQqIGkhvxlFgX1EAJX3+RP8b5tw9ym6
MtAjU9uEgapTTokPFMtoyVTPtGzLo+KOLqsXCcZx9sTxs8130ETtUECNwqLDCdVhIk/hbZM1MMd/
WCa7vlp2ijmfwQFXcyOC0aJH+BbK80zuZNTNYTwsWiwl8HKg2uz9EQ4lg67qOLQ3gVvY6+IKR5ta
mzGEJh0U8+XDTMOVcfQiXJmFPaIuP2YTOfUkgl0FPFvYUf70pYkZNvusBey/PfweZw46vdNmQD/Y
nW/WH90UoEpMYHLnr7G3Q1CWDvPNpCQ5sEKD7a8X6amWwrZ2R05yg725JY07Hjkv88AXNBeBiL1q
Dr9Rreylalyt/moH81qjXM/m4jevHx4AH6q/sOikRKYUWXNeD4MMBM4GVa2LYA4Rw6m3RYvpdbmb
sq04Fzqa2ks3lkFz1sgcNX6P4I+jZxZMdl9LdU4b0e9wROtPOTVcURnZo49fEryXCaFqeS/0wgWI
Z4wcdOkHPcde2EBbWhi4614m+HzMODUNgid2MU4zDHPfEDmsNJoOBBEBgFFL7auiKmyYh9D/Lwkj
/C3eQX4qg7YA3OvQsdxqG7TEOqd5dFhfBhstqbk8ofTFewCNh22ENsB74QmRtVM1p/lzPs62ffhE
udtQIpnXD05SXZ57zXbUuw9Oc3kGGF/dUDYLeKcXb8pb8ZuQzheyatJ72dGAucxtUTD2nvAVp9Ue
TpZmDjACeoWRCRk/DsjMw68E60XiooTH2w+p+IQhU2GyhnlgyKNsdQtH1eVjTuRq5IYWeJW5YDDv
NzQlgwZd8yqd2F0eFgRfGe+LtoKC/Oby7askw6P9pavM13uHNGsxdKGVDjFgoFe/yvBmECWBRDyY
FxMeAVkgrQxwm0TQWqJtu0z4LbdfUip4/5B9TA1641SZ9AbKf/+qbFt/LuMZL/Hfc7ImMiAAdB0+
Tkp7GXtAsGrnJtfIfYSkUeKGQAzqf/4TssTrsZBdp3cZWDPnb080skKxi249+ffKPE8Dr/C1Y8WW
eaa321aD1S4XVvXSZ7o5PUrf4ECPiUms41nK/GCNEtwMY5x7SvT0HOYP9DhL80zzO4Kznpg+F++P
0M86kXfV3GQHt8hwR0tLxT/RpWZeN8fHT5GNGVlkzDWCVlL1fxa/kSs4go0KW7bYL7mFdYbBUfJa
LWpMheJbW8zbYJ1W9bnH0GoY2LKy3nOPEVjO4kcKNYSltIqCpvZe6tkLY0obsbFicFlK4vJyHXsV
kF1x1XYggoCfUKldMI9s/zB1QSdJzb6rXzOG0yzQJVPDmEYZyVdB6Rjm5rSt47MiU+7NQVVJu8tm
eeA8rx6YUNuIh4zhmd13m1WbgSlWATYzsgeVLdnTkGsH9yalDS5G90vZVX2tANsVIV/QO21t7mDY
EMGQz4G/3EIpgnecFZRup4eMJulW2nA+qqn3FT8eAMuBGfczxYbE9DYdRKTvWgGrPfVCyheDPj2z
ZWFeMzHoNCzZrtKViEDgzaJDeYA2LXMc4bMTkLvFl1OwNLauSnB4kNHe1CE/p+x+8Vlbl3t3QiMP
TVXeDSYGH8PyJ4vPVHlql/fwR1yq8i744XkpKCrRy34/yZR1QPw+EEzFfLWzfUbwKIhLbefufKcE
XSSfCRq3UTabaCdGSjz9JG/EDGdqwIOPZusqN2w6vIBVcTvMiXoU/N4jtu6n/ZQ70K3FiZp9bh/z
TNjG8BDkfBggCUwBW2MF3vZ94C0yidNU8l/Ji4on2OGrof8ygGdHvR5hTzPj1ret2dNJc7wCqQI/
0d2UGiFn3fA/F2bDRvKeo4UWE9+7WGM5wgEUZP91/fydVAjQWHzePRL/tfRyhCvC8m3Yr+QgAeyV
QYqcpway/svC1cs15tyndI6t714M+HO5Rjnlrx50y829+cGDdCPsjqYnHORngJ8BPW3O4SKZpNyx
ZZmaLnDDHlZA1rW6S779t5iaok1OXBBYdbYjwUviDhEup0Hy13pDdm5cvrWOrw7r/nSIsrzjHpwz
QRHXGzMvxrbJ/GMWdQUEfuA9LMigFT4uyrIORksTjEPtGw4I4QQ/zqQ63sF5WDezCfqaSVXS5FC2
qag/W+/pL9tvAPEBCrun+tAvHMeAylewK7GI6wBqqJiASrbvXUGcWB1vn5jy+WoIviNuv650462s
AQeTSgR9vBXm8+4tRlbAvSCrY6SzIXiVIkdPMtqH0eKhw3xtGWHvaGjtmciZyUOVkKArS+hYBD2s
L7fYhlG27Rg48Tpk1zRl8L3vrTYUrs+55elXGp2ulUqhVeNTtJwhaI1mAWawrck/iAFajRoWSEVY
S4W1Gb0RNzCc4zoaufF2LA8UxgfR7CBRajm8+Mz7zddZft4RtlpTHCpsRjZfzuGzRAxqkVVnsj7c
eE7l6Gf+A3k4w5VzPWvVU+oD1klDBco62J3OtmbKSV6xKn+TJtTN9ABNk8IA54aPWZIwDYNjNgkM
Z97HRbHAfg1vvFAM/ccEt8HvdjWQtgeMnW19rW5DVj/SXNzfwolwsSQ83AQUGAH+rG1TSvGiogiT
ytBRMAStFqhTkqRjyulxYFTCNE6TTcW8TmJOP8YFq05bwW0imj3D5ad2RkkwAjMZ/ZcKKq8zsRnj
35BcIXAVLm4J2qgG9TiHyUiSPT8irDdigvPblmCuVhvWbUKESaHuFx145qbELDYEHCUZMsCZK8Al
9OMuCVA19GXsfagc6pTW688jABV9VRWDeasN9sEPiOWTSpsUcxK99FPTJHv/bZDfhVV30kdL22nz
u/jltWdC7zcdgrcFqyY7eeFQfS+bXSUSRE2k0ppshLOGWz0miuxn/9hm3L6r5x32JQoF15JrYk1I
MDZRSNBJnr4Yt7ziK2sTV8u22jNzR2XMIH9Wwnf9ZfDaXtDhjODkVKbfrvymwxiSy9W9J1m4hlHJ
HOLHYFYEz4sVKXQuyoIU9YVsEIYWtUreBa+L3B/gbmyhUsuWHnPF/MarnX6TpYgRnq4DwWSNCowO
SMO+ERF9gZ/7s8uFq3+b3N0yr9L9+crsw8vT5ONuuX3ZI2c3Ks+HemSxPH717auIdvFF9oOZZQd+
NhQKcL0loNL28A0GWLVZsWmeAq5zZnD1r/0HftbkcdUgdMkF4iimp+asb2J4x8okGezGSrITALZ6
Igdw5M9/vddux5C+6Y8laR38OgEcL3VMuvq+xq+wmitzkx8rJJEDRn3ZwnJVC+TWnPDHzx6wl96i
5r9i3dCqdala68X4i2q53baNXSsqg1R3mnRLRcrqMyUUGUGRERfwqmG8lae4y/M34o1WBdp5T1De
fUZzi+ISiXK57aaSUYzN9Pgmgi+HHo9E08zLmV4wBMNUKqB1xbPDhi/3LTag3U9i9pVSXTpv3UjO
R0duPJ8oW2Ccv82M8UlddZyNJmsmZAu/v4lVBqAca6PylE0zCdgSztMtXjqf99InnMdi6uFIQjBw
QxKd/ou+u3BjCCLpe0HwxGj93nMeG3kHNXKF0anILkEZYrYe9alnvaCEB7AHLlJX5GMW13SeAHRo
0KU06hJqBxeuOkB6qEIAFECRM6is7ggOpIMCDtvGvOjK3AEQ3oyiiaKsf3u/q7etbl4aZ9VsN/Wu
VeaZeE2u30XAzNjT6jID3XgCQZAbCrTJce+xpVRecipBOlth5ETYeb7f/GwL0RZMbMJRpmXaY8l8
1j+k6fkbOdvQylSFVRTI3warROV84EcePhGnqW413Hyg8yiDKRI7f+8XkpKYo9zAKWQ9HDSIQkAs
aklMCNZnGw26jiqlnkVmee6MuCAp8xm9SYjdJsTjYsjxwkjlZ7sJDkyFOHLv7AlWFyN8EGhsUfCs
Sx1Aeruf/FFd9n28mYxAX2jxjnwZTmV6EG0QGwXR13V52OV75snPXfrSTyN99OEoBXWNmUn6qmL0
x/4IC+x4kykOQ5mJv9XlT9ivtrEpdgeHLpWOFAooZy8l5yh8NN3dVDtiy9ir7jNesT+sRZkIZHKe
zxuR1+bcaK47e/KoxfVGzoLMnVw/9mvYb3abyH6K84Xd3hRsEIwtRW8iZ/PMwmcWGo9yZy9IOFTX
aKuz2JqKTW8//F5vdQ9VshqFadx25CByMLME61p9nVqLnyHTgYrKn2Gs/IWCeaqJzfumML/HN9/x
wLGyRq1rY/Xzg8sae7rruioNzRFqgLbcOsQYeeZL5lqjtjd0C7IsjF/6nZNPWLSfu46toQGnEOJs
xx5NueZcWk+xX0FU47miYC2qocxpLFYdZfZ6u4EMtAd1BdMt5S81RoPquwjTeap4rB9zkYpOFVNY
BgJOv+DT3mPf24S7pj7j1V0n4pOtD9e9MdpWwg+MLTySQkWdbG1J0Cu3aABO/5qwKcGec6DsmcHS
oq05GRPF/eP5yuW0NKdwsDLkDj4edYYgRVoTU6LL2VtvswCmwfQmmT3BKZX40PYqrTD+pZb+BgoL
F9q5fmbxG3DwxVCEooa25IjijYNWr1rg4IggtJ45qQCRd/xSYgrZkq2qWNLYZy92lG0tspLF0UF7
uvy+FAMu12ktKWj5mBDT0wMRbuT6lX89D9a1q9SAddPKE10lfONFySEC3ggNenAmDQhURvB84RXG
shiK9OsZHfrgo70PUxwT8N9R+z4uGm87kinEhSuT5FQyguIKnW2k+4gNrmassmJH2ISZdcV6qEgu
hvsnbtU9JMtux77vtqhLBsJ5/brvlBg8K5mKFtT8yVw13r8DGPDQl5vOywfHnG6cBiHOluA/tNtU
vDEhbd6vQfgnVkUlmdOxh4X3sDcDj5esmZRMq1fojdnmgXEmmcVSDae5XLlFmxaDlHlfb6x6PWa4
q20Vk35nDzdbsuoi3q7B+z8XwIhqbBCb9nSI4liNMCHd3nEC/UaQ4xye9TD56qgXwcHekwiyFD/h
7rLFA2yxQY+UhQD1IIEysZpx/3LaWbezozcTg4luB52z7PgCwe1NBgUl5CYBdgmZj77F19K8Q8/K
zWD2bWgCl6H21n+I8X9ZeCp0x9Hy02g0ed3AEtYip3+ca9PR5vD7aVMalqr1pvL1MF39eZEvN9AB
RvEIY6Zmj1oqGrqYpCV1wUJGooElgIw/zaGHvIAQKnhLpChke8n56d/0zcL+qf2DcnuI4ByvgqLc
uvXv3QC/QNoJ180aJykvmiGfWMbK+6qM52idOwqOIo6aPBhYFObHib6vmCqWvhqMtJJaqaATfnNw
8eXNyWIASM/LI384KcMp3iZ67bsQPzmxfL29wCeV+gHk4/dy5cKhTt2NaLrZBhpeOcVoKLPJbidL
Nf3EWtZIgCs8dJ6LYMUS20cEkAHTPW+U16SKGmZUeFaoFQCcD58mj3cc/PDLLFimi+2ENdDDs+bT
Lbar3kXiuy7inEEr78ieMeB7I73D/ZQ13ObBn6JCZTti9AzcdOx/c/+kIGyuXHmTOogSM6yEAsnl
H8mjup+YJy3TeP7wiqkr97czTHD7RNNadXnTkZgpGI+7VRoLwLgYcvMPD8ihalOqEG3kArZkofO0
v1YGsR6DzDpxg2qNbjzt9TVjjgiHROkPnGxkohSLm9cNUM6xD4NCk3RSxeanr36PmViGotXl+Wue
4EWzV3/4Kgm/o+CDG1Ns5gwZHoBe0idWNPNLzEEexmVMiaX3j+DjklfvWL9ZNJQEQim16VPuQXQk
QWW6/jNqFSlEwHdPMnCDKEzT499arIRe8oNrjQzmuSGhCb9H1bf3/H+NYzjhwMlx1Z3rlgoxvj33
6SYd3/Ue4XLrOvCdY4aduGTqIf2Og23qz7gMNBLC2YJ+1d8QQ4km0BcJcvqFp+XFvop8FPYZDihW
anE6lWnC7cKle4LdgWu2Vr8uv1RvU9Z0j5Mv89++C/HHyZHlopIqXbtuFi8cJdhghGhna1b7DMhJ
ZKYCQYGVEAshQYaiHze37ymVHCw+IB21ddx5k5lgcK3mLUvV5u1xUfjFq+8FakPfFcViaCt25PAo
gAdxxe89xtQKp3+G+GYnl8ANW3GXGy/n/v89uNN5Quz+Py0PMMhrek1sxhJyMnP2bK8Xor5aJyfp
LyuZV4lF/vNGgmysXaEajTeqh2hQl42KJWruqs/X5irf/uqOHECFDcP2qfCF3f719rB5VsNIebh7
risAipkPpQQ6GJofSr/7lWjKvyZegpy5Uc6KTOBax1MjMHtqOaYWSmk0rsP5pt5mC8v5ZG9NpHS0
23eQ1Is3gQjxiLpc74z54f6JEigHSPE3Lwnu0jS1NONPre7aG6gtqBwG2F9t2+Abc1459LHomqTz
Zb4tNMjwOV3dTm6nNxq+YATli9apIYa8vLWq37OVS2cO65+cj/XlC+PhufaEfYsOYte+7kpRRKRA
EFAedv3HYx2tn6jVtkRef6j02+vEWjO7sOYj/dFGYMy47EEuNhvbZmFU0R5QJgN8zZ29eXxAVVvP
T4uAYp7zB2fNqRwNUllI3Ss5XnvLibL3rSr6wp6hVE5VwpXjfQv2H5MeVW039Yv8NT+4GhhQ+TNU
Gqax1WKWagHfvuawWqLNUyCb5hR5WihzTP7nDoq/nGp2exrdM05Hd8QF4Ce7ldVJFaXhHk9Pox1H
8Ot5mgatyect5bmKWJD43QcID3cTKXyhg7+jhe3UdoebP0KLjGg02Ky39l+Nk4Hgcj8QVCzjLPx3
4ThYApKiW2Z6q4UWiI681ZVXymjfzpjc7kXyDqjFptSSRDFqMm8BVmUJXtczgYX0oBDlT5Ms10UZ
ljOwt9CeksnrvEGneyplVcro+M3ekYo9BwcXhyq0zvrt7jgiOKRQp8dNT1noKglPBw7uz+26NaBe
QtlwxqeodBF7IXg2rJ296e2qbGBziz3h9I3hHUItb9aWskykiCFBsUi2Vx8+OsE74Q0ffJKgZsoz
nDzW9EYjzu2XsiwCCGxYrWiW70c2NeTS1dRZlbcoMJkBn4H+FE7C/ZYrr5Ji0OatlkyWw91/iH/R
7gO0PZszNBVVlHeKzMc6lx14Y+DidiKWv9NDisp9LXh87/cpfxHtEMs42Hnx5ZEdJolxHio3/OCW
sRfkfCMLPRM88uAJv9NC2lNcI5v7+e8VBcIEQXjaxXWjpVilZFOW2JGg5/knEv08yuYvH+79Gds+
Qr7vdRWpO27eV+aZmHiV8vFS+mVJ/BtCwFTe5QashD6NqSj8FGqyzNVtk1FxoQtRlGCh1Y3mFGo/
QOhW2lTA1eTzZvDw/4+7bA/Wq7RAeJi82bnw8XkUjwb0ncfQjk92sdOK+Y2K/xiKktaL5K6DQiKV
IWB3g26iJ858vo9nN6k30GNahboElDlcNbNulOt7tsbYr783Ts8VsuAClotBkPum7HE4mQSBdv3s
Twk1/2VaNdh5/4QeLtv4j/3LMLMIpBr6Yza6JROqZ5KvSTC1evseqCf6IG0sbmLEP94PtH+QRELH
J3X3p72Sr9wxlHceWOEeN1QN6szthTOSqD6LCz+/szr8wzU181/31JUxQr9nuhlkBBep/50xv0Eu
haGuNqO5Wbdc7zHvists6IqvZ9GsBACcnnL1wj2wbdBMCqk5UdpwyACpma6MXhJbScxR97RAExH8
0GAWLmEoFwz3SMBF5JYhqmTgI+uNzkhv8kU67RHJpRQzP8ln27ey3Z7brRbs7+NI5Rw1a+gEx3ci
fE8LEMssMyWFq9TJbb956XKD0cJBQaIIWDmgk9yxkNQmJV91nAcrpttshyDzz+HiirWD2UmZ99BB
p4TiEGp9JtW5f22yMVk1bdDLrbOnjZy5iubvHTVtq10OPFSUg9A3H7aLuqFCvsHYCaMiIBWQ+AyK
kS1YyEbWu+KNWp55/R5hvAo++BfTo9YPlWR/wT9TZMgYS02qmbsd9R6YeRQapNghouCEX6cXOyzt
KHufXoferdNZNuC4xni3MN8FdWbBGvfd+hpCZpDbFzDUqJZ014K5j8PiLRcGESAEupTIEA5DwIP3
It1ZJV/0B8dlW1Nrd6itlYwPxlQNlNDzszHSgxwo0JyIo/g8KfPSX5onLC9xvmLYOpOTXPVBw7ul
1x3jOzZaM2cccW935rjrWaLR/h2nqYXDC+ypN9J1dNcowk1ITwGDYFvkvCeay3vCXjuPDDAp7Uok
jfiOwkEOr0iOAcUEYTq5oB3zaczAARxOlhybjjXtvWeYKwUmbke3v+9SGuulAxEZo+J1XUSdVTx2
ESjuIa/Q8ZPDJrKWSoYd7qhPqy7IxDDpf3eSh2L2Gqep2PvSq/OWHFUn2vqJYNdScqHQHEY3iibL
QxLoQaCob2MvsW5+naw8/7KRofQxbG/rINDAtjHPIlNZXdomyusvgw9saEbjquFcQewLcVt1bXJ5
u0TjTx2Zs/KrBbYTz09u0JnngrrZ8eAsnnaFpYstHkNAiVQ/rREI+NQXqu3ScOfsnb+P+g+vyhKn
HUs7pRJ7uMo//MXY4PT7gMRMmndtV1Ab2gSU6sKtlEH4/aQYbVMlZru/zh+Hq81TxANRIvE8DFve
1YknpkNV3/XirscKx49yhXaf+Aw2qh1J9zBX5hfFwYmW01GigD+0rthCsGVKR90s+rUByr9gcbi0
kctiX+kzbf+y8dSaNMSZVMAKgW3IWfEtxn05u0NfXmWDgtluS7g9P3qFh7ARuC2XaDW3D/k9yjik
8gz9bevpMLd/Lk6nMql0Zcpq1/HJ5cCkQIUvcAqAaJaDLctSqzD5YvJYyioHu0Qb8jJaF/tItMay
jiHqV1w9b9T5mGi2cUV1DJmS7HXCXuMiS6cozVgS1h5P65UerxCxmsS8F0SYFRt5uNXRxtpZg4se
62kxrf+K8fqQPb/DgcK/cplhC1aDuZjpDWGkwBusCHkk1nB8Dn/JYuMY+HwfDYwoDsZ4R81/0rju
w27Dx823lAbFmfHZMZLKtztcv/FKUaoJkdstJ60nZYVqcJxifketScsLjcE7mpK/LBlg2vTWhVxF
Y8kOCTNur1yoG+tDLeKTWrcmaDlTwd14a3zS0Sxw6G9UTewTJqrmpXpcq0LCpM2orBSCDwm0BhbC
s1A4NLCtIc0eDrZw0JiibS9XaSpEN98/XhZs0gMIW96XmLDwEOtz4Gjt9fEsSEWzja9Jno1L9o6t
HM8xkeKQEbtz/Sze9u121owfl9p1qI/qOIvHTZ3azQhM0jsqtoXA+VxOxxLya85ygoJLZkXDj5V/
RE+NSPTxsBneh7okE6VD26D9jV8Qy6yPLtphBsDGwCW/eKCbLZRoZ9pp9pGYBO3ag3R3335KBfxj
zaQ8jErXcDDQDJxP9FQ/wvZnkBY96mI3C8ed+D3NeRBqMPUAHE6H1fdERaXpoLkX6vqGnT0g6kdp
btfOEu2lyoH51HuWe7FVgZaLhYj+KhFx/UK+kbd7LRg+UaBNSba6EHIrQ8R+Q6TTyubWBDY4H4UE
piIcB5F8qtCnuhXlwTWAv4grXq76a9py/DUbFsWyEF/R3UIW6CuBFahbiwtqj3kraHSfDv4JGRU8
zLEEYTK6a1ALHtkWLjwXuxCgFjkKgUEGBXyjDZ135PHb47uFTuE9KGnfbMkf4F9MbXLH/BgoDLCq
eY5GeZZ/vbRPBAytHgIrxX3h+TfUJuqwlbPj9YYim+zCDwC+m9y7edV72QJmu7dt9vmLO2zD+zdJ
1Kvskx80Si9OSG6Zrcj2D576L2oEZ1TAnG6k/k4DHkWre705QImQXeTuCELJMibBZLSSTYzMCdY7
80vEV9Vx5LyXUk7ZTVxCC0YKdW1BLGfONjQP3HliMmumxmZbyt+bqkgp2EwdbAERIWfTveyaqY4d
4KyDxzf+xdRQUh0rTMSnmMRSk6WTGdAUAYYmyOZB2vw0w0+OdMOBswqxFnJI6KGl874McKP4frjH
e68MWkSfUWUpxtnBrHIJwkM3AakrqfTwrQa3Z0TVe/MKuTnix6THw8TSDms1FkmLbQds0dN31SfS
boBDZeCRoJEvJeBcNpslfQqrmNOeVkYaVp70KsbDwZMarlx/tZWyugimimtYHk49k6MyQt0jhQiu
geJwy6ajOHZkww7vftUEUCDuxb8FYUdyPbjwVLc0dQVpT8zc92djqzVc6wZfuTAdt+IDR8bW/S9M
nCiiRuk/RCBqbaX29g85C++ezVImKtFqcgAQ4qss+fhbxWDZ/vjts8Z9j5XvgDRB/BiRF9CxuzKg
fcx47F4zNBjnmz3agmSx87CRFpBcRvqlxfckl/cqqTWaziwLdfcK+XJo2LIxilZ/1qZqO0YHmpFO
DqGDq9uFwh8MmlKjxQLznj0+Iy7JXipYhEl4R9vuxFgoDFgr+VOZThzsB7t4K2MZRzARAZ9E9tvA
AU5AjmnoDjLuHzhKFuqNWVM5Wk2m0C2ZzUsFkVaP+94Q+Fp7HhxRSJVRFfmsFxZU9dUf6hg3C4Ly
PQyAQV+7DGDD0hp0MOnNkhPoy7QTHw0858wm3UEoSGbEwkNUjwuyYoeEOfIxVv/oNUnhkDqO6NKj
ybk3RKLrquv0wCsE1cQ8s3pSsdYGuWrnQhdX7RqgIeHFmnIscMbU0eAzBprHyRYOjyqeG48umwDd
0loasxCaHCyxdxfZVxZTYSfEqP6Nw0z4zdqjP5POBZLKGB6KT/iRXPUYGKqB1CgGumevMCWVmKHe
sNQbjVOgrJLDoU94MlhER6Ge/SCTcZlVx+sGoXbkBNNKdubs5t+Fyn8ytA8cpzfBD18UIe+SlfRd
IXTr85bAifNk5sEdWkCXcGzb57xwR62hrtz5zE5m1PwW4JowWTBt/PAFhUdsnUm1R8woqyzVLnOD
L8stc2sxrPb5cGu/HHFqL0xxLYWdtj58qlgp/xMTgv18z2Bauy4iajaRUfH13tg8RFmywe3GlkXJ
al+0flcyTZP3gx/g0yHj85we8uzadkIyRJDRk1G3pnXVRkVaxboFPzkMoqYJDV57LvUdi0Dm3RVe
W8UBmxMxICif+ektUcdA0vb2NZzMlqfTVA+zuD82OIBU67m6HO+CUgCahrLxRKH2nidDC5AGlrHp
cw3NZZrk11cv4jmBKf76a6I8ODGAvVyIgmvMK/4KsNN4KbcVmhPCsaxUEqhN4udApF8IjvmXMnm3
/AcpmHyzwUEMY2i/ebjG1tkI/CyhIcuPkgXAnwYeSIuDIlswohPhsAVp1bW8MxR7UiHd8ONZ7hZL
9kEQbvzdWqCAXGo4Y3bJ2HwH9tcHfJWdSJ4AjQqfXTeduYoLNZqTeWOTGTcoe7rkMJjw5e59eORv
0DdA8jBQoPBO/1Org/Z21s+FXr2USm+m+LKgPw3fTMDJ9TV3kncq7+vGPJizE1BlGAztUdElcjb1
pwUqecLL1B5ARzgTlMX6EGEyKFJaY+ifqjn8MYSbmVCrFQhxIwb9ijru0WEyOJ5sD+XLS3bOddPg
w0gMnCU0gW2iCIfaTmv4PIx6gNtqqB6Z6Yx0QcDK/3CPqCRT+0ZNYtAv82iiOHfAc3VLgWuvbATD
6lAGxVogoBrdf/0R49ZF7yzBqDVWGOpdGv/Pj4UlfpTD9JBtz8/O8CC2LeubPUohU4s5g96zeLoV
s+UHw+Ye3TrPTm3LSQSChi392r4y74Xx0trJd3RIl7KlbNucMr/sRsLJhRXdlIvdE6QITVdaZSUX
m4Of5GVenSBq59pdghX1gaSp8cOOlvS4xVY7ogkxh7o/1g463OBT/1pGMWJJ5YjV92nXd40qVmd2
hZoDikdXuzGA/1NUleCrdSEj+0j1Rec1iGYKFTiLADTZMghyUtEqlWX4d+iLXjtE40uWc2IlslSa
0eDNm4JPj47VD6unZyiZ/16Y3tMzhqWku3QGmaJajmfjqI2deXmJxt7J2QamZ0PU19vy34IeYK8k
02jlGz0T4lW/ZztkTfvf5cz42uxISqrsrZJ5LFZBERz8rcEU582ZmcpeCV/Fo0uycdCp9b1x6t1/
ksqrn47We2ZIxbUPDuUPCPYQf5YCsNoInrtCNYsd5tqahjRiyX6h+h7m8R1qrGDjYewp2O4v9smy
gyRwfIRpicttiH+ZwNveZqJcUFiRntSzPAk51XTiJYwmBsfdJLwPDZU3X80CTVm1WkQjdgB3D3W8
B8KFahu5xsk34eAbmXHMgsv/6QQX079O1dN13D+ub7YhVZJE1RaSyMRZFkWUAfwv/gJ/I75EH49S
mMFOU8YnYQXfHVXrkZOkvdWId5jjAP2PiCPPp0f/EBTumKu1ExEBdbbST+xGzYiyowrRd60x77UM
yJCERqL7tA10LQmM6ch4OaIB93uJJ+8C55DphJvQd/7Y9GNlne2XNM/PnWBUNyLMDpHBuxXhJVf+
2smmPcRfDrdh8c0oF6R7bTbbN+7IaemRI5wNHYSZR6tD9UxbuXSX2njnaS9aMO9E9gvncvpbLGpR
YkvH3Ygl3Ix2HLYuXcZdQI6SWCQUO2ZzEa2YPIFuDIZB5B6+2s+wHq18ho/hcdNUCjPLqqixbo85
nCowv/cTm2dJETByMvKkfdEZRY007j3LAxP5/o5VmcZfHsXw6dAKONpw4bAruI3mmqe3hP9FbyKt
Cfjf1WDselpXp2hrn+WNKbqDIebiya0ldlkqp2aYdmATzYFNBifUNQ76VElrk21jKvNH5vqX8qbl
kpx5hcXm4umrfr67y/kgdjgYLAEbO75brZ3h+toLdIdISd7jtEhMGAqNCIsR6P2tYk0Z6gLOsoUo
8PmbhoSSEYx67N6A061hbqpvo7d/oIDHyJY3f8NRkE9nCFg4ZG4WWhXdIguMljRBJSiB7JOZl2HL
NJj2KsNf5YIhLKW9TWMAwAVGfry3Z7yYmH31DsC0jG4Eg0ZLYbuYZD4x/6TkQyWj8K2NqRX7zdOB
IrcTllQHV9kBL49FjdoVmTllZz8yorUiii55o6AgBFjn16bnc/+y2MKQKwuk+R4u+eH7+XHxlEHk
n7hjoao0OCkcKgTPzgmFaOnBOdAr1EF7bEMwDT5LuRmsFI5jAy9wYMaVzn82//4WR5+wPhXuMxWj
N9tZ138aRgJic2bXdGwu4cMqkAe930wUyxEPOJHV+bNG6ZyfvbfeqEHqSQwAueFgXArh+fTUqxyk
DwNIcQRN7xL2QMFBN+h+4o1ZixofSwjrOctEpO124nhjcpoe5cKnWVv4vcz2Svt6ZHBP2UYMVNzh
IYo1dzA7Ot2skCeROpHrr6cN1YldiaScQ4yADHPKsoZwWaMsgIgZPKBuFknmW8aXTVmYDSgvduFO
r+M4WAEoCr27C5052T8l4QT00kZTUCYFnmXhfxt8R3iGJycTAqiWVk97nMwSHIjIah2YGE2l7cOm
DwLWVbFpDnKO+N04Fb3EdooHTf140GBLo8/ydsKvxcvd3beX4tB/YBo+Ky4xs3n6bZo0/tZ5i3hP
7Q0Ag+kyKc20Uu6cYVFpPUXRD+9Q5rG+tak1KfHzcpfLBC5nnIlMyupxNJXOCcOCq6OZXzhjgwBX
76VN01P1lkw146OGrWt+PthKHXwcyuauUV8LWo/oMOojGi+B85HGjConD8H3gqc0dJeXPop1knT5
luNJSoktVptMQkuiXahjUYJ7Q5Bmsb4cJ7+/BeUsfxThCDAgaUqqFNBGdzIqel1+fFa948WRygrw
r0fjzSl+LJgLPiMIBBgB3mNorb4Ckir19zKkBElfE/4n6yRDS3/sX1QdQKdeM2BHUOxbbKAFo3RS
nEtIxGmDr+rQKwn8OX11mLVuF4H+BGb1lEtT/3W5EHy7E1ZfyGsx1ZYDLI64Ipx2djqqab5u8TA5
6bOBLK3Qead9O5p4O6je3CoEXHOL31WSRQcx955Ls9sm6uqxvYdxtGmm/SqnODm/Sw93CQPr8Tw0
lc0vX5BQir9leer72T1ioe29Qoc5OOpALxykR9fig3hZTxWNH7tBCgKDHfktOTM6phMGbJJrzePH
03cgW2+D/a49lgqyvIru6kkTyEMcUHJwhJjbMzRsYRBjkZcGCp8Bhn1dH3xST+HwVVH7qxof03Ax
5ShQZL/BmGKNi54iEg3R2UDeZd1SuiALzpXzNTkBHQaSavRtW7WGI2m3t4O+G5ffP0NEWBgHKXt4
MzbdxF15CsU2CAXdlU2s9QCZzcJT4TxtQdN71Jdtbhoq9UpkUyy8njlwQLPEpAqreB1+klO/6yYj
kS23mtnN3l+8X/eb0u5CVaRorQ4Vw72ab1Gz/vgBBae74IX4yv31IZz/pF+3wWwd+e/A0ukYG1K9
YUqkNTn3+ZgaL2FiRZiZzjR7JJK4U0yBg4Ux1uCTVIWJSdEow8Gf7gzAEMkao+uT/fg3svqXipe6
n2Ia/C8BTIB4aigwXJZDIgAolQ8P3MS8Iswayl06oaX9HOrCzUk0uUQSGLoRt47BvfidOO8Thbu9
njsEpVeBOwMC8qyc1kY6myXxxaK8tT3lhFQUoVNrlSY8xkxyfHSroCLbffkhjuhA7fl2ovj2MmKp
hPJvuEa2KRYxVd5AZgI+MTZ0PdaZxyzfD/oaF1ZRb0Kj3ii1IQhRWLMNokOn88owRlktNRXUzRD0
oMuRt/zBPlZOvdx1jNx6Mrwk1GfaCS3TxIsI5EZnb7dDKeoXinpt9krr9KIV69D5IcdJ157UP3/+
6v7Mo7H+JxMCLnekp8IURLewvrWcjcgngezn1yFkr5lf5IpRrQGiok+hBN0OMs83YD51X+QdzIbF
ZkFPFR4NUaaEODqhqHr7W8XEirM4bMOfREYf6dpCVDyfFiPtoaxcOg2Uwhq68jo7MNfPOiwDXTNg
ZjWGjNWDgoXUdqD5mQJuLAEJCt10Csh2oyNvgH5xCMbqThDpmLmjpoUE1yzgnjnyu2c6/9TT5ndj
q1h5IT8eAkt0Brz1s9KMIBhTpEzFmqLtlT6F5CZIyh7XE6J1K/kJmcKVZgxs8HeQTPd5C8FtSdVI
yGpmUSeNRA1NGohocTvUOBzAB4mdKD4wyXi69VZQPkDb/9gj7iU0CbgFULUDUcHrk35TwKQgaixK
//0+ITCNAww7CK2G5S+zsZ6fRPhk1btXOt4h4m3fdypq3G40s8rnYjxEFqI+1Aby+IHcuDN2GYaZ
DKUA5DXlaTU4zjoYEwnFCqGHzm40HidalAOvDnSbgd9qpsVEVDww3hnbT5KJ07/2+ntJSteHEowK
FXXUd//pyMUSVd2OgD53VxpyD00o4zDDpJlYVjp2/JqjJM/kzHbYiSTKidOKYPVP2LRT8psEzllv
CFwlDTnsg7M4lQ2Hkx6aq0+pLegCrcKEYP8qxi7kJKETUzSo7x1SNNQ9Q15jMMm+00r/IXjWyxmM
bWjuph1Mg0AdRtDhJNhP/2bEzm/CnGxMeQkGy1ZigPk46qnpKOH6faW54umVTrXUl+0i9a5i1wPr
+x5zHg7exmrVbJl+6bWW3SHZ/rMoKs1gD9cTH/JyJvhLqJHHq81C8iZzC+TagBB5B5A5v0XCmbN7
Y39IxtFSoYV3nxmI+VVZLKzsVgx/kujgwED1BSqJw5BH/kzpbRHmamAuguppyNNKXw6GrjkT9RRk
qM6vjlynTr6MnkX8LHbq5xtoeixT3D8qIJjRus311Xl1CUHNnLQeuLOsxmb5beNNWrbuOkq/Y8p4
s7Ev8QTxrpXjDdtHWkwlreI43DBxqZ+qJlQzij79nFZS/o9NtyLvF8ciRYBpBSMc3Jp4b7Tsg6XW
fZFx0BbHO1LSbNixq/Zum1W6lJpPWAfkd6NATZ3Sn+ChqewwUoXplt8M5fKLlIPqja+MeNS/rotm
RODvC2erRVn+F0c10z+uHA/2SPj9s60agvMXyzYwKyrya3GACw211y7PhVANW0yQwDVoN3nFAzuu
LWOT+wYeXm3qUI2a/t3XimJyM4Xwza4wDAw5pjrDgwPNzOIGhOvXH/si2eos3pBYTbFjLJ+ZAa8Y
Yu098G3tDJTtT+foM7TtwfEuqKnLXNXKQmi01KXiBW0oTwk5C5eEfTgzjkNdKaPNRSJmsFA/PAKK
uwUVw6Gajhd1ixGmxLoxXPRUkte2OKSqYYjStGZzI3nAkgI+OpXSaPLLuIN5xQ99iT5r1L1FvquT
ppC4BTLrikZu7wauIcZzbmgmuCeQov8INdJetJbqqdFaP91nE8Zk71k2ZDPQlNhurb9pYMjk/M+0
k29ew6cBX6t+sCjTpyxU2271cbccXZNJtWJWOLuS11SvEc0AOahW0ipC9ymwL6Pa3wF7It73VqZT
aYPh/XkFTzu93lnLaf4s/JAGgLUNStuXJESnw6pBFVBYf/dTNaRMM5VFECk7mKr7lgEyJPkKIMUI
vDNU7vYB2wVyO+gXPSVsO2/X4NxaSMypRh8698MRI4lhzxd5TqbNdVMR+VE3VctRjJM23Xb5DwrU
SKb8A426dqKClX2ELyn99/WzaB+uwHI9vjrTnx5fles4N821+qj4VCxDfsRRFgS+MLac5PZft57r
fPB1jlN8yEhdIOXGhDj8PdVHp5fu0NxsbZmH9sNf+BFdKNvuplLgPYdoh5xP7Q/idiE9SBJS2Cwb
Aw5CRQvAbK+AaTxUZ0K2OYDhoLaX+K8O9fZZ7PNDu3zEkjdS6FZPEJNR6eyAgu3ULLc2UblcdZts
xcr0bAV1MdmCu3s72wF9GgJBgFL2N/nAfCyZ7HnL/1ljbFutYCp21YXDDKysUtICd2zoTACfB7MX
5IcwrjThRPQPwCodR3GxW2V6jDehsBeNg+Azg6lL4DMWESfCdloELZxrLGr7ppJRiiMspbwjMfx1
XjMtyZKYa7XmwibBtD3bIAb5UQNS0Qz+8qvxCtACZTrNz5VKLNVaSQ4McGyxPDhqDDHerK2ePE90
cebBjwPnm5mav0KBa6qG3LGnVkbr2IOsYJLklNqz6h1k7Dn8s2H03ajQs5IsXOOiQ0/az3cBOR/h
N18xNh0YfWUXN1aBewEgpWV4bD8+y2NVmFPbRrNKT9FuEYpKZDWgK1dz2aXpanMFRpzLohMEzfO9
kky+mufR1jAPIcWsQtXQxFJhTcAauiK4PznD8TaNYlofySumyDO2ohlolyjwG1hcbsROhjsBkRzw
a5/zzrIcSesGSW9QSHdgxcX2NK6sNkG56r9S6fGuHOUCLJ582EZjUnNPYloKsCSJrf0yGkJFtzuP
a7YVTbnhjfLr0jpHltBZFRfY4lizkMPNMov4UCwdESBBtEn/yrKdZTO4/ivh5vXDL6oDPFhvpgXX
FcMlaX7F87iO3rdwNvFCDGixvDIU/jMg1rM9G47WVD+eAuNleMoQCqIIARsqofBYQREITLFVXNzz
oIdy8vATucsbahKcSdM2avcyVLlAHX+Pv8WeG2VkaFDkW7ajLicWh6Gvpktef4/bN0Azg8kxUW3s
Z26/MllInIpMXGUm6qT7SK9xW6KRAsFH/Z8VxeVDrRlYauoJse0KfPamIZf+X4AkmP/63alaJuHI
EovLhA1Sys2+fc3qT69rB+qBCoqh1LXZQnCBXGCfY3mmHE9+egNEGxni2I8XJumhZrWBtmX07jev
7OCDODwRIK/nK30P7EGN2UzRJ9MT8ppgN05XUcb3b2ijahRI+zhlIPTDc1e0sQIU+uJ0gYIlEtcv
InFx354lp2nnOw6wmkU0sLS99E4fATQ1Rm/kEhbGMA8y8siX2xN64y5fHy8hAhOj3P1P2x5NXVha
vVZEjKM7ld2qjA6H61JC+hCl5DMpxkbmIFyeOzZOKD1DJ5gxcGxNoJ4zPor1KJQnTZ3s7T4h9Uy/
M52n7G9wR2cPIiACCPM3jSwSlwza4KjStNAOPGKTdy2JWg/ybpwHDfMVqcnJKvB4HLzqWFcYBt5k
pvu9Y+nbh77t7HDVwd9/e1vhKzF/SSgnJWDJHnx7GTTe47roCDZLWDcPOADWAwXGfWV0FmFQkejB
HPTtvstZjGJ7IOzvyLzgMOavofsvkZStKF8ufWYEDckNcnfmugH31tj2llKfwDWCDhZTupL8M/Qk
jFTWlE83GkgLSXwW6NRAZ2PWezAQvWK6w8454u0xiBtYOR6YKHrWGdZuA+4DOL9tGbvulXOi5mun
zN9KAfCxL9tiNf/iWFh26CEgjfKy/kTEtgBDQOYx/DZ9Nv6uf4B1AnzgsrSzhFniLmPnycWDufWW
rbNNp0oJ1kA5mSf2cQwP3ts6eN0/Cyczqawo3gZHJynMAUp6SQ3u3CERsOu4+XJ33JjfdGy0hU17
weiffVA0sehWepqd2ghGCJlEmAsioS9xKIYrahdXINTlsnEysB5hjS1FUut7a8qL6z8f0f5yhaPy
gDTQnj8Q9XXK8QmTtvOnDqVvua4KZPut6UJBLxDe3l0v7XM2ilfADeQDsjveTTy8KTSG8W6g33o7
Uga5nHNqHs/DFBEd/pWCi6rpkRBr2u99Yl6Tz0p7wxoMhy86M7HXjlvTZKw2Vjp2O2j2/XEpR0pE
3Grc01IP2ruA8v6AJsUNvxnYC0AjZgks8JZQ5oMP1/obQA3updiD7391ZdnaIinyphpYE0g7N1Yz
1EX7sSA2RXInQ9L2qhpmR1BNqlYoZzqCiPt9fSp7ie1Ysg+sgI4BDUS60lGuEgsfSpvDANpj8PhQ
I//30zXgHZRUu/+riKhX/u7DE/C+PTdrBBbgL0jhJBgv+3o+jvZkO1J0ErlNB2ki96bhgd9EnPFm
W3p1UglV1PAnW7f+LNoKUcD1ubMN23ei8I+s8G62o6fNlX3pSN0Rkvxyc5Vuae52G+xsFOKKLtAj
1amJk/mbX66hs2bKxii5wKGQbhfoVbc8LAC3hsuZ6iTFAiZh16hpUBT5ZszPk4ySofBe40XIhH4X
QPrIWyAmKJ2TXMiCFhZZ1/84K6L6z4WZfOCgsff/ybi5DakkGWAjGFwWgXUc74NikjKRYNLnL4M2
QBW413uuNnUw6Fvh1XRaDIZ+0ovTryv4vlpxowtTaXLUEgkqk8TQwtzbGeCUtVCp/SVOTUkuttVP
a3TrGBFnHLVF1OKyb8ZibL/MXv2SVe0K+/0erarX5MoyJrCqUu0PXwIvL35826tVxCMNZeMGu7XB
JewoFjNeRyFGZjgVugCpUjm+F7wE29ivup25Bq4mQdQeRkHWvu3OziqitW2TZonxDuYCsJioWs7L
J+e9CxEm1IM732gvBu5rDbOlWiXID4R+EC89Pk911bpmiU3lIKmThV7qYUpdyQQuE2V6faDFcfwm
ZRJ+r6ctZ3tnNPpF4T2M/ghsw4SzJgZv0kNW6qwCzKS7oIsljbW4Bbafzdj/ivcn/ia3pZcyVOsK
pQK0TK2wuSAn6KatCuLrKzM7pjPc4+jfxBXZ3xZ+Pn9jN8epL9Am5LHRS+oNooD4aKbD33ThSY6w
j4I1ToPDXcbY/kz+f2aHirl8QA8/5BmRxeJLpgseF+n3a3wKjWqUEAftQ29lFlmul0PSb0JN11W7
SR7X9N3p3N3qwJcILEem6m9AmTbmEso93UdBY/gU4t/Hoy24PqIUrqGcA1rJiL3CHb0zcefw4h14
J9FDKm4qf9p6m2fTdcb+0aV132refyJfp6srYXKC3C5ax2NjrfLVwL2QLtsPXEVAnHffezCmsXZl
fpP/UwhT71r3GRBHOIDDIhNlYGzFdTskv/MzGF7dd5Iol2vLhu6OUgigFVdoovXpHHkL606zZpJJ
ZtlZzpBud15T9l1Bx6QiKLs01kXIS/AK9roinJgQIMA1dlDaDeHZ8MmMsSKo6yTNzQD2D4srbxTy
40r41vFU4vSgNtfsjD88QQGVK5Uu2Oha60NfmNHzQov7O0/Ugj1FxVt2rHPHjN/XBguTnSu3SJQn
hccJyEL1d/KOdTDGRvrGi1iPCw72uZs827A+Bx86l4W/h6e5kWPIqU8ak6zcDFfv31Doc73IhoWl
VnoH1jZ0NwOO7nhTOanvYJmfweCIJ8QEjj+4gnFURVPGxb4ywFwuAbxpH/mk2gqW6qwjJh/maN/T
ZuS7Kl0wJ0epaBKisliZN2/Ujb+xoezfNeAKihFdJeNOYf7/r6DqLclK9uJjYWsNHM9ntC2LMTGx
rrKJe7IVrmWEMlYcFPIAByUjO+Flh17iOkLfMeECE5ZYfzfMZWX74be7+lZZDEL4eQbzcjk2RMAE
jQDqyJTWVlMQLa/01u11aHRGlk5O6BRmlbN5RvmOfOo77uaTb6N6adQCIhgLZAZY+CeQyBihf5KH
O/gQEwbKSjY6K2l7o9MU77I78PoSFSje0KCmrTDDImyOStYwRcmuieLOak/1aTw3r+awrvMZx4SA
3kwzKUzcrF6nTMIwGuY5mAFU1Z+uAwAEy8i/HL8vyUsZX9KEcIlaiYLyOhtfuVdwbv8r6aMvplOP
DYtJHUYRPfbpX4gKPmyNRLIjtYrexmJFfnpyuxCmtLkDUxQa5DM4IpyvbgTNUmTUQRYGc1jiiVPr
ei+hdQpla/QVEguu3oBNmYl5okCGON62VJYja/RcfRrFPZua6Lj+9Meg/VgggllyzhdO9XKIQNTI
nP2Oybk7FT8bmonYpz534Ndk9LqTXc4Tt43bzT3h6mJHDw/+KB2iZg1iTR6c0mqzaishrChl4Xg/
Q6FLejDLTtD5GSNCbhGvtP8RoHwX1xP3TQ7Dt6OSw7ir7AMHsOQorwWdKkhJK+qoenIMXNTCJ2kp
oYotKrgPvjL/lJrSGepXj0K5TzOKlM9YXzr0AWaKCbKxoX4xiz8mdnW1+yBq2AHa4+nxhVB8zgxF
HpLXb3VDa9lbZGlWwPUwAbwrszOrGw65zEcqcN99pd6uwEByMlmxMb82H+/z0HTA2z7xvPr1zFOz
O4Q+TFaqLqDmI1qBO5zId2K5NTj8V68G6a+o9AskeswROutGVojFu3aV+Fdd2K0hAwz0fS8QN85B
QevVgcK1FmwKThOzjMzfVzrMcX/tUicz/qZ9D+E9HBQgP2baawMsd1AyJ/q+tM67GkJdGouwWRsN
Si1mYhlMp9Ow3dn8YWfinXFGQPJSWpOcz+a8YluYtAh/MVjQZT3r1pnSmHxHKHoIbZiql6KCEOXM
xT2CtUdQYzo438y7MJeOALlhYt0jIJAfwu5HqNqM7ih83Nt55TUcAz7173YBgck+JRkHDioUdwqm
aTvyFsflutRHZCJSEdpCdpXQIB041dFckp/yNbRk1RqHLKU55bQvDRkPNIhibg1TJ5kF4FL/fCdZ
uVWNmfPO1tZFDIHYbG4z8cIHcXiYhLBpcihYNeLQxnMxH5yazgeYmqmK0i3g7dPXc13Dt4NnLgBd
fSdQMwX/Ict4XdO8IhQJpZ6Xvrd/sjn+A9Cb+HKp6/KEMgirKLAsR8kmHTgz7IX63nT6y9f112r3
Y4IYGnVmCn5GxcUrwn2vPskjaB+W17CDHHyxGvhCsQcKMPC0cDUJA6/BUZbO+JoMV+h0QnFTaGUf
VfM3X5/RT2Fvmjfxrl2j86YbeO/40422k5upBmGaf+bqooaysck0ku4OeQD5xhcKPBblB0iYYyYY
F7rcZVesG3QllafGbQvzfFOOY8JKw+ELIXLMajSsaPZp+P6Rjl0ZrOwqy7eB3yl/aQ0oLmpo+bXi
BLdN1p/7L/dtKlHJ3CxHlVGaCi3lNpLgN5163hCZbK4O7bFKpyS1k633RRsuMe+dekRWdd8g4x8F
JK0PPEpTL6SOJwc4C0IQA3tc/c6REgfO1oxqd4DPTCIeNYR89E7kCSv2Rnv0cKhOFLOOSYOW0O20
0TYihyyrUcBw90HUjvopwc0jQcCSjvjsl9QTVDomWrWZOHZ330sVo4XdxazyAl1OTEAxIKBvY37v
zoxzg9EOTBb+sUr1d7PmM7KxHAcuecvivdRgNeSAfsKqAyvZihbZ7DTNIUbPz0YUu9EhjUyoMv33
edRHFy9UP1RNkuv/AzI5923xVpQYiYFGQVRqdUCL+5KtgWwPMf96XuV2BIEH87SaEefQ+u2NQEy5
/l7/FdYZQh/xzXhaqzQIEbxKGH4EJGmvWbnjgpobD9SthoGHkH+1+cytB1Hxbt8h/hUjH2ZxyCra
9SJz7rm0M24cmMDi82utGRwJfJOhwTxLU4OVd9Br4xt4z9qSPTdGURWY/WaPi6nUAaG0vHFckL5O
f4Gz2jPtd9hXuf9iTQqWRnFWisb4brbVWlJ0dw/TGx8HNeZo3RNiQwL1Xly7juvnDkKys5tlwfFZ
gQqrLqYt78jTPb0MpOs+UYx+ePCxI0pmQw0XYnjvGGT+K0tBbkPl5t10n0IVqhl+NGTxuRrPCuRO
6YJbih28esmFLPDe2rqDzNBxDpYIIlNe4pXltPQoQUDxHrbgOnbY2lOcD5e9ojplabmi5so5DfZc
CSB0DnlpgLkgxvUXTuvExYmjAisOUXBjq82qDSrGbSefCmvZ/sisNp0Tg81oDSyZ1xg5NX/HQTso
83WDVy27DkEAAXqpYIjY9HS+Sm3LL9B9lMcgm31+lNz7zIqkNbFeRDC5fw/VXVRSspjVr67QGkxW
ClC/Q/6x1yMK3sunHB6BGa5yRADNFvAtBCTSTQp4hMWdaDNMXSZZNJ/e4Ljck5mZaLTfxB0VNfLt
zJ3i/hVU4+mDu99GIi09/qVedIMApbbJLImx3szDD5NyfuoZu3/cTuAiJp8AC+51QSWqlL+ICQW+
e/MZ9NGCIlBMVExfKhJU/zJWEa53eBQxt8JWhnaB0QVzGAomQmgGjnMaw9fDupI9EpfmowSChZQn
GzIfuvbtecN1yrUf15i76KEVoy/0n8ZVXLxnVS7GnAEU1uPr3T1rOkmnl19prgc1zMeXvAPpZI1u
J545CZQdR7M/eqgzdh7YYAf9+1mKMU2IS2ENJgYVgviKGYuhAeFoKQ9+5TooYOyXl23g/uJ9Jcx0
C/4xVsI40Y5kpQbqCd/o1MwrZC+2H5mkE0/N9lnoqPkDs6x9b/R5EyYYpf5B8qqTBip3QEHzKEb1
WMeeMs1Z9XdSljIKmNX+CnI631er8EELGkZ8Cplwgipet32k3Vs2iYrnVPub/leYWQsTUcczNeh9
3WOdFHanoOWa9NCvnCqYZJ3rU1u2Li/fTeV9uTIAO7ZEi793yF4baHiL6zw2gwz5MdTZwE5mz2U5
qvhmtrU0e6kf/3Cbo/DrG9zI1zynmy08hXZ5hRTsJf2BlGBWru2bD1Jxb8VulUgKOe+RcTs26r8M
vqwVePiGpOwSQNC2cG/j7WhDlmMI2q0zbaibCWCnYHt3Uxj4Ci0D+a4XYNbEs9d2F6pL1nCke4wY
N4vs0XzJVib0IKTs+FG/8v6C5kzZcftUGLekL+8NkvBWwzHEKkwer2rYFa0rG4X1K9QLSBdPQ7uA
4anfFEp0Vb4pu+ymA8YD4pu9N3kXAQt+bBlzSRY5QRF0Fz6hS4EMUMU/8HGSeshlid4xGWQ2hQ4i
SokgdlMxDYSF6vU+6XRI9RVFsLy6pNwkR5FGE4ncnG/MzkAQkCDi3KJUqJa8PAyXopTAGswf6aZx
KrguqT7Myf0eJ2Azoq1gdqHmVKlpU1FuOI/u5TtmLmplg2dcSberosV2VPf/VHSQvJJAm2Iv+Xr0
3JHUPrA3mv6uFBkDZiF4Dovm2F2PUqcryRDqK03jxR3G7JkLHjAiqg54BqrhT5ERIphOQhR8uw6K
jIn7vAILtlTyPHOzdwYXKnFtX1AUlp+sNjYIYO6XKEyw2aFlJkvTdc/UZPmT4O+Tbwu9Eky009im
Yb6FgcyjuxwFZgbGJHOFvYfITqmghRs2UlFqo9YmumUT9j9yJJgfZzwo9rpEYHgu4/Mn9cxUWshr
nl/sdPpvXB4YQGgT8fbEJUq7QKYpUyYVm9LvMJ5NuXjlmcSGNOdghyngN36HxLjR3++a9SWzYeX6
4KV2WzaO/e/Gk33x+PkMvHyMsJgxhXgdYapBMcFcmp1orwY3sx6B+vJCvkEWVzpcNmoqVhdVsDYV
o926vXFBH+y9pQeoeUiCugwn8Bv16XYGi4LSUDckNie8h6mk6yoUoL25KUQi2fs7QK2V4FoZ9dQH
m+lzhK0sHseFS5XSnQQDOsxSqRUq//YaSoP/nGJPoROqnLMXwbDoQMtFscTv4IuZdFBkFkdIhiMc
Z0dIEs5Flz5AoCGI1f/K2Wny58CLKQFvIIwu8OOrnhxwICeArMJfGBzPYurwEy03IwuM48nqX0Cw
4u2LkuLzYjHG01p1v+XJ92o/zSJbCTawOWsEEPzcjN+/nsayO4cFJgh3pGBCUuVQOV5Fc60QQeHG
vhlUYjuGli5hwMmztVbfpxEI+JxMDi8b7QnnOnNsrGy05M4mDzKEQQFEON+jrYY5rfEE3lBd7Uo0
EhbixlVK75PU4oTJOT9h2YYovf3edp+t3deS7riVbV4/yvDCSXdR1S2gmUslxeHieSKc9yVjt7t+
FPGe+XoXG2IwkS6buGkggdyEuBxMLW/wW6UY/cFOpYA+bg63G4EOBJEXrwqxDMezCozLeVNYNxPt
a1n54uRytD7b9T2nc8Tg+yHZuXb37N7QxRvfvxTzm1bYoglNnrzhPgKIqCoFZYgRzOp1c9WMSMTI
2yRG0sBME8rE4eJ37uboBb7PU0YGnYF/AsDgMPV10Lzo6p+8/NSLBxYA+ZY4qZ55L5n/vOxUJzxR
8uYMrXhxf16AXmfbRUpSJCyyJKuVNNlZs7JSKJfD1/+iscJDr8/87c4sG8Qj3PSHyFtgURxEchej
Wi8G4/9Jb0ABSke2c/rlUVzR50AAGhpCtN7eX4tLhnkq1JNdTVSMc4o2C+/fqAIhGFB6KMwXNmTk
AZKVHzLLz/YQomdpplTiSVibcmzyfff4ejrwx1bDmLPtQj28/ezu1QetCRt9USdeLuLuwhfeLvsz
erJjiQbGRXCVDbU9TxCEVjDnuSfNWpwXcU15q/0dd0bClTCB9GI90mCHfyXnxrUMlk2sNgTd9zZE
JZCGjXZPVkrE+YyQUxrC5nKdAnP7zSyTAQxKNxqWeXITLG+OFvb55nN3IpCVlV+4kdzvIDswhhIs
idBFZydfgh6cqcjO/HaKiW1qo6rnbpCDYpXzfI6QZTeyMqh9nC7qqq55ku5ax4/pMT0a5aXyFELB
1YPnDvNcO+75PzfjjnEG58/CXXYR0fCOynSdNv/N3c0xJ0YX/mLzfQdO8aHe6FLx/OoUL7tPbEOf
V3AUmqiWfWsXYa7kla2869neDE0nrYU+JMLijzFnFGF67LvFeGurV94O5Eu0/PNXwM5sjUcAHVrm
yJsZvBbXVuJl3H7yP5iBjaralE/BZN4JFYoR54fUdpKfnr9UWlBggbB3u5YwfvXq7RVRGfo9REA0
6TDYMdfYd0m+lLBfqpjFFQ1xmNhY9yUHYd6gcnSzFGBMYMDlAD6tbfEDmWQj3iEIHowZ52LKKauq
OnL3vrKGLcUulOJ0stlgr2/lgPetZXUEf/9o6hGvmBkXvW0vzCeeKedvBc4MvJP+fY2ELCdimV9k
Jyy8RvkqekKZV0o2e58iookx1XQqhws67CA7+v/aQ9sHVU/VSUUZjgeB4gvmTRo8fVlhX3LKiLKA
qtlXoCIS5nZCa5zVqxJ3F6+cILBkb84fhcd1liBJ8+HTpLV9j0w5a9I5QO4jgnSZxc/4hn7xy3FD
wBxmjcdqV3zrtymmH2wCCXKMox/6sDlYE/4hF1bjJG6lcqPXQi5qAxGO42lV6LVL5vJuakTUECYh
55Zms9tXI3oyItR2tbZN1zyq3CI5lruZDw/2tUXwKQez3CzZyVSYTb7kd0A8fZplkZxQ/om3XPo2
VQ6p7wXUdXKVVEAQ96xrZaTG76QgxW0uNLRj8lXDYw+fEsS+G1VQNq9XMs7bqYMY4Dw3WS+U2bKY
bwObtZUERvOeuKy3ay64AG4P2Ldt+AbHkKAP2vwezkoTMGzS9Li6JxIg/4ERP5n0plUUn96KHlCs
hjtOZvFVeDfwp02++tiKWn3hjXphpR1knxRtgEpyPoKmalGZRsvKXeNsXkWS3RiuDe2OUg8fkLlK
z2na3O7gM1EMTtjU4fA5FEuOjCiXNPOjudJV8rxDGeilularjbWXpONOEa7XQYg3PG2AE5RWeFgw
T+bk3OAbvqgblKVvR9P0nRtIxPGk5hyz7tzlPogGWlFG88HpOmLRTy+SM7ARgGqKxOvSD/4uLYTc
hmrcfgi0pYVgKamD6kpmeJUVd2S2PSO1BS/7ILg3OqqA9jOZ98LL5SJDeNFAcck2iBJDS57XQ7OB
0YannIWt5DEN+w2QWVTSLjJFkt6PDfbmrCsrap0hUyxwno63kM3d/oi3p5rgKHYDDErIhIrl6Z88
RVvAvJfgMnvV9iKvyMNLcS17MMH13HLuffqqbzDCREkbT/a3l+T8dSmhhllpRjZE0XOkRJqXA6NL
ukUCeksmHg+rBDiIoWtFprv5gXr7/x6lBmkv0IEkqXazhmy4bx1McW1gT+8MmmER4N+GQ+0RcuWL
7GqRGlfFAjJ+Cy63JRxeGMBbWD9Rh/X8ADMqOyXAZHUUGXi5sbmI/ucO/9fu6YtVDQFWjtTFSp82
TYd+ZSK9nFKwLNjCFRwAP96x96SFUHNubP/lQMFH8UBHd69fdAV3xzyzxTwCiRwzeUuZGzO3eeDu
FFw5cvUSzS/t957+Qwhh7qfEAXzTAjsBAmYELsnvHm1bDpX1XAf0uWnaIhEodunhlSBZ/am3k2iP
U+4sUB405ZOMSB3dHROZr4q6CnCHQ1fSXSKS3UWfXra5+Zlj9i2VE9TRaK1XrPU/Z4YRO9+qQnjr
KKcLBiItFn13i27eK5dzrDQ9nK9ZVZNIaG1efUq/KWEIep/soy7PqjE911RhNctN3K+R6OBI4WDd
PjE1nIA3RwRQTBL4URNli8TMrCiUCPyEYNsGVZYF+abL5m6CnO9ITYekbyiRqyocxDxsq3OquV3N
4xsAQ16QprlN2wmRsnIHEMph4Wr1gsf3Q7cPkwtSx5ZK3+l2Yl5dqE19QW1P7vhdfApQwTLTkygI
6ZFwskciyWrKBtQ52HmBe0W2RyNZM1EMnewzxeu/YkS0DRNfWNij0Zk8gVD13epRHnN3CHnP3RxY
1XUtXoxqoAIpwdw++toZ0h+gNAGdIHfZV161FF1qP7eN5Fko/U6K1Lho4ZT3MNuNES0M7lTExfag
Y6t34Wf3nfk8KZoTJ858ZJao7/P5qtwi5F4SE0rgBuobGYVSw6dUiZGa6EgC8jMGV1QM0vp1AaDs
1rJZGXX4s2f8ltcZcjra61bH1wJLG8gPqas9JetxQ4Ip0c9FzrlBYw6JvpfRs2TxbqhnVJFyltL9
joZ+yeuoJi71g6r8RGGYiTYLII/I5r6z7aIB4HGg4jVYlBza9TEhnOZFcnkKJdtW53MQv+cl/4nE
PImLO9iitwtGN0yZOcpzNEjKWJptsLMNozxVBFSvBkT8gREapt26fjhgXinIGoD2jayU2ydoyVLg
DB+LbJ5TiTFRHqVlPqHZdn/mNnM1YDPUCJeqjHCvr9oGFRmmVeQL/GAfLhbEQp3QPu5CgvzE078s
4m4hU9gA2HPJqHhDsfZ7EYXsaIkC3mRsV5xixkzImP3ecBEwiO2OkfYpHGyNjsZ9Et1EfgiM+4ux
bDDR9PAZtJ394X5OQytpf6wbVzjYsCa+VSEwQp2eV7qmNz4+Y8afKTcmtAq3CH8uinZK7RDS3ZWm
DdYOycv02+MgGSHwZWD36MBWXEW3KuulAQkVTubuj09tfGbZ+jWrykc2vyBNZroz4wSeAba+Kx+R
1XrBZvS33e2/oUE14ghMI9is+9oQbR5+eGJcHuSN6hfXP0hrC72MrOWcT7ctzwb+p9lKgJSr8NM6
rExvHXeCU9IApitvlRXKeWD3ZRfKdTGKFGLr4lLhwuq/P4rR7IL7myBooBTD7p3DR8kkgim1F/pW
JjNxLZwVNinTVHQTFXaVppIa3K2cP2n6fE/VP0GuBS10ti3nTJNlr/vpaB1torBA7KbpJRPzLpqF
f6BWlFVdME/vBaL5BcnphGOn9VyztWsiRjeddhLiGMQ/0jLppJhtdP84oKt7adS4BWmp10elPiBM
6lkUcyoJGYvhbi2q1TT+C0BCZJd3noy6OW5Q+3FpauzFcqu0mROw8j7v19kWfxMMSG6jtBKTlxfW
/SR0qjERSjvl2rhnsRtkspN+RP9DJFi+x5ic8xuwkVR6sasz8FrUuq/p6u4tgZULoZJ2MqzBiapS
dnLMMcU+Y5c97iXHWmroxs1hSQ6akiI+8J/Kzq9jUfPqbfD/UWRt66sL6Xt4ONQ4DVoCznYJW+nd
iMS/5CGaAu/gbu11bUdhSPNSBG0sTCiapUFIGXA8EDBIIH6y4QQ0Z68b/ylG9KyjDceWws7iHMxR
HFMFhtjSkImaWnlFyFRahyBAP/PlFZ3mPsWXAg28qxwNDShc+LvtT7e1ueizeRgbs5ZLR7a00D69
dHfjvVa8zMfiMub+yLoN9shWLY1Hccvr2ek3YxzIzVIbJZ+8QZHbx4QBatdPBbTfuRR/f8bhkafT
LuxZjwRX4RePujO6pFmrIzi9imMavlI3gUwLU+Jun72Lt5XAQ31kivNR+briDa08GFgVs5xTe+ry
7RY0GDwKmhvSKNf7jy/xRZoCbJ+5v0Lt+Zw2qP+vSznu9ODF+oBIxtB1zhF7H2MzBD8m4Q5PsDLR
10Et9wgOdd/6qVBX/lRakB7AaR968Aab0K8EKgWp2sBBNIqRC1pt/GVYKg3yqOtGMTp1SjzjdQZa
BWfYfEUNoLJyJdggtY2h2MvTFx83fj3TBqS4tBL/xmFdEASWdDgBT4xEBAvpTAhZjDA6vzYcPHzu
j33nRT7rxVO7jlGDQEVLQtNgCniCEOfat3XADotaLQvb0wQW4+SrhUwPQqqsidqqMcdr7sQ2q5hk
xjxq59y7oFj2gL8P9pqvsnI7n/5xDpaXKCINAt+1rFdfSKx5l+q6XzoFFwZZ+1dcJyCHaLEZ6K/e
s0Q05vrKF+R4ZzrCRz3iK19vde+AMhLp36VDdH8OMCta8BcYnlwIbGcFilwA9sApccZfm+t5YDaA
h9uIsP0fR+BHrbjfPLOqC8dL+5ZM3b2Kt0Chyv8cAouCklH1FQQ/vHqbY3nN5LqjwAx/7duPtn7b
/TkdskGcTLdc5gReCtZ2R1cKCkLlfDqER7m6UGW7SLrWzdFLstBwwNM4b2qnLV92CCo0rxuYxRPx
orOPOOMGF9vInBJtuvmxPqSDOwVhIlox9od6iaJYoBRmpeq7MsJsDJ6Dh8hsQVIeUiULThL6mVqy
RiS1KSsOUJnI4TIDVDHZ/LCvSqE9EqYYqPFq1EENAKuGrhlMx2cXlDDKkc6g/6Qu0OwvPdZaE0k0
Q1CF5DMMHYDDpD5/B5NUkJabXjBsx/NrJMHcpaYxonoUsjiWri92iD0NtoBlsq9EUd8XXuN3L6Nd
XjgdF0wXpMX3SdEZHJEDrtMLqd9ZTGw16RyPHa4KfNp6ilXppB8FbzCY35eWRDI3oaQU9knAANDV
8QiUJYKinJc+IuA0ENS8rWgrTPhDQdqeM87SAzIl5uygrPHfrcLGmrm8yspM6AAQ5e98mGApYneK
KS+cW+UOmsPrH33mW5PEMFGylw3bvfTw9kQqiPOA+y2zHkB3FDZh/OWQYzHCjHADVlFZBN5hXkCx
wD8iLN4CtDymjTFkGqfcmLmSDx3eD41RCSZTv4NcWpzKbwvAQs9hsepdjn/FTq+JGZSTtrAC/Cnq
lkFkoNvFGrqG0bKjljVGj92Uw6EOWHPHhNImTcyd47+8jq7iSpjjNa/CofUYKKtco1u+iWAHnQKe
oyvdut+MKkDZNm7LjfSNmRlQgbXBXFKdNJJqdObbC/7a3Gm5sq1aXc9ytU5b/Twskuv+519Uk2y8
PXQgtbxV4IxTfO++KkUHFj1VuF8ZbK3ReABGGUVJHLj0Zv/sgY5QnzALPXglyzQrLYr0SpIRw8Q/
ZB2YKMz9gIxF1eVX+SUxt7RJvA+Ob6cC8IwDeiQKGMiSZ4/Eo9j5mQtBDXh3LHpWlzmSD+p0M88O
6vgboidPaUWYLNbJ2qhk1wLiTPIqqV4SUFYs1sN1LLds3ijpGLHd/RBdYRH1sKXuVrPtqCPfbQBn
mtqXuIDZczp3FqG7e0Fkw4agEYmYfHyycYCadGGoRPtr2QVLeTWAaa4WP12GCKbYB4/wJq6THA3A
tqm+9W0fbXSk0PzDFDDNxpM+mVk/mF02hF081D+piw/GQf5Wh8PssZvaz2pxfX55walJHPMcj1kY
PrzfPAdsaesGtqvvTNaCLrHNEFUa0ISMtPAcgeO8u5dvAoAqnUms9nKBNuu++YiJFpV6VOk0DNko
GnxDwSdPpeC6czcu3sTgw3/i9klIbwd0zXAW7zvKNsxbOdPZKqJ1LFRLmF9BjMh4k5aEiqlGJR0+
hupTffD3Py+0FCs+xUSKpLxa6fvqCnP/cqgwnzOv9gk6lCjqywzcRRdyVOEFw6Ml0SQI8n9xeHK1
XjIJsshZGUeABx2aoh1FN2jTkcRvVF/Bvul66a5vYs+rCM/WlDqRugeo87GJA/Gye0iQ1ZMm+myQ
6AyEalpAK3LQa2DZ/llUY+mdONaqbqCHQWRwd3a0Rq+Tbl7qpkGRyGS/kBVHL6gErfjw/akUdSrG
AwdJITlMgr1xe5Pm7A2BHvhO0myBQHbuZv/WxuaztJPfN3QnQCmxOymjIJn/mksc1PKkOuElRg1j
y4wb4T7OBwu2GFDWdFy9+jrFjpetRmJ65Z4IyKUYiTP1S0ctleKC0CZslahck/XJBAJUJWXhUGVx
5eD9DQXEdR+3SyKIMEHkIX2gXCPx6pVGoGPokAZV/D28265xOo9dE15bKNdk6FS+BHrUMr+K+QcR
CKMVBTrWvlLiYqLKjnThH0qB5omNdqQZ2coOURYeKG1+iS+rcWkFn/st49x+Mq9hMRPCce63dOOK
ogQjaoWOfeS+hdJH7zqM1aBMNXuQM8qS+mZ+8AEk6qRMDnAlAoaf1BOkKE0GZAk1s88Yq4upMrPU
ovW2d5PqvrXglYFZaC5K3uUGJTZp3E5bNzZ+kOK5hlprgSRfYU0HijJaCtk2RhYRFJQeCoRyphUN
rOYqTS2T0UOygCFNscjq0OeEf/L7o/0iPXpR8lKCT5WP2ayd+zSLQy0PZXKy1Cta8IY82wbgPv+P
wKbdlBH7qJVETzPTart7qNK8irwOLP1fDqWsQgouGFyNIK2PbOQxMUb9aNJPi+gU/p06dGWeg1Zw
QP8UI1hmkeaS8qFQFhLKarzXn4OAMqvNU/De73CH7ukoBqpcFuFmqJgOCP6bQmwH1cTefXUebAqX
/5wfdUDlHdH7STS2xeSFCpPQfxQDzFALKd3wVj6Zuwnsq8Uw7sL/dJNYvw3tAeyl6J5P3DKE5XyN
Xxi0rYSuqcWR5+N9AuIrQfdb1QoPJ8qD5jfKokFebGJtFKGfbvq9EuUIkAdtRoT0TK1NvmHMjS9M
XHrshZ651npuhbcjj8/ahIjyuHDq8W5UlGF5cbWDTY1NxJVEAtODyDmsOytlFMNhjs5A/CRzmpRE
edsksCkFIH3JjmDyACy5suEYFM6zfSPF/qTqzzCcvgV098mwvl+Sf8NrmMb/+4wXCoWdzDRerhdO
aR/fL4gKUNtWlO6inNhPBCiDbtXW4a0+WnGQ4JBqmM2b0CyjxB4hRLjAunRL9XsXO4cQ+sPiB6Td
2dMWV+CEUkjq5weMqMGJj7TDbDBp8gMZlQyNgi8QIlUVfES9NZKbydrGDKPetkYxX2ddfFN8cLCC
3SWPHsOCRiaVoGS/mHZqfFucU6k1MZBzTvAUBYWiRukZbaNeCh2CGBWN2nqcLXWgdPx3N7ebCew0
bZOXSrYf70uwTc7kwGZSzzPqSXyEbNcNffSMAxR9anQ2ShwUBQPimefJSest+vtFygGbG7QKBkYY
hka0i9vLCa3evbpvgV0hdNzROVtTrmcBYE7DYA9sy8ytSjAHR66Tu88lzdl+nJPIBLgXsEEjpuyi
+OHu5vZk0XxDGcopXV3FyReffqWFdQSH+MtLWMuCp5lmomSnjAwAdALM3j6SKOoXtfFsULmKJnxl
mxmpwppa1JCgYibzURd9z7P8ikJ/ImURNEhVHcm1d3qpJxlX3CTBJ8ZVV5t+KKj18K8V+RP8SnCW
saJZZ0h4e/vCeqqdtekVwvwiZ7+YbMuAJM3rAnu0sKBtEnh2ctBlgYb/yMVCarM+uH03VDwCkiqC
Lu28bGsll/joSFvTGz3FI+hm5XnsCh9MoFrRYmUPYAoMnv10WBnwhXlmiKwzeGETCRpyma9xJJzI
6dFCRF/W7el+zqvvBQGMmMghahTgS+kFHu/uFphkLpLC+c8iNG7bIjgcupRic7DY3ilVi+fP9Id0
00AOs01q/w4o+wTP3IIoKk29+qLTLAZYL2Wppv5aQnu7RBYOLpmJuzOw91WB+sZCchUTkhBQZjQk
u/IdHqKipI1ZmrpozqJhGVCoHmU6cWEzmBT39nEvgqY5SUk8ddJNQeILOU42Zz1G4of9zPd8Awod
GStwgweR4FCiFoNAgEn/ps/BLNQ6fuAfJhpQ9wbZFnS9B6Qqz10t/tqlUrjtSK3k3GgF6c7qwDUt
wTWb5CP1Xrur9M6EKhJlttoBYMgkH7uiBkTcXhlglSAwwVhKJBAusk5yPm1JT3SRtsyuo9s4l8Bz
jNmky3zAmEG2S/r0u2+NBlXWPgb4sPBvurCr/VsofOHuv/z2TU8sqYHaP4Znao2wT5LqjDm/pe3u
D2D2N7u3um+3jz13W5e6oM7Nsl/pB253c1VsNeHSXtoXEEI+6KHBgaetOSgMjq5ABTyJt7J1SAvL
/hflTVLaVSh3iqxiUVTSfaWPWHnVstlKglL1Uuc5Yp5wQqCCHp9Ok8Mnre9rOHFW+U+XzSzb25xA
fQ1pnoF+WlcUhk6CHaoM6gSr2QVKbzgTCkl5PrFvl6kQwftty0SV1g5VKnujqhGJHA+ZJZApey7a
3ktDrOVy1lBsTVW+pzyj7TN3/fkLeNXJO9bQrqAOyNHQPiIhbCCP/cn70+aufPqZKm2u/aJ/DJqT
SwKlNdCksMl5bOhbGc9afc3HRDHIKgrJJ6HUEY1DMY5hs1Y4K6+4GiIVnaBaNccyCI3myg6moPBx
VSTiMjMElqGlRhdqjuXylrRABPxnYfiQMPKhCq8VyeIGcqUJdmTYJ5QLowE+gegl/huMoHVzdD1d
apJdOW0EwZ+plSh738KjnfZ5mDb4fRGyhIN06Fjdt2VIHQ3ol/klnzQlRTXl+yFYSgngWSwb/XQU
x4W9BeK/qjilW0rGidqaBZQhGEOIIC5haT+tvSYMvZ+828RKMd9VbCmShDQaagC8U6dBxEHpfOwa
IOZyAP9xp5K5xfMN3dHWW6bLdafFyrBVSaF7rSKDrBHM3aE1xvXbhfIKOSGBJg7soir8By2bwbin
1LQC2yt0aKX4+61hIJzymAmMA84HKsBogLPWAJIsXMv/RqHsT8T+phpLjgeqnA2MDZDmttXTeYRZ
vYpNTrTzhhWJ5lAyD5p1nd/IBVkSij77EvNpw3hDqUec4PjELA2cvlywAFLMdepe1sauQvvqoM3k
r9wvdLW2zxyt3fd3K2WiMxXf4ppf89jTvd/prDvAY0bJTmDh3Amhwi50fey1zzDgInYx/qXKIm7D
tskdFyPTMEfhJqpZsCjd3OFR2lMQ1zy9H/AVQVS8z45Zu4/DyYcVVnxeKl7Of/u+I9o5+TxTWgGI
OeQHIZFS9iRABdCTJBd610wRArIOiWe7Qxgecr+1hr/SmYsY73mPgFd3FuEdTndKhi6jQ3J/GXno
Gbo6v+JKrmihonGJuehN/jVq/5DduhRX/v1jApxjL2FEPsFKbCaNrurlXpRmvOaQoNv24bnzzIi4
sUntr+T9W3IsI22v5rK795egeLocq0W8INY0B3nIDfkpNcnwpW2vNgGkmiPmtCe4IzC/cdHJtDuv
6ryykwzJhClonSS+PLH73OK9feSfdQjifELGaBLYopOoSkAYFScOKoIwr3r/K/uqKKOK5j+cf9Ea
NyqeWDUI3FsbA+r4owMPVlnpgzRlRGMlhmH2GBQrQIReeuszBPmnkNZk4e/daND+7WotgsI4Fo/+
xEx7lL3TZJdP2TGi1CJkJnRBZywbRZEEdR9nVOIjuu5Z6SCT7O1aPLS/z2Y9hjA8mR5EJns8ewdy
oEvrNWLagQCmCoCt5+Doom4EkR71CDEgwH5whJhieMRrGWkTxlGZ7TebGGmkGoNrL3CuUU+Gcgr5
MZzcv9ia8aT/FFlHyhBG4CiLh2jP+3On9EfFfbJp1RN54kadatxBZfAJK7qVIrYPpzwkgLOjUBfW
M+HwRnjOk2eaiMSgtylT3vEQ0k3r485q6brMWLlfuAT6VuF2OnJotTDBqhsAiPOZc5T5WBksVptj
8Lchatnu1iit4sdyGC3h+cBPG+QwKg35LW3ozGpDzz4+xKtD6W612zlKySZKnxDJXqXPQGLi1NsX
/6I6S5oBIUuvaguHgazh5VnHErIJilbY+an5MvayzamNdI6MaVDbafPZ6jz4m7tXuZDDwCyqKuXS
ZFD0mdEVxG0pl3Zc+u1ImK8M/t0FlXEutkcPIwOCjsDOf4nnxATCIHNLuBLP1RI1G+/DQm0fGK+2
TVE6YkMlzxUIC1P9OyHxkJn4X/bwsU/uhJr+3lu7wfEaJDipTbgtehlXC0+gC2DVYYkbjOK8qk/4
k7YzvQbmiEG7D/vbWQ4cDkk7lBla6GPkrNUn1amqmhz3rAFzCOCUvlmk8sD/xpqXPPfzWs/cdTyZ
h9Z62d8qOFBUezow5RAzct/fD9yoBXawnUmcDhqpf6dL1UawYp4ic7BrGx1qKyh0WlcWh6KMPmQn
+6qWm2JpPb8quSJhRZ2D6iOGRIOLeoP9WvmszNcrCbmR+IVu+DODkamtJPgxelnLvOhEnF3M5V/T
93LddHaiYSZhJY7O0vk29EnjWq0H88kCp+PTZY/FNUxqUpxmgjrQfBx9C0AbTweq1PVsuqj054eI
GtC4bK+ZUXbideMyXkZQKyaUi8OQ+EM0HuP5YJQWeO65KcGM1t+J4jxuoKfpUZfXqx78YsTVd0fm
VoDtbO/irqq48/sxavwLj/V85UrUb5XCkwIysR11RhdZRIYDFxu4J5h9RQHSbahaOu5brulO0/Fv
c+pbA2FMQU9h93HhIMERfG53GuhZxZGj4yUy2xzqtuD0cui8TGYUFi71ejQg6UmgzkWUDzAU/0J4
xiYq4MKCrQNPEpdr/scxqX+uBU66zTjpVuP55O5oiSd1gJZqzmgK34putmM3+y8m61r+l4w7eH66
huedTXyfNvHrMGmMD9zFX9PnHNVJe5HNNdz27knUBg6qMXd5jdjBT+sCbphQLCfOyLzOkF40+Wrb
pNsHEuGPqdPm540I1BwJzG0EuoWwHQh9JdL2hV/BVjvLNRTYdXUabx5m1WeEcYsdjOWImgM2CzRP
xxrXEcjrw4Nsd8eierzhD5E4+SB2VxHt/N1St4KVQUJjREH1YarU7r2IExgYeuQwhGIPYXq9RuQE
u8i28ivsFPChDMVmpv4LJ9bPnIHU+0exMYxsMMX/x7W/00Fs7vldIBeix/REGai97IJsiixdFaug
d8KjfBd2yZbfDpcd11JCp4hsd5q9p0DSU27xsEYgrjP3cDj/KpGaOgVqaC5H0+mQMMMAi00byQNq
pOhMSd9qgZxZZaH2TAc6xz54Iq2p4v01jsOSxCGM8Ji4U5kXEXEjmiguNzyWpTJzNu0wcZ1IIufM
Fwd/tEb/2w9ytKRBPhKS9zgL1186kg9gSrnbd8jeGOfChwjGHBJVFTXxjUdomZT+dnlZxIEFhNgk
HTjQyJkXA/2zFYAVs8rASScWL3AUx+6tLzjIztvb/Vcyt4ZDzs+wFP9CYq1s7A6LTXSYzUZEGhsx
iYUag8IVWnybnXvnzl+L02FnipGqXp9VeWlmGQx4cL9B2cAiOwrCRY2w8HdE9HyRFHOQzq82Hyqz
SkizHVyFT6DhawuXaE0b7xBviKapYvtM3/YWVvCNTotlfgAdJNiADe+vhdXdgDr1GAKd1htfcLDD
LhSpcl1Isruyoo1FiNcSmjn2BNio8Ohss87MfLWfwjgg7HD2mu9dPuCEuHRJR41kubRzBRx3zey1
Mmr1cYYLG2c+68kKRqEFV1OKhclrc8qKV+WTpa7Bi/PY3jHQis+wajjSpC+3wQd8F/J73QKfQKI+
/4ipVmDN4xfeBQURY3nKWGn19ht1WqYeJroN9smhqPizbCOCwy8SgG3+DR7qTfqubWAdWXfofCSn
Ai1x+819mhEdSuSzy2FgxRV78cJejX93h7DIUGe8IVPwGXDF3KmeybSTaGZOt/myNxR4xk4q9Pvz
w8Hu0mL08BJefL1N6EHlhC23SBiajjfuAffQ7UnwpQjskPW8d3Cwwra/OzpFLUGANtpyJuPFQH3+
XPtQ0SwRq0GzNwVQj23/qnLFXbCHtXXwhHRP2NnSeemb1PQcx6RUHfVXkeiaWty4n31dlL4jkzXj
82TNIT1G829IM9jg7RC0OJTxhqcRSXv+VmLDR1o+j9ROExzMz+fDJqI0Pra1OmORPr/Y2FM7bqSp
e5iPgLgVixUdO2byMnYQ16Y20zT1IBX77U584Rlzljd+J3tzWqunj0tMJ32JUnvJ8PdemmnpzjVI
gFTSftSIC29KJnn0ZwWJPzmR0ZpKX5WVVJMsXHsTX3GlvMgEIxg1k69nkZThMUHH6gvTMusF0X0c
sn7U+xaGOdGr1zSUohApXkpVjBC8wn6HsiZV0w1QxVveR53I1Jkr4Z4mnqJeqSHG64se4H/X+maA
6XsHZ0hgqifPD706lMgvU7kcvv8FC5FVxheI7GoU9HIey61VhNecPsPfObr2xOzrRdT5SS63UJVE
p/g+dsXMW5hyhbX+tVicAXQoWzMwJuaFUCqpyASP/FYlhVyH5L++TmQ83SQLjV7rlFKyPDyjT+H0
Uli5iCnj/l3HVWamPLZcy3/api7zszpohv1tjCB7KD0LleDApJC+va7ZmhosO6QgWySWb0HmMMm0
WpQfqo4GiTtrZ+hHG0eJhKLQpPUjz3QLh16TXZp1bGhLSeRQUKOkZVnDBS8jdS0XfcW6kpESnSzj
Qnd/Yk+kD4N9Dja1RePUlL9NPldpWUjvRYQsZ391/qjSi/XAhJF7pIF0lfdE7E9cKD6qC8K7H1hg
bvIp1Y+M9uKGi0k3qjbKh7J8PiOYSoGev07jplLNlp5UrvWlhrC/esiDL54buojJHdXWkEUYoyvE
l/DA8Dr3PW8041bwGz7/cDvAp4g4FVowkXPQng94Zjq9hU9p9ydEwPRpiMP3eUV6cLjnXYUoGojJ
uRgci+OP+LrzOHIbRH8M3WLbMaoB3AX2J0Fp/+Pq2rdP6+v576di1aGFq+6td3yh5+Z1tz2F/pOL
bk2ZHiqYJF9iHhlfvm+EPLEL5ujAnuj+hwKoQJVbVPuNmxjGY2ZHDhDVu8Zf8JqKYpl0uz3q/hcX
/XW+S9z4TG2YWE+fc0i80z3A8cuwTXcwysDU607m/nhVhVa5Pe6gIhw9nPBEkTafe+fxi2PmLfC9
IlgRiHXIyD4NwuHv2CZGhIhNUFA4udDJK4iCRwoTyMXV74DNm9V8gLn5OPOnJU4OP98Dzu6/NN3z
6QjHvPST4X+/sUem0GoEjEtjnYAdWCjBsAbSU6gjp23lRJAuYOwjNDQDtI6JfP+oQ7N5u0c7kiE9
mnT9Ln0XBEKL3PEBFPhrz9HG0mBCMOIQfMBZ6Tc9RYVBb8EVLfHEV7eI7LyM6FJMq89zuofLjFJi
C36vizDvvphr1Xopdyi0wwrYI+I4VOOBQe1fGp+1ACuZismcmBscZqNVXt2S+98v0sIm3v85114+
tXdIsvKIfurLZuX0Jq3+ph+Ry62l8vtzsxA/S1zG0zRRAl7+LFaB5oMGbwQOe7cD02/9y8hmFrga
F7lDyyV5h4S0mO+SI4VitMYuS/TG0OF9qvwR8SE0WmKjqUG6DPWC3Ig+Do8eYaYcGILu2H9SaWEw
xHZEm9HY12f3tB48WSV0JGxvbiagtO6ksTleKRYcjGtaMuBO5JRTRVCegxwjrDOyyj9LlQXrhsAS
zdhMF1vml+ZikO6QOO0u2WnYOSaYHD6UbSPsr+3fRk+BlvzMU2KgCXSZthDBpH0ZiOMlKCHDpnUZ
UP210N2VFhLmS9hJQ0RpuXgPcQCQ+Je0tasAWBYNWbJs+g75TU8kdVtrg51iXcPfQLGTqKEaMAmD
8q9F0v41u/kiI7AVubZs9JKH+hVQkXsnq4D1s7oIckgNVZZCwdMe72dQrEEHZE27oEckStu+h5LR
akDURG8RvTlR1+0Zk879nawwdhAAre5chnva3cplVJ3WUc8M7V3s/k9CsQKMfg6Z+G9z1t44pEv9
nnqORFHQdE0tmUYRjbcOcB+NZmvHCO2B8P2wbAoL+xYS2Hh1R2q02lYd44AhcVzPVb3m6bWfgbeQ
wU2YgdQuSLlMqRtuctB9xbXEXicgZI9dbEnp+Pg/tmP76uqkZMd0SKzyNbire+SPCRf9Gekvpv2Y
kRG6wFQ2+ZQVma5Oc8HD00iyWiyGsU6NEMU5npfInQH8J75ol83Vkafx4BCXwgycM0KEgxRa5L7Z
Xjb7/Q987whL7MYbHpWzwk9ivvbuVmpt3MdZee76wtdET11fRvpFyftr3APIeaDj0EpvrWYsdiB0
2O+nFM4h2Dkced2119Wol8+bz5bc6U8/ilNQSm8G52vW05XLboQPSkCNLHQky+aVXxSLzK6gLCpX
8dWMiTav2mGOO1GMd7McHbsHBj8/kUD+mGFXN5S04hNHOSW3Ae2etygGo3ogNMI+ScymoXB1J/0a
p3xl3PmO8boRTivVgeaap0RBGS7rPrD9HPrQSjZZEuVHLpNN6QvgV02oaYj18wCUCSytVbzeLD0G
S5iy5YVuwLsh/jgwrTwp4dXhQqQpeXYKE/Q2I5+V3AlA74dIV/y7tMJ1v1iSj5gfBO/LZ1L/qNjc
pWVJ3UgWn8nP3xqIfKHhTHBSGzvwWHybBGT6z+W+6RFrLQNeEbG0Rz8BoTXxyT+1nYtXH9E3BWfl
C0EGoZ6EHwwUBGeJ+iJ1Xtv2VXy15GQGiiQSYc3UpnPzZvgWXsCuL81U7EPcM1tVUMx4GjWGGGF4
sRFSb2g3gz1zaTMqbLIpYcEL9LlV738Yo5pPb3kx6akTgr6c2l2Iad8auU8vb1ws+CmN0w66hXQX
De4vXukcZ6UdSDtfgZBDIcBzJTNIa9+fuD2jRYv8Tho+MqjFYzVHbJy8zGZjvnDm10GjoKJ5HNTJ
eTtnaLnftT1AOqd3XUOp9BRANR6Qg6laSN3cmpvsqABPg3BpyZJGlCtLbgDLPxw2TbwnWSChOYmC
0UeUSsD4WGgeC0iv+Rf2OIioaKNOLyKk6VJ3RLGCFbJg8Z2E24xA9f0CObr5tCoKjpVpRAiyBLSv
/MnFQOCXkEEF1tfmk3ALWTHpFW1DHRG1Fc20sTxv9GIGsSNl48BDCI5T/Jk9MUSKTf+v4A/85dRy
5QlssNtmm+6eqz1BJtS1HZtgi/hG1PffFZ+3CogAGIFIDP9bnMDweko01nrg58qY1yk+zCwBo9is
Q5IctXIC4TO4RvEA9090MxlRWtsb0yBjVO39N+2TiHaXkBaEgkkUZuPmJ5Ko+nExqkFhlrx74bqV
9IdPkxGVLpHhBq4h/zbopuOOsoPIGrRnLPDmcjch+AMR8ZRDaakKju6gvNrnwl34wQtruOmOvXT/
eZd5Ki0tE7oGe8OqrU4EWKYohzA7R7D/uyEOrtqdadysJCIQpOmIBKQtRoxmXpG2AJ009Ub4MDwY
uNLr4W3D36Z0uyU3JyJWPLaNHrttZle8JjK699tnRQwsDlZ5Uo5Gs0YCygaOn/SFZdlnT6JU04T2
RYyelTcZkvvek7K5ywrYHWDm2a+H0jUZZc5/VJ/8QcCVl5k1SGDGR6GKKfUSlEEDLtqDj3JGCAHo
qTBkIeht/mZd3JABMo1vFOr3LfV3aqzgx7qhOk24iOYyr9wMoilqj3Z351ei3tAHxOAvvA/4brz1
dlZNPz2dVSweJbqDyYKfZYf4C3xugW639OF0qUMxcQpEM/iiJZxjMNJ7QQt8SV8JNDozsS78Foei
QHn29jlQLGnyLE/rmCaHn7wuGOMD7ftBmF+2oi09dm30gafTBhShhKXwpZhhYPx4i7Dsa2OTUcHo
60a9kG+eWcqYROQeoh+RrAo2tJzL1Zzh4oH2D3QYQN0ircGYdssivFGMr1ttz7pkrcE/4IGePUTL
rHPBvmDU1lPvkAamVBszBQDOMx2Fwd758GYDiibFyyWyQWKu7Fbhva11GoAJSvtv+PVdoSpUInJo
uP2eO6t3ZQg2vqfVSbnHHVUEm9q5NJLovqr0w3M29bJtEiU5i0l4u3pPAugv6Ku50RQfoNwPURzj
CcJ2DgUOrNXTKU8Au1dQGjVnEAc81nYizyMf9WrNyYl0fphDZy6+X3XJqd5Jhd7sA6FpJ09dmM8F
iUBg9NYwzvSpstLBo6RwbUbNlLEV76MXOUN1MEPbvczzYutcuGd+HEKrMk/U0pGzm8Rt5u8rIuTJ
QYc4nef61XyltIp61sw8fdumogIzE54gVnCVq+y6kLeHyH7Tuk0wSavc8/I7ZPY7USscJX9JiDgr
7Lif+Axo69piVTSzmIrDCfJtbSMpZZJzTKSN7bAayISSgjs6YOszGb/SCOOzFNm1ff0a9Iz2WwKP
BJzwLoWlBAEbFrDqfJL8UUkopWpQqt6Ff9ELH1HoHCSrGubYYGLWHPALkeZ971iyY6+hWiyx1vZP
gv4WZFco+8jUaH+or4BT+EWoKsgFaznm9OOfEDb/L5zE8urShel7PvzO8PnF3dpl4yeRoJtgYvge
VJ1UOBgr2VCg4ImxqbH5DA6ioMedhPNptkXpNBiHvqwGDosG5k1seX8XKYmbe3r10bD115s5Hp/Q
nBdHOBwb2mAwTL3u5RzqaRAtaTq0vvZhYd1hN+ustRTAcdHvQBd5rMdPE2GvF9ZGDAKcx4/Gfuj/
90hiybtBUNDM0CwxUC5JSZ+DrHx7R6i5Wo2LvWt7fFOGUHFhtLX/9FNMhInUm+vhKF7uixGdAZBg
wNw+Tq8ZOMIDorBx+N34Fc0Ti0zDb6a0t0QN3NnTxgJC9oOX44CNTHSsuc0CnEP6PAs6+zbgqM4L
IRkJ0LUEyUfnXl7BixZ/ZtSrNvZWGfiSQdMGlHEIAKz0F+FXvoQXDMUr0cCc42JNKLyDQYPUbrcS
9J9UL4QPpPTi24EgD36J+gpxrJY3RTJ1UW9B9VIo31dZarYsXOcUD0H02D37p5AAwYIKR3mrzpio
ufsAR/bX0b3QhTq02Miw9unPMP5lc/IBUxIfpISk8Qg0yaygWnXuHMBQJHS5RMP2VwBzsiVn691E
KXYuGbInMoGdW4LC9l+FVesHK9Mdr9PgCq+rAF84wozGoyZBxrt0jAiGVbrP8wjyjZFl55uZgw0t
XRymRUUK46aC/MzK1myjrv67ymyI1uIWuhGDMMh6iPZi9KYBPwpLJpy9eqUHcAMwlOmGknFndoFh
rZELZfXyI7jawOquEYLIb9d5qCz9FHL9L5Xl4DGjMk5AE1Svtlj0a9ddHStLirVUMsAxMgZU7fp9
y3X4gridUBgVxjjvUZFD0uNajWky4mGCrgk4KO0ej+dlc4Z4IJJROJG2ejKFrJ5BLf2TsQZNYNmc
Bb5/RfRO01dVr88KqDZL6W4KmnqAASeEC2hqef+dVANsV2kAPn4lPGDw2y219oPGwdrEHhznD+ik
L0yzDQO6bG4k/TFl7ptXiEUbXKPnP1PbLuik+l+AH1Tt6mJYWBhCeVGB1XIjAy9ZZzCBJs/k3H6J
IwhhLhiGKewjfGqsIYq4v4hKdP40KWYkUfxp5SNrLqXR7mAkcxOAiKSJH6iEA3V8qnbYG3HC5Iss
8IpHUx3/OlDy5YIIpiCNnVswIYKOWtmJjzVYuIGW+M9hKNVlqDjJjlMoqEnWaHghvA/Etq0myvBd
/aZyOOjjgLl5b8f0srt81+KfSuBGoN1xkeiAbTOyfyFjuPd4qKJal960aCtkLCVVbWdkxaVLsJUQ
lxDb+x0AqqaTZCE5yJ/p0EPdPkpEZplhaRqVGXjvDR9LW0tfzsg05/lklSj+w8yqojBfn/jnvgco
DigjoG91aGTKofcA17tDWMzLauAgj3ZTKz6NQfBbJVa5G6Lt3kKIthC42i4mcY+kHsMgGJmWG9mc
kszAELYx2GTKUFlmLnAAOVxLEtclnOo8rnOCMCJ3tDDsmi5SLidICKCHKe4gI6BrMdiI8I0UXriI
fwXEq+5FiYhxWEOj28fdLYAbKFgfxi233zOYqVC1V7hVd+Xk+Y3tUqwdOXoZ9LaXbK2X697eO98Q
MAqGGizFtMuP3KAH9PJ9WKHJUfGg7E2Xr4rqd+Dtu/Z7EkFymeDROo9AE8BCFDQjF6tBX06Mn6hc
slMDBgROrEn2frMog+teHjsEEMwgH9oR8zp/BKOTAt2saQ9rBaSJT0dTvNQAnXzXSiJd73EPO4jt
BXPnpCb3jdbO+WcFn898ammujLxWg1hvQoe5SO007A5aLIMAGQ+ZzOTSuCmtC9YFuSeO+prheum6
uYk3qLFATs3meslXqrgwdNi/mQLKFHzOodWmcrxSdc9OOLdtoQ9CyWU5yv5hDVD1qKLN2e5dOJNK
znkW64JrAxH+3dAcRODLEg9JEvvyjzAgXlT4DQ3osiEzcJbq//sh6CTRTnZSTXBfsc5jGtTmm+Qq
tDEjAfAmE4OVO5Ehd7SBX17Bl7q4lqwL+f07/Q9dL41V7iQ0KK2wRXPccgKYFZirPD6pExaWVlnl
kGxUd/nHGC2UR/cxrnsdwsRWiirxZVhdF83qWqm1OJnja+e5yTIc8bvXw6XaL1gaVWNrclx5US6i
qlWqhqneQwu5eKsXs9q6tce+udT1IXvd6DqMISDN9FUEPOb1/M7Wcz6/gm4quyA7UNl+tZ4TJhVO
kyxJ4OK3vWJ5nFPnrnQYQhoaJaZXl7Hjwdj5fTtCiKCCOuz6yfJ9evnqRMEfj7wZhUd33y3bbJQs
PRfJ0BxBP+5jqRM8TFEh8hknzHn677VUDGfI8/74J61c0Bx1e7J5YtP+wPV+8J7TqPgPeHWydIIR
3ZEjQv7ywk3USa13f3EwZD5SibR0EdNWU2+DnjDy0d+MYlG5aeIFuUvEpM9hKMAsjEKRHjOBNpyf
HIY125KiToJYEsAiQ1eS3dgIU0EoSwcSJ7+G70XHIXPuudsjmbw648dYrqss8YAVLMSOFASdQHzH
9lAZKUs3DQCQY0J1OODiXIw/ROGwOHRgMYrm/Q4UkdXzFmsLuXYlvbLgd9w3yjDyRQegx/+l5oyl
RSCiyE+M56xpt0iWhoWPBbZ2WSiW4z7uMTylt/8z/1WkVVXCkSb9ogWp2QyyDmp97NUVmDnCXf5/
p6wikmAKLzEVWGHXTNAhn4lIK+Our85ynicDE8m6YmH07UJ4Lc2lDA/0fx5F1xo7YupG4wRhyK5V
lP6gMcW7VE6cdkq6SebZqJQawkY8jybwIX3KZpy9gdkp5+FM0ba6QPate+9QYm7R61Imh69jtohC
mdaYM6LG1adMPSVZarRXpcNFCtN3pC/sic9mApIdDbJFi5f/Yb4BFvgkqCV/zhPAcqzkhk5VufJf
tvpBwvf9ATsU0m47rp7QEYxM0yt2bBMKyiSrgfHLxgpyyrOQQY9/DLqVltml69BA0rDc/w+EY2F5
JXFBEmnnsbciJMB6LLQZYNa5X7ZTewHmf9xsY/fH/uVZBHTzQva/ZcA7ltl+cHLjamUGxCJ/ytY0
XF30wr/QRpriaXt6UbGmnMsUTHvACJnLx/zfG+w8S1i8EuwIYUJzg3hU4I+pEc62XbxQFE6YP7Qq
uYrWhSPlN58f0ks8nWnZpud243ovp/LCGLNMqLrt0YN28wbkmtYPRGoBqKw6My0db3Hab/wLR3fQ
GS00sPaBIuG+/Ru8+Z4ZYj3GjS2wLtbbuYa/hQtQ72jaKY7qWTYOBKlxOIG+9fiSpF8COwEA5HSb
JqOCIO/X52P+rsGh2PLFuVJkXWxLGtSvmKElRrQHTBlmfRCz9GGWZo4lW9CcBQfZWMUHUGf2ATlA
uBydy6xpfYqGIO4PSESf0Zx/+0Es2gQ/gNsX1+qbwchlwJi4vSWQzWeN99H+HOsTkgHOow3mJ+4p
ow5C02QK31CmwyAmrLGvOA5g5Vp9kHsjoKJWfsBma2qq2t64IogoXy9CnlswNG/e2ZgS+h5hRuHr
q1QFPHN0GYzlzUt+z13m05vXjSpUIlnLoxPyvlQbSExEDH4DeAur4QDjLnlR2T83FCkFoiyOgowI
kacRJOelldUawIqT0o7nXx1p7gUURNRuPJsbN0UGjKBJh2r1zpAsNOIUVDnGeUbEFUfvKmg0vc8l
DFIqAfc/BXmp69aLrGGnY0fz7m5q3OAdudZC/0jPRT4q3OG6pkhbJeBNyHx+Yh/CYQFSDz59wnTD
TWRtMNgwNBJiWK50j37XE8q2eaRDd6+4wYX00ThSwGwYbxE+/fdc5CsrLCzUoWhvxA2KADkets2o
apneJQZ/BhFWr3oKzGNkFiNqohCkCEETwp2+28umj2mWiR9vS3iX1XY/8nNU8PjtpzUA0ckw/l+J
01JoYICTAtFQOQdXy82ZfkWNnssY10DvblbXtWZnPss2lYsRtUDP8QGsh6hvysbaboHmckR5mJK0
FXsVwJr4BfRD4gByqPaxSqH0S+E5hZuXiidjpCsRWfW8gLS5QXQ6DgMy5LRRTsvGi1q+oTwMbThe
oqvQGaelwKPKmd5/Gl9sgZMyEyJyDkvLHn/EIYZQ2cv+e+Xrd4EZangkQySgmlVfv83johiu3d8H
H6gZz4FOPmNzmhVtKsjQ9mdRd2kgKdytcRK8kiNQOI+eoQZ8TG6QhWKjFd0IlwjG523Krx8E6zSn
AsxvErVVX47TNWHE6NodvBZr0bG0bs/s4V7bc1mB6Ki1lpx7hNRzY2oloabW9BhOLmPW7LsjYaK7
Uwrn4fXkQ7+HUyqj1hEl2gg/8cn/mX5DNr2QnX6JNqJX0VRxWIsKiKAJt+OXRZ2Wk2WCyxv3K/dg
hRjO2BFsmXtZU+SGSgFLRxmLeoBt6EBHI8+jTQNcCp87kfihqSz/7gztyPmY8PKinAiluQOtC6jc
aouJYvHFjGWWl92T+WEeBQht4sEFfdRkSyGJTU+b5OswPRZ05atcvk+QBV71fKu9EivMh4AR/Obv
eYlJ/r4xVe44GaDfNAzvbvc3FNSYdDo/f5Fz6CuvBLQFe7QHkkvWhRjhYNrgFfzBLPFiXATusrNI
c0fI6+S56/P3mD6yPrZFB1Puc7njoV/zeT2ZR9N6DyA4+9iN5IpSwCkbiNJc4kf1zgXZA12uA/vq
cOCj/sCGV7GI1/QVx5kXjv1F7MgIJOO2P7/lm0OG1YcksCaj5S2KffNO4fmQ9nZgtsnTNA4IBy3Q
r8o3a0+RnRF4IpbYEW1AK7fcwxD/Q9JJQhWH0o8g/CpSePJ3oZgGw0JfhPDURDlKRycTgUeam1hI
UTJKwe0OyFA9GaxZ2G1TkcYmIi4qMFXyynsKRw6WLjHuHW8PDo3SZlKTJ9V4qlCIgnZMLiiM8pyT
nWatkvFx69GXL6HfK/fWmkrRTV37k1md5oXKO5oSGn/GXmNUXmHOXadSLt79djONkc1GvSuSyOiR
nIBLxFB8wOCFitMaYQ3jC4aSC1zxzhUvnIMKALjzwK08yIpmW6JIvjB2o9E8SQtJbkeZNn4owafH
DsQHqaKd25Duf4Y6v09W+cIx4IjoD8JZ8JbciKxx6pinpqTNUV6SnqdkzysIesV+8Ba7cGSsxCVk
m0WmHGUfVfqoeunut38/SHFv2hBhBeO1/5pAxjtVQafSWtz7SdEJWPGCzpQ47o+39s22L+B2JZN8
l1j8AwIN/s+ImBUo0z/AyWxUPhJLIY9HMh6xyLFBIW9BGyYjfIkfSs9wlN/QO0PnFJR+Drt9XSTt
gy/QkkqHM6qj1w+HLxAdQb4p1b2K6Cr2w8Zh8yCLP8BWpd0eZLhbdZBqDCG8uI7aIZPUKysCk7eZ
seOTjj89eXs64RZVUka5jqwXTotFdF+FRKnAL6NkIxBUQSafN2hdv04rVFTTVyouD3O/W6SauSM7
MEgx3kWVozRHsq4ALqToaydfPtErNbubn9JugbICjZF1yttZH0n5h+pH8YetSW/geJ9mHgZrPUHn
twJynTxURwnWa73w2SDH795sIT2hi6u+l1hJcZuj3loePU5KbviBnSLJcywxU4x+g+82fmjxSUUs
UtjF/mJaZPW1ENi8Gqm1yzPdiu8EMstTWcko1BjJdh7D+KD1Qveo4QjSepWtNPOQHQaeJhl0Vmfd
Qct5Jyrit+yQWNBPTRBm7oUw6Ln41i44NhZrxToYkdUr4zULRKiNLGz21ngK+pkEIGHyIywFBL8J
I7xP7i6+7pzj9fpoD92hGYZ8/vVjxh5/shOzF9lS1X1Vdeev1hyT1tJqabKustIbRxlrM/5HcTvT
ggZYE14KrYM3eai4XUh4JWuS1jnaQ7rb5gcecXXFHWTtdZh8oJEw50jFnzCK6AXYXOnSJERaYndd
+8MJfYfdhtMSc/9ku1zdcWw8W4qiiyz1jTan+neqt9LwBj9HfSUq4x1aX+tzNTR+MgG0IjQwl29W
zi36DZF84vGrMgk2GZnWkgDgOCLv1LdTR4YInOaMVi+/dK8SfbXGwKObuibzMQWwnyZ/yqtyT+AM
CrwJGmsSztpjoLw8SVDphLftm5X6PLm3cwIZQ9pSXiPXv5W/cmiY7rDDhfTgqj429fxrUnZQlLg4
UbUvnATD2fI0cXdYlTrn1HlHYtpzcpUXJjPuwRRlpuLJ1ZIzELO0hdTPV5Fqw5XxyjZavoFabbiO
kVSlt3iK0LwC9aD2dky1vyxhV3PCWX8yBXt8C7vQze3/3Mbbg2ANFM6XPYl5sA/JBCiSgfQS8nTq
BUirWzIOFXN6x4R6xZkohlsaW2tKvvUpxe0omJ7nhw3EP/Six0zzHDFhd3Z04ccKw4G12nKe6yc0
5eHf/+9EI51cyC9rSn5oztvEcBvTEo2vnrEjaRHHw3gDdyxFAb729vEtWuY8JO2AZ3PnmjlaFgEx
YynoXEcrv0+oGO5nGcQu60nXOPSC5lH7K37R5spgjUc+UANfEV+7jQx/wtRxB6qwX6QIL3OnE6E3
VvIduAmBA4l+UBzjpfhOF29f39dkXVPGZ/9AdTBmcfkvYlAlCkV5f2h1gNcROI++0+Y4NEIA2B1h
T+4jUYlkfqlj1wUJAc6Da2iz6hsWKazDPrV5NVuz1GSKckfjzMwDVOEziIikBgRF/xSXzooFGNz6
GzCmvgdPDBuvPaA4rDmPNLGOO8UbJlmCR3f3wN27b7exok6/eaZyN24WxaCGScV8brXDeh514Up8
+aCAhk1+kO1rKqSom8AhigD8uTd3UTAa+xl+cgCz6lRszNmI07TLVD7jN5CPvUkDMSRSkutelsHn
zi/SZAK+OxIAaX5vrlhk7LuxZtBrAqm7WU+15OQW+uAeOyFP2cWKUwRG5Utl0IpOCUhcC59A9fek
/r7HW5Bcm1uFw7ypzRTzXGEut8aLy3kiYlVNQrfrrYSYxLpOTEtCkPBci3AzUFmeQKRKIVDwkiEn
PDfxa98E1cWyqBchT2xv9iuDWzp4SV709y5KVFd3Zlmeng23G6FFqfp5Cci60MyfO8m0+SH036am
9b6ezSTGOYD+IOpD92gduRlkSzwW2pJBSGTppxl5k58Lkkz0Ztlxti04Ky7KUaIcpQo3csdUWQC7
BVeu/7OC9veb0NtLZXK41dJayutqTg/G9CwTssiYC/M6BkyAzZUvg1x1kJZHur2xoM0+vnvVea3c
sos4uyEC5J/TPfc2mNHAtxxU0l2c/vzAI6N1lU++5V2PDeg0w/26mNrKOKkbaKNw9mcVXLbjnRC8
nz8UcffXGNiyfLkF7RfjwgixKwh3JDSoxSWuzvZgFG2U+XYuEptUa+eek+1BZnKztrh1Vs6jccYt
LhQroQPHAqEf47LJs1h3SY6i9/CFH6qqwBNCilg+qLh9GsSfyPtdGtIfy8f6ZZXIpTdQ9rOf9kxy
W/S4aoXyQ8kRRtF++2aQ+1pscpal5KrEVZH7qH5GyOsi/O0P9hCMHwWvGp8Q/7yu+k9wXZ8TcfGz
tE1p9q8CPR1CyQ9fHeVMSLNmJIf+xmkHf5bEWBpC+DQix9WqnwNFoM6+ecv692jLLYAUo7K3PvFr
33P6HdyVbsEGpQVZ6N5lcFhlHKnQ1bIauhfobW5/7+12Wax4+G+36yIuz0dHVK6dCc5QBTc8ZzBZ
VvXQxTNJZ8/A+u5UTKlvTxVMU0y2ar0+/6ishlbH8Sy0MdublL5H/cBajNMrX9yyi390xAvxh+/r
54/AxqsKjtZKceuGvFcLXiRSYnClKIftDiYCVOdy88xgdfPS6nL+ake40PyAr1IaRmFsLNYZN1pT
jtS/BrBw1Q2tmTuZKxoHDdg+bhuNhVCFHVzLwVwJnskM3BUlBcmQy77zpu+4NAz+ID6JCs3U5Xvx
NLiOxk0AIFaaTFYirBi1HGDNObVuMnGgzgQndCatdY5A7qHXe/fPd4aEF2fC4NGbMVFC8qPCtNzi
OfRPSJugzGSr7bp5g2ZV0s9jCOqxI3A6vJvemwrZ8E1PUg5aKgXeY0GtadRgKSbCL5bDCB413nkZ
2HvVW+nnwPIgJMuYv166z9h8rgW4RoxF8FT9Epyp4GOEYLx7G9gxm8xiEYkoCCvvmRnatFTTDKMw
uewokrfN+I1AwWKnM7b6qLNhwc3tjLAXED7mJa1Z8GK6kOV7on7PZ/XU1YHzvJHzKIjGlCLBcHxe
mun/mR770k2N1gVfGkr7kULqcQdPaUhpTiLJGfPjlVaYMGruDQayw8vw+ef3hOql9wJiepGu1l3Z
gSiZlCF5Zg7xsE8Y8KYJz03+PubmdwbIlClMPXnaD502qF3kbpBHL+x99hK6Kqj4g141V5zxkXCw
Wzu3PjCA73AGGYX6nAeNjscu4R3vFh0eWn/Bh4PV4i4lMIqbhEQrIYR8O3SuKJOcl1fegkCs8vDS
52kd6dQZHD4BfQLHLuAdSNQfCfQvmZo+tqQ14yzcCNiv80T/oSKGyrMiaXJK3hxlU/MsiuydSaHS
RiY2EeMG0oP21MKUzmKpo3akv6CLq3YIJVHUH2Kg1GDHeFV6yoqhs6js0mgjYtXqVBHlwk81OF5+
ASTGRgMTRI5XzUlhWIruYJ6g3HvS/i/8wa7nI2xCZ7J435JAwJZC0TELBwHkiw6dk+jzmkbG1TDJ
JGqXVlZxA/xDB7LN0yga3jDDOqpWD9v6E8gyojdwURrQdFUGnthW3Qj73Olpsxo5Hj6037wbG8H9
rAu/MOrONSxNWqR3qY3e9G7mDkJDtSixobuL0IWnzNqVa/Pl1Bubqq37R1x0/GIsQaUHdvJad+t8
6dVO3s7b/lGWJe/ZYAn1vp8OmUejF2AQVV/wJLh9NDeTFO7W8KR7eaDKvXT87u7HOdGOPdFgKMbY
9ANlP40WZQs4OU9Ck2PBECIbubH3cNBroxaKbTaXXfu7z81zeaaXx5rdxtW/QD5cJdqYwusQHEus
iOoX7BDFIra5o5045fcTedObeyhOhf08zjj2A1J5YoMe7k3k2v6moN7ZE7QWAt8bB9SDQWuZjLc4
5UZMgsV8i+VLauMB0AhzJnIifrdKF9OYry0zzooj1ZamxXOPzA/ru6o74tYnr3P8iOEp2OMjY+2s
g5IjnyN5vpLha4qVBweixkgA8m0iNWDVBzN1kSMfUY8mPOqwUgG6HcybhiHzdn7NPihgByt/LoWf
GkOHRdk4QhW09KItrlksFdbnhKhj6i7Nm0YOL0wM1VvzEqOCHhO2IWY0Q84vg3lew7HSzoJxX9SG
HXrANS/WNuXQOeAg3bzRTIBxrRDu8+PP1++L/fBl+4H4cxDHJMGxEL34t0/eDNIquDhYjwDC0Uqt
SNPsEHQezm8jLekHkOzqfM6ECNziwKh05gCYZAkhjooqjUzP2E0e8CT9M+/B379Mo/87F5kPaWOR
hBeYQ8kzq3rG9wOtQ0bthg6wfUfXYk1nXygCnW/mfJwrHqn8LHpZy0lB4tGGQkwS7/zQ0OlqTdB3
meKYqFjKPPPBunx1l7r7MhEvmlBNWhTHH1diNbzhI1hta6/1ZsNIdmRsYWHuT9EKgVayy6q1i/e3
vZO5aXNd7Axs966mHFJdzk6qxYhH0gJXysKNuILNdPxJHVYORJ1xeuOMdTD/gbeC4xPHks8Npm0y
dd5+tdviJafi3vqmOHKrWNXA0IAEOkZFRs4gu3vrpXZXB7pWLIC53CW2hv6oQ2Vr93gezeQL0Pzn
Pv/UsO1orow6EkQ7QRqxfQrUZ0vx+L5N4WzYPrlm1KtZGmT2jjSDjsZapP+Q56vjM/GJH7wRO6RO
k0AEORBgxWNhONCo51vB7XG59CrRGe7JNDQrAZdVj9TknsuqOzCPOtqyEgHXuCgqWlmYzWZ2xVBx
nZyfAJbPaDsfcEdsR3c7VhHu7y8S8tXY/Au6ntI2Nvp31LqB1mHJJRdbJjnu/fTpWIl5hI0eyzsw
u9sxeSm6ZHod7+DhxeE6AoQa3Og+wZigns2v6l489Ttd7iqep+yR6bTSjGOHY4mppl1MnoCAB4xW
iMi3lgik8V2s1YXuGlq233BlCWu1fghDd9+FJFyg34BAcWT5Dc9B2TNgVITLhrA8PvvKJRm9i65Y
ItjauTVdCTB5Z5RG7m5B9YVpWOeBnmy+Fz/SdybIJ7cEC1jVM8CYI9Aqb168Iibgp8WYclHk2/Fa
uF5nx8yh9QnLy21qQH9BhSwlu+W+/ZwiuvuAa/vQoxAnWQiFQ4OlKsCedDAq/+Ry7vATUEiAf78S
iM+cue4JxfZXzk6k60JXar/OachJmeVw3Hyf1jJ3A5LQ0Ls4FGTJbzdMonxojYyCw7HpYJzLYgID
6uFqUl0Qxu+aIR4Fq7RlCHOoHzIBtmJzGjWmEcev+Rg4Aj25lexdqREneLGs7C4II34ZRbmdNmjU
KCIo5RwK+GHnAXNSGkLTPjDal2303z0LNQsDi4dk9rebDSevWg6jSK5Dhzx0aAQDcfVQlJVP1DNH
q6KhNYbEffTswhLr5uekzw6r6cO2HCaj5LhxJt/uWjLhgnCmfKvPiybdX0IebsKBvkB48ui1STAI
euTZc57RghB9ibXwtu71aSbPTH9HNZzuor1odzYcJwGOuTdtPJJDErC4lovc29SKYrQ6JMnz13u1
KuQFGUWc1KSGLIV1TN2WdittMLHyK7GJPI9zIjlVmqJ41nLn+3m9BPkAn0y2g9FvqwLIxQWbEsak
wyXq4Ka6lNor64/TJUg23Szhk4KryowEvqYmsqIULHFGK/eTYaykzIuPfc6pWtKHWhAI9MMfWGQm
eDqtrOVL3so3HZ/qSTGbMCBBBbDF+u/6GrBg2gXj8V98FcEaVbRSfKlOBpmn0JyNjmbT1di0bHWT
U/X5iRAzVfyjTbtmxtpWeySYyAxdXyrXNkw0ntXdpCgGgfnL7ZD5JVKUuuh88TYHC8wfs7PRvvqp
lshcV+VI2Qj+gyBfRjH70aKDSEs5PVWq3yjgkykW0Dny1dwnZ9Z24qxelipXOzfUJmnJcfEAM7p/
5gFMCYJfOhzAlMN5Fgd2Yw1SNzIS0skMWhhnaOtDpQ8VWSsc8JSXfpoxk//Lw6LLZYDyw6IKpbm1
7OAn94nTboPAUvp1Mbmi2kexCGAyLDY5tvrFvBAjr1OGjWgH8G7LOT1C07I1o/dIRoetsvSW/PuO
hZJ/ofASMuv8X9y1yRyFNYzYKm9PIv/a0TslklWoDj9JElf4C0Vj5tQWTnqihsqf1lr39KkSDbEU
NwtjibOyN3q2DUyn6mnWfLvDFNs1lusH306tZsu9i8qEB+fh6AxmTAVpereEAcPpNX59rJ39MBVY
pthiQMu7YurM6cIcwzZTZFXgsq4HdkJWmS1tFLNLw2JUF/5dwn27gR8Wjfan1ZR9C6NS+k7zz0qm
JHeLh0a16ryUCShvL2ZTuPYJObeARgYI4OflLsKglqgT0fgMQaA4dlHbf/YiWlYf+dGkf/MYs6py
LrlgdzSDbN93+HlfzsJqeQl4tyMgRxz4N4B6Fin9Ev3yCEow8RWg0eTEe46laSAOsiQIfGDYAydw
S5cLpKXZyhJ/Bi0r0SJ1X9i5LdwAZHItQcm3Jkx/J5gTi7sqOcFNY0R79ou1Ez6GxRY7AXAMKLRL
TY17K4QiLLH2WnhHkdqpBB0iC5DyN9sZ2Ft7nLGODjae7xZ6dIMFvKuMhDDOXd7jzimdb29r7YXl
YmKzX8bZbmHkV9YoQzHJEnEsolSo7CWowophT4ov89RitmennELE/K3Uiw0w7crGgwe2dkOvJPzE
TuAV8zgzJHRF6oKb6MdPNBjLbTJuhMQ0du/0pq3a97AS2niDMVELRM4T9aZfqJFD96NqIlhCl3V+
MCZmg3XIPUtMBb2PTqZOlZ55pjEX9QZRaKrtcDoYrCd1jNQDMBfAUWeJk755Y1yXG3vcPVpX8hB8
rTmuf+beKKgfOyc7FryPNqRBWhGN7uiqJqurzU2R6O5H7+jZarB9CesGmu/9jQe9N/etBUj2Mw91
7GvJikyOa2rIt81NdTUq13igsoFNHSF+goatqgIOyWkXPh4fAcasBo+Je6jvaun6qPg/xrMmO0LB
BJ9PYhBhfpYskcUYQbVOnIuz1k8QhveOtPpkkr9T3VNU7+SgW4OAr+1VTA39r3Vhq5I63Md+LmXE
44+BB57uT9EPeP3UF/J0mXwhOW/a1l6rHy9Bk5wC3d6crobIMTZr02hfytH680DCeVnXAOOVDuLt
wnvz2bZHto+Mj73BlJ+bfdS1MpFjkbQBcV5vRKw6kVPrZ7qUsU23BZFqZ01T3AUfdFOksq1Nza8O
PzNk9zbte0kx0eFCAtZjRQ7WyEOfuEaSdUeVCHZevH8J0R/ETdLVVcpgZcXl+PSSYuJ2DYLL3BNe
u8jmgvEDW1CxVaw8MZhN3W5P/Bb24edqSCeghcAqLIdTwjpoXTtahh4CVMdH3E+VxbhfE2d16619
Yr2LwiRFpV+4PQ09d1PtgeN6+nOCaqEHun7cT2liJPMh03I6UQ4GWaUrfRjLUzQpsWE3zr6ijt2e
Mr1GA0GN6fBSCd+TtZkg3HP1/4l3+OIiq4aGg2cZgeAY0Phcof+8SrwQ9xOjWSn4/sLu+rmDVTXv
nHzNrcQ55phAU3QXYWZWwTcAzLmmFxigMxFkPbjSEj4o94SMyw4cX9+GklKWMy3045xtFRkS4KVT
j0bg4XwGbBc9RZx1LnyFZ5Q6bCkWVbcR522bpT8j1RXpfIEN+f5ix5hfRfhq4SBntcoVBK0qR2Pi
Uw9fd/9WrEDn0tiGXLKLZZvOTxRzgYgCs7jdP+invLkHxjyycPS5NLfy+X1GpHyNXXHvXQwnbtVo
cA/jCPW4OnPcc7UYin0Xo4lWGbFu5tLARjMqwWgN/+KxKGeCMd3HIcsJRzjrUAC7agzKfla2EbgV
to3yimVCO3oCI/MQfWWrSOAYQZzWZAZ0x21zv9S4ygVC6YTOwwSFfeXGzKOoZ06MbqxskyQVfuMp
Dbb1/LODN5dq0LebVrgSDCxr5QspP2R1PDgZbDNhzDspN0hkqbugjKpkgFE00Xif6G/8UdQmYR/h
nP86UAx2L6/A+2g+PnD8SpTDJnsqmiwr4O99nTWRH+hgqxexB5ehl1VU0KV2O7luH3I60LHLhLuL
dC083UEAHsaeWBhOEFq4y1nOqH8dyePsydVHzLENHzTwxwQyC6nwJLihP3h26wWAOFlaPRtCjSpc
i3eXbctNAVUFxwO2QJe6xx3h5qIrKNfbBSoMcVQgl6hBFbuSHxrH6OlTJhaYj9Wy9747u/i46MWX
/uTOJoxsvZWLYCNs20v4DAFQbz1TJLMMdryVvtyoGdR6mKT59MAQ61XryZFBwTZo9APyfp0UbWuW
gibFeag1x3ZVMVxEAwOCR7XY47pm6pOvsdktfCJVdZB8MLnYclp+Rs5Jx7I/u33T6pcMCnYkcC+j
D3amVQWIIgla5QDO13u2fJ893Ng2N78rrabJMyr22hBF5OfukIRhovWig5VWp6S7uV2b5Vhhg4PI
vluhycIr7jJp9NiOD3KQnLNqIIInFQoC2R+Jh11mg/NMdyCc77IntsOw8beWYV6zy10VPikD/ova
AJGGDl7eAOSTu9+2nqEAGOK0hcTTYV1WI8iwXOz2Amj2O06ZvxxnMwoEs7RUWmLdSoFa8jOzWLfw
AUN6i26z/uNugG673pumpW/aH9fJlzDcb7mnCwL3yUum897kf9U6co9RdfgfGgAiEtsS6H6UUrYX
Z7OPSU+06J7/CVXLx6sY/S8b48rNah2vF47MqY/KfHO+Kdi8pKEMgrsYj8QEID4fZLo/9mKesyqF
SDq113dgmKDwQoWyAKAjb9pWsfNGEGS7130t5uDYz8VwOnS9oSTXb3CMqEWUHUI/N7/e35pmzNB+
cB0fEpGZ34Jbk4D2+guzvS+FjDs6U94pVAlt4rcGNfxNVm2JCNa32BSefXRkfpKzgixkQ2kRS/77
Au5h6F/hzR0S4Rmi/frum5KZm1gAMH/fji39Pd3xPjJpWKH4OUaIK5L6hvAR3gju39B8yFMUfQML
pKy7CiiwhqB3ZYKGS1sQW8Se8AOkGGz8fjPefdIynjlT2j1LHfJS+upiRuJVTDqZUCp9TeRtGgpX
aOUbbbSt2tNwh+iD/wui7fftujB3+eCTiA49jubdV5SK6HR2Wf/UhFZH3+lpXcT7c3Wg4S2y3zZo
DSTJjtTp/wgeQYVUrnu80oF9lOVGOHMQ106uDeilZpRfxLp4M/8ZKoDx0hHf/ATaDk5jAXUN2K9a
S6CJEidla6QNlpGYWIkvPFwP6rfLioQxyx9Gf/F24OzLM+MXGNQYqyA0PoGRywFjX9UqY8RCHDwW
fZr6EZj+VVqRotvK3XvHIM/B0BZP7qSX8QZoBAqpJkZZBYpDlrCnXHSFYC8E5fy2e3cjmZUlC/64
GpkIeydDW5JOvuDXKkZ5UniKz7YDDJToe+v3Bv/EVvc9eaOLFG44kI7ete1yKK6RwhQ54a/NomXL
ADT/fNQycZEqd1v4XR+j93nBzxvINGZlFUNFxz54vT+f7vShpzddsPECDaARXYpsnEbQmC24b6o2
b1Mls2v7fK34xaKzBaMwNcKO/m1gWd3t2xebyogJTbYF0XRQ+uGrmCohgGmsBJSy/qQVTzD3PwzT
pmFYAY+E/AD2r44BW67gi75wQ4uObYfZDY9eud21XFg5JM4UiiO90GP7u2dC6PClz6ICrDXYXR4C
AEhzF34nuSm5V8GUI/PxDz/J1FzEzxoPbpBmEvN1+XidxhuO01VnulyFSXUPhpCLGyKvELBoY6Bb
mKoesC3AphSQMft7NzyBPnTSNdMo/gthoU/KDsZWn6NMvkZMdEMlI0v7bdTXY/yV5WBdwlovYZ9p
LKa0bHfo1oH64gBaMYx6HTRpw2P1ctwd9FXHZap9pyULL28+EPVmtPcFt9O5AMtvayw/ncTftLdp
hbPQl7ED33cXBBSwC8SCngoEn73R8n22w7qN0oHhe9QQ4p/IspcTPmQOITFK09Yhl0xfjVUeAXQ6
24qoGQydiEuk/2MyVj41fXnss2DvIHrn3/ZJsQ1RlMn++dINtPYozMmpcoVkD6OtoDrR4APBk9eY
U0n7XIKg9m3kuYG3bnCU2x937txZ92XtfAq9TGZcSRrzS0tis2aqkzrIFV3/Km+pgLZgkmEwl1v0
wOuBy5gb+25WgMflPvzTn/OW6VFrktzp7aj+gtBu/ihKJwqGoWP7DmbU6Mg9z8jmAdHmpwPXXVan
QYgQaxb1LCoq7iYUcVg0XQOZrxRyVL64MjesnMvxdPxjsNy/OjkAbkm8ORz66nKeL8tsiGWpGepK
lguJBHPUqf/xhiPBeseUJxzk4tWx9mHS+SVzVeZmg9h16drUUtmD0muPruVNrVAxDQ2yGR+xCFRl
RkcCrKZtXOUtqX+nFkxP2ZyqIlgDlhmLWtx7iUTp8avn9H7qKZHkr6+CqBA7BFgOzDkiwmyfsJO2
4qoM9+hFlNKEhK02KJOWTMJBu2U6a/bvV9+hjB/YFJRJO7lb7rnCLIcyXy97x4DDPC0bth4ywxH/
LvRrkDK8HJivwSJz+NrwYzRbyM9fpwjhIvMvSBiQmHr7AosOHIeni0nMHMtei5xt2kX0gi1AcReG
dqLwl5e+kz77WQ9w7gEkUDLv/dkSyO8w9HGQsf9BInbWi9E2Ol8HRnp6w11bZbGhenUc+6Ipcvce
YaQZl9E+aHVly12PyPWjo8ML1t6NLq2w6+WUnvKnT+pnyACMICZ0rd1IGSElTsBvqQEaIlXPEbo5
y5YOELLVnXVGp9qVPMH+bIllrTSA3h9JvPPztqquyqcNsF+hR9Qi7Yi+mAgZ3aOsJJGZeNvZOqO8
efqqCmn/Mjg2lZx8Cdq/rNWllmcv1uLpNWIXGw2N0NXKlzr/OT+eBgirz9JS6qhyXh1rPrS30yf2
K4JKbbNAmEbSyKF+nY64IVdhtf3H3fZmQ1ym+CdGrBqbia1/6/uNMbG+HGIAFDBMKDuf7/ogN+GB
5WlfYb3wVB0phJowMFYeSw2+xdy9qgB53bDu31kuU7NA9cqKnE94nOHpZ8S+xWuTv/DZRc/kuIse
5xv7cAbZkLnmrTh11T8aEjyGMV12IuyBFF5GbaLjfEBnQGLIHwSIL+lMTmazq5EQDNtAFL9g3c9S
8KJpUCx1O0nCQ+kBCcNALsLZEwCpeGZsfj0SekmRePpIKYe6W93HXDu3Cq9wvnVGTWEvf+aL8JdF
LJUm9D5PQUSNX/+nAER0rM0wwo/FrM3EUi/7cKQrLZ0BKuoSPbeH1D7fUStoz+ahRDPgIcECd/+O
K9bjZQX8RLjIiTcL53/koKzIFaUSgNb7TVjEVDy+ghYA1kgxFlQNEiPG6JOP8sA6qF/GwHffOc+0
S+NRPfkaXydfR2dDgLiO3sr0Xd4rt0gSKZ/o23fiKb+gA7ygQZzxmeuP0Kwib9ThJx6AqXdTf70r
tK3OUc6WhaXtnzdo3PHI6l9ieVVvp5zS8Nal1ZX08yaGnqxHSSagyZCR7kerSdJIvJj8m5s+UQG8
wcIhRzVbKhQejMT2s6WWzoFMDqotGVMP0nSlNNW339K2rx7TZbfNBUU6WaoDNx2nxRZW9SglyR5Q
xSfgimoqQ+o6Vi16ftEWkxWWYSAw3EpoRtpBz4E9wmv7yVEc8tq7qDeHmKgH3LO2Z6l3xorN47AX
REbqaFEOFJRxRnZPYBmeq90cJsuWjAZawLtkDYL94MenWztbcAjyAq6S/4w8HigHUKtGHa8fgq9U
rGkpN+0zWV3mUO88kdji7A47W0G0GzLkwrQDtspFJNBLqCCsPAqXw25Z7929iN3KG/NsNpSuGAxN
9pdiBmtZec3vlVu/9reNkMRtw7i09PWaAVrTOmuc0HyyxHZrSsBC6UjRmTAv7KPlyJyqZM+6OK3N
DLqfHo8T+MAMAN5Mfagkp1rM6Wdj32uu8eJYAtJNF3YXTzGfbaIjPk5im1PzuJn/8+EAF+V1oPGG
G2h6EDrUQe4HyI7flLfX6iqzwrGR4GEkf42rxIq4cuCf44jdoJd6xt2nTiQWHxHSJT5GTVHnno2h
FlrpQfY+RetYyd+EGXYjG7txz4m4sjYvuDdNNTfWN7G/pOwi79g0fTgsInRNmKZk4YtT6q5VYtg4
h/TApyr046KxiVyDDF6GE+FSVKfxvXDOqRnMk3cuNinvf9bIMsKQkAKSQ94qSxnNQyvzF5qjeJ5J
rPMlZd1DmmoMHWQgLrCYYHUJop+2yTdLDOi0bJ5nNyZOVFic6RhbF185OWSrsSuna1FXh6KMYCnV
fb6lwx258+GMad83dchfd0FhVj/EF1HdnDsTrU/5mXIumap1P1oP5X8wHXfK0vbFUKOZBpzxYZwb
U6BjaRAVwFajvs4KF606qpYlV30vujO2RDizndWW5MiDORCqwOAr9L9tl7oXl1IFgnTa98bICNWg
bUL50AoxoNQf57UsE8NPt2TOTFhMHbVk+7U2izoO8i3gASn25rlhAs2YtNW6U4X4a82UYJCP4Dmq
sRZunkH/sxcxm/E8xEM1twHuiygOAiKP58hUjSUFI1uxi4IVQAZBLUZCcyG+YLZwL/xQcm+vqsxX
a3lYK9KdezGQgRyboAHPMeXTM+KMKfHWCmxbyRtu0FheaZrIz4e776w8E8l2GDBGKhNW+8AMUzoI
C3U7iUD59YFAW0JQsqXZUfPatoR04G8PjPJ5R0YBTXEFzBr8x6SYYTuBJ+W1Pb92vNBDbsDB413P
d0sy3njr8TL4QX1VbTsBAZLjCathuZLht/mJ2x2JNO1waM3zewLWoRPC+mHRT7/ku7BdHmNC/11i
a1LGk3pDykVrZMQIIdVOyqhk8pwSL8epb13NG8lneik6fQt4RqGjmr65vi7bJ/yZQYHKPTCKYCzn
QJQmmOxrDgCBT10Bu27BSxSOl+sm7m7eYCkHk+9kOpgzrOrNHcxGp7lqdKczx05j++sJ/1R57G+6
l+FRuoRTgAEp3CuxOdctwHsAVckd/T9eP+EKsurdUAU0pNeczHtO0Uz27L+1DyR8Dny7EOOoICZ/
ZGDYAnF7E5YJfVW6ZfkMCgXKwWwhuoBi2mfSD1KpMBZiMLnP0O37o2mJmnSD4UZptaSQVDoJitS8
mRmlUhjRDysFUt5QQLg7qtixFDDDgyJ66EmNfnJev7Lo7Ec0ie4IiT1HSLU62SRP0RM4r6tLbBlZ
/gXFrV3hJxAHOwsNiMlJ/6Amyeont32dEGBeGgGCEsKnMB37oCTzkbg3nneSGzquTKwA1eP1RAkb
4p+bhz0dzQOqRbL0tU/JsSoDFzr99ef8+VFmKFiYD/UHHJzGtTtYjttVCM1DE+pix09d5Sduj2M+
VnSqamhhsmg6XZoe4PtpeRk6IwPq5xvYAPIEOji0n+gspYRfy+ERe0P/5tt8mRkjyH78/6FoRb/Y
DxYxb+sS02pEySdvWE6dgKkJelx53hAsDssr0kKzeMQ+f1TptFtSQlshRcVzUbufCZ3x0fz7EP7c
SUz7b3bwBgg8O38S3u1LWq9VolZD9DNYXtniq/0zOQPvKD7gM+2lKu9G1ejmYyIBlhfDxIrLj1+f
Sz/1CYSV6+kRJ8WtAlT31Vad475RalmgPCWPqkbYDDPRs73yLTcZP+CzbWuHjBMFjGmbmWiTa3pd
WYGQzZqFnbxURsr0U2GxaD5cg8KBjFRBZS4a4xExkDplu8qfMoeAJvWTpYwyJVZBk628+cb08/40
8Zw/xdc3tFcPEux1xJHe2S0p/DdUky1clhQ4evFAlbvpv8vWSaE69AIxOhyhuqiF1PAeP8xY26Lh
IaVBlzjVk+yVV+PaAr4J9p2RDxfJHmSPh/ex9ZO8QwjzISac+Jm38Dr4fjnSZ1Ig1ErkwbQJ+bHL
BGWHNEiEQg6e04KkWy2kVjiGUXhBHiWhKlPPoR9899H2Yk2Tm6XN1IpP6zvpttjvDaGV21Wde1o1
WBoggpekE8yAt2c8vdAKarTPf9tLZDZBd9wA5PCtdhov9YWtie+kJdFv+Vpi0pQv7sOawObbEYDU
joR7LzBEWtsErHq4Cv2O6rSMQ4R1+auzYG6WkmdlRLI3fuEsLYD6ZzBRnVdE9OjiL8cC+1mAR4t9
fKfWK79YZkMq89gJ12GS3JY6S3G2Sdt1Y9Jxe/34+hV+LPeZuKosMnqwMyDbFWLI7oDke6LJJIcx
6yB8X8UjgWGd5c2kYMn3fDO083ZF9t2xq6zqxPy1Eje1SMiQ9oMhoWddNpAWk+ZcfN/gotAydfb+
tfNwaZHjhB2xUOlkeVxA1rBqXz2+x51WknYe2K1Ueiju9T2izvp91bMIjaeGImTMcgNJ+nL7Jyle
B7I2ZGgC0+nAxpoln1GfJpSMU3C+RWTQwzkzuMiFrcKNIESSlXJiu4rViZvfj1fMf+1eppLMwIDg
prk5OW7DPH4Mk7104BBVjOQZioR1K4zCLM8E63HMlg9M8T30BCk8lkhkrokOPhPHnQUHVJMkmbxn
TQlR3U1kaw9Vkul+j37RJlLmN4qkcNPEz4Wqm5x5VUgIiqsq0hDSPbilkHsw1ST0EFq+bKqyYik6
70GgUU2j6PNgKKpyGaN7X4qUMxWnG0xioBIJarpC+g3zJ0gAqigKA6VJ7Z4Tb9W5zPtaQXQxBxLk
cpQ9pyU4NDPFR8y9Q0hqr6CT2U5BdKQWZ43CKbNAryjTZCaYVDJR+pM2d7XQlKy7cAG5rthqGIEs
zAh5Nt8bVWLn1H0aI01ko2axAqnIQfJlQR/COIW2dRtRCELQfR2hFlWbvaKNP/KuYAc/hwROlxq8
z6fZ05Xo8MfaIzdfXZjodjeS+W8FnC+4uYLf3jZaP2mdK4CK2dU18b31TonhAT/MK3i76DSMdYV0
xGhS88wxznVB5ykh4IkZ1ldxlpso0ESA4qQpFBXUJ7gpbQgYpLt9DAwCJWRorEyln+8wJfvMfhD4
WA73zsT6PcbJow4do2pzC0aTP/bIdl4mt6jgIsC5VcnhkjNGY98bgd8CS8WNyH10s3RuIItrCByZ
/qvbIDlmUJ8c3Ot8LBt3ufIiCwE0ZCzng8wzuGP617WyDtjpJIYZbyF6CxaeXlNc7p6EcNDj3z6e
1N+LEP9qeBBhpcB1/tGkDXcTNUUFmh9+q/aglilxtULGFLYJyj9qZ/aaOgLq+fTAyAfjAAJgRWRj
GmevoGcpskDLTY2eq8EqqyAoeMq7HxOXaeRPWRacAfOyMukpDTwqaYccqTp1I/YT9N64g4mWDevS
LD4ECjLQDgxaVYBs2AdsCdlIrXrESGgEvNVKmobKEq0YGZK/1V3HhHm7/UTM49KbGseJWvsZh7mS
eC/PuNtaByidSglBnpEoNto9hHFvy7Zna5ocALn0ZB4t0roMjXnxmoono4qFJkYY5cXQrplTlMdl
sCnuF0lvUcvcwJDuWeD3y/eRINqTgRUb/0zlnR6sqLWSe3A6BJDan3NjDNZAdYDEyHCOkc4Hk6uF
y1NbyVr6WmFRFl94kTl2c7jp14xqfeQEj/70418V4dUr11NMxHO73nLlLYFGB3kPfVMhtSyw2LPE
ZiIblsdrjuHe0poKjN+AyDlMtQygpHdwFPihokcO5lIBYn9+/BpUI3H+PMe04BmPwxLPZmTcjCwG
9hR8BJkUn6Mlw9Vhg/hKGC/7hTG2D4J3FgbT9im1iI1HspYnXgejEx3XZ5x708nZURk1BTSAGzHg
8iv9r/lBEzqEK9cNILGIO6eqXaQZ9mSbKvN0Dd3C85MFWEuPdlfMLaSGpFMeInuWQuoeTtwOOXMz
Yeq+eukrI1hLgIus2Q7usUWekHsO78csVo4tYntzwVaL1vO5frHW/A0aoOvGdOS6rmT7WepmVFOT
UyB6mrTBQw9WLVR/PiijFol1LAPIWP5YXVuN/VgHVbF8cJe3uyQb293psLwTKOOORmWYKYJa/upa
3od4d3dp2rmUj0mTDXxXSYFQf38fFQgttXm08Jfu1xxlHh/FU9Oewm738g0GIRxh05O8Yh/CANBH
/kVE3yjubJwn50mUgIKSoUCeCDuyMChbivpe1jmGcAKMHByf7KG7PT4eTg+1+OvvUePKlY0bk5z3
Vk4tJkdZ4q1EQWDNpRHPOZlwWHAT4vGBzG1WDf8rVkJ7DXNyPigTnwxe+PhXWzG94zdhXVMgZIWj
xpARYsZQdsregudojNFJWQnnoHypZ39v6TkkcVK/AF8BD5GlL+hMqxTwzmfBvZSC0AVg7pxn81NY
8lKO3geFvZemOB+BGrkBCk/odszrNJwNEQ0NPnikt2yYILtvkKjopx+116dGcs+SAiawUxYMb1TN
UnUX06eYfbHoqGfJcg43evhiFx0c+tOjfdP37wmzeQIo6mCnMwhRpQSCVY3cmSKAk0VX5OXpDhwG
zFNS0d0/2AhODQjl+CFAnVsb5Teu8UGP5P2tElxrsvBPJRlAAYMHcEBkqbxYFpiR85YYZ886y6o0
t1KrL+Ms4A1q8BhOqsp/ghFHE+zGr1aOSwPsfNzcN0t7xEX5+RnPXDX1P0yt/l6vhql1k2ZV+OCx
gIwCi4yut747uulwvIjhjSuF4xnTliN2+RhPQLfSp7LrWqWIA7dzAopOLKBkYTLCFFx46XMeqdBO
I6GR+EsKBCMHwz+/cz0NqtepXMQWFwKCGuk5GQ1ovML2FJ1XF9qEgqVq38kQ2DSExodgy+Xl7WtV
8Bd+1Y3sdWiVSu6MrHLOQOy+ekaVB5QMNBM/Y8exnoKNAV9BJKKik+96CpninHzImJ8iT5PHF+qB
kKxivSZAoRz+sEVvoVmOuZrPe0DB0sDIsxA4LLcfGDCDbGJxtYnEJp15k7cjI+sfD1IcXayaPm2b
k/GtVhiFkJp6P8rVD8lEU1qaFt/ICK0+091+2JTCUw6tCta+QfAisU7BjKiEUbJkyx8zaeSkKjNY
CZIEiq2T7bqfUpzm9WVVpvXDLEi8VAhYJMe2GbIKyhamSzSU2JwUwiHBVDF1LQMZqFk0Ql2BsjmB
NJFQ/OjYPqVQSvXCMC6UehcPpXCfnzds7ntaLoq/nv5MiBNsGfu5xf1pZbF2mg+22Xk4pAHa5ORv
iFtjxNCZ13wcbThLGGGvhhMb/q0XZSfyPdQ5sO258xZxnOS61abHEYv8m5zFWHKaig3AJwJsIfgH
o8egZuk8Atp96miiuYMccDj/2A07fI0QRdm9Gr6DMXooaBUgVZYb5nYHGfT8t+BHJbJc0AcX9/RZ
CU1jSs6OT+FXOfnVFsrGwP/UZnuX2jyNPPkHZ6Z3eIorkjfpwopvhoUhwYaeDMh3iENjtG8WqZv9
v13jJNE8RoiTG78dRlcCA6wz4jem9n94qfeTbRzY4ssRNxBz8BNgR+RlIveFgFTSPZXgJLipbQpZ
zkW+pcJYGepiLRvd+aXYvCGM6iEN4xLFZa9LSvOp0Yp5bly5Wr9C4dBOdS9LLrH4tjcTsNEvYkTo
mmd52YVuDeQpGkY6QkpfE72Ie4WRfSA4nQBo/CZ809HBQ4HR9/d3GXZ0+4TG0juBY04Wp6owrmz4
Yp3MRPmIPGeg3iY20uQpId+PlctRyIbovWHvaf47S5JTJoW2k+T2zNgHP1svO/EakkJ4xckYt2FG
NiS5NaHFXFRIG+NmPEYMoH8odCEy3u5ydV9X+wEZy6D0YtI3GG3I3DsfVfotz6WM0CKo+LeTOx53
EWHtA9B1+TYkeH+Yi9Xs8BmoUPEJtexqkd4fqQOeacDHkKgYV3XGiVjRwdY4WgCx0YkBLZKK+niA
q1zizbandpBcSGL4FVVE9l8har6QuBkTp4HyuwXXpoPfFFrJDofnLXRukK7SVNx3uzlHCJZQLaia
imURg6UscroBuxteebKYioKPyJEUQvMT
`protect end_protected

